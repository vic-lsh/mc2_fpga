// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dtPfyjPt25TEv3r0MgWXwNTtmJ9pHdycsH8DKgY5piwSq/2gkkesGq9zHuv5
1Ace7e77io/5pOFg9NfA2bYqI/TmU1D8piSkrtbpvZC5yWXmNUGWM1y8hmfI
TshnwJSqYLONemeQgO9mmAhvoGZWmPwnYwtfO98BUb7kjaniYWu4fL+j6P8J
AAhQ8yj5CKRCRmDU3C51OYCqUgtuUzTqf5nC7JH2sFCqjBS5WuRt3EKkWb2p
OdqHIovPvhKGhxhGPRmNsw1j95f4U1hhwSSVqLaWsK+1U5jppZvm3Kr4cjDc
/0m1dshMzsqxJ3skgBunIdtoiASyAjOsZyWgETurkg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hWPAvw7V8zY8caujzg3718s+6egpASIpKc0dVv0g1KohPBRl3mtz25zX26om
5XczfV99JhS/fsMtIMAV5e4tbVUARf9teo2xz5UvUvfx26gGMzcdf3jhdRij
BtxcoH1l2s4RMKLOzrEYjIMv2BgecVavkf3lTGZcv0aGQIHWJ2sIFMI0HR4v
fSX5wd2NHdUFoOSYeCxg/gmSa+gXMYJwnklqHjKYS30Uz8gVyxtedANSiONN
u3LZ0My5gu0PUEC5UrAW7CIy5gdIbKsd6keaaWK5KsXkDDkgyBBfHEM6w5RO
r7TeGOUAR49Ce5xmOSSVb1TT4nfKTioMN8n+sPImRw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LlTaG1+Iaf+0FmcmPbU3bk0NQpcCgYYrsT/xLbBt1janyNP7Rgin0VEkShgO
orhW2L+2PsKIuAm7KCM06Kw7CtZ2p8pHcpC5W0FZdaiHy1Gbn6/Ln6//ru1Q
yQiiwi+kskrRoqdr9ypQ5ZSZlFoiaf26cEcf9SPVnCAV1+JQSLvdx8XuVefG
bXsm7uXNwkEnEFARCzAUDhvO4JtqtfI1a7558r+N3NYG3MR8YPSP6F+jE8P9
0sWCLRvQemUw0YLZ4jayp6ZhF4XhTgPUj4t6BR2OlzEuGt5YML5nR3+1iteZ
lXW805TtQCrFCwbyd8NRtMDgYGWok4lgDJ32XtXYVg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gwFZg2t4dY4k+J/NvLXZNezq8Eyojg2qx4LiEMmEvZy2YuTKsBFgDjpH17Pc
h8OePrDqOi9dZ9djsDmP5j9cC+cWOGE+u+zl7nKU01DFoRWSTPYmd9Kv1gyo
GhbTg3NApbu8ijqVRLDXtj8OL8p4eqkwazQZVjeHRLhtUZq+T95xHbu5gNAv
xbuQNYCAh87gmS6YlHHlgCBz2CxrWOn/P6xAQr4sHHYHqx6JmsSDQCqHzxg7
0nCG6lgFx/6UGimrrikpri01R+3ap6v5QZDSe3ujY55/r5p6xp7rLyvZ3bXg
slpzlMQKGIT8Ny9stFd7TEN/ybvGU7sIRw2IM6iy/w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PLz5f5KOM3jyryn1H+o2lWomqawscPHyDb2JuzxO5nlZsCd7U4Nm44NPFZu9
lCv9QliGWyVE4a2CI+DeSY5W776RT4rIXqeoV2k8u/s/kwVvMtLx+hADPe8G
GMag+jlgoylNv7ujqGpoNEGpIJudXmNcKAffiyLYiHMqj/Ntshs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
G6cLBEvKt1hBUhU7dACGsDKJ8qHmCOO9KIYrgkkSKbGtbaAQoLPxdlB7z06k
oi6EtoZZGMPjNAD7/S0+z3yEGxvbAZnxzgQKfPBHekHbvKyA2KIqQo1cjZcB
Bj4iqms5OLuSSMbqLApM6+XLYTSFRwqDTqtQhDQl45skDK0hCo5I+G5tpLyd
Y5p687qVBkOVhtwiVsznU7Sy5lCrOo7VgXMt7Llmfc22FX0xwXXlryXEMhWM
a+XDwCqu767rC08SUn4qjgQpSQddiPHQV4kYgaQ45G2PNnzo9GqLTNqo4Ivw
jqsYdWUsaD9eI2sT+6bhpcMvRygdUJbIJJrylERFOxxUGOwW/e6FXiL1ARN4
pnUwagAn50HmKwc5X5eMa/ekltii704/J6fu2Ec5fmC6k/6vbKTv/TiAxAAT
Vt5Q+JlG1AjO8QXgyHyIWY85Vjm+u0C2XNpNDmnZLF5I25kJbWZzs5RXD3ul
8eV3C8zzT9TWBOhqe2cKD5rf9OT2QZAS


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sJt1Sum44rxJ5LksoNw9tBdg9H+zYjQkTB2MhZwwnZFtXf7D6byLYURr/SED
BCph7VPRa41+3Jkg1aZ4v7lYSif2EUH9ggg5OEvJEa0y2SUpR3kFSvwkFT3L
aIMfz/ISU+5XVooijmJu0VvY3XsAq9lVCsYxp/VyowjkiEM+iwE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dZUf4Kf2skV/kR/ZCznS7bbwhwH2zt5nGpjRukBeQOLsvG03Oi5GyqmCZP4t
o6Cd7kOD9u/OSzxmgioX3FrOWuubm9BbYxxBJejn1T20EnHoFEAS6JKAQ9hH
ydGIBAz6jCmeyiLa/vLfvdKZB5JLh297InksGthk4CUZpE40cy8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 14160)
`pragma protect data_block
GsXrMzAWuYt4y9D/N0z/Bv1+Zvs/wIwtq5fMQH415YFR+pc+20xTrJPY2EtQ
uvkhS4dzELmftWCg2D8zFBTj74b4jI0oXMYV31cQ/fQINksA02rN7uDqatG3
xQWABhj/L8daZkVcdFYEO1qbldIEMAG1Tz5toicL7FBiYn04AjYDhYOEoAQW
3icitreNEmh0pGxN3hrMYoO4XMgVocz+2naK7lWzb4qgEeLxa+ZT4B8/I2nT
tQ85Af7/Z9p/it238bfxd25/7ZYEGyAIn5S0jW2zQ+jgtcX20J4zDqDMrVvT
yCmBSw9kN9tOLvP29qZGNYTJa214BbRCJX13shELeXX/nWbdan3cC0YIdGJR
0z5MJzXzVerc9fa6lnSCiZlPtWGbSIs5GS1LmHUlBtkIkK6c41KyqxJWBXYE
+S3RxhpGg5D5nGt58LaTUjMj15QzkPXWBGUY1vKPH1hWHj+f/i+F/H1cp1Y0
A/5ItiqCvOfyxY3/0HV2yU2GBCpb4uyKzOxF5iJbTCyNlw7GzBIXOtcVDsyM
erGRCcVOiOvM2HHrbv5OhglacgQViMqePKKgS2pliSZyCKA4ZdMrugkUzpu4
YpN4qAeRCcDnqXocZcU5po1w9wS7+5X6z5atgigzWW7019Cfif3wgsYs8yeE
/yjs2UzuL4imOMLJh6EDGyrfNCZ7xoqMLvTQdlHqLJmXV8SWKskqFVDecTXO
U0s5wVq1CQRI9rgw1iTTt4Rd7A877bhj6RcOIYgRPSvKJJ1LxG3JZmG32aaT
mB8hOXGuStawltASTt7U6OfvytawZUeCshaYhrWPrMGQiFlquY3sxH3VurNp
uInYd9A2O+pR0+1apMQqoh7hdn3Rd22X/tcJn3gEEqorDW15sbdvBZ/+CS7s
UsSCYkK2Q2Tqq7n9X093OYdptBqF9Vm3wk/k5paF0iyB/8bOtuuztJE8Pucj
6cM97SyCoaZ+iSPWWKLFFUCeoI0Z3q5d9muZZNV1cF4Zf9ogHxDf0KudV0aA
DRnuyObyHUWNmWsBrozzqAPJzzH+o7AsQP2MnfWXQ2IoVtHU7HSJs4nLrN0A
VFVysMor3K0RKULImj5f0gjOCeKIsTyK7Mk5XelE3+jqd9Bdd+3Jb29+ds+s
3KFoZ4IesPygoMe6dgYk0ywsn3JGrnTpuyad0lg+HeOFQKAn1oLrEHnyG0vx
wnwWGfdJ9QcLT1dHGu7KG4hv2jf96hMRjficsFcGqLLfvdgyOp34x4m4GF6n
O9ZEw1ZSBmZoszMY/YFqZ7K0Mp9rVhsI2GmDbVAZha3Tynbio3P4oFooGdji
ExwnPXVNSsvEjVrEEioZbL//+WZD78Dd/fRfuYgVZB7P5r55str0jr5w1X4z
FbVbEyv2jubmmOxywf0w6fCZ0vYo2xpvf48CPkD/IWS+30HBoOUDL4uSHRn1
ujpkQHuBfHriQIjktIFDDmbiR/kIyWiOHnZdqjVX3/cz8vgz6DA2xhqQbvQE
l33WretbCqdKARCFeBGYoep48RbLRHDgws30Q7/xNDlukidbA6QGkZeI0XMn
dm+IBn3JnnC0RiJ+X8wxM+d1nW689E+KRWVHQbp9lugMQynHKvSL31uFMZZ+
Ci9DospT9VPJxuTO/EWfXv+jzgntKJIMLTSgH7D4DcN1F6T7iTYOqube9pqM
w24B5sKZJ+GdGxsg9fCjj/wXCb7nvaBFPN44NlWt9lncX97LXeRxenmwjHdm
JlhWYR+IFolFg1qa3jSD1CHrBi4bNM9A4SjpOdbtECH2+A+zpvBhQx40hz2q
wCAMFysPEgKF5rag6ofbSCvBwreBpuG6PVZQkQkzvFc0fSewELyJUKF69m/n
JhoiSZ0i3OTDHekraJGSrpp2OuXlPdcnBjJvfDs2NznMRZLuYeYFR9chM6q1
UE4jQ2SxztGMxbwkWxSMf/EZlze5w7PbhuNw4ElPhQ2FNXonJDy8iIjrfUW+
OMquvsxGbngzgWtZn0rXgrdPOCDmIhcnIoRVzr0WldzIcyvDwaRrkSRAwoLX
pQdVVqtqW+B0ZVlkhu1CsVccKdUOReQ5OTg05yAXE96ndl3cGVCuDj4Vaqk8
GYfe7Vktspi60aHhXSq3bN7MV9PXoA3bj2Q1SOjNReGFix5PI7zLcnS7UNGB
w9xHXih9EioNl138pR4qharWz4Hk/JF/2DMEuFVU5BRv7If4PwY4BXut4L4d
dnWUUunhtvLrzlAeeekIaMARmUDcqjB78IoG+zdNqkyohIiWUQLNvUWmBjj8
i4PFYA71xZvUaayMCYsXLOQ/YKBXmchkT98QldvysCX7uPSOS9cXtWbAVrdR
4nyWBfd5W9xWz3U+J2onj1L0dDq4zmNfYjkF+TR0ojSxGyXkCm6eMeUdBE8d
CyZgK6ElNIwtwJmXFfZkWFYr6DKFfIYg8ggYX9SEu74BaSdxnECrP1SIbG3W
YBnZiCMARgdflB2/8GI8Cv1wEW3MgAy8JbxBX6aW4l8mCZqeG4kHxAzhyov6
xMhr39SM7QdAw5W80os253vZW/X1CRJhWIwKhJrKbja6vv0FmLwIOovOILr5
yCn8iFmOb7md4oN9wcDWlyMhlbhq+dyGL9YCAFBwkPYWGgf7T2QC8ppNpedh
622CtvwbVs0KAuw9L5uZJaeMgMD1YZB2lUfRit6bA779jW78Ok44FCh2sTMK
1LTpoJu3MydBatBlqENsxXbDLDCA356BPc16qfoarn6ydaxi+hayN9VWODuy
HbpO1QUetRGeGAKDR16TNASx5//D/ZIi+ms5te8UN+yb7CuMn3GhEU0EklfU
YhdC92waVVKIjugpTsszYrZbIs5SVakEHSgfciuXLNCOI7zoXEofQuKYHwOx
sLbtutessq8WejZ4libEyDgE6bKQfNKH77r7tOOgqi+s0KyKEKel2kLaWqMa
RWFK/rvaU5vHHknCoBEFMKNpm5z5a7dpRtxwxHHkz2GmtuRTP+GL8m5evGiL
G6/Qzv8a+65MhgKjIh5L/bwFjAsYX+75YTCIo5jUfOl+5syXFkScXhteF98g
hocv6lEgvMYV4HF17yeFabYIkls9Ggt1t3Qvi/tIySTg0e4PSjGdlVzgPMOI
KihHg+hUumsW+DrdAI7l1u1jsJ0nZ2q4irCol1ahpf5ch1jnmr+6jw3GjfFF
4wb37PT1/22WwDbMj2hYcILpEIIqp+B5TUxgWjZea1JZMUP3xFI/LD7vvoW3
wAGIrslPYD+Bv9GEHjaLuUnf74mnwneI/hKaZ2AYSZjLPL5VA9J3vHKw3Lt5
CKsyIJMpSBTNOGzbwBiwrjb9NZ43LlSKOCyNcOvHGH9hNiJVfQTS10u2WdSl
BkbPiCzA44rG48TW8TABoTHRfO9/Ot97Z46gjaeJc8TWeEIj4WgvWbkwCTDk
cg8HAkEP05cgVb0tEWa7L12VF6kZoBwpOMsvPGY2ujaC1yUeJXZ/N2t7vQf3
JbubodgWprguSrvsdoYwLhc2wUgBuZugOipHYxmCJSs9oAqoE0WlzvlFMkWN
OMWmGSOPXIGeSgcVqPZv4t46AM+2xyrF0EhOa8Y+Th56FYoKoJezS7yNqv2m
+/tf1pIThZhlnanDtZCvrywnlFrOnnnk33gGA+9eLtW4PsneuDX+sKMNvpcu
BXlDGKBvH6g/2e2fWsV4llraC3uBA0r2gmVXMXExjQXarmxT0+KMx77p+fev
B+UJ0uSs2cNQ0tqpm+0eE48NB3sOlahIPhU0NGU72dMf7u3iQpZNWUCkvdsk
Pi9DEotOLGZmfcjJaWhrV1hnJFTEZL8cg/MIRtc8n8ErOeaY5/ivWSq1yg14
LQLqOjyhg+fHpl3MphJjGCuLiXPWi/H7meKSYV5DP3HMfXEHR4kWfVkLWmQp
yG9A9kO9ANGdxSb3Nj7kpmcw3gYKGIGIXdLjaqEILXr7l320t6IGGetKRlup
8aPP7hTKh6O0ONIx7um1rAWWjkFPfRhc3EBRvPB4/PjAXnGOGpMkRy35VxzI
azZZAgIrbK0zlMKVYVpL+FCgteTnTKui+1IIX0iWp2x7nNP5eRoAwcoy7jex
vvZ5I5AKMEMuQKyLLVQMOOp0HV1UqaPFvJNmFw4fopYeQQ1msUpo+tY2riNN
C0P+oA/+kmWrWNu5TNjHhnFPgavxxgISWijCDUs7GaFjsnnUgsfGfi2Wtlr/
UDjCf+ftU0zegnWl4sI3SB7APBC50fqsEHikgGGXY9IY9OXoStDkFEPf0f+F
QzzymOC7Ja36+JGwXov/vTN0+9cH28o33a9wute9NJhKFQlnoxPoRRxNl89v
Y49XroEDy5bd7y8CeLuq/xH0atadFbkUqFE8EnOD4AWnupjWtIBo9oPXzuQW
O5JOxJBVqK4Jj3rKL9N+u8Bbq3spyouPs7EwZpT8m0VDdiergRmr9ffn882r
rjF7sAhZMaM4I0AErRM2W2p3W/eogKMVcxT7L5rP4fg2FhmbqHGf97MkmTqC
VC9CkCKj1rM5EuZ2mwAIeovC5VYWQXuX3S62QPJ37Q1zlw8ljLUw3GjOXb9z
9PLt0gwMqqsQV5Vl1eVWn+JZucOQEFhcWAlrWbiVgBsFIx/A930CKDQk41I2
dWOKxPgIoXvUf0WGrRtYvPhcQ2cETQCd9pXz8ZBuJlEsTebBQNcjnByj7Hbi
3r9qyhWJ64N//Nrthp42HigGMkDMuadW5QJV6DSlwUVyKZ0erjbp/T3r+yeP
+JB9/dBk28yLwjjcOyypQiZgQutEOMlzURIpaq+uhB7CgfPZ9u+wnyNW3hjG
z7cg6hcprAvvVX7fyRcjiMzXLE0XbWlbvZUSBn4Tvh4xuPUSKwNocj/M0FVh
UijdeoJPoDpONNi5VwQNnnukCdEdQpepSVawgF9T25tSZU9RgslCAfk2Cex8
0lSQ6d04SpMFRMBX5SQRnAXlm5fsUBn1xwEFZcYbQSfCAxGYgT+5gbDiYoKQ
RDM9cMgS0NqFnkaRWtbFYw0aBBsSZBgbyHOEZLLuEUwHBpRSFCl1+pGkW+XK
VjRhQcsIJChiZWoKI32OAWssxr4IpB71/dW/65y0OvCeFemz5+ctLtU+FA8F
jIM4SeW5FtDFqizJiTUGhgrx6YeIA/8oLi9lV9cjjetVDWD+rbeGful2c0eW
amRBxweyBxIkNugLctgwvkI4A4H0k+p9vjoR6ibpXZYsGHxriQ9TRMuglhYa
dIrsRuWq10Uz3dYfJ3Jbb2LcC0QNdZUcPsqi1XWP3OieIvL9boVhmly60r3R
Wq9oG0UWQDbOACFBkehad65NJ90VaSsQDkq6aSknyL88GX4YCWy2gY1KN+5c
aX7JEyGXSLfU5Uo87zl4MQLcNyowWxM3LML9geEx3Jehq/GGBo9sHHs/HMuI
uGyreLjpMsNIkMwXw+QJvbdCrw+HHC6/TwoWnRvaz78H2LaPeM23yclrtUsX
HPYtd6qikV4Y7EBHGVd/1s3DUwKQyj+LGIiS8cfoaEj2K/MgFlDZR3jnDwei
GJabIhJU/z5atVH9PQ4uv3V3vp7ZZlm3dnoNROx8Ksn11nQwkNzh0z4nT3U3
RZmoGEUBS5fIdxJxRXZVCvo50iLr17Pm5ehXCocorE2wz2UzBE/0oL2Pj65m
XmLQms0mJ7LKzurCnRu9pEZn925D8i2rEO4UXdICewxVV8urfdACgK+NKM+i
aSA6/KbjwbHZORzJCoqiB7Mem9hcMHjicNRm5UGt/utrYUIWdXapdGFP4Rt3
OGscRad6Yu1PIM0yJmjhgHYYwbeb+g9hLP+qZbTgRgoG6m5J5ubBxyKz8M6E
UzgSOkxQxtS/GIdfrUsDWmGGUaCTdtynMxN4Q+YL81LzGOcAcsj+M1nWkLRs
af3MKtgx6Fjpx4HVg1tSpQjIsGzMfVpzpm4JGBvUju7m78Ry8ZMhzUWc/wSu
3jd731k76hzSpb31gfsWda7iO89PeiEHkK3lhJ2w3++FSqZtRyQxxqGPx17z
RfURUNWsihJfpMff6KQnuzJS+wVKKJoS1QskUPalYX77ct1bLFZG77h2/Ffh
rDlCbuNtmP6wsM2bTVHLCgDjvZRw2ZcoRq6bq0LKehhM7ojctpIK5bZAaSQg
S4X+jYtimLeHnmM0EhXRCpS5zlsjn3MWpT7mSlyb68Di3QQmeJo9PJOOnebc
IfcLl6n3wqCbINKz24EpmuMUzLx5jV1w60ZdIVyF8ef2fuCxKAVS8aXNrEHC
qq0qYAFXT0buWvzXbl3WxRFTt94eEj0JWPPgZ2oXG9oa10kKHkh432ot86j6
Hx7KTXVfSHTtGEOKrlIDpA6bUeSNfQrRHi4U/iMCcNSY4isdTMDAIq7DIawu
RC7lwRVL2ngmgc5Q7uLrhYuvmJxh+XHhBaO5IC8dT1txjLTmeBPtWI//wUlI
FiEHVoVxo4HtZe0mosjoiIpl/asZAZj88OtIe5Rc9OARrfPLwnGHChMDzzPm
tklySgU/7GJWFSXlnbf+/FSMnb2lR1/jxKrpayG3IvWFH0IOmSJFTrK5dXNt
IdM53jDd8e5LJbCMy2XZ5DvPYzBR7nr4QTuz6oIgQ6KUlUs4PwBXRTvOHwHv
p4qmI6k2rP76wqoHPgFuTkO3qhIgX/ooD2ex0mw2CXRvk+EzKnWeJ9GhC9XO
VaHnuY2d90BGvltVqEvII4a++/X8rvEy9QKTuVrApCtqFKLpAXvvF7GOcuFh
63JMFV2HjINhBGFVDymJLSztPzAsv45LHEBYu2RnGLwh2nebcOp112NfjTD9
tvB4INLrGzidn7aMxWcpPofz0uAgQ0lrguSfpyufrgNQkGq0A67ccizRN8mz
FbAnjcmT3OAF6IwvnDknOF4HDhNsxkYruPDEjaxL5Yqj/vnwVkj9bkkr+xH0
cNZ7/uk4PQIb75jqFYVYYdMQD6Ub9SuPHhmHlgXP6Nun96qaLGjQhe6cymUd
Jc8u+Jy900J2cIFpJPQQFdZvPOH+L8d5sPCcMg54e7rnxB8U5A6GveuAXx5f
RXQT/DfG41EG2skqIH68DEw66fnoNwJploX0eAgrit23NYj98b/vHd+5rWGL
y5cIliuyc+ln9p8SFgYWTemug08/Li4c5eivQewNcpJyvQbo9pPWBm5L4Pa1
FYIlR05rr43yrkAWa2tkb9l9qahaAng8AT49FwWBv4lSBVF8ATRKzkugHhiW
LMh4+RIJtVJ1w/qwA74M8mMy7Y6bnVegnT22OWLeVWzJjlRSUIPL4s4HeZIM
7Z8MLXOTs+TausKJROFi4vxEm1mCxAGMR9YYZtxZ0bBwaJwQ0BzW+nEmxKJF
DnNRV1M6kCISIefPM57b+1ClKSIrEr036wVxx+nQOBDyEbV5/hU/OHQatpuf
y8TfTFF1JRq0yg0WqgdZjHYQLDk1CQw1V+nAwqXQZvpvY0enHA/4t7rKOXuD
foXsnA892QWwa+iMPhqaxkgTqLpbdmym2eeF/Jd6fe/x9yv9yDWY+X9RsV5R
WL+u5g5xmtSnpQ1f7t0bY28Izo/8cpKVavmMLyLCNTUXhkMn9pN3bveEqsQw
1ic8YIW9WPeJqaK9McisluLtGhct5ycFc6nQI+ev12374krw7RXXm+pfqF6o
j/eJKrysz7QWgRkI+oE5+7n1057gvN1niD0XHJmXfeSiXuTtkxUGI+ieFIf3
r4NkByf8mXHfc/M3haHlfQKVBKTKGmuQw7n+FfBw6sXuuWjoO6ofg92EK6Q5
sqBoKYMOcU1+aEZU2nFc7atcaIJK93iDh6j1MJwQr8vBZym42dunjOFudlqx
MVe9MqOlHQuHSBnOvFtkTCX9/RnlDvXj/dEzA1g13+YnFAhpb87VfEw+BTlr
8GizdoJ5mjqGqqIvgBk07+59wQjv2STBZ6Vu0A7s0038pHOBUFGJ6WVOsG4c
jRat7bRWeJegIUPE/IJSWkIpSoEEowfLQ7eOYCrIru97IX3gNw25Gm9RFb8p
R82ilLS8PzYBOim4rc4+89mBUEevHbvOaAwjuCHLgwTLiHJZkDXtTWsQVj6T
fxq/QFmKYIu93Yz4vcPYfpz2XVTJTRkUWjJ+zSpuH+XmVZ6UYPRXO4AY9A+W
q2+l7iZOaKg0NUt5MvtssOe2KtrPmUaGras4MuSOSRJEkN1luMOeIpWpe5B/
GQtMzISL9R6kC7rWwh7DoUr1U+4PXjKWb5nxvJAeoQvpeChl+NOLBQN/rpO8
N/vVBEXZQrXkam4FPaHaAFY0Xq09LN9P1Kg+9aXUnXNiO6kYSLo43r49m9Ag
eO7wnxvqQ3KCqIdz5rRv83y+RWx9ZHjPzSbCI08j6GThtglIHIbDaG9WJHdh
XfHCiVk8u6r0WjI8dLnB8m93U/oTYaKVrM6hyhN/4mxDm8tNDkUGUhjO59/Z
pORSaB5MbVOeJRW196ndTiy3KPOzXrOUT/dhOoTAmoYYMDK9cobnYFwtx7Wy
VkfyZjO/Fi/uTlZIs/6VC73PHw5ii2plUfcMibX1vg7DD69teVftSyfwxJOu
nSs2F8y2eCZqq/wO6wFzhIFQ4itQ/dLh5TtogEE3QLgViQ8alOFL4mZhUhX/
06Zr0h9b4vnbz5DbhlaU38WOX5DqL7DgLDS65wPraUIyA08cXtaxJRiFsLMz
d6GvmBZsgtqSuIlUG/w5wuK2K4RrgdFAHXqbeZG9ZMuiO5WwoDq/rgleUXgu
E1PxlUUqCfaUy2oybgeivyj3jehDHbqxT5xgxzssGHhb6zDDWo7UAIq+8TUr
s022e12T/IP2eDB1kEA1iCmzm4dZNNo3VGP1NV2GUzkKeavbeBsE+3/qhhN/
x/ce94d0Smu7WW+y8UcZYKYoxkvyNzKTz+Hnwb90GSUFfmqVufHTxODbNFpF
UGXR+7lz1RGEXfETD00VLgwgOqfGFLEGd9AOKjTICXxGWv+1Hvkj9zLhrNxY
c7/34s3EgPOOQ5we7OMBrvaKUJPB0/yai53IYodTsMYnvmgRCmShd3M3jigQ
6R01E/uiuqK3ONToO063XOw7O7w1hJwoxMihBvf2alRcOvc6AO6Y2P22vbWL
t/63KDYlfaC4Q6hA0uC1fd245VV2BiAA9hRcdLp3Qea0sPSnfPAyMC40N2UC
HOsfsYv/7YC0zH2XOqev0RDmJaPefhUv+BQ1rfbt+HnbfxaAaKa8f8sZtKyY
382fsAeI83dSGlesWMs1QhAXj/UqZWpK7h/14aFgU9nZ8BDN36xquJHp9zNG
6PKm3E6zgX683fFYecub+xJ/D46LmYSESSuk3BQ8IBCF6CdYFavr4vz81HCs
UDw5hmnp3PMuP+4CZLHsNjLj+cZbnTQ4tCKi5hk5SBmTcH148LgJMrKXdc6T
eogy8efityt7wy+ThTOFXkwh2e2PILl6cKv+SqUeurTS/8zqJnzFdzRlbSGV
i6KnRHrzKmH3lWZG9yV7Es1av9U1HMy9eCXBgh0Zl3aiHle7AW1IeDpgvK2R
7w/XDFy8bjSpdGwVR/XwVu7aSNs/k5vM2Y5mChAS2YnlzehvMLz3IiJRz5VH
u9vfQFtN7tZk+8h3F+s+pYOC7iBWW8oIFPEp+w5Pg1YdQ4TPP82DrBH8yXtX
5i2dGFZ4YLYRxgtQ8De4R1hhXS3h1uTyk3V5yx3rp1UrrvzRFvIVIazatfZ5
+bZyTyho826HJRIJKAczwmZohGMmijEiUjBxN6Mdcc5KsPuczNY9T1JacwCx
AqBRxVAhe7ZmR4hh16to6sZTan4a+EjCK13O10NAgH8rDGJ8GZAftFuGuQqg
jpm76Rq9gXlPT6dcl/Me58/401YWjw1IBLzkST0hp42p3udgFPU7BgoXD+Qj
ylDBPuyIwkVhKUY5vI15nYw8+bQHzk+KS6RPgankrZtEmfUdeTDnXiGH3ufy
TdVDPno78ZK63CIFQXf5Bt25v3TBQirqkI0/cez7dGPncx9FI+sS6HnZixbv
k4Uqb8k4dlU++N63jQdgKUjiKVEqOFW4EoJ1MXatb6HJYCyymeOrTUhEzD04
HA8px81uymbTn2n5WQK4HdTsJmzQF4bwTSz5Rw8IX9f2cTYekHpWA3haCp0h
svpsEufEzxtnvOjSq8QwUhVbCySr1WqJDQTvAcTNtNXk7ahtYcBGG4L4xKt2
EukVCT/YGWTSxw1uFhikkLg6sXOygU9m9EIJUH1ivmsmzQtR7CfZOWwn9liL
HgHHn0SaPSA6X1t1IRvIpzVqC8qknx1EKPdwwxgXGfz99W2GWKV+/Y/U/c5C
ou62P2uC2St1QCUR9ULJYZgzt4GkVn1I85BxsmkY02FhSrgzbFvStWWRAx1I
/nKBh80z1jFiKHwM0OGGeCiLmihtgfYB3iWMyj1qw59/fyoJ1wnNUYgAjmij
RL39/+i/NY9SyTR7+O0ZPnQN2GxrW3txRCIrjatXkgyJu1wLfBI1hv4CtVWa
a9I6mbsNAA0HcumLL7SK49venVB2TXGHRshzZpbuPGrXhxtGfEC2Y7o6BxmE
s0qnlpT057DMSK3AIksVJuNRszNNHjw3uD93DJhMepNMM28Fnf3QaeaPaAjO
DsJkIHtaAz87uYqMULSabsi4nkj8mKtxHQdS7p0fEOrHLBqCaJ8kkSaR3JcU
vU3UJ9myvYjoopca8Z1gLMoYOkCVEJrXX/ZvJySh0+qXwMbn68AZp6FfVmfx
C7CIAXI9BXW/YY57JuAmr2dchEAjswrkAZLjJUqUjkwsjhyIndKSPOqPLf6X
fdvpUQJTCorX2KWbj9kRrb/7j+eBZotowccgxr9V2ylUzkni8p+RRIpuy6Jf
UkP8JdF+GBtsjEgnxn0340o+ZFrlhtycn7rBLV95bO4WKufPC4Gf0mKgZDwW
yqKuBoL3a7lQtRfHkbFh0P3N953x2PpoK+A8osUvClVQM1srAWKMYES5qIPy
imKzEHPznOnm1v4eHssUCrfqt4oXsM8CbH/jRMEF02PIfDs95j1fVHX4Axcl
ahAWHBCpkHL1PhCmS8nyHieu/xvWbbH0sfzJ4oehfnRnaP0sQwCtuRU2Se2p
4iUlfKlcMhCUTkRTWBoyerIuLHqrNzMB2Y176WoQviWdeKb/j1qUwgyTmPJ5
SZBBjDCxZ9kE/sJxvGek/2HVVU7VQmjPedj5gbmGrHJ4r4VFkFikMZJP4wcv
9027d57kV/tOS0fB7+iDFHx17SFzOlAMNWBB0cHGwIyN8kni2EUJjXU6jmr1
RB7uWAo4WRa9MOakEN924IR/qwgwbzHRNfh62hhEgYpY75k95IDlM56FEMwb
ggyyjuwRco7GPmknoOZUY7WUsDiv2d2xzNHxYj1HRTopAy/faqALAB7a11yu
05OcW4mOwqbX1xzFEpt14dYORyYG7yKrFT24VWUnLarCzIhTeTxD+t68G/ZN
e40lSXARpzPA91GbJO5plrj5LChFp6rz6xPTUbAMxJ1cgaWFNX4AuqsGH56R
oVwmG+TZ0qolSqkYYZQgrGAqyrzqBWO5MBXrMCZD4zjNQ/IdqIolo4tdlAvZ
4VcNByRRr2Sha3ZDR3f+zu0ThNy699CMbqVH5m15S6uneZdpXnILL8Hu7XTp
9qHSOALiF62BJn82068121A0eejr0L3OlhVpPMgzNHH4QfiIBVL6j/eF1gba
5UrmaDJUfGGesPI0thiLVKkw9uCsDflsDc9D8DVAUEAG2eYxP60bFhihip0t
gIZlARi7kdqQemguCJQBUFI2eLp9JpYmyHs/sAV1V6cko0/qHyTM3p4D9jie
ed9LHuf34XEdFavB++p4uXJTAOl1VQ+MYW04MQEWPEZNs51hTy1UJyOilSfO
VTx68OjYcfTJIPRJdAGhJjyhEHOG5oJUtvUnUE3neuxi8/ueImRS0qDFzAaf
c8gAOuMFuCFnGng5B/3uNwDlg6LmsG4k7DfnYJB/ldZU19+7ackGWR+vW8Lu
ytlavplDqtmVH+aqQKB6z8GSspqBgBe7aEgxMTbsfOJ0auKscLaNzhnn3tCG
RlhOtbwSRtpWJYuySKNU460QwQte3+CTipzly1sTBXaE0RjUANvMUzAwSaUp
9jSR3IMFBjSqpxCGLGCwLqBRaCvmwzxE9/A3Pv7elvwo6rG2wnY10BsExJM7
kfBiNabWCMBKq5/4qB4EPgUxeCCD2PSYI5oLMssVP3jzVDEfzI1qgf6vVZgk
2eBHREtBcWZrq1AGWCDGp3bvhHxdOzPJLZkbdVHFHCTtjCiE60qQFEzeN/E8
m4zYteOUIfC2o4gxEwglu3sKi4/jaM3w67f5o0Yw7KyY9FWVilQ+4vCxEuh2
uNzIbBfLmROIlsxLaztfrdeLUjL5ytnIJjvPX+s0Fi5euYLxzSSs6FWC5hfD
X5nLzuoAfefF5xLWVuMI2gGbXsSt0GvFPNxLfCwgIG9TiWxhV5Rhl1iiXjlx
cXtan3mqm4fOO31dkrMeneVzXx/FN2hhFFE93RDgFk+NVm2oSnvVMd4m2wwT
iEfe6uuNDR0p871DnhfGeCLnfhrVnKCBYgBgM2xvzS5/kyb4dG7V8qGGTL+w
W5VwS8CwlEuGWhr+DqQRdAl1PmRcQxeEEy5Jyh/6XmiB9T79KnBWU1EY4Fog
JBVP76x4X/WCpKq1xIfnaIgIw0jWv0vLpBF2K/E9XyEuIfjOhJDb1az92yv9
axU1pPefj6Seq37mAV5FK0GuujEq/RNspAIrtRFf1i1XkC+yBkuGxc3evNAw
rMHxpg7TGjRU6kxBSJlgPssHvzHGAGbLsGhyTWlB1cWBRJkV9jhf+/pev2le
exK8GvY4cLuz0Oa0WrRwdcqcLXu3052d0QJkiBKLKDbu/Jcw4oMI3diEKdpd
dUtjdv8cF4LQ6MboALt5G9+ZEWNQ14m8LJAHmSXr4OTfqyVckI6P3U+PGbNL
zTHWBkQ2cdroPZQwiRkoToivG352X/ezu6ZSbImRRWQMylrIeorbfNpgejte
WNXmc+VoFojYtPG9LM95L1d+jWG7wuK3sQDW3AAN26JdIcz5ZTD7gj2RjuyB
bvWr9skd2kgAB8P+nQbdfra9XMzteGpF03zGj1MkRyB/SVCLGgDjMIisVyvp
n5hrt5aPc8KhcoqHNrkt9z/P4V8L5F8+YFM4YBgZP9VUZlbXYJgP5r+QANbW
BGLEdPxBtS2CVty6JnUbWYkKvS5sMVTInwvqeWrwNGsecv3BU8bp6QhdOCSP
AqtRxX8GSDuLWFWB3jux1bVjLojQRtWZz6V0yUVFCpBpxkWgBMNEu39IbOo7
hCTeClQQLH9sy12CNreU2KdnnaaYHRwK+z8yURt4SN5yix5i4pDco14sYa3V
Ihz7/WcAVehccPTozOaR3B2H5N2lXhrqIwnFTkPmg5aa8BHdijMedYnuzYpj
DWb+REcFPgBjf4mvN29jgDOVE4YYOh4n4o3+sCaSJG3YBVJaSrhdVLY5MeYT
15tYpU/Rh3XNPGw3R6r4MtLgc8ZQ36LlkAxne6Liubv36solwKknas5DOuy4
5Op6zWpLf5jJFwkQEBTpNJ69kaZi2IcRXn5Z9vxNMuNuZHG7uk14aKIkkbEL
rziLU67+s33H13tK3oOGojt7Vgf/fzwT2pacRjN4qZRssZ6JrHo9f9Ylccqs
v7wy5lpA8tsDhA84xySRRUxK6vaMxS4XAwps2msGDSYdO/9AxnlkjyST/xS5
0KRkPTWDb1GFZr1irTeXSZiR0QgBv18SBJPaJzwekzrODrLW5Tc10JW6mcXE
YMbnyAgzVT23Fp9sH8KPnWPwW+dh5z/O9dum22WV5pu0Ho7NxvzpeL7Y2URi
KxyMgdaxpO5TK9J2iDCh+IN+YGP7ZH9rydSkpY/9AZaxajTeABrCFyzkbPoz
ejXH9xyNGkHu4d6szIr49KmsDKAXGC/fXzZEoQHMVRkG1fCNUzqXG/+t79Eb
a8NWJoCqjsbyRmhGO0f/G9uLGSCMjyrMDdRVbVHcLqLUnYfnzTsSXdYEwgfO
eu/9bPdvq16xeknWwtHBniFPHJE/8BOmgrgYn3iwNBgwjmOrcebMrbyBHkLy
U4julvfvtzi9Xc8ugNCUwX6G0gZ71g3c0ze6b+gl+lGqmJnBtRBP2fl6EMPN
8NRoWYTUoD8f4hoLwWEywjgwdaV6nve0UJi0zQqwgPLd3HFcf/ZiYWS/fJ0k
keHMOuHUBWZC8cEdfCWYgm1vlqxZcaxiI0mGBxx2KKnam9q7SWjxAIeay+6Z
DrB/CJLmYR2OpJwMM9G7P05/0q5zPATzVdffHnzHOrdkFwK91PZ4sP97OgBJ
g2nkyvXYJbl/zsTQkdyaxRo6DD0Qs0IHIeW1qVV+Agp3ZMyLqlBI17CZgIjL
cIlfeqhd/AFY6fwYS4T3Zb0dJQ5RZiz54jyN3K4p3RETUEHWMbLxZGgKaqoM
BUq84mKtiARnDLESVkIu4eedikuzWTS65EDFxfruGW4sLigE/AEOA73A4Ncm
xAW4LiF6/irwF1ZZ2qIHVEXWvE5OZAqWuD4fj2psoOtH6d7ZdXp0UiTj4nfK
+ySjiK6RFGBvb0MwGh/9Bay9r61vAGlvkLvnfmWoz7kjeNXA4VUq+nxvtAU+
+aL3QNSCznA0AYKiLmtuunLpkYl1G+QyOq20ED6qqSZ/1LrRBg0kN5m7stNE
9iCd9+pep02HfgPCVOcYqRdpwuzWxmowHiOQ//bUX6WS+XTw1aHAWUN6r8/+
EyNcBTt+EIMilmf9ysr8qulV76PD9pUuEcizdSBLVpGveND2gmp+ywR3g7a/
wRwk4k+f19hwZS4D+I7kMrXSLEHlN38edpVGt1PXVlG78iTrccKOPrV95wih
vWOP6kU/CchT8px6BcbhqGDn3UKGDtM3RLehZzKjTqCcofVZ/wZQMgH+5xC6
wqyITp+Y+G9sobqNBxD30k1q1Io3OXbFIS1Jonz/Ujp2TxljnDN0eA8kFhZ0
ZcjtHeqU/30A9yNRyBOl79ztye9B3fhYSB5DY0vE+HgjR7OnsVSBYvmtSDug
ftKciYjbhOoXJWG23EKICyPzEE8Fpdm31Pq6rUh9ZGlfa/e77QpP46wocbm3
cPrKcHMm87tgK6j49eAL5D/CBXS6kMenaUdAoa+WG5mVcLfrNPXMY1vhYmW6
4XiLKWUjzAkWpPMlvDpSwEOa52eRrn7Jt1Jwelm8gh+B2DvuaT8vVC9kYaqG
td5/UVk9/1EAoK62pVg8Inw3S983iN3ibfdybSnTIf4N+kfASnjzIKToLEmu
qng/fk07TRsZU1pqkyejLolxlUCrPcjo3qMjto2kWYQ0jjkhsYw1RgA7qCI/
uaXgwGWOzfNohW1inctH2VGsEB/I779+i2TqVjp8NK/MV41lHbH9UtSighdf
rOEj47an0uZ/3UXtowRQuyF5InerFohgMTrsfqu5G1FKwkWucB73CIKzthUI
1OrOySH6sZ1XxVhdmLX6Wanh+a79XpJ2QP79GmiZqbIKeI/px5+jy5WoUpcT
D1GAfrdLglsp9Ez98JWoBkR0wXDfmaVL1KhU173EaBopYW7bhdc6nCLzHXql
G4X6qmyztFApvVQPoPM9HHgBg4d2QlsACYufE03WudC0EGY77jzbOug79spo
BJtzr22q6TtbpxXc7X6I2X650uLi5E8+V7iEf1hQ75hEr5PWa5dC4ehL33HL
FxliB6efZenBTMXyoHU5xMNvXqhoq8rZlvTN0eK1rXE7gPv1ath0iUKYLaXa
yQQvFgKn1NJg5E19zp6kSAbnXLMK2VtEL2NptYKgHAIDb6s11+1J3CZKAzLm
fZPZT5dqyElWQ0Oh9ouRk6sIF4wI3cqUl8Yz7tMdAE/XBAly66cfoZVCy36B
Bxfx1BvKKQKVVqoTozp4ASJkgdH7Rpk4jWaaLw0vrU31fcRJf733d7yoPXrv
VO+1qzuAmR9DuYg90/nd9NuRHeDVIKWg4bc65aqszYKwiqqX6PYGZV/Hn/HN
S/9Eh0vA4d+hZ+82fE7uL5z8qmR1fqBFJuaeW1KBXq/4iYAL9UobFGwzcrla
xN1W339q+9Sx7h+I1jG1Ad27cn+XGc2TtwxKe4LQjLHADoLFuoUhK5zZ7Hwi
+zoTBpvKgqVNlHsCjadbKA4YU2lLYW+LkGnYpJhC+I046noQ+3DW6dYGE/3c
WiAWx2B80MozQWdaJMsaatnktLdPNg4q7YNo2zZUd9TQLxTMjyZR4xDmnWHJ
Vtkz3JL3W1d2qprwTeMZWo/BZTtlCBdG204/jEkHEXDn/bhhFofbG+2U/c5+
y58HdaLWotL9vcEb6ItBmv87cRaBf9zSTIrj+bRtQDk5ZCb5ytlfMyCVayXj
e1CiN2zQBxbJs+6otf5vqpEHF702lNvUk2lTdEeBvWK92qF1XsmOhAdvEZBY
0v1Ey7Yhry1Yp1+1BuB6CuEzY/vhARIzXfxmCGcbFrgeRtTzLr+qix+KCEFr
GOB0DQxernH+5XWfHtd8Xjv6TSrxAmxhAvdkY8FtaMywj60dj9Urq7ztA3oK
OEl3d3CItFl2+S5sGKxfGBHyS/Q+c1i3yUf/yvYUclEskxslCUf4+ri6s1tO
p4O6xsyDuN9g00WIbwpUtnpz1IZ6hKPynDrZwuO/57f15uX5LqZerwo7JjWO
FvPPrKBqZknjwAVEd7f+v1QJUTNc3td8fKqe4lb37kHdeFr+VvLUIM7Ku1/L
uq5jbC5agx85dXsN7dZc+JBniWSb/lO5jaOyYVjpw8xz1dR8Mj0ShJSuf0NY
F1iEqvxHPLWc9SW/WEzeCpUp0FacEG4hGJhycdyBcfUXphyBsBk/iSf5SUbJ
9LdKLF/WXHUD1dOAa/KqwBR+elKuSl0PTeqPIYzaGH0yILApkfX1rqPu9XVm
oC1QS49MJz2aK2NH+gIlCmGhHrXHw9B2y3rzq7nkEk9PyHLxvR9vvizTvlW7
G/Er9L+cpnAxH2h6ZTEPNc1y77Z15CYfmhuBZYxUYL803CNYZI1fA5HKzWv+
QlDPrFRL1E4ZkajP7hXThNZOt4XG3SkbrxqvuPpAMVGVL0vw9R2RIjgny1d4
RYkmmodhP/5JgPIs0RdxI0ddEq0Rj9XaVtc9gNpg+WEu1Yk2wBjcNW2CeLQy
8qts8AxbJM1D3jm240R0FrLnTx52h1siWHVKYntlDq87xwRLHa0UeXTrdjAS
nd3rLFMQoplJakKqRJtPpNYTQUdjf5peVcEQiUssyE0682kjZp9A+XN6dFpS
VdRegxHkYUGEbHcv2/Xr+hp8wSuZEjH+N8SoUmKgNe1Jco9rh8rwL+BJ3zAY
xhsH21oBaKOhOA49ZjtvGgNeLL9m1Oq1Yd1J5GkKnl7eMoF2v+Ij3rwi6LD7
mCynz7Y0pHxQEjy43W7m84KnzvDk/ewNRPhk/s7kX9rixy7ey014qXkicGam
hGoT1JV+2gl9N7NsWIDwgmc4/ZDl0NJkT5jRhl50TKlbSPnorx+07D8Ghsaz
UwT+zUWQOzz9dVaxIo2NvJD+r8GhsBUfNBddRuZUYlZons6PEtfRCiM9qYa9
dYVoQOTZoem+rLzh2u6lHx9olPF0tmTu1GIkT5s0bo/Hl06mOQ57lJwzhCxj
JnJ72lAynpndp+MDa2MsTB9ddBUNPoZgTGllI+L+XuoASI1faLwTiOUcAOTY
60LCMSwE07Pzf6KCIsmleoaGiqSRexzYX7gpG5z6FM0OMSFPT7VMBNFlT2hF
3GR/v72CzKydtCChpyLfpJnAg7sL/8Q73TrdYblFqRgWpm9jDsImwxgatdcs
WSBFb9g8bFVZBd7dNYuFwG0paGx2FF6cd2ljbOT+GmUWjruIkw0EQgVQKnUW
mHOdJjRNsYgQ9NYaSoGcwWRtBltX5Jo+Ei0OIOZ2RRPcXIVvAEXFQWZ5+46E
yQev7Y97JWO1zJ1zF5hk+tvgCzeMqUH+ZgraRm30kry5vCTDqGmFtwWCx7Ip
z2Je+DP0WLCNgC9LO2RfQU6jNW3K0AkISQDSmU3cSssRC0rbTY1AMqPrRqwa
7faBaj4NNrYinWI+EafhvioXFrmaKToD1e1nTh/HXjtaeqa88zY5qnTdGuw1
RP9HjdTXef7H4GeoXAjW1b9Jqg5zMLYIKLc7VCbGlNPqK++KSyDHH4OHwIbW
j6WrmB1e+oi4+pFFyBlvUqNdjC9c6zph5NyDVy9C7JJJcMZO7aoHFNpLQ25n
ufmgv4GiPDOI6sZYAF6FJTY2BvBzqDpQwYzY9aDKPDf4JtPznAiHfuiVI2E5
pexabPUvUNv9abQ0TRu+QkbKjbQODMDxiw/tmJOYlRNjhf6/kwM/G74wLgjf
m+FUVBMLqR4SdNabBKtN6AAGYeU2IGqfzUVgjKiKlqugpTYtCINVcaMvsgv1
7lJrx9Nv7AC9PCfQ36LJ2W1mqmeEYqDiNOL6dgGWcNbhIKADPkMNLbyO8qBz
LpLGfCNfw6jBqFkmKEjhmV4xh+L+HP3dTdpedGm6l2aPP8OMkG6sK1s10VgB
FhAKK9OBAVUJ9JJGipokiwivGZm0JK79Aq6Tv4Prv4QWILCZV1o2QvXgPgWH
5xJnVOwLE2mCDjGVOkWEXcKBrDed1d6E0FOnD5T1df5aEtEB3OR3zgzEw2ZG
U7VeruVwXD0Ffc6Kg4ViaZyUT6eEMrI3vs1UMH3s0mIOG3Ck899M8tNRr0Op
v4pkNQSzFUCQWhud97OFJrlPvxRIWDTtumt7CwXWk+1YHXflr8ILC1VCViTQ
dVWFcTjuJcgv8/8umJXw5x4APqzaU0Wt1r9VZlvMpGYn7pG943sYt3nH0GDh
0ELv0PV+ln0zA30yUT1HcwOnh32Zt4vpD7nSFJ8fxhEIrZxPr2GqH+IEGfpC
7JLgMtNsYusRkHTzF/XiFHx+NI4nu6U8911oLahp

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Kttctzi5aPKQ6vg9w+1g45z6Da0UaxXtt50QPmQzmLiVao+5Qg/yS2eSRK3c1uFoxS+G6ngDcAKHm0LGGibx4soakCOjaaRTqJmqblCXBo4qigRRJU5sOpNJWGKfxZC9LZLfFjqN04HCQ8ah5FN3P2yNU1iObRgi2dEkx758LbIsGmsSUmn36d6MTHQGWCnH/AC+2pgOY84Iul0q5eg7DNO6RSxNOih+2JmnF8szbMNUemBxaEM+nA8C92x8Fhdrhj7lN8yZGfSGowOnvm/NUUE4g4NRwkEfNGQ+dQe7YHoVQUykpQ7SnJgJxCHmnKQCBFzqm5oABbPvHOs5qsoiqEbix3IT1hI4kERpqtAj/7tRQw31D98iA5TI9xJgoB9uDAFvWUNgZ9QrEijUVwym8/U/kT84g8bBJ5yfV+BVGi54H3UglBuKUVRWGsCQzq9mctlGk56fLUKsKYxLVbFYlA8rQwJczh5e78uIRscvk7aQckc/ASnufqI/JOY01wcYP8Idyq/aPPwzXFDZea2R8q4F4eDpmXfHy/GUaT8/GktZNPjo40MoS61Gq+C3vk3QnTGlsgie6QNV+dF1JD84uPKkFpqqLTslA3zATYvLGUQ56yx2PIn18kAe+XhHQriKIz+T92z1vbgO14N/C0fuBY8aeboJzoN7sNml1VJIniBBFuXl4dprlyC/few1Vjotr6BzK2i8TLQMts5iNkPJ8ga2rO+HvV6qAKhRLN/+9QkOvkQnVBfCXpBcNuttdGsR15EyTDDKyTotN/m+9Zh/pMxkwWjHCethw6iL/737/o8Nyz+D1KBF9D7yapBD1NN4etWJomQTsg93Q9+lUdnE0eUdEi6v22WGK8zYKnYLfwXWoRRrztT+yvwGLOug1qGHoHM1IehxfKiwIvPX9dF8GeWlPDZWf8fCDwvEn7ScjiBqr0gB+xLJTKXYqKcSQw5ALZlNkfXpQ3kMhxfBXIL1gIMvXpyJfDgTXJqgxsY5T1ELnfPDt4kgSfalUZyJPnpP"
`endif