// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VafQ/0Cqn9zksE2kecgTiQinNROC+e77w5PFjjQlDprwibbE+6jKF0ZeT7v7
6Fl+w/3RH3EwuV8MeS6lPUX5CEjuV3MMa2JBljb3Z743Ty/s1xvbrTFzsGPw
v/YfRuqhLSRrABEL63I0jhQABbqaHawsAzL0LnU1wBEVbBJILVPEEIDn3cUU
Ogy3UayWF9FyCk+8EPv2HnEU3oSkYT+X21MAM9wMp9ZRPBVCogbXRhI73d8s
P4HrAmRb6wJjP7ZtO0EAc4SY2EUVjYYrVqiREsa7F+ynWw5YLjpZrI+sJGOq
4vP1JyJBGAi6PMUhS5/lKU1gZIiYS5FkiQxO6hPkLQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bcJZvsAumVuTgJNlaVXhqZImHeC3oiELb5JVCcuw2w+o3CTwccyp03KybJpX
ivB+obfMDlwWDCk+GiBJjrKowWPXELoWZWuIkik1KspCwp07zwoGtEWlSmF5
+t4vYI4l2KiW7/6Nix3BJ0U1jDsDLcdLIR2KbASTse/lNf+lrcWcSuSjnw9F
0j7tOq9xhZ1VBiyPQMr3BSSOxmYVkEnulR0xFlBWano75QMLxqYTF94Lt5ho
7wgzSdcDlIIHhd4A36Gay+tA9i8RJ4dQy9d1NDmfMVPESRd72acC5ukqJM4d
zVjWQ6vaaj8BleoGd3oBo3+aqhZbv+FDB8C4S0mVjQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fq8pe+L3pHa+ZwJZu12r/8Fbx+7S+kAUeGZ+J5oJz6GED6LkjceFXbi/6Vn3
jTKVAmL36ACcrT+Akdl4szBTbBlfrfC+8oKO9+5zfAOk57XNLjQxcsBrucmP
dxz8oeBmkMwMqLjWt0r+UwbCuFDqnLd9A01Ga7qJxokqntHMiDaCQqWzrUYl
ACn/cpk6zfCIju0YPkUghN21PiQTPtYX1Wp3UewdF+WzM/JWUFunj7ZOMy2t
q69xML4cpKMEhp80ewyCpo3lZFpv6/ebG5cFTwIrA7ZqQ+Bx4gRfL4dOruVU
UjGF15Te14Y3tdmQzC2ejP4hjGCUiiv54Fx3G6fuWw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ap6K93z+rQGvfTv6pFRSPITxFlJp4sv/BzAjzui6GpME7tUyI6VBsuo+1tXA
ZhGTZGSTVlKo4FnCJxfLfAmlhydvLtOOz/2HXi8/XQSGxioI+11QtybV5Pxm
Is5MF53pAN8jUeS6us5tWVNzQJhhYaVrRsQfT4hUaVq6htpkVlIUIBMhuMER
R/JXvoGvTb8rqjfWm+j+Zuk/QyrYgpL8kRWngzh+rXLlWjaCyZsnaAs5+4dU
sfPhGWre/fxY8i3i326JmyVJcBSC9Z/YgRWWbhHZobWf5NIDz9HuRr5PhyRz
KEqhPaCDtFU6fPqT5Poy5953BFeXhsLoLNQeVeeGfA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
T1Jk4EDgg6uo36LimpEvWCgcZ6R2gbFxJt2F0QZrG7tD5VSTmfV24dA+Y6iY
rbplqPNxQqvfFBZc47Dl++ZIDdxh5VH/jNcupUVbHLuzVnXwo/lIGMDPya9f
emuIdVNkXZl/H0On/EKPlSmMEiavM3b6lUWBq1OTN+SNVNUXFLs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
d3tGARF4k6r7AkMhwQFIotE5wYTKojp5fmwauBmBtouwj7WYaeAyTrYs//ME
g8kXjbntuJyxM4OS1VCOddpReRH31nL3UA/0m+JVbpdX1QDUmQAalHWSTI2t
komlc8hWmZHdSHgYZqUbbjdsBCsXf4FYCclI5wkxaLywx1t3Uc5/cYjlQKPf
TzJpvs3m915eACn6gl0F2NheIORDOCeKtuJvZY8qDQk0A85QP2Z1Uox7X6g3
q+ze7CPdObH/4tuaJ88hwzvUTtB2eXK+5DMOvOBN/KmPGmPRWuy4dh3EkNIo
2RRC49w598WSCvvAmMbgmRqo42iBXVqz/+NsfNAmtjJPgoEGg+mwWkUgY8NX
Xf8lgfdUFZLI7MB9K9EdNiNIBzJs3BYotvShRNd89l4CVSqQFuc/Fors9Bgz
zW5fP6jIYoSxf7CApWPbSfoGoZ2nv7g2qNGzJEukzPCzrVBIZHYikGI+ZHiX
lmgAWox2RBdV1HPfpmgnS/dMh3pjK/yG


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qacW4iBanpxYPjIjBIPJqLF0mGZzAkN+mX7GgV3fIly27Y0X7Rv/W983dQms
dQMDu+eh1Z96lFyNES99OKHW/41i9YIJX2d3db4jKk/B479WEDqqfG6no2ZD
3p8iKNRBkq+t+/fRxsL+pZVD0jAnnx2556uAPYi1WHwKI8Fx4kc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Nl2JV8hOHJqyl99qPPh1U/gesdWG+1SxTCKaRiGlc8yCzMgqxi9tF3vALjwu
/qEDHgzKNUJVzs5sFEcwOPgQ96octrgbe+OqTizLlWKFEClUzZOdrdxQOhsS
yA0tNyGvtYn8n4YTd5N3UjzHirqPmNEJ/wK95i+noqrdOENOoIw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1456)
`pragma protect data_block
2SKcSmgb4V+DtPT4O2Xfb9I3u1/edvjO9cXLl0RSSDsuQSBPKCXNfUKlQMaC
EDVqDLkwIX8KkYpz/eOV/hTFTskH8Wmoa+l95YlNbJ6219C+arx4jFKWbKkD
zQCFlHdH9k1zveJ/0FHfP4pjmfpwNBiIbhkUmtIUpOx3V1KXwN53m2wNMa6X
dAYlWgAojAovjADSUw+AYDlbXLnWmzrjb3vq4a5vTqO0RgS4kExQhshbvlTT
iDrz57f4TMrnJNJNHaSG+GPAp4redhd+QNzKDxc45D4tcJN3jEaNRIlWUCFp
OslxmWw8AxirCpEKL11og5TC3SXSOLZ8WzUf5dsdWhx+lOQ6GMLey3iZ1IzE
oKnHZGlkRgpKLO/jd2uzV9BvzhjpE8ZtZ03ErVaHBryVaYthNa2S+2iSVFxn
BQcSthIualIMT8Js+CkePwLj+fOcvRIi9VykmXEGJWgTjlrT7SFqqD7KtICJ
LfQhfVYXFQuRLtKpP07XMIMZOT1rVsDadiBvl3EF8poSW1/+N+x7WKJ34OoU
GhKa6S0LiqwlydaDJipieaZd8cgkHWlPliTQ8dhdbgB6EGuNG8KIskv9qa8P
xClEiWFuwOpj+iNzmWSkkhcRIEKgW3T0DvT7TY53OzJRIz+ANH8sotTisoTP
OfikI8r9FRtg9W6hsYbcHKm5OAxG4PFMf9up5vfw/IRHiAjr2POFDq2IcFI4
7miJyBd5fr4G0GzP4GO2qm7qffA5viWiKmpEKPDOLx89dGJ1QGhmVzMsAiTc
d2lQvP7KtcPPITm11HxL4ZuyUv5aCtEsksSzMB7gajDgMtxA/G0R7rZwNK82
U+oQEQU2+AvUVKdg1dtqVuOZOdFhRhwCUna+Syo/v2T0YmqErQ/ICo7lzuP5
g49T7MBPhWP4bi/iLldIIa1ZaPqrpgKUKReSvPZr7uvUfSwDkuajDEdCuQ25
SVEwODBOz5teaJ5ltxnJrDaL1zu1Gc9+4r8nL6qCVdBXRKI+xPmz2XAIaAs4
7YFb40HfmfMrME8ozFp+quiX2NNSc0zpV9l+DFeImHP/NnfoOkcGVby72Ew8
xEfh0Z3FI1C8mQUR5zXwxSGgKJ0lJ3rS1AgfkKwfl6zubi+zC10p+Ihp8zYT
1pa2fKbFag1Ghd7r0ZD0VZaaa1K5Pcej5PWZGcgLbWxM0m4KLfNBZMaqUhJZ
qN/194q5w47zNplMXmxEP3SXVEIsns+9YQreNi3yvbneKryW17LuegZr+qj0
8I4C0scMQ/sKX3Tu1OgTUnc29HILOK5tJh2bJwHjDeg2+owaewMAPH7h+fyP
G/IMrfN6G25bkmwXM0pJf9ODF7Yv4g0Xx9aCXjMVojyvPUBAQ6dz18CVZtIZ
a1oFitCYnVrVzq6M9d3zYSTEdSbOi7bNCbj8otIP2keEZyCTNcWf2qKh+tdO
4m+/NjnOiDeBeFt/AUjQTWal4yE2s+cbAmFuWR1ltP+l9lV8+m+eFABy15Fd
ZaA9BVoP/tZNKsE9qpVEN+mZWohuZFBPNzUWosqwFOd6OMHFnb0JJ8kLyeLc
0D3FXwSEQ67hT9EUjsTqobIIOyV2K4Gl2UOB5jNtE5XyeDwX7kOKE1bAZ1JS
8A8gE8DrSzFIL84wcEZMVjmhX+usiTMXfcYtoETXZbR4eGnDJkiYgZWjGUl5
Qg1JhtwDCsKVTFVCQ/DMw3OIsvcsGWU9DKUrdsi0MRklFj0RjK2zqUURxd4t
ifQ+syEidCQMkElOIVNT7JrBgIvAo8L5CAW6PGQffC8NJD03xNfYqfDvYwbh
yvBq1fddfXxIYb00uXJB/UyyTDZr+NMBUCmQWVEaVp36uSoRb/QXVAZf3aYt
flIEdelmDAkIovI/55gZMJWra3KTgFZVFB+jTQf6Ocr8BeWz93ILnKKGLAUG
QH6NC2guOFXE0kTdVnF2qg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqcTbYtJICkeBpQuHxtKWJ8N6u/9QS/He02/678YfCFbhW2ZDLY9VPEIWetTfEKDVPOqFFxCdp8cjg8/1RPqiV2LjlqBOE/6kEPCDByDhvL1/MxBur9p7Xwij0y3i2qvXEwHWOAHj3g0KDL90bTksMipA3/jMF528XCuH5hHymwzVjsxHEWZXoyM1QcPW0yD4h85TgPurynx5P5k51yjPjizu9EXXkyV4pXdgQ9yayMa/5IgaDAQDUg4iWtVmODX0XIFnIvHfTmhYzj/527I5DXXaWppOdFmWsVsw87Fysez3r9L5EyAsb/dKwGkJ3AuOHc6YPcT0clmnKOCK0kp9EuOP2FId22JOUfdT9G3L6tvHoh8duXIoGa9GdO0Pdbb/6cjMXD+ataVnkLyPSdcmB2Zjky3UZKPWzzkjptdpZVsB8IsI2hdEpXo60aL0ZrYZ7FjoCnh8n/W7GvvbyRrcIDDNF7WehmkWhCZnvOMEs7iK6B2nDMp0mf0W+wuYzNhpjkCrWcs2eU8drdgA8nQZj0h1j1zWnDLn1xBM86xCLxFVovq8lrwCdGQ+u7jWabILQjp0Y2+WiqFhD9mZWWx393Uxs7upMhk4ZqQ+2YqgCFB5x2GbJ7xFWYJK8+wn6eaiqQWG3Wfxgj2mdc3e3df74o+sPfKoD3nzMudHvYYYc4gsT05oA9YyZ/IsrCNnAJ9rhGOtl9pWldGIn4fPTqO3JEKf3unoZLoLmqNfPQqYaBf8L+iFQhwM21MnKkOSoMIJggV7+wBlv8BrjoU2zGJebb8"
`endif