// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
flQhXCc3qf7eHMPssf4SH71a5ixNEdM/aud30D4YxSqrvGfziJHMzrEgmKbG
OR39cYNxKzEdx1qysL8Xc6wc+1fdbZIemBmvJFjyU0D8FFxdSE28qtx1ll/W
pqpAn+3Dmv97icFeJMA9/Ty4aamXHLb3IYAEc6a0GCRPiSH9vRuatTssIeUz
OqRUL8EZSQXksIYjXP4phNP//YsDg66uanRwTsnnmzJuQi+2yDWy4QYGyyBq
dqPo1U6nGZuU0m7gCTaEV+HD9kMJrm1D11ggk4Itgqpk4PdzAdeCxOQXofVr
wrY1P44KZhyn9yABLh2LOt7YkciKYK5pviQHPz9ZMg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
czD+1ZV2AMfB9hFmzQ276MzOAJ9iKYXN3Iv4WCCteldtJSvIlTfrvvbG1A89
fHFZMpCWESCKLlpFmDWn8fAxM0MxOcCNGviAnZKk8TbuRkD5wy2OWk2t/aQf
2Nrwfw8+gMlDvA0oKhVUnn1Ikh5jjHtRSPlyIjZBabScL4XSjShLXn/LvZBV
YewaxWOb1r5MunSjhoMlBMXOkeWSRjIUYRgk/BOHpCRuaXq6sxGnNfgIjPzF
WT2aD/SbTVY5Rgyc0Q12OBzcX7JJYsENlph5v2RLlKPUN74ptH17f64dpKlc
f/FtKmkhgajTO6fEjprWRhH99UpZqZGrfazqMFpGeg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Bxd+OBiGzAwxE/tPiIeFyjZhNaxQivjoi6LqiTeFeBuIZbCdrAPv4n865D6C
9iN1SbWTmk+MogbQ+GpD8TOfrRVNUrc06ZkUEEUaazj0mNUD56MR9rSuYyRV
+C2s1QaG3gk6mTeeLE6SsXn2ytoAlsbvygoni+k6PQwCWrX9aHCURVMJ6DBY
1AiYa4V9QU5IOykJqlIwQkFtcvXMnWV7KdKvg1DLR63+5FMFQEmmeQ4Pizfn
NmqreQhgSaeCSZa359iEb4SRj1IZdPWB9f4HredHjqeDnCP77OEnZb0vwjxm
S0aqXFCGHxfRnXKjT5Yly57St0RrOBHZ/WnblCHU7g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YZtnMDcNT3sdOPZDyBLZ6EFNQqKOyIKl24xyaY6FphmCMxadvzLCU91G0z06
dumeJgE0jIasrMHm07tZWW689r169bkzWGtt3CPsFbIbOptwLBUX7n7ZqZHj
EAfyGrs+5kcWw7tyKOoSbX3wOOWsb1594ksglWvnFIyqe8HmbrYuoGlOeZlV
KE6WqkdVVT0KUX9PmGOKlGh+Ww2MvIcBCXNuMbvhXyYGmlF9zPTElQ1ezzh3
W3mErqjs0qEfes9Drn9bR/t/SDYVuVmXAISqKrrQXsB4NJVEuYa6xI6Z4MD/
fY3QNvqlkzCv2GGCYioM3M/YnxP1b8nz0M2jl+2e9Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hMB9uuuTxx6nO1TU8w2YxRzLkroG2TZ0TJtHqBt/aoNQVl1IE8ENNbeGsH8A
542rpw8qT4aHEp7LVZOdqUM9Uh57UbJCRuzmNxmjIS/TrhaFXH86z+ezbMB/
nW/5DxdkFzfK7MBDvntQzkxdR3/k1scjIruCYksW8Rc4hfvDwkg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
p3W4No7jDqrQOHXvZ/UdzJev1x7FLbacWAPmb/Q2jhQSmd0EV1BsJF5dYd7D
Rg0114xWiq5FKYBNhsRye+DfICjvmIIYTpMZ5xBj6noCfHWB9UFYQcZKv1Fc
nIg5LvZ7ixE+AkbtSWNUA8rOi/EhmCDfH/Ln5lYL01EPpUHOg3/mYc+YQ8+D
51JvlfbW7Wn1ZA8jM4XOBYujlzd9XIYeaQHyusgNHOXu7hJom7zAjH2p5IWG
JWVDI2TFw/xRlvUSpV/su7NtDim2ZYF8Tktz1sAP+s5AlPyBr1Gl1wDlwiBF
KHlwUxhvBAliNUmHXkUA5gszJAbqSgFAKtAFPhJWd9GmLdSQgLmcNCji8Yhu
mJe94p+Ea87n4JjxE/aCqvfT2qNwlA+FRmw4nF5k5MNt3f9prEwLxRf5foJC
GoGnjVC/aI8Nz1qqP8ASU/ENdhd1Zkhyecm24jqX+8SCdQgGmmcPUCw6EEW8
xd0p48tM8r5AvjVrJ2NTJbwOoNH/lFcF


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
isMCcX+lWaOpURy7BNTKIq1KUQIlaMJBuPjBnE154JR769W8SWjzext5BC30
rHhs49qhc2z8QqqbfQ6vJ7A/XmWBx5vtZrwXpbqo7oOtTr///sUQzqWoiNeU
vTVp+loGbVv60v5Xt5fuOL64z5oZjklhKv4ql76RJ8COHV3OF9w=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aTJul0T0TT80fADxoUiqberqiHavhLYxtkNpiMfHiqI4qM7qTUE3/M6tIdEf
H+Uz6r45Vi3bHBGQHhnwyQDRmSGbQE6u4uzPRfMxNghRgthYMb+u7D6CepOS
1vR9I4/GFW+fR3Lxr9oTS2W3tjzEChpSlDLC6TMu/N83n4ANziM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4080)
`pragma protect data_block
lA1MW6QC9ZE7ukBmXIOtpzOhCE8ctHpirNRlCT98ahStjaq4mgBdmAtaCYKr
8SSiyrsWL+RLb/r2u0evurbvJWHyHhabmQEwU4YOrb1mvhmCPDXa5rBoD9rs
pTD2VPYrDxpE7Ixf7KjNFxj5Jjk7awj1WCwDlrZQAIbjNKjRio1wTGEAf6sC
iS91scKk+3bXXoBeWHBf3YD1hK7ty1FPVO4c66+WujjlmKSKYxhXS960dmzq
zRGXQpBFvpXGX0TcnL/25uxzqUbs+CY/nVLdrOOJYlvCPxrcEok8JsAc8O8l
4ZyqNikU9O77TwwNMbZbUwzI6Ji2PO1NHe3XsCwU+vspEGnmwqnjNa3ZtGPn
MTTRGa64R+NPg8yZXETCWhIcU3YCb6e2t38biy81Y7kAlAX4LMUfqxD9SVLZ
4Oh7A83Cbjc5z5jSSxL+oGiBtPBMlyoQQZm4k+M8sShsPCkj6cB6j29q8jrt
qeo4/bg3eNcU0d5rD2BXnaDtJTorIXu+PC0dJYpYsztx/TXVpWtf6+9gF5rJ
Q+Nm+x6jUmM4BNBs3X+U2AtzK3cuA+W8jnuju+fCXDkej4aAp9Y6t3Qxv1AP
NksQJ+EHb0Bqkc9A0BVTssc4mSk3wySF44kbHWhrRml0DKUNFqMgEA/QtG1L
h2wTE7SxjeAm3qja0uaiTIjjhHdB9MfRR6XI4PAeKA702kZmLoQuCgw41ps7
/mOuSkLuOJKhSnNK32lEX0uzfcSXr+oqOc8AQ/iHiW9jjL+1+VkSsvNtuQuo
1scCax0Ar4D/HyHYanCIgw6W5X6o6FBWec8dD0Idmgzt18/LZxFQUlqf5z/I
a+J4UhTIijd8gS1YnVRmypg+xyOlsX7TMVzjGEV5ujCSls5Z7PWPb5plaAcD
iZ5s/WgOF02HeXEpUns7HbrHlUQs0q93z4m2IT3doTpernAAgeptddPP5Yar
8QpPNJdi/y/Y6Y+PDgTFI3ZJ0WKlTrbTppNY32clCk8Q44qOF7kLSBAYZa+l
A3zwV1KRjbgPLm5fsyrDyoooEnJ3cODFTJlNzlvskzZBvKcUdMOeuYM9HyAG
cQsVbQ/mOsKMqV3uxWOLWno5OXzN3bSKbv8nWpabrLsj36gKcgedXQXwmedG
MivSPMLopB8urZzj9WYoZa9GNGZlXqZThaj8AHVCk4b50jWFzdlqIuv8LezW
+Iq1gwzy2g7AF6BS4mXf9un+0tGKldN3mqUVRSkJdtq3rTCJIa0BngMjv4QU
zuDdJRgAG5y0wqZjEgpdd25sXA0Gq0zsAcZ2NqiaKvv56fTUb44gov3Bb3x5
MdV/lG+oNeGWxMLaTCqkjTSiGDu6srkUpYkmAQAtek3YvtNH84FcDkvg2IED
WoHsYWu1zMjz9Qy+ZGFu8PHYLDcqNWdFP4gg5uEDd0bDEBYBmJ/K5Ve+8E+C
gHI5pSadv4Wshz3GOIiuMuv+eCh/gaQIFIguC9NVp3itTWAtsHkK6rJ4XQ+9
+772RR3vzylMvUG5i0RIL1O/A2M8bhQgFIQRiRupJi5U0wTLp0rD58qsf3SN
cXoXb4z2FZkYmNweWb1m6jGk8nDpNhiGAnl0tez+cgk7rjymxeYdLV/EaEhE
du0/dQYPDa+sSPohmrOE3gzLD5USVzpJG1ro//2ly/Su30elP7j40bIB2yOO
qDKSq+yz2nJFwchv/g22Vh2e9jMcAXT+UIKViu7t6M8fXms1eA5iu6knpJQg
t52JwQBlmF+Nf1RD2/gWOPmozfuHPC4JeRXUoMJUVnALgw18g+R8xxz/q7+w
VOJ2SwigQNI8zzB8LqyIUKfZkZE50YpoT13cn8FQNSALgcUv6gJicsupY3pp
npLWvbeVFJA6eDdyMw6Sy0b5krp2PmkYOzgReNbh6WF8GDbfQbdResCsf11a
xF0jQb/VggZtd2NbIa2doQmJ6Ix7Q5rocn9rai3NGFAHs45zbLSAYzMbFd6b
7GNwN+zWi1MWOLFIEslEsspszQnd9sSdKnimQa3iAul2trQ8MxZ85Y7KdubH
sYUtOHwdhQ5MqcNTJf1qs3k3KbGUFR4b68N33CaLVfSkWLEgULHqtoKrBQRf
NxIBvUmfIRZZyvoK3h44GDgxFJEXlkVVmsFz/m320ZVf4l4zpB0fDnYdX+jt
XpHMYAYcOwUqbeLvZxthiKPLrpA49f0VuPV2qUMx+oYtP/g/dzAUajiOSoY7
kpQ/M6HALmYS9m2QO3pKjcPvINlIobt5M2Hw8Q95p+GMCnhQK2/aCu+SyjEY
/bBQrGyyCAmY5eL8sWB9/HTa5bnczY6yNCJum+5uV4FYPJDsgzRYvDb54wP8
8PRFHRPNhrbCK5+YfG+1VxtYUXj4RYYfpkHySKmjLCH7oeWVaWlYqdRORiun
NOG8DWqCSTgBov3B0LCq0SDMrQ0soQ6bJAPKlHargcv9GE6UgLs9Z5z/2mqR
p5RqDrBaDg1/VvrN4mJI//KdyzoHr3xMLBy+FpGBJPwxEKIaTFHTpDxH84Kn
ZFtRXGB/7uaImcbMti0KcjKKbydPBmm/MwY68OGhP8XpeYFwau8oSIfUFkAj
nND2MFHlRdanEZsNc6CnVhI/Y2K25S68hErYOqGWM+BMBx++d3SdIC0QQcoB
R9QJNTqUF1navRmUYxlfxi8w8PnEsxqD8sW/gT0H5xFjQebFq/Xcn1A8K3ZK
h3QnS+O629M/sklLzC5PM/uBffj9uHbuxbk9snWN7rKyW11MhbOoEtoPurg9
gDTxT1oH6i9M5Dc5dcW3aVm6k3U5GLLFiJDvZdiUmO0p4WzIGTQk1/SPFo5v
q0Xp+cRHoAhQRHfpG0lgogR8YSffXAaioX8c9zyOezQyWDX4HXchhQGtJFeS
XNjfUtePkD9Cc1tRCXh2V7GA/3oqpZfK3k7rg2MxxnIu5jeM+NuA3z2pl9Ad
6KaksnvqTQm754wsYKFhIuRLDsoS92KeIQGJhSAhhhNoJLkb+GYDChUv3422
AaxyzS5PHrtxppbwn0v14WqyBJjXFU1I28d/nODcC30VN7dD0eNk2AUrtxpv
SM6mu7F4N2ZR7W+XUHRAg8XPhSwrEQX8SLsPJiEzcwgvlMk4ICUfaXfCklF6
cAwr2GI6ye/KANxs/mpHPNNkrGUXKrW8v/c7FdKJWIB+omYu+hpE800WVUff
T8wyYxMDFzyoyB+gi9LP0WS+zgIcDhH5sMqf6StT+Cx0945quAxFUbKyN0e8
fd7sxnvpJ9l7o5YaecLoxq9YOS/ZoR9exKwF2naOdU4crMCZEbHZIuFDhGMy
14PXbMKb0GSAKrKXGlIrM35uz5LZPM6mZLweZ7Tu+9mDcyMQyfBemp7FN/jk
VSaEbNjCwuDTSokbi2kLrqDK3PKCBmGH7gcYpgkheGb+4F9Giu+oaWPs8x8k
mf+SL3FFyLHUOArG1JeXaVAWpo48Ic68fhsHwgcwNkowztqXuTz/I84CKuG3
Dtnn2quOGM7fCmiySGp9rgLi71EYHGo9DsdQOH0F4uEBy++ZAJ4C1DI9h2cR
5yGcOZNjK+kQE1KBjFFRWq52Ptx7LlFmqu9fufT4Xc6EnsQAIbRd/QYjgj8x
fKtnZ6pjJP2oxt7CdPUk0DdDJU3xtxWgbQ1CR3uD5gjSNIE/gYVLFB0CqA+G
MFeODoSqvj8GZo12GIgXWnhAzFL9qUkhNpjcEh2DXG6XUdAOcq1dLs7wyrHo
EmiHM3Sj7jDxVxFRdWVoPNYQEJorMPWnjngjjDMLgk2EdroOhb3yNTbBiyqs
HNWM9ZP5FckgV3eqJ+USJ9DT/rfoOxnCY9pvD8K9B+Eyowoi1ZnKEbRcnS6N
jD+RoNNHL0GTWqOj2Y5z1d/kwsgjIwXbRIFv8pocWaNAQTfNRoSXZuiw9Bty
nHCaY+7Qt/YCW9hU8boM1CkMz97QLXZ7Y6xCjHcQMpY4GIdPd8v9dxVH6rGk
FcGkLYk5mjCUEtEMb5l9aih2SCXh+xFIkzng9U5aFsTFVQi8ESKdDu4F8Ke3
PpRkeV1BrfOHJITaMl8BSJCvbNODLW40k/v4xz4ix2pJE95YLjYgJemRIzAs
dMiz5ytJUSgVOgDvKZQfS7SnZWOBWqG9FWVjqOTBzUH9dO+rDbdWd6vFU6uE
mimSXtRdHrnrIRj1/yBe22W+JNy8SrsVnZRq3x2V21D/lSuJDFQiN/eT10gz
RC6Mwd/cOg+B9+fsfjAhSUlOjxU3qrOp3YQ5H2l8Ffmrz1SyNy573wjNYkJY
Hy4/FLMDaKa9Vz7XO4iMO5+sZfpHcxMif84JTA1BgjwJBEu79IUs+s97vYfx
QtNzBQeKU1QhQTAi4HjmgzMrftuivZuhk3XbBUJ4WkNs9zy2cG/U+sJp1XQZ
g6YQvsgdGngiPjDvRifAiHqcCoECY585uzDCdDGzn59179uwZTswUSP+KjgV
kqrPmhwiIwt4dJgNr97hGIlfDls2/NaGebqSmE38i8lBoUEEh1HESGrTFOu0
8FsIH86R3eX16DRu+CvyDBKA6Usm+yIlCtygX3/EWXjr8imsWNB0BoLjvesb
tvSYtsaWmU1jIhVEA1sEGCwFMAMp7lzScTLZeeZjHmqqDS0KytQ1bhASVAwb
qh58e1v8SdES0PPsRM8rk7b+AwW/702IEF6Y+YGd0+fOY4pNJdcUJiRNzcZe
TECpWwS0ZCYNyipQyAM9QmwMl2ZRI9JEyzVMopMNL9W6pRNWAZYXDK8nj7c+
K11z4LQeWda7Y4nmEqTC1/5xrouKoEhW4DcZH1awnMXoYjJxH9qEmioqI/J+
q6XdXCBkoN7FLUsJM8j8EgF3l1cSe2LLYfLxwc5qbVL/yRc/NqVotUrJALBn
tAtVZej5zaeUBWzXMKdm1qC8h7J/WCdLm0NOQhTElcSCI/x0zx0qI+ZqvC5J
LVYIlwTkaMBU6raZxqSFZ5kdlmfoE7Xs65fk4RH+lZpKHHgZlyqzOWpCOwor
V7c4plxmvXJTWeKDG/ZO5TkLGn7FbQhS5pp9mSHLLA+JcYoPaPp4wplvdnMX
lMABjZzlEb5QBautnVxmzpuLHQb57K1Zwx223i8/lTq96cJGXVYBt9/nJQgf
oBGhkR+IBMLwdXhfv5hsf9s2/FX2lV7rHsYBhGP6ofd/H7IiAeBOdVIAV7TQ
6w0fPM2xrfHGyIX9ytYHpEO4DCemySCOYhIg9lvVJ9oHywiU7XkKv5ZLPAdF
zOYWGrYNcVdiHPyrnSJ5FRh8WjqrP1BSQa0xNqsIoDio7YyuKIXWtxZwwLDw
fUqYuHyKlWrYE02WehDjm3EXVdBTxyTeO7PqhI46r5Un2e48P/ey1SEpisn7
gXYye3R9Shf6Q69uKBy5U245orAPV3eIi51T/p2xh2gLC0JjL0VWIEzIPjgm
tZdaRehjDIonPfM0Lmp36kgrw74X4y9ZLyh7mniW

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzfRM+F0lZfQOfW/M2Cp/WosuoaF6VXHMAbimbyQVV6HwerilpJ0IR88QxksjuXUTLb4ZDbbQc+xyUBfm94JZLW6764ZaKgXac9qT+1zehIdVR8mLQXr4B1/oBkZBeBNS8gMBwf+xC2BxgJGP5tvW2SvKEpazPXIkRZlzDcTkbsGsALvHNUzit3njOaRu9VS0Px8jg2R40aCXsDM5B3aVIWM20ZT7xm4J8/xJoiYNkjQCxQmfln2K/ljEYp4oSfmMR2SN2mgOWaxdHdsMf5npqAk1R0O7kjp+TLUkCUvaglMHqd1tvjbPDmR33kbBm1akEFCIgua/EOj+5cmyUatXDvTnqOruRyOJzuN1n/zSeudORDxlYwzIawJ1oqraxM7myyf1YtmpZTpy3ZOjv9G5kj2bV8rF9RLAlFXPs+r6o2cq7zAZV4O8c5fKnDj4hVM8CGr21uedbC+gDRbz9sQTP5u2kAoTHxnjPPnb+QsqBzEA1hqQ2p/NTzc5Q8izt5zh/q1Sb7eOP4R9Brm7DyYJ5wu09rJrSB1FXLRWKRf+636WFe2WWdPI3f+GYn3rHL3xjY/5zbtxO09rCloA8NaFb4fBaWDjB0CdslxEm5J5GPzrQ0WbYB5BXyEh0ye1U+inwRN1H8auaEsS5/F5R1fTiSDjbquoIuqmtrZkWjpGaugpYFV/zyDOYwCZQu7clljJ8rEwu22zD2lYw65oDrDiYWsZ8rf+QBcDxWBneTPyxCWnsHzkvDAZQQywAubaG1dSxlSFgJFuV28HZLMhZUotrS5"
`endif