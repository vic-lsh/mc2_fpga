// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
A97qkof1WkYg5UDnTJ8oLN+Ecu8DjFIIYku5y05/cHuJmnjwAzw/IGKZTaFu
tIq5VcrCpigzDsjLfErvwaWRQU3cX5EAcTAR0WSXUf3ZCOCD6DP1/ZRs1S8J
/SGkWpK+BlK7rKz9eCzGu39ulb+IoUhRIX061fR591fySiQcpd/nxFJ+KplI
HaM0AcgJAOZgV2rtaN7cL+KvpnqluKUnjyAMzN5NNt69fJJaAHCYXZeMUiIe
EGb7RDhdHp/sLFrxNntKQZJGClh6NmPBkpIwMfFDlbPAh5lN4M/rUibGrLIn
+kRUO75RpuuzBwJLt8MFqctq1PrAMi6WRczjUaencw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FVuQ/xnx5Im7yJQIGSLcjzoG9jPgnLG89D5Y3+izpKEGRMlIJpfCHls96zRg
SIiGSQNYpIvDptGujbe3P4lgYWOZkohGf499IUGvHCAasMQPT5Tic89tlj+P
UtbdkoZE9JbqDIgxojuqjgF2qKI3cBgiePzDmUjk8Kej9ubKYXWURfPUe42t
GEe7RMiG+fnKYuLRfl5oT9e2QZ4arv2YowvFiZM5eZf05H8PKv59myhrNh7x
B8qSWI7kkjmNfe1S5U5YgDEyn1nZAYkHrcNAh4G0pEO1rXVli1LH2p54HUUW
He/t8DWFuASr7jy0tOBXIBFYE4EZALC11pZBJh52pA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AlsYA+8R+IjFG3onp8ugsBW0MkgaYW19OmRQxxpg/85FED8CdPBsiKxTlsee
5DPrZXYrN95wIWI6lBmnFH6oHydqnASOdDrSM7dkrdQLPdLKk2sWDwaJ0edC
vwJT2cpFx95GdO9YQI2dByMKfozFlLHYix+3pKY5XJDX/WrdpNSaSz2e4gza
QKJ4bVwCOBTqeQu5JNdcne8BgTw20N6j7tKOMohMr7QZInQ6oGQn3zQcBYWi
MHnLaJ00+e0750HWgOpqI4x2n2LZsouYC9fkzw4CrVY/3ud4DfugAKazk3XH
jaUruSd7yYuC2FoTICDr3gfl1icmEBIuPHEGd8i/TA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qgHaficFztecPZdgomVPFwn1/p/XTX/gfi0SvmvnC1aOFNFN7CeqElt3Xo+H
JFZ/xFa39kaidN+qEWPRUVAzGYbVVv/pvXeTKyaG6YhDpNP4mikjNPlquAZB
FYmpIK/bk8u7ctnOZQRkjL9Ag0wNNLcJvOE9gOazlIEj9S/xd6pQQrtCE5gl
GhjlZneBM4KhNe54gnXD0DSr3LoyXOalG2xnU/NEomny6uMLoTqo6RHIR0Wa
mLdiUoo+zSeD96EybzHbfaTbHDUxGHfz7aUrvoXSDcGGgTvh/18EoKUXQiut
0XOFebSodViZ0N15MflXQ3ajMv46KpqPYAPFVqslBg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YjX86IK1tUGX39WjcPac8w0amtD6ajk/F1Gp11LkWitnkij+LobLMzZ3jnY+
WoRkaO52ornRZQB64w/EH/8zGMiGdSKnIlq++alt3GOnCy09GzZ/pTqsvTOl
ZSMUkLSVtxW3CWKkKFMt99LPPz2StKF7+yF0jaeu5dQnDY/Xc4U=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
aFCdeQO1f2VR3uS9TzoMa5muGsdHGhLMTVIC/PoqP8adJ/yACyIeesZr3APe
YXvx8haqfEfmL/QEOcXtek+96y8ud3RxFuiW9i4wYRcSAKcnINh9v+h/Btyz
LAnZx/eth5KSIZTgjD4FqtyoCtwPQddTeudfVbP/1pbHdEhIYfLwaL4w81Q7
qsF36v1X5nmiAgBxmQ4X2Y1QKyLhSU27XiXhbRBD3k1bM2O4pBZuK/7T39Mv
LOVMk5GOipXyR0AEnTvmZAeMpthqv/IfU/QcDGn43jLOegZQ4n4pT3BRgpZl
SGrYRjhjv9b7XGk53mgAYITl5X4rzWrF1CUAKVzPZc81yzrp377Z/8TIiMu0
BcqVb2W0mTwgzbM9vQQ5szgL6bwfHVuFZjpm3RWRVKkNFePOxRZn3uLsQQF8
BDhfUhPWceWnLmczNRbWqo1rpR8JDc15L7VvqmznrTRGaMsGDps2SeuE63n1
c18tA8uCzSf7ukI+487wMkSR88pv7oca


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eqRNpXt8QVCySYRiOmmtDMZg/7kgyeBJ29MwUgWXVksuEambkixX7nuodo3R
MGrjVrSlPd8c+EK27bu8mPwDXUkMv5z+n6gHoNC/7GQs+c35I0wMBGj5Xvto
EZe73LZxECCHypTYotrRJyXzSNh13LLH0/2eA7rys+8eUJ8amVs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MGMfVHolNp8aKPv1oTT8iPV2VKWkrWEXiehc9FwHGg4b/xr0c0ttnwu5XhsP
Fx1dnC8SAikkHO7ijUJKF2fpCKWC4sRgM15lXgYnVhBOuemNM+n8kB/TimaH
TnzxnNfD0t7ssn3oLhniGvpEuz1ktIOUTUkupVw6rlDAbWEEgZs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 95888)
`pragma protect data_block
Ba+5i3PKnf4PZNQuBFOtjOK0kvXRIwsRr3lKGfWtJgKxTiucI74wm3GlMXJO
nI7TyrUrQHCKpdxV1IJ5g7lZpu6yQI/dXIFSe/tqXPZ0/swKvgriN+SXnFvX
1h659IBOiZDuE+bX/baBpnDG0OtRweS3ZsThzqMVO/hXwtr55I/xcIPF1ELw
bBEJiGnjb1HZF387cChLgKG8zl9ReaLeVzejGejk/wWtrROtIE7hbe679REP
9tfx7BQRgQN18EtDrrF8mt5UGz4+jenUO1yRwQCGupR8N2EoNNc+yyD3wmTv
QZ+jbgz1m6SKOuC75Rmi/iIWnZsKZzAKDiF0QxLMQxBmGxGBZQQi+FxZO3C7
TINvDaUOxABiY4gZXwl+FdJ2AnKcBo4f0vg8hFLPeROBLWiUL6oEUNVxc5Vx
0P4+eiyC830jvbCJIVlxSxjmiaagOa8L0tUQU/z5ijlkU0qISPCvquJ9qyId
h1JBnHUSEnhVA70XP0r8iCqnIEuVWampP4KL77htglptxteA8eMvR0rzY2pW
onSEPnZd1z2W/LR87GTGFlfcqq4VFAAYB//n2VA7jirsN1j5ZT8eqbzpsXNB
Rxx95V+K4P2e6rRUkriY5nMaHfWeZRtZPwuhwG5pPcQrhUEj8PHnPZM4eRG0
q20muLdetkJJ2TZCn1xKlOYdDiVSsMFc77bI7pEFXtlUxH8gSIBd+86M9rVV
LW4mTrBxpo2o76UPDrMK3D8D5HW/tlGNmHdU/0mRfiPBtGcwBik10r7U0jEP
jp+lxrSQI7XuDg4mosFGd9IU7VKpqm591d2peP9G+iRVZ8J+xf2ZrBgkeS4G
8cnRi7bLkevAYEwvV1NIu4L2226HzI6qC/9HhI3szH4CP2lxeZndwfaoEpFl
eYNEac5dG59z/ceTof0iR7MK8eglsYyiADzM8GlxGD3hIveL/pcB3mQEN4K9
mFD3Nqb0FmpFb/b8yovqOvxELAgfmZ0vOjP4z7fK8qFz2ibhcnukvUczQCNv
lLPXQjUXkcInCVvHef0lxRI0df+mW09FkcNVFUue8I2ftB/HpgD6PVNN0PBO
erZtZJdTGh2/h1DCV242Q5IxYFsBm4/SGD+NTd3glnLjfi7Al5WPMIvqgGMY
EXdPBgUF2Jn9LfIanBNJJYSAtqje6G+QTY+arFj3OCBuGhqKQViKD7WmEz2z
IS89mnKtRD+nj24yRc0Ib8EtAyKsghQoRcvy1aarZPdWOjSrarVJSiQmKrZz
TEy9WZcAPNCPvi8Zq8BLdijb6+ZmDtZyL8m4l14EfxyBRGjxxCrNHh4bTNqg
tTf6XtQ4UuYtkqWzsVDFU4HenTmGQxWkLQwS2Z+C1o6YaT5zLy9ukBdZhTKi
D7v4E3r78U9uU7eZG5vx0mn688PfM2Ak7bgr/jiZJcj8gX4XR147GoqsNwrp
qTaDbv1qkFZS7vJT+z4CzaSGT0OLmTVvcdd9w+u2Zf4weT+z145gBX22Cc8M
GPVnysVK6GzgD/jL1hhBre9i5hDXB2DYWx3kJ0rA9BCQIzibfiDMpqIIqloN
/GBv5D9Mud3GFvpZ/U+PxLakqzde45xIJdhO82KyyV6NnwHSevp0wkXXx4hd
OE0XIkZq8eGCE/UYvN722Gz3CoQz0OOfns35KsoIC3yrkXpXXZbTGpgP0eWE
fmNOdnmWgcPqRd9aSm1xwezI4q9qgqf4jVf9vDseMAiR1ZfBN9xE8CRermwG
wpuk6l/ylPUltZ59Z1bH4zIUdKZLpEY/bDso1dZVzqgY8348S45uguO4OLny
SOomWH0chM4gkpjId8j2YjLr8huFLxXEDBqyD4zMZdcYcGzCjIGegynxKd7a
6WkRRJEm0f0QETFmB/e3G8LKvJ5ANTdWCi1hsW/ugLY//iQqrOAHIK6+pCq0
c/lI64wfMWX3pIWCqBzNpqNv6m8Z31pMCYV0YtbSP7bGGvJlbGjCBGQPUJWC
ZpfE17+BHP7IvE5iP8SEsOPV01K8sKLZNVN/sYejWlyLl7HfcmS8lhTmX49y
ay4o2d6TNJsMZGmZll85Tp2jmytyNTyZENwen/5lvcaWoia8Qm6iuUHLThbc
cTv70a0EcVh0l6zUOU67bJRs1oBhtWcmzVGlUgtogwBp9KQUPE6ervCP8YP7
DS72VxwoDkQKF6HZQsk9K6XqcohEekUk9SmAvLWEuXmptWDUmn3unQBxDf0Z
3dLhLyNPM68tGe78T4Kd/5FAPPdUbgjIsusjpBU+6dXS9XaDioMsF/YvOzFS
h8UbFb2mhMauQqDovt5TCtz2zGG/dTYAgqQB3bnf8ZFwVzmXs8FlumwqHFHJ
7nL/2wt6qZd3skE6T3w94bExQxraJ0cPBnvnfz7W5NOC6CVgDu8OeqO9ydEa
9zpM1vbArSOf2lCMFhzE7UnuUTaENI48PVR0Lh74PoHPqlizymQZKSbqnTcu
3oRat2B49OyVL3yYc0/E7qRj5OkeU1pnhUaLFl6zwj80yRee4QYEFFlng3qA
Hw4ngsaASW7uKXxjDZHj2lN/fQqDwemadv6/P2le0fryZLPI6npegmQowI5e
qBg7njsPTn5FvTuPuTgti+SBwe21dTW5EweC4mmPMWlgNlkFBIit1SLyPfnm
nvlsGJnniRkPXshQTJRZqgc1jpVWj7uSvL/Mu1tf4uKL8cRhm+Pec22Ll3no
BXUOqujrV3urrq9acPOH8lwgAJ5m8sVxQUHKZiJLqStGR/bZj0HoHEw12PgH
K9ugQEC3pIod8IOK/PdBzNqUPHW79wWnJDQAraCwn67+Nyy0LcJQkN4LlWWz
tDrlbjR4YcB3+l+j/vFzia0PePnoy+ZRsrHDbkQXn174qfSr3benH9zL5eW3
UzL32TF2uNZfVm0RkTQSuSOXfDswOQ8dHDd+R9C2KBsWi2h/XYAgwL4Q8rdb
dL+4peKHAX6R49ztoiKSrJS+VgUMDBiKs4WO3qd6Angcl4Me08fbvX+xSZfK
024N+X6LLjcRqz2TbODdSCzqHW+2EtQWsDm0x8Bpccf4RSN0aAEViNigE9kK
c8fogIILWy91UG+9d51pPt9PEIa8v4lGKMfCkAmpRYrzx3t5cWSc4D3YbwrI
uHgUx9R/AapDW5m5qdqRxDFm8KD/+H56w4N9LVkBl5f181f5DhR6ax8z+sNx
fQovwBJwdox8XiNpeKRwTs0zTQgRwwEx7qH34sUqf8ck7wl2vY91rPBlwFhQ
l71i7L2/KPDRNTP7iYbkBphOkDMaf7AtarTAR26wMy+3wDPO4I805Mz+h54q
d1YfbFd8DKT6YeYeYRz+dQtuEL6XQjx2V3vJG0qJcE68xs/wMzRW9sEJ0MW6
3MeMugRGuIFOfYIeye66wNP1pBAKm5RsaJEUaABexAXKuE+O3sUNK3VFtLK1
kAvUHAYYPj3OJ+iUm03UeWQse3bH046+Md2vgp2W+hAshFJqK42wfWjH7yln
AsqoMR2d/iYmcd5aVvvzGawokkPUXwiEFzUfktF31/eeJeyAY4A8jxa2Y4/m
ew1j/YaeWhp5CG0DYqZrk9zyDgL7sdPINGBhkwvVA+mw8z5Y88yGE1rs/x5Z
XPx14IfTjlZc6mIAnHueTji+6oqAE6IZ+x268pMfJUp77ldonXrbAiQEEtXm
wWn1HkVvUeV9l64h2or8hLQqo9p8dWxVbfwpuJZ5ISECG2vVwYttnphXcbW3
7hX+2ISwiBbLbjhIwe5uDd4dfXKjqS+oHTzPXXVygdJ3++lEyFjyTKtGl4FT
1jvy7JTbl++kUImManiHSp50YqnJVRKkOCW3b2oa9C2TnxRiUXhyrdcbjL8S
8SQvQfYZ13g3ucxJrd/z4LxPaJOmwe1XoU4NHT0cZ9IbapPpalQohaeaM49r
iDwjfWvqHpD0KomV1W6yZSLkt3p9Yf7EcO3TrunyVxtIw75oIcADI2q+7G+m
dNg9q/mg9yPgeti2xMeiph1I3HylQZVXFcnMm9kqIlfPElX1NO4YDoG9lO4E
0IEP30qk0KCb4btBxnCrV3Ma6CJNtg2utUJczQFaQyLwgQJbfrlh4NauzFjD
4VZNEeU7+uUUzo4sPz4bOUIRqRy7kDBuIpoLV4QWFlbxOd62QS18pbiMepRu
2CMxiUkZ1JvD2i2XNfI5J0hZ5gxR7hLgFPtBM8KGzeBFpqWTAFz93VI9TCfp
/z8bZwWfoQyMy8pQGT1b9EXuQFIGi1bzzaMspmpeHpDttzE0xJZHQkxaqPq6
SAsOHUzkb4Czc/SlPiRpV3FWaunH3nc/C+MRYuBfJ9XJb8n8eeCoM6WVW1fd
FzrRe61OFLUA3uBeQBP5NNjXDP3dSmk8uMc7uHgqRJvhJhDpL7OfBKGVbCqj
UIp9N8n4NmKICXur9Vod0FnQSDSpp+ZWlM4+Hgchl9LShREyQ+EumsNcoePF
MvKGAB8VVzeEWXLOj4G/LnWUQn4jgGn0ZIm0EOCzm+6oi67w5rPCV6x7ZmEP
CmEcENcovMOa6Ln7i6ilPYyrHReDtuTV0f0KnzzDEau2D8QA33jK/U1l3chv
w2yk98AqP65frccl4WSPytuAeEVy4ApknO/M5E+dlRHOep315t12ohn/wbkS
W0Vk6JrsXqVYOvQ4ltmzGBzwur2/yKhWkX9owdSNY85tJdlJelOcJw4uZ5rI
P93JQW6t+VxbIqJDTzJya9gjutz2G27T/NzQ+KQJA9Yze2ydd32bSAJOqNYF
uO/I2IokF4h5goGf5IXhFDNy+VhRPo4STmY8v5ZdUNxpQYiEvcSrtnWohr2x
DXJovVD1heA23WDr/KUCA53zzpeyCrnfIv4NN7ZntIntpcr0Wc7UsjT1BPZy
BA00WebJT+/zaMCiMnLHeh8SsBlne3nvnVXYBYnRpzm7J8riXUNMWp+3plB4
PD1NLbv6HDbv6unA0NDuDIbOBog04qmJbvKYiBG3QsJsLnDZnnWx9uMWy6vS
791eF+ebutvqlfoh7wTyDbkThbhQiTHhLTwHuJ1Izq2nlw4jIvc4Q9IgHgv7
4JnB/Lhh/sy9Z+KHApPZeP9lE7NbMfjq6ItMvZxyyKUfzcEShST+jbCIiCR9
zoR9aIaVLuBuq6vai/XKP4UJkzE6Rouj9N3XGZp8ZC/zpjNXiTSCxTBpCzBp
8FUwtUogKifSPthS2+ae0j+Xi5H6brGsiZw6CzIBTZ7zIkUOyArFydFKGial
V6wboVIFX3xCkI840nT4lC+WgKgIBrmew+E3pJwpgqmstMD6X05g2VoCezaR
7gnej/S4wy+5/TGvvlYUAoAXkbeP8ndFAcrNzxJ5mYlUwyqbrQtjXW90MylV
deznvX3pwmPB0g4AVZG0ZKQ/Zm214+eqpf4Tq+4WHhKqtIC0KU50wclMmuuH
T9GTVNtmc8gQPzVCrk7XkbVyoBGRZlO92KEhIRqJNgwY8iH4P4RpbKwZ3FeC
LmIWOuARg6MaYdFMAcQABy5x55xSYM76WynIqvF8tDz53eLRS2QJq03FSRmP
/k7D0nOryNzd7Pu5B5v393PXwPMlQvqge20jCfnRgmm/SeOGPV1qihDe1/VV
QUrWPbKy//9HSEEnL+GpI85fowNuoQf1g3MDcRrZZ0F7Jh5Fnero1q4Z6yWB
QfBgOMIyC0E9EQzjttW/hvr/+YBuv+6qLbC5jTi+ggDgzHMlAOXrpcbIDsGR
wyyQ8LxxQrrljMbAauWoX+BNyViLxvHZee9nyOwaZmMHQnFlWmHuWjRbcvJX
TuQSTOGrHTXTd/XOf5IsSpwK9J1IMqcNEtOHnqCYyHm76vqTk4KeKFcv7hAW
y8gt+6a7Qjli9srOYHQEWnSYiZlgcnQ66F/hpytNOV8nL8MRQ9DAl4A4rFkO
3rewGo5crAuMKVltnyiuKykGtbvpv7605G9PoI4MWPUCiyg7dPZk4qukW14m
KXsefvlUByH6hcf2uxFbu1CMvUzpxLloNY7KTnNigaSTzykiac7s1l7TABMl
iVKUOHaFVG7lK7mi62ga6lCEXNN/YYuYH8SGd7hIJdRgb9lNW4vtfoC2SDT7
DmJGcq1Ok56Dl1/cyvpo9bFgd+L3bsgDRenmSczxFxDudiKnBxJ97nJBJC9u
KsTSzbhOlmECd7Vmufu5sGseTPaJ1VwFH0u8yofB+LMmdsHQHgfsz+IIY0go
2s2kGFuNmHj525KvZOfgjdA9gflmuahZ3nV7lIPajN7Mj/NL0L5D1obSIWA+
XmImKHCWE/+IIJm3hb4ePq1BiDVGQVhbrxxnFYHhtKXZgZrKc/o+YfXq2ylw
m5KVr9vgiH4Zc5vFT/ujhrJTAL5ARGhT0Q/UUkcLyuTumNHAxUVQztVoq5/t
h+/EKznJZ1QaeGHP/XGJQKsUBlvAV5dPylyx7gVv4khW0m8SILMLlG1UDhkk
gkcYv7FvUAyyma/yV4Mdm+fn45m8267So5QsDIIfyl+rDtUd0yFv1/jmmJOq
r1IPAI7thp2eKzOpq/Y5YZnH6Q0SdhCsCejgDt9B0ogKUUuQO24hWglNQgse
Jxv9PgxvEEZ23A8iygcvnrA8ySLb5fJv/+dgwN4mp25DFHcDiD49ncrL6QHJ
jismYIYVwf0DNSRASgsYN2anjYCqJBkjn0aFxTEpY08Z8vceXKqzJrwKerQ2
mIMcxnkI83woHERLHCl7xKwxUiOOn/26cLm7QHrdj3dfhBz6bd94RafNRTAq
rQkI4cGTZgwumUPotbQEXCacWcU2PvGfHLEWSBmjaSyxbtmWXeJ6csvhtQ2U
iCb4NNP6wPbG6EvImI5nVYtG10nqM7c3pW5PZpbWkEGPN54AToO/A/hjvBW0
nUJrT6iZomy+6AeQ/eT6YsXiQGHgR5GYT6GPznjdr0unr+7GVesY8NHzTTQk
P6HqXHRSTMb91wA1/JYhrR57argLao0iYXmlkIXV2MmcbxSj0AuFuMC8xBTX
mdx6ShpEyYg9QBHgQ8/TcxSSU3E+oG0V/2ym049K4bUZ44DAUt+Xdpx5bifS
x2ifByh9CoTOwMulU5WMdhbJKptlM3Nubc/E4K0pFc6l7rWJMJnyJk/K1VBl
42T+KkXt1g+Uxmihrb0YZlvR3LQ/DUNUQk1SCtajvo/stoU8K0JBDrgnnCwg
GsJ1cYlLMUUFe++uJ7v7KIcoly6q+e05e6BgYKos1IpsNIvhYSYXt2JpfcQF
FoggkrMbpfQqqovZ61W7VHLz8ULRE/DvESa+sGFQZvMLlWh5sy6P36GYVbyq
E9RNfoGawQ8+M3Py8W4Np6e6dDykupowQKv2YfgGCKSNZsd9p/JjmwkHMbzh
C41Igr3Ef8/6lNMxh8jhRTcvnK6z2BF3IX7QB+REXRt34pin7PcqZchXDvaA
KJ28NaqYLr00k6ZzqZLGTrFpT1ssSQWTSluwFm7hggl7ICVR+akLYLx/wS+U
69MPi8mSln1jJYLcZUoP9ByacIrHp46H2QlKbtFyCz7Bzk2ohKWWef/b5Gry
Il6G0VX9/j5sehiPhStrQZj89q0+dMHoyRudy+fYUK2IKCOHubPrxqjdTSag
9vEa6g6gjIy15qPf9OTw2guLZZrwmHLWiaLkZ5dkiK4Zq1fCmcIENITqRs8I
Ya88Wnxmjm1SEoKZPgboYXgtZzSn0KVuXWGuX+1dinaUjqDaObDZTFc9P9M2
YPTgpyROVGm9DlR5W9btWW6KS88ebwC6EV0cWT4jRPs6Dh8UvHtOKkztsyJw
8BQMBV4RGwLf25FReOxXtndoX1PzzuE4bvJPnOFWzWlmBlA4lDCY8immBsPP
w1jwsIBp4dYG45yYpM+etCrEbxf7eKYw8KsM1oHImgRGSdMa4Jamy9Tjk5I0
3p8Omac1SzSqSUUrBcdxntU0fRCws6N2DytYuLIjfC3faCG6t4V5w1yXAo+9
rGJPy4PB40pr2xsSLnbg4gRtk33k+FuDCtS+Vw9plShx4hbhKBRHP2Y2JGhV
FgPATuIaC2Iuq09aVTh4l2Kt1s+1GMckRMmseDr/8QSxxgt95fIJYII4Ft6f
uxG2h9bN29mxlyEF1B4PNvVZCilvKUIhnVaTlqneY4ej/9p3R8Ucisk9DrxB
o31p/E31LovZWppqo+pbXiPNOG0AF12sSmIWj/kF47DmMmrvgYwEbk9Y3P+0
hVj6/zpcOGSZFZ9TeTwctjosIjTE6Cd/dVZgygcIiTIRf/UTHOrzod31EIXr
uzBk0EhEZiFT6T7FyHmAY9zHWDVmK/u1RqJv6/VLaIcvv29CSmaETr6VF9mM
qZ6q3AT6yddJy+xpGR4KVaItdCsqwm8Z5vYP9mxLDrwNGHj1OjjXPbE88xxu
DuyR7HdClM4sdxgAmw6EOEbUKF1Lz38zadowsUl+YF+xZFDJjrad9iH+FYSa
q1XJAFgAY46wJ+aAVuwDl/4ZJNOpNCRyRNEkRb0rwkR2FRwoDi3/XInCLc5G
82G2eRT9oJaz9SicFqfnLvVVCnbx4rG3bEFk5v2M7+HW+VKlqmJYmDaM0/Ez
bU51HBxqxWDhAS2x68didtTU1uGyl5FKB+Ot8qGNbCWFAyp7Lw68h7eeUfn0
TguZfoVSpjVZ6z2SogROnS2+jjuxf97VHdKRa3jTVvNkSWNrN8e4LnVVdgU9
qS7eYbFf1a4W9b1vYao99VRC/BLaLiqbI7nBnWBoiW7iZjP4Peg6CKxulSqw
+v2y3sE3cQ9aHZCjesx224F2q9VXho6KVEWZmwyKdLML6YVEiF/B0R5elHRE
uEMs96mfRNIBtu3GWgAsp7S/gCO7GwPm0l2WShjp5Y0XjbaILFUwBh6vj36b
h8UAEwEaqIsYX6NIP2gqpTlGaSqIdh885aWfUWdSqa/wOi8f0voXjDIhrKO2
hQkXXwFZDdJz+ctvdVOkE0ljcarrFcQG1Fl7R/WHbycaPsis4ZkhnDGT3oYK
8yRTfk4x7mY5HfhLA0/9Q2QGyOD3XB0M0Nmm+N9n/aAl9v436xgkaTdWtesa
Ti+gXQAiuxg4wbcSvSTNVL/Y+kETgfljaKS+rxxNKdPNU46C93a5bV2VzIi6
6SCPqCZOrIqz9HxV+KIXVd2E/XB9D9T4sb6hAgQhlFTBvISd6Fhen0FngjtB
ejdmaQZNiOhkMlayrtTYmCl9eHIj6lyMbmjqrGx/h9LLjpbO25+1bBZb/A3H
/XLyghHEv2T4B02k3ih8bb++zkPblSDvxYgA4niNpTGn2qL8rMgyDVrDpB97
xmmgvB3nuVCsD6/D8r9k7LzxcIKkLG8kbiohJHzlPRndxcLeMStCZ7ZiehpK
/VxhfaDbZRLd8yr2auaIbHrn1s4P4pZ1EH1LKWaBA1pWKzZz7W8tC5wpEXhH
NUB4odI9r5MpkwIeTEdpPcAPJOJGcsNLCNDGb1j6ZMm8l3WcXyrSferRA2eP
dk+fJ8dHaLeoe0r0SOGKpisQx5QzkIJj7rsObG+NU6tQ0s7G/jBujrRv0tRG
N6uKpdVGUMwowqHsNf6RFNbAVuY5DO8JDhX9xLl2xK6CU86WousXBZjxb+9N
CAo5422pVUsx0BjdiVg5ic4IQS3QRrDwxfcOzZNiP3IJVSaiydkz1VVhZPe7
x4Sxd/FPY/OTa2VbBf7a9hP520dSuYcdjJWdlKmp7wbEjK7EYuwtCCillwBi
ycoABmdJswZMTAFqXvOYXIwwwoAwa2CqtO26Mk/hEXy4SWekC8m/LT4x3yQx
kbfCukG9qEJeytu31F+UJ7P5tH2Rx9U/24loDr/0etyFoc1pW1vPdP+4Ev9e
koeAQqB9nOcUmd5EJJ0sSy9ea0oJnONTG2CenYtuBgKiWMUjkwuEVR3igag9
Bc/H633MI8K2sTSEui/8nem6YqnCHecyMW6KbJm7/4RQMrsr+XwPA+hjFe8q
i27EiU07HgofZZyVZ3B5XmtcNIt4yHe58cCFoVkDjuAzExyvG57Xdaw6RAVp
8tDkaQ0YGQ4DmkZlDgt6ECtNltGeriofEX+3krzdWfwJrjx0fODnyltW863p
0aDtOzWN72WlVK2KX3F8l9SCx8Bq9zlYzBCvM7XQOlMOEn9sM+IJE2NApUgI
moN/XMsIufcfGl/QAxQOS3eaGZmUZhnwqiHA8o+OCU8rYbHGSTGjiDr5WuHE
ux83XVPOhWLNp39qxl/bIEfMK3YzeX+wTkgC6YMcP8ldcBFopklXRSebjkLK
Xd5NPtbAvHg+N2hzKSxUSyCR/4lffN1S0uCFv33xJpUNNgBQrGiH3HsyqDdS
UXf/CG1ko1+hzcmCdULhkKKHVE02eBqwUdN92z8gdBJnPwOLBU3Vh7BWINKx
0SE/xDjWiyAsYa8yHW8I3eZAc9J9uL9GYIlqIXgq6hCv4HHVKArTXaJIihbQ
Zf4bzgD9u1lImp8z9/9S7Mdmv6nyBRfQeCc8yDebEvezTWzuBd1jEyCUunnt
MxXAqowll6ycedvJi0QJml3+FIhpMo4DYT6z+7UzMQkQp+oL5V0WxUaYxVwi
Ovaep/iScDeT3lW3DoWeqJlSzC5pQL9xIKcD2OI0HrQvY191bZO/vkfvRynO
xMtaeh0FTR0RN4m7ASJDAggPR8iunpDmXSniPol+SUM9gweXCh2PZx/Z30X+
WDwdjCuaAXS2r7Cks0f74UCfCGIQC7/5hMTLT+x2U1t24sKq/FbjElpJMWca
YxcLZYtMPOE9SiTRpjVrn8az9UJf4rHlNwrGM1Z3kVBIFUZDSAaDLX4OjnXX
zUb4ki+BxjL4Kqbkw6lg+btDlkPn6PmcNh+MFa/h7KU7ltgq2P/AVslTY3zH
naiOpiqr8xludPd42rzY3CJPUoInxD+1m0TFOBQmvmbWHi1qjg4GWANuvyN/
oYbnuBlCTiasSSGsbIr9MROjWNkbIFF1wP5QTnMiA1mwMTEkLKjlhppuT+yl
JthEtu0h569QFqoNTbHIi1RsvtcAfHYMyk6mzP6Gz9GOPT1K134HH60UoekU
XgTkjVS2va1qTWfYFutyOAC6V+Sp2QbYsVJ9r4pbMgIZRPp9GH16Sx8nghbZ
gscBg6HDorZhakC8p+PkU2wqCxyI8NpqHoABl1bLI80Mo7xaO95V6ZtpyIox
1QuLS9ERenBul4ajieugGB1Qh4GzgjfVjGBSfqHbIqpH5LbR8GdZguAd0ciZ
Tc9qnK88VprA1s46xIJLtjR19CEUTTqaYWdTUMjdMQSmVbifM1kVdlbj0mr4
ik238VJ5SrFHiYxCPdW4awPZ42I3mlQ02wwyABa4Oi6pN9byLfE2vrFsi7KA
ANX44XnoQkdHYlrLcTjQFcZPwp8PjoIqYXmaBlC1YcGoo0NmgeuSGQO7U4kG
5XJf3H684y5ue+rNJuccS/5JuKvGpsjdTVWV78fht31/1m1Sh/N2ETrE/F9x
9+c1JgZcsuHSD/Y2tLYXPixN5ezfnKcUK9uDgA31oY3guNw+oEQ896EgHhtI
L8L9JgBpbW/G3GqULGNKUJU7t3g3sTWDzMZGDRNFm1IMiizr5CAJBOEBoztW
LbBRTNkYLav8EZlG5pM2DBBh+mlsvaJ2E2NZsoFSc6HYldVcw+rkw2uVVr23
iKFKcAOF2O5px4bVP4xMZf4J7RkPhid3Z9ycbShuU1n3nr3UUJIT4/Km3rcu
mtnI19ViyZ7CaPeuQGIOhab+mPZ7EzHCwT4rsHjJ40w6N+Y7hY4mqgmLrtGD
fsijxVGpCSaz8RLZsDbzIeLAv79IJBURk+C6s7+0eG0FGsUfcMbJ0zJG+Bc7
C4wWri/sxfxmgTUaiGP6q3X3kGXY9rC8SZDuEmbNaALbOQX0V+Q9CqASfX3c
cpx02m+6Z3O+KOcnr+9cn2ktU9wHYfJrY75fPjDgUBgNI27f0jUVqhyGx5GI
R6yDj5W9X5Q+2ogCpIMrRZS3RA0VBs9beXNFOTeVqGL/FdJOk+LgjWIlg91z
MbYFx5U6ekLEx1PreiHLeDxm1Pbl9axufyMEwp6bABeg4dXCOMub0yj9cVp7
31zccch5xFoRD4NGJyJSRV6fVqI3416IKHXqzu1sdt0PlcEmxFeR9k5WyOrN
LSQpjEukqNNcElSjVvKmCvOH+OyWdMW2C//oFaLieB5Ty5BzdC9fwYV3eLyo
QbhUGVa5EVl7nH8xEvYGsVvJXzaD9NMRA93/70aKAGA84hnuO5yN6ZPsRkMP
au5EBNqX3ZeApdzE/utQ8/FzPdvBnvvcsiMUAmI31X8DyPaGTXE+HkBCxUb9
pKvMANE6kh+vPklQJP5zxw+PXQQvkQaVQOwsxaNukWz/LpGDyU8SWPNY5gca
1bhqucfM8Yz3FHPWDwvXhNfBuWAZG4MSbgnPiIqZCup2Ta1OEEUBYFRjNijU
rI4u169b55Ao9o7LjY5/wG6iB9g/n3b8HQAEs1hLLpRjRir6ZRrn1ojPPyMB
xdH7OH5Iqr7XdrIN51v38l2B+zSWQNDs2YS8KoXNbZDWqDv+EToJRX+Fv3d8
+MlIYl1hugMHTMApMS3PzpjImZNV/lHcS4KAGj/9CEYTzUsspSnE1TVZgsPH
F6axiQpMWfFHxfRtDHPByw8+sdgL80UJpdVJJPIPNHexB7IDjHLuNEau1/2b
x0jMpjz+oIHy3JlslKHPUROqwS91OrDHEKushmNoebdel7AnnuG29mUWg4jt
rzVLZn8vmunkQSw5Cpryvq4whrAFhp67OHQA/LndP9v6n9C2IF9lWf0PCqrd
K0WDbdIHKtYPHOXeZVZ+d2R7VvjMy9aqKzbYlU/oqdzbI9A4P/cI5rvMiC64
7Nvz7eBXfae1tyTnECnwBjK2B+iTj9qcIKKMVhn1niAROXVrx+pCFFY/CcXo
SnId4ofqY/UF3JbZBSJehYtL2SBz8SA3CPX2R1Mk1IRdHS/TIYTiwkH/fyP6
JrtFyhYTAspjqXRpfVd1sNSyZYMnXNipKFVP4tIgbC6y/G0hS2QWk3J20UUx
dk+SN+0DBahfTm6HTkUsHkDSd/5mj5yvtXsR+F9H6dOse1Wi+9YUnlcEM8q+
kSm4ugZ96XwN71qhTtdfmW436+bxWDk9EauGPutN57A/WZ6/6XGGYW4qUAd6
wCDBicrfn5qpRnccA8ULxKmjNB8ae+UDRfi6wYbba9659sWvTVSTZG7hK3p/
IUfl5EFeuKCRdPpevdjhAnQxjZFCLKrfjcya9PygwMzQyWhVdCIkcshDA1/X
Wxyc30EcJlpQhmedgwRolpvzRYobMLK1aV42nLADefL7ToXdf8gevz2iI6L6
k13KqIa4zkKt8G7HOY7Djhpj38f1A8cUCFBDTMlBWhYpY0Fjh5/KB3DMPEK4
KVL9r88PG/SdPpJb6NgbuCINir/gmamsSbryAyCt6dH5aXxsAnpn2WSqFfbE
IXwsrYsAXCeDp36/uoabhmzRS3FvvyHPp4nMHKz3wVpuqFJPsqiwlSyA8bD/
lJFhDaLvpLjQTaR1z4M0mzUVEGrmSyLdYOLePRJTHyydibbgTUUJ/9ytzC5c
MYsErDAgtFtpvuKChIckS9sOmL/7uta21BTrwVrI2zSwlO5DyBHNg76+YIK9
j9yAjCg5wt/3RovRsya5UZ9fuKPod+BWFEjw9PTEsFP6L6aDGWumLlqxFFHT
1CVYc71zakt1NmUPP0Pncu7Fjcb2eBgVKg6mxh9VmLeG4lo8lk00WsyQiAlW
jyBAHRd40h2D9Ltxi6H7qQhevng2bUGRz9ZFkhyKz5ge5EnSBbVhQUxsjnps
/TlQBYiP6MRt4nxZYaw42VXRCx/2+djalDlc2FRmFDcLN++3kIT8qCW4eKHv
jOHT0mnxiTqrLI6KvKYqCnFHMcdWypZSrQK4yZjLjhBNcOGI2lX0CVi3tQYh
6ZWGNG4V9SxcVEXqfhV95xE/WIQh52sJWnfs4n+SHcue9LOcOgMS84n/7iGi
H35iMiSI6YaCZi1998Z7+rD82N8IC6MDGlAfjyG2J894PIuFLrZl6ds8+n6l
8O9pkQX7p7epzvbEGJ1dSmHt5ehPRFH1lgLsI7mXMKoQT9NrmKRHxSsB0ypi
+p7PIWezXcDjwSERnZC5VV31vymx4AiYMjhJwevYR2ekV9XJxDT42SWRsqPZ
afpIsGB50qcaCBlS4gKcr3xQFe5rUXYBUrFaQmEht3BTM3HmJ5la0XVp9bH/
ckBCp/vJBfnOXw88/i3ntwauEsZe9y6+jyybFz5UcgLxqqo6w/5airJCQMgF
GVMiitqKSCdT690ll8fjT06LrMts5de++GYYqvabPtiVB7p0G0DuXGkpsi12
Vp3trMJ8eK4A7/0MpQJg8BwlI2APDIvOAPfbqejdFrsomuLk8/jalBXZSZW2
k4BHCuKdqEWEBp16kMQgoTBh1hEjhyr0GCz1HdYrP9vugmC6G9vYBfDgfqJK
1zh7O7SqApNw6FsntrUrFOTLNkrRQSJQPk688+1bFV5SWbp3H/9ZbZ6/6Uhx
+t/HvLAOVO7k/R1sh69CypsObuyBBPfFB601Qbaic3M/zLFHaslnS0qAM6qe
yVuHNTM4kF9hlew1C6NVr5fJG7UzHszQg7y33GNrO6Y4U4fIllD09/1XOg8h
gvOc+NXJEasGV77UDTWS44UX5EWvl0kSIlKUYdiOfhC/j94JrVicpbb3BaQL
lDclbq2sxB7k9v5hBfRF5nIKlps6JsB+txKNEkl7EnOTRQrDHzImmpPG+bLb
1yq/xGtRYTij9n4kyx6d2S2kc81tx2RUut6RaoUagY3lD2fNedYy3QBzBfO5
XZHBjp4uWvHEy/Y4/4qMlPCcoBaSEHG0h0YFlj4Q9iT6l3coCxDLn4bSahNb
s4bArpoKjOj1bbpTtoNLk/Nrj78BsEs5pIB2h7ft4PjMhjOKyzcS3qhm01ep
Or99jOxQe0ivY3+LBpx/bOQW5PZjB+YeWpKM7QpaubXch7zwMM8I45AKT1wV
54gsx2NqbKwwjY21eppuGqnR2mlgeE3BaI7DMC45QO9HbvISGwIUx1wlIjhn
7hyOwdXBQ3B+zqY4MLzZStGSl/GvK0xzlZOPlCqfyBZMQCWsJwZl+CBWf5A6
mYv9ubbvk6rEnLNlkl8DctkqBFJ5MEuMhPtMXb2SLHbBOLpCJVcWyvgpR/i+
kM4NMcoo7D2wf6HEotsVp8g5ayklJVS9ObKXBpcOgUFMdaOXw0tKD5FwDg58
2N4dC38mNserRKwOYuTCQ4mUjQ3xyFshbigcbPeqGo0Aq3hrF2z6f8HHFnwD
+O0wUIwfq9KmVfaLIXV+hHvaCI3eZxUjHs1fBKGS0ZOyjbJumcIt+JD+DB7Z
y6fOCMS/eLfu6aY3iVcknEuVRFDabwn+4I+s0f+Fowcq+bWtd7kJdIfVX+cM
WCMv+2jNCHgqQYRQEhsh/ptjaVi0SazOrCmpNjyrU0OQp28mau5pxKhOladY
Bpzv3FG9E8eUsqT6haX7YmwcFexL7RjDJKUDcpYGXPuxXyFV7k97f9T9eC5P
M4GHC2RIc4mCxNhXoXemM2dQmQno/A4SIMfIts8/OV57T7HI+D7kMLRvF9tC
kAPji2kT0jjsb+ewtO0GRezYmmauFFqEIZHSVwSJJtYVdDbStzsks/3atGVO
pHIiNQC8zkSkonPeqBsKdoBvX0FBqd9i0+DdZqBE+HoSlnZ1Z/1pTiB0MNlJ
YyHFrd5porZENbIru6hFn/RSF840/+2fSsVMj9TeleIYw6gf5JILS2FEQQ07
lN3ehxkx/frZ4oBD+vdLoyHIKTo8lgYguAv8VTIvfOnEs3mZlS0mXCHd8rQh
TUgPdp78XaVKJM5EzsosuFd1RpHkdyckySu0zk5jdiLgSCnrLZn7FmB+iMZ3
fgiB8m43fW4swN645umaepiSD41XSsv6sJSl+0NosuahjLbMO5kEbTkXj2Ig
kL3C+u8boyXQ6G3GaatESrRBNVGK4JygJG6YB3eCJ/RuSgU5OxRZFEiwHxDZ
D76pMmdOaIC+kkaaDYw73fCHb595dyXy8Tfc+R3KI8Z/iI8SAQr+niudKeTo
j+sVnn6JaQ0Ndl5EKFiDDGziFsATt50ug7pGGpJ8AxyG41whSlDH2yaqqwge
yF46dFVCqa3lqNirri/31bNFNoN8DKGUHjNoWIyEH461B6KF6rOj0verI4tZ
x/RpTfL0mwAL98Jm15W9B4CNijsteBFX3qR6fWbpxkwakbHLISj0y1TYa3e1
GWVBbL27fIHt6rpndoX3quYI1515dAsf86BUMqwl0b4wlmxCI3W6/WRCjsor
8K6nL+gEfAgpn8bQg04g7H0xMy92OdVBYNVdsmezZcWq6ooPaAGELKYN5quD
ygrcOw5pyNKiowjcuEAw/w5bbhchSokFDABfFSm5cvi7q42jXNTmdvJQAZKP
HHreT/qbtoVXttjRf1OLXbCO9P78Lr47+lgwZjxMtIMB5xaA+CNceXdzXJ5o
vfScgJUxW1Q5iIvrt3QK5DNiV9GuK0hFb010p+ZPnzZL0LmpgNJwKgsgxvQi
HxaNbn8N9ciYu9gQ6WeberMwPg2oV+0uvUpjr+U9o8MhHam5nNr5jvJHYIUQ
+u/faH+CX+rxAnfMCYeryzGwZBkMzanjglzhT0TdHYZ6e0A7RLm/wLEIa9rP
9jhRVBHVseQyn3gXGzwpZUX2Btgte8UeVC/jGOo96o8+e1KIA+NT6fFpOPjx
+kR+4ft3DMtxATcA19y7W+dCVRlqeBeEYbvXshjB6RPqoyfmhOMdZMnEGFMd
5Vbe3MVOJpAQpWT4c2PVMGGtOAp7GIp9728SyOdKKqHvLgSXg4X228yT+oWp
5GkTwctf4FaHTyI6qMzVvUpQWx3TCWnIOC/LNKw1YrodEyyEOYmGNrN5AsqV
orDOxdOQ0Z0+pSez5aXv4LqXBNag9+AuXy3lAtYPKYh4n4Lce9p8FHg7O9IQ
7equ8yCjKBLX9VfG8AVOMhdLcxguNIgyaiysaEwutiSHszCHYJlOzQCrxGSL
NKBbR2jKlGBHOYJu7lHidZcLMTdA1FOmHL/8CGJETcCVXN32PV4zDXR2wuMC
efnboqE7ep0Mrb8XxaQ3NCDBmKKNeVtZ/YaNn8J4At2LO+4haqTXfYEtwC5K
SXmOt8dApmlQIPkEnVtz9enD6fZkXrDUxsWH7onrrDRYPGQObB2tOpsA8iGJ
gUGQsXUUcwhgHKl/1dV6zmygvMaj2PrwVIStUmczojO6T8eO8FP6r96iYRNm
m+zHc5l1tOAvv1BTMmnbLOnwWcB/E7Pd2MEexu5YINguzBeZbDjp9jFAJ48l
N1DTQs1NXQxYBRB+jLKaVRjezPx4oWrUsr/ctxU6Cg1E2jBpZBraMFdLBUgn
/5B7h1x7tkB2ZiINnLX5Ohr4Jqg9qEe9gWIBMUPTY/5PuxWslO+DYy5Uu4tL
qosMIlhugarJ4RgyqwOvWVMvE3bvq+YVawwMZk4JslzqD3A8ouGp+EMDdtk9
iKQ+rlwLRSRD0cu1MIXv03afKVwhASBdQv1QQrOd0Am5eFwcLRr5TCzESCC1
5ztw9ROh0ImAenfK8SybQxpRApe7W1B+c8omzuAz3ntHp54KNpedFuIjcPM5
3g19/aetLqNgu4r6DZ3qmjibuA6dVTeMnNcw5MumuJr/+sQs0Rj88LmYnxnx
rYrXGXSnQvRYebYX9NO0U7v3a03qrCkIuVCq3MfxC+ziretPApSSg9IKqPYC
k+tvopcdpgR+m436Qji481Gx8sVOXYWqQBbUZyHf2kEz+cttNB+ePAGfrtVv
QMszLhL82OPuI8zElmQiQVpXfSYSBwnX1wD1KceVQ9JdTz8qSF0WFxuHNFoP
P0G4QPQHdDg+Lsv22cP1uMNh2mYc8a08+xGEOnTwLL5Sav2W6uWy0+hU4Pap
i6ZSQCJUddURKGSJRjJnX6Wm3qEM41zqm1tCpWk0mSpLh+VcEY5rCznSbkJy
ZqhBM7oRSBHf29zzHbHDub+AIWEpcLcAzac1a2gKopq8Qx3EYqEQuS29NWpt
nNqu6OmlOQaIEzSRrbw7NOo+CEegy/BAQItDf0aO+cGaXT+I3yHFPA423MOI
dmWOBbbxSuBx2LqTMsn+fwh4JjLWtnosDK02DUdAkhrFfz4JGwzsx3gdUCMa
CKFSTSaCVKj18Jf+Ftzwa9BPENuudkguaOwQePCrv4ryMbDgnmd7l66B+/0a
oQxy01MG+6siDSmr0ekGcoBofIpbk52DZWLjd0MeX+WjeUDy4gtiZYhMqcq7
LU3SUW6vUvWUgmuFNJdE+3t4sAsXqSMmHAk45W4+ebODJKTK+kKVnpyLSBdT
EQLskVjswnoNq+JKLWw7kwHABc5GLom0e/9cpKuyZlS6QexlMJleGHGIKoxf
AB0p0pMbZotqwFFuYLajR2IH5sIa/LuAobUUldiL3XXAJD9XhQ8muxrijRQL
wDd4YBlPV4PAyHRH0/rjeLCnW2W2BdGowJXI+9WJQVzOWmKRASiAQGjv+C8Y
V2xrqsCXvarFJOnhk3ofoNCRcYBGy63o5FKGvY/iZHRIwdhRsP8ITEqfwdKd
ptKz5fYx4pRNFdYiEO7URc92TfexTJVLPHHBl8XLTrQEGh9lvyh9/jj3Uxpc
62jh05V8faLgKwZOvEbE3s4FeB20vJ0NLd/hMoC+Vcc0ydG0tF3qNFEWAiMx
hKzelKm35ulkQ8bcHFmRIq6bFHuZm0oDlUTYTVB+BNZB6Q0WMTsqJyAZkZA6
IhSkiryJnjGd3YnElnkAXTg6lP+e/kc9Rs2ipyV3Lx8mYPFSSN3o1h8mM7s8
GYW51/ikZYUXxjpGAG9WIhX7J3MQvLRVPa6GzoXEWQwU5RWpuL9MritbAoT5
m6mOEurqVuhnSuvb6I4dv6YVsDvGr3WgEfIXoNExFNZ/pIEk7qmFMwSYd/Rp
mFvaJlm60qB4npNzrmquRjmhJqikHN9VnGETtHeHhSYtezTdLtBqGwdIdvt9
z5eNDm6cAfGhy4/veVNTttWAQKPAdCVrEKrV8ee7K8HFUzvffLZrJ64CCnak
n/XsbegwzhlFk5N0j5Y3zA16K0SzY5C84hzWXMyL1uJiq17JMqxH0/7i6eWp
PqF0HBA9q4cZ9LF9Cy48z+GYp9gNuV1nW/py1R4r7dg2BYjFOalqNNXlogdE
gPVkQqLU5u0szPFcrdXHc3I/GNU+zRM54NB+GjORmqbHmHwGbnxLRQfdqZS5
GqT22ug91hyNRKWavvPQCNqOQF8lpdxSKFLGXzsc2uVM1sBSbJC+Dr9SOt5W
611Sut6rEz8/tDIQ2bYU0b3g7gahf8ya57ynMTvmR7K6DUGcheuHVeIta7XZ
Jxkfv6avPJ2qQ+DJtAstkYJL9hWH0oFcA7SAXzY96y4l6N7ag6BStVCDqa7z
dnbO8jT13DUCM/NShJENybY/oDB/vR4oW2d+j1bff47lKN9hoZpSaz4RiBsB
OHdwQk9E3CUo5EILsjN7nd3xd+JQvmZHKZN79EfVtvlr35BJ312YUFnnZSzF
UU/hHjts3yuCPoP6ElCTXYIqX9Q3Y1z4dbZpCHZAsjRKx8wCq0feK4W3MOjo
88yY8WS0hygB5k8vycplM0fBWwRAlannpxKYmeLhGVeifFrKL9eWgSugbPfA
0z4x5712/772uRYHveRf1UJZVtHCig9I4xjoSAZkku2QDblLRVXqXyE1XZjk
OzPnCyYVyLzVNYiq3K0EgrneiocX1n2ROlNYzH2GXYVGrrcLg7yx19f0ghi0
fg8IIp/hALcHgPhMRYRsTq4W+5e+eC+L03wA4ZggtXZB4Mm0LU/R5DxqfImS
/xmLAkrTbHsmEbQiOc6Ecz3xa1mGzRzBk+sO++wsxmOJxebOzX7F+sQ7Iioo
q4qPZT5AsF1DdJQdLt+8/NJezEHCRQ/tjQUbMVgfalkhRyH6WZ50QLWSnmHA
cXKgvk2Pale3X57iDDh2FKMnrSldxzwW2sItjqltyvwnLA8fF7loluNSA3ce
i0P/l11w5V1Hs6GEgSUehyCIH0djReip0vr8d6miinQnuup/enHJsB0x2sV/
CBZi/hZVoQKN/EBXvR5Si+WdPzQpFCPJhRzVytzFOYNhHc+kCZUFYKpLQMEA
EnIH8l0jtKpqvM8Qxsl5uR1w1k1WlIkqdX5e1me5sqX68v6TgaZMlMTyqGJ9
C7M13MhsCz3Qz+g+88tkkA95SFk09lmcCE6Y1vaPCsNeCFAkLzdUR/JOuZ7B
JqzNoNnZIVYiYxvnGc3iHtFnymexYmXS1JINKSkTRtvopdt/BDNCtyFEV2lB
ZKOaRBdVNCNct/Blg7FNnSNfFJbq4971dO9Sv/63Vhi+6ogOAgIFpeWP5Df5
0Mx89nVbZrLDTfSeoIU5D4z9cG3GCiLUoWz99dYzrAaISgFO0V6lzGb8iDu1
XOcSEsNGWa81THDRnEz2T2zO5ityYNRzED4QaDZ00K1xFSv60aCRFqM3L/Cp
MsfBRJlgeou3mn09T8mcY/srF9eKQnJYG1RXkFzyq+gXFNAA+s+7vGQoNyIL
lYYv1KHjY1tHWd6f3gnoUZKwYhDNuNOYyKbt8Yps6Xg9qafPUyJvYhBpvND5
uqcHu+7uX+PAbIIewiz4Qg4cJWgFFG2LwSOmZnYFM1bwpj/6MuPjxtKfFR7V
N7EhYoufIoNmSKh+3KbUSwPVXjIQX+U9+rllO4HehspSBPX9Cls9w4DlSPAm
LJriqr4obm+tBV2uaxDva7rwkCXjaVOpLibT4AMyI5rsalIc0w3zefhfh15y
wTLg9NyZg4Zrm9zegN4ESqGTlpG0DUBaQZcAjnMYKikww4/6lcO3GR87vtVw
iqqx6OXuOsCyvNf1/fRWwAIwB9ejeaL4D2ssPOIJbhUwAS9j73m4KpS0F8Wn
MuRE3zJruknPgoaVrVd17aa5f1GG79UuJIeqFD01ENU21BPLvYS+qQh7wq/n
Cgc+u6xNPJeKIJXRRnTv/kcdndrtsGi7+mdKusUPghBGSdD4pBNEHh2dzSL2
R6t5M15uMj0RC5y+qqtr6OTW8Zq2QX/3juGWsbceHr/I8RHgVUX5eQa0FPbY
6Jxs7rxbm8yrniXazD+W7pV2VH+Nt+jcmqoLdCrEncGz2SwkV0vEcEHPzblj
iDQFJgPnNABG+VVCFUIM+35WrJhATnqy3UWtZSOMUoV6CF3w2ILt244EyuKS
+bY0kpGlTVsVN/byNrphOrHB5cZ/vQ64t3tU8qlGq1p7FFIcWMRpdHGG4scr
m/QxvBlMRToyR3RDS638R+/8jzGPNvRK+xrluFgQw1/xEumGu+eaX7GLQuKe
eZSdcv7stPx7Ls77jsUb+Vd2oJWIim+Qeg26pNq4438GvZXEnqC6+9BSO5EU
HwYlY5lpumAtH7AFSP1++xgY9FUoX/nzx97TG325m17r6Sw1EVAlC0ZGbpam
9l5rUjkDnZVqxW2n5oRu3/VHDEhamuKSSpoDubXKy+IhwbN7+rr8peJ40cVt
jIsLH/uvUZMJIIWmf7phynLon2z0pP0BCRMkv2jmC8fmDkGtm9ms90aAgd/M
NU16Jp/ddn0vVKLRnoAToic9MbOnc3ArTE5vELoBmPeZfXw0BZZ0a48TbNWT
zuoCPxwa3iRMsER1aGpKtZIKO9Hcwjb9euL9i/1efMmutZC+Rra3d21OD5kt
Ll//FOEJxcWy1EbK54KlpE9k61cZtoI23b80oTyxvAHUDxZ78mfWdCSQODgR
cqtb3up6ylpWKX5t0qr0/nSnUT1Nv5+JRg4xY5HMEBokzz/YW4t3pCrccDuf
Nfb5Ac6EhL8LvN3y3FFKhfpIBHr5vu7ftwpHvaI6FIHdIgzpP3pzl0JrHMLl
SWClH3C2/rEc3TgNrPrI//c5BRJuY58Dq2dSrDUvI9OZrzVeZC/5bTrXo0fm
JreFirShIewWenmkcJ9qZBvD8g1MOLMacLc9awggx0E8QkJBrxcIzE+DhD66
kVF6jdLnE/tjbUlS7QGoAASeFesLqwsf9BVR57UPywym45XPwVbQyUKMOXdy
vF3i4PCkyemqg/oFK/oy7fsPGDy+GetEBlp3cyAwnLG/c5M16WXkJtwiBqQ1
5HSmknCGgckPYDBEs0NPw7Uo6Zcxh63vcgk+RQSz6nXRm/VXV7WrJ3iC6bLp
vvOOQ7MdcDM2vEvn8dsQJTAdMrJotWp18/RxDTUR4N5J6uWxaQELaPoGd24Q
9oxumm3w+RcOa+FIya0fji22H3dMaaijqUZq0ew8m4iaUrgCnfHgZ+8c51PU
SDl4B9MbVpvcbPdsdW4hATQCBpyVpjf5Z0fWCWbtmdWu0FYUp1IT3Rfegqm3
i9jDHFIEZEkvFWZv/gDNQFrZr6nzdtvVjzoQvAjWq1DR8OYA9SYaxZsB6QeO
A5bOauCz6tl3ivhPJ5ySa286beej4ZZ1tWPINvRDe6eowo/rtHwNw4FiXpG7
wl4r75+94DmcrFM/+4+Glp4zWBUV5sWx/p3QaWsufe+4KxFOa1E86gloedXW
QvsQhj95wL0A6w6xrjVT56m+hWTVnEH2GtAyZ9gCIFXRFYrGawJ8qb2thKet
Oot1xZNQg19jvEL/JXqYvtr4m7mLcAzyOt372F6KPSnNA6zKHR9dmY0AZ1Q/
m1XlU35HMDlIV9XBU3kUU9f8OeH7eV4u6aanQycLkf5HSE71aAfZwqUbdSeE
iIo/CwKO67KV4NAipOiysb71ubUbsoGFu6+voE+ZWNTxvOjfKdUBFu6/ZVYi
kmFHM9uQZ0V/GsVhTL/lWt7JQbr8twgPXTjWikr3vdf9BX3Pf9+lEZFUNqJK
keGj2e7UQWjT2dGp/7MtYTYx+kh4uOP6mrkdA/76nhIflaaNBVTniQk9oEuy
KCC6h2Hnujh8qMmnXk5ToCZ5WxDaOFkynO8GDmSliF6518ROMCc1RKg9g8BU
/pUA0gfAUJ551C7v0xCevxNXLB7HEQNRS20J1F9k7Km18dfYUYLN96fUQxhB
/Ed4vgl9lC9ulkKtL5Z0YNkMEF30PZZ5jlvGzwsGVq6oMC6AvCwupBMM9Q4S
HKs2VzpvzLdhk0cFvILRIXgJPdDVTGZrcgiUZGLaEhA4d4jk0Kc35suSYN1s
0EpimC0qdzFh8nzYPy7LqD6n3FuEciP3MUo2cvDkBh9vZuXCTuIG/+IP6Yih
k8FO/LVbidUhgjeA0QIvUOd8oX8QLRuFcXUZcj8JXSpRQr5WgqOLZ4m3C3AM
7e1yoTDPKW/NZCkaNRlKcKXd2z8j38GZ8gyJQ8Z08TfCFTPULWiCvmwXnfAn
urPaDPgetKZZmx0ROVzNQcs242Di45GL09nFuTQjveUFsr3qoeIAr0vhKnCz
ULD4nnMO7a9CZbWsaFg1XtV84gekbw0u5VR7Y27C3SPNwgKRb/rMcKIQMDiI
gj83nZN/otR2gTy3G8L+d9Y4stkInNERINl+ey1PJQO2U+R6kktpbHmgE+BQ
e5uhxodgobK44BAQnh+w/LwvYMqlaOdnskFxH4CALmjq0ZssQAryi4gs7fFP
zdpHDubqJ/NvM3i9JCiSJSzlbH/yVtzlktv30KvwxddAPwvBDuqSFLbQkB5b
k4UTZlAkhkfDHHzUK6+E6rronE6k7ZqBd9Fa33ND8NJmZxYbquJfRdhVoMa0
0xzDpoOwtQf8/cqWYIPD9FOC0RGweZtOAt1xsecURbIlm5ErpiU9tUOYwmC/
BYTp+vhbk7Ir0z6Su52dx/1R4a4YfMZWpteBvglrWdFf8PjFqpN7d6IX3OwN
w6igt3tBmZk92OvJEIpI41rJ5MQInz/yJV3e673RdAa8lxWu6g6k0OM+NCyS
+RkaURbTsQZz2+o9OB+tQilhUioTwwkSBSm+WSAviCgbMJC4oSgO7oI2Ss7j
Oxx3q1NTqA98XlT1HKZi0Xd+Ff20q4CvxPKJTUtBvyOENqcMFMf5YsaJSieo
FUrrs9Wz18rGouTmaB/ua0kQwaGNW+AYlfic9zogWfaVVGkCNJrtHOaPQqMm
dxebJ08qf9/nkVXWJTU+ORwqq5/qa7QOPy96dCgtHO6DoOIoSR1+Vq7WRaaO
kQdwmF42gJ4nq+oCo6LXe6FkFweSl8J2fKnUF19g4lamzuN057PbmGXlj4NT
o47kwcL9dhfvI7RlrZQf6GhjJZO1ajllGd9hzL5oWP5gx6zmMxL3DnsvtRL/
uMGa7AnbqTbCIxXsNoFHQSEFTyTg6mvM3z3WQgbRyZNXBPRoWisgYIAJxSip
OuStjNt4YQ9NZG7MjXnov+eAIRxB6Fw+D97XoBtylSJK+lTU0HB31Ad6acOR
KVzKxaLkuHNRqPuD77JBTCpKkUBL4LpedZb22mZmvuX7Cu2oVFESqqr+nSB+
SUyldF7AlZtep9jCafHEvjbfdiemoXyuGe/fCcYu713bZ47aJ8r/4qp/Zwyb
nZpwi1eUl9xQi1JFohNtlMEtvr5EX0OffWLqkHX+Zc4y14dQBVWkH2udDHvD
QtUm4VU/qQYQ7w1kghQeOSzr6wTOay3CITX8MPjsAoZgcJAK5/5kPBzxoZsQ
1SHL+iHlCABBH2dJeZczssbP/QJ6Sw2wIefbEgPrGV14qKBWYZQN82JlrIfc
EtcKEAWDhk0FefgE6K7YSAa39yKn8sCuwufpsvY/Y7sB5VgGhrD8/ueWQltz
Epk9cYuK/J1h3Ic0sIDFEjnXk9T9l9RpHaCPLAs3leXWn/CSshB2OfOCrMty
HBD0lhLnoQwmkOXvBAGzJ4hXBt52sbFobYZ7hl+lqg+N8Dboa26s6eItHgfX
DbriM4aU11EzHpIPgHi59k5RsomMpEQ9d56X2a+BgtBwtRP1pkN2yumUITUA
Q5YjfuSL74nODPbvpJOB/O9GRyMBg5D2G4gro4nHSTzUBcYGHx3iM3v+hVjf
NhU6ChjU2IXeLhm/fEPmaEX9xvUuju+qjdNmKrB4K/9FMk8d9VvYCUyftPll
n+76rZgBkQ1FtJAgYL6t6zNJrz2ausOVkjPC67fNf7F8GM6FrBDARCY8vitk
N2z7KZW3Te4CTfI4UNtJOmiCz+ZfbmAuYTjo7kWUMBSuW3mzBcYuyXVl/kmP
s55aivvcK72XNDvhoBeU86NISkaZ0qaiLa8gKSbEmOTqqIYG1JY4exq3rV03
NKIhsuWQ9ktJqBFHQIPOdBJAn7KUNfOq/tfMQuL6KcnJgyhCg3GAuAWIII+E
vjzZ/zSyTQVyKANyUXR6F1+dYNZcp8dxqqv3O227mk2MER1xBT2j2cUd+ywQ
DoP5lIWwvSUrL/KE2cz5co+lwV3UlPY+s95yvmOIlIuoPip8Zfi0ItmngWjN
vPyACWUtTJU9Q1L5XNJRc5DXh7gieFMpiQ0GxacUbL2PpLL4r+FW6zJxlt5f
Y3fbXWwuEFFkatp0FvQzbMw0rgnU3mkh9e2jktp+V3FaHm6YQnXh59vgkWuG
71Gl7tidZUtMwQttsoy0gNX4yQQZ53sWPuTAEzBXjbQYh7wAoKFZEXb/D0ql
RnqHKhQ021F6aMHwa5CHQNGx6r+qGoxhIJ9mK+2JSX2Dp5mzE0nySb5lXLBS
tUY0uDaqVSasEvBrlseb1IaKnLd01iztAcXrtcnERctaJV6rBwlv57YKBCzg
g75dJ4D7Hr4zvuzs1QaDKAhARjiK05UXMlOa1ya2FMoP+Hi4RFU18v6+4Awb
dfF+sfiD6sB6dydsCcfbnCXOJ8OyoGg6F0nidtecgPBokry7lVbSkcW6f1f+
Zjo9LWwoC+xWAiChiIv55RgbQbHfOkonSZbVV04ZcYn9CXTSx1rlMZMXHBLt
Gu40AVee360w1Af514D2R+9j55FsnEDAy2I+QO5O+7mJV5KkcrcLyLUnzoOZ
VVs9pf7P2UzuCX80WGsw6LJSROFpJDzbRbZGl00XQFbyI/ydbkFBGWXuCV/s
mGLC57ZSwnW4ntjXa/pMiiveuOSSFDwUAiGfxXT15Wxpo8pIxw7UABEJToV4
hxy4qfAyzpGsLO6i5p3g5hggi5GoGPRkWmBkt0yNCVVoog3btmARtUAZRfL8
W6K1YJG8lcW0dtECk934P+T0mwK4R5lSP63doOfUkkauIKPmmvnw1OMYWAf3
r58kjWT1thsQFx2zZIPofkqUIr0L0ZO/EpTMu3UlSXpuhId6rGKf8OscQUBt
pLyH5ET+PYbL1jiMp4nrZ85f9Irh5TyVRnW/k05eL2JqglXiNEBkns3b34wJ
WUtZhw1q1hqSy/scctUJ1vyXDI+XALX2+QtlubQR6tgEf83U7hau1Td2Pf0+
ZQMF3NkIhgy3qwRMqH7db20nAZdfMY4OUaQj+0cy53ALd3AkA55cf9YJqDTs
aM8YnLFqxnhuYPeIWSRspkQQmYlHtzR03PfBj+ze75aujYC57ZdqzfBbU21Y
XWQIbayhXw6Uki1fGqTXlhH++80O3X07Iqc1QblbLgMhq5I4fW3AvO1/FR8k
jnfAUDxV17swKP6ur36IgNNfuDaebFOlYfHmkWciUZNpgPQuMS7ho2cFUlQi
z+1T2NC1sremehkOvGr86n+q/gwsspaplU2xCQuRQ30kNFdWTUDW3iNmq7WC
e77/ygJZ8if7fPdLJHR8uGPZo6fWumC+dqTjdzBVqVJXsdiGQtfKFXtEjVMj
93h7KtAhGjyPaYs4Xdaka/zn8lL36ErIs+wr+Yen3Ds8EYbEyW2YIQZngbo+
2q7r/la5HcgIE+hn5U4Ksa9qaW490AWSvuo+/6IpaGTXYVBg6ggoItnymxet
TFK8c/xM5kDoCEoGqDAQpVEk2+xRCib7AC9vOx3iKiU/eYyTza3fuXJ8cSUw
5/jWayyILGu79ysD4/Q8jAULAAB2WkrCgfyOmpblBR/4pfG9Mj3eDmT0xMXW
zt818bFFD6EDHuWEbwPfY9aICOAcqOCQWl9ivzVRhkO3WknXseR1gK3VjEKc
kp9FeaMANJ6zRGE1m6olG7HO0F1EOWUGXjh/c17woZHRhmOnxz7RTWsCdkW4
38A8zoJpjinIJqKYgZ21Xf+TuCmk/vxLLXyw2SUw+Olb5g4L60IRFUt12lgY
tH+2stgsHgWJ274JKMtFM+JVs4UbqgMpU+1TWnMhBXEBJ40V7GiSOLav5/vK
U9/zOE/KtDTDQqB4BWGaSz6nCg9kCguYHXEzLHDa1K+neeeMBneaxrr3bE8N
ru19J63PI7o8TbhkYK2Jgh7w1diV0DFeBi5wqrKqbuk4gtYl4cKSll2j+fme
pZqZ8+Xs+Xy+0Nk8oV8dV1y4FxZsf1fbEu3Jryw+7kXw68Ffs21PA6mHY5Fj
JfpmeDEsc6Y9+NtxzhkNo7MA4dNCp1igOXJuP/Isri5WR0o80740YWD4f04v
aYlPXNr9BKLdSuOkmg2SJ0cgF7cOBJyg+IDYR24aMO98wb3lNiAIRZsq3IV8
HzxjIsuzQDxw1KXgklfdnRcxh2p65C2JDJoPZ7hNX5NyruB2dxtAVh6AEyxW
0m28+ceyEftYCaNxOtWnopSsRd/CqzHtyHX5B8PvbDR8v7wFkcoYDISfTuCs
6RHAiCERT7JwziKj26cRU/bu1Owvqi342IPLIH3dRNPtZBJ2I7QtW+7yoA7F
F0iUE25/M+AXt87TgGUyCWa6AiASnA0yxR2kb7EWxvkf9KXfTEpmuXPU+EEP
QcD/rcbZXgG26bMNq/pZjI2lhPXhvD68bl8ybae9GL11aI0xR2L0YVNFPi7d
pjOOMlwWCXlUB+nz/ipHhjCgh/czYawebixwmc3r0q4Bh5dw0i1CfbCsFCZU
6MivtcZ4sVPn7LyIcNsA9a9XtBR+A1MHaBJgScX06W8WispCViorNegfeYYC
gRVrjUVjkmiENeVJT7Ndhd1enctRg0jMTGJ2XWBnCrgkKTomiDxEoSHMb2Dq
koa2+52JEJ3qYfQntKhi2WGNjX3552jEUZVR0eWF9ISXcUYy7wqR7e+LCacF
t/PdM5JeqxeRltAdcmN4ZDaDp+iaGDTm5irlbtMF8zpdePFvIuwn/9rwklly
931hMfxRBx2urNn4oRRx5YyYnfLEQMU0fTAVkxZibSHo587rB+pBQgnJzUAs
iY+GOVmti2Jra15PxVeGzkJF9mAshOIcuDXTX46vkjF55QrzXCbMzThg84eQ
wmCDtR/y5zojj4Oymh7v5ufiTkVdlBXi4KfWYanwjhTgI0IBPkFGGsD50/TG
jFZKstPtXcYwnENnLN3rXw64qYs5mFhFMEoPpiGbRsDtFczPtktEpaLMQ1W4
ljwxKWy45nSgMhL2gRt5JV0/YfctHRCgtH787x1fz3YURUuWONJzHYrKgVMq
ALKQxLMVQniAhy0kvaiSZ2D8NbNVLMLjdn0usN05IhAIbub0zzxcT7Y8VJu/
WYz4dDL9iq94ewZiSImzrTNErHyhxlRghoCZgzWncbMljEJZKDbaqIZ09UFl
DS1cZcOAOgKpbIUo18U4c7Ba9yJUCZ17IHxwoxlp5SrJLkZF+n6gpOwQpR6A
PCx/e9GL/YgqHB+hriIei+wvc9aq13k2VaRjiwnH9qdKmJxMQnpFNUPuaccH
2zEvqY3a0E27VcBT3Lut7e4/PpLGU1/hAjEnkY1L9ND7ROqU3E4FXQ3fH6XV
6deiuLQXssVFRFP1Z6FKvpdBHjifzyErL56iMZm0UxnZbgbPKME0xjMM7MsZ
AVk1sZ24uRNTSpHaN7Cty77Jxmpw4FxDrkYPisIM2sfUPhWl26iVS5dSeguY
efsuZc+WKahlNrx/Dr2QtbJeH/VCBX5XZSjvJkSmR/UGqSOCuBK6Da6xmhmm
Ul/ihV6WaD2/YMWn20qQUP1jFxaH0B4pBzsRj0g39ozoS+tDKmeTOqO2OUIc
JUCtbtzf1paDPQDGp23nc58R2pu5ofThcQ/Ps5QJe4eHzCj8mcyFSUTlJTFC
IB0epqwilvxzplFv1D3dVS+ETvSYVxigfXDdLMt9fVsvdp5K2Ds93QvzhaTZ
2fwfwhm17R3XD14K28wZOrXIsSX+J+wSLQw0bdIiFDreYen+WIOphuFFZAGD
j12NQVbZPNTHrNZv3Who6fcCaHySkE98AxkPU+Zj/R3zGHsvdmyEMN9F5vc8
R3P42Gq9/wY8N43eQSqRctimVGze/w2qOB7K6OIMxiGoxBpIJAXlxkrygwrd
gr9Odov8do70LrPaVL34yynfD6ZzBjUOpKExuMH7TSY8GMSvwJK1+W3wiLaq
hTaFghdPY5NfeE+OXdvJsVn3lDTUmndFCMXcf/E1YVXTEf+hZydNe0jlEpln
gZL+3CYGLGrAAv8Xs0xOXR4Sa8ElGbcU39o+/R6Om54dA4kv+zUWDtmpbwAU
25D3Yo6fBj39jVyFN8vjhtSHEvoLyKUTgZe8NwzbKWArtxeVGDYzxUuFLCUt
X/Ji3xbEEbVoDTJuE0yQVBL54YiKZmTzMeEcjlLn2DKVX1uVJc0jWgBRiHP/
t/dMtWmUSeu0sw0iqDKtzaSJgxXrxZBSsIW34R/MpmuDwhBZF9SisDLjMWrf
ej4vo1GkHMwXulZvai+k5LQ5ye7cSNYlbmbu8mQ1t8ycSQcFlyKff+pD2M4G
oy8abwjX7UepcdcTegqRuK+t9pb1OUqpr9NH8rYWtEvk9BbMBIiDNORxhJP8
m+i+P3Ezp9qpFNahylPKNT9WFcECbbame9g9rWA3gLNRLcHpgO9Wlfw8FOGQ
Ib9/VGHLEEMr/kfRkQwqlY6ZBGRfy1ZQxCn97ZU3jkcl63WO/835JPSkYN/2
PcendYMyYpFCN1JJa2ajGgpnLVo3Kxj127g725f7qpcvWfgw3o/ApwN8lWCQ
IcL5LBQCCsH9dUMGSZjYawD/jzMnDrDsGdwqhHkzH1KORsJ0+o0E0EzlVU0K
ZN+aL6SZK96HeXkQdPd4ROY1SjKuV1S+lvgeaLwNSKf0e0p5inVS2AKkgAnP
8HrtCfGVi3IP+ZX8U2cxs24PJDyHsGWvM1mKnR7InrY3+B1nafkVSHXfPD0J
GQXZod6rrE6DV4xHcnS802sfhzNk9VNddekUcco9OSyVPwawKlt0LqDXtPac
sd2fgA0H4V2Fm5yjDreNU8NVjiYNhH6CXRb7TrPqqnRcWDqh9bsgGmRJ6DfI
NwwLYztMK02w7wrakzoL/FcJi2z8crjHWjDzWDRfXDzGlLfIsHiKUi1ImNWd
oz3gFBkdEoanuwsbaWiKHZ6YzdAFBlqg7GHcM1845AzX3h9GMRFwbvRm/mUZ
R3vydrM3aPskX/vJHmqpKPOwS2W/lsk6Gm0wv+hOzNQVExmrxZOqBSE/7tm3
srtLbUmHxdNMQUhiiTiSdvBLyJhdgA4kAO4zq9DeD7LhLm07VaS4b6Wn2BWm
GAVAPl0ggmSZUKcLtEVk17bBDO7sTtL0pvbnCPsjvJtEQpTn8PtNoLf9qM+m
WsYF+wRIOnVe1FmV/8hqiNpRWrM3esuewU04BF8pGUlRso9TOud2H72qZogO
yQWayhPnRf+dwVAjZyg5MagbGSgLdrf15UFqTbs78FMSAg6VLE8wc4dJyo8P
yDEakYAin3LoYbPCudOF9C5ZxC/i+4dkWn1jwkM+9ZPdkYZ9biwUfU2y2qIb
PWUEkcaWJ3mKMC0J7sZCQokc1K+7eQI+PBkQNnjHVylV8r55cgUs7+03D3Vf
8iM1q12Fiafcuogu0dKfSfBHfmOWFMEdM31SZ2VuGJeqJTxWjSN+DBjmyqCj
8XJwpf/zBbBZvYFpcynPwVuk60CACYD0IyJNPAfYULO9nXyG2vz1vhufSBpa
GpIYYFwBFbG7sv01Wraw02T7Y+AKsFJ9IoFMkH4tX1zQ+lr1wFUtptsVBD3L
3t0gndTQT2mHDVilMkE+DkS0hCjUeFtnKuYxL4/xGTVRFskj60FpKprvD3CH
ne8lhu5ReYw8EX4FfMKh9mPAxoPrSg564opLu69b2ES5sZZyc0AAQydQ9Zw2
ymvTwb/x3XKRiAyzFMOQPEzD0cyKuKig/2BdvV6IclX40eoGakkTZEBhjXRI
lvSo3SsXhKhruuH/MS/dVMXHstGOVdXI/FLrY8hTBP8RTOTNEm765PJnIU0d
IsTSYknobHeTP7V4IjfnaU5uM59iAtJ9Yqm5pk31RGiEFOlpHlRFT2UnSJr6
vDMvwv+K69zHWM41f+TBR8H+78CAL6fXu3lX307SVRV5TegraZcXLydZKg94
d0LdtaWHHgBEjdVOao9WY8F687ma84jrm0JE2ioZJJFco+voN5SKuwEJU9fV
93Ewcl7x1QiWiS3yZm51gli6u4m+KZsM16DBdpkL9TSw1XFvi7CznW3TVStt
sQOs9t3hkywBJYJQgOqZ/xfS3F/o+G8c6w0zeSRhQVOnkqD1WJIOkI1sdQMb
60jbl3eNPD6IcLboGsCMf8MxdKdvidZy/7c4NnJSIf+dioL4YNehX8UtjYKX
WOP7orriOu3TdPUjv0dW/E7lytpHi6gHmPmbaL9AGNvAP1plqX7kyhKMZB39
5q+JbEFj0ir10UHrQCKriMYsC/JiGNarqIqiqZ+9BrRx5YdJ8RsjK+EMyNKy
EDR+F5lkKHByJHeeEOwcUW5FWAfRUInmL39oQst274c1X7qa0KqLgC/nbRO2
w5/Ae9gK+nByvJm94u37NzXnN76sh+qRMFScbFmMtJ21TKEbqeukVFwxAK3X
jp+wZ2rC+k4wyn/IkuWhwnpQCEoWoJ+FnICHerED0IZjg4aFVFDq+I7miK+z
e0cHoQxarH63Y93RNoL67Ga7MlWlpg3doT56mCGkX0XCDMOKpfpqDzfN2BwF
+gPj/gkuME3dye80PwhOB0oPyPoNi9Pym5DQi88M1aG8GyPikapRGcuA+SM/
fXlMWVmN+N8gjYfrmMHwggvkxvPHAyFLkr8x03/9ZTzwXxVGFP3AZDkl1Mqj
1kbWieZc6FapQdzFqPqIFbea+NzCTMw9DYdzZzL9fZCxEO9eCQiM4nE7rgZg
q9No5sU0Dwh7DLJRJ7Pjf5myCO82CSJOTxqXw786owzJg/ct52K43zoFTiyc
fpeDUQlxnsAJ74Dr6W2cwq9jA073/JVPKZCFPAJOCR++CWxm/9yvlDRU6CJR
eM5oYUat911WXAIwDjTP9M72Z+aOQEPWXXjpBBgGJe3JFpYP9XCaiorgvjtb
DnbtlXL2OXN/ToYUMLBfmQeXOHBDOSm6gJtV6butFyfUWFqkLW+p6dGJBhXp
cddUrgzF7Qjbhm9XRH2lbr2AU/b/iB7cNWJotIbP9OuCtuXXM2Dq/IN+BFwc
DTj3pJyMski1CdR5XNm8Zs4Ave5jSx2Zns0WDIWGqLxsivxgx2mbW5qz3/kS
/mr/qurKvaWq7YHtI4wXfu88ZGyA219kSEv4YPBsaZsbYiE/e2HgmkQgWyxb
oQ7eA//kE9UqOp/SvxVPAsDxyp7Q5UOy82RtcyJu0tklkJCLmMVC3UeVIrPq
FUbiehFip+yA9drLzeNdXrRv9K+LV3+TyA17OR2/jvQHB4UyqI4TgCghg69X
k8x6m/8GD6dwAnDNYyTmmtQPA2rH0NCQXV7dHcHWM2w0AeNvXJQ4tbYgKWJt
GRKW/vIYdQb8JYchWHx2QD6MJ263gu3BI2rQVRjN2Yps4XgEmBJnZBqxc2EO
bV2fGdoc56S3fJDcj9oWMsdQQ3yqnWnVBVNc6B8IJJSD0m/U1XNKPgQiJ2PD
UlWHYWGJgN3d1M2hDeBZkF5zDQHcKoVMLty3wzry9EeFB7xIs3rR7GYy24tq
8fvKpunNa3u9gopXKheA0iS/o8r68Vqg0x0zfX6JjB0e2TE6c+XG4KuYMlth
/qO9r5ziXa+S2za/+GxYtEwnftaOfTo/DoeDa611l8xzXimBz4Us7y+g19Sv
xmULO0btCz0wKolzqHDBUDoSl4DVSeILIvQU9ZymYVNcK4y6hiMqksN2CcF+
5cLcYAJIV2JWEIfzmjEVTAJ+HpnnEYP2qBXkPLyCZ1Yjh/ygXrbu3tJaLczr
+IqFV6Mh+GQIA4kRyDq+565qdBGYdMHyqhQi+1iSGfCuRr3xCmh4BjOFLefR
goFm+BaBwyxWeE6Y1RJwjXwyOh3oe0zXiPqDM25pc4IRarwnzuFg3IhlLqrT
yhLAD27cAuuKbNzuXJxPtbALibarDbMKJhaWuDs+w4ikVfJw9htYbGgvgbYM
8NINuISDbiDbwbHIvossIlcUa65u0DXb//ohkRSun6jsuFB+xppW/sWjCnTD
1JbF9sg+oltqpdzlRA3XLjKzWioxLa6VvGYDzISG4V4KwnM/pJxfmNujmyBz
fCakIYODIElketbBRQAraBkCRB783FVsbKSkxFOjPzYhMxfoqGu1lisvmxNb
OrKCdmBEXRxyHORXKEcg1mv/M8o0wWGEeINT4NNnNfLQRIv8Z5D6VYl+EBgI
/lgyvBe4C5BfMu9P8gCACXXf3F5OSOVLLezW+waAYvz+LoDjfpiTxD36rhOX
A5whluF84u+Ip4dkMCw6bZjr+h8b3TzoBNVIxZZEPQV0mKLbqosd4wYX/sAV
6luCLZZT7yCVO0v5Um+Luhh6hubUkxHVLJsy5GQX2c9gSjcUGbGSLXktYO2d
7cJaqiUrP4baMYM3blCRKeFG9Pe65Ykh+AlMyZj0d7KSTwnQQmjew4SAQ7PO
W5v8lVwubwR9ux2LilpDDOROxzmd2xntXqX7L6dz+uSpgSa02tVzBQ/Tlhxm
xkuzPvOoEAsWhtVLFgfD5MG47aKsBClRnWcqizyT7V/DJJcJIclWCo4UG4oB
eQn//d+2aUbfC9aYge4emA/+7elUr6rhqERqmmyithb7QLQgr7n9n//aj0Rz
z04n65a41v5muc+XFCYVR1nXdNdsFBA4dB+DkY0LYsuwzxa0QmpCKyy6DGeE
WFaAnmVoeZDMGP/9kILEX6ydZsMp+0zDBWqgSiQlO4jiu7kcdwVisOnLPGzJ
bLLfiqGKkIkXK6SU01pqeaNQ1Lz0OETuGxHWthwc+FCiNWGsij5jRPCdNgvr
fYciL3aWDHH5jM1iJ2aPQcItZ8+H3XImweLe/TqK1Nz/nXBczuYp+Y5CsMWm
Jb6FrTWItBQw38SQkcigcxjNOnNNNk6Ebg+E4Z41fc5wOdkzgyUqBmQcB/t8
VSRPr8QzC/iH6iduRv8/bp8/e0NDnBmUwIyGb3ngu2p3c8uYRGqEgrDsX3Rg
zgStBncqx1RcZ7LTRF26vJgDZ/Vq5G5LUoYxu4AOEFCXH2V7ZszMra6cAMVO
8fhvjcuEYtr9sdSjKda6uhnDTbxF767jt2aJefIh52ZQ01jDTomsi0jub4KK
mYrB0jBHNcFXri+3l9aTejYMT3R9RowDf2e1mAC9w34M+1YZA2NsDaVFUMui
SGvuYsTyWdZwljTj/0tLXYMJQIdlFMseS92YNsRAcfOwBFlM/NiYyBKV5vbu
puKpQnQZJtAoJWz4Yvq5JQM4x1AtAiMqL1BT0eSrrDC3/53D56F1xrtnzqoY
Ft8Q8gel/5zZ/KVAtFSgqrM6bcck1c/vXnZZ7zl5HrtQgAxQea+OWmE3jtqW
NF1vzQ/p8XQPYNySPZdtFYDyGJmlStxkTgviAmG1U+LKxH3FZ/Kxqfo4Izgl
PFgS2S7kFG3cXoD1g/+1Rc0npevfnJpj2MvdUyY163ggcogiqqDJ19vL22Wx
SNeDCM02P44RrsttKBMCYjuY3BAhf2GPpZwYHvJ6wvjdjC7Yjencf5Hyy0Ga
zD3a8BrcEJf4kuzr1P/p9Tdgsps7vQ4avSVbXpoC9v/QRVnPs+JzTyWtGLUh
xmsh2OcD/Q0IweIZhzxOAagOrzSbXgxVqLecLjFIc3sA2DV40I6Dv2VqCdeh
3AXgeeWjQjvZQDQmGF0/JM7NxbTvmmuzBczyIpe8R9GRxrCk2EM3JyHhMziJ
mQJz4NK1kquWrhvGhCYMaawzfus6JuVBhn6TRNYE6/5LcSqQYzLxMUuecQ4E
hTjhVXvPV2Man+6vZsnBKvUwjNeW1rz77k977soajpjk4oLHClcA5EdSQh2l
fHVngPKaqyxqCUfKtbAXN5IFjj4S5gr5M1VtP5PTDV9mgQPUD+XKh/5qeabA
m1kVlbxdo1oNLEOM4Yybm5QY5vkC4cXPFXwIPDCCly+jvyWc6UVzn+jLvHg4
BdNEkU0Naeo6DxVQ96L8B4P7ntObE5BO3wkOlLRwsdfG8BrJf0cT6TA6DutJ
WAsjhdPMZi+9LVeX8v2O07YXas2O/DxUu2VC6gSxjHldHWPeiFRdEApzfFuZ
Xj+6piZMEEEgXV6VHf6dy/HOqNudMXo5l5q9cvkpUveImOlKXQ/RyV2gnXs1
tahtgwLvbNcxU/pOtydRG5nPmOQ7WO2qw7baDdc9waN7QDFq6fGa2wgx/vvS
EGj/g4yvA+icwXK5tZalHmCmWVUMyJEHhik4FnjhIWTc0eufDNK49Y616SxV
7TMdHSsIdtjAMFE+vps4+S2DzxTRONM9GmoUzDiZ6q3RNNu0FZmHEX9PzopM
Mfx6lnpOWTY/oIzUC4AQInTPobntr+DsRfF8nsSco2JOQ7yx7HxO5hw47ekJ
ixw0Y6oXn08THU5joD9WOiXbguwOsDAAdmq8hFNawtKPgGqBRDRauA1dBUV+
l8ND38zo0pQNr+a+YkSkCM2KDwPfdSIBbmdzPEUnr6Nb+agAZH9heKOTkrL8
LEyp9YveEfecBhyIWf2xeugQoEtAEGwu8l2ndYQvlcETEpzsX8p518cqdOoC
HrTqcNC1v5QtNtMsRMLoAAkca1Ng33Z23q6RIgRTqBUgWXX5PfH/1jdLflaA
oH0RbN5IJQrBwQUKsuKddsmRjY1/7ig6S5fIJ16pBSeKVjuitnmOKUkx+4J1
R1ruLNUNUuzIxPxezDRpag23YiF/kCZV8SAkeO8WJ8obpW0amZjR6M/taM1L
syYk/dr6cbR7JqqYfMUwT0lM8y109DDWWne5lt/cJTaXWa3HcfFOcLs5FNtZ
BJEkNHqkPQ3Dpse9AAUZsFNTN19szwlrH93Eb3UPCqsmJzeym7/u9wmZ4ntA
rmfifAJ8eCV4wJu4+xCicdKAMCvqYP9Nh7c8u93uRdSKVOhKMv7GzXDjyoe3
saYKy+k5jSbjSzFfQYGAmc7Zglg4kZECgTAhRQuUeL8bTtv06ZmtcpymY0mz
HjrSlw2+hat2D9YXnSyv+IjW3umvD3VU8FUZbf8mhJWli54tGTgxi9lOpibU
tc/aJwhIIUz43D2uFoqOu42A5Skb076jyBF86BNNJJkAJQGoQLbstKKJVXYr
gHJ3sSQqJ0uXw+X0QdTW05bb85Ll9gchNAoYx5c4lBFSC0nQsBkYXEWoAzku
kX/Nwvs8byw47QJOyYpr3Olu3kvWWw8D8pc+TO0hyam1oXF55+EDD2t45rBq
HfvfnxyV16t0km/OZCi2jl4SCbt8Vc+ZGF0+NMWPRkM03rFsfz7v8ywJRQ9G
RZgGmotUc8e7FPfi52T0Rd8vuveNjKz5FIJ4D8Le7KsHvpUsul8nwmwnrROi
foBB5OQh8M9lqcKOZuQOYWO9sVYMR9kGDe8eMGmeUC0JOY9u/tJZ+vU5ecX5
1fcKcD0VkNiv0TEAFH8zGMa9mjwpR52a8P5ycCwbthrrcnJkWlUqiGr1Mabt
aqTl1G2BFcbJK8Kd9AL/P8P0dchRC/4s36BO0cji/Q8T/i5NdoaSYKjDUoCq
1PSA+cULWN3o+8GAHVbEd/4P14mDGSUHm9GxCxxCDho1+wqBttj5ILHGvmp+
uADD31gTAREyseGDwCk8qWYkF9mO777rffZwyf81aFczIWo0JkHWMYc950AC
uVoTYnUXwf+a1oGZZNXT14ZJ64jQ0AG0p/aCknMETY8mmKWH6/8HPlTU0HGw
Ijd1Ez3r11jldenpBfIYrBB3eHLBKYlb30UPuYxRpQEvqeieacZOVdv+F66r
G52X8Cm0c8wUNideWdx1SwyFIxh6EDEs3vizGRs1lUwzHBli0OBVNce+pGnf
BwASIcv4LNGNybKa2qT6fX4dKYR2Wbw1wngCYkVrQ49UySN2P3PfYazapOUM
hL5prd0MSRUYZmdGfgwzcRizuRj8XwyqCFIX1vSswA9pTHyyG6m/Nhyjmhj/
rBW5pm1u20nPfqtiBhmKN3asY+yTLs+Pjtd41nLGSrMWXVye0KhUIV34328e
sU4qmECb8ekVr36rRcceNau5ZAehWWI6lbX5CUsF7Zu7UqvvA5YHPVUfP0yN
7Zm8I9Cu/FnvWIwyXGGm2OFxtZBnqNrzNPLwIEOcP02EbOoSnjo/j+6+2F0j
4e5VcI0NFYEcVrRCUl66HixmpBwDmBHqsrq1RhSAcN7S8klF/j9S5dIKebp7
4eRjNfrswlwSx1C10cFERRoybJzhAWomG4Jjg9RMZXw4K2sj+P03wXusltBP
rlTypnC5BTzTM/Ynw0fFBEIxGc8QkWqWhnKRSZEHaj9civBFGkXIjVCWyRf6
uynKl16qUcr8QLporWzf2oP+UtTIQMfI2U/gwRnuu+niE9IFuR8S3WrWn9xf
nj0tHeOvW0XM7FLINsR6GN2593ZHgADj8bvFNyz9GX1UJWDa9KBtl3jIaEyA
31lw39bqAvRRZIAIApfFbcovC+eBS1BVlhQTVew6T7vVqg+5YeUZ/5WKrUtb
T2GQ+lFcJBChmUNC/T0DB15cS4mXMKSvVpxgtBLb1/ba/dpOysxoHMs+byTw
y6fv+UjrpKb5+/qkkQDiRZ0RDgkF7p+B9dx0ebMo46jOjOxE7Mc8vPDeIcLC
G0dIfTijaoTsW5S8djwxDoy/4FtEaTOqxjvzlJkO3kCarQutIQhbFpFcVeZ6
x1Vw+xj8CsNVGtbdH+YsExOZVs5BIA1spR8XPmDSP3d+SxDW1RKV59wpYEFb
ws2sQOBA6PYYL1ACCQabWd1I6pCZYQCTAe//N2U6Qad16rCzvTBwphnmg/z+
rKJlXIMS+fvjJtEGQzJgAvojbkHNmrsrQ9VDO7h4qY1QCimbkxxrfieNT7ab
rQH13pdPjg1sMMjh2iVxEfzfu0JV1RXkWdnpI0c2fJf8TMhgXnaHKLvXwrzB
dAMynkanoaYRqsd4cznNdhPugNaoVyetVXiBRd1/rSoX+lBqnzUpYhBAxKFV
rNsVwikd3xNbmssmTlx1PDa+0uRZ4Ny+6A1ef4dxDwNYO7U7qEGSc1gLZLLv
i4OBAr76EnN3LQpOIUQd7dhAowIUFZtTd1bp6Ojb3UuDOLjKQisIuKRSaBac
JkhzMCjuC6AgNiIF0e9XITT56MkZR6I2KGIAQ6x4/0btaUzfZAPrW2WGyOML
NHfUJNL4O35G/59KZVztwSUufb4bO+6QcBDP9izuHrfCYauYzop/1M5hR1b5
3RUBJTMWsnxb7xq5dJ8foSUUC+F+bZ7MtykTVvkndSBvtcUKG5RhGSz4Sufc
B7Erv95CSOOYqRwThKcguaw3dqJVcuHVcnW/NXITWI2JAC2f9gJzchYxHaOZ
HwL1B8nVTswm4WOLRHeVdfMuZ0+Mkh7d8Cl+aA6IJCNpZm+ymqTj4qJSpLnL
rZekczV1oGpAWxA/Z1+KV8pcvnPwSzjadIezhMsA9hY3tH8REMA9Qjzv104C
rm+Vle6TglCFHB5PJhKaJpXPBnj8f3n82pC7fCxWr2OFQyrsWu1T65MluKuU
DRvmenIllfkZrbT3f6wjZJkjYSQT8XnxdX3kFx0rkcfEMMatf9/Ww2+fYV3O
H9mD0kQKtUNCc4oyc2nQ7B41Emiud6dmogRxFnwonqHLKDX2yp2ohjW6PewT
p/ySL97j9dJbUEvnp4O/REb7nEEkeVKDQvOHe30jEAYkMl4CMQckLr9yXrCM
uig9Npq1jZk6kym/m3/3SYM1MhqKKfFqqKpNth/jgGqFX+jDRL+wr952dK1p
5KCkA784tDOxl2PKWaYHMkyv1LipGhqXpMN7+uGQMl8PHbBPxwydrzJBO/CN
G+i2dNsU8Cx0S8hAuLEJXt/Iazv5rDoFwuXGogjGzgsU+H97a5rbjFfUkun1
l+LEfH+6NvzkP+kljbJgVt0PSP+q+2jkGi1yOV6c4pcoeVoUks+62mCxJLWo
9ABpTOvPrj3q+P0pFET9cRI4mrk7e3npgi+/A7qXDJgLWFT7HXsbPdtrrtOK
5UE6Xssqps6zy0APPuQWXTUoZKpPtHXMMd7QBrwtOgJDcGzqlePow4yrw1Pn
MADmodYpdpR4DpdufoXQ39Tj04aaMf2fh3k5xB80maAyCPh7cNDpvehPZWqU
zSm3/Q3TCEPR5nhECAU4tzq2cuhsC4TkWdFYoUJqdTpB164Ko54XHmVldwIG
v5tUopOsENIOzmMiwd/mXKsLT7xYH+Q8HF4fhds3gRu/2qlOS1At9PeMzqtc
WfSyH8+B3vqAirRxJ9n4URy+FhBoRrmiIV6ZF7NyZvFXy6So85H0Rp4qCuSf
BPenvoTfSX/YTh0cpO/uVRvcaLqSCj+AjmY8x8nJxugeZoIM+R2/CmiPnViC
TMJq8yRsMiJOK+SqI/H5iIGKHte4WkEco2UuOpceBKtsskjZ+9Wss/dhsw5p
MnCZ7lkCXvzKjnzXv1PC4obGaPwzECafiWBXPHypE2cR4Vp7F2V02owTX1ql
I/kTms7ney8O/WqmlRbIij3WJMsPuXULLG8/3S2fGAhZ4fKo5s79XppISelG
ukUripQEaj4mJlXFKkdG3ijO4SU/aO+8iOEspxrnX39t881NKanm4M5W+qHV
N1F1xEd01zGUOpPogP6vN9ttjdA91nGCqWhObSpQgdQBzv+d803icVXL229w
MaMGRLpJEhFBMokpmxJy5/O6zF5NzpdN7EBwsjut739omA2xaothWH2ZgZFq
4nOnKqeZKSwiXlhM1CKDUss/IdIufmIZucPK0cc+64Y+z2+YX7D3GggDL5dm
+cCPaQ+s13XwYfLUmmep68BquYn+jXg8szsHMFaYd3NCXzJJU/PYXjhx7fQP
otLxauctep5465jsbU8glLw9NJjEjGeJ1N4WuwtIxR0UNKrGC4+KgX/+IMYI
2ehq0KciYW9qyjnkueILMdJ+hPPLCaOK3A++A2AQPwfld+IdRa6b+xSssXVU
h92hXK9khLg+jOISNqtvDc80Z/by6v+63Aq9O7+WI/UIY+mMbn4Mqdpr1+rR
IFaFgrYo39eCub9RnOiZHiMhoByimFgPUyF43Ov4wiUxOZmwA+/eMVaY1m3d
64OWFgErRfTJlVDs3eoAFTDwAoSJRIlQUo4l1WvKGsOCp6AeCMEl3O+QOVdo
5Rbe+e7uCpamNw4Q/rhnMU0F0d9hllhNWH4GloOzd0v5vqFoD1BpV8wQRPom
a005idjGFx1GYfdeWIzvnk2IFww/h+Xgf9Ne503WhAjYkpmUBsP/Q/02JMNW
Na58bIUJYZjIWEoCITGp6Ph5qjHP3ki7oP3sgU0MjFIEG3coK3CgkoPxvyNV
mdimtf3KIduDvunj1MoLF6YmJqMmQeR0LcWQcevarbLTfJZaCr+lAIXwATOV
rnfDzo1sBvOHz7TFzdw7F7vR7WoPFMmyRsOEzCJN95TXrkE2XhPpnatxT4y3
GMwhVLKgs77VQ7PJgmJ98I2fcJ359/QD7Nt9an000Fluxk6VdIMnh26Ekfb6
Ja3ljxSDOmO37NwJl7hreAdsM6fNHUiRhTyN37UKuAxMrGzs8VPUJWDLYpXG
OqQWk/2pab3oOiTSo7kwXSDhXTpeYK+a5gDK2Xctx8kzz7SUrLyzGRq7tegI
kvusasCwyzpvN0Doya09Rd65OVteYZ7D6V5vOm9A/ykDTuwk2Ue6oyBLVJa4
w8h3uH9D3dJVPn1bRuVaE3yB0qnZdAdNKMGOPyLf7kVW4m+QKK28PSfpSdU+
wcyiSjQRSzTBl7Yirqrcc8E4bS13l2fNzvX473/3F4G60j7zsCrJZlY/tWf5
Ad1kyyW7AFBk7geMX9e8LX60VU3TxhXYsnuowngU+PtkNsLCo2zFJ3oN6fXl
xXt1zHHOMg4IFYIS9pYlo43/dIWqEvhNLpyIG+y0/xCpbd12s+4xOzAYhz+C
RGy+9w6b9t5CFw7xIbNw+VGsAGVMD1RKlI78uMlKfaVxgFaQD5WRkPBlxwt4
pRu1+TQSuQlJcp8ctcbnRmAbrYwZLEafmZ0JfMB40A0xa5LE83IJmHXlidwZ
T93Gybs/bgK835vDyiTHPnvwxDRF1R7mnf9j9HW03u5YdbHcNl7KOHZZS0u7
8ABzay5PMJKrXHcKNgnd5VpQ5IY9LdHpRtetn3Jpph0K6iR3qtSZabFGYGW3
ggEb10qakBvqI75NoTjyyb//7pttNREKGS64Z2Z07TBSYBCbmxVlFM/dUIfR
hN+Gb4DRw659D/4Gs+gS4Q0ElggaAnlZKJXcidAczvXMmIr7alz7yCHpqYNT
8uGpN6Tx3ehysigRRSumJMhT3su0fIVWoziY8VpRkP0/2kokCZgbqWKRuzti
StnaIhddctbtJF/ZKsBCBf+YU4T9HOqcha8iiXuoxb5aq6skhVRf9GQ+2Ozh
+kO0LaNmmSO/xs5LCBY39HYslW2yzHrGWuxwMTqQuHlm5Dkm/NUHnX0AM3ZL
uC8xaDJs7EWG0YfOGzkOjtbNnHI+c2ulxlV4vM5JHtceaMFTSrqIXsFcLVjl
oCHi5IIHs2cZaTinsQ6vL4xUd3U3Fw1sYo2sjB+HUdYioYMtcxHd1cHpc2v5
ilN5c+GHqJNtEU8/3NhkZ16dNPO4EB2ovUJA4N1z0b6fh3hkl8whRTMEZLba
GrISktHev6cbga2vTgAplItd+6CRv4G0BvqDDR7UY2/+TuV4WphfbypCUmM5
DVr46KwPvSDQSZy7tZjk1VEJkOYT4i6KbrYcJu6MR2HF1X01oqBh4yJXPZcS
nyGCgsbRrYyXQfwMg2PiBB0ocwIczBT7sh0OORgIu8Wi8xvPwuFrba2z+Ybz
Ln03ZkI2oZFc8+3OBlaf+UzMASAn7j2RSk2uPMKiSTzYCgNk4Km0TekoTn83
N1tZ7FmEUEWSYk3F/HW+GjjrUIMO9qHX/6p28PsI5L8OFWdRfsyWDdCMJ07f
6Rl7LPo0I1iNIz/OSpyAOrVgoFtDAVCcnfZl7edgkdd5Qk+UmVESFrftWQz8
JAqI+zNFX1p6veAAOtEPEI/H1gbF2kGxRlbXrSMuCyj11IFGw3/B2EEB3XjJ
Ku53VDjDhtEPaY4rqBObKh7baNwxuc5WHwWXmpe2cw2lnU8V7NysJWhNhG7X
BUB3ZjCX9IJeOrUxYOjzjW59zZyt/jXAdafxNXanyHSBtA9HxgauH/CMigRh
tapXxdm28pJt9wYzgEfhISWXSGHT8O6MndYpO2RPjZi+dwgO+NxqBc1MER2o
+wBf3ccDxYkSCzfNMb4LRzZxl+I54X7+VXlb/ARFZ1NfvozehbXVTKjMpulQ
R/uRPcsB5N8AwAEtWrh4BCghOqgD5uoaiNq4BaIlKp0SNmeJFDuWaIh2OYPF
w+U7X8aode8p+rXBPElbLvGP+fp9nX66lA9zc5UW7OKHirY/RLmzdK1vfDf+
S5OjxnnLs4e2iZ1agQiOcwSMXsub0cVh9x9BA4v2FsQWra+hP3Q4MOpj9XG9
6bK8wuLXO8Enaf+rUA05V0B52pybL3Ok4i0i15KBNnUQfLWH9SW7iswPuqNl
gareja4uPChndGyqJ1b29Xq8TbF84MthwgEk6go/Edwn49Zl9rDqazbW3mVr
2IDfaE93+ztLX3nJMqkZcdy7VFNbmMPK3zLrboPU6H7s7r/EN2PqQpoam9+i
jTmywnx65nlNUVhiSgqPto++AQUJNqjOLwySI+UtYHXwpgpFrfTK/ekalM3F
aEqqEnBmWCJWYo6ggXJy9C0yKB/1h3FgHKgi7gSDPaW/x2dqqxYElWpwjD3O
+T05YiB2BN91tMB3uUq9XqZBKNsDHz5yjb9I6MtP8uUt0PzVt373JS0q2zpm
ChtVmsvLyDShiiRY1MPKgegulhDXdOCMvV4q79PV3vUnBhbqHliCPGaOPaeu
rtsUXyLICYyrTDR14mK+SjuHGwx4ZE9Vh4g51DR8c/sunn9Z4t1bK/Gc7jJP
f1HRDJ4PPm5kg4/0gXtBN8ZU8uCR7nL/HRtuxeol5ArbwpuQk5co7C5oSHob
lUxaIbd1ctl/GvWI/1joUJrwr0y+xivLrVqFpxcqJNEre/BqtS+Qq5UJmPiS
MGgYcHAZ0x180qOIf0k0pBb3ST6Xxzi7oQzMJg/e/giNXmIY8nC1UGbf+eSA
C3DXi/LneFoebUaPB/vLph65er11lu33m84bMW/hCxTDa/envV7pVISYzABe
JFlGnCpATIvsYnOnOhlJl57K5rTBT1Dye23u2aiyTAbfrj7r/AHAphdnwgIx
SRI+N5YfJyhhVkAC9qmROhlhCUjDM6ztmC7cgGwpYA5yVhfIz0xLv2Rl26Ja
5TdK9Ny0qMqz3bvZ/vruJVC18F6kR0W9ZnX9t6QYoHcvfPn6R9m/hD8Xv87c
ZJp+VO4ag5WSv+ehNPFYYfRWsQGZE97fyESwSWPnLN99rG2vEw3VG+ZGo7Oh
cl1vb4W9JDcmK7bgxqK9jBxH/aOw0/J7KlEXPatfFkMwffxS4REPi1AK2jK0
u23GsJ/9UmdwZCZvpkUfXxWX8MDk0ae9haRn+73Tp+DdAOv5/7YSyMtbeOlN
MObiNfpfLg/bvE/ADtW095dL3GNwffmy8TEV8+HeBoiHlUn1OHWbNDzWDsVA
U1gMFKyiGHPre3ajtNR6G2JydALEdz40F+P2OAWy5kzamItdX69Z0H5ECXkZ
rMpBZ8JAhj6ru8ErLsLwVp5yAYOVeiIPUaI/Pi4nxzVmZ0er5bPHO5OOYJL5
VEY4YugDgi+1HMMeAqbzPEB4GM4XOnicd2icbqGQbVqtNN3AIrrsaBXN5bI4
+Pr06YrqLS1q0umZaqCSzwDg0d/NvozTEEbu2pHD/Z9PNKh4Udb+O6m6q2p+
2ZsLgoczfk4YO1KLvcOL1zHI7/jC6yKcNsmLy30ybjebYUECkU4ZE4BN9DMr
+ULsBDsBN6NfrArpHFI57cE4IcYnYSx8HxUn0f4GnNGG2xYgDZ4bBpjQUxGh
QtmB33nMNWAYwxkXLZji+8neEAtevByCpvevDh/HDj9eG34GRYF5+gnpZCeh
kp88WeC1TU+1AMQH4X89zJ2ClLHASB8muK2dDj2ItxPDZXmfaYU4F4fLUyHL
UfKpszk679W42Ipj77krQTf9O6Mn1X+gfbu4qzc87eSysg4IJMAp33m1iTjT
reFDMytKmM5uDsjij/8Q+xaHL2em6mV2U4UQKXDkRU61jmj91NoZ+R66QHRM
M+GWWh9VcCPzRc6DXISx1VPDPyBtJ8dO68fNKMClgDuKWEn1Ml4s739qIQI0
n8XeGRDBkp+NYEuWqX5c1ModP87XW3J9wHWkOOHw6B0hGQfQRHfgtyFu2ahg
tRaRjOuiKAVt7y0DLaq5qtv1XbxixYR6bz4J0GdWttXSBabr5gUZoGjIfcWn
lpsRt4ObhFJunH/sC/Fx+8YyUKiVWmTcwv/YlqLjKEhR9K2m4GfAZnxm+4CV
jN+BXICWVYjOSp5qTCQ5yG6ERnYyGHBklHOYs/ZnLYAMheeLOqrw2AUsQh1e
HAc41SQbYdtRcSh9Bh622onfBtnSdm9+w2ZnTaiFI+4OzC65Q7zO9dtkRjAK
RXUExZokzHklTWsvk+i0tc3Ob3wSy1uwVTNzKNMqL72AutCVwoQPUqB/oqfc
0jepbgl1TqatOznmxat7OTYeSEpci1VZGxOCNKHvhbGqvP53Q6RNxq08NFPm
03IjSFkFvh8wuZ6OnXpTD3lfGT6FMpPDyGGK70fPAqbkZeKIfVKM8qO1knPz
5jUs6oBSSsrUrotvNwwxo+03H0sSYvoYrNm7JrOnYnlER+UnF/H7MGs6OIjC
bh5JoTPqOynnkkyFEUpo0uDguQ4ReMtr26Xyk4wCUl1YE+WjL2ugoZBp5cgL
z4yEHfj11L4+3Ruo/CMi8L5ITZBIdLor4r/fpiPM263bLJ7CSWLcbeLao+cc
e+s8PQogxIFvdURNUSysOx/DO3pzIFRrAZR4Hfyr5oTsMi1RFaz+s5qgWC/x
7pbDo/CPCCIEhk0I54Ju/fV7uKql6MRnAnWQjr0eh72lUmwM4oW7ykGFYNe9
vwQlMlvc3jhNUZSFALBIAGiCFB9/bt5r7GXGlRdSwsA5xvNQSjKg4aSeh3BZ
C0RE1PBMxoR8NEw/V8DvowE23u+bQBKoxgT1+7S8XnbsldF9x0DHfLog1vSo
/toXjAQIaZ2GNHXWju0MC9MCM4lpWyk2FyU7ZUbbGOHgMjGlwYb9K+tzuApY
PiBYyBxp12HoNLps7YoZm2A0IPZwxwYEoevu0t6mN2FF2Bn/TVGCyXRJYiYq
GliNJdnDzEoOIhXtc7jH7b7hvJaZGK/aHkmsxTJSe+QatNeCQt5rBbkOyFD0
13K5jJC/SyOJXzL13G3J9HxNHTFmt8CIDp57BQ5RGcGPMzEQom7p3oxk9wt+
W9UgVRT6Yji7t8LzVcFgIKsHRD+InImwqXXc6v6543RSrBAOrZK7NKcnRZTR
i43Pe/bhk268kmoilVpJZt+yXziHNmmo6lwIRPgnZONW8sAuIzvoqfgrPnYQ
KpHCixskSsNp9sF2maqTDwFlp7t76V8oNhRDWpoozMsfus9emyWanq0drXKC
vj+4j7jgVbmoQfkkZ6uBlPaImmKDHNmXNGvxtr25Gc4dEb5kxQD98Zc55qsx
kFr4Scu5NxtjnCfPGjihvYQUwtOY+sPQhaQPN88zpolx7B4FcuPMAcvY9SPZ
S43vxXjlBY6iABvQkdF449x1o3CE+PPTPYlRDtCSydfgs1xxeEmXR69aHEhs
JXT3k1tR3bVpQT3KJqC78rCsXgFfLqICI56vWW+CS7LayLvRosuVtj+B0pOx
GQODfpBQxGfzpnfpeqeQtoool6D20M7s0ZnA2QVlzi3zjzXCaZfwsTEJ/Hy8
LDgDcRBn7p/SQfhvJAPTUBPJIsV/1oS6AlupL1SKVqeuHRrlJn4as4M39Krj
P/J7SPo7jXbP+qTGAgafZKmpF/o+tkHceYHqcKiqkr5Q2vlHlbhEKH9CzOA+
eF/P8wByMAVrNzlaYY+s7YyeBYsyJ7ydj+VIMIS64prFwz4jHIStjS2OjxFJ
e3tz4Y1m3FsY1v/PAtyI2rLtlxa0iNilbecfUCO+zeSOBUecTpUws2eKwpNG
Iql3Vg/h5GPPPEzV2VQNebb1QirqQUUZq1uXXCeaz03A28vbSgLmYVPmV8M9
1F8dN+u3sPqkeX1eW1Uu8ohXg30ocbxWI+87C7NE8DX+X64x1CIRG+wMcJ63
NJPERcOcAOEaqWAwV5wVwMwhUpr2xXKYYlCvEthzSVQ0XWds+JO5aW3qUJj3
XoXP48YtUiqYi7+HcSI5ImWZwjHwJS4IH0e9sl+IBC6YAtwNUIpNA9opc3fU
Ps0wzXShh9moSTc1Lu8wHhxsKQ0+xokBZv49M+7HELC3f4lyV8vE4R62PxP3
ao2pnTBReWhcbBnB9RB6xRPOnebZ6dNFbjs+YS/e+ZauesBY6u2+gbQkULDF
+zQCL6hSD4kStpWLq+6E/mnaWxgMUWv8W3ZSufmMslKQCLzezshIo5ynE4vL
PoS94AiF1KPTvX1oY/pTuOMI4JfyccgVBhp30vlP8TGQ2MK7KmdKh/m5asEa
udXeV6nTHTZ01Z0F2K4xtUdo7LG9vRDQxkLQjRXydwuiXryf9pDg4op1z8aO
imMmIvILVj1WOckB4mfsLY7v2Ie++FBjauAVPxxh0Jro4nsq9tFpUSrwBakC
QrfaNa/98Cp3OxWCr9iM4TIq44nOFFkz22CzEq8pX2yfBx3ubviTKq7bIgbb
LsnHYsX7slT9YFEXFHEQIWLagetJmfB7YdkwsrieOXEsMB6nD5AIz/N1n17W
WEAeTcmx7A1iC68bafJsxoxbOXOxRsdak/f5ImxvDgsnpQW7bk41YNvlR2PR
PNHCuwQSmzSwYRXtSBtemto9R0b23UAAt03Tm4jsoL8IZeHBrYJzhRV08Q9I
JUNLgApQbysXsLeJjdLeFpVhuQBiUDma/rYyGCf/1AoT6k+Vfq2gSqf6hNNJ
KAfigaTkxWIcBWx/wjmgj7T8XTJ6UdVGA+07oO1hpqgLT+Fu2nXNlBzif5hy
0kE8qzQ4IXBRvEth/ysDKL/Jpg2uN3KSSRmx2fNNLDc37vT6H5t0AqMz0Q5L
c8Zktr69z1LTQLGMo4wdTrdjPjfE1HAT+payv3I1J7oIu9/k3atPOPNZ3KGR
PTN33uktmRLElh0hd5Pk65B9jKiygrCVSqhKng0Qe2QBDrhGXNUVkP2cjKPX
SrMjEgUU4RyX2kH4bhM9O4q9FHCD+4irlKkQUiHScwXKeqQ1avmAm7CzeBl4
iEeugKhYSLw3SjvHn/pDvFea7j7Gh6Y56DA8HtccwFW8bIHukK3+2+dszN2U
5rF2kq5Fq7cw/1IwKRqDR/heFHI9zEVXOhCFHEdjdLxuYwp3ZyJvQkn9322Z
CELIjIgSwmwJNFZHQHyCQ64vPUYUITBwhaDqU5tnhhfIe4s/RJJyKvvdTHpR
ghbWGjMXSRHfMMjnIz+8ZQzYJ4N2hCutpmd0QikOaUl0b61q9hf5yp1jydnE
RVV9KKD7aaCruCEEhhGrED4Rmv31n1WGQKqTqybdtKD2RhGGZLHi1i3dlTWC
mSb8P53O7hTAq49XEzxAM2X2jU28p65ky9wPZFTLEYdT6RLwkSzcHg3empr4
4b2gkTucP/qCPk/pgRI0UYMOZsJVvtCYAhpZ4OXELBcaH6kdtR+4+1S4fBE8
ykjXQalpH/vZkrAVBBNg3lP19UX7ahGTpMjHIpWj5QG3vaXIS46+BxSh0CV6
8wHEQqyAxL4tfldM08DwbVLu+NET/h437+cdCGTdmBAL5D2zQknDnyTtIP3a
iz8bT48WUNE1kZfKScGj0TmWRJ780YbqBj6ChaXD30qZ/5bOjyqgbXEFzR+O
dFXkyPoXNsohEgJeUYZeeZmGvWwssnMeCHOIVkotrIlvRb7uRXcOgM20q/OA
obWIfeiSX7lhHEqKJKdYZzExmiRD9+O4tJgh8BgU3ARX5EXrLFQnhiyVmF+h
GJ+9n3f8gEXAwg1tBP5xj3lwD4WQjYWDik5NpCEMCLqiUAnWrAdYLFhEFU8d
uvFc6CZ0upVlHwGxJwFEqgYri+lrJhvOqeM4oKdeGg6ynKvCEcf8CoD/lvj3
0PxzdFOjNjCVeKiCCqr8dfaElWfI/VhFinfNXvwGS/aazR6bh7S7u+65H5Xd
FtUEo+p2rlwRxVBdyrimtysWS59d29trf7E5yhhLtW2y7JBr7AOdt+BkUctw
Ysr1ESULeopINozcS75KSicLezblUPL8qvWLf0jmbCsXE/jD+1NM85SXY8NY
B5nVd04JdRi55zgU07pxEfpYVsuF2ixe+fVOIE0+eJnJAgf4lCS70aVQiAxB
f/+Tdw0Y+r9l0D7fHzDWECTSsiCx8KCw0IJkFcxf0285G3AcS31uLbU4mwum
SHVqIjAlmU1Hisq2sLLjoPh9iiRD8/yMxjXXql2PLPgUgTd8o9L0Khb1fCvy
lOUSfe0vVlCS576z9+Y2X5tLsupBMW4NcMY0JmDEHm3NsNnQN6/NW2yjRCeG
Peses5t7rYFAS7u/BXnwLsL8Ec8TLzTLqCsl2mche7MrIabcJt8i0IzmFSnm
a5qZNiC2hHDr8v80nowFXOKtcchiO8rmAWs+N951Qy1nOcwop0pJkLaHYLBq
IsC9A6L8yIo6BdElzbYWPhA6tLY2ab8BIN4Gop0jWc5f1pDhWz4A2l+QQpR+
KFnB82CwgPGTO8WXFGXmqqUcHmeSZU2PEY8ECWzoj+s//TcBYAXtB3L9b0jW
u8q/xp88uyhR96YV6xKRpqyHAOIofsiV6OOLgIC1RKeqT4b5Ja8JOzNz46aI
bp2ZJVfgSyQpqoAjJa84HpTiHc9JlIO3f59Jc3l+VRaQp7X+0KEuk5F7IjkV
Nlv9cqvduEWXQ4KxOGCQay6IxhFK1S3H7LVXBfvpo4e3xsdZCuZZz58bGQ45
/wSezhtIpu+Se+jT07T2AmcAdvTiQNe2SoRG035M3bwjYPCD1WYagQIOR6/2
8owU21+J9HYuM/WZ2DYAVQQ+eME5ehxYbg6ZnqCy9aFKWfKOFNJolayFQ83m
uKIz+25aHhE09GUvi94X78niUOup2GixHZzvnaTOAu25iKtv1oq8g1g4Co8k
W17uXh/A0eTY95vk20AD0Oq6ca0BR/2aQK+xIY0IE0KLq/xpdfWywpqlNZEd
NB0QAyAbfFb4mQvX+oJGBOqQ4FfGgsQ1wA6GeTtKAQPKx3i9KVruRdQTTZJI
zQvTl5Cr9f1PiiKwHuIit+aFvffkS2ASGfxojvsusmsWR17hnOAg5AljGu2W
p4Ux/i4df3m6AM/FXgWPFtluX+Jm8LG9F1Gasapg5U1EXpKEA1nBm0GMR9sc
bJZyG4Sj05ql4/qFFw5ImPODLAAZAUfPaPU57Sw0I04HS02tdatRTYD/um8h
qpCmIZp9LTa0IdMGlNu/rGKkwDTYD0UkG5utKTi0gtzDs3K9DmQDa5LQV93O
9vjTNkwncWKSOl/N1fF/c3l3RoP6DHC/FbGXBt2+ZsCZyT/NS+lcDIA5NDa4
AzJZIUk8rjaDlr6HmrdPIdxspYOP0HMXr/NMzbWl/rcIC3VplBE/L2b3d1k8
v/SZzMku7O/+kiKRKFCx5NG/xwpSMgmkHxVPWZ/hRW55wci+rRt/TPrMvJ+c
4Xc5m/G46YZWTE9gHLouZ/sCVfQ+qf+iUmcSfrjB+lZxAh4b3bAy+wKWaoMy
KK5R8264wtMVGo88WaOlN1wBD2D5qqHq1m0v9I2bi2rwCCJbepk6P5WYwkWs
8MMKlGDfTbDsuAzwZ4rYModnyvQgCQVHlgjaGMVAvMEVbzLlPcsGMUhoKHP7
vC0fMP9RlrXXHACUV/7Q0JKC608m56QCm9wtwhe5zCJS7GGbC2ncI+xxtwbI
jaFw1oe4R1nkME+96X+Hq+iQSGVZF97nllbAIzTOwd4/nCzSBZUrxD0gzSYx
L4DXey7A+lqF6NSTU14sCw/+WeiFkcOsdA7bwZnuYnlfQhLpvxzP1c3N+E9u
wexY5Cotmq98zx90MAX6yeZVr1Ucm8FPombgUD8UBreLAOSTqaHV5MZTC5b8
Mi5u9P0QBm63ScyK9e4CiejrhxaK4d5i/AxJ7nRX6jx1xjODobw7XC1jFomR
DweCZBwQHRYVPLCOKP+0Xf6EYolwLzJ6xs5bgTyAODCHL3RUFskQtOYuW8bU
koerAwvBoFx28QqypoY8WQhFk2wiy4fC7V+jPi93ToCChm5mPZ8vYY/paRwZ
32/6vQEMTTLRrowTliz/6GH5KeWSDZIp5VKC0aSi2jnW1J/aHvzeS/R277d0
rqICUDfHLPOpXDadkcNmn01EDfDFFXoILSs8FZURL12ljdWAI21YSTyXtT6Q
AWt19H/BIHxZHK1AzF1yL3sPamuoaxdB+D0RSodaOL63NTB4TbTc8PKUBBi0
p6zhVRxIwDN+PK/hCETb+5jXWOWO14qUpCzcz/UQrWDAKpW40+ySsFgGJXvF
8AI1SH7ItZqSry27jr/KD0YYGjpGWVMnq+FdDsIr6pxovovK3tL2yVo1DYkM
ffbX54tbR2cu1xngszuPnQeO6sxxiKdDZBsdieVfntPO1c1i44aqDrfNZLqI
hxZILtQ4trLK4I1KPgs1c2Ng8EowvrTugYWtRVZArui7UTa3scvI/jEEwevy
htVIfGuWLJLgD7BqCVmB13Ar1HhTiY2NBDBmRwbOpw7jGkYr7PHtGqLeDY3C
YipkU7KpJgfnRF793fSqgH3EMpE2CYW9lPVZeccodQ2URgjptaYWFZM6fJFJ
IJhuzU1I81k8+RLwShmjoxNsBLOb24qDs2JARo6EPf8V3a5aLNvtAM1TQNeE
irN8naR0mjEVq/hE3kIgz21AedBxODnwW1jT2nnFDNUeZLjfCkI596T7O8us
2Mjv3piQCyQEv7yB4KGdDffQfYXC93cdOQd4pwhc4fsNZSrGglwQFXZQga2i
dZNu/Go17goFp7LsHTFpuj8iNKKjMX4ImitT0FdlQ45a7P2dRv8x2x/AMQX7
PUessJUOkrtmdWFE30bapvA9sOkI2mee5Y3/lPe/mbDSBADc7MJWfxSV9qJY
n8VEX4xHWkYlGNs1YZUP0rOo3LqHN4u+Issau4Sl/QEtkOoO0Zyqm7wKmE3U
80HcTCeerc8SFr7TQS/xdOeqY0wGYPLj1d+opI05BOBawjUk/D0VN1uEM7yh
M9lKphhK1dGkArmm/dt3PHweNGg7wHAqSvRIWMqnDwCsU6yKvWuLJkZDVLNM
kSrr1ANIJxH1CK8+GJbORl+K1ejS/pNaDZ9z3CItXJE13XF/CiUqsekrUqV8
EqoKyzGyD944QKAa3ObUeViQAJw7EZcXpPBkIc5xEp941Q3GLUAOUGzYZ82T
J0GkvZ/GHWVwYXjzIoiiTNZYx1zHAXxK6ngv+OyUtEQZMDdyFC/ZCijpBc+q
0EXdKN4XCoW0AbPm9C6i75ftgSxU6fD+q7Mp4utPlR0u6YGXY/ay+OkSKFdK
sBDbaE/0mj4qsNTzyp53/tw7ST9s/0Jbbh8W6HD3T7eZ6ZohL/tnZ82638ab
GMCpBZOGf19ha0gzX5YT8/GVgms/A2e6aVkOR1kCYew3HeHct0c8vcvpHZr2
sLo08jHBW5F317BL5AsnUOhdSDiDTjrbV/fw42rDa3G5Nas58CQB/yojXcjI
tdfTWTsOBTGgkUZHXjLsRyaRW+ZyseJmVVx/Zis24RdE2eKvJ7/GJk4wCNPK
jmrQotdxBXdEJ0PB/+KMe7qIefPEiur8oW7w/m6Cww8agxyo7djFGuBZRAwp
nA0MxKFQ7A6cf4wb5YnrlKS9+sp7rzXgnpSVuex57bsRtfxSd+4+Hc4/llGI
fA7I5HUJrvN8cBROu3LOMWDpX7C97S0pzY0WgnsO8KGbDYKORhIY39qjiCba
s5TeK0Ub2Lkf4G1THaiFA0CHE63LdEL8Vr73Y3ZQe9ugzMnfTSwF4bLqB9mp
ggcLDSJ8ynpLUjSa2fetJXOSBVQjr4V6dF7qhxL6IjWfRFlucByupRAeHMXY
qOH3NxJcJy9zwSoGfozITZIYNODeNJG9ndYy6b0BIrT2myoZQ+LCxjM3Z8St
aMMlvpVB2awdRT246o9JwbLN+dn4gTYcja62btG7Tv6rrIQsw0HKwPwuio//
+GNtcbLIrCScsBqvX5EgeEi3f0OR3VwNWy9A8eoagH2Z9+FiBW3F7697hTDS
HtpSPQyvOnKLU/RyddGXrBtILbPQI4itmrQZ+C9tRYIah6Am/M3pVWLZRVIl
5pfhLDoSipPiZ2J4mjp2N+CaVAMQ/iOSzZaUgA1iQmE/OXz9Kc1vnm+9nvXh
ninDZFLyTSF3UOUYa21l/juWhsIHiJX5l4wBgZHPn1MUch4woiYw90YO5jQS
uGRb8CmNkv3F2OWzmbPN+MYTc8cT1HDJ5Ztkr1UKwpnCnFH2DIS8krJy51Yw
t8H7Cq+tjx7OsDMHkAo7W3CpguSpfrY27djAs14wuSVZQwVEzdkGHGKN6KGv
PhhgOF79oQ/oVAdEKwLeyOHrjHb5ATo3avaaCxWAVcfX73ZQH5CFxMlGgkya
q8XI96rrjnCOuUhtHNT2UcUYvfE7IPmTgIRZx23j9BE8A17ToktLzjZefZaE
+4CveIYBqQXZYKnPZ/velH3NU2qXpVBJMj3aCLHHsYT5nfREiqZjFjbmfJAS
vmvy4x9hWHyoyqqfHj4fESzUm3yZXYwrIY2CV9LkH82iv8mBIyUjBAhNSjMw
hTRN1wLd+AvIs3mqCDbXCsw9Iy3CJ7gMI+s3FvURofS84oiPydt6CeXJl95u
X0RsKwBvE6CGiB6DLFECdblGUVfOk6SakLOrWybMuoT5TP9pwtEvyscipZ0A
8id3GqR5IA4ZZ6WB3jfAkohoHDjHbBlLKuoVXeIPDQ4s2tyytiwZ+eCzDfba
Y53Q1bpa70rqUnswGsC/m9rKhw3Xei26jDl6HjLH8W+V2TZy4l0SeXEEvBzY
4pvz3KXi+kIxKWgVjOgOMMCPQTyT7dPuiGsn9knDMqISlbjwRHrM+TLoS7yS
qS3miM8Y13g4Pq/ZFkxjMzdjM0sJeGElddkrdmxOFVAsEBQNz7r39nBQY+IF
PmHmxqVbNVKWFmRTHmGAjeIYDLonlDMzLmMZPfn3Q8DLhQ9Ub0+rCfS5skfv
Sjdv5TuG9pp8wpuseQdoiq2pQv1KcxMxzYg7K3H0vVewGN34vxe+tCLWAbu/
ABSeGyBirJD/uqkOcYMa+0IxAX+7VN8MP01UENout6aKE2c5R+vWboUxgO0T
bdz3Evynd7uSpQWezPvvfxiFUHRmKp2ZGhBfj/2ZX8CN5jDA4tAUQEnySW36
6hCO+1cxVXMRAmUuGAFbcraog4sutqORUsUjCo3muG3trpf31f0GmCKwMoXi
DISBdgwHtkD2z8qe1xnJjmFE7iLKHch92WOnAhfn7NXGv2AkRCadgK8TuCX6
vXZQeuYY/SaCSAs1+1QpBFHCI8IIevjzCw7fAoT/Hl1/G6yShFJi+patXUVh
rvCsUZx+mV8Ly7vxNPHRHi+unWELQmaGnjyI+Sk5rhFfi/rCFuYkXUSrkX+Q
c52w9mRBHLHYU2TBVgANHro4OnbBddcswqGiGKZ5SZ+ExTeFJqrHVNS6qR76
RqWpIcjOaqYP90iRYBUen0Mk12fd1mRD5BNVcxUnKhmCqQyYiRMcLDlupslM
NEXKVysW5jLwinPDmuQOITJ8QmfDLPz6CCH4qpulOb4tQBtKeoR570Heh9op
+o2w3b1O/0cbO01Z6MGwCGbO6CIlgmrcp1saV1yQwuumSssFZlxNUbNgSGBj
v8rNqiw/cbag9r+O+O03dy5yiLww5AWaDqY5E8UAX30PedgipgCMdRJdhfEG
Fs8yMxm3KtBZ4wUYDiQF9KQ7TCSnt6zWmKMSpgbFzYlK01rnvxk22H3Y0QTg
MXAcqMsm86nWp3QWvdSa9pw1so1HzGWO7jmAHBnBpGqHOEXZtJjw9Z1qWmBE
w0EQJSUszXLX6LJg3D+QFhrATQHzOUsagQrV/ZjFMw9bPDBt6UMInBR8qXwU
nuKwz5iPcHOs9mvP87lq7hpmH2xdRys5zfrNhnog1Yo57u/9WuwLHKsw+vCL
l7RNijZwdCTj6Kp3NyfM8jFrpFhw4yAlsaedSsTme59uSNz6xepKzhQ1zHIQ
t5MvghaOGXq2jA1G45v4jHTmlWD7EKSumFv0Nmh879oO2aAzl8Q3fpR0rtwC
0R9Z5iUz2+SUfS4TOy4qOuvMlIc55jRZegjGT2R3moJlnopETyh1Jbs8h7F2
J3awZXLSzjrPz/EXtpoc73OYoH+oTM7GBXHm77TW3TO3CIF/5ePw4X6e/I50
kdAh/ggz4w27SmDDA00A+qAQgM0qaXbK320FAv+kkT2fgrNocjRMILg+iwCZ
W96qlt1jxax2wTJFoCJz43SWz1YCsinu3ogkiatoDFy7+INe6pTrHsBwGdVk
ZPgGrKnuzX9oDVIRcorgjmOqRlQC/UwfkmfZo8nBY26T+UzUUwM0Vl+K5VY3
nD18WJgXCGUj4e1rpYT/YcnSjN9K6ISQFxEfNTk/ZpIlPaPnHN8CXDZ/ZFBE
s88wLWaif7eZ95zc74IpBeBQ6jCtAdCNPJbVCRdLVXMzdP20TeNJ17FQ5Bwl
xS4+lGhNkNlExVsqq5qtWsmj/MnMBwGoR8dba3c4A9XeUgM0b2oX0vSovU3n
L3kSOFtw27hMhpOD2UhbPqD3appz4nE9L7RW7fKA24Iu+kPHw7Ufc6zAbt81
K4sCS2M/PpAs1ehXy2qZp3Dgvwec8Wnr/xZvEfWrMpN8GQEYMxNv9Ulv76XC
n3RLAjCKKLT3sGaeGTHGlfx1LSp6Adft0RUqV+SR3Od8nOIXIm6zbgsnXbss
Ei0ZLbr73/kPZIaV2s83lDeYsG4hnUY+Avowj97pE3jNaUuPupdXofr9CWwM
Qqxw2BlgfphZxzc9sX1z4i50LBGw88uTNlSd7qEqCzHWkYVwVjdLc7fdUGBd
C481aNan8EeNRs2pZp6yfV9fsN9Ik2fCRQz7imWJ7ZQ+xUY+2DIttA6rZhFE
/e2jdhu+138UeVDT3m+xOKi6kaz2yafAgma4mixsbBAAVuipZ/Mycq0/IPQc
yBUJBOx3PWMjGNIpwYvf0U7fb7CXjDkPUeniErW+g9YZujtl/gJYh5TPNiI/
AI8ZMQt/5GDtGanS0ED1y4YRBOJcJ8RY3zmL6dvO0tW6UTsv+rV1S/W9nnzD
+C0IsuoWD1IZTIrMYbMXGtj+EfUFZpIUjRroNRpyIb03lFPuEDnjk+UPP2eH
QTDJsarFBdlq9GZywyiEpcLsphjahdoRM9M3IqPql8OHMEwzsmwJ2R2RRogD
oevQAEIs0fdlBvUkb86XtU48sv4mshcTMABPyM5+qQ+vBBLPQ3e74Fb9khhc
fxadcQAvJHfadIHmJfL3rRaebUiMLRcaP442ADqHelXpcw/xB8LDGZn5lFfS
wlqrpYKuNE8/XFmnCOxWFL/mFRZ6xETMe9qyBGDdqwlBE5RoBEjH9Cl2m7FW
4iCGsB8ebr5hmrQv60e+4JIvnAirZbufOUikOaI4R1fbPRljdNysR5p8/A8I
kM0wxPZ7c++5Sy48iuchltaqo6U6L700tNIiKg74XZwz5PV7zxbQGRKP4ifW
h5LjRqshobpAEbMzc+MMQAFXprKptAOFAdJFM3qM16xRXJ0+4ATo8ZX5m0nl
oQBAizQF9Zm3fyy7XHHVi749C+mUkojoJlnuWt2LyCx7IGF6Lg36XMqcT+v3
wdeh7adMuY7lmqAR87X4E+gUl64Hu4gGP6/i80vM8SiCZNrY8ZwoXexUPE96
jFJOOo//meGjyu/UfgtvTeuwPbtiljXYNQparzSL4BjuUak8uj5CbMJmlADr
AIDjdxX6XxKVZlohJfdlwws3iNZRAe5MHpnJCqWqvUQnUNa6ttzCmhx79ken
0OpjbO3eGIwHHnGnj5F43vH6IYTeanHIvrMTq8mfFQcUhQ30TLhP9NAUp+ZR
FkmvWWKlJ1cOoUTAQVelxK+rRAyFoORcr5peyZapmfvElWM+kyKSRYLoJlpF
BZLfZkt/U0HWwXqQhyT47vWrrl3fup7mOO3RgAwRfBeBjX1Lablgrm/iwD2+
7ON3txWlCnB6YShBk7nQEb8XumrIeZmZrLs13yzdRkryFXxo1KXnGyqg9Tsk
nmMv5Pp4xPyK4IFnLdcacIxDK97bUOGpHHm6pfmS0QPq9rLQskyv/DZ1j5+o
KAsW+gGE3n8zoRUh3apLv0gMim7pKDj78AiFx98mBNqscT7fEUSLmKqEFAQj
XR1l1Q6GDbQ9tgZ2QRZ4/iBF4tn0aUYrM6oH1I7wQf2IPbxMaRQYb7jeMOIn
jwmtVXohL1K25/bv+2zcAYTVwjeS9a0sPD4U4tXgTqb36wuEjYuop0/yjedx
3qzLeBa8WkEVKy5UjGLTFjTtuH5ElSnDflEBt870wb31lC2JY7ni8soYIrHK
hlRJg8LKoNWqLZgOooX396mZSyV2ovyC/lsnuoMh7eOgpN3fcaAdk+r4HjqI
S4fEvxJ3wL6lAl13LfB8kkWna9w7P2WP87Rzc2RM1uN4Cvad33CU43vH2jze
qpXH2MiF+iF133aWaTBQam81RkjCdQcWKKG0Wjvfws2Fhdp4LL97WoulATg+
YqQ8vVAJGiz9lHpQ8KbTn3LvHlGgfbT4HNQzWFz6uq0DvwMzqg6EKr1sbdDa
ki5myU9PtUZeujLY8olmoOoYNw80ocSE9+MqQvEUTcntEbL5azWyTUPCXAgw
s5mL1cOd/0KAt5aggKo3Y5iONJpdTJhYurnjZ3aAVazf7VINq5yX9So45ZOE
FFUPNq9BDtrNMOwwzEcKTtBq9TiUPid/Cjno59brAwoU+pvjQRdsS7bbwEcQ
mjnvddFm5Ly/AWK5ED6keIbWrrmeJ37YxZNtawYqFywmJdCwFxNN0X49dg3S
8fEnldVO41ePfXQoQEXm8/NoJeVkKd2flU8Sjci91EHo9fXgjEywxW64P0XS
9JIQp3c8Xgoea6iLE/SYVG1ctPseWCRXnkptIFF5ftLh2d+SrvozgvqSvSfV
t7AbD0zTQ+Ws1ApFsifsr1TnfH9jDZ9ddiQ2jnpjYtlvkBPCxRAnHxomk8/E
Mk1olIKKGu3U6U0KcflNqYPaGBYdx1NMVL7SHnVKnXEwviHq70aZKQKOEw12
d+inGqzVGGvKLdZL6EZ5qORydf3cn3XCL4f7pOsH7aSTNMUQJWNlMX+ycJMx
UNdc929+dtdx0uf2w/tdXsKMDDqNbk5sRK7/Wa3mD42QpNiuUHtwQDPd8mYC
kQ+Fh4WEH8qN6xfvjMsDWaSyJAqaab17uTRlSBlr6Nb4XfJ2gtfHPuYHghRG
zKYZG+vZkHDXCKJjomRGRTBUPNe/lNB4Vcx9usUobGeAkFGeNRgYncSYDggu
oB4OgLv/Sexf1uxnnQ2SBbKigj8e08NKhREqq6PrybVywzep0TJRwIDkJxGt
urcGVfvLR1VnZz+GJhO9H5eOjocrGBFApZi89vV9ovQRBEK21WYfeh9Zp1h/
oc1HzFCf7F5rsAeSi/a1vi9nAMWPahw9/tB4eW05WqynFM/q73v9v4zEX6CL
eaUCVukA3rmevsMEyqd3P7C8RYIk6UPz92gTAMRvbiE+q5RlMjjpGPqDuhny
Y/Bt7Zqa1IjDPa1tEI7NbeyaQVu+U4LMG2LK945BEvE/pMUUPSQ2RNqS1UFa
YoaFEWHXVWR3IWeswmF2rrFvM/2c8gVsSl3k0nROxKRKRlBLOyNpMBg7utpj
7EYYUnwNHsAiuwZehMiJPmVUiDAiCqrpc2x1LvYY0jOD5J+cA1MXVPBcdNjJ
ZpjQbDPdXtO0nSq3Nc/sm/sYXPsLmbRBglMp9KgSilJBwZuVjKeXTgBYz0jX
tqWuMRdRA27GpQsg7/B7LqAgrepk/u+BwW3g0VfanF7/VZ6HT9pRJHnAhFUp
jVmQ4MVs+HibIBN2T7qVyF5SDMoUhekGaUYG9vCxldnMaXF/CHqh4UqTaWLs
15DOX7t37GvkN6R5fr5VjhA+7ujljCpjI2pKPCx+HEq33KMTlvgFH7IvL1eK
hFxcAGwnsbYELA8bhaJcZZAmrSxGM8Irl5sAxatcgeJ9iWbmWY0Ar5GxPfVN
W4TfdtWx41W/I5F3NHEjilZCUs4OmD2mx8YsYQegiNgYARKu/LRszrubXT99
Jr+bT3kMGx+IbvGR+canDSH/hZDpFm245MO5JRD4KujwhHEnZO2tM7BuD0xL
BzEFWdXVD2p8ZVySWEA6cgG7nZlSHoits2eO4b6hGC8eynnfx6jXfMQdDRSW
ZpTeYGqrQrzXEO9Gucn6sGODBBfGUGWMLaendLtpyZ3x8ydf7PmYVwuMR8+M
TSNgHz4g4d5p2hFuhIF+ZSndtceYExE91vn/Mq4AtNlL2oI9fHws/E373KK3
hKyKC+OddV5tdszenuMDHyiRGB4/k4zQusIIRw3zrnVAKEpmGYDxnZKXY+Gc
h4WkhD1w1CuU2S+EYVRGlZOuJGxrms/TCrKaOj0dav0gNt1yoYk8omjhkCBs
sznzd3NCZ7znkijb84g9bhkVAiNclP21V0Xe6qwMKHDB9J5lso/6ZuTCDOlK
QhXaFaOFH8y8c5upkuErXFgMgWxfAkdlqsBYp+TEu0FXB0cDRm1CEvgSZXC/
7TdUTK1/d6/+hfkXN+3I9oSM/aI47fJnzIwwHTigsS5ZtbzmieUOhbM+herq
4EVraxu4LJxkFMNNdiSIURn5zAL/bTBprE0nIY9uDbB7T6ydMLV1PoxbanJg
iWnPZZLbqrVz+vKqtU6IpPFloD69lNceMuXlRmSa01k5KOnHXRsKGBEp5Qy7
niB/N3P0sW5ZLo6CU7R6j4oUDi7KgA58FhFx7oHE/Gzz1Zw3eBiLbU/1YTd7
89xp3Ua5ybhoZQNUYjBi5BCFZGShExlq+cEbizkJYvd7RQBXUR2UrlK4ywbl
Qw6TGtLJXdNA06EfqlvkRpqMwtTxGFhd1Bew0OwjrcMPaMRRC01Sdpo8+9rm
qcRcbM5sPQsqBQNxhAbi/oyNuJ0dx9lrubHZ88rVtgu7LduIJX/Pl7Mrclyy
LTJqazAKnZGmDpM/ZbrNKIxFBdziN9GN8KN171fP7okI8U5sQXuBdkStkn1P
sUuZ1VbfnOGJUlnzQFVX6wLzz3p1ivHbIdfn4IzwEzI+q6DmO4632MlQowSe
6EwKWCgWHqVswivLXWNWD4POsD4pMCmbzXghWZMp2E8HzsBtxbS+hUDf30qR
mj4TUh5/JbGn0ghFFP1LWKGE17FD68bR4yxHGwSA5iDDg0VHg79dqdBJX8f7
JYuj49Ju6zbezdTcfVjycrbvXymyb57GXYUc4O568grPHM1arzs4tODN7DR8
VudSGqTZGbPJoJ/0n4v9vYVZj0lHnoER3qFD1FmqFbzWbZDJ8j/LTiNodmGz
AJIWEqNRVIAc7g6rWJdbjgCXxo8Gr2knOE0nLbcEdhPZQAWVskYMioPdwnm4
03Cq9RRm8tRKKqg9eLs0uKxHqgU7Nm2jwtaIe5NlsmFYa8aCg5qk5ghvkztT
Sv1Z3gNV1RQHVBC2ubafSXbACUJWKR2PQxIfqGH8353cW5t4G0o07TT2+wry
eqnBTByw6U4jPxISusaUL6AHuBs7n9ihqtaQ0FgC1E7OD1PgUnUrH4jfgid2
iKajYLY4sJFkuKqb+ASYB6/6qQI1Yl9oEBtrdR4ZRs05BnB9lBSZ/XZbgpcH
pUal+2xln7gSLvEJCD5cvPZ9/2CfqGGcYGJQQaowy96debtIWupqanK3PVia
zu8iiH6+43hFKdUL9PZA9TOcTa6HngxkYG3DXCrcWwojnpy9MR6enCy6KI5o
JTvJ04xx4IKKiz9ulcFOS/rl7pmPFPvWiHePu+sWWeuE02dFMXCXDQ3Ts26g
RmEHE2lt49EUPKIAnCw7qAqbEbOw6yEcgqTrFStvbJFBiC5oBx3RtPXoL+bw
kSbFlQzfSZvXriVHbzHPFq3Vo6OO3sfjxAq5gpAgIQgSRhJy0p6s3c0SUTf0
mrOoZBlH2Z65PCDnSdFp46oTLcqD4TGJCaY50AaiwaN04LbDF0rok8a2t94j
lygA1HPIL1lEK4/06El6HLMnzdTDpK0sjdIccfNAg9Ls2KvhwIgmYonwvQQf
j6dzZkK7vi8Eez0mtyh/EYJZWRX36w++Xrt4hrlmhJ5ejNI+06DEbnjFl+Iz
kdbKbC1yAxrxzwHCL4cVnoNSra+qYkIewuCIMmKpquqfJRvPCG3h80ML+HqV
2M8/Cpiq4pTOz9RyCz2yoqrtzihGmqgqcoQJCmw3Gs7ExYbemCsfO/1KqANg
eXwNJOHpP6ejf6J73W8iMY4jsxkmJG5GUfAN1YcTNmNsq06Yk2QZbTGRS5uW
lTr0FCwzg63cU+bXjqTUC361MVyEczrn6ykoWIqjsavm2dFO4MZxp3D0AcfP
2ddAT5qgICboBjGOgQMGdz26tOYM38xdT0hVDiK7Ffx+kzZj1Pd3UKvm+pqO
vmJ3a/03bQQIBzu4OMGz+GtXW3OPHtbdS1/Mz6wpVCYrj91juiqp0dJOFXJ3
vekty8/JFQ4/tSy85c+KtCfuaRaX8iCqWZrDUnb2LPyaFiyV46tylXKer1Mm
X4Tga7jyZCjnN7HLPKz/G6gnmtozWaULJHlRXRBh7QVeBiN+cjtAP/YdikoC
sleSAzxC5xy+gh4cc8dpLs51x7calDfjub1YfG1CG4cKQohIYKigYa27CsaT
YivWiFboAZIgMY3ZogXlV9tLH2ZP8/4ubyDON8Osdcm72cD7W4QBD4pre1g5
dSKNvU5dmySMikMbdQFQPB/t4fuqSehf1syghhka/keKNZ14LyVIW8WXESmI
a9KurvhDimFEVFiFhPVGW1pve63LBCJx/6asTg5Rnjv0ajimTOI/NBTnwmSX
NPAFFG8flIwkzWlEyRW2+geForP/9QVPjO8vSNUyZmv4Yk+FciJvQ/f79iyK
6KgSdGljeJVMoIflCjPBYGe/2qmNsikoVOB51elkqryEDxGY7fhzilJiEdNa
EEAVzYUcsLNdEVRc6l8Ueuza8xwq40et5AzK8vQ35VNw2ls5Y5RC1j8PqlW9
WGqE42bdMyYnQwpPQTrjW14fuPrtUDAI2bVtcPmVpA1zT5O7izDbDRrkO/YD
va+zBMeiY03iP1CwR4dfhab/jBYVe+ms25DUNMLHnW2fr7NZLP351sFXzlEB
3gl3rBk7QV4UFTZuX++hV8iHVpwY+gGY9fn1GUvxGP5MuMqqFjv0NcarYH85
GYsmDt7RY36czpMb7QX/Qqd9Rheb6uuWHqDPd5rvJ9qUYtdFxcSvYiod77BB
SCBfBzX4aK/yafVN4SsC5CbV8hPvOnwfMTx4faHFS3q5jDhNs1fRtYsTqqwt
zAJ9+OEyk9ZcBJr37RcC5NOthqQO6AfZQWTghuN2wHC2+wU//TpQ+RolITuE
VAb1S0azK6GgbA+ICKx74mnaOIVyTJKGsGZqt5bbOBNZej/QkEe5ef4DQCq0
4uJT2v0xG4dT8HrFParR1zNj7IuyOOEc8A+IH4g+w8WoRDgg48tQ88bUHH+K
ejVQdyUe8RaF1GYwRWWJaHJJQ0dhyvYA+8bajnTlQbdnMhhnI3MbfoM+kVfA
Wb37OCN7BQ5Hl+pW3mds+JHa+irKME5U1X+Xbs75ThhDihOjvyqpDtv5h+zb
YC1CaB0eVyhFpZB5gDVhvl30kHczazZQheWfudvKyknXqojBE9Yl6SL0FHYt
quIKd3AEG4n+yvxo+DNMXqs0Pst+MwDzCeb2LpsBfBWA7WRCPou31VKWUSAc
gNwrOx8dnwT55/+P9W/Rvy2z32sBkVTjTzzdatPrTYdtCwABmGlcYmF11xUY
SeK0lwbIWfO7PsQrBnzWtU5399EuhMwEMhE0V/aukY+56sxwapULsmm3xsMc
Oi2radVk0kZRVd500qBqJS7ZoT1Ep1szYA9P0m7mthJeEVODtF9hNkOQFXtH
3u0/X7MorjJQwp43+c4Ur3SPjgVopXSijjcrkCwVUIvSKeDYRK7NIC231cCz
bYLrPXIDOQPj68N+ylSO3uLdeDgIPQ3gcSDdVNcTmvHAxTCuWsYDhe9Tukdz
3RrLK/yl0PA1QyyGPTzTMs002ds0ut4P1ut77lAI6d86frHWU4zHxX2Olsis
JhPeCaC6V6im31mFjtiqaW5uv4q8yD2ReZHdvaOMAROnEf8PogR3InwSHw0C
hTlmfqjdnUWTjPfnQR4MVty11aNfK+iDgMuTnKOrMHr0wsb5TMPnkI2eHPBK
OYH8dEuKB3jIBTH6v2zFpdm/rZzXJMIwulFhausIaimbqrkgJKXMRxtj4MZQ
08r9yQ8YPv3T4s27o9cBgbQD+BxMTJB69DLEnTS0slBytCU6zEV/zInV868Q
XwUJR5+GyQUqyugLfWPaiwV/+ts1T8n7nIsHNhKsNDiVPm2a+iuf9M8NPkVi
4x9MBFuMav8ftw9EmO0xN/p8g1JaWi+cSnaQwHwvsEujueyCw3cH+plLg51u
tRd2GhhFrfS5fOcb1z8oTxuIksrQzVwERAhEE5hyKcD0O81Ef3aNwzwHYLgZ
DzLfCuqEFjzJveBPa6ylNfKQ9ZDrmlTavRxYpPrFVxv1OeEeTxaAZ6lIPRqI
YJBxGEL9eNnSClWpZm1CZQjSvlhURc/2reydcCpXe9g+vx7sW47d4tNEzFRI
Yjj0cQSiSbsyl7ZSbGtIJoRlNyJ0eZm9T8t7XjDHbrnCeXCnLtvlyxspictf
be1OWuWg5coCGcaA6vyAOjcwSFml+TQlBK/BwjHSUjOX6ZBepFJsCxxUGoJr
AlAjYLKR9bT+NOKe4ZvzXYRhwLhE/tZMZLi+a1mNiWUQ7VYXFd7nIL1H+0zp
I1ZDVgu/3wX7LOjF8btk3tDG8ounq849I7GtNOmtZ+Fmah+DUPxAle/SFQqD
rMXy2R8ojpTjopz+PTvJW/+h4RqPurBUIvvFvp/Q8LXYlaKdjckxBDK9drZl
VW3sfp6YJyNd4GZ/LmK9uh8+sMNBIZD9cYiXY8JiLXOoEiBvjspPlK8+wdTY
UwVOU0HlsrfceNQCEjOXJ2UqBxycMBJ2Dvst2b/j0wvZtRLhgh29OdZ0uUHa
mNNYlhY1T4cf17rlp5mS4RY+KcCxeSwpP51EfCTIWsxQ3W6mqPHKm7jsZaX3
r/1BSK0LE79rHTDHPBTjPkjphqKZLOUQC9Qd48rI1j/HxQBDp3XqIuxRVTnw
LflkYOrUyt1odHHWEk+yUJfXasseO1MXCUMFj3Ydx/+NJsOMBm4AEA2Vj34X
yccBUoyPw1pLy8l35KbG5rqiepNrjGRisZOBuB84XnPY71lbtXdYUY7vFWfv
VOsLMyXYvQs4tbJSYZ96Cr9dBtQfdvKXVTvLDvY1QJI5jlrxSdSXaEKz+K5P
rtCv5HTzacvHygAxxoLnW6ottGLO6e/x3kdCbfmfuJx8qHFWKLoJZ9Xk4u6J
34lcFiCt3+bLLFhpQctJVmz5k+R9f4tjmyTLvATtvuJ80847EuvUdxtfTTjc
/3nS8AdedcmLG1u8vni6D8K2Ap1nrg3MvQT2lmNXgfT6APsqjPSzXcSzXDwR
nHc60d6edDlQ7WstRXBhyn8Jp7WWWTL92rSrsgEmyJ798zJL4z6fYCkwuTIT
tPfZlutuSAjGvg2+onrTbci7diyZ4UBfObTByhstorKGSxwyF91Q1lL0IgAL
ljOk7cDRSgiQjB0cBYWeVv2sCEubUZR4f1Y+7LzQMW/C3OvbSbsrSr4WtlkH
sYKZJ7mp4HyzYyINI7weGEpMkVqfkeAUMdIqoxx+NLNMNtGFCRJ/99CvaCYC
vM+pCYJKzjEpR6CrucQpZQoEpMUp7Z+1zAS9Sy0TOq1ifjpTVHfq5woK7FfW
Eqqzw8+tYACJ6OFu/WoL4NM8PRLrH5zHjMJVunfD+KE47wedsbMm6p3ezGzG
tW76a31b2yNGcOdW3BggOIuQOnYP7d6clOaWDnoaPsrKsRQ3bHZy9YKS2tFo
rddpFGifZSipkmJj66sLtsH/4zOBCXp4ky1cf5BsbtEX7ZxolVWs8pebTMpx
9/2jntC5eVzyT8J3tZlLT2vj1zT6kwFjt6UbKoYDDHBmMmjQQ0b91TnZjzIl
VFNe6gU2LDipFsPDxan/riZ5/ukDihJJexxmi558hdo72fSOWth2k9I8a/c2
7j4h3MLm3RypX0DXtWlauh+UHAW8zskAjEKBRp+gP/e1dJfLp19Z7oZYMcrl
yrJsr6zlAL0jswrCbA94cZwsUCvIUsT0BmppbI3Dk2izbI+Dkd75Q2uLbj26
QcpyCALaB6GeGHvJDIWjVd0UjDYOaDhpGgTCtLOH5R9DQ/EOWDlQz8dsbBpS
rNOINKdgAWlea8XU0o7DQqmoOg+3KjhI2wECZWjSs8oktAG7RC0krf62mX2f
OyPcqJYtw89gK0OESCcTZvA9svNs54RctOmZ7xfdGJhqErlYDREawTVIO9oN
B8KO97rZBX9m+zZe220EzU4kmvGcC6/6666ziopUhQEbGi/fUZB/73iI/4Q+
PP/aoEF3kdjPZtMxQjiMVvrQu3XTqS9Q+LPeoqZIh2zkvb4C7v6AX0kydpU5
FrF1wMr2uNfPtcvAyR4WdvB4goDHt04wq5eTrDyAceJWJhLMz/114vfrBV5p
1jdHcEVxzP3dHNnj7Iale4qjC9eY4uvhjnjNKdSzQmyEY6xe0YO20fzM9aBL
IFiNWzNl9bLuF/oZJWdbGI/UiT+v7JMethjUI12Qlmi6bYTC5nouJO63P56B
12raekPh7sQK+uOY/TBFw52SWCDtLC+OJd0jgh0D8OTgcCCuqT79ZynbrNce
Wp5p+Td906GTIl1mIBPJjLkqAKlsbNsI9Vgz/g83aWlqja5EyvOJkihw+DnI
q0o/idVSjo2pTrlyHM+lSsQeKm/6LObewMYQBqHYJVCy5qbSAvNk5uLOcTyP
5PnYfvOQIBRC5OFnL5dDbO21WSKMM8XjO96fZOqx4hq9w3zi+VgNsD5P/0Jw
7Z8XJdWTiUbOGQMQ8copsvRk3m9fN9rkKcina8JsHC2WXSuz7pY3WbBfaMH5
K7W6JNiGblyakzv9NUXPZDsCwXM0nT++Ziq5Wp86xEwvVS41Kp4NyoEsNaUz
+tz+stzzkJf7D1GTrJrrnmiLifsusN8ZTha3NwM/afvA8UsqATJxssq5SzGz
lYUMCGbSj0BnVCLrDML3dP1piISA6z4EcLEfDZOnARaUKkWhKrZVvxMi/u+F
ARy9GvfL01Ys6mWKSzWpGFEAfoUvoOMGuDD5FfI1xtcwUg5ue/axCm6MpF8Q
K8RDXneQIa7XZyHRpmrZ/9nSn5EBq0QQ7kC68mrQk2I8hyXTL16GblWgw7qd
V+daOBkGf38eMrpObEXBj88kgq7JCMwaB2SL45lL0XPECk7izJytwBbKVylM
CDJVLqrxQGrt/0kYqi8ZkMYF1K5yEnR0jL/mkfAaIyHm0ps1aQgqd1gZkbOB
c/622ZNDaBbHbjCGG137QElaGQ9L0/2TY5h4NVZySltmV+iKZE7s6RYD0hNl
r5ubTJmY3i+iOVyby4j8Yk8nIZoi3+JbkxbmZfVrRDCkKG7yQPGi2SsPzd23
MYnEqNVkE3mBxOqvKprK+Jk9oM4cbAmaPn/ifG2a2mJgr2vbNRphtaKbgYx/
soDulkAVxNGD26oQGMrfxEK1JDrR9rUq3SXXcGTRVd5QY/lE/QJuMirUuTx5
BP/TPnN7f121PSr3jZZN/uAdo5mqwxuOnOBFhhXTMlwx5mse5v9ag4Lxl1wd
UuLBa/wfnF8nTrAGwBON0Q7VdGEAF4xc0/Y5d35Pav9eQHJ5rHacGQXe7z5a
1Pmuok8uE23P40wwbP7AHPgMenWSFW/3QLIhmCIek3Dk2gheliyn1DOITZd8
BUXKFULaPDXb6fJvpJeUu9OfBeq1oc1++M9VKkZHYRt6b5sL+5AbWcPJlh2e
vgRxd8OJ5ClWRBV+6WyYFB+q8WL5ZvK9/TcyMOAVzMujELehKm05vCvnQSUb
fVkvkaCQVvds12ZxN7RzzjER36LPUYjN3zBsXjOtoJ2zso4xgIJ0VtfUQ+vv
MbYiHoDGqnQZx7IB/bkdirEolp3p+i4nvj6c0Qy6gZDmEqRS+3od1S8ARew1
qE1QQ6z4c1V7aUtRTO1fEvLzKgneugLCMRrvTdVPD4uU0hANbGfvI170gTk0
CLoEi4IYEiYu1Dephg/akTcTnxh60QLJVcjU2mrOcnzFw3SydnKTLdr0Xs6P
KRtU6e65CHjp+K9qKZPyu4/HTQUD2TeWIOBKfS8wYtNzqqx774bApdUyI8er
sxnqmyahWInFYdal42C+qoWkYrww2cVgKjO5CASIyF6rgRYX0/R7sroptWkD
Y9CXUEDhM+vtd7qOGgOnDK4l4XRz6REuo1aNcrNCzmeuZqDdd8q5J6nnZ6VU
XBdERo7BESnRTlGqlvfDa/mvlIOwf1NvSI38bKh10JyStnLVsWke1LfgQD2F
BY/Em0tfTazpmpFXAl8rkeQTLD8DWAwRaTNP8eocujTUvMQ47iWVdfQe01+L
wBXtebXWrAJGVZbWCv9CfwlLs6IYRh3U2yHLGPBdyBaVIT4wlhLYdKZvWszN
uwVhEOUEE+hYIuy5eQwMlgGiTWoyws8CGA5GOFFMEaz+Rp9oS5Ej7RMjxWDt
oFgWxp3YMV8QuOYiwtg7zPBB0Nzg1YO23soNdmLrzZWeYe+QpBq8SdncbeW5
77qtVCGY+FGjPbpbHOEHtkb6G3F3v4IuvbEVfgwnMP2mPUGD2ISjIkyVCCXR
2DjMmOTQjQ7K/uCk2KdUQXRDi5v/dqgWc1WIgMUT0q2E6ySJlloRRC8QgGmz
J6bKN/NnqkOaEL8TTFagIpuuQQmIcPM2UY87My8CVEstYlQXnFdHuePbmeON
Hx03Tv3nV4cC8mJqoSyfyVHdo/aX7biU7fkMibqNYA4hFaA7d4xL9whLRovb
MK27vVZIZXxgBFNFd2j0eXK+DSQHr5kuYOa79Y860gyyDErMhZ2Aq/LrYxUg
sZOubi8/HX4vqrfQRxvp4hos3q0S7rLOnVbFelUKHdHnnaYYnt+P9xYupgiH
OlhojVwr1WWCAMxzErCrTSmDU13R3xUtUY2nGMt8cRt5AfG7T4fLnMTqcxGC
jpGKwWDGaNZDy7fdL46ADxhFcA0pr/Wiw4r8xsSaWPoayfrutNCVALhlpHin
rqsFBi8FbLDcLEAEIqyKeaz4u4gFaifbCEdDegZ0e64Me1AGeqeuwWncB4xE
G9ZfOIRkLRx4RCAg9/2d8SCfbRJr6PsfuldBgNjZKi+Djf5oBC/bJBuGw1Je
NV4xtHdMM8523ol1NfKX90l4sB486vwdvCQFmIrq6x3VuNkaCJM8fPXT6hR6
J3C/TBlBKEqq/szUkTjxZb+Ccdk0pkA7ZkSV1m9TmKo59BX9B7h32pr1zpLR
FnOssDoAVr6PVxUPpPF1HhueQNucxEvekQDmGWCXVd9aBUSWUIPLQX0+lhXV
qHBPEmOnnzrEVB8suVc9yIZECJeEqYxcUJpNGm3tCEr4ItHGHToHUW+j9Uxq
Qh/5fbrivcSciWfJFqJ2bV2HsVjnKwUyhEst8rCSAsHcQenOnBrOvp2+zrr+
FWzNF52x7HeB7ePYLLVXNs4j/9RdBZYiNxOISS5tyikM+p59a+vMK+tZYmci
TLvdyyNahHjXaMKcD5/IH+sa5OqvkLYx+obbhuFmTh1t63NTogPMbFUBrhvg
Q1hrbvG4iQ7AJpintEKuZ38k2JfaO92sojHdC0u7LMcoZV/+wWPQ9jb3bow4
PV9RQENluzIE+0HaM8lASlwTgF8dm6+mbbQ9Lf9jgkmc64jxhxq2qL3hecyr
2hkyeQCtJQQvS6w9tPejxxrJQTzL7T0SPIU6elZzmF+xSqMcg4ZW48P9m9eB
bTHEVSqnR0ioibb2/4hUcn92DOQM+iQAXm/tMEvqjXSjpcftgGX5IOOl6fRb
MZjX9vDlW5fDi+Qp4XHzk2IANP/vbZ1aeTiWbujrePEfPw/OT9L2PW4oQ1wU
2fJ26PYckliXH0z3LVmN/u06UpggBIKkddU4LHoD0nGyu1nhnOw+C9mf9Cf2
NXzuh7uc00JRvmVRVoossm53Pq7Pv9wfWgIoQscJEkfFwtMIUoLgUz24XMWp
DuiYAX7tO3u6Q2alIlRrmvWlIE5QZ+E7LNQHeUiDQUBQBYU2IVLxpdDGKslI
9gIg2KCOTB49hlpxKiYlR+jEDn9MnMtndOikapoyPQO5qm6z3mpwQXb5Aw/E
Ih6CAt7T2s4dMOI9WOId8iTcqBnMo4VjtRQ6/CYI8icHRLqO8x+lUviFbh/S
6hrmpepiD0GJNznh7yrjLmLtS7RNOn3BdYIRVlrW++g8vDdm4P2Pf6aLtj/8
09ZU6Qgl0tgtLrAD+aX6n8amxViolxIxasakrhz3dfgoWDWY93DnNXkW6db1
eQYLRSpwfEdKA7BoPSM4ui9iDQEBGJuzf01TO/lcCe2L8eNuUvnKYRQfMdpn
OFkyRgQDn3DSvX2CIMT2L5iRGZZma9iUXhaoQLuqnXTZ/WkvDXZkjkjv5viV
WJsO8yiKS4fpYN9y6+APRY+Gcc/bQvqwoSww9AIl+bLGBkarTAPE2Ben2IH2
1P+RQGr1cJF9+vKImeBXK+dTsyWcVg2GTJYFdIZE1HJmVrnr0rNtICnTSWLj
WaHj/E5DJ3b1sCpwXmaI3vv/OSFCf8lwQ6irTq5EJMZAdYS4UdEXHC+iw15P
UmiyQ3u7QAgabqLYvVaamDoWnetXBqsSH5PL0r+ykUUPTwecTNCLs+IdGCMV
7827kLvHdCWpDkN0mwj+PkkVsrtWOEpY5o3kSXq/VLHtpZ73cXxNxN2Gk0sg
7jaskn6KmOIFVCfU1ZB1iZTfN1Y0PaDXQ468jv8flGP8zgW89m3htp9p+cPi
9C8KlJ7RjHnqMWCck907CHGlftLgUoNEuwo+oWMggMv9fq313lyMvCqwbA2X
1DtgD7jyTHFdsitjbjPQ106IP5iOBI8xGFO5BitjdLfxPYhx/AzswyBBRkrd
sxcbFicYR/2JG5gndesw6Ki5MWZCW+wBgReiTLHi7AUXBbcFd1Y7ePdjrhWe
73SygFhsBTnAi/UngNL00ivzjsd9KYHLguKPzXCG+/cYS9ktzjpdK+1A8dIj
lWr44QJGpkceZLBKdc+8aUiwgQGpv5ZVdcjlSwVkdxNIeM8in7t0jJu41i4j
wRj4xk1pA9shvWxBlzl2gTfBeNhVEYl3N/sSjFF5/mIPOUYH41ztFr2QT/ED
ZRVelnezkrYILk0bv/GuMySwZrZ3aUGdvyjC13IxOh6rZ7y8lLaLqkJpCEzX
dd8VdxnQXOBiAHv3ZqMCsRaSZn4x/n5fXowfYZYR8jAQqk7RFjK/dBa2dmVg
u9G/ezYt2nJbOiqTSjKv+9LXi4D2rUBlIXjgGZXRJTCilo2pFdsWqH4i4I+u
8fLqPfUDZ3WwQ3KjjfuaPZzEMWazexxPlwm8W2PJAvGbcO/vebnN4TG0qb6W
gnDHiYTTkaeCDvWD95cZuW0333aZI9mn4MZZGj7zyHSSl2uDREr1qSG9QEvj
GZwxbFTYMKO1QwF5ntkZfp7NhOaxAvagV5XpGxDcbKjcOPepjIM1ytSKcA6F
QiZMVTGNTyeMO+vpo2wUV18YpW/pQzJ+4djmNsg81n1iXx0Lj1f0kAykyX7b
3Q3F1NT8vOqGVzr+8GnruwHUnRJxxWouIMUJZ4gjtWxQ8Ro9nPmMLWvYOMww
Hh/Zq6sAdzMln3wANo8r8Z4zXZWrn+siT93yhJLroqjemiBen1cjHv+vK9rQ
BRQf0PbChMVQc+59jyXR8bQZRNtIP76xAUl93zsbIcHFO0cI0xwy0ae6hhxN
QzMZS+Ts5lZkPDgjx5x5L3CADdrl5eedbHVm4qYcdPyECIPbkqFpDqr7CFnh
AxanZtaT/OXKsUDZzEWMH7XigWcsfxn8BtckuuZP7TdvtV19c8w59P6Vf3It
XAUPo93TNZ8Fo5thU+iV4kmpsTYBmx3bBUX0SBydN00T9SGjQ/T1IaTtnaL8
NaGvG2ObI/P3vimX97v/gtZuU+vJP1R1aBhgjRofRARS8u/EJdiEOCYFXYoR
AeekBeWmEGH0zyIEmECfk+bmglQQQAy5gOJ4urMwSRovuk+t4K03qS27gUXp
C8C4au/IbTQSUN6qfE3FYDYFncsPlDmBHUD3ZRf9kKxxc2RDvGmwDTqUxk2g
nfhgb08vQCR6LGddgwIeDe6O/F4M1A05pgDp0lRKDR+cQYQqkOmQwhBx4q6M
CzHuSCmpdyqEWqwzfXFWRNYa9ZpiAG66bu31ClneK3Ki2s9+fTPZh2fiKSYi
4+rKfx/5bne7LoW68rXxYtKRI8DV8izEnPowrbHywdxzCmDN4J/zYEAqB3Mo
nJNogKPWGKDhOHhu4R6Iqj4Eiwcw9ZdfYTeb6Dwf19zF9wuovN94k0QxAaMb
uvhZmojH+ghRS07Xhf05A9WZh3L00gtl3PXrDqzUgN3F/7XijWCsNMsZIPZL
0pr4mztO1yC1wGhI5bqM7JIaMEWHB0iTuz9TvchL2OWMUJIl/zhmjw1zJo+F
qYG2VX9IISeaUCcGAabrF5lswdJl/Ct527CeFdkZKC6EtzXJE57alXdmMZl+
tFzi/syQVAw6BJeDGxRy2AJPzQpO2oNkx/4pzLwngoQ6Lz7UtsY1q2opH8na
dLCIc7mBc6f0mRkqjtcMbraBmu4s45kqXTVL3ymAntDlO7wwJffzDlDeFSfE
+1t2iJ2GIiKB9QqRRDgb5HCBmT2pbawu953WTHT2fBEjzYPcoA9T7TEswWfB
DNGgR2X2EYbUBkXGWDlT4lSjIeyMFedj37QpIiNhTOpyBWSRuCyE/Lj+zhHn
zIDanZvvE2ghC02xA011CiaLXI8mOtM3lG8tSQMEgJRXHAItNw8V1WyamMKO
mBciLcTf+i4Ile4TykqfweXIuICN6Qt6cyVsVqp8NfybqRK2V2ealcA4IAia
pBpeJrS5Ynyfi21IlycncBIO5VlcZ4pEBbRIpkuGFy6keHE5B0dgx2Yogxn4
WGdIQBPmC79TMyhTfymRDoUsChZSrQTkc2R9rEjXz2fr/uDRNibkDNKe5RzQ
OokyCh+0jSuO6+e7Wu8L1liLkuEi7MmbDlr5puBpkTEYZpkRoltKTaBaqyVO
5JU8nMHkOkObUaETE91co2M2VocidwKwFD22C0unLxW21OCQVZuFrJt02hIL
rUZo1O1+/Wf9kookWtWS4+bxNC1pX9N4QEoIJp+MzHj/kSYnBT8KpfeixVdJ
dyY54tjIlj6Z/4gcKzrNuGOmSGlwN5IdcgKe1Xsah42VFUnlL4T1/Ad6Ru4y
ZXx2gu+VL0uY4rwXK3a1JWXVYL3wwp7dOTxavypeNqJp4qzfd6M3ePayyepA
ICtwvvBa7kkCAebHKddMvjMZYDSDL8R6SeJat9T2VhaZPqIukrlA7yqjg1JF
Pni7OXxV+9FcxEo56DYs2bhW1y060RLX29h1RR6RSmGi+8vwlmB5lqYIHlIe
rcgLMJhXLJSAWVmdTbEUFCn7aVvhfOQPENvPlxGJWCUr9upEPjM+WV3fYd02
ty1wf+fylQ56eV5sVAwRhjOsizdehRA49Nb9uOH7jqz6LqSqLZGQGrIL6g09
FWjRkdljxunsoyq8CgQLD+pzmswibTKCOH1vA3R2X4j8q613o58jFgwwBpbd
98bR3rujUaRx0O6yNH1ipq9rPD8Z44b8sABMZWXgemk1ZYFvZAeGvKj7cj7R
uSj9Q8ql+7YB87ClVqPLGP3FO+hcVJEIykxIerKkcFNoYXFTAIq5NQj9X/Es
orBkeaAm7z7JnNBWqjFZQ0oJNnhpl+P0ke2lL8/vXKO30ESeDw3llQf8OhXa
5tJT4gwxbylImygyKrLt7ZVxqtPnJULfnkvJwDkTxcIKb4iRwkLCwPLmBrIC
UbDapT2wi9Dy7dFdqTkZ9FSHUlgCXdC/CPrPU7OcAK/ncFcYN8Bsxehc/zGI
4hJEJ56yQpxOVUOwGdMROuXtbKvWFQ0m2Hk15//SGZTIDVSs0mTJVkUgPocR
qtvXHEmm0OLPTKrr54o0wAPuk5k8+HYsNDTI1nAWvhi1I3D3Qal3kNMXTOul
6LjkVF5c27PJcNPNeJMp7IMtwNScmyc1WMxt4wB2tQIsDO4B0o9WqkVWax6j
BZtP7wrorIfneXD9acV56+zer0PKn4gtsep2/dlDShskpxxCFRBag45RargE
rtr8ZYzXO3O069jPNOLrOliJyULA3pqSWrp6IX5DDGn+OhF9lmXiD70NQiAj
emBiRXgQJ6ib0U4Q9KBqbfbXhcT9bWvVly0LK2IMHuEAMOheseRgd5+Q8/Q9
Of1FwySQmMuhxq862R4KMDD47KsCIxdHDZlOad0VKU4o73volexHTfE1p+aY
GjVjcVxCauWLQHV77hZ8T4enI/zUks4reIqJqvxYzFY3Mp3k7zH8xE1bclhE
DA0fJ7/teqT3eglJURrGCatWmtZiqqV9zNYV1EsEd9U/B6TdcSbgObAdSYmT
1JaPB0TD8r6LpRsppUcd3Ew2eHH1P+xuE0+bov7ZEyVdKMxGwQEt2S035Zam
wWza0f9rlbrIkqwnZ9mgdBytFsEOG51mIJJh+ezomGw79JT4dozxPeGDNk9H
kp/HHtM0UoGfZHpYFypMJO7/d7HRVpvUNCxrOU8Jgjrtyf2LnjsQ7HEbt6Dv
zssThuU1Dklcuqm5EQShTMmKk88O54ZGhRNzIHzfBB+4bju0zBXsBwbCEyj1
280NqvWIpqrwyH6Wxd+I/N01RnCwWin2b977phKlec5an+97apiuARP/0w7J
dTlF62A6Ek9SkM1OlLFBcl9yHxNBCR9Vudj3a4qH0WfiVADFDhS8BoI2YcyE
zao2ZfD9QqsZvzno8nV7wLuQUS1YqTa6XPKZkMeXeCKLy+DscOVBSMb1zcIR
5o6fGZQJhLUQIgY6+VZ86KlvZ4RW3dUWFQEuoTFLR5CIzP+B7DzGTJMYy2B2
kvRSz7Nyx2d9uZps2KRz8IRjlRuZ8ZdA44B5sqDRq7PEj0ktaAyUzEUif3Ic
Ue7w38pUKcvMY11YY69fgm8mi81M94/Dq8Vlxn12Hp2zubROtAMeKBbg2SBX
o6Dg00t99MhImg3EAInnF+g4LgIERf0+QXEyVJLShjt2LBgiDO4o3XP+y/6I
eW0NHDqhxoKKKHjEYviy4bRqRQuDWut5JhU5z+ZNIzJ9W7SuWZPgL4zOZoOx
/0IozhZPh0nmVVGTpjXrk4/aarEbTTKaR0q7fAfDZm7OMyaXnt6ror02QPn0
I2GtSHI4FTRsT4JO2NXMluMYjMLHCpwte2yAWeIB+7lHmUpxkLDHYqA9rVol
SmGPyTMoATEiOqGk78PlicBMyd+b9zga3K7+Umu2jwVDnW1LW4rluZeWn3At
afMTbcmkmkOgYqJU0R1p76Vex5rfdao8dDbF33UJjMtcyGkzD7b8VO15pt65
gmj09/bwt4DSqF77luGTuNUXIbg7ck56RPWXd13+MuFGQ0UWbK6R2kt0YLRM
hdJdiFRsUNfvgLalM+7pEZ4MJkeuE4LOW7fGlOZq9SgsAPtIqDlZfq/TC95c
jwmVnCQ7T+SGf2MLwc+1O1jWho8KC307gvmysvjekobZj1Kv+XtnTnbLcatd
ck4bdJnawA2nwXQt03yjMOryK6JMUs9SINyBxWCDyEpLA2LtywpGFNMvpnTR
cYNvLcKH5/wdZO3Tf9aTZjoXMd10iKqHZuUBXUqNmUf3CWMSX+GI3F6+oPmw
a3q415QHmecmiSLSmkvsWsKS8efyhT0gjZhDvo5Ecww3cxkoSf7pYozKos5q
QruiN5f78yUM9rlpK0RoBh1/55vEZLrApEkwsmLnXuwFDN8T2GIhd5Gwra8c
3zre1MG5LSPhTryF8Pg/iNK3QlmHmNjTqr8T0zvmAfaznlBHUEYZH73GcTX8
dTMl+W3329RusmBph+AGsRekqYHXTvc9ZWfyvoMbB9ehifhc5LbFUp1G7v8h
4fuKcaoegnEolmPCHzcjh3L/DDmVUP6NHqMCQsHbgJEPKDU/eHlvjIaYmQxJ
VMZL4YMJHfBy9ScAkUAV7+z2KsIpvkhefQTvMUg6rk/1TMconcnPsZ3ioraL
PCfx31OpEyylKr2lTqw0OhUmIOybJG7DbRPo5ij4Tvvok9Db9ibz0DjQv2vV
B3x6wBxa/igHZVLDn8BQJ1l1ds4IdDLOzssPBb6q0wDQ2185zM8LzI8Ng5kZ
zE7hxY3e7gEc5k60afdVuGdpk/CBeL5RngQMQrmFmuSxDOPpbvkaVbJgUm01
SfC1dMKVVayzi8o9lw1w0Xc0fvam7AdxUGs/BMeBFQFupiX2iQ2dByES3SZC
64ezCUXjB5idgx0RSrD7NTSeaktgEj+AIAWADU3szNQTMVazM72msxoseN3e
13H95GieUUoCYn2g/rRK5bzqHaYMmomGdZWEygLjU345O6kh1c8rL6rEVKX4
neQvMh9pNrmA5OpT2/rwO4d5F9xMVbsRI9LKxOTVdL2F6eWEGmCq+lFkvxED
mmlw/+tHzp44qt9OWwbdP99MfkgtrpTpaWzJY513htE4QdAdnwX0mjvFceio
shZKCr2puOJxMrnlT58WAiDZIVHlQBpcY42Jrs+GJvUmG+TEd1Ui/8lwgcs3
KnxLv0+G3AGD+RD5ekfZ/fNyE9NiTNV6bjmtBTYjhYedCHPqsCxe32/dOT0q
qW2ODdhXSJbRqCnvwfqV+UwItKp7CkKzcHqTUxclNYhS4MHcLgtY9oVw+5Cl
8UQTsuat61PRk5E6Cwdpwby8+mYlvjZmFIE2b6/g7/j1i+iqZa0rxB7FgrIg
uiOGOqJ8cUL9Ngwx1MAcXxE+/9OpJ01NodVa/4Y8sysVmAwRRTZs96loo5VO
ZzC0RzWLCYoCZMBfCIZi5ZzVOUfW+jwbsUpFUzvVNg8wKs/R94bewuqlj9BF
QL0Lqzu7NpDSw9xWItmL5rlkS9KIK68EF3o80P1BRYquzGA+bftslLP4S1UR
w7kAJux9pDxB8p2x1BaMglbrYsanzxUwuwvVojxZKKV++PkroGJtE9sOugCN
6vElebBfz7wjM2tjY5O6G1z2oXqXWzge3cJiaGumPmCVLujhv9FK55dh16TI
J6Ky5phsqxZvHD/uKxZ6QHIqdvyRkLP9++x+krPfdTjo/fvsRZ2YVXKanh0P
RPJla08yDiXPOQX9RnwSAUZfi/o3joIkfD6hyegWL6kh+femA4mhOwhAIEqc
2lWHh8xHEJXmc6indpKU8KGN14kjniOKu3/rUbHarNoUQd9SU/cCJ6FFg9AY
0n8EBHFMqd1vKErpgYYGNDePyMUOMBZDku5xl2U83JuTI64YibA2xSTekexr
d6xOKuwNOyFxvH5haSj9viwMlh7bSoo+o79FK63WgRc1n4oJkJp857lb8PM9
HaDG8+dHOWnfAblv9mLaJXBHJ1rG9MZaDRcInB1BLXuk47qhapGUrwUiNCFm
bmWb9VQR+WxpeePBXTsXw+dIr+CT8xWHNR8vx5AefraRkaKKjEQcNz1tNIDD
bEj+zu7pqAJvxURNMpXF0D2wW/rAm71EVC3cXQoIN4aWVoInE6A4CVd1UrWG
2flcVCzgcQ6KdLd9v2Qy2t8Obf98uPDPsNKfQHplxMdPBogbJ0BuifogcgiI
tR4IdPtqjeZUu6KpPHUp1OPtu3XEnFFe/qvGv4rlyyS1fuFJsNLwTQeAgSH9
Kqxm+xmazkaI5WsitB9SN9OyTQRgkPtp/x4cM7f5c2VZPQSlsjPAEWQgzcqC
BQuCS5KTsMux2KYqEOJMyAYLBz0YO5suW5OPrOfv/fmir5ZvUhH7ma3QQYr9
28Vb2qPEF6ldtRZik8q2QNVN2ioQxfo16pMirTPZqG68ibvwGDv54j6u/1mw
+/xisHQXlRgCmRB3wIpby7UaE/mP7fy7X8mXu2nNc4zHPE+FDyvTBfgR/jzv
53vQ5ghXqCjWj+6uyjloMW5xp2OiKP77v67QrmNOktl1at478+dHQJnouShV
Tn5Cq7khR9lTgWWvLe7tVUxrCURzxWKenbW/BWW3AnvmuWgpzjFwGGvs0MFW
oiw1OBaiV4nG8hV3FVJHLsYxGrggw5rCH2X309tsMnlRwcZZPuOMaXmRqVNe
RlQCkKwtDi/7iuv2DSIEzcONb8AD8UvgsjMNB6msyCP6jx+oLV7HdrRRJyL1
kBr796kKzMIuHHpqTF7nbkjoiXi0DOB//ek/Mp/nVbrEqX8B+5GcURBV/h6d
uZMtzkpdaCkQPiRwVPeKRjx8miZZlmDysmYDs0MSV59juJiBAIk//0SCfrQ8
9iYPDOgbwvLJ2LL6aiJUyIuI8pNyX7tvJ9Gi3CqtTRyn9hNVhcrn3vLQpSk5
fIIXLjjplieAK3cpMem2HBH8NhjLEaAP0HO/Viukd8uoyOaVFBK4WnJhHD1N
mIWwbNR2+1ZcK3UuLMY32T5KvESRlAsU83NI8BpOKnDLRbvXHc7BFnQbVO7Q
7ZS+ll5hTnLhlVzFnZ9MYVaM+/kusvOkrHnHMsu+8tpva8pCtwH2ZUguSFdz
ok0Cz8ZLfSwgInf4Wfco9nV7yG9lNHeqEHC2jsN/1NdopLoLXSd5Gi7WpoMU
TkaEuT39HlgKwtHC2YY4uEq+P6uBMiEo3f5MCHTBb4AabsTGP3CzJ6lpoCK+
duBjJ8/f/mqSZ0e4V+tkO7wkBjOFRl0P3GT0LkEjVj/zljTxzNKs1QmYmhy4
/1e9rwNdDavYtYSAYALB/YHy16r48saBoZzAn+pAcWhacJYyQSysM1BewXf0
5+6Nm9Tc5aD5YyS6BmoqOeLxJjd2iLa2YRwvNRVFdheFp+J/G+Z+LkcOUvCA
nkiy2lfg5XJzRkheVOEPptta8HiNiSeKn5d9ta0R1L2ragRlW1mtbc0UiwUm
5ycfwRyA8imTOWPEUYMgj9Jpd5Z3fIXGcBx4Me6odG5sdcIpghEuuaLokQnS
atD7G83536gnByWvdhEeEQS6PwU5di46zGgxcZ3XwSo+ttdJ7pJ1GSG0FTUn
ApGxn1FtLUctlIxmSp/iJr7rcburMiKVdZQLtreSicR3KUiF52I8cB7mLjx7
1fmPh3RsbqNl98hACvxRaIDp8wCwOUVXxyuMOH6SnKW5XViY3nMfYi4Pr19D
Bk8YFpzCIwAXpuL/NNYufDiWhZPumXFubdWAMug3gg6LnO8bqY5i/mHsG36D
dzUxhu8YaGpbjHUZVRTq0HO6Jdv9GdaG9K3MTIEVogVmt22MZj3DL/g/HNcr
vVDZ6Fk/K5N4ltP3vvEfxD0TVnaKGLuKAnysQo01bmvaErdZswxZtYhZKTY9
+HNTKU0wUh5K+GwYTPCydVXdPUeT916XsiVZtlCaKwO0Dg1GfIWnBzf/jmur
CYnM8303SHdgY1f99v3Ax0GBL6c4zBzBic9fqYIKXz2qBCpCEuCpyMQ8oN4x
eEsE/Onqk/XLIL1NY+7KAMeqPWGsmcWsB04GTbgP/ZxeqBV3Busqiwbq4VdN
mDTsoYgaoJgO4mgqq5AlNEnxzJ6VeN0x6FlN6NQipaSb2PkadEnpB3oG2U00
d2ooPJ4KoJm3aBad2NbH5lVG9sXeInYd8rZdMHdQuo26y/7a+Wtw0eGfROr9
IcHxSAEhQCLHLFAscLBI/Wx+3BKIGZcpmFYCOiq40BrIOW0vWJdN0YrO5UEe
Yi0cHNTbvR0rsiMVl4M70SuqOKyD4iQGd5Pl0juRL6K/GPES5aubACMTEDgY
FD1Nr1+nCu+d/hz0j4dvYWftfBZtRXXOS1rcVADpTKxCuxTSaXOvfwvGuScB
paZCtfrucdKmAoBJ5r7aIESY+Uul+ZCUrPkYL8zYnKedb7u4UYuHosEKdjYK
LcrP87So3w/L9GJ8ma4vzRG5AwvwHAlkveOH/hJqAGfayhZ+eUWwbPWQq8hd
h4iLyy72I2mInUav4nU1RHSVsv9vstE6iU+QYO0S4/EIUcXV2R7e4nP8TE+Z
wbpEaph9ZVb15Y/49Gp3XgHABv6R4Za2HBHsFDlFf//QibqBzUSnFErmzPGp
4MNlEdUPSfs6piij2vTCGxTkFM2w6HCDMbbFuC2+Z4qqCK13rLIyX5Ew25zk
nsbpBBYDCehOobeV1n+B/xwZDzq+MUOjzgj4xbbmSj5j/1lxfSx4HYNIBq+T
oFEo/bH8VSAa+FHeX3/uFWN1f6bv7sHVhaZzLSQcnDLFa4uAk8c3OV5rWuK7
6a+Sw5/L0xp/h2B7RCGHNf+SgUGglRIu9gy3FtFB+Uyq7+50GwMS3kjjXD8r
7YJatpOm8nj3f5Defk+ofkD4GAtyS+XxXiSFt+eKlce2TL5tPIV53ex+arhG
lGqdEQdiObycgfFySWOamAg8SDFcx6iFXY52dZDPUm+JDbWnBqB0e3Moy7so
EB8Dpu1VupdN9dtjp/rMTp9LJXQQiz8WOjPS8l81203aY2WW7xgqY9nC6HG6
Ru1kv7kD8UInvAA33HZT30mwwFCihk8dt3Cd88XN3jLodAva8JYpJEmIy0zv
TlXjx5xs5MGynciNRxNN7lbooej1i6otZz7jZqPKOvCk3+9+mvClKi7uRhQE
FNUBlSXFfQUmA2tY3W6qOlQG5oeG4d144e2uokdNpDoXhxmflHLOHvv748YL
dHN6fgMXa1LfWIapg2KjzZSZjIxQolIvWBalGOFZiqeMkZHBivGYL91EFOLX
clJMBrcg+l+ZyMqLU7DKwjFWFs8KCioDgqkTdWpHCgwf2wSHNoDPNwG5p6Nb
/27PNatD6ldEBSkAjydgS025HRbyw0TevB7KPqRK9kCajQtRK9kW0rJoqLi7
COV8XbV0G1CxRhePau4guLnduOgjEhDSk90xg2ppR2X6LeiMiT4Rk25wOmGd
9sUlKIyH+GXNh70Fx7l4BfBdTU7afklnXC0NOfDM66byNy62CGz19vcaUmAh
E3lkEZE7ILdKx3MPYlPUAur5NS67at6BdY+tAHOZyn+T8lywwj1vVRyD7xMs
ua8pXkLGiQS1ZiGHh3dwUDJVNZenU3HueE1qWK4iz1ZOrsUT/e31LaJrCf9I
FYqMiavkiSOh6hEdz5Szfh+6lSkLFtvTIpoaPdljteD3xvnE0dZzXfM0mw7Z
aJmzHaJj1ajcax2NXxfk4EXtTXFdieeTM39szHPDzt4EQsujkq+EvfeFnrgF
Z6s7berVF7wJZpc4OTspXq8M0gvzSDiNBxYZZaUKARSRpKFW+POmW9yDPpxm
C2CXgxm//7mpDYtwegucLizYEnDnXfuznmZ1uZPzbZ0LxKFylW9sMarjOJQu
hDDTZCx97H2G6rTDKViIQEZWQJdKXrinpHad46uO5o0rlCdz+K3usRaPfzCD
xtf1QTt8vxlWcoLovaKeLGXjuOz2Z6SRddojQHxh0UTKK+8G/pWgbjSvvRUc
ocZuFADFQUIM6vkzQ5pXGBcT2jl7Ct2rMowpst4/5TnPjmxrFo+xH530hcL/
zANMdzs2iCUPh7lT+sOGxAw95EGIX2h4/WWInH6KRq5qQH1xzPyky64H2bhI
KhWlgiDO7ujuurZk4V8uIBiZ5hnaYXsY+5UWKf2S3WJ6FRHFDAbG+e2oVzBq
Vc9zcqoQvmyXNbzW2EIB7BCDoN/eLap6yLZF9WGVqPpRGDwzSWKyGTRtSQmA
CBl22JE+yxocKye2dqoGE1ma49+uUu6WSsCTRcV5hoQD4G05/n27lcavi+bw
nHDxl2TDslCGD/+qxirU5HLxlKLhAQa3gZFqmJ/etbCWFJAXLFp4KWXfkaef
ypcCzdy/tgBcKh+LQ0tG4N3gGz1hlQuD7CvYS6AvUCkycUs+DDIugbvVVIPT
0ZBirb6VXh8U0uvq4Q8jtkKs0QOG0aITDoNCHCUqHJCf28U9jT8Ig6TXH6O5
LIBwS6s4aHv2E8HnQvHvpV0JDPji+U7juRZiMp8glRH6jVEWVKw2hNXF0XOD
nPpCXWLFQHsfAZ//k0R1nbjXKLcN3k/lqVcg0WtYcmvsvJ3SNM5puiPT11gW
WQXJNyX7Uz4Jg3ok95tN6aLxJC7PojCp2DIG3LDCA3JgJE2ZzwlDXAa4MbzA
WH76XG5WfyGWX0Bd6B/hXgtaa0ATi8owsKH1X+uO2a7Do/jhKUg+H1HBZ2Nh
qBdXnGRHXZqSEd6PDujiBSo2i2HAxRmDhHU3OARqTBAKWviIGOy4s1+NMXdK
hmAJEPmvDWDTRlhwOo9ZkYTGFL72oiscaj3o9Ioj7jY0b+VoR0g0SK9Bwbd/
AIH/vx/Wyj12KkAu1S9OH/AxkYTlMldfPm0+bFqqQoy8tJuFOQnACiIL3kEq
/NSjmi1sDhyUz/+TOdwallNNHByiCIM4rHquT1PrcPHvUZEcMyAT9iTVg1Ja
NscjPznvPNtbApjbaiR3TFMMv3Sk9H5n6nbe2FrRNGUCFis8JcUpZ0K98/uv
Zs0Iax5fwbGUVwKTP8MGoMaYIdz7JFkbzvoGhn1SKwsAa3wLsYMEPIvNXAYl
xlo4h4yYV6xVucj+6uPOaP0/pZFrBfVHabmTr6044cp3dBrUYL5F75yD00PF
5is4crOuhpr8ptW2b+Rj0e//BjpkYVkPnx0D6YiP3KGnWaxaeBKzGQTkhCqP
zSklSCGpQ8a2o+Ik/DeOLkOiQZqdKJifYP+/lokgtWMMGo2f1ZQnToHhApC6
y5yS3sMfMfS60llb8fx2O8Vcacylz5nZzegRyozTJG5RhNRn3f19ZIUV9Yoi
429pH01jBkojBSplKDhPS0XIf/IvI/FqB2TpS1CTrJ+ydlLHIuYffK2+/Q/3
uATbdp9Bcr5LjW68yRYZ74pzHGPMGG9ETBBA158L9MBx956EvokLqgMTEtC9
i83kqaYl5KGSpjwl1JBbwMxlx3eF3LKA+MLoIoEDbd9OJ7yr1UoZ6sYXAxb1
C6wuzC8u3n8YnVDT3ViOVI95Eh1zHcnvpEaoN4+/9cHsDXL3jHyKgq5l8en4
dLBKo14DAWkFnOOyWJYhRNSl6nvN0aEv6u/j4Zclqsxxzh1X53ZZ9tpHo/K7
cVeqk4wDWsh1Wip+G6CfGnkH6kDULIPSMct2g80JnoN0A/DaWisxph+fpPhp
0hgQmfVADJddB/U4SI/qphCEj6LZaYaMt6CE9dN4UMOCMWcX7TD7pPmXAhYg
IStm6UScoTKHAU8FP100j+NXVYUVrYD89jfTi1OYHxz7QEWMjO08Wb+f02Pt
jDW6qdjQk+4olAOziG3oEjlMh6OBsfBDAAmIKJ0j/iqjnoSDYgGrDDiabV8g
Z+I915Q6AzFdMyCsWQhDEhGGTkTSpFlA020lOtCUVhWCDYJOsVbA9gEUPPL2
UQbEh2VT2HAsdCbkjdkSelJIjMw+R5zziL4bEOqzzVCqI1JXLVqilB74gWTD
N0ZmB3b2CcHDVuXmpmJ3jn4HMrwHC/ad6a6FKPR3fvPXg69xisKe1DbqHiE9
LEFa1deKYW3ZzlELwV7Oz7A3zNd/wUI60DVpAEODeTOAkOg1bRoHm9iMLBJN
/xdQ0mrS74/sF9rxljFR3odlUETgSz6nbRkuksWxIC2w3CTLnczqgmxATuKQ
SAX2qytzbQJaRdrZVRgyx6oqIgj7F/KcjFIY2+Y90APJ2W9ZqrK7vFbtnzEv
pLdxJVZXmozkHiVn9QkUMDK5AobLXVrJnRgG/3hdEGzRK8gD018/2sE6UDjs
XFRc3zjIkzYDwYEzv/CPqMjV5hooQKVEV8npTc9GT2KSQ90nk9xmFjsRcwgg
PDRYVLxXS3CpXU39F1VBNp1gv9pDZWLvezD9Kryr401QfWFqx9sypNam8aO7
u8nzclJ8xCKAF50Cr9CRQ1bQDQFbYwq9VooelkIG3IiijK/UvDJ6wGXIHlt8
bZZUv6sIeatLX3rgcQ4NfDrN6OCiOFXw5VsuPms0k/xj1V9igAFNdSxd6ZV+
mSFaWCsp5pgklsq2trGCsJ53wg9hNMU7ssOmtkE4oU9LBtkOR/ulV11JxZ3l
wyYYN1YfVho2hMTeMHdqzRS/TtvZQnobdDfFBljwRzhFS/t9ztTuh2dd6sCk
zpvlqyDSDRbP/24DTFX6fI3r5hhT/9pgIYGkODTurhsb9ohI62RjFC84DRnm
6nBpyYIHrq1Lrjg/HsCFOg1Y3iGjo/wRbo3KtzthfP2DxOGgHRCLq4ToX1/H
KtusVRwot08MgMaRAT4k4DhzLxodibA00ndv5RaJp0g7WSlnBozVuklabkvt
nlSFjrxwO7COgti3UP1LFOycfFSNOxlxs1RNmPiejwGbVCd/NrD+/twWVdQd
ljtY6hDBGOiJ+x/wRueOWz2sYGANl4d3+sC58PBfOJsct9schIUg3CQyf3Ty
N/5QCEma65Wkr0ZIK8G/L4J1nANlqI4PIsWhP0Yb5jhDSzTLSoXZ+kbJqX7N
tlQ4hZMU7eDfKluGqwZh//iFXvGQHniNgjO6doracWhMwyZ7/tk5FCI6wjjo
TDw7SmNpETk1I25veCbku2mK/pSIrRoDcPuXmLIT3MZC34I7M1TO6qkP43xk
3BNpYr1xM+o3KuRIvosJfEKkj5g4aA49rRbAM+WIAKPsF50kENQvmwMTYMHS
hkfDaYkj3OSVuxwyzAe8cotU+H5sB+AP+ZH0jf/STdt70sItf3m6txv+SAcN
PeRn6hL6KR67E16LkqPLVOvt3qHKuT5PzeNwqDnSZVKLyKssIPA6htNXTPM1
AEokN9O/6Flq+r0tQJlTBgsa7WIgN+dyWsm0LBm4jgPctr09MnoB+ocUJ3B/
8cQo/KPmHcshybrHroNpFa5Vmt4i3i5y9WrsRb+01IpUr16axqW1F7vfkX8X
z8poViCkUjFrRIEwPW49e9jIorO9BmtZ9cbtiehHmXo9Wuz+EJqKDuoReicT
d7bKEScV5Adun6SNCTN6N022HAojgakTOr3hHhNH705O1HhIpMH7lwBBY/tH
t2DaHKUm2NInVxxXlG2M/9fsK0+aA2kGyBjK0sQe03PhFoEwyr1KNKjJYfId
DBDw+QBcMFmHOPQdLreWfwLGYLi4kXC1HnDWi9cLp1Pwxon5/bpPJRplsZm5
5YshtI5tJMtSD0nvza3phP7w/ul8KbiRzRejieeaj5AmmbDLhpDttDeSEVY9
+rSpjczWb/SzgmsZkK/gvZ78BHjYHoLZ6V7epAKbxcYPLZgBjeekW+oos5ED
f3qoVfeKPjnp0n6jk2pfTHlbKgv73Nar95ytBZGV7oK1d0PdIO6wO59RcrKR
b1bkrPK+AJiiBAItphup/JVrzTpSYuf+rNYXsWJBo15HAE6Bte2lnOUYv5kD
ffzpIn0r2bu94As8XuxxAn8msr+nEMTFBuPaMTPbsCsWj7ihOMlXJmJaQS35
TBnJiINCZ6hHakh9mLErdBWeins896+XWhMlS5v+TltagzZqQcy7pwha43qR
C81nLiORo1Z6gnu2L6ZLNWnU87Ra53uqxf70rpme6TRCzENXEjSkbSDmVL79
FTpviykBP8dNrsXWRFObO6F+IVwCqh+ANuxEF4v91Jdo1Zak2gmqvj5Hb0h1
DgMxJgkLpLHoC3GqBYIIvJyD6J266DXwJnPec/joXHMRqcUe/asKH1dv92ms
jcDKSHRIOm0irLqF05TBGYtXDjVX0qVgEd9gbyLXV56dDzpZBlqmhHXgYDh2
uhfjWy/UT0569E0uiBYSUZMG6tDqLrXGwDiyoXHmhsexEfh+JfZ/7nnS0AbN
AJsgZjPerIxM29TM4F51FsBhsLgfmLZYvKnEZCf9btmOGGerdy8Ni0dnwdYt
MOqDdlcbV2pW79DP3LAbXjKy5gFFrkhmpxlZ2pks2WkumI7diSwz2XqEbB7o
FD+ievn+QGUj2tAkXki6+dzPbkjMIVTDjEPZVc8yqq/Oyht5sGJB8jQ2sz67
nCUMSNCsOknR/lk2S2UfyoU9mgRfndjoZ/m+agcdyGBcm+PKI0GMgKfi0zvV
28lJyHyASAxMGK7xXmjrY7gvFfhsWRmMFs5dSL+YeKb7dMqa+aLTxkqzT60q
qzI2alDb1lMqBprr+V43aQy2cR/D9FBOme08BUtjqMbWEUcAnqOisNvb0ANF
FtyTsHBvR3d0bjjTfb45y4vmEt3AJRpo70SaELA5RZno6vMSvHiLnmmOZzGO
p3BwcafwlscLxpGHmONAsGQ0wy48S8RqoiHMQZy43bM+Qb3V/Jl3ICVdGxn4
PuLD9Tyi0gTs7Xbuo8tYF29Nf+E2br/M0aIQzbUAgIC81BMQV+5sIIzac4wE
M6yeRo0IlOz6xxFobLkW6keebweouVzGMvtN/yP0CbxQX/aKKGAjdIdeLvWM
P3b8bOA9XFIJp8zN/rrgaBDfngiGFe680fJl74iS2/cDYRbnWvOY8O4DCm+y
6SDHbYqOGmxHOxhRHCiAcbYN2zluP7tNMxtWuStKTub4KxpMqsMEDT3Uk/TZ
MFDRYXU2dpbtjiRPS24Nub0VW08t0nv+K3BleABJE/to8ENJ6jvgkzko2i64
Gm7tnXay+B4yuq95cWcHl5Ipmwk7a5rxz4bfU9q1LwdnvNMuk4CK2C5cJ+xV
hyzQZZp2WsL8RiyuxIrhYXKx/0WBTmjGHw6lXg4ftsQIOb4d7LLW91Mq1nBc
jMb04B6MzR/Li5zU+xqOp4IVJ0X6sQ3e970UUL4yEr3OXWoYRqWhA4kDoFhk
lqZREOJl1lWQbM9mwMwuy57wh8neD/kflFfDvKrpuFSH2v6d/QVmnKL9d65S
BoUJYVizdb9kNFrvG5nCyZmUx15GBA72YwwU4HErkTyTsAVWYmw9Jj80pvzA
UTuG8T0CNlLgFdoI38BMpZORE+P169ma2c4tscWWFuVWUrtjFzar09qkbero
FyAfIjN6soNDg6x3gwMUW0oYYxmdfbUbLLvKprbyGiR3I2o1Ve92UBwdwEB/
jWXxYEfpQ4Q1fPxZ052CpMc5eHwkolSYTk5BzD8BhbulhaLmbPYO6kUW0d+f
+Xh0E8sF5dx1Kptw2K3M5lG2mtdVvFoaBfXlwF5bJGqasxt1k7jtZfKo5/eF
238bH6j77/5bj41+K9ND8pzo0cj17Unyk69ara3PhxTCP3KK51EF6Mn53WGt
IWcaRiX7NU04iotiwfkqtGDULX4Azl8SPb2QFKEu9YpDwlws4/IaFsFcfqJR
cEiu9/xIsRL9KGBxPhbTsRHxKVJpfiefih0qce9rFBckonXoKlkGt9sBjnoQ
s/ofslK1P7CC7z/kQ4+bZeHnLZkPqbRcnj2ER2JgbBR9yD/L5SqUDp1xyMSp
lliFGbVy0V4psS+qkpnKzrGAogB7HYL1cYnis5zhqY1UHlvPq3DrmlkZAxdM
w8cRYoZCa4x5IQ155ui4/zNz6sTcfpSyXspP/CO9PJCJe0L8Y3pu5xPJARAI
F2PVR4Mymh/8x2srqH9Ghb4oVc5ALbwyPDuc3f5d+C7xI/zJlQEA5txHGlVh
cy92deRDOWZ/JrP0PXTfxcn0TMlWkBGgR1nbXboVvHZuh3q7asnYeh+gYi0R
kLeA8KaSyvzS99Lrock5eXof6Af/Y64ThLHG8c1rXI0Lv8Q0RPLOpUXoZDDC
xFaVVu6NL93quu0KC3WCFpKGRMh0+ZBP0EM0To7PR6iNyC7Yt3EFM2qVWP/0
bTOP0uW0N/fUncsK4wyls2z4ahSdAup+wLEN7Vlxw5ZvOSbRdbds99hoZarq
yJYoBqzyBbw8aoa1VCsG63oNeyfFR6ruyrKyyMQXjRb31N1nvZu1AAk3u/U/
fNc/vLJ8MyoS49FoK1DXBRR3/PpXHCuW54bdGbAPhtulR0C90kaN3x1zXfOq
1Mr7IrPl6ZbfHPL0XxdljJgLHqtFNu0L75xP8KK+TW94EV9d7uPPreEfOu7e
l/HID/C/dabxk29SoMWHDhCW+Q7Fz82Eadq8yxGlqHDM0HctCSAtB1LkAfIB
XDBXvL2StshOi3eTLFRweuUhye5/5e3YzoVRh3scmT92PV8MrDmAUUP8GmPG
I1XrgskpPEMOixpybvrRQoyeVtv3sESyXhzSZzYV01VMhdjruj9xrx3LiJrv
7fwVvqiRQR0BZcH+JAa2X+gP4EV4hXLd5/VngXevIPR02cpJAzE5H//txRLX
HPMa+0GOEv9BBbfcEmSqh0abn4DuboqpD1Dpz/H8nJ5hUIN8g6H9qD1STbPr
DDgPmP5fMIMClNU4JPcap3SuLxX44uWcO4drlBQayl8HjCCvHWXnR+wMHP+P
lXwBoMqNXMhP0pISJEUBPWREALC5aEotKPYq5lg/P+l1kOjPpA53uh1uwzSv
NfOw7SzGdqDP4J4IW90gV6wylYYBbHvcMI8yPAyA3Z1xAHUrD2HiSNbCQHs+
SmwtvLaZNIRaeyfsZm/UHJkETyKrxiE1ZYawvEUJpFwA7u4yreSiEuUFnky+
Wlq8bbzFTuxfnDi0/qUI2swLXKUb8EJo5DrZknph3tV0A8x2oLkYpArnSrc8
lcqY4o3yb2higQzhx5DreP8GCVl5tOQA8l2/E61TO1clOV5ugQQ3vNGbKRRr
WdUSNakAa1u7Wx0xBmVaShfOFAImbEOj/pLdfsxVwQkXRHErr2d0DuubkxnL
reWfTGssQblL8BxZdl6ab3H1UFSIHz5XD7WGkdVOOUEjGRe47X8xYaJ+N19H
O7nXBeEsVAFa15XhLsjyfd320u91GG9+kv7AxO3sYKoXsQp3UdMEYMQuVEOw
vYDQNYxBZ4ktEHaoOZA/sbENTPDWudtuIzpFGQre2L47PIUVXTZGApq7YwId
eaCqXbuTTSqGkobyjlUt0RnbVQ+bAGQwWH1igwDbQWyG7WBDYC64or92zayA
GToVZEn+Nk4rCiAHocCYkHhO6QrvWxn+I1Zzvp6I76Q+v7Sr9+aul50LfWpp
/zHRBh73EefOq4bsOLGriMACNBw8+cMsJoRkM/WguFJCaxk7i/Dtrx5bBuWv
a5ExM3+R4BDvLWKx/9QiQPPXRC+NXSGl7pLpD8nRLPbokZkHqNRsCcMxV6Nb
UCmhqI9aJdkcUzlMa4PyTy/9JXEgLjmCrqHQ30Q9tGWqJ/ccOArzH/wuXQDJ
H+zhxZ1oYlsqpALiUyVOFsK0Bo4nnLdsSwm7U4fMDDxchEkKBpseOZp4vDpJ
smWv26CbV8hu0gddGNjvJCPN1sPPdbtptlMh8cQmbVwUDQ/T4m8/RU/ZfKqw
b8p7cmU6LqidKaGSYmQVjfSWp/W5QQt7RgSPLq0bodIU+ETuVdT9m0x8p9V2
WeHHntypTMfdxfuQXs+ZCrsJdKN/jopOz/AgQi9CaUHUFajBySoyPI9ak1mp
gDKfFNXAIAFIBSCcAGrt7wLIsXC5tk1/Ecfa73tcnEwxY8RfR4aFVU0k1eQi
g544g4Uor1tBgoySO7uh9Ee2+iVwZekfFUqADWIzFgcs6wjCNOpo6+M1K/la
uhT71lrSeIA+pao+8e/PakNAYBS6cplep/Y9YZqkBfuVYRYH53co89iKv+kY
Pcw/n84ZN2qt30mYkZTP6b3VKDDn+1sRJHlTtFeYM9HebObS2fffeOAbaFnA
xsJMHS8HhMWnaC7yu+jbPsZ+67P9PNdCPFOOeqViigN8mf71MlVuBbmfpRME
O0HX+myAQdL4OInc6vfwNcTY5nnOpoxBIVD1Ebwt+lciooaO6LNHj0/xZDNx
EUjVRDN9fPECpHPFoqZVYE+8GZvCm3s2GEUeK8T0XSk6FOAlRxACep7wAVW9
PccgJjiEVnyuL58wdfGZn2RJ4Ok6YepAd0+C2tyycByuCz0V5SU967z1sAin
ZeUmhiwH/JiUTN6bTsYe4LFle+Ue/Ly2X/jWdDVFJ+NegQLadQ5JjmNXgHkj
qFsr5VG4ZpBVIlHtfzFwBWOTPwXyNS1jkIPydyBLnRuTSXOOTyUCEC0ZH9CZ
pjrmCuwb+jflQBGXB7TxIXctp4YQsrunfA5r5dLHcQnTrvfDJkuvCC0vfMo0
qK1RT7rTBFoNIcrFdjFaU3bPMj5TkBlXJsZSuWux5eJE+LRdrqvT0TXXfand
urjZhXm1L6tATBQ40hUHRxYNyq3r/PQzQCA0uOtLsXHrmau9jz5CP9wCsNNX
Dd6tS/JuNXkDRLdDmtRnNm8qRmApNvSvuh1lF72iCXbuk0EBi4NHjF3XtRmy
pGAblpnkGImWGmn0ytplIsATAqowXgjN5TgQC5d69YiiU5g6uXEComH3GQG4
rmKJNA4LE8CYFR82GvpT2js/Gc/D6sstB1bJ3ms57v8DQFhMhFgjc9OYAvjk
SRiAoz9p/MmYe8lQComoJ5DzYLvV+U4MH8XIXuMtB+ov7gOBPzW/Nc1MgbTL
b6FdfdeVgkiDW1mVyatoz68EN+CNJeRvCBW663bJFq1fPA57T/EpYZsQRwPh
kgMkOFYeGnkShT8BY/7Yl7gzTLVuxGRqBH/hLkn7lowg3O2NH9wNf54j1Cd1
ySrd5M4yhA3kQ0HYbLE/Yg51Pvy8mIMtgWuihSWAHlLUxTM3iAUzkUY6mG4T
uS3TgdHKLYv4fXcBQzqmkGGzlfZouVSy0wgY0r/dWAiIVEPZoJANvPpbwhFH
roRMdjL4sGcUOYkGD3mwARdyvKNeoLwgo1ySRTwLDW5F+KH+4BRBSzDb0z/t
1OgYMr5y+kb7Osf8PGH1ID9rY+le3fkhxj3QWIxQY4T73ey5LRRk6d6QHW5s
z2inkMHAIQzaQwHPxFNMyv9eIMFDTrsuKmP1FMPgCCgFoqOval4mC3EuEsIO
+tW71MDNirv3wCkaGvCr55iPa8csO5zWER5sw67765RqMAjXnWiTROTls9hi
I0HFOIPTUZLPBfH99PzBDhlOy6SYLlMdjuafTeOnC1eqCEIrWzqFgzbYNWLB
QGorM3stDnuylouYrKnl4KbtO9IKpfyD7dVgFxxzLCXEtGx/lgPkuywYNfQC
/gMRU5tOH4Vj5PxC7jz66ZNr8iQ1mwFg2Se9Q7qioY0/XvFmY1cg0oDIxgMC
pbt4y3hQikfVcUh8ofgp4jxgt0j9Sgyfr3eZMHxwpZRY8N7+xBYSQV8FFFrv
9U9oJb11xEy/9WUuOoidFQtDTrJxpMzVC/+WKBCmSWKI224k1qC2DZnK2HVp
L8KRElGh9M2uyJFabcWtpgQRk0Kh+SiEp8RXV6rgjrRh8qCJMpd5dBN5Nh0Z
ZDLPF1GEzBftGeHYLSEGzn8leO0KDPYn/IvcWiwaHhmBN9Q4S1DaFOkSx08a
jDvmsAzrSuS+bdlKMuijNVr2hw9bYADHy5bojqWC1CHhODHW9h1ZJKMvbM3x
ab+qlDqNeL8fUYQ16isJbTx8ExHxgflBNyeMo/GCfCC6usFa3cm3iGJQFZM7
TvPPV8nhNP55lVeIfgUfV7VIIJH7NcKC0UhSJov9tpa7AN46+VVNgCWlJvCH
wLxLohIEXnDHvry4x5mIAilFhxUbD2OHPVNHzN8wd78Op1WWmRDUmTeY3jY8
mY0bksJAOBlzym9EVH/yHGVtFAoFEog49LERfR73oyxALM31hPGqo4WAbuOi
VDkYB36an8N3mPusMhOJ8PzyzxxoQ0yw1nr6X7MJlzh8iULZjhHXxAEUNiGQ
ydZG0Q+DbW8AWAZOaiDwrRfBVyjFVM/tQp4CPGyxHn8CdiLCnfRkpKucK7Na
coSfNVE+EeEUM6SF6/Q9eQpQCBAWX+LJRQ3jWpvjsOv1Luyw30vht/F7hfx1
KWJDYxE/vYhi7V6IMW0ZJmv9oyzoT8U4nrVtGcS5VhO/4THRyTh51Wy8Sy0Q
Ofk37pe0taG4HMulIcMMKx7u92Es8n/+7c1Kf0+j7QUY6lQabh+xSEoDZLRJ
33O9Qhs2yvQ1Ki/u4dME3TWbvrbMjAyZ4xtbheJfnvpmXVSTINFXWMbO/gmM
OR6Oo1R0qxDyboYmuhXDTSAQnkZVNOsxqyLXzoKu+X2UsVwgMlFLDEqUIour
JKHTvMynQl9/eNYKn1D31klwwF9Q8/bRZSGdBY5WwNG1TsNGtgw+KvtUkVWo
xX/50azDh42gDa8EPbTF/Qmu1cwjueYF/P+DLk1dP1I0S8fZTbLRkxOn1Keu
siPPtS8mIY2nfiD8TyqdXHwRb3q2aQc6M68CJ4OcT7gNnICmxqD31YovvLw4
fZO0mItT8jRZFBSz/hLBIhRSvAv25ufH/mGxIeCXBu69LpA+CvHrIQyxGsPY
xGGOa1V7IO+8xzb03OEmzIOxIHisMy5wk0TwJr7694gCBMiCy/dBDJai5xlu
JXnOmgYYAcUEJIWywEAP6spS8I7e/URgS32kBjtrbCQvO0dTnzabVC+OSGPG
7mvHMOSVNbd0ff/V+d7UUYz9/xsOjpzJ6Tf6/nd48cnYjiJdf5Bjm8uYxgnR
Rc6rn3CWvPIbSK4o9q6TEEmKsI2ScJXRAP1u1jIhqntNam3og7iKGzmN7R3b
TEAe/zworXUCgQvBRfppK9yT6T76ZP/SFhxfYG8/9iSNUPED2/J+YtKM8Z14
nHzipQoXm7WQLvLCPzTZRfP8U/sidyQjXYcAALD2bUF1bCkHrSwS2+LWCjwT
fJl682JU0gYTHx8xbWiB4sc8Z4U8EiPKFELFI3SlkD5QgMAr6hB1ObG4vYuj
WG+1tBFDRUvX6k2MqDc3o7BZQuL0go1ILpHWMN2CVxCY1dfjn5zrHavYW9xs
LGbItA3kl108l9tzbwXkxcGX8HxEonwHefrn/CsXeeXgIViu09zae6oHNZ3T
+pDmp4USpZe/JEQK4f8NYpdjpkk0NFgtZONQlAqRUIsA8D37wgltgiw/lysW
3i5VF1NrKvxAoobWBVfEkIYW40cpRDbDO958Td+Aw9C8MzsAaoQk8UoLocjZ
sP9u4UVUo+r9uyNKMtXXVxKblJsgxaEfA0DnLhXvJUPpv5D8Mw/60QGwFuaU
DaBx+10andZnJbU7Q2BAkcYfwGU9gpCKRCRozMIL74+I3x/zPt6D3mSHAdN1
ZwAfseOdwIJftXzK+cWHJwrcaGBcw26rXBqyCZ5/Q4+UIlq9Ch+5YH0LxHe2
u3ODoFbZ7FWQUnhKEsBjZvKqTTR9URjwZaVyA+ukqM5i/nGWbdaE5g7pytSL
2RSChn94x+/SK0glvFdMvRyUCiJ0/0gLuL6yfKEcVPClKzXctwbNCyYXWe0e
NkyZZn7b9jB6ps9914dNK/gLAJys8k8BRqxdlEhbGEhlo2N12tWDAdPTQEmZ
XMJ54rh1jpxR7Z8Rg95GnW0zzsegMw1VwopSblH3GIfwJ0+e+smP6L0Xu66x
kQwPvBlnOekq5+UdPBNFKUB5VnE76Da+3R8WJo54rdgbFF4mPmraQGmq88ZI
F8sGZhcwao3smpYhE7em82fyWbh4lCvvMpst4/diJP8yPZa+vHCqqTAoPxnT
OpYME6un4A1GRgZdZOV1EzyqWPpgeIezYgPwvD4EH2L5jHk67bUl7Q/5E9z7
QX1CakvhVxNyP7VM/FUEmjxW2mh7ta8NPfwrvXeOUgtb1YAIySeQULWD03qn
amx1vKCrvOVFY12piLLBh8qS7nx990lQOIid+Svj+AEBB8y6/k+w5qAiVLa3
fdnmUneVaKykiZX6LgZTDW4gyyP5ZESFdIpG9Dz0XntXunWoRz7A3pv/YiFN
ljaiq1qJsT/WLe1+i6fXC9jXf1v4NBO/CmgZMuh6ZOmCX5DUys6+t2qBajWp
ClAbRAsk7H/X4HH9qqh3r4VKRsJpeqI6vohSMlHItMs4HXDiT6peXHFkGtsS
b6H3kS2dXlX+P57X+oX9hF9BZZRzuabMvQo4GgNLQ5C6hpz7+YUAhWLjslLV
k5972jcQp5zFgPqvbaux2wMuQHWyMn+jWzDoktzY8e1pO5jL4cAAZ2wxnXyE
7SXyWLGwrFFKbQEbxrjBPGKtU94g4VwEJjuHCWfyXUp81FvdXTKWhr4YBCr9
rOmCTMQzsa6MBucbC8uoBQpBin0RKnqr1Ci6CaJs6ZZl+6gJZ1FLcmFrlGEE
5q5RRJlH1yC93DhAtpjPwQinEq2COAF4EUi8sh4TMwlSJAkGZcwgdJbNQ87T
gihwqOjFDeG/7SGTTR72NCUpBDQUPyIN1qxp3eesWbpbqU734YG9rfLnrhxs
Q7kKIT+ZAa0FCIJggiRsKpwDV4NEBb+lHSL8SFvqnfigp7jdbyqHFlQVn1cy
oIpklT5FoXF30nM66iPjGh/6MmqevHZwksnV4d2eotQZpIs3HuqwpQmaMjI2
+5qpgoBExuLFKpCeoq6+gX+QRVccwVvUDGDxL740tpNKeENmfTuZcz45KaZQ
7c93qAXKYeXiqkH2cRg3IFJV+DJgJpSTBQ08wX4LqqwofOgGwFt+PBmzr5WT
+gZGm4QKfH14+qdievDpQFi3EyaoJgSJxWn08uzOscEKHO3TQa62pXPe8gTv
7kZRY7s/WjrhgO7odW1z2wemgkbOzyL/Y9vEfa3w/UbEo1XOcKBmoeXCFkNC
lJ2VSUH42mQPRp96HBhLz8NG3SzQ5Op7s5Mpzc1biF9gRXWSA4w62pziO09z
zgXtfCJJ/SZxXXv9ncJQ2fCgOONCrQhRTNhAKQOYRYqgeImmRanI/FqhlxNm
Bo7mDLiDSjsSG2AyRIrM26Y/1/KEjNDOZRlVDo99SK5Jmb7+X0l2gY6TpURq
q8YFNaiT+aKfKG1VZYnYeskbgOiT+gzGSq0TLp32Gqdq8ghILCxxr3z5QCST
X2eONkUYIWVJvqeynp0t0UT/uluwK08w6JEK0hZ32aRg3IdWBypwcwtqAl+Z
mIumb/R5pgSnOZl+V42ZTErmmVd8BWTp3byr0IhFGByh0ww+wd4af1LTaRpN
OSjgVNkGbWdTF9lvY1sMR9bj6A5l4/EBc4WcLAfvvmDfN+HrqKqLFxWxp/Zy
WWFH7tBmQsOezzV6eIR49Z+AmadT2VYX7/Z5V9pX/HfWGz+ibbF6y36sZHVk
wbr4wB5heXZa6RGyc/IgqGh1+yzdV2I3eKuSX+z4D0i1MfYd6fBojsRPUWnv
9nHXOLQk7refTQ5sObX5vkUMXoxd7KrnH6vqueH0ExmX8Ofxd0/vJJUK93ZP
p+PgiMcyT62Uyr3gK1C50UwlNQlGyvlqeoWYoSv6OVYzX42uGld8KhN3W7BJ
gsa3QXyUKu2LgZ6gk0BhQRJjOEn+tOuROPsTBKZQJI/hciR1eMK9kSLsUjHF
94HYpl2HWHfg1LpSKGPGG55y1o3gb8zHhI9+z/McaiqDzfp0vKDKQLABOCUH
M+A0YoKtPWk16F8rJzy59wdxEcxCdoJMCgZZXEY9q65yFr/6/wALMW/ga0z4
2l/IfaLAP4l+boJUTuyb4ftNJn7GFw+TKUyx/a+1YwldJJZdUUf34jfHiq2m
kg7Bp38dWoTlvXODRJIS9lgczLNpOyJQJvs/HeymapPmQVmnbAAXYSNBrrvw
E9ozz16Qj6lTJr1ZxuLe1Ztt+cwAw15daK/dsmjFxU/nRuRqyKscs/vrsek0
ujoFTa62O/2RG8RdEeTcc7wo7ZSxJInjnk4IxWVYdcC1LaXdvw7cHiyfxXtl
AOjKIqTxKv+jEDTr+Ujtgyf7QGKfx09v/Yi2Dp963AacLe9+mRn2A4ZQn4QY
x7fOXiLcvcGEWvlJ9dudjoZB08IeblnIBeDPxQBvIuKkJXG12OO72NIz51Fm
u5vow9gmkIdMzzPHoHqI1q+uXioZ3ierNIk04xcPmTf7yDysDcvUP/gMQAYf
5ICHQl/lK+MwDJi5VBe6xfR/UP+JS7cIqFN+5R6d5TIba2A2Y6kmy8hU35JM
EgBIPtMe/lkR1xFPl0nB0qjmF+GmBQycMBfAxL6R9jvF7frpHXpRCP0G+5qB
82Mv3On/FXE7o1B4t4V9N+MGkPw/wsLLE6VUVgEMTCI1w28upgUaN5tEYYTj
yPx+SJYrc4L0bjFYDv9bu9tgxP1jQqcyv/2HMl1Z0gpA50IRkJy0xO1SVkXr
prQG8NrSmWnLS+2D0q6tJ4HJtMTvim8epmy0uDN8pk2PNGszc/yJC5NBudck
iF5HLXdK77jBF6pAfyHb6lCKZdcMgt87BujbUEVf7+6Vc7HowuIsgmvZgUsl
wkvZAE+g8nTeLli1tILgZU6ZxjRxVPjOXZ+mB+1V+maWHXDzorSUDQbMn4Pl
BwfWkp1PS0xwh6p9AgDoZO6kKk8H87TWiWrfvA0ETQNMlZCXXsTe/AYw1UcD
MRY4TtXCn9gpGC4dbHSAs7hrfwNjLCIrZxarmuwzP63sWgshE60r+1yeI7Xh
sNBfssrMWIf4euuje/XzaDM3C33il9SAJJ4Dn9f8e/J/jMqdQcgtYYdjuSQw
W/+Ik8IEW90DtotWmEd/5VF/Kws4jbsa+96TFUAoQweItqzCSUdAoJKqPVfj
7qhedYLdMG4MAZ3rJEoJTetoVqWndu6P7bAp0tRWs0Zj/dUngdbXn/zs0YiQ
YMI5nOrI4HRlibJ3M7WTxSlEHtC60ZAapRrQ0pd/Ixkzox8KleeFKlTv9a59
XDM9icTyWE1zS0F5U2S9g1HSh102lL8vIhJ8J6SNPc0zdSYODuIuwj81UzAv
G/vqHjLPdHhqr8JFsSNtNVYZb66+8M1tmJd47r0j1chs4GQ0tUvu3wb5xAR5
TzKNtjAObPKRIRiJrYNmtRpq7FKSr5ngHmVbFDlTs8UU1RTvupptGWiAADDT
MMVHkEj2pccDCkEkKP7v71IUf/WDs9N9L8PcTgc47pvuFlzn3B0p8cm8KdVg
TOTuKl8AfGFtknYTLCE1tVVnpCisBRSRrmzfkMYA4Vd8xEh+T0vsvRDc/Inb
8qb/9oOkHaRMR2VdlakGunlBhL+7N8m9lgVhBlCHCOoYSRGCqOrb1s1CjMJX
xR+JWbg6kxSFdsIpVnmDat07iWK6HogrGSDh8a/ZNM0MbO6jbPs0uqQPQ83a
Zx9D3kkAnxQWKms9jfCy3RofubJUwCwyqlt0D+OjeA48qrfHc5N+itVK+swy
fUtSQbrBpZLlRQS5YWvkvUXvQW0qXJCALxN+leELqXgb1RoZ/1qvvNZjvdZq
lPKLyW0qSXJtbWu46EEQJ6L1MRoFovv2OO95c1iCzTjlps9uvDhPwZO2x0Y6
KCYSLJ09LoZL5f7fmioE5Cg4bee37ipHK/mIFrWEME8JJcWxULkCxkgzAPOF
xzgMqTEJvpDdbDITF3d1srwvxduVfbZi4DzRG5kxhVTCZKuAATy3lQzd/SUT
chP08+t5U1FHZmER1lvZEi7LwxA6aIXBOp48ddWdZ2VdNQMNmNBE4dyOboPr
JNYjtxli9Pxqy+adt+dvKCVezg4tj0ZL3lh/8bmd01TirKWXGgaapM6KwWpK
lrHbPe7ycLOfELeT0S0eAFFpEoZkmf25FWCs3Pi+aA3+ZfShYwRqpcoP/5Mg
YuhKygypUdPU/FBdAZg96aeZ1rumOWX8hpFZ4914zF05c5oIXaqrVhU8PAE0
flOEVTX9TT7wpEzYef2q2bbJQUIwZoR4BLsBTLC/3hld+jp66cFHt9nMigvN
5U0ekbMYbWBtXixuESo5iUq1dvO351ExFkF4kAZdnD0exyp9HIkpOrBc/CMX
gv3UvlkgdHUgaLwmStCnFV0pnwzp139HipsNTFevIE+KS9EvPbKFsJgLjpOo
lzN/LXUwvuZwcTXOaXaoVq6z1lr5iCrJ0p97tP1Et/iXZeWpvkGF6kyz747g
h/IXTHexAjRf3N5j6bRu0GhrOH1dDm+l3wSusukmZ6YPt/cnu3rKulRT8Ue7
3mrECzEdTYlTDioXATTmqgyDRB8p98xaEviDUpe2vfIvm1F7NMC9ggjqlmxF
+La4Qq7s75l/bW+TDRbeJlHi1UpwnekpG4IOZ+p2bZ9XmhaFVKJjH+nXixmt
y8+XB6GQSFQqYlrBENulJ4mQnq10HrfuJnnxmULyo5U9rsHpKexU2+X4rQ2g
69c6mOiURz7ajk/ixghAFRecrLfQirWXQFtF1Eo5TDUjZ3Cruj6Wj6b8SuJp
wudNV+3/SNLxO2q14xcIQfXEKhKF/D4QQwdEmcFeV3ZBTsOURvFaKfqYLcG8
Zg4HffWPF69gwY2KsfNADPzLECA5PQhwMzakxwmjF+j9ylsOdiq178OHHA/T
E6WAjHsqd+likzwT8Q2o+rwHuAjAStKo1sDrDVGADIu+j55Ux03CHhcNKL93
YOjXpUkgSIKLm3gBYhURF4d4p/GipOnWlT280KKhAHI+U7fDZvNg/IijMhOS
+stRLGj9+ftngz3lJ1/hS9SC3Q+YOqwLFyPjtSIqU5DHPI99LZZOPoux+1ps
/TVpOy1y/bYksK+BGMnFPA+SO8HkhQ96qHygpH2h6QSdztf5GJ8++dhZmP7p
ScXuz/n7PmtZe3CX4lL86c1VWq70bIGSQbsIRbBpelq3t4cd8YXm6B3GlygI
rN4o7Qa3UzXtUjHfJKj2KTw2w6l4/8Ff/s2woNb2yxaD35+Yr4mhqKuwg7hm
vjXAUe204SNgwB6ZOuCyHwP6Oyp+Q2mAO0aZUsuwbfOGZ1litOO681UOJSR0
HM0BLNn/DY3WvYvqDhDM4UAtrXEvYe+MXZTI0+2hCkzUitsJhAZ9ALSuNxuY
zbnuYdCq7fQHbSdQk2Ji0xBxVzcbvxAkZkG2kKJodWnMaHmM2bkuGkj54rTB
OT07faupWORdUN4y/15423BfMq0tXBoVQlS7YTznpxA2Wkho9aHRtkjWnuo2
Y6njWGJMtLipNZuJoMJdmRXa0/LF5Iqm2dySB3vEVcF1cgPH/6u0Y+IilK4t
nrlg2vkFt33jznLJOXs/HbmEos69R2raU2VvjyaPZu1TYl3+9I+oSQeAkPfw
ty/Xhy5TpXU/jSSNaI4wF1KlP8UV+X6FPWOrSdgDGN01aGtlic2rSsWs8TC/
95mGn/j+g1jheAdBCt9FkdgJdTff0Xfy9+bsrFGkuaBQCSP++ugNjWErI/bQ
0fq2pfJIIcAsRpCVv603EcXmMagD12CyUBLlAuscIjsIsqp/iOQ9BWSbLQK0
tUF8Pb0iv5uC3xoha6HmGH2HF1ZuHTvvIbBtMaLlHQDeqQO4MAwie481dfJA
4KiaESMu87/+VZuS0SQBfUPuCLXKvAuRsc1oEerlFxEPH5y4oCNysLPuCHt/
HGmJqp2KE8rNWV8XFZFidLyPz1BxOf5NwR0CEU0PEyd9U8+54oogyBLKm9Ie
62GqhWq7nWAM2CIj6pT4GxTY6G0QkjWWIvEpRZHgRj/Wt2o1IQ7PH1auwmU0
tuQuCVyNOZEY7ixAV4z+Qu5ZxKPJKP1MXc5vm4fGQQSQgTghNS/l281ZCSCO
Kp1nw9u061irwEygDDbs6pMMSxLKYE7Qk5foubh947/UmpIWtfmGb0Z6eovd
7qNaQksaq/U5OKTgOz0x1Xtk8Jbg4rc5A3Tl00NOn6SHXJewCmVD/c+eIOHI
ITWCrm5tGCYwPUrnAw6hoIU4Hwgi+qeMTOz3/TEOFprO7DTvWIBG7LjqjBZ2
TRfvfXihX/H12RpXGEXYjnlv77A4H9OuZ7pTwHYOFApM5whnj6W7bp2EOSOh
Xg2y6JiFuR7mPVYjRrABDxR3f52SrDwPYvB2m1kqvNRGvuJCh6tkNI/PiVPh
dOA4H9muc+5oVT7J+OqJ3GAe/ATOiJ2qx/vM/mOYqCiX3dEwAfE1AIariTFD
oQ7ZomkfP3nsZQPBGeB1rmB87elpeOxAS/yOJ5W3P0kpZcHRKSpY8Din4hKX
0y0E82gwx7JK2h+OdpSDxQlm3LUqgCg3dJ/nDWf903qf+FHGE0Qdw4WQE7tv
8w2s/ilwRiEWyGP7PWwVdJeOGDxkD3BQ4qYiRoOjuGA/aJ2ixwifJxm9CJju
+efUKtT/XqrRmojgLFmlfYW7JtkkKV62hl86IQsm30HqZLUp56cBOnMgit1e
KwuQ87us4/A1gjPR3FgYdcorefIQ9E6uMSjpb6fZ9qQm+1fwXGvyQSpQk3ev
Lj+wS43pCn694/t2Jm7uGG404D1YJhlO4dN4JwG6QPQSm225lh+UhuxBUVI+
8jnG/c2y5opIp4UwbzlQ4ePv7jaLnNo3wuSCur+0s1ZkjPbCJs91h0Ru9wcF
11JfGiEA3aBr7E2gojmT84jIjc4b+mb8iMKpll2UrvFWiOBlw51oktqA1Czq
kBYKiF+tM4qSEcqMJ5Ko5XuVqUQoHuwN1lZel4v42wz+hvADMtLxE2FH0RMF
MROcQ4g3ljh+fUnoEMg5oyxpPL/ClHpI2Es50Jwe8icqGQ80S3dUxEADvoO1
UESM++f1X/TJKNDc/GnnlaKMJ9tiv0MH6qLO/o/0bSrRUvAuvCOotWh/K21M
VoJNwPonNvG2KSMGACWIzpnpS47TgZQkxgUsMW6xyZYpeyEox3U5KUeYhusS
fcsFK45MYnkzfBpzcSvucq6cvkowX0UlfxE3jM8QkxBmFuF3BUQFMSRK4VAc
lycdhxgckqopZeRSoEYxyorb7tCqG6BGfHzpIAOBUSvrlVThzL7Rah85SqZ2
0puItdNY6D+XKvCM0JRPRqqPatCDf5KDAcrL0E8PXTV2HMD7KHiOEysvSAlP
9MgCmh4FHt6H1V4X6yvhZB9jgctf5wkc4hr9b1WZyP5b4dsup03Vo06zHJ+p
iva11xvRP9m5r8wrLgKBUzw1QHssskHHFhJ5uxP8N2K8CMTYGJllB2L1EBr1
1FKbOZ8d73SR+5TLiHm/UqfgQmRp+twSeZVumDU7r+a3NQEJQX9iJUeJKWI6
IJWpvE87x38pQdN5Vp4sMK8kbE0iGnPO84oQdkWjmJRQkZRSdID/F9eQI5OH
tfFJd+CmReqLX1jPlC23YSq48KXdwZi97FmmuhUsHzyMb4sZtum07xnWGouD
qkq9RKTxqvy+Jl9w69jd9zuDrvQGuuzVcvW647n4RobPo3y2LOZEAGmuhG3a
/eASPiSaJY/ndSQgJwr4pT5kawb7ADzhusjxBWP5/trDpRIdmLdGYoQw1yAN
JEJq0gn7t6bgM6L3MB3uO4deF6wajKFPhQqlrt94OC3a3FzERpsM81GhY1ie
maHT1DSchEt/kK4OfHsNQccQWDbJeF3PNOyxqZXNOqVlrjDKxkJnQ76Ra+Eb
tQoFkKProMzy5xIdviRalaP1NSPu9Dyuv3YDR4k2fSbzqP4JLrUcTvBqRKAm
eKWIanekDdtaookZQswYU0FL7riXaz8OrtEoaNPAhz3qncnvmkQ7hQCjEtNM
aKfn2Zm9pXcHwkASQcRBQrtCeVXD+eeYvB2IQt0wCh74Lk6k/P+eMUXzcQkW
HTD+gSNtbkJ/XP3hPONk9XjCow0g8p6PG6FXQU72EZo56lyIRNfyoby5TcQT
zmQ67mVlOhj0zyYgqiEjTPadAYsruUpBZa1vJbmwP8maJcajrldGn7VLMawP
MqNOP6vWSoSj6WsQGcLXAXMZmsASITp3WKdV+ACs9WMniGU+lhNvIfNMTAer
oFdNJpgSJe0e/3QvIqKpmw5luwRhA5RoOLGiMbzDpVH7MVzeDAdiZUh5lkgM
BfnMRwkl+7RPyGfq3Hs5CJTAtPNbGw6i5afxj27zgNhdYzbdUoqiKF2LjVVO
tz2vPrHPgb7CxVSS4vYrrYqOFe3J2f2A0a/ajhx6dx5kD/Zo1+Bd/UGhVf5C
WvJAv3i3RtNdV1DzZgPLLNs9OcWOIci14KhBDpaBxTLfRrx4VbZ1cniHXT7O
EDvPE8zacNmRuawQkguvxjXeZMKVoEJasxoXQep2FBORIhnkrmRHKA4V1Ayz
U8kkJpXLejD801Oe+zvewy2NEIRRz9GYjT4dJj+55UwPzOxRn6tl3NdW0m1U
TPBgdP70dvJ2DJpaMcAreZYO4OU/HZR8VjXNp6pYT4Ny3Q0FjvTJUrRfqToD
hPH0r3cdHrWH12SM10vuGpIb4Vz5m4euOW3Ba8up1SjycnDw+oL0D+nxFTRA
YJ8T2Xh5Q9uWTWdJIFlyxIYrcBgaY5yrszUFbF1CngCIOpvbjMxZKgycs+vS
xkM1r/k7ItMadxMCLkBTry7DWUxoppNAYfM2+4A0bjhhg/l+RgP65Bq7qGJA
EI4/JfgKW4G7R4Pf5saj1CEmQ214zZKehZ81mfJj2+gtZ0XVrB6LOPSvNRQY
o8ZaX/sKvSfyhTpKWx0tXD1ub+/Y4UHw0wmCWGh1lQaSFQY4ESslopOhXdnA
Bd52yuU1bLvNqRnRH8JhanUAt6ZbxBy6Lre+JkhxM3ZuvA/GxXb2AubVimAu
B2tmr7Xj4LqFANYEJEUmt9Uwj//Pbgefmal3OmTbVpuyD0wtkkO6XA+HFr3q
E6nT7ESPFQHZfmVeLkllKzpWQkK5dBfXK7f5BKDOSkNUvc/TuFXaSdsaFVb4
GitcHcgLzKGeY7Qulvi6zj8KA4Hgzuq/03ENPeU4tM6BOg7bHL3psRzhBbyG
8RPQA30AVVIfLC/MpwtDlRQ82o+rqolx81Nl/SdT75GxfsRSnIritkcyNwF2
itEF2dDPdnL0Dzg81FqmEfBgrtR7I1jQlvPEJRfBazF22xvYVV7tGWNe1m5c
sKUiGpvrBHOPyfcK7nQ50rDNMMGNsmK+wFEVvpfDrpwRS6ZJkagKZfHS+XaM
3T9JXCbZIGggvhfmXXuwDX5z7l5sUDdMXCoqlH220mUuNeBNjqK0He+PD583
JcsZzs96N9tJm3ElNIIgM6vje2Q9wGYlJUeZbr+Ees5UI6B/go3OebPg9/Tc
O1nO188dxg+RN0h5riDPHQ1/i9Uln+I3JIpOHrTCTi2fHajr3zbSbJtscfRa
XVzTzUieb+h5wjfUBCkgnxF8kkK+Qo0ovIB1B10kl8GMKrrlzCRLn32OsZph
3t3xAK01FNyfSFA9ruSCvotcSBQ+jryHaln7Sp8teHDzsZdyNuPzy6Bz3gjd
+pkElN2YukCUuQraayVumyPv6KM8AA5oxIUPMu+up03Mlyav7G/M5DZuNTXq
Quf4EhhFbCuSu/4taLdH2rz0T5QPithQu72iZjRHtEJhe8rF8oATKeNyvDmr
73uROrz9pZPOH/ZC4VdjFXIEeFdQ5WkStlDYq1mqU0OoDKlCPDxTnWLESfJo
EMAfkJYhQKDX46pJ8E4PEqz36hx77/L4panGLpho9n5IHrqS2CI5bnL3CeUM
pU9SUQqIAD9drVUFr3hlw0AhR1RDxNXk/M8fRJUk3dlkfND+8J7sEQba3NJc
e4SAKuh4iPRQiGOZ0K5D72S+YxVYIaMgD3+/pgCeTLQW0RMbWEXQYwME9mHc
cvCPbhJM16ltCeZJiYCap2dq1ZYcMSqSCZQ0KnoTV1Al/3yrYHrkkPk4B9Y0
iixSkGLV3nwk3kg7FrEjJ8oqCxmGZyv0btBkW/BLupPVVsRP/fViBYTl1r50
g2yZiKYKtmU1U96fSjzXKYKgHxo+NTdkgbswXR4d6RSzROUE0L7b/9Inoki4
lwxaeflAFAi1qbwsXzBEtU6dBHhVHCrH7xYEaJdD0FVs9Z8cFPcRy/sGq53W
kmCWvtH+OKVo8WCI/SXALiffDV9UvKfXTbs/gKLCGl8T3wiHLC/o7Uz7q35y
lmJ8W/his6C1qb9WNWRgSjglsoCJuxN3ZvDA4OaaGvZtSBCneVfHZYxenGrM
d3jRmac+2q1BBMOBCpQTkjfLmPL5yBn1sSgU3pSVsV9aVDlm/GPhzmYsGqku
tDEOl+3j4oBXT53HfjL+VKVDqRGmSxMZ81IgOY5ZTi3Mx6NgMCf80mlW3lko
N6DCf0aW+cTqs6+vos6RUS1GDW7vDxyHj2eety5XrOuM/FFGihDc/Fv/ah4C
uyefjTVCIQzhTWmRNszlEvl27aMzIkDkgjS76FBseO1YTNmz5NmdKHnM8gPd
sAVXg9u2vrYj3G9lTWDOJ8MA7MesTvXNwTfhiePDbAZCkH4G7bgtOXE87B3V
Gf5jww4MmPXb0hONyghVpIUz4xfVGNWto7uVSGVNSu9mudWJHGYvfCtTMUbM
xFWH9ltP7D+ob14u8tyRWkgfNUs6xQ27QMXz42b7MSuxGpFNRsfS+gneOPzk
H+B8xwiZ7t8Ab3nEIdddVeEzMGSeKrEaysFsqvaAA5Df7nR5fcRynyQEUwR3
flSYSvVvpCBmsvfUA5++1QMMX9OqWqbDl+qMrh6pcTgawpP4VmkutElFmal+
CFXvUAYoFsOxxjzzDVbYy8zezz7u8dPhrJizyMFJEdYoKZuBaWpMmFgTWJ5Y
xIgrwOPoDyHBaaPuNI7cLby1D+7qpT1VkjRoyHupqTsAnxkgXL5OEDiy9MJF
LtvSQQJ9osALK8CAmhnTeFLoDu7ZE08Vfm7YOXygECWcGYl8RB7qTsqHgOAU
P8CONdoxYlkMfwCrzOVnGfQoNDnAjeH35dc0smBIOubyJZasHRjNNF/wv37S
iCJHcbRI8ca2KYDBCGe0Sb4pb3o9y9Vt/vzBiQkrT40loHNU/5lF1FBBMlJJ
u+VzFcMwwps7x7OAV7ijl/yzxIa93K+0jSyZ/WK7c2GeweMq2OJQAsxylN+m
/SF0voday0OsC//ZJ6/6ceuOE3e58/JrTCEfMq+FXSusn3xXbLm+uvyTU2Am
L/egNqLQieRhO2WcXrqVvj9O0ifkHHiJCqDM56rUymBsNAXazkcpltIuNd5M
7xhz807du8pRsTi6jvLvQ8Eden27bDmnHaHZmpjiNUKYtYMJrk1NsVZGvXHf
VuCvdkdF2vkqXVFyJ5wcSLcM5VzYGqZhW3oABMXfs49fK+zXmf30zhYBuCgO
mvYh7fKjx9EP8IrhfJljnUtz4KA7xHxzccr6tqsxV80v/8Ok3+5zHL5rWhKy
Qa8BggALQC9R2caOePiVCzG2YZQVQAIZuyhzCefKInWTWHD2ukR9izIhryW5
mWw4WtxNSJxqlCcVhLVmgKP8HaByKeOOAp611uAozuDXV8ru3OabEZdG+Pim
T56pKyfb/MWpje+YkCi2WKw7fPunk9w4y8RCfhIEEpLvPbQ2Uyq8qbHlDhb7
+xPFfTtrFz8sr6I3vWsmbQVXEcYEe8TX+W9PCYIqVpz0k/FEGZXdcXpSU/Ay
YbuyLhYrQ8sKE2PgcbZ6tQIMLvtAOMMy8XCt4+sewlqjqo/jAI2emgBmfG0G
s+b8XDt+NGqye6pYuAkSvqoi3cXLpiAWvfUtxhs9IALchCeJHFaTTVZi7AOR
EYqLjmEnm3trs/+gNsjD5HZkxAzL5VlSPIWMmUBvmzxNuIEosg9vPy1BSVfX
1zqoilWefe0KbgR9wCXf61JbSs/SaTgP0k2alc1MJlzl6GJWn/EV3b+gAa8f
wQYSOzyi3UzQ56aPKCncXTKXxcyC4TbqSKNr5TA1nhI9rgVhmn5fV+sw5uzW
bDtxo5cKZVmFKQu7d+S9oXt+JCercTUpG1OiBBZXTWegEGsU6yYYOWzTr8Ns
IREPhhq9OrNYqI1v5iOsBf0CDlwNy9aIo2SDFQc+jjPI/EowqHe7tkFz1efu
MKhVq/A0fBTd7x0f3TBSluHVte1Kksm+Q1uZju1a8ci565KnH/VhbP5+2Gt8
Oz7u1m2A3y2bg25y2UuvOcNc9w4uYaBVLSvyY7dHkEbLX4P+zPpyzTlh9C7R
R2nY2vV8rhjQYzkHJ84+IPtEUz+OPihV2NpgJxmINmNI+kEoLLHnv3f318Gx
DYyWGoJX3uXALc02c77Ts9iVgNox8zRkfNNs/C32iMbpgEkuoHoTPXYS8PvK
4xZBKg2yLctn3nFFDfk6m83EPtP4xeeqVQdkR1+yT36Dr+A2DxJDE+aJjtPY
UOevlUj97gtI8hHVuMXg/e16uDUyS0u98p+igsIXD8qR5hlYfqSvK3b/mh+B
284ymWvF8PqhBdfgTz+omwMofuIzR9IVBxpRe+7pMoVoG0n3sZ/Vp93p0gwA
2XPwPMouLyP3Tq9DQ9GLVPLi3yOuTbSZDGZBW0vDCbK9JPVAsqvBUm4R4srP
DkoX2QYw2yI1P4c0AnoMSKmgRceEeZ3OOG5n++iO45NvUhjYhye6L3OJt+DV
GIxhbxQRh+/G91l3UC0OBSkDMUJbxXrf8o6rqBnTE6nLUqQqXnfQ2Pdfsw8o
ikPEMzN1ZFslDtdFkUsamzwcCod0KARTQtS5FL7JZzSmzL/AODwi8jDHjWLM
n48r97U2Nt1LpCZ2CG57aTyRAT+rWxuEwVAVObwHe+EMmEE986jlpMRhqOt3
11zUcp5ck9mJDXenziacgFGGQmUsqrSRpUOgQxHRCC9msYAC6oNefulEcC2V
pL3dBnBpUnmtXv1pJuyCXS42nMVBeRB+JEM7sIKVBSIDUoBBZzpb+Ou/vgZc
4lQH5ivsV3ZHSbxYRi8ugvA0LmQc1XhsOEPlXXQ/Ar4dTtvBIVqj538YNyhP
2Fke37EpEEdJawJx/Ccn9hlQNnWbp4VwBxP2y8I1TqXZpjBDHf+vaWpM0iU1
KuG2UE7U2KqgO7IQN5prSo+zbeYdFLsPuTzaQ+YmsHOttg6QYQuCADiDqp8S
ua45N4hubb9h8lJmzJgETj5w/k9rfR6DoBOsVc25meZlbXANB8eD70dwUsCa
YjbbCM3ETaaP3iDvHDrEz4JQKSithu1TlamYeraPzw/oI/unwQoe/yASBMXb
wzDgvjcNez8q7Fc8YXpwDxUlFySALB2G8NepDslVjclKFxYp8YyW6/RSDBAI
Ssq4tburyoF4djhbfMbUV1XgLpPec7SknYMQhQiPNsxenH1anCseuYy/rk7M
mcPmTtVps3N0grwi2Gs0jITViNIrWgQV8m9tc4EtOX7gOgEsjk+9PuQoi7AK
thJvFbFAmkcYZwJ7JqrkD4x9YG8yXarBABTNGElKOpu7awBSU0UMRkXh0ow2
x7ZlH5OQ4JUNl6/UoxCSCOesVxOsJuNOU+Li7uatL16trJyo06kbabc2meNz
S+SftIg88PUC+L1Cu5yHoL5ga+Nkp9dLUrdr2QKXW6QshvEDKUMwiTeI7fnP
YlQqdfNgL7H3geDx3SNqL0UOCgC1cOt9oJS34tOEO5JzuFuPCi8q26SZnv6S
8f5HzJ6rxzB4bQU8/dHJf+Qd9SjbbwPmHh9yeJLXBwQXWxT2+6goJ/ABMSl/
FqNNDM28AyfTl7yw5UY6VGuzeIsiNBAT8ORSKvLNdAhNvdwB0IgINT5wzVqP
EKleuuc3I/CNsTSQEhpxc8ZfZVQl7C42Cx2Z/fb9PItW8omg27E9NznHBATt
tFntToDrfaCZFqDOBiSP2Q1BjKu70rZw8Bn/cBY8/ljYQRzpuhvfDtHLkzfs
86IZdcFRX4ReF2XEF/O+BmqxioWx9UZjJteQUq0hBmlQiOTMf3Yak05QiGEt
IPmoZFKEiV+PtBAPbrcEB5sOJRr7np8kp+LOP1twm8rJqfXE9Nqcu3/6vVRr
atdi+2SuSVsfRMHhVPV+3KrdgKN4SCJ5ScuXC8YChbM2YDloKP4RoQfpaVJo
EUWR+lMGw/DyN38pAmYMA11AQmbDnNRo0WN2QBJQy1GhT0U0dvS4goTUeBQu
OvOvMritB4Td7AQtb68tBRPbO3W9AUxwdjcfVfrvsiKT+ODahoSuhaRXD7zZ
bM4l5gdQAoe9Gt89OUiLOjug+uhBIkij/6Zn2LaCiYsTyCzmuXa6W+/uQxqy
hJTeKRn4fkOFfM9qM5G6NxZ3EuXIu74/Fxbm7tdDItAHAnI6AQGJVAPLuCf7
PB4UrfQUdSXoVWJxACOwleMWE2dUUdVMFpBBY+o5I4oc9+P8r5jxpiKhpYB9
POZy/hJHlLer1WWYt4OQE++DGAYmpPx/Wg1jVLqthnG0j4tzdtNo46/sE7rc
DPboNiF6F0BFAv0nB3OthFTnAZcJml88CRMirHY7RnJgB53/zMaoiOBBvGDo
NF8kGbvF2x7DZCautIPPivHnFR/qbK65JQNF21KhJcvBeX18gWTXWWpYiRaG
0MkjSTHj0RSW59KH32NZlwF6VgCazKf9MqyGn2ih5eFVyfKGYcaOzX6XpG3e
HL9DTxhJIaWDPZgMr+kiu7Tk3FyRoGekrgD/MVekZfL7X4/xkDTtPs/LDo95
4rkQJTGZJ+NNtBoq7P/UUskRN8jbfLfTX0GJjf6NucK3jGggss3vXoxu6KR9
YX0CGUdb+IImUNcb/RmxQom5Qj17DOEusDC979xVcseh52+DNOEReaIF6Dk7
zFQlp8f1CZzqNpy6SBunUf3dNjIci7WWyOPZXVWl9DurHqmZl0PIVmO19aTu
M0erLTVY9P5VvBxz57Zs/Hic+AnIgshKpsG5wBpcSM0JxnX2voJIpdbuuOI6
XnbrV9b4OHLbTahI3VtFH0SlGmeZW+WclbAHe4htjsefOYHooAsaP4uoHl+A
TIj2x4DlkQl7h699zHbRqglfS3Msn+0SRgXxL/AOPtEqDJ5MwwNA0GojCfTW
nrwyZ3gkTV32atogHAyKSiKrLbuyXQJGftbs2eH8taBH/Qav4TpaMFKgYelV
CygI2keO7/aXzPNpAMeJQtZSgND8ib9qWd1MHklrwWVnE23ToJ6qNF6MDRb0
iBnSrrk2tr9DV6r9h7L5knXDZMeRhrBe7Kn2mn9tq3KKJQSYZR4fLj8EJG6z
Y8AOXbeSM1Ub/EDc26naD6ActTl5t/omIkpFGNWCLJTVPeqL22n4e3moRhr3
KbSPqLncA1pDvtNRATw9jknWDWSR1ztfXuuV9K7FpTFER4YsYYrlxxLSY/ym
AeuapT9CLho7z0s/fRfPJAennwQQ686kEv4hAZ+HXRPETEcYpFu6xDMXvQGJ
+E5og+Z/Outwl7Je1oDJRvatMRS7JBoTfUqqgx7HYnxBN+TVLEi8LnxHinBm
JZb6d7zsu52AsyW1VhR2UDNCqOXm2Bxzc014U4VBThb9RlQvdypRdJF3qRcx
06jYjmPIunC5vSTw2+nvVJKncFf44o3GT2t5yudcykhMpuxkLJeSQp4b4ufZ
Rf2o040nxWSeCqT2nsA9J1gdg5BebqRpSQqzaWKjjJ1UPUvxx85smJIO12wZ
+K8lhMAEnTOvv7pSf3bUPCM0QW6oO7nOePVohDHEYPXFG/5KUw3ZlUUbYxSi
J+glfz8l1qkUQdsDDlpDetHXQUG+6WybBDKB4DVuKqaawYKDSPDwKgmMUaYc
gMatlATOtsomdJH9o7GG+08D+5xoQR1s/c7Vfix5G/b5eySKdxVhfAF05bc9
Ju24Sy8YsT5BiqFHEdD7U/87RLXxrxRFHLE6u4xKfCY6LsshkngeySYPcJhA
45izYKmidvnTezDfQygdPVd0JxzNf4lpjCw/axAmUCQhz0gDl8rzPHcKaXEM
pfAWfGIskfGdnd69J+n/3TiuKHPRlgMPYlZ1EjfXUWb9ACecv+tWitRVMG9T
ENP7J6HiAmMVted6WJCz1obvJOf5H9dQAOl56F8uKS54tfMp9qew2HggRDcf
0nWZAwjgH/NDSJNduHMApIHxANT32T2zTU4bIs5AknOSV81CrpFyjrEvBXOy
/D3Z+pEf3AbkrIcZ+lNBGs+isP5+5CocojSx8V5QPEKLQz1I9dZpR48tbTo+
NwSiUblBzOmYfycMoxiCogf+HSA1W6tuUXF7gMlyaNkbaHQ692Sb62RKMXKF
JQQ/HtwOQpRszpD58s+d07XB3ftrGoo5fYR//LdkUzD57VFmDBWb79k3MYLy
e4n4uHPIpMH3k+tFG+FtrIkwZRW0OJN7EcRMhEwLEGmUSdH9D11+Qrnbbyef
LIKmvxYhYTWyQEWCGBZTgJrlZakF/EJLI33n8xRbmusSrkt0po1w/gCNL9Iq
hWbmZAtc2gYlyKjct4ENJMO+PVXNHMynhzbkLzNi4yxc8KdMo2OBGpeygDvk
QJW/S31zS66J73rXHJC26iMiQ7Q25MMMbGxPR2gPCrT1Zqd2L7gicmf/50BF
y9LgpZ3S7hTYkXs6Abx++iLkgi0gkmu7RKf41wlJAuhCQVUSKrCxYiZaoIau
oBP6P7N9uXSb+uir0lAYvMR4UFAsYT+Ch6yzpPM7s0nrIFft3Z++brQ1cMGw
sBmBqQMw5NVKsP3Q4BGYFV6yCEXXohENzYkKytfZzg4jI8FUPGoWfTyVT0MO
SHZ9w0XqwQnuuuKzE7JxMorjISHG+I+A1CNzQv4Y3s/7ED1wzFoZ10m/q0fL
0tfHmgIZSmoT//R6YxFU3MpL2vays9lsRWSQzfCQf+T88AkLPFCWV/JY1J/V
q2n9w1fesWlj1QNZ2/syhdsSENUBTyjiTtAYRM2aeBQWB+tSz9QfW32VzMWy
en/6L/pd+QtzzqvI8HVTRwOPqj7oeYHr1C6AjidXwGkg1eloiF4TlsiLiWSd
/YbQJqAhyebLVvRVwmcfLz7Q/WsMGtkIJ/MYy2dWpsNjOgxHcKqTcTPHRkdj
ZIv7VsbWBC3z0Sx5fRu+2aV0HHcxuQ+ECfUoD+6jf80YXu/uEmz3TKNbGeGB
tx+a2YPNkSR1JFxHkeZErod0zc56tAYT2zSj6WHRXUE73buX1y8EHj3xl6Wt
FleiS5aHi2UhH7dM3rQrLv3OprTQzuvmifxeAP9dKg7p2oHaJo2GQmiPx7jP
xSnlXJwMCmQSdfD2O97pXp3uqN+joQNqrEeDk/3u6weHq87ZT4TJ+ZDWB58p
IUBCHeFEwr9GyGKLjYWJ74jbTwFYApTU68/7PeXXiK7CJCLokHUz8w9hJ8o1
BUUfOcAbpRRmukHbfV49iZArpTLApvjQwnIdmL8zcHDu9g/aXkKD3j4ZWOtW
i1FD8CkZjpDkJ88P0nw/de0NVuGoVqC7t2y07Lb5E3k4TrFpgDU/ccPq2Svs
hKAKCLnU+7hbdUxo2SK3THGEFkxQ+49k/43UhzJ0k/9mKG/Xi8OjqBY+P63M
qJbkI+v1KGJf55Pn7opGQFjFQVR8B1GSNaAV+6GXZk6GWiPId6jrZQhQhCu2
AxeEuumzbxU2cZN2ucbKUBbMHXhAWEfJw8RaKZlAhYXoLMKYtXmIiXp+7HV5
f7un4EtU3LOj3yLp2vll5c2b3s5yAefInH6AWsQ6w3BHiotxcLDuIR5wLBrO
tHNKo3RH3/zWZ1psDDb5tLBWlahC2eQgoOpxZ7R43DzKCD2zxINP2Nt5ul+w
Cid/2ZfajiBUI7FmnW1NBoApp2Q+rt0X+6wcmJxlcWAb7HUmUomeAdgHh0zR
v6dJA9IfyRkVBYOeH/mXdgq9snV/JkcBHjo1w9NLiErY2/DLum/UPSZMUDYZ
4L8Lg36oRaqRV04pHte6QON9at3reGfmH+5ubpizW+4YMLQCDE+IXuFiKNWj
bQoCgjcqUkcpGiGK87bWfrjvp/kn4uNpKsjOg5gWFby+z4eIBKxzM+KCm1fz
OOn7lUfkRwjIb1eSu9+33bDTdbKfYNXu78M/FgnmVIGJcuT/B+5WajsIdPZM
F1M9QM73BTn6AvLAsqBjridyfHzS1zvWBV6zwc8CRJDxN3q/4gHCaCBsZVYu
ddFWcUbiiUlXsai/f2GWuJT3lJAsV5G2Jtj//RZN/nzc6lRnADsJXhS273Lc
P07q5geTrM+k/zKQFkSOAs7OupdwDRHkmZPyQ3FA9XSQQZI/MdmkJbA1+0hx
v2033MP+12ce9XQ3OYwwaEwYSkzZ/rYkMXqBzaVClDjJZifNpF3Kwa0V5+Hx
r9piHLipHu7l/CPEsOy16BS0AxkcsaTJtoi1OTxNzVIW2yKBVwTUGm7KQyYh
RSWppjUdoEAWtHJJZf5558rf6Jhy2DTuhNyB3IynU13B0d1J4ImJ+QN8rifq
oTA58QpTCgPBUDCLFPwcMsvwusvb9Gd5A2xLFULE3GB8HT+cQc+mnCSGpjEb
kR9YXTV2Oisyzo4dYoMpDxxeYaKLuB8WSTv5tk9lqjzbXWBI56e1ECWt/Ae/
aVlFRvmTIZp8RhwVlgbGnCOevK66h4QUfSlzvuJC6PxIc5V+ZjVasbbganD/
xP3tarq9qtww593bYhbMzrGY6/tTCKA4krUS/GNEAKN1ccb2xMbNeJecEmuI
vAuTBXbQabo1nx2crmorFx7tfh2J/NbZUdEBxgfJ+UtXEpkF3Q+rzLkbwfXS
atIzRo/Jh7VtfGbsxvLHiy+p/PSHabrf3GymaS7dk8WAfJ2juoq2bmjAsE6f
QDwL36XRT5HnADZzkC1qAppilVpQgzGdyhmQR+JU/QrWI+zdWq0a/5xfDzWy
pczdt3M4o9BqZ6zeNV44xko2hiYgGnVF56TK8Tu0WEKzackXHMaHIhZujLyN
77OLxZgGeYDtaWIBvGnZaxPnOUHpXEaNWKr7kFzP4Ay8DcgtnstQnmKQTvOe
R1djKiwafl28FkzzA3h85tS7TtoKmZSOlo5Bi3N4/ZdsbhzD1TNSvTsMjxsF
Ec7yxzksWMRRO6rz7wyIg9C7bXDO+rRjHUsvWKuo4Nu3qGJaXfhTV7Qr3VkE
+3pxdtx7ZSwwh4U/7wJBZq4+04Mw4OvQDY7rHUyTyKqmagTkiApNwpzlR8Ak
3kvYdg+WR9cTW8Dokqw3fc12GHGSk+7j+1dkZM9yaR6iCgzyWqrJKmW3EVuH
w88JMyvihk6fyjCInPKlZ20lGxveX6PzvMKT1/cYFSrV2Sdj9PUwCxX+gkfr
XhL8l2PC0M33yHEk6VzAjeDePOV2Iye4IvQrIUmit5+ZbR3StVF8CKAi8Fg7
YG+wD+TCBr3JEnYyGN/kjUy28VL9TAXKLP2D/EmKrDelg6nqexpTbadO+jNE
XbkjnCxWt1T+m2K0vgOiWvucC3NvGsdo4ZtQJwrNgrWV1yn3/vOSenVyK5+v
yw774VcrsMKNH1v3BJlCeOAlpv/mpU0CV8IPnI/S8RrGnXrkrnWJZtVNUYuq
mjl5nLMAUOgvtjvF6W/YsslSaAveYxzbtR7uBP2elpedoYvH0CK52NzAECH4
Ry/oCahIg4Y5auq+iYi9C98+VN0I5wcKDhHfCndBU1urW9idXIa1k+lwFQWF
NrosA0p+GBz9vlskAgzWe3vz7SbxcCFf3aGZYm4W9L6FJnOMCiVrP5quKTK6
LWCNPVKvbRSzRWmqQSEsNYjtBFiSFonJr1htIMcn9RSfiEl0yBEeJD2ZX7Oj
smX3fA6SaYu+6gZ0vz4xx37T44nXAd8J0eNGoYZ13NACcpayeJvRs7MkaOtE
+A+woQTWBBueDWR5ic7AQ0ExM6nQdCOK3VbretQmzaS88MDG8y8JqtXHZocQ
otVmbShAkQQvUccL3ePsxC2hffWnSdIlu08x6l/Ch06Qx0D2WKmcr4W69tiz
xGXT9dVVQ7uZnH1sv9mtjmQe+fTs0IEXxddD1NN1GCWEZBSG39Y2gVmVnAbx
hdlT8Utk91zHYsNYMQqUkWS9glivF6qSxmtT6w0M78j0CUYsdExkgTc5r3VF
BcR0d2EV1rEVWIyN1QQ4uIhiYwfvWDULEQH6Wb6CWSbO3yF0kR+t6+btKLr8
Q6nJFQpLztWtDPQ5hYkRRktCLqx4ihIijftk6c6lWYVXUzxHd9eGRDhAjk0I
p5qoyDJ4YxhnxZKkodcWhs+N2lNYpluuJoLcCH/mdr0134WEBuJMl/psTa40
IlmLP5qkih4ghz4Db+g5aYDJ4CBStX17D2yt/NfRw5Xu8mgLH4naV+Bqcxjh
2VqNXWumPrZPH8zbPu7e7QPII6LsbRYejKfFsc+jTKaJEqk2RoNvAl36xmpM
Lfb6lXyP5Fy1C+YeOt/h4n9GTnvQV4TwMQc0xoW+PTcJxLF19XN724eKOMlZ
xycglyEPVRAZnfcJkQTivrEa216UWoroVvanJ9ZQtJi7zMv9E9sck64fzVWv
F8kfbuPyvLz9czr2mqix7JtlM85JZNrEnbml7QylMvE3Xb5uLyKmgYGUWoyW
TrchYQllhcfMEQkJmY96QGiH6G4AAeuOJeSpFbicTGn6bOP1r3R+6bLZbr3/
jdzCJOOb7ZUsZorFFXj934vl7th91gMC/CC4EtH7neyAopgps1DR1zaVznJj
2EUE6qLnAlyV9HBORYg+CE3NqSy+VdjVKgO/ZtGeG9N2HuM/1J+6d/o7k5lG
W/Iv9ggq+80000oR36SFchNzsXm762UmmoGeULOhOljTGwJyFVCodPyOBNnu
IcJdrxUrnJiPuIPWmCFBlkjw2qL2wQSPV4N2wZR1iDBErljwKZzjzHTBWKxM
CAPNo/+fXixjl+BMkNM5ToATttBio8wHwjlxcSsD7i2mcs6KmOKqFETPNYys
kN79Ic0rP0P0czJTAXhvpTr/v50SxBJazenCvxd6AH0AIujtRODC/iMt6LB7
c3ZiuYQBz1ZkhsYdB28C+nrBRVckGQJZvOsJPPNOjOCY8mbBzpNUt8jup2NV
FmMLM+qGnj2697AnrOm01zDUTnZO0ACHPdCVHfaHP8hVdVwtf6Y+SAlYjTTi
W4ckdMcJMZppEurmvE2lUUZYcwtJXbYUuH9u1hPMXU+G1ZLXMah2hYeRLDZ4
XnNZR5+ich2Sr57ZJiRvcoaB1GzAUtLn201nRL+yW2Im/ejwKH9betewh7zN
+jUig1xsPowAagJTo2BjZMYxQ1/i/Y8lufTgV/ASj3jC/SgdIvjZ3gCz8z0k
JL3HMruiTPxWj5LoTn3rRN0D1yVIBg7z52h4s0UJYqHZ1N4SN6dyHmonaepD
UQbref2EukxWjoubFbk0Fg1sWGxhQf8MhEZ7Klv3su1CPi2ku2BkTv/Yrnay
jmOuwvQTd606xyD8S14SXmrZgbKtUb+fgnJLZwnAi8RDlcaHcAjMZsyu1QeI
DSgPRaGwKk2gTtIGGDlfvK58oNrhey20aK43JovbqkRCaZvUf+oBQymKsKQD
rMWSuUw20zHW5BmbEXGHLQfIjGe0sWT78ALwt0ggzIiJVOcoTqVBtTdXlqOt
r48tU0DPjQU9HHzf36RPD0RmQLh+3wkVmOu8ZR7qqvsB8YWhoUuUeCmzFtXl
irA4nUMZDwz+DnPWjPrXTeHz+K3+bQAg+5EhqTgvvimDw8jnAr8OdeRPcor/
0fa/iZ2OLhOvZAw6Fj7WDKf1+9FtwheD2nESHJre0zAxhRfJFtPpGq9U8zuo
tVS82APh3GUcQGo6DsUtuDLDFWqeE1PDEZT98xvylEkym4ajU8LYFXfAThks
Bgl3bzEe+Y/TWLigpnDlysV5zoPOpwWJ9soPR1dVs2nRP87Igyzaw1DhJEXJ
LkoeTpjgJT/g4b/YwDD3TBT5aELEu2xURVdhM93XLvhnlG3XvFmwE+kynQyn
jJR5WjPriW3VE1NA6cQDwf+G/ZUxTri3VfkBFktXktT6fM5vjR/oBEF+PAx2
vtp/HffUICD76hdtM46buHyZu4e16E6JPw9CLD/AwlS+HS5jVeaW/OsRafcX
quM3CYHQTeicF+pj3OxQifHFcmBfzfnt5YIg0shamL6m25K7L89/y56Qjyv8
f0WCac3joGMFxlPYtW/YJvj+83DXVLzZSh06WgKPg+ivaYhW/jlO+g1eLRzo
XBORYbvcMaMnicYsP7ZpBLQw5bRwBso9pU4EJHI/hzqvhgjgGQ0wDlgcVT6y
2qWjjTBw/YXWimSRLkz+W1U2VPqn3Owfbh/6vUx4XaM59fD3Fd2dNq64MPeg
9k64VTt86T7YQnykISWFw6HTSDZXz+4gVE0l9KAivpE1XU1DdnrWPFQFBfJx
JZIRx85ODTRTvdHcEzJFdVWqxayzXwLCe6E/nc2mT8xBwRUVLh6GJV/ojcnC
Yfxi9fJg5dDv95EGWFjCWFDxuxUGXwWREn2MxWKG5hTWXw71kJY5lX74KB1H
Jk2e+aqRWqOwRLHoWP4/wNTNYB9rodzjX/Rkw20oiakmShSKzXSarlUwWo72
H3LwGY5yEuVCRsqClgKsLDtYBlSDpmhrDDtxHJRKz7G07iRoqKGZo4SKIh32
B0qvm5f6kau/JFU6RMsdEylJ/NENnsWr4occ+JW3OoabtjlauaOcO/Cg3o8q
SEnvNoW2m1cCw/75KfvVl2aVvHyScbfb7bQaYCTHii2Puhf7ZBogP/zrO15C
Fn2Go7qbTt/IMJPmwhRnPE+b0q5O8epaQjs3YHSqDkpGVvyJgYt6PTU9WJPn
icUlS9jTn8h4dZtebhTJsvhpF3iFk6JRhim4krKDVVU4QFloV1XrTbsFqfel
dv6xQQIRbtGqVEsHtJTqivEMw8AMPhextgNZCI/DyvcbQqwH96oAoIiGRmvh
yxZV4aNbZ4nHFQ6+OeRymo0WsM/t4CYhdfV8SD2RbVSqbvZtE+DRF3dZFnDw
RCboECQXqNItkMdOueQfCLsQwE+FNjLQnlNNLj3G3YfwzwwuxDv13gXqPAgV
MRxQqAWuo9vMcSlcpDd4raGWma1yPc6T6VeeYh1Ud8/kLAVRq7aR3eIgtbvP
6rkaKZd/vC0QBpn18dsV6KI4cGd7IEWjELZ1e4kKheckTT/58DiZNkDPR3Ps
ijlSwO+/YVB29jDnX6ma4I9YsylrGvdRn8u89HRAVvMl8MLyjGavEXSML97z
FL4BwXKjiW/OQ90xlI+yql8LN5q/s9ao1Ehf8jNIcpM2CM8NEvTzvfTtDAyz
FRqcadxXpTswtCQYyUzwQhldgYpcKcSx60ymxOdXK5iOROD4a0J75x8TrD5m
7htjUelok3zS0tmiCuxPGfcXSsSnuj19Zr6UXZe+C+c27FhRvVHX8S4NmJrj
IFyuS89bYjGAtjTGbE2vSVsE2sB+LFgDhN6wfu9FZfE61l3Sm47dUkdZlAy9
vvlPfZEeJ70WvJnXIKwDRGlqvZENUZkTdMKljx/SUSp3CfJkxM7s9t2wx1y+
NTlSNrun+EYG9nxVRkNlDtEFLF4BNqc/TSi3e4RjRAB5Vh8iQgIMAIE5YCoh
V4MZNi/1NXRwZir7g9oLfTqTQPbUxyiaI3RzzlCr5x3oMJBHUXGtgsPL4YHM
ne5jYeHiIRAO3Cx3E0SKjMQSE9EfdilfoZ/Z5LgNLO1qxmJs+n0eLpMVZtsL
LLuzjxm3ybJNxxTN3AvNT/i89UZ1oDI7rxeLEDH1tifsOdd3uvKi8/2OJj2O
BFU9pUJ0KdqPuaZoVvzuZ39xKDNVdQ1HhlrTlUbouQLGD0KDE8SMOBy/zgIm
+l0vK0f1HuZdUI05qNhiyT3R2AOtUF/79iE08Ll/g20V+rlD/LtYWbc61BfD
BufdrhMANGI74B+UkaSxmErRLQXYzscszMY8cBRov3iMPqHHCvFxfq4Y0QqC
5u80odHw4WwzToiR/KIDNVjPvOwzBHRLDoyXGW4LfeRntK0j+5V1FLcv92rK
6P+3+ZX3FM3qFGoDLYJqI4mESWoTWmNeyqmI/abJcheLia2E65rKXwbiT/2/
Cc0Zd74Y/edLMt92dNnMxJd8MXyCwmHmGxS+J0i1j0g8iq4zgv8NgwoO2D43
YcmGZqnUpiEHbfXFxhkQiWma7y8CPIsLaP2hgooDl8flKkJWZECTRCMpiojM
iwpDAFu9Hl4EuqQeNM0nbbhgyan8tlaOPsq6/5n9gISTtnjcnFI+xzqtI+2q
Oas6QARmVAFSiIc/Lr1+c9a3ggR08lCFUPegVVta7E+m3zTmgQSfM83KEnOs
X7hXV3nGh6Cz+IhKgzVRtR1Wv0LSUzus5LhmhxTEqQA8FqwBIyZhUvcb409J
BaN54IfK99Z3KwJ+BV2ds1+rKp/iy+3x8qq0L2/t6SLhFTvA72ita3+RiXjt
x+tIyA+rNLLQRAgGgd1Owi4NNJhlf/Xy9NhMaoeiDBsVAKKJNMdakTpe3bY4
RcKVl+GsFnXUfpa1RfvtddKMv1rBRRC3vgF6k1Ux/hraEJBnikees++dhKAu
ijnsIhY+GRhpmRo9XXy8vcHXs4MPixXRMEZN1xsVPBNBJAghERGsNah+aF7V
DI6IDfFYBSgN1IbdLoI3dj2rhVAvZuTn0mgmx62IyD63ELhSmGdlT7ZHQvCW
mvfLB3s/Blf2vveQNGnroG9bjEn3EiqW7Nw6qoI1oTPjv3mjsGyV3XH7oHvd
KYJ62yI1SWXnlFelg1/+UmaWg6csW63nS/y6BXB6UjttjmPmo/Y1zkKA/j+S
opIBxM4YpdmPg0wCkavGBx0xIbe3Pkn+h69QXC1KFRRrR090SAGjXGRhwKZJ
MaK5QShGgLBH3DoZeOoiUxti46QluGuvNlq83+QADy/BkJP5rBXTV5R8flR5
HHKVFY4JreNDVd+UHJU144l03yvgsB5pL3O/+j0gv8h0oBZSvhNAh8Le3dB5
pM/MA8f3laHkhD+OMKbX1nlipMcpWvtwZs5qp3hocIrnrss6lLUr9275MHfV
bmHuT3YzjzZcy8W4KnHQudPDlOpogQambu7+m3X6ux7laBxe0h0BfOzjn64I
ir1ZsFeYpCViH3Vv1WMOwv58FpptQehKZU7PITjG9IyMUWk+gqkzw3nHgHlY
bi6k5Cw1+5g3EyJww1m7rPb6T0RzUz0nTfiMF5bxDBtPoyF6okNgWtrzP6pz
aHXFLxC8FawrPo4dG8pb3Hm8KdjANZgNfzqG4/jTYsXkwiZfaJJIXZof4IfZ
iDm6lenvLfdq+5EPZTddy1WQAF/XGDoYcG2gZz6KIbmC3psaPZoIeMFbUFTM
+qHhYRLQXhnArEFD6/LrLpo45E8qrNCUS46t+TWmoNPkHBb8zfEuWfvEaq8y
8YLL5SePea2s4FO4lCF3E4/FK8tTMxxKDNyr9TrW/n7at+5jREfYmvlCdONc
8JbcIpz+zdU9ndj9WWePSAR21oJfaEvbRi9gouHrmM86CWH+TdLdhgVQDitB
cne4dqzm998QHr/5D/iXWXVa4JDk0KGwNkZvJjKp/f/qvdc33icKAhwy+DNz
2UnkQpRSibRluMXyjHDslLBvp6UJw9o3vsimg42qjWd60bsJiPwN8n0YjpP7
sWP1863dc3TJ9WELtXQ+HI6VVBvZeGBpvELMEktEcmzyxukRLokbHSaZ4CzO
4RnAlX4Ikt7jtAajcBSokZAhlosTUGvC9XJ6G06d8YY9z/Epv2J5mZzfT7JT
7D305VimpyRBHGLjF6SOnv0b/by+i19xMkbIhTQTUKMYNshEMvL4JOaPLt7t
QpsQ3s8UmQ/Rlnvsuqd+02u7u7R13wl8bHs+QGfvFBakd+gahENnKyRc4pxz
fexF/IgBa5zOEp3L5k8k3HfykR56Wu0hARx+63nm29o31gsygvOAtbxd80BB
GcalL5oJgB6b3sry+63p3Lp/9PGZcU6IhWXDt+nSE1MaRicmExiiF9xTRGT9
XWcS8PKvgKjsd7SMibU4JnaDxA+eQls3fL4sF5lUhxANK1z+/3Rygvbp9Yy2
xL2wzLBB5hia/Wvu6Rl1xiBpqZAZAr+YZyaoramNstltxolDtM9p3YA1X7dx
udYZ7hCobnm9x2uLPfmisqz3cGwAof8QMBPj7TIoIaMRFMoTKAVUfWSu6Jyl
KRvm6d1eh9FSmqUfWlLvJSgrPDu/w5HwiMdV/us7JVndYAdxdsQsw/ryGS0E
nI4PNM2xX6Q0OreHJfPmPihohaoJH7IW4sWDi4D4phhIfxp4WuB1dyZRHbxV
ZIq1VaQE1Q4yVJN3kStOG07S40GSxxaUJJtbubrcdES999SmVq8VkYeF9zHl
Li7kGZKfgSGpu3O3cOqaaJBIKF4lbCimgnhuVF9G8avvN0x267lDfqfxCEh2
ZXkoxhKYGDtLiEWX6leRML8S8t53m0kW66lZVrEr1a/kJsrTz2w8anwSxrmT
aYSKKomOzNPK36F87r31n3YBDcewejFgQr7gW7Lq37gnSMKDaIO5f1elbK6J
e0ZQBSjx1n0tA7LzuT6mV5D/T7MJX5HZydm986aD+R/810Uo/xbb8ihzjIck
6X/OxTUZ1iH8A2AtRYj1c8PAoBE+AapEJI2POV6gRzqShgE6yByePldBIG2C
TEsCghkAoxDl8wpSob6r4xo9X3SbNDLKop1QEB9NehNThtBQAbZd3WEVKbMw
I0aAq/n1TpBDPe5JfGnaNOEL8h9dFoIa925ss8uJNsebIq0sMlaO89NDtH+M
iW+pSeb1tTI0b/+CclpJUy5S0T6YscHqP77JC5rYIeqHWK+GybH8LHTkllp6
n5pQ4aWk7mNiQc34rxsbWXvF254pBiDEcceoKLYXl3Gw/UQny7FCf3YZGcKL
yoiA7q8EGl9vYf27toCZAzdjht39E9qQJkiO/4Rfv9GAVklfNZmXnLil9c24
zJgVllR7ipvwvGrvPrItqAcYToxpKvCW/o1qBqtvihMwleTeWPHd8lvqeQ4m
ZkZYOL56ZcgG0P0svNZy+9MVwLH2Lv3G5GtISgKj/o+Tb6miZxxzraI0vsHq
DaBB0fBfLtzvgTWH/Y0lOlxh88n/WohRqBnwgMCth4IYDpyzG9p4Mtl1wGhl
+BU1L6HcSPaXeZoSGcfsg6cUvyAQ+RImRfFq+k3oqw3IRyr2B6XgqF9gK7MO
Vc8dXIDd/MO9IqM2pXHtCFCAo2sYezRFV3/b3+Y1jfHoD/xziLY3g0UJbrWM
jeMRZSEKdlZenEyw6F3Gb599OriBJ3Y9mvSDvJxPc2602ZqSJyZajvs4gZdD
bYoFKwUJtWWNX48ne7n4WcTz5Rr5pcX8st5TMoba60YwMNliYLKom0y2pezG
qBV9DIRbb4ZAQyu+dADTJgeq8SjGxXlT4C1tdPbmZD2NrJgGPWH3MOvYWjnh
t4V8EjUTGAYEfcpgNl3zRkpakBkWw7R+7hG0FsLjZKdB4RQv9wAtn7AIilcj
xJBjZj4yP3ACxPy4XEv6RiX5+PD0BIm7AxoLsILAdTfx7yBboRF4SQKmkwrp
UBazSb3m1Crz45wyI9Dbjw5u3PZRcAC3l/XjSUDElnckobe2L4qc3B3HPPkg
0Kxrc6ScCodkSLPYH9xMFjpRtwtj86Iio4CrD5iYATYxdChSSTaptI7Y3zbL
4dvMPMBtW+jusRQtyQMJ0WS+/YQD4aRipbawiDk+pTVnOVZkeUSWHJNpsJYj
lExzMfJr2symtltxJJs6Tys42zNvle1st/CBmFZyFT55MZ+WoMxG5+1UHVfX
WM/hzQkaWHRvdbHO5IsnseJjavotwGS5e2Lm9aRLdGk10tW3dGH8urly6LpW
/Gf80Apw37+7bNhjiA4Ja2YxnqyW0aF0IRdOhof0Adw+4UoNPM8c9oOy+ypL
G0nNy91DQegJt9FDUaXuvz0DVhLJvs0GKaBQWNdbMZR5Yat4e/Q5qUoHEIN1
HBfLPMbJtemwtBSypzvFHxMqY3GI1q+pV5fOKB+XkdmRo+nQZ3oHl+JkL2lv
D+bdyE4zVk1JKyzZCMd747cXrB+jHqXxOYKqRNsqj0s7SAWht9N9ciGG61qj
7HQ+HLdqI/vypjnJ91NbM43hZjyr5P06le2t2tpobgVIHrpolQRZ6sHqld+m
ZFvSqVeViFOOXyICR53tQhQmWnF+VxK0kloaLUzWeQ4TqO3lXyhE6MLRYUNF
WfJGE80tgH0LFvNyPd404q6P+2tntMIOPLWQclX/slZkDbzmzQr4z7zyRIY8
5f+HShEtCWrINu9nuM6oubLhjzYg1xMzmtmGKX2AhZ9jg50ihULbro3aUbWn
vzves00U1Y0PNxg8W5ekM3+i91v7+BV+2hIDT4qVXp6IZaltgk08FxclEeWu
wNDxnvZ7Zq/dOoVpaJzETens/NA+08EPTgbVSIQx2q4tSUaPJewYpAIPqOW4
S3r0fC+iwTHMX385Ep79LYHuKCGV/PLkrkBPRq5fm/R/iOGrW2R2lsstRG4C
nQllRMaFJlNYa2xbz15E2SuP/YY5aWPktsInn2qKhtHayk5ZcS4D88U7zdi4
geeYDZeMK0vl2FwGWPpo88b0KxXX22+Jn/gf/yqaXXvcmUiAEVdtMVembmYF
SHo9zN0rhvNpS+RH8fMFISIFKtMZ7P09Om68duiv/xny9UnYUISXJs4YOk4W
bG+1J1VENJK1XiNWC+Dr0Rusgcnfviaug47tp3A+yQMF8xh7sq94hoYx87I5
zNAvTp2/fPc2uHjlOOQUQJtF+Izd8LyDN5BXO337ZMeWJ28Z6qCIqHDCu9+n
2iVng/uQSD4Kqt1tHH2vfgxtoyhbL+06CYvvF+Jhm08p51VN8uId/UvpHLHl
q5MvHVxq9tlCYG9qcNodQhF/XXUdeY1CFawOER/GjtkiJAtFOsSxh6OwXGmq
z38vO407fJ2JPHFBCK7oeVBIi+LifpO5ySuWDGRPEw15HuyR66sLqmcWjtol
h0G0mw0cx/VjLjTZNtWxpJ08AIIsfKY9cyQJatoB5rSXESt19RC6EshuBUWd
nznveeUIXIYhn5waNomQfXlGpFkulIcEKzpBiV1m4Cz8e/OHv5uZuC2TGrwm
ljWb1NMjh/PG4ZmBj0iGAeNxVAP4w+kTObA3r/ATabu1nS79C1fHdWwuARox
C8PTKKTCVtL3LQQh12iP5s9a+iHyJ1nRdOFEmgJ4kpKfZdSsW4rssNSfzMAL
MYQD17O+QCGXpqQ3gnQd4jChPgMcIHrt50Kc58/VLTuQVsvzYhDqdrzL9nVr
mtjPaKXi6njRn1GBOBjyH8i6hpPuTJx/I7HIGeCwVLfIf1y5nJsUQCjma6YY
Ak2cHCPg/J/H1VFAJfkoZ8b3hpOExkV9uV+8QtkSEAEwS0a84033UszxF27C
bsDiw39yERq6sTblSsaofkFK30QmzxusvTskt5RAPdUJS2SOtaPNl5kYflzq
MKe+x/QRlN4fFzsKIF2qXjf2rGRBu9M70Xv3mMdMeuOjs09//3+N10Cp8y1O
wPjk899QJCRnADe1kx7Oi5wL3MzilTlfNrCS/jfgyvceX7+uGZtdNQLQj/tb
r4YJNoLI6fmCY9w54AgQq0C56Y55tezicnOBoopJF+6r92ttwOnrYUBMIuHy
a8uIa5D54YpVi3CTfUNUWO6SiuDS+wOq0SbL7i5IaJXv/eoLHzI1kT8obdUx
ZMK5PQnnTRxjQVwtBeyYgAi0wQkOJBV7UqlXGYPiG9JpOyiVu2gAgHcJPWMG
hwoewhtRfN4rE4T5orP0jjBlyua23iTN5T7Wy24Xza7twTbVKAtx3tfujJOO
rVQ6Fe3RxHWVrD0GbnDMT4Y2qZxxEipbQw4U146m79a3mpFEregOTN1BXCRa
5PfcdqTz406ii2S1S2qqBDngIKGMK/n805g9Dce3a7FE7gZ7erYLNSe+Pi+B
966fVna/ezk/mXv1Xp2cvqdHrZdyuiS140vMBr1zDoq64EqTU5BGvjTZdZ2I
SLSR9ITs8NCmygJxGl5rcvel6KFDG99AFTEaJGsU96KZx1ldR8BtECb5aKFP
CMmohMfyREU8CTGnGa1yJRb+gJORuIOlq8PYN4YGizWaVBx5Oe1ns2kJBmn5
z2Wqh9wogXKCDHu67Qal9rSKDnripZaw1GXH5pcIpTBdS0aW4qRlBxfwuTyk
LbXYkbAIhtEhcxHTINoAYl50O0109tB9dAkIVO/Qq6hP5MhpVXuVlYrADPD4
rkCMbM1yfWuBfm26BRzJJz2Kermxi7FC0Qsbw1spj0ga5B4z/DU1sQdLq6E2
u84H3C3+MXWXIYQFF1rE8qnKiAbmSq5CiH/8lZM3iy3b2OJq3TSRMrO62Y3g
cx+AVBZsa2dGMoHMvlXRDQiOnHr0g+lck4gQgbI7+yGit3ddSB+4Ez0ijlZA
OxVg4acYCaAjP5CqvkIMHmRU7aRhZxt8AlAe7wklEnEh62SDrqIlrbzC9eqX
rz7uz1gU7em+GU+mjwT8CneIgJ0/JezrmEFh0yoJHcC+K2WDqm6r4S7IK4UZ
UUoHtf3gfmOAVVN71H7iPYzk07JT442PyUfy8FEb1EnoXe3SlCrGgds5Ou1+
jkWfEMlm8zNtoJuFhZOMWiuPWE9W4wpVRXrhqWwPoPejw+J4FajLSAqKeqF/
M8EnN/6IvprAI5Qady+wFd7HtW7GABq0HxU6cA0agp8I7j4xLh0wMlEVuwHU
9l0uSwuWTzE7w4oPk1z3YFDGuRc4cKh5Po8XgO0V2oFqFa3tkVhNeTe5z8SP
jsa1hLbduUc958Goiwt6lLpeT+AC/tm8nRxEzyLPmV4yv2ryCBXpH0lRiP2G
9TTRqAHot6zcAT9YrvO4i3xj1jok4OZGrwy/znC0rqYUEXsvqZqHso547Tsx
8pvDw+ZOpMlTCmGPgeCTTTL5dDmoqLgVRQqv3zobZfB6966xvOKxqi5MChDT
ak/RZ+LJdAfjz7yYaQ3MtEbzBnzXINHtYShBhHn+XA1qqymXUi7+j2n3GFzV
eF6+g2DmSRzpxDbrO42Tb8whiG7p0lsMlKDSdjZYYTsvhd93y01YtThHKmb9
82FEbre/7G6XQvFcXN4qmxfa9xB9kU+suLo2ZMpIj8wkMzObKmA1DIppQEJG
xHqJP++GBhm7xmYCyavg7oNZ/quuNtgB7qLlXM+4JJcxCqBpdhKBgiRQBcpv
jzGkXrNV+wW0A21zrQC2hmXfEPB3jZNe24H5sfC7RPD06lF0KokKV9LJkiNe
2Y6yFaxCu4KBllpJwvOf3eGYyOaAEUwyCQ5Svut4pjDQTb/ZiYDzW+J9lkS1
Bgjg7nhds4Vo4sza5H2xiTkBLgIMXPKV8amvLN+LLAXuZzvu3nygUQfCRIoc
xsJp2Xn7+Sc18QgRmEf7Hv4znBowSyAs5gAUmFV3ytPFhCVj3S0l/3Nwrs7u
WDlvd0THZXRIHEw4WCCg09QjJ+8jV/GZsqvGT5jY6xrRh0NTGhGs1+EmA/AP
MfkB0piAZdFRyN/2QHWGK17YNFyzsNLUrJDYNejlDjo9cf7ZGfKmh8b1okaz
n0qtPc6RrJP9njGj5VaLhKVTcCCz38LUyBycTDhNcQTo38TV/vXpzocsToZX
Pp7BCgMTHdG9JKy5DWgdWpl2y4Gic7LAtN+R1CVzLR651LbvNl+uz4UjbHoW
dK/rnoUMI3Aamhvmx+OLlEwDmvuarBz+s4WzDHyQUXuVjLaNGHsiRSN7izEY
+wUqHK7KO7cbsJhoWMcBTB+Se34smQMSdUWgOPFyYtjjVxCUUU1/2N6yMqNd
94I+2nOZWprB1SJ/7h4aKllzS6sGXHJ2IZWOD1ZSU3q2H1rFZWQUoy9kNucZ
RIFfxaSEO3k5EOfYm4l8nGWLJ8pUdkJdRoWPJ6YlcnTvMvGjxTcpuwGQSUeT
kC0XLZY4tASERHCj1IjiuyockxrMvzHtn6wZk8UFGncpHvpm+DbjRy28QLwG
HI8vpwL708iMkcm7evMiHjKEJQEymfrvUNJr6Df4nD1PuLaCF4xMaoTQSoe/
RNcGs+Ymbf+tbniXgeze6s4hZo1BH4J9g5PPILbo+tnSXRN8OnBMkkhuZVQl
8pULvT/QKfqBQ917DfalIJF317mZk8vFcHBMll8rscBaVJRzbemCQi6VETUm
RWYDdjntkAr/643lO0Qi9GnwiBlDBCrL7PFTN6Iu+P/iT85AGDRjG4XtX7TY
pOi3aw0C/NAKqBwtqE15L+GxoiTVOM9Ov1Xsgd9cXCbQLM9ubYbTAk9ounrg
0H4zI60o3EKX8YdT92EDK8zsTZSosiyxTTi7XRcZQgz/ed+B4ZL6lBPFJZp4
rC30nQFM2oFGGU5I6CIYVqTCvJKgY7oVYs8ZzlZdQbbLoffo3/xMNdwWZ/3E
oYavqJxtNhhT8O0PZytovyAwbj6gbJX5MFoyjtzF7Qi8d7IMjRVtYCM9XCpR
dkQ8BwM6rK1KgGAg9KoO72pPoKtGZ1O3sG8cFmi748WsJr0AK+NkBr9HV/Pd
cdAYOXsFEznNca97MFLLfLyJv1MLwHe6ZK0HB11d2Kf5PqkLWLv8Uu2gTTKm
nIHLmSYNi3zalrsVOS9yVnU4l+FJhs1lc0QK6LdWocAGX4BwxyhjBR2Xx5+W
5LIjbv/Tdsyy12em/5JgWwp0MXUAfsES68Trkh5/H4XwO70c7MDSeCd3yPyI
ZgGHOKznPKhiX9z7HPi7/TpY4JgqPqz09z5GVFVdRs+Bt+1BXEnX736Ku8/P
YCOOYhGRqjqYNwDnF/FmIZb3/1OiQ8/wsMz7Av1F2swFTP6jV6wfo7uB1WRA
pEqzmTi3XzjJGSk1IuPDzDHr/u/OErmgiBIqbp6ANotB6q6ggCbOxZGe9C6t
aD/+b0Y3pXanToozF1Zt/pp8vuvxYRPd7MLOstSaMx9y5TIuQxcR5veJdUVO
om2S4NOags87GVgiAVVKngtigkt1RaYP35OtCP3ouK7SxraKVVLP39/B+j9o
XKdlGEXm0yFffomgww4v1P0GH68A05875whvGXZmAn+izJKl43xkbs0H0jfZ
e3+eWVnxQrXSxW8MKu0DqQ0mSdU4aHs9NBo6xjzqa6H5Hg6zW1c5jLTAi03I
TXrrbUyDCE5m0kpiWqjM8sQ0pD7ijIucCJzjty0eKdzG54Inasv/BVGASHc4
Ktn+n40MQy78rFykoxyhUJc9k5KwRdgjL0VguJLOJWJKW40XiiLEDumVcwcG
uSXnQvcok2oCPFBWg3D4M+ICKSdr0ndYGaFpRuarXp1ac+cLp8IQtUVwH9od
VPZweUl36A159k+PD1pnCra/Kjo1/LeWcXvrMEBomun0yWrEULb6qYUg5z5V
zqiIz8YnINqPThaFjI1Zq5/893KFiMLORSnhZxVpWen/vsq2fi51S/Va9yk5
bxHVhTKqx7LMtbRu+71+AOKWeeCHp7TQo5rl3Dplm817aW7uWgvdM8kwbhoN
UfOheKW1in6F8+52GUlTCixfQUtXFPMPqNX9TgUKMXcnU9incChJtyvVBl4z
wgMAp14qFNzzo7AaNfF3rJ4MxCyCSee6MxtM1iloQ3FLursNINUwu/bN9R3J
z0hi6gAyAr6zWTmjtgBBeZSCQFmnQ5tfSTO91k67jqFOA97tw8w3OOEHRZOo
a7zt5tQJS1dcIJZuwVN4epVIcfXEQ9kJJZvckF2teTHoyB2veOMhn4WfpgDV
PtI1gL0OniXOmiT3CCw1EhB+XEWnnsoW5uOp9r8XrtQuC975vnPl6FDZ90eq
y59D9K+ii7AEodkT2VqSVHDpkCw6exphHrr3sEXXSeqmfjXSWWpjYxI1tD2+
6trwE2O/86/HP9we5tCN31XCYYuPmMAAPdq0UI8lLHV0lbKPtm+jX3s65BrN
ojU3YKMAmeeF+YBX5kOLiU+pj772Z+43qLuk83HUjGtdv+rvikscWCel/opO
lUA6YAs9MvBdXNHsF8iP1ngNsCWDBGWz9v2faFPvN2PFqCqgB9cY7xZEALzn
UHPbgfZTrrhN6g9DKU/DNyDqCRt2u632OWCkUM7WmAZDtZS+8QaJNbN676Ea
IpgTkwQZvJqDpPTW87vCo1NLzDEksaJVU457Ap+zUvTZWgWO6BkdvhPQwxcf
6t8ctRYnQUWpD+txO+oap1QaaY0pA5fD+GHzRVtkS5uPfrXprYm3JHIoCntW
fOv9vBf7zFus4S5KeCkLXfENvoQjeZlgzXcJNmGS/NxzzMrVxFAJnp3Fc0rO
VpdMarrycBtlFYiF9JFAz45j/9sN02yMA3FwCun1rzbPUo988sFg1yQTrrTd
mDnetxWZwyhUkG0fXfin60/0J0hgm2/YaiLYRFvnQ9IJ14nzh+GyyDZRhpFH
ogu7fUtMxvgdzdwuKUUqT5jZc4+xTMJpOpVLyrzXbWfPKPys/29c47bjcJ7K
cJe/HASHEVHDDIIdFbgnrw30P8Xec0Slx2toNTweUmiYBQyLR5eXbqoarYAW
e3TgJy3xECLpmnByiy+meN7KgM6ugGr+ki4wATe7mNakz9c95WCAR8UGhfqT
OG3gMRVbWSgBQ9H10olp+cx6tWDprDQMhN+4tClfUvGeJKmmV/Eg/V8nb2V+
4ims5tDCnp3bYlSG7FWwJ0cnoV+9dFOTxqCkehbiyZr+6DSVScdr6AloRIte
EaCGPZ/12OzWEN2m2TqfF+p5RRIkY3xin+77yFjmcBQitVTh76Z3Mxw2aoNm
qr+xuagtu0KsLA6qUj9LIJz2fopb0nVWfAAVyj0okalcf0Hz07MxIfG1rC2S
YueFcGCkOwXQ87R/SESQfdO44ZJm71knrW54CwCBdV3/6OF+oplaEduJomd4
E0bQHt8bffUCCnnI8oO9EVYb0R/ORqArwbb9dqxfQWxOJQd7JIwm3ftJ6VYg
zEpynX4MwvY8FR+bHZsMGtfjSrW52mwnQBSSv0jSebbVkYFjsfNUYpr7yeLq
FdRY5bbv5tyHOUdDbfC0813OniCjbprBf5tUrzhZI8Kl+NqVPIcGIiCJDc8g
/S/iFpWtIqxERWO6QuABeCrOIYnEVgComJ4yDtiJcxpqUREdEw+BHwp8vt6e
UjfkUA98n1aBSbDUW9Zz+JaEboGsKQCme8p0DVbPyYsFzpmkS6GzvpFeHJUi
NxcJ0eGQaouFXVc1Inqkes6g4zpjsqi9/ujALi0R2nLJ2ew4cJfQPAMhznbV
zEyDMk/ayTd5cCjpJkG9sPQlyTt93fBtIwn/Uh3Civtn0LZgR5EZ0UavFeSo
+8jchQpKt2JtyGdDypg0x903k3/8ZT3sYmQSxY0OdsPo/mb6qrkpGHPS5QBW
s67iyWYnEgOTJN+ikChtV/pYClvaa3L/OT/jFC6gEg3+nNZknmZJT1QYCs9b
hZ8bZJnG++X+7ICREqsVhil3Xq/0QewoqBR/PsMnFNY6RW7QnpDuon2AHgG0
uSnkOPmY7kgBXKDiVODRhgUQajhJDlMSGcq21i6+tkQ1F9McMHP/cg4WnT9s
ma5FA/7oisnW64jPybH2S36hNg2xJ7cXKfDr36kJVplVreqMksGrqQ5j6Osb
k5aZJ3LcLkC66U53m+9igcysJcA4M88e2GIRg+Ao9p3ngThW0+FKA86E/H8w
QEm66e4QrH8+vdyFZvvCk0T1A0eEKfFcduhd89OdhySxLxM6q4sd04aaRLa5
7JkWnpGq4XgWy5IUc0l8HXmxhGHuVh0M427VoqHzorlTrA7hgMXQOrNNAjm7
AgLawK8E4f94+Ko4CyWMsGLV6h3V+M2qY0r5HBSXJ4i/8ZleGwmUiXzXlCAk
4aBwV3sEEdNyXe5E5O2NR2iW6/U/ZCIQII+QvEx8zVBC38kuV6Q=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "sTlVzHE+yhAN9Vt4a+7yJC9Gw9bfBRq6xv9kCe7Ng5psJnHruz9VrHCdetev/ZiPTJdBJQmffKsGhcT8C1xHmtnWp2phLrsA++mCi6ZvsisBHsXsEe07/2w+B8eMNZubT3xnRLX8hyEfcYoWZpsP3M1DFemdUhSKGBtblrC5P70SnbNX6tsPF3y1BZk1iC/CtfkXVJdvvd+neDISHf8HMgQ3zyVqVVLAWr5Qxk5Q0qTkn4wPEV7I9sr6rGAnqqLBKOknP9YgXkaGBJWlxETylhtgOJlU6Pbhc0SZqhMkahXSsWOrRqzZlYPkUWV/X0Dh8wMRlt/+2OuqjdsOKrBkmN2uGJkgb70tralVnYw1gMiMDwaJ5dZBYX63Fm6lkpNOCidCitRUdoiLNwXCnqR8apUQJpkXLv5gtJcVAOrpO5zlhQ6379DaQkDuOJiaOjooef5VeoqiVfTCnupVMW5OgZKGaSIOHl1pAqsjTYT/99EBiLp0UA29MWx6E7f1ryc1OZWrLC0gqlfR1hjkkE9+XYhsGYPeqCv9lYacLOFuALndfEHbfR4rwS8Ed+yySOpAQPT17Wj1qkesVURpNGjB5RJ7Xv6Re2H1AkdqNDJuk3fbvnQjyY/dew8i9n1pbOrBYlplGNVn3VKuuJ9zfPzy9d0qehFgKJw/jJAJ8g0f7uwGn+BDSNmW9VKBu2fLx6Oqr5TT4hjyr8iImVm5e5/TNT1MQj4keNZO4xipM1QDVksmciptrr5s6xzs2IecSef4FHayJBRWGCwQW9GXdn2iANCbuneHjDpc0kwI/9hv14qiV69q/C1R947e1Z8AjQOaKvUjm4EHGKhV9Xm4RJozh1Mq8bJJlwBLI+nO48yQnxdL9t6CIfc0paYcOzGTqJlONL83uEsIR4l77ktXb50Gk+5zxTBzBy2wlHwY16xCBVNT9ZVgGAPsCTUr25fr0X1mMQlbqM1BWQRdAtslcRxwzIMfVdBb1bLxU6GS4oxEDo26nKvEfcb2sMnv/NBsuF7P"
`endif