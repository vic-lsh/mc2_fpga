// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VC0GZ55qsXAbExiRrDCuKYvLhAsS6sAHRQrpsr39ZCqAB1xAtJR4a6gv2dkh
th5Mv/J59BQ2DUWAja2zUCLCIV3+TJW4M2lO3uQjnvefuOO8QOkroYHPBNcR
Goo/5/FCcR3MjhKyDqaHm6PCCivggkL4IBdM6xbz10e2b87tNERvCJcgIuJs
0GLMW0rSjEq7BNHeMugVkEGX31/iKrleHJuEiam90wmAJxdCqbZagLGRR0mD
catLc7fv6E1OO+nw4vTFtUwSLVE2s3IzYnJ3ONe8bgJuOtLArWgDMzj4wmE6
VOhv5EXBJdGGkKOguNk8otFgLITWHxOACKTrTI07SA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DGyQt4x2vcqDNIv1GzoeXnuH1H4sUdZ3JVAab5390EL6wbQ1zarHUqo7cCOb
wOYzz9SyFYFt8L9dT5jL7s/OGezEkPDCrgUQqzIGzxH8WlJjoLT0te1X7wGE
1j3hx68TPZ+h55FJw+aO8hTX4EZ9WlOSTzldCUvpVSqxN7nhAwHfZfESIhof
qSj+sStJg1D7QHPD7p40Is2OS6hOzto4z28Cppho6gGBMXXklX7fG0cnzda8
upsH6DxmFyfk3hFk9nMrWh/zy7m8kS2LpzdJggJsQjEVxSck50ugtPVf8BSV
AC4jmwS9NOp+Vzn3rKh/KrgdyLySLvnw45e0lAjE5g==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
e49FrYsMiQwfilyxiqKgXVSsT7eEvNGnCLjai9rC+wDHVGsEGxFqkCXpPbz6
z706f7MGltsz3DzG8Vel11H/PZAiiuUESnAJ+rEVEspGBykZSD+1LFlHMiti
MzpXVBDmC4kaQIExJje0G03GDT/R1D2DxjicuBhS/IBL6g5l9tq3X73L2Jbn
FFTrQndH3TCjJ2anyE51ZSmpALvgrWwA1GvjxgNKQVrK8v2y/0pHmOh8pm1f
p8CKTQEOPfxsj3BwMDqnTJii4LQWC5xf70xuc5MC3G+jyh0pynPtMSyLMGI3
ltEjkWReUKIyTwi9kR5iPXT7qRqRTcNVIoNyopLeYQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
b4COYSsSrI5Wt5pOAxD5kAS77BlT5Xmdhyfl5ecYEv2OOwRE2vEQFwiuOh5+
Iy8iBZw/J2ndLSxdo4+DG4Ilf4edWfv67tnnCJNdy3XJw68jjRmFWd4qLImp
KM3PBtTIqz5aXGBTKg6xsNlNd6m1vSMkirH0+ysgdRMENJDd3ccfIjx3X060
ZrlhxpZK+ZWQrN+z4r9yNYqT38a9IhfyXduJMDyGIBdRfF4DDrVpIkk8/LNx
cqhX1Zm278riKaPyit72tYT8BkuASRQmpQyLTLS4ZVvTnh1RdNMNIXVTMVT3
D5b/yu3Ba9prMi2QDFhZNPyJFRzwTlyTE5V3ZYlU/g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hZcOcTOyOnPUU1ASrrpyyiWpdZKHfzObrFaBztGSUt5HlZ88z/40Fm7uhYRe
u6VqPG+QSGAFrH3MoI8Kg4dhmzSF6jGE/a1ZdEuL21+ObOXlAsaouwwmh4A3
8ZuYCXXwO+IeT+cgcvT9DZNF61EUmfg7VI/9hkjV9UIA2djhE8E=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
PBkF2IzOdAKzoZJEA1dcsaDA0yx7Du+36ROHOpZthIU7AgFN0bevUDS5HX62
Ibvdkx9uP6gYa9dGp1X2EGXg9YMNXltH+AsD1G+2MUYIHhaQAOgtv+Cqr3D1
JrXV13baNn8Rq4zUmkmX4eBLIiZsdS8Y4jZbPbNggMHNsTxzrvPmq14lnxnB
Tq78sLbEGyNRI901YLjTjxhvNoakJ91c0p4gzm4NA0pW1qr/o9daYD1HGLSJ
rFadLhhfdIChd2pcffLPrllZ1oSzbhcmMuYb9SZyCdAdu4ICPN6/TZMApUbH
9TcKnvPQHH1a4iajIFzkgiDQphFMsgubxr7JwujNS/+FlNgxWImNf/N7bTCW
Eide2HqA4MgwRsPeLPwbknIQ1WRnP+vCQ5suHZmdfk++PpL5IC5ByqLs8XZT
ihsaOz7Gpmk2ilCk4GW7Kq+P+GBQRgGqrBkcEOrLXayDtcO50k5Vgs+Z7hn9
x3ZE21MCkfFLPV8y616R0Hn+hgykKf2g


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SzAp+RgIgCqpsDhKJ5GAkEIe5xdFRF7p70F6ut427vwi8ep2FoXGoxGJT8BN
PwebYHm25nL2/TaFp+ZSu0IH53IHQ/qFQGHLaWugp7tmfYppyToqijXbh0T9
Jh4XNLqWwmL8JNNlF/9GzMcPRl/mR/yTtrL3PEh/Hl15us7Y6k4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EkbX5W3uhbWj8WPDV2c6W1YhAPPduyr6lSFvNJyGAKutdjTDVqO7tdT2VeqK
1EOrUU/vVcpeTaiNZxTsNZoimMaJcxCKDn7JgRTI87qCTLWjBRqjNpdBuO9n
kFAD+neJ5JCfts/d154NhESMDi3atqBQCyfFBM/A6lipYBnNjl8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 46672)
`pragma protect data_block
FR4ArmZJYjqr2MmaVL38foXd15Wr1KVRB1JWtc5nG5GRY9vwBngz/qHjF35C
1CFRU8rWKyskMiawADDn6iKn+dHmNH68nNjQYXGGyaQU14WypvRLYGBI4v46
RbTjbxgI5WfOJAf5L/Gd3PNmExz5q54Na0QthW64d1EM9DsrC4hoqlQZYLxl
4qV35dmklfJaUJcfGLtlDYBY75Y9DM95IMz/cv4asIpw8JWZ9wbXQZj05ckV
ZiDIVrCFn/2SCJFvCJiOrkMIjIQhW4R/0eqh30M6Q4BlKH5RERVTJYjlUOPJ
18a+hNSFQ4tPNA9wFtN41KfFObuT+5Rh0KspZ3jxQ2fhF8WA/ADALdJEwSPQ
X2o0ARwoWWuiRqCMeiCWxbZ297YbNVyS9T3iiMZA2JtkkMgIG3SlioviQXM1
V1feyNe2mPbbLdTZ/GVZlB8Sq8Akuo5/XphGtLg5hry0XY6vwTk+YU115WL/
Q9V/jf7g6z5gjH/NGtRYQRHgPiVXUjaSlpnHnGj6YVCIzUMSvn9hlKpIbG2/
HyUPdYahJyJ+DZgGhN9YoF8X1goM5qctBNH4V/9rHwEBkkUuxwCGeLUAdx6Y
Lb6+06pAe5a6VnyOddCWc0hqVN36iOQrqcIMANlx3+awKXZe1TsLGV2yxImj
1JY+VsgiVmfpWxAf6Jqe+QEumAA2spM1hR7avlzLYbP7dbMyJqL388GKPve3
j3b7iyJz84Rt9j5tyv8Skjxq/hoE+kCp+Q4JulJiGKfa1HJLhJGRB1chugQP
BovBm+B7hRKwboxg/7UCpipKPZG9F9KNxVfuF/O4CW0Wpc4n8D8taHFWUjOC
YGJCjv4+5VCblWgEi9kqJ7wau8SJYxOWGv77NXYNQfT/b+RIJYwxFKUjhK+I
LNsb5Wn28SY/ZGzS9+Ikshs2mrUjR2pN1P/EGzGDqoQsLZvqNS1eifkAN+mA
Yl5JjZQLn/QSHhB2grXR2iffSQeNTFtyJ8q0E9S0Q2rJ/TrzEh3SlHUB/Ekm
NJEyVgIFwKgkiVzw3ZmlB8bhFhFpeX8ia4a1t1WKZxkl9tSPsEL0gP0R97dD
klZ2jt/bDCiQqwfogYQ5WIRRTvuU3yYFIHsdHVSr8tTPl2bJ4u6iHTVdFKsv
4qWuvfciKwnTSbS2yhhRv6913wGs1+LD7NJNFkR4okErjSZ4G7g3SpgDwc8i
oB1OLOwALJ0re3GY8EyW6TphhaleMkxsSgMfunmo+q5U7faC69vMFXEXcuLF
YgDhAWID9S6v6KuS87YrShcUxWHcbJoA6D+JI3f7+t7MDkMI0Sjbj9Mifk4V
t9W1bXDeDHa4Orboi7gby0RQAEs46RrAnshWmiNsOOvYwJaoSA7tDbJuqxqo
O7+oOnOLDq7ZSMtMCBYo+qBsoKVLafuZi2qTHp/PuG+vbrnEnyCE3pXvnZbt
cwkxWhsDR1nKbuRTC0MF/AMgjc3G3uv7yN043YAoren7avmq1EfrYKOEqDR5
eQuX/kj2R+Mw17w45/Ilskkyf+upR9VEr6nL8q6DYrlQOfDoztjDLs40+3Ms
XnUUbLbXGoO16X93MBL5VnIX2EhWBKu1R+EaQqqHFQ1fBYmQ3fDLCsvIIujt
L8cnK062R3lXG2g0Dz6CMTSui1abyN7EWIeSIXSk/+K999qhSSdPEKxUSFX7
AHFD7/Ku4Dksl/BlACFf0xIW9L6BJUHcLmP+OUcveL9XOLlLj1LfYsuRSmXA
Wvaf2DC68Pq4QPLcLUuYp9ukUil7ySOtymshp/CffPZ2CFoNSuIXBcrA12xm
oAgqelDAuuwV7HweAKmds6vtRuwsbdeltPz/qPavQQW2CcaS2x2SDsY6FECL
kLDDQ+IYbJCYAsA5oGwgos4bcpV6RfsqBTtIM6R16yP8s3FYiuQzyQ2fGwOb
aAXOiIgV6KjGgJSRKjJ2WltjGGL33U3RlXGNxmycCJTPPWmH6vHdCFGDqnXf
934k58BZh1g92a3HUSQEBpXQEpHlXJVo3vZ9osK+tzhQqxABXk4SU5IZySBr
Qx6dn0RDRFZjCm0P7SGSrZfh4nPZ1dcGEt28aJldDR9XG/9Mx6XeuNo8D32N
PHrwV1GEMHrcg5xiYiOrr7avSRLD9mBiGkeVz9dmcJRtSG4rTlQ7/scyKOJe
yyO9nnnw1Rrhi20bcZiXVrRkZdzAppgQ3/+EZ9pp1jmSrizoqm24dGo2L+cP
oUZ4bWl8r3kgmS0S8YHC1HXgdiV1Jnm0bva8Jdc5z2SQVkDF7ePhzDfg/KOk
CP1WbrxymsrLJStOBWF+ZPc24PpB5oPa/bk4K55OZPblG58do68oueaqQtmD
GeRxcCYPhBxxrzzVT6tBXuR60LDO18kFkqTDz8dtp/Ld+CrFAezklvPoDiuQ
Aq9YoX7Qm5z9sXCZ7f5t/16TEj0YLiGdSXFk7m/eA/Lr21Mczvy0Rlf3BumT
zxb8RYnjL3WjTVtv+dy+Xj/HjrbZKnAf62o53Es+ub/xHdojfG4aGKFkDNwm
wU5nZeDXfXkmnK9JLQU0h7uptAsrFLGn0t4XNYIVOkor+fC+51U3XAerHxa9
XvhI0Pmc1jxQ2z+v5lyNIKtd0cUmtkCgWGrr+DM+9CSKt4L1SZ4CET7BOwXq
fBGRCsUSbTZyKskVt4zAlQcW05ozjwPICXnOwyE1MMDcpDDJGAa/I6P6hr+X
EhI6pHuh6qiNW209C4YHWsOHhn4nKUgExbNML7LcY2+XhRBHpmHqNLrwU2cm
qohw3vmyo+NjPZV/kbnNCAOHlk8EzP+ahieVNzgxgrv3le75c526T01CFwX0
30G/EAaVDHgA2rct8Lxa8LfOLZUCex6C64ZEE8PW0Ev+XTQ6gdkQV0yrsqB+
dA08BH6osW7QqWaokF38WkhEdV/zHQOafQBArtHcGOBNAXjOSfZcjaZrLt2y
BOWIfjPJpC//+6nCz3Ax4A4jBQrpkJ78lrMyFCs2cVh1CIATTDyEu5BdVwPU
sWWZJjRguUEHi/hAaiCu2wuEwX69nh6eMxW+iNfH3yNeF7b8l/Y4S1hlOzR6
0eyAzAfUwfUQVaiwotDLiiw8S23aUp4u1Pz7Y44109QNIygBhid5lqr6n2Jt
p0fZVAQckwBI9QVwvN5DldopEMeslrtWSfTX9us9QV7wLb3Y6qUpvmsO75B5
0xWLZTCzdXsqMaJxobOYl99xXw6jx3kF66/yVlFKcsdy9eO8kjWGAuZEYrYo
sXiOql5cVpZneQLVYh1XY3bBNPGOQ+BANhJpaUWS/fFDJZpNmpi0opEQdsSi
2cZzUUFmdfCOWhsqAMbggmYxG8+87ua1fJpwoQd8Vzn9zdYy8fx+La+LQndg
Qlm/4f9WDNs/65H+zXQZeKE2qqxq9HoEzbmel3uT/9is+oeAdR/8Trh3rlNY
0MocJqM0WK3sBUYWL1EjHLPEnB3e3rRY13cBYaqUvs6Bk0zdnzkjAeioOBFP
TPeuLwGIoDGyPkyGYAAo8FscifEx2Xx70CneN4CgOpb/LHf+xXRf7XrJTKiE
iqsVBKh9Qp8l5VuS+nW+2wEX6NnmxUasvjIhyzxrPRgYEyfWP5E6BZRwAR3o
6WNKqaErc+4dt9dljbsuCO2kwtZceAZyWUDo3BApw/lwu9BYSmnMJgdz+AbY
v2m1wV6o1c190Ys6XXhyoSSeLF+Pv+LkbLsrm62rMrscq/h+hD9duSVAWhfQ
ZqwbDltYR/6tBubifERawJ40QDSjFVJ7zdNH0ShlgQ/b1y+KHAKEerY5WE4m
LkdmB5auFgydl8K/I6GXOeWSIKEdhaCPJwim4hk+uh1lnDPNTOxxf7SgUDWD
1jhWK93GD7gXGm3DP95Ymkdxx94AgLnLJ5hdRFfWtuUNKyyemJSMPKw5TTBm
vHwq2J8/fCFx2REczkW+GzpUlPOP46YQ1It8W9nG3y4xvl6H04Q/V4iFjerG
yMmOvlT3lCR9uiZNdNXgYKmB9pTtAxVmx1Chetq6O0fq+Y1Z5u1N4u2sEWom
ItAHSE1BBUvnuvyzPQFe+lIqS9S/T1J+t6vjwcO2OvTN16p//KZSNm5obvVE
yuschtnX5qoVqY9le3wH+RVF6u5WMddfz8chfeGXMerlA9n80Mhq29FJYYGM
40VOMRubMEfMAa61nBR+RKMtHuoHZ06OcwKRbnYMv7TjlSLzih/3KbV/3S3X
WpxnasJGP/2Z2O2QDLPjfgx4zRb+OPVsSihpltcuS34UzPiJbx6qWqANucvm
2JV0XZ6yGWTSzq5+Lh5Sbi2j+kFmUp/UDMK1SSOKJgpOFFd7gE+C4sS2I4kw
HAhyOLhmqVzntXfK90D/oTWLnYe+BeECbksMjStIE3Kd60xf48dIzmdC0KOQ
x7zikoLYtbIwsufgdTpzzX+Q1fiHtg1L2xZhiy8fq5rqUXkFs9EOZ5MtU5hY
z1RA3tjbPTZFKdTowGvF7epIuvd8N4XLZiT/srXJ14cahvjUskQgg3zm8t24
yFvY2bkBZ46DxYcoTvv6U8GfXMxhRWRg9zWKgUPJbV5hjcd7uIUHIzsU/Ot4
apBnSfEBajuUEze6vfU46RDj9fc556xumKByTpT7bdyEHnsBPgproAOHUKFm
c0Qg4umNpkN6Vhf334Z65+ZKTjALH6O4W18XXJhfQ6dH/a7gEIHxd/Y4jqI/
CF3aFr0MQURKJxyM30lcwhmj3MV+GIrgdoGzQUTmIGteqvCHKh+e9UcKoTPS
Gj4A4JrsLompgIo2JNV/EaKm6eY4nGs1YlsaU3XJKyaM4wHS/yHhhGo6z8vK
s7XRfoMbfce2s+F6qoyhOoxD65pwciy0YZ13UZrAjUmA7MlGY3eCHmBfb5k0
p+JtUmuWOHvUVhpJLdbu6f5BCIBiReqOqK3+Qaa/AfpS/OI9WiqgcCOUFQcp
r4EnTFc3lqR5dW8qrV59CCp9M7hrU2E73fIJZ4WycrFdYV3V/HftROKRh+1D
yWwMVX3Hk87rnEZw0ZvN1ocHiwNWFn8cwMIzcXXm1+dFA+cfApg8/zR3Pn9v
yaIHc4jSGyowUy1KPh22tj2DUo3fnaGkrLEeaxgNLvT2o8IcabcHyJom+2pi
9i9s+Wc5moa+mdc8r7xHtf5I/CIbr7byvtHZoI891gh5IBxKaddPEMB+t07o
tgxx1m8W0ye9Jj/+YIXZIGGLHo+9tNtgTd5/zjw0p4oqQ4D2/2C9FTyzTc69
CbtLvMnby6cZyGR1ioKwlTLAVRWYe7/AofR6CUHJATyRvY2z+4nvtxUdQYRn
lRkD0N1d3K2NdBxZdIEq/T/8mcI0UG9HSfUaYguQrzbJfh70vlRYPzuSYiPK
WCoF4GbGl+ghaZOxTZwo30MYxvmvbCVdvap5TngrmF2R4CmqRNUzqu0qH34H
GqplHx+wnfIemJvy/QSzgmochHV6EB+HRm0l1v3VXHvFDxU2ki8eGdE8J5//
9Our5WPkXbTKmuE/kwE2LnMEMowX16uKNcHOH6O80e384hnkYocHBAjPGD9y
NLf5a4WXV/1kF42l3H9HN3fXAYaYAYx5RNmiDr0UO+KPOLTj0Bsuopa41XUG
qquYRvnsUFnyFezDLMbgpdoyEQu+6riUHfQ8NGzqrBlBUYVkH37HHMeHWwnx
S75ggun3SV8nVGe5c0jqQAt2EONRuhmsllR86Z6QGhh62BN7ddSrEq4tgEb5
In8ribhK6f3cL1asJxxAYNyF1zUHguXaS5TktD2+ZAjmF3M7HBz8C0/+ltqm
czNY20H36leKqbAMxdiLM9KefCoe/ZMejZT2gy3JL5pMPLltjPKG3hhw8l0s
ubTBRU/jVEjiX2LAMt6zqpTYsUtxiiV/keV8kXIKmj7686SnMd3blLPyT/8T
wybsGx0TMlt664DvlatU64yl4QyRt6b2W01g4HlIjnW1a2Y6jasIi7jMRL1h
8UebNEqXCZXwPilk2w+IsGRv7ilI7f1vDQzjlBIz/fVhW8w7a9iK5YPnST9P
9ojjngQ2s0QLSax/wdxpVLikgg4ECN4j+ys5Gnc6NQx3ql2B2Zd60eNy9lHv
4Tu3SOYG0ieyMcxOOG+coJAcMM2mCYChb1BEMWPdRG3Hsfn/GPHaxofWFuOr
PKDuA3R3ijKXmJDV4R+MnWcykv1AGH7vO3h4w3QjxGFdjWq2Z2nvzO7S3f0Q
S4KI5/jj/cSbZiw1yhiiR/eJuXxJMSQ9qEn63EcaV/ujXqfe1RzWqqLz9coe
i2Y/Z7QfPmb2iPcIuXmGirgR4ioqqCC9wsmQrek2u3IR89RydD3adTHYFPZs
RHq4+pCUZAdP5co1zI6UR1pyGmjKiHueVC/KEYJsFpG1XhPv7nWK/i5EjByQ
8CfrrgyP1I8Y6/RliYtpx1PP+ZULB0+yDSslnbqSDQz123ANNciMJp/oPuYh
z+CuDE/rXaKg30PZsKaT8KTxiL+AMrH212JaTAa3UH1ZTsm+6zB8BH9j0Hm4
l+9fnQPTkwNMN1KikBV32uN8fJZXyOlcw+TWwrGApw1wzPiEwxaekP8VvsmS
93qVRbFO66HJdXgmgBBqGhOq62brw77VcNozVy+yZ2Iiyx5ynQ6pUbqD7biV
HZq0/D4+KByzbr935yn1kTE/WgUjI2QINffx5g72goC3MUsr41rQiudQjocx
I/pGe+xeeXta1WXsG8USLNP7YWhaFoSRIaMA9qpDBeGHJREi+x7KE6W7viJx
+VhTXCSdsPZiFkrCPlhvFrWECMetwYwE3RwmXHJdtwryWDQn6gm4zFzXSsQ8
o5oEWJ9G6lKlskl4jiYCVk2DqrsiEB6G4CshsAF/8sUjfZf3Ti7KibRyBxD5
LWlv4Wc0bUViHJqqDqp9Ddu+CBpLhwny9t24srd7+vWQVxcdY8NoFviphLVX
n4h6Z2HfzJOBz0kWfh1PSfV3LwnYHOkcVoAJK0qrVgwylLLJDn2mzpPbPmKw
7i2AsdBtgW4iZJ6cIW4qcKL5VrVwqYE+y5t9HRQDcNZzadcbsohfQsU3g3qL
vuKZ5V2CHofHwrFcU7Q2HlEf1AcKlxk53VCw0XY3rEbi/A9ThYlDq+SxB36E
4fHGHi3qBIQmZxF9Kt1nBls3eh4AgjrOTD/xti/fKr22SRqUlolUPXfOx+U8
vmAhI+oBKC3H+dav4C7mqolOUH+QW7r9KOnCGKmmEJ23jr+7i45zUeCfg4uq
lqIC9lvtXEYjK/CjMaDSTSHpooIX//slrMbryb4NNXd+coKm8CzEGoXsyIKK
ziO5AZp1UjG4zma0dGEK/KpKMKcFP7odrcepx4i0cxM33AOyawHI1YMxurQR
VtjX3Lm7QxRJ3SWUBzmz8Nk7SNuhyTDjQBA9++TLGIvqOqHEclhHt495Xy4j
GE349BUAtpo9m90V37e7d6OlvUQ7Zv1u0fQ4/FhkeQF9NxvStZpr4l44sjNI
NcgbMnKaGD1uwDnGCrL3oovAvLQDfrSyLXNoju0SsOIHZJvbeKvyd92qBuCh
XQ+Wkx2Yl0D65pNlqr+ejrY2gaIkXzVBNCreGzXjp9BTEzYNJsdrcX8wvQw+
p5KqQTWbZ5Dwn7Kc4uGur7FPvRC+Xk+KP5EJBIassurTroOpoznR1VAm+iJo
k9a7ErlhsImy4A293AiKk7dBhW4M3aLB5hylo268f1AhYvtQJ2EahivRlnyW
yutH4F5zsBRihzUWljx736n5c4o/qwKoGQ7YpHcf0U2vCVIjgXxqnGkLID0i
z3yWzSmUlfYjyaQtq9s6LLh3pwhH8xR2es8QYopHlz3hstsIlGM13DoWFH/Q
dEwW+c422mlegyFiD50gnNibhiuGqSBZ2y0JsZjaPO3TBtcb2r0Pf4QROHkf
Wm566gCWakveT7US2cKlMFUgCD1rRhTfSb+tuaoWkBtitKS6XoLh1yHYlYCC
a3zA0f6s84MzZgoYTatR/m78W3nysVGRCBiH1j3aDflx8xji3RIizecekTAp
BObYa6g/xcuPc9qBntf5H9kuHPmD2r0jL6i3yHE8AtO8QmS9C0/dK11zLMi9
/VkoXxI1kAfTVWftLX2/E/GF3Zu2YCbg+CXBsQU3MAH1w6roUrCbEprVXHxV
0QQhD8NnH+U1VA/bKaV2hR6FUUrWx6/0b4xwork7kh2Vuhl9YNdId9SRGa9c
TcqIIwgFhhWksXK5w/DvQW1LQ+CrFj8dv725jmHg5J03vj6prJtn2c/Bseb4
WpBpZ4PVq6PpTVi/kIw5WrlYLL3FlGG1BfOh7Kz6gcUbPHfk6IYG3t9ZHM7j
QQQjS2/46mdx9DHOUvTr9WyRlaBdFB20wGQKxMWN+H4JpY6pAsY7Gh+WPaz5
M3hOEyBSBrsu18iNedCAtx3NdjYn4mIJ+aZ9IAJqH2tymPj8QqJznToBx9Kp
Aq2bbWcKLpHHI9le+W/flzww43ap9YvvcznfttqsXKYxJjKCE6ILPfnT4q4G
AADwQN54o+JQwtF15L5tugEGenW7xP7ZViAwwqdEyu6lLrar263n3pNqyXdH
fyiNRP07QePMFGT+Ymg0pcL0ZAYw/mRvShMqll26LXzNZ705C93alfbXSHi7
OD7NL8vCrK2ntJxiUh0GalFE6kNbI2wf0MdJyi5VOXuyR1YGdeRIEnSksy9m
7oORpsqPOGD6v9W0HkG7eRPIIQrjD/bksPn6mM++H/5UNA+17ZGnM9dLJ3VQ
1c22yEckJdaAZ/Mtid3HV8rFbctVZQ5187W+brf6Y8de7T8IiIViY3xD6o+f
NFswiIqcAHKGF+p5FqgKROuzA4O3nj88w9rdWhZBbUWyhdNV9nbhM+eBV7Xc
H7xmam0OzgNGPGFeRRo4TuMADxQdBcGzs6iO9RkDSZJlHJPiHtRBIeDdIUm6
QSx5Bo941yL4n4Tls1+4sodF6X8Na/yypstGD2K3efO/Z8sc/CoooqCEolXW
sNmrCcmrXHboQNF+ENoNZSCX/NTnCA+qG8yB9hlVNNoPvtXf3nzEKv/8QpjJ
Ym0+/YFC3eUOqz5QC3PUGADVOK5NGHHgzOtmu8syeQeiKev/M7tL7r1qBdOU
WQagalgms1mxIy8WgKbXrgyVlIbcZAklv3iKM6j1/U2M5x6U4ZLnS1Zj8AAc
Ssooop3G0/SmTMTNhZkTP06TE3JP1olTXIKSSgaQay6SDyZC8E6QDuK0ExXT
h0zYFcihOefd9wIpgFa21qtP0+pVp+aT8PhuOJtCs3Ut1SAsyU8OvOie/Xdq
YsAIMKw55B7oIKT1oE8G5eLI9ZJyxh/qk/WQSF+qKGYz7KDjbcei9Q+o9rnQ
W0k6dM/pvHIowJykQHT7pp6GzZU125TF7ADyMLMvZ2VqiaSUwSdqqClkGbDZ
dyo/HATVJ+A1rPKfbOVPfHEqNxQfjUL9cCUEnPJ7TVu0k/wBNXevQrORS1Su
8VTZnktEYaxDD8VD9pQ41W3uhQvwiU7RtFthljG4seVJDOj3BbfCCcMDmaEe
d2ZrCxpE4ndxAA5J4FgW0gPcdSF/AYR5iPR3UPG4Z0kZo7sdnb7OviaqVu/I
+EYckIp+ULizJmHOHzIKtDP+d8IfC0ZBd2kMXqhAOwqP/OnusAyNP1rfTqtj
gKTUnapkqQMO4no8wdUfNkASfhEAzZDaKWSQqe9H9VbEpRKAvRer94UhWn0Z
SLS4bXNWRoenTaixRfw0iAXKFG4DFweXgFBIDbxouX5lisEjH0+26zUrj3M5
eClA+25/JO1hHHfBwmY8/aoAIsL1baLXWkH6QwsIHgEh+F0STobBbhksupG9
gpoo0xlkCSGs+HCbHRttImcOM3fpdSAHjSZmJhpWxQVwn1d6E5htJOYwXExc
s3cIIwX6F85Izf8omoCQShueldogUzO/7MfZso1aqq8VlYjd9rA3dQ0sBLKM
Qbr/WfFg1gnBhD/P6WXuJSrpVrcX8KKgkECJsmWCNR2DWhxe8Gh4i+fwEdUI
Q+X6ysKD4jcsZsOtII7Jyk1eHSpcC3cZKz3mrMd/S+SEeSBuMr2AJFOalAm4
VBKfKdrBU/hTfA9/skzHln5TGBkVi9CrmdfRG1qLeS+Gf6B4reFjA6R+ENgm
y3wo5WBdD7hAShU9hyWdjqDoI+G/sRCtNb/vjpJfa5vBfyJRsIFMdFd8ye23
JE1tzy3FCVFZ5GxNbpDzDD9YRazwIg0ywmV/ccmEElUqlrQJYJCUUS/CEHRk
+uwr+rGfcAlkEy5Jkzfc/5j2+p7zrq2BWy7oBoViaBi3/TnLqon5MbvY7w6W
1U7ZAe0d7m5SFb4ZcFZik1s+7v939MVYFS+KT4neYOym7qXeBDY3tpdRp7cg
LJmyHvcRYXdylKf9ScJgrCSAizl3Mw4U4DvqWpVoCDtxiawVi6Wsgqz06iap
991XQbm7+U0fVs1gNA3FPF9F7WS4jfmY7ozAJkKbquSurE+9bwVigCpkDR9M
EETDhZHOG5LaKSomBR91gyqTOJhzdTB1aLAUgJDlxbhG32KF276XG/dwsVUv
bRkLrV7oyYGxagpC5FvoAza22+H4DAMhrXQ9hSCr6/Ulo/WcD1frK0qycA/K
VF5zTBdDf9yzYZVx62C01guopsKi4MF4aXtCWxfMXqIRMqfnXVP/0n+iciYa
JTstWKwt2Oz1hcgiiPdCac23Fpzk/5/0tJwlbFSD66kjbRqIc7CAJQX9sC1c
fRkiIzOyUa55molHaV1rIrIxe7N3hcW6CYbdYMN24KGBvzIvQiOdaDLDxqqb
EDwBAlCQMqGCwyeFuDAXmEbwFOu0xaD/M3f7iyMI+tAzFnS3o/RyH+jtOPkM
ROXIh/zbgRrqRc0ZF1bTMYb+dCAWaoxUAl4I+LKG1Y4fwU85MKc6Ilx1nJlq
VI6KlvrMQKNv6BP2CNOVXKM3PWR/UGmClUIRMHHHuShi1EbbYxh4hTrpCmxT
1Akqk7H6jpE4lKGUqQrOBgx7ej1vLyXoUieJEM/7MxnBsj9itHhLcrUTnhOU
SQPKQ3PtuW1tXh+aroP4Gq7k0jDihzLq6/Y9Xcd2P8aR+2RVjkWU6OOAb6Gd
Du0o4BaiVvhmNtwAfLtNZbYRcHYHNNH82WvuVJffy5fp6FTrVz73SOrCU3jX
5dzb5vvhGrItY1gakdh1qrSMiaBpx19EtU0Zj0rp7da4zKwewxESyIpbd23k
oV6fh2Ka41J9mOehao5SO6I6lTaQ5SHyWYy+j3xyQDk6+Wx4745YB6fNdI8v
zjEQEPQ68/6U+LQY2amP6E5lmJ0IfZkZlFELS29tZNCfzJNLp/PTXSW0eNUP
ip/lv8SrhnOV7WvIoFir2jHwjjfQkQOsW2jIOheW1e+6zCe7EVaPzb8DqA+w
FzBBdQFMIPyF/nQvpo+YM081P0s2tTPT1T82LWZpGrS0p0O7p2VBjtSJWWHG
QZK39OjV0t8dxbd0N2zmRM+JZQmn4GCEk+L5OYtip2nuNWQkKmU5LPTz8TTu
rgFS4njikJrEtdgDpJ8swk2PViqiAuRsjIDlT3ktfI/ZYKF8M3F838XyoQgr
rxVLOa/X9duMjwg0pK4fpvyN/sFEqEDmM1KzNJjd/KBu5D7aOu9KvHWf8/dc
TvEtKoYdModTbkcyoWGVYTlizgyOVWYT68fLCMVpQ6CNwGFE+V3jFsGJ7/Rj
htfP9oRdwjzhXk5tXgMXCcjyf3/n1h3uERon5huvp0IkzSk4+FJ6awzgWaAm
Pa/TfVSqbAVtXnOhuVTrkso4hjIDPC9dH1YvmqTdnYbACWDVdd8RZDHzpRoX
cXBs4X+x7CTN7xoDzNHUr5OI8puLwiPrymHmaW+jOWOF7HjpShRybHx+n2HD
dgyHaLdRpdMDfACqeNKpeJa6gQTWjLIFiz7gB/CgnNkFsppEq6geCzxhEDXZ
7WMk3tJfhNHFT2Y2I1U/zcmeL5x2uGQlIylVUABoi+7lFVu4YqaRo17Z8mDW
nzLgZYE4+A9c8jkroBDZazjqrXGVJNHvHEWr7nxlQbDWEiSFsMu/uStDaC9T
oThQiqTmJ0mn++spc5N6gncFlCu+K55gn9+vqpnBOg/vsHYDsx/FxMCdUmhj
pCGxw2qHPhAMuXIq5TGH9KSsokUJr0nWOeItf7CnYdhkauryYkA+iCtYl7oH
EtlYAN1V6Ud1x9Wq7ysDS7mxN7lIwDmDKhIIYEavosi2+3CPwmk91P4kaGNQ
K8GGHXiKsnwLLdXh5rCKm550whxY7MY+VTRZAcS8NNWD0HO40xRKvTRIbuvm
oNeK+nCNHC5LD8fNpNl071SG0TUoU39legU3n/V1Q/1WSeumzf+atBTXX9yZ
00IaW1ov+KxbJehTTPO+HyDTKta50pCFve1PPvuVR6yMHeWdgnkqQvwDV5vf
YFeHU3oHzjSCHo1S/CQgKTv88IFMz8nJ3E/4gHlNDwL7aApAPu8WRNqtArVy
oRY2kw7VBT/m1TFFyt2NILrYW6J5EMa7JTpKivx1U/QXtR0nMGtiyxmSkJF+
A/gH4BKDPSIEiSt/XyO0IVNWr3HHM3EAPCee50ssqwgJt2mPR2qTEv9PAdcr
Qfj6OBB71kkDyD2rgZVg+UUgCLgXBN+yDjF5kM4tS4A2kVzmYv+duhqfStEc
YXclr4nK9iwDzoLTajVxdcA2ob/LlWxoU/iuHguBVVmRM0hYEg6iASYTgmbm
QBBp4q4LMqtVkaozgETGZsoX0qSiFelyBfmdK+umfsbwUGry3GYf19GtdmDM
wGEhRZhk2SQssg2c07P39sUgyQX+oAP4gXuMq3upSmpVKpHFR3nTTYz5/OZ/
Liz6rJOOlDYdODwxBdZZmsv3asyovvsXTNSMGjMWvzuoujDKAwoKZHifp06h
qpnPVzcOZWCGuf53YZhXWyufGjESEBux+V2T3POO4P/MeX0rs1eOYteb7JDf
3RN+YFfVY8kFO9qqAB/Sq4U+8p8IkikEOEwkiBm3aDmHwtJZtj7jw+vHEZMK
YbKaK9fXPg1bsECOAC97ILgOXEOjsPeY8VmgfcwfiYXnNVfjRLc9+uyGu0kq
tT+hwbLVLfg1NyIAOGJuCATGLUnUuqfwr39Sp1w1X2LaCp143HHnvbGJW94W
detGsw1v/bb36UOdrKXMjrNagvttsqwml4CJXveqC2ckvz7hL375HovmjzWv
DvKAjnfm+MJuaKWhc3ADP5IUkQP3k5P6Y1S88up+jlQyGS1ZFA3D2nyCvJBd
nha9e/qzla68Pn26kWOMW0UNluh6oneOll07uLvvEO/0y/eWNVvGkef1xY2D
TfXmMoW2EzFKsTtsXFsJtJIw3a5m6xQfZZofndNLnZQcEyON9kim6RhvdYQI
ehK0cXLzfCt/cuy6u5UtLBfwAMXJ95DyojpYr9tbWoZFyDOkCJAOUyvGUkTh
5wtrlcM6rxprohISn4PadhUO4E17y+r53CiXnGeuaLlnpMm7Aw+FwVwXW1G+
7jDVFi3lL3ps13diFpLO8tY8zYuC2mNke9S3PAG5eae/DPJtmMOx4YAIapms
WuRx1/8utCvQwxtU2KLOpyC/KwRHO8kevG1Hqilf2IrMkLaopycMJUv6moQ1
TN/eHFCYgnJc3gNZzo27Q0UFWnwf9zd6T16mxWFUrrgrLxyUXf9errdu7jKX
i8EaOXrX7D96gfgiUoINZHJc3WCLEG+ocacVYXpbXwuilHxCB6zXc0J8olti
qhVFOVVLxN6QMlKvpR9dWC5qS1rUi8yKs9w/hDRYfTw7BqwBuKB7hHL7rncz
w6fF1K/M5AE8cNBxFuEENvArv7CSSgh8i7A7pmikWdLyYFQEyh8gI3+i7Skd
PaKSedh92s0nv+VNlzbvNjoyvrhtZLRNJ9G7oNny3Ja7qV/v+xU6dFvzhcOt
gp0gKGDasHzrEnItZ04eWjRE9rlx6ETqRbWxWHrWjiDRpCmZVtoqGtp1BrvU
V2wRgvVVOKzICmrbDcjiJUIWFnuANe1Ze+0HMoTaZJ3DHvsqV07ELshDPWhz
wt5FLHufcI4KL03EH+j9OyaBrkuTl4DHqPXXDhW1ap0rbmYPhdy9el2p4b1N
YTEVfn8B8m3SBJva7hhkvTRtYOslnrO+VEXIr5X3MUm38GWV+zMo++I0Afc6
XnpCpHANgUXGeIBUb0I+cmb1WIXlt7ulvI7F5s/MNFd/Tw+cqFtr6x27AQwz
54jEIheXJAnNIW2kfb1qDfmnr+LUVGP+bj33KGc9uiCZiUApCSOUn8cEYKsw
BQynn/pY4N+fQXM90rwU38BtnlUwyKQwumPMrLazP/1v3EvZTyDwKB81KQSI
20GyRgrxp/Qflp70J2mSke1ORHnn1lWLNjdJ9T7oCTK2HHBLiLKqCi5ReClc
yvEesZeH/rvfQsyLtnjowI5ZouMXD6krVieJ6NZ499lf4GZc4S2zjQcnB2RI
IAe24wFwuY3g+ZcUVkupvCKH8rWLgkeHyO4eQWHJVok2/Oo+Nj738mygvnbp
rba3yMnm5Xh69KCPkGW/cuP7W9TWYZ8jooudof4+AIhKSUF0xPXh2gObjGAz
f0AxHUdYS6uh/R8qooS6nsJaLapP9oflNlepLaXpva1+P91WyC29gc0QzjpY
WYN0YwYTr7aTRS3MfcOHcr45ld0MbFmrivHAyuYi2AyQ5fahRDF2tkqH9WpN
sBomWv9bFBqPXZN6G9iHc2OEiEnt2tz2yTnt1HoLB+dh6it8AdqV8Btb7n9L
TcgN7AnjraWJlv4nfMLXfuPWqw94t/oD4tpczhtGMDWeGcwk6FUEf/evdT1u
/Fgfago23raYrfNZg0jTwlibEJQ05K73C5qLMg6aer9d+crUegaKwTQ9LjoX
uU8dCsHrcGvkl+JZBAjbrm+F3LO4ZGqYyoOIqY+b9hZQuKznHmXAxhwIR2d7
P5FjFdg5d7d7hmhlQd5RSer0cBjnp8wXQS+mOtC9ZWoXUjdR63vb5bQf28rS
vCHkBQ8vxuRlnKH8WJCgQebUKI+2dgqCdXXibzeEz3CkmEL949rYprI9Z4ov
S20o4gRF/9Cc3cfmEf/jQXgYMyZ9A0xKVaTL4ZDoWXJgAWEPhGMtLB8RNkN1
J/0tPoxqgXq+BDZRMY9sohPFID+0CNCqvVnJS+y3dCyxqZjJZbCuWW40JTuh
awVMvmcGV9jwqNK8NDsSZyMlbcHdJdBzqPKdyzAMaXXp3E8jxxL/cfew7oPV
ZPRpD5XvKq091qxSDBmK3H4bgLjzjFwVICvkDTagXRW2UkDhjVBv65Ymt8ap
RgdPkRa8TMTN1YhTqL+s8RlhKsxMAITKttvYb7wyBBceBcgKhtq333P8hElH
hiPDQ9RAuIg8tlGObjQt5DZF9DCi/3IGYisvsFXqXJFHRaL2MmfplJchPG06
HPj0SjMKier+ecopk6e7KvdX2c88XLU0vfdrdgctCkhcNMMnpJB4e4vRhAF+
lz2liB/rqw5z5f6nEgtHiSVsmWICp7j9QuDSbGjsOkzvPaIfkHFo/eVYXEf6
ETSmXTM8yh856jvFY1W7G+BiFJlsjZ2hKr8ZYsPTeDsGJGTKBaVIlJSqCD0G
iARAzL9qKiAYLvXG5BD1bLdhPxN/WivN89VBD7b3YfM+mIzYXDwC7EYWlXq2
X5zJXgIqPlgQwGHlSIJFWWSoefVMd2Vr4t8VI9yD/ClZkkjogvY3VCOFXUti
/Jw8calhmB0O/s5tynbPwsFneX5W+RuOXygeym/lYBaUZUn9wLSa/YStZmIJ
uhZ1IGJq2n1KG1+KuqEOEYyQT1SZmoxkg18GUWahD6Vh7hYv85M06Db20HXR
qRwEoDsmIH9PfpDJkROyWk2YKP1yogdFimVLGiTKJ1uK8/t8AjPqYAaIq7VQ
boGdr9scR+EkuIvuqEyP3ek7OmcnM/00BvpYGGvU0z1JiFL9SHAMzafM88G0
xRW4t6F7ll3ouexeVJt9KjQWYnXVBQtJqsLpnBjz2ZcL/Y4CbsnfnsVQtzPl
++jYP9081tdA31mPB7bfG4Q79ph0c4DT9U2nw+0yGa7FvsZOaDscuC+4Jixd
9TgvrJtybTYbmty8gMLQJwvT64OR9g5rPKVvKkNqLpZPHx44BBag0nz6pXQB
ocvKDy966JSb1UrKiWcW7VqXTF0bVIe2gUueAhxFD8thU2kQd/sJi3yp+fmY
Uwhp6Zy9cFDMpXlpXNsjvkctOrnx7ot8sKyVFmVVcARfVyXzXXtBjGrZJsjw
mKeQ1P7Ld5SRjior03WShoNz7QTHA9m5iJ7bsO2KNtAMSMu2lHFnR/o+1hYM
HOeIsUOjjDGL09wSbpunYLFeowstRDUmprRsPXjofDOqODEMUdVeXTQE8+z3
W+w5rsevFdQJd9bbc/jt3YJ9RVFva/glWBrpoxRFO83g/quCtp4gfCt/v9fu
Zn7vSpY5DCNg3Mp1FqwVeq8GkQVS3AUqLqjtRBYNE1wljBzf2oGcs/9+S5K/
ixFWeHPbGm3DsFFjmdsXAEM/ITLk8S81ebGDIyxInT7WSyQne8dt2IU1Ilrf
Pjwtfxq7kSM7g+hSKlr7EEtD10DXBxUClwNlE8Nr7xC/Vwf50sMGr084P5UX
AQED9O84m3ZQUsDgCACf++7TWFCrBDqKroYFLXAGt+jWVokCZibhXJT9d5eo
6ixUhYZ69LKN/eQfi60ORE4rYZAu1YmHx1wLsdvFKAafgt3sEh8VxGp8dNHJ
QSSYFnzwkCN1Q+jnzGAi7toLD/tyxqyTqFD2HlqO+4CMkQCEGVpYLcfRiWBz
22acZo3G/5NFirH9L/M+oPwaPtYmQGI+vMK1seJCIqiUiSymHd7qXyrxWtSp
p0HRzo38b6cbM1u+FdbH7dXK4BQssylukknemq56nf5NKDqZoMHkUm6u6Vd6
8u0ULr7kysZzwAw5QyvAkrb15At89zXn55bHMddM5AiBiOeN26GYfJ50Gxhp
9sZXa93g8skdeWBfr2gqcORvIgCNNIZwPe/X0jMjAE/ifpsLCDKerUFcjq9h
kwa6EJ9dvMd4uWVuhqhcpsZ5YbtZqBgEBALZie2ieA28R4BmUvhBHBFHIh7q
DvrgWuplEyMOusTjkx+4ITjeBx9v4h5oeNdvAM+3BhgL77+M1i6SZR/I1uPI
JDtdtSl21YAgKRaCgSDtvaz4eULXMsrA4OhFp9BM/vb8b4qQB9TqL5nzQh9i
EyQw/yANqeqAPpf/OhNbnAklT8c1csLCscjoSvpn46HJm+IDi/yKxaXgSNsa
BBGyYZ6uEG8KmtiZHRIu4ltsMxNAfZC0m9LurJgmaWYYWme9EreVKqaN1BWb
g/7pA5ekW5cdAJdbx8NkLZsVOwJG+5mjAgKIwm4E+1wuOeiD688wNrUiH45f
BCfp0EfBEbdOTF/V03hllFIa3gq2mPlw1DZC+8y4ktmEZgAu3O+NtZ17YZWS
1b0dNsG4tt35maPs3sTxm3VX9nWdXzp5R2kSEO+lV+m09r1qs9j/SOsJnNvw
eDeoiRJa3fTQaS7G6uv58gmv+DOUIPnopYJw6cGlOTfR66X5HtoqIrvOeZwt
zoZQKDClzO35wQhyjTejuX0HbRyCuUh8KZ0QKBMTeMVzyey2rlgP/Tk4fvFA
3jRH8HWv8FgmIkKdEHHb/tGknXPLfMnu9XACY3ADnp5UPIWVZtFE75oZ/qQW
m5AWKJPZZWguIxvsE2G2jiKGT+tMstIeMZ+yGofYaUjiyHfuipdbbhCBF1B9
nCk3HO1w4r/Wsmft8Vhbx4sDiYF6N9yqPs1OkHHKh1Tjarq0yW4VGvPbxVcH
OI96wo38Ay7mkqLASwNAPX0Z+/2XtAE3UqDEN4xEMLnd8z8Ej8KP7VK/g0M6
OdB3PT0ZNanIa37tWh6Q8zII4+N0JJbKkxPeR7ISjkit5EUB8WyPo1Qkx6bZ
l1MclPnvUL+cMB7isOPU9IjTXePcaWhxuGCzzcRGl4TlPsNpbcq22nFq4yKs
S/47HiIAntasY0NfMt3BWilD47A9bNL5t/pnU40XkFV0Z6e9Q4sFww4fUkQO
YXenCqjm9z2xASEiIICRcnxW9Mwh9qmk5mrGZFzFOheTaMXyBnWSHwzJbZuX
zqO9NsYJq1ti41UxaI3sfu4ktbss+eTZx80/Ma4ZOZDQwpxxNc573jGUllR5
c3qpEgkdM1rpcAjztCneKUS9G3hY3TCqsMaZf8A5jZaeTunDFnhWG3n5lATr
/xl6M4Jyk0blkN/ClzPNXy272oTu4DY7is5pfK1WnXPn7mmkH4CaYXRslxMt
99dpGEsHtBb5zEHf1+ki0LGObBbghPElK3FeF3pUXfazxtCVQVky8lTi4Mxe
PeKZ2A7vANW+1LX44d0tbw7bEulW5XWUIhLbcS0aYxkOWDLdGQ8qkFA4+NSY
HAN5BtKQI9b6TutTuiaIdLacemjlYd9Ozpr97cFS/N++g/Musspj5msRxJhb
mP+twClKl2G0ndQofVrzBcyCJg3GLQVtHSyxE3nyyI2cq4aAwlpkvOvKkSKZ
rMIz6RBCJ9k3VbPmgKTelLNLaj8/+37/Z2WS7medvU7UiD4K4n2G0LKIMEck
b+oJzdiT+SncySpBzQBtCUO1IEql1wawvSPqBC+9XUozUcsRtO+SIQjqIcqB
K1bJHo9eQJzFzM2r9AnliZa7LjxbMUoWxKaIYEd5ez8zRiXv5fkPvjjwDUy4
ecWPfEm0u0Y/xEx4AoxRmiXaqqI/1e8hgtPJSFiBBLZogDPSLG/fBXt8h5FS
04EStmmG2CFEg2mS24HZTebUJYy8m81zGrp8khWGMb2oNy8ANrTWVYLJnZRK
X7iBydTwVua/OLJ5B8kx01EuTndbVLHBsqNiy7HCWGYTgD20/kocGcLk/+JF
ySHM9pWJ39gckQSg3Erdx1iNUibLggQy6swpwvKMFol0A/LNrwWcEwIrFKrk
/eMnZj8Mplcz0bbQ1sAOHUFJWiqpQpXbjLocYRhFzW5/pykieo4I0iQYefaH
tXykVhznQ1AnNLk12Q9n7BpATVqTAfgnkeeLYJVziKis8jt1m7OuZakn4ano
lK9MERPb8uKIcUNtUptz1Gg+x0wVOqB9GpIySBEHT7gRf88u1JpuJK6JYT2w
57Uqk19epnQFSXcDbNV6LeZNXBteSyS2lCY+PQ7hgzc/gas8KyhEoYR0ddwi
xg8CZ+yEHZfqayuZ76EeW6SJ9WWhQDXZN3r+W4UDfCJ+Y19m0x/JndeArUUB
SrqQJhG4q+PtAmA+A5HkY/s8P+SH/4EQG5pwoAUuEXXaxjiMHoxCrm/GVI1x
X+2TDqRKVWVCMZz4g0AlT3fpPLPTne1HpZsjWOXDeZm3G23XLNTDWBVugW2v
QQuFtjDQ1G8eYGwkw96nHmnjO6tBGRZKsYUtFBwNaPXvIdv/iP0Wxffb+mQs
95PrB8S35nmXw4RVi6bKlrzf1PB1RyWnoQc2VYXMYamvD60IcfIOSQyyBWMn
gvoPBxHeeVOmz7SxG7cWjslxfv3ZHnaLu+ttGT9r4MkyLSxC4BMex/zfydUF
wc/t5HKV2fWSIMqUNKuDqBpu2SoENC4RYV0x8V+rZZYAqWpsSaqJCARNFZ6c
w1tE8mIlO1wLxb5X+xmMQZNVkwJlBw5eRY5HJFl1kC8vDNQdpp0NMjowY2gN
haVM33Jtc4+Se7mFAS/ulA8o/kP+UQEu0Fc+0JPkr3uaOcSvFCxG5gZhNCwG
nxQuP2dSY5+itAFFehgK8rXU4PcRzyftP4g38YcBY1KHhLXQBVawlgccsZoz
tE2anLH2pUGs/HhsX0boN0NOa8C8jrqNLjq/XPUAjMhKwOnTQY5hdK/vf3N6
uk1o6A3gfNN5NY/RWka/qA+wuvrpf5KSCA4JokO9gWIlOdGsUFO4J0pc++b9
63oCDKKMH3z1J/WEPM4W2UcIy035K2yxE27Luu5DTKN/mgldFqWJutmV+pdp
lvTodSutdQ2bHkuFXOxaeE9YPYXPMehhkjPtaNpLMXfes0I99jpjTsAlxL66
MNwrxVMiBVaxPBmSDJtWz9Y1wytYnEUTXiY98D6A+LLJtgC9BgWqE6+X7fGb
L3yCxgNoSQS4LWJ7Z5LgrbqBO0g+TKqc+ObYES1q7vCHVOx6y8DBJU8a/NBN
jZGIxmcU08TfauG+99YUgoc6opCL5TxZgc2MICmRA5+50UCKnhYviKS4gV9W
/C8ULGOmtVYjnlhjYBRqDZb6zjJKpLAiwdNpN+vrb2ig7tVHYm9paZ2D9kSw
D/BQzKGjAg6Km50iGmfRpmdj71+xJrwiCRnm2X9effO2l+ggS3cBpWRa7ET9
YsgvqPIs4ZZDzSH4IHeE8MukXrJTpUGg0Mnnx27bKOgZjdLdSzgF1S5MUIVU
KQXO4901ATikEfPOpctEZNqJiQo5nGqRNVWgHZCPdyaD6qtL8Ok4FdziJ8Fl
MSAUKiQlSsJjditRggESZyJ4RGYh7Vq1k79nphXualR7MP5aXFeM5UCUYupm
VfoXs4zqxyeKWYI8jIrSUaRUOOiQG+KJg+Xwf+hAj+9N+l5lkytudXhxC2xb
HoqkpBnh7qrtoHDMxV0NXfu9aKt2cZYM8pDXUGnsxazXvEEef8fGASLYn9L4
5WM2qgAtsGKpSIQfTyJAC1wvU9JHrQeeKnEd9GqHN+DDYd+3Vk65pzGwMZPQ
DHkFcwsAkHZFL6HZV9RoPzBiJUYaGWjaK3yLZ/jaaZ2wTa4CchUh6yVk7ewK
lEEupe0zBO0Yba+6desIzXHlw2ivKmbBosjv9xtMg9rRiq5iNvPa3h8IzBRz
UIuTcUxnOaarGKC7ZH2Op2xlHm/IXlwx4faH/RdavnDXgIsKs9RUCqh/tlyO
V2nOmWoxSGNo0f5GCrxJhmS2TL2t8zEmClH0rP8tppjEqyBifGqTAYby+Tib
BY3EQK7/oqqUjOvxrShEfR28WL6dH86WrEI7IzW0xSvaftbBzZGM6NU+MdQg
ibU1rqNt8dWbu+7eL2SAV9w6Lg/O8Vot7UJewuH/yCT4F2H2rdFDlqpRHbR4
5Esfol/f1XlsRdroyvLTmYp9x7bjtUDTMvmKKsYFpJWM9uArPE2fqoCqk3IJ
WJiAapYFLhHrp41C9dDX9j2+QLOOKBey+TLEjMfuMBs8YXGj6mq55KfWuelN
+jKDLBGqLIimjuKaBWY23OBdw9tiSdmoufUggU4a09yucX6F+2ngPJsczzNw
vWBH2IsNmldHt8k/SKEYFVtehl/11xZOfalaOYdAZzkh6I97tz4RpHB66kgv
KxhN1ftZR5ogcTqUjIUR/b7xjSESA9TRHIYhEmCErtGyOQmXRwBFsH5e0epy
CBLuaQpFTzFAjFGOTwvCal6/yUfl14qJ2+Has5uIaMGHfpbU6bDIsCwkoymG
U525ZFXwzd4z9uYSPLgyhzclqm14UBmPsrx45IVvUrsTDml6uXtE4pwI4+TV
fEQtfMSoAHzIaq5Gl28H7dn16reSQAvJ89kcABcYFAVFOE2SeobEfkaeOHpM
89JipRu+s9ndJ0HKG20iybPP5lpqQFdGXLyHmVWeebRjXYxXNHnzZp8daPUL
1mSBt5ee4w2egMOIUXVRIK4QPxFb9r8YuuiOqYRvrb2JP4IPmp0SR1khK/nM
9vfFEJC704LiVDKb32djazufcKaEQ8RjkA6anKeJv8QoT45e2XMTPgG72X6w
HeH1cw6lNFnzzFV9iYNCuts2Du3ROkE6JaYObAlE6DHMs/7G3We8tXOmAw8v
weoLVsVwhXQCukZI1m5ljfap5hbWeugMAnEzvMZyHqXYVdVR0A1ZeGx2pWzD
4o2bQvDchAGOM+ldZq4GavJIWN6yAKMdCwjFlGDLvW9+EGcpPvEikT++QHzM
RnyRLX1kTibh9pTgCoD6fCUaGfC7tK08A/KmhVfwHCgL812AQ78hhREiMiLn
57U2itJWh5CdLIzTd6i1Yuk8IYMp36V/OLnpQxJXhCxxjT+wwMElUQPKlXpe
Qm3CiD4FfD5D5nA0+4DRPoTY8EtGUMgVCNku/u5BcsGJlRgznqQxskBlZ3ql
IaSMREhDCPwozim6NZPXIuLwLItPO8k1tBY0Y1W4mQazWAg3z7Tq8bb8tOHH
tarlAESh8xGMPk8xFnjQbOeJflT6v6ZYehAFC/9zxlJFT6nqIi8L3AI0tY/s
d0d8jorpVSo+x/uKbA0H43oiLvuAV4hmhRbHvMqvMyD1idJFyuGmjsVncSGc
4OJSK31/ZmH+jfJoTBubf81Kdg4PpcLCVDE9rDd/CGY3p5odNR+3C5epjk9T
OdEP8JelhrLtf055otGeDGZR+N8v0rbM9gRYxpvHRNLlbDd0+sTXWz3k1EBw
5QrxHfKEzOnLUNpQeoWzcnUHeOcmdhoC4gNxqY8nTyibWMqo7/LEkWAHIl4b
gSFCFHoAevj6Dt7pZhF7UFUzw5u4Q7IwQUbZUscgJkKYBMp784SwzFxxjtho
QE2KAm6qUY5Xdp3K3ZM/HVQ+7FsyZ5dPmsWGs9zxGI/Q0rSOVn4vNjseDp0y
FbpGaan9h0HEX7kmxSYMIaJGsvfUWECxrOvuFDiG64TDxJwYlfks5qTICtCD
iJbglPAwIBhoGIMAXLN5BaHdE3FkifFkFigq0daDH00HykbqkZpNrqSILUaU
63I0SWXR8BWaL231mkiWzSfYhhUDShre/fpu4nkMs/58bzXe+iVrRWwsP75J
5Y/sGL4DEwTs32Ptm4xRVxPhlboV7zSdBsDrEc/5KsEMtv2f0xZPnE3veTiR
VZEgi10EOJOSr0PpuOLXZR4cnlXXy5K+YeF/To/dctNaFZpPa1Hzs4lwv+XM
fbFslNONpa1rjJrt1rLnGUzVUW1Foqx/5SSXGrQ9SOul8yDDLDigl0Ireybx
q5lK8zsWgg8M+P3A2/Z4kjST0DoOWN+4MjxxiMnx0eeSmtMBdOB/scFK5V7a
ElhdLgo01XBO9ta9eZ5QKAVEox4vQdrI7guiwIkkn0dnivyReMh0AT5ZC+YB
CfoUnTeZ6MXWDFB0mLMlc6CQDApawxOcO1mmpzeOksGUhed0HSsjK7X4jGtE
cXZs4bfQvCTHPJaKXRUvsTgUC761o1qJSD2Ibjs5xolJwH+E37mc076tgP9t
efFsSpcfRqbs7A0Os0y9nGvROYU0tfZPdUK76kWTdNrtxNBjYmQOH11QxFQ9
/ap4faMaK07YiSqEYLfI1YExhx4wtKfrEOVbW9ENT67QwiWz0T7yguRhDZx9
AZOgg3kryh+6HoYuA3FLacat/KPNgbNYbGfmQj0pQdYL3EUexW/zS8GMlcRN
oL5F//yBXgAJB8VCR0hX4A8LnRUp+aSm+COo05wpyvDPtr372EeYlGcOsnVX
WoxqIHP30JQWRgNrRQ0v1MtX7u1XSOuuU81hDIU7Waok6vZRimhc7sKPT/+v
f2EESo6db82uG4sfD8K5lCPof157+cICi2+DY2ytYfEfemmhV/SbXleKPVU9
cxoQ0+EsSrnaXhXzZBo7sAHojocO+tIiZU4wakMpAoBSdn/mkl4/xRWGvoxm
8kAZWQXtmX1L2kYOuktQYwY/Zkv5eo7aQu8his85gIskpbzyI9bK/fzlvJ/Y
4wa488BrOU5SoSj/36TFSAKhrESc05RrRl4WD0zi9UCgMfwmosQLNrHJtRv3
T2TpP3kgJ653am5m7IDmH0JjTYrf8yZ3F2gE1wfU4fcuzO6ZPN12u0PmYyCQ
JmFzy8IZsChFedlKorwwUTUfDJJE1/kdfTfa2tnX/Kj6BcPRzMTV9xLpUtkr
mzGYKfJLpZuWaWlFhufqi93g16jVjpU3AaYBtazVHVH35uH4ffu9KMpTdteK
i1LflRk1OYI8TA9q0tcKZn9xVeMWoe52vw9U8vAdTi6C9zMPkLSeE2LBOR92
LF50AreGsN6qX1OdbxObUKR2dy1cAefnqR6QIoGE2Rm4cpRSslDy01B6HCae
5h7bwgsrwaJAW/ZgJY1D/5/aC/brJ8HPleZ6AKJ/oX7K5AJbPJfRBB4IJcrz
X5x7ZxRUcQUMCwIAuf37ks0gW7ziJWpxgsXe6rp92sgDzzgs6SzTxkqmGc/V
Ou3qVyTYP1mj+yEeYoJKQ/q3Bp25JUIj7cNfmZCNIG2lRGD++zKnCSrMYnJ4
t5SXDnNGJ+V57Vnz0eWNB7owJ2/q9nTwGFVx7r1eUJkvMsGjVIW2fscsnd+C
4irxJQrAuAAGFwhgqObMyzXiuesPdZFu8rq3PSxldWkPQDvWghVQCIVkUp/i
ch79Gxqojvw1xrSeMUUFsfYQrYx3roG7JW6KUBbUbnfBrCVhxOItWdd3+Lug
E9GaLx7AxXXXd2okP05T6Jw6k2kELKxiHqC0/MeDm9lv6pkAOjpDpuNy93cP
iOI7aXLGPesWiC+8N1/S6JOfm4Fxt5pWtU2a8pgR9eOJpgovKuMEMwUmDIkL
ofOxw7wHXR4f75ViOuSQ58VJzlGkbizVSzAeaNdw6AADohBgu55/lp4Lt7zg
d7lj3T+w48nCI9HIrYq/9Q3D4rIYB7OC7hTIHWe7Zup2ixfjApIfAi6wuf4m
k2s7vq/vkJyl6cD8FNutH1RFOP3SqdxPhM9nrKB/XOn++pw9GGjUbTOg+uj2
peDJIf18vcbFjzsBZSlzofMHyLkNHexN1baxwtAeAs7dY5ebHhx8j71fC69r
KPD5nuH27cBrEkPQdXS6j9C1DaVuXVtNRhyv8xCOYvl6o9p3vlvL/eDM5cxr
9/oIqxoSyKxZPDh4L3gRempTrdsFW/bfHiVHtto8PBKx4W2EerI+zYRxOIcQ
LAKqrWcy3dLwhJY7JXTmufzShS4v9WCFQbG3HYimjm0jkkX5L1pjUyW6J4oy
p2PefBzGJU2lNXt6Qn+uuzVGJ1aAGqfUkEOyoUe/Rr351DHFy81l3xXUMKt4
AVbEwkoijUljkwA7dnPksmDKi2go0kP9DeED4/iVEBxLcO9ku3tph/CXrnlY
mE1jTMwBtxyoD7R92FIm+1mytdNoBC0XxEseV9E9ZdcFAouOQk00i5w2iyvv
il/HG7XhSXrf8fPd2/9um4+dLkpZlxwsNS+Ah6AFPyCpEBlcaHawF5THWF7+
e46/Qle6ko3GVMOQJM8HGKVoiAac+c3TT0ehvc58igilMn8tt/gFaIfY61bn
i5ahX7vGNzeGpH69BTY2rsSNhMPmb02Te+oTpMJQhtOjGRQV3+e0bh9VGQFU
mYQNYmVYWCxtMwDdXoSftyqGFExy81E7k3Lf5H1vravJULCa18nzqiHkfZ2K
yini4DrhAj66zVO4Lvu+5boQAYN8i0iAyKOO5FkBtJmp7z3G5KdGF58FmXlJ
TDGrkeCsAIVpBwtsbq0XPvtaGNUYfF4TOYijOmf7FyzGkF1MtU4qZ4MwgN5c
TaWl5NTa44j9V7CuYyKTYWPbEUYqI82xuAQSa4jfxbmNC6/jNEHy3FG4KyZr
EC6if/8qaAtSHVru9xrVPBxfSV2bvdm0EdJjyhPm0ToTw88g5s2kooppVMvy
dC/mx0euN+QUxcCPWAQjSYPbMyZaTIVShXhW3c4S4Y6ZaHdhz0eqS8oq477T
+T/XcTET9/YzDKf10EeBsAvriNu778kLMwjVMbx1zUu0iY84jnYNoXJHtSe7
EvJSm3e6f7oZtvbISLFYv02HAMtwB9Wb94rjvPz7X2fS0ffLUyRargpY1gKC
93nrOBjnWPS5wf9Hp/Hrk+avkETvnJdXqi7dGGC0PRhBQnrN1K7uUTK9l1F0
klUD2qZsRfc8C++LLVvF1F2JTvRALPu5MQzNA+3vAWcfz+6eyJXS3Ls0BMQS
XWCgZsvpV8TTHRR0jT1IYkqiX7sOuMOXSJ2bcSEuGdfR0OxwVS7FzLuNADR/
0UcRHq2AyCRIs06LjrZV3Y5m3rfX8A7kYCj0MuYou3g3X309RHhtsjATRm+t
PcogdgbbiDwnM+dlY/lvVKpfyVJP8HnTCuQvClY9SCI+nt/YYAaFwj0SXMvz
LsFD+il2A44bG6C33wA4hfEQmKYblr2/30NCtMBvq6+SF4FZFH/MHIHE0L/U
2QEjpGQfyhqZtu4cx3g7w2Yj7BBxdBiw74MLj4IZbynA7xvQTzyeO6LXFaQt
7zGsujMvDc5TWc2d8qZ6RyZoyh2MhmKgUUrJJkVNfYvHPVtgRgIDBZVyfkJV
d8WkFot/Lv4p/anxCcZK5HDeErPqXNAd92qX8YOc6DWj67WMOpyVI25/9KD3
7FCIcTlBbGmLUgyZnTzhjnBDmWkvvf8WnA1Sm/hTzQQ71IyZHahLbJ6iHQ3d
vr8orEfzV4hoZh1Vl0id3UEq84WqF0Gp5X8bF1pHLpVdKTbjR5l9UVleYPYn
o/z9fRCIXgDvA1q6byhQO+LnAUq+XpTJfo6fZcoROcsN/73heo3Ij0sN34gW
vSvgjB1j3MGSS+uHe9Sibe0reaEAaVZ1v5VgxjA5JkgiQRTJjuTAivQfMms2
YepHdNDOmyQeQ8F5o2liN8qaeBbhtAhsTeSH2xLa766N1e1CdXKCd6fGxr3/
1ax5cSMSuq1gttQgdTSZU9Ja5iSnip4z3aEf/yB59feA0EVoxYRTqwYIA/OJ
TRuq4aiPF+PEQ/M+tR9SehiFaZuwt8SU9J09MbStJ5Zxl4NVICAfWiS5g6SI
39TXrOTIJQRwIst6x8S7N1QKxHXtS6aAhAa3Q+NI7/7yWRkLQzA6ZM26AJ4B
kxpEXDhkpdTzB+VVhJAJFpa9+eTsUGd0BJCrE8udJaNVw4vKi7i/MYSFBdoF
hQAgnNLb7KLpWl0jTmy7pwopuxcoFg/q12Ou5bT1R3oa9FGtdJm7kM19bJp8
JwknNQsX8StTcgenKZFdXeDgbdL/yrkQEQvtNbZFE7JKDj69iMtJkNRCb9yR
HqJF18M8iDplsZeA2HfQXlTVzoi6I/wuRPNtjAiV6ymTFZE2sYPkj5BJIXp6
jarejvyaUNpYfYDbihiW5HvoubRbjHYIKxiWw8yLlcCvjW1BwnczwS3yMhPl
j8/aLhtctQFvMyu2pJA6CHdrHXXPQWN/Qr0ueDCtcCuP0bZ4mk5JFdEW5FMu
odGU0xSmam3nyDjh+8Xc0zchDcWpZTeICxOKHz1Mm3js7mHQiGsa4KrhGb2b
oHaz99ihIwZu21yt05YZJnjz8kLHVKt1g/fKPIaQdTi5kRPNnpNWbSXSVy5c
own64YG1nLq1Zdhqm+ZsUtqX6j69GVg8RVK2kk7kqQxfswb6msmOczQgJAp4
qm1pbE7jnzaPuhUbKF1KalFrTAt2D86IdBejbrg9Sl8Jj6IlyRdGcFEeECQp
+b3EOMA4Zv1QgAJ6IFi1eYQSCrhJIJhzi9vEYfjMlnfYrdhoELrGgUH+iQmA
Wg8u5amZE95z3zHCnchOcFAzLgq3A6fqw3iAFL9SWc6IRzhG4Xpzvhbwz916
zB/3MGAI2iQhrwWVCypAUZSg6VVO2af8R9n4TTCm1VcIDnGYNLhOct0H36OX
baALqFBPFKK9hoxdWhHxLZa2GaBuucgyKaZ8VHYxhNKtC7BSyvCSr4eJrjDy
yCHLBXV2Sth0rngEFBN6v1lMRWGveFjEF1kTJncPRK2oUNc4W9sPUNPSyIkC
y0kzBuFDOxwe1ObjuR88aKuGTkPVwPyYxZGH1FmwTrd/9Agw1YJnwxDFY1Wh
PBt+YvIN59mHxvTEdTaAP5gF9jm3t0LVC7cqcREd3K4w9dVfobe9NdACZobq
gpYmGUP35u0qeqIfvE+s6VribUU6CPHknHIrEo1uXhrHLfctVuXCTUxe9wCU
mvF1LWmkPuVQH24lfP9HiHqysqI8B68O0Cxym1+MvsPIqyDmJRCO3Tik2BZC
hV3mrRgvYzW8d8k0nBmxDtjUuLwxBp2ZoYvwb2jIzAW9LgRPb497Z8Uljs+B
qIKUWhmxRYHLH9aEDoogLrYhKgybgQFmnFW/jpC0LTJFORDw09D+yOzsx19C
fI61OGONtrX0SLvwiVmq/5w26JCzJJEP7Jynfi/dYyM/hcFM7Tchbryc5FFe
ueJP2UWxFKz0FcexseKxeNFjcx/tBPdJzwMr7l1xNfmvolyKyU3z8uN0rU7m
1YqLXAAFu9SUzEiz0J++VqlUCio/u91yood1vra0J3V4LjBX5XsfRula9zoS
T0WQEwtE+vJa2ae8fP6N/LnROc5SB377StH/fTMXxEiFR5JwfMxDoHk8p0jr
p8JieM0ixMJjoPZyioyI2pkZsBrDaGQD14nuz55ylHtMzbq/9RT1RPEPg50f
856YO3Hvz2yyQPGAa2714wdjNc2/D08MrD/hXNF5tHr3XQ4TGcUvNqlmYtDl
wc7Lq49g4Lhs1KSGZhIPvBnSY2xRpuSsP3bO/MTW3Dmh8Stls7+v+Y3rvnZA
Ku9dYJ+Y+sU458sWdWAB47Y01qg/zCLuwra66k648VHFXYjRhzUbyKdLQoOD
w7+xVyPaRXJ3hT9F7LKWfZbaSHnO7T7K52h6+LJhQdQnR/gqmARWJMLO4keC
t8tUshjryWnVxeTbmrZ3Z7Qmt01R/Y5u/1eUA4mrP3YZLeBySgVkVxQvYERI
nduvVo20v9U+R/jI/KsJxz5lZDoSNZ82kxR9WtQnQq5ALohoUoG8emUK6rX3
lHlZsecT1xTpXpoKV0WhMDNyMPFgCimUKhy/dYvy7HLKtvBAP2X5HTx9N9ZM
0i6YvxEBhAikExQgPm1f72aXYZB8Fw0t1IeIyKPF+nKtZn5i8fJzwSo/rXMf
CHuFjlI1GCylMgTW5hZGeVrqg4L/zQSOo1dzz9aJSGZR+p+5gxdIzRBb31/K
Mm9qO8YHKLTgqviMgHJc6qKR14Jeg3ItMYX8wPpCSReqHvcuD0HSbkgcrzHZ
sTSHoU6DQtkCiSwvs5HW2blrnZF9CsikhnM5DddjkF/u9zuhxAamQITsnT5y
ibOHdM/GbxrYkvdzy8CluvHtBKMJ/V33DfqQrjWWMTODpi8HDcb8sgcOZiyN
upYsHALGVuPP+hIvv9OL+iLFjxaY4AwH+M+D7YxApOp/VqNjYlzLn8b8tauO
3Uc1VN+NPrFCKP8qRN9TRnDNpoNgzU1m5B28UWge7BtmwcLSAmF7nO0DLTPM
xg05HjLqpnWdifH9ECBr2Fu+Pf7i6Ybs0l23Wo/MN1s3hjDkQYUYmb/0nuko
fKfbjvvLzC4RCWAmau80ikaOFuC6f94VW+avqT4J/yM2hcdlylvN3ZQgp/Qq
R5ADfq8stzlMZVi2iKNMYsIFQOSK8xEWKnZ7HB6YiJaPq1jQJyntWaXjHSjh
9lRbmxMzO947PsGfYoxMtbz7uZh2MxKXhEzJgrMM7QWAJOOYidYINzxs+kmr
hl+wvXsYmlmrHOLml+fpe3ipnwy3xLObtJ+S7W3GmbmU5o93vcy9pBN7TMZ5
UgI+UWGscYeJB/RXyLD73UXlaCyvQgfMygk2mX+dy2qPpQeQBD9HvAc2eEVT
heervxREFhaxSPTMJrW64yIOtYK9nKMKkeuUQvEAqHM/ooEMPO+z/dMIgMbf
TP+pw6XbLgSG0+Bj2uwuza628LQXqjolYCnxTXUk9hckHdrp0rilyPX0XK9M
9yeXWRzGCIfQeyz2qGV1M6CkhqsX0dZoCy5BPM77QXbFkzLdCgdXbRPQZ56Q
qC2Arx+MJveD5YY0FZlIz8TEhf/HeKRwlpbxemt6G1Q6BKUV+8fKNTrWRhuN
sslCmd4p6J1R2+9CeSNWf9TNiySzzFgmd9eUU+puFT2vBzdrYe0oNysUc3El
e47GfA5K/yC+TBttGaz+ltncodOlL3cNXozR0RFikYHaVSZHzfmub3BlRrJR
JGKjVHgYAXwJl/BdWQ8tiFyEIFB8qkVe/hdtOHK5/JidNUWcjxtq1IqaKO6u
GeB5JzbffJ8OThlDUFLfVZeWmxKxo6txkbvEYYXrNYkE8nrlapwNcIs75g5Q
p1qyLN2oqjsCYkwTvO4mkB6mXA91z7G8JSKLTaft6SqFjEcwE6kVq//fbgtE
w2FSZkAhSF1SCumP4Y+fyHFR19C1bW/8cemqzDN9qxnLRM7JvCLmONxGhZN/
yT+oHgJtlWkqb8lljmqex3zZOYVnkPO3xAkPp0H+44B70Chb8xXfDm0dRg8W
3LmLmYkCIkBP9PedoVn9r2n8e+70YZdhB4dTqGxFYMf0bzXGA+HFogYXgH/C
mYMWJ8m9Rr1Y//YiGDLgtdYgaJWRpl5wAbCnCqFBdgjYAboVjjKTpnD2BkPA
VACwmipcISGZBXTsQlZbAgdB7gMSUGiuy699SomdXq2wnkapwUjwiXfHmn9Q
HXOOLpWCBAmLxpjWkPPbigHmrVEZuWfDLvw6Q68ic//aDZb7UmC0M4p4lv5S
pCFBUZU6nkrV2prmKGvRCXGe3E0HsyAuo97qGrcKKmATLVy+i226qkixuuaF
rlHVB/r+qCmLwyNKsc4uLX5nJDRTeGUTVZWvBquHw6MRulXiIuUThHEx0vfZ
ATltXkqpiSIG68mTNrvTjKHQgwP+eltkLigsodULD7rnySrOT9X0NRy83LvX
mXiRwBEv6nX1Pc5Ck4kIadeuIyMtBGPewWYy4n/F+hgOJZgsLaxo1e47Ji5+
LJJmXqlqgXTSd6IfS7addgDrFJdacD3sKedi1gpeL3FX1g5LxPxGR5Zgeina
gOsAu9UsHQhySxkZMsDOKATdilqrisstlrLAHK4byjkMakpRHJxxL88le7wd
gaLWdwY+znlCoyG1CKMy5TqcbG8wKOM6BQAfu29TsAwCz28s1GTDZ9ppBPsM
x4huHFnlIjZk44g+EAgKzOBPbvlCKuufgRwqfjNRxFRh7fH38Eb9Q7z27KxN
r/R1OE/OogzDyH4W5RAdlZtK/FDBS35xtO3nUHOqBiHjOXwI3z35zeKILEqj
eptB8rfSUtY086i5vRuo7u245XgVZx1+btTsdU1EBptY6+yL/oFlSafvywKP
bAYHKiwffBDvYpa/K/lPECVilfCt8mW0munJDDsW/3NVn5qndSURX2DlU8Pj
lz4T/nIT9ZmtqctVbxNcC/9zbdVzE4YRZeqSTsnHGCFD9ZfDhrlehh3hEZ1A
ak57vaaD+eS7TSjQFHtxhV9eRQiKdj7BpnNWNlea121wAJNxM065TTKKaMV9
cztGxirRwCljnAdr9LLKGvFa9RTWrumB2Aqf2YA+rWjQORTBALB/eAC5rCtE
o30J8qdU8BNnICEYmpZass+dk8CSEo3bcgGT5cbJRKQFaD+UJ28qyv2LmZZY
z7eUW3IYndrvuXvd4ShiMwOPCls0iI9GLQ75kGZxYfXa5q1niJ4oWft1NJM6
tqHhgkQ/5T2h9QbYbgcxcFQT5sPz6S8qgNTw/q/4ZGiRXwikvfBJYhraU/nY
aEUB0mn9ySCU6K4UCl1ZlorvU9khlX7arZy0AB0I6MlNH1Y2bAYCxevPgQbe
MIncIOOjMWeD+t7bGSWXiw8uyHVkk5RY5bm0ZCb9VHVyuGnlfzBCTGyYIBwW
w+tGOMrfvTMorYRCmM5zmhAngFx7tQHbqTw8SRzJUKyJQuAhCw3+aF55Vz3A
fv6zHdTHtETseQWpprb5hBNi/0C5iLUteDFZD/HjfmzC1EAtUYKtj/DHeArA
eSwes0kKstjdMf6zrj2sRdOxPEfjZ0e5c/VgH68UBvou6bkCybCllrBbQhBx
7l628IBr2J3WYFgl54tW9Sxe0KCLTqKTaSUBfhTuVHi6pvMg+nZPtQx6AJcS
FFXhNnLcPnSgnILWc69H9oDbTQVkqG+7weBmqWOAzsiUnJ7jCU7udax9J4QI
Tn9edd8lfnVR2Mv4zUIFLC0Pe+8ibzpQsCxzWuenN1UMQ0jzMuRdHAM0IlV0
Y05TlJvyAnZm2A1uWR4U1393ZrVlzASAX14EzOmv+Yak7HS9UleGTxlahtKw
omRjHrHJMkISEKMsdLDr6WTmYVxAhuopqRj6HqKiA79g4zqwFxUSFK39Gaz0
8JU3BgQIjBmbVo7fhCZFEo5VJgtUewwYrl9mr7wbACHi8t8Wlub1EWvSr1DO
iAfDOh3xWYrgmfa2drbBw5ps+ufY9ziwY9uctUaTFB+ycbX3omXxErywhlAO
pAsQ6WtDymPHeevqKzZf3LZuZi6svGN2SOOsbQX042WDxSjoBN1b5ClBGyw3
38syh5jB3KqzhKYnNt3wltfLHCt0l0uCtwsxITVC3A5S6pnFxTFz2Pn/7MQP
wmjkjLLyT5WGI2ln7+RIsBC/Wh3+R+3Txi3YlkmEAmoU4AccJpEyPDL8NgjT
KIIN3zBuZDrc70VtnInPPRXaQrWmOfDWhjl6vMzJoPWez12/wcg8094sRet3
J8OgDYhT0H2+IB2pqhFM8d39pYHOLIdxqyu0DjCIIFJCnNRyKnRUZiOwYTRd
bplxGk+kYfLaL5+8MAgTZDHy0SGg9yWP3m+4QuLi/iyovEhhb/brktUK4J2e
VXIEYAjdIVxsbdX9GDyclNLokBPO85zZQ7OtBsPREtidgvNgYYRsh02JTL1u
kg86nkQesjBfBaPM6lJ3YU554ReVUbEp1kS42muRpXJiQLjttpQa4/GWJPjz
8CRreT4cc2wc9JFyCj5/QtUVHmOMhkkCbSDOMU8YYF0gIKZ7yJ8TG4u5OJqf
/0nLsOCPlzo1qHcWwlaJQFJF8HbF8uj90XqD7z/oSNTogSCSAlJlcm/m4n9m
UH6cHlXL20Ip5pH3qFXMVTLPwDws2nmbC64OxcoV5jCRgW3A3nLGg5e3NODh
jVPcp6d5yr/kV8drM4p9VunRB7OfSnO+vQB9GIrNXBAMLt6p9ncoo9FJmaJK
mRT0S2movwcoXRwPftQ53MxrjaJfKSXid7k7stSEap4VvVa8DSPJkSox73K0
LrTk2tTlbSz0k+vb32dGmEPPr6kSoFki3NNKrTkCo1SOQ+Aa/AHrc23bPorD
r7YwQaHrcWTf24ZmL3JRc8yKjW2Okm74zRExczpdW/C3M0eSEEdXV8CixcRZ
B19+Y5d8QqcffoAm5FJVNr7XhNCBUeWAz8SPcOKI4GGBXzqE/Tk+rDNq+3V2
+vhn4JeA2CixpdbBJuTmPrOheGyWWVRZFprlIWfipD7X1F+6iZs+QYi1xr65
AW0wQCGrSjYT6c50R6o7o6mdyVE3dfUGU1/4D2nCBu7GbhylnoKH551NfBzw
3T5wNCET9sSCgeL5yUYvSofsf0ryk1jddv2oW2GeAF8i0XSS2+JhZxhgq3aC
gUYvj3tUZSfXTZtNIph0mj6f9R+bW0J0L7m8RtvanHenTN/953O658nnOSLl
Jca7fBLipQvXvipdGVbCMvOC8AseydaZ+q/+EQk/yobMktUbIMFlKahzin7N
uLgHym7CiPY7QtQj20K3Rso5E6eQg7Dr3MwFbAzSJKFCn69Hgf9v1P7yGPdp
WqJl9LZ9eFUoaZ9qe+vBvHeB2CSpeOc2fx3Va0nD+p89JwR9s+fYwhD2uJ7N
E4rEQQbXrzWUl2eQ/dqOJr/x91f0S9Iumrda65FC2CDtV1cR3mnsXwxCszi3
Z7nREjfupf11j5xp/6BA6c3nWFBihdBJLGhn0LYkNGotRlGeq0U48uWYs5t6
lC1FdKm1ij4/ioVoTntX4j4t2/MzSKG8R/bg7o2mkAbEWMrY8Bx89k0u4ICt
k5TyDEUx8BtEIhrKVnKyI5qMoXtEPv62uBRROmGb5eLGl//Vz97HuOm35rXI
yydTFKGyUvc6Hh8yEdQlYPy04R2eDlCJkBFZB1manml1l0aEqkiNAsieiqec
dp+SNraCPJ6H+fMggwXu57w4fkKd9yT/AvayROAd4QZXNRIZ/rtoHVLS6nS6
jsOMAhO0uPRkxzW69wabJnA50ltucJ3CFHKganYddKVxu4HCY+7JZKVwIAde
Gf4oDHDPTy4qKtH4vWQMKbJ0hrmczStXtiJLbojj4phZ3L8ECtrxgUwRmeZK
gJGtNghLBl8rOnw/jZTTIOzGaGCKCxJVOx9d9fKJD2vsNXZiK6YK2JmVW/Z8
7nIwY3S9ydVYeFhMYNUfE/EWGWCcIN1G3WgdSMQ/2lDn3OjjAHMr1GB0TzM8
eNVU7yZZBW6vga3JUhMkSK0TRNVr34wkGSBpKntL1cq37shPPe3dWsYnoDjk
q8kbJBfsqcJ5WXohi2nkpNUMtw4zK7Hro/qOHHSDQzb6uByqko8uu6PfH3AQ
SghXCuzVvJV+0PKdvBRDOrDYKAB+aoaE0VUR0ouUC6nGq3SyE0DH0lhAI49B
wM+/jm5eqvBPh593AefIWJnSjeV5uxuA+vxWUVRq05iMkae+YnyVJwJxwH4i
eDW/fQuYood+yeDm9FNgyyQFT6Jh9hITh5KWt7eVQEXFrS87Mf7YKEiQsdSo
9HwqYjeFyzlDJRIAgkh5wD9v9S1BIMtZ1fGWxUmf132ZPBRK9U6kRgwWe05L
zVAd/9Xk9nlf/LERN2WKQkq52djd1Up7mPaNU5dIeEauJeFQMrM2ZzA3T/jj
XHMMueJEs9zkJyMGpLteEOp2Spu1fy7wr4aHi0QRE4gX9UrTH4CSJgrKsmJN
nN31riFor0ek/Q+ZLlk/sXS9DhUiZs0SDCstKV/kV2yO165ap6O4whWZ2Fxf
pli6skZnaKQUjPyeWyoLzkDymSIGCMvqSuJDFMS4Is1XTYdv1ktioMjVhEkf
Lri0oSj4IGlzLID2GeB4d6wzJgY9S5cADgETNcvhDYQZvpXagG4kYRbImbGw
YY/X2tMCtxLlnI/qjd15axKONGqmqtpb01XKsjXSeMxKWby64HLNaWkmcHPO
lXvejOWH1o2Jh7lQnMksHhJX2l4w5ic1XXyUR5j7+RunN06ZjolbOkjekyXQ
rYeqRcXy0Ie3sDYjXl7+rxW6Gcax1+Ld4UVPnY4mwvPcCMNEj084Z88SvEcm
00gW2CdBHnb0EgIzyNzicDsCGjDzESpXiFAuLaSeLelkKAGVE/xgSZmviKKz
/ClAg/GiiYZi+PGGcyJeBpn3k0f6Azq2jqfZQNYt0A7xFY8sayFWJnPEAQcU
aCFEXi//DdD/Ga1qRqREDs5PbxrDFlXMCSmr0aROWrpKgs4yeKxq3lZ0UF3M
FlAl9JAeVNiABMds14qUxWJV+rSsWCkxAWkdhJzvVcE8dC54ZG2erE4cJ3Jw
ABlAczxCAZGOQ5V+DevaPbdYrM6ho2CFIbSQhjX9oC+jMavGjEWsqfHFbyIl
W1WeXY2Yiu2DTkJs2cCcIGndoIXHFcdVRyeaRs8cxdxmhhzR/rmS12vV+t7c
zAFUdAQ4IlidkfakCoN9/IS/vwZ2TEdWR3jxfIsKMNb4Or2NPIcRamDLhG3/
nuAclDUYwmZyipbXy4qumdcbwvLhyJ5H9nQlHdNn7Y42WUjKOxMIHlLms2zL
l+/5dtEtg9RLqAeA7RIOw2ux3TUOaVyJAyQs8+NSkv7dbODqoROM2znmQWn0
SYyB1phpguLbGlSSfnwGpv+zGz6X4VCncmOH9ZaiNfBG89+ZqnzBjDXztU5T
JLebGc9mLzkDdaHs+72RwFkWPqSKTAYL88/R9b3lnmZqxdAL5Q8cEzS8qpX/
f+7pYqd0+PnxGAhPaLeFgG39dn0X+LN4vsP4vVqhaMkU1ErPhefBAtiHLuKG
QScHXbYcYCmdLjrHToyzYFuOX/iFlo5OCBgDWfw8p9rMG0RJU3t50Jt9WSla
Zo9bCvaPYApKI8Cyey5kiJ0tOj1BXYtCxfapw1VqHNL4FMvYI6nuDal20pz1
3qgsCq2JgqvzAlMUJazIZEAVC60EZBMhzvL3iLYYUhmj2Jm3EamYcedCZXUR
i7fl23z5uxQ8oleTTeh7LP8SVGx5tLHsFpaK03yRIyETaUVpGZ6qso7tFUj/
Us9yIC1dPEfajEtqcy4IZhMh7S2fTO8UXgn6kIz+587uRnZM9FcWc1f5Bsz8
jBo+CG27paxp2OMOgY/npATrRY3/DCCokaCF1b5mO54ohC6gbkdksSMjAdfX
lj5pW1GL3p10b9bIRHGv33L2QG/5MUkMSblpwvW1ns3MdLcj74mr/JevtOH3
DVHnX+0tTVFunapN7f+6I4k0XSwYRbUyjpWAYFHXXQAS211FjinxzFWzr+tT
tgKk9rM39cJ+aundeMYsj1fW/3HoIHrFL26yhQtiEwwkklzSt3ayYNt3RfgX
Rc6TTH5274F9VWJY6I239I4WDILajEj8W5jrO9QsviuLIEKtdgn7UxMJPo5i
3JwjKCfHWf4oUz7bAcvWdaoDa0xSDp0pGhxj3YJmEZyDLayoz0b1BgmXR9RW
8uaD4FYdiBZbMKu8pb/riDfT/5p0k4GDO8FQYCfXETv36XISSuGfB20RGFkP
FBPF/Esv7YOrsAbpHuHgmWsy7OaG2vbcQjTL9C0iyQwp85iOjEcKf+QSf9Mw
BKVXByZ/iHkTPXx+EM1rU3qaEzjtgaqNWEarnj5pKjSEuLSxULl1O7ny/wuZ
3xW52kVJlMlFEtsZzTafDCyhw7Q3XpWDNSlsYw5gjL3MSrruSmOuhgVj1DL5
D9Z/staB9SpBpgF71nHagrG0aDpzQy+8Y20G07HrdAT0jLEBfGP/ifwy3TcL
rLk1A2RbG5vuid2la3CAHxvm+Vrwghm5jR9SKQ62Om+U19ND984SLZQJUUas
AbsbIwa7WKGrvaxmOFj5iYscj8vZMlFEtZddxw+tmh68LpRB0cUo4TEjKsp8
+rwdFpGkbRxM+2TO6KZTtIfhX0ZCxdKkHWZSzvfQodW7Nu1+C+M4+rzGU7ie
NKE9T/t75hfkdOPeVsg/3VqSaoRcCwFgdfoyausTAlvPC015Gx0bDCLdx123
vDMUg7C7rs7CFi/oicatlTy6cy67YscZvJR0lF6jk3vZV/jcDhf7nA5FaAtS
WpduDkiF3oQEBO009NJhMWXbdA3PJuJFU42QY5p2NoAg/X9qfsO1hYSZDXVx
GtOaoGvqWXZMmGY6HLwTyW9tye/ntGy02hcOPSh3xyFvZYsArgfk3fIEUB+h
5gRTcDLchGyQX13gs/lKhnOWx8CZJBAc23ZLaFZ7AwZVZbLzZp3TTg3W0AcN
hLmpX16jZMcg0akuh+YIsZafUT7q/8ue0kff+K6/ON8ywJTwYWuhI03pTZPp
ruFl33E0IcvvGvfwswIY7ELcnZ1vLvs2Wh2WlgBAcxbYTC9sebPgrS5XNWPM
KumltQyHTs1Wl+qwm/e/1zzXwoE27ih0lnBESfMQOKdMEoGHsFBoBb1nmw33
0hEp3FBGyyn0N2IFehw/kyJtGhjzTLZO8FUXqz+L1l1sZRi4nIvLDkxG2/xU
0rjYXT5SBp7kfWoC9iGyTlX6P8nwlN46DIC5re6SXuhMEwoh8lQgu/7brNI0
z0YD8+0Xgzc1rNMLuy+t0gWLUmXsEPTRhnjeG000Wpp6Q8QS+ekFb1/oYk/P
J9aPA0n7sZrwv7Ubajk9DffptXBWFj3fJVc9hn7FQS9dj2ix+NOLqLnBiPA+
ezWW0QtehRn7+QmlZP4eGzeEc9n2gYwikKjoqFycWhlg8alrFnbTPsArX0LO
nXxJJP4e/SsUgtDam03dkjox+BqSYZymQXsrLJBvS4h7PRcjFIvPY19Ufec3
1dJzhgD3zxyTb8a0nRrrB3M6NcyIcEBLIic62nVkfHsIHEl52S+GrOLjxpoa
8Tm2Fu8JHD+OcFC2cbPMsXgEoe4eLe7aVkqzXh4Xn5O2lUC8gQ2SfQPLZiuS
kzU+0FK9xlYlqqSyCSw9ZB2Ftm8jURRKF352JZDSNaKJ2b13AUi+YzRn7XhF
dMXR9cPEltPPfdduJ9Tp0sUKOV+wgbwA1wMPJoctg0mOxPjwKfprmJsjAGzU
ouGm///7Wic1BIC9lEUz1X+xwI6DBfTy+FdshgvXs7/iYHDRWaTQo/G6G3QX
8AaWL+GnKgHL74lNcEKEx1NAvqWShru1/ddfR/Kgq/r2z89dSAoYrxkzaZfg
lzJ3tEBPguPx2BUULhvPvmsqnT8NaHGlS9SCmJWkReWZZ70InPzCo+zkYdVh
go/jJt5ynAJIA2nPZjoaktCM8uoKTvIR/FbXQLJvJw12v+HFLP/CJ0XH/mKr
imP3meGk3ylDkGrDxtHadPWpQdPEIb5+kwo0xuxblWfXsWqtjdol24e7pY62
EPk6J6GkJLUSz+Wz3PcbdZKBecDy6f8+xVyUQzaTwqMpBg7Xpz5yxDMpNxkf
S7fhZYvp0MPdyNZ8msZK9Eiq++xTRspV2z12tUkBJtL0l5Kp9NfL0nU9Li3f
qIkrFDs2492z0fZgzv/j7Lq8AMCro4nHhB4S9tEAaGvqDQg1x/X+UjSy1GG/
Q05WapqH+6pZxDEtnAIVW1KYsQhU2tjn14B26BSx4Peheg8OXcXqC5VzuM7+
rp6r+uyV+qupaB4c0YEY3rDvidYZa54SspAkt9qpwZ5j2ygdFCaRjgri8qB+
MWaM7ZG487YVz/7xnLKAxd2nx3/lDqqAWc5Q7pQh+H2GEwAuC23Vx/8EDZlx
zYgfzBKMfS17j6U3i+DUWmxvrmuHpcIEwzPa2fPfpR+DWH7IRK7Cdxk3lB8M
wTkBUiNPAkqzaVvBvxhPTSL9attBSoLBTq/8L8M+gOdLfhGXN060PpmaF1RQ
w33wRRimBrV3O+L+2Wo0CCyWOaSq1pRN+UQck5BIxBFZPJ2afyEnjVHFzYZ6
T/4o4swFCaTOmKDzq+RoWd9IButxt1OID7Us6KW40aO8+ciRxAnQKOaPNuGS
pNVwR9pmhAs/+CiRhGNO5ogOQv+HWCr9GuNRNMTbn2tbbi+fjXCkM3hYSjPX
ViuI2HxGNVnFsJDW6kFSIVceCNUhTSG9hJDEglA1Aar9phBOWCPLFRuXhrmh
sEbFkyl2ukolKqarKOiMzJPy58y/Jxw9hszuRGUV+iWwD8+M4OTjZ8vPOMzI
syVmUPSeldmPks9O244/2s1niVWN+1lOIeJIMkCHjDMCbagLaHpoY7Zh0qlt
5ft7uH5owT1uSLdwP23hoVHXeMhPLrUzl6EpBwKUsqsGqo85pbMLzUC1EBUR
oUeHXQgVwScQbrqUtwNCEVEAFc5Ws23MsGzWqFOtxt5qNfsCAHKaq6FFTvwC
vLaCwAowbSIpn2I+pI8cZkNMF6mutqs+gb0PXM4rbg2vgTT8OCTz7ydHxstM
Zd6JRjCo/NaCzzzLmjnbzV7LqRWox5646XoMQByqHdY2rg29ZWdp4QUAinb2
yFBdrZMVF8DnngLWXFfuWoJ0Ya+wDsAdJVhEDb1pMYA11Pp0hGbdnxpo9dNq
j1AZPEQ0QCkh67cWbH0ZrvhgJKupECR4ghYwu0sInkTA25lQbsfP7YIvlCDj
N+JVdvXrCm9nGdRZdi1nFRtGOrbXzNvjkOARrS7VKC+oYto6kk54LUJg+bMB
8jFsECU/riPlvSSMhvlxHuHxMn77U5YkoCHEsXM82wXlcljeTTLEJ0lImFWG
Qmhwc9jZbG9PBab80cGwYvNNCzCz0h97lqjrJVWhsCRCitH22AtTR9bGWgbe
hPlQ8JWff++fkrTS4x9ywZNb35wGdtWfRwfzpWyjTFSgkXIX6G6TvxWefiXF
25f1SArkH3TRyYvCIsqSdGM+v6qrhm5YpAX1Yo08Ys1Yda25Ko20tEKEDY55
1PbTuJawYp89OgPwrjbB8Y9365fv3ycB7v4NtXyzOPWp0GzzmATle66DPrWy
rExjBwPxuDgBddVJBt62IJ8mUyE/WoqB6WbafGi6b7ugdV4VhTEh9sEusk5l
nxOn0m8UIEpjgdUKBU7VWG14nJ+7183LPGo7PKmCTUepPuXoejlWrnTM3ugv
baX7qSbBjSTZfTXW9NLS1NBIT2dUV2gpw6Vq3XNz2hUrVhNzatIWB+9KxNSH
C/yiweTZVAmYnUMhnOP3HHm7eJG0jviVCdHvNEuSwSupoCKcRoGB69neS/eR
e0mqVQI1GRD3dj14DPFhdljlarKr1bsjdI9VS4/Ntdo8VBgvUlRN3oyIxPJE
bEc3zh5dr/s/jT18eRPNJ7rjxO7NIKg/zzGl+2QHhxW/ZGveSE6ihW+RrpiB
32F/2KWXqy0KuHv2g2SfqBDcaExDPHxDIPRgIwOkiw6BvoJq9WWV4f2dFUPf
77QNeJzjz3Ft4+Nl6V6A7tILiruflYoXeqi8kAIHCOt9QpokCa4irqkU4Qc4
fjCU3DLXrqCvJaQbPNw2LjDjMoMuEdFAqL5C5B94SNd7AHrAMtGs7ShBth1K
te5gDYHCvnkcyyav7Xz1sMPaoGoa8lSkzve6UXGW0C/JAjx7JlvXzd/T5kEx
zJ8RjxA7Mkr/ZZu3+2QYTIgO+4/+0uef4hvaK8J8c8pPRaURD+rNw3UxfNP9
NW2Q78DmQS/4qB3kzlT9a8ecdBYhWDQVfqBNqEh8wRbVXKd9J0E760bSRwNZ
j93DJocT4SUdpXwoEh9fZoRG6tgQ27ofkMN43zAn+TIPmtcDRqCOBSDL9MSP
UCymQmhlnOCNkA6wzYwocgQ7ZWhy7iuEjAvojHuRL2DhPg2K8BedikkAzaQ+
g25ccS2cyBR/eQ7sOtp9NsDZSwiGpeAztyCfAlVUY0JLgwpMCOUxN755IA3Q
DM6JaG0gL2PC8Qqy6Y36fNjzPxMl8A3ZwetAVEg8ok9W7K76g4UBD3XRWR7f
kH95gBlUCwBGkoQJtiPOQKD5W0u7AogSpy8Iq5K3+FFJxZNmAHUgWACTt9Tz
wjhCWs3f15q4HullIU/C1D1/suWUG1TnKgIzTlnGKQMmP+lGAyseCa2cgZh1
+EC0KTdO1fy36biTGVAQJBNmKyd7K/2o1mvD/Pg4si03KY4z8B6Zw3saEhHx
wi8Bt2TRdbfRFMHye/3LSgZsptGROc3aY1CefcGgBrz2BzR1MgwGeZy1OOG/
ENzl3P3Hn5K/e0usjVvhuKlEvJlnoovP4Px/n04mlWSVBu/OZivcXCsqPko1
crA1IPpx8DO/6dHMd/GXQ8NFyWsieuebxWsYPDZ8DmI7gRgsCb2vYwDRSBQy
ePkxB3wwd59YEHi2xdGVzfo+iRi1pt//gngx8hHnytHd7R1f9S83cHPq+2Ey
haEGSqCTpH+eqt1tDWnjwmTyrE414i1wbAyGVckZHHAdjXXMht264brR0m2X
K2VdLHCTJrZJ9oKgfV9X5Y/NZupzzEiDb21sVzXkPQQ9Vn9pfEYFLMoVBCWn
F/uFbRwPLzKUOyhEo0V8li2mUNnLXii+uX0zgilc0XFriTkROXpE1jWHm0//
XZ9Flz4PVnLSwDJSGhmLyHPTPJi8r+QElTHmQRUXj1tuD/TU9t9ew4akrWEu
foOO1likA31RPZitIotpmkUUM1OGHWpgZ36TpxvOx6aImxpGedN3gUA5K7lg
66RmNNzypmwpNTe3GIL7A9tcZ3ZS6oAX6y1BJQWmABeWqdLrTvA7be4FD6KG
rcNwFELrGK4QbfVuvPs7FwM2bkvSFc6Rw5vdWml6iLgVHddE1iW0aNxoXamX
4AvbHqCgiPVzkwZWUAGaZcEyazfH/iu7449oQStFSxvpbRDHif1sgSNTk7fe
KoFRAsTt4VSVMBx5ZNcTi1syjl+PK7lD0Y7/T8vkdQPTIgq5KgyTCkEBUn02
s8gsvzDz6Hj+nDsaVSChgXKrb1N+BMDaVzPvmmcnXzjWHyXqsgDw6RnGjQyQ
y4ZJ2WcbxcbH2apSsy6CZK+QqGJ7lURPGuIHZwhaSgC1pTpQgZLMxE9Gfq9k
r0fFml6BG0YPXDSKZtu4vzmnxESeA1F1598GVdTqW6/F4XyyOrHrexzIRaBB
p7RShcgzpd5oOpZLOMM7OSmvUw8rKCdIhtnyfP056lYXQ8dxFQZQvn9T4w2y
fiyEQYJrFz6P7+NICrnKK2cNmO2qLQtZG63o9usn6Oek5Fh79Mt5qCjoBDl9
hPPOAAd3f0sgic+Rz6giqk1RrTASJHoA7W5ExCUyabTdC85W/kPbcfHy+PxO
Dl6JqJqwAOAmPJsQ147fksLYwG7J5HnuJJ0VIuJ1/fI57G8IcbdFmA4x6Vvr
46BKbI6EPgBV0w7VJvcNwTG2FkRZhPgoG+6jy/cYzcJ/dTovDa81ETRbfyGh
rxv0gUuYXRIt5pMyiEmnCUCurjahbLuQP/dmp+QfEWKVu3y/6OQFeJHIPPiV
FBb2j4e/C/vePuQk0gjsbzVAZBhGDuEWljSB9Bh8Nr1CG8XyiwbXIlR3YPAy
2kCctuvH7xOgUSWpNDQHL0e1Uq7B1Mq8ckp6mtAHL9j0CUcIUittaAcwyup0
lSFTRPGAPzgUlFCQy/h8O8liKshkWb91dtar4RJhpmo6EKa/X1hrzstx3Ui/
asEXm17GqwzDXy0ftxqT8+9Ee7CIxL4ZRgYTxYAM0LubJnMZzdMxwrKJHMJQ
5q0z73gLqQaZBlg9k9ePWS+/BkmiaFmDCh/OWDdeQTWOaMd6ybQLV9qy4yaa
9NMJHRpvfWiGhYUVx4/0acPre2Gyfvmec9D8EybYXAaxMFNBWJrJ3+QmDyA8
qNhHY/xFwASmuv8X5ntzEopEFykK4NyQBqucIx/l8+A/GcOFtTrknhjs9gie
n4XO44kEZerCZsajgIUBUFTyjylyciVq0MwYBi6CA6nCg2tAcFI9Q8zWQ/H5
SKYrsspGbiZSAjLIbuB6Rf8avOV0YicgAyzO8btHmn1DUzekLxYG64eGICFU
W/Nw1Ssq8pu9jNm6cM3JCiEZnVgl6QVGn0gRDFJUPbXUUduQptFiMCNW/2gd
xYJpk6syix6MbVzLHDa86xCQc+aPHXlGKS1nUmclVPhvo+rPmOkfonOB7QnN
WWkUI/vW8ivMNGdCXptI6aLgSeyZg3u3pV5z5c2zMwNxf24fjesdg/6TO/fb
NlpbJS2rm3K+VusMa9lnNH9/L6y6Br5RUnbuBTMjpHF+xGsLdhNJTtnYyhql
/uZs5fmpDYaS6ZagjDgF0ApCJaX+HoEjEZRqYtyB567x4kYn+9hhg+Roggpt
ZgCBgA4xyaKAe4JMLsAl8Q7L9YM84/Hf6SZ50p1C7h7a6IGmHzAHhlBLZ9wg
WbBPuhgATuw2INsFptmiRPPBecz+hDd8Mg5N6AJLBp28EO/IcoUyrk9XOgWX
E3YtHpj75nCpXOlZKMAqtNuZo7NHhNjHRDo3hwP8N8gYdxURt897BU4afRkV
WIyxHW/+K9PB7l/T5Z/ScFvxL0pCdM+lCzyUwijmErS59kbcodirvbxvWKeL
9cjaDo1w/2EayGguGvjuHQh+QX12nLSoJwz1mLscaXQheHesLtzAG7tdNcOf
t9onNR2uYj5o5hP/BOFRZGqGxoZ5uNhuLFTStf0XjcsTZUQitOgULZ6B04dx
oZ/apPlciIkUqT5XIUQHgNMjfPi/MYR6+UIJUZqWxIRT60qvF5fBrtEX1rqO
TPPpqo4imgazJyp91Ri+BteFxc+AL0en9yNQETTDBPWS+BXNasBSNzeEh2BC
W7yon3Aj6DWK0zcKBxQNcm9UROwopMTf62VkflCQ/YDn5CitOuFnD343q6Ag
OuiLxZxpvfXRs4AKc8sKI1AJqAkc2bMLPQ2KzodRb4IAwxFMx6w//vvDngUv
yp1eaZRaOukl4ku89yBBOZ4skMiu5bm2wnk7R+SP6dTsY5RnDyEzUI62EkHJ
YO2V37Hfo3wAU4NYlK3Ssj4vdOFlBVZV/ymL7sQR+khYfZDFIgw7cXlSA4I6
NuW3KfJCZxi3RWJwVI4bO2BMvIi6eOzt9RMdBngrZhvt9c+aNSGIt+spmkpB
Nu4kLukGIRkwsesOXaM1BsY4bumC5civhIRcXh8Sn2MchJqYn602CuJshy7B
kj/epvR1A/jNet+PXm3+7kamEt/myzbgDYyVZF6N96n1UCKj9zLXnAKSFSL3
I/KzLRgSzYXWl/M304ev15U2KcMyJQ/igXhzc/0BE+xGhj1a62QjI7e0Xh61
LSyQm1LXuDMJbeoL92A9zUGybkp35ZQFzgkCM9tjuQYx9fFoBSgwDrtBxTAQ
GH+Sks1f5DZpmGZoiNZYMQA1CNDMIuWVKvSTjEomq0V4CqlBk3od8WWt07Gl
OQYENZmZdyliMgGjW3wxuGWN7cR+P0LojuZGkCpGBUEpuKubD83RUpGgZw+d
wFFIHhrIVs2GZW8y+DXtMhL9/oeUHpDvyCWx6OsulrubEZ3jhebbD6C7qx+N
W+oep00Z3+w4DgJZ/2mU8mIo/g1U/dRcYFO3JJoQCWDki6/LhwoDgzDKb1HH
A1K+BfLLcJc03u/4jECGR7isVl1WHLRLVtshvMkYVvTL++Kv3xWSE6hLEBml
9cxocCJSQE3XcAJ9YhhwHAKUD0mpL4fAhVUHYrw3Ctjx03Wg/ISuRlisnDPQ
zRL+iiqNANOqKQ3Bubuf2QUIJ4ek1InueYKZrOv1IvvwDxpmr6jbOH5mfMXN
y8PrsvUnOJhFzFHWVlmByXnymKI1GJnE5PBTCNjboeHblQrGWjDm09C4bMaT
ZzciEO9zb0Ui/9p2jBEyJjuVcHoh4zw1T+JhXhiM0nJ0mn+Gk/vUpmFc3kKC
KTmXN1muB7KlB5CslYLOLhIaBiWLEB9c2fPFqrBsxFNNqF0xpE3kzEFda9u/
uMfz/5xdPIcnVyvm0NY7ei8ap5Anx1nk52wqazpYUS0D+Eldf39Vy4TwYuXs
0iy34WLf3X5KAq+5Ch4Om+jbDpvnBbapObrez9RbKj6YZYsJ/a3fwWj43Mnw
Ff5M/YCrJp4bJw/x5n9mQb2c3+meuIMqymIFGkGgD5M4bRYUyPtfpGdHQV2W
rJA4y45Y0lmc1v6ZelA7ZLzlVbMRg8G6voB3fdTzSM94KTYxyw+OW9oqT2sg
MOBXYh9MEFN/8pY3WSM5NoZO7xcaKR3B6AxRgPoTP6c8Y0zK+9u9k6PAb37x
/PPpoTb5V4QTpTy9jvce8c04Q5/M4Xn6Bm6XtZDGo4tn5EZgL9J5gBPyaqMq
9qhPCUeIFA+wjiaa+Ps/maoQieqT5FRi+etsTt6eo7YFFviu+tMX8n0TNSbE
+jLw0NO/c49sniU3GkKY86AxdPQ9/BHfUShBvQjhL2QFzX9IXSK9uNnL/f8E
5WVMZnzhqGOSw/va3JtSszSiyMQtsHrW9Nftnz4FqkBnOdj93LigFZscbyg4
X7buecr7k5SPpElCA/asbXEAFVoX3TsKcKg+z6PwKgg0DFzsC9wwIsitMqQT
UBrOJ8gAX4NMJhQnvTTLuUNRPmXh935RhFlRYxCieEVJE/6PXSRZytgax09g
UrH8RqICPE+SM4Ky6f3PGtCEE6diI817/A6DzP0uamf0dyorHQb0l3DtFfCO
AIG8E1JT9rjF28QWjuEoRnXbJQW7lc1ADwLpA3X14vmWeUOPHLNHSRzKdYaa
pg8OzQFDIR+Ubppm2HXAyVOg9b/vwV93WK1iCXdNx7zIvUC4adhjGaAipBbN
YCppR35+pY4H2MBlzUD+9toTd6e0G/Rd1eH/qK+8InQYINmgYJSxAYdZ0eCG
vkcUdrcnuGCflH7qGNvSgkyJf8EaR8uEjxVziO/IwWP3WcnaAD+QAPZ0jHkP
bb1GP8Sxq+49rq8EdINtFlcYIfLdPPklxQe2OsJgQO9Lu7s1mM3/Kr0rA+FY
6xbcG9s1vs/TS4AANGKRPVyFF9r2UcDlV7HwoAlg55W81kdNjhGeQlBRz+up
A+SY6Lgo62d6BxB9RQOrFHlVgaqWoz1JP3cfBwXZTKL6vpmEDDGsT7VSgt15
35CAY/0l5WrtuIEoj+T1GIf1x72IHQfxw7GIH/gHYOBbq5HiZAw7Z9dJe6py
Co3A+NGHst4EEF11XxrAUBdg+rr+Ab7fLgFlIbmlcuhbyelbWgesv47ihEV6
LGf6SZ4GG/l6ycJf3Mo9o+V5ABy2uiNhB0KW+cl7w9FWs3HQVMmoSvY/6ymA
a6vSIi0KryuwiZmKEZtuMfe246ylTc2ePl3bLfJ+4VvtytjTFyH2ysJxXBO5
ywxXZioPVlj2J4s6m8ve9jOtd3iIdrAl0PHoXw0eml4ZQXhhA7wlrba+E+5K
zGTT+7BxKUgqzucebQWcDLCSL7/GdxzlKY2xWpAAAoP/H/8781jdGpMfSeuh
jPqZc5O01qnMvGuxaCCDsgDb8N9mugSTPWRKM3IjkJLRGsEvboPPTOQtvFdg
nHVVfn8A15oBevU89FMxPJaTC25eCU3IYW8xfQ7f/4K/e3mZs1XBBj9tZvTs
n8dRY7aGTgl4/TNFPoflXkKW+mRj89bru4X6Ebz4hj7racG5oyodwhu7RpxC
Bmq12VTYAhQS7Fa/SVu1Lda3yaJb4uLCm3GaIF6rOtuqXH1Olqjp3O1G/n60
r1o7DgjLPjUNGfpBPKExQGmEV1k1Su+5o3xeSMvOZmdiktZkfTRrfxr3FMJA
3dQQLUMcSvmohgsGjizlteP0fwT2sQ+PatIpBLV8vpYCFINLOSVu8jTTjdp/
0wA2ES3uNZOH33CbXMlElw2zidxklu1jTzrtV9D5lwWkyDn6s62GtI7U17PH
Ymfo06JHVKvJRAZsfDKN5sVgTkLPqhaRamxhsStHkFCI20CgA7W1KbyMyz6m
fhF9SeY7AhmqpbRHmYfiPBPgbxOpmgFCQ8SGdvDdOqI9UdDtmr90QOE2pcJ3
C2xgjpsvXGPa9F+lugMgJ86TOk2NQWzM5wKwV6WUbqRnhcqP8qlLRj8KwJAq
AVUYQxvYrrM7DJk7cKynNNvJKvJ8bski/bCd6qmlcSc/ivh3WmqvKvpsMtmL
L6A1U+M5bOlVohjlF05UAdCLHGVTD/uvJh+LSUKZFpR8avN+CHBeBBrMd4eN
ulkzn0XDwsAQB5MdgGkpfUtDU3Iuv62Ts8V8QYviIN89ivmVA5i6HmPqOaWX
w59t3qdAaYK6qXj6xIaAJRxdRpK5PSGHd6mJMCXrs8G9nfVbcYLFIv4nRMVv
H/4+H6FVeOPHy6iVJUHt0iGIFosr+kpk1ogCf2/POVN84Uko0gSTm8kKhbVP
FBkJDanvXuRf/+CL8QLr9gbvPe9hJWhR9PSPZfBBcBdbLIp+fiPdZ05dkPub
DQ80be4OY7BbI3Gy6a5sVKEmE4Rv9zJQfajG5S1VUzrENsIsHEtRmFyiNX2u
oSEpiijIh1fTN8RpH3udl4G43wJCH6FbZTZl7T6SdkA8oHcva4C97bLBZMKX
f2NiMtv4MqqlHxT6rdvmV+S9v30CqweutIbFs/JmSwXEgJ7iLNE3wKlF8UY6
4qRx8zmaIXeV6pfXsN5Lu1D8el4UMvVKnZ85z1kjRI/WHNvyKozqBIiLQ3B8
OF+svKFEs10e1S+Dp7GtEN+3oRIKyd9Mme42DRoyVIZM+8ErFHrFQO3KOp1Z
/Yjsx7vwTRjGNlkW55ZR+Iuf2mH5XJxu6oy/RpKrzN59e7MgXHLty7wghzje
5HM8UaET/kn58E0Za0H6F0ILj/kbzpVJfgVoPSnKC51d99k3+vmbH+wVRGi/
Iqhu2RK7I4DnlphU5DNkHyU3DT6gh3voITsr4Bw77N5oakifT8iPAYb2Q+VM
OiuMYgZkUvORwhYaTexTNc4pcRXTuYdRwtvMImcpAF+cnrbDr5zRxUnRdOeV
P1vZ9s1dnsQtv1qo34MTAJqbFbiJfhWknjsiSw6kbEYtTKqLgqpXC4ANwiSw
BaO7gbs8IGL79ZTIAyEvEvSQyBF3vgayuqTkW266d94FfyhVuE2L/EMUZYaA
Nd9qiZpCI509NXYc7hZ+T7+drs45SRc7IpdVxJ74HIiGJxqG/140pz1/jook
RKM2dFFyqfadgBahdJCWvaqsJ3k2eeXgZTfh0J3IRiFt6qCHkfYNxZAXRcjB
8FVIg8a8KWWil5r9MCOvUmq07q3icoFCk2Ll/cc/Ps8BkYUpOaR4atWzFKNp
5mo0vTk4AboLSaE3ULh44lHJVigBK5stfA7p9OWZPp041gZGinK2bSBhSr+5
QshM6g9iOnibDiLq8XSy3AiE9pDqQi3Q+uLeyVMGBQy+MXc0fjtXIa9OvK+b
dVWhCjoFZpguc/L++xyhVRU4U7TwBqIHSmkLIwlCGa8XNbpTQAX//j6UzgiN
c5xgLoWrCrgni/9tEa54PFLJjM7PUkOA+oK8TEsc/KajmmPgZ7hdaSY4zbcj
ttKB7axJfaHUtOSvWTVmX9p07VwV77El5Sxl0uOfYsZQZv75IeaiqyFvqqnH
1+iaKvIuLoFFOjxzpKeEkzYhUeeRgjGIscvTM3R/9IuTyk27LpXv+gfMzimU
b/dBgUBiY1zr2ODadtVtWmrdifZmfj0xKDtYdxDoDoSG2kebrKbCJ9D4zueQ
6fCx6mCxktntIonh4vb7iVX4A4puht0yGGTfLyspo7EQ4ALmuwq1J7xTQ2Jd
T1J2ryowUXiAO38Vs1TP0/pfg6DWOUMeAa6Ofsz1VbyjZ1cijLYDxp1oLkfx
L7y/DteRNOEIbI+gX7FPLFNstlYAx1gNcW8WKjWgHtvCnWp0Ecpi+5qSzicr
40KHh0GCOKZmZj6rNVhBhow2KMM7fcj1kE58ZKvBrHTAVib78ovogTnWJMmo
ycz3phxVnWitxxvRIz3fDNTYv1JlT+j1EY/4CBxMc3+5PY8/h3p7/BkGKk14
Qsaww+r0JrlWMUQD3YIXX9Hsxo0jDiF5MQX6IU0u6RWL7E7jn8ae/rH4W6+C
fVSto6aIr69FQog9xVGSjzmI54jYqJPz3WqjSi0dPp//RLwvgJFphI9xWBTg
XBNsU/GkyqY21vAoonniVXOZgKfM5IPYe4N5bJ+ci/B7Q5r1SEjTsqW4yAfQ
yoo4wPfxBbzrfhqKlUIhJaNpc0YwXKB2AqfBJ0gIR+z+caWfQynIMeBF9wWJ
xOTBKefSgVVCqrHDbKt3omiAaP2ahukyGOsp0oyNBIkedRLlCldBjMT6Ni9y
C9PQ5VVo9JhsZ4l2Wj9Jrl1RW4UWIUeQiYTq9CoTOp/1UcgkZrA/Bd1bgW+v
77+TOFjBfZK9Xfs7JXTeY+MHN2ejrG6Mim1ut0x+lsNv+0ADiy6HfYFmjQkB
V8bnBG4Nyo+GFQue/a4piX4aOPXqYG56aWaK5Ig6JBmrtZm2N7G5XR+Ujpbd
Sv7ZjZNmcxHoykneBDWTWBuT8IrNWLlX/M9HQZmLqsWXEU3fmdyJkOAZpRQB
zxyP6NhcNCcr7fbg/cYcCDJ+XdbuPbeKUuxwNCqYCzmNV3M1+BmN/nmY+BhH
gFzvQkI1QuRCNX1aZ/261NAQ1W9YHG45BGGSF6RQOL07FxGViS8NaejVeuW1
zw7T0mebk8M+QSKn/fYP/fnZL57oxksFk35CGjaCRS/ncknRao6W2vq7nIts
k07zZAb7QML+3Tg4//7iUaFcHF4e28s1wuLoll6Je2X8hT2Q721Pg/xaAKnw
bDg5Cb9m5mbppQ4df/CwQKfe5fprZWMqcW9TYyKzWvKZRDZHJgfEyVlI3eTZ
A2Ht/bVg9xd3lfAumpAnUSK/5Z2zzZIaQAGn3M/kWXLtX649A+95BP6Y3fCK
COL6Osd5vExht3MVhP6KXgwxe0i5nVYJxodgfTI8Tqu8Ruj1UZSfTf/eRqDR
TDHg6oVQxpLT3WkzibW5tgZ87VpMDicOZ4l4t7SItS8yCV2i+4MSVdNzlaKL
b/VCwnUDQ8t1QSTzOs06bvGm8CaObp+4afGnsjzfR6rzidWVFRHrXLMC13DE
VL1gw6OH9mqHPAq9sJ0tydVBIFK1qtPyGQApF6Xi+RM5nAHI+eFM/Bn2TF94
UzSA+kFFWiMToMBPVDbbD1K1K7u9zEGrDgkgva+brJ9fm2B60OcDaOqCBM0l
wlwfNAadNqpiiDu+iFhiyW4Soi8i/v5ZHVBVLiwFKKmRoN1uhOXqeOv3UKF4
Km6eH7VSjMk9c/SfvsqbV9ywiFGoLXMxIgZLdpI83uLuqfSpxL3d0PnE8Ve5
GgO9hYs8yYeNWvdWcHRSP1D+/RQD+wwaArwPigfnDWFz5NnpooGjJDGhNf9E
qzz0WlURez/dSK1xtXdUieUBSK9odvntyRy7MrFLcfDJSelrhZgycSOEhBni
BNAvcEiELhsvA4JvX1dXvJFfU1WI0rlMYO0V/UIpm58a2ceD2LrwNOlL4j53
8WsHtQCFIFKt0gpq4craXNN3yV+b16GVmERL45Vg5xv834kXZFxzKJHfb7ct
aNG9VrWgon6/wPfa/6+/+/eioL24dv5DSroYnrxJ4jcymr7f9HrzOyUHhShl
/hQCLOZoorbQxOX2N+1WOeX/AwHuXgQUHu/L+lxXjxT3wWNKaxbwchffO567
KYRk4pNLmiZxilwfJUyECZux2ST96phxtRDf30I7uxuXdqEx2RBl6RGaBk0K
p4EqdHLmTbfFkgpwAcDgu2hkRZxPstr3TCbnvqEW7jBLJRWIjtKe2BS15Fsm
2waXRHj+d10jufiQix79Jz4XtGWEGUt3+NhRo2uzQksgVlz3QZJhjwfLbNQD
CoJxz6NEk8X4JqWn7tmozmf8V5dxHN+GkNogbZQpegy5FunQBBqp2S/rvkeq
Rf7eUF/bFLPDZI2Zvm+7K4Z+Y2Z6uSi/D0pAoqVI94hboLtz0YoQdgaQLqQt
650o6TUcFwYgGwNBVbl2oFQ1Ax52wmACBTnefrEQpQ66LQtX0WTdyY2hCX21
CwmrSs41LcEsFfyP4htO+/rjF7NL3nWv3HOQfWsXXMvpUMtwRNLNJWExnyd6
RoqSWoR+gWYKx6LrKY76d0m0lDgXz0tEU8ryLdQOBckLpltYPONkNp6/2jp5
7gTmE/uckwSFpzFKt1sX5ogKA0SEP6Bl6OIpcKSGx8s10dAzxz8FU+RIZshq
ww15hRNFTiz91x8Aygh/G7RZwurUFPLrvNEMV1cgDaFCTvUFH7hNyPrxTl6Y
x/vziHpomPGEdnFTWYAINXg22oo7l0jHrIlgSv0lH6rnBpzEcXD8ead8g8/R
ZM1B5m9PaBBJILZS7fUmryKQqLUpwDuTqtA++5h6pr28ZmA28bw/YY5jpXnh
7j5HvyLEHvPVlIWKu9IP3BIWz/JdWFTBu1QM7aIFWBUM8yq2poXcjFM3UyZ9
ubQILh4IIlzAtAd0ZJbZu6n+L+6OICESmitlTrd/5Fo+kJJBw95heXMT+4M/
R8SLNMyAcgyLBZ04QwiZWr4MuVcxwhhl3/0Nn4lRODJqavZxwi2msfZgZpY5
W3EgTuhH3LzdP1OebMs9FhR5S3x+u9qTYoNfX63Ht4Y9zx1q1KEsycUnhUG7
tQeMhsJOFzdjNitK1fiBbMOXsBmQQ7MSt5bqssh0ABzFlfKntu4eCflGQ3H2
TgAsD5SW7q6sQgYA41L0tZYHznUDt+Da8U3a4XObT9ur5d0wqMQc5Db8cfj6
SiX/PKrVYEKFLYfMD6pVX1zTIRUATUU3hUdtpUNw44ccbUieLi1e7Jr43yhj
aQO3tPWVv+4kiE3C/2ow49p/FqBr0dEApcSewdSvoSCmpib4xMn93h+lBtJR
EVrmkBOgKbw7DsIqY19NguP6cF22QSuPOIz+rMMNjhNIP8r4Ggf87K8/fIi1
mYXKjYqGBbTv2EmXVSKUlPZlGaN18sAfy8vUAKEQSmNkYzvnyxylCkG3AXj7
XAqLhUfCdkqmcQWQ87/V6L1RcUUhm8REYKYyvFJPyOnOPhwJMxH9yk3FzFl2
QbpErLrk9VEiudjwSgIF354NS9VWb1/x003tLXisBGXToo5kLARadOfz9JBJ
/lwyPT9vDPoSb8a89q7bcF2fFd8mKOkEY7MbZWB295WHIIY81KiyGNq0ywZF
L9JKrR/Bwg5uiiOhNXPQx/byh1IfjqthS62R59+ZAcjqkczsohaA57mAfIII
MY+0c4MQZBjDDHgxnowx0UFp9NATMn3EwRU+qs8tpfssTa7iz6mRMaISQzMY
p/WriwFocRM2W1lIMtNcttQTfIQawyEc22QdywaEPbxNJRCcVOsnBHrUanQB
oZxNj8o6LckYwlctZY893exAITgi1jVew7/Figej2popikwpyIwB7kXMdgqF
sOI4xDL19EsmOPQ7XO3zDSKv2n+A4oxobMJNLQ6s0/Xr250AL4swo8QWgJNU
+v8eeyK6fNUkJNTGMqQ/4SwxJ/Et+P4koAeXKQIIbMvDSo/A8yDpIRTv6Gfr
hYGqSY/K9MneLYjwgWrcVKWuOanUIL8kV9kKfXmIwwQXdxE4ZkUjqXx7cGnM
cRIB7IwXXiDVRY3sso/FuXX325tTt7UuTUoMOtNnRF9O2vrRmDLHSz0mlIRr
tofURw7EznMCN4r2IXVQ94rZT4eEY/LmAMLOSEg7ib9fTeCCkBwzgCRx43z4
JCFAGEFyLi2GF3gbCVlLOIcThVyjwxXkOhsWoiU7Y+3suui64+rVk6upG9U+
8+QMBflMRVPI2DQWdlYPmqJ4/O29fOE4GppAItm2NGqkA5FrE7zXuXH+akx9
2NHU1NUIKEfnc8jYInTe4Gcbo+UDOvPn0ozoSfjzZ67gkRB8OStU7HSB/4y0
YQHDPpcsd+M4qCHgM2V41StFESv7p2mzmyNwbtTwlOKifEalDe5eoLxQtSDR
T2+txAbspRvNelOqgZgfMJO3oOtSykBo18JYGplvpv8LP5SYwE7zORkZvINg
/hPPFZuzbqJ6al499UK6ttOIQxFVE/YM6KanlCw4H5sVIYGOq9NFtuA90GVA
6aWNjuhPLoDHtazIM2zmeLgiNAgFXWI+18dEhgwfi/xcC3GPwkYXwd0b7HWq
p6ZIH/W9pXROcHHx2EODXzH9LCT2VGrQOqJeyxvBdxDVps0SJQoIxnSHx0Hi
ygey6bWSmwlRj2sMz2g5ofj5V+xgEgWrlUi67C/5IKxLPlmU74VZZdVBGHUX
ydh2AGQPLCBYpSHA7deIO/kwX85rv2BKqFACpS1M7g82xbblyntOwOccQq1R
eDYeF1ntRQNBjgMwJH5iGCbZjow20eKq/aqCWN2ZIFlMv1Lkkkz9CrcYkaIx
KPmYJ587H8CC6UYtFZURHVkXVixF3XGyIskGYA1vkF6QZCxwu6NbZblAuXCz
/sPhI3HcsoSW9KjiSMFSkxA0TNREtPxcgiFLVSEfkiyLiS5PYHerNTIgUe3Y
Kpdqu6J30f/JJLLWNe/9N+KnC8hkGlhVYyqREh5Xvz0J7kZlW2RQ04YE+Was
2M2kwzJGWihrPzZ3uEvmqpFwNXhQd6cgOZxceRLzYKhD2CYKtcfZVm0DmtQv
gcgbyTQYOKKpMHa+XMEGoi39utkbt2hNzrGE0V3AKIyPBSCZ3Hr1OmpQJecY
iciOxlGjdem9ae8+cWw3Ao651kZYatVcRPKkAKEjWLsMIGZlUiQ2Hba7Tkvw
EAOzwCq5othMTG+SGiLtDrQygAsQLRe5HvdVbhovDzPA0wkMibpVULPkvxr0
nbrM2yWvYv2gi/fIqtGE3sDrI4hroaX4GJlDYZrhbPt/V2GJ2O4snLiYgkw+
GygRFqUKhA+CTneaUmnkNm2BQ1UPRdTXrHXBJof1voiUlpRn59PfmsFtBr/n
Oy3gMZlJD2In2y5hTZbKuX7GGEJjs8vI7YeRiprLoxCibEG+3w6XMrA9jbaq
E2Fy7Lx+trQ0rbq7LjGKjfbxHljDS8q3Y9bLrqpaImJ6KIelWZyeBE5C9aAX
J+a7xpoDjoTwOFnaIDja4987l7dLZzOptwmgchbOcba4NEh+f79l4yMLFWIi
hcTD188hMRDBcSwfwYTIi6PiEYptVOIPYAnkRH8ul5aO2qY97ad2vi3+6GbU
4mQtLC4o/40s3wmrWxfVNAo2TREGBEbZDL0yEq4bkhB25OF3UprO+gWifJ7U
ZmYFTakjL5SM4v5UuTG+n3Sakx13Xvhl30mVOqCx9lCw5AtvUPFPdt/CLOy3
2QR3x1rmeOqNFfPVS/BMFXgjlGTJ3QekJvpVTZCwONboLZU/KKT+v2E5gRwE
i3yO9AS2KEbIrZEvPckHkPgTltKmq3ct4poCh5ixtOiRTPd8M34YcmD+W2Jd
52Lf+5fhO7gVaWwE66BYBkUxK1/IK94HFXMH7h23Ed1afRj7BmMUOTc1JBhM
Evp5BLMWxnPF+LY7Cu81SYLdyrXkvEyju6Sudk7hWQd9OUmhqrzI46HDb38G
SILac/j9KJRnyYyx5O28fHJwerKb8vobgrQyiTNb/g+FyyQzPztyMZidB/t2
NQK0o+A63f8bkVs1oTlIwEqhVLjEdBHFn2hQGol/gJ/OqxpiQefGqq6w++uY
gYtZKeA+2HTMhYSjE6v5a1eA2qerGiUo9Za0jExUW5Jki1Goufo8wo3fWCRN
0+y1g65LyjGM6RpzT8S7jBn1gFJAOzfLlcQHsdGsHHjWPjxArUGddJts/mje
SuLfa7ccTG+x9qIJl+zVej8DsTjYsrSCJIsfYjFMR8uDPoJTBKcU37CLy7qo
l4ROhijRpNkV/lVclXDWu+0CQhXoeABmuyLQYc1TfQ2iA08CxZPwjKUCf0Sp
s0hbWK5xT+Eb7tedgwPchUprosrlJ34hl84o3VkwyTMplsY03IzAigzMGbD6
qpKHXfhhM1txI4qnFRe308myMFwkAY9T/+e249TZ/3qfFI06Ipec/87V85xk
x9gSblmJ8H9yL5WpY5l9f3nPvBwhAeawV4tb76qBNDGs4hn7N/+gPi8+E4iO
NWGr3vky9ARI4so5lq8wKKCLlIuvrpvuWZ2Z9d+1RJnBDN1QHP93dVML6OA0
8kpOC1IrHbXxKSKh14Soi5oxMl/8q/XNSYT+Rapie9Wb/ahwbwgGwxqKUvCd
VqmZ1UhRTV3u3RY/4VtziT0vuRzJzPX7KDB55G7AYL8QroV2/g+hhewlYsyi
O0qF7l7OF2bpXegNrw/PSOMH+RWFjp3pIsKqXwfUgpVlW6jMbtMWGlrVBKlm
e/e/J/uqBwodijCBaFIVPBu+IZ/1090Y3EexaiHsiNSbtTZEWavy2yaw4x5U
aYcZWWCkpfDRBgd21eb2jfrRbwo3NxRqtXbd7KNKYmkJJ7C/Ps9YbTVa1fwn
R1QSk259MSZvh6QmlhOSBPRlsVSMHbcJK+ojhUF5+Wa8RJyQeUe9fAUp+Cbd
fxQT6lXXzEHkHpcZiXIUY1ka7Kcsd9Ru3pI7KbP6EoT7JpAmgfCC9ODMUpA7
Gwq4MngVYOO0CoxPXXunRh8aukQWWlm8/xb2gXo1+mxG3Sy9l4wO1IDaVRGE
lEwu6pTVjkh26FljocshnCnvK5ATA+7YzTzg7SHrL/FE3789zF/yLlQTIW75
qM4dYgg/XkRe6XNlvfTqBsA2dBGF+8vTYJ/AWwuGl0Fac8VUyBhzByqrIyPF
cZjuKjJLcRd0YbtdeGonvumIZdwdqQq2wMkxbLBv51jHfVkwkRtoiDlvxIDH
2DQRxHsO415kYGFNz5Khsk4FFQcYtt+IxmfQ5ebAfTGtfPEnkD/0JWGDJOIE
xCtOoEgKSKK6gfQ6UZkGEH//9J56WXWndItMEmpZtsJYdoPn0AR0kmXhGqeG
FcMoPtGaprKgnLXNOkIQtHE+tCO+4frslYUmQ1ep5NFeR6qgUk0s0tHZkBrT
/9A6NAaMHO0ky/L3Gpe+5aj6/LJ1YOBCYfsozJR2S9o2/rdnshRVv8z2XuEi
8UooGKb0suM/SlOJ6/3xCx9l6h59IwKk16fkvT/ILtSJdEefW0Ow0Tanw2/i
REWsIbZq0KIhdt61A65V0UMGVWrN/D16k0+86Y8kcMiWa2jONxYsI4SxKpam
zyttFekgVPESNhVBdy4lcvqX4V/wWXLMpekKjdvseQ85VT2XFrxATAn4nZbQ
K3lmJbCy1v66edptWsEZ8dGruf3MfsvyOFENQDtcTS0JP8CN84fiCayvp424
rAh8pLABobQPaC4b2PQNWPSvKBxvZ8PrNaJijwW6dBWV7cjdJT/8bTYxwGQe
d1nBff5by8ksiqNfiN4IQy3UE/tpRLB2PCip+TpfvVuCIbET6s3aUMGR4lm8
HIvz5yAhlmDR/kW4TBeoEgq35dipsr/MPz9xJ59qt5LTuqdw8N8VHJ+SJD41
d1Ef38YuFcaapJaTxQEYb6tyXbyYjmeRrui6qKH+xRp7ncbYrvYKieWbfuY7
dhG0zcKNFsF9m6PquQcKY+8D1XGEmdDFJ+SVAn1FVnyx6E/sqlzL1OkA2Fs0
/lmnp9NCtoDSetEmu2zFR9/u78OdAfE0efGSyxH0fqrdFu1FIg+fiUKzSXC1
u4sRrjFZzjVf21LbNUvNrM+DQlfM7Z3cz4KJwnnd8o9nLlTjyRnGJIl7/8li
OlW7WAJpWBf0UOxJbxmjUIinj84r4cKC3+C0aViBJFZdBBePrI5pT6nzfbx5
ZV7LG2BnGIpu2T7m9E6FU4lVIPYeSSWRWEnbR4wUf7PxBpApoYsNXEbqrXfs
aj7yjrWBo5rMNj5z4hkoBzhOPEvBp4Ancxu8n1MtKVmAENlwMbwAHfrXJ5je
wljWKIn0amfLvfP2nKUapLo5KaO1TRZTYLke7xdQTC9a2NnMnFHK48OVOvpp
7AplXim4qJP/YEIS1870UUjNArtU4EPCu74ivi6NAC10weIiKwTNgYOQqEcm
a1JrCWJayVz4p9DTZpdqN4yly3lxpzfHk4d613uEwgmrq+T0DQHEA0t/bDzx
m71QOBtEDB8o+QJ04bZnZadT4/BPTD1PXQx8SSFpnUPq5pZZ6b/K68FdrFrO
6Gudo3FM/b3UCgu+QBFypLEa3Zo1w1Rb7PjYTjNPFMiueca2Cin+ZlDy18qc
hPM4eziQSFvjsEqU6zIAUTWoexzSFvuj1FHSjJx0qH9F+Ckt2OBSfdThbCst
qeUT2+K4Q+9AAh/flz3Wqq82iBf6j2B4fOXk5RkahRs4Cz15FIMjtam/lNWx
BPnwb2z2FXDyjWr4IQovosLJ+vVkrPq864WRiL8GW/Dq/bQRKr7DKH66U5QC
sTgzwUG8izIzsF93eJJMrXzclBfm2/AxILwx9/SKCKwCvm6kF5byRgcdU9HN
0mxxI2m1y2ityVy/PUm3YlE0pBbPP+prJEJxcKEoXfj6ugUUfqq91M4VM3Px
DvHM06EohL0mnIesuQjSSAN2OGYMkFNN5M5D+VENeTJ4IAN9tdmVFvpIHxZZ
f0yQBwZtbw3zgrdGHB7jgM9UOoySwvsm1xjMr2BZ4HGDHYDPlUG9xUF39EqG
5WtYM+CAAGsHrElzQXIbC7VOgQi9m8s39/MgCvI6ApTh4TzG9IgeqRNvtY3Q
O8rX1/5UWpnWwc4ODfIsi8JnIu5xifR087uYqSRkKi3hnDC15zLItAr9k91s
C57UqArl/YJcU+/buEpQ79nRCkG9Xm5o993fJjkwfBMQVbIa5N5LPVl/8R3V
te49AOa02YUnGVmGWdw3aUsONibWXTOmafeTUHKoymy5q8VgqBg/nc0erudu
IIX0kmjXdApKKO4i3GT3yAda1IVtVlt/iFfjHpa+r1WdmqD+vHZFVHovYHp9
4cypTj5RnQkVOasyhlaRnaRoNaVUTfAyyOHCZX1oCV8aHDISKZHrWhBKWOoS
A81+JwERTHgAIoz9dOMSa1HxcRlOn/qdu4HXZcEumUY5b/iSVQKpk6DsA8i4
HQE7qf4MrC10c3M5yn6NiTncxenRf7b9YoGSlKs5H/fOB4z4nughVXU+xSc/
JmBtiomnKU6aHO5YdIrB5hxQjHOLx7xfWFzOpwoyhtbaP3LjdiNfAoVNVwb1
kbajmDsiMy/D69C8OZ74KXLl/na9iuYv/mYE1Psb73hP05a3UxhVILmyN0Rm
rDVBD0CERGAPc25fY+RO/4st6asDcEfD+fkIVO9dlBt7ZIoX/8FDwuFxpQqz
vGBoZozW3p+IeIeQtZ0FGHGbyL9BVnWYAHm6Moxi2jTmm3rbpOjENRgWg9rA
90BBtoyBnYinkj7qr3sZpen+Ur/+x+zBf81tn5KbizlxMzLmuosr61/g7ZI8
xkWLgkJFTkXOQ4xVngMJVNDIu3eeWdOg5+3Nm7G2Ae4GzFOFakQG/ZyFcwW4
vj/Oly+KxMqE2fGC5T9+ny5H/tXUoOCBU86XbCtv815OePMhA8vTLlbSvlE5
h4MnNf/5iRtby4VSny4COHTxM4RBeFBl1YQJCHnS7e9U3G1yh0aw3UnjlBY0
qlXoi8xf2q2CLTsGiCU0t6icUlkPcoS0IHmH1ZlSFP4gQkmN1EsNJaa8ABqm
RHwy88lGVBbQMtQAtZX9WPKQ5MNeoq7gInwnOzystUcffzIWH0zCImoVUH64
KOEflrueRTwNN8BlzV5+Uy7KisXGZ2HRaRa5+iltYGZdO9DXebF9HI0+I3oz
JJt8LzFCG3nMO3A8Jj0kXVk1BU3Ie9z0SGFrur4Qq/h8QFjxMKgFIFa+1atX
Ocdo2CLulUeo29b6wtZIqXqMNNxLJ85kXG8Op/h+cimDuzrclp7LCACfD4ih
r2OhvhtTJZa3ti1COYwkOxlESRqbakZFvUTDPBJPc29b29HidY7bggAru5Tx
hld9dOMMxEQ+8pAGPHSNXiOv2AJWltgUlJ+MY80rID8rdLuqB3K6K2PhKMPo
q4gSH+Y+WtkoAiUoNx1+AB0kiwwQQAHIFgJZ/MRmS4r2WvLq9S5gYk0KW7Fs
xQA+5RonE4izcBG9ZrW4BRoVkQh9ia44zNNcSF+lnF6qVKiaenaFw1nWtBkt
gdlEogT3W+3I6QM2AA+a9ROem0sERAboYLXSVit2575mI1iENyF8sUMbghgv
ORwSFBOjefDC6eTSAPuXw9+k7aukpcfkm+SiL7bH9d9JGh9p2zHCLWaA/Bwl
+E45WFFSGndkaXrSyI2F0wnL5486uoGNbvxTK0x4KFr9IA+Dl5QqVW9hIn/R
nvJInpweU+HfznD7xZtu7KObpmwZjV5yE7aID7ie9O55O/V96whJfw48zMwP
e9pqAvsbwWBte44eBTJq3PgUIjTBEzz5eyCFS5BiWnfRjOXX2OudPEF5ntrc
RtDSSntHfp6qTyFQjhmMqmvig3YQXwYAYdROysblkmjz2/kVEO0p9BDZcGpd
fVFV+dvElvO/Y80pI8pKR7WKN+SP1Ka/bzw8jbGNtoUFsxadTI1Un/6chcbU
il+1FcM1GlzxlQmzBaBCFgBN+yJHLY2lyTS9EPapkM9s0hqIT1YO2EJmLjax
FsImzvsWgowize1WqaRUCSGkhV4htKb5x+CCyYlG5qzFG4Hk2fFyK/Esh02T
GlLohNxgsTXdvdcsX7nsMdNIOxyNKlWJFz6iBX9NtsCyHVSV5RuOEoSiWzYa
erLKpD8ON/il9lEEGx1OyXqtDylBTTXGn+jnHYOBiTTq+BWuwYiFxOgfvyK6
F+u/rrjkUu8yW7Xr0DzPleDtK2R0CEm7ndPTfsRlys14iImKlf0K5MNg1+IU
nlz+b446/wK518pEtAkw3J5hbX9Jt6Q945n4/DSMgKVPDVn9vJvMXv1tdIGW
JIrqE9tPYuGWE5H1lS2ezky8zEVIHIH6FVagfJigZDt5tD2/fL/VkOJQ2Rtj
GSpb/4jSeFBIqN2aDvYudfOB3fMIWNCLEkWlMArQU85f+K5dkF/QekdPGbm8
hRuule/Fg27Z1wYHDbsVDCV2g7kPpzlMsfxJZZEC2tRpvrnuCtoVUXKqINzA
wsX6JBEU36oCJ0jk7lta7ZGG8RkJTEFjAeYyObUezHvW+8ZsIhCh9qtJUyef
C6mRJId7+4+zBaLij0tamcb/3YSXeo7rfYbHcET4eHmImQSbuKx453D9LXtJ
Jqs6ckUYbYkNC/VuNQ18DpI5aflhmDBhF/tIIKvnlfWenZbj3CfCIAl8Tv4e
x62HXHkslX6C0TmFwRkmWcXFqMBDPk1+QlaFIeFOkumMkOdV8O1J51amJt2A
fB71ynqkYFVeQiA50BSXGVpKokhydwRJ7X02uw7CRGBtY2xY1Fx5nEoXS4Tb
XPN5MEkz0zRo5VCDbTptDFwmjLnJRN9nve0kSk1m0mGyjSjCFsNbJS8Ypizi
gEna4QzE/Iu9zi96Bg770I59akJ3WpuF82S0tOgGNlR/xNtT2KfqRHE5wouO
GYmuYET2xLBRbwXvqEDdgpgjV1orFvrJ4MVzggI3YeWFOfLSCsMRQI1sCeAF
ULTxDo6RsiHANu8M2HeXvykkNnyGOorU2W1Es5PBsIhB2FoGhtWBZI3+T3+a
KJDQNHPvFSH9WSUyuLpe2ePcOzzkFuYbtU+RbSsmcH8hi2bgCSE74MFnGLcw
EfW8J7Zzz1QRGY26G7P8/5NYHm41BhK0elD8M1wgKnE0H3B78E/VVcGhi/rh
Pl9AREYgGuaO3TemXWCUGTYMNXkGSC5hFL067N3qo4U8EGQTO+ZzuA3syyUu
RX4POWHl0K9Sr5C4fYolNIpnPlG33945LGf7tOuYdmItl/gtOyRT6ZKsaE1s
paRyblX4TffvcLvSmrlvhaXAaSrClOkbCoQOMjNJxLmV35bh+uUnF1wBcFLA
IyRgynqO/s+BpN/AzAST3/K8ET1oDwGyUR9Za15uUwSiBNMALrYDdur3XXn3
oqRam1fHMxckVLuYJzXbpV+0RFI7ZxSmnCZBragjxKvHlJTsVkZK/gjikpwu
j27A47Q3j9izYZSLFTKYU0EmeBWigZBdimXZaH5pMxHUY7rh2tVPtrtrJBs6
7HD56oM6s67fvxYfl4oOLGGnAnrSiQwLlSuDuxCSww1pf4H8s09/qjsuB6tf
hz0+pqIooVF5f8snEUPrSPXbz0x9E9yRz9evovXMq5KOoQnSPUcEi/lYBYw3
k8O4tBW36gvF3DFPugXtWEHx7mWS9uWH2Dec+hP1zQ6b26mmUwvXPplfY1XZ
pVXU0RUw/CBoAxZUcdwsYl/ncwKeQ6GLP6oT213XHVi1HBo8pCpchHd/HE0O
7UqA9VP/H1QLAXWdkHZLXAsNzl0PbEwvBVxsitX5riFasO0fGpBn1Di9BIJ/
9OMKLmixJSFyfpQOsWBhwoHlHoCJyATb3LQ0xDVakJw3j5CA6fFDHBFjItIU
x58ekGfx0FN8k8pgjFOTqV21ZpNi1ayEuZ51f9CL4qPBFkfETcHT/m/Mg+sM
5MLIcESyX7PE3NMjEY7miZDpS8SCnqcMKmxJ08+5bco9yz/a6IGF5bv3zftm
D0BPvRi+CXf+ut6Dz7Ysble6Om7rmtOQpVr5KDAYopvimtAE85rjXTUKOja/
aoVxBeVo/lJLkkz4D7efTOHHdmuK2vM3rK/MnYra89O2QYdxwr9qVU6Lw6I4
QBpcCmisgGMOBtW9Y2aoNW1me/c+C67/7M7smuAiOLnx3Z6SGG3uL/J0ITj2
+qug/HlR4Yfm2yoiOO0N30V58fqB7ex/IpTXtbkmjFW9fma+J3Oxf+jNxytm
VxFrtDL2gF70waRVbF3OtgYe8Vio/ExU3FnSXC2N8TFXXFGSpTRupsKMp3PC
PpFRSWTBMfhJIakr7IMzUbppqPspGn769xm0OcavW6v86HNzYKB8TH+w06E+
JHb1huYiX6IB515hrLMQkzbN5lVGPi0YA1+OJgAP00y1CMBL41+eW8QDrYtr
h8BGyn830sb08jxvQ5i+G3zeBtcSx9klXinDH9k+uxBV7q66Vi2ZBlpdy6Ui
lMKk/eXkTNt6Q4sc8tbEP02IJzsUjtXxWv4ZZCuYAd51H0L9Rc/4Xn7cT557
rac9zc9+qlXpuZUpFwBJwJIKfCIghMcfozpjztEg+jcCG3j9+jFhU1WweweB
HUP6U7jRBQgbPqeUKqAPxwEaINO4PEQ8m4ErzigQoi8QDOCmfFMS7AANxPoU
lFxH54SWb0uED+dWEx2eelQWgexn3P/oHWMWNeAlFXoyMNJqJcsmECk1rLV/
wOICCvYDQhx4vTdbEypCQ8YDeWunPYtTChBExhRZjmgAs4U4hkPhQMrp6piY
3mk2gwBXwzveRuLEF5lw0Wyixx/gnWiAkm1muCEA+pIEzSjhHZksBqIvO+yL
d2W5ybi0GsPfAYEJ0onj3Iva2IHis1FI+Pn8tDa/cZlrACefnXUm/lNlCEe0
ePcI9rAvEUD0PSXLSn9NUr3AvxzNDQ1g7/tZaChCdNBsWJRlC83E86wMpWa6
yLsKD+nvLRiR9BWSR7NyCnCSvlAsVnrMlxwIRgPQ6yW2hzp63HLyOCe5h4DQ
lpWl1VwFrw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "hmRb1hCms2kg5lxwgzvVC1ojkYPyZtVhUZroYIGDp3nv41l/XQfn8gMXcNw31HDDWBFvru7tQ/av+VlNCOY8CAEc3dS4tSN1iCLWoSLzjcf1An3u0nZDKunxPUWY57wMTkfTn6dFEXYBYGQG/cgNqAwhgy/sA9kmZ+yrzAG/xfCgRlDUR3RpN+hQPPycj5HNM2pIgRPAeD/5T2qj/frBFu5c2+SfDL19Hg79cXZFl7U9a8iYS+SoznTVGe4dEdet0ClO1quTm1gWALJQNzPYv/wv1zKSVmra2JLBiKQ7FgnmWWPACCQAbb2yPZJ6gaZQcjgiZoPLUcp6YBCv5fEhWKHbYZ+4iFwrsuZmFtEZd4uIPsmGjkySgxivamOA+mzHl8iJUxBGRMtM0DzvLhsc4lGnZ9Z9rROLc1HqPTicXLH+8TQltFBfmw+Gax4t+IL897pmKQznhd4r4Nrr8lr7TZ7TNONxZuiqGB2oIopCz0jT+QHBcuWPdmrMUgUVWEhfICJ554kiXLZdd1ULRMKRwUF3BwQNWN2HUtwRWE4KODHTeDOBVq3r+xvjVa8tp6tGiAz1g09PJ6drItrcSWWqw8YFXPihq+NSyUh+jNEfteWYKSb06pSYe9+j2KkEinNFYf2SfpoRahl5xg2eP50sv+SnTfh0wYinfPAnU72pYzQ+gK8DYnIOiTIp1Gp9x2kRvwCXzhTxeXcawhemzdD/8g3sgsInHg4sfcDRhPLZx9l+nBWHJcVUxoLlH21kkT52uSx3WoCgkhYXcyqdFz173v6tJvCdcUi1p5OvS6tyCX1ab3EFtc4gjSU8eKNLaQ2olMzoxOFPg/eLrQ1V/u8LZ+A2ebGhrrntHCX1g50movtcjRP619Abo3brFftSlJFe+SqzdM+tyWfkP13R4DvESJFY2PBbDK5ZpeEgwXJ7L1uxB5kjJghZjnQrV3vWwlq+Xmhl41MNBmT3X4QKyjE/yA05GhWru3aaOLFkUGBfaUEhT1760KZ8UzhJx9CEYCXX"
`endif