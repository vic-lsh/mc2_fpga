// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UuX9xP/vFM059D35U6J5kC4sk91Lfy6HorA7Z4ZNnHnIeAMyDCcy8jrEwVMC
+Rg/agm7LSchDayEXQvVmHAWIpDZJcgP7Xkp79M1Gof88P2jQ/LKk4iJnZI8
388+sUU+bfZdM1W0XepPr1BOTvfO7a5QnbemhMBSRNCoGtxvLiZrfYDwyZgK
KRI8jrlZhvAZeFbXzM7wecuO+wDEGgyHE27/Y/YD1oiR9Hlk3CzCbRvbIFyx
iTNH0bTzJ31+Z30OZQeW+9d0i/FzBux8jclAeGPRWlp1dmxfTv4UXJsFX4av
1k0oGgwO5Glesf7Lltim1Jev0SoFlrC2bNTi+eZxpg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gObbDmAV45B5dZ0rsN9jUJKvqOMAFAFD7CKJ0gnD4PFMF6kz/kt4hZCmxZ9S
QvYYg7Z1QUpcOSWaw8Ulx3rKHSCm3bxQpX4JAwgZs0qHzSlRBGDJ9BVmjr5k
POU/PvoLclqptmBMeAv054iKLnKSWz3aO7tt7AQqNfNOVDkO/pTIPRWS2NSE
BbhmLCxO/m7PM/hGV2GAjD5BwELViMdYq9PWmjutlS0/QTmekaE8faQSC81y
rlPI24Wpnt5H4rPN5WY/apKaUvRN2XzMfvi64BrrJYIsXmE+i86tvVBhUXMT
JJRpapgZ221i6NXpqkMGY5vuGyfIC5ZlwlDFauh78A==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
P4095LgyR/yX1Syl21Xvq36ENYBACQw01wq7GG3fT0gdTn9K6q3oyxqU7nOF
EKr/dAgDQKllKfvYflZuSTgbWABWgcvutABoHpuQ33r2gvcU1UcTl83qF7fW
EwLn/Bw7lzcy/mEY+6oTkxX498ZOZ9BwfAdmadFKn4vhhrDQaAMu2ZJXql29
lif7hKzuu0uZ0XYVi/0Ff8NQHz7zIKsRYc2cxFqaAXfQW8cfyA9ILcVCn9Hz
qFPTHEix3//aUCPRFoz5xtvc2+SU9pFcnKPnKug5cboqP8aQXhj3NbyolFt5
y02ZTlxuT5bvn+k1Tz8O6Wn+t4uChpSSTzu2sia7Vw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jQWxU9ihCzbeBfq2y+6+9qcuJ9IQhfPZ1GxFgL6GiLcqKF3yb+L8D5UmI8vp
1AC0B6fMWZ4lrsyZdIr4pQMgPHjsCDyNFKBuu1gYRrWl1bh3M2bMqYrkn5Q9
Y2HToDEfDm1vKay4LY0p4l8Ninnybt+FDAJ7WssSDc/Fi1mllmplWaxmZuyU
o9lub00vrGCUBwbKFjjYko++5Kn4XJWT0HC8S5cu9jYxpRxgMBpNuCSNeBu0
RHFYWwR89XjeQX/EVD+fU9S2d9eUcuNRRgmQTNILc3VQrgopYDs3TY60Y/Xc
4oUWKovrWG9QTms4LPED94XPpAbEPjaZ3dtxDghmDw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pwCp8xQS3cA6LDqBa3FIVP03LuFVhI6eZinEiKqpmPy90vn724dIW0sxaFjl
tpnYQWo83jOwbrmIKMfAx0oL521qsKB8kx34So9mYn9WqSyD/m1sOJDWM+7Q
M43zGVKMKRZHOB421BqkgfTh+2Di6L8qaeXTmhwoZscVDM9Y4Ik=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
s6J9h4X7+6vRfwYUOEinTBFvVAtWzxuQD8dq4W0EA8ggNtsY7P0HiCdzW/iY
Cpe2WYxjL3IJ6LccEuheaf5KVXqVtDr1kA1suOlQg3k/gczsGNtKjMMA4SNz
haw4vvSzYcdgI+7tba+MDkKC8+m/HNAbz+ZnYoEauO/dFiBks2X5J4kb0IVX
TyQf3AIPz3/6b+ZfsByr+GTBEqcJ3vEIqBY5HeYIMO1eUR76D7Pny1h/xko2
WbPhMUY9PgApOQrSGzD8M85cgYBmHeWX3TAqzFxjKI9bDYhiFtjznKU7ibAA
/pSAXIBhANc/gLnaIx6HHhS6MjK3CbvCIY4NoA52e8somVlvdbKcEzpzldee
0Hi2yeTkfmxA7/oQ2O/lomExLsjshX4KcjeXqa+FQP3cEgjrID9VO2TO11lb
CeqiS+Ls5k+tmcb/CkRThC9aE5RDeKA+3AklFjPbSNBBZ03uj8QkZY38D13+
xDT2jLeNbv3wXuUtqvgo3keTdSOimeGJ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dnkxWuXJ6GGs2uAnGJhrKOIWZzG/Ga51FRBetyBfsZZUuqeygY5gc3W0O8iS
7Kb7TZijG2TGYQn0Q+DAKWk0a1sBE+n28A+3pv2sHxZn3X7DLzEi4tn47Rao
4EyU+O8IbJtmhm3GfG6KPJ2uDDkK5m5iLII/dZUAGg3IV6bVwdk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
afJ1RNXlLOD59NZ6DmNSeKGxrVusl0R5zpiXwqhUc+q/0BbJ0Q8UBVMAbbEB
ihqJXsRrGNjsQJjLdAC5QGxlNXI86Obnsp7FjtL38DMMOh0l0DjPPloRlGNX
gOFTWk4ndlwRSBKPYoGoUxiGkew0UNOZU3tzqjstyEL0QLsmk9I=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8416)
`pragma protect data_block
LQ0sx3gTQbwLMxsWZ2rD3+y8boH4qSymanyKCc6OxMiFbJjMd4dy4rNEPBAn
jGZqTnHJl/ejKInYB/KhoSpS/tIT95ifsZcvRekkXG0UMeWUS5Y/T4keIXEs
cEIQbYL0JEpiZKgPZNZUytH4DojhmMEdWVrm386mnyZN7279S9z4ntcBji+e
jOsWX2FE3wM77s//AM7uv9KhgnTZKYcHlkD+GRZwhT3ADjD0BNPy6zRoamSv
ETUaKbQmyy4lOa6aqGxqgSB6h9gPCxzVKafvb3yv8huD1AMGx6SXCwP+zjJF
jEJirNyr6N3/PlQ2dRCGoUQkNamMqmr6Nwf1YqEjavR2rcoZkgDY7p65Zx00
Gh1zgtJF//J0DL8bX2I+6lhBamywLm/eI2/IkFurbTXXbT6bT/H3h9NDMcyV
iBn1j0DSaHxHl96fO8T2vydnMYiJN81PmAH/tY4JGqvoJCBryXr2g2UMEafP
/QlcfOUE2TfjIieR753NgZiOgsuGAmJGQqwSX/8p5ZhLjCtb/7SArRmzo1fS
NvXXYhSbFQSaoKLDNrQqifXkA5N2VOtNwqRnF7SfFqGjyxCJWK8HmTgYtp5R
uYGWbLUB080i5vE2V7Z+Wu4qokE0V8FHKvfy9LgVwaS47IMFrdStowJX+aHO
mF1v37RjTaAgaEoTt1lcCBBFjP2qS2f3q3Up7pveiQFD09nnJ+EWRGoyysRh
FTaFtBa4hHKxjZpEWDFjf/te0vyz4ezwg9zyr0puM03Gc0Km1H8a3A4BD6uF
sWrtnP8izjaPjfaOKfXGRic6yegpRmbvBkFB+Au3S4WxUJYVE9cggBAatxNc
i+ZPiyyFcoflaU7jdQq4iWKuNaAW3AWNWPpQfjYrocD4yZ5QUIS3oESfjJ4F
5g3ZtegYq6fXfo9f7dQkh5yCTJW8BICI5SU+gA6/icGoc0BRimP2BYHzTVjd
N95jNWklwjsdyWs6nROkQz/5gvJ7V1bFXeBJPO8MRaCr0PmLdkMMKlZWrjFA
GmXh40BOJ+5UHWN+QCVhcE2i4xlIVm+Ccn9DnpbHAzkkKdVGQGanxmIEayJw
EttuaCroewl1ugBMmmd081t9KD97EmLHTQJ3gqiR02NXttGvTtE/7Ddc7BrG
gLS1Ytv8vsBhVgEV1Q3CzSLZyooixLLhQahfUoDwbKmocMGPOvDnOB8G+Y0S
//8cMxnaqecGtsqopKfoCpmHcWwKzI2Tlla9ZgfmGNrMzDPjtZr9r4Cu1Xfp
5cLJDnKt8QbT7zxWBIlSPowJl+Xjg510qF13kBrU2Atr6kXbbzA4kb+Mw75w
Ioj/JbAWlEDxYvyD8sU3Y6eTUpvlLHBQfUVfk0AlND5ZlfnJwk9VF7uvEpEu
ZCvAFOIxOQ8hpEu2JUdqB6NrEJJyjWrpgV5+mTUXb5OT3ykmw4TJ72n5ysJI
to/gBuM0C74gxndw9jCmcVubA5zbGH0scsO7US61Yu0gPfe9eTxbOPbvpKxf
EsB9inlYuXcqFNPC9CaDnnIURVedvySo2sXio3D/9+EMkkFitqSYCTuuAMYr
FGpC/Dv6nqpq58XnMK84C2Gz9DzCHw2pghnk7ybBWvX1wOfeHREtQw1aVq4o
/vblGPrv0adYa52GxS4n0aowHR17dX5wOS+XCmPaiPumFDJijW06tMLoxGHP
a5Gb+b6W3Ng+5SenNHTapdFUaLt2j83XjDcPY3hoejh/nCobOABRZGQXS3v4
kRdYRiLzzQ3ENd2Ikhxfp3z3owvstsFnNy4WtY96GnujkgXiL8fhnpnfs0eP
9343nV8MJ2azNFK+4qtVgiJSTEM4rHEfAFaMYpWraMfjforYFoOEJ7o+Bl0m
q2CrtOTd7K2hT184I45UHXAXAMQc7zP41B5hNPsYjJosFwGWn8AE4jIZPZfw
z0T41zhrc6Ns3zXlTJPDX3stcNacqSfyRgw+d2RfDUK2K6XXmDIScQmMkJrL
DCx5zkQ73zM0EegL0zRLLQ33l5ag8/BDPCj2ZWnrVOkDGNqQFovbPGeuPn1M
uuHoT+rNgojMv5cX4MgJ3UoaHKvX3siOgKfC/pu5j87PCG1WmJrsJG1dy4LU
6r2IswtzktkEeG11dL8xVQ6PQ5X5RKwrY7D3E/5tz9xD7l5A5Iwb1ViS2Syw
2erEfPr+CStSHctBI6s9I+x/nz9pREt9ciMNW5Y+SAMd+M0o8kNv4k9EFgfq
5Y5q1oKVclUKRvIvHeTk9TINPQ1hqqN3ffMDN9Pwdk1d/FHF7o8xVjgA0LdF
saYUvgLORSFlU9zv1g1pWNjd62arck7/TLd06Hu99qA07JlrLMF95iGuh1qL
6o7rHpxDUP0jAMkhL/QTsvyH60lj3IJIKNS0ipsJ/NHhSqef+zUGAmS1FnN4
lpgDsaIRu1Nh5k5RYFqq3j4zwOk4qpcbvGlxft/fvkvRcNbt1XXd27Sf8hAL
vorO4c224+SVWft5W6w+x2kg/NAthrtg1+lf7C5hr9gSkrCEggw+6FzuJdac
OoPQRwNH1SgedzIgpYD717YM70qFtgcUx0DoLQtOzLVmaTzAx8BHzXrtfmVF
IoHMJ/9FVKN6+BO0k0Ea2grGh9uvSMRffaP/J2MDMTuOCHuEnkRY/urqSN2s
75WAN6kLL0yduPAQXaHxL2ymRz/QJq24oJTHF0f4AARCdP8dAABCKOvBvCxh
wdpndcelJhxam0uhMhrPmLkty9DR2XU1N1p5/D5IjsXi0PxEAIvbghkygzf+
4LVK0U01rIrE5uUgdH9DihczX3PWEVswg26NAu+Q/dv7npjz/IFBrChmaui5
mDBQMGBiP/fILVUrQLfKppEabmU3lKHYhslmGnMGKUg10x2p4xHGV34IxBnV
ZiBRk5VRBNR+zrd4uZFvim4E7YYepaNhXellxT2xHwT2nAGaFXTlqr6HHSD9
b0lLdcHgOnXbcz8VMnwSDfJQpKBmhRrC/WCXnYPwdBGfr6dFIPwp93D/8xZf
UCJuxiqF1nt9f7IpK3Y8Yizfw4NtecNi7rBxms0U20Q3qrlkNPPLd6D5XSEY
lnSEJ0ZDUVioSxWJOW6JQzdApLdFSTyJJZNi9GdZhCcctl7rkfrXeaxE/2Kk
JIHEPC8JotbVCwvFet6+huVaTAWrwvU+nY4vFu0nZbaE/9b08VkCTDL4xmnK
hpOZhIeRAkmSXWLTxiDywEGPs6A+kj38kQpyvr3OqR8UJ8s13q7qnQC7j5tA
Ihy1u92uTGrNzNjyK1M1indbdDfFgSd98pR2nV3PiIIeNIeGTOCcEQoNLVsQ
cDz7SWbT8214Cx6lFIjEl1yt5W6wNUpe0cn4WGggTgKlFohlddvW6CFqC3++
5hKKmEA++fE2mxkiTT1WNg4CeZy83vB5bESvXrlVotd6UmAUs+TTuX63Z5Ew
mtZIk86txoImg2ur1hEuURqGUNs8fekONk9xWyd9aFXVoiRLkJRpvCADmG53
TzFn/p2P66I4ATc8t0WnUjsEkUzzVP441tENhoPfq7PNTqDt41eV2Nz+R9HW
ljtcNKOzO3KXI+JP0DmRShS/VK3R6R5q/AgRXGYTc4HcEVycgMziYqTsKIFe
xmEl7sb4dKoSPXku62HTvuDUOwewJpNJiYrwrRp/KBt3mVQS3LjWd+qqS3Rq
5ugasnHdCL0JeX4Rt3iAIwn00ueAWw6CVESrkKB4hxVEu/88cYssnOMLH+2r
VutBW+rg8gfvhhtsjpvEyyFXkQZi9y99l0dKu1jKAalsqQD+qr3xGJY0v9St
IDwfQ8QcZasF54bVuclZTv0NBbRf+9ZspCcFYQy71amOP/uWxwrdVwNv6ehq
AdS6RQqezYc64RDVPg35rZKb61daMH5S5cTnbal6EOT+zlRJG3aSKGWLxl7s
wCZItATu7EoXhfm3FMO+KU74mDUmL7aGKffZXsk+xWra8CSiSaBSukeMtPdj
XQhhjkBCAc7YFUMHBbTzZKUZNCFJNZlEY1X48HAFhbaZjnV8aXU/J3r7NVzp
/6kBLRTJ0DFMlp2baafBxfXFSS6ezdnFcxpGQtpJZPztjmgogz7URkfK8vaF
DNXDiubWJ1gCJHuSSwKYLGaXUnFbFS/mnagkd8qxnaSad4KGho8IzwpkrCJ9
HSiRfXG+RtILHibgEvDQibVtIqHT0v/Hiq2SRJ/mdC6fXb47u5KWqusB0CNP
1/fUSz+PdwHE9c6K6bLz0jKn5+Ha3oRJpBbqTGJH4Gpv/U79y1kShbCYTfK0
Wx0820+qVJgUqGGLIzgCupHrQNssV9r91jnF/wdmPoQHRvixsg3HyqfbkVN/
bnBNcwOCt2glaLsVZaRbSAsWYGIXM+TkCY8mo07RSNFqNK7feTyiU2HMEzvO
ChFrsDGq3fF0J24pXPslPus0sM7voLLtlZEv32KMKsb4WAlmtMJcb1WaXlRX
LkZaVBzOTo8XtyVfG9h5Ez/E+fEzV8cfFIY09OsmoadfzRpdAD4zSWeY3ZCT
ZUwbhKAmSuejSJpiW2X5FR/mMaZ7DqOvBDITWkvDXwxz9MhqP9ksn1k2ArlU
Xukc0wycqzc8dBcw37pEEJLgHF2qhw7tin/h+r2dtV9k7JiCiB59vSTxcEKT
PuT07VuXFvZ1pNJnF4pSLTetLy7uc5ktm5b8Qy03yGMUqnWeR4GmvwtCriKj
b4IgrwSxMf7JDM1T/Nqgeb6lMQ1nHdtZSbEfCGaTexfpUjT9C4BZkt8ld/GQ
NTb250LaXgJPDcBH7618UdJJRDN7/SmAKlhOGgdnaj7x45M70COq+G7f9SpO
3ospaL+BiIYFb0PHFoirweVIGX16flnB/Z/j9yVX9qLyN7rYGzl5Q8S5dT2p
T5BIhekBjvTe+8fyhTWPX2jmkvz0SLsRo8q8n0Od1dfginXdTuz2Ne3YCEoS
flBY/904rd59EFlMtXkz4rOCG6weL25e6DXOeMECbP5n/wLHuMfwhrNOkCz2
2f2UjVLV9sisugsfFmbub2WvEZrKxX7BFjVR8/eBCPLniWV/yXVFv1xRMy4P
Jg64tGIyGaVyr6cjQB4yYnrx0Qo5rfw5jSvWHP/t/mg/hoORAz9B310lybc2
z/ZbmEvoejNC7NEwso3m9dVBxho7Z33LmiNPkKJ+iJe4dltZxVBfApXSuYtc
qYun7sXx9jbE4xZ5pi4FWNidcVB7Y453jX/J2ixdkoMbjUm7IoaDwaCxFsIp
6vyWMcTEOl34tXXJEQk1Xh7Jrc/0mmsZefJ1buYnrp8VYdi8ccc3ZWt1x3kM
S1ndRiAP3lmHV83jiG1KhGP2d6y5PjfqgtBoEMgJZxvpR109KOqcKUqzBe+S
xffquDVLqbSZKA32/sYdkFIi6jFBrXpLb2Uu319oouga/JX3eyc/qE4PNC42
Rg7B7lv/0Qg+fBD1MXJ0FyUVnV9oLe2cwZGWybnjicuHS123h3sHEVMUsk9K
LuAhP6C4+pIBIibuZoDb+R1WHJ+F8N9E8wNcU2ckIxqUUasFI7m4ZQCp8Wxq
oytIpe2I4ThfxtZ/MEFECnPzplshRAWnCWe5znFQMma8UcEg2W0DShL3ETYG
IglXffrOzL2FGBmmM1xhVp1xxACFXz919ycrZPJZYpIcdpankNXPMDFBwxiL
qpqCIlgYL9kLA0W7wQ5fPHY2HQGoWXNsNQExJL9EMipMbrImHiL5G2RyUACj
mvemXDdxrYfpyJblOKMDL2j3D/Ga+54M2W11IfYvQ2l7J/bY6Lk527mDVVp5
2Dp2jhfJljJlBGXYeWx/YSBbonTZ+bBF9pLj+vqOANuZnXNd/5RaOlg2qcPu
FaF7Z4i2S1cC9LeclvPjBce83XImOQUb0M6Wl1epbC6WU1JhgMrHTMIpSrrR
4u4JXlNo9GizO9UOUHV67La/QWjFXUwyx2qKDHUI9GGZr89m9Y4GbuRxaAPi
YtDFuyes5aN0Y+kx5H7Fra78s4FLfCxmrZrEL4DuIRKsDDLUZ0uRVdYazOJy
o+zPp4drVK/YNxwwKGVFQHioaLfrCi/1IbxWOT9JaLiXLqzuY+LwVZ/DbgBJ
dIsPeQPzzNZ4Rn2J2i6RkMbA0NbYhxTh4/bhPy2s3f7DoB1YP4uS3iZ9rAjF
j3GUwrunlGiQ+BfOBCKg2vxjkMmv8apm7KIk3p8gGqbOM0u+NpZ+FR8mX0mV
E/em7SbJRFkoJ9Io5V5kgk5JcMRz3LplgKMyUFCw3x4pG4gAugoxXit3tPYC
qonrWMKO0gScOErjPwLaU6guPSwXA/uwQORHL53f9Nn2OrWGbKoefitveiwc
5u76gzq0UxNNTIuQcY+55DBuEhj6eWtAUDuF5pbe+/PAf5Yq6RpwG188Aamr
8ZB/CgN44BjjDKAUV2dZYQ/7NbJw7QOErcVNFabE4dDImDfmnhTJxZQt/9wj
7EL0PC0c8eL4hRIOgtuCDBEGQ2nkShNUQ6oJheIh8JwnaNbSsh8xwRBbiEj7
wxTrRx/tee8EvO4dw4cDw/XWP8UMPhirM0WJIxoffsvvsDiBLTlr3llm0h7e
ZqWOwLaQdZatjsCA4PIGmn0PbCNGpamlYBtTYJcnWGdWh9Hh8tbJxnnEfW9p
TxhzgcFRcgYtTB3kJC/fndN/JJMvG0p1blDR696uhntvdDRbjxlq4DeJkwk8
/y0eHGqL0jyKxmFTLFKDKqkwG7uoZlqE7gXKdVyzbm6wJfOk6QaMRvgY1Hrb
NQas+rCHPMBM9P2Deo3mncJ2iiB1zRTLvZxh3MWaEuxv9jxAfyxSvkyZhJ5M
Q4AW0YDy5+bZS3BNI1Tbv88w2hxquYLTgYa0fXJO85zwzU8UmUdp7SUpu7/X
iFp8eAJsAD+Yr2Bsmf+WvJ0+9QFRkLoerbi/bqcYynKR/2GynYaKNgWPNG0F
yYitpDS31mXlqxaL7DKM5gyJKnLjgUkLsmX6FKyHPeOMyD+I21ddFr3rVLGy
hUoaM5CSQIOiAT6ZvPq3d0fqwFUlF2QeMyjQ8lxnTcG6xL8t7RT7esTFnv5y
wFJ1Dbz3AHPT9YmjLjWyVwhdR/EuLDkiykNo54zQQ1j6Oj+TjKd0e6jwNTMp
HKTID+CYRtSm+lTqBo2SZnoabrOHcz4/v9XuN8ua864lrj8ddueI5h358h8Q
uFmc04Y3css0s5+v5T4Mv6RkSsWEtaSvk33SrHp8vsdy9BE8Je0cVg50/zhc
IjzzWmu8UlTyuUezKuwJhtEveCe6QDUQrl1Qe2QvuDZURStQKMwRAd0B1qkG
Q9mpANFLFmi4bQTBj+9KPeeqoy33nOrd/M1/S3f7ZnHxFUcXElz2gPxOM3nS
JExxZ62VzU8rpR2E6I1Bkk2dcNzz61NFnj/4WssNxN7Rot1fKJKheZS/GjM2
YxGO/WUG29ir6Sc0RtrCn/MrPO8gUstwaFGEIx06dBpVBL0Bx06JnqnHQmJW
9mvvz4N3tGPSr99xg9eraY80DIP9PEger0UbU9T1ZRroMFEbRQ7oGADfBogB
bgBA33OVEJ6Vmph5m9McOjhsMVHTjKsQ2DlOEhFmb4ueMHjvD3FmUshGPxH9
MWz3cIA/MzAN5jnImbDb99Ei27tIWlbQJC8qU8BuGID7Aq/3evxpnBMNNFl1
GlQXH721F6k3GXnNZivX/SUHIaiUvLPLF39p8DxDQ7ml5LAZxMbIkGucCgzS
smpVoLvF1VWAsw1nG4NRxrRBqIxn27vHtMeMIdi+VBid9S/dJIWphG1yllqF
Skh9SSgT6OUyBcBzSm27CKs37H+eO35lPocbMvHJKe4VTyeWjYuzK8SkbPvK
j4IWjKyAf2NwopPE/OBvKsS+oKNQVzbYUGVg/ZmgfMAlYJx9OXUJAJQi3eap
tArhZ6GXFhQngJxGPf7KbLVQurnP5k/OEMMvZLQ+g3uQo+4yYme0Qyt32aE0
rqJzh4VcBG1wXdR92Ot/GjSnBGKfykpLM+1cXrorb4jKlJabDbww+xfF7HLs
eo8f1bP+fv4PEHbXHVWSX42egLu4LyVEg6tbptW7Y/f4czNEgqLZQyrYmDSv
5NbMz3pSWv2EEv9b+aiQTfwGCx7ARQAH+TYfPZeFiprnsUW3yUVbrquDbMLC
R+cnuF29G8P23uZKD5C3L15PnbVZJgyYn4Il791t0y40OMgaJh7PDC/64hJW
xpRItAJiMjnHRopiue3K2mp+4m0odCNWA4libXW4NPCYSgvvHIe6vqIKwjmg
+/PkLAoQVdlWVHmMwV/ndZv1XQ4CP/8A95LFR4lUEw6+/H7WElwyWverkOAj
YmlIfaD5JtM46XTNFmykW8Ht+3pzEKQutZkfhsfvQn2/oEijJXREdiITImSp
yl1nNHJvOptrDkSEW7X020Exj9cyD/cC/kKU68Jlf5fg2d2SbIRUiiX0nvys
JtTLy8dGq7vz4CMXS2lhzPPK3wO0udrVNz4El6/q43gtg8lVpGJlDigcdTpb
L997/3oMznuwtfW54SX3xsPurOaqccxuRFJfAnJKYzGNFGEewrjbKWhsqquC
dUDaCDfaw2H1nU8B53sFAmFZNCaPsTfYcTHLroexgztApMGYKWRb6SnaZfzI
iOPRWY40g8aU9uZhUbq7ysZG7cy+QftgR5Y4E5cGVQSxskKl7/eu/UsVMxXR
Rttpc3gXTnWc5CqtZ+KSiVnw9fMLkG9Bketm65Wsdx/uKyGPikYJfNcEvAM0
3GnIcWhijlcxTW8Gjw191V4W8NxQwqulZza4WSNleBMSmuZluVPhvgam4LlC
qqo/AKh/70tmwHc+bIOPiXogw5SaBqO1LOMOns+9+LEauXsgFjRmGYyOXgj9
w98fchyjhESp+ikVKRUZeINcbtWZSY+xJQmsV9u3jBNIU5DXUTChwhQR2n1t
D9O7kMtNqftgVH0SmqF27HJLbmsbMrOGJ2e/8Rq8UgLNkYXvzVK84ddPUpCW
TjX6W3BrcwStcWN2Rgo3trWMTEaVTCc6BT/eJ8Vi+DJlEvPlNObHkpPNspo/
0pGNp6DKih1Uc8vu3/Va9VnxszyE6o3guOkZQcdUoqqP02RdNRtKnzXSgyjx
9/Osa8kQJCbqdR1AdQg7oM1hoH2jZsxrYfmpJypZtt6em7+K35HBrg7pLh8j
XJrEsarskaSExGL6tuyzqSiSDuF4fry2SxwQNGUv0uf0je7IJ7AleebnSnp6
tOmNKO8okXQdiPdQ89YvWShaqUsVnRABk4dG2qm7aRBpq9PAM9+DshUdHOAC
bitHDDEYoFWpx7Yk5fpP17CcgxMbJRD3FrrxI6oE64KQ9dbML+Xmff/Ko0EY
PLiVncnCDQQLg0tLTqO7+W2mqeRhfbmN2olF292ptS2/qxzBDnYTabnhKG7I
LrjpFfXs9l338C+9vHOiWKGJV6sBe4224/5E78KuzYzTyNYpnnnerHTBtITO
yK4kJRV0wXf52bvCQKatdMxmArYAZ+wqlcpNpD4kO4d6xSbyN1jeRmM6is4I
YcfLkDLlzn9dhRm5roPrBqKz1dcnSFA6wuZEMf2Szko1MUFGcd6P2tTRXxjY
Wrn1OHhO41nEuD+c7hDLXjWnJ51BxS75PtJi0dFoPvD9ZI03a1GMBse/YIoz
mG/seuYgpzMed8cHmwbuD9MpG2gBu7FJCexP1qNSfQB7RZ4Y5RHtCs/rojrp
7UX7ZBd8N6StUIjZzF3seg8R88Gt8wNoFD4ze3oXrK7IdCWgTT29R2lEPgTm
2dZWFOP7Maowez5L0/VNHAM9w9l7An/AgDP/EK6NQNlZkmnCL6cCcrx8IicU
jEjicImGgtSHqBdhCwLdmHmWHWizi8zDnwFfbAqblZ1uNdS2J/pKsgjlU19Z
FDBRdAu0eJ0EjaHPy9ttkrfgwfl1n0kKuqbuRk+w1JNxjkkgROPUVhtHIjQL
EFuzwYe46QdV2lhnObimsDjx2Jb6+yCKBMYgHvbV0EDeu1PnJncfeUhaoqje
RDunJl4ETqCaWflHUxDQ+XyHL3RRzXTQdSVS0weDUXiwD6sXKqYUlALkJIF1
xDyFs05USzuCQ69LMbcChWWVugDxo7AbMTVeyQ6E7hEXFnqlLhhwgSQplWPz
TS2G3xhyQayerimNQaEZCS3+nkSnwADSFQJlEbQWQrWCij3M15BkAxJmMhWd
GtJr7O9CDcRDozgMUYgqm4RVzuAfFAPerp3lF+dgjO/gUDQXEQqKhQuYrfYH
QWhatwfb46IM99/hzT2DnLglT1kNktSwsiDzUpqyMKfVFcm8PehHYa6euMNi
HdDwZRNz3z2X7EyhWjclzc6sWLXqBC2I3Vq93ZURIqYpPm8bMgMs7v4pff+S
rJYsWAGaTjjdkTSPPxn7QTEd991Ek/8pBRUvD/5hjqjyUW/Wefvm25YODhJ0
VPrFwA8tO+SdQrBrTWfs7gGs6v0xuQYi8CFXeC5DCdcCx9Pvp9gkPxH5EepG
DfYfM5HDGqVlUjAUZQq4/bhU0XmQbP+Ob3TGWEaNukmVte3eEf88avmFMbns
REf0b+xh7naTBXwtzEc8t5dVJ5bHpCE8PdtX+ExFGLQT+bIvReeitQIFtleW
YJNuHCPXUyCrkab1d7sZVqF/ZTJ/cjQE/tdJs8CetjFIHi+FIdPpIXj2INHR
30GRoM5l/MYeu+3p/XR9QyCWn6MZPY4lH7U2rYluo0f4XGCkeey3WG/O8Y8W
NGrOKCyaXG3/2bfNgIPzS2UILArLljERc3eDBkkNbhWXcxh0/s/Ru+xh7G/N
xQq/oyry9v1gxm0736aKXSa6+bCeREUKmfBt5GmdgTYSGWycH/UouwSdHEC6
IXUHn818U3j7mLyDiEklw60xuZ2n0VvmeRXy34vtSoZoV+lf+CAhECPfCJhC
ndYCIFt9S1MxDojX/og2aVrhPYlYdi/OW11STxi+0qymmINP/4hgztcYENG9
EMUqVtGpAMG+xa1gwFfsw1Mf9fUi6EMwDHLwFsXQvWbIBSlTk5zZs8tZlgNQ
v/BniBto+VEPpbk+PS5qaEfcYaZxmQhkeaJGv6uCtgRBwjRB+LUwIXt/r9tp
bqNsZHLNRWKA4HookkKFfrJUpQAVsxPfjZlqp+MRr5+OkY0+s3cdD46JUCPp
pWGWFGH9FMxSgzWRKcyIAEOdNiMG1iYfEvOdVy7VNAgyVZrBm0sUw/ZLjNp7
8LCHYXWnrdm1eybBEXIOCLwInMikXI9efxS43qFt+NZXvS88X3PfBWjpbSf6
iw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "sTlVzHE+yhAN9Vt4a+7yJC9Gw9bfBRq6xv9kCe7Ng5psJnHruz9VrHCdetev/ZiPTJdBJQmffKsGhcT8C1xHmtnWp2phLrsA++mCi6ZvsisBHsXsEe07/2w+B8eMNZubT3xnRLX8hyEfcYoWZpsP3M1DFemdUhSKGBtblrC5P70SnbNX6tsPF3y1BZk1iC/CtfkXVJdvvd+neDISHf8HMgQ3zyVqVVLAWr5Qxk5Q0qRIs90INLMNC1WIPjPjVxIj73PA6Mw1Uv9gVUnfaIT/i2XvEQ52aTkGejr94vTjAMOpp9EvLv1veonvbDZXxeBW8rpB9EJH1r0+QLNmeFQLy0uYzc4ign4CX4FeviJwgi3oLAdCLWAUzmfhIMWLv6bXR8VH6zOwGdNEv7WH9xk7jeHpNFAiI5edJZnqGd7TpDuutsVSYu2bZjDkCi/m9y/JeX8XiQu8SR6x5wryQkfBDJikTGkFwVN7NXVQAfuXnjebigdbEp5Zfey16WTFUkrWlCe7zkF/1KjnBawPo2U4TTUvlWjxYfxUab2Y6fOn2E+MLtFM43R1fY8aj5EtugUZP95W1QrAFtUHUgo3XPDNQT0sli6ZedLe4n3w91TSSihS5OCm1jIMMbhezsFma0rlOxy/tHWq3eIzXFgTRrulBii0K5vFsggkp/K+kZ64n5HIMIWnff952qtwgTiKJS7UbfgbG8rPUGdoz70aOmSFqgpj9Tbumw+0/Ro7rpXH0N9w0oGQmtUoBfR8GHfELOm+m4K47DZXw0aW/nzrsiMyHrj4iyINOSQ/CrUwE0hBQM0yINunaZGEMDvmxjd3ZaYLirSsReuACnMVLlW15UuVNlfhT7JsgZwf16tilqMdDBetEdzbYIjEYFVjdyzq+O29mWYu2KekmIz0e9r55+noMBffMuqDk+7txKzZ5ZH2/fgg4hOHbyAeW23jz4TwA+8uPQ6NoLC9jGE+ILbWfETejZPv9FrS/zG73CB0EjHtsLaGYB4mJPwIBBefkD0Douod"
`endif