// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Tpo/NKx4I7Zm9tAfDXW8DRZiYlWkdjjNON4Tt9SngCiwsUMoVyYbbCf7V7DI
Z3t+MNsOn4N/RzujZXg4aes3AFSiEwM+q8aMS++M4SCKVpa0xRefdj/khb4X
BD/a+sbEIlL/oMKUbeZy5ZV2c/J/Monoru6QVuijIJk/4Z3i2+wMG7nvHOTg
l0XUDyAU4RbxKf2cDJMcYAn7TU1ippX/viQt8gWnzyJhg1neIEguhw4Ei/jq
JI2bXNbQJVR92MY7ZAHsrttTzHHf5utTnZtwcCJY+TBMAF49PHJqJj/oXyZa
YkJsFg1i8p3gnhNEphRSxWGp4U6pMLWltIvpnoy2RA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
anCiM1fm9e/+UH1AGKf7wo9Z+sPwLcqKVofaYVghzM9t634J34pTjB2BO/zD
gIXz4nNz04rEmTtba7OOvHE3AJD3Nn2pLDKq3cLoJItSk6XjNDpw6q/6IvnC
QJt9cTrtt8MvJZ8qlNV+Rwhqc5OQnt9OLpwXsNekp19b8SKhFIsFeWbSlA0/
DilIOa8NxJ3fCAvo4+3yXcSB9gls7IuS4Y0AEdD9N07l59bDvL3RS0dC4kiv
vqxxu9+jXkbSGHcN2blBw3NEuzJj5fFL2Q4gC+Ci3H0ZcV56vkJHrb7qmC75
Ymx9Ld7l1heHeCrQ15M31U8FPIUROyvEpK19JUHkMg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GRDS+nHXm0QdcFi/2apJiJ2g++sTDmWB1xtzBwQe7v4CWlxNRo9d7iuKiqG2
LQprlTXNvR1pX8pedcRVxCG4JhypLvmP+JeqPPNY9Y5ccdtfRQ9Wz4mNI1JA
0QTnqlZznU+mz/Hr3oBAX61zQmwY8y2KllG2ZdmQUvxtXrguGihcTPCmq9xz
9A/XSiBEy8IdOgrPErN/TwAQSEMXrWRhZDCde7elz5/hsWNoicsfh6AL6z2j
JeVn44CDd9dPPJ5iBSEs2g4BFy6nnVCy6InUk5QYsiaXJaywqoq6iAHdncRS
F+4gn7CQ8iDFETHmlkexnsl0yc6K4yK+p0ar11zFwQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
K7xsBCld/HvMIVoHYBDCI1n5AZWF0QV/eXWN8YWkRTn9P5wUU6vqQTOj2kWG
qWNjLgV+kQGiFfdvf+h8z6SoqlRbNygystMZGnkcKzdnsPxqE4ikzXBLs2tN
IpjjfW+3UphqQi5nJVPdDvN8niCn3dWuZYoDlTiMSt6HhczttHXFCxTELprP
DHd+1Muxn4g1Gu8GE2yBqR30kanmMIK7DHUfM5+x14M85Tafg1vSQJF4+2J6
Aub/yoQDd5BciBxMZAhBXqDoDqFuo8JcehatomIZhGQUr7nvILrlkxLOR6aZ
PiLKQFdT84F4YMWjfliXLkVjyKAngS4tAW1OTeh2+w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iO0vngqUUFuDRcii6mf/tNxcalmXA6Pg4CGhT1RSgEpyuFy2mYNP2Lgaw+VF
9RnnzGejIF26WssSuQsOIzZWql5Lqh5t9EcwkD1y+29twINwc6qnVyZ5Phck
zXOiCLhlTOu4O+nXuE5JAwwUnGMhYWnqop8QLMrjN5BOaoVm4Mc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
wbunzhi5sQtMeWnNWZi8Uyx5uDfbdaZqfX5I4idLM88pCRQc9atkgjKKj6sf
2rhmMEfvpOpZdoEKx/Kyk7t35mmPs1DF/NAEeJ9eTLoXgmM5jHIhGDUfZfyR
mQwLe7p7iF0OG4Di1+K7L6BZMpBPGDcNsg7P2s93R8yI5mGBoeq8ei+K5rSz
ZoyiM0jtY99BSc2nn1Q8n6HKAs9pdFq6Ai47A4+0eXxZDL1/HyA5u+WU9WyN
UuZOo+gbw4ZQJ5165k+FpOpMgherX9Imi7jO1T0uaNiGbDFpR8DnFGtJYfvk
atz3gNQuVT8vfAlT4BTiMP8+7s/sYVNzJ+kPX0R1Ik5I2OYjT0fxeG7nJyG9
pu0sysZeHi2bDxqB4RK3kZQxFxVZ1w8fTfMUgIdNCVmh2ZTqiuYpCmnf8USj
PiO8hslKmcMX5MVOr3LD7KR7bOYZU4JLVxgHgQlPZAagewYOqUnSYzpjEFNq
2o9L8m4KpR8iPt4AT5djxcmmhBdtKzJC


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aA7zDgWPo4YyAuIxwu5y5NybjB0svTfab9g+7y6AUKN+4p1ZoapaODGN49Gh
vaCktAgw+Zw0sVq+Zv2eVrXsVGv66JbC2/oWUbtWVmPcn3m+jMuulbrIKdae
WSo3kXsJqpmBrfEB2okJmPscU/veZKgccccFsDQmQyipUGLqXdI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
j95xflSwDzxoVV+HKeHbYe8LTKsy/umFMm7fMrfvJ8ZVAJsMf/6yYlrwMpfz
fLgWU2QlUetLJWAzC+vcJoyb5PTtowKpPQv2sq4tK8N8VhsFowvOZmkQW5uo
fC3VwdnEyzuXAJibOvhcCPPgcghWahmc6cKHZwz93SjsGo3WDO0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1360)
`pragma protect data_block
/z/BtYSOhC6KTI0Qcb4EcDTV4hlf6rYe/vnRuTu2tmZGu14h6WlYq2YtYHtR
w9H5yQpX6M2C2LTyhWb2VX6Z8dT3fVtUjlf2tBmfbXkq6PikzUB/w02bO76M
wVX1iHkEyOmamMjwEECDiGm/1RntMgrEPGVklzivXu0z2F1+mLbxJTC/v+QT
WlzPChszUtkrw29fWZTgOnXSyu+II+8hdBBW8V0SI4w+n3QABwzgqX81UAul
2XJdIX3VDZch4uoJNGFAeH2niHwVTuVG9Vckk2fwoFLwSdediciV/dKTi6ZJ
ZozT3VUdpfAAlYCVWboj0CqmMwQ7Wb97s5SiPek9NtJ/m9T5nY1ITOMnK7pu
Dei2WjN25zm6jKAfeGUxlZuI712xQ9b+2I4cexZS3wey3FVfPm7ELynCPwGF
jRZsnaSvw6ipnfdMLupiXcf/z/QBm2u5kwYq88H1qP9dZXLoDmL5r/cOPRFL
0nH2TXjrskQAo1fsWcrI3ig/V2+vJGdQHWWQDD8US3tRyBKpYYtQOACP1+qC
3hwb33s5D1skx425Ub/kUUSLduFLEN4KerIAII1rxv5WrJQ2RwvaBTr8ahO4
0MuGU7v3lrzFIaT0a8Y3JCrP6L16IO0133/vlSugvrqsOTYndJ3a6ZLKlE9s
97tswNsAH1wkTjQGxP5BsSNSA3030N6U5xmSd2zdVQ91BXovsnoFglNoBtk0
sjpNSuH1cDiSaTzaqHWNfbuwwiNllfRbwO9PmH5+CzZaob0PsuiWo1CVNOp8
Z6+re2iNWjN5oKgQlS1FweXwTUf6Crfcm2L+lJx5UkME1VK/jMVRf5MY9YCo
UHp69fcE37oZhHge0jpHQ066aV4yDcawzdYqdhOR1qtDiSjWJncOvv7Z76Av
O94tMKBZ313PO4l8WRA1hk3jFisKJnXaoVHyiGvYDAGeikMWEaLuUeJzhwrx
WjBA5xPog4l2rrem4lZcHqnARZtNhv6a0y4WmnO10WMK5CNfaNCEzNLCbHXl
LDzGb7gyAVYeicYdEcS+13yH34nQNSLX/KbKA/h79yx5TQmGPyC8gaEoRo0D
GyyQMOrnkBBksBzKl44HBIRzV7MyrQ5u5LvVtgPGedlZWWAMb7ZOMMteQcrc
2D7AqHxrk242Ejp8QPHGapBIx0eyn/RER//xyIYuLtXThbhzBlRcfL0yUarT
R8wsG8rvKaJG1okOEQYRD9u3G9K6EcW03xXYkVlvD+n4kuOSdzAgCWzP/sGE
iLIC5qDJmhtMqNYibSMOHjkLckOb0/VMjuTSDuVvBde2Bd9mqBq2emYZQTxq
sInvTrXgB5VtEL7EfLYQmwX0CVntglATgqAsoISyyX+jQZ39j7niM3pIESkB
o4L0bdZZ7S/cMPO0I4vPHI7DoPuQhzEvbov1QIU9qL12JCff2PtNVB2fpdO8
W6l03+6W8g5MXBoQNldgWAfh0l1A/r4hPCc7LF+7KbJl+qExsiid+AlkiZRm
V6t86dteFWdW1P7DkC7l7foHmpqaImLrTica3PbcMQ+b8vL3IW89jWlNG0FK
qd3unnp7kNg8UhJIQv7PhvF7qfJUpKW9OYupslLUajj1/kUV0saznFvETzOk
NKOUMDxwr6/Fl/Dc3DE6YvlgEJSWejVUY/8P+rGne5p3MCOE+bDgCCsrlAPi
dSc6y28RBivtdgXMXYQG8aSIzi8L9QtcyakII7TOkLxWiUX3YJ/MWgYAZbr0
FnLEZLCNwZPaLJPZDKhk9wjMq+WgUAvEvMr61bxMQJQDe7sdbG6P1pdSGCUE
N2cbJMycDYhbXw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqdASsIE+freJABvVgrKeECBfjFq5+qcXNjaqkF1qywrEfALVp0UO7uc/4OvZK5x2c48jchvMM1ZMtSfRqh1IrPuqEUs2F+eBUHZMOalDZdpo8BZfACmAcpkSEqUvmjR2uI2iA4NB8+jctNoqN5B5pMvS6yjpNYGMhS3HOJMEpBqay6ffutUa8MfDj5on0fdE8TBFnpeUJHd0LXHLb7dnE5UNurPxDsLL4HKIN8kt++1Xs/Ntpz2D+A8wBkNIPEsr12WmqZ0hBW7ApHdGIKbvFiqL48ACBJJdXXQJE28zoBeHcLbkfES2wElVj21WTt6SylWbbE+USUSYWHr0NR6KWi8XZwXugYdDgMc+Agi5kB6VRUEPcektodN51Ka+T88Qn+Tgkn8111I4tab+l0nIV9IDKePEZCCNolhMv6D9CYvE+96eFDYfaIbKMqx+tHZNopeiwjQtwGzGwsaPaPSM+TodN8GyvzW9ApOXqs8ufj0x6IPKM52dC3HWyTsWVyyQLdezl/7K+pWigmM72hLx8kAwd52CqNf4CDY4EknnBDRIiC+9UDQUZTc/u32WJFJR4lvklkXzOwYidw+psKwELtGpOTE9sLP47iHzi45/M6B9zgHQPQtJI89gqeNh2LRQqMfJf9q5EBk0/+MaWsySbXBu2DvXbybSXjlrgv9OzivN6+OhPOiEmk687ZGI1p0Rde5m2zJEoOcybpJDKOGPGd22Cp96RnQtiEh8ddZpBzfoIWG7PayIStr/qkvtXCjiZZthWlY/mnd7hpDs8zIsErr"
`endif