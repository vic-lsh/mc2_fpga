// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Bdo4w7cLlA2o1bLDgkpuvND60LMF2tuFTj0jHCwQh+VmKf/mDEj8q7cEXWru
KycHr4iOSAgScfeCFS/6oX/WbQFPwP9b7QDORf8RRAaxSuh/T10CHDg8KEQ2
+I53qA7aouqRq6B3+atatiiM8m2EMa07VjfN2w48OJUS1eR4GYGjhZcTPJzH
+8015xm+sN0WNE/oY+dWPMqI/A3q+U0o4aZmCBi6r6XXC4iVOAaNPVKk3JhO
sEbXMLoV3EsctVClWC5xrt6XRT7BE0ptPyZYtvTB+nydcJ+d/e40ikiDBwgJ
pfuvq4ObDgzDNRL+JziSGh0K43oSkgSVG3/eUKlR1w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
K7CQ29mCalPGMSr5kZCCuVDvNyVWZ3+BHVLkTRelGyUpGos2PfPq60zCH5Qq
XnGGxA36W6olSDwv0CWmAlHeB8syAMtP0pX7OFY5bgkdmdOe1nlLNTd7qAJA
+DnRuzAPBGQ2qEy0h1WtLm6zI57a7iskhR3hbLkFm+3NcAYFJkxt+haryMej
Hk8I6q+sSBiauPu7nIfWhd6r9LzdMF7r1ydksrnLKAebrZVyRBsu15VVSM/q
AJ/8W+/9tMgSG8A7EgR5uTh/Eg8GVdDmhiwSi6Dpq03BbOB1XvScUFlf8b6l
YGwVoQp3ahKZrDC6wNg6V1Lx0QmxWZajKL6HoDOT2Q==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jeykebbIfoZsiZe2fCFR8QKlN1f4fvW7mZED+k8eJNR67nr7qjK83W2DR6QJ
BGttbklduQ+Fl2oxyozTTx7GiQE56dGJjwICSZnUg48Bb8ryafNDSdp5GDoW
dSgTxOD+dfrz7U8lx6QaVBZdfR+/M56/WQiFT/I/MQb8VJChsZgoPwMXfifk
GsKtJELKC2RGvCIGf094Ct+yBs4IeQVWul4f3aaqnI5/tySCQxy5B7tGoqdz
diRroLP/TPa4CIV3dn1XW1lV8SkF3QscZxu97/MHNMr+93mEL04GyBbwpDQi
RuW9tD4qOqFdG7fbrIhYzSTzVSyP6c5TEpwU66V3vw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EEMtExo8jnaJeEJV2jEZReEMTTByg+3cHpVM6/mPz9G9ZTO0Okadqwlwd0TD
54B5PpzkRQJZ2jiNSSEy3EgOLFdg45fH6Og6rzH9Gb1U3WTABYGAi9diuRap
LsW/pjt/knqFfgeGWRNJE5i8xAdTCg/hvqJyxWGYoctYZ1VVcifbbTu0dvyZ
mF5RwSpmTYdP1mOeV/M5QA4l8DTIGYXswglXI+OIEQs07WYkyW0V6spekMzL
mo0RQzr7xyVv5AxVRjmrzmOPKXC5gQP9D3fkmOkHftK86Vf1VHFur7mseIQF
7IP7e0DVPnE6Qm/8sNdihRxj1WOHE1Q+DMOmXofSqw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
e88f8lckxcZBtzl4ZcBY+IJjq3l6tAlLzdj3DoO8RCgVq0PXMoav2ff80a67
k8TAi+MqqcU8h3CPA2qI11jxnavYpi849UAgveC9k0jkG4H3Eht14rUU1RMW
NUj9f35kc0xijEfMc0cL/N8giRCMBjaTE7+VMeSVRtEVGWjfSPE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
A5WTrTPNcl8ReD3mrhKQNeru5g3USEK2lVXDKMMpFV5EWKnKLTT5qLpKX1jx
iRF81kPW1lzRQpqIs3k1cvCHpeqQaWCTe/K9qVvLsY9MjBz4MC36zFmrCFPf
Y8EmTuarexA0N+kc/dlgT8DR/a/IDK+aHwlJLJksjOmD43br0wrgcmJiFXlT
yE4K8TVvuvhxUL3+d+leEhwr5N8m8bRquYtw+RLxMfqGz3ZyxN6jaOQ5ymoD
wvkFx2WKfgNjivrcBHTvUViKLVAtwsmxvF1Yr5pCMJKgNPI1Wz7XqLetbs7a
cUGL+4MvBbb+g0gytqd74v1Dq27634o8h3DDCOIBA/gTHWNSDHH5J3j4cGgq
bE7JQW8uDmk/QIRUaVgJTYkbNryrYaIARaiWBgTsRDRb+5ZuvTfUL2iTaMy0
UKsm6hzn0Qd1dY+ULEvZLbTERZDhxtX5uKg2nt6wxTaLMmeYBOn9c2aDBlTa
XKNf9RN+BRAFNJIyDCXyasrsPWUmrrsO


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uFJ9XZvM8qk02zTL8Ywz4a138jonnf/CxNFnhOlZAbmy/XxqxVpxNT498Cn+
/H/HEA2wRfO8rYYciuZoOsbduNzhCMpIpoir6cawUQvtNLl6qy/+hPzgAiFF
7jvKg/o5vKKBiWNIw0JrTiMDJV+43INAv3kqLRw6YAovFkjYtXY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Uo0TLC+22Lq00BM0ekkIp4AdDMHup5sFTJ9CB/MBmsHAYbCg891YYn1p2Wlt
CYT0IQe4reN/vdnO1BNAqjWyrCnqblDrwMPqjVUvhyDzqwoFJvykYGJbUqFS
Vh+STYt7pIW+F5PYkXTxNaEcoWZGoRJQG3pergc4nvWmM/MWPzA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 32352)
`pragma protect data_block
fXR4rDyYkFsq44B7vKrk3LpqX8IrkYcSxK23Xu1cd2nSfFjWG3pU6Ihhvsgu
G80/jCCRLCReW35BAfJEpdaX+j/JyKGFmdJ5/qoLuC+e67Y0BQ8kgikSVqeL
jFq2R80eVRyuPBkPckyIaC6L+PCJenOYAdn/ACAbZKLJ1JGU6bGQjAakTXMk
zr1/1Avh7QtH8rhuY2+pSoyjdfXx+3chjfW+xyT5fB6ua6vgWRsVqyqQklcZ
KezDJShBL/++zsEBJnD5msW4iPvTjNhjMNw/QpRFbzBUeQ388HWDQi7MdjZq
Xe/L5YPcsqr54vMUZoPHlh4Ztfv0Mc8NzrM9W9Wv4qKrzBhSapojQ5moa13K
P5WxILQzr8mxnMrVSu/xxshmHOQrPzzblZk4sC7ffd+A2FN42CWV4cT2N/UK
4p2scP8GA3GUSwAkLls0Nt1XieJ1IuFo5DSRtLQEsAP3Sh8UmrBch8KmXzCD
0LCLobUnqBUXEKiGlkPal2W/MZ03OHHEDeuJyB/XM2Kw1XeBxqrEbSkJURue
aj+OWE6DetCyzvg6X1hHCpl2khvyZPNDgD3hWKA9cAHJHy0ktqo95JAw+SZy
Exie0DE4g/AvjUamivgAkuIziuS96XQZgpvOOIuILn3FefuJQ+KX3G6y7STy
6v+gvixSaTbLpoO1CXta8SIDD/lHy2ffHEndLNW7KIUZwR044AO8EYbgAH4c
hgOaA87T2BrAwVlGKU8CsI+72GC2I5reDiY8j/0zar3HwTzwWQwXNy5ZWQWt
gw1SL8evuKPF+6kdXgZP37h7mEUgENhWyjoxHhTQ73X7PsXaPGAjae/Qptcr
2u2ITrhDMIU/yRCRGDbguK1MgeM6M8ncuxAklsX284tjoOTUtAYG8pR4/CJ+
DRrWxd55xD6R78M0JJZcvBVmwyf434kPQ4qC0AIMfr6lnlAnQDLbAxD+hMUc
gZvnmVTi03HHFzMt+4LV1xVs/vrCrjRZPeiTJ7AKQ1OTu3v2mYHyjq7ybP5K
etYgnbxcoPnoecH9P+2AJjrGdKb1ZnGpge87EhYRJ4L1QTxsGLZRkGP1tpfr
UdVPkNFJeOxmtTSjP7GXIy7I6JDQNf64T96qrgYbBkokxf+jpcNybZdPTy62
QxCcEIwsoMnrGqt3w+3Y/UAH4op2AXTU+36xn6PVtH8bDfm9YuOR36p4fF5v
jyZB1/iyaQf2gzIA9Hb1UxyOZyTE2mymZkJWEsusHzn057V73RPYLQEskPC2
yg1Tsl7NwShcUbVTidqWRyG55SWxZGd+ly1v0IBY3+7CEebixMZUjYWltUaH
WR+piMwEHn3ESLCYd1jbBOiXVVPFwHwLuNOmCSq9TKwG6Rv7rVcXvucxrFyD
UR9YGcOei8bLJ/f0xbldhBuGh0HUgbbfSIdyXw5WCmuSX449OUTjSXGd1Uu8
rBBOMjIGnMqnhRuoI0wH6YT2E/9hZ3rs6oX/QioTketCg4S6uzFvIonBjknr
XglOMcsYzAd2pbGwC6Tn905N9xdg0DFe7Y5k5GnYaXstEie3UiSfTnVMu6K5
jlnQEFyznbzGNCt7ML0Wz5mhr4QCX8l/qoCcjKJhElfi1dM7W5cgKujVHrj1
q/Lv4T/MhALz+2jjDuhqknPStrZkkYlbe0dWPP7jhW9zo2QvJu7ozjeOTOsh
u1MXNVjduGDv1Rutp71bjaXGCAQqMScye+RV52tyOWLTVb9Ec8gaunnJkEGL
AwORBQgWsk8UevbGhOT2OQ0XoJ6uXsEwQpRq89fdO0tZJGYVe/8/AYlMgpBS
12FYR83NHvRHeGMvYylaD+SMisU91LIga/KSkCJ3VsU4kKfeLDSD/Kp4IPPj
MGby444uf9qPQEEGAGnfRkalP66wNY3bdi55NatKLMWe5JxQPHEp1pl9nBnX
N6Uf/rUiHcrprqSurJ10+MttBf8lQ/FnOFHzHYf09dqvMQYFp4iZhdkGBLVy
I1vGSptvL4rZLjiHgB99V3v4mHS7HsDzPff5JzZJ+Q/qOiMBm1iJiyPK5m9L
4AZkbn932kNid1PpquePWstWkm1PfnI13iryT2TDd3qTb8Bx9yvChuyA1J6G
d2l+SjwQrl8P4fjpneDD0ZrgTcjaDV4uWSRkgYBj+oFwffvCzhV8oigiSYYd
calXSTtxKdfeQahYrPUxhAdU+cx05JzusOS2Q1K6WC9IYrDgKfm3vdgqlQqY
H8FdGkjKTFbfSc9oskW4M8VHgn/QjyNjjJDo3dMvhP23MQy75Mlr0lLW14RR
J5KG9OTXSgx71i0uoM0yI6w7xw7MxWUUlUn2y8YKGlaKQ+b7bNfKIqkpZ3hm
p6ksQ939kTjuPvLoWJFhcab9sgiENKW7nMdObQRCeKb8ZO9qSTyFqaaFV5yU
4/2XlbrS6DXmrK+9iHOnKOqasKYeUj5lJZvxvx5i2selBsCKNvBAX21nenIK
5eAHeN2ppMDePjxKNWPRqKDUbE4aBakbalLWvd0qP6pYrOwA5X7Bxgsfi61C
Bbez+QjwwCU1ImeIzJOt9j9+JDYM6DlLIEcOUBSmD/WcEtZJznu6JQBMIROk
SwukM3FM0NklNLOxNz/2CO5uXOq2FoiKe4l9KNKhSLsmdMnJZcYcEODnQAqW
c32BJOWxRMyQ7fjnVVBZodMVKaf2ZxZvDngWzqfNCaQGnAnUCFC8fDMJRhdu
QLjmx5anlNUAELPgPYPzO/v7gmPMfd04FMa5oqqSEqNiIrDAOLMeK7Nrzk8G
XurqjmFey3K2Yhw26YVuqq25ryk2yeMfssMV0Wvp70A4o8VvXFbVIk3VYt/r
WTIQ2if0xa8LUsisQxAtpWOjivo4J5aHwb5kg1xJJQCZIqK0hwq13S76BDSI
dg7XCALhBe3broLmTbL+qSU5JxAWyB6/PJZVnWjnx73dNCZUzIy7mCi+N4g9
rymnE05bQPwkrTjvh6MBZsgGEk+O5ob37J8tZrb0O/7tLxEDehcdbbG2b8m9
wymeOKOiY6L5qa96jQOcChfnYJ5ivNVbWUHCLpF+YZk4YaJDztdBLx10Y72M
wRos12TS87COOtqftntEq6AqFhMVZZ/dlU+tpwbEwc+g9ziARdJYZCfsxBZY
Ki6s309zU05KX42gBymDTfVp1g4rg5MPE+mDrK72pJ+joPrMB2oDRywF21S3
plQdr4hNDgQdagJZpxBRYixKAN1T7pRxMeYDflq1TwPSx4asNW5yTzbJGvaq
zjeidGdhqO/H0XKv1RRBvvHFVCOyv26h6ewdUC/QubDTy2CJemYKSaS8AsO0
7WFBmms5NyE6od2zuFNxPavOiXRxU/uRupzj3CDtsP+4R3ZRsX0wXxdna+SD
FPFfzeucR4szebecFv54SkqdAfSkE8BqWvj2STrq0WrjFBX8s5VTUI7j64Dl
tSkc5WRoE2iCIzijtoZzucsxHq6MVJqiskVRxGW/yn6GdGZ89pctO9lVAP4z
hzB5XKxLKUZ2/bv4fEa740w8q3Xgqh1OP6K7IcUY3WX1QMJXsLrn1vCq2DX1
24Nh9s/bDjrO2mwVwfGNXJ70yDhiwr6o2zlXC42r848EYAHwSyLjPkeSHVTd
MKbF96+7Cj+OteSPcv9agMPFnxtegHZK1ZdZhT1xU1MzlJjzTuFZN17rr0Za
MKGDYgS0uDE8Q0mhtddO1uFTBlQsFYvB7/GJtKQj1IsmV9pg9uG1Dg2AQ168
9GVf2PFa/Ith0smD26GTnU93rb7wZ8AJQw7cBtXQ1OmQzvvrguc8SmYxx7bi
UTulFjnRwcUXiKgSUmDPXzXLmWQXLl5zEvaKMGHkTlV4PB5Xnt37d1NFjhCq
iIKkFMp7lsh35JEqc9fAH5Makt6HroX1+gGkW3ykOpI4v/RdSrNcJYpJsc9G
/eSGBNur5Gnk4/OIqNjKj4mQ/Bx6w3jaejdBoM1KdR/DcUVQG9PICcJuXMA8
6i+8HqWsm2KXsA06fmDA6LCZzuDxOGRGs2xW+3eCUtidaue7/b+8+ghLJnwV
1BabVhNB0lzlz4pcCDe6rxFB9ytIFV0Yrue/F9KVeHoC838WyzPyXy0fsi3H
J8WQjvJ22WXvXMMte+VfYWCQyvcNzuZoB5sAem99YBKpqfptni0VdyJ3Os+F
w91Stf39fxKWlmkqN/edjjq/eCLCVQqjFyOoMKhoSmPb3K5RttcJhJBwcSnR
giHSXMDTdpRKTFP0glA6DNZwoQ8NpqWSfYMTyPHovkeX/99yo0LshXmWV71r
yDzLzDJ05ViBL3N0Wcp2ZNmVB2Ch8V51a39i2FbmQd4+65LIRqI+U/mJkE2O
8RCzHK1sHTJ0PGxlCf1LhmNCIFdfXCdKH0pElkt9RX5SDu4AetNogKoYCmx/
7XVvtZLFhruVRaB0eE7lXE+Upkde364VZlOw8LRJrM7k5gJF3asBVk9Whu6A
tcRNoFLgi6FZCDFL07HrTMvgUmbd2k5fYSuQNJTC1ID4uNvdsOJxSdmlbWuG
uEssnZ+GGm477xR14x8+z+Y8tfsKgp4ZPkTDENqEtAzon5Zrjwsu4a34iTnJ
QIg7fCofCVP4tkhvHYhw8nnTDc/dpSWC4eW29CpI3ycrspotRzoUF2f+7TSO
Ssg1OZVarjim5BEjyOZMPR9Gfp2bMHta7DUCJwemTYyw4yqZR3Mi1Qfbj4bF
1Nly51MES9fHaiuo+2DJNX4yGj8VkVQZSlx4c6E0UXiaxCk4J4L+dYRsUJx7
38V1kBHvGtWwCKS6xxbRc1JUX5HnlFbnbq5MzvZoIDSwzeOJRvskbNNTzn4N
CYJWpu82U/PkUwU9/rrDwuZxwLuH9DoavcBrg2kWbbjTO6knFzP9DgK1Eil/
3AeqJ4crUGOVW9yCzH5z0i7cjy33Guagn3Rz99hwBJuPZKCTeLP3guvr3//w
ncPEnjdsMvhkrWqPx0F8NTDU3GX2sFMHUSE4oKXB5+Ii3UkVzFjxLjGGjzp1
He+gByAoM7m49CrDWmGHo0TmDM0mQyecQqrmIXahtAXt0O9oMPzizKZzdIMe
Q3/nJX8ljVdm2CJajHgmDJ2CFuw+2JnxLHtBoOCeszBz9zLY+JMTsDJcSv9N
LETK6y/W4jPol+OdfcOk+ehEf9m+Ln4z5o32vXl93P3bIzGhNIkzvVQ3Rz3+
tI/r+iWpdBVbWb1ChvhiIb4ZLNOdCdlOCNN4rmKz8ufvUGPSZ1xhO5fkvV4H
FPnIfwRlGupAbJzzIHk4K1cFFWrkynAFYUZPxHMAok2oe/P7YmGzEhwKuAVI
7tvD4fwJRBtytbRNpxugPdTSGZhtGKIYogf1lhrcvQhFhvODomTEG8ObRdru
rvsr5AXbhk2oUOKiU8dFGs++I6rdOZdts9we4rwiLh7/d7Stj6Ef/+pTDe9L
O8Xc4QLqQrdcpe7OmCp6K16e3yqnxyHkxyInPD4ueuRA7pmrpB5wAT8LqtXr
kkv9ECUg5MDESq1fsJ7hggns8oh0aQcl0xBTSWsSH9Vgbyqb7kq9DZkyUVVl
/EJJME7qpN63l2elM1pPKHwgKEeVO3q3HtUYS2pQFYvYu8BW2zx8NkbFEVPT
R8oB4XYglvRskVtmkGVPBnBwQtUQeO6wtv3cGSArRAwFfn4PMyjDhGp7ASAl
9iReDNtSEU1k0dT3MX9/wop3y0LGPOAiT5TELieXAFX2blWkwzlBy8wU248S
ZChUPzHVdSkl0tiw1N2HuXao/+pIF9ng8i+dxXmnHhxB2BejrkLUups2OBTb
78WErgsreF84KsT5MxnZc6EL/lx6KVB+KpgJJmVIOEWl2qoCCN7w2bkQDqIw
ShpBTM92P9IlPeEsOfTxmL93hygSefjYFs6lBpfdEL7rN/e6JK7Q73dzC+Bj
NPZS+jpqexRsNwjW5uIs5vnPZaqZyBTT7BOtb/R6DqJt3JGHfibvHq+od6CI
KZxau0Qcbe1uesfTb4ryTAjMojM9FX8phsCVuB1QG18qRfFAaDa6iR3HS03o
ctR/rme2AR9V/01ukA4tWRxraRgYi2T607IDu5hFd9P91zWHiTH/9v8QnxrT
AYywOVbl+/mozPtmt88xBLFuhatBRpKM5II9MdtrFCef7MlOhvEqa8R7xkb1
BvhqxFI0tDF6i8Wm+Jz8WCflcdcWHrhxalxGv69hbde379O2ITBObm81B6Db
Z5SHwtjbedeaHnNouomzq7aeRp+uWQBPQYsg0L94FWm/hrJN9Qti4z7yqDXP
pnAzpQvrW9qczOJBdt/lLi/1KsoitSWqtUSDFPLMR7awNBwXFlGl3OAnCe5Z
QY1APwcN3qTRrE5Zr16nSnwcPvMPc9qkBnB7UJ4zQhaEebxCUieZpaxHlMVz
EFbzbM0KG5+ddeLOGklL4W/i0Z4OCLONSVrI8ReTVpP5iH2oE2ef8C6KoKZI
O832oJxWIcAiS2XrE7Udbo3+AQss0TYnrC4sPP0whAfKUSG2c/RDPPVJnIRg
SJGLfhYMhNNLQE/zKTAimUXdQqOIe70ZdrdUKz30/uroutD8c3Xlj6K1ql1V
TDdEyse1GVVp2vyIzFFLtXETjZs2ygfqC9clMw3DKo5j5Fr3BblZaeZmsSud
J88jhd63ZvGm8oImKxYX/Up0BX4ZzZDLsvqZZacvX6tT/3JSvrDyqUpolJbn
ImPOok/AqgOC7CXYYN+E+GBaAq4wdK/NWUmJb575/kIpZ5TaCy4mfmobV1pO
Q0H/d4QvOGzASmuqliYqwlRDbjfppwp6/pF2ec2yuF905vrvHC263v78tiqr
sAVD1X4MDl89P065YmaLaFtOmrP1Tg67KtKczoTq9y+dSTwbkfNWbxPtLsYw
aM1CsImatENv+LuJb0RsxTqlWELwEbdmoBVZIbAXAvWtg3ZH+MYUGmDWfwOj
z/A5Xz8SMSb2pgNBT8CM9NKroHTY1v0uN+rvkH99ZLZ9WJ8w2kEBpxnQEAuh
YaS3PuC8IoVGigccygRzJ6EmRZr2BPOOuLwaWnC4YK3+Kccqhud8ODOpWy72
yoFalOYoZqluRroHFDKyh5OqFvGCb/PnmLfpNHj0NpNi6gTHFndV1bikxLQ6
OBqSAQplORjS63osFEIr2sHTmTWgyqmTlH7arcpAjUJV+cfGMJUZSLUKZTdv
eGCvoLpWU5Mbge6ATUZtgEsqs8Kh5DkOV5I8xyI2JuUgXkxLOO15EUy3XXFe
DDpCV4fNdfrhIgoLM1p2JdAA5FA43m+ncQn1uxIc1TSkX+4mYZ6MIbILlqPA
yjuynyfNqnDEl2NrN8yy/qT2tk+s1thGy1T6tr6IyCh/7vVru+P8jO0HWxDl
INmVIIYT7Odvazj291OMDa1QGXrClS9hV82RULuuuYHoXbq+KtfDWQPwj2PW
qf/ObzQ45iUq6WwIxNQENFwLVYyC6Nsk76yu4yNHDpxvaSYD+sj2LHK4btA0
F32fVxLc279M2SuRYVKsotD52AX6YzIhbVfNqZaNtPbrmvrz2JqLFJgmVQ/T
mTyGYAseNMGpdjsXVvKADYYXjhC/NweWT6co5GSGWLrv6zSH44FphiMPa6ED
GU4586tE6yfsfoT058Zs7McQFHXd6t6mgnee6eMJkDcp0WpGLEP/a11P0VFN
ORXG5EhMORneHTZ272EPA8Ir42OYUdlxG5JxFoefBy9WCl0JsMmN9BFURVkz
ENrZ4muyyXP0vygQ4siadPMVT5dvfdl50sDIJsIag0Sw2R9J8f2iRTi661Q4
1vdy+2Ut4Dg+7hj+5XTa62Hcs0kyVjy0S7TFykYXMOo9VitA9VOgJ0CWJjs5
oMKKzZR4CAz3SByI0OOIDwHkII3vMb6ybQB00+4p4PS4TkB+hFP6VWFTwHVN
7un5QfADe8i/AuElh9azP1hnd5hOWDLQG9z+DG8w8sxzcNnZlAp3e0w+E9mn
ffnDL8I2wLoSQicTnCTRN5XGfDTS6mEpT03g5pJEBRbbukpLfSj6/r84kN+J
QxbxEgFAgih11bv733HW35uH/DrvyPtmuuyplrPwvsohOeSsnmmMmV1ZCG1S
vJHWXw1qOjfkisjN7GX54kJxUVeQUhqITW9tRy7Y8A354eVfzKngQ9IMiTES
N6HY1Usp1/KKTZcs8m0jzJkv8upZAIo4svKZJV/9xoYDU9/1oACZVUQVPe8g
CQqwKFL6uhObVmLcIUDs8yGik1BzkFfWxJeSvGI2X37ttcJsRIiw+oo0jawT
ZXXnTKFoFKhqTDHHAQIj4ZHOndnjkC8pyLtWpYDer6Vjw8rIggD0fx9P2Xzk
COS+6YuBGNdeFtvUsE3j3k/zX3NtxxGT72YXl61EX5g+7inP362iMzNKgrFv
7e4xL4oBI6Iat8Lsf1LUxaqpY5Q5nETWULKwTJCEUyczWCOdOrrR1LgommUL
4qzv8cRUoASoWS9oR/Um3GwKdcGGf0Jb2hAtmcgXhVlS3FCLor5t/LBydy2t
cWWY75eiT3zzVg84Y3RA+igxJ2cTBOZ1ct7QpprfW4W3xw9+UbqnX5kyjLmJ
nbnCeObRmo9haqIuE/vBwBdd01sGGVyuDrSxJeE1IClQd0aFYHtcSOcvXwqd
7O8utbHNIL5ybPJodJbO/mtTrVr+pkzwKtmMocKaLYs4C/hrlM2DB3/MAZpQ
LnbPfLaWyfofJHed5IfSM1TFwsc5WN5q42sLFbnsRWAzZWA2pWRCNo+JTTit
GiRPz5ivW8KjUoPrpJ3zuu/ZaxYO5P30slfodSW9BIXg9iJyd2fla+yduIEv
t0WhwEEleoFAORbOllPUzH8+pUrHGI4EAjmsNPssK9djpbJCBipl+bWpFl6M
k+DpzGp5bpsIsaSWFsf/7CAyMQ9qGZmYzfLkF1ceKq+i1OA9eDl19DOoStfH
jUSepPV25KkGcmaP1sUjoYyT3Dbuni2bwRkHd6aQPi5F/cRTC5wDIG65UIQb
axvGoznxiN6QmOLBrCPAUMmnp7LlA+ZzIYge9SQojdRvTA2g79GguxC1gRp3
WY2gc5C2Fue26Wvk/vttqZCyyC6zCMv16hehNyeA5dMKufOisQbe948ch8lK
wDYnq+VuJ1ZbYLmepmVFrj78Z1MyZXfOtNNpIhTWF5sgvex3VlhBjI9szpLf
QAAVEGWSZxWY0cZxUPawPPuOE11oQp+Fx3YILChijWJMR86RHgyOYkPeSiN3
7ArVSw+qH8bWBkSb48hoZzndLdsPPI2vYaDxAI5AZ5iHewBwU0/s0pLXvVWh
kDvqfebUrqFJC4A/MyvPBUKffel73lujja6ZOKEnfgQMvnIAAy8V5RJvM1UP
Dd0WsvMjXQMwkJ/pjnOJsHg7mkEmYt/5bd6Nr14mA9848R0Pq1KBqL1fjhXw
4eSyc5FWhObaL99L0uvUGdV9mGdVxOLcSS6sfaeLk5m9qcoGRCk3UIRXkegy
XRkbDMCnvSeM9a1oDeq3/RmRELc4S33SEROs6bKNDfqTi0nmJ4zJteQ84aTX
PNXMFMIoi3l6VJCbMEHDRmc2u3kLSl2/qmepihb/VtaqgvVHbMRiPGlBhGa5
GXF+GvSuIaNor/B6SKd2v/ALQ2zoQ3TfpKx0A53TJWdUYc0iB5RNXzWpTOp/
7+4GCAZ2twdZtnx7I1SSFshEeT+fVwWuASXuaxjbuli9TbiYE6toQI/adnTV
xP45EdiRcniIj4wKWS7VVY6XYcLvwFZfcQ+9QSKrQuaK07qLoZCbr6kt123C
nq/qgIn/OeYGhpPBGhB5bDK85D5YVZIfVWX0en6IJx0EhieAkSkesO0YytBz
n9EZttKcTEbDhkuv1p3fH2UBVcqeKoRigExK2oMtooCzGil2r5nXXtFnUrRp
USJYgZ0N3izIfwtTTk6E7NjDTroMr3y/QNFgWU1Ro2ogjZT+AG0A5O2/wL/y
OU4XbOs/je3TGDPxPPSpjY7rfv/s+0FolE0QNRXC6bdJxhbuTmRzNnWq+Ca+
d3Dq+DK+b7soqHMaBDyqC1Xy+snlGThbZYfY7ncgstD2lxb5hyTIj1LNEpEh
VX1TG1Ih0fSAU84sJoOSmXsEW+iThwtXo+q/V7l9WGlOiU3rkQgIBbV46Bhs
XAe+h2Lh3+7kKjPtzzOFAYbnmlcN+kAG+hO2L1aXW4sjL27mgs6HaXEGuem+
rgXX+MY4/h3aS9o0+6CWpDMo52MP84sYlWEguxg5etXDF97iLefm2gFDytHi
oh/BsOrz5wY8T9xkW+snAYjfOvgf92ifDfJ2S3hZe7tSLgLBnTFOTGSMpm0R
OArWe8pJNTYYWmtwlBRx8qIY5pOMbDZYhEmpeVAkOuXqXlPWL7kT/VVezrnl
C5WccFj3khJpDnn/dcg4MWGbALhmbkoJztvPzYDFmM1TMankyvVWvJ732Uct
Kt/GuHu3+dy7wGMPUl1OUjwzCQUZf7uYx15JLnu+tYbM30zTqACVxXlF4+qT
MvEc7wzE5PmX29BGfD01Pjg/8MSPg2gA2lN+RehNCwMXD7aPfFM9fWPFbayM
8vULIKURatNQ+GEwtfEiYr68hsITFxXcrKJ95GuEJr/Df8NGWXm3Q++WyAGr
HUj/84FjY04jv4Ttntp9MlOgU+3z46Ug9yOIAKdGRLDs9WKII3SJp2siPISZ
QNIH+KAMUld6/gP5fU68sgs7nXx3KKPZQjIgQXi/m32MXoatVk68tTPMcp5G
gbL0Y8abksfdwZRt0etj6X3MvHnRzR46fR5Gr3JaVVchaxdk6BVkhjOypjYc
CU6zlzahtgt91MCGV7faMf8JBvFA5ZNWdsUXAL7p3Xstk3AWxYo8HNy8R8kR
YF5H1B7Au9eNfSuOnvzuyZ7SGrGFp3DBhd1JtqmOrwcwOB4v4jOErtfalh25
xBGbRHTO+j11JF3wyPxVQZQ0C2neC1ZfVLIE+rO52Hcb+5B0ljlQN6uRWFLw
ggbC5ZQz2t+I86/NB9sA55CkQEfTK++R6Ykgy2SZ6CFpDl1HD132ykj2G6pd
0mLCgFlLwEZqIwmpkHIo/vF6UZgRHcUR1HSuXgC4cwXj0aFrBVfio9j/0k5j
soV4P2puD0MX4S8Hq7DCxfsCum6V1E6XgB0EaNS7SNrDG2lwA7ULsH3XjsHv
WZhDqZj79vHpWgocvbUE+mh4dXQeo7yvb+6XYb5K7NpneI7UX0u2sWZsvGNT
uYKbBFKASdonlkeYSd5eEsjPd+yntaknTzV73Wmk3woun1ztUNueCD85xVs8
3bG1RvjdtC5OG+B3PiWtnXN5HC1I6hFJX/dXndhsVovnAxGrzVHOPnbGYrIm
cVpDdG6mQi6Pr5l8vLO4QPnw7Qwf83c/AE39OswPP2Wm8/sx0ubPHtLjOXs0
CU142Z2otUDQcg5d3uo1j+/xEgZkA8OBXyK1VscXAru8K2pZNOZq5g9yVEiM
OPmaO9u5GThIK0s1bRmdYOLELmXNq6o3A5jhGO475lxfdTEn1DZ1A2nlOXq0
0SEap++sQtOVNVuoch77UrTKgXepND1c0y1iLA00wtVXpSlxGSCByxgGYs9U
L8jNxI/QxTiPZT+o44uOGLD+x63A1jlZZC7/IkqIx8I9fvzoWcpiAl4GW0WG
/4DLUMuu02cmHXYZicpxGgbJPMVuNGSmgv4myjKwNpHXw72Xd5YP0OYoYd3I
2MIp89pVptkNXeJUgWcUGFB4TVHqP/9Ydwj8m+l6sR2nz9+yP52SXA217kyF
0jOk4ubs2Dp3ksamO4IXtJsoZCM+n2ukLzqrfQOug9E9C4Lj8GH0iN0qgHqc
3scocnHt3BXoxzljC86KDgA24u4cks6Ic5Ltc2AQdtFDq0JdWD/c2iPd6kxv
rwiZkBkwDlcLe60H0guvLqtucW6ghQmOilzXOu1iXobvIO0FhCaP4Ogh3BOx
+qyMMa4hENVzd01ATXK/PY3PpKv6H3Wccz+LAaIO9vlFjuR730rZxGStpDtG
jcuw2xWC60VijkjskuiZK7/VIOtUs5b58/RCHFTMGzJamJIloEKuaDpEcFdy
iOtNllOgIImBBEjZGJkRHDMcAj7qQ5JyIrsxUeYw0MuRHep6ybQXAqyNTKoC
laUqIzjpDa8aSt2TQhoTE5QRjiEvPPWf/4JWyKCGtHVhcbXjYCoE9eMA68Se
EJ9ghagD8KTXUj8QtUQIrvBb/sRV+bOuYdwGX86sQIwDgXz7rtTu++Xlq7Gq
Cr1yxK8TX6GEUVCqdhGrRp5WXhV2cenEC4YyKU4r7LhAxnU7G4o8DtBZZTjq
gukfWJpzyCnF+Q8QqWFEuGUBYKq/nzJgMU+N8m794CPrah3MeATj1V+QgAK3
FThFbcoNGDfNcGJxDQV0oZVFoIh0K9g9uK7jym5qdwwHGUN7tQioU/V8/vZg
57ISDy5pDSwAquDFevvBkY9OFJImY4G0FXpwprOKUfkkLzuaHxt5sQ3yBLYy
aUDaAsYLx+qb74c7dMoJq7zwkV54T5gCiMVHp0S/ytPaSAg0fkVARTO8njvM
MfYlCdh2Q8ybvmCRtJFVHgvHIC0p+YzKONHADwWxbOwC20dnuzFFdZ2w9+O8
9zayiVcs8fht1ljN0bL9tUbJT/seYYHayT3m1z578ih7A76bpn5G2892dByL
cQ9bRN/dQ//L8igM0wdBXC9z6iaZA7ywWaOx1RpPPr/xXiReNBPHfQazI+gO
vVN4wC4SBD9PuCxsrc84pTj7DRQs+ezU58wUqNpfz3w3kqryNs7gPcCZmVjP
NTE2KjoYo1JwOD3rwWw9coBPvc3dzQnErDtJSVtdLKhQdcpIlN4HbfBIELSk
5S57egm/EDc+Ji+p9WdPU0tpOwckVF/jSmIQKH9dbu5eYkydEDgBoe9vdUrS
coD/58Gg3+VGcWqTKiAoMa4lxUQ/8RMCMU2tUkxw4FR2e8Bml9ecvw+Y/T8e
0rffy/aDiQHnk8BhlxieU4Jw1JOecFyAa9yQ5SwtGQ7CvjKaO/t0qPSSwBg7
ZJgVvLERpXvP3b/GnsBmZA0MlGlyKzNholKjHEyj3z3Lab9NyAh8bCU4AN0h
g3sMBOBWooG7tWT99ap52LAsrpVTYmmB1xl22IsQjjuKsaMg4zb5VQ5vVei8
nicqomMB4duEcna4jLG9EGumYH2eK0Qbw+LwbafiCk/1buhbQSqZsiAAt6H5
8ootck3IpE2nJ+edpkDi0ey2zhBsIQEqdjmFOKfG3oGIdtEm6mVFwCgR8mmk
0YZDYIRgo4PmkAGLMrfRvH9b2fbrLpZTGyx/MbsvHyvBtlUlL0lQ+V52NF45
G5PdmCdqAUxJt00sKwVyKZPTM0sh7J/cj0O9mY9EA1SpgPER1Af/O+xhoDbZ
vVnOt3R8GHoTn7xXpe0H7choWmOtmOUZ44rJn8xPmraOXuU4npFcY9KUDcth
VQq63G6MD6H1GCQVhmFwAWclzBCy3I8XMxAHs9PyU6h3rHKEnnUClAg18OG6
73JIijzYIZkeRGYxuYyi+8oB1EpGDeatle601DwXs1hQ3etqHXnX+xxMGidW
fPKChMeO051SUHefXm3Mp3cWQNv+xGJXlI4/sD17apGF0/txs4IZGBi4k2XE
uhRFiwhoFWIGlgEVyZswuRlZBKqBKbHGBO/fMl/PDqfzlWQ1lZvAQx0a20Z4
VNu5LCv8vIZ5r2DWB2mP23EAsKNy0b6j41rBt0rsgP/WEIYQeQEUjoO/Jdbi
8qDlyeGtVakBt+S4QctUjVjCAy05/KUQujUXnQUYFBTuiIUNnvJtZCSvqbH5
UmNt7H+26T7msbkplpQRxAYZClPuWSbfSYN+2mU5zuNiwd2xOPo/TD3tFByd
tddB5c/RlNVHx3vhTX6M7V/9uGYZF50uEVpGkBmMhAnBevzKl5eozwFuyZpC
b7EieIQZm6DB8wkW0YAQbkMSYpI+oo+5dPAB8IhSJRAzhqIOwITtmUSBuhnx
X3uhS9d9i34o8/1DF0kJp8rNItN6uzKXD9pkflNKmJF2+a2DzJyW7uQWrWLC
lYMrqJf3UDERPNAcvlKtTAs0uFpfsJI9XwGtIxLtuWBzZrZt3a5wdHrDex8F
gH91pwAvbAtr4FENh3UgdlyfPwzghIDtIYrAMDBV7FBuq9iTxmmzb8AaWoyf
MUKe927W10JWtF3t4WbYSO4ZLV8xrQYXf+ZMBZ3IJZByAlS6fLKSNP7JWcqp
VSN0cv/k9F5diSTKeocmomWORMFQHCGsIl0cnP7iJ249iYUzXGjHZG3HB4DN
9lwHVG0ycBfwIcKTioCWKhV4Y4bC0tv6iKw4nxAlIYsyl1D2WgBpllNX+qi9
O+PFzcaxcazZEE+GwJvkCo6D2OHUN3FFdfcbJfazwZo85qFdy4Jpc7s1Gtdl
3kM23wnTNU1Hcoqo8GNR/psFfJmyl7S4iVi/qnoUjkEKwuLrbk0FAMSey8B3
2fNC0Lt5P0miQg0fV+RP53zZFmeqH1qYIeU0hfSnTpjg5rFK/iqYMgAKDKqw
Sgk/gQj9FikzQ5dgJosvRaIJYRGprNGmrmFWs6iDMe8o8OMHfH9Tjh3LIAXu
5NQWR76lg75yEOob5gxds03Ak43h6BOAk4lD/N45AnTROhAuR9tTAGnLCzYb
tQSgZIdaf+jLx0xmNWG3Zmdu5IcBAYSz+pbP44+dUhBlqlBP8v3XUMCQNhmT
hv9S6mitGmChBJuZLyk1iSVYTl7iWHT+ZVU8M7emcdRdJeID7Hggof6oUe8x
cTyiPCLE6Gjn1UUcI9QBFZvBVm6oBdP8d99aJXiQY4UWHjvlnvIbx8+ZtG0C
UHgIfpcxI+1kERo0ncZ2AioQdMgTCXI8nSkbWRGlO/6TtjzISj3OqfCJey7Z
2x09fAYhkKYyIk4PwzBnUvOcHbl0ERiMtIUQRWG5f3G/K8C8aUnAoBGXezen
qE8w8UtuL09WQTCBiYGL6RnijjugFx1D6AnbtOONGeOf5hTq9RFJqfyWoxui
HC6IK+l3TXOxHXMTnQE735JAv28JDucp5Qchj5k7Bkq27MI0L+7snCB/QXn3
AaRc30Dll53E0jdh1MHKiovGItybBEZjQaFqkTgbJYyscQkdmda3Qv+m/wD0
kc01emQn7LV/u1tfGl4sHso7KTj1pCuKMEZSUANFwjde4bcWyCBXr+9qvCTf
xLhGaOBrYfCqwlkqGB9r1LLNBFwd2mD3wp36kQQ+VuQ/s17bYTs8JIs3rYKY
i2QBbbWeNUWR5zD/pNIKQInfXSIUCYlDHJeCQV1WyhBGZ3Qy8RBHNZfGrT8g
obF+nmBRpL1DBs7CN6FV/JHBPjvbRrzmJTHFAaL9vN8JQbROqCHEgZEuEIdM
AgFqWWsD+AYSKa5Mdk+mJEkOyI36uXN/Fs9naeOAgqCU74GkfO+P7PNJsFVr
57sp2FqJcVSvb9B+ec9i2Ku2EhgkhwmrIatjrtCnzUHPflDkMK9bT1LLD4Si
Ct37pJq6mrL9SgTGczfxj/fjwaazVCXhwixhPfazxVtNVKu+sc13ubaMZmTP
KJspxdhennRFiSEI6CV2UKjiA+UXDpL0Yzx8EbnMQ2JC/IPUY+KWpI4IxPwh
XO0c44XSHOBI1RT96pmQk3tgV0UuhIR0qipE74d61ZUXsi1KTUELeMuh68/q
O4oYlqYVG1DqcGy1pjpVIjJlWCgjKgGekyPbOzUM3xkqSnM2miPnO0JvNl9e
JhGRRA1EUR504Ofb1LwyCCUucA011meOYZUnzk2SeO3Eo1zOUikI0XXqNyYT
zVJElmof/98FS6ecvzhjrNFPCJ91Y+/juWH06XYdXkO5erS5eFo5HwobaHFW
2PLoB607hLI5VTn1JNv917W0ITyysBtd63V79SiG4b6dzbJXap5/zbb7jrbK
jBI6BdUAtqflBOWIpOJ2RC9Y0AYNX77t9/9TxLCvlsElHBRd8LFjpkwYmsiY
tBOJVjaE/rTXMZsu41nGigSgAr5ynJyt0SuxvmlhjECCXFTVC7260Gxvcubs
yJMArnyk1DK2emMzMQ7zYywfyxQK/2LwVPpC+HBQlXfW5I1mVfNex3enjbdU
RQf/5HqV8UhQQE9sKBxwE5SWBBI9HPLZqcNNTJGwOulrkk6xv8/x4IfATLmB
GdyQIQq5kHCnUjJ3Wru+BCtGv95f6puGyNuV3uNr0olWSLT1QDamO9IhTi4w
/XQG1MsZffNvohhToGxkIzKpdTAqtZv5QIpPPb3xS5WuX/mMed4gCjjcuUuo
ElpJW3i1lKfGFoY6egMYFjRzZtHyyJpPi6psZJSyRz/BQUpT2L3ucu+xevaP
N+mjpVV6K2OO3qJdifD69K92awJSCnkmO7y73soDqVmhSd8IgjVwUw1QYjRH
tTKo1sN0espfukZeViw4LmPKEmo3uxcaq4/NRrq+VeXsk9xQ1y79mXIKZ2um
RkcZnh4qjahn+Mnd8lR/EWyZLtc6/tdLwQlj4IdOvYxCgheXMdLKsLsxBq5G
Ac88RRNM+Cwl3PIDgp1V3pAb4xavaPylE8lEHXxKCKlyUIou9D+WchYU2laq
xXeuK+oHTXsBMvkiqWbMqxeeWHmAQ1dkYs/jmHnW3dNKf6guZ9nR4JLgqqKa
nysd+YqA3IeG0lK+oCNoMW7zGxnYHh15Brc1FNA1FmVdN6o5Vk75ssb0NcHv
kDH18LOwYrT4QYtLe7dpVnD6RLYVYq3Q0StZ4ZjVwy/OF4P0lITaxE3lRV0H
3kEvfOUbVOGICSC8OVAxXgn/sP3r2uROhYNlSDnl8eeMbP6ciYdzmjCfxmuP
t/iYqdRMUFEyDoaydrYKJYFFSra/aUVb9a852yDIxRnvYUSCQBXQNErzK/dC
pwClvAAnvktv4LoJoPxKTEG0cOmNdHJbK2C9J4as4i8Ybcgv4yAMA7KGeDfc
wHc7ACmgRZbYp8Tcox+ldz/9mcA7dAbJNKN6D+FgctwD+NAM+ilMgGKFcT78
A9warFkrmMJ+MwKSpuChyWjYzSK3b+Ugr6l6UhmAYjI0v4PK1Pfe/FfTDRV6
ElkV/GKk6Yu/Mv+CRltOcgRMtLNA4ABcEf2Uhy2YAxwdV8edKItWWR8CQFYE
6ngRPPVzoJzXSQ3f7eO5/nHe4p5h7SrxG/hzni+DE+hUqs5lkbJadykHrb4d
LoyUtm46uWkjzR5OLaL9XCCCLjSD4HG0LBYJe0UYKiTT9R17Eea8s0k1Gj6Z
CzQJTob0mTUB+vbkESSG84ghNo7mQBbp1YoTQwuXXHZ+5FkLj2s3x8Ingu+B
8iYDB8XuK9nPo90HDi2+RUuEBs8Hyd6SAS9uLeydp4x0vDqiB2itEAjSX4Bs
5pmDDHW8Gkq9jPaPkAFE1+Bo26EvgApfgBok+BJM8rJeVp2UWIUgImDxGVWM
zrnWmjxzVp0DxnDj4H9VotwP2AfOBMTYtwGpZgiCvn9Rji3ZQgjD3Qq8PQBs
9R+puOVU8/f57wxKvRi4/BySBaOrsjU1s+WD6IWXBkcXzXTyEDOhrEa60iII
7rcnNpOX/Sg/My4mOUaiaux6Zg+df70Ms0R9V0BIzGxU2G+3jLDMDZoPWQI5
2QjfhAVz9rAEurr3eigPVlPFUtPbOyg9stJbd4qiVy1cSHr4OrfXUQyDx6LQ
u2mVT25PdaJf6fo44gG+m/TYM9/f6qzbITYaCqdJ7MVPlfdoZhm0/dqIvpYw
KIMyeQKlsWUla887tkjG1YEzHIBMD03A90QhoJV/Qo8I1/QaLgkS8mtWHFLg
6gqSzvFVlvi6CBT9U40vHrFQK497ZIMT9yJTNEpYihU9+8QT4e3rdl2hD+rN
F2Ls78hIJWZ1uE8MkSDG45G3thcZP/mAo0YKq9xJu+Gko/ktijrd4RItZCOU
r1WidzWMTWgRfrDd073LtBZOLr9L7lXgj5IZu3TtHN8Cuv+N0PqnJhoUVZLx
Lub16+G1N1pRJr++HxJJTSqFB/gt/E+CrJdEXvQTiDpHILIX5oKvudVkBKcp
bN/Jajyqj7xVlWDTTHHe8QFVbcJymPGDQAwpjfzVXU8IKN43l2eIoxex7UyC
QPmcI8MndL/imPBl4tfOnlmNyKxRyoFBnTwwiFQoeelc4eLTGhEWQg39Efbb
oIXSqsZbsknBG7HVM/7JNyRIPOaSfLxTh3XoLf5DDBzGeHKxBQHktbs220X2
Wc/nxe2aVhx2LyJRdKoabh00DovqpoEdoa2oAnxomr3rGfcPI5R/JLCtIJu0
gA6c/cI0wtPmLGjZlpPpewXg12N+w93NDSYEE6KbBg+967E5/Cbb5UT1T+EM
iBvE+dWiwsuCMsrlf9RB5h6sVMyiLgfsCCyyj+byou7EabJiJYCztVWig2WQ
ctnpR06HcQiC1PVuKojBhfZuBQZz+rrANRQpbfTsFQ4Oe8v8o5T7sOhjB4uT
TLSyjbYMSj/+8IK0/e4XscZVX+ji2/tdQ2VFr1cSVbsJyskiRFMD2i+5qaVy
2XcHnpobIkViWO4Lj1tUsufIylZs7ap+895OOM0lGYIaokXPWzWscm55rzE6
lK6BK1bEJnxkA+K7cbgIRciCT8/Gba/nmIwL5CFC8egmcCOpqiFJwjGMcH2g
kWRjURkKb9eDINXGK1apzEFvFX4FCrbw+OkupzVj97JY+w7tMVh1eraIkkgh
+XzrWwUayzBACv5in+ioouImum45rYM5ricdamUvziTy8UWzRiYDTvFy4htu
csW/sIK9xEDeiG/ECZNkA0LhwQAOi0FHsII9tY9jTiA6O/tWWcpqdwbC7iNE
LvArdR6EaGk56WPHrB3aogOgXuT6OxUAIt9N1lLxynv01Qrpap2gv+Vt7Nxb
jxMFDJ3Ms/P3VBNdQUJqagO2OOc4qlZ8Z2vQfSSiM9YrG9Zs5iN03xxCKwHJ
kMhoowOYUcSwkRDfZWegaEZVvZgCXMD2kQhW5TN+bVZAmjZ2EsbfuOsuEQHh
H5BjHrcMnitmJqPsn49mdsllDSk/2cUCM+oOGqVSYp7NWvOAd5p0rtPhlXNB
yQgmkR3NiWUSYnwpDmuiwtAWNMvicRTQSJYm7iDZ2HAGz18PLiy41TiG5uSV
eJKXkBhMdnscWVRQagmK3M3g0VC0M15nIg0sDkpsmkBx3S6FrdHrPvvcfa0L
FfrsgBvaOtp3XLIoj1qGTqyJdDRPR6MAPuPDWFKe/2aes4rIIbxwxerncte5
l14ApkI2zJjrnYS5bSxUyzIJ0p+QxEvmzY1zlkGsqUryOJzePuvTyCq+9vuT
2Flzj0GOVtpJuoDQDt9blqCFpe3+/1cf7jWFiy6L7jPAP5pP9nRwNoyaUH/v
Cjyb0LNMzpVDD47jo1UKbwF8ipACUec+MLRi5DBCP77AGthCA9fjfEuEul8Y
5PGtgxmpZwdJcG5NLOlyAsMh3JLbNTbPdSui4TenD8DrPwiKjv8F9NAV5DOB
W2PL1FR26YFniMJ0IY/PzL0rFwEmTqRuXNLYHK6bL20ZtHCD9x75Tqq0gqXn
wqsKTlLgkDtSaYdAvmgo2nHUnGdFbaQHrwK7mJELxeowurqTW25E5INunn2H
fq7hp9dogGVYfR/OyT50xCMk3nMb8UGPbmiLV/MjG8PG/FWwxMXv5fgc1mjo
k8HdEmadrnRwGZ7zFW8Tpn3rTgq+lugvoKdr8Ao2dU+w+wo9AGpbEWN0qqQT
pHEt+Xl5TTwIFll1lNySPm039ngh2HojZqy15D5BQ/tvqQ7nvTBjzTv4u6PS
60SPupNudPuDO3x34uwx/kHJ2VW0ASpq4EnrMGX16HFi9xLdHSqPIh7scCzQ
fryZgi6Oai7qWPy3K11NhbKykiEoyIb6gRrRwtEH2xk/yLokG3h69kCQj0mt
8X6oTrSUIZf74exLeB+AqFHVYkY/RZBg680gWZUY3c35sHKmHUFkay7tjP4D
YVLuiON6LFKnObZ2tYa3zD/+Bz6ajN65g+TVfOvOtT6oFAbj9yMGru4Ekihp
0zKNQFdYYTYoCAcSY5CUWNrHIZCbPrJiENKE+RYqtzv5FZ5b6Nzg9QGH2Iop
n90+FaxRj08EbxPlSNdNEGauxBm2lVpAvAOTfbOjbKKHvugH5CPcDt8A6QQq
DDUhRvRCk0GW/+Bv9XotDSriioH90+uSJhi8kF2xJyOA/7zA2KteAOc5AMO3
aGtcy4/XqZKcUt4Nbk621qMzPEMxEjNCyBRWPbZw54LGW3QXjD8QdUDzZGNb
C8fQIWkovpWoeTCvc4VQgAjTV3r9wBZKJI0e3mN9EqfWT4K4yoYQruSFdjI5
DKBa9yQJhl0HLL2ybAiHca/kzqcEvCUuf9592YUNNlK8YEtwSOUdb7bnJR5m
HstYPMkHFyHle6AI3CuFoCdr9avtUVOn8Nz0p8DsO2JcOyXc6vilTUVhavBc
FfXddBynfSf2Q9NcNhBrdzmKWdRlDyEN2L7o2uR7mNl0OxcP8S01ikhU+P4s
rzXp1m4/sh8ZxX4bwG6KSgMcHUudqwBHKSknXJfz7+M0INI6URF4kBjxI6hZ
9KLquYCtB75+QzHg859ArzoSKPfe0pYO5p8OvCewo6Ef8afC5WsYblfTIVMg
mKbP68yreuj//1JIy+ITI3ro0d4PbbMK/X9VXfSNU2oeu/M+9hN5UPB+nk/I
pTeuH1Y8khQf6rf0lBS7AiP7VDbh+Mj7AVPQ6xJYDaarhY6ol/Z1v9/cYP2b
rQW6CpGp1yhjG9mjfqFYAu5gV02waS2/Z6et7zlwNrsC0k3M0pl78famICCu
3mGgXwR7gkwkz9Zel+Y380WLsmqNvBFdrKXsVrVDRb0+XdEJV9J05wT6qnO0
FQQZYzoPDe955QP5QZjAqO76j9Hv1EgrBi9VgL09y0tsA++asC17V5AV0q6v
OBLs9p8HC50g3kQRqvRZjB4DlvulBmBf1wtT4xIcUZwQWm/9/GN6e+IfnXwD
jRNdJaWGBp4W0EzXzXkihuuGhP1GE/p3uMTYfLGSQuNl3b8jvQm8uQ945ECW
t6zwBslZyONFdKgeENAdQWS0Fb54MZQXQLzGMryCbbFaU3Z7n1zN3aC+CVyY
MCAd5F1y3Q0nAWrCU3J3M0yk8PKPfnw/LqXb4bNUijpx+j0q9AOwxd7gpbpI
2XS9lILa5BWli4RYrMas3r6oft2zTY7FKO+hk9lmKGKFq5ZoVAlJBhoqBgb4
Wn5/vjii9v4tJ+uc6AKOA5XEVlb/mh/STLNVKgGFKWqhcaWNRJqJC6HxoNsW
G/uxBKDSMh5im0usTBbAero5ZnFSjiwblqjRqz8w+lr5FKu1LFaqWa//fclK
zYMb66OUC1EXKnSQDdXTidLGdOB2b5+dgna2At+qeSrhy2PHs2D11eDiaUov
uLblxkegEiKTtqKZn3gMxH+iE15RBM/vycAtP/7G0yvUYn2sNcfb3swHQMAG
afhErAzradRnLih0t1sR3sFRkC2zJmL5OwRTRoGTgI57fJcfqGYEwTV5x1h8
hfCTTP7FZKJPV48oHv76ql78vR1/J8YmEPobhlbIwnjkTxTNoaEXdjVm4+gD
eGDNqkVaGMd8+5ZOGRPRK2cYAYYUHtjwhh7qMCeglWgzKB+Tjv2Lzq/swGcR
O+gR0qpcVCx2Xqnefnt8/i5OW9jyn1umwzhBtBRriZ55PW4RyX4bctFh3USY
gdRg3C64lg8jSE/yOQj18FaUY+fm1bjfR9WU6WGn6sbUhYphrAr8slAUQEx7
xKF22jRUlRUSyP+0e1aFLJXVpqXEOJuITD9q7MUKQSy2M/hL3AZCGHFCNvCh
ZTXcWa/l9/0sdOysCw4yatwxa5igU5PpYDG3xsic+12XSuowfLXkKHLLYB7R
HRYTM+4TipLrRLV2B9u7jkpIkrAmFNAu5yXn5xZHQO+N/3GEwVJtHWeqxWkT
JcNT1iScYxNVwtk64Cw8SGKZ+3do8AzPy0YdHmnXuQjsQlU8w85JhC8JWmUk
HPw2mpikZtjQxacNSl3MT2XV1wUCcmDx25Cpe0iOpPaAzSt38N+ES5USjFyB
f3coZsQPbPFFuy8Ku1uUDJZs/boG0hWdyeryo7LYonlYJ7QQSl/sN27qKJVZ
4U8Aiap8WZbV2tPWHuiV9caKSqfCALjuDwLRRWUVaPHf0JnnMFPaOm7s/vum
0zv1m5qHPPgZukAY1hqT41Qcl/FItoBSM/pljiUYST5IpwZ9epunyTiZS8LZ
r2ayA7pnX8e6LA/VdKKw7B/M89BKchCejMZi4UCopjqbx4XYuCglawLF/QOP
GkK00kpVWdITZrivorb7uodJ1lOWXe9qctocXUm2Do3kI9pFZzDNJ8tBMMES
CjTL1ruuSrqMHmCXDSQYYECrqkXLR04laPGWpRE3tV6/Lpv123YNYb0XR9/I
yies9nXkEHlfF1/hsUvSgkJcY6YEY/SdrHcVsCvlCA4KihkHxQcAlMHQheV9
JNbKHbwnfBIQ6FCusEDI2REKWgguKBD6wq58SaYS9c4M6SjG0kQ+E8BnhbHf
4I5hGI2nOm88QVSjsinOL62KhfsAy569yiCd51o3tUrJXuFcly7xxMyRZJ3I
8Jg/mfdB1FYrlWzo681F/ZfTdHGXSv+9DRNciECXiWcRPaGsor4nw6vhq9DG
3NMWYoG+8ba0NRcqq7tqNu4lJyjselc8SuQCF2mjJ67JDTirt2DrYHd7bWKe
2/4eGrD6JgXXOoaIAwi6D8oFS5RT/TgBO1tpJORcCSahm7b3cjOgN5qiSN2n
taLcKjFwLXFHDHkt8QilzXE1vNSXaITq+Iyhpx+N6eb/gjQRo8TCmASere4c
Po4xflM02Fn43u0B7u+jXl1XRciXj1msf3iVwgrKweEYl2YlI/FfDNXmQAXO
h+x73gvQ0gWIf8M9nac9aYszmipiaVDDdqq71RDcTpRIY3SZb4Fu0cGjL2ZO
oVeHYcPXGWVTU1RR/mOa+mdr77btiyYDauLBPjPL9a8ZFh89VhD9gom35dbe
EGUtKjk7OTENv9kC9MjdYgw8+C/tnblDqjRGglhzsABi+AvDKO6ddKsm0TLu
SkAjx8D1/fjIDJ/RUH49D8VK7yD7TxvRgforkkcNgPs/TqcpJZEwhwU7BdL0
pZ+Qa2g1A700m8ckAefUPOblO28/kYUE5DUrwVkU3+okfcTZG0/jNSNRXO6h
03+8C2cEh82mASC/GrlWKTeLXMYu2neGSNA5GZOvetUYZ736pu9NAVY2CnIp
t3i9qyBY7qjYUH4kA1IlVw/BboxSXWsjBHukSSqheq5WWWnSIrT+mESUEDO6
H1BAC1afeTNCXeLUh62iT7nwRT5yhiZRUFm3FOif/3qyA2Y4/dxqfj6aEs1b
wkab5doXmRmFakU4cB2x/JgpQWxw4rAeHSBSYdLDZIEar6VudYlyROrWzgUb
Dks4TbDiYLzOSg0AWs42v5D89RNop0cvk1YyWgpitkQQhb61BDlrrmmwPUTQ
5+5H3i9uolqwfAxH4jBTYI9qJH7se/ZkHE/zkotjJRjcC9Ro4/Nq7gIi52Yi
JjE5Pfaa93cCFv1EsUXbELwkfvCgMdEBGI9UjfXRwKfXVaxK71Mn7lR7FwGi
2iY/OHPsCWwOQ1z+YQowqz6+fdE2MDw2siy7MS7PpvYDE+0YBWaRsVHb7oU5
08/NNNssKkXK/Fk2P+mhDipfe961BebgQ1VZU9XC8fW2LZBGD4btxojT4VkY
cYg5mRQ1HUTfR7WroQGyosVbTkwQFbyuw7W/ISkfWzbsbpizLiFvUrvSFvEi
yMHm9eZ6l0+pQ2wcTDkuxNlA29759p+L1iDD1Gw4+6xCgZIN1f75teRPA8jO
endikemYX3mh4U8BkR5/xtAYxrH+Q9PTfAZbi6kLFkZXto2ibwHZcY96oCoB
4NyBH5xoFsanb5WhKv0ahi0xMMA8iIyNu+rhFooVliuT8gxLXbR8ZkY+qUx4
TOJCwNh0tKS5nNUHGXkhhE3FfA+RO0G6bile6Oknm149OLKAHzhscaPIoj7L
uirCClRpLr50OEfMn+CJcBkDeX61d32fIU1yGrR5jKmhbJwB68O1va04hyP9
EIjw0CjRcUXA6oNRd5nxclE1t8Y9m7fy9cV9pabRhkBR4Jklehx5V6c8XnsH
5xy2I4wwsftm7uGzES86r2D8uB9iYs9X+TXA7cAjP1X/YOSNXTyFqPU4+4+2
KKgF75ANn/NfqABKPWarto9+rZDxqQtcM6sPGzsyHMEnKcGjvt+DfjymsHmp
JA2qU9T7cux00uyIZ5aIy1BCNvcgnkq+3aaWKhLj9KZfAQ4928cpxYK6vdH0
1PqBizZHDgj9WSXH/JMwN0ZnXcrNAcQJ0HoXEpMRpAz2Zce0YTYTCoH0BdSR
a1M0tT6fJXWzAENH2ndMUZDCNCilET5lUE5COp9MGuJt2//uuF07T1pSjfIw
mRtnlwROxo0omAmPTvkrj7P0ItJZcX+MAoNFA8+UMQrOFG+ICVx/4phBYKGu
rfuWmwEnU1EVXirS+hfE83WrqVj7xTj4gPRnKaUGOTLAtcA2/W8q4mCT8pJi
xECBEWrgfX0lfavuB2qdFp8QngfFeX057jEb7ynsAlqYe65QoWOVj0PIzxTu
F02Q4gHYntJxyLZr5AWQVi0wjLmNSWcA3Oyj2RC8E9nd/RzieLEs5ep039xz
ilVNT6eCXfR9iuXTtLP0GSIMXjLwkAyh6UpuwUBRCP1pk/fXSr5CSdRqf5/Z
j4n/eymIXec7/BVO5mrMbYBSbkUE6PPhjSo3hIt24K3BIkLbj4VUgkxAGlaP
Q+UmbQ/luBdzcgSNQ0BRC7AkvYH2ZrDDjficWi7S8eY9WmRMx0CMUfwbrgaL
a8t8i+6Zb9JNXJ6qFkvbaq85dRwWKIXPvPpeLyFGZQf1uxqNXU1jnaclwvt6
9dRKbwhwImNIB56V6Z3uvC0qvIVNLkYG+cwcUGqavF1sv0Jsozex/0f+cg5c
X947zN7fkryslqdF/49W+AX8xSvVcSmVuUn+LzIKepcW2PiJXeedyXVqqlBL
MJXpqxkAMZIKwXIAoxWpWUfbqU5hU2QkJFf+hgl7bfwoe8IHt93QrQZGm4Cj
IZeb+kFGEmDiuXkU5xeFgjIumkzPytWmneuYHVjjEoXPiw7pyUaAfekTiFw5
IS6GMasU5Nv78x3+Hw3S98MyOfVO+yxYkDh7wB/R0TCQCsOam3zBHQ7gaB88
BA6KE/SHBAE9fuqEv9tA4oLqq9I0+fkG++g4jCZLIl602c09rJInAwPdfr/+
eQzEhM3IuXIGHFCTTv8iBNIQkmIGTp+/iB+fTwmcVE+V9T3uTpBBsSZ8vL1F
WjQQkjh7a8qUeaNjtRvc6pmc5R8rVLZi6BTDAumKzOC1tjvBNBePOkWX0PzD
6qmjYnLz9q1sU1Ny8XiF4vY7sS3LgV4Pi0yMo7OhRkPagzm+YCiC75Gnxhf/
e/AADwDx8yz75QMqL6yT0MIQT46mm80/c88vA+A6tK/PVyjqJfkM43ia+zrn
j9mc/42sYaQPYIx5EmhpX9I7YdaMzf7hy/xmwKtVqFNxl8IJ/fX8WRI0C1GE
1OTeTTrxOmBNAaso158ESlzehCBs4ccHffS43tt4udV2OFoNAsOALB4gXMpb
NvHO9KO5zhf03gRZNdBhj50f5vjYcIGiSDUoWkl5O/h8TEIc4+hl/MOGc0uy
wvygiACXpcAVEZghvw2rHNxAROlVIPPRejZy/FRxnepVw2jtqKuiOeJiu1NN
SNwnUKeIQPEXPEKctJCiq8JUx1hxpH1s5gRHYxi0O/VZJTolgJ6WywZFIZAo
jobDdRNXyTwGdy+NgtbyWNwb+pg2UvjUjEeZoYepE/jPIcjK61kXYvcMe9EP
fy6nkU55KYNsrewJayF5TjZUDceW8g2oRHGGgNHvcGZMicBZx3wjvIfkj62j
eA6LGlpYQWKJ3MPHYuTyooYebGRX+oX8nzmu4aeQ2k7dxGTpPOHUvh1brtQL
18GA5NW/HP/evssCvOTB+qNqoq+LzexAn1weZVtcDetxkfKEujYu65Pu6yt2
91lMCZlHvJxX4/GwY3aZ+DGcvhuBJD58bP8DuDLSKmUap34iYanAO1W+UdFJ
e82E4ujDSZIQVKBRgLJ3wOl+3+9mS3B8KEot1/4Mh4Xa/dFkyrBuSYzj02Fb
U3mT/qY8dQT7INipCezNTCpDygU6GpwlNltROdFOQe4cXJ6B9NfI8u0LZV3A
JCZWPZSyoWBkdpt7prSmgE9Zn3ECrhhtssMQJsUEIDDfqWbAMvu5rBbQBxJr
xWMvUZks7ZeDJ7t0Y8J5Te251hEGz6MSjLCh3+SagzNCGoa3Iw/e8c0+hiuj
uoUMV3Vfs+9XmDyxmN4A0QBatmlRu8UI4BMklhQKs1PrMQYqPhcm/uerD1rs
89YglsMIgTZLSSfqOanL9bzcnffDvrIdkR/4nRLYT95SnWkIu76V1a4AKjDG
ObRLO/CJHoY1PJIVVuRcapgy52QrYWB/ygdpw/RHSwUcYE+Ej2BkBWKe8Y/l
nNAHsimHLZ9eo0N5kdCRh68ROFnnElKrl4fP2OLRjF4XD2nrnPL6GZQssEgT
uzv/Vf8u03y/aiy+nrZWNxweoXx0EOphixmJZWgxu2LeWrqTe76gEBX+1RKR
TaYiuJ5euTRqUglcsnbIwE5ONVhpg7HEdAl2Y8Bq/2t0oafaRgZZDkIE7Msv
BBH5C1O3guyvkxZ8Mdvq5siS3vkpg1aeQ4Bk+7Z+4lI6Pv72AZAHraPpqe7I
CIhjctqlWs+Yb0lh/vDXAz/P3dUy197N23beggYel1zZZYhxthlyvS46eLU3
WMmutzz8YLDsk47fOTbNIk6iMe2+xttYKKIyxhbX1ZqXXHCzcW5UcNkBQCNP
nko9B5Y7l4je6QZoBx91hJttT1tAir5CCyheOTY1bwRsngEmdGpptdyn/WYt
jark5cFM4dWVyRPdHSIiq1vAhbegWb42hPunlF3AZjffSNFmkG+Ij9nP9EPC
a2TQeoyH7+e4/hKhK0/Gfg9O0hTu2SiMhjurMlCIpM3yhJepCWVHmbVUQouq
Jwbc6yJVAnS1xCLpz+nQs3hVPPK/rQurSNBoiBSQNaunrrNQDL5+1CRTOBt1
I62ulKZPI/tTaVAJA803pVS6MW2lDwJ9jk+8sW4La2+RJ4Ax+zS5YSmzacDP
IFs3tizaLeiO3u4TOcTQb1aBcL2tpi2BXd0y4rwWba6+g74umM78OhSuN3Rh
PHvbJbX0oxcMY+Gt1b0Tzy+FYqIRX43ivt+VWpECnojI4oLe45Vp72dML6Jm
sn1YMPC77PV9WCDQzh7wyo2RjWf8p8l832jW6wJpOX4g5wzOfWnsh/+xuJ9F
EHZy0e+0AVY8R+FICJNUDiAieEzziwbEM8Z3mNNpFZId2zaX4v7awfuspEz9
I4HVyXVspbv1YY9WPhjnTCcxfuhjq2+1QY42uitvbRLDaj9RY7KNl4kNx+ct
kYW69xatzzjwxbFD70UQb8nlc7p5M5ZmXKOiWg1LxBJBZQcYG7xC5Nx2ihB4
bsryUGIs8+vKCliodlESZNZmErsgexCwwL0s3QFqaU3TK5KvWz9xuLbZ+RXM
dM82zEgfonWV3rjgJWD8bWyJeyg3Mu9bEL5mGXalw56PS+jpZfuQyu5DttoF
KHzbN84PD5dzSQ48yoSSZUfWWupl+e9MI8UTRa7Bqkb3I/IM0VxBtN9gDXFu
+MpsSO8thI4jOVcjGDJZ75jWFC8dPw/sgxV9qyx+JeoDrvo+VC5MlXif741X
6Y11NfGf/xtPvQjFbV50Yj9hGOusQsqpTseJ10HD1ZdBOWqkOA0M+SO3uDvD
RM4TY6qxACV7mtur7GfbHc5M7bFPSo99CJrbRIZWyy3MBVA8ZVh+6YZaYmoA
VDyMcU2q6adqMYR9e+UnILacZiia2z/9dbxKWOOzL4xbZGHgZEJ/JiSHyD6m
regWcAmamlHzJA3/eTehnpvAenS1mPh3lh9R9HKoOu6SUfmj1J2zLaHDRtVZ
kWnTzJGg/Z3e38e8Mlvlx943ZzA1ngPNyq5H3goeockPCzNgV2YEpRE2N4s8
4sDcr+SylMQ1Gyl3IVkbs/YpfaPVrRzgQ5ggwslBCE3OYv1QMKNzy430BpMD
HImSiaHpYYNLHHZf04QA0DHRY4Zm9XfojigEdim5+JqATAjQUZyzEntMjRlE
gnZ9crFB6LWDqX1LKWWL0xVoCcLm36XMmhRuwinlWkhQfPvZYsoREUIrdJz2
V+YQNQMsDOqQ/G2AhLGZh7WR7xYuJp63s+dZjZxvcxih4pv6ZFi/uYJ3jmgi
ZFnJr5FWjIrAGTtEBIYJOJ656dWrFKfz7xUKpc3US+fnkFFeaBH8H7IpOvX+
WsgvLce8/Lkzg0D9She2XCcfUFTM0wBVqC5RLhWXdfcg0i/FqpYN/kMKCZmU
OLJKfsYm8aZ8GBgvHuKBzHpzBlzV/kp/q6YeMm7d4SCBJ6hzZnlViTogR/xT
nIrlyYAL+07V1s9wWccAkcYll3BHyOvoRz9t/AEvgNJUZOH5iC/6pU+vTvUm
H4coae/wsA1Zs0ByAR34YXRitNdW/uXAnx2BYV7vmYFkGNZ8Czq62OsbUpf2
7IoLERiN9bhbfAmrJ4+JS2B9QRp2F5N3rOxOgrHVOcyvvf77kVSr8zTFqG3b
ytj9k+quPap20Hny4SLcYFhlqMviwN5zTBxWlRJbBxANSeWthIRBnH3nbfTm
oz9PMIHV4YrTyaj8/8oCWN8kP07Blu/I9E+KddrsdLaa8ARDDGuU/OElqIuo
vKzPgg9gIObXf3kEfz5C0NNmyXrwieelWtpiMvXE7dv0sgBsOMaq3OvIfJw0
9TDP4TYXuaA3AKWQ6Bab/ZRlXYkTTZqwvUgus1KbJXyC6FWRhLzRXYUS0BJe
i8GQsHtUNClGDkyLm0nB1vBLJewcRpkgkRfSTo/lpnCNxeP5yW7BOydNH9ds
tnP8DxYTAOD5iUIgI3v5KOXAMjYRG1r7hECli7ddI6zOgSMTB37QP17ejW75
U2vp1qQq+a+kD+tWLb+Is7KRRn6exGIhwP1bMP9a27XgpuitMXT0sobDSBzY
kvap2RS2uBlFTrhGPw7Zu4YDffJJiyEgNXGX7cvz+NMAtWo4R12fY5Cfmy+z
dkA883OVP6LulIBnh63s0O6V92xg4kSZ8cpB0PiJ0Nm7KhdILEJfB5KOqWrY
qkdINk5i5ecXGYDkrE12NdTv4MrmIKS9wE9H8tUiL2ZCAtq2w7HWtAO5+nJz
MXuZYxo2MqpxVPI7tdj7vjqUlv+vEqAPXdocCmlvBEBt9DYMof/GnpuI8cPY
0+th4vIXeusuRx2KWCrZ6NsmpsE9dBBLCYA9YuV2tXk7oI0apmUqNyN4++90
smL4Xt1hiYKC1xnMJfj+GCjZv/a8QE+BHe5+Mv3MFTm0WKxxOy60PuMqmTLw
iJgkwl2jezdlBQB+77P+SYHgQvx6CQuy32XcnXmn0YmFiK15upEy/15v/5N9
TUpcb4dOjUDOMzWBvdtpbjyzxv+VK7q/vVoeZig5ebR7fRhaAL/hHOXVBAmk
sCnYU0Ti8MPJG5FJOCvA40yPsgcPgJI+iUoSGDsoLTwvnNDqXTBmjTN9rAAX
WjSUryFcsR62vHEwtgwjYk1L732GFRSMDKCLJ4QjWRPgcu5Z5TAbx7TztVN+
o2NyEWsjSvhMP8PZzuJ26SzWv6b8pbUFA/F6fGMHPC5p5CZA7NNU4QouYW6R
dPqvIu44qYcqixVOsDj01EqadB4u29zh9PDiolvWlAsgF/3uBfE5Wm/rsi9t
uODSKZ4qzCHMiJUhQ6Igv2Ndw/9L+aurCXtUWNNSk7IlIRpKFClHkDl63ntC
N1OusnxjDTBrRIjIEiIxRLMSPG4wZQTNDd54+727GTtgvnrngM3x1kMofyDS
VDPjqCBPTBUXb5fZ5wMqV5Opg3kJW9ErtNODVJjd8hiBn4FzL8rs1VygpwoV
q31tM7F1apDori4IjnWjK7VcK7sYk0dKoG9X3ZNJCoWP8iFIF6flvH/3CgC1
U7WyTakv3kq+KnYvGmtyLjeK0JJU9DL+/qqDlM/jTwre9UU3mMxg+E9AXCZX
hDLxhbi0Iho/3Uf1UhsLCSNxGEX9VqqFRzXY+CvN+Hu/zRviEu8zsB2hSyEq
hy3/a1G67/A3fwwixyKiMxYDuKk6WJ1tVEGAhxUOhUTr8ubQThjCgH/LHvzz
AuojZ8j4NQgFlya9XHlorr5q4M+3aT4ok7ah1+7r6jo8emTMrusFnS/za2o4
v8Ij9RsISRbmPDmYtuC3EUz9Ta2Eu1pGmWLdUcG0E78Y+RZDh2EXeqd1ONBi
o4YEh8kYVDQlzuLL3L5/tJIQ156df/b6ZSJBtQ4BrT2SId48LnqFa6LtzLIw
BBXoRFrNsaHsNVWdOtoIcEWsOMJDoBvbHeJvv18hdbKlVvRHbIM8U69LwMCI
Sp0djSYbLTUSFX5drVb0cDEYHwx7jHJL/OxGToll1DYZDx+63eMpVX81cE4w
cCxCfrfzwwCXWL6YDyIfxMW9nIACkiSdMmjXMDlQP7L1STb+ghJY5lWSnC8s
2oY7ktEM0uaXb45v82gP8ayj5/EE8+AuvXdEuPpE+3exClO49xOLf+HN/9O1
gA6Eflxi/57wxfn14NGP/LCdlNHWwky62FEIyqRPIi88rk/YSvhOLEaoIJR8
BeLWl9UzV9NkQOFXQQ5/wER39NJ2AtPOY8rHFhe9o3mwbcCeTjt0Ljv4srBo
MsHYMBt2Qs0wWbMYNnDHKIcXTuf1dbRvD4kzXXN08FrZi+LJc7ZN3+tzHYNI
UWaab7QKZYgiiIyLUNOeAJ1K+Ff8ALuCc5XW9Nfc9N9ccBBszPdFJ/FExk+Y
VUFTl6LG4Lseog7QkPj2eznQQ9L+3SpF5x3iumFyGDnU6bMADmj0XhNJAEe4
y+ZhgbFokppH3VAw5i/OcE49mcGt58Crr6CzyWQWJz8HKmOPbDfc1vMphRZO
BlqIxNivkpWM86XPpQUVZP8be9y5HTaaix9nhKGM0r98Eyne8gWKG35BNizx
gtPH9BPZeR+QS1uhP7A3IfjEy6dqMmuK33LlRDEM9tv1ZfJniAETIomzinGO
fw+FhT0xd1VGFDAMSS3R19hp/DWLCXjSlM60n+jtLQpreKxyIqw7hR4+lxwn
7OFBnGPZ3O5Rak8lDGo4u8qWckjQF3cWHqRHxp2/2aP3WZUVbCGhMPSpJSpt
upw3TyZvdEMJShlRNkg9OQcKjBi4oCFoubFe2JAXpmM5U0N3Rv0eWVNAejEX
mNpWKFm1h/wtJCHMGdkyP2bAaQv2FubarEnQ9U3fiTlGm+1Q1cZZkMrGY2st
r7ZnQY1b1K6r1s6Wn51mZRS/Mrv2mfAvFOnD9dRLtDh6owowAJWVYsi9pXDU
dQVrOR00bJTNCGxEXQhf3A41Hn2qi3jOrNUOqsRR2G2kHG5LXLpXmXBXB5bM
qP/RWHlP/uTF6etVfXRoUDyToRIUkWH+XR2AKtYP/+68m+Eu9CRorI4Eu6r1
eD/wFxUsx8BAY45BNvuwVI7fEdVheCEypA6mUxB6sjAVTqK3wFyHtlPC+VlP
8pzTAelZPuuzH3xxvfyC7BWQWWkZ4VLjgpR+TcyphNIR1EJA1my/XnVIBaKd
hTrU4cUmO9965FSySkcM668yvYDN5c2aaUvGDIgs8y+0xfBw0ETxnshz3d62
7o1JCEEDBrTgNbRsW9UYYcbHOQCTlncJSPQsLGD5vWXPU1AHMSYsbskaHrEM
yY7kCT6aDJRDXg5UIDr46HpNo8XqrMRtrePWeGcSoEoGW9WaZwoXWfoAeL4I
vxex7Ur7Byzq3Us37uglPF3mFNxSA6Wb2HiOhXPdhn0TcxflRm/OxhZgovU6
uqSOMuNvvJNw/9vnGOKxmYJ0pkind+Pr5+hRNtrvDv0r5Vl7OcD2UGNPHsf9
+gfKB8yUS9mfxKg67NcnF2l3242ZdT9FAkJMceWX0Vzvlg7Sdx5Pa6z/45dS
mC2ACcFT0dmW3qC4jD0GN5ONhyxX0E7MGdR4sSZIaoHQQtK3OXx7/5gyYfLh
aujyISZ0icY9eXzuFhbeqNslpCyNn1pzrhbf6IIyEPD4vMp3ATAayzuPRcQU
J/rvGYKKBCqLdgUd75dQ/Lqyt/MvJZgHdYze4tORWd4EW2f62OtcyHIyY6WK
Z8NHAMeK/9T0rtD3xXorgQbQmkVxtKgBDpoj5Rcd4oz3kTGdRujcC1YYxQ4O
wTfpc35IxLdpaYsqArqBA8uORMNx8xyesGcxP/LNUedEU2Dq0guMCggkSgVR
J1UBB129go18PC9Fwhnir8CUGIzgu/ARS4SZCMiycPWL2haGEJJjUzr8pQ/B
DmgFR+HRUR3Z7B8E63auYOiz7RewXjN8TMy1eMJnxHc152WQA8McBrqo3YRu
V1jlGac9pEj6UrnDylA0/dlVQzsrxi4OjVbOzrGGzwfICful30n6qMikQEm5
FXh+/fS/TvlfTeo62XiQcUCXT2O2g2Oas0XSifkxa8Q2I5JP8NT5BsYb5YtV
DxFt2WnCVxgTANsPoLO2lN4Pu/aNnqtNaaC49dukpEPYlJIF1/ATK3jNqt7h
S6BQQseqP5jXrx471YKWiSZS8BaBM3C2U2U29r5ITKtM1P/ZZ3Jli2KXAtWu
XaxWoU+vmeBzNUOfQ+lVh4OzlGyKnMOpa6Sh8PgAuCdil4xUOOFEmTW08wQk
kFRIjAF56eWMYiMAp7ecFozR9/YUtpGtNo0+ogaxro81dRUVrXvZg5zw7Gvs
bOFyklU7C6oa+dQsrIu8h5ltUreWg8rsQT3GIAfEQPDpAqYUw5v6A27VCxWE
FV5L4NXkyXmRH3A5yZq045j9UgFwmymz13xfCdvyhJGTKpzvLarMc5nGYC6x
2v902CQJa9dUR5Avy7Rwzdx1PTfpNi4rly97pAtYFOdfh+YOnU5k/raUp4QY
+DK4HhNRpNcFnTvg8Vk5Ej8ca1CsjKI8V4JZd2Mtpyqv7p5ixfajc18Zgrwq
tl9N/W0/Qo05nkzkNktElYg/M8Mv1LxbiCujMQPkwBJ/+HkXC6+f1VAPeUlH
/Miva5WVBGwxjTQG4qX0eXLYWKVknIB0/t72cUJmOIwYk/UqRMuHj6u47iP9
jJJ87QN7G8XtiufNlTT/OalhMQc0G8sLLPF7/c8lwHkoumllqiZjRyzldAlN
CucdIrxj69pr5ZMXDAuEWpcuzSWHhG7TktHEqHVkT6q0ljPE4ZCaRBRobE3q
m2YHbv/lIzKqNAOUNmO10hu1irsYasqgNX3J3gZDSFJwUErXV5UTW6gAYUzI
A6WY6AKyD/4gG8x28GVmtk2BUSvtbrhr+YJq0B1As6XMQbQC2HDcPNABmpYt
oEISI9FKdDNxlc5OEnLOgZ3ChyqRBnl6jIJYywSluFV8zX3f75Px7VG5k/uQ
9hx8d2J4SvzXB/VJSBQOKvkIQ1KkthTyKbGxJcs+qSsgmkz+EVgss3jLbUAa
W/joNdVDYHtmkqwWpqbQmJpRO+SgGQIgcgqzCqyMYszP8Q3/jXFMOS4bDrFf
xw01w8WM/4ZQE7KTb61LHraGxOkExBha/7MhC3aei21SysAX53vhms0k6Nwe
nShIaoLlT/7PRSzyEe5mhpuXOIIOiT+Np6jREvsWvm+iNkuhiquCujxkb30Y
HQ4H2t2g4ruULFfTv480a4gDWbPJmzh5QteoaPFPKsRYfguOEsHHnt3XFaBi
kgfYbH41/d6DcCinDLhY7wsGQn1HEp7ou9zVeBTR8rGYTSR1lBOV9redAWbw
eaHLIUW9zt3F1qkmwagMvTnhMYkkuqlwGvGiOR4E8D55Kjnw55N+mruobLaN
EJ404gDNzLi0K5KlBZHjJxKfuA+M6+ZLYWh22dL+RtAD7j11O41i5G6A5+DS
9BV0zgDj9tra7R1bBjpUcoal3ubd+Iu2Orn6g08aXBmOKv16SgsoMAll2svn
wwcJ3xqvEYEMgQIe2FmI36pJ9V9JVDfpXjf5FYRhYlP+zuG+bN5BSgOmB19+
BmSyJt0y/o6+TEFspusVB1EOtGPvdUP/2H2NzTl5CKe0dVOCQ7Z719NWHhkT
MIOLwlnlP7JA8UaSZCSN/QhAjzR6J+BkSlbrPrjbpnvBMJ0MHqx2SLQUlzhb
9vUFdEnFyyGyoSMSqdai8eudb95Cr239pO5QIYy01Mmgx50ErTai3ksodx8Q
Dr2bKiT2LH0kIxTuIS9QQUHexj5Txlh9lrerG/cd5QOuTj1VLfaMS7hG10An
0IF+VxEZMzZN5916HiJlz0y7mgxxl/QJq1UbEdWDuC79FFNuKxfwcvQhpMpz
X4sE6+H+jNXBkl3gXgsP2ixCZxF21Sahjh6Hb34xX2gy5jkCx81BjiHV5bGH
K3zGwX+KCCy3qrN9nzjM4mTW8clUSvlNlAFodoDFTcn+8SgAEPsXlINZoaZv
C3rc1SEfZse92oClo/xEHJxc98NToiAHlWb2dMCK/PcTP+/4/BXYCslWFxmC
HbFjibiFeyHDoJURJiRNXE4AkZJNJ3HQ8UKOJqYE82UwYNW9aYKMaktYMZBn
m5C4lYu0BeCID1XxPmB1qK5r4P7inWOGTnC1MREKUq6ngUL3FFsltwJMvflH
5GFpxHDlSqcnUgrnr22mHplTF+TN5L1h0fq0Sknr8fWB5mgOi4keN1E9LGYQ
7vp4hbtdotbDEt0pwvvOJ5qwhgGIzFAY4fhOlAlXK3ENdr66MjoydLDaOQxl
zbghsGWlLfsJb2mtWTqv9YLVgmDAghexxrOQ2Bb0FMkCOkt7una5cjQwIyVX
2yv8e7/zd0iniB055V1YubAinI1QUEAxvo50w2dS1KvnI27RtSrvUdjavTAK
YYjtTsQf8BR7u0uWB9FsKpW3YiJ9lcMhER3eNaJakeBvtJ6s8dU3XCx0T/S9
76BMs2SOTGUQ4U3XY7saphjrHRN7NHfaq4Obbc4OtjqZlwxLeK2eb1ihzunT
qqMY89X5RHxgrGxv10KzT4ppoqRBuyCcmm3eR9rS2ZwYZWNa9tvyUOrXq9im
LXe5U2eetihhy9d8DrsZpL+TOcdyqQe5JSOwMcRWyAUSY33MpEGu4t6gde7r
0Lgrz3gm2kB16F9EGD+YM7pqM+KeoRcPolT7cIutIaO6c88OkWEshSByNpDk
Z0Hc2bf5g8RMYQynXEwyNTmhfVe4+xf3oX0rZbwRWc0iylbC58/HzGsmb3n5
R6fZeAAX4GJeaJRGtPShWoyJAX4refMAu8loWbopqnDQG84G+ZxZeguF2Uvn
2gAOswRq3HkjWeI+XU9S3setxc38vQGPZ+GjnNf0hb964BofXqX+kajKlfLC
Go5pkhJ0nQQhq/N4WNIEgQzJCyrqcCbr8R9MB0ri+6unqJxVKtkVbQ9aW/kL
7uAWq2NqDUYu04OV611GZIlzgMVCv976F9MFQzw0hzyDwzCZqwgCtN+tA22x
zkYNb/tC8zFIAiYEA/6LUd9vrT1LoV+sP/i0g74IkqiL8EV+DCdyDQEy30Dm
GMW7I+5Cm3FsJy9BkP+s4HT0jkJ7qaxijRCjpxFIeL1HAvUW31vrVPVfQqgd
jDJuQPi0jpP48LN2+C8GNWBXTMu2n8deK3/ZUTiSkqG9RVIc+lYDkF9287GQ
HqqKtB72nS+SX9yHlnL6lJkorkGLhHumgIFX3c5YasLxIzGCdGSWfCrJD0Mq
b/P4Zz7RrdFzJg7z7oRZZgjk1IFxOtcpnayG7q/D0i3lT1DgWPvQM+J9c2UM
7RAXpkcl6VImidpEOwvsncd10DPaB+t2WRFVFR0krdCIm235Es0ecg7zv3Fp
dTO5T2m9v6J0pic1LtNPbXS09vVp2jy5sl37roJuNE3Wrz6PtxZsc/OyiC4s
nWQXNuiORgcKOM9fwzXNOeTmaB5oeOM3cEeSwa49HRlRWrCT+InyFk1rY2Rw
0ndvx2WJy6lPJL0TSRU6epTjuRmtWYLld9qOkXpI/GZ1fd6W1FQQOrhtQlq6
Sp+3gryvvcJuSIlFQM2goeo7mTn4ChJvFvz774Mhukcrnx7vg0J+OQOcBZ3L
mqvSm5g4NUeu4yK3dNQqNpHUQzkjz2+pEtgvfwNOUFHmBxxmSZP+HH/v1Hh/
SE3PQvMu44Vns0cbgwtWBb7GSSB5ZbKSkdSKeeUv4k0lu+FzfsMy7ReR5cyo
xqsTfhITWfs3hf2/DCEs3E1n9Ws0s2NE5AdLyl8fRAeXGxHM6r53x3e22hhn
L1FuYGmuqPdMUcJnAGuQ2GxJbgk49muJWjUjJzQhxBXIhyqKcA6EoAcPrwLY
Qvejnr6KtyIdCpmmq5WnmmzCyzhJMwQfoC5IsKLDHxtSYEDsYSFnO34ZT8NC
oQukfoMVThH1S47kNcTFgD1WncQnT1lnOcIs+31U3OYl00eCSFC9ICjfkBHd
A3FbV41QJOBInG3Z4iMi3vsBFxGD1YBqEo7Izz8yUHb9lFYQf1kz8lGq+wz1
W2/cUwawGoNq2uhnvfztm/qejxenZlqAttk7QwUkbtKkBnBKXoGq7DM9gqkd
TbTdPN3qHl9ynfv6/E7b7CIYatqScbjFt2UM1oYehDydTxdB0Kk8mFcv6jYz
Hr/9Oe55ckPmZtpA5AE74MSiIxIs8ASxbaCq09pUUR9FatMhxrgEmNzb2MLv
2K9BmwSVvlUd4yRESvwBJEi1tZ9qnJPvs9aAxO+cp/xMdFrI1lc3S1HF8U/x
7jx8VZgtm/2y0UhYnbp4omdBJjFMx7nCLdzsrIr4aa0r4NZ8KbF/ONgnrHMy
RQDYWpOIXMO9cGycCsSUvp2Rhr/wCTpuzZNIr0pKs2FSKHjb1DxYv9SAody0
UijLWpdw/93AYg7s7RntnFAfoB2i5HhQAaGq0AHaJ44XHjSU6PoAgqBgl0y3
rEqGBgfaMFu3L8VrlusgopXvb+t3+nWiVFwk7Utc82aAPjtcIQpOvPr12blZ
oqYIqYi8tpjBga2PowVURZzVd5Zr8vJe4f6vhxXQeNZK6n80m7LSbEZKow79
9m538p6Sio08XkArJVamMeD2XIcM8RV+2gjqTLAorX7Hnq66JubrcpmWYZaJ
m/H7NEJoTULx+cORcLC1UaC4SvkqoJnsJjZ1ntzBlAfIuOWsvjACRjutjNor
Cn13cuRfXDtFd7LPitnlVTnNaY9QV0l3Fw2W6T+gJHWtOhXiYgD5HA/Wmoyu
pLn6uxm4bUWN+Wo1AJ2y8V2Ez6TURmn3WOgguZPUT9OqgHhqaUj03v5omfEN
SORtOXRrsb1a/6vgYZh8pXlgdonRN6etMjw2ibukbQqb58stFw5kOJS7cpAu
d6Zhn+oQJRp9fAXwA/Khlw9PXrqg7aUupcBNgAhqqOsSgE5y62mrh0sguxdw
QzYzFK0YRQFzOjZiZiw3XftoN/DrOnjQKuCoJZ9cTf2i+33+pmY6trlteXmg
EVxmfaNyunRfPc2Jv/M8An6wDTwzWK7Ib0OKo53S16pAWXcbwGhkEgYXvd0m
s1Ik5p7loal0FTmVVj2IOr7xOlQ3l15BDoxe1BgnPkBEeR8rq9h9eFYe/4Da
YZdPVMnQI1vKIBkbrbuX6W1Qi1meVeyvtcWZIBWVLt78WHNKm8zsjoD2s3EI
2i+9FaLzwPGgpSTXLtYsmqZRMdhb18yiz5oqH5M8FjOHbg4oVHiz8/8/5qbY
nWfCAu/bzx9NGa3U2zS01e/s621Nl9VKkThX5AStDTPPcJ3E3GOTHro+pPG1
psIKJXsn0Z3R55I8a1Pnkh4iqtO/+X397rQUB91w0VCiTIvWmOidr35AZYk2
jOVRmuZTmPQ4mZJoCMWHo0a7y5X8bB1r0vNmowKeSJE37FUeDxZxqL/OvZT3
wolk5A7/UHZ0Dn6NNirm33x6WLweQzG+v4wRWEhOOA9vbR9rWB8S+fHXJD2U
OWdaF3oXbQXve/Vc7MD96BeV0ysr/uWcgbXHenxdyMx54IwPnmXgoxDLS2jc
2goO4lpbkW4A3rSsd+4iUPFEgOKugVFN0O4PTjh5SSQJtpCo2pYQ1QLgq5t0
ytCdaadfb5OLQTuCrpoETd158XjcoskqNuQfARXfJXrCMZJ3DnwJlLgOauNN
3u2ieFwlNXkD4Q+vUeGpJSJZ8z5d3zr3P/OCHyqw6Mem6Y7ksl8D7oanqA4z
3LCIDCRzEKupGUQ4v9cNLEQtHGsDT0gUpg0GiW+7H3KJpneGan+KOlI2LECU
BB1znWZ1OJkZJdCxaBmDKMEvglwMM2ifdNe+Y4Tn6B5VstuG1+1Txw6If4ui
ZDmiEU0m0pYXmWm1A5pZNrGZ5jc79Q9pGbJeQYBbWljND6SMCW6OCxZWzHJ3
CGTlwCEZ67EFzsXZJ/w3syOYYpzTAEo3Pe89kRY2j0Z0JzyC0lLUSqkF3JRn
eqBUkJwZGdE+osDIFc3kapHreed2XBrkitKyu6vdGgV9l1j55SYT1couX/c3
dRmkFn76jlZclTOAR9cEnQsYchDyJvWyS8gAbzASJ2BWsvCL+3ei4cnAsJg/
u68kAC4P7B6ykPpsXlIom24ayZEfhoBJnchiolLg6sC9j4i9kPj7oTD7tUFZ
ukJDwb4CpW222NXLtDjHMARKSePabyNEl/xOgLihRSwuY/UPi+9jVfcchVZ0
l92iL7N8PaDpIZ2+qiILm7TvuM/YSCOIqkyY5IPd+hQJuAZa22ExG+8dSC7V
V36figlK3rCjEm5a5FO3GZKaGomirXp94BFGj1ucThFbsRKBGSFfSNDOP7VN
xg/oNU6cQBZwamDxlE4VdYSLfjkjS+Mi+q270HtcfQri4Q2C/c0lS3mBhnRe
DYPIAIEgRYdgTsD4Tz2/cd10Ekb5153xhMoJ+9dIB3E3Y6lWQmFmQYcWakST
xhhmmN2CXyGUf6/T3K0eeM2UNpoYa7RskkCj9vO4KuGcYgV9k8sApaISj/wm
J4q5P8P4JcFCcigv8bCKAAs5+1rciKY5JwaBF6xoRE5OV+2hu/ilqJDYR8Qr
hbjpsyxOIcJ77yVbcI11NbiNkNUFajHzyJG0VZuYGBEYO1c8zmVe2U+2WJI5
Zoc1FAGw/eq0dQ1UMk69wactSeojS1/0KwqFg1XVujC7XMxN21cmjhkrlntR
gZaIs1xr+iQLwmJz3dm9GeLJ2VvK1vCCmflh4ZpogpZNbbJlBCgQ4GtyhU0O
VQcBAqbQsJRZKkHGxrTU0O1cFln6xgaj8Zm+BQi3xQZz/K7rQ+gNFYFKOACG
Z+BDFQht7I8on1LPxfx2WL0VLkT7Cm3l47m5H5xytrMwIoN39uxz5IeHwJ8n
ArhIJj1/DbA32sjbtmdFl1d5THz8Y/caNQx6y+AoiGbLsY6eqKtOUzsE/PEZ
gfkA5k2wa1ExR9OV4WzPns++ERva9Gy+aIfE1AnqQZzuMDCXYGMxJdEZVAFN
/lm0qfv1k6G5Zbh1hSaKvs9BTjh/JoZWBncc8bqgEIXjofHZ37iQZAb/ZR5C
kY7W7D5okdw1I573fCQw+0HOuQZeAoIafHIbdosX6Kwo+ku8iB+LinlbO6ZC
Q4INxQUosA+a0Fj8nTM99h3yTXKueHEwJ2FxNsoDvb4YqrQe8xdqcbp/pvzy
n5JJomD2MMGOpTJKT4thMP2n3Bk5uqR8n1ccMFx8c8ke5t21+dipMOKyo323
53Z1YUaGdbhl2VTM9g0mvIHc5yOJt1nSDJ6P+TvkjUr/2753al5MhnrztMJh
l0rAeCPSPSlk0HGcuhrv6YTY6Br20b6dRX9czrVJGROAnnWN8QC+AvOP1nBs
vmqzEehyfo7nKa4jtiKeSCb4kwb7LqdT/tERHNYzrHQvdVzZj6c/wUtw6r4T
HmxaNbCS8SZh0Pf76XiLxGBZ+yIrAewfchf2odpLxVcWcIRnfRlD++Sy2j1k
Ic30ahrUXLb4afQsIvX3/lYgBfz3OCt13kZk6GK2kOnvKyoQm7WNjvPD5xp+
0ZMxSq1HYn7bjbNfdwXmCS5nJ/dN8VEO2E4LfLzb5dMWjrwAdl6xuMLwBlFh
/QTNt7Gb4n4HI9N5NIUjcrQSkpCLbnew6zZlahXkm5/fF8HxWsP0wFwuhdjS
N3/BK2vdr84Fi3MXk9jz/a1ilT0GRSGKkzZSRewPuFKtLCiRDdHgIxuFF83C
nP8cairbV6cmS0jQZpNPZX15XuXIYnr05Tg11lUN/LLDhsALsGroUvZ/QlMB
2AqaDsbl7eg6aDXt+m+qfqFI6I323LfJK2qXnmLJh1gFnnJpXn16u8xo6TM6
R7ruaKkeYnxIOiDeFiVG3ucM6stb0XnXBUf5ehtI1xDzF+8XfWBp7gq7PFk3
lNcXLC/taM9gscti0LnG9OG2AgCu9blOZfWnNmoNZ363p4+yGfj8B13iG3Iv
YXWh0UAB4zzwLn3RgtO7yZBguqKfzOqO2zdiDlQ1lX/hBH7Jl2F606KwN+6O
dZFe66Pexrwy2TZG8RQdfbw2k99Wk2ptYS9riWn2/NBtSDhXbTxf875IK7GK
VVO2kFH3U+Z/wvJbGUUAakj/WNmV4atTNd3Uipv6aPjKt9k7oPyps8iiGMmj
uwqPURT9i7GOlF07fRQ1kRXwXBZ8ixL7NImr6h62BT43EP3PZyspRavqFE9r
kURCiTNlxbuRKjeHf5iyq92AAe+2hvMuzp2v7FFbfK9MqA2Gv72pYdruQEWo
kbL1+zR3r01ucvj4oRWLNuO4JJYNhdAy2c3898r/om0XC4W3WwdZymDbYNn+
+EtvA3rGL9oed0UgObv44h6VUbCBtp23D9B/SInciXRVVU0jYw1Y2YcsOgNd
etl1YgCy+9jAmiRV68TqNc8EfUgI2sinsVJbOSLowC4bWVnf6O+seg/IJZ7U
HPlWu6NW4/srpUUJk/mNW6nhSE/ymV5hmfzeGWYvMSXhw67FBoJykqzBKSo1
leav9JmS2XnXL8wx06K7oTA5nem7wbj/R4Qqj74jwaP9SLCH08pXqqVLqwf/
bEn9poDALvUY6eGW+N3DA4BYvvRj3EW+QLPjsTH0Nq06yqyDUAn8cyXj9xMm
vRFLCzdQh8qtT6JKF+c1iq3Na9tJvAFF+DKHvrO0JZGO/EWOC/Mw6yzvDRE1
4VH0s3KkAtrEYUrEERak/E5CnNB8y80G3IyL+niIiw9K9ELfGgb/vzfISFf3
UYeIjwRESn2LmDvBQJw1vfQMbzYkmW28kdZOvijnszHMpa97kVhB6NgLb0RP
HX9NSOftexoN7MhhByVu6JjhxevPXCGbzKTESATUlqDBF3mY5LjRMl4XwkpU
IU3dgn5nC/bfpTaptukK3XBn7ifP4R7+e7lSHI/pvw0TapdF/jKvXk180mFb
b4ZTQTzLTtUezvo8gI0lApkUdxApE7JvsfljBys+azAUvnMtTFjs/gEpemm3
3A0+SGaKfVrVWlOay4W2vIagLbQGvJvAsdPYg5unzAUwpPfnbSgA9NvDd3/Q
898C/Ac+onLNoQ0JnI1UVKBvT3hRPOwIrKXEUg8fC5UNBnJMHM35HeUEKQhM
gpKMdxyDEcz2IZ65sS70ctPIMVZ4Hw8hKo0ecvXsv6SRVv7DMd/PRK2CJ3Ir
iTevaaeklofPQBdkKRLWyMgwDDs8cz2iAVSg25GviwGvIcq7tdskb+vtno9N
pPaS61iErRWbzfREmDxYU8YJ04aXYBI/Yvri2CGZzOY44kOx0jlawc1jopje
5r7Ea2RpHcX9mgNCiB1YCwEyToRop9i2YMszVeTagsz2HQwV4FrtoMtKRC9p
cvCuP7yAZSILxi4Egq5B++S5utLIihNgQPZIxHzFjuYTO6FsNG+Ln7bbjFS9
ikmll/dLmDkGdjVnWbKGaH4MF3+CwubiUSktRTyPTl7dTnc7hlcOE/LncChr
f1jDa9xtu/GWVyxgBAGvfY/GbFOOwYyV+55NnL/2Bw107kHij2r8rEIh4S7B
1I490p+2ALc+w3pMpssE/ps0cnvJYmHToPr0KA4Nap2d88/1E1tPhaXXg9cl
GEE+swpPL4QvIea5Nfh7gvfaImIXU4M8Q1ZPwab50bsgQnu9QarneWNhZoLP
wfgqQ0xMaaQf/1gutyFJJw4Cs/p1TDNS/8c9GHzegDwe/oxvv0CydX3Ijen4
sEpwBwmDBUNu4fqyHJxwyi1ZCqfVb8k/yFKic3wcE9LlFfiSdG6IO5aGPtxI
oJZXfbNapfOZ5vhQALQXzMZb5ifZwjbWtfHRLvq9yzTzkUQ3g8BbEJOmEKFx
qalR9m3eADrKqD/Rb9jAWgXsqsgPCl8E6aatkUQxkPMNOrQDrPqAVQTxHUIw
2oZjA3H9bQKavS79yBZSkm98OOqalxxzrb6+Xw3XYwlrV7AhjG3ZtWbLjbdR
APsot41WmwMjF1tue8XDa3UbBEpt+Kwh3CIrCVc5zbMnarYhyWfVkXZ3Ci+J
zNje3qy0IOaZMTyVJnsrNxdXI5rCQHrTa4Q6OgvGU3MdX7sHjYJ0jQJAWDgh
HmB5hskHDQnw/oWVyXzfQme7DDLfOnYDqbCPe1XxCrKyUZl7kTt/oUbaoBUM
h5QE95a5oxvb1zAgCK2ZKzOOwl89rldwwHwaLRAPE0KKlBihZneWZigZDVug
EvT1lRr05ekhYxnXnvtwlrIgy4q+QEwjSrjwkNhql5MoYewtoyV1gigGfo4x
2pVvFEL8GmCDtHgF2nRCtiyhMOFrnRsG78/jn98cpsW1KQhlZpS//lBLYx9i
i0syIheOgIP/xmrTgtQOv0ZRloOflpdtGwLjXgF0NU9XttBn1FF7vhyjRhpF
f/mkAjuA7MmOeLB1kFkhNRc8TzD/FZR6YYI1FvaWn18eXxP4wqTxfLuXFCzo
cUHSZIsByM+qYvyv94VmsCKwfpfabrAqu765xI3jrVueNgjV7kPCrDrruDwb
18xeOuw087AP4yOHY9nx4QlQi5vn8XSuqAHy8SrKOgM60rJwReFjazDyoDHW
11RdSsKWWiPBVLuLfIt84Fa9Dg14UOe/NB6Sb+OxAT6CjaZmKepyx/QjHlWD
5sNMmt4ukt0hF4EqEPvaV5POK6Wkv3sAwI7clNP7V/CWcKPk/pDG4zn8JvRW
arXMuiVd1V2H/do8BmM+j8g75jDhtqTUbHMytztmS+zv/o0Z/HTwEMZh

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzehCgVkviA+W8vYo16pPLrsD7wKOKdNkWpduCmt0YAEd6Z0KKWhDdDUTwz4A/toQlEmxSJ3aDv73+RqK1JIJoIKjw3cdj3CIrZ18JxgtOVVXv4G/QCLXaHmleRh1svs+fwSReI5nC9rpyJ6UUOM5+EXiE2zMYeeIrZ9FEQhAHVzLIl0nU4NaRG7ySFrQrtQSYJFm4lKWB04ndBRGrWHiQg19TucfiOuFDihLQw0FTGoL01Tq9E5yQtkeGOnXs3uTUsPqvDS3BWG6q8drHpo+jv/BFgMVzpJ4L72T4DvOrBXSTmlwDmqDJUids9QB7w0Btazk7qa8fGRIkWg5UnuoLAZt1gtqFZWv+jbwrZEb5EaP2iaRLqPa+DoxUzn3Uea7UFP1uSM0tonAG5a2y0d6xNcNEni3eKQcf1Xf7qvIrz32E9/v2q1TRT1ggk1XFl6U0uriiwDE5FyaUX34/E6A6kWmpVFfXbUa9eb9EvzXx5icHGjs2EFrBiFd4fmPVps6ZGUTiF61z0lYR/YaGc3UcoPsLOYmexc92GoWLUoDvizR89Vlsycw6yz4QA7cAyMqOtt9YCiDkIRP5YVSAk/i8UduRBn5vErIhlgAKH0Yir2w2WxBus3A6wIeS/zo3sTls57oRwMbfUF29rLSEMu7WPkeEDluLGqlt8AAryZ9NftVUFb1ZyH/e2SuLONRop/D+U8d/OkVMM6YpjPkxZUcBgeCT52rBQ5bjUC5o0fBrIjotkzZ4m/tQwoX6Sxcf+82RJ7MG0jhcsRwRIY1PmdGoLj"
`endif