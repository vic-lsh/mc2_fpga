// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AIqOD3RvuHPmaIcCrLy0MxPFDWQyn2x/ZUfKJslL7/V+GV+/jfZXEblcor/Q
O3jIK7np+Joz3ruCoX/ePOR4lJ9H3NeJhon//l7qqHA2D+ZV82UmUzTNaFBW
+sxNhMYoeVTKMSEW8hvy3Flz64aP+T2qQj1Qzu2pqC5sq1cGnczB+yLVIcIk
HGUOSHk89MEg2rm2ROWCr0/ttV1Hd+jkB6qA1JFoKvytJDbSCUCz5r06WdIq
J4M4OMt6JBharY+3GAaiUwnI8SfwGN18Xfqww7TPqyLk1cGlg1CGwLU/mPQY
apAje9ZiTAoggM96h+LoyZrfiXYg43SKQQ4F0FM7+Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
geN5lojcjF1QkDfU+JiMQHZef57Y0xX4kgt3tzkF/4U0Ya7obQjwGOEIrUhq
QgnWRaOrx1aaE+fZ9FoZXoYFPxFtMqelyuKDKEIIhvEfibyWie+pjDvGWcUE
IkJkY8OZP0nr6pCGXNUzJzlPyAiYxl6Rs6AyCoyTfuq8IjNzkMkWAvUdhS0y
8j9AlxcA6uhUTUNXIWk8bXxO32ZfPS9/4jpR0gQjtzS+m5+GgxuhqFxIzmaJ
nsRys1OUHaPBePlmiwXbbqxvAWWWI37waYAAgeAcz12/RgFfgtB/LF8DIrcO
6y7G+8kSxILGnPjOieUFKpRoKa/RwDSOyktcX57ucg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EbpNCX4h1BCgU0+Pl6ERtJLpeEQnOzMfmEbteEjoc+9lmkj64Q0aZOjhwXiB
S7v3BnWrbXSBLsx+yCgQoBl0vfjeyXOad9kB1ckQdDSkqlEbibMp2smReuKz
npYW7pUoVQ8c5NPQGxNPPF4tmzoUk8177UoIhjAWRLutvsZBGTaFzY/fjXqz
hIBsBSFL4fbHlYcCFCEdLh2DUKxiS+JWIfvhoJ6kaAS/Oqic1dy89wqqsxSt
oXfJwUfO1KRbcdBbUMjS8/bgz2wjvLzg55yt43M32LKpKstcSs28Krmfduye
Sxvw+KRoff5mVa8dDoe9LotjA+++z2XNwoVM3qTuaQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dM4LhX0kOeA3A5ku7m9jE7CGpNKgRVTIzyrzEmQDSVav2jHTaWRHeqQ9s/IV
vh6z0AVbPhWZT1tgJ/cB8zhv/HzJ+mRu3mxC3OR+zdWTuwXgck+yPIihLN0P
bddRBt21HppOMknJzi0yvrOfg0eIkIwZgL8MDLN+EFTNI3f+/cVMUfztFXUz
g0o32vUwfjm03lZ75Ju9uSHfLb8sfEcU526iVA+5inPOvypLJCy2mJiR8YFO
qz8eIm/sftE9foTY4Ag8S2v1g+zOAwLnUwuuTIOIP24GTwHGy3ehRa2L0FYX
LXBsbXBYdNcTzTEGjEI0FsjLRN57qBfnYrraiJyeqA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UR3QJQ8QKckiXI4s+DKnm3G4JB7tqqwMhGdZcD90WbIvreMIOfGoxcd46xUQ
suQPme1aX4WeRabymI+D/YrCUvmwOAYle2SGMo158sC/Y7WD5AesGtNyP6+G
GSJniHMzml3etzbaFU7gi5y3igX+k/xoWudiztw4ffJ9nCoxfyI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
OtLzVsJxLiYRWyoDB6IOk1/HMaRN14KHQ1/PwHobEf38lyq1YGK1UvANdUj3
mdxAF2hMS9rJ0LfaOvwHfGhFEEDZfEyh5AjNeuEVMv5OAwlYWXMfy80KiCPp
OZRT5bbsNd6tq+TD/Qbmn8Lv/W0CVBh8i/wBRHd1F2bGJEFZIMdQTLhdpJWm
k/J2ZFff11Ua0JrsiHtk3RDEmtEzXbTcM1YhgN063j25CzCZpj4QX7Pd8zB1
uVZyVDBsByCz1XPfF/eWJGgEpNnEVh4/yr4atYB4c6D5odUVq4FOu/jNnDzN
9aGVz1qL4DCvDQ2bUFcqkjOhk+1EOe8k/ZXJ0hvbTg3a1+G8oZgeWExV8LVw
caKMUeh4D4C943ALOna12RqIhp8ClUFgc535YzVI5p0WEjiJ9EmDYGfCaqQa
td3LoK+wVMjecI86J2BNqdGvguN9HMHI1Cz0DKnY490aII/642Cui1r+4xKR
9By6VWWqxsSRDvBY4xTC21W7ynKQAEbF


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mGqVG5Bi7/Y+gYoGlDNXTIjSmzWPFM4JCN4a1IoOJBe4M7JQT0/2xc5YaFkL
sWfhlGin4k895R9ku1ekbLE/zcc5QbzZnah3hW1M0fXfnMOKqPUZHTXObJSb
BfGpsKmSprZ7BOxBOS4yL3eDr/2XZytX5WXHYW1mpxVGforYIHs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
P6sjr0+r7C0d0d2SDCtNqL0jwXJpd0JB6iolhDp3EWgldZLV+t9fmuybH+EP
IuFDC/Fc+Tu/M9KAvp8dO2rNOa/5b9pzF20y+e4Nzlq4I2jh75wnVx7wsa5m
paBwHi/OF+Snuaz3c2s9MqpdzgpUlGs9w0/P3UhIeNI9B1kiqxI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1376)
`pragma protect data_block
E+gOidVJlhsjXoI9pe1lzmIi/RBcrk2hjc+hR9tauQTsOxxvSkoLEly0D1og
mRmgm0scLCedo8nZqQfTHfxLtUkD5BQ+mQZqPDwLhSHL0APeYI6ketAlbsq1
m5HBJ0BcaogKmuJCvZjwYMnoWWpAno2f9Z8/MqTS5zIdAE4fjcMrGiGDIext
gIkatgqThJAwduHTZsD7zSadm87tpo/GqPQqfkwQHuH3ZMGbjhLiWA5Vvcqg
pkfsctD+3mq9IJaLmb0OXFmwG+p8tB7F5cYiKJ3Jtsg77LA3EptLsxCtutWN
H+zqXoVgyG3lT1RFqaiRKmKurHGAu+6UL7aE4eUVOgXctuXBBDCv3xE6fVfw
472pf3eIk4KfL2k5ZmwpANjdGC3d7XkF9K++IbkYoysi5htFGgr9wZglbS2w
btlhNKJrPSHbjpP1y0rqyq7roj/6Y1JgieXFbWIJM1zx5pSBki1jvdz3XXKk
Rw8PLGZnUo9t9JObJk4iCWiHFRpqtS5OLkMME7aI1NFFexlYEvgGxvF3M0ql
EKg00+tg9uryyyHfqS+zViSPDoADWKEjmux1rJ93rNKIPI+536YVqVorY2G1
I8NzXWJglayjyDROyJC6RuKEbLQD1ng7u52Og6A5UtqJlYWxiX+risOIKCNt
h2CD5WZBu/LVGYP02jG8JQapBBRunfG3O9rCw+wEKZBnuaLzi5HOpSXo5vqj
Gbr7VAtCdnaucAML77jADtSf/jWlBZeinmyF/+FGAprNSDkJGqcR40/3MINg
JWbqGDlMC20Y+e/s8qDMK3+ZqMIm921dhROSIJYm9efeKAl1PxFdxmkqyofq
1xq34ekUrlqYrEvKUAXs9FSR1HB9RdDpxBKVOtdYMB3W+YZVJ7L49Mh/xLFg
cMb7EfneEvt875iEUMIGe/dMVoqnlVH25ogVtbCeXCQM5cHzSPtt9ePnmqHN
cScO8Ci7x+O3C6oWuXQWdzCF8gHWQ5T68zp9ikr8HS0riSlZYC405wI0k1l7
fap3oau7MIz7T4GueNSJTqeqyliNUnEARGKIRJ1dxjrM2ibcmzFdqKxXxYiC
xOze/shlZCdE8+kI8EFrBdjWm/bYZCO+Fkc7IQvBOmJcth2weP3W/L331aMx
XHfQlF465/HHYBBQa8pX4tE/SNUecNyejLgArV6iVwLfHpnrbXRu5Z9IRIRE
qcZ3Ma7gS4n7hIWvnju5A/8Owdd6IO0o22iy7iABeDwtDxFJn4bnRxuAMiUq
jymSsyfZsK5Lw15XMTqepONMv+zC38guW9UPRV/W72RpP6CCOzntXwo5zGrG
ZenmRUmUcnKD/VifVxPByauA1lzqiryCS0WmA4BAPrE6m3zYDVXKDPJLtaSg
/QuJIMXcxPAqFDV3YvU2C6jr2z5M9R1JpSplN0v1lELunW6GHWEaV45Dt0Iu
C7VwbW5TX9etQW/Z1Z+j9pwcLPr08WqMQn0oG9uwLXMDGFrQwSHtUAU9Vrxf
6rPPS2vmCGIu7XzrIazpnzSffTLxUdWqHEvmPHL1uZcKb2wnQIU64rfXD2Lw
N+frB7E33s70dElxaSFUlsWMov9E7DrfcOpDhiLxjC54e9GYJqft5g6MPn0j
mydYSx691k/5GbDh38WfBQj6z9jHG+Lna/kklWOkxHZuhRleX1+DZ5iSHSIz
Ip/uVhkY8boMabAzq6jzH+HBB4ZKbak49ddlHyFKH4uCyvzerfXUgdx6MsuD
2/N0UxmQhVLiwAWjMwbpCYnLcT58Ou3sKNE86ygCcD2KUOXvqVmecJpAd36k
kxF4ICxiGv6AveNnS5whfNyVvFbzotlL6Fs=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqfqeSjF3NMz1euhLNJUGPJkkWj+vce10XO17Aoq6wWjBDl+5itQY4isqPSSS0m87U8H4pXtnqxkfNro2StxZukSCJa0XobP6xF+JKQ7i1hor7FXYwnUBGhnB+/k3okFAzP6pWriKuNy8p0G2CEwKISQVI3AenY7kb4UG02Hg93IeeYjdfzOtmUdCS1/iDU1zYWH1npbSIsy/8xNo5b9bfZr5gQJRgSQ5YfhMXdQxf8ZF6pu/MfcFFgT40VsiamaEmwfc5YapJz1VUcXs7A1J899i8nTYxlyQwiCuqOPoZkVFAWBnWJVub4yF+nBgU0ifbnZWHOSWgrvYMJ864Vr8vVDD1ge3V7SpNQK8kAxkyX2O7IvdhsGYhmAXUcwu7AX/ludRmzxQ51NYj5MGlSqbtu6WF4SMNLmVGaRUvkb5ypeO1mNnu185vkH98diJUm/xZbEKxLwh0ipLSH7WCYidpjZj4gq575Q46Ggh3V0knICqPVYtil7A5a+QY0UIbgNH7FbmDSgdCmPHfQqOm2Bdvhi35tT3LfeHWg1TUDSGYS3Q7/nPHUiaS5jZ/jziI9Jquu1G2S8OFOHhEFdkY6b/foAHHzd+fc/8C76YKTG89/uGMBBXvjSjFzQ5Tfrj7oLM+3e9ejdMT2rttmm6y0eBg6CROG4p8FPE+UxFY2klsw9qB9WMraHKqS8GtCBbbCQZmcPPScaZNl22H41QX0SQbvm2BZjyQP8wHYbaaBfURrBq5RG/Rs+84TWYF8NSL/e1YR/6X7F5QfbwJWZLUpO07Mh"
`endif