// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
h6uKcb5Rnf5VfQOIACC0CJZY1ZvnaHf4cTaoKdJQOww+hEJiKmwmtTjg82Ey
RmbxXl1h8OWDjo+WaeSKuSw03aLAoE9rhcWc8GQ62eNKOzPdFzPjvZPfZH5N
SEpbzT9JvHg6To5LdXUFPBPwH5GtGgo3odJQpGg/bZ8+ipwR+0FAeSI4w5tA
4lArkXdWZagHNOno4znjWbwOvS0gXsFCmE2RLSp5Z90edSUhOzy0EecHc6zx
ShA0wcS0S+JYyXI1ok6BvRRYwtZ9mT54BRQiiG1N2oTzfxvXRrg37p/4hdBh
K6sJJH9zt0xJZdh6fI+PWG5gc7YGoAtSH6JBClZLrw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dW8QZg+EYBCJYNvDOAu0I/CnrZUf9oXtRTy5oPfr1x5lNM91TwEDCZAd6iir
p8W1e3ZUgWJbASNwtNj6i/zMtTGruYqb+AiMnO4g/x6PBmLcaaovOE2pjUXO
SlIweDgCT4v5KU8ZGUG8IHcEtf1uH7FMZV9K8FRbUpPWAZVREnZcLKDegygM
UTFTLJQ0Z6dyvZsUlKtO21OaLEf2khncoZcxzcySH5yryXT+KKepov1Wt9wW
RFnM4655E2nzm3u8yqe7BLpWqQjreVDq7H5biHXJsdK3uOevrSOplbWbjrQv
VP3GnJ4Vv3Myxk5/K5ZhFsYW3rm8fndaQLLCUF9GXQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
t5PNnUoTEgnfDdcnabDAbl3mtRkNPhqIK2N+KM3xiiBZhugzkV3wVoajs/8d
DG46Tx/9M7fIZuq/ID1gY2lP+5QnKea9xtKuesCWcAlX97+csQSfTSsuJGZA
h3HXw/OdZs5hF0Z9OL6alxmLyBMHKL7YsSloNuymcNuomCPZc7S2WRsFfb43
Kx7UGqHP6WB9HUk2f1zY+aToeGmIZgCB2fUVN2QT5WIgptPtwtdXdj2f+97/
DmKG/yCROCwsTNTkDKV2El2eCzM1uKaIzQ2WX0le3j80NjhdCqhSkYxOkyj7
XZ+sVHORXFqhtQ2E/kfiho2rJRUo6X5e+Rzh47610Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RDFQYw+GYc3njxK39Lbm9b0M+6GfkjhoDuO1uXnYqnRuAsSTJC8cOzyeEUdB
KtW0PBzlscS+C0+m4gF/o7pyZXbynnyrOSt9/mc31WaosGX7goCMPCtgXfGq
yHPpke2mUjsmzX3n6MV7fJTVb1qDjFCnk0CsvfqoFChKwQpskZc9Jq7D0FSx
g/Lv+qQp4P714d0iX5KvqQBzyOSNPmIcA8L0Jns1hZEyXF0vvO7+R/u400VL
ee0hJSy7gq+ZNiskWDafxAvO/9T6xLTuKNT6efX3IbLXCyGOcBXc+RrHpyNB
xQatXM+AoFwyBISEF6Psnqq8NKEUNJ6O1FoigzzbvQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KANqXEEW2Iw4bUprStvh+qL+xigdW8nQ4x/1cICcHzkjnjVLw49TUmxDpqKX
djlNOUswmX589zK8UI3bWFZ41vD/dBNNdkuzZta9v69Y/kvbutVaksxFHMf+
wXjzomQSY2PA/SLCmgwZnZryKEoc3ygy/IFEOXC+tl2MYGYFlMQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Ifgd0s6BhZZuJk2CEYEn3EiKqahF/JULtHaxvfBs0R667SFcFu2k8KyGaIy/
WgPW8LcuLcMPh4vR0/rQOMc2iZJAg7jQqICgbK2/66BhN+nLqk8hvhkGE5Xx
RAHx/z15oLFRmJURvZRrAFK2gwaMMr6g+y+nCMxNx0sv7DTTIfhZC0DRV4I4
otkeK7jN/GPuYDANPfoN0HPi4S4Y0vJW0syTJVDycyXGxq76BZIhGFzyksVI
hwvuXvlQ1OOXCGlTOzQppXgEalw/Y5KfVa1F5oZBq1IY7QfC+gNUS18gfq4q
BJ1ib4jEGJ+gXu3JtkqYOSWBu3WCvr1r1pk/SVHb2wVrG5xxTrXxZfWzvH6c
DFZFUWOAZmHQ02DirqvYIGm3gNkBJN13ryIdYK0RuP2HaYFV8wZzjL04R7MU
VPEICET3ysjsILFxaUiGAMNZ9QkqsEr1i8FOegsnKEGIh1Sj7S9Adg7ikjxS
iE7s1VnnK2YId6Kbefo8GI4GTxqGpNvq


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ruq4311hehjjaRQnQM0df3DfaHIXd2OWCp2FCJ2VmuVh9p4FdX9C1GKf/tbf
XKTkwespo9SQtgKXoD0QZ7wvoiw8DceNwtnHIhLVOPUoW/HbvWWrSWg4gRM7
cBhZi4bWA7MleA2GZn7tQs9i0UClwINzS8f1Z618SLP1H2Cu5Yg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NTJHSr7E2WKyHcUuFKSj1qgJsg7O2sIuLexRf+Qf6NyiDRiofzsN+CRSdW/z
ZcGbVhhPvIi2TfMRfB8ztZHGxtWsqYyjaInZCP04ecPS7lCdhCiotL+g8Jqe
yEIEmE6/UWbkq1rSTz0wXDtc+zgZGVvMr/zf9NBCSCVW8sCKbsA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 172208)
`pragma protect data_block
O3xgtPNPn2ROTuEvSkG9mo3fz/AweC+ZjPQ8Ejo5WHTwO1XZwk1JtQRVK7Vr
63WDv21CGlG79UkBOUk6RH9CWiJBrUpPRfOBgq8c5ZBuvDoGdN2h1yxw+jOY
ODTSK9e/fiUY53fRSvG0RqBjBnW2R3dfIdSYpKCWE52GNusI9RqY1Zu5s38B
NHqd0PV6FQwdgNlJeh3C5nFnr1rrLjkpouw2l7x00x6OkLOvdsemFXs6tuAM
C2v72IeVerFHJyQyhEJm9I0kWcwHqAv6fJLKoErIfiDFU2gSeAPolaKnlI6R
N6QCDc9KN8NSdjfpPsEkBkjKreBFz4MYHp6ONcRzkGnMm+zRQWY5QceJtCOY
V21/ht3nz8CG2yyUHh5/Onacie5rlLGzDm4nOVKA2i3T+wGT5v2DR3i8sAZJ
mimr1uKo4DRigKgYEAKZUQNWQlElEb1Ndow5sl034UevAxkUNE26AEqpZWdM
isgaokkud39xG85UivVkn7fo5oa78MrRw6KedXqAQHKZycTy/liAHEr4Ndym
edLFDwi+zPgUPU3jaBSBEk5sffNQsNqFJIcIgwCddHpS4RMa1CKni6DKMqX0
z+7vTA/AIaT8dUKpDhXILXhrUJRfYA0y5bplNqZoKquTNl0U9dWfa9JDanEq
amS6/TZCp8lfZPDZ5YnZqCzcGlLYbd0fYnaEca90akx2XjHJPBBl5UVB0T2I
/Tj5vWLtQLVwtZOqXeq1kb5lloJ0yreGHsk8as447y1pR1I16zd0+Z46Scew
Fkd3kBHcLCmwH7dykan9sf52OJ4FCGmn7D403hUWpkw7cTYywZsWtSxNJRjv
lxJptl7cYCXXBVhvVAZ5/BDYeHCpEdqP4tUTO9nrb5V5QIqezkf4ku4JlKFI
gXazdYxO5MpUj1mxiy2WBBiReRBA9jUEJvcgq4IY5YSp0xyVHlPzTjH/YFMv
6XaYkG8rI7qrd87gCXxXjst+arMF/VLkpmUYUSqPwp/o5sp5rpf40tRR5Akj
7CnUgciEVdO8o34MHlC9Fw9aJehU7xKx3NXjqMPjjMQhZrx08ILEBSZWHbxF
iEr831r27JV12PyvC1th1jyMhS9uiGgJqn77UgVgG8MSBseFTJxzR12Xf05a
mDLkn0IqedA1CSdUwJUGL7e2SrQ/Ewq+6LmEb9TuXtYuxdR1HcimO9vYIwSr
8mpXtbsrCUwtUzifq49l0p6U88UVKpicDIhnMI2XpSOkIcORAnyhtoWxgZUS
KbrmkqNNdMI6/EPW1IULMlJclBy8gu4uSTqvii+qtwrIsSxfiKJaeozm8q3r
lIQBwY+tHKutiTdt3jrRwP8g1lCKoZh58gS4EKokcuXfuYcqS+NKGZXX1ugt
6iSGKtfHNEvzdyE4NNaPfe9wmu0+cR/37dXUhuRBgN75/L2Qi5dwiAk4wOlg
lUKL+BeSKgXLOq9Yq9k+29d/KfbFxS38yvhkNHxKSFc13N3cLi0CFk2g1J7M
7RRvUP/HGKH1/dwDmKllPKIfLqu2+QbOFnjpSzPRfxh843miw77SkPmHhgRZ
tf9Jz/GBO/yAXrBphwrGpBWwC++MpJ6xQVhGduV19/epMhONjfPtr6YxY6KS
bSMleTpD/p3CUR+AnfCw9BNrZ72BvI+HHPLDYVuQQx/bh57PzUqWAUyrD2yQ
bQDZ7anx8XsxDEDBiN88Q6/eqoje1eR/iBaIDq7yi95WSi8d4TSDLDZn6erp
yj0oc3l3yNf2g7Vb54OuCzM6yX+ZJoAYWA98ybCLBFmmvv5InDzpm4CHwHrO
lwdhnIOfTbcqrMU97nZFb0xV6NQPR0PRAZKY5GZF+TNUGcjgbjY5eNM9eqMd
3JdMEI5u9OCPbudJzvX3PAaHoIj4PKQ0F/hDjw9oYIob6af/ec+9E+/oMdDw
Nzpntw5Hgl/v+YQmgTfJWifH7GA9uL3CNmqI4WYSsG0/01TN5ENZGGNMh4qT
LXNIW5ysVIknm+x06Bymc/FU9hRvFoTEdn9+XE9yQqvOt7pKDLt0oGAvNPQg
TEp7UmRiMKeKeA5LtUa9AgAZSLAod9GTLz3L9CUtjU49VPWJ5xDXVVJ4rnRW
3c6nhFmd0wSrfxqdpalX3+BsqqP4mAutGCg//jqMHHtlM8WTiQNjpxyCey5W
konQqKr3JQ7nQuQPLz3DZ51FdS807AznSxLEHdxFdqdfP4VO2K4KJAsbWY7V
O2SbUh+gbaSQHod/1T/cBQz4Ze8P6SRNoWjN2AqCgUBC8CAMihcJ9YcF5qWQ
TsoL18goLlj1czF+dMmko3rSyplIWdVPHBt8yLSdLmAGYxEtTvKEUGqH3G3C
XBFen03Y7pt3I9TlfQXaYAdHcOjaCAwLX92wj48ORwWrDWvud+JJeKXl2FOW
elTaEBOTAptK7Gz/lE4dfgAWm6x42+H7/fivMmggKICmcbD9oW6uyi6L8UNN
TNPqhOZQj7UWMnFitjMRoA3mFl5RqO6Y357cz3r6FcnufMb7QPF+QsNH+tUg
fxcMuB7hofqcPyYBt20NWNRFd/XNi2iwoJVlAUITpaIJg8SXMCMAfvpa+e72
+sRXc2l1BfBGQU3Y+TBezYLzgUuFylXSSH+Xiuv6Wb6QwxaGc86wUe8aX39h
nMq3cpiw1OmDdI6BkmidxyhwSq7Q4EbIqc3a6EDt52ZweoH65WV93T2cPf0U
4TB7ABZg7tQyTnFsKFsC93zIKQ1qNXqaonMQDDc4zsSkT36NEIaLCchia886
tyJZFDY3ZxTWj6rvTEGRM3zo2fxx9gSv198JrxowApWuazsnhtIeFNRDX4S6
pkCrnaPiR/OdAdUDvI8Q45xrmE7T1COtUKNGEesqS8u5dzJyzHFfXOg+EqBC
nChvmclRBXIbC9LYuBTu0y2idAx6xDpUXu0wFdhHyefxr0x3i9viqkfunKNQ
DQJIPD603MyEKDACjqELUqg1X8zZYiEbBL6AjsP4ZS06hjQSETQqnRKJuU3p
Ad0DjieVn0qP8nlB8qdr2BbVKcww0bZ6yNQdlHhhu80pEIKks+C7mz8wM2it
lwIG5jTx41L+Vjk1BpNXjVsuV7E10/oZmGVX11ibExVotYtMzeS2520O6/GI
eh/6roJlUu0y0BwnolslZ/6hvg4PqGssTieTcbtdh0EgEvs8/JYUmHqmchFZ
AOsBAzmUzC9+YC7NRWRijAn6aqcXziadCzJDTwETloq6mHCWqbQPM+McTZdE
Y1S2eopBZyqOq33ktpWmIx0AIyqz+ZFIcpJB5mIC9ec7NQtf6cEoTD4MPM+F
c5j7d6tSC/Wp1y+9BJ5FfnP+IqN0kweenKFGoGQmT2ZIPKo+p6cr5ahm4CF4
askMrK6LLJdTJ+sfqPtA0A+gxlUmdiuOKtTIvWpoM/0m1S8HCAQdik04Cg4n
iWAoqJSCFgp2KnCrWl2HNttVlosz8RWMQJbOULbS5fDlCGvhOgfBKttXBF6j
b7rpFWGjO3iKgm8VG89a+bFj+KJ8p4ndS4fWdqgG/BEw/GWLoqwQYoLO263d
59WAOM7i1DqUbxC+lEazWF+j72Lrlceg9LNAcv4QgRL/P07CIudOd/csK3C/
N6Kl3Jo6KZ9391bAO5gWakSOXgngp9+7JPhxGjMWhk/hvqYtkygix2ejH1rc
pcXJdHL7LPr2kAlyCpFTg/DgbnWnp9cdh1P6+Xudy7k2L15b3zL1xGgOXCuN
fkTXV2lbeTFCjpj4Mel07bj4foW9x5MP4st8wVzFga820VdqAVqsVgXzbZAU
3Vtfd7r2/7u5SjtuemedItL3Ay/Vkshmfk58wNNxKvDF6EDscXQ9nYrCd3z0
qeBWPJLgaiPANhU3fwcRqbbLUG0zZFR6MkbEnW7HeNAIP4l9BmNM/Q/WeoAt
ed9pfBz/9xGI4zie5Rdm+09BNVceNBXZy/nlIr+GDBEILNQfoXvF5/f9dG6k
DFjSaUddX0FtIAUn/DceqEP5AP2IPsYqG9ftDPsp4GoAQT/h21YGDz3WY1JO
kF17qoxiHe6EgZ+HLnEdhrY4g0uf+74AxpwkiBrV0YR39MINVUskpz5lKXYl
BLGl5bCXBD7LOZtkPnA4ipDz6qAuDxIWo7fnwIF9r3bx9u07Cq5Aan+hIxFa
hIjoQhXUarsmJlz43mjSsRA72GToyaLTOtpnppKFibepQG+FDmlpm99lLnG+
sJIbfJTiTP1sSwHNCgDBIaHC+U+k2i8/8hCt3pROS4YDnytfm5t/l9sNu2Dt
E08pMgWZJ2F3DulT0mkAWyItUZW5pJj1dXJxOD8Tu/66skYyq5AHHfaGyg+o
g7wTE5u3cEq4iKHqJftEyATWS842vZAZUsXKktgpIng0Udsjkb9UnFRVu7jn
kGkJJ1/mvL71wyHxKd5EjqaVeNc5m8r2bZfCDBN9Q7d/Rr/LO7XlIbfISUwf
ixE+qhc5YMYNzNzVwT12BkbxnHeYrwCc1qIW5SbXTTPMkrJtVsy0SvRxlV0U
yCNRcj9anNVFCoG/zSka7NDrNfaZXpZ7KIMrmpZJKaQVQ+ZIgU67RQ697kra
kUpdI5eiRzjDjCHGyOBDD2RTFaXyEJtlWKtLnmnMmh443mqUZ4quE5uLyPX2
ZtRR3WsyTCUmgLZYUh1rBNK1zyFmVnvhQ+1x3RlCsMntFjzMYWFt5LxiuyX0
tkIFmktogBk4V7IZXbLvdJRB/eAL93Gth14ML+2pFlDIkJFDU38YQJNISb6A
/pD5vEEp3vqbCxTv5OztcapyuIZhGdhKT/z3iuuN+t0+jxoRznNQHPmh0Hb4
HBZNKB2kkkqaNulnWuisQzLYeKsx/Lm9W7lt3oqHDCUG/X0szz9skBc06ks+
bhwXMmeNABSv/qH7SpPcvNj4qVjOYT3AtLrHRvfufK6pOPmJ75bby9FKrTpF
h48tx1tkVl2/aFInB+pP7T6WXgeU/ewaa4Tq1pxBCeECNiAj+I0YSDXYBvb1
ogmwzVSDxNLvbwxuFZQHOAA8wOjnZrzrDucU1UND4/4F4aPSc83bljt5jtL1
3qxYS3PC/dkAO6ev8PUcsZHg/wsklSFu2pYmB/tdEN3hWtDA5hJ6jkumpQdG
0wSWY2aooOA1bRpk+jiJ5j69US0QDkl9wfb1R0UwxwxXzc0b/1IL2LhE6vpf
1sag4IeW2PQQzeL+QWN0yb03Nwb+xzn4G8E40l2HkWcfiZV+hHUY/0ohWcc4
KZUpiROvyd0P3v5Pw6RgxvwrT6EytTTeFzgGLJDBPE3IhAnC9RSYfvOpEps4
5BVWBG+gK6Sv3tYiqptO6ngF45NEB7FEqm4IWiUlRSAVjM9QScOtnuhuzX35
s+p7/+MEIlo/ADMOo2q2YmBctJUeamqxR21Yn2Or0tAQUVj7l40Ecrq3JQop
Q3EAjctabtoL4S04qCEzPF8E7S7+Y5dHx1Re/bQczd3MjdtjDjhXdAikwvRZ
q3AvF0I0ODkbBJkoJKlvNyIkUrVBTH2PwzBtFa8/KBR6PfK1ICJuFP+03kK2
HYxYIt4XHJOUf1mExOzUOOYxOpB5s9KNcoLNP+a0tVLUTOpSb4l7Fg0CCNmA
3UkLQSMe65GPdwIW9rDKmyNeIcsA/jN5zJ2xCTs6Skt7KyhRd3pLvE1y7zOW
DfM2tqzPcgfpGItntqQ206YlnFuGdwEFxsUgmw1RLz4CCKKf2Sudy6PHT6rt
73HHtPII1P+D4BbfkfjVjnAkE/D0C7V5cso3OonIqSZfSOrxM0lTYzSFLiJU
4ie7XQCiWT9dm4sYPY6lPMcOgSuV+Y4ghRmXY0/8Ghr5Nd/+SdkQT7lS0FaB
rJ2sTOvbM6CUGGwlk/3Z0rBnO5NEso1l8lcSJcAuzscDTcXXKbPPg09GuY9o
4fdkELv3PhI3r76Q1rfp6Sy/rfJvQRy6ZwaQRJIdsz4Fi5D8zUoq3iiwhIO9
AC6i4Xc5rQhldRJUWOK/PBU0X4rS+N35Pw2EAUc7vXN+jqDAOxjaI3P1eCSR
ZljzNKdCEa9ygPp3Z3WZGv7ENgZ+hXh8PiUMzUpdGUJ+z+AIBZWppNBDaPmP
sJhHcK9RaFKvd1hLkbzk7ussWsc9P1u+VUjoU2pKeVS/V0ITcIfvdmsdwPW1
So+dURGiMT7iaj1iF9t2W9OStYKq8Te12wVIa3NY4jUTidUIt909aczLnWlb
bV7j9OfX1yxi79I0tLYerWU9dEIFqNg1P04w4oEosQoRBxpbBM3c2s9NPFC4
Hmtvk47HUjs8KG56z5ka5xQzO5uRcOOIfJij16py9eMHZAnI7bbv+Dvw8IaS
ibPTgGu44L2IfVTduNKSgykeFA1AXO/ps323xwOfSS6lLRbdY4sco/5Jifmk
zKsDwWqszP0MVWKGLWEVS4rEaG9LqGQdFvfgcbwIj8nptumTJQCRiEuAqF2u
Os8RTiyAI3t3nYFndfP+6jqZ8+Alfqcj10zq6DkKPEYGZShwJAfjU1updJ7M
YaHIznNi3ww/VgoqW+vX+lvBa5mew7BG0pGnemed8VHpSoOncWq+NSUuaFE/
P4SXwKVWH1uSbu0I61FzudmK19DjU+DWArEyTKQtsMLAuoaU6KZX/IygG8yI
5KjJwr6/4HzScvvIRHUEqm9VEiJ2uu22L2gAfQx/OWX1qqYQFzp/zBjTvpVq
X2kGzZtiVswxwHp301AB/bWRIT5uv6sLItl+5dx0XnveFNpv2uKvRDECleiy
H0cE/iPK8R8IR2Px4oJ4Ng9acTnLIKacC7jKxq16bLkqqllClBKfdWJigrBd
DC71Scth4vwnuOFGvwW9uy6dy+BrL+ntb7Wuqi5Wc3pHyY/SMB+HSYVcrRJN
+4YSE24NfEKhWuGkM1YlLIxi+4Q4vdd1AQwvDqPQAVZFOlSWenIC81Eh/9aH
QZ0YZTWOYOJU+ojEHbqekLOLu06W9WlfKDKgzpk6HcVwsamMndfXZFdHlD4D
pt2CJoJUyPPAXY4oOj4GlrgGqkwpQvn+UzkN4OyTyO10us8JRboWW85Xq06z
darT37FAgOSIygw1jO15rUqpDsnbR1VL6ploXYPrg7BF9Z6DgVZ5dZRP2qt+
8oQNhNIcQqUIJdzG1o4GM9ZObsH7j49BGc2Du86gd7TWwifoaN8Zyn9yVgHr
qJJOzZcH1eMd1E8gsB4Y+35+7hTfXg1eQGfYATexMoM8KG8slHSfNX4Q3W0/
2+laLEqLzivz5iFJCUUpYkO6trSKvUVDz9JhL2slxAXJppEMwnP8r09r9Dht
n8MK0sVrSZE28TVU1F4A9TyMkNw7s78+k/iGet7GBBc0lNf1wYal2QZDm8hz
MCq8JGLTbS4sQEK7S0Sw4XFJsh9Rd3DbFH2+F0CUYzPZ0yT3g52UGQV/F0EF
u7L7ZcwM4dzaUI9CGu7xUUMVTg9AGWzCWryF0N1dnrYm3nAxR7lh8b7LCGOu
lRjERWrX5ACDFLTYcIcAXb2PS8ZFvQZFHgE8cE1YmyWvoomlmhYH3UuYlFQQ
w3CBK0e9eXpjmD7WT3B6hO3vP/QcKXJHyXYM5BbU2WqJ8A1nRIxDTmPSYofG
Wxb6QULlOJeg5yUTMW90mQ+Ug2bCA91zACHJGJUsQFB9siQbWii26hb98Xg2
unR08H+Rctc2R36OZCEn5Lm9gg8O4/amXbYtk8thq8mIoLuzS8dQufmpzLPL
PcDhKZxxbw//cmKAQYI2DLNQOjvwlqOz5FguY2pPtt3/MMW4h/HWbmGICO6a
x+xwAXzfjy2bhIRRmcMRb70hCBc/uM1/AL03mBKYmtXbHu9MkFcagWWrypJV
4AWbnLP9WsRzlc5uH0Vx9vEHMljy6QSch/d1d9KCg3MFZSaZqhPdaYd6hRsR
A8x2bKYbF7n7mwmuXw25Nv+lcFc0rqhc/HsPezL8PPZ9mYidfPCLymrwGgWd
0wk8J3iVI1WEaWItBkAtwZVn9GCu73o812dwf/4pgW6DWNcRkori67kE1Tf2
wAigEIAvnsddQ79aUl0hCb94wRNpf5ZA0UlZu0XLdrozsUsEVX/ir0UyVToA
jl11DI3DPyFbhxMr8G4pAKCo6TGVLlUklnf2WoBMxl/BWuKPhbzWrcArXbPR
qVx0iCdTBeJ1b0SjoeOT4wVuP4jmOxtt5rQTkos2PoNP85LBvPhTiBjg8snB
xB/ifEEBgxzxbQjR99czkX2g3QF7wf8s/jHFmok8SAGN5TS2Q/OQ5HuDupag
EpO2YtOvUSCDSTfW0iQqcKwx4tgPgo1iDdb+6Z+FtFKA4C0bMD9zr2ZwPWSY
POtAQ+9zwohFywEnGr3tel5eHXDYT+5NdJ4v8yZuFVoqWjLeOY/Fak53Md2w
ea5b06H7dG55d+QlSzxusNIxBqfNDCyfI/yN0IxdHqU1cQdPUaCF6OxM0fSz
bQVYK7IpLJ+mzlUtVYpbFKhdJdy+bB8JY3roKVZC5DwQMcDhdPWnUM30yjxy
wVVKVjFh/UcIp/J2MM3pqUs9Bjkf87z7rmLLKQscIvPozpwamaww01e/psNG
naDCI6/5WNIQrnamQN2qLtu6oLPD576U1So8Nt37Mhc/QwQbXsF0Y90yYboR
Ly0DQQ0FluV50txc5k4acsjTQm+K6mbvelb9x47wYvYxzA1YJJPytdOb+2pS
hemSaIXvDRqYAE5awsbkSSBy5/ldYyZiaa5/oqDtdnTp5Mx1T4g8SuGAaPKi
QG4Rvcc98z94chEjgQogp2cbiWVPgc5RbCr9SFiOokqib5jRAjfBD+kuvGSL
nXj4seyaNUrArvHbZkJhBos3TU+LyGTDCs48A6n3vJ+2hyvSVKDRGNr7rHQL
1pHlsmbAKKPvJsSBDoXoBALMMyUPUnIWqhFYcOlzIm592YyHOoegL0fPdLCP
pKFizlu2HaAF/wWMHqJSywmJ1GhFPp9AjS+d2EDX757FakXLSJUX6dajWLp2
ldUUsYDnD5VUS44Mz3ncUGo8SFfsYAhvsAoqEsPSo8ScMjgQcDgg2ZKhVcFy
P1legV9vU6RvSt23NMhB857E/p5/F3qvCqXTdLVkVaftndTPtegfYztp5WZM
evy57t4H9XcgTr74cuzfiQsuFQYMr75XEVqjfYYFTW4dQxeDHPGy9QsXTU/y
JS6duX3NCW8y8ZNbQbUlbFH8k4v9PCPSswcK5iOfwa5VIluotSMmqU2tztcm
Imxi30ab2vNTyBedsbuPv5k8s06gl/9rmATEn+xDsQ3Y3EqM3eKrOVHVU3aV
0lLuz8v2+SteQ2ZhxCTRe6YtwC1Pe0Ay0zadvgGQqVBX9yfZP9XNt/pPzUwS
UuJQm/BKbHbLaWCJunqMMFkvvM/Xe5V3CY+KWG4vL/QBGBOOHwZ7wHZmzumU
jXkQ491cWC/ZX+FhO6kxp7FANS2KonZKGmUDkD3NldvnWk6BNSUghr6G1k8e
bQphkhSS7kZsesgtdqkeCjlH56mFB26DfcVNoCQlFryJka/Ywonva4GkJREU
8YZ98/bmPOsmaIWCemrKXVpSuIx4H4Va4rggKRUv/wXpYfn+uyMmQZ+EV2eN
RjVgO4xPO1A3uK6yICeAUXyj0X5pD4elNSjP7smldrPL7aQvhlXAGJkkcViK
982uBX2ZhwZuStV4pGGWTdwYamXnS/5UorYD199RYnBrlSrqfZQXMjt7F0jJ
D4IUnVqhC5UCwHivULGTHA6L2SEcrPZxVBHr31STxf3k8UwidrYIxQPC16IL
3IH1GbJYkunGaoUrT46z7OHonBoUrHT/qKk+7Rfhf/mWqhFyTMJ7jDmZqXr3
DvGUGoImsnJOXx/XCOpt15lBO7inpLLykwvICrN66Nwh71hpsv9rXso2DmxT
IXlQOs34g48f4Nb7lbh6le3hAyWlPnfgOg7nD/vY5NRT0Jsus/AcYPmu/1iu
UXi0B/Xpr6L2vRGkj01iSqgCJ9NdWv1EN8jUyUp836I+1HL1FS+iB50P/CBe
KtfS7mS5X27O9N23D7FzqAYLeSR/pMq7/WbmZiQnbmp42utyww3N+e10K5pX
XJP6tik5JpGx065N5uIn+DWUbNe7S/d7NMl0zeYwujpMH0q4oXfcVxYVjqIY
5UuNVdIFC/fHy2/Gf/VCCp1rAP4FOCryBbTlz1+Xyy+kUM1Hf8F4MXysQk8h
vmg21O03oC7SxgblXVkxNTEqvWunQkkywo4NauM1IP5LX3g8ucREm0eouz7b
I3s6bqczjVfOdTcdNZh9ai8uee6k6vMU9AJdAMcP9ghUmLxjCul++UCfGPlO
9i/5PuLb58LE/2xuzNOfLIKYFqtBVvRmKqDgrOk4d6Wn5PiaK2LSY0umd3t/
6I6g+gOuwdS8hVr2WA4uh4w7qsQiIQCs1qnsspaXsjCXXfL8HyAQNjUJzrvb
oOZTGkG4BJPmW/hVkqL4NDpN7w55d87+C4Rjv8QZMJIAtoZmwPJW33Do0Oz6
3TM1TjHzGDurueTGsUyl8jTVGDd3gmNQzYdvIGkdWrjdcMVKEZfHekgjMj/l
vEv21ZAo6VXqZTi17UBREjtFeDu5Vip5y6Zm65YElUjjxP48tcG4pFzFHtQD
f4J0rapm0XcILSabz8mx3eAIzeqhtuR2/Ck9+n8BUhmNhWBcmjdqLdPhr4zM
7xD+1Eek7bBT1bI5b9cjquwhvCmhbVL0tnx9idHH71sS+77jHY/Zx2nOa79i
lsgjH2fuM/rx1VWWbO4eGpSyWn8ZqOz9cMRr5CYOBtF12HJ6JLbGuKtGtNCQ
yPpwC0USm3ML59gjuF7Lzm6V9MIyXHD/tCvuyauXFZXiW1/646ZNW+g9g+ZN
M0X49fWPHkTm8ZlsOWXJs5OcCgrlyYgmPsnHJvtZ8V+ohdD0ITSak3XvHvHV
dZWRZp+qk+kzLlxyMg5A+tAXNOfxxjPyfTaGNCiHK91XxjRTV3PDo59NpOjM
p+/W1vjdOtdbX9hf3y7TBrb+KQhNBW/ju/3goH+Kltp3PUGo5wWXmBiMWwu5
FbCNXsSs3bFA5YBQ9eDtcdYOwss9J94dJPkGuIHBUQ+m2W3CL5FubJVPbHWi
WbiGTPOpn6wl3l3+VKroofgn5RMm1abdAowbjKnsNBVviKDP1Ndlh1wZpMCO
G4P4O/L3esZZKzbLJ/VcxopwxPJBr+J6jyo8i78Bc8WGDdAqIBAUFnUrJML2
3l4upiFWmpE8yFLnpF3B0b+puRdSx8sLKKz05VTQU7ze3HetIZlOhht5CAH2
S7mJBZMQk+fvNfqEdL1Moi+YfN4hm5TsCEHWNXqznkpN2PCttt520ktQzhuw
uakZtTJQSLXuA9U3I/O5pQned7ljHXNS/n4YbeYSip8MX0kzCLzqJMj6jRIw
RVfuCJkhtXVzGyl0Pey8OA7TFTIx3tBDWdUHT8SZvxSuupKh96a+SU3B/Yg5
6z5CeSI0/uUEgB1OaRpwQ4DB1YAwAskF+ujsvbqljKMxqrJAOXJ8jrP5/TyG
fo9d+8HC4a51gJNhDW+3N+70D8bzqhoTwNv3Y4EbB3Df6HY54GtxPOUHj01b
Wy0NYu2pZRtJp3hpC8hE1GzVXSLaCuFvrH7g7pmdS6wZTcsCNDmZ8Ke/OTvS
1RwRRYu5MeUDfQYgqT1bHnWGNgAm4aSUyIiYJESAhN15ZXW9V8r7PDN6NagP
Kghv3pLbmsy6UXB/fLWxHMi3Gbn4VMfVQ0QvdzBdgr9wdJF4FoJK16c8jVj4
5iv/vwEZ0rm5cWMWf1T+VuwsWtJMR+tAkf7kvs5jzsOwUoz4e8cDSzuWpio3
LhVvWVHefSg6r/hZMTsI8uduAxBMwFye9IGgjcnVSAZFajyXeTDg9UBvDYpD
ul3nZDqJHRISijslD75zsyGiFkQDv9VX9RldsKfvsKJ5QajS2ByG/ElGYuJt
RRzR3550cYBWy6jBhrr8LBUoDKXKavpFJo+mmaocm9TTX9IDF8FPOkcNrlup
eTAHVch1rJY6qS/zzoySTLLpSMMfwC3Qpfb0R9mSzKdYgaGwTW/mAtG0k8G4
VVBthnNceQWqz0oJkRjkHn+PJ+kDbmWf6ajQDA2iKmD2iZX4nkMDxceltSRi
ISGIO9yCKQL/b3wN8Cuke7JphCbm3N7xQrllPD5VtO9BS+ogU/c6WXv6h9JC
mis8IyXYAEMPqKsltvd4UMMNzKEVKnlkPfoH5/Z2x7VyqbFiLTgYy7RI8iax
1bbiONapElNu6LvVJO6W477LIXfE0LOakPbPwn50M5WL/c01e1fsh4uCBRWC
9EjSN3GJEXwQx+2ei4tMBcBdd/X5bSNuwIJHnT+77u32Qudevb08ZrWGb2P7
py1tvOFM3H0X9PIWR8Gb6LP60Z5TuRBlCyGG2beoIeovwuhfYqNG17uIW509
WiR4yzqaRYNzD2Gv20MNXfZ9HQ2mhk4q3fHzSebvlqp9/aKWc6EghkPfFfKS
mL+ZJDR4YR3oAz0gjPZwjyu3wju85ULCZVwBWIceB1s8NaYdy3AF/njVdZaE
s6AcHhHwbzEhBNHfcPELCKbRA6HVuAoEIr9ty1xmLWiDcjFm3lMRecS8r5+/
CuOVQlDTXj7lU52/xZ4+uvcpEoV4E1eE6NHU24N4Pkh9LaTjxUoFexFN8sbx
b0/xWrMWxcPfFdtgeOBuNliXZE4kauZwPRumUKJpZgIyb7PDTs3xnBWEICzQ
hDuEio3dCwYzTylhNra+OnZlVOTs4W9K5X7n7zgxa2WNuliBtRjHUpwCwnCV
l/EYPOSFd3giYk1AardQJVbjk1wHIHnvyiOIbtv6I/NGCe8UNRgZzXc9k3Bg
8AIokGrfqfuoJWORMCMwMh2hpeP5wP7GbDZ6trwJp0UMO5U69vWA+Et0NSYc
UaENFYn2RzzGNH574rcSaZT8vWYiztJ8piEuFo+drz+oee6V9k8thf9+MZkB
byHj0ZkA0oNRTu4I/LtQL7hy7xVQ6AmkseJACJxK2uHy6lsVuAFAXV/07YcZ
KOTIFR3h7gdOIEPjaayHbzAy4UkyNQ45GQAHv7aHCccRm4wG6Jd2YbOMj5VS
XJ7cc/oeSti2ck3kWf3PZvUXMH0TJNGQCxJfmceV5PZIS0xdKvxmK+WB5Hwe
4NBwRllpn7l9MsA4rJQ8t0FHblWF/vrSK1fhEeSlRu+71i62iEqi37im2XCj
SqyHbFKRV47fqSyc0Zu8krl2b0miHo61ryH8xL7KLH4Mkj5J5rBV6Hcoj5Rm
V86Cu+/pmHroBrYmfRGKrb+gGawyxAKArlA+YSLNhVsR/77lUok4o4Hthgv1
QKbvyUdSJnTCxVHDq54ZUvHBSgeSKz8h3tQ1yyLsPdH/nkQGj8Zo15Ous5Es
F3cg8omm/dot1rQzIutJH/lRulvd3+y8GRTVnyNA3WqkjMCcUxvao8aP18nU
SPlzctO3cfpLnLZ5KxLw0suEh6KBcIaQLl5ltWeLKdya8fGHLjeQhciPi3CW
DvKcn3ASSRG0dsqznDmoj6oSqTPTpEqcvNzBUyrTpu9nhJIC4+DXRs4czdA5
bBHDHEw5743RaRFqhr0GFuXP6TmPcBv/DTXeQb5REc+qNK9MbrIfuqkr2jTx
LzVBWaoGSc3v6E8WYZBa0OjtDgjqu1gez/tDQOlzKslO85ajrKVhjZ7q0J19
nUooDCXBP09Bbx6GBrkimZchO61oMcl8EMawI4vbmTaoseDo/8gOZ76fq/vm
5DclLWurm/OrH77QUsXW9oI5SgsgiLjLcUZLhwSt75t2+Ua+3iC8/O9kAeZ6
iSkoibIvbqUNp2LOoRWe4CcJG4pSF4vQt2ibMkgWERvoVSszNT2r2HioEjo+
TkfvmEv2j5BzlgNpXuRZR+3ToAdDT5pEKT4W7B91ER53xkrH3bXlscNjQPVX
zjVoC5RmzqfIQ3keTVicKXEeV5Y9dwtK1JmRs76lGK0F22HkKPJQHjBSbw5J
1YzqQ/nr5pCxvdyCgIB/NbY8qcCWgajzNqQEzfDS/dUA3qjEC283nIWMJuX5
vPpAIuyyNxyRSgGux5FqWsAK4cZgULWeEq4hltkstMx4/IJRcv8IRm4BX34q
XiGolV372g+lSMkqxhEpkMbC7GJF+rOttGvA+w5OSXuGpK+EyvHKnOKv3rGM
1FAr3OCM6D00LY5IgMIkgf/y5R0u819sAhcWHmnMYg4lSLiYSRl0g3K56spr
ExoysnW43wS8YNmOMZKLFuGjEhkj+eGvhkksBYIUCOuSdDundSnbyC6W/FCN
FGzXtGZ3GcnrEo72HijnGTAnS3Z7Rf6LDOABapSEZwa7naIqacNWU0vdRgEl
5ZF8lDf4NB1b4JlZrPIQf5N53T8vbH2d8IlFLjCJRJK9QwytKQM6l0O6sQd1
Y8/ILgY/gooUjnMKIUyRF6U47JpMatDwAmRLAUUNpjn+nSHo/5Bqf1e9vf9B
ytpvlO8vI4wl5kxIwCjzRRY37abG0wLJA+/ay+1129NEs198cMedRjSc3GgV
lJGhzbhPwZZ4cQZSTgHflGi2SIKcqyuXfTEjQcaJauc5r6JIUCQ3jUJzqGzm
i9TaK7cS5t5kObM2tl8+wiZ18nWY5ITAaHggQKHN3O2pJVuAQC/gVZ88MQiX
SfmWJu3IOYswwuFFG7bDiHw5YwrEP9neQliM3/ZLIebK3vVMGTcYaF8ZB6vX
I7K5aORA9CwvrCj147N7QBsTxtLFwWMXeAhAlRjJLXc6na5ukOt5NhphdVGq
/MaDlJUN2fN8D5yVtUQWrnOXcCAqEJLX5dIaO3lVm6tjtDQlF+3NdzdlXMA9
bmcS4aHJaVH8COiHq7h98S5S0VG9ROqtqxf9CxOFC5KYsZl0c2LkO41YH6qP
GASBgYT6YzL/6bgBgn94TDtMwZxP7UoCpWrRwnUu8+SmVAHjEMvgD2NaOCiB
M8W1rC02fpam5SchT2wBCgGHx2UfZ/2JmkywJfrOWcOA1KeNQUt4PPxFk0ip
WFfKi/0mWHSP4zpGYbzuD9rmdwZG9Ik9dx6Pt8OHYyUuXtTGUNdTPg/wEFy3
QUfWRAA8PJ47dTjcaqtAOrprPtaPF5aKkFEKf2vhNLoWxZ8ILa8Vo8al8Coc
6sHbWHpsfDNZGsJxEQmhxukECMANSin0vUYzy62kA07xS1GdyfDzzPEiXond
rfAaBJhRsfHDJ20vmZ15eeViH+89Ms2jXgTV6b4y8ezb05oFe8TSeYgraaoA
ntqBXZWOC6k8y6agy+pbhb2LVXtpS42IduLL4SSotUQpXDliam9qTGwjGRgk
a/K4P3nR73/ACA1UP4EhHhNiV1MPGGvaq10HhLa9iDltYEaqDR5ImPZHCy9Z
QdrYItDq6n8fNsxcutDKAJRTji84rXS6hYbm4fFwZMSQMAKWHqNlqrhIJmIe
6BUeX062Ih+6NKhS4a9gRZdRMjwfbGb+/d2CtDZCyhBaa2ZUjgeONnWrf1M7
WAc8/MraMzohhJy2j3GKrgpAX0wHQTTyqw+LuR1jPbBkxv4ot+07vApmygo5
3yeBt1knMsTGpk4vtnZMJn8LsS2REsvV77wG9JAbmy4BHusYH3ynW45E5g8/
AXZOryk9UK9rROaz16lm7y06n7EyaVQoOYXmiARQC7iX6JtqyJppnUAznFDJ
EimQ7rekRgeR7+pWLj+D0IpuVh0r6G7+tNSUp6gQoUeJp3SBXPkCLiYABjd5
l9KigmMk+wbqC746LQZPxMxCOvfNBi3JBgqz2aWBwmtDIwfOw+Epy20AY2Jj
eaS9TnHQ/lwj2Dd+aYM1P5k5zCTh9v/fEpM9763LFk5gP68bnkfe48usITWM
1zXixVkDSga97NhVedRzYt41AsVjaBCvvBMKYOaP40BmIWi7qDu/5YxwrzGw
42x+o64Rqar1SkMWsgcocUXGpJaKQSVCKt4VOKXCFD8AWpW1X7AyQD44tmdc
Vejyyoh3pyHJ9lN3WoAjatEkhcr1ityXuvDv+0fU5dVft9bobcVjIbbwyktO
ly6kVwYnAOn0VBSo8p9eofAnIaCwyZIhzlxKvFbbFYMH+1OEJzL5TO24fnWj
cVW1lnV3KjIcLgMIf7ArAMKfcEEmmIZ6DmXJUJ9zE1rYnMNer6Ari6iLOCuH
ACqDemdcyn3bq860oT1VTlMspKCcHFLeb/BAkgd6xvDpWNAQP8VnZfJNkbQp
juEOcISKRQbO2SopkSnsKs/YXSQ1gP0hEJ2STN4EId19re1NbPZ00k9+yFCC
OqQ+cMFRrxbxt/41N2j9mou1Zl6tQqH0VT/3orAOy/Mu8wc68cAb/bV+uT+1
w98bVqDlzvwHtR/rq6McVPlr9PiW1GgtcZqolBQkbkzuBlrdUwbKAfDiL27s
HwLVSI42vQNx1Gfn1SxGcrjWwWcdZB9ojdjN8PWzXTgE92WJdR8dQPbsHCT0
HKDJWsOhp8msbSGsFifJqrakwlvUJ8edWXJtlzXqXEN+n9hTRx7HKVhDUWZI
d0CZRY/PxNR4Okr71S6Hrg3BSuniVWoG3RtiwbKtNwCwI3sSyYPZMN9fzs7R
tSlI16ipfbvpxXp1LEEbFSQmjeyQwQgo+s2CmrddCPV/Q8FIP+FdGKUjYdbW
L9X3bElGODG/VwkydTl77M2d/dyUDgcicDRWJrdQo5W8XvJK3dMbfQ4kDGuK
csu0u+CRK+J6ziHN7dXec2RAgME38cgSHVnhcmZqVjTH7e07UH+oSfDevZf1
jSNtSr4F+KrBhvdKiIgHVKPMKNIr1fz/Bjgpid+GzLZwd4XXPDQw5AdSpKuM
osjqxK/1WnHeM5hPfsBzjQahPe1v0mGNiqYRjS6xWG767o7IoEVJQEAIw1uC
P+hKWIjfLujqEvEczBgTUusiDPZPmlv02QUhc/VoE7J20ai89rsZzEjjLk+o
qTlqQKh16yK5qaAeMIvIl/Dwzf8RZ99I2rlHb0JoUXC0cNIiCPHTin6jd4Bs
8WHzy27KmgXO50ao7sfMdvZCWz6RhBLdvjM3N0X7PaGiYYwCx5kxShEZ/L5L
J11zwFnlreS7zs4YJn7kU0qKcwu3g5x2UDw+7R33Z4EZc5JoQNdzb+5virc5
7OACEeLGH6b7gvrBJQx+r8bBmm5l8Vql7X6ulIM4ZhUCzxSabMrsZpbeD8Bm
tGconcZv8jpJjakXRXnOSJCREi7/+lTgDchOF/p3mkMxj7UhQMrs5ljQ7Ju8
9theJM2GHjSGr1bYyLIq0EiAX4QVFDzYFrchrtGMxxJPoyVJYyVfw2SdaDOv
kgi23N3q1rEDIxekevrYWuR0MZKKB4CFTo9Ic9fqZNZ8R7Gy4sgn7+JAKmAt
m/EQN776bMmDPpqAi0sRIeQzHpKywSLEEDUae0PtaHLZjGbbNpqK8te6Vat3
yvyh8pIEK5F7JVx9Sa4Y04iZ/MQTOE8J/5VJDqAcPFIw31U3Cuj3Usz46TjN
DfnpWJ1f7FJBYw0SGml//jJCDaHKzjigo8SWWqCbZK76koTYLXUm7bA53GC6
G/KcbUsDRZ3Eg/1WMUwZ99mBegMFcM2uoC0v+lzWWv/nN/3qeK5LDf/EK5xq
Q1NVVidAHk4kE9/yJaPelT6nuDKYgw27X4Kyure4OUcWLMxNRf5rQjIQcItW
5NYuY5M//QsH+mOqDKD+Ld+cUGd5j0f+1Am+YSBjyXw1FOn0FlBSITunxGXj
cCK5QuO1CsB9eRcEjf4Je7sssgYu9aMBxoozRQEs1ONEpwtGDT6zjvq3ab2x
xeSTNOd39pulyzVHv4TjAXyONKJu/FrOl7/4xopTB//zgLYMCG9HUJ8heeDv
VgkPJCvRlWT0GDUkwuNh1li/nWTYqp1P2kswzKRaI9zl5cYUV+vstF5EfgTs
LGf3of+fOx7PW7E/ELpEVKSFC17xAo7CPQdGDUVZdHnJJpXwLEq1xBlqzyvG
IPuzYrHuPTlNvjKdtQ3dV0FVb25kbX9p6jsjGaoTKDgIEGGzOrrayGNi7q1M
tkZS82XoJHcEU83A6HCEg7a85htjf57VD3rMKQVbnJ9s9k9jowXEOWWUMLbZ
wmslKM6R32VScpsEQlVLiej8Rake7fUuIVGyg2T970VZOk9OW9BEW0S1XxEP
U3J+X1o64nRbjR5mMeTQvnn3bUnO9Ge0XbNssQcfVomQTLteTPG9FUxRmV7l
s91vN/EUIHFROkRIys27sCoqKuIGzzHN1ubDIsFEsH4NvS7/z6AzXu9bvXs3
eAxIjUmFGyxkkQt5fo4W9LqT4hyVX46wQnlF+9P3hvJWLXNZXy4x+qMM/eMN
2i2/EkJJo77w75Yx9y3nqHR0+C3jQugADoeriZXdUq5W7PNdbgf9atbQ6BLJ
lB86kNEmcMEbknMKhcjpyHRxWZGfroPB4eujwy9km4hLWkiSq+IpnugkNZHH
0fFhZh0YaDAdKDf6Rp7Ch+F23nu4Pa2RRGsBrsJePGVgCfsVaUXl5xaZo1Az
F0pD2dFfSmy5FzHw0peOHL70AS+MzDW0oOdNW7WCGcObd9MtzQ2JE49JK9MK
S/C91TJwIFCIQWCoSHtwN4z7BGCL/F6VQ+04oBw+xEe2g225hiHkjPdC99qY
0bUaYjYP5qpuiDeHd7akZbT/0mej6bkqhL4kW0yd+90yZV+3sS9hmtNCGvlf
DHeckrBgAcZDRma21ViGLZRNmH/E0HKkE11U0xhrSR9w87TR4KFlud3oqh2w
e+JftU5lVv2UfT+NGRAT9xXA4DzCgTqKuCBphoN+4P/3tLwRg7UP4anfRQ5Q
xwBwd9tlatctYpAn4K9SL+QmImLTLXggg+KNqmxJh/e0cs+Hv77CMUIq+Kbg
hFBcCWOuKA7SdlLBXuG++A6wIpkykiF4TRj/HfsLoUbpDr8o/T4zX1nm9V4U
6/hKhB+Or865D8+qVgsREqCZSfPZLnB6L+mwEfBDH68CUWIpctN4V9clRBs7
NCD8bATPn8NKS/3gHHxizwDaAA1dHNu3RbWjaMnHjYDObFWvI+gdG+WA9JGC
GOHM0v9eAdvH8OMqjOlNRMcj2/5zHkdtsdzJMHgRxlq4Paj7dH2HOIp6HpYQ
Mgf0TD15WPGYHsLDSio3IBP8xOMEMWMCdJbqwSylbUf4GFHTQXk/3KQh+lZq
MRtZGYgyrwAV5ZUyS02/VuQBi7o9zSVqTMarL/KNquCbRALcO4kiVj/Mha2b
VX7m3ned+uoz/IVI2KiqIUFsWAYkhgzKy0twjk4bBOcfKm5WKxHFuA2wquIq
+Z5EydmmArIrCeWq58aoMlIiF226IDw9srZaeuqWGTa8t6ue4OQ4Bq5xydp1
ek0Lqwlfkuyh/wZG5usU81c5xli104mbQUe5NZfZRD54I+7FyhT6i7r4HTFX
M+LpwAuyr2i+d70L1tLA73bNauXTJmldudHhdpK9d3gAmGrMUYUtiRn4EVGH
wz6y1ecFCpJ1yKktzRARBRQgNc3GC76vuJOSb9JeYct3QFr1rHi96dLgXPHY
x7fHqXaQRdq13hNl2AZhm7eAbd7+8mt/5Z1sS0T/+7sZGljHrqapGd7zl0Hh
uOQbaVzhaINSVKDmEfMzuZhhIzb6G4yfS2Tkhc/QzFMUwyA9JVo6rRIvy/Zx
WNcbEYda5Jg26J+BSixRPHUVHH+0/P9QRtR9eWS3jUjxQeHnjJ6YErQsWSrf
9vxtrOBtVvIpBtyHLEnZJqoXJxcEECpI7TDoQsqyr0a3gBl5OUWpFfnfGySX
hiPneBHtU6FaestwCx/MdXFxOgL/AT1UhDwGw5uohjbqzIT4x2LWgl8NYVkT
e+yZtroKPA8tGGLPqBjkouJ0Zcmb09qSr0NUPx4Ti/oloO4qR5C76gsdkSRY
B18kfItgDR5Dygl7imIHUvgHcnzzN4sUHU7SentWiyBFdpxRDyUagDctsz+8
ZNMNkBBZRgJ/EIkKGHrPWO8J0LAFP+dKjyjybnkvUOMl2RkOtZUmCIUD2f2F
mWso5mZ4cCS2T/7o+UznvowVUc+6qEwPk1BVQ+GwXZTYTy/3OAbj5j91eoji
vMHnGy5+EyQRXX1Ahxrytn6tIwIl555iXnUofd/L1wwldHwS/SBHYB7Tq5r9
H0g9XbRk6xrrhojoVle5NbdNWVxkog7TyR5wyandSCfLZSIFnH9otaYdBBM3
Yz+drAnI3Bg/D6muAfZWxVMCoyh2x82+aJ2ZgPm+G2iN9PJ74kp8iyR/knlI
Nl2hZT5VdA7IC9AA7oVmkPt5kSolxQNI/lRpxygzv5qmGEtX0oGrlDZ9qL7D
TJCvUjkquyQU3WA+yURrzW6dfFTk600/s7VGSjuWCWxxfVZ+VDiIiG9mDNHm
WeFeL93LT72vWnX5D97snXMIBMGRt8/Fa0OZRYTen2+WJ1gjrbJSbrWUGYIw
sCVR6vVYLdYQO6KPR9K4XilVhpO0CtKrUxW4ThD9Y4CbeSUabXShy8TvND5J
3ogU5TvHMZF5mhNZfiGMJW+HwPdQsgnrQ/mrYTfqdLlwfUeqg62cQXUn+yRQ
K+uYKbt6YG/KXl/ny8THfCJGIVSNuor3DfwJQR8931EEu5loUoQywIkWkUzR
0p1H4Eds4JQx0qYl85khzbpNtR1mL3zKiAvBQiB7flSNDbYTASxwc4815sYl
hySHoDfPsqf4nHFvWrjvqcOMdlmfKdpbOPDGWtFZVPopbn7GgtAubqXkhgrQ
iYpE89NSMg/1Hr2G73D7gLja+YR+UULmCT9FaB1ahjjL+l2cz3r2/ddVRCxX
LVaNWEFUhrgJHN9gAuJsaT3tytCjcRLy4J9iDVaKe7pmrozc9ODo0eZd33yJ
14w7g5uKKkKSOYREAyepaxEZIQBQu7hqF6BIhOeLgwMM+XoBu+X1Ahle12CE
IirTV0UZBjkELfXc31PJyNZjjOVf4cmCvm1CKyx+mXxW1y4HC972/OayFlzz
KnNxY16+9+mF1Y20rSYjhi6FpSFC03HsMGwa/QjzEqnzTSYllpvge517oWLT
BqhxZS+krX4N6lyklZudi11FFwCRZrx5t1GaXpuASw4QMcdddfnE2ckFN8gZ
61Uczzh6KmxyghlN2OiZ9mxkK/TBL+TnFaRxciQITXVpoDNCWQ0PmBH7T/pO
BMfYu8su0U+k+EDvM5Vhac1b0TolYO8h5ixDnqVDP/ZUgcpxrtYOqiklaN+2
Katxlkm9D24jIuWTO/M9yCT5Z66PoGDxDfNI7J8MQ2maWjoVxmuIlkarazLp
v7QLb1Y5VeSB64nDGF7GGOgWkYxff2V1xaTi9m+xr8sAIeIpKosDt4ANC8dZ
9N/LjleVRDOPf+E0jmrcOCEl+LRLcCLVcVcgW5KOh/mlDA52qy/dRYNw0Kl+
jyeEowg/LMKopbYRGOsPD6aIGr4A95dJWGzIJA7TQs3Vc+pVQU9vvTOMN5Pz
brMmK7fQPtR1zdBW1pZAPHI5EDK40hiHibYR6ZOpzc4F9tkRQ8hMIx0CXVxu
ahD7AStALlK7EQ5Zh75GUpCZdEKMSaOSWTO7fzbGH39meOQxcYTFLSHmPJMt
UJvdJjbKoUI45mYRq9VMK6YdTpnnR8TaYSSN7M4rP8E8qeg5sE2RUEqiLXyO
0YgZ1e/59lZq74riUxdwxYq6k8EOw0aCsb4EGfsKuylD7uL8O2QgmxsdFzPh
0j/OsyxaAoMCUbxCAIEXl85Z7D8llPbV5FI17s9lYdUlOisS0XDwfdTfsZJ0
DLaqlK+VqzB7j0swpolvCNOjzDxqIMwbAqTLPGLWNUBoFjr3ltY4rJqNXSc+
QvepFiF3TL/5bfV5rUUuiENqPnYXNia1XBWAcckFjQo4Vns6LEUOQsJDzT49
zmPdeNZEhGAKgJuBFmkBV4R3FWHERyTtLF2sQH4fluPbvYxiih7zuWMjGLRH
5crgZQwy/2oJThB70WaBuVpJfxQvOdXuK9JUhpv+ZTbhmW8ToM5NpGKM2Ebo
mEaw/3mFcp1bYbVjfcX3QP8rCFeBKZ213lXeeeqiy/AdS1GHFUolqAm50Qaf
iA2tOe8wmgkIE3sSLvuK65R7W4yO/o+r8VwexESpDQhn6kc1Dcrg0ksef3NE
T6MCgCK3jyNbiA+yo3Ath1RHQqvwryglMwbwReuLwtiOSvlo5yCkGb+jNNFR
RUz9qg6BpEyAgu03oO8RgqzxJqrn5nXfkRX7Df+nr/vZUyyN/ajinpkH3qaV
uz6U1bda9JC6WLiR5rUN7zv2HEtiKR7RY5KCLKCtp2XMhFLJuSOmSMD2/blr
sta40Z/lfIGhnwE0HaHs0RC3Xdosmdb9Z0c0++iTsEx6fziF+SPgKMsfxRsn
8lbbM6r4d1u2wQdW3Dr9OlHL2g7jF2T+fKwd8qxzDy/MelP+f2LPH8x8yUrI
4QTGvDkDlicFpz6g0y3GUo/ykh76mUhmXE55FdX8lAlz/xd36jR8q37QaxTu
bfnTTf5n+4OXx9qkK2c2LoO5V9Wu1BvbBPOLPEWqsBc6042snuZMLoIVZ+iQ
Nlor3p5p8eX2UoV1uFcrgBbnSD18EJddYEJmaBv5tlVXfimR9Ck2pffeMovS
91rWGhn+n8oRyf+EV2JVNvQJtiWXzj5dsbWW+AfGmxSrHBAyxawoFxxUbvJR
cJAeMZaqlPkg5SBDu5BDdCQJgAFlZ39idPDLHwW5xeVvD1plj2VTUNJwXm9M
SMNEefmGymefJiJFfNigLu9u4UH32c2d1hexg2tN+WkLPW4jUMrvBokRoqdn
SDRD2K6kPQm4qoMxm+ZNBCkmehuk5Xn7AHG8Bgbdlue1BgSzPhYAQBtzVAhf
H3Ug0d7MwPXgGzGq1N0wJQBRy3cwh8jm6Jp+ZTl/lU5udqI6cT3x0W/vs6Oo
4//OX0CPtprZEPhFsyUD4FX0vNwHnRcX7zlOzQSXCkCa4zS6DZdKFuVOSJj8
dzwKS8+TVPyexiIPpXwaVftmyqQFwXBS/JA2VDVAIg8vCPUf6iIW0MfFFCcN
RqnjYtY0A2B8xmbfyiYnmUvm2AOnxa6D+ZHWOCgQW8ef4fSVECEInlSfaHws
Oj3crMThHnWULGgG08ahYLOycTGTv1gvDVG/ozPwthU1ZSz6dgmz6AIxEUau
IAgfSsAjcupWHtS0FupeKLKxH/Onv6ljaK+RMrtsOiUIp+wztDAX9pvy32A8
mBBK0GSM1nMAcwW9r1+nU4Kk7h/H6L+pzylCMEuOu6XdGkuQxPHqQub6HHIX
ZRAcX4Sbbs4Z/B7hciD+I8uEKflMzA/Y32xVABOUZnp6qdBcwohaNtJnuuMJ
KG6AFnZ18yFVBX+B+OPsdrUeursikgqDFg6cWXAFPge/rvdNE1sXtL+Cu8vm
XQd/++0pw1xIDPHbnIc2BvspJ2nrT66seTzo3BNptntNbr5WkJlLnR07lJzL
aS1ndGpvdbsthFLBl132Vc1kTZpg/H2rdxkZmUzxiY/ka/EyFmMQYhY+6Hwi
iB3VxXBnZ1zxLbNYsLr0ukhQWHBvlRhLM50QuV/e2+kUs2xUIOEaoc0xTsZo
FST8fqncTiHIeiNkWCvEaFaWRTOncmekllWG3ItHgrq3lN0mhdHU/DANG1Zi
8U0ka/QxprEZeNKkc498Xzr/qVFjiWvq5pFnpu2PoCQwywFvAtKXN++feF0c
2m5dKrBgbQgald0CMn2rGg8zszQYp20TfeOmQuth+6ozaBjr7raz9kIVoyhs
eHLRNP2GD58Y8i50SVfaNOCbsbF6hjv5tmn24lxSAj96Dl2fwjK5ewEb2JJ7
+LHvZHNhRwl0puXobDDkYP6qxECI9xrwCPbJ0UuJR2qUbGloZk/sR8dOQjT+
s+P3hdIcCeF6hx9E4bgwk639M0Pxnk9tUMYAOb3PB1OuEjE4FX+pkAIjUbyG
JMPLRp0jX53HHHg0Y5SayLsgwHv/51PevTtsRn6PIMP7zQu1cpEv6JJ/qYgQ
aRdNibRbIdZDLMW5fgvcXtpvz983WLFFY7ZQyAGqcjge3INK8MDvGDmHt4Hr
HK5n+hFu3jpnVnvazcO4BbFeWW5gq/iQavWIz9PgXNaEUAyVGdxJZy51NTTP
pHnq88/oUAQrWPT4lm/awcuIWvk/1TFEUBrIi8iI/Uj6kWuhenxRKTTacBf0
aUupp6ecmDmocjHGQ8ujr5CKByWB8YrWpIivxCrYHgDBzWb6wvpnLxsC1Omy
lsvqnUjY3o6WF0ybdftUV7AWEf0/bCRpFoZ61ca8L1RR+sIm0E0+cdOhNtMK
Y95oCnPiuwkuR3NiOpznRHRpNh/6GZ0Zzs2TxJyPtZONG6GaYdSLEf5fnc/f
SQk/gkfX0vve2BoygDpZPEV4TkZ4LLLP/a9jupPJpZDnDv/PtM0kwWUTVejo
c468AcrJxFhSCcVrMH+VFRkLPdUGkrkFZLWa6BfgPWnvk25nGgHPDYHCEr8u
FXdtyhagEsMT/6Rk5UGwXuSYMfaF5jDpb15yl7lc7/BLOyMF4DvoN4wqADT3
iotiuESWRiA5MeBlDmZjDOtGuaXMpGXdWDwvo71PuJeTPNkcwsbnrNtm9MsP
YHequXoChinc10LZVsal5wZ4OcMAo8bzFvl71JTIXNQnEHQH5pTHgOPPxlJ9
EUSIfvyghBbKlwzgy+9bCn0UisbouspNsxGz92Sncdkp/0B0QGvd4EJaPuCX
2wu2WanueyP/z+5Xdeqf/t0oGuxDaqcu+djn4FFmBj6nzqowflSmNQMQ2GMu
V4X1Ke8JaDTdzh0Ueo8oWUuTlJ2ZgW0a8x75j9xAtFaZW1VllEJg5snff6am
0Ijhdabe0W5jswzwzU4/pp9XwQ7BZ1morAWmsIIoJ7KyldxR8VVRgWy/iba5
k5Ol526pY8PnCUhe3mx5BbFWhvVaQv25a+ZHW29F3nQi/qYKjGrN3sYixMEM
sPY3DvTMKXPUx11JtyMRaF38M6cJAZSAIMBSkgDVp4mK04xQkxQc3W61hQP3
RAoNhvVOvC9A3Az6oWXi2r3wZV0O9nUzCun3gN2BvDyJRFRfLh9KLGAX3KeY
4QZO/r4KnLkEfbg1b63QTl0oH9ha3c6lW00wHKFLet70sIEEiN02aNEjnyW2
LpLf+ygmGdJtd5rfGBH+GchQAmCvyilNoJ1tQ8LJFBM8oAQPatni/OLRCDLP
Oi34SrvQ707GGwLD6/tNQINW3JT5CkRf6habCo/gzKTl0ESkf9TnUofs9INv
ODgL74xqhSDfyugFbCqwxM7H045jaA4WnGWE62RxZ2qeSwycoQF2uAEiTrH/
otlF2t6CwmClbtU+0cqxyrSYZ2IY5KzO8CuibI1zlWQwsp3B27jifjyNRExy
prn6yyWBtW5+8wy9qL8KaDC2h2INRCRC5uvbspLvAtzLaR9mGR+NYPZheV3I
vpUSLpb3+wYZ6wXwtYj+0jIpX9s8hQFHMQdA6m9d3Vt6IsR9a47PM+WtBOZz
cu2cny6X1pkxr4eK3YafMYJpjJW//YpZrvoHRCYlkYz87S7ng5f76tDFySvc
Zw1Yt8qEMjKmdc7tDpy6BBA5Ox8TZ+C+v/6/tIBY/U/rTx1f7D2de3E6psJL
2lVGqi7PUudEBG8QBpg6MHZ3vzCxqZSsb+BWZZl970KcEWz73kH6Fj8/pyMc
4mwkGZd8t7UYvosb+uHQEogSRY6OrzGe3EWIa5N+ZzJm4pjT7dQK9p3vB6H2
vYL+zqOFtvdm/P88UeVg7wrg8aLGmrf6GDUCNWQ3QHTDRNyuUM19i6YlXmvf
RADhESr0ScQaPWhG8FqY1ZK6noviLk4nRhqdBopUpfiMtib3+3IC86zGk4wh
RODp1giTA52mCHHOmi4YIzvbsLuJS8srR8XOlairtxaWS1pW9A6uCG0rmQsK
HCQIvmyXVDzLgooA+bF7UEgLShKbghEXUu3AM1Zn7150rbGoR0gqpXxKZNGE
yc6Hj8R9qhWff5qUXFKNgP2E1KGRizJKx3wFnVBfagXMs26P+f4z9dGDRce2
M0VmfNJgtZVXUSd+2I141FbUIEUAnfCWlrjtrYnxWywE0RYLVVl/XNWnd9jg
jZH6I1kq/DyCKMesY7pDIkFurytmpcDrvOyDNkdSYU3ux5c1l0/JY7oPvupu
K+RaFaMWlRg+YKjfP8yZp6tmoBF1lVuw7qIBynnpQI60Vm0BDwxzpdMJecXl
fBrR7uXrRtVNn02soclabAxmDhP6wpAQlp6uC8mBCNs0R2LqlpoOqj/oWzQ2
HcefUMjDdjmFvQKjf0h2vDjmgbuuNvoP3xG6O8INFB4WAR7twj3g9A0HBUpW
SAzBc/MmLTbq8aimNQsSv5qxmxm8taEV3HIWOoNFir7lbdeiYsJsd/O7Y6a0
BLkuE9oIrGEYRfZq/dikiqDFWIgVKBVS+FBOyHzw5n26gOk0gE5pxcKzWBoh
fCaPMDtZFreveyIA987cml4DqLxKfM0ZH/dFdlXWgiCIKYaB5BEpMNIq3D4c
+DrXYhR9/DKohIeXH6JndOQ/pwnipa6VG0sfki+8SbHw1CI2BpNBiQlREsTp
TxrS4GgAiNc3FoePol+7sU/9zUOggaTlKu0Ky3Iss0iHQKIK8P1Xju1sV3Qp
7UVcy2zSNvTBMWpDQHWawyC3JpjgiD4jyllkt8lRfea9tyKKZ+Uxa40Jejzw
FQqNcH2wtLCxQJgdkm1+2ftZr0mbPfYV6smahr3OwOenCWyMJHZ0fKbl1Fas
F/Jfs13+iRgvWZoQYy94+oYATG42NVGt1b1h5nzt5vBf9VgqraGiXPglnWJd
sFjxeWhstFqy+NvaWlfS2Bwc8ByJCfjiMdq44rrPeyWjYYxN4CWnf9CyrfYT
QtEIPFPYfyLvfuj85JjW2kvxyIu7+Rijaknx5NHtdzIyOxMTaDFT1xGozjKi
cspFisRxc8s0rJocYpKO8aK9BmSYywEJ50HoveJJKIztoqNJMU5rFIKqs6u7
bA/CWf2DAR1pvTw3N6ODroUqjdfF4KB7TAmAe5c2pIfvwI0jEKPEq2EFjVCy
fgGQKp4FPPQsNK9bTq2EHaV859qP/LiRLi0TzX4B07dn+8kvbyYJczSyjE0t
HOm5B31ONz0Y2/OOIizN+cxGdXZxiX1NfDJoOL2dMWzHbGly88Hyi3sBBb/v
CA0PBAxaJNhCY0xcYIot3imqRiuENUKvtROfQ/Mw/gHBHsm/HgTkE0n6HsZK
xVH/5LE7dzrFNMS8WsQ1tK9bAPS88HhCO1wIrP8lltgs/a9bUTel6yxICIE4
oJVPQjD+VNyUe2TBI7tLhUYcPIDMpRIwrpflQDK0aJO6kpZndY89iqvEqSqh
tp93f5TEywep2FrHG+CR6IEsAfNdpBLgVKaWj6/0rb0+tRhzGowsLUt4uUj9
nbOwsZ2Ti37FTh2jC7NggeKvAJqSS9AFTKtM0qIDKjsLpCo+tQZokj6obXTH
5pTbZno0dOzXUQcHCEFPqHbJ1+AamwTOPfBC5Dd3UY5WjBNIhsWL4N/XuSGD
BqMKqDuFUJmqiIoHt8Dwxbgj2rx4ODBj34FzQsMOd7GTe76aD9e103FVrVKB
FEjgrl4Yin96BHVrqUp//HisCzPauWrFOPDilGH3mB/cEo9fCXai/SjnvkEr
44obzfFNi35JqG9nFvisBdhz5wSRtEVAvkDqiVxey6edTTNlzkWXweQ0T7JS
Ukb8Q1I7ivn6MxuYdn93W1fWIRjuNHmjs0SwhuevevPIevPsohxwdEKE46Se
v1fi3g51alEy8wtRnThksbzlHWC1ZzjAZbbJwsQe+zLnbPDTmeBSxSvti21a
eCm0Q1xQopfMJ3uCGBtMiocC5CWloDPMdZlZJ4le1LNmUEb1qw2Cyy3srxuK
5DGOtjU/G53lMqkxNHif4dPuTqnme1lkOZHh8cQhcip619aG5rAucykzLyuV
zS3h+LH+3uSvMfxikRdvOqfWaGwEK8v1qIzbQveTYmlURF9dpYNHu7lTF14X
+42dOlurlHXCEQLEX85NfBxbmSD18qh62yzTnJzhKYP7zIlUY+mChDMXMeKs
Qr1z5Xyeph9yzePEotf/fSR2BA6pRd+zBjOxYljoSofC9ZXyp7YCbfdgnDZ4
zBjXGjix9YEC4M2b2gBfGzlZlF1yotegB9v9jHHQQUkVKmsPmcvoEOThQRQt
8YcYcwohXWJ8X9k5TMXnSv1+Cm2D3HHGbYE0IDIkms4olS1JmGgfJ8JBO9ZG
Hke7UUsl69c/C+/cWszMXMRJIbrnP06u6j1GzA5uhIpjUnkGUmzYUI7D0uci
dUDITXoISagsukAox2af7i8ZscHs91vTMBlERRwM/7bq9gxegNfq2t72MfKX
bizEAhuyKkzEhRStoKw0iQIT9cCm+odKKqQIiAvOtBQt3CIr2XQvVDl5aFhv
U4HunfAYkZTPi2SSeCq9D8q4omJ7iIs4Ig3BM4UYOGx+T5PhAFKT8/pDGdSL
y7CV7WMS1P/+nOGGnYaWzPDHNcePaQ/L6OjlZVtZxxwEckD4tmt6OD8oFPts
t4W68uPhsoOS4L44NnIF8oGoN5ci/Mpdc8kD4pW9RYiM632I17GCeFa7GooZ
jcN1AAOQ6BOW8uWUgjrK8LX9ySawGS/4Z9MK9UXCgdhb0n2UsnoRBzwunh4/
tEzBx4HZ9yNPsrQgP8ic9u57X+INaGINnzCXYCJb+6eP6ff00eoU/zaAtSTP
kB+LkyQh0AON7rr0Ylh6nC72Pmh8HaZo25+T7NMR63wpVq6FpPYLcn4yhGPP
8LO5a3/3UwpqlDSGBX9IXS/RTVPS8fjSo/9RSNpZ+RdMCTvRxlWkNualoA8b
2cuEMiqTSpS8+vVCNjto+6FywDIjaw/8h5IGw0lGbyl4xnSKFa8RpIfjG1c6
nDoy+l6lH4CXx+W78j2pu+TnAATC/z6UTbfXTG+0O3/uEr4kgc8XdcpE4P83
OxNwIdszryWVZa2RwgrEq2I69uvVqw9HbkCjvqJbK8UaIH/t2G5IdaxxOkr7
qbVsK89Tc18MSUWqthPS/dfv8yEkeNxBl98qsyE9JZb4AIsxzbPb7J//51nD
byvgYkT3G4wp9Wp2/SrzPQwztv0LcqO8Czsf3AxjpInZqhTmJsw38XYw5hmw
fDzEKdvaUNNdd9q81NgsZy428yZPdY33V60J+iZjpnxU1uwjQPbRt4kHsWxn
KM0g/GonfQBAh7EcoLalexbJhPyYEJwuyJBxb2X24GMRqMC/IQ8Y4C+KLq/u
OsFBdhRNnjs/Z4y4ooN0iuYVij1iDezszxnk6V03cw9ZvhV1qWrxf7ZzOCiK
+O8L/F0Fi4JuZrq0c4UXaYRk+l81yXNBJP6aOqg4gvvFzUSq2peSIEspAPp1
G1NAwaanad74zAIxWdnvtc/F5VLEjIpuLtNl3eBIIZPgLVYyH4CN0agV6gW2
26jjpy9H3FO3uiNFYjusQd9yhb6vtfyrM07SjepF7PRlRsbgt/4U8fUFj9VG
XsIxoYljU1+r8Hf5/I0XbDb63Jml5c5pd3g/COiCMr8abAQulp/1h1TsL3yj
rPB6/oqfi1Tz5GsVZtZ156/75Z3V7Qz1Gjr5I4EStPXGkm9u1k0BWmg4B3Vn
i7A1kmsWAcdGgNxwTlTW9EX6cgwbX4rL4pK2GfhqpgpqI8aZNSZ64Hwi1CX8
y5xuKHSlhW1Msk+kCl8HDGsHzyCnx+zvwT5EENZ8swgzDL6vkSAcI2H812vI
Q9Vf7/jAPVHD9b0Wy4vn4QSRgzMdxrDXmSd9d6MiCVhFVbf/n3NZlmSxEBoH
+XtZmQqVmWUdt5dh9DlNOQF8NoAQ5CvpoWGZK1q94qq2GiKUt8+wE6poKyFa
NKSnAKdHVYuF+VTHwHhSMPzUIcZqhJrWXbgJqo3pYPWsGFUn853F00ARrBPT
GkbdRJ2IeYh5Uu3pPi92BqkFJRDv6jA8F1aKIlxw971AoP/B413Oo0A0QFf5
Kw1A1XTS/43Qtl9S/IL3WAf1Dvou2uWJfEpYRxv88ELTuCn8iilrTpUt1I9O
dbAELPbF6Xu+o9QQZnfNgLcNB3/AlaFooqkfAquH3MLCkFnW8FedwCozIvDn
f4KnkIuSOP/YH5MrGpaNZXwpHPT9qwd/RW3dzFOkExBjyVrAqJEVC8xTn5UL
S1s4q6jfa5Tetp0rVy1XVZtm8krj8feIULFe5ZOqouFeX00e5WJHbHElQ8/u
NwC2Qz4Bx6WhLyzEiMPbrK/uoIrwIQf3JvWLfCM5+ZcDuBm6OwPDQLLB1m7t
ZSfv/KCIRDwnypZ97Aj6u++qZpTgFc96vSf7D+ik9+znUHVcxoHKcw5Fbqej
anJQ5DmnEdni644/P3fXTG+77U5sqcdxZpvKWcVPKphehvDDuCOxlNatgQcH
DnpHdlHWcs/mHYKZkNRFOryjN5P3KuPpsGYDdEtSvrpBtiIBCu2AkmbTa8z9
/qdyaMVgxsu9UetCYr22iBgrTyCgG1o9t552ntOJmyjt5G3EbBOySx/m25oY
sU1ygmNrTyk8/72CwrJtIyhpzFjZLGpqpEGaOeg4L1ALY7oNvH1vzvT75t1R
A62yRAoMNG7OjyKqVzCT74EhciOrpS/KmtUQBmSpYD4t8nLoQ9tbV3t1YiyK
DpCG0KgwdbYZi4sjHQKO/uGJdqGofuYZOlT1/XjK1vsO7sj9/tezaCVlX4ht
kijSAngOmzbvPQJV0RasVfYZUMa0VHwerygS6dt19RElJ0z5zIBl0SZ+IXhB
OrkeuOgUcPwKrFX3X+QnAjJOI2bldSmtgNfVXJUjoIsNGIlZcKAH1iELt+XP
jZt2DNQxTVmLk0UgMaKXQZ6/CBjYPg+itrEUTv/CW9GaaA3KCiFmxjyOlAXB
UWr9MhOHcwBWDpTRQmRPYaPsHzeWkX+wUT3zGOoHkClDMx4knSNMMbRgGyHO
UZdqFtMw33NLPAn5xAvNrePDueKEgpKzUF4WXEca6tXrVKO/+UPggu+TigDf
83unwV1GcUFhawlo/a5gLoVl2dTgERB+6/7ABNKuoZGI5hIazNE4mYxd5pD/
8XfQUURTCWL6PbWGEhgOqY01nQwE4Doj7uQ9MWTHWT3/ubxtsaEs4C/+PP/d
d3p6Wja6QOn2ce9QBbBsctGNCp/NAnqsm8vHFkDfgoJJJcrAJijBiduMfo2u
p5v47hTahOCic0XkeKP6rNoaVCQ098sEXg/tS9x8x4edf/6brakGhz59+5RM
rd5r6ugEim9OrpmrEqZDdnzKROmR9bCYAkFngpNS1Ost0t0+OkL8Tqtg3yP4
wK3GDJgAYQYOUDKnWnEJlUlX8pFvQqnAUfbolBmrOqq/MkMw2xPZB9F/zNzf
pc4VM3Lh2tRoDy4F6R8d5Db4oaxjLzQE52sax3iY3NojuBAhjeDOwnX8xR3R
Cbotq92jh/Ef5G65qF3WfqForsyGMsizcvQnJCXhprBaS/5UrvxN2kzecnVV
KULktMYMCLQgh4rpexHyQ+ENCMY0GveeUg3PztRIcux8AmbDi2e88ldDQ0zB
Tb5ZhaCIZ1rVDnXgJ6yyVBR5v4uN6+cxEiY1+MNxuBbWgxqcv7IyaybxBfEW
nxRQp1CABcZTj/lYb2wZaK1KHAPyQ5s8QTOPWxWvoeY51OSeWqz9tzjcSNQ6
xyUeoU0IloHA+s/yGjL5rSP9CKT1SNhvfxImRJavKIH9ObKSMxFoVnKm6h92
lpZCCB1gkCrluICnDDEos8dkUXLa8zK6GoiDE6WlrhfWAswe0mjaseknNOIq
IM5BsyObE3bLwMvQQabtUVXx/pI5MGvtFPXUy4a+7XlRqbPA45s2xnox4yRB
6LiwwV8uvYvQtHBXZIYZb/AJYkhPo7o8K3TZCXXLRnJG/kN1GHULWIzzxTt6
g8t1RL4YZMeQKP8PtamU1cpmEdzMQa/VpEDmZppjif8X25bEitKmeZJwYkqu
FYicheynW4ONG413YlzcRI4d2z001VD25ZJXqOvFyn3jV8GBtG8f6Ljv0HvY
4hRitW7Zq8SZ10bhArK4c73FamDzmmCwsPKP4QtEGUGszJPFVHFfZ+40ShGU
ruP2ElGurJKAerddUjlff0xhmKoN6BBdr4cYe9TCN+At9jw4Ll4CBBJ9MdK/
alle0epBgOgwW5YVm4mequZbLFGe/34H95FRrG1cSJpi+BTmguGhUKNnHnoj
UGFtOacdxi5DTlEMC0jRvEu8JVd1Dw7gXbc5pXTeJnMzh1I9Tc9YghGvsB7E
19G5psyUFEh9KP+k2eVsEpuMUGO3+l4wkf3/Ytp0Xgvcs47HYuYxgdhGxoL/
EPINSBOR3QNT9iYSh90szsGVQ3d7/VMI6hkWnNqJBIQZzX/1FFZOUCseTMbT
vhyvpO2JGJDPFEXFcg/Hfl3iNfQe4BVK2YHocgG7YB7RlOJ9BpWzs/zUpFpk
EMmaUkAmHojSk2t29xW63QUgi+Kby1JW99CjPxNxu0wkMQr0sxBWoWCGkHYb
KlAlWZVkBj9dTIVhJeQQmITSOkhnX1HQv2//TzXTiurYK1xuq6EU262UcNWX
MtaC6XPjIHq+fwepSeZB8XJ7NpJU1PmJjZ6PwCDuynhRGn4RTFfKGHg0qb6w
6LT3duBSoUIXU1xKD0hoY96j0jhWo7iVLCjxNM8URnq5otrZPfG2H/LlT7BO
qLZ3FkrCVqL8UELYLZB4zWDUZU7LKEUHpuOc5K+GwVHA4x93+xZdFab6UiA6
krOD4rgRdqazuSvwuECpp0cngVtP8NRrzqDVqAaB1MQT91bkLzp8hn5vyuyo
t8u6jUGv2nEEozoF4bEDxfMc2t4vxgFQub/cD3CWYYjfxChCNhTbdG6Gbapz
NpChuyFxplwQTkw/bur/QaUZdlrM7MvVtoZZUe2nvPpLSb5aX6S+1XLu4rSD
3AwPXwl0nLHMJ+HtXBgZqmLOH0SD8gazOcFVHIv8LgxvIPP8HIPK4ukFw5xp
3xzO1KEutYq6Bl4T6IG60oQNAU7M0ZqdkwdqaGPag5ZNTu3JxcxJ4DLfraZR
TiAv1YVRMH4JBnQF+hwomzgloMytwF6tezGFCPAgTUaE6gyXq8ZxcrfItSzl
EnYfDedsfYjtYyysJ2CvIhSInClBEEkp4ZIdzl6c+Bf4Q913ujGR/7m6AOxI
3nF1lgwznprULvYs2+Aeb5t194qrOXrGzkiGVr4MloUCoLfWfgNkXmVo9MAE
gHMF+pBQ6++BaomlYvd86Grl8PBPZ2xZEGl43Ig7IYYuSTx2bvQAq3lRJCON
IfbjI+Itb9OIkN2qx12qcCoxRfj+nqvZ+vr0Dt/1vj0szostXEj2pqCvI5EG
AalGlOAJU2pMPeUSycPBR1IceKq/3mytwjbqamvjOP3+ge5JvJ23HaSti5Qg
yPwkhPqyM6Zseey5RsSnf0c9TUHMqJnKbBBXjXXRo+cWiWPvQOMxEamNcM0p
MBXkyYJZjl4IslhZERbdlbGGuHya1zmLtPQpQreX01HblRS+5WPEOMOLiXhH
I2Rrlxz9ftuMN8683J2lK0nQw4VBRWh29h+xDCoGNTG9ej0ogqNEHt6OWS9f
a6N4vwL+IDBMMtLTJvBRuG8DX9J39Q97pjaB/b8VyEQBV0Aje4RPncJxvLpG
2Qml/CeN3eFfGsFTYH1Gq+hc0u1OWBuCZUkuk4N4Q3dhI8nwEL2EBvTRJXo6
enM2BRorXsrMOndDU8R5qI/FejwC/suzzgVXjeOBR3hOtbla/SfcNOsyehkI
+lZObHtX69/rv4U4WWSnMeTX2NxrZYKFwHp4W50UfgT+AXe7CCpS5xm/i9a5
JqSKqOpwJ2DqEvyVAkUn8kjOJfz6EBWESPpsHNmkPd7gd6fwnh5dYGhYLujj
/kKWAs8AtcWxkx5tCLGNGYDDWIQiF/oc66rhZjjaC5qFkE4g18TIXcFkZRA7
kM6ZN0nigs0+Rpb6Sg/k+EyhTgeFe7xr3+X7NRjkuusEG0MYFuupjpwk4Bun
nFZBoeJaQmcy+XotJqw88II04z2GbKkJsF73H3zQOXLCV7fuKDAFNhyfNJH3
4yXG1Y7eM1Nqz3mKTwOcAbODPjo+RAQl8xzRY8erfa2Cr1GYgFQUTBgtYQok
vXVkAzNK7ioVaBClh5HzJXO0Yb55NKJ9UPYgTsYoRmYRI6yxIL+kwUs71VJf
UxX0lM3J8hzqL6trs+9nuH8lkjRDhesM8ICmJ9O/xIXXGOV4FfaZaHs47PTj
PCHJ9HXorLkyO0Y5Hp1GR1IRX2gZY+wMJ0SHgqto9u4Aj8IvS86PZvbtCPmG
wlDQtUBQ0Hzc1KtCFSlTuh0dKQmf2bMQ1Wf3RVQSQA99NhzzAUi4o6pgaQ/y
puPlEUcnrStZUe+YNZbgiL8eP74Tvn2PVVHWDicpZ4yaj+t2LJfoO6uYgxdo
cMuAl6wULB0zHS0af1cEz6EBy78RX2hiuF/30SXuQsOGVqulpLHbVhf6YmWK
aFiXvWRH+vF+Kcb4KmTIUhKFmwYO8KFjSwSHYIsuiRQ88ku1vife4xS2d26d
zdy8ppw97weVlI5KhJpBQiOBrhBYzhV3om4B33cA7m6MRvsORvov1Oji8w3o
eik+cBdpZ0zPa5U94wAuuLaB37HoTSGU9UCx4R+N6gXIa2U7uespAr1tSo3H
v8/6TO6yNEPzfsD4b6LQhCK63CaAoncDrMvtefLYZ2H/pRyOvfMVnKBVHQ9V
hLCDVrMa3zm/tbB7qbUyjEaKmkrAkQz1KowEZGd0YlDKFA3lUCuK6U7sJUu4
MIJIFLsuHNFL/mI0mjN36G8rxMeOCoCzuGZvbIua3GaZ5AMGIGK3rdO4MeTz
89IBhqdZRPtLt3vtJ3r1bmZ4dXc2/OlhndsNsRCZbB7/f2IZ3sZkXk4IlA/q
o0ELxIxgIC6M2OiYNbyRcTUkz8+RVTRwyphPp+wq5f96Xr+0KQO6UHrzzXlZ
jcxFMDA+vci8cYO2r7wBiym0QDxDtuor2j37nyJF1fKweAhprlZ7uFpHRreW
VrMI7xoDBaZZGaSR1PCjlshFrtwt3kVil3DXnmgaNib3hhfcrSnkC9WXjvqF
8Q3PxTD/wQwP5V6K40VD4bB7a4f2skIIzJQk+Q32/GXSaH6Ossa+Wy40w/Fd
U6Y2cN3kQ4omaCpielgXC64Ro2HdrakmlLskkEr3HQHA0cCaObsGs/wQM+9O
vX68NWiSqWyDD/qBAvdbojpvC/peYKZuRnNhgaZ6WmwfcWQs4jm8APmXxttt
1KYdmVUgC+J/zu7hKVLEE12Wijgx+FSLpMfcMYv5SRhwwsLRJJZ0EG4w8WWe
ZCflQvm0QL21hh6QkkkLjzHwleKnRKa8VfNNUpWjgyExgD1QZ/vZwKnzTlwL
C2IVOcVymtdnclNO54nn/QxLGUtIfQ8eqblmjtd/N6uqijLDowqS2iU+EY2m
YD/QcD2snCuD2F3C3MkwSbrn4kdQ2cGWR0X+jndAZu9X8OmjO7ZXyJ5aYMn7
J+d0gz4aDeG9uD6vabnOLMjMfMa34C0Mz0Rwr16sYxt0VGQkcPG1X8CqUpkX
Ou1oW6fNyAaI1s4r85yGhqibXVTD56e6BdiR839qy6C/xOuUKVsI3nSsOH1/
GrMpU9lMZKKHrWqJsMeMQWJelZxwP355gfBvkUGPCBY2DKh6YUkEY4vhW/8b
4kmSwiJLFSTrz43dSrXCePTSB/NJaK4vldt66WeUPQCLEXRumpfpG0J9KB9t
FpuRU6iHZg7WNGrD/kuq8XSJbx6Dei/pvY9GNrNZ56jgOaMpzL65tvdkpBES
3IoB8CY0fCLcN1uIc4d51Oqvrun6JQbbGKpiKKJqhw4FrJLjz1C5YDY/XhhO
BilERFrSxdsaWmEfWwbwTuufYtz5lbmduze6ZSlI+e1+e33v4fyEb1nKfrSZ
9MWhdzScmWvC1/JpIeKON31jNRiFEplxxLYT5ssFxLZi+Pv9apWdCXVRaojR
qN/P/I8frCl598Ak9+tPxwW7gE9DmMyPXSizDViPT+SIaEwP28+eBhxqQjrs
VCqTQnZYAkDmgLJ3Fn8YfMKo1rCpgeGSJMAC+2pdvhC877XBk9eXYsUfsIzL
1vp1nyBVL0YSxtf0NfGYVhxGDHwIA4TbS+BMeY0jYVr19xfZCY0RODE9qydw
UGnK7xCqqaW2z70X9IG1PJWQvjIrrGH/Y3ZvZKsHveHM5jCnfAxfU8C/Reuq
kULXMoFtKoljp6h0dBGJMU9FDgM6Dq1QpI0jkRbAEbVakYNog8mYtPqyrKCE
vntnDo9I+IpHZJ9tBCVOuL7XgxEBGzx4bZs7vNGJ6Aepwtz+RbAmUZDh5Gav
yvnqjX7cUfTXbVoLhh3AeC7wym6aX7fVBno/g8QiRsd2I+yThLSx9TDR3+gy
A3WkWrb1X3/vNnLIWuM3lsaToTMbTJjkpwdSVxcdrEH4xpaPp1x/NQaiXvI9
CFj9PBbmbRDi1t8fj0eNOTxndW1hhp1yO246lO6zpM+0GzqRGn+AYSyDa4l+
l9+U0hYCD+Y9fGvtbhsqILSfWVWP5aEKXb39XSgBL5cNhUrfXrj9omtmLOwk
zc0j2blITgFOHKGNb4YN/RMSZZyPtYFChcPdGuvdUwfGq0fpeleH9dZmxGCt
cDPW183Se1+5h1zLastqN75621lzDTBGXHelMN1uTsxd0eyGT8A3JIxvdBOF
F+ye7/nbHjD9mdRhGUFrt4bpk9puVwxUyCPGJBwG4yKq6Tadt0QVeDD8cAes
GwYHXAE8YD+s/0pOnYoHq6l3eaVbBLHSO42rQwbXY5PLQjqU2tGlgkKshuwv
LbtsUPLU6+NvLBeVHGq3fsoB1kR2zPrHvkm92hkPIzRVS7siTbFfrOUYnU8U
UDOIm9GIDMeF2ciX1ikFhhc5lNJZQrCxaXjr4y48dYP7VRymM/Fmx1+kqS99
nrg5wUFQ9GnVIUuPtO2zfCbYa97qTNb6pgyqTwPpZ78s0HXRfpD8R+ZO6Xwq
RFbzly6Ggdh8OwjukE8iRHvFt41JtOIUPwn+/kub2OpBmcsGtYvje4Nlo8dW
bAFiN1pqOfGU8/QWMAzOj/w8GiyxTnkEXMFC31bqHf/UlwaaD7eUvjWm4ktB
Z/2zLO80HYrwKPcYBt/mrREK4rw5OjZ6Bs4sxxRt69yoQGRLoK5ACp1Ormrh
R54q4m8KRHPiIyh9Qarm9M258hGxQpJpfhyD9FMIt17zxqHpESjKL6y5o7Go
0/nn4n4Sen6UqQ0lNknSqfQDgF+Ucx/T5R4DUA/aiLESnn67g48mTh2GxL8A
M0klfnNM67SEmSdvmIrzvSmunCKjEwZxlJkSrOJAMvRW6sn3LikxzMT8Ld29
xgSDPfcu8jRK3iX7MTTMsTC7DUAPwUzYCTfYBzPGaRdpAq0hDKMxquqkRvjG
yVWtdSOrgzX3OtzMR+uogOYspYbFevzN6qe24Cw8Nl4ef3T5Adc10zDcVYPT
Dp9q7iahZigMUBMpjo1Vr8JaYL+kCKvFoksIGdgmD2HVqu5M83U96DtsbrXM
js04sSEC7N76D+QpKhNnTNpG484qNYnZBWsXEv37tThPQEoW7nNfQ+qUwJuq
TxgLuwttXzTw242GBGy7vcKJxvVF8/j1zXv8Fall8WZ7hcp/aaBC7FsL0vs8
h3S4diRd65yizJZ4mThZgDgsBPdJi+BNEuaoQ4l9TwDCflR81/U7q1L+0Wn4
hunMVBF2gIwiaZrvrBksXiGZFxTtV+BAWXOWAHzSXoYcorNPngd6pmzawTYd
o/G6QSrJPpGFav8IprFJRzzUKTGAlLGavdPEQNYGLLqHssOko5949Z0UehSR
stDc0YKnmRF5ltIxfhTXHQ9Sg8f/TXpdTOqjpkdXICw41aRqpcrZzZfD/XpO
e0s25DtP//fvtmW5+72+bkOXIkP+6ykHV69BGTKqIMcua+5xBkcJgaRRpDHe
C6PCzrJnpehANWtxJIXpeP1QyWrq2JpLNvsuD+Adf7TEqiSMF5xBIapKOPlh
Kp1nsdVouLJbQgZDIAq+lBFZGe9uGAxZvKEuxEo7VjYYdQaco0VXdqQYj1tE
7zgep3zxluAJBeBYraDY9LLKeFIByPPPVnE/IdJ12MofMeCwJ5dvPaT1SsBL
QMhzkm4+ich2aPFizBFJDkVQ5mDEP85NTtpOQtgU8h4o6a9xu7dQ/RsxLNjU
ay30z8lHYCBxHRphUss2mQ97jgjzs0n/II3V5n02tvyaq3kqmpYdMH7oaysJ
mUoEEmO06ClFAKdwns3gDp6zSqJUCFi9XmaFnDzmeq27y3pDYA1cknGlZnzA
r/MuxRMkpJVyzIS7DfImdboGQOk/rgSXEBNvsF9SP12gUq4Pq5BPdrtoUvoq
ylF31Lw+CcgOAhtwJz2kzDw8RKn3h0clM5SZfIWIEOIYaPrfWhZuDBUzwdCo
xq/5ooAA+jzTByppEyn8wUSUtK7MMQw9oQePjPrmo+j4GV+uL//uvgqVRUuP
oQHzC4JoRc4VaxrxvxRO525jt+BM6Nq7Us6oCSK8Nh24iXzn5EM+hey9o1ln
DPIjyxqvmwSbNjhI7ZRg6GxoXjMTpmhQVrlQLeEViF4WzJGYTSTJFsbqPvVf
f3FE7CXSKgC6h2qk6i9rDj1UsEGPylw5s8Glhue3WKo8yX1lxOu9qz6XOGxk
qF5ZMSWRf0svwlulLt45fN6xKAP23tvtLIWkC6veAV5AvaJNrqaVzIZymVLt
YW0VjklBE3Nf/LsaNDtBqv4eaMyd3ciYcAis+8+VE6YpA/nVPRxhTmo1IZ+U
mch+PCzOaVNKa0Beg8nAwa6xIDbTMC3NPqy9885EZFDrLj3HpVVLEFzF7G41
LpA1v840sod2quxfJir6ltj9JyMSX2HzuyBKpX46tCnYEV4zKgHYbsD4SioB
dTXpGbFn4rhnVyfKNQ9fvNLHhVOrhnWW5Rm/zzDLUfqyoU+tCCUSsGSPu4dx
B9R7VbrFLQxVuWyf0qvPEmXOPR6j/7RN0zC8ncABvx7pplEZV84EwgbXahdi
g1tt02FLnTBwgh1tIegy5uQ0Fy2MglPVMLYt/TkFw7UQzA3acsT743Y6BrK+
kE3lUNVgiteH3AcB4Y9uCRXarRPqXLfBYMjJn7qvZjOzTQqenjx/9yUp+xz1
xJXgCnGhOh/yh/fBRy5tzIXyuzWp2vngYlxDKnDRMGzIpik83WSj/kYSVaxo
omNeyC8CmbrU7pId9EjftWqV2xqawJnWh0K3TBi0R3irCx17i7XsvpyaXnDr
jUHb78r6wrhJlIEJu0iHcf9WZzrgBqW4FeFE1HGpvEbdgxh8LxfAfYeOQq67
85kfzK69mMOBuXBhivkquYb7XqtelsbVROJ52eA8/GEzjISIiCr1ALI1hNCv
bEWyatdTbqzZfz+5xBbQG5xj9A1Nsf7Wj2w6AhgBvj0d/apDZYdVpPQmBTBT
W7Y1Q463mA+iiLQOc5iyDgnhrOvecRfCoSJU4ZnRGTwpMpTrk1Gu0npB2nC/
ikxJeNJAvxEDVbX8VlMSsjqy2Xicv2vnn2Hdn2RdxL9Ku+Oj+eGFejZFBoj4
9r2d0nu9OaITlmSx2hnXKtt5BuPEZwwBePo83ZjvLS29oJJ7B5+LojpVDEmh
U1Mf6XWjcFZcn0Eu9n8sku/8F1xRdXgndrgZGCOfXQordQNQDbpK3ArfJwRh
IMFss1Pqc6/9tRkfdRwxUAaAbhhlLtOANq7tcpMvqdGYTn3/ZB9CYMwnwKbT
rEl7vu10imy2p0MGBjD08NnBjUCdK+qerjHJCBVj5Xy5vLFg6L5Zi2rgmdDc
RaR6ywup/9WX02HalcZ/eGDDOsGYyNDaj+9aSRJ7K5yDyQWCAqOkQXX0XMiE
tjAgxALjtUI2hdAYkMZsYMawzuXlzkY5il+wihWbxYi6sVgVHYXuaj5ivtV/
DTgRw9PTy/sytmDcxtY2TmF4MmI13yHBaU+ZP+9RzOqVwPNiRU2+C/DweTqw
7a4NXiWL9mVd8f9K2rOnNb8MD/daeYRDpd3h6qpltfS+i3dMxiWCJMMN+Ne0
+foHTYTjirdW5gIHGiN873rbSbnuvHmcvHCps1eE+SaCPt8oj6ThNPRdnf+P
u0V8c71UJB8Ip3Zp2N2KSKN/v0a70AuZrZBCjqScv4YhcuzTy8jbUy6vOuLg
MLJ9c79qBLNIoZdf8l7RDIjb9aXpU8PicgXhGZP0Zx0zkS8LU26vtS/smS1j
e/0GC5Fwe4jlzyYoxPQ6Pp5hS/Bmp4omltdpyuxtTCueBPvNmiY3z+cpiJhd
E/fSlY3YPzZGRxhRvou73E3tdzReNDbsazoJ07zj6+dsahXLkfNggFQCDNN2
0Ke31EyDtz9Zp/VXDz3gYaviMa9nvCwKSvau7tn2hink3IRA0Zmh8swj88ow
tT2qFIy7sVOxlcZbHSepcwm8lXRi6cPPFj6lgvAuGgWtkP1FOHWB3j2sdnhu
U5s/NE6ptYp9OOqYqD/7WSIUh9HfdFlVhomQpyLae0eDkBe0WAb/7kn5MH3i
GWcm9JnWApKfQLp20m+sAPnp+vcUk1MNgFQUb1yjOYi3yAtOQDVud5QfJbVj
GZl8kAjNWRIcYlrD9df3NKryGTYDFnnjkmI71qYEcS246MOc+dRYASK35ZBl
wcADV4KZJXjypC8e1gT/LJy55Si1C8pEu1KBqnzuA+Mi4zzIym5YAMY/YulL
UL2Hod/hPjPBLsNg7pP4MjTqpLkAYAzIS59bp/Ff+/brb5IIU2/JrTtj/O2f
wPup1q9FAXdtkJ1Eq82cGIBrO8K8sd7Drp15K+0NPSxC7S6/wt9LHPSrRmSW
Yq0mI5DedFkCXz+wnWV/lWjJCywd8B2egkzweb4ZiIRNDD+lw6/KEjhkWksb
WhXIsLCUJ45iq2YxQVaxRYuo67fZRvH5T1+4vuZ16DkjMzzICHaVB0jsF2ht
Oj/3RYv6yhGK4BQcGp+UZPsiuZxuarNHbAfy20pBm5HHXmZhYNOHk9upT3KQ
8/qHB6u34MMA9tT/Ab2qa6kMzdI8pSvvjQSolcvF+gWKMjxt5T3lhuRHf0hh
X3dhl8NSY7alvILnkuIMoP+DOX1W84c59gPUR9xvgz9M2Tlxuh1rI+zXScA7
P6Ob/OZ5Pkht+bXxGErJaAjhNNEahD+mWmlur5Ozw/f32MYulaKBki2Uwyco
D1FwbEQpLsDuRknO+dpLPGCBH8jgzK03yIkr/e5B5jP99gSlkYj/3NRj5oN/
cxmdHnoZePiVCvBUA9IzlVO/ysjdDLsNUvv0BHg9aRNnvXdtsJOo9KdCd97G
CzAV/swqgaAwV3Qg40jXY66kFtKzUmSzV0C4VB9NfLzSu/AVz0XhbO/bOtA+
9KwUkl81QsVa3Sojd+sPRzwUKfkpe91/YZ5x5iIuDrZ1Gw/d10uzEL8ptB/E
to73XTA8t1Z6ONtlkWClO0jddBtRwLE1RfeJxGqKuVs/G2jW0Sb4qqhXLzNX
gonNApnZJ1B6TKn5GHHhVnHJ4vNIERt9BhhEKP5SIG3id4uT6BPnGJKNQQwV
QUiSlrHS+0OSMsjsCpuuN8Z47Yrhm0sBnhvuqGcFYDbxmiQRx0L9MVycJ0ry
Ccjmf5uks/357DTfV/2fxaYmdqYSKBcmHdrl6GHFMoqPPukkRBFpJRdntXhx
Bs8A2KGTYs4Lz86VEgNE5cIJ/L/TpmyVuofB4y1oozWCKIJ7d3WBJN7Z+iGD
RHjyw1ndgcnGFe4qZw5655tMBKmcv0rQSJ/aiv2pqgNP4TaLIn8BVabQ2GXs
/cQGWCAWiR0L/1tmloWl4tt8nQg52s1UGM1n7pY688qkB3bQK/CtoG9W+a+J
f6F/HvMC1LSY9xu7TdevC5iXRscD30wAcEcbd1+BfMXGpdRSuIhgIAwoNRGt
2jbTVeOrrNsRCN2O6dLiuNQkJ1hqm0jC2lVZb5QNSHuLcHgp1TkfMbXrOn8H
EUSYLjbXR4k4NIMrDpJqxwA5QJgwgoVBebrSIF1tJ5fVi0XPGWTPLfQfQm4P
15QBvOJC0fCx5tFwAcHhOYzVnJKYweZNC7OhzK0AFddH7MM30xMJwrLQcJOK
p8guX33wMQfpGqOmGGKTPt6Btv5fBBnpTcAhkH6l4HOm7X8AcoPXInyVhNpF
Ypj1+a1wvPwZ/ty7ZmKXMxMkpP7wAPEyxJ/4rp8DKFtthedanIEYUNHYMyq6
ZvMd39j+i4nyZe7RSiE5h3Hn/02kxikdSDyUE2L7YANucxVm5GmrmAeQpt1y
SK5mQ1wbgIwFA+Em6vQ/vecL6to74T/RSxuTgk1gHU0nPSnkTHYJMK3234V5
eD7MQvLyj+XOUkUDh9Veki3KO0tlY6gcg4kIHVgzz1cqCa5AZbVGu6kKr+ly
9WdfQu9qWXeuOZNZkeWEgD7YN57hoyBstk6HWpVEl+6QzkphRM8y+VcrfSxS
b3zov5WCDPWyVlPPgMWgJkFPhkMI1cvyzfNQqpzv5Jwu1YAc+PFAN/A53XZC
3CSEBkOa1qbHGQ8EsGIuYPjpzWPLH1qK6w3uT1hu160P1Cirb4DrpyBVrP4e
VqI9R+j2VoA26VWqtHeGDaPuo0r1xAAZgCDbOX5/AYYNY1IRz+txG1UUgk3X
R1xwYJRolfpNhYApzDhBKFVJVGjkItTgWFg73gEsGh7RjaModxpuhtYlEdPq
QUKNaHtYbfki2QGJdLYw03wOr9aOyEZwr8Lyub8a83B5awoM5dXzfSwfrVDI
Zn8IYXQVlRnX6cH2ZeTlpvLRBTYcVzbjkhu7s2DubWw/jJrZ9G6VtzAcepIY
YoJtwi4COA0hakCMq+s+qPLo+tPpEZGZygpl1OuXzCN17A31LyKk8ZM9xuac
DROI0XNY4DU9h5l51pbqj6wQOoXCdIWRtCNFtKcligWYkdbXoh7xJaDU6UvI
L5Agr1EgKeEjrGjwu42pf5RkgoV94GIVXEkoHkeg4eqO+s/7E0lPJsRkcxwk
PgIlt2+1sy+i2uvClSqMYMzGlBOGdZzcDavi5n2mPqBhgh+nFxsao7WXJkQo
VrHaxbAWhXds2ARFo2mJuoRR1sfmj42Sc33883dtI2xWFv/TajfmisCEt5Sy
geTBd3b9hx/cJHsglMDYgN9vDzTVa1+o6XjKnIg4RTfgfrzhumTYpnyflekx
uN/ogKv+WRCuz+Rnn3CNch4nTpSgseaiuV2nk1uMlywZmo4DKO9xqQv/B6fd
Z58iRlHAbmFHLOJi4E3aHlc+tAvMh6egfEeaazzo2ZE6OVZmsyxBMUQnQ83C
74Zi7MEGo6otvIEVvQkjUjNYows152OiuKec1YsX1KW55OdHU5DNHJ+x/LHg
iX4+YU1ln2AVzn7fPgWGepRsXNEx0+bhad3/Gt3qCCYdAp0lCN8ea/kspKPV
pTB4y77sXKWDQZTMP45fFBVwXHOTCfwEM1rxCwRp0PWpGbhiW9m65zCM8JTQ
Vd8FSBO7Zeibwh26HuN3leaKMeKEBk929eYaSo8AH9zMevTlcqGlqx2i7N1R
oFNQ/d+SI5YlMqkoK/JgPgBNlFghjbMlUDVfI2J5iCdRMhZ2hyFh+Drf6CgK
Ts5Qa193GBtDtAdmlM/zcQo/yzc+Sa7S1Z+guRDHm/Hsu8yZuJ0qevv8MDt3
TuJQydTQkxkxVeQGolLtqLPBMxSoGDxFI+aQlvPpS2z2L3tSO/YtvcCRm5k7
rI13G2OhHiI8j/erWrWPLqLiQIMPeKEw1x+Wn9ycIOPo0lej4BTEQui6R3tF
YYrDeF4IU+vGsYqixK7m+SsWAGy0wMWVF2J8bJB0WGgPlCeMILePbKyl/yVC
alH2YUGGNp8bgPmeBvOpzqM32teJkIZWd05Ht84+F9/VsFVZkquxW65Ck0nU
CU0EpNCKpS1QxPgow9QUrrBO+KTYVGpnnwEd+LZxMdLe/r9oyqCsYbC3reN8
rf8p67YonPfFVZ0a8DkH6/Qo1vsVhknon3Bmoj970BQEIf1xWYaWMNCVBr+G
wLO6YySgkwCwrbxtxuX8adl8/YbXJx613NhBG98LUI8lLZJ+GS9fnCJT3HTy
Bj4QM7JPwG8qAGh6Pfh1mFw7gdE1jCnccIfxdFzCbdgabn6TOi0UzinJXX1z
9ipt9h+JZOhSPBfIILVFdT9DGiLoSZoQyxMsE5v32xwYNSl80d3A2dy5nc2Q
XvB1UVAI/YqqvVAdbfgkyD6vPXwvYyZxfyxwuTa4BwYfqSEpskaf3cWIfe39
kKWTaBlMC0vfY/fW/qPoB8Pbo96ZzQ/6bz6ajnCxhGN9xdA0VaeYPfWktmTq
3hYFu/o7JfuPjROpiI6T1BqqM8pK4jvTiMX35NS8jZ78R+iqz4g6FqmAOk70
0wl0ea9VYVlS7KEZsWrqwIP0zgGSlF77fllRPIHdc4pwWhXmMEnnMJVsnaKm
CDwZMUEouxLbLO2p53mT/aKVk+5H8o45cM/ZA8zGU+b7E+1cygq7iNc5/fv1
BqYcfp4Gw+X6FVZepg3cfw2d4MQJ7sllCeWZmXaynkgbIkUXmLZ8qXJ+oUOO
lrIg90kW4oSf6eb1gfFm35NWw6ZEOVgMVcwJBrI9SyctxD9eY+RU0kzaNFG/
xbeiDXYihfMmWlvxvRNp/TA8gCRLqxaNfFgwPMVlvkhQ8Fd8Kpsyj+G1rcgG
xAz90foZegRpQo2bEH+pRnJtzfn8DzZAxgoOCE3Ym9fO3jfJoxuFidlNASSh
tIauIxcEQxkWZZd+Uf2KW0LobEEHyVkVHTNaOQVETDeltb3K3/+QYkFgNWjN
mip9riZtm2EA79MsbDWICPTiZlEg1Sduuw9ujfrPNnqCtO9OTeDXeuyPtmyh
QDrDNkanUJAVdsQ3Y7dwFPdeXrZtc+7Yw51ye8+gAFLbUh/UCpZP19Qz3RSr
gM/DDYXhehMYLus+AGWdElCi7GvvHgE3k2EOhU5kamHnCeGFc8jNBRjSeQCC
yWopgnoKKEMad+W1euT7mbrbnocZZftGp8284OHvRq6Gp66g9Y0joHUORoLv
UGCF5YhP+i8XVI3/dhuluftobuAbsxA28iaBWh50l6wRWRUSngTdrQboM1aK
WfUIxCqdM3c7zUfVTL1brl/poJej+N6/qQ3cZ3WXYvR1e1IEmrPXfCLGdXSg
h8tM6M3CEFNvDS9trTbSFgO4JatxuTHAA/NzeEik1ZovbeE22Qc56QJv/K1d
f1sXWHM9kdlknHGQIuPnXB/3lFbSdv+9XzQEWlxYA+WsrOLM5FIy/Y4hnH5A
2T2L2POh+4HZy/i0utZJ6YLR8hYdsiAs3L7/977Apwb/yLJ5NFar10UFOgLi
2PlBo3pcNNnMa6Oje26yb9vqS8jIhupuPjFCqF2cjnhjv6luzfcT2GhPQbGw
477Lpg50FdA+saw5LozInuYQHEvucTeJe9XsPiNb91RmH+yrSjAABJTOQjQw
G7r/ZAJlinNgumczXc915+2Vjro23SselcLvXfZJcMaC6RFhNP9KfQ1/MOCi
IZ6KuBMQf9B88SFof5OuYXAXiw9eHSkwySTM0hwo4riNihesZYUMDZ0cGjo6
S36NkgahmUPQ5lLIm1kJSGisfjk5DTK0bg7RcOJg5o4OusA4lpIPF+0P6jIA
KvRPagCj1L36upXPD8gOXDWpT2yxlJlN0pGoKmhxPsYKkGTLdB5tgIxq8tET
YBLFMz7/+MVhyV2jEstWDAq/K92VmDXaUwRmLXD9oA8jSnKIMrd/TRZxWFiP
Mu4rOGYCviDdmqQotXjXM1bfjbh1QsQR9E85OKi3IoVHIK4kX2SS1sgjgf3X
bVbkSCd3JRi5Y266zLSJUWNA3+wBN1QqWEVGqdgGLqajmAKsL9m2qnfkMOgM
e7LYq13c4bkixnMsaGYhOlbjKa61+VkgwzI3GQo2jiPBab9NHbxXQ6JM/28D
M3XAgeStlc3v7EIvTvf+LEykk/NYFglNosnz5uWQr7SHWz4NEoN8LfVpbrPA
CsaBNRxFU4tNMefiOeENxuMBHUe1rPk4/7aKWV+Z82dVQqHwzPQFZ6498g0E
osNtsS3QjnGgcCGIlUxbuGH5abvF1UrVT4bIG+dMe5lQgx0+VReGFZbz9syJ
FFS1PZxbAcEAFaw2vFHaX92hcYMX44rxjYwTg+81EyKZltuBr6c7yxqLdZk4
SyrKIVx2vw4lswCmBYNPjWaOwPQxSY4HSh97FwtFZpMpnd5qfteOLAb4+eY6
64Eoa7aaYU6AIu19AzizwqXND/k+N3vE4nt85sfMyE4Qf42z6LGo1ToqVfE5
Jew3y+Ppdq+qC4pAtO+f6i7HOwZ3D+RbC/IBYIXDvnFoEzORtMkkNJ8+cO3O
8SzQrRQd+hui5xRB5qHA8hD+KzOExpgP3AXIKBQSKQ12k7JCsMiNCm2Pe6Gs
c7AxYkMvLt6Va78lR5TO6q5UyDp1TZYJtZFIc93I8fyGUBp2IM5O+fsvvcyu
PiuUJzAMQOfEMUFks25sy3uOxmh4ftY4VJilTc7raiDGOvUoaP+hM+Ut/Xj4
PcZJjuX+ssXstHOVgoX7QdecohvLZTO4j1B6o3Cfjls8Fdgz1Ia8YOgozuHC
F32zn4Klgp3nPguli4WuPtnUHeY6oCLHsRgTGxxx/xy66vi24J+f1diYa2jP
zW6yIT74X2SBPQ/adANmLs90jwoooxv0FLqguMoy24/TItrI57x/Q2sU8RRq
6+j4Fe4TghJDLfflqh/4NnCQLxws+AnEv29CN9ikCj4ME3AVxO/YHn2L72xI
ld1woaHoc+MbMrUisgJniUAw44Y+8E6wLaTWmm695IOO0O9rVQiE4auUkWAo
r+OhGNjQp8/+RWZB87nX1FY5tnA6ZkQ2csATx3NISMy6oZTilrzAwDp5dfAn
9K2qyllbiR0o8dq5GC3cBHDtKz/cYad9iu538Ht/+4RtU3PlWgDISMfe40qY
Q917hFp4enzrhXRSRlosNufmd9WJkiU+rlEhfJXmbWjmx8YpS62TKy/fKKwK
77g6P3yuKZgxi/KftX/v8n6D39YoO/+PhYiuXRTyfdUyzNjmz0rMt8qFc47s
F1Mau7KTsg2/JZjIPljfhNgUcUbsX5NL5b6WHN99fVc7WqWOMvyeP99b9Oeu
Lldx50MW57YLBIbM3PEqrSBOpOEAAXCAXQpoJGkvi1MpQ+YFOzbPDyiUCpZA
F8GJ70UNLJ1ZXGXTR0/jJDdSjyhPeKydVVJUXJrvx/MmanIg0fwjGDKRab05
RujxAR5Eso+4q5H55G2p54F3Dq0k0uIG2I7xkd6uWFIHmRFh7f3aiCNh43iz
Mk29yU5mB6FpFF8HyTxCLqIzQonSBmhCxGpjM64Z2snTRvuol6K4hNWdojEi
ta1iMIB8nIut8cXPyQJIxfN+wjH6XIkX5blWKTsJvLDvs4R1BTILpTwATO3R
Setvk/F/sAL4GSUhUZE9HDxMjITfNtw7H/zfOgp8vN/hZgZtjW1OzmVoQtOz
1lFD5D0WTtKHXP8+o5I0uRNaJKNVgYkmNgAqSas1czok81vhGtns3V1KEBv2
QjCCuGN5Hl14MoDr2W8Ak8Qx9c4ICwCmODKbXk5j/OY5t3QY6s+ThB0WOcQg
VNwjdlnXeoO31fB1NpnM2sLBUNSQ8rwBcgnnHq775pYImXmRFh8UWk0R6P0c
UX/e7OLTklwXrLXKi5jhJqvRSqvLLj3KZ+lJPlolzTR77IfalckaOkQYBSgN
obDY/MYMh3pTDD+zP+RsNRcD+s4SRGGzn8cBsXJB/Sxs2HW+oZFrIbzKTX/W
oBG98x758i6n5VRt/8qhBaYIs56k+zbcP2AXrIyM5VWLpg8eavCAY/AFnyjf
Z56JK15e1ebaJnCRdIGfxPUfNFn48GPYC1HkiAnNQJLsn9+27sddJFByA0Fe
W8NjKJvGCH/t0zoxsIt28vqkTVxPstpbTJMpa7bG3LRwez4lOMHg7lEC6OgF
RgE9jZJ49616Tz7K7XbiurZygUT43MVt9Wpo5UDUdn/qL2FG2RVFvYMpscMV
Avi/78x43RZG5rYIjbst+2506lFqhn/7LRxUMikCLrU4p4nkIQNP7yiO4UW2
tItrXeqV6pyLnbShNWfa9C5IkUCHs0/tzpN7ajGWVyLcdvh/PmNN1xim+rRP
H3G2fQfcO9Lnw6QqL+YTAhghElCz2tS98aFfVdBMN9BvFkLOg2l+CpOmIT/F
h3vjxJjfwhX/duWJwqzocTqSPEwIR65OQT+Iw4LY5PbQYe1S+HdFdcWElSnE
WOLYmgaULOTrP3U5wMnsApQYoa/qI5v2jfbN0l12eCkMwh5rqEToPmZXxpry
1J/fXSyFq/1CJuxflgN/PkeU7jnwp78thiKZeK77HG/meSNDqQrPt2Nzrg2l
DrmQh5+bxD/VbAOw4HhKccCdz2+nLEuhkr7TqVuHk/xL3Al2pRHOtGyabiF4
xS5SnoYWfh3eoJukeNJvDXWnCo+5C2x1ERrBDZT34OYpqqOQ7yS8AbWuHQIq
buFmmAPUMBRIz7CPRuGFkbQpUoRSmLHggjjSbazet6XwGWgkqIqmZjhsSDKt
ZX00D8eGYzpeW9kkdLaYVEi2aLN4VRgTsEAPAI0CarJJreOz7USovTzXybAn
ExxaaHLOJ+J0Sc6jhRSCJx/5/kB5cfxHMUYyPrOaabjUrgJZrC/dOe4nQ8Gr
MF+6hRr2Gq/ZyFGA5p0Qo1XZHoq9jU4prt15kc6RArdMjzfHjUhMs1bbdXeW
4sSCpZXSU4RViCW8NipHDT3LtlX0EZbtEPX8L6UJhqdF+3SzN7ejQFF8x0zD
15rX8Oe6egH+QRzbjOOk0c+fOcfsUn5m/sh6BmeYMdD/zLx6lHgsTXi9zQHH
ntVT7cI/nZxzk5LwzUidpsLVsOlqsTCecImhGygkCnrG25MRKeoril7EprPy
qkzRz1+kfxiPUwy6zKh6d6il/+jlZRCUgVxDnM8f9XzHNaVc6hUsbzjPgfoX
Pw3a4LAKUXuMGwqTxoTgiTU/A9ZmfBdXmo8Gjfl4soTXhFY3RPlXn9+53m8M
BizlowrltAVJrP9IcZ+cDj5efy2lOtn51kVeKsSqX7+u9eRqY3Bj94FTXLjc
EHqb1ByhUXJGFuUgQVfV5UbDu8lQ8Zuahbn2RXS0Lw75povSS6p04psDX7hP
Eamv1B21zRw82EjmOVh0x/wWKN7uBsuSyVGm1Ic+IHNx0YgDB8conuSiKE5t
Xg22Egc+2zXOo5U4+voS4wRYAPKlve5uP8KdxeAjBIeetAyao006rqBKOr/1
99aW0hwDa5hnfRxmBBEpGPaVt7oQ/j0ivRInlkyFIhtoB6SJ8K/Gt3bCf/Mc
XMnaroyPJ+IBTYOyBBEjI5qCE+mdHB63ak/h1gQFYsSlylrYT1QJGY55P8xb
u4WMR3O/Sfr2EzK9rpwVbzXjsOn91Vcam5kHro1F6Nxgq6vYr81cqtsr6z1B
LYI6vE7QWtlE8evBM4rrHwM+2Pny8FGd1o0e84/1n5Zd8lVvxoG5NxidBPhv
UNeOC1ZxhOj1J7iDwmKQE7x7jCnQeQqKBd4OSt7x4PEVSDPO5G99rmIWRrtt
3q0jOvvkKBZXGt3c77EDFo9AiDSIUYtkN0zqk3q1SnB+MBJKPARwX8pt6R35
6yg5QwMm6IvoRFyYcCsv7UJaBTeoy91zRJCfiTjsfMvFIBms4IThFaVN5HxZ
gq8y4KNUv+Rxg7jdPF6upQ9eS+/qwGSnNdLT4Yhl7jWoAUZ+3ZCC4RLPN8oR
GvMC5pyhkS4KdYcncyqNUPnyzMXXUQ6DWyR/ZMwhdp2HOpY5gyxK7D/1e7od
1tODdBVRi5Zsr3EruXEDYTPNBJbGP0afbpF6SbWPQOE3IMv2AeBG02Dse779
+iWZrqF6ezD+JOv4Ao6zUw0hUXr3w5kTSeCxf0KdbBUXA9wOsLVhNY35A63r
4oDq4HXyM1/HS9u96YphsuDj40y7TgqL7He9ghFohgU+yKC5M/FeziFUqSGI
BdZjUJmzQz+8UFWYPhiykLefPmCr0NKSDueArn4JfUiKsgvN1E0c7zuiRTZr
Ezz7mey+VpgzFy2h/zgkOYGO9OJlzBJbqmiUSuy78UyahlgdaJL4xM/W7Wnw
+U11sdu2r7DWxiKrWMm2Tdxe7KBVnIGZ7GWHsYx7BPOt5SQGX5dYgszwT5+o
ACaa9FdQzZSXdzPh2uJ4ZV70rDPJK/vRSjOisI1pKiiYZeCeyvaY0zZz1PTH
Eaoqxzcq79SS2OY8vLDJ9WW4/llg8od7T3no3IGFmVV/VQRjtlhJYRvgbHRI
inXwOouCcs9qFE8Io8XWJOqGXiMmFiPNMCMQW1PuZpsktmQ2FXE2LZn+HLKL
IHUaehftHIztJcwW31L5krNYOJOsT2ILfGlfIm7N6Uat0kHy/9QS1wlbn/Qb
8OGl/3TNfQZcB56WiAkk2+moZKVWTzmxy6JJZkpBQJ8Lrdl22XUJxy0NQRqL
cBYaG24acSv6yW6E+tzpIelzw1d/rRj7VnpzUaIzzKhLzffN4OTS5LrDKyKG
cLr0mBD0puclf2lJjhhOfW9/JSdgcE0phmDu1iW5buWjLaKK3zSdomba0szJ
qnv9wT/YzztKzAL01FkmpEmtf67US5IB+fEunvZJeZumCouhw2d0H8dg0w1U
DlZk3HN4LlA3z71Cdf/bv4IcO2uKnsyqHkdiUI/uZ94PUxTBbkh09YLtqRtd
f+DqE0zUq4Q0KRxtAP4uTNzOEeF7+bUOSd2hmKTbS28hcwnBhPRdx1N8o+2V
5gsvA2wLfT0ovudB8fOwM03Xwpwy7PZu1dn4SFwtgbNVTDEpt0KRx2NBtNo1
SnMj9hFnQ+pygHrfJlRS/rZ7cWc3kHrOm4b47J1aNltj0+O6d4vBc3KQoQG5
YyxlKSVJqan2EX/LiwGRUW3e5fszz92G+y5YtKHd1QpDH/FEnauO+GaBVhO+
tXEiuvLEkKeidEHk5tbhBoWXVWMUzNz0KjEG3juf0/zNtF6TSRw2g3u3h2ND
jvbKMG70m6hDm/1YMkQWI9UIcujK5F70I4N9V6lBfNgQBT2bCR4bbhpjhU3/
FZ78pLE93992kVX5azQqg4dRH5+2t1HAwiIe5S1BXyjbiH+B4TOvn8Et06rv
+B0iXLzUsy+DnWXv1xX5tyumcgC/i9GJ/MwVgsrNdGkw5J2G4gOEl0cUQ2DG
r7FjWHNbfOwiMEwGNCwoXxZdtQdjOOj0iE3YyuWrKZFp39XpNlDOBZQpnnOZ
6EjLRW6xtncR01/kYCIVKOpSbLF/435IIMgIQOmZHEcUUTdHcPXE5fZZTuAk
VRoDDOQMhBFRMGGiRZx5JcOA4Rvc5h0heatS1G58acwcC3dw5s7RjPHPo36L
kTENSM4dxyA2nNChJ5acEPS8tmGgdta9/fh9Y3OCXLKjrcmqiCAhp8TgNfMX
tclq0MXEuWf1J/M5YDKaIAeKRyCR2Bi0Y279LofqoyGL9BMrcbSjnqbfzCAA
3S9f7ZmsrejOHWbtOwNcZ0DjqCtTXPh7D2e852gjREQqYn14PliCOm0MJCO8
3zILg00MA7XMmKqIjphrUFmQj9zdkomgvMU8NLEAhDiFrAa+wVHKC++f9Da1
NMc9WVBc8PddlpNaDXx0nvpfrs0jvJ5EiknJbybpg3Ms6LxazBD/ZkhVzvPJ
k1MOuRgqoWNl/v7AlUv04AD5JSXCM2EeIKb3GDcjzDHdR9voPZuxsVZpJPzq
hdEmsEHC6xCy7J7T3kHU4eAmJUZEdB1iQ3lezPj7KBwa6y4TGI22c/jWSFCG
3MBfEX+rSxA0NeEcHAOzVen8EKPKdoWLY3U0XzG5FzCk6FS3sEnkCJgAGm+j
LobmhPeb8m/PCpRNWzDe1uIAtIrLbOKFJCfNbY/FydFheyyQvW+Xf26hy6pu
43nvswtRnbFIPwAgskIXyXWZkwnmZ9N8L9bGVFLsCms7IHT3o6j6/jzwnvT/
q+kmalvpS/pHdLNZvBTKVNBGRxEPS78KiAk/wntQ/MDi4HRuwp0wVqIKOKWY
gy46IvoHaT7bl8NyoKBSRZESLIIb6u3QLvJkzzVxmSFocs5nzulL+q8UOnqm
E+/Q6e/cI/Ju6WPLWLEZRRIR/k3yQOt3VbEMgJ1tCUyLpx7wKtf1ZtW5h6oW
DiMMVp39BP/DyIcfxaPRHNEDMx2P9+2f4uB6B8TtDxobrekB7Ff7KVro5iBk
jtL8mZ+VxEg2MMTRSmDCx1m+5lkqricFwRg32u49Q565ld7lBRp5Lj+2tHkV
ngHBtdZ6xeN6gx1OkZwAXDEpjCOMQWWPDRV1Wlom9Sr+rhAqcmq9F7MaWL/4
PHCT6eLitZtH4Yhv2YSsPIEJxyp+YkCoEXKXeOCD641p1ag2lM6sRcMV+jEp
BtE1pNLf1zfMo6q7p26Q5resaeNPGyr8lxddZZdU/gurJNXc84oz1vBBWExv
7HKxQqFM9QvCVbphW+oFMSB9VcmVVD5qZdhuMr5GN2KAp5q6RQXOnbKOUToI
6aLoryC6A8CkVugIG0vqcDKdx0w+MWivU+aEodTq6Ui355fae35L3jT2kJF4
hZl3kCDmHL5I7hweFUPaRw/eqor7hnOjbQJaM9vkmB8wAdTfbZY5ydPUK+CF
SFM92IZjFVIOLhlyqIjnG0qxwZnL7u0eyfpvkOLsoTkK/4THOHm0IQ8CHl9L
ow5SMYuPVcQ2XnTsEu7OTCPv//7TP1KTszEIo6tN2Uv3ILk3BGaF3l8T5LD2
84SXPib4/BTotQ8+gmH4jMfQi+aebYAun7xIwdUwX1n9EKN0wbUtWaTQHrFP
f7mg0pTEPb3UmOwSMaemMMWI4qEOvN86Ed5MbZjfEKhGjwOH71mzc55a/NG7
A9g9uVpCKh0yyYEQfyE2LOQh43ac2Q+si6v+3ambX+cwOHsdbfDldZJVsV3c
8r3+lUPFX2d6zDp6gUanIghUDu8tMb2GQ6T157ArlTV8VfoQg9vmSc6zOveM
Q7eawhlgA/X3k9WFGFTfsxL+HlYDwDIaU5YEC2EtSVIkqPF9/yy0k6jbHcny
K1uc36msIvbvS+l1NZn/yykb5pLAYRrsBHT6vvEX9NMhixqLXIkrkYrYRZGp
oqeo1GTCsibulrgYGbqSe0FQGShHrlSANGJLAXEcWO6OVmk9G/XP/10VbHhs
+MKFiH4LZ3WejdoH2hPwT/TbIBWyGeaX87LTop7tNi8hREvbMBdRYHekLdke
kK2xYJXIEn0kjel73QEBKpdIZz2GDnCPIhCq8B8VYnFBkZrPhFx1qZMns04g
0DIOitEJbW5FwM1Pxj1UK5DdiV2VwO3P0LCFAsMY4Hze7sKRna7JITaFJG62
G5TLoy1e53jwsr1B/XYiIxdu7M4KRn/+sSSR/0x3asQvruiWAaS/inV2x3TF
TrW8aD2MPdptOaY6FgQfwTO8WwBOXooz8esxIWL4+Cri3g0A0Vn056s3v+Cn
JB9BV6VkcdfCZ7mUsMCO50viyBMSsurRfjZLl5SPYJ/72feYgpJi4WtuZ6ji
jjzqTe/fwHYqnh+5IBXeftj/f4HcXeCWvDvirqAvQGLN3Gir1jYgkmFgrkXV
T/SBPMbY8dGMJo2N/qCey9bq4IIf5Pl2IWiwdf7VHhAsdMRdso/waB5wIgjw
Fawyq5Lh0FC5HBdG9gLTrCx7T8AQsiJ6XGknGsZfh/DACavAeq8+Z5jYEhDz
7YzwTGzORa3vYM5Gut3V4fp0g+xjLGFIj6mJM47eA69H/QJXfb/AN390pdgt
QP5eGZPyfog8musdH34vPZ3vr+hHz5budvh4mSdinLEJliZQdd7FyAYgMus1
4J77KsMF1RI8lOsjIBgqYb2OLmCy7ICp3L5WknDWKFWTZOMcPHss7U8B4pfF
58ak6NzYP5t2/ZGcQl4ua3oG7KyDtEczPlERu1VdwpyWk4MvnCi1INO2qFHA
LXPyMuF/B5IsK4L/0bv8UyQJ1A54LH7FFjE07HK64KFn6roNXL8UKUIcTC6r
eisSIuWYhHMVruHfGO7vD/50Utebza9Ut5Rdfwmd0ggtHEuMb5Fjx4H8BdB3
KyRopQDNWrGkigeWu+11hnwVeJW4uxM8ZgJEovRhltVG+cwi8b3mBd4p4mes
aDNORpcsxJOBK7kfkSeOh8W+dX9DMxup9rpNz+Ob6/X5OSbrIZ2gUdGlIZ7p
8JiOUZJ7pvrVb/35hHSPiXFEubOJaE7OTfb19OKV2E46E7Umg5kXf+g7It8R
S68BjTR0jxNjZucWRMfrDXM7FiZ1XD0RKmJl9NVaQ6JiNwSt7KP3nFCpjdEG
AFsREwE00jZXUNfPE7j7/efGyzQN1zMCDWanR4urNr5WCUTCt0v0E5aqeQaF
SaQinLnIE/Pf06+qoL+++tNIAnLbCxQUdVTV+dawdXYKxzj5gjnXvN2CVxT/
AYj3mCpqAjJ7lt46OF8QdQHcm90s2aMoZqQHqEiRP+VyazCyGe1WvvGiERZJ
WKla1TZxZQJx1Tzl69mD4XZ8oFWvzJMzf/cC4Zn7K9sHBSubVotKsICdGF8h
FFslsJh3UPUq8YA5Z7ag9B680pht7eUT9tFCWFXGt6RGEfdRkSVABID/av7g
kbcbNMQ1AUdvoYCu/vfZqY8BmAqAQGBA9drMj7XrCSgG8ksTVREvwmAx50UL
/ItpaEmIjLQJBck/RCYLtSZf2LjoUWhHPjjtBxMr+ZxmshsFHQKctPX6Pk7C
JkOiRsbStge9MX4Ta+3R6QeAA3n8Kci/MqZ8QUku42l7YQJN+pcFF/SM/LXC
gyLho/C6rQfQHOKNMAUuKmyuVLnPEW00bPIDjnqMgOydfTGIKTHKikhZk3LO
nxxzJ38pYEHzzBJN9fC2FEP/KagJXG19xhaKgDaZ8SQt0Cb0zpkbNnOn/V6S
lc/Gtr/colarnviu5sj9f8mKUJro5aDYYxAR10Lwaydipi1hthQwSc0OH3DQ
31UVWUWujU++oGK4YP4SAoDJVkPA6aP2X5bwHRncB3zV3LXEsmvNGQc+iEwD
Rk9d79lGhD/yuWEzBlVr3+AFVkol/19ieUqGKs4v77xEwcMKT1MxA3je+CSZ
WOauXKt0l0YU8cloQhghmeWR/PCB2OHJ+tVXNFt71IMUTi+UDa7PdDhuh9tn
L2ghOZf71CkCk0OMR7Ukvre6Scfa714hrwKfDrjDxlWeIDZEPl0rzsUtJQFh
j/HT8MR29m6uelb8QfUZdkGudgAEjyniLvjsXDEzCMShI4ckLKxOliukxq1o
/5J+KJxmh1tZnEl3wkng8gSQ/G1cUfWTVjW4ETXe22b8eTJSNc9j0/Vye2rE
/fITnaz02GLZbEcuSkeOMs9WLgTz6BEa8sy1L0WynkOS/WiTxB+prYuJ/S1r
WvZl9+0hKfbt1r4S7KAKdUmvpCyicEQXbtdyyqYyYkp44YYX40Nr4OgyqIsG
Xbc0LCMmQHkK25Srcfgn1HlkNHeHYVWMf4mXEhBSX1o4VNTTHJTHifM+WQnD
ePRg3gCQXb4soK06j6VtE1EpkVAwNXMso/UiCfCV9gztOmfn1ssSrEZ/2gtX
evl/OjlBoXbkZb23yoQy+0dv7EYJS5wqxUObs4CBIXKE1q12tFY+JFr2AmLs
DV4EPXlNEjGT7zpUWsAyz6PtaYxKP6rc+Mq/RZsKXydAFtb7aTtFpyTtRRyq
E0CVfQGF30AfOpD3KOSVNR3wNdBFXfxNQq6AAfWfJ4urztelRZzwZCJ8fMC4
FpcPiYFi0Vl7px0PRBvjAqBDPMyh+F5HEF7dLwHmSTLtQM/GiLWG5sqrFQRR
X6xnhlkkXYeOqxf7teWGts7mLyaW4ySVntiLzTyOGmWqCepKWxUpLhwx1CMQ
f3AqNj0Zld4l9GvwLwkDHMMoj4xoGyM7GJ6e0DSjowhznCQ4nZ2nTBB2ljBu
K8JYWpM495ps7QCfz3nHM06D2BxHbOQ+HMqZFGxo2+y1McNj2NKBMdMK5UoY
WADgAYRL9E4kDcSguGzuwWyoiqvjWrqj9jwUovq4ZaKtT2wH+Q0aRwalBhpI
qYkYBhjJ/P5axE3LZ9Tn6HLzgcpyW0HDC9io3M9itgI5WQcDk0SyjvwrnRxZ
CFAonUeW5ATJuaRTDMrccCYlSlSXwnL5piwbnbRQqyN+XMUJlYbLLx65eO1T
s+3jd1vqmEYXvIJ59WDa50LfNDOA2HeOpiyMonQE1Cv6y3fRgeUHeuOzE+ZK
jb9KuIz5pNTth5jmmQ1OD0Zk5k8sTocilZ9NmZ3m8Dc28vKWP/6Y5CmSx6ip
HCVrg4v+oJy8mFMUEbVimRXaH+EdEMHT+BCfHq2W5ifOdkLLrzjeqddxBXQh
mzh3eU0OfzX5GPCUANRvLWaLWAwXQ7h8ZN6Zo2b0dRNKwGcotn+v4wYCyqJD
jCWGfzrTklHEH3X94z5FFltEYD9LxHwA+SFrP+Dh0NtuAb55Pjwi3SxKXQMJ
z0P/F1cr79XblJwsQWzGPwbaTgyO15aYseofpR10250kSVzaeH6epY6QFNuS
ajzaiVQKJOzVqXQT7ZEJNbpTHsP7rBt+X++JDlt/6jg2D2rGY3u8DDUWtfEs
IosyK6HcFIUMepdxT1tv+xNoQA3ef5iVyxHQP/bpI1Xm+DqRdrRfOVHzkp4w
3ifHCGiEOFk1BDZ48s+6NnoXY6n6GKpmL8/pjJ0xDQQS8rHxh+DmIuVAeuZ0
zq+w8wgwwuchVmrGJiWuqZH2JJv9qEfMwhnvdWTwwI0HPQqbozU7WM2K86wb
zJyhnn0KAZBwOYWYr3zUy3zO4asH1vKdc+M9BRDXj2Mhv01ckJTrMBN6VBog
sbN7ClMbLQcif1iMk/yrSjmI/wm8Q1/3lXpKfBWxiovv7LYs2qHrtu7r8So2
VxhNG9y5AQtDA0NHSK40yyhjtEvy/BNPVeiu61muItKn6A5yOObJBFlUKk+c
uvNQaWW3EWPKrTsI2FAIb3wEXhNVsogc3UstMH2SE+/1TPLWgl2wh46tRoDq
UYXceiCuZdW5JcYoHo3xUz6g247j6JfBMWo0Egc2H3NvKx5jU9XXS72Gm31+
6eWOEIz0PnLqLwbrI8K/ba7vwLJ+TfQY+paCC9jzIdjOu0o2oeKJDmYLVX97
n4OpXUZJi/tzP2jKrNcnlx5OMNpDTku+z5jR3rih/8t/PpTZss/pvoaShlVz
djjilva3NxR4M0komY0v5zUZMUsjxOaw8Vjn5DEav9scRGi+TwOcNPBFQamS
2PPnalOo81agZK4J2tchCGh4OyQxX5rYGL19M+qHzcOzc3A7ghoyRnvec6bu
XsQ95h1EsSVhoTUAK1HnLlA2zQKSz5KcQFvxmqDjNm0GHcsZ4PRko0rCPQVj
A2MJoK/anYHE6iFg7X2diV3WKbjI/GiWYDJRlRZDYX8XR8thHaNsySgWmdZ5
hgahlHZN/e7G1l9gBWnf/Smruffcago47dFApSjaU/H+B/Zhl7zysE5d4XvQ
S47ritfxvcNfD14UGp94M04w5e3bQthIzOiG96hcIRAfZnjuR8MS3l6nTsTi
jqw6vwNIU1+iH2JR83oyhKoHJZc2A/Wr/fQwMBu7ZCbFqnFAQVsF+1H5WzNP
VakrT9zL03N8wGZmtiLZmVt1O4GuJTAaU5FvUMprJtQ0+zP5Jm2mVaC/J4V1
E1Iclc3H9z79Q0ScHey9FRl2YIrtedeAug2i2yYoDGONGfr6suKTRi7A2xCy
98xP3a9c0bYX1WtBsyVBYYSoktAdRqaNTsAKyuyTZb5ejdV0WvEZFz3tsOtq
Oda9EQiAZVhMl5pCFgZO43joYnQU4dgXQdKZCbVjsdGevxuIuf22GPKWqGv6
Jl7F3db9fUxW2/l4rlvgBxtd8IC0m4DmcJpqui6XlCFMZnPaPdfPPibKTBop
IZ8LdPJQkFdKtI2I6RT93+ckC0snnA2OS7A4RewYQ/kyRJvc4LRVy58wjDil
9aWOwdGcRP4mm6U5ULu1FqTjPDKB9omlSfd1SKdVwg5R5yI6zVcLD6r1qVnW
fLr0TYFarD4rdtNfXBT/AYT6h5dAWb0sKEbeo5Il70VEOIJsbrqcSY9g7TVc
9c79kBiP/fZyVHRZq4Fq5Ze5K132L1tHAw19SmiBoDgGX3ZH+gAmHG/5xiz5
llpAi4YYQoz9IgsHQDqIOam60AIrRBNBIk+xO8J7zGGzEeQtqvEIBu7hOCn3
LwCiIOQePe/oN2c3DTp/ypKInKYpZHfNOOLYZkOOPeHdoMi3MwqB8PqX4RIU
LEJqLlJskXE59WMYYFbhiCdYmYuL5JhTmVRl4VES0u6kI/4D1utC5UyovB4W
Xt68LtCp7eJ3GMPWkxXvMLqhAzHZySIQ6fQNjqisU9bxxMuhtLvu5lMK5ubH
rem4yY5bmrwL0xJoZSlBGlJuwzdWcnGgqTQUya3OCWLlnXYM/F5Y5EiivXmI
p3y3M+o4JHhOilVbx5d5qsJFeaQoqu75+uakqF5yeHVgkYIxbx5trUSAA6+U
FSZZ/95yCKnCioZ955Zw4F6TxkDhIurnG8G0VL4LLF1MENtpQWmk5p0upd9r
8/Tfu7pGMxFE/gwIchNEo5TShtgt3orkXgqMprRjGQ3o1V+OQa2Q1mjLBBEe
cfxjAycJMtToZbBKDRBNJDcUc7SIy2c/3A4iQBUhBk0WFHzZKasgg1pU7mII
OHD41GPBZ/3alxX9edDAaNfeLjiXnNRLnUfS+ORJp2FhzcwAaGk2V40zCHHL
A9YkFEQ3f/PNM2EPR6ZXfXb+vvfHn3ZC7aB4nvyieDvxWWjFNOGt5gXkaLPe
/y1/OQDqTKOqaFBAu1cydbn0lDHwdXlkBAP3/gmIb5ydFN+a+V2rUwKAKgB/
2vNpn7tMYDrtXESlF/RZHNxESGvvRwemzRbFovQCQwi3Jpe85YQNDuTho/UF
dsYXpnNIVcN/7u6MreDgEyJsreJXlODK9a2yQA13ZUjiPRallrljAWzpDUh3
l9Na1uUFLOh3ciWRcOXUf7GG1xtbb0QmM0clQAsHjxJ1YeXP0LxVNVysWOGF
VplU8v3LECq7pUzSyF8slEk4mBUwghmYopMDpXotkNvByQ7ebiowgVCav39c
S/4LLNylW37R1Gl6NQR0nf5v9NOXtcjiBQWv4xzbLWKP+C8QnqKEf/DQg3sl
197JwEv4bqi8uqoKPYqY64R/2cpcaJ1aelnxTvjONAyFRp5RJVaPIjaURRnB
ZWXxduOEW2pNJuZK2shyxwX7mBDbPEWL61S/0ANVzCWiaIuQqfhKILx+ML6I
uLE4P4STgckS0AaPpBSLHHq0da2M51THxWMWObsavwTfRja2O0wk0M0Lktzk
P4PMwwnR6Qj4Ck8UyXGWIDYc9dAzMj4fY7cxg1qUxeDoERNsIRXD8LPDG9UL
8nFzE45O4HloHRV5VkCUUilZL/YPjrTr+BMsKaku9ReHtl+sYcPayUDWF+EQ
/FeDqx4kB4xUMEo+1BMuuhdEAb5VqTLzbMVCR6yLp0MJdPMBoEvzNSeqBCbu
tbSwWg+jYvgSjzV7veDeay6lGgNoYV0UP3Hl53jI+B89Hu67gioyQ+TzzMDv
2Z6Y8HL7ODvd2tFVbBHRYqcMEwf6w/ZU33DKWhavNsMN1nYhh82zv8XYC/PB
KsXhzl3h+IZQQfn7zu8SUonzNTnari504yVZxP/c1c3+62wZtYyBnxBnXXAq
WZN3SGh7fuu2C2wA+ZD5U8pfLs+ojo7ySICo15+hhGBcBlsYbeS13quzDU/U
b6p9CTROnPCvH/MBMiOyC2BGvarn8Kivip4x+WKuvzXcqsACRl5BAFHyU3KV
D2tyKu9w1oaBkFP+yZKyxV1FR5rvkpq3tbdDo7kwcf2CrjJmYY0i81XiQysT
/CUGFTXbA0Ctc7KDGfifyuzKYACoNEYAxHCRxuHKhWOYU+SVhBULBy67oIUF
guBvrAzP6G2qKPx9rzpAOjdSluo6ZWvf2rF2ARChJBNXr8Q57U5OJAoVx40k
Oju/Rx7ZJagSuAdsQPlnDZbj9IlJOxYq8qnBjvVks8O7Pe8mS5AhtkeB/71W
5DNV+9GXjEhW0OhDe+8ktM2LfxY1rAATW3zZBaHfwvq9rsD0MP31mdbocjaY
rZjUN7TsgmqT49+Z6k6PLcHhtOvACPlsax/A3toQW3SKj5r1TucF1nSZQG4g
FC+IVL6RGY2a/dcldH3kQoZxDPRH5RCXvJIyGLqqDSCcwMV87t2SNEbWg1aF
iF4lMMTgLN8nW63Y0z/j3fyGm7qaVyRabvnBy+3lXzn6jFGERymVpTljvI0o
98/vezPruo7jzWSklSSgkj97D1qsbwb7Slw/SN9iyoHuIkA20hqGcaxP89z/
j5oTSFqJ/hkqxhC+peAhYDfbIReZq/yjvf05PvBXgV3SZ2dLNXS0ZBJvm0GG
vK+qZqz+tAxUbWj8K35DLuVMkV2N4Rt/jAbv9PpmS1AD9kmfzXRDwOOB61PE
zrxsgumBLBTuCwT+52ZIaGlWC8KZvLBZz+HTLF6ARj5uTCxgsejm6AUYy9pt
5P67OKTuflgfIHoMKwANq3VtJYGNXu0NcqumPC7Dry2eaYqubp+pfwLWEE8I
fbJKfqBxnSwz3OziPkPxSh2P5YDceMz362wVhGf80hRJkHoovS/0VlpQspmW
Ytg1PLRcVae7aOuM5XHikx7xhl1bl3cPUab88MbKqn42sLzT6VmCzWR6Db+S
bpvN6zUO3DntiO3rAgQZg4h8jaPL/EGHRk3SXbo0IOmLpTR7cOcYeON50FQB
1U+QSRBWHEAzzVWvoVhWilus2D3h/vjCvWfX+O7FDBR6WpiOhfsfdidpYgH/
365a+J+iOPP577NlIRZkOB0IAX3b9oqnd/e9YVkQSRoGMAqAYCbwqj4aqc0g
OW0qFGsGoBfRRqMmdGaFj6ndVr1nK/ouBEuvO+UuwixmdQJ+uh9wkfsNj6ZL
GGtqhztomQxFhzhjUEL9QUTImCea9OSHx0UEe1CTJZAg8niB+S+eJOlfImyo
r7wX9xbnCLyFPZTrZUygotWmIOgdryQyzvLTassTVjVwmPBCd+t6nGo+MGIu
8Bmgb972pZ4Fio01EiEgqVcxaZM+CG7290OQqL6lppd58RMj5StUwYkuzF5k
A57V+fGAuXTdzeAtnThlnazsUu9SQcnSzFrYNcgMDrtf+pLkKIpKp4lVEO30
XRKran7GOBt5eeS1Xwth1CiSoSp+uFOi+tTyCIN+cg9O/GFPKzBE0L3po9eC
nUqxbTLzDuIDk8Qqn06QTSO7GCO1eohUChA4Upg6VgGIribaz8noWplMGbkT
cRWnppfwAozmym0OnVJ+ZjUXw5OV/nnV4FrOaEXXfJ2cEbL0Hp0afcluhpJF
4Ply+R2q+61fTQOeo9eMlmOM+5fU6mmDK97AKbqglRgH/mZMiDmXsUQq8Cua
jUnY59n56ebJvHLIBoMYPy0gdM2Ub43eQ4MkBhiyQjBRFyqpWWpvnQjgk+2r
FI6Ovwt0qHbV6R4CQ7K31+Of02+PncRPRWR2IXESkslUWV7Yy+LN2Qpa7Yw2
7k+TMO4sXT+CWMaLWIh5d3/xpPN3aEOoBKuwb66kCLAEobeQWEkOkXi1fHy7
F1Zu+5dkdZyPDXeVA6f4+99TV8amHy4FFch5obm/y2ut+k4wbCO09j4zlRKc
t+Pcf0KDFJgem4+xhOp/OmCZhiQXzGetvAPymAR7VWZMl+2NmEaulopsaQ6b
3V+eq3KaAyaTIdv+ovmMU9Oy2qX96/w3qjBzswHG8k9HCvvhJ4kudwa5Vf7M
9XxLVC/H8N+5JWahQv6y/uwi93eWb/qE9JEII9szLGR/lwBYs5Vhgq+3Gu1j
oxncQaGngOt2jquIqWUzEunSsJZJ2kXNw7XspNl6u1WXoGLDMIxB8ky9tTq0
w6Iqj0lZSUB0OL7TAuqjF5mH7qHMbPZ4sAF43KMEWJWtk8mOu/uLKSUsTeRb
r4mgmnqve1sowOPyRFncLk5rFmlaN+XGRL/M52y0vYWbYgyYHmdJFKXnbFhF
ylcByFHHRdx3iXyKSZKS9/AoJ4s9AjKXtq9gIp7HF9fNWMpQkdjQjCdc5U7w
mhucErQlUtVTTB18j5GTpAL3rEvpJ6o93kpQjSuhYWJbElC5a9GOwTHUiuoD
+HaHaPXDqFZKc1i8hbGXUf8hSWALN5wWwFBKtoTYROVH3H6etrJKUaKFukje
fiyWEF2UqqZqL/HfuyuCdk7vSkHVebhq+B4mf3CQsIiGjrrZffZwe1UImbPJ
yifrexiVHfwJVskYhEEgghzUdFCO4vWE2FEgUyeL62PrOTqsaVG7P+595zSa
Xr4X8fk2Pbymljl+cXVCq3iM8JS9mAbhhcJCxW2Ki+zcRXqYnDGV/CuVhtaC
c08ZqssaP6yUmBsigsw5u55JtbLa7EdcUXH/w8LfQ96LHlxoHWfINkv9FHYv
ForAR5dcI8uOZ8bIdcrQjOXcpfAye3LtRwZpHB2/LzEwuQFMUuH4HP6Zpivi
2E2E5t72riLlxwU5dRv40U8rFog9if/rxQsj7wMuc24uWOVZUZRWVhG+wi3N
7S4XSIvqvEy2mkSJaU72hmmbgIzIWcACmA1UhaKMbBFhFy64AZcbBOvO/7mE
Zyr65MXty8+PyIqAaWflU1wcyZjB2Y3nNqCfyEmU2qGWAsFb6VOrY4OmfcZr
nBsa44oFd2n4R5Tf9XJO4jaGxfulw8YIJvfKA/NrtjxVHD/EFt/6vHEoi/sl
YdlZC5xDQD4QziaA2QR0VcBA/0GGV5CL9vF5nq8Oc4gvrIHcZJeTsBc7gv/m
u/d0T7/oNARzZLZfYOV3y/FlhaR/xdXPPNYQUU4xagpPetuhB7NV5HusjKPk
1/noIsDxMNNpoXpvgnWSmIHUiZLrYLDDqh6TCldxClZUN2Deva+m+/BlLGYU
/PqnZtRMuaDZaZPuJC4PGCeGrVN4s9qbxmJhTlO3US9vF/nXesfPg0b7tiOR
qhWnuwPh8ibGBdpJVkKd+QfAgkyPsL/hB/2IeCm7BmKPIKRt+vaBAYTyBTcg
CnKGGcKJWo2QGboVrnCIR8fX3RxMrSma8hRsD0OEnfvkKLyWwo0jZnE+KWmn
2BGCmf5E2MdOjr4PRPtOkZQ0nyK3n6dIV7HyEda2zc368f8cvQ6D0HKQVYje
JuYHicIlV9cWCM9z9j0jht0kZUtQLocVWAdUx2TrGD/buByGkHapTHr2k2Iq
sub1XzNtyZhP/PRmUvLFxmkJjLL6ipkduwhZVG4leGy+Y0RIENT/qJ7GAIHE
1tzSPqeinFfOyEwD3lL4EqTfQHtHK0FeC59NVwAUn0BbQKgbQXyZlmEmQNxC
JcN6slx8E60MqKBhFLWmZp8Gk+aUgtn71VVvg4H4iEr+pNmgRvwN4A9lT4i3
FAxCQM5G72XTORztzZZsrNuQza740wZ4CNraJ/je+O+W+sZl5du7lHx7R2mZ
DwMhmCcLKwQOOKl5VqxD9ssVd5jO0q1vQpMoB6rqe7jEpGaYOHMDXNNEDd75
c/2VslW942VCDjvIsVcsDa4MOY9ub3yg4IkKt0IWkdavvpzbW47aFDgg3wZy
ePMzU2jKjRwqkg31qezAsAgRL3HWXZj708YlQbeorr1/H5HhMKNIs7MYphws
9EQx57/0w2NLfxLUBFIOa/EhSiz+Ee0z5aBnV7hikaCm315mfVpRD69DGcbi
t9ntKHadhwWCTQSPs74TchBOkjceKO5iCQubpJfPT/RDMMPZcUthDo2vUJqJ
NvQcDNVOgN3sFu3q2cRzcygf9Eh9D6YQixLI3APJmvTP3Bqib7BjV7OOYa76
UB6rHyD2MWwyTLk5ReDRTDAm+pqf2t9z05mEkMt0KtgjvkB2qF1ogMal3sJQ
2iq39yymWCPqy67Yfi1zECFuYRGTu8fBkhNg8M/QBuI7LH+uwLMq/hhtIm3s
uVYVy5GpD7ZKbQIWl4k18y3lco/CryRH2Hbu+QVNJC/X63Ebv+Iuqn/S8oJn
O0FrIovgXxBUjde2ZMPx6+72QDbF6L5uXRrnyZQdOvgjiPExZHaSOLDzJUuc
6E8qUPbL/h7jy+Hj5Sryl8QIjTMFszueL0JKpNxOsK8OHcgRdV5NjPCutCfj
LEpBGgIDGE7VSsSkeEgpl+KbGyry5NmMLGfvVatBQUD4k4DshGVShVoCcU2I
oXh//KgiFizxECk4XfL73QFwOjRnNWOn6YoRZ3ctaW1EEkxtHpkKN1fhRZTE
QSm4spwbldL8PmHv4IF0zi5xgUa6AOoFzSucHWmM8fCMph52NenV5kxJVXrv
iLwlpYqKKtCvRfcDX+P5twZkuKkf7qbMhuv27SBvU8+sd74wq73dONZTXvRj
njY7OH29fFXEEiuzahGgOut8g0jySjsv0PmXpvtQmEDsuJR6ReAxkZ3Nlyb8
bbMC41yDGdwvMdYME1U+qHUi5850y6jf93lyoynX5g6njNrbVVDy3VTcqsrJ
RBYzocdmW9jD40NU0N/4ZrLYKmx3nlDpS/h0mnYQS/v2yrRz6xODK5WimaYY
hKqVg9IRmvIZ79VrShSixcclocSOjcn32/ZmIw1nCwpPH1/W4mepJysXojgW
rS6XtdzCUjf6QPFk0lhzPvKaSGDJWzsGsKMzY5rFY6qXCFovrOn9M4MtXWlt
2PLGMNZpAoiDcX2HOilc+maLVTf0cTMzQfrN6WruPj0xPAhIzpr30JFGYZ17
zwOeMkUB87qUqrMGVpozuvXNUM8eB1ojm7E+QM6ynqK+IftPKo61o+tog+NS
Kdza3UVuyVHbOwnegc2bq2PTxdTsdGa1E58796VKGKEIPqifd66SLKvdaE86
YqC3/BFJJTSCMumKCtQPhpUvVi/3npksCAO6Aa3ToDj2u5URWfmOJR2WfHHt
kpZZYIncm6y+dKQGmrSHC2wbZY81wPEK2UXzv+CfdpkdR/KAGeESIDzVXug4
jMn3rqweQtspKfnmB+8GgodSyln6EofApD/0xl4F/PmkGpNs/xQRuEXJap1K
VfHrtfPUPlEckiApIVfOU/TNaaCqO3n3N/IKDsp4zke9g1umpmnZb5IQ4sAK
Yt4k8Z++qFo5NoAzyUVXEHXLk8ZQffgGQIahaalr722+Y20uKKYYgmG13QKG
UPsqMSRzbA2uSpZI7Qz973MSq1thDn0qx9WMzjqET5PynRw5/nlbUqOUMwq+
nw3+dkXJKvOqwjzBqZBgAmmfZQEOg+Z8z5Lju62yNlsrTMSzhmfUvry6KQiL
U/FueIfDfzSjTRey0KVG6s2ojGHiq0WSATUMOuWPt5e2hiKqevKFvKX9qoOq
QMzbET0UvV2C5iToRGVu1eHU310Jy1QxstJr3m79zDKzrwVySqeQi8WhjojP
dCxpIGESJlUaoAxazldFnWRRHYaNXFUI4DXs0XewyRwC8rWZsCdV5x57sWT6
zYftUshzrGAv/BoVUWGTphvOpeccf7NDPa161A69yV6rljFq12FBZJvcer2M
W967CK3ZdT/6kr3zQofCIYUp/ugjpmKveS3zLJvEvg+LlT+gnn/e7eDHQkAQ
gVC8eX8ZYnJw7Uh0y1yL6oS7kI9notb2OdQ0m9+umYA081Up8vBhPgnA/Khg
RQXJPCEt/OREBuNqB5Wp1PnKWoKZcvOBYSUjxdfVfzrtV4/yy4VwgN115ZLZ
G1zd/KI+qHrHmdu/AROajhEokAnX1ziTzo/aeiqRHa5Uy89LbdyTT0HBRcY8
t5uLM8LmG3FOMiMRW3Znhw6ZnVCaYjVvkK0EdlkMfSTzKYvaZRBmmn0q72Rd
XuawLZgU5+WEy5HJ+5fQ3CZakHvAv6AKjQ3z2prY9q6Q10PUzOBzM3dYWMMR
o6vN8gCbLxqFSvocmiUIfqXzsE//nAgaLzJ4c4G5G4aBTX1hjiuAI+hDHA0M
X9+4/IfuFLi86VZ09H233v8lSaHi8jfjIfZ0+FnIWQOlvAfZT4U4iAJWXC7d
yCGB5lcmXGZ7+AjmBRHSpW8A9Qqvg8WiaOLqkdQi+G6vuXYQggHdTiZfl3WQ
lChMGiv1Nnd4bdAXKOjYQghukpo9+C/3uDMqpnvdPsR++3e/ifqi+YkEfK1y
8NndSvnXCw7vJgFHREdoXdrDQ3oslZ/tbMejVf4LbXlwAehvjbIAWheuUu6v
ZeEaqvw6gAtqd6UMVV2EHKFCN5JkH+5GpH8KgjMJjPIR9EtsnPJ/Wgeg/b0o
ic3xMkCDbwzM0k/x/KEfAsfUARNRyOBUZGWffucWB3lRB1dnd4UKe6y5qYEs
c5q00MSQ/a3izIGcfTRx8fLulz6jzAKVOiYGbkrThl/BpBX7gms+FS5EjbLy
9QS+uFxpYzfOVXxi8HrHTMEgU4jSaZGkvMYnz62Buujq3iYqRsNSEL33BJDl
Rxmipuybo/yDEleN0nfv3zekEKYLX2p1GRegEAHRxzEqEifQgfjjWV8bPoQT
nyyBrKEvDNvwh0afxSLSaDllSDo4Pu/NCnCQu2MqxhsHgipgdscDNYTYBbWD
kQA7ylVRXiUETWcvoVk0L5yFFNKpsqTCVpSZj7mJUj7+jneuCRCx6UhNyrU7
rPuy2BIf3v5MX2wB/IV76LpsbWvBkZEEx2b5OUyIb1jIuAGkennyg4Nktu6V
k+NyvF/Bk98zXJ9m2I+asxUiAdsl0SYLcTrmedmYNmgVbL0kJvSWZNQyqFQv
IDRfVC+7qLXCARXqflRuH47efoupw2Fahf5uPNVkzpDPSYBik6jqHav0DxLj
qGCiTA7b06uRfqgeEcVNy8qgbvRtjOT2378DdrioDBqT5kCBSKkRg9dmq/XB
ef833qOWnUVB8I0E/453z5/JXuBccNqkpoESJQFhqZ2poJgz8YxZqfLh1XKs
CaZo+2+iEPQ48aDd6SIxL0ISQKagi03RAlk/gM3WSx2N4k/X3cid1Q4WRhrw
dvIa9CCKEWJTzOETXYwDfo7ICAy9OII3lgjMYVzJw8B+Bq9elEqhulKncby7
ZXtdrBpgHPVOtT6yUroB7H8zeKI6+h18aq5lOOX0mHVFBGmrxBR5IFNUWY6O
eM0VR7dmNxsQWkuyPrXuDcEwQRA/xLlOUZ2Y34kGVR4rakqUzOd9ZpmkRrue
gQhbicDeCcYa0YZahcTGOuuxnB/uD6Sbb/xrOzA03MlDc7R/ZVRFmninrQ7c
G+t9wmnXKl0nl5ghkb7wjYqyR8e1qCJtlmCN/tzXgm2buUvHxnkvsGoJ82en
Uqb7metgHGe4pfeLko12qWFdAM9xMZmptEBSq8gDhWhQ0jQyphrP8T6D2Y90
E5Ezg6cv6kmDqCto7+j5zenOReSKRVvroknqMUqXN3p/T+uyd+wiatJVglQ4
7hpDnHbTd9Qxesbjh4tXt9N2S/WXBv5zlrn/32k1/LMToDoeM3N7mbw5jP7f
QQ61Wm3Wn2G2HQkBX6OqI2HVuFrMvJDt5dpP4SM5yH9W2pPzDydRfIBWdrdL
V9rGm8N1KWDIX/YpF9TVPWTTL7XAINW6+ZevDRwE54lHyWEeS7lwozopCdWN
2MgRaZGcJ3/szS7JVLICgs4SyCVZVRcsnwZu54DugNKnG7UZJLouq3Sii/MD
z+7xRa14bdZ82mDo/jrKUJvXzQk0o+6F9cvzLGV8pQsxX7tfNrCMjiYKzeE8
YQjnXbfTbpIIVlshy25c3KEZ30AXR+uzagFm5PmIUOsOMTyb2+0wN+7uTBPl
pCeJ6sF5QR+kJWijhT1CkXEUxwzhoPgGM4vwiRMTyZGWvqfeBGiTQjJThWrf
9e/D+JUBQ7n12BZej+L4J2Ew1VfW/1qqmzffwPJdi9A+3qmu3r9YSJ3axhL7
hFjqLq0RCOQfOAl/3F0MZ7Z34ZFEyr+NWagtNrjpg248i+gp6uZ2ZWRl4D2a
y0YWpuIzeULrQ9WrMMSJ5cu9iD+Q9d6skosCUOPvhR23HgaWFvYVqfHbEvuW
pwxmpY660i7k0RXAPnqnN3IefWFW0Zd7Kg+H1xB+xzJvaxxw/q1GfDbsZ9Kd
jnYQiiiJJmGQqrRACK6wTE9WspXnXmrwLkyUQZOIKwodVQr7v320jvAQ5KgB
SlUPcWdEeSxsScQNJFeBpXbH6ck7kn4z5afLx91LLwbsXo11RVlg/vz7ML1x
yL9LBj4QEdsbNof6vNlJDpWA6233NVbF1reF/yLl65upKJIwsY+1ELXZY3qt
QYVjeUtgx2mgJbo1Ag/8pe2c+8ZcmZHMGS44Y8vgjjE3rb8ZtXeI0RxoFhMl
4eQid8TNOselxXt/JvaWs71W9PXnV5b4Hy1sjcLv1H77VC5WzKJavnWCXtwh
FfcQRljoE6y0QfY9rjSxcZpTKL0825nk9M3v7LLoFXcBxWa82vY6oJhWh8qq
XVMuKfmoy4xIw+TJGjPHR0ZdqxE8s0DDC3PCmoZrgnShIGe+KdpaQ4GxfnLs
mxrs+OOBe0SylhtGVVHydt6BSJvz3lz6uPlS8UKsy4c7Ns1zlG7w/2wHiXU6
LDWhMXjccOEQRpbZ3Ytk2s8wbxV9uwz/2OqPBdKDa5gbcNnZdqpBLTch13bi
UYkYy5B9D1vwG3M3gZbKVEI+FCbEKaUiDNDL8nWIIf5FMLO6D7heFIJTu+4k
AIIoAKedDE03djGlCHWdlwLgGFSayhvV8Ap8w7wGkPwdOVOCafDUotNxrsqM
dxd9Fs/ifyQ8gKGIjB9PxGB6QREWFtK4AOj0PhmBr4mpcdLz7/By+71OqVQi
DhSigPc6Vgp+7jmo1swrN9wfATG5my2B/6qA2c4jmEyUzqh1z7XJbcCMgp2j
wdJezBenB3xyYaRJreimAG4hI9KfhiV/zgdu703BRsyeJK2ILuM8he8boD29
zDtAQ+NNgDIjmJGzYtWG93abcEjdQRg8sSKZq7k1SOXwdiV+P3kW5Vs2cp+h
u+X3OiNMJmd9Rrc5tbKczGyZd9vOmouC6b1pDBmRK6bwzOdaxNcNA3aw3XTJ
9Sr9jmshN14YFsl24etsaX6sGmUxKQrn8Z1iWNz5w5l16zGsMGiwxtfUbUwz
7SiuSJYfHKZzA1pcdFXZ+0Dwx9eikRgkJPzVVqtul1qOAQpr8ttvB7l3Gy8t
9YdKSzEyH+nQOGkTiXjMfmmmSqwd5ZL6iNbi1ieikca8oct0HgUsKk6lMkJy
qwanyHrhgaHzOLXY5MvR4ICdgYxKcuNnv/0tWhoqs4pMSAeu1wXXat4veCoj
fb1sPX+jiA3PTPeeqC2XZ14+CId0WAcGK0tuRd7eFZpyjGP9BH6F2+d3Bxqn
nXgqIbv+mZu1BU7cAbPeXtzlgP/d6oByUh0DrioTdusQAyu7ca8y4GmAPLZa
6Nj7MQsflb8aCxj8wzXFjN0sZLRDEMFIGf1hqE56H9NGhcc4Y0JE2L/pmwrv
oLul7NWHAEaFDKrNcofywP+rd3yut0xxU/GWxJVRkWb2svU2hIYPikuqtJUX
R2IdsAt5OO8cwrTYqiwnq1xrf/qIEPS6RM2oj1yp3j/a0oSOMu83GNpEg0QK
yAEBnP89N7GDQf7KGo7bvh0abOJuge9l7rVB2OUaOYvVexmuV51Cc1x4qpNh
CDIJKGeeG6BA0miKTEadkGqfThTUbmSGUA19DiLXzOHMDjFbfHjAHsIdf+Ze
K4hRsDxs9uK7//tA/jrQWh2ilKqfnqVs3G/JyOOoOk2GSSoEn3htSHlmFm0U
fhGhLPwoeucVlCY4LtHMTtdVpKIAmWST9ehNQJbLhSytM5PLJHcexbaU8D+H
JpcefCmgNtT9x1O3BN+K5N9uPQG11Jm9EWLCCZTc+YLNssgBar5/ubg6+WE7
gWT3jqz3CPOPJilH0WiOPF85SVwDrzDasliLEn6tYhMFilUftMC02/iFumNH
7a1VTt56MI2aeQdEehSLDjDm70yYtcrWFmahidlNzIvLCFTgaBPydil1hpKX
qqMl2O+jJ6KTJpgDed1OKq7T8nmADldFu9uZwBAXRQrqnNMJCw+fE25P27qZ
/H6ABdZRZm4YIzN3ZWrS6nITUa7UhAQSTta7BwSnRw8z0XSAF6tKNUSQuKPs
2ozsVjejnRJ9/Tv2hkTbVLiFDID8iu10LlwCLyTW0ZYPNG/lusIO7WAUfbzy
KfXzgi27npSoaV61mLYL9StuyjLVh8VErs6ssDP4eDhRJUWZUJ1VjruIXYQX
4VD1/Tc28sHyOO6xCdc1B68e4sOsYnega84u7VyY4bBRoaz448YtYQCRGk/f
U1HnZkORrLlXLs3zQtlGUl4PezjMkeU61FhYG/BDT8wflWsIZkLPy61cRGXM
uDb5Ue/vlOYCy2Q4Wum6Z7tEJuIVvoVIScbe7EWkBXJuIrBE0WJ+b+8vBvMV
tMPqSXFnkFEkX4cqPfJf5PFsCQftkwfwNL6mIbAFQytM3dnPJnPUcNc4EtHZ
8/+Z8NE2W1rCUjvEitobeyDEg7x7/D2HOM9jBUJSM5sPCS25vc5hfmTmCyLp
pWF51ZZNu956JOAKvc/h1xkRNNTxeRT2fFWc/0tY9TI1tSTDrqRbGr2xQuDc
AwXrUmPlKkVH2dLpannDxdcLG575GEt0Ls/wKq6x37ING0AQCMprVurnHnRg
YTK5qSgFcZaweZ1HMp2OH5cYX+wVm4Faz5pjPp8TPo4KCf9xW/Lr6AqYG0yt
7sdp88IZaWB+ZaQ3YpDpWuWY8unRbi/yGgk/dOWww1MCU2OMBIVP9HRDzssD
6wzm9p737yppHOCSrHvv/uUQTIzU1f3ltseb0pqTiSYLK559u0jKaB72+qka
GEd5uFsKewVrBR79/kUI/S4g5eb0Qig13qO5epyyUwDB1LNiceOzGrwo5HgC
Onmq37WD745XE7nRA9MOFAgduKee8LJUqEJPs6FrhN+l2mb6WSnQcSZb00zQ
3CHpyBWNM97rRUq2snZ3VZyVuaTB7zqy6yuzMdb68cTIaF3/uECl/Ed9EB6a
UeFXRTq/2eAmT0RUIUhTxpQOW51KxCOA+5J4/ADon+n10ivqXLBvTT1hPDqo
iyCQIvPdimY93461kpUCO9WWqffpD93fKf3s2cpVW6VUvt+f8vi0qMVTxaH5
lKGfrbjaOwvpQmMtfKOTPaZzWw8uQXVLxiRy8NBW7Iih2i2lqddaG8Ni/NGq
P6B+WoBKban7JqzsAsOSSbv2+mDdOftRjH7sRvs2uD43DiokZCakWM4z49bH
inSMRfBWLEdev7ws6osV+NqlJzKvsQopgl2eRgFElake/e/YFx6FAzTORVc5
tBlbHaQggUMt/ZYBapd3ACTCvLJElWXWBdxMjOOdxrGkwVB4Fa+rhRg3e/cK
GtfMo2/pUiqWnR9kGh5ukmxjyHu5VJJRCl3vrwBJl5XE1j6A7xpy4xSbXb6f
pxPGPsOUJm/WhYpHvH0+owaY4+Yn6CaTxEb62FjA1lhojjkyudWgY/dggwS0
LJctF72MrBDmSeJagGn4W3vogz7ZQ9wD/WBvKaBzBwDkSI5XD80OA9boTvQl
Aq0JgoOixdDHmDrYy9KePvXpkLV17DjI9BuL1Hm4QtSFytCfCbkfdyrVPqO4
wjKb4kt7eeXKzceaPNEOyerBZQQEJJj4HV6NkTsgEcMJ6LCYOAhGasGAopnI
hb8145gEcUbTPW25peZtmpWoPoIkcpLLKYNxKXjdXWGd9Kphwhu+zaVBgO49
yVgUVGxq9j6/m6eJfVJOp7XnRDp4LH5WHyKJGp1y1FJPampgM6AORbHJxBjm
KSqhbfp2wpcZi2y3QJ2Ht2jUdAWvvqlsNdz7fcYegjTL07kEUVpg4dMXSgU5
7XUvlHQiHd4o701TsgVOWx0UoxttX4vJIzcjxDrc0Q9qQTYouPKj59DoMEZE
FaV65GttZKol9+uAPJRAoSXC3SuIPAzl/JkVll3Nw4qLYB6tGW54uXOIm3l1
gwTqXi0GhtRd7IAF7B2K+p9hmZnF1tMt+VxsPsEQlvuc2ZlDktILpmYo0LX9
0+n0Z/lxJrr6amfSng6xQVeOUJjAM7VXt32vIXopyfmEShaUJIhmLblc17qS
gTbRrG4u+Kha8DrSFVY4FSxQZN2OGSGUClPsKJGZlW1CXbOsld1fmfDqvCoK
pgPZdKvQmBwtXFjMGqjckfJgTpgbkSE6zjbr6vVZ7ZHBhpFs7YydhX4YcM84
cPnhNB4LzxTm31UQPQG/ZxHMTlktyUv2jUBDYi2SGvmCsM47lG144B7oraFf
fCSqh25z2uzgKQUi9fgyDYWhXDuO59iI5bLyO8PIqRm6yyTlCwvwcbhridGE
Ks5CmHugTfK/UyQxhn/H0F9MfQOLi/FXhWwzx2YtJZ1eYrlvCtP+yq3ayI/X
/G58byxACGg9esXZc0/lbhlF4p7imyHNGYawsEXeG9O8dW8S78IwRKnYcC5n
tZG3lOj8I2M4K9oe0Z9B/u5zsulaBAcsSOAWSHnD+RkGy6Ic3Y6nX8Fghizn
ud1qpVcNn9V2sLKvhd7l3jBtPy832tP88TjUSbfWWyvred8KV5s5Q8FWkJtb
yQID6eFhjbmCEWVo6aKdlywDxmlJOgO0CX3NvCPEiMGZvlg87XuFZxPH8OKh
2faqvgIxGBWX7HLUmKUgs30vBBPpoABV2ujm3aotHO+WU5vQHN1x9brLwnE+
wN5G3/gxPHqLriG59pdt/cmk3V8khxKA/3Aq2N5Z5lWGbMHFcbAcfrzPh+Wg
eeWGnNdhy50JX4hSXBYdBQJvFt4JiWeSO9Gj5RQQDFlFD7VJvKcdUxbwHw4u
7qIqPEpVjjxmQ9iJGx/vodo8Ay9IlNBAOu+DUDpvYwvq1JYPEU/b09mLF6iV
iSShl9nq+j6ahvRvB7/Oqhz2apUaiHTaPqhe229/FqDzGHoII7xzA6vKcWIi
ILkGlQxXHXLmJcmkL4UGbGYOGjqmV4mf7JZsVX0zRZa0mF8/oG3zErMtipBV
KuxVCvfxFrgpux+9IrBHMt9oOypADfBczxDCawB2l3egxE9x2W8q9JFKUALy
eHCBIW3ZdUB4WdbEilU8vrLp+NKopphBn9lo7EkeCD5q2zHlwVppuCTniIoD
8SlPlwiBumz2LPExMHm580SjJstye5GCzRLQEjSSVNwIDd/sUVKEUKa/I6gb
JrFs6e3WTp9A7jphbbp7fk3cWr9Jk1bk8AfISSyjEvCdl4CvoJeYWNFcPcjT
aXTusgDaKCoUeRlSnMAqSEPaxw3bLlyunBCFn3Tp+FwForypNutB+ZfxxtJm
fXIrLLeB5htrVuxMDEhRMO0FBYt7Krb8g5v/6NA8n43mAXHnGeddxa5UKvPQ
H6H/rUSSsdOym6M/oVy5EKBmydw+Zq1B1q0VkWOR+k8zxYVBHYpjygCgddwD
z2n8OZVxGl6cnw+ziiplFT/8FqBVTPJh3qeqmAaKlYR0S3MSzDE/Onajiwbm
yUAOqCTrzJlFGzmSnYlrETyrs8JLk1VXJH7YTaiaRf3Wb0sE0lpOFcnbcF7l
Y5rN9WJH10MI3mlwJH5uIH+5ONAIFelQBOoOzBYtB1XZBPZ8qnnowAeKiinB
XhRpk45Wni7dXTc27kI7M6EOoi2w0g3VeTHC/XI3hl4JmWX+fWiZBdhutdGG
V42/emSRPzGf70MPAI5NEHdIuMwhTQs+r0BqhFCUledSyHdHZEzMMX7dP09W
tvUDYOyNDckm1I86Q/uwYgXb2BMcYvffk6Bt82g+FnqbtVTZpWmWKK5e9VY+
4Qd70TKxPHSIywgsimCcluIbG6j/ztxLyxIJKBb/6nvV1QApe+hQ5OLFKqwN
cl5zkJ0jcO0UskocpuGpCDqEKxDSWTfjmyUdGuB35brc1/gzOTP1GvteIfZ4
yqlb21T2VTrGxUcQcdMeWTLkyw1B57UY5OXKfoMXDDIWJpj2ooNP5kcbvLRA
N+XgPKUssRy5fGOGGuCAuLgcf5CsMiStx07+p39c3O837YfBBv1yVCsnKwYv
avMJGKzcn/lv3MUM1kIKUCw+W9Y07EiGSje5vmC/BewIehnka4l8WtB7uBH1
bOGflmTdexV69+hqiN2VKTMpt9d729B1np2hSw3hbMf36mpwdnLbiyEw2CFP
TxsPvaksgepjBMZegwfsD1FTMWeMcyL+w9VMDa2sIznHl14Lm/+chk+vG8Na
dMlO6rxXk0BDgDlgR4ARHeXuaZqR+oGbGOOGv6q1EO2CWoRysV7bySkRXoyf
LOmmg24OaaB3c8xiBsx4bSR1pXrt1xqDNn4+wUGNIy/CEhwWvE6g76995t2H
bf4fuQ8ifIN61zh+r/kt/kDv+zAcahA04/OohZefR6YpKHF7NVDdjCnf2w2m
R3ZMel03ES/7R5fIPJDZzGKRA8+C5aOGTdh/89F8ANflJcDVW6VHWk9nca3x
GA2xLNJaHcaRyJlCwGIIhv0Y97xReXRyPDpobAAV97nIn1OqE95hXlrroA5S
r+JD3+fDMTnpLpN1DAS1kOwPrHp/ry/n2kIcJmGfu/0cZ9z/GkVYnnXHcXjM
wbrt/5lDty7XvrEspusSjfz3Y7ban72FJFBcukwYw9VhKV4Prx5z2imdBR+N
lJplVWXw0m8WvgxTxDyifh5CBNWhgQdID0Ny7KYMTufYWCLAxvLxTuYisYlV
oAyBOICa2Kz1LbitOGyUyClftM/ap7hcdK27f6o1THeKIYr/XaVptW32btbP
YuxJGMBdVDyLGasa1BVBG6pIX/v+vFXLW/hV4kc5idGG192tDbSTBvfFMr+y
n4hu24BpQ3CIF1b8BTdWPm4bEkLp3ZEWvUcgOZvHju2gP8T2tYfaLS10wI4Q
EwveJDcCoFknfR/1u24Oxv44LqtK/GRravz2kYImj1qWNFSR03UQbwoSPsSO
8aiAfJGv6cuNnpe6mUkPySs4yLXwBXr9bYi/EyqlHltCRRjbX7Ci3M10iORq
2YgJXnWmqWlVaeRN3EtSiKj6TiqlSWvktn/iqy/wlzYx8jDtztMlySh7uAIr
wnlNigiM0WH9y+hQ6SDPutaLH78HV/v7c4Rs+gBGjdHdPW0iyzs8abz6eB3n
DphHQ1S9rBbdP9AU8DQO7viRPtVGMHHQx+D2XSl4sLFeNIKKIJXYYZTNoBUY
daRmITx08q38PwVjeeUjpfoUHRX7dAwpC0IV/oekgiDaIH+Igvy05QqjB6kE
J50ER33LJuBxPJXsacGTmZbAc4ZkAJ5x8EMMutM7yjICw+smMCqaSiulxIpj
pH6ftuGHEBedYzq5++TJuuNyhCAGhvcegausH/12C+ZvoudgrPl2B7vkvKex
j9CGTg6URD0IoQMjqg1gk7Y9v1PDIxTWm3+oBkc1RsJ7r3FnRXSzwpBNk1jz
3s2qXnEZWmhc7UrDAAYsbJYEwdABwW49MGpVbU/9UQnJcfvngB7WbxliG/Nb
UzpWOfprf2m7+ENrkBjmijKf5A6yeMvaLwfk3QjwZXJso5AYPyNjKSegjro2
1rE/EcvEZ3TrZsuky8xtGzx/t89Iwg0JSK2aE4Nyi1Wwhd4qxww0Z0IdJGp4
fm3EZM2Tk7Lf0GWIQv0Hf/iIuwQfYhHpR9SvgZi4zmrKdAGoGJR69Ngi+yI8
qbemQ6t6wJDiyvL5KD58GVjyJ+JJO+9oJw+0L+cG3TTmVivajlJeI3BD8SzO
UB6VSXAwLXVf2wi5kXa52iqhhNh5kZWGQ7loJgxG7lZaP5QtmOp8Rd0V4IWL
9wwcYBN3pKgvS/oP9vwI7MSjtidHE2ZT+ciI/s9QLkdtAHYkBu6Jukk2JJ2V
oKi7yCMuqAshtrxbIpq3mtc9IcB99nsfVN4IePde7glWgOSzT8WhhNwF++4R
/QXKU9RaX9ExOZACx0YJKcsfshS1uEGyAwQFJs7kd00VDiILRiSPE7D0gg1Q
1eRXmKyvUen/NJcncsOcLGBx3mZO0udSN67eyOKVBK0ixwt7Y3URmuKwtlqT
nbmuw7e4m6AaJp+099arT6eIwU/gpA5Qw+cULvJ0kWbpHDSF+XBt0XYuuNic
pG0gFs1yY3ejBc48Ju+GBrFBQQYT0GHPwghrXPqs5jgBwlgwNKIfeeoTxhOF
OsELdvoYZ9otJKHHSsIqpssvxwSm52j6VwkPTesrQT+NgYBdZHrHPtm1vjK6
Cz+mqmkMTZO2WL9ijGAg7L9iJkidX6soy7yVTSvm7InuHEmF5za3Ayh+F6pi
Q9lnKxqijWpPS+DCPwK6ssmV/iBtYvn0AwlEvyyvMvO1FdxMTjTs1s6zljh+
vmpXrL78MFLzZJ9X/YGppEFfLbC41Rsh+kM+0ReMqq282anvsa/JlyvUkZvW
MwJvErBxH15fxClDBLaG3oO/caWY+Euq0TqkiTYrZcwOBX4oD6mVDVMzMdu+
qKKyBIWjb5Y5z9TwMRJG2jwiluNLdcxTnnhN4I0zwBnNfAWWL8WgUm1KhZQm
XjdlI+6o+eTlt4X5nk9/+CAP1vL20VTRP7hDhTHu8f9iAmODlQzAEs9yXpph
lSd8yollJVyD7rDYj+wyUm6pYyr7wPFaRBV6WOurBSuFqKOToeC234xmI6JK
LTaH36s+VdbFDFxn99syZuTpCi1TAeRRX5nIEEZ4GTHKRKce/cok4q9/82kk
yB+VssbkXncICXOSINLUPgJ9RPe/vVxAdNpi5nGXem2LFtaOprPAE+c00FwL
iZpzgMMY06pk3ZrK7UwI2YdNQmAYeHeEbjNd2vj6jT/8fVeEhqd+ZaduFa3F
+Jzz24an0hQ99junkFg1BB1drzZf3BN1AXd3h+kbj5FxIV6nMfVkWeDiq9qw
zO3ADJ05ar3un/lF3MwxTqWA998im010NSQpM9AohOXmTejrotWpuudKu6nn
2bRqjPCM6FydXVEhjGpLbApty9Ttwqe73akrGTwnXVLdswEDfH9HJxbb0tIz
cBQh5aT8QwiMRq+3p2JnKONKaw1UutBybqvn5FoD3ob1DP8aOYTzqI6ZAG61
Hs+fkc3ylrvM29cej4ceyRWu9UQG+YqxTB8PrMJzIuKidy2NaW/f8/Kwaqj8
fL4RrBeyWEYvpCfDZLI19MLl4k56lr99JSntBJJGIrAbMpposatExvZYoOM4
N0bdqxrVsv1gD99yc7VzczWJamrToywP2NhRc32aBMTbQfuQpGCwuUF1CEb1
6dXAnFphB0i1NfvFJvlo2W3BxSW40gE2VkkGOg7G6+6A5ks44HJPGQLPDGf3
x/MhQGRm7pxaWbSAIXO+zVAqtlGhndxzr64M3yAFmmdJwwq/d1YiaaMRP7cW
+UvslrPjFNc+4EqNFWVZUG2oaNYzGzqnlOc3RrVBZPitETw93HwxSDFedxkM
XimbWgT53BB1F1Ec9q51Ps8HpIIg9naZYstz205lfl0WLFnNI6Had/e4XZsP
MMndbDyNDiP80ryuEEgmvXlh2zgt3ttlROJDY+4rjNS0iJKk3wizou9fbU53
EyyjZQ8lwEBQjxYWsWIHNn6tdrFflqG4sPky9nV93XxsxgMkKAqQXjSW9IID
SP5PAzFDPlQC8e7PcESvEw3MbyXh3xDcOi0luGHkj2mu7iYP33nBI36A7LkK
W2aT2OaFnSnhoQeFp3hWQ8ReYtps7aHUyJYMHiJtJHhDkwAWhaPjdPA90E44
JL5Bto+6vqDFeYVUBZa4gi2lq1iZ6bh8AA39ODSEiH0/gV4CGcP4PjXgFCBg
zyg5B9Fkf9IfOIbxR9HSufWgz5i/RAvsFTuAGK6Pl1G/zySAnx3aVxcgNlFy
998LBYn94mGisgjkjLLyoEPFyWIeIldTo7LjSvq5WklL1uSKEhCnD4j3Rch4
7JdxCK7WShsRjcpKOkPyYRU33wTAFDJQEtXWzexIkdpydKOiuh5irQ9PhoAo
z3qqvwN/mgLOvK8fiA1G0TlOtRn2cN7MkWqOMwqcWFhvdkjEWzj5DEul34PE
FDKqk1ApsONGcURN28YOXHT8qZKILuxnZ+p/P1YhoiL/yNmuGnvYvAIkKV1M
7Agwhg71N/S8LQRg0XOG6eUSXKUKtMQtpY862XCnLWkcl+W9hVwLan7/GdYC
mzEqTfs/rPh+bzYbxe0SPPdTnCxkg+legkeXlo56xfJCs8BO/JBYhHu/xfoL
t5kayi9QwBKTWVa+E4KIFUk5Jrixl5i4alpipaprP3esIhhhA3RE/SubktCF
pkjvfn0T/fQPkcfvEKJuz2icBsfYF23wnt2/7tr98fBwF9h598SiXTgUvVnu
7lsEssZhkTwD1wP8mFpO02HKuRRYk8dJy97lwvnrxM2+2csWosI5BJFYQlvm
+pLoAI8LPxPergsCRXW7dg7RfhwYF4wdD9iaJdcasyXWJn0mXudsafNUBd8O
seFwMIP8ysYb1iXUUsbYmjEUB/4ZubNsw4GlKc0TogCUZXIkSBz47fR5r4Bm
tx6v0McRIv6QYVo7Q1u7e7HCCU+q+4fJyHsQgxXYWAJQpkQDFKhTgVnQQmzv
AmDyRkoayUyorV/uYYz+dRDZ+wodsX8dWbeSmoj0rhwC/W4AlBd7BppKrgrk
Yln5Xs5TqAJkgQ3x7M1qP3xOZmusUuZin34QKDRMKTAZAzl5SdZ4K2N9WRXD
hHCc/tW8L+3Su8WEQt9rLg5giluSLxM7VcXBd1Q+/hUf7R0DOtt0yn7PVOCt
37BwXXpXhysz7CtR6N5EZjoUIqhHYVbOkFYMBIbP8aV+WFOI9SfgoEa+VCyU
OwiwxgyT7r3DU7u0Oua9nAjokLOEampX5iWsaFeoXHLV7YmwfuJZ4u04ckAa
VmwTrhzX6TpUoXTd6sM2xmz125DzpRBXtpYFMemxMX+X7QBAvtMqtJDwSR6b
FnNYjEMzfnKH8wS+AkCcMbGjv3TMMlXdwI0uevU5IUL9x0KiXvga07iF69fH
FqldTaRG++6IeG1/p+FOgKpl2sDIXk0Vm+pTCJH+g9lcD7Dz/hKmh5qFWXmG
xfp/k1zLuIb0lpeSZejrL8TarFQYJA/hfMFEjbK361woza6ILYc69rMzKiUo
QxvBu0e0d2tJJy39Do+iJ/yV3Bk6+rAJ5NTPCFhs3u1w6RStjZU4skfDVF8r
JWWHUckR/GYfT8P2H7iFv+EpcJtCUF1Z4irKT6Zq+QmK5LMJjtcxQOXk0NjW
yr3+s7NOFDGD3IJTKhDXtHJb8Jall7XLwLYATpHaLHYs4ViztDiLiTTwa3hM
xic6KfS4PB0QQMsHoL2p1BWX2HYJaB430BastfEtj6feCq587YTjuWFLAUau
LptbLgzQP6BnCcSrp55uAIrcuJTK5vhsdkUtb3UGoaQQ3FduChYsnFCOWXeL
pRDa+zFf8C89/qCDvNiAC426AzdkyTJg2nS3WTXoafLbsPyVdixUeHrSra86
+lXvmSthVLPwvgx2QG5+6Wo+Wfen7WsPB3u8BMGTWObxB/Edbp2EU8OVtD2i
3swJsh36CAdafUbuyw6tyVCExX7mG5Z0D1W4V6x7/LHWznP1kCqKAnMiRpfy
2Ng16SZdM9HYu2nCYuXrj+f0JqOdnhvv8c1GAF4itwG5vW6W859nql0Niocj
+nu5GDCmJTF/FymwNEby9swNPyIv+ktZGzflMJkavR68VAWzyaEgVbp1dGHS
S9AxD7cCzFWiZzxcuPY7l5U0vKgq70gA1wicv6RCichs4vBna4fdW2jaL2Vy
lR54l/vDWp18ftfUrw7Zhuyy9ZExcUOE6UNMzLxOH6Vhmf2NXzEjczEEGnBB
d8ArffxxSXePbhgkHqxgOk7oB7d6mot6hDbkuTDUrVcSa/CRt2P9wJXwZd3l
yolBlPfFma0aZSo05ijz0eFBvW4Zr5r8RXPI1GYpxj6CGp3CUTeN288YaBPs
dIVGYbZ0fZAUeAvLJS2U7RSkOvcJymA71HnOb+oWrh5Leib/YzPJ1htUF0n4
9BmXbKKMtfYwO7zkxLN3piJBRPAcH+t06BZJ4D6VuHtwHps0eAdV67aFFJnt
mEVq8PUw3UenZ608aa4xTj1KHbKY3pb7kBvq3nBHveCXx2KEMVgDyK1FHiWq
zZQNDAaSdic4a8NZgZz/Qlco+llxoULn1RhgwceeL6dpU3m+YLIw+7HeuO/V
JYY2OlQEiBFbA3Hh7ZLWUGDX653Or61oo0ZEneIYYOAzHdr+Juo6m9G97JEt
ILJy0VqInppX+LO/mOeOPBG7nII+5vyrCuNJm+U/GErv0FEIb+GuLlNKh+X+
Phk7pVBl33urudobgpdwbqsrHWIrK56Hw2ksVf/nsfCYjSKnIEC/+9MEBUOm
+eFiFspxvf69veg5OPVgn+8a8njU9RnedQQqT2rJO6eBaA/1Yrp19NCyN5vf
WvDmJARiMLI5ekgyoM+OevXzTid0O9fSScPXFWFLjm2Q9iEH+86d4qd+Hzbm
FrTxafLhuuohHCLJFjk5W7iJf50xBC0b1oiVxCtuRkYZ/kY6xnYWy8CwdpZ1
6BzqCnWblGG5ZVbpQ4dufdRyiBPGTDxpgc6f/sirg51Nd/RkfmaYP9zjWiiE
i5pHGMl1b+afcSkmDYSNXoBfgW0lNkKurrqeuL4NyjVpSyYkbhWX/pIEM2z9
R57WnkU/QwhHb1zCfgvBTW2ekZ0htSZFPP2CPw9Wo4hl5NXhv04NipHNRaqF
RzXqfU0LT96WGmgNsk+n1D7CdM2UaXJ7SSgnLNrA1idMceyXqSJzGMA1TEJX
FpEPoSEkOiehpuY4SU9/kIxrD0yWboo7l+dZDmyEErzGTUnV8Vq6aVsD8dnW
HzEXcVFPx7FKrhb2ATVp+PeHfR5asbuQulBHkbd8SM4fC4gBnTov74zTlFoq
/jhRY3TKiZ+z0+uKT1z/5YmLfPcAI6mEWjrBLdghbJf0LXXMYa2YfRgrRp7v
HXCOdxGamNC6e6oKyhllAzR5hzpF1pWljt9dwRA4d1K0OSbCUNvEyNbdZLMI
NnGbao9VzXiGNeOcqUOh8aRe1xOw8NaLvFqAe59wNUDRvRTl5Pk1dbawdXF0
tESGHT4PZjKi/KH3qAgcmhTcEbMjoN8iQyPEBC70yqcRJCu5O0XPXmsWVZHd
FdCzENzfiA06CGkmsHXmHa4Hk9SNtdejgnNXCN2PyGQmG7RsItGaBN5brLW0
VKwycTG4tbDAA6i3yRDfZ5k2JcOQ70CN0WvStgaDShxYRNGQ//cZD6Cbx9oV
UePlQZVxrr6NPkj5QmRrde3f4xg0viCotZwcZUHiRm8+oiqAY6utfcP6wFxJ
i8/zXdW3RXGQp1FQod3gFn6OCG67Obv1clgA/Jf9n6pN2OrkhL7Ear8bHuUo
P6lYgWauj3nVuWy3OCtP7lIVhLk2YXxQuTHWichG77SuhK2S8NVxoYS1PaD4
+NNvsk+wdeHW/aK/qfAy0kqZ1MVA66ZtWcxXxfw969+sLqQ86BkpkixT3oTz
LRiRemEBZu0qQl5SaX1jHv6rVV/zERzuYmjuOAPnC4vLB0u+XcOI6VWxi0O1
TvyRxRndIV9spqT1YcNlaWKxdRZGQPDV/pSXgmSOhLNo8yfTuW4UvhrCxL7B
31v/EFe5JTnrkfRlnvflqGXEGr/MTgZr6kiMv7XNcBHEL2ty7C1WK92RVtAq
EkwKyc0OTK5holrllb+lOaDVRNIu4dSOmd84hfRGIBT3SYZxaZS3WfAja8A3
ojrAPrTRF+oXTNgugSuef7a8cGvZ6zQSF8b2PFqtrbiFoQJ84/D5ddGo1Z+N
srUZZ3nxqJggYzPV30lXLDH27wMRTV1JZZZJMaahRrczATrYSw30QafRyXiV
CNoRkgn7VyajovURMETcF31+mfIfj3ZYGBqmF85UsV67QFmEM4G9aLOdi1Y7
qno/78I4ONRsTYR6uSFDwzat1KTcHpulcOKrUj1daHMvOXimfI9utHOEAb04
SnEFP/tdhw4axQfxwuS5yXpVo0J1G4AipTeWhsBh+iVloRSVoic7GJHlx6Ax
337bu3NRqt7PvT2Xm3i0VYI0HoMwmxmk8aZTHxX8wdjUZfOPX3zSU+UASbiY
sRE/OMzWqo0dpLtxhaflqvsnyyvfG0ZsfyqFYh09q15HThLxlIZ3qVHZDWQO
woC2Oxz2hOGLe4xkE3BjdnPWpH3qeSvzDGqEd/cG7IOozG2wt/EqM8GUl1M2
FVvRKFVNQeZxuyor6m7XgxCzFnwROAQkzF98bxVZs19ilO9hyTDS6E5HOVCt
LHHeNrulW0SVnM8ikJqnv3tgrjjUeoZdn1J88hMZOdIg9ICzaQD6uJ5pS603
9dRnxapRNnc52gCaCPvvJFSn+jNWZkg6ZkFeWhB+Bd5HWXdoB381IC942huJ
YrNHDUVN1hhurjHfBR3x1YHxhRqv67ZTzdSolMwxuSD3jcMRaDy1g44jMjkh
L0v6FkifZhyeDicLt6LPsZ16u6sD/XFaQoTyJLKBlJKnSmxyqeS2OZSZn5xE
YWSOwT4zPvRaayVXAn5cC/GIaZeDmDCPmRzoQbR+6zexOBH1ojri8ZJfGXL2
M78LuiGKS/Tbt64HQ930JhYlTW8nO6B8Uur1+QFjS/VwK18Fs6HHaSHij0g2
9011e611HU8CgAX9cKjZTrs06ugarlH5p9HOGIdgO8ImrTlW7ubhzTVRrYy9
TmwqTMOZjwRxormSZAgSYvZUbSAQ1W9i/R8dNR5Na6QRe0FDI12HbV+3nnkE
jzUJBuvzUWcFRvM+LCIqG1fELUJuF7f3enkZYk8zJYpJSgVmpm6h/b1suKuk
jj8evzJAfXnm/CpDSLOBGCfF5ZPFgakRoZ0o1dh8DPi8xK27rD8KOZXbyXPt
K+qto+egqsUkSRF+gTkoDKWwVs8Vv/H6dPoM+MKKO8Tg9830jFnNl7q5oZQz
TC6ZU14iWyRVqedUKnbKjR5/xeVkXSdjpIiIpOKnx7mN3gyTcmgzd8JzXsdr
fJGXTLL/q/Afcr4A1Bxhf1qQ2Vl1yS/9CdeamEkZPaVr7+iHMRcRvLGYJi6W
R5NYr1eOdq75uyEDosUppYC5yIZeyIYkMcnRB7itNgZm2VHoOPz6CZBDWw9N
zjnVe28LLeEJ0hC1GQuNCtDmL9knq++f/7V4GNSAsX9Nmi/3pqagR51KUHvF
+oCt9uqZLCj6fTO2FHnm+gYwfnnL8ovoRH9fI177qs+eoshyhhj4Pz8793dz
6Sh4D1bn7bWBHB/d2ixVj58rjUnkTUmC5LhFh66qnhzoUQplZzKeRRh3hpTN
dzUTJnJjvoknwMyd4LbjlO1VFFRRiv5U2vHsxl+n+hduXICzzJioE66zoTlV
DFnkUCjyRRqtjptnLkKw5fB6ifOnXVEB+dOLxdF1dr0s9+KsSrRlPiupk/Uo
cbYDA6OJj5k4l49aVEnb8b2xdcJFzjZfzcJnhx6oi6GpRr6E5ZdrPUnS1ihH
EgMuYtinV+4Zl/gbiBG1DS8e4xnXYrcg8HdZrEwzNThh2bXfZZotPpP+3s9+
Z/1GkFDM6eBwFukxudQHfWnaBABNksm//tPBiLupdKKAJ5JnJkKUcTWS4PaV
oQi3tIida50M9wiyHR7I8IbR97Y2MkMAZZi2ZZQcshjWKxazlV4v25H7D3J7
xadrB6Ftd4LUCsgh0Cg3NwdKTBGxhZv2iHi/fMc8JXEC3CoOOmFFc7ddasya
/Z9xamlKsOR7/tMlLxxlyfrwDNGYAdfUDSQVRZGfPLULphJVCLCA+ut9pVVH
SDSqMR6uTydaeUyzwAw64ruxyUwZmq90u0xlpxgJqmwVtwdwPXJvJ4wibwib
NU5H/tqPwHXR1ZFiWf4S5Ev2ODm7UJD/cLEhp2pSgBP96SZqqj9lRt8h0dnZ
HQBWLrWbykeLtgtRNzwyjrh5bq3mWfKclHmiSt1UpUpmcbLa6lOT8guVh9zc
wEkIYBqUbiNdmxD/X67/C53BNoKEUAFqHTCXyFM7B23oM3mafa7dF9U9Eky9
pafcAFlYLpzVrNgA6S7xvt6ATXnIKfe6KeeQK8FID5OHtOfA4TZkh8OLurcW
ZH7Ua9nFQrImHRKgPVSxQrwSCjQ3BO4TXKjRXfGoZn8c5pHQ33/q3LzxB7NH
naW+sLNGeFXEXiaS06B+Uz7CsKvOySNWLBsENvAHcZisrN8CKnL7Q8uLo7uj
5LoBidzepwbodctvgKYROZ0xcItOVdpZD5JdLf4TKeFy4Kx2j8xfpHhlDu5D
rhk7h9YaMbjKJyXKnwrBVwB+ezEHauHr18S+N7wZoEky1FRt38zSAJ/elfeJ
8d26vtOUf2dym10kRjB32kuMXm8HLBbpxGa8LEndlFoyYeOLIKuqIz6i4cRF
WaKsJz0O0MirTY9JdeqDcFwtJHr2rqlhXVMvt5TRNBCDO2wuFUQYSn+TaXAr
2Izc3b2oPp4q+s3d7Xqhopik3rVN7oWcR6BbvSvI8pSzrZUG2yUi3jFiL4Fs
0u606ZVpB+WdeOopmbAU5hYmz5cBpIyVwDF0jcx8c4DIcVEMHtVG/XqTJrLs
ucxUY7VLjYpOeAnCBIPBgoxtUZBeOiaRDq6FAJtklxJLiGmYuKDB2PCKPTJ8
O4MobcrCgI9SVRq550/YPeMkHCpV3Jn+7JbHj3qUTh+wPhsUFPyIV9pkFh6X
gw/RWTq0qalcgC9fX4T16gcw3gb9X6JWM1zQMchgvSkIqbYVOb4ZfzhB6doF
wS8Gtp0efEf7BfPcYBLSPUbaJcZd/gMPJ1GtdRMrjERcJzsjL3Yg67a2VGFW
XsDaJcZdW1pu6ju6uayOUaE/0LK40nbXD23Oo+ef3c0bn72YPsYa5/urEQil
ljUDmMM7y+2yZRVTkn5ObGMJt+qBhjNyIM1rEmv/hzqgqUfJK9b6hOeNaDZO
8447cuGTKz8BJXjBU3DUkuoj9wdawZoAAIgOkTTIbaPDq7myJ2r6x0zZfpDa
ARy9/JBPQf3eXbUb3fn4MR0knMhYMHJ41HNPazAJzphUJ0eZfL/NhB+CfkBx
mO/BYQyz+lzjRYS2VLUt3iAnJ2oV6wWCmoo5N+JHGUOSlk899DfT1dURuoz1
wmv8ZIOpWIfAasJBzsLAMMXc9uaERF0vdx5XrbY8uAXPatT9BiSjMLFPSJhh
MLeBzFpDvCxJ6tYWOFuB6IOJ/wcpA0TdfC4v+q76qwF4M8Wt19Ks6+XsXrdp
/FyieF73ZwrFQ3nZNrPrTILdO4vFiK9m6crl8n+1BuhV5WsW1t5p7ujISbZA
j/9edevKu5JL32Es+tmZgj6qr186hNnTaBIfs+euD7iV1SiH5PKps/0/XkLR
TkmUho+YlX5I3KCPHzkntrduuUz/9nDqERoEIuHPwwql4pSUZoiT+a/nITNw
FCmKKTJaUx9MlBOQB4d3eRMW7uguT/G4nHiY7tHhSG5Gi3AVrMrs8vbBYNMo
NghC/gWYZduSigGk0NHFDmgei+eCdLNeY7/jtegHmqBVGQFEVe/1JapfpKV8
axD82kUXMQ4uaEIQ9QDGbicbwfvmd7Wkbkk2Mq9Xj9QQ0F6u0H7hzQBEQLFW
3Mf0JSipK1c1u7W25fKQka7VkSh0rIWUQnD07i/7FrV95Fj/KljKalXIJwi+
581sM/yRLBLBATL7FvCPF5vHMN13im7nNKG0BU4jJH9lOwhbL54kUswBsmYP
AQEf55oFl/f3yHkGqSuDcQG4oOMje9XuD22U2DjnnRoWttwogzDOvXgYlxWS
NtDL56z6hGPvORW1HBvaUjhSsrLH8ZY8gaZi9CcNtC2SO1gZdo3N/FKwGqiW
aKq3yg8yNIt5uuGF+DuQYfOWyaExT+KgWV7+dVJg6XP2kWdUFzBlvKBf8gar
QVp75q7wHLwaqAtaKF1SQIi1FSwsgGdMktsiievw7TIf6drQYfo8M0HzOjRj
qPcpz0SGELOg1O2IRh4Qj5rwPQcJJx/4mecWcfRwVzLYVzBkXKBpeiOaaqOP
b0XXCPheuhDBrVUnqE7d4I3G6usv7KvFeY4Vtm8lgad2MZ0qs4m/lhJrciWj
kLuGMBr8m5nNpdfqRgDAmzpS/7Csi9jhpU7y6q13DRcNt4lgZjW9PDNJGllI
eJLIadlQNvJo5OdjUYa0Mjc1PHUB8qV4DL7t+egDsC5PFjVvJxNNlGad+U/x
4tgfheciDhPvBt/3GDIxV6GeOMCkhfySnlLEmHf0Va9DctAyyA/Q2sSinX5C
A4mxG6b5TDwTEWVTE98x01lzUGG4Umt4w6W925uY+USbS4ojbbD+va7tn07b
TW1fokpBdqNuEAcOnW6EvBZzgvRYQRrXc6C4Cuqzm5MBKYU+g2z25XY0C4m+
fd41E6IJ57VuMtTi7UurJoeoW3Icluay2KrPK61ryXMgIbcrCFDraQkuzYld
TcWVHbSUxAW9CaaD54fKcAtY3ZowasVqED3dkSb50Q9DHYJVHRuxjlRWyQls
mUjrafz6En93fvODE6T7EYWmUUqkcX7hhB9tK0c4wWlk3DzMoLzGOgAulJH+
z8nbEDvaTnOvzF+oScZJJkFKOo9cB/zGoQRqLgLxvFZTmxMnKK86Mhp0DiLT
N/BUDlxg9xPE+8HOoPTKDl4dmO4BEMBXKj5TQq/gGwGfJRPKMWLWUAyzscoZ
ZOq4MrlT9BXuPmdRXCibXouMBi8b66sWNBCWacFYlarE/TYKo1H/J74vdhk0
lheXGWejt5x/yHKo9QxwEzhugCK/c5blQwyb0tBMgHDbM8LRU4MqlnRyeAxQ
rZSRcbuRnz3kWI2ZxLIaf5qFEt5WE6sACh4OI17Ck64CWZbcurW/w5Dy+0dX
7+EtGn2f2VZe/yyh5u+tsZxiXBjYSvWb/1LzKrfwPKlEYkcsZnw4W2VGOzEW
qz7QTW94lfpW2h1PShOel4iWb4qU0IxZz7pp9h8JrxSr02m9/0ST5RGq9XLt
EhuzgAaTlurymUVX2p8I8tymvcAt4hC2LZNrr9ZqBWe+KOWz0Seq1BpQBXh5
2sSD/qKG8/XiMbgAe7j20+QEVg3vnwQ0DJuLNd0fMfLdBq9MEF1BKyvPwjud
NNSlxLhfv0baoRpOVpenu+i18C4vSCGf0x4BNaPs+SpiIzT4S9QlZH9lQq01
KWkXewS1IX0k/6dL9hfPgf+l9TwcyF4ZM6FOjmOENHCKoue0ZHpMtb3W1jlG
u80pHIGxE49Pg5YxnFy2qMKTLBL6TQB3M4r04ASusmpTu+s7vHFmb3B9CEq/
av4g2teAe2ltDPutHhzsIkQwYGCusnFXt75nKcePuh4kZAcx4QukSaE3ySeq
mqnau9SV+S0zWljoSDsLYpXmlVxKkVi6A8C+dMFJNEBbYIcJdTAiDkL42J3b
t3QierNrhMyF0qbdXQ4fhsS1qyNdnPtJWU9BzZBIe8u7Mk0dVkKT/Jd893/l
YAiujtPVuMUkDbyAfwaXTNPsgCeBfJ9BXbz/xqu3aRLprGp9hwy1VNi6mDop
ggypSvZqxeeL5dX/auvKeVrA2P9wSTUZmFACel0Byl1T2PRECH4j4ntaZtjo
PF8eYKwM4V8aF3lDjOTddRSlUKi6r3pjMjn93ng0HcFaALcDc73qaI/pImfr
clp7OM6n7Hb5pbmb5sYC06caSmAUmbBd6jhx9vfHQIq3MK4tW92IU8aCJfnl
CBPgAaq8Z3tQicavJ0r0GLdGvxkwtAKa0UGEdCSchOH+NyXC/j1AexDspH4o
ys3Egh+56kI5Ntjqk2z5SkA2LCZetdE70y1nGk05vIdc+ybs07rqjA8egfuM
0RdqT2aCkqRfFV3Bvvnj8mZZ5DLH+lFJj21EzPFGhPcCc/OwzGxiFq9s6NBR
fi/EVQB/i10WqenAOLIebffAXi89nysYU+2h7tVBisWINo/8Lf2/mHKKgc9z
1jm0uRTUWE7lE3yjzRr7wfD8mazW4WyadcySkHQmaV0zIx9MAhR9Qzpwr7Zi
/162bPoNV1EwzFNwIq0wHgPCKavRe+zuGXC5WHutcYPZzp7m7zBesGIEp/8p
HyxJMTp1xQo6EWq/ACjn2vIhzwGwzD0o5zQ7Vj1anWCBqLp/XqFWt+nY2zmQ
nwD7aqgfkvVP27JbY+x1S/ls13+zVZniSC53ToxmnweCWaJQz41Xexty2b53
KZNdCFbfUBFtAu7rsKRUpoFznN6qZxz1RFU+aNuQq0f+6V4BpZu15jCV4zKy
R1+/J7v0Ie2yjuRehuuY7mlKQWWsnxbHrrvLRV+BqF5IM7rReWFZW15WpAIw
h2dO71BKv5M2N7Fve2CIPRIHvoHO/5RvhyRjJSG8lzb1uDCuiCdilS1Tugg7
xOJHXnNOZMgFvh9vQltLRwinpvHTpxH/JOGl7RQHyGxvogWLciVKjnFyBlH9
jh44BRx0UHEZLc9FUe14zaH1IhahtkeYM9UuZGVZEdERRzHtw1upxmANKxVh
gRjezaaFhBACvOV4qBU6b+9vRY3yCXsJagKPUjPM460KQxtsrmMwJuWithip
/Rg0ylQ51LMvjdGz3ZgVRsk90L/PxKfympXPmexFFguFGTR86kK4g7H5+2Hi
oBxxbI8FGcb5XXiy/PRkkTUZE7nqepqcHjK/a07NcHdX85n7AaiAkbCAxib+
xxll8vJrTQMI8K9F8fU4M/65i0lG1Hx7oyoZWgR2n8PUkqkrtVUAbXSuzVFK
g8CEYgiIl8Gl5wJS26ROUDHJvc81KJqb1ThFHhAqW/3ytNmDyV90jzehr/BK
4hasmuILj/bALBcBaTmcC0RlFUjj9XJVFuKnB5efoGHGlv51REKVuMkBjTxe
t/5ybGodHIO1HGlREGESYqBiBIM+F4Ig+BLkvZn4QVTvY4m8+BPw9C294bXd
pTERWnnyXRq2dcrBRPA3V8gdurrMBCGcaokib1gKSAJq4Sy4TokcxnkLm5QX
VeZkL70tM3cPZ5gHLk+Cm7W0CYQsjpfsC8SAmCrBS33Y377bxqQQ+sHmkf3J
J1kKRL09RxGMxTXew3w4q4P2snsGbwCnMxQ2ephr2YaXFREBLiRGvND3D784
hyGlavFp4xlX81yvgYqnESMuydfUhVPTA2M5DrJqnKu1pOZHP7LN8UtG7h5S
UIfefTW0DFI7oxXHjokEOoCtN8Se+4rLby6XXWq4NMGIXXQFPIUudpQzx+tj
aRc1dwLGum6GDAx8PE3tPW9JNz9utxALbTJZ3iykLsik2nQZ6HM60cQm1DQg
ap1dkt5ZQusAQjx83YJhQuI0NXjhCJr7Tw713FLInFzlc2L40lJy5ECWPDjm
+LEBFfrmFfSIaBOkwVw9jrSLfsiQLbEv53Z1grbx5fXtzu9vdzbsmSntmYtt
K1PzLu22Z8ewf/Vcm78rS14+1s41cp3OHzMxVTd+UCoweKgI4FvLDnqFbNhz
O4up8qGINVqEM4eOqkkGgMP8d3Y/4T4XKhHlhEEiIEo4C5J0n5K/fzPdqaXk
1SHwnJFHynZwwtxP8oFh1DWC0wG1dg/iITBrxcEzvpD75rVC3oGIS2yLxgjx
kL/tYAU2EW69Py+78lPHwRaK0gDyCjAV2T01ng8G5hlHokS0Me7C8yRx8/RG
oIIRE08yRmQtTaOHONoIL0mm6ZM3PxJe/Y8WdfG14HdSHbYMuzAXJLcp1dcR
NoJuisDiyt0vPhFdL0Qt78bi0CHUeMROSz17kEDlexcO4cESkKCvpUuI+UBX
b+O7eVw8F0fB3wXcnduaCMVynX+eRIyPwFoJDTw0CBoy3b8qLanmWZpqlk9i
dMnfUa2TGnm0f/VBszJpkOgwgMhlcIXG4Cc2XyHGU5MiBnR0Mxe0opRnsJHV
PdQ+gPf7u2I0apTdQtm2ZaP6fMvIoScDZNz2zKau3MWUC4cFX87AVET/WIEr
lfeZqDlJYtVNSX8PlArW+GJ6YmIyFSbqO2xI6L2NRG9TWjNb5nY04nE7Gfca
3Q/tY76GIHJQKSmCa28iQr1uE5R7AVwGWNwkc3zLF5r8vpM/H/wuOUxcTvZd
/EVdcNpkBqainNmvTR+hx6vlUJcDuvMucN41vp5xx5MJce9S9iSInbRMmwIs
ZLIs1jumqL/4B6NG18Tycy7ivA2l3cD+uBmJaKHll6SbZKixh4L4Kdrj1hhJ
DIucZZ2BIzidwK/vtebBfOrGnHd3IXj72s6qLa8TGiPZOmpUzOHwaLqnxY86
iv5eBNCbODSLYOx5OrIUHaaJ20uJgmyzjShO1QiWqBIkiFcB5OJr3YkSpCdM
W8qQd7BvF7zaKDbFEdfMY7anfMAsDKkMZSR440Q4BElpdSGUdwqEjyfGgm7x
1TsKxAwp4qzXQfcBOU8ne6PNpFzcjV/jK1v5teEFhNfs2k2pIH/DoIXpvk0k
eFhdzBq26NAS5FjUDaAyzrX6y4W+MSf/+TgXO0Aa1eilJetkD7YUbDPsdD+B
cbW+dRDxp/A0LGwrZgnlSBjTwb+z8uQ7rqKWu+IQFcNAWB+HeMu1IiQIWfjN
3xccZiNPUEAEC/gqm7iBBMWBcXaSu1XbnFF04VMrFWJCBL2FWjm3DrSSbguK
RirGccz+NCd95N8yZcSiEN6ux2jROj/8ko0Vcf/RjHMQZrvZsZEwdbs+v5fy
aWoBI3EACUe6cntq71WtGRXSaXxnxuHQ2cN8aKtvq4g4+3lMTcuAwfvvLcWV
pz1oYscsfGuRVS4q6bnSuV72UCkyJ4i4Tim+SgiDgdhM/sTdzIHVjAI9wZ8g
Ir0B//1VYPD5Nu8Y9faltmwwjVwwIcTzSlgb071k6qJLDqwg/Y6NISokXCi0
63Y6//y+3GYnocTOCmLi9TK5LgaJhHrQPG93nkCPg3axVk90uZSYa8lYj3ce
pArdLmR6RGiLfS0JeXC37sfownSrXUhsmyAPS8sVLpbRl4YXzpNUZvPwxs51
RiRsumHeKLJUF+tQP63+ktXwSw15owWgrtHjOlbRMed4tYlH2M55ZhzW8pj6
3ce4EyoALiZJol9EWK01cRR+wp/rNXtTlYAjSY+I4iHWZrN3AkjbfAprmpiI
e7l3QHf3b47M9+ltatkYb168v1PTLgV9pGYS1M4svKaop5A0LJG6c/FqA0Z8
jhZa97h74j1/7kAsGjcRDN4tQJRDVcq3Gs2Kf1JQor/BwDTmCE3tUKit0OOT
R0bYzLQRu5iZbPzzTdczQnZWZgC0f+TVx+/68j+PsjW+T2y+lrdysJPCHtbG
GmuafmB5EeE+U773158unlLXO7vHb92F5KkQZJW9EX+yyVoQtlw2c3978O6G
5GfVEcKVb+HioxmILrlEma82MTCr8ZSJFx1mA3JxTmBgGl6NCG39m6F1JLNc
KsGG55duRH+U9qFh5qucr8X4V7mzUuLxuBq67za8h3lNRygqkpsLOXZilUEr
BkqtyqXQ+4iMJVFl2Nz8yG/KhvkREzsU/FP3YbUNJyEpYd9X21FtlR1J6zDe
NMHADiXN32efq/pOFwBcFs7fYmRl/HccsYyCH81mjDPXCkyWbln3VzCNvaud
ssVwT4ndX5LKuifSPJ/aoiwgHRKfeYNwEQI+6wqB9TewS1nct5FJddXJ8R+M
Puu/TTwHDCIqXz/tuuOa6Aqq400Bd7c4sZgVqvENFf0crJO9/k8ly7mqjtDk
W3y3xqxQriP7UhX4DHRkGKkemnkOihf7puVmGnPb7FpdjXrC7fp9DaCfBNT4
/e1vloEcftT4IFEv5rQdULA41ImcG93RGNyflpxGecAtNcO7Wb2PQZQtdjaR
P+EcTDiZXHN/ElfINxOhi8Sg2cWFw2AMkSb2mUbQI4aQUpk02n5hRuOsDDgp
Xua0g8GhrKXYG2rvaATI/LFpqfSlrH9n79e05csrcPCtIlh+aG61UMuU9P42
873ZR7lFgQ39tVOy0JeVEH1oGaLG62CShwJcEgWfuF0PbLZqIDWhTqucgdBi
GYTyf8Q8nTHNgJwMWmUljR3M8+ULEuTpBdJfgxva0m+SpQ/Sq1Or3nqHHOSt
kPbYU7WythsjD25z6X9maLykR2pqsNILQQQ+gY5DL6PlgUral6AfflwvLoHz
vZObVD4sp45reeBcqfB2nDp6jMdm7Oa9XRRjP0zVt2vo+TAxzfAjovSC53NF
ywV6GC2uRKpM2CZLmJP3Xo+oJZssBcW/4SmUkw7R4ZnAuMzlILSWYR8u30LU
/JbAYcNO8bhhGXBMjuplNyBWrWmmRWlIencNGtBXOi9ldo+tX+J5RcggsbBm
hEQxbOeLSrxuEtl8sb4PrUjmMQ5HWvwvXSP9r7oGxgJavInMds9TSmKILaUp
8oXGS+YwYbkMvMOv7hWJdtifyFHZEMSNmVTzXGuDh3qracZ+3iXgXU4jRoJE
didh0cyk3PqrXyb5DyCy+axHiFt5CzcCo4hZ4Nn+dhCdBRfwdqP03mLku6f0
Zc4uF1rfxoSKYSF3QDQIGa+4orq8QucFUpOLfw16y8oG1GrAPE1klLkdcrU4
1g0dvbu2D78/vFvieQne4V93Vmz2UkK/qw+u9oj0WsZICKsTCSp+DRY+IbPJ
2q7bYeE5XlOCPg0PepSF8R/m5uR2w+kziEHhQQRGqu6Qa5tv/gLqJqy0dchV
vvEcXslPZe9KA7xoeilu9d+aX4CQ6W/I5qlQ2c8rCq0z4GEQIqpRuQBJp7hQ
8tRrriSWcSCBrpvrBLh5tu4vJsOjtLEsS7rx4YL3Q3wXJEZrfVDs0ywNBCtN
TRBnGJuuaSvfcNnuu1PqM0oW57U8W6mGZhOIAn7lln49uOJIHLEhobZI5txa
TtNpuQJa+Mu0utrlf2jmWd8R2hjtfpojykklqc6pqiqXACwYmwucWYDV3piH
wdaaHp86sJJ7laT2KrLnuvSMA1NlUz++6zoGZCvwMiKkFdEsxi+nzZ8Dzeta
VOBvT/MfB5Id/QyVXYDMdhjoPJoqX42meGulqkyURwSRvaRf/6FNGXMweJSS
RoGU2eJabe99bJAMHj1OU0QsznXTaHRL1vFEGaFsdXftznv15XPRNUSqG3wG
HknynO+0caFAknOADB0pSF2xee8EzU2XY7ZV1eE9DmNzf1QQhoNmTfBlfhLU
SZGWb6TSrGkeEnrQd4lLeWPgKdatd1GQ8yh23cKLY69004H66a8y/R312Ssu
IlnOZDSO3cFhaRFLfHw5M1k/Pppbx2ZrFx42jM3xv89YhKBJ2P8JJD7p4yKe
8d9e+ue/5uWg6FVWBRj/aNLYpTAQePO62vCQ7Tx4M67gvELHhCXV6S1/9nvh
uLUvbji4E+HUolsurHYhz9Xq8tM/HOOcG+zvz1mto1TxjQwSdQQZA+CSPY5/
nf1lSWPIp88h8iklsKfFyYRwpdcw+qxEx2sP7j7uixdKzov2xjjdKU33wQtx
4O6PrOVEXy9p53wUmCAF2Ct8fdEoLXCSqr/Pqyye++0G2GGhdAuxj0o7GXJk
tiRTopNr+YwrqhNySRA/xxxblwwb+XSexDVKsXpKrS/H1ypyHdNj1A5SINSm
X1t/32WcIKKcfs6ptsKeJJ6oA1Bh23ca/GsjP1lpunjxZPr+VWXT5YwDVYfX
VLSxEbcjtMBon73lJl6aCTwxM3rYmW4JlSoDdoti+XZHfb3d3vdmWqaGIwh3
YpGQhj41SHag0MdUf0SRF8jPW6BmvxeQs+webLcjlSiUehfHWFRPQCk6URXt
YYm0Colkh+/3F5niLzdnrDV0fatrUm/Ja2ATTOIPK+OmF9NkuGCCKUwaKAUn
tsnDJYA/3f12ZyNeHA4M/6dK3lZrE1icf1eSae0p/Rabi9N4iKf/4eVrkx91
hFNA+lCN6a5Nk71vCymKehvOQTkCzyJH1UHAsN4lK0SdQqLULpffwgjn+lsX
EkFrmmPEJfAqCr9+vufYqo3EkPp43EkgblgWl7uyT69TX2hprS+lNvuv+v7e
Zxa2S5NSA4jjqtohhkunE6kzOTjS8HjQ/8sd0c+VULqjdlSyLRO2YZbjdivU
zwraiypYANfOK86r8mDPOzRjqIx7ItW0/RW5m9LvuPAqT9NXZlA38Ih5h8W9
6K++EWc0d++f9QtnZeLtOVzXpGxNOF2IBALjSPRkhYks1L6m6WhpjzQc604k
AFkNSGFGkzQi1jQpMsxjYbZNfm6SD4uOemveY3lU21FGdMkYyam36oEV9sT2
R/tzgdzBgLjmKvXBLg70HFG8HjhAxdMJV0QVX0/t0hpo6PQ/5a4JK9h3SeKE
XQZ1TOPzGw3qgJ/UBHoiOEsMmHlgN+ksdo+I/xqwWc7GAxr7VYqWOhGamDNl
aluARMvbvHwjKSn0wwvxVPlzqSuucv2CDsANd6POzTT0rYUYkRhrDlUGjjQs
3NEGFOiKfs3TNu7XtjKvB+pAXI0RuWtRcL4U/0hTu6E2VLVHVdch/HC9+72y
u4o+ZESelIKKLi0BilPxpz4IW2vB35+W9zfZnY/bdg/0Vm8Zg7hwni0ELWy+
OorI3rPu3my6X/JOvU8m0wW/yR5GVTdpZxaq8/DK1pIN/xVeqBZruhuoa9Jl
8rYxaxAdH7Hi9YZeV31LsYjjXzO03XfUrpH8i11y0l7c/mEutA50RcObL26g
EbyfTs23iKekEwoOPsSH4iq4yeI8P21IqVAwdz7uEYX+ouYTITwxucyBaii1
BdjMpypBbGkZ4mr+elNJM1VvBIfj4Lt203HLJ+MPDuSDg+KX2gH3ymnOAM7Q
tp7kNZD4Kull5VtQ76mZ/+3ylhGyOlD1j35+0UhT6BOWivZIm3nGzmm38cGr
qnrwiTHwtX5+8mXKjkwOnl+inOv76vkxvAVN6YtpYw7kjajylX2hRwL6pfF5
I0EL7Pwz1m9pCca+hh9U0Uy7Ts16FCfJWe22PwA1O2hDzRB10R5LQfZaWQGp
uL/ovTLdkaw+REEBxrZ/NBDVeGKQufEhhrsbN0pyUEWWAevKiZGBnnA0ctTU
Ftm1btLWTrgqGVU1IjAjj85p7teQ+Ai03ES0sSyIQFXZhwKLtk8PR+AIncXr
ONm5uK51Ipvz/8mivOQptI2rc0v2ZqyqADoA6SGA8awcA/h2QA4mivQ/urHD
370zwHKBVAuZmBcL1tY1NBUZGcWER1PCKdeSBSsx6FBxO3DQ3dGE/hCQhZlD
faPN5A6uFHlJ8M4HZkf/CzmJ1SkDvFTKt/q9Kx7Z7uviZKRDJLoeYoN9Vysh
uymOedHJakikwB1g79IC6v0U0KORNO1XjpMGGKw7wQrCFWTBeLnYTTTmtTED
O9IZvjT+XwpHxASnAU0acoTSkVPoJ8MqJ1ShVprSKgwAFMfsaxEt91o0o7GN
pQ7eUaEmYmGUAKzzBaX5/SWajrSUUMH4Xb5/6dcTfcl2lL+XAdKLnWwrwgDB
tRHBZpNFPlmSoJRINoHc7hDVqFl+RJmjHUWSYbxyalhFiSdsT0JSONacJJ4v
+Hrpnt+Hu/s64FRAEzpTTNJ0eW23gneZWbCrpy4lSfZXVWeiHBT/3A6LoPEW
MJQmnJBu5G1F6l3YUPaD4gPTQ3zc1sfNJaanOJYqDebVLU9Oj3nmloOgmDmR
fK3ehhePW4QAnbePyDlSuUgs5YqC3yzVPl28W9XdeOTi50T8yce1brfQvUuA
txeX6eisRGTvRBa8stQGFC2p3jzc+VXRFraty9b+6Ctyp99KPM8r0+VKlXH4
6sVSPD7IChSN5YG1850fBkNL6B3rAu26/kdF2T1M+ck8IUpsSMvnCfSqaGnE
xVqwUNw0YYqE0WP6RPM6UKrJIjUZ6CV7bybztXqfqKTj0oxkmqKAGu+uz2HK
aRuJhqPEbs0GmKLwRaGnWnD/TcaiANzopJCIjgqSM8Z14VjFj/Bl7UcmD0g/
P9lMjQAFXkGWMEZ8BFNofsavhWsXloBIi5przvqv+NpL389UAwWL/VVkJJG/
DbJVpH+6p+/7cy96Glx/AwQXINcDpYJ08WEQ2MlZ5JDTldKLMKN0l+CZOZiT
znnXfL+vKV1WkaNk42fHSjLjqMTY/B2rx1zJvdWuIpWrDkU4Cplyfsn/FNnF
TAFpbqGFTsjYbDJDH4XjLHOagXZvFt3FAYC10zUA8acItmwNtVkmjeAkpw1W
uI4cPs8fA9DggfvhosMZ0G2A1eetxZAps7XgxCN6Te9O3dj4n+Hd7ojQ3y9M
7g/L0/z7ULlgEcu5dLlpZWDVPC7Qv7QIsqq1N93D3uuJwsD0r3aDvRF5Tt5V
gGEXgxQFxms/Pr78avxhsQCuwUP/jVd7lTpx0c8xR790/Qul3cwW1wKChgNa
g0zDAF8FV51fQnh+mOJjBjA3ZmU8P+G29YGVVWtyZO3BB4J4rtZNAzbtAKaM
kTCiXFN6J33oKJDsOOBDEDQoPEWjTH8s1O60ShMk42mzOO7/bE0Bf/JPqhqJ
1GZ1hjRaQK5BAS8U66F/KTQtiaVsXJQ6CJZ+D0YS5Bc2OtxsLfdMnzctp8Lo
ejoAUf9sQZFJPWFRXVW7dOHaEJRvch//P2w4D+fcQcEH8/1DBLeTFctrxS7t
desfirJB4zB3/cVne/gctD4LWwfvGRGIXMXQidkMiyYvLc4rMsb+/7opv33m
8hYkv/ol5lJOwdRzyjyoGZQjompK8pQ2MRlhPOEMS7qDbCHGbJnVx0gEnUN+
KmohtdOpwPHw3Yll6aClxT4pSSg3LQVkDBGfQc6diWW7TkotBtbHV1WdS1iP
MlIFAwOhIys7lGj+9Jf9L4e6JSsVCyfHp+gQO/hM6xzWqZfcpkJ+aCm3/h1I
HkF0VkAsOpirn0l6qcyrgN3RBhjqpFi6IMs6edN5QhWobsASEOEZmIyZSn9B
SJPsXy35X7/xM30kFSaf8Usi7Wi5L12vGDUFhMzs4tAxIAwY+LpzrbNOo3AB
Oxba/GqCkmb/aBpO5MpHMkygsARVg7IS/dTZd3r8Cklmh6k7YiehOS3r1UI1
zIayyDMd1jfP85UlFsGdIg4p6NUeN8ESw6n/+nJSTaylwn7ygYtpwJyDkhTa
rZp4UD+SJ0OO7Iz8teczlpVaxSeRQCTs0KLB/mK1MGhOZJBii2ZCeAejwO0F
tyB9oO/+mVBaNoYfCVeMOKDJ5LP6ZJ8CFR1NwJfR0g5Jg+MACRBGHSo7NBBv
cjrTaSTcjYn3keOA5X5Gp6sV6IcPa5sSH1gaqW93qyt1Y6aos8VcBHbwlFaE
fmdzIyig2lZ+L+3PRSwS1Ql7CwLLe3uzgn/fI0lnsk6XQwwps+g3FZDFIVaf
J2z+iuylnpwDphbq5w+g2Z17iayr3kGDajTjBcUKjgyqUMHzwfrhFSRxQh5h
5Mx63ybykmDSu86VNsPvubbO+84lSzIm5St5b/4si8F3K7EEhISGB/f5oTXX
/9indkSVgWZYVnTJwS2xOcCx/7NuT8RLoIn0wIpKjBX/KQfBv+qBNPkOl2ar
+B1GW2HtcTHXi8zAks1BQyRRxuwmDGLHSG6Azq+lo1slhJkd1n75w8qMfQV4
nZl1lBn1HiKoCqprSTWok19qo64EDPQtn48V/uJeEcOoKjo24Pr1ht7of00E
wb3XN50bw5QQNn/ulPllt/Hpc7SiLaPtN0MJaXEA6OB56RIZpOfStFM0H20l
V4DhLbL8hEpVhObkoli5eZBL69EvHFMy53MTCiaDpjOmVcjMFoTliDKJsA93
YX0FkSNsMF2Tj/QmoJptsmATvzUZ9wL2p515falduTOtK0z+EYRhpK/bC+Hn
K4Jos64cO5yYMu5j2EvyuFkSQDtTezBUKrlFZAY+Skka8nLvJZjSYY9UoL3w
SuOtt9wAaWG64aSFOH3m+iGQ6p37aqYghpQJUkKehhnoX0OTigj0N0zPzIXM
accYHvzbiZFxcOn9wudYjUDUPVzs/EfGOWuy7spuq5+58wuMsYjynDS441fa
a7+qJtvu49Mv8Fzip6/kwOKGESPis3AjhNXRPM3+8Hkco/OcZGfHhVTpVPsd
6Acmrk6QdDtAtbMWl8vJdEvq+NvrTpzwyP8RE2gg13EqUGteJDwu8NrnN259
MPCLLQUWNeNsCtrCKwjbZmVXb0rh/YjGL5lpI1QHZwMxULoYCBJ3AYIP7ssh
3tY1cu2BL3tvAkukx1zBBqQSnMG7ozoarJQmjqcLzEeffFHr23Zo0Bwj1bA4
cRUt1ooZUGlosf2KMkc2tyTdkQ+f8SIq9oeh0SpjwBvk5C2hjfxzKCYBiHeo
3+3J+j0D3rQuxEl4iRim7eZ54BzVw4QkgLF/NsrtWT2aQvqm7jIm6NS/FFiR
jxbnoyq2ZfknnomAn1+JuSJO8HUI2I1orjsO/Aw29x5GwcqoHjj3GPLKJ5VV
oEnx8LgfUgDV8GUkK7H08H2FNZXn8mSV94c4/AS4T0g5QdC4HNE70jzQ9wLv
r9Noa98pXd6HYVRkGVYSC1EvBueCEgVR6axf5fuA18aP4chN93feNJQ8bjF8
i51ZMV03H/TEognnJPFffSSrbHWycyAzLuPP1AesF7dx/BjYZ4QGoLnsapdE
xenMJ0Qsuj5pQfq6Is0YwoZzClYy8PAtSBl666KWf0fOVtkLSXcOz/u/c+Is
QaU82aJyrMUZE7ecwZIOER51PJ3RYfT9m1oja7D+NLyznVQ2JSpA1y4bTqFD
D1P/FouYM0nRdNOclS3EBzTJDy0kVrezOsDHSlby1OXtQSZ2Kwpt1XPSGn01
vp5UCOTQGuOckUwQARLmkE7Vy98lL6T9oxMx9dswdhw6Cy6jHe3jxLOwqEPm
bbogydoAKC/ATPlSgaG4wX9Fq0w/vCc/l9nQwb1dLiXCyMvjHFL9o7R3D69Q
5DSp3RL6ebOuPmK8aNw5fgj2b+8BAe3j9iOJADoHuQEOTATioFLZn9CzMpV1
V+oarqhiK/7l7RvslKHCVlPNKdMDr0sTrFOVJb/hD2WJYGy3WUSxdZMhT6sz
MvywsHOm2vBCMu7vL8TVLtOLblbRxQ4whUK7w4d3z286P3Q72qDhDYodhxG4
Hxa4HQJjzmaOJKeXuPzt/3B2tWRGgEZ01lxhBD4yGppY3aGXxj9yPojXCipL
QyTmwB2ZVn6ngtJ24BvOjnK2ML2RDb5PG49ncBH2+NOuCFWFeSRmLib7jCzh
/42s5eu4cd15D8fkwcx/gd85Vw4uUvNA19nWRWmLw4Qx91a3jbWp/k8absBH
7VMC3+stu4NZTgLKt1kMeRsZ9z4JDNbu9U8jtVTNdurbv7Kt+Gj7mbqePfrV
IXjMlcKfv7VORulGMTv47DNyzJs/Ovg7GXX/cO56OXVIIm6gJK47/0ycXoIA
Nnfg5PxnAvJ9bKBgTWvvXyY+mXRdGlq66CBV4kLVO09pEIqwwOCxP31xjD+B
UltMnqH2lfoP+RmPn01hQB04BNavvgtShmJ45jdTgszaQ1+FsLuRthYnitLD
7Njs9FDdTlgOCsk9JOuX/kwlcnzb4H2TyMEbNEwvUANZwOEWkUqz2yKXJ9S8
CnJLgMt/2m0bTpIBVaw9yA0zfBxGcZwiGl39PukFStWAjf2Lz6j+vryC2slT
1tu5pXgiT7uy9WO7AkBLqRAQVVSX99M3SXRvPGN7dJKaBTp5okn+Jsyv6OgF
4tZTDK4L1ReYZFmxCSfcndH5bPiwo7CETp2AMCWBRgwdYcjUB+f1ZLZuoHM4
s7D6u6hHov5kkuV7Ha3aAOH+N4eND9LZULWUafA72DouOu8YizkzrBs+ADGr
uuzXD/bwJ+jnJayN1fF2JYLv04tauYXWUyHbVUp1Oi36+r0DGb4nIsWLA3ld
vTGbPqqOtJVzh2RCHROT3SZ4gmmVI9DAWvr0fcR7Nz1F5+NCPTosnZQrJ34O
g5aDaEVqScRTBnQo1pM4fX6yUetJg2QqcXy8Lg/H/0fHUFZFbZh25wCV0DhB
mKfC82V/Dy4Dpc4FZksISreISfKXug8jpZQDQyeYbwL++Epy/bQ1MGjaX/Sc
q6vFvk99jgslNMTvcsk3D/BtG9fD3uIOyAMKoshMXLIeV5bCDH3RBi9y3iIk
j9HhwdMoq9TadeGyUHJA0E3AAiMT4hiKK9ravDBqFSEs1DTdRLqTS94aBjEV
DrBaGc0aVuStWcafC2hKvtnU8SF8q7ITBZqtoqUc3Q/mkaQ9CPGFrdmLSowo
gGEP/29Xv2Yp2mWlIse2lQektwn2IHZgdzHW+GSeYc+8C/q/nMcWHNmMWVRv
aKRxAPIVbarmQfDK5ZoT7Ff1Q9mS3CB8ZVt9H8lccShidzF/3iHFG09uELxe
koS23PAuKFTOWTeHSG1VRU/oi5ekJTyw0KD+xoQt/KlKiur0flbORaR5hkES
4B/MT/yTQX2wods3s3abHn0lkQ41PTdPHtDfjBzI+idGGJs3nlcpWZhkBPes
VUCMmNtV04EPFEAhe2iyhIpDcstzuLdZqvyMm+v8+m1Pnn/peTm5CnpJK5QE
dGFDiCh/yiqA0+H7qD7b19VKsVNFwJrXQX9l6PME46RI0vOodt3Hy4drWNNx
G+9kmQoLii+qBLVPHNxLBV++Tr6EsjiG/8EL0hIwcdGq46l2J4rPSr5ClfnA
p8n1Xpk4KUre9lHv5wrP3ETHInzyRnG48W4062O+UF1XyysxBN6WsodHml+q
HX6mWM1MRI7DLouNOq4Z2cz81FsAtyHbq09LdmmagcJJUAOfT4V24jLlKE4c
L9KrI/JW3O6FqO0RvqQ2iXZtp2yfQJZQZUJn1vwtnlPHetijHfN5ahri8Y+c
f5zkKYqMuOlmAZU8aW+CJIW3HMYeu45oQYGJka34jiOxRwEJ8KD3CB7qjHWO
BKMPDW04lQVre/hnA/XRX3qKUtrnERf7aRzTi+kGPLpreIjI4CV3Pv/lmxxq
F3fg8k+w20xltcdVbw15RRTaiAOyAaIq/Gf1NwTxCqpx5bkT1ybz5wqnE8gz
A8AucfrEOrrpNZ5bmeurjC8RozvIAFYtf5wef0BsdcuIg84pK+qBx5ir812+
ebNSJCvWiuSMqaDIl1kcVWwCwjW3LDffEiY4QYWw4Aaml8Qv9OaJACgyEfTO
uvVEKnO3GPWwwtY+OIRNNuATbetMSAd+hcAqxk8DeeT9KFBEJHNGPD9tvo+l
vzbktNm1/aL7NEMKsSEquC+c1e12UjcTh3RoOC9UiCWu+I8zCcjaTlsVr7Td
24QwUvTz5md9xTWBPp8ySfbJwwLXtydDFAfnDsG8npMNSiWYjmzERRCY4u6P
NFBzlSJAvOZ7KVtUQCCcaT00MEGZ4juNijId92vU4Dy9Tvr/xtM7nJCCEK5n
7/Wt+7gij7QtvGozrLaWLMmyTl2qrZjRY70PsCcmWgXaUxB+t0MQq3JySEsf
6QgQXEbLPuyus18hzBKjVKQmp+ffjY66/ZW3QrfzRexkuFi1yqM83Q7GW/bK
z4S3LXeHnQ153EbvgTsHiJ0GBiEItlHc3YZoAo85u3W6QYguOBZzsBW/a0lm
jdZfG/aDHlDnOVuTHGnoFsFForuxR5NXLKxTtl+fD5SfpiQWq6TO9FdesdXO
SBwoBeATdILoqlu3T4US38FFLv7tZ6QiUe/cMjj+Nssng0gRpUmcSBD6QScx
bzg7pzxPUxr1HIDMR1TAr66zCgeIqKbj+hz0+eQPD1iTh9VAtDAwQGtMt86k
hKra0/yUOGiNLn+Rn9MSnXxhOzbWZTM6Lbeo+16De55gXfnD8c+lhCm2ZnSJ
KyN0Bw+/MqpjM9a+1JSwna6gjyIyBgxh+abt7EfTM4P1CVrHC1gSu77qZH6H
I+Sz3mVg/92hhVW9us3eyEIX85FPDwirN6kzKIknq2aGr54xMtXaJNYNyxF6
2IsuX5AqSNzQ05ZojbqitTRSYYzutw+mNeirKRRBHJcq5cCGW97Ps7m+dEle
9yZRUGWN2u3zso9GOLUhz8p5ec46zbZ+yaeu7+Vy9nI9JuzuCOyjc2E8659e
bACpyigw/gvsarz9WumQE8OKA7FEfq11KAqFMhKFyVJ1ns5NQSo5iHZ5OCG+
FcqbRiLpTD3E2BXt5CT9HsuPKWkC5BoKsGu3EE2Z2yFJcu7ZqnM5c4injd6P
UlJc/8WDgnmo8mKMBMH9xayJ8kKeXHIdMXEJgN19ToRqReStbJHqJh3x4Lq6
AsuCvGXaKstjSabkoMO5VYRjTxcd36D5vvi3LHaTX0eTNK0W5UFdYDTLmzvw
SO8lGaQxU9zhzXGOp4xT6k7Hu2X6LIxJ3p8rHTXlLKmgwA1hLoy8oF7jlXdm
PSCc5YfXXbxLhuSoQSFesDS+SC39g/mko2GyYTWnCTiomzh//ZpMCCP6oPxb
332XpPironRIrjcpnqgkWcTLPsXRJSlMhQaDPqfSx+sJu07H+xRMDx1vIAUY
ItBCzOZljoFpqc7d4EyKCR5PY1p0TnFfwh/AqJJVLCLndMUJz6FEb1duXO9i
9PEGPLu1GUpaE2sSSsdO85MrvY8mbbC9QNCKPzS/Isxd5uUw3184nWZZYYwE
AGg7gB6uURq38yt12lLyuJ6aCXvbzwKa8A8QKbhn9PBfprWzvQWyYEHQ0RBP
xIi2/8tOF9ssRhm50tqtCKwgLzbrBh2TVPDszw11uv9mh/OoYm/hUsVLAWYH
dz0kIPFQfHM87wr4Qya140W8heLdXC03qZ3w0m7ohU0TtvGcz6x8zwxI4I+a
eI9iYxj1s6wheaUGH7HynNUyqB9hz7mjiWJIZapM176BRNkA7ZqKmnwxI/ak
ooWR0sSq97do04Q1JSiOA2ymgZovb2W1rBqSGzEYdIUpoIV1YD90jF4ommw1
zk+D9AHeGUBLoSN0xPxOvLliJsdEX6V85gyeTQMUsWx4PaQw1OmJKJN2U29S
Vociy7n2NfSwP7uvVohebT3RMk7SNIc2XyYUAolCVplVi2rTfZxOC4rTiM8I
ycnfPdyQw9wi4HJX9f37BMiY1G/gzvlLunbO1sFGNGPrCv3dBXbKj3+mVdNI
HwfCPyr9WGwCe8DLR/h8ez0xvmjVaBRHGHgRVcPhQaFjJ4E+HAMpBX4gCyzB
2kl88LEbY9iDRtqkZIJreRfho3w5ckG2SP55hbamwuevO3yzKUJg61wKPnpx
X8slpS4zZN6XN2A6Xi2dCTaNrtJSpDzVRlIwkCVNea12mb2cshdErq4lfnMF
ZuQ1sTKMIAa5M13T4wob/vo2wBSd6cz1D5QHlV/B8RT9hNkTuz+pNroSwo1M
zWb4U0A7CyP4qN8paWbByf+IZbagCE6WaRkPwA7kOEATTlakZj1WVJsJIMpO
LaesxnF6O7YsHUSSgXUgKmTT5RZWY7sqMbufiLOZ8xR123jtm8HPNs2ULHiw
uoZNpTCyjjbCeOguMfWmo28caEDaAhOt7hjTwvSXFsnLBHyTCQSOnEYp5M1D
C3EmDPascFitSoJokcUCHBssWPIgd7okpwo/HeTCChKo3UQ1xgGtjXByO+GZ
40b0aeEVeY5l0zilbNEQQkF1YACk6vgda6ekJ7CZHjDq8/599jFq811RTXeX
cYCLU/Z/oJTndNCVvMsnFr9jHca1UzyhxaAQ5Hw71VQgXqLA7Q+Q2NclfxXm
AccnTdL705fUsSvhymVYZhdq8r2qbqWAYCt/fXGxXixxNCvCk+wZlJbRyenl
Hop8+KaFJ2unhKNEGB7NuwPxHFcwUGziahvC31msI1g+o2Vyph1hY1FdG40w
wQAxuqxRkhVgEzsSL41JQBGxVClWEwcPfYT0Up4boW6dw0Uv/mn532Nmpfcd
tyAn2aXRmhY0I/K7UWa228LT1zVmx/cqbexxzKgmIYgLQP/GTCeMjWTcfzj6
CKa6WhLgP7XwKtTB7RFOmP6/B66m2wXMOfTG82pLWJM1AzKCuc/Lgv6Eh4DQ
xR1gSJNj2HZMBULech4OgE/e7btbkUKXUsBhQLOG5DvWNWIroKUUckXR1rOk
/7iJpH9YCnnXg25G8/n8XDbBUc2VZIi/fIyg3sDpvrRgjjmik6aVzqC7BcvL
poeU0C6S+j3fhxvQxj6/+YXhHHgYvvDpOAIbF76sbBt8DQLiRm4zkbBqccly
hHMedqmY0wO7AfVO5BzP8AJBYf2yV2+ZHM5GDUY96fmTAB98/izqS3Nudgua
x8WJ8oGac4Z0afil214tmM6A2W5DZeaoSYQsZMK77UTE5GGAi8QCFS6T1y1h
TD15o6RxRvQBnH1KfyERbH3qw2lKzzksjzSHALP+L/l+u8+HvJBD4/Iz/HQW
dF7d7G0vp8UQkuIRE11wLiZn1nY2ouRQaNAr92fQ5RYS5Z4OlPN9jjabhu6+
a4swC9ulQd5L3CFC2dm5EX0z6Kl+vBYN3GUbWCVdupKncDmZ0F2JYnRaIsdH
qQN8YOkTEfjVuOl1MKIO6a4f1oHVTKYb4gGX5FeK/lS/1SdNQ49HSXWQWEld
A43zeIUV9NTi8zEYAPuyHl4nqYHNhDb7FswMLc5O3UrYrfKQ4yM+jP3lfWyj
sicg2jToAL2+28K9CNqOQzt2w5Co3JGT1VZluVdFxUk81A6yutI5L5zG7D9f
aziZhKTHgEArP3Emenb4AUY6TwiEGh453EMAUFYMQup3/h00z8JLjbvS1boa
zxjyHyVX4+fKlBHCXsltv5Z/6LxStpFU9mV+hmGupdoBaFPBpEIiGdyi+gcY
UhnuLjhDxVrPtPFj5c1GTqEtbcZcGH/qTSVdlHSo2oZ7+tjWKPYfRClfnsNZ
k0a4EpXTNcVdC/5CYSmhPeLGOHN30NxMTik0jhVOR/nm1vB4yQwD2xaMn45B
GAF06jx5sqPmQ4ABiYVTaPfeiPSiMY4b71P4OzuoZQSM+iAj+3rS+khSMxLY
9vfNUyw5JQcCz8HMtr63yg6M6gYyXljfzsoCqpnwmBs45Y6djmRls+4+bWF1
lj5X93Xc8OBnFb1z1u2lmImBSf9GNbVD1LsFBHb+z/4/S87UKOTvd8WfSr1d
DEVDi03veY/nk/blpKBhP7u8jvdhjqrPbZDdxRlHbDaXboiIGy0JGNmVpQ7l
N6mcKSRLIR+WnV22WrP7WDSb0/Ulm2Cry/WP5JBgDl6aKVlhXqDEmlGgGLvZ
9UUmas0wpWHv7cWqVZqKpw7kgmi4baYSRQa2ITmXEuZr/eRSWUfpUpJvkzuY
PkoNYhBYvIBshO2WRDJjfhGDGBmxRSbvexruAd69+Bg3hrpelpyFBObjmM/l
F3sr2UhDA2vi0Q/I/NRr9Vt3FMFliaA5d2vxkQC+oJMxHkJ/gct1aq0kWzSQ
WPR2ONXSwG6sPKOK8DoR5fecC5mXFKEaizbgT7rP32TE1PS40N5wuj86Ife4
DgucMXJSxJtADrJqPIheWL2rMaUgzhPzfvJ1d48lQd+OqYMz8NjggCAFTvLJ
S5sbm6uoz2T7TdkJyNgTVD4rz++LW3rPKOn5SG2wxarhtTdMsRVqPtwk1Hp1
gXEolN+dJ2veS+We3C2R/Ty4KnOVVLp7RiF4hByRKUAXFRXyhGNqE0vocPMZ
q0xbxecX2dz/+V7AMAS29EPbE83FObAAstNqeVRdXjHBlO45lep3WxLp08VW
5/AEkr6T4zgmt/1oy3uR3KdIND8fqjYiLFzKW6gC9jhUwkHuSGzMSQI1aiHI
W0bfuA7a5ZxR+KjuZfXY2yrggQQ73TWBR5M4qff+1W48+wC3wm5jQfiAgAbS
7iOQg0GSs9xd2UG8EFPzHUc0JBWKpVGVgNjsO9b0XFdwOmW7/g4rgwmNxUZ3
iIDudjvOGDsNTVVrABjdSBQ54TPhNxVL1HQ9htR98ZKg/pideDJ3VbTe5++A
kx51rW3z3cPn/icc+sZ5IrBaNcrJRuWZ53trH0TBMOReav1NENrKjqQdGwtB
6wirNDCH1Px9gIJleo5IyoI47XPLMS3Eylcdphx6cX99h8O+emyRkQBgOwOB
q90zLJZRHcDxYs/7oAvngkHXfKPjuUeW5W+v4t02SCQHgvPPp0OiTmmhvzko
i7iBTpDM+lFsm3vlYUK3UHDrj/U9XQu4gNmx9wVsXg913m+YFdLI+u2bZij6
uuLAei+dLVbE7+mH8YjxBBSEOk8xAea/mhXZxApypRoRA2rSJj0UTpv2AaAp
ZbxqkxJyd13X0mfu62wayfiE20Tp0zz2aXhgq53Ja1kGbMiqHqBiNODeM5qy
/3WmvlJCRsTQco9727MYWjJJKh5/qjNj2VjcCSAI5EL6WbWoaJn4bUOQr+2o
e1erNPXBo/IaNZytvgFvkgGy9N20otawPjuuLh0UbNgSV9IlKRmzqt3VNmS6
SY8oK18b+dF9QhLEvBVKL8HT+bKLnsVMxz97cXlrhXIB3BbCr+joeiaVHz1f
mvneCyvGraOYFXIu9Ji4W4ZOjo8lgjDQ3nSDlfFdukj5VAvosz9VUC717/9t
exsQYq3ixoBjYkqxfpvgQadtGG1TRDCB0NhpzcLoh0pVqTndWlMX2D8ltH2T
3D2qLMjloHMm3uaha/TeZ3IhdzAYsWjSGQSK5nKo9kRYqTMB5R+degLEc1a2
917SUp0ohr6N297etD1lIeJxFwXlTJ1h4ncRclaJ8loNUhlLmkAPNKUOINau
02emUD4JurcxAtJk6/md0z/oReyOuVNpGQ9Hw7b47Zghgb2UXqnAKSkISira
rhZqyNhYrUCl/Pazk79zI+nv+/aWx94ms8yw3e2xx3da/PSiSkpo64ad9SQm
jTt8Wju8qPdQC/w/7nRNTkKnvDjhXfHC+lZlipD89AnLO8SeyNGleq//gS0o
xzOFa3altjCOSEJZz4UkEntpZh0R9Yfhl9Bo3C+7rU4z3i7DEepTotdNyUpW
ziZb04KMmUl/IwuwfLxNfKl0Zvwu9M1WvMpzHALQ5GZhLM1EFRtXL9AwQiBc
I4eLq/sWBweC0IR7y+kdW7+lNR8xxYXz/OyNaYeMGVL/XGuMW4FY3HM/Lzcv
R61UdvNI0npjc0wdtkivUpxtxKLau7hvu8hJ9uL/1vpVwgO97idne+E1hqIP
0IgJro34r9FTwO/Owvo5MnsKeW37QcfQBnI4L7QeDJ8t+d+avlroAzjTJ6kk
HVCFQP680MnhELRe6BOTDk5YahAcNRIiwJ+TXKfPs+M3rd8mPNzY+XTlJWRc
OEOjrjQ8DtO63c4DX9xX1O4WALJWPHpHT2lmDE+u283BHlD0Wzy8Dlar+uWO
fSUVenXaGL5vRv2mufsdANjljlBbd9S9O3wSJaH78VV6h9z8GZKbUhUkCDsb
7ymzn3n4Gt5DwBdBNQoDeBJ1W30fN+B9Lb8Qf4ZEJyBdWy5pp9zFetJISY6F
EcOo/hbvecTzsxrMMxaLE7o7PZU/W50aBtQLo/FLdWuMZobxMl1s7Zr9Cak3
p0efL7uxg3hMEgtBDvcISUof5IjWjyt4/9UCY1GxNX9wfv3nRiXG0gI2Wi77
TprloBhos2mkPwWl7BEwkAI+15BKIjFD6bDIysuxutcYReZCLrrA9c1QkOEL
28ctjl+oAZ6r/UMeEDcLJMyGd4a5Iwt+iv9sFbZBZowTi/48pv7AdRfEX2hd
7xu+JrqV0rRslMEGJwcJUF0yxCkRdGUHS82KdV1ezn383TxUeeutuhO2l/fK
FkDjZkjISvZEuKz4jM+XS4swSJ8RqA8RSsHVIZGAKSycUAAGkB7lVrsJl7y1
GYWnH0itCWq13TTjp0M7+vtaNqmOUF5Z2emS6RD53lEHPbp2AjIGzrrtihhp
jkpTQZS4a+kV2G3srMti2+OaSk25eMD/D2XdvUS1oxVzv8RM8pp3DcxUMsJg
6f0JCHYFZfRu8B5a7GI3c1NA7EpSwag9AYwZqFJDQwXWtp7ecQU45prsw5pF
Yzb4jKyimxsPDBqihmvin+GXlBxcAu7KtZB4PA8mZYrnGLLeMTPw824TpS9s
Qj5230kTcQkmbOt+itVI5dL6rBC+T804wzBDv2koMhWTXZ0jIxko6tLAdMST
kEiRvYan/Sb1lTgzbSZFhslcDpdzPwTED/p47BONyQfkVDV5T6HxfXO7U0Vh
JHQIifmQd3nhPWgITjDHiSyBe9UcI3CPTVbHhN60KbqHOx76qbr/QYenE21q
krjLahS+SHLWXS5yCaWM8uqs2nD4lJByEEDerMVDLrcHKfUGHWnn7x+GUdGS
pe+l4Rvnhc75tVCHmZJhu8Mm153yEwvvjk+WvAuWY/KmHpR/8E9skOFB6NNt
iIClW4mMYY3Erj0EUi4zEMb1c830DOf7ekS8Qt9crXh0tjQoqcXhRY57U2W+
YlrF6YJOSaVyJeWVl7k3FCr6urNXQLd4R6rxqUeBa3IbzMGaLbFkiYrDyS0I
y2wHhmQH7327cGGo0XPwtQgo6Gx5H7sQpEdTYGjT0RWUMNdPqXaygBjDm8El
T00mQFnjwl0u9Rkd8Oyip6zJCXUzZ1genXEQnMtVLKIWfH2wTvWUfPE3pLX5
MLTsOzRIxRCDbpEtRwx/+IiJhlLYg5L9+gnfEmo/hHqEk/cqWuFYzjt4c9RO
GZe0tQu/vjySobxEBqLwAVh0QWjjtyw6o8T4F0AQMdVeNYbWEI3ascN/nMau
wjclI7fOkOWeQzQW62gEfsQFGwXBA7v7WQBZ5GrrGLjDSsbmYOIX6gNaqd83
HZE5kuc9aTRj8WNp06J8sgRCCLIehUBZCMhvjCoKAtemo7sbxO2qcB6brYk8
kH2llFngvuNzDoQnbFjcDUcxfwOxtR/K9L0IRoDXrjFc7BV6v/o7kdDAi5vS
UmeLMepELL+NOZoXFSia1ih2J9K+C/m6K/PR+kKM7/XnGJGQoIaqVYmKhhmn
tXxMt9iEkoRiV5DfKosfmHgLzcyZwPaSbdUaBdLa5mpZlBF4cyyAU3DxIE6Y
3D4Ee9Om+C4XAfzro/dKVH2QgZ5WNk/jagaioYAPE+N9n9FQUXKBQKbGdsa+
FHBGmu9amaHN2f8peS+dlMICmuSWn7rMT5pFpFI4tSCR/Njxq22mNZ2AMjA2
T7epasLFU5R4d6tlab6l6PPx+qUy8qokyHbTVC7KSdKjOBBG+csR6EXemwpE
GxOIVGfF5XWdiOjqiPFbc+ta/bpYpgnSD53yHMTiVK2V8QKBRF8KPbVEgK9R
zO7svYVlY6NaYBMVRjeJogRPab2TQTmCwlEqUwUfiLSMvaHCpChT2CNGIGpo
iCG4JkX6gEbMt3ueX4dpJoHMn1guWQV6yu7vPacRA9LNegdhsQT2DPCbN1hj
qtUWvcMZD0rM+bo3dShvmDODmXzT6h4DntisS0WyULyG+M8iVvkr5q8cNiCp
WyUd1mkadI0k+i+Wgjljlw2/8xez4RbFVKjly72Iqat4EvuNnFyOT5fQK5FE
dSzxJkX4GfjUo8bX3pJHwwfE3cM0gCrBZURC97zyqPh8CpKEOqlaR3w51EjC
rMYHeUTTm6yESBC91jQpF9YKBkzlAcAADpQxrhmkV1GiS2AW7V7ykcJXRQtA
YXck7cTLYEFoNBTanp65/F7Xql8M0iFfGY+QSV6WhoxIiW64NwvyfEWYfDDk
OolhNhUFhNT//wGK4ki+kIrHD3tCxXRT+DfzjqtvfkmCfxKLirGgQlv//Dmv
zHPIibth/9Q9OedYriE2RqBKj3Uzakx3fSyOE5h/vVV9FK1UNpSN22rU4El+
uLd95vapXwpwl4nlTiyYl+JDgOmmKIBDcbJvoNeVvWoLen7qssZu4OaHnGVS
t9oZUC3ocX6N0zL/OKK7f089roFPQWfHwoWwcAdRBaMHa5m71HXTrLzfC3+v
L5bDKEmzbGpT67JOtOzmjQEXcrOd1xiHdieNZKBGMDkAEKFJwlfvWqwAKzUx
IfqFxwm7DypAH5tfhcIOOFKbEV9caDv+OCOf/XzR3vzAwP/ZjQDXqY8kl4Md
W9NUXdaNGpOnwWtSyvpZ/QkuOMr8CoB/lteTPT6znHJLGgwZet2ELsrhz5+S
b94HNDz73GUvLHVua3w8XsbpAdU3UjMlb1QhyeQJTxnUuCUquy2moqfUGsdJ
hSsq/JtphFlqmL77PRZ/spWFl6xc6jU0WxZyAzI68LRmXjV1tuCBDOLRzXNg
OBoCHMOL0sYeifbLCL2FAsmFiT2MeU+KEISxR2cJzXfyo0SvWma/7SJd8sz4
Wz2LpSq8mbEs25u3Tl9p7S7bBPP3nXqH5S9r75/dPNWx68z9qKEN76593ZKD
SaGL02xv2d9qEs742W1qgoBa0oTno/gjNVt1ImAXhwpArvid6kkv3tiMSYV6
CMlEkct1iJFUHaGyapV6+1blTKMeJaCV/yM3j1Ylo8zC2yPEQ1DxBz64hBD+
2LLi3kGKSm+cwZplO/BQXYLS/yhR8DNYnR/50is3uxjKQnOYnGO0u+d6u0yj
mcqke6jj/kw+ahKWPfXU/gXddKs5QzeqkR9ButmLJJGWm6Q4w2Pqa+7DOCVw
ChFRWQwEVn6rCXebYo152Org+SldCnRVPrW36Ei7hLxAFIxoSuuK3SXCpIS9
ioQNssM1uVJJfTeMEhzN1zBBhMBeOzkSvJy2lsRwyKe+ca8ThCqteWega3f/
hc4s4I73Yy7O0Jcf9NoueN97kBKXGHVMfMFCiumvumn1qMn6fM+ijS0tDpmn
OlmOlUgqiw5LZ4wbXuJ7B/771pllEZjXCVpk9s4oAvQ3YjkExl+w7LR/u0zg
7E9iJ3AdWl4GSFqppDJfqBDAcJPTXcb3HQmWPw2jc8RzPoqOMc6LDCDEClHR
S6RXBzQOWeJ1PsrPGZtLb2e1z4ZXzUxGHFNadg88sGD3a/PkSS5J8siG8S7p
1ZzJx7RpIQP5pKTykg4MBPjB2Depz9rlsdf5Atmz4069o2rjAUpPEGUHlNot
HjNfYAVn1w0kHUt6IDwgnUVts7jRwPMlIlJelRbHW3HKJT85m9bgm9OxTZ7v
COz8v6yskXPsog0w9PlLy0WjrDGvrb1UBbdntw5KSlRCh5HUS7nd4Gnyiv4H
Hbdp6D2aDiME7cSFBum/PfzD7YFRfwLN0JqRifcRFUAiZKGTjVeUugq1BCYF
IfIme2gk3b2d1vw+yBRNzISqKcP97oRJcb8l0mNdrrEYIWY0U8+UZARvJjkt
ZTKk8uX+S6UPN9ylLqOAgq6/Q7DvGV9WYZtOcG1V+pYphYJoMMTyXxhER9OF
C3hAQ3KXjiPsJFx7oAo8gOrThtRUOKldyqd0lgXLybgoY2xDXbZWII3d6e6R
xeWu79T4A9Z0XGwaiWX+1Qwb+Ij7bXlYDsX2frMadz9zfDFiINTPxDV4apP/
mt+j5tq3NSQIQViSMTxvCEWdXrtlqcQ0sv0I9CTCIFocgirZV3AIDLRDOIl1
teMfHEf6a7pwmjugUmlBe9S7qtJJUk+FO0Hl/cvtx4qsVOCIdPGmuL29tdTg
Fv1vG+k7cP+idEUcwC9PNA+9uf49uJTMFNbdRvHTrtZwL14dE27DJPPTb6Hr
aUQItYsNqq0WWUFkvzqnhEhOv69KiZrFVbYBM+CzYFrSDvXy8s/UE82XFZWB
muMkycNNGJOrvuvtB5IU2CaJ8AEF9ZXIUGICJJ1wwc0yp8bzk+H+0l7UNSlZ
avraBdVtiud6ggDXhdnwpeJWO8FNWXby4JKKPZnu5rDKuJ02o/mBM81NXnZF
9ewdOiYPEGi1bN9tlFr9wXwfKQcgQGwmPyQobRuW+cPkH138Hvprp2O7tJva
e2iCySZf9nmBmV034+DyPAnZHqCPMb+CQAd9u2Dm8yNjawBzRb3bzqmLFPmY
7P3VFw8jNkYfaa+iNciZvgRGM32ZyWbFB2Q/9aBZ4hQUg7FM0+DvoroyRokn
pxOiAURGUZZTox5ZmAlQskkVqmr978ju6GltgFUmXNFs+RKyYkEm/IhvAEVY
CGOx0Gv6rvw1/3BS3T5Bhcn3ud+JzHH80ERGIOAd2snBeI2R2NhztK+UscaJ
s3bfXtoCThcSwaXzDFI8kSGmrQS1GRXhws4hI/zAiuHyEZarxTeuL5h6eeaF
p2+DOlx/nqqS7wocd6yrSHCwpCjwc9pF1gMW0OWdMn44Ua7JwbTSe0t2cbaw
mtuSqMYMfZf+nG9YyJhF2cBu8U5h7ns56jgkxQEzI0nww/Dmw/6OCV0iBHrO
mg21uPDOB+pGhs76WNCfywOtHN3V0o0kvo3DJ4omTIiXA8HyM2/ZssHdVbcm
K+mpRrnuTpl8iO19z4Yra+fBv1cNfgw0Ia09adj+PY9d53D2AP19eF0A0nIQ
9KQXJf8Xx06axQHA6Nqdd4IwwbwvPrwKsSx2Bczj5SOOuEMcIzUoO1TeCf3I
l35uusXT26SkEm9SGOoL1vj8haiVd28bzzsR+3ODPz5d6XKZmr5pVfgT4EAZ
iuo09Txo3mqH/Y18TcTDP15yVRmBeVGIp1KTTn3+lCDx9WkVvGB2DgHdaeVq
4CnkxgOWy8MLQtcsw6DY/wUhfY+fQAulLdS4ifzI6kuiHoHQWwYZU9Z6lGF6
5gU+GJJd+u1t7OyKuBNnAELM1l0zlI/Skdg+7+BsKDsTkQISrSfqSvfj5y3o
T7nI0iWpNKr5+FKdbaEtKwgKFezVxSBwOgYILgCSGdIR5jrZMJjPWAXjeHn+
rC+hY/3MBJRVF1GvRb8dMjPB+8eLCFtP/x/6SzuzoxgJh2lYo/aTZV7Blrte
+xExFJeuTl93rXHbWOVvU8OUWDYY0SAoq2QM8nJsYpHjIdb8RbLbwQ87fCLQ
1ZKDNDoj6wo9r8TZTNADuttZx+cNHM8WVRX0XnhI6C7DX3p5NRnBipGonSKz
5SJGJbhG4jd2Iau9OHPD7CmsW480SxHnZdzgu4EiMBrOF1KAAKWMd60lwavZ
a0pJn6YvZNQ9Mjl8VkDi09A/kYqd6inEVD+gDx1QXPq/jdhXHofraPPgy0TY
ZIGuiNlTDOK+8uLt0QrbBlRFT+fCnYhPdUw6RdJESm4OtVlImKlU2K58V2nm
IfP70wrZT8Cv2u8LtPPvuq9RBBYTD3g9Cxj1AU98zJI7fsDfAtMTQrP2s2yf
3nEXUto0sRKohC/gDtIcgbmSAKc/fpOOmCyYRqzxKFFFCpQiYNFPcyur6hlz
DHYR68/RP75CfR9SvYO0d7tujtEATazFwQVP1QCRkbDkmj13ZbkWAgmIYLPc
mCOdeAiJZGt46g/i+1btwDynrigumXee42ERkcqhTewWFFk1S1ufb0VlEddL
VMuJjMrmaijp3VuhvqMffA0KGg61ytPp2O4W/ebXYzB5DAGVwNuFYeaERlzY
vSGJAch/CI27naAbnaL1uRYnCd6alDn8oZVL8gGpTHWIo06/e1Du0CLS86sZ
0fmx7QSQ5EIlrCDt5q/thj3nn+maAGDfA2EKSOZb/gG/01Ub2QkvO6ZmAyY9
CdvOGHQ/FpWYD15OgY8a4e5NJVEPsC5SR5N7y38vbkrXg0rnExNs0HVMX9Dc
+FjvzL+XXkuGuTD7HwIvrfTYAX+oQ+2Zj/RS9O94RlCe6Q2SDJWUFo4nCXNi
/O0tHunHnKTtwfkBW0g15Igpt/3ASITzNjkHnaTD58kiBHzx344IA/UtFpb1
4Ma1Z03r9wDUhNTIg2orjqaSNVlmSi9fpCPVm6vg0YiAI6CopdP621wO0Dif
A4Ve4hkMgrFjZ1lNh3bc1TPHzDFZVtfzhnGPlUQaN5K4qY9hgGis8sZsikvb
UnzKFT4uUHjANvqhX1ACYZxf6McpTosUVigp3HytpnyHwjsTXkFRy5Sn90hb
jh/4l8h1EavnmaxA83RSDWvTB2gAw5+qQ0rvnGuzpOKU45xdOHJ9oUTqWoGF
/GuPQp6hugfDr1c0OjXoYbiQf9smOhAATbbDu3WdFh5ALu/jBkM0lkYwEQY4
x0kKNVvEigjWY5Nq5vkfEbTZOPUt93Y3N3pt5Ow7RBsdL/jR43Thk3TbKTOM
gBXw5rJMeE2lagk7CYF+s0FGX85JKlEXJhwFPHtSTQGhPEVK7prKuUOJCEkM
l659IDci959VnSX+t5Jmn99mKTVsD4G3gaYEOTDzypMni7SgDO2ntt7Wcs4+
zwJa3gEnka7hLHBz/urNs4uUBTNnjYA3hln9e0xQik84/JLRmcoov53okZcm
k4UghrTzjbjabq3+qfJ/RCVlkPZVSpoEhx0ppUrPL8BsGtFJI2wLU9CHx8fn
oqs1hAirz68WFZXdWYT/KG3CAXandW29mGD7JZ0bpXYQ0syH4QZacSyj1U/O
LZhSxUgyGdtCx+HmNYlRE1PI1r/curMTsp98QOQBa+1IIFETPmJiBFuejmPc
cQ3+h/x/wwB+vUzSYOzs/tWhido9khB2XqKkP3OmcagDB1FwKibbeVKSo/nB
HZ6iue+G3796/aYXR51id+We7ZCW2isq7YduysWIjS4hF2E7mBb/fzQD+pis
QMhiZXnCbfN+fojuynLwMvFUNfPaXeJvVSMdE4uIosimk4pXB+OE65ZYcqwG
GmLHq0rhMEz6CKan8EwPwmbGzAPnzT9ipYJKfxw4RCd3K9YFKyo3XL39Fv9j
QD59lOx6X7zMUnmQqnBP8bGpbemFX0FvFgkJy6PdveyI39cwEd4ULKiO6Mim
lP4BQmBVMAm/1yQGjzoLSAaTtywN00PWuIX03EWd9C9nqdzohForHcOl+Uw0
tA7w1xRONmfsh1i+ETLixIJ4Y7W2NdP5NiO3OZ+2MRXbBLnlup/WAJxqPFxa
Q0tGsglE6fFV3KcZu5cach/pmbtnZjZiy+C1rrIiiIe/hHgnYeQxHOGlU1wM
ses7X0wIW+sRUnl10v7zg6r5np0HYdFGRhKkNx6O/DlcRRKYZz+FP5gk7ktC
/ECJ1dNn5BMjIo1DMx+A1xjmM12bjXONmJQHRd/mAY2DykUobm4eXjSZ5GTH
lCay9bezr4S1w0IYdQg2PSONgf4RhkaQIKjXMUztUJPNeJ+jaGGjx48/ugoR
a561qB9PCwUnbL1aSagc6feh+gye9FWiMyRSEO2WN2DCLeo6313XPSg+oTLF
wNwIn0ut0ARj1ElJD3hZ8nXgtYOaaGvKwUG//uwW+JuYbPa8GoqW0rXc6nAK
RssuRG5G0+q0GXhluCEtcg5PErsJKdFLdZ883BCqCpcg2PQfdAXO/gI/t4Xm
QlDh/ScQfyPWyTASIrDFFHtLYs8iIiDAQQUA46WAJqkn7vlrh3FtIcb9xdb6
NB8DY74H/rcKKuSsRafLzrKIXufUECxE8AuUTj8sQGnn+l00AniLhe8cvyQr
cZDWYCEzGZzKKffn+vUHiLP6S7Q/wE7kWq+eI7DDi/snwou3i2r02zjKbu/f
2bn7CODB7N5jbjynFt6E9WqZNg2QH4sq+lW27vzVjB35P5KyBjeXgnelNN/K
3yLFr8xp5mi9qbyxz9E6a+SddHOmSufqBnaWbPkFtzjeu6js6Hs0SLZw6j4l
9i31Mg9wn1mpYMv2sQdtphypWsfvwKaYREFrWpn2AxG2/HSmNT46bW8NQdVd
p0n/zCTjTn4hfW+mSuFL1DbBYTYLKPN0oentTRh8EfH2euR+YzwD4Gxelm8N
Z+nS/abeVDDtzHDcFSu653Tbb9KRXSs2BhiC5mbie3mWbl9w7BTF5VeSUR1C
Xx7WbIEMKIN6TzdVyX8xYgfvQc4+Nap2io8KdUwHYgFIgdsOx7oO4mChvibh
v1AG732byeT88WcD7YsNoL7WQW9qUvJFH3jMbRDv4fZd3+VllKR8V974XkyR
8Hx4aV1I/uXg06PMw0Yo5U0z+SaBtJZ4nWPHp0uFiANvUT+rj7Cis9UC1a16
AGvEokhDDFL5Q0YO9bR8+0bV6xrYScfYVzkBd0TymjpdojK5rzWwVLNSjE+E
pRmg68DZ+SOWllNH6rsUfpHLF18OIppoTllW02BOX/5n6jj32QW5whtdF7BP
+H7Ww7tUM922RRs8dQapFWtvC3RpC5Sr1EevrqJK7KWsJzAs7Qrkk8z14WFb
prEMSxK7o3e9Qj/1izVz9RLVmpqEK30g8e1QERjiN/AMQIHxa1oe0wocvEQp
OO+UOOvnmvsMRr+fGZ276AJ8g8XCtDC/pLLWOWPxNhjVNdgMRNW11lAs6uOH
Z1IVwgDjpgm4OVTB53K+2DqO/qTtWLlcPR7RwSDJdPJ4IWVYSeuY8jeXA1tW
KAqENI/36Uf+YC6xummiW2Y8DuK2kqSRedyqLeEF3LIvVe5MFwcvhbJErh+R
bL1MuAVmIkFt0TOkfQtkOxQg3qslsVxa5G3v2Cqer3f5D3p75BPhBz0IYKn5
O9WWLWPwwlkpn8lpZ4vvmL87QEYmW4yynZzylXjrQcsbbHN4++J3JgMOl+G6
O4d19sqv52Pam/BSLWHSoxju7qO27rDMThnoWiIApPNE8qSmNIfzcbIE/2d0
8maJmoeW680GDHm33HrDx39YEcJKPaEXm7kjnRRKrjsI22D5dkWJbioJCV9S
+6tih+TRMtgVijtqDXMRaYvfNTfBAuxzvIp8o2DijP8ZT+06fVjQ/YoVr6AF
f8eCT6n7IGxdYwULfm23NOMpzQBFIkRjU7ceKFgzP8UtTmfy7NLbwGNiajou
uuC80ocykV4hjOLAZpZJL93hdMQEF0GIBFBXAh66Cr9mYed3NNXdrlbBVNMN
U0iBPP67TslcV6jQOGBK0PZzCjR/cgQDOw8zK3g+cPlLGLt3KCLfQ9jBjOt1
umWpwt2hF7JWXEeonHKjsPlyodnmpSGIx336YM0R8iHZDYLv6KrlQ5mUcMnG
o6bJJfdJA1cPfmCOFNAIAzJR9P05jY02Rx1GLFRSABAGrckrnbQ/Z82nwUIS
L94spNobLPMkfoc0mv9tDBWtsNxXUBgaEkr2SRLsJitWobExmCLNxceKqWXS
/493rIeotpUuEtMGOLdzwG520TXgNJXv/VZOXd9wQ2wG568ycEr5EbErw/Jx
NgeUjrYPi8BMQdJIOHo8QKqyqA9Z1PJU2a+FlgRYmRXgStc5o9fAEJ8Orplf
Dv4eDfOb+6JBNxtXf1rgVMrjoct9zh4IftGLdaQivhCcjQfYO7pqSR3KHef9
RC0UpTh5REJ6DtG2RRwcic3woOdEIZhME8bQgUO5gNRhULcl0mIppdm+eXVn
sUqkG6bHmO7kNfjjBwoYYNo4BoflXu9Tjn7j2bdMQOrrI9psbhtpqR55TNas
jdd1+jl2shP+suGeonxzfhAJysJSKyJadueud+1NhLyFO5MyGNRrZ+074s0I
/4DVQM1b96k7BjPUb1usfLTKx3E2ZGpfweWM5/DeW9tpTczAX2v3kdPUKqXr
FRdVVSsJnO94fCDmKQgsfIFP8Wm1lAk2UbglczXJcFi/muflUU8SOcahI/v4
AQaaufW7cnoCnQDQPfGAPmYYgG1ldZut/B8axTP4+NYwHzNOI3amSvfQ5i8c
WroDO+6g3sQto9+Uyi4yMeVcNJmcTwWa5zZ3FNH0aH5DeHf8geRGKV6RpDN0
ZcdMDVvfVQQ/BfmLB2AxfvQTH97NMQSsFdvKAR8cadsEwfRX5TrUefI1zdVa
kjhiXDFqw8LN33VjGVQJQvIn0MH63Q6ZuflPPB++J3+AsR5uR+KDiF46OQ5M
ljIehpVVRDXwpaEtroM1D8S0wnJQhFHSpBS3XSmDbJKVgvNCAiXj0iMa+Ome
lcvtFTo2JmtogeJoIA4cdSkw2Og/oqrRtP1yb8Qip8CQqCl9PANwDrFYhGtm
pc13THQcE8UcB1CPlWyyNPLs7qaHX0PLGdmD1IMV6oylodT56wa1JC96ne6N
BxnaN+17lpVHZ2z+TE+NUyyyZzynV72mcKKojyTJSKfzRt7Jqf8cHgyXjbs8
ec14Y3rfQbulMZgecK6EYCwvMB/Pj14ip2QClYzLqdBv70R9kkqemYs0vx3j
WHzqcNY9i2ciPaQaqvhvtHm+4iODwfpHcnX7n0yF+c1+fUxRSVHiistq/8/e
OxnwESk8K/OuUgos3QmCNvdjojC48IEIsEK3ZL+b+cUbi7uwLESa7Ph7xuXM
zM1GthM/pNznSFPUcZ3Ur0omj9b/q3uBlKw2HqoySs/79QldyR8YftwRSkU3
aRlY4Qn9lmTnhUP5V+wrs6U8K2q2lNGo3VyzE6cNtBb0Z0sXHGmC8mufQSIY
NEZASTakMlc17jV0uDC6fdC3d0uxgmu0SM9KMjS/qek3UOMCSj/R8AjV8cVF
c7FumGNfoof0ya89uVHe/ZhFGbYH3vjSe8ObyQMjvAVyZi051F8DQio8dbAv
ucrC09itQiMRcZEB+z0h2W4oY9U899oM66mj4dGRJDqH2pWmx11bLsLmk3pJ
f6O6ltvr/TC9HvetRTwpsVyt5c8jZasjGv+41y9Fk1Ao2mQd1Ksk4VidT2mu
CATu8B2P9k3G6AurGd369OfqeeCQP7MbRsvZRbusCQDNnt/ywr5OnvwSHBFI
zYdbwB1uu+W2Q5fJ7NI4Mbfb4UiDmGJ7G8VCimlqKFNEvHuf+mmAtHmRPdPe
97pRODzR+A91h6vZdUipMAq3DqdK1xGAeJqWSBaXwgifn22AxItGksDJcijW
YfdfNsda/NFQoGrsN6poeP68DmnDmcTgtMbiPJAhrHDpi48Vf9Ps1CiIFdlF
pll1AiZ5UT5l/GVnhsDuqiZaoEJgXB+pLG9j22Wj+hZCdeWeujmJeyueRoNx
mT63YNafBOZwtTvQmG0ReNkWSW1l174Sgm3NupAZclO//V4v6+E6zoW0sGOL
/ddQlfbiVl/iGzk9b+5CZU077oVzybxhB1nPvocMhMXoR8x2CdQrosS4SmIL
Bye8njBJIt5PsDqzFwxsVqZkzx++D+/8aNZtnvsUEtUrRNTY9FAZCN7WfOgO
8Yi8HSIDs5ZvqZ92P1gEU1SpOvpixll8YcdDTxV7sSmHZMDZHBnC264TitTu
e5lwMG73KEBH1RqNYYp18gLu5GgN1TOAN/+FruUEfAc60KkdhQ4rnjIYf1Oh
6DlYyb6IwBGHtCXHQr3lXyX+s/WZ5iAglw8uvqbV34iB0YuFn/fVb8RxkIm5
QUa9vo1JdvU92L4FUBSbpL5VtYr7FLcBhxhX+xMw9H5iATG4iR10h44oPiaO
Yf0QiB6dDrmWpIbsqqrKOMf1OgR1O7W1zo+8keQhOuDxvRP+MH2Lf3nnybnV
tH11f0JLZbOPOpLOAr9A/zNy0s7chYpPTIF3Iua37SERS0EJEheiLT1khxkT
GZN57/fa3jt7xoNERpNN6KKdR+VuDkmkdibWwsLIY+UcB8jzXdvElss2iGXI
NqORvamBFJVZ12gv7JlWEDWqzIV+XUmHGpT4yonMM28lyEAvKlrraJ212yGk
f8iTCd7wET//SAqjcLh0aKPZedw4CQOCFPZWbV96ML8/JQ+YqfasNwIbbPoO
Mmvh0XGbSXb76uLDFOuCs6odRbmMz/xQJg0dLSbUF2unAc74WvRyQJjlE2o1
+nHku36hTEmZoNcxuR2QJo+EcPo5QsXUF/abGgSfKng9TsLxUPjKbyinhqYi
1a94qkPlY1+YldgqIwmyTH+NN37RLYC4oh7LDrmQdrBeqVq3WBPMrdtVyTRz
HdwMz0osqcXu7ZYTMKs0Y9Yc6uv763MlAIIhogVmFbqoZYTwKXz0maeHfodg
0ZO1FZy6QKmEMs/DoTkx1cANVlzNxBE0/kt3TFfnkXcK9UmPqkgvPbrPMKK6
fmEYM0E4DRTJZlLyqfFsfZ1JWWfOo+sGNX2+DiDjafxYYw09sV0CcWRluQGE
5C8eU/sDVKCdNQl8uq+99Zu+K48jqdgDYXbcSE7pD224thsP7SoQnbrHoptu
/COOc7FJ0vDZkgIYXOCodWcLTawEKc4tyRhCYQH2GAbYhZDXSqSQRLyfy1z/
o11c0whueFjylYtp+KlkoYERz7KAFd9UtyJ6pDgs5RzsVhR8yBd9Giqgy9ZA
eHQbYCJASvd18VnfQvyoWzOVSqCfBw6ueSVexMBrGu/56RwE2NGdxa7Rc/zi
ADZnPm2D5rdNBJ+hmPG3DO2c9Z2kyWR4E1FXt3m1TrH11OK+HeCBbHZSs2D7
NBloW4LzLPnewosEHItFBxJN7Ke7FG2rY8GK6e9Ua0Cudm5HvsdkGFtmXEmB
2WGYZxtaV4j65f5ox8JIjj/Kej0Sn29oNyS8DpSoou3ksmVd6TC4+CEzmyc/
bc+UUDTpGbn4PEuOpKiaeg0Il2rFmRWVPIym4Yzr/iO+MeYSKoBEr96u1k+m
p5y40baF4lZpZv6NpJrb6/7oPO5uOWRVHzXfnIZYH/pJp/T6859IdRMoxxv9
yQsxCu9t6HygFVvYJUruPzz6tnyNmCfFCEPrjiRCVZm/+HYFV7r+ARVO3yqF
npEa6oJdxX6BJp2JMjUSUO3ruMtGUnAqUwcNGYnuBpFoYhAFvxfXHBHqqVS1
Z4X4FjdyQR2G1e2Z2H/ur2N9VNi1v2Arr8xeQ9u9WorXuyRK4DjMgeFPZfLq
KmdU2aq9vzomvqvGvGCy6KXnsx0U6pmDguf2tANM8SnHUNxTgSxGqgpCdsZ7
+FFcF2zf7WYK7LEV4/MbK/cNGFisWPIZTQKzf/+SLYNmOt9PlRE064GYxBRK
pXJRwZ+pQo3XkYhK59Lw+cZpWd9mGG9J9yBH6YJnQnIwMog2VL53PfEHZahJ
sUQL371hy7/OnAGawxFddTRk2rFitBaT8JuuhrN9WS5lZrNr8WXThVvbH2FF
GPgicmRT9JuLBME/4LbYNEWoW3vJLmVeYxXIxZfmqyh7oBlhIMl53v2wKlqi
w9v6mn90aefjHnpA0H61p5De2MdC4O1GwN/hSZu8uuv9nKzpfBIvU16YjEpA
1e+A4PEjmPXBjwxtDjeJUEmKeOe1TePHWbiF5lS116OLFfWZnqc3E1GUtu3N
oljkW0lK6WEInNIuT13CXlKao1ofDmLtzzsjMUy+SBSSudtt4sE7NuSbaRAV
jJ9cAxn7aGFZ7m3w6/6YA3MSLvFuqRS+P+xS++pzO5IyashebMlk3Ubjiqex
Slx4IU9kCpVL81Ic82p/IZXHbs+KRs3/gJA/vV2IxaLRCn53AirgK96VnP95
DKdQrjwu3PycVfrGnT6AJupjNSW2zXukjhf2maZ/5TqoX3IQb9FJob89zrsP
suGOUUekO9LdEYmMVZh+jhuHl/RQhAGihgnOEBwdkUwoni8G871PJSst1/Pm
veCZnp/NtkzPSGcGIWFw2FV35tls+11UcGwePC/phfAeb24Z2oMYap9fmXbE
p0eVrvPkkz2+pnX/rjcWNEnh6Ms6nyj4B5aQ7POXDb3a1eEnQxxv7LiYqAy6
QpZvX+r01L0oIoz3whvG0N7XI7GAwGCONx6D1MAk4jrmAxSRSLOGJlRO45wN
qk91LWw0TJTUEVplAKSSW/oSARoHfEc3QP/yqeAHqc1eWBM4PwhpWSd8DHGE
T2uXR5y9d0+CVCepzCSDkCmgrp8P0Mu0TDDQem1KToF4GxJercf5fAOnpW5C
8S2F0DQeRF3eCKp9Ivq+dJsQGlQCfkSgh3b+bqAi2+F3awIw9k7ikrQIFkah
kWVCZxRhXzONwEUtY2ZPBH0Vw+8OQgbayqeU2M1fpmPyxR7/oiak9puy02NU
A4JVq/4a4hjdiiu/LgxEEbX2wSNqoReRriMbqbrAm2TlHvM/i9H/Bb02tQfl
YYd8zkq7oYRBUVehH930h+HcCE1vxFOhyk9G/1MWLWsfiKjK9mGvDLQ+DAEu
2QfWx6sNa3wq1i4oFBH0FGSBuWRJQNcpLqG5zM09Wz+Okc9VpKYIBZ9B7Mm4
P2lL0BEvapvDl+3NSKEIqauiIfkVvTyNRwCIp09xr5xzz9bpgcwv4Mn9fdGs
xgGve2tUvItacUsmry0MGFSZqnuad7aXC/SQ97Tnmxv4k9NTHaE74oFcrUjZ
RZ68baDR3RxKZBFgwa8kugy/9w4bSTyAH5aB+jkeBzXgjshVeaHj7Two3You
HSCyLUC0Zed6oAB/7AdxfD8f7QSqsQAGaRE6pHUNMP9rHlUr/JIFvscD9EDg
qU+Z9CCB5PRfmWCwzq5Ss6nPv0gGiQSkL6CmVzNJjqEz5HylSM/Xn3e0PfQG
nG6n7zCwiuO3k5VU/UuU8VtPvfXrwJZLzGHZj+twb9P3q5xqyZiat26ryFkI
SayPVyPoKH4418G3T53F4TV2XfC7qBvhfB95HaF6MYm/Qzp9E+P7vYqb3afe
rkAk/ybftjYcYV6MV03iRHrrqZYe6obSot34shgeSpSekJuiIo4qULjUPDzq
L1uEtWSxFTt6PxzTQcjVeRcKFSuXC5rtcf4I0UBJPX5HDEmoQpAqywtpptc1
lUUZhL8V4QDQ0R97Ay6OL4mS7F/S11dUbn3oJiUCuN/kompfzYU/t5ATjNFS
vR6zi/JPbNK147E7X3MOScqcHMnK1YNY8IuaUr5PulASxqqkYRnYNy8lzs3w
aOi6jLxnFZd2Gy00zv768alkmzC1KCpIDFuDW7fIcCr10/5h9iQ18ioZ+zWv
VMSC5RQaXPb0fHwV8WSRv+lTg4awt1KJmW73UDB5ZJU8bZSJ10PVM8YSeOhX
GsCh/tlNKdLf3J605LAPmW9/gSr5cT4t9uK+FSoF4R6kOuzEhaonxllkbSLP
+CQRHHK0pEnf1ZjQr7weQsZvWVyNy0nZfkJDChzC372LuLPh/5o6vB9Edg42
lN+LAIPtiY1FZV6r1WiAxGqZOuYzqZjg1kXorTYQfcZy0PBn0EJLm+iYKFtk
o3M8ruqLpu51KjDmX6cPmxuE/rQI9/jZPQcZ2ZeTkl12PEubtiQH1W6HrtnA
0QzzBaiTplx+oewaY8qZBKCpqDnST/uFydF8pU3xM811HC9vLlRYGIF1Nb+E
IqE/3le/agP89b5TRCHPZoFNukUbQJvz7QxQYKXRKf7wVPiKVuIGct8uKDe9
oJIb2vfomsQgX8dhR4t0nTBVM62U1xg0B0gmxJb6PTxV4dGeVmW6j70gzJFg
IznUwJNDTU9OsYVcutC8Tk8rLCONap7mUWhzPiTGqovzgn1OmJIzF07Kttju
PPlLfx0F0vEdlKQliob89iTnrj4EWN8iyoY4Ne9ARUli0V3K9lPZm51XmPt7
/R5d52BsJkUVti2oT7cSeVMbx/dVfEuz7SBKCu1h5ozfiMbBUyGFZZ0IBrKo
+AxLLmyvHDp/MXPULogILzJZHTxqpqCzmcXemY5+R3Yz+BO8srh9UB1Uypjy
T1f5pPEQKzzIDZMym1wBrLORwsAxJN3TYQUxNXqpUCimCJXzeYFXgqrvPfnH
8FY1qd0G8D6PyxkjR6Qe4mRI4wLeKO+e7Rih1j9fP3oV7lJII64il8QIdac2
66f6rN2tB0uITvmYKFs8OqVEIaKwBvbEjIWk7b2qW+B0oTemjheEcLfixmRD
ODG2vgea2U62fgCEY5ApRkW6IOudci39SkD9GwRfUllM4kyId0jrd3zK/+UZ
gsKKvksfjK+h7VVO45Wtf7ZlKLsaGIiBW7aeqcoS2vRr+BznuHyBTdslDTuN
Mh2nSiQxnJNm6pZtvzQXdyVS2LeIR39DY4vmLtCngqsykgUw5NQCL4lZ90r2
QSsowGXOXB2hW4xuGFSYDzMZ6DLIyaMtc+W/OLwOdWeFrYRgcw47zXNxtCvl
RBlwvxRf5ckHahFnuZMV5P+Qf1mzv1QWsLYCU45ziNrUFszWl1DjngaDkFJF
zIZoyJWwG5agbyB5f1NrdNWtVfts+LKlaibTr7QMPjc3Ro0qOCvDlRYsKwVj
ug42o6JVVTXT+3q5+W7YqSjxrkBRtbYyCNueQwEnfebJw7eurfNUNd/WiXjc
DzREL7CWphrsupYzJxNLaV3zH9pk2kXITGfkyD+xCDdqvEH2nq134OrTXFPu
QlMM2qY/YtBJgYs1idyz9FMRTWzlP7oipR/oZ8IpRTvIrsGJ550xoBkEoopj
bOL3F2s4f0cy3c/r8v4uonjbSplrMuJj7pRexRZDlbdnswfLCX4bpxeNiEca
WQCPt2PVFpSnv/ymX6pLO+ah2PgCSlr/IkdCXuBTmt+C99B/rYbFo4uiLx1s
H9K8eJvFrQrmlfIg+HfkGUhe5Q60DQ42QcEh7J1yZ2V6FQvyb/+hh0tcGGGG
ul6LZrhxvezQTSgFDrJvau5CT9HgFeYOQirPWIn8muALh5B4lJK5i1DBGIhi
3NHZt7qf/EfFhc1nKAohqGOp0IHTYDhR7y1G+GkM1FWOzxn3HEhGko5gR6nM
R48h2RodXpStLQpB2Y3Epkmu48INA3hSjRz9fjRFyE1dXKYvPxGUTBit4aSi
Vl+Py7CzxyHHIiZUpoRCBe75x++zk5QzNUL52sk/JChAClgomuJOudxCsH7V
DpzT5j2vYAlvA8CZvHUh9iC+bNXsOpRh1d6VUTVq3Yj0rTDrp/hcaEX+GHtD
UNRtHalsd1SOR27QPKpWbM2+HULvMfj4T0LLhSwT/FrKFHhz1L+nHlJ34Ci8
Pq4ydAZMiBwItQ8M7pTIERjuwW3eTazujHkLcorXFvFyVsrGKPNiTScBdukK
+Ooan8mrzqWFY0koS3cAEKcOC3NhUMwjmuV/gglteQdsIhhB//6EFoOk2Gtu
RJOUEozq+b6R40GRNq0KReuFm5CtYjN2f1Y6ma/jAhAczUlqs+3L9QwETjVJ
Jb80QXkkv0uaALWj0179UTfzkPfd83eyVjysOTu/b1PCNqrF3fdjn/YWLZqM
7v9RJDwZGOguGIanbxe++MLKq5j1MCyccpLqISnjIoBrjLE6W6QkKVteYQve
1nKQFBk2cmX7oeWzB9r66fXepEcW5uo4y7K93jvwqZkx8UpQeMXI/tkrZGFb
GngLxi8wlF6sbX2VwyBl9ZWXGbo3zIKtBjCkH+gIt6yUcSzVy1AJ8vvqwjmO
SnNc463YIwZNFu7t2AFYh/jOWnW4hD+9jU4CyLs/Jr0PbYqqS9OWYYID0nIo
KjxiVpHpmjD1qFaaI17wK1jgN0bZXOp9uT+19PkOVmRjJ7Rns2fMuNVMN860
48LUT1CqXlXXEVBqKeHSp/t/obkdi0SfuYZegK2EOmjAqbv91NCmPW8ON5eh
XCeH18tUxfkL8qkxB5wKoY69fyeCwGBMfEE+F9v5l8qizSVlvYySjwDojpFA
GZ5Ojms7xS0SC4RInmV514abIE/mZY7L73AEcoIrmq7LAoWQhVZ2GYJtW+11
8l8RMD8wGmB+gCT4Dkh/P5qshZ8vusKvkQtJrR5Ejaz9oMd/z2q0ZIOPjwUJ
cV3DiMcj2W65n+wABI6mHwLqeM4WGGB22/dOaEo2NELDTfWYAjsgnt2lOrGY
DuFlBFp/K/e48kItnZwLYbs/BV2AnvxPniTYkusB+S4cN+lqhVniYvUbaD4V
9mDjU5XP/G1PXxHAKWajoFp6XXvhcUHF6daRnMVfvlw+Px7c65LqVLiBvcvx
zX4NCHsGHvsFCpbOEM3ChC5W8NvUKmmiQ2Fwd3dT1sgDg6y+OYkGPhIMpfK5
yPIz8n+sOvh08fxVGEc6PmnlHYvywaWSs5pTQM4kdr5+OmmaB1D+Pv/3853Q
d9gwJuDMEOGPK/sllUcjYl5du4XYKyNFjZ7TNMQ3qKXMvQdy5nL3o4LmCDik
uD0ULq8qWM2Ud/fdYJ6u9jNrNAp2i+jln1ym9V7Ikb4nTYHPvF9+hY8spcBF
DRPpOXBEQLOC9EwLRoc5J31qbDA7jHmCpyROiCl8lruC0+MsiSg3mjMh7Ohw
cTZw6XHW/Zy4FGF+uMRzfUfuRsUQ/IgC+W5Ig9q60GjfYKr21uniLRcKcZvA
Yo5issmFed0N8ju3lM/1K+9NpxWmI8ERpWYGsU49pe85mWV7Dt6FESQCvcfx
/ahPbfJRd9ozgraucayMgCKtCzPoD3+OSikylYvj77evk/ek3BXzO4CD1s33
mYrrINDCXnsQkZ6hI2tQ8mUQsJ+IXXRjgdN8QNJS8eqjksAheiTjEbrqzYWp
LSd6iUvD7ZHPONZRwe0GXjSiPLFTw5rOLTzFtkJTAyTmXmqkMdlarDOUIW+v
NaWFS6cU24aBsdqA+CqxcyHlee78Ty/wZEH5Q5yP5lOpO/O3tBKZRsfCsLHo
AlLdtgiLyOVMbnc8W0xsnqPHmJ4qBe8LhEC9LEW3BToNnnKXYAigCS/wKGxU
8qsQjqm/VCOPo3aPDozNsAC3lgoV/bAnqssvgvJZHwuaTa8Vxt+ecSiEXTQu
XBzJ3v5/NJw512816GQBJfnmSqWCvel0RFe+27XwERWEl78sOVe0WCqiLZS6
YeYNUxPKcOZwQ3KFMkDQ8NJRr4C18hdBaVHQIyjRl2qJMDvH0HxYcM/IdEuj
8Vt8AGffp2A/PxqNot+TwPylt9dmGaRnDTq1/wuCYbZ+AnWAptQgzxiRkzb1
l1yESjyXp5AAYslvTOV8GQb9RoHVVxkNZGaVhTqyKXonqReFg/r3qx42vjp8
tZhDrSlHwQk4jUvBQM4NB1XhR6diYHWr4Wag5+vof3RnENvbaab/w0MtnA0a
XJDLxRp+9DZoDR+K6OCkqx52AKxdAvXVcWdR9gBxg0IDRPQ21YgGRAGrKfSu
AHEAfAlBQ9MtB7h9CB+06fY821M4j1aeBS/rf7ixoyUF1RSd7BvU2Ax5ph/L
sO9HqiP1aiGXBAtbKbu2u2TzAGYM66Nq2a9tsgRLaKBFx7OmJjFIciNWtjxr
Gyr/h7c87nblnlBCNG8Hcx3R8TEKpY4UmtOiwutcWIi7j9AirtX43n6OAGnN
DAOyV4WDPKIuXEngICVDy157Q2RR1pxsR+1qmOZ+qMn+KNiC/KC+BnH5Nmo8
2Uk2pAkZXgXZGl6t1xHFKa2Be/gFZY2pVHR4ex+D+dklQacRPz/PY4XI/mhu
s7n8hv8FX9TZQACFv7p+e2jqFCu9jxDrqNwm2gF67u16eAIDXD6RV9wfMTWq
2QQ2J8xOuNsOeKOMA3CdtAcYdJPJxEZStvr+ndDxG+u7EQ2rimMsyrbmjsyW
8njMfd7BQvx4E7BSya/3Z+aCeiCRe1J8WP4tGZql2/U7f8v6uJTStiImz4ix
Ukaq7ODceJUP+yn47rpLt1qGrZNlN3bYS2a566u+2UU/hrW0tceeoXfa7eqO
URpzQvoDGqbF3ghUurpjBsDukwzr79PUHL2pyn0N9GtMaFSa/DDki2AUcPII
P0IFF08OgWmadGU9FW53/ooqG5ajff5ke0QjHrzUBE6+Q1z3k6+xlcyKZsqT
0rdIz+D4wa8YoYtdxCpLsqxnyJTco1Y88TtA0G8K0smTFY4eavq04T7YJH/w
rKetm0QI8yurCGt4Ldr43dRctAQ+Fk78KSiwjsU8lC9KY2X28+975JriWxh2
FCcRiCK0FxBk03gYy6OGnh7rDh54ClZYMZ9dIJMieX89DQF4a3X65HVYZfOG
gKYaa8ibJ8Uwo9evLECw4UUyxAaH2BH37MFE6sfyT1qpLrVl3j4xM+CqUIzP
VVsWdiGrCErdmNAVjjRvTtH+gIhcH0D/7D9CrpwjVlt03OMlyvrxF3fACD4C
ZPW8ifdQtpwLvkuD+YbIf77E11tn7J66HOcnWqaV1vUt8/FE7daQCx1pwPop
EDdPuNc9zT903RBkEbLk5HdB5DkuTxp4+PNCp17rXYx66pmi8WiY3eFxmabk
uMBdbr7mcrEFk3sHqa5f2QSUl8B/i1IkEnRdeDLlJX+Mu13Hape7HWd9wNea
/MTHv1VBBuLP5sTgIMSeL2HyvsHRFKgb/ER9ked+KsjxicJfcP1PmRRJCIJJ
DcZyWEuBs3PkETMrrVWcdmtplaaK8ITGTo8CYB2PY7aDUjAfExpvHP1m7vco
IeCV43Ni2oqu5Hv7cKtcQYX0aisgw1HgVJ/jdwKCqYQQ2F8RcMG43OY85Mre
zPSb+8SJjr4KJ9mz8DWyryfrCepvxD05q5Amo1S2d1MNFUopkVTW3O7I6VY2
CSRPdSvYwiFgPfs4AEJIguXJzRFZOXEtyo05hnyGLqxnR9KLqMSe2pTA1sas
ONDXxz63T7F7xojslsRICivU/Phwt+4vn8mjkiZsGPPfIO4Zp6UGpLGxZGMk
53R8r09YJEwyRnKBhcRiWEHkPzYXQPF+jwm9mZXQIuDVKT3zgnbrdmwa3g6a
KDmq3BgR6XoQAffaCN+MWDQE/FzdMSv4hIDbp6I4YmT4rxVYmVx7Hu9Fvxea
doaBGHPbTTLa0E+QdoNZUj8IO+LPZe6xAB2jdn/rjzMnJvdsUSjZUvzqNMgx
5+zaPSBLboANSXS59pqCiGY0Y4yWGtv9LgXsSA02FO+Kfw9HNJr67xhKyd6B
t2vGeDG326ykHMjUwjeZQIGSsD6h8tBkP+S8X7O1EPsPrl/bRi3jHi28CgMC
0KPNkzSUXIxr2zeFvwuTFr7hJq75ptGE9SvRoWDfaQ26vjDQl0SixXBb6X7j
ws/cqGRH+xpWZjILVYEBvhBiAubFFqGqf8U1ykEOFYM70lYB52snYUIVKTWn
6bLg7efCeoynStRshlNTQXGvOnNE+H3CYHqc4kw77EDpyjxyEYoDKyTsqIOx
xfLlydJIH4VI59gSp4fYgHXkSk+EJIbYNaclKtJcMryh0jd01Y8O0NHeGxSJ
UKj/I3jbO7MM8GrCMuCKb/ibhtWT6jstPic6g7vo15g85zesxul5SCzLNEiP
2qzAqIDd7SwxgkqLFaTT2cBOOYBHpIH301JFnrKuGrT+sZsznUPHZ5eiRV++
VQs+l9WYgURlqvJoyo017JBzpOiy4SoLFUQXaP4gJHUrMHSgqvnCUNUhZHwd
0x1E6pgsDgnLvHZIQ3bEuqikiaLYWXRQuB6p26p5lUMNkVniORzaG9iizA9D
cldEWhhS27MV3d3HY93IoPVS9UEFalpdkgOsBYbxnOdL6vS5a9KD53YPMdTJ
OMsnSWctLjCT8wa9sXOK6FNPaCFHKFxhD85B3ILvuxR8p2MLFN00gNc2eGZk
2XobmxWPV9VtPNsuTrPKwNShb9/h8BSsQ4ryvQsvFFq6mt6khBSDPWiV0sg7
5Thp6zQOqQ+FDUYPMpgcAXpZkJ77hlKb/Q+cvwOJm3DOdLCekvkNE77rLXw/
x4g7sawvZaShY/DA9d//kqzJdOb0r9sBhjKpDqs5C1V+oQvl8qSJgw+CiPhB
V1104MkTeEgFGdYoq1Q1LNQIAKDzLlNDslQLW0nrPHDlEiU3R6dnWB+qsoUR
9IjoupBtInrQXkyYcInQCo161dGv45cMVoffIqoHGb+dFtAO7vy6H/30aRLG
xZgIRl3hKOEZpCIMb6uyNAYB3JYPoZ2l/QXvWxIR+Yi22ViUwd6ZQI2PtJSk
BE/HQCiyZ8u0Ov8VvS6en2Uw+zVNf7tabLbD/FEy9ttHqeGGpj/GTYGk2ljg
h72I6pd+1AK0b19trHY56xdx7OnejpNcIbhKG7XI0qLMUcvwoMnY/AbRCscS
FB9VqgtH9BhUKolSmlEChHtqFDRKHXxkbKBQ7O8jSKPOzB74vDVZAYm1qDIU
KCBySXh+5U1+O+Ljh5b9YC9ogOmdAV32HYRNLrcdhMDpc2O0hF3dTbuR+z/3
jSqCKqXRrLkqHAp1O8BaGIoWUD3RJYJ+0R12Ny80rgMw36NF+mzzQ2VgxVFe
oG9YqzHjocuqY2dH6tuABIB3XEjBN+PGRF4RoIrUfbUweAS8xFdv/7GZYtyY
63fO8oqLgY8oZP+d64Qt7mHCZJWMIbz4r0httYPf6lsoRxXEcrJ5wbCsWIZj
u1A4eBCehJjzf5RvnYyWS/uC8v1ns4IFAhhv0TgYy7OvOq3buKaymbC08+Fk
f6rpJ24RjI4eDI0170XqXoWcpQLnINzFKx0zUi1fIZAPPuRHZ7mW6E6hCmul
DPRirWMFRXieNvjX9tZrj74GlPFT4lx+BzCGI0eQJgVotaMkNpNN1ARqVJHw
zHrOOrl5K/+NXnTkBzXon7JqiQNrXfEgM4STN0kwtd22/xzf0/e8MvxT2sjI
rC0aDQZCJKfHUYH2b5h4HTlwSxCapPTjZljVyqfAzzf9Ipu693mnmwDteMWc
EGUdw/K9nIGJnn79LFw7PJf+2xeqow1BjhjbQYa5baEHgETOW5+VWMGud3qa
MdfOwiKIuKUad+839NFLdE/dSVRU3SPkicHWC3QIpqHoQVRhLiJCtncon/sq
n3FTuAywon9UYmR8DxqwajoFbHoxuO0u3JeLXhMerDwAz+Jfq5fx/CQ4hhFH
gaXQYyfG5SG9ej/8SpxwQWMSgBjdl7STqEgORS+mcBFVQoIdbbyWHKua6xYv
iS0Bmxu/EIgM7r58M+tQvhmu1QKHRzAsKKCpmHNWE926r/wUm/oOR48Vr8OA
LupgxqCAAa9M52Ya6Ir85q1F3dA1Z55Hstcsdf5G0BMQQDK2jD4fMVKwJFes
JTrh+CtkXGhKKhY1mWpUyxTpi0ElqOf6YIWiy4raVl6u/0nPpFHVvkSPybEa
ALp2yaxd44BYVviZHtmDVNoWJGuY5cfmz/X4jcsm2XBvVuaYvs8Hlt1aF3a2
gDRAE/Iel7f+bmXuAY+h5bvMJncqO2sTc01YwePHlzIBowmt56rx/HG7UdP7
qlyMHqWH2z5bQ3aiFwqSXtnhgJEsEh47YfC8Fp6Ypuideb35JWu3K6/5Vmq8
4FQn6F+HzVtWqo+gldS+Aw/R3vI0S3SnhLHfamzaWBJXDyXf0EqGCyZib1dG
P6s25A/C+VA5wNEjwmfR5NWz61/BHKs+bjqrVXD1nwoaWSHOKhJjYIMVPTBs
S3C8AuVcgzqP/q6CWbEb3sDtI3unl1Kg9GLE25Ns3O0rUf4ksDZHLu6ZxdLe
tZsUCElapUe4I/K062AB3o8bByCZf15iC5zwrazireb38gTqPHm+H/LLTxIJ
rWzi8uSBi36r8EuXz0SOvyaEEM2sVmXmRKqAJUcXWyMtrH7Oe5o1IPtjsMHU
40pYp8XMnifzopJJDCAR2jHLEqyBVF+AuQliGGogpomDm+q6YMNRBk5snx/g
bf6A5rTfvsKGpmBwhEsZ0dstN/Pasx7ki21FUUfNP4DrKJ2uAOTy3/Y0In/L
to5qngMnW99cwjdBOjmX7ozeUIplaG2ceRWMPdrznS7n6cqA3WZ5SN2k2GEw
ejOAwKPRtxvYCuLGOUvX3zvtzthMlrhvzuhuU6qG4SKQMb2AkshbtI3rta4k
BXFPRhnl+I4E/228JNduG93yNdpXJf4P1NFmUHAKdIlo/aZI2ppMPBNByCgP
H11Ujy5TJ9pLnHaKEtmiATgmxqco8BY+GGVmIcXYM5QGXBOnq7WS+BgdDiR/
oLSMoVo9/qVdvjI8O8nksDWvIUsJalY5t5gIfhCA0/9qrklzaf7WWBE0sNwU
/wXLX3Ide63YgDemGbPQzNwY5bqOcqZGnCA67mPcvSmRVcOtCy2T7Kau0Z8+
m/LleNJ1PD4KNDEcU+l7Z/4Ec5JwldI5oL32tKI4XiVLa4JIqEgrHXkzeC9k
Fri4EB3OHj9DKuqaKMpLFtW4oAzyoZaI6kKd1MlfnnPGgpvAkYYg5aIDVTiz
MtxScYKm4oyPXQ9YaLmQW4m0K5pJJf/jJ4BPj8lkAd1nlHFIWCXIRdW4Fq9y
rH8eLHjpNQ6k9rJjXbpofUoRjnw0mZjjJpmiG3WlLmSDmNY6jSyZsdj79VmS
k5sG+xNWlKJrcPoNeaPxbJirIwkRCBK13dDBKxobCfKsrEJkxpVFE/I/vQ6/
gxOuVIHCStjMTQuuOEcFwgljoHderi/+sLH6K+w+05HaKlw4PUNMgA/uf3k/
v8A51qcOItLdrTWgrUN/dr9lfoX64qMmxNSfIxd16jJtf6VG09dYdsiYMpAE
7tRsf4iII+lSdf3Pkcf1FYWbbbVpvcjF+ORnGdJOZoh8QUByC7JL2QbpORSh
c0YpDrQhBz9XUOYA33wdevqPOe0nJwCukGgLhvIU8xYPAc4zTh4JLrzZFFFC
ahGN35O2IBZxVgJGqVLmrQpZ3BuoljBxQrFHmOQweyNYLIiM3s5dvVB/eCkI
pSWXhnqcT1HbiwC6X/D747SVlyVgCjfUDJADZuUyL8oeBmBbE4Gu+q5pyYsu
lnSZT0WZZOPkZrfsi8x6TjUdq5p9CkBXbGF8mxrpEbvJVLokdL0fHNY6t6V0
Qh2DQ/QQNdQlm0o5YgflC/+pIbwm96jNFdgWpBtfvcqZRuQNpD3EFBW7/4Kg
9J3JIV/gvMHdqM1Jh8nG0QEsSALNIZERygsTaw8zRMdPIczemxStw6JUSehT
ooxqvGQS2kf9QoY0hRSWYdzVt7TD3BMSawhWC5rbvHD3pZIvChO+POSWeGWM
NbvOdW7vo2jyX4iaAozPch/AZYpAQQA7zHx/DxQA+27gEgGZxUTstEs62qf7
No5BfFG5R29h+cbLl6vJinyEl7bR1Xr6Nej4jHR8dwv52ZyVeL/a/9G094J+
BDR1XB8Bp4o+myOLhuCT8Ut5Vl/waJD6LPIzv/omAHCpHBARJeDh9LSvU1s6
8c5YXxi+3vUq5wecMSJN2felrsPYrywM1feP2paVnqBoqVJfR4ri7rpxPJ6c
7z0wZlfBiygwjDq4Y+LkuTuTsTwJgmQ1dWQwTVLOOLzCANmqaa5DGZwHzfxz
tWGExTc3KdfI+gMEBEGc0AjM5i82MsrmbaOKYbAzVchkceuDWoV7KYuJp8Ch
mIXin37+6t7+u6+Dw3BVjOcnvq2a1HtcpznG8s6fa+e4d+BTyJM9H0TABVtk
ci1vCy6JDlibdcdeeB1ZjmpWnhNbbq9zI0BOKtV+MErc7V6e7bZRhaFxLyM2
tUgEs4Ps6wrbVABfP5T4q4scpV0IlSAS94cqpJaomG/6qJnzGHSbIhW+h9If
eWmO9yVd0j8/tW/YdBf4MJ4HyowWFmkiXr8x3nvGBQ6lKBmUNJcvA47cPdAg
NRAFgpwqqeoYhHqBdyJZ4u5QUm/35jVnVEvitXinX6XNG/Dls223TO4oVGFA
pUKt10ToYPOybJFQuTQVLMjEyUio8UK+D/MLkcm2fb33AUXoDLuRt7sZBa/s
jHMx5+XIz7eGTnrfUdvgIHb/SmGH0Lm6EcCF7mw6KvKHWrOAEoY11uBULC/N
7QyS9x6wRJBq2qAM+KOPwhJ74+73iXDCSjv2LqIcV7GmaMMVfcJG0E9KceIK
LMDOwzqFOdvvSJvB4ZjEOCdAbZ6Ar9xyv/nOCguK3PJL6t3r0GSFYj5TLDhH
f2YM/yOxr4mARQyaore1cQISmfn4N/JDnf8c3D9a6M8FDEaoln1j4rdToTmi
ckjjYUZlD8GkxbX+mvYQjw/bH79C6peFEVaQgcQjKdPk8Drcl7fUW1oWP4pN
EBg1DQWg5aqVwco25OTKw8cW62dhQiEMnFc1qxv1nsSl9/8rTo1AbzjXyHC7
ejSPbP3YhU4oo/Vvr7878mLc0XKy8S1XJxoEE0r8nSsvAgmzb2nzeBkrMjn/
y0uT6bzmoNQSJXlT9K5r6lqFMOiZ8FGuYpgaePOTRX9bICk10S0QqhCB6Rnt
DREaLH5nfDqOvsxGeoVHYZp6vsN4bcKJIgXM4sep5dKb2yILoghbYjARUF3j
h4wn+XJivJLZ6GYS7giuYGzOjp+qhKB1ejk2jgWvnQFLf9w7kuVjQnwW50Gq
/lDDKoDFIvW755D8GE3VRawhqffPNAIv+L4caOxy3AlPMgbV8yDgcRK5l5ij
scv3helJr0bgSD/FGpo9fq6NWjGpZSFRCkvos4vwD7+BAfKHIZ/oZ0oGKDmH
BqnyZK8CprANNVECWyorHefawJqqdFYInaQAykcjxqNqHACHzuuJEqzV3GSm
JWoQaeSEXfna8QhTzcEr7OBOSz9MBOZdi4eMWGgAiu2rPjYFtybmhWqXSNZb
ymOPpi9BP5SuC9RlS+1yNy2cMmmOevlS6O2gCotFdtYJ6RINdwiK9OFDSt9A
DdwodlO9T49lpI3vtyKpg2PYMtUiNjJ6dXRC0TmTIHooEE7bh1lqrktmvGUx
fpiD3qgkgnTRV/F4FguLPNXw3ELeJuqsg88eujL6L1v7BZVs4ent6Jm2Nms1
ppNl4prtx3jTV/Se/BE2NPWd6ZFOtOydJAS4qDdhiy18QV3cgmPKeBc94Lg4
hWMXir6KK10LvGnnylJmhZh0dL/a+zrGI+YzpFYOEaiMNgN9WCQu9GhWbhVJ
2LL64dS8GJcvlnuemE02/hOyEw39z6KlOhcfWNBoeDAcnoyf/+1XICYOe5kz
WHg20h6xQGKCBHF8145Cs7VMkR7eGmhwByJKRpF7m1xDKN89tn/nqeGlZR54
RkBkuORiVE7FUSl1q4/UkpuLSX/o9C05lhQ2nho6/rCxu46Uvx8TqMfvtruw
p8ill7wyKCqGLMrk9bLzcrtNWOZSio9FmkqI1/5n2lmYdX4pXyuCgCLQv0Pf
P4Pma18xyRu4WPSUqGAa2WbDr5TRdFvcQ8tL7SBc7Xx4jUlAkl/Ohnbrkn+8
ZvZq8vqIZOuAGlsX4tvTpyA7L1nGco6zqyZju1ae08K7gAonwvGViDc577KG
ulss1PEyh0uYz+UePQHc/uZMtTNFngTuJioDx3Ru2BxfWedngQfxKHazZ2GS
X6jp5Yook9ORhmbAacKc2QeEhJeGkbwJFbSqksDjCV2QMV5yrNOURB06OIuH
wzzp1lH/yvqk6NHF/85Iu+Pp1AKKw2JzP2SSg2n/09YCIgPWGIc2nG+eBwiQ
oKut3iu1GKEzBxgL2mnu1Uy24BCOSs+5TrSwxlZPh2dm/ID31PyXeaAw9Ape
/dcL4wSLH+nSH3gCsU77H2V7HkWaYqxx+nJ+euNQfm4zf4Wl2FlmTPKTTpPM
/G7/2aY9bdNFxFTYPU4fl3hwzKaJotDnyY8j1oHwALrin7KOyti5SD1Yl0OT
ga+3eve3EmURg2QqGwBKTIgp5jzyH8MPUqMf6ZS1zXZmDzOOj+29g7FoeKX9
zgaeJQvrhjnLBlfd9ReDZwSr3fDCjrXsfPJk4/xk93upFtGzC5YeoSdfZC84
rlS0rvsCOoqQyAKv5BP6EGhKwf8O11kGgNWeF68Cr2K4ib8f1WkKXjT8tptw
9ZyOSBjV6YaoDj97xJgjYhWqgll7JeUzZNMM1rnReGZnlzdP9z+glf1kWPc4
dGP2dgMSuP5DXtjACMsxc/Rbm2H/1lFwYB6OzHs/ZLvC8vSEInK4MG0/9cWs
OV5IV29RZB+AyQfvW1SXuE88jjtJhXeXOi2Qil+m5G3++z40JH0Pno3iDG+M
pGT45fHTtcvAt3JLgsegYgop2KTgp2oWL7filtiXQEGBbtFg4cDgjW7rCkdI
y+u9+oQb3lQB7lQuWZkDQFlj4obYOLWiUWH+nk7Zf0xaC9jKZag1AVXzAqCi
JgECLu+gmBTMDpK0JMITFrd1HwuVOei8WIghAtxXHwPHMM0bRQEjtXEI1rtC
YG4ytsZzgAlaTX8r1hNiKJAK8l8nnzK1Z7+comVdv59eO4baqAf1L6CNgeoO
dZq6sR5sIuWjNCNl2o7mU6PcBnGS0x2mJDVm+4k2vArFlax5j7tJMdeu1JQB
3ryVLB18zVj2LCLar1J6XEsAxi6rzlrvs3oLfuVrT65M7/Urs0Y+IDfUSops
bngFkCNEAFtWo9i6/hW3M1kaHbfSucsPA/+/dlA5sSzSqa/Wjrl7hd1qoYNg
ewBbLW1WpUYkqacsfuHdBmNvksemvQrXctlJVjHmuouhV5H+ruyAEOxWI3LV
UGKRZhxlpnQJOYDRlqVYHjo/a64MKZ7YUtODeBUbBd4dlgtwgw+Oz9GjUoUx
6m7WM5P0hmxsVJ9rrKhlX9DlogJGQvh4rf6MGYscuEscS1hxrxb6tn3Or+TZ
/MVTeLyooShczBITVFfPibYDUSYsd7ZUwFEDaErIJNbZk67hAjftjyo5df/x
0L7RgLgmoo6ILXQGSHftORHxjMiQ5O/UmaRkSWDhcx2VdBYv1RXdzYIOcmoP
6/OSrAj64DraemxFO3HaiQYX9ddqjnvkbtvw7z1+wT7oVnxpJp91u/F3wdVf
wFgkQdrgaPqOmfGunLZZpwFFNeJ1GDSYyxQyxJ6s3J7BkJY0hZBps0Jo6mGv
RpA6wR5/loNQ4t7YqpVtPlRPBeY1RWZw14DnSG+VprV8FXVKrdTWk4FOO//+
XClmV2MxNCfevYCZfxM1Cjc4N17vyONF/DkJtVgvu9lI+GUguPgMtiU8n4OB
3Q+iVquhOJl4/kd4P4Oztg+Zc1J/coHw4TWa8DkDB/GzutR98wFekkn/GCr5
qjkWbG8mbq2BVPoYEs1j+xhsRhQP5K+yuFjr+LsRykj7+1JxxTyaZTwt9f+T
QiRYc6eqEKkWsSIn918Qa5+RWdJi+Nsbboe/rDFc+Lh0XMwne5RtG8uM2aD5
V3AJCbH4NlsUaAB06pAC52cXuERSYIQKUblccM6jxcAL1xmR0/0xspcGuls0
WlKnvd9c+xHR2SSUKnIRuw2ubTQRI2WrcWdkShW4V8xZ+crVoymWxS6QtlDB
WvGETEKgF8VbSPxZ3Xi12mllRes+r/5cMEccA2jg4QRUpUjZ/7tBCfcir8e/
wKVicB/bqYbhvN8OTHnQ0ty9kG4CDaOtrskq46/zzQTRjG46dahUXTu4sUsj
qA7Oj3bQaPS7WrE97Sq0BWvk9Ve5xARONc32c1QGvSUI1hZpauPkjtAaMnuQ
VZ5tI7JJxhBUDXu7xYicK1k9HnoqZahE1ZMIBUMFajz3DEWFlK+sz/PN7U6N
G8VpyzVo7MFM0WlSoc/rL8V3huoiicHreKUxOldqDT1abyLz82s3qFeLX5yX
oH0q+E7nBQ3jufZrHzoHMIBA30dJvnJDM5grV+6i87duXsCZeuj41WB9je2w
DAwyf5n/3nDCLbPRYj9uWrCBjf5bDLqWfglW8gB0aRmmp3ojq+sMrQmd9YPo
D0ogoAeSkXdM3tl4bBnqIkJJSl4qQAhCrdxOJ1Xr68tO3ntG2Dm/6fCx1Ge2
gIIngWCS183H4U1LfHd3UaoZH4J+EkXgXMrChIBLYMHelwkWCAQauCjLj6y9
1Ed1h23DixsJCC6IxiIU/xWDfD0ox150vOOfiOoZj+0BYCULvb4TiMCsyINC
wA+vnOHuPvh4kuJb6jvzjclGfTBNLU7NZ6my8GLKr6VoLkXbWhRr/vTrS9V7
k8bI+BAU6lMSnz52Xx6pNQQN9Fq8uIzMsHhMxyX/3o4wivLsjbxsoh2RFjB6
hPjWSCioZqKrHdrOCG77HDEoRLPFK6Y/2VonnDKL0U2wnw+CK+cj+BQO8bU2
9eyYpi/EOQNlH0c768n5QZGx963QZ2v7/MPR48FiV3yRs4/8T3BXlXAbr0Kk
3FGPtfsxs6Q9IYKGyFVir2gQGFrDzePwli8SRQGXagmYywjPyGF/jVGkOvGp
4nRpxivWrBBMG4FvX09t/JMcmR6Av8QM/UtevUTsrDx3oy3SoTQb0yH3S9qd
M3GLgNHf3O2cKdM39V89LH4Vx0or2A/eo0xfW0y7ypG0VUUWcUZ/pZII1UGe
hPAJEgZTWINhSxDazK8cZx/3mpOk7OXf+5KQL/V6TBrMjrMJH6qbnloM1CST
V9T9E3hhBYI9+5SNd7hT05l+lX9CU+WwNLDOW9yIzcEjoKqm8yHxrr8b4UIj
iCrGrdSJtkcENldMTC1nspHy3PskvXOxKwS90v93slvJHMWZ24TurrMti/Tl
CqYAeHeoP/IZH81IZtUdbfxaaecqG2zQV24tX6ocedEwm4g6WmjZGuwFm91O
/JkCPRip8nVWVD0uya65946V22Zoiys3Pg6LUVTFWSAws5Y+Y0Zl2irabABn
0fNLiSmzlCGOgiHbk4N7N+qR9+kOVg6zB+6PXaukMvydvJ6KHCYtIT1sD1DS
IxUXl6YgA/Y53vF+iV3DwLoT1+7IHwXt6e9NcIe1ydkNeOBF+mi8Qhh0fnG6
CzPZZeuWk7BiL3xslQVTmLC1NFUkTO3pgmNB/Rm/w+5d+Hv9y39RMGbOCp5Z
cSPfy0Pdqp3mSvhLPPLlcUW03bAi+P1OdyRhhh0UNrH6CPiv6ewyiP5XCmUQ
t+SdzikdVjl9UJoDoe1cXu09Ikk1hDE4KOtTDpivlazhfO35ekUlVqNflSqk
KOn5Cy/kWKxlGzDedksoXTIg0U6EUH6PC5p91r7IS7Y83VMcig5bhWbhDq1C
KtSKPXij9u0/hY+EiLHncXUQbHNTq9N+BdNJGCx69TmL2Rq92TOQJvFRbm2W
oZUewzJeyZ1ILikf1wHgMjaz95umSLTP67/Ue0lazEwYkbox2BEifJ9XC6Nt
takKE/L8Wi1NanUm3OJwiXx0L1rhGMh0udJ7e4q8s4xe8SMAbJeCkl+71759
JeYTcBwkccwRcov9efb2Y9dL4aJONK1d/EylW3qX8AG5CQf+EdIGZrUD9Xio
hZiv1m6YwyOwVposNvmWKD1kuOCZJI47RFSep0uZFoVYjm911mCM+xlx/Xw9
c29HAi2TXN/IIhhJb8x0i1s+3A3d9eNQ42Ei5qoPfrZR/ux9CqCtxozUP1jR
Oi36NCPfHJJMijTDHSWTaDlHFWnlXdMgQOGRWGw+kYCctn5CN5VniC4Ogd6Q
NQ4FOL6AlUzWlZPg2XZNJsFJpQvx0Pty+7/2zt9KyN8VZMf6LSRdjlwUw7YV
ZpM0iMaodTv2P1nKfHyhiki4+00543QYCBxYuuAbBj6Jj67EsVqIkxNDzrdr
548OCGWcc7S5W5+qL5lR0a5Vt8QTxjYenuFHVYNdujcIqOZ0oIkSiMI8HQUt
bKLLno3RpuO8mQ6tGgxXfRd4BSRfmInDx6EKgzkdenhx6WqxyMSXkuTrXG01
l4le/6gEGQK6xnuQndVVbOBreYsKX0vk9DUz9HzDAQhGDKWYqPtu1VbY9Ccb
zm7m9aiOJH/btVy1PhCOvr8zFyji5SwOHFhHnBIzPL5686HMX5zWC4hXy65b
goymvF+4/zvY/OdCRLlNiLBGBBSuHD9o7aJfy+pvEeCB9a+s42k2wlrzlVVH
KWZ2eUCDr4l7RM6Lfj2kXun+xysq3uLDk8giDZsjR2PehqqLuZPheOZdKsAc
YCrYvVvQ5mBKSVvRjr2A+0iyoEjUmo13WR0NefeDwvS+BHCWdV2/tKQ0sYsa
CJCBe8qwgHh5uX4/zMtE1wBu2STfCtM178MhRBqtdR+RJrts+3wxGAqnnexH
d4qtEoJlSvD/ZDe7/DbXEZpy7NpHW1IkbO2OGq7EZjrhjuZ2ECx6ILww1K8i
0tUT3lgHC8U7onlWTl+H1TiedstuafC7+i+lO5aeyIAkaFxVuRZCmY6mB24h
zElogU29nHrNAK6PM0LGZ1JhZ8OwtzKGoAkHm7MDmTlCeXHlHThqPEFk0jLv
Kkg3DGGP0nx0IbadXJGiC8xlt0w20sQc3CTfL1XlNn10fhUkfbEtkcQkFV2Q
koZLSkgqBP+J1SjD9K+Krj/j7ovtrnXB2iGZCkkYmqdfK4KOPM+679h5Dx5W
xbWVD/EO7lzTlzIhh/KzFypwOtIng19r2Ng3YbrgbM2DBoqYXREmImu1DMjW
GZhwkmivbnvI1KIrJpEHYDWjBITAHV1zHVgcTULnNYb590UBSGOwocIBfMLL
YngPIRZc36yHlzyURrx70uyc71oNAI3TT328tcCckT9Cb16fjQYUTojHBExZ
7p2Cckj37EmycIxQIY+Dh1UBhyUNmT67eQeocwnmLWccnMXmceycKAPjkl96
gFQuIJWcOdNNkJfl6oyL5dfvAkiO4v6FvHFuEqd85ee9YQybS1hvZ0KNzsBQ
KD4RKm7a2WYrB1yXO+QodvsYS1CaV8JP6u6DS3Y3X/nDYfMhqrJswpUafifo
7UDUozuQfD/wmUhCd+PbRRNS6d06R0IIuTmx3SjQHDD+e5h3bwyqT2J0pZ97
uHB9FTIFMNjVDkv6t0h5BcQWjBKxyx03swVSThPhGi/aHyz9fBtiPIT5tXkS
7cplIQ0zG0h+kqkjj7tj9AwkSnW6PvHzo4K0tmsjvqGBt1J6L2slaqrWvPHF
c7Sqv1g1mgG4S3fEt/tilKTiCbufLPbYZQabcKkibNLZVVpp62NFO0sGGruI
anhaVFhTJi7UBHM2H1BXwA9H8wCLCH24XahL9TeFclf8Z1Q2dCzgO22plzg3
XhA4RxAzRKd7DECHsbnfvgZQQIdg5Jt2upTemN9OAE9Bmyy67c+sj1LBZCOw
vkjZlzh0kvnwzM/qt8ukITQBdzSJsYdBFvUzi5hqDXdmZkYB8frAmutTmu9S
uiBuwoPZtWDa2pJEDXzMrjxi1278kseiyz5iJQ5NOtmUU3QhLp023mOEf9cu
b8lwFfxvh/oPIfDdFtPH0buZ0v74YJCOMwnnceI4B5X6LGB1FI2E9sMwOcGQ
TwLuswBFTSTCho7EBGhL19hIIiZm4BE29QMSDXxcHSHxknuVUi6ez9ejIf88
V0fB6bGdZcjDPLNhI6L403HSARr2PO6ndiPLOLP+iq1kBhZgl7zAPsKZebU6
jo9135SqEDqYeqUcdelL1Nkrmw8zpHukE3N+QURjDlW6aYZ/xrer48zhb2P1
4qUk5ix0H9s2FYpEQdEtgBJ6fk88UppAuCvjQQ/850DCwOXm9OHwvtqlVREn
p7yAZFtN06PZCaLaABFDcgyi00CR91rptGOkJNoo53mVzwaMzj7RkQG16z2I
0OJ/vYfRG9P5xUrrjn5m0pcKGGVJ1leatRSl1Sy12SIjML+lpRUlE+2d38yQ
c02OAZnDEhPMBIWiYHItrPDIKKTaiZQUkRnKdjIlnOQP/03cT90ONLQafEQh
lAoz6CKw7oYUnY7K97XBVv0OZEO3g/KwSrvFIwR2PuY7Ri7uSTymBFYaUxPN
ekUtcVTfC9RP006LWZo5VX3e92ckCQj76AKaEWBqpAadVGOYIskPqeLu6Ql/
4BWhxeBJm4TouUxui+Gl00sqHRpSHh98dm8xXhjeS8Lxlm55CZw9NSe8rlZO
OSpCGz+x62HynZd8yEC/bQsuZEjsDFO2R3GfmLy3dvO5BzEqUxIixW37UIfy
jsGeO0VI6PUrK+Kt7DJE81slAbTLt7GtpTrha9vrcpGRTULxKlnK2RATkl+f
YldrpB45a1wDUB6PXgKzV3y9bmlfciroNK7YbUz3z2QKVubeiKon/yeO5Yew
BMU3CvZr1eqWBVP91Z7jlKSdEFBv3hAFrhKxikNOBRxkxcsYjbMH0G2dau1o
7jQyzpb/g0/2MGKkoeM9c5BX8u8PHlErHu5P3LCur8EEhJevGHz7k+Xlv6W6
p8dZUFzkLRB/+fM588EfhO+obiUcncoMuUHMPLxXSXcUrhJILFhMlv0VHu+T
pWJDQ99TxAQEgx3PrHt4AiAHQPXIbT+/WUxZPM/kE7lqZN3n7qxmtwMnKq5+
JNnlP4jkrG6k+mGD7M3CRghCvsaB/7TUWefUWVhdLAB6h8l8y6fhUI4wva75
AnY18WbjCNByaEZcRoZlLJv3DNt/bytB5OXZw0aK2UnkfLY978GNr9DBExDd
OICgkuV94zGZO2vIQuYMKKRp3aR3T9MXs8B1vJURHJPhqqrziu2gwGp0Jm3u
J3bUa6pRjs8YrlUlkyJh1bjpT6wbriEdTe9B2Wc+Ts8mSSoZmNBEloIorwu1
5Kvd7l9FePb1QOlR0tuBMnBJ/NOFqqGN8nNZmD3RebSjMATPn4YXqvhLJBHs
VgeqJgZYmsGFHjzI/FE8zdarteGgwyRczUL/8wVtM6QP5VBI7hg9LALJl+KD
cJQO2sXoP2wgXqwF1jsdzSMPfi/ENDa/uEebTtuosQW2y9t/3V6cyr9cmp6W
rRG/Nmf1tpxbn0lY4BP9S6n2a6rT7AUbrsu462NszYfuNMrT9eU5aEpgaHGc
vTQPwfdQMlYDjTHyi77BP8pQ1D36ETR/lC67eW/kqs4XyuGhSMAvr3AIozoi
p1CEdrqItQ0EKcOC1A5dYL20bFrhcImBFZQ7yFDaSKGt3VBuixNvGXdIOh4/
OyhSvuPp9Tt5P1XTWMJAJOsz4vdsyI4Dom4qzADxlW9aapKOmserF6xHJZnb
MF/mcfL5PTio5g3J/iiEdFUkkiu/xLIlqUT/gEVhGwNEHziwBbfxMPdvJ7ko
CcefWksidL1H0d4B2eIb2zyVQjegRctJ8KYCXWFmdrBCarhxde+oXFsFgdZZ
+GFnS9i7m3YTEh/gpr9Exi5ovqBgpnTmkzA/B5o2D7z2fY2ua2b/4h/uKyaO
3JPAhNlHydVGh5XUxVOEq5/u74E7s9mPcxObqreS3a2iKN9E4LFQ2J+VuCeL
RA3vBzUiOCQE4oh8/aKnrmthZyBpqiGlVD0ByVJuB+h0qMHZxqn4k7KcNk7M
8AlQifZ6bLTXzI3PVqwKKhpEOP9IM/33qyeOktzZqGZHPhqz/WiWKCKpiM2O
8F5eTia2G9x1yqOcnSj4BaHdj6DcwYLTkdcMYJ9W7xChuTBFR3dbZnGvVqEX
ULFVG/MoBTpSuzLWZe7/y9POncyoLAiGa2Q/EG5ALJ1jSYsOnhq1C4jFzj/a
yZS7jDnfiB5TG22F+o5zfH8T50CF/J/vtdI0WZF/R39vzKogROp6JyZTVnmf
ZQcIBuFVYOGwePMOUYO7HhhVxwGiTh2Qvy2cMSjXWz5eN3LdX/27kSAWQYDU
nZq3hEnJoNhXXQPuRZZYrhMB3Y2w6N1U2vGd3NchPQAqyiGe/wg8hJ991m41
SPl92kYLF0FL3v87Lu5aQtmatjTJdcyRtRcAD2g9+p0fX2WLCiyZalFVptH9
RxSBJGTODUG2qeg3LSHmy5M/s7zim8BPteLljqfXZ8QAU7hIotnUjPLI9to4
AUy8F3VAWHnNPuUZqOQ5PlWzvO2djwvnjoRai9fK+a26y+UTw1Unj3T6qByL
eDkVUeVXKFHIbR4LwQrzB0TuhbZQPTCPbIxdd0vQMIdIxL1oGv8skQKXQyEO
wLRi1Kkz2gCxBw7clQFOytc6zBdeZwmtwAlCLE2e2qQAwb3kSQPLGs9Q95hc
ujWFkAIKygatab7QZdtxeIlXMdoQDe0IZONMtwj2/CWq6Tv/xy/p+4y78C/H
DnIXsvyocRNyBXbF0iTR8Af8Ydiu8JknyU7XPUNoITjEuUtwWks+YMXhzcgP
B2jPUeTagZvvgAYf+1ZnNSzCWvgpuvFj+uxId3fIMjEUUZuVb8GG8D744K+A
taZ6iX8SEumO6lVnoAB0Tfmtea4Yv+xsroRfo+fdtn+81Sks2fM2SE8kImej
yBIUnu5/ZVSUgTIggI3sxIW4iG83LwOT9UAZXEEZDqgG2yP/9riHoaVZExt3
wRfbRm6QUNwmSg3yH4YfQSOszClKs/1Rp7BNOqgq18boFbvvLhVnjTwfGykT
uzzdYUKmgAQ79j5T5GzoVbMV4Rb9uWp18uTFjVVsuruTGiQAnjbXoJY3+xdN
unxdAEQ9QiAjRg8gVFEvIDgSf0vTc6ypKMoQ2NmQ7JN6zmzAmVhWD9fM0VtS
n172NKRxAh/BRWb2dFe0rLSPYq66fIvyt7X3myuv1nJcJgzznUNnvuCFrfP+
9kNhBd/ov0jqXaaD/iASo0qLvNi5zVyFMmaOzwCnwMj8YTy1mNMWo/Tmnlkh
uO6gLE8LsepLXxqRzcOQVfqm8rWAdMszC4E8fLMH48SCUpcqsU08vsUjKxYt
jEfZchAxAFLb4vGOWhhkqBp5ox5UzcOAoCKfZbuDgi/6bKbA3ouWvgQMEAPx
TNlrltb9anc7IzOsYchkQog766f3SgKtd11XwOgbZuBz55ueCBuLHSDsm87F
ykZQD8OzQBF4izSInWGXXjBMMSHLblY26b6AEMluC6fpW1QsWc6X9JriJxZp
1FMNo5IEbtH0j2RUxlqcsh5i4MDEZRxlHr/fSnRzxEzimOh3H5AkMkgBU1kS
bR34NrObXZgLPdwrif8sWx4LdpCt/q5AJGSuFBWTYvYzqnHNoE4sTzu5xnk0
GDlMMQHm0MLwvZOvlAoMJ/s946a/v5ycA6j0KC2pfBw9YhUDvjGR9ZhfNiFY
cEFTnYp/eHOX+J+zYa5yZOAwYtKlX3HQRepxQgXYp44l73GTrafkkbHi4Hrp
XcA3Tw8DHD7qC8TYrCSn7HU1Jo/3Unl/n6emHMQDBMzGCB+aD1WnF+ZLNaGc
jV1cnzm5ZZwcGDKset2MF2hrsu45jvIPvhZvt+fbU2qf9Z+GY1l6OYWN11Pw
pQLr8I5pWjJpypvnHHWix+KnJscJGH9M83xvuwtmrnidctdJ1yzbwuN1MUMt
L/Wpfc55cLzkSvUU4iI9E52vraY+gcswz80D5Om93nBNWrE0WVdASdBQT2Cm
kqo5DeRL6fz+JUYOAlA48GbOylozWKn3rhqYaM/28uxdkQdknbaDe+m4u+s2
+AR9m16nGwNeumLaHaV6fVQjQLtVvP/2iGdaqAkXKq24o5wM6nnaP6EMnuTB
AGmB3CF6n2KAvLq91ZzGr9KwqH7hBpiFfBrkZg5KGtngAWF4vGqEoXhmMUfH
Lvn74GZWUx1tqtIeslaagcswbvF0wI55GxVnKBMxG0e+ZLz9VHsnNuZ4XwOw
pOPe8zwD5guoZezST+bKQhNAtW1Qdfzcru6PZsFnhAlXe1IkRjCneTmqU1Gn
ZRfC9s7DwrIQkuP0p3TIAS0AE299vyP150Zn+fRuWPRJz8ARDjFkZeJyHyFc
3D7/RBhj6G9skQm3XcXcnzfqMohHKW+aEzbbE2DhOdjg05KzS22/cCjgD08C
C4MyqI18eMTkxqxY8CSG07J3LV2fGhOWumzRk3f24L2Afd2nT/1sEtf0d/j4
6tKt2AnZoKVPWN63uRkqwW3PGZma4VFRspfFkFzuT24PbSBHLhPE7y99uKKB
VkfbvM5LDoZ1uuNXFh9sjE6UmN0X1IHhkinYPkgi3rhECTOG9O6+uWCFpKtd
RVgTnMcrrppp88lVMp3+aFhMh0hsP03l6mGLQT0nm7GsjAaxv5ZRNRgayBF8
sntftKTVULewUoGd0D3oLQPo6WarafawMGuZSJqKOMbkbOLEp0dl05WHt2gu
0bvrO4xL1JNcrI+2dspmjHTL3a9OkyAaghRUOJBio+iU6FdPXBT5tYTsrVnT
KDMlpHsLppeXwKW65fs8qcc48vuUd1Fpq+SntYgpGbZc1j5PJhAQvcljV+zx
lfWCueAKDUeui2LbgMemVbcL9Di2EIgH0ZBjnaWqUrtwDrTdhZdCL/Pps6SN
KjmAuL5E6CaHUKNzXMJjXQUiejWhXfnH6a+Ss+f/W3LHFDyNZB+KC2+/cytG
bBq0ixJcfdzxhMpjFJ/+jHQ79SMVLi8e4oVvd28gLhIa94eaL+7CikXZ26f9
ee2/Nv4bUbCS+KqlVMdD5irbOVZ8KSLKuRh2xS8OlDKmXvYE9RBWnaE87eMV
YOXu+WAMYQW9bMdEczZKJc6WnrYiUzY5lEjnNeypksbR7gs5iOD9yjAw408M
UWwZu1wnnw2l/tdoG+LJ5w0+OAGta9RVsYyPQBkA+Lo7Xh/JXRNr55v7TAFr
OKlI4s70lX7Ui2zBI8pEyOzoRrlk0XoWPUuhsNHkv/fFxz+v9bqHo4LA1zNL
wYo8g31Onu8Z/5YMLJQpxEDzBZ9AEekJNKI2fxy0GhuAQ+jSuHA9zzVgyWS8
PQFEgLT4ZRChVQmf6OkgmVslNJSQz9FiiENFd4jDF12E1urUGqeDpMUJPZkr
O6T2TNz9gfYhUCQyiBCAOgUmLbBqlZ0781xLzSyXxGTDkNp+PUBZQPG6EAFs
qHpxgv3cG/w1vrT04kWBxWLyNnMPRdwRzfh/QKK23VoDeeZyyZnlVilnueg9
SLugIgkQzdK7x436ecRB6e1FDqF8TONvIOBTeFtk1LeD1JTLGxSqwwmSkwbC
3aQg8ZuIxfGpvEqJUSW5f38nmFEK9aSKTspqUUD0+Z6Iv/zpO56RtCRE8QMx
JG8r7OnNSuNBUg+9CRKIpOXoA0VNl8lIwLkq7jn6n3uk5CdI/v9exZkpSHBq
JCpplb6tAa2uZlkOB/YJsZdZTP2xgSu1VpcpsobWdnipqE9WZQY2dvGG61+r
ZrR9zeUPwikcYc/UTKDgKsfLIDejvk9J/7yNxar6jJb37C5DsQs8f0TdRyhD
A/7FAvxbiO6IDGhnYSBkVdk0R9W+kspcc6id6gK1i+atu1k84sfjbrvX//JG
4hoPvuhIMg+h2kzrjW15uUAK/IRfySXTGx7ZtVgodTS2dXPKn0bWBUH38faZ
DSI1E6JOV7oS98c8hm+vRKZnzhb2a1R6VQyhIdKLqh61kqim5ErcJJWLPcE0
LVR2N/MppFRbVel4DrRIoOYXoM/gbIHJQoV8rJdJZRjDgX2+tzNIW+gBIDKX
jexFuqGbXu+2/wMoEAgSeJ9NK8Zwd1kxdohasNnUm/2MUWGOXht6o6dlvfjM
0ZCnhwRddycjXiM8MK54iri74Tol9aCam820oJaCtBcYG9cga4iCpFN//nIk
DevHfStYqbeN3K5y48dwOk3SoLh0Htki9CzIKwfxls+MJ4U0K8dzWJA4xI5J
/Ac+P5mpfowWkBWaOyiWzrdcFcP6tAfBamzQO4tFJ0f00+axb3CyWMLolkXg
Aab2W/MLLFdQu0fz6PRR7ta9XwQzv9KqqQarN3580Awz6zh9gfhjqi/Om+ij
/1hRiScOOpYj+y1VPfqh4IBpejJO3v35G+XdxoyFDJIn3l4S23mgu+F1d/iX
SmIqJKjPqSHB1wAUJ3q2QLLP1s4xf/XRKgnSbH0Bupr/GLZ9SufFPg3aUiCh
Vreix4i6jwpbpyBIAkqTSdh58mj2svwkgOnRhbWVRf0kAIaVtUAUMrUvxwkL
Tw/XeVp9b9QHsmgtctGC86QOivCm0Af0EvqhhgQu9wgR540TMbrvS/whGtjS
K70Z6KE48EI+8xsnjGGjSONPPXPb0asJH1xMkdSGrUVp/CNLZIHTPo4DZ/cd
42pEb+xdW8oTkCFIeOVLaZQDtwqJfDo2GTMJ8Hn4K4BDbGNRkeL3z1WEH8HE
XIYofJnMUmUr8ok/jgxQVjO6sH3u7qBzsazahsiUemWO1kcmaieoBlJrZsRS
BH+R9nS09kL/e0CB+sXZeW4q6wkFy7X24mwhJdA8/CPQvMXas5IVvVPI0Xwp
lyWRSPi9ftY28LoocfmUFYCONAHLnbsVwEo1x474SlO3sOSxfM8BHrZBKcIO
MMbS8qb5PX5ri6WvJIpdxL9uTQl8nAr1ExRRjguX/n2xFtU1T9K1+5cLhG2V
Y+0WlUHdrWbVqR6jIezbAECEEJDtvatxDnaiCJHVNrmLuG1gByH/Bnh2uvK8
e4LlvIYg6mEwrkW80JYKWjThHiL7G5TntXCMP5KHQtbGDTdMlgHjr21Qnb2C
bVWyGboxqUL0/Ym9Nu+a3Y60CME9ODQSbvJDGJj6QMrxa+mF4vndmdZkVDvz
UDHVTJZ+JZgaOQCVO2C1kzXdoyNhnVFiU7XTt/I+YPINSfClWdk3XlmwuJzs
c15wgm9MPzse8caYLgX8kO+1ExbD10b3vCTgzNp7BbvUHIEwwyiGFDTU9Eu9
JPraXXJhkCIYutKWu6tQ9fLSI3RKDZknlwc6jJ5WhO4XOELgAQzbnskosW2X
q2wbVD8fODuU0aEEKxI/IYlSkOmdXwE1O0TuB/e7WkwHyFVPDD4ZEyTDyObL
3E/RKfNmOpzLW+UFkClNHXPAcrl1jCr6olxpCWU4fZwtPFOZPtK0ze60E1KD
BXDDrqAhKkKjKXxv7cHimGoPYNXkHdlVoKa4LFDiBAl4MCj01BIACEgx4zmH
AyQ8EO3MS9h6DS0FcQQvYLwgFvPnLgIG0lxO/n+/YW8E0+hRaaTOPZIi8ayb
rM0AJ4l7GfRMc3DO0R+n6D2HWuBwnRgerppWdEtY0HfFuhkGVrafW5GjzFtq
FaAKtelFSriAEp2xxWuAHjz2OBqhrUufJCsO8qncdVpjRmZdQi+f9r8bwbGH
TloXmfQBlCZTDCS4vU2M2EdC8uALM4U/ePQm3meooKsWFADN3Utts67ZPNbC
hOdyk5jJkHvR8p2rGnfmatWTFjDXjbypqheGgzTd0t9kEMec4qKvNyrTaDI7
OHCGHPwowx01fdlGy6/wRjdgnXlSWOcx0E+zbdtmCbQGXvMa40a121H1ZU8d
7HTHU+q9ulfatp+JisdG4knglyt7o/B7epGH1+2FLTyjmdzN64MnPeOotn4f
rE1oVJ4XfjyF/etqH41asvtI/LJmUkMq0xT1rUZviQWc2cqbTjSkywy2cTR9
ePIB9fUH5rnjy0M/nZg18jC6KCN2EIkfTdRHrNc25aEE4xYSBA4n5rSA2rSI
uxHPWbPqGQ2T3a2j+IGCGt1tTPKmPhtAbDlv4YPKUYu8b6kc6aeHbR1HFXFb
LrUktrmNJKc7KcBbCSkmemjh2Tpb0H3YtSrP20AikQzzTZkkn90ymCPrO/RE
StKChjzjzqSe1Ble9L3ObuWhO4gGIVz9j5gHufLns1UoLOtPGBYCwFUDBkB0
u9MoIxvd2TjdKo2F6xTLfUDZ2VMSBuc+H/3cOHlW7FsUUER2id7mVRH/TFh1
gsatNEmfX2nf/59zDpCOyvw2/rMsOn0fkQ69KzxTHxf8VHJS98EpeIrNUvlm
LcfTtDCyQT2vNqTQwUHy+dlKxy6Yi4NUIVQ3fTB05fqEZTgS3e1fLM9fOalw
XRQKnZOjDYPSB0WlndD3DviljSCZFM1/9ilJmvVPwCYwgEKpFbuKJOUOQXCy
JppKJeQw6tDHDl7msfLYJ0YjBJjTrYcJicMipj/hO6ma6wLkAQ2+Oztyvu5e
LVewjxqczH/MM5BC2UzJQbIwH1SohIxI8Aahl7Wz1e1jxiIwYwjBE87gfg3g
ciWjnsy5fIvAniK9bwZva+m9ROxA3O/pOKMD2ORlfclsukt5c20M2NUtE3eO
taQvltVGK7+bcEesVAcR8EsxwH4mB1fFLaKeaRNyRLeo0uUy5dB8m3H3j9kE
0MNR4JIuPWVyP6MlJofGgW3TnHtvVXzGMOwgPkBPalLzyl9GIWxDCahOw/W4
0tA1c4UwrhWhfrI1G5bkgwSR3Jfk8BYk5+8kD2xw91DHyIWK9EeymjMrhfxz
a6eyr/wyUTd5bB/V9qT2X/Q26FejiUNKUhPLNyB48E3Wu0VEHAfaF8Ayw+MH
AhSjo2jjcP69qLeQLdEt8webqINFF3IsjzpbtTgGDmVKsQ4IG00/FIo1OZC7
uQeN6fEK0yVK5t4DgTNJcT80VYA8+TfujzA7B7jmVDDE+L2P1Nr6lZvXuhv8
Bnbtr+UTn6Rwet4rvnzBWFNOsTG1/TcXFPUwcBuO+Huj3WiSiki995PfeEXQ
AzeSmJSEqHd/W4+TCIaxACz+wplDwWUqfZyMVNBEBAh1+OfBIfPmv8yDduZT
t3KVtYRqx/EdLdChyJ8Us7FDUVtoNE9spg0lleCUOwiFU+9cU9B5Ftfs5f/5
2CRsSLGJZOaODRPMsnJP+nssHUiOzsSiriv9xUHBy9UptP+uufEwIEUSX48c
O8UeHZ6muYvhxiNLPK+ncV4I11cpGQkK0JiHae4ypD7hDD0iD0SDsUSdiQaF
SlPLNeu+5KYEWZ+bBSMxL0hBu8Q4cR3IoGVOCaKrSe/WG9xsl+kND9OfxmDq
L7klPb3K0KHhP0hcCv1PzpmlKvzyyX9GxWdYZy2kdg3cMBWMoZ+G1H+JVb7H
hPR/Phf1JWt3CNU8Dh1KVSdxLxlRWR7UlJmyJoNUahoYcW40jWSI53uupwyD
cM/aEcdZCFNwPxAbRjVOau4Wh5NxjtL5qgtOqFswdg+1hWeWyo8rAS94/AuI
uBzG3sc7ze0f6GZrkoFl41BMklDLpYDf18NDKTdlvYT+fAFthpEQn41ppx4U
TunA2aE/dz+Vv8gd9695/PFlf+mot5iUFURgjCmse7hcEM42cnhjOOkDNJCy
vT1r+sJ5PbNCdeuiqUSYRwgq4QHrshIMdO+mpqNZccGmSXnmFVxEOiNp5WMK
sxtdKEakmRqp7xhY/Ybtz3RH2XMoe9lOXFfr61mvCuh+4HJskeEZ/85+0GKJ
sX2SiTCcT9n3yTJe1NzJOqhU/mSfDCErijw1QI1cako4CPBjxbm5GdVkX5i1
3gZN7E9MbcJakve8uREhMxnIEmHMk3MDlLQNX/AeH7FV7foK2VICWEEeRAZx
Lv3+A00GBpV8zqTvxSgd0WjoNu25C6ZbYC4AP4LQbV5U2tl43YSeQA9VcsQz
adZ8y9KmNdpbNaVCqmT9Z5xhBhznZY2JO9jMQLC6H7LKzsxLr2QiQ3LG/OeH
TsHwetKfjwsrqhMBGNu1g5oL4z5lZPT7U/pVROEDLhGnT7uD5CkJk5nCUFFK
0+CuqYi8C4ovQlU6JchVyZaphZCAgy3CwFEnEt5kes9x/oOTJiRJR2fHzROo
KOzrcrtZYtkZlH3lNyiKLHIdtXFF2iX17inLB+BL/MptQHFYa9C3cbrHaWm/
7eyj6ScSk+hE8maoMOnz2/YA2uvN3R6JazJfUj4xu+PEu3mwmQ1XqPez8fFV
XxtN50NGCVxY2OzkA3t11aghBdPduGYM+E2TZV7AGXIFBh7yiBvE3+z53pxl
vrwOJ2n9w8D6aGiU5q5Bo/6Q95I5nDetIuJ/n0ozKsEfBrq5qWOn7mvBz9lp
q9bBfOFbYBZggw+nVxtl1eQLqVikGlTMaBgC0qmKDJVuWNWZC4y+2Jk28GWN
C/gPEWpZ/V5QCed3rnSksDPUyT5TLP5z8dRz7gWwc73ImGH6CqnlFoFPZTDi
piS9vfH/PlgoZct9LI5sfHzYQPSPPiSnKDhiaU3fFTiXzHDUf+CofjSsIvkI
JzRFoY+mEjddAqedNwXWUS/ReuYlvqMUeEukd4CbYdrQOwWziUQXRaJbKYdE
6N9H10zwNVlZ6YTvWHlnMKNrs10xFp4ZHIe8ODaIZaem7g4G2VkS+dRaEFBu
EH98OXjepDKcxzXDa8aAJeVOu/ZiStECtxfr3EDFacZBAcQmE+td/IQNJ5ql
tlGCdusR5WAm4QcPRUs+MJRtStCaYzpVcR/8RCcudPBIcmgA0C5OYojBTmv3
P/VSvySiu5XzxUk0wirHvnksEC870ZOIfTOEfZntpjNEfbxg9dNDDcuiDqIb
xKa3AwW4H+XYo6rLi8pn3UPqK4+nubU7+9lbZKxrUeIKYiyipvuxNNFq47eJ
uIdJSMKokdT8bZ81bGdfzjjBZZrPqIE505WY4ZCmAsnN6rqqGPwAI6bx6wAq
hgnDa9Ccn2BsjMoluB+MeyDYUrrRonLr35PWviFnPDIg9VKntzjOerK7otqW
kFRZWwsAEGAKUcgZZ4T8ConETCmehE7uw19AjeJcZsuXnk3WSHYJgCkJtvH0
6u2yma5mKT3XvIxSQcNDCjkPmUjbfizGdDgN6b8th1k6L4TV+EEdfZwYzUtr
1lbPSM1CPrM206ABXa0LR8YYYwRqsq82IFTyj4YwGmIJIHfZxYbOD8Fsj9kZ
hDUzthK1nGR7nrDBM8E+j/hW8R7LpPIv8dDBShjRiOZCONsozLt/oSXQIVOL
R39aiSqJgKfHedp8OohfBaavmohuymaELrsmJ2nhWXt8Ls4hoGmg2l3NVwwQ
kSfDAAEMp87YWDqfBdLUNLs5vr/dHKPpN4Ab/+rTtt9HnyLCo1aBmB+KOeGw
eVId0DDCCDyMRVTt1sM4vQeqs7UbJDTljfNQFf/zLiuPU4lywB97WoNA8HE0
1Xz6NEHcLu0vt5DUuOiS7fiuboDteySYTypa17K7FsGP6uu8W4yaMriqqcyg
l3g6sPS+viB8OBVQdcFj1rNCTnRLT5ukImVmVKHWPQaQQiE+iCTBSOt+zrSo
vHDm1TZz7G2ZMdKYiQxxdq0ch4T6OmfE0TbsmlTBYtVikdlJa7a8X+GJmW/s
UvSDhp40nkdeDidJ1BwZRYyzwDsTr/bM/qnb/JVqKAloGc/7yazaZHySdSgb
P3a1gb0wOZnU9qs5Piu0hbSiHb+v8qxdlWQD23slF66n5RrCKEG9iHC80sGz
rVQYKYNAa7J7zMcWThtSRm0G7LFDFNhCkRxaNA0tt4NTKI/6VRYzyObssEyX
1hOsj1CLb+vomuDkzH488N8NInk7HZiiOIVxOKcFTbqpvWFskx8x3e4XTSk6
40Ye7meE88L6vlD+vaRK0JKo7xp5j9egN/K4yvEuFcY8Gkld5J91zTlvDdnM
KVRt3p2HuM9ug5KOCjNUogOZjxZ3ArafLLgikdqM44uiSadIR7Zk0ATnggFk
/3rfyhbtHqZ3vPAOR1PrUDdlaZqH2mQVfnj34OSWkJAcxU4MOUeIlVFeb4w5
cDiU3vbVBcuB7PyIAedmfnJ4L0rXcWc7YcEcpB6cFC5dOQq3yZD6wLXKCJfB
YZM/F6URfdaKR7XHBuJndw40EFUa8snyq0QAK1oftTuwXkGqiWmx1g8ym4By
QLEBvBWe9B6Qlm2nECZ8FvOvjplsXTZoJ+AZDU2ZDBVWlE5r4axsfVqfX7ER
EpOafw/65kmR2TXCtE2V1TpLwK/uonWQgVvjDYiVEHIamyZ3qcWhJPxlzOBT
LUwllbtV5xOwBzO79uMNkZ5+IdjhlXh7O+MTQ5Cmeg5ZI1aLgJ4DsPwU2OKE
+46SEGwkcaQAdQVJP1FteM05ZuVUSFzOURnNZ+YwBKu9A2EFklXhY5CP6Ny5
Lf4dfslQ1NwAW159a55Sr0zPGsAfxoOumZRqdNkbCdqU5v7v74lNMJmJBGFb
coisp6XrXXUSQUM+ZLgI1Wpbk6mfRFPU1Bn49IYQJ3cvIpMQtNW/tw0bFCOO
GN5fIh+8uxslxDoQEleQ2kiggCAHJgWR19CFWSkQZ3imq+PjRT/wOFux+Qgr
FTgTLVz41N+tLK/iNezBDgnOF6L0m7uRjPqYV5G6Ics6c2WbDG+nQP8Yrtxb
mByFBUtMz2gok50/LmWtJ/OLh8qK/sBHxJVHRU6RhJEqQXf92yuQRVOWJ3Lm
tK18KiKygw1EspEtJ7IyKq0sTK/71IWZPIzXvFHJK1p6IST5e8E5wGpCE05K
iaEvyQw0RlBM8d+OTvAIoBJrUV1cByGblbBRvWM2GqIICMr+7tKh4r0FIcCD
P40YSIzlyLAl2MHmle6XGLEUVNGl5R7gwib1S3IkHjvKfmbkzXBAyljaYhwE
8gV2VGOwY6KWXpWiygHIOtDuJjokutXH6umdINRZj7mMbRILyXzNfiYTAURM
EcQlPSibwp0DRVTaCj6wUliKAqiMZe/JthuFmedAPYW51OAEt9TW+wDFZDsf
LP9gcFulbxpC87hqA4RZY6HKrA25OBazqD0uyRJ+7OBlJaDqyY8Fu8xfguZT
wHr+swLuh19pCqULwuoTZj39SZjMY8b8M5JUYOeskUhBjgFmETWpw1Y6pm09
PDumsnGT9UhSOfwyqGHo4+tYwaeCE2CSdcKrI8M35q/qpbSFV03tzae/1NQ4
x7DTllg1D4sxzibnXzsFS1IN77HSwtdpqPHDC4/dhaCDlxFGl1yJZ9rRIkW8
eOMLMg+DCzXEN/32qFEmOORQKWVp44lGNELjXgMLt5rMbwrqebmy2HyKjSd3
PByN+J/BS6rLLxboq/+P/8FG5kXgDO6ORY1H268zDtVe1SXxLv1RbkDQ4/IG
w0DCyrOLeYcc6jj1VBoKvQOb/uwNFy7cB5zkrVEOwtKgVAvFF/UTFYw8hzg0
oydyb9yB+U6M1Z9U+1rNDHnJfIdrCo1br7BIgGMUjD1DHZp9QEaTDvhIGrQh
mEXaUQMSeIoMW3EZv1CAKQ5I/JfP7hjzpcx1STcfn/kcp7fgz12grDUNVhtP
5uhEbIkSvNFFmt4WCKzplMxgke1+NmmYHbpCBwv79R3RbE6JuKCDC5RBBWi9
70xNe1lDQngbHyv9nTLuNM/vZJT0FZbcWxxe/teDkfTTS76w+vwcgaPmrQKl
gEIIqAsLF3ZVpu+nXQplVCXP1PxWFfqVmcNHiqQGzdgXpguWuiOUVf1OY2aB
dvZ0dD8Q90cz+6KpXiL5urdp4qzMgq5FmPj0Q+ynChpFVfL5yN9bgrMWHJJT
PzbM69hkv8ozkaVSdSFIr/O6ngTohmTUVjhbd4g0fXH/qe3rV2nrukQ7aA0X
y8WE5/9ADEBplrG1Gg9bLFX3uroxw38zN9H4CSh3GgMgoyU7P7+ntik5UCXf
1kEprCqLSasIgxtqlIsNhCXzZWiJq2q5KRiR8iFPrj5BjXRuvAWKTYsygdYV
ny/r7O3lvNxC6SO9LKd+lJbH/BR+x3HmgdlsMwjFdtaYbVBltbWjrXJMO+yq
PcPM9JRAlhTdCsTZydsCJR1BnHPT/Y/2G8tRgZ5rGp32OH87LNfV9EnRHoAh
hVfSOtysAohJfOOCPTNm3ktwAaqk65nM3q6+YOUu8j90kNjKp2TIirRQRmUZ
qX+YwEWjPjMPy0MSwVa/0GPVvv7QimLv2Ic95GYZzAl8IYUi+bAZWgsdr2Ni
p8yTWjZRL09RrgPJ/QqyzMnWc5JtIrOd4VK0wFgLXLWqRKYngmqSgJE+SElu
mZVBntWry8oG5dYNA+oRN6CocPnu1BmRyjAdRUyrxgVFUIXGowpeCahd5f3W
JgO2jbaWRnChE4hYZksd1owGDVE7Oe4M+mahC1jQJdt8uR6426rlFRe4kuqT
ZRkvwtsuCY9ymZaCmUHh+jNztprPs0wuNBJV8Cgr1OuEGvWWLERAttazaP+n
Cbbp5m+BSOYHpS0A1lp8fuZ+l6KBohLuB/JLeveMG2jtiXH3U4IEefRDniwt
fUasnxGJ/qOpWOkvihkwGZDR8D62LxrIxuCARNkKhnhyK2eU58jETSjh0WSA
+7QPJp5IT8MW1Mb7/+xod7l+WUDl90EaLQ1v6yVJCjZGnrl03NA5nleyJC5r
UJ9ysXhZy6GxDSfsLDIT1y9v/ktWsoS5zVhOvJ6R4AXvxQ9J5f0prk2spXLH
pDnnXzGrgUzz7FOqm+4yy6E2wvA2vOOBnThcAaOUY0vkkL/U2zGK6uW1IGmk
wNhkc0ammF+b1xI9OR1JiZg4iDX+fRaxGdVeRVfNnGvswywPCP6snUdKKt/g
cOC7x17VNy1JjuU0IgWaEv55Oco9r2nZU27KK/TXQ2gSjAwfBMpcei6e+E0D
jfLJj/ZzqHp6t+8IPSIgpedyXXoseiHeYNAb7NMVHNFgc+DkbrEDDfMkALBX
2Ahj4p+DshikgD/LSrfmKmrqzN60WXlP0OwRZkdosYU4rNKw/SL350eMyWBJ
bfX397BCaP0n+DVYwcatZoxTd5PLix3PsoaxZ5zv6Ld+6FTD1y96G4eRGnWg
WCzM5KZJBOnF61O6/CASPPnzb5t0Z7jubcTCzzWpWobI6iNeLHK16D243ur9
ejKI5DF11CXPDkkX8Rug+j3dfDpk63PQAt+p//5Z8HP3+XFY9rDFl5ddJ/Yl
x4Po79jOdh5TmwDU7xfkj0VYg13FxTFJJUDl3zOOxxnTV6tQ0XpB5unHbmlT
ZMzIvce7E5TSueQDo5SpslFiaNHDjXzGEcKoub6eXX37cyyOLXuzECEDAkd1
mwjtRVzARE4ai3cp31EZLjvqIBTpaztIVUKzRI3XuuU0drw3Xx9ZYnfLZ8NW
DCSiOH1SmeVD82B2n2TcsLSjDXQj2U3FyFgxwUPEoA7HCoHidn4g5XtfBd4M
QYSyhhsUraTq4vvO/MAlYvU15yGxXarVFIT5t45k/p6umn6BSPg9vPUERn02
O3umPTVOQrb07cUWxHlypR5vOYswAVz7q5S2pBtgjkt3tziIxRhwEDIOnqnF
Gjk65ya6OjxUutTu8CycJfSRhmzU++i5SpzZe28a9Scp6489x+C1SCX0iPDC
4vHz0uRyVR5BOK5QPT7PVqTb9dERdA1roc7mVdAxNWFvSakGWq6sBVjiGdl3
JwDDTLz9U1rFljPWxSe/VEUhg0izBvCMOpNh66rjisqLeA1jcPT6EAQrwYw2
NwOjpjon5Z3jSIlwp4r+EB8J57ioahGDdY5pl9LU0lYpOrwtccxEH1XanMZ5
0UH0tTAXyX4oQcx7GSU+hVSVB/m5d/13zlj3VHhkys9wZKJ+k5cbuG7t82Js
Ks+w00lsY9p5oV8okuUrklG9LpNcT+YSeVVBHGrTRhEeCztAc2MQPcVV8dyQ
Y8VBvw5J3/v3lBtp6H3VcZPalOXrtmP9qjQvNRBRD29xnOv0y5UsYShTpj7W
KJO2hYe8vLj1iRGbcDF4tg3e7oazi3gRE5KEV/p1mwRvonj+9Rap0ENfPxKY
BEJBwzER9XS5PiTbqjFWrav6ma8b4OxKozfV6TtwZNI++1tocq8F6I4bHPca
bVwxobO31sfTC31adMlo0xbxj/+Wh31I4Wh93rtrsRn6k6x/QUk2TUU/WLu9
ZjCqF4etZoKlGZEOGHuLRSN6PEWwy0aAei59HPzOHt2OvE2eB4ft6bUAnuA5
oDIjUUFP3QC3Pv56l2T/8T6RMXZKPBIckwWLygma88Gv91NHHdOyaQRShpgE
Sqr7OY00MxyUKnpi475EygPAPvYF/xKtU1O8BP6q/mnmLSnVsLLjWJiywmE0
jwtw0jPXFI41D6ZE+IfiKjGVhsNBklYtvfB2bfaOhtP5Q8Zz2vO/nLSWzKhQ
uekUOISMlpTWOvP9JeId+fybwpO8690Kt68mvBxgPgx/x1yU+9pu0FC6YZvF
NfHNH3fYiDDQcVUx43OJt5Hr6r7VE2lbPi6W3isidTGDJ6TxSOQIYPgXVjSD
sh7XrfEFSBl7gk8YjIqIYJLpvj6IOf0Csgeh6DZUAD2Txhp1mphbJxAs+oiP
nzw94WOqVqHd5ZYJ4dgUdChgWoSrlGU9r/U+GQaQV3MWozxyu2cQxXF0S7UD
Iy7jVlkDH5fOF9nwYSsEf4ziijYNqtdPZK7wnlHOVIIOmk9m6KyFlL7hAyhz
wPKPG3jAeE+P0S8gzEFvk8m7RtfYn5Ipk/S+zT1OzNjFXWr3N95dklISS/Hz
Q0JJKJxP/bH6dmNdOryH3LayxPeChY3KVEyvQBmm+TgfzDtABWwcfBfTzfgU
6INI4X16oy+YIpWdNbkOYDm9F5P9R4Ea8F71SGx6HLj3VlLAHtA15PBmaiEf
DFk3G0agMdOefjvVK559HYmhsbuRPvDU06utiwPoeT7LrkNP1RZfQGpiSRm8
NqA8Ebn3wga39iCX2edoHDS3/1KKVQCbCbM/DTANe4+oLarZGiY76Rza9kvr
LrE+qP/BIov+6FbDZFg+EommERuJZlkN2YKGDOhf5Vq9iggJzKadAcVTau/4
T5K5UIt9fqwKe9cJzAmrSmmSvsD7B4CYorG5iIWyafIgv/+9BvhVKXwOCJzV
ZsdnFGG3chfdsBVPnSqTbML1fuHhA4Xm6/Zt5LuhRqg9ZT3UEitw66JQ/obA
6aEjy2aDdX4D4Tc5lLX8g4RiNAKetgnxy1UbofC3cnnJY4UcSo3SIcqbfU5a
okoKoCvFSpKGC0tENE6GM7x8ubkqwGvLtpDOBThct4s1TnXq6/6ZZig8/qrN
LcKfTUgoOKtHdHaRyvV5coLNWrxA7v993kLjGlqWHEMQgT6Mzp7ZkQ7shX60
6MQcf+bs1Lbyp6D687evHoDddukVR5v7+0EyZ73X5UXV69f0RWdhU9gYIKPP
1B2U/7KTMDk/1qUIWwx0ILjSYr7fHnsrCo47zk6F7l/1il1r0iwoFUJUTdbb
mtnAGOQ8ZKCh6Z+h0JuYE/6S7Qtg9o8HE4fdMxjii2PJ76o4qgDf848xp7QV
z6hAUcswS/1w38eYZPEGJ5Kpdb36GrXmqKONNQ8Vu7IqDTT41U87LFdCgJ/I
hRR2NZVMcT7fQEanwMAGBfODHH+wM4Aad52409pkXjLlbROokTJSeq56b1q3
BdVbbFEQneGD4Wgc9w6MYP54z1apV7m1LmhAQs1Tcg7R9X4Lk28NL2uisPOZ
ZDMUSGvYOZSfRPEMpR2JAfVFkDgAovhuLNfQFNjN6b43kS9nd4CCioshYgKU
S12u1MrWGaVknEgd2AgZUCcKszWutrNwgQa/CDz2W+8ZJNWqAYmjF1C/MMX9
3slzP6uQb8Hjo3ZrE4XQl74JVR8dLzxg2dEug7MXcC/10uM8z/BeKdZHk603
ALcfD+8HddCTn+Rbkh27kKILkK2MHpAGTtPCfWJ5sYaVjKJu1/gBbDUqWy2+
5wgi0OVe5hZd1uGHR6FNc0Jq3FCY2IjJ2IEzIe/6nAQxi+aqK2MqZ9i8PgXv
kEkfhnJjmYcc1adw82Z/P1gF4trr2oCDARGbn558e0dm33NjCBRIyrcgvvW/
NT1korxMaWs9C0oZwbe441bzPiWyA+vVg7BQAqkv3jili45dUtirKE/Srslw
sjeStL9q3+cGt31C5MEFcU9TjCc1cvhxDsJUHmQNWRfWSZ4ckQohtLq1waR6
PB0WmInw3YYNb+dbjoErlmYpxrc1CdQbrW3p/b8l78KQO4Z7Hs0dl7e4h808
YxMQKbDtX/xWqIle2M69PgnZ4HZkUu5DFj4khZoEAYovQNSdP8awdDHFGiJh
YIN2mpC5xLNUA9HWKx8a7IhlhBDd+Jm/9d5yE59RbfT3/RfEcq+Te0RoOHCG
XDlYGXF/DHPbw0/F8r5S0k5Ou0yItQp5vH9DW58A9nLkaPJQxZp7GbNBU29L
Yq4nAip8rMVTb0bafWmnYARGekvP916AHnGsxyZmkRRvu5Rhw8x7SZbP8qyO
VwnfRgI8NF300evBeGYo/GqRL54MXcAHTvZ+zot4BgU6Q+tyX1Xui8QIccOq
XwYGEbEG82yqUUWPeihK1iZX8qac6mDKbnvRxVBUCB2y7g1hmQanuWH+r7/N
p++0usEWhDkD5IyWYalT2B8N3tHdawrpvzITrxjNIx2sEWzF8hCvsP0dWPBL
RupIKwWgylGATK73D8QMTBD3dH9M2ds/Mj/aiw6UtfHvbE+vkXjUJUcb2Qqd
YdXElllYqrn5iR4drewzIjLmy3saY8MOQVf/S61iZtoFGIFOKZctKfFg9YKC
VmIZP5pmtztWtR1JdCErkoUCB73YzyaJNP7u3eNDqGtlgmBgySMoTICCUH4V
ggkqgFr03btQfcDmPkMV7lVaWywB6ASPiXGls8oh40gDpz9G8y9/m/Gfem10
FeKCjfF6uIIvwp1cq1KsJwQ5PqOFsvPCC4BgrdOon4W7S02Nj7/0VXYlJqBH
4pe3JVTRNvtaNlPsrOxICMyz9H5MVxTGOw+22DOcEr8BECVNUl9E/c5beWdJ
NQzTAARR5+hpAD+4Xj51IRaW5nLxyv52qw3wLAeWofkaTA762KikwHAfk/AU
Hiw0dQXqEmzkSRjaZQv3l1uR9sddAqrBf0MRyUMZXWXKPz3Gca9xIZqncel+
Ay5p+44O2TnWnvhWchftjTNx+G39quzJqomt4OE0S/3dE6BXwvo0QKFEgnN2
DC1PWt3BP6AGS/Hejn/p1x384ku/DiU7IX9/ZZWdTlTYZTT4LBCVSAQCykLG
VlL7hL9G/MDe3f91uAQ5hP4jlPhmwxOVgehrrEq3igs7QDeVTBmqLKEERUst
KXs+OOpFw0tw/RlyGIqX5/E13F4jH4DvkXLT4eULr25Kty6DIotlFfNqGCxv
oaAeIbC1iUBLqPMPdkfHokD2XyFDbN64z1VZ1r9y8PXCBexSfV0dyCxQsYFj
Am6AHrN6Vn88oGFl9GqZ66fagaUmg857l/FtCqYYBTJtdu8YcX1UDrX1Vp+f
NMugki43pOTn+3Y6wumy6GBMe2SIrejB/BXRHs9UOjoEpFFXF9QjHO/BbxoO
JkgAQEmAnk3a0iNxvnbKHXKB16ryAxNJ+p0PwdiM/W/dHvWZvFpciZa1Fx6G
JWJYDSMkY8rOXBvcmVW9Mj0/9lHmuJAOZ1Y8lghfRo8WTGEzoYl0CkaJSJ4l
rnCJKQbTJcqkigrBNkfrmd+Zpvb6RHXk1uLMKyXJIpnRTPbwDHiHM6wI3JsT
kzyB6VO2fjnvOlBzYJnsBMLQ9zeWO/SGFeLCIEvlC2bCcDM9rH0wKI4iKtDG
4vpGW5TfeiCd013fXMnyVDAwUz82T/Up29OGn+dqwJdRjO0TZGjYdWiCl5p8
vY4zZP8KjzvUyD/sl1xtqaRfNeFRMvIG5VSQYpgYppNUyu/P4j2Dv3hEb61g
Farm8JJoS1LXuXd2RJIgAkGmp8N4RXwzkAoF9BNFJ5lP7rq8eHiecJ2EWSib
7Y/vCIfadW2CMBJ5tocna3y1R5uRfasEmGDW3oTjb9VBlUBcUJt6LgZUlsGW
0MGc4OvCkYiWM36eYRp6OY3R3BQexh07+8jT1Kc5s6FH13XNgf01VoB+/mGy
Wvbk2T4RbdAgR/P7xJvMQBv9vcqLXDTJIslG+ZzZHF9JCmATKjkL+h06u/FM
1dZu6o1iaUZZllHWP+t/rqaQ9ENf65YX5EtVTn1LgIv+RbeluB7bSzVmJxwX
u3SUoS8AjGF31evs6Tsk+V28BzkDVzPkpNWKKlCJOaYof7HmnNiiEIirB9WZ
HzssknUrmMjPK+crJ/pZAtSRIhcTUq8WyZW8qLumb1vLnhJwu0dng+ABZkuP
wMDZlfeXVOmg45CpYTDAznVbNFBxTSADVdxv5tHN/MpbiLdC84Q3GQx3pRZ8
m1SPZixPRIC/vcWZXr9gcp32rs81f3mCEf6KgULGEoELb/scTIALlYxfSEum
SspFwvDf82RPAMh1JkU94mk4nZxkxjpJFPGIscsrg+hOHnxlaac841H4Hnak
ie/sRv4UYgV7/JmsFvZHgbc4kLvPoijM60dwfupWtb4Jsvs0IR2KKyRAcvuR
orbkKtBl8P3ThO3PI2t/k7q8EMGnlpxPCcMbzzgMkXDLEM+yEir+vOJmHqNM
KcdrcYGiLidU+mwxmkaNkH2/da63hWUoME6ww3L6ibkfFTUfezmBi268n/KE
pfhtLVk6iZ6b7OXil2l8EJjBqI9Vx6Cv87NZT1h1U17hhReYZ/jvaDq40mzn
j9sKGh9GQ2RzqYNyAZbRqxgMY9ftnYIslqYqHsaVbz/szZBDzYxTSnGghE5K
hyPASdAZAYwhlnM+J5ybjLXWk/LG/I9LWm/AuXeAasyLuWf5aqpblkWLhxoG
fCXMbtGbtBbDnVG+qceDAGcYVIel8yKuONcVAY/J8h62TQmKMUBzJpPdEXrG
luOU3Z+z61yggXQQWHH4To8v6a9uaRqAbdZfGRcpGeQMQOYVOcUu6D3wwFWL
6GnACF9/FbzPBehkfvh5zd0fp2yQ+MzdMNhdRDBiExXHcg3BpvPqPZp8MCWK
5dexwKqrYk1O5WfNMxSqP/jJtpgRsTsbmWxzINzE/TW8ZjIM58BLWrFWaZik
n4c2a3P8KgUE7rozvp7O4gqs1aWHuVLD+Y5auEKs14MCBbcpwcvM5CruUrjj
MxuVEDPJEhqOdt8H5bRJL+qMNPc+Apn496meQxOy65RHeTjP6B0/Nl/0vWvh
pv2MOYQPLWss/WyIH27kcXJGcrlNlPZI5TJFcnSwFfEPa3R9UdUThAr5nTjd
ODI0q78XS+faMQeOuTFM/wbgX+qcktsdRzKfkVcADlcx6Dz98o9UKXx3jCZl
5TBXEUDJUuTol8apfnblj4+uIiZerSm6jPhTMtZRp2VJWsynoS5wKG5vE/by
WtBhsvfvn9h9aik943faKXSfQsGAesfAp46Q4bNgXMqcIULPU94IKTzKTzZU
FtpJ0BH65J5xkgr2O0tcuNGhcJrfP2qF/BZByx9INo0VEeojtAAto/cjjFOg
zi4KNqoN/FMdTGWihI6m+WOGMIZ7SU/1/eb89UcMPjypoDyPB24S0+kXHp1u
t7k2viC149RDUwEbHxbu8Ag/hLJyeCbwQryp3rtV0TqEvF92hZfEzlCVxjWA
VulE1C4miIzHUGN/0rGSs5n66XP/Pl7KS2+p3JnGs7+9yOMjAyKrEL7LKYK/
79dLiHOnTEvL2UCPr8EmCeH/vFCNUoaLHsXJ6C3Ph3X9L9ngDHZ6mTw1SuFR
0Svp5hR/Z1kt9tayIzw2Pe1OOcpnAwlBc33+dCGsuO/E4FsbeiYMjHzch3va
qjncxRJhwzs5jraHismJ85bVnTk+yhc33WQH+OKfa0BKIkJjyl05TbttdLTj
NSpK+WZNcsDnrp3nItVu5BsFqef/Sa7oZoPCG/iIQvNF8tIC6u7vvk+zuU68
8W9PNeQN5vc7MPtI6QKTkCLavUPqaRbFuEiBashA/+3B4QYx4Q1o3Ip9TE/E
JSgW+FcmUQrYJoaXLyMyQIasMNCnWUwHrpC8yEj04Eo9UxLc0GBvlUxCtieY
pv5pbyeERLfj+DjqgCcalzfT64vjA07Hgpduirv8GZhbHXXDCLkVa/vv1Tab
5hR/MqlZX79CBcTcO1DK45P5ho0hUh64264PP/IxvN4kN0o9kmP7geP6goMF
qc835utc2gVnM/fzwV9drbGkluy143zoIvBQ92mUSbMuUtmLO8Yn+m8YaCb7
QGWzYBKBpXcHnYKrInRhV/Drd/bUAlSxEbOfEriQvWJSIIt7NBrm+/x2PQbn
Q+Gp38417D9uEDv+WOtltHJYl5JPc9h7pcFWQu0lBTTTbnhAtvIWXFG+6Y4Y
eiiBbw5SoE00FeYUxpNelHyye3dDZoqCcbfDwGeXWuqc3i33Uq5ykPgQ4/Oi
AFpFUegKyWu7c08HPCplqWz3pUgaDi87TkCCys4+yfspnWFvZKHn6SnDC4+z
qwvPAplgv9z91OQJLTf944btvpzTfyL125/MjaEtd8uyJxGGB8cyVLKhh4ps
0cGS2kwDum5e0R0IBATYdo+rOZmIjiMDJ7ucCg+ChkDa8QcL95KIc0+jihpG
f9eacn0bG5NzSsb3jANodBt42+3vYaHmoQFuJYnBLyx8dQo+Ami2J8LB/jHJ
B0LTAW/U3OKYTMZnbdngK1zZNC3o3JZNcyvCC046VekHcPEOQ1UEIS1G2yS+
4sYqaRYgSjGht5MXohwaiWeKZwS4sqp3IsLtzla64tmPBNVHf8RID05x4k6x
I8OmyGn6FQx7P18f1QXkKbbLoH/yD+mnRzpV3rYRzUVaXvDj4pgohFKgTE41
1yVWpC+0fE5UbMlHwAIPUREF1KGnhpioqjct6gVF0IVoHpdZziqTVp3qcwqF
2zU8pdxiwtmvOvYqRk0aC/K6MbjmEXw+2hKAIfnSlmhQIIDKcHeDla8tQoBb
/qMe83uSnDdqm/N9AE4UbdF2l3FS7i5nLs5Jrlhe3PlkAooVoiJeZxcdZybg
F5yz8F84LvYcUEeqdsRkwC/ET0L+Hs1KRy854WX4bd9r0+IRMaNsml0HRJtk
bU//7hSBeGhD1x9mOjTVIqAawF8g2iVewAtVHEqXmrSxOEu4n9ysVBhurUUh
UboXtjUoUDWV1kpcHa+pG6l+/nQaZPFWBMoRwqrYr4Dw/xMcFuBMqAmtYy1X
IGYuk2t50fetFOfi1y0vJ9jqxgwMB4/dfNeUzqU8mNQvNWXNSvFy/2FkOpq5
9Mld/dahssLF+UcmQovBywPdzgeN+Uw9sE8giaXp/J2ypOLdU4vv6Cegb3Lg
alJypXVVdWyJ+Spppkid9/BropF+MC6omDuq06/P2fvaboqAFUY4Z8gzjWbY
SiQxPm+Py8n3fGd/F/veNaWgagWRGM1Ia/hmgZG701PcOhi0h19amcl2+GlD
vDP7QDtOzWA5dVwSxQzvpGUlBpsEtApW1u6867+AifQiQXXr/CtrbsZ5oGmm
8uYnkdOuX2y0/aTF9HSLhN3WlHHzzl4KlYv3y/vLwOs8Ow88eSNv9ME15qAl
Yj7olaVKj3UKiu8GRiSAWe6Gzdh7QmURwxT1Rw9NMIT161DQOooDUCKezdeK
4yJDXLebFm9wtPOTmypwGpXA+1dngp+/URsK8bW6I2+AU4wpquMy+udnS0cP
yQSQXOlCR7gW0jeZ9IGs7dqlmEFHS3g0Crst/K6I57dAocs/hma+DWyzrWBh
VbQMQopVJPCrNx+gotG6zO3LQE0m1WIuibhGfNsf2Wlq4XHIBZW0nZ+UlJ/y
DdJiZSHHic/GTNveMdlzBvYOmMAeqV973nGJezTtjUi/obu7+nEPtQ8pLJpq
/6bM19DtQIvRmOaftXVkvfKiw2nLevtlp4L2IZfUh0X+LJ9ReeC9bWQnwXQh
XMLivYiSKwEowcUbfNXRE2dURWkQUfbCl4hMNtAQaTWLjIzxOEUdoJZbHpSq
uc5YaeMaa+tT/7f2nB+R69C3cezS5QGjD6EQ00X7J34MGnkNj8oO5l6BjEsP
27GCkBkSoo+azw9lE+esdD8RZ82h+xixb06rMbQzHo7DLkjpvMQt2453Mm+i
atMVFwYGG4faUAotX5g2QzTdJLVLoEZ+WN+tuwx1EYR3XSWEqvrS6qSknLcb
RGDlm82Gcvs2wZDbOsemN3yhFJAfFcZ0Oo7PgVs01RqfQfiEtOrrVKh6j2e7
Zd7GiFMfR5iNviWDLD4SnRDbLuj64TgIa6XTfI5P+CTJep+pGbgWEWAALcWC
lwIEdFJd1gKCKvGY+QR4AP4A5bEmOIkpgNYBz8K0CwQbJX/HMtHxGk7wb4iD
4RTDssbzTeliiUCrJ6oHhrGfn1x+HK0RWj5dUCCPhJ2plag9tBna6kD+N73q
tvoLLizqLgnYRqoX+ZfBB/1oJd9S0VK7WYSJc6IYd7zKKiuAaiKXMqQKeZSI
s7XGWfQj2dT8Ex38Ie7wHuJwfcLLad6C4tzF+6RGJYw2Xdu46hiqKqcZIDk1
OqdH9zcrhOjiJxuDq3/YvmmtyDgqI29zFSYZDB8puQMCOj7o508/mbjvVeG7
gDPOaJBp7PyKXaw3YRuiNQM9DHYcB+ru8VRnkZfDzifoOYkU1b/MqjXlhY6U
3pQPXauFV4I1P1tYPDXpeoMO8Jn/EH6AJPdAlJ5EruD2VEwusYujOw/DtecK
hEko/Oe/PWNGXP4MudmFbVvaIf7gSMSP8P5cW8BHC7gVDRLvYkocywab2PcJ
hCAZZorrrVeUKXNNnWiETH0s6Rj8skes31wKDgv9g81L4r6AG1sgt0l+ywbc
D49YxGFPmD8EGnliTyBWWIG4qZSFSZAaDpXoXw8nnEKGUN4Lbl4i/6GeWmI2
2boy1Y2tIlRTSaFXcog3SkuAhL3pezbh1tpZk8JJCKUj7kpYNsViRsamPqIq
GCE6ooRRw76nLjOScVrQPtxBbY+LcDCaxRYEleclA5kXaPmtsLa9bMgj6zZd
y9QalCUdZD8cbpwF3EqDUJNCf9Pr7XEwYODifMnonQNccPf+Q1Y9HjZxYAnT
l9sZfZ0+mxOho8dERDp40rWMF9Ryd/GVNwc0V8ymePOg2lfB1m2Hg7fl/DmD
mbb77+eUiIz7ezgUGS/DuoyBiug2GnPnfPXdfa9D0+Ez9McJ1ROm+CKAVriA
AwdqRe4bwGYtB4EYdi1Adk1Hy36dyD6/r/o4hUhN7ukXT7BsJ0JmC82qCLUY
nJ++1nUjxitOrc4SE3WtFX44GlaitFpmg2tUErClk52CN4boxEqYan5CR/AF
vaEeDGGcO+DyptaeaI82t3g1GRKX8YThcfmnNvnNmPrIGu+qANryDWC3JkKC
/hy2Inc/1YxbD9GxPZHcRmPD19Cvj9+6wy0vuzce//GlFtoaZ9UvjMffXYXG
YXygCXyUl1j3YsR4Kq3PS3FNk/HuPzSQlZV6x+bAwrcaADVBi7F+3NnccBN9
Uu5A/y5+nladHnVN6mNllAwRYjgoZd4nWW7StREpjz6V8fnBICYwC84TI7WT
H5r4ClspLs+9Ek8y9w2BP8cQ8W6srZ8CR29WIuHkNONeN9E1Tkbvi269gCU3
ovjoVik3ovYIPFGSZNGptwWUGMAW9YanMPBq1YlpoBIb32BnNzSsHn3h8c77
zibddQy0H5YMnO4s6sPqXn6d87Wrh2EoM1CBUnY5gyy42/D88Z5LM8PbON57
5C4HhvLyuxJSTNOuOBmzFYWKkH3vsQ20BAm4No2cI+uK3a/sEHCHYw9Nmtpt
O+XXphxb1K9CvgKEsjy74HLWtXuGazU7LDJGca3+Ni2TjVCZbOIE8uTQmBB2
4YGaJMRm1MYx4sjHlwjs7UeW8HKBl0XgJbOY6q8/zZ4LjzGQjzZfIS/2KCzY
Ie/B4gX4XaBsURIuWxb0UkAhQ/mYRDe+iT3UEsOw2BXZvF+4kaNMWmgWxbKI
ZWrNE2DNu8TlgoLXKutO/rcNIZvM1fQ7lc7yqMLtPC2tP9ajKOK7vKKQjinD
UxHvaPFy/Eqx9tqtNv93MQPuNPGl/CRjW3ujxCOYrsHv8lKqq8G+HfdsvtVo
x4YR0FJ4FAkl9OCYC/mUVJtCiA6vQ37BnzuHqJkppGpt9apls+RRqTTEv+DS
wlijpTdNCl5Q7nmefkgLIcqRUSGSuOmQkXfTz5aOrWJ9Bb+0QMFsWegPdLh1
gYOJuDrN8nLrnAXB5PcC1oeAbeEM/L4pEsCuKAIMrkFrs8oKlqC8+dVEDqlw
qT+U2ySLFFcaDW3hCZEX7HYKYtGTfJ4WjbkJ+r2DHHcDozTVxKm4yU8tdLIW
3BhuRxWSWWS26LrIqda+MKHcKuOqWgvwRIVIX/9rz6YUvjyA3ERKV5YBd2Wd
4ekslz/bWYgrYF/xBYsjlyoaXeZwaLzEFFcxxPRT+4T2kuzuNeAigSJ9+3+B
mPEJM1TPxGeS3FoTz70eRwpMeJb//T83/TPI/mCP2u3RYkxfM7R9KRhotBjb
8mVXQYJCibqL2G4BJbNE1qenzFqLXYxf3OhUyOWiyeKocYBJJFnvxmCzkpuP
U5qi2dYehWD0LNJy2c4Z8KWZLu9PRfwcGe1siY8nChFERgJyUZkTLSxXTX9l
ZSBDwUafAIA9/g8dBpxrA6PPxbOzdUl5NLKE1hJgs6Pnv/4eq3oZMAnq8G/M
4tAxgekSCQVdtY0ufUALxy2hxeGaeURrZZMqt9aHinz9ctMLjdTVqPy+broN
o+yyAsX/pfMu1I434+0B1APGZkUj2fyn+G0IbWdDml54ik10KxGA9Zzc+UNP
NH/H5C05xygNspy6+Y86eRub7gy/FyBUwhzTKrZpRAGb1XysjORsLr/cougC
xuocymc+IVDPzrFTiYFR3fBtNLYenj0eBmyHD2/7t7RBO2/GdKPLDoCidkBe
WAmdqdDE2+XCJkahhDPr0UpQ1wcw+T01YOjsxaUzM1Fc2ATmDJM72GYyyH1h
APlgL1s8c0PxYDGZhc33aBZeEEruwTA3GnBBLmD3EEJIkEuBPIYmOs1WdstY
g7apdhuBcQxAbek1mD79QkjqiAKEtiL3/OORN+BhotD4aw9RGine8niY/mUO
v8vPg1Ff7t2BFjhFmsRzZein4gpJLGYFUXJOv2DbI0IBpM9tBMWETB7CbGUp
MhMD5XjUQvumB86M2rOfNKr+3nRr17gqsaimWO9U5siMkmzd8iyIlY49rnNj
x0grAnM/Ug8q8j4qlmQq8uUXKIEadSJ6FYeJWiLy1IFJaxmLlRO0TqSxoPVi
/7vjk/UvUAxBEPw3X0FiFzFqAfUiKcZqf41VEq9EUfwgwRokn1R3ArEIU55A
zKwfGfdaXoq9y7fUesPYfKJeAQytK2iI7cau+N74bthOThP8PTlhvNyN2bKS
q5MKsi/a9nFDm2iD++uZWR05/VJO4o0JURraejfH1easJFgZRHs4Giin8p8P
lOZcnIRokIg+fENr1DfsRyohVgyZ+ifQ/uHZyxWRvTZl2JuPWoBE5xAC3NRR
I72nHWQX/C7su96X1w/q/1dYWtCru2QlqdxgGYgdVbvfxLQdkKUY/BFweoQP
MIt1ie0O3ni2AoEHsU/KOmwGAeWJfQ/6yTbTff3+v8zw9n46xC8KaHMxHyZz
9BlMt0a+w2KPlC65+CXK/SWFvZY8DnYY2QF33qDaz3xyQDpX2bXqBVChin9O
6Lk6i0k821p8Z4qKcOhLZQ9IbvpP4hQdTxkXESAwDzCgPfdpk+bNXgoRaAk0
Voj/KFAyqpQNXTGlm1bylMj88tdsjPG7eSboXru/KhBy24z+uWqz28y7FHQh
tvtXZiTCR4rAIz3Y5Ys8+a7YqOI6LwqiojE1mz/GVMaae5YImVI3Ire8Ufnb
f+39EZMZ9f388Gmq7KQLvfJdqVFIRswm4EjGFVW9O/uR6KJykLKFMmJv3bqd
CJckMvCRU9jBQKqEz8kQ0Y2/QB/KyBdYJ0XGWNWeRnZ1YEF7hOh493exy7eu
rIT5UnJDV96BRI7ZkHCZz5oSzlWaOFAp7s1DfUWUrF96AiU4/YoqU8GP/vX/
PC7V3HJyPTh9HNMynKWmQJQ3w/moOUiguxKoqDC5crhUJRdg3eQFAdpYwBaI
SnOJJRWsdG/rEzbHDjyXSsgb08xqxdOD1yAwETCcPs6y9hT86FDSNjsD8zla
D0Olj0hhNSc/SmBVr4cYoQIEc9VjI62nv9r73qN8znyNltw6dkOWSgD9s5Ar
ZeXWuJO8lu/ZK/D1W3tXpJNbtLrh+SWxroOrcR91Gj3DWDdKWqFxmaaOpuv2
irzH8exAP1StBiJPDin261qYpzfqPKo7gszEQYKTC7VarsU5SKxz8hjROGqM
8a3wwunlt/pWmPW31bqNHqzzft+BT9lIqKzGTQMFsbg9YmAT9xiednYHAQPh
nwiPdXg7AY9CvAWqCsrwsV50eZlf6XqEWPepXBdOVF73Zfa6eTdlZJdfW5tf
8CvXT62NpPa3lQi/o73hH7v3H5c4DFgE0TsZhDqb7p3Qjh4pnzZxIYZq9h0f
TjT6xFxq6AFizZHhqaHmqTSOPstu8fWf7JlU9TOl13ydSfqTH6eNNBP+aZ/6
BanrZqjowynOsxHdfml9AmCySUAtJYzLWScRR0SkMid2iZzltDntgX7POZP7
kkocGO5d4JnRAfDdJ477UpGmXn9MWxkxMy2w9lCX1v9OgdyM7JVRrLXa1TcS
VSzMjyJyVxztP53caFJLG2/cSaP5GJKWJfVpCrSdUHDuZRrdtSn72VbF/DNP
dI5rR1Y4wYuNah9qgvf+O+LelzqApK+zDRMSjbP7rRDvHHS9Z/l375+tkcaE
uL3mSpc89dYBby2lUSL7GMrz3ze/8cE8BSWkZ9tqwxN1Q2dQl7rETUrOjDl3
jIWWZb+eUD1dBLNCAtn+NtR0HlUYlC/yjl/w5ekAcesPwCju06ghpiAYxGNt
3MKFjHjfIvpAEH+ZOBK3tH0gd0bvchyzAZ3nx57q4c8e03WMPKyHWTBPn6MR
GnSPMdIOin9CfSzlnQ6FYUxKtInh0VgQO/B3LWlQc9m/Jc0As0Svk7yoGnw9
8LVLeIu0DA9c2iqfUDAdcfAlSQVnvagqH4X6BIVWv9FPF3DpUjxB4W8hRTfV
3VD/p//+I/I+rxAeyf+T9BIHTqua+R/tlQWLDCZiocDb+aKU/Jjb8Dptc2ME
sRcBo9g27lcHlx9D9hIUknvZdKnpujQgItJFl0w5n6LfjmA09ToSoGtfcc5N
K7psg89AgyqJopZHzr2vug5u77+2yIXaJJE9MQ72Te9tvEuuaMPWMuGsvhwT
DYxLEVvEFO+8Hv+GOQ9yYYZHfFK5aBm1LKdtQRVzHz44lKdKS4izPuoaCBX1
ROnYQLuOCqLRInobXmYUxWB9lI2kWI6Ksd5cnY/zF7vnrxoBl3BX8Q8u/q8H
h9vHDF7QW8W7xncO+Y7HclFthakiaQ/XTtimL8ClBkpTuH6X0L1Bi+N5UlPw
lG+3FEpUnABlFmkn5ZV/GHUdlu999WjbY5sqaxMd85+xrEldUDTayzKaPiSf
3HHsKw76gWN5DkelE/SSU0AwL+gxfHAgCEuXqTN1VW+5MHM8ZhJFZi1QJT1/
Easw+DZVriv384BWEM3EGqe/KofygoQkqir7DBmKVWP9Lrf56RRs8z+8T7ua
/2PRJ54okjqpeR2kYVasWpE5BUgLjVz+8oU9nCxeCkTGfSnpkvhtnlQlW863
VQYipjmwe1ADbkK3akynFztyyXUd7bEdmdVJuRCq0rQGJhqZHP0c0KYv7JB1
HARxyqtxJeR9vqDlCiCXQEGR3LuK6A9UIPvOhOthjUKr7HHZLuFNDt9wxLN8
1m4gRjncYcIF2DTh8V2shduAVP72vet6h35mJaXqZN+aM3PUWQo+uugM3yqV
hEJgoSOxQlXc8eS9kNPXW6JeJ1pV89esE3Vx4BLyMM5FI60JE/fhWC31s6eW
dvkwoF0BcKcj3ctowy9jZkt6osIGUmn866nOiss4jlH0GthTTwdPkP5UGeg5
DOpOtqJ3rvk2VyID522bOl3prYtve0xy25cr229I0MujYjcRa8nfaipOp66k
klzKXx13AsgR1+ryQA6c6ULg1diTuJDZemHfOwpyiCcB1+0pgSPEAx7MAZyv
ZClVIlgliYudLI2Jmj43OkbdwOxCzEMpcffJ+lACA1f7XaiV9noNr0gjO82f
YN7NYny5wTUiUsivsXJHHfd7YECi2CKYYvDzGD8cFNEGNtL9pD38HHWPZSDA
wxXqtc+xqN74sPfEe5Fi3SbhbubBuB1ok1a87mn3wkme3WZslKD2QT9zDwi4
xLuwsTfK0hDbkaJgLFfLY/YGoDjfpe5vYCbXZSKm36ubDwjUsV3yo5hMaUGh
WncA90vRpUyuNWkh5OCeFPEOy7HPgqTLjAJ1+0bhA9GFoXj89s1LEzOWDMRm
DpXGDE66ohuSvcChtl1ENm2/6h+eoZIuzvLMCurs2g8571ZjhHT19V3yWwxI
V4GL4VUD7WVWwZPG8Cvy9ylbN5sU0AcLc+ed+y5b++kJsnpTWNgsmJfKprhq
+mEAN1CyBsX87+7zeKV3W+3vNnz4EBaDJR3gdTmxEJgLwXn/6ZeXNug1mRl8
rORCKBs+8A13eIPq+uLCHAupvmTg0Xhh3wjSZXvAzDsAw/3ODKTFBmxWVKK4
XdPpSNzX1Estf7QV7Zryxs8zoScueR1dZsmNYJcWcIdB5u3LVFSt5C8ZchmY
z9U/jPRSvH/n2CdkTKBBLKKYXxuScWAqIT2Gpl/OyUYAD6tA3ie3uFCCxHo3
b6DWIopYob1OW4Z1nsLIzh5Dfc2zHtZ6fl4K3evq5QWzvFfYOdBRiI97bjk2
t0WuMYPqGOB04mdMGNmGCBkwtu+V+WfjjBMOMrLgLii96iT4CKhJOub3A+SZ
gFTcl6CxxZt0C6MzaZCNLbxqUAxvaUwE4B4rjW6GHccFz98BH4TNyRYYKdAw
SI9IMPy+u/eGI3e3z9cwUR/B7lN8Euh0qWdEvtOOJ0d1vEWGQ8OTu3tvDiBz
8XnDWtILP8v5k3UZUhw9rKsn+YBWq+wfN9FFJkL23JRhG59uVMQwZiX+VGWn
TYwbjIUqsfA8RlNUpdPLKFPQTkRlqAUuqzeqQn93MIpVEo6sym0o/TBitYdf
K5XwkhyG0K0Y1f0WrP+7z4nTkn5P32I4pfJUiuosTKSpxJeTeL1PqavVlkWx
h9iZ2pFutNHxxuHwrgBdIW/NC18Y6CBq3VisOAKgiXI8A2LEJyAPCwT5ibhy
dbxr7dgYvtS0z+MkA5BTbyd2jf72zY2Mae6GhSMETfgB6eZuFdi/eJrA1R4F
md7PY0RutoiCFvyfFBRmQYk0wyKpzYf1vs0kswj4/NXKPH8JEzU8Ypw7NQer
OY6Yr73KAV4UcKvuxuEoh8xSJb4H59rBjJnjozKopTY7EBtkyrgucabayUja
wddQP2e7uRdbvaB9ypwCAeihDgbbMgyvxWr1wpwdciqPtmnYZAZaCmXETKah
iKPyuvdOF2pVVlvAATBsE1T0IkaqfGJaG+IfMMf0QTbwghzTUKlldMLCRDuH
31nZ4GLuz13VnfRchd4UJtA9+/KohMSL4HeQ5/mfxctBZETJdXq8W+sEPJ2f
oou0pZHkYsVSID1RDFyebYNBBVQnk5MPbJgS4GpsAPdEf8BZzbMMrcFVEPZa
leBHIMNBnmX7de0QGi4qtTIrGLj+7a9ahJWoQQnGCspLin9X//JE044TDsuE
zEujistIgzdJJGN4SLalBRlpI12Z+Kx7cQlAwrG0Xn58v26FTCGZJSkZ172L
97SPW01YNJF/tekvNhcHQ6AUn8vwRHC3pDnQtFLfVsvGuxVgyM18seD8CaKi
SQefxBsMFgCM8X9STlsmxsSp64EvEXzPfWV8xNgkOQkvPjNXn2TkxViKFPKJ
SIb/6e65pSbNW1Xlopl5caYismnylq1RbFfdKsrAFGfKBR+LuKaRPOBMGvj9
Cmn8OWy7U5Rf5bhZ4ORpy3yIYVOuNijGtG+G4ppkIRRf8BJkM2JRfWOrbZgH
eS0vRf065fgbhC5Hu22gp9v/v86YZ/eOvxjY/XB8Oel153VGpw31WbYxBck4
pqiVWB4YYtTdf4F6QWLPuzCl+DkTLc6Ztl1Ix+EVmx7ewnV+9qCTuVWMsCfM
TG0JPCEYlAHXVCBW0NK8iSRwVTkooE6QSLvKV65fcBFoFjNjZFU0r0sCoBHp
k8K5ImrIrXIx6rd9D1yfLO0wcJSuZYC/thAlUzoMS7rNPbFyFbylRiirKMIZ
0D2ZIXrvCuIDhd0GhULvsiSqFY3hPWo0JdX+ixG6EP6YQ5YWhZzJkwHAlg30
oq6NW64eFznCyJgpO8jQoGr0wBhXLRx8zV0JrpIh3iDpN9nvejtcUad5B5BT
0FG/G5Py7SHdFi7wUgxi4gUDZNz/R7fDKYKU9sXI8cy7mRoDEAA5fijwaitu
BYh098CyCjgYC21OS52nN+MVSVHflxPBKYJ60Yx4I36RaJ2YrhOsWDehaL+P
xylb5ClykGcKBQ5ToS2gN0BmRaZX1hYi9NNBmvDEp4CqQ3LqZW2yxmt2+E6Q
BGOwL/G2cNAva9K8htUHRAEzMStRRAsm/rwry1fjeE6DMvbo5WbIg3vfNCw4
8bBhtA8QeXM/VHZmrOEXaB+MvvTlGCpzypf+qwUdyKHHKegZ2kcAcQ6i3Yt9
dgxjhrGKu1XYjh2B8s+xK09flP/faWON1OPScZV+gIb5sYoWS1SO8+WzL+tp
rkUnKZmRBCw/BK1kjs8OSjpFTrv0Lt1aDUl9lrldlJwTtDFZK1tcnXfcRK2s
DfAb/yLnsrVv6zU4aMBav5ZetgUfIeP2l96DFyFtpen/elWmcRZ177QxJJ1d
ecm5zZ/TYA1/kIZLb5eo8Y8XaW6NKQ6WWCMstQXTjSS/bDdYpfmvCI5PHi4w
53M1CiHytEvPVxxr4PMbp+v0yHn0buIJqpKa4GSzD6bOx6aRySYWZuCQggTs
bvvBzmr70uE+bmybzV5dd1+HJPMQEDfsqPbNJU9rTpLXOBfhwnTo6dxUi7Bo
zEkVXnHjC7pLZuVHFGjCtXPEblv4Lym9liktmYby9BkjuSgy9tJv2ohIlT/i
UZknqRvCFdw6fVyyCUWHN2bLYMNfSvfl86JtDqKTqC1M2Yc205quaVfSJokB
9/o3Za0iOPAEtUB90KgSnyIlWGDEekqDAdIYf8246y48hg6XMw8E41amjDh1
vjWE5zHhtSRk6vXeKWz7wNPPtF6EHoaOfRi7eOakoSb8YN0GLpioAEflcdcS
T+y5La6re0n2FWF23ffPsY6IHXWy7B13x6x1VRbMhrrXuuCszwg/m/SIPBrX
IrrmTfMvOjSVJrxz/ijsGI3R5nt3J5RC7e2uuV4u9h/ZQ2W5kYarbEO4PabD
gPEcgBkCdBYJqGm2+7nyyhO247jp+5gt2gY3APDKfGSeRJV9vCJrVSntxh2l
6bW6WtY4koM7YVBnwx+oA8aOcI3Rq7HXJdBht3hm0a19DQDA1GWlk6UInroc
FLMhxOB3xl/ARkut+7BAw2djowKWFXoxHrXyikBirdNlhFp7IuWUt9b7J+Hr
y9IzQdmX5qNqH9RJzpaz22C1QKGHgxLl70SfdKTL7FO+nmS5CGBsuvOPHEBc
AS1iRj3IBXz+2wNE45QD9x+p4ibZ5FX7Ek583/7s79gKxCGkTCaxaPlnaysX
qFR2bBt9KL82zlppEBGVKd0lx9n1i3h+KjTZ1SspPjY+JcIXUXkBrlYtTl+Q
8gRVsaBu6KRHKfFWQm+N9DIGKTz3AKVr+o1KkTIRa0BE3OqMPCvNMAtV3dOJ
hCFkhNTC/sdAF3i0fgEZSBSkey/mwHiAdh3tZEm3D6norqKR4Y6IzRUQA+JB
8CWC0ULNHXj53MUHnJa7Zgdf/4/6Qiqi5aYHQUcHySY955juZhE5cz3Qoo2I
1qVLMyGf8WQWMpCU7D6MDYd7ZBer1TG+XzlQeMkCPEkc4FcJbeZ+mU0m1ZHD
C7+Ybsg3ItZpVE2J7Oz1cgE1XM1lvjx5EWf7XMwEffTHlOhrMmoFdomJI3as
Gb0skyrOnzufWcY39bPmTlOTLRbFtRX+YmssxK/RwEMoJaFG2B9qNzBDFWWG
wJ+1VYlCP9QafTyo5pBI7xOY+4trnnRPcXq1lkjmJIv2QpA4nOMPQ3ErQcBi
PArlXzXQtrNLlfBb4KYO79b6V7c3PEouOXI6KaCFIrej2BiooTCAq3lbjdx9
7cG4LI/L2roF5RPCukno1I7JjAcSsD7X+va3dtHc6YgpIrlrTp9y28ic0oIu
+YRzj6icFFdYVK53LrIhSVpmkqYJN8XP+MLAfzMFAEykSF0QpkYmT+yD8EeZ
BuEzTURRaN5EOteKtR6y3UzUheg7l3bWHQKlUiiNKZjvCSN4ApkypT3Me8ML
jAo2zMJbkRCWMbiqtOiz8eh9znOcvKQfLzMX5Mp4g4wMtafbuUPU8xZ/+7ty
GSYMabIVyIdqbo1WjpkKCHV1swEGTJTrciFJXPoy6Eo6Bj3EIsQQn1+wNqHm
aOPhL33tKBzFKzIRPdYjWSgfm6h53nNFATuxHSTktuS9Jcu+TmD8bLSQbqTK
Z/P6GwlOzTVKpF4Inj6XMnqXqHR1ZSbS7TmDrHqpMRhVegH8VUr37Tmy6qUt
XlHlbhtJmoX1BqZ2x6KJ8Q7o+Oi1A412P/OHJqd7bifzJQjUzGNNKZINbbld
E4r0DxnqF5PlVHdE6HFauA9mWOaT6dkS7uLzfEYVti7dYLve5nsX5z6CWKWa
/OZIqw8lV39iDgIw6wD5ple3LpFJMPM80xYg6aYVqbc57z8L5EoPmGTyu4hp
tS04n8Geld9Yd+Nqn4O/qWPCRzcWNuiqItEt6v3QGXvg4my9vkKbGLG6onPB
3RzHKZS8SpVmkfLc9tOpfIqbzWQexn74jdUt7I0VudYDs7f73KDsQ2XtXNGU
ZGzoE4c8jwWg++EC9I+J2WuT8bpxfb21g4hYJkSwQ0a5lPhS0RMRuDC0vGwE
Fkq37ehvUoo9cn2VpkfAxkTdCV35k2JQVvWSO8NXiiMI9fG5wdTYVgRZ+JJw
MVnLkaJLGIrKHEVaF3aejUtZLQo0LIw9wMiqAGvozuOwMY4pdKiABL4zhVTk
yrpotpd4KqvSXewnyZaUt5MQwav2vCn8L+Eqg6fXQ4SP1Vkshp/9yzxOyuP3
mNIAKIVtqKkw/2u+PfiTzXFV82oQzdM2yKHWTTWvzN1WBxn0s6YbS/+yb5Xm
UfIzoRqp+xIj58xPOE+CX0FfJnIarGEdEi3djJec21xoNKCFSWxN4x1Fi4OM
mis5k/oP5lIujH4fjYuhA4A4qxt/VA4HrynCJjbz0SEdfDDBbB2FhbOsPVMF
fwuBM++G+uK8pJ79NqWZ2IpZK6Yk/6ahxSJ0Bflpy+wei0MAXvUmYs7IWLc7
q6SdDOFydfXwDgSNYX9xeNOwssEaA7AaoLKxb5BTPVVM7RL/wxheHldkp2Dy
faGlyJihNVT5o3THSePxS8i7vONGHVQ9v8guD6IUg+jf8bWpOxlpJf/ZUEsE
TkNcSeWbO6Y7W8ksSMEy7jn2XtaFJYeUz0nPv2z7k4Hqi7Vs8Zmcn1c7tD+w
XBhgSwhl8xLqdGfk/ruw/XIr6gENAS9hHdtr/hv1Rzf9h/4cUyyWVhyiRvYc
nc9p5IX+noTue9wa/AV6t4ldl0CXzX2svCE4FIYLL7RbkCqSzElE7OfZqTpG
A5Ldn6Q7Iz2ooscXQmyMY2ya6c/Jphu87md8XVTDAhbGOjoxC805mz1ZRUln
eNL3HdsB6N1IcSyJnOr5dtqMP+fpTbpihRrS4UWnumTywmgBLeVdVfSKD33a
o6fPXFipBu0kcw05YpwcYYe5+oJOxw0d9ci+LUwLuOh/LjM+sx4MK7shHek+
CWtKF3odsI5DWKWGBQ7YlUQwGJp+8YKhl+GhjW6mztlo4N12GytUkX6mllGH
3WUxoSUFg2Yp/E+xMXUlJVpi454vI8iahEWGmPaoyLCLco9RbHISCMvOLY8y
jpcdOStZO65WcGnMAlISKJYfCBAvtFkBLBxNUht/SsQ+bKTlk4PBazzJSsWM
QUraIob0ysRff7U5GwPM1CSQqWHCzjMK3mYDDRxSTjuW7jcxgoaqIuADcIZr
PYqnMXnopkrq9xxgwcSC2MwJCEPyf+ac8qlvH9BvTfRaJODGOYxFjP5kfa14
EZNHQYoWAHCQ1NAqWPJ+e1elM63Uu6QjehO36tHMA3V6S5wyXkAz6dqmEQXm
W06Ga1tEMyW6bqYluJsAjZcGffZkj0NmrEVFAC72QAZ6ZnKvetvy+6NwDwsO
hVaC41M2rGm7F+ehtH6LAT3GA3ZhwltRPmhd4O1QbHzX4Jr8RNYTTF+lSLE0
d2v/mt/+zuYZiK/eBGPnuxvcB/7MS27EKrGB4bTDc1fJJBFVIeXdHLpIpJou
JzM4ZMrCtVhTnJ4eNL5kB349CuQDhEhuoey7av73JWl5tdY9nkRkK+XpNa0X
Axxa9PW3g9MC6gDAVPHjynw4/YnVxvK0Dt41PgrlmBJ/NN3CNp7GsglnZrfa
hshray+/B+dwAujYrJLBExSEfjXU7qrpSp4S5TdpNNDhtZj+6FhyvvkOXM/N
Lk3yBhlSOEEKk9BqkbU/jV6bdZI4w8UaWfE+k4evh2SxGJvgP730ZouxbIQi
n/8D4nF/kLLjoHzJim8oIhVW6eukfv+9qJeReQZV/2MTd5PvNCyifr7+705p
rLt6ydGPh5UBSKO7LmGFnN6Mg7vOKFLfVkd/fZRrfe5LlmFQBeE7O3TSuiSo
ibkbXhWAI1m4WMTqmwy7TxeJgKmbKLSOqLl4q8v9T6rNp63m3Eyux+sUgmJc
ndsVjxs9V3KSjSRHlHvkmTTfbib0jriSYVq2XjdQWs1ka6gIElqZq7/JDAEF
iJJhJnmyt+ZlaQmY1bFY2DDP9idpqjPgzJDPBnltmUMiMNBeh26MegIr31zx
EUAVzT0+WIbln+BQn7zsPYJF55vI/9Z0MQYLXSwUZMIrOdnp48v1zT2cMndS
seGf7iic/4QOdQ9UoJy4CcWSZMsmFIQDSvp6Us/zZKIP4xAV3g/nXK57Ol5J
sJmpelLsiA7Gnr9hrA4kfDLU1r8a1e+G5Ep6q6ZL2iD880qjbW9vYEJyr90L
RmtvvDm/IwYSXorPG4GVkvJFczhbQv7F0CEqffoFo+3GImr0HNrEpDtuD6FX
TIzZ72UE0eFW+80+WjhoXzj5bMqIxJ2jnd7zJmGLvXGHMRHlaJJH8wFUjYSG
0ZCbabbUbtaxX1+CxzbWjir1Ra7PX4eN8u0HU4qNLxVEMJrYORtngHBEQn3U
wHjqjSwBniEs3Txsw/h2/6YvMEJ6nEvbhh02NAngTODKUob2ZoDyFYe8o7Vn
6EZCCGHrzCmnnQTyQ0szy+rLOhbJFHsQlsgG/PmtJ+Y/goZfuFtT0p8Si8WB
XsyRtu7VGxaxwsgNZOut/ibkmW+2k0AdOmEgdlJ7crjxJ1lFTmcTgXjhDb4F
G615lwD764ca6/HYAk15EWkeYxfvkEZOq0FyjwhZ0CdsyGySINEuGtMpoldl
K0Z+r3mWZvX8ZnmW0Zq+tNLvr6SXm2EzsEAvNhIshE+aqWtRZsg4UThMrhWz
wzSK1W/ZgP+SauXqaXCJek61FIcxmtip6HqiKGhnAOBvenYyjy2Uh4M39HIc
IxcCTvLPRc5UOpoWe4zCsSODlQ2ubzGbjKCh/RWbLKez8REhEixP4YTH/ykP
fLxHiRCyw/GUBGlYfuhK2m+eeUx8OCaAs9X03MWWQnVuM/t4XZAfpVScY0ns
JFq7w4wxylIx+2PK5mLaLYyWjyknx6qv+S+PAvPyOX7pwmYP87ou/BDryu57
b7KxB7W7KezianVnDaDy/LrL7/9mWUaAvnjUCLl+zElFNZ7ZSalsDOMBekHn
au/CPLAswOC2o4/MihCs0Fy8+3/O7b3FH76xSYWnx3w5YfswESGtFSbnJ0jD
qB0WyKSZ9WqVCV7JtE6dzY9O/mxnanTqN8NNwdKUoymQkiiBtCVlIbPbaFDD
dq//RG6kSm2O6mwNiuIgbQ6CVoUlhor2n+Ft6V3YFpKIcfRWpClOt75RE5rc
6v4cgkEHA6Zl648PW4cO9j5ZghkASYLYQjVhOzs79X1bMuuHPbdJN74FtnKQ
Fh6h7uIF+EyFUAHuGJHofLX8bAiKwXs6olzic7wc1UuDM4UT1xSzEMG0mqC/
qXnAwdH7fr3yd6eeoEkoC1iTOkt/eaVEzQGaRZrCz/BPdJyZkKHetru7Fsfr
qi1FM8IrNlKaGVYXa4LzcSyvXIVE3vgeGyOjyl3N3M3Rnlan0AWkXe/9N+Lr
RNjM+zVGv0oDStpP0axaPup95yIVhd++Q5bB4uv+cFFr3kS78tK0f/chR+/R
abTnBmH45etMRiKICLcIBG6pSlZiK7EvC6xZCgwbSw5SdR4hN4bN4fXlGG1u
4u5Vk8zHNS5NS6OKaT4k3u2GUsfKCBAJxCeHmFpfswqPbYNRVi4frvAyeseu
Z0tGt/+ST0pGFI8G7O1C9t8AwsZ/loPnOfKKZGJAJyG2SoNp5i5yNQjCUiQY
ZKerBT5F+jQNKwwNcmPwjNIfwnXwdDFbgHrCT73W7ewvh0xy4UZLMc0L7tlf
HSwx6JKTzaWvmVDcg/4QTBXc8B40dspHaOibCRz9Mb1L58LCMorjcZ0GXHSp
1VwDvrO3iiwmTsJ+YUwuLP1KZiCem6j5CkmssKQVab8regb2uKZ7ce5pmGJC
+G7RahQDBcK+SPHeS+F05qFqw1V9wYCpf/hFN/QXXqIHAHt6yiPZPG719asx
tMNf9wnIuuZmLvIiWa3NoIe4w+HqcmbtPtA2Eywc48T5YRg/42LTPZnguHRq
X/DuEuikBNh2CrA744vhx9OB/ZZ1L8NT/HDuuErD+vJtu2PA1zvnzog/79LN
qfzAUaNARve3J97iyMeRBIeMFl3HjQhPUJrUhTLmGVvycfXMmmO8c6brg43J
znVYtw7bRjqVOaJ9jo92+IQxBuLI/Lv3lB6mMJCE7axHwbyV+nXJOh+U9vN6
2hbOpx+Ru1/4I1TUdS2TTRCD4KVoDvLuK1N5m8i7ZT8TVdJOGsSORVAVgTbL
uqy2CQ7jQDn5TD0sNCS1uSTo2czgvDJ8nV8kDDYqWHnBO+Z+UBmH3yj3aalM
lmC377tI6UL2266eVqq+F71EoFBwuGxMKm6eNOWXVerX2hVQ02OA/bzWGS5f
oq3AhHbBjjvBtBzhrupa5Guf+ToqVLQJzbpNjuhPBCwOryNLHMtsLIuJhyZc
UUi8Za9vy8eTYEYKbsJ9zpZCo3J2Jwi077Y21xC1ckxsmFp8yA8O7CE6GJwj
Y5BxjrGCynR+5hpXf18ZmnP2je/nH/nWIwuIOa0yvVkFXjo+WHoh18ObVS4E
FpyLQHccruoHRGj2rqTkcbQUYrhlj6PGUbPbqDxC59UyLT8P/E+bJDCzX8ns
TvCriItARM5RQlvvPTSWexfMpiFht50V/nqqLw1iyAsxmRiQ8GVMMgDdozRK
BUbTtWkJxHo5Em7FNq2p2g7vNVa49fSe5ubEdhalFNe8ZxE+XepV8TLC7DaQ
FsO8yJw9Euq6imek2Zhac/ujp2iBlclWdiZ0ptB7U/lh6qCL8XugOziVV7gC
w7sH7bA6zC+JVZl7BoZDMLXyYRGrEVA62MZKCgoOnm/eZptvX3qSPQUsTCLG
zUQ5RmPFxBkDn+2UkeHB+FLLl9px74DDhbUP13m1NACBMyVEoX2X6DczfMae
EVv/KjSc4njemEaTlvTIQSyVCeLjyKZ0Goj9Y9JpHeJi2/Xwf/VHzoBfaY7T
bDPfGPaXLElr0EZl9hW3HDevWYhnF5b56ilqXqKv18VeqKVhRQyNEI+w16PU
P2tCz0vbSDHKBKTZ2f+GHBxZCokKVXK1g/Ikpod2TOtCc4mnk8ew9DvPzlmQ
vIE9te9UdoHXbgqujE103P3a1lRJc0Ts739tlw3pDAf6t7pzyitbxhuxNGTG
E6jz6EYFGZ3YtdrqO4fZjt94MGoVe+tsXvhnra+VyCZB7uIeRhFoThnL1WV8
o3cBCyVg4w6NnaGI+PNY9Dxb6uRXKyGD237L/4dFIV6gDRGuklJ+GiVrZYGZ
9h8GG+uE7REmJqajNNOH99YlyDQXXzKggTYvYsRB2TrSaErCasXTFKYGlRM6
0xVHRs7ZiTJHmvTe+kMUwtXqyDdafIMYrDme6V6ZMTUOUJZbL20U2ABFiBM5
wat+eimaXjgpnf3pe6PZSa77RJIvIrCx7tSKn5riUEXgWR6csZ64pVRt9Bc+
l/2smj1AKk2yHUZ7+CkbqRHO3wwZs0wLIJUKyF/54JBD7rnCOf16wYd3xJm/
rlFdBXpENGUXkAnyiDkq+HvYtfGrn+2tSHfj1tf34XGbvp+YTMQir7I5Utpk
Osxmuef9/hRcB/w1AgpV+JaDbbn50RUH62d51rMe03IG6TNx3oZ/ENx+db4X
oy9vQZXqGN2hd8ruZX4oupWxTd6DMOKTGDG6ebluajPlpgJUXBIEamdBFDGL
altaD+R6yWJOoRCOvUCgFHe0cAi6S9dZwtyJ0U/lC9yuEQUhXy2YLG1xnjsc
+VOI2TOlYMgixgsgpH9x72H/0Tr3vdjOpe7dweBYCYKbfLAt6MHfHvm0jU9U
+hB+sLV16zR7++VVGIbRvDfUPy+L0tfI1nboAlqZGWwpy9irkyiENdhjjxR4
x/meSitmQGGhgwpvVM5W4a+Bw5xc8S1FyL2Fq02s/vvfwi96s9/ynNTLZkja
gM8FiIBnBD43BzqoxplkeVfQ2wdzerya6ByIcGylNhj2DbnGFCWJI1QK897V
u7gyjqIjhWnyh58xY6NACVRrBeXaXDtVsbv/gR3QqM82qtzs2L/orunTR9vd
vfGGN72gthwfP/u7qtG9+6N1yI7cVAhldUp1FOguUj56K5hKeYDfx9jTSig0
U7NABkYKW41OZBGa95i/jbJC+E/B5UWrFdBPg0GgBUeX+uf4brVmuIq6Cpji
hWGZ9jL0g4PETgAT+UScCyIstxu+E26eLlrpthbRThyEG6F3bI5boStyPm+Z
hTogpzwiAQNOD+FW4J6/KzYq00348kdkekZ1TumivRhkDTGUL1uuFhR1faC6
/bcZ2oguoNlITLemBhKU9R4S5C1FIFhibCvzKzaP5a/L0XNsdiJk4h7OLPpQ
4a5cd0S/RWnFK6Cj1zvj61dWOfEI2in3Ww/pjxk4r6FFOzOzlUpJZIEyNX1w
kJRM7qfqqInVjIQ7duCissmjOs1kvuHb3qSE8rN9H0gLttvw8ecuuv925A24
71pGk0v+6v+AempbxVLJ7T9DUqyQRPuYWGxx5iIiqNVb/Xntp84fPo0MxjoJ
2qx5+Eszy8LKuxLW67tkjIGJ0zzKHmHd99tbOSwYxN9IS4BXEsE881C9tvmT
nPp/5J7CwKvU3pYhOTYOG0oODly8EpXy7Nss/Fha/+gjmAFiiwKGqYXstcrc
XcBsMYYmBDuR663zq1kB3/Bvu91USvdoZjGZOOYY7d1+/mMYFZh5ksF7tP4U
YT1cZ7YsusSq0F/BEn/yF6UN28JmHlQidLj9vvNj6zETk4mNtaEPL5UqVAD+
LPNFgc13zzj8KvRcG1kFmcVvQQcZIwFb3FPjhzjppltAQHLcqvtwZkt40rpo
12aIZf3MsgchLzKDmZ7FzcPTtVEOkLLVeX0aMFzvTZklVXcn3sLydyzkJLNE
ptNVSEzSXoBWpRI8l1QymX/CA/MKZqINS0jlTbxrqAGdijoeAjFIl3xMNohJ
/VLFuqcMuWs/7zHEEckjOEecgbazuccH5Q0MdcY/AW3WpUA1CGRwLtLdhRlY
8j+t41kW9/4orbIs24EcRUapZcH9XnwTQiY5Zkv1SpATWZD9KHeK1U6t7Gl7
SuiKcwerwVZnh2AkadFInwNwnPmnKvgWNqV0EtA1asamwtqF/xW+i8rmcYDM
haXz3RllGoITk0efGAsug/IcsE0rzRbOHwNKmiMJCarLch8rWvk+nBDDedrk
oYqYBwoprNWU2wJy9geFATc60Ginq53l2Yk1dy7hif/lCISSLEtbBAzkRoJI
yYDNSU6mFzDdlxp5p2DXPHDHoRt0gntCf4HDYSZDtlMKqQc8kPCBiZxI9s8y
1t8yTQTaocA2o7XrsY/0gmORNtFx10sKWcDMcioFV3LkpdTRCShqM84Qyvzd
afWMsPooqKfoZeqde4+WfDecODheyh/tS72s0vE24TpZBSpSBAwwfZHWUkv7
MbLl2mMuWsfLQdBZjcZ+EdSJn+Icbr90ptsE5JImFGz+76Pbk3fePFNpRfes
my4AkAl1mvZrtWWTY4HOU+RylhtC3H6YC9IJjKH4XZJE6btrdHY2E5XVBxF9
j+7eq0OT/SfviJoxmp3sdSAimqtpR5ArhnjH2hZZsNtAn8EVRlBqL5B6BENC
EjT4/kNFexVYnVGEdBcLhn21e4MVpfP3Z420pxgOGjRQdmJ3qgmsSp4OentU
Ydedo6RLDo7ABqLAR06ZyUP5uMvVktQwMDgJrD7wONZMtO/aBasdfoD07uvm
sTZlsHBxjJ+AGwrSR47QYMnGQHzCW0J7KfQkDM2/WFRIJw+TYhpPz3JHnIBk
Bhl4bZN1eL7IbpzMMEsQ8T4blnid6ihaUt9cbVGoHTxp6i3M/PBE73nq4mtr
iTx67DwhQDJI9OQrIQIofmnpngFhgHoMh5XXbWriuH8kWAYaMLbo6RrHkFoh
qqdeebS5LZWuFcAcX+PfC4ChqvRIKgxgndzNyre0an8+FtTrtzzeSmL/HpFD
ORVYjBVEAnAMsBinsUi6zE3x8ZW9rtXwEJ6qdTnx1jiBBrp82t9UVokAuYbL
napQlX/Gh9520TLxmjxDBQ4wdKY+7vz7zTer4RBhEi25T7GDcj0Xt/r3wNls
PaXNi2lbePIrXe9iS3GaGBNJ50TmpOI7CUGd2fOiZBw0eputqzeQDmclqNuG
FnuXjKTYHulPrNKjVZPD7IJyMHDXZBim47gE7Vn94toMbWSgPM1M6NdoINgl
WC1mnZJuajLWkYxUzXlOcqp4aWdRXnjyiPjP6w/6R7HJALiproj0qnxAYf10
fSZ4o6HdxtpiZaZyw6OmpmXdyL2bMKMAuUzvgsRWmKKy1Au0LqScIW71jtMM
AjgFMmm7pGqGEmWA2NAQojQThjh1TqMwx8UaNC3YUKaq/C2YfqbYLypuUl3v
8wMAqiWU/NHA+tkq3oHMtj63cc4tytoHAixLl8McPCbUf9c1LYS51ZcjIaAT
OCoyaP/sb8MZlUL4aGFxT3cJRrk/h4rfvWWJRVUW6FmKi8B7Kb1HiD5u5bx1
GHc0YDhcWm7piwu9WXRp83XiVSA//jI2BFXD7tDOlxi+FU9PGk1/Q7XX20UF
73ziWllxu8N3MYqhV0BMJS5iuG5P8CH51BhEOo/0p/FopRVzKP+W6lUbBO5p
hj1hx0GsTfAT6zxNO4iuoXkXfZSBh+ANzcD9dBfBv2DZJp++GhOLoJhxCmbY
Y+m4gp86/BbPBCSiA/DWfw4sHE9hTQarS4KXCTJVZrhyqPBhH7n9h8tmTZEb
9YWmmaGvHVeFTOwqLox8hTlyahJax/CIsE0N8jj4/aV4LLAIYc2k8Wc2nrOH
gntA084hCYCmdQf7KdeC8vPq3AnekS1Mc5NXz6XPSxL7WrtE06euKN0zl8xC
m9+yrtl36lC2pG/7MlOwS2NNS+FsMkwCTLfyuZ43VSyfZFe/VjSN3LNl2+yi
EptKq1PxLIXxBbR15TdlIyyQgmeRMZxZ/hkVOuLqY62mn4z2xbpKcWEUEj5j
O7xOpkLLOrl2pPH4g6yJ01Yf+fw26YJ7913tO7UEEa8oR7I0SYXgoE+JEIIp
/dynLLIWu31YxAsLTTH5T1SKLT0iXRAZom4fGp6G/Ypviv/x4S5tYEXuF27N
+3TiRRSzkB15Hnk77glsu/VZ/+whTsWMCG+YNp1mkr1qQcCItjXsB8FsxMZs
+O5zbbLDW0Ru5t7rviYWMMdUNpQUN9U8fLA+LnZXZOAK3i8VNhRnSNBwAt/B
RDJLxyKLNQFkMDwXhsjXDsSMJbMEuSlEUOgsNDeo1qKS6RDkwpORIVG093fR
7GmhC1iBz1t91SY76MO8J6ZXlx2uD2bLYkqVKRlOW0oPsZXfb29/LDumbVpl
8lxkckc/RvZStwLvUwTBhC+T0hkgA6Sqg7gI7SnHRm9oR0NoimvMkGs64XDu
n6c9lc7HguZB1l3ShU4HUEOYoVKecm62ib9O5JnaM/yUvUmdJMipmUaMyCvx
ifdSZWfnYRES8yLDgT1DJBfYmzAu5lCHhXxFA4lQv6VNPWFxpuA7Yv8iHRKD
ngVyA8hN95qvAzZFS/+amFmzQFrD8AB3pE2iiyh21ZcQhUw+pxByo3IQLBcE
6xUbcjuSZRhj04e6i47tqr5xwBozi989DlD6ibvvJq3zRlp6hWqbwXtnkpLm
iLWQY3kvhMBr/T5jBFiTQx/ki24Rfi1FZRSJvg2MaMKp8PX6t7cpgQK8iws1
5Yvsik44lOtn+xppeqhvpTl1x4nOU7B5FQ0EJKFePbYOoeP8ce213rodGUNK
gqav6QyIC4tj9gw13GJl7nrmkZycEQTL2MVoSgUzRFcfXQLpd31BMTIl+plV
ENf6OmSTKWJ9Jr4Si3l/v+9zFeYSU45jFUjB4+mUNKhZH8QgGYyzQSGW9frB
Qrj0L/V50fkErMpgLZSzETwYkNCMMpGPkAdio4uXRGhFp7qCZ6rmE32qqncz
mN4gu5exdy9kzXOuTo5SVL+NKp5qMSSi73MVJ2p8wnarKYusprLdEdhFNYww
btdffhF5LPLk9de5Bd1sGQZFZ4+fniD8ZtZa6DN5HTesZLCrXdmxRQlYcDLL
6OfBwFYnj77R47cUS+2OJ/VCheVZOGSPexwYXL6nPHfsnX/cfQYkwz4Z7oga
P0R2Lmk0egZ62BhzMs29O+xtKEsMvD9HYdsqSBo+nR9tz1A20IVVegGqAJsA
f180yUh1qVPZ+rk2gBQ/wqR4ubGVlQDQVV0t1DS4KKL/NyagiV4IJ5NAcTIq
+Z95hXDZml0ytTn3pKrXpDQx6Nkz70W962sirisBdirXWjf8eoh7C58UeBR/
U5fiXcnR2Pn52ztedY39dCJNs6qeG56MEzxUQrZXkVElIxSfhrdSRbSeIpm2
o/annOOARovlUTl6NxX8kwsc+t/sKTaPLEGto8s8hedOtucw6gFXqnQDLsvb
ocT5ChlaPy8TMJCv2Gdhs0mO+FUkb1XmMwbWV9VvrAniXhsz/ibrtKNTpBsH
Z6V9PTlYNyTSQuHoUnoJ8UHpbmJloTRvGPijV6IBtYDFcGX7EYDoR8++lXXp
SEahqm/zn4DJNDTlV0HsCezNrXTnvvo85/aFxcKYmlPQLg042JYm8udvRhnY
w4DopECymohruKLaLthL6nYjxv++/9rFn4I7t41gW09fuK29mvDyJv44cerF
4Bhhpkwsr8IHPD9gzBwqRT5BCkozbiYIhZbVetZr1sUkNKhnxJWAaeSJlioK
gdwNWQrRv62bfHDisThe+LcrrGsOiPkjUv60axIxIhxrh9fYooYfT8XN3ryO
mb40zCsvNaWgg9dwy/V3UliKkalCwTWjoSo0jh0ZA97GkwS6mvYKcaoRMOJD
9bHvXietcGhhBdZ7SGXolwQnB9pU1NxW4JnDRtljvlvpLNX4wqweH8ddIWcb
ZN1vMrakejxjKOL6Qsa0s8dPaXRhZXCHtOCiqDfRUzAk0vjkM4LLtlE20/2g
dvl1VgYKvwdK/4wiHhRRNJ1ovfF5xim65eelOrRGhKl/lTxwbNqci4JERHpo
pSrpqfz5Oqm+LZjU/D1GxOgrpWgL7nBaayZHHerLnttIHlv78j/9FWgMhJ72
dHSZKvLRjTDCJzzzvhHrgq8nv4WvfFYxJygOIz5wkPMswMb3OoCwz9Alj9R5
Zafd+rtXkE2vY/x9JHVhlVL5yRjdap3LA9ZcllOdiIp3JiN0U3psT+0DHs/A
D+fTspNxJtoR2JfjhqizYPlo6O9zkPBuwHv4pRzKeaNLDeKLw1tms3S10+wx
CpO+w8oc7YYLxfTbNEUHmO+moedDq0xeRLyF0wm2rXfnztCsTo7eUCyxbGeV
9rui+8pPaqR/trpi7Q0sFZE+7ix19jCPuJJtI60O8wMhODVWgTbCcqrC1AEO
a/g4dCcdRl5nidR/QkLAd8FSbnePtZbLtBAp9o6uyBd0/88LrFwjCHBK4vus
AJlsj7PDwTtqiiHIsDT60oG/UICuczLwi9k2VJfIAvKH2VWvRdF3QymmeL0J
DUfD5PPkBxXnOw0rCJULPU/SmMDYTuXrzZdpmINkDGcdi46q27moy8rchRnE
yodgf/9XHtVrAm7xG6u70Pa9927EhtwXPim3ZqbwbU8zvHGHgatCQS5rkFvb
NQRjmF7IguchzWrXtAEufmQZA/VaW95PeF0JIxTonZFlg7MQs0ukM2/J1vcE
cYAK0PWhshnhju4CWU1v14gQhVTb4pYyUfY1hdszrvEmr5yWSPK+6f2X4Al6
w0mtO0+jYK4t+n16srantEBjYL0Be4StWb2YhQj46lg2HqsCJZe/CZddVE4A
jI8R/yMu5qNDBCSV3+KpFbCqGPvSCZET5WsDDU8j3KRVKd0rlJRGQUbKKtMd
10/kT4kC5zvWGM93RChcYW8a9kSC5R/PymzSHXU4vowVaTBL6O+q15rGLOIk
xWa0cjQ43gYXmw8E6PbAkz9153O6T5Oltlfy+Pb/uD5qp9f5BSQjoY/I1ccG
sMBK6Qnl0O4B8g3ceAPDbCycRePpEJ2gSw6UuUnhBGyV2knIZHsRN+9Ip697
bjwULcPQMpgLkSX5pBeB52q0vbv+9+9S4hC1FRNtRqNtYV0eNJgQwnRwp6b6
DzdNGopWIShiaVTrt5SJGj+ybuB2AmmV416f2sc/gxv/Zjjjlot6jY3Xth5v
orLhZFQWiZ58d/eWj5SRd5jR3gMm7+vNOWIBXDUVAx0KN1JfXTfXvPgjVRbn
hqFB/io8LCP7612QE2ZtDgEyK2p9VzSIs8vNrNpFg7BwcX/InrPZwTcXx5ad
0u04SkKfju/5qEgVFC/oIccmk6j1DZ7z3D6J9r4pnjTesLCtNWOXpkpP1nhu
yuv0/HtWT3a3Dh4kctjTmZPX9oSPz/flAuGDebkgj70djnXjEmoadUFgWpsH
trfrANhZpVreoPb6KycD0gRtlV2UttLIczGQ+Hxb+S/f7o8qiNakK/gdzT4d
Q8ExdaIHIICXhuO+DKW8/WDqXo03C0tkcI76W/vtGWqpHiluPsZzsDpAZSFL
sMXMjv49VUeTK9Xw8oZI06kRtlhabyhBlFJchi3MZwz8yh/WBb6axYRUeF7U
TX4OZF7ZcYFee2SNecP9/l+P/UVxnXmHSHxEjd8dzfAE5fQz1NYoSrQ+XtOt
406XqpBT+LQCnUnOfDxfRtelivgu6sPbD3sjxRwXg8/sGKvUMZLWDxtkPp8v
pkWOcNbHFARzDtJtefyPQmhmsOFToJ4vFmIe0dIYpxIre838ovwp6zbi1UdQ
jN2QsJwQHDsR2oMWYpqhRBj3cTVmyj0XUMMgtRwwyd+BmlXCKKMG/zrCwiDE
pLSXXLMlaxnA5Dvzx0v1Sjo5iWLmg6WTLUzNQDcnvTOIWAzgWUhWlv6QT6fd
CraQ4u1UlzuBAWCT47ttu+IOvZDLR3eumgUleDUner7ffbc+MRfRKOCqE7Qv
wtbkYWKO6Vwaoog3c8Wccax8zq1+gniXx3dnP7r7icJDbpbb4T8B3Os+uaSF
skR7pgRa6bFIW1Ialvc0jfTXjax2yiLfU6G6HmjWkoCXvjC/wasbUQ5E7s7F
C0JLy+gv8kPzw9VezL+02IiY3pDOVgfAWJoxnC3ThNUtAlboPWkZkECRoLwE
ICwFD6BQtI0PJ5XX+GFcW+ljYoTFyHylrEpiEMoqZVXjtWlvJQhzkOSL/qgq
b8rcJ9+TjqeWEyJc8VRgbMmL0DFAXnvqMdPX5JKvnuFToqngZtKcTJyp8IBx
SAtYMidYuDeA6P0K4gnZ7w1wbdFuJIzATcDY8A1JBnX7idDA3rjuGrZY0dwM
Fn52i7AcJ0NpDF0s7xbCcs+2Kj2b3VeNL9rbhfNHKz1DB9/5oEmJEl7xLvSc
vd0NnEMZ0dbvCA0Dah76dOIRFIg3j8LuBDIlkVL88+0OMYBYSSVK+FuZmxNZ
vm5UM534WFgpyFbBDWUigJTvxLY5i0vAur1+SbWb69h3qpvdBlpZN4G5MskB
FQmMAHGqHjN+OZYMOwktdIymYusOqIbBBhHU66LhMIMp77eQCFlnIv55OfYJ
a5yklGD+w5YkJrgoDpEI0rzVgYkSSRseDP9QeK+ac2Ez3nf/pNxJwPSHZjOr
5Qqn7RZVP/h+BgBgfC+zygysN/ozKUrO/LFORhKQKnPS4Nn/pJMe9ggBIGOG
6dE/RYilttmqYv6F8kCfbTWdkxsDDFdcRqLbNHe2N8UP8qCskCm2GPcAOjRW
+47w5Rh/lMK0AMM3YAowA0KSGTVK5ee3t/RairWcVuyIKYkjxKW0E8SSa3/C
03hRK6WAeRMI2mWR4hd6fK6ipkzDv08cn/oIpk0wI5Zxn2Df11frDvomM3Cr
klYIsV033hvBa7J4uxHEKyMM9FFaegonYge05iBDAWFkULI+9PKKQitspoAB
s0v5TfxkrGAOO/W/dpnoLqzrtz+4+l/wwlDJfU70qttFzfwV/fwrBIbL14hG
AVUfxfLe9LRb5V/2bKDZQSOlFZsHVxgbADl5vc9NVeWloiUBQ2fvygmysayf
3QvuPmwSa9cWbmZ+UXYFq0T19G9c8lKznSPnp3fgEo0F496Q9cS6PfvXzlwm
UUNVe585sIWiA7NtspHqgTLWuQBiLhYjc+R0q848uXicGxmOmG0BGeMUnH5d
2zrExgHFvQBsyqBNiGv5MbWH5ZeA4xBSKk9ZQJtnOJdZbYqLeVxs7uvJRk9+
u+hNQd/kZ+K/za+AX3Ls2Aws69MyC4hESSvfOEc/TpwcQAl6oK7Lpnq/it3a
OfAikAbHCbfGdYyDeX5XQ2XK2gCiunrJOHKUH5JqUELovmZbicvTGfDCUL54
f03W+SXnTsXfH0ulUdSrftNxHtxvklHvI4+jmBD8ky+H+ed44O64lUveFaUb
tEWQeqw6EzmlaZi+7SfLZPsrMpi99r+uUr2SMakQEdNKD1o9jl9zCnERn3l3
htHbGMb2WUFdlHiWnaJaL4P5Wo3+2sfrJK8xUR42eal3hVVDqsausCQ9UwaM
HX+3gIvKyqqZAkO02xwz9tgWLTnmL5MNs3AUyEH3N+xbQXdPQWBCRxEHTdO4
ag/v/nXYJxjnpyOLPk+5Hi/9HCuBR4ZGkjQTt2bAoNQGAgR9aaABYyC8JBpV
bsW4ZekDX8NmHZMyHNJg2p8COrLKCao+QLWMtObqVqBPACrnfY68SZYHw/Al
R5gt7xCc1M4NHcMLHVq0V8ibrML+FqhiLWHFjuL7RFkuAOiGKyeB552lk6c+
psYvETvWoFO4C+fM24+It5HF1gIc8lz+ddO5n29JvYye8lIjFrMrYdd6NQFt
cZmdZSsmNDPUWXggIoGDLezkPA9sHNBzx86gexPp/Wzt5lJRZqtp5b+lqh8A
mFyzF9koz+64EcHWyhcdZdcqGiaVNig8dnlKMUinraK9uHynuv6lOL/wo7YX
f8vPcrEb7G0JSF/YJ1d3qO/AcFhFK5ErCwQw03iBHbSvnq0Xn8HL1fA/mpXt
DXqk4Z3rQpoL60YOFOZ1tSwBuXNeogYP3jQ1/l1MGM+5K9U/2AV5T0qmi5GJ
Nckejx+lcHnsiatw5V5NV+c3auZL3zkFyb66DJyUJxegFrOSkBveOzjS3LK7
vc360F2RkXU6l5YSCfK9wX3uEINSvvZrCivVetTXOlWQqDAKFWgQELTWo3Km
2b9wTDyCE1Hn0pCj3Ef7q6wTlzSRAI9ttNvTcY8KxnhzbQpYuE5g37gxerx4
oJlAokaZrTbRs6a7hG4lRqgWvwhX4xgALcpfpcB8MUDtBvHBvAaLTePvvZ5d
lE9xqpPCklrUTEqzrmeewCRLCRNHjrODR8Cde7B1ZbJWxEk2rl7bP4c1voAI
5LkNuLiuRR0QjlZLMrsKthhOmVAkjrvs8RAi997NEuCDwZJIS1MwoCjgfFuU
Kc+p7oQXF3wWiQBmf9jnNj7VuNEa5/vewY5HG6vYEb1ZY9rvb2vxLP+ROLCH
R8YhjPyRaluZqbwErq6gzrk7m3rIos4uE13hc05SQD+QqTLxVVJufnUE25qo
SsCU58GJ4JdnrwrdK32EI3Q9hg4YHgE3CiAIK5Pt7Ooz8hFb9O7GahREZbTW
xstNG/nvr/yCpIm6JKsUnPe8YSbA+Ned+TYcbxDwcpwCYuxBxPBBSWluzezq
0JH5GgjD7nn5V3d5gCdYeZKRzS6etRTDYncse9N2Di7ovMQHk5dYZmme/JPH
B+sQUmaqG7+HJthYvZ+5DBxT3XItjSv+reh88U2ryBJ2f02sU5cxad81SetG
vyL7BqxkrrKFFgyxaoOZOMizgxGpc0Xx/pLpIrme3oDbQp6NFwflXJ9LZIee
+msUrb+sC1dH3QrAdrRXSsHWcoy0JCNbz/z22ahr8t4gq8qPNEvRATyOmfop
+squhMZpIN5E18zrcMarB20tLqA9gn+K+yURt5bZlu4rw8BKde3DLvf3k0on
3TnbU6NYfRkj5U1vh9+o/FZHO2eE04j9L4rF/j4zT+LaEpLiwoJFI1lxL07g
ebgRVulu8zAjnaT80vCAk8uR+yEzh7qqybdk9/KKo/ojQwUm3Krtgn5DAeRt
KleGJKI47hqniYKmNfPmccTjUO8bO/a+KOg/PlR/hscly1LLXdWfwQYeydf5
Vr0qxEGsVLSo4hzAPHKCgcCj2wFgP6DmsPtcND60O2v9Zqjw0QS8PZT4vGR6
085YNO0TjB02LMUXxVu8zOAZnpuYTQ5B3Ytcq9ddbc4HMZTERhwJakagNF8z
A4TCOK8MicoT5+Tvs/zlkxUtQi/VOq3rQt6Sf8/QLUPgQzbnAwnC47vzK2wm
3oHZWfBMCdjKufzg1ocMLdB9kg//WiMzwnrlZJVYGKzSJN4tCW5M35QoPkeR
oPasUCq96IuCAjEh1m4i7KgT7U3D25H9+3FSylagGXswwg8LH2MJ5fQprn6E
8OU1KjCjaRh+WL2hCZjMdRrg2ZMAZemst99SWX2gRYRDiRoFeQdMcn9HRfYw
P6cF0aTdU6KjmQfIJqNSzBaE0QzKqeK9Wd2k0Qp1RrP9GJjvrdzuWkrtvo8j
VtpCJBFmhEtsSQE2Bfb5Q3cUi63xdtc4VEofwplFzlfPIWdPC6sRIXH6uk+s
LQQmakUKODVvXJF3MzXKDpiCJpdqC6mIPS+rw5TSyNvU1yTlMwjxrX5h+Xz8
5lEzsxkuIHnfBGffcc4jsbwpORYlMspIq3CK288sVAEMYXw1GmvsBBpJAmgj
T4r49zfqS8AFkiBHE6JqyAI/MchbujH/5Du0d3OZVMPhhBKGoCQ2Me6ZOps8
SUeVZL9VGORPnxGRxBvGyqQtuvljLbNCyhycYmhizqRxnKY2OS2ASzTUOJpb
Ii5M7QQBItUkJPX00fLLeP+VMeU8+3STtl4SdKvNKAtpC5kg5Urb64xiKamC
bzVEWrH7R1KX3xhDBsm1HPEj9h9msqHLon+bLbb1rtyGYKAlXEj6rtmAMVqn
G0x7qVQloLfjek/Hl9NJYcQJDDMlmxH+GS0C/brysuLd5zBYDhZD2YbQ4oU9
TCT+gYua5XPzzo0tF1Kmpa7YN21/8864h29dS9ZEdCanX880r0VTA+0B8yho
93Ahs4OItERhYQ3pDCvzus/Ri9uyuSKKIgnnAV4/orJB7zqmORVxk/8Mis56
LI5eYywpbmmsCx5zTYH1ZmncnA/oa39WWWeoWzwr9kHfOOX1cKUbZ01fsBdx
xjMLnUQn+JT8JBb2zI/cAR3/LQwzV89gO7x5QjaO8aAlLKFknyGbspcGBQCc
xq2VxLEfJUgLB/d6vPOfYoejA0R8dhJHqhI+B52odOXrc8GskktgLR7Mnr28
NDbhfcbBpyfwcGu/bN5BQ5QLgrwa7yGgrE4IaWMMwAeXNKL4bVeB+9Q9CH4F
shTB8csarg9PPk9qghFsssR6HwBW5EUQ7LwiRe1QYqT7ZiwraP3v0miVuN/b
rxqfBr1THvEYQl0BGL2MzVOMHzzjDo6qaqSJT6pqpUTRPOZI4AueNt2nuBki
C/jTAOSyH3XMeGuvnoJZ+3ecJp/ewN9zLHp5wVMf8UEBRo2svy1/5YBjlqT0
SFVrcUSyakHdOmeH/qSwVjCDS17w+Y8LuSMdesaRQytJuigbvrKfUriiblHd
Ay6I9Ugc4WDRF5bC4zOt7bxkqE6XLjoK2EqRalAvwBcqvHIR7FAOpwGZf6Nt
EJMcnSt4WyZzPCc38qZHpfzpckke3OiUJPUuUOzZ7goECZqzDGWGUofUOfHB
2rkxSHdrTnkWQBIsrqJVq7TH057i6wE1dqcd41CwCdAXZoJRXQ/q1/8BX6qX
GdgCaS6S2s0m7Sbd90n6hkxtislXX7tOXRZD2mKEaNRP9zIax4V9WM5bf4WT
at8G8sw5vBWgJ8FjFU49kjqvAii3RLCAs/yhMw8bQ82dQf4G52PWaopJKEdN
l9NI6TO/JOq+faX3+/oWjAyhgZofSWMZx6f+7yt/2j0VORS7wekAHi4ntv6I
Jyvm4/SvI0+tAdbY1DpA777BOYCyvx3y8/1VQb343lPdYnX+oKVLJOuah4Xz
HSvTFh1tpy6X4Ltd8V4ymuSPkg9aCi2dzYAmC2aal/HyDeO9mT4s/SAg3vwS
Iq8E9T8OiBa0RDHBCscBhstSf3XGlOemwT11EMdCMYmYXvoSC2loVnZsvqKN
WGA8TiN2XQyDg+oD97H/3b4EhNqDud7b1T6/fOSAKjAR/4Or1B5277D+CiNE
oroNDCRBIcMiF8y3vpHQEzLuTJ+2VTJCJ16bfH2A/Ixkgi/zFdL0SQ8NDl2c
tONZ6jk0zaMzF/tOy/9EEaDarf5U4djlyeqjTRCI0iFJyKGB8NDA4l9F+Q/k
YdqWG4gYc6zP/C+iO7WRrwX6EnsE5Fayg2bJIkoucZlYwI9FM66oEPnDM8rb
EAbVLfcFakG5mcIK6+WrqYRTI5MCadVwUREbywcP2uJ1LUoCEEXIZXFVhZX/
jkhf00UtC4bRnZk/HM+bdTyfsy9dnNYADe0YS3HJOe0x0lrUMbTXELF4067l
O+twq4WAFhyjLf2B+HFAsYMpcpep8LHwqF0/pqo0KBCst5cuXIzK1x0jZ4di
nTK8H7n1dEBji893bDas2frdQo2HeIotlwJhYQ0Sneyta+0qnwLHoCFP5Ju3
1yvCbUMrmKozJ9eBjhMgXCa3q9Nz4AidbnGwconBsESVcANii8AnXJXuTnJC
FrJhuYlc8Vk0pNvxrxGj0OPjK27WDl/aGKUF5DOi7YhxmWq3vnYjyqWm5rpY
Lsq9qs0UVDBDaS2d0j6M0GBqRS4ItXkTZ5PKRCIOGC+OTJrKYBXxWucBjuu7
o1k7f7rAiPT6Bx2kGoasLX0wR7vQ10XYPRlZVwe1TIxLm/GRoi0Uz2ITXcf5
LvArzwUvQ5gALAsom3niE8prRWXyiP0MY6b03iGVHG01SjwsLJzABxBZYEq6
iMvsp5eRD3cFi+xR8Xvtj1ONDoBBAgZXg3Y6Dn3GJ7g8sY0I/AAB9H8nXGii
/mRzFcrFWtQbuIMS7xNg8GWdj5ltuPY5yWeumRwJ0/+B5CUOn6SrIHsOVWcg
elUG9g8Bi/g8AhJYizoJT03/ybgS8v7/Pcc5NJvHAJbZ0d33LW7BTGBIielx
I0QOa9jhJOe+ybpLS2RCV9yLDjtNlrjtAtCKnN6tNo8/GJ8sj+a1Kv55t4qE
zJ2h7eN9/nszvcAlxyXlgnQB++9a6d2WIIBcqzZyBeaNxJ6WqVqi57pORPyf
jw6Vq3gv2Ptzd1gsro2ooTMnD/BuidsPW9gv3vpwVHmjAEhRnLELNR11Di/a
kiInPYFuzJ6OX7Rn1/YnjiHVABCVWfjE3iWeDB0xxbQKtXBd3asqKKwrRyU8
ylkJ5B6ko//N8lt/D968p2JGjgnz52kYWyGsnLqHlgIZicSJjO3NLueCfNVT
mQ8fEqk9krO3HRH5QIG5oCLk+kIc8qU4DNj4dZsqG+66CiIFunvi6VaFkouI
YE4aZ34P3oiN84P6XTZ77Zm5eeEGTY5KwyDukd1q1pz5BKIWKU4buLi6gxxf
hfnAITd52IbvMVuf336apuTygN0GxIU44UA4mo2oS+rvC9CfevM1D0OHscpg
cWVwkWt9xQ7HTRzwE1mKYBFShN5/NYfewyIAsqETJvud09IOx0QUqT58MPWF
KndFcoyWFHgajOVfT42OCVtxwytUE8FYg4uGd9RlpHbqW++k6A6+3XHjOyhO
cOT062SvvFJb8Hgb7uhn2aBSyStz2OQN24k3FXn4HrHmvxgWyXyTW3PQIxhM
cW4SIXEu9B8NG55t4FzF8vHNPW5zbzCbB/LzMNoWr2TkSL2rZF7bOMsQB2NP
LOcdcMVDGUQ6Kybu5bDh4LSNtuLMvJKCvAX3FJBJKOwCcVSNlA3l9Z1e7jTf
84dMWQBr8NGui1qXMWFciv02bfIORBK9/lB6eK8yurfVpNhDTZTwB1M72/ht
+JKalp9Kh4n8/fK57B5q4yr2XyQwm2AtG6rrgiWhvr/fVgRN6XBq7fg2uXU2
TNlEepi5Is48LhTKOxyaWnUwNTLVy+6JJX+8pLWZVU8Nd9AeCKIzvoRnoGRE
/qH3BEcZQtmNS7hEe8rJnuGLuJJ9X15VaJSKE8ZAdnGgkOS1Yhfdef8kvJg8
1UsjRq7WNpvbkma9XTlICUg42sZShFnmS78YyzbdFnHydwQQPQ19Sn5YJoyN
AU1619mU34xUa6av8OA5y8hlNk1ezeKZPqdMJ5qwWkBHDp7h4HwUTRgqRv3u
6R+U/DuRp4w1ZpikZduIP/PkUwX+MCH2p3GApAraLg22a0Pl/n/mTbQEGnbb
byND6sI0S1WE9DsK0g2HhZkxG3BhmkyvXsf9C4wGNJNC+P+oR1ChWBuNX5Sk
ITV5BbbB2BD0aP/COPow6+Lo5kTrahNmhbrXPSfeUyuYEmbslCiHlTUtlMAM
6lGOh/kWiRBRrYbqxVPx9jhY1HsxnE4h5TUphFOdcgK5SrK6tpT7r6c1D+7i
7NDBuVq9xc7NhQUo2s8/BOvYs5oLt8BeGhQ9JhrSWd0lkqwuQfmLXWz8a3Vf
20iPIrDoQzliAf4d70Xbnl6vGMBGc92khCsQRn5ma34UChwzUmycNUgn7GUp
sn504WCN5HS21sW/cTqwKSEHvmo5KBrL8tQQZfQP9trx4XrDy/lo15mAflQ5
NZNJq86A1rjpckz74egb9B3uXTlZVJvPTSWSAQ7p3JPRy2WMWueVNbqvwUbz
FJz0lDS/NY2nWCIIvB6XF2gUtWs8g0jgQV074s2yYnIjzo9i9esD4IQoDeYN
9LOErMweVddxzbswgLKj6mGt6mCkAnzBBXICXPebY5tyKTJGi0o5p+5fzitx
R9PehWt3TGKp0uJYgmRzcE8vUufERI3wqlxNj7Lh3fPHHRLRO38+YL8a10bV
8VN070WcxkCAuFSWZwUB8FVQcH5fM+4GT6idwHZCvF9sckf8SbkAB5i4negz
fCADYcdu+G4hekf9BQT8EYDKhwr71mEXn+hRSwMmwuUdD3RNtY326n7UKq1i
L1AcTLJPCy7z3uugw6XZ0my7+2u9tWdi8bXqjN4GVGeRV07LdI5ZWu5TDoh2
z0I3iGcXUSP13CgiAVGYYvnIazntPNVLTzq5ZMD2jOwARNJn9L7VLWoZ7DwD
7lj6jbWF5NyoJKLk/2CfSbKC4tZCgULNf4P0McX9zzy9mhEhXBu2iBhgYlnp
5G3AqZtt664yuqSXL+U+FhQ9eaN1OOtlVwJ6aqSD7sgI0r71DSRMXcdkEMIc
iaiqeXFaIjNwCiy5CayOL8U/e7kVJ8O1LG/k20of2SL2qn1vU4vp8do62Epe
Z5kNjTv725BLlVlVXRuDT6ukGgyLMWBDYvmc50menQ+/uMoRV1EtDHo25N3N
0IJLq5CbmO5MGwCIfZkGH0o9A4OwE0bFMOjKrE8BbDEbkDj4Fu9DEHWFC7Tb
Zd3eJklPoBolwCyLLMvFcPBmrLRBD+PCo58Fs5s92C77BuERd1ftg1ss/8Uz
o7PXMhtNwYan4+bp/F/VOdwg1o744KQSaM/V89xlfwMpN+gNdwstQcT4fQaP
njHNTmOl6S4jE0DY2XJInBo6AcDw+iaNIFpvjq+7uW8tGFsqX0IZ8uMk5b67
O0sFvxN7Oy9pFfc/ZCBKKHu44hOJ+JVoraHIjHGTHFmnvCVVDC8DoXMCjpF9
/dt4RcScCz6nDYedxkcZk9K81xigInXExq+NTPOHibZ7aapKtBL92GXDNb7z
eoKQvqVIVrkLNWaZ2SQ8xm4v79POsIIJJ2v+Mcwe79JK5hZEZYDLmMPXv1PR
663TfWDC2SaY14QVr/7WF4uwmZuOnvwZA7f7rbpflFpdV9CjkuRYx0h5ilZB
WK3SVJ72NS/pB/yQpWbfgVWOlngZ1toIT4falNoobh8tGPiF+fpX7tbEg04J
3NJB+8TE9tVx2sclPzq0yWHHxT7tHceK8+yH74dT9ohJ0DrzkjSml76unRz4
yUbZPHbVX54+mJ8Mglp+AlRhBeSSrVxMLmGl/l7seXuDnLwm/vWz80UXiLAZ
GdL1xsBxFGXHJxWQoyiLsXECP6Wx9jCfIZ5mwgl9vlmFax/OOI3BStZsvXG8
QmJwTG4Toa8iGX8AjrJZW4M1Lfk6e01+14TzHTawpwZRk6luKkVQw7GTMZRe
/rGMIjbjeRhQA/T1xlek0lEkz40G1+twHcj1jum+JSNHGmFMBSsxo4sdAIP9
aEChCUgivyvIbhNxFY7E7ff9CJJXBOeaG2OCBVafK7i8vQ4BrOh35E8qvrKo
KCyPfRnIq1dCtBGbe73N8wb5grpcwG352+mVNFMhAJpGCQd41OED5ED9nPVl
3KmiPELW6laTw0K6y/5UQ4+bTKRF77sDPDWd6gruxb+UzirgoiGzuRACr3YL
W/ns4k/AMFg/wfDcS0tCuuXbh61X02RsuUt2vhK0leJO8CR1E0d7ixHFusX/
5f6lbVZPS/i62nYMKPXebCrNgr8IYdj5GUXrJrVuBdmgrnph5loubEgminx3
PYtTryn5V4WEBoQa7glUe78L57BlNv7Aa9+TW85llfrdxGKbOFvd29geBW9O
DmJEhHGkSCjhRb7eQBTuPy937K/4DQUoFhH2jXzDDiibbMfaaNXd5ToYn6Ac
SruZwPRa/O19C8NShfI8VaL7D0xNLJ8LBYW4cX0RMewKBiFuc3Yue/GMLlQZ
vePNytsgNnVmkyuX0ukt5BHJfqCokwUG04BsPga5F9POb1GJAmftw6RlGCu8
3aNm2iYv+Uu+AjAD5m3KwewuCBZk8Ul5kCM+eNSV/VDB/+qj3aheL8kGwpfF
0q1gHC1LZz89bkTUGnX1HH5JmCy8FO2tTUc26c82zKPIKQOJCcBSANT5EMMS
deJdABcyjzDNso5d2nEZ3EGi+vLp+44A3x5Ek6ldi6KQWrEzsrGvdHTA0UWr
iVwaaZIlVARTOydzDeW9BMwbtNcShRoL/OHUuGXeSAayNVAXWT4nJ8fHvkgY
XD40/i6ofY8PMIMzDehsYBQ1spNoZM4KQKVe2MNRqfNFLC8Z17Wb74c+hWjb
35epz//KbjZTokZpmH4OPUpXKXN5L8Kz1jsZKBZP/qawqgDF+VshBuuPQAWY
utGLsUmNT3CZEPjsPDhXhe487DzWa+NsDSYOcj7oarS8DOdxRNN6uvpWFHds
D60pC4P7umzKVYkQXDNGUroMw5KZV3pUXdaVvh2biEdTgVSRK5M0D/5waYRF
D0H09hxBMjVFbIgxiCfopJJpXrfOiQNcSF+BOklS9E4m7VMEIoVL135sWh19
xn9XrajmEz4x4W8shvul2fquT5ODtwvvXbNn3nKxST/TLVNDHcpRqXjav3lx
YeDkV9G2rmv6689Zy7B4KZPcKbUjNMK2ZizXNxTiNVhOunu/LwyoGr7zGwtI
zprXIMkHkaG2BfEAAObaBTH0qv6OhdoTK25F5tnLpQ4FSOyPDAMX8eahWSkB
UZlLNUJf+A8zfrugAwAkXXhFUAEOepu2s8beJaM5ZVSAzYpQ6tArv6cNQyux
oWrt6R81sHAfoU0k2llrZQ8SYUsNl7Vlfh8b+HSKB4VpO5rHrMWI3BgzmfyP
YpBh5mIxyyKvfWR9+rwI4fe51/QWhD3R1AY02UksBrxrhhRzqpDu9M1+ZcZT
zllEG5Ikva8tsCq7hBgq28TiejheXNcbcW+egqCmSpyJZw4NM4ibW/k9aqzm
shZWbq4mom1VAn7FAJsqPfjTr3DrNO9CL8bMGsEtFEbS3kyD/mXkpjmSQ7wA
GuecJsz5AOspdKuffnpbXJ7Sf34udK2vTJ0rJB1IvYEJY4A2fCSvNHbSSdwp
l2wMpZJ7E+hTjJBGQQqFHlD6bIMu21vkYK+l3kZeVziUC/OWGYTOlqUk+nQq
mwCiqYaUi33Z/E8uibc87b8lGG+aucC9RVqhL9Ht1dNXjAEe3zQ/xjClds1U
Xt2G3yrjz52eyAeVdMp9WUqC7umwTBMGndyHsI8A7xWvYLlIUOszcxb50kPt
MRvwxo8JBPA1pbNHqmd0fM5E5Udo1Yp5T2090nvxDD1NmEsqBQW/RUp4yFpH
O4KP4iucgeaoIo8NnYjv0apA2jUy3/BjpECDDc2XZvcu6oWlXh+gnKqBp0XS
0aP54/pR530JDh2aChSbvCoaTl6Mvy6lugikcyOc4/4OxG8BrEykncgrM0Mr
BQ/dInBftRCZ/VTPuSF57XmmTpNe8QdfK14a0MGoihgDRR5OmFOtrHiW/0xL
n5ALS0A8AyUF8qkLzp6/TKN0pd1MQTbl5POao5iBiL+y0rASwP9r9B9i9MTq
hJB0jhF+b9fIV2UMldl+QfPgHkDVeovr9MX27FV5sOK+uC9t4C3sJBs5pn0p
4t6hSNmqRyReRXsBvHjUSC3eZl6iCC8u54Ir9cmO40hhbrkPfXJABYew9ea7
IBa4r/hhb/Po2p/ht85TtuzjWbO9PvBkxOTVHpztb+Jhmw0kngO8KVrgpiIF
5G08kzWo5S/njPuxfoymduWULnyUJN86dFXOGQ9NoXDGcMBK919JLx5BUvaC
nbfbcOUjsei6qQ3vaJnEitJiq7UL+VEhocYViLCmbHrPGQAmPBqonaTJXZ7s
vvMkhrAwkabc8T2tJRKbR3PqMM2DMo5jYNqWlkXMM1zCiSRNWN907SUoKLJQ
xPThhW+ETGMKxTGZco2IGKWOOSep8UAxTxjT9C4jPOoBJBUg3B48JPaDc3ld
hjbxC41ggrxKiCarg7E2xpWiZMfiVKDc+sfJaW7BeRnBH3NCIEtys1EL+JzL
QATmm+dTMsi3RBCv4D6DQPJxSvACJJoL/QDTkTfJPi+KLXV+XCcmyCAk0GSd
Dkfp5mKRxkr2Hjqo4oFWuGBiYOlGR1byiY0F+UWG3WlwF+IAd9upO/D68GUd
qh5T+hRciJejkFkMpQy63slc5CFrruidAyp3/PaE/hoJlcpDIM6zxkOpPdAo
Mfd39OVtoR5Nfe78gODaDWbr8HpEjUTCx3W2qRGKoLIuvJ5tD0fAHTVVXwfi
qGP4AfzT3nLioETFOjhfJV6dQx3/AlXPjudjSFyIFmB0OjaZLpNsfNryAGVL
gf3B6XQDlnoZSKQMMjKNra/V5YhFtE6nBgB00xwEcBLZ+DHNqqUmzq17Z/R+
hT7t3HRjwZT/Agrhed2THhU/ixsVEiqpZwL8eBdiNh5BQ8dz/BSZy1NhOeWe
QWkXZmt/W/07p4aqsm4ZBnFTd3t4d+BfLQsKph3sN+1b/fG1jylcSeUV+v0S
b6R3UzS90tv5MUfrWjPjjGEzfkuqRgQeXKjBfKWtjmR3oYaZV7EFfXzOkMd5
IjstjLQaxndCiQq6iK3xsYLZD0I3SY1KuPpOpa1jKw0gJHNPBBO7rflcZF20
AAoTOQBtkAldPjCo9c4UkiHdBnKoSMk9roLtmlKxDQSuNs59Vgp/ZATqQh6z
l1/ESn0u++VP7KWL5YdOdhH4jzN7pAbpCMcZcbOJCJdy9B5Lojd/oRxKB0qf
euUxMWyjyfGPUcUrB2HPSJF3Kt5orvTEh/v/VCvxuzIUZpI5MXTn/ylX6Oki
EteWA+KR9birNWGpaivlgO9NuqfyPhc+NClZ7+ODA2R87FEApB9UVkP1Q3Sg
4goLHkjvWnvWUvoiga1IYdA8yTU+S8+15VnyEV5R+r6Ef3wdZVismulL3Z2C
Rjet5AdxnTMEzvNd5h3wic1cZVm979ch7pCIUIB4oRIt4UTwQ/R5zInGYZMV
4cOhhAHbIYuQYO937iVpmWZJDEVMNb1d0kNmQJJ3W2lT35vmI+S0QoPhehfs
f/v5aPux6f9OlH6tNEh7bXVyvX+iDcoWUQwT8UdRCDwV7ZM9YvX+k1b0KV5+
5abP3VjANSLyRrvXhx1vTBkMKjrUEXjaya0QNEMivKRPNt0HNGwYxHIexFzN
IpTTjuuMVmTvD3LYmi9KRYxwSf2L8Ww8MdA7iGZZymjCARJXc5rnbZVfJmNL
3OiGxTBUnNarrh/78oe/KzgAuAR8C3nkP1+Q6laXvjE3xv2Ox7oedZv4uAbz
4DiJZQnSsgUdYI6ncB7t2bAM1vRX5iIVlRwdrLn+M2rwFV5OHPxsq9b8lxos
9HrFkz4Nlwk8H8oLgQxIfFyAChrvFh/R5NaFjaSwkXAwZeOawzBtTgK/CKME
bIAjm6UqG7ThFIPzZapJlB+R3rSUgKdziIhsEQWr3pPnssUN06XcXAI285b2
gjOviWOt+hZ9CFoe8zklQ3NVBT3xXOIrBAyvlB2ePwAUwhZkSroP4eQygHGN
yAEnjUfPclcfS2sbyEYMvFQT3uXwyQ9UiGnmhuofnmMZow5EZ+j31HZ8cTE/
IkXxp+SWYzMwpGBL+et9CnugFiN+bDr1zfR7tbld0j3UqSaV9I+nkVJuIAkd
c/ArQvaSZBlXDsA3u5rK7eHR7mSwZG5J2vC97rLQQKN4SMjU+NSmbGwmn2qV
yZE1i1OLXDRIxj22m+O1Zh4TgcfdFid4NKQz+OY1wP+hbIkm9FCr/f8ZrsH6
fgb9mT/gp4eEzF+OyLowyF03BaOxs4Sf2ohZ4EvcrceYMU8D42+aM1DjxGSK
W2i/0AknqHzm4By0e5dQusRku8BtDzTJ3CgDGbQjZe9zBjV3n4goY8X9XdP5
qj5fd4RzNMuzgqhHJLRU/QFWgcvm1v9zNtg+BtRVAoz3BiG+VIBYGCLuvhI0
RQXkfcbZPpyjq5Oe14dWkz+AJiyiqh8cTC6BOKKpBFz1+SV73+Y7Dtu3gPB1
hgjNJCbHh1lSlVXLrvh/tLFU53BdNPaH44mNQCep7/bTg9iHIGAqIqp/Ryf7
CKIG5+mkuOTWZIiR3xhaWPfVQR/xuqwyORwxb2rP5wJIyKoP3BPy5ooBPvoN
XyYdbaEWyX5jpM+YRekk0zmFVu02iDufSoSsLaER2TNhtNmoZuHsSwxjVA2R
/o3ix/hwKBAEQR24pMCVqL/i8xjP1Y1imwy5VvageUkuQl1Y2Kdf0msxjFCX
TtlRrYC0mmFtGqgL2ChU0vdMZ9EOJ/ZiZkbjvZjPnnvBNEDjvq2jtlAttMGK
Hc3fx4Oz1BoOEMqAcdxjFBqjCUveTKSTKdkophUok30Zgz+avimAIZn6qz3D
25mO40aigv/HUElBor/tFgG2NmkfYu1YSrhhsPZTu0GPcyBf8svWgTySB5Jq
XujxqCrSQD2M71mWL5DBNWInjSusaOsatFyjmEi9RIOFCZKiWPn+x7PJiTaX
O+lBeco2OQxV0fGQ7BXN/RvcygdM1lHpH7lt1QbqcQJgVUuHeim7cXLk0XQG
PCWwWfYzlaXqHnsTkdkuTiIuiQkr6RPptM27OrZx5jMeoXayew6aXJGEn57P
L5GinOFZWkQ3tOiAY/2uVzdOd0YHhrewAw2klK1eNq+yP5CmlqZIy11XErS1
ogn/A8oGEruy31DLzx5RZ4iIDR+yj8x7qxBZjw3OE6IJLROhDGzq+V8DAz38
zp1oTjavUj2svfzwrfZIIrCBtKzSCw73rvF0RBgOajG4RmKQLmaH6fP7SyTU
lbxt24f3xXgHJn7r03ZP5HPRcqiFL3/3MeVJNfdIRoonLCLP6zVbTcDi/78C
8TKvIHT+47vfoJFt0B0Ltxb2m5fXj6gPvGeHJhhw2kcqJU93vZGMfa16pZ+W
lulTcqegzvk+XuvW3FQ7hD1A0CAsOlqNu+C8mfhG4iTxFWpDZRjkzG7z62dA
QKU6AmMnot99PZVd+/T+Yxpg2QURodGvgZcBHFsrZPJvlIeRUqIiyii5eEH2
b1Ppn7xaW4yVzsRYG67A3WkMz3GEtcFhFZgzLk2fJuO5M2zzQg8Ypy81Ykct
HrgM2x0LSzIlCyGsUOmy/ttvJUdaOSEqK/mdoCTdPDZ15zEUQFbQlU1AbB1Z
DOqLqEJn7ShzQhpYWADe9xgBIaFtWjhBtTu5FfKfE5arsDRN2tYXphtGQ7Cc
sGTmky+OIIqfr9gNDuojgf/fJYwt5lR/in5w/fXMtgehxtx/DL/T0mgeRjy8
WNkV4WQ4FUFrmzJJgBmcoaqzOdqH8hp/WUMWinUlf5VzB1FEL0Hnvvc/tuDv
MrxUPx2Ju8vjLDth11LRn+011ZJQoqYNb8NVlPbxlA/wPhDwz2z+DX+AT/Jh
py+NqpZYvz961/oWmDdpsPhneSSgTOY9ymh6prfPqItxyyOgjkoOIi50CT0P
BjjqY+6Id/p+TgtapEGuUIqmjYBYovusu6RHa6ZS4n7eH3ZgRiotsbhL1xTY
4BL3y9s6C5+Yb29WaAchWdRQV3NLGe6v8BxivXmQ4T1LKT9mRpH5WoK3aQ/O
iJ++HZdk9nAMsfiNXg20G49W4O1OBX+rJ2iwgsAEH2n+pHySQzKBC1I/O/hP
GKqioDQRUrNzQmDN4jZ04K4miRtthfhfTPK8zMOeplC+0Yx65aNzfM/GjT7m
pK0v3AUtaKYY/xBHMO+ffXJZ3OGFjl7Fse45f9merP+Q0zYSqUZz//3pKvTJ
g/kNwgpMlJgPNDGckxB9GUvU/zUTTNOi1hBxW5Ok7ER+Fhq97r7cHuI/rAlz
c0tRpQNRA8ttdWXBwK+/cv/7KhtHtbpLc9y779//ryZHb1XERX18I7S4vgA/
e0GxV9qLGdbtThOEDcO0IZTk75QpvDEQqD+DtHz/Ty1kBd2m4NFXkWsVng/m
1mSwfml21IshpbRA5ObokR8GoxFbRNhTpwH+TttDMXW32hrGPmCJeEVnn6nD
cit9HYaZA5oVV1eq1miYRrDEfWUsYIMTE3NxovMZnrof9Y44bA1LoZva4ZZ/
+lFj6GJmvWd+qU3pwimSg/mOQRzW0ga8WuNdKEbrGaSzpo0Q7m0q/tw9DP1e
WwyGilafZ+goo+g2KhZEt1atnvk88hwcxmZhYLhAwqpLHSoMBi1g4SqC1Pjy
xj0si+prWz3jbcR+l15wso5wCUkS+Lup47yuLvio+/zmombtkQvAiCCUgVSQ
bnTL9/DE+NSfWp36MAfS7uF+EeoYAUujz0wMOCJna0GMvdeI/UfabeVvH6im
mpVqW/cPlX2MyrY21jyohQAY6730jXMsp0u3//wPFbHSm8qQZl0lfWS4MDEZ
0t88bN0Yl2eoeC6UTOJgyeo+s8G7xQJ01IUaf4pVBlgauCA0V8hjaCR4nAhw
tbwa3k4kuF27E0gHB6GQMDzsaxdWzv6kj4T+7jDvU9eyWea/tLWhQxeBYHVR
LrWS09mpt+IAMA17GbQcqSwMV5evMq4jnn4e+zb+nn19+tRW2lF5Wpzlg6+8
B9I1loMb57a+wlVCjU1RfVtiROoE4DAXtKkptBXfqed7MHgxZOQ1wffhpuVj
+XAOJEmHdlOHbFyd54Krje9jBwTpdpAMSmw6lA4NGeLihbXAbUFEgsbzdSHb
GZESMUM3bDQaRszpe1Nct6NmS42xP92FxWlS9EPeNhM5WBsSIANzyAFuCS53
hnaqh4Y13Ug6iaz6P6xokVP0bfXZryEatsVe5m2MtmuWS7fjhhSBTB5IaCY9
YS6Vt/w/LWFV1dGs2NmKT54lvAq1M5jX+18ncBPtDtqT8G8y8UI152KpdJVU
+xtllGlZE1D06QeRJlzIpnmUW6B8dnS0gKTEpHZYZtkbBJOdvzvLj2kwDKRu
QoNSf3Nxl8Y8XC6BmrYIE3GWNUifIeDmuM4MT++RblHE8CCTrVezPutGDH3y
fMugNIONx3WTGbUf4osqRA7ZJNiaGT8rmyPi5wWR0hqQHaolbKuLxB/XZfvy
VfdIJBMJu8ABGTjjqm6BexhVDyYlNVDliF4zXK+8sM9N0VSvRspTVJGT4kSI
/SpwrBWfsmW48E1z1Ov4G0Ze8FJX6olJDo2M+RXA42E3xK9dCKWsqElcmJQ3
oa7sMaoB2b8T3nnRhOxtfg6xqHJVc7XWfkEMEqSqswqrXQC8pilXxU4hsUXp
sN6D2o6Tz6AfW0ZEVZ1ySvR4W3Em+z9GdUMYX4BmovJ0jqDaNUSRIzWcPbua
n1w8l47xRaNEXA2sp8EJ45w5U4qewyEdHKEhPwfAx17UqRUifT7hPHAjSlOm
6VmYGGLAtIWs020BdPKb4T4UmyYmV9hz3Xm6Y3ETzBYv2NWN9PHipUldy11n
NADt2Fn0hbyzqxYLceXtjXzo26QNyH4Jk+fgtjArmYfwIkN3FrUoqeKDoG0D
5tSoxHKLototnEE4UINux/MnECswGN4yVLtGtKeaqnE+ch22iDt89GJQlNaW
+nq+Mqjl5Rmu3RENSlkl1WwVNNAmw95YzU9VWrof4iZVVeMKZHs6Na9DJ91x
0dbvPJ2fpFrw2v1bL5RHu9sCk1bjV7Nsfq/HF/Lh4z6/S5aOcWF/L+loOvwg
tHCJXujH+/Uxl64kBPcwpW7DIQ93tpoa5ACOmyLH78YZN04o3V7XekKCSITz
h66anRq21RsTrrW2nJg3fyp2ylkDPVRoG+GEAVqBkxsLfnPWMUWj4nM8fjna
R8D1wxmpLCtObYBc+aaPfR0Pi863sjRhpBvsguVZ00BtYRNr/qINtqo5nHQK
dQ1k9p6V/2v9EiXBGfNbkRxSix7yarYIHGK5e7bl+ZM9P4CRQuiweCEGiLH4
KH5LWEZuIRc7ecNIB0YxeiWOcTecAqfKe/Fd+6MdwbUTFSdxEBmu3aRc+MSX
779u55GDNdrsBBZcymZxHGCQEBK8SM4KAcsaAzzetzZkgQZ8NIxCLA3W6qtf
j1c8rYpgQZTJplXvaVGYx9+27+gYdVP45FFI9MqP4PzVKellF8CZB/EM3RgX
FGk41Le4EfErP0FeHtNNl6fFqZUULFLMFSS5+qKI0vih4ywjUqE8zYT1WJOO
JwWvhbKCMBMTAZ6ODdbwrF7b582rhE8PRmHwXhBQMpfSTVOwiVf+MVJJV1XO
w0GwKsZi447RSHgj81RJ58vBSq+VVJGb5hudfTORq5p4UPO4R0i89EiDtjSd
EiRqORlAewcJH8NuD/gWAlPudiiV+PGf1znl+2WkkzTOWLXhW8gjZDStkK6m
4SAMyYT7g8M2yLjKzUmR03mQHptJ2sNzPdAnDuYyAcZKeEAnxJAP2REf5q5W
Kkn/KzScwYdPWdd3lGKScDqAdfDd4RMvXW3u2xcM6iiSy6kf6dhcndAu2Wc6
0xI+JbaR48zTeEw2kDg1SzWdDANYQJpTYuSoEUcJee525rfbKLAyYRPWlQnR
q3IsbKWi4Xh6orPWrcIurZaAt7w67jXQwUoYQ83SY/vZNVap/eY33EpfEP9B
VNSKCLKPLwwJATstG91P5FESXRNbfgXASMBuN+FrtdBwk41bSiQPbTp7/2Ij
9lY4RC2ALIimMXL+hzQtDUUbndTCujHLA3DSyyRCh01kNDAF8mcPgTK2Gqnx
3sllPnc3NoIS3ytxoxyNZ6HPpKHiKl7a2X1lVvTAS9d6nS8jpsZy2Ry0xuyL
mGszQsnQ1hUJT+oRiZjaKiTSa11ce4Rmc/wU8EiIz8vVeRphefEBUgxVpDPE
tO/SUyCAprrGQHMcCX37nK+ODRtWplEsmWzx12wN2VaQa+JEt+Il9eH6YAGU
tR2KWOYywz8N/W0BEIjkakV/imC5RoWNognpy9OEAvtAtM/tCzhdVak5GK0V
A5He07jjiIxEN66k/eV2BkvEJbaRY+mxtqcMYGp3Y4SjL4ICtzwrju4z89rh
9i7Tghay4xRbRol7xAxqMl5r9IS6zPvRnXD9LGfgQJfQXEchnQAITKkJNvqC
+0QzcvJ1JDjs8Rpa8BJ8+iPX3eUESn1vGxc8yXxkRoUbfpr8WdDsigbk7Wri
gG1VB6AmUSEWQuwh24vO0ZHkiEADqb+IAnZ6pnqIn0GJZhqvtQZ/gav7y/HM
L6aoMl7vcBXEYm5rhJl2atDThekYTg5jDdzjRUuJOHRsD1aOvVNWVwg4lD1l
pC62Wi1EDZ9TuQq20LoBmJO6uzPUW46BcMM02vwmcjnta5h4QGQ/g+d/RAON
djetIZ7R/woYROzaR4nw2t2vo926AAKCkvtvaQXrzJCzbjAfMZpPiJb+RyNn
sEzJlZGNYKy5o96bzz4ulsYiAY5yL7bGW/S3jLI4D1tuVI4KBVZf8HPYyPMa
IcljcA+O4KZnZgYB3rSjyNS0ke1pBEdFbQFXNN6VEOmpxkr2vvFkhYIAoyQl
7YmydbCGZgpBkGDyGn9FyWd8in3cLbbRX6K71w+uUVrD3xNfSIARXzf1SLuh
erhwouujFBkpyPef6H37HP3DZ0e6ZS5q07eatF6eiyWRoIjEMLQOp16KnQbX
VcfoedjZgLypqDxTOdwJLqQY0heY8DK3LxtKuXeIRI/QXOsE2xMtG5VMMMGl
LnjccI7u6Z3Ape2YNFv94WmPL5oKU8wtqas4XRGU91bbY1cVM6BnRZqN/J0u
ZoEVNess9XClS3j7Ren71U68kCdCmwsND/0DpwV7WtHEG8BPQQX8+XQH5Oo1
SVpdhcSEdO0LlnxRhn1pwiEcMwHBDYr3kpTeZL/SVBzUC9L+8KdSYIhrcl0M
s9FBV5UT/fUuKutvI25n3lmE46n+YoKOXnvl1MJjRmkhek3sE2yR0kSneZpJ
PIchc0kpZYhyJvmgw48UFh7IB6FOTRQihhDMsFAQHM8V0SXsTZ9Y9+E+QGvc
+06UGlGZrFPZHUn/2OChzulOj51NJjS6rjaFqViTEnw73qXHay0Ng+ZHtFk8
N5FIltK+dIadmEqbg3MxcnKZI3sNTuPqrKIaeplg9zHKv10XCp5+Xtvuh4r4
B8SoNh4mb1LgiUvuIgK/IPsFgBP1ZsEUugLSHj2eb6OVLt/kiHMML+P3kNvw
A6UXvQxIDI0sKoqQ0dIoc08BWL+/uhO5ZtW8WxSBDl8GzQgFpQJZQQ27HgKc
WaeyHBBJbTOdUePCMs0NE1j4S35VECmd82Q2cn7nWaFJsrOSe55B7TZhSt8k
iXxnTVD2wp5fkxGz/gBXoNDyIAkpUvSs3CqYNcH1nELDeIzjANb/u378SByK
etWgKrE8DN4fEGr9ehRZOaYUsUxFrxJOk5aO9CKt50ZDUPyofdWNYJRwbBDD
dFnL8WOzd7toxMEQhvjwx6JpT+x8QHPTTxA4M4iXGEaf9Z8n+KuK+SxfJdHm
v0tK+mk0tLSimHXHostRDpIdg84HRzzmkM6I5k30LVvqf3QCKKLU8GSihOvb
JSDlZIsBXk8yKFveLMzIV5K0AHdA2caOxzREBVcWHI/p6Sw2cKXnDlF4m5id
l/Sk7SBLtnONV8+T2gvYLzkiX472hjTqMxz0MZtpyXl+MtGwagOLA1XjsF5d
qS8BdYJxL+QAq+4kD+dCrndzIWI9nALLzr4qqgDXW+WhIc0sEMNJtCtJJicu
MWS170AetqMiPUNKjGqFzYDbrNCJexLOp8nsKEgTLlUlkoteamG4uOO+OarE
lKgUmL2kaMfDl6OtTuBdaXAYX61uqYUcOJRYq5gzG7h0le4uZ/EHZHQi8p9y
gdU3b0nuITWnUgnuv90abYn/Y3+5oZ8jTNAx04sx72P3WUmRkxafu6a32U/P
SMpMJ1xSKY7Oy9EmigwdWDjvpgyf4IusdA3888ExNvp2bf8rgUxkV+yqloKz
DoY++o98jPcm1+8rXk5nv1qPwmDsReFtsZ4LbwRDi9R3l7oy7cMPMCZVpqje
9O+v73pjZdoID4Gxh+GlkeK1ZmQrH74xwc4/O8b8OepOLe49rpgWpShZoltD
8UzArxraQvON0ev4aA2TPd0tiPm6eAtV8TYrgjZuabA7g+mDqeiGTGP5Hp4K
Zy5v/POg6eEpTe9kVQuyUKLCK72LfKaBPU8a46qJ3MjvhjDpjR7i2UqM82n/
sp7POaoC9ENSA0C+4Kmg/t1Ch32spDsue4R5Dh01A76K3FyeBYszyTznWljf
0c0D/gF9Qkp7T+Jic4oaOkRZZO3lsj31doOi84TJwyfIy9FGEXf20WWvfukx
ZQBsDSsrA1hER9WcWHMQXGx6HBGXM1yWK3tTv+XRWtJd1q8J125pAuOC5Q5G
B9ANWNo+AuUSQv9VyN0CoIsarhbIGyFG8EDoNKGQZQpDxM/i9axa3o5YPYg7
k35qYGYNd5jZ+E49EqPuYthNKbEkDIaaWVEosWf/hI0hTx8bPVb//fI+joZb
02rS8Na+2rf4+r8HOcNTvrg16PZe6W9P+T9O2ZqYS76QNENhAIJrS4uwHzzQ
o+IscGtbu53Bx//qNZAvzuu2N7WV4aZqmZQt/i9uPZsFWbIKZOTzyphdxgFa
jzIJUETuUrZAMvu4JXigKI0bpFz+98rJ5MFK9eO2OutbsuPedHkcyfDJCTxb
uaLtXs3WwQfSKbQHzL0ks8J94fhmifB+thZaggzqnqVBgp3BA/QowJNgCVum
eshkfknqAlU5IuhSLqfJJyhtS62ehK8g3gKVLOE4q8cCIoxnxQBtWIOqmZQG
Rusc1CFDdrCYiT3ts8ro4U8ZM9OBsKajBS/ClGiuVZmtWsOtW47hyBi00yWW
Ru+2ckcV1FFK/bzNKtpNGICHVV4BW8yF/VMHwbDgodOkBiKxsEyDPFzcAvUP
ff7t+m8R3b5FuIwn91U7wB81yU7TCjBGA9NVCvJzJtkSob4Ae50eSWPoVIkq
XN9PDwAc3QjrSvI+zW63LIiNA7crW9GsgwwpWRUdWPsjuU6HNGZJ1j0I1Lay
q3PJLhYxVLNqQmp7F0twZl9HQImDKosH0HBvcFNbNlPWWe6Cpdq+4OARDwuN
8YCW1SFWSYDxOXbSnmDRK00BkLibGbT8CkNQH0CzG9LPFK6SH4e1e2qG3SK7
tVvb11yjvt7eogXlIfx+61LJJDW5fROWGrmZpcXz1Vwgcl0ivMfMdQDfIFeJ
SOCuhsY6Lu/wowsaepG1URj8V9mJ2WkShnky0qQMXw9uCb77T3poiWsJ/gAr
r2EjMz1Azdv4p9Q2y+PLn0pVb+0fbNkAtYvYtfltDugWdE9ws+toxyKZ0P0V
M4ErUPDcX1XYXP91ZnQNLoNPW60hKaiAxmvGVUH9udQ3P+uKdwTrPbrBi8bT
26f9P2VL/FpGoH4XzdqGIZ3LD6m41INbRNbqLs4RG/+1duYEDa/nu/vZ0wLP
mDa91fvemeC28yL1EI+mHa3C1HcYjcuy2ZxXH5TCY0CUBV3STWnAelmjp5cO
MSwO2oI11dpj1Ex9YhHNA585ZRSugspy5p6HnumSr3w1QgQnCTUh7fg9oWyG
E2URdwgNuQVR+tO8tywyWHsxoQR+q+Hw7qynAhuE68IMEa7FnjJQ7UTHlXJC
+YYGSiji+Xa8vUPs0DAwFy8gC5323JaPqVMWWyCrqRMVPOcLYwdvVjk6+1ur
iULbacd6W6hZrMDMGGpS1NsSjuNp5unjftsPEV0REgx62jlR2KKiRckhiwwP
FuetAQfDltb+c6biTvwTe4Ucrp/JoeTXn5oAfnKtAOAfPuyso0JjWBDQfik6
2x/OWAgAIxf4ceTCrHrA8shc80pfu+G2WgqMb5rv3w8mEQPdG/yMkvwjJcUM
nhmqJe3Pb1x1Vp0QOissGjq6zDy3IiXuM/KoClX9/fkFbvMzbljq05W0p4FH
Yrjdo8a6k+jNQ1YWyvG0Mh0R4Db3U86+7aqhoimVd3OW/K92XEEMFFkqFBxl
3I42ttqagpxmJAjJ1F0kVELiAyW8w71qvxUsfhsPn2pam0favRMTPOh2C8BJ
C6qv0p5uFouaTws03cwuKP/WSItZoUmAuuePyINOLRsqWOkR5fI4yTP+c89k
D79Crb2RR13S4NCoSqUedY1q2co2IuO2tuP/MEstIY6yjSJVj7Yz7bulgoKr
hvfTDAjwjAjpcdVYK45CMHWy9w9k5L6wlfLjwLFqMPj0UOTG4fqBQG0Kz4Bv
9CFC0hGzZ5ZLKgKpSmjOklMcbjbjXwbNfB906uDoc/jqptiI8G1R6X8LPS9r
lwlIP/aptNz5wlnYDEN5cQT0J57xSe87F2Evx9tvqYQpuOVXg0p9bMvRMl+5
/axahvv++6vvQv16GSGzCYZPiCw+1lms8NLLaMUJ3qe+S9DuSOcrFeBV7dbF
xsKjts4F5dbtKEEOJw4KdYbshT0PTj5mIy7jmlneV73Qohp1dcZqzmWqpV9Z
7h3+FHuZPETKMcLlKrXao0qqPx3FJG7OOpcpY3fWohIIer3sHB/+LxNZ632l
S/IOOiH2XtLcpeSazKnnRiRtrPlUrznmcaTlXznq8Eh/d7vSz8iLmZQekewl
5fz3NXkp46lPK2lKpMfTcKPYccy/EX8JpqU3Mt2CizuWrn1+jI9d4q3V/PZU
+3VGIS2x2sFWOKNxP/Hu7cV2Aik0mNVk4pki98jLccwlKQacqq0EdWtbV2s5
oDneLKvokUChJqh8YNqVUwkKMCzQ/2sVPIjWAtrj7HQ73NkmNpRdaMnnDoJ9
wFR0xlXPfv0TDx/IXR1pHIcouQ5saUgoMeCmq84nT6/eKc6HQoXuTeBJKobg
YXbr0oF8a9ijXrtwJwg5059rhTb9y/TuyIFxDtOVd8Sgzy+G247qE+tEEehZ
pfgihNxy0LGgcLvErE/BBbZbQCvRJ91hAnlxFCc1HyNucWyJOHFpDVs2papx
48nfbHsG9GRaMPp31VFGlZgw0PXaaF0y9rX6i6oJvPQiEUVM86mDmZSBanp+
2uENIDIU9WFOxuOveU9gt0Puo6Q0xjte0UHaaE0BZRQtFv0mDNr4jR4GPpsw
xZA/VvvlNe4/Z54gi8x3neNbJ5ZTNfJ15kpAHDwJxtRe9YY2psjLANZyJGsv
MvCVd41M6pMs688QIIhBDoOG1BwbYUm15QAQgxT2h5mtEe/lhaGQit0uZEu6
YenRE3YIPF+1Hj8GiTgTGtSXqhwz48g30zUszl9gXVa8j1i0sl82oFR7X8i+
KAmqYFSaTagzuhEieTPV6cpstMYIrANYmeQ+Imecz8GvQeBgjY50UTxc7g2F
wL0pKW1hGwbkdBbS5RuetbHG2SliwiTx4MH0W2eCsA5G4p9QAc22bC2PhiWz
MRfizX4JXPKgeyk2aERqNN94Y7TrJDQHAWVt7Wk135RX3t70lCAW4ABnHmm1
As4mEW/AuQ2XCqbdHsjUhivx2vLyaAHKtAqZJPobz8fulZwyhUnkIOccdYX2
+zj+ftrxQRhz075NhEEqb4+QMbfaM1vogQIyI24hiPVkqMaU5atjz7Q+jg+s
DKRzQG5mcikDX4hOjpmSiwboFxaSokt3pgUPyMKSUTWj0OW6cpW6lgpPvRrD
HTpt4cLMjT8BG6wqklEt6qy3Si5GiPH8sSrZCYsTStPpy5+iPh31BFgvN4e/
H3dUTDGgbBpYr9bgtcIDj/Ea2jNbkh0/f+PZ3srk4k1juQeAqeAHat4I39eX
NiCftcjbttmj2APPHEiTYBRnzB2WoU3w5jJHS88eSWbsoYItYxkaVVzJQXt4
TMX7ggdwTInvV8iduzW+hFxmYPxvkdjf6/cWxQwmxodT2qC4fenCBjoDujGi
SLtjY16epJ1Y6MfipT3sHHvqdo8o5gxw+kInYI6XuURytpe5KFWPbPMAK057
VAP7JIoNdGzZVQI+iRV1dS60juyjyAf17m5m4zJYUOmVF40NU+MxqKfb8BUd
DDgPkLupKQ+XFSNmg5BJGdKYJCb5LW91HVk82b20vdBeBKbeCi8BUqozziEC
lOpHy1XdqTtmY7vRsGlQsUUovgAuGJ5w/xPEz3+8S25T38Tes8RBjm88LEtd
MPwRcKK24tcL5NaNFoAGweGCAAFUw7kK493YcErdcymZn0b37h1jGQjj7OTv
jNZKeQuOVIyUPjvA4uspxEJOAx2DbQNDpZifYC1jqH4QOVccEUzFyuujtHvw
U7QAy5hwuYNLyqSsTl+XZ0sINfPdsdivfD4SBocolmys1nI/RDt2t1ekgS9k
wQ2SRGSGE022UTfgCy7HLhki8Z6OC8kExwxy9sv7UWhZqgsSgTDTZZ2AAeNI
qMfktdAWG+9LdyCxGtBv4cezgc4kX94A0kCNrL0IfeT5/PlYeIUMJWfzNbNV
YC19Gi4Va9Bga/9cUUshFvYSCppsEb29JWkXYQNAgWwAi+QweuqDLE6n9yYB
FlnE55BTHbvX6Cjj6vUjn++1YOizV/lwFnKd62ecdXLt6ZU0ij88Khqzo4vV
+60VKoj6tYEHlRxCRJ7fsaF9zh5eTbq3V3sVSUa9IzoeekAPwPApKQ4RxkyR
1kAroQH2T+DwBahKnSGlwW8NTUHwKLUNO8PT3Vb8yvC5vwX59eR3ftdrOBGy
YbtxSM2nUq68N5WPbuqC9aTyty26MH1GJ7e4Hhsuw0vut49FHYKJJp4kdOln
qBPvT/l8+SjQ/s4YuDAGED+7DmkNCyQTeaYOVllFAAFnr35sCeKAqt4mgiKz
7T0ou6J7nhC0XTMhLdO9oev365/kPOsmOmkMAG0OAUowMu7F4ts3suD5dkxS
vpnOAHC3/dFmL9og418KBlWgl0TuUzU/5lK5nOTLgwGwhU2hDbZmbVCRGNXp
wWd6maq8GkvUlVXPwJXp3C348S9BsuA1LAS4GBQANtcUH9Rt+7iTNNqr6uWG
DCwBZyrgsXiePIG6hD5vvMYA4sTgjPNBb20BcYCvghNhC9BQ599vVGlzbX2Z
JF9bll9Qr76bnsYXlMgMuUyEiZ+3HOm8/T2HBU73SkMXwnK+a+mks9RXVpmc
7ksKH5Qz8XY8Rj2S0SyO7NkOIvseCbmgxIAPSC3yY0+2it9KwKaGVbSwN+Wg
PcVFu2q5YifEUZzoRtMDgrmrZpx5V+XcE3Wl7xD4HCHjsBUuDurNYsnkxgPj
4YMWXK2m6hTKzSaRM0qgMGklZQHH/YZcDdAdBLVsh5vHBYVVHxdCwniF65Es
q0Z6svGuwKVG4GeCSnd+AjR86r3sW1dZ+3v/LV53XeuVWAhQxYzjhRCfvGlS
D2LjpIupJBuGA/fKj46oSy4+utHPo7oHTG0liZEy9E7oVagQCU16VL9wx4n4
xwAOiZZKef4UXqFg3A+I8jBSJ7GA4+Jn14is5CCpIRj2er9hQmBq4qZtubEm
d0SHOAX2b/hS230t4ALAGjkfNIgA/p/G7jnD9wstrLt+n7ZloQwsgSAlYB3y
rl2Ux3pYXUY/+HgQetiHRboBpTpqbcGg0DX0ncs9XlJ/7i8rehI1C8/JVmlg
pF8pnM2dGfIB6YztlviB7bwHyuPHqLWwk3IOo48czCfmVeiHra6HaaScfDBO
o2jjLPYh+xOIHVuD1wZhPzcR4DxTt2uGzEfUWmGhZ6tX9e06STQkEqJvlBvW
R1VVxV/Hnj6fmbx0bZLbjjk337HL0r1ryMptmP4JHsb2Nua+7i4DKDvtQBPf
ZS78QSQtfiIABpnqhkx7SYv+hS5U3hOICRH0msytgh6R7+F/Q+gYkOMrh2tk
nvZ9YXpyjv2Npx8dwVrrht83IiPUgFa/7vhTvpmumlpuWBuXo6rd61N7aIvS
LlU+jHYQZt0yChOTxi6x5MRnZQPcXt932LJuj7C7Waux8MUC2kDcW0PB6UEd
I4aJsiPHv2FN85TCKv84RTP6veP3f8IsJCANduTa3lqoAZiX7IE+e89dD3kN
rxvPFQE9BOBVj57SsK0xpTZBpJTFzzSSGrNfDKJBDosdyoQmMVkTT2gXOXBi
vGZ92OtszZfuoBY2ab+avIctH7qQvkBK2lFyUQAs/6bJqS8y+ZPpfbqLqv2s
8Tz/tvAjXZOl6tqP1jOSicjN64oy46tlFhBjInrzIHO4uzZ+9psGcQUdObi7
v72SwyPHR9mUDGfJT8qyv17Tx4uijILj04I6tnSy5YzQZKiDQ4wYAa8U6X/5
YGVCuiGQEdt1Kcad4UHRnBS1YHVo2GFG45goCo1Oxl1jEq0hA7usoRU+bCRx
N4/+TccUa0XhBNOECTLr86zJ7abD93kaSyltPBkNDmqiZ04o8koznnBB8jH/
Co0gff2v4004fpa1B9W0TOy79pLR5nJV+5uGDjK7Jtt1sSd3oadmA6foYmx0
2ja1NZtMl6OOpVbQeRBGysWp3wPL3RfXIM/KUcTqzRoswKzFPPq67cpNzqvm
xuroEVgFzR7XDwcDHs5wX5bO/gSnig3jt1rH0RofCRfr+EXbnU51/FAflgVi
+r0gbcsL0HjowpHSWWrec59PToQji8nZw1czz8O3T2jO3wTGEt+OaZBQaxUz
G7zBrviwCs6gbn9MoO8CYzUTjhS8607FT/1S3cGaXvcpkWoj7oagamzh378/
CVx84LK5EVYxzDQyiqHXJQ2U5fj2yJH6QiNT+lZKpGTbcVlCa4ZfeGUFwtJy
Ca87hVKL94rHPcPIhAjJMTtWBHHB+yf4ROIQzkP1MeNCJfLTl2TdRPMh7o3y
T3qHqULmR1oeclYMokgKaklNmbWzz5DWb4f6KbU2DdI5lVWlLUROgjKPaxjz
OWZ3inu6tuRpjYOI3ycNMdRhpy5WXRTPXUV9qd6OmXqz6fsykZ6HXA8J36nO
GAOM7ihpCl9KLjvW8yHNDgGAxdP011AhZaPX6PNWhy+6gOnBwcre5Zo0FxkC
qHdYNMt3l5RR4lh1J2n2UYTFV5clYnf7Df8N3Y6TDCPKkaWEbrYV3E6ULw9X
UCozbJyg5nVry2Q29AfpkJbqFg8OmWo4QNsgJZo73GWyT9G6LgHdEoZ5qvfC
39GHuxm5ams3gaTOIv2OGHRJcKOdZ/6GDD+jdf1SxnBasJNjVRdYsRO/ilm5
Qbe0FF1QIFF03sKDYjuP3B27AA4i4YjCQxdm6YBnQ7LlyyMKmkvW9dFv0HGb
xjLqTuUBp+ggMZrSwcZ2JIt/QdYzZnYhi/GDUy+d1bLXV/gGRvkQOoEDJvCV
utTxoozVP0FfuKfgKoySU6WPo64yDCTrEP+zBfea3m3wiYTD2EDUrI6f1Pid
XmYKerFUcdmwvREI7I8y9+fnKts7yDdfDAR0WxHoCli+7cggwiuO7bhs5Dhx
sKHve7Ms1f1OqgR0fyKrNXL/ggQsSVCD5QjMucMfKMN++gH85CNks4bL0aSM
b97226ztQcVODbRMYG9Np1L5KB04AxmR6YGERsp8HINkNziQaRKtvR2sMkhz
4TSbCaXOXLCc1ZosuiC1Whn1c/OipeD6vlo+uVkfQebzb5ViKu0Hk2ijTr4X
LvKzqIVnFNitxAMQ3v/kbtSDtQTV2S6ds77KnNqRBGeD42wBBfElUZUj7FFG
gMBsEw2Q3dBJEkCYTQhhz0c6cA6SEHAx2krdLZ0CZJnqVAjHurszlb2I1euz
PE4033CVHCFlFZkee8IxWDvy/yHHpfkUh1o0vdGOb8Wo4wAzqJ+4uChP9IG0
EjPFDDJA6z357de5I5tVG0l0bxIH9Nm1v/xCuPxLrYMCS8At4ONUkoae/Q0l
Ga+qcK6PhBR/Od6Cvl0orkjDideoudTmMyUQsvC6vWC8BSOp/EtKXdFmkv9S
Ek8ytyZcyWKvDnccSqfVU8S7uC9CTEXA7XAIuEzT3p8OSchbYfzOmljo9Mgd
pU2RTjrtXvqoJUchIcuTIE3Pv9qXBUJhLOv3Pa1zkJVGObf4AxmuiM+APOvd
8Nj6LIZDzs1AtFObgXdbrT/8+fgnTNmAvQd+zbpBOGPXZpLGio3aEb2RTD0y
K0yqFk4AYaw9XWQePFcRkaeMyPhTstcBbsLwOK2pu20H+Jjf8mdHfp/kLsfj
0T2/UzBbO/iNQI4TyEE65dj5kp76eO4yK1M7vbknZOb3zpkeFgcfrKrYFCjv
n2DJY1gUxTrP2N+NNSLizRfpRiukZwJabkvzEATQ8LwvWzbwXLjQh6S5Uaj+
/1aVHqOYxYmvBKehLGvpCz7CiMFaee87TqhWTySrHQUuioigJnzpikYaoG7u
fLkfSG23bLn2ur9aB3wvyzUpfWOoMhm9qcudfeC4v5AsC9hpaXfRk8RjfuD1
aW3mSD8rZYlkArNNmoEDoRS9oTmL1ohXCfQq0nAMaCD/uwVYL6lv8hcn/s1A
nZEGAK71F7n+Hc30yM/hiVGlXDmNRoXBC9592Cu3TVovg6Fh8UHMoTGVrrBI
396SYq2bVTQnDKOwJ+fhlzfhImzuWznpwVAypx5mvFcInFUR+CT7NBdzkQhI
XyzMQmQ832ulURkI4mS5acC0cvVOMU0dJ5PTA9OJSJC2N4cPEe61QPivs9Rc
Bo2ncL6AhZLqimCKdfNaNHp/6eBtx0G9MSaKTlqeWT57bmITG+SbVjdo1mI8
tv0Oa5U6ZFRLSHTx7w0Dai6XEzzL1Phx5uIWMKVKSVX4xVP9z9zS7LmQaMN4
9llIAMy9evYX+8ZrMmoRuorMLM9dacAQyHmen7Utk2GOqh3vvgeviYnJCZ/t
5C5MSrezphxrHDV+pQaOT36fFCRpJ+Q3HmB41SvVcWs6DNmzNhV2O/pHQ4EZ
e7DPB5fx9xhbDrg2QzxZyajHXW0Z9Ix4IggDm7hP8Pde/O/cyFIylQ9fdyJk
LK7Voi+yhXg2/DAsMPCDZHTStr/x9l1NvyE/n5AyJNku7ONiU4m3AhEhbA1E
onTFCLteGfyVccIwOF0pNcGz625qg02FP9SYs+yy5XnkjqLAsjJdC9bqgtdT
EaahC+W+awLOKBun7pr/BB8wCJU0JynbyspFSg+6v0gepFaUl+U7i5DLP3A/
zYOcteqLLhYD1SBVPOy8wQOP6TjadqzZmfkPu7j01Z5JrSO70NbqVFqOaUZD
Zw6FMitFtkJsl/Isea68XFUMjnepv/y/7jaHA/oDQRbQE+JB+beLP1GTBprU
8IJOBAPMwrezDbddPqTnYpB8z2eJZcUrZsKMlVQgBRM8TKck3pak3sytkWDg
P5MaPSuMoVYV+d5aSXimTTsjutNk+risbksWgpABSLGJkjJWoJssoIcPm/bk
MhCM03ImTxNdg9d5EU2gUakgp7zkYKBBnBIv+iAN4KnotTUxYUpA5eOEe6Wz
wkzkNVsucMDnsNSFmsZI+yIepTut6Mf0IU5Sm+tP4Yo8M1Mq64DTZbx3INgU
usPEhEXEk7NRCOA37QXSsfSuKhGR7cpoEx7OS4LxAQU9GgtZbEMjrLRtw/wN
O9+PhIUDtWoH/XecYs5h4h2wqW4t8FbckSeUcmSyrK6vyA22Yx51xwdwjoIq
sbH9j10C6kqPGvYZjSE6HmFRGQLcBCWm2GPH152AFMt917Blxg1/UDLx6rhF
eFx9uopRhgbwQM1r4qsnf4eK+BeBt7EH7ees48pz1lNkBy4uIPi9sIBZKutJ
egdDH8GG30QSUTRRsprNuA8wQY80mkVHwQyhz3G2dLa1i4zORsDZijhVvHGY
PJnKHltVEiiTWrD4YZQ/9JKOUneKqpTzBMiX3KVje1h1hs11aiFDafARdw4W
mIzE/4XfpurUbl2C3jVfNNCt5tLmowrj35xNsVKdjY7AgGEwJcrsNeq7dnbq
xx3bFTVH35IigPmm62IVmWBMmYtHQSe8cGpQ9Gn5jcknen1A/vcmEAsKuMb4
tX/5JAc2/eMoook5PvvSJPCtivNdjhL+Gu53v3GB7lJ/0GQYaBjqk+Dj3Ez4
V/bGFNVhbOqPGVWs0vHb4dT1YIvvW7zu3GQ2yWOfuYz01RzEoJkqT4Gnk0LQ
Wt6i26F2p078BEn3wsszKEjHwzKbTwe6AoN8jQ7c9Zi1X6b6Gv1sfAroN7u3
5KNNnZNhEcDPFLBk+ZjHMg6hstlzDsgTF6wohYLhKlaB8OYZPSaRe/agBd5c
fV0e0rXBuExJUYl6g6LD5tG2jpfWBsDIqv+KyHvDo5aVjgFfTXpctx8Hsu6H
Vw/7/ay5nQufv9km5wnN0ASpBHuUhWH8aiW7L7tRgi0b10y3ZKLmDKEQBYjf
PelG3MBIIFvcIfcLdf2JI4AwDCKy5eX3OSen6orFoPPOGi1YULpECDDj/Gpm
OCciHPRpbwENDOr5LmSniNZh34OK56qaQUaty5hchVabbkce7fUbdjv3exTU
JiKYvqQm1Ya4/3eZLgcNBfTt32lCpnazLER5yTCQ8mhtXI62LeDZeVoL+UJW
iTIggOsEVCBPTA2uZ/eBok4ddChboX3eLy65hwv7rJ7Bvu/Kf6npXauSoHku
Y/UN6ae2peO6iEvATPaihCGfhtPNQLpUfnApeeoxET7ffIWa16hCzDefMq+8
ZlcrCLHgqe4mzvEVFNvf8D9e+WjHkOL7ShkQAxlqa6ov4HRl4uIbVfqlHnBV
ub2ESfCRunKcbUlc5HBJziNfXtV1dZZDcxTrRFMYaICdfqtYzEcQ68r7sk22
+B1Gr8Kz7sgmnA6FQrv6qvq/OW6BReBigTCYqaszXuD+ZM3wnQycXV0/yRD4
OaVoqZlZvBkEYdgwOKeAxiI/jtYVQ+btfxzx2bN7pVkMtTK3WdQiZ8mxeYZZ
lqKaFyChsdUA8Lun4n+pGRFZA0p4le51aIIutbom/ocN/7jVA2aQIpCoqmDV
vfWk0wbVsT1za88bWLClTXGek5kfhwNZPvNVLytOSFrynmrEvcYQO6RHyS6T
IejncNKl+A4WVlYZqvo7hSgvLjUAq9L80Pz13lSU9pSzEaq5Ca6mw9s/mtVS
z679pGtro77/zaCxHri0jjC1eox7FgWxoeUMEea7xd61ruJ5CAkbpnl3cZy/
L8gys7EccQLkd819j4KmE0jPYczlMbgJU4eKLRpeFoRsibStdzg6cx/p6Y/I
lhp3evZNTtSgJXZSgNg56vmbSA/IDY0Ard8+xN3u/o6Il3yUlpaWCLu5wve+
OEYWrILDIKgpunwHQOONlopsWWDi6n47dudOkO1sqgeB/OdPptrgdZaCVY4Z
tVerLc6cvrOv1/fvIvxzPhPulNtY3Q1t2igxui1kxrTGV7p0L9FFfBWj5tvS
EQhTJUV6gxUr8DXd3PEiVHxuo2ALNJsFOBzRIYqGDjjs0iDuZZYF1ZD2LMck
nnY6+N8C2uMVC8d3xHtegPlFh9+5xQEg897BKib59QyuNp041Topu1s88g3q
A3+fzw43NqaS7PqYntexmb3jcMwlINWmLXqxjonf7plBPdpHdZPJ1XizR4aN
FH/gsn8S4ViurXonP63p5xSrDBg6Eis/uMO8Y4u7p19BZtfJtPC+0FocZ0kU
dquZkk1wSjy2hk6hnVHu2xUwtNfWWKNqUE+9EQg5Ghnlex4dN9TZ6KLUA1E1
WXPM/X92N1iitxunGqsjA5reHjCswxZJr7DMQY61Pdz36cefgJ0mv29+P4Br
iD3n+l7kjYCdQa4JNxBf+epm02i4tMZ3JE/eMXBi7/KqXWDROUdPtIwshrCV
H1nDOVBBgdiiSD9GQwFj8S5BIFbdUWErz1mmydgBti2o0W3LmHqmnagBYOWW
zxNei/h1/hqG1vWIQevDCYdVTWXBNpc14P+aBGTG42TfY+oMs2jAMi1WkB8T
KhLeuOt95IK/qHd2eZoaSuXYgqTDsoakbPKe8ekko7/Eb6ih+seej1PbMXJx
YJ+P6MQd8l66jr+CZXk7koOBe+je2IbBImr9RsVu4Gd1aFwV1aACyQsHDWAj
VcE1ykSvcGIUFFIbPzdFcOpxpam5B69nCNNwLqei9eFnKM3WdrZGLPhXYZHf
Gf8/X6O2paUBnB/9fMF/jUD+tjdfAeVYgzaS4dGiK5vX6TGsJtEtKYMJKNFM
4k0mtAk9JjHQ8bcmfb8dlDJUjh4O88exm03KqRPt6Dj/ERGMXBvBKaQKpJM9
9SP/Fu9ljRJIG6aYz6x/cJwb1jteNO41bBYum9x5T5DEkeEGm/cZnlibLlfi
UrpBeIQzpT4kcUqfwcNxFgiRQrcQbBo4QyvLarIJF2ybwc+Hs+YTTSz0Fuab
xMD7F1y6NoelR4H99I88DSNd7bwZ21r48NIOfN7a+b+I9bwop0hj0S/jjrhO
ZVEQKDwdiJZzGnO23/YC/L24n3h573v3X8Rfbt1DxZrQI825fbVvGGH5+tTl
c75xM5Sxc1zpGG3kSRKMC0GeiUyF7F7zGqCO7Sx7C48en4OkjO4VnF/YLwe+
g3mIfPcHOc10BPrLJb6ZT2MwWFbF6+rUS2UdAntQoiwvH5ZFvfjwimLg7V9i
hbvo344cSeDy99tWjgM2+B8sInyz+1tU/0TVAbc6VRumS8jb00PyuMQvvsdk
xoNSykLlE4pk7lXjGgH8XyL3qOVgxaajlYL240boYmB9Gjtji6txgyvgfeSH
LF8mWGXaGSl3Re+fdjMVzfdm1eBM/bitVI4wteIo3zsj6Vq7UTdl2+ZLp5O9
78nR2QiU2KBFBIG/HIAECL4Qvbgr8ihW55sNANW/Pp4uVxZH8cYO+3cr9tli
BT+jCkpPZnJZHK5m2Z5u4tVM4tn+ymljxMIRBNaAaYmIvhAZ8FmL9+lNbW2u
Yb8Y7y5XZsafKm4pG9hVrBg7Ji8rAK523AaEUWPnmy10njHHPSCuL9voFGQk
qSekC3W/A/GX8J2PmqKsfz1iwi4/PPvRGW2Ga1z+5XF1G4C56d8vmSJbS+0b
utsfjxatj9o0TyKQLrVE+HbfdHhPtybhgsIbb6nRak0TC5fDtAoaRHKNSCVF
79FO2lz0mrHZe1f7UbeBhyrcr3IBGCzhMSp1fZdcg6wUN7uy+P8vJxDFLSQ5
bkJVpFihktH3twnWCC4z91J2kHmrolEerP3MVFvrOIJzgwcdjPU+PE+TOZTl
gpGogdEzolrgNbON9bTNgK6YGx3Dl+l6HxFd0T7AaMWN9t0EhvoadPsrluD6
kWrNQTcPGgTGQl+QHIqpIvXR3cwhQBtM8+RR+eyqOpMvLqz6yCgbQ6x05CVc
JCsseUgtUsLBPOTaWHEAN/51e39DJiP3wWWl6j5PowdMW5JDko/wMsrxHOeG
DFF+DqZz0+TXvQXF4+2pUwFv1oRvbfhMG99q7tMfGfa4v9FttlUj2/zNfAkt
ULFUn8lZyF9Ol3qjhQ+v44S9eKbrhxFKtDcPncKe7bFoSwzt1bASayy7thgX
NIz4EmnzyFVS+rQ5eWazyLEeVkBCOQAVdMeLZtNYCDMGe3xGiGU9D1knMowc
pkTXcmAE/HYfhjuOiLtwWqOKF9xluw76/l62vly0AqgC3AHuZFoJtgzY+nvl
yWNylqa+NE8u4rnxRdp5McpamQHcDAantLnfr6ZCmhWKQ/jmV2EWEuBzBWk1
sVs80vTdafxiMfVijqVwIiqMgBWng6nQbMdHU5myqd0Nts4BpY+TZKNu0O8Z
1yz10hznUVkU22Iy55Dj9oX29Of/afoUjmLYmnlB7TOw1kJVOFge0tHZWgLN
oFpY3FJgOYEURE8ko8wjlsWFBhgz/69ZnXxE8dVQKphLVCDpXQHeG2Zduo9n
BVEM3vZHfRucUXZj8ZPL6J90jtDJSDGMUxlLdu5GMlUhkMCxCzN9nnmXm4FY
YOSvNcy38jCDavVXrwwDu1svu2unlr6M3iBlORJznY7uZKPTWpIEZRjG8Iwc
2sJ5WGAVncvFcE8UM5i0gBxcUZK9RHaQtfeDxUqlxW5jjdznhxRFA/71v9FI
6nvBg1bbQeZw8kLI+0Y2iNqKAEI47DdheA76p9E3GSA3Y2inSBDLh8zWPP/P
jO7NhMsi7TuCWZRoLo0bfzryFF4ApRhfTDoZlPXQy9h6M/I+xr4wUl/OXGU9
HlsiwYBXy1QI6YMB5eUf/aSrJ2nMuUGj3KXUJ/OJty3zQa6NPdST7UNnLarG
F6+u9HGK1qk9ScG8TiCIO0AtlrXOXxpgils3OSGzS1f80BgTOqD3Y18EzdB8
vcEe9SZjXRvS6M4sNJTDmh8th0o/fDlwCUmxTKFxkhsfVjtIpmJOtu0wflXX
nf5PCNDnA5x3S+2wSJoBcZzgiy/4A8pjRGu6PX3o3KSroQtzKeGmwFlycogG
4v2le7VVcgNSBQ17W4mrj6Blquu3cn/15YNBOT1o6WY/2lmPcH60OvW6fkPD
kD8AYpKMt7ZZg8hhcMuYxtjsLD83JVnnm5EhDhfUhTwOsE/aNh+6Cb/42YqE
oOKfIj1QXWG0pORWR5sKkuga2qFI3kdUhuEGeHx3RDbTAEzDLVqqDMwZL/um
v51GVgkq4crdyWpk7z9slWpm4c/7Dhedy3dqBDyA5W4RsgQNqUvAeXyjcP+t
RgmHtS2uJ3aArp63s9pudmbtUBVQVdwgAq8QR2TjRbsrtI9qqARvRhg2YcIJ
TEgzatNcoox3DhWFH7jxm5wOFgN36JJVYLuRTT2cGquF1ZRnUEGoF62q/Pfi
THOcg8MW+GIZRQyBemcZ9yaOCKYZ3GbO8GW+0+he0q5O2Ei+lVTjX7OzA1Bg
eIIn7R6NkYfSMIKaUDjx+v7lfOevDKtl11xno2hJ0mkPQ/p/wvHetYpauHZF
OP7lCXnzcCwE8zucBWYxNxccIPedIy/oOFX/erkRfCKLQeLz+O3wmKvJDZJz
zgLgZaVIPe6n2/eAmNvzNexm5mp6Gzp8cIwvyLLpbuKrHYhnYU+X63qwXzPI
y6wf3dYR8OyRAthhAR5RKXaqS03JlEFzGCzwSqpix0cA/zYT7WB1o0+EV80Z
0C+zrBDNWapO0Wyn70yMjPjPfD7jVEZFU0DpS32c672fXS8NbqS5j+dIzefA
vj8/mWbsQoEzr6Br7k7wWoS08NrMGLD+LFVjUjKyhkJV89P0ujbNX7IZBytB
aPu6T2jWC39M9/z364lj8lh3cTbYL1XXsZlxH5xjZkoa7B4xJ5P2lXreXjy/
KmDJ+lv9Q7frdgWnPIkBFEzfD0kbVba9JinLDN+jsMKb5l0464Z2sa1M9EtX
1fMG6lZFA4c2gjFv8AGXqUwYpMtD/SeBJ/NYgJtTzVVINESphAl0o2OrDX7v
L+Tm2eWaRRhEG+XPy1Ay7Oor5bSbn3MO0gk/wx/I/sVpDOSJQYa6FDrC4cum
vV/pnrthnM3yH/VyoNmf+jIdS9vtxYZiYY7KPlPQCJdnoQS2MEWN4/6uyGCE
DA9VOcavl0IK5UuvAcd0xTgqE8MudMJ6wfy1FXJHkH+t5UT8c3YW/eUgklpg
tF0lRUKMBtWLOiRKJ1Qk68XqtEmcgQjuncHUYhy3AXOOkIoPtUfWTsYMPQxx
Wy+XTWh+8lX+WR0VIOKyCG3L7bBHkZyWTTJ3fPaoUcUw7eCAK6677Zxr0pQ6
xELy7mh+xFIMDRg5HwvS8gf8THyRyXwIZpb0fmuoMH1ijNHyP/jKTr7EO+Vz
wXWvEOJ/SwFn62NAz9trZlbup1tiV7O90M2fkJchtfko6ItJXpOET+TqgkSP
3k1WoxKeLJIZSudKIh2hgiJr6VoDooYUFVLf6BcvF+l+sFIiX2EfrPuHuyxH
y4rvJoxS2jTLnQ/3KSAEDrwqiGscV4JMi4ZMzIFY1g4V5f+PezS+5wrWeFBo
ImwV+PCTv3O/OR4YBgMmoGaOqB6GaY9qlA0YBkDwJ8nURyKSc6tKP5B/iOrb
orW3fownCiMwWHlZa4TAzoyBuiUI/MPUzZqgqG0JMv4vv7yS6eIDgJNamz8T
cika+9FYqMm7ACvApPQggWcDYPQuQubFhKQ3rrc/a/6933I3AbnvPY0ohij7
o6Qv5wVDsgTSwZepLIWTvVllWnvQgk//2fS6VNicD5LTglQcLHSIw3eAMIhM
Lx/Din5D/cFrXnklk0ELABPmirqO379JjU4Pj/2pEEOIhXa2hm8eGzn7Vmg8
L1tmL3z3LujFAYWF8/CTET9z5PMKNUscx0HlLoh5nxGCLa9WIZ3Lnu+DVBDl
48Ry6jC9mrLPu1nPoibxxPH/5+pYYPuYOZyXp/6kV3HO7LLTjUafeQWgew1m
/GjlXLT6BNdgnZ3xhVVRayWFTh0qYRDuY8I4ddjKuJotsrxRmNI8Qy5iXgyE
ngPPekamRcsjeaHFO8lMpBW4YDC4wvZkD+yMNfVl1FpaC5YhUCfP5ro0QUSd
66s6FPdT/YgKtUNxLkpMAfKUvG0Nd3u4DtMzHcdS2oZmC+MlIWKG2/Y0/F/k
sCznWv4J/qT6mZcoTKa12oxhRMoZtzCTjvGyiHQ30GMp5gM2uYdSklaTQSeh
0rH/5uKQPy/ouoSjceI/cEoG3hnOCEAZfbLMyiSzPXOwi9hUaRX6QExxw8uf
EGdCiuTBxgKzsL6KBMPApoQd7xjEmZcwCtdpLoVOBNDnnFW3wDkJ49jYrbsO
sut+jC7xDQ7HDqhC7z53qGavH5iSW0m+jt8ZWADPPcvu2tBx0YNXMZXX71ey
Pm1Z0/lx1dr6HG54pBNTPMAmj7SXD9FuwiOEB8gIYe1papIOBDMQNvSvlhJg
yUcuOUrN0W7EtWJRAeD3680brxfvp9HlhpReDinjzR8c6RU8Hf9bknvDnjr5
dNEuTMEM42uAzuV/N5Y7gYI8LFdLtmNRIxWIh7sPg8wUBfR0Rkp53jwY+pDl
7AUkcCb3XrlZND8Jww0V8yBT75vzsgzzuD/Hyye0S/Jfk8qKaPHFjGwsMJ2p
2ujrud1Z2LjTPRosG/xygPkKbARRFikM/TzKIGTXpIZXU8b/qHnT9B0wB5Js
1v5QIopsdxqLG+rBcg/ytzmiEL7069J8BeraKG7r09ai+ECI1BtTs/emAoOA
SatFVHgErY262D/LzY9at/YUAjA48wq9SE5WCoOkRdIDRBcxCm58UN1O4+72
Yy3268yMg3IOnviFKw1BIFSoiW6nKYZ5yxtisrv2R11N6fQac/Rurb1DbLjh
v15WoHJUYfF7cUv3hg1/OittV/fgcmRAX3gGEsSCruqtJbGch/RuO/bn6zjg
LNcdmbBEqxHAxiQaNfDxnNwbHIFWhU5Y0TzUfpCtHuWiLYc1oeOFDlGgOzB5
g0d3yC3hm0Ga2SMVg/PC1IQVkiaqyUQMNDxAIEkGuSkMqRfOL/nqWLMt6Muy
qi6IhBMdHEe/GdQjHoRAvFjgYevd0/1+At/qRf6CemDkvD7M3b6OZVUrmR8h
/5TZePQeXx7+wk5ZA46WSldMjy0lwh0OjEReUB8qT8paGnDtAtH4xAbq6X8N
eVu+wkek46eRLWJBidVABxpeESAm9aoSxu7sYzqM1khHaJL9ZuFfYJzIB35g
lmYPURkS4haRyxG9ZMwVgRDM/Ovzfnme0onQRleFCKnRghFnEFVj4UQGiINP
bRmGtuKSCIuAyFUVrV+vnAwk2RyypbcsTU+itFNRAJctXHHMtr4OJbjted5P
YRyhL42NpFpePMSLS3vo/QhY+Q76JQnlrhMzTcK8m3EZhepFAmY4i0LIcuV+
QqiD5PwE+CDM1/1UTPCOHQY4nWHg1qTZhs49GyMAdx0lGvOiKiT3PGKKbarf
/hOJ48ehUbhDyesMXNs/LI+CqPSuwzXXXor4BmsoeoY6kYLElxSm/UQb+GMu
fD9H+i+jGaN/iAZ/IxH9KGhCukyI8gR3LhSqReYYNDTpIc7H2kosP6suS9qL
2831z48HWtO7JiOThcEGk3o6eWeoy65Tx3ak1cmLodMLnHD11PKm5KyZOI9X
w2ry8HcrmLaTYFXDXQ3kWKARa8X/HmihDRu0R7b6oQuWgmL/4fH/jwneIQrL
fCAlKRIX9jl46zAbZ6xT7S2vgesXapxiJJ2QS/oYBwhVDcICSU3ZFJrttZCY
wlnJ7DdcM9xzExF3ljfWck2nTt62hPOOxHKVDnIhXBgw0HK11WvkuOt5qttX
k/JD27WkmqIpvowjYCiHR7VId4hC+RuLdxqOft+se6K9O09bG+A0kfJlPtnU
MoxZbwzLA0XPAUXAvB29TyLbC2xfvSg3Fyy1nThRHFpla4Pu/O+z/yYAsxe9
MhXXAc4zkI7y1l2N/9GB9wW/RfcjNdEh0qPF0WPe3P4uOPJa9QPy8VvmjjSl
zQ+ULpXHrm2GW7QANRsDOscwPRXkJmQXNaKjCnOIB6+1OmD7eFXKtbj1hWwf
QuylsMAeqEfQplWAWHUCDx4lEkqmEWh5jCmdF9zJyAhaF+jCNSPBsxvcteUI
MqE+FzX4xWZJ+aZFv9i5RaQSPDSm4CkOjiroNqz05algyWLKq/0P/tioQLwT
7HAvDRv3OizLazy5yUOXONqJ8DTi+AS76EPiI1QGvc/eR6hcG42im3KX0jKX
7krPpVJpe1HZ8vYaY6Vg2RifDysARHnf5TffSRC9TrpECFfJbAh1OKAWfpuf
/MiNKchPDSGVYEXCaSLoMvd+hA8yLrBgtjTgwU7wFFVZfwzN1TO6qg4rqeZU
EMyBupoMr9ffRwCeifqrG1PIfx3EStsbzIFIAnxsj5/bvu+8zAqNYCQNYqzQ
aKRdRHlZA76X9KmvWFuYC+/NtOKgNnPFd6b1FXe9xZ4gETqnzVcaJLJsT4oR
seKh4xDmT7A4ehjup77wG6nOqjG0ng7a7+vWZIZ4bKy4lSWl6GH3IttPePDC
RRHfQWkZpnO7vfI1JJbXXSn4hrd0eXBjx75CxUHCXuKtwiJZ/jrj3QsMNJze
DTKDOIih6EafI7qb3OVs5xmhUu+2kNAwuFfBDDmfo0Kq4/7ab1/x7iQtI/Yq
Pz2dgy6tybiKIbOqL1gQwFhYagULQshlK+0/U5IUpkPyQtuwblEz+J0ZKaBh
avMSL8cfR8bbWjogGT2DRdqLevcTiJvIoBhuvxWiGme5Y33C+YJs76wacPgk
w9v1D23aShakPX8mZCvftccfhFcyqT84vYZDUubhcIaRZw3FVv13XkQwMkLx
HED82hUsnSmdUvB4uIKs8JP1XZ9ktwMizYaVqTGGVV6xtRi++ivt3sl0dwH+
pL/UqgxYfJu2VdCtkkl1ZAP6RCf8DbfHTofiXFeZu0r2kJQ5v2LX9WK5VqNC
3sEkXpvN1RovRADZDeDZPcqCEtg7mjOi+CEZesxoA5zd7EKsLwWhnc54HHiS
xqQIHI4TvtIvk+EeM1NcJYXqGjVyYzoOIpzQ+a3jiXsj+ItmzxCquwX+GED5
u8lhr6lwBa40UR3GU3sW7s784FkiPOxS+NDl2R09/7g6uaLLDNA75Y/FA7ni
Yw2R1uMdBP3nyE3U7cd7DnfLzXNJz+RPeN1jAtZSrj/s0PV1Jugj6F8YKMaw
f5qbUmsF5atKFHSBzFesF2utyiB/fKf/m4NCSkWnyOcGXQDw3DDW3Elcfyl0
PaTKfhq6truSI3InVNlPIINtTbkFsJKOee13MRm7mFE1qhS8Q6UKIMDe5Z7L
RJ1MqEkGoaTJJzWwiq9A7xGdwT7d6sHPXIhxiZchaJvf28L3yZ9H8NT5yjbO
fWPCuvHBvpyIwAO+dtPyB7jzxhZOpBJksF/r6G8Fs25E87Og54k97Z9Q5nmL
W9jEV9wlORgKQAUSKHhU46FkKuTiX1vkL/+7sNJmGA30iHRQjGegF5t1VGRU
zQOS2eDPu6rfgfJQCkN5SEn5S3eY9ZmHOiQJgErnbudZMY/CFek2PQj2bfpM
PsZV5a2TKSCdVTuOaj9Br89NosyEa133qO9rnxe1Tg0jKmsWHlltnNHRREzb
tWB+C6+vJfzVaWJ+dNoMmWBUjUu4PtDcW4J41ygNW82mcGvq4HMGrztuwNmr
fbtbnKiEbSiRKTvTxhss7DBNxGyszd5rRSvO3Sea9enO0PnEkOpNtxV0TMWD
WP5Ta03vE3a5th11juqpXG5GDB++W7jiGQzrHIpFhzxU8qvJiYPKKktTCGZa
K6O9wbVipjq5W/P5Gbr7W3BvmfbL5gZSCAaV6p+w+2lac3j2lb8DbxatlEOc
ps4KmuuC9DHZQBt9duMnUrFIVD4OT+JrNM35wnev1PZsMWs4tq1rBXm7ku37
c6S7bzxcFxZ0MyhiI6v8yeTfsGaOxdWlZHMooHMNNWGjUy/W93Ie0LKPhYgT
e+h8bbIbCH1q1xOpjwxkKk0QQ9iMqH7fzkk4BHV6Si53a1Sxk7BR0rSNF0Ox
nYYO0qXAUEnwWkM2d/CJe2FkPhNpzu2+VIj6C3hQF6Bmn2pOh6BkRfQhaD3t
RHcx/u1QsEHb97hxth5V8cbLl52s86qIKBF5oeigjt8jdcpXA/6pOypX8xlT
TK7yHoROV4sN1ifcanXH3oN75b0pBlRQw/r3I13KnNgsOFIkBQaPSnmgcfaT
vNDb9QJe0evZ3BDT7Aqzfbhrf7+u/B+AQlsxpzi+Mk63JjJqDEaWo29ql4m9
ysVsuhGs7oT4tbj/Y/sFM4kLmZX6Z6cHMmOdAIQq7PAJiESHmZbZhfxafGfF
d+3FFVa/IS+nf6PT0TYEdjko8HLXjdwuGnQG40AtuLdYAHqbLM0xHD2va5yr
9mDTexUGvz1/D8IZliGv3ZKcQ5m6Mju4N7FHn6VVnH+PfAY2gnzVYSGar/J9
mPHhJXPLmgjNAznVg9xGmd9JlcWnoHHmc3NSdx+Ra6fWawg2dl5qk7loFGZY
I8faHCUSyF3kZY+VzEr479m3DJovHt5aYWCVXcZzYnMYWYJO744=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+EojEp2q93tF7Nuhqar8kEv86drq3ri/6E6OFMJAsIljYWw9af1sNw0XZZy01X7+C3gi6/+Eme5oiBPU21PX/m0xqoY0PLGOx1wkBymdTxJVbNQNOpmxLcAE/RYlPv/c12WBHWxwkmoFJ8ESpGw/NDJrhNXjPKzAVKzsKKBeuR4dTMuFo544BWeCxdU4q4ARaa+VOm/2h50V3h81zaLJR6P1bjOLkYBcEbNAQtJUc1wHLRmFKsd3AFve5f5ShyFZ08Pmgzk1sm9l7ypCuqKFwxdCqFRNutafJkjtrvrriY4WtLHpDs/UdCvMPXQG24mwDv2lsP5vN8qeODV3mdk60F1RA1jrrmqH9dy61r6HzXzJV3OpeKzCZI0B1JDr1nFniokZAgiW4jrlHa/YiTFXKvlyIg+zmYU7LOrUG6lw6e6n+z3Mp7LQT9tbU/y7y4XnEgZOUgoYIOXdsAaAto/t1ieIVzBh7ZEQq/r4tdmaHGVqMF0IoSRcbPCzPc0cMazBE3DQ5uBxX+8NATIC57E7ktBiZYIbDe8ZFRgd1/VihDC9mngmmt+9zTCGb3kPQ96piS5+s4ag22JsZZVGqYYivxwlv+fgz9cDsJm5j6GOyv0KsIu2LDoM0qJtLhmR/v4ssdqVYSiuiqqCZOqH3fC1xM5SLIHY+wOHGcSntjFPgQ6TQPuJ66Dg0eaef3qSLiUBCeMq8OM6nNaM677j5xPbvPamUFPvdq9hLwX1mhMm0aMc2aKd8speGKmRqKqHWd2xEQsS5nQefn7sgbG+7+cLxwPZ"
`endif