// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ipGkPdy8NJk6i2KBun/F3bEmyxNPVEBkRPrgapvovkDvVclfseRcl0hYAxpW
va1qoGjhdG4+zvWmmdeRJbWDpljX5KaKR0Z4gW/uqlhpgZ/qXQQacBMnrnax
SDYIsb41ijtjsgsD7poAi4oiY9Lx1exuXYi2YfCDQG9xmJp32+Byrywj0l/O
dIPlgNcrtdWktvJh8LwgZS0Q99JoRmIvXMFj2keBazS2hxzKI4F8bYhYgK7x
jmPlar4JcrO1oeJowIBUFo4BWMZ3THbl2p5nkRd9BhraCNlPJyLCMp/wKTzr
nsXCZmFDeJAXFosfcTtcMfUt2dkyYTSK+UwiTpStWw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WOff0tXyaZrbL9hgNHayrPH9PTIDstbMBmyXlMDlzS0cuIXbaHhaHUqMdTeZ
RSw15lM6ws91jsyjRnejS7smYqWJk8CFJTwJ89IMlrddlHVz2iTibXkQ7RIw
1WRcSY3tXMQmHYARy/asfiE15Xw7iWRnulwJ0Gamg/X3m88+1dm+Eo9iZhnV
oHY9Cao78x0G41hGnuCpvP7ZrmM2wmfnGRXOd21KCbeadyt+GGSNdnRXQiOg
tj5aVtz3vQB10wQGBWbS1aBS1P0Z6aXlEBozuKB2tU7K5om8S26l5sRMlj8X
LjJFtRXdoV/87ndyLE9rESRXGgjFeQLvbTEu5ZOB/w==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
K0cPentFgm4w1ohB/cS33asGFY/65aIs/GgUoH7peQ5HIVdZxqTiVw+iBEy0
kjxIHgQHSja586QFrq/KV7kyoGoW/6m55G6w1G0gwzJdQ2lyvLbgUcaiab98
/45lOsxjlcVA+IfBzHW0Xwz5vXnPBCsSx6zpcIxQuluQkWj4PJ1W1pePr2zJ
b1pW2dye/t3VcOA7IarDPD/Z2aMoSVgw+Zk9vvXfJjBs4YXktJcaCHbrPuY5
aggeVh0pMcNNUseZbS7uf+1yVAfJl9HtpioQ74+QgLzv3rkYiszV9zfccAJE
N2rsjVDs5fw3sPXbFKg87ajABlqTw8vIkMxcIZrTlQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GeUCPE+xtBLM0TQFLWcoSV+/xc+l/cf3uXoWuRNCuKBh8KbDxaO/DbJ6bTKk
a2JAtREjrdlKMSyXPjWTj82m9XPzgZ7pTckWnxLthO5X5ECG3sKyRBeMNeZH
QWjdp/ammgc6s7W5ottmpo7JRM9TI4D7vmVHgU9JJJbLCP66qrnwHqQBTkq6
0IB72gNVlPg3qvKKsHIfrf3uyUmJ/1NtLKFhoFktNcg+YnV+qPbAUHYtEuJg
2IsoMh4vJLGCP0gadKJqp4QgYs6a7/A0eQUCPtKsnoqSCiX3d+RBg+vwv4CS
i0dOhSGtThl9u0T/stL1Hji+65ohB3r73K4YMG4gLA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Gq8kwf5U4ykuXK2jIcWeCbdnb88oyWkWUUFj3T5bFzDErOQXiRz+l64Fq4QS
Fbo5wOf+f0FRTYm4ftAtNjwNmP6rFURIzlZEIy2FCv/P5rOIfhJUie/rEFlp
ta7u8/7jYsUQHZ+HlHEVvtRgPXyDYXPCTNwlPlP4vi7cPvF+6ro=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
IIn/+dWdi+U87HMvaOzOyqys+VF4DIryvI5914zRe97lPgVfOwP/KUojujcf
/lzwMbGdCccrzrgJYWlNrR52jX0AARxZN+HXCZKp9meJqI/J5TxEi7UKnLgH
OQs2rKU9AGo+IE4Z2nNZMDjrhJZTPlRhYimfqr9J7z1eU3djOGuvCezEdlGt
cuwscfjIRN3qDvPOmmRz3gDNK9QZlRLKgWjbEoRofbniUwZod5elOaX8hx4Z
8wYVaUyUhRL3FRdq6PXv5J9n36kqjwSpn42FREEaG+kRsPe4mJt11zUGmEBk
EXzMlYFUVOGicOd0AUJHlid9Tffjrfhi6u+cYa6l7VQviLhGmSO1KZorf+Uh
nrulH7QjlSLPbSkJEaUy9JBk4mxIOJfOiVGDwPnKS+zy7mZyeLidWBHgfExI
vk32QinvZKh+ICW0FX4uCjPOihdTzQqcizeJRdP6uUUu7QELDgxQOxM03skk
L84Dqm0ccTWebt2Mv6K3yNZOmGnXopRr


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
prPYjRWSimemkEhj1Ty+q1tgxGKJk4JLVGR8Opdq52CUZg16UiK/5ahFPgi9
0qXhUBFBdlxfflMkpufIiNJPADsPc7reNMK004siOwlrchqBP5cF/sEJ20TF
trJFZXV8jC/6aRlIAOQ1SP2tyRzpo2v8w4cqRF/47bDn4lHRWNk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YYAOHoQ3xvamVVvjV51JzM2du7i6iDoGoZ9HMrB728YC4+s5PKLxcNiRruPW
9fe/kIKcz6urgQGIvyPTUrAx04479fy7vnh1SaVWfvLIYeBTdoHq5PfgEybd
bpCAQIiVF2ZEtGR+AFjwkwBqGhvb5gSUwpvzkJNQOtkklY920RI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9008)
`pragma protect data_block
knPXMIZfAdTZz5ycoZ20c0V/JWK+yWTtsE3Hl24yy7xMXcwnSopIDlzaRZGI
DGu8i/rbtLQwRUOo+tEBenLqZXNh/vUKnQR1ez8aHXTN7NgXjJmbPBjhcbfO
gJH289ANaMkLOaIX9kmhwuj3cwBdLwkp4AIqZRHGY03/VD6R3YbdD3M6Sdkj
+I9ryoqwdeKpr1H3Iw8t6XS9F9QscDjEd5/AYxgSmM6/hiXlTV28HlMOK6nG
CNReEKraAWQaS9PzMHTpUzPXgiTsBxDCXmedtj0yIMoBApCfcg1psiTG7Rpv
VUCHq/Jqz8KTekJNCpFMdYVQf3TJYMSkY4phyUPSEA272/sOClsraMrQ0OuO
BXbg58ZtF3Ln7gaPsPBNaVr23m6ynYtMmfaj3gAoA2HKTe3OG2AqxJsQCEeW
bCGwKtvfjYnuUVMmi849Vwf+WidraJk1s4EzvqyHolWLxAOQmAzj+pQXJZfb
NtOOY3veddW1DUUFs8GtbBj4ebymsVaLSR8J+AVmiG5XgjfvXFs4wYl7Co7S
lb0svJ5mfPzkaBRL00ocnTAaPLNM52jTVr222GpO5R1l5ROBBZf7DQggJklR
VEs4ANH7efl4qkNrrHWAzQCX6yVPjO0RKI0d6n0im/m3cEOMZutvASe8gqgl
myxn3Opt8BQP8asnC2WJHlWr+3zmz3dC/MSBc2bU4Xq5A49FyOMSILUMXxDG
r/2fwZxMv+ur6JWcf4NmYoCEV2eTUFj1QtwEs+13XPFsfzn3beRqWoZvgoVH
0FFxBtsZVzmooMrKH5oNmoNpHIvGaVJGRdhgc4CKzxqnu7TfwZJkVTUxOmvD
yQfF9KfrdKLnMZ/SSzGJmH2SEFVtUCOVmTtUaZpw5oBB3hdm2JRNXH7FRYrT
HYKVMXjHQMYj4Ex4gQmAn5h+dqxNA1lulSPEvLzEeNxJG9Uh8sqS3p/3I1xZ
uN0Tck1CTxkzdlYc8T8a0taHxl7e4CTygJkf5/dgLsZOiiw8j+3Rimc/9RgY
3KhfB1NNFrqqyHmk7rhud6x5iWtXrgt/tnQxZnTpfChlbQNoGpOyeo273wYh
3LiO8+m+DE39MbzGHYsKH1R4656+xKD16BJRnzlyMuP/i4g1mJf17ssI74rn
NsTMNFg+s0dTL+hmhjacRCK2zklBn9UDQ9I4gkaWWR7YdO3h82nmbWwe/z2I
ksqyVa1VYh4vT5IxaCfICtZj2BH19GUqiCrcglChF94QrquDLrxvTWXpCGum
Z/mf8DtgccBHOV++g0lFmtOPcXQhLgx4kIJzLm1t54hTBPBmeSZhtHVjyFJr
Fwg5rQmWLILqJttQdSTdeA4fOaIsW0cFeh+aeEHZfxjyPEuyLbUL3e/j2NLM
/n3jjn/3vN9nHJ9xnG7bevCAKytdKo1hvfIeEaz/84xahrAABUVPmrgA20fX
kSt0JpdiDwKwvPceg9afgoJd9YCwlEcFPsQG+vMcpUP6A9zrvHKRam5DZfZj
hCK1NYdC0rsrhC6vmtY6jWno6eltGfuaTg9lgybi0nOPFaupwivPDqhkAHbe
KEjuOdHA75Wbif0yg2yl2cVWMD0PxCSVtsduvDZkrYc4+Kzmd9f0yBelB187
UkEUpkCLQZ75rnYY/Y0XwJqLiXfFVIz6YTsSnEB9eGu1Wl9NlXsR2DHD8B/x
+ncql1tgBuN/paOm7fWyhfc5ibDuw0c+IwbnkUx/e4yVNvj/SPQbLUYYXHEi
5xp3vAn4CPZzXQF+yw4Iv7w1GOJxKhM0n1OFmeRaeHa5N8ZQozRjo3D4bOjK
Dho7BTHnENuUlAHpf7kJiaBeSLAvVRS1GG+QocttNuoR0ZOvrrJbYi1WKtEe
ROt/yy0uBg/4n83182lwjSCzHRKR0os6K6u14oNHR/Zd7IploHAKgJSoOxp7
cR+o2PJX4eMDjWEbooNJb9hBYV+rI5f0sVWNl255zFA2UKHBV2iV5LEjqxZg
ts3kbe2RiS2ROJKAVne3kFUMCWHz/2oecb/xfN3WrIGszsNsk0Hqal20xeBz
0DEX3NUEIWajuEz2AP/mcfI10P9fvn1+hoGzRzFdpkAWxPAJvEqW6x1GA2sB
fiiuB/4bLv47sXw9SBOKVG2yQFrEnWJjLR+bRqpI9XrUano+1kQWA8KEHDhL
TnHWREUpQuRa7fakdYU0w0u+7Q4IHLdV89wu4JZ83Zh1jS0BNJGvGItKoABb
BYeRRAo9pm53ZfJeL3BRgbbIehEL+z6gn84FHArG7mPfkIOklZzMj+6J/Hts
EEATOalfngHGL3sSs65Q3aVRhxZbqZzMAaF3SVqkusYKADcEqViZRJidMlIF
BVwcEgevMWf4CZwNkZjobYfWF3KkuorVkakpud1sDTOxPAytaFPrYxPTihs3
IGhLDjXIkreaJ/Q29Ky+laKGPph3zpV5/EWnqNHFRJgqeEmTDqVr9JIfwIxD
k0FrGV4fX0XtTD5gfvZKH6kMLeeWYThkUVPI4u0JJZ5MjbNFv2S/KgT4mRhq
uPzM0FZdGYsxxJL//y2REmfUGejp90XkEUjwkQOxpZsSjT0APHeVeY5FaQ+S
2a1DiHkjfy10WA8w1/QoQbif6S8mVZwOs7toBJ+r1sqnMkdEpiaxjqHuWF35
S9a9JzG8JmMJRdjrKjSs5dXdMUK69NNPor2NdmmznglhqRPsDIHIGTA7/fja
ZTsbn32Qu09+MEweMNoHJASOSXwO4F7ENhrTccSIdqgGKMPdxLoVS4P1oZ07
Z3TrVNdi6sT7d/jkZjBSZ5nHWO2ypsNQa3dJWUgCoHHmKpA+XiQWicT8zrnb
yWLbkZAsPchJzaNfVPeK/50q4AQd2PMgxQifQMfzJdyUHf5qWce0XlqwmJa/
8mM/omWufGbOILxG0Zb4bvYWcjifpWIylmhjh/c3/xcUEY+M0e4r0zVSWD8q
EFUrfn4lFvFe9csWIJAJUj31SWQWY62yBNI8gojpoUmU6Et0oVJn2E87pJFX
ydENw9r+UK5fy3itJ/pndXJYl22Vm4OUaEdQHhiLVPHtGk1KOMkTJyisDwsG
g/GS1T5awn4tOb3EyeZ9wv2m4/JrKZ6HxwTg7fJA82BEfBOWVbRlIATNN9Zh
T7XMuAAfyixnxmSNBKWrII5gv9ruA6QAjVVaBjfOAbVEzgdMFCkrmrfh7WF0
LMqktaGMOdWrNvXjKJZON8GqomOKtHkG5JYLMBnQH4Mppn5KdoEACZGDjrC8
xFDD+rcIC6ndl4GjPq9QmSqK6CmGxj4628rbLDsL5LM1NMo0A6hZ7I3gaxfK
rq/uqnIE8FjLvNEY5z3z3vXQjNehhnqyHRSn6aUU6ZCu1AKnQTnW4rXKaT31
dHyjyzXDQSj/DKpk+ZHDXHPCZ9fxzf5u1LaImBEiw6c7taHpvRcyO/zvbJEe
XlUAFnSv7grXRROsA31bo64W1te54mG70VQLAJ7DkXU4c126h9lowF8KNkP1
rD3nmaoJjS7JeZ9eDRfjNagbieH7tWJMI7iURiFAIv7T8NqloiEvqW9HCrj/
E8yUBRy2pq6YnroNyiH33mZ9qX/1RUiyROu51t6LQO0NvmNwSFj3X3Pf7T8m
QYzSQ7+aD56FYDIYS4Mg1uuIi4vJsA3g0dGk9iRy4okNTYIvHLDHvEdMrxAE
3+rm3R5ibijCDTec8On+h/+VQEHQWgLm5XVtjDq2HHWXGK85kapjFaUKpfV9
DsSu2qcempHwK9raaaN64bn0u0ELrThlksUR5YBHSsIcb2gfxPfZHjFZ1YUw
mchjkK/iaP3Xt/DL2+e5hejsjiXR6jhZAxztWP5h4ox51ZOiuxI/XpTZiVD5
xM4q5+OGUhIHW6pOR7ZkWfw2w76mTkvSI49tEBagiJI6yCb5De90kTEWszXW
2Hv2BM8kij6AHpL104Gk9LAPRThLi6usPNAqJIHduXOw9rJ1HuWJVoMwWrw+
BolVQsPoZLa2Q9zNE9JOc9BwKwzn5lQFCzvk3U58vAHSKn9Fy48nKnYsW8nM
z26STS/uIR+sABHtKocJou4be4gtD0fV0o/ZDKLW6PLFyB1eQJUj+ipBdwAs
2q7gNbLv0KiRE4VZc8gyY75OZZkz5xIDWjzpxrgBOO04CDKDTR0yhx8VGwb7
4WmzP8q6/s65ENJv0U/KSRJiJBTCuzdIYIzpwO8C3ohxh7IFsr4qpZh5Gegc
WShBE3s40gFvH2dKwByIrOAlOL2E0EhhNeDe9/WzYpBMPUFgNopy7Ome6LII
LnDZsd/rHXleXBEWdrjWEHljjN5Awn0t9JB/F6Cs1pvaue2FQ24I3R//Q4ZX
NV4lOchzxip5mVV77Ldqz+/e64bmh7bco3yMQpNVuxedahYKiD82rZ/GAm0D
8X2qdJgef9kyL6zSF54zjSVICla1HL4e8oRY8RNPOR/GLoI2T7r0hAjz9mp6
rYaCC+kGN5dIAFvSgGGl5R1AOZ6aTo2JJ/eeLzvOK3DLYwK/DEkpTB33xCgA
dEoGaiLV5Edgl/nFQTLNsD8A1yyHb1bqcv4UJ1hR60+gS+45txMfFesWMC3t
CMhb71vbeksrM55jihSN3JOIU4YLoij2lKb/xglRBafty3qUxnDY/KLjiEBm
+YMoG22FEgW3j7mlBqNVivJrC0HRpZym03TNKsqB6HSo2IZpar6AeazNtGgs
yPQGF0m3doUiK9LJHvlemTGZCuU7zF28lqIFVnuG13U/2cRvcn7TNJpuIq55
LiBvoevgxKc2eByVl0ySOWTlDjMYDay+j2wmNVTzXgl5/xxM/y81oCXMSB5+
S+m3tzfrWAvA+9oAexFZQC+ST2KApy9KZo2h5RwejkME4i3YtPjnbefuiBDn
rwXz5X4Mjpm1TeK6h1ieZNMAtOrKSVTvXTFpCaCHQiaDU0iiUu6yzEBvOTAi
DmlbeXrv0p++A4d+yBHJpKHXFAQk5tu6YTlP/iAcy4iezZ5OD21SYbibRtK/
3nmJjxnGAd7PIbA+aiaIUuHZd0LomMSFB5J0Mfldt7BtCRDQTTuCu7gInGTd
n69EDpxEjFOPAC8LTrD7gOxsMePGA3eeA51LgDjh4d+eMDJMXIht2xR6piaz
xHH7DHZEiVVwg2HT9AsuX+n0pZ6HPSZie3k9uqWkHLJ8PdCdoW6w0nQxa3mQ
MzC0N7B/z47ARG6B8g+XhdlwFJadM6nS0PsRwlGs0UF+hMJOodH6tmR9kztS
qnHn818fWIpg+Rgt0CjpmvqcIr0Kki68GhxPYBZeawRkXgYQJ0BO1PW9YeZ/
BXTT10x8//ejpBoNTJ2it7Gc81CjEGrxq/Kkg0fzJvqJvi/2IywQXFZloZPO
GrTDYqYmgBvsYTUqKXF8HK6TeUyivDU7TBXusF+2z/v11FT2UCljcdJc/djH
2SWWVGVp2kyt6pO7JlIgD4kJQ25PO/+JKX+T91CcaWOoPEVpBgRU3/RsXboh
ncs5Tbha7+lpGGoC86mfyDZi2ZfSNOjNe3XHupKImB+DZvDOLhZthrjAPUA3
u7i9IA8kIkN5y3N8YC7IFr7PM2GzCRAFIDtoG6YJ3gFZ//pTxrXdQrB8uZmH
5PlkmBlF8x2j1wsjV82y+zDOyynH4P3yro+ZhY113qCtoaP2y8/ebB6kYCbm
FwUJxKPHIYCGWR603krqZFHyimZvIUV99IHGEzkiOJPog6Kp5TRGIAtiFqpH
ZTHWDlTtYljHb/akPg+PMTXSARGKlOGw6DuUHWWmfSnHE7hrZ62TneNUg0aW
J4hBJWT/a9u075/2IwnuPNt8jqAcqm7UvOrXZDFSBMZetJERhjKEFvgMpzpz
eU9HTB9CAsLRMo34M12nSqyWc4c1j3kLUsE020oPlyRtY4tSiGjtujRFJDow
kmm8y+FBwNh45bwdhvMX8HAyfF+E7Gr1/1bvOKezb97unAvGYSXbGZ4UCpVV
4DddeR8VQN2A1B9vaNoto++5mZasERNdzGZxC1TY6CW7tySyPsnNQ7fmohsx
jfqit9eHanYxa+Gy4q91nmRsREuk/Iol+yYQjtVAy/cWvfP5ljkTRXJt6QHq
OUuOc7CCl2+uGumtFRfJ0J7qBAw5B0tqX8G90jXL6euEAB25sd4coHvJTBo3
+TDNl4rGWpNP8Kw4dNXvqhEBaRWLqWP4kd2dbyMqEfP+NdKLMiigg/xaIsMR
+300k4irlFDve3bJmgAuzMlJTdH0/2IVwkUdWiGGEg023RMqkebtkBtlbmoY
qxMR3esFy7MR3tGa6J/eE1w5M5LvKaLQlvflWyS6TqpWnpLdqRexlX7EpSWF
jdeV2VIGDWMRzTz06Rnoob8Dp3yzTD5Vv7KKNy/ykG+Bl8j8cjtMqF+IE4Yr
ZbM2qOXylzuRazjQnSYdyOYK7gaOy9fbqXrkDHqKH+Pg9pFwJKzXKtR05TlE
xaIaL99laDVUX9aWstBdUtMf1sSynWoWq00jefg3iOYyTvQl4trzC9m+8+W+
5ZjzmgrFppTsT5DN7ggh4/JQhapAgh4qinmO0FjU/RcAVho7DyVa86l2BrAD
50UiiCqpPOPhKbLMp3KDCQ8cEyBtVbXsRYhbYiLmPGuhSgi3fGPLER4DdvD+
NEOefac/IzuOv2VfTTwmNU3UWx+/20pqGfNQP3CVP3+E7l6ZzkkjRLpLyaWQ
NPtQleiinxC6DRTtIkym841gaJYcR8Z8Jn4t7LBvIJlFljPNynWAtQq++Ceh
3Yb/fcvBB8biumP5kC8eNazbh2EhsGeUx5eVavuHYZF1/EpfGQ20dTKi1G3c
Qn9GXYwxLYY+xpA22qkkGVmfuLYPeTntYifk4w3mYKVpm7aJJETldV+LzSIG
om5nXirXQGQicv++MZhnlNUroupluPER7hNdfvwRdSzQpbhwHZ9w6SAG9aSV
dYHXBXyFA7mHMpr/VMWaRG62qZKqanInF61xEWd9o/67tTdboz+BIWHb+XSl
/ENd4IibFvIs5tpRVBAyvro3IRFKRcSNFrDOY2i6vjgC2VjliFgtamdl1Phz
6bQhMKQlkfSjmpQbq8NIeNeRnqvcExpCjwyH8KW15Zl6Dmgl6M8/iVrqYJCx
gqYpdf2f2e5R5VwbQSKQYsacP9GdlNAHC8mzaZgPOQFT33nFJHvvxxwyvM+s
W3ubgMRM9C2aGbuhTNsbYBGtXPyuYTM97+MYWD80TRE8oYRW4Npeyq+bt14y
pUHZFs76kRZTwp4qZcy7ABD15D04nZHgAZksBACqnh2siW9AN8pnQdXrdM75
qGFLV3Y1pFM3dA53y/+R9ICICwAXZkNq1NbL/goKKdP+MhvmA/Az+RCH7aBl
J+vrFcgXwaB0qooAHJaryv+6nRitCMcAZ+DimoQrUm73+WntQOaiAizuReCp
mDST2Ux0YYsv+lG5l4Q80pNQ/9JM4h323IQNXdV77KJho7/jCBo6EC7M5/Pp
+gYynhFlB0xoTJCaqbX8p4FD0DpGezf4gGhvYpV7gdRoO6/GfPOU5XLPNHA9
k8VAg9lSg5+08rTg5B2ksnXVppytjJ5M5k7Shkg9YVE9AyQgyWe+cqPpHmb1
vEadyd32uZ6LFbK6+GlqJWcpvqbXGqKDsINvKJ5nFQDe/HFQjKacZ+OiDcka
TWBZvXVdq6Q6pVXtRliRSm6VhS3VMYB1kWtOkOp2htVJ5JoSI4kkz36tih0n
7O4RZ6w/k+Sql4/DoXJtZ+8iS5gJy0fMeBO/H6nc6AxAykfhQmOId/jnNqxn
XPe2fe/ArbvLECJ6VxaB+jaJ62cdow3hSdGMxBll33vN8spH6vvWI5p95Z4r
WSdEf67/hOIRMovRdGqO6FU1jREDJxBU4yqfnR3ZKfX88ZuZf7/X0JVGCi95
dPOBCCnGYMGatAbu9lCweMSecHuOXm2yDGGKvFPdrjwT3MH0N4Vd/bT3mGNV
WMrn8oMstSjP8xEpzQWBduBzTqrkRDIVHGQTduZn5zidtrScEYT/Bbou9rHy
Mc1G/QsYD1J6HVqqkv4Fz1cIhaqcUA9bOJIgxypZuJ88g2yzX/h0efPXFzpj
Gh0xhm+qTD3bv0R2O5OykmZ03+EZe1L2QUSrwuAfddmZ7lN7xfod2PzE1SGX
Ht2d/VYdIMEtOwRgJvkitRg1mwA/xg0KtSEYEC5MyYCyj5GYoul2BXJec+RE
kr4Wbm0QVOU/lI++HUnO6dEMeViU7W3dzROUAJ1DQmWklYieD0rOO9aiB5/c
U//sMILD1A/5kcUl47HMX4t8WLGN5X64A2rMeQp8Pp6Roh0FHIXXLyZqelqi
Kce9y83yakqq0eebSwUnR++NlEO4wowXHcubgwI0p9X4HJVciNmX0bMu9YEB
jGGZa5dvzo9IJcGT3ejS7RMa1K/2TJNoilmMKkQmBeFB7T5b29U9YJVYXrLW
ov90NzAorHOMosfez4KKlNvlvxQpN1OBDh+zvtd6TPg1rPz23iSCM00dRUR2
S9A/aLoiCDumDZqtZcPJz/0MJNtHZPoXFCrfXYVhltLwfeOlY2BsySSkJLHr
WzoiYw9ZUhycHVPTE1RRVwwLiNqYFuHr7NtxBXYYtsFmWttemHHIiusHud1/
rNZQYyoFvBWG+diKk5mp8KeDzE5x8JF9OZsVCunz8ZsaCh4OdQlB+fPvuEC0
pGmc9bQFW5gN/RngYD1kMS89Uo7A+oxw0ovMYu+AX/2pN/oVxmSAEAsPTshL
Eos3r6BHxXdsiFe22e4bbcroCMJ8xyUZwYJe9R9K02oRzK2gM/R3XYkJcThc
ogeOmMsqcl7pPjXtckGmlQC39JUZlnUcSY/Qb+2vSwuyfRJyRNENFvma0HxT
USKAcTm8THVuE3KizEpxIO9UJLtr8G9YKx4vT82Ppln2A+QhPk9Lv7SkimKp
dA0UAp8ClTQpQxOZP192lNVPyGm075pm/R/QwUuTAM5HCtD8pFM6FgZ5cCzp
KKcTc0V0h5sXfymS7foGlDt2ljQPk5mZJNJ90b2HLW7Ub7LPRoOKtEurxjcv
RUvKFLPRk7yIVkg/PIsJkMUmiOq5yZLcACeam//cJsQF4ypJgaAp2+8aAvuo
uJduTnBAkfmQC64nv6K8becvhXZfYNkgthoFSYct6zUpIngnpdHN9faCWcYQ
vGYfwA2ccQ9G1t/3NG+0pGzZjFMV+wXQ9vyTBhty0GdesFQfEk6z/X5qXjLp
fJgzc02TseOoxO3MdV648TspZFxxNWMlNmRtqkU89+nJbN4YI4PMIbRIQwvp
2gUSkgss7PiVrMs799NlnQ+cPrnsL9ovP0gUoAVZ/ekB8ZQUNZPpFJX6+4NR
PFutUGVN0SOhmkvzQ7SVcKSy7UBnbs5xGqCA0OIpCHRFxXKWP9Lktmual6xq
/85QF0ZKAvUpiDPrl5g9TcXBwMnlVzUza6AdXEPHoY2FsQIDT5fSRjSOFtVr
HluXGxEuTjcapJ/5i+wZtMv2Hmlz9Pz9LxhDpKmfUA6Vqzou0X2h0Wc8ZiH5
w3MUmbXEitquRWp0AZ8g/dpQmmtTEL0Er8U6nPVwoEVWdX0PMlCn3HNz7JIF
hK6XrIn+p25T0v2mYzXS34zGnEkhSnt8APlEo5OYKeeF1rKMyFtm9mveP6s2
Jq+mSkAv7Yhu+jN87OwVdqe7crBudo2bocB6c2Yg+EzEdd2fPZ6ewQezx+rP
vqjK9Ru8J1qkZfw5vY8bWQmcTxYb9CEASd+NrjpssPToomJ7P3pT7Vl2Jt+k
RudzwisW8LWkLMz+p00u6IbtzyErWhwTCXCbsV7vejqH3Yz/W4qhn+4ETor4
9MgiUde+IBud9pvfemeO3B86xa7BDTKHvVRLvBOOv9xrt8jsPyI5/t6Tq1e6
xK0GUmOLH/kUJRutJ/joYqjjv/ErLyNrlooHX8BduCJ96wn/d9pMZp7lSKTB
W7FGCD+QfBjKuuWjrxXAX6uiHBwIvo724Hfv9y4mmgaMWYaemdZXI/op21WY
wFnIzvmWEhi+82LHnuBxkklegByHz1Rer/x6h3OXR2hhKykxfhsxi55d9dkV
CAb1q1emDeCQg/MValMyuQ+7Bdi8UVukwgxwS5K366Ai1oppRKK+clTjZN4P
GX7Hzelw552FipBD6E9LxapKWmgtqDnGudeUsjSNmf7d81xBQ52r8E4QJ2Ch
yIDeeYs0WmYAXd6X0VtTyCPiQ4eTULLuZ/z7CEeHDMjDHRAoJvxgowlarjgY
ZWZBbQ4AS3U05/lceJNf/b3qyMsA5/n1PMu1qAnvCFAX88cxt17JJrbVGV1D
fI0zCjhbWTIO/5ZwN0TD3gEIaIId1wLcd6rETlQ1KG5NBO3qa/ypwTabox2I
5UvjMUFryz4D+tnNDn/UDv9rueFTelHaRvlH7REC+RFCPfpQruirH4UeJQ5d
0hrAGUDbzMk/J21beSs537Mg96XZYSMkVQ9wknqI9dGgPlffADLhWlDi9KkC
TiuRfSE+pGF4MiTd6erhlOASmUbieHc3zDV9kBJ30Oz+z8YHoj7/zvUWizHx
qj451ekWyLgTmsV45Z25sEVbJdGhoiiywbFRVbpHc2lPebABLp68SPW6jTGL
Pfg/x7ptkLJ/Gn8Gor7VhMFb9pz056Pm+KqNbmibSPAWB5KqRuoKwwv1UOar
w1fAFkBUKp58yqxD3QrrMXcE0XKZ/YHm00Q61Ob/iv9fTw1cVFGBvserzm6S
4E0alP53xaZ66g92M74MK6uhRH0lf7wTpycONTKVETY0f+DXRWn1RC9HHQUg
P3v8kxelk3oFPMMaKnKsrl+ny61yYdWky/9qc2gqBZAIvyobb8NgFqXKLYYb
JGUV9I0kfXHprl4THrvk0ZuqS7VSGCakqCsdtx1ahMCrHNPrXvflIMWlW2wy
LWESv2zHYWLRBEuHR1w5s8cubFcuC5MaeUmTan4WnrLLUcMJ1e2ZhfnSLsDY
XXTVDQkduSrey2jdrirMSr1VNmW9AhYeP9ZGd9+4DDufiwCPv7voqDgE3DR/
2V03AOdouxpiP9yt1e2FJoh9CnfIlrbTKUFzpBM08TzuCLcNrDXZLgmekcpb
0467P3W5oTonFkbn4URe1rO+AWUnZaJKNh0tESOSPvQs98efHyIJchpFdExZ
11qkmh2r5YBhUeaO+zf+KX/RSUxWMOGxuRmOPxMGZFYxpb1Q3VucdZ0kM8F1
8yfaqNh9UX3BR5y2NBDxvwnOMIPqlL/L7LCUwT9GRh29JiCYc10+aHY+T0e7
CH5AZqUAMH05NcKAoET4AjEv1AzGouZIjFoklNfI4stX0EgAcwF0/KCEyNUX
ZKvd7HuMUGyoS3AxDLGj3DDOfBH53SAU43HpX7AMdddHIosL/zu2OB2mZmjl
D3AWmMwgP+zc4Y48E3PaVziw7KTDVU6ttudJgxPNrxuQ5Ypol+em2UMJ/K3u
1ObisEzzAxFDV8krWYbPgb3+5uiSmeQ8kRWsulcqXEGNGGGyOCYTA9I+W59X
GgDwUQ0OcTQGi+tBbovkKypZEOESYn8LREksfdz9I27mskZQQV1E+keLufYS
hfNJ8QLhRcq8eOajVpd4MOnGPVtZU8FHXyzEfPoHm2Xk/G8pRORyFe15u6WB
+cpf5E12CFZe/+1KLu2eNXy0dNYi5fokI2FLsAgs12FFHoCAKuAqaUiMbGyt
I5l0wphVxiRXbif+CoWxqHC2UfY+MO9EeOLK3vqd4EKRS5xNwCoh2hn7vkaU
UeQxPfdeLZZWB5dYb1MblitmNjdsnxt9ABq/E5oop68SJC3Wx+bSl11ZdtEg
ypEXK5HqnqASGeZY1zH4oqB7hyjeKFL5JSTHQFnef7R//gTD5wKDtKyCCJ4V
Bsch89cQ1hWv68Eeuh91KQ6rLj9L77ZIW5N8T3zTn8UcB1h18QoFKCabbBxW
IptV2p6qe7/+m/jFZJ42E5osC/6wGHc/Z4YTRxI9O5+mmTMBr2KCDF0Kc4cL
yAEyF2/aOqyX8zGP3SRzZOnwgAANqHjK8oNGe1aUeszN9WoVuz+iozXheCff
VnkDm2AyxHQ=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Kttctzi5aPKQ6vg9w+1g45z6Da0UaxXtt50QPmQzmLiVao+5Qg/yS2eSRK3c1uFoxS+G6ngDcAKHm0LGGibx4soakCOjaaRTqJmqblCXBo4qigRRJU5sOpNJWGKfxZC9LZLfFjqN04HCQ8ah5FN3P2yNU1iObRgi2dEkx758LbIsGmsSUmn36d6MTHQGWCnH/AC+2pgOY84Iul0q5eg7DNO6RSxNOih+2JmnF8szbMMRQoiJ1XzkjCC+oSzVQgOUFWmdwwilN3HWgclYVsjQVQEzFufAadR/lo6PW9yLmgxUKFtXGNfRnvUsnVEHrYmT9ERwb+6WSBgDgBRLmFB6HVCwY4JlAjCpaP85NptRyFis7ClLVXf34hwO09uFkcKiWBVXhJpn6484Gnwo3J4WCag/TTzwZZaAY+R56mFfTZ0JIkvdclFIufZ1ib3vW1KN+34xHl/zAFXfK6GP0xsjxU52sVQUCaEHEcfp8xFjQTt93XCEfzA05eWqwhcVWGjvvYQB5Gnt9/vC3hdGA37u9SyfbLzNvj7ZspPWwCvbpKFGo80mUEJUePBQl5IMvZfPF3cbtFHfJYWwLo+CShvWopqw9XvSqkSeWNVkzu2BE12G72YYlYLU4/Rfq2Fxi9K++1Pgb3plupvLnLrZMPz/gWWfik18qd2oWWocEnSxWi6vpeafkRuE1SyQ4NYxcUzWlts3rsLI7baMCJER8LkeGgobKY9YB3YfTjTMA250cgaKfbEKcUkRb8iP8spRMnGYUtO+gMRTzxbybbKX1/kHDxu7KeEZR70ab2jnjq2SPSiwDkHwaYTh7AVGeNwphv1W0pGfy1CtwCIekue3uI5tLbnyVG7qtI2+mezvVtX73vBkf+rfk3B3h13a3aNrsa+9bA8oOvnMCllY7BUTJkkRenF3Qe+NXjxZx9JBAyRWrsPxJcycr2pVxEQj0WE34p513RHMVGRtkGCHZtb8SedqLxBUdc3iF3lvpy85e3kUkaWao4//lHUX6Gn0bHmem4c9"
`endif