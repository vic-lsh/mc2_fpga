// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BqieFAgGvmgEx1iPOlpaUm3+o1CR79sg5aRqgRyeL+GPf9sKeMyFrnDtPbWN
fBeHWf1C48WiwieRPe4KLdtNhkf0oLifQb2V/Ee7DS7K1vbeNTyLFvwZr2yg
AZr5zNwcxENaHhExUjHXzfJtwGagcDa4kZk7xK6nRbCqjcaOUFeeMQtNObmG
FNb/FBVqv6RthtbHOTsjU9I92nl7wdE4cWKKSD0l1lOOCCkhfJ5nJSPh2MGE
t7RRKLA0/k26/dZHY/wPU78jnukbJVr0UmL5hOxD6WWUxaZM3uTEQh9Vuqta
AwpU3viscy4BR2opbVrSIIdVSOQSbdArmbkcQiaPYw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XO0q9Lz44VozxAJBBmnRRgh89KwUM46t3CrkM3YNjtG7ODWMIDCDjJSW90Oa
/SfRDcrBGwCVxwqma6qPjiksF8SfCqc5w8p7YwHB2XP3tEVRb9tZtYQ9QlsH
+ZGzVydGl2XBQG72fWwjUB9CsNifuKVraVCYjiTEXdfIwrq5G4BkceVcqStw
FzMH0vLZeOHWKITbTHdz8UgtyJT5sAvu4oBa97sc0lX2q86lKaXJMq3dFBzB
TgXUUpBgCPDwJZKuV40B7aIv9JGSgAsLQQNWt1s58mkeUWjytHe+FS3wdWB6
gQhmut4eDg9i12YwIhS4DfB/xtbr3ayznYEG6mnVnQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gxC3Fu4k4sAqgiZEI8/8z9lAEs/QatfEHgl6uHcQ4xRFNkBhUcyyXqag1SBv
W6AjEXy9QRrtZvfobc3rvsDdgtSKfCGMIS5p+RC5W0LGWfmwOiqX+6ge0dUo
ejQcDJn6/CZOTzWhWOH0JNAFWhJwT1yrsQUe5G5mIzueWCBQ+XMT+hjf87Le
2hTRNNdoqk+7D4Q4BvUsBCynhjvahoGx1VmZ0k04wG9yITmHHbHxOvRh61Ji
v4Xs57kZPusybyd4orGstnSj67r8gydl29vGTZzySpZa8JRk9Ei80EiQP9Ch
wOQKxqqOVPV7DFgcuaeRwlB8nLkis+Npe+PBDAf9Dg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
csgco3aNjMUZ9JwuxoHWKIrrFsbT8y+Ozs6RH8wOE+SC2ws3lHQuHp/n2J8v
YVbzX7NkObQU70JO5AHYOLBr2mq8ulzwQ2mqWaOt7jVfKRCdczdHxnUBs9OI
XlFta906VNo7IkB7ZW+DLqZf67o1BAF4OosAtJ1eEdtP3jFE9TzTAJjqU7ss
cdXqMegiquGHxY9LXRnpKbTp8kpPiKkNAuEIqXJ4vDTLmUQrXW0mLDoRjDMQ
DwKZyebxfEd+Vs1r3d/2bXxayNMaOY6U8zJ10np7Zxz02VP32zijUuIo2hNK
SUWR6ehh3RL6EupHUaQR1qRBA18v4516MnFpql/UaA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kmiKr8OrKFTHH2HZD7GKSsC1IBSa6r/d6GO62IALRBKulx0kA1u3KGssuWEd
5tWB1xBqTSLEZ6vAUFuI1sUa5E59BftJatZQZ3dn9qq+Xa3Qw5MMQ8xFk8JN
n+jdJEfS4xAf8Kb+VjZYL6N24aQoeS6labv9qG+uL9SzcOg7MMk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ryCNBzQQ4xsdp9kCtrfRn8uC6mw0VOqStLf178g2xE+R5eTxYXajZg1F6azI
BZkK+59IxuLKCaQZWDydhlK8X4x7ko6Av0rV/pJRXhxXxTlqKfgbgqDji4VV
mnFN+z7ZU8aTodEksnd+b3YSW8X5DkhW7TvwNWwFmo65ZvMTw+KKpWvqOcHz
viAfbPMtPbg5hK2zYYlBbc7eckqJR9VndYSmZBUXUbRg9ca+9HhY01rqBYOM
6qo3YPK7N7Xv/I1DPPmO8eB+VGUqHMXh3cXzCHf1a3VADMAhQX8H+iWgzhIb
eMkHvG1BrnAfWjV/VgH8t2/cn7F25YO3dXmQO9IuwYMY/zod0HRwRnnIvdoe
NMIA5uRvyEP5INFFBxqqez1Lvx9FR+y7YVICxH4AuZeYR8GZTeFUa9TvLnnc
W7EnVvAYZMtMEkmXw/Yu7M/36JJODL8Lz9WMVcOSy4gnYMhq9Hj240hpeOVZ
O5fNwarwZK838YFHGFrxNj5xssG8pypw


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MNfaRWxHHcVwbfPvSPLRRGkid+VKjlVOs1wi+ml0nClgZ2Kzoz0akfJyBnvW
IG+y2mGDA0oJQLB0Y7FWY8p6mLnoPFoL8wZjvZ0Bel+WGITQc/ZfjXtRPXly
jazzBcnBmbZ79CGF7fPtlWYEsPjwfOoUwdSl7XOTCmxFD4m9mN4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PebzrVndEZRIkylbh8QeecWj+TPd8qPmg68E/u968OzHzLUaPLiV79vNz65E
aUR5JpuwgS/a9rs0LZiBDcWQJADMRjDgAQFXLy9dv26ds5lRR/n2uddl+435
/R7mPs9r+uKeuBMfNtXjrtVszx+NCzKvij1zTaA7KHVBvRzSaOY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8464)
`pragma protect data_block
o3udcJDyvuoQfN6L1XuA3xz0NJmZ6gadbxe27iEgxfyAI2+5aTM475xSSSi0
ULpYU4Re6aL49XPr+dMi1/Rzy36xngwQwn7H7zI5n39BYti7fQpSZqVWDtuJ
xkpIwySagdhFfPyGveBNcW5hZDRpjZSPjaV8iAwACRV6EVQKyoXzWtlfy7S6
v6gcaiBnd4PQVkR9IWYmDUqUD1Ja8p3XwsNdgbdxHFotQFVx5oYCV1etrBVm
Ydv+ZCLefEoC8jNButogGzxM3JwnHwsridM+HoAiW4bLskNAmbnMwOMTOUuS
ma95UP6WrO0hxUaROt1B8lruA3LloM5fC51SIC+BYonc9WlusOl1g01aeYcV
YWIytu4TYAcmhvY6bYoZgp/Z8Ow5sq2ro6aFQWg5KSsxT1MRu6rEituLNodp
SaSiHtpcOFG6zxafcdhm1MLLSWDdeu8d6lt5su5/9lDeXQnUN0rtn4INRQLs
U1uVSH+KZxCMS1YRcAXXzCU2cbHCTWqY7/EMMf83PfArpbID7Sc+qBYzUDx2
hf9E0m03lxsezaAQ2s85UhViir+a7ex5hoiVt2oscaSjfHmgT8XeJxzvh/Vf
SBWRpks1SPAhg6vZSSX/WQyfJlUu+slAEh+XzyyxB413iIwUGhZc96GHs4Tq
ZSmpxa+XRM8m+hQ8Xz/JRPJfmyc1QyojTOR2KzPHIXSqH9xPVGRwjv75swie
kMBVgTKnik0Nu3CWzgV7SHPYng68cCP3Wcapn9T53REJptTAr6Wxm2jszhY/
ThFON7aCFz0wfRFJwC4LgQoxkvGoXhFCp1wrN1o67eCvIpwvu29hgD9r7QI2
pDni9wGAZFWjBZlZ92mqf/Kg5RtpIrbFdDZDAHcO/VOntD+2WMp87YG7pHAP
ef5tScwGW22yQSt2/+89Yq1I0DnSm0BbwRSxIlXXKoDQMlmuJqARzm/x7mIT
jT+6Kvk169P+fTQKbQnE0XnHCSokJyFU9zGQxehwjSOjWnaR8CU5kkC4SqE3
3srPk6vc4k/qtEasmJEqQtSLOFmNZoDphLYtWxr3pyuwAipcp5r70LEOdjen
/Bi0CThigS4aYdnawJ9Dv9+KDXDX9FtaRtc/VW5ApBAbZbL0YJfp4QbiWbjb
c5xB4gWxK3mjFSKbfQqhan3oJZAVeeGW5Ey7lYU48vM28ldylHIR2WpfLnx9
5e8BUfvJjbBrizJN4W6CNMLVeiLxGUP16788tTirRYVv/LTJ7Xr9VYl7dNWM
RAycPmMNBzWJOYsgoC+JQxIz8ABLPjC893kw8+oriWT1EWiHTPEjiWYgIu3N
Cz3dppbP0LwP/uJiox3i7dv9xMOwIYp1aZ0QOh76di2Kya40TDU0zcOUN37q
q/7RqbB3fi3fItAiBSyy0j0Em0aB0cOW5i0gCR0tLmw120G2Z2yKIzprhUTF
V49LwzI3UXgtpZHmq4Zn0kkO+E6n2R2iqC2AK9gpvikplfp5unnzKYO5EfpT
JbNVCDG0DN69TdmIQiyapmtdKVvAPKvlNJo1v/lQdDr5NP1UfDDOjll4HuxZ
4CVr00OPKOHgW34GILytkm9rmDztzBtDRaOasFwS33C7cYAYmDYIpSdyDUW6
pHWkvxqHwPkIhdOexRS/AIGc211d5bFXktHDCLsNpeAkcMPTPTBsxqVvlGPa
LJ7RnfgGN//de3dnsTPZ81vhK0ZeyxlfdwYELHpM9LErR1z2cqhcRnCCpDdR
ob8ppMVexka6URLuUHrSRG0MWd2dUwjFtASYKXYld/O7oYWVXSX0OkzJhbSa
YAHuegoeYps+cnVS9WsG0q8Ozj6RLG5NEJBc1ImZOx3tgal+ORq+UM92wXFU
POdfOQIUNWV/gHZfplq2na9vxofS4u5QKyrq+g+yBijSYQ3doljdyihvy7n/
coMm6ilJm8sJVqor6vBYw5dm4ArBlb8QzZJ1xQpwfyIYWJqOax1Pn8tt7mvt
E/1f759xKO1bIvVj7hprMpvco8O0u+N2w7OKEfVJ7xMT9J0UiSSYmJE130R4
JzHyKeewW9z0w/YHIwT0q7WCAaemCui7dZcZfsmU86iBvkY7js6uNQA1f/Mo
wiDhOmKxxZrur+q4r+ejxvpYYwsFoqg0CfYtim6w8na3HUT4+Xe4NsOM6/ou
GM972B+m48t+Oj3Hy9O1P50oVlpj7uv/oDOZPKL6ut8bEhZenIm0F0qBAePD
lkJ+FIojVhN2UbYj0UGhfGV1GImCx7t0T2qLRgivEO/A/IPeTkiU0TOsDuOq
IgRI7DgZspkETlu7kMFCIJYr89lwci5h9Vci4LonbyrvuppmfIL+gwWhdMd9
vMH8va1vDSDU0tqYqblc3swLiaVDk7JhbibXxvzONhT3OPpgkBNvOpuXXRUM
l7W6EPJTYzVGow5m326tvX+aWq7AyGI/RS8TJx9L83oCh4zNtXwKUic1JzRR
XsGvkF7ZiggugXCP0Ioqd09D8CsTuVC7TFxClKGoK+wqY5zPD63igJPkw8FQ
AbWJ2uoT393Jaui5tFrtrG+zy0rB7uZWoi+rNRAuafswvVNS+1zy5agQS4wa
ZxcPKbSTrgLkFE6nOLICN29qJ2+9UEW8bIhiaZaNHoQxMPoWVZT7RrZ0LJ50
zsoV07RB6emNtWd4wxhGP6wOYPFYF0BUi7G+LnNZS83sihhRa4uV+2TC10xt
VNX67K6RbZGZG+PDlb93yTYG5ErW2kork5/9nxWUjcrYLE8kSr2gglME2VMv
spGh0NvMLlMFky9NNKTreeNIDpjm+cITr8qXUwXM5cm7PqTbX2tuiZCCjs2e
vMbwybetaYKaQASINmCssnL0xn/mGOuPq+3HEXAFTWF4lWzwteL1F7jKhcUU
tUYiUFRoNfehzkXkYw0UVDrp+I5RvPPX/A4hdSdnp9WqUSSxS3LBY6loKbah
kKYIv+hvNJNCYIy4B5HorL1Psa2C0z5+2p5MZTb5aIaHFzt5qAEn4r7clJnX
499Cmnkie71WBO7wnwFh9gZ25TNlOC0AKRYy25YXZZN19RLX2ohIv5J0jbka
RAux2jABIDNF5eJXWImmj55QHlxjW8hjo8M+FSjjPg5jPIVrdSxU454cuDTd
R3OMYeYV93TI/1vkYMShV8klvkW4+iJHtnPcHQsmFEqQ8MMUtPochaYOmmlq
wjUO1+LmBxFaQ5efrFKbpPE3FoUs4P1NbzvzmG5XfRRF+O6xt0AxEnn88tys
kfWNJY2amtcOyXyCeY6lhdetCTBJmtnKQp3Tm5DSruynB0ZpRh389xttP3jC
yJuVzZLDvMlP0B38IF5Y5SEy6mFWThmGutjumh0t749fMzN6V+8MIW4OclYx
ljfVKViwHVwOZyXrslSHMjiw+3rHyRrcwLC/mMTsUCHGSY4LN+C/OkYtbN7y
S0KsGD/MCD9yRxyL4CIScyhVHQSwZ/Udpl/3OIxxQ8b9o+HfLJMOEezZpDe+
fLwOTKMXeweRE4ujRae8byARV6Sqsn4suidAPZ2LTn9yJcayjGwMDMJFjT4p
xbqK4+anWsCUUYRALpO1XnjwpeYie7Trx9KAldNuDhz3vqHuqZllLNo1Vhof
uRjsEBAVlxqza+0kcDLzwl2vq4j2dbupJn5hk4n20eZH63fjNMmJlMclY5jF
IevwpJ7vEoVKZ7CTJrc4yE9CGUQ67c28Byt7Hz2SPsfs2XVOWBmFJ84Ttxgk
LZMIHMs6JuxFEzL0wvM5QyqR7SCwmzvRYE83gAQBoRKYnFooRrlEm0wOp17Z
pSofOUn9KdqZvwiKR1vG72XTJ4QmfMgEdpK0bvbyN/MAkmpp4++B087OilqN
mN3JaYPG0V9i49jzt0v6lD+3YVIsnkfEHGxU3BUdFxNwDlhg9y/rpoWR/P/+
SFwIzk0akS9TSWo799XqdP2tDgNbKJAZwqDwBeEWfAjuf4geSrBod+HWVjDF
KsBlMpp8BQfwUtHSCXMIQOCisWco+N79CRXlbgGPZthQrmpeoyQpYAhfQaOY
ClIQLnxm9P6OQnNXKFZ4niWh+gTOq+MfJrGLUPpBRwhNohXTO1+P4dzITovQ
tabjhX9+gpi38pTgh387xzISRAcpwhneR+lPVe1uO6i/gY3d1zOHM+FHstUz
1CxxiThBxoxzvMY45tVqK4usBQrJosxJRf2+6C/GhRcM2YxGPuGgQBIr9hN4
qN314PygEr2pQ0KiDG05j49mM0fK3Nu8yZMNuVmLG9oSNz44Q2mopKDDSX3L
yC1uRQ5XuxvVtuTriZ3kdp3+ilNmF7Miv599NOYb5oYnGKVw+6Iz5jaS8fhy
LkTnvBL2PzdRfcbm4pb5Egi6JwZU8xGpgRwzr9R8he7haotFBCCl9fJNu71n
cqULwTCCkbIEDq3dpSKqcFyx+XwufiGpz2IMkq05EKGZ8av4U5nQ6CFoi851
irfhpaf8ufTOlciVBAFLhRNo+qDOoNa92jmZj73SBqBVs8yBt6daN5elnlPn
K4w8zknGGOXvVKN0ZEg/Aq08Ht26Peri7rKcWcg0Wi7UrsOFbZllhtRSP/OT
t133MKeUW/vEaZtdqWc2a1cPZv/gQFKfAyedvR3HE1GMAq1pl47ru86oW8lr
gw3+b7sgg6F+HIxHZ66Jf9i7RFdcUYIvTqGZyUPKKgCHs5soVp/wgcwat8YH
mnSe4WqpZA9mKeceybus3XWO+tEHLET/ep60XYy3VFSphXX7n19pRXVaBfvB
ZkUSZeT2yjd4Z/zeXtuivQeLEAVSzg7LMQ9cx4BYt9plyp5N4onovfqZ0LSj
GzMzyqLzuZFoSzVCfhdqZqdMFQ7mWM/hvLEt5lkV0Xhmj4Z3+D1OTCd3j0qL
Do3vvRYbXi/S2NRddX/uN8EyMcxCANnttf9DhWIAdxcT7TlaoH1sWDLDDGpM
gSVDNp+YJaYVjjpfQuNele5QTWasTFy6ze1rb5mbB07LUZx9bLN8lfCnZTv0
89UDY1KDEFBA6+/wAAGkwnhWCdb7hSng6ie2arnv7+rp/PLUTOQ2OkXMzhDi
/t+zI1t2BeNMDxfDKrVFtQ3+k00+UG65iTAAkuqI/G8kevNF8sNI3Kagyjz4
lwkqd6te9zhHMtQ3Cdlx5nmbROocrENgZnB5q28mLi3k0ZFZpsr56e1sTyDe
tw/IbmSbJlJbunK0P0APhI74SP5Na8GRnitmwRLCpxXXHwcU4DNRojGcPAnT
4xvrp0YLsjo4kZIBfdzVVbGGxSGk1EqQyhKCzmE4SLYp4az0Z7R/Qph03m/t
w5xy+B7I+6BmMAbQE+Q0PO6AWesdWV39yVCbIPTbPJvH+PJ50Mz8/JfNfAP+
inv63fhdBFR4dC3HhHx2enW+fHBTKsch+k6iX+tm8gyEJewoSlmMHsDtEmfz
lrAlhWuttfCxJYiImuXd/6Gm0Q3eHimPA+pjXsJbTweFPCQjMBOTagPJVcQb
cwc5kguIghoBkfOViD3ph8oCNrMM7AbEdqQUl2f0P3KWgfFvlB3aHzcW7BVP
4yNRwPa2wT84v1N8LYHqeL/f5TlI5ZScSltWlM8aDxgc6VEHyK4TK6DFZxTb
q5neNTbmZV3I0Wb/0slV+T+1e2b50K7JVdeejENWT83XZT0aOlhAwRLc/buc
E5jWN2rOR86/TRrwYqSGdNHIF8PKP7L7/Z72Qh3UUpBxAhaRSRP5cY9aySah
JMM3cybxinvbnDlRxb7l01gnv1KzXLHcHUC+hNrsrVpn48Zes1HHiW3oxrkf
gXUQNQrZDZJMSipY+EugoEP4CYOlgHVX9KFvjaBSkBuJyqQvxCEq3+RYaDuU
Y3hadbdwFID6jFDNNSshmA/7lsx2Q6z+pAiwjW4AYiTux8/B2KH+eRxz437F
plMg5le9Ce3GOU9MG7Sm33qSW6qYzjlHG8OaPQXuCVR3fG9edoUnRivX0Jht
8him8WhPNaE7CYdjMhT6RAXrL2Z+pXG3pzlBWepAa57JkKAeIWiV3J8ry/1u
RWiKC4gDug0qhupHdAl1eG/im9af61K2IiJ07GdH7JLvOtDKUtka4JF7n48N
/90wE74I6Tu8Xyt5PChMrucqo1v0brxYGQpgTYAwn7IBkeslnXt6ZiqDAuUe
uHmYQzMFKgMnWtbN7ZvvV8T4Eo4vk2tOW6pJgg0t3uH0u21izSzI6yJok1ze
z41JkMb2cb/AJOAKkPeq5vVkAIk/Ys2uTexxYFYszhcHC+aK3DpdgMfC9BH9
x9/b66PROWwWmmXQa6wz5PNOTQqpPlv4NOhswFVFCm6Xj1ZbpZfG4odQO3eL
jU7JLUIAsiYoAgcgt70Wh4T2kQ5FIIMn6rAF7D/vkUqd0hMhXcfAiPTRi5wd
rRhzQcv86aegb54x8j5LliPB+SkMou+DxNxwvqD/RBIq/xdlVoJmQZaX71CT
bXPg9sKX9zfVVH4K8rFQzN13rhLUCR8UeVf5EMz05TUtlG2alyCQ0EVQwIXl
a0SKdf6lxg5n3hhzFKuZs/b5t6+Fm6nQULmQJd0PRHpKtcBgZc+pMcrC8pTt
N4otmmF0Qy2R5WPAPPtwwm8YbpU49/U1XbJGA+6syDus3J5cNw0xGpMzqUNb
xNk2zEycDycAZ0NRoasNmQEDrlM9G/3zhqQRSwVYmPUj+SAHpNT8ReDce9bj
1PJMhSmz3sGUvQXngms7SwbhHczS8UyOd3F+RNKD6Eo3WD/lwnQJZDD5avOM
tGbTfn8B7pNsV0yBeDjz13QpXdtgyL9D0cCCe4bgsVVPg0nybxvyncR0WtIF
0kM+YQ1JFvls8VpS+RqnncPdnrQP0pu3hCFB0jQMwn/Wg3CBoucPn+8TKj7u
UDPp/FyixxniBZVfqNLMrrVVccxtuNEvhaoFLp93P02z5S1Y+45We0VULe3Y
PnUB4c3/qL1yuaKFadcL+eyuh/qcX59UUISZCRwaRiKgOrnlhtl0E4akFupO
mfXhouKaphUQzD9YaZDTYJygg1rvyEmU0kZUjeKnSAeuoQvqBkmjIXHcdHaW
jo03PkAfm1FdhhGORyaZjLQkefvrNyObXyPlAV3Z1fsL/sJDqsdbcILb4N4o
7I9uLdzkrZpA8FhOeMRpjIt7Kz0fAO8Aa8KTi0ZP0XK7gjUX7UXPHXCR21/d
qDe5HVd0GoiZL4BTl7ncweBV8vhIwkfZTFS8PHRqenfNwNL/voI6zcNDpLe+
vPusoJVPRMymwXcWqMt5oiL3HGIyT6GY/4JcJhT8HoB8iM640dct+FnkdPOq
Jg3/RmU8znWYhgoi6Gw37iqOFBwzWrARqq4sXY1ZYr8AsjsFgwVA7UvEGpx3
H4QwmHT5TpNyvkgtNhSPwllO3I/jRaVXyZeboglJxUWLk+++TQjYtZF39ib2
8+IvtKAu3XHQX5sR3B3ItfDftgFldbKDud9UIiln/rEWUpLQsdZUyVNNXPGQ
kheV7gB1lXPO/4rQjrpkPgLsd1MXG2DD20wkZ9EXzrIc8KXJ5WSbyulI7lIs
KVCFhWtVhDNUwnzSmxCHdGmjLJiJ5pQhD0lvSQhCKVAvRUImCW5+Xqsj172O
MAtEilBHqdTBUycQcYHqnwPPw1s6Itnn86+fG0C4XTyOp9AeyON2Ad7HjPjV
QTc6YulB6La7oCXGCfWw3U7XKzM34wo46wXvaSRkmGJ9XQhJVS5qZuubuxv2
2+r5o4YEiSkTxxds5RyKzFY+Wz5FUD1H9qYKr156G2XDdCIC+IFNahh7buUF
2Z8kKcKhSH+U5sVBpKmHvq8tGRZncbkoS/B7iG5r34GYbDGDqZ1d4A2t8JaB
908vtJF3HxfdnbaizIMBN1mFaYo9TZHpioNEzpP111MJiao1yD7Kzl6Db7tY
m9jxdH112smd2J1EM1SamU+tbaqwsbgRn9/Nrd4aPLI5IBZjlnY3fx+F6kRP
7qNBKc/FjT+rir1n4lUoV3Qr6PJYWWpZXYoKie2gMQbJFu8AcSW7Tx7O3Lpm
t7giyt+hULoVmSNIC5VHTmInu2A26bFCLXxNRdnUMQTTxDMykRTF0YsUIDym
SyDWA0SXIg83GPPHq0RYQaboeV6WRXcf4hCQCzmf1XsQkrDq+y9NrfhL702M
emnVTfeZrpEuksO8X+oxrSFGKafJn2ONaHyKBKHqFO9QcubC1jpZYA/U9tij
43xNu1U1qVWU8no3PXgxY6qKFuJ5K90VjVv5WgqMI+BzTUNvVvZa74YPTrXZ
vlBnXevS24zmGIUISPGILYm8tHg4gFWLziX27LCGUkvo8gvSfRAVBkMQKDs0
G0n0FS1OEGIl0dlfzWtdbA9HdB/QPzwtea0d3XDmUYLXE2R3gL5VNlKKk3Oo
4zfjFlr0aSJifRJxz8aSPaEWW76xDIRTgTLriMpTqSJ+NlelhRWJtqFATNbz
tUbg7ZxoLNJp+6uM2srlxdAOux5dPlN8ZH9i0WNBFLtTbhkcpuXsARdVLwst
czdV7Gh29KVTRM9FYXzKFyLtC3EkEUwGyITMswaj/nlXG8ppZVWcE8m93Qwr
TSkwmpz/vsbPauTSdnVoOWKkniScHlGR3YZrh+KKC/BUGJWEu1YvQJZxrojl
J+N7KlERiN97htmpk0VVc9fVfjDppm0Wp/XVAMcJM9mctYJuDxlbsUs2F109
LrC3C44eqN5MtgXn/K0ls8r3734NywNGBlyN/D+rnN/CVqgkZ1tVsaGjSFRw
HJSYuNFQ/JyYSdPh8ypB1Vi3kfAyk59Q0A7Paudup393FLJFc6ezftPQHPwL
vwW/Q/OMe9sTV6SfmJdbEIR1fdywM876Hx2uDNDqm4Sn5Y+g8j4rfwZnNrq2
WWMVsFvxJksOVqwiiwZG0a+xs56GUX0HCioDmlsxQrqT6gp8idC8aiODE/Gq
axOD7nz5QS6LjaILBA1aQtxGGA7pXkzPk4vr2sfWMaMhZqaQUM35SVURI+h6
kyyF3XMj36oMXT6dpYOwP5i5IA0UR/AlYkufyOvOTkjp/XuK/d1AjMwWInfl
A9k98M+nUx6TtccKTb3GzK6TxObgV7tnSDRWIag+gt67mgnD/1XpTQRJaqu+
icZEgELtj50KaeeKQpYwtdZeIl1pxU12Q8ZinS9mN2E0oFs911Y/hvt8ojls
t38WZO+0vaxqvgeIk1LiepKvbD3R8hzfNU62IvYOIYztCuSI2ERuSkgrJgJD
Fq7v6cOXeNUla9DxnwoExbKtJAADvwsTa7hPi9tg6iQI1/GbVtblHc6Ho+A3
8AFRwD1ZNwL6KyjlbCPc4BytvXHsDqLu6sMlrltDUB2uYgD6kOZZCmk8SGDR
qiUa2o5C+4ZLyvvyuAyKiQ94+VNd0Z46dJSZiV8N0m1KtjDvD0on58UA9+QB
PmNkx6qKf3WNra1SUzcg8g1URrU4zyKADRgQdgftacMARunKgCSi/FmlYsAJ
2zlW5L2YpF4wVGSVAHlS+Zq7CFgrO/oQuCE1/DAo3UALGjsxyQA3h+UsyfF2
NuW5lHpfWPxoUIOB+yB6EAbzVmOUVD1P8NALLvrQH1c6tnaJjdXG5phNaD9f
gepBNvZMowttlq2c9Co1+MJDw24xd4UYHHW7Z6AtyNbd8mWvdcmPKK6nvBKO
louk7dcsAIS0uIywx+zhQWM4eRoJvm/lmxeREjCUj31eHcHO8aj1Fu0SGLE5
ARyOz7COVROcmQxCSCuBveZ3AB/1t6SjX7oZkMFGjv+DJ6H3v3+hL7oVe8St
3rkQANQeAlishMmTDaNBEgy/LWOD+DTclrNAb+xBdtfIHhflCcSaOvU20E7E
rKeSCD42YIqVRzm05SP/qeoCl19NzaZkYiGMUGZdRUiTwBTEe7u5WQcqefxM
30XB1E9CaF1j2q1iD0c3RWhKzOZAoGQsBL9kx+UXzKtwqM/tun0QfFVhzG9D
gPt/AOCOlnKTjoF7ock2qrqw0yCJwHAworM50avV7PlYynpf9qgwVUdDjnRW
AQkfui3q6zaWxkosyZD+4VQpxOvS5CO9fWsJItrXk5k34bfCbeUEnj79i6KT
WGiP5kihBBLdWB10i2Zy0LJSvsd1+Kw8qxs0jf4rG24udIt5y0jVmJVZ7lQZ
bSLxqYrpgMXpSBZqtsNYZBQtWJXgDKWAnXInmsC++Yfa3pLwH8j66GvSIbX2
+DJ3q3q9UJtJiyfjJyzPMlf25M1aNTp/5CIdulMNH63mfpfGLxTb2JP6vXy+
69j2pG+Gq+0Y4+mojP+cGyi2O/tK11fLwYfWNOAZFovKvQqE93tLxuGx7xuk
/kR397iw8nzDagnNVRwzKWnZQ8o/cOzH5akx+nIcX0fvdz6v7GenLlxjZ8ws
d4f2Qj0P5vP/4f5N5LW59H1N2tef0GdMIMPjD8Wu+lQv5S0GV/Atp4jk6T3z
/ytjH1vdSnoa4tgJWREdZWKa+Y4VA0CcR1JCney54qTbrdhwyWGg2Xyw407I
Z/K6PxiiIc9MlbezgtgYMAQR385hMAJ7CIu2lTbbAvZmVEMlBs4nfpWcVzXD
XJjpwNxb+7ULZwpthFNn65zb1ZLQjEFRtrBDehCl85aDxwgg7vowupbEZ4X6
jvQh0alSW0SpIDCSapscZwpF+LbWWjn1KvxveDf3QRVkRGZ1eJUc1LeevXKk
4YFQkvm5wfjz01JzCgnKt1jmT10WaQmOXQCSG5nfclQHif1DYd2KzI6pZtVJ
ButTSxuEZ6Dw/QogEndZXe+7nEFd/SLpqWiuAo4yeOuRTL5QT1+oR9reMiw3
UnE5L0DdOkP/8TOGasM9stenUt0GSJ2zVifS82j1/8IZU6uvBEqxBjTiTBNT
HOolXZQrTrGTZWP6NRQf4+NwEmSZbfYYurBZ2+RqSUGLe4GwhxL811rPpU5t
dOH1sXp9IPQ2zNUElLEmD6vlXwa6G9zMxQgVknlP50Lkd4/jYCz7eNqjNZn6
T4eFhgCnFKv1MZBraVAc62ZVYfwdUZSOmuRy8FLIkxVoRtQDfm/2QZCOpTEE
4CYkNCdb5sFdHAdr2XYJoaE4rgUwAcAYWhSO3khrPh3spRosmjeUku7FPLUt
/3pmCUj6qB2aCQxuAbsjByge3Oc82kJSO7KW05QhqM2/0bkjW7FMvG8kOvmg
Rl7osLe/RLHBYhBi9irUrhasBBtyUraE9p5d8jHtBz8YGz+Ha5sGmGWndWpo
L8Maqbjg8j1mqRjFir/CqYNrDr23+kXfG3MavKAAimHw1yUQe7DVqSpNO9Xn
LXKT06klpSq36fr8eebskggfwLCCkkeJr/Ghjx1KDTjRhEKFMSUyK1O69DEH
EuthCA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzfx369IR4+CYTdta0EHkUI59ceVjJ6a4SuHeBm+oFsjseaGDKiUA1FWNl46VKVnioG+TpBim0lFT1u/ZWWEdL+TJaLAaBwP/JfVymQtJTe9Qlivott5kGfxALyNikbZbJ7FidsqT88ps+j4FEiSQhLLjOgOPsJQuaK/oBYZb3q4IMc8tB/FXfgIu1PgvoOd4TaxN1AFeVYL7/AmOqfGyIpkiH4ideH7qwKRLVPxvh/AHgNrcvSOl+EhcVShKfds3e0zwRVga7uktO+uoenUhGWAggT/nlOepjWihj6ZIWVXzSYAtvp/Y3asfwxJ5bVedvuOGH2ODMWGHg+CCWeBGXJbC4psEfssBgE0K+rCGin2K9UthTQshw6WiTkYGChI04IF/KKVPgxsWON0ejdpG6o/XY8X57UVYWzlQwuizYU8I5iXA8mTVnut5bfu3a8VmNkpc+b0yjd+XC0D71J2as+BPQ9+OktP4imTMDKS0Gvd4wqreTVtyhzhzOJgy90o0iclFenoD0e8o8dsGKk9wHde0Cmxag7YIG9T/Unu8pOEtIghXPIr1LNQ8AnoVLCqAZPAL3founmldV6pQFriqwc8nPuPUDG2K09v2+X0BS/P0b9zxtjCNp2Hy92yRPV1JyDoWDhONQcqO0+huzQl5MzjTDLwNdkjlpBUn8SbQEmS5QVn/HOYc5RpPiL0eeBPfyB2cb10uisCT8nfCQ+AcJ9XQ2F2ZvXnapbOZONTk1pLCUKTjqppNSQBRkP/3vdHzptmrX7Q+mMQcN62QTsovmgb"
`endif