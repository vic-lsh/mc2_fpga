// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZBH8xFjz/Ggt7sP93WYmJn0tjlsW7kuvbwBxAAn3SkVO9FBjUXV75GcrDgVP
xiZuWZkS8jQPj+RGl2TpwDT3ome/Vn1lfPjtuuE9iMMFlrICMJCbUlr5oP/5
8WQXUSuaAWBdmWXjP8+x1iLjhdFUWFZdPaGxKefhtkDDUIfaLMLot8LoW50f
gjG8/3iL0ae0gNbIciTZiMzzudF6pGXRiJUYK7xz4NAVWSYqexBKGtyMbLvH
dvV3dYOHzOwYq04wIJ7vAtfOUB1tjpT+8g5ixeY8fiXAfTEjQaipLQdMA0ih
7etgCSAd0fEUewHjgnb6DiACmFdJHa+2xdXoyxCOxg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KZFuEdH+biTDwB0Qm8Pj6qQKAvVB7Z2j4KwmdWA9FJgJacySI9WQnT75uov/
eytdr1iEzeQD94R6tSWueb/ZQ5xSvvLCX9OtAaIAe8LqSzRh7oeic+vNsOBx
+QJKkWWuKSAZDR+DccwODmGNjEsjsYPYRoq5DQ5kr/VwpxmblZSc+V1EMsUI
ngRTr667iqD2YWRRBW8Swx6Z7Xe4gj5n2rt0Ivok2lO0lYFYKLiPz3oGC9/+
qkdSvWpcUF7Xq2rq/+6rbeVQXNopks2Plz9zM196tfpFz6oiBInmA+4myivX
GwxLXzEayXNf7+2h0IkX0xMEgLZHOJS0NUYVYQ/mRw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mNkkbnjGBqt6eL2kC3ZmvXSh/HVTdWIb4I/Sncz4+BM3FpNcBzcolaxGbEAT
PWXgFe43VUp+wlNkmJLeOlLpBivIQIXp3frwHUGBQ5+aSlAz6LPw8NMWf4th
bq3wiHkokP7mo1LLKSVUxSG2899HaNEdS4UTVMXUWvR6El+ASj/mFsqbPB/J
+1xuVPMWglhu/rWJbKhut6jMeKM08h8kv7sOsmderK1GCiKI2QXQrLlHvs85
AjqA2uRWml/bvkNozwZnxjHyJR45BdDNZDvWYV5F9vFkAKKVnjsw08DSe6tv
0QjCKsBUzR/E/49aaRyysZGQlpoSBNUPHvU/KaI2ww==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
V+9SpKh1xPBdNTTX8ckOlWfpkNc8pjQv47EdbVm8e2D21RBhY/YbTrTDjOT2
/Vvj0died80TAiErJebyJFQI4YEt1dKHXDuPNBwAVKt2SXXhRlHZ07bxWZa6
93wql9UOCqyHJibxfUzA1Z7tXDn0HDFufkOagKYkg7mqBpUUJPB+ApB2cWXj
gKjiK0Z60t2sxSpc9c34ZxwMHd/BxsrCy3uImBT2TpRS1KTsTTlhA3MtY77c
fGBx0gxYJndC8NOBGWVVi0pdrviFFuv/uFOqExE6SsKSv45ONW4RdRC0rglO
I8m524Fz+umZ/F7QnwEgZ9LlKLVkjnFsjQv45n3UwQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LMAsWskA0KEfLq1gUTqc7Y8KTkzZKtYPyApdOfPhrZ7YtjF58/4NlaB+U6i0
pPvWdi/XOR3nsyzNpG8JnpPzl7Z9TUCMRDC0r9Rc4lFX720YeP3ElmxKoyWS
NC+OPe8rb7iZ+Yvv55WBZekROi+LXIOY5zuhbQlZCE5cdNKHqMk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
PetFxQU95H43wfpxT301irFeJToJYTQACdZxfOzglqpn/LtHW0UVpwgc16aC
7N4K0IUUPv17Tq9w5Qd1+sf+sNxLj+I2LGTEUGajiU4Sria+bANqcLnQnzYF
luYzuWa2CB22l7ru1r+Dx5W6o2mCj2EBtyIHI2tq8doIP6kWL0iF4fhai3fW
xoOM/DefVCErU+aNBdkXSqPlZaPkXKhHaMdWUsLhBHGbIEoNQQ2LIgB/F2dB
s+o/GDCmXlZ4vhUEAtVPaUf32MFDIu+jL1MZKxNMvbxtqvZyRCFpm8cTHNsj
RCC5WQ3F6KUEzf/Yb6GpF21MnmKVNP+0y4+78f398nU62wJXBMtq8U0BLiAG
Hsz0xSmRJy6QLvzD3XDl8r+MKhEqebf+pAHMxPAt3H9Gi4NzlGiULygnOtz/
vFQRAQcM4OqjrwOdotxUox1epkCv4Ej0fPzxkPH4JcdnGi9N12U3vp9HycB6
PL3xj5gYCakexSxegnWrBc5KNRxd/QXg


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YoqXONBULWts67vVCniz2hqGKj+lW/HXpFTErm3DFadR1It4wD9tMmlbu1UA
2f//KSdVzWMvSAHiTm9Gm4QO3RAHMp5tZVGFfJTaPzYEr3cahIObR+l9oeil
86uHHNjYfU3YMuox5txcpW6RZzU1Y05J4vYr80fekVhT9CW4UZs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Hw3WOIaVcptGKHUHpQ33rSUUZGCq2bZlPxlI+mtO/D5m2SCYwNVLNQNNXZjW
Jz+R8vEs+3o6qmFpNdsXyPT/4ccedHeqaloQub+scZoSSaMFTaBYDIaiTmhQ
pYHHL5IEwvyCr0t+lfTLdmSLPtylhcDamLqCZWPSrQBdVugZB5s=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 992)
`pragma protect data_block
UJJCJXKi68UZ+tfJ1aWSn1Qp9GRpOGJG5841QgUa+H87EAXNflgXqDC+R2LC
yWg1qh3WMDVvKGNmwRi2cTlqy4Hzd1bM61fi7KhkSYiNl3x4DEMahEcOODuL
4J/ZWDI/uGKV7OKWsWUSREQFhiPebEkE1svJmCbJa2Gv4YYYC9Z8qaaxlKUN
4S22Quw9u5md4dzNrWFO2FwepwhEkhowb3ZS3og+qPDpolv5jBI15YSblE1J
dVmcy8LUaqZUvZzY/4gFWOVIuCDIOvT8/fzDPTbNfpS0Dwp6zixyfghCWQaZ
x0FU0VRgtexm91RnBeNJMEdlnfXkXcQJmnLt+QpMbH96GQ5u1rc/+hvcIQvn
7qxMYtYMorqaFpknQ+yK1S0tsAepcrHUQOfzg240x7qZGJQtrG0bzJYq6FPh
Dz74jRoVH8V1+yZXXF7DQANjNY3ZeyowhVnijypfa50OVnDFuGlXWpS4Rdrd
3py8vqEpbKYvqcQTvCpoDxZNs1oBf96XJG/+9958sbkW0XlUBAMZdpHaO9ya
MCmYpT8R2nllJSNhpTTk+q+YV0rjJA+PQBbqmv/adMiy+MAEm30U7u6+WG2Q
2FBI9jEdFQsqmgKzBWxCfucQ91pVuGS7QNW9DRmj+Ls4wEa1J9Chku5HUUn9
cKGxmKX8eKGmYnoKlt0Km7eHMidLpvInuCocwfxB+pGfzsPBTEJGr/Z5oodh
/Sm6J9cE+g0Sot0IXrs69KyD7v0zno0OGu6K311MmpD9AIEgX5UjozsENpa5
KK8uy1qXuvplf+uCVpUQbOVU8jtIMmlK2Xs/MfuNJSuhtChAn3EQnbXTzvlT
klXw8fhGPGdDkDur4UNf6PY6Wv5NUCFL63ozpgUsGL33GwoYxZA7Eg53FGff
Ki0qw9PQdx80OQSmYefOKWCBD840r6g8dEZh4H4IVxBDE1iEPkyZ++TV1JaN
58MAYN2353EcTzZpWDimT6N8MgURJE/URR0oD5XIYpYirbtKVOCiViHR0cy5
IF2DIFI2WRiQxLWt//jCj6UqLMcbvbdh7275PV8BCvVRCXoxAupdKxCp+NFP
5yi18hJaBVrYlMorS5ivEKuNG5DYyP4N3N1jA1AoM0iwx+344JZ+iBL5EVe5
ZcW/MSY4TII9X1L7uvaUwAqKBYy9BL0R/Pa/vgIgpfaC3jZMc7FJbCXUZ1aa
Sy8/USyNhLR7QxefNmpaykoDx2zjSC7WMfI4z/S43qOt7R9t4Bvu2V02Cqbr
UMcD3sy5EIL4l2KqO2P9kljK/E8UwtDoVIKKkzRbWnIf59BcB5IBnf0C8s0c
wi8=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fidd1oyAhusLLJ6+7Y4fW+UxvqV+8TisWbzB76p8J7jCbedVkgTXiBKrUzNVBIRDckfBwS/gk4qyrpXnk44TsazVN20DO3TdF1x8MmH2pGcTjxrJqgYV/z3UJLaYPiY1WrKUNRPOAuHkyYvfI5GoAsKohhmpB04sGLV6+cGIymx/RXK+eIUgAROf9S5AOXsk1U/Lqv4gR7i2yfj3c/IhJWMX+Ld3X1LJ1lp+Ly9OQoy2VNv/Z5op99N/Suv50pOwoTjgkXEH4s6iRQzW9r7UAh2f0Yq6ExicyZgqQOnFgGmEB9eMdj82ummDa3Rsy9qe0IWTrXkr+bXUhISsD9C4Kpo0qTbdIiGr1y1pV0AyjOopvgXvpyKr4+ylB0ZaonwMwPj1qYL2wA7pSLBBwARvYZWrESaPeHaQbDAwWTfiPvmSv6WuTD0WxCM86GkyEHUziBN+oPzF66gn0YZFfxLe9de47T3xTWWMDBa8U9L0REkkfKhHQK39DBxnqfwRrcAsnrHf0jMRnATxGM24DnLeNSg+czjPyK3QM2a3wl6lhjxCcoT3/YFIGWyvh6i1ZYrktxQXYJp0BWCfCuLxD9rF7IfuRhg/G8YshWhXgwj2Mg68jwERURXCO8N6o7I3JYhrIzTcias5cAjDLoDHsdGlUgvqt4vWs47KUQFnU9o79sgZPBJDClTrse/IWYUqym2J8hzB6KMgzYYRenaz5mRJgqTMQ6/bng+cU4Ts3FV3SLyU8VSA1rHMc16/y2VCj2/QA51ZCwKR5260nwVz4aAPNessQR43fJWOQ571cFThe/uyxlYh2cWvLi4H0aMnR731tzAAhEtmoEGTOZ9wwABtGf2pFdlnd7rtsuVYgHau2AGh8+tb0uO23hSkdMqwnIlynhebOG0pswP5Jo5kz6NXq7uy8ejl1J+X79mpIFpmQEODzpZFmi5IPFKHQVaaulEOsJfy64o9Jgo/tDd0VbmYuRODErusNavZwdEgzIXiZgi6JbLUQrpadFsTy4STx37M"
`endif