// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oR3/FKkz22Ubf6LfgrILCV7Miygf3PQpbKgjA3KW13dD9W/EIQ1c4ZApF3Mo
WfMiwgODxPM5nhGBPT8Y9YE48q7UMzTmumycYGSvX5ihhNjxlRDDfXf9bxxr
fVIWkZ7cIDxtPL5kE3FIdbfTl2jrn1Q85JdcbBycfzhph/Whed/uqUWqqrdg
pnl+8rZniLJVFNQEsPVAmgnraHqhk6ThlxUNIyD+STdQzlGvb0RePq6zI4px
HYZfhbq6/g/TJx2km0QJhGoxzu+U9THffHZfRp3CiSh1nwyEzdfsjJID2XIi
t6slR6Y9he8sEKtch9wXpf0scsTXvMViCeyhRTs6lw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pP9WooVdwXr8Ho/nkkfIzqis9g40o632LoDZXeyiAMke0mTVp/S49f/cXOjC
E/IovMn7MfaXd7OR4SKk8iRkIjpsB3RYkzAb45WA/hiuTVF2jN13+JT14bX/
BO1kqUT24/et9m3x7CJVJJTFvNo4L/J0h804O3QiTHHHvk9FVmYprhmVikZ0
lcbL0PjbnduOIpKTqlPpb1NhEgDfmBpkiUTu2JRePcAVBtRFSTFhjdkk/Huq
5+gUuCH41CoSntDEBT9Gtw5i+gdgCLmdXC+emweMvDLJjkYL9sKekpXwdX76
D3qq3aY2iGYC1Fb/2LpLwSlGc+vkec5MI6KhffiFXw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Yjoiaz1XWkKvExCJeKkQO6QJ+UNPCGRdV9Z0/1kwQlE5fp/zcwZkIb16JE2E
fBmXj1EFD9vhEuGXHGGBbZUGDRWJyAP/jJkNGiPCe1H8Ztxr+5je6HS9nmpb
+g+s+YWJFimzVYcMuzTR7CJYKxNY8BZPMiECDt8mhAnX/Zc/i1e8fHuTx3R2
BHbAykxKOCNnwZqTigN0hSO39vo6FAgVKNRRwNJsd2PrDKEDL5OKlv/lFcO2
wqNhec1NgAP8KGOz6dLMRJsoMW3hxhhHtTAb6sozJzUQdyE1SjqkhHaxY0CA
1QSN6hKx2DDdyvCXa+KnMPHoncNee2/acQjEtC8QrQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VVsjRX0Sz0X/u+5gboO3DiwsWLv6WeP54EILgU0GyFCd7BTn56enI5vYIrxj
+F5d4qAyUHmcKMUYKSZWZXCA5JF7N16A/r6o2r81/W22EZEynbpzm8d3R1PQ
CZdQTBGB8RKpgm+LnwuUzch5+uYxK4puCRhtK1Q+zh5gjeQ/TdqRnL9Ex6X9
uHV0bY59Y68GDFSPIUhgirabiZShZkErPqJ1I1kM36TtKR7MygnP4yBfszXY
VAlWM8z5XvTyDTueV3zRNNbW7atmEbb7RbtiEuYV+xGhXgYWhur/+dRR9xmC
RkYmjtKHafH0FTs+NLLAqicEIWLCBzlk8QOUhyNxAw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
r4oLxa4M4VcLhyxNEia0E+cYPEeVk/Ge9m8qXVKIe8XM8hpe87UZXYphiTa0
+CnjqInBto9HcwEA3Yusa3uE+/dlhnmjpBbpGJ5eaViKrQ+F8efyemK4l/QY
MdUlVYHjS7LchO7Dbeajjc9J/Ixu//SgwuUgKiXvQdp2b6e6Ts0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
yWnja2F4lJIeO4kLBy5EhzV70Gn9H6GARU2w1UrB0I45MTQDERyzhUuAT5ht
6oM5TNGHWlbOZsHMNHBM8GOYSJ9+ig8FuLNN7CBEHCLm6kKYsF978o/pKTJ3
Qs4fF/8+OGQmrTy119Xbg5NOO1tfb+/lLdVhk40XgEN1XMq6Edf/CeD3et5L
AgnzMxoNLEJYHSVXGBboLKm0z+kmmNmbrW6CApMVeljs6SVi/5mVyxG+aqtG
7OVZthz8mMWj1Tog1o64hKN3s9UrCRHdgM3n7AGUF4gsHDME/YZ/+SWPhjvs
cEWMQSC6eM+ZZnXBcEsSaUJQda1DVTP1aSCIzfwk3e55F6SPSDypmHTeeHJS
uiT2ToqFXgmxt9JLMFHSjXtLHM/iuhh4BymNqUB9lKYtUZY+zJVnrqit57FH
3nFa3xXSJBhB0ZfOWZ6IdrEs3dQlQy/Z6Ltvw1FlUdpwSBPF3DZjpCGMFwQz
UV13ngIcL9YS8wP5RnGKr+d3d4TYumT2


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
q63gidOU7N5t99rH9o8EJLGdUZhf7Bi4j7BdGT/Z7IPG0hX44LdNn1QNlzPv
0H5Z9pmrmUqK5+XjR7NQuT6SYj0deED3JSxbds5PdjSBjcItIObVkkt6CDUp
PeHwEoLleV6tlTU7PQWUbmXp46Xa9JWZ2fXCg0gF7kx2lMEnAsM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UTx7aWIWTlNwNE7ciQTNkBicwTECgfb55Adz2UE/iJLFc3YGhRIQzO+yuAMT
3cspzkR19wzDdXQpw9zVqi8x+Ab2JuDdPYnnjRG9gJbtq5g93luVnSpBqFzz
m3XtWMCelMZ7rpy5JuLZ2fywNizA1JkdqyzxRaSQRnOogNcHZds=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 150352)
`pragma protect data_block
JeyW3QWfAV0xI47BeLhNhEUKIfEGsNWQ7oedo9JdcwwvRwOzSWa+MXhdG3kI
cl9UUQztqQH3VpgSZxYuG15Qpc2aVYXSYUfOmq0m2oxTGh7oD8n/V+U+GHzB
l/GFXl6OYWHSI9cSLtlrUy0E+HrIj1h+THr2s2TKpmK50L4+U1r9wtHu7odw
QLS/t8umn+kpbDyrFWtHXva0L3Q1GD2U1NAIiqFeb3A6YihQOK+XpT/4moAn
MNpMOaqGywpnlXQ6oOSVQtijWHYgLCDkNz1Xx6GdneSYzb26qRaQEcqwUDb4
m9FRpCMR4Bu5oX53GrSwWXjxQbbDeKItFSGaWDFGjQKzlSdENq9XOF84xOw9
CXiRGSlcQYzmI+d9fh9ACENjXYUGU36LsK9RGPELKvBdLhQjSBMdBG+PC8c1
V3mWF63pjSaZzW9UXmbdTCsP+w1HqCYDayYAzPdHHqVd/9mwmAYsys0WYFlJ
RHF3h/Ga0fb1+FU33tQ+ToZ06rYoFDwfEz71EAGjBOzRLc/0sHFnMO1CsYRL
E18ViMn0CQyVKeOHFwdiAkhGUVBfJdmpt1CCqDcu9ecn9R+nTTPw6zpma1UZ
ERbNxDXhIQEfo2blXrasc4lu9QH8f4F7QNdV91dy/YINzWLIn3sGZ566XFtB
S4Pdt8BI4RbZREuNlj3XKegQ5lSVA6hGI/VoyshbZBSHZt9hMk4vECPGQKy6
EEWmPPren0zHgczywGWKJJbXn+jF6rf9MJI+isE7w2aUBFigvOnOWcXNl87C
jbI++chfZ1OsprWr0nIJXxnuneGvfup+21aMs3vx4EP16obm4pjxQxnCAsE+
zOUK4tL9oC1FSDanYieGMNm1B18RfIWBVKGNvJemblwNM9HkpG3qAG6b7FgO
aFv7InkK2coPkbYpialM0xaPgiKyoVDs2xKzMxOi5FJ7Vu8GRlyexKkMrfED
h+0XEtsVNZTy8nKtDZCusT+WdhAFlpLomWV0WmJvq9Nu8iXF1BSgVqzbFTO0
w/NASvBWdvoh+4DQSK0AQunF+GCA+iFqksHSIljvFONBYSsDkUv9RtZRTVVy
KP6seKYZMKdfP5jawbbGV9A2WI78XKf9EhALAORswF27N1uABbeQLIjWU+Mt
fxwmioFkd1iIo13h4FX5PfplpJ+ZGjk/fdGvfDP71uObmY+5rKyhf/MGkpfN
o64Z+2WdK0Sqsc+iaSQ1F+OVBJmoK55tts7Qn6jaO87Cxvwtpvt5iAo8EyZI
8+48FIy0cQO/BKihHqBLVx1w8nxVtnNszoj0tf4s00Ldxq3PB625kanDl+nw
hIaj3tUITcjq4ehr9PvsNdERpvOEzrDfrmUcfqWEoImsIQuPAfD/mVmcowlc
LonXfPEIl01inh4vU9oWiR7YfU19kbWCi7mjLMzh6bCzektYCHGk0FJ3ZsJ4
i1kM2+BZKrVBiCzdJfnetXVV9difZjW/qxQs9w0kCjUfK8r5EP91sLZBKcWN
KZcbd3ZkX5DWmtAQdGdNVmZu1d4PXxsmDxWbHwoH63YP2oxWHrLVnA67gs5r
zY+mbmQ/GElZb1wE4rdz2Wer4/1NAoIv4RChFN8agFRP7WU8CEJX/OiUYG5c
/VsvsvSNMAlE09mWefndO384aW1mghTVGSFGZgjwOe9TvSeftENhgLHUUWo6
Job1kVvs6hke5sQHUF9kn9bXimp8h0iuw2+MTwbox95LOnFtNlnohfx9K5O5
iPXk8hN5B6d4mpwJIUz31GBJvRTiQiFCcrubT7utJ1EtNziOLovICyxOGx+R
rYTVnL6RBVtCUznfFNy7Lsx7hSbZ+FtGOe5H3ISMfRomo/qWhMzKATN5JtyP
jPjLkadizjexgIxKmLHx2QDJuQV25A1RxuyNitK7lDmxAo7y636gLFAXmTt3
Vl0XwcaMgHWpA5FJWlq2xZnqjyJRZhO7ODvii4nOKl/bb2JHzbW9UBt9B7pz
57CW/1+nKMkBq9chKod0WuNXsRLsEW+E5zTaKKCZ7fN5crrop0W9+ZRyFqmM
IccA2i5j4zrhBX80A8b5jOCuQwWosaVRwrAyo1a1l04m0eUfj9XDD4j9nAAU
EljhrH3OoN2HwORffvZx6lODBnDj+JGZXS8TkNQCwD/p8BGS82mVFCR3hWbT
TKbjrJShgHmNHDODhYOV+Z4zkOOKZeZXgUlQnUUTgl1DT86TFgiDsGbDK5zg
gJU9HpHcaqEJfpsqOLgkIFMPNIa7v4wVnj+aBCDMdxFD/tVXUktJS5VlIR8Y
FxYEvWLheCX4Kc2kYXrEojJwiqVSI+KE4Ag0ESXAgcYeB3KVFcSXA2y1Vy+L
CeaovKdIHo2YVZZHOEFggBmfm+a77SByc8u/ihaAHuSBlgYyXWxxiU6qOntG
c/oRNgPZ/7bpTgb2pmSgdafS7ydJwTykMNzVZSGFctp5EnmRXUTNECxkbKh5
Qa3s2rgdxWlQucAbNOerst9LdCvvqXXUuwtmhQDEv6TVTCTYlBhOfQN2iG+Z
gguIvEpjf4q8MmmC3F+ouLmlHJGNj6l6RNUD4SmojwtFB7QG4A96w5DlAbeK
qvfWIoDjvOxH/j6PSzy3A+rouWIipV7WEJS1WSmpGIolgik6Lw/q3RwDzQV+
FFQDO7MX8bfhVVSfTLGGyVA6YKqxy46SpM++iaJUzlmeqpyIInO/N9n8O/W8
/21QA4YmxfTPHQ+FPDoGsmXjBhu4wDQrHqermJGvAZ23M083/3hFFEIe1kho
2eR2p04ClUHEBig6QZCwzWY67hVlGNz+DYOiIsmP0z55AsgetDBaBcR4Fj1r
czD6z82q/vB+Mhlv5rnJYkFfqbmAW8OsV4TyUysq/qjHnRVkMOr3DvBhDC+I
ICVUGPC0dnlNi2CHsHpiwPg9DL4oUapH3gSKWTNCwcW/A4Jy+v7cYvaeEqDr
PwlN8AVxtkMnBDAK6/UVRnVfCcra9Myxr/0bXwMAlSWSZZasMaWmV7owGaXD
JdDL1FTJ7daEtsAnlZaMretImZXqFWEIZiHQnDYlVMcJE3kZJNUh3PDyCEm9
bFpiHIayuQLvkmqzt8vq2H3MQE6ZRmp3LR7tI5HH5rTKcNLpQTIBgsXD3rpf
15imqPJYOaFCEjEFCf4aoJ34roUAg7tzIfJVtNedwwADNuPB4IcrlvwOmHmZ
nAcdG3opGJn8SsbY2KdL+cmQhlPxm+JWDxh0FuY8AfjHArtxt2VlmmXuK0ms
1TcdP4p3J9FygFnnjakQ0OgMd7e241v2b+TAUFFNw26WQ/jCkUCnIB/83DLq
SDoWry3pZ6UmWQ8Ei66/QcHtNHY8vpMHa49sViuUHh2iZTGCM4tIh2Xln65E
vcSqKJqvzhz+wuBq0e5q/BVFrZ7GtIyLaiCv8dmoEK9JDKjNGUs7b6HWU30v
HLKjY7adNfIFVZXOjHpo3dKSZxq+KnJgXXcZbC3uXj4VuIIRB0fOXyTB5A2E
PNqieeuOwX7gNyohoqjP5iOw+Zo4eAYm2dlS2xI9m2ABlbLbz7Krkd8cJHjT
Z2/uam2a4PT75FiOiOXeOkzKnEXXirqRzslFbd8DQSMYMPvxcEL5moTVNzyB
mF3LbYc/ol+6okPEhCruaenMSG87U2k6xtMRsmN9AAWv2L2LZvfj5qPSmoGl
giVt9rv2hlXPiTc2DuSpvBAw7qUS0XswM+4tlkTlUiqbYlc9BR269SAYxA+V
SvfkHFuwrwA40snVG+YZVUGNscZXAENvLBxyU/u2qfw9bt1U+GUeg8028Hap
qHM2h7VYdcv4jKXiak5+Rsn6OXVCJeOlAo/gwLM4LXobu6yhXJxYnWu4K/BH
dYGhnHR6fZdqa1Uoiopdfpn6z0XImKZTilSPmHYAjZyO/VT0CBK26GzfTSL9
ayeNA4jdHVkledBKPdonrBxD4DhIby0x2D9B/7ELJhasjOKls+hfNXWmSpiM
vmB96EmOhFgXw+CmVyCIXxsA4Xm0pYhUdOn6HPrrDLteV1KiKg2QQ7kPEqLI
6W9IaJ1Wx5/YANgkq919sRJp9x42cBloN0SFVNEpwLViKaxL60nC6KCXU5rm
ktWQQA2LS1Zy/dJ1HUKz3svkyQJ/FP3C2j2efWNzqupxFyd6h7ZuhIF6jKWM
sWlZoGvtCZLW0Jm1sSaD3BmMIPAw5zKFCOzDW9hUW7qQqgJjtTT5dxXuv65A
4ICsHJfHBYiIHZgwkjuiHq8wFh4ATh4Sr1Xf+G8s6BkPl88pGGNS3a5P1PYp
6rRcUUDeYhl6GHZp75x5Bc8qFDtujzdy6QIZINN/bDK++vNWBQwWpMBH0cab
FyLgvfAsa4m8nzG90PRpB5qwxxqNYDuKRIZAl4UTNyW2xfBC4J1qTCbxoLxn
g9AKrldSOxEyiscYenawoPmE5gZb8dmJNqjYLUye/1L3WcYq2XlGf0rCpT8D
E+6Cv4cU1XFiNWwWABZq9xV4W4rob+6Ozer0TtqnwhmMHKAqFguzMGa6WFPx
lzK8Em7mgZFGPAihWU8jFFdwVvN/a53DJ2s5HLow1sLgvYbFHKjbJVOi1uUb
r0hYEGgQxaeNtTmhmE1zqXcio+sgQgXj7gL3UjCLwMbDDeb247BQUw7t+lHY
RHCA967BXEe9L/CodBdxP6DGGKOQlI5/QD1sS1Dvt5kmeaDhO0mNKewlXTy6
ShmQFdk0ByypdyxjzH3Pw8o47xSxDHb4+CuLe+yodqSBcJW+lrZYsDEyg0fe
IrRadv8tETjetp4LGASl0phyt/2RIQ/xsxRkcuOIgF7jvrBvQueMcDUxFqR/
uL+6EsjZ+HNwuYGefFDIAAt0oQXqYM1dnUqDHKHRVZVN2v/e4RjuNRUxkhhr
z7ypow3T1xDmjwwMxCyxtFH1EkXeJClEI5B4RExFN5VFvXiL8yFtOQzoFPEK
c6PV/QxSC6D80TiUz6xbyNDX5PalyafJql4wEtFqLAbokHnwXO8Hg7k+I8ar
glTDhMf1rSkL0nWEFLJgh5JOuzBZVHlnuNvVWoqVqnnZACg1D2yPbLD7jndx
XObRu6kwpq2aU3hZC0SfY5OoGv6kY7utTj+Eue+pbYaql86Xp35Vh1M469IS
oUOzCdFyq0q4AIgsYm9lOY55mAysperlolYla0tpmUVNy6AzN+SyG7EnpiTV
HwXt/YhmuDq0jb09Q8saiEvM29i6IWs+VteCQzTqGdP2IvMPzUtNJ86IP/uP
tCfBa6oa9VfPxfhcts0bYztB9qUijMa27Zw6PeP70KuvjisZpjKXAq6B/UMm
5tKLU+N/2Dr9MHI+g5fncKM6VLoBUJFvzknJWKOweuF46hx+e7akVoLyPkK1
SWzwtOce3WOQHOATkcMB6tfW7FNvPfAnEQe6gYRTF22d9tiCt8IJaYiALsJC
zaUnP0TNox6Fc6P6T+RyQNQxVE9fsWz0sIWV/z//TLdrK2KTFD1IKRHolP+s
I6UdzYWx85T2MOTCz7Hne5GRMLgIUpHcLIL5OdlsqQo1dQErIT7nfIcabSdr
CIMfzPt1TQ7ccAIMP1jCRW/b/riLouco3SiaYkll7szCBq2H2y8LyiZvfOvP
frwjS0N/NDOe/RD7iLEPvH9bTikKsIFaFHgwR/L5CuSmtIztEIoeKrBZL4QK
cO/I/+AyUOpKLx8u9SYAffcRy/Xpgo9LjJAkMuyFHsOoIhbHJTVPXSBS5bK6
rramE3gSiOPUUz6Sv3ePw6YG24oGcu9SBwdE46tNs83jF1sWsQfCWaBesSby
/3oXJA2s+NCovhDNA9XZeHyGZbVMwlGRuh1pqhjs9pvAYKHvVO/0xI+svjmi
cYvvlNF5He+LTssy+hSpKD+0wms8xI4958DKRqdXbdT/+N920XXeO7jGyp1g
VoOJmnWH/C0jIX7CbGIm7iax9RyD+319Et2XV+IHSTkL3/qx76/lbKZVRhqu
yKnj3Fev1dkpzwpydtsqHxGzPThLQDmWK/KInZ3O9eOPnsmM6lCoUx9ax69g
2ejYDMuc/bSTbKcEPfeoipQt+tzKWDWS0UPpQ+1J03HPGWMLwD9UQ8Sn91Kk
IR7h+Rofnp90N7fwnUDC+Kp3fPgMp/KRkgTHkDkynU22ZDKx5PwkkeBIU3JF
ZvOb3+wbGGFXOXeyg9eeO51Sny/9WeCDIR/Cxw1WqvdJPAz9ywYVLz//KoQS
qAtPlVR3ESyF5ovIlNBPHNXqg5eNrYcEDwp8WOGDEPXSNugoVxlL2G4hg98G
esccwE/m8Sjc9mH2vbYQ2grr5ElHfP7Omjt3ccOw3ZELVk1D5kXPWPzdfykc
2RRA2IEofaqTjZVPc1tw+WFKxIzMOn/b4NjSeU0H+FQoS7fHssDe9sK4zUlD
FFkMy+se5DhFqZMMx2LlslyfyB0U0AXcQ/dwD5KKBlv+62Ug3YhEGcdU9KWn
KTDVuWbWXlC1sJSg5hnFrnFXA6UHb59DyT645fmF6MlTBZXgufJW+3UwKYsD
8WgFAN1IrUAhH/6ni9v/z1I5KCIDVirTaQp3f7Qq3TzzTAFKhQVkIhYt7bY5
E+hPDIy1ByGg3LZYi+ybFajUYKOcwfUNpYTQPzDVF6f5MH/5tcFF8ASCFrQE
eDr5NOGsrzhGi5CZxT3NssW5xhN9NT6qLTtf1l20hh76bLHTORlJ3DJ56lRJ
JREqaZUenhuUH7nEMO2fjGpbboCYGpzI0e3YrX7StnEfT1R2iMgE/wr4bDeS
NCRUvovFoGHZvkMsYtk33x5UShO+b8KtOJ9dTZj7Xo3cPF5JJUoHfZ6Ktodc
lBgIVKBFIPEuDz1pkKVN8wQb6XO4BAK1ndCEhx2ga70HRYXaOeUXLYEvuT8H
yoDKHUBn/5ctw8pMOFHSWEinkR+hmWj1+VkuYNcUSkUdPqSWWcRpK1GBYXv1
d78fiuUBRctKPaBtbjbA+v1CQrx4UATVVlVLWf9HR5vcM0lZwN+16egkyHXn
O7nfhL+cNAOaBYffnWWpA8lC1kv69pLHjUu22yYskLAh4NNJRzq1gdFGtXoX
C05mUdnX72a9mbcWoon+0nrOd2YWGdRKiubY+aKuMSPgFLUZm8RqgeyXa8fV
MbMkPch+5Ot+HXxVjKFLIT1uS3rAzIlNNc1x03SNuneBE17u4dWP1ZVj5W+1
WDggtADuqSXq/chJmuDaAZenMWC2Pnqtlse5O+g+8OU2uRWM4+KtSGv8GZQ7
g3vN4jYe2DsrWluolQdFvRNaFDYLN37nuMyxoyDZcixWm40JAqhm99SF1KSZ
1uOleXA2Iz4EIg8zBJoRmSkkk96H3XfH0Hs+Xa2IxubYEsUS2iuG4IxDC+Q8
9jk1PhH4LjMm9FaAlnBkXRTg1Sb2d2qn7R84xgmLubrPI2ENaXRpWbo+NZV1
rlnAvDyjSwB+v8bivwWlfnrjuH67L37v/UhlxIUDJN4H4Mj5qEHNlwmQVJnP
9KcR36ebVRdpo0X9jqBsy4Fo2vvS0Zzq5va9PMIzVHmt0yTIPwChTZ7ZgbGk
NVC28mTFz+dkZr+R1wlHiZh+fOUgvZQR5GAxdPPvXzMee6absab9TkeTcQ1h
l7lnZKO1LO0MNbyHUIpPpCNXNablCq8LUVt2z51doMbVOU7TjURfzmuLa6cQ
QJm/K7O5xscEyN8X64D6eQlzgnUoHeh/IA/fOaLN9RqO9xB33lQ8H6FQP96o
zV2VeiCNZ2RJS6lQMV3E7iFBfoM4z2v02CNlBxvxNx3x+Tbb8a+tN/ZQPp76
kb52Cw8kgnXnpkR+FOa0CTvo0W23Fna7c8ozGyMncRjc9bfqZsjL0GoE/5Y1
8BL8ZXB0LCLmNvqH3nISLKNc2Ba6ZnSTBpMChfIAe0xON7v61WtGMDgaUFpw
mBCmM6uCvKoeu2bqrYeVEzAeyN1GelermfF9Zl7jBfRCqUaGHVC9pmbk8FSP
slJKVLoUg8ZNouN/fimZpIOulPK+WTDAqz+cuKHvHNghfZPMuWWXkWsJ5nRC
3pmkZUDfHu+QzywlxPYthkwGjjiYIgD238RSBX9WzdrO/wVKBPuRyx6l02H3
VCSMQVR6GcFXUIcq6VzNlGK81yql9VRQPABy14RkejKlPdLIo8OTpAdpoDzE
L47FP8bmVcNyWZf3yGYhyI+pKHJuG3/SD+dbbwg4lZy8y9IwLcX03/1QU6Gk
C8RCODFF/+8LjT0CWdyh951L43yh27+V0qLY/iZQuom0NRQhORkoYaFFvc0K
1WZ98hB5e+ZacGNouMIh6SkxDU0E9jCjXwkmpRw8PnWDvc8xWFwls3JKC50G
cqJn0HT2G424AiNXJEqQkGGxPXfXhP7KPAe05CNfwYxs9BhUolK0WpOXPLh4
AcArICkDd7fsuVpHnAb0DVzhkqaIzZh10ABSYUdsAuEx8UbViEag0b6Bpo17
1yV8sk8MohK4YkkadSWqfUvT9p6BK76KzpUY5wqERuewLydPx5mY/jqJIVY9
VRiH2FC/Rx8WWdAXSu7hAr/QZm5iv6dGTSRsxN6rrWJOhCf+DKG/aW88nOGb
fLMAGgNmB/tmNUnSzL21wTuDZCOg3oPtsZQj1RZEdno8lWcioorDDUO3gJu9
6D9K/OO8R00Gu2ZGlRh2pJW4bgo+g48LDg4nkop1iahx1Cg68n8o1F3nyOsd
LUZbeUVmSC/fo6RlyDQEk3rJhRUMZ8wKv8OLmrb8dZkBUXvUzQidUtOnaGvE
0BqP+BfMIPYDcnHhjISawNfafy91/IvaL/ppyFdkJ2+t3L7I9zLuResu9Hca
iEWMXFMWGwROL5xS9sU9qNiQhcrr9QpwJmHmKS+VST84daARFNgukV+DALkU
3FX1wjaIDuG2z4rc1ClYxU6ubUHAlWvqpMNUP+YGey/QfK+T4hZnNNxlyiKR
uiTABnkIGMKjU24PI5Ao0lfbL0vLlrVbtuqj9Bn6sLIUiG/murI+1D0A6oUW
8BBoSP53jv1mAlgNgWZQSgiwY7szW8McmA8flGOyaC3D82GPP7Y6nsk6CsZZ
NVIr8qqK71uHz4CAYEIlBHWwN6KUZL2b3lDlxRjOkFUUAzmvfVQGHaGrJzGl
Glbcn2Y4y74iXfqeuwWZH1hrDVSowIQJq4TnAoCnlJSX7PlMHjnW9loJp7g7
xcas1glKUDjttBg91ZiN74ATzAgu+XNNLgv072xKjrR3ajP4TiyFUpNwX26u
Aysw+XZtWuYSQF2p55NfbWxev/Bt3nECvazdxCXv/fUuB9ECSBZ/0YngIuKP
hh0UKVbF/Cfr8cOpy0cjbAkeRszZBUDykHY4Sp8XaiQcJpmRd0q/fA0WRkgo
A7TqhDXXWCT/Qj7zFd/Qjyrv/YRmqQoS1sKzLsFPY8UdKkubLbxe7op6ViQh
JbyckFlmkA2Cl4ylB5IbBhmP1FwHtvboQz/5mRFdl4hfaxkXLghOtweeF39M
rb73QXVDhGUlrha6ZXDME7QdFZ3MdNiTG38rZ81Ujdy9jqkueUmBbGEyqzDm
L3gAiK0Nypd1x3L1jD6pCKKtzUeETUjfPD6WhwqYILINTpAdqTHole/QDvnH
zn2nuZXfrHHAnzhGkpyA4iy1pcB1OsXR/y5dSoKSpg5Yi0NPfUlcN3E4NvSo
EHXksYkGkuLDD4cvCoLHL18SwHitwtgJor5dDb9g187vacN1k2156U5bYAcT
eRqR8DX89Mz3swkFZ5J5fsA07CeEKDANsAMBwkKi5mLbB4gUZ8aQc5wcxvLI
vz9jt52D3I2S9pZoP2WdDGRGrx1z0rHXoEVUbMETzInp+QQJvoNndF0CiNjV
5sk/GOgESTiD0Z8UmuBST2V03WN6AfcDJoEuJd9nurefWI/ssQJqt4FbB5A6
2hKMyPTeY9nKievAQlFUQzHOiqx11HnAicWASHbTMY6eszFdLYqabKyB3Xb5
b09DaqxfCfX0mB8Cslko9Q1d49iWJsMwmdgZV2yShdNFphBXgTzw+cxiM5aY
gE91y7kBxTAhgnn762jn/pyR6v5X6WYpXUQ6wtfxLfs2ZqnZYE751yByrVU3
5rsZBV2NCJJJWCz/fi778O2AvHeqQ9ivGNO/matTU8RcP2decNI2sAHSYZhr
U6xiXKdlj/mKOmNv5dZZJhwRHUQZKu3Pz4mQoFxoZLUcV6CDAjsBDGq5ZXfg
aTRufGp2RMl27xXz93pVLxOUaabMZpDTtKt2VQQGR37gYWZyPbnBLXmjeUmf
ZFS6aXWFkHrYas8QNRg3v1r9O6xPSXh71pBAVuzsAOuTtAAC2rwXfjf0HLJd
g8lAqdr5na7DsyrBVNXnL6m3Rdi+v2N6msNc9U04U/0wkDBnt4eD0oAge1/A
zTNOoW3iE+Vw6cD5E7aqWifdzZfJoaPiRRm593bOil+t238bQjx334dbsnTA
5lHPrrGvBEDhyVa6CHce1rglne6X7rp8nuLgBSZmtAwZ8LpO+RA3Ry/F2pcY
Uhdrg2HsudCMNgo9WSzXdB6aGbr8Yt5v0Satc6Dc00BBuPiRvw6y55uPLyA+
lltF6Cq7A46AFWDCL0qILtggFV+8+Qwwpo3fUjkhFrFgWQOKfxilEruyyP6Q
7fdq83Q15JZ78uXgdZlcuAsAPNrIGw/D56dHfu8yMtXbkdKo0DRpywVA2tOS
Xo1/87B0OsrvcST8MkBsNah7LWCxqG7u1ZqOhMCiGiYp8vgG01KxeaiChNxA
FvOkndmLh7tojZWl/I9ihOyyn026AkTDa5/Xg214W8Q33bmr67/ugl/A31WY
ycfOUSh6jLBUOxnZ3wxBWF8i+sAOkN6R6LM15Ypq26DnOSfdw1PO3A8NsIHk
tetB7xg8rfds5gTPM6KEXpGve6Q9pOeQKkkOvBHCrtwvujgllo0gp4/Itc36
/g5mIlaGZd8vDVc3NMPh3J6Ha8UmAWOGZWo5k7RUotPUQVOvvAuChmq/1PDF
Sk13057dXCsS6f1YLdBVagxcFidWRDcWHbucJT4fihcUHzrOydQwVWPSVSnv
5muRI6fDRdINohqvs6mEDNuWFKQONl2g+mBPXRxDMIHdloVOsDEMXZ7rsD8j
Tc4+TPi7YA/93nrA5eoJA9MBBi88h2wkRVSJJfYg346AO8+aBtEkJuKSFpsQ
a4TJOxVt3r/sF6zcNhU3YgRc3nIpdtaZR/UGTQETVCh/AtaYihMSV8Iq5X1e
CNIroweLoHeBmEMgAdavmSUaaQ7WfNJAsAodWGDyxEs90S5LS1WsPsqZgntx
gHLUJY/H/KMq2cX0Tq3h5kt7bPdv0Lf0+TYQpxcX8dUEgzJ6ZaTHoVKTD3mv
BBtxWPGRdMM38tv0QKaRVY0MQOltwR6ZODeKJK8H+con+g/NL3EEB3DVGuge
bTkaCBtI+TqB6vehDSmCd+JurhZhyFvGLFC6hK5XWUOmeKuPacLcpqANIAGt
XHdvcUEE1oDrJacBl6kwet2BL4q+KN3lbhuZreHrdskSZc44s2DoX1J5qtnT
iDFczVyysWBmLSJ/fr13qw79HO1ZNVQl8bCw8kRYileFVBIbCsYvDuFjVOIB
JChPY8uP6IHYJG8dktqIAjD+cYk4DYaZBNSDwjAMY6Tb5qDrzd6quYA3CTg6
T2zKfy2sTiIuk4b2zbV3FbS/vKm7wPZTToO3vEcAKtfYLhY69hSkettjGUOj
oOE8f1lPmUSkwicFPl39DYQ3OoSEilic02uTijy8V67isED4srIJaTZRdk8x
74VsCvwUsdQNpE/Ci+8/+dEzJ8+/+NCyKIJrsrvn50foPWMPCAElz1UDnujZ
D08xttKvDetfVOvDVuSHGwVsSZoaOUMUFva3Kh5zGSHcxqPeyhAJq4iLaHsp
Nx/7X2mLQfSbLF8Cws/S8wM30FG/bC8kt0ijC18mkKoW+KVCiwr128X3KAOh
7cIngs0HJar6ttzTNiOBnc6eHdU2KjUIUxdQuZobDLKoAvJlrLxZqPagvJNG
BvXNUp+griUpGh4uBviJPqbx1FYBiK5447BC+shxKCn010rqkCjgjFiOnrth
dcm6npBJ/IGjYPf7pcT/AhDCZKVE1sp5n/ZpjOeJG8IBu6R93hnX3BdrBiNE
GRChH7psq9mva8vSRK4cStim087BDYS4jJU256ujTLJyMiKaV3xyLCmzBMXs
T0o5EAPcL8bnF8NhdicbE+r37eFTXTmYxnQk6pyREocVXNgACFQ4ZvZoND8v
JXHHlLrY3PCT27cC7AhDigDo0F9STYorQ2bMMjYlH3AtpxBSe0Nav3m2EEaa
beWxZjjKBNp3UHU3vPsobkmTdEDCsbH1LL6eOEaI//xEPo6gxsERy5gG8esX
KGXFgKq69QpjSqpvnpfiwC6CUxsN5K82IUt9yW+UDBmFybvQ2JH7k7f7MWYd
HIfmFfvhjpCT7aE9NgBRbXp5T8V08lKNwF/f9SjPvyI59P/AfmShaLc7fTp3
KhOJVXdfkTK1IGWSxnYFd3C79muaLRwaZiH7P8T8yjI+kBloF5BlT36BRsu4
uvlQANStL5nqCwEGbED+F8iw5IL+/nexiucvJ/kAHjLXc6JIr1sE6yGdeg6q
EJrSb2VQ6Wp7gAbU0NjyrWxIQxVIFxhIoORB6umuBx1Tz+D4LZSIDnOG4NXo
m4oK8+Z8O3VGvX+l4+8rmG1XxOqB4q7+M1UyY9w+uh8bfeJNqjAo9K+79q1q
ZnLwVjVrbbXM4HaKgekmEvcb9X0iNrPPMMFEuDTFy0dGflL7GR4zrp+mu0OH
y3KoSVe7l2iVE1AAQsSVRBDi/N9GC2IhNSd9YLGey+akOkJqlHy8qEH1vj7C
wpkwqOUZEU1P8XF24JJG1mUIuNrQcJKcDfstV9AtgkLCDa9DFWRZPYCJuiYw
QDg8eJZtExqoci/8jRZwMgYo+o5+yxgKazre85DgC6h+w7E4FOV94F2v00rt
uxhac9BuMt59L64fRXCvOXkPiaArWqqPjs9mfN+slmX118cHYmxTZgVBXlBD
G56Tavi8/votAAs6H3zsBIqEUMGxVB2jk2CiO5CabOK97mWtEK28mq+ywHtc
y5O0xUxdYFt84vqgs91TaFw48/Hc5co08Hshn0vSFyqn2yqCfL6KTxieYcqR
j3SOzQYh2iyzCVOp3kz6Qt5o9p/9o70pePQDLgEilCbt/uzzWBUoDmtXYi7R
Myibus0H5hFKhkelbkHLvWuAjquVjCrqDpkMwMJCUH2uaeBKjHnHyZQ9espW
4sWSIkjIhR/iEUtRdpB8r0KJ1KK/3wD6RKwta+/utADLrD5Y97vq2RmU+fbU
4K1Go4aggj/LtWcwc+0YrUat7pN479tXZa9frjwDxPuoEG2O/TFIUDnCUHpL
HfR0559Gv0ep3AIHb8covQ0if9bh9Ibyhm+GPQXYUCTFQYrjLSZDCCisaGha
C05MEs90dJ/G/NTTGjpT9NeMEy4AnakT34uAIDClzzuXx9jIPMJVk4y8HAyP
saEn00G7GWShFuHBEJsGfNfz6nOvGd6GR9HhxRkYRD/e3CDbBOtziHH4YFeG
KfCYbcOwPGFJpdCQ9Yztn/dZEHRiY43S8nlgI19DAwAIU4Rapog8vEWYjGpD
sX8ASS9ICLFu6sKJS/SOZYUKYW2uf0diyueAuzOYfoB/vK6gm1AtnSR3Tgcx
Ce6t7Z1KiP6wZ4GgYKETOPvpdMLdd9ImLkJVHYHx4qI/9RTgXhKtj6PIJOfM
4NmUrirBWoi5zACRjXjJ2SYnDHJn+HZRmf23TqQ2eNH7BecLl2DTzElbGDcO
kQ08mbFjilqxd2rgoi9MrDRYEh7+6/FfsAHo5yQGoJGGrIjhTKTif2D+UQWl
qUElADGVelLbHcTBQLQ40niuPNY7XZstAan+SsLsx8wWTQpVApWqYvV94fAc
pqKKVVfoDOUwDfXBavK7rPVz3/n1yU6H56KQ03jPnkXNZrJr4GaxIDYBUvkU
aMF5hIOzBv6etYfIadE+KMUJU4N/fMRmhvhxrafkSc67tH75kR/P/iYZHQpQ
EQn9Fr2i6BO40cGt6NWH/I5w4eOAaRHcPi5EmFMo2z7vOf0IPYSJxcjeBobD
vWIsvN3EEoQHEh06mfzFYr3wR39HDqoLIFX4EfEAwlHv1Hl+H41ppU+5IHZh
VlmlbpPrAw9wvtLZoZRDj1VONVJIw0xATn/iRsuSdHjN4TiYHNvPgZvKxS1B
Q8qMYr1xyYNYe6ASGftzF1xuV4wSSuWySg2q2G2qmrNiIkbvnxBTWmEwTRPe
u/iZTR/nKJrszxQTvgFy7OI9MHsSKsKWb4Ks8Dhd6I4G38odGz64jG8JDCKi
Q0p9aTTUrESRMVh9xfmPcroZ0WD+807JuwkMYAYepc0hpT1emsIqYqt88+ra
MZ0ZQ3nnsregAV6oadNMAOs7qgS/OvalfUiAs6efKHIj4aNUgbuIxeoV8Z1N
j/SpmEB21Gfwhi29ajMOsYlEsskSHcNvENaHlNcNYJdtJff8x+0rsNTvPdSY
9arP7GKJ1hUAmWIjLCYNNZ1zDQkW0+m5REsEwq7lNN0NZ7TQo7cJYRIu8g5l
jYPyBgyG4DBzwR4MjDpEhWXK9y4XFHeWlno5GAcypBdZUn6psYZZvAA0aemT
QRo3MDZNwQUqxW7nVae4VIdg1F81ftXVJ6eAxWEQyFrRcfxjuiRT4k/Rpqzb
92c1tFakm2B0R9qdO9cVh+OHAsWgabBgQ+q/r2V+jJCxZ13T1QUMTEiekgug
oRpFG+g1Rs+gwy96cX8+DByVsKtZuqr+d05u30UVQHfrDu9D7Xnq5zK6AkjS
XmMyoVMY6KuHJHb3zy6xVO7ZsJqH3PbTslsnOv6O25gS8+cR66r59buiKfU6
WLlvErJj5UAVZC9fyORpQMKhzyTK9IOSEhZTPkh5QqY4rG/kgd35fec9Gbpn
5ebuyY8+rY5fZJnUsJ5wOemMCY2y92xeJIUqv34ZaE/3RWPqMPs6MHWAHEJM
BdfC8otrmY+V26z78x2bpUkv80MN93MshTRf2RrS4ak0T3/fW3MVluFuNRwn
3AfS2R5QBS5Bb94fBzAYkDboIs11wtwxRPaj7Yf3gZVUHsVE6MaKn09VkZsK
I1L/qq/dbixvYgFCgr5RjIIfoixB3JAAizzQ8k/P8BCZ5l9qAF8NxllAb6cR
YUY8/HE5yfRMYp/XyaOu1aFx0tLleNYrJQxjVEOnnfjgCo1h7nRhk+AT1XE+
EfSD+5zkfXgLh5AlTo91yDXztxqIjIfxvQrWUSolXySCdQMWz41UHf3srJ+0
KuGBKCqUJSEF4OClURSWiOTh5H8Yb6PNnjGNh0yFYo1FfOd7oQWgNYsNR+px
HwdI4PjepZ1izFmCxN8S1YFYdjmKgG08KcRzZJaDqZHb5NIFKBKQaaWyioAG
E/c6Po99JLpl4KlcSHRj91Myp9jE9o1Maa2USK9Kr0A2jp8F39lOJNhb+ivQ
S3HgLm+a38GtZr1l0brEjaf7hFF1oaZ3I/5K4p7rI5+NSlO4mMKjjvQxMy+B
vDYVgtUq2ri/Du6niZvM7M3QxpdttGznS0KTlyHytolNJF+prXAAzIGfXJNy
5K2xTTZK9Z+zTFVY/yT8M+VzIwopEcHMcpxFj2FXx3Yt5z/jGn1AdAnJVhU3
RKAJAvOwj/smjZVtd5IIc0JmfYPEZUx3T0NqHeAGStLxsGZEvGPrwsUFPXWV
6HCw/GwxdJHGxWKjmnEmyeUq69WpDWK/L2826DOFTfecW+Ey2Pq1QVxZ+J8Y
W8C82k4n4Rx4Xer2Ex0mQ+oJ0PqF3bIsVWJBFObODAqbVdDCBWyxN5EFzwub
rOLj3jfNYPJlrpC8yn1kAEIF12MwHBGuT+B3Cq1x+WrPDBz+vb5Ov3UvWt8R
N8a1RXRpkQ1JB+a5SKDvs2C6VTikd/vZw9x5rK66RZdz9+mq72g1NOJqm2B6
oCGgSaqBs4s725leV9EgvPCz8Ndr2BN6UIrAoZtusTD3m7mt9GXJhnUE/WnR
IMTOU954eNDLvj+dIiUpTaRo15F9d5oCgzDHLavashJ/jkUbf2aP9wxa6m9P
Hd9k5tnFTx/U3hoRMYbd3MERAjl3n0Tm4yLnaceT5f02hZuvVYf4M/ig28ba
FD8QtxJsNsIpfli5A2v1IjyD1wCsK+6fSm1zimPiXISBwoV+9zFp+r/2BDe7
fdPEms9Zj7mV5egC+ZdJmmIRLuSln/GuydBw6P71OFV6p/aiGxUa2+XZ+RrZ
crDLLHCDsfKGMu4i5yPXGcDC04QvldRgLncDpk1+l1Fh55NgagRchqazFvUQ
bM6JwTbtuKUgEhMbdLYbOC9xZSqMSy3R3GVAn+1pzun03jWmobCm9TxlS/FN
jeHz2d3t3UmbZLerCYnbbQ9LqSFJTzfzwdXrPojSFAAzslcPlayVXEc3cY1t
/w1zVJeB1bm3E6CygMHQol/moAXv/NdjE+yhKXSUl29wk/njOs+chINTf+wO
Y56SO3JXNxAP0XYoUYwXZ3bBQjuDoMu7O/uiLotOQAGBemDPIu377Fm2WENt
f6djYCb6c+BmkmV6B9EtIbTIWhcQv8agR1hPJi+RbfG8QXPNhqDUFBeQktGR
FXZKlCFUABl1qqTpmu+tp2zwlLdJ7yC91pB/kjK4V44Zl4ql2YUF6VKj4Yla
MsVM6kl81Nynu4cusvcVYHZYVll1okSE99bJMETfADS4vxGQkxYjDkLDQw2z
28NbtekwsMSnB6ya+7a42XooEqpctkCN4e668n/Zw2mV0gWPbSfagCDdZVWt
wNcVvVz1kizT/5pOJI3apU0LgNmPM40+cASHwebA9kjc9ViV3DzwDzstchMw
6Zwh7BVOVTWkvjYfuFTY5GTVgBCINnWpDyBHBJxtoZK8JNCFAG3Iw50vkVDA
SGBNhxdnZVaZKUcDK3AujVhbsJvnjmus5ffw+ex/nLBfHr2iwfpY5OfPryDP
8vI7b7P42YsmkJdbahCTGEJTdpauEJgsvT4vlechX2tQszjp8OvOqc8kzM4I
okUm8r0/n5IPU3k+eiyNjLL0NvvyptZ7o6Dg5kd3ZWjB8XZvMAj1kvm+wP3a
U19+rO/fg4WodGa07xvyjDqINxqWk6us8eeLJUJitFqGzvqI4aBTET3xnQf5
T2zOC54ERPrTHEIFN70iyDQq3HHuQ6sliUceo7bduU9vG2GhhhU7J053HqnC
UsnCQ6Zbz0TCnc/MmaqgOOdcPMVPIiqYEL1kFY6gM6pW/nG17s7QqJOi4keG
hRbh/sa94np/JV7yynDA8Bj/lew2yrnDJUY8nKce64rE7JbzS8FdHAR4jcZA
HxyvanqltmGqFrkWRW8hye0NVsEbTlV14GUElZ+7dtMGCRKqAKQ3VUrbqjoC
BS4e5FqE3y0vfrV52VCEJXoGDuV6gtJYYTZ8bqHXs/VKqr2YUIYomZj8DpI2
U6AHmjQ0FSLEISnGtlc8KQHe5TTTp7Vq06OazGS9z9JFG5oHzvelRm4oAX0Z
OcxuDJ7LTYghfxYQpIMIOr6VfJmA5pEgiwA3mNZalZT1TmVDZ60sLfeXXHjC
1faJHe9eTUqFarCZ712I1ZBaSXtIpqNdnNmJX/smuGliTWHo4Uj8LOsHLdrj
UU/mni8dve6gabhf1oYKsFMrbg0mhx1NDusUZ+1NNY55MWulmOCwk9fFQwYc
aXp9DvCdsCqnzegUDCwvedHQHSncZVj6bPpvn8nfdlKvYisqpYDFdbH1CmaC
YnBO/c1p8oogsstupQeChGGNGy582jl0BeQoReDTwYlOFethzdCIuMtv+bd7
CH6g50QvulA9YcOlFawKNqCqnBUxu2PW1viYPyVyWuRjhGWOnUL+f0Fda8r3
0tj27vclWtXExs46gKlWcFWsSzjtj0DG1/Zf5APfabzd6cdnfZKwV2MBLLXG
1lIIKo8HEdjN2Txh9LsrYsRBLkyI1r6tIuz8WSETsgTEoCdN8g3Xt7nsrt/6
pH4dU3eUP/zx3VAos7XJOckfnOP28wZxYJXf9TI4Suf0RRi2rFq3BReAHd50
4FlquJtENdSf523rhgX7FrBT1HqfWsNFvayon9oETWjALvSTa8CYy2SDlzn0
qBIpVlwPRVzZSbq3VPSvYV+6Sd9QT1xJ3YoKr1G+63BRr+w8ASEgaasznCcR
qVCwXgexmkrPryqkQyTj/DbGCDyxhXerAqi/cInqPNLK+G7cFGOX+ohzAVOQ
UwbpN919wPfeoFbBCfcqam2ui2VhCZO5D6vfWTjPqPxZFU/oZzm5VhyVAr7d
I6zKcFvnXIA+LLdV8tskA6jQPeS32YKAAbeOQgiiaPoZ3Kex6aAmQvLcMgV5
Tc2YvePumOZaPNZ+h+bdlyCCMyADGlHPcse951WsA+VLdfIsa3UQ3C8PZyhJ
4NtR2lqB2sz9eW0a9+QrWopqoUPi6zZhoNKZqTfRGS5/fUO7tvjiV0Q3JkD9
8Qp6IKTpI8kr/x9LVEycanYgT8OXzoYs2ApiMYP+xRS1f07X/oaVU9c0fLu4
S0lf8roMXoXI3FvZN3C55ZvZqgQFPCjUvDqt/2r1j+kq7azFdGDHhaM+eRDk
kUSYQWZXau9S87PUG1S6qZUifiLUHYbxw64vErLOkNPIFPkL+DhSyj3jG/3M
eLbZMyqCJ+ET8tgaTvunHp58NY75D7s5oAk1hfAFc2NbFh+B9hjoBBTa9DS/
1oRzvHGfn8yH3rKVvlYUSxq0yuv4DkQsKyMrLQzpiGu6VgQLqHyEg8ulnbI8
i2Kum6EVhp9whRp43B1AoPWxfnc6xmffDoNNXB0DAoC8wU4NZzlQvSivshPX
Shy73IU275V1lj1LOiCeptS9RmrLjOUfIRYGA0Eln/gwuhgCGlejOVyurnB3
L+n+bMDooFcr12AiaPTsCwfqRV/kouImKBZVgO8uuJtV2//W+JaDgPhUYAcl
bQYJPdzNT66R/eZsK8V3zNSyKUoT5A5shwyr6wzcKWXtTGmglWmEXk6aTAy5
xumaBykfxyqtO0XNP5ExfK96mc/XnSApjTTfBUIWw+N1+/UVbhWHGgdj+KPQ
8ovHvKX7L202XjVuNm/xowPRwJ5NZinkZO1YoGSbEGe2twmqWsGcuZ3yBiLz
//ywhLTd+edmR14cXU+rduK9xqz+brFHrZH0oEH2Cb8j0aptmvAd1F029S02
5W/TwvcF7dk3t+FjgdaCZKG1E53Ly9kcjMjYq0s0GW8fBXDACMqq1s1Y7j/2
9Q2xXt3XC9lnyhvAJNDNWyE5EuW/0Pos9450VIpoaPEdZYoWWR3xLBW8l61q
zm6Oa+Vb34z1xN5CiSDRlAgTgpLLBZCf2YFsvV7G9cEMoSIyRvgx2n1fo5wj
kbgLurMk0KGuraZDa04nki/PVR++oLpEUW2H4zcYcZ5LbvQ5G/USX3RM/6W7
J5BQ8+s8GJglP8OAMWw9iHT2AeUTC2D8Y80NqG+OOQ7xtrKadBOWOW7Uykar
+2XFbVGOSeVY5ye3uVrgOcRm/e5gwqa7ytAl4PH8F5BXjUio4Bpf6vgYdXLd
mWPoJP9vpw3BXv7V9XOAKYjn1UAbMEAMc684yM3USIvwLnaITRl8mIGVADlf
vvUmhSYyht29d7ZkNsN2VvW65BR6TTuYa0CWqVdIAjcELlsikrimSizZVVbY
FX4wjzydL0Fmxfo8fdhGT+Wl3nvDYudePo+5nFgjJRtZVxSnB2DWrFqA1NHZ
6fMj93xn4XPTAfPKO9bzOV8XwSF5cFttf4JUzFyJUcGcd//70aY71KDKgzMC
lOw9ABwjY3d11RB6RbryGNT7wEht50O6dU20nvoZb36tu6GPs9OINcFeELSr
Q9mw0v63O3PWYhSgZgka6fGUcR6PC7YG5NmQkcFbE5Z8ai0Gra6aZ60ljZ1j
tWwatuiphgvdlZpzUahXyq59mlYH3eg0ENPuMxkd3goTFxu85nIJgD/rPb3h
UeR9vedzKJx8bJr9wbXG4VE1wjxyX9/bgxCCl+tem9SbC12AVFzYyJ+UIXTG
yl7DrHp05RVoyvTell79x8rmdjkY7DmetP9SwlFkwvH8Pz5Zx0RuinfmgyEw
X2pD6mKxniXQJmH3dJ6NnxAAeiL4MKa8jfMOqQ+RIOz0Hb/dWgmsvUFw+Bha
XkK7c63oYfsH0+yIBSPlCh4zpYQGo4v7k5Dy1x/hMGxb2yfTQNJMIseCYiCK
lnfSWNfUxn7yO859dQYN/Z7Zr7nkwTT0qQ4mlFHH7pEaxt3dfrl1sLbxms1A
tiUNXM+EKWtCi6WDrbmnpMjZsmwhTkRVvzMwBbYWuONoviSE1evcotMAHdOt
T7Y+jH/QxhavYaoOI5ZBOI3f0wCpibB9wLm5L/c+bXYoLOzT1j/67j+KFrz+
RqJ1Hi3Y30rWO6ComUdCulqZWESA5HK/MtqqGqjbNYnyR4rPO5O9cwm1jjri
iplN0ZQufgiiGzic6MvocAWJyKEM2RoVHN6AoCUPTmY2bvt1cocQEEEqcTvf
0PGMaDDK0YPkC56BCjG7GTB0nkiyrnSDp/s6xyiRow8NWOpgxNTJ6brA3nj8
hgD7r74UPpLiOarzU9gn/bojOKqYav+gIotot0MDFnxh20+O+tO2dKpNhKqy
7S/RmIgKebwmkRReJa0lb2PhQlFHY6kz2mFs9pATE3nBRuyGsOH36Xtbtjvz
/rezDSsWC7GTHLXmJ5QA+HgM2lY3gugLvlG6TrK2Rz0o/W9FTl8+T6Yuupyv
5jGuu09Qp2UgQsh7fS2ZKgd1wxNdQwnxB7yvIT9U3jJ0dbm3Q54/3GE/ojrj
7PTmX8bs3ipu7iZc8+o2BdSAx8TgpKob7aIwGW9CHacQ4fteDVwndAR1EYCU
CroBLzd1/WSyrCFab9cZgKQg0xtPyydtvugIcYTb9fGiDmc02LNfNh5KTDJm
jgOQw6CBPZBlYiWZ0s6w8XRpwZNyaGsJKnL3AqJIpTxYOd89MCvjYdVi7UIu
Y/v1zj6fpsuxEgpvQ/TurYjKKPmy++EqRbwbaEUoJTiBKe8C9P6TK8jIEjHN
EpXHJTDgE3NGCQ7iGyOoYoB+xQUR2yB8KE6EY69HNDiWSJ1joR0KmZE+h1Ux
zUbhSDfTJ1kCWRw7kQKBrjS4GDw4pe8wp5M30vUmmDIrDBI/SsqJYbXtX0fE
8l+ob+s3UBTOJT257rnStF2pfeTQHG1kY5dYNUZ7YbHV9Po0hgE6tvmW4299
nAxX+jYvxuzIiyTsvSPYjAvShV7mFQOMGRJlbArs3xJ3E4+qclTbtaz32Si+
sytT0MohWTl/gmAZE14Uydm8uDo0P5+GB6OS+pybOnNmaPGwnFTxO4Wf4PWD
8UjqHwFPH10Qn+yHWKwivvX42FZb75DMrxJdLQs+veU373KEXyc4zGu1192v
pbCHPiQret+1a3I0HX9hQOvebM1dqW2E6ehUET0qsVeGeRJib8jHfR9Lt3VU
ob5auM9qt0MqbW+r/54wEPRmys+yoBe8T/WrAsmsDFg4fx3OnZOGV6qq/8LV
kLbj0rxLUv+kaPZneM0Id9VWwhNzNLMRRxtxWceoO555mwNxXHfCN/3o50PD
1GphZ11a/pKHQIwsYQjxb+eC+euwctLCh8jPMjVP/VkZmqsm+wzcraStAFCs
+IXtgSN9mwF4CAx4zKc6++25z07hL/2G9u7DKDYyaiJEMYajh0uJxp17c9sq
LXl9kSzfzqGm2FWESWP//2RyXiX3xt9tKZeRAaRetL5ekyrGIwMlC8KvrvFu
B0AIbr+yJfj40x/binKUatH0xE6qHEbQF9mJ08+I2cnwteLY0tedP/5rMop4
0FOvywvGsKSDvjtiUCnb9gRSYnnCIcNRl1aJAgfCXdjmG4XzjODq7ukWBe+p
UJ/SLv+olQDQYpRwUqVAYrQIm738NCz0RXRLHCImXNHhdVpLdX8JKhkZYRsd
74X2HnHa5Mu/Qs37B8REReGnA1notfcGuBkDgGXWcgVLfTk1/ArSg9KAH4dx
iWdMY/lcrgsgwK0ywmxPgPTBv0wkqHGqJQBvrUwFET/Rv6gjia8zBwMGrjde
2USfmIaVb49UWqtn2ubo8jv605MNiEz4zxUITyTn1Rfhar9WSACRyCXXxlOk
7hwg2UGyBwkfwW6v52KsT4D2ZiKy/+CWUop3cr0Fm5uwvRAmNRomj6suwuXY
uueaoR38gzHMEF+dHpYdwqOPU4uY0Q7oO4W3K/gKtvJ0cReIkwIRNl1nYUGL
7hlHjF19cjiXS56wmzybMY9Dy2mEMdbPDQX6bfTFplW1ISGHjBKL1uKrqoPa
RfCOFe+YGpqDdjYsbDBbP1yyfIugr1hFxYxxCrEQfGdOlmuKO5On0cm+R/9V
PLU5XBadb11lmOSXUCHy7/kNkY40iNFcBno+6qwCeYG4Vq4ifoss2l6B5gWM
hX2RkfUDF5wCxjZQpeCWzQ5hyh9U8Rd3iRcg4gvSJ77kShx++vBQHJOeIv0d
VCJ0gzvNILRA4fgrnF6lM7hKTTTrONlT4AVY8RxGsuRLqqeZU8y0puIZbMUe
5Pmgcv+J6XEBq7lXcUr85apwz0mn5GROSDfIrIWHy6pUqmKMESb9xtCdZPIj
zYHLuzclYGP3EDSFK3ltE0F7aIEAHSG1ZFvsU57sEV0t90aqftePrq0YMJKd
rgIgMP3bWgQUPYA6Mkw1v47+cZ3mBZ6YbPKgNm0pD1dIQ9XOlkJPYtLD0SuF
IJpqzoxcYeq5Nl/tw/fhnTGXY0NvXNz+YQxZiGhaghDxgJeM5vMGKR2WywOW
v43ZVFTvvJgrnLv7f1xq5qN6O4cYByBNs28oNFcGoqPYKUb1XrzYl06x1OF5
f9PWAKGcBbHdVQYDIP/Zs3z2MA4nq6cYoaalfweDKhYGV1Q2VaN2Fepc0xvL
H0HJnTEiBd3Kt/0PR95vw9ahGPEyps3lakjx9jObrznoefd0OS963ao7tnku
73URDPgEq9YtQJn3eBu2OAMWBeLXCmDy4qxdrpDmd18RP2tMLwSOYXc5Kp+W
PFY7VvtEWWRUatUmlZXLEgVOEW+FrL4byyNtWp1cMC1DEiu8RSiqMdhg93u6
mRiz4l2oDANGwKCvxcH0IxDoW5JgMjHEo7c4Id9WdI0OwkJ1yrOuQNDww5IU
nW9LPcVZ6/1B+oaHJQZvJJb2O0JGVqTLgvCTTB5S9JsWmG+Q6+dk0h6raan/
32X3iZKkstuQfEIdc6UHEvywkzbTKVoUVUuix9yhC976uiUgIjzmP6p40y2Q
9xCRfHC6m9walChgUpbFpwL/aopC0EuzAPQ4qVkSIRfWLSM0bHIEvLAhV0QZ
eJsikx8AfzT5WRTUWor1N9Y01uat+R4Mt1a/Yl1tzfQKSon1lk9Pe2ASflFc
6l0DxOml1BJ+ZRrXdDKNaYULcagoy8DoCJjTcz+TQy4TrW5+f24/EfqPXuNj
iuFU5oFyr/GAgwDtsSipSC+25+uvcZn/o5vLVnCNCaBohU7Yz1aoiqXE+J/h
DbRjFhOZyNXMFXqhj9kGGR+rEQ8J8ra4feSFDh5OuZ0H4u0RFHiEmMtuDP8K
z7chLWceZaGVuGwdwv7g+PRBZyQpfnrGEVwWacFLm2QuI1JPyOvpi21afdEW
llTMqNynH4HwxjYVnbbKWfVr5Ij/47j+k7T0eiN+lh9ZYr3/2A2uDKyuc8ux
d3AHfnPzU2UGUMQKK/v3p/np97GXnOpiY82BX42zTWUCsDLwn/m5tcrQQtbG
5ij9eJalyN8bbLDfPucWXii+FsxoIJicFncT1yrYU4anIx+a5uFdjxDje2xZ
A8MtvAwZzpyts1+MJPceyNH9022n2C9PL63kLPH04lMq7hkuuviaGhafpXN+
24hpCwp5h5UjKgyUGAZbD2K8Ba9lvKkXtDtveLFMR2jYLmSMIcqirTZxsTT/
Z69ZJPfPjKx23+6C1pAWvp9xsRsjb89SkOGpQS2VIZFym4BrKNgDAxdlltgH
d5LDlDYRZE1b4B4UqpRRDZyjYSV0U5xFIB0AJO1jprBIZda+hcZgDC+5gQ+y
lqwWrbSsbLVOz4km0hSmo3vpKK9od5j6hDNYVVQT+ren2u34dx1sDK5w98nb
RSv35WKoodT2L02qdQsjieOtEbaxq1WXc5/WsBtEojUA/oi9yjocXUm7cVb8
X8kPOMfSe1xfYm+dI8hFrHi7ZhfU9Ku23WMjzgNOg6wkDLJcP7JKbNi/cWRP
7l2+rormZLPDdmjwM0bxCxRTBED5Qz6KPdhyvN6odHvRL5EDF4wSYTLG4AbN
VAzoAFqI0+99UpuTDYv6ry+hlx5bH132/5HpxRv96Q5mKL8R9z+ZOywrM9nS
ruI6Jfj++6F4jyrVz8Hrzq+6CldnJc8y8ogFKeVSyF39KrPQjHlOkk/K/RVC
OkvIjWFev6Zw78eciAYFPwor6/j8Qc5iTN2V63eT3g6mPa99V0Xtfu4LpVo9
gTS4ZxChP7XGfJYc8ERaXNQ9j2uVlyge+fJJ5/bQwmadoz7QC+o7c8Qnck7u
RjC5fAF3r6mcf7MC2FZ9Au4HaEMpBPDOde4AaPXngmZwTBW7+b56th3ldNJE
NbWonWi+ZTgop4tUVQ2hWAFvIeTfVQuBCmxTzLQ+nczlUtvQIIQDMphiFiPi
WCc/y189EFnVbA6YaAQr+e5nNx3Erf59N8CrFakaMmFsZ+Q8F0y/zOl+KUbF
z7GSf66q+1ydh3Doi8XaniSH+/goXmELW+byT1Vqwf4DuxtKyvg4ANFb4grR
AQUjMGMTYoaazs3hB2sHZIMR8t6aUILuXm+JECggIRKbxQhwTYAvC/K0MxZy
0QdNvcZFTchmJ21TVi8wiTaULb31bKWDhxGWNz18u3T2j3357tw42aAfr7qS
xX++3hTXo9i5vO/sc80Djwk9LSgUTeh8O0NZl4c3OLW0TYQmSsfuLAlydyot
5njekzVwFuvCtjbFNqVixinYGzPwergjyMvFi5fvnVIagwfP4zI04JkTj0vo
FphFBVh8tGOmHs10M2EsgD3YHZ1Y6E6Gi9SdEhxgLIAL0jM2CdRKMHyNTvxr
WvSBpi3ZIDzLPE7WDpkm5AwQguLPqZl/22QGXJiC66mFFqhKM93p/sT4vjk1
AcLEJf6jmllBo72lVjzEeZDhW20Z+K3fHYFsW2wnkmFc9JJZZmvH/rE4pK9r
f11+OdrWqQh4h+WhZbB27XQUR9hP0mxiuoOXX+bfbcUou3o5RsrY7mryXPkz
l5awkm418VGfOtXgQ5OegTlymtt22mrTDme+Ne9Ylzj+vTccu4XHhtUz56RM
EiLk864WkOhioFhFsFTqoKvUpA4UXKSvRFs1+RokaKVTpNNcOCXeE42GIiiw
zr5si0cbPj27AznTf1HmngJz66ZJuc5cEvu5aG+owve8XdVFnuEATKabimap
QcXMeJFB2Fz46LCq3w8gdcQ0oi1KNgcS2LSt0Lsz8X3H1uuSH8J9XVAB3zIe
XQb72ZnV5P1bVEK6GCeagEjNcw+rnfEgPYAQsDQFku8IExd34haGJ8RqpTgQ
uMWTHF421+tcURLUmzHr7oZ73uOQxsb+edwT1buGGXNXVlTPt9nPklzCgHaf
8aOUPfAAxoefdT8d8M9bnxC7NfGlAuGTcG5e/OkRAta7n7NXkRLFxDObMRKF
1WaA88BxkCIIWnKiIK8rnyon45BIpsCdWCHpvFlQCnG/5zm2J3D0y4rr58Ya
+nkSpp+8s3A9AsySE47IH1mhqzaWtIYVIAhkoc2p6z2SkLKIyyaxKLw9JNR6
bhKYXNzkOT6Rb7uFOgE8YQ2oJPuCLJx0umTKSP1NN6556wyswvJaU6XDCXiq
b3QgmTjG8twHeuOcwcEzx9Yyhx7KqIsljoMKlIyUdb0R6HffgD0X2OtKzUKU
fqTCaAIclTOLK4721HoWGcEd2D0Efpb5qhHVVkpj41w5PmT+BnKeA1UanWrk
/yBvZ6UG8uydUIcUxLwBvfxPqR64Mj39jD7IqUiO3uQvTWtpeBko4GALeuh3
i9N3QZYXkppcu5Qf60xhQhuSkxZ2jZpMnqWbleiFtatEnuzYRFu7mfOyAcI7
WgDroaQFTz17Tk71jJAWSNMVu50gTNd1CW79UB4/IYGSiU0sTfV847DOJqNk
KtUdA5YFaTgUS3cVv3SNrjPwX6GAmVb9ICywMiT5WEwR5pKs6sV04uLq0LE6
BbQwNQ1SNnTsSd4gGxBu8QiOVGNUFLmtHwedia/0Or7t5ot05BpiY/druhsq
IESaHNcRSpBwKApSK/Ta2TwkgrS9GtUQ9UZRJy+VOpE/qlTV7wTbIvqLllYY
EAHYU8xeG704KNk6SOGF++w4Eq3ygfmIh5wHC4WkPcH3lBeGq/4NT8TSaJI0
upW4EfpHQ/YAtqM7gTwxz6sAutLvUyf9wIUU+WuUr9hWXsAGGhZ/8JDKPbmC
54IU7C04B/L3OxMGTie+VYuv7RUvgGbKWuHlaFOzcpRmNyEQznE8w/C6o0db
NhYxv6JRiqsSqfLxSoc401ZGg9bvSxtKZAShHfFTpzEa3SHCCEfnl+ZV071I
0Kuc8dBCOXDsoVlRKlCMM0OHBoGnyttCsfRSaP+hrzQoh5u3Krs0mml1YTRl
PrhD+8lXg4OMNpwVtFpBgcIngMfGK9222Cb3ArHI4aHaE0+pwXjMG76mEXP7
Kqp9PN2pTlVcBSK1kf+KzMAewdWA07XffqK6nlnyKdnnJGulWEJo4hH/iOk5
lN5O+h3/i91N6S7aqKHAjXesODY1GERKLxfweHRTzXL8LVG+d7cNaMcs9Dnr
nln6ztKHUHgh6NlzNus/LdnEvr+MyNA6pqEa9sg6sz7uZQWnWwS37psY1ACH
0eroDQu+XE+9bzQtQ0jZgRIG3E9Ni4TpE/ERda3g30pu3U3a5y4lSGYmpmeo
bYqWEP7eOAOq5WQa14BF3vz1WTvoZoqSxKnBIAjqEEnLqyVy1tYnLkId5DD+
V0x3jFyjpwtTLFrVqv58IGNCm1AvMsKU1WSQ23Vy+ClZ01u6FzAtEpO542VW
XMx/0lovbIEpZwXU2/RKRxl+Vt5wtG32NF8j6jkHyQ8harihcZjKxxyPBcBR
JhcPYucPJPXC3w2UTqyZzBcbxnTADOcgmwK4aXQNZvAbykoe6UwNwyX0hDp0
vBU2UOFkAVSfipg5oPg6ePA1LnGpjbzS1n3M+h+zQup5YtjAwwO6t0Ozamg/
pKx4ex+SW1L3CSnCy6XUjV6hkvSCHTzF6hmuR0QUjR+fIvsWcQ55yu2bHjtV
VemXIV1hHkdndjQImquCN0nrQLMb9vQCVb1mMUO+3u7J50DpAZj9GgSm6asx
0LylDTbvQZTUxnC58aQf/WXYsoSMdEUxUOpIikjvSOHD5XX/Zp4Yuq90Q5z2
HtjFhXpfPrwxfSR+vOK4fFKY4uHnCSUeeG8NNfpYZLVxJVKi6VOWCyNZF0DM
YWiiLb6iF9Hb+EgmAsrNALTaanCMXWa7/ALO3k1Irfd5g0gMKAKVXi+b6dUt
12svuaqv0/s6zCxq2QbM1OpxlII6/2Z5qlXl1IEL2JcaPlYNg+38nq0FMNjT
VCA3Lgp3hFKeQlIkcJO2SD47C/iPJlwmzfAQC0Evk0gXNAHMdJhAkALcxm9f
MLh1CrKEHyD5c2V11rcxlR2YqK5OpVD9nq+Xux4wFuUn3DoTIuxvzaoTs1tI
tXEx/ykhApWu1IjuHkRRU0ntkJ384fUBnYxnAvBOlG3Q0/RfD9hGGPevDwKs
u/9JJZU3/LZ2GzFhugvniAhc2UhkEO/zfjfhK/1s97nMsneMgYlXL71gfyOI
I7TOgMUF8neUEbeXwyo3KiqCzBHyaRNWEd2ZFYaelAQuTt7U942+Y4vVCpni
+HwoLrDN2vKix9b/iJMqu53Bpk9dxEzmhOWSKw3qX4R7t5dG8HG/yDyjrpWz
JbWrx6fJWbyKRR0J3m8IAndcXbnQVVyPBfkRktS979ydViu3nNKEDRB0GKDy
J5bTULAiOyhxKrt6Q3NZcoH5HCYxlZt5f6dZjrWKOGHcPHYYh4K+SBQgrsYe
zvYBmAiXRtVoWUz6ErMf8j7q1j45LF3MNkkSGVdL5x1H+Qt2UdMDFQzUBxKk
ClEyKn8J6nLnkhyFHl3agflFD2QV+OH5+cD4vSIirQcds1H3MkcmUe5TeWyf
TnMmQnwPmmXk3pu1jDep8QD2wHaUT23yDdeLlFyyju2hPFHbH7QQ+dnrOLSA
QdRZ8M1f0kYfawVRZbqSTStxpTuGWrBbxSUWipJYTLMz3sPhFFqRM+Dq5rYG
PrNnKwjBxYGK28ldrTZT/yvJ7HadBaWJLBUv7Sji+O5u0dchKfL/vMGEcVU5
0cnvna5fsAoXjv7MobGKl9YAEtrcDTNOS2VoyDEGOKSVu5RKSZ+LPs3CSjZ4
OMRd1N/Hbk0Gndw8BiKhCwVpdzRFvHsm+6vlStBr5qJ/Ut/eDnteie03Zl/I
76wYqADbiP3y4LvWj2HazGszPsUHUbHUxqwpShpC8DYLxhZ0r6eGrCymBNkJ
55hr1VRVUvIORs8jqMaP5jLG6dCOrOgkjJGiZKS1jtt2LE8+RPF9AXgAnLC7
hE89/3M/ZcmNS90YEC7nj+4UG2D4mK9rhBmNQrM16A0NEXbWDsqYJTOTMrJV
S+nzmUdAtH9ySNALq2EtJ8ty7J++usR+DB9K78icf1OhHa5CikGGOa+eXxio
pZT7VO0wMD95MMAQLU6IFiBHiEcBLC4wx+s+bKHPf6koICbIADvinGt8isNv
Vnjk9lskvKhqx7/OB0kBdMPwvriZdn1ZjiYNGAD4OOatWTzRsXdom16XdZnh
e3VMHXpwady+wOfrv4XcQG61eA6jHhgxg6fqkDVSO40m5YSV1WzowNjz4yIg
dNp0btc/Uurs7oYmcJ+uEemvdRk4N7PaTICN6OYe+t5BasQDDm+XfGZ5TvOD
YRBII1crTdwofXv7C949dQRK6CRTUwW9ftmOP3ROoyEF7uSgvAw+ZRkoh9yh
gBSqrHToVwAOUBbk2QZfMK2gGibpA+fOmB0DAiUWA3zSbw47S29owalAfJ4I
q8aBIkeKsjuCXfJb2cvw2FJwz9RFonu0mMx/7FcC1tkUDrI7nUIHeAlqpc9u
1OCVhPbYi5hnNWjICYVBwcLQW5qB7edtNPNuiFu0D4tG1jO4a3Pt2xzwCpTu
onB8ja2NqgRAfsXZDpGM/woqvfMTTEpcRyA7PsKIE+PKU8fwzrYQbg/l/oQ/
65VJH3cIudXYfx1N/+A3SQac7QhD1FRovnlAcPnAMTZJi6qLLBy8+5qrD+0u
7A/Zr1NNSC8JVW5QEmBOLCIdVbdrfECQxjQaaUwYiEZKLkYA61J8oIxYCRwK
iaARESnpYtyqWgzC1mY870uxk2mFBBvIYhO7oTFHyPCCA38nx9be6ZkfQQIp
EHLTHNAJbkS8H97V37kLcA0TF6kxWSswu7TvGBDLPRAzODGWTU5oZnpBO9ZC
zNVeFWz88QPSkKq8g/a8oFb8qWy6sDDpsZv2C++0mKf6UogvFliST+XNav7x
y+eGPcEMNPxwA0UIb906vzQ0l8D/4QhAbfm35RuphUZaod9xDQGEPXMDMvVj
0GMfQuaHy5G2l/yOFkyatpWyxjBNezDehrja7ONikxM5s/tywjcDFE8WcyMw
wB1M9k1Q9NRmAdunMkh8l/cu6OkpDrHDuI7Z3dBwzi50sQA9jKs0qHQMSAzH
3/Piqc+gnTV4eTBxYHjbbiX2MpR9DnKdbdEz1eU843iDM2XyD33vAvNFfTU6
BmlCfcB7IPu2WO3TYzEsnEQne8u0p//7+S/PKKOIyfVRgJ4ZcHjQXHtgMidN
hrexu7jOsa9Tc4BwIS0DHU7uZV7Lr4CZiSPujxpdnCd4YfZzAEVErc30dJSo
BhAKZs8cNIjRT32OAHiqYXJeNYjVihibYBsgqS9lIWJbh4xxe9ZahHeToMtP
tqP3D8O8BdWrQ2fArd9r6HNxfpCAVgVGnVqYOSE0I5mXqY4a4vlv9/dLLiJa
ch4qO7uFxeSq4/Sm2qaYzYKkJhpeQunjLLYl+72vUTxWl8FamJ0gjUK5sGQD
zpyYhzfCO27aXwv9JK/L7UZPA5uC4gBDyFajhD8h2EgZ3XAN62zZm8Bd1Cll
K13jntFiGuRfr1fiQww+ZMBvfofUaVDI9bS9yte/yqGnUISzv/E1A1aDceOp
iBh1UcKAMRjAagFOSHBTejx58we6KtuOtMHpYB/6LkzlTwhm4TzBJ/67ZmY0
zWaLefMJwAHDLA7dz9g2k7CTRMjf2xI/K/g50PJdgioCGHqgCDYiQBwP0Yyv
W2ldGu+UxgbWjcl6YkQ2KMzovxNd/5P6L3//C8rEL5Nf/aPIxWEYNjqJHDmm
TIxZ+RaGcWR1kfb91p0+yosgFl6yugO6VchV54nec2aLcrOnO5TwqOvu4/pg
G46KmkR2SzVvpRfKI6zthBfiO9upM5TgnLX0sbtCMS1+mhwP9ZpPMmxZV7U0
DEzXM8/30tnfac8t7FlC02dMS5EDhI53K1WeVdbVzce8RPrbFL2KdW0+kVqh
gV7+B4UaK+2ptVffjGccpgOykugebYh5HaZN7T0AD7a7mq24tgMcvMza6uox
sgGGM8k8AkPNOgRQZUgQFwgPQHhjYN+2PmVTkjSfJknA93R0s7d7+cfN7JUM
+a/1Jnt87hha7fNNnBKEzLhxWASnx3irSoBgCPh1c2LCEY6PnPdwC29rgnHQ
jBRvKbMkxLBRl2JU95NlMaTt+VxPOr6bQjR8xvfydvNMoju7sNA6NdaLZRT9
ASRGkwOP4FyNBQeRVKJSeP71kPqJ8HZr+kJoHMdIBdyvIzN6rfEZCvRiPHZI
uZ55mjQ5trLpHPTAEMHFl23NLcke970ucANZfwWgvZHlbFqKw24si2ExpBAS
6gOxjAqyJfS+AhY4auLsd6VzEGDZZC+urz88kAXplFYSusdvlyGimywHoWoF
6I4dbouMWPlTlFh7dnDxqkc0LNRGENOUP+UchbifoYeVjTLlhVDX2ZjRyoo4
X7+QRLzClw2T8O9sJ2Dx/Fxgc8ChjX3YwGVYLhl7p62Pmybi74VfM9phNDkW
pVt2DTW1f34jI4jWSPnu5IvOSQaPfHr4aGxKGW9RzfGpHPwDX0TSjW77qvjo
zVDlxv3XUTU6Qgp/krdw6Uy3oZ41U/4lhrbdM2J2K5mT1F4cdy/WFaDOB1n3
1oXpoe9T9ZvULB2iGDZcNfQqtxEfyrrVasyvk9t+Rez9tr2/ZWPFsnLMB0fW
yaA9H67WSFEh6kQvOx0Gd6OooKgUJv8wkN11GFqjbsqjSTp1wJ8jFaeJwdJw
GxXLoOCVujh9/YC9ot2GuN9CZTjaxNCow5CNfPUPiuGzL+hcQCbXVc1tPdsZ
mHlxFHoHVw/84hW5dGTOt2CNK/jtY54kVOweA1UYISqrwUh67WAeUmQ1sm5w
gs1EZES4sfF83dRQEEcev+IkJ1SJLIZ+d1egd33jwflaba49aNh7pjg9pW4j
E4mq1I6Lw3KKlZXqSgjdLFEW2OpZYsLah/+y/V1ewBRXNXGiXhgWxlJEqEpX
8IJUX5datYas/goUPAwqA9ADMfmlAmnknWS1yfkkAuasOe1k6vTOYR04iXry
y2ts1g+XsREZnFv9p4urWEUCAEk8YDPwkw2k8eKztXVz6Jh2xiQPXV7RLY8f
qoUNGwvQkcVNjan6uiaxVTnownjVsFvsmibjB53z8evcIf/SdyW6Wux89xyr
cSSjwXcmXmO5sNmYHfvsilRxh+6mHS23yznMTU18MWAD5zDFWfk7lOtqWv7A
m1HOTVppB98V+A9RTQ6okstJ+IvG3oCyWWlOEjW9CB6YlgtxbrDh1sSdeyGU
ELUUP7T8pf/VN0bCSZwZGgX/mQjbIxLuO85cY6GLvMZreuXaNqEEtdZSoU0q
SHl8Igvv6GrFbqWsmEO+ZONZxfcVjbC1NnBiiasUIEHXxnAGfzNWuni4u5HO
LjApG9Sh+arsP+OKW2S1QT+co/MQFEpjHEhOpZsLSAyYhb0DUid/mfUT8myK
KyRTN5RVkPL6aoJOhZCNk2nCgNsXSznQyoenS8+4zHNthOy06UOTVENJD/gs
CUjnlxSVzChhj1OtmGLehtEjqLDOKUF32RjriCHcO9jq08XLyzye70WPbLaB
ajlTjs5mXnN+6H6FAFTAIEwYS9T3QC3d3Eg84zUzSmHzBKQ9n0s3CBPmOEZO
KtmVEMhPzaHM2BuV2xkIqcFLgzTX2LUWPp/7d89wkB5PozLQJAdWu1T8F9G6
zgHZ4YMmtCCDN5zuFxDimVyzcFk8GIGTYN0TndOF1cv8GA2LxjP53l0qEGeS
jCW51m8wLbv9FNWq5pCU0S5fZMUim89f55qbDgdrIorKy1G//wNc1qH5VL/3
JzSYQbFceL1VAQ5sN7DhnzXtU5YY+/3k/15RcnF2Xcf0lVKs8ACJLOx+g0fO
tZ2sByDeC6RTYGgNdUCSdsPRsRm+8fBW3Kq/NGciy7N8itUzu8nsw7/QH3eC
KTRltyOegy2T0ryBi6V7iOwB4hZ4oakxIo9152kVllnsu+qJFeFZrB6vYGyE
9bgP7M80DQ12yP88oP4mx+4oQEIp0R8z7ISVfkt75vfy67zRTA01C99T7mJU
j9fRmByGIwpMbMldc+JWpDarkgixSMwdTdD7l8qv9M3jwcQ9p1z5OGK2WJx0
LvU52mqRRCc1wyCk2Yr7+mfYoUJTWrCJofs6I79MDNmPfQbZoeCZ+OCvI7zW
ZrYC9P/RR/yw5+ALrq9Vlqs3ruWZ/bKAs8v0uX8Kf+b6a9W/Y3edJNlF6xPm
iJZO73ECdz6h+cTsC6oJp2nVhEZPoVKazT5Acxfo6FNpkbKR5g4EmaKCtyIS
W63KJbwVnJa6gHfm/SEFmchLOMdztDt2nE9xWtTyICNvDZ5njcNdWLbzvPO4
+RtnGgsnUSDcSDmzjxDnKC1gfYiHbJcAalY3VTX8dc+fVSYQT76upI5vB/wQ
hwxudvpSHJbnrvoFYOL5kjk6D1aQ75NfdIBTmsSMoulruQ98uuUDOwzIS1iJ
q90IOH0RMf03YW2PL5sVtB7RH/Dbmrg/XLswNzAfMWOwJ6Xf4uD5Ld6gaX2X
yg6Xb9i+AwMwKxmzJIrTF3aMmHyAoon681RWGN0m9vQW/REnbNDSoSoVgpcp
SFzeiBw1BqJoQ+BExpQGQiLN6fRdaZEKD9sSFdO9VyMP73yZsbisrqlZb8az
27veHFj5pwu/Inyba86VPbpL1ySKr0uX0o3WMEklN1xVp7s7u/t6qw1kHEFa
qEUuHlPZgQOfMcY/dWi4RQdezdv0afpHT3E7BsQdBNexFEapG8htpUocNWkG
czNwz7mrY1sOVMcOasGRO91GPqax3pOTRYlFORHB5gg7082t59nZ97nrJrRq
XlqITWABWdpRs/Zbohzaw80jgnvE9blIn0WL0Aka6Jiuic1IBif99RGs5t/b
ftm7ynM3lpgOiagrve46LfDAvgLIvE9WCZtt2pQYCoLE2n1whcQQDOxRnevv
Kk3Lq5zsXN0FMm2x7pUTX0J4Q85oxZYHIWPcyQNefZvGiCuF9Uafz98ipae0
MtqCEL1XMCOLhExJH2J1VF+ww+N8BnQAEkHN6qrhZfJq2BEkYe+1msC8HdWg
DyCoo6YxPI5GEvEJA992MMGlWbXsSffCqh660LCju/ktLreLR4pf30bLSLG2
JisnLTloKE+z7kPIwFDEQ29gp6IJ8Wy6PPpnTixen8Zt42H4JVUChMTiYKyq
aGmAaUAeG+ZT4I4DBwDd8d+GvmJe+SZOt+mcvjn3msDV+71fXndpKuOy8wpy
9Yb+TiwR+NTnp8mxGn69nEcGpnvM1ZhOHGCreXgwsuheoVYAUa9tasz5r5K+
IIwxy0OkBDYkEKr+DO9KgoWXxRRwOMGxAXdT8d38Qe1XyODWcM0m99ZG32Fl
PkXjGTRJcJmOBcvmeO5rNdPGibXdW3fD/LRfMxRUb0efD3qFQwN6yYR5gqzN
nyh5uKDQGTFTBr1MlGjx04lct20uHyi/+YpIgDkWrM8eF75vxGV/3RCvJedM
uYtpcDnCo0pVKdUCbDBt0Fa0fD7A9IikAB/oXk7zd+MD40JkxSLkKJmIdHLt
lJYuONagK+FaPx/sFpZ9FaWPdXwL5TTboADKNEEE0/aYMKSRxWf6cUD2JjJH
xUK9dyEeqyAGa9JbKzin2o95hxIizSGwAHtS44oPVuTR18FqJ3VIIN84HEHG
X+gzQnPnWS4yxteHp6Tuwc3BBlqL+fhUHXiR0LuJnpgjwYj/hgrguVuecVeb
KBN+WNhzDSuHodYQ/jt6qingqFRHYNwTn87yy8UAZrmi9kHicRaHEfo5p4Rg
o2xN5LMBKMZMSCT8Xw1Z6F2XfAs5M1xTlHcArfO90p4j5ELwYzgDu5Yh2MTc
K55IOFAWNXkDiUrADH9kBfWYryRN9SiaSRZG1A2s9QwNISt+ZEcI8whRMngm
SkdwIsuBt7Zl6e+MBLsldt/1k5SJm9+lSCdzzubPHoKR+5JY1rIPpGppj1DV
b2/nOsGyzkX2dLIG4wb2WZLZt8B+TeummeDChnL393RTxlfll3JX7oS4344n
l3r+Kw2FiRIz4P+Erw7wAzGFvA4qbWccHXmNLpjJf/MXUso2I+gwn3FX4c1+
Ff1lXwwf12ulIO3idJELdrvoyhNA5kjZB/UgzJebCYpS8bxqtba6SF9BsM4j
qBoyo3+Ru2j+xxqI9w/P4EiQFN7SM9AxI9T9BxTgk8yJrQh4IakOP1CTiaTV
nmJopCts9mBVJVKG3ZgCzdNu3ioPHPuXMjUFj+RBbqrS0mideM1KLYq3JKVy
477L0/yXqu/XaQTY81hmLiYX7Ht5G+WZfEcSr/XLaqAx8NmDHKewAKZewpPE
JBmHlpfdOq0qey4k6tIJ1v5qpdZ0CWAZXo3j1BGnlCJ5Ou3h1rA7KZHE1Nyb
f/5otIAWVtff5D8VSQbEkLJgoKHWDHOis4KaqkNMP5YFAdqmxdOtH7DwLwh3
Dz6skECHd1em+BgT5JZOxfKsbxwccocE9p4SYf2K2NmD7dj68k1zJ7ldikjr
w+PT0WaocsJCIwL2wBAw28gwIhjk92cnZhT0v0oQqxguygtT82l8tFeatTB6
vSBPQnilrgDYCx2SeYVjhCxRAq+ZOZWNxAHZCkPtU16ZalDPTBiHzq2YsO9x
65jLYOtO9XSywEtPak5F1iYENuenhRQKIbBGLYcWSWUT+O7iQclYrO4AnAAY
lZCD0qkDnCamZwdccS4Fyx84agWtyNBMpP1y6lBNNnkAu5/Jvsok5VjU9g5e
qDepldYkMrqjg8CZzW8ZdcOJuZrJCexaYRVUgB/CA0s2NpfPWC6mMamHWmX2
x+z2f48wZUQvU01rJicyCSKoXsxSQytYhZYk9m6IJe0U4D95fiZiYJKANf1h
i3netja5h/v6Ppd+njxZB0UPI1l9iN+L+FHFvRPHPw8lVH188XUICt7Cn9+U
mgcgkiis+OFkLDwCCTXSXORH+DWrB0HoydROerLllwhTskaoF4ifdsfmtwYT
pk0t/gemSfqSI0mvnrOGhJs+WAMaFbFtozNb8mn2ql4J+FBbL+VQM3B3Offs
h6FH+WAgv5mWevPfmp9UsijLu9rkVd1oLv+c6sBy/Hhi4gHY2DjR1JKTM0ff
gCwJvw0cR4ZsYeVUQ8uLKLJGjRjQG7QC3iy37m02adoJRh2Vkqrv4Mm4t0l8
fhbn7Db/rvjMTdZjDVFgr7lGCnABcoTkrl4DSi3dQbnoadVb6oyshSemL1wu
0EdM1+Le2pYa/4mH2qGhIjbBYaEtuEKnYwmV6bsQmCeLU6IMbwESpJBOolX3
91H86/thtP13U7IAyikwyPhNFsPoJ7/Sz0lljaNSoQM0BxC3fSHaPSlf1HiF
77cNASvjPuYA3Nuxt8VfY40F9wfeWDuHPiD/OM3XGqFrQSLFomUWSETESf8c
h+a6eai8UohDiym1W41b6C9I3x32cUWyoTi960JTtswVhLSDIvwb2BwOsjoC
MEPfzDcLKO7hJZsOYKepSTa5pXQfDwjug+qKD2EvLAuT23bikaJNS0QfCEDu
eIHHqi1+fPL39Wi6aMWd9fouREDCYKfd4wx4Zgq/1oYPhIz5luBbso2L3wbc
/ZGM9dLrofcUQMbyugwsUw3wRrYAtW9jH2YrTEE2L3kXunT1XMYlIxhGzW0x
iGCQZDkW8sE/Px1CC5w605ptEvAP/6nwsiBarNkUkPh10yTjQqMAIvLNjuOe
Idn0aXVWdWXLEarp2dq14b83wrF6oBZxToVPDFa4v/CTZ/TFagHcxnN0XFEa
RDM4bFXr53gNFjqXXr5BlnGEsAwMLvY658El/9IKVoz8rNBeYyTWgb4V2tOP
DW9YmjKV1zqriRDCZh+QFVqsIZvTZXzYzqgqzqzXsvM0r+wOaR4upjqM7uoX
Nc3n1cZ3fwdG00FDKFvWQ5Uq1t8geyM8cZEEV+wlTqngaGBMMbWWAuOPebfu
FyHhbrRzwh8ZfKKkHQVOIVzjiK12cBfyipWz1VJPL9pBNHmRO6KJns1CrXiL
vTXCgxyjQfxhoF6zB8qR6+fwmE0MRsqj7Qp7HeAhWpYcQ9O5NqH+BzGcGt56
si18ykUEVrDPkQqZFcVPq4zzDspvTY7sKBuBv5RIntUXl1ePgLccL3VbQQLs
Nr5pR8mpnr+fn9fX9ys3bl5ts4SmiwbYkqcAR1HEPUhwIKZ9q4DvmxFeGY0L
Lie64RiVd98NMcQDWeFDt8V9+6/GbyK1+iRh9nCTSHnfGS38nYc/lsKrZ3fI
ZD0Sr0nXPrGO3qqwhiBi1SP1K6XxKuiKKSxiFvCxq8Y9lcNbODtOHBDEovX5
9tgx5pD2ae1fjUr/xEUPO0JOwa/fKqcfaZB/SctE+aH5M+czW1c7Oi8ZxH0B
lgc4S8+shXtrcxXkK+DU15X7XQL6yYBpy9w2axBoOB4zvjjF8HUd9cx+g1Jk
QbMB3PScejpZIaxDpD9Ikh4DR1ntp9jGvCo0GqBNLTi7n78CMcx6UY5TIChD
CYmRESOMQlh6pZxII1zYEOIL4by6aibKbmdvE5IESAC4muIz0JWz1EXRto31
HxgtIllNx0w5pHuiC/8zhjklffOaCwdbKuDJiksqYffKz09i4FUjWh2leMNi
XIPjYThydGtmpmdMQMv18+T7nziLk1Ed46YjETD1warNJ3I7Qg931ECuMG4x
URDWKvEh+p314+V1s/oqB1jbySvHaia9F1wBXY/XmDhAIJSQ6acFBFLGBbCF
Hs3y3Zoi3hFYUFLGtNsdgFYm9UrHTXdzyMW32p7ReibuAA12wI3EMwxjWMvs
sfQi6LaMM4RKKRA/XT1+nVZmv0VhoGpZNWEnE2bbPwrjtqNtud1oHtW6w1Cf
9/SNxWRiNR41Z2aN1FhsLt/mqOWNfxWwYdvXMVwJTUFGGpv4kZHK4bVRWj71
jmrRgGtAbovu9TW5c9KaP5Wu4IDDG4/IABHbSdNbbugqxyPJXybt1SUU+gAa
AKzBTL+UAYS+MU3YUbk5Yk+k3quUBg53Q8qSvkBci5nuPOn+0fe8WkmJRuGv
OQ9wJmTelTpSVuXQxszBS99MH2b4m6DE45aoCcZBcCVaQvIwhJ/JfJQp47Qr
ZyJLxZOXsxXJ6AJ8778iUY6yObsorwJivwUURUAbYEOQwwLrM/7lspo2Okhv
cIuw17vH7ZPdph28dj4stj/bDcSDtjNRXdunozIQmRjq41Ll6YEHUyWWAusV
bHewGqdEF2Ngd4B+THiZwUHxV7oVHPPsWT15p6eVpyLJyW7GmqQ/h4EMtoVt
Cdy6WP30pGdmwDtGPJ3bBVVZLQAki1eM1sPmQwwwC2F95xSFGI9X0s2ClsO3
diRyeE8YVesOF+hRfDLH3O68RCWOBD/XfK6YIWD2jkpy3tCoWxMcwwxXu4zh
jcZZ0Aic+fGJG0ta0q0kRSZFCvbisPxxUD3KMKUnssz1XUC/1Uf+pcSOP92I
lk0880F3PYlOp1eX/h1l57hoSh/AcaxfaIIbob8FarUlP3ja7F1uLe98orYD
6AolxO5Z40J9Sef7WlXT6tnFpQku1FyNoCwI+VEVgA6eoGmGV55GKmphVUVh
JLj7rpev055pBB05Z8KT7BEUXjNDnife8VOW9pbokrQGI4vXbyJN2QXEjTdz
4FRIKr24/vZLf/9OEMK5+OzwfSwVan7OUz8905lpA/ka4fpasefDw5729nZ7
YWQoCdCbFHT9RcqM+0vp/3ZPiHDa85R0a4KtZHzrN+9RmBlc9cO13ioFKa30
GvyVwgOVVRu4bqNzo2uunBl0aywQp9egb/vKTSwWb3HZl8/mYsw0xa3XZ/Kz
m1PukBphOCu4PDMh8diqXpW9DVA/jAEwIlL4VBtSZdeqBTF5vAF3px3U42v7
5opNvAk83BuWTrIoQPFXaHer0bh8f7rdxG6MerKvawoV7dvqU2H4DGZQmvRq
JT5AzQeQd9/naWmzsyeOxMk5fGjWbB69hixb1anub65Xcrno9G3R0NiVznsN
czr/QGHll5Ac2VCVnGfXoMKMEUBlU8XohX+GbD5XapACB41PQ9lOI4uGMrpT
6RuG/E1saYVj+vaIL9pEr/E9oqe8G6FIW1zXCuIw0Zqy6G/loprVZ/iZ3Iey
yD2+iR2U5jMSJVUyuOO+v6ZZpshF1CWb2BW7LrNdoFIhaMgXXSI4ynlF7JdN
QjefceKdV5go8GjZyQwxT/kfT+ievhHEw7KdIYmDGaCPlS4IhTPfdeMBDueu
cKugpMiJerzhdkS0oRDLVdvFHVnmSB5m4gl4jpBeCnVfd3nHCixcBZEV2ptl
1bjiJ6aoBVf6fsCZUhOhwicXjKhZ5c9obCSv/qHSNQ99b85Vj04O/Ik6H4CR
/ktI6WJehP8UlQ3EAes297SIzZ4rUBJuNSIyU6Rfhz4pO4uTA7G78MRSP+8J
UxSsWl5rz3PlC+kuYJR0td/wYhcHWieOm8LagIU+0ZkuUHhlirs5P7yz3RT1
C7J3lcNVEeU0pCIDoP0IxBqN/zG2BHT1nJi2kueOduydg57xSw2NTN2GqAXM
CNqKWSYAvDT+6kCgOC7GhZ4KkpouGyIyrY2/EeUFUG5Tur9a1B9XZQcxgI2k
65uWkikaAA+o64bURQIK5A19a5uzxJbHEuiR/zFKbw1DSro1HFCZJ95Vinrg
NsxLc1bJAc69hNBgaAl6EjJlTlkQloJ0W+PGhckvwGmt5PIhRi9nqA0QyVQ4
Fvd8VSIlooJ+gW+sY1dSQYtgQHlcZvbvv0yjh4ztmlqkKMes2JrswBqPcmyi
bNkVSB3DIMiMVUfVROVf6IlqER7O0+9V4r3n+dbtaNfnnI0Spif6+1FQeaCC
ItlVHwTvJwngJRMV8NmazKEU9Gqy7U6bni+zebM2wdadTuL9zpDoPf+VdGFN
wfH5DGnFfrymkDETVHwHy1r8ggbNaucuqyKIqieccUnXx2Z364DsXqwiK7Lh
kVRxeM/NDBounO1misewuSCK1xoYlbBghIh/sFELRzRqJ0ZYPq7lbxTFBTWc
faCfoFPpRPz+UwoKH9A+jSFpXs1+SQ0TMo0n0b97++aoZ4nkADUJRYlzy23k
ZP0Fbu+irV12/wAIzDZfpYIAcBKfqI3DDT5CiPsKwBWyqJlp8gwW5qe5C4Pb
VgxoO2sAd39jBCoNmp7gmamKerzjbK4SSaZydwECei4Y9qedk3j4w5RKuXM8
o/dhVFlKWIQCoe0q+SZH1kIlOAdd5fu5Gm3WimJeKCgo4fo1FSILCh5ReAfe
kRnfG4BzWnutQnXQAueQbSHdGMQLAhhRM41/QUw4hAa5OHxZ+szVdubonpr7
lUeu1H8KP8srNTQdGW1OHL01sNzqMx0kBfJIVnOV53vnyUjSQtq8cYd00CDb
SlYp8ohutmNzmj5O7UK5mDKRADnjaMXMye/GIIOsQfhH0kncSXVGOLthZpKe
ri84qOYZWnnbO+IbuG9N7VwSh1S8DWU9LN2rHHmMvDueSJcltg2RL9IVzQXP
vE76rXCr/93G9K3lQVqQOqsHFTIDVciY4EdhZ6Wih2VPYY6jFjcq9Ks7sG5C
rFDFi0QT7AKRT2opzuKdfEmj0zSuBV5VPYzvbkVwSVRobFc+xgMuSrTLsguK
LP/8Iqc43rP2V4h5oQERjjxwuLSrdwDmaZfJSvaa94/N62YIyua22c4Oz9LN
aABszAPH5Ttiw1DYhlcsE8rLoGLZziCulI+nmhFEzGKnIWUQdblx1gg+Cywx
a9MlVQ4JbEL51AZcIBZKDAqaWCNlCuMKZR/GAQYyZrPgRtm1sq2vJeohiavV
XCjKWr20IxVIhYnvAj+cmqlcDhNzObwdZv1hZ35pSYRDOA0Nr7FsrPX2LIYX
7ETNe0uCwW+2N1UcrDhpgmUiD977Z73wLOjXecu0whElitGHHa+BIfXQ6kZu
0tcnqaWrO6Tfnz4aS6WDIxbRde2Zl7+1eYzH25aoDUvWys1KgUKOEHfFHkHw
Y/Ex1Pt8tqcmZ+vSavyQfRVC3MuEwvfo8ffs4TUhdytQ+5wYHwhvpkxANss4
xy9oxH7EHqnn+WFU6QLWV8yKRfOQAmG24PIyOoAIUkoZn7BjEvxuHbkJv0GV
aPRrdmeImgonaQc5Zr95Fy/FL9cEB6tTuVCLfe4xXw933hjY0AupZ2M7QvfH
Sy8QyqL8VViBmeUtrkvyCQYNLuf1U8pwiKKuVpgpQg3BJMHuZvi/SVk+DBPC
6NjVPFtvJiAfkLnBOw0de8TEtXXZ5HEM1SYtH4q05jivFcx4Ypj9qElLUFKH
Q5qkrJQy/fcwc11XpMKsI3eZF0tv/rLRiqPTTtlCDmXLymTQmP3zJOPOJ4Vr
NhIuz+w4xHATvUm0nYbtUoH7FRcSjl/4G6aHgd9h4VP3B08ciZFWTxk2pEsw
c25zKAb7ao4nCw2cyZ8IDjtgc8UgPTGSkwpMXKMXXgLTJI7UmBuBrohCjMKn
OI2x6E1ntKMK1WrGMXItEVkn5kMVxAeLKQuRdN6+LiO0+881oFCsVrmXwbHU
GxGAhG3dyfqdb3uA1vYjxbBL5wC+oRDHLM8SJVRtOGHIv1lYPBErhavrLTfr
3f84D9ywYOsHLsE8oIlSOm7miieDDe3j/0quIaeKL/cPIMY0ECMjA6c6JiGF
alGnpfp/JFVrg/qZ26NpWIrn5hINPWaa6v1JLfKMcvst1bzdfX3bRpX1cu5L
gSKedZ4yWgpi1yupABUScDB3/UWrQpl5No229m2ETxQNI/4FdDDCyRgk2U+b
UYBYLMbZ3NlNOHHWc7x7rET6MtGkgK5VV/POx1JKuvQshS2XIr6K0jMmwCZf
XsXmR+4KVQCxDJhEO64/QQtc2GqG/1Ayel8/mA04tRwilHkKHRU4nsD6SIE8
27zYXQfmDmVrKe8mS1cj23TD1nz+EEv5vD/8k+JjmK/7ZmpPUh/wYIIQSoey
bvyrps9bEPjsS6OpVLjcyN9OVxN80zSWLpPi1ZsxM17CpxVK8eBAnUfg3xQx
0yPxwc9mQNLZEWCnDhff4NJEarHX3M7gF7PodpCH/GSKvb3kOjfhNYAmE6DR
2EGvZDCOf2nELSljPNzkRU/XnTcrYhJSFmgSj7CZERZx4phfC16A2MgejelN
Uu1wnWbBXVclGlJEZbTvbhz27JBwLXYyWKaZOttpfrKUFERHyESrX5TBxuLI
ejUfwfIfzcfNydOR1Xc3QICcVdRc8U9LlhGX/i8fHj2cKZ/p608E7MIWJlgJ
BpEaTRzOCpJLrIW0S4k1uOeepc16BWKh+c2kzN6kfS4dPL6nfD7EqB2G+5Qo
2EdyLzRa+4YnGJeP2tDYqf89JVS4+S0B3XdZLNMvaY+l2yra1CtEatV/zuIh
mFYhSUETgcwbnhSii2MjGzidvi9hPxnMYxu5NdMLpvXINHq3sVmHgIxbM9ox
SQfxd+krItk9O88QRjKUz7rrAQf6ivWgCLV5VLXO3zKr8FYn9Pt41/Hl4GlA
NW8kqtA8wzLnOcNF/HIzrXZNwhsO78LYo2ncFmqaorv0xfSEMKz4aj2ua0MU
d0Q8KAVS+eHqxS3ayp0xDv6H1maE/GqMwShMcB6ycYhg2++9CE+PO7SB709h
2GJR8z6gx3sIIUhmgzbv3tK4mN0VQJ3XB8X3o3CdPfouhk+CvcaBZYvwzCrQ
XhXnd0Bm7VAQp0hFJep3jtMhbeRKTBvkGAgnbw881Djvqn/2YlTP2ZHhPUDM
x0gvOs9RabJWHiaZTGIzf4YN1VPYGvck5C5pZvMtBhQQl3rM9m+GrdX7qx9A
+l1w4KjsV8RspsxgfyCGlbFRoGQLjRgYiyLs/0tLcpSNg9ZurmkqBhPM1QpP
AuxNzWC7JmoVN10cRGKp/ZR/T8Wrqtzwt21JV+irr/FZkK+wmMF05CrVv3ns
XXlOQ2pdtFcVHaYxtcMfjambJUm8ouEb+lNaSspXlYOIPaAdK1lnvxQmtHwV
0anC0QukJNo8LjX0tPc7Fpa6XMmhu4Qz9nq/LOTJYXR2b7/Lc44qVKJTImQA
MSKd9dsGHxLA8/dJQ16ojmxC91eHOExoyM/RcKzcHyZ/OkiU4ejxAG3rBJYG
C2x9q6pasE5gXOuAXzKMsUq3YyCNJi6esEaY9gWdGFCCgG5jIvgQ5611ql3e
MkamTUWmVOmNBTXYZuli8Vhs4090u+ugOaRI45xEf8o7SgPe2aJWOdXYAsnj
WiLgqT4aERbJzK9eqXjQTm7yZmD7vBQjlA0vHA3YhR3c5V8wU/t480D75Nak
6MSMWMQH71VrhAKfOlNWkVETMrTmcMubQ41OZ9570oCprwehibVBAUaWaCLP
NhmCnqOBBPC5GBsODlLXD/C8M6xYLTAkSIbE8Q8AKL2QZTZeew6e1CVRuW0A
KLTMmgwP5eVK976xlZsXjjDMPYLA2xI2SZPWvXaSLy2MZCyZ27bNMpqRBxtO
hh6Hh7NLHlGkjMxaUaB3YsNyNFBN+MRdNn271qrP03rWzuo9G2LyO1egDe6U
DBbaNdJBCmKRA5IyfEh8YfB1fOcD5JQhAFE/qQ1SM2g1+c03scO/ddiGEo1M
9wbrrG+Ycxn9ZWUC4++oZ00SQz/q0v0MZv700hGA55rYuEdzVbmpUyZt4hg/
tqoArudBXjgYEQYlJIcWEFCTO287YRMvbzEapaaWxRKaHKbGzVXl+Yu0Chjg
gUMqn5jK07k2a3wMa3J63l+YpsdomjeYueUXjJCvxb0hnnme0Gyo2BLE9T9k
MLTRSII8dOSKI6sbwuDVehkFNdRxBiwgercOmAr93Mg3rcj+43Y7R0a5Gzw2
MsArlvTDMmnu97XafebMNNM9UIJttU5wKDO64rrpq+fxqe8D4YrWvXAXYNPD
tiDWv58ZHAoX3ZNGTCYutQMDzh4LTCnGtCTFJu/nuMKjqQhjeuC4LU1rcuF2
zqDW9qkikN9C+yqz8kiP/hDLi8OLzBmwARUBQwdSUc7xvD0SVdUcelofoQRH
jibbRfNerOZIqlQ+Fewrn0HRVS3yQchtD9NDI9D0dBTm2Q5LLOf8GWKEtK0v
nLc7PvxAQvRIzum1OqUxzCGmT1Izs5MfnEyPisqi6U55qvMgDz9szAabU0xg
rQpZ3yTnVom4kaO3i6e7/YkrGjgRhiXr4nXSGjDZmLzC7LxpiQhzTspAXsb4
1PuyUz/MXpsnONGPX4jCExjyJ7jNm237qR/iygNmjlx4zaeY6mbYXndY0+B4
H5gPbVBZ8ghQB96sdJHA2g1hn4ptGkFO7r9TwH/FMwMhixXqFq0MJhFnp4Mf
qY3mhhghFZdX7ty19XSmZL+U5+Z8VKF0AbIjqT6h0ECf9M74ka6SzKxbt45I
Oa+/BlnZFffFQXqmMrwzcdxyXwI6AZOIWpP+F4mLaOoubKoY8rXhZ7fZlsZv
MGAa7nzk672hNeZQYIu88hHvgKiYdTT1NJaWeiqK7RzcolSQMeEAbagJy5br
9oiVSnKBRuZzz8CG2gaikfT63konXg6MBNepuwEiV2GvbLGAivDp8k00sufz
fk5Ka6Z5luecy3D7MOMGDilRvVjrbRO6e8KyaUC6buEV28lZtRZ3w230irV3
aYr0GKe+iJ84NnxgG2v6Q+h49qR+/RhNN8lRSv7DeMqBn8eK6kHl4ThYg40N
UAgNPSFnXDBKjxbgFKwKEh9GC0p+LjCB3ZfAkEUWvRgYBoBTPKJmdQdoo15k
BWyBjztZ66NxvtUFMf3+dN32N5LRa9Y2CLa1guPT+7Xiuffag98UakL6Udxf
07birmBnYxvy5uOdFQ1CcAnEsZ2UHQ7uwRQCfxwysTwWTk2Vp6D2QeKnt1PQ
WQVpcOh1XSRcclse5tX9uvF9F29x8LdNJ0gjw709DUN2bqBbi61GqBmOvvlX
Z7r664/q8SN4/7Y3u+4W5af6VVZ6z+WHpcILfV5gZTIoJZYjSkbWOX/ptrbB
gP2tsNJbho8UJ9rhhqZWcuBLBoXIzNhC72nqeX7EkIOWQp87gLgMbAePQfPM
FleaVaKt5RgjNQZS2j51nyoGTVO35ign6/5DvBWu8LMHvKLZq98OSMnI2hn7
qSQtcXR8BTKHQ/k0sTrkO3fgYZsTwhmev2K50AA7o8Y7ZwDy+YZxvfEW7DtD
OpKmjJPXY3IB8HtXlckcKqcmRNdqskMmqnLbkc22q60gJCIXreFyI9vz/Kwj
QjcNS+4MKwfdKB8i2KFvnof68b37WAF9i8r412NUx1cei+40EKYQ8o0hIFl2
JG7QhzmI66CAGjwnf8u9FieryAXrcB8U+ScaCiT55A0JN9kcLujqK7Dhe8YV
hJCkCkeuGphPSWX8E4bKqQYZnq/Equ8d3G8FFNKAXdXcwCCah0NuiAh8wgmT
5yb2IpFdINYZzRHagsXBN5ytceC5H6Rw7fAEFTCqbhoGOMcItP5ArmeDrCIA
0m36DmFHBh8NQSncurv8/+4PeKr1jrQb+Q8AAtBpis6sNR1f6XcG5dTbRG89
+C7fxFinsJZVFeC2iOLb3xnr70SP6IzhKo10gIrn2jP8g3cXRWNGCC70lDf1
cqvjBXKm2qS3ZO+C0El7SoKIvqDXLsttUgBeiDli0OTwRSc56DOHCNukfvyw
TL0q6m1x+1LsyuYqWhHTuMz/5ZFhpPbP4ql8URcjJ1YAiDdYWHIVD+x+uhSD
DknekQV8QdJ5U3ybWyPhGuWQmhYjBwJqjxG76wRHGnzqL9mBE9G7GpGYZgjb
SR00cIkWldvZ8qgV+zeXcjK+fDsq/GKZTWf+OfGmmE2kiOzycqnEqhnmSROj
d08cK8M5ZbRxxiesNJgu11KxJQo1+N6pJazcTdLv6TtmpGEjpSmtY5Znz0jl
VV0WfxerV023tJyXR8+tujzEV0iy2SQGg3O4JZ+P4zeMN88qYXI8xJoavu3C
lGV6p0tyCJ8J6+oUuX0LYgjI+vXFIuUBcDunBIQwp/9wxxdgHXiy4aW3auMx
FtHswpA8QZOLzbFXr20unF4/RDwIbYfRo1KhAWRlsJEkPm6XzjfScA6SpcI+
bkW2ckI3BMZ8py+D9341plmJfupRxZUNnUxFcTuBb+iSIUAC1cdxwDDIJRYD
aphR8eaKPygnpqZreg+inChLV8BSlQrbmOAiUamv2RA1DOLPnE07AsC1MAFn
DCGNev8rmEOPZ38GWbQlvZIVwJYqKlyTh6jOIQfH2FjGvwclKEGVutz5Pbor
jvkgrOPcIwdwMewsPEkmiMha6hQ7ykP1xMM6GDUPUILCkZu2N/7GVZTF398r
D4SdxDsSEdba00x+tzHltr9e7EDictoUeryi8KoBsDnsjmt4UizpRBeScZBg
B5txGFqmRxRYFHP4TiDjAdedRSkKkvhh6wOsdFO1F8gc7RdqWY5DKVQlKvAv
SNgNaRacKtfu21StrgAbLn9M/SwDCNjfJJuvzH2XX79euuvdhYzU4ofW0ol9
oodi8bxPSPuVuzcR8a2lq2haAbCXJByFu3BstEcgy1UkvmNLYjyuS8M6sCrf
t1s9UJezjvzR1P0636ekuPHwpAQIBxIUrWVIZfOC4eEEeGXcaXJlPuUOtpYM
1rKtEhaf1CwwW5GU8UxFP/nUXVQ5oxyeQ5GZqEt+h3X45/pQVxvH0VXdp/WM
zyz3wr6m1x7+YqeHISu3PU26mB0BSWIgl0ieVv422qIKT5HcytnD6LQG+kF3
mPItZqYN2SFFoPR5D8hWcChAKq8bXJ4pKFnxpghFIcp6wKPCBTklAKvlmNzS
7WScee2L+EJDwDxeS3Ts4Tw96HEhzhyLYr8xcXBWQHjhJjq40NtXwLyuYDRv
lAHyR1Gofh/tnUr4Awmq0IdBXtv805vZQRkk737BJ7idG+gRquvdp2lyayWR
n4IN/Akgs4o0wlysdDQOvNL9uHuS0tDZBs8JHSnj6Bdf4ndaqo+prNaIbiov
m5Wjck/R+hvDfkMW+eX621qUFr0BiYnyQoDVWujN2eg7W7wm7zah+l7MOWu6
70YnsF0g3dteJAZZNzWM8XxZeshoqnNGW4bdTY0jBA0u3JZSvvGS2FfH7T0p
IaXgE8KBCmMAJ65PTbMefr7J0TBRfQO0WyM49JOxVSsLuRaUlw7M6VhISmcq
WK3xHtRW/MpGZ1fHRiDeL+7XzDJ9SP8oNgpDcfIsd3aMvQ8Z223uKblZP54n
N4bKHx5EIfnZ9NBoi2QfFSyZUBAfponoBh1cOC2ozaDDF/zYKi/D3sEPzVSQ
CPpTjg+PZjIv71ahru+xUJYz8i+Hk7pSJSNVDdvyMomz6K+q4L6AIFLGqzz5
HUDx6XK/55WHEj58mXWL02WGMW2pufwnT8UVehqyalJXJgvbyYE6m3quwCJT
hx/hXLdfc8oK2LBVUatp/4MS8j7I5ipYbvT5l7kr+xfG6PRGUN3Y4j7SZxkj
qW/RJvaVE+5bRq/dXx7pjxS+9VyziJ19IZZAIyK4S1HPcjbg+PVrr8bWcEla
/3krfWfZ68xhvA7LxirgBx/urx8ZIPuYTYUtXSXL7OylCWhiKWa5pAiwW57G
vmf9OMmJElU/7aDrOkNnoPiInf8ID+ItuE2li2eaAxnDidS2/nMBkoiVYZuX
mqn4kcHFgfOYrd4xifSRsIW8j+NzEOXx1XQI4hB7YcTn1LycAtS1ADka8M/n
PIWdcLTJWN9L/Up+sv3GlMNnN0ig7uM2cYaYlDSNi1MS84gFZalbBwKjD87N
TIcfMwOaYpEy72xPVdpS7sJpIm0TAxTtAZQWl9ONy7UAAKOfOSxjZA/IH8Xr
jLm8y32COgTNk89hzzGXBxSrArppe81bFs01+hVdzh5T1n1EiGLrBAmT27l9
2qG9aa3GUtXehGccRSVoT1z6sWBQIFgZbOuQhr81aLMgLqva9OLHw8LhNXQR
AE+8tVBr1a4my6fLFuER6ejFa61SffPjbMqkcyDxd+vrsCLC0Nbl3JDfxWpi
aGrVIyIeoKcIT5swMbm8IEXmo2AosJkr12bSjDoLETTtilyxOKP8XDxf5Ow1
//OJs1dZjVXaC1KKmtllS2o7JQP8/RFbqjnb1EUaD4NZY1eB8V0odWGWsQLk
2DrfsajsI1uIYyNfCc6L6zvZAnZuoI+xbhYjs6BNaCtgjGwzdUxKfDvYpgkx
aNAgXReYBgMI7PQrlHcNJds3YC2RVhUX0y3qtE73iLiSjDmcqprVIus/laeO
GELoTU2QPRzcvTJAU4JVIxbW36J3rYGJelbFy0pMCpoHCcaBA4B5zx5qCGRU
EjJzFoDwhynDNQlDmegxB7AYcjc54CkIaOksDloGF1RRCbeV3LtyDy29MaIp
54GXPDcEP1Kk2lIpxEVGsY3FxUBKUJqCX3Rx39gQEkBO7XAzqYye3mcbJ/uz
E9VopuseC4rnukdx4/OBkt3jWEgK3S0nxuJabuaJEDYsKRcjQ/S429CZe8B4
6X3SfXLJOZzdH0r6LArFzXYCxfSzTd5IaPdkp8cWm7CG/EADamTG1a+99YLj
ceHVNGYOQE/J+I0uKJoc509wPuteXpAenTZSLeXnVCfhiUbouVw7VDca5so0
aaKgRyXMh2LPdobaVfn9RDzqnbyns4r9VGKbkJ1dEP6sspYN9g4H6Zu3D0QI
hDmtKuRc+ECjGQ//Z/3wJbuaEu5DlIpkEmrwX17HbM/pH1wLN0tX2oo9IxaG
NBRR/dMYLB95DxwU2ofYSCJbMLcF8Z3rVmmd4/+nQcE8a878onOSCQammWQM
TScy3sHWAxmQu8d+ys9a1IvrKbhAwKVQcPV0/0s32zvAK7G/3rSVbwq/WVrf
9rcpRpxyX7pdIzhSLXv0mzFz/iXSTElmykcevVwtlUT/REvfOe8/MXKiQktW
sYPOX+nB+mAfEZO7IeLjw7S/ELTcWZs41a2jF3YuaqMOsrr7vAclEtFMxpch
bPNABh46SlN3SoDiAMRNKieJGzt1LgbXY+T40JPX23L+8tg9GvSzWJ2AWeeY
dxL36dG8VuPj09+zBlNAa6eH+Az8kGJiFSxBIGuuanYLpfkXvmd+kBLe0X6W
HI2RE3bSeimkHCFxdzne+M+OpnqefeXXi1aGk8JMfmu9Fu0CmCCEe9ZFG8IR
crxWZSWXNkj3xxaTr4U0sr8nx7eWBfULVHUtQD+i2DrFXv56yzaaux5kV0TE
B3Xr2+SIsEIkartIkz4QfoQ5C3mhBIiIaI/Jx76h6wZZZ2g29yIdbuKJaagg
6/UbH5rKHwsBxq0077B/JxK46/uczMY9qt6peA4q81eHjM1HDBGywnJxVZAq
E/UmIR3eJo0mziCGci6eJYM+kyJsl2Yt3erTEm1IBvWUIbnIpN9hVoKb7fKs
Ha+SV5lLPpQCDnc+guRFr+hWg7GlS7VgvoLrIbKG8ZqsPIfzKRT1AsNw+raz
2FQmJmQB2T7pzmk69gAKa1DcPfOEjjbHU0a0E2KmY+TepWqPCNsVB8RMCDit
Hy1zinfG/ASxn1VA+JiytXB9Vrg9jEWRvj6yGd9C3ROJiegcAOVrzPH1EK/n
SRt3bI9IMsRRnzY3s2V7Ju9TelqjutKqCkKyF1HkmIGUGJGqbWJXWZqBUvV0
UHO3lt4Kv6xxuiw34g/nshc4u+Vk+niO6hJO1faaFPqIceL5fy3+0UfTznLV
Hh+W2Cj+VzfzCZDl7x/SLaMvFefTVyGnKvCtXOl2LJbrl7GWKVjop8PxZjGQ
PyqcRZF2yu4xSK09fHsgDHWcX1fnK5QwfF9Yfs+vBGW36oPbaZJPO68Z0KZE
fpE7aCpz9ITbthtfa82mcdMqFH/RCpxrGZf8oogBeto1/A3N8F6kVwIZkmq0
rmV9I8kh9uT0Zn2UHDjxZ3uno2ktT5ew0Cr7m7ObosNmcaohkqUWhtLDdFXw
KH08lmho6B9SAaXwz8feevjoDuVfgdmgEcINmTd8UxYI84sW2bD+2Jvp/oEh
bcd0t4dDf0NmOk6ZqtHtF2TkigNd/KZSswyGs03+ZU3ROi4nZHGvXzTnXClo
7o8G/CWdR0BaLRerfT5dLlOB/XFCn24KaLwCuUpHN9qJhl2cpu8BdFJtDBsL
4E7zWnNtUw5aGq1aKozOZRnv7O6g2UMgdddfV76stwQ4wwvBuXEHzaD3Q94F
4l74GldSpGhs0oeRqTWhgMwRrYoFv2cb73IbKyrMxUUK1fus61+d54/4AStR
e8qbBOymA3xh95IGs+ZReTL77u0AY5UYUNJf3ueMe8tXVXy2JHwzIB/ixFuG
muVdPqGA8DXeMfG4a0R9WdUl3YBfRGBg988VhDVcCG9lg4BbmG0c6sVUchW3
lyMyngFJ7bO5Ap8UvVJITpiOMe0d6wsDypA/43WbDP5FNZpOlgPhPgsyGepj
7vDopQZ/GfuL0Kn7V0zvH9e4DDbyBN4rgqB3asSRka6cN+5HdecknjTsUX1D
3Rs4so8oNCPZvsOTI4uO7/xL4f/Bgve7tfvoQa3yeyFUXfSb7XRBhlGxrmLT
mGWEAW9vU7w3pej7NxNDo4vS/6VuBu53VeIbGFoZCvHpuXiEDaZRLi8K5E4D
DdsQGeNLMB5/Q4aAvCgRbrDfzaX1lmyzNRBriadqXGHRBhWVosXY2vwYfvQv
LoLjqQLMx27qksY014d5pIzgI4Gxhbp3C6wDzPdAB5OHirOZHJvY759wPyxk
D78Fh2QZL5cBpNOqvfCfKGqyDcwE970xDC7lXBUUmVf7doUCJOA7OGwxAIc4
J2twLMLYqTaXfuy72t4oY6m5zEMnY31z2uqbArQjvOhkaRPF3A/MsHQ3MiZE
9zZs5aXMYeOAYWUoP72MaEFePDn7N0sQWC6ub7duhnrlQCP3pcKlq69pcxfG
LS/r3bY6+VB8Uxe9gTYHHkndXwryBq+D4/Lw3m9QO/U0M6Cd5E/gIApBk2Aw
8PuNirkwLaTOfFrbT3d4BG+/3altOZy7tQrYdr+82IZ80AQ20ajVwAGWjK9h
1vi+/CFNknCvVkOMvpPQhyqiVwYbJsDBSydDO6KpDh+OykaO164BN3fZDSqw
SOsQgnFT64asUb7GqB1GxYzCp+4NTfD0iw4UjBZ93T06sQRvId0Ljxm1UFZO
JEOq1LHHrsk5G330NaRHU0LT4QXS7ugxCPUJFRcJej5JONVN5jxGea+DV2IF
2joTSDOVpAi9SRxuhAoK2jR26VYEOrpTw33cSi4pqcB/Q+8pfLECckKJ674a
sOXuSxSHzJ78nbq1Z/uok/VZkw8DgrHi3EBUNK5S+YqkI5LUf8CVnqzBOcJN
wpPbIJTPJrX+6Ij46AE/lHTyM0HcutshRInoC+U1tV61s9zgEjs2UyuYSjEO
9mqkBuIL1nSEgXTVlhGqfvLbY3sEcuEGKlqQiOWe+KbtaES5tdqluTxVcnWX
lwXPlj91O/MIzfdgyRl6JJ2Z4UjKOgFG32oyJ/rxV2lk8A5+JlVN6q/OvFFk
FV4QXUkHQtfflZOmKzQxpdJx3nWMz9hENptDLykkMiG59jISiL/2H9N0fIhw
jO1ZKc3uqphqKA+AzDY3vITq7iQ+VBzSHC3ovzGLCFwMuwmQPNhmBQ0gdNF+
SeLbfBNjHcuTZ2+/pa2unZ00rPSn6HDC5lYvQw61EfVhy6vQL1plQx/jA1Vb
Gq4dSyM6ddamfOd5/sAY8g1NmbdL2Yc2SWdrpn4Zj0ppciTjs4piuvcK2sMb
UpGfrIILmyhOGxtVfrvdvSPW0v0gbhme0XTUJL4UAgEW9cdDA6vLrHEtO3yQ
gwUQFfnjaqrNGnsXM8TbhW0scg+PF+pUyJ2q7r0SCPfnfXYCqh5lz2nGJOD6
ph2hdyZjW03kli54xdEWatAKDhILeC1ltLnsC4mphOCDJ1nvlj8K35sQr7UG
hTefqPWg67oxshbuxT+cuTQjyiZGC8Y4zMa+7HMNYFNiM0XbHZQDhFGZ6+tK
AqmEoE74RGiYidJGpWEwslqrUdXTm/xCP/lENcvFZBEgsY7Sqc28FRcKHeeZ
7LvFh3k7lWic7RhhdaV3/Pmt56tTbucXpNa4+UGdTPlXqb5cVAqPI2/Ekhod
qmb4lifSJXrossjCCaLmn2BTzieKTNeWFrhMBmw+sg5uD2mH53BBat8QTo+s
+w0P2WS2nmM/iJWJjadQtosQFMzo7NwzcCfCmlwIN53VSlTjPEQH+wLNvQeK
wMnYG0WP5fy0+ooQKGQLktCE0NbQI0Nz1yGJDvIPcsEidnhJlKxFy7bn44Ib
oXY+XhD4niWfbRB2aCjIfFnka+uP8WbgXLmQISZjmrq9AJ1FrQyslWLjxoe1
66VYLBBFmpmi9ORI0iqb/Z4pDlmVwv/hDj+huBqM2Ch67+C2KSvHLxTKdFRH
4Yx61LGY4iHSNsxEfVtc9Qehk6d4tRAeafDlWm/NDR//u+AH2x/+G0hlrbWw
0Gxy4T+ZtHWzSfJn4gmPDKTslkRoHS5abHu5Hb8u7n+znmTlR+lxVVitgB9r
OgBEYLyypYSoUH2881VnEs+H3U+KUAfQiRURRIh8367qDlw1TePioVTplCpP
Qwmee57UJM8/To4IEtJX3q848M/ofAbQmddMHVqpTq2nEkXLD62NbYEWpf7A
W13yNsJZOpklN9OPmOFgypdnjxiD3SAA0fwnelJLdyvvZgIQrB4f84i90C6h
Sc41WxHDBI9uQ28i8aZlGRfiBySP5WTmRMOpyv5W2R4u7ihi+u+II8unPmky
qHoycle57ugnNfb9VMA9XtcI5VyRh50Dhrww53AFpAtb2xQGIY2zLJo79eKE
5P21F3wycIqjU0HkFl6+pSGHP+ezzavVEaK6YAF7h4m94Lija3CDrr8VoL5R
RGwo4vEKZqr0SMXT+fE2uOEnUpSgbggjgcBZtdkqOXaIAiAFFdCKkvEFS9wb
DFNsoD3mcQSopaDwjlMSsADTK3fmMCZNzVRLTIrPi4udumuDQk1JQVA0pL0e
3846ioj3wfQkJIx2m7bVLB6g3eqw+6Sj9s2nY1emPD/2OSmj+ld/jUllFq8u
besJirUzDew6u+bkilR4UmMMp1zdgBDrR/8JXo07vuf16ZX26I8J97JzNHkU
YkTMqxGA19TvWew0oNRQLpcv/q+gre4dUQ6p8HqkbeMr2N03I/EcAKxrw/q9
izH4U6S5uuRipO11IlqwQFx3+kyxhvITGvfv7i/nuuxAZNNmhOUQa1U/x+wH
bZdFGEc1NMy9zHxi10vypFrLp9nHGZ1bjgY7tVW5qky8CMukffo/K+TYj6X2
IgtCDkHTkDK11QQ/4abCBLYyEc9axRqbXiXj87lEcOFju+UN6Lv1qtljQjdn
vG+lJGkWI+PJRq6gfMvMR0JVV8PcdIJjuCPdlHgTQ8bNMvHWHoYerrvJu4dH
F/9QEEjQD7VcjQ18Gfov5l2SijyMaN8tRSJLwt4vqfdDtPDIqwpbKpvH3Zv1
kXrE+54y7cBjwdFWCytAqJneHCHJUTIg0RvY/CH3QWzwlda7sh33LQ4fW02P
oBy+5Zr6rIKhN4XsXpeknK5fZgCGTQDcYtAt3xbXwbiYs6hOgCdMNr5mDD08
Un7yoML6YzIBE7qk/hXSrzlc5ZSg/YAfgBhI63U1/nHEorgc6OabIoq5HJgP
j3RU+3OkEwZ86W8ncxgfNyaOa7ctgjd7nEWV6OZCQR45b0KzWGGgP9Zca0Vx
eQtd5NDSO2UOWQvGy48SvOzoG8svBPTj5T681E3OXTEhs3Sj7OPnad81SnEE
Pv7GhxsiFeCrwEGUQbqAT3WomSbuYxDC3SqC99j55AqgyNAVyj3lwZVoTNua
j+MeAPT+AZ05saJ53LJgwUiA28E9BtArrIVfdkMIaQ/EejlH8SmiTgAZtD+4
drnSEt/GCEL4BBAso4LfggoOWcNaf8hQ/KTRJyjBUdcvx757Qy4JYLao0eEG
CoZucgYV5ZNNOzMt6eHhq9es6HkTzpUW/SI1d0M1pcFjoivZqP7o8w6i6MBk
Zex0DLPgrSu3bmsUwe4th9N/KT1SEebMrdda+yzVyWq7R8WLo9FmPfcMAher
iAMsuZvw2eld7AK1AZ+HLNl9B2xgTScwPKGCf9XE3DWqywcC6lhylrI1TKEJ
XesopkFrhN2CVCvxJWbVk4Ntv6Ifd4MI+qjRdqII103YQNPpEyfH6sCQ8dhp
7Q5jTqJVeHW9fMBXdf9qZnozbJgMLOtwN3U9Pdih/t9PJonRvUmdBRoTGrY9
5grtbHO9JTcufgWr2vWlFB8AAdkwzrh7avDdbaYRaN3Z+mvZKCrBrHYLY4EH
V46VAZWQX6M+PK/8NxGeZ53jGk7U9/SWJ+Dl6n2eD4/ipQD3E3Zd9no5fSxy
sLPDpw1fWjAzXhpEoT3yVCjlvin5bOp+2Fi3WqUmojiZEEvEqPaG2aY1/m4y
fbiwt9dQH7iRltp4v9ksYOKhuKxfWSAVMIwkwSW7ZxRDH7unoGKmmX1ut8Oq
twxvASubWftK31NJ9S1ZRnNGZ5H+Y8ocLMjweaWT3seGbj+Eym4ikmvZndsJ
HTAWvbUXVCokrgbEq6kbZDrTTfAMVEl00WtPB4gLDvNMiX3n5di9bL3hFBmp
EXUERie8C1wPbSdwUCpO31uxIvKgH9qe5OVplyhFyRbgiPaB10lPGs/b2wZ4
lE3jY/DJE54qNrMH5q3DN5W4k4YoXIZEWJuY5gHhPvIvm1c6IXUw0z46gG94
A4EbQGunMpnVsLEDv9HP6JDgRiW3JIovRdRjK74N5iSCZ7cGEOtJRToayLVv
OVEKUZJ6MnBEVKB5w6DY0FkTvSNBGsxqdFQ7bVCkkI/7blgVNoKYpq08b03y
G0KuqKoS/T6ESBFeIXqxVBJRD2m4E/brLDXfxZzruELQKhHR/AAaK5SEEz1+
JSVCRygmB9aui/MPBnaDsQ2Ye+cm2iuxswSMH6S0N5SJozRYLp+vz4sd3MPS
KqSZDoAsifx385fyBAxVg7k30fo1Cl78jD3iFT3XHIi5Sofz3dutajT9VVmm
1YMkgp8iavNv82gEr2d4EqdwT7SCHaGS/aqmrCxvGo2VJhHPWUhd8AsgW6Qp
gPfSDR64cgFeTohaTU/mXiFbfxZbbLxN3GTIREEL8jHaQa1gruU91cvNpYo7
YfOcnCBOqUVYsFmH/QZU/DmrAA+9nfRDouI2Ks2lntMY0eDEGP3WN8UWhE+G
XXp6NJspO/eKnjfxa5iXoH8+8QiuQY44emWcZJJxnXQrGK/ho3QX0ht6t/gc
dF/A9kTp2mzUGc5teZlv3y+zjJmbpNS/GKh8bc4V/8Ct1ym5pxwCze+kz+rA
zTdZiFZEG5tWwzMQ5Y4Ptb4zbUkvygez2n90Mk5ojsxYeG1XK8Qem0K+rK83
iLVERvkn7+cWliHG7iOszqRQfE4GJkRIXYI2VkrKkfaNxWrmHZMNha0XAIbk
E5JQBXNxhH4t2iax6a7P0S6C+cD7GphERRgPGMLUwGx/4aMfSY6YBDz4Zsnv
jgOQVIqkaWKXdNgUX1Hw3WQOohlI4T59cyLGDzjxYcNYpSRY78TxS1v6VHrs
bVCSon1+73A0cWjKc4/epf0GuZjAGZ9+Wee0dNvIDJTzujKGCnr82kIXZ5FB
cxzExOdxR50UhHeNtePY7r6GcZnYop4cO/HiIO/xm2XGrnkxSaECiCwK4fhn
D9K1m2ZWpBVP/ESELkGRA/bAw6DxjyU9HPGCC7iS773AAAINmuuEdD+L1Z6M
PpupOY7ON9U+4X3fKV/1aXElGJbpTljM9l8fAcm9R8fyKGwCpEF8xsKTgsiA
qReMZeMeLCI5f/hN2khnOw2miXv+qMOTdobt6xrT3VXCp2t402Jy0FSrxPVb
iLhKIyDx/WQCsDKc5zGg8d1HaF9i5/3QYA3uUqNd3LOmRfQI1EI4MJaYIqJQ
3kSCsL7eZWtRXggLP14+vZyVwD19NWfyE8whw9JaordvYZF36svHnxksYhzW
tfr9p0x9LWjdRV2XOV+VIE4FUcc/5EEkuo0UOdJMiahB2tYdB4APfVl88hDu
MGgqRUS5RtqfLQDYRd+oa7SNbWMw7U5565XJmP8fyLoqn5PZ+8fpyNZJN+AV
jpIA6CeihPe7Q20p64W32eMfJ8PfiU/3dz6trIrL3MKVwa9MxLIRA7hmaQDw
O0Ja8hGqsQmgD5dKHvhUs4UrNbRWD42OLqw4GEg8pxmQTiVsWqeMKplPDKGh
RR35YWU94ULmhCesbQvUzIF/zmfwnfDeXQeY63OEewyO9945pNOMgfPq6yx0
XMxuJLt0yJiu/pjkM3IJZKmh10pVQHbXyt1CF5O8BfcVgETyiPYaoWa2LY+s
FyBKUwh/VDtDV+zVyvl+u4xc7gSWICOEjEmCOCtSOoNSzV2alMdOb9IjSbN1
6hIFMA7PE6CBUSqjy7qoDTy82C3OqKqoI4mDh73gp1YLndxbAGb7YgcQkLQ0
YXiUhpMVbfKKlFX5tgtfyPTdwGOpb5Vszgt5qxzHWBP33q1b9OLTWutVEuzV
6WTguhMCkYeMMNySTM7rSc0xJoiISIFEp7U514i57a8/3sbpf8GJQAenYK7I
CznhN3RD5Feok0KM+oVVMlCy2+zVaAjEoeQZBOZqdFZskW8R/TO41FI7GXpU
Y0NN4LWa8STMWuVDTRLA1CrpTGI+P0a222wIX8Y5xybXSL68hSUR1VztIxvP
/lWJ6tvsoTCLoDRDQXqO85yXczE5dKeWcHWxSUX8TFbdEXQVG28TCrtHYh07
IhuONkZmLeoUYesU+l6ukGOg1JAc1bTBh4BNaxQA59xdkUsLKi+XovNLN1Qh
yXJTWjNuUfemNCXWj8CGLFLXjWKKiN1YUl0j+t6aX/PGq7Zx8FVQEa02R8e7
nM1TR+jW1KIuOIEOY44TUHfWw0TfIwfXCZgI4kJsKloEWMEV1Rl+WaHXjVCL
cEYyfLYh3rEIYon8D500HaSEzdLLwG/4eQK67k9E7+1Z0ZSlppGJc+/Q+pea
zdcbe8iVWNf5v4nZNNBF7qKjjtDXtENJsGblBM0nFFm6qZO69cMXbOv92aJe
JjedfrqyTwfCTzxRRtwA173y07OVaNDqhzNr9rsxHQWNT8NUZmXJU560iRrt
1ft/pHRr6MjrpWMx0ssKh7SNOR08eTFijmAuAHSCSwzkLKd6HTzymap5oJoy
tYWVrhhn3nBrFqznZWojrnRMKCEvlyNlagZJB0UODDqhdCmtoJ5RklxclCCg
kO8ZVrVdRiWvJReJtBuv3dgOvCoZ65DgEODooM6ED5Y7vC8uG4p/AI0ElOFo
jDy5K/Y/ooUzUKEPhiOAs0xGH2M7Tm+RG7DiA++Rqv++12c0BITDO0YVNki/
PJUO3P9K8ygxG9SXP+/soeLK7fT4rkIKmgOoofIMI+z4FyRFMCP3GuwxRvEe
l97LNn5tXvGqBoMnlcrUc+kMKoDOJ9VbiaKeNFb2Ch2PMmbC3FyjaHOEwKNi
fAo8diRQCZL4v4cgRsVwqHGPOnQ3WroSqKWObUAiGLmuY5ExjUOhVVmS+Nrc
bhpbrB8E71iibhU8XdtSa1/R6eD9riWIANj8fCIMk50o6HHlo6v7vXMBsLtZ
+xoTtj2LYvRSMyPMYv9j2fNkPZpEGlSDJusgBDQhh4L/e0oxqcl8UDxBp0Tf
P9bpn6zuWDJPjHRzGmRQquPo2KtroOKCRIuSA9+Eeb8whB6bYr/4YcpY4i+7
XPmzCGlyN8aYch6Ubw2t+jXpevuOhIZppCfChKl6KIDQNQ0Pp5TTKgbedCBh
5VGs2WeOTmIy4+3iyfHi3mv51fK7YlVrbnYQCFTFB/eFHGyOhe62R++ksMYH
fNwh/Zx3GVJF2kDsnWMj3NrE+uRMKYT1dmmWW64gmEjfrvJZcSbey1rbnWKx
tCHVf16PqB1oZj+x8VYJIqHSwcgIhSATKPa6QCkPMBlOGIWvwPCgq9WWHyQh
pxqcWSuRiigDcWFnoSPO4EqdNoe9vcG5szVtzuXMdeK3MMScETu+jODxmWoN
rKYpwPKaLUA5l+SLprsxr9fglkvWh/qkZmZoPO58WewbUpnHlDxdTWosfC9I
2/mDFuytcYcdGUat2Y/P7Ofj2aQ7Z4fQIRsZIjUUj8GyPDquEoyW/V4M1VEK
qml62N0v1lSpGIRI46QXhE3evzq8Yq9GU68yAwEqhRw3eiQt9cnVDoO2dWLC
u2wEUyU6S9kpbQZDUHELpE4f03sMSAlIII/2TxGo4hcAl5pNTy2ouv3ulX1t
4TQ2/IU1xTWyfniokuYU/9enXusPIAiSNilpW1nzDwaof5efEUot4Vss1BWd
wWbme+ezSzBFFe32mcQccesKT3QQY3vd4y4zS6A1/63Lq0sVSnZe5/FSRaYi
7Pxx9/SWPabv3ZM0I/y6cBT7GftPnhvU0nj+6D1x0mnEWcdICO53Yk98Luwd
ehkmsGlIPDkR84kPUnztx+wYff7YRZ/PpxLe/aXnw2qQm0esjvtdOO4+q/Vj
Vhu6LWzkLYEfCbiEgEo3TMa7NzzxxiEp8VJBPfnWGHpWNJvu+PCygI4Y0Gk2
nkSdjQlmturQKbRcyHFO8OuPxovHxhiD3esjdghFCOu9c0y9gUwPjQTjX0m+
XrRcrPwNzWSjmNfYbReocgzeQgNSvTqa+DqfmKw3Hx3L3ETES2P98sU/oCCy
1z9qzD6xwle32ZXImQGH4G2HqT7utbSqTX1LUlEVFATrsRYaMpB3ZtveN3vd
/kcmzBwfuxQdjHkhnbjD4cJ2A2gbMPqiv9ithSr7K7Cd1s43DX/H2LKpA4m+
ITOFT0z44ne3jLvO21bV9ji/XW87D9qalEguao2dwg00Fee8SFWG4m4llojY
tGtbWVBOEcWCwn7nZ6ltmitdNSQy01JPBMy4henH6SwtrLIBB7Z9mVGr//7X
FRhJGxEGsxdjjcm07BMKnm+j6ZMVjz3wIZSgZKlWoX5wKiKmxLd62WmnASwD
xlv9JaqesoDdj3qL9jjnzXQ17CEF5aIdREBw+BGFWtFPmrWZ1vmvWlpmRb1i
qqoc1NSgh52lQrdKmk8oAu8iGitk7Q+/ZGAf7r+SKfKlrv2DREfo3o599xwo
GzqHcICK6VcFOwOXf9FhoufQeK62r5y4TBXkHFxKwoiA/MD4JDUeM88UlYGR
gA+g2gWhEMRiDSaC5ZA8dpmSo1nxS9o30GcJIeFK4MiG1I/cUafwqvYS1Mtj
02XqmTeZmsnijie59bVJbhtVvf/7rfC8/71F2yQAfX8YmZ7X6tNuXsizRw0d
pJ24pEL+08WH6a8f/EshJ3DS3QHiAPFt8zGvWleXvbGwpqo8+skzKkRbVxTA
u5+7k+XOpOYf7LVD24skg//yHmTrnttpfBeJIBzyWA/NFzENMRD85pgHA57S
CEZkIdUyL6TEKLRU9xdAkRRFeSZXrwIuNnK/XQ7o+2TJxDcQvYZS++d5pdWS
7RqNMkm26lNuZ3QaSGbDbsFuwWM7705q9XoHG5jvSsXURX9TihDWk/Xf9CT4
hP60T2p7UfaEMD3g5aigSAQcoOI2sIuRdTMxhg6Jp4iChP63Ux/I1GZj4iUZ
b+rvFBeygLYT6Em3k9V3GQ0LdPWd+iYv3FrqQQGFRcZz7gjOnPHSt22sDy1J
9VhcmNISreZmRnRYUXWsUfGMjN5cFMBj55WrQpqY5vgHIw/IbXFL4AbEOH8a
AUsDdw3XH5o4ORtEs/PcDG4UspFZwA/IgYvV5glA8MDLwIMHR86nPbgP5r3k
4Weq/sJPZlk9Q4nAyHpl4464vscRLz2l6mucQLierG2xsDDeG4v8DVeN0ZyM
H3CtJ5o8Y5JR02PT1CXBLUb18wGagC/KdK4XbhR0uKi5y9KUffbSrAR7q4Kb
BacXeNF8/56Y4pDIDHhWbQ+oWeghgkJcXjP+/HnLkgR4k8fF9nkW5Tx7npls
Fsn6bHjAQMZjBxi/cvIBKAt7RUyoIqcNjH27fC0RG/oMAZQ5sECiXTDWKljj
hG7ZmU+RYifEQq61WnpldFJkMcQv5cfJ8SBlfteXTE1hrVILWwoi9VDChyjs
bzC+EPQEHW8ZFaQsWCYTlvXiemO+QGqURRSFpN54SbVuhYhP1Q7GNfF+zix/
sYY73ge8l4CjQCHnQ+wjl+5Ap8BEMZ10FDH2IrcMzjK+hnKGv9yWV62DFdcf
W5xmAYwB9qvrBJQZP+TiCSK81Dx/Jq8K/JmFec93/jBeBDBGRQR40W27pvg1
tqlXGK+Rq6wrs6E3S645/IeXiUEWM3AuFXspp6uHwAgiW+j6ossdwAkecrtM
pPdKCbSlS6FxEBA92g0rzRbsPkVM0gJtuq6MKchp52It71Bhs2uxLxfYDiEh
NtnBlaXtANyWknwNyOH7GCXR5T0tERjXVaExZU7M5/e5nAYqLoBnROAAc7ZA
L0PnbyNgGWSgV3kC+qG48bYU0LdWRciIIi1u3nJH1/Hti1PSuyuw+dD0wyw5
eeyyF6nDbPBST3hL5cuAP0NM6Dywkj3dRWw566KTk7S/qiIf2lW1orvdJ8re
jFQLYXAjAYcZ0A2FgzwAuTHv2Em/ySrkW1Jgk2W3jJTWp2F3BUmrgmv8bQvq
dfr00S0NbFo6BpCI2WLgB5KNBItOwh/MV1qHqe+byoxe9dAug0rCRckKf8UF
JACvIgW4ZzWIor5+I8X0kILRC+Tb+3JaVemxlqvYfxrkw1zA19Y7RK+AmlML
bmj5GiRHmHazA2cNMWOy5bSxZgdF3b7fnPYFLzxM0n98ehOknDPQBixkA4uR
DW7dPlqxBo4Kn4OY2Ou3QfRuZacGz1T5G0ckPLWJqN3YdCSYzfhyC2xBvPZK
W02NN3EN+VaOJ+F4/Yg0JNQA6KJorjrKx9E+jxH+uUqWqHJqLb4Ssl2nYzq4
9gM22yHVkkgx3m7HrMBlXT7DR48xs60+L51Y8TYCjRGnM7hb4EUdrFUy8RTf
g4bp7dW/YG7Mlp7NCPp7dd7Q+CkcgzhvkkRQrzBO2Ccy0yFRbFtP/jZSfsgB
rFupldNmSOo9FI6a3QYtKG8FXfAKzp7lyEZDFIjpctwaQ7McH6elWyL8PQVa
VQg+omNiFOVYnHlK7sFHA70uMaOyEBZdY8UHfSOoIoQbJyzig/padM8FRDB1
aowMfqpPjvJwG//VJrKLh6LEeCcMjt0ASS0tE0ikWPj9B4ovsfDmb0xdL/8E
0cw6V7aki2h+IhL56VMi+kC7i5ZFy5myTqN0d1Jh0yv5l9cPK9vRBowsCMY+
AlvDq+Lz4q8NeFzjJWtOOMMGSIsX0sQLt8jFhwpbXSDocFayObyKHLKAv4jc
x6399rNBuzIm5VItnozs2Ee9V/b+2sXlQoHI0lC4uVJhBAhP3wyepRYOrFkM
scjsjCj2gwqmPHbTNEyoJi2qfKuSCFwOSiE4Wc2zcPDV0TnjgJEoOhorjhxX
GmCHBU40jyeZFUpTXgn2IJ1JQSLMieqJH4RGV5Q4t90ypWTczCf3DWTTF6nm
ezzOk++yUj9yai1k2YZCWRoYHrsulgsTzZ7judpacGK+8aPsQmF5lfow9u03
/UhqVFkjHeMyDahboHK+wXHYkDbrHp2vvlq5FINa1LaobhxcPVmmPvQMQhqx
KUcuVuuL/cUbQIaxpXP8Kkz5zL976nQy+YU7b+wZLvbr6Oj2vf0WLk9tmDRb
CUb4dabeTOfhEtj+c0DVlGZtHH9fKU7JKzfC3/oSHgeiO/5F+ZHFXaTKiFDo
z7U8AhaiCGchSIt2Bwu9u0aN1EXexijiwWctRC5JsvEx2YKaw0vN7JyCIxyu
Z8clImeWWsaX20WNcMMKFI8IrACNARjLjrj6JYj/PetK/Z8HUMwa4/+XCHjg
CfNSRnMfc2H+ybzS5rUvdUWSrfNnH20KgcQCJ0+MNzdtDesUxCKAjFtfTOoJ
eXu+PMPfqCAOQPITqyrc2Tv3UzjWhEgGN41Ee1bD9lTOugM1Hi84KTWmZq5T
GXUromKEpH5GYgDaN/qhLcH2BS0q+FZ03iw013Bwd8gfbwOM5Sc25PU6nm/L
cPZ6iXPVXyyIq3Ol3nRgnMT6iEl90wPlNzfYkiHS6nMTn1WIdfh5s/hIyV+x
btOe1GwijrP5LKK7m+j3FIiZN4evv7Sb5JuxBLIBJlW0XBm5/3xbyDHUDerS
sBIaGMvcXmIgJsFLFkJikC962sbMjwK+VgaQMj2ESIqVPOhXwJ4RPdM/M6+F
o+xe2ijFSPnszBc0mCeCldwtpbzPOFs4rLlI0DvCReO1m6JgPpjYlSwHVhzB
P7INhx7X6buDDV72tbeSGLHk125wKsVUr8W8McJecyGZPKO0zhWUOpV5LvRY
t7XJ0epepxUASIXREieeKA34gFFLLrZ9XNyGcZu1u8ZJBhjVV3GYOgN7+08w
roINBBGoytBjZVnJmK8GjLLLV9D09P94y7AIIOTOwmEu7uk+bLU76ZM//MpI
JsBmPmBLuyutd5QiZF6O4wwlPbPnwPWQDTmz+ORVEQYTsy4gJ1cKIxjkbaK4
3I3gfwBm62/LvgVgjd7QVEhWJRU0BnJOIyW4ZAkcXkSueNkJZr8N7IDGh0OH
h1PJzKXPoAsVkEaBT0iy+Hqx+okvaY9FtcQBIG3o1lIsZP1lJCVA3lCCj/J0
VKeReh4P7dG8TiqOiqfb8Flp0tF+zKfbUQt8zGlGown7sRRCl9y41NOyIQdl
29bPFi5D3qXKlHit1gegZUde54oPQxuUF9Lk/DwwTEKuwo+40iJeL3Y1dQu1
g9VlD+qoEpvrQN8WhfFHeyjt7iWjIhUSx85Vvf3MRE7/tRSDshYCn4bFJyQy
UxQql+BZqFRHGmUAy6gVhQ5YMiyFwC+wArsiSYGipox2QQwbZi0/Ypdd11ZF
8ZvfalQ/vU+njp/BjKXHvJ19hGjgPu0sbfOmH/K/LrOT2fWakTmzAemTqYgT
IprwTU9OkiQoxvoL1x7VcczGO56oCZLNads4v/384UF+zX67br5rIbB68GNS
5kyPXAD+rTH3MzLb3UmuF5pz4M52VHX0AE8t0sRHRAArhSLl+rEmNb7i0yt9
v0m7JUmJwuEJ3vQ32C8aJvdAUMtdgVDfiqTPo6oKiEkr5RdHIkTY+zuxSDG4
tTqASNiy31ad7Vb7r8yapbFm66ZteqiQhPkgxG3b+BuGRvHiZW6tLYljwpQw
EM8UIEF6cmC7ruSWFxj38SZ3eD1f48aYRbHJlVvptzjrQQUl1PziElO96LzS
FH/Fb2bKx4Ij6RsxAVm8NMDFfGI4D66vC+uhMrJW14vGLb8lDJHhq5f/Vnmh
x1DUrgVy3TubGxmbcrgnfQClIMwSb5SCkPpHv8QNkLnUArkT78Zg3+7N4Zt5
a34N5UYDmdryNhoOiWqAJMsyF1k2AkWEHy5i9otcFZHUZreo/Jsjh+XWhExR
qVdjuhbdSR90gdbdOLBvuXGbptMuP6nqKeINxbmD36/icU4UW8hZrGFX3pDh
RVhtIMWYibpfILC6WqgZq2ksc2PjXvBaUOvk5CZvii5nBHtkAbeNQx37wGE4
lD/9Y9tyWRWEIHvj1mHXtNNKOCMt9/rVZ9WxU+1ZIILGcYXaq05Ot58o47Tj
4LzyYDYbHcXLEFbmtAJUmYJyKNCgBlfFIKbj/Mg0nh2QaQTen41R3KZVmB4k
eoClM5z8fzo8Ph+hFoB42YWWYtMPvw7ewuCYKOFmN9nwRq/1szrOnxTfonrG
RGzVvbdSgD3JWOj7X18+Bae1L3GjMj++jvR4MljUi8TCUnS8tSOPh22hEdTD
bPh626KQTGeO20io939FYHHyz66JdQTmdWZ4imz1JUWQKZxEX5jeHwJbRdkK
ix2ThFmvemy4HPYva6itEXJPPbZrvDb9UsaCvT7rR4gWjCKCaCl+9OIA1p6S
zz0zV+wH/9Zpi37OfHAdMYsY2aob5r8x1fB8XzIoQvH3rfLvJbRtyxHHFxqI
JxvpFZg+XbmPEvK5UIEWumyU0S3Qeuyo5SiMEvYwH577a1DBKsrlfJIL/lsv
iXmiAr4/c3kCFT1kRCRPmHa1/Tap2MJAVUqp0eaGtLpB4P3HJ0Xi5TQHrhDl
YhLvGvPFS6Km7/hMJoCcsL/OVMIlGsu4PSVRAaLF0rHksWVMuuDLtMRyY/YK
K8kbV/NevhI/sih70JoshL1WQ5Pc0baTZHLIg7ERgU+5K8gmh9DiMQ8RzFTz
YSNYkBSEjL9S8py3Uk/0kWInk+WqW4UjkIiVekI7RNkNigT6XfDN64OYKzuN
+TqOlCv5Aolgk3Fshw3dCzRbVQcwRaAxkeoiEJNQgnBScSb+dw+cHl4v2B3F
OO8b9vwSmEwPg1cph1bMlKP30zc5hW9b2hKJnioNjdpP3PUaTywDDqhuMCbH
8QZsW3n63WnadtvuHXFk2Zm8K108kHOSyVhMD2P7MONibMUjCCGWQTzITUTm
D7I26NuQ1EpCOinsVqQSI7LQWp+NMELavxDxMO587YntQLPT/AWHuqaJ5sTk
NW5nGMaepiGk+pRtUmtff+w+hgMxp0bxUeymWsxdFtrvX6hjEmPv1jF5NJd9
x6J5WPw/CqeWl/7FvRyhpjbZnx91iNTR1Lj6S49e3r/Vpi5KGl+XjBSxahky
KFsJsABRqmNTdvsf5nKrXOJWmqMowjmra9bryHO9Avt6Eahq90jStP+jSDiV
U+wshuQpDk1YENqM1iQ4Cnbrad4wksVzy1XX3gKi/5Y0FiaSEBlfvjKZ5KSR
wOP8N6yr21BgsB5Pmk1gYKr8I3mkPXHlk0R1m/4Typny1XpDXzxpX6jcP3Fr
/UUbjjgNnC8WsWVdzzY7UAvwgIUbY3uLHtGFZnoHNIgYoVpEPG7sfLaBE+RO
yw6nvoC9GtFWYjV+jnrUTpqFB9fyMxSR77Zo20ei9xupEqfWE4t+GfkDjwwa
Tcg+DP1fKHNRH3jF5HxHxCDxi/94Kho0UIBMxUvdiBjuwgnR9wjNjg9GLhY3
YVcIms/4Ud4iQT4tPDhW6kXMimID24sbtKFZGtKeUXU6DaRn/n42F1zNcKHC
sReXh5KrFJKRO4tHgIjHwh+d3HapxjB8Etz/QvWmQoyT0k21zF8S4AQ1QMUh
EyfICiUbSO3c3h9aPP4IZGxU9ZEXO0wPvGpBGw46IdSvWLXJEYEGdxh+9p+e
Hfc3kLg0MTrydoA8VUQLteJ9cJvwkdiaPWoCPfOvI6D4qlzl/Qo10d01NwLN
njQlJ6Q5Al/LjIyHACiDC2X8qsP3mEd89Aywqaa+/bJv3RTSVesLaTcZ6Mxa
AESnc4k2pOPnJCo5wsZSF18YzutTwRlMVmJ6d6opt/aJuJyJdU++hnAtg7pv
REyy1/MFf0/jxcxD+hU7OydIYA3kztTZkkRIlNxa2nek4/FvcxnMt0GHZSWT
GaIMIhTXBbPXVqTqe2sMwpced5sucJLV1Jzc1kD2eRskVp9uUBw3mojGblkl
g+PI1yCWruF0QgbX2/yvk3CKvatuy0cjIYgygfXLxXTVsoYl2zGZDaOHWXWC
NDuCkr5KRm5hVNMvzi2FuDd7Qwi2JXRgPWH3n1n+rZgGAlIj5i0ud83STN0Z
yBuhWIe5gHLX+RjxtE2Sg8X2GUby2gP8w4RKK1xovqCsZE/or4J5vGK8YD9a
LIPdg6HYogyBcfjD3SBoqVU0yWORrUxV3s7rNoK+Vu4E7v0XWi4tiTWwAzrj
hhMHxMU4zx8isXJpKiJiv9Qt8HNzPiBO9V+iK5JeE5I5RImpS6MTSzF2v7uz
sKKW92Hfb24aYpv0VJgGnJ6q3dXOewqGTHTbQbd3O/G+yUjE5UUhsPSqDpXT
pLLpUZ6SOvDhCFppwvTOHQuUL+AX8pW8oSXu9FU6hWgLxiGDla0f1DsaktBE
0LhpgG7Iav680h8idkb8GHfWfx+/MEDksLojoW18L7PFxvyXyH9Sir2fflCx
ZM0wO6DdHyGyYmYb+8NVq65nP2K8+d8r2BzVq1YUfMQw4G3/fcdVWW0oB2qY
TC6q89J/Q2OMrZQhj7wgPB39e6lkWy0uaeXGSwZHv7H676gM9TMTCzG1Olc9
GkgXMvBd8v83CladYL5l5SaxLPzk55DDFZ99ZDxYkjtttHH3/xgt6x7TG3Ur
pIlvHtubOzgmcYmvsWj0vLR8633jLdTSLYFAZQX2iNP8EaXjZz99dBFid4mp
1vvva5wAhkimt/48kfYCawQZaUM37wekZUSRsoCrOAaQ9BSdGM9D8RlnPTaT
yr0IRiGGqDCm9yVeb3Vlq9EAXLMDMQRTyyhOuO6va8LYvYz/cT6XzZhjlL1w
pPLfPXPo5toeeiImecRNFEx6X4XN9N2kCwph7vLZnZHNbWhknPTdzUkXKMUU
d891zjybves7dUNRjoSqfP7++0+ZPJzwI2FBzzk+AM+Qt7xX8ggw3TGrakcK
tY28WFy+pgfbwSvLNneJtR4wn5PT3m0naYP+450AT6ewmJlfcCQsLeywL/M4
427jph5/yirVKJxXc8kNfQkwNa6hR7qqOLJNGKoQQlf6fsg7Vv8D3kDPYsyo
N7VL9I3opgGSVfei/h6Ar/RWSRctSitY9u+vy6btrfxKS7jFyT2AjaO7MRXp
ysswkilUbZ3u4a8aEjzZ/5ZC2N4ytuOUVjAu9Jqyf6NP79LnhbscKJ1ZBLzI
qf4bLxNtumhHJKlOtvwfJMT6thNL7joUJoo/8RBapQTWuQkdJ8aITifZq6nK
HCb457zGmJfpHNNb+Hi54NGSJFX3rBnyu3nJfCn8K1vz2XSvu5v1n8u7k8AD
vjO2qFCMVyHHbPFSmYqDnRAPeu0t9BvM6HseR2MAweOS+Qbmq/GhvP9pO1n7
o2NCyeBn5+SobmVUQ6skmp7NFABbfKJraWvoFbD8lbgXI9irYAQ0RKPF3ao5
xhS8QpWh7UkPMymUbx3K04MgBefkjw7YZbiQT45bb9C8w/eCxhsdgdN2dPCY
saj1Jqx45eDEqlhv01oo5nOS6G6eqEl7PsbeuFZNCfFNJ2PBAgG8uiYK3KgR
9HnKNiZFY8HcaRVMb12iUtD261zZcd/IaHXN5B63YgixDc8pRUSyLkB0maX6
CbumZ2/HiJPDmfPNgHlDk8ou2IxWjxJwGtvOy99D3eRCYJBWNCBsE/2UE4ym
FlJozyOByR1J7h/zzhCoEG4QsLRKZQjsxPTPywEeG6NKxlLdDM29Ve5vN72J
MZz63++nhAEBzdcsjQ0jj/vtL7cLNXHa0nPYq+AqY22CcgkcXdM4CU6EuuhT
Vvy7CbaZYjLMgwj86jF0KspyBCWU7c5LwixjcY0aoQHzVTplOHSYWe8uewGL
FYyfdqsQKTGM2b7URvJuH438ZIwDY8SNO4gHxmrTmeiorXwoPvQcC7I6FXqz
ysdYt1u8PXnXSuiGmj5TSDZsbFjIyeWEtQneMZD1FufHtI6bXB+5/d6jZ2BV
nLeWRSnDtDEgGUrruWcgStrFTin6yVa+WwKKrVn5R1n3IRaA8twCYWoU2lSF
5zuYI9o1+UB9ar+O1lG6W0zvC7gPdBfrAtvXp6kq+hXyJgstp5CJXUcLHDJL
EG5qKethP5M41g1ZlOY3MLJLTnCH8U3DKIJniz8nzYHx9J3BnA31D1eT8n3u
seG3GEEoPhD59CR/qcWezoFE2Th+cAT1m7Bo124GX6mPlkb0XTYg3cGgbbmR
l2bdByV0bO9PyOcjxsubqEb7656PsHBZ7sSUtHodhUmiqZPDn4Qhr2SyEKYw
EmyDhW5yEhReRneCCnMBh/77rGXSy/u7bF2UYfVv/Uf/lnD0GHLrlfKT/Qud
gpkziyELrzsZUHBhBk5SyBqVk5c4K2Ry+zv+S3fVJMeRndFVEgGyj1SQInSB
6D9XSmGPwmXQlSM+ppYetwVI3585yXuRQPFROfkUYjD/hq0pgLLz2YxOR1m7
ic/wdkvCrD/Vgokfg8d20EpC3pUxSshDi0fSeSBhnNCNaYaI+iasrC7G6EAR
f0UydbdAbU08YMWKryHfsB1GSjLT8da0RgRa3PiNdvQf7ldnSd2EtGXe+uEg
IAuoKqWPLaNvJy/MTJCn2yxT0v+KvznQB3xfychk0g2+wan2Vpc+31z4xctB
p4J0gdkD0WlLujuatZd33Ra30NK7/TxodUj0YJOZcSZngwZeCk39shIZUw3S
TeP3Q0PKcxNWOGFxZzHmKtvNWweICbreV+yFnZmwffvRyiLiuS4MLr+vWIP/
0hLCxviXt1nyJvlq/v+AkrXvycTes/53ph58eBh7Y/IJkFY1pFEb0RO559HU
H8Q8h7eeUpDJeKLAhDkPFENr2dUW5BVMX/Q3OHWGitVlLgatWxOtMAoo2L3N
0XFR6V3RE9J2cuGRXvuDiOfy6NwzB9ycbIneArlFP/ViPeO+bC/wBO4NdpDy
dhE2WiuRhq76UEZkzjV301ULGhgXupTrNmny8tD75UH1YJaPKgUZVlc5h/XX
ADa3z5wXl2PAgMgQgLvRIlcxL+WwqkjXSAQ6wmPf4nb9q1cGlg7jOo0smHi7
JZSM++UrwAAkKLVPpI4+Y4Nl+IVjZCPZlEHX7ugu1oulLFiSYAZqqilTWUgQ
3z0iiDxMEupn262SU5Kgd/vNk5gzIHOu1QxV+83Fb2v7UAuUtHncO1nI7DHU
T92EjoZL0noKhqsT8EdBwGyNK6ROl02Y1IbF1mMO4O4GlxxIrW+NUckoBNGY
WNx/tD0AYjJeydQ/tAzlI0TLVXKJtqZaqc5+uKk2fYJez7Y6y0/JbRNZf9ku
zgNhkfCcQSRb/ajo0FKpEb7uyjix4ZqPBkXE9aEPnjwTu30b8YqW6qpM0IiW
iJvhHB4NboKa/R/RR/vLYSGSZ3+XK51+RAgOo8RBNOEYjtJH7fTeqmijOTpp
k7VggAjpksMWzM0Dy/qZpFNLfDhgVwPebp2XdjOvt0S35+Fvp/3MudGhwFyQ
dTAwpeY32DZdn42d29JKn/aC1uQblnZKTsgst51yy2HdX50kMj4jWXNGPW87
Bir3TqNIGlqqL2ERnFvcDHGQfsl3pDMbg10jCPm7IxH3LtKGcVhc3b9j1ViJ
IAHGn2dP2eZO907qVPcGNxs4kPvMFCKDWtoimScNiV1QLIVwpM+XTInN8BKt
3eAsAiS/nzFhLWB19GqZqA1HX74X1DgPlfGekUXAs6EysaJ/KwHh+eLExn/7
76FrVDzmLAn6k9xX4khjbQHoaOdvCfVMYG0N71RuuZSkm9uo1Wh+wHFXDDVy
dDXDvM5WROQIcn+KB7u9q6ZQxMAH44fB/26DmVcYP49TwcV/tBZp1vobI6pk
9QMgedFhtVAKm0VkieZHSG0gOB5i1I4TbVEQyoZzWJAPYf1S2YsRG1jdq4Nv
DYjwPXg3M+UPOKIMMBy3GmNu68wN+GBxmA61+bTbkY0uQLzRy207L8ZEZjlQ
68B6+KLq0CooCm1HbOoabnvCit5AL1KsaM7ves2ADFBReYvD1TZStjGW3xew
1XIHXMcA/xVDgtNAKOy1GCC50TkiTneSA8Wj1eUBGIKakTxjGCXBBu6MDqSO
1mzDnRkRDFT+mokfqtUtmmWm6KLIK1LGF7lDJA6QlE5+Y+UYWM1i9917NmM+
hvwIrjEVWujYdNv6fXLhnd/yDCFa64pIZjSSx0bbKZt8zlSQCPSuC9+JJ6F8
CxtTdJ7SQZqOmwR9wthD8fwtn5lw2DrHi9wPoLGuiGixAFq6h7xKpZjh4hff
jwCJ9/2kFD5ipb+OWiZBKX5P3PIxOFs0gAseQtGTSI+Q/vltc1Hj1TXQ+03X
q0FGyayXdBbbYcSrBBt4zfZQ7XQeo2DDgZOCm05/fcWlKfyLIroSIpOcfH97
ja3sLeo2rsNw7ck1iqdhGHkgq9P8dTK+FIfUjnoreIW8KtR4HNWNv3UCv8bH
zvt/gpSSjgFRJOIK5Qet+LXO8DN9WIXJUg7ejoVA8Y5Nnf/8eP5pSl1DMjsQ
rwQ2jlvLTHecp+t0fxCIF+/5cPdHpa63Dt5lvn6jKNCddZYYeZEgcZGc7kwq
pIBkVZhnrdu3L6kTOBROQSC0AI711sASi8cgamuAVhdQEMYwZ+snTn4L5S4D
mV0+P+1RnFnZ0jpMwDxMxKk2uv0SbWdox9j2DjdWex24ZPPE4mPKTD1tvZmI
3HekOBrWgJkQmvtNhDiYa0lqoZshlnXd3yZz354WXMsDIAUItRw5VI00GFPI
0lCT2zUPcQMWp/Kyq3dfPXVGqm8ywUxlWhkr8BJ1ihNwHrW9IgI/MEmEBhb/
96zk5/j1C9ijIcjLB0mCr27vPlodSb4jM/XDhUe80Z4NfV50B0GN14QYTL/2
PzdKwkdLLIhiOvQcigk/RofYt3Oe3ixeFjjUEGRM2+u1ZTBlI1zFs7UV1uz6
y041ZPUCmIQlv26xVomNDc0KEWd3/uD1VP3vqkBJRUCxVSpz8DMxvoJgwET9
fgU1uCrbxGsmM6iX/qoEs7/ndTJK49snU/Gy6MWUvE8z/AFkhNrzLTR9bPXw
wKT+ySsnatgCIQK0AInmsAujXc/c7ShCeYeqTwHI4KYvB/aBB1SLnXRh/mMg
JQQzgd2pqVkLVQwtXFXijhGMt5NbG3HkAHGwKNno/SFXMBYeLDaVXUeLmDnR
X1ZINwuN8WkUZOkLiou3VyBaOAy9zZx0vCWokTMx/BUgBlk3lM0zgCjDN9Xl
rmNwJ0AdUsp43bREADNIRWzCuI+GGTHFKTBmrW/geMCjbefpci7oHPp4Xtdt
sxNiixfOpI/Nm8Fz4SJ9hIx5DE8N4SEVrVIs5mgembs7FolRcz04nNhk2ZXd
YzMJ8pMOC9akOxIFB4oXBSTpP1PEK0Y+I1/jUOcPqE9hKLE/EG3hitvTdbnn
LR5xDcGgHTHuUuZkiTY2nz1aFHKXjnGVKTzjx8GLAaCVqvVM97klIrlphjir
FCqkM/Q9fZlm+8hjHSh4AqCJXyBXRCYQLEEBwdq9HVz1MpVLNmEJo/uFFslW
wdR4eDpfeQnO8JfEaTt1Vy42gYjiUSM1xz7TI/i0wjkb4A1eZ+seXUZ9zaUw
PtFMuoj07WDOHPFYal5Hd5kHf4b6CaYhbj3EKqIR3YTga92rpkMEXc2VUTYt
Ffc/3GyVqhqXNXFLtWJJl9raqiej1CfnNTuqE2yhXDNSPv1w+BE2BLXtxBAY
NDMe4c/Kf5d3/XenmWcPsClhskOSpathW//uPzKGtrOGZE60YQ3haJYCzyi5
bpJACqJxQjMVTdE1hlj8VSqEsW7CbUOj99oww/8+e+aMUHIg9hs1F4xb02uC
wS9HKb8PLRbOERJM/DdLcFzGd4WyYVHZvJdXH7u2hWXl4FwKFMA/UPBfYkhl
kW+d2AltPQ+RUycvgaJl6PH7ffG8YMcHiXyPOrumYZFFkI6R7tQsq5anuTd7
yD5PWDOrkWqO/HOrXFzx90x9P4jYDxRzk5Pzews/TYtciXqDm5/xV4rT1UAd
MwuaqJ371RQ7r2jtV/s8Ij+xSj3+4ME6b8oUR4YvoA2LvCsE9UUeIHdOLOpD
LJqrho3xePhH6sV6MSwqi6cVtheocwsKFQN1s2F/hZoOVB87OUbpyr9ftlkp
UOZDYt9J3bG7K2uoxqdLWxQtKjbfGqJh6LkA9QxTGpFyNqcIOhe+1YAXZFps
LtUSdeM8f7DZHZii+knbLysk4L68+ZdFmiQemb44lenjmStm5QyVKnZsJnaA
OCRB+Pgcl2QCwt7AVUubcCNH2Pw03StVKdi24IjXP6+8MvaMmP8srSyeQNVJ
uyYnBjq6S4m5gc0eKo2E4ED9aPqFPB9HzIljTL2JLNgy5Di/cib86ph+iCOQ
rc9JNMiQuniBtXqDUdLpjLHm1kQc3o5bv2UgCm5w71pBViqATPcOa/bVlJpC
LZRINsKJ2qJ5orSNpDEOF1in1SINf8Is7xVre2vYRbpGDdmrnb/WHvI6fIyl
NQLo12yd767CcLPZZhMzheKYPc91jjfhjOWegy9bZvTMLLMmSJqNj/Bwg/n5
NDs+fytCc0r5OhXo2ESGBLXzsh96PKgFM93SX71s0lYQeTUOvBmSRWAzrppH
J4JZcj93LK3Px+v0UZ7HRcaTpDyPAGUTKqZSfIvtrCqP0uVrVFsPVL3JRMRi
fia22zG81EUpZBc9rGkYIAIUUXJob3DdYrqpEtneffdl678/fXEw1Nqmn9ah
G7N3J51yrybuq5vphINtaWdPYSsxIA47PnB+lna4g+hvzCNesVywktzCQapB
XRThsRXkB69U2W1pfxmnS0wO+igx4r5l6cErJrdLoLPnhzcStnO/fPzYGW88
8KMdCJMDGtfw1aB6OoT2h7hJehLtyT7n630V0recZluMVZHTnMmAQxywBglp
SGOCk4YFfURj8EeN2fTgKCLgyRvj1DRcHhtm70cUboY2tcDf3pco1dn77hK6
5ZQpRmC3+gnKw5jfiWy5/1kJWwsx/FpvJAUDaG7MiynHwV36H622AmWVDeK1
X2QZd1/qcA+eO/WcGVOG/iMilShKXWaF06n1eR5VrtfEO+3Ww4MCmAHCI8U+
KMt5/RhNNJhFxkFC6YkOC6Li1cRJSazsILN0ji6nYyncJqtYuA4nHPozWdN3
B2hFRucMYaaSo2JrDY2Z0hgBl4QrExaU4mwvnOWlqFsdywn6eQsL9O669TxK
tYx+KvOyOL5nTmDcfPDKzu9m5M+TGaKwWHNg9bVJfj1XwBSsoULurS9mlAhg
rpXEKEWc3L2fXOB7r055kvbGmXAzJlm1g3woze+lcsUgYFFGIamJOqQXfrz8
Jceqa+svV3YEZxTTOqnW/tBC5p4T+tCwg3QhMrhqUiUwCHTYJ9dA8KT2RZXj
qbMG4IEx6IkGzeqOqYg11mT1nax2f8wm1F+iS/AuRdBtNPEJdcN1lHwVcRVR
kIDU9NXpBVDlaISQP5hZPfsApFJJONvA33AINQw/NVn+rdnn28OzKAcAJ+GZ
YN08JZdYloIVfCK/z+YEfsC9HT16z86CzWuzqIXjQzjDy/TU1fApyhZJIxv0
O8kNr/ilEd59BavKvVExDRp/yl+Oi/0CfBcIFCVBkEAkWmeFdcQ9oZCu8SsJ
594jXEooc5VgwtKUaeiFCKj7sB3++DLMeiiFT5sQIXGapihyg2ECoqRHoGUT
h9GmB/ZHRMUt3CISNNhwbX2rF5Tg7Mov6Y4p8AOvNAwvEoPK4Vr6jPuH0wAE
n9rNneaV/6NsyWyXE0Cn9IqPDTisTV893TMKUObSPBgHpa47ae9I645FhyA+
tmYBx4+f+vvkAU1Xm7rSQebL6lML93t313pEH0+6QdC/AqjR29d9YK+K8JdD
fbVcWQL8UDS+/viVKFQcVVlshGuA8shEBFeVREQTTjzsJjZlm+jsG6/NUewn
DxdqEdb5hXS8ylAcV8PosUrCs8MccicThcwHBLsiYSbcL4U6bjejZGm/rdtO
A9gpb2cnxcZqRmxAaJMrwIpI0TvtQwy4UGCpxe4b4aWuvtkwGynAHWY8AO7o
jE3bzmTKKmrNi8p94UuNZdnyFeRK0Au7aADeHX9qT13EuCiXQzb4XD7olO5t
Xuh/eOkdY+1EjlpAcVeQWePE30Dub3cHeieFiP2h6BHgwzQkHOzsZ9mQ2VDq
GVvYlILX2vUL+HaFiAc3MqSs7Z7fhZjxR+T1eZ0uxEMYBUCeaNpUjT7kxWEA
DbcDXLJuqYW/EqcCs+d+DcyOKe2Z2OKDaALxkLPk9n5+SYcqnyoPNV+gQXjg
JfHjFGvHRPcDCCjjEu4tHaT5+hYqsiNDINAuYlfyniRfRS3noHc16QUQR+bu
xGeRNZ6ETwPwHSx3zYdzZkMBPyL4LAkOMp4dOswKw/wz9jW0+G3n8EvssFLI
daMGPUvkSMCn3SgtgyPBMhMRahddVGww6MeWKmwO+bdNY1gdloYM0xIDrrgc
N2jUTyv6QIfdJIWxphssOF8aGr3x/SMA1cuiEWn4zFR5kBER7uhrGbJHPMY+
uz95aydz6jxZKxgeuI5B3jTn6uscVLDNLMXYYetlZDyNZtN3n6HcWhqApYvg
NwxqgzldonX/NQwoyP8C1JKi+FcCMo4VTFag2AeejoKefSKPGCoXCdW/V4AN
9QPRtFj57VOpqUtm16QMBBgzG6OTv2/qqoHgo5+Ysb7MXTinGwJ2KCnzd9d3
BdzzP1sk7UU5SUOQqZqog6hnKUGH5gsMY/AsfnxTmCrvao+qe2OsBfcb2rHI
FU1T5d136Fe7wkuyZRmN570oPl6C278PWcOZNnDsiTYz3pfthrQ1l192od2s
GGdur8u5aHdel6n9PXuCsDzIxvZxTk1C3lwy/aF2Oi0qXbUwxAkIYUQ47EMA
DTrqEgxWcfEllZ1GETWd/q7ZD1kVGBXRjROpFGsGDlDu4QnP6B2Yq52NIWtp
OcwXgLo8behd2nHwX4TaeCPX5vcE7eqMZ63AEbf62ZzvMYlhAlrETesZFycf
u+0mOSgGSn8itPYONBxc7E9Eh5EuTUOUSmS034hO54izQfIt2+dvlzGOXz5J
PZIJNVX6CK1d2XFgcZg/Pse0oHR6nQLgkklw/pbgD/GRFiqNGsuggSx7Z+wQ
cbI9RMuySLg9Z5Ds9mz0cKn43QCDR3VXx5PhfWYSwwkFqEZR15EqrZrdeFfN
xblI59swCAObwaYuk7NSDFN0E2rVfjKjwt/umrJmQNuoR7AMiW2bn69GcIWp
1nM2Fxee/TQ1PEGpdyscca5lFdpKPkX0DS2fT2fPNyKr5YWLOgytCJ0wXZry
q18sctGf+xPKSW7ojY7uLd5qWT4SMV1MzoOSGvITYgYGWii34gd8qBn8oPzY
v23IIQO60eG1/zpO3LjHdrV9nCnMfndcU5KastJH1CpTo/gt8FilyKFpWCdU
qXzTrMBFLrUvuS5J2XoyC3MWupRarRo3KDeM1u2ltWOEQZc8yxSBk1m1W8yT
SHq1AWka06VFkWdFjYJnJ0pmTckBcdiqcuy287xkwujphGm1mY5zO7emLCmu
LgPI0umjoJ3iREjBjYhiHj+sBcKgSkQeEl3ub4lLbZkEbP6BiWVnSM+zeHe5
Pj1otFxZrUfoHCz3tb1NepVfQWzzgyiI372DT2zZ/atNdAcrRAnx3xr7+kCb
a8DsL8H/hG0ejjCbGBXRaXu4OFDTHIEteX21tOwZQKTV2mD07R/qEImGKqIY
VBr0/krCn57pX7l8gZJ5umW4dhZoq0/8czTarxC50uTuKPbUx454BZa3col3
7oYxI2866JHgVI2ctgzjAvsuDDk0EC1Xl0fL+TEclH/05XrkS1DOU7H1FFz+
315qtfOGCQTKjYhdaP7AZQZ5z+2hbrHLZQceq57dJBXuVu7ZdG59IVIz+FNe
WwUXf1FcpzcAjNi/Ssp28y/U5ABhxqGIcYnMghXCJeq9xKPcJgSMXO86k+OC
C4UPXQvFsLQzjLCpfrC1MrOphQ9zGbNdP+vJqYlT090Ub5sOjG9JVB/+1BN/
ejbLMWtBlVtoYIfiWb5icl0ppJGJQl8MOADpUPCkttay+n+ekFCfrDxLMaWs
hHbVARblaAP1xYKc13GSpzKiGnJeTk7mIPlO8PGLOw3pbdbplABE3lOhTU7e
c5F3UVFvMmG4gwUq9ndwncGKDJTh3GBvxbgk3kPchd+4N7J8jnydAP9UpTzY
SYv/w11RnGczeTFUeXi1zn9NNe7OI9C0jWhSoNE+p6Qxe9h/ZxS58SE7nkH3
mmahBEkIDgavPXqQt8D0zkJWdUk6Puc5PuEHTDC2DXbA3wS/S/ZGSNGOsdA9
IA4E0fETTnVz203GwJvvlG3adon0c193djwxpIABfLBx6+6hJUAhGiUIsWqM
qe9jGOXGfKwlsmL0JiG8bTZvKjagpN8y163PS1QLcHucvUXhWj0MJzIkBSNA
1XxnKW2/4ubjS/KzRK/4QlrEHZb03QR9WEOVV3/xrzW+Oxx7b6bJtTAXfKXt
PL/3ZYyqIjOi2+4c5yf6TFmw0cCYkWlktnhMVKQt+3sgsRR8d9Me3VDPF/Ic
PTM4CghxShN1tWNrMyEt3k0SVq0kdMK/EAXL92LxrV9+bXiF+ptX1kth1wfZ
3h9nE+rKFGFOe7AB0c/2+QiLxKVqw5Bn3KGNddggELp7r+QtaGmFMjVmAH4B
bSx4GEI63CQCb7xugzxqq9pQqXjG3wuWPKeAT6oFj1GGFjOUl8owuzpVn+f8
Ga1ntP5iMk2JmI8JKLRPoMRh5jnQxwFGBR1/CnH4ph06o0Y7ZjOM2ZTBbk2P
t0xuupKSd01pKi5+pG1VRmydrXmpSJWa3/QTNxccUAinUQnfvYOHI0CuqjlO
14mp/fes4/jzfsKPq6erN5n6W6t5ULMTpkhAscSBhzBezo3me91MxNUwzaXM
ZGjHHJFazzft5woCfjpXnpxsIvaAjqlMweAQoZ7HV682M8Ijp8Hv57TQcUu5
xA/kF1/546CUwCNBWP0PG6ME+0WAITHCk3zIOL1o8wehC702MDkVXIN9meMy
R0fFBt4p2yqZmzPt1fp6r83g+P7p0HPWnVYLKBxWYxypw7WuyBynkARNhqv6
FlOiqKc3is5qe+YxlbaB91S9ZfmHjh+PtuhifoUx2JC+So7FB59hnX8RUDLN
0U15QXd9qPwRAGltYyBBNe+P5Yw//jq7gE6NWhp3jPWH0KF5+5Q0GfngI1nI
5CRqBhJauHxWKLgL0Yrg5URdDWHXGmRvUcm9TMWCMLti4omPjxj2Xl+lQmHR
0pmcALLYN7GRyvjAj7G9FPk28REiw5a5D9OcBu9xsQZbqqLbVmdSpJ0WsdsZ
hWjLMTSSObnbehfm/4iakMkTVusPnA87JLf+9PUdRD12wU6plKyXsqMXMwwe
hkFpGQTKzEq2i4LeFHE6lCMrKUh5+R5O9bsB0fEuOtoOEH3xas9YGqb/xp0g
Qi9FwZTp8S4MOco1WkDYBTCUclX3Pyld59A3xj//V+X1k+28BiCQbBksqdp0
Dx8gPTSje0ku87mtrL/ofCN4IyUDDAXUKftzeAFmraOQDGM4E+vV0rlBOMAr
5+aPbU4vd5Vw85fjRWn9oIfL0L0NI4Dw/L9jjPulZ4CpFFtqtWUaeBeSnzjz
DTlJcnVHFbubCR8Uq5s2Z02cs8kK2CWOJvCM9XWHgPPNbCR6/fmt9FhNt9lm
OvvkGsCu6gaqx9rotYXem5EkXLSfSk8gdYa012/F6i0lIH5IdP2/rsZjnUJ0
9iIvW1QEMJVBMejfJ7iZPVWxZdemmcM/4IibeGBDzEMuTf69gRP8p0kNkvsE
CGSCTBtikgQSCx1k0pk50cdjw5Q0eSv/1P/99UCn6/T5XOSE76ZdjT7FuUcS
2/Rze0QqpHNn03X3WGpt9hgFcbeTXqU5Ycu7spp84/XVbdNuFRUstakFV3vA
8YoQ1i3t0f2Eu2u3ryp09EU1Z1+VU5r1Wpz2JPfg1xO1QRkqv3JX39WxMsba
xYZ9IWu1rjdx6wrqAS1loMu+0nMbbzkVC7WGNZR4tilV1WKD6h315WRqisjc
KGALKqWQOy4HdfEq6L5vPTXRFHxOLJNsZd57G9pFqKPSKx0iSsTby5g/jmHR
ssn/QGX2ff2igQhSII71WqNy0ADAnnUOyqvLy+2saLE+rnN3PH/qEKMsgfyo
6omVQkJYzF3ruZIdyKQOW3HBRynMy6nkNYAbBQeyrocoIXYD4U5KanIoBp6k
9JNcZHI6PI+cP0N8YoO42oIByLve5C/mmQZQ4R9zDl93Asexd5FCDbO/Suba
xlmfMr7oYGLMBmxAFVms6gQ0/BL+ZSxKy+TTQyUaMT13ubzsTskmRErmO+bv
833WC/29zjbv8ula/NeEUn3cUCvC1gbzLdsLi6D2nq6c/2tNMsLW7rDBe1xE
pAsxg+FhtDsCSuJyTHHhmKiSJFzOr31Bj2B3+1fQDEqrDnFXlbC0ik2RWcXE
4HWVie/0zr2cIldtob5OeDFehe+fXFLD5MjGAr54tu1sCgn72gERU2e4g1/D
4mBTOQ5dmUPimA3Nzbyn1kFxUvFrXjOnCi5J34TCE0u/+jIXnvQrxOaDlV5r
K+VPg/VTESwZ0i1+70dkmtxL60cJEpNFLwUJE/QZZPec3SXjarggHVgE1zbJ
4BvzGABTcsXvnFhECsEcSEUQ9iBeDfvqqU0cTofobnuvqxvKtr1QR1FO+XCI
w0I3Ej6jNSifkE/2n0eNTAtNd8wZOfzeHRmKXDqXy1nheR+lRRPUTRJHOgrR
Mb+8zwYtVInCquFEkh4NUwWwbanRSPF3s2rZuJYPkK7VL6JNH0qKtNYqA1bf
XiFedQKGgdVrJcR/Akv2V5N1O5HTOo0NGwdjjXoHoz63ozmoUXkgaBzeYQAJ
sdWioDLNOPJCQFf3EbyVwQUvWkrKVCoRjNj4juRsPd12Ab3jJ1XozBvPu2J6
CCMTum/V4WN80zNnD0fTjD7pTlDlfAyZyW/dpbKdvD6Az+uohyMaOflN4orW
RkMQyyToHwZyHOnG6QWKrGgdsp7N7u5u8q0XCysZAGEaiDC5elvyqIbzwDS4
wk57RDa6sH/jawLRSDKJFoJLELb8DWo0OpNsPU/hmnKvcHjULdykb6keX8rS
uWjYGZOLS0o4iUjCw7NEyNjCKmPxwyHCuvHpyesto2xVHwWIz+9g14goaAiV
r7203yfkPGC0eK2aPZBf17k3/3e/u/HawyTX8I1xIxCrfD8L70OeO1JEtT7M
Q4JJRK0NzUCfvatEcBvkhXu8PA4B6C4d1lJU6uyxTYFW06NAzbRPVd0jYF59
YTMbg5li+sheEgUkp+QkOT7iCx59iJkE4mJhDHmMZCfHVKpW9YIP24TJMfKP
WfkD9HpZp1xynoLwI/72HxAcp+U6nEq1jAM96IFqk6hBY6NvgqGQ2fOBrjvx
bGbLfUjgqG1ps3I2dSaTHGEK5Xd4qnBD2j3hfwfqL+Ez6Iydd49yVrd0h+dG
jBYBBM+qFeIs1j5Toc/L9HUqjo4KF0DKKbOK31HRa6JFHSE22M5IH3M/9I56
niEBS0DMNMuaNz+RhSoVVMl7hMiLCA6VoXpEqM80xC3v9/tQkaWqT2TyJhkH
Qywx7SrolQFWI+ILT1wvhA6qYnlLxG4+UvgazRvcIgYQ2CMz7HMTieQ4uINL
l1LMw7n9S4hmN8kfnRybPc5H5evNMq5jatYcb33v9ttG76ehCGUPHD63rVnh
DuweSOCGd28sV/iWDVpzi4zv96Y+xVW6vgHNk5guy0Cm0/gE6u90bkkuTNWN
ZwNPOXsUNXDJBOEj6HbD+qFDyH8uNOJ2O9H8fBg0YMKynYbk7r3tw2HZrYup
rvaOpK9y7F9j/unvCKsxiSMa3+/nD5+pG8IEhoGqC/fG/znd7SgXCcllU2F+
GG7aMAZQDQ/by248i56aCJpcXM0oefHjxFacfTjO/RXLYfZTPFLZucsjqq7s
9XmnXz9rPOFer28QtOJn9wqEj7OquHfv/KONjg9l4MW3l9UWMQA/LBGkQeF3
ToD10xfUOX/51JmYDiTFHkSuVsTHT+plPdmOQ7AvYR83YH+0oqIBT5QVwv6E
Hn9agm09F+zhCB4rkP09j+ToVpSP2kDRHBPhqlXf7poP4yMB1cJpVhYxLoqi
6zC4zmXFz3+ONmE+8JD4vVhe/MXx+UIDj5hu+l1fmHobSrS/4EteBRzJLAsQ
zi/FlyH18w+3Jv/1CjaLbZDQ5mAgOTyGDV4U2YbDVk6y7NQzbxENofjT/sa0
3gOPVzYUQKc/GJy4suIQUIuvkLeGh2jZjQqAJsh5qgkeZLIkQiw5XhzwqUcJ
EoYi1+7E4XKqUezXlk4JitaE4xROGrfH26tRynmWYSBwTyhyB3z+B45uSFj8
YmkeAZJx248APIebP2mngU3qL9UMQM9orytf4S5mqa/+gMkZK1nZgFKGLAxU
D3P5Mt6sIVSooMoVui5fLT275naqA3qKYYNziD64dP8V5RkJHrnR/jlwwnLr
k+xmAzmIsQigWPIOWJi99DoTh1x83WCV5i84KX4fmgYKAU5+FTLzDe5kQ1a9
4zmAaj4tpbk03a3RRi+1QM1nvPNLZ7ZQQnyoe/isThcAU1i6OkOxY8717c+Q
9enufcAUwRjTh/2dfXrD440ciUEwd+IzF54TLTyf4bYdoL3J3viZ1nIPXzCR
SA77JXaVRPmCeBNzk9Y+4WRHQisqV5BtpnOU4rsuyjgFr5M5HXt6AhrNmrOI
vF0nVOSp6v8UN0LwRc437RBNcRJ8v5h0tzpCRMvMC1/qMcQBuVTGV7lmz7Nw
iwtFHcnz5NzWfTcjgr2z+ZebyK5nX0ZjOQ0dqXwSJAaXevtLz+GEAPwvfBMI
tgwBhabOANaVmEGRBXqSJEMAuzV+GJRy1W3JR6BlavFYCACcTa2R88eV5s0z
zJnwrNA5pjiFcRHNHxylPYd+QTI+5mYDZ8MBYYSSVDMcI/12dtpAcJrmv8kz
FnTEbv7V49tdCRpOc9UFwwTMhRQv0GznvfgzSZ0V4GtQ5K9hZsLZkoyKzn1q
in/Z5znnhnk/4aK8pKLjq1hNn9uDG9LBQn9C2H8Ysez+jQWbtUYH7sy77EMf
7Lk70FZ6NNZqRicAYQEat6t8ARhzuPV81liPfPy9hvc6m8G37wiu06jeAy6A
O3jr+7nuJz3v/e96ilxR1wSJvfMT5VK4/hh8oa914g41/HYchr8G07wxQzx1
y8jy0wtendSh4FkUxRivRJJymFdlHqJTltLf8gtmpee+0f0fnoJWN3SBQ6Im
1dkspoUE8BeLtqfZ1vvTI5WVKvdKdL2pjSNi5NdtNRMpl7jz7akAhYWYG3H6
WNOXq4ULhRV7lHL88kjfcVoDRYdEQ2f4RwOst7hryJNi/se6hsNKCsu376km
DlZo1ZNU2+0ZW8ck3v8AdRfw/VmJ/nsA1c7vNQ7LMwOJ4ewbiVl77P59uHQf
k/RclR5ojHiZkMgT6IDJRoCoPMkBO4aJbKOCwl5lqxA4p6jFXxX16mUhq3Po
Nu7WAq3oIm7ZrZsvYyuz7fedonL2aUU7bEVf6TaloefTKKXKqSz7oJPVaMWe
W5WcVYasis+ism+MB8CPQnbhbHuwTY6W16U9at0KjaaKPVHK3M0yKASFWNG9
Sw6UtxwIYCi934BFCv6sh8Kn+6KOlcu1u4n6ELGrrdtKy34x/6WwS2+ixmh9
aA7FDi1/+1Ef9eLr1NkJrqV6VCymxK+6/uNk7fUUPka2+c4Xc7xYxoLBRlCE
4sF9F6ErTX4Z0rt1t5mX2EHmC0CJs4hhdaYQ8jwws+VL828KVJqizyR8ow7B
huujpe92VC7fzBMqJXKux+fzIdJAhph2j360TaGdNbD+ph3nCAwPDctRbpvz
/9VRPKpweyH9VrrSgt9AFzRf8EZ17xIuLpwWr1sujRUCsLZZaYjXpFqWO9Cs
0obBwZM3GywiLEaG4Wf9yUod+FI0BdXOIfw3C8tuhd/bE62Bh4fFdJZ2fQz8
egZgrlECu0MWdbBHxKVu0oqkc0Y8dkdCHVqlIfSUfYHBmpB5ihzASRx3s3Bn
YyHr+JmoYQelsHT/S/0ZYBne+Tq+EYY/2/6i/e1Er3PE5NF2UQ+tNhGSWSXw
tiPjJbgbp8K4V5du0kiydhTit0Z/4dO8h0Bx9a/SMX6I2TnB6qmk/Y5LsBQo
F3NHZdLjjmxVbj2noDJCk8tTRaT6tM3+IgWTDCOAWm8RnOHHdzuhUlhKd2Tj
C5VkHe2hhVDi1ldIlm2syMYKCQ/XYWtOyG19dNJrZolW4jW9PiwXdritsngC
1ugEvtWDq3jWVou0Gl5BWSbhsUXt1kIdciP5kZM+vBrlMBFT0Oc5z5oQqU6U
kvAX/H4ZaRJ6PvDUXES3Zk/xTfwrm6MmGJHaT1ST9C6xXHKVONw3F68Wf8BW
WqyEYYMBJ8NXtPLah82pig5U8SL9zAO2wSC3cVfsukI72h5Sl+hRS0I6PAEK
pBC0MQyi8lhL10dBR4NLiel6GqwemGoH8fJsjBiNhQbwD+OhUYWZfOqsBLmA
U9AsBrkYq2+JBJwN8WcwbjxcH+v9wCZ5vZewZJ/F2y+BsIUbUVrEAItrzJb5
i4MVKquX/IFv8ciZkWpnQUXm4zfYyiOEETVP6bOlWwDowUQ97kiqjXnaGozw
lOuzE5iEkPBatrfhiShi7NIGS1ccLnCqQpEPNWbW0uhJToT0iiHuwhyl8RdA
yI7uwGWULlDiG9WWvd6J8R9W+HplXmG+QNb9xsboJ3rmW4WYXF4bNOa1K7EM
xUlrGsQu24c21naOXX4x/WJ3eLD4WLbQAwWPjeocIfZrUKe+A2mmcTYEmErG
XKFnRJVYMcgv+tcuVbubDwxll/h0fAJChLUgyZvVveSihrt7Qe70Fa3tpemi
YYy6UwJNOx2yHbaTGer7XUaaDZ2/RdhXrbLoSGgPiIFMJy02BiawTVy2VuDB
FP8lo9k0pfEvtYQxnljS0AgmS2Du8Bl3vnDrgHJ64El2qQT9syj7Rgo+UFFm
YgujvdF8IKwfIflGyxl20kPGldilfjJ/i+FUlksWgwx2srnLipFScbdWn9fv
1UBrRcUBmiq+g+v/d57xsV0GNMpf4imRpYjAO9J2zEs8SDF8hf8sC5HU6fTi
plxGG9OgDZvnjYqAaMJeaSN8dbWDZqw8GbCJwCJClwuAAhuZy78kRLBwP/9u
Ay84pf2HzbBWUkWZPpwr3YvXAW5y2lr2h4ERner+5S6oGwRY2vBXMtvghv4U
CiGk+LTEfW8y54+a07GR+yvlrIe84UBPYVzTvmTbVFkjx9siejGViID5iJOc
M5mwv+I91x6QsqG9ndUS0MSRmRMd9o0s2KYiCB6s5DfuBlujuMXUmxJDJlTv
q4PAUAnrmQhHwkEw1j2g2e/a847fHeSfLmOngSZZgVdSlmCJC0dP+f3/BPHj
NAB/uobq6oQhiphwdjBK85Tc3jh9Kc5IoHMW3gjJauniXR9aHdFbfaNVzAqd
1rcoMvHj9w0Di0ipKZOyQjtJ+FZlTGId7fdO6UmizpG0QK6/HZKqsNYwqCNb
TmDE/pZ8T22SRuLUXDj7VV/T5LIC+KtUmpma1v3sTKdH3LpQtQHVZIePPrVd
+jr5iRNXN/fpSaOgIclELazrZyVA+hbAYB+puFOUl1RRnv9jZ6D2L5/hyz4E
cbizk2u/3PE0hDz+BGDEKRPwpF3xEIBnAG1YOM90xuoHairr5GYnyN+1DGIh
IPTlsHz7FzUzuqcYkc7sk9ZSL9Y+hbasVMnBdnj9GAFH2KJ9437tGgBnJDpI
+5XmyCayNmmJeqAhGR+kvT4wzC+/s0R4JcYusZvDd7QTqRrMFEJjp2+gIfXM
0E150ojdgF+VNEtxPS2PsSLBp7xuf6E+UP14K/Hizre1c1ImI1orZcGOEe5P
kcHVfrhWxS6OcdTotq8Ua2ox7AVeYCgIOFSCJpRBVWVuR/fLS+VPylBti072
lR0LGpoJZpTYmCcKpSIze0iwGbgKvxQOwIt5+GIL0MzHpOuRtlJ+Vj+43Mk/
uvU1qAknDriT5sqrJr7+VZx/sBpE/D9GHV3B/unjDpupbhBnp4KkuQdqHgjb
w8TyKGVFFQlPvnsp0On31xZdJ/BTZNRvHgeXPyyHm1+9yb1/69TjhWu1I/Fc
WIf6OP4pP7ZA6BtB0scY3CKBABbffi4bOEhLfNfkTyiT99c7pHm27AUlw2/H
Hpvm2dw2fTpxavDgK/WNxedZc1KwR5AnSrdTMWdJFbjjw+vwX6zXy50U1ntY
zzyCLj8FyaL7KdIDh41vNKvTWqkT2kT20q5q1TrZN5c2Zf8DCKZy/9Uz0zKi
IPP+TsVtTvIdbo5rbXWRsYzzEgyXvpUJR9vCamLAvS9Q1OufKN3LN45yXHEv
8VC1AslrfIoPkgpOZ5Hi5r2Cj0JV/f2m0+4lhRkvh3tz85qmhb1zotyJ0kTd
w/sPKLqbLl83BLv9naC8gd1pSjsORqWstbGLIwRiDyNsvse4tZmMqnv6HfQe
eIX5gV2zV5u0WHmej5LEuve6MfqS0d0Q9bboV3wQtTe3yoRlcCn26VHO/riT
ZWmqNdr3dAk8DklLQDlKbG0fI2DvI0icpeHGO8VjQGn1Aj0g/raFTYMWozAx
i9Fm48/QGATd2YHtzxacgK8gsnOFU1cJolp1EInGL7z01rGZmxEFdcCFJY2v
EVimCG/FFyoblhmryRr6ICN0PkNUGXbZwWLoHvgnkvcFzgYcOkuwoofjnDfy
3nlu3Az3gMgSqib6luAlm2+mEtjeYa/dGftLTlXwr4MG0FlvcG0pPOTSYL7A
wMpJgiG0nH6ibaXqToGhFWwBW4Dgexpc7oSp2gwEp3Nxx6MIIoDGd0VHAPaF
fLOIDMB2ySjuItomREIf/ZAL7D3DzOkwLzU2wsbAbie43GN0PcdVRClGMvza
JZQs3Cdqm1nA1hvlezXai8mC39x2VXqb1Fbw8sctais428pbeeD9gfLrkJyu
l9RFFLOV2Gw/vp5Ayv86mB3fu2g42dnD0fuimXOR0x5AQG7Z7rEGYavnzdkv
psJEcIf8qmoUXciJIz/hwl2kpkZ9IPBjpQko8sDIi4HWqOVFbl2liPZB9LD6
LLccJ8pw8xipBR6XDdImski5byZ2n46AKa9y5JcjO/ge83bHWON+bY2LGO60
hT6yK3kN278jtiAx6lWVbzsPTUqp9bmdO4s6wQw4U6t70U8dk3ciE6NXXRca
MCxXlS1iemQ6qPdQIsHBOwPDfFW/6Z4rgT4xTU+W+HlZwlRMjSu+hD69hwwx
WMc6mn1oEpvmczCXlU+Jg3P9+SXlPyig97pj/uFdxKd+JbAOaCQe+Kw6wGHc
1KYDFamwBPYiRxiYOC259wcX8zVgAxBQWjAoZKwaNzAp7cV1LO6bbJZF+4bA
XCIuWxX8In1L5pULPPwoD77NvBpLqpekm2Fp/rtCWh8PnjCjZInaNbWSPrhQ
89MfKD0PObteF88bR/3SfPxGGbYhpEJrsrK1qGwtDidT3o2nd6P4tG+dP6xf
HUrgw4B1zhtrSH9oNtdIbS8InaebqhrMTou2Alu9xfGQefHpkd37e82k0HOe
BVmAoXSV9DkY/35Ujz5BP95LcT5kyA3dRlnyTY+apMHl3alD/5EML5PL20NG
l9PYFrX2Y2+bYgk10mrn8tugPaLJmhKYx86RhIEDQEL3NzN0eczhffGif5Tf
gYkhEJbOxkiHzzfIr6NVOSoHIqYH+f2I90bHH9bT0eF02SFQ1KLRwmvXmEpM
jXkbfVqFeD9Kfoyd748hHJUqJUTxvNEkLPmMHEVJqAFFOdLrSlzxCGoUNc9D
wET5+uvYNWm+qdskSYEaslLfngTe9AWAI46yH0AAj5F+A6hSY6PfDdIu2G9Q
yXXc7ubBcxo0t8gnCqQlQrXbXAPSbzWR6OhJZ7k718i3GlWhIUogWNwzN8l1
IOzmkSbO0UYxdkQRadGhhp9QoWN2oRV4I01DtGOTWCkyCNi/DaAqqsVsyhcd
22urBUEMt1qqsFolAWk0sAn82mEDsd3qB+xEO1aAI34PvfjFIZq21rtDYUSy
G2hnH5Fgd/YTc6SpO3sRAwhgB5duxbaiJX5GPow+DBRJqT+P4hp5bJXAHKoG
J30UcUvbI4g6HzmgGds0fYrJ0S7sk/wcO4hJsRFje19T9FMaOUNkp29FCRRI
yqxSf05ZhmlL0Sw3RWY9cAyU6iRhk/v/LdHfXCOt1ohCM4J97iUzNLLAsd3A
lsi41HmCYpSGs4+uu0P4JnSujAfUGVaOGGyw/gBUgeg2S/8n4PYg5ABJE2CP
nXPw/An86dACJjbzI43I2ld31mvguh1kr2rVo4em1vwLam8TEkcBUEc6w+ci
9glJCsydQ6SL3aiEgSXmfRSu7IQPfjMMfrvOKJthUC/8st9UMOr238UwK8i0
+xjYz09BjChNshdOmygMqFXlJN4CI6tSjDfF99ZJPhRiBNtLqHfChdziknNj
9c/aqMU7acXQN9CP5tV4aB+/TtAHSPL9o5DZiCxytBgwTHh00wl9IbEqkufV
61yHcmiNB7tqzzPw6wbonXRTIW7lzjQzdTUpWaz5biqtDdUt1bvysdiK7BuL
hLcvjdyNFc8mIRz/1FzhVxatbwsBSOCXgYyAboxSaZHOtINV4XHt/crDI6vJ
BRy3R3PSnvODMifFGtwGa3+1cvtfI9n1vZb1BWiozHaV9Auy82HLHu2IZEiR
IiBZWeS1AwXuFqwIGd0lysVxoqvr8BS8LXOay/nsthNcyNjBE5OD48fMt1OR
nYAooj46S9UpeYAkVyVgbRxWKqORlcT7F6axS5NV1vBAP5gIYsN8e3+eEG9l
U7che1ZQD5ZNLqVYCZQegLXM35ubqmzlGTGy0f1808xWQeEU5L+vkW9PQUWx
qNtVprX54vCNl9YjsAaQO3aNQT3tzPn/LwgJ6g8FjK4oHPWqYWN00b1aSldB
YfKdOsXWVhigO7wqbxaP5vZm7aFySi+ih0oUDLFNr1t/StDd3LrT91L/MY5u
PDukPTecR0VCu+oAcIU+niQW/QJjS1SnP10zSlQnI6wfnZAzHxdNshKX0G6T
InGhPK8BdzYMpNtwX7RF1iW/UxhnJPTCi28mTc1pb535or1LGJl3HDGNH1oA
49gQ5kszdYu8d9Mo8JEzoaUDKudqTG4LdUfB1W/IkYS7ENqn8CS/dPapKqSS
3Iz7G/du7U76+Thtb/HlvEKlrIaMcd7uFa1qORMRZZzFgcPGEb7I1xIPWJ1R
ath3+Jbgtl2TyKw+79RqoFl9JXbwklrBU7K9jOQhMU9nUVVa9zdzeUqQ82RX
6/i21y+WN9r+XmC4v07b6WhUO34W3b/TsTNz1VBNpF5FE9LkiWNjmuqbdERc
Ujmmu2lyIVydVfLk4lNz+lCeaTXjuGbMO9vMinFqOmf73W85Si29cFgzOf2s
xMoKlLX1TtqXcluBdDXnt4g0YX4c+RnDNnjI11TAmJd4SrxTle1yVWkvgvFQ
Bm6nrLG6M0PfG9zRpvY4/ns86M6zAC1ezhc6tEb0HDTajqf/E2Dsw9yK3KCx
I5i4jSM7VVWOV6kJGTvVduoBqg+QZhOqsZB5S2yFSDzcuyTrMwimQsKc9ss9
Tll/1Xi4hWeV3vMaZPlTzo7HpzHposu+eDPMHGPhyDhGE22UHxcXGHMDbXCw
f1CI/1Nh94Jo032QfioNAHJha9MqgxcCJI+I8gerrhzP07cjdz0PNfQT4j+n
PocSDZDIrMGTiBi/wwlt/fPrdznKfJZAfTw8lQuBbBK6oJAhgnSOH0FGmJBD
S5zFAJgwMysI6x7aGZ4ct8Zy5kIt+ds56l7Oqa6n4k7FxL0kf4caJXpE93+P
XLBtdVCHdAHwytucEkuAr/SQ1rsPeQCw+I/Cj0wHP6yeDRN7vSodj8uQL0qr
r+TO9qY2hY968BOEnJ//Jcq/sCXpaj0llicNa20YxE1nM6FpKA0c8ZUSSGlB
kXpRMGIDAmNxuGXCNlQ1EPNKlvgkxyiJdRoNUtqz/H6/u4j8ve7fHx4hIBK3
axtcGuKRWZHh+kdAMWvrl3fODhtBf+13QhFT0Icdoi91grcPqeTqTJWfHLcF
l6xq6U0z7TOV4edk/UEGDuEv55gfwKgqe5ZdaBpwsQs9rlTjspGCDhmg5F/j
HURpWbn8ly5G9GHDrM2mPGwW4J9KSBP+9DMFynAbFaxMMTK5gKATyqKiCaWr
N5kgt+qUGeYIHPnU58yOkscPfn/SVteuihRwwliv0d0yZh8Qs/KPZAOEDL5q
80VFcv5mHsrOI60Bb0/FK394EMC4jjrDi9kanwW9gn0lH6iN9Jmm48bIhP8y
35ST5tS6gAnvSaxn0GPjnO1SnoFfyzbzDlvf03x06vMvds/mZfeWqXwZDWLb
v+KFsf6H7vTdid2NRmuDDNVaVkRRK8Y9ZXoUJJ+GMOh1zGFpWRJhZwX5RJri
tSOkcoYibpocekaAFGR4BceKIXaXRxticcRPnkNdTPEISjYePEullfrRjrfX
KP0XxVlPYDG0MTIC+klI98hm1XLLsE8NeGisopAeKku73Ij11Q5Hp4JqxwFq
DPNONcFLjRfDVQdrI7Ngy99OjGyTmIJrJJiapowH/CFXefDMgVvJHmF2axuJ
ETk0aklfqIWQU2WvLccnLuAJY5qVQ4cyUA+N1BWKX4A044fxiZWN0qx6wlUR
Bs900wcJxMCULA6v+YzqfT4IcXZGmOnVPtE378WMash33n4v3BTXzuEcJ46d
tpkR2f13WmputZ47e09l0kpJFNbb6Jzxvowqw39CMbKWE15cHblwoZtCb52d
4T1g2Lr/z0q2dNwoF5RTCgcHUOvN1Xw0hdtqUD57foywuKfqMeJ3m77cPd1R
/phwpQu5PgjPHY4m69Mf0D5Hk5c7AopByUlnWGlP8J9Za6oleFEKt1G9ltI7
0o2e34+JjJYk6V/9MUaqITSPPeABKmWT5zuOIJ+6p1NKojQzK6vFo+N/d8Fi
tq8CEJtJRQGAJPy4xT7SFjBIovlfIuwbWSjEXGgs0NPhaD79rZxjdTx6pnM7
m//3AGgvbTHboTp1CqzILvBIBm7oZHDxVO9y4/X3aENFnvho6IspkpvHP3N+
oKbhmIRpDBGlAcAn64Z73RqRW0Xpyw5qeR5UXD1GFqkEUAWbJhtzNi7XCOyQ
meCsDRO1OErVtJhFnPu0An/zsUfMopGD5jT5g3CBAWcKLWA42mqdQu2oQCtJ
6jKvMKNzLnIiMullI92xnwCpGoBdNhKrQidDd/T7oOosLvG6av8OhNmW+kfW
t+H5h23Al/6qURigo5V8blCPVdxKGDQCaPBWO47SJAO+cQQtOw6w/oGjE5un
uyXPlVqNVBMRXcKh0XNuda7r9EMAWza83yUSUjqlLGqYNbyYsJzJLIrqR7Qx
M16tI1mpiSgBrz2+Q7HB0Vf0QxqNKUDOLPVyBId0dGi1MpRCc69Sk5It5SZZ
z8U1rLu01IbzohnMIqXvbKD3juMeNGwDJ3pu37qChz3TVc44tzpMevu6R6hs
TPzl4VsHGDgv27Vfhv5oVYI6281MZFRWd3QxhV1H8X7o8DgsVwt4yK9s+vv6
zYUsga/WeV+0Wbj+mn5dn2xxWXsuaVy7crIi1tHZsVRyWdqGUySR3FDh9L0I
jYDeN6gZhMAJVnEqqWackD5M/81r+EBtePrj7BRKP6hNPt6Bc24I5h2pOryS
4s4/37CpOKSLjgeXB5Jp4AqBHZ0Zyz/BTd2DnucTPmxgOAe/r61Jjum6KFzT
aWKbGTjwOXE0pQGT2BZFRFglLih5/KMl6TswkTLg8vLYr02ZAS3jIoJM5RdW
z2g0B2UjqyB4tCwRmhrmTm0weXwg75oV1QCnUEEyK32z0S8JOlkrxxxpAZjd
xtk+h/xWIMHOyFTDEn0tyHztTRtrbjFpcTRV1QMoCpe9yeOgnBR4NgLw0Rw3
dvYqrdJ8qjsbOlNlUFVZxY/2riG0F3++w0oklXUuqyovlDUDZ0SEGAp/lrr0
BjgOaCBopvlzjquwlVrUaAGOk6KlTylBmmOS7OLZHi7nalYYO6jarXEGRE9p
dGWqbXReVHUTiP9qRP1VkAXquzj13F9aKkVWXh7uzlP+Ei2I5EVY/TNKGme7
pBFXJIRgDbanQfxbwRo+wLeppkjG07Hw50aYSucruWBr1E8naaZOs+fdOKRX
TgGwe+TTJzkX8fDACGbhkYfjgZpgHItzKUDQifS2J9RIJgbIDl3vPs39YVnr
7tDCdhG1WgdRgeRn+u1WcXxzcsnN0+7SBupfEzfwfcGzcLTRuartQj6qf3V2
GKGmp+KPOK0tnKbd68SGb0WaQMfydGj1z4gSxFjXPdjpRWE7638yPd4lP1L+
COm6pByBHipzyVYuPn02U6BbYPe+/LX3P6SK23JjmzeCVwsT/ys7vvM6zBc4
jLh9CpT3u9wnq1WvkPSX/9ucoUcHNHP1yQQB2ESPGmozT0/oAk9TfaLxuIis
R0WiPyjI6g0PSoJXK0oG7t5rIY6F1bg7tDgfsthNbN6tx1BmV/JlZNDyDN+R
PhlCp4DPaVvGcMzTPgVejJwIjN4m+VcYVHytQtxY3pVUAedcPiZhStgjsQzd
EYN49+7iHGFnrm+F8rVU77xHHfgtUL4tdbE/zGTwwjScmssNDKi+sxaHil+2
cgUvqRmXmGh4EF7oJhziBE4fySaQC880wv2umoC8amUqbSYMefiyxdt0Qjib
uYxX59R0MoIIG/q1zFJfhvE+1eH77kafv7njoIQ+QpTScsVsgBY4igy7utIT
KM2rU4w5wSddHIRzH0uMALKsFLVSxms6a6nBM5itXOVg7JkoXM/ltsJ/1sBT
/OeKA962gCaVCw9aOywpLt0Q0pg34XFL918B3tSXPprXJhJPNEgcxFJ4iJ56
7hRB4+erq01U5bYYSrI+6FBQL8VSC8Q0ilhEFc1EwrRVZYlGJ78GJJSg1xu6
SpPyxyGfIyHBCNapu8kS/0Mldpw3aHw3lbPmIwn0/TVWUMavoHnxkKjjs52n
ANXbQ4aS6S/L0jE/hC1b96j210wfYt+AkfKkdGXdVWqjVXnnvtFGU1BfypzH
nZRlw0eMNXwQdzf9V8aZ9inSP1kEaY0ykXpRoteH1bWzig/op6rKKyVfROR0
sxU5YuaS36wWLRyieV8peWfNWkyOE0F47PQLDHCA5l6z+fVxJhhDV6fX905j
pvtOz1HM5t52qNEHu3AIYPpY3iCegIu6MegkEKiA5m+6ehV2daJfkJ4MPnVU
3B7hDx+7lOCjP8tF62W+8ZuNNg/kTcSBHwImpnnzIMMiKuc4CiN1heGlUAOa
DSCqAIvLOXOQuObIdOz6gWqUpvBOwPaN3xj0oKDGfpL5UBAuL9+C97t9SgLB
cx/xhPXHuvjA319CntuWbN3FwTTxa1ZdpBBFXmYhCahr103iNcJ7VrgCKW+r
jAUvnmDfhSuNj0jOuKaUqsK54J+mx8VbtM3au5pIj2SlhvK9i13IFtVhaz91
S9pEOk2hwN05Z4ysXdXQ3/yOZcjxhJScNcHoxwxQnG1RqvE0EWK7VzU06i1R
ddNoLcJbRacEvk1zuTBcMsx7UUXEaiyXDfQSAhJYKYXloYPd69munIkuLPus
WssNhJV3LsXRJpVX5TY31nOy1G1HqHO/0M67jiURFaYN0ksoBwTryXTpw5CW
9vtj47h6Z/xHAFAo4Z6EONdw4yXv/cHlx0jelqop2zdlBejKfTFbKuCTSNUZ
urgA7eldFqLEPS6vfYuohgZGtXNoPWid7J7ku+74luJ4B7aHpWmAetXpHl/X
BFBCCI865PYqe+20GayD+jeuKZdUdqCvHXITJ0Zr7+jI2KACThA3D340agYE
pw6Ck2fzRb/MGWAxOhpfeO4OIwUps5tdAE1UQIG3mdJduw0joJc+Ca3rJavw
kCE5FfkueF72bUMNKwgAD8Gqv0QRcb+gSYQc0ud/uXEfh0xwdM9eaRU7BCVV
n6MTe7HtzlylTJNiv7ZfZh2ZB+BllIiQ1iu9VS/yki7jFwYcIkZQ+fxMSHby
f1EuYNOlkdQMMszqvot68IzXEKKQXuGYmbBCpSsZPuEjEQx3+mlul8L1+NG5
8PfcfbAckMhbli/N2swKiFee9bTjOWeV2jWws6vrWHYgOrAARliEUpM2jbH5
Otj9yQN6rN5HxasugXSfeuRERHgTKQGSlNFNfOli/w0KwJ2bYii14aJNR+Mh
xkuXOKpmu+eHt4oOJnU5yTU4SfjCRvz2UEOCkv7PI5H9y5IDeTR7b4evM83k
5LxrLEotLmtnc3lyxOiO8YbYZ6ggVBqJK3/tzS/jOkJexBNDUVyFgiUabGit
m8xrxxfgjYm124Pu98fzE9+I58sV17DLJI5g9J2T+aRZA/YJou53E78ijQPa
mc8cROgsrwBv9BscPys89itmnWPIcPtbTmFAuzL3E5FEW5/e8M3AlrCazxCG
aVP8+UynTMQxqbYRcByN1fWMCrNY5X6wpavaPjD3yD4l/zi3HbRjpCmyPuRC
9heV+GUkjKujnq5HyGLpzf+5RjFP2XlaguadKxZwEyoW1KHLUMHW7hgYaqsp
wAEGMXcASZm8OUK39mLAFE4l9AWwtVKmkbcfHLbzB0rkSXAvtVHEO2tVUzgu
ilYzUGhGZrTzxqzLRPAreh3+r52wFZ2hHk8C+KR1TftQOT/mvGA7RYdi4t+5
K4PztoFsge+mKF2xt9Su124hLVrLnFeEkW37OBbeKC/yeOIzb3H8FrQmQRNW
kNv5oQKH8d39oTjlb3HdT5cCce02MWtL7VIt31zOB1iy8WAyyKexZ9jpwaEP
lka8bGMmJVjWo7PHy4FU3gu+mUXvY1ZJ80E5JO1GdlkmSebFw8/E/0+iLorK
b8cizVneKbkZn1GU1mmgBxE2zLzl0EK800bkJ7VJvbKVK227aNOaMLpE0psl
jjbFp+htgUcDIZov7ubSAoncjgt/TPJV9tqekNcv1m/Qxdc00E1ykjPH0tSB
FudQbVltaLjOz7MES1NxG2SEg9NqHWll0RSK6uOR/SbE4hL81ji3cimfyTgK
myibMSIA7LoQcrfcp/ghUItbrQgeqNQWHRtcMSwE9ZXVErjiMehlW8EuHyo6
BXyY/7PSIFZZM9KBWqepCMbvxGdVYRSCjdP0+eMcMiOqX/hwIRQNQgMEN2W2
gWWeh15yKAFYKprV8uprAbkTpJzsmtHNWI1rjztP0ANwUTKCu/s2qALRDwYj
1zM2Zw+HdijyjLqBi1/lfwhVIv4uCgvkxeovDYIXxjQRamEnU0r+iNaVd2cj
pktWaRWhgbHNhnhxKpon3mmOj3lwhD4UC7tKfwHF27NnZoQ1PiiBFmCKpJAV
/UvnzCW5HUxeFca/A6LFbFUq/AmTTcXFz6GuSa22TZlNbLqcC/YmhoHOWgAb
n9MHHu3CeN/MMynSknIYZka9HmB0mjhlSY+tzCfQXUek/Gs2nn9pBdzpf2+x
j7Zrfy+YE62wvPNC0Rb3UmpB2ENpd3gMeVFKctVeeD/cGFKOiown6XBXSW94
htop6MtvV0Qxn9RFOe4Rj/0yTNEpINKS9xLmECQ5sAXTOg8+EYU/BFLkS8pd
8hGhMAHnBd7KTUXHNO6XERYuQWTFveW9hU7xxwMYH9ZTKl60jI39dCtPLTIS
T4kh8rmNjMdHJcwojzu04HZbtNDNWqSI8CT5igz4uvHEC7TgZfBMprRC6+OI
gln9FLjZLHFPWMFz0LA+2ShFEP01+yi917k119i3JwtsFI0aQUYhpTJ2jTWe
PLLmggweNP/C0Z+/vZdnIM/lUn+Hh7t+/XCAhiHcaJXGJm3OZuYsStn5WgyA
4ipJZtjleKiFaazove/W6lBeRFilQ2plmNyAVCzSCN6JHIIMmKtoNYcssoWh
hvOG39du0coUnpkX0MQ4dANJBoZcFMVDQqQK5cMi2Xq96O4mFLralvI0IljY
hpXzANR6Ly3CuVALlkGiR3FBLp3M3d3sJvIXouSxUHtMRpiRG+c1LEDt57p9
8advSt/AAPS9FRUnzdflywoU0agJJ+VmNYz5syhiG0JseI0PnrHa98T4pHHK
s+hgpavsMzZx0Dp3q/9/+HqBqQdU+DfjF00UFKsF3iClHAlQwr0X/Nh55kT4
YKkN7ldPkMulIZJ2eqOpVz9im3uIbCOehXYpvONX2VtM78bZdJ+AlKdKQ1Kq
IqhvIkxOvFr6fqcAjKO4DVNGzixcyRDgIDQ7+bsJPtzUhwVeLR5tFVfw417V
ufa7xDHH1wRQC9TzPlFTtn/mgt1iVRqeftM/X5AsgHzymXisIsl9X8yeIEXw
HdJHatBpfrzj1e6fWbXXEWldOwUta1wUjTtDuF87YM0+YdNnrCSEcV9XV3kl
EV+s4e4sFlqYwkJ6neYPhacXGf0gvq+q2ISBFwWc4R3zWMiwXuw+7KZsO2Ml
6I13orPePvJ9YDv40zFHgYnuLncTls3jYNpW3nNfmGiPth78CA3EBVkxcLux
iIbhVVQAFgJ/wNMgvfcAbeF8vI8O5DrfxthMHN4m3NdF3BnNMn60egxwCTPq
VdiXzUKoF3Ckz9qcYKZSX58qGDMjemh/k7GcBAVZqjYFoQtnu1AIylh6zaz/
kmn0AL/0z3a4k7tm0ETuvSGYNDcTWv1c/9XI634RYEtoMEJqlkbdKkBoYD+Y
pETYhWAjzpYJCT/kZg42O9qiqiEFmorSHkPOC5bBXV0EfMfyZeuI1dHPP9U+
HGcKal9KunmljK1uEXYW2dSkAiSR5Aeewo8V5CupisA7y3R5fibXzfpSN9IZ
297gmbW3R/7MtpPZpfU9b2JeqhRmFg0ZSFeghKWhKnwyEXJf6FO7TnpETMIc
B71CKvkmuvmky4LrgkTcWOUfw0DTSQMhqV5XoVq8I/z850rgpZej6pXdieIX
cnkIQ+3HUWSEU4utdpsaT9SQRuCw7FXIuBJvRwVUZluUvj1+CSErF7wSDi1E
DVFXlX5Iluuj7rkIHqtdvxo2b7da9Co1RPHQnsSl6VbjmUx/styTE/Qigp4Z
WSfgs79aLFE54/JwZ9WI0fES+fqhivtKS4/WrlU4NBxC7fmGDunwEndkzcaX
qBSOY4qJx0K8p+cFlaFop9PT+zrYihbZWyYymwoS4jkwqJYrxdXqotUG2kj+
qWQNnZkITmSxAh6VzHLchix6oYvfbKtip3fbfiEZbsiXAOWjJ18xLoA2EZ3S
zSovnVqP4UcgrTz5l4Ov1cH5p5U730wUtoJlX8hmRYLHPq3wGM4Gl7O2SztL
kZbLxu73y5nbqC96HWlx1+Zy68ydBhcS8xnZE3KptYTMSFAN5Zsf6AGtOIAr
8jv+15ZSbkjM0s/Oj5sk7PT9Dfnwab+a3MY98tIC+dEuowxqT3idRWLzVOEf
4PRvbGh1glg8Vgz5/AgV7Ua2CC4TpntIZmUKOzFMN4/ZEqFnOnYvdaRftGk2
L+UR/OKKHyts9HUB9xiMLEBt8mB+et42Lc3qahpiDw7HR7SvDcvBTrEtFN+2
M/supEhW8RzbPGarRiNiTWb1VhHJvOLPovJxXh6gzzfkObw8yBSVQBhngXnx
gxPKG5NwtBaBTc+nRppLPC4LsRIEf189NU61MrCGQ/bhxRYFD9pl5c4Toy8b
MqnaDKR3E6f0kLsbo13E+PfQ1RnwiZ91SRPb5eeFEpwiezJnSwzQlxg1VSOM
+qsXNm9Yp8d1JUV0JpCdPtqtSV7S0buW25qbQ+cS60HUtQA1nFjMA+gNvo96
VyMO78k7qxvyqEsF0MTpWLOi7TfDunue2Cj/NqfumucXf8uVCXC40vz7xqJy
MH6d9wNJU4iQ2RwkpIViVOrw+6hrrdXJmtbf6glnZK7NqfxjPHKo8fy42cqY
BhM8iTnqBdgNvjO3D8n3gK9vjdqfI5I+inn5rqHRcfLsbOrArVfpEJE/ssyf
SMgOlCSFeC3N/ejaQG/gU3Ky9tgLlXtZuj96GFISjvsp+nUL6LxsK1+Vv9tX
WtXU1I4eUd1CeVOBUVnHAupWiXfFM/z84gduIJGigmil/bqEPSPh8vlU30K+
xRvsvtHovJ0JjOvAiAffcYA5LCxJLMxwvJ893k8jm4ogHDBds7jPXz7iPxrZ
CfbHg5TDTXqLwDLDt0jyepjQlSiGDQU9GiRNMUxVBNuuYMBASz9nEPAroIxI
ACHl2i5xkt+Ydh+uPaefcri9iA40FZJt+0sDjYdeYVUQpKmgvqoRjHnrjA4p
GB7cHHgXE5uJKKFOWz7p3+pWdxjdYPKLIC7c19EsRBk1JsJn7ENPr9KMic/4
g2zmUY+GZi6WsfCppd6qu6FnjlSL1Q+QUUfeDWVQWZZGpMChpqS+ORp4wZfv
cmtNNgcKsUbCJ8K8nzXsKHBUErwKt1IzoHFOBBNvu0+mEMe/9vM6khbPq1w6
meLBRbyGdOkqiZ1rCR9UAaO0fFz2Yjc2jCh1/ByMks07T330Mdrpt26HGn1q
bqWNJh0QwzJyFBU6fVPqzv0XNke4H+xZFXPgnEWfEzpInVvFGZTYKsfJ9YRV
PrL7OB0Ll3fgXn2nSAfs2TqB84I3/7dyT19seiJMIeC6/nEQd9KDRx0FL/0a
NkY2jlTqyBTJGrGDEftszTzYLGJ02/LeYR9/V30i5F1c1A81OwoNIq32uZTM
8ghagYN0KhlAT5ZiUbzRMYDq4kKou1a8qZ1AZfSancozbsKm7gGB4/gNIzQ+
XNefOeSs8Q0oJDKvcR/GZADSi5yEL6Zqo1ESABtaryRi+/wvNMXAB/EaRS2o
jfbmWKjf0J7jAEGuTyEQ8p5ou0T4vvbqYbNHHen26VFzv7WP1Nf1qZav32AL
pkHFp3XTioCu8wCE/GxX0yHJV7ZlH3KmFVx+NpY/GGLkIH2loPu1xC9ya2MS
l603mXgP2/idiyZF7ULY9nVBt5I1q9/+CGaJilJw7RgFZqOA4q2T+H2drL2Q
Sjw0e1bnMA3Hr1ClhAWVBMtGQaN11ETHtF6mczQy7Fq/xkhitf81LSQtT9i7
yXpncQqo0H6t1hf7sjFjapY0vbfvX8XwStBCNax9ge61h0L83J9zwThpe93W
Yg/NsrqNUiEvFNXwHlq+z5OSD2Ho8rbz8stNwz2m6WdIWCcWgKHHCXc/ZA2R
RGScdlU05OtFSk3WEIXgFP/LP2YpPUiIZt0Id1w4OMQRTVYIH89ekFS0AW9J
l0/xnoV2G/pUyqXWWmurNusZoP34F7vs972IXvEaed9fMvMxMJtM18ZBfNqF
dJgVP48Gz28f92CMaKXitv2CWPQDuh2FDpvbKIxPKvaUCm4f4EpxTyHZom/9
1QluJov5IzvlSAZ/kbAizgYwgogBM1+klRSkZ+1gVsFkyi3P1q/VCQ2IEe+Q
jWcTRGsF2uGz3MsqXS6eKetXxg4PzwfM0WKZ1B2VTDOsCvTkoAkQiJULMdAd
LXBt8NC0eUDcdK4YrxmBuwpWy0u7LldFrnpNrAhlfOpD6w7QVwIsESh1E6pC
mWZl2WwQbZkJvKskBPgFmc3vmcii81DHp0fBaUYy7b0MUzB3jvyK+gWCmtBV
kRC5cz64ex0bdHNEJ8vARAKUhJWAv1MbhI+kdZlYU+N9D1Vjib5BNj69DSML
cgUOfWW9DOSxEfOvL6E5qo6bWHJE9T8u0mnbJ2CFV+czcbcj0GauqQRp5FJu
G09PrxFiUHi6MAdJhPUGNywUsUlzamzbcnjJiVbz4sttK2PJSeQwIA9yEK6x
a12EBunOt9Y7twUk68k623kr+0lTPTtUoVI4+dD3Lv2uyGQH45K6CFXMbHZC
dv7mGdL5jxB54ezVvbX/MbXWDLUlSbsG2uuFU8ODQeVa7C4sdHUbE3lJjwQe
Y/+nhjv6g0c7cIpOgDydnOTuvvEKBc12PccysAq7EpOXZ7BH/VxuPDlQnAx7
edc0GYNQ3Ge02wDHW/64KcbjDywlQMyw5YTibt8OiqIjNytXjhbqeve0lvhx
B6EMDHzpl15qqWSXHvTU6o8jwz24P1H4XUa2vgY3T7rygbSFK8wkmkOiKNgp
g7jdO4zqWFUnPUocgfn8hxlSqfjDHQ24YyqsN89d8YgDFZ9C0V4d8bJUA9Z7
/eXI3M7Mz5eE0dR11NrRv+HLY90l1WIhblXJl/QLd80S0HSyMWJM5vJsAdWj
+3yQiTi7wRKOqUAxnZyrjcc146xqWyFEgECuCdv+9U7zF9pUOjiAKFhPk048
igRsH8jOBlJD3BFE7WR8lnxr7T27HZjsXRnepVVLqgqbby2hIDFUHWlD/nlr
UH06EuF3lJ86GZudn13CPKJlPX37ko0zVCHkjEmH87xS3QmmJPPugSMZtL+8
Evlwa8oTTK42RM11V738Ubs4k2W5gxCMRw6Ocu1fqbPCbUCwD7cWgH3WvK+F
3PUFtU3j0Q0iWxkeng82cZWfCDmDZ2ahMwkesJsiGfrDRdNzdn/5lsOJsOWw
vVbYWda4Se1BZQUGHAlfIpnAAuv6Gu02FnEKZ7Xg7H1KeS9E6dFw9LUdmZqT
jPd1+5fHsXQtKjM2DydLPnYAMBodsNOku9XH6G9/JinnKIA83SYdREc6udhp
nVZ4TrZsq4TQzbjxThIvOvHaDm5JmzP//dZ6HUdd7XQqVt1JltHjvtPFPlue
48idGyoJPRBjGaDZurySmXRaVrpHaQyXa/RXINOcIbGoYZzajLeiSOuKvnki
Rjqj0/G5ekGzGqe++vS8k3EoiFwbXk3iadSaL8BLLDixw7HyRqEvCy3Jm5al
p0UDcrmRZ8Puz9vwmaU0GmX9+o4vTN78xe5x8WAOGu3iqHUDRSNGg7HokbeB
Ejnv3h49iV3c17lGdmMuiKeClrjplF6UOUJsZkhK/vznDHj4rdaPsc/rgW+z
5+DRnwgpiDR9GxrLvGEqyyLwOT1vhh5+1XzB3DNUroXkWJMfiN70na63BHPj
zuoTj6Gq7izcbyVFWoeZl1ttxvhRTGqhrr8gyK7ManzC7wmGrnQoFhgASKUI
NdGRp4BjX8IHzzPMPdQKco1PgEarU217pspo5x9QtAyhkJkGgPmu1IExt61Y
BomGr75fZQCGUQqhAr/JqmAYh+ljatr6gMU3Ugcyb/HvlYlzRPzWIHCmzdI6
x7Fe4Ax05oNpDQFAHjq1ID1wZ87eLyF9crw5ZaRT4TchwJ2FzWLXQQRCToPk
5i1KT1X84pP9C/2KVwrpA79hvdRWehgKUiv7q7P4zxcX3xv72o8IDY/h+QyE
eVLsG590C2a66P4FwY1QmqUHKNqokXBGyZcoyNk6gGTtaptVzkenTBYA7PdM
51hJ8gcR6gxIlgzW1hpYbgjWbqlYjMuEAPiVxDLRSjB1wTI9iephDU2Nbm/f
CTa2dhQGkZ5t0hYce995dh2N9YYhWlY5uEJ4ubvIM4PdgwsuuopnLlzFYPr+
Rhf6ZP9y0oEO4aWgxii7fQ8/UL4MkY0A/iXzgAbCQvpvOSOrltDvz9FXsORz
DsjhozMyqS1eTIRlIVuz6+chXkM6y7fUXO0/Aj1z4VWKPMEfoaWwa7vag0/e
S3FtCc3kdrCCrUAeFySn5egD552NwIFvEvXqlIGdNrIScOb9oYJ95a+NU5Dl
TrxMvGzXDM2J/Ua0ur4E5qu5r+XFK4+Bp3yYuXzAxuP9mwRBq4wwl0pPDMYd
snfVmFW89Fkqhsc8SjqLnxLaRCbyreDT9ho4k2bW4fDqAH6LYw5tCbvg3it5
GTkGvTOHUGn6ev9Zm3+jM7Yi7qQf5+WLOEU9ru/Xu9ywV1TKTzX1wHVPaZuC
CpXm9N8ys0XNpwJGi7nXfv81vlNUyyJuipgwM7FY1/h9pK8CY/ADWOYgP1SU
Qx8SgsF0kXfQ3QysDrBHHDfflhvns6GWA3yvZjldqgKQBmNpmEBCsBnTWpJI
qnJl890UrBufuYp8xCgnp4nQKiK85ngd5hsqoNsCzRzmwDvvM4mzcqa488hs
AC8sIfVqOd6a8MQ8obJHVkdokrjNQSIK99bU18WE/dw8dLw7EBdn2L4MkGzl
DnBO2FZeTY+ZnLkC2y6CA4QHSg63wizeAPg2RXVmi5qdN34b1zIAvqeA3qjL
SLPkJ1UxfUUVVuJqgG+4JUZ2019zgUE76PUSCTaFT70U3tiI1x1alrJgMlXF
Q/o895UcYZR+O+q1yh2xiIWbJuAqxjSk1mQuAdX9/cToEsdZjohKTi231dqH
xbgmjDrRL5fxC1cEMopKZlosW1mOfKCtnLqXfgCDpJzfxixyFH+xKt+nMThA
T71qZoOhC3iz+YSX1GT1ulcLObPfjHqoMfgE9L0Mmh7cpuN++XBG8egvKVmX
v7RLxVi6T5xiGlsr68cfw2wP81GUHpVxWYxQyEsJVTDhPpNOuEt4rE2z3C+K
DwlpsCRluTKNITKt3nAyH2j3+wneszCyzm6y7IQ9VzkH4QMpATFie6K1m8yw
IblZzlkyhod6HuahDkHAxgb4XNKKW7BFE6NHNN9Tm7ZRLuU3GDeo1PMjmrZI
Qg039Mql2qWg2JUYF4iqZQL+qA6KWTk5cL5r287Jh6/FyRXEGJNu1FJNs37N
EbHwzBmyl0MBUIYG2VFxLZKY3gLNFR5fuQtl9TxbEeOjB961/LmglEpeXQ7f
JzuY1YWeTzj1cUGG4diJZ2X27pNAUMKcRFs1gMvB/ZgS9EOnbWgTzEIp9i03
VCK6GM3mZ3zU/kRP7TnX07hb7t3gG8WSxRINF8EnK1piTz08HOLmNt9NWpTv
w8KplLW5J3MT8cOuLSY27U5kdnkBp0OP2fAKcAwdYHku2eZQOtNXyh5AsKt7
cPi4W1PhQKH9iNRvmprwL6EMBzpwi6vxfClDpcI0zACo93J8GKVZseRXWypA
dggtqUukueqiWxDqo4MAUYqwsH4Pq8Ouu7b5tekySTHlf7HpyHdIP5dp+ER/
BNnRWdukyow/eMH9T47b1l25J0bqtd5e9e8oQVX6s9/3sXFRirzkqVOwm85w
e6r59XXDRN4tN/YSYTBvwPMXTJgzXpvV/3QLRmQ0DPU7+7EM79tYGFSkKrIQ
69409Y6LhU8xJicegdDS5socSYrkQ3A1TV8yFqJcfXOAZ55Xk5j9ODgwJwVm
qDfQmEcth8uaCJTb2mF40w4yaKZ2ODhuBcXEPgRpeVRo1DJG4piIxIneonDM
kpYPwOKjPFlINtX0bap+5U6x8f3vBJ0IFje5J3ie4c5oCNtCwS7syGAhX1ee
W/tgBdVQP6IbwTiExeICUmMu+GZtOO08ZItsyEMSlc/MyTwghoGWH3Q5vTeK
KqHsre8Z8cYtvEmOPurkg2+x5mVJoCeyELZzJxuAfXfQ344cyPnxQIZHkgxi
IED3v5siZMgAjf9xrzdaTZsZwHoz6wd+qwSWDexM3HkqPainj7dijsQiJV8d
THn5K7krYOnq8o6YkcbZQ+dzp2fNcH0mrf9e8trsGbHVdUXaetG3Dpwey/nL
sMyhwnaAECxbxovq1oBJyCFCflNB7uw/jn5nsTF+2xhpkdEUM3KxnQVJxUK4
mF4hudyTCU0VOR1oUd5TnlLSscrFcOpoJKUtjFuot+dErQ0csq8rBadQB4FV
n1MUAKITFliuVjNhiX5Xqi8BSa7kDnvIAXtp2i6FENYB3LHyxy4vwCcDJQHp
XkhIdr6kk97lc9rCPO43iJ+AYYs6di/WHq+m0fm5o5XovJQqcloAdXd51JXn
eBpSrbfkQXvzxszsmGyFcTdpzcG1dzzFaAs3YtstWknesEBK10TYknbGDIkn
pn0iEQub0NxdE3L2dgIGH766z7H70x188EeEzF8bXo0W3RZTa3nKCjxzTvP7
awVpCg4Okw/Rz9th0khhhkHDqCQuzL9yMrZ4VC9mES7/ioClO0ez1/QOm6dm
moSr5k2IN8OmeYKLZXh/eFT+iXFKCCaFE4YCFZAM1qS6qLn6/ejRfM8Pn7lJ
lH7FQ5PX7IVOHrixblmrkQFeDCbPajqyguXc+DCo+4mREEMO3vrOOBbz1QPO
6czdCYVYOCFlL/573niwkZECAvKendoZNPFMxgCoEEuhAP/qa3KhUi1/9wVI
wHtS7EqnkIZqql3T4HC1eVLEYXquMZShYu8YyJOS6D+ecUmZmx8PyV9QHwgs
BJIElWamOiuBO9LpowAd+9JAEvFuwIxEBiQMvgVcFN2OUOU23xnduyKpp+6a
ke4UkzPQWGpY9GeIhXaHtLo+R+w+Ky/qbj/eTTPufymDItr3cCGIu+pAWLZ/
TpF8d0uNppGOnI8YkBYRgCJPhYAakenYkC+shRjtvhGrKewOtQWt1nZCF/Vf
fvTerxPwZNbdjPorjC745q/s4GrBhfGBL097nfxO9ZPJUdVDkWa+jwSOa4rR
OSJtaEUkS1pmaMtdY3u5rxLltYuEq3cVNOzRG8W0SEXj3Sm7MHhHBp3zAiRJ
fJObWJTgL65pcIkQ5MW/Rnwzix1TDMpLgAmoSutctGOJidtEE4mAOWF3BhGR
fTQzWXwPKQFR+xeethLsXJarKg8Jew6ON5rVQab6FkLIEe2p5ImjLfqGxkC8
v5kw86sXOWVow8fAx3WsJNoCeG+8DDdqSbzdD4ERw66kNMRRJwGzA6rKO+Gf
1cdBbf8sxFeEwPXrKAOJpG8X9j6GF07lomOQPQQXdBR6dXAcKvwVrc86Uiux
s+Br+1Js7TTqiOkJFpavT2FcW9a2OdR8dJobMz216Hw3OQAoyj8QpRZ7sP/C
QWTr3THA8daRdGNtBaoNDHBaXzprM8ypvHx0DNRmrz/NUyrHV5EFIZL1I+9e
2L4rME14yHmTyHsUoJwRpQK+EjEf7N3POO9ed/DpAPuO92LKMEOmwOFzxpls
5NPeYZSOsq9BtG8ZQ4qof6y3TmAHWO9JiYZctfeeNB4nAXUJeklGBMELDtgI
yiS6O86F3KkDL5fSw5kCUQlm+4TwPzM2usNx4qqw9Ggki6HudQVC+DW9UX78
Fe4aUq/BiYOAmnOjAURyLJF6KAnhch+DyJ0OV6ouC4QgeN3L4blgcyq9Kelg
03l42zvCWp1gU3bGXfsT0BfdLAlnA7+6JX84DLJ1U49Njt2w+zGdkOo4zoQR
zIWFrq8TRAEIvuKkChsPzZr8EKzozyHMFTX5/z584rniGPj2U4x7IiKU7MLa
BT+GgMwGpv3CKKugkxSOORvmKU4FC9jKRcz4BghpTF6w9ORHJsArmIfqZjbx
PP3b7vzL/ZCPr5Ssr8il+OheyUUMcnSsiqL2fV4KTRGt5bVkGp+a/scdH7Qb
n3PRSEyImI+alAhYv9QKRmEaovgIGh26yEZaxGTb2BkPbc7mC/KrnfoK+OrI
aX9970MBNz+bJqmk48uyY0Rb4Hlgd/SSrZjl4NA1Tpqi4n63exBvsvVWACeP
dDYRCXqrmnnHdXwp33sOSMQl2BR5NAOA7oU0eAs7GKUpz628STpwUQUe35bP
X5DDIQr9Z0GQdsWGUKFObyKEgvVY+47xbSLbQSINCirMXpaHpM+TOs3X/C6f
1A/ugQJv/BN9OqcSFWKWcqXBdFl+1IfpTL+HaFJl+9fzwpJWByZA5tWazcGV
iiyPruE3s/sCd33GLiVFJDbxa7zRKqrIRXvlTyZgx69qQF+QaFWkuSQAT2py
M4hqaklS1e02GJ5QTuEK+m/SR7HqYWNhbKlg1v/ONTlR3EboaegLnZgQ4bTP
7KsmqDHWhYGzbEXC6eCvhKnqHyAwAc7ocg4su3lWzCubR3JqSETKPkkKErI8
cj7R0CZe3XRP5ZTmwjM9NN+c1hwIY3/8pIJW0XDdEhOVRx8urNs64YnzvBpZ
9tmwp9KngeejwHor7rBkvQnyQve5yBth2pBDM3LsC9pPRpHcuhwkPvAzT2w4
w2MqF1DpU+LW9fBrBNii6aP5pwnv4dPDxjuq9A8W/WwzVzeXqQwiAgdGfeL9
YYNbODitajoJxQi8mUgZ7p2uHKELd0M4AqyDNLLA7LEeIsztI0VzXWmCms+N
+lVtQKYlaTpKYJ2SsGHanbC+KzdiS4FYundinsyrPe4qj8k+iBZ9q5uXveLK
UcIHQYeVl1WXYOTVXLimyyQ88GBQiQlqqW72ScTHLPXBrULt+A09oZqBh3wQ
FSKJmDe6HKbrPCXmGt3qPf6Bkm5bPSIFDcgNyW4LkcRdeAt4NGo62XXu20T5
lJHYses1pVnJcCqMxHTGljPOL6zYM7vLppvHGCNqCd87sCp+VIIIeE9iestF
NWEQdBLbkyXWuoIUf6GisLWPLnSQ/hXF4N0FJMAJags2e41p9rKi906dQ5Nr
n+99FOSy/X1MHA3YYalCYQVyhCd1qjm6cbZq3SPnJIPi7yJrnQ4rnNKC0Zpl
LKHUrMofflQAW/x9AB5sVrE0WErgoh4IaIrRwcFq+0rbrYNDFnjFhZ8XX7Ri
6yzVhLrrDbGA6/Fz7cN/fOYFJQYrGBnkGoP5TIUwARSh/QI/dWX97JKH9EF4
SftQpnXhH9XVRV1xeyHZTDF8CI97ElGxzsixu/JlyhvZdVpzeA/xN1oDtGU1
OA8c1DW1GgBuAUJLhpRa4eBQ0bCAMUZTgbTScB9ap52IRLt+D5mWYwpveppp
UImvcUxxGqbQkDeL9X/uaZ8evZ3isjvd92hnQ4Q4QU+MuGHkQSosck7QIOTE
jvA6+XYAIzmolGqla9dfyOHJjQcN5K0oMozyNzQRrUpxwfQVxTVvpfcydXoV
RdXlnPMRMrQsVNW/2wUtsjCFjqeTBQZKNvsVpK+1cT3RiTe2J9iWyWtR3nBF
4eqGDZ+uKHqfmKUfZzA6jtB45QapS7cg5s6a6TalV20T++oG6qOlrjP0W+Hp
f9tqGHNoZo/3cQaFjjS4JbcfsZdIs3uGNVXq/DwjElOt/clYLxlr7YrPdUiS
CrTs9/2qPhjglhEuU26cHEJBJSqqsNr55U9MREAPPwg33slVELVqOBNFQVfT
kOHYedaqi67CtkEK5aKLBljZwCdszW0CsEqZcvuQ/6MeG6A3r0x439XmR/eo
+ycuGD4kth9ZT277zrmz8dBZIjyrIMn2OY62cvBsvyUc2zd7kOdevVn9U3bH
peOjC50p1tC7LcFIk3KMU7ZUBj+UVhpX6uRBQJrQQ+l6x/hXNssXkUNbVrkB
0ACf4/uDoWXz+lMKskxEjVM2GDvoPYLCDlDzlNMTwNmrBlSmmbvys/RQlbqR
FIEr672PSNuHWf8kGd6tXUtsM1dSrr9YF0sTk/dwm9Gi+V8ED0osa8ZwvIOn
VM7D4L5OxJbRjdLXvhsB75OJ7f8Vtdlm5eCwWRZGPA270X9NnAVNzhdwTOaX
zYG/E2vG64IwYYwsRC1POVKxBR57XTg0MTZHmVeBfGoMakkdt4AH2bJTIyDC
XeVeRBH1z58dF3+yZie6PJfr8egAbSgf1mceVQIKfzjDFaIQypsC/RcevyKj
K2OoeUpAcAjGUdQK9egOBNnJUnIUyHmutrE8bUiEJSvV+0lWMhrbpnTtbgXz
haON9eghlcsIBh+3j08STaJiRLLuGESHmBK8XoJPTVxVDy4kUSmiC7IVGAF0
P9mNLyJfxhFtwYxxm7G+G+nIL5l9MwzNSQPgghas3Og+P12SCm1r6Y0N+9Bt
8zDlGExiE+mqKF1uHh4asTw6eCnPzf13szTyg3nEylgvkNW4W2VdluHOZgo7
SusVw5zLuo2zcRISElUoLtIC7A4FI5JmcsCHZA5fzGBGWUprDnFwi0hf/9KD
OijAo9NgdlRq+SDwchlpObmFe5ATyTCKQnZvgRRP0zQRFL/gJdDdZUd+zGgV
FpufxMdEDXk0pIfEj740qN3I08F6ETDVXxOU+y4iM1TC7N8vIE5FIKD7DOQy
4PHnaTV6O9Eb8aorT7IE9W0e5eEdrpPZg7ck2bWELKA4U5zWJ/agXTpzOqtk
njJsTVixcQaaS3yX6gekl/+pDS5b8hE5rH9gNiwgTApj6xshHoBayn8mzQB4
NQasBM88iqDZ7v5yQwjHrPwn1vz2gex/7wxDZkM+CsFlUqhoiIHRClDF9Tk6
RYDxO3DfKZcWPnp0m7YPr+dQLjRdJRFhGgFYNKpGWayhjsJ0ugoALoa2v25X
n1hEiq+gGVegN5OWbBPe4Q/ud0cvjdXfzVG02RwFvwIgufet5FqcmaNpEmRO
RCgEp7947Dp1XBr3YuuJ6OdpSoIW3RxmHKbzjkHx0nQsNJ83UKGCpStHn4hr
vNVLWHMM84+7KhZy4YMC6pjV+eVnjYY/NJPLmwt4cqlcdcEvIst0j7BsC3qB
JncKcN0K6Guq/0cvW8d1CKYIuYuHXlFngFPVnFTPeMp4asFCL0J7rN/l8m/F
DVmPVYKr0R+WgBT9auih2jv2X/aq90LVdcOKdG4KcBQ3yyxAoWo6cZ/ht8Ob
ZmM3ldhu51Cj4tTDqTouXCHbW/+kmG/V3I8RE2n7SzUeUhWgSjzOtIS8iSN+
zaF4CRlciAVoDS15oFqO1e1L2h4LaRiCyOWxzJmLtT7BUxfOVbBarmjbiCoV
qiA0oG9fyLgOIypxlH5BlWYxRahoFU5uG91dcSboka0qmmIrk+R3mreV8NPq
Sx5+qP3qyLGW9CIaykjO2+Hz9G39tCBf8rJ5gNt1tbxICiwq7BP8jcXUboxV
zjyx+cdLy7Hw8GF1J7fEeCNaVb310PHv+bvARnWg2/4Q+8IPSGNFkhoq4hu5
qzg9EZi+sFjSMRo5x8yToe488K1o2y/l/c8cEuNbKDdJGwz3FdIZC5hLt/39
lxGFqSJ/RO+bh3uzCVAded47TSUHhcskRbisV6D0yAejBpFfcCVmfjcEEoVP
VA15LYZ+9ri3EfRRZAPY1NVHhuerx50zsT0qnrrb0zPyg7RutxKwEtes+8Yf
7b+i+nE4EXD5TM9LoG7jEl4NSAD8rEG2bzyeqmI3vOON2mrR2IGyiTtVwDJp
pGwEehVXXJauA5cBoguh0zWMwGQnSreOfHCv31IzJISEwaTSJitpNUHBXUDF
2IYcToZg2GiD3WE34ZkGGIS+WfGZJdw1Ya5k5r+Gi1LunAtuvDzFE59oSkuY
yZP5Rjk8zd115J0HCsuS2rplueRGLhC8S3c6c7NXkL5lRGAEpyglbcNsBdtG
i36TCTqheuvkdajNGZdOjr1kaYaQQSzNBVlYEDJ0/jLKVjUzf+nfZsku7pyn
0gp7l8joU+ISdX85F5RQ20wVagsDXfwQsII0XAaiw1G3nt2+7Wozlk/7xJ6Z
SbDr/h3MB4C8yFjPb+d8SqZ0siiP7500N+cZdxXgzDZXK2eAf7kphCCsLnPc
86ezThjcmttx9IlO6vAC4fLwnY2t8tR1uhSR46WlDYUk7QfTqmJTySculeuE
S1LtMnaCTIKbYC7R0bCxEXAlxQwZqG8yNaejYezQzXvIqm/Yijro0NIxzjMa
aXhtxGA2+QMHhuCmP1Snd6QWul0BSi9lqzNexQ9bE/fSLrwLw0kHHnYsdVtv
jfpvFq/bpjnm7Jg6Jkodh6MZYx9dI29eCmTXFcjdtT2l5aX/AkQqV4l6bKDy
9vs2hT/p70jMWYd5sOsI3dD1PIgeq6B9iNJvwsuu+sKJ8IckZZdR57QSLi3p
VKReNODUtNpxxvPCWdG/hB0X22r3nojhRrduaKhDxHGLAsgMauc3xf074sbU
ueErPfPqV39PZIVgVSuMK1XufWIUIGvpOWKZcQXzKHonsOuTi/7SIV+Odrs4
66rLQwJ3FxKGhMUrGiIA7yYYjFnmap3ld3VPYlCJ49w9EzrN2wom6LGFLDJ7
gTo0v0exI9Hvx/O4sj27VCm25Rp/xpzd4b/k2Lv4JBfORbZN3PxAPiA0wK/L
kY4dG4HSPnV0mYHjVupeah1vZAKq6W6uLi+tIBtWvHpirD8eJj+onCgHVpJF
qWPZNSFofAgam5MIiUltt4lM8qj1O7NrzvCnK7XwdQgLX3qyn2KtNaMiWV8z
ApG6yGELER1gABpLl3TOoKoPobWGJmaBre598L7sJeAS6NtlhdT4t9kAS79m
ucD2fU0Z7352o3YnF6313n9dHNQYNXeKBfsww4EtPtY4VIYgT7PoRohiRl4c
46bsDEzk+dfZx6nyOKtXQ9ZW8uMUkp16D+1Rxy77mFg7GsWFbu7vfS56aZFl
0piQF+3pLAVR/grV6KRhDmZymXcCRrnFdq8C4+oadTshHGRraTyGTdyyFXEA
0DZGhFvxpGiR3IaH9ShAc0AvWaC5fnpRgQcS9WycYlKXRaRCykezQ5dKsGOP
BQAcOGewgg2J3usVz9B5L7ki0QVt1tkoTz7ByWm3whBFuV+1YfbL3qZIoMc+
A3fFDoyTpRDilTO+UXemH5ajdyC+o8h0vAeOWH3LJf6V4raN0TmC5eemlqIj
c27E4Ql6TXvXVnBIyeR/8wvfDFGrqjTVJ0q8jdOjf1j8wEFAjnzAowd9V+qc
88XbfDlJcgN6a0m3irqO8YpVYdnnsTGdlPx7wpvZgx8QJZZ2SPGTPZ9dxZ+Z
p2b9jbxd5UVAsHuQLJuOzn6Rd9pZoyoCw/rpB/pz9jqGL7ZVpNnos0W3ZRaR
hLpZr0aHAhYMD5MSsqXN9ApR8o8HKO5i4azNyI3Qcj2CkTws2qxzrYo6Avr0
U0XsfCCfuTw3ruulL1U8lW6w/3bP5JCzYOnV9kbCWWnJSq0oEMeFD6cKJy4P
fU8dPK8lBIwp06vsi1t/ijhmpyNrYGl2W3LMcfd00m4/92PGh2Q2OvDuND8u
nqpVbHFkeJqlD9wQWWMt7KGqasjrp56rRdK1W4tHrhaVbkR2hCsUhRSJ/kcB
kXGf9vS4q509eSlL7pWCOj/AAQLPxt244KNkFx54RZBXAlnM2mj+IYZqEh8Z
A+cTH+VnNP7OVTtyHSU8ajJoqiyR8L64gkTQFq148lQ/nmFHAXGjBbAyMiMn
ImzyyciinVi0PcwyLJ+xBiJhPTs6KMUBL9oLGNYQFS8Wb1ErLVroPf7VKSqo
T2faXegm/7NJgRb0jjPF48UuVFjA3h1S7SVRVvqTpuFOADhWivXge0jhbJDG
gEpls7B9yxVYRmnD2xelY0ea9Rc6HY5e8W+zVoRkS47fHOCSIORPppxLWIUO
K9ODlB5+E4CYFj7suLusgUBMvJ7phfpou7Qz1R0TNo6LDxeysOEufu/PnlYY
WJYKV8bAPmHxRTt7wick5nSB0iIR8GlQvkT2u6MJqj/uXkrelUkT57TZv6Az
slM+0hwOapNUJ+OBTeqeGOJuwjFGXncn914VIo8W8B3EWdblrD5kEC/qLOVO
61saIFZ0W8Fb8duIyOecaqh+gBGbnMpgj9ANE6iGTNu57C5VTxg+pCLvy5Hg
3ftyc30kojq7CvqAvvRtOG1kwM2NhX/VHO/62/aDKOdDICb5Axo+MJCgyU4a
2tAiaXvHNzBxHqPCgNE+VWszMJvS7aeMut8zG/4sWhP3/vgQfNah1tZ6JbL6
HjSN5sOyg0t7GXUtwnpgJ490lXUtaAzaxqFoAHB2eqrk/MMgB54FffT/59J5
qeFfE19CJ253b7lUZfN8Wj8P3iq6knGte6Dc2SBAb9leSjRRsnF1F76JojMJ
hxTSi90GRsEhMCtTv3LW4o4Ve/MYt/YTXHOp/3+fYkG0ig6zSxt7WsB/V66A
d2zb8OKPsMP6l55zysE4h9hfmuNV4GYIcug0deR8jTnGii5/oU/ZA9BZC5Yh
IztBqiYkop+j5PWMzVM4alpDEeiteJsVZ1T24ykRd9xgr5pz3Z8mVjuoXtUC
wjAuBFarcKEib9G0JPWGla8T7g8oCLrwIw2l0z0IdzFuqzi8rQqqKhuZ4HnL
XF73ddr8LF48QYrqzoP6SELbbkYz6xnJsYBP3sRxR8vhVjuDmz7PYtrY8R9a
N+CH7MnloPECTRRDROjmJYGL07LckuR2uBl0cIiJhGZS8b0GRWIGCy42sxsq
2GwH/6t8gFLwlm5fZs3HP31LyjCRwGe+jSW4ke4Hk7kdsOQlf94Hvo/oCELk
vkVa/TZwA05iEngQjHjYpg2D98Mt1tk56vOIEWlykNwShGK5RZJzqjN5L2cU
Y1frYNbnV1yTCqZ0tCiN9fx2siOPnaHb2gDfBuqsGSynTtbeDxC9YJKnDWah
gEZ4wU6xS0KJceyOxzlxSX9G43J0o3RLuxGPF2e1BWwS4g4zzDm1uD6YP0me
1ET218U/Pn0Q5CdqEjnIwzmCK6FnqIvL7xeD/kTjv0C5qvB4cZOUOCiMbeOk
Pw/emT9d7206l8meNUiGwuJmisDL75Hy9FMhDErq5enzaFoOcOByuANz55Pk
jKYyoghlEHHpCucY0TAisf3VMA/voIdjF5LaJ5BFXgIN6CAj07JU35J4WkDm
1QJhJQcVLZ+q/QcsG195UVCT1h0n6VzEVfV4uR0Khr+9zaQofXk/0Y/l1K7t
lGPUAN9V2yBkM/aUVrNwGDmemQ75uvAlQ173BgOqF4XqkWEkCuzXg/Ht6XR3
TmfYN9+lLZKHGQWU1YLzBRT+ayRTgeo4YYJvEbx6lIazlT6vgNvZm6BmOH5P
Ckuswyvs3m9hBXE+mXJ18XjkS84uAV8HzaXGc/BEtFV86wWi15yaWvJ8QTvx
Lzww3jAy81mmqnIWHbva7abi1LO3P8SlI+GfvQLjDKSblCoC7KogmrhRjCf5
2up7G86mSop0XJoRFKdX6YbcAomGExXHlYjAqU3ZSXYn7rqSsvq69Lao/iu0
zkhvoiorgtk2eFA//I+v0xFbMTRHw3XapB2Sshnj/S5T6WicmvXbN60kaCo8
1oIiTUAIzJfh/QA5e/dmkIG6KvQ4RiF+Ei87l8YEQMU4gD7Ve20xnOf9KKLT
657MNa+3mDwL/mYggSvALxIy+j8JEOJ5q2Pa7GZdjsnjIVqlwg+5j2SRt72Y
mmafxwgIJzTFY6yB+/7rlns37oFyUi7KJ8V2k4wZTwp6p9KnDIf3gg6eoMe7
kj+gdT/ASMADGwhjspqhF0WAiQp4gp+kQhFjKNHOVjjC9w690aG8tTGO5e5X
3z28BsArCF94PCHy02PBtLnOFCiUA7Igh6TH62A25r0ZFsFBwakmzdTIHrS9
JtW0aRfiPAYMGXom5UoPI42vDHA8lGUeNpDrEFDHsHtWVTCyhPbUpC3aQi2n
m0GrBDr+0EkH4DICYj8OTIIMgwhwe56x4zPB+V+Bk3BicSSGyuO+SHmRLxQs
kitp+LLHclSLyc8MTe3NIzDUjC939YNPqKJIO7yoDsuNZDbWXaMGAF292XA8
4HSmz3fKH205SbadUi032cBQCJLJaOCAtnhwXElKs3zPJhcJ4QHGNwB+jNt2
GoX41SYjZyK3zs2Qty6Y+x4azFeywEjAN7XZEkv3jrvxV4/Y7EV9xYMMLWGW
xYcaZZ2O3xjZDfTkn4Mg16ffV4HaeScvtRTB6UPDXDbZyaVSgjIqgz4RAvzw
xZX+Ljtk8yVTSMIJRBg6R3YCkH0HWn48+4fEJJbn8cYgkc8v2kk1wdrKuO0v
bRZT5qTKqQfx5pTZRM511ugO8D39eqNEKoWWbVj/UbZ6kZEvj9LoHH4QfZq6
bn/Ccm24NkGzhZY/A70K3eEtjIyQW6KThMzPoDtkLYphXw9IDJMVfOb+WSo3
mWW+NVhCXeC0aeYj3R3c3pV+gLtNRKBwfzNGmAEpzKNRNiGCN7hzv531uP6B
kAmzhW9gCfY1DFsEcE204hz9N4pJ1gVPcLDAwixvWj2/F68ayZo8HNEHDIij
TNXxTuxgb6aTrxLZWO7fqpCWM1u42desD7OcWEUoDftYhladP/vgIgiFWz/Q
uTddEqSbmSDKxa3+AlooxLVTF8DzE7cUjyuRTv6vfpAoAdNwlnxXYleGFcHc
Q2yFxsMOaJxtkz9vPK8Dnyq0MNaDwmE2ehdMBFAptXwfgU3wGKJHEXV9DlHc
jFkZNmXr3cZQeSWuJkvR4hW4LJEO77E+AEouMsRJARZ6JeAMR78GT8LlwAP4
HKK7whu36nJ9+Tew0+8HWLNwmVVY6G2YRZ9G71c1yTeTDdIq6aAAqcDJJZ2i
mqZ6WyC+gEnMP+uSzqwqFgFKRWQG+e5tHZUvlSxI36/8R38BmmWoD0ixbURD
Yuxl9c7BhZHbrIO7eURWhRUMqGRpO7Iwfx6WAIwdKwcFF9SwF6rWqQI+r9Lk
pY6hYq/jnsAOqc1bETeBr25W+nZeiIn72hhBSAzuhPTkqOz2NnUMhE4R6RgZ
kzXnV+Gwbs0i9ggNt82V4JwxEdm3PRY7+BiIIpAIsns4HAwzfyo31tidxXVA
4osn+Xre61flCnTwbCJMrMP0wDY1SuDAVczK4gpt4ALI9r/5bpN9bEwL8iFo
jtUoYh7bEojmyDu0tNJaIINLxVUzkq56E486L0OF10sHg1GttQULV1xyoXlE
kKSadgZqDuWpht34SgzddzwiKt6mUp/19wG/ZaSd0ppu2dQtGnLfvrTX9BP1
izt3usNG7hA2tGXIsVSevhJWPsXmCjjnNXYWANwLSTWYpDYnoH2pl0gcLoVP
nVu3oHUNbQPNJ1fTE2Kchw8WL4TIncaljAzr20BYsfDkRAzlmFYC5ue7qeyt
AT1ywUcyeqJ13hVkvP3p1LoQDRPXISVuLQak8hmNbvKnkZx02nf8pbCGFpgK
pSHbNnItsSEW3yjr96qY22lZfj1bwyhtOo+lH5MdR4btFZOKRJzqfMKeSWOn
RcZ34qUvoKy3EHCRWsFzbbJHaWBCBs+VCYIS9B/fzQi++KjFHsvcwwcKdj7K
swGp2qUc+Y3/2OzigrKOgJ1FxrNnW6pclVZeeZT1Lf0mavgIfgg11NZKT9jK
vE4BsN1ZBDxMksKu0KYeORfyv1rN/uj5MsPz+3lflugaZADZ54hYKcE7UQ7K
WcAjLfjOUuM4xwJ571H7wuZEs9OwYZN2681IE2NamNC3IwtklSN3lyeA/p3W
exQiyMJ+vmSIAstpqLcnxD+ZhzJ+CmPGkQLbmDKLSnPPkb9gINFNHn8fyCS/
GEur1s2clrtThhR/WQqHMClmc3ZWUBP93cBqAZMemPC+G43vUs7cfP+JIxdR
ZQuiB+3JzuaAByQmSOwMqo+i9mGoUMl8T2FRJTznQgyAVyFa/T0jrz1MeqAr
0u5DeGzhw+b2dcElGZ9uovSPewunsr6CtMnvFeGqqQdJRncXvgtQftKkfFU/
JGa71IKgImhyyKI2FeOisdom1vpC6IUaX6ydbOV3JGYh8P9+aiQAFVpnWsOK
p+rA6F4IFXsihkD1pLEmLuFkCPV37mPGn2MkoZ+RsGxtVynm6GYkQ1tcGMEY
0Fpvpx8B9AhCHW4hd71Te+2wBaqwFq2Dyxq8SAJhhXzC+pKD4Aba3lvmdDh3
PltlmsLqgJm90h6EzAPNZrLAzlpMFIIgbGmKHpCHntqC+W3wW/B7XrEIIE3A
F6alEOYbQE6Xee/5ZuwA/i++P/yNrmysFfZPSRuO96wwjBrtl1FQp2kVTlIt
aQs4iuO+i93g96LY4erpEj451Wvi8uBXYQKrMdkHP15RVmCm3+Z4DZTsUp5D
45BP1sID2JkaVcN5bLrrxnxwgMi+z9Bn/99K7dU+oj7pbQdpngdtMnotia0t
E7XG0kK0xop2VM2x42uHZCFHgsFKdt0j9PFQfQjKy4DLneCS/m7RdoEwTNXG
0jOG2rzMXAx0U8vxQs3HOOA4Sw89lkgWJ79MKi8jvf0MFB+czMkkJWl5djmy
ssF3Y12EVzLCWHJ1/xJcitnJ+9uUepAGF0FBB9Bqbenfk/tydTbklBEiOtK8
BgD4D+CVsi59SjtDb390a9343Z/PIostoYzNobG2z8XqFMoKXSxLQrzmo/OC
SeC9hdE3U6W/UpGCo/nCLXNPt8CNqNPlHoNhLcHwmcix9VP4rmQZ/+wqjmCp
3nKmopCk0DIGRiZ02XqUhceawsdVvT3q2oPAj2C/wWdbE2RFMRNgFB49bIdq
/GRJ1cf7TZ5UPQNPpalUQRZq7Az3WmCcDwPEJ7f+7rKftRHK3FVB5fHMcJgo
N8bC4HZt+piBYEVrzftR/wnvTTZ+8veindwgr++GHfkHyGXugqYzW0U8MdP4
8es4pWumJGWd+NeDvWber3rP8VrvQoQnaTWZOJJSW2lpJgdCOXaLlUPtiWLW
wiS47vOJZDC+BNHnUtLOA+HoUINsG/qQkaZsb8hujnSl91AqjV3ClJIs14za
D6RahimuChVH/CVl1Lzrkc8Q/tK0QAT0spJMunPCB7FpIs87hGjzynBmdroU
eJ7UH1sb//gL52CW4AcRsfxBsADSO6ziDLfkyVSRY3KI5tcKrNiThTGmqN3B
AT5pi40B6d0n2y8jpewXowl6jjm1gauDyvrECQ7+jCH0QL+gybm4R8T5VWKU
3TP2/JvMldUcS7iFvWDYSo+5XySbjR1cqkTiqGcRpeTl8oIwT9ylXVNPK30B
bOYi3jxAMJ+4I+0ZJzC2ZIAxk9zQFgAkd4+0z6LMP893asNskTC5mPXG7qxf
/ZTX7+bLRgVXVSE89X0oW7Ga6aRD3WHLfzcPkGHybQ+g9gLztpmO2izb0jTH
gNEtea0xaecQNDNvCemRlDA0V6j7Kp8fEvenYWJGrFlMh3ixFzrD3dsQmfNR
VO9HVm5M28tmQEjrPRuSxXWj5hdHVqGYA4m6Oa/i6uxt0ikx1fSV6AB6tSPc
lvAb4yXxR/XDCcS9QUi4VCxIp3kVkKpCqd86tpUrD7Bog5d6IY6sD6EF4BHo
Nn4wVzH3MQ/R02inI578upKlTYDpr818xbWrw46kON9uN40Mkk8//BdAvHht
ijOBwi/wcVWM9SvfzpPyAye8OOZaWbBPCNHJlp5Dk5QQfm4xnTBOjo23cODe
u7eErXKLDOCXy/CvMTWbOWsSIBGBVAjJne1h3txxnHgDBJZIbW7Tmeed6/Tv
Ib2zUHF0leNwyIZ4Y5QfV59KuixmP3psr0pDZER67wa3zOflbT2cr7f0tfX9
Bo/+mu2+Kq2CAMoAeCjuSGdbR1CisJjzWGS8EyUlDh3LEa1/OSsgwp9OAtIK
f/VEyCaHScdHS3CI5U/7Uc7AI52w+zabSu1CfFeuNxFp7KzrM+X3+lA9bPpP
tKR6STc71wi6JCiIrVzY/Jpe1rc7zXngaXbAIAd+7doXvKrRF089PTLzFDAO
qY+bjndTfd/ZrvRfX7RU9JpQ9eOCHFe/s3ZFNnBa5vFw5yaqqe18ET+r4Q+R
vayu2lBYKc+9N1CgApjxD1n6ooajUD75RrDSVdC9XzJR5Teo9jEeQ4r39qpa
CIuPUtbcbt1VoB04QozWlm3vVVwtjANhhnF+EMFe8Sj8b8K0rsEIyH6k5oOp
E1gcZ4LRJgIolBMWXuLKnTq2Mxh6dcXeqIdMM7ial0AGWAmS4TaKsFQQUD7E
HYW2dkl7KqMt+axJQoY3szzfE9HqdTMTB3Bl2uqugZuXFFPmx9+4lrzgAsg2
49+d7K4rpU37KnzEteQCfCv3+C5a8T03UIOoY+HLEUnkTrOZO2e/gj4tCQ7y
9a7vPwAwfLStLkyV52kE/lkm8fShknKDK261RtWeIxG7Oz9SKXd0MGITtATi
IWx2AZbNeJDMY8vvxi7HjyxQ9ui4g6B4YFAl9kOm3GWBPvardstwOMdJvm1n
Dfv1NkH7PpB2153Ig5gMeQmapHNLDzLLPFHswdCy4q1Y4HJR5PPR+Gei558+
771TCCtf4YsOL2ducLPNE8teCT9QWT+qYC0+CKQ/HcqTxFRzC3Wvr6pY3ITd
a4r7O++nwh4WfiGCkE/5P8iLceVGhUwCkRoQs2vm5eunZpEU9E169eyKH3SV
YDMGjrm4YY6fzoejAOO/h/H5saMJKNHDfpb+tDbV+28zGFfDEQwXmj75fXRQ
YSHgiEzNnjK18zT53paJl+K0R2gqN+c63P78gQz/zNFzVxfmEDNWve0siwom
DCjS/GOF7Kug+A4Rc/YVUyLycGI1EfpVeZOrc4D2ZszwPnTTdxJRD/NAz/jG
W/y2ruIcCZeej64XWRrYbLhH6ADtq4caERIVttZwprii14xUaO2hJWD/uce7
xOaAXitxmv/2QbPtXcjm68keCdiJPpk4pmMH+Zz7ejbI40ZXF4OKRQHZJVG0
F1Y79k2mS8UxkKvOz9G+paTM+8c1/5Hk0Y4s/0sV/2ezObT7X39EM4+I6YhF
YiqsVzJrseiBH9gr1OnNKb5ImYfXMIJjE90GrzEF0jlbxO4vZVV1bh1qZ/f9
P3LFAr8+xkaMJ/8KEITP891u5dU0jMmqjMcjhm5j8Aj2YXzHIaotmVxdIkEN
/eejWocvug1ZxxhiItfI4efaFenLAOldXIEghH4PFgg241w9Wgp5D+FIj19s
y49gRfm6JKSulwv4nZXYMp3U9kDKaJnQy0lyze5PKXxQlB5ZVd6n6hUIWOBU
+RDlU9+R5YI151Mmb2flOu8ahNkAHt777FjaeLyNKg2zpY6GAHtt4FBqVe3d
dxE0yhNZpQJP89hwVysIcRQdXeLtOaslFy2p3q4kb/AAXSgygppFbojgU1NQ
XNMyTNJEGwBH6GFuMJvkTDq/6ohE27oVo8MypfPIGZ+zobP+PCVHT1fYcPuz
082MPCG+uMhZIU7Iiz0MnWt5kXxUArfDUqDZZYmu6t9D9EcSVZlbwfyPJrsX
U7x1MQPx4vpJEuCWI2jTyIOX72dtT1/M8jmeMElTc9cf6dRNmsl25CxT04WU
74nC+rX9VPcGJ74hNPUYxuCeh2g3EfFybIO/HZz5ueurL2VO7rppGrXkdbQY
KQiyIvHvMpo5A9ROnqtJB6EPK+GwyFzuB72dRjAS/WRgXMXCBgnHh+nOl0AH
/vmg0whdnQTMFIZAo8BMLmncaN9ldg4gWMbxoqcDUDc3uucdTpdhqiBuM37Z
PfqNh3m4kjqUaPmJLm8opJtHZf9eHpybdkyDD7MvkrFymU9MYdblSXfT5O8I
NInofg2Mqz4YUTcVjRqhPbOPj5EbaHa/fHu3U/WcB4br1XOKz/A0Ix+7YSrE
2OM7VbrPLReoYkb9DGpFRUynEeypNXUFP2uU5W2fxGA6SyYpJZGtkxATMZNz
vifB072/2OmfNqvdjXCLY9v1Pa+xGA0L4xROUfQT/10EXGcg628145BTTZN+
Hk80Tk3YV8zfH6RUk1OJp98v1rFBl8kyMwaks3WIlaLqbN0Z+1cmaadogMwX
k9HG7Dz/5yIIr5HhHmV/xhactEsWak+ZToEVLxxcrTqUDvu6YRJB68hT/rEY
JJkjAw5qy31uCU4/qSMxwE45yoWEL1u6XYddJgulwaySlOgam/Tp9FNK07gj
wHMvPUuudLorN113fj1MIy6CVtgpym3VrU09CcDP09cxRgssbacXSWTWtl46
HeNpbF31Q0mLfjPz4PuzFPZIHZbsBfhbqoZJ9nCshK8+2LL3k5W0R6gV+5Eo
n6377L4rvfWqY7hiDn3xoUc5yrRTd3C8U/HslYmUcjrQTtvWoujDQrPczDQC
Py2lzcYtwzIWb7khnfGF6xadOSw3HWWRbwxrfaJOiYT9qsdKcDbP0AKkkfgp
nDycG3oGXqw8YrjRteeWB7rWDoecOrkCjutN4yGM8aDjphWQcV8eCXegV6c0
8MISR7ResPw//wwrcb7hkTOjKFJje8F22akY7IA47EZo89A1ShNTstVE56Ds
2EVTezANjvhAPBDC/2RLct52bbk7Pczl7O7mqmAFHk4uKtSBkSJWUdB3905I
wknXKqR9m+2XY+2ueu/JdijaHb+laKCjUrDuITk/80iZiaRgKqA/+mwvmJd3
Ac0c+GFwlnbAWwme9nI4ehUQwZuPlnAbi9WhMzgYr+2QLnZa7xNmvgwHZjiK
GtfonR9XhjDJ0mOULN2JdztXk+PSPPzG0CpevznkMA7LLOPgdysffZc3QcSl
A/r7w05aNwrjWt4SP0FribiKDpqcF6l14+StkL+tO9vcayqPbmDGcfKt5RfY
/F6vwQ3g7OGApTtbrjCRKDnJgm5P/bFgCdYjpBfrj8dySCgcgLAydxkgE1N+
dO+IdgTHRDYFH+jQ1v1iUX2KxlQS6vyY3UkoSRrozTiqSZ0iKyaC8E+8hHV7
aE/+WJXqZiX3oeMk+dGGjEw5AuQVbRNkdgSpB+egCs2tGXrNc8dI9cgtjsbx
wJLGscWtuM6AvQLalpDUh71ZWhwPsWmUlQb+EJJIh/tFijy4cFs1c9+bzC9C
o2DmdemMlPvJECg2rlFTdWswlq57OgEIH2JyWoKCtf/7dlDRrOC7MeS7vi1D
fUK38xX7gqOp10oJTZ9wFnVAkgEFtvzToYZDFKBDcjn+31aPRNnQX/i31hQg
D0ty1G45WokIfYx5JaGOPVW2OEoMCmHN86Q8+0p3kx53NB692ZJfjAavgoBP
vKlYUmH8DkZyKHc06ilWMJWkmqF9uTlDWkg9cIlF3GdYkUYvDvDb2lia94AP
lsRo+PJq362EcJzwMs8ZuuAD9R3HFyU9g5wBmu2bbNus0p5GK/733e2/ZXw2
9Wq3tYOt6Gtw1htvQNaH7eu4S1bnGDzy2HkQi3NNjEpHXd3V/i2vaKWH5ZBu
ZQkta//cg9NWO/DkOvp8FtMu9NAhQ1FuD1gT3vp9kUt4mm4oVWOeN6sWES6M
jSanFfIBsa5Fl9HQMYgeQEyS0RyTDFU/303g7n9Vk2pWYyL3NzX5IwKKO8++
9AiY+8eXaxxA0eLqnXXv1iFRCKtZMj9Pd8UGxSDEe/jb/rZn3u9y2a9KQfj5
U9WouhQAuuXopEIDrlVNom4cq8JDjO6gQTMnaBCNWl9+SnAshdzHUkCaX5km
WZphb9iL2nWpXzzW7ofNlRaP6YJENGV/5HnG058osplzp3GvhE0LG+ZWwbkB
OL6NLcy1Ky3ciyMTvarTmaI7w9h/GNTa/osXRjMbw7wL2T/4uG/f04ptFs7Y
e3jrEkO8/l16k6S3D9i0zLGVw55GYon21TbvnsnBfZAJnVKAPaZcu54Om3Y/
uQdjJJTo4urOIADgC/ggsCOz+gqpNH+tmGv0KdRnLFJGbGw4av9d3gHeioG8
DonGl86QVbjJJ9+OIfxkMJ5wweCb4ZNujgKj/moTzfNXv9YeoCvNqAqUD/Wc
gR7MJjp7dpBX5w/xAYWVEk6TRJrfovdhxUvzdetSv0lfuNLxbhOWLxdvv8FM
yeBi5+3jfl/aePmKAAjTXNTKNIV0+3+j9k7QoeA6bbYCOk5/aZzn8GB3Gtlt
KFkAgq6JY/DTuJ8ZgyUTZNJD+qKNtcR6orGzzZTery+0aQxiK+fWy5HOcoZd
aiek3C7UekTIxboIjc/LPVrNa3DG4FyuTEBx0I++Bj+mJXR1U+3I39ppF+0J
gmQgTugN/6gPwgTGwEY4W1Af4F2Bitx3MQyL4O8oPJILqxtWJNJ8dEJJCzbr
YHU/ntLTs/cWvufDryvYrJo19frSD+dlYl8j2XSlVScdjZYmotAwK1FxbJjO
2YZiClDW0Emkep9+mH7IG+xTaW+j898OIuCwbS0DSINB8JC/sPGTFjxLH3L9
aQoQWlDy5+o34hWr5EG3b2WEsaTYkEfxocRWigtHUUr7dgvaKHrZc9uvHzdK
FeLuBx10DiCVMo80N9Lwp5lp0hnbm5w2WOuAPkG+nuyzaU8nuTOPJ/ngX+Uy
gOBTtfPSd1yrKXoK2AdvgaV/ZpOKOpYmbe3f/s6qmRO3p9OmnDyIrtR9GbHy
p169r3OF78LPjJSPQ9Hd0mZCJTdZOwSiE6cJ5XJiCd7H0UKUus9tWuk0AJ54
rPAeBAuAOXQevczy07WRzZIjcfFuD6sGXSz/roghHHmkUeHEnEJQcdXilJgO
JXYcKWjYVCfvZyfNoAFaoMBWAK+gcHhNp+eI3movgUGpqbKCoHMu1rWnBa9b
VoLpRTGmjGCdQDxTU5DdZBtXPAzwFVaLxzNmGH79aligCe7+S3LGNIiQxcDJ
Soqv31B8441ozfl7/5hWnt6p90wNxFqJ0az3Ux9+QuH3YuPMK3pD9vI+sFqy
JoTmIcDsJd0401ND/UguFYmgzlDs898vLDfZ3nmiytS27dxDG+6znDBBZ7fd
ffsHueHdne13sZtHcC8t6/1a0b/zRFP1HvHld9rjQd1X2mBuuWlw/XVMoVXH
s9LteisdjIncVMVPnIA1wt9IMI78bqjTJQm+aSt35b3wCqxCArK0c7T2K8oA
s5Qa+XTCdj+/A1ndT0btAe5nM3+g+Q8Iq97UXAjfMYCbQTWMm/c1ll5PwZbk
wpoAZrkHYGfNufnJNRcEUbBQMqKVHYadqqQcSnb8AMwpxK8rbJP/9Q7OSYsW
3468pOoLm6d9AEFCyKuC3udhqQBdZPYITn+fnmrcK9/dziDUwEh/mAUkSWtO
Ms0X3C0EI5KLoxawpuGfLP0KmL5i6mp2LTMdu7qoTxtzl5dBXvaXMq6HuytV
8EHo9+N0Y5RkDSjk3/tUnDmUsS4M8g/wIOaia8FVbngxOnojXohK28OiX1dL
LziiZDMLrIbof6T6kmfV0/cKFiwmbiNTcUbczRDDJYBHXYxXDyXZowE/z162
QrsZSK4ReFQqmoQjOPuXYz+B6AZE34iAIB5/LcmgRjLps1+XjoU63IV8bgB1
jWFvNuKo6tTqs0HLpgd3H2bYNE5eV4oBJqpEEXf6anv7jyZCO/k/FaD6HfKV
yQeskH3pQ+oDq+fPBfqwKIAujyHdF6u8TSA6YQ3Bvx3674cYByNcAoITRUFd
Ed3kwca5mI/KIgQ1URVouaUmcleHTB/gXl810dcOJ9AdpG5wt5SK6UmKM/HL
GxzcwzvFhbGc+H6rKxQK3W8RY2f4uAqY3I1Db+nQJU3MWlv/jwIxDOQ2A76s
4XjWAzNGrhCWX2EA+k7SqjwuwmJs8WHmSe4B4WarHkti2FgXi75s0JtJ4QZQ
9lCtUXSumNPHHKLh4sDAf01rchQOn6y9j1Eye3JpY+4/ae6TylYPQpr0Vah9
xXVaQGO7QgukTFEKaMmT6HQo9/L+UYBKAv9KE0YiNYNRikGz4Y5v/bBiES6I
fytRgovF7bJgKNte44zrTRphytxx53bpeDo3aq9G5dH8JHIRS68y+48qjVcy
GjwhEImi+yYRe8HTdnCS/FQ01Zg9AJ2KdvwO9Tjq+VGudVqhKskW6JxjsPBE
d4CgQhOCR/ZW2er1/IovLE5SFgENNLbUYaCgnDdg/JITqhi+JQReabRkGMZn
lAbhAYI/zadN8RDt9DldA7MEZDPUhWNHKc5lqjVjw8XAxRgMiMxyHz6JySxp
WVr5wvsC4PC0Ti84Q4SoMgUCjGXgQgXj75s5gDTZnejjZ2W+ipzJT0b4CkfN
2lVxTz5Is3ZHeYHUHPVbvGbgwZhCDdK3kmuhG7twQNkjqviFq3PchDfxM99o
pDSJ9/5HoEttTfarV0qkdKvumRG3LkA+2Ao1Bvf2fb7wZGE1QvknV25dr7p5
ourA1yfRjb0UwwSBEO9VMVOKtPCq9dV+AM8CLwQF1Nj1hCmsjxGZgPfv0U46
vZEX4TtkQ6K6pwAc6rhRMav8WCd7jhfXRjgG1HebJRSW9zbueCF0WboLATVb
Rnv74dSZn/EtSRKEZf/nCxy9BMrmT3pK19sN4arOi4Yr6P3E1+tyeCBKqxrE
o9vwP6/ZC6rK+CHBjxewtV8jWePgzk3lbSOCMZNyha1U55iYCmkHbmW0m80L
dUelI3PeMHOeI6ipU9UwNA2HJLmE1ZZSghkF2ugdhXpZx+u2ubHE/CGaz9mZ
gE+YKXYgO2Ui0oUWkB+s6Mede7hehTdajlL84OleD93gR029ZeijuuZh7CBT
X5DBrCNoh6qL1qI7h43+AcHtnz6D6gmDf8Yw2u/NfOqjdWklQKewUhkWrFyQ
2JYiJCJzkg1yFYBCWIWE5x2eTu7bR7yYkBhmJKjpnOGbMa8YM+k4+EqAQgiG
/brRYfTu9d5Kv6pfVH5GRy+6sGH+ExtuxNqujTcQizGYq0TveEcmFrEh6Oar
r/HAxK2xuHrPYOYdwhfWAWD0u5PNpWcc6/YJ63wYryol6ThXvf99CaJOztqo
qIzcbVTxJcKZfK88/QAydISUYFK5HULYQFoG8aJcuKJh+v3dMZKSqJVKeEb0
wqVScS00Ieqeg36VU1xkclYvFjmaYtyFKd7LzGJGm4cRnKUvGR6D81QeO2Zr
pv76+ZCeJlWMVn6Pz4VgQ0WaWyzVmWsdg9Eu+oGSFFzjebxFV6nPfGi3PSyR
Ul8MICBwSRZh3DecFDZfUat98hJ771Ek3TAyFDLhfTWZLTpmY5zzTiHe+PgU
8eDRXQzQrg1EuRPB/mzgvRpbSZB9O73GkMF7JQzYhAH1BDWLup97I/7rF7pT
YvJ7AN/vITbmbdlmtTmCBIJv8kbMJjVGOZ9ikTzy7M5Q8jcP5YRg17H0sYoa
SjHwiyeZxPbzw3RnzbdleFiqp5wv212P2sbURYzNtebtZ8TOS5EcJ3zbYf8k
v6sjq8nnF52iq/GLBnSuDy1yDnVlOVhpHZbLX52ZFGLVhmyNLQj7SXcsUo4J
wY0oGBqsIbDOqE/D+qVDPZQmOeYBGnVAhba0EQ0Jglq48AwqWfHesXAL36QY
cl2S/UHbT8FZXiwnR4xZ+FqMFGLmzEN27ASLNgp8wiShvO3sgP6M2Krg4q3e
5t7/T3aF4Dqz9gGrglvRmr7rV/WiJUA+V1YZgHdLPMnPoc++w1sVS7PlRB+V
vxMzkNlrokiJNwS1JKS6sMYXeZvl38XOQoIIidWy3kugkvBkRxGRxGbGfuJe
xyoakw4ZhpLK7yKXzQbHKt1mZcaOOGbL6dQRF0yJWZ4Xef8/dlL3ovmrVyl7
ire/MJBtwXekgk+DfR36VEt962sbiftD/ewUKffYTUfsmEmndPfbpYCDoDf2
KyYdWx4TQETHpmyPxcII0vStY1ZuXcc14qHgIMu+Tqdb/tzmGYmuf+osmMvk
NPSNwh2GxfC6Gaxr2M9lguIRBFKqVPiZa0V6wTLwubwobSwHcLjqYbudDTNX
LyL8yhDeOGvEX2xvf1++hx5rDBR67E7iAnT84U18830TNNRVES+a5nqGVqSG
zNcJ/KnqsoQnCvYIZxePAVniX/5vnQguDd2j/KHQ1ZxF9mLLRECFAVfN5+43
m0CbVN97UYZFdLCrrznNwAh4S4yTSxkzIDeTJf/j/QytuRos0861DIKqQW2q
kr6St5w6TX4qWWBG6I7QeQxy5YMnE/LCXal8HPptnTEKY28u8+4gfKlBn3FI
PeQAudhh+hGuDPXEsHccZFE44Z74q+/1pO0ev0Ukb8uKhxapSN9IXsLQ7hMI
qAkV3OAlEz7jLMuHF9j4/NGgv5wUQ6tsjVFYdFKI6kSHyOFC4N/njW3qLmwn
cHUap7ij+ZCFj20/6NB+NyUgZ319GrkOf9RCq4PJPb3oW0ObQtX3/q5hanC8
Do5EmsqtKJShIVKrK+z/7MACd2X1iObJJdJ2Qo9CT18EgBnGrw0lpH4z00BA
RnwMp0Q9JUqOD6Sg4AdMLrhj9q8/Nm2AlUMfwUhB/0MSG/9WBLFTocyFJ4xU
NMFs652Ci8dtWd6n6OG/q6RwoJXol7Fhfmw7abgOnbezfStcusDsaCY25l4x
usdOBJQaLlgQML0EpJ1hfQcw6JYhOBuWaOZANYQz2xup6wSG2J+pxGOfwfHM
u/Q0E9bjFw89KAOyFAND6E/qrxKCsHFmNs5uq0EzOuYplkuv9aicbSefj99/
j30PrLzzdJkBkiWlx5cGHFV/6B1LV5LIih4HvWRmkgsw2NRCgMBD0k+2qB0H
7S9L8/4blg4JLkIcQNr04p5x+T+X+15Bs/FKm3nsvUD+4WdR+C+SPk5imY6/
GZ8oSuPhsepe7daAaugtF+oaNHXw2lul1Xrgnzx6kbx5RbO/2YfKJseV8JQx
l5xKcdNMhqd1jefbI5E4n7fPz1Rjr+1aSivto6TXbJNO9YquS+8JGHqGivmu
aTZYfGwWeKoNkZg1EqBRf3mTznx1ZKkDPezDqfB8xwof4ofKrfwOoioTaA/v
DLtsGdI4pZdF4M+BFXJsu92Mvr2XAZ1IZObxdk9/nC8i87go0LMvycd9yXkR
MVRLT3ZfYNM+GxRF4C83oG+YysB7QZ4QG2edqcAq+3T2YtrQG/S04ZBVpnzV
ugr0Eoglnguawc+OFEu7IJ4vKQ5e8PaUFPpVHyNcbNaGGBtkL1UVQ+F+t9av
iWFXz46PGOZTyHrTFngCwXAXXkz8OTC5EepNOqddG/TsCMkJFrJgi4pkuklM
ApGBCvXzR1wS1BFnZEMueO4U0HnXUwa1WjUR2LIsYWoQvF5h+YE9/2SWCPCd
vydmDgH1NNWuzIEdBcvGCQy44lZ30ZzYye+lU0XQoUnpjF0BSgXvANBEAGjY
2+Y4+zZwYvqK9wNKc9gUNNyyucsHRHSPAmOXmlfRPckG4WZfCRBtWmH4FOy6
Ah6th+7S6CaTCNoz09ipnAzSIfv174HUr4ir6WkVveVOyp/pocac2tbdn8qh
6okfoWdPBzFZLmyIrUKZ1z+BBOjITSB97297TGNwCRziHFe2ebGMr8nW8QVj
4V6nVE4NMJc1AdxuO/MekSDkV6dba/iVh+yRVgks7nqCtF7z+bvjbSGwcF/C
vipq36uHGKs4JMINN4nDH9dwn9WfRV2/lh3yZK/CuFYirHpAqwphznLpQdRj
OPpDiSeB6kSTNQsFXtgmsFxiNAwV8PHf/qfRqxYDQayUfakvxV+VIR8hOBNc
LUpo25tNa7rKPTVGmnn2GTCIDWFzFYWyo01ILdhpsDeMmDOyj26ZHJMrTfyU
Ebvz89v/57IjQ2N+DXwTQ7FW70FXkFS7OSzwy3tsPUQS1ifBKUEZSd88/jSR
RV6ULukvZuapyd5zh/uw/fUjlPHImogzsx45hk3FC4VSz5bVOpv9DzZysQjS
zFC4I1kk2ukriOGZqt0AEz56n83Xk6b9A+0X5ryGKyIw0izUIuf2bL7Zv13k
VGL5s2FVUNgjDapBP3GyvaJzR0x0IxzQisC5RqR+7oiC8SpVNYdiHySMbaPx
+2JVHbOJw3XJmJAgnyYPympqt1EdFJ4PlnLWsi2s47GgKwoGzejHi2PuSUbW
BpwMHYhNeJahbnqyyKaHu/TTh8f4OiT3MreUgMhyEIz7X91oeMfIC5Z9V8p/
RVlg8h4dxOpn3vEwVPFSbxGhhjt8AsZTPXJ3A9jdzN6HWq2xP3N0oypgZGgI
QmNcOThunb4X2LYIcyLx42TNl+YmiMf13tZZ70sXoGkhh55KWxN7eljfoYtI
So8L0n2+am8sMhJQ63GvlUcsL0GVy8zhiL3dRPR78G65Z+6NRGm9f5y4GfJw
rZc1PapLQBGz/42isrIm6Ns4BtSJezO56ggqvP3wDZVBYg70pHvDbsH9ettM
LRinqd0YNPtB0KmVMOJeH/i3Y66RFAypezPiwu3LmuOURHn82zvsdKqXI4Hp
HKLJpcCrk9pqQaWg/jswmxOeUwV9sSKjyo5v8iJHdAbJSbVPUnc/evG9LQMH
tuPZbl3m/do6SpsJ7ImF9byCje6o6SbRgg/ELvBinJRsSN4JetgZz5n4lRwP
hsm3c9SieLld2bZUqKf5uAxAX2OytWB4d8lnDd6VR0LESduxVJSfjxWz0klO
nzqEf7PmxQyWmYUAicQiQ7kigdytgXk8DvhCYHrjEE1aOsf8vE04ASapoHwR
0/rhUQwcM+dARADgEvZ4lPnK6fh/igvKki7pr13skJ5m0oTyb6C/+lFbXeWp
3uxp3JWPqtIWrk2NmdkPuG2H23lt85NPwsgcHXxYnhUOSkve3mjgYaLjFvMo
pLE7SnZnIDys5MtAJBJImMTHHVuLwhnXYIrC/k0FZRe4F9ktx3pVA/B/zf74
1SRN7pu827J3VOZk/5HXCjV4qt/d8YDSM52ETSc8322FrcFa1wmj/1caB5St
w2fsCbX0L4QnGZ9fvBARocC3PKMGZYxn6NOLwZrsiYFNyo9IfYOhzkxgV3BV
o2YhhkFGlGsVE79VO+vgVvTt0Je3rrUDulugppsfAZ4WVJdyLksiFj7pt2xS
sMcfA35d4uFwwC1vm5Nb5WFr86rg7NxGzdpt8/7ZbPjuzacN9K8szCMQWnOR
hZKQxsUTTXzECF7yXoLEY66bsOPMV+4U1VLp9CS+261PkX/fv/THz5JacGT2
BdGb4P9LxxHDy23UaKm60JQLxnDFbIDpmhjzgWOrz3gRyp+RbpBFL3pSmKgc
DcOTacawo4cFsDOX58QUR9jOYhXOncCj55Cv9/6875jyRN2ZNHmhjXJYcCBI
1AV6qYpfdNstkouEWt5vIJ5fzCD+qrTZyw6+0ciJ5nSNwD+Qny0UBczMpWUT
796e+yv1TpDhUMbgy7TZa2FaW581N6WDj593fF4+DQmQuIFVmUtKcv/dZvbA
WW+483XMMLEhArgFLOJV2GvRK++CLjM1a8BsuK28LooB+Hr8yNZj5rkt2i/R
+4NGyS6w3fnuAZlraBpOurZzGu5zXLNsvvH22YitJtV6c0cEI221GxOOEW2m
xXAFEABHTXTvI3uhXp2Mlty+WVxf91OY2ubZIvmn3GRg8oCEswwlGOv6Jvwd
+Fo2XNW7+KSwDAGz2mX/w+pzKsMZQWWxm+6/gSjsF5rISNa6l1eZC2CBUi1m
jZMYU2AUF0osWDTpyOKjmlkzRSFwzbxunnzo3qkUEClIsQmfSQyx3ARpj5E3
Hk4CLmKHkcsrymksp65R1hAAMEP12h/H3wQ/BFF2ueFNDQQsG+PPCMC69/II
jJB3L3FrrXbHLfIuiDZJw6u+za1jbTKWPNu6oRGD1Tckde1OWT0FyFkj6zqK
Uvpyz34wc/T99mojgnjgGp8k02EyVfP0+3iQT95/eacB9XgxE+dlpOE9AUFT
MB7T8Tq2a6JR4lzZD5fp57jIAbYqoC0hlLQeod5JiyJbI/vQiolqmjDy6hhm
PVQjh6Cou5fMyDdY7CoKfj/we+zD9bHDuYu1abj2cxOjzBzHDDNc2NSoM4iJ
pDchezdNgsSVUNIFGQZydGeW1KFl39tKiCiL3drylZPjZzs2b8VDUpff0Exz
U+t6c/pAqXt+DkeFEEfIaPBgO+IbgeJqq1U15og64Tsb5X0GSP32iMbImpRq
wHcQqfwdhXoHQA+gWNqHHYct0SU3bgh/DrVLsJ9LmDZmYgeouUtGU6rQaTFl
41PcrV82b2/bqtFAFxyLN79L0QaK+2PgkXEYU+f8QDAQBiiUBhd0BhSRYMFP
fsZyonZB/G9AvsGf3sqi23cBaZ+9eg40yxj8TETN4J8K3SbTLyujU0dnH3oA
buaC813WW/v06u0qr5Qvq/jq2XWafRvDjkhWaOeCnXNJ/OEy1v2cTPb+6ztH
pZ5BbWM2NZkAu8Uzjab2m4NI0jWTA2SGVDnwIa5V+ViBPkhRtN80i9vpNZ2a
EZ7pse+CE9jstF5Y7VHkIeGTIV4nDt5Pgkg7c9Gfhabi7GQsj5D00ipnp+hf
i49yM/39RSHtZvoR52ThZv8Ukdbgduic3WP6pcGIhvTicB6wScwXMEVDwiK7
sgurPo5yZ3FLDIq0GWPHJ8ZrLzkZby2YjvVidV6h8vhYoWbJ2qyTjR+XdhwS
oXWr6yy64eHjPFAv6jNE5qNLfMR29jzLqUMuTL6u9aJA59nmxDiMY7PAWaWA
GkVGHV6oK+1YSQsbSipO0p8I0MraVlHx9agoJidGn3BQSJpivfUTT5wb5BxC
WUH+c71o7FhQJ+8Tbb310fYauM1oUE/9oDjxuK6CiRTEBnpa4qMUwESlyiyR
ZpYNkRDndjqHq5PHb1F4WyubfrcUlysX2vpGwhbo55QB1t6vSCOyjeDmxDrk
yI1XGY/jHMzqTKzckK9Obu/skvcRLFa2wF0XUXoWBVnHxT84kDidD9xX93gW
dMTsSIOomykJahvcCwvciD8SDmg8rOizf49XRV55VHL16hh1a6Fk8RpNi1tn
OPflQakx5V91EW+zCvqmS2Speyu53FU05EseKwvO2nHyxUTwI0wfpEIjwYzw
xNu1sGrbgJHBMz5ak3wk7Nct6CZYH2ddxSCklWWBt90N0pHmoIChDZI6LI+1
n0t+nQR9Z+7SF2u994UPYIaJ8GmWPSk/DhAH3XgnpWTiH2M7qr7djo56Zu/L
4aVdyukIJnIATxBGhafByc0QLY0P52JjrS1XUQVF2/9z28CNhFuV0unKl6Ka
jF57OIREBnp9gVbtfqU3T3pNJxrBWmqKFRcaqC1cCmItn0tYpl7lxoZrXgMK
B0O3qncAfpW/MrbxjZLUl61EPyDivfeDDVKpg8U3wm0/JkA/7F3c7AQvRxYr
I4oAZ2zHnaBTPROzKhBqciszwLX1/WTF3nVzDA/xf93OQZcQtMpLs+Df/yB6
EibN9rB4JYv7FjPI8z62l5B6koblR6RyRdo006q/fhwYfZZnHiGIOtsyGvrq
pKH59GX6Gdcs2uddARTwWV3Nfgxw9068I55UUc607YWB/SlBBtIXUuVYf9rt
QK/De5suBfSuyAQgcaUvSzRb9nFbf5YPUfjRG6LS/qONirRWxKkqItCr4iKW
3bAAdNWnz4QFwqX//vwDg75tb7zCD+kFmtpZQTVDjFUvCGE4mzvmD9SnKFbX
+FNdnqavgQ5FStUcSn6NgLotwER7oBxOOMaee/qqxYUovohcOoRMImLaOLk1
ppGR+73jx5r1ZFe49endLp+fKFNDAj1uPNNVVkSRV+CvRdnadMEVWzzN5QpB
J/C2olyNVib5vsgkJ/cihHZijgGNENcFESpx7nPYNffbHF5QewFr/Fsz3KJM
SNyVz9EY8ZbCuVwBCRsXonRyCCY2TFgqNwEmIuMTHS3lEqOzFt48FJPhrTJ7
m9PLUJ2Fu9WpRcS0dsBkmQjhYIyU1jwxTMplxnerKHJq7SVk+BwkbyWWIn/s
nSH6LVRCkjlzIdUqPevjIJ3d1POlg/S8jZp4DV3kYx6YJadqDhuJxK6rziYs
4D41oI2jEe7x+vPKoWAI8mq4EmWdA4yR3VqGgcRW+eLVc71ynmp28Pl6EVNn
GdbfEanta/f2MwrjhtH0P1Y0gUleoA4U0sC/ies5uxQOg7n/jfvoLJm1LHj0
8gViEqphy5xxsuE3fqRVHePoVc20Wf5zRuOBdow+8sUXNKmXLCQMLClYUTLC
HmGFXiFEIDA475xj8P3Nu67yVQYlJYGXlOsjCVb5Xqz3f0vYCxvk11iKQris
DQkOjZuM6Wkg7RN86fiL23ckqxsjqzN6dU5yCjXZYraGJBybIN5C5cP7j7hS
U2g8GL/kpGxoZks7IAUYVuOveoHy/embfRS+/jkz8nUYR5JM62H2gcIfnDSb
BiECneVutTVuFrEzjSJ/CN2IIi28K5Ob/aWL+SAbuRZDF9vEhd/+hdeUwgYk
IR9OV3G5zB+Z0gG2XjakaHbJPsHIfytNtQGAq4ME7OHc+4iJh7ROp9QYnjGd
iniB8OpO8+DUFz6zxJ4SpQl1Y9NYpQzPHvCxaAOhv079lQVzE8DqqZILH2e3
/XQLBm+I+pJBYcK5hdkFlNBqBlQbGuprvhHhA1iJEOr6l8TjLTAHZtiHK+pu
64wROz3LQOVkvfbHWugBeNu93eTz2gb+/tWrUcruKqhQ2fJDRHAMNzqUiwMS
RwWx+uUvJwkgo4PbhV8NBNanHPiqlCAlVKS0jZMUJCMkI2fvxjIXOv925awJ
Qot0DSgBFfhxrBeDVZ/raS+kHipRxFydcMwEVVOxklZQTGzWlY2x9cy4ynqD
xEv5Jcax/Z/IgNRUEgNU2zPu7MFTjfg3KKp7jV2ysfM1gwLOUVgN45G7jSTV
X4dCeNX0yU4zWQBzQ8khi3gPe7fOG8STSTlt3NwCCIZOb3vS2ygH5I8UxU5G
Rj4y+mqmqinGF1iUNFz1T/q077g8C11PAq3gB3wfapznhMBnujotm9UEC3Jw
jKrPQf5j2pBepBEjzcoi4eupaKqelc0dbWIQgzKNNR0SNI9U5Q/9k6KzxBKg
rLnspzfmbpwHPeXIpacvlv1goyzv7tGWOVw8dTn2vb16T0UnQzb1HmtrRMoR
8p1XVWJZxlmQkhtvtC1cPplixbuououCSLYSvWWgg+GTsme3zRsbd3I0X+Z1
RO+ngSzVew+qBfZEfUPZo9ccMV/AFo3VM2V+R1y23qvDLOrqERQcBPrvm6Y2
0hU5HIIB34+hB4YhPuvfSdl0gCtrviZ1C90Evu1dgyDi3YBmG4emsBU491m6
b645KBDX1PYFydo3d2I+7iyqPwCOHXfjV58luMTkL6aH2kYfJirAQTC1aMXK
u+5uQtycPYzSFTnBEEovui4c65WuF33fK9xkf1j99t4GOi6A8T+hHMDTPKUE
l9Qe8k8qSTp0WypncbMd1Iw45ITFlFwZnl/m24ickAXIe4xTipNQf8I7jDrp
rSUhs+AiUbW3fyrVx5qzAEEEq5ge7ChcVy1hmLazK2R6L4l7r0yVwCohd+do
UA/iQmrhvkx7nRbmTRqVVXFE6QAd7S7l7+o0pe8f7iUoPFvtvM8QMWguOg53
+FIcexYgBTfE1bBXaiKpzEaWSJkqCCmUS2VKv3UEStADfZLoRjR8zQUYKIAb
TuSAjL8YmZJuJFxIruKB5Ev8qRybjfhqt9T5A/MFxTm32W55yGn8GK6z5hDo
7RQadAayozP03g7egrZlfGGY2c/NenQlV28WvXA+D08LQLGNYxereJqAxZjv
hy1MZbwx/IVwD6mmOUlXYNKD5BY/kVP9OMW+BX7zzuNJdaimIMZq95hWJFAZ
IZriHidrsiDanSO5A4c0GLWTf3Il/e6vR3UeKdtZ2JLllc0kkVv0Y/dsNta7
PGOnFy5aTfUMeZvTX1ldQG++G3jSpK8e7Nymf+QzMH0THDupJWv2UENQmBIl
cI9JSJobNDA46pj/a03BcHGvPPOZ0F3g5HCg8+WwvQH1EwNi0bv6zhx1vkda
4r9w0b+SeDpoDcTM6sqaJb9/kfvW+83QHBtPYIPIMEALhBrhgZFXgVMbOKNz
ts9ytButtWNqtwTRoETxKzdyPmfgOcHbl1aLvRaAlJreuprA2jdDNp9u5wc4
+mEDF//ljMzE9Wxk0+uOOJJIPeOWDYeG9qAiaNw5pk0RbKRvA8yrMsF2hdye
mZpIN6g1Qjw7pXYfJ6eO38VToI4aMchgjspr3HyukvGonuqInUbsQO8jOhqM
mKrz7NPqe3R5ZV7W4nixH+R9urQlZ8b+V/rA1pxxhCsiX7pX+U4ZhaUa8RuG
AaOl1QpGjbLo7ijLyhMZLESn5n2iQRfavQ6bmQ/UQcLyouPXDCV7qxEAVJh9
5YMBpmY4PTw0tHm/oxuzOP1tTFhNoj3UgS2LjWx5XsmSW1uOz907Njr4RE48
dk3zgb4/5HiolmxDR6MfAlAqgfaujd6NiGFhiryjc2yjujRLhlaVX+uupI8T
aiZx03vhhIctweHkxV2J5nf0+jRH3wozLvRk8eA9D1eC8no9KfluB87VwcCh
jhCIw4Q5y2YThVK63zLrXn/JQ07u4lMICiVA8ZB7gbKyvWIVS3NCIIqMOP9A
88LM0Qd6b5P/D4Gly8jHgVL2NGmq5DCOOnIrpg9N0UicVLrdLTQdP3WSwH5E
5gR4lzc5C5wiE+owoGd4Ye3JYY1bgYgq1pRZtNZfC0l1RaWEnwySSZxn6zCc
5b7g59idCL+gwFaeJmNwjoOysBTbmEr44Sb9xobEyFA/CmIxX0TsqJ9N6mGZ
3aHpOKSXazLbV+RnOEgmpmZkc5MgGCcuf+PBeO4YgJJCrnAAuga3bIVf0W3c
+i6Kvf3PeSizI0GtT0A5iNmrrP0yuW5U+lu4X/Kc6aB37fgd8shDgPH+KAWB
TFYeesjSqsmsNvCsGzSswYDoPZnc91U1kB9mN59FjFQOE+zGMcPLnIcpLvp5
aAghix/Vste5G2dSh6pjNFGGn2zCX2GfOtSMp0f6CEblZocgxzLVylR+Rnn8
O7fINVnRDvnkB3ufE8p9pKglXfrRoolLlN36AiUmnTSklsrnQZ6zsoEbGrXf
vmWwrVI5k4yOL0fpUXJ6eEfzKN8U2RX3a6AqLs77wcHDgTBiEsRGSRGjmCJX
0VBuB6Q7XfZc+mafnAaQmKY107vEX516Zu+uMWkiPU3NCr9rARh1dkK/NFC/
lyH3ql5b4VRBFYzO8LYHXqWarkCVFnUEMpt0Fh57pZE5219pFbLBeQvAHBry
pf0vKbTjoG6/5Xzoe63w69E5nmD6MTRWw3PAh6D+8sOS1guyLOhKkW1+9wzp
5WxFm5f2thI7ErbHAlD0F6g5i4LpTCxEZuAJ0r/biML2tYoVLg2Sqb0vwHS/
InBpHBOr0Y2cMT2sHCy7LSbA9x5Nt1xNeg6gyEiCMm+zBNWMMjyZqAdQZUHr
ve7zpwrw005QK1ms6m3vbO6XKS0y7q1E0+0p73gfnLRcjsuSWNl7VWJ+19af
SBpNQR8vt85DcPp0DQ1CxJuXIIAjDkNUkcQaoXjl21Ou51idvvYA+CYFMC4C
K/OFp+CiNVPJPcNJzo1+zMG5pYidI4mspAiW872E189Do+V/kEJhcbMwZLpp
F9vO4BDioQpOOvxtiX+caSMV08z02a/l534ksC5PQLU2V2MKr/qrGZWdMdFZ
Q/ttD/vF867/PDh0qaZoMhzs4XwAIfCD4A3ZLx5bmfnnAe0LHf2dQNH6wpw4
3BJ1IM3SPQvxf0mwZfcSmGT8uiMwERcitXuATGt+F6keQaj7pTPDeWR06zbA
+0O5B3VBK3v22xOcoQ0dKtrksAccT18LhKxUCZbNOGL08ODD508k9fEaMaqA
+iucpEC2PgSDEQzLERlFKMbej2vLQNaz7VZrEgS+Qb2PXZCgm27Y5+66gB/c
Ye8Tjdv7iyU/LOS1oPWf6qfQZpTIi6xmQahaAcwSIZQMMviP436c5BpcG3PS
1l3GuGBx4N5WIdaw6vCZfY0qW9D/Ixdb4+z2v5yLrAE/smdD0v3pXnMCxtA5
sDtxWp7S9/i4UXMMRec7XFY12k1zpNoP3DX6ZTHl0hrPaHIgKqIp2YLtS7Fs
HNAtdhfKln3WGZ+bYg8/JrwooIAd4Ze9Md1tNWeKw/yjd8dc/89uNnNNF+sI
E/+5cMfzKBrswwlPCX3ki2pdf67X+CDrU3+pI9CiG6VvqIKVc4q8sAORiu/H
DY9ZVAjU2cZwArAcDy3Zv0YKXU3CiTvRkUk924mgQ1J44LT32mjSWRbJxLSH
30litN3Q/7q/J6kJoWr0KV9raafOTanFRlNiOF5RIMImmFUN3bc1bYOZi/jU
p0+SjQWYrJpBJolab2sihkHePNDdmQaL3GWPLm2qO3xmbCQfHytdpAvejPXE
Stexmd0CHDqS6+sBeqAHqlwvjf7HoqYbNYkAdElIg9hf51UDa04IGOpqmfUv
g9v61c1pSm5pbV0UfIRnVfQhVxgmOXES8s4S9Q1ib18pb2d5n6jCZaE+jHDJ
E+qgeHs4r41A7gBfbFeXQa7+WvT1gtSjzRlO184iYo+qAxSTLJohFadIVBk+
K+HG9aZxv6zUaFJNJkUGCQ/HVR392Tmm74b8U5YwMcMLg721eiPf9n5rYxV+
S0Yr/p0ciZTFaXZGL4SQK63fbGBGPTqcR+9kWvm3yIOuKXfY8wK/EegzSX4V
WB17T+caPwZVIGuauPqDqMZbAYNmBhUWumFdfU0yaIUiBq1NBS4XH0qIdckT
hRcC6k5zdcjqtJh1dM0wsJQUe9DR4l5OztX7MhyuP9bo1diIL9/h+UgjUZ1K
Mp0FF6bu1UoHmfDRdwwuFlMazMAP36TiIv2ysrvYzCwrKkCGq+rUln/uJquq
yVrW7W4Xhotq414BbC2nq3eUY+fq08uX6wkmBRPGuG2MvEM5eCaDhB8JiWX/
hzSoc/v/99XSzwL1wBBYNcMhYqlKTeaQeHwn+mWaC+hc8Vcry/oc0fZSOjAz
gg+PEM6AzRjFdmMeDDPPQR9e32NNN49dE/2h3gUwDYdmlez6AROKOozbN1RU
Apv/xXITpLdfSIQD24u2deS82W0+JX/hzHlRqNl0RNPrd7k/uhpVSZMUVu/l
k2+pKk3TL8d/DU5enG60gBfQQDw4V+gXv5NkweRcfRbERZENu/PDFlTIYbXz
T5QlGLsGgMMDape70m73lbPqKPL1j5k7GM2paqYDTIKC3hwd8V+AinRxBr+Y
RTuQacTbndaiw+hsvgvBs2fjpT7cLtR/Iq6yRLj9rubBxi9O/LkegBn/cYkR
8O1slzyNCWcH9FAHJioXR7rOBJ4j27bxdK/1XDSUuNIGG7duKyAmutGVD39/
8pvWrXWazSnz8kbu/Kv6Dh/TuWethxYZdiJVHZPEc38cz/5etUBGNL1FdfB5
v4kPXkcgLk52q/HZOjQNO6y09HDH+VCksYwgoXvPS49msl0mweu0sgYbEaaF
kH1yMdlM+aGpOvSFpetNjyn5FXpahlGGNeKi/Hx+BkLYqMp/Nxz0kMXVUokn
NrhUGKV6YNXAVVlKuCPY3/k4xHqLJ/jZd4vhl18VyRr7OfUVDwTClSzMnafD
eqY1XkhROOS7hZqBcn+KzSFsKYRdNQwpfwe1kX8VF7Ws8JWQOgRaF7+Cemo2
NSo5YeMQMEZrX/ACrUPbTxDxyGU5Ju5I4wPm4MdCd29DEFp18Bq4G941w3Zn
ro4/jijf8Kt3nM3sPCsQLTEw1mPd6OibWh15ROaZMlGJFLa7HDcOpDxZYKA9
9nXfFJu/n4zNOgCvk/CqKxoHOB0Ro41gom7ZkzSXi0xWU3IUSvSkqds5K66N
0YGJM8MEY69f5BfubrOsfEZU1RDC/z4jNig0qb1WDLeKrtrI5kbscl3guuL9
6HQxU6cDBngMcbfeGY0TuJVow3gHJjbjs327jcRaItLyYUDTgGgOnBIGZPSK
smmosi8RXqsmZCEQp7hxy973AmpmcuIp3vyDh6tHzaojN64HwysGzcg/W42D
B1aMAJ9aCekEjD0uIgWzpiQ6l+TtbKUa0uAk5diNyTcBMZS70AVxICqrdfHl
IZemvzLvkcPSZrWIW0NvlUpf9pEWc8G05xgDum65GgeBimLooeOO+IYIrvLf
c7su73FauB8PCTbk4soad3rViFhGfaupNlEwNUkedoL8hdmrQdMBsYf9P4V6
6SvrBNzRc/EEb1EZrsOWP4/BtswYBqVxk8zUsmPh0RNdTUovN/swog4UxDBl
aV44nubSqHv/2noTRE2OidQcDdk1eLlXbFZcnWNjFC8Gu9Jy+v53q6z16u0v
GLY2bTzr23mrWV58+veM348uDYe8i2pcvq8w/7Grd0AFEQozRRTJKTWoV2ud
qU+PdrIXWaDI82gsvMUYd0JU39HfTglg6m3+IRzir2z1RolX6YxeK5YyIgX5
LnrRsDYw+rF6gVy+17ZKi2SNCPO0rfe+8Jb8MZkoWId6IEbzSsCiLazJu8re
xpOnGnPo3d8VJyR/m6iW42nokKXk9Bt+mPe5t+sF268ueq8UhXqbye2gx0fl
yszQjpbkdJDbBRnqFE9OXurZiFZBUZ5gr3F+/mpEe93gR/hzoEotEEOrDx4t
lC0kc6I3H5EsAXUymanprn3G6ZMXjAuBSK2x7LiJuBodTyjU+dAbBkmHyQzt
naXXHk+lOgEwAtmUpc2Cf072+WFXdtBBNPbeE65ib6sfjcKLeDGuflnY67II
8nfHOFGHYXjSHwrN4m642wU9XJPZOTksiNVHBWrH3UC2XTxDAZO4o7xKQCJ6
cZ/HTuQKML/3uGtoVTE9JjfGee1B0ypg/P2wP/CtHkrgU0Ybqg6miqJkpB98
M3asWC/PSC8FLoexmPU02L3CZX9ubNv2iE1Ibf0OvlCMfCP/odz8d/Wx0tV5
/u073+VW6tARjwsYtWE539fCuliaAKvXa3DF3L5jrURPxWF/8v5ij2Cvn7dC
v2BK4E0huZ4cOV20wO5oAsSufRVuTC+R0YGQGViZJ6lPBQCA3vIaawHiGodi
qGIHuan4hdmZYXfxT/y7K1ccmCwiMIisgif57LMXZi/QAJ5qZSjg+wnXJIv2
yHZRZnBzLqQTBTGQnHnKkjviWg5WeENYDbhFQiUjUXeqJU+Ond1DOA58NBaj
tYGWIu7dUgSWdI20GAZy6sTh+y24yQGk5+bEpEkZj/pUtbo4SZ2A3oCxSPr/
2g3rMY0AiIXivA4kciCKnhUe81aefvRiEkuE+BHSimCuTmg/su3vVJT1yfkS
OG3CbKCg33QUKukQswwI4Vsz0D5styUri8uw0hbE+JW5IpAWZWGPpQX5mIq5
N3MnI6VcEcgO8A7FpvV2R15x0UkD4ajTLomd/XyhEYOP6WjpbJ3/ihtDT3bN
wfK3wXWRgeuj3uCdmMP8lEoVl2ZaFWeLhPa721xip3Moo4iIk1ukqqNMpehO
g31OvHmHtSBW1edDROAwx2ibokpnQvx/3U4IMuN/Df72ScXphxv+rHq7HlZS
evysLdCsEY7y94/EXIW+bV0Cac0uC7/V89EfeTQy47Qkt+6M6iOwCcdaK6bA
ONLMs0hVJDU5ZYT+rSUake1co8wvTpxict5WGZHmoODlF9qgeXDwddsJBm7W
PF/yeoNkarQiK8uvVNZyPbrCupb+7rRcevG4L227gDF8+hmkB0DxDImOW/5+
m+CYZ3+310wSLijzJOInGlJ9AN6xa/bUPrGCova9gLz9CHYyxfRebNBzqZ4y
b9JuZFM/rYBbuVFZSFfbrql0UXB6c8BSNppsDiiaEx41GaznRs5+3Lq48txY
8COWU3KIFFBy1JJKKlDXP7GkunfH85rACZZN9ZXUw8uq7pqVtctHfpKx3gna
p9EEKiVPtBpgtWilIQAYlv2yQHq/gycSh6VXoVWKALzgaGX28gBSx1bLg7X+
vi10LtnCgVxQmSec+B4MEobBY/Q4mfw26qEGEqglnPG8839SIhrBQmOUsMJN
ddZFqhd2Ic/P5EiAM93yTLkHKZxULg8J88iKbJDeoka/MSXB4rwWDwPSUaI+
Waq/fw9CliOLFkg+ttLPdzTMW7uKZrlhzmAHt3D5O9igJbAVjH7Ct0oMkatt
jv8B8pt9D2PBs84WvmbfhsX5mFGaTLzTIP/4Gna7QzZTIOidg4v0T4QwJ54E
b4J+GqdOA3n7xTPGtdsbuEN3BT+f25QN5rDz227YYQL/D5vtA5ZQ5FFull33
BdlSbG1Gn8FlTz601Y31BTdyMZ6p3HMQmhKHzPQMX/V1D0ejB7joxLLvHZxc
fQYhq/YtOtu1zWtlOxV0RmWFtOVfJJ7yNozS4Yu6FfcFBoDa4XrXavkSXRWb
ptR7tKjSvWEyUeZFWUMhCc+oyzGI2+guUU16mZfGn+3/GWQDPSuaJNQpslaw
lNzLbibAPoa7b045mocuL/K4sBkj9dFbaEx+6+Dkv63UyVDXNgs4Ywm/DbKx
5b06i/x40A0hE9WZ3/gzOJs2rOud3b5z4rd59E5eU0uIyBRDiljW9bW+Y91X
1mdul0yVD06KpSF3PlCCFMMsKToZyiV7S8LDkE8s39Dj4G+SbHvR2iBVT0ZI
gjVMuL9YtXpUgemYF1Mo7z1Ve29JWVENydqZa3BAoiGbYt985v0e99moiVS4
WKzGy5MLhJOClqwYvwqwxkhK+Y2UUNRWE5UJX+6FfEQqShDr3PsWvbhruRpg
qxVEc4dyCC2HKucwC+JTzLvkPFPe+j01kVelF+F/16fn2GVPNQ8VcZz3zeEP
ywcQZlHwjm6hBN02rwyQ8Umm1/OYBXpG8JugQUFb+ae0uL8CG1eYcogineoq
+Aao4D849BS05dpJkgV+ONkPyqNloGERj5G+Y3zMdzku1MvurOKI7wal1z2t
VCJ1K/9vRAE8U8hXxLlaBphUvGE7XV6LxQj3OXlEXY0cJ99i8tarIFhKNpej
MlP+W+wlSsI/Asr5n562BlEZB3gWczuIFcln99k1NoxkiNc6nGsf23hDUvNz
v4Ja2mYholEMCRseZXhCQlmNmrkHlVQRpwuApEbWLvU67S3Zwo9nWv79Ry5o
ZwCQPY1muX4tnco44m6HJSgWssc61MrYpgAq8qe9/fjy9N7WR+etZTfkwQaF
tMSBuEwPBteBLXeB6ySLK1Ou53LW86phPM1hq/eMsjY3KcAZCKGiIiXG2hcS
S78+X1Gma5cPMFq8uOmMSFHjtPz57aG50ledOFcZXdw57ztRs4Yeqyt/WWIQ
0pSj9RHfKLntbu3KEAo/KX02qqT7Ih4hjL45PqTfZ+6W0Rz0eDg0kvtItkQB
O4ABfUD5WvaPuAKdvAgAayzVMqq9KOqVnbGLnMjc6kOUK05e4kZVisjGZSbl
S/V4/WPMZ+pOVLbolJVl35chj9PIl8B4RZa90H/ISqnSt8NlMNGq/ZfKxVwK
QuM/5E9rhxOblQQdlUFGNUZTYTJFKz8EFzwfEBz+lOWOVWwbvs+1R4B0Rkvq
ttRQfjcEz+NuI8mWhYdJzZ4lz6/pEotZg1JCOP0VBTGstj8Os1nAwKusY9AA
vc6ncVLe01HNlDpauvtmKdrY4RErKXttEwfk3Gm/+gzqwxxKyExm+oLPVbTe
lLPI+cxTHzi/9PnhEQZIuTMSpmQgejNPzy5+VfnSt5cT3Rhm7Mf/ICqL+wSe
MwvOHlHRl1dErSRq3mIiMzXpq2KuBBN6uXalRKUt7NoCbSYMBRkL/VX357aD
Ml3HQjY7oJY//lsTZ+oRGGcDKMvGcKvZ7mszZPmnxUA579YXVfceWkNZSH5H
0mccQogmP+yHmYq2rCC96TDUIrW5cZCf+rsEaJnoI21nxkuwTNuZEXvYmnC9
txnF/ZqpIlJjtFYQEkCKytQP02P0xONeKeWv6cPoiifADcMfIsOCTmkR36+h
M/0O3iXDS6mI25vwzar43KoOmsS2Mdsv1Kl8SkOXGkmxWftC5jZn4dVvbWMf
UhrRQDlk/TCNDAFoHQ1lmGrnDbK0TD/wh9V7CQKfyR8HsuT+j9FAnyCsoWaf
Pn1mX+W6MgQFTTDGFu29mDeaShHqIItv0iT5ttGTKbGePF2iSNY88UCVVN+S
AZrpLjQTJfeJCIsYyit/RAiSeut0de3cYG5u7QuJLpYnJ2lCu2WfbkyEORq4
4GMmeMnWRwBYd0oAG8F0tVsJNiOL72s0VxPjlN0VgF96vS9Ou0A3CqDs0zkl
DjiP+I225VuiK0xC8itwXpiTQ1wDMpKcYUE0euSnLpJRMej4JygHpg8CvEpb
ng0c7PMbAnroz/OUbZKEzeuhwlAZXndy2jtRNvrbb2ub/B/KyzsT+xQ9Qu8s
p8JeJR74qAxvEYWTTP4OrNXHw7/GzG80GKWHwAQbFwGWrXkzt2yfPsBExuqV
dqzNPrOnKtoi3Ld2RcsOkzls5VmxF2p+uyRb4olupJu/q9OLrBYTAzG4e3ny
lfYy7S5HWXAxqmVo7ABUJ1i0NcsBZ7h3rUD9EKBxIzI661laNrP7gt84EzpY
+vtHT6toeXFroQeifxBgEUNw7pLFS98YEe1n9qDuApQ5Vt6e6fpNmKBSw4Zd
5mLrVwWdQx3z+WPV+oD5OwMS5+ll5fzshxmZdZ06fIyu8E7AAQYMloZAlqYk
dDaLgN5AcqT9PMOOXJfSuzwGcCx5N6TbH3sZI0sbKzelNvp4sriRM2TFTBpJ
p/uVP0rs+nE5OFNINzdpV4eIoa9CKNMmOhx3XXfQ91tPaJXsbjpsBInfe8T8
HNyZuAr5xihmG6NQf6RCZsxmdCDzFqiTTWdP0UgPBzFFNok9QD5jEvAOJTta
JWFNhbfU5v4vYvTVI3EASdcgrUDukUHASv72T/c61wIQTeBg03YQAXZySHRM
OvqOqKPKWqh2BPmqp/TgeJXELPtPFIZePsg44F6VucJY3osIEgZalJ6Z313a
CQ1CvpPZFCoUdxcvysDyyL66Os1q/oolxQexPSW+Mac5RdaLBEeEYrip9Fnc
NsIPFYWaOKCnnKVniIzuoZLp2Nmw/+OEG79IaMTXyEJ2ufozbifg2seFZQVN
5vDy1BltYHcU4XMDjemcBi0C+X82xzpSQoywng6/05A55Bhmu66vK2F1lwSU
y5/zAdWBSDDoG6Vt6XnY7jB3yBIOUy28I0bSZEN0qrYBultSDY6SutifedCn
q+hnTdzgW+LDbluvYKJfTme1/xkjfyg8cpmkyBDXMmolbDvrt/qYVjWb6pe+
Gr0ukV9D4kYD9uCEhBDQ0+6pBr93VyIxTwQRhv/utsR+NVN7Vk8rOqYeOu5C
RddjLeY5wvMXoI9oSZTXXyDBWB6PiKyXC6QOjDE2nSm6g6neHvJHI60zeDSr
6qLBYna1tNQxvJvS2epWs0CEdbQjZ9iMnxdI/MThgraVnp87QKSLDBnnniKo
oA/+UbobG6N+hLed+VfeejxlirkzFNHSe0G5wZhl/RsJsFUGbra/yM8CgVot
CJuD5pXdJkXcUstxgZ3Vfr1kVRp11CCKshxjeLhLTZPGLKnYcCPcM9/KZPM7
I5xeWxMWOVbGQI5l3ruqIdeexRu7z6t8Q47/IglutISECaihnk8eLEo7fpEb
ewikW85cmuUHQqSZPx3xLq2nkNoIITJxF74LnEiiLWySwQbbTbqyeJaySobd
ZYJLquqI9XKKKAu5J73qrnFwdPviiqmhkY31jkjK1T3OQgkQUVNuzdAhU4yK
Ng0Gv5BeXsZxgbGbGqXneSkKKNpcBEDpmGBUBHSUUnkDaUTuXB6TRjoOnfeT
vCz8+vvvzofxxwJzXsif3xpvKyhGpzb6Sg3Lffg1jnGk+l74JX8kSqd00wZ/
UGAEozkLr2otSZ+4Q9oykmO1ZSBG6A7CLDHwqPn4oh+EZCGO2tVoy38d9Rv/
bt0VSjFppQ567etzsT5v06LnfeQS1/7FVZ2GNv86sB/fjmSyvONTXecC6qmA
jAs2KJfO4HY7ZyAaxcfGTVdXNukRZOz8bcqR0o1G0BU8KGI308daxpLWOYOI
xtUUi9RoRQaBJ07BKxjz9VzHW6D7KAW6PKXDkcE0URqd11rSdk6lSa8LHMxT
BiVjMbBnhsdJ35NV5B+wip8yVZLtwnrW6+1j/Aosqp9MaFZ9KVAG1a/8Qu91
NuYZRzDLPmuhhB635aKf7+/IjLZt5E4w2MLI65ZQ7Yw2Ti6j6a2zvbBSbBRv
uhbLfsSbMZJOFPg1rUQEDoqdwKghgEyTBCUo7K4pE4DP7vJqoKYP/YyAm5Ba
zqX31dEp5FyMP/mPnQ1/Lj4PTAiP+V5TQXiOhduLWBh/yVGUMJMiL+KRa1P9
BdsiM1wrjWSwfoAYJei8RPjNZnjsYl3SD9MYVofY8anHPljzRRNUABce5AJN
kuT1XVrefWy+kPB+KooQ1FLTvDeGVroUbHUzfr4f8qg+78KPBQY4gYLf2Pcw
tqin5R055LLkU3a5fBQg1kRCg3Jo4DU+W5kDZ7aU6FxsfPcTrelXBPET+F8v
ecUCXpjvoE09hFBqyAxpwLWxyZcOPUfD4e+DE+ZKy5VfdMh64eaCZ4OkFVbc
XsjnEcLLq2B+7Xopu/6RZHtn545ZG5TGh1dTNTO+xZqFvH9LnKVeOdtZ7xAH
YOW+kxzJX8HppZOWwgFlTm/EUDrzxd3D8pSD5hIxY7pcZhS6nJYCy8ATDfFk
bbdsqhG4krzIOFOsnhC/BekQEUd42ZVmahoWqVR8QTVG7FBuwicLVj0TD4AU
FUEbUvuWInTTme5Hbd1xQP3Kbo8UZQrmwFaPpg56zENu1dueKI9j5wcSsuFU
e+54OYogpZoHkl3OTSvL4bGsz/Tv+h1xgVlSPeB07HVZR5TWuuB8mXI8RtOW
Dh5FBLLAJ7s7yk87GIztTWp/yFid0VLEEBkRq93E+b+dBjPTU8NCaZptLyKe
K6DWD5faZpTKqe02zDz4MQLvorewhto4eZCPXfCsOQejVrpWIiqW1nsysI3U
BnuZt24/IEN1j3ZiBzPpBUFm4QmFevu/jLIKh+5cf3/kalAixKAq0ltCg7aI
heaVAVQuVJB5+8F5zg+0pWd6YPFTJAPxaokEEQZXTBUaySuBIpH//9NQqr6w
RVh/RShrkdumMX3XqHRyTwtnpfp531PdgTNItHR00yaIz3CJlRE78TxlqeZ+
hQ0TDxEW4rUGMNou5a8RyCYlgUjR1HXOAEfI6coo0lVw2hYkeXcAf4DH1/Dd
g10hm9nfHa7hW0ushbVrWY3weGS98/5/FrQVGvjjUGbDDFvKDjtwNpeHjXmp
bVnqd8GsmJnh+7ojYRJpdHNTl8A+O5TFBJtbWD6ITQeYtUmdFdMU9pM02Fy8
bTGSFT5xiHauheZFhjEnNSH2LXdA1YpJWSNZFnJ1Glil1wNCXXjaHBQpmF2z
3cZ5DhZi9EanSyFeZp9R9pA5fnQA86u3wAiMNlD09OYZUAAYJGtkOsn9aBhJ
+0c/9P/yUIJxFKYlJZaQfxmVtJPHOmIiHwQK+rj39CAtwMU7vmC9K2qodYht
hwF69vZGSqYu1RGKzrL646WVoQjbMIpnMv8V5tZ56AP22nQXF5HldWDOIlSP
pwGaYGEIhiB2HgCW5KKxqUsR32J/Rry8jfD92sGSW0MCah7gMJBC5EfwneWe
ddkcwu6fNm3wULI1FNNtAp6aLN5+ADjAqFOyqBc8BK0YmY8dfZR3Aof8g+BJ
7KwY2AGFIKPz6jvZ9pkVt68L8Hzwytx4o0/DM+rfUhbLYrN063v4ajW9jobM
t3SgX0mOXcAdkUvcoklWkhYExcUi7N4CnfrKd6VriuG9GFYXN6JvhnDAOClO
A3LVcGPvRSy1VR2DzQxMyLiBa9MFvcRQV1RQn5tpyER3vPDnw911Mxdcvh64
rl0F87TONUzbvQkSnodOs1194NEFGRtNMh5KGDHgClcvYGQ9CiqznzJqYoVW
s2GGdD3dGsBbR1Bt5gBgjha5EXIELGNmtZANf1uCMOJyaOHyIj19DOF3KhZc
Pg6xvUanj8FQS7LowaEtp3oDuESN2Knx9KRuG4V1ibo0IcD7g6M5oFv3knXU
lzVIZ9mtq78srh5S6o4dLdqpAviRMsd1tj95G1mlsUtgm/mDoYRmH6Dvb1oI
cIxfZaW1rvkSwD+8H6/J+0zLJID83Mqev0oAuIngVguTkeUz11wXBLhEsbx3
nwLwtun4XGZScgwAUTfRzzkuXurbMf6jI3S5Wca+DQ4VPP2mHAenBCfYDmWp
9IkDeinKH/XwBl1A+xV0zEMgf8L8sMwQ13dfyF0PAwk7gljhcYdHpPu+Zg+9
3zIop12iqHOm9xgFuNpWsxJKkxa6QigXaZcgQZemnHboUESQN08nh3zguLAk
UFT/ojcVgOwQ9u37c9VHZzGn30cw4rtPBepplRURmkZPwkdxJkVAdIAJpXU0
z9DC7UbRFTQg5kNV6JAcELWtLRx4SSV5gVhcCn87+WOYLyREv6FPH3LC0NZR
U0uGd9/5HcVzUrIjhpLzhTt2YG5tmOUrtq2siEehubWiSW1ApKGsZWXDpwAr
/EeyDmRd8o2obOB6coY8ywPBiXPUikUWwyaAQOEvgtYuFnqRtp0wIgt/0o6e
QlH56i2bBT5wJaCIeTCGb6M+3K5set4kmaJjrmSWTuDeSz3/rbpm3uGGEda3
oXtWs0BnQE2D3mi1vZcNaG8Nh0ZFhgmvjEeOkOfUZsskGbbZrn50zC29i8vO
YQwmp1aJlakxUFqXeHZ8qhsdlkQuhOH/Mk+KrEVQY3wh0+gQJokU+mKIuGUC
f92G4m0vKIYc9OOGDb1lt6MShzFsYdrtdnK7qj7VekAmLP0DGyJiw/U5Gybh
GVBXACnZeIv7tLcDYAHbSPssELasyLvkY7lRZjZe22fLJXxJ38fcESmyTa1z
ik4dMlhI2PWmp7qYGcYr3D64GxCR1/YflhKEAWqO9QpsGAn4AN7kkDGPYm1p
ijnm93bRq1omfsnw/ZMl9fT6pB8YNsc4IYUxekmI1AsGQRtg+VpwAijJvZz8
BBoCF7iqqUmfbRFWQJ7yCNk1r+Ccj+pToE913GaKK5l8t3VUZoyR3AMJ0q7X
lyt1XSiCAKD/9Xp++HYSf9d5XwuKrKIUiIr0M86EfwLuhCu4SILeqmJT798+
6BBXKwoD4NZuRJk67Nr4z9VeAhSsj0VHpTrrshUL107r8Deanq2mayQ7MVoS
vBBqF9YcJL6TWxfOrrgLQwN8MDWSH+DAO/j81J1ywxkGkh/JUTPoOcpRDaoC
npWT06s+/tR3MTegtEIy89NzZOxJ4YZ5NNw5TElAOr2p9lLysbip0SQeLxlV
qUh9dBLYK1jODEl5Bb9gQfOCMeMUcCGcoHJMED1VcQWHCfVDG4MyaYGzg5bj
e6wQdsEnX3VocUpoLLvuipITYSHuVh7OvTuDWIQ11BKVkLIaPBYcrLptcy2I
NzXMMSKDbHoOTq4FnsDSi6dH6Z5DKZj6B+FrocIsMu6NPRdyaatdGNe+iCuU
JTCAZyCa1YK6crdEckR9ao2UWus9UM3V2JWAq+nPOTxFkeW+9iL0o0V54PUR
PncH9ejg7dIc2ytz0vVkvHeKdpdXmcUSnLM1+fvEWEAno+DmPPreUVm0GbiP
bn08tTuzgYVR5Y+Fbue/0LhfNXCAXbm7oKPSN5EaKX5FEdb/xqDBrSuM5aWS
MM/gq+1Hsuz9xZPqQ7p4Fia4VLQ7MKqT+Md25iBtOs61eF6gkN0s+lN7wPAB
qAQ3aGYINyKcP7tg//Or7cYlEz4MBqME7TFLamaFDW0sfZt+GngwL1ZDkLDb
WcMep8CuXVsCdbPqO1zEMiEntPFpCMq7n2Oh0tV5EfhBrLUs1nWt3ZmZAouW
zh8hbkB5U7MUD0rq1SQzGXMgN1p5vEbNcy0HquTC5LaHmm8s3nyCsIZYDy+h
qbnyAKPNjavTtYQCNAt4ID/HSkP3hug/wo9me89oeMIKqq3/h3+gqQ5eHVsA
gar5oEpuFJ183b2+WWEse0JL4V7iyPLVJw2lQht9RdILV8qaPmvNKFUPrsMV
/kf8MxIufCaVwy7i9Gy9la/5TOSV4KX/zJI8J5oDF6O9GVXQ3G2mIj9p5KQz
y8tOSxNhH5HSjjoYV0mmdanZoxO44ju/DamBYnVw4KXgjH3bNPpo+SYZggQP
tCN+DnzlO0Dt0lBU/ESxmSFDHIRC5wlQd2rnTx6ao9QDH3YurMSgR96v6zqx
pUT379A/0LmxdV8gk7c8PImwyt9R/F/2mN2EDIp8UrQf9CYNJtnU22Hn8g2e
l+lF68A7SnGrB7rKqjTc0AlY0do+UHvdo/sk5v3xZbOBR/WDn1NyIddCiiTQ
Q+aVfQ2fcMqo+yh95N5pHnMHl9xKLChLk1Ya7uyM97IaoIbkX/8ymEp3GQ0d
u6DlLBjgpt5X97IQOkodzX+WPql9FscYxnnmWL2ws07MkHVnmR6Q01ldYOlb
gtKkPUwNmzIUbZ1AUy4JOudzVatySAsi1r2/OKvybn7xDWMVjvNUoCmULbjF
xAhO6GAm+vsM4BNYKbEy9Tpzq8AAubFILnX4WXRijXBnnx3yWMFRevuHAY77
7VOQ6UmCjFJyJtodJG5LjETMFuSF2POXuMSVAIMB3LJpbWqHfQwHeYWXehQn
fBmX52PP+K9VPIrv+Ctf/lhNUvBYtZVV7zx9x2TJhEZ6YEQH873Y91Vl0HJp
8aVIuymHCJPcMr97Dqb9vQgE8muvQVMKwyDWJe9ZQvbzy2z8zK/tUcFUgktp
LAUZfvBGSm5ah8f3V8dE1UaGytb0LE2tcIYCfj2I134MMPjxP/+PUPRFvquv
MtTnsh7qApNbeMrGq0E90mopguoplRXbnSagrqvEaEdUKF0cSO2ri+GRx8Dg
J6FD9ZL6W7vu26AA4QmVxYdw4LxsbijygXcYLjBHo3gsnP6J13NT895cfHIh
Iav8+77gcbqiYZ1eted1Sx7EYhz6/ONSIARIx212IQgqUKy9+nOzdXFHsl0D
pCX5ObwCddJ1+LXcRlODEjgxhkakMT7IK0NyIFXARuuel+PJd+5JbQESTA2/
I5ppU0RdIyzhRq3/qEZZ0EL1RI7Qd9uAeCq2vGs+FLrW9dg0JaIhDNtAfscF
prk3k7QwFeKeya4+VcpzfFiX0DKY10mlNXpX5fDAn+UGrddqIuFopTEpHl3C
Y7R740aA7gyz6qj1vxtKnCd1LF5njRobLPmHfOF0COsm9Sd7vFM+nFWF8yHR
QnSufb8mvyhAamAzcLg4o+a1BgF2ea83XnT2Iie0basgOFtlvGm55xZ5My7g
s4UDfLrwMJ70As2p/wNuNtUQRvNrfkcFRCMsHMeSHmN80E46wCJswcxEYRta
cMS51a1yehRIVJnjhhv6ox3fOMyzZoVI16WTzPKsDjL8EoSoD3q98ZwVRZO4
BhxYe+ChPeqJ0HJEJf5nWyP5ozvAnKO0TOAYKgu2CqPOxn7WdieZq0krSa/E
oqd/nIE+oPqnoegO4CX0xLLS73uoMj5+1fqMhoHe4lzZn/dZJFP/yV1zfXJb
fbNcO3nODfksgNzlqf83uIvyC0JaESvO86mE5E8F4ufJM4wSwoBW9fX0xzTN
zVGeChD+lfzdmiGX6kk3WWLG57+dMnpv6HzJZF012lC1qOfcozMDF0oV5pnA
0BvIlulMim1GHZVkHoOVjRZv7UXYdwYMrrwFKvYalE/YEmiBINozQFLdElj0
6VfVz7edIj6xTPxRWwirZ6jo+hxnRuDdipUmsA3umqXjNcZhc8ohE017PsKa
3WQaZnlBJfGa0OylYkLb2SM2bAjEryVZsq3qx+2U/pPQoZLfZn8Ms9qiioeG
jvmkiRdDtF8tiot9gHzcx2CdGSWuw8tKxpI6Kt3P7RfQKj62cEl6NWj25jcp
Nq11hEgCnJfkKeTkhocQIyHMBDicUiBQcXRa3eVwbd75sypY6zSeZwpair6v
PUfp3Xxh2JQzXuGQgdksC5zmlmvg07ufDpehcoRy9Rb3xxi5iMZN1UQQJynI
KdWxyQ5D6G09HM/9PYpNiVP5g+hPJV3QJN1PsF8Ci3B3TCAnYQCsRbRvhoAJ
ThTNyV5L34gxI+nVHpBFUms0JPbiyaG30hFHnCZ/GtJzZ9zeC6j0JAiCHpNm
lIIGQ3UwoE90e6RtINMol4hmBOvX/TnA5eTdgBMiGPrnLGp1J+q4xBallvTd
a3wm8OAqdeuq/8scAhE9Xn2E/wJYXBtriqVg2bnTmbdOGtZ/PcX/q2CGjWdG
ucJxpC0iFjuNnpQMdSO5raFCol6WKi6M6XnDjPeRUY0If+ot05xzQ8gCLGgQ
9lyM7BkepOu34lPU8j6ieqFQB6YAezovhpduL4rQ7P3dAJUXwHSUknEwfmW2
b1Qs7SGYlusAhkrBHtWQ4HrHZ4sZTbO0gbsvnuLqwMTSqMr0JvB9e6b9mUSq
dChi5Fw4nQTuWA7cFj7PlUPLamZxlt5EYT5Cw2nUwf9uTneoiwajkoG2vZJz
4xqnCJdPX2avON4x4ob9k4cJqCtqK7ALZ11lenzhsLa+F7/CR0TsKPOHfGxe
MmmaRMHuBaqIFUUQGfWSe4XNBrmt0Q/5zAcwTvj5Wl8qsMzDZ+C0sgwVbjC6
0YyJuKFCODgUSKDpf32SwbrGu8CZT4qCY6YLuXA8NpH0hAlI0wMbMW3fMmB7
SEQKQFGF6RNBQtFE57Oo7fX9mzXIX+kyrSBwaZzo7Awowp2IpH3rXiWlqOV3
TtUEOSGEhbLTPXN7MQHl2/ml8tWxgN27OLxqdfTpo7anMVpHH8aOteRdlhoQ
lfcaIUKV1hSaR3ti7obV4vIum3v0JCI9PgIW+itLMHKYoJ5jWXFigAHKPM50
Rq/PTYyqpqwlfMpS7U4I41mjkw2MrvtMJ9aXtAtKHzIZG570/8Z/Tn6BUymz
5/zy7gpTy2XeKDa9unci20SK6/3p2QMyH98mFHejb3rvNls/qO7hGMBXg/gZ
NFwU4kzFPl65sdsDfgUMBkM3S8Wmqqilb0u+VLQ5qbosDxK+1wSi40s8K2+N
kG4Rm+srT3zYo2UQy++Bxhe/o4F60Nwg63EhSDz6NCh2Kf5kikvOBUP7nvak
XYUOowhF3ES/531HFWmLyec4/F1l4OuDEX4sWnIB85Duf/t5CD9ViTDgrdBV
zPKkaCGngOvvQ+s2JHCPyAMKluufy5cFCidx68vxC8frddzzw9tEoMfndS7X
PyPsSejuieawZ3lal2+w13sv0r7uhFXXDYeuXgKVDGN1A4nPNRPRcgBw7fzw
bMdQ46BlrQ8CnIyRno8YMngV/oMl8Vr5L17ckBUApeAh6uNlwWeCnIhRNm2e
2OlO6IrT6xLSpPRoczwB4mjIP2Mt2TgfKJfP2HV5Ob69Qiw/M0iziNttzGdu
9fZ3fn0R5CUuqyokp9jDnTnvZRdDmiOPvRmVjbq1dP4p/v5BvQZaLZIZXesm
gocQhlMitPY+mVeUQ7IUqBmwYqGf8COtPl9dOgjTliQwyibLJfg8FPU6d0Sv
USQI9qGWL+2aF+LsoNqNRNlHlOL+G8NaWOetWjt9F9I5o7TrvdhyA/jwg6hf
qtRRXrBivDLPcOXg3stDAp8Hy6ZtfkzPT3fKy5SDH7zZJaSfDdhli2qqlkZt
5Z/d2to1sEH7SDybteVZrC1qDsY1MnBx3dB9JVSttbqIOl6N1PxX8LNoO5m4
Lx1iQS1D5AKacD00INcX0OR2Qd5NHWMyYWvM8YCSrppUKvmiQCJrajRjNLzn
mQeySGQodKHjrjzGSn/Nry1v9gdndWN7Btdc0Vc9vH8u5fStPKUjnOWBJw7H
qw5kWzse+skdDMxhovI3oYYjun/DG49HpZXEaTqT6yOTAd7RQnhGd/z9/3iI
xsb2C8tawaqD2pZOuOJ3ZMWfRQmy1eNty4Ob58lOeEivYx2iPaDYMNHJh7yp
Dlvb3dHnGvaGEIHjtvL7HBdG7Vpn30ZTAkmOqJUMylNdCGntDkpSmu6iy7j8
IXEDJxT/YOj8TxU76DHFMAaDW3yS0ck15sZfEYIgGexGQT+C7a7t8zEZgnCA
wHNbA8YgymuwOaxbkT03Xa4i+2poN7AHTkEEpDorLBYE+TrGTlpbWWCSrd1s
pC3yBhgjGCzIzKQWe13rjetgqnprYfad5DeiKWEyEBTQ40BM6eavFSH57/LZ
D27WCniRIU6h0sulkucZVTIjqdjxbo8NTOQxq97vi3XAArNwj+XHqbf0U6GK
l238BZzcWo/gT8kBUVko9SWMHH1TS6peauU98qBBkNQp+yb7obE7whmEVEly
w3BvSOTOjGHS5RDdbkTSPInZDiFS1nAYf5Tjw1k2gRb+xVfc5gTJllwTKTm0
ikL+nX896Nb9UyTmKRTl5As0Jn+j+Dv/Y/wRgw/vTGwZZ24Q1qK6VVlIESEj
8ekwUq41F9Z+1jcG16dtMIGzWm/NwX1OD5ctBzT2hGUpQoJgRNgQnI6lc8Fk
MR+6IrfkHX2Thynr8TCfvIlFEqTDwpLpEKXbf/Im2fir1fK0e8awJpPnjafp
8UWd1wnZZXFns+V18ww+FjmptjI5mLHHLhsTFtJZrrB3QKl1eI2QB1IKFfN4
eYbJb7mdI/+572hdO24HFTLCVwML5PNcOQMOTmQYNHko03RpN4wIv9v1s3Y4
A2r00zktW+76LEetO0VadiYXvhNES8M8scMOKRPxU/WKJrSE5e/hFzIkHfSP
JIdQoYToeg21fFxsF23vFjEtYeWAHEaLvHE3HaVtCk/207UDY9dzPgUz/ujd
nDUA2Ca/hgGlH3lYzYDWoXDVgE0EAENf7nEsHAXSiNjj4YafmlgcHjfq7uB0
pNDPa34GxLthpkViM4N2mHfAHF2z5Oxo+Luydkw+/sKhrJtWi6t7jM6nxat/
QUElyZYvPmuAgfF+ZunZ0cz4kl8x+doyXRDLumheSRRebp7RgrrOuANMQ6kP
v6THnkVOrBprcbip3Pz9Oaa0EnxPsaZW97Xl7JnQ8sskq4SLNTuQQMzeYNI3
gdhqjsjrT2lZshdgUsGVVGgILWxlYD3V5mSf+Y9v9qzmn+O03G6ze+PaM4Ow
kiNNO0X60B6LBNHm/BBJTX6rH2FY0eC9k7kyPahfXMaX8Cq0mYs8rX7YRwhL
Fcipf9f0WdwuhwzHkCws1En0PucK958YHHWIwcwxQwEGFSYxWI0j59zXcT3i
8kGTIhNDW4d/eqUx632wm1ad8OppN8VNzSRrXACZMaZbp6W/kK01GPcJPPEC
2NsWjg3IFfne4pPovILcN645r6VcNjmVKKXXkOgym7zafKP0hjKGMeSw5e8r
ELQu4BxSv0Rva/h/N8jJihgjQKq1DMOYwTV2Ban8tVJ3We0h5XryoSltSet7
6bgkbF81TN99xVDNnb0gYnBqKUCF5TPiamzmybnOMjL5px574Djh2qaHrDVb
JQ2fuVS0U1Wr5kZRYDZfQo4VNuxL7ljdCaU7wQYuRVpXOM4v0uOq3Kb632EU
NIytWNA3SAh280YnkZ8r1hQLb5tRbPCxtfobv1/SXBqYB1tD7CYo8EcjkpPa
J3n0AhUVv/up5M5HEyscFFFWn0IfJVtkDcZMGyKRycoL4+qD/DZyo3vWtItX
kzC3fppGUD2cOyR0b/VPBPDZPK+Iz56F9OvHcCfwiedu2rz44JOA1ymTHLNE
6gkZz2bwwDpOdqADxK1xVJ1W8v20Dy/o4/lYKVM98CfZB6kAiDarVBfUYj7Z
EHOhB9tgqvdoe1/tqoAtnChs6gUi1nS/jV/13OxBZ8dATGQMb13xEjOFwg2M
6QZtyX2TNbPKHfgd1w0TTbCgheVjbZ5WIBIC+VaP6Zxg48OcsBUr6eKDgt03
oES8ULBMMw/BJV/919oUcUgPios1pyXFcgRKttfA6Ukwzq8SF21pU/rUCCul
nwv31YCrKa6r92z5DPUL5QbPOJWoFJSwxVhhxJNIMSYN+SW27pVs2q2wBMsR
oiDBwQ3Qaor/FCvS5ou3ne6U26ENF1hTWdGqWALI7yJLOqHdA70XWBiaZteB
SWQV9P2aXGhqqHFIPYzn2+Vqby8G0zkV+R7N2QctYzkhWqXoJSlhRaj7hvL0
IoeKpSTr/org+wD479lzVqnnfkWqJ1BvIs44MkCAw2f5fuTQ/pGGae2jmk3U
i902hME/TgHPSAgnmajbSXS7Bdy6oV3Dm0rCT6hfb13VfMWVQ3eoB901jNaT
5M7Kv2RAjNC85EY0tvnDjVZgSqqvGgIzovytU+EcsCv614fD4jcnXC2Hz7Br
sUbgl9Oba5Dl8BOUzV9NK3o9/m7kgRTAeGUZOQFtlcjTRn34twu3dmRdYy/4
gpYiTnZNHo0pLWGUxVnifqDjPpqldfpb/LU3sn70Iq3R6bDFm8YsUCEpn1tb
l1NGM76u58/OQqzBrYxzXs4HepOPkJmL9Ixudt025KKltMkcY4w+dTTQpsSH
iUbwo9mZzCxddVUERBNkLAVxAnAUOjVVsdPn5vdbMxJjsBRk82pSicg9U19P
sbFP7IsGjlRJFdg8u2AMMZ+bx00U5wDQP9csnhl0n/VcwGl/WGL7Eir2ASQk
+z43VfF4Z16WlTzARzCjCLPpN1oJsFFz4mWbtJgrbqeXP3zcIXrNslsl1VLI
kYIWlv+Imwpd/3959X+QWqd/RhqDlpM+3BA0vovGxB2ukCktXyjtbbZzP1mc
hgEl3vXEoeBoRXMRYbD/bM8L0kKZZTRLZzg06sPP/Oma1fiTCwj/HqOAQQFB
C3WK2isbUrtyiPhnwN+9Anbf775OxQUpC92uI+dF9PezAbKQV1BJZNXO2pN7
BsryevpvqnxmDR0iXF6WM69gmc5ogZVlvH5+thedd52+iakiyd6iFEW0jxSo
vH8u9w42CINpU2UefQxuSNFA5gdRGoSuWP3jwz7VS9lo7hH4FJCPNnNruqWJ
hL1J/q0y003dNh31UnNe5+vAungt/Rbgq4ahuhpQzehMfECaLc5SGwc7Gyqs
NYDoUQ28zJ5Aj+AwuFAInwGM4jDpwDpJm4ztIOd9V7XPEP9nlyz+aKHUDLT3
zoHoTeHqWaj6BJi964QvzgBKgH3ojo0e9SIEjtafJ8CtcjoE24iUd61hltBH
bOfx8nfAqLsA4rFho31Y8KjZCIfyXumSFGa6KA208+X6vy84lNS2R3ez3y8u
p1+9gt6ONVVPwb1uqb2P6RZxLSkk1MLGNBSecMLNn6n96nFTkelOogxfgxqK
ODPmkiN/wx3a2jAUnlbmxPhEcmkYYp5dMITOB6gqEXQg672pd+Sjso122pvm
KcQDwKJZ2YuFTCsbpwd/HU9QON42T3CEumGYoSgkeT5iKvxCaUgrKg8gmdK2
kD5up5dyKNBZnbM5qY5SWkA6SsgOvFlK1WuZlHYKoPnObTKZIHX1Kf5paMGa
sPHY7w7iWBUJ6BkkogkRUttpt1JOAwf6dPVjASCnVNMw8Q6hG24mCTIalC8t
bX0X/6Dlx2WaLN1Ojw1mq48OGj16ez50lDExN3e3NMfUXOxLrqGA4a5NeoSd
eV8pK5ti/CesZYWK94Goj6EDBk84k2XYnRWDgPcNLRhbfy04FQ/zBxk4pv6Q
mY9Gvhd+sQOmW2/p5AhlCZMtJvzaoJb6RXtDKRtu0cvD7aotTFQxqyOi0RwE
bYFB9uwbGjIgOYUNW3+rkJolT4rIQYSuuP2Wq7Y7yE1+dBMw/pABds/2cXrH
WbOfzxc5w99QJcaYk08A4+VLFgYpaE7/N5r/9WetJojXWAsaU03O1Olh707u
ebNgBPTeaCrPLB4hUUGmAG9L/12L4Uoi//u1x9UNe+cr3leIh3OFy+2Rb0Ix
IyDex78P7zKHWKANdX/x++t3tMFQzocHFLbUDZv49aw5BZ2yk2jrufHfDkQ7
24xX83CE8FOzQIjXyePDtqqpQniVo4CR0ceGC86wuDzoWjer1WElj3/P1r6P
7fvn91SE0tja8LvpdiJC7dRMDdujN58rOSFxvZIouhaiuYfQeUCSr5LU1wZd
BrNUcxCjqInaFYfMvW7k/6SK4YvxDQ5GQ9CqY/0TLI5XmemFME7OaGHS49WW
7LQyYBbaHO3qFHNG/4C8uwIwK0lhU5COC20DsY3eW8OSTdWw6yGB2TH1Vddz
4dq4v0oZTymxtxtAbVV/wUrUxCfL4lX+oCYejAFvWiMyvqHQgJARcztTjRiq
OjhKg9/w0QrXqnX7FA4flpHO0y3XM391AJDkFFT6zc9O6elCBs5RkQb4byUY
UWuXgEpgBWhNgAFVyC2n1rZy8WQdZeV5iWKMkt+kcx9zd0I0oyOrhFfC4e//
Fu17PnWJBoLKe0NsPI7Nd7jrE0TD+7aPnK4h/weQamMxD0M8wpJ7XpoHft3u
Q4mhj4Q2O/3wXEHt6u/GlQmbB6sr65FUvro86dmX/XeNEba77J8FECLGcle4
ExI5uQH5A4PXDZNc9/HbdL52zFYpGbncBh1JhtbfaKuvw8kYoG6dVjJ3esD5
UEMyM+A6hpTwgYLgl878KyPwA5a4t+m5iQ/+gNAfb4+kdqXsoEYpCwXGm5UT
cU1oRz873cCpuUbg0xYzVjiSp8/H2Mg8n/M0w6VaclPIsTrXEsJjau+e4Wbt
NL6midG/ykTpCz9VGQ+/hsZMdjPfSx1WnMG7m2T53drRertZBGiGElXYIK6F
W6TBCU3Lu15i28xsLrqP9luL8ItSQMgnZCTTPhuWYHmn4KH/zzO/fmUuVQqr
3NdSMWZ2zx1Vl7pGUzUGSAiOtz1vK0m0y+P7ekGAQjHn+O1/8VCb/o+qbz+9
iub1codsqNteOuRw67fQ/5TjCL5LUwKsQ/C4SUP5snLrsRu0Fc/vmbgAT1FX
jybmyQs6jWFGnYALWjD4Dc2G6VxJ2BTGJ3yxxT9Uj2wfUUkWIUuTFfu6S669
O0A2jB7yW2O37hKNdecSLf2OrgHuuTdJ7Dx+IyNH2/uPiS7ay2JmzUcFvAaf
8BStOuUAPk7i6W2Yih/CH91tq4leG7szp1dyyFIlVLUDYCf+f9Ea4a4QEqR2
uizSe77weFPajDZhqy/BrMQxVYur8c9cVQOKjwwn+7zyr2hhDdljRCSM/N2f
zJIYdP4YYcbWqJfifz5nPshX4bD3/eU23nFq+vDizSoGq80JADhTAHcBRxbe
+pdvq7lEoWllZRZ9vuf/Eep7ZLTFRc7eiEMpOA27rxjAW1fSLCl1zrDrmQOl
05pF0T8KgxNkrUjZ0ZXBbXDd+KJZ2W3Tw0TAX4UkHCEhxmMP7Md0vQdZktQ1
8Epg/IaTzCVMJCwv0YCvx12Eou/K9txW/XFK8iJgAe+Ke02d4r6TzVVjGXOt
mxTduuq41gZ/EX/WGDKzR84ebE8GYxX3wHj3IgKlPsBdoQDz914PRA5mZlBm
Raoy/63Ubb9HKcJBYTUJxBA1PFDomcbMIPaf1XNuBH1JXtiKsc3kytYMgLVv
g0Z1X3SzFehRlbWZDKYI1hPnQ6Cs23T4JbY99Jtc/xaISvWTcMhF84ym0ZoP
HeTxkpSnKYIm5+abfKJ3wUkesEVqNRlpIkRzQUWCynf0ewbfW7UBSrffxD9o
m3jW/Gt3CUgnA868jbtcwBk2ut6jypN1czEViX/ZFrRCSN6+8Tau3OBn2KXU
SW+27+JTzbCtnxE0wE8OAYZf5mOXVzhwusrcfr/rImi5c4Yv96RMFHkj4z8k
ix29W01nx7vJRRFdUDCv00am6czg0mkxQ3TD24qt6ZEVLw25wTXk27tXYagu
ysygeRSOTnkKF+vhg/VthhvPYCG5rxOwvQYyqWfcHrcWVk6pEiVdWVDfPsof
UF9e9vD8589uCSKWDfpLvJIwSltmWPRhn4V4DtsAtA/yHtOMJCiQ0tEikUEg
hGaJQ14HKJ6ZMIO1+lVx38GYDcTHevXpOrk34NL+oScXdGn0lTNOpLZwG1kJ
6h9DgZKlgiYqNsHlM8PFNibHwZTMjg9l3e3kOLUAADg5UeSQusz4tuKlb28e
Ml4mUr1SlPQ8l0fDChhU34vqzOf46wI+9hDcaiB37U+1zYsv6GAIzY8yM+sN
Hton6HSXl3MI55sIGhErlnPCrliyj5/7BwOjiIj0R2bywv934n/aI8cFmUoT
/qU+5bswcrrSMJ9IQVViLHbgqAvdM+55SSZske3Bxix0ZCFjlnRAce5zvk6B
HCCUU7AnArxaLzPdJeZTIOuBcYuixIb1KZQzHEJJdemHREJ+ijr5W+aufwbT
LJFJat+lA92wfZ/emIwpFc831Re7Q12rllZ0Iua1DrkOQKwdke3115Q7Sd7V
xLPVJdwEoORdI9GYlvDFw+9CpyfXX07aM5nMZ71DerGR8oo3KMZX313uLPxO
vaR8UtTcB+24VeF7tJJJ0uMfR6xy0ja70sBOTyV0HCD9z1RT1VcUULi8flFT
tPRRCUoKVLNjfnpzhW73MsTM+Rx5acjg/heweYvXgi4YM3eNzVjJQPQ4+uHV
5VQ4LK7vKOGbwrDKLJOOOtiUjIqBeEVHkS8/XMpTXk16njPd1eoJKbZYp2kG
FbXs498swsRI64CWzMo5YmrHRuDq+26byeq0YgIAn0N0Uoc7hcHDXA2tQzfG
uIKI9mz8kOSw4QGtEFG2rKiFmWdbui3b2bnqm0rEutSfrJQOJ168C8XgBo5C
14fJ3yH2+1qO0pXOw8pMhIird6mHaUX+nuBXxe5mQYqErjwxzyejGy3GzF+6
PpnwCoV+fLaYwTGPsZgn9YyrrJqJmphiXtw+oUlItq086KAqfzhRge9fh9yT
/ZMVVJbP51EV9fYBT8IpY3nlARvdlX+V+EAZ4KCxP+tSTVAyuAIlz/JHfcra
ZeTgfPx0sz/Gap1/BanrwTkqFi8wecqnxWYrU+zFvmX4uFFXNh9FRBnIFD4a
WAfX3I6P845IQFgGp9Nhy0HXVY24YJGMGY0K1DY3FoS5gJ/Oxel/SHbSJnvX
U3ic0gD1itY8m1G4BG+F+7GXteaoMtczHiO+JdLk2Z+S/SbanNa83yYdVs22
rUyYm+dLTJbYFC6JruM1/MKA6kLkgkHxgxELNeHovqT35RZE4UNf87NnsCvM
jrNx8A6C3trICjcc4nOThHOL0+szfOrP0EAuTl+fPWEo9kEDY9B6SJJDZoYM
Ks0asS3oBHtDwh4XDb3IPkTBDXHAt2s5GECnFbSK+sEhOx9nju77upWI8FaP
8JSc4Rt4+5DwjY//sue5fxASFQQwKeAoQoo263/jU2PLJMaMdlV06UT4fNqT
a+6AjeayinRpSWcJWxhNv5PNEAFitrthBzSPwWDj+6kdbXu4nPIDbqqU3Kuj
MbQim4mt07p157ezmGuHEuMWeJ7wAAD2JG5iluOqEJ+feqdu4HOGPujpEXcI
5Si8KjSGVFXZlF+/058tuju3SGiEPfRTj7fywPm/anjV7oHlv0B1RNkIJVTO
S3XOUdtLV80Zlxxw2KDU9c9VXpCBbT5Tb235tBo7hYnVhUvmPWm2qpJzFFO1
V5VQq+R6CL0kq4uRlAp1JT7azczcUGqePHPRn8RKTh6AxxI1/clBO6HbL2gY
/eX/qRO0zEAwN7Jlw2hSH8wABmIakAFIoE3PBcou225z0s7s/joae9FYNIHC
mmm4cgahHsnyzHTPy15xPryez6XHIqOp6JMnCFltmd+dtG4CELf9i7KicD9d
k6rNnsv81+tMNj75R/242eM+cGVmIjD0gN8/L+Iocxlfw2XvIN0F2QnDMMjV
XDGGzKSJz70uyWZzu6O7q54EPer1OX5YdvwGQe1lMiwj+c52gLi5luy5zSGn
qI98hP8Mok3GFrvRgtApaYzLtxWSpDESC+HrEKrWz8OPUwBnqQ1sNo6g3Z7p
lgiK/1oFRn3SDrYer6rjbdpmq5ts6j0qM6iOdkrXY7GtT/VlhBXIOzYvslY4
CcstikRU7skm9y/sgjDBP85EQunFb50JlCTcvMKY3E1LWhUatjezgALALhW4
i+fmWKHHCIgJbNlADymFSTJNni73M+zyXOB1mIZCQRyUmpcgy9p7nmKVCvsh
M+Dd3X4rmQ50pesDTFaxQ58JGwd+5PDYvVQON06/EpAnKrKOf7CCgihCI6t6
3w2SvVcVmLjqWMigGi9g5a8/5uE2QGItOU2ZzZT2tM7k4IsB+b6JcXGBI3Iq
CutTGoEe7xgQoV05hbHvp3+0PIV1AcLCS+FSLfRGxwOp9IWvZPjcMQciIWch
6SPbxG1Mx7P7ac8PPuPp2R420OVU+ckvOyZTCN1Npf2lS+IeShIGX4i1Ki79
kVeXybU+fK+zhDuguFhL3HVMS31EPfd7v9b1XVuZ1+avuaRXNnHNttNaqzdR
sNFjwLnztKBuyXZdJayKa0lM5pAmiN7EWkPF8J5sG8/g0cfABFbLVN9UxPZ5
iziWHkMAKImwwuEajZNeu9SDBBM8WpaG/e8QtSn2KH8brtpNlhCPU0VYcf1z
vlFkZCnxlDR9BhfMTRBERDd97JWj0YnYPv0bLTu4V1Baz9DJRxtyN5SKy8bL
4TtdseWOeNDFPdZnpg/44OZSC+Jj8ugvDpsKiLSq7B8Q9PBc8OenMLFiTJmd
BHYLxhoD6SdTJcziobTUG0il9ex4iOsBv3OWSqYmAHVKQScN/Bxy7I7h/3A2
cC0AKqfEP7hFIn5X2RX/JKHiMNgXR0N6dZArQCGHZP3qpjaQ7SPeeNkbg2p7
UmcSYpSdUfmKArE7zknanoKl9MwnGs9M2cUHBw635Am9Rvf9eyWPCxEEaSLy
oBkaSJ20W3hHRdGJDhhE8PMDveAhhRcmhsV0PPqoCqTas5YHDT6tztvg6R5x
1W6Z0rbqy8oqEDmLWBciDvPI8JoTNMlEtCwdiMlbM43IXsUugX5djjZBUddK
MRBfVUCkcTVAH8IiQgs6T5iiuxG+rzNDwfNAi9OcZsFmbM/XblifIUOrj3cw
XYj7AykkyfYMQRxPjZ5PBSMb/86XutkfhSTJRGeFpzErP5ZX1tPSAWHCPsfK
Xn7L/clAKbz3MzvIJa05ZPUDsNeA5B6r//SZmD30xF3bxAl6TZ5pNuoj/WiK
rgUCG4Nfqc0ar8m4mlmmBaBeERHxmj9Ru6jCpYODss8DCDFewBbPx8Bc16OU
KDoOjNNPgQt/yH5nbmBUDwNOAa/FbrWL48Yh+wA8Tw5hfhL6WT342GPQrCjU
mBPAog/uKP4aMjdd9acq+J4gjSTZyIVLqYYS+Ps9nacMKTV9T8eNBqBRF41/
hASthRMwf6WYNxkJqcSIJKPnwxpE2dk227ySGQF9JYAcx2ehrIN6HthGpeW9
fRqNNMeW9QXmrUTJnS+rYQZDowDNisuN4vgzWcU4a0v8yktPpNZolI9eHANf
8Jql1DnALBnPPGHCEk6AP7xbkpXAvgjQnuFufYvJUI7RJ5V4viq/Pz1mv+W8
eZ+S3WAkvCy18hoGPkR4TBFAUedQgY8oyq6ArcANuRHmDEy+3l86Bm3wfvN2
l88VLYdwi8L0AVEU9Y0P+pE+Jjx+I8yv7EkDlRuxdeYD7t7Bs+6SD39KsR0s
yp9qHum+vgYLLLWb5esx03mRMbZLUrFuW6WK8yeGe/2eTQZMIiocjvGYM6H0
65PKFj/wmMggtftCe6BbLd/TrWO58/5oh7aBpfdXt6VX2pGj3stOFf5pjKny
mUGdH5zqqGdATx5ycVG76PX2g88jJR2sIsNwbtkXg48A/XAg4/h1WspMJmHI
bQjAoBWmAqyPxNL6Sf0QtQm7i30mkBvXRTg5cKrgfmCZg++lBikjsH6ZDnEd
YxXwA8k17wEDm+TCBs7AbdiInZYkmllx6876OgLw3k5rHI4kseohrvxArdh8
IaSIQNBjhANGbuMLTRoqup3YZFuBv1utkn6Md64v5RLJQ9ea4iJ0afppztSZ
ymeVBF4NQacdXK5fy2W0pfkdCFoA5PE52uvoEwXBWCL4N3jZd8PczpPDncj3
Hjc72Yrn+y4VukSkiKVkoo5p73w3lEJv3af3KPeq4oq0m/exiJwT31XXqFI3
m6r4pw32OKx9EetQwTQuYYCNu6CBTwsvJ9K/ZpsDlqDgNYKqOARIXRaeiJ9A
L/ttXOqkeavZGQr3BeiqczxIOitgh/sJdbbyOcCdbxYS9VEwbokpSePmN4/a
A3kAX1gAQjKPoUd2vWbvSBBhFthf5UUdgcQ9UlLEN3SDfZHPHdowXkY62DWg
FhQXFvg/02v9DVLUFgbG+E13DnBbOodOkzTsicSyz/vDInzF1cXeoqltw8rq
112mJTu222ug12yVV7g8rfRVsC36SeFqL+RIMb0CIxJdg5/xCYEd55OMn10E
+CbOyUBzinAVOgOrGmuA3GhmVPAjxL6XurWU4MguWZNyquqe96lzgjNf2FN+
GIdv37uANXsloLrYk28dGDvDCNlqXCtRzEmfDqDIopX8VfZFn92FH0+Sfdmp
Fouo7MwUT/1NH9FuqZSm5wy/U4RDeskdS0BaXxX6wPNPfopmyaKOL6MHG/HP
Sxt6CUDLCX2TiVQQzvU/PzcDDOezE+m6buzychb6KWJLqpV6ypFlTUaJ9bGo
fY7BPCNPvWRSGPnXY8yToip88LycINtz2XsVecUhpQSm6HjbCtE6Gq/ndhZF
s2Iy7qjIPlNKPaF8S1Rzb36qkePKiMW8DitZdunVccVME3FNnVB71QypAnBy
xZMdI6ISjzBbV/pOtoOzgOZC3qRGXTtYqI/v+q+CFzLJTgqTV2L+sJ1ZVHkw
yA2tDoEtpToBYKwyp92732pO2ClnYZ3yuanySS7DMKIpqhnWGMmRhXXnY8SG
OfUvFfDe1pxZj2t4hP3DXqUz0N9Lfiw2WLfL4aSbLvgX27tJrZ9F23skuTRk
qkiBdF87ILXe+TaAv2FKDcuIjmcQe1TB3iJW+XOeeE0pPbDGH+tODQdl26+M
pJSBAC5dyaZSvd0rJNyCKHBwnpVFWelQXDCnZurTc09L5WlOBJw4E+36PZiL
oqzY2M3MQkcXGcrZxu2RI66iyONJAae8uCvjnRywPfmAC4JziQj/FPSVL5c2
3GitQfa/JiZ4a+lzQcZ/9QUMZQFVQEQEZbCsuvyO5y7hG5rU3Bvd+rQNDWux
tB4nwCaigx/VSwXRNlUEJxJ/A7kaVmJf6qahd3B3dGCO7MqiSLMagVHUM/4M
Gb9i0Iq6bqqGYCsHXrGwhoOY5R66N+Vmv9MPUQE+X8rxGkAfm6ZOrv9F5kkf
9CcFtkrfMBxjgI2S1c7vJTVhLrF+5OLd9DBaTIu5fSVo/5PWrrA/UTGhPkhq
ceSCDOYNaYaF2XIH2bN8amPfcto7gnInO7auJO7Bk6gK40D+nTmBNy44GfVb
59intFs0NZqbzQxZUp4sTYGXYVvA7yLA5f49HkndYhiXk9O144a1u/pkzieP
+RBnmniP9SHWdjFFDtRard2uMa3NRY8w2FUzq0P7mWZooGpilv2iK2ZyIDzj
y75nd7y2/mYq1b2GFgAieEyyB7wD5HHuw1qanqNIYEdtsU2prdw7c01ZgENc
nYeNkyvSI9SwXC75Dq97Y1S8qBjtzzcm7g1NSyJitzeZKR1GVCvD79BF+Ekl
60pYaF5+lvn62ZNJP3qiStTmq5kGFD5/TmcMX/RLfZT/nut7xvUhd3w8/LdE
oEycO7b23JaVbcL5TbUFeuD0gg/A0eL/ZW26HMxmAf35YE48NOQR3qqDsjFL
LpmWJ9rR1gdJvXmgT4TlBwJNM80dJKk/FMbMvd+MqDHbTDWirmy3hY9m/9II
Ne8fkE5n6pXpF3qp/9aGFkQVy+A9D3K7iLDpUl+Jla0XTx9ZM4xI+ORRjEae
QCA0RSxNf7C7poZkKYc1ejrBphT9AJLqpGL6mKq3NxAApuBlAR2mNynadRqJ
v2a2734YrtghdTBNZ8SKoJMshX15tGQaTbQG7rt4OQAKR3wg38xQzzOZcXDa
TtlUjRCZfuC/LtRbEEePtUSP1RJOwo/xFbA1tXOM+WDFkgU7UYZ88z0K2F7T
1i6FFIOKAgVAJAckF62VV2bRkDZ+l0+mt3R8c2gFopcTAsG/11YQ4d87lj7a
uaSW1RbfwXuOHGlB3XX8ngBR3X7+etkmKP1lFEpJnahCCuDpta9YaqIdE+a8
/uOdlvyPPQmGD5Nc9841FIER3WTFmehdXGQ0eXypStb/+D6Dso93PHv9svvu
Lag7qpHRDI3yTzEtViTdTummIYwtNQmnwTvGpsFR+/aTUPDzDuS5WuWtb2fB
iDvlNK8z/+l8jHC4NwPJUd9F8Y3ljllaa9Cqc/GcYwz7WeONNgRzGfeVAyc+
Wr+PCVp62Ioai/31jPFkX1gcgmxfT3aqKX8n08f2k02JseqCz6JNFXnNnKP9
Se13VkHHDWs4BqEKfB5tfEUB0GZGGIOMdcMDcs/oR0bRIJ0Df/v0rh+G+aUq
8HVkehHz20CSB5LC2w5+MfUVl0FMu5l1tCd/Josl/yCXPR6rtHVVRO5ADO6q
rj9HFnPTLCFH3vW2m9Fl6h5OE5+w5hsOGswzvT7o4bztZKbhjP4w/kWtKR0M
BOvO01ofX4hsuOFXNl2uszDmgRjVjmU1l71mKGbSJw20N8f29z5gGSf7tIrs
3LT75/chS0S0ipMGDNO1Q2yhPFpFX1tXzfXPxNx3/WOlphS1iQQEVGv1ILzb
gQkWF7/THVDsD5PCHkEPWARM3S638QKviuN7L+5PsiaernP3FrvZopFC2axC
KNEJ2J3xHL8P5wcgJimhOWvvxYsFKu8Sq8gCymJM5VVlO1rIPAShz5jVgIT4
Pxw9BzfGblletgiNxLAcustSwgUtSYecgQXpqtVbrqgEVdPhgblo0UsygDtS
IK5ISeEZD9R1hpahQm15YODq+o8PYWV+9aUhyJXZsLOWcL5vlQo9OI2bcLoR
Ov7vJtkeLJvB+Qc5s8cqAPnC+zis0qZTFQiUKkXHgv0nxLbTNTdVfCtxnnos
MQQGQ6piST0R39z6Ut8Q5otoTPmt/RTgg8ofmF34BpNB+faJjt1ysbU74N7/
xAmShNxO3740sAgNyj2Ofv2K0Vy/fiy59bG+I9dCuF7EFFR2g9gEue0HYy7b
EWvdafhkPYcX5ooqCZGYNDKt2wAs1cLYQdVptWO/ax5iKzWJD7iBx8nuqycC
ehCj+mUz+no7iLM62t32/KrWr6236uh47pOdWKN4KKh/49/c1GfLPU0YgqSI
AmbPa0Op0bUTOryuo/QvIe6EmMScE2zykcJqPYDpGltvYVApjjSig4mS/Q0P
LOfYbjVRxoE8lzDKVHUzV3LqraUL+HszQtMazr7dltY2AwvsHAK0eQUNg5jL
EPztChrWjUbHxX95wzQHHMcHGnwv0YEXKJ7bhM2qDTFIhgrC+XF4zJpLVHS7
qGNuB6lK3QRRvn5yGSrBy9dcer4FMsUDkgwC0nHNGgbvXVIE9tSNjZpYPEJH
4RG3aL3e7bkEW69DfZXmkA641qD11hbB+Z/NaiqtpBRQGBe/QA1Ygdi8u1ip
jIGVbvdpGXddaK8WH1bTnaHHxYt4su8m093M5VBUfqY5HN1AD6uwKu0GZwBL
I1I2jP/Vw4Tt2BSEELHnFDi8B9JKHRQZYImbujo1R8c7r7qcaenZAYpM0g+s
jVUb42AsVZzshBlzZ7BEB0qd6BF57s/eVfQLM9/IKadjI9EUJJYixL3vBwkS
1+YnT7qOc06V9zcnSb31OMh1q9DbpYviN56NQq795zLIiNptYdG7NtsHgl+S
61xfwei8o54egbeg7xmEIz4M9yJy+yT+tSt3E8xnf16crvsqkIxhwC7fkQ0Y
bfqHo58QGdu0EgNn9oB2KGsNarj7hVGW5YfLXIek74yW43DSpLDjZZ58J3cz
2qwTPVDWXV98g0mPE0U7j2jJalwvxbKok5DJzjNZv5oTZat7elOrNUrqmJFX
AHuLNpp1YTEAa4QhA4Rbv4Fsjgvep7GJxp8LfufPMx07WeJQ9Ho/ya7hexVZ
LXr05MG2OmvDmQA07SkXwXp3rasMCVzQGFOUVY9m6GV8+7g7050guLFgXJ/7
ts/Qz7rc5Ha1pCtI4Ynoxp9Eiq3RU12jC358Kki53hV7/D4fzvAw8f68zGX4
Ni6rTLAKLvQds6U5pUIivTsK7KqqGnDMYFicEnFNERPcvfofq3p0NwEl0+9u
w3LPPF0VaVbI+cJhR7saVF1LnN0bJg9OV1r2P9TZAchXjEFyhrUvdCGvzE9P
sTC14pvEiMUv8HksYxC7BXOkNr7wE56wbgoWw5bPnFtq1pd/RU9GwJKxVDrI
U3qt6ogvZOWpzWy1BIR1yteQE3vAwwjwDutSNTyOqG9c+hNCso/ilSlMRzKX
0yhzspkPNrgQwwxGgKMSr7inB7P0W66mEpTGKL/XPO81AbHJlP2jFQy3TN5B
7U9tvKbnlC67i8abL6+4ElcaWP3Yz61iWZc9WxDCo5PNaxqu3zn99MeJQlyJ
2AxUINvinC7wGgx7TwKDxWH1MQ+ZeFNcG8Q7HGg8YycyPdPC7QIERhvimUAt
WnJF6CR+RWPatYtt+qFJVRWm5aAvK2TnZH7Y9gbV5s44HtYcoUesmdOA0ekP
+nmfPUWQDaXWjMGX0q0963Gdi1JalYmjjXiF9JVNoQlrolYM7PrdhQ3cvoHf
kWa6ULUXhXc1ILsfj5ZCUQ8aJRpFDSIPTzbp7psIeoJbcG/982TbyX373C5L
Cuen9hGQU6GBNXh0RF/raZXSFbSZMNBTxNMa3n7t3uEEbAeqVfYGafzFactv
9Gl8KgpfBw52wvN9yNARltzaCVQ/ffsOgdEFL9mU9VzNTuMUxky679xJ6VTI
c9svm2VRXlNwrJfkVHBt8JnY5lq1pkvvOoFmBktgAfHO4cQbnkMAEe0LZbZS
KK/5YJa2B/SteYzDwP+KPKzRh/Nf099XbcXpDCzm15b1KzccVyWsQyFZm/m/
g9o9EbXsH0okOIBmbnzVV8d3JJu1DlRhSeKQNV6VABPp/JRHrB4yhLSTlhu/
M+DS51z9yCDWZfdiPhIRzvp8IWW65WyNMWCRrNrOXd97L4XpilgzCPhEv819
en+HCznmXBS+ULI92D1H4gG2wMIfqgWCBP802EpeUBulUZLeS20BT2l7FkTU
Wg+ei06rho7yTT+qLSme1vj63t7JR7MSAV1MIRJ+bH9QBES7yLgwTpt0txrP
FYFiZFPzdNXh7GqwgqeJF6750pK2fm1afqq6c/heSs9hIl9GzqX61qnqdzVd
0Ol4M9LLMg8PG9jN57PEibRouM/i7eMaXdPxZkkeAs5nw747ID8YBXo3+9sI
TiQdcm59JLbPaVM3LE7rU2F8RlelvUj0Ly+KAOYnRItbwSRSp6ZpF+Gd7HZx
HdFsyHMwYx93daVm66XJTc7I+uI/TTmV2ZR8GPthhbXQOpjDOD/ai3J5NX5r
p3bY0o9dF1pThgnLBCUH/JPcfNBh90Nc4cCu7zsIXcEqkJd9bTKIfuq6G5wn
6nwAcdZziPzkFjBuuYsigZPENlth0zOgiKXzNIz7lJjv7lZcuNXpu2pMklOS
Bkbm8ywCTtjrIgHSCIMsuv+fIBEILV8WeSk0sdklX/MdlM9zQSzOl4ER+6Zm
Y5Mk9cswCN+oFlgGEYt0nEt5rbeXmQZvXkS+flgXKEO+AoPVWn37rBktpCSu
OOSFDCeX4O+aD5AQnvkuXphLvjCJMX6LCUULv1RwjBz0gRZiFKfwb2m/mjdc
AeFfZlUT3dhgciX2vUMQeeA8Dw5DmD73bMCA0Va1Xu1iM9a14hxwC57zth4g
ocwfZzKghpIhYzVnHk4FYTg4XI8qN0fFjVhOaD8EPDi2ixr6cc9juXTc9Bo7
LMD1ianQbmNfEX31AJ5AWlfoQpq+xerfzkREvHUS6w/Pm9+b8t5bRhM3QINS
mNH9PzelMcmi5wD1IMy53NIRfiyTOYKo6DQj99mFOzF3K4pzkdIVKRGv02UH
gQ+APIP7oIVCmRnlTiRhk+77cfRq0ZIyu2fa4wq9oxiC7S/iA9mAhLO7UHa0
pWrxcz+avCDnyHOoGnAIiajCLOnVwVxoNATxXP0L02/r5dpFhBlQq+21r6KT
udqvV/RwrJYHckJzdgAtsnZg+crURLQlBmCixtl+TeLD2dA/6yrKB9KoGc0X
364HD+Xe0WXV8jldV7sGbNIdjRopDFB5mIROp0DC6eZhXENZjE9HMUXIM37y
uI1NQUyts0ISbpTk8x61Xh43sDUV3R1TfoJGSTMtKNtKMmAcl/3+7DT/qSJF
WyFT6DhDD6LAQf/qdTqWVkn4ENqtXYefNcRPH4H8SKMGapK0NULgZXzbtK3H
PfqpImTufzW8mx/h11GeQTPkV11YsQFUdfgHx2Nm1vEdPHcbm0ho+ix20Z5X
ECFEKhL9GmosJPUCSLwd0FjmCMkeG7DUsquSO0xfPPjRZC3L/uj8RTQJxmV8
mWraFZCQErrZG7gGr4sQQF95y/XuJm93dvXXao0yoxqGHe7Vr8hoX2rmqcWa
QQsazf+DtGwmL/LdC6FRdL0ul3DiDGGIzpBsPYh8prVgl0wu1m1s95ZqYxFV
34L+Nekp3IxGeA+2scqwyD/lfb3p4eGagS7Arc0LzDV/UHuWNNoFioKJnqE6
eGGgV3e4kK9Ev/U6t3kh+udFgUVfI0RzkJHjTHE8kuw+LIajA3Fe3Na3/Rpz
uuh47+BX+cKrqxr8c+JasAmltm4VmCVnYHqU83zWVCikxq3VmD1lePRGAYSF
gBtDyOykojIpWl8bm+h7A6UhMD6f0LNThoZ3hcgZbj/lH7GmxUmfr5U+RZdU
ek/PA7DJq8k8chLSMLOS0s0WAP/7f7hwLd87R8+WPi7U01iU/jhZouQCTrQt
xQeu3EM52I8UcEloHgJU+3NpXMqfYQdkDa1RfQht/PqKgexz5LeHGW7tW2xF
5Y4+37y1uX4BZInmJirnLM2Hw9e+pkiSfCj4fypX6BbGxTnppZZObX9hhPNZ
IS/una3rMuKukbl0mlbnTlD4RoZn9Qb3Qi/pwUfL+92OH8lkuJ4oKWRh6WjU
5cPRRQKDm7ZS4Ycyl6Ya+pMG/nOsT0lqtSFsJ/ZGxP0J9a3sP0HfRVqOXmsP
OkHATvRl6Tv7oaAr6zz21bszKQ6tVA21bjLlmWUKBg8CIUoti6rjvNGbj964
NCe/+oYnt4STiPS99uebaz2lNUyor4wox8vppybFikkv8erC+5GngYOwqIaH
AIh2fEc5/Nr7dYWPLa4apc93nAKI3I/yhpKksiRTEEIk1uiYDDp7N78bh7pR
K8PxVkgNpfUu8B0YUK4lWo4TL4FANBONmJ7o0yYKfbuop0JlCvZV+A9Spg8N
rjY5lMFfBCC7OM/g6OrgD7PlDi7/3eAkOXlICKVqG0PiTfnR517SRjyG6O5E
wFrUjWhzWyQ/5RZ/S3dEJ5UCFeEHHi2pg3Lmv+PfriqnNEG870Tsz6hzhl8r
C01v4XHfXnKtee9EGZ5pgW3wH4deuVxTjwitoRv1m1hTzmAHZd+oDg3551ML
t90WjRq5I71hBKOvD44AJtYAOfraA+js5sj81yTkGTmm1HxAPpv1W9l3jdQp
msmtGZydsVVPHVsyzAWjxNOzpX7sC46VhDOJs16TVcnxI70PFETQoH8tOcSu
pBaoI6rcSe0OVomk3UhHKuRjB/aFH5wyvVhbwYzkYibie+CX5TCExMQj+7WR
YvWX+huEEXXQJddkgjgVATWABBNm0+43zMbcbL13g/FKFgXkTroSJw5R11yo
+raYsxGoWKUBjKN8Bz3YFOWqtLldyIoSLLfzGGMD8n/nTKXXWehJU7AqcBWL
4x0f1u2Sfty/Yio1kOB3j6dF7mV9tq/mlcsa+KGTLJWvB9lIn6IOjLOv6yae
k1eh9GGQOYC9pHnr5vlpESczBgjeD66O7GNlBv0YbCD1hlqaSARUPcw+GWfC
sZs3Iu8vrs7ZtKHYiQiFcAjWT/+/GPkWBZqGXbqZa4vfL8MDAmtdCgmg3Puo
DjdcTAhahK0TudYTGoETLK6Cs6nxow1XC2TxqdJd5/l57CM0tQUGzq/IpkB5
f1qMnrrgqMo1GhhoJosWzXLN6fjyJnIbCEU5JRnnCKpy5Ol5HwJzBMlQSVYv
jMVelpY/fT2f3qy1lNrwDuejspY5xxqGDkEioAjwxHiUe9clNxMOZWjx6KQr
4DcRquNbu5qztFf1uM583CBOKiI9Ul4mi79sBCtFbwBpQIkwfvwQx/0U7FL2
mQn2t8IHWpLFKF8dH1ByywE0qsBwKI1/mIAZrXtXUEpMJVnS1uVW8QSkutox
6DNQNNRccCn9+m16NvNxDE1u6gihWtiveH8xEzXNMT9FV6Ai3FSpK3wmEWzS
YlgrIXu/xE7t4/cu1hMH9PY8tDUCfQ5xr6VLnagTAFIUaKcJ3tORaTjbhwvH
J178hCwJjtJFiy1iRUo/VvoHPdgRL50vCK4yK5VHJJBeQYOhwIDXLy9zIhGK
yLzpJKbXd0umtrKeE60Nv6KuZL3saea5YMUYHMbM7hMZS9EGaViBD63UtUpp
YyK4PqzeQxROt8yQYqxO0XdM77cmiEdgpzESVPtHFzMAXCwYuOt1aOh/Pj8J
QnVGJDpNwvCtpUhm9yc8oORmCYZFxFi9vPUplM/ODs0gbAyoGZYAUIiW6ut2
Le+wg64q7kXRlGvI5uQKhD4enxp+uYGumZNKWrbWJUrAFyi7BaY2D69BZ6Zw
Be0i2freUQ6fdgwwMatS/pWvNJ3KMO573kvIn/CeSUbX2IyrdhBSvRRUTXKw
kmZq9fEsPv8Y7YfwU69y7JV83sUzhBIPgHSL/6TXE/mn64mF8v1+AzUXhZNm
eDPJcuo0om60AjArGftERkG1mtWHtV6r2rMuaHmwlv0+5sZ9B8O5zz3oHg+P
tF/4zcFYC3kSaipYHYdnh2BH3oCQ/RYPL1rtzFbvuv3hBTfoQOm8iKoVrhYD
OAiZ4Lrqp+DYZLXgDwnpGmVoc8d5WryEcq8R6G1ikU+RKHi+ldhS1h6bWO/G
WE4ofnvjYj0jse7VqFk0icwNS78YEy9xXB6FhJP4LFeeprE3zSe8cDtGdWeo
2FLHidhhBnrMGxm3c4z9SzabdxUFOV+n9jaBUAX9ZXooZ9vqbTWouuE2D5xr
rKukAz037ROY7J4OtGj1wyh8HoHR+C5jIR9hotS6+cp3nf/WrOr214zSca9t
B02aCAGRrmTCfA1fuhVvDPeO4OnpYpvLfX4qwuTuZX6Q7bpiK94IpB5YW4hj
eqGAhqpqe4D+WSzVFZpdOnjWCoFtFu3sExQWgaMSJSkNghw+5rafC2XHLDcd
ccw/YFDrACjXg5gtoLrEzgDBx5krvyPeJqLaKMiYtQJznrxWQbpFKQFvxtZO
5dwXzRloSfY4vaX4zAebFSMTBcd5vxfJM40FF2q1xrmyDUm5HM5oIG+ZTOOa
4XX89NPERI5Haxh63wmaqN+yzWioZe7KEqzqbOi5QIUdxIQ4C4V93SDd+kWE
/yIbu6Jn5i8j3qeJBleZWe1ozd11F4RTnJJR76wVROdAI2pI07Cy0QPJNmCX
9YfcGWvH3tJqFLMReWkaCvDIQBrDqoxKIIc+yaTDW4NlcEIeAUUyzckof1bp
FO0PPLMeDK3ByPZnnnqT32fjbjqWh0ho+mR0E5A4avAfb3xObdJOg6N0AEBz
360b4PccNIszYMFQ+Vxf2hR+hrvFM1kDuXjkEc+1rtQrXpXgRQUTDxoHgY7l
KOUMmwmDkDoByv39uXr+mnLOropsq88fxJTEbL97Bos4siyg9wsYQA2e7XZK
CLBUUAh9CArSmTKNQfQvAtSKNt7bVve+W/JokFUJ2X5jClpipWh26Po3UhEe
NhXHw1T7PfrmsPinjLeH4zyZbBicFMWbHWqOiJUJI6+RmIEcbLxehllgizVt
eYiND00TS1by2he/uzj5BLKlMxJXFxAQ2ugJYf8b9xhCRk8qUgNFXHj70WI6
Iv6VBnyBapqsGBEcY2Rp/RsMb/URer7p0EAgNbTU98lD3izguECaLH2/dOod
/VcjH6evABXeDWzEylOS5ZY17xKuBEKzbkuFmAMnXEdmtGbV2LqgkF8GqJnS
HUrepMMSAiTJ7FrKwmxyqskzJeqKtsLoW5/FbuloEM0Mw+t8c/MIBmQ+HS7b
56FCYpmSLsZ92YQnt6kod7dlc//+QWTsWayclJ02nkCo9/gRWGhIU5L6Cshv
d6ZHloXxBfDjuwUts89ALSFIMwahZZVikSRpZ6z3j8qgtRb0PNi1GmEK5+/e
lvP6ddkegtNzGJL7xms+8ourmHtqyJZkZUCbI/LtmkTeXDkyAeu38nj3xx6N
4Gn8OESTJZ97XSpz396pbl0RCFqLNvlPgsAcmhCrLwlm/eZ/u6jZv4d2hOtB
5J+tzud0rsgoVLZkQf1x0TU+mQXZNytfWn4WMzDwdliJKFvWDZVkq1VHJZyK
k59Vf88YpYcB/fkLK/+3aOge0FYJgWxsVtFFY5YER38PgsQrOZuFDzuWUySs
qM64PxMYbG+HInkodL/EVDy+d/ONPV2rOofkRj4Uaw2LG9YJPJcmVqIYxrON
1Uom73fiaUAQwU+EIN9sgj1B6bto2DU33SDADSqkT8VAOOGxPTk3VRHj19Ko
RgKrlkMBXnhrvhDxogoqkaVqkGe/665fqWTQFGhFJvsUPy4Ssasw0BglqnS4
O3Y3sGbPpHd/IMFBVrVpIcf7mCUdOjogwxkYb0ekbyR7EsUFWwpVnAsovqct
Zv2I2uUeeDvedBKNnKCqaTzcZiktWXhIUeyoHx8AiBIVuiKOIY82R21RPnfD
pq6AqmpB+L0xZP4DnIckJcP9ZgoPx4hLWvtmSSlIDnCOPS2w3YcDD1sBhCg9
CS2KvB8SWKN0KVS7EclAZDmDO7jf8uWoul9+XoEqnnawTSzZQRvwW1Pfmy5q
e9WrC/uM/IrN4D3Y+TL8StzTqQkvhHcVO+mYMJ0+KtNLecn+TpRlqeEDCU1u
T8owC/h2SVqTrfnVasYV5EezjLdyYv9hocYMjawVAmAXKfyK1KOAmsow7xrW
VT508jsAGpS4aMs7wjck13olcUc4Pz4/I9nbIb+TbAqP1Gxwwrbuu3jktFVw
QxSvfUN2fnKzYBbQp+sa8FVda1T5tmxofVb2LVGJvRTCgge+kfc3VcKdCn2u
/UtMORezwjE6qw2sNgdTAAzmTDdROKhByLfUBEBPXaPFBEnuBoBGVg6ommNe
czkUyxgVy+3wl3CCH81AAdNTp2CiQQcHqvdfmGNH26Ali/rVhyQEG48iQlhh
9ZI/f8oQmDsqkSk7AMKmIop4w3UATazvDvUhiDdp+vMD407OGLChnLla3oUd
n78rLrrR5OpEEHPShemfBryIaibM4qkNAslz9tsmn0e3c0d6va9fCnzSa8BM
Y11iNKzJ8L6ELADLGZaALZE2/PZQxXhXjZEaFqPr8oUWoMLcGliBur8vGRdG
VYg+lwZO+WCPafICTNwB3283uAnKii4kYNu9btRhjcuCMMAUv1gCMpbvjquC
DTsId1nXBDUUEFx0QOqO/4yF88I/iLcEK4cXaoamsdXB4D+MelybEUc8Ni67
SBo1I9gSoUB6LIOHJ5oV7gI42G7DPKiMfctQpFYGK0jkrscQUE2mYQjX0owt
6r669I0+qSuAlc/Q2vLn/uM5OdXXEODInJi31nzo+cGlHIqeX6D0U429GrUl
fWG8gVernqCDuZbrR70QX0BomkXkonIcx8Bdbx8qRHZZHa5f5WyyoCSVE2qp
hzIsk2qKZQivkRI6rILBc7rnEh5zilfBNfMcgvYPj1DHyy+9xz4mXdpp4KGC
x9eTQ4ceR34ugZ5Xt954FXp3/VnNsUzV4SCUyd9jVByfiFG0b9BnN6WAYjqI
xHFput+VDm3gktRVeeWFsjC2J1OZcGTVGxqicd38DFBugUh+ZBUE8DCCUTCh
AHpG1Dx011+hOOAaw7i8UxCruTai2gPNfMIUeG8EPPng4euKHRGv6BRJNigM
KcGqm4bxQE8lFwWk1sqk2mrCvswnraQvtBPE3TSxImQCFJfslFROy8c8jYvt
F/FFnFHyll0B1gbVDQ8tfhAHVGs0qiqyO5kM6ew/f6x3SQGw6+2UZ/7Qw/Q0
7Z1lD4HdxPYMpFRBGijKH10XGzz1gU/1MLcId4M7F/HLHhPLW2hIpQIuRyhr
i6+9Im2wfuohdYiBgj4OB4zXKoqvGF+OgDRVkTCfj5X6U8VeAmpwUU59af08
+qQpwl3pYak1Cp+LE+XGaizgWyh6pFRh4mdmndFOPYeM3d6tHCwOayUsO3A0
QMKDU2BvHAGZqf4qBYab6CyOzC0GtRNy1ApVmAPfwZuUlGLZ+0yK29WzGlge
fFS/vRO2+qSv3Fy0T8gYh9Iebl4j/jOkERz+ZuXYoaXOlmYCaCNfxjiZP0zB
3HGOLsPf50Ic0oRdUY6YIcqG+ONyS/qVy2RMJyzn+1MJeu/MndJxQyBNEdtb
OCD5WujReG1EAzK42Ap4+MnVFeKG80itSdDdpyLjrL0GzJkA5VEGjniCEbVx
D5EG9yEHNp+tnzFYACTxWQJez025jzlst0MCBrudMYZKneHwoJ7ZClUi7rAS
TewDUkAdFVL4wnsTT4dHv585d9bK7va0L5PSaPDMpRf553ErFPPZqXc8L6gv
tQvklX8HYQqhaBM5g/eduh+f9ZpIfjfTz6rqOs261zoOrrCS92RVbl5opFvR
IPr7oOOfhu7zm9lrCJAx6/TN8swheXifbiUJW8SiPuFh/bZ+hFOocHZ0dsvb
oEIACJwNkR+KMNctjEhqomK/GXd8te5zBqlt9rJ9d0Bo0rfQBudq9tl0wU7d
L2Ia+bhk3Pimt0t01Wmvcl78sBzVey/7AmkwDHCGJJCxIjXUPx0JmV7u/iVX
e2cIelFtfG0ag/WTyUpm8Q8ZE7Lq46jG9A0UUzZOSlcXooy/Yl0tkko3d/DS
dAA/KLLuDRrX4HNSzkedpJVQyPeddkzpRtbhSN/ijYbXUTUxez82UW3+/6ug
o6UGQCkpHEMHgcWJWgy4vCJNV77uAwfhZmI4SeZu+fo7Dc96ZBXndI/AA5PZ
zbIdBir3L4Q9xq/9ovSnSKERkQ9vw/o9LdcUX36Sgt5qEERv44hBa+lqhODC
JHgAMxqUMsx3uD2xMhl14cg5z5yTZYYKCDPLtOFvUh3ASIpRE8Kh9yHdK7b7
6lxPDnmX/MiJC8j2DwuTK/24G0g5rg72yPY6A/7s3GX+WkJsGNqU3rIWASkg
hC/LVp5vnTgcYIiebHc2EAnSzUmYwGo6bsry3JHnHKayRcMQb12LTqRJZXUc
OGJJpWE98Cf77teBgk93n8gnmYTcICqCTkOhi6sZlOz0LkaHX7PxfOnozjck
BgCGqyJPW7/j5ry47a2YKpM1EGQ+NgwSwQ6fwQuSZtXh9vrpGEWmMoWrphbA
AfC3W6rBwb6JkI0HdNVRP2QXXNwtV3dhal25M8AQjA0OfHSE0VM498TRlDW1
rh+PTQUtwtOdtF+9JjY7yTYuvtoJ/48+jDSbq7sywOxnXA0FUYlOhQEoFlfi
iqqjBEf7rGFQs6kXm2XETRAlfD9o9yJd1+Nuh5ACjdOIuJM3vN7rbo3UaurN
b4J36Cn1dRrJAyZCgGn6JGgqHfIkHIoMNETlwPuRs3WScBYZ7V0lVVU/QGZi
V65qdEXFh5wD8v3bNMGwYcraJnSBMrR5E/I3RLCMg82m5vy5RjF1TLC6jKm1
8bbu+Hdp5Awa2V2jPa6RTk0/hy1X726OttK2RaQLATFxMhu8cqwJQMLTqM8Q
wInqZyYNde66pZaxoPSMDl/KnlEbW8CpONGEj+1X3qad8fuovcxoIPY/dcwZ
u7MN1qV24NsPrH5Rimmd/3XHsa2AcGjg8kxKfqDYeY78LvqrSmvtbMbbeTWD
cQNfNFc0Yv+QdoeG2du5Ob/zF2bMJ4UsSdGaQniYLXnBiZu3AX+ErlhTXpP/
7+LRAE0wgQrRn6L4EzovuL7ei03zNLbFSLrV7bhq8eWYjGJJjrDrMQaT2pMc
REW3/TmtclSR+64JPa0Mkn9xIut5ekYnQ8181YBnGwLMBa4LOD88zjkZOIul
TRJxLTmUKypVUan4j7wTAl60I+N0FKYs0inW3dQitmXCe+iojtlnaFagccy8
UCo/83aIjJ8Ex8e0dHsSgeylSI/HEshXQ+58r27Ktz+XB6zC1yYC5mkkkFtd
88EeCU+580PWsvFz3ttCQORJELCf0PYThOwumkUPSdeRH6uAtAcULKoBn7y1
UzdmqpIJFLCkm1f3OoFGsAxtUt0/ihNmLNVsyuSDKxUmBhjFebR52U//elHz
n2CeEtMayYm9mXnouclQQ5l56TmUQL1jmSsVlgdIEM7UB67hVIZYfIrNkPTf
jKEmhTlTsRnGhyEsUwnf03QKgVmbAyO9OaoBkNQ7TVQE7U0H3X3lGKyMIv24
ZKyyPiV+rUZKGmKVqjjpc1L3IPFueq//JtVwTMxeRGX0+a+n2jiPhYKrXWvh
pkQXu2LrH4/cqcesRNlxAKtgmLRtQILoyqvwQY0o+hC47lmw0SFR10e+g90D
oEmNQ9uq0dJXbWoHzrgESBImbt1VcvvXWoTa0SQO2bRxj49XAMDKyBhMSVf1
DqmFO1Rhbn7GfKq/7o+Ym28yC4I/UwTc+YNLudy+LN/w/jvrVvHx1iq1n7i9
9qH5OTh8bntVEGOWXxGPwXom0epJfrHQ9R+CxN0Xd9FMtJDTSavLcVcz9jnm
1JhgKgCTvubzitOl4mF4psMABn6qbNiCNj5IqisYaAPgySygldHV/0xRo8Ae
KmjnJuRmB1lxNugqf45lFIlCXo3Um23i0lORWIIozztEPf4XKIc7FhRFj9RY
AfOYa/ALNz0hW5SzMPgI2oCxyFGSrQmhezg2rVWEJk5VRQmfdlUkz82Fj1I7
KBnH9Bpl3Txh3x8xao85psSmXR4aaNXQSmvGOrRRuHAQiwxE6oFNRTpIiKYp
snC2Z+bYwVEMqqhr3vezCi1kjGynn/y+1XjuNoykGxRJITbJaPzYCMo95QBT
xXqR4hLtWfDXKUAhmIcLeCsqEYvukt+2vx//Wa1FqKLyU7nt+ANvJPUHB9Iq
LXTWIcMQd9cKijP0xAMQF1LK9fi0Fn+GxIiT95bqeVuQiuyQ62I8FMpo3fOO
XW4Hpm0uXJoYCh0X+Lj4bhx2MPPyulXeDO4YzB/FJHFplYcTjiJxMQCeGbvK
FMr0yfQtTvuKbQSblr4Z5ZkDRODQEDbeKFn4YXdcLiNWPCwKiYH47hv2xrgi
zGmZmbu/JZY+hIGYIEV6nODa+oE+XHNEzm2PDbOAlpBd3y3/XJaThlboZGwC
BRpvpGQz7Hq37/Z9Z8Z3UP0HdlzjN23gC19uL7GjmVrv1z9XtCKb946OKdMT
tsd5kkr0N30csTEqfJkyXd/d92FuHUc5TAVjQ5kXOsiBB7tviQDPTGOHgvvV
a1Z38OebYq2vNmuSZjQn8qPjFOVzi2+b1B6TDMlFp6q0SkuGtGEs8qgY3Ts0
sQmIkTMqWhAFy0hcdRrdaQfxqchhuwkGG0Sg9p9m6YTH3yc8+TVpSxaO9VuH
3SQfzOKNAuENCnAaMIAfxuOdNeeUvukDW4mOL975asKP06NKUSHLl8JdRi1i
nHm9FeqV+AlhlVOemjX/TFKRLS5Pe3/1b9ksfLOrx8Wcq027jCJ9FsS+a7at
XBynb9qor2/rIPnnCX9cvG4jPU4iodCDDrwp88m9OaLFKXbjPc2Vph5DpU8z
OVKZeANaGErVUtZOvsJl6NLBBXO4yzIwQ2WYP9qskHP0XO2eyM4BoL6PeuNu
iagBRS4/x1dWzw6fVHFy0lv+AJjRebcgiqCKJJnnuvupu+X+0jTjIcMB9sv9
edQCzcL5CkeShr1ZyLDey5ukyxuy1xs/CwyUmrYCx1xNN44jKyYhL3+QPy5g
l82w9+VeoO8AivH+sWrL+lzbO6x5LjnBKUNZKK4MsQSz3pHDCFveT2r2dvyR
PJUhxVXvM6avkPhTspCstjDbUa36h/OGqyg4N/oT5cO2B33d1D6J52O8iaLd
5XArEkAL1hWGoSg2smLJE2/vgoAF2DKGiq2lORfzYX1+bbLxybsmiA9Bm3jO
vJLsf0b2jjQxD5AtNDnBmzKV7zVPA4d4YFDytePA7OjdAlPyBJFD1OYQ7J/f
9UtCes0K9rR5S/Bv9O68WP3t826CnZFs5SBqPzFapE5Ju2Dxm4tWJDzC8bpW
pljTaVL4QtO3LFZeQop7MPzOckOoJv3q0c/dwb5HXxPfJlSs/dREOgW8kOLT
aN6moGJtEMAlQMn/3xafPfGQeIdgbPkhTIIy3pITUAgvKrFTvQUbGXrn/Brj
cTqueB+phdDiIHE8cuFi8owjp0Qh3dIaIv21KbJBwNFjWerjZAPffzaWQ3M8
vP6BhH2PQj4XgtvncPiXrb01q3xaIAFu2pTF4S4sm6vi1OdVGOrO/CeySLMj
ZhjooOYdmg3Q7nuiq5N8sUaxsviAFX8Rtx7vShBmztnxPO8ZOolmJATbUmXr
Kl2h7SSsWvtkUetN3QQj4CpyRXwznGTJ/YTVEhy3n2VqvPNlj4xkd5dsi4e3
jdW3CjGoDFz5FRAVBRgpiFjij8Q/QxZPXZI+OVe3jDBLChS8Xy6EYdwkg7YP
RzcsrPJlPNHCXWlScgRocZDWZcQoH0oYDoicKuhwYKxrPPgVbl8PKezhAP73
cq0T+dzGbkVQar7ifCPNlieKiaUBkSzpzDB0F7/OXoN7f8iEWKIx34HjYHbJ
l1Kzvjkcvcs5dpzou6kdJzz68UF0+Oo5vaTje1rO8o5oNn/cCJ7/PmYthPZq
93v//Z1A8vtxAVaDuxWYJcz1NOqF9v9uuedY9FvjIQwJy5FIQTQnMZE1tMxE
EPIuUB+qfUERfIz+NsAXV6zJsfVgidoc7DhU4hUdq+/N0kIkofND+C6ZBeTq
AVoGkEOtqllPpgKxEGBRfRRYsm3xHr435F92fmVxHxE+lkxDWy8vM4eLFy9L
MTQ+PBafWX6qYFW0ny0qMzcjf9lZEEXijsllKywfxi2GXBW1XgZ4Hk94FsY3
CwWU6JdencarGZ33E1DQpDHJy57bfDUYS4AyOINun1PtGhHg0lQMXczaU//o
P2MPeNMXzO/Bb7+ebjBu4/CzxklEBowWvLUvmls1tpfi4NiB35Bcy5OJ0SCr
uvQj2CUodnO5T7qPh46FMdIosMsqB3Ra9HjPn3TcfOnv0gka1V3cq4qXTh6F
oW1e6RMO/cgvrXA++n+uVzrrQgZjKNkXMSu+FnB+2IzNFm/9cM0PgMO3dy7q
HAD0/oEWvGBFiHSVPGwW/9TcG6SYhnP+MV+KWIWF80Q23z+Ej02G+g+GFyVE
uoXTlvbM1aCd7HPqms+EeG8dijBkpiilCRsmT6IlTej4YXQcCIuEIn4pWqeD
QT3VYErjG+5FAuURUgJHmdBgcv7KB/yWEbgBcr8fgvHDsiPLA/y0T57n1Drd
0UWsCDuVQHaRup/xwdHAF3iX1js8J+B5Qezwr83ALRWjXTrMTpmeLH4mx/Pd
nZ16qaYCbpFFItc3GycQhkc8tPamZtXSy7LcJKWE1Awnk7iy8IPhEH8KLZn2
0UtCWIQ/BdjQ/vYsLNn/3G59fX0/KibP6QsUv2uIoxT1keee6U2Z3+Bn6iQ4
5T1wc1eSq8J/KoHnuTp6HkhsVaeug7eaz1RjXY6UfV57hmZveCdwcyyZegEX
VIxZuF7QJ7y95hEEy3qgnjiZ7M5sqf6LGuh4iLrVHuEX1msNuAcWozMdGYZ7
ditp2Mr5K6VMB4GNChmSKLqk9xTZEEK/t9aYxjMlSkC9B1gn34H7wcfnNYY9
xu2D37iP4tCA94fQ1QJ9TttkgFqbRU6v/z3SZHdfrOPRBRnCst6Ex3bw3D2R
SjU5eAlBNI67xL7Fg3Cp8ZqEVS1ST4WbQt7OLgTzfAz6NLXszuXuS3s7hFp8
OPA/TFDnGoK1iO/AMnKB51M/3IXkQx220QSVD/tfpHrbhP2FUn/7/M7QBjPh
r2U7KlGFyT4jUditnfJFXvV5lNRx9dfSKI8LGfCacJyUUX/vIoWixVWoldvx
Tu4NHoPxuKnqccsNMiHS8iOnM3PPY0Vdi5cEXveLNYtiOAPhMv6dT7CYbx0x
tWIqpD2VpeIjs8ztogu0CNTymIXS97Lemoh1CMJluAZIfcFvmIkTWCdy2wf4
ggmOz21CgZMPmR2QOed0/hsGuoX/l0vU9r2lzb35jYAAW12x3FF1o59Il7aT
o6HZWctbgwFPbTaMLu5/590UwMdcXc1NXTWzTVzT/21PJcW57w5L/Css+6Le
4SLbk5J4DBNlaTHFW+tytYCnxWT6dgK0Vd36hY/tjnwng/Uw8lPu6rwEzCB5
x3bhOpThCSbe1rATVQ+avEMk2xLyTkSl5zo0vUd7+khVP8Dv8ot7F7YAMbpN
kW72oTUAFBlSsjJptFgs2KYro4Qt71P4DJR8DQriacfV0bA28avVmvyLLCPf
CtW6+REEgwMWQhlf62yr0O0GXSwE/dBDPoLscn/bsDtZM+5dAxFTELWyYHqz
jvaRj6prhz5VCT/kDuGoadqNzLoNipCcgCFf9HxSO1taXN4/w07ARDM76YDI
72FrPc4oyYoJVpHuD+MAlJLPup6DYACsdnqj2lRGKlHW8KqUYEKUCeiHMIJj
GQCBaHVRuqCAL77ftu/c3Xz5l4Bi5WqnOqZYGQlrPF4Wr29NF74jTH9ilIeF
Y5dxy9UQ4gFdjLXWb5KzYsM4ezrW4DHKXs4ffBhSwdX7XDxMqZ4KRSn5dXkO
c/TsaQw1ooxhylMJDU5xoaunnqlKlQw8K4lW7euUFf3IzCiDfFdFYL0rdxvI
giDgA2S4oetBjBWu35z8jC4RPjwgvt7RsZuACk2Azklom65we9G3m882fLE7
e8Aij8CJHec0LTSVscxQEuBtxJJgyLaLOG06OUbS3Pki3NoFvGi5g+1iYVXS
Kt+KlHMJTvxY0fK4YaOtrQ+3CRZzWGyB9UTd/1EfFdq97wDLVStAC1XfhWbW
U2p77fJwd98hyCcBzMpxmp0GhZ/1day3HKfR3S1Cngu8FQOEXwHDtmx5mkI+
UHvRyc1wc3Ph1LisFMyVrAmIPYG2WlT6l2MJOOr8Fuppsk2B6B/4TKR17BrX
QXrm4oIK9xzxvkPvA161ziQW/YiTz8p98TkYiTMqo32Z7jWF7Ia5Kkyvl7N3
TnklqgNV/85kJldrzVBWYqhSlgfiM7EXZH5nuepdI0CCBFOtUbcSGdK6/vqc
aeP1EnMy128wFiySt1p3rKCuG5DTCoM8lLm5nQ4xq1W4IUZyFz4FLspPD5vA
90w/+aTROf+u6hA6X2aiZJuDxObV226l6OK4120cCeECE6xc7dEv7qd39lk2
PLVOHeArHiRvWxWFnFKX8JbQjsTWjvJNWH/8WSPGGOnzMf0r9c1gHGOe4Hqp
SyMQTIxRa2ngebxoiEk6+hpUlDCcjyPMUKwAR5omS8KsI+gJWR095oqL6W15
mnn+f1b6iox3dOFkzu9mCFXYrPQzhrpxJ0bDRgo/sqDFJgx/wYIpQEDrKdoK
NqJEm3S/DDn4wQlDuYJgyFiBrTlCBd4k/HVYZelGIYyV1dIh4ZQBcjnE955a
BM9UYm9uPOLv1IZw1lGRKghk50EJr5pgrOHxf+6opz7x0bYCJT4Y/VJ1qesf
cwuWogb5QRWH1QZMGhcnD+qJTUaQLQWieSEKPz7T3SESbq+Kv1xpdjvEKApL
gf+Xn1/JcfUKiJmWbBSn6VJjrwGCjyzL7vDTDr1aExT9+POv5k5US+HjbzpM
rAjYBA0HbblFQ9T06VHizrRAlnQoXtPkx2Po39/f7fw42lDkEA+02XEX/sbC
Zi5sFnAXhuSq38bzJgoQS6hxX3RMlbj+tqg1qadXFH5uPREKGEYsNl+D/AgE
muhb9kbgTvVO9MqFPICnk9nP3zEIj++Kewjo07h+ZFBuUaRF/2SNGwC/S9Vn
gfqZ5Z536NS3I1fp8drluBeOKkCA2sAAW8DBvcoIY3FSA29GSFnBAF/A45dH
UeifcevRtoMjeZ+fi6ScITTE/l8J1bslQnzuc2Zty6fCp43qyyUe5PprHsXS
2DxFta7cCNFaTSAFXwbVhmue6h78vwDkB4aj1ExIFy/aIg8kISyOcp+hh0LS
7Ipchh+4+Ny7qbHi7vpMM6gDyl86F/YS4xQmfTwYFYN3/Oxac02ZseWFzdKH
hZBUp10N1qAc7uemubQUCMk2aJ4mXpsygxTiOtsoXBPivmLaiAvldPT2YD0V
Di3lc4WohiEU3tzMaPPJqS+bZl4w2VhE38NB2Ixri+uKdrNBU2PWzSkoMB4j
ogm7cdGx6PKw0ch8xzyrDM1KPtJA7MaSDaE1ohvTRVYqUnJvlWQPoiEga+qM
QNG0lxcevDwYmwZmRUpIKIJsD8x5InN95WIwtwsgmjayrsjp78ebD6K0bbPe
mcoQfiRX9HmUSsartfnb7KfJB9pgPcbT4TOQodQmSuysvfnp6nnQYgU2E4Zd
UXmYiZa61y9tY4zY4k+OIZZYytTnNaZhYlpFMSDzcrmkN1AyEA7XCGi7j2F/
qx18284u+U4sg50TWdatbJppC5DC9DCjfQ7VnWw1/6bS8NSCIj7dSJV1xVJE
0f08UFyEJr4qnww1xuKGsTiFGCq/T7L9EM9PfE4ZFdweizT5DMVctEgzndYG
/zN7S7RX6LNu31PbnEM1YZ5uWEx28ZIaEUhXZvq5V2b4Nc4nL65Wpv3j1gif
T06kjMoyq4TwAeLU345Px6CPkZdYriI00PjEIhjkpuoDncCqmdEW4f8+hdHb
HFnnds8fJ1JJXotRDDTB0wHhHGyzl0QYkm6EYsORcx8eByIVmoZ7XDaWYrZo
lebp6Cs+O+QNBCpZVIBBIAFN7GDOa1pR5fNnfBO46sRhLVEv+eN0nYwXciFE
J0sBg0w+AK4aIMnJwxA0yoNsOy3ibwR56X63HwiI2lxQauEb6vx2lDrbcpfw
Ena05ueX7mjP6MRc6/0mpoRPyJXXg6TQmK5rHNzJ4BsTKwBU7Y0xyuvWaQDm
8rgtwj9kchEpQ5Dn891bfaaAzNDjvyOvE/QKGdhQkB+Dr3Ee6qeRofSM1JDX
d6yPp56SpZC9kOVw7UXnNPdFSy6UiwuIG2360dbV6BO27zBA8TWIdzTMqNO/
gu16DpG6dpeo99i8q/eCiqR1OsctopJioWWT21bXxHuUDg88J7kX5LMHdwVW
fJYSF35uBVDaehgv1vqKESc5GPomLFOJxOFRSDVCM3sVmbZP9B5V6VEXQa4+
dVJ7PgpnOe8JQNLGhxK7RkY6NCFCO1R+fnLxy8i9+/xwViqBlyiIxF/Ecee/
SaqRcVMv0VWowWrGDA5WxuRmgpKGMLIGSosGybPpfuEaepbURKPsrDsRcRyV
p1Ae2EoXXaY+F+ufRaYcjhFQLick4eGfw9U7eX06ssGL8AHUbCgIcCINek4e
PKu+vT0XPqw9qFHsNWHkWJmPPLDYemEYa7j7HDITvzv0I5f3nVW3cf4x7Bx6
HcD5rSSMUgZG9Ai6qKHlEFQOJXri5W7P/xt84s8BRrGz7WiKBEWnDEIab/nL
rWUMVe+NQqqS/384a70wWev7pfrzKA58FnsLfBhiO4TCkZhJSIhIgY27GCE2
6DqhifmSSsvXKJRtaOye6inpLVwJ9Orj0syU8qoZ1TZdkEr0SYKJKjB0/PjF
mRJoaeVHwHWxMjDzqb6vQyR3fnXf/c0Xay9AndkzT8mOJ1CXdNU6GBNMe2SF
V7cnWMDs7LpUk3CAPrLtOrL2/vmmsVGgzOvn0d8Av2zzW+6Yx5Y2Cfe304wR
gO2f98WNAYU6QSmGz0MpJaxZDhgrhjIaMbzasZPPMJ1/MrXyaszGbbuCtzDv
6W/i0bDAonODRzZH1oBCGoUOjQLBmT/Bko/vLapKRHrC7CDAKsRtOBJCw8ea
KJ0aYGqmOlhGqbyHXbevQme/01rjFDCThMFt4Vm3rS5LXZkFs249xpu9tF7f
U+ihnNlNOTygCgXLdNuw0F/DhSAtJcurKFPk4seyKWDxeGJUQlU9LKzxBZ5K
vP+Ms0Swjl+EOCVCE7j6AqlXajJ4sNRSzuCf76SzH7UgL+f0cQ/r3BqpI8hA
9UdG6ujrpTfeRYuHMaRrIwjiUU+l3uAmhw7f4WkZcqeRjrc7rmjmKxknaVz/
m8V1zZNvpIx3HSUeF+7K1nFPvlMy7APH67rNR/lIy/byBJO9xhdduB4T7Guq
hOifDfEzvOTCWS+3OUF5CcFAeNJdK2eoukaoBlqyBAXmwvvBJJu9KNT4kDr3
LvSLUmBlgIR3PHPUxPeaka1nFdmtmmKQwB6dgwPuthwFI/MphueN+IhA3j+Z
2ZeAfaT1SJN0bWpJ0oECjeD7AriLEGZ73RIUKDksgaIiBqbutCku4A8vs1lY
/Wh1YIkJ6Y3ZiMRXnx1d4JIIY+RT9CPkKd3XxdQ8LoLb20OsXi09ndewTO0Z
0lsO0U3oX9MBKmM8SJQN5Jh9mTODCzI6vRg9gPT6dk9K87pdbgVf7TJdQzHx
nOFbD3OwBcNDupzdj6E16rGzkFW8nz90d1szbkM1DCXDXp5DXlnhdRev0GFD
UiYFONOTVQnoqoniFm1cnDyerm0DHTG8cltoXtt2kJpdn68uiK0+U3WwRUZl
gea3hpg9R8GOWc/tZ4jZ87nBFaf39dGcPbtXECrARZ2KS44UMZ9kc5CKeyWV
oY+uf3ytwleeDQkQvzUHbI7D7MdQacTOVIzTlnafap2JHj8a3GY3Z/SYo+fF
FNrZzUDRygMQiKD/ak0V7QvSPpdwg2bDrGu3WlcOVgxDLOKPggvIsfBiTqkj
uDpWE/X6pPP1mP/l5pvG1qJVk9KRIp8FDDRutBGAvQIVII3AH9oTfxU8AjLP
Gfu6fLIlKEeR7M7yJfcPMNJnVJFwtrvYSgn8d3s1v+8+qDXPTSDvgHEzHA13
jyiXGI00AWsRPXmrF5yynMzbxwT326E2Odys/Rvd9O45KnQumVHREvmZzhWx
k3XOpW9/9Ph/hUjoSLEv2eliqSixfNncix/Y97dj6DUUjQq9FQF5z9Isap4S
xT482IKLvjmb228uKmtlBO9ek+g+TG+jJ9ZwTFQvw7y+cLc9cghMaAKB4W/G
2aRlJOIRi26bXiPzk8PuAyU7a4VaGZO1ZO3754/y0qq2H9mrQQvdSWNYH5m2
ZuNLcYtn6Icyy//KHOlL86D4YO8DuKcJw5Oq/9792dUxta7DgP3v/pS2XZLC
OXNF9ldxYAaPD9O1wK+E0yigQ41EKa1f/jgA3iIs3fTRXJKT6MYHhfpGpvXW
K1pOLQNJao8Ux84oHCJxx2kK7xtg2N6SHD1XLMAKwj4owuLRy1aYUg1OJ1In
spo10nUx1YUv0uKiXsvHUEsA+ZNopHztWTxyNkqzNkZDywt4vFQGTTKcaS+e
/Jip2eEITC2ad62oGD3E1VJEMcquVhX7qhgKL0lDLU7JUsoiPSctvwxNTxSu
fS22ecfamQv495Mhf6FWxjFOqtQk7/xwII9uxqUS5jfW0PuEchpsvttTBbWl
hDQUs7pxBVRpKb5EGwesliikVKIILloCUJJvOVU+WfjfIx1Knx5uv3LYTRvx
yOrhcK8gzaERIXBER+g5EoWg7hbg/n+N5DOziw4Hqny0fsi1iNRyrC9OrrDm
JsvRjcYnsDLu7V0MSR3rkDqpyChIVWWjVZjqMzN7q/tus4UnLZN6WsF2u4/3
B8TMEYrHf5hfdjq6hkUyw7UdXMxA/yc/Dq78H43K/f2IG7Idxc76SoQ852vo
ALnaiQUBmn1viLDjAXqHhQiInHJNl88zKrC4F+AbQXLT5um6Ac8mk/FI9t7T
pdyO9qCL9ZUQ4wAOosTa5CbztqnHqCD40FtZoHK00lchHGJDQCB6nJsr+B1p
rK06+i78UV5+kDw3DZq4G4C2WuQ9X6G1UzPtKzXrC61teLWEMbdwnltcjhUA
hu64PGuB1LNhf0dAYpxmNOpXv8fIiInCSeUV3cSPnW0fe2KsrrbkrBKufMDg
xSlCx+c5YohYODIjIgDo+6E6fax5B5UACx0/R8WX5uqN7XTfsX0pEPADedIf
7/tvNb6VvbzvD5VjfadFBjNFmFfin8ITXi8LnKyuyPu7ClblYwJWJeqV/JL8
e9KcK7Og2H8HaM6fLSZMYV8L2fI0lnqQzlSbs41cCqrULzZgLXSXhHKa0E5K
mahMlLo+lZt4zEfWO0HVzAswWvGSV9E495bn9dbgdPXx/+N8bc7XvCVjf61O
pFf6Jb2Y2GY9N8zMDcg6UWuMYdzp5gfLobJmmXzXfKgUXqE45yOU0WOWQUQp
JivrYnZ5Tqr0sP8J0wKJWdqwpZuJksvhlFOALrKKvTZWxIXrRB48C5Y6rYj+
gFF0fH93DlYGEUh5ern8r+xggTeT1QdqTJhi5HK/3UB+fjTKU/Kt6EUBNkA4
V8VlXy639xLv/XT2ZXu2xdAhBV7+tsXYr2T0urCFWejcswCk/FD28cGFRFV9
kgUAKtvl7n/ubKF5q2qXFDW6NebfXAQh8F2CM5Gwc0tQgRNkpt+M2L4po2bN
7iMGGaPXLunUAd9S+1o473p/mJpbDVOMS/eSHjGSnn3qzTgDeoZhz5cunAx7
My8wstYk1ZkkLUoL1jQzMoiSjV6fRKnxKCl11D0CxqxU0dlJNoC9M0AT9PU8
XBnal+7nkdQZcE/noch6DKs697PQ+f0gjI9X99fcCxWL4adE1MLVHaVskg+Y
/5RTVbcDj39vxujXCF6biE/+l4cwLLKOehRcSCxHAv9weXtt/piMxsqNNKjQ
Zh5F6XLtQTDSgkQx5v3BewchC4ftoJRqrPL9qW/4vZ9oXoTFK6FmgbIda5d4
oyvpnNPA20P9m1NwS8MrklsIJT0PHsL6yizOZJdSIm5YEVmZ8mThdbp6P//s
vBn+Mg3SBJDmi2T1L1uREVFqm0uIbBCn533c79G/9XnvgqIKG5WEN+pilVAV
330uBBrXa1MYBQlTcJfCFt2P/d7zWO2fiGkikJFcyncmkJOKiSyye3EigTqz
z7a4OhgstTFwHyu6y9VBucks4trTu2FiCkMin+sSevc7vKR0FRo4J8m5r4Bo
z/6Zi3kHI9Z7zigbHqUI5PXmCdOPnZNJytnP5wBTYKhL/epHtVvu5Ojfvs6Q
Rih68FTqV3O+cojoC02+KQflu6c3rSIeocCvY4EJKVjA5vy7PEUG0rfw1fTb
KFwa2aWlNT7FBOIB/AyGqnJdtrRYT3Sl5M+mt3AZz4N5fk/KkKXxnSXX3T3L
mticgaQsMjlxmJlM2qR5K5THQJ8zM9+cB8cJTPZtuzbWZB9xBNqqmTq0dMI8
tas2dL2wiRZjfx4Yd9O3UNnCYPrzEqLF2IDkI5LTkUzfysrOB37ymHJlu3oH
yAHDeurXV/bSnWruPLkN4o84XJxQes9TaR8oFnWN6HNa3M79yQxM6b+DQuvH
I7t3gZQ+gQKxNIrhZquQrq1or0/fIZMZS/EQUesi7XeV4B5soaT9avKaalHu
E562quRIjKCTLqZkbm+DOqaZYtwYwiE7K0nmTUg6irBL7+5mvjQ7JT0zm3hc
qDmmOPFvQektxNIE29hlcBh3l87JccrFnfMAA9H+kR2u2F8dHJR1zSuNh5CD
NeMDZyigJLGdHmbmB2awE1RypDETpQenOLcgJLpNK7lnvSS5I8FwQWWLU/hn
5A3DIGpw6LFPZr5adwkJfPyf/+/P47MY6uWGlutFXMwsS7g52FOnXKGQpOLX
PU/bcoACOe+Vmzt8dDTUshws6XbAe5FKkIQrRtdqkThNyad7aN4hXipcuHRv
DididUTIc9/OcqTk7ZPqiQuAUNdRPp26i3nKtlgsz9QXA7ejNoKCYNT80+lA
RMpcjMqMH/kSzcZ+kbXZxNar1zCbOOrkSatLEAUkDK+amHtxbhAfzXD6VFFG
AimzSwTw8+lxI37SW6GiPqhqG88FSHeOX73wmcr12bPY/z2Z0snd+4jP3slh
HW/DbNOz7up6hXoKYB4TABXuGRtwlvhVMRFvm88TBS2FChHmDVvyF8Fn5nqR
fxmm2BSBR24px36AzWGKJD/G1f6sokXiMjzLBJvHWXfkrHezBAxeHZd3IxzK
oJugvMnBGOwu4mzf1fNGm1Z3yRTLcdt4EjrVRg2cyIGNh2/Y/6FZAEqWrQrI
VNPpNuomUrx+ssVgkgui8bfg/AmTwos0D6ARQQMQOnJdu9/FyVvD6I3CAPIZ
HspLiEuafvkFm8srV25skM8m0SBmYaZSwMVDLSsenhhW1nAhC40JUV1zSYCL
M4etq0EKdkKd8kZwe31SatJ+T8QaDaHA+7KBdipOCffqdxf8zn7wT5EDKi4r
1oCpD9BxhVtznTf71na9XYqBNoXxMKzmxQP+1FMIl1zE0MK4w34h3yfdaA1p
X8sbmhY2gUt6M60jD6mNlBcfAgJYeG4voEkndWi0Qcbfbb+uDDc8qgDRtl8J
AZmzxg6M8yh2OlUyLgR2Hkc1tzl3nkev71+n9hcjX/IUIrFg1ALbkwwcjeXk
N+MdhBmDEP2fv85fqAdqxLLAE+ZehyEyXEYG1YLiKVNAFPtKhFHbP8JjwhMy
SPn5oQOXxckqaNGo9EGZk84T4GRtIPNB71pTAwxexR/zMpQrVZtwvGH7P1cc
HV9RdITSlUIRU4sqMVVU7sItfxO0EtPGfAq6FZffacD+SMeNLmDp32YkUaWG
UG+OFKO+heZCjwIfI+HZbjyXmANJZwIX2f0HZh6taiP3S1fCmVujDUFg23Ze
fa8xooka5LCO8HolWp8xW1m+eb73qxfRFOsvmlg7f2lhlRDubpN/jNR9RGnn
HXMwYIwqBwHBOUST7PZMV3RVnMMuj2UPucrj/gPNZEyFZ1TLbZaAwt/sEWZk
tKaZVx+CcBVQ7d2KMU1DvPYqXt4XRuSmXSkMYMjvfEDHPV5Npu3VfzTy28pr
SopI6CM5vHwoIkYP2J1X5oluqLdn62M6A0LE0cYpyxhlp1p9VtHyNbJQN2Od
TjSql68F16iYcOTjwUZOLGdwuQhOEY6+bkV9mXabU8uBuPob29psMPifTSPF
vKu+uNUj4EccLmS3eBQnl49fSYeFpH6QgD7z4FK9KYcUHpdSstQFFFdAyeby
4Dk7IoyeboXIWswIKEgxgmRQMxU7g44HtHAy27c4C9ffK1Gtr3hNSrlMKwly
q+LFOvap1Gy8mSF9194J2Pekh/IC8QiOybepPU9CJkqVAWpW+XmR2XvDtYI7
IPLFi1YOPLJhssZIrQXInllBsuZ5UBbuHHbN4mamI+JEN99aELoEx6Rr6rAT
rFm9o8+yRgiGp6cc/epWj1a86VNsBxhyB8FOVE8xGbtoPQdCvfMbw6boFWDl
sOONzhGPwoKCezP0lnewDFN6ZBN21NAidiHazePWD58Sv5mI5nWBsi6R9E4c
wjuMc6gjPFzMqFYFokiHyW3Ta2gPqvMiF/+w6a8PPBwAyKZV4R/BdSkMJO03
Mj0vqt2A95Er2xfmM/Hc3iwTteHEFwDyYu0wYyOFiEEdcLFssil5P21syerY
4rRoRVvNuCSQh8RmwKdmqH8RF8CsVrtlpT3C/b5DMATb+RSR1hrFpE+8H/Z8
7JLL6b7iDKVNNTRN4Yv4RlP74Aar9X1VXySn0LdfTEjLrG+4YFIPlc0x+rNH
4GWIGewAIgtjyrz0n3Q1qDnqDR+TAFasI295uaLRhwtYZxSACSqMOAI10ZML
YTnci5Pi4ysCD/fVinmtyKXUWuu2pTbJtNufwEOQCjjtig9hWdw2+rWxSY89
69qkt/MGye4HLsGxzRD4qjGoPEKg/+e60T4m+Ce2xbrbWbOYMSQMDNWnUVnm
KCnxyofgqI5qfCyDJcXwShpPXnhxA4KCL2IfsOij3W7DPZh0exB6Fr8hQcOS
C5+ybwmyMZ+TUUZ376hard+bdvUczl5gcpYSdb3gS+Be8SUUD/CjAiQnvqsg
hln0+qtiGRkB2Qt7FcziNMc548mZYZztZnG6qZVIgNGQAo7OBLFBWhqVokYc
G+a+ytNz00JMXRpb30co4y5MqcSzn6xE2IemMuYD2TCSG85jpWaeCTisZeuP
hTqxn5ivFCyl20N2HXiNpo3jSQNmxsoXJ1aUgvnHZfVRiHXxZ1K8R3d58Z5a
/bbFVH0FZSKm+s3iOYRzmPu0hrr8qbascFooPbYfH1uriiPzpwXwQeNtCjSK
OmUGwKEdBBXBIt12R5WTMknnNd/tspoIEr9GAGroK2LQmNGn8WGulmLjSUp0
nVqaJJEHc0cJ+PV5zMv4gI/5tbxJqHt8RoefbDNKW0P5+Z/RMQUvDbDrGWa5
138g3mcl/ui1EH3XR/jBcGqf00ezu+DktAaS9Ksxhj7FM/ldRTl2LWfjMdWX
T4RhRIpyOy5NT5eAtbZfZkgUIvjE7WAAafvltRx5HzSWAMytPsz9iAUOfzMI
Ie+p9Ligq6U/XcfdMz49JGusTV5eEiSqsDn4INgQhNiuMdZ7YAKkWDRI5x5Z
m3PUeN+oTsi9R1ekBaY/V6uYrM/Y8hZ85rhamE4JTdpRWGZ+UWHsIpGgJosf
6lF7SecuZlQ8U7Gc+BaFTF0HLADP8cN5cN0HTQ5tZFwr3GH/3nMbiJBkyWIP
kvY0IRq5OCFXoiQ6T0L7+RF3X5O+fy/LdzbTKvG5M6bHjkpqLIpn/SFzRRD1
kPMbU/3ibzil8xeweirV6D0M3DID3AV75Zav1wQv4Aw4pll8bPc/BS0ubsHZ
9/9pIkRRwcEJ76v59y/ZFD14rLuzysGZgiZAIh73cTNS/7HVIG6TCEKQ3qKS
K8Hu8mwHyTo7Qiqxd+zakEOIxIxpQJq5Tv5XV8LsKUKteztHv8AB5/+c2oVR
WEMsWfF2/oGL7H/hZoFX2FIMQkU845jpj1NR14mKzClXzrBmcOo2pmB2E1jV
sE3ESU4cVg8ZVSPKTaPoROtannHAwjXRNfHzSfbrwIi49dvLJK/oTHh2JiSr
BY8TXrYxq2Zy7u18V8VzBFcmE8rOY/lw0BV6+AcxaGdJAfif6M7tLtXPsYBF
BpfV/iE5TLRbOqsriajR17u97gd1YMajwEMCromQs4uJbSJtQYQHBSVcC5qO
Mm18slkogGHsg0QOBYMAWm7/b/RrlAeyiL7m4U/pcMpBmjCVp41j3846Tl80
bsvNdNksbvgkvd6gDT9e+aIfSJHFXOTLo017oEg77BPimRd2J48SxhkLRf3I
69Yu+Z5pQV0L1ySfBYlEmDjYHb4WJMENlu+IkYis8H1IWDKAecpsRce+BTwK
mXi5Ds6/XI0icAwRzYWrUC5X6g7anNScnmG7M8IRlIzLf9/22ObHIsnd2bZ1
XNOiIkt9v4euHHnDPZm7xlILzHlbAbAKI3JwZyljpkrzUITF5o2R4AKlaVGh
x22xivqiDHLWIgYAIzY6u9Q1EseoHBdi57t5gKPYnknGMn4+bLmdoPvdT8wV
636YfaHkLBRUiW/dPFotoZ7poSaZeXNaEKPkQn3gHUyA6+uepipvFNzXCWGf
V94WGbpHnm3knuro8vo+AeXbQs7iVzNyK9ToKhikQac0TXk2d5rVf+o0F68w
KZR339kmnkCjGvhgKd3PwezqT4Ti6dnpbLs177E0llL33rTVOWNdO1SUcnzz
PwWaq3XM7pS2MAx5jZ9SWrqq/Lrmnm53P20Vi9gHtHZKL4kyWcCJPU7CwqJM
FY3AM4nHrO8vMoKew4hCA+pPwGGetibQA+l2pOcTiIGpFvs8Zae3+sD4dLJL
uc0+y8Dslt/V7hkxOUkTckHooFCf8NKS/2qN9sLgVMif06kQSoFfx/0woTCk
P/cEliOkeD8klUt1OufkzAgTwykunZZ07fR0PQVvM9x/l94Uny0W8iAUyRH3
HfubSUcb68raqrsLJ6OCcf2lXlC/ScRf7VRz3/aH8+Av3+LqV3bIy9xUrAE8
elPmin7NhKssJ+JKA57EccBHV04PITRxhknS0Q570JO18SDxvtPgtkr/Mms8
DGMJ23Oo9UUxeE+muGuxaOcyr2LdKL9nyZtUAxvJHnD+6ScqTpNHwXXwGkzy
tfSa1rwlD36oiHq71n1cZGN3OG2JQYwVgIoRWsFxoMsIiAGhhsIqmtxeFMKu
xsHUOhzLhcTRJXRB9MbudCFAb3tZ+BDVEj1as6tlaGE1xUp1yZo3td63sTv9
Llrc0PjInd9GeJNc/7KF5ghFVWodH23DD37EtL57uyB9Pf0A1hipR2dUoF/w
H/GvFMfPn9zlcrwwTAmlD8XTcRfYirE5TRZhpKmEK4Hr2r43v0uiADPA2f4D
jLBXLHDWhTFhrJ+SWvEiRgDnhYOQgnNauu3eru2k5rwm1yZvlX2mGfe8bmqF
lvXTSgqbsFozPH+b+pHvR/PZyX6rhR22FHfbLrd3jNAjakvQ+ZwXcRuEF326
Wwx5QnwjC1WM2uGHWXy9yrxMyKn/Hhpo+45nt/wvB+f5Un1sJIYYVHZX9n5u
oxHZ1xD3QE4kG7BdLWkRWQ7fg28GjD2cxFtMzLiS7HGH1HP+gye3UHP/2c6q
X/uJ/302jl8Tmawm+s3D3m6wRM+SfBNQFxn0z4Pg9DLj9cvopdb91ALlLpPs
Jf9BptGx9TCoy1C7dXMp4rtw1HrqVXh2ddNG9ZWjjXd9o3aLWXVFmKfv+GRG
U9Tbt6LvYGiBoG68wqv2TgUTuGMhoYYJFWyWqs1pm9/xYVZPOym6xKpblVAe
p6I1KwBwB97wU5086MBZzpHAUgFUmINIPxCUIYhI0xMci7m9lhblF0d31/9a
0GxQeqHfvsyY5kmH1EvGA3SApDK0rmYjo2Knj8b5TeLfqOufNUyOwz17mUuD
ZIC2ijb4HPARLvEclt+7nYp91KpfNVuiAfSX97oQv9OlCO5bPRO5/juy5dY1
YnsrJ7L3mimACen9PqwROV9JmaNYPCSMePM118DlbOCbqPWnP2fzKIjhMsDi
nHGyH7RZxCgWS/qAJtiBZoFZty3ln+klLF5f0uda7saX4Y3fnLGiqCiv2LLQ
7fWcHZRZY3QbCYHBMBqszSRL7mM3TFeOeRZwCGoDxzyj0N3zCmxxeIqb4pCD
oXMiwIuoLaiHrFYj6mYwb7TCnWLa7vVtfQd111nH2L9NS/wU/n98FuCwB37B
TQRlXMsOnaMKM7dch+H9mN7OR9uITndC8jpjDD0rhKC5xh0NqNTpGeNN3J0j
sSot2cOyM2VFfVlHHlOlctbtQNRU+jPwRlwSvO+Jf8y12YSImWijcKNu9rR6
P1yfK2J9laSB3v/4xBoeUzyqJVYBwqEKzt3a0JFbbVFE2mxJY4dRteLqsahh
njT9ovex9xGBnygXwtqQZoh70iHHNwXpnx0Z9mpMkvz9pmwqY+mQOERlSYF3
9N95deOyNCEUmPS8an3qsBrjQYItO2N9I+jkO5XL/9zmRw3fMjvnCSa3WBIS
gcSojFhvCXYb+zye+Ygvvz9TT14p8bZmiVjan7aVUtMnjaFf7kqrtfBstqGB
t0kHpZ2VI0NguhaPdxz1euvXfXJbyozcNzYVQElgupH6a+YV5da4Rlsyfjn4
ohg4kxZxxTO7KUErcEOIVcuQN77RrYlcAsDg5PJhWGjYLj3E8eKOaXU7eLUE
k4skscc4QAF72U4zecY9DBGoRzVQbf9AJC6+20Qo/EbnhSXlEoGXkWWJWU5h
0b88dc9jWQV/vU+EXns9A4pqVdF/2Uzzukj3rwJXz//eZh2z0gBXyekr6W2P
KHw4vF1zlaGWql1645qk42M8O9PxnuoJfUYfK8qQKhUIRFdNXX3XQ6OF1dQ7
xde5oQLHukPxWrzDre+5tMvvXNVLYJ11aGxN7JICVerYKZxm4zQwznhTz7Z3
lF0+YZrYnbgssQGgbTjpAxDoHadb0kVvEtua1a0og0TMmLZzEQprRx55Pivx
6HIZC7VvlUE8Ci2fzNm9bL7g4D78l85cN0WvVHUsIsZvsj53VEMf9iw9+gau
7ZWjljuiTCuBXwAXgobEZr8AyzjYXrMYc38srPaPxIgixuc9+IWG83++1VOb
VXBRpHVkFZF32K/GXqfvNVp6w9uy3oIbXI+2lXr6h3bFLK7tN1zz9pBAiYur
ePQQfUCLDGNJRFz8rhWyPrOED1yz7/4yoGITiyaq67CVxb8qGREL7Cm+iTNd
ULZE4ProSyAWvVm2eNi8bsFEM+NoeLZ6sx8qy5umT9sh5TsrbIzqrGLx/yps
p+yJipVKR+vf+kyWNJXfPidt+QfqtoDpThEcWig2LWyOFfhwxPgUdVHGgUNW
kW7zaVikK/Ihu5HUeTA7lO+HrnDy9tG0kwj8ipyD16D2aXb1aDWomeKZy/8x
Z5njQsjzCQV/OACwn1X4IZXps/SWYs+ZezfbAp83B8f+Q4bKRiqORbztpAa4
c24h9c5C0rOy79YVpFQu+rIhit+4GovWxaJKYAfugk1+9L280HisesC+a43r
19/GO1KYeEg9KTwZiWvVZhfg/fWNi3T2Wy0GW1orcY4zileGh3VyEDU79m8N
Z60WXKGGq604pqrZpxVVFF5TkRZKOmj62Jy/+JbC4rhzy5HNFF6M2rFQThmP
ZMLk1fiSiIGVDQ/7pYFWQSGeTnv19OE05ajA4pO37hogtbijarFL+NpVMAa9
kvv3GgX/FJRE/6O2hOMCwIajShPDXRWAg99PoHl+0cEpswoLVIaBln6ZcvRE
8JAz0FvYwATJhMgAzWyL598PshZjXxKPsOBSdsmPLy/lAQygQyQQVRA6qEZb
yiNVn7slTeHW2AK9M7C7rkd25HZzsW7/4ymsT8AHsJPF/v8oON2LXdGppZA2
tfAalaKJMPiKOn2+/un7gTOtSoWc+KV1nGXh3tcvm5SCK/R5R+Y2786rk7oF
+Eue4jymoOJi5R7dCaOFgx3lG6OhtfsEg/vJ0HFuDdvSK/PX1ObzXXUz9b6r
C/JrIhdvPzAPRdpK4pGT5dhtHNKdotBZ75pn8yBhA8kFJfgAYeE+j7Kq/b2N
2Ocl49kiH7+rQBttSeGkM3pmdlfoo5VMSpg0hDQ60nxZXtpQYSeDovHFrfBy
kRn1ic1mgfnhAqCTphmZ5TZwiSQpfexox8Zqxf1k+B5dZURPcYrPimX8+QC1
1HLM69c0SUfdsoY/WeIlbGiP90pj0kMYcQn1z1vyuJ7QYnAjYMEduXgG1azA
YtQF769DHCxMpBDk+HUdDEyYEuEo0dg8qrXj4yNmoQXWCM36a5uAwWFCL6zX
eTxagNqQ5sSf3/xVGcnlFiW7ahWAEmsFuST0neuIeDcVrY+Xo6Q1iIj+fTsF
XAoUuC7Kya/UZB5LLssuzDcMTYfFIXhJ1AArzeGKx+gTTygUb3+KICvSxuj8
30PDJS5IEQHaEfIK/LjfYwlw1Kv0WR8M1j2A2l1Quq1u5XFq5Ds261C+dHKS
3VqzHaJiUQil2XO0FxEI1h2yziAs+33JglpO8CsUvthZt2EI4t41XY8d2xZl
bFlPR3agqsmfzLjlvjaVTlLrW0RoW7xjD6Am+UViK58LxJ1syay7kO+tJq35
Qc263+cxsBt/d/scYRAN4XKus126B4YrdGRktpyNGpP99Vt8Ua/cckEm3H9v
oWnOOO5HeboYnzLYWY4nf7Ln6ZHdr7kNiZIJw1znJqoHhz3JyuOK2xyoH+AG
wC2daqFcLVf/RWTsbfBny1ETYfnAVCib91J/BFWW4IVQBDXM7Ux1y7c9PM2U
b2hQIQLlYV7mzekzeJmEctdc/0IpTR/WrycMD5ir6/58YmFt6Vm0O3RtMTSo
xmQ+2GwoDrdcUAoQhYByXj7TIcOdt/0Api+s/Ngkx9I9n4vmnRbuyhWoJK6N
qZAUvR70dH178EJswQr6gL2Mlg+p3IuMKiLCX6D3+Bk1n6oq5ssbpjMjbk21
ugAqQ9m3e/7lGwmI4Ofd5drfuFrzcF5otZle8H7SpYoSaW++eQFy5Jps+6IA
25OSA/ao8rNst59snOguakWbQHX8OJgBCyGXyA3GKGl5UWkEdV1GSCvA5LVf
dlpYOoQoK9pYJdis2FDl6IAT1/GD6M9h2XHzjP6ONDWY1NHkyC4solDFMhSN
IfJX74MoZy2K6hrO7rRWvK11qD4jkXfShBhxd+L274s8II/DjAi/vPWGNB1T
CoYlgzwsin+868ByaRQqKWl5/ryxWuEzB8/2458KkCByzH27RXKsgYaLKAww
b5VcJAzHeUmoPgXGaQBBf8Togc5dR72k3vyhjq5D7MBnky5q/uBZzCKalact
bLWPRL1V8O+Isbxp9HfRaClGYJeXHXp8ANfpyyFyWW2uP+9pRPX1fRPXYYad
q1YUqoVxO/XBRjG1g1SFBo64lBO0JTwVj3QzLJJAsssZN0FMwl0Y+yWY+Aun
vMXWIlWHQvtxSC9MUlv/kBWfjSxdX8mxXwqu/KLG5CCv3qDBzEa3aGfFbdcY
5DxVIxan6xUGvGcKZzUSLEc6y+sPheAHjH3QiyWMuCJVLx9CXVGg92knsLUs
8Y3XIPo66tRMrhbD23ufgzQmotDFeRhGDSOyA5B540QwNzAOXLNnSGk9wvnF
z4SobZKSr7mEZ+i1ALLmYL8Rp+KumIAhq2OhjhlR3GjB+LmwFNKBW2dSgWok
wxhG2/JGIVC2HmOZ5MX6VRjabpC2izu9SGO0CnzErQwckEkhV2sj8YB1GGUZ
JvT4jNDzB3fBHLsnlt7TMFchbFSbU3iB6bb3BwoLKmcxWV9BQaZvWsQ4TnUn
cXF+zUBtQIGV7rrgxZtvbwvEJUAiuKa6gJTn3qloI0QRvs629i5T4bfq+8r0
lz6fjGLITMUP2Lgfjt4GmZoTG6RutPnH4S/XEEhg+a0vPMQYlEombt2sq1XS
z6rvZO61QAcuD7o9ZTshGJ6aBk8Evsp+Bqal9CEwY3jalzLYISPJXtHN/KrH
6NAHtRVphhKguSCzhSxiiyE7Nf4BuOBtQ+t+kHltSg4b3G0ycPJd16JIMQ9x
0H4WP57Gbr3zuwSUaks7KF4EVczo05LFHlj4EDAEkYconwGmU2gqVzfajxvC
YrAVKZp4zQe/vTq56YL2F5rNOgsWYqvTtXJ8c7YgONKoWEZgLtsvs/2ZUCv2
gUyAMy8hPXzEuZTruTe3vs03Hm3XODFG4ou1GgoKuBLCn1rJHotDY2zM40k5
5b8omCIUZF5Wi1cpdEsPbu0z1wsLHvqmg/w/XzgSzUN971oHUCUKL1EbX4Hq
DFkTO8DBNg6XRqGjsMSLrcKMZnY/VfKbPq9LMxEtNVTPfMzKApxVvHS3t/5q
pGdR2iz08q/Vpf1DXK20P8ktUZLajTHD0S8tGbFf4BQEcglJr/YX+XdapAsF
L5XGreJTO+gqbYdf4CIi8ITD+SjqNYhh9ZOx8/8f1jI9AGcUg1G3/us9n6e3
0q30hnFT8f1wh0ShLQ5Auk4q3NaCrEOv/r9cEJcPCwCLov6ihsWpCAL7VWxc
8DXtOlp3qBsLx48FiR95y1WzyoqpgCZbX3l0syuV9IBPHk3E1Gk66YFOUXp7
11p/9twtQsKh4abtytDT10ydD6XZcjIyNUZxhwX10g+wtdb16XUku6YJVuhM
thtSQmZksm2pJNi0PEKXRY2acOhRW0RwxhuyRP642QkoNXP9l31/Un8zLJ5X
K12k4ifefjOGMfli+vSg03oXIzs2lYIm8hTgub7OjaR0G07TcnO3et2p/cZM
tIdcIPLbGXddVt8pvm78DP9xSDieD7nC3BLnv+kpkkkzTeggm2wu1iCMAzb0
lRbRiZtmVd89SLy+bmy72H2uPeewl0LJM+KXsRmdaKIJMKTGwfzgc4mkEhmG
tJSb1MtcbZf9uNJgq2zGgpTC6EHM6p01OP2mb1stGeC7wdQS6hkr5Wni5I5e
EqjQZl5qV7d4teMIrhhWDsh5kduFQ60ZHHGbIN9HBPjPn3xVt8w1Sli0o57b
66rPZANRnCsrYGyaMjF4kB8Spn12h6vyMdKzNB6V3P6qnyep8jjJyBf0lw+x
joArRxZUaDTJsGCk84Rhs/3XVjCfm4A3ZmaAaHGHNtoe2EwZD346mPtc3oAz
utfEnsvbckSVHa18ACnw9dfT6TqNzmnOM6GEHD7AZyd1KCHCe8QTMxRDP/zy
Gjq1DiRTqVbu7V3Km3qLaAqkmjbaOLq6eMNdf47QswdpKP+Lhk+jvLRVNFzq
HWv/4TEaypgmIEu8YSTj9WBGpYrMR/obab7HcJFYVSJy6/q2nWKUW7yc1rWJ
l8DQ9/okHOGAdUhmhF5iITZd9lzkQQ0ofdjqoowp8QUpmbdChuwFiwhuqFVI
5Lu7CzmJWcJ1efX8LE3h8K+/OQ5qYQghXdGiryJGcq9rbpQUNp25cd8nqjGG
e9jbnSIElOoBdwPBhsqmRyYmT5cx8hEIMjEHOhzvPfEXacuzEtaQXr8M+Y+P
lsdX7XlJL74WWKEAr4Il7RbcbcppaOM+geKAKg63AaAdKNLONFA47urcWC/t
ovhu9lz668Ej5q3/60VXmQVLBEOQA3DqxZjCo5cfZmiz3+LBvF5HpWOYtwUz
tgqsujMlO+T/r0gFf+ebYNArc/zElEWgmZ8YlTT8IRGb10uO41+hZZHWTdCD
xNophWhYL5Ia+umjTfVDCQQ0T8pafVLPehuvsO6mgE5tZeE8ndjP0p1Id0Tl
jeMGc8RqcciSjzIP4WR5NW7T67e6ZzGJAYiP2E263lj2yuN7FgvE6FvLHilh
4chqJhnx/ocqzNVzCAzJaGYht/MG+C9+rvv1k8zydm+qE60/UQsYV/QV6P7J
Bq0NP2+WKW2Jop9rDtZsvF96f5wVMPecbnI2Gqh5clTGUqUoExev0DTeIAFv
k4ZYhtaeazi9QkTVU8utrrotJ7RRuFmJh+/GQ1YRuJRMLTezWW28yzIeiOkO
9aUSd0Zb2xwh5cUZpHPtRFlyZGIlFIiQ2BhofmSUTp6eh/0VaE7X2P5D4cin
fAxp89DQIvlVfHPGl0Yd8AqBm7iDcIKSWF4XIzGnqRyeEoB2GAOFeu9FQWoC
htuld4j0MLH+1GKLsirYIw5ek044/yKsuj3sUPwHjFrCZDgiMTjNHf/kyf7O
fm0lSQkh5I9x3l2iJIVoGVgtv78cVZQaqciI4OGS6iQ+mgLqeT3d0RpnIs07
EpszJE9tx06Ie5iHwOADqgchkyHlZKEnYrb+EwgpTFJ/DIqCVLM58zf9WAGz
QegSBOHPUHhpT2r8Iu/gpZ1aL04WNdAXSyBcvJc1Y/lxRLg7d4XGk5RqMaPD
fIOFuQOHX6kgubCbhKyq0tg0tFOuTLMAxFiCdPVRk6XRj9KhczO4DYH4Uxh8
PffNujX5GOOuiIG1y06CiqFLdKl4qdBt/8WgZjdTm/5xcw+wSyVuD/tOKFaF
7jvoujRKjXQXyErc87+TBP8AIqx69o74OX1YlCBogls5Qu8Q+0LFbM4a9+0O
R7rnv3wKJ+bbNiTROeKwtm/dDVso53kg6+v6VWxiJXTLEpmf2YJVq7Bxv235
Ppk5zKPJEdz1P8se69sCFS1Myou8vxjIZv+l3TCxwKQiZMmjBuaZpgnaKRK6
cgXW2xW+FwyFhtGzZVQP0eLv5WLpdWWeiTz2GM3zW7XUiFjRPfimSBbPiRQ6
n3+UTDlRL9+hSxyQuqJd2ulqvE3Z1OyOop458aVV1xK9rFEi9MZ608ZMafQF
TwJA6dah3QnNrkokoP6Qu5J3TtP07+NH1ENF1k1kzXP2vtm5qbAxtv1AYU+u
hotK0HIewnBwQAmgON+0jRI2fj+3fWGv8Zce1OxIwKsh/wr61eX0VuNrU3Gu
/CyImC5jyxiVRA9PkORb+AfuA0W/Wi4CDyrG8lEgMYjBKM2h28GbD5n2+ZWj
ik46MZe++aLwQbkgnzuyUPUrTE8VJDBWVKRihE8OoOlX5TvsVBCt3XrRSDOO
DRHznA0N4GYZ1qPBC1hoM+/80ZUbBdFEyiGBLdBI0ftr2DHPX8xZBWENDKRk
ACe3gFuF0aRFneG63ErP6PYWulvjnKDiNU2Lebbw1b/W2fgE3mECc8/j9+F0
5nYWtQU/dlaZj4fhCIfFEUHTgpz0eSeXvWsxczNVQqnr1jRrRCgd1KprL2uo
S6Dfcd9J6x1GqEh47681qpUAFbNjBOPnNZ/JKLWjfR8JfRRHunoJS5VVHKUX
ZMczY/8+WTDmiTSu7yoK3c6b856NI/+XR2pt59w9KTBk5O53dxtRH+3aXVOQ
f2cfhm53uTimccsTlns6RRoxBjBvRMvr/3Dv2UMmVUncEzZpBUPBiQKI6fn5
HlJFKj5efX+BngP+aKyDps+g5Dyk0h2oeMd3Ga5ZcOnUX0QBu/0YCIaafrMk
HlYQGjjAv6uGgH9YCC69RmdgeAubQG/7q9f7IGfmJ20aKHp6IukHrh5xR7IZ
0kIgW38gIyV7jZQZcxfbVV+IK10aGZ3o+ZagAAMImRuy84DLskJpa1VeIVfa
yQazdLlYjONE84Qtw+jcAglDGQcKvzyKsy6HDu6B3o+hWA4LJ7MlSXTl/u/c
Y4Qifj/0gWs3NEzgrb7FtZwsCyFCkALmTxtiB3Fhbq8KVyNYuLgR9ojTY+id
ZLzHvc6gkkNtazr8a7WD4G5c/GCqJ8JsvEeHP8PnI8DqcWfPg/HOZP7E3akW
LbJPpsJoHp7yA4rM2jRO1qxl39MQz+qm5LNAcJrBnQJaGS4UiSwShO4mlIEy
A+I9VPQ5VcpAy5r49V1nenSp19fcs0A7ozKo52bn+e3/2ZRGhQbP2Q1myWIZ
v3j94GGm1S6xC4cEMELCRPEtmW3JC+7sykgqfPBcd7nMu9N5UAUCngctIqnn
abBiKNQxBWCf+4p4uvhlBlyrgL+r0W8B+2/FrF8HKRocqqDiAWqutj7WWfJh
Pkl5VDhOeDkTdnkGrBJkS4zYTNQUK1ijtpfz5OWTLXWzV7zPxIGc5ipVM6fl
+xl/lfLQG0kKDNvatpEd7Uo88WM0IuRjwCBCI5rqE8/fM829XY0FKG1zNaHM
WaRfNMMI9WIyvgAsLHPWvQldYyhBKhC4Hr4oSNFtw9aTc8PPmDRMjBHPToBR
hDvFgpRkNqijHH/JADAxVz7JcxMGREbE2e/DJ13Kyv0zaR6YfcK+UIKwcfNH
6mcXX2IaKHW1tcvS3BuzeG3uo0Pk6/OGqokDjX1hc4N/XXmj93ba0GJOXrRi
XQa1LoCq1gf+fW4hq9PNqHGpqWdrC9sJOf4pHNLvdn2FRPPtrD27SyvAO/lh
LHai6KBXmEeHWRQ2tQ7Xw5XYBwzbflFrJswCMvcTNsRKce47TOCUUUtpK1fE
ydf+SA5AIXIfnBjBGNQQLmaX5RmGneN/YLfEXqcWx+0JcyJIJnVVY/IPYVUy
ekhGBtRG3fM80wEOrB101ZS23/PX4VHA8ln/O48gmSy7S5Y1m76AEjQauwZE
k+N9fsf/6+B4ONNw0IP8cILoGjoXIHyuzyj+nNHL7GoCFVH9odmBwDkxpBND
EcaiyT+Hj2fPCfrX9xQvjxVmRRBzoqDAy+izRznuiLO4nQB5hGJ0pTapxfHZ
y1rPvEBsS+pDXl4CEypls9naxhT3T66V+7xul9SlSoYGNiYSqxVEq1kX8B32
9W3SrCFUYfi65s6LHoe0sG7lY9AIX6y8JplOf1lhr2dVylJETu+zODAObSZJ
MHqBiKWAau+4AtwKlBNAFOURGy8ecDjOyb7LvZSucJNVoSV7jVUDUHYdGhzM
8e+oaB/GtnJOKQ3MVHjHFHRFOqBVRQkWne8kWYWMIIIVDHBCuUbf3YwTXydI
+gx3GAJXRDuyICrw/M4qUi9wXT+i+TwUue+r+5gVGIGQTlTIyZdlKXTocYSi
UON1XzopVtk8MQhMr4L6MjDE0DDlc0Lsk69YYnKvUMH6rZsPZTGs4KAaNPGw
xBI5ue803Dc+DnM+5kuR5fdiKyKMPBwH3GSgXsFY0cetvuMjQfjahqOxwrfG
rdnnb2swTbraNM1l+VSVJQpwQbaMBYz+Im5UGibaptc39eUxKaUZPINxYwdH
J9CiL7q2Bqk5g5Wv/6Z6NWIkRyLlED5kBFQ82gUfByAm7bV3ldsrQ2Zv6hze
4vqxmihPf0RPiy8K6NZ3Mn56923mvFv7uBvNTetFZ43BmPVtMcgtzfhSpNtI
WebfVtatKoq8gxBm2V64dgwhCSJjl1sOTh4XlWvOdE51wMMcVYVI0jFLfKKl
ZA98wyYqcStpLg1sNpxOC+CUydgamfqojPxGU6I9s5g2y5pY6kE1CGQgXrMk
RqI8pryNvGECQgtx31POO85paMjTkHoPE3KZxBu/6sJc3ENEFyX1xsnX0QbT
4b9jCpDxNIb7/eHdZDondnYGR4P/+NfQOzTvbVRWBTolJjd0c5jJ1jLw28/x
3GgUYVWx/x0Nsq/SBFPw6caOTb7cA9Nso3c7hErdFUWU47mCNsSl/R//U5q1
4ZTTZsbl0HbQSVp7Wsk5JrqLjrGPNGj/1r/yzIIQZCV7wjgB93Dw/LWP9We+
KjTENzaCHlZPN64am3RzIXoDXYSQHl0BaZUMJb7wYFAUC9RGtYIN1KYWCp9/
DB6zcf5IWKfmCiKz5gz9/XukzZVdCeF+sMzQzgFOJtskAdGcLzFoB7XYl2/m
/hChpAu5MMdjQPvsPOeagAChypY1aRG7Fp4LIZcknegXeLTuUB+djewA9Dev
YHZNqhj3sML5EzEHD1+S7IuWA1CXR5skEMHGoWeihNiheMdV/G6Wa10kShWh
4nrasNG4+YCLXKQhj0dut95FXyvacNf0TBG4NJYXrajCxLp7Lv8D42hdhsuu
zDI3FIvrPFIGzRrLMecuqrwR1JMXu4RnXb6KarEMtM8dfShYvH+YlPMYJ2CN
rScDDljoXhut00NZm1yz+xJ+R+sAfTQBU0k8F0l5YgEtJ2yxr4YHZtGC0XIi
7bYGl35UaAt9eBInGzRJ3R0c2WrgDuQmV0snflEBLImCnWFY4z57zx07mwQi
j2mc07SVxE7g3WXc7RAivjGvI4nej22xU+PSh443mi2XyaPgQQMG5fA89zMm
aPMjUjrJw67qgIGgG6iqJCbQPitW5n1IWWMyc6PRG+3UCVvXgX0mp1rTmjZx
MBytVP5uLg6VlA+dRORlVgIYz6wNMQ227Q1sUl5tpxhR7wAzYWx0fxiFxq5y
1tx+NwG2wrihWxEHKVZEeL+NcApPq2TVOStQkdUMYjnfZqcXCc0Z+Kx3AmpY
SgbVnQEHVmOiC6R7Wie+c9oVybq4fV70Dlkk8NsKKtTL3jzWHs+8SFP6uOUu
clCMauw/E5PqNpOWI1mZ4Czwtg5P+Qz6s3EzaokGw871fBepdJgwKD4Yu1VO
xUHN/4rvX3eDzMCJHCTBJO6JGAnU1Wm4HGXHEQiTCWQA3ujTYNpIlRUduvSZ
OTNi3QPShHPFDP3WjKCT2zL9Clyg1MX61f6fly15y4oaZiTXsBVL5XqZm1kS
tfX15w/bkRHA2afBTiQfxsIzhvEnOIF7sRKwaAxHTi0LpIBp3tYuEq+2P0+R
9Sw/To0jBppvaZngumOpnqOQ/cXTYecAEYXj1Y4bNrVkZb+9QQVBDoSMYzxq
oVxrnnNwCk316jKoZYPEh0WDKDYGSXbavIymNED4zc0M2Jf3srPB1eIYutTW
BOabmJ1U2l+pAqiA72+4a4y5RpC8pBX6Q+tVXFatWk5mRMN+TsspPX+OyR21
ew7swGO4Bsq3VHQcOegwsDOH+NBIukvNEXbVV+SvV53cK2cK4vOVg3Kaf9yT
r7/gbnAiJESsCYnazRiJnNZD05Zeu3lxAomkqjidD9Uo+HMA0JuuxRXGMRCD
ppqiLIQ/86Eh57eEy2OWiztZFhfLwCMhdlv9FNzLWgyj/w5Oqotq6j/19n0Z
vxywJEtXX1/z7kSpQu18wjaXOMfGmEAUKkAnIzm9kfW79qH2n+i2mdBt1C3j
dC6GqQtV6jX/+0oI7hQ5gHI4cxEPgS2OQA14iOWMb4GOTyGWkpvQpcpZagX4
EqILM+xBTXt3vVErOL3TZ7/ABLE+qiu9JhdSw7OCUiQjgouElXKbDadB9lRb
SytJ6HvwiNIvpKBKhf1dlzLfP2HGmf7M2cZUbAeHsauXeFLUv4qVYc2PiqUt
6H8BSsx+EzeD0n+ZK/y1Hgv5NGxLXHFhDOPASNYR7FVkBZod7ImNnPpKEByw
e/mLPijZHjajZBA/c1+oX2z+MBV4WyiApQaPs9Hu4/rnxbqFLdk/E23d9mFf
WtIuFS81U0EsOCrY9I24Y+5rTZ07IU7gwoq0kePZ2GI8dpAbfYEyzbWhJdg4
rlu8lvVI1Q==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+Er2+WD8PQYFVhZGqFXLU0wT+/qqtXrmuQhU6QHrIDT7Z8yylEcDYHAOVxQHm5rYtM5xNLryTPGmFlu2AnFfX7+oNWfilXNU4q597738nZnAoagoGYh0vWYGLicCYfGWWV6lECCRXMh2qxNlOzNns96fk8RrcqcowUVmpwDoZ6wFO1Pgtz/sHpaRwNvdK+tyD3EwagQY2SbDHfl+N8DzRloSkM919mz7c9aVGwLPHDbtHfgyK//SmJwABXf9xliFmts7wmoaT8+Ic4ibQiPkFeXoIkj5fg/SCn6mmJw1GtgHbbM1nd2wd5Ib9PNAPspK55T9gQJV5LMJxbJRmynxi61dFfGZ3N4FcGKoRCLU5nCCgpcIpKNORY1zzWSQcWyeSoZT0kswfuRYX+LPqofXkYhUHlgjK3pDCpzc26H4WoPaF3e9C6qY2XkMSDINcsrNvukKabtkvIkf4qOnievFy4cM3rGoeOlBi1NSrmeQJ3cJTxuk9BiQeFEWGYRhuU8TsdttkAKM6wd/lc0jGuHwIWrsOLulii0H88nnO++1/7cuBJAFHBpUXo6W1gJkyukC4ciiLNFqCiM3qnbHpd4tc84bTfCMHFkqxcZb6h3iWktPCzBppS1XmaI7Bw8zWHJcOlc7lgd01maSmnzZEU1MvRNwdpJ+jr8WKp1ouiYFPrnajSiKKJsg9tOJN/BeRmLwDt58d7keeudVufVWIGSUXvRF7DpW8RWXyOygRoCO0CIETKDMCDG23PD+WRk3t9euZrr8zpwqSh4HT2Je2P2Y931J"
`endif