// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VgaWNqbBpLxiF/80+yGxGY89T+7GD+6knWlDlH0UEn5jAk7MCmXKeQWdV0aH
BVgXiCpd9UrH5zadtznRiAmEa9A1Hh1sxz8xzDUtxXx46NL8ymSPJUDU2YEX
cgmOSYuvG7jL4I4bZfGXWOFVtD/vVGRVBhtUpWrXXnszX1EEULhUfiGwxr4t
q96xqE8YTCljYUrr/IhAiug89sc+SCVBO57rgHdmyTmYXnzG8CSN/g/TMEjC
pcZ4GxnOebxyhEMHCa3LbIud2W7U/LhxvKydgzbaivNOpLpUbC3gMymYuAJN
te485zZWtkzZX1JYGeTDiZ43tsJsuYzy9EZK9ZOqSA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IHVALsA7Q7pUz4Aea9wrgeIjsADUiNaTNj8+o/KECTojlNmeH0JaIgUrTBhW
F/bjUTUfFHzxmllGIhOxv7kl1m3nmhNnWBtsDmON3f+ahsDzmbgxAn6fIrKv
RDkGOLkDYk+jCv1MhPiVpDTXCqzFxNVrx7owgNgoIR44ikR636Oe3MRrCBK+
x4CgpKcEF5mTjoY0lrpPIhNZ4MgZTVcUkvNxTSA/9NJ5Jz1xGs4xNP0SmFAF
g94GS911BdFSyT+2ocr6ntw3ZFRZBHSyDGwA7bPRl3dOF1/4OfDOVhovyRa8
zp5KFFAqGIiitSXPM5C8Hk6RHtg6YgATBsuYL3NE6A==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QdyFdRIvHyGYBtogeVxg7qEBfFeeIT53CBTYKbCMETCu3PeATTEjuBmMe5xN
E7rulfA0g9MZQ0/M385pT8ooWYLcnTg0eGVueLLylA80WJa0yOf38lOfh78Q
CtBLrq5WrM3W/k6BNWtIaVaYxBd+l9sphtk7h9cKG1hiWRD2i3zw9BnMY2uA
LWM+S912xNYql/r7reTwwJucEtJ7IccWEIak0MbmaP6elpKhSX+YKHRS5H8s
gWftd8DUU1Yd+7gWodrQKstR2mEYznyC/jDW+7nBDjE/a4CD3xrj+klr/VVp
alXqrlkhC0LGnLdvonIFiFSKmZLYJjqyJ4pTmoJS3A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
L8H77mAUH7s89xmBcGYbKO28RkUJ/yVPzHs9SOe2V69r35yT9tdRByM5Xs57
QASrXzabEbzUn6WkC+uFzUyythIJsNf6Y7ZMSRprQCH0QRzfiK4Qr7BUbk1d
N76A4NwV8DAjL4GOh8PRLzn1F/M/s4kvfM7g9AqcPiKkvLHkVJUyLnpnbpzk
0loJXoUmopBki2jFEZMrO6CL4jriYhVohnnIChUz/zI2YTXHv92KysRlv94h
ISIUNxSwi8PAMRK7wKjSA2qQI+n7BSnJ2bO7RNLfNY2QHUVBJ2sKhZ4sUMjW
+6Vc6HrWFrfc+JaiX5O6Ir2IGtgKVj4/l3mqihTNOA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EJEuqGyVCzVSitcUYR3iu9gnpjkttS3mwQz8bhZVawulUM2xeOSbC/gvWWoc
w3t0omJOWrOo/93RL14UGVkOn7Xd8pinwQ44hjt0zb7eq2/B7NN/zVf8RqTK
1I2BNcVfwO2yFYk3Zuw7TWV4mJzgdrK1dO1a26cbc6ChfauRBmo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
VV6LSLg/aOevTzMj1hlFKnFhQQQCG4WMRZJ2mCgyEGZbMepcjVIjP4g+TnZ5
YFoCnjlEsnOYQrNvAp7s1zZb/ZvrHvnjLCGh188HIWSKJQGkEqSzuPEZHVpP
12KNDl+zmnmIK+MFvTrych7qWIcE5bl1JBXFNACrL//8+2kLTSjABRlsRLq1
3po30le6LvhqT0TMik478dB27uMEoCgLT3dPE0h1ggy6xXSm9qrHTaRY3g2z
bLnVtnZJIrXZIkT09p93hayVifJGgB3sWqqdSN8ixXjK7rIHswpK9/YsfRTc
K79tQ104WSdB8iWIEhXFeLR+FqrvNv/x2Nilu2oV/GuJr9zmnjNF6bBqHUoX
27gEc+l41D/Wk4B5NXhySFoK38a/bbtTHa7fIUTAjc8qb2y0g82sealuBRQs
diWZSelSqis/qZLrsfdddVuyiJ7AAVQrmS/wYc0bSjDnlkZ08ZgwbaEto5/R
lfdCGHKQIabG3iGBr6girsORh9/xwB63


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ab/tf7xBLwtWFnfdRAI7ApACBKnU1k/XnO8XKnMXedxgpHlbACqt7yKtuN+W
LtUgQuVaO2EYR1a9HnHGY6VjF5SmcHUMuUz4ejyKlVykUq7zpBRGnLJgfEGV
ADt1u/s5ZdxUCrIuMUJnR1W716CdfFhO4ZJleR5fzTZUbhOypF4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JLG4lwQXeJ9F+nY3okeDZyOKzoGUkhlc3YVdEKhshAVF6gfpotDI4a3ZdXrG
epcz6iAJ5hkdVybwnRXwUeaYkwJALoXExoph5S1YSu0vNN5wKLc66qMFUws7
VlUpsfeJAF6IolUodcNPy/4+eUubgHv/qhtM1zmrwp2So50BPiE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3120)
`pragma protect data_block
XOL5klfAPT0oyElL7XvJWOQOZZ4AgOQd2NhUa6w4Uctl2L71eePP/zUV+Ud0
PcZIdLmTaB0ki/n41wWJ3WTomyHKs2rgTRuKLPXiiCPQg3B1JsaWDCC54vcO
nCAbJGfZ+LAUpZgx79GnokfUu+DcgwYDD3BP/DNvB+L1AqsERraeXdkdTRRW
hWRbMYxeDfLzm0ss7sEjUWN8jzKkbYVSlVqPtAgC717qhdvuO+KAlNQGvvdY
ojlFEKKBy072FDkq88Bg+UHfTFXOom29T1xsuqJRxoYzW1fEY5V2xla+WQpJ
GY+f+pE3Rcc9QQ0fFOZe+RyClqtcZepSsPKCXh9+P8chrKZlZNHmsglkUliH
sftc25pL//btfsz8ENl6jVAaxpfyI1rDL98g4H+xMmc7fKyla8whLp8K7RvE
VI78gXee0IniohNXqAt4pCIl21OK860GjSsFewozwaYkG/tD++1XiSlcozSt
JXPkJjLa8YzLeL3rSseTEiQP/q4ej4YSgJ4dnaQOwCjLTKjCCDc6MJBsuw/q
tG89XF41AcqUNwbSgyRAAAZ9OQ8ikZ5XBK9BPUkvRP2ky20rH8i9fp4lh1L/
68a8Wml/izVjmbe4mJFlKnn3Fx6KNhq2nz8ZBbx9DbP7+b7UeEd5v82AYJbq
1W2GZ+R3GiFyh7brWlS2UfbRKK1KMzLQGrVEwOOqaMP5PeWlIy5tUo3TJiZn
nh3vAeA8mU2a+tPL24M/iyGU6XeNFY0PxaP1jomyZ99roishUSet3f/MJOlp
lEwSzFByhxJOZqcC3cb01AMTOd7gEUJyDMSDBX7E99BAR4+7SQA41+G9RkhB
5bgpUoe2ZrAcBNfsO6rvWNJb/d61JJ1SxkniXT+Ev/cYmzioRijE8WiES2GB
zX54JulQDzL0UWVhmQJ3CKKJ87wCFLLr1FpP6T26SfA4+4GLKyX963QWoT/8
z/gzo5oQEFdqKOGzUrTFwDkqr0cGh9d+0qpVwc0w4rcOZWZVRQARsgTbLr1x
NMCCNV5FkGFkdz9sMsLk+IBkHneWE2mfYBlfaEPYDFeVx0ZfoHqvD8442ikA
Si2YIyh3HS2QNslMsXdi93EkP4+t6Y4J1kh2x+X9tJcsqeD8GVljD9YGNCIY
fv8BIgKiSAGBKuZ//Fb12RboKaO+aco4Q5uy4W8ZpLdtEdqP+5SJI6xwqS1f
FnX2Ok8cp58wnDIIhCI65mWf0f2jBS8XQO5OPSXvqcs0Ue7uq1yqVVqeEz17
8a/SusJgSjVYhwKMtLmb8VvKhfE5Dh1pp7OvheQ++05gWI+886ZPWQOIipPr
TrqSxTwsR7TLxZRNF4G4uF1eWuSclkNJFKQbwdpAhsslMu5knMz4NNP7bZ8L
HHdL/vM5/Y2fZ9/W0ceCWzNtTJlHGUu3ZPwcJomJrjoMXpCDhbydTGUAewDK
udOMU8gaWkbVXN5tC/iEMY/uYCaDaYlOe9KxvlET/hrKxyRmAd4rr+3/BrHs
xiv47ju2tL/lROUri9+bXtf/Soc1lEnARO9ihbfrsKd5ZxmRs2rd+Hcdt/cS
YQ0clLsi1mv0nejmxAbCIFVCyvAZQ8hj0CtPGWUjGZcJjpaEdbxPMQS4GGuU
CaAml3iLOmsjkJVJ8+nL8gI3bin/wPohtiHB6iQTdV6ma4ewIXxtI5oLCL9H
GOpvxmGtF3kwmjZwhLT4eVrkDQtVQW7jZfJJ8/I5co5IS3MQDTyHGXim0iRo
wnwH14Qvq1qnX5b+mRhJumFf3pD+P+ojXhmbWeYdXiPcLsJwwVcbYYSgFe8i
ge5lWuolmkBSTKNARrw4D0mIcwvoLq3HS4rikmED8wH6MmRA3zFZF5jKi1fM
LTUT1YCG5WP60uMsw3CXrGE9ogYe4dcHqMP1N6PPqhydaLXDwLG08fA65JTO
RUEnAmA1TycwmSNQz8QyMmh6jWD7ymDfcQdvCy+OSKokf8wLX54jXqSe6Hk1
4sBss3zeVSRh67gIpbJpOswvEsNxl7L2XhIVHamlw1G9rhoBW2bR+23pd/PN
XvZpFqx4FUNy1jwBFxjxjv2EN/nY3BHPYpVNP9tXznqTN+FF/mGPje300E4e
W6wR82lT/VDLpg9Rpyol5FAiM9waHx0/NKKXEREPAVqln8nMr/byXi3CHB3h
O8bZtBWSkg4DL+hkDZQfu9Emor+tTi3s/ipP4wEawp9uYem86y5PnDbVvqm0
+OBkRXwrC1f47bWdw1h3/uc5wFtypP8t01CKMLth5duM0S//I6ixMpQiEVGZ
g/Xdqbq4rGXUdskJ7sXghLLjP0L0kqn6y2cnu3oQlcgfcTKkZcg1s4WCzS5P
/V2lh0QDoJrid0tkCjt4QKtO9hwF61eCFlrWRfcTIsoCSRxPQbbffr2bNEdn
ZmDULLycbOdCfPuVv9RMBKb4xgN5rbLmop7YKHV7axZfLkazyTYmdEtsTcgW
sm4LkRnI1/jY3ARtDTTq+tGddW40KAuwn9s9gp7IOBt8tYGtU88ejNS1HLH8
Rru/TmKVg/sciBhLPM/DaA1XxBs6dtQx+WIMiVLTabxpYHZ7yo1skGgTTVmj
rOFvBKmMFdHFivDz5kdkuNKiV72OwIM+tMmGW8nYZg7t1KMOJ8r0aI2z3jej
Z35XUxPXEdd80gb5YFhWsGgnizCF1pnEZBivWDgqTgpVoLW5fcaj+n4yXIxn
7S8rAIUNFBA07uLP+aBugMaIxxxYbuhtAvbMe1hTnvp+kEzTtEy4F8ipHQIU
KUCyRDULGYvQRngrqMLQZCTijztXApWQN4ZG0BzAH9vrxXT3csSw6JmqLUvK
PCfLHw2A342AwawZAxbQtbboYtxyekZRH2cWy25mPksUBj4WBma2T64EWVAZ
phBihmhvB6XHxBxGSnevjcRuAuQtyBuemYsl5hNg3l+bhfpGSckNBiNYJbWt
HobsHUfXio0XV/U4692mtWnAo8/hWuJ8vqdjAM9dhd33Ip1Du3xvWb5dn22M
tPPX1BUnzppVqawoonpyqKxY+/QutToM859ODMr7cOsC5B/LYWI8fsRjWg7E
J/bWBlbCkpKaRjRL2Ed2GgSEQgsdlkcU5sqPLF3AUypO76j+CcfNLiC8TCbP
gOwo1wNc8Ms35PX7fKwMDVvq5UAfmRPHNJCkJbdQUKmJmOer7mIHex6XIK+N
YXoSKkPiwmsQcYj+5bBfI5SIPbwal2R/RnZyAjcSoffIRiaxhrR51tNnqWtO
LdDwutPExIgax+29ZvutEE02XuzYChaZrw5gpwNp50fC81QwCeoQCbfZ8+B3
i2ycQLUkHpyg1a1J+GzM+Y1UbSXAkHSx4/lhsWKubm4THLF6oxhLFu7VpYab
Z7WJuEFA1YJLJOnFyMNzH2QUbUrmD/rJhzVLJ9c2VgrE1Fy19bdg4jltBTAN
Q0iqbzBhK67dZGXEpqZ3r6YfG4IcPRTtMo8rzA2FWzWC4TtoFzdUpeamZ6RG
mFoVCdpMP3Esygy3MKBYOsYPVqYGJ9r/k5JiIi8gx0BZBztHj6X2CIfl+Nsr
lDmiTqf0/EXQeddcZoZE4msw0L3fYYJOY7Yzv3P+pF1TDAZm7RIPQchh1wNW
d6xtnaP4Ahzc++H4MXhcu2q3DkYqp/g9hk3B99M2e6v5OwceEPCr49zyRPoe
00d2PxuFx+Mc1BKbEvqaOngq0YB/4QBImIO5LBdQV5NuBxG209SFIYudoQ9C
atdWIvQdXfmh758NkWRVvNMtD1d3nX2NqIG7kdnwqiQDH6Fr/jgq8h+T+six
dC+eE+yp9mi8SbmuV+28KXPWpCFd3FPe8x+FXD0TVNpX/OyROqSlbtoUHQKK
eoVOHXThneiAEOGH+yRgQ9h5/Yf7o/zXzMD1oQ3enInzVDIs3+18+MHq3w11
3YCsB68y/fTiqB8qC6qtcXLnWXN3j0rlbpY7M4QbdKC6yTJP62IObIn8IkuE
Y0wq0/udYLdEFZhnsFv+IUfeLCYSE210eBY3Fq97jf7YI3FX77YUOlbdfEyv
U0cJlrle/38lCcCj+wm/lh/NTZ02ulcPbW5VL2kg0aXsbT+6bOz517iBdl6a
nPRv98V74uit5M1Ngn+bycEAjdPZKMvU+k9Aq7Xc9SxO+bCCM/S/a44ZK2H8
OBJ/HvaMdjZf+RWFA/up

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "9RW93T28GeolckbYRvHffOsKFRFmORm+azyCUYhudrVC3P73ufaBfyRVMCXUVPfCA/gVx4qupGWo2/MTXHrbiqujt9kp6+gvryDIvlW8esKlSeDbKqIxzhLY+DL5yFAjg+mCmTKnMSoiZ9J0N0zgOO806IAkac+OYN9FbEIEFuaO+G41krhhxrcYAZ7qVX+m993ig0jH+TdTkf+bgk6VV++svRquWf4VNDUj099hz6BAKTOqBA7vkTSgs5YY4GuMHU0yBGnZuTgeez7cNg68tWvia3Oxc0qUc4aQ0V8EjmeEREiqQSl/2AGsY6++rRSjtL+zZQ6u6xZEB17l+V2xOkLaNuW0/uw3C7Zjmzu0sPb/4p09m/5fjlxabBrn0+VKTITt7jaAoYhatmk07/XMky0+kQ6PH7MvujDi3l9H8vsykWT5gXO+4SOcUstEnDMW+AqmPmNtW2buK1rUrXNI3jrPCwCXAMOV4mWMzgYQkHfIOvnEy7ZB2CMQ7bA5IZO5PZbR06Bqrje8WZyQZ7kBgtnImPa1hskKygDDGlKUEuRSkkawnu2C1R5w1NyVEV+b84dc4h1pnvNrRkNzshOarmIn+aVurHYXH3O7zK6erSOPmBlQmnyRlHIfAcf7XI6rXGmLl5j+gd44iEQEqglHyXX23bT5VKmGBOw3Mm8gnO2egtVsydxZoAYHMAYp8AsjP6Bx+o6YDXIELw9Xp0xfJOpdnwy7kZ0LDlGFfR8Yc20cF/7u3/kQEV1RtlyLqOgIbwkF+jsfmGufagOVx1aJL2IbNJnzfrjVq6a6tDzYcsQeb5RXWlDrsPCakRY6P6t6IQ+ONSYNXBR/gue5KvMIk8PrCp1T8U5W0UNSLRaBxgxIODeh3Y5M/W3RXdCL4TXkHXUNdxisB6BDVraGvnTx6mGZZOnYR5tG7qXk/ZcuveddeGnznMcCPkA1XDmOTiVt6/NqSMNI20yOAhz8hdo1cx6dP0op9SdeN4hRxc8GeJ4Y9i+fEcBpBOdsQRsXDzK1"
`endif