// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gKDjgCB6QUd3n0cvRt+qkGoRK2+cHcWAq+uop11vfxJc86XH8eFaqpPjiOat
A+EcrCWcSU5OmdOwYoW0QI/oJPORsqMwK+Pf9CnBlq3dXk2vToFRSar/Lfgg
WAAH5Pto7GfKyokndrCeY2RaannWbe1tvyGuDABKVt8vuorp0LsSQpZQCtEX
74VOVVAOuxyX5jwHryA+crbmQr36WDO6vNM1L8t5JBC+gXE0azIbd6mfWiTR
j6Cc7jhnn6EZcvMFtfwkyerK/+QXFNYK6K82H89yFroqa0XhZrKHivTO9JY5
7VEOXE+UaLqWGPotJYhBmVexNpUyjm/eh1GSOumnmA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
E5cR5p9t8uKNCztLHcsHiRYGAHWLy389TBMSDch4SZFiQek11NuOU6IuZbg0
RyuskCdmUil/4V0SJfQwfSdxp2nQC100WgmIKGJlD038HVUZHTqIJ4PBZZBG
HLtVO4Sk0ULtGjp19IMBrrHjgJWMyXOxIWylbpnBy6Xa5iHEL435+Tat2cli
IhsTzYYCzutU02j1RS2LVI6YeNRKRrolMu/E1jyVna2bnL3m0r71MeEzADnI
+RPumwIw0R8ohK8OUGOAjYaurzihyh2f4msFljTCiUxhOtT2YP4LIDkjzvId
y2FK3PO7YVXhIn+SJnjVBqXweils1U12IVPTjRxN3A==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WsVoD298gWjzG1H7puAREl6+ep7n+wU5Gy30BvFSHDXJLbyGjm1d4XDhldOP
j/hg/q9nsDm/xy3euqTjth89neK6LRq7lyuw/cZmSf0keodTdoUkwmVT6E7X
diuxJKKUB+PKnvayseuXP+IGV8qwjq7mceQD3E+HE7SoteCF3SSrH0zDqamK
RQdQCfDqrHfR2avXlfN0x4geNC+Z4OeCt9o99IzD+ExkiRE0J1smfp3g3dzE
f4KJYvBhLyXvuGeJZ+iWyyhpNGateubyoM87EmU538BA7fR71IrOFShbp7xe
l8zEINB/feENxW9qEUhwqz6Rz+whHlLGifvIA2YcWQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CqU5KzCKxDJrcJKdDGVxvEnPH3DT8BHAuDh4b4YKZEDcDrrkzfDPG2M5MqaZ
pJ2ipDytOw9sqgz1Q3RO4UVg4QFQc12XJiOnMOQrWGoOnq1f3o3cT0xgKSb5
DnsqHxdSw+qCfApjrmJwkabJ5fFKCrCR55QxZcmTQrNgxL8i37KiS6PgKyJ7
ZZOPMZHnWdo/JYPa2fbjhKkcXi7C0KxDvNAISahXewLF4H0FoT45qvqM5F6J
rjmjlg/lG3MtmpFGJH1GzQzNCBFOhWDdXTv/dCWpDuFLiMN5bFtffLzmKCnn
/gu/5KtXXle/Bs4cdQ5dB41Hs2RYjzCHpQNRv+hKIg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tF9HuXe50+3bCk57DQ3a+zwPN59NwMDHIucidZ8I1QZDsQiYHAyZYg/sIWcK
yd8IlOxVxcJbcvEiRZPMW3VCAP14BP4zgfdIirtFphPu7UnUXU2lWaBNfLz5
rbPieW4BmWUfsRjfJlHl45/CGQtpN4WpK5GGJUU5kr7gEWe10oY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
JtP/1LEfrd5CgfmaKw/xKqNQB/9UTRQeRm3b6AgU5lIvnqwAQsO29pTFQPjm
bb/c9gOfi4KsyApRjTfSBVvF5TDQlsgCb4wfxEL6QYmDIUij94Ar3RpeL9Vz
v59uagDhyvBEvSuGexBrcS9O7RAD+UM629LuTvUbzBnvNle6J9HkMnCp8nnI
mUGgurJalW5Xrpk4G6nnshBO0vCXP7x0dXZ35o6q1BzZaPZmjvSAwWYQuNt+
9awiT32ahOT/C49dXdrwq8vqqljS3HJu9zUGqFDMxyVDE2zMsKIRf8lSEXJ/
YoctVutHPHbeTfXtTTEd2W6l3txLOua4I2hAmFFXaELdEq9yi5WhSCkoC65G
x8rfXdyz9zllBKIZ0mxwbxvu7DtEzQLn4bidF5wHo5FzAa8MhBJvtc4RWKZx
314Ipyb7qVxerKaV6YvVlfm4ggPx9xEnZ+A7ucWNAHKov9cfU1xud1efAe1e
sK/1KupYpa3GSeU4BMdlFXmUyhwTKjfD


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dEaYgn2evj7wNydm/COSLQCtFhCizE5YWRkb/vcOyEJU1a+7zt35skWIG60j
Wucc0E6cvzW5jNoGFeowayrywF6wYBFHLq8zEq7ZgYaQJp77V87hSNHzbgEw
OP9uvKCsBJ5JPPC5AyuCeJTdnlhFe0zgU4tVfWcmBcIeldeBo4U=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rsEsDuS+eLTlOGpG95Ovoi5jhmNODDn7K6HX44qFzFUnU7NBKBD1wyhzWtL+
I39wybqGmbRwxwGWPUJX5AqHJFp++5uVOmG+WL0Jzbz9C1M2L+dSfvbmln6w
ILCbo5w1g7/VoRxe2e+iIAQ+zbCHiVrX+VveLjMhmFVq77YpFGk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1280)
`pragma protect data_block
bIs3VY0fpvgIGbuMTTB7jdSF3wTL+DMrozDUWPGOYP1e0aXXGvd2Ak7V8EmX
NdgVDFSmcWjIGTvbumtNId1X/YT2GMjELibzgaz9CZ6nle+YTOi5yBHmVpcV
v454uOgoEHCs/jJuyuPh3jZI7LH4/ryk/qYwTByYXgmjO1x+Opb0k/XJUllj
IG471yGj3NYaG+iPSE1y91I2NsRUL5puMr7n0k0bryoWvM3oqu722KM1MuPA
tV+//kKUIiiK2c8Km9HQrrZyro9EL9x4IzY5KhtU7f/QfLvSmP6hX24e7+iZ
OdY56rgrsLUcl/9BJZWjpI3rJgCz8PaBVD6XctkxlcGKALSVxtQYujd1hHMk
LclEJ09JKcXLnpcUmPUQAk1ZjNe0PvSRzOWMTojOXEusXwoXp9FamBZ8TE0j
RkPTqLrIb/Yj+FpjfKUsAsPK28rfHg34/qfE6F8gWm0010EXUZWA2WewzHG1
qM3BRcHscNEmm5KEnrp6x1RxJoVfvosyqwMi16eg9cqiD+lhYtg2ry/j9CyI
wX41xlssLKCWbujioaxQQHOG+H6/+tUaWR1y+83ESPUXkggc5Fv4DyRyn0mW
kmF5Po0lVqWsLYtg+gk06fklBJe1jBMk6xEJ3s1AQm7btrTc4g7gWQs3rcNx
UC3rE2muTXDni5aX9UU5X53wwSHXhp5Au2M3UHYGbmhovl3BncZV8U/BX4FK
M6Ce6Cvz7iCN9mwfOLFvt9iQNkl4AZ3FXezMhWjJQzyF57pG+ksRGMV5dhFG
u08ae9/Ni0xtD8l4pI9Pb34f5nWQN1rtnCr/8saTvuhCSNbJIj1O4HQ0PERJ
XcCj5akKZN6ZDI5YJqpGvuLgr24jO0xj1RdRq5LlOqJ0d2E+QtIwyfzQcEGS
YQ7MbFveP9p3Nt+x2CdUOsO7nhSBnb5zLCwhTYXjC4CKAMylZNkNm09dfZKy
n8H6Oa+BeMbTBMuevGl1CO+mDyvgs4+qP/C3ilUfW1cYTV7oAewFRW8G0WfM
l91/AJ69W5d6Bt5j8FeGCVFkf32zfDq1WIGjyQex8m863h23vLKxGumJbGFX
pNr45hxrir3ZqFd0uBKGTec/VYQXQBQOty0i9eHwfGei3mzDRp+X7Mqo/Lr0
CREqYNr+B1pOFH9ki+k+VkaAteWTUnnDKbeY/1Dmseww4UE4PLEEKkZ6RrV/
t55AA3YzauixkC0gMaxQvOXRWoHT6r/naOOT9fYjlE1kFg9QuEe841ZmQa5B
rsB+e+ZnNGBM0ve9VRxRtU6kG5zTwdHdRVrwxe3+Doq18zJByhY9e3nwzDqm
tlhhsAvHTbx8vycmwzSK+DwDOA29maPutJwaRPeLafC5hxA8zifTEPGkK9SV
bKhh7+DSxWfNAU8B1aVNlxuIfyFwsPsbQZpvkJY+Sf8l6LvfP+D6kGBl44pL
DQHbNQRgWZM64zEYSvaZXFBIyv2EPX090F1A+9mZn+6q5XMrleYZZbwmPzVH
4rYscNlC7kXkViaPT1l19aJlPAPgj7qEnnZYvQ8xJ93R8vztmSJp3AID2IOe
eNgWq4HhmyNluUg9HtdK2IhFY0qmBaBxLUlbAlUXu/VzINLuWEqAV0v3VgKt
L3zgKhtTtrWtNlG8wKlKnSqbWHc6cZ7oZHbvfIwLa3/B2tHmbeWPjR7R8SfR
mezIb8nPc6UBdU56tCpD2g/sggg=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqdZnmGrP1KWfB4fXiSO+0EEdYkvKatVW91AwqgkagY1YXCMR5B7IWWCBcRHNNjsQxUF8J1ccfGRlDHcFiuxi9bXurzU6yNfCzBjlV6jsJc6u7v/5m3UtHRfjWRngSjtnTlT7+uYN8MB0bcMindDyPcl8D3svBzGK/aFVv4orf9yDVPTp+pHmk7z3IHmRo8z8mn3gDLpgxlDsr1R2kU0RhnrFyDIMqjeMX2WiQXFTJ7Yui5ew2OamktxtUXHHAjRnILXQeiSuHRohUluq28ZnokYMfmoAtBcA2sium6SQzqHUO8HR+ELG4eoiMSEXejZUZSOT8lJIJQcRMzIIhVFVPBYaDMV22CLv64OJBb2cLtn48caclhNUCLgybQ9+PMPT3dJV316lVLeRVF3Ea1vPHzsbeKwgN6xyAFjVdJS9hwfr5X4xMboYQG56drzC8ve4zcF3cjJ/AvsP7OEITypORv1vylPYLZCQ1omwxMEvTiV+L2rvZF3kgZ965xyQxI6G1v0M+sS2l2JX8JVhdbIwxYSIwog8vWTi+qO3fwR7f6tvMEAPmwqsQms+HVW/8jERkbhh2DY3eayVCW5MXo3hZ0MeYVyPUaLQQ9hUTy16c3wp374swtoOwOCTk1VoRL4pTwhnzXjtymTmdAbNsE07tRBFubwA6b4ipEzctzylrcdUXQbd1k+jcTmSRZjhXohJPK11nF+3hh8bwYWxiBPI1enTNfDbGOeFdtqTJMBicBpHK4lnG5ukNVOq+eFo5tpFuH5v9Q5EQzu+cdFhSRbEnTX"
`endif