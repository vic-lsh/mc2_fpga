// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Yo/9Q9hp+0D33OyvhV0tqArpdwGzkzmnZfue/px2KGCWh9kzLlpRBFGUcI6E
5wB5p58cYwial415E9OInec35aV+OkgCPcYTC2H6GvL8VuvWU6BIylPX4bRh
EjlCHxI0+eLLhfzB7WryteXiZWKDSAlogTwpvMni2q1VAIvNLnSzLUO4p4hS
kagWRQWUOb073ctjRI2WbGDVu2zwysF2s6qf8ZvyLQr2Fchk+QBSlQQwAZHW
6X5RknaRE528542K95ycRYaWP6iL3hW0s83E6tYxJ14b8fK+T9BS5CY/9CCn
i2N4NMXEI5kX9jXNs+Vjk9bFS7icH+2iE/gq+Eq1UQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UQoVxaire6jrSPNM3AR2dXH9YVUxUxpNb13cKba94q4+ABa5F/CmuY0bFoJh
SxHLQX2OFKgnF6RCJFFTbuIrJ+Zd7b92kYDltOfLIknQLBzGeaAsWCPPkb6U
JL+12lTjs/exvtKiQFxNmu0/Xe/lHd3RU9gaFmiJ6x3RJ2i+RVsYYS8o9ajA
VCQxEPLB2wc9Tdv7oZuHLaTQKG+/r27nQ2YdjsmBIGn+xeSE6DwtXsw+dtv5
/mA7JH/cHCH9o57nVBW8sgAxE5vWLSNMCke5+6JrdRRBNmwCXiAZxr4IbIbW
FZlnUVMTO/8wkS1or5GRwhrTkupBQFNJSP+r1j222A==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cXY7SgHNwlZuUhi4Hfmi67etdBqgHcovAthLIWE0RmFtKq4CNW6F3HNyLkZj
/gEu3zgYMwMVc5ZMrR0KVGSK/XEqDjlOj8h25XiWlhLQpn9qNukzRmaI9Gx0
u6FENGGCMF/q65/zCGW3cRQgoBJXys5gamv88ceT+o8ZuWmW875X1s39xdPi
jKZfdE1G/5sZ2XW4QD0Z6KCBJeH3H/9+ZDPHvvyi5JySRSDHVWVvkArnCDzT
L+EjKAjfFyuCc/wn/EzK7TQfURx+rMlQMj0LxD+NjIrFNSiasjoJdzDWm3fX
5TyIS4kQMge0JsegE8UDbzyo7UG/UeVho/L0iTa9eA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bXTau24+LLi1gQtUjZH/SZ+twFDKecqDf42b4uqdUDe+PWV7JKTLSedtJ+kr
48OKyZ1FPiL3fevyRP9qjEk4+BiHn/SRsjrPseJuiCFFJk2kQ7xYYP5lBCTG
HFNMbYCwN6xrew8uENtL+5FNhjf+9VBRUXGyXvSVMCGowQFwe7T6efKPwAbv
LvA4PWWuppukzWUmSba+JnB5llwcSDqCzMk3ny1EFzkFPy504rajdHiRDwSm
ri4HWDa9jWxLTTQzLPYQcK4QSHKm16cL5SKi7nNiaYCWgnOErHAGCkb9eX46
BqZ1i/aWM4xACo2hLXn2+Esko+8yAWrq362c4VsVJQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XcYrkboOai1yaHXgCUxVX/v1tevrk2erbfrgUXjuI0LIe+hkJvkF1iYQsonb
iA8Si5dI0/to2o0/2vyGml3u28JdXw9fWrGUHatDW4AyWvxFksJCMFO0e6+n
UeS5hstAll+PCa6WeHGSyKyf/WLehxg95ZeaR1eBQSh4N0Ydedc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
vGJCoPGrrxnJswj5l5DQKeGBUI/I/MeNZTxgNClx7nFiLvRmHgL+y6xAdewH
Fk2qFXX/YrnpOFMDKS/jNowej3bQ6Hno95Qv6h475Cd0zU/x3Y4Er4WptGJi
OWcI95rEBhBBK1tA0lCh9vBFNxBVTtueBPmlLoSz253H7t0/oudD+/oF9avV
IC/Jek/iQHaG+Bo4K+XkGIYNDxG0HzHjVCWYVauu/RlYw6LH9YHB9Ec9Jq4y
naUIUOqAZ6tw0CkfH11ENsxjIlQicYqopvAaeN5kVqUWSVPEjz2cAqZmnyzs
lPsUKZax0wueRkBeotaMpQfbqI3VZ28SiCBHEYI6/xzecgjD0um6i8UwFBHE
G4wkGZhT6NGOHxPYHNTbBxtDyQ/FfEoGv3cKETx7Qq7068L5ayI5DBOfb5v5
+91Yd7tti1N6orG+nBl6S/3Z+2AUB33eanZtGmZcXeNh/dUWmdCUWtSHjSps
EbHcASwNUFF+vHzXYGjEqiyxDcovVt2V


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
g33Fj6ZsdJuF0pAE+fw2UtopMkFXmlGOTd8Ws4BPlwTb9SA5wKEMYJLLpPrF
4veLMJhpBZgfNl7MFbJCy+4PfCKzHRPzCOlh//idLDxd8YxVHMSvRh3f7hYT
j3pPZKhyVXTd1znRXUq7gDh1dQAvixlL6LTiC3EQf81x1/t7mxw=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NqulsFlT3v8Tt/lzSb3J/1PHAG/Qqh+GE61StUL3zOYa96dageGVlOpW8iLZ
QTNx3tsKm81Gzluh5OxrOYcriaFxufA2OkwJP98DdGJ7Q12CfBDj0XJrei76
QjPfOjeF4eoUqZJiNxzkLbTyam1S0G8PVshKUw/a6zmb/wKZvPI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 104832)
`pragma protect data_block
9E9QpUg5RZEUAX/VuoA2Nq4BIwUGkkebDn6Ff3+YxpESCC/xpxdAVExMT2SH
1PxvC79RvZxdHIXUtWtd2JKyJ6h1k2sjiu/uN2jwZRd3/tz5Bfct3o8r0YZ8
0yK003UkdwnBLiKCMJVe7zB0IU31z5Q5HIOJxTDvSyIuLik6SIwFkx1U83qj
F1pWa06IICIjwEWolnelHs9OcTW2hS3TUgJCdz2/UmHK6tQs6zXz5HOptL7s
Mo2bwM/8/ZZS6LpSKVK/5G4rVS8602/REsAxNyNRiRuDJkDkJrV0sAxQF/Ib
G2PFG2SCuhmSBpgTZoK1gpTP7pS1cq7IDV2MB/4PZbOA05CgKq5N9A6YeQLw
mbMQRpbHJLg38SS0ogGKZ03BQMn2qiQoU3OMmBOhq3b13PK9W15vuv/S8fNx
tKuYDC0e+xb+drJZ3rNMTZP+o2h3HIsMDEn9VTTKhO+/KZDOu3n8+LpWAQNn
atbQVyWKSNKjGD+tsrNxy9JuR0G3XGmdt2qdsTiNiwnfXdHsa4g0L4Qomrjy
yLkzmW7U+hXBH+w4r9REs1RQAUkQwGgJ34k2FGA8RQjXvVDLZINn/+6OszRQ
JLOe3F9BbpHirEeMXC64It/BL5cbPg9TB+qeTpNBlQXmn7hem67iCtfVUlun
yHMp3sF/dL7cyra9FLaj8dbC1d+rGE3uRnyc4PUyFyl5BRyCiJ418+lIzqv2
nLZyicvV/1NWwZ0FZg9YsTZn5+TVR+0HPJzNUK5xUPedaqQ/Fvn/DU8XV9dh
yDByRsZhp25Oha7+E4PACm2hZXMSI3a4KggJDVI44kvudDujJLqABND6YcL6
TMlRyNhLtz8PkCOTCXykRMZLNAOJuXXdd+eW1gL0t6H+ynVPH/knz26RNSKr
tCpGPflqb5g6psD9xQNmjHUEuryxn9GuXSmPP/QcbVrejo3JZrIjp6udNSw2
267BHjc8Efg69In0LUnGgQUQXG4qWSTWifz5t0eeRrwoEDPYnJJFC8RaNvYD
/PploIE4GVhno4Iaq1yjRwiv7fRJAQy8gFYrUzXEMsP3QeSpNISbaLEEEX8+
8i3ewolzUZVATaLtwuQtWS2dzYKc3GCeNSHEJypiqmeVjsiQKZllG4XzQn68
UxaeNPRY65raz2W0a/dtqM5xw9DsM/qY277BFy+EUX5dhZDfQw3B5fKCYXWl
2j7++MdBx35nv08q7fE8H6cSgW26662T2/fMGoRUJBILapOC43l//1LvEhRv
Z0uPfRv1IbC28S502yXdGD+QrvWzJD8IohsywbhZTgwHr9aF2hXuPWM00CrW
YhRrEKGh01Bg/FEF9IHQ1RXIGGD/iTof9t4nqipViWPguSxy1NYx80tQO2PO
08/MhzSrOkPVJfRSiwT2/ceo1u6saIpBAbQIBvThFmqAZUqglXaffktkwoFD
0sPc7U2LomS1bcbOZdvCMFqdxSSg6PLcFgoAd13Cx6q56ti5BLPPgNpI3Uz7
Fo3VHTL8AZPQpzvgeDp0rtDbhwL+KLHQJhP0ibi7884as60UuDXFgG1dNYPR
ywDWY5u7kYV4nIsUBoUYFdQnIesCqcpmm1Yvih0Mef/XCToe334+6+TZvg+I
G+plxXA8h7UDJ/IyYHYHxcnIi6DMTJ7So6YDeKTk65XMS5T5jR5Hyl0X05co
5IXKFnmcXob/GiMC9lkAnmKGCVd4gRYreIL9ksASnzBFlsob8XFERhMgYd8Z
GczfRA79pc4S5EvwzWKDeqWCDFbF0CJQ8BLgOdSHYtevaI/55KU2gT0QTD+Y
5IIK35qF0XQN1JLuj9jgTpSESd6WaIz/FZYkOBcWhbeFk/mhOPnGtTT2M9Ou
5dXClKSfZP+3oFWlFbUTvFMQ3C3URru5h8xjgkyxKM9BHK7FEXKtIBzNxyDi
ak8FQ+Q11HEV4cDFVa1wQIIX0XogmEWGdIWtr6OniSTcPPUVgNQygtQt8JIA
vJvGRKNqi2d/WJMFVZ1wRRbkNQuTx53ZPPNLBvxlbr5w5YiDq28hYmbrhown
atExwrKOoafytmmWLDk0XIc50xl3Nk0Rkt1Faq/wtrjz7TuR2cblplg0rE6X
lBAKaFuPK3NPODUyNaLQElrwnji0TNXzlAAaZJZDbzlAEbRU1C22woqdm0h3
28Y/c16PhnG3jOtiIcYqAE8fsgOUvPxu9SB7ZCvjYZ9BvXNT9ljzknLO/m3H
8bJzrDVUTgGeGERnF1ZXNy+kiCvCW3K9J9rsBdxU5b/BHlRfRfNs8cAFpX7Q
QQiVBWAeqXV0IxlSF4fcv94BRcqq/U9gbi0+whekq0zgfGGxfuoQLpVZjqqh
uRdMj+CTjVMq9bmDXBO0zGpk0plif9tmG+q06pxTjcEJ7i13FLHixiEGO1ax
rOjCxO7p0IVfoBFCklqR7+DUKpvkHCVsiuK0lvccQstAaS51i6coZa4SXI7f
sLtECbfVzk6zS5Psl4k037zNbroA6sEggXYZLejUaPOVcBE/bl+kfkrO6pDX
t95rLFzJTcchLpI9/afrueIug+51nWJ15OfYrrtzKQHufMEpnznjXKS8BSBh
lQnavMGR3YrbOVvVpnAbwMTNjGXUlkCWFGQEo6NAJfn8Dlpo4sh+qdFXfzQ3
E6TO1mYRCi9ZPxCfm0ZjXb2IPXWLu71WMC1utl67Z/k+W/9tlCsFTDNdjMhl
S7WIoUfANlu8e5iHQ+aIhjaehpXVL0VhMQun5sfTrX8qWqp21eFGKWniKq0k
h3oH7EIy82QhaYJ8heOEoC1lJDGhoIH9DmwefthRY52KvNfo+3eTtGYNprCT
JqUN0FcS3D2Xu45OcPv+ZqgLNsiSoTqDuiYYVg6n4FyZvFkpRUgvX+5DWqpp
7PWH5fV0kvjikap8TyU1znMm4IHOCxzZiGYW/Dz/OWaOL9yFYN3gWYiCe2Oy
PlJRLLC7J4vho++dZDgaFsbNcL4gmI9uks+doZX9xrcZUfU7LQyzxJIxtves
AGOEYR2qxhpErlFDWFevfXdOQzbobWspdaNCMm/VDK7H7bOcDlpfZjLdINMm
l9dUWhgH8ILRzahLKUeuuGwkLjKnmAKvbnOYKYai2bZN+S13Hma6Khtlr6U6
sDKDcqAUrd1N7iay9EiuQl3gJgvuM+s9KiTBckrBA+soxcJ+7uVqKedhgw2t
dgeSCvBjeddz9ysvYUl75LwM846LZGdsuZ2K7LOK0i0gNexEYnEJw25g1LwB
gvkRSXPR2oxmLTmO8wH+EudgfiN5bwQVaobF8hE68xjDT5iEkb1puLj2nnhU
/H/9r9YP56esdzvR/NGnx7fjcrPzMVv71Pvh8XbBrDFNZnQhHBAjTzwM5zFf
5vg0nmKnkfewURzmc+MBhqQydoxC+63bZIbnspKaWoCNQxysHHD8pjZ+M/Kw
O+5GsC97BAKgf0CnevXrbfJiF1ukhHquiYbaMcWxDxMWTUf+y9U8Mp7UQ0+1
REPhTYukxJKEfqmXff7WHvCAik/30Xoh8V4w4gzQB/iVo/69G0QcKQgt9kOW
FX35sBVA+OD3qb/ZRY8U2DPcZOEJPtqa4KMWkDZ1vycajaP4cvlQEEwBoQet
sVozE8rvCsgUSISsg01Nxq4MkdWS5FyPbwCRjhOX0icf3MJ3s6ivdRRARB1O
tp0OFxJxskcw55bJTFI9HSKvSqUMG5xM3ptb/lGBNoblFNKIgtjBJtsBGZ9m
muiz8jGdsrJPefdFcFGtXLNIuSEy30mT+R5FvEpHX9WSM6xICVFrCK44vE3E
7BgXoJAw/1USkQhXBLrYQjSJmhC7TGl6whM16rwibWGYj/8pTTJHimsVGdqc
3/0dFqPY2PqfJIwNzzSvDHfTeAogElW/RKVBqS2WHtpcOeyWe+se7Zu/iA3w
3sNSswXyiaC/wFr7AHY7AS5V68jlVzIqT0xB4+l/56zF2B5FQQmN+bxEaKy/
pMiQikc0u8GaCivOmCErm2TZy3LCkXfufqA2DeSkm16tESIxdZNLjf/i9jgL
IjMBwcmM4tUP7efuMCOp4zMqEaxpHPMCI1lkIQrtbqw6wnQZBF6mERTxDAGD
KOtyRLUfC2lV9VWbzFC19I/EYSLmrz9adfod0wJI4hVyUJcWuwL6n5ky3Dsg
vRInde5EdKbCAzp6mV7m2mXm6RQk4+dXralriTpBqb0yrcc3JBGpVFDf0D6O
ESdNo5QgI0Ii+Bvayh3kyyJunHN/qDgJgpLSldq6s2SvPT6oHO6KB2Dziece
o/37BfvHqW3I9QBPPWhoi0j3GzR6Yhm1A7KhV6WeYSUnW0i2JBRfJNBzMCto
Cx9oFfkcaEnS712SHccj81NCMb7MVPVeK8tteSrrcuvzM2jh2FrHzRv+pp+p
DdzfC6t3IBAQju71SiYL34XDY3FrQU4ZXiSBWJ7VlDf1bp5d4Ae5i4eBK43L
/7G9TZF3gokLE60/iHRz/laorFmQ1AGvVKiLM1z1KJiRVek1W2B7lWinoyrI
qWS3lgKMkTOCg3zzVzDLoxdMqjYFPNzyHhzTqjujYGCoUSd1wMcXg4gjEfZi
kpNFhQZjSba0VBuahSw6ymcz7/c7EBg7Hneq+ZiDdJAi7ZKhY2JM8TLNiqw9
YgwsgOZWwvO2VPzYLxyl1C/s3B2HbPEkLmIT0ZwQLP5yGlzoQTlOb5HOZQGm
gLc6U55oLmC7IGInvhYu/mlch01m3pNiEp2zD6eiutBEc7BJthYNNp10zapo
jdMEKq8tHtpaAL3E19QCX6CwE+r4jigWNtaiRFmbD/UDsUJlvYfkN8WHLoEC
ClOxvBJNTMWCMJtMH/rPNVydbe0nZKF9Lfe+L35GY3QSj3Ukj49YsapDQfFl
F5l5APh2KVCqf16Bu37jbzU1USxwEnbww17azdcbCsBLowtnaICWmJitrk+Z
V1xRhBEuubBZefSeIpxw760AhdgsHTQ+uOexk0gJ3vJPF4B+ua9Y23iwx80R
DQL4af4tqAw8hqJHxUSVPEr+1sdBbn8iMMM4HwvTw2d15zUY6mK5JcvYS6rH
MmjQz8d9RQKI6eooh7duYzEAdKdMjraWla0TqnzSCzoe9yQ56iP+hubytCwd
6wx49zopux2kbBXzA5ZCpoQr5DMXwLLOp90H7NSf8oPRgHi8w48MFOqvb8Ds
bGrhGrHVpX891y0a2Nzc/uvEnVUEzWT7Mpf/XmwiIg+v/LASHm2s4Q17FSkx
GIgCOTliLvcVi6U9XtzMT76BSaktXXwqRRf0btLnWZcr2n0vpDTsnJ08JZmf
pJo7SGtH1nZtFd6Ah2LeOBWKVJeNj6MlKHQd0UFXOMAY05z2R8Tn0MUuh2gb
Md1Kubl3fcpCj6I74oKINCaumB5xTylD/7Fu+VMMHdXvBRpp9V+0HXRdksYp
HWz7XhJwudjWNkM36hGdrfav/wwkM4vNpgJtQdOL027aVcbEq/aKAzOOVksq
dnGS9aD0Fjqo09AFuif8VTfSTG2hTkNWTE937x4cRge/A0yqk7pRO/iT4KxK
rDiOF2+S+HQbtCsicqoQI3OMluatNLqbmJeAcwCYSCwd271XbN1ViHUIAIRk
lLkkYpszMJMKsqhx+WlLaqV+8rHoKb4DV3kvdxGe9YFKwwE3srqHvzxKDlCd
CgA9pioObjgPs+s4Li05NYGoRDVs7wJ7QKr7Zx0r5S6sFQkCmbNuzRtz/N1i
uoXMibTUpSNAdxS66XObYpFzefL+PSeiAqGGHWAjuerDfuKcs8oTSHqac4qd
3bOeYoyINI5XvSeg1NuL85JIqJ/KpAPZiYljwbmqRjSWIrCA3Jl1jkcFrrkG
097KDV/Rdf2IrORHfmbgvsfzfHZAyS8mUOn3gXMqthmtmvX+sFd2G9fc7WPy
VQO/LFJkH3YJ6kPXPmz/56d6mqWeIr6HfSIfeGdytb15LiBwbl7+cZSLN+oj
GmGwOKdSicqjKCkf3ZVRESNQfNo3r00PfEXZZWFVZDhRo7D5/S9HXx5QFh96
FhYObxQCma2CAy0Ou1JgSIDy7yMjS9icUWtandUeAJRjd069V9Hkny6vK3kl
YRG6RFCACdlHVtlzjdLItyr9Tf1LHeolKKPA4aOPbkuxt/7hSGzOYlB3KKd1
EVQJkWsiN7p0i4hpoz3eeARMJRrIVn3pqRcvnfZFLzdzmJaoNfil8+bBE0d4
uJF4EnxxcBgW5l1hQyodwx3zsztH/zWrMDsLjnJkgvKawM6R7AR52rlRHsCu
0ieQd9nmMSeYX29a9otNMTlxfopK0FdhiQE/h7cErTvwcNCU95zAhoe1v7Qv
VjtxvHMcZ6Jl5x0YTkPjNg0fK+9kXO8Dvb1nreK6ru+dFO/rt1QtSG5j1gb/
A6fGJITdSZuqwnVZs8lKDkZIS0zeeZr4/1eE7153w/QCM7uh1Ib8QiIu/hT6
dhXIrSHC/Mz1hsZNFJdAM66lg/ozo8YNNg0S2U41gZVsC8g0joZFdFDY5UXs
z98/J4YCH+X2YAmfeDPAEK3p8C90G0Z4FaUsELM2JRmqs387g0YZU8g5A3R0
Vo/EXzZULHatwUYb4c58R45EpGFjue0D3vWgacSdsum/aPItG+6w3GpBjYtI
AHuFoCD35lhHW8EaYkO2b4MNCj2xXBM6PHKke49yt6s4ZoE7xxQRvRQFQ5mg
6afkBatnWJq5ajTM36Xw97WrJ6lE3fLFV/PfyhbmN0Kp8kTlgnalDGEHALws
bv6t0f+TLD6Uw3lR8rGqTGxJIN3tcfSh685XbL+DT9QUSW+u2cWRwXYOv7+h
cCxQoc0/ValyDkcbZ/XLNEDjp70HO93L/VgVyRVq6w7bzjv0iJMyHdLIQYQ5
+pKDn2JKSImr5TIZwxdUtOTR+RgCTrQNTK4jdvQwN/SQVu/bbHv46OPo0Z+e
MJGJAsMt45k65lxMFFDMb2TJduTc/4U3SgdYiIFzgyfkQacyNi/MUSUe3bvx
pi5oQG/4EG0d8RU3Ahdj6VuvOmkML0aZvrXs9ot3j1CmaR7owhiebSfLOx7/
b7j/kGPJo39ec6oOwrrCwKhcqqfOVTle+LdATl7whLTNUMet7wcqnt0KPrfA
oKelkylKeCL0gI8/TAAx2WKP2ySrYVfNKtLY/iXU3Wey54f1F7e2xEa/QYVp
hpuHum1wFNJ1PKX8QoSGW/LAlWlqhFx4bNggzA4yP3YW2KAHesbT6QEjL2YQ
CdBbnOZzYhnWwFCcEu9rYjkZUpxMSI+1w35QpTXreG3/t+dRQQFyoT2DZ3gA
TjwpM3hCi2QMuObO3rSpk9ZmFfPg/AA7U70WmdUW5H/qAdFdr8eCtZraolJ5
7EVneTCQiYtKnQCJOUOdpTG/UnUmj+XUcYxBXtx7nHx09/zyrbtr81kyrTSP
Bu2MOLOOy6hBmqmPdShqm9+QlOp9CB8a30esEMjdYHLoaJQiBnXO59kEQuaQ
SDIEOxYiU0aERAIYzdn5SXZidurlrozcG9DM9MIDDisvb9cjOzi5o5Beiwzn
SrwIcj650yuVQJdd0deA5Bdadkpu/OyU4h+05XvyX2Rm2U+uFSU9+HamWc/X
HrZlZWp/7nOHMFJzHJzbPicTpodnxgoQfKy5FlJjI3kjuGGrKdOT3s52NIcE
+BFiEWYMojk1KTr90kbihg//DTxR+KmFqNxFzIdX2KL7oqF0U4tHe0uQiO8h
YEL7i77V6kpsDU8zhgi6cplKKvMwdtrykWmHpq2BJXVvwerLUzwJgL6zsaex
owzL73WTxaHLHlEmMPF0Blr0R/3gQVk9exgGdUCG95OG21Fyz3jzlV3xv3pD
K0ovaMEPA5p878DL6QplviIOk8WBsl9G2nwA1vqu69IzsYuixeMYjoU4YWh9
kmnjyrbM3uBh3gD1Xu3vnmzT3/XXdSGRUWzuwEpngC5nyvxgVCeQ5VJ6Zk5f
8j+2w3Zd5M5q8pdXXIuH16ExUre6yNdEYo+hb4TN4pXcCUpTTNAD1zMckJJ2
7VLHXzCZKxhz0H/HfogdY4tnEpjzxzPOi7i67Rb6FE0zzyLU6j9mjwAR4npz
uEvgQlVX/LrbgtpbB9/QHS2t/ImtmnCdCsM9IXMjUwFTc6kh1fqexN8Tuan5
H3IQcmu+hHTZLIKkfsEaqYppyLY2c1dh8WRZdi58wqaf0T1f79C/kdEWzxfF
c8J2jYE0ru7UcIAb5pmLqskerX7PBDx5vhB3E3rQFMIzPL4cggyg6aGPFxQe
xcMw+22owUE6IWnwa3RBm+d73rZazj7aCGoeNJRr69A7260wfzN/PvFtSkRY
LYGbzwC6+YpxkN/iZ5wYa4rk2hMxjZzhs4H/DfxI5fF5FlCEU6gELEbSC3Ix
X9k1xsm4vdy1hgG77ODx6oQwOlvhVWLOobw1lVh0zU3jyRJBk+YiFVfHmTzV
Xa9lJB00uq+stk4jxFlUgZ07ncmsTQ9YyVjGTWwubQt9zDUfibe2CpkDSd5g
HEGiXVv1M4e0aYBL/Z+n6ox66H0ukelEnAS/IezqsscJWin9267l29qgjgdg
Q8TY6zvbu9Td/9tMSADDcdWCStxd/af+sxEIvBhdo1AHhke4W9EveKryHSpX
Ii6a8chBPmmn57JpVRjGUMI3jilRAFub2r3bwOy/Kpcbzlbyv02eUPDO07j6
/Ua5DEI3AVWy56E1WP7rxaOyCxwzYbZuyAhewP2TCiRoP6a9XlROVZCnWn7H
HL41QWvSOetz189iZW1h1tMZxmyfbKeOrafBSzsgcYxMZf+0b318VWUgXzSg
3RMGS1tw4yZamMIbEBF06wbmUNQprCEHJuIpSX2sA1ujXqmX8Ws38PwLavIp
F6uRz8YHUGsv5z1UwZIstbP54HSRWXXAj3zwtdL7aWf0aZKunQmeojiKEH7+
9X80IhhSDX1JmBEuH81eCX52Rs9XgluH8tlfK3RNbHDGQariyGl4kUCr9jsU
tn+amWHflXKSoijCDyn+yXPeMITbI5WqceJOwBhHASme82Y2A9T42boijfp3
725Tg9X8+B/i6UqmQ8VcVR/iYVj7dC2pH7e6UV2eivktgIc6LTpwBYrNU5s8
TVBzXNUJReuYeGFsImqYS2QivrNnBfG0dSiqYeTF03sJnMU6GAMXQlgOc73z
a2YoJpRzLT1xMBvqnzcXLscip+4O3lzdKD8rJPPjStvMnOR1UTg+iFMcrPz2
LiLNlDQWdlL6hVqW34+RJrIeovISxlbZvHcbSCm2bjy8NU2gpTyHE9FTWvzX
Q/vtQpDi+d7hKG79RnakByaspV+upcb+WQ75NRsVHCwj5u7LLYmM8BpFNTiy
hgrB7t/F3niq9uwWYS7tKksICAa1JWpSi9fUtXZdHxwQ1SrXoz1o2lx7yjgy
4JdnQ4t0R1UHrszgGfL17mIFU+/WHsVSFcRAnrfc/4daI3CJhbR7Fv3oekkH
A1WJ9DnCjn/iUx2cvmfxvse/oSIAUwlripEIb/gTQbMspXmOxYipAVAc79w/
DgdatFtl2GSaBK9MWU0UojpOL5pgtztRCEb4CaZcvagcTt2RF/ed32dijGn9
qvVyDnlZAx7sYC+98CsjI35cBLC725HnlgWvZ1ovcJd2a+IcDY/d19YeHbZ0
cytqUmU/eDRSk2OfR1UcGPAhJPWpo0vxpIu9WDOcUFLVuxXKpoai0HRdyflJ
ACP4yHp59UhzMpxPoE+v1J6ZQ2svBkrx/iqmwoX1Xk4I1zW5hu4HSoFo1ij7
f7nUycWU/7Tss1QPwQQu1Ppz2QER0rf6hX58+JQXfH4Cm6jk3aPSlWa5JXm0
qzt/0sRHtYRu9FkEO3EDaP3yy3VPBB1PrQneb003xwwtp9MWE72UXPUGiT5L
dhyYnqiG/Jgv6+qDicY1DciCXlF0jBooFpt+WCW+dmdV3PF6DqFcLrH3zyeR
ultIc1z7E9OJ6LJxXmhojOL1PfLb3CbicYcTMtfa1IcUtPt3ejE24rcXO4uo
IIeHZfA71mErY3m2bNGk7oxDKeeOvRq086ukqWsqG55RMT4hc5DWCZeEzAfs
qrTx92Bq+OuOBeg8kG79tBdKK9K6krGsaz0xOXCsmuwXepkZvxGaWfwKnlGN
4qE/qEDAyIysFlY3A60/7NyHr/cAhyQZoQdK5BugJwYqWLMGF66X8AOdMOLo
1uZJUXUaAQjQlgYxyrzfwtPsHtjCiVbLxMYF8akE95q2C9+bSPvIKkWIFO34
/nkLj2Z/ALcw/I//lzJsctRFeEmwRINjVNtootpoXxg7RlQRd6gE34HOJJsf
sKj20ssTTElbLpRqf7uOXKa35vDnZ8jriN/JCEp6G8emrlUs8MV/4uVN7Zfq
hmDiGdrZTFbjsKoPBtpgfQLONU2VB2Z2Hv0DEJq0nT651buWBhM5DFU+vZ7/
2Nn4Z/hyJQyBgRnMcTcRBi5Qe1Oe97IGPyiNv6oJlyiLmQGu1bNbbQVFB/xQ
5ZhEqHPLTDuVFVL365b1WbPZtbDO62aFuiJQ3/e6OwBvkpJGk7o3AHpVEpTU
cNSfyTqtvyB2wzDNukkAEXc6weJ1+B5610oPYLrwHknL6KdhGDeied3YlOV2
84yt+sqyY8yQ4SWAR7bk9CTETpL2rUO6sBJxR3RIlvSR2Etdz2PrQ3/C1uvn
MFVz6zn4VLCEFK5pLj83WkjGKHaWcgPbUArhYEgcsvsTGM7MdtPYHnUkQb/O
z07VWoDc1OW6Xjv0kcEVplnKuCujaxN2MmIiFgkHaJDiWHHoTY1vhUUcWomp
QmPPKRAu8+4bvKDEymXvmV/HCyVz6fhqeVVonzqjBb6Da1fmmfamkxRYboHM
fikeeeAabl/DRbfYVdl1Em4c4eJ4ZyLADaEXg1S7NhEpNJ+h51/MOAWfqkxL
LOCticoDSYtLsFNDlTVANnmSolqM/lnE5xxscj4KWpnkOAsSZvz84yYBgHTK
7hnTAPXjKQNLthu7J9XhHHWLn8cUBD3UVlfzEMxC2esOTHBX5iJ63Bz1m5qs
QfUDm+01wreAruVZbEBGSmWUglJSDDcEvOKGF5/xgce/1CPWBp02JkGzReG7
5QdLGnNzJvdpBe3DLl6QKbvY1Q74moQ+ED3tKeqcJCnfmsBQERrvewfjNip/
6i08nSRzgGCSn5OgYVqRkeNlfejMkj1rQy/Mhcht9biUNW4jCVw5rijgfg9a
XIRCUg11ZushE+V2da6wQuSt4DEi4BD0J+zU5/bAi5rZ8o5VkU4nym08wFRp
qdco0Dxn+8rZEslRJzGTYxqoZYEfzk9CGCG0tNf8Hr/rnpNKEt6roW+ZVLOZ
q+HajdddT64yRjv6us5nBGXudLD3JRFkglxmjGTiBfe1+a0cCpeO9KSV18mg
ym3ojuEqi6N8D0uJ0Rb3LW9DMLcotiTJsiE3P9wMRpidzU26mzU0uejnk9pY
iW6DkMgTWn3/NlAUShNpTBhKdwJcaHBxLDLp6XhjonHTdqYBP8FMs77VYZ6C
Ff2ukUEh+mu3zQt2jHBGv0xO48G0hamdItUCKZY+QKMVS15mOm6ECMiizc0F
PYgUnwfxCxgZkki1SVPWB7nsBey5xfgcoh+hknUYH2l5dyzCjs2zwAt0Svny
MD6ONHcnbdMVfTwzENtKwJrIJONFDP0ygsNfbzoJfldXJzAK7g4TGtxuUiCq
HZUHEQvFdTTpeUKsCx/fENpnfGv43to5NoicyzDdtxMeYBsAqW2sI1VBq6ws
v7QV2pHU49rfEKGJBDC93VUrxkiuCT+sDTbewxtJRhpqirr7RTN/pC5aDk7g
3RAxvwl9XzAZbyXbQ6YGkg3tHCXcrzYrCEFB9PNdiZht2kzGiP2MVMHVVwYP
nxkjEcq9P12vml5PyXPKYZ6Yw3/bbIEJGdNPJlSZqdkymfyWdGbe2SmWVXnp
h6U9LeFMkcOakgl2f77vTQCdYM0waRWv7O9ERt8h7wIUeEtOjQwGblIwOxr5
AAgex89mcru6dpT9bUlQRWAH063Auhyh5PB/xiFtN0NiykZMYRykZ/DwHvJE
BemlgQNftQ6kBxtPmHI7FU+U5DzlSzfvmKCgOrWuougGXtiSb2juhxuvXHdu
kcJIoikxrZLwjSKqg+PbueLQqe2ClQulnQDBY7Ki5nA4io3GO9Aw7wJPpFdr
JItu6Ph6rDZm3Kzmyo6RGVYiJDIV71lZnQ7sprnDs7P9BPP5Q1X+l6JiV/D/
IJaa4HpIn3/Ycf5ck0x3VRXPpRGHf4/Puw6QKfHkH7uZoeqoljbdy3Chrslb
AZU+D0NDKobCXKiQaDrccjvuT3dFpsA1P3zdRLnIp5ldDipw4TMuwvNMAWaY
huknr7espxe2ahOqaHbAv5hB361Y0G5ktZy95WccXQB0pC949dS2X3CYizEg
W6i5cY8KAFkRpOY1lODeK2fFvaMBcjTo4HlfL4MSXXk34l+z/cHHvBPcTCep
QwazDjj6NFDPPbtTbu6+zkO9Hwq/wY2Sl1n155x6UQYlxLVNEZnBTELSSdPc
uy+92JEmfHCX0hwdEyVg7HQMnkwX/rk2ghvDt62YdUTeHAjFJe0D5HOgTIX/
xBZUkNd30EVW2wMNPYkSW35Yggsbym8SiEgmOoZE35X4OerOS642xnm6rJbF
KvuJI8Sb8JV7o7q5MEZ1aKi5PyhV9xO6CYgSR8/Y8lfsNBgHwmGx19+yiq/2
iMQRIKncqiATIGnzgyRfb2ENahRsjr82jrj56wMgdbd1CrU9RVtXlrJOIffA
WRkeaP3z50plSIoVvfgxdthKhAanMQlsgYi62AjgcVZbNr/KJ3QapdlljjI2
RlCc8VXvKao1aJCw1fXQPgWqEJHKfjwd9CTIrZuPKk7QEH2tDayO8YHK9IbA
/qPyvF1xHCrpbNYLUnrAOAjbECqVRXe2DPwDeaplS8gYaeSIwmrzqYoJzFNz
Oc2967+LamgnHZGheX6x/JAxanjXAlWW86FciIBvbu9MpQ4t65seK4Z+ws6n
ZzuIfsoOKtdHRnnrIbFkyyjZmYKoQCWbUDpU5xQN2B1M7DFrVqUFqqX19Zdt
DENroE07AtjuG+l9lu60fSd68aOeY6iwGLCLL+7nolM4zgG2/rsYDXXiNCX7
jTUvBFYO5441oU2dI05lGXaJkI+FKdIo9Rlese0+eWPSljnzCL35DNN7c4yq
6hgfvlrlcV8bAO9boJWcDv0dwXe3TT0eTEQDjSfqi4BfXpPv5sQ4El7D+fo/
x9qJMCCgg2uiXe8cbPKRUiz6dg33I544Oz/vtB/ziNYjrPWHe606g9EVUK/7
d2FQu8fEK5ZHy9YgHveExlVwTTzD3SUY/zVgSxtKv0apjMmhafkBP0ea2DXU
WmVLhMSqoaqADNbtVWdbOx8wwEpoJ3XQZABwH8HCSs6Ei82GmffmlXiIyp35
ar38iHEfp7gtNviPplfOFzYvu7WeS0CXn1OtR9c0USJcTIOH69MPo1/SxNIu
3ETTryuGGa0OzuOfnLF8TxQU59xM4GzApp/xupQGklyQ4TLfC5Re2wHC9mxB
rkjMfChwpJicLTpmYWRsuzhFe+QmmEkc79aoFiHqORn73EYZw9Om26Ata4p0
m7Mg7fo3DbekvDye96wyqISvWeMUTE0FyMeWNOiaZTNdJM/0beew8wick3lW
Yi1g1pVTRUeWo3Ysd9L9kyZGmmlCDkhBD5owINRcnNy6uETO76qveiLGQ+mc
N6EpNVIx158A5wZwW9zZioHJNG9dqdxoxFZvZGRchtKIbnLM2Bw45/Gc3b5w
8jOISspLxYmh+B9owioPYhp9fJ3oWr+oRpvNEy4LOWLQgohO1ocCosue7Ibr
y3yVFJ0jKWUkKTH9o6rZ3KxRAeY/z3tdEPl1SwUwV1g/UzX5jtqETw4w7jE6
vr9N0eGT0v/f9l9LJH1myX9p9tO5trSrvrhh50zu87ksAj+Cb7E8liEt9miz
HZb8E4hbUIqJPkmqxs7vEfYxia7SMd/oZvAMp3rIvsW49VnDrBUkN6I8D+P3
4ebG2rRacLp3/OobXI2EMcBoeyLUvk4Banb9tJX/xdaHZ2mVixKpsFDv2mbB
DBXnfv9Ode7pYfvq0dZSS02NTwsT9Vgfq5c3B5OQzOf63Ly/KGRSf0LFARxq
JCfUiEfO2wuxcN1oGZgNCrUQgJlV6NtoH5DOvZuSj8LBwjI1xYkEFiTOErGQ
DGUoHdziHT/PJFiPxtOrb4kHqSFuNIUoiU/Gjx5WOqZdWHU9HrgTWLT3FH6U
OPeEoB6uufAVmyijHudkkhbLG/SY+p4Dc72fnTJ0DVnXrRwPwTUD/d5hbSTR
p5WSJm6op+Ou71pyCfzQMvUs+eRNWQqVNeOnObhC3o0WmpSEZGTyW2xB+g7u
Hu424h0ws6UzgYFiaSu9RD685eW12BwUe7IKdfAL+bNh8wavKz0lH2c/Oh/l
lAYU+JY9Bmn6ieE7ezbnzjFbEQG3d4opUt7GolcCyxK12M8wQ4AlSl5r8h4T
nSVF9ypF4pZk8gaw4G7eVIeZBXMR4AsTXLJ9To+LxESscfkJQcDonl18jIZQ
tIJA3iTJTgL4fQgPBfXHOmMx7W+gIO9YEdE+RPm5MrFtYKqW8xCdzKJdlh19
CHoIiFA3+Vx7NHW4oxUr1fHk5jxYkI8tSUw6s0cDxYDzi+gxUqenPmDXYNDR
E29HMEO6tkA67vojid9ymguETuKJO5xCGpRWpIw2Ip6bIbpvhtQhn+AP///6
s+ha/wMovyWiWqBUI3TNDsv1JiidlBFcRp2KEwyRwYjBo/jqv15KO0V3VKRq
HWqyXcjiYAVPdFzOAi+ZhKRvA5LKliv+E3VfXKimw8j+UPpA0upC/Qe+lus9
1SUn0mUv6cRT50Bi9cbVFHxqgFnbPdNDQvJgzn9VEb6PexLFr8FmY1VLxNWm
YCibZo7hBibXH327OunRO0vObm2Mcuw5nIUYlAudML9EHj5gllgDRfe8U1Ai
b4pSGQQ3GOh9wyPFzpRACXLVpuBvOaJWl1jQrW7FPApIaD6eMQToTUN8k00s
ERL2HuMqJhIC1uujm0UCH7vh553GoBd0fB6wXKc0KrPok0Dk6yUxkJwdAfHH
Ugg54u9YCmPpsArpqF/K+ON7ncO3asc6YwCqSz129tdeeJ4GOMNO1KC8dTda
dqCFlzF/utR9CwWF0ZOQlcK0ETs/MNO6/htWi8ZlAimAumww3DhC7Or/X3R3
zvJcqBE3UGnetUXpL76Sr5QdOopNcxagQ1ZE95Aq7SJcsJReZuQfkL4cpye4
jA//5VO1PjP+75K3mP7b/zuOFGItHxefaNxscKkxqjw1u/XUriAjWLtVKF3+
LvT+nt6/zWvnY/ZJqM3gswITaYGujH6iGKSN/LQqtw6yDDuO4HtsXpmzAe+t
DI2HUERIUQ8CJuyo96Fvyjecyf0gSret8qzCVOaV7oPKWmcO/Bb/AzMyLFl8
dwFZXVctsUsIRs+4YKLVTyu+kcpD6oNIcP981SVrMtyZs/AHC09w1frI0kBJ
PGvB+XSvCVdqXXEXuV4zpIs6phwqWolmhmLfIx7Y3wxASJtsc5TeHBuUKeJM
OFhTlb9AgzgaEdIhPYzwPdx9s0QG8W8WSKSiwfG0NFPBpaR4w0qw0VFoygs8
IbAx3iI2iNK9DJKE0EPQWPiRX0TeKUZStgvUPxr+eilY1jvdva9UsUtUsCbO
LuBEdH9V9XaQ8YSmMNJ+l9Z4IjO6S/qkRQqTMsulhcR54aX2HJTBahM3ZNs5
eTukZTzcHMMAQWRJ/WSCF76kW1pHVhgnEYWb4C3bdaLdGfnmeD45Lti2u5I2
Nj8ZEPJd3nQ1/3nsgyb3fAGNLUsni1qeKUtuoVhRnFUIFzp4OJFDe9MzT0CE
op/KP4OZJ3U4EO2NiEzvx+an8BQ87wzD+wrkDWBqPLBXAgvx8xFq7JAXglwT
YRWhoyxvHuBiTZvKrpn0WO3ajd/7suCkdWD/DEPneSvvaRPsejMzApthnXGS
DTxTO5NC0w/it0qOiaJkJMv1t8wD832u4IkpaD/Pm3QlRlnIlZl+6ZH75g1T
6pMUfju737z7NH1e7mVGubamD19uudgAUq0V7VU6VbNPLUrF3oDQUcFL9Q1V
JQDZtvXcgBaJQ1xq5fb+oEdN+Xsf8Xe65M4AwPvQlPHBiUEfKbUFGcLLEeiH
J46076JhfML2Tvh/6ZFoEQUz//quMeVH9KHyS6PcrhcUriS7mzOKgYgPz3Ho
ElVzCAn+vcRkNXDrkgMnNtZWBpz/rY30nm59QuQHPHVH+JQn0BrhjJsGj8tS
PeqH2+kjT6FMUXHtpqdD8212CcxAc3PyxOlEuTJi6cUbj27ZTM7OaFUyJQcs
rykHzM9cLnTidxnSj1c9el9SlQ7t0oTHtaPxRiq5Rb+9oRWctd1EvRmGgbZM
gmLb3kjXJfOku/9c3d8aal2vqHdkqMikojTQVr6NVCCfidT7Y58L76+xltic
lSoaCBqltsdPL81DkJ97K03H+fMOPqe44q17S3DtRp5u3gS9687ry9nkBqUH
UsA2k9Nm5z6qJl88NpAiKtXLJt04zLytftSbasuxpDF4z+A/lwD0NxFTWTTm
mdgSHdxUToFEHxaIE3/I9O2dOzsw1cUDkZ5tlimqfPjfuPoZ+PHRcQpF3KDz
JuigLkv5Uwo16+ePhkNo9uQvRhiz6R0xWP3U8MZvMvmOe5Lxq9eF/8SESxQE
sumuQZYfl437EE4D3ea26EcrznSVCQVuTs0pqrnArDRQuhu4oqfuen42pYSh
jiMTQvPmHMVvObRzNrYtSeT8y2+CpGc4OPKzUpD/adHf+UohleaPzb0VTfvx
xlHGyMvcVmMua4BJiP+OJJU2AW4CTpDvGLuLYYiXO57fw+7zYVJZrsA9akHY
v4TQG/qPiZAK/92FrropgsMukIWjsfSsEGt2oHMvntbeuQq1ohPi1btyT9Wj
d4rSLcCm54DHHO+xVf7+0QoRjI+fe6niQlyqE97dNbJAeCRcj/P+JsWN2bQ5
VEDsvcj1eXryL604H7HakaiJv+X/ge+mMEDcRzXOJRVrWchgMSDi8Qcyeoh7
QiB9QfHwPCaqonUplr+UZjZrFUMZh1QGEtQKKGr8mtBqBVsmtlQdALsRrFLk
XcAXU/0W0TBZU4oAig3CZmyYcZNvgE0zDr+ry/Eu983T0/HXMwrNarboO/4w
vVCYbxedyuefN5DF5Y0+4mMhvaxIJtlcb/nmxZgZnQo4/54wd3QKDYqzd+Wh
8OJHzFyEviU5N3BkerK8BKnPjResLkZGPmTzkmrPNVsG/dXK41cyGhQ952cI
9AIfOrgJvzruUKz0CxqLN7dFlwPgFajW/ROO3vzdfM/xX8R5X1Uj/6SQ9NDE
bN6z39wGhmeQ2mrk3yObsqUIjWbwQbH/RNxdWHedpqqaWrplydkF6baVa+lq
2kqaMkzIx0H0ueNHsZduIHDB0QoFdwv/9k7gr25+k4Ci3CmXgM6Yml0Ys3rm
nsjahi8+RlbIWjK7/sqrbweJnVt3id96nfc6Ck9WINToMBXyt0VcWmxhw9E3
5yydrlnAyyYD22y1UskGQRVDvnHi764Ai5IQMZ3hyUFCRIUtWKgYvyMpBj7N
FnAZr+7qXd5fpc1WnqT7CLwchIPG/Ahp+3qZRtxbVaWPhBJ8KJpdy2/KWyaj
l25Ce37Kaln8VsV1yQGEsQVUjWFDlZwEcCwPVQ5nWrEYFkD6ShAua5xHRTuE
NQowKF2lxcdq6kB2oZPLuUQ8c2yMAzJhV7BM/HxVdn0bEqWA8aviu57hHbGV
keENfzK0zy4Pk7ZEb8002xDzxInj/Z07gysvXa0F8pO4GmBc05eFOqSWu7Q8
GoSxixhm8sML7QpGGrJz+NAzJdPkLQk1iCwuNTQl9p7WOBBF5REv1mYXlY5n
+wIZ5AqsYE9AshmbHAMmwgecQtjjN13cNBy32ClsqpVZhtXpOkouogLf5/5l
7RHOFOHBjeR2f3wL7VN1j5OiBc3GFirx/gMJPcv75TLqQBocNvX7RbMFW4xM
mk7+LAhVHmoTn3aLRmD1FZ9cwXdWtaOC28ncC3MOO2mUeUfwDjaOXXx9pnGK
mN3w/CVol7nkyahZF6CbjhJhf0MF/N7D0Eq8iwHhYR2TmHPleyZQd3ZkOZ48
50fNmWrUTheHcAbpIZhTQ73KodCnYOWhdpn9ErJfEl3w1ranrITj1fWMe8n/
IncEvSpG6toTT9L1bs6Ao0g2ej4ESUoGQz1etwQuyep2Oh+rV6tp7iMYM265
VNQkuG3ZgTAvLl5mSHYs8MvWE74tAJbaefXm9YKk09BG4D1FVTzEKV7qLgur
9a+bR/aYHKFzx+UIUUe2hRb58IE+l3RPn9uOzcX/LTw+wWWQuKMrSR5FAvaJ
4nk78HksDNe8bQTnee+tYtNgT1hzBJBBqI4qYReVcsA6Q/nqCW6LanCOCZ9W
Xtev9OEOXRY0G1coPqgb7Zt3V7sxeZyXFhlE+x3/q8hvHVXIdJFhNzhiWRvR
CQuJDuqLIZnrzmY9FfSNaPfGR0tJ20yga3gMG0UjZUakXQjQ8n8AskEWIX+7
YqHBObytrdg7TpSdVGt60u5U5uMh2fRoVMYAaMCuPYMpyhQWRcfTBZX+uEGD
j1DTIMUGFXK5PKBDEyNumOFgamflUevYv8xUUAYNOgUpoPhKbjS81f/qVLcV
UlpBSMX7qAsWKEaaLYRNY+ySSb+24WtU2oYuUaKUe9uzD70Gx+7iylVJks4K
h+nZN8X08FTOMZ9iuhRo6yBD480tHH3yVqErmlTxSUGRO+p2rsJBJjSAP7sJ
osIrGmjm/w8ucHRfR3ZAbjyM/SdaFfk3sxMSs4piHNWk7inO6OAU44omVCt2
3Xs8TNoJpiK6r3c6i6Wewnjw7uTAdsoiAqudK/sYcegE/N4H7mStYPpGfeIr
FJkHAgvXZ9QgjjqMPQJr9/maVhNM1PrIouI/JK5s72RYykq41ZdYytEVXGD7
WB5Ht3iB34LlV4PXII039CDlhA16Bi3YIYdvGYCjJHdWxrXOcKAkRs1PBUv+
jC4fRYdRLAB4a18qj8EOu+GkJeKnIbO7m01DFKoIlKj2I96K9SNt4AEdzysb
gYqZhkDEJvqBWmSP8I3bBtuUbyefM/Mj48OpsduPpkwOSw7a2nKjKtXSIfVt
83BJH+Mg/qkFrABk/G/GvIauttWFDvyDrW9ig56R/pU2qbMO0CfctndBTqEz
kzBdwked0nnbH/gJHEJarGBSQwAU3Wmi5Xb2JBpRaIF0ekymifMoKVlyHiEI
3d12ytl1CgtbQB46B9NHfRHr5iOxB2WEzsZH27u+M5K9O0gWYYvfDqnFU42d
qNbaUUpgL8UWrE8x4tsHsqrYuMuDRDYZCCrmchFZc7wFYbBNoTPUNDxg27Nk
3iLKsRm76aOsEY1j5SCqd3/9v7kyLnJ1p8GxHalHOLLEdHVTBeURbXwLAyl4
4KUtAfIPzwclv/xKKdfx6FA8Y7FN8TIrzm8jFQ6+NRlTIzMf6es6s8/y7Gjy
V238sh31KDNFudldjBLi8xvu1QWOcyataGEJpqQpscW7i8JhhvNVfblXzeqK
DGlOqrkHtNoquVJv87xGw7vMGda3c9X+7+jzFLliEzqRXEWNkov3u/PXzSvW
Ltvmx4LjijOxwSaYkEgyvUB7u32mBNYfhiNVCQ65ubmH3ZQFDyz7Tq0bZZq6
+mjvEyugQZvsfp25c7ANdY01tlrd+DIbQIWo+TF61SpOnDFglcQifGOMxC0U
v8qkzQup+ef3Sm2CJUxRV7ggkzsoM2Hrzq/PZwoQucGQ6w89FSt/3CeagQzw
29tAl22UxzY7Kkk5ZlQqD9eEZJefqA3apbqgtp6QxVdE0OAFynuc4zqFrXXA
RLpQWK+PCyBZqhgHKPi+kdO58nUfPttwPPOqfK5U9heKc0IzsO9r6WUiP6B0
CEc3QjSejCVZQzqtwNCodqAMgH3wTuoRxnp67ohN7/HSNdafuN6lE2nf5n1h
NCMLHo3ESB6VJqLMTwYy+Ea/W0z2tC6I5hAU6fSS6gdsklBoOTQYJdCIb33T
//qdAf/HdOG57crl9dB3hmbbkisGdpv5IHoJt8jQ9BvZcZ2IlrXnyD1P2bqL
Ja4kmQ6z7pIqsFhsvjs2QHlcQhVZxXaMq3HgeJo5m4Pd8msQ1YZwIjfZ7zXk
7pSn1RxgLLMnHh34i5ueRmSQ31rwAcyDbsfu/7+Js9TFRQB0AYkJBG4IhUNP
7j9zmtStNg91CHAEUobUPlkZJwN5pu5gz5LiYdOJnv9B68KY997/8KkVUyLA
KSdr/tK7Nu7sgyEdf2jAGJPWNiigqfsARR8BhWwN9V8BN25j1inEO4X9w/D4
+lZHzS8NeNTsSp3IrZ6v0Ad1ndPKZt+NZnRyBIv6thtlAGxCMg05MgVvsRFf
IYOyrn1lPBcMZXzEZ1uGtmtWdc22BYnjD/PVdA/YmKHnbgB/wCmIxPQRs333
kSAgaKK6d9uN/2Kj2B7ROvOSnptMLCTuGy1x3fvi5rzL4qrmYkgBpNuOPt2W
3YJ7gKSpU44LrfAH0sdP81us9f56BaCW8Qe+/s60lf6y/MN/dTh+yNHrDDsJ
0ZWCracNo3MUcXXefwO9slJlVnmIk8r5ASIHKY0bJK6PaK5fAiLcqEfVe8JD
xc4oCqRLtb6wreluVBL3CpYvH8beu+GRPXVKYYxCMvb9SNwKxpLXiE/3m9US
s5QWq0GnPbFOxJaguoHob00f63nRroLmw45zlB6LDU0+lF8Y7t7ZN3xwC37x
bSRJcMc4TSmxG4B+SQfqrPEWBUbJUUI7q86Oz9gFBcRX22zxkgYGdG+dZfly
+YQKZBL/gdeFlEkKTz9yrUUizZye0dWlUwcq//FeqU1paTgUHOYwplsnoXTA
6mEDxM6hxH7SlQ8xdOOaIu7kugcJLUGYqwIZP7nAom18ZBqOiEpUb8wJAfKL
C0yuI/uwZIiayhEgoEv8kcqMq3lsPr/dJgEkPefhCSJB360vt6wIIv365/N1
8VEEP8jByHJ3CB1bzBE3ksdGkQcrI8Te4htDTAwz3A/6MHIuNyVDvvhisS6W
p+QQZIGkQwrIb5pfKniPvZNp2Ux64t/6OBGOmj2/Rwa8LQIqz43LbyeCMl+q
36AobcP5+WawBMo5+ae8k9hNeKRt6xbkB3D1ddfrAYyKMJYExSz1zIxTw7w9
uCGtO2vpT9unM3UG9Ne96uwMmvS5ji6xpVUcuFXuDzPvLhrDMef37u28PO02
bJMS1Ohs6NvvZgGWiD2S9KamLOvdfERYGzJo+DD7cAwevlW8STLH6zc4mS3x
AGNMWO24FF1kKyLFBeIZiTZPXjmBd5c1Mt077rZdJiQmYpOw1zibJtkKR9K2
qTPPR4NySNOrgJ2VAk2GyAX4cWyZGQHnDvwYfMO67p2Xag90F+8hdwZq6cWz
Q7AFaUXfobwOkyN2pzWEH5k1ev0lt+eLBIPDTXX5yqDM0J4+uVhQSYKHbo3k
62mhEVecROrtA3d0n6B+RLGKKU911A90raJSejpBKiw2ev/4FSb9r3kYbkyj
3s0qMTH5rq0yxrM61MkKNIv9FXBXr8Yxkqf1A/Lrmv90jdorwFx07DJ8OlMN
Y1xsFuZ43Wwve18QNOK8cxCvgl3gHN9nQFgtlYjHJ4Y6lPubeRFCe4BpKpxX
Nre3uDpbzT16xzIhg12j7PYR+/HBmsHl37P4rHtLFqKslTGS3ckKOicNHEgN
aX1Vcugz6ULWnKWN142cUHEVtbTj2KhisKEoA4VFAdd8Csm/fBZk8jaHN9AE
Fi7wLrq/b/rl9Cbu8ZLZomJN+C6fmWd8ToEjD84LUszIRdN6K+LaA15xUyCM
3wWcEP3pjQSNooxVU7+1BsAldF9cZQXFxgiTvEYtXMqKQXZc9uu+BKZuydn1
i47ujLuo44B1lVPNiy/62DGqNcxPwfT3ED3Iy+hRbZ4H69mNMKCZNANZeNUx
dbhsKeHKBDuxitOJWc/OVgfowlQesut84sDwi0EWQXkPH3SpjjtdX3CGG7nN
lnjHUwZ42A7wbP+wqvnIeQ3/RdHrHmob8bbiCujLnUgEyIlPGzvNvFN/FRU5
hhvDBSvCZ3/DmDlLBFGKCGvdW+Qi7TOIbfZ48JYaiQXsbAFLFCU/rMx5rw3a
JGrfTD0siwIe3TOebP9WVXURcR4szChKvibGYFw46efqh2BZYQD8swJCNE/u
fz3uJqbRVBzOqOFq8/EpUv6Aj1oVQbY+o8+x0+I8gxdoBjLVCi6RgrgLg4T+
TlrVEeMNrbNebZdfiSmKEHAsi1QvcXTzSxEFKNKfQBfrU6hR0vLt5C4Eqtiu
WyYRARV6om+pIbI9BS89J7keomjiaMUwV0e3xKsM1/IWisATrXUrLKIDDcj6
FoVyU11I4ogJhCs0RHmW3YRJQaYor6Q8sIALekAxi15KCKx8DgBqxer/mN1d
3siK32aetb1FjSfB6WM+LLgnF/Yeq6wT21B1G3nkqiYq2+/PJBPVbbCBG0jY
WX/PNHSSDPhq/rx5d9L+8/jkUc4HLApISlqj1N415MNhuE64OBca2Ny9BHTJ
TOIi2BJksUIBMXgCzjzeRJqIKZcJz0HF80SUw69DdtlPpzymRh4f0uxe1fob
0HpwnyquzfSRbu7C7ppRxwZwMuLGd3YdRv/mLk/Y8LKwhK6VeJ87K/M3lK2u
H8aeoML7OI4FAkYotwORJLmXjV5ewenNR2KNGcUxG4+vKWRQUndTQbkPeB4R
A+wa64EL9Sh4zsCSEn/FrreF6s3xJPoYxVTntwd5dC7XIKecihJenEAuKm6G
9uViy+LREPFsuWfXkJVE0QMsFF9pyidgAJdjVEz3msISB0ItHac9f/fYDUgd
C/ShzQ5Y5yWwJwH7BiH2/uDGyNMuy5w0G1zz3KDiMH/7hjPO2EKeteaX9USs
Ojw+Yqlv6Pp0HES9PhTpsX1zwOTB4wJLlVfP/i3CaRhTsgdZCB4zxmbek+Vh
djC04SNBtECkeA2Hk3oFbiHgmuQJLj3v+TALqfBEM5PvcEKRspa0vz/hkdOn
42jJURJLDZaz8P7M6KszUOrSyddoWD8cabJ9REXl6hj9Z7LXCbqtsTRv4bOA
svKoJ8z6cUPOadsGA/Vglzhm3cfddpDM7oixk1u/l5EZO265GEQj0Z/vv/uO
2/Ko3FupHSMVtA7/h47qUyDNCAnpYC5m6scXAvIifE/H+BjiYOPVwCl/N63O
ETicLVdn8ByaKG/b1ffqJPI6/fxqnbIPPYymp8SwOY4B0XZF+C7+6UPqammR
JYnew+KZlVCgRUjhGfUGW0utoxm1JYxFoVp77YJpOdfs21a0EM7qyAQsHvmt
A2D7SZdweojLX54y1hsnr+loNypIgOVQfJblW/EsvNVenVLxxL9tdN3zsozB
pptTfc+3jHzBTKC9lBz4q+K6WBcLQ5qunJMELOqioFojn+Cfi14S3Rwm7ZtE
+EDcRKyx5N6cI66g6aj7Y4x4f8GeJ+ZkLKoPfhMwyinChS8qSouxOoaUr9LP
6yG0Ingp2vl0gxVpDZMrrJC4io7k9eN9iMi0Aw99gBHqIMVTiGAbRTtVlYsC
3I9cbmhqVGVjFhkpYMMwdLC1L3419vGBCJLwYJQ4ZY4R5O1ggQ9xa5QTxjZ/
WvpCzZ5piAVQFMjoOpLvZ71w8bMSZuvW3iUWqBJKdBlEqemKSX4fnD8EqWu8
FXukcaXTUeX+EgLgw8zxuujJHZSEk44Vu4sqcgHDs7sZ6oIR0uuvE8B0Te3v
M9y8tE/9E6aEaGiH36dgUzprv0X8eNQIVV4rVoIQcI2g1RQq3V2lBw7qYj04
fGcZvOtdiUbUKSosPn8nKKqxJyjzSBUr1Zf8bwYUkbgRTQJFx8BuHERRc1lc
9tuehtQpXEew0D6nJRhJe86USrXfSRa8gSQgNAqGcjosU3dKANaumipvvtzc
65ZJR0XnxcA+pCgtaoqGGPLV3v/h8AZ4gumgIV0M7JcqOSDu94S7mJRNs1yg
LJ4C5wlfNFC1epCDK3Di/jyZ1y603wT8x8aUmnvRbjm3OSG+xh1LPV6tQNDF
zqa6xXWWZNeYP0sWHanueKHPraH9SD9+7SGQy4QeEKandIAXauVr+wLUVnaR
0KxNtncLddvRcLY0UIh0Re9Oq6txq58V+iB2q0ibCRyEbdmWJAX6YLIAz8Gc
BHCwGew3MCz7C11YFpptZDC/+Mk0f0Dv5zPZrffvpI91lXKVLrqi7asU09hc
QSwhK3oHMhFN36T34uLTs/iwaFpD/6KcPx/2bdGhCRNXmuo+KrBPuFl/Y0pR
zIpMefWwjwwMynMp2vgMlQ0wAI15SbM6LnQrPLkUnT27MQ4g9XMoJWCIPORo
3lokUQtO2rlqbjbem1pXpIiB/gOP4VbMibm6O1k9XwJ4Hd9XPdRNZ7mgtxlp
HBeCQ53SnEAWtHMW5QBVGRsa0aHZLVp803QGXduNx4jWYB51ckNJ2W6YXnSp
5IUjKN8K5ahgSreMaK5oJlgpXtqbKyZOskwh6QijM2AZ182zQa7jEqy7+5x9
rRT9viYOLwsNihH+20SZ0/AO3yWUi020MnidSjzraLgloAT7wI5IpVWK8+LB
K98I6YE2mSqSXMu0y7eMgXxgmMo+rwWtrzFNhd7dnfjWwQl2ihNMEJ3apVZj
zfnaxv/t3TghbS6Sz3XJJ074iU2VoRTdJSwHPpp+2hper8w+jpTytiNq6dGv
wjEqPuv5Qn3RddEx+plCaMjzH7MNbRY+zRsm7sBN3u6AlBRQX+ORkRJpRfkA
HFEywsQJyoii9evH5p4MvGBhHPpUnXkERtGSlQtFl8QNPSYoqmPgts5DgzE3
oTfBQBgV6Km6s7tBDxGkxC7ZKGGGvZxpZ55YFmnEMwA2xxHjSfSdiHg2BOn1
p69HHx8UIwIh2LFkHK/9EKsOMd5hvyWyf8pQFNC4NllxUewmX2TdgJ3k7W1T
pXFW20SZ9PGC8UdH01y6h6N5kTQ9d9H/IarN8FqvlZcytVbJ7vtng5L8o6Ov
yYuDSkNHGx+ayTbCnABOASIelTzVyzK/PixQwEXISpvEJibJB+T0Vegz+We9
lGMlXrAOgZa+LvcY07+r6hCVCpftYAazCJjtyScvbwyb3ldg63+LCPHFcln5
ZaTtEhZPtWTx/qMutOx3hTxAQ/H27wMzoA5K9ePhfdRGx56sATgnBZZHosRr
3vCT9fz3ZMdOgYqtHdAjqBplzSSyZ1idfpqYeDPP1mu7TQ4KMyuuKXghgrum
kz1vX57w5Qhw3oOvOiY2I7ZJ7JrjUP5cyyvMh+ZzxLW2ApaIdQur7RbQ8JAE
IXjd68pSbxLnJLiFn7aL23AIyGEk4TS9eiu3QmtTybT4dv0wvuwCAs43EGmG
CVwvAlDgkDbyRR2Ur+1BbenqqCtSAV3T1lvxRtFa+gV6jL7F1PDHhtIzHOru
dPLi7bUXXJA7GXRNg/qrhlaANsJiiSAgEhkbzwESrxYUcpgYC7Y92aijcDDt
IHQbdAzFtxTC/CaUaNOaimbqQkvxbgCeFYnwW1AeSO4Nnfu8K9arqZ+T2bIE
XPA1asc7H5TkX9ALktiKhRgggqd44ORiw769hdIc5PFIlP+0BafEdaZlorGM
dzSnnna6eF3yB1of3HOwDc4IbQgISC0kcfiKTV2qJ+XFSoWwKj5LDQqMg3hO
hcpOILe4emN5p2Q+XDBn3v+Mk8cn0njThQJrAHugcEBA6Af+i31ZinYiEVOl
72GCL0pHBLye0FlRgWjzxKj6tT0Kob9RS5QC15VxRPxnP30J+RBb0kBGC7vL
HuITA8fPWsXdicbu+gf2Ln8kBmOsylxi8Mcjxpul8wNHdzaxT+SdDJUwq2/3
X/Sff1PSWM+87Pft7K682hwN2G+PklsO2KldUl/KLFPVIE6dQmApBoZVjduu
OWg3vHjusySYmDXgJRDxgrEdhlPlyHezT7YtRai2j4CaH8tr1tiBviGtKK6S
fox9+d76Y54ljobOSTneikEBTFFWXr3K0OkJ35s881G1B5LDj4lnpgXmOo/6
jD8LB4QuIN/VHoykKGBR82QxidZcUoJxU4s7nSZt/NBfrA7HSjwQZRPg624m
zZTZZSnmuN/+yzurXUILA/eiynNlWcp3FeNihYkZSJs7v5TNNp5g4pf7mc6G
lXxkTc9HxPWE2fHP87vZjh24w0RTCRPoN57IjnO59XWS/ozRI0uzucJDUxnB
RCQhri1zA1PxhU/LRfZ7p1Sbr5z22ISB/xMRANNBhjDTLx7m64xJxT6vi5NP
WFRx/rcc60lxnCfsF+w3y4/VIAqudu4nlFOqXru4JO4KRkJt5MkAYoIhn4+e
hSE7J7zCfwYvini6DPu4jOToBTvg3TPr3j+qPh1IMHkNnctvEkxTXRQ3S2/F
QrWqEldH5l13OVJpuqC9A9DYmwhdAUOG2kIKpt6AbwOq1tzNkpq53EYlMcbe
t1sOJZjiW/QBm5SinI2SMVlObhm/cVxryoHVr7bBPS/HZbTGFu7YTQUj3tJe
fONZQa4wRVGzpL86GKl3upvZZsSbFx31lXqMjAF0HdQFZaEXHKPYCi3pfnxc
6ZJJxmS3kCBkuDMy47yd8grWk7csfUXe60xi4cmUz8hJFnaRmVtAz2p/zYD/
fHedjKSaxPQ83JJa/KA9v1Wz5+NGHHQ707RL9J9axwQl6X6kRGPhOri804+X
4fFWgbiarDFAT/wxiAobgs7bKDGWcd34o+eibF/jpty4dh6Xwri3pg5SpWdd
3T2EtaCIZq/lwLOk+Des5asMQC34T11RLZsFlQ0yDebbrcN29ESCfkYMh+wj
eN+3Iv9TXJ6NDR5bu5+1FeXt+VfSo0VKXkDg31gJwbmXtFhwJwLoo9ERjnjK
KN0wHc6Xxdbb6LSFjQlL6nGBYWNUWhlqTK+qMpHUanuxfSb8ogvnHXvs3MUs
QneOjY5WVT8h9MfmJTIdif6KE5z7B7uI5wnH5978Y3IGG1Yc11/0zO/Gg7W3
tihUh3jh3tOEuU9Nd64oFjf1uTWn3+klVhOY2/ANKWeIuVLj1n0hx0k6Jz+H
y4nRnkIHgjhXyusN0ltLcIHGwOnEXF5OudJVZYro3WwBx2MDt96lIaFHN5AV
zpbgyWelIKwfzu9kBoiShP+MHt1nTkhHBZBW7ZM7+KbZbjJZD9N5DPVh71sF
esKdBKZO3yGVN8IO//wVvlVO9Xv+TVahjn6F0fDO2eLT+V3f23Vt0EP/An1i
3KwtTH/v0G3WdBNHfQwx/H+E21/5pAvSXob9tspET89x2hK/grAnMNe7InA2
kAHmtb5dSyGPSHMFQepspJTMtBsrza8r51junyAsovSNV2qn1Jws6LTIjx+a
h09iKWUP/HwTdw+GFF8OVMVDZ8LR6YxTs7kqA03E6w0NkBLGkg1QwwXR6Qqe
HDqmXdHW8Gcyprt2P6hGpanvYjio2Kd6+gZb2VJfw9CNyYzsHzCTZ30M6WmV
GC11w7AEYtqqSwHDs9/VMctjFmwvxkQlc4TF8jOP/bq9l+tk6404seuhHQ80
1rasJ9f811SBPfjNqZR+BoPtC9Wql472AtFe6LF9JtK0DsP9Vx4J4fkT/EEC
bvSRnHOL0ZHE2X/EECqRWuvS6SKpl9KusiaBIuzIgNktp7aMId5dDXZmvL4i
Ie3qu4x0WiMFf6hSuNJf/2pdtLu7rgaewgwsjBov3RVMpJHYbMZT0fzOVgoR
NSX0plpmeva6dmfDGiwgyUYBwKSt3aIeMaH5dp7rTPYSkAZavMzUgMwDPlJh
q8Pk7L7TyDGFVStEFRAzjOyf0a6SrHGmhF84Eqz91mBR5SNJ+I4ltxmbDkez
fCYCsVoVA0g5E79xh1BlW09LUO7+W+ZcTAkzbcPKYcxMwaye/yCqs1UTDWjS
wx9VNk4esvf/lQzvb0RKQLtvddY5IdNm5fgFBQcVgq8jog1ZvafwWeaNTfLR
uzBBcE9wbyO202nGuqIzjvLQprsWwJUw5O8XL5cuFDYxuCkbIX8XiJEmCtvk
QG3B7HJ/I11qfbb1xEO1YGXBAENPhhSm/RiqDh0dBFeKBbnRdjaJ7gElUPry
I7qpIY2N93DaKXskvgxjozHfZuYgeuWgH1q1ah9bX8jbLs3NIqKS4j540Roo
9WmYjMPjnCnEXZ/PVvSe9zy76Eqgj/TSJCmJ+jPs59V7yGuZnAla8xGEUQMI
6B6GAuHuTz1P6uAjfAYNEMdzrqgyPzSczX1b12Tp1NfAjokJBtqQ23CLx27g
dP1IVZfcOgbduD0d3lLPYm2o6cP38T6kpHCMqM6NQ+GisPEXp5OhuNBDU0hN
tZa1P43SDrJzdFv9LyFyJFdDRY3g0q7CxCNKNvA9pKmGU4PiVE4Ti5HEQFAf
IPMP0dPNPQjwPF6+fp9s8KVVKNpCrksW5SNgN6OrdMwVBI1jMGZzfMWjYNSK
dSHvDzcKZfS6/nGjZI5a3Y2DhO9QN/lhZ4GzZTIb5Z/aT9KZ/wHL6Yo3AVKI
ghtwqwJ2TwNsP7ZE3TCsiyhpypI1lJJHnCtvtSPwTuiSYRmE2CE1dldYlOFD
6H45MEIrjdn30IKBVeiLUP2+0kiG6HJIVp7C/isKfG+JDRwNpohu1LIPW6ka
oAB2IJ/PzWI3k+f71Yg2R0GsfGzO8M6hdwpkTeKT4LAqkTizzzvadgO3VJAj
OszF9bI5jMUED+EDcrgzPioWB8D7LMNOUPM7h400m9aC1lf0autHg/nanAHM
RwXuQ8wthBXkgGUQLB6xk4zws5AQUUhXAPBbUL2akMdnRaN8/LP5eFwPcAA4
99lMDbdjVcLlvJBXwWQdf1lFjLTPp3prBBKxAuqxAMcRNvYhYWAuaXOMpQzi
f2AIGMLYKouDeQC0xR3lwEabEtGvpbBSd/aOHIsVF7uCzObIkuqGm30+fnKl
4xg6l3CTts4TJB1QAcM+nk0V7mz3gWhx4gj24GPJNMu+q7Fo8TKmtbwSbwwx
iRVSJKAi6x6cTlGgQyUzaeKY+5mEXcxz/az+QrCbPFgYu18MAf2XVq9JKNNL
8EAbBxPBe/Y2GUHIvSSYrw8rlR6IfKlRaL1JGkA7xmjnawAtYXCk/6fSdq9T
nRvpjUjUS9UB/s3dMZ5lb87Z7dth5ANALqZ8mVYQuYD2Y7OijDVerpKE/1vH
l8jlUvUvoDBSA/TLmq4i7nTqGRhDzwmuwMy2I/768258vtFQkclEsoMrEp0v
T9xun1BijgvDkgh/S+6zMDs1ROskbHoeafD2zhdGvTXHL6u0Im9Hitv3KB9B
PowGz3AQPeSdamgi+A+vs2ZU6b2Er6JnJ12eyE9YtouME5J2s4psxrWlpFRL
ltP/Ry72hwMF0ATILaYvGo39G5o5LTYw3rSjNrjBDgaBFOvYr5Bq4Egy59jK
e4Csic4qjGH3fX4qrIVoDzeQQRLSyA7PYocsoCUPa9uYDhiWmJMKqE2RubYB
rOs8vUqIJjVRi/4PqzXBbOZLXPmot9FD0wPldHAtGVm9HTWKh8M7ryK/46Dq
uem4PcNZKUDhACz6GTuyzxhH5ILnFsHUD2uiclbPfdCuxrUiH085Q25wTZTB
Ze9Jm9N6k9gdv6evmhYjRUvUDd99TVGwXeSoMzBAcTxz01tU60RIYXbNnsYm
sIzju8TSWNdmUzDtv5jDzhTLdYDW71tsexpUSJUx1xNOt8GlTR92Z1Z2l6dd
ajDc8SpVe1eO9tz8qMSRjvX4Xye6hfPgrGaLU3g+ITTGaNUNF0HIKiV71o6K
alxfmv4Kc0tT7Sh74kcxznqwH8oPkZEyjiBLq5yhTpkRdz1yHQ6iqzRwwkRt
2f79mhArjrroPn6OQqGLsc0ZeKDVNqDSLAilElQ8f6Z1ilEUq8zUuSjzsBBC
Hsg3bpRHLaLUl1oIat8Wa2FpUwwg4Zo3hcOneq3sYhAQMD32AEQhSlBnMzgP
ontVsCGVpha1gH/mCJpyUpdBwjHN4IoqV/qLoNjIGPw157LR30UM2r+Cj4e8
GSmhmb0mk/PdmSUkekMKD2SF9UAlXtM3/fwqLY1TvdN6yUKcOTQIP2dQUt5I
Ch0yXqeiv9LDCFpVZMxtn3UexYvduwvxqboDawn9HznMHGj+Hhc9jmIAQk+t
DEXAGGbNy5XDqCDO1L6BdUq2hUMsIMkDV8elglNp37NbQitKZXCqPyXr7n72
LUi3KJ+hDMv0MXK/aa4E2E8AIXuizyloxub5VMGodb1WHr8OwkEcm3fdV6dA
rfoLfVSp1AHio1rZHVX5RC/Rj5X0Bq2Rdo4Xe3xuh3aAqOHbLeQIzkF39ISl
4DuXLIS3KAGPgJrVzxmsFXEpqbm6OJbKKEkorT6O3gTCxXTvZg6ukS6VKBTj
Daai8xmDiIBltOdiwbqIDKsRYcR5V5eS2aSmQwJTT6FdR6Zz3SrCf+LrxS6R
yZkFMTBTfOzt69Zp/N7yRPiQegrZY4MB++xyGvLqkFDaLcegc5gOFEnmr8He
VBV7dneqZkquOq9nrBLaB3kqEEwPW2UUj8vmnXNRwmcNX+WdVLaSD5+DI8/a
ix3+/fVjfM4MOaoGBoyMqr5ZOT5T12DXXZNE+BEQS9dNrx40uVmzzgOu7Lb/
y8E+rKuux+zzyk9MfMxY75xEleQ0hiQNyc1DP5vmIoAIRxNZdcuQ5ZdUuSV3
zdvAciQ1iV7ddlAvKTCbTCKT2qiSRQHfYC45KD1ayRiXcIPBxotIws/ue620
2JxohZ3W5i31MVeV7fhvgj3Nk4zfYLPWnqDz9unoSfpfnTR43wlcZr6ac8SA
jg35ufhhNFX05u9NuZpYAk6zhjZEi+CEv+Muf/8/zoJWzZhMY4mLA00j9CWJ
FobEo2hNyoVGwUFbVmXDkDNd4eIggvJSj34NW5AZXfLXH4RROOlDXqmpWPS1
33QQCV2eTHENWvLvrTN4rB6RULaq85dX+DQjiGgimlKrrpJ0qqQMUgwwVkAy
w502b2D2yRmrgxZh1yF5LhbSw2PRCjFSS03nlPBr/2lmcFYfW5NI0OwQzyq4
+oILyrEpCRXbDld6mmqCUg6oIPzT388u65+PW79wenzUBdzkdBJ+USDrgcuT
GCPcsTgygEQQ1FEq2GSVzO5QYceSdjdZEh1f6cvwzQUaZbyhWdQhLlJUf575
/D6b54LnnCPKxzEBme8UgJsCniW7aTa9R9ZuwCOVUZMAXVbfEccb8YwEVEBx
gMYU57qDc2TfnZEBNhaPaPCm3cyFlamE7rg5ydEnkJwKwxYeuOfkkVdFnukx
PSzdhB10OcmoEfMLwNE5oGzDsN8Se2BWa0fZK6wgWI3XoLz+/yqnk4K0Wr3C
3ld+gduGb8Ji7ndp/6o+3NWV1PKPT0rSiSgFNpTm62apXaPyeeLe896h5d83
YXfgtv6VKqAo6hAPXUwY8c8YVFSg2AfHdUYrqazhIie/OXFt3BWQQR7re7P4
yQzsbOiZq5nm+ZTnljdMeK1ZKTYoLbMot21K1DmomdztshMzVNoQv8bVg7N9
YWaS7TE8MVagtHX2LpRRX8h69srMrQ7AuaDQJ1K6+NY1brfCLUco8yq/2zeK
oJ6OuaDgUWRWSfjhilKd8al3/lNhaB/oca5gZrUnzMUIF4D6ZxfAVV3vSTnS
CmjeR3CgGrrGmi++X0QaFyxTfiLQHD0FrY4VvuFc9fYZpoR6aTJ3ycYi03ER
AoiUc9VRRGwxTQhjB1GChQmCHhMLwj/XRzXqTqpZRlLf6UXjgW5+GvXL6b2L
FZKM3QSm/PuzELv/DqryBTRH2Mm/N5zolj8AJjbYE+JELHBaX5xaE08i2Qof
17iO107nKkwZRKlaOLC08qpxNDQIyzWiT7nrjclkUZGe6mPoqI5vjbYgk8zw
jdphK4cZJuP/+QSgvOS5wytvlcWur9ptlrops/LYOSAXE9lD3Otjoz6vx+MX
rfukWTDTIVuEnQlvBvdRX2tBbYZJ7OOFWoWw/nzsUyV2bLuFL4130+sytAga
jk1hKpX6rnrMzuAQffkKhszTYtq61bdsY/+k+Be80/5ucyXGAerV3TvFixSM
t0HsAIO/CLPdgPlBzoJBASqmiXfhbE8qDhH0qt94qIwnG3hqg17bxzlRtpA1
eTFL6uvZm7xUjFWgWu/UkfUV0+eQr+/BjO9zPrfgg0ei7QP9/7WfV4OsYbsN
dP7H3Hd+MD78knahj+ZVH07qKRkzqobEk6gJcebYbMY6DU6AgwvBOwkfNOtS
bQewwsWM2cY8LNC0isCrLLrKWx9t9iSzUfTxnsbEnGGxo901ny2+gIbeoslB
yH0LUQYsLUGBoN7wE8+O2CMXQ8Pn0qrT2h1b9LDYI+q9cNnwlH6F7WRvS1Fr
tCDdoF62Q/o+QmX79QHkTT7oVVM9xFfD1BoNUOBqDg5hnuFQP2BEkSosC8fl
XCgVsyIJ2hpAuMHywd9VU12aMAwvsIHQewncx055esl69xGu8ttAQajXCmtv
rxxGHcAUwjcU/LIDAGPSv0vf56XfPNKG7fnOj8bfRcIF9yvH2UEHDxnJIJ58
Y2p05GwI5O607c+tyV6euQ3c207k9RzorrZf6UQdz6J57Slo4s90+dxhsWGC
zfzgc2udySsOmkYGW8lDssA+EeonLg+udmLE/YKfOCV2qCpA3d3xaVDgNK3Q
2NV10NaZVQuVW1NGyfGjGs5Ncxifco6YB96i96F8zb/1CHuFtuMZLgarQRA8
uOD5PNBt9KoS9j1NpUNDJJE8vSdeS2uGKl2twbf120BC7dT7RpCzap/XAtj5
7Q0or6CRyomeR922noeh+8pysD3k+HU6YHqelaMoobiKMVXD7pRFr6HUqnuT
i8EL982ODoOmsmvlX2zFtvjB4ZQf9KnVC7eazH6oSBn6gUJxQYtfssO0bFn0
MdmvqkDxDEnWRVWlxIkl/dqgKyGujfl7UwatpcYf/+pmMnKv9kBmGLVS0HIu
fbwnAdEhCeiKVXBuPglam4lpbUmL1f6OiazmTpxgffyWPpauk5+WG0kL9t5f
/zHG61TKi968nQYakmldz4DIGHxDHLlaupkgUokPzi5J3ae6g94ipgljn0bz
cAHq7OLuMmradHzU/HTopJ9EjrE+TUacH3SEtPLpIRbSd9s1Qc5rKi2+/VD0
6wzAbLGogKXsMkwS1INTVxDdf+E6EVgPIoYnSBshD+5nXdYvKnLmtthA5ceD
ofWrgjmRPQCJ6A0hfvWajvL4u8TyT9dFZHQn6dC2uE5DHQH2mkdQg4I/bB3/
kiQAVXp9mmgNJceXK/NuhrngAxKgzTqFYFmG96SCqt9t1Tukt8Nkqvq1u6RR
8WxFFRBBK5MV6auZpM8sTwxcPe/HN/2mx4h0BR6n6FmkL+VBTvWVzZmJMyMM
grKGG2EluJ/8VE2oVLpMYrwAaMEvO0YxcBzBhAGPd4mUdtTPktP/vh6AB3Fl
3e7Dv+Fl7THy2fydXMdvtbVS4YRCwhH2PBFMDD/oKIGDzbTPUmk3RYB2hOf3
fXEw8GPHFG3xgZbG0SKbZlZ6NJ/OF/LaIyHo62pjb81urn9jk8XMwJq4tDET
4viQRsmgMftF+wNVqhS9na2nRnGp75BWMLf6uVDeYXCmXhW0hEIbKluiskRj
RS+r1FkKD5vrz9tBpliKbK6Rrh9VDwYpg33P89VBERjifeC2EgyBr/qKD/RM
pOC7XP7TjW9WmGwhs/99ZFAksgKlbOjr3wEaYTey4fS2l+by2Sg2SX4+Cs3J
BZtw+PRSRKNWFNskzXNy99O+Wc4zha5JIMMsOVnS248csl14MQik0T1E5hgN
Y4KkoT9yzja+iALKQGNR6fSZvKOt0U6DWs4ZfuCOPaUaeM8zp9niLt3jLuLO
SczveeayqWKINuGzwjBgwwJpJynDiDYwsV0jxP0dK12NpTLt5Ch3SUwANQyX
L02gKTX7gLk0BeZNoEm12HP+N9DX6no5Xh/Ph2QfS/lyb/HLNiM0uPDHrO1f
SE29Db0Fo94p8jByzhE0D+vEB/FwlOd2JQMuBsIXZBuUCL0rr57Sb0wPdPjT
2J8LwLSdBf6/Z941/Rufps4RHVBpaObQiG4uOA0xP63J9WqWZOm51rOyoe2q
6jF9hUlPSYgmlSaqp7e3gK/vjekM+iJ3HNuEeuIdgK5sSkym7rzNVbM+mPuf
vPICZIucMwIxVUJvVfXTSev1r4A8JEmxgwtRCkLtsd4AMEpnlqqYZKFiYAbg
LgAvUcogv+s4U7BRFduvwrhk9tmxT5MBplEu5dCgD+rkniVq9DGrDM/wXDRz
/Z5QouQLFwsQjdGmhLTIIGIJT4AqSxdmXCWTiKbPrLDJ8LdM+zYiFaT5Vnga
37/yS3rQRbhRQNx2XbcMif86OIlKe916tPwkG2l8EMN3hJM/yVRvgvJtR5i0
VBv0j5lr8sao7Xnzv9Sj9KVgw0Q18XMteZWDSsNK0FTg7W4UfL+Ij2DQ9GJU
YLuDJSXNLezEGbrh6T9KqCXgSJUff3AAXQOsRy4YHT8OY7/kbP4Ad082mV9k
Ypunaoi6C0mRbNRpoP94V92mjNJ5oNuLWM3J/duFhG+M4onJLhiV3xJuiT93
HUV5Z9biD/tvrkmYDG7EoeVt/hMJhtUbAQP7lZ4HKtLGSSniPZR+Ngtny2JQ
avc8xXjR3Djzd45WgBLh5wTSNO9o7KeXlW/fIdupNNp+IVDvjHfHptcFXjPk
h7kthzvcb8N+mgGxE4xhZ/wpKKbGtvhWxN6ora77JGeNWEx6zWy+exxYyFZt
2I1BEMZQHrPOr7HPQMk1D+uJy5is9OaKYG1KG98aYB4dTVN9NsRpIYidLRlQ
q1Tz5xXl9nLZQX8XXf6DPehRm0MukLtv9cMJTmE0KHUJkGPYuuigiw4ilqBU
j/yM0PJeCBRrYYM4l0X53ClZrM4FKYEFFBGP+uPzZMCA3KPncdnmG+u7uIug
hOD0hU2lF3lYLcEA0hx2edOLOuRwdo59WxaqYSvtWfct5fE/V5LmMwPpIwZ3
zSANgcOITtUfi8ukYUM0PGjV4wv+JQL1GmlNpsM3ePz3guPqccSrAWcxDvdp
Uy0RDOqSD39YbTTxtbGNc/hRQbPallPAwN/Kvxi/Jya1xiMVUsyQVUKLmdOA
50IuHO1E90yDm6RVYEbcxy7/eOyoWg567wFOFBDn4tlcLWmJdzra3rcL8hV/
BKkqp7JN9aty3V72zS2L1jXkkgjjwsy9lemBG3ipulFQEqNnh5mU6WiRBBbT
WSGqLA3kvfVYdM9RREMy+SRD2dJJvEIpSp6CsSGENljrAYXuBzkrGa4r8sDC
cACu8TziaBqI5Nsm1xU4oFPwcKG0+CPejx1EI7LAFZXNIand44XJL9lT88hB
BoBwTjlXLonPY4tx0JcwN47ZrgbIAuDP7ff4k13Uq4g0I6M08VS8UMPy1nS6
xPWj1x0VlyB/0OjsHAPG9PHPsKM4eVria3/6FyVx2uNx56rryRPpJXOtCRCC
2gobQQQIhylL4sQlRn1FMPZ2mF7jdpyEhbk060EY4puZZ8dEjjnLFF9tnpi3
SyapmksQOncBMvq6XeG2RG+oLcJYqu+8i3aZ14KyWKxQp37AjZrL/b0Ixtbg
4HnyOEQOFQCsHylwrU6KFhOB25BragRWvNjDJmWky+Gd8RQKfPzfPlBiOiX2
1WzpRTc+MrbUEZVMcc67bgtgPhJdK/8NvFF/PufiViWmbUBUItdDH8+GMJD0
kgaoWtTo+37sFhAQgSUjH18oojVMQGFHHKvbqrUqt6CUz3SRe/3c9/9GPv1f
zzTl0KqTyJDRQOs3+6gRjGcFS2asc8W2bTJcaltgrLqUa8Gp1qNCYWL0Jb3k
s9B3JEsJUXr21c7KFNxlGasSiJvP61VWfmeaBHX97rRNv6+Kkpo7kwz1eZG6
FnPGXyk5k2vURbYjW3hJo3g907IPXe9OXz1h41LB4qsw4oek3Iyn1C4Ge0Gn
fZbZV5cYDyumC63Lru0ySb4VO0nT7pqNZ1XVMrQ+qtbY+D0HbKdMPU9y2QOR
vWOiUy7CT/POBka2sew5I0SWUF/zS58G1XEzW8UR/GvYorBy74w9VpKwr7nW
HaDGJOHz/mBPiYdVVODc/h44uI82usapJDLgRqA6qeQ0JGsIfOG/U9fie3sb
+/DzEnrAScQFwPB/zKwB21vp45u60F/w/v9XbIPK4gFwZ5qiM2ez+WUTiJx7
4WtpX5a4hp7q1BiIT9dVJP/B8umuGj+GXZXLnFuUOfdKvIsVVIFTUe6Zz7OO
DOT1eCwrTV2DVnFd0yDsptFNwFfvgGHMK91KZBEVdz10837/GRkfxfBtMvHR
D9VI/0cJ8OnBm7tLF/UXjckR1YSIxprO+vHFUjg6M2J0y2erI+RQz/GjGpz6
85LSgk4l309nEmlzF5sn9IUqU2jnlHfK8qmSPzDGF1S2vEbBEFpuJgd9+2jb
/UH2QseQO+t6fw7G3xgGEE2T6ws+XFkGUqA3/KgwFXMp1xna6F/BDUTkNZQn
RLreeU9+dcZM397HiCoX+DezHynATBaSm0pgSII7teLM3SvbP+Kr6NQusoWm
kcVv+A2cjCs66aR5PlECs/bys1WatlXfp0454dGlajKvG1UtHSiXT0FJQVXI
6/4tqvI4ECn/vLDdcG2iRF4Dyaa2SZoh2EoSfA/RRZhXnGWI5v7+wCLNW6/9
tfu9DrmWsnZc0m81ga7GD8YJxlJzfNud+CFoIvyHiOmLlKXQIwXvDxe0qVVH
qgKIvjXq5+xiJWzubt9QCz2nOm7vXf5MgEwSOjpcZdTinO9Yjv2f7WOQmqwF
UIEmE3JahQDHuKVzH2a2NaQ0sVL7OWAxo0qBltfGrS2bXMCjn5va4OMI0XQX
0a5EAh0dN/ZGFRbVvjGFSec0l88ZEhztlaTLj4UzbLokm4zBm0qIEL4Ebyhi
+QaZI25V2fn2KCaI82esmIGGFDVXIUKFvZmGWz7ilCUEFoDWyG1ybuDHBp06
sv9QlmUWEm23WFgpSscN8jrZRtTrp6tsj8Sfdx3hsFTHpEaSO6d7/tU+AvQY
1e1fTx9wIl7MoxDbeQ9Lh9DjWcUZIZxBS4InYiqEjolWmDsIaizg9ZHdO1lX
bvN9ZfSqB+BwYbhkVzidXEUFe5VYHUPR+fadoyDwi3nDGP2X+5HVQFhHzWOf
ZV9WnKWCdHigYEELromt6G5/VRwuWXq8RaduCG2OQ3WYKTkiEZhTZu20bnBa
FRFE+dWAtBr/4azWzA+1Tmy9avgA56y3AGpb00OEQN4655I3i+Del1zUC3+C
M3K4Yd01VJNTZD6msJsVlIYyShq6brWjKlFjdQfOuNlulE+Ywzk//ZXycoEs
QcP0/Q6SrbkylMQrOKN4Skgh0RMZr7yoUQLVGg0Z+nOgmO5TQBvUNHcGTrTB
xRuLiosKoKHjC3XKbK6O2JRIFqUdhXUQWrrd8DNBWz/wwn7rKGqUAW9tPpLT
jYOwXE2CyDGhX+EoxfGltr/DTmVXo35/tDEKcNgICcGz7sKO5XRAXFeOAInm
FSaGVD0aq6t4NV4yfJOY0RqcbQpwn4JnBnct93wOVxM9HryklEZRew0DHszL
842p2tRUlkVtWfUt8A8tG6DpeAMJilc+dlYSXN9RAsdwkWK6BJIl7laBOJEO
HZgtWQDBtXdRApBMcQ7rvvyHgS86PQnlKU9CD5Q2uqaPuBBxm3/hVEQLjYPI
zGMqgB+UkZLxxZgT35xfJTWnJO5z4iJbk9QXQCSl+QxeEXiIxKCN+Sg/rypS
3+vZCHu1CyDy49BMS5GZdXtR/va6PyguOb3hwUHv4Bh3DzyGCc6kW7CAjI7c
KmYMzHclHsI6eNlQ5mzgMDIX/YWrt1SZrn8Ke+YTEDkmxRkkKero1/mWIuZX
XbnNT2umtkqFwphW1WDuhwnqvxOBb9hMGfC99FwTdxVHxInf57Cs15EKNfsW
IBnoZKFvJtVQuYWeayDOnibAWsLX9ttCU6Cdttx8PSz1p1zFBNtt38oRVqNp
mZfB4vhSRRbIxX0LUY0kvn/ps8t0d4Nogku1jsnlFAsreuNu72fyJoqb/ZRT
egh9tIPpFN0w+qqFZohL0QT8SrRQ85NsqcCk6WOZhId7x37sqQxXKtXKmndf
4JAyFg9KWmkOQN0nS7JMQqveljN7uRF7V+WNMkW7mLlyhSgAhuLNcWlmPuNZ
xjT1zaBq1Z//0utFu3S5AJpjwPuVolP1uCc2fM4JxySVpZsmoKK48XSINCjP
QystFiUjX+dshuwurGJ0gWvvilqT8zb6nwJSqD/k8xg/oUwk8cNTOlQJLEHO
KkOlBjiGBNOGilsyot6irQIz1AvH2t7w0xJqGSzn0kgflYqAn8tWoRZpnG6W
6oNcTnzOmdGsrhtZHDRUgIhdCenMDQkFDguiLnc5L1r1YQWuApYhi5Dau0rl
3FOB44mQwJGWxK4BQK2WPdmZhlqfXaivQkdO9YUuHBQnSpJwDnJgGCa5jit3
zasdRnPHhfEb3scCjzGmB7KMAjKB7iJWErdINlKMvmm1XqqAwptGkRg3wBtS
2beHkxDKm8bfoGeR0SjwRM3Jj1KjRNVsxbHnrRNSqhyFPVd25OGsxOf+SIgn
smT6HlJ5aZ6ekvNjHdTlhlLQOslQBZWGVeatqfyJapfRHu/UxAx79kYKmmlQ
6i3WnqsGqXak5Dwy8GyM324DWFE7Xx1JTo+P+Hkas8TwOTDJOrcP6XQDipZy
lWQRKK41dJd7wZnlOIOGGDf1QQmYcZym/AWMsB5Of7dctx12QtuFRRELBj0q
wfAVKRP7mHdfiqhE4LJqZYhKmYP5LA2PI8QySvTySGs/Lt50oeo79NEB6pN8
7IXJ6a2nhC3T4rBfU84M8N0lBr3+VsI2dS+iKhXSNQTJ/83Fq+flsk5alspL
0qq3PpqCGLIf2G2P3yrrgeLKlJeANX0h1ImvfKAH1aCZulHz0QNM2YbnFj8/
E0Bnhg4qMNbyKRgocPiVOnzdw+N8mkb6avGcNmuk6AdK8dfDRjXdVezwfKyC
wYgzDUw5/Bm8eWzQyiRniEHLRzMDMyYCv9XWrd/VQv9kaxdRK0gdH9AWnYPY
gogXmwxuX8Z0bnrqaNmO/zDwhYSr20kSskb/zWQ1q3AlTykdSf561NQVyjOY
JRLhjRdSlxtRsxmYbUqUKpTw/Y43kdrqEhKEQpJQ3XrCG3bRoHDmMa9nj7W7
/Bcp15rsfQjHnE9tmTS6tFnwAWG1X5A/sQjdmkSZswq4gElPLds2vlWaRjK9
eOj604Yw9vY3CgreUqT/wmK0mWjmNWMdp+KPOpNVjL1KAJx71UhODYcR8pji
EDJBTKU8vCh/Nyl2Aw+smm/yDorBMGE8iriFN+lU3mCbHhI6f2fsYjt/xJAo
uiA3S9XD6LMssi3IN+jqZnjKD63Umox/fy/NSPo9/3itR2AxzDe+t4bTZhum
B/Yrxz6T1QbEOuoHzcrCrtvQ7v45FeXLy63FHwtGkz4niV9OC+Zd1GvbfJGX
tB60SG3EIT6wM1nXCbJMEYeF4nZeIzP+MmH0KoBKDb+UssXX01ptCRVVxPOF
uLfL9LdMguWuZW9HDE9YFk6lJyoF6ANZLcfGPUrTjyX/wPQC0Ar6QEv/wSIs
AT29+yGWNq6k8mqNGB1SifTa/H32XN/HvxZYdK5jRsV8qC3Eh6K/qqIezoUF
fbgXM97kOVSI/WmL2TwQ5N05XaYnYeiO2tWBVmtGiGWHRnjvCDxUZpJqrdZk
nqPuh6526I+wwls7+ndkQj6cOZYYMXIMBUlcarmo5fvbu1EFiBKIV7yN8/vx
Tnt5BQSkklxRIwPoeqAzrI6/SuLd7m60AffiyYVL4DWxhtjyoL6aHYzAt+KB
Wz0W795YOS7HLg/J7NU2AS27c0hEbur9Ra4BnlLmooDgXr5k9d2M8BIJC3u5
E9s8xREu9QH6iq2xkOWoanlTx1AN4tzbJmqQdzDDhJZHjuqvpkoXJ3dfrUmo
c01dsP+Z3ZCKb+IcD+DGj5RydfDSzDFPkZe2xEwLT0RMCTtGWvyKgPJG5CVJ
VXQqPP+GAgpuKE6fTnVCUUxtc/4d3Vqsu5mA7WQvgQJtku8FzWGCIkd+wj1f
fX3GzK/Eotx4LkLP/cTzZkwcoCgizxWrYA8zVvo/1uqlJotpdFOaJ8IsPC93
kipEC8TgIidzjXJcTgmPNarj1195Sc5FmrpDIlCkNZu0DHofqA74CmqOhShQ
ygaXxwTzsTnzhdVjv6GQcuDGg8JVP3W0qKHHeRe1ZcuDK3J6DRV4h39H+GI/
fYTRg4HG5tkQ9xII4/4e3SGQkmdHdpIsCphv6iCilFgxqP/xPSnKJvCeapeC
o/DSJoT8bIg5uWhOtkudlFGtvmnpWcVGnJm441pQs9mdODhD6A7KBT5lad+q
ExKdb1/rc6PYBF8DsQxsrKawYmHm450p4LlkHVznIIczn6gXn/3N9Npu6uNs
bi7Mu+FfNUJHHeH8Y9kX42Dn81EQdtnxSabKXQrGC7xSscEr50RvJ6IZZ697
lpCL9zCmgXBpu1RkaLYu4nmh430iBJuayjcfLLPqjJJny1fKzxuU38r5Aku7
u70L0gl7JpbiNX7f9CrVyEOtkA4AjYye0z3aGElNfRk+oC0qOpm2AAUFF5Un
uI9twekwr0il1a0Pyfex8FOdoM9tJYTu6/hwFMfEWT5ZjvpODniF7OxG60AX
UDqxhGbVz9K+fsZKjxJ8D0UG1wt4Bg1nS7hN7tqZMKZiZyBHr7ZnnOLme07e
zeeUFwS9E3OGUkQog6xvRu1rKc6FA+qS+GKvvGOpFk1vtpElVrVfo/OLzmKH
AiI+CPHdlYhsjmQ+77J55sMGfrdkeu3aH2fAZdMKHKPD7eg0ssRTsd5Nwjg8
h9wl2OU2VDZSoRA/g4K8vpNh+fLgvS2JLg7pYBBH2J+GFC5gFe99Xy4Y+H9O
xwKECBhMoneQFMQxSCUIJINc6PLZ+ke1ivlzhrewbitcc3DvtfBIihPv0MWM
2RWmm1YO2xgrMYTVJADklwB6bhGrZvDFgP4/z44nPs5RkE1mzmVZb06mouib
ZtrSJUqaIl0UwUQvngU0G9jgWBsJ2S2iRj3MKNJ2C1DioTAEFWqIW0s9N8oV
A68wBvpmkUs0t5iGbNdtTc3BI3ucIPXMJhubdAsQZsooODFYtFzP/5vQ6MLp
6oMG7GvbTARIuD+HRcJElx+3Wgst8sJjnDsssz100XeT0lOMgGxaYeUaRQG6
FPj4k75vc0D8gnWa8NvZrjrdJ6q1ovkVhZHxj1i9BpEdiUyHfqwbSdK83WF2
ZxnzsH5h1sMj2P+cgEP7wlj0BuI5CXVt/RhSFrS/gC4nod+z+GxboDiIu7g3
DSqYHghwpM5bUDxIsVVQGxSfS7wf0h/WOqhC0M2f+spcaZaLhVh6k74GXzMt
hPuYOBOdjfI3NANBuLyBv16OHGjskucjrI88Zlgzceu+zsl9Kr+++AHBzBgz
Gz6QHQMtNabOJD72PJ4JKW8XVB9Rg2FaOBvOR/sjRv6bOMiBwmMxClIY8jfT
XNgYZyS49SVFQuCCz8L2n5p6WrzQBh3zkzLdKWLi/Jqduygsp6zluzbx1RCT
/QE7/CS7SJaszA0v5VYlJTVvHFbBiuQ3qLhiJIS8i1RozMWamCjw9Q9h26jN
+AWffUtYOHKAsxJHFnj/YugsK5E6V9mHbH5ynSNdXQ+PtvfgR2yCBqZme5GJ
pFtl7Ba1ag+YRnluejbUOOKVoEQ89v1zmh/De4mOlA89rUPfJL7MLI0gGgAH
ZiXEniIRXgBF17kHb15y8PD+hVQnr+eC0ok/0Cj6rJfVbiGMbt0rq7KGwN8f
yl9cuK8t+a8BlIlCClSi5935uq/dNm4P9Q0333lPyCOlc17Ij6NCZcLD6rzH
gZhgOKJsx3nU+AKFb7GcvRiuU/Pl8DH6Gn1Vcq3MWI+6XbYUNxD56c0vYFEw
HrKQ7v+nLA4ImeXbwH1bdxx1CWzsIi+ghFvSNvzy2OfX1rJCRWHgQJOxL+LQ
WG/fpJM5flrr6rT0ts1O7dPn/7WrbUoIVy3MzjT3LPo6YN1QF6isBCb7NON7
okVt5DVeq3SrQ9Wf0izBrPcQ4ZPZ2KJowXEMCWTUIPYQ/tR49wk+qIhsIsRy
y3XqeoD9Ux63YxvKYjWuMUvbd6kBxGG4qirWCA4SzGdVDBQGft5oNCmIieP2
W8R66Z4ABTNVvVUxVBDjG1Hckauicxh1qVhCn7pRWAArIpIS4qqHeWliK1MS
99cQKhjxjEShKtEeItKCism/A9Ho3lCVcQ9gQe3sZZyn9Xob9VZrQJ/N7RGZ
Hzk4bvXM+/x+rFoHsYqBAKSM5BuDezvKB7sj/gZae1I3hObqd8NIfQCzdlvb
trUvob8lyLR3TmW6d8LZbOgeiDUCO54qUjDLQVsOVGwyKT5oU5/dUAIWZoZR
N22pm4T/vu7q6CUurOrYxnPoHUNNmWIr9uEMR+tdCk1GX0PO5R2TAbqMXKsB
14rbhgX4rL3kIj9FIm/jIQpooeGHREHXHYKOk8+XHbA5V/+uAD7QQaGM7r33
w0pKQ473mnKmQs1nS5MlzB5NqVbc6wBcPJATN1Un9rqPzbj2WEnVR5Mb7Uha
0MsJ1Sv3bfFJk9D0YGLG7E9FG0cg6gG+yDX9c0NNedYKOGxBhk3WBOkZPP+B
KBOIhEAKMJqD1PTw1w1bObN0Gh2yQVKSE3+ZKJLpzekWBHrI9L4CZXWd7VTb
QBULYl3cVWi76HHhWSbgbiKVa93pWFyqaMstuWlXS1O5wd2ee/dgoEgy0el2
bcGEW7UW2nDqWHbvlV5Q7r4uhkLwaOaVGw5MsHW92JGVzgTyw2QFBLqRreYy
+rRx6p69fiPd9AakMTI+dJj30sU1fRYUQo3XSCqI06gQpn7P+VHqlGGn+VFs
gTnnV+Krq2/ijdQlgyNcG/dKbS+7pEHdAoUCxSnBzGUKh4o0vXeHxVpElL/5
dVl7rNVa5XEsanza2xh5CQSb22M15v1Db8p/T5nFuL6ffiL9VwZ4xhR30w21
iZ396g5PXGg0Z1qufIjVM2pN4z1AR0Kch4pI4ZbIaJR3OE5O4zv6aeQDqs+5
84mzWQPWlqClE1vzTM31uxU3uZxpZww0keuNvjSomlcFJDNZpVHB5ICcd0Ko
oKEQIEoi4zAv4b4PhTyHxPkM6LvsjbmDdCHbOYER8mCMMuToMqM1q5k4gwEX
1i5+8UuK/ep/EqHtVlqb+K+Xt7KduUHRingfVGjLHky36gpGy9K9rfbskUQ0
IThGR5f5PsY23TtvhQ2vW9arSQsNDivU7iXChOy7aAp7jC6kdw/nN7mj5LTq
+1pzHVZK4qe75dC8eFsphgdBWUHWBLd/j8GgRGrTMvWI0zgNE4fPTeTICghj
hquI6zurcvZdTPAHW5Tm7NXmzr+hdIT2c8KNnpJ9UIN1C+/XPZyIFpoSCb+0
dn+EQ/YKUavs0dTvhSC29+xTjaEJDdjAfEKVmTQ8wPgMPXFgcXJ4OHGHP/Ea
kwhjGnK+TbgZ2sCuKDp8YTIaNXC0k9Xd43aEEQO8scJGQdHEWHCFPiHcoHAk
CokzczhIUONZEhZYGgSeQEpFV6O49i2/GZZGcc8jP6RKgvTgpUHmbe/oWr83
A1KIWaQpdFUE7IQEGKrV2UUfz39bFYtv0ZyblJKKUamPqa1XYcvohjowEfIV
uAN6d/ZCwWFJCgPY8bMdybWkhF+p/tj+bGpcZGjSQt2DLK7hbgThCJ4WFYPL
befS3U+k8a6kvy1OgxtfVWy+CGYI84bODIRi8RVB7OZL5zWNinXbXr9BDTlM
NHygHMQTCfy/H6d84OQx0n80uq4i/p+Hpw2L3XIrgpQ1fAgu4AvwZoCJXbUz
g1RmkgVtoNvRRmXp5l/keyJlUm155LVkPKOU0/w87uu+FAUtdpJFhIsiYC2a
1gEfnxwpJJvZOL0QFaJo/mK8lPkWTKP+DYOinwVbqkwao/u8p9lHXfFGSMA9
FwxTSDVgmzSwRRMbL23GusMyKk3GMh7JCN5uu1AmBQhDNyoQ2qUaXNXmd53U
Aj6tWX3wGY72s7afwOLzB6bhVV9uKskdjD1qOYGRW+PG3llsTiKOG/o8ne8A
itCwW7gn6woD8aWkfr5WHJHuOxy97PtzDM27Pc8N/WbpHZ+SjnAdbfp1/bYY
5feiBVMgRYTRs/Upk+VC2fLqD+mLABzMHyy7Yh9xZcZ1zr1E2qEZJn1ZZt5a
trCCmqXIsuCIcT62dtXLPVWEpDHwspKlwxozsN77o0KE41TLnHoR8kLvCU+j
AlymtnFRlVqqmpdRfVOTJI3dJ3J210B+/JhD/oN0B0iBk8pQ5rd+UkyyT6hR
fAvFyRCDsTnn1stygMzlKUxpIh/aijjtyhE1GyThI/EoxlftA4yYO5tTnDbE
AVNNfNOFnra5j7tJFPimmZhhlUXiZKOy5ImDeie59XOFkpLpl7nyCwXlDVRZ
gfIUQm5fVewxOqoYaIaGy0VdtOlz7jy3D47q1P6mJL1JNim6TXqf+qe1gxaF
+olFN4PJ9jpt1yBa97kC5Nh0hIECaWeMWalo8AEdYc3p0nL385gZ/9+iAsWt
rIgnvhp9EKQGjEsFSHWi0CcxTmCDANcuekgtlYXqN7AtMlS70mnvi/8/cju2
qW4dAY9jKa3tRxAiLus5rwZwum2oyHcNseu4A5iQCBbcWPx2TdSp9KdejBVG
FkaJcvVxLagLlHMf89+ZwFo+DfP4oCeGMB4M5FHgNjUaeJqVVH9sXdqUBxeu
GIawFH95dmM/oOihX/+KdCMs1Ee4tdkAbNQR5RUErEVHBi2TACfydrVWW/6L
DmN/f2TUAYAftB2QpyPYEEaft1svmLNGINsiBSTIncTOXtZTmEJPCrfIbUjq
bu3tQUBwJYBp4prmz0AP6kAbz+1gdQwTeIGri4IQoZaTSniFfYi3NdXNF7Cm
d7So3Iru4hdhZjFnOJU+3sxTNAObIcPgBx/iuCeXz2jhCNij5dFvk7IX2eTO
S9OSpQCuBqjV9ATjmT+KL+EzM4axiahrBmqEv5WsMBDW2HG7MN92N7Uo4dhk
SJ+qoKQdgG7yiWjgkd3AHuPCYoJiJT5pQJufm0eYwbPUbSXbPTD0DkaJv9qH
JRPvVK1oclGA8uPjRXhpfipE0NoCajQ8HzZDN9TUPvLZVrEgAoo/S6hABiTu
2iE1BWW9z9j4fLYO/n/ecpOz1zQ09Pa9ZGbKna50B5xQR4k9iJYDWdhC+RD+
dpplJoc8Sm3WIcIgV7/qh6j84D/kO8viWOHRsIVCv0UYKpmFKJKXjvuO8lAq
QBI3LxoLR7KI5kOocdALgD0g5I53GcRF7KCmr6HPQkg6ceyO8nNup8P9vxvb
7JXTpY4aSvQS737M7WcJI2yIYerGkXPWrS5gmJbJMU02KxxZjQTVWLASzpWR
EZsiR42rVjEjazh8zZMNIqGZ3EahjHc4WsDg3zaSLbiJBJOxykpenaG2Qzp/
mCj4Rf6VJtkfOm0gRrv6wXnIDxf235oED2uuHoCiYPAySvMHXJcdz776EZHQ
4GvnhPmZwGV/AxNUF28sNePhjzc2S0HiWzByPm4U0CPJJ0MOOdjAGXt3R/+u
nwbZ+ZNCSnyyMnH6bNfaPyY9LbpSzjRq8QTxKTxSy135Fiqaqvqk7jn53Bz7
A8qoZO+8/4VeIfMjtx+E8PEsaesBQc2pDbm+7F9aNFCuD9et2phdthqyhHw4
wBKtQWVqKzRIunzItLQDaVNDf2kD25XnZFcCB4YV97cBAKNSIjO8woBbmPpR
7NA3s5we7+zzpDz/PhwrDlPfGV7ZV+/JyfOJISNGUBaaAAqkYzto29Vlab7e
NdfSTNjdP/8n2y0TZisIm+i7GWEgGKaf2EX6dHmYOEugKuWNYifjYKD8NCXC
IbUQP4eEydJ8rJKEqqIl9cTTReCJcU8o8pSoBVHjv9Hv08u2YJV1gafUiD5A
nonBpeu+3RHFfOUWgAQ/ZA5ZDTbJ6DilkxzHNs7lA+9DgNM1OYLXsQS+Ja0H
yhIZOaL1WC4amvEvVmNLJwrgj5GnAEzqI2mOKdjFM7GVFL2zCp/6Yje+yv7w
pSL06Kxlh+i+7JLaJZbNnXnVvc23kligZ6+SGNG9zINCjvQz6/6qMioFIWib
TFgtPhh03VbFjdk2SbVxaq8Lt417vdOagWSnnRxGl3PShR1PnYpfhDVSuZe7
1glVKYDHqDZqYWgLHNSw7+y15/V8YZrCs/nHsQpXO8RmvEc+UMO0ULoIsjJw
4OGA3rrBvVhJyTaf5ko6SQw9vDwbwJypldBGkbekd968ZIDM8cS+GJ9dm0Rb
DoD1lOIrZQej35yojXOThxlk1LS5ZPH1NvE65bvYOXFq77ibKt6HkW/J0+Me
g89Nfz01Syx2Sa9eomf2DYhzHOKbAdft9w6UmsYmiugY9Mxr64p4F7S/cSJo
/tm/un39SjpKDai3PVVPqViR0bBncedqVUb2T1taJS1IE+eU57AMHTlNLFFH
deoBxP4o6yO3mLMqNNNWvka84YGym5cLc07cuNIIQUBpU3vrjSMi5t+yWeJ8
6YLFkCSiqItE/MPaiItMuXWn0gPaSgeV0DVLbc/burQib56s3Tpt/T42xh/+
FzuTI+zIpSeJFaZ1zvz36H/Vops2LJNM1LW/EvRgD4+vBEcklkmYfIjndqlf
xxMIT5M+9x16OBFPr9YKE+xaH7iqbzGfv2wxtRBpHKUl9UASPH17OjZierXw
Z9xIG0jYo8rbzrkNOS2S+7CIIjilyrKbZg3kM7Di6mAc3Ujv41o3oQUiWd5k
I7pHz4I/RmBUSpYAF9Oc+FRz0lJhNEa0AOX0kPDXFJ/tg8bwQzpcS25LFgwN
SodW47KYQbzUM1olxpzxf2Qkz8Je40XMcTnKp9W67eLfvH9q8UuD4ZmARUps
620+wB8Qle3tV++mx/uL2Q6uuOKK/I5EmBW26rR9WwStr8Wz5HLrdTKO2SDk
vqPLj+0eJi9Yx3UiCEPoSawvEf7iktZ9v+u291EU/K8O7JArIMukbepUIraO
/V2S5e6OboZ7VcoBRw4uQZVdkuFZssAYeIytQy1r3eF7qXwSZIzQhKTlamYl
i8nqEfgLSePS8BEWTN2j4uC4dI+FSEftaJdHE/CgUlLVRuOXUD7E8TudmVIo
42E7nGfCd+qilpNnkYydCMS7R9h1SGGWCM4EXetNMefKjXLmhMiTo7k4y2D8
XY2vBPhDRDkivtbkkqCf6pOzebMCy65BxLQHu0kAyUTRrhBGyr0sqjjNY3C3
WrHRdbqY6xnHeUAfq/vKg6Ck1DrzKex8YiCqchjHXvxkNCKBTkLwVy/Eb3TU
ZdWWMQ1hU/L/2jk98B2rbpEoxwWw/EMhnEoymRJ8AYN3QDmkoXIUp/RdtXHL
+pD6WQnWXKhAlQpSFLmEhPECo1AURvyQQXYmSa9OqolcFoV9EdncrFVeKTPP
PZFPzMLZyF1l1UW+lXTLp5EkjxZ6BAP95GsnpJPYCdAftAmwZUyU/xPFgeTj
AH2ypqO7a6By20YP8USvQ3voKSgbTfvRLYGuRuHuNV+61HDhMnmtFbmtixuw
KM4E8yc208SLIKZjEviuIaEL7cCvPKQZhZyRn8MpJAPGi1T/iD3epuJDvlUh
A7Yw6VqZ+kzo5jVBevHzFN5/93ThePfkjBNDMDWfdYaFBSeFe54kvcP0DhBL
uwjlqphcqNvi+2cds6btsq6ykKHDExDgJ9Il8bzLhrIFTHJ+M/IP+Te+6yvV
gFRTFYdI1f5ns9QEQRGqkFmkJhgf1dAr8HQJo8V8+Jg7+69vfffAwW2i+PWc
gLdr4VMLStOzFbRtzqOErvkHuDutjofc55+YOuKKkOE++8m9JiJ0QYm8sFPv
zpr/hzjSkqGmARp1stWlnvyffzofUuW0ynQY9a3GTt9SuvgbL2d7jeHUxWl0
YfnYq9jsywPXMLH2kbkYKiCMJOSyEowjn4tnQTGu29NogtWdiQe+jgeOn7NQ
dv0pRzcKqPj2yg5lee5UyHcGMDLHryiSsPf4dpXKZZVTfl0iULw/DPgtp8uu
9ZNP8Ad1V7Mg9g6sufOS+4fuw1Udel569o2B3Vm6ph5N+GwCOiCGSXK7QDjm
Xs6tBid1e3giyFebo4qlA9euTyuJJcRKx41F1OKSmt8Gbxym5k08PTaAiL/N
+VZwStpwePoOx4Lbcslw3XoifuIRHukSOugJNqDArdiJwvCSONHOU7C/vCSR
39VebbfyfHCUjBsZLGc9nS2OrClj1F+tQ4XfN3kBjRihbX595cgDL1ulibPn
CN7kmgy5Ly4eAvrWQKxeF2l7Acvfo1AziXYE8zYBNxXAKnc03AHcAHfbTPWj
tiLFnMZK+gQTyRwuQdcXYgUuNpuMOBVVbow/boB63nTxV3z4VBWy2nEszHTv
hNUzSUS/sErrQueWLZKxEf3u5KRtL+lhGk17Lai/XnyVLuQlKR96XCn4895B
MJKL9c4RvT8tdMJhy3GxSwFT8aBL3IqGvRKfhDV382fbkbJabbQRU3OmFqur
EosvBZscqAh6y5RiJXv75EUS6sed9s0hRbsHo3v5sjRpggDMV0W3K9yUOmm2
VGPqI4PNCurZG8TUBVbqwRpRHZkMWVttCsYamJNW4dODTlZagxTFJ8On+yWj
4+BEGI/0RqlEgFr7WuPwX7CqqXAncpUY6/jjpcm36qZ72oqGji+uHkVAnVkA
Xo4cM6f8btvfWI8jbcJI22jnz1s448EmCguJLFY7OQBKRRuxRlF1V4n9msHf
mvp5dmoJIXiB9cSQBJb1Z5KDx6RKY0Ep3l8Onn1cvL9/RZjcdKKkMLAXzQam
rfwfY81Ya4FCSKXtPtPrf4JUm8GwQW27KvHHWou+7LayB97LuJVO0pPat8Vk
YDngB9b2tOSeYO3IjyS3Ik7ziZBbr1KZVbcfE1CKRVQ45zDfu0ovvDjrRcpO
uxGcnLVe4y2xLNqmqfB3d8E4TstS5j7AeHQpbDCkpnnnTVmiXckywbuf6jTx
gmPltxcDZFU/Shn1ynHM7+Qo7Fg6DglSCJ2akV1X3hJpqf86KjSUn0WG+DOH
Oj1v183hAux/t3FhZ1RwNp/X0BBixp1ab3PWQ2ah63MJTIbbAQatapYkbHiW
R9h4hNJpVcchBv3+PNSy7xy8U0pBU7POxMvUDb1u4Wg3G/hwwo+PV7sESSbu
KMCB6uauTabhAB0u+XKdhbjfskeiUJ60YQWHEBva8cZC2gJhrpSi347e9E4K
qjEnBRwBCLglYoF0Exlpkz2+YD3ZkSczh8AGvJwm865yOhhyO3/9sLCtDgyo
g4tr5+eGZaxdHknGkYvGuonwXx6Fvs/jLQIa9oOboLBqgX7G5/lADuPgvZEn
jJpXvoKVm4ah+BJudfRJoP83sq1eOjygdye6u4JrNFN/TRCDHQGWu3Bc74uP
WWA17IeeTy1wraqsH1aFvZzGPlsMucYqj+/+GtYGQ2Zh9IfTqOJ2BQmjVBPM
sNa9PEmZvk0tGzaoD3XQTYYZMFu0WJ3xfTWhiZRdGLHe5RL796M1lQRMaGkD
UUEnWkun2gXGrf243ZBdL0iwVTxM5SKarIvZoa8EukUUK9zy4aNA3DfSDXc0
etfU/ktCZcX6ZJ+ScAfMvuh+LgUgmELSm/1pURH4ZWBQdu6zH9BPDnMio7cu
CrArgkyfEthNEP3oar6lMGD4+u8q08guaJFbDirEWa21HnHAs/w9biiXA3d+
iivAQ3A5IXxyQWGACqyCmgxQnRxrbQeaHSeH9cvaeQ8SoWcQcDbT4DQ5by7y
u/x4pZzyIZVHWWu5fcgcxxJC8DeZ58Nr+oLeOlQVjnWFgGeb7hQ4Fjk8HuxG
cEP4K8/D1YngPNzjqQqc5Za15gXyGRXQK6MfBotClRjZrxhrlz3aSTNTuiN/
1cVtw/HrH2IWbHtKN8Ju+aVw+j8oJsIPxMbmCGB1NBRwG6ndP87hqhHRQtnR
PHN56o642/evKMQK2d1dx5Q/adfm3YZY+botW0RBmfCxhm/PIg0gDoNEUVbG
UZ5IPwvJN8RJaTZ6U5USMvtFCg5iEsusLo40VBKsuCOeaqFx3YPSoBclTkmx
3xKeduRYdYWK0n8g60uAEKhneSchaz0evnDJx61khUYdYjWJ5TdPhdzITyE9
9lZV7zkQ6nHR7cyHUunLia6d07ULN+nAAfR1o8b5XzhAI+0ErhkpIVhd5CGO
wVotiI660YEUCM64kzaw4iE9OFqvhmfFtoflsPrzNv4dAR4e53bRYCT9o9eF
Mj6Au903+tXV/mdj4aTJsFrlMv8rVsacqvHCS45n9TvEnFxhQuwJQpTT24Sm
pzHr9DovsCusPWPdNt0hZtMoEx9PpscHZ/sW35K8gjf/+jdLpC9twvi3h44p
KFv5YWoTEKQps5D3Zw0y2AryMMuXJarDGZ6KJAaq+i+lY3AQZdYeexbMXluX
I6uJFpeLyYM1fNdTa8vve2zuUdj3D+gU1Heq++9vvpv2pjyPf/Nfwxb4mvKV
UA4VzHzJNpqeIWH2IKgZ/vBzYx7A2s5l+OPpFtc2KT9JPBSa46J1Je87WjUS
4alKn54CHiVRY2Wo/eikAtbH9G1gVFQqidQPyVwa80MR9KeoPhiYwpsCUxFj
Hbm8o41b0v/TIJi66YhLku7dIYjzuJdq9Hf+gTLbEVx5sVLRXG7YbD2xdXqa
6oD6xqbGIpNUZBnKTKzbGzEqKP8dxGkNsLhWvWBBeSUE+9E1moh/bEMMWo17
3evjk7K9QXjsq7jsfOMiHYg7h58b86+N2o1bn4yLm10HKUXJegyIs457AoGp
PYD1K6D/pM0CE87VXp0Lu3qJuMEs0NwYkzuOamq++kf6ju52MUTv/Wp5xca+
V0ne0EZD4BzDybqkYbYhc1UwcXSiRRGRiks4oCO54qupSElg0n8ehOmpZS1B
z1i0Y663JwtFlBvB9THcV6iRRyntwcPqh+y5SbZIF5x9thp49z3vDtwz5g+u
PUTMKEDUh4GANRIUteWUU5yN6E4/9sMa09TMaIEYbvkjxQfha0ElMA6t9KMb
0u2JlqwrjUGXaH1kttyJTrb6HevR1IObpYsKT0Q3HO/6dlYk8JdYQE3hNt6p
fMHFMJluPiC1w0qERIJ1tT4FOnG0TxxXuS7AQZcyygahRgKmjsswr7q3ghY6
XMVQuUDXz7bnqZ4NVCA0lWEch3nU7QZ8m74BxxQ/lEBr1wRru0QAE8hx5sjK
CFaJdw3z/RWcEXxqwa+ztYgWuiFj40adMlLhivpBtim3f7ZM0XDxb6NFwDWS
Qq+eH52AUh6Fx49FTtBK1E/Bd2ZX40FA6zB8M9muMIAnlVHqjoaypSCco6dH
zu0h4s9yjeSHU+6OqtVOgC0C/QvZ1ueYWrSMu9lGsKn07tVfB4dVsjmi6EQn
drJEz+9ZtoZYuXdJ46ADVWfvfhE4Nzv7ZvouwN5njEqYd0g/kNm9HunUih54
X3uWXx22tK7ELSsCLEEi/pmGMjK1MNNkOZIx/91FNdcHxiZaPK7lGYx+tkID
plcCvQcEB+9lafdl+iWrnLphPCgRjkQ3aOz6IObsiI8DO9GU+xOkbPuns7qW
PQx+93QBpr325gdm/3QXPAa7NAnoP+KI2Ms1pEzgDdN3oPANYdvMT7e2c4tR
pwFolVC088TBMad/B+MNUnD0iXf5syPu7T0/ftqtJlGuaTqhNeGakdxswjmF
AmjmOz9iEy+MOXS6ezRaSmGM7lZldsSPAKQgqa0X+AM6J6ASbmmGZjSGVMR7
k89DDYwqxg9acBVYh/vrDla6OIouygRIzF1x9i5BrFhL2USBl2bwpuFdUfI+
e+GVmL3yYTC8v97oCBXnzh3H5Fko6jgSEYJhPa20fg8rxgpkxaaY+ttSxJqy
EwtsM+6aZFUNyXrrbF9ZL0hUNy2KjdpTZ568jUSZxWRXv0a9kkftQcD+2a1f
kQP5TCc610Yw1A5vqL30Q840v5+WajhFzjdn1Vh8ZgCp6KX2I+FUoEeCmHXk
6oSzr1qboZa0oC2viM/TlkoF407vomSgLkH14zs7Gls7yAr+pSjkBw1IgFja
9nMOdsd99xg5x4sLExrAf/D/BoCNW36eErOnz2rP5jq4cvQ2dTyyirng9SfI
or+h1GXdFHx3vLiKE8Qbpklw1CSf+eqtGXWMDC/y5zuE0wHTFA7gXF8P3YhD
9bvODF6webXaBnNl6qrIeVUFRM42Ga2NrCvK7NXYkTr81GFRKmLvYODNiVMG
l68XtlFjeT4LwMqHIpUzia3EnaJ5B1025kGzdWxqtmn7x1WfV3nGDWxoMmsG
CFnfESjq1IAfJQQ8aACOvFHf4wc1HgWGFjTqEgV5q5Iuv+hga23YRbwkXChd
Vudz2VWjBrwz/pb9VEQbuM33fU8rwRv/PLiMJp86nbrDWqyz15tA9GveF0u0
eqSnN7OO9x2iVRbo0TJtz5PsdmcnZXr2vDKS1/U3sjf3R/FhZfYSSRzIyUSW
thkeGXQbPatN/NuEIvWzQNH2sF9ryt/3fHNRZU7fscakr3NdRp/oxLifL9vk
nMMdAtfPvHlM8BFR5Z2B7HqXRF/q7pAlSGJPzSFumJeuQvqexGlxEV368Ygf
B6pfFAZpRp77D+MzF+2ueOGaJjw7CMWdXYl0vILdHa10CVePb49FmsvPGkXc
JqTtMtgxAboAdDqIq/OqNI09dChtjyuKwtc5rLFzjGi2CnB4izJeMziT+5h7
VviG94IXfqSear84ht+Di1aSMVSPecELFFOJozXSLMrzDQYRylrVqRQvLEQO
i4esed6SwfI+g/fRKsOByeYI8VBC51wmNpLdv4joEHHDwGvOHCP+KuzzPvq5
+md2L+vuVYI46sqOwSgY6en3Zh19vU+HvLZlusUy+btxCtWTDENogt+fkCzc
ndNzHsjVOJIXZ0SDyQbbriLB6QmTVEjArFGkubdNahFGdH9YtM1R4lbd1TGt
hiW8owFSEPXH/4H5eTJjDks5Xeikr9fE+peuoTxHC60fgFm414vhoIBNKq4b
zxjMn96YWTM8yNWPPt8vMtNrCMdeSzWdVz0uU4KAF5YgGOGYCQN5ZJF74Z3W
Q1OcPZbjS1YmxtcpjcjwAwooJHU9eC5ELD3AqERtj7kWlNt65hMbccJbWScg
CE2woHzM+Casoynne565rNYESVN2bGA/ktpViY7vPmPC+HFcoQhxMeUiIDrn
OrV7uzB3lBJGUyOqxIJmOn8m93bmxKCFkfITXCqG0bFr1rBDb5tm9TrIjUkb
OyE/UIjGPcDPy827oUOT0LqVvtNX6vbgjBxAt9ExQxAVX4/ozHmad490ASJE
uWA8UEZnOTCd21BZyaL4PhZ8L8ARdKtIbW5Ny9GoV32mJ2P+jcX7Dwit4PU3
agjwsEzEbMg78V0Q+EL9PHGeZM744CymCk5euS3ViZGllXDkSRaX0ax4C6/K
AwkwzxMHHdVbaSVvJMjcTpGeb+OG1/HSgt3O81iRSMun3c9TTt+uflOJ1onB
GrwnK/CmpTGaEf4iu+doWQ4di61kwXaeaVzObwtV7PZtxu0H/HQIo0w1cVbG
u0yxXARJSPd1oOhnIAM5ManTX0KAmG17SA3z+JA4y++1/FEUDpXZIHBFZWxo
C3F4BDSBEFSOmchi7edSShFC0I7BfIqV6g/3Ekd4frquCo/JS3ViulmcxGtK
9bnIjweqMiVhrAC2wsq/qkmvfE8NFy+0fa+9uA4vlpgURtUECgG9cfEUj6TP
5bJ5cjzF76F8C7bAmsc3Tt//xUoTrxhopSIVYdCq4gSZ+jWl4oX5e1e8VWmN
grFaD5kre1cEeyPEAi6rZe0dILPI3KrbY3ijJWwhL/k1IbhjDv6QAyDon0ZG
zUwvXn2PTIcTCpluo6fb77iRMqAcogrQ5MdyP0HCzM6yGXjPRf0YQSOiX5Sn
VFbFaY4zJGozsMMhRIXdwDEu1JnabdcBX7u0JYlvDJjO4u33iRpRhscQz7dH
QR7bh2MG5bKp/wZAHaiCivzlhlObonAtiSGxBld+/bB7seLIK2RmPb+GLXEI
SGNUvZJeKC0P8z/Rr9JkkEP6T4y/kJl5vyg4IBJ9OzQgyYFzfwZ9Gug6Y5/Y
LC4YV7ctcsT/FXJy1TXTSqFITL04qEatYngRut9gMdFLjVoO0ZBYIUykGcWG
iCeZTanChGi1ZmoNnks84n+mU08JdKRy2L6equPTBbLEhHApU6b1OpH+WN9x
NEZ/Fn7uwRvAaGBMZoifiYk0LaHqtkXwYz4o2B9ltKn6YhckdAIKfv4h7SAi
vZWxkqGOXQFZG0Dcyw0TT5Y/mEUL1ioXV+0pBHwh4ypCPIbYTkerN7q0at1w
X/yiLNI4JpQwO0R02Raw8DVGRe7J9OJECTnqKv/8VHw0dNy+sSUm6YaMML1b
UJkz35TlCzrk/ldDsbLQa0c/u9xMqSb+wId4CYqGnYNU0dSUMP6KK4x37F12
FPkPw9sZOD58fr0g1BtFqXQD6jlBI3FUXDTTAokb54dDmcHfZSAratJSxW0m
chrd480m4Xa4msR8pct6HsZ1jgrFFxbW9w603+TRNACyZhz0j8j78bgvn4Ep
G0ESRmkCx8qGg4dJu3ofevhOvFMq9SsjkUj1WImds+H7Cn9iUV+h1h2Dy7Ea
y70M9sW9Xo8AGxGnvsA+7d5xTDtjBujGiqPc1ucamW7anX1jLsVgqX/IN19O
OFtkH08WtFsXgp9rDOHXe+nC9syYSaEo5CEUGU2fQ02xUw+O7jeBPQO/PfUW
Dg0n5h7v9ZLvDkmROdErZSdpcTQbKeazx6r95NfA7a+IKDq9ak8rackUyEAX
bRGcy2+5fveIE9DdVlgZGnp4TM799hJLslOyJi6vfoZ3xPwbFZ4QpFXeTA7h
GGsdTu/6zQUcyH5XdgnK0DeXkUtN7X/elsATwdZdud6wzEo7ePGjnUZOUoRn
OX1WU2Mk+JnN+vVqElRoDkGrUjqV/VQr4nv5Q7SFiieIQF90K9EG9uB3am8j
p5HcT6fzRqGqdzBG1Co5IFAnljr/D6CoiN+QiHxHgMeeVi08kx/X1HHXf7SQ
Fdp3hCWHmmBmTpcp3oVKDPn1BHxzEdyzUzad3Fz5p8J3GgQw2H+lmN7+D/OR
7ILxfoCInlHFtgBangFC+6/Wgt9Qg3bj+RlZWBB6v/wDFufOFkLA/eQOX8RF
ieX/Jird509rh/ZUs6pNcbPRVZpa/PgcfPhlG/FNtjcv7qYY4mCupKAdERc/
TgE40yixQo98WRy8c5FYoS031/BdsNQyfKV/VpQbIP1ze4YsTI0BzkCwB2/O
wPLJJJ+Lg8I6kLtxofmOBlh8PIaXydRqAQTfqO1lzl2lF2laKc2CtUqFaZ4t
tWoKCbIfZptcm6tlWjzdVuMFwkWa0ayfP+K/mQDwUXuhU6i+PGULVXtKkIqR
2weiMQPqRMIJy6I5fmOfdjd/rJTfdk17EYVSaCbwarx4VORzAuZWpmk7lyEv
Mnod7x/2jqMxPA1TaTm0F5GNEzYUkLGACqvOdgf4Z66zvudRXmqZUzWN0KZF
NnqdAsXHUH7xIfCmpLQMCluy+mCG9tkKgAfsUD5p18gcyid4gyqLDgUJJdjF
WQBzNERzH3LiHrOjmSx16E4R+u2uEybH1tyd667jit/eTkmHfOSAMoTa7vBa
ISx51Zl074HNznRds8MJuKwFA05Z2HNWFODq+Zxbfa7y2qlVHCUkitBjBUJo
kSxCMR0N6x6j/K5j8yWC4R5JLT8AhcoKDO5NxjfsvY5iimBWikvgm8oitKBd
g67seKptQ0Ngy/bMfbtQtlW5ObvWJalZhpLpadh0ksDuzju5LbcXM+1TmnJR
wx1/EFo2DnM/JnbnzGEeHsXxSou9/m8aPwlsHy9ZZepyTUaeYujwDAnQmg/Y
onkEscrLKedEkQt5wuR5IPSyesbmYpUXzBrOUG6+CWCeEp9JqTo+sqkMWsr5
NqWojO4g/RX2umEmZEWhcjN1HFHGZKneZild3cxcXBWNRlYUdqPD5BM88t+6
tG/2vwA8FReoaXO1F1SXPxDndp5k6sm+YGT9c+A0t1EXZYF9NbF1JTrVSSRs
YpzKfAusWvvnaPLetc+585bkEhAHXxZaz5/TTg+HJApq5tVeJL5yxCcbpXC6
7VTQ7UGSLy265yuFWKHDImLs5hjMo+nd4X/cnJityJvo2DX4W9b4FGtKo1BX
Twg+8lAnYcldspoRkWgLks9AS0A8hbLqWkZYU1a5faQGhfz/n/CQH45GzrcG
UOitUMAWPZxoPZ3mli59zXAwwkdlMYeiuegjddm0KgmeqG14Bc2av9LLdMY1
+R77vjvyQQ12kMgR6h4JZqIAitseB+uO9McOVtW7cl6Fw0GGQJTqwai5htco
AmW/INzSnJZtl0sZpyXewYloiMhXqj7tM+yM6SpzCO62N0x6MG/X40wZXacS
GGlTk9RH3Nwu10ufwmE4LX7CeiQVJMzR60dESDW5JsMeoln3DnY3qfEpbU1z
ar89wKvpsyJ3io4vGs0cfY1f+o9xqfvgsyRwDYjVBSjrWi8V6Ib1moaFqcz3
ZJPnzK8tr3jioi9DAMp/Mm2S7Cy+ZEfohaReTOqGG49wpZhbwfJ7XWpUwHlX
a46YJY4QaBGYAFgKYQZgfjQtPotdOEsjcmJ3AU0fr1WD3lUZWE272kbM6rtr
8ZhyD/YjuCwmrpXUhY8zvq16Ww2jBeHMIlQJW2H0g65pDt5rViN48V5R7/KW
qL0wrWqs9zUX8MquKzz/aalXAr+Rbui7uzXMxUlcRrldr9eagjqtKFMbYR0F
odHEhpvntmKHOYlwqfz/NwIS6E+3vqCH4XOvHjqf5aDd0S/5YWROYtNtI/lY
qslvQguzQBRuWa/sFRtlJEPaVIgZ98zjsikk7j+1J29/uzOpxGCE6A//NsRJ
IdonaH1JMtiiTwe+qCorOTO7s5xmRtlOhZtAbplwaj6NQI2hghmM5ZbwIoDV
eOclQmEOvd5Cg8Hw38OrmSpVsNNK7FWBXfBbCRtot3Fj8nFy1b6Z0GlTkGcA
yjmQjTCWAdelriWbFmbgoo3O5PCdU2JPbe9/VoVg0H71PebY1Koqkt7+ekQE
AFrBslYJ6hVq2nUktHXyp3FvebyalgBUz6b/KrKAcXwjL2xpBtUraKH5mqEQ
jNlF2gkwZ+AUq+o+x12nArHFc9lmbVsTxNXdDsBAy+hOTKbV/gHLoxPKG8Xr
ogtcSfLugS8P9WNGrnCRJ6jWv8Qx/V8Si5zFz4ZB4xUeiOv6fHSFDDi2B7Wh
w5Vzg2Sbs6w7X+btGZhnmInBII6JgsiMWjcEllhV20TqK5T3fWJr5wTiIPQt
sKqpikLI/KIELFZbsmQ5Xhir2EAqirrScvXwd/NR7ySxqKUc/UfnmbP55KtF
b5Avc7FfUcQLqUztciO8206XShPflbc7xIL3w+GgJnQdTOxygfXO4fs58xmT
2ktS2UvpkS1nIIcderTZYBGVY2/t9Eb/A1BGG+W5tRvL7urbqj6ulQL/cEwG
3lC7h4G1CN6JIZUHCkFhvsveEGQ5aKP6x4X2QYW77wNzg1ayKeGw00LJqznA
pM/27Ste8/ZfUMZYeC99noJ8BElU56NQhqg3dqcng6EiYgUJ+AxJB6KKXy8n
CwiXH5KquzqkWJ/FsfGvFf2mt4GoDpOkcfdORa8PV29N6QAYjBEk3BUNI6Uu
EPHxATKLqotd8R2V3k+hXEj0R0Rrgljj42Gx9HOqIlSOpwCDFvmCR6mkuAOG
64N5mInYtFRPX5N8pmyloFlZeYzyknX/ZzzU7SkK0BpMmhXPAFodanyrbRiD
1fMrksfq9Vk2ryoS6I6CVLQ5ogGKAkbOD1FceiHHwPLZvnr3Mz3Dhy02DpJe
WbWO8Nfjn29XW45qj7zY8ZsM2ONnu+Bq7RzWqiCKmJ8npheCmE6JUdWWel2j
l5gc13Jz34vzKwRYbRDlxO1iDpH8SEJJRG3ISyJiavxpIiD2RAUNvI9uN4z0
mcLlESURvGGTWPD3V2SqslsHPtuTgZTPkg37JilohZ4LQepyqXca3xNcUXi3
7K+PZmoKjLlBF/bSNx9AJgTHUx8JQkZJPjUc3wE9gIBFiVfNsTLdOWZqsvw7
CMTdou6JAevag8GYs4xllBRTg/R1eaAbcNIX40JLm6BiTFxDKF0sqozTlgmW
RNGAuGYw/xqJJKXS2j33IhQbpIN1E7vH9kkPgELhW7eLXLdhClNpo5BZLLzE
C+UfiY12sgXU3y1aOuxeJi9sukgUPbcJr36aY+R+Qm+VarCuPGefnp4bwCE7
W/VkyKw23KPkMHTev9dVppEijYkyzRgZzVzu4MrFseWDlPhnB/6MnJHZtZdl
YHsW/E9FAFQc04BMmyuTRMmwn2ZpEWQllWp/ndaAV2//A7n1PJBLoucpEMdi
v6HANE/2Zu68rQ+FMYVHmu1y3pxVzXl/Jdnz8lMY8CQniaFYKluMM2MoPZ53
7JBhbtGRs7MHRe6nHvpWuzGEgFrq4HC5pL4OIvmHYBJygE6ETyjvdCgNS489
O1j4eEImRtF8++JPz3NYsHSd2mQ50s8jqkDsdy11UGIbKUtc6S/RqtwGqvtA
oILT8k4en9OYeinhpMuxyDQVhYkBJ1Ri1BQIX4IeUpeMwxzsLVvdrGoeW9/z
7hZbUY7H8FO60yoHoIjunh2bBUHxXHqmBR5f6fDD5ZZ3DZpWixGwwZh5a4Xn
Yx2hZXvq09qcvm3yuJEoYTI3nnAuBhwwTM4zzQPoDZPgTz1i8nFwXOac5YqQ
Y4GyP249ogi28UGl3gr2qdHYekFng8Qh8qsRjDP0UC/olj+7RKNHjDiJkbsV
3mXw07Bqf3F6pk9OBq0FZNMCSYTmGyIREr0e80WIh2wtxjgA5D1DBdJiKmuG
K+fQQy4+6CxvUCjTsZzcrVkl+pcanXllfxtHN/KgQYgqFtpION9ScYIx4+S+
+wQPxJlLx0Ow5uuU10y1UOMBWbjIYXo4pmXYnhGTc1m1TUmw9LWawlrWL6Jd
JXQiO+d7z4GvPPRtrO5oNmKD7AWpKysztEvLBWyu1+3DBvht4+jkRolYNWPD
JXn+Jo8Ww5w7QE50dGweEAn2qaJY2aj4d/Xfu4z6Fm5YwrSUSBX16+K38+1G
rBFAjnzFD5zIYMVza67W7h0pZzdAGlw/0RU+bbnJoOi64LwB56ePlbU4dVAV
al1InXnTtOoeQBtJUqdsGBL17pw6qshIGdvzpzcgmvwYOE1WgVsBwFh0PPxO
8pmFCz6JWtqShpMO1ixYt8MdT6lJoTgwM/yS18DhQcwcC4Xqt6iWVxuqeEPh
gYTX2GGv05KIq8+TdbShmpr+BLw6qpxS3hr9z4z2XmtPdxEYDruy+GDVl/hW
dE5Z1VgxLn0YfYMgtHj+gpwqY6hX+SlHWVjEslusGGQhvc1vjUfqGP5EEC0P
LP2Qm6ZPdcRZkwHY5MnHQwc3VrMrTJt4mI7E5nPJG8ydSweI3et4jCD/yBNX
YHE+dSxQlhSw0by0jgW2X1DskszfC9VvWPLJ7lvUmXM7hMa7W1aYmrK8qXRN
BdWqVdtqR0uP4VCuHhmJdXsSlhSU51quX60Wp8bHDN/D+3q870zHqISRINuk
ax3sQzm/KrDOc9rqs7ImkPuvcMJTOJ3RkG+4iOl//+Zq49Yf7I0gafbUzXDL
JH2AH8SrvE0xKVvBSsyiLvo+KuJIwKDzh3zp7LiPDX2tJ4d/fQoNQh5qfZuH
M41BPYkboP0kSN6T7JlR04pIL/JApOCzX/HktTpkiPpTqmIVE8CQkkdnedMA
EHgT0P/3CbHoRyy+qUD8RwqT+hpdkA7bfyCUUklGIspuzp+qEl8E6kn8Vg0v
9j2re8O6h8RLhi1TbFSmB6OKr7Vo+RGidz5JLoTW041dYld5nLtyg6N10bgd
hPd+klVe3l+5G5H6JprjV3hoavxuTQ+u/zbt1V4yG5wz8vfDlabbd3B4GeJR
Hcm3Mn95cbgoo6GOwMBCi8zNmoXMCtiVj7SuPl7lADYZsWt89wBjg7HVUtps
KUXR8OGqt/XWGlcmtU2icYOHKG/5aUoPdNgrg1loYqJDvuqmXHwBpzsRa4x4
Af85yEAkGardUpRNUYt7xQMW3jYsCkz9q5i6hYGKtEf/M83zrVDW5AFSyz/t
9GyNfAE+MjyBz5jHVsWxGe4Xd8DDNBwbFxp5+Jbgr5mQ6bZFPBgxigsgfPjg
0LXAxFSVpweJ0Wl0IGlGJ2jCtw36rPPHvkxgrLMdHHI+3u990FGOSa82tVl1
N/673ocz2oX6RTKeO0YB0Zn1DNF4fJmBRyt7ArIcQalEU/RtZtJLdqJ92EYe
kxsMOdhzFFtk+omHX9/lDT92lkxM14O92YGTJCwpwq9PY6xKD25Wepu5+4cN
eqNNDi3tbD9L9I+RxDn/Ge+6bSgEu8WuFClXwQ1NNXIK3vazUlUmKnHJoY2t
3oqXgfiEtoD1xhLVd132cG9rBOUl/V0KleDIU51A4zbJ0Zg/2DUpMx0k3QaA
Da3luoPuT/J60uOyjvW+kyuZnrQqAMYLaEl7+NxOEbmujfsDLMWIzrkhyIes
yXZPRqGNcDcWRc+yyKF1Kq0PmS5Q6Qj68IggqtN9IFhbwNRO9VaBL5ZxU/no
9n6W8ZXJuSXSfcFySkxPsfdPgUp52A8MLnxXMUuASr2m837S6EyrrSa9FLdh
06RK8mjQqAe60i6Y6SHQsln/OTx68W9EK8YcB8j9G8e0mONvhOFxBfdAMHJD
ybIwswdSx6HulV7DiMHB/BB4T1PVWpmRklVAsxR3APq3eygZmzfkjL0IvIvS
kKc7JGARJs7k3Z+ynRK6D0OoJry3CXmxR7QybV9gq0m6FP1V2ZfF2c39b3I/
WBjaX5POTB/YksTGJDiJ+wF7sEqNwq9Hs7oOrdtuPFJ5228I4bnqAzEsH7fc
0XJ+aw+Wi9u36JwtgNIXKRuWl3BH7iLvUVza7lsk4RwITJN4YJ+SKmNSPeIm
aLgrN8MwkiLGFYtuSVDVQhvmLywAYf9cTV6hI5I1shT9MFn3z1jxCY6aoukA
7PaF6Gzu3g087w37aynZ8ISmWcEHt2B+EeRTnIbDN7K3pLdP+45qI+GAwoPI
r/y2AjZ9zNwZYV028OMgyD2jCOKkM59y5Xk2ETPpbriV7QB/0P1zJdox3cSo
4MXbGjVipXK1xQ5ps47SR/2C3DYuzxvu3viQcRcs9e2QGI1VktHtmXs2t/wk
zPHK3gdkivil5SDYyuPBpmGNNGpJYP53vfJ8Hcq9JbtIkbA8ofSXFGBwMijJ
W5ZXV6soDBAmgTqaOLZf1zwnDlhdBWfJ5/X5Ss6/eWv/wi4hN0JyuS2AtEbp
7vHx983RP+18nBYQ5pT0iyXQi9hiMyWgqdcGZxrCoMkWDpnSOclBknsokot+
ee6ljbUF09c0wJLurkjZxcYm73UCgftcpFWIuhnlSgJbxTmvqAnTkumIenM/
+ry8B6BYORiln7IXKODlZALQr/5qR+slNFdJ2wfIdzDKe06G+5RTz6tOwhHi
amX+Ka9tfSKgSRTJK3blxLcw06/RBw1YP4+iNR8d9SUSbI/BNKEMV+aC51my
sAlNinn6V69FaNoilhcFVBqrerP9O2CIy8ZkrrZAtc8TnHUnhbBrehSTOV1c
y6j01ejDcKHUlIXdoMNxLK+x4cRWQasKeExwyyIgNFiIyV8ALFfuXIGnk4A3
qodpWb+UIOdIdrhjysGgBEQkPS/waHYIApzHGbYg5yt024/0c4sRnyPGE8HM
AvmoL53lIIY3HWRUFfk/wyVEdcu4FOcgDFbN7W6nnfq3cbrXJsQZzUEJnMR/
CDkfxD41q6XiMjOIUHREF8mJxGSlbctTaRMtlgq0CwouoFM4h9alTqvMPe6H
G1c1VyscWtS4Ize0SBKVfvpuODqEYeTe/qdgoc7dWX4TOdSptesJ9gSOkFaD
5jSVk5NmZbBZ9feN55Y3z2q5wO5rCG26d1Zl9zWBhwYXr0J5wgd59MeAPU5i
VfxgbDbkrvKTfv5mDunWjSuN8UnRLZkqXbpTSg5z3U/drC54Ww71QWU1nlp8
e3wHeslch9adJTFZwPiZlLjilO3NeJHnSntqL3j3hSplWX7brSqKBQGKh+S1
/G3aD+11t5/L3VHF1R8Tt0QIjimGZdhQK1mAL7GLAOE/UWu5pE3yCHLgA3zh
mMQDV+0nTd8s3A79jfig2lhs5K08eBb6psl1LOsH7G2Ev7CxzOqLZG2730X8
twkpZfij4dXiJBjMzet+cy41ZrdDw2bsxq+Z4Knf8Gzz/0rIIqUioCfeiLfo
FHwN+Jzvz3jPt/X73dDufksz2iEc/9g5VltOpBMgio0HLBG/oBwQBtOCJolE
PZXL3CvkWYnCXLPekvMJ0HeSu4hkfvrcBlVRuDx02LuLbqI5Q2x9CvHsPlb9
5XW+lsIO3U8rqQvHOkjiTg8nrWWKcGIuOgEvh1M37gAeP6MniYb19bIy+z/a
uByysEPvorsT2hNWNa1omJ8gDX6j8ibYvcr8J3A4UKLlKLiUQ8fQS4ZfXV87
g8AzsS9K4b2nCD8gCXC4z08rAfihzm2TrOaOKuxQS22Zy+7HMdgjlsbABx5I
NgW36qx/xE/ToQ1tQK/hJAMHq5PThw096gDWZS7V7Sg1VGa6xxf2AHPhdHBf
rh7LNdzk9SODzUDUaZwgctXRNpgqp/Ws/qvgeXTvYm3uxfS3ptA+7+dlBJDA
zzZuNvgjj8tjvhEsjn6Da6AnQgYsk8naA2MgCGheJ+BUbdQjKBDpG+wFLhcC
i5GxcSiJQYWkjT4ph4qEFxv52A5TJLguSSIu22CTHyHQALFgsN6SLUDM/Axr
kiA9Mu0301X20o2D4pZnzVTqP0HqrKRVXrPqO5gw/k/aoFyGcIZnsuQ3qIDJ
kkoW2I1wTiNDNaZ2Z82/aSx/CgDosNKVj9v2QZ5To8bHflTsBMjcBYUNwzvj
QD3u2LvZzEddZXj03WcSvEn5vWC6GkjYay2zLduLOQwv3+MlvP+WOsWfK+mf
wOqhh64KMgAne7JjIuyHn/wqkMlmSIdBS8wTCGXDK+GodIJFuKq+BECADtDi
BtBFf2SPsf68KpD0AixLwk2p9OXlgA/tXTF9eNu/NXawwkLQyb25sMYJGhZP
kF4ZYnxzkSuf15mNMG3zn9x8QYoowAFipW6TUhdGQ+FLheTj8RwswDtmRc1h
j1Bt8cyWld2p7FGFJ2W5y2U0NaJO9snAgte9iqc7FhR38pnV8YjebkFYn0UQ
VSU0EFWE4CnUK8d5VR7Fs0wlUGznfibGKxTzQZSPsuUkam4iY3HCaMImMpy/
1ULy02b3jTSj2jMPfUowbogpTvsxHYmGX54lY0xzRBMVGNLugZnTGUcPcYo2
ehHZLDzr6EBDL2l9c0e/jXIpOe9i8ss86eEpuaZ4Nn/qBHePCBtbbHp/OoVp
IBgevyhUclnSOjEU8yF1pUf8i9ABttBRj626jGLMTnCNZxlZrNw+6JRWjArB
iX5OP3asR+YIVIEqC07ErDqfC0TYNkG1wj/vuy2g5+GSWe7oWeaoRaQQw93c
SFtKGS6H7Wd3GBuTuiHWU2r0c81lJR1XVU43dI7JRUw+uB+/m8lHqQWSEdkB
Gg8RePwxo2Ix2FzbSwO60ZK5BrNv/bAW87tVoGWFX2XH6PxpEcPjbr8oiVCA
xwj5JnnweGfMUHMdlpP2mQQ/wISm7ZdJEbvZPbvmCkV3xxdoAA/D7cti9yOm
QbASCKH/xwN4WT3LnQtsxOzNluk0FrN+5kSkuO4yxCKnsg3on/h/+Uue0+/+
zMgFUVcR0yoY9x/1rw2+txrwYpcAvownfO1+8DUlty1+N2mAUkDZhcy/mb2j
4m+NjnodMu6YMjAQ4aFh1SbFIr/sVlK/IwcUOvOad4PdhzG13gpTCOi4ilZZ
XUajmB+8gBqoXMxV7JX/W8z4GMCqr6MgpHPEpM/AwaUkcJckOW6iTVxP7kRD
QcGk1M2xlJK9OtPrW9Fxm2GzS+OthA4idmaUrqKf313WxYgYo9Q594ict+Q+
yiXnTkG7GNb2Uc005C4BO0XyMWjYIobCyKaFaMPcj6/K3Dr6LFsfTNdRR0nt
kz88SbLCpfpuDiSbrASQwg28w18oIxRw/NNZfNR2QBkjOkBzSkF03a75BXbs
lYQboVYBtUNAs6PlFW+lBkcJvm0q5b8QrHegXGaL8YfZquyGFF4+sPU4l9IA
eTjj5GEO6RkhEF8DJiobHqIG1Xu0WvvJNau06ZQLDpJBWcOsQptNG4QxBhRQ
vfVyA/Gw4JEQH0bLfMpRw+eq85qZQbo4tWtQAc72ueRS6CF3ss3COOmUeq90
25GQP36X8HzRQn/GDjVgzNMA+kA5EuizgvFYj1zU+zNQMTNYE5gNet7hsCMq
5ZqYaENsT1S8YLBrAGNBUGbiGQgMXhOOTukSvoHWMmnPY+kC90N9MBpkpq+P
qRm9tvBiIuFbV6/AGcF1kUt0/3bONvVGWuTzoJcLxxRKWCH9do+gd4NSg8l+
oXnWJeQMheLPYqEvcCt/dSP573yztc6U40/ymz1PNHuv9Y3Jt5tzH3Uxoige
IpkflfDD9sVE0HFvrfn43iAuK3UYsApxBiX5/zTdJYEIQbbWKkN37qBtabbX
TwqRKnhOC4QAOaNTGZssbO6WR+cjTjNyJWGVSCB3RbXt1PNChxnDLpedg715
WLAu3BSTi+yQncslKB+9/KiPdo+wcV+4gGtVLjWFmkXFM22fLSKzLpEaW4E9
7Gygru4cXezSgsWwcYclJWm/BSuIvhXIqDs2iuWFhbsKiqPeVgZIF216YT+r
jWoAa2gXfbQjaAYisfo4JwKutpn8Aj96LgCfNeSvIcijQR1zMtDA/B1u1ULo
PY8TGqRymMsJ3HzDfRs88GBfJoM6jrZfF67Ezr0zD9LJfZcRzyQP3TXL2PwM
OP3Lwc3T6fjhYJIsN761P7naEFoBZqdXJlAgFIcAZdFCtB1MJjn4L0pdvTnr
MbIBP1YHDWVr6IsK8H7H91mZm8yJNR9uC8yXvmYw3FslH+gH9bHOLQv9hok9
fc+vCSDWIbN1MIqa7Tx60RGHPc4KyNZDU6b+FquV1ZYoA1ETNmuwUZLFZ9/Y
TaHGVKreDEa4UsFaz3mLW1cUkFLFPkNEb81zxwrwWIgg605S1SPgVfpDkKek
5+Q/V6ksEtnlE2GlIBHRIe+HuYCWxIaRQo4ArI7o9cWvtsSnGucsQgVcLYfy
T3ewOzvo3dM+PxR6w2YGy0VjQOBCgjMtluyoxkk+ebIO2I076jEnt6y8zb/M
01DuWkR/6dpjgNLcuA+feZA6pYWreL9JGqLQYyjfiTEdklJkqsJzS+8iK1u7
USuixf6fiRpCDhy9zevOWc+DyfksGkofiH1h5bC/6Is3i7eCMtTyb47Bo99G
bQEJkVp84V6ox6mD/3F6ck/uHmU729OP08l7wV4DPHM2jy3Gjv2OC4gQYvhW
HUOF1vBYranf15OcIbO0IISZY9TztUD9gmnX250B7Jes2ox0s4tzv4pz1iY+
h1ndB3QsYAJ6/6U1LlIF4Scw+qRbbBd2fr9hVNZ+WIr6E4lp95P2V5z0wXhS
3pt/8SvcSWPpTdYCpcFnd1LyMlhPdUWPxdCYaRgcSdpSkpxyc3PjqYS4V0Rw
Elnb2pGa9TIW/A8CCenF70QEmSLuwAMa3lVTdqeu+XMGw6yx0JcKc+hOrMRo
GRRu43ulwe+sSR1M1JbKfPAFLGRhlZMkBUevnUBqhvaDttXdliunzQT4sy6P
q8gTP22xbnYSpD3z36VdIOLJkeiks1/J7vIYKue25f+yQgQMQPFMugVWgXjO
W/dswGIt1/HART5kgHtncdriypdcmv+oeyVfjS3IHWAWCP50Zytq0DUg2lI1
wYBgEbLR83jt9zEaK3YdAiH8B+jyqRJ1qt+Ac/Lp5hYClKu2h5tBdce2NbQG
LEvrXm9Wk0SGRrU+ezXoyHRxTI063zqRsbjeA8Jihr/D4NHGopdjrm/zy/ov
Ai69ipeUjDOLex+zjB6mhq2Rgb+bFZ5r6LVycSjDy3Tx8v0RHm48p8ZNQPMX
6vRKweYf+K4MGaxJdnRuVsevvHzeuTaMzFjBMFvBwmkYi7zp0/YPgZc3WhM2
netih8ATuv4vwKa+t/t+StvSFxVywYKhKsQ8/cu0ILUUkg2ks2kGzI8C4I6x
2nKp5yiz/VmQQL2BNug5hqywdPECUUdVJktLt+/TgvpKQRBrn3ismycNj4gk
HPpXuWQjptIBdvAFe4SSC9/1hUv7Fq9pB/SApliU/KZ5UmJuYoS3677Q+2f7
tp+ZVmiDtved+Wq3tB24LeS91FS4IBcjv0CR9lFVVZ5tS7ZPX8/DXwrwPSxF
lAz322q7UcKryRzNRmYJ5zx1401I1Z3WOTKnkOkQUHPCU15i7peaJrZO6CAg
TVVVdd5yPFY1ICW+tffhq23hJDnkkW0omhtlvfXDJLTcr2Dr7iDSrzmEF1Mc
H/Rus3WkHKXwMyRuu44hdlBCcYh2OoBRBRRZD1W6hl+OvYjGQzfW3L4qfhX1
DJVWsfyF96r4+qn8VtT+3JBb/p+okiIoGG/xoOL+DRLGo4w4dHMi2vH+BDYg
DpvLAwmgXPXpRTk1ynu5S7R7DrxHvTklc4wBJX1SxqEKz2bryG8rQ8fYt04/
gxRMWQPNY4QOYHDAL1s1QunX2zzSvznvE1LsIJNhgTFEKHup0k6yqxTtzybp
RJot8LRZPoIJmh8wPIH5MLV4ygM4xOnh9Cz3I5wASEwtQdyi2W9b7T39LUJM
j1wzgZKF2J6/F9s+R4zlvu7OC35at7DRrOQmbgmWq43+QMvr5rGEAil3gdSe
OxaHNLyANRq/HSm4sBRlX7cM/Dj7Q2tFYIo48Ic9xYh9ldhGuupLPX40k32p
mC5U/0kFN1Y21RB8j/TFrPBlPxfmEE8wy4v5jILPzTeWVsvO3oSmKbwqo7Dm
uDBzNbI/srxGnjH0mjxu/AkWGRiLT8LS2Pdx/IgVPlNluZJBmT2csJo2JLOL
5dni9ak6V+Q+6bmHnhXaDmk7LjT3eqZaAc4EFbVadUc8kfc6Qu+jIiBjQp+t
H0wc786fbXU0l/iYlyUqGNPXElZtN9HYdQs8vLnZTsVJDn0ogXDDs2Fk5VpW
SZZPX8hbz5P8PTRM1dHp0v3KQsEaOmnMueBFasTM8vMNEvz1E9/Bt4hNFoGg
JmG/ZUh2EYLais/j/iDXcYmVLbgbDzUAVgDndLGWD36VyQItwQ0thtrRTSgx
hNYIPNS1ZPWEM0MD7Vnm5Hp6dvTD7pVqk03Xcrkm5bEji511Qe48z69ALQSC
dFfAJbCLsywODBH5olK7sTnuP9/rQPe9mDT+73DV1uwCZLxc0qXOE9iJPv3Q
zzw1z8ZbMFUZfudeTqnYTwNpPzDfVkL6vz6w2af/PI7htLziQLGOe5FlHv0f
awVvkJj7njEeJymNvOGLncKrVzvECkem/pIyp24WMVR1pr8qoeJNlhC5QsTe
SOPiIAMCnbi/t/mSyQTqk2WZ/Y5CI9OSYdwGH15xBHHvl1GRXhUkGuhKtZ/x
139TugfBaA9cwF99xm2AvLGgSZ0VZgolDNVTTUtMUfIglUZEYT7lH2o8z5wq
2O8hk4lW2X+/SpBOwb7zfGyRf3mJkDURbDMPwHkpUj/S4cEL0d90JhSn1k9G
PuY5TEbssdISlADXxDCO2ZfBqjyvMnqp8yPe4E+Bcqco7+UO+qMkh+mPz5cQ
Efx85/C9mgrnFG37R1cFro78tsH5PGNyREz6feuVXN6KfhSUuC5KY+9BtvqQ
9LL/e/k8d3enBQ4WFQrmQjcv6a5Yvfms1yuI5Mm62whKtYEoDeb9k3P6HnVl
oNdOyKjWqvZTSrExF1BwzkveJaKjMe8Q3RhJLgsCuLSxXvZPu8bAm6wRpE6X
mCvFFuodd5uAjG3YUa51xSdrVTIlVL56J1sjImJsvR4wC+PVAi2zm8o6J/AK
HWvevA452+1ReBUbuJD71ISJpGXjv0ArQn7rrDNwq7ge1FHEpvOfSg2iwcFi
c1k3Q0/j6MqIX0oVOc+KxGo05jiQS+TCxMYzTVPYGqf1EJSgqhYxKYDVB2zQ
31cYyjy45EO9Kip2uYDGnemSFDllHu8IgoCzAyhtImY1lb6yjCpycMlbAF2o
RAVqopa7Q1YQqJLxfqB9IcR2APePvFmfyGxYludqG1sp8w3DPuqOHhGxnT/9
wEi6pPFQ69n1DqdmLv/K48RldVPgAnowt2q0A4zlNIiDv0uYhPdXr2XObTz/
+C18+DHCSs+wjt8f+TNUAn6ipt45npwGrXVr0Qf+ZeiqUncANda2E/TwVw2t
L/wPb2dodhiG6JO/rL5dREO05e+isVmHP5jpodcHTbp6/Sjo+CPANVVrrwzF
rE4ffrSHjWN9Vf2v8ESQeU3MZNaCOiB8uClmouoARbq6WxTqel8UUNaWFrUw
mDTY+vWocyIS+OOSuhOTw30yUCm5VVyDgq7uhh0PGWwMZ3F2Do5YWXoMkBJr
DCWMqpSwBgmXlf3s6rmrngukPRSCFVjyd7twqWLfDcS8GiocM32MKjdTX/bv
PGdJolNSgGbsT6FxZsAU8SWtHr3koCrOldru+Tye6bSRSzGaIw1LsR3ouekn
6XFRkPtdEbxM8Pm/Ji9hHiUVHWDFXnaUC9lLCCrSAot68KYjakUAIcqOUDZv
w8Wcfl4Ew3t1OfaG3hY4oPuBkN9uLuTc13603y/EJoMDWHiKc2T3v+0lh6sO
q/mySxcfMkPD1BhmW8tymn8iSaUK11qm9uY9fLASdJr0EIPAB6DAqaSegklS
nqqbQhKnNH4WrAkvNpwMFJXKWH7c8kIvaWu7B2vKfJromZigWxUDjgCjMDRr
ZOMWLRKmePZpZeNKtsqegp2rjW/dlwrsvJGmf6HFygImMszn48ecazdZPbRV
5s7nqQFANy5P/uVPTWDVUZcot/biD2Hu6b8uKbgIcvSP5s+TLWo8wqxVGVVt
k7AK6w4UQZad2gB9Eb8T72Uf0oo50lr/L8BmNNUoyPbOSQ0Zws+TgzJPqtj3
LUNMPVfOGSNVUbMVNuU/LndgRPxfsdBpBCrcxNPfOTYU8GwJlpUFcNZgo6n9
F3Ye6TQGHg9i4w4f2+x/ppS6vLA/7+SywJm4re7e+yljACAYwJ/ikg2++46I
QoPBOWqqweNpwv2RGZuGIoTnen3P0SExGZJYrywE+jpfv3BG+hRF4Odk7OYL
CV3OkpmIqYNU3wew/8FVhRdSgWKm+pb/svV5xgMwJEd2DGW3eBT0me16x/TR
wfSNHv1+UcjioPdEqDs9l8JiSklndlfveG+doi+CfPfG3VfuXxCc1jpMxzFM
P0YCk1naS/0jl23xD3djIMtm7F0KIpPc1d17YX0LjL9O9Rwk34Rj1r8DK0rp
d/6WVCzgk3ex0ZLL1w67NTHPiX+XGhuwH+E4dsZhKXg1LUMilgmS22TZyi/H
GwcRQOT4GqRnvZpbvN/3mlRnB6HGxePRmvJFE6AIVOuAA0W2FWlxvnEobo/T
jWsf0zy4cNKUaA0+nxPJNfhbJKhfwxtnYY6YrFmrDilCc2fYvNLMgkNEuVye
8X6n4ib0JZV5aCppLIAjVWey7jZMtZkxlXste68VsIIoePn3aeHiFki5Hzdj
NDO1ZTotZdIGIxt8Vvd8EshFDJ2L0cD6BBRGay824edaudt9k8IaRdf/75B2
pmq3mHZT8d9yiL5y0E0BxOmAVDeZqDiCz35I+w8kTR/OsSV+4FohICsKNHVq
r9OfTPXUu0UZKaVDS6yiDjEc3CkH81J++OTYWHWxvSVVlvCUy4iGwriiOtwB
KcCxPNgRhwB50QHlELlwdV2f+b0I8d6jMgjRmR4fnS/APEtGnfuilZAEk/vs
xXwaURSkSh9arhjmgfnbCMr3hK+ICnyk0+/gwby1KNmDRpJ8RNcu2NlKqYFh
8WcVOUh4rNa/FGeCl7rtuB3Uy9+fPV60xk5dlQUWZOgxbxT4XM7UE5tzaZLh
uhKBVLPCfTUC/HUqKkbPJKfmzTpMFJqkA4/K0Q//DutldtNdXSnGR8n7jd4l
Fr5SXm9EV1uCyK76zM8+xpPHmmXpbtCg9mf62sdtaYmB47ecLKTHBujKJF4q
VnqZGoZbEB/TUU52JTPLavJcoEXuBk0HwbHzObGaNWKvAoJYwOWk++DTVWkb
3gNEjMMv26Y9+Hil7c7+Rly2gKdtSg3hTT0um7jCktx6wK0Z1Sd13xy2QTJu
sKCxQE/XE5z35xlKmU1eorMJE6oWjZSOZ/+FX+WpnpHTH89h3SxQsMWGWgcq
x2htVEpqWOWjvI2xT8uYdpcSzDN1Oi2QDM4OCoyUb3WiwA0CJxu6WkHT6NAl
r7oKYXdESduilTz1q5z0KRE0AvdiLFstinsykX9g4b8gAs4EqQ5ohtpcEqhN
o2IkdR7vMx0vtKCQ+6u+09bMQ395U/H+XayoCNe8EVFyKdPrcV9IzDiiid2P
I1oF0S2dq0wjJXWoOh2SBxngkPm6Szvh58K7HHR0Di3F1PmVBfEiJSAc/qry
l6JlOCu2dFnpLLx+/8aJ151mtHkqhQSFkIwrzbIFo8ABauNlhn0B2UY4Sp0C
P68167+SLVvy2bzBxS3ulAkX0OQfyIZoSUhYqpPs+3JyXJehnT1eQFAO8C3x
83u9zdizq7EBQvHeyvao0UmJn9MTo7LA+L2igTi2rATTa2+W7PHH6gVrRjIk
L/6XF859woXwzBTecpYBOE6kjaSYCMhCJNH1UgPZi2limRPNZwHkXkAfWIVM
ayMthpBujfPJoEQ0nCx9nTzyMoMYUCN4y4Z2eHylQlupl5X2C7qR9IkCTN1j
pXIojD+lQZ+nnuG3uKe1PG1zHvTdk0W47sdClkN6CPQjisx5vmMTteZd9et9
Lj4g784fQ11G/Amq8hC0fcASX8e1ifAhLmtzAJXnKlprKK6wKCkjoX96u39M
oCwGCjrl2P6z5humwqL3CyvWQqHkIA3g3BfTwk0RP0thb4ZCrqU7xnDq1PWg
gEEKvon5ML0/t0Ypuj/M33HvVNMrh2vQfvj/f598+q6a54dLBNorY7tyeHu/
/MStZs7pwmoRJohgcN1kd7bN1gFf80wGjm21G189QZaHXYexg2gpF4t3sNaa
o56AJcYdzg23vnLDSHm39+XokLkQgw5wjB6sUs5STIU2A8QOfBoRoqdvGi0K
21Sub+RhHHaCx32bbTGmjlUqYBcFdAlIT11MUIYl5wAy9k4e5ptQfZ0MKdEv
NrfUeSE4ahJewdobC7bqs6pip1NAN+pMUg8EIr9lZpYmYbCq/SZBymUj7Bfc
o2CRWDHUh/gs7S1wRvdytfzNg1gucHy+eYDMt3Tm1va5D/HUGxsPqS/Buwtg
0c6CzzCeuFqtN1GrhmbzLbpoQEBLh43K5fgOyidCsQ2/IA1sGOF5gbkQDwXK
1w809XJjzvXsmJ/21BQIopSbbuy2tt39hpBa5KjRn5IsGhOrswAwIgPBlvqk
BjM1b99hfm7dAhaSZRQF2Zvo+LE8jb1WU/gjg4Q5EWEJ0buE6LpzzqLRPebC
FgDmrGtpsW5VWB3at8ysKD2uwNyxi2Uu+EPEOeZrjlk1udYwkOf75JMNq33r
ViEsy8zkuBBxe/vBulTCWk6BlOrVlXB1ukfsqVUU409dNlZPG8yrv1jy3S7v
8G1fePdmP8/2RC4LD0VQa1aGNXdsfXckX4DZ46ZwjDffkrjL9XmlcFaEOIil
GY77odWtPh3nRCC2evefrhzn7H0a4YxowpOX0V2uaElnBT88Yyx+0aO4r4xy
enBzUGqquR0Bs4oBdP3y2qSIqVHkcWlJuH4BMsoQ4EWDBvNRpZJyPHuziR+R
KLZf8ur4vR7LtkWMwiBpgIv8DXpIwfP8hv4LPFqpPshnZIN4ThmYizMAwHPz
RYtaSjX8ByfVJRM5gFV40duYFHdri7Ux9Kq08HpGe2uFNw+CoA561wYZR9WI
7vUrhH+z8hh33BpOc5b5CHEumNAoMg8DBuj0oKrzixiDS1TlOm5xEvZELm6F
vh9mZo6pjVf4G9qRaX7LeDV4z47z9aIcjh9cdQxaLPjrSKg4H81oi5dxZax6
a6FIFOxokdNfowic+k0MwXZK3v8eU4cP9mf1Ar9ll+fjuMJgjwb0UE+GB98s
fg9xZGk311f5emQjgKi9P+89VSyVkTcSPtK1CRGDEHmsTSbihA9zMRje88VF
IIqCDv50v+qkg8iwvgZaYM9UC8qqx8TBRX24piPMZIrwQj1aEg3bWF53xL3D
vkpXQbc5363ISqYIJTdDajZzQ0CTIfJe52wpPmpm/p84P5a1c9C0xF5wLQtM
uRHBYomMQrseu4bku+uLWJi6wHBUDlIrnz44GYRq7HRv3XXHs4jX86ewN7CW
CyAQfR3cGbEtdAWVy1uEPgeiSrc95HppJAdRH3AzCC1r1juxZVJzciq6qM5C
Jjgsbk1Ww0k+2/xm54QF+FrEpMkzmZBzRjWEa27Julmvrxig79L1nbkdk3Us
o9NgNsWK/QvgGubPifu3wfhS/XloTYyRblbVMwoRPnWpGyYgotLuyozfl62F
4kDbmCD1Gk5Wv2H2HvXO37F6x7VrkGb7PQvjgBUhQy2Dhqsds87HifsnllQn
Lb/USAzIvV8IoOI/mQOMmwxd9s/Cbcm+b1OKD4FBmu0PwEfBc115Wkm3c4wE
1uMrQf7dv0m3ZDHmPB1Glr7GwhVvzLcX/KjeGW3ocLhU1rHfSQIMEG99dOkE
PT5Ynj7x/xxf6pmarbAvNu5mn74DRdaGw+s7ZeAcF8WdTaWRIN5KbFE4RHeR
A8X9bhJSIti7yAlcZl4PFHo8/q7sH+I2qPsSKWin3cn4lLhx3jt8lNdRNjqh
u+hmrcvm5ou3va2X0mEY1XsV/YSzaUPMfCuBkfeZ+qGp8ln6bzpIWiiKL1XF
mDiJ6arD0JqBzNoM/GRfRE+bpfZ/oYa4D3Hui2HjhtTtkN1ZDP0ZrMSkdqag
eaDHlr00NLLTJmpERbKNe/olBJPODfhOlshk0vZbdp49WuldRChvAeQpXddw
sPeD6cTZ75XbnGmgQfnXiK8nzo+M17dpvMXPhw4OnxasnxVf0Iz8GWOkEigA
RxNe3omiFKp4p+jCIPH4BMQyXP9L42dSN6CnTC+2G+AsEKBt/kM/FTfFzXhl
X54n9Wmh6DojEHJOfOcu0npIbuSkGRt2fwUE9DBIYiEA+ctSDy2DctOj6pjp
mkqRWweBtTFqNoEGlrcNJW1fYeZtp3b8ZNnatroHPH56tCy5COEk3b+gKgLM
G75sJJRK1rE5AZSY05PfFso6L1QIUaEg0tjcPwldFPFhcRfkspBkl3zoHtJ3
GYr9BbQcmc6czw3Su/AQjr78tGU4NcZ801AWhZtdzkUu6rw374tISL05OgRv
U1cwJcBycSHFVPZH9PKvZQT+kpxriJwhhjx46/NTcnmAM7fP8H5XT3Y7CZjc
zx+AR3A2R3uY5xH/HUxuBTbV8XeauN2GHjbktwvVHXJtDIJ4uhzXUErC0WcT
/M/uxJMwdnvLbim1iv9tcqu0fv/nJTLBI3VrhiBmAxa0cxJTwayJhsupZpDw
MuJ042blWryxkZBNUR9TOjHzrQ2DV8PT1C8Vtv2sQDfGJxceAgQ0oWxxZuTV
DGXr5m3kQVE4R3RK78bJhIjifix4SJhC9SPdtcd5kLcBUnv2+ZH0WdPOUawz
f9gx319lKmBpufwiIDsqz9VIp1MaX0xj6ZigA9hzMJKTmgMY4iCxmnxPODAD
QnyHKYq/TJ2hx/F8UPsHeJ7XNdVuffzjYzAlgfZh+myOxhoU20dWJe4p7sy3
QB5opi5vVfwVwt7gBKG8JPZ6W/48RXk9W4rxyOOMLIFPZZAuDU1Q6ePYmZX/
kms8Ou/Wsh/KDqjausv08HUHQOJMHqAqh8nagJI3C3ZxYsRY/S7PyozDeVB0
oigJXIhYLRFrM0gD6afkNDzjvcPYeXmpbelxuaFUjZXHMF5hn84A2k5CS0ET
P8g8eWlvkILBd2mRtoHuFwLuMq438BJNwzb9Z6ezK7mFpI8J8SUROA5rZEXi
geHK95N+wrCdb3r5Qzn+pbH+b/0KzOz1ySlPoq/E4N1HljOXYhkYRbzk/c0B
qYfigyj67AAmvoAaWwkR/Kk1dj3CtpBAS7G0i0g4aWhrD5s4I1yqdLPUEsrP
geqO+A+Ya8hzDTNy2ykoD0qv36lWI2OXSda8kUHvijlw370r4T18BeFJa93I
umMwDG4ygNVjONvsghPvOm4ZB7BB9WTSD9BoodaI6LIEIM9bvrSxKbCpvAOg
KIG6R0rAJ8MhMb5TPwzxgKnSs2SPZpcohmiC94/fAvVAR7VneX7181YM6BF7
HriGzCHh3C+ItOYVS+TjzH+iTG0rxcf0c2+xdnevE6Koh9FH3o4/Nut7JzNI
Kb//FLMHq6JmeoCASyquX3I0ewJAFdyRr13CPFYIuuGu7Ww44YEZC7ErJG7s
WcnU5H6c0AyT9Ml8fa729E3//nDHA178AK7VYSDnikg6e+QRrb8nI5kh7hzT
s4rF9dk0BMoT+/wXNbBw7uHKMg7AtwBNjhk8cDwS52spb4rLocjFof71rcrJ
uKBaaRBxyf8WiN0SJAOEM4hFG+f/vq6Fy1nmojvJK4MAkGxgvLQp0jv3XoHb
qagxVHYNMBjOuQVqr9pHwIXHm7x8BuvpR6at93WOy0oYRnOo5Vi/RTLQRZtW
9cdNpwUsSlxdoqO5PZlU21ae0PZEwMRQC5FCf9jd+FGfCsBH//rw/fTg3q1q
to/9rwEdKteQDoFuy4vRBsIJZZYDHhdQ0rhTh3jELecY7LRE4XYhhZ6Yi7nH
PC5sCSUgqkJ4CjGOfLqOFEbvo9tbN+UYMisk63vRvK+X5vwTZzPUxVXcRknQ
9O7YWY2Os2sLbmaJY91YSwIxY8146vL9s7EiDFwR23QA5EHilF0Cbved5jgM
ly0TzbjIjLTiNho2VFx8+ZiUmfhnjlY/58EXvXk1Rf8StavNEgrMtI2/0M/u
VHyfTeN3YLOuJLn4dqH7X8FUI2kNPTmHLrs9WU06N7E2cQtsfSPBpUzsr1Rn
utxfX0jhzCH1Xxk9qZo5aMR8RbYSrO2WRC+0zjL5iaX9nJy//UgfayRekRZn
ftzOBJB4/l0Htthb1J6GlI5syPjk4r3RKAY1btKfUop2ZHxl5kGa3164iH4k
KMYKxnB1VUzN+q1dvmxr4yZYSk2HutWaP93f/0yaYO0KnxIoFrDoB371kPcM
7Dw1+JOheZJGJZgpbSWsT7gg3rOJDThykPEe647umc5cd+0ql2i2Rp+17QuA
6VFmUlK3kcodci+d7itFvPHWG8z6lDV6MoodusrVT8VX6QOo5yyBYlF6I9Uv
ajW1Fyde5GXxPTQXspHzY1neohTTj5Thksu6Z6m37j85OFE7hoGB/cIBx3rd
U1JM4XisfyNGdtWtclzE6rXcnrmygWfJ0t4eIY/bhF9+8qqRt0cPBdu8nhpI
tus6XHGI3J/uoI6JyRHDgfTFOMEi3lQ88BKugBENPQtmjzNQeCGhzCp69S77
WpHE2n5kK2USdVAEYnNPwwfKBh8qR9dXt8x5Vme/bLP2LieWYQYJAePZTuvi
wi6yER7C+PbujEnpUaXgHSQr7CHItvbLEdlSqPrpn8QxN20hIfavjYSvmId4
qS4MVuf1weA5BcLpzaKprxTdPUaZp24bhGPPXkuqM2RTWNYPiCgsonVfCR7K
Zhb0AMmXiHLR1YNw4e+1X0SWeJ80HTTNbhzAkjpnbseIQsHl5XxKhbtXr/So
Qc2xfrFWSqdUocWo9dTbEv7vm3dJHL1L+Dvsv284mRCUXoG574X2TDMzOe+F
cCCUCVPKfUm+HjH7cXX8ya0XboDYCcNSrUgPKtmI068rq5Yu2TCJ+N3BSgHR
3S9UpZ2OEI/FU9ifHgrdeGfQkGvvhxQAOge77PA6RyeorAjTyaQ/AI7w4EGM
pV/O/NrQHcNG8OmwJPqhjjvMgUzpGON/+B0VDLTmxD/j1hhlZU8x0aJnDXaM
8WzXINwS/jMSRSl6sxhv/fxoDaZMPsnnvtzYPSb43ULUrcxkwsZUo0nXNDzL
NSw96hi5sR2aiR2O7aiSp36Y5i8HIdP9i/mk/lIng3kN9wsdIbSaLHk7lq4t
FyixZG89F8HOU6ZxGPwAlItqYj+2v95HvQvjSCfno3pteyobrRhEwqfDmXP/
rTQ2rfBg1ggUO/FgnqYh3rH4Mwy5ZffCWO+qSx2Tq+zHyrh5s+acSVZFROZM
W8ygJkKUV0aM2+0tWVl1nQr2VseQ43DcCXfTqDYan4yqQ4Aky0xwannzaDAn
HQKz7nmRsX1SjbuUGINjjgT2prTcTVY/0kgsxBqgluO07Ds29BJImymKftJi
cgPfpY5U4xXW4AgVLl6A2H9MG6eRJIDL7xeB2bTBcPF4dUhk0MzOEOr84nM+
bTLSnxg8gmOOBhtVRuPCRG9HtxU6YxqgU1vCF6Y3rtvkbCXNMLYxSrWwpp6w
if5tEyTJg3SvqYUnel4HMkfIZ7tik/RNQz7ciPOLZZDZfUhvcQUQkeL9nsDD
Px1QPG9tt9xkiNHY1Q+HAnG+kvuCvxUEY5nJP6rMP6qXZ/a7Z5vKL03UGDnE
SBrCjlLk2n0/07JlbrN4d7yRKlgz3lAk32MwbRvDr4h83yHnQEEHx1L1EYvM
C7ohD6rxZodS+0ay40yfXANGi+y/lPlQ6v1AY/WjuPIOlToqT1f07RbAcQ6s
UPIaXWD4609gEv/MmnilNtjeWQL7c3ofCpdYT9z4bCPR2Gf4KwuhO1jNWgTf
Bc2/dgVMENTW7QQfMwnftNdZiMDk3OsJFhnX5tkWx+kjdREewxmpCKo+t+QZ
KL4QX3E/5YHcvxoNJ4g2Yg/j8t2WL+hh/OzNepRwx6bsIDNh8ap9LqZ6sd+e
5BZ9qSV8GeHi5WlT/Ab4UUMMc6quoIn2Bju5wV/XPBi84Io1KB2UVzgFcNWy
V+VYic/SuRqzA5E5XfZmKRqjUBW9b7JSQ45LrtXxvLSfI4WYoTkX6Cb5IPoG
5QHxT2Qkjb0/TnJ6pnuPUWISrxN8jJHztAVezkQUmR3nD+7N9/CnWB1jS2QS
IGEq+gwuYh2rzkaljPdzJvzu7ccSMnG6VboxRL4PRJBddnltDR0HW6iJfoEU
Cl3pXyiTsKKA37W0bqrkAtq0bv1gNFV+lL837aX7n/RbfkW+dLDpCe9T3IML
3HGvCg61cFzlkP4pgx11JSJYGZ031dJRUvqJuHeCF7utw3QUS/sOnipo9dUW
681ddeftOUKjscP3KD+QGTUzI8uR0fzlWlQ/sPY/z2rkDQCY6wxxs6u9CCip
rVetRDzkKuWLg4vuqjk3AA6Vs6gDLV2iOSqsHzaHXuIJUzeYS4fUJInTb/kL
KJ4agh6tw0Y+haQln2tMSawmzeSD/yIELbUo040DMlmyMnoIvehYmQ70q3zt
8bDuDKt3HC0tUGcxtHyjUl56gqRfxTdGExhXNLU5R+X9BFme+74Hf7oMUjsu
ANv/nEj09HaeddsUeqKl55i+g5B2qwrP05b4dFv0uOSeKxkfucE6bqOxnykW
fSLE7qSprTHRUGoHbCpYx08rUkv9hL2E0eg0s4IkLf5JNHtVDWcW1QYp838g
Rh2d8aPfHvGTtJrp9wlWu2U6lrdS5GDIdcL5P3aTK8DbLF2/BcPP5N4YjQvr
k1QitCD69wGW6kq0yvNTXb7sH3DZCHcBEI6vugyrZ2xR08Ir/lVQydMZpxx6
78ykvs+oO6ejVq0o7iXsMwP3uGPG/q+FuXDBIYYSkV3ndXW70oesjI3aKX3o
iS9QFbI19tLQj1O6Fq+kRWe+HW0UqP4xyBw3DBL+taDhMC6xEequNmjJDEnJ
G/517IvP/VnFFy/LIuyfkyQcDQg9ypW8IucrDkJZDiXWj7MT0DYHyguAGQA8
rMLhZx6G3ju9YP6MR9ZJx+W8JCLZq5/NFUytrfAKD4CgYlszlUqn6vaUSH7a
zJzmBemIMeHAtWhHr/alW3wErad90N0DdcHlbl8jDWrdRaSrntbWr5pfKhSV
J6wiWDp+3QLxiOueUmTCL5C5YZcoTICaKTh4paLjOV/0xpiGkZ4mTkCrjzu2
9uqyrX/CJRZPy49iig4XaaIFnqB9b/ZksDwLUxtYuYvIhbKhmo8rpy+Qvhq6
LPua2D9KmZM5O9+BESs6t1YZdZkxEeSXtTz2QmcNH0M8IDdNAhUP1qpeForr
LVR0mg0bIpoHXqxNNUaohhFq3/m/urechTZJIy5VEkLNvojmM335oKOD/FO/
mlf2zz6qBJ79NvOd5wa6ta586rvqJZ1mgo5FFYS4PVEAHTq/+/4SW3PjvuC4
imKpL5CVLXg7eD/Mt4pOfcRzwlYixHHW5nSu+mQ27FAkBwISgCC0i9dF//zG
2v9HYRv02eRUgY33GtUBwm0SP59SexF56TMpuedgFcKu3+Y2YARIbl4alro9
AVXIswkwlD9hVqdS6fXnyc0ctMJD+eb+CrZ+EqZRr/Kv81yGp5fq47N01vJP
kOScxbJT+SQvJI9d2erM9jjsi7aFNnXlGgHAiP8NF+nxNmRkr2qtLqjUYmeu
hXZNjTv9yk7lhDimK3ZQh5twfCi6k9ZqW3fRpKXl83T6BhP8hpjIG4WWaU9y
Q0dxmrFt5zNLOObiOMnap1hyMRUkYHaPwsKCDscF7eEcK2MmQjitb6h1oV1z
k9VD1QN7pRh24cUY6ExTt7q181YFotD+NhWzHShK46laAjznC9gb+1Zki8z8
C+rPJCHgtIFjHquZ/2pLrPqeFfbomaFDoTvCIjOi5YZ97xMutRqamAwpqC7V
e6EqAE0jypzUPRQPRuIUsoSeH2V5P5103dpHbALtkn3g6TGNjCtrcRuJbDQk
p+6EcQlL5ZrODMENtYHl47L+ctCZy/SIDr0e/EmJgecibmoGJMPT6Wde/znQ
dMf712gG5SAOz8+AWOMXcUDAII+IFCJY/MWDMvZEwYqAQcfCg9RyWW+P1pcJ
JagXuJIiOtjcgmnyuPUcATO4deBsIwXSXZMO5vkKSqTX+OlwXfqTbOdiJ3XT
6X9a374ZdpB/cxQ62Svri872s/yIzC8jsVlO/Gd6Gn2kmT0dQ71AyX6wITKI
0eZy1b3TjeQ9iGYY5AJaC7Toev0R6D4JL/SXPHXh2/kt7FdP9GoODKJnEcrJ
SovMd2fQtjRES0m4t6SebKbYKZzmsZWQbhPl3uTcDTxfR3k8ng/+hNmzDdT1
/qs2bYsnZP65PZ9NNimxHMsfm8NVAN60qKZdN6ilvI3mIKhGbsZeOKeOuPd3
z64AMVImY4PHHQSY+hWOqul9nR9qdB3Wbz9OWBQhY4oZNeI082VTg093pu/9
/I9LAXNg6xKzDNK64CGzqL/s5dAMIhKb/q9YXP2wqM7O5pMvXRnXtayOfV3N
opn2j24sREWRTlPoQizLrUSg359oG7IdB0Ep5o9YdT+4FMXJNLRqN/VWbG9b
Z3afp5xO0wwHjz0diy9kUpVLOnVeZSpiXSUOwfQPizqnVIlegZog5jsT4ZFM
L8t2WL775Y6GQWZvHTU2SClrzHAWdK56iXr4sGlukz6ctsvykWbAfdkdlnYc
Ck6cuWYiSCAAlTzQ38lirPnju3SogAzqYz78Ay5TB5LNoowmsq2u2IFv0gED
V6ZapwWhw+RTSNt2JxWahZEioVubpbK5aNNmOTjdcqY2QMYtw+KH3eaw476Q
x/yrhlYh1j3wxvd90OugJW1elmFU0HI+Y4XAjwcJDc3eVt40EbWlBMRFeokF
r7zQxhdXPBP3+D2jfstFoOG27Lwvl94PKHAYibcOvjkupipBx0zcT1TQ4pHp
14fx1GsBRuzi+XsrB8NtVr3IaI8w4Eyyt1aUaKfkzcmcyyKy+HLUeuPAvDhI
LuBf/N/EwRBDu/LHEu65rsm2hUp4UzrvqtjGChuGsXrtNCenn4atkyRzBHV3
b0XN07Jch1BtlomWB7LU5xpbtZZtWPfIKtoaT8pUN1M6xJkxSbeaETHev55v
tDnt37pSB8MrmBQyFsbxksb1uswPYVPkvEkFYTt0bXCmHMVw0i+cO9G2VHPw
eO9yZBw4VBzPZtJY1NZactRMitvSiaoytWfRjq+xoOZCvQKI1+I/7sUKa0Pn
CyH/uHBedyRt2AHthV9XfhUysL0zckWFKHxhG3VxSCvJ/iXjAwLXpZYDMWBj
3A+MEOIm3wb/5B8MW+POHWMXFoX6XkcyXyw3FTIE754ALLNyQo90h/Wd3xpA
qZWjmXlU6vg/PuK3dqutDPMnOcwfafoYUEuDim6TbhRlN6CqQ6hTCULDD6Yh
NcmY8AC+IzJv0yQZFCR7XEzUViBXjsqTmw51hQVv3q4tWjbZSdm21edgeVvr
epNzz3Eca3V/O9vS8Gs+egCWN8IearJ31j6LbiICncOf9OITST8MWOHwlZBi
RYZm8mLjqZHhO3YkEGpyt4U0OCPS6VZ58Wk0xyEyqCnetk5ZgEDu7T5z/464
a1L+0d04zI4Rdr2O3hPxUwquZWS9S3BZFk3GyfgDv+eALompbZa3eCXLkIs1
WULLclrPf1VUA8exRPiZSp1Gr3KQjw5maPh3KhaIcaFeDAzTpf4AqJRD29Sv
nkUxFWS3jzOEEKWBZh7UM90g5w5qjadf5MJ2xiOAoIVM6Wp3x1W+weVezy9/
8cioV2pXrZhHwhRYHUJ+n1cL5ToVx725SG64a5B2uMCWq9GmWg8t4eMY/30T
4fyk3G1nbKWDKSoeUzuJX/vdMX59To+J2WoK0kOJ6FkKYr/er29tFO/qhTJS
2gfTczzrxFvkdBrl1Gz73AjiY/JVRXb4XKp8avA9FEnPOAtMxrHpwon5iKLU
SDxz6TQ8GoqnPuHiPnfx8cw3MUumPsy/Z0II0SfFN2jDdghhilpCP/NyAY1o
483cpFSqy36C1y0pGRWP4NjpKjcA5MgzbzUs9FfLxKWi34ASmpQBSMgWJ/nS
ErCib/eD9/NnUCXmeCk+09NvZFPRqxsMAMLkxHv+rz/s55gl2hVTQwuWW+DK
nvtYK4xMa8Ba7hDnVVQH5iyT0um4F/vXPxHvnbCK0Faeg3D20fm3kMgltunq
WWRMFRBEx8EJGoA3s02sxNeD08AQvrKgakDn1T66zAPmYHfnHivPsPSbnh83
hp4UO1vyQcqUkIzWPR06WORrNvSGhqH+I4s/YSxyFNw9ZufIHPD76KSeqtaQ
AX5SqnXDPR0mjaJSlKsOZstjBstV/0AMzfGtffiaD6+K9yf9q+0Jt0FlpXMs
PNhbzGDhiKzMauozdHu4ykX/1o864GALPbeAzKaSDNDY4F1JZ5mUrJgVmkEJ
qN3BsQ4DcnWqw3yBAy85OXvavWm4hcZwewakKef4rlcqYPPNi3O66mQAnN8N
VSkLqLxq5Y0y/U8u8QXMp6BT1E8IfEU7x2GGyStSvcT10KesCT5VH37r056J
g+eXADL5EbJbCD/Fh7qkZSEJHXCbT2JsTjB9NlewZHiwCHm1TL5VNgHbg+P2
B+DepHtwnOKZpI+XgL6CINcGgbWI0MLlkm+vja2aIE8BEMdgIWwLAHEICwLc
uL1WeUQRlFnCd9rAnr5h6FPgbegp7qCkz1DzTusZLIzSVbBG4w9I4OQj0SH2
dL5OxDt2BuFsErUIrJSsQJiBqhuJdtd29nS4zxoRS/L9QXorFWhiEftVMk8E
FtyYLuYycM2FfZ/gYbODX92G1T1kPYiq8Yey84awhRH2u2MjnpNcOTKpB0Hx
cm55gN2IwK6ZuQMdHo830tgp9R2SLpDmidLFUz4ew13DdXXP2F9A8Gi0r8Qn
hq8xVmW2DSKIRITEXqQZngAW4ON1ChB2qG7O6hyFtXKTB86A0etUwzEJL3uF
7l0PiJYQvafVOXPZPUYkJR0H1UA0Sm0I9NcaB5qOQdzjQ6SwudYZ7IRu3Lsc
5DWU1zasbdGqv99au1OFT2qs+TvTFksIZ4A50r6r776z0DMLVxMV6eiH3eGJ
+O3aqYGvYo3g7KQTNqMNC3Y5JxbqW/UgNffwT89EzVV2XkeRPfe4W3NA8UnL
a4bLrUV4IobZUuMmDeIq5Mext9SaovYUBa/wnAS4A/vgkpezMALDr3SMULdm
xDLQBycToxnXXOJK3gvvhefFYeWnxQwUeJszr7oF3SZpORq6wwljhZzN3QD/
9xwuIefI0+ekhaVLTY8dw4vxGstCGryDa4ZX5KqBfZjkQVQM9tYYCi9THq3t
PpUXHd/laVyz+6YkEaDmSkBEIXlF60Pn+ERxr6dk0yRterptf1BsO9FCeINy
BoHT6ouFHaeWjzfThV4yAZ71BJ6wuavnoy7aL4DpJDEp4EL8JBEP37BHGv17
KRdHc5wLp4PiYQi4cGpCIKmgxD+wxhI1xy5KpKzKOXLK82F3VCOpMFb51ETS
1udpRJsU/jKWo21gJ6+za69bgp73hCXDsq5i5WINy+RdvFW5x6nNllddUBUI
bAgla1CsxOSase3o9lt6AKo6beF0Ult6rBXZfLtiC1T8JqYuXje39fBylBA4
mY7WU/mKcBxPe0CK6hKQJ0jc3eV6bOnSSEIAf9ZFeZREJiWO9znss7gYDd5c
T4/V1lMFMpzlkhSnaQ+rufDaCLiEvOXpbwn1kQ0Oz+qNaYoImEC+0bqaEFKz
yQc2oJB7riT368Wwj9LrmscUwCW1BUCEF95iGaHcWe5s5Bgzk5l/FLRqIuZa
j1gmi1FhYbdUI+OAhZ7oziAeSpoCOaxGLrI5Y282MYIHbRQDTHj1N217eSY9
RheAEbRcnIDpUFrqVN8OSmxyXpYig90rHGTd15PSF/46m1T6vTrm7r0j9mhy
A84gBdYZE1j7tnDDW03DTr3NdTnr/QcrPk1ywee7H/YiNhRAhqWwMIUOgzx6
ZWMDpifyuwjHwGIathW26X3Nfqk0+uf40Cup1me2O3EcAL1D1GnYIKTD9ENR
/vQIIVhq6xvQU+gQk6mMX1EurTtx3Ylh0VmCESP78jTdCZPWByxDE/781Gl4
20p80d/VxKlV+iSpWKxgXF2KA46WqW+BZ1ZOdDQhEIH+g287duZQWrCHQOGH
xEfPENwKQ/2o2sC4R++uu3hReJMh4Hv++Emz2pTXUyGhlOSeI0iTfISP81Jv
rz7Tim4BENek4QfdCdZUgXkW7R4D4yZ3Pzc+muIsH4/ra51QRDZMMDy6Daai
fqmRpswUzdDCn2iL9fgjyLD/D6M2emKFgTR+NumRi/5itX9f8GTG2Vx9nySa
mfZRMcxqklnO0dESCHo+xmmGRSuumO7AOCLhwvWEQgbIds6LPb6jG0dwtEO6
mf3j/HnJ26jrur8WDyeO7pJ4lZcilmsDDfuCa5rbacQCi/5qY+bKISPQ5J3O
dQER5BQsG/Kkw9CqgokHgGoDioM8oebReNGB8Gs3GFNVdl1Ab9AnsPE6ZUj5
Pq+rTa4aq6EMnK93JXIfKEXLma+WVHQo2Bgq7zFk6Ib29eSv/2C4SwaoZBXd
Vt+dfReCY/v5mSFdFjDPxN8bhPwrro7YTsjRCuaQpR7aA3JDyHs7ej76rkmo
rtxwRDvLL5JjX8NZGs59CBJpDQQi/piQApkO0tKOyZAutlqd2rdSDKXNfYRJ
wk2ZJQaZLnQyhQxYXt7GDYj0YI5n4VC8LNqcFhdP/y1aZZHxQ8mTbcacoZ7j
bHRP5madiN3lJAm5R5nExxB01aFVXzb5dGLyLXefYywjbJDgEKcjMiEqEkA2
+XzKH8WYfYbF+JI9p8Y0jqfV2JiA9XJbW2V1mhYcAfkTXzk8ukbbwz8skIyY
qr2PHXIkCeZ9PkMH7SWtKa8OQRFjmwa3K16slZ33HxQAkjZrQ8lNcV0K8+ZE
Ft7XX8V/K9mCQr6D8Gwf2pyVAx1lebz3LIMHSSZFuZMAfcnnKE6iDnAn2QYs
RM+QCGAHCR2An435if8SVTdesT5sppFiAfQaYZuf3UFNAUN+lXWX5O7JqlKz
6h4msXPUCBoH1a0dFNPB87phGwEyv8cvK2ToWhB2fhVENMDxiTBMGLCuKu0u
+DEy0Yx/0bh1mXStsEPUa1fG1sWGOVQmKg5r8K+Qiirjme9DyiaEg+UrTU7g
S8V0jjN8WsfsakY3JqSetq+8emsCGiyeK9D1nax7S6PXpX4R52tIeeB5Vet9
CZSikxmoOAF001codzheZxnvMdWvnV+okowUzsHJW6o31+rdMuV/wPVpKeMr
AfsqxgMj7BNrKrltE4le9t48d4n4f0+FXGA6P8dlIpeQxurwOwstBKqIX+C3
n/E5e+Kbjfds1JJ2CBLmfMyeoCbHsHIEWB7bkWSaXH4XpzxUdo174DFXfveX
XQob5zk3kumE/EgtEaN02QhXTX76I3KYJeQ0+wx3/eQbFxStypLxPPb167JM
XBhUv305w+8Q26fvdIDqdeUQjLOCwWmF/r9aqXmb22hv1FdFLrb1HaMDlGLY
2p0EBXkmf5nAwg4Yi8iyinb0NFoTYsk1PQp2QTSaA30HkvSMbwGiBZ1/I4j/
Y0Qt9+iFJUobercsoz9OSQ1mZdahhgeW9f5OqywlQgpaCDCkVy9MzJ2S2/vV
K4NLbe5bfK36BKUui9DoJfNKFurd3/1EUfeD5LbfN1ZwLs02jw++LEBdJEXg
13fQBGJQUYKYxZU78FkiR9HaqhsEzP/BTF4i7V3Gat/yCRT/HHqAD+8vZ23y
+OAq2UZASIOi6pmSxq1T0l/RJ1Y2Nf40nrNfKQpbZPoopgLHrcycyj1Uqi8w
yVSZ5UHV53zzeEz6zXO8TAq2Lq91GSCWNNjFOG/ZgtB4wVoflacmKcxX1owc
xovGn6bdcikWxrt+5M3Cx+bVn4crVG7mT3HEjpYDV15l7/upqRJI7nJd0Kk0
/OXUCs4JTHoGzWyymbaZF0rqbDoA882YgEjWRyU6kvLIj82zs96wAlXS+zJH
MDfPEf0/p4s3kv0+K69D8EYo0m7biV2MNgBzmg27S9+VavmuioX1Q3oI6XC0
7/6Y+YlxAaydma5bMP2Va7d3r56l5Hj9BMI0Hzv56cZ1qlXmuzl/7Eu9GJym
UVDkqHAik4kOnWah9YjR+OnxkuaKkdXK4MYn8HJoxOUV0DBS8oQchmFH2UBu
7QCzlVNWoBPVu/Ah3Rcfl3Gmpogbfg7w0l7SsEAj6DbCIxl5qvq/E5359fze
HYisKFCEY7I07LLJRNySoOXPnEfBe5mTJj01LDF7vzegM/55OK92z+LyYbLt
OkL+b+pB+AObNA8BJ6MBE46VvCGAPtS8Kf55sirytA+V/1ckRUzzHAEcIc9x
PgWWZGFs15Oqrv5bOWT04XXFqAYS4dlTEi+A8QAB0Z7fRCKpgujSwLu/P6kz
h8lJXdldlnb8DEceYg2xGrK25+FeCVx6RQ5Yj4v8ueSxe4lySvngNo2F3xH6
bUeP3FqYym0TlEoysqQkNcbKe9knJc6JYzztNKN+OpuVv5BadYrCbV4QABmP
rFuDQ9xtEU4TmvyPkuWDRSZbk9MlxjkecUjf+KLsi+fZJsIZeePNiN/rFhfu
tGbZxIXQrwSg420Rc7QMopXlvSE+rWmtGWn9zY6WmP2/pWmHZ2f6jTKQIX0D
9Ar7ee8BRWyyDwkrT22nfosZWAfEqiEnq26Fnv0oAfU9zEZaua04Tzprlhyv
aRBCbYQxdAdVAB+RwID1HiKLKTxq0r/LZ/R2KtoiFbhl0m/dbZfpkGZ6qJMi
VFMj4Wz5uRfPDafZZvqR0B6Q6dD7u3HBq6R2JVhlPcl5/lEsV0fHVjSujcaC
Cd1wPDTUqyutuGlmcCO2+3xRgLw/gW65nUSjVgy2+gpPhrfsSDbnNXzXBRbq
MrXGyiu+1mXax48DKkw7BbCstRPz9ZRW/MzfRpsWT+OXPCQBYe+YjHo3Vl2j
v+DaxURti1rBLMq19i6adOe1/HjkjxaaPYRZiqgAZD6kF5UN+8pZ4pc31OP9
U1EtxWuAVipZtxYzdDtTD7AvSmav24PKhycSMpVecQO6NTygAH/lgPicILaI
emDhntIQl0GE7n4p8btjyBnCksYHxkiMMXXTvJ3d/5LTeqQjfkUwB9UuVhS3
WQxJR3U2JwUxLMlb+YToVF6CkZlTi1DzVLIfMYODrc+Xa2Sk8AvujzpdCxlR
aqun9lx+Q6NMWppgoGzR6TGOjJTb6iPNqW9tBvzNlMb2gzmutllSE6jrjEgR
jjvAIwf6hxGDcopXW8ViTOtDTIFWmG3std5N3F8dchiG7ZU6XU9k46rrnIZ5
3f54Ko1kYHSsL0VTLpdmThME/zivQus8c3NuKy9duLzyR38vNDHxgj9J6izk
yWwL8eMn1aXTggQ3zFXfM8krvfw20QnuGI2M2zIbHQp5W0Lty3mq1JVe0Bd+
usYa92cxSrDs8byr4f6E56DlY1PFK75wR/brk53E6I5RKv1vLZj6BzMOszQG
v8rm7IXT01RMW0YgS6pEH6ErGI6K9y0942dIO9DX8zPR+DdAABYfJFe3klbw
5qUyQ0XMi3VTWZ4n3q3kdM35W/XNCd2rXs97LgQeDfUrMwbDTk7KcRPfvIVb
uw+ozTGYHGr6v1a6ZBf1ZkqVapyUGCN76A7Wr2tvKaajhNlcWNvsgY52GeHa
cjadh2rSqWlh21GI6WahlVmk4MJy9lFGu3fpwloe1f+5xtrUGpqlx2oK2QOq
AgBlxrZBlW6YaXsQhARWeHTx7CwzzS0uwxCN3zjJQLxstNXHLcbnq46EIMkl
rvX7iUt5GpKdbTyK57zR6VNmArhSBm+AlLW6ai/DpzzsCHX5W86wjrfwVeeq
UWzhdGA8PxQfnMXehOvkH1h0h0RkatVf4HYhfQexL795TqatF+K8LXJUGcgO
Y6HHUXnzuHMaKokPWsUtLVPd5RSpsnLzdCPaR27qhniEKc4rXYgf5inZLmHI
iD1RYaKXPUIkBmdhOb9gsjv7cX4TXX664vqktj3Q9HoEcIxzDGFSPX2/4b5O
4d15K1/Lg8nbpQJRVuqdWExJ4rdbO69oYZzNaOloCXvbIxTRNxf/3GhS4Smg
OzS6DCJIJ6NQG59urCILmSsJhCKbbM4rHrpvntHOowk+HO0jblV1gWfBrJqU
Ulr2AAJrl1omOURvb0VKHODnI4R89uhcBXmssgCHSnCdx4CV+6UWkKG23+vd
ZeX+KE+0yjY75/+ZXIBBUdrnXLgrkkqGJjD0YXmrHFwVvbewz8OVnLHGFHEp
TmJt7yeFtRXVUtAZK5BAt2CNTEGxJbEOoAigv/NMmaC+ir42BJcgBJIMTWrk
nMGq9SX3BHgP/5RUHS93YEqDsqqTra/avzmY01Mb4davAljr2Pu+yfPyWcyS
JTBLwyF1t3mL7yG1jUtDhfedcyFLEaKEgODC82eDyYLbnrBQ4SuNgEqq7or2
W1VOlYO+bYdfSbJxu1Db5CrhxpJUn2vPoyMkDpn80VfPJstAsTmOCTrLkF3t
Pup8fiITmnyixCTVi1O/4HE+8h4MyOW1VtFXUFr8HzqM2O77eMi34R/Jquqy
34VVPlnO/AjRRhzxFO0vOybNeVqRRZqgdDFlVqoaySIpq7eFtye0tCeAwvOC
K6IVGWhQxAn45miifLZVf3Yf1TWBuh+cRlP7qybFmAf0AjZAporFroRMdkl6
p5nHwxM8cqpCYoO5GOxsia45Zs8UgZ+PHsizkU/U8CPrD3i2lJmZfvuzUKpI
eqfTkOha1pK7Bz66g7FhZu3lc5GdtToCht56D/gPNUrA0eEgfUxLYtmw5D7X
xAIUyHmiNfGCuuiNNEjBq1DLjqJN47yTo2QaB65tF3BMHHHhjOZSfPqfro+z
NtSNEkJ8c3lm7+OW+XxP3h3otExkqkoz1Q6RBxt88VkZpkwmkDluUJ36oMCy
AnFZK4qMCZ4oM9RiRtbjRiDMVjoBqafaHuPkkzH54pSyZwy+6znovpTt+QF/
kytli8Tv1yuSK0oEiH0mBCd9QURZgRc7jQZlflOpIwastB0Q5g1X12/Ezg8v
AXHKMJi8kqGO7WBq7i4zaXoJN4+gGwI4wCN8amhCRT4s+L3daIdvyMCMneHb
X0QvspPO4moITQ1Gvz2TXuYeUngb0FNBKYhABauuLJ9nE5MotyNdAQWm+mVd
8DXwVGCMWZC55AI6l/AfzD45lyzZIf37hTQ49sjnX0lbY0/f6KPiAV/sPuDm
sz5A6vuK+Rz0AWh9R2PQ1yrKNvFdoUCxo/ID8VsQ6wWTnJuVMuGRiZN4slix
kOCOWuwYSRRCaTVVJ8QaeECjih9OI/FNq+xvFdfQnkOobqJK1dpm3HoiykG9
Sk9JWftGOneIuSKKDOUVMKES/v+pJLaQ2coHBuPVtIPHdwOY+d6A0LA7UzRQ
mwnETJkIoXfoJ9gZ1bU0d8EJbe7hZt6aKYxhig5m4splDHMBvcKZewxuDJ9f
ybCDcLb/gGQQqseXbONrHRWVzwH+bm14rGr3YgPZSgoTHrXt6Fjm/sG4QhEg
4B2GOekriD2KwB7jOkKDnSxX8/VNtqJMWKeJuyWZ+Z6Nph9b3DdJXa7DC/fG
39003tJ6MOElhOwN/RHSVRMh9karHNhKwcCG6nHYHiE2FCGJiVxSxJvglvN0
ztRRQTUHuM5W9lhM9J0jS7sOfEZCef0fTlsj0eIQ/EkhwmLpMg7Ei4pFCpSV
Q39LbFmE0PwQXCdra8tAuqAxVvZmt/0SOm/VMD7QRYrmicCiDXNyqmtsY+0e
hyPu09BTsX0Ksq5Uf9Jpuu21w/ap9bxDPTxWjEDv+ybgFqYU4Sv38isle2Ch
x7bSR1ONYn/EmApsBcrXPICIwhO8B+OpjO9c7fGq5IyB34aTbfBzG7X19O22
9LV6OSvJEWmb6b6uXxyDHoKzdg+iV8l/rjNvH5X4cKne+eRNqy5eUazACcGt
00hwGvItoY5XivKDNSwfJsxBAOPa9sm1C1dS9b/hNe+URhgRMhu45H/HJ7Ku
nC1DqTxeeOdHoP2I8I0RorXe0S6sP+C+aMI5rzIrK8WXRC824Pau+XRBhdZ8
pgUMF4ML0BDGazz6VMQjbrYe66YUbLPMAiQ4Uq0w5t4LlwG1aYpdNMCvy39n
9gxFIrXkILrbJWmd+mRmXtilV148OYd3PkeEvi6H9yPeInRa/CCCoiILsGxf
3GB1aeC0372nRLBi9G3jhzQnjTSa/kaIRyf1Nde5R6qNZUKP9pH74nbtshdV
AgqCgf0Irl/GqXSMUewtBzwhdHt9pybjb4xvxPh+umXUH5JII9/oZ9hCnKaL
YsPYLpv/8gWmR5u3l2ViewfgvoSVoVl/YQMzVgpDimlQi4LGoGnafsK2kQF0
s1wsRnKr7Fr3M9tIfKxO2yKAJaAafJY46ojW2Tv2oiIPGPj3repFz/w8gnoH
ml6mZr3YCabM/uf2kwDW3lDg4RLCMUoOyGLLj2MJCAAspU0BFjmRc2snfwAX
DppAODd4JYOHtFJAMtLdbz3/FdpPRXLNVvtQO8AYMd0OyBv/Ox4V7vGTWpKq
Gl5NX0MicpBz+vykXGnV9RkpUdJ1WSuaovldlLHTfPFweEAinREfI1ZLL/Ap
rasYtWMENJLrjPZub/iIMSa6ra187KZBgCXTw0Oc+OgYTPZGdDIIZBlntjJW
gsgR34WE6TyKaWzQNy9e4ym2STOpB5Naf3tqG9pkg8xE7c9IdLwhFOm1Lgwl
vUGqkFdwYwUH2A5K7KNJ01Fj49s+XBUFZBVb1k8P6rhGTR4skLX0PRGMYlkQ
wdLDhLCOARCd8lEw8TJHVn2hRvtVV0jCrB8cFDTSdXoqmTQNsQ/bUcgYzoUa
RBV+5csJBnTLo1Ebxk19FSxOJufG56pfUzDrOnrTb5DyCqjKemkoDqDQ8U7J
UCToCdlGEjkqlg49JAV3vLGOtQJPtmfB3Rn0sYW25pK8So7ItsXAjtNWvRdE
xwpPalbzIE9lAhUzXwUL6sjLp57cZdloPwwOfHeGa9UXKaXJfao37VNm1OFS
cXUDMyN7bIvTDuXLm2p7XxPXLeD4JuI98PQR6eGvvH0kR+dGL0wIs0LDCmOP
ziYfCgYKLo2seSDGU3aQInQxJ2pvu3tCll4wx2eXmOJ2W1ZR4rRwUs8gMHff
ypGUQM+5FFcV0yAhYSiATe9UktAiEcq+MOUbLjVc6cMahuKz1TCz2EJZYdF+
Ssp9h/CGRbuT8N+OAUs0ifqtRE2xquVCnIzmX2gBhQ0cY/knVKLkp++QCheD
ueFg1gp6o5c70t/VH/d5H/QWwDtd/kOQldLOUfayf6ceC8DWUgsbm8NyQiHz
+YzGImlNqqJwznvfdUHoQYoFoYt1TrXUdZEDUuTBbW+Ng9o4K56rtdxQzqq5
57AqqTzW3bY79NA/hn/nK1Jv6SI26AujoecETkKFoStSbJQqTGpoVGJ9OZK8
+i1BeQ7m4zM9XKVU6GlLadl2PHBZWUv1BizA2+sxhYpGJovz78jWI0VDfpCJ
7LkxRpcCmprDVmxlaqIuUsKtFI57uxmqZ5ytQsUUYKSRthNL/epap5PCQAp3
TdbICJKsbSzKsAWJUP3OiznG26hHERAQVYWuywsOLH3tSznnK+8nx7dtp9LP
FGJ/P+5g0/Ti9Pggk5RqN4j/O/e9OP3Dv3liRfdTBI0SbulyuJkH2O/eun8I
GfEQVLttTtQ1ZKQ9Laze+lKnelc0MDvAgunVHEht9Ta45IQH6Rai8/NON5w6
8JNX6jBaxcxVwle1RRuqdBzzlt58C1toI5BQmRl4HemL5K06GG0DzHLf6ZtV
0MHO73mRBACysL/Ojxf355ljzIiJsyP7300Iv1w5vgaoIgZkKxnp91bR0Hbf
xVMwsG4X0ZCveQSZvIRVwAUspWAjOEwujLE5rCqLbOQPvZZ6NQhyIQuS18aw
cCYAOzP1XTcBkC0NRErtf3c+pxkJIFJEJVf8ZXNuQNEVQ04i94V7GnUAgMjV
vbY/Qd1AnOibcQcEAiuNIu0rpMkMeEXYR7v/aXPHCMGFyHgqp7JadrXr9L2P
+cJVRt8BU8m7yix7Ptw2gDTHYOgbe6Jf98yOw2bHMEVgdOynX4F6cFF97jrL
lWvMZEPQoCDObJu/N/81L+lKfri3g6WBryCC3OsHBHQjJWk6SPFZGhaJuxHj
mgZ3ZuWSYTnWhYLLeiK7l/ImG5ajwKZxfg3+bJ/MD1iGiHOO+Zbkb6coBogQ
jE78/aZjZBl3+pe/QMeo69PNADHq3Z9FPhgD+W3LdRorup+wqUTDmvRFilBE
g6NI0tjNO1P9KqiaK+hqeZrEgf0LYIhdz5RkH5VsX91wO0RrZRWdXzZC4zjp
65g2Qk5+A/x1G7bE9Z3iwL6+k8kLArhAUiV8jnKotZZtilKdBDxNVStla/m9
T8fm79X7Yct5cH2udGy+3UoCSCvrNvkupAPE6fWwV2t2q65pfKgUTdQAza/y
Fifargh/Orqeqkw/AKiZ5hXMIEARIbvgTMM7h/TGBGODWKeZyHGKscvNA+T+
DEBMcwZDNF4kvWgeEm5s4w7Jj+W/c6lxUFV2A2X7CZjA2XEunKxeyWJEuumJ
ATNDhZEJK7h9V1oOU7mvrBST0uNulbjiaUdrb76sitTlP9oRVg/cr4KmcKZj
rZW2m8kGKdB3JskWjuT6qP0ih0QZ709N/POQbD/IID/VoxjeTyR2R7fk0Xd6
VmaQCsaiklEOgwECg3NC5w2mOAR6XTy2pJekYTzRCkoKilDMODAaBWLy+osv
AntRISkLYnJgCbc8pIof/wapRr43RSc4irTray6CKtL9/bSW8R4Fk40fNtJu
tdiMry30OESOB7mpCgLwbgI/yFh3GLFnf1lyfhXni3YhBVJwoL3Nul1+SWLF
NAyGAEZhm0BhVHpeeeE+of7p3CSRx3lUUeccvidgjYHZW9OKb7XZn+Bcd99i
DHHBCM5Mda4LCVI2YVXOn4nsU3FuIpgnCxrGKoeEB2yp7DF61iqz5i1cp3ds
3qqNGRKsQsneaE/axdDJo0jhVfaPFS6AZMeTSx4sH+ApcuSkjtl80aN46jH4
XXR8eVMcoNS+yFWOZGOWXVD+Rw8eusP2dcMAdI0CUp5NMNRZLZR3fq20VIJv
S8er+bb6iqm01u5bL4dpd3K2+GEwcaNcN9ueWiXiqGO3+Y20SJiDo8P7TItJ
gOLuU/O16RE/gsIQ6XTCfoB/ob5jyLrkxbB/W7TyT/GGLk1Xns1LMYOjsyDN
dqpn7oKbR6HfFhK1wAdAtitBuBZZeQAr3Fx13p8IyujIGYJfB0eACrImUqtH
m0EmSIOjdNC4nSNTZnD+X4TF4tGwId1pk/zp5n7vZ1pkoHatW+6iNX9YBEFw
LfgftEHeDRAbZ8tXm1N7ETRx4o0O/RDh1uyXfnNsj83vKiBk23hJ/3gKTWy/
glGOUSJvS5V8ZTIAGaJ7EthUXfCgOrWVkIrPoiU77zMslfWIOTXCX+rcqsnd
jojhozUNXiwBwiDwg597sNaCtFXTDnZ2FUkPemyflPNG2MvvVwtU962uninn
XWwIaXvX5CyOQihQJa6+n/ZGR26VgG9lwVB/kBY5DT+NsYHgE/otiuizpCKr
beiMJRW4JvqUqEogdE/XIndQ8Cg19ItsPZtQjHTXyOSm3C96WYoCfrmRcxLZ
wUm869NKNAtkAfzxt2bxr8xQYYgpDsf6pnFeLOmBNqTCnUD6NZbEonyYUGLQ
mHtjZo23iQe1jAI8Tk3eCCezClmVJPF9SLcPn187FJsbBxd8BnTEODdsusJT
mKE9shbi43jdqtFe98GBPSg4f1fI3JVVxIR+y9uC5VntH+2kNNwdAWNKEvsI
Jc3NWV/X5YxhKYafZGYxCtX3GfG/pv5V5hv+GyqZ1w/MS1exPpBIPs2rhShY
2BwUcsr1uPgddaNYYYYnA7Ti3gF9wxZPetylyob/E7SG8d63UzfKTqUi8LGM
wqaB9lqoZlROA+OSSvaCG7Iex6Ur/5dwu7uLcPYT7x+Sah1w79WDLOCYrMBL
0IZy9Y/24hnRXh+vfwaptaG84W44w7cwA23lFH0dS+yX1rJIu6GKG8pntPob
O0LeDU5mXnCy3gyDiZ4XQgrdHmydQvBN7LRr2BJHG3c/CstxxW4PaUWIF3gZ
BGj+8hZrxVcRkRmAG8bW2JqjGAvYMb/4Q6Xe1z8yKr/R8lE4DHtoSx0MFyDj
UlhJ0Pk+uU4QAPDhrqyi0vERH4XaRpbDZROR7MoTw28bHDpRRbOS1rrjd46p
7QLQV5/3sL8+JvU4Xb+JjbE2rfrckeJFERZS+oDBKy+wkD9m/2Q4yuwhjaq/
gsjlh5ztM5rrDv20goXnHelEB52dvD1DtfJWu6v2f1WVtAOM3novz/xBA1N3
YCwnOzloeqoMsZC3vcQR+HgE7mRL7Nr/DnQ3nv/rn298WdxbTiGLqSAWAbpV
v9wCJT+BSNHalmj+aV4pKTQOFoW+7behn4x1gPwS+2iL/a5M3BFPAJY6XsAE
HCs7eJIhrk90BVeteOwxEFIsshlyiwbKSKx/o7zcgYzcPvlr4MBwaA1AxTLt
4YZjI7RlXUp7c41fz3cIehyNjvGkBS3XXcIceYvSHpiWyOMrKvmpDGxgN6Lt
bDpDxaealVNOPo/gjQ99KKp8rGonw1qjwGaV6buumoFeANBVn68uYTU6z+6/
Q8uZvUdLz+wNZUxR7X0lTdSCDWnJBidihwd/uigU11l5tz2JwAJApjuNribQ
r1t5rcuzQlZ9RiFAQLGvGe2UDCzIp7qqypSHAmuGfh32a2Vcr87vwOF2QfpV
TxRw4NJTU3zmZyROJCj+0G5zHL+WRjtYZPMZCUJSPOxWT8ncdMXI1hi9noVn
8xclvnuZjy5NKBFuPuKqHthT6fh+scxhbDiBngiwxWyS22ZmYeptwsMfqNX5
PmHjiOBMt9v5MRdtL2FDSaBELKv2cgnLjRrM3KqdKhczzobFwCHRQaE342kg
hznIHBH8Qcjojh9V5QWO9aZ0Eqm2efom0CeOvzOmPnJCFov1u5MlkvPs6MNo
VNnmTGSAXAmeSPYwG75OHSSLza03g6QsUk0KTn37b8ToveP1Pal0NbCkAi6Q
ALwe2Tnc5aFNbyw0eQ1Qi3DPdh5XXPyu8Ulny3ROnJDCMKi8+z8KBR78A51O
kOpF5+8ptP2Axw5TuXvISO29TTEqhWJzzgb5pM/IqIBlMjAQeChRABrRc3oL
sxBqvTdxfQKJ0YR7GiIbyhxtZVdRvZCTzcWkokAoDilLu58DsYPHzYGS23mx
rq16OyUtnMM4PbhJ46bAiDmSETYjBWgKXOGGA+E06Us/QFBe7RowmTTWeChj
RCXgo10kdYPUfVab4AdVP/OteWNPi6lpYWwcX/29Z4s+x3ZSD3SEG+0ddY96
1cyd0ZxFnShpQrGXEoe0Ph23HBwHEK3KjJ/UFctjw/3v7jaKgROhZQmr3Ih9
STkEfc23jMilimPgl8eLz/JcPK1xd2dXBcSjZghLvqKb/d1COL7/JO8sUoxI
eEMPJGD6WVidJAlBvOhoznrdJPKcI/XcxlrS4lNRpxjduK7RBhKgsYmOXF9E
yOQx77ohcnXXWfWMN67mmB6ZbpayR1wk48ytoCN2b4qRFvq84WP30BdUkq2c
VMHpx1eU+myl+MJmrQP9mFpZsvIa5eKVig4QeYFwqa51o5CBQQN1E/thCT6z
V/MT92G/yFpmZkPC1zi1ANyiHfcKi/T5H6X54ZEeFptWrG7Mi6d7GP/SJzHb
pzYMAU2jS27hd2ivuievlK8h4bvjr7eFM/f/58wJXN+OXb6trIY/vdzVAByg
5cxu7tgnEBhd593zYtz7SxVUtV0t/T8kTEKDqLz/NGhGeavVKKKDWc9EJKhg
WbnKCdx82me/UsQA6ZRkv3bpnYfxoerh7n2MLrFiDJrVDQxs5hxMFnvyV03i
4EYCglnkYX6Cd7IVeysWMdi8FPlu98b6yN+Txqn8lDrzTmiPBhtpWFk9wwsx
8G55QV3xHx2/nMj/cZlKuphlH/ADfABd4ZKMCVG8qM8NwOadrnUbJXYJJQIU
urHcqrtFvcxTBGKTuwVXQbR0oJQNCT0mKEHwPZVnz4weQCbkWpkAGlim3xKi
oaT3BH1tzyLyX7SWiT35+uhwTbdLIj/Ah8F7bJgsWKfguTB8VtYcyPKsrJrn
fAPpX0eEafl4d9iFbpPEeiXPS1pMlCSWKq09GHtkzp+AVLseJpvCcj3nG4Tl
AUsZGlpvcVZawzHbPSYSojJEvlg2S27RhJ3wUKgIun5oTuhv/vR3iqgES1DQ
QB+6m0HFz/Uf59EQA3BBSPwrdY9HHlAMiMFD8WbXFnknLb1AnGKHBdT+MpB4
6As0qpZcNeA/728L25k+22zPa7KQXhbuESHw23GQktB+Yk3ufeE3t2JkbOBk
hm3mgg7FQUVJPd7iBRaSjPTCCozbEJjLL/ndtCijYitUsWPl89xsi1de/hAf
LNnNwvGloYnQbAoCdtxNG8pXaQnEaUtr2K2500CLZi3AdFEG4pnXJsnf+xUd
R6CVYKMxQkpak9qrZQ5u2CDz0JPCzsfRxRQ2yzsK6BPGLud8YOev1HQfAEuj
i47Bf83ggLLL6jTH134Eu/FQ6GdoRcZ6kx9z5J2frt6M3konuqa8bPoVDZLb
KDqmppk2sGKfqV1S5u+vgRz5kHtivp4zW/9FW0giy8P/savN45cq01k5uLxM
cmn/avRCFZnSsruZrdHYusX5sc0IIFU+OxUx887zhyWBM9Kqgk5Jl9gbaFmE
IV+g+P8nLpgUFFkPVBdSyjiU2RkNwzulroNzg7aNixAA3c3RPFqVlqfG1rRZ
/h5YIqzk6DntZ2ly5k3FZTpIAqCBkMVhjoCs2a5ZxGD8kMj8xBOSycSS9tF1
j/FIjtQ0Qte0o+uOlnN4LEE7U7vFcQiDGrcSJ3qgqEy5W6DJYA+SMsro5IWZ
eLV5y9pLCgEAhk3iBIGtTh+/aM0xqDNQc1jlECRJIV0Dy35Z5ozjYMFWdxlz
EyvlpggVvsFZmshMBenKVCH8aN61FXvwCEBf1vHtzTkrschVsZMWcjfGb+4X
2D7N3U4zK+w8ZLcwne8JpP5CfKR8zarONGffK3S+4vB7ZEaBDfPVoqPdIdFn
2h7eJ0ochAupxAdIQT1uTt6f9toossKrKyeUoLeSis9Jq8FIrRd1op/OSAyT
0nxzP7fI+gHxCQwl8jCUDTxe597K22zjKACYqYX0o5zP5AOIQ9RKBksHPIJ9
qiFdigN/7c0x0i7ytzUAnNvpMdxI9X2RQ7ERwuZViw/zu26ujskc47Kf24Tt
FXtIJAd15uuvG+sDGlS1ZUkFfmlc8Wsy4mnG7IVniIeuYRHPimDQmjwcA0KP
UAIVrWjmqzblcskKguo8bDLxgQx5u6WHdn4EopPzvNJ+mUBZXr/BEgi/kCMO
Fw/UxbODFJZlezY8Dd6LvJFWSXxDQUuGIcULvMjZ10CSpxa0z9oRYdGA2mzM
gKrOvd+hD1YGNxxu1KkK83dUSEP0F/fB0bRghZ63MCvdfSKhChSrxfF69LLE
aZibN4cvuJuRmxanYZArQjCGoMYuhdVZhzqAZ28SrvFD3oj/kC9CtFXiKwB8
p2ZPQThDPirSpPd9EgRXTrJbaBg8WG+mLhBhNSi6pisX6G9TrRIyRLbVD1PE
6byGPX1SrVYKV+oOroJJKANF17cEe4/Tha7qcSghwXmE5mGZGr1yZX6If1r1
WIDTdw3uLJ67MAuRuxZ7qLLV5j3BsBwvKCyDU7Qdn35wlitni6pmnFJxHJi6
YPrzLcU74PcgwHF8DkV/mwAJ5ERkn89G6bXwaj5Z2gF1xNt2ej5V21+FTHw7
hH5sQXY/CF3OFSYgmbyoQp1y9+U1AyyYN1rQS9Eza4dc7ee5ffCO4SEND52l
+xDHJ0A/Lu8loYdqcRvn2+VoEqlD9/ASxC/zu3u3a80JyYNlshiW6uA2ALTp
9mjEZKuxY4zmKCXXVMSWEM83pizV3Mz+pps+LV3gkrvEccthDzeGZlHyBY8q
q8Xxc07RvVJStEVdZAlh/KGIPgroIGz5Zof2LujlDxVtY1Xthcx/E4lfPXw2
SLv5C1SSSl4HwgtKON2bpAz/AMwP9Zr90BMpUkDrknEeu8Ol1vP1MVkkgFfj
CbQWNqi4LKJcg7VM5tEqhV1OK19+Q6aB4G5fcPo06LUFzxkrHlXrEunAS/4d
H7B5Fsv4FoelBfYhBA+SV2w+d/9reK2il3y6Us0FYvnNiAxsR1ooFoYvL2/U
yHkDFIuOD+E5moOS38UdQUnMRiuSAGbdW0oZln6gAEfxs9OhFARhXwN3C5Is
bFvQ+jWQp1DqwFicKzE1aT+HDM3zoxfE7k2DwjN6Ik6V4flLVEr6I0bQnJWH
Wh52Psc4T2e6uESdmEejPIN5p3Yq+q6juYnhomd9NXA84+r3EVwBVNCW+eYt
Y75819pYt04So40rjSunAtYZsBn+IaBJgg7h+DyPW6rWTRzjX+LO7kQOBtPX
7d+BPoE6HHEdR4uaf/hYVnlQv0gtoq14Aj8W2u9zK3LVdLSa2SSZZKA83RlU
/CRDVx7S+/kmeKFd7SFTAdgXSeZeSrDZL/anVBFDVn5kfaxQDu/7eQQwCG3c
RMsPfed/LCw8xtMi1ZdxsBp4isCC9ll0QvyUtK7/aXPhHEkSFnBT7K/0jQ/8
BWm7lIqUygmLMUQI0gaewkYVh4UCsQyjikUpG1Gn6Tmket+MsUF/MQKVH8iB
VInnpOSze/xiE6GCyKsaUgsEaSmROBe/whvQUZRFnRAIkKHufVZXBuGYdhiR
tML2Cwz3EvuHonucRWLjNqEmo1dCNWEMAU1Tl2zJB1jKWMAUrO+VCyyZkdnW
epf66G2ESFTsjZNk0G8xfjx1N/l8GQYhsiThJnXw75lKpt7p/AN8Hz5e8Orv
fF2xEGC/mglqce/l0Sx+KINB3E8EKxv8Cw3Cuh+EsJ+3fjMGG6/D9QT8wnkq
KQKFCXeGGRXyQC0Mre08RB7I+gpNhXowySsJvsRSFh2Cotl6wCXisD5wPEyC
NK1HPgnaTckyb64nUmvKIesPGgUiR1XIapKZ5Pp4CViWVRlx8ppEyem04Ufl
rgndvj/Mzv58SsVSHSfa0U2CAHyJDh5y9VHqU5qVsXRJJbKpk8lJ70iz4W4V
Lp5paVTF3oGjpIPLEHMsX/FFHJdsUeBHUs+LIfWXwUjDQZqB+TptpvFuFqXO
f74VNCz2mqi6EAkks7ytfJuizddE1k2GE0c15dJvdgW3Xh6MvnFnWqov3hTs
Zu9/oCq+6b/A511LIfHXDp5T2voVx6y/mNFAIxAguqi9Fnx4nFmdg9tDWAWS
KwDvvhsLHOea9uw7wgD5CXmkfYyfynNUltAwT398//lK3xeYzZx/w/9gwRfF
W/QIlgJY85QJsJRkuSt+ByJShCmDZmsKXDIvmYp41bpk1Zenz/l////y9Ydi
r01n7FVDnAZP/SAkX7cef7JTx12d+BTC2U9UeQ6gm1u1bLHil302CDsIBhlY
w4L60N6dxmyRLkRLbdOuqQv+KHHcI/yVf1Gr1aDNBH8xp9xf80vywNxKqhxv
SfnQsgG+9KVTz5/pUAoDgoA4szvoClbpmQCsnIWpdBuuJmyyc/AzRsPBuypx
jra9FqeiNlIYukByL4s9dUTVNYymuBnsjb2FRKc2aYeoobJSaUsFCl3F9Oit
NVneXVs3U/dRkyiG0x76c7//ZyPKe+gj6KTpm2jk3ZOQWYqzwUBjwg8Pz9OH
U3cjl0/1kEyqODy84lw4IqHHEnOVES1Eurgsuvo49pSu0dTk0wBcU/YTis7C
/s3q4g6+F5pG+bsFi1sRaofYjMdQi+OX61dxsd4BbNI0wW9elE30ENp+BsPD
pbnpIPRTDBd/NmolwC3B+q9RHXPux1ye/PwOIGYWRiKUHd9YdO8R+vJVvKhf
kVeV9Nq5bwhD7py4kSYxHbt9NN56ze/Yhdl358Ttje2td+Urcsgr/Iw1C2x2
XgP4JQzQjVOxdZmCDjv3wDwBkCqySAn9ki2rNcQ0AdPHINeOCo8JYjkpb39m
yhOl5m5JqQwwyJMZr/OsVmV/82vtvhQqho0bgWK4LsmzHR6483k7qH7hJPt6
+HiKF7pKb03OPxYkikrraqTcq76L79bxoA+vCm+2CfJuZ/fOl2af58pYhlnZ
338pjBY7pZRxxcfW582gWuhfbToB8yyYeA2PbdNwJ/XvhnFhbIroTNkiSRQe
M9AkDIZ6hxOqcAHra7XOZZaTTtBCaFSPGN+29vHUPokZrSkePvfKunq4Xi6a
Dck1nfjn4RKmqwiR0IFo2MxAzBcqzlf1ra6lPGJG1We6fyrT1jZd4a+ZwPmx
pN0cf0ibHh2N2nTAVD3o7uWV4kbVipEynelI6U61SqA9n6wVNm9WPtaU62I2
vck6ISykLJ5XPc3wQyOv3/RMwEig5OyVh0/PLQUbeoVp4H8KTDfGPSe2VzdY
74UJvLDH9tGEe8F+2gsNpG7yWRusVZwwNHqzPLmlFwmCfDjbWS5sw+3Xsp/u
LvEG2Y0vy+iBriqeD2zVPxQwcHQJVWrLkAh6ld+Sr74mQqgxhpc99rdkvHiR
fjYz7AH0Ezyxl3H9zy5PDk5CZ+y3jlRjNUutZaINyUeFWDtqE3jXNhBv4+SE
oXMBS+MJak76eSwI1sZNQyQGaD5oITehGfRQ7W3G4PmKzLaLKTE6BhHMAl+u
YNSU4xfEcKacSiiIoBm0v5sFx8B2VZXgqmJjSr29uQdDr1OFX7Qx1sZZNGp8
iRdeIgiQrsHtoEdmgGdLDTtLzfYaLS0OxLepMRAi0JAxERnIjaHBx0zZ2R2m
/84LnG8N9OV1uJi7F8b0e/IMpenF+liKBPs+4hbCWfJw3AZ0HLdS0cd8KADH
KMqgHLfNOej3hivJqkrntFpO/MJzslo0F9cAEIkhlqvahb/Ncx7LgeevfQaK
UXY2Y39TYpf1NFXwIrY3komSJHTxtySYyeMgLKMCADv8wlyjdnUMnieo+miO
EZ5ZalucdkpEAqipNwkKHTCrGAPtCKx+kIZEe+BDbktCR2Qk+28t0Bv7NBD0
xMfancOa5d+ava2+41cXrqNRr/nQAhDy13k3D4YVUeEtzlklSJyalLI302d2
x5XQSNYfy8ePw4GG9WmC5hmK2rSIuQqE5ulwcUe+a0IFzz2dKyznmdXGlg3s
g+9pBMKHB47zrE5Q/YdS2FWh/GgxEWfKcfdYQHtbN5Xwd/BYckTEhH8cYMTh
KWERJzSVwFxLhm/HHayBfhDjx4bXpU0tluLjdNEjI+hXUXM1D1sZ14XhJgIH
fdXAjI8vVmPZzCKttWitqURwtu7fYTVW+1mCkst7aIHrWvjT7K9O/3P9w0hw
W9XqNpCEJ2ehWrpURhlCFFROJJgg0Lx3AZHpgzU45s0dDo2ngHb80QE4TWI9
HQ7U37q7mHWET8hp7xhlt9BG0DPKxufOoBqSZ6SAFCuWvJKQR3xbTfWmBjkz
cBFq81Xln994gfCqzs7qChJdQ8EiemdmWxyEOoXqE4ysF0g7ouOxjACGtqOp
nEW86m61gPSA7MIYwMbVbmLmXDnLC36rYTCbhw+pUQtIZCXqVGih56/jqUCy
NoXteIBUCdyrh0DfNeJazH+o9OJ+rff24VnGbOd3gGlc3gIqGL8Arwbz0GxD
FJ0KavetsVEQMcSA0HE13unl59Xelt1wC3gbiRceKYIOKpM167XOeltInjfj
j4oE4vUIoxTYxi8hU+xOVHjHsbBrwYthTwSrut+SWCE0a1Poecqm+ufNrdte
0TanGl0Sv10U5U9AV2mhL+tsafLIhjzF1LlENVkzAgzjVrvVfcOd26jGEtma
eGXFjPpDOLneIR8HdXLc81fvDJ/+fI+1mix9r3wkkEcR8LiVOBCz4p6ZEoAB
P9H9KqgNog+K3Lph6W8DzygU8tjzxqocpeevk6aDZvVdD3ly9FlGHXLdfbX9
+hSkLYq0oJVZDuOgyz71ZG31lmZFP8toYK8fF75RzVzVsNpGuJeP3CYZwumG
cc7AmcaPg+8LF62cnH4Hh5pR0kHqsMi1xmMKrFJjv9Sxe5eEPh4vygOkRwxV
Ic5Z7VYUGdnlcYGx7TrBmntOzhzewLQj+36ODPZ1SOAUhqUt/Y4gpLzwM/GN
NOMZU/yvUVVuhEdaVzDvn/h76D3fdlk2mjm8mdACGXeb3+/SHruJV3pJOSpA
aT2RIHzVIn/NCKxhoXVFR2V0mPAYhnkRPH3yMtik2iJlnAcpNHFl5VnRlv5u
NloesmVbVrGlNRWd+o6uLimGe+fuHIEV5L2J0s3LgjpgmUUlV0VO3HM0i2JJ
Y/HstDoxuOnz5awoQZx+8YqPD1Gh3waOvu74//t4NW1jNRY9z1LPz1SbhEGd
BgnMYSjTIaI3YmmtR0IH58EkSVEZNIZbYtD1NFIqy/hFn1uz56/Ds5xkJ8zJ
8vm6O2PVdI/uRw9dCdgZAYB9bTA86jOukxbUofC52EqmxnVbeJD5Om0BHg8v
c9CHpM29MkH8EGs3fwGxMQfLqR/UYSoAFf0oiOwjTTRsoUDKLlP0njwoUDbS
5PCyokzDT+gSU9OovjvzVrVYBGmmeLkX8UYqF12xn1l2T3KJ7Ki4++wj8yFm
AOHvHd7AD99+IcV8n1i0vCClmclcBCgd9+W9AjuvfI/1U3eP0gqreCXHw3s6
Lbv/u2OE9Cs4p+aypRKEIJce3tS+Ri30etpSn7QgY/SRX0ECChyat6SchLaM
b+hqqkFz0RZWcug7FIxjqSQMONJLM7KTUQTIRXe7mqOLlf9lqHJdbOQkqaK1
M8L+kbRVDENY9of3X3kQfSnf71yFj7Ic9smuOBDJa0ixF8vJGadUfmrPzNMH
k7OFrH+wBdr7lfdYe9XzW1x1uQ7MjNfqS0palkrrXeJfTOOADvLdfvHGmCUk
WS7QKEEHZKwA6AolqmxhQqMYgS0jyJg/IJFcXIu0nUFmNF4T5n4B1ykCPvYv
XFfc04VPjVEKZqTpXevb2T48rZmxfMAkA+z5vPOC5G6z9pJfWTaeKh8DsgPh
6nA12hC1esgFAsB/nyewXWEHi7vjz6iAI4QN7RIEVvc2fKg4+Z7gRVZqjmOq
JQg7iA3n6/IUXf9FX6IDLEtykqG6SPEZP93kRXEXhLEUd+WJzIPHLCS7pgGo
gpT4yvO2w/p7t3K9N+2RFit2ohiz6i8/o9cNE7T054wc8Oq1h9I8IAQJLmA/
qe3vys34TTGytWQrNQngOozugzPHENOgp643DHriWxit9ayFbgXxYun20AAA
abk7KCiLyRr93fUhLr/jEgDNoT0rL0B/TkpaXNoAnq57u06L7M75mKhSxg5v
So7N+n0GEqqIiNJZpYrL+GI46pMjD67K8nlM64SOuXAXzGeRMH4qcNge1u6c
g+tq8qHjpLA/JfGOpePbk6l9jol83fso8vcTHeVewvaR5qjIAa+QaQval2Xf
7yqRP/PgaSuO6jDRI7UfqSpjAWcUC/hTd2ChpYKqvOjbHFGSiI3HHUYGn3GT
wrgYXxFChlqJd5spiyWAf2jv5/Pd5KXJ0Cgmrc0+qdkloYN79NNgj+m5qZQA
hBNmkoqUcc3jGik5I4H3JgfHSqSJHH8nv6rkiDF7MbDIVSWEJGknX/bpdgZT
5sy/ehCsgcDjWvAbyl035BXgWoL+ESftoGd0WGKFRL7FGPoVTILrn9jNniZY
JzyyrNVnQb0zcOs/UNb7OM5Op9V6vGF6mHhX9tjC3PvHhJENhIkylP+J8T7P
rrzd1/U4+tQcMCn2wYxe7xpFcrHBMeaM6BqgYsP1OgQIcGmxrVFaqNCgiwe7
Fr5xJdTyfea84fZf4DCsNm7QvCONHVV/leNM6QI8ViyDi4Gokz+WA19uqi21
zrVkdPkNsCsZpwfBZR4bAAS7L4A+9e0fSz3HmA1X9b5uurRbWk7gL31CaQfx
nlYGf85yZzPwz5yoXrzqbX5cM2rBR0xVdv/x8WTBNs/T0Omu4eivg/yFYmaN
4iF7JhqYAX6CSIP4VMFhiPj7pGTwNsAiJ22yfYQjIqnTnv7J2ym+zHm2zcke
M/uM5y21t6+bq3gl1P8Sw/hTABsq5pMUPfAGIWKeZ0BZa8hzsF0RgdIBzHWY
TSF+ABj1A3+CAAZhxWkFUVceM8ZgYGyFse9hEFiKlenxEutLhPVC+Drpv3wq
ylIKq+GTm5oSvynHfR8xjLAjum1goAYmzlkXIUUgzLiqxKTJg8d6bpiB/x5j
04slfEcut+axK0y4D7+mJRikXV8ikhlLSYP7PNt+k+P4lJabupjoH9oIIFWG
6QdgbkOVlbVBgAr0mO6hlUWV/hHNnD6lQLKkQBZsrCEIgoqxxverfxY7O7qu
Wdyrn9WOfRWPKMSo8zNWSca+757kWC3tv/jX1+7kj/DCVKWGvplqsv9huQ5N
9wKt07GQXNwxfA17k6PTj6f6OqWzgzfjvV7qvq+cJduVcAHczsKt6TMkjB5w
rpLZmm1YYlEFnyAdhZ+IAjKXix5oM5T9NZVo926i09GFiyt/6Jta5EFaWE9h
3vP3g2sZMVHiyw6tZi/GL1kuL5lYch9IBpBZOZd82z90foCd8mjsoqPHQJz3
5pwN38Osh/z50hOc6HTYF3BiwopOF5Yq4L8SuWYxW+ERBcAslBkUZkodMWmp
olHu9za1xWfT3FoF6NOziI1OkN1iXRxoLpvPr/afnqBdxgIuTmuyhCXSRyPJ
LDGxdyiqK80tEJQnl0YT006y69935Pg0yqUdKbkjB5wNcbVMGBSSnvDlMDn4
YqcgxtsXj6j2k43BX4/GJ1yvQOr3BOlpKVKgYXR4XmgpYzYY/u8cpKGNzO9p
H3SuZEF0RPUb7EZzw+NOd3YcJVrNcnjikybCQtrScSgVhcEXsOBfqr86wMqj
W5/W+uzyO1373OH0hPkPQwqUX4TxLI5hHwXcfOcepyWYJq3i039eNDchBcUv
JXw+V6ID/LZRaWQ8g//ehzMR1RjfBS7HjmxodzXiyJm+2yfGzTMwVpS/Ndik
E0ztlFZ/7b7BtuYwPANqLkjisktQFaIh5EZM2FNcFDxgUFTBe9d+Lf4foSWt
/F5eDHdl1mKpkHjeLRFafGpt566R65Q7e6GhTBX3FWEQrjxwBcBq6lSJi+zw
xKcCUaMMxNUHQbJJKj7mCXqo2f/e5ZWAvrBoZkocLmzMJNEVk6Fd37RQSyP5
kp+GvkMkmx9nBv9s2EznU5sHjNAx/iz5R/5Yk3ClpHlGyim+N02SHgPFeDvk
r5Zs0ErAUQAa3OqEfPCZg50uHdJVnS1yA4Gy/xpTVhh0MFqiDg8NQJ1mtttc
70xnx82WYLe1uD8k4jMhYnc+DkxERD1r5Tiee7ELJJf6JqAn5aeJN7r5EHvT
54C2CsoJrQc2lC+QnGnjw7b1m9pkSd7bP9+lUWak+UplOAw6fQplKbXzvzIO
o/lRn+JqQkIlNUdztYHp2rX8EXolAmq2DHBIV8RTYq+YhOXIVyGtTJnimkTu
AoxKgxcfAQWAIjjmGYnJVtP8IH9z8ffzg5O2/sGr3btz+d2zEkQb/RV3Fg6O
9j8GGaEQZWVCDRrVJfsEaFTJW0hQqqI6eFTY28w82fZmUiIYg+tk++15/uvK
ReaL4eh9aqdSiR+9fCxJVlJba9ZBNZVJrOt6hv4vpoAigBR/w5XHd3T8+ujU
4dWZku2XHc/tQx7ht9SzfD9r8dfOkPcAaIlNPfXW1r8eqjgsPWkXnZzZcZBj
hMy8/SgjJmoI2rAyh1KjxADaDB3PV6QKoH/ed0ROHDdADSZMPCFBFdHOM5Ht
57Um3jp72K4LM3uXBSk2mlvB2BtBxzeAaZvHq6vCdg1l5yjOahd0b5Hz5HFF
ACLvIaq1m752yLTrJpULWFq6Y5vmMWauzRGgTRQeZKIbvS4+Npun1qavGKUL
bepErrP4R+Pm51tyH83lpSi2FRESY4j7a4eIGb/vNldpkZbznxDFTNXCxFcS
dceD0bNsW4wKPpp7azQ3T5SxAqFqybc/wxfmkVv6p5zaw+raQuWZgfLO6WEN
DZaCDq2d5Bbwal4ZGeS+iN6G9dRUe8gAAiPkivMMf6xdbrVxM1hPdZzLCpld
EQ+V4VSVzmTJ/CNYBXMVRQBM9DIhvchBQaIvzpM8N5peK2aIjeG1MptOe+/K
8ZteqVJgdkqtWxlNW5UUdLMoZDyj/+QnWBc3vug3zYXMRhrp85VMBuKPY6nS
VOClIwft6WDkF1s9Wh8zVwUy+Ua9XmRFxd3SqfEvT9oh2KRb+xAMYssioq8d
GyWVN9/EucSbNiKdKkYnSuy9MnHtAIk0QDbknPDuAq2Q999UNJOajF69UES2
zK3K6J709FjtoneyEtfrrNR3toeav6+Cq61I6oykuTKcX56CK3qLO2E6+AkD
940Vlqh8k+3MqM2rqtiWvyr4xODkG4xh5nsRmvK7E9nvqj7aCLgkoOS6QyWe
2oGUaj9tG5JD2wc0dezyMxYlyOqrWQ9aaqoSP+zXzC0NboqX4BQNe/ewJ5Mf
wixH3Ef/Dh1lHosyUHuISz8ahHR3q88CtYCk81MAzMG3VXvmL1lsiuTR5GIF
StrgyhPmp4Cz55RYD0jtFlRz+L95WjbOleBe2bVLMNsWJxXD8+UzewLnSkUZ
QXCCb3pTVWG9czbjH1VIjVxJovPtwHJ1gDdlXGrqmmx2sFZ378F/HWmdMcOD
GCmLt+sDI3HL770uwc9SBuy8P7ioFWCJzS4s5orOrHxMLXtueuEXDVpe6FwG
dLYpjctrBDxTqmPpbls3ftpHZIOZoHL1SNd+mVwoxmzmBcO6S47PhL3kTlpe
Q11dVm+JVcNyxsWNRabCLfS8f9GzXdOT+AlQTjIAK2OiLdTeaElZDBKuT2GP
77Ar31SWJDsqdYvI8PF2OcyXEqJ8nt996URSuSo5MSsYRgVL+cSHpS6v0MgE
HE2yvT7MMvKWWATOC1AMVVUYV/QjvXSK13SNWJdSf7ZEiDS8xlrJlBmokESZ
YP8RZ364QjqusSc6FSzCmFySlj5tqC2by0YTrCswVFlWZ3wT6J1jT1iyJqe7
hFWW76GelGbYCQNvkb9sOO1if5D1F/N1S2qBCSjEQ/0qOSWsRx/+9ycwEMXP
lbuSKy5tq9wUuKM2xTHDQmMyYlg/uPFYV0SWJIcI9Thuy9XaI+rWBGVe0pAZ
tYn2WA1vPqk2jeRqgAXMtfktJd7vGdF5c45CxHu8TQ6r9CGyAoLXhZp9o4a4
RTMejwA/+MLMHI38Wocn1NOJ0kkxJkuN8s5l4F2Sbu3YO0NQBxZRtBNRlyBW
elQ64VA7E0aPpjS69Ld0+wqCCqUy1uDIl5VdpTYrfMX+xr9+UB/cs1HMdULH
UU9lZ+aVgXyIoVR3tuLQY3X33YKN4KOgqVu3FK3U3xE2CANGY9dcHbfFxw/L
BxvhZWcwDpENk4KjlhYmQd48PfdV6qfRtNYKfXvYZnyK/ofNVwiSrQUYRGPG
S9VojwC7zdTuHBWtjmuj7GIxtTZcbKaYQ6539tbPbfySPPR3GMU7sOf8VFw2
gKFxGsc1v2tURRH9rry6Yndc8HoDrinuhQlakfbPRdwHcFVK8uyjS4dVnjm9
LgvdeISpPv69+ttQAFWm983pw8IoTt6qfcIb2uxofO90DBTecpEGNcOK3gtF
/2G36BA7UoBEtGPCubwEMxeacRI1tzw1HVdProURybBEoZxZc09gEb71hmWx
2V5U4BGfVjZUOTn0Vr8NnuH3L/MI9IGlerpLFzJjtQFBNIKbHovw8Jadsxk2
aY1ObyNO6Lvtadq9f9Ssf43yumZOjkLO+HtTQjQPw4tk7CfoEkmBL+LUnJsE
4784IWb8v2LLCTT56Tg1aJiUaU2QI/soND2CYdmudLMVeZNh2FNBv85RDGFI
fBLLabbsXqZH/R2lC/lOUT4i+5Ffr3a9t7FhrudmaSoqrjsoRoj+kg9EsPZO
kCt6mnpaLC2OOqD99MYt/Gf2XmYxSiI3uCAoAC8cLvNmtPM3nOJZXRoIZ9e1
XxJ9JAIfhMn2NGbZLpBC/HXMZLtKftEhCzW/X4aw7rGF6/m3R102GI3Qs6D/
/Zo9/4LulhnQzMUf33p4p3McfNG44N9cmF4lEAW+ShDS4sKBcY34cOkrTcIz
gpoR+KPammvDEHlJor7YEylr4+HW97snkR8Dpqw8GAV041+JUJ5NRnhHzGA7
ZAxuKhW81KDLpBtg8966CeJ5nmekAaP4yS+mDkP3cIzgXHFYlyN9bMouFvZx
IL2+EG9rWcz5/omWj9CHthYOLMrQ4zABUREsFixys5EgfPtjuoVMBtnMDC/E
ydc9S7FDh6CZp9QQ2wNusQEfwzJbCEXlaLzb3EqABy59rJPLxIaHxJIHvNLR
IkSm0XpIL7bYBHOHQ/liQQ2tDEqGvV9WqCdjsG508kVFCUk3zo+JWlcjXqli
Wvyb495tH3BwQXHVMjGqZuF6lIEumghbXmQjZ/M99PCMMpbt/Pl3ijaTsU5G
84ru9PySpFEePn1LQqOr+LsKIFleDSo3i1XsxuTCmhdKq5VK9BWrW0ONql0V
Alfdg3C4rx1w/hRDg0T4biPiqs7R86HiEBXd70bugMGrpA80RPlFC9lXVgGt
qS5TGlTcdvyZ3pvOrO68kPF9W4l+YtUVjDaOUzYzVNDchM1tjkrP6f2t92yt
VmpT22UVcEKb84FBWqlmspPO2XtFm/wBzKjRMeppLSzV12OYkZzFK+TMbfdD
6b8Fa3/g9xo7njrV/0sqSblGNyF0QsQZ7KW29zhqStn4bFamnSrpmodvTbuE
GNKOxnOnnp/uZd3gPw6JZB3gXWvoPs6BlfFs0Woi0qs3dJDptHd4tIBEhsxS
VfDazPcHwVFR6dChS2d0qjB22hqC/Uw4rK0c2EswikJ4uXTxHxknKVQNDPL9
eMd2QULH4bbDNuBpCK/bvCF8LkMM90iz412A3Ln21D0kp6umDSlIBi1EVvFh
ojqOavZWVSjeULQ1viGjDbGjEs7CFA9lGG7mQxBiQ0Et2YhsDAoNoJtDq5sU
MDrjq64oKK+SZFiLiPY0mlNQndQ5yZCLfeOkC7pdJmIP0Us3fGgtiCOv1704
lL3mAXHuSPj8SlzujwvJsTyG5IX/yEF/eir+vvdnpt85Xaj4mAvM0zrJifhh
phYkOQ/26olVVYx72fiBcGZ3hE2gCeNlY2CsGDCjQRQkvlOQg8DLdVJ4/btX
0Nh6Vdq3ByF4Va8s25tJ2lVCOcn/00uhnmdRVJD6Dr4D7dRREoM2QW2+F9fS
rAPuOtYBzMOEbw8suXxw8d1GsxC2jFghOiVTQgJt7hJGmAz7300GXtceimX8
ewFqGL9uT/dC08QGdU5F2Wn/FV0LEeqAtlGoNcS/1MBThPUqylXigZGpI2k2
0qlrjMgPZL/OhXsIuNeH7U8IHVLAr0TfI3gayaXRSRQkFL1vaRWJVMmEDDrA
ZQqVPV94azNCgsCV+7MzeIh7FfbSswWpW+8As2cabSLZqwQ1SjNR9sCaU3Xi
AeqO20MEziWXoPSO2sxLJDY7t69tnDLnptBhsAXirsvP/LiisIKX2st+y803
X12PFLOLA2QkGlu//SWYeWrp201THuMjwfug61bFywFSV68gBLKADBgLf8oS
Yz3kJn6gxPhyWLbwfB3BLcE1CS5a6y7ZcqXo4um69ub52xIqo6PnlJU/nFeU
Ny7Kksm7urJw452cmIJCtJLeA6q+0e8e6BtsvKSJzA243qfN/2VoYwLam55t
oKa/Crmw5Dmf9qAuWzHIhJ5C8C41mEtkjbGDXCQjN7gBF0lUUmZnBfe9o53t
dBrvD/XZbCy4IqJ4LTYl9/oatYdNBcDYaqWh1SbKePWLThChNXo8kXk38HUT
WqWO5L5r0TOPtljwKaJPDI8y5g8hAZto+ArOiTXF/IC+GHqlHMt5q4V0zKwK
8Jw6kInRLl/1ltp0H9tACNfZs/ZciLl4qz42C8X5dAIaV3HcszXLsv24J4C6
ZDqY5E2ydQJHiXO4j3WMovo44BJ2hquAlk9hwJik92r8bJwd0mnHPfk9gJKX
WMQzsE44dTQ3XWlGqM6zAYPpMlit4F7BSr68D98SoFyr5vfGwAsiIoPjl2Zd
K7AdXkyq6NN22EXpK441StxfkPH0uHffyy8sX9+3AZS3VpGuKzwy/zbaajgx
EFCr2uV6gKMLjNpSD98SoxvcSGkr3bZpnrv9weciw8pvDazlKq3rNVHLnF1I
5hd2jIegpS2fv4A6eWP1cJcaPCdAObpl6Do9nqpcxxqtS5ECuBh5Nohb0YWp
VcP4Su6W1wXbcpeZLnh6bo5XHA8tPN0tqj7IDFUDZv1UoX/0pX0bHnQrERJA
T/idVRbDmtbaYidEkFj985+ZGYdtla/bKDQHWa8hXfZgNacT9nYegqZnOqA3
ysbcCyIuSawNpuTfijtiqnzYMcpFbq6MjEdn8Lt0HFDbAh0IeeGKEWuli3WP
Ic8JWynuTpqcqWDPbecB8KXNtmqpOM6wwN+z3qk3hpcB7UleVAToHu86vDBc
C6n3nKNj7JLicuYwLsXjl6YXc+pnjN21HOpBTYCYxNikzKzbpkqPAtPtkQn9
NDcecIhueFZGXteo5Im+bKwujFmgH/Dr8S9sMiebuAHn4RXW8Kw+wsv8lm21
wFCYvnnLm0NNYR1Daq1d86JN195Ul9R1GCittC3D8Yq5uAxGgGebx4riZ418
pWW14l/4mSo8aM2zqhUAQ3O4J9WujvhAKBPZ60hfxPa0dWBdTwmdfbBLAOAZ
G7Xpy/O6Z0tSKIwioIN1stZqqGj4c49War4siNkrGrqRLhE+3qy1Bu/wqSA8
F4ajTaTW/0lqYlwn+L4PJ7Z/jKbvB2QnZRNmZeLmT270xQk6wfPwagK7phh7
RuWK91r4mWNRZN+YAr8vZ1LcypkWbq3vRG5QSIMy4Qbh6sYGUSNQyUKF+hOV
6cIdF3z6bV4WO6BFsf9BQTQiYa7SrCclnt4d1tmcgM3eOrJg5uMs32aGlZRN
UBeqgnfmX2ILUjg0wiokgaisG3XA/iV2MmKEk5iGowIQNYkjDtx907EAyNoB
yX1CMUcfON7Gi8Mm0NWU3ZxhFjVGH00GOdatNSY/tbRP1hKa+B/8ZEiBgI54
Rj2teCv17pAhkGt9x8wHvnYr0aE6BdxMMStXfXNLxaKXgCeGUUNZaqAmZDJj
MKaRQpCuq8myik8BDA7UIqyIUFQS/CekKDFBxMsn5zKLlqNozgdlVtZLZOec
lZi+Fzba9p8Ggd1m9c01N8fh798UQ+je5VsQa5qmD+kH7pFTcuZ3pv8jD6jg
1D9cKN04pdWbc1kQZqvri0gMU3gcQ1G1C9N0s2Eai7hDNs7o0+HJcLBfnrqL
zNcMUCnCnHuLXXTJf24n8y3V3FPjxiH4QMzNyEPBzJW9MlTNCkidn211FE4U
PzvjBnGdhgH4RT3Gkrk/b2OZHjjusjUxU+UEhuaC1eJC1F2ABtEwcHsTjaHS
1NfBi+adINM0OEV3RHmHGZUOJ7OKBU4+NUL+oSYFbzAqX7k0vxNiudqbf4yP
gmYeLz5yFKjVe6+XZrbiuuzZRNWBvbr19t7mJxzHO8OyYFC6cbgOfFE1LbPa
wWxx0ldeSvRPZIHo1WOXEdwq4jZOKXOxlF4v3yvK33vzJJzE+/gdAilxLk1P
HeB1Rp33NQjzUeFxlBuaGBxnaGgyzcgH6QVdik/gpp3Ybkm9zTNCAIShrHcC
uES6sWoPB26p0N6+0hDXPAh1T7T63FG/I1cIPZJlc4KpO1rRD/aKaZF3L0zu
QNIJt1WHUGIFG8wdEV5r+IrDagNFEdX09nGR6BILrOfgltvOpy7ibQ8//2ON
TUJ9g4b8K7YC3T5m3Xv4WbDaPd8GPFNBiZSfCypizxtZaDDTfTWBaEZoE7wz
W5hhv+ymHxdsQg0pJ2FaCBO6moszTXUDjB9ZZeu3yJ6V/vYRr3VvGPtJtXn/
dEKfRGvh3qrrojQpOeDWq7TQoEo4NBOeIan3vI86LsLBAIEas81YbmdLVkqc
fkqr3eMXXRZ8k7giRme4UoXERf9xzg+U4yaYulOEah3GHvdjGG99OszdbNA9
x0ESsNjY2GvWFYUgvj6H2XzZRfnNOnRqKaotdbOq3syDR2EuKHJBP9wJPbAy
piRz+VjnD83hqbQT9tLpKCJ+KZ0ceCh5rtpQKbcjMAM3g5ZCJ8xcn9fZCDhr
vh4lwFqZPrG1mXkLFVKcUAHO03KQQyHbLkGt9FNTiP4DnG52LNM4E0wp+Wq6
OZoHTucWYCyq496bCpc33b4D5Dip1RCzLdpM9rYwf5uUxIGC1FueHLpoMkhq
GwPgr4KfCjvzHQGxJce8ezMpKu46xHDckqFouRIEmu+Iabr/fW4hAa2rDpRu
OTXTFwktGuVE81O4IkzBI7KuVErRxXRRB32PnUec6NKCQanyBZXh1QL27DC9
aLd8H43+1jHzYUd8QA+TUghBg6zAHBSMGyEM2TQY+rvojJ2Jk5WTYJlpILBY
BuOKXfSQILvtWbXMxCMoYC1JuKI1vXMSTujUbunCO/J9EtMvFK3qrrNeBRc8
Ns6cVcKa9t2KgtAE64QufMVs4cnO4x6L5HBhkf7e3Ep1ces1S4KyWlbpHk9Q
vkHRw5cZNcyVlIfieKFB9D6qI8l15CpBw/8lPfd27RjczkL05H+ORsmHgAWb
SsvcTVzSN38atQy0MAmczntE35oOmHF+nMAb2M9Duz/iOqRs9auFz/lNeIGu
aG8jCK6QRXSf4rZTlFCUavknUfZe5c0a/khSnbHB8I/4g/2seBIRGOSAQYF7
wQFDT/Z408MOnQJiANHoT6GCd6yiOBJ1MeeixowRaS3hHjQX3G11Z2dGy5Yl
3egF2/kePODp9vN2ffXPiVgqr4tJMe1y5pNwV1ipa2SWDcqdOOAOi38uljNI
wQqgQwaPwtVkFwf0h1obA3UAEr9UdgY5A1KegvcYF0a2nZvQblIRQOFE4xGq
VA032TnE8tO7w/QJbWDr/cQ99G9siHCCw9TNZ8YSEc35yW9TPk4BV9jzASC/
1mC/3WWb+bIcI0n4d5Xa5ljczF323vbSiTeSq7qwkIlaXCgb95jaEfAqvGdO
+u3nuEu76zptKAdSUSOX2GfSpbUH1hpSDm0MR2yO/XxxJRuRh5Cw3VbC/WOs
FRDaQ+nKxHlk1TtAeDYVSoJY9w32DvXH35UpyDxAUed474X12+Veh3ZWtLqK
tpUw3CRXmUla5Ae5WAAIoypCXsU2bieU2NKtUj4SAPrg2Qhptp/InoLaBRDs
xILAZTMc9eaOiP/LSMpNNEPHqSaEMEu+Ywg7g3hartjDrUVCUOggyGoWOuX5
sEcx8bIcgZ6EjjLd69vdFZjtXEGGvs/YyOj5X72DyDsxTZ0PsSHBVZJPBj74
nPlSNPwsi4z25RJEQWSoVF8nqrrvFs+KCqEDOAV5ipFu/LcXT0IVc7cFetqk
SNypiV1ZQsvtGKEAc2o8Eni/W7tTEYByo/ckCSYGaqK7JWzQnzGNgNbrPEEQ
JSE7/IoXt+bE0Py4WW18qCMgejohzSVC8C4E9D9p80GOb58gqcJz2luVfnhD
W2pOP2x1khDHke+p95L4JTbdTaq2fEUUzGjAIf/RyJoKh+Oe/TZ/fH6BenpN
SK2OS3yIO5nPo62BP+13cYscbD5TiAFdzlacPiNWsD4PQtRrMMFa8IpzHQzB
1QjKclPZsl4s5wwpLAJq+qyJk1aTE2j1PkaXsgnP/WGbb6uWSB5Lwb51Ym0z
zfr8grdrgBL4dJanQLS6BHUjt8LPabeWHQ1lMDWNaUNKjcKwvGYoF5tgyZ+K
Dj/Y5ti1PICUMWsG2lj/3rLlnFSBuzJgfzFrshIbyAchLODB/mvc7+TVS7jy
aFNvZYZomJCt4W1AL+TTPlqMuqJhgy3BuQE+X0r2mGg0s8GgNUMjF8VoVHV6
tW2Esdk//FbMosjOWNIUVpRex63rH08Mm1RZUHlmd4z350/sk+tPms0j5RC7
HlgNe5CP4n2f/IXLuUDjrSz8B7i1MjKYYpkKCDVS/lzOxXPLvLw7Fz/w7yC5
anDV0edVdd/GnZ5NqAvUdQDCC83ZSRuhfzthLan968XGE0r44vByjgoA/JkR
4MN5ECgiuXD/vAYJP6hN0rSER3AhIM/J7cuErlCMTVGAnqBSUipTfwyUqM8R
6jhu8MooYEjKiFlrdVCEoUA7tR9sd+6AbeDd1rvlaGjaqla8HVzGcOMFGjuB
jhtaiLNQbEvSuKMIP7/pVDLZyu5WQXu8X5ZMtV5s++r+7np87co8At2N956/
Nhuz8ptTEd6WS+5Z4cyfKJx/nPP0I92mgFjVJRAOOgxjWXjFuuvaNE4LHR0c
Usvhs7rxuJ2UQaIQm3tswIzpTrPBUeNsaJKTy0V52f5UM0r+QZPmZnjET8Do
FPlH7pK6f9LYqeeeVqQsadSPqtfdoKu6Gvxd/x6i6tdrxJJTuoBczyeFbJNj
xNZCzjrkNnoHX4LB67nSat/G06Z6i1pDH0mGnjnkWu2Uea9Q24ZR0A7RVvA7
bnMJF7QYo2GyAPtdBWBBHg57A5UQ4VvYwTdOFDVhD7HaDjrL1Kqx3H7npNOK
9pIKSJ6ZvcQDe6jIkDssBa/hV7l/7w2ZVgViAY/lgukTMljUGm/PfGdETHXo
9goBd2janFuKffo7JOGZwLag0f56hnoFVIxbR8W4KmM9WGOOazK/xE+RhOiP
D13Zqp88+rcINIPW9xjSsED++tuczXC8C3BShDXB0aWoAm7GgmpLuQQnaURB
FkBHfX20fzGQZv9v92PFZ0HT1tFW6Yu0I86neXMszmfNKrVvcSSY7iUjlRxA
jdOwIbo9zRCa94ZjT8wFFjb4my4SN+anrTnLlS6wOtHc5PSG3J/X/tjColGK
s0KGU7FbNMM70IelQNFaIJxh/qSVmWV8ZSWPKAcT03/hW0gk4OIrGKMURZFt
FtlxBQY2wAhvYj5qHlOHWqyy2Os279jjgIdsLn+UqueDA9A/TYe8uDNdMrdX
SRaqZ+lE9N0Nue2Jg0Y6PsZwt6TtjYLBnYolBo6veDXR48bwQJyru3Onam6l
1DUAMA0BUCZQY0ZnMGZYYvTx9Ro+0hLV+18lHqNDQ15EMEezqfQO4buFpghK
KhDbdlsXbNvP/Dz4ICYcyW69pYxRLWe8tdtBJsTjn/41G2m16PB1wpnsCJRT
H9+ThNbUviNfE2rDD6lFiqmcEBlvgRBw6Hda1uTkxznFArG4SzwQDU1Q71t5
IyGZSfm/+s14YhGP6afdd4+YbhMNssn7ewfjwN46RpIIWZUF/q2FMuFhuWu4
7ABmPJCkmJQlCVFSyuTBZDj2qQj1lSSTWx/V3UELMG+tbsUurqviZHJLoVFJ
m+V5L9zIpoqjV9LC6Lxv9v/B4Oo3ffucGhdBaRnEQDqDai3ZVrFdyQEFlYo0
GwV1GXCiLMQTGodGGisbPUXSHCKPW3g/KWI4xYwWDfhrjZMOmjdCu9BD+PI4
v08nCohsgpwR9gVi/9/R/Jch0O9OEI0Em+oj4wTEzGcPAVvRlYDtHppUYKDP
+RZ/S1eUGuSsJnKg026SyGa7ISLxd27PX3pC2kG1LDq2yM96i+xF/CG7/ppQ
mUBeIbLrvmpm/FbQCUlqFP1IgMsLqFiJ5Z6RA02wHmxj1axZdRiDdDdPrZOC
WiBtRVN8/eCImLQBH77ZbFBNwTzVA2buONUneELCQqWUPrYyc9JndQPxq8GX
D4RoOPVexek9YnDYXNOoFftneSy5nrCRgruqPI0wHtBg8QFlLyhNnks0OUgL
0miewlwMBWdSMjfSY+lEXi+EQUENc4M74kC6eETKgjlbaiJuIGFe60ON0KNm
Q3Ws3JYq2h3i6xx3EsgQp9ekq/EroapJQUKjsd955rRBe91RLIPoxDLg/AUO
CzPIkhpiuuUVsQ7YTiOP4tpIkUc56N2qh1o1jdRu/BJBcY4D5cr2JqrZbE24
lX5ofEJxLktfloDDhBM2MCYQzlM8C7zjolvH1lemJxyHT+syHdEhTvBBRwOY
IiYBS/OAqFqtXumU2c/YCbuaSk7VSXxM+V4KG0T8kfv93JydzUqvVrFVKwQ/
lldGTLjtLZaBlZuT0GFqzfnVvGQvXUC7p/N73gAOcr8/gSEq7R7sGbC/6qoS
n/XZt052BN1eggM390ASr0FE1xOTqxQJoxl+IAJM/GpcMx5trhbR0WKNoeQ+
CxtB6H/crS9jdBdj1fqmNmangNMQT34mGPWTMbCjkW8CcQC0vXKX3LA5AQ3w
Ft5pcg8z4nmdVCwofYiUpv3xm12O4Lp7pZCI4auKt/Lqo03b798G9c4+iCFO
ieWWfLyCKDzi3GJRMEzUltWC0A6qGXI0OandSVoCaLlY1Olqm7Z+59PA3AU1
O62E4espDkIKItrVyIkXGGJY/t+Sbgox5kjz6svi5mk4UKbwx9Qm+V2TwbMX
KjkAxn2nqtlbMac7jvrprjnCeJfczxMTFKiaCH1C0D8xKFNtGhbGLPif6Od9
zcUSswtAckcM4ec9TdpxyluY0FoUDgQCEkCCc9sMn6ObCXEBgkBXVqGOuO6k
gluGd/ctSyxc81FBb1Y6prTqvelkytwqP+bpVbGdJPUWwSZscUOOHC+WyTwR
W1ZGPP54ylF0Ao/j76sb4fYTUZ3SfwjLNE2vqITI4jyNpaqUB6uR77pQlBPA
8kOg8LYR/tiW8gJ8XezhNu/i4kWT8xhSdjRBQiPFdvsjNcOCiYW4Egy8yatE
Wtpm5WRUYvrp5gY9qS5k/4kzOXiVbza219nR1G7DBE5GXFqSFz8XEpNUQ6cP
IQfhDUMnxQYFYc6Wb/P+C314I8PI+WEjciXVF9LiXG4GGIKaH3bklDj42jha
No0u3p0IzofgPYdBGXyNMIMeELNAQemULu9TqEDyz7u5z60oDpTxYsw5/aQa
rPnTADSYsNvL9oELpyDKo5vvTQTVxi+ETr4YTvBJz8aR/ndxR2ZR3n57CR33
wZF5JYXHx+3o/RLmU68zbX6YLkreVgLfDmYjdH0d2dybnh7BaTyW/5Im4tJh
6MUbWtp+ajFMsGqXPh38f5wZcK8J2KnoQPwcYrZarC4KKNICIM6abQTiEWbu
2CJhEhSverMHX7SPWI8R6vB400z2MqGjJNgQwB6swxlbZ9Uq24JUHSCB/vqi
LOVimACIiVEB7q/B4rfIe9+2kww5t3t6mSLfKDMtazwTlvsfOgVjJfo244vp
oyeKIuG9pCw7g7DGcqSkveOXK6uvBbdxH2Y5m5r5Q26mgm0aSJaqfGvw3D/x
gnT32y1UppQkpiJJwLvTyCgnRayyoi0hAoQ+D2BTswtQcCJl7A19o7lyuWOA
7FQcL02hp0QO+TFdJ8L0kHCi3M8dJ3jFi5b1TN/kkIM6fdvX4OfW/HHhV/kl
XlmS8hKbnQD993lv9pbssRw9SzkQ1svOzWPKYSKLn8C1dcjKz9sR/jaUtikJ
ZscUp1iXJsfHaxg7oWWyPnhOWlljEHLrlc91/4EZCnkFnoy/OyOMa7BIEsus
iFtIHHkFE66SM0x17HCXnf1O0U6WdyggkO1QxAjf5tFJ+TvYYOk/4s7jBW7t
nV1GObR+V3ym63mkGRkCqtYfMwghZxgRwmK763V25juSTizXtIxDEWNU/zf2
nd/N8SYulpDloIiEpA4W9Z4f05mk3kknV3rC5fLjyOErNuQtJih6Im80Z0df
7o+AV4o2Ymx0IgOEIOp4QD8H/Ej0qtAhZ4lAaYjw8Fc/i6nG3Z0cxp5skjCj
eu/s8Dyf0v5Psxjr9TwzeMZE6Rti9eNQcgpDxONZFDjD35RDYB1AHm7/EWeF
mdv5Zj1FnBkQhNJMM69Vz/UPWmPlqmUgBRcFzFM4sn4Rv8jKCImtWpx6pnL4
6eS+LrtzwyD/8rJSA7/WGmwUrzkz1umEvGfzocUOXq8iO30SJz4I39izM5NQ
X3siUS93QlkXLrA7ZNkTCXm73ImvTYCLhURYwfb921iGRHE2sst3vxNo3H4p
YlV3AwlbMFWKcUlSbBFOBWYBlUYl9beyaTso1N/p+2xvrOdY8e2icHHNwaq0
yUE6kAKngzbiQw2g/lmWPS5ZEpahgZDGmB4Sq3m+4XC5A5p2oInIWfZbVCHS
92vBSAwSP/ac9gIBe+UNpKXzmLjTDYcrnCcWgesaaSyftuh/j3+G1uoWUHFe
FFVfTMByQKcP41yju/daILOqSmMN/lB6oWQWNZYnyryNJpfxY9Ufpl5bHdyM
nHvvTUsR//rDfE7O0wq3xq+cQjUyNa/dMWJNbTrIjAQeI4agmaJ7/CnuIjab
dw7LUr0bDKya3IS21e1Wwn1Ad5gOwWJsztEZId02bHRq8yz0YNZ4emp5k0Xp
BIpLJeJllGJsJ5EDo13yiEYOdX1KIOwPJJ3inmPIDv4MJS6EXTDMNJsbZINz
sFOG8PLSaXTAfjYssY/MKxIYiC/YWsPwnfw3aJ9kOfuZS+XUZPyvdCjax9/8
v/O89pcO0NFQDNg9lPpN2m8HT0xIw841EHx7ceKns81w3G70rdcmiCdvHYNh
rxUHscN3ITK4cAmGDDU967PYGpIDy/lrEf5UQiQ1z3UNYDLD5eCsVXGV2Smc
bh2JNnKI4mU/sc/SMCf5URrIU+wmaveZKQmjRUR11NZMQZcO+ix3DlxAkull
coNk0W14dFTtWeP6IVlcXn7Cihd6WvUxp5RN6Vd5X6TxF8WZqWbj2CWWsr4F
GFK1/WRqi3IZMNNoJehdTSRel97aB3CofsCdvV22IJLe37ssLvlDnQMjYda+
7CMR4qelGXCTX9OVudGNSwX2IoGQmC0oQocg+JlqMGgby524wXzX4FduThBO
akOP79VU7xcsQxWjXl5wovBMOIyjl7sD/8QkqPoJYLSK2tRikBTThZShJ3B1
C/W8Y44/9V/Yn5PGd/A/qGs9ilpbEc6xDwjFDdqwdRwZ+7zZpCBe1zBQ52qT
/KAvpinEd1FYgXIBZVC/JdnTV+1PfOLdr+eovQEzuR1YNfiuyE9wsZIV9xGe
kzdfJt4wSbA2m8y80xGE+dLAUPWhqY8aJ8XkNjuvAYUusozptqDV8V04IyGc
lylLxtojtTMxrQ0IIbUq4Bd9kSKfoShlGKr7CHm4Ye28KIC944nC7hv3qo0Z
A6cxGDMf3d06k47mzazGDa8t375Kpo0gyWiisQtq5pqa0dpD0Fai4ZM6Nvg3
dKy15bDBdykFLX6AUFiYXI48QHZX7dSlNmcxeANKfzRU18xxlrt3V9igk1ae
dGnqhFovV8fCfVJ/XT1bdn2qVBBeui9NP8ib/4a8T3NIdDDNbegwoMP8Tz/v
6AWRfDAHzVjCceUBLw+gUSZoVJTZ6REPMYy65S4KLw8ko/HOQKuzafzw335B
xQkE+bpRziyk2bemRoVduYd+noAa8d/HdBHVb9hwgDKfMXrvwq7l+Ud8Ffik
6tk5zNHt22PUYVsmdptLTJwDGYvDT0jtWzEQvgt5ctr2kRvL4oCMv8PnQkHa
aGd5AFQBJsXddttPrCgkOmVDIobKWfZU2B0i31eJL/uRsQh281MKrjOE+lk2
wYuAXSjvdmP8c/eHKGjT7zswldlreFc+Gf9iiUlT42l+1Ouajqr36RUzkaUI
gy96lQIZs7DN1IL/iwCVSjLTVMcRwbr8mxMk7IVj3DRCay3ypACpAM/dpiCo
+lhjG6/uza4WciQdybd/VTq/SXPi2GtVFv11tab7hW77qg/gghnqLudMN0u1
FRwOajo9meFBj4QuQ0QIkDonGE3TG/q3Qc88vjULsJqqxF297aVoke+oJXFZ
rME3Qji3L3CE2nTtqtEFlxdxNLY+ECQm+Lhd93spcBPlZPh90iaf2miZVXI5
r7GtqKWETlFd6/3qpBgYlfXLOp8GCcHL7XyVNBUyQ3Y14Vv91iGJkaN24e7s
Lw44IY1dtIsiM8eHpfNWftDiu7aPLi0mJjcsn0zfeqe59mhQtlVX5+eqczCI
9OI29Eudvya297N+iNSHs6F2PqW/A9odt3Is6+6MmUbEy220E4Wj+/ksHBSQ
U6n+hhtOW87evInlxB1mcorUgeOv9Em7c+xveWfhaFZNbCCA7+oDf0QmJLly
ibp9p6cdEYqIW638/I2/6sFrwOvXL8iFDewePvjDpTkDslh9/DuuSn65Bc0F
FY39cteIRZ06fm9dsBMz0CZG3mz1dLJi+OXcLXgrJ0pJN2UeJFoIeBdd0NW4
cocDAL4+N4auXN1Wo9tukqZUsXZl5eCbTAY0NWoVUtb32m6PIt/LoVXPzOBa
NIDsY9hzrRm1x7dMGVXv11JLTYdCzK7DTpq7DSA36+R9FGODHuydG19xTlAi
y+Xa3SdH8J/uo8Hnb1DrfXLohH1ZoYbv6uvB897B2yeb56muUeQ28YalNuVX
9dJoQLCOr2R4ZBmYj8eadC2c3Shku5Vt//zz0gRvTv2JLEpqnNJSibaAm9Sx
jvlOYzV4coKp3qfcSI9DmQt7ovyzBUa/aMDlRqpJJyDJQGDPCJGtzToIusbo
XIfjkJHX8qyjxsSnLQLujH8zurzBzjXtHtlRk3FsJHMGaFlxL5lKZddnw3T9
5257NWSfwOgFsjy3SOY1xkD+Vyrpri+3zloH7R4TDlz5YSwvj7QaXQutoZQE
1dooqJDxibQxLsPAD7AvSMj4MpoPJpIwcueFiPr1AbzVixmNx75jLrUo3kPx
hISnePFHugSGOlBxkrzthO0ZGRHR+rrAdxdO71SSoRlMISAP1sOF3THc5iuT
SieMrQF34Njs+9thMGVVHZKbwZEnX6xsgc53cLSQUQUzTiJH2ZQsG0KytFh9
BzMBQ00sO3/QkGoOhTCjRJF51P/t4+eLSiZxNaIzCm1YQdw0htc/EoTCkQje
UxzXVAE9vht136+nxmiUvoBD3bp88aCrMBz2h/IzCgvMGs+EO1bgU8Uiw4J0
qAERue4yAl0NyWa+Aa9RPP2Dds2YPINLBoahv2C9TqmRluVYZx7iV3/uWRSF
EKZoG/SN7DAGk5MJpDqQIY6evfsaTCqrYFV3VY5cgRcuQDmiCw2caB3lY2YK
hZ/eu+yDl8WALuuhyYzJ9BBU+OGFsaABo5E3iLreBAblW79Q/rezrPZL98bb
dMieXOg5Vm+dkC/lOhEehAQRLGJcymf1/evAY1B14zpzK1JqEQIYdu2zxffD
HdBOIv4mYxsVyXgavCSnM8/MbrvaHzPHaa/ny/RKoLlWMqHqA4KWGF+PA52Y
+l8wrfcCeb+tmWpg7OeQ1QA6ftFZIUxCl1bEjxCWb3rq0oP+R0XZ5WNVMjuJ
nKoD9cazQTRRXGnTpF4yDGa64cHLk7lJd0He+Zn/jzBytvyk3bUPZaPLIwcy
QdNoJRoj8Wz2HhWWS7FIi7bBAck8GggZUGggxyNp/APk+zfUbHYwC1YR26YZ
wNyLEM9+3tHHIWF3JKDVojMYrGQtVRuiJCUsczg1NNfP/fIi2uDxG8BixA2L
YLA1+ilLiR5ZPPW085UumYbaCQ77BUEetl+LtAKSsooPm7dl4Afqvnx0dYFy
n4wWL7zQZjmIcYURHOd0RtHc3q2RC0QbGvSBZzkMv09usTrIW8vspVzLo7D+
QlZBuIoh6ObtNomSwIYEjONouV5EJeVSO75A6dDnnvgm6mDbPJlXDe9Q1Wj6
xtuxMIBw7gLaTP5noXiRATEYXvWc4i0FOBBDWKOG1DJW5shmL6OTpVUcipHt
rOXySLwrAz8TddQlzCqmwCI1P+XDeB1R+A+aCu5K4rFkuT9nbU0z/E0u6LxG
BgJiO+ohrZw0pBVzkbCISviRpNNshY8jA5i9us39IlHYjRhpKPjZbZRHKCca
WM+3bOSdlCI5grLtisjj5ShdH0Wz4o+p1W+M0R+t64Ogv2SPs4ZtpUxE+eth
xRBiwQi77+pvsOyeVg1DZX20J+mX2pSKvfcnEnx57WOi8UNev5H4r3rlSGLE
2w9haTKJVROqSAVziwXXZNp+VopI65JZHbIIee3UudCspWJ110xWhp3iefpJ
US0B4+0aDRPA1kI+TIHo4R/sz5rmObES4zx9I3IgpqkxnjtePGEj9QUDHQoe
ItGI0esHWZu8OhUY6ACwgOLiIlzrPpXB92F6ALWYDTNzrgJIqCOhdLbLA5M1
XTP0RwAByaxs3FsLW6nniBwGq9Jx9AhJIZMt7XH6+6yPDuPIka1KEOpkkoNR
krbV6TwIvvYRchzXdAxLw0LJNiv/q6ZcdosbXaRiNFNzs2SHdVZRydDBXWH+
qP/qKlfpsRRlTJB6iRhN9m9kdvL0zydETS3fX/sGJ+p9KSbr4znT/OVoT/02
aE5NWSwzupF5DghjKKxTdfCnzVAJGeFiG17MAbnJslTWw+yx9d9GWT8iczA3
Pch1EfLItaq7zrwzdJXgQucO5fYJ4CPPzAK90WFzQ7PZjNxonE9BXIkaCRLn
j/U3Z6zlEy5zKqODmatCNkz8EFnhv6A/m88eNzPfLrhN9ha3VrGyoPpD4Oiy
bjWBuNL0XbXfNNUKCwtIiQ5oViKBeqwyuuCxNIi/Oljg90LOSHkQXbZpicrg
2ZmLuoTCwsp8PPuAGxN9L3dG3n33m5a/HfnXrj7S/IcpptxcRrGK2G5me8nh
neVfRtuvepSwt3iuNgiHF6WEV0eHeiujkLGq6QSqIbHJ4LJNai8BNcYir3uM
kgY7tgbtDiYYxczNEL8VV8O59yYAXwLgnmii0HF9UP3+yZM6/UaGCCJJNs++
+6y1SIdpfhurjidb2Fgzde1A+9rv6Dwg6NjccA/pmDUPzPZ4ptK64p5BBMNN
Do1TrBy9rHV6Nek7i4/F7bTNI5bymas8YnGJYotVylmIp+S005ZuRTVRGXiQ
TA85Udfcbvkh0XXTRnZc1IRwteMJSH5/c8w7B5rj9MJUzSeWJs+A96SsZ8JA
OoZ+wfgu4WvlAhXu/4mZG/QiFLHMSY5l5vZyPBL/4/PjunzDG79z0L9snUT+
WLvLwX1j+fwwXws9o4uK4o0V/E2rqo6PqIAwVwMqPs/rUKX3IitZy8Ka/UCc
6hdEgp1p/JjShDWyIAwePP0zbReVVKQtRJIKlyrhtzWvEuZ7ir7hMW0TzEkU
rzXheqpeQv3FwVF0ROzdWYg6rrM0CTokpjubHXcrHYswy9jrc5pWd1VK9xrl
64UIj+O2F6k8JPxc50xs9I4FrpTAH3sIAeJgXVg3dUgm909zvE4SNTYe6bZq
Og61M4ycTtRwjOR8YLk8y3+ONWT0uzE8if0qk+DhlBdcZ66kEYQYIBvYidvd
EddZStfeOxzhs0gZXIRkmeJ1Vr0k7X8BVAJiO7ovEbjAQ4Sg1R/n2ivH+K33
Wdl4tzFvwHnqu2FhzA+CLIp+htE1jUvs5oZkNo4+zhafciLlmUDunpenv56C
Jiz8X13nG9EODIKhXHRnpR/YjFRMN+PPk/TDh6MSrk7mAVb+N5L6vWmVpp9U
eQXJv8AWQy+T/3qgvpMpscfdCSt05e1pEq3Q4a8CrtsU+ZOEXivefEGxyIEs
LEV4OXst3RpAAiV9ZDn9xw3WRYXJqYnMt3VzNPp8KJlXZzQCrE8SmnbBzYkn
EdN9vDaRCb48c599hIHygh0BDP0Iq/ez7VVc9XWKTsXblHBCvXebMWth0LQ6
BeYxYkUlFgrMQ3y4gvms8UFuAetmQFwltjIw5mVjy9IkuZvHUOPeYCMr1I02
oU7l4gHZOFce0qkk9bToTKkNsSts8dzBBdo0HtlVkf0BfjlOb57/vzzZaNok
v41zRQd/hLmE2ViPcQ39NGZvbVSIVT8sQ84w5U0dHYmkRZH2yvoXK0Yy7P8C
TKRxGtyPUbh4Um26762AoBiGO5Wl88nIAVeca27+jxmKi1b/vXqKVgIi3xeX
KXFuDIhHuYAZSLFDqnaIUl4C4do3X5yVn+9hjxfgiFgmivXplB2vgxUbdYuk
ozOXrd1zSbufMPIndYJEWyPj+0L3OXvHtW/gTrEujp+0z2b29xImO8TRoUD8
ihZBBRweMIaSl/YQDNaFyKyiCrgY7FcfPitCMzWZfptNIph7z7WPziX7tIRe
SeRS1yTZlVo2raFHVNY4K9QpePwgSU4FwlYSdk8IQRNbCkvfRB9T2GfkPrke
G38hD1+jywqpbZas+wuwwG4U77jSJCbXYrQeYfi1xtM8NOzw/YyOCTePD14x
i2wlqHH37hFKUc0rAWU75kKIdV/fYf7rxvlV9HOyoLIAF45x/Fbn0zXjBWNj
AyiqleIvtZood42NJtNV1oj/lKE66vi4sPL+8mjkYgHJk4cuA9N43JULgYLa
Z10eFurDSuGUHXqvXYvneLNVa/73hOrmeL7RTDpU0h0NtAMRY/MLQVu7sC9Z
MtKccN8wQ1bxT+S/5V7KOhqcV0u+AuwzRyxOtjLJukOGO0weO/3bS5oVBIos
V+EqTBVtDPTd72mDBhkyx/n3QHKq+h/T02tf+8Juv04Ckii9nU2neb8Tqnr8
MQ42aT+n06fIGw5hab24KZALPKDfAI8w1zR3/dUF98kuIbwJy/SSEGy3fdkB
M2fRqxWZ4NG/PfRk2PgXXOBxVWETHBlxdDODSMdu42J1CxCEUCgVesRzTcqR
5/Rx/ROpZMivXpo9Nmaf3M3TQRER502qhuEZcsKA7Kb6QG0IwtGSaCwCIUAB
/yuVV1JHuD3HNSiDBwlRMrIb6kLpCAmXcmC5PEbyVaO2BVJtRuqRnumCOpwn
EdErU0/MaQNa8sa3lKjP4/y0ZwwbiWu4YwvP0VOo/+KFp9LXpwCPi3oPdyjm
756+/A/HiEtHjG5vhZ92JC5n7mIm15TN8lK8H6fX5So/35S6XwpoI/pLpX3G
OrLTkhgmLwhoDQa2JolBxjgOddEYjz+MraBmrINPMYUZkxTMgTePDj/isWtX
dXbKGEIHHkJKCJaoL4hX4IQtTpzQbVnHI8q0oUtPpP4E1QVyGYjI7589WhZO
OJc+6D6qKK+9Euy2oUjYYgcvUZak3ngr88KAqLcyB946eAvGuRlzcmQjQDyH
xzdT93h9qORFL/B1q8noWl2bgZYzg0nSffPN+TBQYFXvCzGalGFP1ya/yav8
y0VFHtgEQw2AJtUdToWy/5JZLBJDHXLeUb7ZhnVIw7oiJ4Xx6DKgwjpgi4fR
r9slnjaDt792efoXoycA4Vw4n7sCvCmkxtHaMzOBH0v2gGrDbepf2CBM7Kw2
CuEVaZUIFlO7mecG+T8TdWNfswt1hso71H2Tk5HNMgqNTxST6ue6gnU622D+
BbFZ5vgJqmQfRe0CtorUBGPcqlUl+D7h3Rkm6HHh5UrHZ1YmK0UoMI637u2n
yTs6sOmdu5QXHa7CLJC7ijeXOEMaP79QFRJCkNR4W6nVP3XG3X4KVF6Swbr4
pE5Sg73g8zr6ZjcYACwVa/augdzyoruqjkriPo1mqxUdDJUANDUPzg5aXaPp
HcdJ0YBNHCoEC03kajZeUv3k2KxpQHbg5SBaBHxpE9OSMCI+V2K2sbXJ6Msv
Ujq8MgiEnjltJ7U9N8PglDytDLrmKGBgc/bHCiUh4Wbp6K3nBudo7Fau5svA
+NhEViAT7nemlsi9pdJtqcRqcr2rGNnyYIQ9FaETNiCoqEcYLOZV17AUv30g
ue3P2mLzrG+VxnWFK90zusFzPuB+F6/kK2sUuLkbUujBbyqV+BqSu6sA8F5+
W9x+IU6rASRqlB4R7U5Q6XS+oEFwkRJRrthmuPgWacJPzb1Zjbpm55leVQj1
+6wBaC0Jh5Kz/Y5JxOFoC1A6EW+RcoIQXoeRCAP9easnoi9A5tJeUzEMGO/y
xD5P4h603fwuAJ4JxRQyfCuHVYSwvkHvKybQdO0DjHmxlrkdfUWfx8vXUrbV
mjnFqP0TaKbrzT3LVVzDSwfOw+uWJtLIYKCBZWO+3NxMOVlvxXOO/2gwPvTa
Uh82UZJjlUH6KpvdkrxqqX/HGzuQi1qLlYJHInfCV2mAEHryXbAufQAthKQd
aCeHNbHmA8usGdPKejvhbPg2pYvW+qzuCQBDDhjX2/aBDtD6vzwQdclo2Xy6
hXci3nKSNap272Zv2W49jz3kUaFLcL4/mv6Dd2m6WB8GssmBIWgBci3lHl5l
AyhzV2buRGwSI1wmnFlcFGB98TplYvTj4AsTyeM1uUBKD2/5jczNa4Yt20Rc
EOsRISdsg0xk+wyKsJHq4Tvxm4J57WqHlNkUISVPxius81ui5Sq1VY8BnpMs
VRMsEZdfvGgTCzbpP/uTR56+op93KCkz5OyrJxqYc3IBd/s/LopzMLFpXl8y
Q5sAnvkyGOsg9mq7WkdARbOqOJ1WH6FB9ZX20dIaPPi7n/rSxWJHDTr1UH+A
8rjm44733UiQh4FQti5KsxiR3xN6wbCmEeAaUtK8zPGQVb0H6FeS7algWLF4
fQQF36w71jGenLWjQAfeH19rXZUVZIUi2xMdQl025ySovuXu2vUVv5qUxwNg
eYi2MAjqKni3JfsbxEI+5ltdkjsxuRyJZHs+fsYOAHSI/HZfMN5LSgwU1sMC
q/3JFOST+gXlMFAVP5hul+doIViS+ha538wmXhIJk0lNDuiMB+OGv2ZT0pEa
jb3J9FxtKSx6Lh4MFv6DBLy0aA2npYr0XBLCK1yFyMBNxiOxKt2T0dpzXe3N
0quZ+ZLJTmKy/2aBV+m1hAmKMsEn4wWVLS3XG1k21+KPdjJrJoKT+2mD43XQ
VCfKQIRHnenJckMsd4ViO7KEwZUukIjQSITA3UFkQFVjct8Wlc7ZI58Eknya
YUWyCt5v+oo8SlNCKVP84zUczr87AGQ1wUbZyavG6JJ+JAM0JRr9Vt75DFoY
WMZTFgZ95/f6/WMS/4/mCZRZgMrgd8kp6YEEb92fjq4rVAlI8zh4jsCKCywL
wRTNNbbK1NWxce/KmuX5CboKqWzu2qrk3RRYgE2CXBYqZ6iItNHqQ8GIaqi0
m8Nip8gpN6SQn5ztUter1+Xh27bADZq56p/AXQ5HsuXcnXu2jhOeIm7LUhTS
hQKDtxpq/TryhFb2ujsn682glYCnIrbSBlqmSGDABwy3wCpZVqou0HyEgPiF
+lKIQyQ2YDRFR/vEIkKlYGbpjVpV58pV+7b24nnngbfygtW8wFxGMrtAKFBQ
CBdtpqKTwUxNp0h1Xloe2UYqPfosY2npiVwUw4T2WzQQh467BjODVH/i0Xh1
L5KsT4SjXOcGXNvstB4v7mFBpp1vjreZjAu75tkrK1HX6cofnW1Qcdhl+OoF
ljrWEImpRBOCtpPwkoxwaG2VEUq3FXGhDGzfzYbkdZ8blDbc8yKASF9dO+EW
g2j0AyjSTHCoHp0Neuq6LmL5d8uPEmzmc/qoLUkdJwuOCfj1Zqa2725+2AXq
lRSEXEaaBjdOYV6pE1AVAvnCe5r8IbUZi7ywmgDLO98MAg6XNVrvZsVa9i58
8um31xUCMf/xOGFL+otSG73wvxph18TrUJ2X0edlNTpzrIdI41cjb5OjpGuk
vUBg4rUHr3jsptBdLUDKwJTkTtH18I8QrcFs+4SfPtnyCnC3TQBYJvPlw5Xt
TA4Ob9+gWsGWc/gnYR0TnlLOR2HkheX0sr87TZZRe3UFzZMvppdfTielZefX
MpjN5mZ6090hooUqRbMeoETJ7A8XxzPuwEtPKA2Ia63MdbJ4zd/O/jnsS7hK
zjOFasZrK3l2y5vO+ZWKmSnx/G2FizGXCbR2VLWysG2FZdb4BmwetqhOfrx7
ESVNa6qnKDhBrfOSBlSMfzAzvE46XK30KunvMe38cRJqxtn3tBouYvWlGDZK
V+vwvyJTm5rTmGaUD6E7FyrzZRIASCnqWcycwhFbs7LyFugn1ZAC16HaxLgG
zC1mLTB6b5Qkkno4RQLiHET4gnc1Izq9ZRc4okWC1FVwjkHOLvp7puJUmg7c
uP8cFpLl/8jAGbPo+VN+hMd4vCcVXLAk5wWgBNLHO4wTH/pe0JIxcxjeWMUw
bSuAfMbvqxP1i17H1vOIbPvRp814Tx4MO1f9ARHdzVhzGHynpyS0o3G7pH6E
rnwbH8ik+PCto5nU07zNaTa1LKBLsKY+EVr9Ae0ugPHcSlyAkOMID4pPiEND
XhDmehEPYdcdXdBv6EGZhkIY5fA8qwLyCHdW3rsOfoL4kcOAkZimow0/NTVA
q758a1/N2P0BL4DlaQ20VKeKD3ehb9zmOS4AgPEhUrKGCbIiv4pfmBo0FZV7
ObfSeTldxTRtkyEEnvFVUKgSBbgILIhEBDP2xFRhsYvfIUKDTF811weGPDvv
tBqubd4Zkl5ruzqen8mVaEvFGHQ/lvxkb1indETSbsv8wNX1+tb1OEr39jCV
x7LvtB/U8fjT/2gLUj1yzyfZDtqL2PelmrbvhSvtTDeL7avmecT4xwQ+Xd5s
BgrkvAFxH5HeF/Cmd2CsrHVZe6DBR5GebNR6TBKxvpooxZb1eo4KB9bxd6l5
iKvi5wmQV69bdtGqNnM9wbaVI/vyVerUV3JsF69AGHdVa1h/2tF4v8X8Yxrj
romdPMr5wJIq4fQWAksOEgTgFvYBBulyqXbascgNGA/YccphypjExPff6B6M
TFXn3Rj/M+JGKaTs5sXKiM5EaezNJA1UPCKyTziFZOrQaBh30DBC0O/WnJ+u
HuqGSDkR8HaBnWC9K5rLyCGvl0LCLj/U83wFeL7NQRIT7gj+8/M0QNr7FFHX
dWGpybzIhDKPXCr2LO4+Ft9GAsiRykXjMZbv5MHifQZ88mxvP0AsUkrfpr+k
eWvElkSMPNpNVFBvJcQOjT34NrfxWRFEgVp5BtFvg9RYh6I8xF3ic7LfVd3s
LaC0/0HO9O/5vkpySxnvtNmacRP8OnVGChMi4B/Tt+zgnpbOYVa2Q9wwxAgs
O9rAkHKnCHuXqJsi6OTiMFYAgF5O+iQYV99ATxUDqw9pM0+BvhZqLKLj1r5n
wh17sSEjKa5sWQzE+Ehi8vgsJG4VzIksGrTXCY/E5ZoiFsR/OrjA/4Lt4IOA
4iWYXaCC/h2T7aKHtURS5X4pDBEYmd9TzQ+dZnbvvr/WpaBW8wIjQKzPc7L5
91oK5HNm1xgP7SbHHNr1hBLd8ihswXgi09zgmMtwwS5x5E0c3pBrABBWkpPT
12in7ZvAle6wnx/qytra8QPRCqtUBDG1eZxSvySNDzKKzMui4aBitiGfS4RE
oL2g52A+JjzoYtkYTtcrIBVleYFgkNuBd0K+p5c93nNZOVrrcJ1Kwl4qCJxD
3foxjY42MbHhsOcYUIbKRjZHSYkxpfx7kWvlc0JMRL/Xhi2rDg7Rbxui+AfE
8GaA6xtQty6DiSnosrmrygne/2Y+R5RvPdcaQBX/xAQXoEm0wPlxIo5loTCD
RYezj/bVJ6+2filce7sPuU4Xlxsezy4OPj8VI8UxuWLZfk+c4CAMyGrkZYp/
QMo0XrOackFO9foKq4XVD0LWT4gBX6wOvwFmwDzKNAGt2OsBdDDTVJG3SF5o
WI9qC4WG+oNYcD58laNLjLBsm7Wm5fsdj8pToe3Owx+YbxGpV5kQZO2zfitP
sM4+RT9Ps/jXz69hiCX83wYyz2qocaspUgZeGfzIFc9l3Rr6UKj8D7Q932mC
tz582u7uONiqTZV5koz/y+EClaaUGnfAjsxvrE3BDw/mXlVuJ4MDiort1c8r
5TrQ1/BbNCM7yIFqNjQlUVCYKa0GLTuXfzsP+SSDVxZJJ6Q+iWOf97V6qPIh
q19IonIw4zNVkdeqQqUWlI0RNxWe839/jGxxZKyk0ccqfqotPCFskXbQ9ofR
XgXY/03mlTrSJtmdr9usvA37/N5Fa4PonSwmrlBOuKhSZOB12q5S3UGIZKZG
vevgr/AAqx0WQmMLYcjxPp9eYcHk1VgqlAE/5D8MG4Mgi5+0w383iKdp5bCc
QO2eLQTNqg7120U8P6KEz62J5CCjdNWUVrVqT5ZvpBQg2FbDzJgnLdgXbmIg
XgVfDMX3ISJzsG2de9oWLGioFQ5NOc5JTSljGZWKCrUd+H4nqfwiFAIZyONp
a2R7Luvr+Ck7uN8znwRigW4zOO5JExZZ6pYIE8eUIwriWV5lJwq0ltFtZYU+
XRVV/Y8Bb1HjcooHXg7C9cJdN3TFUfCcsETZTSHWWyO5fecni1wCz71PTg7y
ah/Px9G+L4kZ1UWYvkFS3nLHCL0OzlOXtO1e1CESkOa/M6WCpf/06PPbQo4j
huMv18I3y0wSxRGbHIXGrRhyZ3sQqgNk5F4YIhNQzXBuWL+qnNINBBo5pJUb
LJrakrENOVayAVaR1wAJLEduozI5YFKe8izVK3F0dcUyh/+zzJ/WBofYBDNr
kY1LBmPUz+1ABYjrE64/tJ2UhtNFR/QNBGUCp/sI1oJ+Ep/dFlnWIwR+nNv4
pQ9Lax3TYJUR13knf7f8k4JFmHqxlgrqIbjkWoaBr4J6bdNQd2K2ESw3n9YY
nI0qefvsuLvE1dmv4mv+IP6ThrLfI3jTAuBBc+xsduniwOtMVQZf4pBKNpQX
AXYXBsqS2XX6jfcelhyjy2BN5jOE5DnPJXTVP2QsuvStlxRfKad9+ijvkb9J
PnY+ve+9jWru9Xi30Uneeo4a3BlbnJ5U9QVQ3b8ppM+Xju3J6UkZP2Kgx9Wu
sG3+OLjn0DAL522AN2gJ1pezdvkxgh2qdFX2jx5kufFW0CS51KE2viAY7+Wn
SA1//28s3It6lQwC8G3VfP09Q3keiFguc5Qu8pSzOpjmEDW+woB8jxKse0wo
uvS/+52TUSusM2SfTSewSdy9JaanAtg7aUZQyHk2kavdm6/uW2P4YsHiSD7N
2fYUcJS2C7w/pJV1S8xEpcsWXKV+adlutmcXY1JTFnRZTv2vNI74WHazYmvJ
itGg/FgB8WMJ4H1KqcTKvBDdnFCioTzfD0lXdOGoh7/ooUawhdjyU1s89+9w
00u8U3gqKq0YGorELl2grsECfPE7R7RIMvdyje5LUrJNHSbu7iUG1vj7rHZh
CM4gCCUBp5riYexxx2/QiVJ1kkrWzeTBg2xf9w+kEqyEG6Ywcu06rWAaWwlE
F1uXfBkQkgOgVyDf5t5QIU1w8bwG0o1OG0K9662Sr8r0MWdvgjBOrTAuEO4S
IkmJpKKw+pMaDg+1s/4vVLCDDZ1PPrnL7dkFCUdJ4gdB1GYqTLmHjg3nIm8q
QdysKaJB3TeFJu+yO3E7gJ2T/R5vE4laTXJKA63mmiBgeEfEfnHtrCURAbWH
obx2hoxiguwEQNJRacz+vM2gSys5pdRLPZwYLHQvt6tB3H9OuYyql44O1vB7
gGuefjrp1wDfIz5EdVj9qqAg3VTPReUedDUVQsXS/J8UPnNbORIYvFd5yEQ8
lsdhd5bHfSkhYeyy1mOMYOs/sOULkL5gVbW71oW8yomznrasN/7ghdM0Clka
BrRqj2JF+07HXGyvGJz2hulgHf+XKjTG5592MbcfmE6bgv10pkyyjI66+Oc5
zzdGSOjgDP11+ntdGJNVQ8JoB8r7fKiitmJwLXfI70wJxbKhlu+mWXS6Na5/
ATM9lhiNcJ8XAIEoiGH7iFKvTy/CHe/O5QyPHoGbIrIjoBq7ivuyghceTrA4
ZvsTX9qokRtKh+r7BLp9fpm+L1qhra75oX/IYKQiSOhgYpIfsUPW4NUMimdU
LbpOvzq1I0O1NrVEKOuGz3YDCkDstWjR7vXVEo0H8W+H6vdAEpZYSJLSowT4
NXU/TN26OsF9JBCDi9/uXrDgwfeWf62yh/HuTWX8cFU3DB65gKRzxW5el0rL
bJBm6SQjk/mQigACu/pgQMw0tSL/LNRpB4e2vFX998oEoQuRMhvE1FXOJiat
QDoP5xVmeP9q7ZMUiZQyi3V0hW0xFfp50xxGICObpBVaj3/0uHhPIqIK9CJg
iL0jgRIkphiaePPvvly/IDcG2kH6xiatnZyJojxuIDgl7pgZjW9WVqkWByL9
C+T4rk8DtvoDutpmyRNNT1zJ8LIwscmwG9f8T6DI6jf0MoFE0MAgHIyuBmq5
kFE35x6tm1BCztXJcSmi3aGD/w0vR9y20tKvVugw5v94Gt7W+Tm79p+oMaTQ
3vxe1nzq+Lp2/w2i/92TjQ9KA/8wDiV+vrstKnsPs3qjOVn9n9/k6AzbyCWt
Ya2Yd17IXJoPYPy6iywtOCHinDVduVj84WzAN4CmP6dn+ikIjyv7WAxzn+DK
isb85N4Za/QHCgNUSZ9wQhXNfJ2zglmjsWYo7N9/87quqdCd+4lvJB+bkU7d
dlfrZcWcx+Hq4iHxxu181w2gXLsR+rfh3t3GTV7PN8qP3Hqad3Cqz6KuGN7j
Pgys7EY92aClbDFdNDSKWebqC9sbs3UkHRmgTiosLqVoy9dOr4WcYgKZYD26
mJkin1Ww791AheF5IWnwRKid0dYfrflNm/wKnSVo+61IGSn4MY5IxBRb25Ah
ZLZMTUSYSkKLcyxIYAxYTk7YOaON/5LX8Wf7bjWZDWKdRXWtsg1iZ1d2BrEX
oGzHcPJxQGdA2SRYHfEUQoytsOnEWqp/dcR95nVCF+i/ripjEUcBou7jU6+V
CEAM4tNztH6SnHFVYdYsdQvvlJREqtuOt+PAWPOljD6CoRGNlfZpImsA9HHo
gby4V8s5oBOhA1ZfsEpzwdSMrgW2dlqeLt+xkD+cBDqlcn6Cwm5GXGEIj5bS
T3oA7SxCRLXhNIWg0sIoxhQ6zTFJNQ/kFYj5X4tIjgAjX+YSnV4BGDQ4uYrm
XWTP9f11n1i8nq+8PCql+6oa1up1x8n5maXrX6ig6+ikwaQCHLUTvKUAN+gS
iJUnPuMEpduJD4F48cGg4BAqxNVRX+XxfW4PAqT667ChbD4FqEt/qwXkYb3A
TOJbViwpYgtopDvXiJ41guh1zVHXbwqocG+D8VB7gJSpTxULM2gpUbrhpmk1
PkAGh8xC4Bf7xQXH0DEYOzpT3DpOjXlbNnmbqDjR3WVcmXwdlTkis3H1pKeH
sPuiAbruR5peFMHzqjFpYlIUrnG003ClelcPNwJSPAjKikkSXQi52plB7wTu
u9FogBDiLSaTbKeM8amJE6Onkr+8Ff6DjRIM7ehVYHx1sVnf0+NkboBkKx/t
PxV1IUWBQhCbgqwfBltdQ/5ouyNOt7L+dwRSADl24YPgfmFjGZjaxKjptTfA
A7Oln2cBjYa7ceBtv3UAQZMSX35xoO7+Yn4TF+hik6PyN0iEWoHZXdXP3Nfo
9jTW/QpTGCalFZ90CMbwoPrsR2YqIBKg+AZ7li5VtpqvLqMyGmS8SCjZJjyL
DNOFAKHY0ay7mLJhAqWR8lsGTsbuTIFDUkQuqoGmaflZUeyKfWSfS99am5Wm
2gZ2z1hO7gQ0lsjDBPGg31ia7QayjqhdFBEoIxkgLfGJZ2Db0xYoQit2QoIG
LbFdTLKn3xIJ9Evek8doyeGtZhw+o4jQMypnED1b8HzUtzNEQWZf27um7sMe
j/umrcoQgST8wXYtr9y1Z9iS2GhKcb4sUeTT/qC//oI8hI34lEQaTc3dO0DF
Gs3mkQBTaPyEnaeE4VBN3vz+KpCDbRn2JkKnHlJDKgzP9VvsJTtAhAsmRChl
2x4+GTzGWy3D2Re+csYJYTnAtVe013h+gmM36ZaSgzI7cbuaqv1S6487o045
e7quZPk0Y0Rh8al4wk/zJa4eAkRvFT88GCDDbZMwI9/6O1lAYL0uQROxFhxA
G79+nddUILh6EiqvTU28P0O+2OfXySaHCEqrg+Du8cBpd+KCnx73wXDo/rLU
SmEn6nQ3Rgj+9gRepQkzw4Ym/lDJh6K4Wpkz5ZP3tvvxzd5EutPNRsrpei8u
RJ5tg/gn17SEYcD4ifaBlXVJgjso9nA/GRZgnIgI9hQDWSSzKRMKkYomZCiJ
NnX1pnKNV3bDq6lX9t4W1ckBxHFn98izhMAOrQLoEAp2CK5a77Y409tFSLXR
q6Db/LGCOoKfAPzc0AwVpC04n6A5Xq8VyyUMrcjiDm2voPMao2OOWPTmn6bS
qxQrQ8KFlUfKTI/s8GP/+3us7n9eed2VlMqWQwyhVTuTgN0hgL1fZyDuWCvG
p35xYOg0qYrqwB5eUPJbrV0Xs3praLslJu49WGeuyG5rDwAZ315y77fINKhV
/Ax04cX4oQ93OzhJRVk2zIXniiVLoKPh5pg/7izfig8homgS1Ecpl0IZW1AG
XoDFyjUxybDBdN/XjTIPLciA+n5htRPCPpZuucM5dqygJe9S77ID7w7v9qWv
3kUE+bFF4j/bGXQrdMm5JswX+bc/RXGAwqASHUhHDeUeEG5SZGHycTvAOaLl
T5UhMxhuHWc8rUQqQ4ahWn5NyaKG8LkpMTeDK0wxdVaL+yKFH75to8vYTZGs
JXkzCAH6L8k9OHZmS3/GIpdJrrxL09+ziywUlw75GCmZZjLVp/e5C248DQLf
BAW7OVTuTN/VlNtOKk/5Lv1z3ioFy4b5jkXArzpOH6t8YZXamrbD1YITSNEU
8i/8/gwCYnWMGJfus830Y6g1TaUo+YeWVqlF/TkAEt/Angq/qv/2FXX8chJD
WkzWa4q/0aQA/1puiGIWW2hdvOY7sLN3qOAkIRiQ1roCd6JaP2m317HgKXFe
VdMFJoikwBEAaBhTENfl2TE0hdru+WyWG8xSAuH/cxaLlDVW5Gjz9Ur72hU5
2mBG1zYZrxr0NPUXf1mlroQnJiyzOYawvfbBvZmnZceQCSgrUBrp+KcMW+XX
LJXbhInnqUDj/us+7GK/VoXKdUr5vpntQwDZsTnUuYlQ3n3y8IrP5WsdR2Pc
vZJQQLw+Eg3hdKifDnRKeOgZuRlBkzOEg4k7jUgj+utjC4R3Qv5RuGkZ8tTv
267/etua+1Jt2CKg+0Z2I0I88rJRFrdfMYUXfA+LM7/WGrJzzviXzqJFjHm+
Gfc8ZUWoaB0E7LwUGoLVYfoPAz/hRhJ3uJtpr26NdZoKKw2t4uFt0tDjZJVo
Z8+Wl5wR+MlPOF+GeUg7NISVLSlGIQQ08RqFbPMDuLxBfRdffnvAgdZePg78
HUnTT+AGwyPTA3o4tE4EYs2S8GLuTTR3uxnOZUHAk4EFd3+0LKANuBebnKNr
iEQ8Zk6qAVruIoqydFARjJ3gjdxGAcj0CC5PYuXn5e8XM2wuOjkpzc+Nl7it
zQY9+ZQn4mdV6TBUTeUguFjYQkBqIi0ELza27uBqeEwBiWoP3GyatR2DJ4WA
MSU7TJsxLe6qDCoaLg9KPnE1Lia1xfXAnvoPFD7yAke/oAh+7udbaF9fIX0L
D/6vEKfRf7zSFjp86SR/b2WAmDABmpQ5vhFazP6Fnns0B3NPm3JLlT/R6APY
KbnFSEtzGVuWItDcrAL78fP9Co1xtcqz3vBqlAQScOsav/CfrLXYdbpU94M4
bnSUzUcq1ABvWwQiQGDNf/h7GOtL6fcvMyYrp4uKyMIB6diPkwGffwnbt0xA
jr8Vp+9k+oktxB3ZkNV+N+NerSPw/3p/BYrNOBmEobdQ6JGiuy7PqjfqjiFt
9mlrM+X+TVFUV9Tq+p7wiquCa++svZ+d1CnrZnxltp5vKWYEgwd8Jqm9vifw
LEi3h04MxqY3Cap6EO3fHZ4IH4hWS0rjfnZEPlSajgQuGwfY2rTYJxD65wcI
4fRtlm4x6rl8sc1BFsiCxGMSybeTQ9RVquD8fOiR8kijzBdTsvVU7jmnzD41
xcOY8l5bM0Kov95JiouTj51tWb8nBwvh9m7slebatxkr+mVERF+itT26YiR/
3Ih/iJ9pfw47S5ihcE8d4mDiXz+pdXJBGs84o2WPKNg6D+uz1W9a9jseU6BZ
Py4qPQe5EwUUhQ325x4ihyJghix9kgCayX8P95NSuO00BrYxm2tW7iEArjdk
03A/QGWOzks0FA1keOwqVsKj2BfXCxiS7POnB6nfIoV0pIk0hoPQHrKnrSo5
oXdxsWhiiar4v0O+MpZ0z5Szs7sWR03IfwfBRFJzxPScqkszsxnfgt6dlZtB
I3uolADLxg556Y2gNFRUX/ctQZGPYc1mFYC4eVyVVe3f/T8PEQsRhuq7Myjy
dZuEDpCVlg6paKix9EnZL5WAbuif3HZ4YUkVDutvzANKHUVd/1rPp1cMnNch
alqwIn/v39cNJqsq4XB1QFIokdrgqUS3nb9Jn95EdFAmGfdXTZQURFLgWsKV
thui+D8ANG5gmiNQqoTggXrk5WlfiJISmNp8X2NzDzOvZy+MO+JuwYaJvrUQ
IR/yLCdL238ns302iwW5+qBGxMrsp9CTns/G2hHIU1NiRHsmhMuBLvM+pefy
r48K43wCn4HWKyqy/vNgDP1qL2ZRQH3IY+8nlnYRChJQkFQmo+US8EGTLp5i
J0caqSEdMMqpApfY5XBJyrKb/ug0EVsJa0B7ZBXxpMqgfNQgw2L3FBLGf8XS
kYQXSFWQDzS0EpPOBXDWQCo5XXq75k+wCn1dC1c8uNlFbUn2lPRxn+v5O9HG
FSqwH3mzcWdXK6xBkpAV1TajbWB9hHti27+wy+SL/fIL7ocgrw3NaCkKiYY1
CE7QXs2QNFujthgu0gmhOJRg05jATpJrv0Z56LO6cL7R0vSwwqmLt+OU1VJs
z1XLUGCM8oBeTuyRYhJjfJ5Ck4RZ3m748R0s9X/MMLsHtEJCGnuKIg7C5Hag
xh5Wpc+gyf/qN78B0Ik32YcYyHXB0T85DEZmY/7243dHppPj119hXHFsgp08
pNpQLcCh+kzNYE+737pgQ1EOGvFG+YFk4m1J7G1q0boWuwXcSb6w+2uMqKIp
Us+Ma85d9ff1z2N8UOPd2LBQn4od+p5w6n1V8WQgLSSaq3meOYgX3SuopgKF
NO4hvx/sVfO9QfaOlQac3uv3c3iGxGrOo/dcK5lZ8Hc1VDzyqIvdO3ZJgWBa
sVmJPKsM8+bD4meqDK8LbY/OkTvoNGC+ck1eLyouEmwNMSG1lYT2t7SrIXGE
4Tr0jMI+lQAHR3mfiVU83kj4K584gQf9s0ao1yVRM2ScoVGzeyKciOSrkKR1
DnVwTwiBguZg6sDJiZldWZU+48NlgnXqxfG/fZF9FXcgOxUWNyXQkuHJ4uyy
J4KgQk9WnC+aviSDH77bFTEmIiSPBa04FWLlpgKUqs2z3wv9Vub/JMN5RDxw
AGX90m/6n83Xg9zlhpErQVOeLkrT1oaGzRI70WMnp6A0uCoqKQ+1Jv/cSGl9
qjqMyNZ2/AJYZJpmsfT2N5mspNNzGBo0tn1MHZKNXOUtsT6RGJ7pHN+F0cZv
t72s6ZrEGYYq5owfSn/82Fu993Qzrf7prsuvv0446wtcXRFfMezU1rz4qIK2
OQvGNKS6um8ocx0iIi7GTGX8yPkERyVGLP1+IeCWQCBygRcMbpVhLcPZxJUk
Ak7yDsWVdd54umOlYN+KH5nzx3fdLqTo5KOKfCiEok2Y6eggvZixhCoR8GFr
m5yzOd3kEfWr+83LmX18CM6/cV7RAJhonhXuh+XxSRam9FIxKYylFEl72CfA
pPfzwgVM+kFfWN4hDaoY7PkDOEboiBDeNstA68H5IaPb6hmYx9U0c51ebsZX
DRYd1DgiVggUtsSJ5aIe08FMDelwFODH7QB0QC/T1hPoys9RI+63RHADZcwO
OcOVZYoC3qCi5Lxcch0chJG0X/jgkdzpMh9+sAUMraI4MWdmHq+OrjGOtklO
fP9BCBMLLm0NI3FbpZjentLLwmnDIIQj9sGKueCjZTcUOZaeahuhez5Rijmd
9kaGFoeb2xBalhte/07SfsoiwPquUwLDw6KNL8pDDwmJ+0Cdq1w4GgsYVAEP
VobNmS3qMELdBIBapRXnsmcaRvxeYR6pReBa6Unpq2WTxpVcx6yZJ0J80WAO
ALB8NltOf1uKhei3ep4/agVnYtMHwRIGwKP43mY4eNJjxcTaaQGa46W+t1Ye
F0+nMaLz2fL3BwSYG5SauR00cLNkA7gLhv3mlopCn4LnaV3kI6ehxZhyglDP
r/n11lY8397EE9IAa2uL4QNo9aw4zefe11oixXEPLScztoFPMxrMA3rQNCI5
kw7x7lx7CHfFjhCRoTRKBMLQVsmjByRsBpEb3QErn2V9JwJ5adzXZqzk1nGA
Gb0KKRWFXm56WLqBOwreXrPesWpiQntBOWalG0yp6txZuxFz7eSvoZ3wAgNQ
YO0FAufELpgonsbpAN7/Oit16kZ8IMZQyr5HN8p4OZ85NCYO8bDJLwOb/hTo
nRjl6FaPO4j+J4cHWNLmTe2kTElqpcVMFFEJhgJn9EiPrKrysJ/pZQX47bJQ
5bEJqilE9xAiamPfjsqj9Mx6amHF0VqpCTtBEPLYW1BQHbhqJMYFHrj//1cp
B8lIRM7jLMdIG6XXYRN20MklVbzuwtsWreXmImpHXZ7enNFxl9jc4zPD9sFA
P+ehsv43dU0FVWPSMCTMiFkAZceNQEQ6wLcjftVhilHszbF72FpEU+z0sAXZ
DynsoiQhw2CvSiwsSEBC35CJmJf6SMbGuCWhvUS8J6IaFJsrh1XgAMSZ30Xi
fAAt2NUU6eVIiFHfZLo9+gU4jzjpcHTdAypsO9YA8pMw0HF0dT6VuqUzatFQ
CY9gD7M36X7zY7Kg439a6zmyotOMkvSk/aXGxNNHAuGq/U4klJOmpc/GYW2D
TQbafITptWtR6a9Dk0oNHRJOujTXkfLfUneyhFFRG1cHH9BVeVIaXvra4jJq
rn0oZKynjIFHgUbf+g3FdP6kuinr4x6QhesHtq2KJMnehYh6p0RF1knTtR0J
xrjyo7Wg1tzG0QmCwum6NGdZcWlyX1NJRssBgmpMNGyLzccwOswivV7OsSoT
uYEHRIs/3J3qlGi0ZysmH3w3IcQsAuI0si0qEcLmLBF58tEP8UNCLedoJu2q
aL4jVitQJ1Akm0jWio7ejew6HHgHz+bcsSE1TidYG1OL+pCVPh7JCv7w8/d+
E149LXbQqqiuvL7XOFiDNR5VQCXDO5BKIkeUK8VF7sz/CpHMhRaR1XkzGziC
Kl/2yMUmdN6J3uHQeupHwHQMSruapdobebYEBH9XHV4RvqIAihyMrAF1w0fi
Mviby3CaK+devbHbh3J5khna9b1bJJcVnJfvYVlyYQCpBjqM1Ohu4y74COt7
s7mdQESLqzzt0c8Wpf9SK88J0nDxFTZ9/etQbCy1MIrj0pJ/SffTCl7F8ADe
xOQzUTM3rvk0BSRQQbBumRROa0d1MBKiRML7JtkZPAH5+isM1q22Nf7ff/1v
rfWkkxJK83wlv6c0N8fIUi8kFD43mCdty7fW4RXHGm3gxd4Ij/w8Rbns6ff1
Z5F1EULLsGyAvKRYigMUEE2hrEyIlTzjFm9RKBobMZv1Cbsvdh7dcdw4/AcE
L0F3GMAuvI+EgQyQbUOnx0u4CgoTl7woHPrkXAS+sejKhFFbqwUcDiyjvXf6
yLsFYEt6875IfX4mQlx9By0lAwkyzZuuGxAOq2prgLQpJ2D6iqtz1gAYihCC
pSYYqmatT9I9Sn3awByIrJkevtsbN3uK+5acbKOCAr/Q8L4vnFkrTOBBLrqX
b0seQ1WYr0NH4kM2OrPMTXPznZBEsZBW7d0LU3VcALTHsccQCerNFxC6BZp1
7LlrKaQov8VtwWWuyMyXDIs5ajgiw3Gi6AyBdZHjokRnKX6keob88AmTM816
Gji/iTXdEM63ab6yo91gnD6iX/FIpeNDdeApcwMrjXqmxC1fczGf/ehA4uWN
HwSoJBwNwi4PGf4jAL+VekIer5llidDIyPHtMjLWSeoYZZZ/0wYUJ7TBn6Qd
v2//ZEaHv3Wh8GYVN7ncnt4vs4kFAlT4I3mtSG0EEoqfZ81fvkWxbcphdPRo
twtl+xGuHI8EWJDThEjSiyZp2xAWYaQPcQ1Vx7bVqyrLq7YQ5X3uJ9KpgPWA
kRpCHGgG/5TG4tFd2WQm95UuVexJy5kXp7oLgbQ6MHjIe+ryhTeMkU5MXXPF
Ldpev3mEf9r68gf1yWadDagqd7p+Foyv7UTr+HpB/6ogiZr1ARKRGLr10DgY
EpEgout+LxLaFNG2srm9Di5hXvEWtt/GZYE4vqn8iGxJLZHdKwOzviACud2w
H88/52zdIJgCjyxLGwXHK+k7w2g1ca7uSJfz3P6nIjf3I5T4LGNcNvHW9svn
jwGEDrGTQDWpsJoqIHVjLRjKvG5R64TQYUOTJ/ToTSKFbsqesm2IwRc46wZC
QIR3iITraBkw9dix0fQwuu3iflCqlGgKnlxF8kP0do8Y2RIxovEPsMg/x4pP
n4lnubAJS6qYepWBKb1vIj0pC45pl5sns1nXL4dKDISeIAJ5lYxoPSCNoKPa
oRfk/KL3mxnT8ASTUH13G/YUEYr69WorLRvWjs8m9ZUmKDUtlyYzF4b4zeso
xJkc96acGBvJuaJZp8XNIzhSu09X4zAxTTzjl/+b13Fy7GYQQTg0Wmulpk+V
vNzYplcZCPrbYqWi9d3GRbvqpAIHvldYFPJ6EAVPGHKgeI0cK2W5c5WZrP9R
Shn/9Ra9EV9bDdiWcpOQpXbfDkTAutwoCcco0RJCFoaoRzcW+nxgx057hBTP
JyajYmwoxKrmdGVghXtas+1TS3dFevhyAJQEN1TRyCJrRVoTY2yZT+Ft0S9h
0Xa2L5k0dlb1//LKnGyVI9vFjYrDU+m21na6

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpeilKQgCf+Aq+BLK98mFFWiY2UZnlQhTvX5Ev2w1nt9fDGp5h/LLd5q4nwPdoOc0rjuW9hq7y3l1iPRJN7ipuuAJgctzDWLxtgoBuY9eR6z9Zyl4cO5/cErY78D/IrkUtcFd7KeeWLFyDOI0KvX4zij+Q+EwYLueKgDkEToRbxwQoiLFZxnDMjGFKKDqPwwPQFK9jsEUz0lEWBToAj6pzS1LNyquYU5YThR0zMRAiDprZQmA/SB+c9PsRIWma+Y4yRl1eh0m7BbrTQyii0qlYkLDUNvrAvLl4T3aQQeUAcO4xRkw/p690EoJaDoOvf7Ul84PN37hi/lgKWe6QHlZiPxOVmtb2Nf/RQbLf9DjSJH63mZaubQLq1/77fzMCzPiWESQkhgZotp65qHw3MWrYSCZhHycdx5Ap80xhQBXgHstIO/ZG6bSYzGn80I6uhbelEu3Qmf/cMYrlWDyUMqaZ0JUH8xMOOMVaXPM/Hk9aY7CAR4zRqz8tqq84SsNciwMdxK0mmAhlWjsYhGpvr1Z0+SstXu0+bFGh9+tYt0drorOEsnvGaDEeLwWgDUo32gQw5XQJvkhQFUa/bHRxvcr5gCVMsgcI9O3RN6zH+mC/Xu1p1mV2hZxIS2zwZNtSWWbOeYpz0zOjrfNqrKdMEnWvOfslI3wlnwLE6mmWXo6raP5Xj0RhlG0cVxUP5yVNeCviA8xyJoAx02erKXTtlJRLkYlcUanvnCpj9bgv4FP320VjF2dXPjOH5UiNckJiAuKRSkaysdctmByJH7WXFuxq9ej"
`endif