// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
zojJenNdNaIBCF53Bv10iZZ1n9nWlialiIl1hpAwbWd7kajV6+cGoEtZMbYd
0OWnvmHws37Cp4ISvDbNnnow8mj8kXqp7HYRLKSA8zL5mbd0VBFLF0ugzA+A
j9o3jaYH51+POLpr4D260rPBaQMP8Mv4zLmbQ3yHft5Rj0bVSAH4fRBNCryS
xyl/0C7RvFY0b0KmYjB0jFttnd6UmnW3QpaC2Ssza5HRSsmwUkTbz4XE4adn
cFPPeBiGSYhgkIyYpVAJIr24mPvmvxpJpMQ47ss4gH/pV9BrxMTKcZJyh6EO
+dWHXrl95bpm+GaNRGsz+7u2P+1b/gXMFulAz5jLDA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PZKL1haBkeklSqnEjFGBbFB1yh29DSPiRJGELRk6LwkuIbAGEV2ELO4BpWZt
YeOD7Xjvs/aXMqkbbGXzChGeQvc8sozNGxGL+9XZdtCI2PBKgdaNovEbMPm4
GpDlXg+X435xHNdHVZmnpVfr28iPlFlntin1C+GkymUYn78pdW0ELERv+BjK
MP2K4xL0PRDaQzhs39E4zCw2BZWHCCyKkND+QJOWg1d6xDg/018l69+AHoJH
O/s3E4d8uh+brhjmNK86Y3GW3Z5iz9tjeQVgv6aGkTTkOhEAFYmzr49K7Adm
I6jUlvOSqCBnJa98fW9fA8836XjdH3z48xQDEuZViQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZmGKwCSbKI6WeDOU+H6FAWh/TBxXDscrmcfeKgj0hD3ta+6fs8c4HeD883Ip
5Xaaa44+q7QH7d3B5bVMLYbL+3rf2w0iURRZda/djQXPaFB8pfpYzFgCtkZ2
SIeJgE/Xfk6uRrxROWDuJvWbYjPBBCpdMedzTej7HJ7HyYb1EGnaw/rQTpEV
VGy6P+7GK6xb02ilAG9IKlNpzW3cPfdAE+0W4OaadZcjHBM7KQV33SYoSv8r
IKFMEXioeNEBv77f5u42xIlJ2LOxL1YOpQ1EMTzi948HBAWGT90qt4NU94r5
RIe6c89RyfyliuGsY5sBz10I1tRYf8jy3iNyfO5D9A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
m3vEMQBytMUKXIlPNY7GaeWT1GCc+a+x3kORWr1s1YmNkgreFRitJ/bf2/Yy
xiEuAmJQc0mz/rYWmcKSUzlvWSqPo904PwF6IeI8lAfC63r0/2+B0wHAl3Zg
yeabDoBUU+xSCBL2u2EXIU3teZJ72TsCFrWZsrSO5IOpF3XDBKxa3wACGRTM
SD1VcQCKWtS7m+bwv2EuLf+7+jdzK6ZLGZ7i6wzCc+7GoR4kpJp1UMjTqxVv
Rc681HVbuI9BFj4JMF1Pque+G15/0DrTlf7M7XDqcr15wriltASX9Yw8574u
O2vzbqujVjB+yqLMJVnCc/X0Fvh14hWd7s1q3zDWcQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FvOz9VXa21rX9fQ4m32f9QD8WOIAiLidO9siTJfaONaMX155x/oHfumF2s75
EXzxVGnJv7+Bd7ui//qzzNPJohXQg1l3IbLSq7bPO966AlG34r+lVUy9Lmvf
zhw2sEMAE4RGmJkN0fKLA8TClNI6HiK1LYbhjhOuGWEy0YUuUKI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
uq9I/vByHbGqgjmuZmtn60mcq9/CMuTU3+K0nVoHv+LJmq27q6rUbv3sv7i/
aeyMGHWHf7QaZqM5U+ODA2lejij6AqkdB6mGeGo2vSW7q0wHS87f4ipEqA7/
0kt8XWX0g6orj/eYsTPIy1fUCR3lYKIumdgdSePY/dTG7geEBW/hjh7iQAtv
lu7Cy9sQnNmmkwAbxbg7sKsYg9bmgCgiXeUjrGgoBjfA26ov8Kj+W3VlFvts
UDJUpNAkjOFYo2yED+kZs6Xr05gsOUD38XRlCd+pHxz+PNWKh2DVzeNlYMMg
oAK28HcIzJHMZpHn+WxLP8cZZs4vsyJWKEg3OH3ocNOwV+Ifjum9KF5yw6YR
tVY0FP5/G6/Zh5ueMttkAs6lgZMFFLTQYK/qSWI19llAYsz5/mjH/fbToGTH
6iE/wkWkg7Mjso2VUPAFOHr6Lh5q5VurGO7tAjvAN1WWEpE1Rc+U94CyQ/ys
Vu3T6C5qBLDssb1j4AKxFHVLaUyGJmOR


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fD20o+1YeuegN4BxyzwDvXN1vEuLwZ0Ui2epxOO9gH+6Ar0a4xZ1JF8YAJWE
D5wRy0qkJtN8YMkd9mVXmFsLZYugiZRIeLFLnFF8q4YhZwhW/PnKJ8EN+ksQ
OzUwCzH56JAJj0X06qf04y0Qen4jTR03GS11yuLB6ZaB443ePzY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QuMukNFH3x2fjAEN0YCIfPn/NyoFbNDELDnXw1fwtprGNh4oS4f+xN7xr7HQ
sSqzBMWH+uKtpOFy8NZdE022fHMpMuUTRT4X2qztDB88kNm48y14MhaDeveZ
Q/R0UZdvsc6qnYS6phkUIhHZED41ozy/mk9EhyBsiaxY4Cd3L5c=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 58080)
`pragma protect data_block
jGlSj/BKx1noTbXkUY58dOnq7UJpFyTkoTLbZpBgsQK/yTE2Xvu4iS400g66
Fy4g78a1tbtQjUcNVeTRrH51zEB07IJRcLzrv0U01CEYEc0nHROSh9sohfep
rujuIdd8K4ju2y543tm5b+dnEL8FL8RZUaMp+njbOn+/okt59VS8yDQcC3Bx
ysh5ESfi92uX+pt632P7CgD8JC716Q7Nd4EhBBfA4nRWFte7borQdfJsxy4S
2pxxpVY2TJu0LVL9gLtO89Zm8F0v6dD5lvUqDTme5thAZhJsiH9ciFHXt6ji
y3SCuhTRzmdums+2AWrqXKpMCkNQMhuq22zb4yDdgbwlL8ltNuGq/+mraZF4
GSBEhPlBuEyycsXhO0orzX6mUy577ewM3Zg1iXbcr3DfxjVQB/CHoyhoQvt0
ZI2qZTRnB/XExQGDNQkdW2NwMA3Bj0gYB98bbrkp7MauAaS9WyDiTs3TpeHb
aNFjXNCIlPhC4kh2lC+sU+x1mUnNIU8U4T6OAhQGebbe00jTC+BdRAL5iwDE
asAyViTnJ6AyUaDCFyx4cVVo59uf6RiOQOZg3xmiP/QyVn5aw3ctRTJ+Bow+
1nKfskmtQepuwY9OuGAm7rVXGr1EoNi4UsSVnueg12FATXrU2IBorKvs4kt3
5cVS8oQjUPovVZZ0u+dz4ptOOYEn+QMshsxl27PeuaSGocfKh7AQ8CcXdXDM
aVtLoA4j7eGjC2kf+u4g5Yj53OXf+sMubon8621FU6mdtLzjkqLHXOmuMpYd
2Cj9RUoOoKZm5s5gd6b6oGnFiyfjcPJSZX8M3whoZvEnWRHAhQ82sg0/rmlJ
DZwmrT/6dZrWwKpiOwSdkCNrjwTVwdlwwUHwe1bmqfiwlL7HVzCa8Mk3TBYt
AT8IR/ikM4Na7zZsRK5xEhSrjEUBU6iCd+w32GP6o9W9zKxdpXyGWlzdy1Xl
h0d54Wdau/388FbyHe8lFrahwS09l9Z/WFAq2LMNF5vwPoUjmMeB6kE5AaUi
fhcjPmOU4/GsdnrxQqBVkwPntw7qd8/x0oG23O6SslymbVliZz2uFMyzBrdB
7ASmwax86nw+j4yXWarQZOpwu29pUHN9yU6Js6OBHimm3JA/wwMkC7RMRMI0
nstxlLecaY7HRJ+INXUdc4SJvFuPqbMdIVFKoJuO2nPPcyi011MYQViNSI6L
j3G6pJSQFiLxD29pSAOBQF+1twSaNbwPJ64Fstz/IOkI40k+s6aLCSxe2nbL
JOQwfZL10rGHuj8LiUF5zk27b2bBCYULYJVL7oaFaQ6MVXGvp1Qqv61JCtV0
4Exw9hAAS9ogTmHlDjBcV1ZheaMUuLzoqKqSfuU+PHTv70PhJ0ytmXBGzjV5
7SAwQymzXjuc4cbldrghVedaVQT9V++1CNrtIIwbmgQyHb8WPH7xaUq0Izwp
th/VO570/aMBxIzVLLfrKSyH5hCFR7YwXjDyv3Hp/eCqq4b/rJCoLnxYHwd8
hI9ay6TSjEWMTuIjOGJGzLsHj6I6/WJadlZQZq7lzMn/UG2qHkPtbch8RQg0
uRS6XtRdJxVtNsicARlcYvN8XnOV7vDcKEnCPPLipmbsW1sHy5oYkIqzbvt/
97EuaA96Mm6p9suMxS3pntyAYYQiTMLtnRNJR39mav2KG/IPzJgpYpA2/GI5
wPxHjuUgkeeppetCiyZNAQsotH1utB3LPb7qdpCyAhY0HtIMnwDazY9NNvd5
CnnaZbfJXihZGjavmnWkoGxe3fRY/H0M9wKP7HmiOf88yTUQZFtaZ5NK1Guk
XhUKpd5F5rUqQLs7DegO8obytCsM9Rn9vZIhItsXd89E6gR0rdAKnvYWymmf
5HL/8t2AhQnjrZdm3GQHi8jc9HFmELOpJvz46g1lwMVmFPr6NFdO5OLysrmY
DeHk8CCN7cn4RhAtFqnlmm6+SXQjo5nQxwJNdgipDVsGH26FzL0JLSLfobHc
cTtg6eUGz91v24Dwp65kz+ntDYmOOVNZ6KE2XOOASJOIMqJz4kS2N5DNJ06k
zREYEBvid84PIkDTRvDKPxe4Z+4PyHzgJUDhAYEM0+NeyybrVvBy9ZC0ZhNO
HcXjuVTRxkf3T8baro6+T81lgpDZA+L4RkKcr3tqnLA5ZZnTJWCGs2e/LzAH
hDnQ1c986/pk7kZKciukyytR6g5XDQTZUyLXIw871OL1ie3WXf7zhLTZMkX/
1TaPdYAkFPiphSOlGyxI2u4ApMaKU1eHi3HBbdfSlOo3/XIupge366dSqBfV
X2IujvUOCHs2ETPSgNmDp7POIXMoMFirtaqswjOGiaxiwZ3EFQEOA1lKAaKU
5fGh6XtyH9m1N/hIf25JAzxVnchR5cxoBsQB5oRdMythRE7JMfuEg8++phHR
4JO/5jjnXYn3hod0YKoXluAcmSuRiU4aFtPs9sLS6jh3c+OROwpSBxFhOfhe
GqsQB+gej1AYP7Jc569/rrnbJ+1rUlq4H6/8JQw4tNZ/9Ll5jfs0NaqZXlem
cuG/nGIoEEvfZt++75DQN4FrdYk5sRSWy/hlENXpeFL2Ux/gzRuuCTHFmEoK
iI0/O6A34TJq7l6wnicA/YjXos1so9blM6m+4nuK8Zj6+FKR6izapVayqXjJ
9QGvn5cdO+33dGRswRACa00ia5qYe3v/iVYOk6rDeX99hNvuWPFyNq6SD7XE
yPUonGubhHhK+x7Rbl7ls0UO7zbnV6snDj4Kkr+XpSwud+faCrJj+Ar/D0SO
Va2G4idDPZZ83a/O7UcR8U6hPN9oZzWQSk51YaKG5frINfLJKe7wMwyxihef
fJ7wTEjK8kaDMc3M3XbPZ1DaDaPbJqluUhD/x2op76e0L7RI/VjbR6vYvIgS
ogfnR1MuQvAPN8IMLm4yNzsWVGFJiX1D9VdymrbnG3YA0s+xcCITdUVoam75
LWuT7sWDLEFcgpdjUwh00OBRcR52b8At7emGFYDCEEkxrqP02sGVnYYzDTI9
KLdEhLvde7DiR6lEY1w2J6p9g7s7MClRJvgB5/JoL6KcAHRUmBQL82bgcR8D
zT6H9n5BorS2e8VhDfw1z7aQ8PxAYfV4fda7etFkeXi6ZaMy5pmNHZEOJLER
ZlklMwvOa6OxNRO4w+uE9v/x7MrtQ8rCpoEFeXPs7thQqRRHB7l3SSOs+u2E
DfVn7+1W+nFPhI/KN5wOWFNfHYy78tmJCosJNz6XEZXn/M9wqE4cONVzsxza
ROHsmKOPU4UzZl8KqDuzqoUVw2xkIIW8OZn7BSOBAN8QrbnmPPmhNryQzVx1
B2zBVCcXbubBqapId2e5HG4QY1mRSCwSyzRAmtdtu1gwnopwaNTsIGspe9AK
I0qYL4tV5TX62C8Ob75xWe1Shl1jR3JmQ/onDL3VcEeX5EVebTEs99y2ueTR
4LI34VyA0405s3aCBN37hxINt3NPdJR39cWpq7nAVHKF+0ptnsxg3CeDywQf
Bpru0+GdE/cliwhoH46H2S5g+1weNzNd51aNMsUHo4enqpjxc91CWQh7cVqM
88V1RTwt8BKQUY3M5xb9wFjiCMrIQFkVLFoFIYGTa8+toq+UFS65y8dVkTR9
OnQwYG7oBQxj2wF2g7gscsOL292KJWMtEMSjpT6LJ/OmJXngmWd+kjoVf5QH
Zc16HtMg8dQbCwKZmuEPz0TpwYuM2bXkM6RL6p99sTCN54hkXiYvD2WgrXDf
vrzybv3KO33JRPszYfZ/FMRAKwEeOAzzlZMhak21X6i8U2n2kHo++ao8U6bx
wG4ecvKHEedxtKVy5DdfVUTzg0raG2R4hrEBrWTTl+ZJtOZ7LQJH48cwMp60
UMbbPWYMfl1IPWSS++qqXVPM1ingcP2OGmjfFhGhlm7kI7saamdYirMk1Bf6
hgQSzsEBQ0qDSimE0MMRIdwWEGOxCTiJVmxtE+A+PwxbWQleruelgmL7LisB
//h1EAwXFD7k3jM9gpB5KbgyaTLQRnOYx3RkMsPovRC8pq+HrIrU54CogwPX
ivOTeAbf0CiJhvKXay69yQ8sSwMpp1hmD9TG62SoLqgMPm/DSoi3f48uUFLU
TqGqV+7B9r1uvP1QC4D8kabyie3CFtggs/KcxE5KNhkVmlNd2hr31BZfN7So
Ece/7o6jn3nIBrPXZkgE3s4xXghWh2QVE/KXBkITeeHWkN0vVPiVE58NMQO4
uw8h4ydSCZp0NXXa3Ap/lboVx8UUfVJ+ZJ8pUBHnn8Tcjf5X8FkofI+Ux2AM
uH84wGMfHs4wnqZO1NwIwA50bMqGaffjvepbzOVkO+OlffWt7ha6s7/qPN/n
XRAAvpZ7eVe3DZaw8RHTk7LPKHexedgFdOY+T4mVsI+IBDFoHUMQRVYa8XPy
SNGrJsLdMqijjJxflX0mqTUuyAQOm/sO8SGHVrQS6mYjC+jORKnsIT5+k8bB
6QeJ5TcN13KWkIc5Ahr4+tBKoeQ5hYUQ+3NtPLf+xFaG1PySfJ2Z3sOEuoO7
A4stAWzhGR9Z3Au8bePrb0QGQaA5kUoORfaHD8b7Zfe3XfEF/D1xqbIA4IhM
AIp9nfUGBE1GqNsfWYhupHA5/TCoJfOYKSDgAeVKV8eSDDRFvQmWhy4nNZJd
fOF/2vf4dBzlUA6kbi4eJ0BDnoGVvu8jr1WJ4Z3tlYK6PUhsr9gmmKsivVqW
Vch+l73LGRTtJ0QfCNs16yzaLEU+zxwyqOEHjm2dlPra6ymOrVvCTSweD7n/
ZtCmGMvauUG5zfF/9R++Bxt2Xx9AMB+Pc+RFK5ERKmziX6OD5dMxmNEpQ2Yn
3074Huogkrsj1WP0ROEu5UUr0bwDW+6B4uTpkxxSjPjGqomD04Gcr3isCkJ6
EPmfHAUr8L9qXr+AS2nOOg8F23y5E3pLvPO03cyq87bhI/iRH08TcDstByFm
DwIGrmOLVvMF4Ola2J1Lmkb8cAEiiD1ITzrcE4TCEjEZwLeClZbSk5bgvzJC
8Fc4+6VtZ6vTfd40PnCaB+RJSMAbRG5KeRgxDQkqvgQ7Ub6XxbNWLDhW3u4O
0Qru9zuKc6a4JhhGwagExkY72EHRrgR0yjjKg/mlzuMAcwIXTSSWs4bvbgk8
bZgufGhF5DMwEiKJQpQyUHA14frmKRjcA3bm+M4A5eG9tVZee9r+nhYAZFQH
5un9idN4sS+FlJyWvWC88y+Bux2V6BM1p6kz7fQv5m7POyd86gImx3CyTHy6
/JFFUYLzxaxqFCc9nKXDN55F9w4Dax1eBe93m9gJHz4gLVn9PGhMuw+3JS2T
xNXRQHTvIQ94uEeT9QY3vY6H12u4p7ugg65XUia6+HdQgMGSZ2OibXtOV+Z4
KySq0KbK6r5EA3KVBgGju1sK7U3bGPuFn0tBG3nbUwCPTZen4bd0lv3U5LLU
hEK1NEyLSygaq9NX8m2z7z6LHEp4vERCGQWsFfTA94XXTOUWWtCDPMMBM3jm
LdG2vlh271jFFEC0wxxYye9XtQFwaULg3SjK6jrt4tRz6t7iZwwfB/xVsngF
yq+3PuzdKkSct1/vlbhrQcBVfr1jl83ACT9UZbX/++EC+pBL9yddSGk+Q8rk
HYwfEeD9nDS3oH59D3V+KeTnvbEVC3O4U5KljD0Mx7mbKe/Rqs9R2Fx+ncXB
WmBughRywvbflUO1TFtc2YFy1VSxzE/7n2ozoxeD0GT2GFR51c48x+nwslUy
UdRSA1hssmeVwQi3/LTI9VAHUj77J5R0OWvM3MOJUExbd7FTWRcYAizJLRV3
Vv8/jYjmveRWUA3hh0h+bVQ2+rD563BATkPKEPZ4AKWcb9rWsK2lMnReVDJc
LOMP0yM8YOybY/xe2r7L9DE5fYQa/KHlyM3Y3O/V2DcclVQpNu1yJih0wYGE
DR1u2WCDb6EKtcaOQZ2+qyqGzupwVNJ9gT/P+wiutk5JoOmogfbxRXvlg+Yp
/PZ40lL57FObjvVPYPXvEH3hL7RG1sNbZ801uaDikaSIGrFBnqYqpsUUhmA1
5QP+gmEOAjRIZvDhXRPRcUbc2FAkxk5WqO5lUqLYhHMIv4psM87a3m94lyam
SKdbmH0LIh1GBZqJOBUp5CN1bFoMaTw/VuWAM68vz5K7f2H9u7T48CZhybTB
f31olnWLGEiujQ17bSB1O7BORMHk/X5Dd3nG7e/CW9PHvA4CR3Gsk4BkUNrT
XagndYWGTk0zM2k78bUb2weyu78EBeLrjZnEnNvUq9I27HDuMw0LsFNKmW2K
qJCYbNNMVZZsj6ws2WFN+dtUuDhBPQ+YRZJ/OkFTQKJjDTYsfnQY1hTwRI+p
MY8Jmx4cfQNvqZFmjLdeL5eU6cgmh+2Flza3SeUos9s4mG4E/FV+SusNje6w
Q5T6VixGKBqg4dsKuMRk5zC7Qap7TaD8dJtV8k/nSHPcD3moYTHK9dZ4Jmd/
+LdxBSDZbyHtmkGLjTbeNkzzfqvvID+jNTwdVdF+K+l/Qk+/nemrrWno4/o0
rf4VJ8uUjep1Eyc5A18W5UeAZ7AOGs/VvouPzrOMIk9Lmvx8Ylc5GJmtl9e0
ZvQ70V/nZ9JHy8RjEoLyRinLHgKxkzpkUI8WhCWrMsRZUOXeBGI879BUhe3w
ucyi61rFQnC00zx8oDu3CqCZlOhLi1MS0DdaurirmKDgnBHJA8bIa7+N8lr8
JkkQVNPsOrZwfmeE8NHt9K8lyqb43aNo0IJlIx31YEH8we5glM7ijqmfjavR
D4Hj+n7yJXR7tSUztZpBJkd73+yJ8CVK15g00/Nh0p66+rThdH5Hibm8oL7m
RWn7NX9ZAMvRJsKTYngPj7C+Ds4t6SuKkw1mH4hs5zkCJ6jmgT8EbaqfNHAz
PDhtrz2Yi9Rsc4hixH3qcC0BpRLWJiLEAqifgR7obPixHSFJWuphYow29Bov
8QeVv5tGqePDn5ppR24ZtzDqLxLqWsmsClhiSh+dNc4IEDI+F/TGhmd39v0Q
aynMkIccfbXjUCDWvGDDrIb78eYhEtBLdpDmcXUZILQYhJ+JLbdsTiKfoS9T
gXBD8YWl0hNJ3eCvEJ5v4Fl/0pdHkwK/4aAP7RT6OrVYT7b0m29G+J4r8bT0
S9vGSquEQOfL8z1EQN6hi31qXcnFGaoSirIouB8U2uWZYRaKhAEaePX3qEwU
jYf9u56EfdjhAVNl1MtnKosrHMfY5r/GWrgNIqKghx6t/yairCRenutGtD+J
V+4aMWb5PFtP8yQ9uB6G9Sz1et8Xf7uzEBODOU3cElHZ/27VbNkjiwJ9UetO
iEw2aBSOm1IVm8dgqcgAM3YiyoTl8w1i0Q2/vd2HzqVVM09hpYpfL759qCnQ
89Hk9IifsyxxqwhkiX7E6O+fIuPTABOai1cppX071Hv5vm/yp3oX3u5RqF7I
HBh1uy6E4WjK86soS8KBGlCPiyCsw1HJuhtrEC3FJSZK96VzxKdJ3Pyvc4Cm
cWjkF19LjiuVGBacRe2HNqwlhS4w2o2ZmFNRCKtjWLaAHPX06zYmvQNCidAy
YQKBvpYiHXPB3BpP46l9P/RB1X36LULeJCgYKZ7sOSRsnvmDLQZnoBNra7uu
ieESPciNcW59q26YHfq6iogneIBa0w7Tjtci3k1qrlQu9NvGPIhIOhLB9iTB
G+kr/SKi2ieXsV6tdQzm4kx3QQ/EQaHlo9msmCdTMYA36GdOrgQKv6VISuYA
Ix2kJd4Os8DeRBW77lT8dclUX/pOCkc7gQ8xo/yLeP/p5Nriq7bChMUtsITl
GGjO8IUOPZRYeQg0cr6GqE5K/JAMGKVgvxzhFUuCW0+DbkFMzCcYKp/QBsCX
sweTqqOIma9ZEcyPwy4R5UfuqjY8Wcx0A5316/R1QIsCp7qhMHp6ye2OFfkH
Pp9RiR3jUHuz8n3agQvFVQI8RpfmlGaobESlQdhQknimrC7XUIWd8NM2TAJu
u5A0J2/qnA8NV7KivngU+6ItTnxcM/O8R2DBPtHGOQNWDrvH0MRLYC77i0ha
C7nk8ikqZP21M2/kPj32m4blLS/7eTwuis72jQzgi/n6z9EcYzZEYq/G1zDc
HBpQjH7QXvmpQ3aS4wq7yctIU0uAzRA6AqODlOq5lS9GpiPAdPMRMMbNLcTW
nvO0Z9kRM10P5pGP2RhVLJ0+L5S7wQvK083f06Su+Q7VoDUXsl2yepL8bD9I
TQAugmjQWRnCXAWbCIQSUgvWsBVCvaWynuQP7kQPcvsMGndpM4uUjvLUWxFm
YJd0jO38l2v/sjItpSPgSG4euinLRLnGzGITa1UCrESiFtQGvXvN0bdsnhVK
fnKnO/FiW3etLoQTrxQduSnBl2HjwBTbJ6ap6A6vt3i7PW+NANjeRw/v+UPa
Y+KGHVgp/4Nw+sXFFrEFACkJzmaSLxntlG4uDqVTnFT/BM4lQOC3CcgWlled
Jw8ra7mlAJMLhbvr79/baj0Lp8dkBMWYQTRytTrj39OazktlG5n0hEkRkUcF
QwKZCaBHPTCacZrnf4dexxUJzlL5jF9qq5Xd+EdQvoy7oqr+SFPh96tlmH7R
/7u4nwOvnR+DFa24jtci2ApGZMhO8dChF1g6qshC0ZtizsPuf0pgdzf1T4UW
5WP0m4vQbmoHr6xJGApPbZdG5ZwQk4089pG4S2nVPqjbBxJRvC5iRjglCSKS
IIh9TwKDPLnO3dd1HBgR9Oho6+GcdTzmpSj+dkSt3bPZ8N6g61ozEZRmkmMQ
j0SoZ7ZUJBrblsBY1PPdNaxhDXJow+ECcEkSVdo/p4OVSwqIxSf5dNsWB0rC
9lF0lqpnpWtj/0FsUaPAfw9xcDWLUZvUtIgeStIjogWecT1RrDQN35gJCj/R
U2Nznf0VNGuZse3xbPkmNCQbnETULR21iffOC6UEIjG64U+I8NHwcgrkBmS5
WqGbhfpv8LiS6lxjVeWEIES6m4i3XICpHyblg/ONZgzpxaZ47Opy51OkjGrW
LsIGlkVi2MRXex26bSROvXeirMqmjqwnTLY1xLJcw8JsFFGHa0/ZJEbDtWY8
6JxrZ8aOGXIuNLraRquWsWvJpkGANJiA5DMIMghhhiSIMMf5QWGYUkLCkxB3
VJa7frD9HTkgw4scp3fUKrhVfPNhA9G8L68QW+PzkIhvHU26XnydYeA1Kk7j
E/fJEBIIJPHaawXHo8ah6eRVllcqJBwjeSsVU7jW7LSvk6EMCmfeJReYttmi
WOg04Ns7dnBL7igxUxhkQC44t/sLqKdSJePbXKFphexvMYO/YvjHSdfN+ngr
vDO4MKHs16YSXCxulYIZQxrYOXlVm4apygj8j+xUU9++m+OjNUqLmE4GjsTP
Cd/yTr0T9NCqghbWdFhwmZ5Hm7jf6Fjw2zTe677P7JMV4g5LT7dQsmnMy6f7
pWKFc/dR2N0v31Htg/TGXCDm4X6EOlaXqOb95M70rxFZCYyr3q9VPuWSHZUA
dPBHhYqCDYM3yns/Myenz0GetkGo9/B+KjqBznTYJDwDYHd+bmzr3Yk+Xik0
I+/XbEcRD93NqpTsMsE2+pAuoRPa0obiGp3m9B+EAa4cLKKD427Yuc0F0ar9
a+5lPfzxyp2Qq6oQBceebs9AT6pPnEruNeFSVTREMSET2kAE9buN5FvqCSx8
196X3V5kYxqKjdryu5tsYccSEquqsFreIMga5AIth8xLpugnKlO+wt8MWlYB
yNBfVEBIEVEW5Df7Vfxh0qRpLKg2q4zA6V/86+MEj74eJ+01mV7xmK58X4s4
E6KyFVIm14u4hT/LFe9XIWIFhOsaxrTCmllKWF4mxa98ZNSawLMkc8v9ErA1
g7YLO0Q88d6wmg51BGjeHjtZzel3PadE1SKiIeDne1j1s9199J8BRaJ3O0a2
dJqZ7a2JRwB5U2KEvhVQTrepNaYpoE0v7wMnBdgF1dunnPuavIUfC9JPGWRN
JrLarIGZb/8vMuB//W8UCMqwYnAtIROGI9h38ok+oNI49k2cPW3iqArmHCA8
5xVsKc/5QHVmz1kFjIjNncEeyAi59m9tx1Bj8/Xj/8mFRDpuYGdiqcUytgpy
+vgB7fNy89LayPnp1jRoeKbDbV/t71qh/eJD54qKjsAC1kSc7Mpq4LmlPqGS
RWmhKWlBc4o+OihauVPmGtqjiZYLgW1ng8/ohgYY7ibAjzFuY7sXjvDL1iGW
JC3KP2S0hCLqMCfFrECsMVwPCBb6ihhG3ngHARJFnIhSnjdA1fTrLtEr5Pka
2AzVkqpiWKl1g5Ejf5uuGiZJzImPbTYvHmnps5ld6ydCDm1jWsb99z2dS7f2
tOkgRtaAFRMkumiNkIrKraFJH0OiEGIRBdilZXZi1DtxEhruyFh+Y7IojhSx
mr0sN5mXlcmcsw46xpUQw7I1jQ9+ipH4q+zSGR70hSb6WKQhmgAZpCJQaDVv
mBpSXzLbjysz4ifMy7cnoZw42XFGuSIiqltjg04KEcMTWcGsSusz7yez4rV7
wVVBLa4WnRgD+d/W9ns3/QIXJtjkAJtvQydj+SFlXJvcu/5WcQBE5N8xn78P
X7wd8EtujcDBuN8a3VeFYgiwnIpUtcj00VeS7Jhizw0xIiBMcWFrHSlgsENd
u7rhLgwie4ySgH+YbqPO7upD++jlxAOuDUcaBSC3cu7LRKFCY2ZYX/jQ1jh4
BiAShMdtC4RscD7/vmQEofc9IYuqn3srFFEKqb+Eip0QJNSpwGSe5Rgs0Vfm
EbTNadaEsF4gq9GaAZxlAX1ptRjLvYJ5BHLYDYt/jjQsGHiKqTLbzRdY+qcX
9cHl57N8CwmXcBq+klOo+TbbAat/mkt6sj8Ok/fUy1m1GQE05m5B52oWrUkv
jED/RBL1anFW3nPkQknFQ5UfGoa1U0fKaEcIVTuA8nj64mlMvbBadot/eivg
MiMBt06jmh0KCCr4TmXMyShEAj8TzL3+yoeV6/3k+i6k3gWA78PPSC5XAytr
9GR9dIdGbRrMaQBuWYFdPQZqHPZxFE5jPF7rluf14kDZNlN2HoR3ad/JUEmO
gfEE1xTi+f8otO2KR3TjPz/H7MAyxa13fImqyVtZ+V+olyOGcOY6UC2ztyo7
E823JnlpeVxZA1tGfoGp1eWynzypEBEGzGcUxEGkiLjp8dBk5OUVUcHPwWmB
Ujl2tHCZFV56VecBq7ROtISN89JoS+4Pb/Adl+R4zb+VMqymsCaQqfsSsXTH
8iSHeFYJIlJ8mjMM6S3eSWX8Y9tkjmDbF6/g4Trm3QOFCD6G49g/ZIEmMOXd
D3oMX0ZOavFD1PiOdVS694D898gdH+veMUSjZ2u0KHrAUkLIlsPLmVWPyG51
7hNSUz1LrpWg9cyFSrAPNtU1+xb6aEvaOFanB3Xfk82gZjzJgs/AMp5w3ukx
OhWon3wCuaSFl+NuRxeMkLJm5LMY0emvD9Wqug5CyqkEg/5B0OVPHiqruD02
BOy0R4+XmRL/3IFR4p8Q+t3plS/GngLLYVCBL3VCTqd4KMPHcQ0l+My5JF8J
vfPJG8/s/oFhMhOq+Xhukd6M90n+FBN+L/QN5QHc80QyASCAdHSytJSdAyhm
zktWW5HHBb6b2RkEZngngXKbGjlFHvh1FcDHtcMk2RVL0NzCZCdJ+rvzWq7l
U5b1wYtuxxfcjXdBi4o7BNL1bISlABysl0EoIYGXE6k934/GoNhZCjZ7VhpU
9ktp+32KWIzaHHFSvxAWV2uCTc+Ak3sk7k7ATtYCERzM0dikauUFi7eh2UxG
dKLaBArPugAwrbVmAV6Lo54Uj0ajFdm1XOEOQ2nLrkj/mf43yTa51IgY0XzI
B+O9wpDpzUqIIwMJzYTXvNA1iZUnCAUtkqNlhS/jGSTnnzX8X4EkA5pM/Ebk
JRlSPA0d4FvYs3RvoAp88h+r/XVHMULDgIbmcyLpnB9fuVniMj//zT+XV0Dh
CCNzpEo9NwtH35iB76ID/+pHWGWMGmvyIgb143+Tvhvu+vi1eiodr6NTnB8a
HsR+ORnRevU3WiGGXSQSrEbUh5Vqs4VH7Szq6v9mFf+p1ARqIDylibxT/tHn
FCAJxszM4jfMGcMlTugt6aQQFj0PzURSLy81FOzz+6pWWC2ZDg+6PeZO0ArZ
U3KtF79Mu6T9pZ5TVWff2LRPtfKRYHe1pTkxhXB3t6RKHLMarUZsoG1KHjlx
NFw3ZgO2LgMvqngLjRB9343nIAi6LpxGBogcoWhVJp/s8fHCadXYh67/QxDf
uyPS56CTnTzsQxrEBFT5m+Y1pkAyzkKMgQABLQi/hbGVOTtix6ZZ79zlAyyj
dLMKdttNiKP7TJVjQkmyX2jnVFAw5reGhvungBjYrpY8QRyKPupDwUX6Y49W
qZ93nWgCCXqmYNHkvqrC0KCdWNbTEIiUUU46pUBx66IRVQS/R7PUPusTJDCt
khgCT4wCgiHrGOiUAO7Bf7m1SqEFI5jz3D/YaBWEbzOyxc1h+iCjWeN2D4s0
dbFIAr540NuQm0jDkXYVOZzFdHfZVSBXfdld3hGmzuwTnXHMXFFG3D4ggRx9
8mp5KW3EOJYrS8OfUXJexfA7ftGg3pBMdrFqmhOICsPKTe1fBlqfk15by/kd
WpGtydY1UGvMH+vrl6Rto6rjiCEVQVTTG1ysX6vT0B9sMlWxvJhk8UHY3x0m
VP4a2l508gNGRI5HFj9kGLYPnSckCqA5Sig54a9tEP2ZqfujAVCQnor4gqG9
U16wrQM/nqjjE3Mfw6L1B/wNNUdsyEnSRw+d73u/klYCIkX5zw2QfGyhUhOb
dG0pDdB8xTl8+nco4LTdTPboJXPag/lEQJL6L8hKhHIzFKjVxAvouduCUNCs
iocXw/9Vsrnhh31VR5PreyGFNYZ7pjY//sa50P/VcEIvQ0fe09K0zgLrd9zM
y14ov+jnY0Naz0uQrAFUf8KqlSRmlaOkIILsbrDzKkwXPTVzZi6DSmtBt1ML
sBDaIc4kOGVzR6N3I53p5MvkCQMHISgbg7RNMVK/uoN93uNSn2fnImF9ocJK
N1/qL9QK36rJUbpHYVip/ik90deKa+4aGuypb7RqsgcDz1BH8xQWn+E5dmit
YQAkAY3Vw6h6l9dZJQgs8fcbJtYzCqnFU4GKqCgvBN94OKLy1v7o/X0ps3ZE
R68+ONt9afU092OIRVPmDIi9ZZpZTjXpqO9leVLXp4rkUHf1+8SA7uDHoywG
6nEBi916mvP5R7V8QKrwyafzfAkvOwIID8w4o1NN7f3+olL6TTv0xsA3zlJu
p4tYB2X3bNP/bae9r33ZMBJdkznpe1HN/e2AH1EwfO9NdXJLki2ihwjpammL
oHfA2DWqK3FplV/Tdvwak2kgfRxq3VrHg1yJgAQf/U+sbfZLxhMUe+t2AuWF
c9+w/HWZW5XX16cdxMzrXz+6ZSs9s5VqF8dEajEIans9zSaewGpKVJ7iY4pA
De1YY9hepZgM+C7tWkcWZLA9g1o0qU41iXX0wogp57iisZlriKVO8R3h2wRu
KOEVatetXm2tO+k/NF56ekRR3+9e4ya4EbhyKKZJ6HjxEWJrlWMWy3QQY1Mc
KzkGy5hM3thXKxNMdyoINuEVcEEJIir+Iyzy1AM041JBMfX2qcd+4x+CfUyU
nAqdqbnr0Rq64nNQYTHZkEtLb4+Y49IS1ZYAdzUixrnnEoQzRXQzpW3BBC4C
1GRiQu1KTtzd0yXsq3ecMwxLQ/00TmYLraOQNHmmIs2tZ0Q7Ps0wt1DC5HcT
uRU6+dRm+G21Kx5stSuAs6GQe+2Mqa2wmXX7vWO/4mlw42nwZp7GLm0LfRQh
DCK/wWrIja1JYrzGfEd8Pq5ksvSXCLKZhPWtALPeAAHlNRy9/1qZletimQZ7
ljuPHcXC/AkN0y3l4GKfCd0wR4oRnZ31Kl4FYLtBufEtaV+B/JnbuRgffwlt
MIq8mdChtmDI4NoiavRtQxUE72NCNx07g4oTFSdu3RtMG1b1m5lO1wnNwzTp
RcoAgELnhycXyERzsuozVdN1dloJuCmgOnyT0UYtwKpBXgkei2n0nHWxwuMZ
2pYh4AqFnNmzWe65UzMAyYIAgKEF3x2f+0s7jYaRdcgdMMiO+ZKa3+CEjxTi
p8ic/m2pJ4weB/JuB3qN1LVemSCW5CKi8pdN3sQjnKAgbjJNhAaEbVigmQN9
dJbW8pAW9Ju8+Hkx6Lo8UhfdZvS4hsCynDPYv10rDqwqDus8Re82omsXs8z7
Cx0QXQtBZiT3bTTHEvj1w4OUSS28Ag0k1LS17RP8qoqBvhcD5eJV/+a1qzHl
9jI8bi2KtTPEEIiekJx57L3GC9v2WAwf+M47rmLZKrZpUa/SY9gnS4hjiUDl
2N0cEFgSkXmTlv6WU5x2aEQxrqNMkePy/YFLwJMw1+FQ406roh6ISKXyumnr
wTM3HinZ6aLuXFIv9SpauoXRGCey/gbAqX5zusJDONgZGaRuEm4+T5O4vwPa
8p5khtcy5UwbRoAvVh2vKtJFpUjN+IvM1VrKY8L6JbCIJop+48/SbaXubifw
zH2TGGEd6buctgY11VjWwMCWMHsVWAC1D3PrhtsAVCnrrVU7CK+Ra1k10801
0WpeqZyB64JpwGSUPR2e8p19aXhGJiYkzM7+HnGiThNmtCMRrZatxtRSHIPX
lUQGy6IWEVSowErTLbNPIhvSAsYkdMAuDEEHDJaI+Y1ehRy9MFWlhNtpK3rl
Nv/7gZ12u7RqX5TOn/jVnC4okW1Kl/p+h52Th8uzxcTXnvek8piyIxKCOZ7T
y9zWMl+hxMkg0ZhlhbN3HCvBPvVoNT0Mso4tRqQ4mKfsvdXHJn/IQ3cVrQDK
3XxZRYBmWzyo1G4jjjHfmHBDwE3KPQ+YXu2A0aADjiFgzuzrkXY06n5w+3g2
J7HU+YSe/3ykkie3OuyW7Dcs5hAQIPqNXNBCuMP4tUGl/oWFMfzcW9929McL
5Eb+ihK85s7Lw2yTSYgxR+FDXL1Yx30zPn8MaM7a0pBGFKuiwJyOF0SII4Vl
3WCg9/PHd4SecvhvLOJgtitVbZZSzjIQt1fxcxSv8xGMdI639H01/KDXJFTb
ha7RrTZjuJc/peTWam9OK5QdjgDHqoZ29hqfhOl1Y8Gb/Ce+HloZ2cLREeb9
hcVjZi0UVD1IEooqpxlypRkXBVwsWsINTBs9+GOKyYZyFqOsZtdEs99R06W/
39evoD9kdHxTAHF8I+0LKwDZ2oU3+L87H7AX4inKcWSzPqx2ztQtFKv33jyc
xn6mFf/TysAdFw/tnTQ7D9aS/udxqjr+n4ggmfnrENo4Cz3RKKZgpJeFc8YF
QoRVmGyCVyHvSQSVJruk3TMSf8A8Rvi+SU+mm7IGH3tJtLib9zLjVOP1D9ex
74Q8nlkIOhk11wnafRPqSKftmk+VcbAI2ObtUsnyV6eUCjOHspSO6ACk5pEz
NjEgQuAwLQ4M2clRavDV8kwvKQv2t2o0nM5+1C4VJ1+tZEwBdr85dI/5VG1u
fymy43d40/0lZ+qoWo+r2quJbf/Mph+prpEMPRPT2zju6Zli/V4nzFJ39X8x
xxf3w3Gvy3TtzqFEWabpo4IiL8ji0MZcZjH8Ndfv89iXAWO4fpEj8v7oHwPV
JyVM7j9nUJIjba9eP3t1uA+JA9ZT3Hf88e2bqGE2rwyR7P828PrEFDRpKBEy
86mOGhoW3BCLxzg6Zy7/BdSV0MVhXulHiS2F2sDaiVf91LQEqvmDbvLWlgpR
pppSSM0cLcBZqlPgntWUSBlY00CgWXFK6zx3DjqqfFYHx478rbgEdMXY/3pg
zoTaZRlWi3tK/kfPSE7H/jrcTRIwCty18i0zSj6PH8OAExlLRZhOVbaeXl8R
qoWY4ppcfYA3woYfwZNBvJ1pJ3HjXHAJba0lzcNCeA+KZaTe6BdaN0CN/6ip
Xoe4Ihete9ZzCw9PV4u6g7F2M3ve3Nd4GLGcJQO/FI3dWmN2gbyC4rGm93jo
lKgCjPnaUf0IMZZfhXjhD41HzR2/WWLmq9Kgml4aWdnCPjJDfJa2iooNDOMB
m21I4yQSbgoyd3DBucIMzkQmkbpWPplyGZQCUtv7innWVZivOl7LHY8AQPYC
P04/qokN26SlslkO/juOsF9mb5VSn9bo+susbs8NofGYvXSAFtsvyoQ6Nmpa
GrZ6EFmJU7MvdDRMnKRDlNRR/FoVn2GDOLLXOZjGBd36pHER2gom4hhF/i2D
bQHJXBuYLEoxxxk1dbB1ycUcV3j0tFuNEXiM9Mkyx5SzLNxswGnSGUdhDJzO
sEO0DG0tEUP7RiIG1UisZb8JNppu82ZPKJs8RzIVsQ7qf9Uw12BCDUVTWbvA
InQ/vJ+y/mbPZfi69ubRWcN5+4COsaZq2r6OY6fQ4xflp/IT2ssBuRqTVxD5
Uk6DnqR7PBtHaMu12/34Y+Ocmw5JAz3ZnH37W8+PTdSXWK2wKZGnE/SyCRJZ
ND0iMF3Xsljkw/iF3E3hunWk5zzQ9IrPAQ7RKT7Xhzc6fEe58LFGnQqhbHy4
QK0b5T8Xep3XqgaP60avB5ayf7vHtD87aUfuJ7/opYh4pRHle06Q2q898gwM
2FqDkBw3G4V7LZeMFcds5GMAOU5FgsMDR9vhxzXEM/2yYYNVAkVmALqxjk+1
mHhOoDAzqVhwYWS19sf1/zHtKO3GKK9W8YzP97UofvVB463A77SwbOuH/h6i
Jmy5kEIYOKRPS2yy8Cu4EYao1iwzXV5zO2nw9j4Xse/QMrm00pPfHGNWFwnW
7R1woSKBa3X7Fo1dIyCNz9jl545EsscXzCEULUpDdQQkbMrpHLYsNbQ8KnSf
Gwb4/dNQTQHJ+eXBw5blSwrCI/PsLdf+s27GLsoVhlkwK0n3lHefFvDrrsX7
cRnmMoE/I9N7rjzMiE5cigruI/QltcBt977mFTKljh2InDpdY00eBj1lx6s0
iMnu7gGFpQ88qciyCVYxmUC/fQuN7G86wtKFJAZigEHpvjsF1P2MwvZxNsfu
9/spDFWhsZR57hyA8B+Xveky7n7+Daal3zX1kEPATbT9NZAEaHzy4yPJanpL
95D1mHE43QiBQJUivpSi5DtNpxDKwhHW2dKdUHt65oJr0/KCA+YO6inIIL5w
Ph72IGpa4ofKLEz7q7iZh4IbndSulBxQ4EO251idJvnB0C7ZKlWTkax6fzOE
6LyR2byPCGX614n19oB7T+qwHc1tw5UEdR//mBp7ijV+Afmf8UUgGMdiOuCx
wHnBMNHdcC4RTdGG4fzHmF4PcGsyPBkQdsOTmNSeS0R0eRDqaLHAueO27ZiH
/QMEL34dXqqZQM+jMepXG1Iw8pE+GiSbs5V+i4t4INmHPl8TCA0ENiDT1zGY
sONlvuFjl9nx9UxyPcl3J/UTYB5lo5phv50VNIZIcoI5OXdIRNjjpx8knKQf
pE5VjqEawuAP2O6i5ugNpTFuA1HEMUk9qLyYvABgJOHVMy782rtRpJ8+IGEx
k5wO/HRGb53zylt3eVA2hEPviVu9/PGfkFKidrr16OnA6goMfRB1xkdSqt5e
XszqVUkIOQXAbrqhaWAdxgGd1oBb06JbJjXyRHhWADco+/cCIjibpBAQQp0w
7cFzrj7okmYjkUc+RJrxFtr/o5P8t17GoN/4YsqiTch2D4qJrl3Piqbx/oO4
+DjL22zmPMA7CFTdcWdwUjXPfEfMCxW8q2/qYdO6sg/F3QggIAA5Vf/bOIqH
UJ8pKn61mDCNZyv9iXhWfMs02WzIlXCbpniUxWV3QTyHWdwdn61kGfgYTg2M
7/qmlaX1qR3KcEO9hcO+qPaO0hjSGmPYFgcEzzT6TAPf+VC3lh/nSzZLgkBB
u7F++J/nJqIPp7gmDSuEtOHKkenktv7At+B7EFPAVrLAzSoHY3UdYkk/kcjy
W9pG/PRvIkctROyfoEbKEnSPjC3FEUqoU96sSOKHB0d2PW+blPMSxapQ4Tpy
jnk857hr6CGeFOAK6TtPjfbKBQUqqb2td+ouLMC4FAbnWRhfc5yocIJEI9tM
pBE3Da4ReUtwrtYE+4exG4tn8FWbMOV63od0OoYNt+7qiZEPmBwhtzq9xYXu
alVGnBdGmW2Tj1MdTPhWv4iD2DyIZ6Z6ZaJ18Y+6YGp7iis/bCVPoJTvX3cT
tm3nFGIwbZCAB21VBzVhUW6w68Yx4sCz2XqE4PJZjjUjm4iU7gg7Y64nyA9i
bq5lBMAbwRIoLDFKyOs0JxQz8yTRfhf3mBFKeHjg00SEs3UJNWpCh3KeE4cK
cHgZBTEEto3Q+nsfK9fuGw4dUKVNtHrEfT15IEnvdv+Z0vLlMlLOnd+n/SIi
+ENGS8NkImB600i2UH+6E205BaH1GXvS5hyXR2d9rohcBhuuj+BBdL+UPZAr
YKGWplFdBltMC5BKo1vAAjnm7sL9AO4vEqW2Pbr4nZsjbmHaqhVE/j8NqvjT
OalREjWI1lCuCZOAKjMFzQj9bQR8VEUtbpP7ucYGKDi6o3qnwLhtTU5I6yhj
Z7kPgXKqCLnKoH8zLePAc3Ey2WLeQeuCjPuXAUhT0CFlRcSeJzfKG/wkjaMY
60Z4KAswCfbR34X5NPixfM5dFSnKR6C0ljXzlu0EUpZcuQDpePGhUTJLtub2
tyHT0ba4Ci23wUaba9umDRrsBbgDiJY2BSWAYVb/iA/4ifo2sK0xH9rVUfwJ
LOzzfm7ljKkHNGsPU8VAnM0HLE7fCddRBcWJHQWnli7Dt0ZI9vAfTH/ZjNlZ
coW4miOiZjH/g4OBlFwDEkz019XkYwARgyNh13HHxef3iIsUj28EZwmQ8K+N
dtDV6So3hokhDemUSk4wcCjlYhFhKo1JSM24JU434LY1cXpR1TZoi83XJIkT
iNYkfvYTlBKgOhRb3y03IhJXO8ejtKhSKIAODzjdqmIu6GtSqn81kY+B2Lff
PhQGdHGhxZbyzFw+emrANyCb9rTRn+2gkxR+QKusE0LELlfsO9/JIcuY8UCB
zkNz9FE9FSPJRM6fCEYGdjwcan6lCCT+agNmp7wY7Xtisflpfylllq7CuMNq
YXj+1Y+mWtT3G2EzMnoMKNP5D1KF2Sz5txfajbn/E4vd0zFV1obaZI0ZaMXN
qFknJOZpWsVmK1XkZ+fFWnsJE/zX1Thl71obn+0GAA83oeNl4llSLiYzAFti
lMKqH6vaDYnYwqBKmAZmKuSlEusRmo3grUvCOnMxR8fpxhxHxY2AThnt7V7M
9FXXYr7nWA5bVjZdQgmQVPN96M1405wglu+J4Y+J3mXVnrjjXRxJLx/8Vw9y
bhr8nHSDDexBg8c47WQSLDkCS9dc/NiL0BFl1321B5wrVPUdM5udBuR2ni/r
2Y8m2NWfzpCpv1C8Xt02kUSjVoc43xCFURPDMO+pWeV0E0NLCiMLspUWHEg3
7oWwtRCKjOlSb8H4ORIkJ+7qLR858Vwnq8Fj5hmEKfXoOIS6B3vkz5k75+fb
EXWW4/02awCHRD0CNdyj05wNPj/+wn5vHIMtcbaCgcUHY+GdLkKY8/bksE0T
imCn0/WJMytoBdRTcDSASp5u70XOr3IVckzn9HtOtI0rzHGSUoK/AIJpoIAt
8LAlVDSRMujvHy0kp3e7Xmiw+u+OXW5HKd0NzleABV5/HE/nNjE45IdGvWn6
rd0hfx5fdMbMYuHgMakRLJweYI6wBm7B4ak3Odwns52xs9FY9bB0LQNHPZNQ
3bQTnUzG0W3vvF3D05UHLPwofL5DFXUW9b5ljpYTVd662Iei/CfN0jJMng3H
iibISjJgMwIEmRY3c38uELmAGQVA1hYwM1G6m3NhgDjoRIYKuC46nagCinu3
6QIpnFSiQWkj/gUuTFosh7Cw2tYTHCtrOyRCZeGRKSbSRvOrpf5gCTbm2y4Y
vo6Qia400ntnRHC8T1b3O4FUBqmFohzYiq3T/TDR3pNRYIzaLjO0pCKjEUuQ
HUa+BuQ+r3bGksYYXrT/lP4RVWclnyt8q5C9AUZTIkOqKO1k3khbY5TdWj6b
riFwpj7HUOb8TWnCZNc18cprJzRXGQqpJumok6EdR7EvImG9JdxuDJHie5rM
U9ddah7EX3jY2ZxBx1p1u/b7vVtrbU4pyj0sYyEiLet8KWwoJk4n14DV1ZnK
3WCAQkP3tZJVsBJjHdgKJ8hBkeq/sgV5GirVM1KQDoBGoyRVAd5NkGgWSL0q
zW28NUuvLZ7OMiGjJUvhlZowE8MxQehIktJU0gDNSgQAsSBd+P8gh4yjl3G/
b13Qg/ABYADDdtu3PdneDx4a1hcCyw/QvpoxhVOjrTe460ZcID/H3/+Anld0
gOIFEommWq+oalUg5W/7/t5eMbmhCOaNZ1HmRSW1eAB22kFKO8wNxT654cz2
4bI17Wwfvh/kcjzZV3RXsHPoFczNE49C1qbMykmpo0qr97NxaJWOcF8a9XDW
7LjgoKMxT47Do6NXwbfLIIW/J4n91HSi3mIAjEOefJkeODcMj7cg9QAZsZOH
my9aMUqKSf21NWfz7Z1xGshj9UAWrfV1chJb6k+Wz+5eDOeSpODm5uEsn0LP
3iDP9YCqaaGKwzhEQWgm1Ba7xHMovhh9vXLr2G1ds3LoTChAfmGrjY/EmwXK
mmQOr0N5756eeREMb+EArgDAh/obeMjw3uhM63Yh2wwLL0U83kOR2S8U3LO2
1J48LDAs3bxAro2x7wMEDWPJrVprehcXrFny2Vwpu+6pUw/HEdmic4yvavCO
7l1oulS7KY3w20JClbJ87D0fOjhb2egbSnOGKYakLyAwE1+D7XvXXoFOS9dP
H9/6pZPJ6mb4yDS6SsDZJXEk/YcnjSMUwWpaXp9p2Q8v6iKhgtgAfusKCdj+
nuQRqRn8udM3raf59SroO39E7P8+55kmHKr6NSlCuzK5P6kqFqqd7dzVp5kE
gnAGYnLYfp9S7pATDrU+kGqZKmdFgyHg2qWaxNn6vVFNX5x/5S8OGklIvbrg
DsXN6PdN829djXFmS3B6UC4Dm9BRpxbmyb3ztYMNw8cl3oJBlVh+mR9jdMCa
rvrYJn7axWa/Z16iIN3ma6IPrpzi5Zse7DHVJqhrK3eq7g/q+T5OEzcB2mFO
9hsyu0IlStvDVJWryOzKervvgiZnBJJQZOUEU5Qcyo8xNxAS/gd8UlN02NDt
G4J/tszikCL6YbcYD1KSEjpDkxvfS6pTLPCjnZ2yN8y3CqDf3SrJrpgqTO11
lEguuN9PgzhmsV0xRzVc8Tdnyh22DT8HFMXUFxjdtoIaYSXhH51XpVLiLI3Z
jpx1JPNiGC39EJzrnqIoWk52lc0s+VFA6nC6sDcngJstqkc8bSfNS5yjfm1r
jhMJH8e5sATVS21RlXmqB9CK4rOs2bEgFtGk0UuLgaybxmJsGY1MX+qkvzzN
jroO7pi477YsdnLeELXtwLuKY0IUy7pFJIsGUlv53vbL/NsrFurt6JgPe/QC
BFCeWBPVsZIsyy393e3rGhdCY+sIpEIExEyqWkctQNSo1J3DrIz21UR5izog
QXjw+GFN+oKo+eQa+PoA2dM3fYSPXiDFmyFkNfuUy2XuAzViYA5uCp9OpuQ6
TsAOZcmG4KZcjlLKLgn/zXn5tEx4gdpVNUdGf7q9/EFMpk2FvxN/W3SmY+gd
Kq9iSWL5vYRB6VRoR9/UZ6NAUCEv6cHF9Gnu9rdjgCCmhpJQGyt8vi55j57x
fA7UXR976HJf9iIE+apsSsqWDcwI9/S8GeIMjGGOfvoUlUAanQCa6urbZdeH
C/3tqIbd/HBenML/MaMgt1hsu1oslYm8/PoMV7VqhCYWG84efLchOZMPnOyq
9SC8N7eQ5loROhuJIwyzw4UdByAfCv/ANIbzEnB67qmjXo+aAsx2A3NIsq17
4TaUzkGROw8/tk4+YcCBbJSJYXfywR1Zq9QqK3DtSYjy12+t/B6dagdma5BI
3VhcFS6sYQHBQRtbjlRH7I/tBTVTYGv35gYZnxb5UN+n2fW/5o30kGgKj40e
yrcCP21rFyMz0YcJnrdwRzwsUxUmMZ9NAO/7Zos2BhDlxI+Wo+d0+iJfyFBC
R6hENxZ9xIyMnQoJ6Uyxkr9aIKP2rH8q+82ANx+UyRQ5Kxz8Bx6vjfZqc2Nr
9dufYY90cUotI0yeHxJ0NPcbdYYBkcGdwKRxEjeHnuFha/n1K6WuN9+uZMdu
MQ2ftSqkeriShsQLKQvljC/O2IsoqW6R6X+JrSMOjYhowGaExkWsQ3nxIbKU
TLbAfXxnvs3URAWdsK8QN8Obvz6p607KdRaG9iFX3u0OK64s79s563Ju7apO
P1vaiQjFKbRZO2kVqQykyphChczY9DaXEp2PKxY9v0HiRtQb2qXNnG5ROzRS
nauML/JKdN0F4tQqcHu3G44Cwqpfy7TGWLl6LOcpg7cedEf1GEDvBDW2j5o3
p6agvANgsokUcl/ewtGXjbWoElS8BTaT3wecP/E+2tWPzzeW1DuX6dFqNSmb
FYyIpebbD/bKLVA4Y6rvMQjo9otKaQw78SAEefpE3c6mHXsWtEshvYRasfmo
uA2F8WELXYTAOY9YebYpDXkc9smkIfKI7bhEWTMaKWZhZt64JStfH2BdPJac
Fv8Cam+Agr/jH01SrMuviv+VeUaItd5NxAv9ROI9xISp3iGxTd0X6Shkgc5j
XNHva+tz4xyUfjoVgHPr68uTykQmAJ/VUd8K/xqSN2V9zQmof1AfRaDqHh8x
t2ZLdcF1F/5krlZ+mBuoLglLPmGXx8HPX5zw+KX4YQHtFlREdld6l5+0fPue
ml/dfvyvThtu9avkr9j0lf9LPVx3751b+bGXEDBFD+ydsV++i5wOK08rhPOo
yd7kn5Pvxdd4xX5tvaNZHppB4GMH+8UhJWa933UcIE3GPAtmRnPeFwVGunpK
DWi/hA8TOHLkO/MPP9zJDHvLsMlTjNIZa4ARUJjXD5YTIEH/ScuFF+DGCY+o
hrBM9MXkjMBX8MxvTtOTt+t2oJ0BXqgzGfiz8/HaVk1ZIfQMJsgOaMnAQ48A
13kDIiCwmqT5+VoHuqeuOw8VhPnBeFxNbZ+7jSsdNFvENTWKZXYo3zOA18Nc
eBKR4uBAk4KBdXKbnqZKYNFTPOWSLKF5MlyiLY6RKEkNrOSWJGQzZP0/2X21
iejjMB20BdY/vcVs0zZuAorOgNw0rfNS6XcvBc0Xg7vjK78uKc7/tnazRqiC
a7b/PAMjyBWp2GF0cvBHirpvhglotLOvMONyP9+3ef9WLTn7S3N01oYzWD+M
4P3WcLg2PbUvXFY5SUOCZkkddeFQZtvo1wV0EprsB21eq/cSHXSS2Bds4gfG
MfvzsoSclINTBY44gVpe1kOewM151XNGznvDIJboboBN/INRDVYpNIiBpj3H
1kePevA2BEUmiUKpxXucbVHcD9jn5VYMP+z/h0PcNaYf/Zz48eAUmNVqPSeL
MRQR+HgC+Hh3GQ5c9vYY6aOtkBGGoNZjIBrO/3aRuPc3MH4Si5bJ93gy4w04
BJzZzYD85kXWPamdsD2i4zLTALSIMmWLdjDlHd7y3ogWeXzlqHrPXVd34/Wx
msSQcu46vBKsteULe4dT1xaQu12zqhpNSpzFPi2AlbA5QsZLPUzR9ISztVnN
lEuXMabvqgFpKluSNme816c9JiSJMljtVUQ2VkRZP3PrfF1+faM7RICNElxg
4Gpv8uv8ghV3SPwJYMepUHQ1PyOp064uQskOhmCcI6ywqMVWXId/efg2y75n
Tj/KrIzLX0+fveUXSNNXvymwEY3n0ZqD0vD+oQcLCtwESdt6vnNp+DZfLF8u
AiUs3FH4UwiRFI5U8cmu0dCSrLKd5uaSI16Wc/A1GGQurmNmth5sg9/dY1MI
+gGG9EF2PI+brfVPVjbazVn/v/ULZzMbfDxZNdNpXeCjcxocDhmC6XT+9hGC
AMJSx7yFVjQj3IVmQmGqiPVnzb8C3lsBdL5oDojMEq6rX6CdVeojvixC66rs
X4vijzFAGpCVhVxBlaBF2Ye4s04ZndeJXJL+EaqpdPZokhLHBkwAuQP6cVeP
8fBeAcEfyY5ewS1WDxo84OnKBTo8E6+P+4k6BDdA4tzVDEG9o5zUTIA1EqRH
IRn7zRsZilrLM9SjzqJm9KKXVWXrMELmVXk73bT9OU0j8Q9SDUtoRsebPKDz
xQm6MqmDYtrzDjPeYw6DThUWpUMPvqNY8ldMLp33l98kNIaV/7gmH0k4Uvwv
l2PjNf2lILUuzEpKirpWgprFE6kx96WE/PPCd/kzym3sJGhvQCn3eIY2ZwGt
l4EJdKZK7CC47wzrp6LJBDZEYyBTsPz5kQtVkqNhPaE+XebY/LCWieFNn2c9
6ADrACV96sxNBkB46xHiUi8B+8aW7XHvGjDB9ITKEyEw9Cwnod1ySTzWuH00
7qET2jkAdQ1GlDCW0VqsZF/E/3mRMt+aD2hxCYrAu56LRzKeo0Aw800d1/Y1
Gp6MdPB2IzaR/zepzyjm+6r1RG+O8WrYJP4AaVGkXRGWRxm5qi5TL4Pvqa4l
0TMQcWnFgTOJ+FjJiOgDJ3Ffdj1QOb+aX89jr6YjQgDbFvGHoB/xY25rSFuO
n5YmjdftgnvflFm57gg6jJYgbE0/iUctCiFbobkccOBev6YfZAHs/+iplI9W
BUOzbaEsIZrUA15wC57Q26IbeX3+ZHaortiKgKwGELgfDf7lCy0BsoiQbKyd
/iMW4lDy/omGS8N4H0Et8ZwcJXixo7q+wG4ziNLCnbqo24kiTEq+cxNFy7AY
493OOcFUu34NnlO9ZsNJBV8DX2wPhG5tYKK+qwlWPiUCOB+3JFP36e/BM/75
/mo74p4GCIFK3s60nHko7Xyw1OH+2ZSR3eN+O3Vz5coTc6/KIDDDAFKBmEJ+
UtzpK+1Hfe+dPd5xB2FhCW6vzVtWz2+eONaGzoqFovnhgfM8QxUvdJ2wuXF8
9J8xMewHfiPrxtneHX47Zucr0EyYV5VMWmBZ8vdcVH81D7WUx1e8ux/cvE7G
+woJkTpx20DU64DJv7JzizC1TdUMxKapaeD9sDTe06uslgyXq69E8ysB9noW
9Vydf9eoPakdTAR+KL7qSnAGrG7SMtD33QhTEG20tJVrPna0xUvWjVViTbP0
LANApkid1pPyuSshalYxHGuQjZT755vdTqBn4XCBeIoLr9rqjEYFDXgGGYGK
Zxo8iJE0747J40qOmZlJCh4Bjho5FvDOydmtN2e5S9DFRX9dGdFq4ahB56nD
d2Wcgabc1EKLjLZ3n8MpMMXlwWZQ0wEa1OM97PNaMkmdJqAjchGOtuIsZXDg
34JnNeCRMRqd6jjZIWyOX00Cqcc/eETxGi0iMsXByAEMBORX8c3KZ6QoEQQZ
BMFzT3SWgLgPP3jSQDKdegGHPgugHmJsNg97XbvuhUonXrUxo5CvIaSyIlrM
TfM2j/svOmTFmKtfwShXiDPAclRf2x5grfzqOmMTiStuqZxRhYQnJUjkEIy9
h1ky03XdgbW7kOiEGkRGnihHEy5lEUyqZFuX9nsOw4mXulhDN4f/mNaldDdn
jMZQiQ4UP25kyyiABOCjfGL9qo5FTYE7VNGyKEcEL41LIYcMxNtaIK5zCR3I
l3d40V6AQWVwJA+KbQGXtuhwV4S3CM9zuea+XheY4AzU7N/AJC17KIyrBbNH
ENx1qtyo+iioEMj2gqMK2oTFCfIhdKnFi2yFH6rAnm0c44yMsyklXnjhLC3U
6EO0JsJQDrRAp6lIChS/Yj2WQFnqFvvXe6oCNaLmVQvgxXkfHQQWL7MLi6VD
YQRk+Z0pVj57l27Uqbhg9W/DvEEbIABkwFvFOwFwhTBWZX5I0yh76ZQoILG4
Y1+Eqa9ZIVXHLR8JCdZ7obgGdegk9/PKW7srlbUav/GA4ucYsv5nyWP36vJN
lCqq+P1JMVeXzaKTGPHBVRmi2asbFYpix0ElEjlC6dY8Fe/pmkj2yU8uO+wT
9iUuTR5fQJMqxvuX0bju55pKNzN3jQ+h10Bo3UzqDS9iwKyFNgZytGHab7OM
oRR0pKkJoLmq2UnDwQYQgTD0d6bA1H2NAtlPnC5HgM2wK54BH8P2U7blBnE8
vgaOkLkaOsPjJfjTng+TvZszFgrxHNQSnkaOR+n8CjHALWexSC7XUksQWWsE
1mXW0NK23rtB+KPWvBZ4gd2XiDoy1ELdPOM3aSJhPG6MhYyfzKGKjgvrUp1y
sMuWumOQeXuGPdkfaMGTx9tvVnzMwuaGKdIQs/6iUoo+xKA0evIxIye7Qhb5
t2neS3zaCqpR/PXnuPcP8DA7HmqYBRRLVUlZgkCtZ1/UWPHKonuQjDFeag9Q
6FkYoNIydESX/9oS6l6rETyQTw6f2ruXhWLduqirvREHKHF36ZeeSZ+x0+kP
+/al4937ClL9zDWap66Ubn/qqprQ29V72Nlms7zc/ZuYrFDv/CUnvg7Lhihf
OPchxeG+hfVBcKxjQ7HIE//8OydXC2sJjagcpUaen65r3zMmHhElZtifJkky
xYNRa5IrG6eifHxn15j5m0yrEKx05FvGWoQtI7bMZGLHnKqWOHYP0HGB6Vb5
cIt2Yn+sRy9JI6IF4/aMHOLfgFg/UNmtV4zG+xi0za2o6XDZhCMIlxaJCioZ
8Xlecxc/8sC7E1lZ8Nk2Z7zpYkT9EOEjDiT0NSMhQADvQJr2IlGlUEpVXB6E
OZIEdjECtu4uYddkl8QDpuky3ikWVp+xicpXwHoFvV4xfVHxBOSoJlcFDgoZ
Hkf97q2LUXWHcM0LY4x+c4ZPDBj+lLUztXtUt+SyANWbhYJHQgxVoo4TN8Si
NFAMePcg/chC4poTisVSM3rCgZ0r7wjHAKflAuu1075mOpjp/vC5qSEWCvw/
ncd6kJEIfB/3TRBrGm6BGwSzE6caqwKb3dxqVmbCx+I313X1l2k5NbH7KR5+
SlwKv0AuZIevvk+5x1MniEY+QfXGo4IUCkgPYpsz3JIQvGIc7d9RNfzftNrC
2aXJM9BNY2BtwNBWjkxCRKZwsoCeNcsr4S2ue4iaN+hpz+aAKenfGi551Oca
7CfzGUptAMcR4057svOOCatg5SgHPJ05WhR5UHqKbFjaz5eJqYz9ZcLHFdex
QgvtBm8QceQuP7luxjzeCsC1GXmTbcvn3k9/ePrlL0I0uFk5zn0z2EgmYbZu
uijD0k9FsZBBwsqyWEvRi9NgKJSLzUpJtRv4oS+oNk65rx2d6pIjKYoBlnlz
AEzo5Hi35rJzQuH9g/m9FmkdcAVKD0nDb1MsirnMG+XB5iGC/+HCWDSh7WHz
GhAjHfnKV455bkqGSbTw7q3vSF9DAT0GBGc7LvO9z2uYevU35pE0UL5j7c+a
f7iX4Q4R2KCiC+5qttaIp/hoWEgSTI9IZoh18xSZQZ6doFMiFlvfuBKuNHlz
ZEum1rpRbI+4cf0jV4ptIA/a6QHGdeH5NSlxpP5oHkOS+63rUU2cz2EwXO/+
orE0pclXkfI7aKLU20WtRwFIcjVjQ9Z2GPcRElvciVGXrPN2Lm7lMXP4x4Ie
e0uak++UavyKCN96dap6GV7Wyz+fwjLSeCuR31W/7yXtaZ1ldVRT31DrpG3f
0cV4d8LaykqxmvSQXNCSCVnU/+RMB/YoyFrjN2mBzyCZV7yVadh28GUkKCCw
NA3/G+HZJMplzFhQwzr1ioSEJLO9DMYgHW4f3NEnMD4zbObxaf+rycSpW+Tx
ILIShUF9QhfHkytEGygtO/qJDu1+U1dRN0D/0hTrdphccuSIYyP5WrLTMZt0
za60LSJTaIBTLapIgIDEg295HbruFrzoq1/r5LN/aec27haa3Q4s2wbiwssN
409RLWXjUUXybp3HcvyVTFsVPPghVgS5tju+/FOA5tabaoK1MkOI2XF40Kc4
L8/ncYq9tdFTdLHZhuAhr/ymqB1dWPvUoWwj2GRIrPIqtqb6nkwC5MjOf7Vg
RoCSDG5a3g7rBw7zEaZjstnFqnt7rugXwj2J+SSZ43KeMheTZhlELUrk/+Pk
m4Vd19hG/T0BLZr0r/bh54pGq+DX6tusQaj9yGlb33hctaBYXACoBmjUCRDr
CbhHTOVMIHt0F+EJ+Jl4fkraBndS6WaOwAh9Mf3xgvgvkJKPcr7jru+OGe1Z
FWtrtlt8dB4fKbNz1hn4OsS6V2kHFQvVhTt902QE9CpFT9WAE6GXaergk9bo
5rRaCFMrFilCwCWsJGBDSE1+laAFuxim8jFDg5HZ7mAhXdPY65CK159XrK1D
zEo9hN304KlC6Vs9vfJ5iRX+bTDgMlqP57P/VCJ/54hjwejBnQzRwl9fPM2L
CJR61vG0kFuSQIJG4Q+VXCTwjNOT3X2L2kyK2u7kNI/adO+liRQjK2B4Q5gY
x5LABkM8k4H1sG5kVrlD+ems5ipKEIv+sow3S5GjiRn1CrcbHdHuJ5kzCU4s
Ph/uIFWCIu8foa9KSSvbx75LySKk8398sXVS0PZglI/0vorFERdU46CI3qkk
pz5ljDxpKO7ys1vpsGsYKjq4ko8TxBt43gaVzxDqndjQYoDGuQjpyYJSOAUr
NxvC5gVpcObbjZo9yuvfmnjJlC0ny3VCvZUOn7fZTSAaYbp+VZ9zusKGq10Y
KAY9cu4Bc7vRLQebm4V/jxI9CGFbZS+cEDhqw3b+AHKDNGpGlDqdC728btl8
n/s6Hpscuu3iqWmBgGQszWJdS++fyTvCupzVK8h9CFliRdvhUerQCuce6aCb
RfY8oWTmqBmrVWWQ6SvT4sg50anr8OSDwYSF3LxuDwVLMGBsZltToAoIjXm3
b4+zGU0Z8UxKpy79uePaZZdAw/Qm+T5Egz2h8erlqvbrUOErv/ub2dVvZoe7
ftwyrjI0bduCakGkKVRH0otCKlL8Qd6Idn/+H24M5v0Zs4T9D3usc1IkX/BA
VO0heRAukJbye+sqoY5JEgEnwGzfc8qG3K8/DOBAtUzVGHIp9RCEVHFxHhbt
GWRO9fxrK8X6csGXGXYvUwz1/L4pntIT59BS6OgQA/t42FJkadumcuLHTDUo
fyNrELDo00UD2vFNIxnCsP+4zo6nCDz47TgpibOeR6Hk60gR9oGvY4uCil4K
6CU9ut0eQC4yDBEDKLRFS5xwxoccYMYZQ5X7V/pZXAaCqEZkt/UJ49wuOYUN
eNSztGc3PrRvnTW5F/v1ZmMEUtFyLC2beleeridmEiKRZQxtLeXf1LBN9hsy
G4crxxKPkeKZhTgqMxBGWmVSIlLumsC3qhWmEQUvty2VuaUQIgnVAKebwmmY
Xxv+mNZC4oHfVpdahJBFkkwAd+oJQUzKBGxS5AcWyZx7mOoaID8W55Zxwx4E
i4wMaJ3x5OyYbqwlMpasol3EEsVWMUFaUgNombLnLtffE8lCK9vrioEuIikI
M6qNCnac1WF+Zf931f4Xl2QhL4E4PxTaombaQOR2iBEI46f254FNE/sPZe0U
yrZwXtrIlSvMQcYFpilVoJIKD+CW7NnQqooLIduN00ftba9sTqfcxSpFmzQA
fa6kayWzUVNK2ey0vfaJzn3i49vO4VWclInKhWmjR8W3lc5Dur9b5kvnl1uY
geH+ReJRijqKXfc2jSZWx5LCrRSD1crIBNCWKlfBV2wsdRoKemJmMNf7MiMI
XbpnjguNp3dai4PK/z/27QUDERrPdLe+kuLmP3NTjgWsadgybJjyfErbw1q4
66JoCGLd2otIuKBaxybZ6arvJdvL88Q0dtoy5XqCik9CSYsMEDqXM6DbLvh7
nrLuTUTnDnzkVj/A/IPQSZabZ1IHArXtzdIiM2CO0xTDfWzF8GVPjD1NCkWG
axQ6mZQMo1vbV77hKqGDxIJy6KqaNzV3mCjjoLRzFF3kYsZuocPkPKOxRJKm
LqCr8sSrBPTEehfqrAOkYDp66OGCvHqgluGi2/lZslo0hXHqwELhOrE066cx
h+YVXo8qGMmADPyp+wwBe5xI13lrgXrCyJtDs+JGL0xgQsGFZ9O6avAjgmQA
nd85yJkYn633K1wOliC668XDLuZA17WkRZwwcOSh/APnWJFoNjbEQRqUYaUk
bTLAdZZL5xEK2d0eqdYThNlFN+WSJJ09CxO1ssGDve+/T5PKobpyfApjyjUl
zg6xSp9TR0hD1byZ5vQnwv4zFzWOCI+ci3VpRwEFgxOvk6BtnwEDpQKTrth4
HXsBe/jplvKywFdZmNNzgmPcBHoM50SStnHMGxVQzA7EygWQVNnP3vU1W5qt
fWJn2yW852i0+NuffRk9QnetqqThtI2Y9jKxA/PD55AQUQJ1XEvtZl6qjgd0
XbPbcxFkqWlG1fP4aP4MfpACLXYt0x/mqHQ/3S06yTibc+ek28NWOUQiGo/R
96ce3xtH9lXZI+ztoT9MP+JVsu45at1ZwX7whq8F9DBdkYmBiP+OFW9vxtNg
6GS19Yy+ex6rwCZbzzDDI7uT5koOqy3d6KF8y8awQYGppzkpz/2JQMnRnMoc
0qH5Jqnk7bHUGaOvsKW72zQ7PH97jfV8JAKHERbAcPr8J9YtxJ6yU6T3QsAo
/Ey5t4mJKo2HmBFqwT4DNK+7Bf8zlf3r+QCFl4uqBbpu0Dx0u+sg9CLS3yle
M4RIR0GybVw3XL3qS9UdD0RNGCD+aY/Keco8bAT45i8r1VticxOFhieGfVHh
y7Ngb+HUNyuO65dOMjud5J20/rwJ8bl/ZQOHh/nomfRscYx622XO4KJQJhny
SpG0ovzSSAcS9ota1qvreH3jRJxuP7xAFpcTfheLV/tD0D/IJtwr1m5T4M1U
nJBLtvg4UnXZpsFHz4W536TQo2sVQkJ4jNxqg0JegRoOHAMZ9MvR7RKjNh5i
HSg+c+bbSmIYFQ9Yq3XJzWER+IN8V/tKvzXdz3xLdy4xMjfcvbK8jzwlEAwF
E89llr804rOGx1di/IL/yORvEyiAu6PN+NmoAgtHmClSWKUlCzvc+61lidia
0c+fwOQjxPnNl38oBwf8v1qgnVXC7RZ914QC78IPGhV99ZkpRWJ4cK9EiuH/
OeUP01sIaEgLb1oOX58StqmqkypDTyIqMJDbwRWm5Ip/w6UbJ4b6fG8vfsmB
br9gcP6iQ0XdbLyrTRULJsOAN5YxiklRp4p17maCld5xR0fwHea/I3iW4xfE
SrD+CGndGoaIoPwCPqOYHPe8n/Waz24Wd+K5Ng7bhBHHhpyYxspAp51l5b1c
w1yO+l6Utd5v2t8wMxjUJ8zZBGKXplsURVHZrKAb2ixjSk7qDQxcu8WzEPTh
ivhy01BPgMhnHfUCpkXEIijgqgDLKXkcDUg2Fp+wbIqEsWM6WQ3www0PYsmD
+uMIvh3H9TlpfhdHVtcEAE+9gl6BhpdSQ6nLlrjkXb02xc+8SsaWGi0D9imr
PHXag4g1v53uRx3gXvkehkEQX+WMmlHjuB6ZLwyuaWY0BI3/DwjOkrLuVWKH
oXU9S4kylCIDRKGDRTk0XykR2/8tg0dEU6cTbk/2DFG0rDJle1jfAugbAyr1
jAJD1vzlVeHj8TlHazRFtc88jM1xkcX3mFaA9lnw1+GJit3P+neEFg3dm6xd
/z3m0DnTiavImekJyTkRhrMH6OgDerEBLH5upTGFYetvxzbM0kJxWJ1+KRxo
vUfJR8pSsLHf6vMN9gqWv6IheGkhHK0oE6+PWtR4RvpMcd7x8hl24dB3nR9K
sLUMzTlF+erEJBSv9h8hMq2aHZyewpwic3dsR701uLtkj4tWPFpHNipDLvNX
PeaS6FmJbK/7e7G+Z2fbZgY2X7U7HrZyiqjjFx5bMzBuV12kVLRzLoNGvyCE
k/oYpAuhLKbp+IHvFTQ/sPbTtOjEWWKo+oJIP2W21/81uXOHGYnY/eGRwvle
ZlTP+ywWff2rdePpEe2qM1B1OcyRnd6YhBA2XF+/ByJY5czYyBSiIoX6gXAY
ONZVb2RC7f8SGuRkALi8Y2h+FMiAVfGViQKHNsVIzmTAZ0hA6s5HHlx5Ha4p
2PfHGWHBij7g1wLD1yyxbF6uHZGRm29JWdc1jXshsjnOgwuEDhtQsi5HzN4o
NpSo5bta9u/w6LSB51MGG8yaxkvF7WMGZcipQ1eOysftqD/ek8+7uDZfpht8
/SAF23IpNSowQPgizEZA25bkSE7YYIySnFixxhtx+LGCbq961f6FPAepa2NT
lPkRXrZHX71Hgb2lGq4sNF6pWQneaOCOwNEhJf/8gD1EzCpAHUppotpb7wRY
SUxDNpmzOO1mzvGBnRR/oIJ3NHQMQJXI7kIollyIXtfp+qvAgAFCJ74W1TQ8
+0pLnwE0lNP6+IsZt7SInI22JIRPMlaO8lzE09liTeOjWic9YXdyTZdbBKxc
1ZjTNSh//x+Y5fFLWiTDBKvucEcfL9bmJCPtCwbuP5ZfC2ccfx5nriYtE2QB
630d78mTBwCc9k7fzuJhPesfny+A8QZpJEoabDA9q5LLRUx5QSSOblXWFOI1
4QEWN4QZEbnm85QeTyg7qZLieOq2I81uHR3rWyPwy6EabyXCzNVHLLNN8CQp
XJoKBlZgX00tJbfDtT+n6cni0QB05SuEwVQcoZixr9OZ1pGXkcvoepnXdski
epKB5YcuU5/2FhcN8xh1GAOhkQkvw/iTQk23/qjzBcOu2rD/VujR+JaspW7A
s+et98g4yYuV20qLlxFQYtRPgfKXfLrTKz3xidminxrDdp19GVR6DBiUoBnw
Ay2Mg+mVvpBlO67p3s7nPtT0pCEu2IEx1cJOSi5v8kgnD7gmWu1jtvhHoWRo
XePasgdpyu7aRHhtw82UbeLDFfaLNZZ5Lar9DWmxbpljwVoa7/bjgxA311Wi
MAcdw6ysXY1p0Yqu9bih5fib98LCCHpzAPR2WA3oSuAcoBf01ISPiW8DaedZ
2YKqVxvES42/lX+HKNkDptIbI4iUZIWaNNA/puxM062cSE4MOJieSLN77Qha
bSpk3tzPVFiEQe1oBYtgs2Z66x4HOxhz+orlTbu9/YAlk9BbhuwdKe7xenTV
CN0zg32a7bKMvxFqsGVi7P8qynie6eUTsi+IHH6Ma28xd7+5FhHnNPQ2sG3b
u6CdifEzlenjfij33DNJN5pUMcKw8If/J8wn+yGCtkPGbU9FfOtxagqoUY04
6eMFChIfmUYFY/GKntvVWN2stgUwbawGcsoNIDRURGBtvaKV0nvHi49C9VAV
FoNCNhNkxbdU2HQcM5DxvRkPwVhrBzzQZAj+I8E9rFk0KyZrEQYntXuDBD/A
JJMjF1AoIcI/0SgG0rSKYb3itCluHA2PnOKn2/bYXd3HW/XCmNvjEoY9Gx02
S7KxdTamWzOcnm0H/s8ziDbDJzBCIkbtrVsPe6r15ezQ8keMU9VQ0p2MBL8i
bAoasJaMDK2GDpJUCTeDJgqpxBEcysgaTKkfNyIKPaWnKtV2lG11kvSElWAA
mSJIlaE/zkiFvBjBDwwE9rhVtg3BS1IKgyYrXq7IEVQgMWaTxf/5CP5yFZyh
te9mnFXe6OoTanhgKp/DGU3DaclBbPdmgNwbeE4zS/0UptK0x7VKJTiIxLaZ
ZKeCWkAJcWwp6UwHvXke+SqEVw/gRKN8PLE3mQ3UGLUT1OxiyV8gDvxxo0an
AF5YgJVqrFfXOS5Rk+UTnhzieLfgqjkJ5gmYW/GEwqQsy71V+vRM2dyj66WJ
pLzh2vdYItTcdKnUI5qNNoxizGj+wAUdliFLw1hKOfhy2vM1kbdlJ8IfzWS7
YY4GuucwmObKi3wW/aSVaDfuDc4Cdq3WbOSDe1EUwM8vf5R8TWze0fjrAoMN
UbVnIEfrFxJqIY11HmkDiaT9x3zlXzbKeW+IPk4TM6PO1OmLy3wdM+P/Sj9C
T9x4glXRpQi1/SiSmAWniA4+BMvm6v1sdX+t8bBxFXPXvZ+C3u0qtdC/3dGj
ZpvlhNo+1oVxRSXmw86PG4oF6OxzSBH9jDupG8RGagygUTc3B84wqcMvLdm9
hzfFghTPGNmAXRFnpe6i+oCFTyymxmAkkp7TlIKIgDki2AnctZ/RXI/I+Sv5
FC8gI5mIBPaQSBl+OxYbvRWrbGz2pOBFQqK/OKaN4amkVNMXmz90t4UE2w+P
L4ibAGJcJRkuQFdZ+Xm7ZgGlrDef75TOgn8cF+dsbL9aRC5fHA97Y3Ry/Awm
phiHjrZHuriMrB5ajrqm+mr+AUgTF4wBbDwYOtJ3Nmi0JoD6aqjCXq/6jUrm
GnzMYiQH4Qqvren63kryuHI3KS7De1Sj5msM8nyXkBgwxtNiN0lZuXYeeSy0
Xj5NwxDNqVHN0flRzpSGW+LABocTr/gP3HAuoPk5B8zj6yb6viUTkkauyCnr
wKlsqojNuSa77aMmbWWTRxh2ou2TSOXNe4oyDRMjBD2kvREd1DGx1LBDvy5H
/G3dkTwcCX8/PREqYveZ5lgJtz/DYoR/fcy2JICGQaWKvnKrn51P2FZ2d2Te
B5L7CVsDOB0FspU/cm0GtcoSQqFjc2NciZdde7YPE5tT7336N8tDjxonnmD6
LLttEIIC4ytMumLakzIZxFC6EGzWDt7OIaYO6vYwmKFJxl31LpSWA7YxB4b4
DrUlCeNFH73XIIklgbp3OXpMCYgT14/aGL9wwX/VXzbASztI2OlVYKh1p5YF
iAL/yaIv/y1gbnGtIkr5cXxG3GloL1YRDv5EBO0My1db8vF3LqBxnC+o9gYS
ckxE2mWR+/MNLG1cA4aOU+50Zctiap4A9+ilCNIrDQxGhJZYdvIvkouRCoPS
CF8LWXsLtC1mU+qSuGmank6yhnhSM/OwH6Fq4me4ilQ5R575LA5CGHvlcs+q
eS95WnT1loUepB8Ju7H3lyddAYjyyWadiUSc65/PJIvWoAMj3rpaQyR164SJ
zc4k5gjoqxuMGiNT4kbF4ecixuUtmlokhx+N+/1/Oobe1FvlVqu+8xwhQ/oa
BI1QKK9hJ+sty0u9BfDAWFqSwv8kMde8j8lslXfAA8a6uaOXXBTolAeXgLay
02ieui17u71/qu2WbX2QzPiVckNe5HzG2kSox3pywxDiCP3QNId+atMwAC/O
cxBgeNeP1ZlHvGBdcKmG/rpHMPiK7OnG2TCbiyIgQMH//lBCZ3Rb1MaKExfV
tXVQKkcNw9pPaFUFUcADl+RDxs0zVp1s8Sy8x1q9a+fWHJ8+gv09mzoN8Jt+
tHM9jkjwFJ3e6L2eeRklreGo7NIK3YXrU3iuo33ty7vFivv3/svtgFSRd0ZQ
nxQjA7LqHEcMBtrtbWxcdG72+5yvnRxqw56W6fB9QlFTB2DqOHUt/jfM/mVr
QfKDJ62/kGmdouB+bDrH/p5BNVAUUouh/s6LiqXyw1ma7ENfl14o07rShe+q
sN+54evkPeXygsKrfzU3f+R9CbPAlniVyJpyq1wQQx9tqvowkyopd6uwakxM
7G1CZvrZi2OuhmSWQqJVfo7vof10nDEzjM+WTEmoNCQtJT8FcMLP1aTvR3vK
devk8pxfjmoByNuN1Qon57CHHADyruRJZENMK4Y0lU7L1nglm8vP8jx8mqhM
jLsGmx+AMMeRGb9hq/Kp6jGHpDIoBZr5TPWuaLNirKbaHdNVe/IemaER3u1a
Ldj5/r7ZcRYSGX09Q/IihTgJ+oNp3A5fVmcyzD68xxliRPV6dNRb4LZcf6GW
K1C21bx7Zak2w2QadnUsylka7JtiFwDaUB96znNNvxYQhcskaJQ1sbq7wLOm
D2Xit44bEAVxxTiWBOWg1NYLvaSdsYvRJwWf4N4FPS01lCCvtxIup6J5naCy
0YRbwbMJj0CIMO7/o2Wv5uEZE5/fETk7Ss02SFCLRy0AZvBtfQlC17wn/UrM
z6m4pLJiP9Mz30QGsDXqYVpfcLg0e0VQ8A9DzAPupvrSld3PLixp+NNYGXnF
XJ0wOpbEYOqTW37BgtFWNjASiH7xGMYYIkbXMIOCkh/zBuVSH1mSR2J2ARwj
Z4K4gy4c/3Q7zjSih3HUkwGXKo4KKsKNucUchd2Pck8rbu802G4c3KIcaMgo
mLA/Z0q6vwZWvvtj2khDUbtV4ydVhMdOwsmedjuG847sZ/++Y5RLgyESaNY9
u8z/LIi/rGBWSEZgODHRX56KReGTtyelFZ4sjCfLR6+K5BiXvVTy1Ca++0mq
wHIf8mIaVpTtnQNUOBYlBohe26PymYCaQgDjCKdxx6pKRAvyoZmdXjO0aTMS
Qt1tyNMDpghXwl9f1/L6M8wXGSK2osWX9Hhj3Wukj6VicIRtgFaJ9PK0KvRZ
0lpDSaKW3VJuNqAxKzOZP4/ivkSsqDFH+wmSQeMAC5duA4dLL8An01GGeXsd
mAoVexvxPk8PV0DC423lK8HjSBfDdVRe9Biahb2DNXUTVMsYTH1rtrpqQCUr
2ZyGsbDWV3F22olG4gp8ypNF7qKq/VrHTb9RJhZ4rU6kZzLfeTkj0Nd3ufYK
0VVbpCBUDwcB4rqLke2MBa0oQy9hSlAORJNZRiGq07mBM+crpuu3SjdQm1mu
nQ9n6UK/hIyaDG/gOysvrgfHHFLn9P1rqpZHANAk1I4bNSLYc1MrFnQorMHi
cb45Ycb0Clzmt1itZsXBNhOFzHWt7mBdcljlYaUq+s6MiQsA8DmrF3A107mz
4lgcz/J+LCZzY1W1SP+6s03QuHE9UcN+zrCXuuPMIQJssj3g8zWmTe7Ph9ja
DRdj+/bOlAi1Y5XAVDAa/CcVzlfRylqR7VbD47wyorWDpXVuHusb6ZfxzEyZ
Fm0/KbvoxBNpTSp+TpbySnBMpSHP2WUIIBKuFZetDThTxxo1ynONmSbpF+Mh
7QNe80Yq6fihvwwJrlYvwpzJG+DxdsGKlO2c0gYQrEueqpvGvhwULX8xQXYH
vJ+tFj3ikumtfUHjmpvL672vS3LLGy7f7nqUZXzFtZ3qUoKKU3q5tArG4eTC
DhP5Bm48NngxH1A11blU7kW4eUa4xgxyL7uMip+wo51Sw1ofstMZV6JoEZ6w
62OzIXoooZnEfbWlgBeoi+q3hzWgoAGFi1XdOQm5A/tEpSADsFMsaFwj/dV9
RRAa4AXTTiMs11E2ANsNz43JviCPXg4G/W6R6BDrXJDkYZQ0xm6a410H5Zj+
AucLF+n0UF26JjrEUC/ASTrDwonCaUsu/3TXTWM3ReT324PBcau4nm8xtUoA
sPvb2B5jAnD1FajV6kYNf0OHQEtP1dMk+tyPmh2solnY95cLF0e5jqUqKaUh
666akYs0WzFMyJFITNTOtWb+9Hsz2zNZdrwii9zzMcmNwBs6vEqQO4rYQPTT
64ndWpXjDyCD0+SIHMq4sxhdBM8cCWK+X1sTOKKX0SSZodTARIi0y+z6xvYo
XAtAgnzz0gA2vSdjA7ko2Mus8GdzN5lRhFacdkVLsXmi07GxM8ZS7W1KIwHP
V8ZU4oRDKuPpB8nGQMzC8gQpZ1132/IKvUtZS3ormrNRso5hyF3mH/poJRn3
YDlz2tPyrQQdHj9zOwaWzTqflNVAXdQDpOnWRLDR3TtIALTCNsEcnZTEYZIQ
D+A9DFDAlLKVCoX1xBJP4oERmuDPJLE7XzkUHjy4hSdAvaon9BCSNUNl/R32
OotFi8XWkKoJEqcLeS1gcS5wYnbBoaKu68+b/iYeSbZsdFaPd2Wa+6tIpCpm
JI5XQjWK1TWLTZO23KH2GBzDiOF29qcNTQrBfFt/YZ7X/YSBOHRcEykmx9T0
8QQyqxEQxVzlWNj8/oPlfoMCRKtZ9KV7rbN/JBNuLSncPCsegtJmv9SCC7ch
IyhQplP21SDHStg5oyQzVahUw8nOFT2nCvooV6abioQSPsSSVbHGMzpgLZwI
tebqTf17uFZvPrfL3lSl4gvNAXI+HfS+575Rn4rZA2D9Z7rMqc/GhWJPZZSi
Ra3yv1l3TKctHCyH6Qjy1Ks8VDNB65Cuxdlq7tQyGMwPILSzwAbiYp7N2VEi
BEGMZX+4FlaRYh7dmX8oTc7pHlr7rB50ymKyCa4UENjo9D1m/1K4uqo7n1/s
n2mYBgk8GSEuPwXDmgvaEZum4XLiveiyafsbtN0qBc0ZQ8GKk/hIu74rPNnd
ViuW/F879eN2O9AEi/dAJze8icTxbXSUBvSFL0rYam6Z98BEaRGCHilNNaDC
zcN3vdbhwB7pikIkAaPbXWrmegDNsvL94vqL2WyXv1gancI9XJAAWG79hAUC
Ajg6UyurDI+S04PIMrabJcG/tZpuGmxTaEBAwTzsW8Frem+eSH+xyvGnfovd
Sa8vvqiqcHbTCWmPsUpkoor026jLbHLn3ZX+5UgNvwKNy4/5JdR+sMSjetbb
bbx6Hlrya0qPKCFfI/hCzkfOC4HmKiFqQsq+vROgocE0GKzwNh1FCOyRleOW
AqTSVx5cXur8OdCOMig8PE4cLK8Lv03bOQuSrnvyMtn8TQFDpR9oJ7If1VYh
kEa3J8Bf7HuataydEdm8PlOWKWFmJkx4Hf7dT5JH0/4rIaX8TyylbB2OXCh+
tYDDBuTcZQQspMI0BYOClxsfRUuWh27fWAt9v48CDlTnyp5DE1MYQO4xOYOJ
la3x4yJGKXq0tU4m8mMFdu24c3IU294xm8GMAu5TMcATsi0fsbgYzxc24ut/
fJ93Dj16KowhG74gpgmdD/fpwi7k9AOMctm9gZ5oTdG92hiZeO81zmeSeXxr
jqfFYCcTMSYaIKvV5emX9Y1TarfHEbgAW9hMl2VvziawhOI/sGNpcfFJhMQ6
DVxgxV+S40gxvUHIdxOAIqgl2WTJfBQTnd/WMxdm/xqr0A8x0M54l6bYW2//
3KU1vkb23Qaov/36FiwHtIGBWGwY/uUYVSouTeAp5lOFEHyt2iL0b2korOQP
AJkIGcbZhnB//mkBxiLyhZ66K/goCT47ycTAIFI4u+n1G9i9NTC2VOboUays
PZ1jbga+GIx1kaC+t7s3G9gyGG+AigdfYyuZtHleyu4E89syivGmYBP1a+D9
4KdxnAYNyDuh85mCO/nvA4+EhM999mpEBzOzRUANjS10mBSFno/2NAwJy33N
++FekKuTVD+hQqjKFyuwF8QgggEmgfeVnnR4/+hW97okMhjTHtHSsUdNrVKK
Gjb0vHaCZ1NQxpUmJspOpH6cYc8CeKqgND5XLxU38UAuOXsglHe5AI1Xzf0M
hCOqUdgEno/ipirkKo9l0VJWbg2ATWhXoNO0PpuZ4KNApvxhlbSzQdlzIBVO
MiYje2lXw1hB9jE44PeQoGwjXVQ5RYSnp/5S7e0kIYWdWf5LQllFM6soqQo8
83E25Ma4iZ/jiXHuTw25PKNVChjdZvDGFYIydz2qMCcuxSG1H2zI+I2QL6du
0BeIsMUrHpFJIIZ4eae9eoA/WEEd3uGug6+CyvpYMctmwQIJRMau/9Owi7iP
hNfi9YiFpRd9bUVcet54YLgFJidKVhkC4t+1Mw3zaLwb8EtT7Sw6EbLVNFJT
1rsd8lkteHUTVbDGKeOW973KbcltqpkOm9C1ezMfijTudHmYBFz+qLJkrP0g
jJdM7s838+Ye6+6Rz315JrMu/Qhn5Ti0Q5GTFTxCzfPFmrZH94dysouMxMni
78GOP0kVjA/XH6ZbwJq2XmehL0zpMOzUR2WDlkgw2uwpc/7FekllWw4T+HQW
aSyWlogCeWLFW8S4hFlBokXpLaCadJ02JD66OnL6ncHQ2/aZvAvr21nPJk+d
FiZQaVuphRtsYWZg7N/UHZDGWiol98sX+Gx4zZo12MkMraVDOhCxIpFnUV7Q
0QyWEvpsEzkKXtsyWQDimZZydfVhQincnLEpAQW92LqvJx5MUNAWPFV96Qjb
7ZqqpEnD0j50UJWpa2tagdJnjvSpdVN/2PnqLkaVVgJr1YrbtBTHKPWOo5FU
jDeJCaWUhq1HR8Ro0tTB0zDA0OcxlTXi3HJrko3DyWCWWMLvICbLecRAcn8Z
kV4JVy863YHRQUkFlNA8qdHYfcNG+emeklKo/Kyuft/gkSeED23hwZuu0i4C
KE932nNCZYiHNJttX5QNnN9TNIhutO9a3+MUsh36CDWpjq3Z1ZCY4kDEYEp2
EGi/iONa9cw4Hi9K4Lbpjcqj8+gKUKJ7CBbPHprOWzcCqFXhKenD0C7gG+fj
hheSMqUavwDG8Lr3TFXv952K8iW/Pkn2ZlSkGpqaWYvu5FunbnxhEOWiIY8L
Sc5G5Da3p7e43Z+dCgWqj9pWAJJS6m5yiQQ7SUfdI3Hq1JARomYslApaR0rQ
nNG/0h42hpI50y8IjCLT0nPIy4hMvvn3wfRj9V7U2pOET2NppZ61XPCPFRlJ
eXL3ch3EqxlsVBNmryWCm4o+dww9MwJg2KmQtU3cVfykBDlqMcS1FOoioWNd
hu83ghVyrRCejpfe1Nnz142gjNMs3jJa5gngP6noY2ExwC5y4p3+c0FPk15X
+p1QOxpsCbAj//s4s5z+Ud9LcpSMw+v+8gnOMaRAEiCyO2VwPFRMiI+COM8z
C4ISPnjOyvAZVqiqEU5m3GDtw1ai9uVAoZ2Ayy8vMefS0xU6HXft88oysUo4
uG+/dTiHENNygFer1K5u7JerYXvNVfBxQSwv0BIz4Ksw7dPfd2qwoNWL4h3S
SjQF9Fm6JWzAfHu/Ui5Ejsl4ZCwl4qDLwfB9iEAqxM+MituFgJQalE0R35Ia
U37DzFlUZQqZ8li/CSUO24rZ58Vcc2kEW1WoJ6UneIHj9A+nb0aloYR2o5Xl
S8rDiuEaFmCeYvSrMe19wU0gsKStvaScEsHF1fVlbLtuLv8bUZ6GlLItsTnU
jKSYRVg1K5lwqdPhtPsinGMA5z/4AofG6Izg8DF1NeDbyGYv/fymFoMvIHLu
rb0YlX58AgKugzWs8/Ozt/AQxGauwPQyJSAkGTkYEs6NCkJgVk6JtT4hkMSf
IzNy6ueOeoZIi94o2LFPmppAuhXZzC50joiqsHB2YLyCV4NXE3dpR+hvYIDM
zIqNDWlb9A/KwkOv9x648IK3j/Tl1f0p4ElN0GevSCZcBseo3DHx9wxyPB95
C1go+87fOZFMAXXPjUV1MLjX28TqkbLtEVn360WMu0DEmQVePgwPQwEbYzJB
1EtV1Xu/uib1BDJxU2Pw2qrFMzH7LsCR7in5MZgBBd6ahTdOorihxS30k68R
SPJAzkxge/z2XtbKMwXZCDYX24X4zBMnwAU0UPrJWdaoabX2o/GTQT2TQbol
7y1HjDs6WxJSVn/PPG/jvzbQXT4sasZ6DVQbWPvTlX8EcjqfGpTu8RtCBKsO
REarMJ42RX6pjQv2EFMmwxsL5y9UTMA3lvPYtZpgr/diR2ovHZ96OeCMkMlB
PW7eMgrwrEnf08a7T9YnCr09XdX8tMdjubg8NdGkW9i8Bl6sXYawZyHIEIhh
r4dOoOoYFk6zxW9Ptbi62mdbVF8WNHpuf1C++jYwx52xcc3OfZQKYWzDlFzs
orIrfz3oMNZB2BYnMI1ZUM/m/xRUPn4/uALRb+Tmbm6m/4HiJbUUIoN81EO0
SuZRfyhwl6bMuMiQLWAbEl9ZD83KsMJvbHQhOr/KG1XCPHqHv/8G6dA+5UwD
jpd/koN9IY93gVbdeERxc6BrpYXHjsNyiZvgCOXMdijWpZsSx4HRT1dFvkGq
cFU0lsrDcQMM0OOfA72+n+dTUPaNiUJzC8BP9s6bhUeEZLGSbNrqBfS4yOZz
DRmhwrV3thODzlSr1GKa8/k1MCctdjlSHnctvYACmYZ7xvv1PaSIzbJbsvYA
1uR7995x0pqHELXStLtCkR707OnQt78lSWB0empVJnuUPDbI7j02QHdXND63
6p+2qHsBLYEYu0C0pQcZrEKLIeI2xqU7LC/HyBo4m05rlhlerMFWOS7XkTb7
ujJBWW4wbOZsUxaTPiwRAUIYV9hL4zzwVJwvt+0yDj4zHttaGzxsE/uK2Rgl
blT+IU34ZYeiOyEWS6uJOIwZORxbJfBOKcIXvIror+9R1NCS3j8OiLZRwg5s
8hEyqZNJrSi04XjZDHLiNdiLbI9SDcmRNY5OaF022waiTBUTholgaYucw53a
UJFNj2P5FsY95eR2Lkvi8R6afwY5IvAfgdlqUli8oq5qBVpaw4SXeg48eWrM
G7NP87qvgeprLDoKDBvzB9sNXxW4YCwCl+p+44iTMY4Gb1kwtjmdlIJjux3X
c0XYCUUuLN3GHaKirEiMx76A6Yu0pb6jP6LiyA2JaEaUleMp4kj7dQ5bR9jp
aZHp+j8FMJv831/XhPJftob437juCvT0k0Bvi7i4+r+w9nFLARQZcEI67e+K
UBUvL+J889VvY3JAmCccrFxlCiMQDpm9f2pRfYFt858hilC8dpnKBBVnMl8v
NMnEQQDonJJFMOE6nWDYjKmMlrndExVTtKzKBNA0KfNBc9M9HFmEujFr4jZl
ds9F1l00rizakz6nehyuP1Ii/Gkl46SoMNZ+pkCDlbGok3RVuxwmLHS+eY/g
d58LJ9Q1Yt8w1fC1BbGYpvQ0Dnlfat8AyZUhlR6Ww5J4aclENLHiJLhJkLcu
wKArpzDRhSJaFRDPk9LBjeaVl1EDGfpMWyDKrTJnhT5Zx1PZaIOwRvUagRc9
eWmfaIasDuY32g87fpv8Jl19eHBxOuPT/bQC4+akERhZRkhaulQok1IzMj3r
oDxRsbzSgkVegu4yGa8TRatQDNnLkWuK9PRCnUfalYqcjhxfz1Vm7HBQB/hQ
gGq0g0HWpWIy1yRH4dwpWg6o3c05VB4az4j8D4O1Bw8XchZ5A6slXDtQ1yy0
ZHYiUZzvobJA3byE7ruaejvBt/7Ms84WEbLaosA8G+1FfJe8iOOcJShBQjqV
J7POR/EwpkxAs89iFngvUnwTzF9ePGJ2fE9rACqX9dUcLN1A3nekxiz057cR
L04Ti7MIeMK+3Jp6bI3X3yM5i3B7avuz6hC/Gj8HKuJY0CxPggq6ytRRsCkc
+ugZ2SyOBQPGm9CGnmR7rFy54niYF/GLRh65WgfoF1NMaTPQEudT1dsxBh9A
cZ4StNrydYbx7hq/OSWjFTn42eLCUJzmzRrF7NrFdB1Ulv9yWJXv+6JYS8ae
/qh6u9wi4i8DcGZj2ZXxCPrXAnzKzYFpPNWLa/mdGvoOusDtUYUuaLYD+fiU
WtqvAqrJg6RjB9r7UVO664pL2SNYjXczfFIr8BqZwCavIjHo+kMZJni/aIva
sa0tq3a2Z/bvfcVr/aPNY1VeZdAnDTQJf16hi9C+kkiwx6Tcer7oHoctPZJD
wW5mh6YtZ5lppzDAJimqEh2gEKIPXO6mTMQvTxhhmt5PXNunMcC8PbU6vdiF
ELbQ+cgp31l97EoXvRNg7zuDIj3e/NrKNY5EF5gM/ocVDCWJL3jjEPBjcUxc
bZY5YN3uaXBrUJAD+19Eqwme53AVit/F36grhXuBTInXGBqRFo7ruex6QlwP
ahR+9fLU4T8r6fxM5oUQVr/6tg+AZRlVaD6TZ5nCzxoFqSEopXtRrt8XEKnr
nlsL1Q/jd+PKmKQUsCYDfIHOXMx3/C4pfgEBwIL/a4KueuGMmybZRSzYhBcj
qfJkpB1fBCcEVlKMeVExHhxIS2aOwEOuwiJx4lVGR9U6VrZ9S/cMcF6Mlj7Z
XCrar4xZ4K8oEwHIEAuVzx5LZ2FoO2zHc4wz6HWGYe+z0D61XjLlEXkxLXgl
82hxbnHpjboFu7a0qixS+c6kO1gUj2r5fhTeZDNcbRGNMPFoobBcjRP2SZNZ
6nl9BlvUpv+2AUViceONLkWoASOtlIFWOZArTZJ+dDBVzfAL0XgTdSlDdmyE
3TPUSigm+N7AJFmxXwbpFeoiFsPF2HG0YkShVso9EDpqrUukhfZnCJ1xtg7M
ip8LBzWI7jdDSY+jMUId3ALroaZiMKYEtbSl7ixz9ZP0o7lB8l8y/vthieW4
AkrJWSRQg9HQ7Fzc6HmPYaUFaC1CSVarMKGBe9gXGraZNhvSXwFNCnweHX19
a29A/jtBCEkZP4uoSfM6yxjjmz4iNz4HW4pr4B14VMQttBXJEWLNCaBoFhwz
PoplkluALiF/S3IsiOOjOli93t/OQ/bvIjsxoXwqo62ShyWIlg2aJnBVYLfO
hV1GkAHEriUcJg3TguMu/wTUQsK64rPfWZl6pgJaG6Qso/B9bvDRaelk/PmC
e9BsYAUZwOrkeHGIZDiVZ7lArVbA3swY4++sITw7G6DL81iagY1uYZXF0uSN
7Ar0WXueY4oECkSwmt2+ZvaHEtQBQsInZjtnvM+EMb6MLR714JdaDb4vEqMw
ya2IQK6xyhlcPqgSei2TJaemS+24CFCzgtZ5ssdHtjdhgsi68UCWOdCK9lLZ
Dcmt5tVOmLKFyXbA3H/i8haBuH8ImbGk5vigUPtLd+B9Je/rCR6/fTXNRKDT
YfJILyih7rugCh/RR9vY+z0P6g87t0osbaGgFtGKGeaSFnV1T6HAbRGYFZmn
P4mgKzhe7SvV1ZfVBdOL1F+/taMCW8Z3XLeVhgXN2/vj7Kwz2yRgoN90TJ5q
ZZ3f8di0HgH3oN+9GPrJZ/Ij2Oo4xojEI/3sWddc56/MmnOKqqV0NiF6z6p2
RrAiWJZq8WK/8YlHoY9FZKWhXWjWG9WGerMGSD3bNhZ4JeCtiJiktl2GnHgH
L9AfqsO8YPifLPqqC4pKOK5x09jQ+XEPuoyG/6K3cXIEXVJTSvzOBSNswaQQ
rYifTCmHxVw0KGt1MASCMZcUMdQG/cPu+L4eQXnn7dGt59COnfmtM1njnmLz
Kt7WnlvP+zktzuUe/Kg0jX9EWMtOBjTZe+u2KtjT41sGPRaxOfPGeaaBrDJi
gbnk6I4Xy7Y6DGfbsJn/n88R7p7EVHnecuBD39Rn1uc9QWwVIAVqlVAIzgBs
5B8pRAB5L8mXwiAtNvhUz7H1d8103aVZM64fglbX0QjEh/GdsHPOoMRg6+IO
D8eUq+tMkhzzbsWOMOTJq3pHBnZ+q6wfpyCNtSVEHJgX6O6kYLZ+GqOo5sEQ
blhhCBR1ceOoP8b3JnS1+Mh5oqQ8esDIULf9zMYRXdynhJj6Qbnxxt1eJDqi
XXrLOIAc0wWO+Mv3O3/zYJdTET9but42aVIr0gykoayX4PpsAxeRVd3eShDo
qrxoWhr77dbq9OgSU1+9hn8nYOLTWuxvcUOSb8p2o0/8XycdIETA/Dqbp7Hm
aIpB3MjeminPhSi/e/tY/gDs0NbSFOuY+WhwsXOqK3s6VuGIJ3YP37BK37N+
gOxoHxxJcIho+1EK1+IXkpbjmIlQVU/dyXSPdF9mUqsAH4TsIwfFoU5diu8U
ddtCea1L0GFgbvbarjqKLGn6ePs8cBO35WUpjbxMEvrSi/sLwyfVIFdsMvYI
g1WGB7YfsaZqzSVmDoBmuruGtEx/V/zZIsOmPAXMXYg/NTdnZmF78WsHpn0d
s+OR+z4pWiVIpKIeDc72fXirxmuF2UVPtYGTfVr6OJnmBmyF1DHrkFjci+YN
Hb2rCBpEN4SizNYXWVoAtUaCdeP+hEdMhBYX8/MeO4a9C+0m4sXML3oSrwGr
95qNFCWrkYXxpPx09y9La0RGUl5B/H3C0PpgEa3yBcooY5KvkRxvx+xZfAs+
THiQsMPMO80+rOY2GNsXuesFRinuEAaCSfxoW7t7eEXiYKqEcZnJ5uy6iJXA
P1Qi0n8LMuIdrFzFtOesD2PhJQLWLJcdkwGTR+lJ3lX6X8E3Np6ZugseBU1v
p7OHLfRgfRsu71eG8GzE8C7wLeAZsbsSGwphH4hfxClVVNrF/aUiHLa00Sn3
X4EAgvvoQtgv1XpUMszHei8OFLPfOJz5KBVyEemrPuI6+ahx3lt3nVZqP8/f
66zLaQIiot3aoNOj4GUnsJIYMup37SizfYBU6P49wLAuO+dtNByAH/8QmzR/
8yUBjNFlk/0gQBGqTRxdqQseCiDFIcu7PkvD76dXKEF9Ut5xhtQOxnbydIXk
7Fn2WEZNQPnmo5D0/9xzpiMdHUSIeM+iuEPsFtHmG9bU4c3F8scHnIyhWIvX
6LEqvz3RmCnp3uRF15AFJ1uL/WJGYELu6lNEEMmwaOyJDWIQQG7lzk1oFecx
02TDDbN8sK7pVPon90Qu6HSDEnfI9bmfn2KiEFZb4gR0kFiOHYM2qO6hyXHv
MFIz9723KeyV+HlDrJLJWTOaOT4+M9e5qwP4UuUKDMyAF4W42gY39ZL4ingz
m5IUFnhwcVG2CcoDON18dkFkCZucZbv035nHoIAJQ6uBLHm20wGQadlprM/M
pyo1ZMNgFbyCtlJJ9WhyJr3tYXXezbEgmYOJN4sOnvt74lJ08XPrl35YCTLU
QexUvmScWBm3eyulHO4mTITL+RY0qwQdBeU0wkXEGEKN/idyAxld/DIgf59K
rUwSLwdCV4bg3G19YfoKOcJAs/mwk+jD02lkNK9l4K1EbtnsMojEWEkvj8Bv
YeWlX+FsJwCGQznqbI9qWDPtgCz99f/WYmj6quhGMDTmr4mEiHyMG128y2a7
uCLjV31E7cwLr60wMiAxA68+B3LS9SqFoKQWA/YJOuglIWrIa6l4rbvmZjir
JLNCvY7gW+1/863Jd/xpbD9WF9dDa6dg3tbHgJGbFlE1SFoo8QoHxQi+wdFi
Pdv2rDXJNyGvJBIPPYPcebdep+j0p7g0IgJJKTDb16P7wD6mvWYYLbL/rZMQ
r6CwVA/5AJ7iiQFUUj7S8Z6/vaOu66q/GEWv+wAC3hO42guwq6GWhf6qgtkb
DCk+R5b5UrmWyPsrZt9QZARPmMn+RrljGCgi42bs4XavxIvt5VpvsNgSIkgb
mU9H3tW6Gm4jBLKmuaKFS34eVZ7wOtt7sDEKUEXKan+KKrpt0p9kq3XQXk6+
AyeV4ftnk6gAC2Qmo++xN5lnWQmRWTFtUoeEp2cRHweQbiqNPXPHYVRayU3j
CUkQVyMK47t0PL69BafzTphyGnbhFAReCdEENhVMA7TyPNz0sUWuRxJ9mGbJ
G2LE+VhrLihxjLZauQN4DPj+CX0R/IWxUjVszd0g80/i123z+nzWr30n0Zr/
BNmxv64W/LDxZ/BYazZrcPuKFMtndrnFAczmBU6stVYw6Irw9ObepVjgCs/O
iCkqIanvIW5FIiNhgh6uWF9imX+Q6dztxh9P52aBTmZloSUKj01IwB3WmYwl
i20ELrbJojmtrfZzONYi9+Mb4vJKWNKCg2MqrQVMwHF5+aWP3BWK7niVtjoj
rncOkfmuDJG8HBCHHUj0VdxW4mttC+pQMR4dcmzLkr34VYm+YkK3/nLmeEal
zCMtcjrNRXAuRCsLHak3BxQxCzT4KQ4SDUQvwNplyMyzotnb60p1i2VLbBgj
OLCy3YMufFhOMP1fq9rhiqvTid3rhWlFd4Ahhss+oJu6ttNXDAMy5RcgS0Dk
9TphNdBgAgBomRU+iIfhMWm2dj5spSc76mw8qokSA8saGSy3CL+2yE3nn+GD
AHFXkrzpM6+dkIUjJrTtlDtgmiFSItKQ3DlblrZloka35TI/SByiWLd3Ettt
Q0a5BYrdxKWZuvy5rPNCXqzk2wEWUxRAxHmNlne8U+F2hfkFGbtdu3TMHVRi
I+fuZqosCQu85vXkl1v8+rq+T7gSSpvLZ8Oy2trWNqpZMo5uD1bh5dEr+7XR
PAQt9tsk9pcNbZ5haSjs9inYNnoNY/k8b9dwyrY/+Vrjy4Ey2YunA23C27x2
h60CMmGqRZJRchLP7V0ewgeaX+l+GPMtzVs8jncMQgVCqey2Kliqnj04kwi/
GjQI6vynI7El0jhg/88NdeYfGuhr7ZtIuYG5NaKgWIzIRbbNhwSFQ/qOF3C6
kk04JoUz4PAlguOccI5Uv+gDHv/18sdoUGt72bk3F/hcuw5pEYCPnk+KL5HJ
JoVyU/DyKdJYIDBQiMPnJzcgErur57TK2PPnF8cTboRbrxWDQYl2tThAIYlw
LEd3TYuRcJ7Q5V7ez0GZAlFNxoWs8FuOXmshA1Au8r6bnUWzdDmFT7p70LDa
4BMrD12rpqbI8tpraLuLpurUVDXeAd/h6r0uX7OzlB/8nvwlgevcFbz9/Io7
Oy+rAuoT99pn85Ax4OlfVhjlRhjXF4MAs0LSxDYGurR4NjssYmdbPHCgvjgH
Ib9gx5mni1dax3VUGfn6tC/fNZjwhhs0S/tYM95KCS6ZXo5O0egpX+hVUk8S
kZoepFEN6q/4I/jqcGDsNWOsLFvaChg+ZTsRu7T4Q/uAfFTR/CnMNvpad2kO
jGt4epvzTIlzYPqWXvYAMKFlgB1xnygemWMPDO/mz4pWVNV5qsHDkHGHAnfe
w5xuJ8qcDr+aSbv4U38FsJiVCxtsuWuKKG7GwcbaYKy0TCEQPei9FVPjWk5R
u+Skr5xzJtz4ML0fZ4xx1nmLRq83FrdcWuJ5SKWpF9KJd6oGEXzH4xNxQ2uL
Bw7i2gVW/Sdez8cUQ1/ksUII6HPORAHhdG4/XgcgkC+4A96jdlmfedEV8FGG
JwZipYdFiyn5bm57lU41Kea4ciy6tEUJ/OqbzpTzOFT3dZNXDHgpGJ47wdsS
ecMyEMLFH7PjD88e9lhkFD1Lg5DvjXlAtfViSd0PgIAO49CXfhCvLfbTkEKf
cl6HFsed4dVwI5y3Lo+Pduh6ve6tBx1+gwXNeOuWPBnysEZYuxoC6n7N3ZEx
vN+U4QjNGixDjZ4oQPw99Qxz8kwAfc3ZtqZl0KcYz2bMDe02eyQm77tyectn
UuC3YmISxmeCXp/zIeQGJajMIDM/BgAR+6/kKEoM7arl/SNwqRftQSseVJr/
BNJ5QsHdwD6+QQTTJaVFzMxnIVHJZ57EN6fptS4K0HvrHmDs9JNyOyfxaKfS
AEc6LtU2GiwLUD/u/Fw0g6DZaDzuFPjHKY6B3oqxC715BFEajGY7fJsnihXb
82u3zzM4h/03W5ul5aAIhkF5Mwo6AqZ4J12CPMPJ1ok8cbAOufqJBe8UHeSY
TRRzRU5VpR099xytV4DgJq3udIRkaYAwFnibellbK46q9OuQXP0fdFYhJV5t
lwCbw+QOg86OiRrQCptRuT2B6T6NZ7rW+w8hcoxWwpSRgYnkv5RLurChj3qk
bx9osKJhgTuXVirYsGl8fkBqi+wqBkp6r+KNHUJsMJon3O1iij4tYZ8XGsJm
0kyYW04p7doHWNkEePq21wk9F5mZx75GKiXTqaEp/5inScIlBsOdob9Pa3aB
jZk0kEKSbBfSvV2f7bOOpBwxTDuaqrrdcU5+ED2FkT8VbKAhxxJ/rYbHywyg
y6zNb9WPDjV0knFFM+cDIknwJzq1Yn9UNw/tblEAJyV65S4lKMkH2Kp70d+S
aNoOipQSvH9kRgCrbwdD5VOKe4RRG8OpbOsqD1Yc0IXjSxTPVfiPjmFZlGa4
iTVPaczT0oB3yj3u2fR2QAyXv/EO/0SBT/3hGQ3nlvjCq2HvnstYBOCtBst+
uvh/PrDk0alwO6RqxOVVwWnAssmbmzlYMrWJxBZcUKxaGVUazv9FFrV0MdDE
U4/hkvo2iPPtqBRKoETTYgcHvo9WD5zWJTN4NMRKnpbGgPaiZMpwFQNDtojy
kmIEXa/AysmHQMB6Vi/Ejrudzj5mvlqOtYRPYBYB14JjauTpRdScAE7yZtCx
1g2xeR1OolGQ7JuW5BwTdKWT2+KGf/lY9ZvQYO0NH/PHCPSmNyBwflARhK1x
ThY8JrUziwvMRsV4UjLXQ56dl9lUaCwGVNuNcmN/A3vamsSeFQlhs2WXWbFE
7BR+qEha2uJqoVKx7s5+ZB+aQcbtWUKKQron8FGUn4CUWjm1G+8tmBaNMYY0
DwOG05rErd3KnBjf3Ya3wcS01UBnhj4P7w6iPU9u4xeFlPqbwaEzS6sPCATJ
dOwYOyY6tpqw00gnocbvWvyG2b9aVCUfMoAiOOW4DjHWXe9suE+Mh8B4fz3Q
IzSeK1hG90DkWMQhBJ2ICpiHWQp3dHSdgH0QldtOptmDDZEC7MGkzbvBgjrn
ngurSCriVho2rzW46Z+vNC6sEm14ue2KutsAxzriHVNpQJF+s858rk3TSz2H
BDFfClcRzY8lPE1c6TP75GSY5OoK1hz1bNm47YtjblGQIpC7rSBQ6wMQb8tG
cIwezCdbN2YdlkX1jKVYDkwEdX4D/aKSPWm5PKgOqfkxKXYHi6yVzX5oKuO6
ZRjXnCNosyEJHmCGePY9Fg+2O7JHYWP7sXehSbhxPYlP99IMhvWIpJm8eIvT
mcJENVvILBNM+kENlW0EIg6fJvUrmznhNdjtDSR/JwzCY0VagLS7R0WvZNHD
DvHb3B/Awh4lRxCRL4SO9+xZ6zNCFJrLhYkR+S5a3z+0IV10n2zg2z4hjZyj
/ZZeZOMaR3rcRVWuqYw4vVoaAyVaJ+JzvKcPZNYqqKNahvdOnf0Dnyb/DV7C
vNRsFMQXdkZsL1DBsHirqmOlu0ItLFQTxrkhTZzuSLOO4Sm/BU3mnfc0XkAe
+EOaQ8iYCXFgu2A3KtLeF7WdNxIaEuz9GVU+6fzlxzsoW4ZMHrc04PbOlbP9
inXcgONuxuTrQBZlrrFD5Sx1ydj2+z+9Zop9wPTb+E6Azsj82Wxw891GIA3Y
TDC0IbFA+XHyLTPoWs6/F7p3llJNaFiKYd5ersLr/h+vJHhYJ/+Bdkdfypy2
xTsqLBNtOytADMesitru8xYdTlMKL78ai6TWMVZhpoaqCZQcVEMRcljPL+7V
0BlencnjXpLlhNUOZK801IVdCdEjTa+W97+wJptByYwEsqmgfCrcltngoYdO
TDEvwfjXU00zrI5bHLKlWSvtPSYFs2GYY+Fa+xUXYgGX7+i18cLq0c9s01Gu
SNxOBcAIir1OrxTEGU4cOpaU3vCk0A7FvFf4r9EVIexpUBPc2P40Q6GIoEtM
984BLcaM/0EXLneiCfYfUz7rUN772PJDD5m58CHYURlTGuciX52jZk/O/fgb
1QTdjV1BJW26OaQuOSnMefOa/ATMfI6Bj6gjq1wbPEVhPnmQtflcmCKgIYRk
YGj2gO6S/U7V35IIfTsz6zVNCsoS5kPGZFupFmSB3xUXCVTuAVLO1WSiC/Pr
AjQpQMjVShyhj7IqGptCkTqy3uiW3XdzdOfi4z3oaOn16/VZdARmv8oJ/SKA
NhW+AZs95Sm77Z2iItUbdQaKEusT0D9NUlz9Iv01FEojxfIIXHB0f0HM9zPU
Jg0OiDjR1d2PzAIllfQzP3cHRs9WTHJE3Ovk5YOS5ooQt0NC8DQNjn7Xat4/
bJ+J2cJHf6nFnsXJpyis2mgf/t63gh++VTMWQzC6rkJxXgQ4EmCN+WetMfde
gR2iIYmlxej1AuP4b5TXnJVjRPaqHhO6SQ61d7uj9hYqCAVnsGmbmYgErOYP
euy42Cx4bFBdQcw2E6K9adq1p/A/mKy85/GZf/Meg8wU7StolCF0PZ/Eo56/
fVTjQEIAZQVG8QZngXtmJdggxmozyQ0BraBbOj0Mwo4aXOp5tYspNVbA0HnP
ksJLlBx8A5ZoG89Ufyh8Tlk1wd3DbjvUjrToxToo+R+6GebO+pwQPyzNxrSe
ltrYgL72yBDoR2UcBFKA0zE6cTSMCwt1j38E7bbiW621wrTLF8QqfYwziZBX
9zNsnGXGqmQUBLpP+YWbQ4PB+wgOPG1/gLlwvay3itxtU2vdX9MK/dykFYWD
H2qBCgdkVuBfMza9DGTiH/1OQu7Yh4E2pBzyt47xuTzrELGXccVbo42HWpcT
tmSGB0UPyOa4LF985krvPPj46XGTFODdb8taF6fWFT9iJuYPzOEflnfWEfmd
TISSNwTXUl+Qc8fzLj4w/XkhnmLE+1qqZIznl+xgj9s14uu/OEBXxoSKkqZr
qn1LRS/Bqj2iqL0yuGcrr/PgFPNZ0oAnJJ3CunWN2cAw+vCUV5PeuS1q0OL+
1EASIx6nZYGeGgN20ChCObwin2hx4ZLAO8lwBjVK5ydXPu8INJd7t4jmffnX
s0ZB31l7P6H0iPy1SrasNQOoP1+FO11FgYiHYftOS/6LI2OdI8x7iwqUhkYv
PFVfvKn6OzadczWUGS12QBZUUlHEcZpGK23U0l7Swa4u3VeEnWxOuOLLN5qn
yzfczZOmFQj0VyCi6xDBRvSLJ4sVItc+SMeSrjalPFVo6HSB3QPx8J0POZJq
pb72XyWpTbWQcq4xlwrRdAg1JYPlLdh+ZksurlB66YcZxkhrIuiw1btbD2Px
vJB9o8rPzE8h7Xixd/5WbJ0TtzHVZ1F9I30VcdgcGFyDYbykNY6mvaF3mcEw
zuWoGl9N5ND6Y2yE4bH5rRPairla1RY3gZkULoDKSiga/pWa+cL08kQn+Gn/
7kdKda9EWM3a0g2A8lYnLN75Z1K/OgTFinRqNvam0v0ZhJXUSIPqdLEb15gJ
z/Mqmv8feBUNE7pgq6Kq0FuFqdkTn6kH1VAyRfficR7YckqebY2u92AJO/XV
MXNN1kZyACMupXUZEHCJm7JDkn5T4eEvJ/1IhnxMpgpLVCcWNJEH2AUz34ku
rvizHVN4Kf9lVn6h3ttNYYaApMTwGCvfvendcQC3uZMvHhP4W6EjOTuel5ZJ
RKoMZwRq+KyLDdy0ZCepkJtKrK3Zej4IxH8Mh5LRnb/ijSo3FlOmvcNqeWLS
t8AHZ0EMOeabBuk+ZjDkM+miiV/oDWWThalr0+3XLU+nNerk+KXfJkqAFpLy
EniQ05GaPKQe1NwNZawjbBwWpIVn1C8mH/nxyOcm2ndAj0MLNDRPcTKpVY+O
0Ytc8p09eq8shCLqdimtCCc40tAYKXwAF4c9EnK4NT+pP0sPjGIHY5VDdnp0
19ucNzVS/2c9W4w8fbdqnl7M6mHbsZl93SkBRgRW3Z6RYKz7XeB8uzGj2CNi
IG2/vStHNXQ8ESscnwOFTWfk85Zzo1k2lkdpOVWbdYFJD6iI/+Oyp/OrgBdd
8TLrnRJpgJ4tXVOJ2aSx9L2DKzJA5+Z6dT8OlD6T0euOlBhiyuG0pMiELVCO
wdwHl430I+Rg0nL1+7n4I9fS3G/LjbSDQhfOBp4/SLNcZsVuice0OiqKGhzQ
HDsmS/YuTosmCY1mwWOwS1xVICLNCSvzEhkMbg1kja6S/SNNPgh87eVndonD
6zpm2b2HYYxfCbjw7npm0bo9XMgsZvW3fNp8XMAb5mKDONLS/ecMef2KT6mA
AzL9Fggh12LY4Jyp2AlaSpc/pDbveLLfx4Wm6CBxYNncxGTbS9T9P0MgASmG
/QdO0sRlAXhh3IYe1QnZaQpJpPcyLFVD5xR07yAJ0yuxyBffm//zmpn/yQv7
lpz5/kTfz9mTtuEVpYoZ9vwepIzpXGA4/22MnBsFa3QaSFxUejp3MzG4QiqW
sGAYYp2+z9VbVdp6cCVkJVtfUa8mGxbRZZOcR0wK8qywG15QlBwhb7IJ1LqJ
j3d1dAZL8FzRiKkOqKcTyCdY2En6MzWqWfol+YfkQZUQ3IxTDbAf5dtwhQvL
d1p70ba6+xJ7XutR6zQRPsNf2e6zlIBCJpWzcGMEgZzkE4bqobEUSGBbWZRC
Lns1iikgnb70dvv4bM0v0kVRGko12jJB1U5WVjsOyHPWWDjbRx87ZVp3gzkO
F+dbBUDQxkm19Fdu1E7MR0J4sIXBz2ET2NrWFnfYN8aVO/DeSKpf9MYLu5R2
c741kkh1Pl/m12CjlINKqwUz4cLGgC4THoOiTbdkUTI0y4g2ouk/8n9dK8GU
OiewFh+/1TcqoQQBOW51ygcnSGInkAlB4d87PXhARMSZ47hY1pOYfqCe+mNR
tJzVDhyp40sjiYdAOqBF958DfWBM20XTYrnNDmoUTdjO9bkM7AndqXDt5wXx
Q40gIIRgLhSUGHkU9l4iVTzZgmvNyOa+5jetx8QB3eC/vTCs5HZr3A3LKaYV
nxKNjK5Q0J6rXEb2gJ7pq1lFe5V7+Yuh0N0tkcDv2GMjUFSPb2EQm2ApwgS8
Umh4Mks08IfiUpF58N+iKa4F1QfIbF3nAw8jL+kx22tDya0NyDT/ld6Fsgh3
yLRzH+GJSdAbEB42Gj0rXx5FH7bbki0D9Fr1TDpxh7mkKDSN2k3Hk4rO7K7f
efu8HfjEENFmhKA9LLQqkhSbuO0Gb/rYbALI75RiUoT2ynT46YdkrLnHDMtK
VYJGjyiNpIq1/oEPFWih6jo1P+R1OpvkS8W54B3Y1v8YJ4330lYoHdn7wMV6
k4Gf0T0PlHNNyha8yQPe6cAcbe7uiDIYDMbYUHbTTsfSybgBs5OdJ/YLGvUW
lJd5qSlXXRQ7qN185qfv3DIIk1+Lto2hISslQ0ttDnNjBTMNlmf3cF2vaaUW
bh1pzJ6ohw4KvTogIjZ/Nd2lijjlFdHVOLdg8eE6r8w3A+mTA4swqxYzJfoJ
kNBLNekhdScwsZJoDqPotttXE9SkVKVQeNwZErpvcB1QHYIXeZWmPzk8p1ML
3/LF49m+oULfLrMHxPeWRuQZrF8gdHZ5v/X0hpvicD3AclqPw1lU8uUygGcD
46ANLat+/z+c8MXc5ZGJHJm3+4TsaP66YycjNCkupD4GzaiCVjZdGqcyH7jO
Dw5u5Dy3tWiX83GFmL8Tf6+NJcNLJas3SNNVe4QBxAdZKublH2Shxhh6AbYl
ywpxPhV/LyV9Uo2/rFhnxZIf88yLShEaQukkRBCCKG89wYru59izDAnUDhQY
aQiEe/zuf1vYFMTjKo2/SVmeEcs2H63tDoWFVvXdHgipZUFEa7w/lQCnhOMC
eDsZZG2hSZJLQWxQSnNGh50niEDh5uAPh9O6G99roZGxjc/D9WJWwyIUL4n3
WkT4or/HNYw0rCwLg3tTcn/0nWtK+dWDyfSw4Q4OxH8XMrcCzsXn85O5eleN
4fyZwohCFzvNU33U+5gv6YxdXHj1AtCjkYXJ89aardMJA6/pYyfYlc0lsWkn
irZ/03FU9dDBVMU0DicBK5wz8IrRtBv3pRLyw8vGH/hdmiuSp0rIlDxKd7zV
u2F/tTrYc0iUkeEtcAb0mq8DrJkt6mUIIZ2+RMxD5d0drTY7XSvQM04cEbxw
yRqhVnfhjUE9V27lj7b6e0zjKNv+39ziQLxQc/eWIzs4r3cc2vBJr4Nf7BXe
AWWdxhN5h/1/yn1OGj9CUJgvNZWf/EwvtjhU0r3oQGsuq0F/bKxHJEHqn2m0
x9IADrdrXvlgB/fGoE0EAUPcsqr/SLLMHx7JQpa3CbWQhpuKRDlP9WnuTjCb
5hUMeHRgmDgu25/KNx3LD0tUqhICMOMk3WojX87nXKVOi235wOiV7hF34NdX
ShsEXMe+TCPI6iPf5d1jxC34voc0PGOXcnltW2dxxq7SSnQpPurmP2/2uvlD
z/XmncovSNwHRiqmnc//tThRnYkXUU1w+WmjnCvjibxV4BzmIgT8AtV3d5lo
r+Xp5fMI+0quqinefhdLcqbRdySJdhaUcaLoJrltTZwr+JAY6ZWD8CECgdb3
zzk0ASxu9Cfh2cdLMUFQr4eTUeHklBgsSiubI1Zkk2z51Sp8600VXYPyf//v
9NHi7sYvpXPGbXpqh5yCOt+mMWqs+W59DHxCHbemv6Nwcaw2bG3C/G9BzHBu
mHLMoiNADblAIqfyiHjWXkJnGbrVlpkU6D2pfRiATqWfKhzAcXw2fV+ngrnq
nHgO5Vc5oWNsgVUEXyrOfzZhwvbWBGu11y/xCQUdvOctIaZyn26Vj5vWrwg7
yqSPCjDyRGE+1ecU5dA0D9ZOw9oFHvbNtSt9nyIvBRtUN0Auewv7wdKDF9gM
NigdBtlFSpSQmjBXHIPAta/TOZAC2BGx14k1Nxh8sB6DblL4uXOz+OhNojxW
rJLRZpd2slXP+X6/g6mHbZqunsyQBG7lDhLsoHpaxejrPuKcV+t4aGCk3cRF
B9kXGNkBApPknN/ASCeQSkkTrody6z4AO8vf+XZs8UFhSVNy8VycjYTTviD9
8maZwQJXhApYU9n8N/f0ARiYLWm+/w9Lu7MKFVslKp5g65P50W3eEm8TZeL9
y8gl+xOv1yXoc9guk7jNs9rIvpy4fQcSCKOPLXbIv851Rc5tgICj4rfkwvTv
hEd9ZTh2CwMBFo9UuQuWsLwZ+Y0Lp1XHhDs1HSyETreQA/Cyo6Za0ys56vYi
5CWETzbPkEtjoDRnj+slamylW50K5lZ9DF5wk+yV9tGf2O2umf23aGKRJlzI
rTia4LRFgDwz7iNn3/iqm3zpR4dHqwUKrsy9Be8tCfbdLfJKUcely5CuWRMj
BBmuSBXD956g68oNhXvm5QONrd9W8hriBhYzJJtT4ktyIHhtQFPl7B16T9on
+gy8PG/ee7go54+wUzgWNqvYe6t9nNq1hKYOOuNmm6lHPXqGc8XpLZAZnE0C
E+V4xdMGe1N7TdrKfVJO+b86vzCHRfze2VwuQ51m0kHgBZJ+ho/t3TpZPryr
tsNERNDbr2hyCSjkE/ixaE9nByNfRl9uAvhX7QFENBC/PGXiz8D6E7zpyLPe
hNbK12gKj/41w/CTBANCOA4JUBfF5rAtCd8S3/pTy53wuk9UVsnWFSLxie50
P56qtPUdpCSj3E8wUm7GOzbEfznnMlOUZVOZsAbA59RaSbxzw90QkBZUzboT
meLtPVN3aj8A6Nl/b9P+yMJj+aOomym/B0ojYThw4JtpZHuu46dV+OEfLIKf
x2Z5JKmOY1J0Mxvkp3lBFZTOObw4mHWYErvmN2GNsNcahwFUrSl3kd9/Y/9h
CryRLrKRLdAGhm74MOd8WKatti0n1M4Xrkm2hPq8E4At+F6rC+iNsk3aUBsq
p/eRIkr1VWaHk1MG7zTrsKC/Hf75msMUzbObucBFl0xZgExCJLmbVwNLuHjt
RSXr1ngjzASa+K4eTshBfd308HUxZY1HXw8TCwZrZ2GH8+dTun2r2n47p3jO
ur6Jps0zPNqWcQhVfzesVKBsoznS+3tmVBZE1ULk9tA5MovS6WfYnwCOnLbN
gypQWsvHmmy1nJ58bNcSuVyhn4KRyqHXfZMwYqbXEgX0YGcKzDflrO42siyp
za4bkQqxHj7o2HyUAKwkEbTgApTqdQtIroEPklM9dehK8G8pKgqb7540j23y
5jeT7ROo0CZ4nMUYDoy9RInIPFMW59Wo+iNO/zAKmDQMygKwxMzLJaYxA4aA
jPMBpYIXX4hrx9M+46LMB2jx8Spf2Oj3nKFastKyrpihxEBWLzu3hMXe05w1
ju9Umnd8AJGAAWZXSWvWVq5U5Xd1bjJV2HUcl0Ps0f8sj5w1kV3vRph18Ndx
GBAxNL1jg+dLSBTAnUWzzMnF5CBgIHaWmpBvQPzvn6o67xbR5ZbsqoFmBXW8
PRSWJLYLjpyq3iEoRVh4dnf2HXQPKdvYYbqUl9MXtaQI7OYYe0oIJGauNs/k
sWHmzPXXDIXdx2LyZVpVMbufdDe5KVNANjAv5oRDQiZOPVCly8YuXK0mJtbb
bH3NJAmGLCigLuwu2rIqY1A0OpzU7fxR/h4bC/DiV5BsjxEMBdUhlAzy5bta
U/JumtYIq36/1Q0iNcI6GdwUczMP56RDg+YM7U5LD6YJWrSz/XO4KBeS/5rL
uVaIKu5uYfm90mVFZaDvfvDjnXW84NwYg1MZZLcgWjyzTvH3Bo5ChaniIU95
HSGZRqtHnAy+Ozmml9ivElCnE2qQ6mU327H/TSe+XjGHDJieHTnWfG1hLed9
Ks8DqZ8Fz0j6mSvVpK+/+sTmlRrdieosoyZubwkpFF6UA8jYEUb9AM71dI+m
lBF6O7bboNKUJTSWOVBWvgDpM85dI6URwx09HCmUs5WiHlyatge8YyXKva5E
k0qh9GYdO4XuNFdCz2Dzu6bd9la0O7GEnRuipUzIoxcpDpZkQoSAUuRtIjwZ
WcnFICpz8yXIFq6xgiZKUL1g+/YF9w2pPaqI0ArT4sPub0x7GstcP6FfeSbG
iTb0iILFZrLzPu9B+m9mUh37NZSHao9kEBIg594Z9TIVeq0zNBmIXLET6FEz
EEALKNahZScED5lLej/a/Lt+/30895rzDk5Cuu3Q0H3vb5Tr1iHRaunqrLCA
3rf5SoTdcsRRciARP+yvB+tFyOmBs5uFZ73jmDG1A3p9QbxMrrzHVeO+FbWj
15nbtTELjPjpscBm6Q1jYN+wkZgt/eS8BPrlU4XNOaAgBAbqOo0cSjJ5zsWW
Q/cZfuXlNi13PGHVJa99062uAuNUi4A7riPyDH5BrwkZdL6y/0S2N6EEUmRB
olAHk31ZaD3hYaadV6Yx24JwUVZ7j/cPt6ES/ZvoWIih2qbZWAlP8Am0foyR
9ONDdLTQvMSrLxMO7Cjx90hgfUxeYTxdfgjg00fO9cWyqhEcxRsDgzNUwFxi
PGhE2cgUR0Hcgs9GT/OJN2ay4mdyNZe5VFgTnmw7TTEZaKAdGjJb/Uv525n3
l90XdthTusGuamGvB3htYRJ3ISbZnj6KzgoT0pwxl9vtx3bPDxVSQcKojhTF
HO9euaLdLAiDaq22fs2u6FkoDhXuf2feq1qu59q4s280JcW12+KP6OkkmQGV
9VeYrYq5pCghHCwhIqrX4WeDDfA1GLQVfGu3hGfBYsu2IFvFIPm4HgwolQfs
ubWeKV/WW/m46Zmb0GAFXti6nct5BIdwTcf/XtoQ+MGwUUELs/9pJd1PSUtj
6vcrP7lRMWpjI7qwsAfjL4h+I5zDJjd9IQCRswTGCweFJFhbBmmRpLSyhmSJ
7WDWHUB3tKwsadwXat5hzGSeZji5SyGZdSffkxboTtnvA5cv87PrZ/g44A9V
B+/rqQi93zVgXhs+fzi2cRUPW1XRWgENNDTzKzocF4pehK+jAEp7MfWO0Boq
KQ2FSWNHHBMKQIf63jpjrZNIaff2DhEbgr+Aho3BHpxNbRFl9GAaOGZZlRFl
JRjgq5kb5YyGa8XW99GGL+/RU60Wva+BIO6G6rUPftNoz2uxEPrx028duXUN
DT6yAbUMlZh8gJM89HpnKDCiayOaiNIsrO8ADJjejMaEEQf/BLO54dXeiQvs
45dPynqkx4W1Fa68hJV9S/10YTiEXhe6cDnedCSWfeK21FGoO+WQC/wxJm5O
El8RdElytzRfAX5+nRSV4y9t+2dOqk4yBAUeDHvu/JpimHrZ6v9Hm+7ig7jn
xt4fLqbXtTfC51qsSyz9WUPMOXSnW9EYX2tXMqms49dfBQNblnid5F6c1SRo
rEqMIq2qbm0/17sjVdj4EhBEfz6yYY39f/rTgTQeFKCmuyTuJp4ggKm8hGke
ujrb/DjZYW5eDCrksout9p06dZnPiPwAOSmq0AWaCgK1rLa47la+YSz69rrF
8ZWn9AXaMEAdNtJknPw25TxDcZNB418eynudqr1Y3n+OoFPS4s+UVNXQuS53
5YK+HtC3YkpgZ2SKalypCjI0PYe+k+NASnt9/dDxBnJ+HKa62koptsBqG5iP
1Wfh7NS8ZRXdo9683j11TtRSVF+n+9QdZi8jC99mcYZnJKRI7SQIQuPOzPHh
xgrsqisEkD2qF9L0/W+QbGa5bXIqV5L1InUpd7eyFO7MdBiyYezvnyTxUyYL
mlCzYLnje/RxoG0LihQXf3oMiGKN+mMer3ycRPww9Cgwq3gnpRu/spym5M/I
K/A994oi0dkmqQhyj928nU5zs/WKO7WK9InJ9rffhtxH/qGzsbCfkogqcgPH
syxVhMI25qzLEQCQ0cOYN6mzOmvxurj6TWumwpwDhPZDr4qBl1750eezeUrX
d/j1e3NMjzvRMxINlB9dsElP1kZhks2ZrKLZFfD0KV5Ot54I6DSIkwOJRlE3
WyKwRjeJ0id9WVIhLP7inW68LKERZS1zNTiEQKlmOa2iCqC42WyiHhczU3lS
VNd2o77AgU1oibwnkhBmX35rlXs/amTq1vDTFNEt3t9FVnUqVtC1+8xbGTnl
LAjannWeR2pzIyE0yNrKGP0zJH+klUpMvknm0G8JTEwfVn5U1VVixiA3XnMH
gNnQ2k8pkAQou/V4UI6SEXLFzggN7DOoefWciNAd2ws+Y5lE1lglQbsOTkKh
4WK1eiqpMSJmTzn6lwXMGDKYSroG58Rnbl8nfPAVDe/27VdbEXuofHP07Y/2
1zSfnzayhXslCVHggwNNib1jbdCMWayBAxOWucD36wY2heHCG/L7CmOV3AoJ
hCjOL9EUO8VueBV/TNS00SvVGpc4egQtUpWBvMiGE2moM7ePVyaRXPdkWbLb
1VQUhMrTphnAdNrgcYW/T94CkdOnbthVN3D5F35XZxxqYb/LIzhizU7XDdbP
W3CFuJX/O6TpXZtN52NblIZDnD+AW3LexyvzFR0ofGw0F+IEIfq/7NacANGt
jllnC3IdeIdidYePrtZkGBusqeltglnZ9z4+KKtL6utkkiJ98FXu1VW9yF46
rATXefqrmEtlW1znEE2tO3slwB1o+RYGJz3h8WYDI5iYgLmBggWKKvFp+YjP
M9h47vlpK1WIcl3GpHDA/n9SwueS1sLWrl0z+jwyclbiKKuCZoqqWjwo2NCI
CSz5K+e5DbBoKTLKZ8ar9/BeH1twyTOt4MbkUP4wIhBn5YE67jeyiXe+Zele
VBMnzsOO4qR1CubQDegTYaK9k/C+9ZSH1HoA+UEpYoly3nHxzlp1NaN4o/cQ
8Q2ZsadZ6xCQQvvF05P+qesE6vC1Pbly5H+d2b4EKRvoSxPv/NMwfupueF8P
zOywWNN0gWnVd3qhPpufb2PERiAW6gtkveJ5lxzpolq7Bno5H4FjP1MNp4oj
Sh+fwcr67FAiKoqrCGwzCdu4w4p4+g8sE+F9GRPKwiD4n52kRE5g/MFFCAOE
jH/dQO1e3/epnTdEV9PQ1KkSEy4MPHDzWouqNUZPvK+PlzDWflaFpvOq+jCA
pkgjBlHFbV0un+uET5YaMpKdJdzmoVipoY3/kBylC1vH6GApeWbFpt3Jv/hn
7kIVRwQ9qKroaUeZJahOZOpsnzM3NKl5epMw2FMVG7pkQYzRPkL3AL/HOoRk
wiEFWzArK9nECC7HFD2P6fM7g3KbvXcY61qelCZU5SManeEy3X3y+Ess+T7x
G3JLpofTJWOd3KBSfv0dwpqry5KtyH7y8RG7uAdL2aD8iPqxpgeu3oELkvn3
9n5W2FiVr5PYhwv4uo+KzIkOGU40yes7W7tbS8uoYG4h1qH6LGfYKQ5g1lXX
2JopdnR0pz2SkRY0lnDgDBBatN+nVtIPhdZoLofsN6ad1+XAYjQcAhnP0dv2
AeDwgfrcaKNvw5rXKBUiMM+9nMZncrdu7Ki/prpwYh4jX8Y4RM+AfuJej+L1
xPnzb7V8PbRGH8Snizfpr55gnJ2u2Te61KoBohc+xsPUpjgdBgG/lrvYWtbY
AAqZvwbvnKpuJWAn7o0P2P1fXVm7aNU6iknJI388iNx/jelHcDNfYCb0kZ/c
3IUhes8GN7rGu8wUxkH8fbeYSvjSJCyXXu2IYA7hzQjSqknjhkXG4IbOK3xA
3xWeXxhyUTXISI9HpUU1/HhM6Bh0c1tNmLcniFA70nliPeA/36T4gFa3+c1Q
VZKqqghuRuV3+EzJPlSs1/w4y1eaFlrJbac3/zV/m786s1gkwjzY7oE639yB
f4Q7KfDYb+s9h5cgpTlVlEEDTiAxF4ZRonyei7JMBLcGn7Hm5jA0bvjUL+8n
F8K7/YN41rWMYmtHRf5VVK1mTWrzVpcDkRqtaidhyOtvISMB7oZ23wnRIF2T
W5em/Xa3BkCA0/D93/P82xCgSJtHAnIqc0kCQgQdsdNu8kFutLqg095w9WvE
S1IsyWimUo8A9SlxSanOcpRb+H4V3hxiI92KpMoUyd/XuIdNuj57ZFpQQ9KQ
OYJdF2Q9JfYAPNmzrATgYv8NfznK7WZYDzpehTS5OJUkd/n85nohHDV0aMm9
tZkgquZUEG4iDtAEppXASHt7LL9Uq1MPq0nUhtnYgY3k5ReTHYIWslRF+eH8
Wlg/D8l9LD2i5n/Tq7HODIkHNMBZWCBxuY1L4/+2rNBQ+8U52wW5uEgoo/ql
nGQ553pFWUcxnccIr7kgplcJ99wCn8+FRjCynHogImc+2sm1jvx36EgnQwXA
9SgqJuAnY4R2bMj+tQLyWGccgpWBr9wWJ8JShSNcOXiTnRvhF3a2JLXfC7h8
E37+5rF8svoN4StWErqhe4XiHlcMfaFgxFVluY2SCC7C2RqfZnuxNuHaJ0JV
BketH5OUGGoNyqpp3kTR986957jGYl7MY+1kDn7UPM+HzCL5fSawtguaMnYX
Qc2YbO2CWxsEdIocNvlmRQD40C9aHvU/91I2aW99KX4K2W35TgfoQOYuRHc1
aBbm3b9ZKWx0y0KGNyb16wo5I0LjsAIP+34aqM6sosNJvkaVKBku3skHouL2
xrHZrMRQJ5JJKGGKl7JEh1f997CglVqIkg9uoVkUeQ0rrOiUf4oXkqvQBmeD
YSydi44NODIhs0zQlwzuL4LiKz0SPx9C5Wv7P8il3aQ3uhAHMXGUeScOwT4e
+h2Ebi32gYmkNFe2CIx5YMCaJcT0OOc8oXNACw4MdIaK3j1LI0ZdUC3en5F6
0/MSaEs1lW1v6aT6uxLAAYHT28rVGZ6Kl2zs4emAQpjot86NfsSHKFjoT+QD
TJgxqrGLQ+1CYMkgXei/RJT8M2dmXgNryqr/7mYM7NSOvYzZai5HSyJFFIZH
bNB4E1AiSUg06Y/P17IhuklwuYou0kNYn5Yi9mQItBTYAPkCPCHqEy8wbDxt
QHSZF3wtcHU9vCAu0HhejL+BwynQlBvylsZj2ZFY7fWn4wzyG0smDgd4dn0l
itKpivk8LVctAp+YC+673xMIdOyRZkqMZe5fEG2AUxBTwxw6vmfCXq4l85XN
2jf9f31AXpsiWTg5Nh3qZ9k9JeZ3TuQZwXnQKvLJUKEIaq35TDwURxGMZ6sN
XrxttJKqkmoeAXogPjZ05zmf4WvmQh0TTjbDmXt4zEUvG3LzTmLJPCEuJwc+
aJIR5NgE2/HyI3Xo42Jm0M+cE6pc2tvSkDeg4ksG4Va3iFBKA2FCmfn9Or36
ZRR4gAQy0O3PEBFEq3fT0ehdKD496BzT/V++34UJX9OYglaasVJ13DlNJpEF
Rp86j8R86sTXxJBtbYVnf0Uo6VVEXky1Z+QP1kSHZLHL3Ezh/5ltRqJ9J8TQ
M4aNxVF5X03VenKFlUEGrfuM5T9UnlUN4ri1V+RnNSYzG4IiM1FWE8btWtQA
9Ua+8HxWdtpb75aqN5Vc3+4FjJT1hHdSIl9Rh00zasnmVC77Vi8LkxbR3e9B
iOxKImP09DAKpXdD9ItTkaVBquKyCu9IDoMJ2+ngnNiQ0dSxmyXGBV+IS9dr
VZBA0X4gjjaIi7cgk1gNjpzQwnpSQJ7Vdgnr6NnRa1NlRsBtCEjxosmhyUnC
8PLLMW0tdMM4jng/C+9MG+1OoPD08E0zd3FOwD+gSqpUBIWIS8Vp9wmlLKXe
p8tfTQ+HqHuLwjqITiN9+ieNVzkoZnfKcA+p5WrlQ4O3ngxOqOc3xovvGTIH
jqvnHnjjJLl3g5RxT9Pf0sdRAb/uDkCwS+52mQgFdNxGOYVwr37BdEdvNSXq
QdUTt+VouLIxX8DDYBhIMr68Se0g8lWEhDO34g9JoEInGHFlmImO9LVEkIe/
a1fPqejikfHFvWFk1s2C7cykzorNWX9Y/igJNsoAWE3/W3nEtgmQNgXTeAgV
LQgVLnY4IDNHJUKMc81HyIAIOVSEobLOxdfNQdJsRFsDlQbq7PtPRe8mANc7
bNn93J0xxVHxYgHqVlDN9QJC25Cex099bbBjUyI8UEinkFlgSe39iWMt29BN
gfbS1tb3Rei7m7UbMbF9eA2Q66cBHJKwm4oyWZuHImqwqmqBdvbRdejUmbIz
Tx+ON0+/PZVzMtxvwsH4w+bm2jXOQ8qKH9FSsSpL0i2c3WGP7KIntOjUCh5B
iOAYJiKprez9tFZ2KxCjwnuUSNRHkPMZiLxq/se3ACOKqdFsFAxkFsGUZQMg
pDwKdJC3WkO2LzPAeySVuDZJabGu+i+jtQ0tKrYeqAoFFkYfAVVUqsg9kG0m
cNNL//LcEmDHoCit2uX3+ZWlxmZFv4wFQT84nf/AApbqwOnGJuf83TdYqB1E
BDlAm3YVZo1dtPSA/iQleNfBij+OHImbI9ZjyMBHxwJCqCZ14+3Kg4T433qi
zQtzbsjRe3vIjo88vUwwvYyQOI427iCbsTAgShek0UQpTvtUgrWY8yGQQ1hC
Cfzml4ESP2DLLpmKC2NFE2j2OXGWNA++WX0lfpP06VuZlz65KkmZ+Xdj6K/g
F1yLKOfTs6urlWuI7KqBVUXfa4GdhhYVyfr3zeyo16xwuIeUGPzGD0kRrH10
pqwJxgC2QfVpFRm0i+oBY7eWWknG+A4rcqyRvFzcJhamGS4febpIXTyxC3ws
2x40vMpyZwxGrjly9I56oq9xKRW50fSneY3qSJ1nZfeVOY0dCf/ssmt7c1QS
fcZW3JRkCUYQ29Z4QvHfyfGxxVRvdkNu5Mp2h9cvIDx5m8+VnBYO7VrBLRJQ
QdnZ+1d/N+QMqlVT9OCUpYP63vQLOjS2buK48yFCQx+t7XZ2vMlSk68xDhDE
4J0JGMQgcATUnqvPcHWn15t26BOLo18rN7DvU3CLgeOk3Icv8T6v35qd/Pe/
b2qQUyDSRKX1v685zNCdkmDzQYXEGmYg3B+yWkbjp6hmxxHI4sMHpOpXMIF6
dWxy2eYrdsa6c1H+fH/bFmmJiYGbaxrOGgIq8RAG57c0QWdVSdg1wjxsaB34
Carfh1JLVDo93h0I41CQzNhXXhCETytf3E+LimFafAZK8fND0PJEyCI6JcKt
7uWl3+a4z/il7fVTVGEU+8xS1Y4IYdlckLSyPsQ37sDpjyn3vh4/e51SDVJL
4BFJGBef4u7oIzNOOeZr6c0oXGSdqMVj3wrvCH5qR8JFPVutAq38KRaiKmd+
udNEJHA7twMsn0TtvEAeC7Dg6rpKWnW/s9/vC6oix78f4OfYsuFOoEzdvQR3
wVFnCVBM7uQxAubzRCzkVFZ28YkENfMXUIJumjs76tNJeqlvbUE43OkEEC1V
faE7NTJNrnRX90W9eBZLcEWujh6BNMWCXzXaG9JS6SxCZ3s2WlU9iwGCr9TR
CSD0IBThrIKW9J8nfruMCNpNGRPMXvBnYb0tBP8Q5itGFhvpcXaLO/kmacnd
UKalKW9uJiAm9z+Cp141Er+cye9P/d4WDNnINVX2Sb59H8lDiiXDhRglmMGQ
nAN5Y0Ck4E8GSPOMm6jxklVdmCw7bTStILSpVNOgor3R/C2IK5vd2318VnLa
9Guk029xu4Czh09LIebmJuw/ep1dedg4k5XxKzuBJa0bCONOGA6kIOPM209P
VP/9QGaLPsub1fpu36VwUghrYw40PdaDTY8b54pIRhlo/6DZVxUFYjT8oVqH
r3vlsrbPPmkMuyDn2jD6s2G/j0J2RDdBdV5RYQ58bUKNOBfTRrkITUsAU51X
wUkZOX/LC2i+SiH4u8Ue9ZWQr+ak9tR/CupXoU+pPLU8xGx0bqBsF6f4AZTT
ELfKxSI7U+YIC0gCJE/zr+m812sy5LRL8dKGU4Smdju1zQXTatpp64ERborq
yEVxgTDUBEXs0hvAzmGIfp+St/9HZMJv6VLUpO3iTSrA0xcEkp6tw2/0OkHo
HNbMdqNhXKi+XgF05xup8bbKjJG0b5wirudAiuw1rAo/0VyGH7N6xWmij38u
GqsVXmCz9zYK1v5e8fXb78x6sYlxMtsOl8IASALWyCD6LTcEwZuFtz7sSDb7
1vsT//IfIld7sG4WjBaHGsQ5G04Vv4g0iGG+yv2ZJXMn+GMob2vxXyjw1TA4
eCF1UD6M1urjn+6bX3P92TGvgTvBfD/x7D9eCLt+lBoijIeHLoJFzWJB/95E
2DZoyp8hr7I1bujFdNDss0H9LzfHBBp1DuYr6pvZgI2Pi+JOUbHWD1dlcpJW
MG695E0G33/z1xOKYrz7iv2C7Zkd1N9g3PPkcrb07YTzO2XzIRCLumjgN+Wm
FOlhnd3wczYGXldJTIGA7dEELF3/b+abvR5dqhNjU966bhn/jsSZhr1o2EZb
inhYpSJEJzvxHXKiXhoE41Lsp0x5Q0tQw2lkaye/45We8ujILKPsWFCSxV+1
YungtRBCyjftpnXECcwo7EiAeFF3q8QhzFbICThCDFL7V0Y0STRy/uY/n6pP
4/W2xHB3CtfmSfFutH6S68XTzrsGAyOxgthxK3xfme59wTpyXchCEAtwCZfu
GBmOWYfnfvkOG9GLPpZP+9CmG0EPAx71UYWozWoo8uGfNJKXIETsu+qoMHsH
E+p1WFBO/0zaDbeqe0qFJbCP+Zcmb4R+6vVhdpQg50DtfbFRnUONGZJ0DrIM
Zz4HJHZQvHWVLA/OdYYWuJptPvF0VyAkwdShVeyfPyW/mXKRqG8RTan+3dAs
MDx6YsYm2Jz3fhovCdTSxUwhBg0lx9+eqi1kIql6ltXHeFojF9J/BxuPmpio
WeOq1kI+fpNj0XzeOCo/lfFgfCu0E8UDxsasJL//INGmTTYLm2J2OKltiTHY
p9ODKI+pev5Pk0q0fLTdBUSNYGnWjpNk3P1wmKp994UB8ekaM9HSx28g3RIy
puv3otjXP5jpXv7ZAwdY9fp1Fd+TrWudKEMa79NYidVMZligp0x+ak9Q89Rn
jHxSgd4cxqxTfDsGtcpVQflX4kgxOduddhgyfk/J3f3ADCPfyNDxkDvzsfGA
cwkBS5GAn4vkvxv2oQXqk0Bo39ME993mJ0MZWMIhFu7jVG0kM0/dEzFDGmLG
c1wCpFXtSta/vyyVNC+CoOncHcshZ2/j/aBxN7CpFu0Q7ZYSVl+W0lILOZKF
lMih0bRCK3iLDjnIo+4k03Cc8rI9eAFDaC2cEwgpZk5YOfhD1g3mI/z9V1jX
jRBAUPvnizwyBuqbBposQsL5WVzVrhdaikjxWeH6003R3v7bioI6YZw5b7wj
APMMG/QB7W/hvTj7+oqUdO4UcYFetF0n9/fHcwfAh4q89TPV0Y44Cz5Z7gJN
e8HRkuzkxcoCq2ia82d92r12/u7hftF3kCL9ZlO+jnbXjRADc83LF16OasTV
ikfrdU/y9LAJHFkAY6Ku0V5kmesDWuNN7K3fhhiBTLYCYVuogjzoZCQrA1Da
CjCyJ6pfE0wsxAmvnjTA62ZMWvC167kzdEN20F9cI/BAoaVJQKJ8Djyh3QVt
s0wMJtdxbzSQYfB/Ti1o/s2RL9DXSFM8adw+mgG00TxPy4D2p0AWXi6Ow54h
Y4N2FKXWtoLY2jqDOJKsc+Bj/XXoZY18OaNEhXHNKdVuyl7nzSJs3fbQPXXh
ROWsgjgOMIw4zQ4MW7Y8URh+nwdehIXfWBxXETxqGGPechlm5jdpWxM9MThy
MrfwVodI688MAwGecRDCNgM31kCxO4+qHijmr3gk6b+bCtbN13pGOHimSNG8
dFU1316UrqdzCFMmf6KBjYcRM98wmEeythHP+nlVwD5cVhC9UjxKCJa5g4yx
MUg4ineIQV0sY0Rt2mUHrb9oniUwn4Usilt9omRiRuj8pY06M9UA4F3ZRodC
EOPfih/Sqm0oEcwlpUDB6Me7GE7RGmAM1pbGzAbVIL1K8rPW5HYKi0s1DDs9
RgkNJbXxqYCZAnn/+ghI6k+4uLHdMsZKUh4hHL3l6ul3srwkXnea5DQjyB0x
6DH6u7x42psEQz9hb06NOYzBFcOXmaohkV7pt0Yb7v2VS2vaO/zx8/rg7FZM
W1hMWbktEPFEtyleYlddgyapQmHl7fn3PVaQQtvgf766yXeWBFvVsCTZH/+5
ANdxZa1jMGxqVDyNlvoK4Zlyuv0EfNLVip8EX9tkZgC9lvpc8yUSvdj+M91x
3rdUm8sCOuHlMF1Cio9I0im1eYA5TFV5G6DJcClp6smHWoiHSSbXuBhV6OCW
qQPFV/D0McHuKH1i2kxEmaQc3bGhKYXRAelmSer46UOAo8+BawO0KOOB0Xjc
wAENbfyuHQNBsqu5TQID5BNytWHyhgzLHH3qKePd3XIy+B5SNlbWPqq88nOJ
+MKjiq+mxaw/hNwUKk6sYoQz89xBdEmW3ZP0A0XCiOzgZGxh+DPDbUVNwyos
RvZGJMs5/h0Y8SETaA3FIIfgxPz3poY+O4wEySqeelQpTET7T20CIBUuzYf9
Rurr01DGnRRRh7U4Q8HfpR49C5BJah09hyD55eXIm8vAodNG+yEG5cIOdF3H
4eg8CdaYB9x6fOJxfX7Zivwo7Q0Xa+JSgSdE5hvG0dixNZQCXFS6ydZcyGaF
749YXxJPdki5rDBWSWqVOAb8ldK2TY981fmK3bwB87YneUXLA/2pQLNCcQIP
T8MTSY0ZZFUFWLsR9Z7Liqvon3jjAN5MeXO13oHCYrBTc83FtHV5YyRb5n0s
HysunYLd8fQXlOy/Z21PzXLPo7Wbs8rhg4ALldDfsJrzk0BWbhon9KI8mQSY
fXO7be0xmiRVinvKRroUrLFA6Ahej1moe9H5eqACMuuFWK6Qimzb7c3wxb3y
O6z/qfnuaC/7GFS2vnkERbBVD7VgcpJcziturkqDWqpbWc7h0DmsHN+8xf/R
gZRX4OUxs/5j1uBX569QeaqgO5U4ghVaAqZqtGZfD6iJVl3WUJXjiNBrgB+8
4XKxEN2c8Jq0fhSDSJyqrjKGOxadWBLVQ/KNnI7gY0C0Onbvz+dYOMrScV1d
H9bGLO87UJELjaZQ6m3PTKe5jFP2bjd+hHo+wxqucpOqjnNxkvkmDd9nWyxW
nWNaX3iWEYzJnelXNuE3Rj/HlLvlRwXH+Yp89zH0eyzBRVhraQKchWOmIKRb
1r7ySecvCfI2oelIJLykoXbycvpZBf4WP713iMi4UGkP8v4yXriOIU8W5orZ
ydjnhqNOomPyUtvwB7/Mq8EMoNH1Tgwtde9Nb4Z+CKGFx1ZrsfcD8asLMiWQ
YWb7v7ntxPsowwqnadEb38hBA55ZXXfg4971W6FLPkj5p0zLtftlw0wjttJo
olRPL91I01GyDtYL/AMuTXXAilXU6kJPuTVJpNnoy0gwSG0Sb36FyARfNW++
YqXZ1FvuGCSJeFVJzOAr4+qlQ3dEns7OtUCHXaOop51dQXH55qEQyNsFV1kQ
PNUtoU/lXcli3C0VlioZl2DEOnGolKUknBHAIjMuuAMnDMZHhrhLVD6ruoOQ
ysH17WSpM2VrOhAG01ip6rtJL+AIv9ST3Ut2E0aywpUvs2APQAxfDjLp16JN
08ujTyzsAkJ1Fxs3e0fwFE20JTqFhKoRji8oXpj5AOo1aPGzlfGkUi2arF7S
kk+evxL5jUBFCO3X4X9uzBFtzjQduALiDhhWEGeJK3+S9iF7Aerwp6Amt/X2
kYTJp5IJvfGjopjjUhMXoGmKA8gyjehc4ddsHMlTT+IHT1Q7qjULKOeUQ5Tm
Co6s+mV9Pt1V6+rRovmtbe9OLcWoiExAde/W+bWFaUTDIbUDcnBwYwwprKAw
Uz8u62eZH7ouQFjQuXsmA1qzLIBCA2ZfMeMAYXbQK+dtVuJVI4rzAum8YEV7
/qmWajfqNuTE/F4nlPEnl57CjkLIb5JF6E8BRVf8Z5/ljwI2pNPS9tlI89L1
KfRS7lL5aPS2hB34Uq9yB3UTGhbP4gnTpfpNs9w7ZJXbpcjfaiYTl94uyCUb
3L4S2nWbqzBftI+VHkP+lHO6PWqNYO7Jt4Oo2tAbBQpWz2VPKJRSv7729/BH
hxRu25kO1Uw9scW4uX8iUI9NEpHv4XL/NNoSSYBP62qiheKmxrls6/PP3+uG
zzcsuFF+RZYvjw7DGAa8Ldf0GRTKhRLisaP3ibTXwsoplqz0V0fuOvrvK8sy
uhgcpMS7aJPvAgRosHrPvyadHKZ1fZLfr8vuh8LC5x9yfGXE4TlGvkWyhl/T
bF1DY+hO4EF0V9JjnxzJupjxs5XW92jEjbCbYbqmGdCUOf6jBKUR1tg/Rjfg
a+s6lC4Prtprbl0O17rKqa38RV8/LSBcwbNdbEeIuoQX2U8Qv9ItPeondUwv
Uv+jwTwt27EYcBTjkdqp+JhyNTQu7mW6oDM7CRGvM+tuSBDLk0urUwY1WkxI
PnK0+IqsmoOiiv7SkGu05HRWuawEV+lYvH5rRUR/47vCFtAaRTAI2Jof8O8q
UshLbrB/K56ND13gHh/KOLp8gBJz7CLkdHh/AAWzomZtUUUukytdKaNFhkYg
cHto3Pgztk3zpB2KIgIPq31QE7Mah4+bB11e1Gpil2wGir7hMTP0nJZI3FHO
TFleETDk95H/jQYX3ss9lhb8/9zl+BFnJQt2lLVoaczhtjL0Ngp8F2KLBLIz
K2sONiY5WcAtxj3ADbT8t5auyK9oTrOGOXtx10ayseC9lQzJSGSAZopzJugc
YNCL5Sel31Nnzn8rXJyhJ3j+vSjpgG+9CpxpOe02QiK+VsF1GtFvlw7qJ5hg
IZZuUwMRhTSUptu8kJLxz/QokJmHmn+XjpZfgwfRF37E/sJo7Jk8gpcmkPX3
VKZOWi7kqQ8k/pQPibQvNKMa4PLA5dFesZ7kInUJYGTVGV0wi4l/Oeq0a7xR
naM9VxFlUag0DJk0g1fMsF/DtXPf/XsCAzyZpdBdU+lKW1h1gTev7OGGvgzQ
JuP5PiHgih7fsbY6bn18K4W1ci+NsPQ2H+fThUBEzhn3rl+ayR9fps78TZ3L
D3zjkRLzo7kXLBPibQ0Lu1c8BF+QF1P2baFUc7B86cq9siWh6uIRpd/tsIDv
dNNQio/kMxV6WmCsYd2NpDd9AY8H0iFeHdLaFvjCyxTV9cRFzScpQvmR+tof
27b8T1NmgNinQvddK2LNhjQFvZGF5znkFn5+wH1F2tTI9vwhSojHSvrSHzJH
tnhNp4MkwMuu8raOBHW3H/L2itH4SyvGHkKTYOc+rTDLMCgVUa0VutQodGdp
OSm80IzIHjJETXMFoseMUxviANWY31I7oCVXFTCpe4UAfjcrYhOFJwlrlQp8
5wmKf5Scp+TYK7xwpnDDaoQZ3zq0YyBUDuKy3GXPtpp53EJFMjNrOdUn6j9r
jDhKcxgBMe5EOqa7lf5N0KIFwdYgOSzsujmgsQUIq5901zyygalWcP23ibzJ
YIz7b7QwJZXSzp+dIRkAqMWF0G7HRjDFt8jICFjya8Kv39skxFAhTas9KIvX
9HnleM16jnxIgDJ7DH9/ibnRDJSgOlqAvcgWEUxVkFhcs7lMHOHyPnjMz7HO
l7Lyd0/NZbGETtmqE2CmkhvhlutrTAFvrp2Oj2AQkkgScjHsij53Flgookdz
qeV6wBQAOWomWwnCyNy7rNKPxwZgKO17n4lZZPpQQwkwcY2gVj2A/wVIkPa0
x/+s1lZ2YMDdBW1fuAA/XasXaCSlOcc3o9bEnsot+PeIHZfCJmR8CpxQUDLy
TpFud16Cq82pO1MIAw/uwhAKY9a8ziw/R2tv+rqnvi3LchusgLPRHpy7sJbi
qiswNMB1tmN286To97/7D7ARS1pIMCw65+eDjFF/KeboOAnvCbqARQL9tvKQ
BxvrT6yDT0faN1+uV/wN/2DEX1pyq8lmiqoeTPgKmI2BZt87n/0pGOkKz6OO
Jx6UxlqW3hNG7wlocqr9/YRZvwyE9+/kApk1t3Qx+0TUAwF2Cd2c+9+gVpgy
/bqaMCPzbpYi+AaSyTf+WfGG2vQyNqQI4KsU5ttTaSP9dEHGz0UCOm3mibJE
Ot0pOsv33qWAb0asmXl2GTjCnnGKH0fHTu6LmS/iO1pzR+q7eYWVTbaqlgY6
i3ZaGnwN4832QTfS8WrS0zNbRhJO7pa0wgZzsI3S+OymEDu58o3FAfvrDPcV
6bz9FUuf+VtWBr1HTT+8L+Hp6aPGOSeoBOrageJVGjJeYgPY6NWhtgejfxs8
2RTr6MVBofAp/VXpLMxvSz/ldlCm/sMSLWmfg1L4bZkGNwgjNSy1FDgKR1K5
YzqAb91b2rz14VDvi9YZ1FpRWjQl4HPaqjWlMWNSWwNvJUZ4rdTVgFu3Xqor
F9iN4WMmXArsMzWgwhWoXzklWHagnKi5nrFgsHA9850M48WlByASWtq3k0EJ
/cekIGeu2neJAlx5hP94KdPghg2zfJrC1a3rT3qm0KqAdzFd9DrjXWp9lo52
0KKIy1sPAgnNPNg8h837nbwHWXK6djILWEbYWsrbxTUHxOXoauopP7tHEgUG
JHktgEoHgKn/0r6ceQZIhLkm5zoutQwka2LcLtH5nazWf2UC+mW3ehQUK30i
hkMNjDOJNakzNn6G9eoYTnL+YgwzOKtxXEHpED34GbkO1oaZ0faRO71rMwSw
Tyylh67AkAG/7n7r0wL87M5O+zP6FqSmY/ftskxB2PVIm27/a9jWkK5DdGkh
rUHu3u5ExYBo8AHalVKgaefLGhA7d3ejw2DDOpTvf3QY7frUo2XKyRLo/V/K
R8wXeiXJZL777di2bdSULPOaV12GB2hnWNjBlofncACsgEi/DUPsFhdhiX3H
SYXdIsiDhHIMv00m4vJhG3r6c4OskCcAZSHUwwQQIebmKEOpj5vEPmZApb4u
/WFZgYOcMb7tSU410m1FyHbmEOryLpDwCdy0xPLb/I5lEOWYJxkuOXPfEq+F
rUFD+BM7ibRlGz5x/su4o2qUp6clJDak2bmaYHg4gjYJSey5JKNDCZsKnIsu
o53MIq09RkptIVjeMQ/XPcF6YR6o4t7iUyOvTWthig2s/es59huMJflPpV+1
tAbr157rWFdM4FG+g3cLFYs8WplyJlwIdE/b+xhHAb5GRetYb4aaz1I9glXA
zH6nRIRJov2uInd4MJ5ls+Pw2Id5D2o1T0iJp+8Lt2bhHbTVlJk6pS6ToNLq
AxpAWIIUGIc2r4RltV5R/i/tcoyPf5yYDizr+idsiV0arokPsByH3PD1P6SG
EODU0GL9c4RpAOIKN6z7h1nuF2UranXIFYTLKUWHGa/BerPxZa5p0mn16/vz
BVbMrw5DmNEpaEWyx0fISaOM1DN+ZrDyI5gGsIxskmhEin9eeBhDjWLw6XMT
gXBH8Fz1FgltWZ3pDAKR3iJr+uez1rIVryw2VsJNr/A4vu1jQDNL2X2+w8lj
XiReMOj3V420xZGojRgEq1oxzO7D+iEk7TjoN5eo5KQGwhWx/Ob1Nzy2pcbg
ls9LI5+WwffVPofDyD6KNvKOKrLCo01sOYeJbT8nkXffuB1mPn05XUy4zNyf
ZPPLRb3xlMAMUCIPPxiFsidl6QWRvRsnhff/03R9mjZUwEc0Kdi7/A3QsE24
PhCEseVJmyHGYomKTSE+FpJGmHiXBr3ueCiVg/y0F67KVGIzOla4ULielxg5
n8f+oW7rgIU0LU12B2PvNTdcjm3CWRN7fcPElutC6HiWyMdSPrwP9YM1pIuZ
HN41Fmqg9YI8Fs9lGLSmh+OcZ0RQ5yQCoVFfHgP7BHKeChztJEdo0YlFgFob
M4e0XCFLhYo8z5GQTH/vYhbPfXN3WdwsIZF6BEkIDdDM8gSmu710pc/v7Fzk
Mh/DgbSvho3fHPOmd1EHQUI1DoFiiSnTBKAj8UrTG8Zldvd2GA1AKs0eLkEK
KQRMK4yIVJ7cfwPgXgLobHoCXXilhmE0XI0PS2sekhiauC2vlZZUztMc2LY5
BrK80O+2L4pZHJaTtsCmJTCE8ldsOa0HvobeNGz4ak08u/FKTl1FwxEsc4ut
YQTVxx6Q92zK8alpy8SlTFeW5jL8PqrKY9hl7bX7HEaROzxZKf3xUcfzkd7X
L4QXHQiC9C4dkIdlwekKmmSiJSYTy9t6uvoWSdQv1Yj83+U2/gkQd9oTIgSc
vU+AZKuXzwdEe+6pMUN45Q+P6uy6u4h9vvW0fowO9x2b9GX3eNneDml9jzRx
nosfAj/EjFlUDwpF50nwGnvr8DtV9+58uqP2cTxQfP0G2MAKcvjhfhw24W6g
9L+o5pEvg8RDX4YOpA8I8FEHNpWrKl96NFAETOREcELX70LMg1HMShZEvxbg
rysMxfxCrpBJ8Anoa1Dq57Fl1axVLvf3tLQsaHMsWIexf9x76BYykDs/znAl
PSKFZ8QSJaOY4lmA2H0rlNXgmxTPdQSYk7DpOW+wzRvWngcWYE/iPb+tge5b
Sby9+8qOuElYcN9ECmdDeukP5QMR23p7jI2NU/6BUik3ttM8rh0ouvvrRLAf
ovtkiWuFqBvndozw0Yr3df/M25sNK506K+5HclmnS8S6Naft9lUYSWgz00JQ
P+WXEGIuPxq/ZwFwCmoFtuj0NO6jRO2XUEzRhwUTX+fMpWTZOAN/+k9Fyzbk
F6WDWL7DG41KDJrkIJ70lgSZ82cnPpDAev/Rypo4JueuK/8cWDZRRoB5+sHh
uV9KhZP+GXm/BvKQYmGG3UpwsIhWxyuIi/H05aRTPtmqIba83bAaGXI7iKF4
NyOPhzRwmdbXB3dF/U90TbdUpxZzX337G2RZdQMFgNvqhpF/HkeR+8CWOSEy
WaeR+PdqXOviCFcbxdgBAJ5lBbR4bEs/KjAnpdPmicg12NZHxOL+hckuygra
4DBVWxH3tVnbyKba5bItJn+de+kGUa9T41m7Ts62y6UIHW0xCbHVVaW5cy4T
MdpM3yoBhZNndUPwDKWJynOR0zUYuIo8nBuk2uGvRUbO6XPvFgeoO+XKHBy8
KlWj7hiE/Tg5yRy0Iwhzyt1Q/wp0NE9xJYLGepLd1QwfziRbYgDr2DLKyY+I
Rx5uKBB9RUy2CwoC3HYu72t7Ri+RNr3pNgbHSDXxt/cXxgwzPzEvxB0AbopW
ZMmpogetFuzTCYFC4TFxA0xmp8BnztzizqQBB/ipPPiJ10IcxkTAYbTsMDGO
Qhj39W/n2eJiDZLxCtAqIKj08L+f+x4wZNOeonjbe/wETMOhSBrrDP/Q2MYE
L82UdIYHbHg5DpzSvPMUkZneFttjg6OUr5j2p0+hd9quCy3J4QPsjbBz6kE+
AfeM7+oVTiijH25ZJ766ZClkO30naiXdH7DiV6p9/A4Nl2wppLkJrWxxASjp
C1gQA8Y9ETF5vyNzuF1XGNx10FE3lDSotv8tR3KJbaLwLL9zB/MRRheF5sTw
1EkqDRoIQe0P9azyLY13fRjaVRouOi1p+3I0oUJCO21I177yjpy1qjOhFmAK
MHALnEPCf9g7IgA8iJYz0z0to9+wMnDHs0vBPDJiEnQvVS+Q1hDW2jZVsSHt
DW5e5xtiwC4NJMVeOMUfZ+HcjbPjpXTzZDCSUyDJVyHavLSxF3hv1Eh25JHW
iPH/f5jQ7k0RvlC4QzplYkk0hCZFaxeAlpkY+3urOr+xQR8HAmGo58AJLbva
i1uc0GqglOj1U4D59kO5W9Qh9j5A69R0oR1lu4/b+lLFIyiJ8CkYCyCz8qA3
il8pb5aqbc83xjrh60un5z7/YYt+j1W2D1mjtO/j/LLYVA1pvWHnhMedNeG4
bXp+KqOud84LINCsbmKLA84VmIsRhHbpksX3V16ApJHCY2Mn9VBe9daxnrP+
o/i4eVzx58I2wuwr2lwnsFRg6MCQAy0a2iCzL60iV75lC8X4kuFG8XxKRDsN
pFTj7zo93vgtmCwD349JzKU3SNe8B7L/NvxyZ/k/zukibDNmDayHczNb8eyB
bR9uhiWsoRXJiqsqB22RuHJl0m0L25kbWxeALTBUTuJoJeD7GO9GHt8aHfg1
s0paBfkZ+2wzkqAqM9yg7vf2Ayyqqpx/rrSzV1/eu3lulT95AxrRXUtKF32p
M9/cVzBWAyW4wuTPdjxMhhgFs7v4YGW8hy5kJqwEWrMRpM4k4mkRKEqRrdIe
Sqtn9qmbiJrnHnshHEH6nzE3BrykShqx3VZyME4T/Gi8JQxodbrGGPBujAbY
Nc8LuNBgMAemnteA9mxVmUYyLyjJ9fw151YuTybMCU/V/lYaz7tieI3V5cSC
/w6U4TJfnx3R162z674ASWeMmzoF1mzl9tRpzIF6MyL5XIOxtIRjUpHAMhSm
vmFVlvHvQTkooDdlsuB3PefzWNpU9Gnq7abiFrpDOoDxGuKDNEXG2xPl3zEC
zAM0JTLAxuvMc9IAUcVBev9xE5tcUEJl1qBn+goxhkgOJ+u6L1pM0xjkvYIN
L6PlpIpEm1lbni03ki4Guej2MPdh3f/XTZnXut8c6jr1FrBGAydVGXKv5OiY
BOYKYodiq+aNXvoGhaFUxzay030pnPVpcEN5OEdXzEk+WgOp2+lT+qUQdiGw
D3s8hgkLIJR1M/8yEPbCLEiZfrknKPX+jvkJoc+MnhITO5J/Ks26BS/mMwy9
UtrHS/MACYuD2YQ3GlBuaQC+Qjdq1hMUoUJHoSssvtWhkCCmigsgIvHwGaHQ
u/rwqedp1FWFZI9lHoeL2Ct8ZRrV9Cl57n1HrgQZFkej2MMZiujpcntWcAIB
dwUtEDdvDfknvCMFUDM8Q7d1I+aIuAcmwV/KqvjXiw4IpP7mFwusdaYXWTuB
W+NiJ0uV6sZYKMsP0sXCtR1wTFEQRaBIJHqWAAGG5Kp+jZBoWzrNuQl2Ucqh
Cf9oE2FOnuSk6/zx1hoJn4PsljUCmBaWNk7cdebUEQEM9l7XkUFMBWr4wpya
bcUaux4vQ/MiWlVxawNmTDjWsIK7202ugUFSPkNPlBcSTDXXUqqhfxA13a7u
21bpNawRUuOk7kYfG+PA34OXDmKVbTDr8VSmSu41UXQmgBBuWVPMWoU1ji4/
KsopMd2sGrOwRZiOFY37u0+7tcSC/arbY6YioCVKSVX2EYeZ4xXmRk6dSYkx
S+karI4oZxnMRJvGNAdqX2sdLeGgBEpxXu+UYpqmVbqbALCrOa6o6yBMMaaV
A7IAgS1Ptc3jFFNDReFTB27ZiAtZt2D0FKlh8dC+XH/FW/7tW9Dv8qMaSkNj
55G+TCxik22okgWG48RAw/DfaSfGuUq7btB/KQVl0uLTmhB6bfHC3PQ1Lqe+
5FTENOD9uHUdORr6+Zj9l/y+fRFskVgtH3P3j0npVX6FlFA0eNRMFAVh6GMz
w9d94eKwD4gF3I4P7b1GwUkZtY+X0ZQxMo2UM6XVU3MEojPiTwaQyQHAz7YR
Ng3WiqvNbVuEvsrGh10anhmzb638GoUvoU052Dh02Ek+FBBjxAWf2c3ZzcME
LTKMmO0udWjDopTeI7QSJ+TkZyEdGIjBj1S3oq4o8hEPG4fC3bkmLzdCcR5o
g+yGs7kt7PN98mNkVSdOiUhBbrpmyQhHUsFGR+f4VeppwccBQBT08wHTr3NM
HH+K3G4fDMbS/FyGMo2n69n24pyvwMjvYdxWMuTAEZrdZkU/XV4xxYo8Wdiy
Gxnl6ebbKvfZV6susjqwVDxwv312HgNsG0xsZYepDct1Cnas5ECzwiMYm8LV
bME63/whnt9Qt/8+Kei9HjNejKh4KCkrm8VzzcWDyS0JA1sSu/b8syFRg8t1
C8kmo9wz7Q+A0ly8fmhJMqFO3BUFHm/d99GPB3RgFIQAs2toGveHJTzKeyuu
AKChQqn6Hkj4q+wQ9owVGRVEvnqPOrx9RmxBtMmjtRRiPLuE4sdPISLRZPKd
SiPOgEItIsz8kxrDKQg59WV6xkAG3tbLo0ylntRpRhkyPqBtaRCqAD30VPRo
IWFnN6tBfBV8IQ1F4MrPD6HZ3MyEFhsK+K0cHdX/

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "B40jvh7ud/ahkCWXo8CJP0S9JYnc5+J2pwOdONjrEnmjRzb1YpxBEP/gM90XdEQFf8e+9j+GJABVN1VA/EUgHmy986oXHU6n9uJJjaeBsR8h22iSaiy//95eH4kKFakRZgkZDqWp0dX7AUTwRg4vZKk0rom9cx0xsiuc1Ki6fTzxDmmuuNW+yyxk/luKJogixDl7f05H1PhFx3JTfD9y6cRFGovJ+RtyYHOBbLpk0wjvZo+edItGRXVkEGWRw73J202qK//Yf5cjq286dpMU28e1wVLm3cs1bhbUqY1L2da9yOdeFOuBWw8l2rqEgu3kTDAo8QW0PlRCbq/j1ubbHPakCptdeYXsZZ9yWwMeAiGCvl8Cq2czRdCzUdT/Xorsp4kUDIXc1bNuoKglYsGiZN3ziIiDjJnjAsVnuiYFVQ21VUwIMf94C8USBmWhRzRI28g2h31Remjkp7k7QBe7+O1L+ENVIJ4yuZw1Vml7mc63Kf8/oH5jlPHcqf7nylAMBf4EcN80jVTfU48NB6BZcIwVJfJu9xk8qKDu3NtgmSSDHQjy+qhL0pO0bt1j4Tv01Vs7/QsFrlGz4/tmagm7eU9a6JgTAt24OuXFY8r1vTz/cBcb2SmGhSvTthvCCognktOpifdswfzgqgRW1Gafnb6IwNImZaiJrMljWjt0PPYX0pe8zNujW0v7G92r0cqFsWUR8r06YQyu9tvaD7hNZb0j0dNQyEyQfqOchpk7wSxFyKwc93zOeQjbAtL1Eubbb/PQRWjWmkm0HqErH2+7jfZpIFhXEZt9SZmkn7GiGZO8h/eyZT226Abi1btTaXkvr8SC875R9UFK/VRzUvIcfrgouFcOjVsVpHSCihb0fPtmjw5aGmROXCMnIiG5axcE/SKxMmAYqI3AKMpBwLr3q+W3yorhEsgEI5gh096b/XQLE6jcSnIjt7ecF0zuQ3HRMCje7Kh0zd8aOH1oOMYo7+kfTHfTGrbH5wWYvLiz8f8SCWriJSOSmvhZ7mdYh+nd"
`endif