// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
0RqbYsFgE0wp4WjNa63WCV5Jssjf+3SWZyhMTZbWDOxlyDf40+uKomyBhY5S
dwUqtBu/UPulL2JnSwwucUSQM1WHL9f7mSdMoxedY5VcwVi0+f/TdSbkprAH
/Qrok2ytTuM9Jnwtz+hZlJyddguDtUlHCV+rcN4EicXIOi0dFxZtqVQXVjgM
qMGLlCJh5lIFQg9d8PZ5+Zkh7lPxhdplQFeC/aMMUTSOIsj3SPoY9Ywk9ffB
jrXqkLDXX35V6tRrDQr+LSW1R3TtUVVffMKzWGCALXn1YRA1eyi3IyhePqzq
pbpK+XHRVawqeZtdqXhycCNJlQj9KJomenyxfnV1UQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HhLMuuVkLx7icdTUnzJEZcAi7sNftL9JBMY55KlQvBK972pYwuaq84tRadlS
CVid2kZHzUdZZ0MhseUligpp6IKbapyexVgaOEDZ68KAsRNnppZIQFMnglZr
7sh9UuhnFvTuvVGKVTHUDfd2ObWV2ANu5o4cF272m4gkGzxbJOBmYHzqD2Yy
iYDTTGqkOLfs605JvXYhhmy2kwe7FcOr5hb+hs0IH4Amr5fDEgF6sVAbr1lj
AfKM11bthSjRqA4M/faU5NGnuGkVx3qg+iawHTLZUnm+nVpNppOzt6xS29vv
JuJ8qAUu7/wB0l2xOWhWGf7ya7qHnZmTEC7dIs/xcQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
L6wetHnN4Gy0SqDaby4J97uu+9w4wYSNs+IjckdLCnnhPB/5AsFo5yH94gGu
U+RKWR0DJhjX0c+KvHvzkgUCT1RrhGaQcR11SA6y63bgPBoHzbkCML8CLEmi
3DynD9LgRq6DCrfqpjfUb8Zu1V7rCvIv+kEVQqBQbwB095f2UDCm3lnawKsz
6vQhP/zOnKlfdNI6HjPrGWEq68yownzEGIna5PBqvfxWwyVxQljYTDhYjtwt
UcqYHjd0YbDk1FVf/j+KpiB8cp8UyQCQaB8scdwkMoYwaDkgnDRCLP5gZrkF
yH3NkRtxMO4zsogVR+KcfLJH/9qiSVsbGb+t4TGQog==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IAYJAGtusCJFc5E195Ax7hFFCdvAlEGZGQOtSNo9LacCBLMFYqMVdI3iftqD
jCm6mgz1+u/SlHugFZTd0TY/ESkYVm4yeG6uP+jzlK9MGESQlm/Xcv3OONjs
w9q5178iX4OMgWwAGWpEeLMHxtYrcEOIQsy+lk75kc2uHdFRJ8vfAXODC9W6
2A9A2qB9ajooebOoOoxLHqGT9D0Z59q0Vncw3GNTas7OKip0iWAEMN4g5DNQ
QDEXIluuQ1ZYLfCxv73TQeOl9INSSivaAOO9gI4VnKJaDzWY3ZHJuShYLWot
PHgLfPoVQKks/Q75yCjGpmBbLVtWJazb5+ShUJQiiw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DVwTd+Nj7ivat8ml81eYCtpPhu24KoaAn1c48CZB1ijkj9rYPCYeh9ht6J2/
OWqKWVDhQoz19knOwEW754cpCPv9alVZ/SPxs0IdReIfu3oeVFg9FKBD/CJO
ezaHYyznTYtafLWyggamzNhFoRsaQ+AeboF2MQqUGmKdLOMCzhM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
rmezvlQzrJpajQNxEmZ/ykx6vBHI2a4Vho1bpxBQVEIXAH7AuHU6wo962+cu
C0kuGPCzmwnsZuI70FFPQ2I8u9dQ8a6erP3Q8AhA4ZUt9WEELkJhVV+8H6cS
gR3ryl7YLlnPnMB3yKmsx/MB0w3dVUXLIAZHbiXGYT2p+nkyuWd26kWj/YDP
FtJZyfATfN5ZUhemaSXKRxvkQmlr3meD3ks220zPfnJzaXuuLnx+bD+b7LCr
xh5ZnW/Qx9aBEPGC75/YYBXUIeqOmDYiLj1aABBdjPEiBV1+8Z3yBH+g4b19
Ti1HVZTpMPq84wtQZktWEdaHL9TIahtKxTz7E++M1iBztnaJ/WEGTEqfemoS
T+xMeI1p6cV4x1oOdJntf1KNniTHz8rNr4FYiP27cSjQZLiAczfZ7DfOCEcc
3LfrQ7J7cfY/TJiLAid7ZfArYQUeY+73Oyw/Wd5BpGVMZg1NREOV4HUIWZ5S
KqgsJ++vCKFHPTrELgbhOl5RW43Fp1Gz


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Km/akenAv//4zmJ0vQqkIUxlJxxBk7hhGM9rXVaQ+vkDqs6w1L7CdiaUZn28
eCjbFMYcUpmI+y4pVr1xKXSxejRO1vNs/Ef86c+FLK6dZeK2fuwIvBD56nNI
PobHaxaSnb4iLBwL+wlpKHRbZ8symkM8DrxXfyaD3/m/dn/qPRs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bV31mDglpqXLVZvt3eQ5+UY0KFfCUsdRQppY427KcB6RAApck9MrkPmgU59T
5QE8JCUz/EhXg/WtIbYkSFkorL+I7bf0oZuLbB18R5DvNPNxMb28nRAPo8iW
RSP9rx2eb3Cj6+ypBaw2m62sIpIKAuQtjcsAhJ1EFp9Gtq7P/Dc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1376)
`pragma protect data_block
faWB/TkrLO7UgeLBfP6ICswip8I8QRzZU/ipjShfz9+/UnGjsGwylu9Pz9kr
5UB2GoTKK+/kdhuDcn/KtJ9zfo0Pozv9ttzWV9eOXjrDmFiZ/P3MyNfhe/1L
/hA99zjoy7AliGnmPWulUlnQXA+yAkV2feFZJ9CvtSAgLOyvuZOLOJQ3EY41
Ccj6e/BSLMNHi1RYxGdpfPPjTNdOI/ikc6P/fLmMuCmoTTxZ7H1C1uhElvx5
yUHTCyyxrsFIFq50gXFmDueCtFXJAL6gpUTgjdZMnfZb7ljWzHqzXLglTiMV
opWG1vGtRgCDQHuyRfjl3zIy5mje63OoGfPYuFgnmD0eEai8Q0Z9Ox3ehplA
f/1akvYHdNDOq4LNC3/4f81DSWieYYwBfha5GIIJm4u2xJJT7Pa2B2la0jzz
9nVmlgsqksFDzZaV/mZFCIcIxU4l0OuYeZuqK30jFiElOHONp7Ogftmfr1Im
DaGzXc+U88xv/VBK4T3839krZs+3NyzQ3Iec7Tte1JBAfioRWzmM7H2mpSVT
ouZpAqSw0P3Sj7BQij0nXImACVBUtTKQ4hnUjuFsh2fEcpwitYyzlnUITqG9
rlCpwOOPyQJqsbifJiaCGONU/w93ODqvEPAWOCIbJ1W5L2kSBgIkiAsLm6pO
MYgQwX/a+w26LYxZqssrytX0O/5wZ3wYvuI40FRGKVgXPrykqaIXobeBxsbk
tK/L1oqLfP3c+0GXq7/55cBiKcm2KZ85GLS4AJ6t0FABZHyMIJAKQgXtlRSL
8geDzRBGh5hHL68NZ+ix5zm6PknEJlhisg42gl/45Xon/DrlzX719cE6pe59
UYCCxjMY9QyTI4o1UNmO7KMy3RpAvA3FbWbkF1U+acsjltA57lCjec9yALFi
cyBDxkgvJ3o9F5v+QOXPsheV9tyBE2SexfbMk39GL/9kMkUmvdZ7kVkRpW1W
H84vjzrM4S2XWvL/ZwpN71qiZKBSoMiJKUpACW7meucXRPpCfVeHz4Zha8Z6
Vnk4M3v9oGt+48jqU+tbijN9hvSarg4yxwABfWti5aH4SMMkn2XeqDGCSZnj
ymYeJTD4YYx4C6zkq4nl/DagBnOqPl4jbo/rxGrmTJQ/Cza2NXDYmj4bMgE+
Ouo7krWVdNIL+1uvCab7aseJ2NxwhazmtecLVCPpsZx9hvOqTdzgPPoxYZOI
cwTuPtuCyRiQwVG5l/VmT+8k325rd5X6B0HQp14PQKxoinVna5+QCFxtHij9
dkxgZuPLDIr3jEfiBjJKq5T2vGjKg5yunGr28Mr6zG8y5HWOy7QoFIIbNuWE
yU6E5A2M7Y2+Z797X1n1u8/a+MkkguMENoaqXnNvq8gRsaJKeN7TILSyAd4P
XuJ1xE5CJ35QEXP9jLXfAmKZ5JUpoTmHxnECfwB1d0jB2JZ/0T8OloXbCW2O
KPpeyg87Tkv88NOfN6HNNH/hmtDdT9aeV1gCH0J3ld4BQ9gFun8KCBupnfmP
tZome8nJ7H2hQIjh5n+yxotEItBI2fxyyOQxE23u++G/IjhBv9sdT0PRFV/T
6pNJU4/tEsSV0gdDBYl3ErtBynmhV3/m14YhHXkiQ2sRKnffGJuRAKZuZ2fR
4Ku7J+itMnnWRZu5Bw9Tn4Sf8zb5Bmb/p3xTTAbhi/9/cu/7nqZj+JMg03WJ
YXD+1v7zrTDYPjEaKo4kOZnilPwKI0L5KvLuyY5LIdTnekdK2l3wD9V5MFIZ
4jz6DC/g87/Qn+QxW7Jsuk/8MuNcb2Kt54URXX8XtHHhJRkeNBMfvDAx9UJu
5ujzNjR+WWSDAH54osmb351fDmkRHdJs090=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fidd1oyAhusLLJ6+7Y4fW+UxvqV+8TisWbzB76p8J7jCbedVkgTXiBKrUzNVBIRDckfBwS/gk4qyrpXnk44TsazVN20DO3TdF1x8MmH2pGcTjxrJqgYV/z3UJLaYPiY1WrKUNRPOAuHkyYvfI5GoAsKohhmpB04sGLV6+cGIymx/RXK+eIUgAROf9S5AOXsk1U/Lqv4gR7i2yfj3c/IhJWMX+Ld3X1LJ1lp+Ly9OQozJ4p7qcSpIspKO6j/f2bf18vLe1BfyQ09Jde89do/xhW/KwujLwEhQrKWgvlSQsHu68NeA22zcLBqTE1aL7Z+Egs6Xw7dblZGH4SZ+ErK3eL4ositygoURCj4V+A5e3xLIC8s3izRjPmr0vJyk7XuUBXqDDHIAKYkB9Sd1ckl05uoL/p0VqmxCCLgwO34Rv+6DUywx8lJdfh3geHmhLaGSfQwE3KxS+Z7Q/d0UhH3jybb+e3DwwrjyruH8a4rzYJzzUIBCpR5w79M+UVSkuuMPYOQNM3MJKvQpRlH5ZncCnPy9mfod43mi+0Xso2ZFkab6PwuYOufWirajV4wRJ6f94GJ+PX0vMRsmMILuHUEvcph3AsqhGPEa81AJwm8igU99NIQj169TX5tH1PkPqcSJxFm6sQYkpOboJwGtmhkMDWeQ4EiIahEdPPyEWeT9vHnlTsqV7F/CN0bdRln1crQyuAkjwBHDJ5gwIUU6i0/l8UYK64x+6Qj6EgC9XXpQJ2ooAOrRDwgdj287ujeW+qgXxW8YYJiTnW78pPDlPb8O87vTX7DxQfd0IryjjAR2dj4sYaGYa/f5WGXjsn+iJw9983epWGcWB8BbW9GhqGt6ciVeI4Kk0iPbzq+E0gWt2PyLM3rPdQh2IW5RgGBFFH8Rq0JRgFmZ2gUiI8AciLNTKo2od4QElLSJqTJrskPMOO22ISibBpcfmw1V6LH9wqo6C10KIg4NS+1HOJN/+xKJqpA0pxImxNOin4v9ENGAT4p43Ry50gaFx55NXjd7KrDo"
`endif