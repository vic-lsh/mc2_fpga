// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Bix2p2VOeVEMeANX0gJDiaJnw3OVTGuGr2rBZaCmwsYh7ek1S7BaCZ4aIuzX
7xHS2Z/2dgZA0lihtYPKtheuCRNqXBnO/CsbcsOqnRg5gjot+R2IfdHVrckb
m7eyQFsl7+ArMES12jrWUpgbmDuXtO3KiyOoRR6jIAVs+tz/0ajLaHxyflWv
/wdMURKJHymKgbU68VORTx8ubi0hphsZJbfV3aFO4X7cVmZYV+dAH5lfdreA
sN9P/LbU7QyhyJq9j2yXmD4RNmdmrZnwCDNFfeimT6Rd9ZacYSPANwOXCk9U
vvu5npx0EfV2Zq9aHRN8obXWQj8mRAz4+/iQ9AN93A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
O5Ke14jYzWfCcHFQlv4vmWUzaWWN8ELfb2ekIiFVFSCy/5Q5QCobV8h0kvEw
MxR9t5JfFDQANP/71VJ89PpBroqeqjpg8Ve80rj8yUjC0hI07ATTJTJMkq3Q
YxKKL1SaG7gJqLSOZqTtVFvC0bAOUg1tXJmB3LCWWlYJllduwv7hjRlRnX/n
Bpep+63IJIX805znLbMOaEQES7JrNsEk4oilBIzHFrbGnNY8DIQS2BItpcZ8
niCUwPv2AB48JrA+O9MT8Y5dL/UGfZQcqTxVO1Gmckgtci7H0U0BCshRQS7+
aCDtis5RFyzxO17r5L/xXVAvI4LRv2fdNcNMuHLOYA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
P2/iVlPoV1uGT2/bXEdSHZ3AS5Po23pSq9c71NPhcwB5Hfu7XTRUCMU9l/ZR
s3i1QbEoRpJ+HiOOG9Ql5x/+tyUJsYdCA4W/Hm7TXWdm61jvC8PSoO9DRf/8
ewZ3xIOcyk9dhnUPSYSHjwujMEZqxtM/GBRrbE7TU0iQX+857jV/yW/RK9jh
C5gF5CHxKZlK8LV4QuoFUq3htAF7CND1mi2yKe0Yead4k72PaJ/JGjg1DoPc
NubwdxAmKDcLFht9Lui7w94IdaVoBpqP1lj6mlQ/n4rNFYY+IuMxk69ZhHnB
Kkw4dvWS2czAWcjKfb5S6zVisZsPuAoAXBD4w5w69w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pLD9gjDI0GhZqGkMrDEYt9OdkatnQfaId0LipLRYklO70bi05PARDgdq3jI/
et7vnENc0abKkrTDdahJtkxF/hs5mGHq5HuVfxFWXu2I0Lq4XY1QqS86lrn1
tiwsBEXGsEAA6IvS9ByzjpgGqFXccyHtixIgDcokWpmB5lTP6wEbh8k4LFY3
cIe6xvk7dgXXCRSNka/hUU9v+WFwd6hXFvIrEknmGvHNsAQ1PfX1NwRXoqkN
rW7sRt4E8YPVZbdOiYpcaUDqgk6sjv8JReust98WwAGgjd9n7qRFm5uaAE8f
zPPZGS1Sx1vfgwQiVMez9mQStr41MKd7im4cqQk9Wg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VAp6UGiULZ38KDKq5wUw/CLmhwAp4T+JZYUUbtyvMWylcYGx/pNdi4nYxDdB
mQlzwhqFDBZouaO6v36HyO5ANFjNOTzcEETHyOUb1MD2qHaAxHR75sIxGTqE
0Dx14a3nlA7qpWfej5yJAC3zgNXwbuLoj1kzcozW9aQsszaP+zQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Akh85b5RHMzmXngJomwLFmZFTHRzBIHuIsJ9NO5ODLO8nJNUWSVR8CcxWp4K
1K09LEgLe4QCXTDkYndu1Ha+qoBEPKxuceKtia/CkVp/mw9bLa5wWaDO1mkC
pKm+09u5fZaBXqRXodIb3t+LP6xBS2bDNhstIwg/BDcdiVs1ajBGLhU6b1dt
xfGblrEd0fvqye4bheBwpfDxzFu09OtBcX64fTU56mW6qp4MODKj0/Jorxwe
eNLdcTXraV32Y4Q29K1R4DYd0iFADIBR5xYYViP840X5k2hYOCG2/U/uVD+q
YEzG49TvdJ/rhla2r/xwHuQFC2KTiK98gO0stoS6X4DZuOSMXsmpOXO70mj/
w5+kWvwe8JxK1QEZ2DKGMoFNGFQXEwvZ+xyP9ix5tNxoUgZo7O6tWSMggCp4
e/N6A13NpOJ/j0E1ssFqi/a25gJDoK+Ds7uPQGf4OfducRVE4Onu6tIhpFBZ
iLKa/XAcVvXJHIqhNlLOZt+T+9FIvDA7


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rkOh6G/+j3L7feQ3GSQMaPTQ1AUU+PPdmLSnUNiKelhs0PrGd8Huz1zyKyIp
QTiW3KzLH3YQ98kDcXRmMvVhTbO3CmPcltWBpK/gcMrUk1vOTInqXlHQZb7T
XcYXwhl5YtKPDsQ0XCPzxqdOVrGy+rwgo0mOSNCZSYw6hRsuS0o=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uHpctLcskvl43nnKONAhAIbqeZ7gIf53em08KRikzhhdu0VvVveyhaNXMXoG
i1MJ3eZiIXSVhwtQEooGp+LeWhPbd15GemteQ9413Bohc2b7nw4fjUhA6dVb
0IlJnDcAt1SrN64PIZdaEjPfXdzC7JzK7kheMk6HdVXjcamOX+Y=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1024)
`pragma protect data_block
U85Bxn+jrb/vbGVMDXewfWmerROmYDRi2U+0rvvmLIsmAFh2imht2ieLegSJ
bphU78KzJzyGlBzJvdYK6HomcpF+suO2W/WrIJZWYKTNQT064Vh5N3tT0m8g
9DgQsW2yQEfVprXBqJLr9L2GMgSxSX3n9M+8Hg0avy1xCYFWzdbhLTI0YA5Y
nFFXJo7V9T7enwRF1sZDeHU4HZPFE9w6rshPawPB71sbsk8QWXpbF1NTKonJ
vMPYSInN8rX84Vut7T20o4sj0iXziBHGsGYjyc+GDS/RQ9CoX9mJuON1r3UI
5kGWLBlDTNuvCfma+fl1aHbCdjteQY/YxKAb/aQUoin9p5HGKjw6foO/I8sW
dovo5T+b39zG0oUK49Tol4uIrLsN3uXoZselHZSVEBhei0U0TiMszz/SkyqW
YIM6fT59FOXLS5X+0Nh2uElLCU9wHy9PeYDMl/ui8+bUXwMDtPhmYxZ0k7w2
tZB0TnYukYNmXkMhSyVEgx0ROt7IsmQdd5iLFyP+Ya4qj3YuRZC1aMpbrFQ+
6774Y9trJ654B7kOVEY1xZH7Wv2QOs169NQ2hR9QCIjMBZyE6n3FryoKAraF
zCBKR7ibXf24xclr+3yK7x4RbOZ6n6bazH8WuCp1bO+UZtPFPVi8THE4fmSr
2TP07qJiv3HW7Xt+u5286DSUVGgsf/JdZoaWhWK5N1y/tXPM0EKI6ydZeabd
w2wEFiwjD6Z3apK3BeSG3ouiqWsgto4wSrwoKnHYt2dfRl+EXmdtn4Ziq3TT
Zo6DVovUnpAOSOWWyCU2XNJYQVcAN8hPumfsVV3gBP5IPo0xisVrNLfWP5cx
w8BTPCreSHcXLcNLlT2wglbubjuycaiYtdj0gi0PGWzPzDOtqGPSuqYnOvON
sykg6t0q4EyEeClEf1C7SE9/ef2jTjaw9BBus9LdQ7mqFqxV0PIB3ZTccuBg
qKtXLMsnc2Qkxlv4jpnpOM6ho6kGBd87OBRq1S2NCN/LT9SKvSkpLZDDw0AF
hFygfIm6WMzqL29b7Rtufczk+wnjQI7qOGWN1Gd+pj5G9hjNlqFu/80ByctZ
ayKfqbxq08XfX9JOJtO6uqNC5pIAtCiK9EsYe2AHgUsGoH3EF93G63UkLJ44
gr9Mw7vn9iP6PUw33XFzkUUQNmby857UUIdncmGka5K3t9CS8Ryn6p4Au26C
iawKfDE45VtzkdOW/rUNj/81w4tBJ8Dd/UPU/eF1CrTvFftUS+NzHl52K6Hh
CjUPGlgnXG4ZrtUnVfcVKlBwRIqY6jLbgjum5fO5LA0lUjd5gE0M0p7IUXOv
PxUAKNrzfDFPHUMNJAiAugokInVGkpL6WS/PVZdfheqwjw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fidd1oyAhusLLJ6+7Y4fW+UxvqV+8TisWbzB76p8J7jCbedVkgTXiBKrUzNVBIRDckfBwS/gk4qyrpXnk44TsazVN20DO3TdF1x8MmH2pGcTjxrJqgYV/z3UJLaYPiY1WrKUNRPOAuHkyYvfI5GoAsKohhmpB04sGLV6+cGIymx/RXK+eIUgAROf9S5AOXsk1U/Lqv4gR7i2yfj3c/IhJWMX+Ld3X1LJ1lp+Ly9OQoxuxuw6FJswAGvwHs+Bb/A+ukplfeXGwq2wl20SauKvg46/VwD6/y70X1zYIRr88eVQPP3xEN6uqeG4qV0u3QmWGzm9LpITAOeoYScHQ3TSvcefh4RE0bAp3cTnyPLDcHkBsVLxZmzVhO2LwT8UqxTs18KFinrhOq/xxmaR+BW6PTlPDOyqAM17yHSmSAP8von9O5wNGaWEXF6csxZuCNQZ/uAhufa3gtu7wD2/LklYfzNmu/BjoDQEmtBTqxjA/MyFWMgM+EeNVzYW/dSdIIlNEnBfN659AdmItK2a1l9EE0RVlbIVlod+6rrWnrDN3qq1lE4Hn2CHWKvu9mVdbQBWve57x8uuDGZPyr/2rZsaEbR2FuffEex086soKhIwSCL7sen2EnomFLx8Kgb4CVQj4LorV/tj7Bc2yWLlwcEvA/qEdPEJATSstrB0Nrkj6+/afP0idZlw2XoPXzUop5EBrhKH1nEEDyhb03OKbz6XbviKREmXdRVhocbBlyXgL6ARaXjRmBQJXEJBz2rfi/9hWiGqDZ1OiUX6NM+qpxH8l/GKFNlsHSz92XltzjKqkqkSkY1kHvp7hOndVbbeIyDi8ZeyoGqfhShCjMACjKFKda3Y7k+JAM/TMY7WT/wn/G/K/+whrJ/yQDg5+EmuQCjBlkFC8m0cFY0ZglvvVpsG52Wk/PCUggCLwtdizOzWyhgoJ8IGpc4nhmHHrLCMeHqHapkI3imuIdixJ4eY79suef8hASS4FaQQOnZcJQ7h2AI+8vlw05v088ZavQlxz5NG"
`endif