// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
n1jP922JkGqT5dOcbG9thc7m9VSBoSQyBxDvSu5ayvGTNvM+SDTzl0DeWwd2
3ZYzlcUrcoF8NN3rkDoqdxyoVuhWZSWUd0JyVQMibWQtVQRN+ae+vJ57+j0E
mWRqkMoQ4EWUrQTNQQxeVHK7T+T322vNImdIv9r6ikPfBHnSF6QQ6yuU3Ja6
LGoJw/KmCJPBWhv5XMEjPfLl8qL623+6q5se7X9wkhm6glT+rtEcNwTJRUIr
AqI/R3/VmUDCvkYf2U0BaUp9AMEnwtut3dhmQDbnTHva/x6B72RZqB3H+5hS
E1gsfKaVR6+AFLIg0iLCm5Rb4ICwySAPZxaSKDb3Yw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
h6cs76VOZnZDxHayGc2hcdE55Rs0/zN37D3KLjFth2hcJc+Udj6DihRq+ycs
HJCweBHl0v1Dyp3bZsw8KE17HZ943Ho8rP7zG5e+pAmA1d7HYMGheF7EHc6B
h+zOrimE13xgSswNhlC07soDCfPtxGLVMzESqDqwSyIfmnFgIniwTV5+c9Gk
2XMEgBOrxGFdrIdhajgA/NL+FUkfje6z1UXRSz/MIQ6xw9KcvJiq+g2T53cr
YTsBBhldQag1B60ck4R7WfGVrQU4idqaGo99BMSuxNCYBNNq6hL/yR+Pcjh0
h4/9N/hC1QJyWp7hPqMQi8NUwPyzTvruHbfLdnUgLg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hnQGQPUvb6x5FvB2yG2RMIu+5TmAuoViAq5lDrbR3oPGCnPTwDR9jJwOLS4S
t5LVDY3dIsq1hH8wRwf7JJTvie/NzvNPHkmoYneUrzYVpq10Ypu3Dyz7bxFE
5/MevdDpzFgqjZwkvbhgF2oeYEAptiCObhnxw12xZSQXERPo/D94QhE5VqxH
VVJ4G2xdZ4V6NVui9U+OpmoHFG5ZDEOHiCa4TcJHBxOG6KfwMg8l+6uO/c6N
H6sOjjh9lrFeEeXNb5kKuxKx4tszjLeuN4xNTd10ztiERQeP3n2RSGn6K89N
Hl+ROzedm/OD2nnHqDs2Q2+B1/C8gvDNPArQXctVnw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IkHBLlicAGFzfXRpQUNhwrfcOMSyuFmkNqid8FFSogCf5Sd8EGbrN36uRTp+
BElWCsrqGcbSkqtIIp+/P4ANunrqsYqSEq8ahuw6tHvvZ2qurh2Tk6x9uqFn
2DrDMJoiF1OE1aYbresV0Uduj+kkkh2sHmFImh9F2SeamCHckmZV/IV+/MKQ
3H4DK0jmQ8diQLUHGILUp2YJoeiVlHUpXijvF+wkDjgzGkUv7TGM9lKRTbao
N3xJijIAIukImWEzg4imYpFe0kTz43QdWqFCzaVTtUf6eO5UBP6EilgRlFRS
Pr2GU8rfguPFxm2/azZqSagulQ/W+ypmhDUnQ4fVZQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DmmGq88wsiggsAb4HLCcc3r356laBphyCxsqeHc/YS5X/PcmpbxbOo9SuJym
V5HcdQcgCbc55e4gg9qYZs/KNQVp7rBsEmVdu5Peoxhal5UgIJZNt3W44o6s
xPGt+J8mzRxGBaRj8I7AkfvKHX1tBuqeCKILT9508UMJ+4KhAZc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
B5BYmLMWyUAD040VQClDymRr/tjCI1EjSSJYzX3Uc7cFt2ZYPJrn3Slq+/F2
XJNOwH6pAXb/WX1EbjuK6BAQuo9jPNPAjOdxTiwd5fbi50RJ9cNrV0V+RopS
7JCHjd6NgU2inbUMQ14Vq/BZza6UnV+4PuctQTcORoRUV3r6o5Tk6swcFoQW
bnfkEnuyk9q8QEjHAJhQ7KAQehpHCPpH+kxj5eQTObRknOx9myGokaXJsmJm
EWWModK7etHERgneHSeWJNORhAsfP5E22HxPwZYc5Tw0H1yV+HiVfUubfluy
SQ/lEnKn/C57/Sxy8tv+MSk9jg9SFJkU+u1DM9ckaE27CPo+SoAuw37sW7Lj
tM1kfNW1uvx+N3IOl+tj3fQsM3setuIuQ4GIAcz+Hk8+RjJaOOVHCx3kmSA+
iG+RSKexYRCqiGXPQTD+xB7JLPignqXyvaFI7hDZkplL6wLOnCGBA7uwGIU3
8fBJelpd88hGenal6fgl79eRGv6PnR/Y


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KDdMRO5sdNNem/zv0wIQq80+gomAVGiLpAqShXGromwDxslNo9jgt9vL6KJ8
7QBrB2dnJWbce3nSYLCFT1bsZEme7NJuR5XID413392Ng8RMM0Kxw+qnTCpy
lz+aYUdoS2kYPe3n/x/25LQnF2lYYjtFtRkS4UYkDxY72JeX4n0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gIoNeOhi+617XfhCNaIDtM8zD5Wu8L3suISv2is9bjo6uGDT/Lln/SJv9E9Q
ftdHcQzWXj4tkEHx6E1awB9Pg+v1dfq0BuTBtQioezLhpor0hBAZGuCs65C0
ZCmHk3lUvp1zaOHdx0YL7ReeQ7RziUsNl0UMH3X5rT3zZdXc0es=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1104)
`pragma protect data_block
gEPtFENGVy5UWcDOTlJHbcKtJSq5THjbqMgKdFB1m37IyMKZmNS9wkBl4Q0y
lo2Dr6OVsxhFJSBMOur5ILxrfyE5Q2gKuH1ZtnQb4ATsGGWXUHrb0R2cBKI6
gQgvT98J6cg1z2ETKdry85fGb4DXT8xV/M3brqwncaZWuFB0kVZ8BQeZEGj/
Z625SaHglo/p5PGGtWZzHNB2G2fmIr23a59yaM2YEB3q9Mb58bEONj0yrp1H
9eXwXehIyYZ2G1aN5fNJJTEAAkvs68B23Wh5qf+0lxEwfXrvzrpxIDhIODHL
v1jtYvJZhtfrqRc0CIAcOClWN1lmNYNM/K5Rn9SZTMMRKePZyui+E1RKbn+K
gGekbCFBa9knsUdehwg15OomX1LQawk3/9zrP8taI8yWsc+9Wzp4Vw55stmK
PTBgaW4DTY8aoklEyZIgFPSyDFhwv6ANqh06fobJ3kEBNdX1RAzPzRVE4Jw6
XcNB/Cb5Mc3fuFc505I3qmadvBlQwOm8qcf2NrGbnItSkxrJqA39iOrWLPBh
/mlG6jKaeHCwIpFL3CbN2TgWRgzvpUKIQo3FWgf+V9gd9KOQlKHhNg2de57/
i5IcLazMY/wImzFeWnRiw5oruDwfd5Lu1RObD6WyqDAAnP0XtLykQKZXfO+a
+f81tIL36dJfvItct5va/DeHbHeDXFVPqvMzK+NIIl4bq0aQ/7bBWq9m7yOe
ZsFSVg+REZ+Zd/IB4hdueJ5im46ZykKrtGiOsoOGjy+Y8BFkmqZwbysGU/Pa
GVEb952j8kTlGJc3qHvf/09dm4AOcmp7YhoESM8CwvqHyoEq87QU73PTPZic
vILkFZLFHWD876u3j2DWoCYqdQrhx+5mS9lGIoJhmG5kaE3GRC7b5wEJu/fu
r08sNwmN3UZPC77tZ/tnbG6Ot4spOkK5TEC8rhIYzkJv79+6RMCm4+ydek/K
wqcBPUsfZEZBm1pVqd1UYOK8fc7vuFFr1SyEhEJMZYWK0TPs5d3g9LbpPad/
nwzu8UqdUsXr1I4t1aFQov0+XGdUPvJ51ABvCliIawri5vMruyOTd4jxCyLq
fSMfiCRydN6tAQdHmHn3bGejWptzEeAFnZwCr09Nl5+Jus1VS9XmQTKzw6a+
DCqd2P+yhNdDERg0w2IojZgifWzcXCbDTwsxQp+iyp2i4vHehY+QEY9KLIwD
xlCwS901BwU4jlb7PvJOEEIm7TO47fpw/GOjaH8dTW2MUSchKcNYm/iXn/hj
Og/4V+5q8vluRB0/UnO5X2R91rG+Vqpqed4IB3MWRGY8Vqqjt5AP9qec7Ulp
SK+Eud5F8JuNBQErtb0o2+cXiaWORuKHkulYR8ORQCkb1iT4iLijZ0FXM4Jc
wXBaq3sxrmecQIBAqAcJRSY6qIUpuIFSgI1DRDRAdlwyTlfAUkCO3J6ek1R3
LFKLkuqznlu/skN9ZnS9cBs50R9myRJF

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fidd1oyAhusLLJ6+7Y4fW+UxvqV+8TisWbzB76p8J7jCbedVkgTXiBKrUzNVBIRDckfBwS/gk4qyrpXnk44TsazVN20DO3TdF1x8MmH2pGcTjxrJqgYV/z3UJLaYPiY1WrKUNRPOAuHkyYvfI5GoAsKohhmpB04sGLV6+cGIymx/RXK+eIUgAROf9S5AOXsk1U/Lqv4gR7i2yfj3c/IhJWMX+Ld3X1LJ1lp+Ly9OQoxWQs5Q9QDi+FsPhd4lzFIo5YGdUeNnjTWgUHtdSapa1YhI3X/6+v+gUUMjf0ey5qTEeGiEDXllxHwAbtSH/Nf463P8vIuEodD8/1SwxNEYgGwGA1l65SGiyAFooIstlT3mXz5iyBOH4baLWcF41k4UYzeGB2TN++pXieyITgQ6bBg7M0Tk8Qo/R+ri+/RSPC/vS9LDubix4SeK8RF4L07ZcPF6uposGZW8gSPK60bEnPbqF1GKwOG/Sl/yQACJOojaatwVI2hFog4iXLmWCZOnHRmgHRKNQzDU3cvGEL5j6PiqIr4XrVvBtvV1Rk/vJgTwpcwzPJXh5gcgCMjNG7Nwy/oJYu3Ej5aymM/Y8S26GlmAzK2/44EVYSpf2mM4RUBvivmwY2HEyzXy3eE9b/ghFWt+N+bMFuic4pQewEznZPWrOX34mOhOZ5MshF/UOaEnRlBOsRCqC7jA/eNG2U3fiTiQZlLyQyoa1dzNaK0doVKiytgwCY4Uq1CbXlnl7ZZBRp5Y0axFT8SfXanhpo4vsJO5mcOSnGvjryCY1kofCw1pqLdsLZc9KT0lVc6qCzRkxbnZwDmAs7zGSaaloaePdYofja0ta4OLP5UzqHLhZ8mhMobM2r5gWcV1OoiKPkKyiYwwh9GA0op2b5HwQVzOMl3ayQvaHbKviaatwZrSGHTUCKRdd0PLNwTDNZNnb5T2ZwdoIVx94sfTSCiT55nfd9+9idx4OYkF1PN7jhmctySwBYAnuNeCEgPL+fLJQPHBVf60pr5YN3YuOIwHxHkd"
`endif