// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
t9DRPDEjrg7niEDD7dtMr4aVSdD9jqBY/12I1cJPTXDXs6vd0OrahWiGt4Xt
6YM73LJizcEFiiuAPXmbi/BZrkXuy8sEoZnRQbk/LnRHPyGQYnBC0Bi6DIH2
CCf1DweVivM+l2um1SCbTx39G94ELwjT+NwwoeFHMmOAGynmc+jrP1RU2yLe
tK6eamuSqI2Dm4oa1nTD0rhQiHqlvNk1qDRFm/BB/qhhnsBk3jYahI/Xw9P9
l8E7UBt1KsaG0vXexs1uhekn4f2IJLI52AtyFLus6ls8pKLCT0EkseSbUwgb
SRc+RYyecwpBBOlftUkY8IAfEmrD1FK//9fIk438aw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MHRHIwnUERdvDZZ2ZsuKqy1L3Gjixy34bP6qJv0B722abZt7+9gUnfM5+ySk
y6a2MqOjnOkOf8jX/s6DOnZN9pKTEbYvv2MBsPkc06jgycedGj7ReQ5nlz+5
aAKFO8LwMUDo56zOAfxY/+DW39FJktoEbxMVIlW3BBZ0Y8nzXRmDZIs7O+78
FeQEptP15dnZctoqqOYpAm1aMBSgh/4/N6paLjQ+9uBSuzohonRWk2fDVywI
oPsrjkTDtlzYCxAY3zgeu/6Pf3k2iBIREXI1HfbBFyWCyMihs9QrOIWUuxzo
9JLBvSqtWRSCSoXJIL+QiImvFX5JrzrIdlWbkfMbvA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UZ58HxVDIQfNhBj5XuMN8ZgqM5D9dRGWKWv57MwGCl1J2vd0KVLX7PSWUnlP
gkLNeP8C42jruXoueXpGsV5k0ctMN79BCRhBA2vsizQ2r4KepXQP4fyRVXUN
xZIB2ozHUnCCeHOTG3t6MKg3tiXP/HLb8pOptAE8tL9Tvn7TgD/cxgDJlXJw
CtlIpnM23YRKSaC296hKHNvG2jqoFYcopRZkDYefz6Lt44jovPee6UTV8XBd
62aFCaBrMq29R0HHllcepuakN7ZOeDrvmH9bc3ZKAnmFJwLdr+WXiWj+I5Wx
8/sBf7dbA2gKUyIvRvgGId8B6IzCxjEoiNSXu7rNgg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Rc9zeNw4lLxi+FxBlGdGjwbu+JzbGCoKjpIIotUdMGkE4lNw8A9mNFncIag2
EjGWffpzCT4UMxPCD60Q6afz5T8wV8GSa77V922A7sBGFB9TfAJZHansWV0K
SxeU9JzoNtVfLPqy2dtg4qtD3x9DS4PV74plgzmJCgAa7Bi5sjhr3y4Xmqy+
ba23F6nQRxaayYcZTUWBepFfQivTn7d/QY569sCBIk6ude91o6vQad3lvDJJ
84AVpJ20UChSQiGOvXLja2Af0YNMkrmHOcxAIpaqkmCAC/83kc4fM1zZaHgv
U4jwZ4Z/MfuUVx9ImkdATcdlMW/sorFHlcBKNe/vOw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KDCGmbk9TpfyE6NV7W4kQWAZNPoJx/6b/IKkxIYLBU5qojJ/78IS8UIGYFm0
hczdENj7KgbuYhA1YhIBGAQbEFKp2GpiExeQ7nhGStZbgZynO9gB3IQGy5vF
Ie0NTgnRfmKrywmAATGOnw+I/CUmftY3DwzbFgGiAwN6E3GVasM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
W7xreEomXAKKa3F5B7Q5fEacpFuiZKxF/Yi41Rxi+vm/DpWKxH/qLRnwrrd/
xYsek47ILb3ZXEu8VTFgO5/zO2K3hO2AOItGmtnHIdj81jnxzJR3pg/7dgj+
PGBrW+Nu5uBOjSFFxbEJz0ePSiGpd8sLmKtk44E5HJSpjkVWX8spuFhW+qtD
D0uD+YtKSXavEY0byfGmzGuDX7tJ3DR654FCMV9yZa78946CPErmRkwfgISg
4NUFTfocadDDTbRKTdzNRicte61eWAIiDLk5VUp9+N0kvJIroLdVjimJbJv3
O8Zb7VaQkA9dgKCNPRZv07gwXoKMtxxaE/NfTAUKvRqevl4znFoW+2HcZgPS
h/bRgBcQNNlMNmrCJa/zCw4eF9rqde6VjO/6Lze+my8JzgauYeDDINDQ5fRb
f7Rxg/0Ez1JDUkO2s6v1R5zKg02UvUTIuq352m/EkgSlRL2b0epGkJ1c5yi1
JZvEORSUleGrJM4ScXdAzeKs7t8Cpkd5


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PKerADqUJOeEBUV4Lj0mWCfmtwBqqfJ0U0oS3g+ji6lKSR3Rpil8oRI9k7LC
p+GHhMtzn0XkGdyAkB0dsoAsQGZ/0VBVF1y5AGj8LMG3Ehum87gfxg0n/WCW
/YYoloVM3eScHbWAn3QH9CIa0QtuXnurWsd705lNMyaYsJiLUTk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KQPOHgbtJNfVfwZuoBJXjBLy8a7CY1OaZw2wL3XgquHZVUufxbDGI0ArHNh3
sZvr4x1ynrqJj1bL9InEP7hYTxH4VEgDahvXmoU5cSmx3Qqu/lG3aj2isAyP
zEsnkVVR5x7uZqUr1/+AUg3hECL81Ku8/DGe8JgKv5xlWG9WYCw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1104)
`pragma protect data_block
kYH9z7sADMnjJfT2Khe1AU2/JUznKksyJUjS/HYqRYzxUnH7nJKIQVJNzlRY
tF5WSrjzJpMCTafcSsspo4v1TDgzBfNQvecJZRd/3R+L231pfF+GxZwt/q+5
jll+28NUKV9n2eyn4/84FAa6lMMkxvB304iM1ZO0rS3dueMMKzHm8Y2FbHOp
AZQv83xy3fICfitvAvetkjy1ujoJa1QEH/hrrhht3QjFbYTejSYTg/ApN3bj
7PjFODoGg/2zqjB4lLcCB0TqSIAeuFFBEKhf/nIP4gSbCyghF5qrSfyUX5PC
SecxCfUXpW4G9qMZaFxTHAdhu6ymeYZBzYytHwyVEQZ7XeK9uUdieO0SZT9z
GRBERxWZ9lv5XsCDRouqeTJqLHEkVJcLkyBMcnSXi1AgMLsutqhJ4/9DsEwv
55NQipky6SIlBXxXTVvnuA4IhO+cj9sX02OqBf/baYVT1rDhNbe4bz2hpOcj
drR+31fSux8rqObkkffMC7TqdwXl9ze6xcIv1w12eYZbMOVOBkplOJkI10GG
e9jLs/447Ppz9Lea+nVVwmMIlbS7e7J4Np725m62Wy4/mXcOkpm2bhKZMoIO
KwmUbbsf2gJ5s+9YEIOcydycDy0fa6X0MDX4QaEkvvlVNn2soU+K3+nE4Qb/
Lb4BCNVS+KzZQDpXT3667gDDBQqnUxAyh6/m2yI77ANlNYupcr0AV6+s+Ndc
LOU1q+G6hpUdRQkQePI/Vb5iV6YiNREz/8inAgzKMd19lGUo3xx+mx3R28T2
pv29J1gXuDD1M0a8uO4vquLyjyl1yNWY3iADpGR6v5S+09VbCwVMvXpJ9hOq
UHRkIhZHDlNMYcm0GkGHYDMYzH/8Z1Wv0eJbJcajMy+aKkb18+LOPADNQNnl
WBz8/CEyYDr0A6M9AJeBCZDQzDNDprQ6VHCAx3gUpiruCEF/mpUUh3m8HHxP
9VQMJVDw9gFw4FgPRq/unmHluBaAwR4ZXnWmwLw+EIrrvKrRdP5UfB454LN5
7plPszFedNXMBjVO5MyE/KfgfXAZyzoa9SV39Eutti/1cv5AzXD/cNWucN+/
6DapuKYsTEdKwHcYq5NC6PmOR1X4njeZ4Foox9VrmjACDar1+yQGZNZm/Nev
b8sOJJz30IYq7RfkebRUGb6f+ZL/Parr6h3pX/EhgzBDRonpe1JqIaLdnn7e
goV1uilyMt7u5/W0lWWwJIkoJDMCuI6BzqKIyKzTRxfGLJMESFF5lBSEU87R
EnnAN2zNQ66vyIS4x3/4hojbmratSuoqrsJKavcWNaHX4G4sb6m7Fo+NrE6/
Fnh6rv5bIFVoEHb97R8W5csyuthmMtFI/Qf/Vr7r3PeSOY6sbOUy50ND5uT7
tkYeJWteDs2fW0rMnYCbdRprBRA0/e8KV57KWdje+VakBbGzHRkMCuoK+ZLb
sUp0wL3CRFx0remP+H8FGzLWOY08yW7c

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fidd1oyAhusLLJ6+7Y4fW+UxvqV+8TisWbzB76p8J7jCbedVkgTXiBKrUzNVBIRDckfBwS/gk4qyrpXnk44TsazVN20DO3TdF1x8MmH2pGcTjxrJqgYV/z3UJLaYPiY1WrKUNRPOAuHkyYvfI5GoAsKohhmpB04sGLV6+cGIymx/RXK+eIUgAROf9S5AOXsk1U/Lqv4gR7i2yfj3c/IhJWMX+Ld3X1LJ1lp+Ly9OQoyIXZ9x9OTIsyFwhxN6GZihAPEpliH+ai9Mo9ugPTmg4CGpD+4TcMXO/FDaFG7pjs5+SixwfqO6dQrxpGGJQuWClRg8g/IxzM3ooI/DgMa9PIqwa/T8njTehHMdGhvppLjMe8s6SbtRkcguQ8jHInj9UaYGEEJy/kFwpO8ziVohuegewbKjoOOJm/7OG8rdXtdlObV+z1SPuxEPK86oqNL4Ui2wIwMfaDv+gAbHKcfR6VSYJGltHfskVnowLM1Z2q5RLHLNp/28OVihGO9p391Ck67LbK4r32mI8XyTTD6Hg5eaSXOn5r6zTu8mwjus1km4bMh+eSs/GJEGkkJdyGsQN1N2q3h9CYFUVKRXnmnfAjPi+BdXmAh4IctZ6ILUFlHbEpIEPURYBneqbXOM+CuqlyX2FunPKlOjnAQ6hrm235pHoErt2NOlcL2AUZGabztL6VBUUo1TlEfOLDuBzoNos7RT0QXn+B5lnzTEXFPPi4GdAF+qKY6Y5vD0DVGxFkQ7sfG6SkyL6qiBmt6yLt0dd1Yp1PH1ZaoI79QUuIMbQQ1VUzAReP8qJHaDHxP+9GL4igGkL5Ghz/jFnV/2DTA+z+wHRBvexRTgoaX5YiXMBM6vBoK3WZhXjHTSnuDmPApjwHXTdLoZaC/TCEhhg+5jWAGonPjsQH77ObHnAE5AbwdLsMAzopK1lxLq4hOxLGJl/MJ9r009rks6d3Y5WNIX4ZokmO2kvvULiMmbKx0gcczF4T5tpRqlF6jc9c2wrCl6blfxXIQe0gCtNymLOL5g"
`endif