// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aqFBHMoQ7proq9c6N1aW08UafUHIXzOAGQPqtroRhVbqcSWDWhnb1QThoTbZ
zlUBTiNXkBIak2BUXjqaq5wEW6r2Q/MGYctSj6fXdnPFLxjOG7cDr1tS2ldv
8sbQB+Knskirj9hpFQ0tcXLr8XwR1beSwg90sZMl03f753yboaj0dTW1KUSf
Rzo16+gvX8J+Yb1JNYP+SthaQ11Eq010ciFXtkhwBOpSFqUBG3k8Nmi+qi8L
EjWvWEU9Nf88XI2JA9kVDx8860FLJPeMeTzssNmQuTe8PBP/Z4X3X6c1LUNS
5ZdweNR4vrK4PeuN4uh96WO9962yDGBblSI0Fp+ZBg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Fu+2gfp4rCqva4uIG8orJ5tZJD0VSf+ROfsS15E6hn5AUGxIP40aAwlfVHoF
wcgRfT1ProZkDPwXGf3r81awtbUhC2uBm5a0VljpninW+RpqLEwnXfwfiWEf
dAbrgUF7eQSitiWuDRyN3gnOurrcYYsJswtNMc2/Q0PHl3y893JbESCwLDcx
pka/F0Qn6sZywg2ua+jgZ8w/oDKcDBjj5zk7amBIs8eNgsZJiBHb8jdpxjAx
6jCb6XOy/b498WFvU+9uKqrFwgDFZq5oMFWjatrSI+HxN2t4pReaknzAmJPa
Kcl6olj5NKTZ/AzuOLmXOtbxVIJb5ZRvfRZyWG683Q==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RWdcTM2MPy8tGfqzK0/O57PcsZF1APOosO228VLZXyIVj7f/5Kf6Nyq1RyZ5
7Rh2Pzp0AHU9JUIJOcyDjNwbajO5XsTFXEPoNj0nDj1u1toEUPaaOJv77jRS
JpyjG3y4TVZdKdHkPENTQywNyvavQzjH/FIv5pbZJV4CM2yzH02NnQWwmm0C
FPXmNLoyuL1Xx50BrTh5rRs3E/eKlbNY7MAXQ194QNwlpLUAW4mX3a8bUkP8
tdjYAXBt8cL2XYVhEPFFH7POltpq0Pi+Dp0cZEUTLx8kOA8qcW7rI3pKPkH6
sI6GQ5r6q9KxhU131Xh5WzYwFv1dSh4/leCR2Ta+Rg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
L2u99+GnwhZCQQ1X3TyOnxZ8Jkscth4yJaLHzom+VhjjPGoEGQBHV8N3Aj1E
p8JSF94WisqxP6dlcQXRvHTVd6JAg1IdG7zfu2NIfRWDs8QrPgP/laBTcPqK
XjyaucGmzmoTKridmXnl8hkzNry2Rojo/vW82Gl84KAXvdfBqFy/dpPB/5n0
VmPMnyb7w0LhRbLgzglw2ZemAH5eVFVW8VZQxy61n2+YecXxqsQdiyIijWi2
Ns3UEtNBOJhzWZGkiWP2QcBh9Qfs4+v5YVGuNrF/m5UxSbKV2ECLb3NktABy
fLSeLlCuIWyHkGX0sSMa8z0ZseMv8QdZstHqj9mJGA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ki6BuCyJRmwSm9cC5lR2EDAyWFNml2g2sV5EMHS4bzkEFizZ5mzsyhc4QoXI
iQvPMUgfz+5IQDzvgC/xCYXk9Oxd9ni2SsWfRIFDJFusCPXkVeAsXVt3K6WU
y95etcnzcZwAUsJBUr2McgIBT1gUHotr0EKRo7gOpIUr2Np11Lc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
MEWZsnkzX2RLsQyjJMs3IgKmzTl59euUkkfa5TixmM0aIm5AFZll2/owcLQ6
mCrG0iYk1aW0AQsOGrxM6U94qyeYbCVaX7zhnXwKhmpInnb2QLVpTR1EdquF
p85hAdheqgPOyN1XqjABqKuEdbUJnHRE6lEVhrPncQoWeocZpIRZRqTlqevS
ERBK15Fuj/5Ww0P8KEhDfQyZErSL+yVgZRPRFEMxuN/xWyGREy4cOcMnQAKt
7HFameMWRrhg6mR4dLv21DnZ11Wcn9a8I1CBbtj+5OWnw29ZEEcDNvvzmjAc
niaQTNOzabvIbjL4eIz403z9tUOG6hnExON9JIi1mO8ao/+zd1hh/wD1icSL
mti570balgQ5NPh0u/npqWyr0QHFIJuX8J5klRcwVLAwuTHF40mIWZ3oh2nD
yRW3bdP4Kv2fTOJ+YVF9R845adgQH4I/iAVV8VdxStyRYYA/YYAcchZcsqbT
tMLNvyvfeiypviojcmaDqU/J84cr+6dJ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cKrHxdCt4jt7femSXHAPB2UbKWKodJzi8Ni+Su5DAd96Wp8mw00wuLXLvtEW
ozHuGrbGn897XWbmFTxhHK/Ju4zyjCnP0+MJta7LrZ1lGfm9H1R2ic2dym6j
oO2ag6ftBlAFisG1dmTFSlHVTob163d5N6fLkaJ2eKgV+NduC/g=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Wr0uuUuv0IjI0Mf2ygkRcwCiiKGsNHCSBtsfrkcEyvwsfYPJH0JMp7YAqlnv
e+afL4NGVyNOovuqjWWkTIirWfiUJe5SOJYzGcwCfUUlYGfVqTBrF/vELbEg
YkTAEKpNob3kOf5sg/0RlKlXRNbIgcqJLU+1yfhfIvcknS6PugQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 103968)
`pragma protect data_block
Ty4C3FB3YHnhH05jzXyX0kGmV3P3jK5WvcWEMkwc5o6JIttbnrWat0InnyIw
HDBq7ZSSAPLMuz1Aqa42nv7nV9gnlb7ZGDqNAY3KzlrhApzqtObLPaJTHd7s
EznsYRcipawpp/HyEwhpymim+0AFc8xf5uL44CsFUKMpPV5/fls3FzrHKbMN
I4i3datFXVJynydfWiTSVX/8RJBptDJOyra0wZFJJ4YZQE0t9ezetNekuPu5
2m5J/U1Tt+y33yWbCoOwIPtRNPKsm700UnO0SEF7sSXTIyCM7ncJTmyi0U+M
eXFhfhnoPxEwIefDeMn1pcOofYfyzByoZqmmSWR+Y+zsPIIh1ZdGtnBkTbXD
BS/H2hM82JqhkVNXpzu9nohu2fEhLiDnLUnn6+V+Tl5sPvVOPpz8lXVC8ZBo
2vhtF0Olb4UNx9Px06e7QfwX/HCh7EMVjpSWxYfsrbby6IIaccLcxX5jDToA
tUMG3ooNjIBY+ZPps1cS8cqhLy/6jcwtVUJRxQuRPUBsOc2jotHpKv5oUyz0
cGKBLbumQWghn6XsxfIszn4/JzwxzO+o47dfRBD5i/n0w6kcb6qOL2xng/U+
sBBSDDBJXTiwbylFYuBIr9+KWyxQNdyXa4KJV3+R9Af/BeMTrtrP13McHxZ3
3lC0hGrnv+V8R6Ra7qWMaRKfbqSNuasT4A8DkwmLZ+Nd+dDldiG0Qi/oGH55
5vePssSI9x6s2jwa5Cn89WahgH2AxVLjZrkJvuJxkrjvcbP16tLfiyYdmtfh
nOquxUUZGS8eWnGvMz0a/flzmbZp3QAwKchhSxuiDbuAzMz8XEbv8VBAARXj
9dLv+dUG2RaxPZHGOWkuyEmDGl1hQIjB5AsGX81Oc/qE35IOcesrstwk36r7
2eHJW9K1Iu6a7JWAwBxhtXv+dRdXVnxitz+mJdtbYI102KTxvCE2bxTxxRtN
TSzHCNmkRxff9HdhyaDHjY1eC3IskVvg3rspqXAKVZO35bSN3W9j8Z1054ia
6hp/4yGWlF9xnlJl0pF/XxZJ0IS1t7t3wFEodWwFwUFNivDvl/02VFxWVwBo
ydyfLtRfQBual8BAVF4QIR+hEFgU7Y1CCLuQim13ioP3ztjsIWO/HmzEAjUr
K18jzHszQk+Tt5voeSIklXHj38PFCA8bAsDEeQfBq9VY4HEv8273r/xb22VW
JjSOs9/jHmaYbZaEIQSGhsjulDqzl+FnF+28MoXtdjHesjIBMAmE/C+j17QB
29qtiqlPu19lcoGEEuAPALPw30bzIKDySA6VMrhAutK406JlAT350xV8ilIR
x1vcLevkRhzpKeT3XdtVASmNeffJNezUfYnmpz1G1Lsdanoiermxf77beAHn
UR5F956OU7FxffXctaQWqS/gcTOMrhXzDj00ewjLnlnGUkYqKvKjQyDzR6pr
YualneLFF+7CQPTBBeuIhTPYlpfDR6SRC1+gyqyhDWJgUiMI/aHAvTOw3V9P
kmAzOf6EuTDelsnRHKNFG0DB0+neMQhBuA74CQWaKt8d4zRZvk8k9HiTeI8L
C0T16Fnf1ATFsITASDasfmtL0qXAzr3eAS9/2Bi+zOx9BF1CrZloUG+GNJ2h
d3KtgrrbD9gb9TviaYtM7NaIXPiW7tIb48BpNYnVG089fcG5+SrRn+plLIHF
zBPasAC8z0ERB+7Zasnh+xb9RbzVY1EvqAWqyrQsF1Dmwog5NwbyyoMvJ76E
ykbRdWdrkCvLDY1IPY2m+9fb9H3kSMZOAaHLIhjP9dkbO0q7I0FiS+ep7Y4u
nDqJlXe/b+QpnxxMncESAFrAJs7/d99IDGWYy50H3CVcYeNyk+EAtG4CBeFs
gK2G5SOw/PxxT/kJ3z9n37CWzfcmLJDrRLNe4XVDnIWolF6a1MItClNnsrYc
/NausLXgb0tIkK9QB54Yfx+0h2WUgEs6BwCvrgCbGrMYKyiWZgI7ArPLUGwI
aWPMHZvFvpJVdOLCE3A1/EoGcNOsgwAEZW96soXXc2y6Xb7DEZ5LXIo38IPF
1FA4kuzI3HcOUw7mV+ecOK9z71Pu1XGWKNa/zga+sPnQX0m2xNwysjoGPxyi
LfwK96DUVeliUVRhp4IMGW7pTWn/Z9Ke0LAlBUWcBee5xc7/qnjYbgtIq0vV
tkTLhCaC2qfiMkK9PDaD8J+wy+9N1g6AzmFa/sgnhvSknxArH4U9xx4ZUG2u
t+Tkw9g730v9qERrY/uHEqtO3FM3L1A0LjvpCncqJOOsAZAxkFQRsOP78zIS
pluc+0r6m1/rl3z5uQFfdsZaCxkOzstmgpzkAxTpBGZJCanO+9d3w2RsedCm
AAxztzuLsYRnNuDoDHc5pf4fq+0scKI8J7t1M5Lg3QZW2EryBuiw50edsHGT
TogUMfHGK98mVup6o4Xl59Qx4PHB96pj83/Haq2123AYaFxBz64HJagc1qkY
Zu3UfRudxuS7s85umuAzVYyOUiFyrzM3XHuwSNbC91YHbC9HEExTSARPWw7u
Ukc0iVYHSRZkZ76vmuZRNEA1fN8sg9cUScrySCA+APf5JbJdeOdynQSbzWel
ChWzto01yDxLs3zT3D+zgkBYX9/c0u5sNIzaOJN7KIJcKI18fbu3pkbE1CyL
ruS9G20R+yQKfZO6TBJD1oRfnXeU47+FACOSoG49ycbw0y8jqN/yLuQ2g5+T
L1NBH73LK427nfsLXMV6xcyqz8uknohFnBZu8voE5soJ0+stU06WlblLvFol
5VWS5+QvYomwEye8quktMXXV6Qj+oh2K0fI4CSgWoalpUE1kTam9CV8LSyYB
8arEesDOJb7lah2xyvJUDUghd1BQ7oAkhygtUrdfhNCycFoQxJVOPNjA58Qx
tLV4zeB5fw8VJ2MxfeXMkdaciOt8j7lkBLDL4s11fa9zVRQGv1PKOJF3olls
FmAeebrltpHRptv77B3gPWo7yBmpIaymgp+Enp0JfM3XAwPJEfFDt/eazUvX
AY8CPooUHXC8p0iVjrfsrAamyAJ+R7bziA5oNTzeg20vSK26ob/YHnLE6FZo
IIkpvmYluDfNGQ5Z9ZO+qLmgzN7lSEvbXg0UyTJfUh6mf4MNLwNnO1bwEEqE
sH6lwjysyLuwzyLevdahbxIavFJd3jymLC8Fj5lzvSo1Bm1jvz7AzihKNwOA
GwJyP7eaoVQpRJnepyGPtUjeF0Tf1giaLtBnSf8uSFJTD29dv1VY1zO+wTi8
J7aQUPG/Nfj/DyqlepN/aDSsb8P1s1zXRzLxDVbkN+RRrU9QFEKvlC5sN50O
HiJG/NSzUsNtwEVFO5bd85UyFxLc3TqpA/ZJaHSyjHaovQHtr2ylDAcT+k9n
XqRhApj72ojqIhB4zv1IxOsTwcJq7oZuy2hwC6WjxeMxiInYakmaHV+rJmaU
6eldOMzEYWE+3TV2h4JbKE9eoK4UJvAWhU687SA6vjQY09wztxWmO5+mX4M6
mhk5dS0tEgRqNwmW0+LArZdTW/pVlbY5rTKAL/A61isYxw541a90THoxFs4H
6kQDe4FYCEAPJDfJRwJ7WclWX18LtaSgjB2HRknr7M64Ikjv1qe3cu2TUyAR
ktaR9PmF25w+WvsM0Rfhj4Z+b5igXGuYF8nMMGq0WSAcRFG3DB7xJJGfOLt9
ZHbvS4HwlCktKbhNNhWXApTXmh+tegb0lOwXI2OmDRSqpQq+Uvjy0hbn7FM2
Ra1bCfosihymGDDR1TFOQWtuaLFVuFeK5DjQbjaw2AarZvBl+uhb3rE2nXjX
UK2HvqdtuLDn0Rn6I2XKueMl4ADeK73J5s9zlTI2YwDYqdVt6i+BMNOxZeZ4
tnDoUazvME3ah53ULiF/nRQnbsd7lTNuF9Qox+rgWTYD3rvRYnuOq/Wzopu1
pHPMwN4xD78Ydydm+kcprwuCht87hc7zCXJXpDxPp2V5Y6vWzhvAP3YFXydf
GCLe5jafe0NOIGoPcsUnHKbbEbLjEcCnU+AXA82qjRzJEwf0G5tuyFD/RK0e
lybbKJhciMVwWeb7Wo+ZHWytOyle00BzFfFEgvTyt8odLVJ13wRHvGcc0Zal
z71LvQmyN6LpEwod6Fs921ew8zUlybfquLz3Ytrgs25StDSorJ1T5eHwgpSD
0cFUsXXJh6Evsuzpy7+8kxrdW59Z+0J3U5C5ZMwnrcQvpktHQICEssKVNTDI
Pwx2MpRK9DA/puGml5gZQiqG1c1aDWJA4PwNuZah73Ne7L+mvqipHEdRZrbM
bwOWVP+9aRRzOXTv9iPHyhgGAgFyFbMOV/OXAQCtBXT9xpzvT1Rykr38o2Iz
99nSAE3QySCjk8v3Thpwl51CNPRv4qLf8cz65Ip4CAcdyvF+Zf4bV35I8jPz
+Ji2yMuo6d882M09QSwMVXHav2Uc9F0P8ICV36Tmhyw68Qw/noG69dsUNZ8w
ad5Vm/XQM7Hu9WjTOSgf+NOcWSgixbuCnNwSag0uL7bi1LobAC14IEk0Jt2O
rzzJ6LDniNC/4d+0NKer8MWEE7Q5kjp4unqTU4bUvAqdAZvAowQQ6asbKpV7
DaEGBAyU2cctGX2GnqeA6QPueAGR0+lMJj2n0HSbq+PuXFm3EYBT1X5hH+Z/
D3ZHn8/sfIp9lauvg1fQZ7OdHlqJ/eH1PiI+jFFiTVn4IJsjgmHerma+EvVq
mYMbxHCELShXJFfSrQnc9q8yRnro6vlA7zXhn68YH1j13YWC8wBFOT2uNDpl
yw6H5OnJC428RQQz1pxmeBOsEq/RWWMqC+6w4HnMmM4Ho6bogWVuENZsuhlY
JZcsA+H/0MySYI6tCgBxqtVz+N7ULc3DVxCHBunzxaPtzxK/RaE8L4r2ur3y
98sIbXbYBtsYp5P1BB5W0wgXypW9iFj+FnuF6/bYWyFIkOMf6dPF23NLt7tD
kb4ebSDyI+8Zkzzgm/cJic9Wd1B5vzbj5xt56yTfYNj0KS8MEaV7Nlg8bfrL
ueRhPtHAEXxczk9fqFfGohdmmq0Q74/T8NA3B5t18FXHJpm3OrO7H3FE0CqT
Hty5ar/9lH60gjrvjW2pbVPX4MC2S3MgrTZXbUv0UK/hRZns1pe7tq2sgRWU
DQHHCBL0ZKteX+h3MZnWbgnZ/7k2jU359LOOgUSCvajnxlllBPj0kH/Y4Spt
36FhFJq2f/qMn7fm4UOMky6InhPmoM1C9yvM25cM/iJsDuEgnHBHyRWIIN+W
9G+UIY5nTMB/AnzwuSz2VSqCPdkRdBl6SgmufJTEQ+vHVUp5pvdQV2hmfEIp
CxB684YSIq2aGbxQrVMHz2nniaMvZHFSqUr3EHMAGJARlcVYzOxdEUIsNC7u
Ns1HPWISD/odYqSMJMxK/f/+d3nNiN5OBLVmHKoLGGnLuY/ejT8+5A9uTkFS
7z89x/7pdW+Rh37RFENv0044MFRe8gKLxYO+Fq+loRO9B+Yg8yWOxozGw/qv
PKY9lznRzl7SWmYSNyb2v1idN0BVmkus0/hk52X8TcuvI/ihiThuAGjZvADB
Ke+TMxB1V+eqz9YdMwZj5CBoqZF2ZdpWB73w2fiYZOiniJ0FiioMUuUAN/6V
LlQH2hgFRI2/IxNxwX2/9xT2w6OPq78Mz/WfWTblvwMzYKMtXIRZfGy9LO97
evuSXRlB9BkN+H0svQxUUysxPYkb4j3K5EQXwswcgymG0F9SLYCMVpZwfprJ
kz99nv/fmUbok5UoMvcE9gI5eBe58eQWfr53z9hIZ9iYEh7bHuON6x2CdaVH
GFu/DQ4BRCfg2Nkc5qgy8IYtjMF6y5ZxTsYsj1RHlg/8cfsLKpm47/UGIYv2
MLbdj35eO1xn2zcnV6emQq8HmEqm4f4hsiDhD5FavbqF+/Rk3yl86skmDRNP
WOL0MucqnntR7YrPY3q5XbcGhYFZ5lOn9wXZLXlujbMX6GLEbhA8/Io7bUps
e5FOnP8+012drFzLLgd/F+Dzyge2HKWKBq1CqKooxwC7LRDxiE6TG8nJgY5d
NaDIDPN1ABiihZyU+sc49oaaFeWF6WeDpnRlVB25njB4+t001iaXYzELxrQz
APawRRm8tWSiAKw62Xt5B5xd3js+ClrXx0BzQaRDKql3GMg6AnaLFVytoP2P
4qTmIl5S348GeKuEPNNJYfURqhYgiXYZXiROkk0Lmi4BugDRsHLb3G7uSZrU
OMTPxR0BhHpgBVwOwZoDeDPPrDmcjPHKnC1jwmy7g7vCbblzvej9dpEPs0jR
BQLkK0BXAfa5ZIWga2jEkEVVr6rXWCqmVcO1/LqrVto+mzwe+FczPcBaEEC8
ke5EdoCqJuufSMrVXovmMpQXVI5nbO17YUCIosyAlwDGLAdKwN0g78/2YG7d
miG5eaPnAvpuELmZIJjTVzGaxtxPo0tn/9cq1gKgJiqqgW6aHLqdWhNWn5Q9
ftPV7Eqo3pxv2ffOImVlWSu9UrO7gaubrLMMKCoOqip+18XhLlw/5fG224Um
VnfF//ZVc7jtr0d/V12CbQsth1yHKJ4RLnhhnPqE0Ub5Gk4Z1PdlNF2UGT6p
2apXgWtcH9/HxLlRfhD4MFbdgQQsJVczcy1DBJMkDPcPZEnKA9y1Rmj6Ujn2
cxx9k0cqOTBTT6oHGPOLZjA4hotbYl5ewseTkB/uBD0GXxmMaVi3LVX0SIyf
OHLE2jj5SkfT6TDTqmxUTSQeIh0sZ5+KWHdT+MVwZP2OeaFEkDDHLxnjH1ab
vl1KIlR+LojKHMtgQ6Bguu9BdQUQF0LrIFVJH0IZ/AYIcciOiQjj0fwyHUGA
NtmKozSiIylyAAubqZC2PmKuJ1JE60UU9pEHaPX70HrElCu7sygMFaGFtvn6
3zlaAWmjB+Sq3C0bl9Vp8ERKt80yq4+HVbi5RrApzwyTvpScZ/vhsSzXivxs
2uofU2/hXeqBfJivOIRGq5ZuFB9qOCAOoVjOfjUvR13HfJzrsD+RbEeKTThq
3PNJoDRddkIWnriiRGHbxRS6Isqvk+iIPC1bpdq8UWUiZTg82KoaWPHIQIVv
1aSCNB+BOtCJ1hiK26qhixEcV8iZG33LSlLU2Wbplh0tUTIZmEdeEI29n3JM
W72U+0GVGGEgv5f9WVhgQcRu5DTmydfELNSSj0LwE4WzjCVykqT1ALjV40SY
awRI4RKAYbrGcV7HiVWKHD96IuxsdMfGkc7baE6oNXbc3WGkMShRk2oDftSD
aKQizXcpau5tuXSSNLuQi4z3hv/Fqa/LYEiAC006bHIQ/j0VQOUHrtLRrgOy
72LnzImJcH5TdfVBwu5a6+y9rc6+t9Hi9NS7FtnGsmxWUSpJmhOLqsS2VQaC
e09Rwlb6Sd5/HdJ55tOxtmMT2JfmhlLjyk8og/H9RFYkzT7wKZ9n3K0Ceav7
PFr+dnccpJAfSjCEAym2xOft8wARK1DfZ1dBKxTFLxbYUjIdjG0LKpa2tZvD
uVcuw0cYd4959Qe4ThGQcljdlnion3pDJWQBGauSanvHiyXI6kSAM+13XTcS
ZzipVkaGvB4TWPz3arpzubxvy0ZiDtyQJHYdDkV/pjlz52qhd1NRKZdH1oJ5
tUq3Qr+6unEGzDuvUPFROWo9sWsbyLCreW1VYrdsdRsnbmAJzoor3pqKew39
0J2cwG+Jla9eZHIrHA61+FvYLUbkaeE8RwcDknp9bMSh3/11HRd+ZbaO7sLn
J5L/rb80yDlhLPSVBMwrzmhFM1uLuIVcVY9QLusUa+Gn84xoYCkp3wrQtp/l
Ekh8V64K2jcit++wXnh/QbMoKHpingPPHhcpqY/U4bXRmX16f0E03fO/QpNf
64nAHwMpJY3KEuoLIBCT3TzkwaZK7SPKOKDgHdJRmHuWoA0x0SAu6UYvZb2J
X7EU/mBNaFBlHapkhiDRXyeGMvEGUJnyOTAVuHe4T9+ncEP5SDIkEpKWSqHi
iEV6/pXSvZAtxI9C1lnkbKCxWc5mEWXPIVlR+MvEX67+QaT82/0TMsP7MFQq
QDPeY62TgJnrOQ6xCgXxApSQRXwepfNNzbBDorj9sx4D3nckRR49xt5BBduJ
KUffwMYMWT97VTRfKGRIYsSAClWgdcNobC6V/PgdjxMYYlpo9V1pvcGCp0Rz
I2zkIWMu4cWoODnxHYqtv8/tcDfQb5V00Al0PFwOcCcaOr5yf3vya3H+OTqt
TDtEhNNnpXudUYOLXfLf1zHcNSkEUbV26fxQ1OmrBUQuwOvdOVx8RPuREC1J
WhzpnkVbZyy7YH1ObnV12EAJQ4Mz1PlOgH5VHR4JNJuRuTkOSDK2viAVyqsR
8kuxLmLf55j9oTCNiJHE3DjVgoUznZXmz5WcmR4eYTcDLWFcLWgbVcu+Yo6r
lq217+X20io3AM80eBSITP7+mcjbKiRTOWo33aKF/7qGSlxGzk+Pfhd8BKEn
G7f06FLEJuVtuxzMJBtZPJZRhCdfOyLMXKKdomUnOJa0vovix5OfBjCJrdu0
ol4SLDbM9uw0AwrDNPJNvUV8fjjLxhkpMLD82otGnsKgYu1VBUjP5A0J/RdZ
QZ5+KPI3YTEUYwYvufrVveXHaMPnw1zlAEyNLbBAB2gFY7hv5cUqf1LW4G24
TWgWnpoYRJnkukwD8hjSirUsze1b1Cama8m9sKnRrqaKZtkq+n2jU1DixIWO
ekya8TPYLDxkGB1/oUZwlSbvoYrxkps1uDIpf5+98pnwXj2C37Kq9s867nhV
hUeCC49ybv1jCFj0zs2YDhmvphG8ny9fzfMr9CCezimCNbmO9YaiqCvW5Hrq
hRInc+PT59LG7MQSIQc2grvVSNSO4+ngRFUTNaD7Or7qA2Oitz+lvTwA5R3V
f7zxCgvnuH/hGt2YGfJdq9FzSDA7kPTBDyIsiL2LfJ7y9JjWDoaoRtpi6Xqd
GwFmaBFTxC5kEL7F8HSGJ+cMD1MTLflewVLYu0rnXrDJMg7B4aSTo0A++G6n
jjasI2fJod9X1eUoxU+OlpYlrfCq1fm7+6QWVD8uqg6LNaqYSUnGM/DufqEX
BJX9lvXhzNooqyUF1T0gJUaAQsVdBztNzKF+1qPc256G5gNU8+AS9nu9Vpz6
Ncr0Sj0cGlMTQ6wtkGlW17c4j+HrS2QwcxKWcwLhw6/CE08bhyMCRAsPe9/n
125oPW0ZYKjYjC676LDyCfM+ZsQe86KknT0oTFmdQRreKFxuNkMb46krHzml
uZRJxYuawIM+Bu/SyCeAVEDbQOQAlQwJTAq4SntWvE7TSl00cQAJRx3ZB6F7
GgCUAgIydEFlcpwd5jeLdm4I/Xq2cl0uBFc7ss8JuAIqE0tWGwC+rz832btq
5gAiE7IEjrDpe3I7ZChfmjpc8VlBr8fWVwOc+VzBmIUQ8XQv1r4/OFMgNBRJ
O3ng1bwbntUSTp9KO6Lkh6BBnGznJTjteucQ2+v33t67tGSabJbuYVao95eQ
2h+9J/1JOc+7mAjL3I2V9iD9FA6gPeNlUxdmyWSEHGToS8IIW5S6UPQM0tkH
qfpDwHx8Ryut2yB+8SKPc2LW0YJH77uSPsOhY7Pdvg1A1SqsfbcF0jJz+ubN
GL+bD86DwLcNqHLYzXV8lrGtBCQMBci8tvLwaSV3F1mkq4n0Nuy5gfX6nsYb
RYgk2OogykaWLW/ilt9XqTMFQFxs9zfZ9gUdgcbdm9IT0zMDTHWG2s3PR+K/
ctfGYI+P2DCEBmZIgluZhfevlGZ5AtBgoy68fN7LGSCjsCv22070mzFxElSu
7YHaBIpNFU1DCt4wfRUECjJZxCDejlRjdVcVX9qyHaNMtVYrB36mhdQIM14I
T1GhsSxrnoDmLFh4ugh5PYSFDTDghvgrv35jZ5QI6uAJ7VC7Ks2To7I/EER3
M30ztXQ78Ry6cbrtmWIdIDMjgSCVxfBmsPzHHGvHr3tk42trmqN5S+idGg8K
vozfMLJagYqlXQgzrZYCjIIKIbMqJwFxlsadffcH4BPwq1xwri0vCUb+Mpiu
6xPrv2Yysj+14vLsZmQ8x3KcMCjofRfUJ7TuSOOX9Jx+14CCgaRhPfH9LvRI
allzP8Ilxm6X5ZKOqH2VdSTpDw7xAL7HoVT3VEl16gynmELHJC9KXFMJjK3r
fVXemzHqC6JLTh1XPK6S2wr6SgvvptpUEeHyqcvsf1A0CD+DdTUL9z1eJaIU
r2JAHPH1Ntti24NBU+qecszaia9we7vGI66CXa3JI/VrtqrGpARtYP9zQLHK
TQRYiMutgXkL8K702QFkNyqMyxBlZeNScXmyzxyjQbMii3YtfxzgVP87HyLZ
uL5PRSfy+X7y8MTBv+1yO3znbvhexZbwBrHQpY8RbORZMc9ry8UBKNHYjQvT
qumphtkOzywKBQcYlrFeRzOuZgBWNyzzP4HqhCY5D3/X1pUC6YA05HdtRbkn
sC1MAKV4W9pvKlgHbCnkbcCEIdVfuPanyu4V8yefOx782ieTCmNPjdwQMIzI
EE3bPOGYOpI1WiqUa9xuBFS6MIIKt825qNyQKlzanMjOBrb9Y0hPNeVaCaI/
D5MWn0/0xFPFSBI9KRLUrPDm+GmcE8XlCs06idiGUnRsJaIJnQFPld8LOEeH
qWnHMWENbMxbkfGpiYkXNwyOZLOYafsKltlWVX8Mi410XRYg6gMgFy/dKh1H
/cZX6WQm+/drr5laE9Uq9XnFVMZvCyr0KL/qGJ80IWf6dRT3zxCTTwwnn3jX
TbX/lsMvWTw6tsPG/axWQ46jYW6S0RnpSgJ+zA/gezp87fvxNcn0RSTRFlaR
Wur1gtGtY4Bd3tPd/qfdPFutfPOdTzjw065Dc3FmDCqhtIGs1wBH6RZleqd0
bh7iaWRqSCAyRx3RDg8wRCK3ZwWe3k83+0tc0P7lzk6p6CviiF7/8Txs1Ce8
XkY6QsKdA9D0Imaxs1Wrs5eXA/Z4NqZBpzi6cVVJRfDIpHb688Mu5J6JbFxM
7urr4DJkTiT1NuAPBzOJyW3g4GAcKqX1GW6Fr+gW/y6yAIoT7ro42l11jqCb
H0kwgnbD6TBYJCHnhLiTNcohpA2JDMUpoyjwk9TrVO2jTgDCb797akUolLM5
oI6lQkmxSyBEBykBx+0sfZIVtqMq0W/r6MNRQXzuTutWMe5Os1r9zCZ2FCQV
8HQVUTVTiSrmp5IWm5+BZpRIzZtlFvNH5y2TrNao1EUwjvtTaXQ5owG/nI+u
kGUq+wnOsUWIZYY496cOYSNYxYgONhDeKY0apDBUlu7111/oXho9ckphFD9E
YAL7XVEMiyid83cjUfNFel9AGQIFziZsV9PgU6tkrjW236WPyvIrfM8x5IlT
VbhMAt/Mo1TZjEp+T58JEplk0m2HhB06Mcrgd6r79qoFW/EMyZ1zL8NmyuAI
p9mhuRMwWqioOGqiWRD+ikyHNj2uIynVPZGNCCET6aTspkbuICEfEgVL3/2y
cubzGe9p0RUpYlNBcz5QojDu7tGy9hh1C7gMcXc4jKdkli87sGSHiDHNeWY5
cXrtoqhEyu3cyevY5Dyc82MyLNzAnaDJZlMQBKb+mYeRlHU1eNbJOhYI37eQ
O/O62xsVIJEv+HRcvWGVDn6zXJEHUzeX0OOZ3itvW/4yEK10L94yx3zSGVvg
ShqicGKg94pWjDU6kGS1MrdQPmiva6YDkT9rJUV541fzBohjXqFHfGuOV7A7
513W/JrehM5+jC14RnfvbYc4ZgDDJMsUZkHcsJo27euBHj5LYCTCD8nHUsGJ
zyJnGJvnL1MRiSf+feR1PDoTytIRXNibA3lOdPqLKX36iPoAiTRkBf4C5RXm
YVlw85n9+aui0CBuppx/625TEf3/N6/lWLrYdAZX8JjtbIhFG0iHvaLTa7ye
r05aCU2Y7/LU1yPjA7tKpQnc4z25P08FtYm2/bra431Dsn4Ta0LsOXKPRUI8
74Xcs8/VThHvQPMiW8yuHVg8LIzUrgQSu9LJt8DLt7kZUuJYJU2rXp2D8DFT
DByiKtynhg8ybRLd7ae6q5hA0DJ5DvNGFGKHv9novXMZ9YPHpTVHjzd9dTMw
kQdAqyMeyluLQcbmct/2RFMxQlbOgglFEeLveU+OVMSSuknywVSfaoWwzjQE
cWrO07u4QSWf35Q57gUalLnB5x/kKPdQloHj4f/ejyyj8jcLa7Ub+yRjdKhC
K9MM63ZxPGSGBP3FI9AbFhnfr2IdIzzArG28quA2LOu7KSn/JmSTLyJ8YPen
KUM9zLiVv+6Ba3YqkUaZtJmDojubF+bFzf+MD0aRrr6iRQbmPKD0tz0Tlz4Z
w74omnRuUhfKyauYu306/kkwC6U2FtnbaGAfcRnwj6EFJokrX856gAd+yb//
LhBmhPPVIJDuIBm/4apJ9Koap6fwjILc2Y+5Aa42aLyVxop5iZfAtNVaUKcx
1J5eFLG6eKkWlb8eTw7EwY3RMBi36gRvwOfHvfk+rUuEzmmh0KLobFDfPQp2
kUg3/JN0q9k6+7viBkukhaJE9eWwDCgbh/gLZtazKJIkAmyDQiGtFBU9y2/V
4F8zyGySaOLcqK9lKEJSzDlD6BXT3Xb42WtvjWYCpVi2zrQMtjm7AQnlwF9s
QQGWBGG/tf1KrIrrRusqtK/2oFusESUp2UWum3vAre3Xu4+HmI7Ds5ZvhJuX
Ge+RaE6YVodJUvi1CEYjCLmAid1qimcFO4SBl+b+9CaWjSdS/UBvmmy4kzEy
jkuLnzaoEYMa4mmjKP6EXE55PKX4puAdgNjKvwn+ZUrlFhKG08vFsoJE3h20
F6tLjLBHFVIp/RnCHGJC8olwse8KYqATs4BXs8msmWBPJf8hOUZCgJhkw5eB
HS/20l/yxRvnKp6V/UeCnqekYhMu+oLcoJjyKasMCHE2tCrFyvS9Pxd9TSB7
7MF1LLTuUdI8qu53/JJhXOKNvEENJ1k5k1K2yHPWrrB90Rm/ZOerIbhldSHY
o1oaURKwZZi+eu2AzKBsbHqjt222ohui46nHD20vMahs5eFLk/cUY173By73
rDpsht0yyMqI55ARQVUixxnaZHm/Ai+nZMCLknAOSnUQl6wUaGgutUxfaclK
mZp78MYKB/iqD9L2LHKu4/8KrbY7l6tA4kjxEh43l5mABEAfcmIyJ0DXrI1V
KSov5hWXRH/17Vhgy0Mc0asx/yN/MMdcvq8cvhiYdx5MxpM8xCo5v6A2puk/
qsgcNN5ku/ynMWFF9YsJDRgz0tq/gQN5G4LLiuedCMxTaYfrBeT+xv/GogLR
U5lBuWFf7BESlvPObYVIQCdGsOLFHZn+twY8eIWn99n5dW3885lRyGj/Dmic
DX6pyPd2n5WnEdCc39yisUepFSMDwT8GkgMCvv+oqdo07GhZT03S9lbON3I3
6fv60t3lpZg7D9DGmPktwh/tIKcesJzqS45B2yFM9VY2HUfcwgcmjyi68DJF
I6dDRvlG6TUdmjl9wJJ9QK6/KxtKtfNV2pykoaI+nRZ5NVT24vg3Uyjqe465
U7Wb1eZFUQnc2MtY8DoxUftaMBNvxyFoLa8f5qOk4Ye4pncL5V7RSyMhyeXE
yrXMD0Tx8m4GkPde1Vrnl0lJOzk333NoULoKLR67loOOaoa1SNpEDi213ehc
J+omxzy/qJhmPEz3yzZZmmMjrBXPV9ZjRVN8zaEvSLd6ljuBX+GcZ432OePF
Rut0Rv2NRxhK6y5OcSqVG60EBL8A3zIbNkcpgX8rkv6Y5JoB3L0s8nAfvQYP
4DPIuK4kgbN2FcAU5rfANgLTiHrnh1ktE8erK+8dDEzvxTb09QZ7uoRpRBnb
8h5SUv30tPh9N8ZSMLu+Io9uvCFYxe9BeZwfsGRUAwbe/txxdH4EfIGCMLah
+Hsbi6WQUFlxKcNJZkyxmVaoQX++NtlSLaaw0gnn9dt5XcKBfQv8rnKdq3NS
iKkDuQqDiFP9NLCASNFMwOWhGnSbeVTsuinkAIh0+qW9mqYMlOetHtvfiytr
3JsrOz6QSRHaJ7pU0TQliBxHKO7M62TEKyUkra74vM6RO1h/OvWojQnXFCtW
gspDok5ADX17azqcV48OTP8ohlP8XbKU4NmGPNf5idIPZ4/4iBMS2/nyJpyc
vxlf57V5/eVMVrqmGkTV1Qt+s7N6ku7UX5KJmm8kKDs/5xR5iw8PdNXNT30z
+OOnokajpWEvAEQ8PDQbMe0MN9LH7CRed6lo6mkB40hTnoXFpASbhP4oWwJt
lV6Ax2V1OxHHj/4KA7891hmo6RhKGDZLY1kyya9FwfHcoxY1Y8c7jo6PpvrU
YtV+4TzNe87Xzn7xDxqlyaXD+KMedjGCcB4Yv3AiBW+0bXylUNfpCjxdxVJI
3ltk0qxUjpDgob6FV+vOOV2DuWsiU9LIk29CAom41SGxIl6EZ2otlEiEXJG2
tQf/57Puke0fN67zgNHgUgkNh+gSYfL+1VjEAS3FwvKEDDr/eKD2uKyWt5wr
xRPsTS7XjFY0h8HoizwnJ07OXYMttoXKFcoCuvLZdZuVIqcaQvN7FgSdi4ef
iKXtpn+/jbN1jxYJa5GOCgdIQsbesRKYDxeMaO7mOBvDGtUh5K7ovLY4UKhi
WcCI+wEufiWldziOFBdxCmNTAvd+qTjnNpH0yrmUpDBFMkdVPLaFxdkQt7oW
qBh8agYQTDGgpTut0XcNijViwDUmGFl+5Byb2E3lYYKTIkE2ewZpqe7GpXUF
mYB4cXADsJhc56LJRQxDTAc+vnBgkg4eyOIhAF2Vtqj9b4anoS5JKN4vytzL
OYwRp9L+XwUsOQDKUUXbSe7ybZx5oev+ev5nO8N8CfIdiNZ6eXYUsDukTLpD
0LFd/VkpQGl66LpkDe8QpwVJ8dGvPdN3oXM8BSUtYsTTTimmWc1CweQrVhR0
cbXFEri+F7EV5mh2Mh4t06a6nrWKamUTU+qZiFdV7BLUvOfYJBi5dsAtO9lM
UGIASnRikZ+KfSPbau+XUP/Ebo311IEYYUn6Y18KC/iwLov8pUmJ4T266bfR
/Gkc5SpEHPssqk8i2OseMjftvsJyxKat3x58VFZvfg/TFZOnj88msuLDr09y
xryeYjCh934wixqhQDBtz2hsuCTU9PD7C17ja/th9TWekQ1mJI/lyuf/BeX7
DPA3X12P2qe32muzjzIGt1K0AP+1eNmqdpHCR1ec+Q0zxZT0hHSByN3qkMc0
xEVnyVCh5RFVJl7rxBh9gTNTgdvRvX2RT+/AqTakc5pXMUPgthVj/PZH8js3
op5NPzzXDzA6vXCsscREDtskkL+/c4IGLU+gnQtqoXdRis6TO3072WYBUuHI
HmwYpufe5OzySCeENaf0HAoVCwhC32epdTJrr5ta4M/JpUGGs/v0sPR/YjBI
SXYtpUu/ClXGRra7oJQE/HArrlbCfLdzJCBvi/nnG9f6nUtPt+WUBOQ1HMPn
WnQMzQndETIfPOmnQ3Fc/0VNCyW4dp5RqXJraLbusQ4alCOMX75CZiQFDlWU
9ZfrVmAPvj6+YYRQbw96DmNDiqyK8sfjJIlkLbk09Qbu8LBjVM9LqrGfFPQf
9zKSElVfwopAWuYypCa/zPFdXywdY5l7nl9RrvAtVLR9PEX5RjNgS6kWJ2zz
Ja1tfzYax5B0kZnhXaNLo5vPXIhRngvwUPKfILLNE91MjWQLEUFymgz9wk2Y
0Rnv//EdlYbrKGNWjJpK/rqbhfnjGVM2BdY0s12gAPLeDFB/el+kSRdzt4MN
Ap0cM+EKuiLAGUkN88IEUjZ8XiJJhf5jnlLbqHhPqyO0XwkURY/LRsYbEE3S
I7qyWN10mkhGajWA1oa6+gwPoOkR+haORqC6PcUqLWb0B9SrXl4AcY+H/1vc
e5K4r/FZjWLTpmeTMgPSyr9B9U+xGrbHaLkK2MTbdtwEOIViRPAACDYkIblm
2mo9xB4n1sc+18WDOvaqgDYPQ5ukhlB5HLY+3KcZuQhcx/oKOCIp6UPzT6+f
c6T8DMEweZsGMOuZ1W9W059KSBgJfu0MqHs5htARGYaA60wu5lGDNK1cK6em
fwZ1+EAv1m/hsqo7zMPfM/qbNtApEJUoLa/Y8Y2WgiT7KNqrTNhrBDysca2h
xB05XrHAEYeLF7svkXG9YcnQRuKyjyTtY8LkKKvJj5/CSKxlzZw6sRe4p+VO
+oI1hgme40vV1Fz9h+dozeRkCNwk/LJ9Gse6Vxi2UfHoGG0F1nJ0rFWNTh7n
1y1/5SRF85zyGiVb+D3WgVYviVGWrJRbT/5NN3S2qjSYhZmBx/pQsAiuuE2P
mqooG1PpnWzB45emlXz9yAly7xpSNuMIRS6lu/of2W9oyB9c0tB2HWnj7MxY
hz9mzUn7+XEaPM5XAfI9iQnHtR/UwKVn7PGigRrlkGVbfZv+VIu9AlaUCg9I
+Ml3mr0sU5RfQW1Uk/k/FP/WZsuYlSotVIluaZpMFTy/ssSyVJcQqe716rqv
QeGf7JjySR52UMFEWHFN649M847MbvLatQnuZ+dReuUk76NyF4NeLmu6fJ27
6QwSnnCw4qXXKKMm4WkX/6LvSiu6pBjd/zjRVKv9+IoKAy9Z/NpdL1sWsTAy
UJsgfAWCJ/DXpFbbfJWXzrvJ5q+XQJRw4o/p89CD1TEXzjngPjaegXx/y3t2
PvImyrzr8zKRet8Gkt7jqpLhgSrtDSpEfP63WiS01K95rZcI3kO6Mw7f0Bso
Ek83r9Hh1jrEDdKFgr7WqW9Cs1R2enGRsAu7WZRFfIu/7Dg2kEeuUbUjz4aU
HLuGszZV+4tRFyflTxmFNnfd9IppFnOrwJzcRK6gC+iwrYjGPTnr15k7efY3
C+09J3i0axgMoIQra7Dp9VU9BfW7jf3/dRNhz/mweu+PQ/Y7Zgg4X21cWbOv
tBKtPwH1XSx7ujwrXHESHnZVSB3vZG87jc2Rh0gCB5Li4+dQd+P2v0uWde67
46+WXifACRyle4uCISz4FKfdD3y5HnXZ7nO0lgBRyOtpfzxQCVySU0Cm0i9r
QjqP66nVKGl5EG7BtBmc6RE2TjPi+6dAoSnl9Da6ii3QOxHt1zcEnBRYXiRv
apCKyuBRKbHg8MeAM/KLeyXFXzflngjWuGEPyi4N1DUguq81wicpne/Y+eWX
Lzh+SlF+eEnjPOladAxFd4HhNwUf8D3aVTXGQLwWscnEvUfZYlBz9RJRTDoR
qNUh+OIExtY963NMfdvZ/4gum0OpW1i6M64BQsFsW+YkntoCHhFhm/WMPb0U
b14GL36XR0mz609k2X56+bgcBtNaCnss9E3bTadERtTvttQ27+cU0f/S1V+h
7GBjZr6nZyFr56ckEXosVvdm3bYHjRDSytZQPhoYxPDw2USOspg8ZJntGiuQ
J14Q8hIyxzXLvZAVGzXPMCBlHftlhZfwBaSJeKiBMRE+r+mdRF9zjBIC3Fa+
eki5f4lfYEyOwu+ZHBT9WQfM2FTB1nC+HFSX9Drx/C8B2SjDETgqdjnF/TXM
y7qJ0S3XcXk4UA+0WC6ngLssP6tIeNqIHF5JcW+TrVJ/r3H22fkLXErUpW5L
vWrr7VhFxwpZz44Pxv6xtAUITJ8D8+dJb9h7TOs1Y1Tz4TdL4mE7bYDbD99x
HG9m8AXNQzd06F3At2dHPggX+4umZRObe6hXlc2e9VTMSfw2DS4/Ak5Zt/Z3
PhRV2/9XZj1MJ6t6oSvLdn46yBJOjy/dKq/IbFSqQ2OaSQMDU7k7taKWEPXw
u0hToPgFr7AsNC8aqG4XlTa3MFu7ZeWuuEgkX0VDI8Ux3FmzaG0D6Qmz3Xx0
Ti68Ubhd9gwjk8Ei2gjFceqosSSKeCADRy4Ut5EOPJ55EiBkDWBjmTf01HKy
7Z8z0D/8v93hbELy8+TXL6hDvMqmsBaxBGLtSD46s51kutf2OgTl/QmTuqfv
5U4Jcxd1s/rxAr6Bg5KA91DjCCdVXZ6Am1IWbxt/OZNqkFRG9RXR//TwX9BW
ma1/WlZdcbsotNmP5BjZo4JWVplHT0taOLxXX11G1NIR7tt0Yv0IG52R7cEm
Q7gaFI6u6kNuXW8qPXtPZOhzyUdWuQJSMHAkoGOsHecJ0v+r6pxCwyNJvbel
ffosKoyrVNS6b8FhIvyjUdT5sT3UdavY/i8qLF48PYXrrsNqcm20QAmwiQIP
q1wq5jT6bN5oLdLU8fcli3ck6E9EC7CUGdOEWSxhM1BhZ3wXYDKPy4wag2wi
Wc0d5qwNo9+3eo3kvn2szqDhT7Yh4hhUOKiwdNSaKYOiogeeicpO24Q0LLPg
tLQfQQgQbFbLFOumwuC+6bAemL3bu43jRCl4d1Pjr1s9MQx0/yM90Q0O9hNH
L7JIEkIMfdNKAiD3OXf6k820JT3UyFFmQGdiQdayiQDK9G7LPn93xkrViiZB
MNLo3Ejg74MGIulgRY0fmqIzXhzHnWnhAtjp60uMJ86SQoEez1GiZKZ1MNcg
JKkiGCaFUkHjGq25lFJCxVOCx8DO0SzSfv0sVexHqLoyTktJdnKNyLvbPRJc
SCzd9oZ9NkvU/WB3t5Zqmf6qE2NVfeAXxqpefbOPmdbwk74ojd2IEDRFe1HY
zPergpvBTRYqY1pksYMyA3Uao236vBMPv9M+xmvG1OcT7jyjgb9RdJw+JmVO
CLVP283ojFu2r+EdRqkTDlYuY4zWRhV4cPnBd++hVvtuPqZf0nps/OTtdTmi
avwmo16XGVYZzh4Dn6c5A2S9seqPdlp3vNwugNM3dvakSN/MwRJjabUw8QDM
Aj5fkAZ0fyKR9YSkwUkETleDtil/4ODKFBXAuPhgenQtMQAir3hab83XSWHc
0W3PqUSBn80CF0bLmt5znePG0Y/Dco+FWDAiE0pYMaxDl+P5Ybej5s/vuhw8
Fj0RrTai9ugSls4WiHe6C5ciVfsYFnsSOvHTHdQUe+vUyfXeLgp8I9pOYeMx
rhEg2JI5P5HZoarxSZMoCLXBJbr7zLRaXUgrP0g9sR553hlYYesY0PRvMvXq
8S0QlIZW6/XJnCXXIWDww45IRFjzblkg6kAjnfsDZ9ou5dsvRJRdJkXlw1gc
tjRchndPvCL19SB677SR/5Sh0lzqQzejtqt1qyekfycpdZ8sCPROHEFzUa1l
FcmXEH6r+SVSVX61h3v+ULFlN3kv8Ld+7TsA56Wa6iQm9AeHpYlX9EaDVOFO
cHcAuTwzdMLBEbo4T01+L+PrIXRhKF7RMUObHiuFAfR2B6DiYHf59naBCdi4
B5TEfaiCFjKoGqP+Q+rZ1Ekg56GX4YSa8rleupx9gVhJTJVE/0U8sjOjYPcX
GfiMVATIVM5bxTi7VThHMsqd7hBtmZKEeAGlEvVnzR23/XKLC85XAJudy2Ez
4YCBwetCBvZ43QN+QgvVJZsKcyRd15DQNv+fRew8zrIdJkxLlt+oLFvscuCv
rZI/ilw00MSXNxyj9T4EzgtSyvJYeMH5smXJgmP57RblZTVKjqHPbxJuhnsx
FsvBzHsfeu6l7cuI6+U4oulZUxiXqSzvaRuDHSbhLfymeTLAMTwJw1IopVUU
TEjnO9lu97mQx9EpN2oaa0VJhQ8YVus1LVK4wQFXYYj7lAJnGLqcICAZB9c8
0eMYLDU9n2GxxBruOlqT0QU3rSNGjcWCndybPg7yGgVRRGlMKuvAxZCYiSFx
P3xl3G3uNRcFad1cqxM8Z5O/Gcz50DwVvown9uLdK8ABlCGWaW6jxQpfOQ9Y
qzf8oTXVKrayCi22AJ0H0msyRIC+4aoD16sDD+Uf/CzTLnBNpX0TyRo5y+Yp
MJaVfJE7fRYcmV8WijfoI0pKWadxyS4308eCoTMObqcJJ0jVxSfwBnw8b7hL
1pT1aZvBQjfNLZWmJgIedvpM0ujiTuM3p7Ydh+3AkD0YJGLJWb+li/C1OixJ
oVue+mZytJ6nX0Dml9ibXxQ5BYo5UO200fcHVyTWeZBc0cPt39JT9avlf9VJ
qA3C7LktMXQ09eblUHDgDOLbApVTiR410066mRtGWjOD3HDhWJI4uSOYexey
U72+bpmua1CdmQCmFj8tS32BAjpy+2I1xvO2AsAyNgqt47OAZrEyUw+LdRWW
iCXBKaajWlsLXHrDu7Wwyx9mkOFAF8JqYIS4wD2cy2kiaZcQ1P9eZxH9wDHm
K0b6PqUwMybGO7Tn4CHNN/+DpDTYBgDcD+KtaiIRZvB16MpLVA42vB+jKk+H
QCq84oNnRGze/9rgBJIkZT3ZkomamGs2vM3XNU0yji6GkNS4X2NSEOrNgaX+
yxH+m71XMZrrWmY4sIwPeR7uJNkUVjb1gGIjGBuvsnayCbQ1ohSaojnI4XMf
wFRQRXJ9KDKXbM3mMi0awWVPXiBhyzGvIg8jcBMiVDohkVLfcEg7NtXB67z9
DS84ryqqQdePEuPrYbvvFcm11uW1abwVioa1DYJhNFxn4xPDVDI4wUOBWAI5
wAQzmdftINeDhlVOpiiK0b3OrvB+cEd9fORDqVfPs+pnuSrEaFgKiFfzSLE/
oT+/KTKDW11vzIK9kSFNv0fePeBKBD/JjQpvQYgQbJTlojIGbY71OOX6lbci
40HH2i7zh8j+t1LGKgWBq/2SNOekKJKUx2dovNW1n6eNKx2lJP/mA55NbVxs
jHVNXr7LsQEV6c/ljg9fhAyAHrwCDNJjbdMkeodRTBs92/x+8UM1mUSqtsPz
+LEOVHrXFZq7PcWct2URkbNJTlb/Q+uWosErkBVMpoH2auCgicTMbDRWcXEt
axUeur1iR7W8BLZxzVW7dzBjXCFZm6ht8NqhnNwZ1E6rxRwr5s8Xsx5sQGU2
4FdqeUrvPRdsl3IlD8CffsC4fnegJsVFU2RwC6u2jWXa2CVBeMZwRSqPaXLc
OUR/ucGn5Ep0jSRpE7Ifb11oFKgWXjMEMnPNtOGxoXzVzqelz8Sha8rYgGQ/
QFovsgCK/lo02p2jkyqFZsSzHONRTVhIrHuCQsTHM45H0ao6x1xKJUYOZZco
h1GPQV3s04HS3KBO+qBkioysqsb6mhupDqni+xdNRGPWWr7bgr5LdesxJKEr
GRKmGIvb4tk0iz3o4PnRRMDHRCrEKhwVSg2mBUpu75N5M+Yn9YHYEnvALGXq
E3gbCXkKjK9q+ytL7u2xB64EntWkqvg5uneyK/3E/leAdRU7oQGfvwi7Q27R
QmZjhws4YuyBS7z3IusZ+cgs/3/F7ZlpYT1c1kP4NpSh+aofJkCDvf0yUEFD
sVdqKqS9npGJv9W9cuy0HNier0UICRjRrJ8VFLjmImZTYT3GnZ2Is65iilm1
YPlgSv64UEPjZ0hK714KHKmkpU1bNspwZ57U+4HQ2yZ1Unyq2IwrCAEnCA7W
LymerYEYVEIDqGPBaVxPRfCdXzuFwlMHwaDQ7pITlBVMvhnpjKys2ZV+LXNZ
ZnRF0NCTipTeudE37L5tXMTJk2eLKRpwJ5f7CYlcal9UcK7+RpBo7UF+kvmh
fInh0PHNub5qUwyRzPzqFS7+i3Fhj1/c1al9rdqfdJnuR0Yl/fk2OYJSAZ3s
JO6ZAwdF6MOCzdRX5ovED2iEJi9Z9f4SUhtVUa4Di7rGOfXojwic3iAdM9wT
yoApYOul34M+oU69wQF7X58Rc1kSfpIwOw3U/uanK0UmC/KydRFRgawCZOvq
BcpXTCFEm81+K3MhUYVB1joxmfheNickj/87olobkQQor8TKOqDZnu3gx2s7
4Cklhc76cg5GNBvNOA7Veg26fH/f8KWXNdf7zAUpmEXpf5kI1ipYskyTWipO
zUXCmIyghlCc4CdG99NNoe8KP+UuHbqKVqAMM1k6vswu1ylnYbNU8K4h5uh7
InKQ3yO2D1tFHAgUnfAGauUiSieBQ7lD0CPSK1zMCSQP7N05bfRB4d4EoqQL
Ea5BmRpTm3xjAfh6QqiGSogiO/HNch+qRCadvlCPakSKZahrtWYr1kwugp2k
MYq/WSjvCNcPVR+CyynkcS/VXBvLtZmSTUr2bZZT6ldKFlCKmi9V3ZpVHIE7
zZpZOBU0VN11Lv3kUxRLxJLolx/nxvuvWF+qYd/wS0F/FPD3RjckmGK+7rsv
CbBm7Y22cS9c8mRX1dOh8LAWgUNNQnK85jKQOc/sDQtff22mRw3sHjEg+u/3
087hqcj7TBY1XCBZYe1WvpafegBmdLki7fsAa6m518gJCMZP8X+AidxiBLyL
xIib4doPugV89FKYQtFcdF/YSOew/MkzfHwZkTu+4pe36vl+XNJk4DJ6fNWB
dYTRzufWkpB8oN6dpvjX3OS+udmU/zXV74yHokanUtshYHUB/jPFCJw6O38E
+cBF5W6+3lPVlF19mK2ms15SfUIZipmDgVa/qSlkIzvE+Q7FqcN7gARIOKlg
JFtHAraf0SVT1C4+rGm7btEVxmCfomOoRPl+fnmMMhqv1zV/AXPDkzfFAc17
28Kqh44kcgtawjCwPDjZueVuPCnK9/DlhlD+XNS9NGdqpO04KLy0hFF4GKsr
bQfrIcKIx52xgCiOpxtsjFeAtBrnFvRSK5z8GqNava0H9Pu8ymtajVyGwPh4
bAVgesOvFZXIcclowGJyV3ARNb6K6pnafsMxBW0WqXW8E47VeQxB1DoMoUcr
hE1m/Z6vEaQCazzVyRtn/nbUUfUASeoiR5JY3SVWOR1PqBl6F6TRZgzilLDy
0JA/EHgeIlZf0VAuiOaLwxxYo8eJns+C5IiZe2wVxPyBhuxWsqBRONVjUSGu
gwNw7CxFXpH+Ivjth3R4YtEKSBsiAB5JBHIk3x4RhayGRA7HEK7EtIkrkCA1
inAMZavfCqkYWSlH5GtuMKU50491hUO5QhAOQ0+bj5jmZChQUYJbIRgILkbO
xCC0xZ5t7t9QYSktkiU6u0ji+jqpcw2uiNslswJ/Cqr4vCwAzkGJ40k0slK7
VPZBP/FqPvclnwEllbgeZTS26iAxIG0O3tTCi1DzbSbTzJ5zj4Lf5JQF+3ZX
wVclu2OyGMnUfhBwsjX3S743u3MUuDoAmx4WhjGGlG9wyFjb8l6nAhRolWxr
M9ivJRlx+2OAa5SYarfvi9v6iDa0ZYrtbcjrcxv3jFDkia0xmLMhHDghBrYN
Eh5jBesaBjsaINPWKFFdlPcExUJXs8UfV9A1fWKFrhcjj9WeFpQSyBz2wMK5
sBokdeqgM/IDyveW+1WjCv9ZtnMLcVHQQXty/zXeMSH0w/7iZyWawRHEh1j9
cnVwB0lyd2cFAEvtd0Gc21RCZRHGHOIO6zmuf5HYDV8Mrn1wX8Y+e3itPBr2
Pvx1iFLGysojDZ9cMVtMMgJRRnPbpqxUvZ2ZQjI9pNlMr6WFvmVSniqICL5g
ektE4h0gT0Q0RfA1KVXYaG2fOVsov4XOuvQ/aNN0wYZYn/mCfkfCg4+vV5In
8l3Hy4Ci8KO0aRIHwjZdf8S5ZzTw823zMceBL4VHob8wkn32WmaAZ+3PN8qr
ECt2GzL+P5yDUlD+mknh2xFpaTR+uoGAIMqqT8EM8r82xwoD8QEOqeSOIZm4
5pkIcwlWbl/L7RQZEIg95cbK2E2WXuCyN7IUT1MjueyzdHBUNoc9YlChJhqj
rinJSNThfFwKY50RFF9QhmY2NyzRxPNWRBlm1TUpaMcgC3yNEvecWA7X9vkj
C/xVXjHu3tHypKTJUohtnMQZX8OTDlaE7El7ZhBWUki8W4KfRjKH+aFOH9IZ
n251sTzEDhzjii8CMBgu2OFHZ2ZDlFBhYofnmcgg0eijAtR6jFtG5XGPqob0
WVtePuB9BapIWnlISvd9y7kRegPWfV6TVyhl7O6qJUfX6gQv0LaGQis39ZId
ZikG3piBQjia8ZU5TafcK1FR0fm1+nI99STEDZ197HOrcbNzWutVauK4BNdG
mMVeqUtIUsoVAI/WkfDNTTMqQqdeTlK0CJmwKfRWYBiLrTpWjzCxxW+QW378
kv4A2RBudpbwR0JrW61zpxR9qSMCKTWsVoJxhP+lY9ocD9rmyH9oepGjaECn
cV/RWtUAKf8LQMWN2Grho5oFkbCaV4ldd+pcmhvrNkZHv3bawUrKrK4yy9VK
g8br8ZXJfaPVOCaK/LIzzwYbrLdXB2i4abQk5sZu3gsHfHO6Ht1Flu/eGeH/
dszj7iEVcfD0kzK0a5CjkRViWcOYJqnPbtUfPrwH25tWEJQZB9DcGPaKs2sx
9oDwQ1sPa4gSYRqBcd2HqFv+YjLtjpQxpIEef1mZ4cwyWFTBqd4vmxbrE392
/6NHGQG+alqRdkgJPaLvU76E8YFlqj6VikNwAFnj264TE4OKAZnKIoI59n0Q
O4HxWZGgXswGLU9yhTiVxNq7t1+xSTg71/DvBPiMQNavzpTjtOenjh2V7WOD
GZU3oYa+AID/Z92yAY6DySc1QQZs2uk0wJUbGF5KV76jgHvi8Nmt2BBn1lif
t8zPwyu3THDwe+vXkc8Q3w84gJ/cyaNlpNX/22KmOaSb37UDr77Sxs22AT+x
hDhVH0KOzd/7PO7V/Lg4Dfh+J6NJcjlg0ZXK4SlWn46Z7UkDx0BN+lRwAh6z
e5AwRxuyUAHOjdpBYzVDTgwjixaHVcZt8syNVL6i/VKKEUjWOKWA15fQdGFZ
iehPiQ7cXI7xQyvkoT5Bt5t/CQnTdCvbhDk/EVh3q4aXfL6XVvUKkxAWXZnL
puidqX+ZYE2vdVA/TQQcJbR/oYGxU+FkXnTMjdAULzQKbH3bgWkxe7u04Wg/
mVPlHhtqdVKouZlhSmGli43ErndFhUOq/f4CC8hosoNaB14aEd4OvxsQQIYj
MMzBJoNIWFKoM37bqNDnneANuzTC6bjVpPdPeiHQGPjpztPaoYw4WQ/M6By2
yfSP05c9Lk58wtSDoQH4aI4+uuNGFu++bvbZ0nRT772tYsL7KVg47D3zlPnu
rlTD5BF9qawlT6lxksKJFAh7TDTrk0MINOaP1tddSBTe4eH3OfzSnGB+412G
wwT1bTa6enOe+YSxB9/CloQ9g9jraUn4GIWI3xwKX3T5bI0pUMUyeQGqgf//
sZCjIiY9WTv97JJbasfQuAKoUSLA9S95NSE+tvaI1EjuUYN9FEXIPrIfAG7B
iS7JZu+QxxID9MSWXrmsP/BkeT5bTDJnfHapHi1JbJ76FFCRLeihn/kB2W5B
ws549p89NAj6s9BAEp5HHktbndZ33JSi+NMkUYJucyAOlXQTrgcuwV3+faH3
4iQ9VwPweRoUqI8ID2niGLm1j914slNV33f0EEzIqXpvQ3WGs6SMBMEYXisJ
sZ/8XO/PnRZb/FbO3QZtYqNNR9sPmCouc6VNtWH3tCWACCwxTQzvdYnYCHrQ
HxG7erB+ZacU4w2vdrhgnJpTk3dfzfhUnWsuAMMJizTSVrnihzKskdUuUlfI
Wn9cNY5ZfyvS85E3N304lEhbLr86/8hsmuXXonfWiiY51XFTnUWy8QElcirx
rsVJxfv4uy60HLXggqsyhSP3OV66Lar/xyF2Xhv7D97HKfWsxznYC8Dl6LqT
JHtsgahJgIL8eKakkSBqt6VI8g8bLwsoefa0vP1jdTzpAVwfuxxwKxVrT3cs
8WGv/crLn5aDdWZYnaTabVytHASW86rc4boxwOCAriR2xlkYle4DEDMYgfYb
J23Hz7wrYXbGPErTl5HsR0y6lhTBXiBOOtyJT/GhYSm0AQuWo3ycH/9WagGq
LKYKyOlm+KSXbnxUUS4j+0bUtu/QxsF4r4o00YA+UaY2X+wlk9dzbt6wyEFu
Sk16YkoWoixaW02y/Htjgnshh/WkF1Dzr+UjAtYtDFXLCnIuwApFNDgyBoub
WteA+dbt6D23rH5EkcGlzaBJc2xxspCwzVUjygI4iThZO9hUFQiBDetd2eIf
y8dneIGQahcQaanJXVRV33JELSJAUfoZoJysfBPuDAG7wBPZXmdz5IUHJT/l
UhbcMHVzXCLdT2Liq1+coc3Q+vnezZst+kVVwTPoUQs68U1K6HLDyogFk3MN
Ci+PUkjih4Zz5XBcZb7jSEnC1qfWg872i/ij2SfLpI3LsuK2o6JjaGQ8OUB8
SEaAO+ZQaGNV9vnN4+eXzp6BuQOhETPVyel2o08ZitRVjUGAy8nhFGLFc4is
uVL4ET5X5LolN3q+q8QOtAdbmpFLDvHQe5gwfT+x8P6mJ+XwQUr/CgU/GZ+w
5djgtmJ3zajzYyWSG6O6Lc3wKbtvoTM8wYhQWApPZudlzE59AX6CHAWPK9fb
byzlIl00CQ1fWe7uAtEkCUxL0j/36OmGgDFR1YKXkqCParyOKeBmXjXRXr4y
dtVPlog2tzl3rtJk9UhMhEzBwalQkDTQuS3b3SiPFMylapHicV4exEBiUPPn
XMw28qZYxVemJB51VtAdFAyIo8agzy8rwQYsVUns21JK/B2bhgr3YcMznIo7
ze0ppdilqBGceJZrBW5Y8cn+UXjmDE21+wrR3ooq0H76ZQuFXe+e3HhiixAW
Y0kWR3AX1OukzZKFpQxxo10foC6nugodu98jps2jOTnnuBJWRNHWoF1uTIa4
ioupE1PU9OGEsYqTbpwUHhVbsjdw4/KZ+Go7+gBptWKWLXgj8TlP+J9q+KDe
08PGAUhG83/nzhKC/2HfpTOmy878G/BT7eDyfpbqHScr0DLfHZ9ik8qOn8Su
S9IMxTUZpNQzT/1w0svC+WxEHlx1+wb7hHaIzUzu4mFXLjNKUyOS1HrLgpUj
A7FCCxcD+0LRisBiuYa4uP+tyVQ1tquHoXspVf9IEuEnDYbdpKqXqRrDTHyv
dQPsXIfsa4JPZXmruEufheX2qfE7qoZurFKauH1+k8BeemCgTl9pkyAWZel5
mNCWyRfOZP+RKe7w/B2PDTys3jjztA8o0eWXoJ7+lWiyTdP3VsGy3s4nsKCa
TjCKSLsL+OOPgVmrd+NueGELLS9IQpzjjXOaRJ+6KO0UPnNV8jzuE1wT6fvx
QmhU3Zc+A4g/b+YWh51JDGzlzurZmr9nlcmupLUbK4TB2peQhMnEAhCsHdWB
Wg0VkEJN0dxgD/4MabXEe/tRkqFVO0MjojRLz10RjYeBohtk00yVvfIzlfxf
mQnzI0jHzSiSE+3TOlzS/HgBQcfvtWIdlsVMoeqOSex2jBlMbfMdzPn2C7ld
+F0Xr82dQ94TlPQR6pN0TYX+7Eaq9/d4UtAOFObVO48bIsazaALOBiJxygav
jkLrXFSEE29Zru2Tq9SD/gVF8owmlScQi6XGi4lnkrCuXj4ro7encPsmq7to
UAHihE9d5OOCajINdlD4Sfyc3/vQ0fI9eQnt3fPMcWGs8KfHvB2A9cEcwNI4
4hErGBHU2H/BA+LzhG+NKPPCzo4Fr8/dbJgpP33q0hWnHpjybxBgElGQ7v1r
um3Iwu8U2wce5nWIzh36S5zR4eptKDjFR+rszSTIsdyoIFu8zUifAgolyJjs
J8RCTgOchBsQ++/Wj6BLnp5mIU6v+wtIC4HQULbYdm47pXhx/6dHoSq9u1bH
/Q4cDW1vNvjhry0PtqrAddqsqxddEFzG+JPUCTCsS2nZJP5Iteq3QkrRVsMO
B9wU3f2tjmpJ4au5txsN5WH+3oHSSU5ln70n2LFG5U85d3qdJHC21P2ou3RB
ftHUznD1Jgw6JEOhl49gO2jDBNyi2QS6MRNn15Lq6ljO+lcBR3S6CjPMeP6s
vljkHaFQ6utV5h8UPDfyHy5v4YgX5IprzfC5RdJwoM4BdXqYjpljCBtxZfEZ
tKFdF++XeUQ38vSpCqCPOqCwJL5kbbuj69dsvbSMgykITZZbFSK87dm+Rx+O
Q0TGKPxy7Wa8bQKV2X8uUWXWZ3zbt28ynN5UFPVCdPFtph0/asO5Yhrhz+QZ
luHO3tnZjZXV7u2AxnZY8rXm1HZBnSFQqclZFJNU3q8KzV3N+2+qWIiA/4Fw
8VE7a0YIgi7aLQCXm+WQjhrZoLFpDPDHOADVoQIv24qmIeRSzECOw6wugkky
nZxEG0Dx7kwWFqXxhw6fcBjf6V47GG7XcLQ2B4AHgqAUCTJbJm1xl7qUmSVv
AAPJuVYznchx5OSr10W8f9jp5rdECrDFvHAcBjE/E1MDiM6jdekQ0rICG1jt
LhMrCgXLMMgEeaFDTuIVSe6BNjM5nl38v9hy2BiqLoGTvyFjZ/QZR6J6AZgf
mgBmel26BCuQ3aygOc1Kn1pZkjSABvK9H/sTujmkgBDE/ow6YU7mDSFSIuGo
eJeAgrOySjk6aUN+CEJSkwLc74pJIVl8Oi5BJbNuUTUz/lvEkwTAAYxmNmEj
xX1QcsWDfnb1ubSwyGyOv92q8srQgd8ih8zC6P1qtKuDpBNUYRA0lYHnNCgP
ljRSvjp2DwLel1VDYvshP2syIx2NlNOzc5DfgKvoRSF/mcuptAAZgDf+Vopa
DOE7S6x8cCfMWEIbrofoUmDaNvrcFMBeBiu80xm12NrAlxZSdKXV5aOE1H2B
z/SlZd02uiBK4VuT0pE3ucLWi49do+i7cizvR/q9kKB7cyJmoA88DkVJHdfd
Fc8lTs+rj/GdW9rWt5bjzgJkD2ykcefgab25eejREDMdP6uY1u91OzRWLfh3
Tu+Hw4tgaMWziCZwZDO0IvTVr6JzsoScMmmBc1bbRSOeGmzD8x9s9ym7Szzt
9m+tcWpVTd/oK7/ugbLAal6urYe30wQfdI13Ys9ZaJjDuX4rFUVzeNdSsonq
GOSd7II9WKlSGCZj2et98iX8Gk89U8R4rsZsCI/TzXxbaZaY4YuEewnLZ2f8
MeF2DzC5p7ok60QMCfTCum7oUqkk/r+US7oYS9ij88FDZbDTpIgQAdKnyNfg
7AYrvxaEngokhsGdQb0LwIja8vRmCABjQhA0WeLShrf83oYxEEGdYyWdEtd3
4yAoyAHGRNfK6y/OVyAo39xPXJeIqJ/hPKZ2WbCyKXrRYKED0dr1LKZK3GIv
e+MyD/GMgi6yZp59v7ZUlA81Ys51xEQ0EMtoXC56XecVccD2zj/CD17qSTu9
vV3sNxC1bkIMNqN5dtzLyZHOyW7ZL8kjCTw/5XehgxJ55/JLOCSgBB1na6bK
F4XGQEvji8fQQf2LAbq/QEDf5I11DFDgk2LlibTfFJLXr6Lzcwp/V89mBA3Z
2bYKqcdriss2MKtPzdybmhF1uM6fMgQtuVobTPKYd6TXUVdiJxZPgJpAJmyA
kWJy2Z6D6gvL99QUz2OxRatjniCew3Wcx4opohkLl0urdZem5z6Ai9hkmX8d
GlFnZu0hzac5FjvzovWDhYNkQxQPiXYAxXWJZlILzkPdjpRfBHWZUkUZE2Ko
nL/qbeWlSv4HYdrKkaYbAS3yZsT/B5OfOWHLkuPENi8FitND1Ztm5RsGQZGr
PiotP5JIqIR1NTqAtTPXgXRjh0O0O70DHefOPf8gCpeGPXxAaA/MACpYn7UO
X0tza7fYuv0inlo5Tj1/ADVwgfkTTn3kexX8y2g9pXkjOE+v0rr6XxgDzGOF
5AdvQmTAhFnbsy1+94KzEj/6DTSmFR/TXzUOmaFwd1L0w29tWqKtVNiBVeGH
gkbli9MidHvRyI6Yovt4N2u0kQW3w4s+GMFOkVj4zw59QX1B0I1gIIyYKkS/
4uVDD9SpPsbyRUYDpi4DY8In9P9fn64uM16kIhEmjWI9HYyJqnzgHEIlGnP6
vB1YwM5VJzopmmiEeFIvwd357y5rn1gYKILT6yFsWm2aYsyqZ2I1w6vAfL7E
awZdMZCRCBaiJTeaiRa+l27+vOReMO1NgxPdnuc4/pzNTyTihq5B8wjZC/zU
vMD28pX6oUc4V8+9ukTmIk4pP/blFamdAaN214NlZq/+DvWDq2b/buf/IK8n
77xUyLpV8/XSa7B4V7zE/7XFZtTpcwc5EATWNOd/m2N/Hz6HdKryZW4nXl9+
yNENakw70h6ht4c4bmG7cPZ9hC1T5G0gnNSJh43T9YUI9VYaWQNirzkonIyU
YXYqauWAQk3K1mzaNHXhxOztKNr8K1cfqdqHBBevYcCKWqK8hSv708reLm3n
H0gDsnns8OnXKCuUvmC4Io0gO27Dmo6ls40KcDUbSIIglaVYLjgbqz2gTcmw
bBfTWBi5xZjHBRmiM2h6tJqpb2Lhgt3dZPx3MDudqzMjkks0n2XV/vPXO/ct
KZCn3eYqySz007V4DF+qY5O79bhbe/GACV5Uro60q5qaZeclXOFkU4VVbxKd
oUtVlfV9nydcFsot/ClqXuIGMNuy3aMY7McQs4e9eSmxEb6PqiY+gQqtv9MK
pFLg2jiUt7V5HwQicobM/idFrzXuRx3oqVGEp1BYKaJDzpzLTnJHI1wQBX/J
HpHacVtaOo0o/grVax9DbJdUJoYbROUnFNbYGH7ac3WKRm3VB9JKBl6PG8JS
klucM7TYzl/JdGIQApM0K6sJG22/Tt7XNq3L+bOtc8bqe5IcGejum+ApvLv+
fElmXgEsZSjTq3zC4kaDP9mSBfyx+tH+SmVouuAE5ZQuFi0gN2T77VtQbP7N
lWA8Y4TvcKjInH4P8O32JB0qVMkGxHM/T/18zzr1ccXekRbXWPheRyufRCf3
hLj3M7St88DlWOEHuJc5rn6gZohCCJdxhIM1HQZZ4TOir+LogumIrOt+hCAi
zuhMliDuDphHtUpqwfeHzUMBwdvkB4WfQBgU6T64Dhjjl4gh2csPT0/8dKRG
Bhe1F9Iujh6KAHv3fLh0t5h6IZ0UHUxiMrXJ6+cBVkHtTdyT2fthdMD8x4Uu
Ya5ZbQOtksHVRxlebAVrIOzGw3IGPBKeE0Ek1gvMF0sKar5viDkr+lx86Dn0
xojfWRaSBygO7wxAzzZU17UqrvYq/z4vsgzUTkcNU3RRXf1J/sKq6crpr+fK
der3W2tGlj1hmnMbnWZdF2fH0BFgc1/SAalZkCRsdWvyu5rAAa067fxATf+I
Q4/yDHOGuzuTjAOCN5H/KaPhpvZCqpPrm0FvhsDd/ogH1pOYhl3m7feLuu+6
Ot2xgPwhqGOmLsUc9OgKX3NQnW+TedwUzC/K1vxWIQ3lJBipgFLkJEKMjMMn
lRJllKW5fLq752pjMSM9K69IfgZxm+eHt+Z7qP1eLnCf58mHJxvV2NZhxn4R
tC8bo5enjjY9zapyQXALlxfyyHXv1ivOMqAUzPmp3LY6ZHDHCN5I7oOz2gzC
c5Du3xxFRQbvdIpeChaQIy05+l7PxEiv/UdZxQX02VNcmHO8X5dfuZv3hP4y
lgH+O1RKOMcNiQlTgmxe/rNY8caTmxmp9353e+Z/P6ibh1YBGqNwQUd0iW10
RU8u+0sSYcdWlrnB3t/BbpU5/XsFfDNBpjWPAdY3kPzWYaGhSycJ5ilDDXl5
phwF52mUHVxs3Z6KEKIOzYqLi96kFMTKqJAdlG3SuX2vniHWx5KF8ZhbD3C0
kEmKFyh2hAa3VLXOUdSU16xrl2ezXEdS0KZSzFnMZLhtx3xOOz3qo8rCJI7e
Ljxa9lcRfYN8Xhs92uwv8fp7CjQW41y9UY3L1Cfk2lfhwY1I6zSd+eHlzE4o
XnFvjkWeRMmPqiKU7w0OkS06RI9yDYY9RxWZUTHIycf+mO/zi76JXK9O1Z3n
rg0UL83Y2TYx38QTzFbHSpqabNSXGnOfvIbtkkvf/OgyABHsLwJ2tHaDI1JO
29YprRGWf5+aGmGnUZwcuFlYlz6C5bUD8nK60G4MZEkGSPo0qbas22g4zcRV
J+Je0Am408Ab5owD0QZmprqSK+u/HI972ktmaTEAHDjaSBQgx/wumzOI3Phm
kR1R/UYxQ3oQSzCwuvW+mNNJKc50Y1X0k66RkaUtI2x8mQVg5e7GLVmsd+2L
8lyuYgax4PQbPV7U15VI6Vhc/qjceGEVwlxvgELv+xGSynmRUUbdVyHxpdZh
98BKOVbmJ/GXggDRM5Z4pu08YnIbxug/4lWMB9bGoPZBQ5DcLWfsK2B2lpjJ
s9AjW53QP9jfkUkxGlM3bR+UO6tmndfFZAJgje2N4gVKgf2tY4VB7tJAcuni
QxbAQPRoqQKUxuNDvccps01e8rFgnKUFzgUKT8+9/8VdTpKEkXxzkL6q9tOk
zA/bMHWcZs2HCVvkaX4yLUtZYZY4abXrrW91dshfk50JS68GG/6tSyFkdpV8
06yyzmdK/CfE+Jw5z16Hce1K4BrmV+YRUZJO+UjiHV0RFUDmrOUab1HNUo0g
DL1HWabti0Lv7cmehuUkrgpeJn7pZReL/ejImg9dUtEBaiO+vEWc+rYGcawe
YXLeYWSL1jvg5CiNXo6hGozyCuruNg0m/moHPobGnjxaejS5jXoLgRN9UkR1
M6Pqk56kBy2y5VUeHui5q2VyI1kDIvwFYyvkIsdhH30C2gogijy53fjfykUL
Ei9Ld3tSFyLT6j7EBkbOBShFYKZ3KGD1bF0ipAXQkTXclOLfTFHaSYSVnOl5
BRnyBrACG79jda4Y19rlPfcvrtJzOuZHk9alSLKY3xXnLbE7Nsvg5Qp+vOWZ
DKJtQm17ENW/H2LFuH0M/fiFOnEO0AKFLJJWAk7OpLk2fxRvbqgSduOfbDxj
+n43yQG3v3mzK2T7+0HftTDFbYoNEic0egl64bnXaa4LL+eQ6fiKydJ/AQXE
cM5cVifbvaIs/GvMj+A72kzZfjgBfyTB+0qs77migsfABDHxZFcAmDScGrgd
Qk/WJC1hq23ocCkXgiGFvFmlr4kTQBbDapoD9eWzoOjD5uMlpaT30tAPup47
U1jlxxYP+4Be2RVbVKbGP9418JkP2ASBaNu6YuUdE9ISfq9DW1aFHa9JpqKQ
3E7RBbITUrraSFQkA4MsA2A/Na4EXIsNUA6EEB9zR1a64dBhQCdQCwYqJCMP
aNvnvbWAS7f/EyyVkm+h1bGQ/V3mLjAvY9o6xOaqYyUuRsQD22h7mdFAMsAe
CMN9bK3/UtvJr/EYkEX00AnYFqCvsVYOFBROQfpDtxGQyp5GA3FTs8i8FfIZ
Im3IkQm4x1++UWaP79cYeXxyjBWMbCnrPPrm2d0kdSt9LzZ4DEXmBzSlvMmq
jVr8ctV01pIBL91JWFBPo9e6PexkNMyzo0JD0h76hlNAi7aRECq0uH7u81B9
o38z/mxADrKmFpwER9i5J4fCTHLUvybgEebrVqOchIh8eVKSevv50lXCHr1A
dV2FwHsual07yTYH2JLWC39WNZoGffAt7sbmDPccYjqlwi+z0K7oK0sabcK9
jvvIucKCwQM0U9YiSoPIOjxO3bMlQLrCMDCX1WIr8TDGE66SuvF8G2yLVkw8
CaYDZ6+eUoZxTDRKCHB1ashO70X4ipkofe4XbYrTp2yVVADN1s55BhmRVgub
xKFANT+TNO4dHQ01DFwYq4Rfnl/YPOLMYWaCx789aXlY48aOwtbLeb8BpFj4
YFnJfCs4Z2aWER4IH6Cv9iyZjlzOgvTYtIXZFnEhRzFiNs1/XnN0ImXxc+uj
OvbwQ5jkTjTu8n4YWHadXbx72og9nfb7FRutYRp4vBydTZxFG08UUUYGnXi7
aMJycbdXtqEBLPCesl0inYeVSWvrUKedhKAuJrW4eA/bmVyiwflztW+Q48+c
DxXS4ZmK8sxfo7iMiMES0rtRjK6fobHYjnFv1WQZ4QH1jcrtn3O4g9ht62Ya
GiTE8N5NoFXbLnhJ3Pr1Z5m1GV0dEQxufLDal9De9mBQB/an/6hq63QSf1HT
E5uSK1XDNB+WalO7/70bP6pKA1NESMdn5Klbi3h2l7pJ1EnovB5RwGjGYWrK
3awDpgur0mRwzMuC9WDJljIYV2m1ClVRf3Xd9uLkcD6RGKnv5FLhjR0ujTEs
qxoQUAwYxQyKRli5GA7IOS/ABtJfjvScxx7db5TopomP0fb8jLJYz3kpffVL
sI4NSOqrpvAqvo6DsoBD8adOC5an+AVhylTDce7kTihyvIq9oGOLWAJxLefB
GBECcLJHQRJPafhumLwNkVBJyouBORbDq5fQN6y6zlEQwG+2XKJMTs2hYEiG
23ay0HGAlBLJ4ww1MWOZaQmGR0lpFF0QspWvCK74AYJzb2GTobv1kQ2HASs/
4tHTAqwgmeZR6f7AHW/0uZfFTpliyK21ffNjdTS/rfzich38wGSiMNJ+h/fh
+cTWBjzwkQa+1Ace1aKxOIyL7Ah5araggsrnl2SfIqU+TvrVC9HVDV2cdRBN
7N3OfUb/epaaMJ1GZPqlDXtaUgGSBFux354zq8x9kgMvM6DdhZfiKTpurh7X
rhHC0SrEF9zkOFjSGA7BTGN/ldvo7nL+PK0Y2dhAUIDMBdtZuYlqvwq1KrVw
0aZrVOBGjLsv6OEX6wYRSGN5FvkPrd5OOybILMuof4Mr02obnz8qPSvtWJEi
Z+Vv4C/VlGsGafgB2EyYWoV+mvyeG2KcRTQM4GFqeY0sWOq1E5xz3JfBprSn
8nzCezuqN4p2N45u3AHBZHomh/d39BzVgB77myjPi7c1/VNwK+dByH4tjSnV
wBaw4EBasya/inU/X/1MXgtS/0i1JuciUhMy6YJdYZN8ouV+4XFKOpikIEuK
4IWPC9tegmxsIH4FjTP3AJuwUvQp+cHADfS2fOrqv8F/a46DBH+Ama+GCrQ8
WKrNzV6GuU5XGId1s2rQqyYzhepkmgTMiIiJPET+J6YSx7Bev8OTcwQFjg3J
4Vx60R446evmp+I2GhZ+xuvTHolBLlLmuOSX6aL3Jj1w+EPO+/XSISgawVX0
/H1KNCMACG4OB2Bw3XChoGgwAt9Xo1dRYd1qTiwG1cEm+iy8NDMCK53mTf1h
obtcnklrvGUkilEhlZuQNhph5fYsdrtERJRXHpPGEU8lAnJ3Z+fxeNu1XE2j
jvyiwAGqqC4wDaMuuCeNZ7MaG7yk7gkj+oI61sxxzA187+092//3UmO8Z1bk
QoX1EMMix/UFHxs+vyaN2QkjOMP2Fl2ZXiYGuNMjkD41O078yX7OK8eIp83W
XWSGyKNXFiHsyALtneuzDQOAfesT1iD/jH/xJjiIgTV2koh+KOl8o79SRiiS
WivtTBLwB6t3UkYbUv2eD8PwFLrAfZSDQxxjvdWhixSIi9vJubazRHozluY1
Ri6XqzOVEvwlepNYDzNsg1CF/WpaxOZWuGsMJJb+0E38s3hl5PAWRxeuuB7Z
Y5qCM508UdxpqEPDUEOWU/VlFpSA6naHTDKwE7/1pEmlGpcjhsuhQn/o9Aus
VRFhy/Kv4ufsAOj6nwTNM1rndRRQBpoxsB/voaadPpi0W6tWf3WTAptIKtRs
CDhYOKrm/bhjTMAzqusvIfwoJYjpP6jvYovHyK3GU0xEffbRoC/ozd60daib
TcSp7xn6VXc6tPR6jZBDXiKat2kNHuHApe0NUN6PJVasXALqlF6L45WwR0yS
Z8NZW2LqiYpidASevUGM0vafXehQ4K+YC04sFKk3zs20Jn3sDoQ6dzMSFLCE
ejRwSzjSYzNmecNECXBKf3oWqiiBdov6lQiq2XQUc1TK2gKrSKkGMcHlr0mM
Hyi8Gf4atEw0mNPXw75flj91RcOFskCIgL3jnD7yJccC2s3+4xGWqLm5BvkT
Kf4D2LNElzF7QCrKbprDpfKdQFDppt1aokgnoCHrj27ahLB2m+XKcQVAnWOe
Vahkm+gTAkoVSjenevG+S301Xd6DV6zW525bzjAIh3it1kKTywCP08Na3Zt/
WLZET8/p61q5IVMjbcTFfLerRa7Q9MqHqqXAPBts7lDHJXZPecbIsD+XBxMh
hI/PrUhN09waVZ6Mmja1+x9J+vaPxRnvFqdTQIyplFTKjLWuy70WoKv+ujo1
qMPl0XPWxRahzMhdFEWZGjVDoADScd12HCau5jI63RNG6ZfKq5nUKF4TquDO
i21J306/UOK4kkQKL5NsPXeAv/qkDFHxeRGi84R67L4zUotYmP3BEiQDTdQX
CHaVA/LYIj0jwymUC3zHH7o8b3MBoHDg6UT9S45DrPnGjoiSzuM/95UVWZia
QSZoaxX544ru/+exS1OlOqhspUcM91cwd0sAzRG0193w7kutcdKir/BHWnS0
yXnVnbszcacCaYze2BTz07SIKvsGngoE2gFqGt8aMt+ETWW/WJBBp9AX1jzi
rzPgqUfvJGDWK0b2caLCB0S8nQyqTtpciMC1GS873LpCSla90POpZJ3mGmE2
miCqnWEHLCTYdikF1sownivlgIRDDMZTrOkYoNnjN00vyE7P5BPEqx9mflPW
bxn9iZReWh+y4BurQhzr6hqLslU3f94CVKhAkp0ZwR+fzAuPvU60IkqwYKBd
PhmsFu+DVWFFml2bg4F6Aft7mNTXDlRgjehBEnn7j8ozLlqLhVr1omJF3tSx
7jffSU7F4tbYjiXK1etB5aee/GbzqtC6R4XtmtQHl2cxjYMEpJ5MBDg3+4vr
HaORwMASjc5e9pc4o9f1RS/w/Gwwae76NsMK32Cnzg6YdClOzs5QtVH0qM8q
45aQ8DP8FqXMHxapFUxyjhuKzxc84TvuIam3jXpW7zFf57TdGyaEGKh5PidG
oyQx/rY+uW0EkK6LkcoxhGOhE41FpFintMLS3HsT6+yrKog7sbe4VkbA5GYt
IyACATgJdUUQ2skOtaoloeedpwuIc1Ewj7P5lCXf7RFcOBXDbVaYS6Cbxd7c
zZ5ukzIS4Nk8Od56r1x5H4jjfSu8XuBX5+w62/zP/ETQrhgtjl7JAeQoPJrJ
h1HZVPpspOh9EBAW2DXMVjfHfehoZtMHXpsjMIBy+GkWq4lIKM4ESYa4LZNi
ih9bLM/s4bMI+5lOLg4M9gXpIw0G/T+r1MCEmF1JsjvJhB1/Z7nXO9+XV+Ty
bisuRrwTqF80y7ZGYgHDYqJINk8k02x1cTydLMtUTvxKcv6zocI9BDwFhNh6
mQHKA8dDR9qy32wHvp0FKjZWQLEp1XstRvFGzv+kru2OTwoO35rzCTmRb48I
nHZb9FcIVuOeSZ+AnotR8la3wyZyX6B9ms52h6c8w5sWys4xnx/5w5ghhXlD
x9WRgw+JYDuqPE0+SgaIxUPBBgfNPCx1yh+Cp6SVV7VYTP0rzeUbED/5Zpby
shZsBQIOBZgkBnUPGStqFeZmkMeIwooDJPdkKhqDZwCoaMRKORdFJtDOkrZx
ONHHjoKFwybY3QP5rq10UGFHwV/ggb82GbiEfbGOHfJnlaa3W91baHl8Bp2N
vk8Ksd3bYEoRdCEnsEVXEYqXtZMILrs/bxqcEPF8042sGb+G5NaTqoC6AJ26
0mwBNor945NHcSbxr+Zp+rT9Xnql0cbrsAuUQZZ8Vh54Dyaq2Zna9oqnubYO
wH9XX6FaG2OcNklA3oEecnRN89t+NIcJ3Q6fVnYXRo3jG/lrZiXniILvnWTj
bvpfc6ENTCt42oZAFwkiWAkplo8JCYPBhXjSF7qRJZfRBj4+PdOnitH5s7BI
32ULeEhX5XhD6jIpnUkPDpHmf2us7CPwz3Ve6xwbWs5h6tPPngJOavka8nlq
ZuahM8B8HsFFkMcdvs3GbMKFPNpDpRPuG1qCWLUeyx2PEzGNOCCL+b3WDqhK
vc76Op8DxEiHmRZSs9EzyyL9APUb0XGABc09iIPMpKLyZtMkUqxeH4p3WHNS
IKaTVNrQFCdwGvsddjvjhIlY1KBob/FHSRRfH4twvdzwZIe8m7PPET2bqABM
lb2zccU6OULQBu3GztbKso+Ctx7tSTkthLD5KzDyFZJdNBGkMML+ghtIl6JJ
kdh5DIisY6mHyLHlrxVaLvc+ZIWMbVNuGILISnI0gH2WFx87G5LaNnj/i3W8
n5BbC0vPimYu62ZPq4mxndy05z9Lev2rTu7iYs0IorGUfhydyKqtzusMALIB
b3zaA714xN2kZOK4th3NPNYHe0id1sVHbLOvRaIm2UuLrLJow1XCjuypzP+5
T4naM+0TRW4ZtFD5dowtV/2YTnWsA7dzeq3mNjkLhht9E3CBUi2QEARLkvVu
GyGS6QWICPxqeyX36E7q0sINxqk7Y06CJhe23VrmaYy1d5RZq8AwkleXzdxx
2hk6YLXFlotFXdezBpEU4F7mo3zkgGQAb+dDmDcBBGEc6k8RXdPH6qIwYuWg
jYiAIKpoB81Zxjg1EfEw53Bg/Rjij3C93OcE6d1FljBLRtB63igm+aj2bAr5
C0dhnyureiC/E/mUlqHEdivWy+zmJRQs074LYMAwdA+0kpuhSvyUPTGWfJr3
d7FLoz+hzHwmGA0V6I9jW9ClW2Rvz54i/jE8123aoJZa3sVj2JAWfs5tqh/Z
eMx+WHIAFob8P/LumvGnZFpiCg4awWG1QMexgBi8ds0lVwCOxd6T3G+1PeCO
hOgMGhapWD8/U4XE9f78WePb/zgUNjwPuwX73JyCUWPs4NkQx8EIQgzh9d4L
RCxhhdoRfAOzphrSwhSnQFQ6TAzn317suftVfuGNbGEp45ZmF65kp7gaY+0a
1DPNdyYbZhi5QHE2/LreTOtElGz3+n2b4qikEhBMDAVdvHapvzbrrBQAQL1o
bvBn6b9lljf+WRJhfUsMxq6hAABEBjXmpguROi8YDl3cjqvBURuCehUj+5xj
6i/4gDmQ/4NFjzNxjz3od+ynvLKMZNoAqXCTUyRqDDigyWhdF4zXFeF2d4Wa
p3emeoHEHUkD6sRvaL4G4rX0UbKiJZA2UnOzcP/nMJEC/8Mi8UTf95CIiouA
2Jfw9PHfd5kmRyxiSKKF3LJmaqwoFfrktzBgpmG0K8gwV7s2EaNkhlWDcOTT
ejFMA7yjUj7c8x1T0B+CN5V+6MwtzkV9W8Ik3xFS93phxRz3ar0Ee4rC5K79
wxEnBImkedcVlgZWpUv0Ma9azMuxSf+V0zdfUiF2Zy7xqCmqWAonnKS2IEIB
r7rXHyJxL5P0l6TAvz2Bt6odc3W6JqOa2ZN2cbocKOYxfz+o92tleWqrppn3
GKVd4utTNv0uq7vQRzlmS4raMOk6YdoLxycbsZKCcSzxQxe64pPq21d5suMG
IGv9Il4yRpPaKyhXpoaWqNnsTC6VnVzbsxCtRy6QpBF6emBi1g4vPJEGzAWe
O0juMKZu3sLjTi8CsYt3bHVzu1jnaMYi1RsnZgpkqbH/h9Qooe0j8/gpdC26
5S5PVkb5sR+9Wm/LxpKj8x1tuih/jfRlx00LOpK68Wo8eVeQxMRcStvXzT0D
XMLmo2hOwm3aJgMi/zHblu2KI25VEyLi4LljO0tNpz6uo3Fms6wPx+ltBhh6
5laJ0AhquqviJ9Q+koi3GXj681xCvpy1BIindDKeincFuleZKSaw5887EQNI
t/UQY9CTXxoZaxubG7Ob2w+Qa6hmAVSQpCnAzXHi2Te5dzVUq7Eux4RVLR7L
utXuu23m0+HwSPSGxxiEVB5jjrsMCd4dF4l+aRZBeLD2RVlgu8ngkAapfUD3
rRhAbVXKjcdQ6DpRZNUNAq7vw3eQT4MxBQ6/gQAYvYvQ/pfEeO7TOYLKvmv+
wX88LZ+8CGmr0nx7IIUKySS16dwiCkK71LgzYf3FMJFqtU4KALJ18S2j8/cq
JX5QiECvVIshK6H9s7zmtf6dSX2X9NQsYsKBMk2gVEpgPkBOri8COskzbiJ5
onpU/SOr3hAdfLLLzzV0Aa2xhC7EpywNqZpUSLdRohkcBT+lxCJeqfRHdYnO
PlGeelX+8E4IcITlqvGDNmAx51YZ2qVCzWWBBN3bFvso32j6PMbMqRu8PPA+
kljLUWRPTlff2v4LMo6poTGMTenfiZrWuUWOsVvWOa5FJxs1QVI1dGz+OAyS
l18tLaWuus6B7YU03wG232ceTQzaDR7KNvseZV9mOEsmk/oz3xmoda5xZpbh
s25f9H+3pQspyuLtz7UFQQUtsQ0siLvDduqaadnTvD+zjOvMx2ITPO1WFoB6
RyNuv0KAbXt4CKJWbYve6eOidg8z9d7mlsIZ9tTvvQyqMlkSQS7uxpFzUBfE
n4SkSp5DxYbEmIb8wcA1Y7MPx5kb1POGVm5pCqTSw08fTgaVWEpljgn2Ll4a
U5OB2H/o6aZxkGd597QI8UrFS3Nl0aLEDgwsWKZR/xxAxdW5YBlfBAnoFASj
KpGh/kYKNPvobN1GZU0KoaLX3M8QeptaE/P5ceXAj2MtQi2wbPbgdHEuxTk4
ETTZy+dgtdkRafafeNYtBw+s8zTvTiYY1T7FsQIjB42/j3Y+L5IJNirsmQH4
m5HlXNOfq8UlLU+nB0+ZEGJ0wfSpYtpc//GvVecFcAi58cfzkIT/g1vzgJWi
Ms+0lm0kSQ+b+ywT4w4uhUzucFXV1i0GrwUcAmvzugMKq1UEaI6hJJcMbDTu
xyIyLJZQeeSVMEnnHK9XrckEpFikIW9t4VbTZHIONej3dhbNWySMfsvyED8x
2fsFFkdxv1MAYy8AjazEn94mr/FXnwYbI8+O/CbAYuueHaLY5WHHnWaoTYf0
tkGcPMUMdSP5oNon7P5cdO9uP0tSSRYSfOmBD0me2yDzoTNkX2m/LJGh7VxV
v/kIjCK0+tu6/CYq58luQn4ucuZ1HkZ3jP2hDLHjjnl4iFZx8vL/12IiIr6X
uCGztn6DLfcvoW2KvJuVe2Zy1xrusIOAmB40hNQmWNPh1rUWpwh5+LGpgutO
hJTJhc3iHDorKPgN7I3j15KRrroyZVsDaMhK7R9u5rFE+cRmpXyddsfpqkDt
WpgapoAITndSLHY9MsBXnSyY+Cd8E1JVmml+DYDD087RBhqzFOiF+ycThNhz
g9WIVixJuC1PqR3pYlS1gtddc0Bf7KjNR2LKQ3UfB+3evNYIwRC85XPlOKny
qbR8YVHzuI9crMaItiHNS1zDmn/RM+UZRujcutztV9Sl41NIBNYqhww83zCT
NLJprwxz8/Q5VI8y9jcK5UjtsjDTTu4T4BJIEP7h6LUurb183TpqzVD5bQvU
qYbIkSjatCJv6lQkL0f6e+jfhvoXxHUrhaMWIYHbgv0B+cIqxwiy04PzPwyA
bMtwVXW8Zpgt57mlKLF/a/Es3PgJVNBHqhQmiM50Ap6CACXs7+ijN1sUZndH
QBZtIx1nt0wvkgsCfE4iRAllZMXVxN57hgV5lrJg7dDEjDr1Oz8vRyKz4PfR
6+/t4lHJt/KOiDDyIv1IFLk0DMc8UhKtLzavhHntiFxKmCGwCzE9pppcFn7W
M9hWzMkfTtqaYpEL8jA5zXyS7irwce03aShdNYf/M1iFA8OmV8VS+7/dWpP0
m4nShBK+LRLOrAUp8nkvbDhgQSqrDrpFEwJCS6+oUW8em+IiyS9WnNjJL7EU
biyeQSPKFjFbTzQbbI1pFH3Ps9wsED2/JpCXME9IWPAXdvebcY54/FzPMnzz
+kzJ7thUZzZwd+denKlT3YtKS42MkEYm9K3QCrlD8FS0TyhMBQN654darV2U
24GhYvtODaITVqnMdTFbYkecA2Gxjjp6y0tlZ1H8o5prHEIZ7kbsTnH6BETc
w0T0Dtp0c5AIkVBc700b/hk7UdBPRZFTTk/fe1nZ9YPKkXhEcKed+9kjVcCP
Bs+td8lmjS/5fHj/91vujDE7DyrU8EsEuHLZJS9DDxkq3VqodYt7YAEQpYnF
F10LPDNYn2UAib9FsW0Y5gXdYt2+YpVDLNDU5c6sskO2sJah47DSdcgnD1D5
WlErbTUcS2KmHtVTbkwjlzTEKFGbsnCgo/ZjUS9fEUthugxWtIBqTsA3g/M6
YIKyBHMJirXsmMZDPcAABNu/ofegQK5ieYXLlopcHyrdL3C5CaHbOuJd3dP8
BwCMDJknz61y1v3JiUYOdxkWI3DUyyqrIKI1gJBtpHBBj9OZwOwE8lRt2zzG
cwyHvwhxZd8GCKQcqQs51eFfoBP6IaqZdQ3+mik4zl0vwlOlnJ7Kjeyc6NBY
NtR7BemcdiJPYj2Qj9QnnQu/aNU+jliCoPwwXh/50Z638EV0uA6aZQdpMcw4
agx6rtuxvEh1suMNgSqItHLqdgrVUDB6LETRKqIBMQu3KVEVQYhSO2H6yAx0
JAmSwWbWN2etcUgk3T+rNPzfZMX1a4F402zn52UCr5t9N1VD7C1x8zsqB+XY
DBMlGWJgiRPsyhS65Pl7ONwc2vPl4rT7ywu4AwVBvKsfoB5ers0mOHpq//Fe
ND8Tg5fHP8NxqtQjenifRZEEHwZxhXfThOYInV7c0MYiJBwjOmb0koev7RES
zHS7mudXiTyM8lfizDJTKWW2e4+wLZfAtcI/aYoyOX+bTo4exbbd/E9VRSqL
jki4+4wRnQJFfHlBlrZSt9yTdQSbjN2uIK3jOI1oDBU/932L4gDYSdJPECWM
ahLQnq/iGBaW9hYobO2T51e8ZLdp7fc/4+qLphW9zoLIsktubi3nnaedaDBp
XntORbhpoa7kD/DLf8ezkPJovWirLdiOscDCapS3YSxCOlFbVAZBZHyH5Dw4
dnj1tS34+sjdbNDQnh32LF2jgBoIzfxpjCj7TWMMWuvvOmU2xIw+LemO9aX+
0ievYMPk1hPbKUQ73FbbPH3dx4iVtqLqu3sedN7hDr5DEoK2sQXs/EhYLS2E
eP1UPPSjz07Ge1CotQtPtKH/WoAlY0FrAkK0to7WlzC74awrJEEKNnaYgX4A
HYcsNfqv/10/oafVtwFbh2zKnG0Ou6TGXtdXJ6xQCHECMckpxmAEzBQsNHvn
Wh5aRCaczlYshpqaimrCisI8Yjl/zQdGtfngYffanAyz9nDpjv3IPr0HXJVG
UopmrFfrcwJS5eZCVLeDdP5/NxJOEceEYATwOSd2bCsHVMwgwjv6SIKG/v9D
WaoG0MO36RgASD2Du5/qX+QKsuu5fqMEhpZRvuiL8ai9KvsEDNUjh/3qrgLY
/EEvqkeDGVOkgvveNVT9HxOzj6NmwSu1HCTjlI3aMwXZ5TgcBW34GHKvp1gv
IoapC96RjtYblj8SqFOuO4CW1mzJ0Doe4gvSGnfyW4jvrQ7h0LO1qYj5Q8tY
X+wQg+UEH4oc3w1AStiYDg4Bq4yVdWmbNLuKMmXfD/u9NEUHAXpPyCe4a65T
GXRv0iI5LmgLwYsAZsjx/1MAWBTk+SQwoNfV8/HOqp95FaITo8k0ZQJFyCoe
MNaE4EVz5H/TWLTYF+6Qu7J2McsJ8zU/bWH5PXqWhYQip4661NlCiCgDGJln
ELwJGEshcCLdS/o3FYz9K8T3cp3X4iC2Z1L73LjHGZnpzqmfB0ZfPsNsiaZY
//BOHJZwsCzQG6/lMa1svve+DikOmVP7lwS5p2AT6j5dd7wZ/dpUdv9LCqe8
3K8zk/W/paez50yKl4n1KkJm4KJ8WRU/tKPOCoCfFF6lxTaBE1HOQ/2T3JbV
bFd8iTcpR1ocdGWQEAZSvH1KYqtEMyuMlSbBwfo7yFsWoTnYRq+P4cNRJRAe
6hmZ5WajbmO8sZUawwQS7NxBO3eNIDbBP7MjO/Vw6cQdAXThsyxRZkYQ6ANC
UZ3YBNdO7oSngfBb80JaL9jHeZLRtevAbVFkqvl9E9HVm8bjpIRKdqdjKPaT
pwbV8djVGEy835Hod83I+DutmIzeJ4qb6b+qAz0ReWamXK8Nb4Q4CwBBj6Rk
6ODI85U18wuvE5dRVREzqKjpR7S7udH59Klr6HY5gVa+IOL/07Q/FE3N8Uo9
V0ppQgVI1CI4F90GLZeXfteuNccR+3/J5L5SpYffCIRxRopcuDVZ30cv+4vN
dyiFju/JS+LJ8UH5nAlP75d38PSxvwsw2Ufb8qeiSjH1l3Qd10Zy76Z0xVAh
L1oWAzPHK6s/qB329108rFMKg+IH6BDhmd6yE46wfklPdFAX8d4wYQJwqx2a
23pCt8l4Li63Vovu78FQvbzy8TOcIuysWbgedFZHw461JolVQ2H0mjbBc8Rc
0/+86UeQm7ShIf86yt5Z2lVfyL3LUORLs4oWs9leVeIriHZN7WhYjm8HxhIJ
lrrfbtyRf4H5LN99r6G7wIO9KS20Ehi28zyy5NBxVGSeKdNcXs9yuCW2FKKS
OPlSb7CcEWjSBvzr18aRk+GsXkEq72XzYNCVddFHekGfXCJ/tqpa8Foh2/t1
jI0fyS1r818++Ut7sdqgeTIUpY77DHs+YoraqMoEp7d8ZClrFuKjYqoEP2gx
RfFNl0IOm5Iz7suihGyd3E+JGRGf1Ua2GVdqJSaR6G0US4OjPkJqzCwWkNCq
Lcu3yKYUKIEsgNVJolJNVpctb+A95wnmKI+Gx4ZAgsf6xl5HfmUeKsZtQodI
qx3m9uRxNpehmbQ7LT6OR1/wtJySEFmtaZl4ei1cjlu81knBtZ8Znlbla5zw
hz8P2qtjMFmrMUheMFTJniAb5lwevJmz4kq8FE4BBLXO3zshQo7FCGIHOLC8
PlasFiQ/dT6e7Wubq5Z6anKvCyjSNK7Lcn1lvhIlFIsBr5pB5bJPygcKdhVc
EHx5tKwsgz7S2r34fNT2JkrD9bUpS0OPuZzTzV+z9Bk/izL4aF5CfRxaRQW6
wP2St/6XRX7AyCWC0KCPXmIip9UjMbLRV0AUNBp5BTM2tTvX1gf/tilg6Q28
3RU8bNP3wrvjoathRPka0whFICicwheluuiH/K6K8BwRLlX1jWPAdKOh0ygj
RsCcM21lCN0q5FIqLNglp1pqiD3wDe2Bg6qMeKdyW9eWDsCnQiM1U94kkP4I
CMehVU3YZm1or3SN+APi7AbsGoMnR1JtaHWsdnKfkK/i8++1Ym2nD6Ik1cwV
nSUNa/Z/5pVJX5WsOjKHGWlFJcpuQlVPMZiy6L8thzuzPWHfUTVZN8nBbxQR
GOxYTtLfmUg5LIWvvJR8AJ8/LQrQGP2FUxhmyVbHakEahgk4I8imBeHzM+6k
y72t6WE8c5vVbiYZU3VY4FuU+YQ4rH3HLbjLyIVPB1vOcktiQcrG26QXRg7T
yUZJc7HF5gry3jpbSfKkKfVinNB09fL3Y+clsOWsgmtW3OWZrYhN6XMrdwzs
31E8XJ39qxYPmIBkmfLgr0LhwphJEONoysmTIf5HBDiomeeXXqrGmXQu/86d
SK/e0HzVVZOerlnDWkNCchfyRQuWbVc79yjgGDRU95vB7GXhO/76kTNYan7x
d9XTOm+y833YwGWAsdF6hMLrSRUpt3+oBPI/McU4FmfNfjQzRGYoXWb/58AZ
xVQzA8Z18aP4X9ys7NXSC2EYGL2Hwmi07z0jzXJL0Q2Tcs3h6XKNkzf2QNua
dT84l4RAF13L53R1ZDCJLTCrvq4RayRd3d61CNaeuYBI/Hpft2rTcaeDlS2X
zYo03JykSVg4K6dD6ShCOOMXcySXo+OEVVMYnKrBzF7PRTtGEdtJXMa5R4kE
eLNsmo7pcERvqHgV0Vz23J5X+eZhNg/BGhUj5ZqDq06OEDz7co52NYY14Tbf
OOmVaIPObL9VfSYwQvD2CmG1hv+bWJuQUEk883PK3hQGZ6xjJsAbRIFKooau
WM1DeDi7Y2NKSdka+FDiz/GKIK3q7y7MSn86lR5zmKRc1wwXs8sKvJ0D7Lvw
9BgvyK266JKdB+6YKtlMh1qDQ2pydmkdaH4JakRlpbCtamEelOxYY+zqlq+A
rdcBDO5Qz1jUeM97zz9k+n9DqSVdh8lBULRO7ACYL8tGvfsr2hjl0tLmiXGU
c/gZwdhXwOjVtIPebnOQre/61qkOZQNrFNUolfr9zKFFwv4zU7ottFDS+4sw
X9nHFtOxcPUjWpG41Q5NcFlFNSbVWryD5OG/qsOcdHxLILr6av/lqKU2yrjy
Pwvbc7G5BcfYg75kwhmEjiA60FsCCdy1/eDEGHDC3CDCnSyAAgTBS2Zx68U2
7MIkgzEvxc0I+sx7gw44KupWxA0A9sww4mJMQ3IBUbbP60v1YhIU0SE4NTkB
a65dBecy5sh+jB4awPZxLUpG9X8UHLCiWs5bPKhD75oGGhaXrpGvH1dRTNBs
eY+7fakl0tXUJIfHlLQ1UmMIS8Cd7CZli8oH2oraXHU3vSP5e8LVmOJGuQL7
KLkWQV6P8GqbNOAR5gPYCmOGK+wtBHuYUVH8o/q/b73P/gSnbxWBN/HMgbNz
I8yPKX/ouhjBPAy2ptAARgOCrhTfjGk3oUA76JyHrYIZ4cwAh1Oy3j/Zc1Vb
BtEmF3UlOblOKee1IV8ET5ppSqatglHmOQ0EIn8EQ8Xhg72O9O5uLxkKaMYJ
QOuNdPtaxr+5BQIAC5cb380tUA3QwL1SXE4KwBb194122x8hdYQePHFENcS9
CnbvWdKZz4gia+eDn3JItPOYMZ33HOd2g74s0SS4PrGzOinglvfJbgQrlDJa
ca3Mr+/EYW/TWBLCn1AQAPgLCyxdXioMR+ggmblGARfwBjpettZSqlsNrasF
XB0o4y+bdef4XFagS91Zm691p4W/Dv+UBu0zw5ec4lEAmxJMP1mAlMPSO7My
I6kH9h0uDP4KAG6k75rev6TUgOvd4LqAvrRMf4C736X63fXDiZ3gWRx9C0My
ybZwUCrMo4KEO8l5P3BkM5OM6NuX+lzPbWIqTc9uR+bYzaW8B23qyEX2e5g+
JhWio5+zcwdCKzeoIBZw4BJA8pgnWn6hx+WN2bzIMmc6Ouf8QSQ1Pq5MoWM3
jf9QTThHvElv9tFFEqnaXgZuROLfJ4SHJF2bkWoQPd+LuIVD4NH525B4XB9f
xsZe7rXr5e8/w6N9scNtXZHgV7IzZmm15FO3MQaZvSanxI29iuIPt8mq6s4+
i9wk3nbOo8NoYrsQBWov7Tv7L6kJ8hKnBitjjVJeB/wrs5tX/nLusXG5I+3f
EXVOorpQHscx5ha97rI4O091Lmaiu9zT869pb77ZciwSGwzXeU+RfqoKC+YM
AOXqjFStNhB0AY4CWhiSF3ZiU5Ifdh5XRjvM1ND+8c1D2IPJyGMwgHYilWE5
7EwBYTqZoZ3QoY/Vl7mpB3wLOpHoULunhC8pX9Isy7QWoLmvXYhw9WzWuN3Z
jBpCdJ8c4lKVq46177xAv2cQYk65IDl5LsoH/j04MgjNpyX10oVjh7DcXe7L
+rfALWdhV3X17Uolk3GP0hDrG2ZyKSqpETTqMokRsEgivsdwjFF5wH+dTHl9
wKdA2mFDlDZczxoRWBOsmdCbqTihrivZ5cH7Pj4YSI2xWciQWK5QYa/UO93s
1Fr1qYuqy/K+e0UBJJiskv4hna0C4GHKRxy7ctaZ9oDbKaBWcUfx4hZf1Kf/
6kj3llzL4FaAk8mRR30oO/vLIRzWeDUCjrhR+RrLoRJjnCxEhljdebhhVx1E
1ci0byOooDT0jJM8I1H2LPxvDP+ke70ZfHOOQ51X3wvn3FTsRjaCWGXEDS80
eY8vK6fvD1Gat73ejsLz8zgQijRHGsNATwjRZ3V0JW6odAq/WXXoNQjQUuKk
2V4D5l0YDfrVeTTkyQUdBWV4HIVw9eTr/nzYnJVkpbZGL8AbAeXEgNq5FtfM
47oGIkqMbzlvAVfOeaFZ9t2J9xDLtyw1b9xOjcB5YGp1hitxEij441IbebIg
BxB1Ittmkzs9aTecKZHHP62cb/lZ4EypiS35zuC/3o5qwkwSrHK0l7KM9bs9
K0/5sfXBgjtA0BzvSeSrF4o/hTkW6FC5oXLQULRWRitinpspkJ62ww+nEdDt
AkW/RYk7uZBHVsgBm3hC1U8gWn0P448sGrQ751W7BmX6kyyxJKCqvZ7F6VuY
/XAn7kMLFfu4P46bEkXmY76nQI2NEjPmxljY1w/92XhCmarIHL93lthPgOub
8qiSO9VPonE3B/Y3P8uwkBf9P69jH01ww4RbQQWr2x9p0jh1PAgMT9AI6UNP
Z5giBbgorfcbEiNYIp5tW3RLaTsvR19QKd47C2jZ7+1xrQfFUMznR1uJk5E9
yo3dIV6qsDBRvNVjr95uVR5AC23NkQfHNBVuJlqAPfNiY2jbEbHJZlg6jtqn
wVmolGNlz9b4uuznb7beGPmIc6fXnEC7u2vx4GkorDxQ6psTPl7v0Cl04cbe
Y1Yskerp/el9n7HV+gc9Y24pKFpyNZYD7KUF8BPAnsn3Vl2YZ6jbQkpprJBA
/dQixV8rPkl53l9052UKIAFzVjoRAaQ9vBi81HdGWj63ZwWKD/IcU85XHUfu
8wtuh0p0c2kKLswmirphZg22aYaV/Mmn0htjlkT9kmYC6Q2rwoj1nV28swek
IUbIAJhmYgbrUENao4RMwxAVMEcGFQA+8JKTb5qEh7uLPhOjUb5X1eP30HGL
YoRjIQaKkfBuGZNK5iOsYPA5pRPR3VoYrRhBz4asm3ldkxzupWoTmHDiVccq
slxZLLMxvPNZFtq4x5DytmZj6NLDl6nSK1AoZNwzMJM6I3ESqZTepy2NlVWI
ov+hONg827N5c5MEOYM9d0QKQawBf+vNCgAeMExky7zB6lFENYfpJRI5CxPe
AAH/4fjHrIgq3ouFmrR3MW0CrtDOFBys5qTUAwLoTvpuI7chMYO/u1+grfMA
G5ZSvFOPyDs3pDIp7fBpqQYDOUHRDGoHzD2dKWF2q24YCbocG3ip6X8vhg2s
x4Sm6AjLb07dVKadJlN/auvifQGR0laMzJJdDwUqgUjy0900Ere6Jvw2xn9D
7jtimO4Subw7Urcjf0Iah2to7XHUJ6DzCs+O4tb4fhiGwNIaFW2zs5Qifrc/
9BTj+2mZZZEJJvyfuQIZXCsOXTdPNUureDQSVpzg6mEpSPMuGUe9cZa8koJJ
SPRMSetsAvZVs0cOQmX2LFl0AtinAIa4+m/HcgUfaDqYGX4WMQ1l7QGyhcU7
inIVyQ/mkk0wdVWXWvgq0hp4DMGTedD7OuSQ8lh+j4tDVm5i8k11Aw2iJlq1
jHHDXDm8FUm3x8aSHsuKqli19QWXsje/8NVm9dwy+QrFZIJ8jSfWF+A52kvd
A8L0ZAQoGUQ6ptGk88XWPnnaAX8rwtwZd2uNiAZ7XL8odUOP/6VBov56zOYi
D+r0c9CIvRrAVRu+ZIq/AYM+dmgkPr8I9AsrBDZkyRNlk/n0COwV757lDNhu
8Em8Au15aRHUf0shGNEtNM3JDUvIQzVOxLuYjql+T2B5nq0jvqeAfr+IpECd
u3BDQPVRmDsu3yWiekMHI5AD/SMj4WMhT5IQv7g7kQNh5bRwxbmFaXoPjnLe
mnQsnT9K6L6QpF3g+BvaVjAY5Iz7PcivR+x5a7VaT7i9LKbt6Qbty592EmEo
E4tpNzbvZiknlyU2wwPZek1y02KPIREMI6GDfT+MJ4RU3ocmDLA3F98snC9M
fMSCo1i94aaQPSx9tjkS23ejlOxUvS6v59RFjfIJwYxjOvDAxOfByF8TEqqF
VJYxUDHrSEtrrGr9u4s69tILAW5MGRD3aCxJqfMlhWCyY/DPlZZkp+/0S4Lm
etYeAt4gZhlbl6jV6vC4N61jXC9kqYsTE9sUJBSfiUBkAQQoPSu16FAQ0uAX
3v87r3m+1MWx4ylc8wHUD7XMSmkARfFIyh/LO1kycus6maICBx991KuvN67F
57BtShFpLFC6ZaaAJCpNFsXxzrY3mb9fm4Qf7SgQ93AJKY3kd9Wcdw1fgJGg
JVHk1nvinR8u7VumAjm2y4096f5DjnMo9IhotZikUQ5JYYPSfDDTvIfOhGkm
2o1TFVIOW2DCLh6kkU5D2P30FNAMUESKpUnU63TIarrpUab4LNUEJY/BIxWv
JcQgmY8CPGSjhYgHIeYCvaUFwjXpOb+XBO9eYb4Jm25ylMvhqnU/4kBuE9bx
pR+yfLaZI3IWQGSEjATpT+81zKZupBy+iPKKXhx7hgCkEN6nDuHfLRh/jSMz
nT9ANWfJd+2tEqegcGxYcf0eJq1OyqVeL74vfTf6V0EAp1m57l1rCuzsN54H
G0VWNMXs5tZl5r00pvBOIAPPNKuFO0HPjM9uQahsFgqbaJaz4qHh81KmS6R3
OyMbLcxjqWHgvrqstws9O+6GCsBrUSauyIDyE1dCmn+obkOsGfmxXW3bcpSA
w2jD5AL/OhknzoT3tuPh9onIXTUjS8Bij4s9lukRSK9FVq4bkuWYl85jNMF6
W8vu+UnPFNlpR9lR0DO5pK1nbO66pw8kNsm197D7bj00sG5uXhtAqdByaATF
NBiBR+Yoov+yyEb4GRCD7ar+5WrJXbTdIZpurxt/HscaJJH0Egy1dwkh8SnW
GwQ6crptE2ECGu0XLjGrsGKHko1w21uuNjUg3r1HJGkwDG7WnFjnGgn3ZHkN
l9bkfv0sB0fU211E31o6XyJhsRiXt3jBwf6hjCxyhadGp+HcohJ5JQK1MMtr
1JSN83LpfQ6r6A2X2Xy/WhvdNcMvOdE5YKOXAVa6HmS4kd59NwMDPoRI/YpM
LBSR/9B+TIW3Gq9Tlmdn1go8ZgmaQTtbAc8jSvkxtQ7+ChuGPqlVWnm0J18S
6R2lgFuCG6ILPf9XPOkpWMi5ef9CVQHkx9bjznUy7BnsFNHXUKf6HbbI4RYe
vi8rRtqQQ+BgG4XtKIbSxCkWFpupqMR0muihgC6tCQ8x98rfo2xTN7Ux41Fd
S6m4geN6QprySsqR+mSBOLDGbzqgSUDVr6yMN4vLqZjg3rP4w0kuQS8UtCyb
YwzceMTVCjI3qo8iY/F3FqZSDpm6XYw880y+gtVwrZKHHMutMRWTf/onIaWh
X1A67M8EJqbMGIAIUeYUpyjTjB8ioPgfJZBlKNPeGXrZaVgOVgI4S2ARH9mk
M6zB6GKZ0MGgS8qGspS2ezRKyg/N0FeGaRynweF9SyLcOVCzK4oEWnt+CJBq
KzlqcATH1nkcoZYPUQi2dD4NEUoBousiPl+DjEOFJbdCouPjy4U45RLLwIWP
NjsFyjvueXOBbbiOOM8PSWzPuQ202+0Um+3TRF+ndFDIXmy+kca/dK4EBI2W
dBahbq4mX2W4ZEvpu5AXbzk9MNWrZ1QLJRmwrBhBhbqIf1vv4zzNTygqvhSI
jNY/QhiKH3EaLybff6xoXFIG+vLPf7UiswkFDDPJDE3vVj33FGqsrVSipxgk
++d90WgJKu4cmEzafA7041AXlVfVWTeiINtPSINIK1HXMzvyH2Bko89bMH9h
B6TMYeB93CYNkR+3WFL/GnGttBbzv4Ogdhmk6nRXPxAV19OPaErZyy8m/oLp
sraswz7cXc/z/Gg0eQfsrAw8teHzOayJcMB5KV4jssP40ZB7+uuxIlTQomnW
VrNrUu0I1M2ivZjIXidefk6VtysnPFVDXJzbTPHmtS9rWsETgVnEkJ4P1bUH
9SlLYz8wDROpC5SolG0meTH5CsLW8o/nE8QsXwagWDZtSbJgoUkV9yiG30DV
cDeHG5xEabhBs7VNaQguc9cP88zkC+VjSN5SLGGC5O3aZIZ2dzsJwa7Hoa18
6CoAc8t3sclf41Ga0vKVI9l5U3VRk4a7p5iIg6aMmYhKAFinAFna2/WFmc+G
IcUCV3Do7hIbskeSyvJuUNuAdCWiWVDSJbBJ8yWroOol/kK4y0kUIPa+6xcu
NfxLXtX1eRYzh6wDEKzMQyyFXYCZ5mCh4cKojeLbpTv4ul5RHV/TuIRGczkT
cvjHk4FDKOeEbQgTkM4gH7sakPlyFywuttGGS3SnKkV5TN3tXPds+nVI89tx
IqJ7ZpGHTqoaD1tuB2wOJThV9F59KlDyGRKPiW4DJ9fR7D4hqRx1F1KnlHLi
cpXoplaJkOva9UrB9IOcMzyxjoy7xFABevoyPV7wXE52osY8fuX0Xp7cAv1s
d21uyrU+yzDkys5rcPlSx5i8HJYbVfIKfW/Amu3IzWOo/OxLZOGtQtZAhcC0
B180KbEt+VgR0jQZMJ1jbo2mcMMPnoRY02r+iuGOKGOpRSw9/iPfKNgfD0j7
oATagFIvhTdyZxvZIy7jzNlhgIwHGE/9kscyo0hTFwQ4Mc69fzdaoWRVD30H
15dQpUsd9C7mHiqGkPVZqOm5bGrMA6XrRY/XHs4itF3yMRR9yKBNk//dRPA3
iGbXR3wOn3z9XCiocre/CcVyha8oZWTLvYgL5DB7knuQnTMmtGCZEQzJfzDh
gjXr+vSBLobLDSzo79dQx8hBItPoj9d06erGnhXhHN5KazEAfcraaYJzKNbp
Ss8wc0waoAJoiuxSndXsaRN+3WJOx7mjVaMeSkS7wZ9jEidBeq1u3Khpg/Zy
23kYjc5GDOqDER1RhCi/e0H6ewsyN8C+V1m+Hek54tgVP4HS7G+O1IOqQVwL
NNEPuSXpAWmBqlT/Mj2m2ZuecmY0FWZpGRG23+isaYQUDH61U3u+a6moc2ox
p1ly9wwONXQKnTDXCbtgvN513jMAjiUKY+cdQ04nZFuyBq8XXSO9wW2P09Hj
hYgCGYDPSQbfltsJWm9ZNH9tNQt3hqdIfivftf2zYSV+B/BNdwClMS9yPuVQ
XmqlaNEsW6v3rjSDlYkQ41GyWYzYUNiIGNjXl4Cy1yGy090OMZ4UD63AhPbq
ym70f7klgFD+1LrdyvMqiYyylIW135iZ6clS1QrLtv0/AZfzkwSITWYg2vj9
/Mz7dfdlYQrbPNqxQ+b/lSL1otJTETjkZcnBOFUypcZHan6xZU4X1hEyH+bv
hclOZ9JQ6P5xpCxh8oKKba2HuCgw9kEVMDlUai6Xp5U+3rq5tTSV8e+P1906
YtbJ/Vb+Tsu3TX+zsiRIMcjAxtPPaBxaOHGR9VcLPjECgEDBoQBaB/OykC3y
c5BNhquQGGxbEmAId8f4XOg9XppGv3JuTsYsQ5Pi+6pcUmh0JSngCXBgNdIx
eDpSrFifEArcLkrdIu/cL6F3ZBof9+cVEvDMqadqYrjq8z/edBNzVeYAfrk+
HC0RLexXgpW4Co+ImjDCYXAPHgO40bWJAXfdbyJK15ReGIC3aUFkuXGaao4E
qvsMTMjjJ+NIMAXYnEG9wZDXSZnIE1dLqBnOGbJKuIzdrP/PG9kgYDzL8+e6
M6tGhrBzdOr8M/F5D85KUzj1oxQZcQkoEWqAuZt/2/57yVF/syJC3HKve7Al
Xsbz/hC2m7aUAvd75cW+dM4qgRQ1l7fpe3tCm+/0u7wEtSxkmmk/FkCrgfz/
7g4PXv5QRvckFEDQZYqWgiWGH23Z7/anW9knK7jSK1+5uvVPi+5v3RvtFrTl
oa5dQ20konr0UZ5TN+F1RMQgHp+aCn/PJb15wDELPc0RUtQEG9Kt7jrNxMNI
ivrg1MHSMdCXozqaClk5CoWbX+cumhw4Aw4i1p6W+k2gu4ezDRfNUDXrZhX0
cnF8OTHuQGBA1mHxtkeRv2/+WiQ65c1xVXGkq6JAT4NbXl2/KIui1R0Wlshr
i6xUZcqbt13HbRhXreYsLVpCXgkkY9AUfDZCQmIQPHQJGk2CuWh4GJ0uwQgP
N+fEGSb4kyicdPZ0kPGyX0e9BlhMsmGZe4uns0G4MF3YYEw4UEzIguaZCKHK
8I6RyeSrCcnGpmrrG/F/DMWcclAD55BUFrkwqTfJxqWdLOIMgO/gXnFGZeMA
C+0tVCDxawkJjSjw/n8xBGrXFRkhqAqYseYV4JnWzR2PtxSwrJjRZ2AZwCQQ
I0P+Dp7iV50xFrRl2RaDc8OXpB5Oavwyj9joDoY7vduD0SZJl6UPj8lmbOH+
g8a4Ebi2MWST7GlRbcZXNhhLOaF1MyTBoATauO5kDRO/miUkJ74SGVOnjmCo
vZRqiXCeOZrFmMu4TxYh5HeY9sib+V4gMKM4CzyBVAxCC0sNsIYMidcmphsf
ntIPqwSmV5yF1sOT5UOXrjgIgpDuI4M+L7oauB/QquFWAEgaFrMsXNfodF8k
KQC3FkVCGjTSg7c4J9zhB1fpqp4EAMj7bV829rRLGasMrffPt1flVxuJiSPu
bvuup52BMJtr/Iz/NQLtvPCZaT9hWotvXmVixtOdy+x34ZbzHsIei7xDfyJd
u07g/U7eBWgkTnYRprD2Dron+kmskYfwGQulGs2HT4dxzNn79Qdjyo7mNoxZ
Ufm4leHPItaRe6m7cMhjjW9Hl61DsNVZN9i3Jgy6qOGFeB8vLNMEk4MofyDe
oxOGVA5zau5ueVTNVftz+TeJF6qu1vpBL9uUzfnetgxmwwFyUXKVBTMMJvU4
76AiQLO3DxrnsogfouLQ4CSKT+vY4hxSJt4l3D6AZ8c4Hsqhtrd+KgzZoc9b
QnkUvW/4TgwqAZ4J7TQxYB2EAo4GGxrYmMn2gmCAaDjpudzG6mPXDsYx+xDB
kGit8mJovgPhQ2Q7m5xF+on4z+wqYoKWE4pM4rrEfDga9arZ5bcObKJvb8Zh
Vau5XdDk2rT5/cuxVCKs98sfZgCEuJfaEaz69aSEYp5KTtVhLH4+i1xLUb0v
uI9ofSL4mrPDlSQapL4mnhBIyFd01q4Yn2JDkElxl+bm4t+mm9ZxcJ61hhmf
YzcrjigKq2168N6jniOwqSO7MgBqjKGem7hPEwTss2G7lZ3lfu0ztBT+i564
p6y0+oXTkW4y2feN15MpvWOJXL2iEYGtJomwkfumpyGSEOTwuIX6GWyUUoIU
tBmcTK9J9Aafs/2SpvwqLWvRcGF4csPuQ+NOENqXT3a5HVzaWJ/FIS4NAle4
Uycqcv3pSYGu+w4QakO33M8Qgh9fSwp0cy12mtxPtHYYMQxcjN6vFDmcm/t0
QHeEIMDbOqTtLDDl4qkmRvMOGV28vAnGKJfVRPJanUDqJdk50gNXAS6TBNeM
f62AwxTv9dlnQCZkLXfYocgq7X9nt/LbdOHfKhfjpVqFyZMNuPuDo4ropckz
t4hgHApFaYDsHXADq6GRqO0QQ/f6p49kXpmFlknr7MfZoflu7oN17GMaODGa
PSXu93oyzCrb5noGwMDmniUbe7wOR8TRXttD65EYbNvsAsbhq/avqrtH566P
24U3AvpqUDm0449MTQfzx6lNL6ZEsKhZufVq6+lT8M6+xSbeRsD81UJVkAUg
NWNFJeoAQXB1uk3rwUj6VFWpcJPa0w6Zaud+7rNvd73z1L0pKeR2h6ZUgJyZ
lcQprT8ST0JW0B/2UWowhTxdQzyZtaBAgV6APWEkLUKPlcDV5BpuGvJJ24if
lG+KLbq1znbQcdFu/CFihM2fbTatUNdRwhb+nZdJ7C91oyw9z7LnDI7jU7KP
eJyasrj6UBr971tiEIUq1Z3ZgH9VmtwqOzApuc5Y8apirAmQ8Eqv3JNpktnR
GPlzacfHTIFw9/VcAKeOviBXPa0tceJtSmMBr1MOmP68D3pO1x10kEtvh4gF
R9eE15SzIVyXDOjzqluGAkXDLiQVXCiTd/wSprUSDywfH0+aQ3TYdCM+pxwA
Ah1YK7pPY+BUUYEm9nfoJtvM59+CYanpiDm7womiym4AJq36pDgVDCfkHTiV
K/cD7cy/fKRb22YfPxsXR0GKv3KGlxyRSx3EZfE3VL8yW6DTFO1KdEki2jmg
G3P/y0hw9iTypFt7cKOguTAMGJ9KXNNPqOZf1sx7M8parMgU8PBcyE4siGz2
ALzuQ7b+eVQ7vTutUZJdDU/7B5qMihxjY4RYLsvzZTKOxZlG/jFSwAt2hso0
gm/OnyGtFnFlm0nTZSTF6tyEIL9EtIytgQJt2ITD7vA8anN/M0XpWFdgIC+Z
UpAAs5doaKpCcN/G6Dmr6OhqVETfLhBgL12R0qjPqdDSz/U8fCPuM+9IqpOZ
4D4RaciiVx4wKgqGb5mV5NKlvOEoEssZ/tsiQYzF1ZEwYuHu59yUI4MtrjEh
Y3XmC/KtLNBNOP4SIzhgBXVdMPAGOG1QdQfYCSeOUsn+VMFvzXKRC9xGO9nj
N80eUUgUEcvw/nagOL2ScNZeLIKAitf+9pHNsI63rmnB1lerP5hItJ5GAqJM
qutdZssJhPXaT8rnaGrswzIBOL8q5H4T73vJdU+yQepVwJ+xH8hKohzRzlFV
IhevsNweC5JijP8ZniWTlN0bz8UjVR8tMpcj7UnaywuxK3GP+fwhO7MjVnSB
PeNccrVfsEhuD9mQ0TOtT9vlDd7AKzAl6ZIKPxYrGdAvnQFQ+EFiK5g4kuQ5
6MSnts9jOx92aZFJ/oUiyYvqLsGIn6LnPchEMKS7IWmFWLNz9PyMnEwQzTQa
Kwj/POGCzfwBHwRylAJ+e6UvEmJ6/o3RiIfTb8g+o7gdKQs2fMyT6CHOAMPy
sb8YYRp/pGe19fiPcZ7ViYE3B/XKhQGQaDmW5ecQlTkQy1hHKkZhYj5qfHe9
Jh4SJE0SKVHzteq3E/3Kcv0qaz2QfXTyuLlNflxuZCWNA5X8cF3TUGj6yM2L
pQcIJYJJkvlD0rjHE00Z+bMj0ct2VCRERXB0F/wPusAdLlQnrWEMlUp2RGnf
Nxqf5v+AXjPytop/TWVRr0GpWjwDI5kZkquKG3NulkXchebBUgET+IXBcizZ
p3qj4KkFHj7vhOLR5lhiUVdfyR6FaNkP4QC8W0uTTM3IVyIG9zUuKO49IFdo
yj3H6OtadHv+Q0T9+wQU4D6TiuW06bEhdDXrMmOhMXs9+FQhz8JobWpAf0Dd
cn3U40diiZ7K4Bb8IsHNGQfb6iOzGA9oxJDenNBKnrRrWP8Y/spYElAkBXQH
VzJDT/gRxlO6oOrtaThbvUTQK7fELthotpka0cQeeVT+613XIlPW9qswR50N
ZzCxsbPAio/3BwdxiIvjQrT6cNJ9DqzPnHR5P5hd8ZzysGHpBeUAfBy7ESoa
SE4OxsJeFGF2YkBesbLJG9DtoXrIRt8jRUDlsdev7XvhWnlw+Mqpw1D1OL6f
BD4grc4DUzp56YOF+fFNiCUOCXAVugE53oRwpQuAhyB1RRbXNIZEbr3T3beN
k0PANDsz3gIF82HW2JAk19dhy1plU5rqZrWzDlD5VKAJogmvcysjfPqLGRYX
VG74FvhFPGr1DqM8s7i5zJCSbGLtMnknx0QkwRQbXTRjM0nKWZI6s1gNst/I
73XVXmIJot2QpeKOB+5UDY9X/mKF+yN/kt3eZd4IdAUqO8OG/UL/EVnmKhcA
m/N6B5PmsV7rRyH7x2rhTuVz2fgBxZFBPnXgwA5zA1n4oK3V4TgPBaXHvgGv
cKwoJpXDmjcALdX7al78XX6Ewq8c81PQwngIXBP2H49W4o2b6gBnSspPhs1c
E91mJVWtdP37b8xcQWbyUvAEKBC9oPxsfnMCLdJ7zvs+dgVt7qMgC/Zzoloe
MNwyLLt36vRH6vx2trhDA2xtEtK9wpBqAfWGoT8heMuhIh5i0S8YX/xKXkLf
xfIzWIGCcM+L/eaYqNTj5/7N8TQJo7pwl6VvrazNedaGIZxIr9Jh2lbKmP2S
iNVywYpfHsUIqJBXLNhWQVkprLa4q2dXiqKN/Vp2oG3JHGK414JJWA1Vb2WB
N52oMx8Fv6EqSRQPsa624rCM03o2rRk8cvGyW7fv8CZv+HU/Zr2R7OpQuWzv
graVyUmotaLtfFfIQYo8LhydWQ5lhokTkEm5AwbsdHr9Aew/ty06R/p+cGPf
Ho2GM/e1ySGtVuPYvgCPkdYdOiZHKBWBdIc1bys5lNcKei98E+MxZvJ5YvDS
/HXJPp8yBCC3UGnku21RCGYquUl4W1RbS/Ex9wBPkEfcvdOYYE5Z+AwqtkSd
0WMbTKd2aDh9idfw0CjRj4t9OHaGaQXu4WJg+FHw0uBxBcKZfFytRynaQZBj
NvE/rhB1LcaG/CBhNPzB0M9bD2lKTesFDUojh0OtIjpWU6XKnSnfQ6ipO8tT
TOsdqMEAMSW0BqvzBEBPqcBj2nt53lcc7VNxXgLSLA6bJm0NkmyW2pRlw3lY
gKdxZdxk/iMKKKe7QSI2E6wiHdbOsPzeAPJMcFZk4eA3BDCqb8kSvBvve29z
+v+2oCUj2ig+6KxgrqZBSoWxZvXCKBrSsdrv80vncVF+ss7mK9C+rs0+ocAD
Gj3UfL2P3BmELL8r+634P6EodYEUq6+qD5iqqtk//+98vmiQXCBfOp/1uO6P
Gke9qAR1mfzrbDuIy2A/vJ8YO2LZ78Qr6yFdaAvudI533xl1lpqJOv6vUBqF
ic5ppOxnNV7T8515/fUfvm4r7KBljvb75sMbqzHMGfX2g1e3qJTT1VmGzpQt
PYcxd8trBQr+QmQCu1Sctz3KOuhXPx+O7E+2RHttb71Uhqw3YgnmMh/DABfn
f09rYpCXiDlv/dv9QUYncnFbSiflfnNhYtrp7o/JlD1MR6Oi6ozs0pzAkEXk
sTXy3NnO9DdDlIAdHSIp8tLAGrRNChOoI23E7bEH3OwNCWx0+WIs1TrBXDEZ
gE2r6DcTykQVq5LWIo9E0BTpLQfwBSgee4RaGrEmbknpDl6uuiCxj5P0U86o
dmNZsd9Ro7UEHchkBTfLLgFq5unbLOTIasufTLhid7QVAbijNYDqd+lYMcfJ
xzUvGrr8evkMqERT/H8VX6EB8Wzd5Xo9nCU7ngmSrm8ehhoENydFFHiG4tqV
/ZG2llT25fsOr65GFtSDfax1HekNY1xKEFzLarV42hP0qSHxdShMzFBWsJP0
mmzzduqnlV1q1Z2tK3l4gDpTHlwwI1rYD8zezrenzp1xNGn7qWMvZFt2HIfb
NqZT9HG1JUTi6Kl5x1r8r22CGEgfTvoqQiwhTB6tj8chGtf/jAnmtYr8X7S8
uontc6S/iH/G7atK9gQD2ZWbNVqCHO6u/dI2n7VlJcEKf3K2hG/QzHF/1b0v
XFEkSyYK4+n8Tmzq5OLrKyq50Em7H8mOgFmZyZDp4Xxqzl3tKNOusDihRAiV
vl9hpp9WxVGlCNNy57EpEwOT6KpiPfHD/yVzhRoIIM8GSnezuRU5eU4Cd+El
Itt0IAa5j7CozYCRDstzPQqrcK/DlaVDd9yk8/u8I/5DrBHSbAoVPiEvklDZ
BAE7PGKTFnmSjbkf0TH/utiBPR+/j4JBo20z1OKfySBUMqi2sGYurEJCnvhg
5rL55dhT0IDTMqh9+jvqB7iDdQLOl0DhBGDBZgTX7kuGbUY/mUSFkrYf9I6S
I+a6yM4bj4aLa2slla7+5vSzbUTr68OgH+liQO+zqX4etZ8bF1XdQ+RbR+yw
TZ6DJYUVOA877LODiwazSs4F+dtpVx3vMp57otaLk3WTNq/4DlSfKq8gq8H2
6UiIce/1iBzlhW9oYyAC6GUFnM6/zeWBr0Io8p7fbsDDgSFvujwVSF5Wz8lj
0+4h8juhDrWpZPL+2i59XlPdiIfJ0TLWwudqDTu1a0tt0URJrgbIMevllAiq
NK9TfwQruL77Cj92ndZPMis0JudM8jtA/hNurOSAa52W6K2jcPrvDgkN2OPg
RgtM7jkUqvfDNjvRs1qijDUo7t7SnCwcEaYiOSP/ewNmdlBjfEzoeQXcYOnn
OO7iz+9dBoBIoDMTOTFh+V/emf02mT1fCV5sP/7brOYBXduPI4XLFLzJZ3p2
64yzkyhy29En5gUkR6p370YBTx/HKTFPPDc3k4AwAPO0Wr+xAlXPjZ6Ypv9j
K7WKpzQ3DjuVVfkzJYm+MRX1MouN8nvDENf4sigTT/pk2MbZ4VE1mEsJoIxz
CwGPLnzeYfKRJgrdpcUUz/qUu+L6yfD7587Gb4nekomCGQXX3kIZYcx1HPg4
g1/aRqy6bgsU7zbkD91EbByhKtQuZz+aJijhHOmmSQL+KveAsW0TfMuzCVak
k8W6NkCQrwanfDLpUHymqttMgKB3m9xTd8fLgu0yV08HQlNSKSqIsz4nYhNB
RGShu2VLPWV3sQy+4ayR7x6IG9TgeQ1mrqwAVqMBsqdQmW+TvB/FV1RidhbB
Q6LhjzLSWi2XxI5o35lSnkoMorxqbD6NZrY+09rjJnkf0+xZ3dKeAGDOSOJb
x3zb84Leg0mf+xn0JUsXET3ztTf8Vy33hKFtsAD+rC91gwmSCa+b5CxO1te2
VxA8uD6/tJR42SB88aTfSkIG5ZZR8ofz7G6h+WjH7ryQjtSkxudx8UNCU+lj
cfB2AEWxESiTToLS+ehhbJ+tKmTey2Q6pkHXj6mO2L+EOhIHztfjSggQf99I
A9lRuH7EHgsh6QGGZKGOU3ImNRaeUDmUsdaoQHyjP6HxrMkHTzSooKDrPwmR
/rBXWP7hdUyJzB422nof+Bk5h/FJrx4RSwJmqEUoAlWBsVx7nQyS3BuuUkZ4
T7H6mVUUT87AErUwiiW7wMIbSdDGmj8kZyikUgTbpdRc4XH5RFXHvQCDjM7i
4AW9Y6jbAXsXtr7zUHW/kdZELy/LZYDHyPealBW7GAaMGkTAn7lJH9IWWJ/+
zV0/46gy90nZ8JOjym4SZgEf8xHkBLpVZWxyxW7RvnQ7YAbBtqmMhO1AuYyL
yQ8NMi7Occ7FSyOnfeCFMrzdRSXqitGqabqmhilgKEEJgO8OvgbJ5gYD9rxR
1HdnJymwurXJeTsvZyYBotINEbkzS2cL/iNjyOJKIvY2Ii6OV5m1ccr1mIIF
sC6Nlfih1wlQLjCn4hMkJzlesizI4Zbl20ABN7VDJWU8vNuuawPu0oxO0x3+
1IwCodPiE55SQkg/FNHNtTf4M4tpZ/Xz16T1MDUiA5c0P08oplYP6w8VpCAg
0ZsWRB7ScImejFM0FAsOHf6MhQo9umxWKWUVU92zel1Csh9wzMzLd2v9ZZ9m
o/OqlAYsMuguDRRE5gtychByAcqZmb6pUGkjNLM85Xfgtb5e5SuOYaZ8wnqr
cEjf5YVKboW+e3hnZoIQrnX3ikot91p5Fp+bNVz1MU8cP3ZVRlKb4MlzdhTu
cQNjJKvMHSlymKCm949CAXJqY2S/w3L+rsx4eHzPoSymXMp2sRnwzYzh/Gfq
Dsf52sV01++pJXYw7xtswTpyDZrYFwY/tJWfHenJ2cNmsMT9Fede9Yj6CTGS
XrQt6SZXDwotxSGTMPc5CHmhW7AcYrkxIEr6qxUzC6f7UvPO9msdXFgK2KhO
ud/Qa1UcDTgdS5jkyGmNk9pFBtEFd9T2dKAIcNKXnWfDBc2UZ50Nz99epcMY
uAiDZE9ja8w+WlMd2TetUb0AQNJpTalc7bBEnsI8hyzEDpSTBEW19TljF5Hf
p+kUzchuVWI8tUuMzkPj14CcXp/QJz3UmBgP8TKKIJ6m7pKnokMsW/JzoZLN
f7vV/4mToL9Z3i2k2hz4Kx9bmmYWtIgB9/gYAJ6PmEDokQcrcnjnGxyQUZFH
IaJW0kCP1cgntn29MIcTR40guusHmITOTOKcNMqv/gbq5/fRvNwIT+qR5JSn
12feBMdARDKXr70v29N+bOFpfoQF7LreosjPA6eNArqXqHfbTm/DmOejLudF
KlGi9G9g0Xbj2hGSYgQjT65J8zOwwC9tZrpYQdVdBa5kUFLQXbxv1PeQoWa7
HQMpMfRsVZ+hJky6fiU6HCVd17HmmwCcnnrOHpwEPhRclpSxsuTBtfOfc1TE
jMT24Jcnd9G8oSOKBR4iMYznuyGqV5ktj3nZql2yRXvKXugcRXlZAEzG47Ud
h0ju3CQzojfxY1NgeYdCVxxLRbVugIyvuR3VTIiiqQAJEEKm8z3vuWJ6L8Oc
K5nCRjL0RI+HJkFbbkT7qetlcDYvkph2wydon6z5O+fnW5ZEBFdZQT0jRwCD
F5KJuPkE2QGxEcoE8JVxQ+4yPeNbQCWGzP/Vg28sWwQje+95HSsB5Duuw3vp
6Au0OAI8fl1DmFUC8mRLn1ptUYGChm651yd+hFhw9uS/4reXSsu9GMwzzv/P
r4HtJn8lGjENJTbLswpkM3DsfxTGcVq1O0kHZGqrYh3ZrJilP/mmPgyLNo9P
mVlMyfQ7yRQCm91JiIDghf+xrfm03y1Dwdk6nuy6+4W12ey+naL2KW2PNMpY
oVF4lGJVsDvYUc6+H0ZIw5G0jacHDyIUwyM/xQ5KuX5EGZnAeVFwRF4+qz4A
uXoJarS9Gk9ies2mG7fUGGGDQlr1jCyov77jYOvdrY833jTZ1p4zYvZ8MlZm
IG/8D3JKtiOrQiKk4/pN98GZo3xhh20aMN44RKdp+6uwWU+YfeImvDorYSTr
Nz6V6rxlMtIIQ985FsusVpZS2CgAF6dW2AYevLnydQO3lzy4aJjlKONDosOW
UnnDvEQS1XtrgLv/b9dm4NziNioHjT2+r0VGGavBkD7fIRLSRc67UImi0zaT
4Xac6AHZi2vHxC3DuqFXUrekwYYNI8IEQ4p7NbnRJBqNcARdw+UDfu0eo6CN
VLBrn8PSyvRUFKZp0Fc2ValgT47jZv+ZNm1fmh3c9iBQTyPDSODJ4Iv5qQHh
9XFDqprejX1e7Ru72snoSYr/+27IiJ0X72UDzXiBpAznskdqZ7xvsNOuEZ49
dfuksLbMwDGjI/EQ6ewNncG5CYVviGPXklLDb9tsG8fg1MqVWQyLtR6GslT+
GtxgcaYM/5/7Sixfpkw7Itk6MtpGNsCqkWvB8psH1ulOytxy/ocjtTQNQmBn
nt+cRi4uVXtJEn+/xhI7oORPLf2ctkECsFvH9KIOGLudpkrp4ETcRXQp9U7a
Ll/QaIctgTkSZ20Dx7ItvIoaTsAlpDB1vAs6NT9b+wtbBQA/VwLaRqYf5ndA
sD54eRlzxP0DbbDktPCwn/9gu/7ZKLL2iqIfc9b4R0Ii40sDTbqUSDIu5mAk
cSVeA6imBVMJnUI0B/MICWtQUyHrFQS0qH8oaiwydbyp4RMJ0W1UDtiK57iD
jb76jI7dKDSS9eOQRDgJi6QkQfy4kbh2fPGGUNw8xu5ZWA4OHwgiTKeHglOR
fkgvtIZUXFNnEVAj39P8UWi3DuvL1dk3w/IbQeY1BEfLYwbfsrnymUevA9kw
GRtylZx+jhcNWkUZxc8lA2yMFlxU/AGxdAyUiIr/R2Y5S7Ar+iCYKC4fJx09
PCc1CXRPszRw5w3olMwO+22ve1u8sUikPQFvOwa7UU1o/8kaLSGssD335fbU
m3K2bNxm0XvoShimswqByWLvUgBsGeAEZBBb3dL2ryIY17EIYAJI0oAsjUQn
AtaLh3h1tKPCtNBRBYmuCs2hhiNUiqvIcxN2nHWrDZCq4cktCheBt3VZ3N0C
DR5fCrofO14Xm8UCSjEoZvlbJzdqDM9QDAKvzPNroj4rJN7MqVYUpHYy8jS8
0BjE9ogR4KE4qM1MxweY7tmAOMP5qUK+WavIvkxEfKq6VtxfTC/U20xcqxdD
lN0bf8HsfcOoPvWP4Pb8ESktD3FAJ0oB2If/2l0vONhVN3BxPgJym4k7HjYL
P57DPx3cQ770OsCjZJYQ/AJGAlOehwx5mbYkYoF3N0QCr3jPKwa5ae87bQJ8
bp0pcIZyxBG7cVZHdXQ4p1CoiAJ1OlDwZgYvM+HEZ/wv/Oh6fY6uBQZV1ICs
2ZfC1vOheObniph5vng5d0Kjqbwtti9Hz0M8f0Gyusci13YZ0Qr8hB/hGox8
+jogCFajYEgxEQ7HWJdfDFcJ0l2+yM+Em9PYCvZvIwdy36+PPiM7wGlFVdBM
/kb4dDxf+6uoXPWqABvGZVeFLTY379bMc9+YZ/32rhZtJKx1SWGfK9G4FyV3
h3HcYN3ALJZqcQoT/nUKpTHKpioYHfq+Vl0QN1uxpjP69tOqBlcb6nJqoVa5
YsqF+QgZDsfsMui4VUuHRWpgtIVMfZr7dIFZoTLr83l3M6VAQnawXhb+c9gP
c39Xl+FElCJyhTytORs4rhe4YJ+WkJ9OObnJn0vQYAYZhf4ptregWvqfswvr
syHaf+nk07HPbugLI+275ToupXQfwXNfahUZYE75d62xQiiqwmGr+MuSRML0
T4wpuEjDz5WIOoQvbHxL+5qIs8PG2Ebze68wSsOODcNn5DAFVanaVxEzWN/9
hGoAlmon6Ii8Mkw39ajZYJOYw7xEynBE5cNiCjww7Z3thyr4xfwX6RsJm95p
e4Z8N83Q9U1FCnXde87hWVHaqw/V5zZq+XM4VzG+u0SHqrvIs+L5AmNN48eB
xRJOkhSqP3rf4mn01/0PChtbLf6Dp5gdMyoJyIUdyPrJGActgFKZxzGU3eiz
h5u7WK5+NJM3PwbIyPrsaSpzvrlL8ap8NyjXpGtc6erbfJ6rdvcEz/e/eJJd
eRquuLhGfCQgF9nb5I+HSaf4ey+6bYt4pAUQ+bOzYzPGtbwKzE2NP0sNzR9u
aPG7JFa8ohMGyQP90/4mgCJk/E3ewQBoe7UurJoFg2Mc9Wdk5KaKocqk+8dz
wrQrx6Mq6jJRRD4EnbdLdzjsBYx++DTZpW4Y77CVVYF/w5fZfwzN1TJHzpgC
xBFRgISn0KwpvJjzxpM+hxW9fOwUcUAEdaMLkvhuVKhlBzwDpfyC6eogL908
9dWXPy+5HLVb5jr8mbVxsODFTf60fQSyvBIVJ5rTJDvkUAdwwT6VKP86BeFi
EsAGM0miXiDlwJc2EFBtQ3yrS2y1ohmleMCUGC36+5Vk+cM7De0Kfzui6iMl
mHRuUEu9D/xGpZ3f4YmYxbbWq4Gc8pn1iH0iTgjiPaWoZ5B7eqhr21T0CFgR
RDdl2H2FB9fpBoy0WmSb0eaJbmxVFHfgQXcdLboPwW1mNhXAQIhG7I4SPvXv
j2BByFyaLkOxrEPtqEIvqDaLFFpb69HtXVsWpJg/TWti+uOfSR/9TSgOIKTy
pSxnx+S2B4x6lMf6fag9g4NKtfoo5m94mC0Fh7ZA+zJyez+Yv91jcljGUTMQ
6gZGzkuAgElQKFzhlTAq3LXkd69RHKuJ4hCWs5HcsCRkVFD3MQHnqdL8Yzw/
aXdF3Zii9sUQYnUL4rHKnV44DGHMwXl3kUeXcX/pqsVIH61IHfmFtEYoV8ti
Mw6GmTBlvcNHNuUWwj5djJVRYmiusOHvAL5Ad3/ylPaft1S/klXKtZVU5btT
l1G43xlMJuFjSLi73uDEwWjYqst5GK4yoJ2rwNUMoKykTS2q/dzvOuAn9Mg6
iKVu4sEsL2wQ1jhIkil31uqXQ7/NcJnfm6PAdyKWwS5PIH3wC1YHc8jopuFf
hcxHgnYykvVdPo+3IDJos0vZRoEpC/AwnzWiw7cJ1jB2YuFDexTbqB8GRqdT
9sDmanAKNOgaSGaDOyMSE2ZrtCcR67XT6RPpkFYytiSC1T4CipbybmJRbKWT
7W1d6iQlO8JD6VlKeq6tkmxhyVH8uqBint6LXrhxVPMI/IucnzyKPCexikov
XXmvDjSU3FAjBVOa2lumg7+52q2nY9OM0FoSL6y/mYkX3D7JKOsJ3q+Oamao
pcpLamrxYo2tBcxNsll411J/HIidM+Pj7L/2IwiVg3LoxTPejvx8Q6C09sBQ
Edv+hq0KTnvttbQrNhqJO7+mRq8q974m06hIj4bQ7+NyGZc4t3nWBiBWTKVB
8Rd5RiZIYXwHc+TP+lvIlpU8Z7fW0nDdVEyTSkRXHdYMtQpw5Go1Hs8mtjPp
wXsu0MdCQHqEROhv7q8KWsf4JeWiWe82TIdQZ3s+DyfgH3yUuSTTEBoOcJSN
eJl89feMa6VtOMEjHttEARvrIXtkk49zCcZTgzNJSSdrAJLw01XOe4qu/7UK
8oXGH9jt//UdbD4hZMTTKC8aFcCn7FV8GlbIHY7TFhRd+mc/ghqTQQqGUAoJ
0Sh/c/SWAVuY2JZPEq0DxxX0RvgSIORAD8n9UcQRCwYJbQL/zX8mpmNyl8+Z
VWBy4GaQbavsH9qrVUVr16wmSCs1W2dyFwlQVTDQzJ53F3n9I9fvlJ78sNvE
rN5a6M9+q+R4VkXK7TWeRpXifCI3Hdb7kYCAfOL7SWLAYO5co8y1vKxmgOks
MV/vKmMjIOJklPQ7z7Ev7cRxoU5Jzn0NcChJbFQsKa8FwIiyVku5gxP4FFla
QbinKy3S7wWn1wBnQJO1ky4WIQVczPGfQA0HSSdwLblTS0evBA4hUa9Z+PJ/
rASXJnxEK/FfOkyqu5xWqZgImSesTx9okhBY2XlabRolrG8bXckZxhMEt3se
OUd/R1HDe++DOtRrWDFc/tZHMMRhUAyAMqAiNsyM907W76Tmq7Cc2JsXqLcR
0rYiIlaC1i9STeFYULErs8B50IsrWE6CQTa5AA/KAbpr54je8LBAs4xoHrfp
2C0GjNhGmiRq9sxy7nCtS1KSLJvebC2/qwWN1bkegE4cWOsp0u9GusxxIIy4
SP9MeJQRmjBidC3Recy66MsWW5NyyKEmwStfhcUGQxkgmH/mVI0/rOSqoz8x
LtdagvanCQ8HyKyIyvskXo8aDCwa40eSZY7lg4kVJj9OQyacUCD4Znl8L7+s
PZaV3yIkg+9WWBfnuK4qflEmu9Wbc7kamFS9II4gw0BOuHSxVkw1dQjd5AII
Pc9aiZBPtXFKj2GBLayN5DSn/gZkEHroKSd80h4fBOGxamTHztC8pCjtwwca
CLcfPDnIhu1LxV9eNj8EsKYL9pTznj7BVkqva+2S59jzYxjIoXcf2iS/jD/o
uUgA3KgUFyPqIMsw1W41soaI7VvEDFojdMgQ2KmLOp28NKAETwxub3d/JFtT
xoQrRzEvHdR+falzHwYNasONSwGVOz0+L0Ra/zXm9boVkoMVUM4/9Sq2Mslz
U/1//O0trfm0KJTlKHJnHv0zIvRnxjWXVww+/bzyAGbIh6YZYjiRXKqvwJcj
3zcT18/tePbxIU9kX4lX5B7r82HINIjYvojQEXtMo43fMm9AvuQR3A0c4+KI
LBiU9Wx5mNMnMlgQ4YuZcSYNG3Hy5Oke7lqckTHFh543yOSwrjtVm4xgm9UO
/pnrRaT5z+tCQWTNW3nQFH5gYA5UOf+dfTBBkeaPyDieVURoLQilD+09loHQ
XsfHEkAgolKdtF/LtaxQOUTiYq9Caicbv3nKDQCKwCAH3A4aXkn/w0hXq3eD
kDEibcnLZvYz1KLBi2JbBW92tPz6XJS5BZDW7T5D5kRXR3AECrGBKvitCJaC
Ngqbfw/G3TuLd5lUdSpmQfz8Wvu7lbb9O7zzRnlp2gnZSIsYKzUx40TJs2+2
yI+QE4435HaKrVUcT+vL/d1B/9UHa6PSCOK1quHRD7krGKmVYEgCXERHrMFn
K6dK5TFGjtBCAPjXMrB4rrHweJYG3wsDtQxAFYD2ak5sniTFHWRcP2yjLp3P
pI3+DyiR3j0Gm17TxgNa9vnEDl5eRUyANF8vAkM7KDYV4Iz8A+qqQr5b2SU3
QLI7ms176v6g+pifrc0fZ0mXDeDns5d2CEi/VFoRQ/hTLYbXI4U+NPuO1+Uk
A8l7tGfCoTutn4+nAKN9AwMlqPbgp/h6D59QZ1bXAwJuBHeVd3t9QYZ9Yr4e
O9dAjEBaIcuWbamjuUD7+9yqXga0NjW4P3YGvbBt4JYQraKQG/NAzyd1rCXK
5VtQlslDtek+9W/0M4N3KEJqwlWSjkopk5C8ZeZ/7VfPI9m2VeWIfcyYoBwU
8+2Gn2m/PYZg/RnPvpH3qdZcYF+mQYZ+3NN6jkB86yCNVt4e9e/IMQKYlvVN
lPouhVcCHbSfu9w06jiaR1c9zwltmASgkVv3ryeIcOB6f45CCT4IIXSwkC14
ja2Y2hgyaUVbpxYpuBqRbgvleOeDfySZFUSoedQBg6PKtqnpOZ/GNHQS4w99
kDZH0FxfkRM+DBtd38i6MdOvLCoQIY2/kDsR+tx1lykKBvRfQjK/4wG8Y4TW
ppuOItO5cYKzKp1ZVeKncbtgbtAsxZrcetVTn4AydNKYcCHMzF6d541xCBfi
/YUk3HCG83otDO61PAtYmf0U7Xs7k5YY2R/ON2/YTX5psGUjlczur1cd/UA0
9Bc35v/aYRDlnbTktxCuQ+cenmUmMErJCNtJLZToWlux2N1GuZKWvCGIil0H
6znPJ3ecFxCXa4rmhPpCpsbAwVKQm38SaXNm/5v5dOCUCiKOB88HHNwq86a3
HTQByLj96jqH45Gf8Wqw7GgO5f2yIAUdNgWFqR0LV0uHTfCydqhXXpLe9+CG
IGtMO9/W/uvixWKIuP9I+tJbf86fyhwRcWRrnZQNEMh2D+vFC4zzIUQeVUMv
Gr9sakcmoTgkz8G6eKnvmIS0lo8NEhPcppQhbS9l2scHdulnFF3pqWaqFaXE
yXDuwUuRFjluuJRX8FTRc27G78m4V+5InM8QysvSiXcqD989jumMqRbIaUeF
F6zGIi8TNzAjZRueABwS1hBUxOO/v8HZBkWky0AHP79j6RaVocq5haTJs2Je
qeouFFZqGYxAtj1kDGK7T7GpW7iVJtNq8OQrzInVy0EA1UnyC/tEDXqQeiKB
g0gPzL4aHNqbH/kTjd9I/p89c+VczKAiCkaZz6kkJaieVn0dGyCJJ86+0JbU
2+BEHEe/ZW5LxkVVvuMzWfdCw2U4VvuYxyqiChlW60pMXCmRB8yqkbmGMBO2
4iwtYPtZ7SrYEJTswE/XD7iivwmK6pXeMz4vGzVhTFBFRmYcuUy2Qv23RNWm
3lugo6TrGHfP2srPvSgpGpfaPWu71W1uqFFLBKdC4HATns1Zs1zjkK5LjbfA
2HF3Zvja5nary/yMqkJwZyDYyLs9IclHX5RjTsb7Du1CAGLX/6IfK3/KqG7V
dJ2K0ZO4Jt3+n6yFUeRC8vC6hxbVunMaIq8RnxlVBbYEIV+nBqWzLfl4tMQG
RRIG6knJiwh+wtk/74P/F/rc8ctJ0CLj/igbIU89IEGfI8kjhhiidP4Kaq/2
xcQoSk7O58DIZnQFEFXyjVowmGZAvtF5gKuvXHr/K3I1i/BDShZU64KcN88b
hZnwY4Pgu3XG+aoIHkV0eg62AA7hbhiuiIE9nkmZNpsoik4oGthGQvDi3FG+
6IQkiCK1kTw1Pcf/745DkUGqnlbH8Ibvuww1dHWyPDYAQ5aUUp6DWl8YrLPG
l+OdOOIU1MjSjZd7ZRB9ug/+Pz+jNXapxvJ7SFdiG6EZ8ZZsiaBxYIwd84XW
qYTSn/+yu8D4+GE5qPIC10ZpAP+a2aGRspGU7M+VbkHdlyZDw7A9bz+e/Lho
BGyYRDTocO4Xhcsp5xZNopToFCLIIvJ/wt0njt8vU0OQ77+tTgO7eHfeigJM
K2l+PCGVuISNR6u9Rb0Hj7BGPZazBV8pCI/7S1RvGxec9QqOoSJSn9QDqM5S
iYXIWfnb4733/iwoZP8pGhEZXmE7+VQLuNCGbq8isHKi8Qpj/pED7loanyDu
VOVfs8ZBH/YjLPophD0fv6DixxpMkO1iB6RsBaczrX/aw8aoBMIlxQKDR2l8
Eg/beuYJ+ImNhLGYafojtgapBI0ZeaRbySLr0kng9gPPyakyJcxF3YBjtT12
NoSvGGxbExQf7i3Ofqp1nNk0WgEit40l5hWzs/sPtNdkeoqWgyL0bfzLvuej
8hEXKJXHXIlOl7M45WKqbb8wadkRCt+hyE35wWDp6BaLuzcrXnxK4NF9wVlv
kNnbdvwxxLkrkZr0wghELuFDraRIEHISAc3/DdujfPUyakCq8XfDhjxHRh/q
LU43nWr2Fd+nyMoqHE2w5XNziew88BIk7jdm1m9OKeILKv5ZZum2tFqVwJ5v
IwBmDDHAnc9bBTe66IyVrJisQWXz0yWcngKr19zfmO6xC3Srf9LXFUlTltYz
Vzy7a6MKfJJ2xoEnEmmsttUa5ZIBh8PY+ZuOSlgAHCz0TA4aGvOYqxt3titL
QzYka7RQ3Lfh14M6VGfpzkyYDx9YJPbIkUpYHkBwmo6T7Pj7qwdAsPA7X0RU
sovDC/AURHpK+HIvRWloqkU9VlG76IHinPh9KAhCBjbY4bRKrTiu0nhIXpur
UAc4ToLZ/HsmOQcYH+u9T95HTMu3W5Zgco821u03/EWgiAg3sdsXM8gUny1y
uywriz4sZ7y4AdozbULvwwatlSjIAiwZuDAROWpFKeoYj2H/7iJGj4ypiBex
V1bZsHkZ/qFm75SqDJGg+Z6Gasv1k2Kp4xDLQju/LFvs58uWZ8DLlawfnb9o
ckkYM8/ZSsdw0XQzvsG0gJ1RBBEVh6Jyg7yUPojDiAkxio82eJqQSBkH4819
kUymUFbiwDX/1IqpB9yE0DsJDTpwcKPZLocCCb9qL5fXDWJjxkUigAu/hc5W
sKOb9QS9xarSJYc9i63ZE7SRl8wFI+S/saqB68oS/xcdAwgSsO3V467tUfhP
15LHo3tNW4OZuuBg5pg6TDZJtWMC+na5RAxc/jmDnFzTTyOfLlZIcGK882w7
mm1wxYQzsQvB73/PJAeJTbUYwm1f2ZgV3HgQ915YG9ZUqU8jP1dCQlP/k/3N
4kx2vO/S2nGfzQWbahK4f6GP4YQR08nxsIYRxiOvHiJ4f2hrvraBkEIY9Bzz
N6iJ4Tn3a1VjvTxmxRRuknZakzOmyiLNAZk7rz5NmtY7tm1BTyefeeKDJs5d
IWGin+kMErQg0Bbh9eZThqrILc1KGZRzjca1rnNx7RTgvapSxd35X5lZvmFM
gtebVpD4fxfnTBW0z9ONiNjxgq+uSZbFpagoPN4fm0R6lKOAhw8kiJ9sirSR
+eeSKYJe/W6VHij2IXgpyDl9Ub+N6KIdrbCP6Vx+eP5fbHpluHJidgIWctYc
vWENDlIriLuHGP7Vx+CtjiH1z0Y7iaV3dCNJjjzBKQbiWSDMLyJ0HLpYMw+2
TfLNQVAB/lxmH2xJ8185qHrKgd1uncXZ+j8UNu593mKoKJibrQW4aCPBnVlt
z/GToV+HDBe+hfOtZBsprCR3CaRFSJtx740zq+OYIwbSyHeqNSZ7S8lW/y/2
HDH3bVjCuVAR8SKmzCjxvSj1Ims7mudJcalB0a0hg37oh1Xnclns0U+AiA8M
ZAmpM1peKL7NlwVF2pWSEDCiUujEM/naJRKL4+GbetZyefxZ5l4jYc5+AEz4
EGs590T//s0IkgllqLuCbsiehyBgok37F+pi93sdqBAPqdsyA8cqvSHJSpzg
Mxv1ogBlYpzlnmooOiNfD6vmIzk4RNgiz/LkGdzhEMkrs/IUBQq3ZH0hfr08
Jyh1HblU7jw01xwr6FE1/MgAEkzMvggbXL/OwoIEe4VaPCfr0jWjW2kw/a7U
ksARWD6Oj3Krvgzkr8bgr4gSgYC87FKBl5Ai5pHIuI7WtOzxtQ9A/A0f4XSa
fow/IXmsrQSTW2825Ht26luO/VPAWGa2oGRWqkMcVSYI9lctLEy2Fy+sT3zR
qy7UGlAxFETeBusEVT7jhrnNdWlf1Y0nlBACwUbln87sM6CW7yBMqMOw1HUn
WdPTil7MLt0bPvHV8g8f18Az/TJDP494ujuVQeGrOtcFcZpGsazgz05ynWOe
6GVM+dnoFpyo6fIyWFfxcOPczHbs+bhYdByR2FlCoKktxshJ2oWpz+Ptw8Pn
VoDF1ajrB+MFUqbYe0v9+eiZXl1gkWc52ORMWNJcnO3KWdwk/TdWAshIOF4B
a/Wb0vk93h1tZHwq7u/VSigj30cu+n6i2tpzsVpb//M9L9BKTfz7ZKAp7hdN
VOkkSFGxdYKGNP6kVGkQM7GMja02jTmQfIVUTnQtI/Dw+bJIjzzomPPwTzhE
Vd2M3U4nWJH72wQs3KRmj9eY2tESWGaLkGu2SJQF1Pp9Wnnceuc0EFVUK7v9
1iGqQ3OwZVay/31PDqNXLdKBubRRe83mGC1x8qXSp75JtOI19fJ9e9bd+id1
RnuBHEtm7Vl3ayGXJoTvQZp/UanHz22xVd+ZsGRYlozAXEUsNwPgYkEQowdp
yZQP1PTkQIS4SBNL8vc3o2wNcgnHooZiuRF85xzXIZGz4+F4L0g3s5ctC1tN
bDaGKTWpX8r/363egEgmxWMsnL7dKUGSvveehYuzRGE6EGMwdesZGEbDLD6T
PH4LD1hSemHewHX0gdqmaiOw1qgFn7Jes7/eKQcE5K3mm3v8S1X4c7mtgeFa
bxnZKiKVnr9WqXbiI6htyJYPrFCtOSTwtUMZWK3clE8fee0sI3bxcBgTtXvW
g7DQqdl1OjolRvBCkj84n7PtUlQvLo+YUFr19G/7GxDYPtb7ANiIByEY2SBp
DnJRTCkMgX9DBtncoKtzmXVyolADenxDd3RmXnGu6dvpg436lXOqqYdGafp3
4smXF4a3iYPllnvPGCt3Nd+wi/3WcV+XmQdqccYfZ93KSCNzJhGw4BWds0Nf
418UVDLUy6V17cbAMwXyvy0Sn22D4WlO1h237ENt/niSAd8o6X6I1xzbmb1N
RD+LMUIETdhZY+2FFKnW+R21U7TGnOh7Ka+3L9Zorw2AzxL3O8LIEkAjUcR8
8REtfny2dY7Qhduw2nZJJ1yMVTsj79ylepF4dseBa0EjEEh4+SPtYX/vnH8K
YZyjRFIg5yr1d1bB+DHFLkiXglyqQuojfnKKW7lSJp2P7dsFb56xP7IBhCt6
Q/Tc7IOi7nx6eHLOhUFxlAg+Ham4GjpGY4QVaiD9wK/hl9hbxA099H+BwxwI
j/dHujSE2zJuPIjWsdKGsJPSndh68pqQtERquwuEX2Lu9B548AVq0OwZaEQj
DcE8KVBnWlbi+an8zybXeUjj2w3EJLjLA/gd67nipUSc8jvQzZfImT5iAIvW
sw3gAcWPLUJc7XChefTckOlVkI4rD+ws9dOZ75JIrx+I+5CMZXLgU40KrwM9
DncQv49P0aZSacLKk9rF5Jo+d6y45lpJyKeQOFFole6LWl0d2GzA/ke/ns/9
BuTqePqU3HlxD7EfJDrHei7ttmui2wQTcqeFInCFdugU0CFGHm9WkenL88+w
qyvFT9yf5auBW/T2Pnu0C6fQy4UIBEh8YFP0SILInGDEDbxTJgiDO/s9pLPv
x8PZ1ykid+y8v8atD9L9KbAhDwBzC/NzL5Xp+GLnxKHsssMzLzkiW7aVPYSu
yUo4uBDPXVrlUYl+K2t6CfCO2F8gD9EYKRojJwIuC0V2WJLV7r+TIzfS6Kpe
NpVTRvrefZfBI5YRiS9IACxE2nvVRDeRDk2UgyKeBYJPzFtL89J7xjrYsQG0
Rj5LbVcgAFDaEopKDU32rsnD1d37E1/p9suZOOGGXOMMwy9wCuWcDVXLaCTA
j1kL+ugO/t3jcxHKt+LDNM8wjdrk2nq5PEgzDCp/WRxTYnnMc9MQ8yzAXRzH
UzDaWjgD1Thj7kN+QQ1ZLrz4e3MJd91Dufy5n94jnOQQpyBnCTIxOwfUQIlT
SKRo7n5kFQZfQfQL60diobPLE4/v3dQ9gR/iMZQVb6XqkRDVDCfqJwOltkIw
lMaQAA6AHIntG/fbN6YNKnZe8PcUaMuEzGTG3mN4Kc2dg5g2EfZPJKJ+ZlPd
4xNabOeEHDnPWVSMk4dNQ6XG1k8XlLn+AM/ghZEWDu1h167TSDbBLXYY2K9H
FjR+FqC9nhkM/Z/bETeOcpOlsqS0o6vV+USewZ2JGlE8QztO8gv6mfFBzEEz
nJQ7ZiOZ1E4ILFS4wAbkwkjc1PhbCmUkU4axmFcDJMrGeKaOXTla3tKy8tF0
d8Jcps9fE+6AmNDytvpPDtMr2trWT5DOrBUr+7o9ujlj/OVDliKmwdJUiZU5
Nkd4LBlDcO/9mqgHAulT2stbsW9I7buPDMzhbRL9NZp1hVY85g0gOJS7hCJx
inMMyjrwr3NkhQUl9+0nj+GpoQWEcPsmTT7owhDtLrNKlKV953HZ/dOkzFZY
NXNT330lIqbB2kcvK8LEK5qELkzd6OPIys/OPl1YqdSPywQt0K9Oa5NMwvJt
8LBPGALpABPz8YfSvizNo1o+ie59BJvGhjfSsyZS9c0vTuTOORX2f9enAmaS
0qy/haEBMn/7LUHO7HadP3siwydWWWVNMijvAfPrhnIobI93t+ChfWgKJVuK
/naX/psebrzhYPQuYO8R5qT3cNEgvUYLMEr38qO+H9cgJBR70zO5BNgH9LJf
YkQmORQzAAN01v2q2TWqaT2erHhu6XZSIAOFnOZkQmMYmrs8FPLxU8meUu+p
3djIx6UjLzd22tIcRFkgBsAsmFOV2Cpxy5erbLtTEGBamp3zo1cUcrDRLlaJ
nWcS2iHI7A2FJmwNj5OA/X7EaPA5aYPw1/VQekuyvNhWIqiKT90l8FKCA//D
6UsRFMYUk1lAxEfmPPApH/ktTG8rCrz3H+GhIUpeleywtnAvCdEJZefZf5Ub
mU3+up9DKiz8dlrozyazt4mOWE5Ufd4O3VIwuYjKGhvrfRSuno5SlEuf0yfL
tsB5EOSF1fjYzIppuhUU1ogPRqC/pxNCr5JWq83e7h2/FlwPg60xZBq0JLcd
Lr4cKMboZOfS/R5M6c9c0VA1hsrKxYyLI/IJDRK9gvJ3YiB4O4tqemyIAj2+
+fCsMj4g8vtERCNOfl7yTbQJF4zOIemZLrbM6Mt3lNzH5m4ADlqtoKPMoy3S
TWWWXZ3p35Is1A+7brsllkI5dq1DRDzx2vnjXt3+ysIuRzW6h69sBrOvgLwq
pIVUih5wKsi1DVICLHgVJrCgCnmN1Y/N8NYRh9jBx6fmCghQE3YUK3N84BGm
ncwFbpiTdgFm/sGYknEBVTDfm41/ZRwmd6lcDD5U9t5RmtC55urli52FJn/I
XjKalyODXubRSx/IYN+HoY8siEjXCqO06+aDJfSRoRJ3WKYXreudoxnZL2tz
swdPWFefPr0/GfEG0KmgZQbxjJ7fXVqc5FGZmmZUUCWTdgJg1e4TA0gXoEzd
rQmg6di83VZg/bn/2RLgP7Z7L04FpToeVL5GR3P+rzjYgHnjD1epyta9GwtG
QUa8m43HWS0dx29U4tBYo4piZDxcGyyfZ7sUZMaSEXCH/QAPxG0qUhTGMtW7
FHL0oEODxMhBjQv6BtcmOwTCl4rhxCKwJuo5t0yx4o/reALASWzxcvFlNfmu
vO1xwfXIn9PbB8Zkub2CHM/ea2DLo3ns/1UqVmpPNSQggXqI4Qa9+nVLxvN8
vy9Qs8WekxR7bP6CR6QZl+A3JraZuFyh+db2Elsf4qIA8lV/38MXDZ8Lactg
dWj+cTwwKL88wbdDxp3gD1sY/Ehi0bBD9oFgXYzEYZf11JVmPLmW6mhajnln
T9o9xS1Jkm5gQ5NlWZ44gZiReWzqyTiv1FvCtEiHjiXhulHE5udUa8/UvvHd
tWybHYvFJ37s4OaPwrTbBqNIptUiIfkBpAAG6/966ShjgvlujzE4ki0bkTnY
afb46Z7wYtnYYhiHek1oMOfNGzs3w47Osk0C05N8R9fpPjrcTnQZkhuHv0eA
in5+gxBawKdqW0nLt5XnCBudn12XqN1L3yzf5QO3PdFlNu79dLobOmMf7001
1cW+uy2V2esKOR/VKppeCBap2WLqacaMdq1ds1fykcNv1/Kpb+qVxNKLOISu
Fl7CXYyD3+4OafgTSgJYvTLV6NWeOq1lyiNKojB2RlMzI+T66FE52An0c70/
A10zGDDb7lhcJLx6rj76SokR3iogY+4MlguCDnOVsaOPW2nuly2WbB11kdtk
2F9yjEliMNpP3PweAvQTAYlopGSJkcvluBCvutbIuS1NBzGA5pXRihvPzWjN
H0/seEAyerXTw5uq2CaMNOlt1u/rfMsrN/IKMCambnel/38kHIp1s7l+NM+u
1QGTalRHIJVduaTkdwrA9RRuaWKcY1YWeX0Kz5C/GsQYSFbQkwDFw9Cz75Mx
ndwyd6B6PXWlktd5L3BN8Y1tluajVdkDSshs0t63I76guNA4xHHuO3Dn9zAI
CHipFqNvotMM6ZRmS3SlzJg37EQdZ4lMxggW+oY1xnR4OZwjPwALY1mpBHxs
H9IkxDmCytUj7ZMlTIylX9bDPJM9coeP37DW02usIf2IVOy01JtZ0CwSg0G9
3JehCu4d1jcPH4xnf/M0vvJlA2sBXlaIkDTP3gP3hZeGmM9PXjPk5yKdp43y
9inH9/vJJsBBJPsUDFQ+XQeJUaiaLBscX8OnD4LxHLyMX6yfiRPGpVE2pfTi
R3occW4DPoBb7FYC0OQGkDWGmhhWhi14bvAaMzThrv7rtzUatpiILwEbQkPd
LOXPOobQ77gjhWPordP1dCgfWM/XHu1KWFK1LCYZ3pR2jOx4XECHonw9nqFK
RprYFOZrGVxIL+O0N4DEEkKO8eD35hu0eUVNlNosMj/Juzgixjfh/64xZlKr
cB6bKWc8gcTMrVHvfFxuTuVMgblbaUyMhKAYQpE1k/FEaccaULZVewUa1ZVl
LC3fVTQ1UIohlKBo6df4K5vlcAgX0rkqeSRHa/Bk/hA/lNSbCflT+Kpl09Pi
e7tzFJXsMzHc/t1C5iNHxf6pzNTt9Uxs9KIYfDLiMQuM+au+aUAaCXB9xqjG
OhS6zhoql+SJxhNHJXoti/jWrN5D1R5ccEiV5qSUTeqgmgK9dz2TGCKgxuqq
MvUnOXV1xNsXk/P9zYmv2KsymwMLKWB4Csq6q7hjgisxYG+oT9e8Zdm5BZ5t
Pmx4GqOy/K+fMkfpcB5rvuJISKLTF6NSY0VENtEnQDc75pQOAq0CuCpHmCzQ
rpE5YdbloorzvPedmcop8qFerymitlBhXUHqzV2NtMa6kNfHy0T1gSWf6m/3
jECbVAKjYLn7/9+f8nqrP5qzRWUskbAJLR1WeelSCS48GFkgKBQxGBOqoh3D
faBIqK8k4aXamJrjF0X+HWVAEtAlU1IlYDs3lUo4MBj0UjiZjI8KBl6qJMWu
sPodsW5zooccH1bodcNCrKW+JKmr82PcmG6kT59iaLDH2+4C1cF9h9GuIFy5
6LOAN6oNaIc0+WeqLPobrBRuBsD/Y9M9LRv5PTanQscSqWG78Wp0Yt47MuJi
L4jPcrur6lIyhLW8k/1fGLmgNRPMkC8oy1ouJPL0h5T9sYlmN1lNIk3vk0g3
1OJlnN69MDwcKaJw7T9osbSh6qgV4kZpbNYDnZTQQwWGyp7AcJe6zvvxqNjS
Wv5eVvsObwj/dDfCX25Qn21J1MUYgjAcqZq6WSEsKd2yUsJiWYcyX8QSe1DF
WspUoMoGRC6s+F7RjQ5Isher77vrKyJN6yISmns4ZzpZ7v21U9b+vKHWAr18
DPXAlTuySxCiGA5LnRuuQYNqpBNLS7s09jB0ke5T7HuKWiXJ3o6QaM0e10GP
vuFBfgHa2arwV/WFAme8i/zdJ+J9oQV52LjSQc2sQkXDL5SDE9n08FxkM6JS
WG2Sx1shyYdx/wO0A/zl5EtZGa8W836LndWlRpEccIMNayslN6g9wXMY60C8
VHHdaFYtOiH2fEc7L7DYTAduf8u0/DsTDuuaGNlieoHXx3FN2SjGDhGH7RSO
ZBDxm9fgf56kB9qkRHbTmW4YdkDnPGE+dyw52kC5G2/OHR4T8PWen+5+FCws
T7Y08g2oqqjJPiTsIX71q7xI1++h0FP/VrcZc7VuZzwBIyGOOlZVHUHTmynP
SZ59pTVb/98TYKQ/2Wqu6/E6VtcEupcR1Q9+jmaPcQK1WroSPGevNXcQMWap
XLiVXqA22QkCkTQGTttn8b3Gb+LZvXZbYDo4tL+iGEQEkLStOvZelFoYtwQM
8bNvDMrnq7Acc1PzzQx0yuVnNAPWX97n+wV5Vd6hRuPkgbQXwf3zYS3B0m95
0xUvHmQEpSS/Ay6Jkh0kePPKgf5sA8PfUCRhtEOj9PQnr/ryP/hdEJ/1I8Sy
PPySM1yrRpWFuOvSlv7mwchrPDXRsnpvzHwY4qsldCUnun/1bwiDjaHoF2aM
KpADqHNX5MQH4ZNRu68TI0DvyJF4UtyamXJ1MWe2eJlGZR2N6QSQlMze7/QE
M3f5GCCAbhqk2Tp6SjsaubSZOB8/7X1yKt1L5O40j3ao/KwxVnZv2deTDSZL
fxSsnxfh8mTHbMygc1At+XPOysoRUMjHNtyE4Zvkl57CWqpwgewaIjhSTzWA
ZmMzo7Fmf5ZB/CpW+fwKIoG176tc+wtw11H87XXCr/6enOA4e9Y3VAISha3U
2bSArItAgpsk6RJOg0U5L3j0fN89NT+YxE1theCj/Fcct8WB1AlMBD1Dpn79
HjptTbfE86ZqmKCThxY/cEBFpGolGzSeFMBW7ln7jrnkIKVdwKxyOAlZeNZ/
F3345VoBTlj+qzkx8h6BJkFj+L6j1tkBxkXEONvo7rY1K5lWaZqh8zoprbR8
GDiI9+OB+1EcDw9eTWPpZ0Itx/E5h97O/1xYimoaqZ0RKYvRi3wrVEKA6ndE
d1agCIby2nQAqkArvzLmSz36yY46ut7YfMwKWrN/XaskSndV9nCnVNFi/nfQ
nzWetiAbh1dv5pfLfRjZaguKW+W2rB/shTx5SgthkwDwV2kJJAifVnXYcdZ4
LivzWij4sodoUkm16a049aqXKBS/2rTRAIQdqNgy4UZCTc80OnHYWa2QOY+d
vcw5MQtyfVJORLkUka9VfMM+A3O/pnfplKQuFvzraTOon8nohc+NMeSkLAir
h7cn63qNpuHDY46gwOrNXEs9+FEAVILKKtkw/8VFoFkYTfpF9T02wy2qcVrg
BzUiuKYm7VGCrQt6fYFUWn2IKn8pWciOLOGJwldnty9BTYyxiCGjcTW2hqhx
i3euGMkOoMTIDqXkUiO0LkyQ4FYcITvSZ89Io+7TBq91JlurbTZDiRAU+r+R
7FFs3Lt+CDpN7Hijq86KHzbNlBm0Kr5v4YK0GGIPdBw9COpwAPSTjWtbLKRA
86+eL0XKqmZBfmLLVnraurkM+F5vJkVOoL1ugD/hWCSeHOeQ5X4tAb1hg9b1
PFXeQgLQPm644HZHjnGzA8+Gn7CvAAAHX60KK9naIDlYZ2ADbGCEsqnKWfYD
zv9JGmXwNh5pZiRRs7TggtoF0+9DJnAQmV96Yz8WIypLEuSm0/R1ginWS7eu
IZBnAM4jR6RwS3q2J6FaROxnruSpUQLpry7NeAp4Ginb5p884ZSfEJnl41nR
DtiRaoP2hXQbNma0mG99thPeGAdqJHd2qfdf/OXlFJnrFoqsLBOhkM8Kh85U
l2IeIXeZwJqW/Ov4MeFjHELUBiz25ImAW/SxziYHXwjhhmhDStQLO8UFNdpD
keon1ai565TRmMu4H1+ZYnPwhtXyPPTFa1QtVzr+5VOlm4J1SvKUpN2+8a21
zNYurQ9kckBm/K9QQ1EdZovdKlcWiCKvDCEv+JCqs8kQIuKHl0/eSZy48jAW
UjbhuuSXXxgL91G43vlcM+5Yg1wK9pTIRoyyRTKqxbEz2TTd2SKoXV1WUk0T
XDwxENTxQyesBgoRCaz0KX15SF8h3241k+UjQmxcp7aHXOFvfgBHaJON+ij5
lmyBziNjs+87e+xnaeabonLe3YJTXtX8gXjk7ZxOUfGMdFFJ6/pd4jfkzJO+
4WMEWFkc/rnX0tWJizUPNkNbU2v3D39DcVZit+a2671RzZBONW27ludAJ8pj
shvcS0jIdNmzIOgT1e+gRc63yyEBTjlciMThihEg3K4xX2ivz3yn2/1OcpFW
frVBroDPtOlLu0kz5upNYKjQ/hoC0RntFLwM8+TBvr6reUbXqQoOadJAXsLs
K0dnw64XalQIlxhzv/vy0iJENOBvso8Z3fCPytCr2pLqzqbKHgYUK0NIu7nr
u0CDp+GzyB5u3HnZn8K0EHFEGSQvF2eBIOdsEHiwkU7LbCifYwJ0TRIfc1YO
Zcw5y910Kvox80IxjFpH1XKb41dfbk+TYL/j0Z1h/QhY6ZH4tcvD/OhbTtsZ
brmNH6Ihy3OXiVr8z3misD9fFl7Fnm7mnVdro5aOYFDJF2crnlfAggv4I4Am
27pgcSCGhhX/LDv9FVQOsUBaDJKukuF6PXyk+c07MuHo4D3rk6XFxYL47rBo
Thv7vZ5noL+3m4Mlc+ePJU7ka9WNVXNEnReba8TXg46gs1RL3/rcAUT/uH78
fw2v7DyXD3xJlK/6yimBLyMqINGJf2uYEulCv0paBSpcmKDBw0YJARKqT+bE
wiP+3eD9y0oS+KvXPiu5qvAshb5xmMcU1mWO2ZDXvEDvYvLWW0DL4xnSXd7w
5to4ReKPqx6Fq0bLaiKOsJ+TxOScz8D/m5AqyGHQtPOOCCaIcA1BOI3YIyYF
OwGRVwm7OecBH0ZHq8047Q4k0Ct/xRs5TQcKR8PIreNh4P1/AhaMo4FXoiV2
8OfugyiDHiTk+j6fp8tJh48Vc7rkyxp5szBBx5D//UNI4nn2VgM8xrS1c2bi
YRRvcr4qS+uNdxbCqPoRR3qhOiNAdKrv6pGV4a4Q2oJsOpR4KtKQXndGEzRg
7i+mPfTP7NITECDspXr48W/YTyHsbbP8IPywZpdo4I/mw5zgwlywVOcDFPcu
M6ADaOG7N3IQRj38Sna/G8FdqEQmvj+zPi7V0phOOfQgbvAWD/0q7Q6mnxXo
Um+JpT2BF/Sk8FhlO/Fba03HLYuu+++YAuotrkVyjadmcnAyRbYeSvpQuIk5
gONaemAcgFEuUtGkajJ++OOhEu9hY4Uo/RjPc9QxE5bPyU7l939CiUrjP0/B
kjY9rwf8gTM0EeVqlmA6UtBQ0leRXMdNddqBlkmFDxAX186UykrUObzrOKe7
2iCavfTvwSkXQFvEmlY8W/yj5Ge9NWwsxwEIoCsJ5ov5YZx+YvtH8VZoLSud
/OnZRd9DJbtIwIiiyMitWqa74zE58e4Bfz4R0z5X9kr4OuVoRGZsEB2EPxT7
enBRnlTvNPS/bWy0aRKKt8uXedqdHuKh16tCaJq8BNCLWJBvGtiEUjOZoK01
7gvBULUu+Ol4Coi3isb/5p71G7+AEECmColOreCAttHwnqddQWnmTpbm4Q9U
Sz83Kk7VJToeteWhXK+2jh5sC+Uh2HYxrCpikv5PonDiJduKLtYCvqI+p6mU
+bMwzMYaYhguyA9Q7iyTg9VCaxIBd6cu3x5r5BrQYL16cnOdWVK/ZTm6dR/8
XG21mCplaeq6LZS2ZLEKRSk8zGtpLWW8b6o4M4RRGAT9o0fr0hDQEH/7eZWd
MlG5vuUw8X+Y1qYJubNcKOudZkResp9fT5ac35099GXAMNAA8G/RcCfuDsF1
J8+IJXk8GBS4FgKTvWET7azQynJNY8EEjP+NSCz8dmfhbLZ86ybAenSv+FIu
eSqv3uX9u4Fro/SG+/q98KQQ40svkFc0AYCmSuRI3kJlqkTicX0ZI/869+t+
8GOqQt9IuV6Jd7FXNCDSNjs7+MbRNFZiF/XBJvYny69EFo+Jy8f+4DJgyNPi
+xcFcg97jVNelV8cA1mTKT/ie4J7zMugziJxBcEglvs68+IaAXJ+gXjVflyU
9FAEUSzk/HOeE/lYv7BgKwKtcR3+8MoicZ4mwPDvq251PVQ8HhN0bYe4X5uZ
2eUiuaz5Zd7WQuafk5J0mPGFiufltSr3qk72WEkxq2LVUDq+GwR5sjsX7u16
6BjQ1LDOpsu/WGl80idbZTN9XEhibhVPJ+88PlzHG+wzaAjNXCTN4EWC4HJW
53jQ40ED5FUgRLSTQMUdsmhT9vv+qBb0xIrIlTw8Hkhj4CDjesIsK0rQa/6e
HItVylL0dYZ33MaDEuYwH0KIUz/PKAHWkfzN8ql9x9xwDjvAPrCGAEXn0DfH
fmD/aKHmbo6KzX+OB+N+siWvo8XDzvFNusJW0MTV0jZPjcGUWhtzMO5D+3a7
ZoDtuucPoaxLHrauTy/nq0lAcWhqCNmBwYD5I5ITl6y1iAULoIWdGJJYhD6p
hnRcTsPB94zNsUzlNz33T/cHXp7d12qOV+io75dUcjeAMzXYR3REmGA9b5oD
Mg4IP97YdHoOdyUJloMkLTpBS+5DKAtnT/SUT9xW8Bu3g/PidfowSRBJmwkG
mHeu7kSnBQhfG91Mpx/E01Y1lUPko1lSmxafhlq/k1LOzaRkEH4mwEUJSLVP
Yv/BCZnRl7I6YYz3EU4diaUuDJuTVOGiyxvrgnFIHcoCISg/0cBLg2xMy2dB
YZ8ZBFtuXBuqOFc/DPDWjqKVCHwo601e9vGiYmkItbZU3erxe4Xq6zyCLLAZ
JbmFTwcEwXt/mmqrbZo2YPD5fLn5OfR1UCHMym4K7uTmXtlVL01b7Nt6U6CZ
6C4hqzqnVYHuWj2NbtdjMXuS+QYUYlc9LHEI/ZIo92YjgrqkGR2b9NNdCWll
Aeagw5VIeWVWsfqIkkf83YFt14yTU5eTPePhsQ+GW4ouJwt497vq3LFTO4I1
JOCkj3CRq+4plJ3n6dJokbyPQ6Jdy71N3USxufcPXjhxSgAbwxOkkGNpXNvw
obNlyTT0cB2Ikeyq7+nIKy8ob8+uYqMCNwNRhl5hrEtY/8cXjVn3FZSpKpGe
a4SeT4u4rMhixeJXBkPTwiHsMMsdMXa5YFjbJFVXzCpvAwTKs9YEr+I4b5zK
8+mc3KDG4YV8opAyjrxaScTc+bGLnS6ELet0a4mM1U4GB8J/Bjp/Z7vtWqKz
5akw5y5yAgl79h4abCl/qqAPIWTGLRXmsLgrqS1Uy2Z+/Imoqf/CO6ME5y36
pOKoTBTG05XQLkVHFMyVyi6AG4zOVFvZGM/cVVd/u0cEbKuGSSPV4YIWIFuK
HA/10ymd11ZQ5vlntTSZInse7yLpYp7mORKb4Le15hkRAU2RgsSZshN1dfV3
OuGsz3COs0pnuh3vKUtWmQVTJn8JAI5dT0OI6hpdYvApjTQxcYHf/2Fqeq8G
tG/oe49H16sZ6qrP1e6RhAzXz/gP1KnWY90RlwIvA7rGSwBvrwQ/0DsF1zz3
T8Osj6TwPzZv+Mfk+N1KwFQmcmqmY8EcYBz8n9zGzzx+CdqknJ6/LntaC0/f
IafSPgpSmlstg7oqsc3mYgiAUroCMfUsylrq9ofvHOxiVR91n/uGKEBXp0tr
4ENTh1CAoSQsCoFkVucKX0cFi2hrwyr3z5eS0yNM+ozS+FXzZU8mR5b+t688
77mjUkUshekqvdQjblhMWFtDPat2M5DrkTMk1RVukuhPPkZThuvHpxy594+x
1Vr/RQ3QGfAo9y/faDKz97Om1WpI5UW03RVjT0QAnpkGgo1YbluIqK+4NnkX
ZSLNr+6jWvwiwzcDfeG3tSf+7kT4RUkqQcwwUVFiO+Bf3AIjMuxGrzvJapHp
ADVh/gYWJjhROsT/OYe+l9NfgV0wJAPR8LCQN+cJWTXuJ9tKCNJb4P7S8+pV
5y6RUt9aJpmitgRUHQZmaC/ERxqdE28oKvbSZb7BQ5nHuErEIRyibbstZsBR
1i7e8HTAti9kcc9FcLX6t0Jo16QaemNIlYS4n/PJgdMmVwoQyWEPWMyersE7
QUCvhy83JKcQlJwZbEOJfw67/Lt09vkJcr8NDrviRBxKjXXt/WAbGMuZvR8j
wXrbnpE5sv/XQRSydlayVLP7OUGXA+pHGVopudC1jdFtf1yUMNBVFxJF9yQ5
5DgKscfKpFk9w7gP2iZ+KR62s4BASjaTBDRZP304WRfYMJMPKRhdwcmUzHGI
b2ViUS18s500Yd9jvvcMdefglLlGxeZmU0bzpc0+r0JxIzTf82RHUftI0jww
pRlDcCCkgTOEV/4NybHsNIpV2rHoWt7ko6DYgWkK4uMRtRehXcbiTzhNK/W4
/rUbSAqRWLL4B4a28vF4a7kzz3/GcL9Jgel7AdQgPpEKxhlZv3UqgFUg+LPO
VWLvKbHJNRfxSZ/mH2mHUeeYxtZdG9LgFnRsVoa9qkVWEx+GO3FkL4fyCsX3
8PKWZwILJaIre99vmaLWPIAnsnTRwqPimuDaOn5UcUkGm7Ov+fYOk4SKZ0GW
M2eTcTc6EFMoaqAcTssiVdLeyS9bcW8Bcow/y3BUjhANq8FGROu8Fix/Drdd
cj5M0zW+sGudmDU7QdzIHPkfYTXCZs7HqA84QFjLR7zp7j8PXWLGGi6MfCSV
I1pXzUAQkQ4GseocjcL6jVb/sJAhh7hfxSm2yYKh/o4gVA1Ix5UJ6MwI6PyV
OMtoFyf5a4BuDeQI9ChWGbHZKqBYqATfhvfCrlC34DW5idwgGhDmew1Il9lw
VDJDGHuQXXtowcHyzub9wp1bE4uIn+Wiyw8Om3vEQhkXkm4vPLlgW7fPDyoy
fQ3z6VLhUbY8G1Yy+m1tLArei60oXL/BDjHTY0tfcsX6ov/T/A70GZwWdA4B
cKms5Rxn8wpJLmkaUj1deP5s57Zcx1qqIvaXIGjGBzfasQOjiRGpiGIKJDlt
6lxtqTRJsAsNzFCWotizaL6nJ4Fq8HbNqXaxHpULlSz49pGJ4RlrNgD5nCMa
FOWh9MW7RhuEYQTrJdGZU3Um8CDurHCuauxfmeMndesJlAEZHhkNvlBvgEBP
WPjse6ydukFVkEy2nFDMrM3arphq1Gq98yahy+yym5o2/rRCUBElrEbQ+A35
EBRDfqZzb8Pn/Cms/Bg7Vf4ji+jyaDQZ0nWvziEgGASpyDfeFgbGXmERwmRE
6tjYVrr9d3YCPS8D7woArB/s+4VPJOynXIn6g3BRnG68Jr8tZ8UAIiw1voSI
zPUUFFpTEw+h43WtYTz9d9wZEr2r3lZA5mwcZD4QcAhs8bECc/G1sD3uPwEt
NmGbN/4RV0Cnfi7gxwUlJDl0vnLs3UMUbxwFou33M2AmdHT6q6GTHvqY0f5Q
5z4+fbsAO+vqtkGe+bglrBP8aAT8uEXIDKX4XzwWY2QyheYCXFwZZXdNIKSG
mBFrmn2kopGDYZgei+9Rvb58VFEZXwJaEhA5A0CCsSIcQYByY2G/q0S0twYi
GVHU3tbTPWySdcf9h5MNAaUnUD9JJJHZxNNt2qng4Ts4SSZs67LCTNhwXhX6
wUvAtuE6pPHEafjWEbjVyFshu8xu1Z8aLLOFBt/aWQqEA6OeXm4TELa52hJx
L+BiJnnc3EUOo+RMQquUW86J4uVn8yBiE6kFJ5J6LGq2k/DF+E8ArXv9476f
ESjo0SIRhjuD4pFtfu++j7FvKPkRK3OHg/8pIDP1OtlXESh3+1Uluyu79g+t
54yKb2grDd8ZP9d0BehxrPBnlBDSshqbBytb6G8fgG3peOkhGbJgJQHuzfSf
TfzhrBlhX7nsurX2HF3XTwWlFuaJynSkNzgSZVwK/Wgd52s3L4lciWF5nPog
z8Y2AAtfdGiIL/rJ+R8bX21Q11uOMpQaz7MN2i7Tc8HvOE/UjPV1gMdy21qS
2JpN7xl/i7b3MS+Iru1QBcPhQilU9Akb6mEtxAgR+oacvLpWgsjQb4BeHAA4
NHGNvgNfJevJ9BoZJdH5bgx1l9F8RMKcDDU4yd7Yuz5cFMaQRh+NW8jE0/pJ
l/WjupHiB/glz+Udu+AB7cnRtxh40wxLHF1gZjJ03qXXc9XaCS9sJCKSvvEy
pV8eWKXqNIWfxZSCGrWxxDr4+eXT6G9rjiRagEoc3tfYZ+rZkTnMUSxDskHt
R7jx6EjNpJvesyZzjeBppozIL6O9FP43BoyCLc+pw41cR2r1pVftGa1d6bLM
Hwxm/j+Xk7QkXF3EXm3D9UwbQJd++tCGx28sb/gXCoSQPfnIe3dIpehpTlep
brQ/ux+JxngwQUZcDYGc8yo6ShdmVGaTCP4UF1IX2Lt+d62oJy/GxJ3EgHOY
F+iiPH1wnv3QLi7h5BYlkgWJShVYO7JPYmqZIYmBWnJ53t/ycxg2a2kDhLkl
Yo+T1gyKhQcZkav5yRLHY95upi3dKVdOM7X7PateJRqILracnCPEi3wXTpdY
79cMWnVxjUW1EMubbpHKWM2bjOPWKme21z0WnUz51g2ruBWrUnwLy5fD9Yfe
VS3k9qAQAqvGLiGgQenxH97nySqTdl98C08Pq1SexgWkTpB1vNtlBNenXgtP
gVmzR8Q71xUBU0G5e1kgrKqoQgVFGzrsNo+BjJ3OpBN26g6VNX1E6Q5FiLdu
qisxnVZu8hcScYjHnW5yVtrVERULC/f+PMJMLVfUuNf8eStj9qn85kychRXv
4SzBIVaQ7qPtQWB9YNgUJ5s6MAUQWznbj/WhNAyB9955WR+Tc3tieTdRV3bN
cFTclnJyiu4RYoH8KD0YKB/Un+EjBWxy9OPCorMBKHwqjpYFAekFNycV3i8f
PfWEvdCiuxaULcvcvRYk6usy1qqCx5ERN7J+W9/WByhKPXqn37oPY9oFo566
CxEeLQhQw6tNO2eZGIUsAdYnsE8Hk5AJGqSWVJpZ51Dbc9NIlb7mM+ahXt84
HP9Q8xMJ4PUf0rtOZu2gRejU2eSvZNPwCEUq1GwGA7q0b+zW/tBpfSPYzrJy
PqddMR9FSw6OC1qm5rgoycplf7jn4yvVTm6UDYfblDf1p/DpISqlF7WBgWzB
8IarwHrRkfIMy0WPAhA9j67DdR5OQkvh9pdM54hZP8Oho4P8PXHFoK8tiBCk
njDzrOXfh+ZWnEEN3SV+Iyj4LSLGUwvQDxMOoIRJWki9iNZ5YbiWg463lFKW
Gqm8MTQOwGebj1PPTp0BJTxisXOVH3wlhT95IdNJuMmiIzr6hOojI3Bwnpiy
VrJWhIBGceyZgOn36SG0cdKMHqTy8en2/zwT/Cu41eOnAADd2x0zE8mNPKMQ
7cmgUCN+PoIoaJOvhY96ot6Exvcnmf8ZleJYRlzq0uGV0XE/xSyroxuOqXqh
xqldqUhkaD555yad0FnnfWWTIbZ4p1jHXOiLjOxrcko+0PtvLr86YmRoGVS8
ADN5T8ERc4Zy5KMTNwYpfB2YdgAK8H9uWUl2GrXwLCQgNdKy6h1hkkHb8neJ
WLYLsx8p2omPdUTX8TF42aVtG+A8HN8N57mpRCi4q2w82sfaB+Y5qfPftGvF
R8MLJ6Kg18FkO68bnoI49oKH2zmt8IDe/XnsOn2VmsIlHgvS1FD+tGPXNAjY
XWsTwXSqV2XGouQloyAhllvpKKhC0e6yB0oUuobUH/rZMgcLxLwX2b3XDrj/
ZljTRisandnubwAqI1W53leoS2UkL6EEgH4ySVQvW4LsgkrwrqT+H8Pd7Opb
iaHEaWa5b7RWB7a/lttgvprxFhqVuUaVWTX+QrSwkx84T2j7zTR1PWMHgQOm
9d4kI0XHTE2/ydfsuDD7gPNPu66sFrxl0wwxaeAHM6sxIRhR5Z0k/JwFJ4Pa
XnPg576K+5zuDzFvy0xbVMoevPE9AQCiMip2dyKONpsK+R/bccu25MCoi7u4
AAaf8HnKW+FDpiuDXFvtj49jkxKmODarx1YpjKLIZ19Ses7aFwhG21jmKLbU
4KiAJwQdCpajOL2VgCR5u781efA6QEdJ5fk/H/ZLW2aUzw2HPbl9ggpDYDEH
k7EP068wQBasget6ZkZDwSYRdxZTFzi4mzY7HnASFgIMRauVUjSCrHu+eA09
bc+SB7S+HT6Qo9eq4AQHWG0zUI7uKOP4wQVaaw6Jy8ePOHe1mHce5v+HKCN5
7OimXQDPX7mpp05na1N+0LHtKtCie2dPaBKU1CgQpE4/AtqwP27eZPtFiHTI
jKgQyEbT66mHdrPYWD2Wg5hEMhcQbrUMGzS2KRFOES71VYBH4gR/eaE+Drp9
u8SjjpoZOcTL41FDaGIbrscL/C3jzYoSFxnCtBwD6NpQmNBuYWWCkQw2smpZ
g7PUf/wVu0a4X0DFw3Lhy6aNWsctyN/hM78N3VFwbB5+OdH1EUePCCW5qW/Q
aNbskWjD2f7F/j19huBz5nNJ3KKWeOh/Q/ddDtdwAxGC5/taVOf5wmFXrA9Y
ec/dbr/1QkmVbG1Y/UpUlzpFINlA4gGScFV6GSpTqSt39RR2qUX4EM78WLoR
I1drEgRGn2tJY9NRjFxCL1+77oAM+6BCDfhrHN7WvS5cu4BkN3hdH9mNAucC
5sV4bobHizFL5BWB4VwXn8Bw6RdBuhKDytmL2Xf4TedUU1ckNi1LBr3w4YgJ
qwA/lBd0glpuHhM1h9P9OdELEPwz/HCIbGb6Ione7ut0p+ZjJmN36MQ9N1zI
ScBS6k12IVnTLGyeAiWj8C81oYxHJAo2cBrTUO6+AX+56plwgzkZ+BTrrYeW
+zCFFVzAR4huiZN7iSaObLJfHcrHP79RcqYStOjbQmgFHdyb4fY7Ch/KTxOr
h6Jl3aWqwmykmBNu9DpVRQlcG60O571fnl9Ikcr6qXb1ITZKYNBPtXJCknsw
GDBJ3LIZnK9UAX0WJMQsn5xccR4PluGboNaBEaJJWqASwNpiF2CnyBl7X7Sy
1V/3RpWpuT0SaeeCw7tiK1hpvXpZoSyfbtk1SyRDxPV7h+lYmFaWhHC1lKF4
60q7z/xmQzf1ot2N03qm8csym/EZ8E3y0NPLzc3zqP3I89KM1wT0i12aBDbE
uL2ma6vqE4Qo1D0k7v9h74Sz2g8v+zoDXsL1DbeH8CxGzZUh9NhTtqQ4mbcQ
z+N3BSSKYYGQExgOv2eNaLirF8Mm7a0kbSjkCg7WCG3eE7sLiTV16rusHrAa
YjEHtpxvgJmgqMw/gbpk31jtoc55OL3eV45D4i0l/2CqUq0Zufgx93JCptLc
h1kANl2ogReEyyWVEPBCG2fDS1egqBE0btPYGbE4yf0rGVrMcO/zMf7YDBEV
CIKr8MsBw7nFx9lZ438Y0UFTR3fgQ4pPa23XjcH85h7yTDSNecGEjkVCsX1G
INHZKCiM/eQXMMgpwRc/L5dMkkvj2ZuCG9pRpsFuS261If060U3ZBrILlTzp
tAcWI3foQkjA92ZvTUyGTUMBZo3mon6NlBDRf4IAZl3/sGpeHiOIZPv4Hwht
diD8Tsp9KYFXGQdAHbqIyah5VbkOwGG84pSwirD6QDlPJGBCAvj5rGGx1C/6
N/57VBySV+rnqDNBB1Zsbg7glaPiOB/TBXutSLa86zDRuhryMJmdXLbWJtim
mkn4oN5oZl7WXhaiGdyGPT/2zjsIBi1IzHCymht2yosqCo88D1rGuKgPjDqN
pTXsjRPzmSxtUKQDrV2hIFCK0t4F3zjXqP0eU3zYZEZdWHMzvlYffAJxfYBe
9+mc+1cGncQC/QwV+aHyjClRT4jOqTrsRG1YJpq2MbbirKcNCRYKxlp82gvC
Wr9GZ0mTkKMHtGldp1Z/Yw23uoTWmxFaSAobLOlZs6HWE2iapPdw+aq2uiny
ESHgJbtHMuRP+kWxm2VYyLLK1JIwcf2s//bU7fg5G70uZ8U2IYP5LQDkZyew
HE/IFMTsG0F+cL6dGhaixVULd+an5zQOVkbawqJLDtVzoP5ZieNz/TA75hDb
TGKA1AfHnVM+rMzGpnD+zosV1a/abmUT94wz+8jIb3x+ZMs/vg5uHyJC/Gzj
BmWvNeDik/cifESKDSHh85fEJI+9yPfgjNed68SXtao50/smQ3knU9Fr1Q3T
jRS3Otn8dE1DdLIuCuAz37RxWsnCNetTKYanalU2+3z43wg1tLfXMGCPKRFu
CuDhi9igSKaoAx/TeVCjMcNTcYilXByFQPva1JaXUg2tmwsCfATE5VwAoUDL
MBo3XGtmSK0bMT3bY9edVRkWk6lIfGe9Qsg9vaG9zSPh5rEcJFV9rGg9nww7
tLyEEunsQjW0w4nsBwlUCqehmy5HM72B15gLcT8eXdNcqcBsfpJBZrgZ6spf
+lJ83su923isoNexKXxnmaTTjMupAdw+a9G0y+WWpw6OTu6X4JO49+wjjsau
Drqr7PJal/vLAWeQgMgers1W55668l1BSqmHOUq1Q41LDj8yAZOF0M7dRDdy
Il0fxLElK75uUN8lLb70Cv+1GjHJieJzPW/u6o/Mpow0gfD1FYgaXrpG06uV
AuwE1s5PG1qTcZUDIC5Sm/7hBIgNE5suTwF5ljb3pyCeQRzN6IHBDwvE4++u
fmTjVSHmg8rNiXj2E93+JrmmCYNG1IHwb1z6aJvzeKbRPS3fIHOcCohI33I6
0X2E+/WM77PKWuWTqtAZH34l2x+kzF+cg7pU/ml6RldIsXlTxDJh1RmczK49
cCGTiu0Kdw0N1ASeL4BYhdGY20Nb+ZiwKA7vn4NkKP0UJ+oVpmzDRfCp7eC4
M41yCTM5TpBiPALWKry16Jh9qzmMUj76N4xUs/0zKzB/n1u6WgHL/UwKRi0e
gbsFMFl9UIbo0MHkQ/XKKZOHoc7cAGyHstkb+mmtmcyuL0hD4JTySp+KWEiQ
0h85dcNtSZ7Aj3+N+b+9WeYdadU5TLrQRIb83ql/MEjn4WxRVYAskPYfhyyn
Iq0azSIdqS9+VcTVKA1iKUKY6cdAWUAf+mJaAl4isR52VWsgO6V1aKB2EbXh
VrQTjTF4ft3Gjbb+juFKzxBihX7zDEQztl2QY4d7IbFAreoXEeDupnK+tyDo
fbtGzXTr5jIpvvhCc+vhmyk24eO2h2EPvjYBk+6ghjNVqGHuRv8Xu2fbOEyA
cl7FKwBuThkRNqooEi8lGBLWHuW7ukPY+e2M31qxE9oUZXwZ8/PwAxZKOb50
5MvZMbWpC24HfK6Ob6hs5hQhYvYwdSLF4aoqpe5OXqjChIgLHEaQ4tQh5XEy
XrUOYX8zpjWDm/z8IsnCOXML/X1AxISnOOosH6wFHIPx/7Lp84H1rvj7veNw
zCxzxLbhGorBqbPVTiITQ2+LaavAQ9gnoLOAiFlEMfYkiokAhkTXYpzTxItP
Vea3GEds6FtA072jTsAKKncA1Jde6NNjKne73oF2WKC7/zLMoTdHHFHGYAw+
3SVWICWIumsQgnqqo8usqZQMTFLr0VRCcKrfnGW/d3Mj97WDjiAGwjzd8303
VngWWiqoogkanndcqgqeeQQnveEwZvCi3y+8T4fL4pt9i6jwpJ51ZHFYYPx1
/ym/jx9WgsdaUGxhpBO5Q/RogWRds7mRTvYJ+ROnhSQW+blb+T92AxP6IDpg
JIoJIfUIQ7KnJVCJ/lEfmypcl4U9q4fAsI0Uz0AqkFq/0IEpv65q3IjQCYcH
u0T4Jjta+bINbwSzPa/leKpPFHwyCH0vUTiR5BjjkCa5xjDDDZ7uPj/1mQu8
pa+5OVA4tOK05sNdNqWvGZE+Werzxm4WUI/Q48q87nBHumEfixjbmDqdrdIs
yqO0ism9ljX69kkEI8c8qL7r7m24taFPjI9NUAL8yrkUO98/EjERcVIitiu7
XwG9hfhk7VN+J3ixoGL3u96OP13qEBTLl04FgFbnolHQkildHDBRR7ixU6YV
2GOSvBaQrJjAt/umuU/eZ3LmNf6edYQUvU3VV6JxLDF0Y88vbKCNuA5r+aMj
8MMKHAOQRmCI+GlxcbN8KCIWKe19UK95l//p8+nIp6ynMC3yvnrcUCtdoJTO
a7t3Mcp2j0dSgfuW7dV/iRsQxSqAX19dcghGqqddo977uzDOgJsIhKR+NV0t
3LxIdmWG4gARFR869zgESDd4VlZW7cF6YM3qLPn84UDmB6VJwTxmOmT1/EIe
XfcNCKx4bi2y5vlg/Twn+u24Ek0PoubJ1nS+PDDkUIk1sf9cq8+kKbTk7l1B
BaUSC8+nkpsCg/Y/CfSQUoDFW8Y0b2YzO7g9TuaKKFgO5pFtgSEJ4qN3oI+V
74dU1Rubk3zmsn+0RlRq6AyXhL+QCTdlr9qoFk+bZ+RdXVcjPkNfLf0xpgqR
IubEfPGv4i/hJXg8U+FDmkwo1WDD5z0aN4mSL4pknyRSZXSaBZ7MrK6xJeZV
GqY1Yro3KZbxkHp0hp6RieZSY56FkobG20UeSNpvXo9sviDL21cV0imobvFI
q1w1JsfQSnHc83ktK0KxkdfNUnUUMuiFb0y+SLYYEDR9Zxnv5fvAeOrpVdS7
1dl1vv6i+D50bfYF5gxgt2kRj/QGnzm3R13cx/oFh6H1nUDzVhxLm4wqop+l
BamNUarUHvaKnJiQZlgCNyZ6mEjxsxeO7DBFliNNR5EF5G4BcwCMu4yHXoDx
OnZ+2qv6/9RynoJj/E6416lGrpjba8r95J5VfbxxKsCz/GmnMKGA4t1wWDue
3xfaWmvQBu+lTW+sgPj0C7yPoh0BHvcGO4nzWS5mWB8MJX38BjmvD/ZzoNV0
m8cukiAGfeT1l24nprzQG4TS1Y3/bhxb4W2T10Hl+MJb5ldOSuW9DzR+5PYB
2gfUqrhXtIBq7e7jKUTEdUcBr+4r4EeFfTSJEpHXCvMsvCsSG1XMM0ISCHWu
GW48MRYNVcrG8o4BMpNRjKGKjUaBodCoYcLnEpYZf5oiQXB1P9nd+/fcOc+i
wibr1bilAp/ECaUDxBPF3dfiGIgLbtRp6o5fk7CV+IDAWMGAyNlqmPLxxtrU
e3+jwcguc/px+znwbxspweIwnfRmVFVSN1ud9bL4ErmXfEF+m5rDjF1A48vZ
mbjKd8FaEfLXxRfnyTzCjDC9Z+ac+JhY73LsO256Pu+Z/ihhAopqFby+m+Gx
NZKPpShIMNcBbDIe3ZGsm+ahUg4z3OoK59ObIk6oYX8NyZzcoyomZWIo5WuA
75JyRp5f0y6FuXkogG56WkWrflPJyrril7iCDRiOUuZtz9J+M4zwhHUZQQLd
LXuYhiTzSFKJNjHiY2cbMeKQFj9vWX8aoqw3rEHPmGEeaF7a8m5H4uh74FZu
U1t2eeargKI19vSbCv4C4mReHwgq0xFwVSn6Hy0eOB+Oqm8Ayzhxj+w8LTWi
mjysMmieYYncP5C7BrMxq67ex33Ixij+eRjSkSXoXGgTvFZvQgJ+M0+gUcZH
FxKMUB9NUKRAJPtoPU2I0VvRI1PzjjbpMnds9oGdwhIiKrsgd0tzS+CtpHDU
lH26hgg8W0n2K5wcBAW+Ai2Y9xGCMN5rgXeR5tiGWx+uEOhZwFgh60O8DwJF
lcQ+EyRGY/TCSpmo7ELZ4lKSscac5F9od/FBkj+mcolthTQpFUD3QOkr4Rj2
ZBlDYW6ELxtc9ZeYtajdDTWwKgHdN5TZO2bbyfFg0bsEYWyq6JvuecYMRVP/
fnAyTJsgoDk7i+JtYpzeJi7wBFLJgIsw3oWNvYswaSsJTQcrQ7of2nRj1Inu
BDhOjbkvkV4GmIwpz4zwlGSttMRF+VMevDGiwD/SkKzp4QkcS8X7wHzZg1yC
0CIjWsFOZUWcuUQ4sVttsQ08gDKAprzOyC0fJZwzOerrrlk2+OjONrRBofs0
7x6lWUiM5buVH385EWT9Q3WTDArFkW1itwbyuKRRPvKQR9yKbG6T/uKnHp6H
h/sKdDu3CwdN6rd9w3sZHM+Y8Qo+c7ztYfSJyLy+6fnPZdC+fOAxcRSMedYi
aJLPrzvmsS+44sCeKX6MckYp+60qtA2IhlcnVcbo9gOGompGN5uSJDzp6V/b
hkuZpjzfbtVN5qo7eENCPApYDIVYcUi3CPGi3C4ZaCyJVV9ipTix3IKeB4cM
H0O533G3palJMxJePpTzpPBM7jJYhrfqhQAa4nPXc2fRXF6N3bBF/bN/ff2w
vqbKi7UtMGvmrr0KpAv9OlLpNW+sCzp33VlBtrqrqw3CGiY4SXS8JtVt6g+3
AECSPVz8epVczRK0SohXeC2gg7izMOaSyG2XwRtOjQ1s2JP0iWgVsDzUsHas
tzon0yHQ0W7g2nY1muwXQYYr3DbYvIjbApyZB1TliQEemxBl6oMJwjR0r/EB
LVf/3N+d/5RCRVkl63sC2ffQuvr1Pm+D8n+CShfdM6jRCzcHgjHXx/kIKlmU
KxPKXVXm3bgnLcUWZH3M7vQ7OjfVNYnTQAKZyK1HZHp+JMQF/Zd61rhy4dhC
2RmQF472OdMRtJHy/8+laF9D1X/iv7Cn6j4Oq9rPIM8EOhdMw5IwSHbkXeJS
DFF0KL6TeQEcV4CUMNjp+nodaxaUaSDh7wi/Xq6xI3+47HCHqMbSwMQfB186
0uEcPPtyIeeNvlQV/K2Fe14eWdlx3PgULoM+ae9JGdo0JelHI1C76djzXRkx
t53T1sswekepcq2MAeTGem6i1P9pKBeaSjEvMDTLhGs8y1afPLj0o4RDy7HU
PofQrIELsgR3JaBU/e1x35C/hdylJh5tPZZMF7Kfi6sxCBMKKfz7eTVSEEqi
UmcFewjJWU45DNgDcQeP3amYjIKgMh1z0fApd7FgFin9wFxRK8e+ynQRiI9t
2Q2LScA/jfOYPjYFL57mFvFNAn95r9xajUSjDFs7wwdoezgB6Vi7GDy7ptGq
YRUqMImw4FTZ2CjjQwP+/kDXrm0bjpRqmn02Nbs8AN8IbMIHiX8fWFwsaCa2
PXxtNw7J3MBT8+RqLoKLyFN5BOvue8dCwStxL2QE+BvdwTPr+FM1LhYMLaW/
w/jeMm347HpEMgdgg4VnlkproxyAIlg/BpeT3HDuRMJMO9z2zF5CLGs8wZFl
DWmsSzdyQCzR7iJyCOYrCxcGVxX382kZ8ZjdJ2ST1Ff+lbzmtORLE4xLIBk7
duY4JAnaG9IVVCx4K7jtmjUJ83DTGQe11uWGDAlw29xsGcTyecGQ7CZVifB2
up2Brp95/zNaJW0ACzD6IcFmvwSe2seUPwBCqcHcnldWu8O+0mHyvIDePKBo
5nMn5THYgLd2L4DayL+3Vl1HnR1AHLAoaxN4gdjmHigRMAwPr19uQIKuN9Wr
lI/J+UTbeCMEFOhLsGVTUecsi8vNBaNh2EPA77tzn8dzuQGLWzUcy00jsiK4
YKp7DnVQqyW33/HXT++d/XHI3de5W0Z18wdD/45Alvt3IxE9ZM1TU/DpVCEo
oCoebt1e6DxPYOKWFG2uDRBfcC06ff0kYkn62GjdO1h0tnosae0Njiwu8ZQr
kSEW+QzxCVX6roVvxxL1cQoISSOZTErmGI2e1d850HeoFpRnU2Xf5vGN1ApD
8OTYY2hK6k5pyI3FXzB/iEXSP0NuWOStBrDt2rdmrfB69cNQIaDdTyl01PmJ
JphwsFzEmOxCIv4/7Usf/7uahjqObt86xPBJQMmY+ASnuz5FLOPfPJ/cu3c9
2lPX8PVRx60GVp4+d2QJq6HYQCVcFRwLhTYhI/+rvd3YNCO+mdFZstMX9CVM
8lGwOrnBwo0AzIkZMpAPIeHIuucTMfTeqTGSPkI7KeW9DjXVZ4X5h3BZk3re
IcfPjcs0BGXVowb7HfYBbUeLcsx1oyc53eGNZ+nXKjaj1nbLSP3WgicB1/zj
7Ev9pv7jxP0v1RJ0o1zAAcenfTkfRJJyGeRSzHjDfnDu8Rrp68yY3t6qGa9/
e0NmNRLp281beQgnTygT0dpN46G6d5Pj+FQSFb4NS7qkc5AvRL6X1e10F3Qb
5hIQBxKth4NK+cBq9+rXowP8+LrzhcVJ2AiYV6wLV2pYkcXbw5kVRfkg0FBl
7gbU+lYXxyyyE9ntA+KDsPXUb4TpS8BPERy2CzhYmSl/RrjekHx4DxPhDCJa
XJa7iAl/bFQtAvc1qWaOcc4t44omsSE5iPRZXIhHKhlKkWXqCwTkqSOQczRg
cOBZGEYFjcNxFFOS82YJKNOr+PftXAo4Evf/tUKuU+Aqabza7upzL4nURCon
MOmXnjw4RkWpNEJ2lWcpUSufnxZD2M6CDbHQEM1KaTH4BlhdkcrHJeKlELEl
MstCKisjx7CGVv/5WO22hTfWu/prWUxA31ewI053YXzDivEl1L+Fdi+yygyj
28VJyF7yZcmjLyItQ1dJmvIZkVdtvFAoA0s/NljpwKS7YwLm5G8GF9+EbtNH
ePlLbGH6vwGatQGtzg0SSRTXncaM/m7fp++iOBaYgzqgvLO4Y12ze0vWbeAx
XkzJyBtPUYPwIJAeiPDONhRiFUZJuSM5Z8PxSDADjuRrWTO4SNiGVSpkV3V/
j8TX9ilXnMOrYVfr+6kWLWdHRppwraz7PWP1MvtRqo9Yz06G9OtQhmnyTFO8
mO/8HID6hxVcrbc0kuKCA00TQnoEz8XaO9lJ1xDEyqiQyOpkYS8U9fxU786D
DbJOMRfdAlXfVhyJXwlx09yhH6Mx1QtXjjCXCwCPEa0utgtW5bhBVATu9FiE
Fwqzwc+mP/7WHvbJNSUJvYXNADRgG4ytnxyiRrcywer/kQ2/0U4Vg/rlUjGe
/672XxlZv+59dZdq8WzXCs3BY5M1rOZ7hWsDQHxXR9THEfh05Q7U789J9AdP
15dbewmecXq/RDd0z0nE1NjKttIKz5pX+CH1BOf0jrI7LTheG0ThyyOv5/5g
nEdTW6JM3Z6E8tCmb+h5tLu4tuqpeU2U6eGSYDKkxRW4d8mjaTb0/xrTSAMK
YpgkIfKfeCzI51qaoKHPT7M+sp5k9nXFbZocGQsWr859Y/YacFhKkxu8TTXL
cb2xuDebea43gPOGiQDy9IdeyZWAF3YX0ozQgoeuiF6NgGryAIhn9jnkLvw0
1tLAImCEDFbtqgM/XIx+YPWY88Up6Fr6yUHrK6N4vgwXmz8Qq8cypmMP96Oq
W/ttr/+/z5fZcjDcJvQJMtQ7O1fRzmdGwSl3Q75GvbpWEe2LW6D8k/bT6+jh
c7CeTZDIvCtcQIG8FnlavuOkr287Ntvwfp+oqloBwEJ58BS/iTjry/7x1SA0
Hs7OnmOan4SPGdojjSTCcsoR/HJND6A3ZxFhKlm/S0e97KfowrCIo1sYGQFn
VZB0dkwebHb66pLTxyZQRBnhBoLjXoPSugqqGMBKr4whqAMhgfAiuy5ZKclp
yxCE1eAYTATqUPV6vgVQEYDtWjOWMat1cVJB0k1hacOYB9RVIjrXz6mH4cSh
XRDurm6xakxGf9x2R7BRRrIAWqL5ARsRrFQ3uveheAuOI5stO4eeq1GvpeUg
yDsBbBmwmlHGZy/AHpnRFrMDCeiEFA0CedKmmht0XTYC8zB2ZBcYd6yr9A7U
pR5KysAbySfm/P6APfs8LIgqYXoMVv1PPjbzdEQyNYLRU+P0pMipD6Ky2vtU
6fCGZMahk0ZTYFxahUTRWUCcaYyOMbMd90MFLEVPZoZEBiCa/ggWtI/k8sJm
7BHK+fH1TguNGZ2aFvE+vNiYHWZRbnOx4o3rgiabxGnKuPrz9XbbGEx1hPGn
nfbJr9GXukurWos0PgNou799f8NQTIebsVc1w+IfTPDNf/NRJ06WnxeimdWl
ymCvy3Zl790mDlPJQF8XKIHOdm5HWCVLOXaZ/nFwvaNcO4w70Iqs2cJlM/he
cpmSEkAtsFM9XWW8+DJy2sMKh9fHpV/HYUu/Nzpp9s1sefVnlU8SandP9fv8
jm6KXAo2JG9iUw2nG8lgveE1movOqeg5hp1093UmmPd8K51zdPRpdQIjmMIM
6BYCz+YfM/k/cHjfBuE1eEcKD8u0l34ZaurtqfwqjvDtBsmIzci2gWW1dK20
U0YxEsbrBuAJLhGnbasHYPF0ww/8Bq3g6sbovGoYC/CM4Xh4wmLwcWbZORlG
JRke+YulbAVsjqf7+WKlk/qcuo997FhmOT7cY2xlfySOvnl5znfmY5amdGVR
8uBocWWO9z/3mO7Jsq6qyYmlO97KiQ9ZJYe7uZQbTEupFxinWvuMeUpFMOgF
HFLsGfcHVPKvlknmrgb3Na8PhMaZH9pw669+IW6/7/uWNg3G/MRTX3fBedOR
FIOo9N8EjNe/CpkcupEmkVpC9/hSVp2mgZmufoZH2wYkpPABLzZKPDWcmw5w
7JB7ebz7ninT3EzPf/+ltYT0wCZIZnmSvo6bRAsUZI3nO60Hnd6gccK+ZsQi
8VHNDMw7vXfxw+vMp2hU0CaYTRCyKWnNZzjFc6EtprWdW/Wm7L14gbHs1azo
dIjryLiblMVnxI91KOuC1TDwfWhPs2iv5OBuNAvtJGNJeYJQmRH+sCGPqvWI
JSnd3dYkdOnCGZkt64GI8YeVR/Fz5NUhhg5xx8OhTJBqF431VPaKhHoj9BtJ
e+UVlxLY7HZoJF0E+gezu1az5Yfr4zACw9weh6hY3+HBqDLE9RmknKgTN0co
Zg7p9ubd+6Ws6Lmo51BItW914B+0oHRgHT/2iA0+FZnNyR6FnjnWi/N6hZgS
ckUXyy8Jqdz+8oBt6UD3ZFJu0gn+NaL6e2VjedkA1t8l5rFM6cTdMWe6kruE
BLoRtL+XIfgn/cqrv6MWDonHYXuvEydSyGJUl0Xx/J4X9akvZwtcRHMk3no0
2wOyLsqDRcJBvt2I2N/oY9y+y/RuRGWd74BDPqbsNjD47uEOloI4/fvvn9Xw
vSIW8l08DkIl/dDGfCs14j3Ln3t+0Civuz6PMukf2WdgS9BAasSpRDpwc+1s
mxog95IEHDSRlhNUD3U+Kwnv9uZjKA/1MOZkNWI9fW2jTuoIVC3MX2axjaQu
ab7P1ul3mS3qkc/zhp/tyjHKjzaWKEC6ARa6tj1P7mEMpHb5pKsIgyaKplYx
+OMfLQHgmGvk+S9tpWyS4lCDy4pY77/vs18Vb+psKF4To1x9Y2aO1JjxvEpl
baQtNrPhQqMCDYGYvQCyl3epFjmgZvj0zCuuwJHeOYnXOa0+pZeKo/PQ2wzg
RCR2JZo2yXO9+jsLmv9kWtbO0NTAZV1b7lC1IObtF3pyyP51ns8d5aiyCQy4
v/Vl+CJ/vHq0sOqy3eYKW2qd7HkUNQ4IJBF/VU9iZgAA1nrLjxbKYN5PM5YB
6PHXTxRHbzWlmyUjzJdGA2FVgAlQFvLW5YTxJKN2glgS3yFkUnCA1KyDTvS8
MIoYKkyXAWHTnuMWD57CJtWePXq12ygE8hHqAqtait2EHagXvWBIAeWVGJCm
wWyefhAaVQMAhWWwHAvC7Ufu8FfF+WIs/zj4El4e/m/GG8TPSgKqH2rkD9Zh
jzeP+zvgjTVLQC4Y++gV2g4XTTjMxDgWryQkHU1SHxB8/GpBFcswl5LWV4LZ
5Y1kHEe2DFTJ9xcjBpdJBKXoJH8ecsAYdWrw5QtPbVUO96H/FqvFnBlElI43
giWgS9pIyhXwjQkR1C89sGhhsYZliBx3NN0lcsAlMCMWI3XX5zs8dBmblHGS
AF2LivK/cdl5Cq+QkQwYDsJ1ck5eivm1ySdCvkNDyHtPX1dG1O3yLb/d53Ka
ByuCiTDxqMVB2B7qHSHcvTzdtV6Y41TyTFIEWirHs1w7GhEHD6pRPbFWeLcO
XYmSwr4O+EqwtYqI1xKv+NqD0sNh4Tc/PPo1MTcFM4s+dLFPpp4z9V5COazl
ZgGKuZufZQD+UMJ23tB1viNMG6Ipl4y76THcTL00x79Fpddh70yWzhfAPh7L
blrKgZ0XnPEtrTU31oMXaInyPeRErSWHynT881JjgxwjgEDXS673ix7c4JMl
k+K7cZFIdofZN/A0lavUBv6rifvsbVYIfNjdf0V33T2Mz9A8H4m46PozwGRh
8hqDULOKklSJ2m+IWAf+1z6/UZ495T/033HavHUS4bRmnjFT+yAjHA79gSRH
dh8JxW7hGUfd5HU+uBevcEGXAoJCuLS3JbuXVQ23IGx4bgA6DWBuyJSfdHD5
rQv3Inowrg8if09ExsihPXkDTZ+Mb9mtGoBn6EuDssMqyTT3HnJjOH0p91gv
6yZcN2co4xwA1fpV5hxEi0wdYh7xTVhKGyqoHX2AbESb8Mw/SB6WGfbso+Z2
EMowLBaOPULaiez8qJCnAvx5EluSix6RJpACTGqghzm4XGXxHifgH8Vux80K
fKZGChlGVqStQoLvcmqLVCJqH3x/+m0MqazIOLyjDZ3QZw54D8ydwEAWc8/Q
2Yw7/jgJvNMqHPEZawWrkn9dYg5niAfDLBbr27O7X6pg5QjLmVcuN2K7sign
N51Idc2LBQ/y6QYIQYV83fJRAAbEiMdr38ApyaN/Ao4sipXfAlj0RMM+pCD8
nrucSsNhd8d2pAYBzoYGD7WN6ssMs2KiCsRZ5OFoyXgQcvuXy3IK6RpKXqLR
Q5rzMPCWHNBEKpdSH5/393zFD1+eVJVebxY5IdUgYNgD1W1mPdT4j8WCxz1+
1KKraowc+kF7HB1hpLhT9QgU9qD/tu2AIF1qMpJmSd8BvVoBPnYiONcvjsLx
CeoSIJ5R3tY45BrOixfJL08rezCpzpGExm/N/Xt0j6nLDcbJbgWdGqifUAea
It70j2YtQqzn71/Z6vuoPVt7N6QDjNMkOeQWY8/6RhVPf+bulPh4a6xRVTHW
qYYwvfXhuSU8hKqCiu/Mi6Hf6Ce1GOrAE+re2FQMi97Y8f01OWkKhyAdDPyY
meVWEcsQC90GXA/AIG5//DMJckXD9D/YXn0I0MttxbfknUSXfPJ0BbRDLAI1
53NfXb9sFllTSxJW6Vf5/5Qu8+d95520HeKj3HRTc1TSZhcqpQYL9XuMJgJ0
R0lkeFlrtYEYXAt3G9SdmpJGHu9gxWPmTBG9YtTGpa+FDGbJLBXv/eeKjnAh
8K8yLreh4bIEXIcdYmfq9GgzfbcHi+fR0iYVwvv9zfLFMXH2FmQbYY1WMqSE
DLHI04JY0WzDLSPfo3QmnemhfF0Rk0C0OjYtBzfepvGcLwQDJrSjVsPmR2Zs
4z1CcVa+P/FQ0Wap+GuTT2ks/DZnjrUja5+0Sw/oHASgMg2lckFEiMZLFA+n
Mq3SqTPI03qqbIHQm6CYCpMPhAO1GBD6APZdqd2L/iuJIp/M1+9GtHCCJDBu
gOzhCMZGY2wJW3lMIQBm9XWF5fGsKlFSNiynAwq2TGsA4hHOyyUgJngAKHe/
ww4ucvB3HLw17mp4fjxeCbBzghpY8I2A+TIhH0e3/twu2XjIRcQb/GLRF30q
QbewyAt5njis3iAQHz74uBDrrjKJvtbU9xzt33iO58TxT10czcbDa1jXlrMT
Io+EpjlmR3Fmm9YoBIo0n9+ybTV7L8oXLUej0iiaUOT0BD6PNHj71PEtEKrV
VefP4SmS5tIas57AWTap9oac9HRiJsQwzkd8jcHDrYm44MMjBEVJ9KBAPPe9
2H3CgIf9p79phOVWii7Hq+9+1P2wYhzQsGf8rSXl8pUMFZDXLVNI6mzFahKL
dniiV5JkF8unMTqmxwAASPl7Gir0snIiMGC8K3incno/f8B3r3NkFganK1bG
5IeQQ2pQR49Mu7zn9FlVa9qfRm1Oe+vBbf5RnsLNphzU+OV3WfoPL3OhGvzz
Ipv0AZlJbRdye6sGyBwVbZ/n+m2GdvKou511J0NlytWIaaYwwKWhJacL5pXp
xV6zWLlwFNIFc8IFWK4QIeGYFAzpu7WQdH+s5xRuW2O/CdG6qqoGnQNO7gAs
8igd/9oNIH0QGwuqbF02nLol2jhrKai8XvrNEI6O0mfOdVchUTuSoJt/ReRi
ADhIn3yvTvcsmFBzVpipYfuvfoW4YddJ57BOZuh31hHnxeduWZaFOjV02N/s
3bXcgfn1XOq4WQ+H80LoQ6Seo4XbNFWjFVntvYlr9uSHeq2N8mKmBS43BYXv
M3k6Ye9q4ymjjJHx/jNJCptPPhC1Y8U291g9W82w8KeEx6hHe2i217s6DQ5p
ytyOJyXsdM/s9Fcsz/HlgevZ7guQGG0sSjHmHC2SpPqdJZ0e/Y/hG4h/l3u3
dNxKU1U8GTJFO/cTOM+sL/JB86Xrsgveff3fi3h+oSsCYlCC16CfiO4C7s9I
U9eqhG2Vg5LXxjboNAwV9a4IHklDxDVUeL9C9HMKzWItXXQBu25hA8bWGz69
TSvyZCmvaoKGsu4UT2TvYvt0AYUBDtFBW1bmX4PgPkbbqs1sc0/oTwWx4t9v
RE0/DN+kvvlbFfS4u6AevqhYcAaNWDyHX/mA2sRXA3tt/Lr895pMS/TNft69
BgoI8q0bJmjL4EPgps47TM4+kXgqx/xNwH0gpiQs9gaSxSAYyRHY7oswX/kv
1pIbWW2U5+knsx7j3BFxULkkkDdHdr5Y+SXh/dPfmOJsbwJC3zf0RtmQeIAj
5LY+lG9ZsfzVwsYizFadpbt1KKL8XEPolPRR/6Y48KJl9AMFEthhPgs4WcBA
8pt8e8LtBAZO9Kaq/0D1PlVz7itqf36M+peKMcze3MkgvNqAlgysGjfkyz1a
Lt3AvfQ1Yy7T0EK/EcMwym5aXetl6Y9i6TgGE5/T42Rw5gXZ5xw2+KCkj5zY
pxuXVPlzpaAn0WUMwDKJVB10YAba0eB4S/ZJFy3ivqB2hAwnT20UYTuBHblk
zSR9Sepu8v8S1FKRicDMSnDJRAz5xXl4JYt3r2ik7IKRISTDGHj8xu7jGaaA
dtBfxBbrV+vIO5TzrehGrtoR1av2nVEnI1OL1harwM8EzhG0FTocA2C9ybXt
uh2KIWk0vsjF69ZmyEiAFMRKHG9V01+vCIWY3BTzD/hsQZuUJf2tc0MJbtKe
HTwT4UvWog+VaX0YTlOBmbTPqPtdIHs8cuVZpW/lem3UTSSig4XNjDnvpo73
Avf/bxsDIuReIib+CXm5zmZDG/VYY497/nqFw/eBUyVgDQ9AsDm3U/CuuBb3
kw1gVTRualawRjNhQBsE8R1ZmnBgrWHLmT332g36qKWpp9b+sffdyyo1ZkS2
q+hXLkxy/58m+H/10b6DMjJdaiNwpEWPugHJWQgD2XtPCXxKzBvyAqett2O8
jzF8C8xkXq+N86kUp/rNtm2aTImYHEprvoGyy/TZq3csDhUwji3ZGCLbGfyq
wVGqa09fQZgwcgIHOCYACDiXt407z5jZ19sEB8pNhDvAWF3oDzFlu8UOppPP
I4cxVeHeRfEeRpMUNRchZD0zsDnky/SgZoV7miT/2kjkorI6IES81X93cBnB
MEgyFg4PApgcDInhL3ZcFSFQqwLTQxc5ZbDhYk9MEP+MhBhOfidEpBri//vc
37u2uxB8FTqDBxb2T3ahQoEKh6NusBHShTQ2Em2wq2MkVWSgGkNdN6k5lDzE
kUj1dqGfOEhYhnN6+7zz4yfrYiEcDVsxLdX5I9wz5tDCw85Po9xii1UpfA5T
wmFapkvszbYnfwD4/7gevbKrxRrzL/4DfwcE+JP8QzH5XQjvbSpZL+/Y51SY
e44x4C1JMhDmVeAYT6rROtRXvtgY0r1MnZsugtxaUP/bShI9DZh3+xZn1MlJ
f8rjZ+i0u5ku8qGFXC22v3w8JALOcxf2RePS8faS2t32vZDfOhwT+QIaKfa0
TGRMkuB2imSPkQg6K0KuzFwxYvz6qpsq7KLM5XQB1ubQ6mkxAqc2rYrhgQmd
7phTcShSNHedjAFF+BJwnIlRT5JW/QYYI0sOliznQIyiKRXypi5rhBhHqwug
4Xsr2LE0o91txZraKAHfMyq/FvrqVyrXPAs/xIm/FepfToVONDaaJ6K5nr3e
B6h98n9ruuaGuRC1pxc0HJiH+ku46JglY4dBCouTMkQkf0zkGUf9fzhGyU5z
idcr1/tXuvmdnrJbT9JgQ3QE4eXfqW2wxZEP6IG9mh6cV/VlBUrPkykF32u3
OUphvxbtq/5lg1xDtHjM1tXTj6bT6Th0yGudtkgTOM549/jK23zN8D1gc77C
K6gPQEY8VZbsP07FGm8QviuepUJzH+bBY3/5bosuzUcyhgSWZZu7NMZsuaPs
16w+4a/huVmB6v9nhJJMexfU2AG4KKl8MjJmJFDS+KBj7V0EuNvl+uzc6KWR
6HQKrUJ9/OeAaRVbL32leZzbvPprgSiLmdOmBsRlAwG/MHuQR0evwO/qFdLF
HN0pTnGxNwm8Z6cJ5wIwgyLWSu8wC6/cVZJiBqFJ5pbzzdv9YlWcPWk+es/n
VIvK5ssBb+9VUJc1HOYWmDItdbtzW6usno9SD3v2wIvW6qVDbrTAQ5rXZ9vZ
vKlWUTBdTYuYM2W0kS0yV2bVMSRdDt4qgtYBvpFjWIfAiswNBVEYDyNhDXBt
JENh4yZdVGtioI8jyUsTpnG54i/kwpTiTkFcdwXci3loSiXEEkxMxg/bUYxH
8+MR4oyWF3ayM13Yo66tRbP4BjtJmicLlj2aTSE3cWeQBlcopyc25j1ax5aI
tp4crTEDsJ8/4PZIpibHnjwcWtYP96oCvIcLSRK9RL/AEvjy2V3xLXbQJbSO
/bDDXe/Ae7V3T2jrAfkdWgp/lLt+aHuceK8+V+QWZf01Wy0EztJbjQTgwlgf
AFpqKWUXuAqN4cWXQ+zvUVQvSCFyvMp92w5mDHo09q7UMKUL3e4Nr4yR3SZB
SwiubnC9e8d1b3FNBXNg2J/3MEWF3tRwvHvQvlSbitLpXfVDvzeNYBWy/UZw
IyJWQAYAOiqh0fw6sXmjRC3g3O+l8rhM0VOMwckc7z0ee+x7aMoKMly8Gu5u
ebkFFT0gpQPfTDdbUm89CW7nSPx0R5hha4c5iK+Fehcar07TYk8Jlndar+3r
CAcgOHoM2M4EwzXsmAXuW4AQdgps4XveHd3Rz89mhSZouuLPjLG3yZDcR2jF
abX2J2jhwr7+xkshff7qrjGaiL+giCXGiE3Gwszu7aL4nWZWYm0UBeey8kBv
HpJokCEALgYmHQfVnT4pdza6PfhXfHbrWJV0P4qla17RljdzCGgOCwiCETcr
/hZusD8A7syfD80NLaFhnvVn+wZdIB7LX9PKSejkEmH7rw5foueukoeKveOH
rNNsbFmDzguE8V558KmtzDSLt2emgPVYeDfIo8yoaShtR2ZomPI5iafT0M2l
Oi/yu8E0vqwyv3iC4gwB0J+B50GGVqqn5BWBS06BkLmbd/6vCN+OvaHNkE7V
X5pRELikf/jDmY3SEaQuv+PB+LysLArR+lU1isqOCOolrGwo0putwpPTbcf/
jaojmz2qBj6bHqywKxccYzqp78qL8QsMa1hUYHRh7y9aS8piKA5w5PByxneq
e13rX7HHGdwDyxmULQ3+J8bGHBS1B2r4EOaxiuNBN37vcdPcTGgGVIqT72t4
jiYTDfs7lzL/ip7mantW6M8fGq1YxjumLAzavRHE+KUn5Dg1YwYt67px1cZc
NIQn7Ndo2rY0ANGZ+HYyPcOPMQbYSVow8JHNcMtgw64BnGQoU5tmEfYgj8u7
ZR1T4zetsUDWKowB8+SdDwltM6pgO/4TXZZ23B6CxHIy6IBXrZUtTrsgy1g5
6/xNu2FoFIhzzbyAiVX6UAZZeQjt18nOg8ShmuNzTqje1gG3S0CaX2Xpd4hl
bVpdRLUUAYTmwA9xGUFvXOlBkFHyiE46Qb6RCFXWPc0VluhRMVh3n8L3BEjN
BgmvD+0U2z4jzpeVokwAzpJWjD/iOpPfGZCHoh2e2+fjKz+NaK7OEuKqSpOs
mm0U8qP2/bnCdYbRyRVo44M1HGNR2sxIQ51JnKYXfmwP2HRpB73HzdAAvnbd
hYALHbiqdJ14dXN7E7nJhfwJO9kz7tp/qkRBfEoYTAZzHktoIlAwGULAFrB/
I6RkdQVYK0hki2o/jADuPv/IXAl7KTDtEVB+vj2apdPNWKNeNgGs633XGN/r
7vVRIxE5t8+ODRm4uD+i9Uy7CUJm7yv579eE0uFAtoxL+u4DXnkMc7mnw0Bu
/otOaLPC9mwIOmVkmf6xt48Hp43FvJM2q5SbvVy+bVlImtRjiqoG3lqfx1Pe
PzCLgZ+vJMuSwiAby9RHiqqNB5kALhfLo92ZGfHy/Us4LAGeUzLkWJrs7rIn
uGsPT9+KVSNDQ6o+pYaqFmcM2RMuqkXU3xvVoObBTBabuf9Au9o4GTnEmkdo
mrYm9ObM2xNCA2ZKSTh+g8fPYJBTlOXG+VorBEbqsCXISDNwG5JXqoFjCX5T
iTT9XNHE6PkbD7rVrgGp9aXuzDjPgdsH/0w2/rjPvbz+Xzr7xPfXfD4W/Os6
n9WHvVX8OCujE1zPvawiDQspamEzwyGHXSrIQ9bOh+iXkod5F9PQiNirnsYq
Q5Wf86rLoXmf0B8QNU97OsVPXIZ7Uqv6pkrW7ofTvqTk3vLlDkeD4vRJgAXX
+UnfMZYftU7wbV1FPHAIfeWXBZaOZkhbRJVVmLg6hbuUqoBvd0iB9G8ryAso
33x2Q2lXN2Ju241m9XzytBgMbJddcfvwt67S9RfAi8Zij1TPvSgAEhoBjWGf
MqhZyutcYMKhUy1U7W7srn+UOmnEMagu2TrHjSkj7Cv6xjt6pZhCwlIDpA4V
Tzj7TjrqyjPh4Y59veR28KzdYIT9E4ldRrg9vUUig+EFa3f/0WUtKxbHCdXB
Z8S5Qt4qtMAEKuZOUzG+EWFLg3iTYiYWSRnPily0sjdSx/iiF6QNCuvc6mBz
yaq0VNoEn1GbFJf60Sltp7tejFn55hPu5KtK6Nah7NzTxf0BPn9M0o/ZiVi2
FH6rU59mgM91yvPx8CURPe0qfva7O63fn70I7SB4acXozFwJIcD5RN5WYRvD
M/rnbfYXtkTmDHanb/4e4+fqKA1PpcrOZ/bGzuc8HW6ssVNrMEEmtkBxlg1q
4rOVAo5OGWEmgl1oCjqkRlPo3YohJlZXxBnAQExbvwV6y1MmJGngQqMUZGg8
bqgdnXJ5Oe9rFj3NxWNuwNbMK4CThCIqxg3sGICAjxlU6QwqIznIXA0PuCoq
MNQFJPvJKhG4MihcV5IWxZefDb2Nn+YKF120v45V7oZVqy51QrYmxe1a4vGS
gK+g2Wl7+M8BuULXege5vXK5u7+Z/SGJD0WVPyJSrkxwXP5VZ97Mph21BIyM
7j2xOxwwvBPvvsozmEI1+krMU+ME1t1b4jSR4NC0o77ywUW9lFWD3rCHAE+3
YbSkXSihMnQqGO48mTuS1Pk9HiaM6710ldiP+Pk//FYTirpBhOit2+Id+Z2Z
0yXN0z3wGCp7lZg8JNVnEQs7PuaOqI8Tv8BuuQXBZh/1AWYSrFgt7rJpSmra
h2uTbkLYJ3s2NCDp/pQddDkBHS0pCVQsWionVJMBhSfRwsah3tbEMzxAwecs
tqhI/1IQC8YOyChTJTT3rizySyKb2aJb8cq9mpz2OJrQLgIUQh+KwFHDTWj/
4nP2cmoauildVwfcpdgMk3JTqqP+CkLoJaGVBEb2Ig9LUpdOsI1iKDcugRHf
m298nvsi5h9G+tX47fqCQoNIUgHsXZmXZwhUTfGlbjrkySLCOV4R9COASAoC
wqIFy3xKyjEC8/iNb0K0o3ioFxhEAb5KO7/IYsqhxPpGvDOSnjFSNuQZNO06
fp0ss/bhqPac/kGyYAvJgTwrg0IkwRZBAxmjYiBIWAsvG69pblD752M6EcI9
2e8qgoBMu/1tHe1EUA/3LPOwoGLNr0EhmiW907jOgH69817mMk5hlmgXYi50
cQ5ZlISJxL68w6MrYIFZ/rJGIv1hz60UttnPT9aHIZPF73hROp9IkJx3mJbZ
Zc6mj5M0CRjvTojCI/G08AXKSTL8+8tBI0s7+KDZ76iLIaBKP6dkcAk5G1SA
MUPnFQHYfTEPZxeSdur0ZyUo41SnA0Jwb/0ooFdgOA3PaCFyiNl4OvYjJcHB
c5WL1iO2wwLcfaAB6dL6c0icnnYhhLtHdowURhhsx6jPlWPGYg2xqrgmob4M
vm2kXnx+sWY6fEJQN8CHbuukFTXFioLPCIhva7M/JF3nOARhITGplWGMZJPh
h8blQLMXdQp6jNlXIhNGLv0tg5JaEVeZWcyZQ3rzfrkrwiYBd4ENL2ZIyH/V
MnSUQ0/9EDLQzuO/P8QyzTOFDbglk7aS9+eOYXKaUb0R8VHRwHFZSyQx830Y
qN/5l52A6pedGPDH4xCBqWxjyNakmegMNS+InEkpyqXsXZvXOZOFkKwSjBuv
Rpk9oCC7kNTV8bf6xORzONvfTijd9nrd0pyacP0i2ab/IkTh1pjL+1PBEf3W
ZgE3shYOy/R+MaTpAmERswtJMtBK4kl+v+HPmtiUvQG4HpYwujco/pb2lLpl
H28X5uvBSkspsogXLNrpWN6rh+P1Ax/qH6OhcnDZ4+iRy8Typy1Cj3u8ezLQ
Ciumpyj2HV6/BsSi/qQhd5OTBRgrfK/cFoxEM8q9D0dgVe3wpMuVWMsy/i4L
Ii/Cw+BYfMk+eziT6EvNXr64PeBKAJfQjy/Spkx7Hcdfz7MKHY/LDlgDZZ8M
C2GHMD9GLXoSc6oBFnvXpz5DaXQKR3+yXfchj5weAk2AsdVlf2dg7X0UeZxh
1NlhlwAY+gesrJS4rEg8BXKcgdDzhDZL4RzYNZIkT//h3vVSyzEdu6WkrQdw
Q58lc4aLkQ747KCSRGUMAGxNWyD29CjpzsAVQweY9HHbLC6/LsAEnh5HH78D
tFraW0jhPA87VXcLBXxbwZCO0Th0fVnagTL7u0GKRBLYke11MVWEnpEMiqwc
7yVA/EUnxEJjGXN7fFj9XoVX5t1cbxQnJnvdCb4WzGAQHCCchjlmDBhQOu1a
F9U96c13qdh2cfMdEpKhNtt6R1cMPTJUIF90Lz5AkvHnrm8YqAmUQ+abXDFe
Wdr3qkD6tEUdkQfjLcQvuTtqdsAMBoDFbj3pSq58cjafl9V4mSyIXmRhXUai
gahzutLNkhxYqFSm7kY4Y/36v24Av1dyySXzEBiOHaaeVP2HkrtA1RJUY5Nj
XDJVVFVq8upBJa4KHVcCDr0OCReWOCuYE9CydqmhiaGijZDqeCIXW4ZJ+eQT
2sf47uzVg0wxHiEIFZVDqV60nrhItMeq8c5+jykxphVePexhacMpnkEk6ZCt
LjyiCobeEKv0OyRzqPGjZT5KthfroahhT1U1PR8aoK3wxn8v0ljSUhhcbL14
4N5Q7+TFSGfdFfud4ugTL1S656DjqoOyTFK2DqmazcfPiiQecRqSslwtUN+C
K8KUprrsn8MWkB5Vd4jPFNrCWcs6P+Mksq5oN/6wBTgD/XINWCtWcH3uub95
2RHdn/mjN89tscfQaquKMD2h6D7NY1yhwsVkgi/Loi88974EYmQ6TkOVe0WF
HRldbEKMa3nuDEOBmElARQiDUemAD1Y2Fdt0mpBVdhOiXsk4pOwS60b/bJ7K
XGHY8wZ9yrmKhJTbtT4hND6YrWRvopqoOmR0vLo++mNUbu04K7Y8BUSmbGYf
W0PRjnoo2YT7ErOaevMIsxw4uvqxDTI3FTulSxZ1Ds6Gl4VlKgkfZrNTpimf
xImSojyDQrGeU1ag0LcOrGLZAd9A1hgWlPb8FLPsLNBLAu3TEjmoYrY++S5f
LzCsTInf61wEji8gxC8VG1hDJ6iah/JzTdEKZc/muMrdBjPF+GrCUSyzrgIk
Xv/j7N0+mGDya7GwMtbgcOOL+uf0+Nzw1aylGSApiC9SCQNYVEk5uJ+QRcOB
Z/a2X7xlWQzPug1x6LGKLzuTFjD0m8EAmJF6EJ7V3mx7gZC+gN36wJwVDNNJ
Vd3wKGPiGU21qZpOrIir/M5cowB6H6OLoRv/e77vhWBUvlBB0EjZUO3VaDiA
4PdogbibPnvw8y5Rxv33Wa+6nH4OB4JhsCc8i8n8akSlea9SE5nunYGuN5lD
/ZeEej/02R856WmGGl8mrb0zEAesebk79k4JV4rax/aaLhRh2FZdnp12o/wT
fEevLoVf0tWRWR8lwj9QTNoPUUH3UqrM8ASF9aLQAAoIvKvAWF9R9oosG1LS
z87rc+jOuEDnpPktcu1+42urMRJBIbG5l/ZX1JBmXV78xGLCFS36SCdbY3K+
KHqpI3Wv+vBGptAukBkL5pDAWInpzbWqshezfc4TM9qDxfHsKN8lGnIm8gEa
lH3PN1Ze+qbsKwxpJzLugT+RIwJ7LjVgi8s5Xvf/+X/Jou9SK2pPMegBdhrq
3j3Jb/5svxmLsvA2Wxd5aludBtGdwnL6V76SRnCCITNTB5984zofwwNvnPhR
fR9aKk9oeM2y26CbuFw2m2vuR/Ly+mupM9mfWw1kV2YiplphT50v1tCgin3z
7ABi+ayAA9PSn3QjDB/FmR9FkpcTvZwkaqzTD+bpbCU30G7Y2fkGp5pdJG71
oLHLaw/thdngbWK44CU3mFcneERc759N0Ike/WoVC88+C9el8Zy2iz+EO/7s
oyn1bM1Vzwh56TKHBTk2huyU18wsqti9rSMzpmxiya+YhDgZaEAlyhWJeOvQ
OkHJVM7ydIAAht1p+RzfEKJ2QOQzhYAWk8WBl/6Im4jTlUqJ71sbUO07q3y2
KQU8iSHKzajVRe8xYIlNwhgRk5v1QepaX/vNf8JFu670IM6gb02NabSwC2ZK
eYFE3Uibczb42ouPjGzLuAuHvA/Vyxf3PNVVwM+IiEijHA7IWUc276ATXW3m
pXSd6/4IjDxd/JsagIS8+XlTkHMbXUQIPCrc1E2hcfTqgl0+FcDJwG09w22+
1feOty6icSW2R96/V9xYog3LU9H+XgJfX0MVQLfY6gBXUIJoHFdY1brAGvEQ
/CWRotwz8YuyKH7QkDThe+mMuEAJNyqOkxWsgWYtR0RomcW3EqimrX8RWwE7
mmoUbP/RS9tFHxijs+i9WKjNwNkJQLz2QHMRHttaP0GLa8OK9mZd04CQT1bq
yiso+ZaW6c4u5pgv4EEUsV8g++opFRjDARRglwf7cx65vEw0FbXFjPiUpJDY
hjhUXRK0pzYe4NZ6XRVFBIIDvHo/WcNIGXc6K+IQl3Do8Gl8bbW+lJIBFbEW
qPjYE8QpueGyTty3StleqJSSZH+dXTkb5dr7djvimC06XeJXVAXJYv95Y8WG
hSChsuvA6u8gpFH4mbBMAgCVENgSOWKUaj1bcqkW+UnafjLkHp7hbFTGBP1B
1mnEpGWAcBNev0NDUV80sIcjK4RXQPhZOFGTFKZ5/3E2wI1TP3NJagXc70F3
16n21Uh5yt8ME0pCXQhbeCiFafEH1LvvyKLKLTQR81dvyQWy8b6UCwPFKl1x
qq9cr76PKOrQQT9jpJ2fBe5EtzzYjksSx6R/9zywmD8v1BONTnndWVpSGxLs
QTraEEtK3xmjh4FAIj6kdSszknn+tCuQX6rHD92Xv4r3YD6N7U9hAHUya+fJ
2gMrByaV15L9g8oOfHeGdP37YFe3Bu3bAl1W7/7eskpQAa1RWgT0S9guGHy6
VU3hrsSBXpbdaxQHVJUaDKgK9vtu3yIRTAKZ6Dbivm5gYeChvuPIcRbQq1wc
aoo1MYF1L6HZIdagBDD4JqJp0d0BcSuiJGby1clKqa2bROU7PkiIj/Fd/muX
odJ+4LXSIE7PCm6sZSz0iplf/KUFhnkKWboB5yErONpKOz0sCJsgr24w60uY
JRoFyB7v+hMYhpoz8BPOkIhni+HgGygVpu8L0qvQ//TTaLtxe87Dpux68uqG
1XOp+BWkF5EK0JGX8C0sF3dwa3SjI2/q5cjaQ4KyHjFvUGewal/XkQ8Ad1Cj
LgE4YhojOz7NFdvp/r/qZaGOe+iqMAxIfKcWYlTw8USBwvKGobNf5sD0ZCls
uIPmZc0DGNhzT35i/8Y1hB6sDkXbLionLJloTqkqE/F1Bmomivu8CcwnoSE/
wSIJtNe16VRh9K2MMFM6g9qBuvC2EzTUxP/8sfnfg+rENmWSgZaq2Sroh4yB
MqtOQ55xxwLex4tnQhvGHZSFv9ReVUtPz46/IuaOwWLK5cM0bCJumB6R4DYv
rnPOY+NzokMp5xsW4HPatDSfT6lIPOz7oi+3L4EqOImutPHTz1o20eYkIc3w
k8z+e18UANF7VpxXroJz14pNvd0Tuv/le6ZLNMisHhR3XzGHUHJK42IlMVcL
We2ugkoiC3cRBwIBnwxVw+fOQvHJFqF8sWZSBquwcYJd/qwO3YMTVuwcpg3W
ijvxhG8pULyAqZmwkOThcTyVhYsoKjHweUuRZBeZKxpE9fDYxxkFE8XfwQuN
PD/28hf6qQtcOfniiOoauc75U5f49qrM65PFu2dnsBcmrYSfLMEPQPpX3UjJ
O07NPqKSFzcKy8Bl1kyatXU1cM10uHp6oOLOSX7FXGPW1bMcI7qUuu3370ti
l0fYGABSSxqqfCgtFeI15oE11MCXdO2TKBFTxDGDlLC96DGOewKhZ0fOcYr9
i1fPtxAWbjbzoAQFHgLXxxCJ+0Slru+Cm3Ff9WD6Zbe65F9GZyKwY+JWcl9P
vbzdY89pxGt5rDSs3CEkAeql0T1pjp0qb3IVfrOKZYj1XRAj+RKt2hwV9K+4
DIdhFLOWSJzlIIXiwLlFM1xvS5TeIvNZp7YO8zECugFnxNxkBiaceS9GaqFx
tCiNTQiTRzI0hviq8SPwCHwg/CNTuuorMnT+33q4xhSWDA2cZ465cj9YDJ+z
MTXr2g1tGyiffzUC3ZfM2Mb6B1b/yQ7sA+tolTVTkUeCovVO4PQYaG5f2k8X
QnpLO0PieAOXQ3vAbpe/9JdRMtWa4qOv/8yAxfBWxgvrtdYeLMyYHdRd+uP9
LrJxXvCyIQLXh/f03uw9PetO0EtpoIDxfg2661MZTepnGZjyhyMoyrCeKKQo
dxtdWekpOlftDXJ5Jmuw4f4GyPnTlcjnffOl/kF94bYeIGGQ64M9dFQcBLQO
0YZteLkoqPPPObRcqnHptvK7DR/V+P+Tf7X1r1p7RzfTk395h4nTodr4jtcS
W3SkyrVWib5NKZnvBrg3q4S8+oF3/OOeY3dU4XwVa+SGEfE7ONw8JnL+kEkB
NYAQTfpcNahRnJ60k68jVOd1E6U9qFmFxog6Oseikiozj68HcUd+w6kTUmNj
9qD7Q3rPK3qiuxaKYoK6EfpZVA/T7r5tId8zMuC9O93zCHVwagmT8wtEqax/
pk5jfdEsgvhMm5V6OVTatRNXaMP4azAu8FJOBlQw6EePKpBi6GR1WU34U5WM
AjWoZyIkwjM9sjHlGWtk514i+hwnzBJlDYyGG/0cuSwYJ0JvYmwitMhGrrLy
CqBO+kfl4wl1eCbh7CUg3JxcvWyTsGJ3LrC3lbA0xPQpYut6e0BH0NvWNip7
WnhvyWuVD1RyVRNqSJybqVA5rkgqMotwCPslh5782EfoAzArKJcCheU/0e9N
6fT1ZrfQKKZjg6bg8Ejksz39FISjK+nuqoNBGGxEtQd/xyybptWEffsz2iaM
czdeA6F77ZysYi4ej6mYqmxET9lq0AqUHtuXVqfo7BnVthp6Aii60Jl+8E+h
52GRystKobL8s4yo8R+R7lU4LB4So6IykclltgFVRB5JG9kl5PaFFWV+FgOs
OzWTlbux+r1QIv1vjcZvq+opNAYVxBeFat7+Bt/avA205DX9kssdwN8FQQCI
rso5BC2B9mKoRpBAPtrxlRoas3q/VaoGynRh335EOrAtOQDDlktm0BI2rp5g
fhM187SdN435vpDlFKeMPJSIRdJbJle9D/UgkVZrWjMzEdh5+ad+QzlSstrV
RlzpuG/uZxZEFwH1I3kjkBQ3hS7h/DjPDcQJ1hGhdc3gEIHPUfAMbhlb9QqC
fxMtk9x/UDU8D2Yy/Ctz2x83bV751hfJleJ4Y6eEMLzhrNtYJ42c2z9jagXb
EIQ4xyZZXZAQ+SzS73HxHgxCFuOK0pLlsgrKJVBcijnPlBJK6j8q+RoHWlDv
Z5acAnFqsH0qOZxrGc48yrWNW7dsEm19E0VbnOin38IIesaOkiUDwQ7T3LUe
eUbMdr22dZcEB4pkeKJBLP8LIhTRHWSBqpncH2DzOo5I7pi8JMuR0X1j823c
gyws1EhpuIg6FuRbRbeD6fiWyFgr1qSWQ3g3hSyXW5Ctnw2R5QRfbQS9WJC3
mzbgUjtwexN/zbABkPFiQedhkOhTbZIFwRuuV3gLyoR3pZbPGbxmNVumVymd
Pj7h+n6e/DVon7p7Xg9xwyVJl3gNKdvJVJlw2Vo20EzuZqAeH2J7X+5JMswV
7s92l1iOOXqB0m1LGsQCYB5jWbaH4HS3VireV3TGIJEBNi/AsQLBvDyWBGfj
4n1QFfwBXIuYM178hGDX6gTluttnzrE/tGOhnEHWE584uJZeSgEYAIw3f1JR
ErHappZ8sJHYCRfAb9YROb0vuRpwFcMcfFC9M65emNqWICYOjEW1Z/MAAqp2
PzTgaL5jtejMNIL5oBTukai05a67OucTjM9CDYlDkfcX9yn7zRwPHAfmEd6/
IYVHCK0mfNRJM72e5IVHbEdBZ+6BG9SrlMexxn9m4pd5u2If082PY/4cYQYH
bw4s1Ja9LmOrvOvWCYDeMPoqnyJphQ3Qs32H3vLfQj5RM7SAlRySqlHvuiUx
PAa81mdmDFjOomayMXvDrZZw9Dy5h3DsnA5dImzoNmZcAH/Rcd0b+DtXfBFp
5tHlG68Jg3ZFOdimVoOVuEuVcuG14Ma3JyLmVfaJTZx8yExYc16DCaLdb18F
rfvEsJzlmsjoiRXbkMOchBPFD50SQ4xddP3ul25s6IEhewJpdFWR3ZVUOlgK
xlI/ot1wmW4s3oemcRgISO3ET6H8yqyZ2/5lI/B6AVY/AxI7W7lK8pii7O7d
Ueq7QFrbfu/UKI/GUnyNd8wcaiPNpck00Q01ofD1Q+4w/7P32phAXyeysv7E
d4q4a+L4tTcUnZn2+bjN07Nskad4CcsHrpqvMTs3OH+6gofQxFviGUeo++oq
K9J9IhyXfb2detfRC8O3qGkDBVmTP0S7gwwR59s57/UFJiYO6S7ip1Ze6KLD
TZ/VIlHM7b8JFsl69MRq0g3I8m742gDh7f4HbkhwoHpKpUKfyRZOOww3yF9v
YYbTMIXgWvgrwhpV6B+oYsGpnraOn9MguCgyjCEtfYzo0101tySMITTV7P/k
ibFMfJ+MexhlfEovaiGfGAZf3aHQDSe0wTjMGkEFGqMlOGfTdPUIuxWhLxu9
G9NONMQzT+dfEMcknGSuVzSbIIbdreh3I+67mK4x52RhdDaNaAjWt4CM6ruK
F3/rpGiCWG7d5bHbrpjMMXeNkFu9YKhP+XEDeq6EZh+fXY9L9CvEuzxRfIwl
wAhxxOqBTg96r8yWXbZgKMKpFnwjQoWPOa8xKXZi4IwaALAyq2xD4FIvAHWw
+aiIaTDXGlO+lNQd92Wbztv/nW7N4xfDLfPqfHOFrZ4a198VJa4EyLhSRspB
53x99jpaBEE/QYUabaE8EKU7KTmcqz4EwV7b7eV/Mi/du8hR/Opsv1nQsmzB
hwVog5f2QhKDjZTxmn1bakn/UbFpNw8JOYsjm+XIvOqf/5EhCBPN60pacCLV
DwJuzkjRBR+kfgdQv+AsJWK+aRnA0uT5q8CxpKEPzI8PN9cqlUk7GrOU6cBn
gbY4T1koi/duXXMrLuxs1aHFa0hSsxA27t+cQNpUTY7zyqOfN0ce/2Dj8MO5
t9DmVmvIFUHZU+5gABuQWynYNMOa7xgxSgGi17GjhbBoltadQ0sNaOx9xYAo
7V8uQ4pnZAb0GJdOYU8NWqNW7Hxm90ReMYgJWxeyLtYMUr99QTMxwzLRcHWk
XzW2blS3YsyD8yi9mCmDDTBsIIfYz2Cx0NKh9fntNeuhIObfTSinpLtIYnbw
n4AI5m/Fsv9g21OeRbb9Wqh7AhUBeDkFMyQzyajL+3zQg42ZxOcD82x+VNzz
YB00x6/M2XJHSgguOdVG7/YoaW6h0qPIp9YzsXfn8K4U0Gbq6oAtovunKqIM
G6ctiGZ/WOH96zgpddld7WTR1SKEK8KKW9WVamkOo2D4nxMJtBBZulyUtRpB
Ymb6vLt5C2iJtO8MLhh9FIfw/uU/ef59WFRtLnhvjo/1d0hJ9KQUFPKHN8LU
6qUl1NPjxC3v5ceo0EsGAl5Kg8n8YkiTJU+WUWigidQKxWzg11ZAcCvp9a5K
hEEy7ngQ5t2b4Ooqip8nDBpbQ4kPvYiENVuTXz2q/Lqm/1n1LyYZ/ykuppNG
AoCB6BkSIpDvDtXIazfBaecu7PpmxqK/D93U2ZT1fcd71dX322LwapaXOSLy
EGosewH/epsYZebIk9anBKzC0QLkHs6QENguhQv2o0fySYxkjMBwscSPS6y2
4Am0roOLUVUALBbXkp0n8e1vlnxtHrrJ88AhP/aeNVk3A/Y4lZu2Xlv1zy2v
Nx0gWuSlhvFcFfXHUV7nRhIZajF0WYsfLw2M5ye6WfF9aaz7LDeM74SNz0qu
GL+wMfjQEW8AXCphLc/RMlZx+Scu47urYU7+D23GOcMyHxdzYm5Z116r7Khe
vPgkxYhkHjJKDDws9i9ahGGrA4/gi4cUAnDP2Up8gO1GG26ecVpMpYgRiENf
fo6SlUbnkjDqDHp5BQC9lDKhxx6U66J6gJGHzkzFvi4/SC6rItTS/FaTnSu1
FaL17IuNtmfviTpYlIloRE3cjZU+4YDxCNEg/wwDjJQkcjFz4Z6p6Cd8/ftQ
qP4yIoPSn3CCHHDtogmuFVEajbFKirvQg6C6lc5g57ReIsNMr3GEgCL4P6L3
d5rtI3gOt8meJy9iP9rYiHADsjRTxZ/YfP6IzpLOKMMItSO+ZalFI44nUoU7
SdGnV3qVIw009dqsLH9qzHON9Pm8WcuC4oEvWxS/DzHdllN1ChqlB8EQ8CM2
njPuvpXlVBgLHjhpeMKWfyrmlMKDoCt5kXjrFdRBqABgz5TIkHH2BDQy65ba
66uuo1V4CTQGnZ4zO+gnlPeWYtk7z7SQ/tTwyReU3w96n6mh+7egYkJfTB9s
OOgavt8DkYYAzdQJ0oH+l9W4sx8YDVfPZ74xHjn32aOSkIxQmrDxRtp3Pn2Y
DEBisuua1uoKzYHAHCueQ+QRbO+G4lTEgt7SEpLOontYdNP7nBqwqpdA0N6r
4DLDklEmYFLdjkLLH6FU01RDuqgZosMGrElt/dLA9/qyRg22xD3U7GDKg0LI
AUvWLfmDXzXraFFFKCS4OUe83cImAEG4Eu7awhh8WBo4x+gEDd2w+FRqnwGb
DDk/8c37xDyNTtws96n9NxvZGsKzSnIpe46EtGV+jT49C0S2Aobd7jjf4QXs
OKRY31oLBJPDWjrxtqF9U9HEHqPQeYjwSyhVVBaXkY1Ygslfx3LQJGoWeZmX
aQkcuVBVMWFhZ1eoKVOwf/+H1Z/7PID0xeN1VpY0KWrFkfN2O3lK8kZNxGtT
XypKqt8UII/RAjZ9DtYl7GroSrCxgpCDgOEiiXePPFfyBOaZmMJ9L9AljDMj
caYJ74b6byFRbVUwLnl/XSrnzCAwhGtTP/7aeIeQCRrDOkLFge0DAvkTOgWa
J+g72D5CIqppUjykCZYZdtRGicmAU/srG57cmIL/R6ke142Wbdu4XjrRZ//y
+iFYikF0n0uq8cJSWfmEzL7tbZYi2fqlJtJGGJGAFu/NpuEJMVcW6qu2pL63
k7LqNf311dN8Ub8K419uqLsd+ZjMpBuFPKT/rvGtYfqkWs9kwYqOoFx7MPFX
nq+WMu3WCyfR39Stlctwy/cCuOd8LEsMyZEkCGgf7dQeHqe0OXvE4v9/CZ5f
K9C8b7C8LyRck5DaMVgB84/gXT+wf1nfqIIHBMl+T1dcsGar+9dPLKxBKoiM
CafhXCbaB6S9Yuaf8NgB97WhOQdNE/X3W04pKt4ICGckb1RzMwj1FWkzJs8+
iI1vpZyA1VV8LEv3j4+HcMVBgLcH42ow/zPy+nLCPgWSKxlTGM0vgQwO+kWt
4m+hmREiD4mEqesy4n2gwTJjGFCK72c9NvTqf+fFZxXKQLr+xoPxNOXeDc3T
DmVvVS7UDVSd5BQoXWwyQ2rs4j4+RA5RSYAyUWwEoG6rP5xWh8E8XCTj5tB2
9bPv0U8Lzpt3MsLsXnKKrv7B4V1NCtspaOAhgCV6bEZ0RtbNDiPv6wNPAdcs
OYfwhe5SvRX20oWCUJKD/C0xlYLJF2XTWl2Zra8ELXEIsFUdlRO3wKwLIYkH
Bp0FsD9HywLcnV+hqO6oSPKIdDNPJg40aZulvnPSqxHItWstiTtCCvGTqxHC
nn2LIFWvGiV7078153me96eJ69Q5rkUkhVMzHjjuYxanilmt6PP05Ra01IVi
N8Roxm3OBMmwHHI4dFJQiYwqiraJFI551HVYlhhsm0nZzxae3x0l7Ha6SpIg
aIOubwpBPcieYM3qPnzvq6829m8J51SC3wL38Prgqp4fi+JtGKsONyfg+rjh
DC0YklOk7mmJ7GbsMdIwc9oHqSTDzskWH+FyXdUVnZy5pL+6Ww+kPOkXaysk
1oSAJc9ur3e56QU54lNRHDmp9x1Eaa4bmtxr3YV7TQD5T/L+04I2mKcve+U9
xJ9a6fTWxVJK5z8fhP9PaC/d0wwoUtHSuJcmptwwnYihi/ttWTOPDPn/yXfH
H3Qkhiihf+4y13PL+9MniFy9JTGxhja6aNlJ7iELekvSEdHXX0vBTb4VzNVU
b4AcOh9xHrnO2DKzvCKdXohnSxUegJN8IAk//7pzdN9JzhO2Ene31A4PpI+n
xlD12Exexd+y/xdAIQWJXTjFdA8phrnLK0sjsnAX7ZmpLVdWD4dPtWj7FPJ/
WXt4T+ZU/WgHgPzRkI6tS1iGz0ZCZBxVp2W8PM5BhKsRf2M6Om48mh8p4gRa
BicKhdZLIwkUPbwuCVUYntHsZxOZTwcRBof+mxH7rgJBCExPXU3CbVZAAQxA
aD6NEDU6TqTR5wOySFG7+JXXUILRqO6skjlga1JK9Ii7DCtsRHtBpgcq+G0p
VGo68Aq2/4eSiKf2rW0AZ62dZktWQsKAi0om/YLf38Qj/6HepB0J+SCo4IbG
5RLFv0dfcWilAS7LBVZ/gQMEr2Uj3hzTjb9hqjjSCluom5EWNWr7/KawiFst
2RmCVu3sAwLtEWWF0L0dHJ2izCRR3Ya34aumMJcbJl7cMIQgfMloVkl4Wm5b
PtEEvZIu6Bqbw/q9a55i957rXBeMw3RWcVBm6eSIg4u+Lo88qizq6m19V03y
Xh4wmG3LoT9MnQuTOSyn81v+D+0ym+ytnCFqP3SVrLveHcidi7oGXFigusIO
9z7e/n36/mTn4aDUPMp/mkHiqkZEI53jAdI7bqSdJhQVuorI9ee0T8+AAVjb
uz+FrhvEvtZLiOVF8V6OYKS7Tz5sQs5AmQb/AfXOvKg8NRRoEPBexZREwvpI
BNjRd770PKBkbKaArIKl0t7N3Hmyg9jbCIgtbgxoPjwqfH3djB+3/aM/wz07
yZRSUwJ2OF3c1aj/38clD58WizUgeLsMYvc+UJAvO/0B7otxV5S/P6YAOGS9
z1zXSxOxJJiFJzrloZxw0hxWRkHgoJGdKeCSOAhvOpw+AnYzKmQaqEt82k+J
uo8q2uTLoBUwcPFVnmfXvUgtA5hN2qBFmWlCalMYvdK++OMTnPKhszLTLDTX
tP9X11WaU3LsoKLiciop7p2UOg87mQqxq0XqXueZZxUKitYV5LIu7OVcaCXo
/7jwkD0rB0s+XvfFNHCoUglx5mygZQLQn39Th1n/6bGVx4GEKtSsFQnY045p
o7rlH3NfeeaY3s2ZPV+6QivOdIf6vGFZjtQOhsdFQ2QlaXvyIJAos2g5r9hZ
U7lf4PvnSKBrqyc4clPIpvd5C/VzRcgTjtkYfWvZycuo4oyEcJ4/XwyQwMda
w6fWF7/ihy8FWGSNP/kzpZJyniajMEcxkVMngfgqZ2tn2KPTmNu3JgE5JPbQ
aSbe+dwmgzkpvvn+ZKNXqPZT66946408OKdlPxlh7waD03GnwXdi+57DSqr7
fmNfOEWhYaKqSkO7kax6jJv2ucCjGQTqey/O4X5WFQUzqiSUvw+kBqIAvTTb
4SQh2o+0qgwYznXuJKizRnRUqd4DY1kTola5yDb1JJMYaHF2zpSewPU5gOJQ
OOtNmzw9LhTgkkj9IcuX7R9oootP4h+/lbArB5znrwSHi0XxPOnFkk3cyUvP
+/6zizzn8jY+MOAn67TAKaqEC9cTUlKY3oXRNBQZHf2B6kpm6ENWxI9N5alp
8CXiCeeHdHsfZwYGERb5lrBEow4tXqNxSFGnbkCiT6LlTwzZFzVyb2gqa//D
3rFdIlkx2asuaRJCwXLEarlkQFLisDOKSoesr0feq4Vjb+OkldFU3lt0Bxn7
fVfrd1Sd8ZyPcrwPV7ejOD2/JMghVfC+le8UDOV6mvDsT/WGhbS9dX7P7RpS
62MFOkUeE9rn464x5MEFOcCIGCkqQhEDuk7jfWSRS/Qs6DB6kqWjK0RMZKbw
HxvPXXKPEONodRxPWV99U5A6qZtJ0EKUzUTdlE7sl4wjlwpMlardD6kE5CRs
8LckcWTljj8k7uaqJBi2Cel3CfEkQhjfKV1vYVXE7ecw6rUb+QOjntkAXiIW
WEGglqXBI6ynUi5NcbzY0v3gz/2DOD4Oem3S8QQC8piYsJGDyiSEhv/MkKOd
27cjHHhP0p7emzx0bKHpVgdoQ+jsXKuw/W9O8WyskjEBtEClwuFcb9Tw3Q0Y
X1kB/HXOYWPh6us04YUK0h/Q7XTZg4ptsKzW/xNBsoq3X76achUa64liD79W
cti2JYrU2fOlfy7ST+3OfYZD1vZhWabSewx0TUdSj4ydVE2s1AdsV+GIqOBR
ENBkvtQYUegr6aiYqNeFaBPyn97fM92boXidenJSNeYEkZmjuSKtXj6+CE+P
bPjqe+ddel4OsYaqGzZ8BsgZlwAx5CtRfzNeoNBuZHO/xm7RurGZ7lUwxk6B
mDS8or1yXGZ117S1MKdsxWAlOUcxKo1Ycn6xvniH1P36fUXzV0bCE3V4ujh4
h4FyJQDxGgAOueK/iAudfQ+qB6F9A6vLluJ/IZwdwRPi/6JeV1IVsXOQbA1m
0JYUp9VlyRPjTZImJ8gTLSZQT9/+aTq8duvFU0PuUVQGf4QMD6m4MOmiOTt3
7zrFb24TcnNFwhxWZV8FmNZr4E5/LKkW7oD1fE1jPKxiiGO4vNr9nhpfb9mC
h6NoPF4U5VsXmnh+Zq9ijxROwwah5VdfG+xQuUGBTy8dfcz2NheW1s2EXcLD
bzYjd0YIrK1Pm0awY6PWZTOoLbUh2ghyPT4/GCLTeHM+MjqOzgleeIXqmt8X
HIaq4t5RnV69y0QyuySrkxifs1FGnLWlR5S0WgYz7cMshSVsdIcYMdLXmso2
zOk9zBuOXtwvxjmoPZ3dvrRaUa2VPbdjsOsvqzq7vVwEmZYRraksYa94XG8j
6b3bbnZlLWe8zg3PgrvFwrsi8So+lphVdw/ciJlfBBvKjALrKy+2cn46GwV0
q+HoHb5O8vm7ClaumOHiVSTalIj0yxypUPnoc48IMQNI9il9piBqXrat3DMV
BcopMl1FyRLfbbhSIRSMSDixY63VBWEdobWsFtF4E8y25v9VMFrJ0eUHDcJb
21m0KDJfuoLMnsxhDle38SrY3RSrhsw2iLIjNfasEjtxTA5jYW9UVB76Yeu2
0Ql6dptWLcXe4Bl4vKctsr+4+Mo8o5ib/+ymuSc8j1nFW0j91u2P3e4Eommo
dYQ6TVn/9m0j37WKPJ5QRC2PClGgcJM6tEzxz3sPlnChiS2mm6Ov3RW0NB2o
8xpEWuYhKRBXb1FqpYW//EeovvJUkWJcTCqZUkepbanVi7ykvp8g/IIwrhmS
pDIV4DPkGmJSITg/cZZMirL2mfKDCm26GQZ7jNqyh2mcSp+xVMNKeBFZV+Y7
wcBktPw0Ie9+I8Q8hAhlKaBrOdp99qHPwvuLoxroU8yRFtI47BosGzOcOYlT
gHyp6HWPL6Fw9Z0UaHxYjOXBmqeo8I5ubq67dbIejy03nhQLYGLAHt7opmBA
ASadaIoBrlY9uyrZiCRPr8sJGHNuMrFTsk2NO/LpmKPmdnBHdDYup3NexoC/
747Qk5gwzC4YlmFPGHDRCCQ81kp795SCF5FAmXgceAoS0zSnHJZEncVZR5zR
S4VIz7nxVj2bwWZjolArAXceuvdTTI/HZAoQefRRsNplaRyjLqPwKqaRlVA4
NXkPyDPFX2wviHoVnkeIkT6trwcsdTxCB1nj6Iug9zJM6D+7Df5Yeag/XSR6
qi182Uq4b8KLdUy4fxAuHgOfshw66Qa5unumHHcLCC6j1Ar+zweRtT984ln7
DA08370+ETJRS4JJ21wlxVJEeH764xvP8Re7l8kM+gpelT+cqK3OTXcb1ycU
xnA/G0cON6OA4JDMNsmQ6Z+gPhF2779QabEjrenzH9XfvGpJ08Zt/sxepdav
6CHAjodmHwoUTLRtZUTq1W2KKuhabOmTr3w+CbKWreFeM5Dr6M6p/fxMXMz4
u2upyuj80riQG5bB3ggk3r0GGusWNIxf74RJ1SgfNsFGVjQsx4xGCrFAFwXq
3Xk3WIHcfwOeE5Wilzz7Tw6/jRUXydpqHTnN5Vp4ZZi4YFAZDf9zMza4QqAz
1+2uluvdc6gX7KO/3mmR2wDvpUMdC2KuOjhcYDN+Ni9tlwkxxqqgzYDfR7yj
3sQXI8BdcQtqbDpYIvc4Nf8DetHZxcm41CR5R3SDSsgHT6jJS8itX6FktZRz
rHAVZP66QoXe/y+c8Tq3aSvGyhsyWJaeaUD9r0r8xoKGexA1we6X92mLVmMo
0o0uCLVD9v7+o07WAZPJm62AM8dTBbjAnmEWBdufUQJjVM40lxLZIqxO87ay
nIrdyMJMl7ckqYOhpxoRQ7BAtuiw4yDYY28mqgvKMqrNzAbQ8dhXv0oScWAS
1OMkJ8AhcWuimSKscR/t3E8Gejoi1uH2ewWQoY5aNzKeeXhGYpHRA8LGt2T/
74P6WOycAPyoqMZGYXoNlTtFLgA/MylyaoPhTsVs5dMItd2UvDOt1oH/m9+r
phhFYo5/BW7kAEiSE6nslqwVbMcqEa4yfvFgkbDbUXlIMX/q2DHmDraFXcxS
pJmn9piBDOUJhXwpoX/3gGDDRGTwSBhPclhDj8vHzBZNYFlKxwf3cH1JmvTs
6JeYs1pceNcbKzW0dU0o94Gh/JGmcZulAiw8j22SN2jAR21q6VA5hri2TUct
UbjgJAixPtDdRFdu6WSONltdUjBrqWHTIn342NMi3jRZFcN6PwsKTpA9QJPH
cmXO4QfwLohY58NBtgJ1esrincQeL8alL9gRyWGfGO5Hn8FJQLuV8MBCBnq1
AhrR/5/hMyVT9S0QDCxsU7CEYyuVKHSemJxbIEhyCmP5tshTcsysMF+M+XYG
Zqt3+4w6Clk6KguikChnrkk20z+sibCaZ9ra12o2DchXjtleU2PKk5LNBrLP
sQiWGxK7feD826GwrLv0CN2J5dpzjLSv7ylNKwLm4p8ML1XrVgHbX9SePo1z
rRePQGQeIS+5CYhrcvUGLRQwoIhj3HhuhAjfXCYTab5YHbn6a3wiVsuguDHd
wMYI0moCheHZcmVQPeBlHFF5FKNhtWJPVp3Iy3DXwsdQzAGPrBVWq6UE2e4F
S+7XNeCNfn/NC0k55h9LFojIZLnIYTm6WdJm5D3b3mqTOD7OXJElwvySi2Ap
pndXhUtJa0FlHIc+hWApaejnTq0ldhgyucSN3WnH70BrrMknwJKE7Vlf5AUJ
SlTBakacHPPFSRGBrEjyy1FyuRwjzTOa3sdiVowNms0DDZkiDZW54+ZbrKQv
1+m21Rllt6xiNXVOcJ5Vgumup75GyCxYqzL8T6GdGMTbsJ94JSJIQW/+5V1P
XIUa+Msf8HXITWq3hUCXiY+bj7i+UtTfj0qTinTqYcjWFQMr8QexQpCbV2aS
1t2kEWwPbXzAm7MqJdb8cNiasU+jRNE0Nw3kP6fyOPsqRY2/QOLC7MfriMg0
+OOwtZ2ZpvHSalfK4QTK5RNO/0Bf36P/YSZpl9Pg59NwEu02iJvmbzb2zHax
y1TN/glpCOTQ05cS5p0DOVreX5NGkIM06ZbxaMWg8geicQfizX/ewvzZJiej
UFdjkcQ2qS2gZs9wzRG+d/hYJdRG1NF0Ju1c5tCv2jzE/5CnwrW6vdV4ds1S
ftj9qMAiO+f7lqAgucMeeVF1RqUUmQKtzU48NCGOegH5ZOpDggveGX9+XYua
i6Re28Ekdyw27cAHrSoAMF2eFgcljeAgqSbXYOJJB8dkUpMt3UmiJhMiJZfE
NaQy40bTHK4FImb3by1Hf9+y3Na24OL8GddSFu0ncyGmlSU6B+AgW11Eioxy
+rtxEpBzuYqGGpKZ1rhGG4RK9tiZOyzNEKx3qx5CsS8KyhoCtklkkBsnuJ03
fDY7fKXkBfPF9e6Q/ZFTgc65dO0h6BCCOEmS80omJhmS68sBZrY0889KDY5J
z0WqJqukPxvp0axzyJcDjSI89LU6j5DSDdpWntuqloLh500SbUjhoQ/qqSKu
7BjX+HNvDrv/J/oPy6aOU3tM3aZyXEeVkYhgyfkBrLoyL1qc3TgAf2ilUbIg
b1WkA4t4Jb2T5amxw76iIDIh7L/3vleuWeLHXhXZGnD42n4Lp+U6E2/sYgEK
h8ILSkCddE4MJLKwKSY9VnGQtzErzVj1/DPQBUbqwvwxNJ7LYyKKRy7Tgtfz
lTSlWqfeVn735zo0qRpo14h/kk1dMa5XHp8JP2Kmm+SGBRRJaKfPj/wA16LK
Rng+Ez96Jj81402c0QstnLB6qPXC1zA2YCjV/JduDoEy8DPZksSNPXcXWnJU
ve+vt2JyHzl+r1Ce0Zpjt8fvpq4tOxU3qOh47xaWAhRJvSzTGTtsTZsB6F+b
2NmMQkr86ToTgCiJSOY1GhYWdrtn3jRGXy8gQKxK8hcb7kxNWVvhtSRUKT7z
tRjGZ1I2PqMvpsl2IHnCGmPVGQ4SqnFGgxYyv24pM0Q/FJ0yoOhCyXWNRiUA
7zxP5IdF8GMTFUe218+Y2FZgyN5pRJmyBIGhNw7ph3oBO1T2NuYJNADLcDwx
rNTapxZ/uzfirStgruE31K+F8B4VxTqflOBym8DkfLRpgHFiZnBo+n3R4F43
JWEWDcHx8bR3VKtDn5W89mEIW1+BdVZsmynIVjQYgICaW74v0KBRB8e1ktlG
fpKbybGtZBlPKmDx4R8Cz49WIMVzdBeE+w9abk+8ApGnp1T46WHk47eWUMl8
dIdj0hg4Ioe6l02VOppSa0Q+vPxHjNbmfh7ga9/2cF7MuPDRRcEhA8J++vmx
lERz/UsJhvGR+45TspR4Eun7CJoBt4RDTHJxruwjt4aJJh+0HJt/InfHbkA2
VAJ6dndiWo0NgSuAFjXFqU+nwJBSymuoPWOayrUK6wpNReMKDx0lvOnAQvaK
7arFljv2M8eUh2jfn39gYqZI7+AnP8mT80lhK4kAjVAWFyuZB0mDdpwidcTk
qkUGmhXpVHRuirhI4eX/Lji5V/CaQR9Uig6cigLY8awTpAX7T+rUoKr3ErDx
pn6MQLgkXQAuV82kdXYgRchozbZ0vnNCzXVUg6GPSH5iJ68KKNygEZCEr5OF
IofW4v7+cPmKvNRb1/De5YiogqCDGDaw/rb05OSADNJqeC8fj93tx9FldtKW
S74c4RAR7Gnz0hNK+bLR0jzC6YdNisBewoJD7Bjz0J9VDcyGNF/AGDDBVlee
opha/t0d1RXcubd3e2byzeXtqzE8mktWMf0TKl3dvDn18dO3txUgQH07x5GI
cv4EpF2C4H2hcCYoGGLvdk1uNaVt0EworamNXZXwrSk4U+hmCSGHoilrrmCF
MuDIa0t98dE0MR/QlvIsdQhcEctB1wmUb0QAJXwqEk0F3Tcst2+HIUgDNtmT
LjphaVxaGuxD00B4rcunLA7LgP57R5Reu/b2XVPZqeFQAW/fmTu+ICETS1z1
gbDrvsuY2fPvhoU+jViktL3t1CPqStD8cMk2AgFE2ne9Hc2umTqvLdeKHAAD
GAk5fzqoIPhMmOjmQ0YW8dw6DIV3vtYrsnQM/5zWDX4DblHnOir2WLYukDiW
Z27Jm8Q6mgbI5rMAGeAarqC+w+6dX7Mw0Jce9K+SMxReErzhl+UmHtPr/0ws
/MSZGeHinrR7pvMjK1DVScCT91bSZeAvtmpY5oySF7S5605byQzBi/qUo4z/
ArHd8Ocyr/tn16Jz8PhVR91EAuVudopZ8irBJFjazVFXjeUpcEXUqj6ar0TC
8dPzpzSrpv70rtsZngHQT9tT3iDRfotqzi9Mnrc62UXmO0u9GVNXWKg2ncMt
m8lp/sJfHW8moOcy0egx/o5nulUpohL5MkByqBevUVd+zZ7EMAxTd+T7S9Ev
c1HgS1nyVO6531d3ENb+UoHGNKzP6ErOkiRv9GAxx7ekdb7U5SqpES59EcEp
WO3jVLjjOdhSfIkrc7WylDPMHCYTIX2UcVhzbEvAGKcmSpDpCs1e82BG1htT
XXV67Uk4QXjluybUF3FvfX/0nTnBZqWz7jCcvJ73MayRSM8TOE4HzoEp6quR
qyOh3tjcjPHF50rjjsYu6UgV5i1pfLGvLwvIhYM5M06Q+Yxj7smdtmAvZmsN
x+DqHZlKHVYnwKAvJ9J12Rv9eB+xfUty27MbhXdJLGsS/nH2twQAx0EeKUiV
8dh3C7zeKO3DLBZSZFhcpKIXg/BnMdvDkpJWFXrt4nvwtEliBxKg1GCMY3NE
zfNjZrKjWEczYN48Lz80MwoBioewbb+reztLLgORWBfaYbuzTQAjVMnhX58g
39t6IlIDSgIW8g19Y16ThXFxsUYA83U3U5glJZNFx+MwqS2NTS/YojiqRtZ3
i4LrwljTf1aywPnFqGt+T1s/U6Cuv6eYF5jgQyXDRAI4U00shaDZbAqeagUU
oYJveDkslwroY+r5JhVNUyVwXomzr8+oBTpAQNTQiYKqJyiTnAbj65GyVnPM
xNcar482tgN7x2Lvdqveu+K1r9/WB2GfPZu+fla3bQ2WKG2rgyvV0fATknMg
nygdlklbVqC6M4NbcvQluVT2Sa9YaYXYmLk4bVbE4+q/9tQ/3ZfuIuFYM+o7
l0+n486mTPmHLYpDi2wsUKF61KNAhhavYGw04j5TKCAGz3AJu6RjAxp4nlK0
bWoc3h+p5lBNCrFk4qh61Hpu8gTjVBh4DMgeDraWqSlp8RTC+zJOUxY4rKkj
o+qPy1Q/6EEDiHdK3CxQl3uXZ7BEdjZ4oVk/+qvR0ZKEztthPhDl9AFMY/H3
R/BkU6STppBha9yOx6BteyEN9uZzXs0l9I+vFU4nD9wva9pPzeTJzevKKKEj
PikIP1OgsqAEr2q25jXpguY8XNIDswEXZaF/gMXSU2veumejfWdXFQQULxdS
cOrhaqLB6v+rF0QeLgFR3A3VhhlVdOOlB3nPi4caCZcGGpcs1WrmbAc3T0/r
CsPgwdj/NEeBb4vPHFxpEWXKeWqDXjNTmpILG+lbJg9K1PoNmX0nSNsIRd9K
sQip8GA5xo0bH+lQ7bzXPoG38SamqE1pFgAGvyu/Ount01RKq9EO1RwD7kvS
QJLD2BRot4ReBSvxJPIQ7EZmu7+hKIt3WSCLM9wzW6dfTVD5vXffewwfsDyf
AURBKqSMN+zBmdDvIHA4EW3q3lTOnbttwVPvsw9i+FR2TV1iMRESimR2GxRg
spM1GIw8dI6ERHmIO/iuShnRiLWekM7OuonmNo1C8YTDncxpfwR5CSggW4ly
OpnEUjeucuPyIwpJLGh3WEriJqSed2QeJQ6acIjwktLa6k+masCNBQaEDcMR
9sEefnLSt7nTiXpdvQl5YIDKjPMolSqX1McgC1okUd3RLi6jwD84O5cvcpyH
Z6UNabIRWGkPxVCxY1AYMjF3Lr2a6ZWm54pe2joH+FtIEBAne4/hHFhCKCfV
aN5kXvKgYfxbpAJMcstaBXwzzAgsFUfbuHQBsHklp6/wFFKORbyU8VEyfEPl
SVhZ0AATnIEdHhVeUJZw4kfKDS70y1p7cfEKp9mMUYU9ZztQ5CNE0xVajVlI
IWIQUjmmU7D4l/JICUDJZ44mhMn3VCMLTg53xfxne0PPx9G/ztlCF9q41jG/
Z2kH5bxrlehpkfXhsys3/cu5CeXE9OCbOKSVFSgo3QAdrvr32fTkS+Z1P9CV
8lp/qB7ISoCqbpMA573lwPGpMZF7d/o3N0FxYgXGnj+GNms+ZnXCeubPaVPQ
dv2XEPc47avb31xfN82SIjN5w1hWGyMnirvOKgbFPKK0MQwGlQ8O39DwK/1H
KKniYUJCa9J5ljKwIBvmeppT593RTUctymKMO5V9IE1iOgHV55tw1m8O8Gou
DW8eIrgT/SvA7nXGh4EwPGbsvPYblhy6CpWPyLXbcu7jF78Be6YuqTLKdfh6
mt8BQ69CCPCOCcZXztWBKliPWJQrs6a3d7BiGT23px/dJlgGTfjrhFS/qVuo
YGUbs6ZqnWcfkKRlCwTZNNiDkYHPt667xQHTkEaNKfAOs++/hva1E/+e7R+i
CPvIDccwRkpXQGwLxk7hxP+hKW9tgqJ82/7z+zPMTDATtfH/720bGdnRoaCI
yD15h1a/0mAAGDQU+8SLdlc9JfhNIc4UfRP3iMwwCNF10ElWPQ4IXRE4z1rO
s+iBJIiPXE+UVzAlwNLltzWGE1A639v0MMQEAXM+tl0p2fzkqxja5XZrk26b
cN8sTo0HqbQuMDEgZy0b29ftqxkigb1q7OcaXJIkmjoM592gSVsJVwq8icas
hMEVq56KHYhxrsQ6kyzGcJwM/u3kgK/ILFsS3XtyqbQyGMhqZNwmxw2hh3fT
FoxDRb+GbccmuTqJcLoZZGFAhdIp1nIw3ZG2fXIonWHXJnesa4z9nuD58Opi
t6eejGv+uJuttXJ1aNTxWKEO2debwRT9kC6+LpeQCGt1+kGJU0w/4QZR1lp3
0LkfIee69I+3GWea2thaCv7B89lOjsq7bqcrry0v812BjodvzScoftzFPP3p
UrYug8m+TzUiSBZNtN5l6zGaL/Hbv98mag1Dr1owEECG/H3OplbqszkMOb63
7tMgoRX3TYpZbIcwBWLegCC7t8ncLhwfBM/HpYxlP6giaGIs59W49WvSMZ8B
ccNU9YezEnbu+oV8xtnsP61jI8FTIyaVklGXQAkoxa4wDqoLTx+PVi754xAd
nezMRXMguEZgG3G/uEytIwz6Ew1Pa1XGZpJCclYiyTuD43jcLJY7kenftOXb
njjsd1hVNu3/zkuQ0Ql7q7fzfskwxaICYAD70pAfGNSls2mfeHi2vY18w888
uPhNIB2soiN4M+kO5dsQlZaBZ+vbfJ2tsYxfAE+mQ5iQ18S3CHi9sUf4gfTU
4cxaHugSk1yfQWWVgA1I30mghnh5y8bHNTS69+ZeARlyN5pDct7NwE9hi37M
9trXnH2TMOEPEfHMZq82L6xC+WfXI48Ic/C1hPqt6mqJ5JJaTsPzKydCNMiz
BdP91i94x8DY+k5ra/WeaxD1zomEVjQLGuljXs1cGYqVF614lj/9Q4bobzJB
DhnKyZWTVnL1fgGsPU2BEZKRyBo1kfGbQTNMk49HCjDGZ3jyPnXIieKjDLdU
NdG0g3WbeK8q6QmVYOaMNZwzGRWyUIAIJsWmAjd8C2CBXlnqMm1wk8lk7NZp
Hy/KfQqXI7Xkf+BAeOllfcJ+gm/jaer6nGu89UDIzP7ssOcKwKMLXBJG5UUZ
zRH9owza+jxA5rrEQxG596TGoUh1TBbL1OgXxdOxn5B3G2NRhEctzg0NuWdy
lSSCEnk56xuVxIrQtAFz9Xu7+RD1i0cyVKG2JjJzv3oZ2AkQQLZnu71QtZtS
MxcoTDsxreYVYsElIKDzxa6UMjsMuLrpse5E0HwXprDsqrggXMItHPRJQNJr
2fjO17lIaoCTuBACRm1gbGFgKyO/cga58GXqA7f3NuNUzQAXxwoX3Usi8GXS
G+1qd04OE1nNOX6ZyPAiUmtPytwKWjvpn5rFS2tRhTLYUhCRiyXmUHZeuhbD
VUvnLCcxdbsLkso+y9nTN2DvcZ+rUmmz18bXRSMtF/BDa471IX1imMyy4eX2
qWsTWdVSp9WtjIyLkxeWLXZNLDiV8BR1filI/qPiX6P+yei25B0nUbHTueCq
/nLIVTLjpLg7gLver1MhcmM7VXrXg1s6Yb2zmAnoY89VImgHbtUXZTuSO0CL
a2vBlXyB7UzJo1D5zpQupaKgDpYECI9SdLIZbXIegqej6eDHPsKXBY8bOHgT
FSyDOOgVM440KUXsxVEOZzI7XF7nc/Nq7clcP0Xr9VVWFTQauIxEVLvfocBD
Hnb5f/8HkvYasseB8KqEH/aEN5yJvbLGl3tSJFKJGnLuKpO03rZrwOHXtJor
RSG0TbycT6D34HLXEBLdfYp79LCquOL93J8EuJ4bJFl7S1XfQkevQygbJZ87
WoCvk2KyZbuhzmE+tox/MGGciEwtxd5SAadKJyLv5QL8OT1ey30UN3AyUTmC
YA+MpeZomDqYwzB5Oqrcnbv0hUGoA2MUSNre8k0ZRbi/k3AuAc8HgKTnbonO
E4T0lxXTYu61UPoQr6VTkFsCFDL38GdrTVGUKnsfxqIFVcucPYVvGYB8fN6l
hY4c9w6ikmB3Q2uKXrwuz2zUW+ytsEE/6ICs62VcFbAsZ9cygrGHLEs/mQlV
ZcpXbKdFJa6g3gPLaAUCepsMVg+Cr7zv1GZQhFh3ULy13V22166HTIbBC2uR
+hYl9Jzc+4H1j4P5DdZmb+7hUlgxmni4PYZXHeH9/lbw6P0CluzvFRZIVAVi
Y87SXizqyx9AB3SkbkhPjRNClLQY9gWF5YNhrc9En5c+LRb4xlxRXkoHn5wQ
A/iWbXV/HBcO/qxlQOmqXGIbvZkTCrLUpMjL9GEBWdjM7IK7mydh90MfR77/
r/LtH27lySht5icAmkEyYIeRvkv0rBNiQIDHhZRjn5dL4+p/u3GFX0VVtYLL
o9BrrrZDCrqsr2f5fW5vPjGAFWWUyJu7IIrNTNgzlFuXxbCR8qAGA/VUO6+E
IesC7tp+IBSH8SwKm5fryaQqrFY5dB7AAKnSY1f/YFhhpdW1of7UpSW7uCoV
iJUJEJJxhCznlR1+t++ifrG3eFYzJ5CZ9/u0Z2QZmFKbOw87fw3LgyjzgFfZ
VZIlSAyhnkGkGBf9gh7621tC7dlB9byo711YoHu+79r0mrNsmvYV7dAzIXrS
dhTt0WjYkedIfrH14w8vF6Jk5UGZDz1iO3NKkB2U1FTIEQEAS7zAl9TmEIY7
lbnme4NIGruilwnrdfPwCaNcOEEBxBOLStXVbhbPv7JTr9BdYODMmfg/zYbV
FdUaZNNhNV9djQWRUISqBCzAqjv1Ouaoj89vPIJriskWD+yZNGc2PZhR33sZ
kzSEduAzwFxV8Sqp7VqkkIUJRsxdIrZhiqJqcOS6ewch6XY4z09SS0kliaVB
osimioEfrBJTLXrXQ+EnzxV3643Pk5jWGCe4GfaoiJkQsN6es58T0ydcur5t
xJUpx/SYTrZu5a3RlhngJo8UuoPqJU5KcuYRWQIbJ5Ift3FESugmWK8GcaK+
wMM/U2UiIBWKcHKZxy17eqQWXoKc5s7k//bFhYKvTFCOZvc8rxZhMusuhHJU
G5yThLYg9euNHy1LN+KplcvnigWyo+/XxQxtt0WM8AdkmBnWu906UzX/FbFm
B6WEUUHEkbTqVTQ4Jx9tQ6r88VZ/jVbbRlvEVdriuxjpx0hZiWwSxlOZiLfZ
NogjEzapTj23Dj95bf79MLb8jdHtiV3etfcVmMYspTqSsSktaOh6XQgTR00L
tHViaNWkzdFXg20FRpilSdMvfcu628oMvr1O5cYqEX2YU2aZvTVsSbryIxQB
aWSo9boInEoIjjhd86DRapqALmaynA1QvyB0X8GtNWa8Fy5UnkhP+bJ0WCYR
/mS9BF0Xw6fVK9hdOH6zvY5dZV7fJKpc53FnKOOgapIfj7JYmqywNQeuqV84
2jB9uFuXxChB1juawC+BSDDbOkeJjdGDJ54nFDeR2SzCp+3GfAdB1ImefqTK
PVbimLYYxJsRviqt/IypiH4rELX79tTawrX4aV57MholED8aOexoko77SrdU
J92VLKMyFHdEk5Kll2FltnS44GMFo58J7RnWjrlL5J2PD4cU8wBec0Ymete+
VI9qwpgweYqVDsHcT8ZnyaLjggF7oCb5qPhZtVa4hB21c9942hwupVMgb70r
ujmbkO0oWrUyXO2+wWk3ggFZyFVYlIuwaQQnKp7uu++Rf34i9McGsTHrKfoB
VonHs48r6CfGuC2ZjhPK2sr0LxLjjhP5wCrfdi8Nxhe/zGzFcMW4Po9OO/HP
c/TunLE8L+/jj5W7+9bvZlqN1d/ruWK978IaGGaktBMoGE85W3KaqMZbfUBo
ME/32OuVFh0K8GpXbbx6mgT9wQTIpVs4cKw70AnyqmlG+GmF3NhPseJeL9qp
pfkDxe6DtMGwpWpRF7/O4xp/R7Wmr1iNGXXmK6Kvr/NvR6abuDmSSyl7SmOy
ofB+bsRnpyFbEYggzl/LDAc28pjnPazmgM3QTRaI1UOne8YFlViq3acroO78
Pl++y3eHOVNKMZam3Iywwex10Tf6lEimVGpzpRIRKR2CbXdlh8646b+HVqYt
39LeD61DaKqLCmF/+xCQ0NxvcjyBGm51StfVQMSlJ2bEGc8zuYoHNchxpZyf
27+7ChbEIDZ01NEqzwRfonz8vrO1oEn01HvksaBtSG4caeLnHcwyMeV5/uoG
szPgNU6ESNtHWvROQ7AZQm7wzapavTpyc/4tQE6BPlMxxcMnTpj/KXM2HBcV
bT8WnUZsa/vd0Ykyn6tALhD1xakXzrztr32PBgY5ZRN10Lmgy2mesk4b+lQ3
pdzlWzceSJVD+w5KTxjUsja2ABoxzXeuR6MnfQcYd8w18BBfyZZHqn0aMQX/
VQSrv3oRaeY3dc0sEb40HkQQUiztH9mUHtBcg3N7wcdVs3SEgACi6XJa0qGo
2z2acfVwUP0ZBelYBaOuS9x8jtO7r0014HX3nhCylTZrF1TuUsnf79SMrAz4
C40XiQxy/pPK+Yzjbr85idO3L1yCRwsp3zKx1IT6wY4J27TW5CLFO1/mowui
agEhsYzCCZMAPCf0t8xgXbMyIdqgIv+w0VUZuf9Ow/GqZCoYtv85uZcEWkwm
y1gk3urgmEz5iQjWJ1oHeC9YZpVzkwNWXtQlE9HlXYuNcno832FKzcu3jNsz
nRj7IPUgNi9GOHlyxX7wOEPuJpVZDywCFn2fcnKCzYq/3enkyc49ChTX/nZB
rlFBukaxClwYBAEm39BZppw43PQdyD1fOXDRIUXTDzWucmjDIZZoqOl5ISWl
wmcXaLAYmWZ0r71XSmId705yj/I08kuM+Mh8ugoBx1Kino7RbkKJFTKPLCB2
FYkkkbHNDUQSdLSk/zBj16xR75rwybxGEdTDZu/ypvoIKXlc0OngkkDuHln8
nolgbppkZjuCXYpOkzph5Kmlqnp2cQb4IVB4vUQ2WqBRRlNiJMdacdIh+Yx4
UZiQnUpyiISVUS2U4x+axAxIi/uRBlCFClooIREwasDQtVdJKQO5gLucJIjx
G/W1vaJI+Y6B1IAbzlTg4ZpljkCZHtHfZf5+4Wi+DyW+/fkybm+jZhCkg8Q/
PZSTtchDORjWImJv3lIMSZ1YcZh/lsegqBGMvt9B7tl6THqwLjHmrwreigE5
nJj/xySKhGrGnO6zHyfkt8cngVHIjdVyUAzenmpglGYOKzEcpk06USxjy90R
Q/tnwSCQPSEWq40Vv6htZKLPPhU0UOuAh5KNBd8Fibzs/2ABrDsTeeaz8bmX
5r+TQhCZYehWsEo7ZbUyEEGQhl5aRLddAyDRWikjC0kNKkjyJR1G4sSJEZO7
Y6oNFmFdcRJXQVFAPl4sAu0WIjP3mJpZhaPcRlhqMpGWWEc92W1MNtM0uBm8
61F8QBnOvpfkyzDTp75Gf+4EjVlbYg0BsKWFKpECxAi2NijTsTUkOs/3drau
ZGY22Rrd03efRU1HtWTQdv0J9Z0Qz5DbcpLwj94bAe15S5Wf27oDDgeM/OAI
Fdb7iM400XJurcHFaHBhjaohM8NP5vkK/gLPCO5eI1FqPD/+omUyUR1P3i5W
9dipzkNMJk2wN2joRxDkh7lpZhZWXhq7oKAcLZ6z/YvMbVKEb42gWuAa6hkZ
jt3mQtBAtPvIiVn6O/WFCAONDweylozQEzBUnncYTN5Gy8A3ykEn5g8T5nfP
Z//4AD8obqUkkycVJjADjE/0e1N9hVdI0wRrPlEGjwizzIEV4wNcGO/6uKPW
O38yWkG6Tb2QkTjoFzUTbGHVBXY/dK57Ad7qN2aJqVjL1xBPC2oC1I/4cAu3
we8KibUS1QqoQ5nPICyW0w16/UNl9V+hfGOGu736p2d8+ZQcRKtb2KhSXO3W
KIA3gfxVrtsOr2MYNhIIUakoUc7UFyIdKMqwAfIOETQHG62tUKWV0+pFVKdt
pbZ6kR1PUYQuRLEtjf0kW2+EG3Lfeyn4Dg2yPA3/c8/3bJHBmkKHAHWoZwb7
LYKXbuTGXT0P7fFfkc4ltZBlhXC+Q+Rok8VShFl1wJHgFI/qR9k7oLDs6FKy
8AU1JS8T0Q9oTm6a7lZ02feOxMXJe1uCwGuJFtm9IuwHTgSVXZ5sQRWRkWzL
+99jmtf3EfVDrsxotXqkTyREXwsJWRpGSDzxRETog+3Ixf8rXGg9LMra+vGN
KFb4i7Qj2szkwIH/Dmjb/nmnDgNXcpkcZqilpdIiitU2vlnfP/exXpK1m/xV
NhjcmeNPHxHr8kA4m6qbDs5Lp7EtjRCxZEXq/IF9z+elcRRxLbqI+0B6Wik1
vVxmZ7s14pSd8+DSquaV5Pzkp+r5i3sxIgWVzJL7hh0JbO7PkQDhtMHxxzHF
idl4viVO0gmpS40CIlYbVpkZLJEqar4PeXN+UDbV7mfDr2jJc7LYYas2jYH5
hyu+JHRp055HRqruAr/ZICQ2DtCZyRKXoEbfQ3Ipe6trj6v4CJdfcJkf6fEp
g6vTkyITbx9pYfUU4eXUgRh+hQ/nF4Y4pDKli6dKdng87GhNXUVCwf5BYPkd
dMS33sJKrIk6yotMvT3F6+FORVF9Hl7p/cvyKlcBLiRnewGLjifBaWFoPD+P
mZxw1ISox2ukM1VemyT8/Usz4V5j+NGKK45sccoY5UVTUexCwqPuarm7RHpM
Fk2haoTbBy0p3y4+Bx3IpyjMfzhs716FuQJcyutlfg0OwDN+Ronaho5OsUvn
2oiFxEVlAn8ds/bp3YmlwXwtXN/HxMz/xYT0cFZkZ+W2F6WXN5nLgO6OwHL+
7zjGefwrWYgqEiubfuzC9EkLyJEFkg5QhqzaXvWwii7MK+oNvQdzypdq176U
nG1z6Z5Ph0Mf40GgzQEfD5Imbjls5ZllgPSwIj/xNDkQZSvgWjyjEGp4VDVz
wV+FgR0gPbjhAXZVa9486R2cHnRVbt7In3SDIn+KQc2jOH9aav57n5uCBRb7
Y85dtKtybsDIu7dSBmc+4bLuizizSMro1yb9WMl+dntJkvf0bkVuo985ljjm
Z+ElRg6QvzJPrxr8Z3lNvT5/hkQMfsIF8dR+p8WhwfPqo57yWp8Xzi8QPeSU
Rgo5vRUwMQEQGHh+uVU5OlF6Vp2oV7WuvkSctxX2aR1LbcMggyvIgb1W5oZL
N/DLIi7tivv8KS1wC7F361+FSiRaDIreuVBVvYD3mBeOWbMajQy2IeapXmKi
/lZn4J39/EHGRrKBId15OQIna7ZqwdhEBUiOwjzn4EF+HP3UaHu4+uLj13ga
jAu2r5hKyKc3Ft05RrsaWRJ6hexqpwbovrgBGzexvvO8ZGe9VIZc7DNRl+FY
WGmdtPFyWxOiGsf4GOMNSa9q3Ix15DfyYfga3RlPU0/4dkaXX1UuamklhDzR
ySYl3AYVCuE5MArAN81io4oUai70UdFwNdbgn2oDLVP9cdxI5SW1gbjKl3Vv
UOdVAwdTr2+bYumtQdvjEvN3f3yOSEbLjtPLy9Q/PUdyQU7E8sZavoH+t+wK
ahHu+n/bpdDhmU8lagTzcjieT+9ZnaTY24sNGQtbxcMpVejvYimQnmj2ueSy
eoK3KHYR2OwrqdFkWk7bSG6t0Sk16+Jx4mkYzsnorp6Q3S4zc0eFAmdPFfBt
kftuHX79C3qKW4s/OuutHHAlmHtw14viNLhiy9809FHxZ+rThI3cJBBfva6Q
N8U8UUYGWDFsG3UvPc85yrQHoASSihGZhYz9NJPzHt1fAC2dlvHvek6NREmm
v+e7Sh80XD/7i4FukpHQFoIvd1FSXPGs2eSY64rNBg5TmBFGbWwU77sQHdPX
dtKaZYxrPz/7ZF8zMCBIKVlWedkdHj6BaV9PVD8YkKD7fC4V0NnVfmkS+v/O
htQq4uIbTR0Gg6oOUFRslFK1OeD82l99oy2N+Z93pDqBYUQx5TZ7mFnM7tmD
pGZ8C4268pvQLIPjNenCtP2kmpMsYC1I5HwxVznDlDtwnTcMRvl57wzuEsjT
JblgQ8r+b4cZ5VsyTYhCHFWGH5EcBISm+ZJmPWGOE+GAMelbre5HeZLkE5jy
PiBT4Ejgw0KSY+diNOHZYIUIiKKCjJjNNoUGgNsp8DzA/zPAjYHA/c02RFO8
mFoELHNTB15V6wKW/ljO/slt+d2B6UFxxqSP/+51us3TG4nGft744bzudraq
wrXmkGYlguwIYuG9AY7icPrKvZTtdAgHYEAN7uLDiJ7U/3bB/WHgPeqDPIyk
loxniFMHqFUk3WhS81B6aJFQ9y5+gQHcr9/gYO7lMzHMcd+HrcoOKNNzCwCW
vqWW4VaxSiXcwoEL44KQWTY+yzBu8DOmOO6ijM0rRTZZeeI6PhGqELl5sbva
7FOhJSfFjQUeufl3d/5ywMRCnFMVpMTZt5Bl0bKwcVvD79TYMc6CRSNSEOb/
9khWlad+HwDz1JpIse4Kpvdb9/c5cGB8h9T+V+oGHPY90ETJu1AOf1kHzxxz
/zVWqnQgcZZqbE+YnZbnbhBucjp/2XyHcd1i4DKSkSmzJrbd+ydGpPZvUCxO
p1saSlTJbeLku691lQLAiutkkFU5G0+TfcgXf0gITaY1G2ec9fkWndsbdU9/
sTKkhn/39sJ/lc8+TYSUYPbU6FrE5+722zjsWtO8aiaFCFQ7Tm4TXPeqh8KI
7KMjsM0xZlxzFsDS4N2Q1aT7Rck6zTBWEwmQrpEQAxPrS/Rz3rcJm4pARubB
qmSm5kRmLE5+2ZPsi5og5AitVQkhtlTlHEcqzf8FUG3Jgv3Y2gbocuyyL2sg
u4wmS/rn7r0sIE0VcI0HPaPP/6hYanLw+IbLBvgpFGBS/2y/8FLEidC9eqng
YwkOTd1JIosk6/tyId+xOI0SfBpCz48jnMVu9hLJbiz0f7mm3Faw/3q8r7cc
NGgDWwcYnfukyo5gRo0eP9qrF4BvD5geC+9KSU2SOsU8M6umh4VLD1qcSfp5
JpLYT44L/04ircH1Q2+oW16fpsoNj1F12EHEIEeFtp1x1hT13gHECl8MdntK
gkrBPijIryyZci+kyEmKgj+Fg9AJCNyVreJtsUhjWVmCfioBe7TAZ2C4GBo9
S5SWrb5wjQe4KE2+lqdqWNQ9f87ZEixc2XOyeZ2QIIpk41V1L8hjZ7gWOwhL
Ywt9GyvCH0FjLWTMVV7X4PJEFYZVZNKeNNiYnhIIG1LoaspwftjlzmFqYhqL
G0m/+zj6q3/8PiRQ+OaQwXDBq3xMsu6696igGdgfG1R4r5+JRZkJpkOGfD8+
qBqKmOOh+jIcx0GprRSpTSniGBHVPPZoI/E12+KFlFvv2kxLX4G5VJwiQjaL
KzfYgnmM2l4atTCzfqFSttLNB+dvkdhwIno6/ORXEWrO60CgOiO35l0yxPW9
20dRVtDbSMiYFacNR3/FD1BTvBNsN4MZ7N53xbXHHnMxm2trxTE7bpv72Q5l
X4UrctLh5dmZ8eXGd06mtr1jj5tIfc2OrGnA8YstD01oBx569nj6ZrQfcwxL
f2+iqdPmVW9vfx6r20C4mDjMv7iAXjxCKYK67A2b6VJsaGtQj72DL0cbfr1r
ZMI/G4sWkhjO1FaDUUA7bNtKtljT2IZuc8UCSsanhpJ4fFXhZEBF+xu7vZkU
5d4NfcAGuyPLeDy/sgBg0VmnWCklrp2SKNLKf0F+Tfe6iuFhFdq4A001xLcC
g5eeNpMHLbXp19mE+h6u3M7OEWtZIsq0RLnYVMi6jWoBQBiA3LraDuziZ6P6
KCE5jC/vc9yWz7cu2aVJFhvv7OJAvWUcPdUvBqyQXxiMeN56N6Gwlt0qRNRt
6T7ig9Sj8wFhfa2yPiCRcYvbJ+yaSrDn68CnYqjJUyNDmpngFosvyEfUnLuC
rhBVVyAb0wd2Ud+OrLNBE8XAqQZ5lSRLUr0yipexu42ygduhQiacC0gmrYsG
mv9KeCTNCVpAyMy21UkaqvKvrl+NpC35dkIZGsFUqFL7kD/17Ye8rPhaqh+J
pqqWnvMnEXFrfhDUejWhqCGrmoNKpf1Efe9UX7lVoEYOICWtZgZUy4MIvGvA
pfMuP4elyMFL2CewsJJk7wfeD2ccrCD5S7HWjD3NTeIYiKOAC4kZaGoMyXp1
DTBoAN3xW6hec3bDLrMmdFeL8CY0Du0dFTwpEQPRQVjbizdHJpj6XxY58Zwn
YA4LVduHHSkpSsozjTKGGPEh+txzBGU8kEFS8KfH/3B1P+M3yAvAjPv36q0U
amF7cSpm7LSj86Ys6KjHiWsvEBp1XanmgjUaD7yTg79g4K7BIjxjTQCv1ch7
6Mkcbjgi4EmKhMkyWa+KR2GATunjmmcCv7QgC4b8P1n/ypRP8b6My0cPBK9s
R/Ygpq+EKyDAObViparNinXwanLqJgnb2kMHlyk94lJNzImZvpv3nvDMbRsg
OZhx8DjTrmnWFl9TYQfkG/bJ9INVLExRFmo/fAKtDVLIsJYZBTCROep6rbYZ
OQ9ZNJhcorEoNWs5jMLJ4sNbtaV6Re9deG+XnXBBrlSplwcpnhjdEGD/nCDU
22g+3PzQI5lv4zE6gOH5HgZiZmQs79uprkWihAdRJDqPDd93O5dhTS4bkGqO
p2qfaG+xRppPRT7fi4KYUgEmZrx9PI3bqEEndCfiotVlDndfT/2ErT6TzUZZ
DHGnd217zaQoZfcwDlZzMZ9fN+WLOopNt7mw4dffKR6myEQ4SJCaf+dGMX+l
Qsoy53O2Lu90MD0Tgrrrb1JrQVH/fZVUW6doOEhz+cAhqxbfNtuSGFYV7vwY
SKspFt10Y04A0SqLiiCb7lUrgY66f7uLLaOEuVNUG4U2/Z86JFKMbu1Btx6B
jdHND0u2l3eksK1jmCh7Dfh7RLxZuqT+i0sNQYwsliZutlvvfe5QiKV27MgE
nNjVlZNvraqWYdShc4kjmVNhYFjHrL846b4CZhQvLQXo2IYFrLEt4YDvhBaV
YVEnFqOPdOhB94uQPc/p5CG2yUPu3f6j2n3258jyaRnzvIxlDiIdybhJrQe8
ZcO1qrDH4kz5EHezJFDL7KuEUZnPnqKl1WVzTeloaUK0VCpmvcANDrcwfmor
HMBtwTcPBTIrH+pf0Bzhg/4FFE4I+/tzT181ttYLE7VOlN1ZOihT7SUFLomq
/s6g8ggkSrupGgw5xVrEW9fTkM21+j6uUmnIvcxaOE9ojJ9TZw3zrTbSvQrZ
mt1KhONCsPmzNytHUTZtvFlL8EgBcqSWmxEDwqHYiYK6GDaOvdYj+BolyIIS
KzBBtWfKdR9aMAP5f3Or0Q1ih2TASTLj9RvvmwNHPgegRrsukNJCvVvTsrfc
HDrKBltIeFlgvf5RT7vRwKR0U0MMzqFHW454WLRnnezEZUMLjf84KnW6hwDJ
jGgdZ5Eh1qFudJYG6mLbwWlQ

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqekSgxxtcy08SoGOZS8JyWAHpAXPa/mTYVFAvt04WRPlZqsdGkQVbHJAIeLM0OVO7IzZApH7y3WRS22/dqFrVPWvZ4arm42+ZsDiBICFPmwOPPUaM0ZuRqTISP03l/T5XSZvDllrauUsWk0RWfzimYq25W2WP9MpHB+yTirSlZuXrXyvuEXDgDn4hh3nmEUxANjZxcoXSaZs8UIuoLdQTaQAQpTaPyBvpAxB6xrymVT2SRJj9VCg+Oc5+o8j7sjVp8kDaMTSDCqr27x+feFhY6SgMlOJxDC7FeLmd/W6tG7f+URkLkjR31uJtMoIl8RHhgtETnDiFOo/n5cT8z3+CB+be3H6vjdHxQieK4D79Xl7AK3rYHXtmUXPv3gndarfqybMyxtKmXiThQ1JffgPK7PSXUugux7yJN3EPMtyg/SUilLL4azuDWEgGaB5IyGuWUp648JLcX+V3/NrxzJ6fUF7wGm/Cm0iZsjbJYprwcalFwC/90vi4IpW3p/7rVA14lJayUHba+zVRUPr/9WvR8XoRp5V6kpz8ms+lr65W8qdS4E3lqP8nP7qoX8oHBn+Fj+Ic9TnPpUMd4T/m84hkMd5zwwMOm11ketPbXztThRZkiL2+FQuZwILKXdNQ6vakNEb2fk+0qhjRNYOjvDakxEPetA8v91K5E0+wAN4pVddbxrbAcvIkCelO6QHtETfOJ+IodRbAjs8HgC/bKyoFMto15MGAAVygN4NkZAG8zdMBvPvUoHgesoJxFOMwHECwMzZegH5slTvXiQbIIuf7WY"
`endif