// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rCeywPowA/fmvfBtH9CyP1EFjYqUyrTIQlwgc5Gkt4h0Q/HqVDtBSdlX7Gim
iUlJ7vgDYPDrLj/DBfxLjVjmwwEddm5VrgNGDtGdlWtZlXD1TNnIfxy9y0Ep
1rxYnteQndncz5MXFyXEfg25LKhsT0FAwsp6v46YYXlkk24M3kATBD28WMyC
F4jnNAw43EwcBz5uWbSObpdkwDFVdK+UCU6ECtsZekBULSFkeHb33S86IjDA
RY7sV0NLlxQgsW247iUpa4+KtfNFNdEtUevwVhWZKL5AfI0JlhgZ4WBTyjof
BsAe9KiMJKSp03TxH1ok0/brseDRgGPMqmd0plQb/Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
df2Hhcvxz6FdW2sHQtmGLJEdKR2IcWECVRwM+2lgZahOma4+l+CnLfldbp8m
vFYvuf6Hr+3MLuwDqKCcVanTpbj2vmOmUKbWQkbFKaKmKMijQ4sDvakXbQ0X
LIwacjKis8LM9Gs90y1HX7FvlouVgkb/KMh98Dmh9ty8WTifHKGywLWsHEH8
y6rjTgjlkK2fCZw4fWGAg5FSnx6pkf96DsI3S5O2TnOd/+3dACVvpSYhuFiz
E+ndOOoCqMyo+yJqaZhJpXHB//UBUuUjF77dwg1tB4KA8IG3kz0I1GQZzAqQ
yOpBGFTnbCDLMRgD7Gl6AX2HvsM3iEpv+kJ+0ivlMA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
daa7iuRcOWcIikm1VOgNCvUsEgEJWULbbPJXMbJVMud82iVfSuOPu99oGIGz
YwAa/49zT6E4lTz95CqdotUEvftcqff7RlF11sdB2NiBA8SQTM8ZZGsn10PI
ZMCo7tgQDDik+zvM6rJKDI6ONJd443/I1FAX1nchuM09c4fl+2totGmdMlJ7
/pxcxQBFnlDUwyWNCk2pFtsfpdGvpXakfQBkqd4TPWJOgjFbgxh7aPWTZtEu
YRAZiTEc9/yCfGSCQftxD9iAeBbBb07QDWi5ny6hLRa+eAyb+IPk48jC+eTe
5r7uHCNmdoCdXgwpIAwffuzDzQGoIijeAZ6TQyou+w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Cg+0jMv/nZJ49e+MUt+RYuueNre4f6ZG2sHxmq4gTbLxpzbNJUv1F40rnsUf
51J3jV619Yk5wnn4q3IEy1U//vMI55LMAYJDTdExk4tuK7Tyr9/AYdcCIOB5
feoaM8jYsp561B5/Lyq1x7yywbPBO5AyVHcy+PCj6EjKzUII/HULhDT9px8C
hOO8OGVkt9b5HnC5hQOV4TO4LVw02Y9A5nm6p9GPAPg15NjREwRZq4yv5ezM
Ih9HGxzAFrfcXocSDBgJrPcyzTE/AO+3mXYbJxJboch4udpg0grBNAbBhSNA
xp/WH4y5FWM9K5Jb4W4CndLIet1Te2LbP9krIXFrRg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eFDMIOnZqz6Q9jpYwg3P+Hy6iFQV9I7lnTXzwL8KHLv/I+3z9K6SwT1QMMEl
3HTj3vienHh/KxDn9kW2hf7B2tyn7YuFrJCNx+R5dWljZ+/UrWD4fGH4VFh5
rv5QagRPtkoBZ8Rpq8LbNh6lkhBRVT7Y4J+o0xoCH5wiNGnTeV4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Az9qIL2ctZU5SH2ISxFwEOrGYZsLOOuSow1yLorcWXL60y4bPybeVjbqJ9gF
ppNV8nq8R2i/gZ8CxMYwrn+f5SnykOtYMii8C5WeFft12scTRKRpkkRD9KTg
3VI/A7gQ/974R7JLct1mCx39Ts85bh6QytggsVS1FrsrNbcQ3k9ut1K75z/a
t7sq3a5stXAAXdE2I+KdUWQS/g6c32+kuviS6v6JLb0/bmArcYkX3mkUBBMT
nbkNo9lPaNWUHyfnT+L2jYgKxLTwzvh47Usu8GS674920q4+ZIA659AuvczZ
xEZrAjrT98o6mALDZCWZR07i/MNoZCCuj+aUmkJfkjLd1pvjpipRJwZYJKY5
c1qba4dVtxbRADMPJ0RmkFkwnpJW9M4boq+14KmN9EU/+qbZrBSbMYwiO29j
LSn3Vr7BKGcLZCqpoB2fU2fhPwVtjUJRg5Tje1XNTZGSwGM9fOq9OyWXKn/X
i0vasnLzdNaQHW5YJk0G6nOfWwffcEN3


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PKw614k3leFt2k80kSVYXCHOAFxj0PP2+oRri0Mpsqn1V7Cvp5a2CAkXrP55
6ycIQzisj4p1/Vq5IzY/sP4/ou5Z8TkN6SfygPIYvRfSHGAgmvCdC2NVZK/j
HSlIGZQWCmiTwI/UTjzJbWWTGRw5jnzqELPbkB9i9At3z9F/WFE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nOrVaokcu/r1ONq0TSkrhJWd+pXM5X2djsOqmkyW5Q+L++9L2Io3YlvVEG+W
3d8OzxgV+CWd59K/XmNzRXLHyPFUnYPS/CwYvRkd1ptaEySjdPjxcrKR/pLN
uCz8ksMd88k2pIq6dWpc2juRnNru/bcOO9kv/H+2LyL/p6PGayw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 133632)
`pragma protect data_block
SxayTe+IOrTUmHyxqcF4dmtKvSHe8eMO72jX7yGtqYHRLJKAgiKOYJNuGyQ+
Ch2T/a7O+HxOpe3hP7lQo+dyBVdOlsjBaV2Ij74a6sD4O+YDnavPk7J0XOoF
AgJwF7M5lcjYQ3zoeXa528NAyWO9tBfRzKCXbB87umBFfZx2cNtM078zsnIk
FPIMMrB0S6og7u/gARPdTb+jV+JTZqH/POUhdNJ+rRXg3mDhzG82B8XGSuHh
IsXPYmq2k+Q9bQ/x7CUA300uP5CISJGQIlPStreLnhfXfHdTtw4I1bs4DYmr
/v+kkQBnXlIHw3hlGE+GgV2crdn+JNlfajUgKip+o04pzsAEYasXn2/Ybccb
Hyg+dOlTH/sTEupJ2lHiRON4VhitUcCRFaUR3NZp0NeO9oObFmhv9i4uBdtK
qVkcRuLowWRXTWC0/jHYnwm4zW8C8tXToSDLqZdeRCvwuC6WYfWCNS8ufnIH
Ckq1+ejt1icvnoN/4DcvyChhC+7TwG6CyIgs1IsaPAovBh1PruAxULTFPnGW
fGxXgO7IsCDjBpqwqbsjQvic87HDAWk65coLBzGz6tEZXdMFwxlsVngKK8jd
+co+Iarm7SqNQGQTT0apanu64F8TQMrvnF7eMgfxubVF/uCKkcMt+EIDtA1k
oVwZ3cPa75fMwqOik8iR1wXy+UdkwPBzP8TpXfQhSR6LzndjJEknqLEa/D6l
a/kThERiFqdO/lNpoUKM14oqSPxN0ol36Z7YAQ779pMxVws1MW56KZaMCwor
J5yK2mDQU9s22xFBL0088ghpY5ceJS7CvIwloLcNlI0fcHDiSUz2Q57RYMlc
zsw0zUpKmY0QGlkrsnnSZqkrML69AGCgquv4M9wNIqvK52zy4Bm+rdx5A4m6
LoHUB6qohVVaqfC96IFtCboLLWFxtpY/Iik4rdXOGW+xxYvjFBfZnhsX7J7j
qpzdFrYERSGkVspawLdOlBTXuUDfq85sgcYaT6FObQyNqieId6L2X8OAsEqg
7M924SqOWji5HR45RkIsaf7bMNd4wBCEZalb/2y5OO7GWhjLbNVU2NuzOlGS
qKHLZL19CHWze3Xzj2Iw8l9nhIidvLqbPljpoELHTS93Uqi0eu7T1T7Pr+Ca
xlccjtLXH1xfI5kd0RwK8qrGoLQACFRGO4AF7Oltv3eUF5biPWktiudWatSf
S6nV5McN9XtRbaRDlf4YhVB/XigCJy4OFQIa2Hv+sPTrtYtgGoXGMBB/HtfT
vKVTdjhW6D4x52VQHnJoxSfuXjWLmj8h3ABLGfNW6n3vrH3f429ICe/o3D4I
M1oiUhxBO2w5P/70GBFz61uStbengVYD1+c3EFXNDW5JKetlxnCw1iIck6XL
M8Fh8xzg4q8BSwaPYZ/iM3LqoYWTN28o23TOXCj+X6XbmfQ+B6m4IBqhLzKa
gZHbOiJX8/SRbAjX/BR2+DIxJsAnzY9fLZBet3u2SF4zf8sGrIc9LJyTWWmW
JehM3uahUx87aED7GAX8Dl1O4zJRGfvKPesZsM2DBEHQ5HC4uVRyiKCstetp
w0URC/wAbw8+bjysDLH0BN9ReRS6BK494lZtdkwNsd1AhHCBiI93Xszdjq4+
LVlu52YHVOS0iw601Du1f/jnfjhum6xEuBV0brRUXEFhW7+KARjaEk8IILWc
Ir1kIr7Mnp2qdHmOt7j95e8LAzciVASUJGNmvR3ykvAywwqWc4erhP3Y0zv1
tQW0wv1dDYNDfL+Jxi1s6fBFBiRcp91uNFkxFohr490D8KCggDQLui4OCd2O
KYvEsRoJo8+DjZ9XLaIP8f4wko+DbZFTn0JCCXVd53fChF8jqk1epQYnU0wA
KfbE6ngm35HVc9m/mb/xlSk5Vun3YUGcy8qSAZoA5z0MbqyAxWwU8fhRAVzM
2VD+/qsBW6crX6+UKmYcc+eaO0F5YzxcoBziSwm3CCooifGmZN1YIMAA2gwl
31yCwUbXfkvFtb9XnUuK5fDXkRiMTFIPhI+mL1XehdJlvtFc+4Jh1Ev+K202
hVTNvnElVk53qzc0J69Ysk3C0vi5N6xGfa+1a2lK8CA468swK3Y33iqYxepQ
dCh+ZifKeVnLyVSuC3GYrCoZaX9BP5GJBw+J1HSwmRGjo+0eOZbfNfScdQJG
021wm1Fd9r0ESewDfE2Dh8f4K5HOo1jHOkAtawOSMgs8eiP9Ke8voYIPzGVv
H9zx/6JjasVfGhNiBGCq3C7nYxtp0CjBrA90R8Eqz5eCP4AXDR8i9/SF/Mkn
wrd6UNNqNRQT+2McycKC5YiPN0yWESXZ8c4mUkqIbrSIKhjJR41bM6le90T5
EWG7JUAQV5Ljwe2PvN5ffCYroy1QFB0/p7n5k4yhlNc1AIut0wJX1UjmHGiQ
slsItmyOW8WMnl/8fexl/m3bSBNemhelrCResMoX2UiGIytXVzpsW9csEi8d
EBaiyWL+UEr1DTgl39PrLyhswntgGQCzLJSIopd4aqU4YKTBhwvN6WMzyPO0
akBq6EA2qealmEnsZeVbz9/wTWxMLIdzwQLoYygN7ny91O/To4bFixjKLk9R
DZFKxWNHXwojWXk3brPUAyba7KMSxQ5ueRJiOzvyxPKqL4GJi5Idx1QmgEkU
hvqvtGZedPA6/m6/GmqB+eBCExebk6ICwXP31Jp5zY3u9c30ar9yRfzjJyPE
k2B/wGhQKmyweXEnUebWQcoxgyUrGmh1St2vSyo88/rFbxj/dSixPBoPvV4P
DyVGcTJA0dS1GILdndAMrxfu1Lo8LNBsmlLAaiHj76zlEaChigWcfPN4wvoT
AN3LJhw2hILvmdoiXTdDIdeWYmyrajlePh2zEEVtj/0agj7oXX8/jPc2V57P
ah1gLCvAj+I2dGA1B1w6VYkr/r4/YOVwufRE6cnFCS6F+MJP47pAVJB94CpH
VidHMI+SaWiKegnEku1qM8RxD8N69x8+5wIuOnP+V0DoTU2hDgI4J/PyPerH
E3QCSn5+wWzHctMmGyvS5tZtyDnLYihkJvEPsB+rSy4UIMgPfZZKDMZnu2WD
0jmzq/wsoHIzTJNumgeAoDgGujFCdS8wYDWmNN8yNdfBpAq5mvDsHjl6QCOJ
t3j1kyGzaiK138qRXUxtbMLo/oJxs8NPd3B0U1qVMgwbreseo1SY2LLpyuO2
y8534daDJE3F7FYBYzK9RotjzBgPEsVQTVb809SUYhx3sK4N2GcnIOgH29DS
uzV2LJRqYBiZH9hKwLpIx3bPfFGcSGcy+3wTdtLv6jhTfvKE8INhI4eMg92m
/IXu0JHSX0a3Q9QCk8FpiYD5v1m3lfJjtokJb9fyCyZ7gjV9Zodf8i/OAE3z
Ic2XRVWco0TZafGGWPE1UcUMRGQuMtGfLii8h8rMKkxViDMPb6jeZwFlW7R/
5daesdO1e9pLeYHbhaqKLVGaySLdnZLY+XmNvKKgsQxNh6xMGKU0tBHVkV+b
fUbipZmUUjQNl/BqBSF3gEGlVcgKu67OmoakF5RMrZAoD+fjGJJ35ni1cn1i
/Xkk8eOvygodE3JEOtm42S9lvcJKFbgEX+Tgl0rZGg5gxRPLk70LWForxKP+
YNGdYdONI010JDt5giRDEEzI3v8dgimbrsn47lBGrTbfJgW+unS4xIS9D39Y
F2sdVrqHdq/hHpbLOs4TdLk2vc53msSwQa9MsRMXUy7fFlYXVUExjwFrFyx+
xT9aL3qpZeJlzw1RVTrGHwGJ2pvklOMEKSw6cG+5LZwf5mos0PQNI8cQxSVc
54PLLLz+xnJwyrAPkOnYSo9fo5yU1mIk8wT1XP7SLcwvQfDKEm44iOmoIILS
VbBeFFJpTwYGGV1v7JSMLLRbkHZge0oI8JH6buqVO1LnkfqODUs6KovFk4YF
8VONTjDPeywTZmOUfdIRfxkb0HhIkukCea4ib50dKBjvAnW+cOEP/XldDTY0
unApg5rKq6cxNVnhXJ0SQcMxGpFcbCggOEdEB3+CT9odQc15BCdkhfCrntkL
Nh8IFu5LVPO1K+g1RZPcOo4EbBUXUDwuzafOYuWKuUy27USgwe2ediHbhfgj
p6HUYVr3d4ySbcBIKmyP1fCmOZKKF2ybIUPAqKx6wI3L7+V2vWzDfbzW7bEb
J6+D+nH4OD7OZO9NLfO06yuD1tA6sSq+XolnR8U0d/Fit+Mdp7BrLx5Lt/WM
ci23WcuH2IjiqX2vOauvr5QGsGQi6HU1htP5Y8S2nbXuaBP0So/6eRx6YFHf
/wjkFHLKEZ68FH+NOzrrUu1djw+wRQMReqXzQSWRRPONzKiKlfWYRpAktbt6
URJYiNK5d50+Kvm0swqoi2mAWe40s91dFQH2CssxaBFeYuSTwq21M/SLDfOb
YzSpgd07Gn0RFlBbE/szvom+1hbL7gKzVgrsxgDxgTw+0oNYN5wzh3V67yUL
80gdTLloCJioCHvvI9ThhfdT000GDffaWtzlGnPDA7BxhWcK5oaqAcHQFxpJ
APRFZvosdD7wOLwyqvIE4Iycm3Dz5Vv9PjMhovniDuXujsydcfv6Yko+5zJK
FYHg/D5iT0adaBKWVhPZnOKgVX2YJzFQLkkpUPDQrnag3//r8WBC5gl1bhAs
iSQUZadTB972ke7YcUc2NBIhdweQTt3T9W5ecsajrXEN9xvFUZx1GMwILKK6
u6ZQDt0/VNubuCReizSC/n0Y83bEoFAGiIhq+JfGaXKbD7LZXJqJ1i+3HSPy
2l4BlRKpVPw1F7bolwub5jo2YBNoIS6izIfBl4HG0kgmZ+Qe5iRrVpDHAe/o
pAaH/jmTgEIplNqcQpdy0vcNlH7tCN5B9rwNlzhFiKpVlYRVht2DtjimuhQ4
6FuZmjG1T7uhVedLFHqotcJqL7WmSc5HdiDUAtb7SMfv5L5EgBUzu3UOkSG9
bpxLzzefMaW3gTKEukX0iy6ytjqYPXFS+P/YxvjIN3bc3WGub8tNB/BXYMvi
vLbw591u0fqYyMcghgF/7eTo89ZwTH/NCMD03qvhz4XuoiPmLdYFzMJZJHtt
A8Fqr2Tb8CgZr92N2P0JVJE6qt8JPRWVx3EC2X1j+MEGgOIoERBQZQVlwbeW
pGgVO0P8GK8ZQVWsdHv7H7rQcBZJzS+0ZrBpRz/k8oF+7edkV9RZfciu2bZq
zg8GrARrakg/QfZwQBiivkAZPtj/AptRzBs6Ta2kzBQJAVvNXJPT6Igkt0kq
rzA0txE/LlzdKGAjMiO9d+eQTZzrfrCrVxkh+ZaRENJGgcg/iC1yqnMkmdZ7
r6I+fJkfHshz6Uy46jv59INjJriOQq8KlaMETM/jxXGsS43V2UMpMkMpjukx
AQRZdeicNpzmeVtvonPjARmQQf/ZK6vpWG1J51NnisVK8w/+iayu/KgHA/8Q
BZeCbMoIzMhIVj5lRXHiHqKxXO3rKvySID7VpbPIGn1E43u1YIaOi4vfk40r
al0ICA3TRwq/jRRi/thzSUIHwjxL5sEx0XQnZWnN2dBQEB7ODMrThX3ZMw0t
rRjtc0GqJg7Dzr7BbkgYgh4By374ozgXESNcBAdJOsLOJd7IdnRtg12bHQhl
JgtnyLqScy6FXqHHggy/B9ojcKsUD8VxxpFctVb6Eb247PP8OZ1lmr5W7T5u
6XqKb5jgv95cRe9vocH9LlyHbkIyCC2Xne9eoelboEjAEcTRLXbb1k6C/DB4
/byDKvrjVLaAiTC9Gbqpkd9P9DAoYSTfhscjTmtp6AzkfF1QRSzLg4qSq6+v
7OcKqERXkmWj9H0B5wK+SvFP8tqgRfNiZzoOfu1P93EikR0rNVMDIVE4VEpi
zNOqpqnlSiJZbvQQzM/6pm3akYszUvTRzDJLhA8Gpc6zPiaE5vp0mbhHs8n2
nVjQWXsfYK82UYRBQnKIMldy+ypTHQZNdSPR2ygvwIXl5Zp98lkoxYNmZ8df
c5xjgSPjmErmadJd608/qxVYTvBkBAnIuHnhx0AHQPs2QKND12QKsCNcAan7
JACZ+nTByCPQg3Yqncox1PSP667xQmWAK4iCH2WcTClenFFJIRicVL/ZJHCi
A06GA6gT+641nzKvM8954LvDhRtmAj2tkG3zvci8HM7orTpAPTZoiA+DoUG8
ikIR2Qh+lAgeOXpFhtKuQrT14A3ySpHXADTnNeKtyFrZDy2LgtoPd4WUyCkY
O/fKKisXG005XgA9PGe24Ytt87zoPPNbuB3/uy6vjqutoyqf/aknrV4K5p/o
7K2hVRam58PFh/ZK+caO6G1NAcPbq6ZM6OPbiJTfVEkKFJe+XnrrcMm9oT6P
BRMRmBXHGbUea8VaNjvLu93rPLqKZKhQFGd21OyvwFsdroazyTd4TJcEoFkT
oc8T1hbpGC9oO+N/5aYjxlarv1KkETc1c2f8GxIRXnqdWI+/UwHvQYIPTXD+
AkTZWh2AOjHzZuWr/CKEQ8eGPFP2TMg7L0j6JIdcQhigOC84WTKf24v8xfEs
wvgmFXxmaAYqHFvGZ43wPsK/myWInqqsc2PPOiwX9DKwIUcPTtVHhYdf7hkq
hgBp+ssheEsL5/opNdBxA2ZlfNgpG9rz4JfIgSP0JbmDFuhkwcaiSta6GHHk
UuBw+sRZWNUvcu8cxK1LIalESHAHP0QTsD7gWaxaWVV++ZOb58O1gRhDw2m0
YsW5AYzFmYBicxATRo5xvVOMaqVXJoFECPhG3ywgR9QN3OTnXwgyyJ1Rfiun
azc03/LmRm36q8YKfdgpo5jICncdHbSFNJEs3mjrD84F/OlVYvTd+ZQ0JCFU
NXzNokQXnNmnINBuYVHym6qypGVwbfxI6a8ZNIPkeG+1n4mtVOTIZ+/KXk2K
GIwX0Sj2+FZ3YBAT33gkTnXGsEq0NeOuezxVNxhTI1BxdHY8IY4KOYy1g2cU
Yk74c6So4iwEcKAuE1llJkeLHvoHUmWJg2WfJROjLM7iMh8tos3bQTbuKQAT
wrWop22xEUTR/awXvp99eYACkH/VOXSrRbxnSrAPwszcLlpy39PCHfpGDMS6
DkagHbkwJoOJgK1Yskug7PLJAvhZCCQ/abtark4PJivwnIIJMijRqxAWH868
oeDShxLzPvLg+jMGoFPqHqHDlrZkuAPHi3HSt/4dcYAhAfqdv1iJ+llJMqCj
XwNSBQpgHYxNI30MXVPS61378PmTUH/JzUry5NADs1gj0ROVePcT+t4uUlKW
Gq81ZpojnU3uJUMqW0z6/rztkfLEDYInUhoFTE8gTWbspGlM9cCMLK/ISYDg
bY+PE4qJejmn9CyWYyCqSVBX5BHgtpUA7VJ4rlDEl+josOUieVZYvvu9CSRW
K90Ez4Tr3ZHsbUgfP5V4IFDSiCBjUr3B5FTGyDonzZ1hk33U/rZdWp8Xp6Q1
D1oCLZTBhV0GniYh++quRjDJwBQnOgAndEQeSTxQZBgAuuLcqSduVA707XPb
WI8SPlrxUY38fPDDPAkVJ3zAH/QFeM9imsPjA6LeT80YINP5rjwVKb0DYLKL
9xGK4y9uYbh1xobxjUiAMKILO3ekgvXjBPxAIggqGR6RklpFC7Px6cfUcSga
1xWRkAUtLehSg3hJE+CzaZpnvHAMB7fI19aYwiHCniaFVA5RoShEJjsI6tDy
aXriuCkeM7qhTtUoZE1eB0z7hMqkYrsNpC6DA5F9HmEOJamE5Ua59VqM4W3L
OKc8zRUzj1PxTQsCuYg71NhRGoQG/B+g8XudF2ybRnDIYDsGxiXt5b/0yWzw
5ljZjIU/sua9OGYevAiXU5d9/BobFI2jfj9sFdqyobKgHJcd735EGU3P6ArS
9bRCoXahYsZGF+gSczVLebXjj32PqPqIauBchJ/figCodZ8K4Ngzxbho2Hz8
maeZhUsXbN3JtYXGnqKcJi0+Dg8Rdx7Bk80/LSCcdp+cl1NKHCJCJ7Yju5UG
Mrf6Lu+8fHigYO0j7/Z2V2yAYGPugl4ksACtAJMHl3PojWDfB1tXuqDfMdum
RTnSbGhEFbbzZhU6zWBdKg8WYXPaFwYbG9Y37mU0qxdm3RUUNaW0zj9RwBPe
H7zjGm1uKHP9Qg4LOlKEvrKPeC4ABOWzzwcaQggO/T1YZicoVZ7pAH4mbJxi
FSReaA6RhHWl2VVhFbEw366NIBYvOFU8odJvHu2lJbkhus6Gao8+ZRNiTUaz
eS4IqZGSEZQsJSh4mrHWS37wZvj120346Kj5p6AI/HPmm+xnXm0xmAXgjVbK
Y4I7rN4qM08vOMSgmkn2eSmiUFWr29d+6yNeCMlf5ehEetbz3EoTBdd+1GjS
Aoxx6fsZ9r0Y5220ZG8rfryk3bDQDHFq9Nx+QC0o2NkCl8kd/tWkPfigu6/2
NlTC08bIKgQGE3bEbvvkUVhz+dX8sW8J81yOn+rDZJ1uYJxCtBxgg3tLTlUJ
MNsT9PwqaAhr+5reyHh6TlI/20XanFhBlHejX01JNZcIqIsYO71/hZfYnn8X
giRtuQ5gNsu39d/WYD2JpdmPidngAH71qRgxLva2Defh2NYTLNvD7nmd/srz
WzHXfrle0FwcTbJwQagwvzZje+UIRt/kHbdTe9V5PbwTIHhq80wUxthx+7TF
qKA7E66PFgOvnYCihBhIO7D7ofk/5Kt35/V98rR4C1YrxVS4SHqiX6OT/QYf
Ul9HsTx91qhb/VCFw4MM37dy4oUOhozVN13SpMU/pk+Nx0Zw6ItVaM7L7Zri
u1GdmJ8KyP5sIYl+ay0f6wTSSrkJUDhiIMBDXhCfP37OA15UQ4ErvvhUuszT
uT3aTDBIttqQPIzk6lmrrsNv3ojbcUdVmi2T/eVsS0mw4bhZ4zXdSSztfGy/
owymaVwNkdq19aCNXOasFaEyBEUkpJNCWnWxHCztdUyHmnBbuwSEYAUeMnGX
ln3ea9WYFGJTyGgPdduGW1w3/+OFwcOVkn8S1mQIsxSJ3Fstce9XwHLMC6I6
2iIjqrzH9ukWvEUXh49XjDp0GCI7KoLSSFnZcQX7ZjiHzWKkHgpKU9HA+umN
KSY3ay63BKo4hIjdB/NqyC8n4L5Reu0oRDdtUj/viB0veSa8bm91FaX3RAlF
nTC0oHwxVx/Y4Ojz6pjWlImgXYfwFuij59lCrpJClvtvZ430hXrDsAnmg9QU
lmU/Z7kvXuJvFwwIhgYVOkQyVHU3nfjKPPqK7bp1P3pkDAjRyoon0q+oW+4C
nCTt2oD8AWsUwsQ0OYUxOGcRlYLpW5j2porVtZ5x0Tajhfdp3YsvW9cnB/v4
cehOO8cuX+XaxMnx3OKtK2fEfmkGd8PbbTVXLtd6YS/Bm3v00KbElG1ZfFUQ
X/opYQpmCfjPBlMEC6sjykcPZqnUo4VDzdZTM+ZPxdCz+q+f8+C3HnoBsiX5
ndlms7PLHI+Niq0OGzsTZoMchf2SSAovIqsSz9eJjlMuRIJUXUNiWj1d7wQB
O3OCjXa130YZjZK/QtiQEvAHdy5uaCCJDPG/ngsWF9xCS4VTZ5UdIB775Key
oZBl5sBgTMKMif7FM2O0SrLqIEeL7svmMvakOEM0xEvJX99MaRFKAI4L7mbo
Z4GVcrUJRaOo0Xh7rVy80LfDE/XhnZtUXpCF1SAFJlqZlwYY+PLu3JrWjkgt
Q3CGMzIj+amfWlnRgvQh2AlP8jR/9DpZv3auZ8pNYJA6zgMDrz6a77i7TMI6
VF/0w0oGV5oTVt9beA64IZI5xRAyajN+Dwv7eUcZi6QPZ3MMy3tzeMk6eLCs
Q0qasNzbsBeusU91rR7URE35ubJbL4gsaUojBciOdC3rKkab+6LpbXpd7xkV
wSJVFNn5wBWb7nEn2TvYAaMkJRULQ9hTRqy0wqEK7k2RQDMSlsNjLk6FI88B
8Knc/xa4H91cvPA7HSLDYWjags1R0Jf2VgICIVzM67gNaS3Tzat3Ies7T6lu
oyaYHmkCXaHd/PYcu2Vl9SwE8bY3xyRRBWOHdDhAalsU2tiZEBi4+eoMrb4a
+y86Lr4hyXlEIOJiigsk5BiZfyz8rnVGioAQiK0itQFwf5/n3aEgtCmARYAY
31Kb3aI8uc9auoAiB3xz/DWvn7OrcBtFGE2M+RGLxXd5zSjLxsbeNrD9AiSr
96HIDImhPX2XSGPeqOEm4AAWS8Km3ptVFlstbFlpUFK84kI3UKUUWX2klH0Z
C9e0bDv/bZ0uzUnywfxRpHrFSxphwpygJ85/iXQUN4c+FEGnnqu47l/Fbxie
msg5l38eULfu3lpjO46tVIPeJdWezLeX2UsA0MKzHwQ6LXuDG3UtlPXd3dsm
LaEgYkBNdkbjFlrc1rm6ijhEYjoDhaWOfEPyHnzABYFXoSZOk1EZMWX8dR0c
7UW7W2bVeVziaGIJ9TrLOVv0K9vOS5hczqnkmLF4XWzR+PRxGrCy5OFuu8Gq
DJvWSwffqAzdInF8Ap3Os2cfBpSJ5+Um6LTTm3Ccxulenx5+LYmj9l+rxLlj
JVSj16Kwg68ZOq9ThqyaZ9RDjtICT5lKyaD5/Ii2l6UXqJPKrshLHuVES+D7
+m9vLQN3qNgiqrKibSj/hh6PqK7bGnvT3Or27bKLeK3uRPQpq+6WyNN+WySw
lSSlwI8GIxjX3zfXVEKsma7C+53UVikwzZ4B9wlchho5nWltJCxJNXDjh3+9
VPOpJV46mdLtPjoNKMMWUzgMwJw0QUiVoh+jcVx7JUfg3XX8ku6xLhrWJK0+
2DZZcjLw9McmBz1cFC8Y/3zZi8Ia+63hWm+A3RjenT7d06f2tFN9wgG757Xa
rR23rO9HYL0F8z6roApaqlqHUe6/jEGD4BM3B6kxYXjHrJplAo0iSdMyG/9B
NKso07Wd59DV3c6mLi18tr1T4FCZado78yfM5KKhG7Cz/pZhubBXO/PJNPgg
JTnNEM+BiSPK9RpohtIMkEzOGf1+86sEX6xGwkpfMACNr5L5cxEYvmg/EmmD
UJfa8fMhkIjdYBGyg+t2rxhpqa80qbFIjZhOjPWMba/2B2yj0907/AZoD3a+
57r462jTrsHKdLOsdF5d9lRZl/+KM3vSwe6t4J9N6DWEbQ51MCa965JFP5G8
rQWnZxGwx+2y/1A71MmgeRYxeMZGSBMMgPE6J+OD9SHv5bsDTFf2csNZC2Cm
xv1BBuiNxk4RyUROK+dEnG5G+e+ej4Yej7uI8oSHI5ARr2Gr3wvwgRBx1wsz
Do7OgBbab3+maJO2x5GWGqf7QN9RrjNsqLkHUTAVI+jbclyUJMn/hPbEY0nr
by822ptNLM5jWyC+Rg1LSZ2rgdc0bCf0r7JjEzmU31wuvXGbcacY8mBESxTx
CpXzzyNrCbTDvPERQMn+0Ou/wYx+L61z9pK3nBE92eJ67C/kh77dvuSJHWwl
4fWltZv8KaxaF5UVdVFqu0w/z59R91QzShefxoElh4QhNT1UUmGsHzoqwys1
dwxGN1d65CC0tcZVhLCmecx+qQrj1sPLoeM2638FdpbIRKaZoEA9SxDM0wz8
WYL/x/6eFugV+uhBhHb3nwH6LlDx9iq7+X3mviQ8JIRNv1h3Jk8U4md4WLBI
iuQm306NBAO7dZsNQpXQXjhXMoVA6O0Ro6kbc73niZPwXpDup4fuxEiOFHQE
uguw4Ha6H7DkAfuhYCRYU6S0XHch6BiO8zkDxcdTKa7LIxLaJ/eUNPUHMvuS
Ob3zCJFbwozGZ0Fb7hoh4YvweLbBuNFT4zDgWM6O1WULN1vukYFhbeeKZTR0
ic2gDqSI8enw7mWoIxMyQbO9kULzUIqrC6+GnXqT9WVqz6/XQkrGzL8DMjVo
yNl9voAnf3zsgwctuqpAUjiX9UBqFwz9VvvMDoSI3eZSwsLYgU9WUiPnyswA
Dmzh7HyQL2AkbX2X4pbh5ITAeXDaeFwAX2vT4X4cW5LrLz0Fs2BJbcVj/045
DC+/C0QWMKgEQG0aVtOIm99FuxpQZXLiJN4pQNH3rEVePpeVfys8aCp5wDDU
CYQPspfDs0Tkr1uyqDeM5gUDzszR9CuC4WtXljCjrHFpxLvxoGJ+NUnq6WL6
oNT6n47ehbQkA/kD0oDKTJXQTK7OsAgONBzQBmH47sX9lb67IQzgFUmts0xi
YBo3FTjnLNOrLnVPK6shkUYG6oWVTIbwoe46snCUDHhwAcoa29pa/YKhKSGf
+KvOvYVc4S8r1XCXrLs0AfVhlJ/X6VaVXTT512cAygwEveUZh+hrYTz+yGmq
cj1ngyIbbY7Q3dFUydfy07wXSMVHKaOw47dunCPduHvrl/ImtcMNawO64doz
wFZ+GpE3fFGPICmjVTlpnM8BqAKK29Hq9J9YL7j3orccAm9X8C6Y7zO2ALV3
0Qdbs5WE7y2ZoYRV9nSSsVtgzm8rzSde6wPYK9z6qMHoSJCn97595Gq0jCNK
FTB14c/EsUbK03KhoqnADwZwUbvA5FU+JLYhomYVRXIq79E6itLMhtxTWoXn
Texly3uO/KUmOJEtMGh8g6sMffuE8IFszyg2kBMM7bYfMDoRj1OoWvRkOdU8
nBuIpE89ka+PEVLgROfcv939NbHXTp/5s0VRMlgDEgp+KTsSMq+xBqrnZTJS
eHJrBeWJmmeQG+SgwAyvwtabJWm2eMQhtiKtmqeJu5zqSV7qhGOZw7E8lNbG
ACKfHWMOdITWxIRuAxzFLMMNTnTO/3lnLwMc5xdV0XHnv9MxKurDynf0G9HN
pNKCVAkjpjnbabAXI4EpGPUQA4FvCiyT+to4AjCvi9DTFLXfJU2HGbsdHuRT
VzFE2rmnc2hJ8V0dTb3Ml84Rd9FLNanfGDHNFmW2MQkKxlm1l/m73s+FiZLl
ZuKUH6aJWJ/83zHKt4rYk+xi4f2fEjn1NVC3AVhSD5iqtTD+1qeWMmd7LH6q
gmSXqDlB6YfrOoHOJ0GxuVPqBII6/+7Z5fURP6awjMfbgiLPEcABQCa9vEcr
yOQq+ZNrVjrZ3hErHEccwvVKlKTRFySqE6SvIjk3zmv6OO3wPJDDB8xKm6VY
BWkV1hCjAeSKWVG2Kw3VIRKGHAj3Snz6lBAHDhXkDMnM3k4QF358EsctAako
X4Opz0r/qW7GWNCbSwCqVrmANTMssbFpBcpkd3zLQVRWvlhlzKI5Qq6/pL1d
6lrb9b8X0bHFp1ezGFBisHpnVDex6vCMzixc/5IXiGCsth7zBWIZg+9zTqi2
7FpjqI6ID9mJWY7wQhSZV1JmAMWuUVSNx4rItzmRynCkV2J/C0PEGWPyB5fI
dQaRGJN/C2S1xAZpnnOZpBGnNbRFh+jte4Z7A4lIkMtwJ6bEinhPzOBiDTB6
TBjUVgQMd6udprkdBbEuS0+wqoTuqTJYUCWRtcEzJKr7cBeq4nVtYmwlZYby
iG1oHEsa8oeUFOvkHXiQeYav+4l68tRIxEud7rrtJSGr0fg6uL2r/dBpxT0S
k4eAnxUm2CG9FdbqS+lDX2kyY710WA3bgYD3L54Zo37puKJLo4tQKBT3EK+b
M08gjbaDEF64mJSnLIUAWISLJAVoijQqr5WhKjFT9IcWByYviI31keP0Wbw1
me/pxSEgWXUNbB6yLPoruGj8nnO2Ezx7PAGJ3N0oCnfj2G92MVcOQuIKq21m
gyXIK4whV6lba971QK5Ft+z1BOPvosdjes1YZ8PFaQ48TMTioYdqYWaV+Se8
uBxocdsNlcjM8NYDa0OAVwVuOKQFqFyVezpwNwJ5rSzEkiaVqS9ONTYCD+Em
r9ZDM251ceP/a1Zh6R2In7y0YZYYUo3GG/j2jW0DzQzHSO2Nqu4DyBjV50v9
h27Iyq1kxV/runDhfxeNE33FKP3q5aUEkGmqQgzddj9v/xjOMQ1xWvXr79tS
w9Ot37GLNp+moIOG5DYPtp+Lx7ldgjghMCuOKcqPFiMStY4wLThn+t0xc4Sz
n+8pwcST4TVGeOYJlKANG/J070yVBRNsD24g05ErTfU03dLMQrpcxqt2JRtS
9kB7lVdfxv6F3YCyFjW9y2lOItVdmPlJITkMzm4UFGXKIcWcDjeQSWamnaPH
FwGr2QZE1dmyaarvgo3OFpWsvbEdJQZLbKdomVH7ljpbh8GpPlxsfJ9fxLjd
godPLltopIarsFAIXtkrplnYidp48OFVVMZ3SmKIAtI/5lBQzUjW2mNCiESl
ltfFUCrF6acc3qgqfAAeO03deNcQvK55peltVjCGFZFalj8jAeMdRmM2DGG2
3yJWTNT5ObmXcXIu8a/AjRQQRPYMm/DTKyhDVnHNo+NrqBmouE0LIqNERprl
fbCNpOTs3N5sXMdsYjZo5GJKY9m6+i2oLbK+OWcEqqhmaSPRGC6L4E639/io
l3u2vGwdpCLocSUgV9BdUCAS9L/xPR8fz3360z4eA4RXlzHk3Ewj0+S8LbPo
3V2UFjeoBRunYrf73VEaf7TiuYwfROBIQjoVNqCrcysB3dub1f/+qzsrUrcZ
7Saf8UtDH3/gfo/coRboVkNkKwrmUYkh7szCsRJFA33pyiUQGlnxvMSgada7
t2QzUyaTzBchYNI3xyApx9wHqEY56vYvvTomJFaJYYv/Lcs0a+/uzbp6yfQt
3U0KMFXRkPyf4R9SGL1k4OoRjMM7ta70AN68t/i5q8esapUHr+PAuVfDwj3w
7OPM2a7sXg0uGilW5qzEhSDJ4iMPrlQlu9pF98nzVsnW+GB7yksRbCE5SuG0
dcg/pZ9Yqzg4P3ZrJlR0bOtQOT5hedAcxm4sPTyzIOBA7unxDLxzHvD9y5tL
16xY76+pW4WZLlvORakhu0O4R0aIo9sAd5q/4QeCJErl5cCvpMKKFHL0Py3m
cvkl0I0txMbZpHzUDuE2tDgt01Rghz+HjyVM8f9TWQRJ6jgagTG9Mri2SUYs
r8PXz0hd2rkrW21w3SPo01+QkAMeeocGTPaaKYSm1XfsI64xuNd3r6qVf+rZ
EcNqb0keycyMzhZJ2Rlc9HDwifnuqKixrAR3ZL1Z5znpyGjH61BU4bHmkaw6
1ppxAoKXrPQKQxVgX+1hPCm5htZ+gTOwNG5X6sLIkkFlDLOfGjfCEMo00hDb
C6cGg6NUQW12utztmdf/WyZi6rj6y/R0B8slFieaztR1NXmuMaDE1k1YCxLK
aFKpWqgC+u4UZC6aiKJLugcK/eur8dvJI5UHxoBKmMsAwz0EqX0hV3CaJsOC
uDdQCJTi3WSmxyrAZ7eHTkaWrUMWGIScsYJn85SxQz0rxcJTqJiH06vvC3X9
KQ0VOBQGoM0ziEhiZSkO+126AkDkqVn4UDgRatDiZkPTFff/APP0/5i/Gl7X
FVMBzdMRJy2Z8vlkNeVk0AzLAfPBOk/mDH/yNR6qri+yfJsFa955vNCJnSFv
a1UmDlooCFYTcF3TxqHvzjtrp0I20y6ZOKnZn4OlowmXW70DtudC83BToWTu
gl3OAu/OSGxCxop8VPcpatN+3Wi8Nsv+T4fgvHkUL5EbBqVozh5EC8NDxTa4
BUc+UfGDLpez5JznCdTcLyfsNyYtnFSHlyA3XmtY+TbB/VuY+5QRF1m4ePvs
7snNvEeFmFsgrqmbTKphPMtihDgDnYzH02jxyptHTHYD8Ys9m0LHRfanHG+i
/jP1QcpQxr1bBd1+567gwaSIA4czc4VJij5e3oErTUoWx3Lxz3/0YTyS4t4R
E2IyaRxFpdEoFOS9WNKaWT9KTTxmrlGAw/Q6GrZahdmgb8/mgN2tHPHKHE+q
2DEb0TKTBR6TEJedAcdyGeQs1YSaAAzx6DpNRduIuNWlQ7pSBQDuogoBwnpb
3AMw+rMGOYbMr3mTjfCZ27N62GrhEK9N29Gdimw3wyJ7b/z/N8V+Z63dyy/O
mUecF3kQ8hSwk+SE/99dmRD1cOLFOHL9v3mkiL2BByI+lyL9ow1C4+nCVVaC
nD30FajNghECBLOAS6+Sb/Yb272uer7k49ZePwNCfdnKnBGHx0WS5of/qbQ4
damPN47JBBAhJn6sgGodlmEmkwxakSWo0rjg9bRcb14P+wlHXttncEi7r2SJ
S5xXeIh6HR4NHAutdHYnJ4B0J2/r3khW5jG7y73eR3kpdG+rxoYbqKDQvPbi
p3+AoDOXk+aU0vW83nqpOKq7CmS+Ton7xh7op31E163EjYz2AOezsFs9T7HA
hsygx5D3VbyUfpn1Qxs5PWcA9dYzdTmMkSZlOkAfwNQb9uXlT3ywNJUxwvwZ
P1BvHHPh3PJIxdyNEp2/VrghJpY2LT6dXWQYru5kIEWTm/ZvpbG8+xHJPOT9
mc+H8LnVY85Rro9JZqAe2ALX7QPOdqZQHNvTSJXLG/s4LvAFUx8OV7EcjhJO
m5BFTtxcaAkbyy8YV2PJclUTiDRmpdnj3QTgsyALBJP+ZnpW+4ak3fx8SJpD
9vG+V+eW86h6CUMKnhTdQ0XqsSUYUy7cy2J8Pnk+CWFcQgFMUF3FxJEE3BUq
xRGmX0bJVmKzZNLpkgb6CTGJdSM4Nqabsn7Htb7izDJsmmDZJDq8/ae2pshI
BqFSnHdJtyuS9HIaYK/DNWZ1z1eZJE3MraaGX3XjjL5pDbbbXQPf0oblQgNd
EQbwd5blao2oHI0BfiIuVRxjpFJldvEKtlxgEtzJmComi0AU68VUhrgyp/pt
X+HILhCBgdR/C935Cmp1BtSsdQyONpJ4/1t1xpeFxUp+ExgzSIk1nuZSizOW
NQLHZa1WbEbs4aCVzsQUVDA7O72glqjMrbQmom1JzX9x5QZ5NNIHswsoRX3R
PaBodzC1Dp9x8syseEVtXepM9ihwO0yf7RsWKDi3teA/LnQdSHexdCNlSUtc
5uqgi2+uUTWnN+EnEdgNqTGbH23F17+904HLlwnssYewzqwpfJ1T056qxJTy
Id+rQh4RUSZcVoUJCpnDVVSBan3WNEuEP0kflxjqgKtBF6fXBvQzKcbG18EY
CicqUjdYZOv+Pq/ILlkQ9vxHn/hbfFXGn0+G6oXsKZqolCy6OCKf1A3WEQd0
JU9hxa8SMNng82VNPH7tAaQM2zLykboganI3ULBPKm7Lj8iSXhQFX70uPAG8
RxV5VWUffwVIoLl4Yry34Du7d3VwVrLyjXAmQBOrqlvC59giSpRh2kOF/Gid
j32HUHmJ4yQOlzeiHtZu3gtbVaMHInCinqD+ypyg21rKTZ9kBIZfx82S9m11
Rxhlzv0dBjcpW6hl1DJd5CDP2AmnGsge8PCE2FG9AU8iISCc3TrB8znrr65U
e+JNoPTE2n4eWjHnBddeh8kCRXkt+r6IJjEGMugHRee+czTT6QFppLgqplm3
84KUw1zdR+wBh90v5teivoLwR+/l4VgYp+lvOAPyo7Kzg5DlKboLj9u23vLI
0Z4g43GYrJxR8njB8fTGNolRurfz6g7CsXnWeXUXnvYHlfLrbD0ig93+MDzI
FGrC5qXDygmR1NYlw64eGuD+0Z2E6Q8kDy5/V5rxVqoLAAAza+/W0w4zFWv3
38GU01RgG9X7z9R6I5qnLwZUpk0fmMGeScqlGP/4n6Cwy4l9TObRhjP351yl
IdPUhp+q8iHIB0ymiZfSR7MWlSgR8gSlqpPYF6KPDIzIOokQqa3/fkEYjRMV
8aDEtSyEOrpEmtol0Cx3W74Fx29q+4NzGUTfU2YyUY6yRVe2awntNeiZAE+1
exxbXg9QhfwXDVGNVeepsle2yqce56Fl8VQgdJ5pletdi2Wm+JLvNxhVxCri
2oTOqGN7e6DVpCp/44pLvGVl7FWjvdb23LFRqmTaWD0Fyfpx/akdHOqIvCgn
CEN29k4oZAvjR2YH1TJl+wt5b6BCmWotQtvuBCDH1ch86pQ9keYDCfo8SDBD
kFgOb8Iik0/aa0W5aVBnFx+6ZCkCo82ks1DgbsFAjjEY0LB9DJAlWrGYHVMa
Kd+K/qv3TQRDdGkzgw6KbourSfg7IRSLvBry8hCXn7pTIHZXkSF0HY719Q8F
dSD6VM3XWgXCNRavAzarGFE9YxcNiaO0ywIXjLlhnpQBW8fcS3ZAkiEE54rL
k1QyKB4JoMRaqjlRr/c3NRHpcn+tSyBKpjlERwfy4lEw5p1CUEWWlh9fj2+1
jAA0e5EJ6poJJAF2XEbf3ta1MDjLgioFscEHjLOJFgAJAlewOzkANy7Yb2+N
rbzRN6/sJYUNT0cOHbYygmMbIsVjOeEr9c/0O4xh2lRN32HxRfDa+M41827t
tiGb4C7CMxlt+06P+v8JG7pxLEUmFNmiMTvQctL0NQwIjFvByxevMnHPAZiY
aSzFdbVjPok9ANT72B349Lh1aLikTZwdj3Tqraylz3LNhXbbvP4H/enQyULh
z/0qw1lgNdyfK2rjQ6oXfKb69kNmVGkiKeIQ+LtNF+Vh3mHGqmawiMxUdM1a
LhMenN/2avpRifab8gAKhvHV2jZSAK6lLyl/zNM/w6SDvrJMCGerzHOrpkmG
3p/KAtH1+F3mh99LNDVLwcFY++DK/9V4LpvtVgGHw3hfeeBvaL2GFpv4RCY0
p6hS73OGi/QgoYfC8r+L3iWGn07Dy9BPmT8yVGuz9UWWHNpaUY1o+Bf6yuP0
wK6hlnQRx2ATtBxqmkOwe/1dN7gxO/vtOhq9EbUNrIjlpDNeTDfFFWUdg7Q2
LCla32Wvo8fQtNJPpQt6mvWVhycFO+JWP0Fuswm7TfmsgsyygohpK57qlIlL
YZAuHb9qv00BsOkzxh4/iNreza3KQe240j/pVEAPjfR0sVJ9hTK1HgLjHD9l
zP6u8UHvoMooqasJQZl+QHw3JCHxlt1ynuXmuaUhKCZhvuu5PFTRsZNsWnsn
cg59m0QH+TzJhDUZu0NnsG4tJeEQXLkyD5x5DL1BP03DobJcPwDdlKyKjkJw
9fAAPSG4gYmZNgm11zJxR8/JKEPctx9O/s6pqsvhM28wvM2g2XJRXGtYpmGB
3xhHzrVWNa/s3LiUvIVB9wZCJE8y1xtvZCXsiWZLZ2P8vq+xiYyPLkTeDEWe
VItYys+Qaw1/O3WwF8Sei+0EbVPdD4mGrHylJMcbRT/hIFeXKMqznW5l33wG
wcxK6eDE7oQVSqZ0VP+hViwk7RHUoCOTFu7LFvOz5f0V6e12ttyrRt6AZKw7
so8nE/hgE17BHSolsa7OspZQnTEWZ8ShdfOSnwrU2rydVxbTJNO7j6ZLchw+
FxZYhx9FkJ765drwYf1VJlE8Jwvq4Ll5S5ZfohUoeUfZjcFpgbjzM96fUh/V
oTi+TlR/eHmqffLQmFkiLOgq8SDt2/9rvAcK3uC+YwhTU02PfzNIdcYn+Q6Q
fotJgsbprYIaftU9hbtXSJylr8KBQmd0NOt4YjHvtPfj8Mb8SBXZs1nhxnXs
A/NOGTw3fOHWa6wg2xtAxIZHfI/IUda1K0tr1RymwcDAgyVJk+KusFOVBMcq
fJxNuN0/2av9zbNzWYkdgGrJ8EHnZBaZysm8Lk4e54Edy1LPuxa5zjmv449s
pdLjnvE3Y9MLiwTQ0cvKb00sxu5rkwMaYjEp4pHMZo/OhmNkhxcJ+25HZLCX
9jFtaXUrX2RZPi8fRKjI1PXUBkm1HW60ugI/nUsHf8CY/NPXXgcaPvfmzDzJ
0TwyK0tb0leNmwHpgDnF7NLbCPltqAbBDq7/hBv/LwRXdUaqAzOH4pzwcXA6
sosxR/mrNmIUHeGxV5iW8GbTv8n6x9GBXqrPOT3uJLsGLsS1Rzh9TjaiPuTc
SPoVtE2nttKnnA0btzqLHQNKVQgTN5zHTP9qDv/LFoeiA6HTfJVDw+rNCCNe
OPjGoOYlkDTR5BZ13h4Pi63NRvxx7AlQ6NjXMpYsUyUK7nFCsoG9ON0blKfM
CChH0OCcYqIojNplHufkQAPa14iIvx8NUxaSkKkaM7eJeAzevLEnxmFKsDLQ
TPvh0r6yldU6ZXQRJ9WiomUaiazEAeGme0TNdKiu9lL7Uj9gVCdUIy9Tw4nO
X3KZOTXPE6Xz3p87RTpPxGlIIfgkF2UOfXEb2WFY7UFxkPfDyWcfNczjhrCT
aU92pc2ZtMKmKnYWIKBoJE8Gn1OdTZOzOY8yEPHv0Cqt1YTWUzj6aFbox30p
0MjfbtViXcHSIYdW0xUomFLAuJ03vYzvWmhDwQukwQMpxrsYevsEnGf+f2bW
1XF8KmXNMmUzrIV6gDY44lA4J9K6li+rVw/qeqF4pnpxAvxfY0ow/3RbOdry
nDTs5nmFMur/nRzu3fYPusqJ1WGoRvhU2oI6LwJnHXrLHpKxsq+VSWU/prwk
YJhql/EBO1n3GvicGVV0/W0S0v0tfX3MdrFfgdK7nOJLOz2kOmqUnq+hN/cg
nP8Pno0h41HyS1jWn62X9lhvbY+KJdrfl+Stx1qnFB9xL0PsWATnvIUgPiDG
paKIewivsKeq89C8+MJ4ptLepE+7KHy0aaMlhvc6+WwyHpA67+6GNZ8B9+Py
UY6wzP7U+JXLRN5LGRtWT4G9sAwvTTVywI0IpARoWb3XrfhQtX4wavcZ6ru/
YcYXF8HdrmHZ4Wze/jFcuz6YCXQlBJQ2EaIA8iBg5K1RqkmDbKWyNsfQv/y5
rSpZZyt0vsxByJw5PSfFLodJe7ruaU+Rkh+ccB693+0qTB8sjttuIDqJtT+2
qCOGippq1Sr7xDu0CZJwV8ZZDZ94fyZADMo4XMI8IienXc5TEZgogG1U3dm1
L32G0faCshSf6lDY1L475Kl/CvoZ6yEsP1FMAsHar1nlmmedNsFG17+AV2tV
5qpVqZfKYGqiCa8sL7riNOOmsxbtfbSEYAoS0FCJaPG701wyx8bb6rTOJYso
5f449jHeg3mkD1tYDeCYg3A8jxcs3vxHlhtaAR456caPtQeWNyIcfx2X/z15
7LQbswWQ6PctbKwt7L1z3BUjQQx5+t8ysMkDDw2LXCb7GVtWmLGWbd5kpQQG
0DkKqunmce63NElELr2XT10jqZahCR8cbfhLsGkhfSPuvYCz9BShcIlK+SZM
7K1d89l8H/MXUY270Iao4TfrxYvffV5c1EQ/spss5Eb7hKPgpdpj+3XKGKw/
zlLmooWSkIeC6l4Nl3Y3sJyC0h2+Xk7Z5r7zFYJJ4G74OgMXwofda11lpPfl
orpsYrMRA+qRbMkbLDy2/fP/FPyvcCdSGYdy1Lqtt3YeR4bdXCqi2oaBOs2h
EqFZyh74SkqK3CP3TBHH22y4skTSfRy50l2ssmmibRUwYIydCWikKm8x8FwG
KmsUwYtjqO2nwCzqtStA5CeHSCI/yZKR0M3LCpSj9XpgwEgyubwOSaQnRX29
5lDcV7CtWEd7f6/HXIPTTPfsebbYszbsYmRnuiZuFvKoxsqoFdKlLPao8TxB
nptMyp5ZxdF4MbA4JyWqzP+QYiV9xnzAJp66BJekOoUhvFjeCphgXVnG7sF+
IJICwyGCVG6hVyBhe4FlmxarWDbTGe1Ww5IhyRSKsH8SHPolyHd4UCOxQfy8
SwNvhOnka7CJyL+TeoJG+gb4XVLmgmVybivSE7euKZ8f/i2yiw6S/WTbd2KI
4htljXqwiIIK5Zo0M2tLsOug1mPBHNggkBT6lvnP7nsLXm6MveHqLuWgyDY3
Y0X24ArAIabNBBmhOgTByAOe3qHggZ+0fJZEhr6PJ9TL6sR2H/CPjG7gEHR6
2XudbTHeTAiySlQUT76W0Hee38sQlozUda8Yfhz6hpDYFifXYnOZhzF4UpJT
TiVTNeYkJm/OsYP0wyiVC8wDgv8gAG/YT6I/hIsaeEN2uzZZHaUKS9W+vmZ9
Mr377pJYinqH0Px59FV2fqy0XXVZpCy4re/GKfmGJpI01/uamRhva7W5z3bK
OSFV2B6k2tfAF/xwtyiA6NAyCiKXhcFp/jmUpLGOU2ZMcPWbjYrJYjsqfdBm
yCrr1pp7eQp9Nj7YoE4Dl2izGWoNna02ayJwx/nR55ginPjy5OgjP3OprVNR
1amzHaLiQiUw+fuhrqg5Z9v1u6SNQqYdaVOnZLWl3Z9BSe+IxXwjVQ/aimqf
sWTc3Wp2v8PRzLKwoQF1IwXCo5gfumhy3Ea8gxGsNx/ccIfGD6QLzZ48F7zY
5+dst69Mhty7YScAss7BqEMUoCiagRilMwuGk4pjmQ/F+wIYVEQKywbhbrk+
M0AKedHwxtFslqlcSTxE4/lVzT+ClycTZKXEHkt1xPTQwMfn/bxtL9UejDWS
wezCm1s4TQMoc7TuRXiE450GcNChB/LJS9VABDcuXvv3w7IB+f+iIfXhjHe+
3BqueGwJySDUkXNAro6+DgXwnd2GC9UafpvVYV/6rlXqjBUilCNV3VhpoZ6c
Ii90ZdGv5I7v/g4wKR4jgKy8kTJzeHZ6qXkpk26iG3hMZA3J5+iRRQCiI1Q4
Ir4j9VIFbol38wsOwU/VZ/eWUweFn27gdtzXTr/DnNJ3s5TGvimn2Jz8SbJb
s0dpvxsVBp2rvAw+sF/2zlm2Z2mCHn9aFoDOqiKXWoCwYz3gAi7Gm8AQPlUU
tL9ZCd1jR/lyXAxUYe5ozIqRZe4C2WBldWs4jpJjMLVoRvcZ+sWznt1aREge
LEgR2yEwF9NoY9Tbi2eSuakwFy4Pv0tMhZkIKFmC7ZaF5MviME7CxMHqjnL+
c6QYZJHmRn8u2xyMzkS6LR+DlNo53v7CXNvi/CkoQdFelfKcYJgLO2m3K5mu
CAK+IERqD00XGNefvmrNf2CkuTC/qUaJ4zH1XiBxCqVI+UpcgpMFQNCmrjc0
nXPLaTutnOe2uh//e/wo+68jmqoGZiaEOgKUeU7K/TrtqDG78owepQRSM7EB
1JLIWwPJJounRb+Vy0xbTbepPTqUM7OgyYg3lJxW3mjMXOGD/LEk+bAqBtW4
eo8qK0rZzuYKAotkOTlDws11NZ8LfNw5HZvPt33eL+EKa7zr1UGjNLU6EV8f
GLiUL2iBNCqNIlZmFAkeKJchqLuiIwTtTjKWauSNnHvgCyCz4BZni74fgUjH
zJ+9s/Q4bHIs+bP2DJ0iy50lCL/U9iGBYTVVRZ57dA6CESRGkWYpYGvCcyKm
GLTVhA6MBvM05DMKkzwSmnByU1wIgCo4XGNIj7LZ88t/0dCVd+p735JeJjdu
5qQ2LoEmfqlcReyK8R/tQPMLaeApW2em8o7l4xfW6eaVMWlYIWwmiv5jiD3P
rzHWuwDeOPypJdjChf0y+tlIILjK1BmlPS9/i+qIr9NIRShGIwesrq5jEUMt
5EcMnG80UVBmBv3mEZ9h/mkm7IiCR2SX9MyzpHhYc92f6BBfxO0LSN8ozPpQ
48Eohf0+23Evx4VT2YY+U/hw+a33ux4v68h6vHt14sLtbkqb++Ij14IH6eeR
36Kg/eO6nrkEj/zyingIt/w3SCQiFSGSMhjnyd5U5348kHsjynloc5JC9DNA
fXoQKf5XHukUEP4MaOaP2Lxh3gVvu4AcsqCkght9HJcnmnF8vGhIeCn3CWEJ
U3UtHwO1rbDPvU3VV23gYl6cWAwP2DXIH6x2EEOW9lAfc9dKwjye2ulneoO3
/qPYPeZg/3fYjvGbScPKVfbkVBV/AcIdHnDTvsGe+t++OvnHMRxH3rfZZrGy
DyKtOKae4WZazzN7+pM+3ufrhzsqHLXzKTviE6K4TFPWQTKc3P77VGk3Sn//
LQPlWPRBlZtZr1o30WFSmwwGsgboUpwgxb4/qm0IJ9eO4Ca7NQMOYEbLolHP
R+hbicrMH6snYNufHqIsI2x4QbjB+rKgXPQ0MxmVANXnL4KSh8mkJaNXQK7G
2i9pfQEMD7rMwWPr880vd1XNMERqn6ORxi698+hnUxDjZQHndbR7cxDnJe4M
5DgNnStzEomu+TEi6GoJA4pXhADBQAE/LAteXTXd3Y3PiKoJ3XnA81auZFrM
V2sWG4hslhpRv5M4raCEeJmDP9V7qbk907bDSmUnOS7mgCd+9KJUXK/B+1zE
5gBZtimaK8i3j5IofoJADWtgWyp2ovIDvG3X3EFzkMCG5c0RNycatdckOMcU
+0nqO1hn/4VnBM9Zv7b/nt3HPGjk+qtrnpeMfxyzxp0APPmf2AOtj+bdzVFX
HChBmiDXnZgZKWnQbkCVDt46omJQvpId2hi9kTHu9+QMP7Z194Z+wMCGyYNE
F3RX16EFHanrVtILw9yXmIXCuBZ5heETibi8tzLTLopSWp/PNR58WfPzjI9P
AKJtzMhK4/4FEBgxDm/V9HU5V/Y8755HWxfqa/RwFkHpCWHfYVTmijgnrmOC
0aMNs+zuQjf09eIr55NXJpo0AhzW9/oZ0n2QQOTDQYHKYJDHZnVaeTlP/Kc5
Orp2P/SowhFbQ/WL/TzJbN7oPbkh3qwTvz0NyH8/DwF2/PLllX++EixDofe0
NKD0Q6hfOphoqnbfKGwSE2VWxrSGc8fe1BzZiGtQPhBTTZYa2MKTG/nEVvV8
j2+dduh8KKHt/BBD3s0n2pb6GqxtFtzXY3bQU9WeekC6J/yE9FyJwlqe0G8R
pJjv1GAk6e87exuev6XBPb5r9lEKJReVxbquseQYy7vPY0kQcdnvzvxLj6rl
RPztb5IqI6SzskRhxCLKJ55gHjJj9bG35vqi5KitjGRSQ2J42UiZYtOV5hTM
KoWqcAJTnot9e3nag+CIEK6EaI+393qNRjplykKfnunqI9n9jqgAaV0bwsjz
I/mpZT2NxiZFZMnyAw94PglbWpGnkdZyIUNmrlIzed61Pjovi4Vfp7E2YOc+
tplcS+WIctCm69K/dVcBvC5K7XXF44EKGPYPEVLy1l5aYVPiIs/QSQ9OWQ2d
fvbkH05aud4B1fjJYuqeUgLo9Gy9x/IAJu3Ch1m4xZiKa0rqj/nOimKfJtmR
2gkDftPjwdGrcMWx9o6aDBGF7cYoLjmP11UPIattJcKt+2h59Wam+jkuqUry
4sS5Jiqv0mxQXFJvMsTRH5RzSceBkXsVeBzGED3LW74hQ2xq7ffnaFxU5iES
WJzLnlXkAykoEkMd2cR3LD15G9X2Tr6VWdQjxgbsjLoNkQT2Eiqxt22p9Y0u
OSPCCRKCmhZ2CLA0eUt8gWfvijd+O6/bfM7tCj5KXGNpiOm1obH+Yy0EVLlR
0ZZA6Pgg66p+nw/SYBgwN/knJZjF2dXDKjdw+F1THmJ02ajr8V3DZY7aBAZX
uUEDnD9vOJHKxdfmYB4UkkUC7p4BL0ptH+IXga9ZzH1Bjn3YJbUzhUP8Fyqy
Ic+gs2MEUCMcMHW90UDWoL+fFySw2X8Pk2CtdVJLQw/GV5eJb8/prwZjDGrb
GMqCijYKizUsSzb6Wnv3HeHQ08vH4dKYiyYQVyTBOAoJrm1ZJCRYZIEZjv+D
tXZVGaFuhIHjNee6scYnqAQ4flaEFRZnuvx/cRP6qwQ9XwWEbVXTfXp3bMeo
oZdwAOMprARgBolQLlFqtpk9mvC0rmvO49dWrOsxpTAx/atUjHJ6iWCUFzmK
OOJrUqUxsE4LFs3iL87WfT7aWCx8Em+ZYuukxGSiqkTvv3RHmyapBmgvhs4Z
xDGh358aXxlhYanN9kikNRQ/ipzNxUS3dAf8u/IZQMOUMpxHsSzgAxkW7+sr
Ip6X/yz7KWX78ynO0cpHIf1tLfsO5SkfnNq4CBDwpnfaAKTSg5AQbuIWPgex
6OAsOXPYItki1erah8PdJ2+Q8EQL5CRql+7v3hyDgXaArX+yCUVr+r5KCU7m
Ywa0jC4wejJHEP/o0gL9giZ2OgQ1QoEsKQ3KlZMVcTWbcorCZs9OfxsnvzWI
SCTyhlil2DUnYJP5bs7bN8yEfJHFJjasF5kDEbFqgOyiinYii6HCidSH/xSt
ggTZg4UOxoVKKoDqkSXu6tVyVhW9ygpjdJZVegZzoCgIoCmyza/FyRlUA1RP
85LGSYkdpzpeviTk3hoZb4aD71nlrNZh32iLKu5/9Pb/Od9254fdfBtNbAg4
k9c0pMhm8KGXSYv/m4Erhtj2m6C/QMwwwCXy/9TM82qVp9H4ZPcSZZB0atje
Rre/EPGa1eETjo5OaxQjf3CMEJLUNXnhCFwOxUQ9X4tZw0Oxn27qEO8D6cLZ
vpuY2TFcQpx40QM2UGr7//0kaRQ7yrImYchHX47bF2LxHJzbIZTiOGc6yuoq
TPISDt73OpXNtAz6ROyo2E23D1EhUpybft/oC4Eq+HYLgGkaQIgHohkh97Kn
PKGWOyjLXyYjxHBfXCUstr6mZoV9fcfS5vPrzH8tspRVBWIMUOWDI6kdLbUM
X/+ajTqmuRE/HdoYmyZSDQmqK0pIqMLRusEP65cTxS+Q1mDkIkwV52Dws6SW
gDMktHT7mLD2AMSFoyEpVtY5BBqzXCSGAUMiiHQx7jL5SjHeMofNv97LJpSf
4sgICzwFAO1jJbSFqyBrSDathomXKWwFe6QTois+IVdg1grwjJGKJSXWXW2u
AZposDQb9PD3BSAfXnansjEg1Yd7CKTrTmOYShcZ/Zq6+2muH+054kMTi8ZV
UJn11vOX+MgWudfPT3qrvtx4vmjYAEEsXrIcPWeZZdIBR2eiWcpP9BSKR4Es
9IBUirzEaLb5C01ZAYzuIK+y8WQjaOhQzI1JD1sj46AGSidH+CjJHVCDkSD/
heWDwGis58X4H5Vi0TZHcBdtU6SEo+WL4K5e8Bm2rre4Qvq3VLUTH99tSk77
Q9ygXmNdD0n+CimYK2Ws3XFGCREDVJnzAbKqT6L0Va6xV3Tm54EIHjhoTvzV
uRt0sD4m2RI+tDin5s8Ax404AmRZc13AnU0QNjPEWulfVEtZtPgZNt826PjP
/+cb0duqpIOmXesaxbnBUeaVaGU/W6fCitEe5M2mVagH4JBEMk3djjWiyHB8
Sp8xu1lAFWll/RQFN8OTeqU6QFSvqeU5R/nPfdRG4hCdDaWE/9PN5n894PBd
lxVoqlT6Ht57Asng0l5H2n6KNMiHPQjPiEpvccUq5hVycfXVpIpJqasLb8B1
3lShUvxF6duYKBknVJozOGl7+HoyYl2Uko152owGJTdoOUVga+e/Ft8s+WCI
oY85gFRnHPQ41g31NJydDLOPVbCUnWxfK0Loy2iUj9Ft25EkzMnOPlZHmRYV
fIClrKQ0GsCvDZ0gxQfDJm/lKSa3dvIR+q9gw+XKc5a72FSzM4F4IUyUqMG3
4laPiLZwTOjRn91ukbWw6SE94Vi8wun5Zs6eh00qWfo6qA7KyAEV8YwojwYY
eK281iycvNndvtql3s9VHsAQRLO00Cm8xUb/SbzPTm+TEQW6hxutbvn84E8f
Q46MlEabQvN4HnEB0ZRmm9Df27VVt6Y08DfC2JYleuJQWyODbEIc8OVDAcEq
Jv4r3j0Rcye+7WZHCscQVAT5ILnJ5bTr8TGTXzEqUvsQLeCN4x1bClPSnaRo
q3VoN+i5+NE7AdaqgaUBm/tAexrlOykQ8OjLbgl/wQqG+hkB4tMC440swz+Y
jtp9us2ktqemHAnpA8DRicQdzezKVW8TWC1M1HrUaMPWkgh4Kt5x+apEcvUX
C4Xxeud4I0iGbnW6y2LJRZo6sB8zh3VBNKCWTc3J3dO1wtjBypsx2NEfykr4
dtJLhT8LxC70g7l6CsNgQgauLf/59bD6NqwJ3uqBdeaTKexT1/B/QTjfRATt
8GPBtTIUF4HFPVdGmtL9AMgBOP6Q3m+UR/0WpqjfqHY/G4wh0ZgbucAaDwoR
v7bOLg4UCAdfv2C4UxhkblMRwmnV7y6g9/kZCzb8gQxCKPeoF/DdLSwnUwL1
v7TZV3t9Zu81MUyB7ns1a3TRNE4HzgzfADQ/3Q5OtfEwDhHGODBzFB3R7KPR
WX399aKaAYF5eeEat+4SpwKxM6uQqD+wy/iPGQntxEIdCE5MwqVKkqKioMiy
Sn3/Glk4DJto9I0LKaecQ+PY69N95qAs+6MWD8uLfpCOflOGYXpjVv5yEruA
bsR6JL1zN1JUNqd0zuSg0kIodxxLXpPXojq9Np3PDiCTxJR77dcZ75QbU5Y6
OxzfGEjSZOjUSkOCohT8594nGFDrRgEmxl5u7vgFtQ6iwKPDckxyibTXdrzk
0LQC9B4stGo0d+pydOM7HZAA6UZOVDUNXaZGrojuwyWM0oTeFT7tSBMW/R9k
8U4DQILNuv3z65DxUPkUnE2bHKLcwaSBi6OZ4rqSHpbLOjz+yvs64uStVLWu
YtLsKqovQHsClEZp3Gxj7hLWaice7C7r57HiNDgHFUHdpQG/KfszxpsP7VET
iAAPYHMneFEFIoa3iu2prnBl88+kWt/aJYHUqIWdrcZLGsFPOQ7mz+n/+gfs
znA1mfUk7gqf0RDaoa3JGo430yC/8sts++CplJhwf1JVLBnrzQ56hM4eBZY4
dlkseVXLpxJk9Yyu7IB6toqxHaFwLx12jFbPIbpQLGz+F0eTo4d2BQgFDj96
U60BUvqH6cvP/X194slqBuEdAoZVoKE6hqtrDw9lJOOTBGCX+umycEl+5BAX
U1rXfRmUAuGIUStoBe4tSFRl0kh1c/iMZxjmO/1QZlPF9V627HlUhd3+gKPj
QbTgI3+pvbflbX7PnPQcf4k8CeUWBwD85tikMT5O5/pKVtZlxiMyZ5kwgt8U
4ftFVb1JJswKP7rbEqNjq1Xuh0cEWz7OecKG3hJ+DOxFuzhs+QjUoqRWw5Gr
nqUTCWLMgm4XovagOsqNroN1pLMxp80b9KybjTM+ciWgAvkO7wiQAfP2LQzl
CyJBOABvKH4kQqk5w1qI/GFrMfUDFzJl3lFAhEJIFGAcovkyl1x+yHJNtI3H
hwiBgC2w7wpTPl4vDZFt0WC4ALxA9D/PFNCNkjKRkFPzEHfQURlBJvTBh2Jk
tLxzLic7RysnZdk4I1oSLK+bd7z0yG33wt9qRlYVruCq5A3amORHRXcKsPng
h78+SU8xsOVVNz4A+eGCCDUp4cU1ZEGvFN5vXkg/Hi/amYICptRzuyxC58qe
oPkQBWC4JFAyIhf665ZM/D8/u0KNzh7vJyAN5Xwv1F5cfIB6xwncWXrPLDdJ
bUNLrBRopMj/66uTCOk8bEamCY8mQP4hFVA1ZhmhMUnJ8pHjpjp2U9U6txDG
EXJUrDcn0EysoAmq19L/mli3g6GHgtaexG+O+mR95rKxJZtJrRZ7XL3ZKTuu
ReUvpi3vupPI55LsbMk344RdL2bjl5m34L/knVmftXorBbHR/jiGG48f3mWS
bFPFGRVK1/cgCPLKgjUeXVBmyZLdbXi6FPyo8r7qQDDCsnFpS/oy/LYl7lXT
77lZ2H74XHxDgO2arMqQVukU0XFTCn7xSosSvqYA5YfpaMBx4fpLpr8CWQgw
HYazkZQ4Bc0ZrExUAgmSefPDXPvA8rigClXAa4UTNp4J2t+dQOQX0dfTZyYY
5oXegq1tFpT+culiIvt7dHwYmrHhN/tyfhhcymTlTV90Mrv+LP2Hg6ivwSdz
Dxmg4lj+T7F6oh2nIQM0QwCE+2PJZB/LiD6XAbyXMknadJOxkqJ9SSSCdFMn
y9BPFZ/5KD6ZaxDggit63XGtFRuNuHlIgTvpNwNIDmN5EEQHsblrns5Aei59
ku3B+baxX4fK0S1YwBw73uR658Y9+2lfXm8goqMHuPlYIgYMX5wGTf/8UJ4h
f0jfxCE6dGHdNp6VRZp6oa9cN75i5lRSjZ6rR997W1HzArS9rLiRbplJt1yZ
aaxogm35jv1p2LArFr50Va/STnIjBCGfh5XxqInyVf0qkRqFEFhQRXVz02Uc
Nt1JPIy2ilo/ydNDoRfwLpZTLcJoZ4Z18pwI4owKChzUtyNJDQGi/UfvxhZk
f/K9jUS44C2VVSC1OtKldRm4e20rhnNDPyxNm4SZM64u5p3mQDsFBglO+Qpm
s4qCKrldt2hJtJXhGG+9pFUHiFbMYLPH87qJ9FC4Pg6hP06Duvvw2qi9G+Lq
uoytn6Ex9ef8ykXwthFj5Woj+BfMdO7Uv0xOHt4pnSgpc2oIKC3RuyYsNPQ3
9nLG7SxCw+cwQFTyyz1p196d55CMqkQ+iXTY/fMoCLhFxyg1pXn7DGhtM0Dh
wxiwVPkgmctqZAbCyOXDrgQwm0h3gJ7C0AiVN0plAUqLMYh9H+uF4owG+eUJ
2eFRmIwq7RYFClyqEP3RFFfhb3xE/oBWhe4T3kTtp5rl4VTQc6DGi2H0jw8q
JU0I/PEHvQc7aDn1zcfR7lqWTNcPRsds66GBHbuY/QmjqBlfsT1Dna8LmL+P
rISdDS2wBoCzvJEF6FYH5oye8lZinsNx2qBFOd3Jcx7gwZq3CNjqzCebwnoD
D03KqG9Xon5oD9PpD2MlgGMO2ifpnjN6AbUKvERe9XvbTjB+4ZSOPI664/mm
yGAE1yRwtx3OEplpEa09o3Yk64Jbf6/PurQPqWlBpS8qbr1Uf6k7sH8GYrVZ
KlynqjyZU6MuStPUQ7oSBLATK6uczUuV5oy//roOPIgz2FaB9c+4SAt/SZUt
oCm2+4F8rak9tO9Yl09mEQSYeUoVEoLkwbUx9oD3ZbjpoRiNvDIhhcFZVWZY
RzLfIQHm9KRjpTyrxulA6O4vcPK2tc79gX9rHhgBQYjRUu2xMO4+ID6yhRb8
J/lhYKMeoxpt1XrmMxC/f5C/iIJre45If/zjjDxEfR4YI7ZJvQTAzzaPdD18
8JhWD7SewYLXnPKVj8G6W4s39lpeyJ1qdYGNcE27nblLQlbrW8oNSKc2238c
GH8ouSQHXWNjEn6wNfhE3YUGR/6tJif+7rqeIKveNX3d+FUqSPPz+swm+wlx
BschAlrTvjElaXk07OixeGs1nQL01F8G7TzNPnXGLQVOlosMeSfu9yWwo5Pf
a7EBp9DrPTPWZhzLFzFX+r/dQvD0sgQpXQQEoYKIiJfTUnOC3dsua25353Kb
io8nIWTdmwQriInRnSEcMXT7w/8pv/JPkUxYqNJKIZS4bGUuFLG79O182Zm2
ad+ukIeKBF54ncqmepts0+QDY/jI2wPRvEYSPMS/mSKaLNGojNYt2jmD1llK
qvZllJTgeEnI3q2QowSf8jqL4h6wQbsBzTCt/swe41G1dBX6ulfmBBco8Z6Y
hXVKxx+Z7nDfblZPafYoh3GUemoLQcJFkNNi5TtP22i2OxJVkzsmektsWAx5
NfNOJBT4xtV+/rpqOgzNr0Rd3lvtAbTQKn6zteLkv/BQChZgHT+frJyXBeEm
+VYA5B5ON610iKQDocnxO10rQdYHI3qYnAYok+2I38qYANDt0J6ADv60pSsO
lH+ZFb3+CfIpyFYQAUs31TPk4eIviKvOT6A2+Ki6E15CZKtHRjyWPiHDq2rh
HC4szkoWNXaqR4wM8g/Bv7cVy5C6gCxQLnjdhFvzy3b4EUJYKwP1eFD3han0
izbn4WBtRgFY2T3vYlRXz2MjXxBAzi8pdO2R3kubOad+uglIRArm00yTeVuG
AVC1Sx7MScX7QalmKhu7tuO1pES60iMDotQWE9xrlKAcw5wV1ul58YVNwL4P
esTdnWANpngs60oPI4qPBkmgKdmC4ep+VKJH23hEgJyQQajGeOUAYm4hZgDe
JDsXpgyBSEScdntXcChZjlnuQjtQHdqV5gmOvh+bLZCZ/kmQwKEugpvhTX92
t+pkX2hb+9yJUMan9ZpUO88ZRBYLVutGTjYL3MLfkEV3PEaEAetgOiyMkwOO
cOUIZ5aWaKgH8chQqMDQ3ltIgdGQ40hoXrecrjQGaYoYbEuelGa8MuhfhrfN
jDOL3NkCTzZozGIlGYCjy6kouLDBIw9GJBB2f0hotaVoZf5a8HQfNPXLLnau
q38uGk4Ga1XeSrMei+d/WJr6Z+tInXAH93ZViswU6nDjmzL6RSUZLkAlnWD3
zjeblNi3k/FZGaIY0VuL39XroNqTVYLJqDianAafbl+vEqibDImpnbOgqm8c
o47zu7fjCe87qSK+1lIBz9Yq1B+Gm4VgjfJx+A56IQv0+KpKuMztt6MOyY4D
kx6B9ECLRb7UuYyWOVFgVPQQnCQxs6ZsmjUiHX6Hd2KBDYJDsWI2kKBzfpFn
eCnOHyzPfps1CHPAHhSYvJmMW1nrK1J8KqzlOVoRjJQLza0taCKr9+kgDaZ1
FTOkMeYU8VOBKsnsp0HxN6t4VRj3r4WLbqeNFstTMPQ9ZQE/SlmnVuxE2XNY
mKHbXyRppC7+9cIlVCmI6MjUYlpcuyV3wGFljGc93+rNrEDyK8QPBxVdHC6f
vpbellhZtkH9YrLeuK4c0qIk0EkD0ZnXtATeGbrOE+MvtjQuYgI+bCmR/54N
KbeBm2MJXoShRMiAT93v3Ktc4WC1ffLWPE4tPKilNAZHx+b2cddwcv6kV80p
0lOb0bNSmSvoTuU2O9aM0+MKDXjhu702LdMN+39yKGHgoRFppJ1XtdQhQ56B
ocwZ9nX/FyIptAv+h0JlHNUrQC7fJCCsXB1PCjHcY2srN1bqnweXHzvg4P+8
wUv2uJTatBGd3gnOC4X5i+MQato5xw+FpdXB4CS8kkzdJqvhg1dUb+kLK7ee
vNDBGsmC7g6IeGaiE+npo6OqdHsTzwB6TTwvEDEAUgZzFMpaziUykDBGxXFp
6jOC5Xt05oJ2Tn1FAvSrLxxIbMhxanRPkOnH8zlNxPKDCUPx7ooGtpYe2HWH
cAPJ/A067d5oR9R68DkEf1uxWJSc+tE80bYLyxXmUm2Ay4E7vMcN+beIh7uC
0gXqEqV2Eaz5mwMQQp5+DiK46B7TIfZgO39RfjEpSyTE/UcygK9AUHQATufA
2nksIl8E4IS60Ny33AowFIRLjxrJZn6fE/YYNJdvbmovq7aOc2nDpZoXLc9U
nSZrp6qmBEH7nBzO1JPnbHo3m9ftuisYT30wV8ZvxEbq677ePsDJzXamEOeL
e+Mae9FiRYO9lV5hevKDPohW2+rc8OqNXmGTD0j2v4sKl+J5eJ9YIdsuBDVA
t0OZr6CDCF6Hww9gljUHnwq9pMPtdq/LMJlpfF31gbwv8ydYNaW71ziLbv0J
wpDRxOxxvhCQ5TfckQCf7hgvMeyeiugfMe4Su+M692NSPGT2Fv39GlpHwjo/
hkSdIY7jLGTc+PQzmj+44e0wF4OxOhXyft4l1YHLjyJVTSU1CfgNF5ENBf61
7alOm4TFXeExA720Qq4TwTltMrwmL1FqdZdwebr07IF7vz79kBZLpIfVRw2k
H8WLJmugh9hpjWTG70qpSp89LlvDYarGKyeUpMUZS4KYfRzHGi6nmhwYKV8g
W/Mg/hCGmRoZEKp9h7dHF1ZQ/I9u4IDWsCsz33YWSUgV+0lTRjBH+HWXjwTk
93EErYxWANyv4fscA1oriV60Q3Ckxb2a7i/pqOxvRbS4SQIUf9te8yJxxQfr
aRuOCXGS3L2jGt+6Nna+M/Iizdz1EkIavpJK9jeLtZ++yKaBh4oDi0/BEnre
tzF0shYEfLtFgKHdD/QNpcTUEvoTwU8/CEsy0+0EHdp56kkzYLVos9p6tsRL
8f5XckcMRuu8FdxNVgrIwqnjmkGMZtpnhzlF9QudYIJTXxEdoOzA1AoB/t/+
87wE+9e84oYri1Tnc4IaBRmjWml75LRfPI0GjQZa0AUH8h5RmnpmTK0cWxSK
3xMOUeseOJBx+ARb6CdZ97XmoDodHJBiY2Q7WcYkMw600its5jPsacvpMFQc
2lYzJoluo6C6XYj/QOSG/oZql7zkB6Zl6ZVP18VrCGUf3qPKmVehBjvHoIM3
5EoxXrLzXsgljw7oYH1XbT0xnphvk3onjbfNdjgewp6GgpTX2vgszO28PNK9
Y5nCJ+FETim7iIbiRwho0QZRd/TTNUaTtD7WmYVqTwA5qYwJaycXrVWXD9GW
KRBJFvw44ckM34nyImTtULP3NjL1QXOATuHLFnQkbk4hGkJCEBzPeJVXZ3Rc
yY+N7V/V0h/lE3w3ONwzdxX1bSLLsqrNkuAC03vms0FQXUKMEp/QQH77Wcy8
uj45A1+JIFsLX6Ws7ylT504hR/8RuOMIbfqxX8i5g1SHv+5V0++dI7PbzHFx
BKmUd2RET3fCNPWlu9PPMB98vcsG4+chm+PktTaQgUv+Q0WiPc1CAr8dG5/b
nMKC9pSxqaR/dzNDaJQ1IkyEWZRmVuOkXYACpsHmYRgtI6m/vbqK0L3U2tjW
7G0OC0tmLrE0Kad8+XKbfiJXQS3vWY9oBUb2Fbl0KuJBtY7rnI1QHyrPJBlg
pvz23a+Vu0VArgWt0zXQqJCq/ftHkwQxEUrG6HlmGTVNeWyfTZiVi/zMCMBt
K8XRURfkX/aSFg/136AijMaZnMYRcdvz1DgfEJvYPqXewBllwjFdtTAYPYtc
DdDeAZwWhY3yewukIPVlg8X+jZT5L4J6D5/vGNFgQJxhIOgAOl+0I1J7ns8p
8PJtajLEhwr4p2cnzs2uwbpVLbsIBPEtrl8ThnJ0aZovgs3eV4jJ0pxvqkZq
9AaBEj07hhkJ+d5c2p2v9TEfL2BpD3HnSbHCC+nX3x5sq0ULJronOUPDnK8g
iTQATbjpP0nWpcJGAbekVwFT7raZU84NCsQ11TNUnqGQpUTJjpg6zt/aBwfe
AfNW05uAjPuJYPVsNM7t1m1exKUeuMzP/I7LEE8gm+22gdy0TB6rkAtjkAQd
d7725SG4hYBG9UcTF0etOMMlwhUF72SY/1eXmHL3Jp2Dxw5Uf78oYO+x+ISr
Dk/grmkf0ugGr/kj2Ly9wdLq72czFKaInu/pqVeUKjW1V3CNKNznEOmc1OsK
p2jcsU5qeYPva5U90fyoP2+B1Uht0HCmghMteExuvnmA2BupM4c1uNpPJ7Vn
DXlKUXceKh+7M7+rG3mpXEaXjMMl0Zc8C+OPoa0c65GwUZY98MwwlZmYBVcj
TApT5cs02cSqczoxEzBQLODhTfRph5kSqwLQF/v5xjUx+50953QSU6H/7GBJ
RAeq/L6oLMqdwZNafMeSrld+BD16FGnAApiW7LHUhlnx4LKConHhV1jP4N0e
v6ZSTcQF2TGAAevGJP1hq2MRdGk/ap3rgvaIfYTsqwq3cfpjMgDsGN4Pi8KI
km0o8+SFF1cSHokm21XYEzjJUW17XRf0DpnIdXsnm/ejz64/1xp1fOHpswxY
esng7wfgMI4x62WPJ2ilGwxKqHO8GwChy3uYpP7CCg+7OEvjK5o95p26tMs0
Iclm4JFG2I4NFYPl+UJ1MxCwa4dKMhWdc9zhRbT5hbx/P4IqS/Gx+5xbAOlk
8r0bR3jiY6eGdIOEX8/kZyPxPurySRxv9SB0WKkdZTOVznTNkx/LbyjAH2br
6ho5IJCzvwqADZboZ/t48t8qe1q6cgiVv2gTopO1MszFayvhdgPsVsOxAc7n
gGbMEFYmm6whA8r6btoyYsOaNUxg4JP4Pvn8/K3bw13cuq0MxMQH9aBrQqHQ
F9Ycc2IYXdbABBk9A0IiscmLfGVf6l/DHh6eELAfReCbnjDT42WUGqlI0Qbd
npYOwzfjHAnBljhcJc/kvOtFV/MX6RqPIFb671xzqZaCMCjux5fQPA/YbiQx
gaHW5d3eY5Rgm0tIl/b2yxDN23hEbhX8RjHmaAgeIkiauOGsenNtVxhq9IYd
J4k0FN5nuqgArrRGVAxaMTNnDcwYgT9OHtzU5/ZgZQLOgmaJOaAaWjoDFHHZ
j5gKmLzdarIbidNNZwZr9NbrgaDNdz09Slm7/WPzDG5e3sbSCYqW45G4/Tak
THEGusB1n2E0sIahCLc4cs7LbqSNv1u/4+Em9V9cOh0SicP6U/VVNlMWLav9
52HqxHRSKkyHPW6x927w3/TahuQhkrojJB2Sy6evNnYmIWJPBaaGDtclvAmH
4TpORiibTwwwiBqs2ZdR1UMFUHBMvAwG4P2qh2CJLyr3r4YwOtKBQ/ZrHmgi
bmON9YK6sIDralo++UUoOLMy1m+pXDpWD8dG3j6LkbgulWd2Nrmi5Uf7FF+X
RkJBqiuEl0jKq6KpKmgMPGapHs4u66HbmQuWoRQ9P3SL2fCRo86b7joAEiSV
Xvs3ZiQxY5fxVu/Scbf7IOCrWSihnTo3x7WpWhgxb0p42zRJ+yvRlbKyb/LX
jFGskgqTK8iYWW9BcdRS79VpEmYLMjkUmi+ArON+u0goFwAfZL/YtTTCRWQz
bsKzYr1VTQJu9ecnQ72wn6X7aNu5aO8F6LRUVECrJo6yz+GU94cAOyp+Geqx
iBOnQymUcQDn70WBKfoo5MONMnK553Pv+OJYaQq0zN/FjgViNv2mnG/IJ4UD
zMpv5LKJJTzP01lQE80tWLQQKe958DeLfILcfkttQIYFE8KVBGk3irQS01VV
TwH4VFNj9M/md8SCzezgPv99g81ZCw/5/KCuXdowjVCpiQdsTQ9ZMUllQx0e
4sj0hD8tbZl6EhShXv2dxaA+/XhoyiLt2knGA5weXXAfASzDYSNDxiKrKF2r
gED06fcKD4LOOHHTbYYouRv8YZxL1Cuadj0FD++R7q7JC1WfkmI4Qi71wyvu
6BZb+TCEmgGYk2/lub/TvoJbAmsm/yCAAtcTCscOjNpUpDV3Q8zYgICuMI9k
yutDvOHHk5d8yu54bErBvO4kYUVIQeMv0mFQ5p3hgM/7PrMogtx6/425lIuh
muR28Y/zBTNBJzgdtFYg68YVaYi/yIXiAs2x5jlwSzO/am9hOT37K+oRUkSk
FTpYp/CaA9A/TwW0y1ikS/MO1KBNcMmXffMJhv4v5qbUNeWDkDqzutjB9kRf
+5fk51P22oTYvo6oiCLa5G6A8ZRqSRNUshUZK0tSluuwwBDIFc7wiyrCGrNt
B0gwXMNZ+ppO69PiJjXfBZ0Bi8kUWtTu17udN6ewqpuG4+njEk+dP0aJO4Lv
1HmCw0PGGGmLtnzssmWQiAlpscGYO+ZVgxY2jdteY52dNv4S8W93a9gTn0UR
n2EZ4QVkgJTWxnYUZkdqY3ZPvAYtap6SACc1W+oEYbRsY+k0Mkbwh1oVDokt
+TtDQk07lE9vXzqvArNoHY4NoAQCHt+CQ7TPp9vH/EP93IuxlP7rZU1IsZJ/
MTDofvchL2aZrw5NcEPj/i6tDIAjNN+Jh7dEoxz+BqSY7yCIbB5jAZEj4yie
MGph4FLTItxc6OvLPW+qrJva3wvaCfunEszn+r+XYbW+xDyBXm2nZ/xVgNro
LksosDbX5xJbS80ZPKcRQO7/1gjLyIh6gBslt+Ha44vxtvxod/mUyVWt6boC
HOX7a5wQGCUUEDJiXTC9JSjkI+yg/h0I8HCXz0jsdmti7hw56BTKVTQImavI
2lRJs3qL4doVg8lhsdXLfyML89mePCUWxnVHurLrf4PTS+Kwe0oS1ykcfcCR
0iOO32IC1YgAvmSxoMcEYZLMxVOm98YFoApbb5EUiou2SQRuuegDcpSw+9rp
Fyk8e2ODkTAlNSzqOauLBbaUfswVK9f6rzIuUO3TLVHVT/+IZvuICDjv9so7
qrs95TCa8seJ2AI4iCSymgMOz6MIC5BnbYKzI/3C26GKC4NK69/8iaXpQkg1
IXac/XQvXfeTVUj+STIH+nLx1Enggbdnf1dBJ9TNrzQEI+Il5XeIdN/tCJkJ
mosR7BJsOa6qDuJSGl+9wy70z+g1nJUGpRKS65q0jWw2rHDGq+3joj9j5sOL
TFteqrVuVDoN91QUw+gPMiLBaXJbdLXw04gjAlsdWMNdo8YmTmyuTVd7UGrV
LPfRz2rPAaYTGsG+FM3F6jRk7BhXC609widkoq1OlC2mE33tBn5C8MFyEQZw
btqxuqkFtWxhYrl0t+idFxsw5hOMAUZZU4LCKKaABs1q28BvabWzgxqgfld/
kaPLIT6hSHKi/pWau7I+JNLEl2EJRDjXaGpcj64Fb1CNsOBWLtKKp2IkkT7n
r10SEno3k4zVnoJSruzLTMZLI30Bvlti2RHJHZeu+1Xo+JrHxVUYoDjIx1dZ
vrkbP5AbEGhrl6hfhbic+zgheUkiRLe+IRA/zwnzTUVdPsfenv8k9eRAK6+m
F1Mghg4omSnC0n9uxWG4gMtp7TW03yIeDMhDumDIBEm4XDNGtKE3GHJnsA2E
myNvvpbNONeYORJN6B2jCV8uX6les/hsgjX6iU7DjLqRUgBHC+Ymsk8iR5wu
3+sdWN1rCrGApBdJBN8dPm/wp5p+Zsn0VfLniH16Zl8iGbYbQOb921Yw/eI5
Fyvm88qszuJiZkiGc5Hm1gtmMyzQ+DEAtF2sP6IXdeugshz155rSUzApVDWI
91dcPzGNyh885KrKSUoL5+1tDj7NjcanPL8jRexENA+k6YrNyvCkI1vy9QIv
oRV2Im1/RnsEZP1qDBL1ZfLXKD4u6HLOPr1a/emPXgiefltHogyIOjc/j0Hy
AzX9PHbvx3mAq4BYT/YLmChl3a1SSQJV58AeIAsjxZYwbfPrpB/ezpK8Lv4K
RNLVWgGADsMy1xp7XlKDPq+bhxZqdbVyJiMFxapb3COu984qpC6t/4IiHLhv
BMtSAt0kwtZL6VpiyLUxOik2FJ6BnZaOmEf+U4SMIvvg7uxL4er4Rvk2DbcA
Rq8VDnwfywnjsWfPq3LEQXqSmzSxlzJtI/RtgkUBdhJkh+s64Iy8eVuEy1Wr
CiNAuJoJt06zbT92Sy2nI2/ZFNgvqlBoj+F1cYsHXD0A1lAdyVDYxigKHXmB
vA1wuk//A6TQs5R+qCaF6Ib+ovCO1X/Tm7g6pLn7j9oHCPw2R2CqBymowPpM
8CYgeuBozzweAr9HbX8JzbbGSI3AlX6G1dE0D2LzSr5Qcb2YiZQNBPg/xG2h
yHNju+0c1XN/CypGnD1jZZ+LvwxybgKwdeBTzvb3TbBzdUa3XfEN6mvnRGV9
2uXvU47kW2saFJgAAYOPUmWlX5GqjisIp60DdorhWJLDTX7BecsN1OXTxOF8
okFU57ykAem1AZpUMaaD+P/urbwMESbclJ8dXaXIxry7+AM73zb0AjhMeJur
mHMB4eTIwyvx1Yl8L/2AKwuaMLp3kjwrCnTi7vYTOvmShVDK6gzN7KCATxgO
jQtj3DVymtQ14DYWAu7G+mkwApZ9eLtU0w7FmaibWvICfOPBSPkIqug0yc+d
Eej8+uwU6As0tqJ4Cy5l6w1i8gUZd7FZzSG94wzWvdcfY5Kw0vLFMMrVG+jV
VtJxj6YdxFZip7b71Zum8Rw0sK6r2gXxmWTssMC20HXddav7ENDh5QDFmNIu
F86JPKdxh1ZojuEw7xL5nm8pIDcI+ZXiKltTq2Xhn77lJUCxDhLGbsNpoe1Q
kRU5+yo4UH9yLdqSdBNJdUHxsgdX4xma6vDynr1LZ2hA42mE9D1KbbwvtZpU
jHLB6EMoYf5fetCA8BSp6Al9wprJamQlQofFzQk8xbcAj621ghHvm6t4ISVH
49UUQnwBjpFkkJH9g2yZHdZzgQ5kRGl3G+kneGbKpNEw0IRFyU4a6L8sIjo3
pJYhfQB0+Y5OvO6pgR2oAyhpr2IPnBo+akBXlvryBQWVSYeaw9+9nj4IPzrE
7PtAxpcJ3OrucLCFqjJENIMbR/MOm8N1FWWw9r5/OIAg1B+JFS15yx9Tf90+
38z6m5GXOvfKs4n7jEaj5/V/MdNhX8l59r4PbLcPO8f3GROwivSRRv3jVWkI
dA0s8hvjxTKGsd7zm9J0fPbZUFkA230NXJ6R3VJCe8jixi644CILQmixhEnu
4CRNDDnb+r08HINjlMwsQsaDtfJWKTbzeynPTu5UytQNSFIVtpcfyk89jMGs
bejs+mIEx/Khckb+TLMtJrEAZcgshDXwK4EuB480Xm8zT5tkyHKgE2BWBXPX
eSea8cf17Sm5ka9RzUdkdoFweRa+/OB7enunwO2fmxth+ELmSDOdxxX/tKfx
G4NNxTaQHCP2J34hvEW0UROHGeNoHITM2ILdwbKvo8EANHGHnylcxIKNUpFp
+a+bViNlm3Yn2iV06pCCUEqrQ3XZAjaaqlXUEEwGiVQtA4iS1S5U3ec6odYT
4KhHXmk7ogmTePgdOeM2hppBHBVNsLRdOLNFgtj4Ivs59mmGoHg4nbMwz9Wm
7W9Eem1QoX2QUc9LgcxcOw2z4MGT+8AEymzSQK5FZMzRYog5mbwNvHxv9Pbp
Ox3SOBET9sCBXq7Q0Vu3fQm7J2XQ0mua52TInl/+Hxn2EReJPSAyfAJo78M5
noj1UuKbIrf0tvTDey63x4f0mGQgQzhyXEXwtxjtP0KeHkeMUcmDDzf5z1oj
5awL/DeVnXI7RqswwH/CPBdtST624+ZzkX9+qcoA0SJuuiHAtWO24ytMzpFP
pT8nFTXu1sIHonPYCNXxZ9rM3tp6KK9EHGUOtWxr0tWFwPAvTywYTUTB0hcG
vBxmEld4KibYzulsKevFPfmliesixhn92rwtDaK4Ipp0r6+PZPz1pZfs8V2G
PVyEPMF58U9YnP1G6voGl2BZd8kTL9U5pV0LC3iS0EbLCwlQYAHsTmCob9lM
FUrj1xkujZgMVwSPHk8Bl9IyS/1q90K3ezr3bcS7puyjPrr9DoJ5ZHdatlSA
F9X9ybeb2MSsi1a0RcGUL0VKyoAvuQ+QTVdB5EojNDqZh8IylHz1NMW9SHiO
88pr+8akZ6d/QroTAuUF/aemEIDk/OPb8n9H2GGWpjtTaDKY2pdnB6HVmmMj
OO+08qh4utF+2FOu8uIPh+kJFVDUyFekiLZ9ish8ZJ8+v+VOVwpNE3ovDdVZ
v/uOumOZvBi8jAc2+LJ2XGw1WWk82/08iaWKawcWUEpuDtmugD2yVw7Uzrt7
HTeZvnwHOWRMNQ3NkhAMDBFMfWpSeAudqcBjiVA3EnKPUJngfherid2lji9r
6HbELb4rcNSRdOPOD6qR5n718jRr5VogvsI+7CNKCzO49l9LnJNJnfvGtIFW
b6p6mz1jmiNOZgBWTAJ8K8BuXAcUmyD5vJRjPwUCsyuvKq5Y59eij9pkdjCT
RgL4WtAyWM+UrA6TnF3wq8HcL4HJ61lNQnFSGuHdWbTGyntxFC1zQgxlwKsY
4lzHWdRV/pkGue+/0AYxoNUyJphrOQ6tLwxTWFmJspxlSQABcOsE/h3i6e0Z
qS7dKKedcqpZPrO69h6gSQBB9a3r4KY9xflOCHBaszqdu5SKwco/rEeP+uDh
sU/1lrUWhTxHPEmo+Wi5KyPg+30mBLHmfHtuJhZGoD5iWHhCeV0W4bPxgZR6
t2k1VN4BJ2hpGv6gPrvK62BLPdypqAzSk7/bz1IjQ06i36ii9VdDmxIIX5sf
BI6xyPuom6KDJPjfaUy1ch360Bo0lulvg84NWJ9Q7GAGfCd/uCGJg9P5fjNc
wMp+NqomipNuY8RzlH8rE2KNzGjMLOOIEv0YdjWnB2DDlo0EKz6V6HUYgK9c
bsr8ewZPQAyZy8l1kCOY398Qk/LhUtqoGGZDtAItP90Jn7DR0TLI4Fhn/0zw
ctfQhbQHMQPcZpx6EU/aD+oDiod3tDVG63wF8z8zCZs6r8ce0hCVKv0mbe+E
zUdyp2FLWaVC6H9DcGh37+34zXu7I8Jypu6o67HMCW5/c9qdt6NghtUhjzMU
ecTDVoht08NeVOcIAW2GrOfBAVtZcf531aXdJg+wQfAj/JsZ78l+/ChC0CwF
+lSY63wUp+ubCjXbf0REQxdVOWn8WfwbEOwzBOUiZ+HTDkd5W+TlKZ543CSC
7p4sLaGoljynrtqhHz+lXkcPx5ZoQO8NRDXBBcU6HXqrKuRTCvUa3rlbENfv
NTtTDghdE8siiALY9J+lsjDpbxl8JTVWtz63W62qXWRL1yIGmV1Z5LzTFeXC
P/oiObNc66FjjGxM5fo+A1A0CNlaVQiUFX9UYHPX2bOy4LHWRGMR0i1i6trU
Mom1jxCdvjbdsrZqzOpyvkAQVchPvoIy1sNkV5SJ+vPj0DMxpr+qLfCS2kH6
jfAu9hNCVjdQnnT46yj680x3lmKEgbebRqvyI77D8GnrGsdCRFekPCxZ6fdw
NZvf/9CfeUfo1dVCuqcCAJxrZDoHX22n7l33uY4aQ0VnrH0JumOM2vprS/W6
33dms61sv06RsfTPkFKqhEGRMHFKOPzXqVLizWf1vzKH9fInNIwX9h/UMkwo
quNwPqVHFmvbBydx3PwTwievAVVKst+a+82JkeEDGQJV8Vwu9y9IgiIQ1Xl+
pU0Te4qXBUsHPd7cuxaqH7pL5Zh2kwbt320Gna48RFaBhf2NDPP4jM/COQ9j
53OmjoE2FTvhRykazpwQul10aoyQpRkvbIiXilL+kCk/XAG7d1CILBlYL5mW
4XqSVJOHfC61mJh6KDn/7+zM+ykGrpqmmjQ11fnDQa/pjfb03qZsm5cIdyek
xFpCbYn6WOIzHdCyJBWiJjaWohfpMfeqUbUXnkA1rIJAPfprTL84MYHu3Hcj
OYj6d06NYYfKjGYv+ncUF9y+M6EvZpZaetgLs/hFkxHkDXMiJ0XuWLThaGe1
s7dG8a5PbAAgxO3cCbzocacXTKURq6B7R4RO2apUSLqIn0YqM5QvHtqUQjWZ
NBiws+OjbRgvjyDnEQaQWEZJaNSWT8kfVsjOCbP02HfpNLot+dRPtvfOD2W4
qSaDaTjlcW30sabstYMZYybEqeUOMCtDmm3fAVFASkcH9kwpTEqjmc/ljxRj
NCPFh0pvz0TvN9hcoGqSu/2uCha46uXwIq8NHStkFKGGfKEKZh6sF2YR8G0Y
ecq5XiBMullgjWqRxpm3j4fuy5a3gUxT5CHEKW6mGL89MfzW0j3lMyOs6zO7
ZfvpIWhB3J6T8zg/ERGg6dDZxfSkA9U5PByxZe6TTXnmCkH+BPHeHuIpGEUw
dfC8fiDZWtcD2C3M303vvxB10wqBfcJ0h6qD23M9pjza5nE5VCoC3+xP3oqi
LUH4xz9zybVLav+x6HU/KjkCzfZJnQX0Neu+h0Gv8HMeK9xdQbQR4Hv7/WME
Q2FN0L5pQnHbYx5y1vFOwHrulXa93ZhYzQN/HNVOW8ttsvH3hUc53drVdfCj
ZtPNdyLx0RDNTeYcNETEtzyRO7XL82xGl+4a59CJ3LyQxi3ZXZPMhAWBWlCv
izDq3lVP7/L9TCNdBgmuVCTmkWNujNvUkFN2sJKKtlLMqTmoWXDGpgzU3mC4
Fwd+/JvADvUlaczn1iCA+UY4ihN7W9FL8lPr3KadKBA+Dw2/4UrSJ528pqfM
e3YNxgGml73rXHJEIREZy2XscQlRiQFTNfyXeJMx9933UpxJOPs9I8wxfHuW
P/+OOC2wQKqhhpPJ/yxq/OzODjqSZ2tINs9tUztiLWZ8oY//GPtOkrhHYiHv
L45tOStaaMsFWY0Vxee+T55P/YMSYP6ig9HT4xuMFF1TJoDXcXBL5lD3m0el
zqT5qO3J+gUW5D5XSeMJToBQodJP2bho1jTHtJxtT1yjB/2/BDaW8/acQ+d5
Ytx4/wpStFW3cxAwpqM4ciHImvvhKWeDn4lLXe23M0NeMmxfnESVr78ADeJS
XMLDWszHbT6/trs9EIJzkbKgJd3PMl6TH2pcSrsKLStBe9MPUPM1+qmLxkLe
qKIfgjR7XgfatpugcSgEuMw0rtU4i/xRlb/xaVTNLS9NFRd08HhBlR7YEAI2
g6R+iLzXqhKYNtEeKKj3ha8aqMvC+ireMk1jpTbB/uPCZrvtLBpaM1i2YGh7
InFX5YZ3uA+wLPqXRzpYaYIkrOCxVldfFDuJlkvjkt0TrUJqxRlpj1oZ5aH9
pNm2ImXpIKU9NqVSM7EICB+k1k3r1ZAIb881NnZs2qWtsYTw5fqijqj1S7cd
yOy6uPJBGyNPUl549h+Gr6a6w1ln2aPB2sdyWsYcSiXY3LhJCuNjh6Ils77Q
Il1kJ1iPbyHuJ0u28+4vSCpxbrMuxp5WvbYCv/8CAtK9bgH+CgIS999Hy+1S
78eKncdLz1jznqXSelTVswmE/rRZKIaHgbPZ4OBvv0G+95aWUABx3u/iIRuJ
PX2uAsPwcWjs3Jjxo7gaLVqP8gu/OpgCY8gy2zsbOspqc7PQD7musP5WW8XX
OcNCfoeB9Ga3J1uIgtrRRIQWOmUQX7lCSLDxi2viutlZrRDBBi2Q00HLqPAF
Ur3oGRyp7XgvthItUOyhRHXRfvJgb72lwEGx5VWYUMDZqX9ZwHRP4zdSvGBq
gdczAuo9/LGL864QX5twccVeBIzx9DrYM3PEQKb2T9Y8qxYx2sj3mI5bbMMN
3r5WQzIu50hve5WHzYEO0hE75N0JyvOFp2Pjs7bqZFflU1Bd1SSisYDOw3eV
2dI9mWFrjJBmzdxXOj3h1a6RVIH1ue1JVD4doQNSPRrV5D7vYL+6WBSDS/ff
Uh8xScLrw2NxJd0B0qy1J5dWqgKKn+NJlvYF/xFZUzp/hGI/Q3LMU3hmV3ed
2tnakSprgU4zS68r07KTlkmvAV+17FP5GtOmla/zhcreYUlm6vEBmtRwnkXH
aPaOTAO4s8CBdRb6eWZVgDDb4eAFr35e2m9tK2lhuzfztZPFQ8aTrbxuuPzr
mh2GUhc6Pd8tL1hT11OUAXIjwPHz7NWv6Gt0rLbaYqJAZjCRXZd5TNJGOT/h
ac/9AMu6hhRO7TyCus8VUAervTQqAu5AGY9uUMA7ULX4q7lqVQJwwQAM9JbC
yYr8sITeb8CrxQQieyxEJA0kWFZDyJy2pW0khudRYwPCp3/KZsVWY8fvChj6
FNvDZzeCLcEg4x7G9m6oHZwvbdStxp76rdTUYSLeZUNc2KV8H/1O1Ghzo0LS
bdm/d3ofmTrXhRdzy3IaFtzTN5wvw06/sH5XY1UAoptX+lJtvbNdEScEsFlj
V02qPMJgI8LAZswAN++cSxwpfuT1iT2xPkPaPbM3ZzN+kYamj7Qv12GfmnLe
U6CdYvWFCrfHUe88nj97jK/E592T16q+zEsYpIUHQd/6ts6yvBj0qgDNzXD0
94ecILoMSREuOfGR71rZOqSEYU6psSSaT2wn8YNZDrXfpqFmRX1TgNMSBiwL
2eRzxbDMIN23yzdFXf6Ef7NMz6Titk/gHr00O5WtblCzF1Sl7fLEb3oPFkHJ
Jbq2ef94WKe3H344Kt2sRnfPYcxu+RJJlm6GXBksaNeOutpXy935zOH+znUl
Lm0n0NlMt3sW1agp1KMJog5tU08dsDOJwreGqR26OS1W/dKJer5CXdEr03Sm
dnIch286pw0cM4ZbLNWnRj4Oqn0kloz/JQcPSqPRl4qqslAYsLZgRwASUWOC
IiBmCohK09fGd9ixNBnoCqSJ6fHtNa3VIn7Vei0oIxNhftgUXahvJ3w96Ac9
CB3IvA9H0FinrQ1BOpUTrZ69Vs7y5vfW6AomYd/MMRbE/x0Kcgnj6DaBhZam
PL9pdAWbyiDnivjDAxIovqK03Hn6z48Rj9Nv/VkWkDwUaK/UCfEt7bMMLP+S
IHIamD3tGpXfsBGHP/FhcAG/7q/6kjwu+rqNF8VIzKyXooOTXReOEWmnFyOI
jneww+itmp4cEiMqAS1R0Z96U3Incw9DI1ZSfkWSlM/gwJ7za91qH6IbC3oE
b1g0MzFHIDPEsORLMkCM2Tl8GeTkCkmW2FGO/u8HcmxY7Kwv8lB98OQziu6c
BN1Xoyawi5s2kXpKAgLYrhsH6gXqmpUzAMDWGJXVFndTcmGI89ggD5sTYr70
VK85yTBNGBRg3YModPEcnjHW2zU+/Eo9n593tDWVW7RjamVUJAql+PpzbXEL
cRhvbB9anCcjOS5ROcQZnZutm5GVEWQ8OtXxX/PDIEafV7w8vL+JDjmAEJfs
JyNzes2yM8M77vol1nX16dQ4wuO97FB5Um20LDMHs4X/jpn2IX0hYOUl+EHO
UJsYg4RNme4eeeHutllOSsfS5c8+3RlNZSvnIq7lV7IAbrW3hx+wJfrynPo9
9zNbbiM4mqchHftLu9KeHvOQ/ll0dWSojtPZnzDKBhb+o8GfCgSFeZfUBtFW
VhWTD/nCD3uPASMdoYhOQloE2FuXDNNPbPk+rGwwzhZlhWqeeaRQ+h+iYKb+
Z2Pcf+i0yaeKZa5o3s9iz5Mhx8a9qS/if73Tg0vNO8eOQ+Z55aqW+JYZl+N4
L/5VNPrVo0/eFqjf3rGeW4/QZkOMGg7+YkNqFOu01vGIqRuxL2QQMtgKdr1a
qYTGMwiI/on6tuNn7i45Zilk/p+yB8VCnsjW6+yrZG2ZGGVZj47Tg5TS2Yh7
r8XmJWJKqoMPyEYJFuYn8Rs+gPEbULapwhR5izdMa6UELCZVoi/mdKEOLs+B
uox9y7abG2pAyDEbhlGdvUZBasw79y4YtYVbV5s8vBv5zJCaKZbcazugfMIL
TeOyaxaqPzoZUF4KFVteLrO4rS2iFMmwkpGZOVgQdzR1lq1cGMzLLds/1Cpj
lmV05dFPWUHrRNhdcAVd2PYWZ/UDKtdHMDEJsxLMt939UKutrD3AzH0xnW4I
9Wtr+w7C2lIVOy3tTzJC/Oywon2U9dW4M+zCjv5uZiJbs/0e/c2NdjA74G5J
POetJUsSONZwv2QKxg/xr0XvtBig4BGBxar5LFLtNb2bqylyoSqPleNuj8EK
GA0NOco/57AZg/TAV2CUlOfzzXntKf0dhZbbEfI3X4M52plfvg7Pz/jfrhiI
f+6GrV/RFE9B0Ldm0J7e422phn8FLNzvhrA4eO7vvLlbs2IdCMHx1JO5NB3G
y3qNcmCQKVR3exyWAxev5lpq5eUdyhdCW8ozX1dEBEbQBSt5ylcrfPE0hIXC
7wZ8vMIrlS1tGxkOV2ZNb9Wg9jdPce5rnMi8h4gzBXQ6+rl2Lu4rghJE+K0y
zR1MGCi6W5LgHhAou8W8vnkkrQuPJR0nJs1Cje1m9ARneCoyXX4BpYYChJp0
PLFiY3JcoetWkrj5HN+npINinSIzSlp+jCZEZNWpumPmEmu4QZmidS0HsYEJ
JDXM9W4HrjRcaWzV8OAzCTrMj46EUVxG9JxpAqPOo4reSsDq8Wk9W8ctmm47
Iksypd9Msf8BRmH2TYm/Itb/3RGrekC3i3BJJVPYkvF9LMN8gJluT47W+iC9
3lYxcSXt5sSokR/xquTXMNGz4iDSsYwxUAcyVluSdfbfTmDV3TL/gVKN8St9
UiJP9uNZS6hdh4/eN3//hAoQCgWcK6S7KUDLIFe8OYrsX94bphaYZONtxyQx
+OtShZ39M80HuhN516NCmx69dahVIqlX42PLnfvWKHhD7k/9Cwle6LumREw+
6ziPyn74+RcgxS2ppFn4zkeDZyxizfsDf2lve2fGHNJJJRaNHgsJYWRGfCP3
Es9BnbQqL4CDTV5i6L/f+pUMNYaT4Hp1EPgg1djtMNOXfIZPwk2idrv7wxVA
T1NZjHO+FZqpC/jXmQdHikEyAjQd4QZ+A0mFVDTaGxkCJiSq7axeq8eyK2Ch
rxkMR3WyAmevZl0IF7JoCw4IyMAuWmIuYDvJqKTKhbh2eEB9ll4sf8erxglQ
m233MMSTuWLasr8cQeYGaxnXx6cnwJQIpGuB+3f0IdZ+WD2iSmtCd43fkmS7
7W4hkDX6Vz4e+njSwyapIItrzK1CD4ak1A2dXEbJAUvx622IrlGQKBTtluip
GpUekKm1A71PvH/7dcFVx01t/LdqixfK6dxuzXdVbIk3PnwAjfUn6r5jFLVF
jgeKdSGPSTV3EsS9TcG75oqRYEN1MycmYqCpSSNlZukyyT9HrBFnZIpzh7WI
mW4UCdUidkAh5UR1TFUcLAp/WVs9E/zznPZTuEgOOoXmi+ych+lMKtPDHL+m
UrXeeFwR4z9EsuAwqSJl3kEA6zkgPAlEnPZErnOnFgXMpbGizGb/WKc6aQqR
1GTVviUboRb2XGEcJEf+F2SWHsJqIkDhMmlyd0LBGUT8DGt1OAfHfuwIe1Ph
zGE2yFAOOCxytzYx8w932Syd+pqKw7f+HUVfAcd2r1phD/k1ZESLWFbjRviV
h9UWXpv1CVwWtaaB+I28bEqHHVJHGtXtr8nT5hG1dnNmY+KRxUWskRXKOglR
NPQ37fRSFHgj5dFlOFEzBOSOyReookHj1K5YroBn5EIZeFpmQC+mgZR/o6bt
mRxziYE6ZpscNkNVmAbYGQNBwofm0Rte1tJwjBNrHrvgPVVwrQ8s5zmxYOyf
RCANDwiCtsHw0WiWEIxFWC+aypczy3gK4fbPTosKAC1SfvKnoxWkagqBuH07
3lYp0wT92/2Qvu3h7x4CVJkYsoeXwbNYBGmdtjbT6DX2fcqXfp2Hp9MK1Cm8
AjyZnjZ7BYUwQgYl49wNxn+YidHCzbZ74zHQZFkpbdONf7kcgmRr3Rrw+H1t
hxMi0dov4NhBEj3IA6pxRSBY8tS7DTRo4g3rjGtl6R3KglXsMnuabPGAIUej
evSCIHwYDshdeJDyMfdymW7i/4LWf1RaHyJnafO3rheaMvzFI86Ohj5UVE9+
Q2/eHssZwygNVEDuwu7uRQuSZPyVotYIFYxKqL9ux0lMaqrO0bK7h+nvQ3Vq
A/RbQkCWQ5Lk3j3BJqJWuyXXlndoH2Gw6Qd/pH1ccXknw62FQ+1qwvWaAnmU
FZ66c566FD3/Fw51KFmN3laqcWEDpE+BPJzN8IoKwCdXGuklGl3oONYiLfO0
awZ/EG/4outV6xmYiUum3zn3gvKpaxk55YYZmBZqyyrlPR7Mug4t2jQpxRUb
AO1/bXsEr02Mzrqfvmtx9hMub/yEIOCxvDoxOc1hJ/AqJXZ7SCXb0TI2NvbY
ZRl74JJWFWIypAlSb3z96x+RjpVVQ56+70HaL5eJdQ0qyvgwxKfWqv0jFRHn
fbvSZAtek7GaoXngQaOGN4ByeVcWrVYTiuTyKLjPZUa3kF911ARaWkwTlR++
1YfnrZbFgR2PeUw85sIblZ/id5waaKiMPKlnt8jvBqoaALfJD95b8advbZcS
7Oz8/1cz4KzCnVzO9AARjcPBFOVo7UwQPTOb7FAD41Z0JedaIERQhto2WAc5
4vleq5OTAN9nx6LjK3otvD829JVFPIfO3pY1tfByE11Eth+Kt9v83siJSkVS
YdLIXHy1Js1v+dSHLILxDI0NNIUnU6maN02t6ubSuDKnL7ojB02p+s2+5lp/
f3XO17JV2KMm09yjeAL89+ZtDaDyY1znkCx8SG8tux6agLaUTcZYUiTriEtq
bcbniBl64iRRsrHPwJSY4t4Sgk06STlhLXuuXdZ4BP6an2EUzONLF4Tk9jpf
USHKQhA3JjFJe1iyo6uIoH1X5ihrTZ+YYITNp3fFjiNQATicnSqtAuNqNJes
5kw7tKUl462dvwbaKYQ/ZZxf/mdRYH95PDjQH/5+794l96o6lzvr+8Awoagn
v670k/7x+OrJN6FNuTZoITUxs7a5KhAPPhsqwDKCTV+zlZTU1OVf9vuAOCnv
IhMvL8jYuUH+H6GGy9AC8/SfKnntbELRq1cZR7h5F+58QsEWPFgtqLdml28z
a5AWOhA3AFBxLGjePHovJTg/Y9Swyo+5jwwc0/+0Mtg9kfuLdeR0dDWHfJ2l
t8Qv926MKZeFSz4j9nnrJzd3KwbOhgAwJrLBi/YSDbaRB+IKOsWPc/td1aVl
DYW1baAGrFChTaowRoacEEHZhlZx4wxKbGzIbKjJEuqcDnp/diG6jX7RUQKR
pr4FRyfERLrj4W5JO1/qpNCOWl2d4Bh/1cvNuKceybjmy0zf9OQuBerCa+g/
K2MuQ9Ox0QBDqsbNkW1LAyt9wJVg4SVxXiLKwjjk12+fLpHXyu365cX+TgMf
CO2GM16E5zB1IN3EUJG7xI3+YIsTXoUtRW/kh8YA5tZu/AysyanMaZ2V+d87
hz5PZbTVgr8mlXBw+Fx3gKpknNvd/jtr8O1qmqAhfls0Wg8MDbbJOIka2R3F
GnxIdasvQlhLlmw33075qX/IAIGlMkk3OAalGxusHVRdFUDqI5laP0V1Vtu3
R3rWh0cVJDK5z+CK7virWK6hw0pUFMaMP1oL6k1EDxD2ZWkjK7n0a7Ed2rzn
5215fqBwxZ7hNlYnrP365YMB24pWnEYZYDGJHyuAp7kJYuYWbF5FrvngPd4i
k6HQ1CRryNknuQYdghyq+RwvtUwTpi3t54Jy67qIrNDJ7Rja9q60i0J8kUxp
gzWKgQrK/0KPj7a7jwVvW7b+pLQAF7Umlyl8A2UAwYKD9GJGz0HQ38JFn6is
CAftaG3RAdW/oEkCtfRz88m/X9zzsa9MPoMmbjYBqDTu3cTOgDBn0FHc78KQ
cr9+hcC/us9/kpA9zv55N16hXQVTY50AvFMuOBShfpBOoUzuLiq9NJgRED4D
Yf85XiZhy1fmFXs9gWSo11sSUiKdJbGO3i2xq7q+0amihWop6JdWoyeIsFSg
4+B+ug3Kc8HKIjbpasLJmh5v20eUUBXdV8SPE42Xyw9aTHDit2QSmjQeCrE5
Oy8VvH4kvjz7nlXBrnTRwFcZIRaT39JVRMbcqcDMSZsXiStQ/J1XJ0JNQHrM
m+A1C+o+CEnAoyA92SQNziV3SyAgEvBxqgSS5Hf3hXWKTCW2rY5DxCDwPQm3
Cew6O3GTdMROJc3paTgetXk9wtxY2s9KqxBpvC+BNZEsWCE1LU/mxStXLsI0
d6wTKDHbpCJQ+uvcneLwv40kmci3gEi5lL56x/+ajY77nHqsmzN6t/Ld/uWk
wSIHSQCYYVG0I0n6i68UlfATQ5qNYokDeKJBozja0g1dAiMPlVUdQj1YID1N
ATSYK1RgHDnwa6kNsuXHScmBLAZrtWwcJn91XpVJ3EoW1Z/OkmJpHbVtFNKT
KjrVpg84kfXBdO0XOKSwPt53+lpjp51xH0HmFbuJeyFke1F7umoXG/eIFz3s
iKIG/0vssBgmeiXGQj3SffGY4dNVhN17bGE/NpRwZwYjZLJdPjoylq5YLS1O
xBUPJpjvQnxRReI81yG9Pg9MJDW9FsCVZjll96ZQMQJ+iKPJ0P77nGjBi5Bk
YbYJkm4k8Tc2ou5XoarINzyCvEe/2pBdcP59nOD3cYCyvaaM29hu7Q2tJhrZ
z8oOivnPCVmI9GWsqa9rOkevBHGbV0YIVLp4d/ZUwq6GMK+kjzfKxh1prNeT
jlrXenoPaWttKRKWOcH+wj6NMpOjIT1EMospW6Pomcx/km8gLr+GcUILX/L5
j1JbF01LJ4hP0cTNhXu+On4Ns9gBz2S5UXFMwyUspKO8QWhsDKiGqCpmBquU
Uub3sIgWzrL411l0B1pTPqX/RPjrO3gG8+dJJUK8JJQT83xN8Tso9un1fSSA
h/yJkL/+bXJFrPOqv4NRUpRKF2jWSdwXdBs/BxNplvrAk80Oh290ubxUaJFf
LqCPWFTo5HPyBbuPF5MEOyuOU1NAKQ+RcvgpCpkjh3b5NUUWuEHao65yEJ1U
pNE8lbnlXCEGUshYrDk+QCbsd5of8zMABqR4k9DSaGmtnus+uXuRGjUmjex0
/r+ogEpEWXwR87QOFQAZahmTwNuEJS8KMI1SpL1gEtAaOT9/Uz/4i+LnzQFK
uYc1636uKY++i9/tBOZT9/dFMFaHyCKBacK+rumKnn6oYja+W/pl5jq+Xa+4
1BaBO1y5wGdMyMteCCrQX/oVpgfvgb4TW62rhMJKSo0yueZBDqiyAB3AIl72
YJ0K6mY70zehpW4+oluGWUGJPgIuCYTxsWUPSZcizT2jzu6cAU4QbX/8dQ/j
ZJXD5oM0khHvj0eFAv6iA5SbtdYuKV/X1VsJ9hjA6wgfx1h0OOvEm8mSMrGM
bUQgeRHktRa+zS9OCiiY3uLo9U5As2kGvKMOvoLZ3Mhx+iWNacMkLqBurj7b
aAq1LDq5Y7aHPYKFA4ZuKG1iUrpUOigvtkjr+wvSLEkmT3f9yTfns2LsPFme
sE2LQlIF0zps0eWatfKgkBY08LgC4wJbnr9d1Na3c8i8qGTmEgIeNr99lPc0
18wT3hZ3t/UznIlJyveOK0vvw8X9IUV/E7SotYtclqHd+SaxjsYE12AOg2RK
CUkaUGi1Sjr0LL3y4y+A1BNgSjiANXzB/R+1XD0RygmNnJ7PjSYVts2xvKBr
vY73+sTAahGAUKKgBqgHPqj/GFUSSS3cxEvi6CLURp2vH+Hki+RuKnVebVDf
hbmzgKUAELTBB3CRg+qHV48bwqSfY40msdbnAr/4bVYRNTqzbk3YmJJpLz5+
kOzw44ESy/cF3gHMSYcQFoPX7aCWF3KbwUWP5gRQ/DmdfdRFIGmjozsvt5rS
2jDrMT9pf0V00dl1AHM8sLMFgalB8VPgcFSaiha15tDfuJIsZ8NSgbEKx54P
QPTfC5aUtSb6Qq+INU8VqxJfpxJBnFGWOybneRKunVTfZVlLv1TsV+xNLj5Z
dGUC4CtpJaZMejKr2f9uGASMwrd5SSSHMgcbJSlmaRDMXfImSjkiA+LqYESW
q121YkUq+d2lnnUqrGY2pHpnXkKlOaNiQyY6YZgUYLTjQmF5uZjZ6YysbvmT
OM9jzllIyYjcYPnZFHyAKCUHqqnUM2G6cngJoDO9WzjE26aVLo0tAl6nghs8
PzuYm9n032CeA6NiJRKN9+kkbrXPKic2C4lYbkK+czYrawAJ6lC0BCPG2o+6
Bz0pzmwU9+aOC3PfhnDO5UAx1NFLjnOQk+GyWGoa6obI8+biUvRyWftNkbCg
jRAOwEdgv40D1YcS2SgSZH365D8imxMX/m73YbeGIQm6GnQwFg/MQWvA+hi1
I4XQVyv5vjdJHMlL3wiqHirFg9/jv3HkkTVxoMA3gV6Z5UM8ePVHfivvAvOp
axQsmIpaTH2qY3WwWv474ZUdn2ny+xMWmjIhlTohvzpSoDlUniQNP4imqxS5
gadERUXKbkswb9/Qzua0fMSD5xVLEAyrT+fz2+jso/1TSkgZpBDv3nBPhjVN
KwkHLdJLLXLS+PPTrep3rR8E2nWs419Sv/Qee4bRzoOGggE8s5GdCVIQVIkH
yN+IsIv3Mm/6t2aPKWrzAlndkdK/e/K/DXciIIimGUk04lISbtw7S2FUP2CC
N9XSp7fkukvQ2M8zBHMHobk2MvsUrRP+9Ilo+pHL9MiEiszM393imj2yf3WE
0+cuKcfvzhYZucq/TPlmsEnaY6iXGEa990V940fwr6oAFeQIGuKx37oixZed
4e0x7p58hsVazm6sP/CYHc2QBDU82BgmXAvGGvGIMba8CEZM+Nq5mArA5MuT
McojuxOJ2OVMoruYeGRmZuoE5JqHKrz3rwQZSaj/L4Xxo6qI0zPkJBwweiIR
nwTnVNq0ya7h6EoCIhWZCFojE8BXpY68S2bQfFYg+GdhF3ORDpeoZB99S92R
+//haxCHdPdcfr5/olkRj0LTzpPSjL8ycqtTOQ00j0+feSVarE+fCtHD4GTx
9TqYhzCn/i8NoPlvSZ4uE20XCk7ZAeHydcQ28sclg6yKvg9KIQpHfdb+4BR9
GXQSo3GYFxm6KayAxIz75PSrJaFvfX3K5J6YC1EnH1+fNprKv+Fi+nDBi2rh
jX8xl2EV1mULpLwlAgdTRmvRZ8jhprEtzt1yi75cUvxciFDUv2l6v1nnEavK
0DN+AjW140TkuUwyArydHKAd/nEWQItewlJ2iZCg6fq2kdDURySSxac1MBaT
QwQExDI2xMaZfmh6ftZxTi9gVKJqsigpazoyL6Syfl/uMFD6ywdHuvTY8chv
iLENJeyZ/bASm5Y/8RvOUThWd6ZzzriLh/NmSVlzslfRh9+3r5+BCAD4wuJE
yAZ302mUdFWOSPzPUVjJn8w/db6jDyy5BEWYDrbbrLjT/a1aaksgTRxz9qES
GmJv0BGrFMB4BfVRqILxstXg7g3/7s33jLNuf0/YVvNsG1lPBhm74K8FPoIT
lM4k3wbAU/uTWrWJHAgdOXfol5zwJuIwxxqH0RfROFJ+D90QJs+US5PX1fQD
ot259wadzg1Ze/frjtWoPghg0yiW7kZkES326PtcO49nt9Jzv1lSOQgagwwS
FknjYVeoO9jF7fLSQEbzFS4qlBKTJbjoI6+Gsg2fsB1axbLHSdrjbu+oeDq8
DuuBKchHaDfElWflcwSoZXshvRxb5jWjkDtSSgBB0jd/tlGTtyjIKd2R+P6G
eHPOET6DwcyHsBB2ZW97+gYeuWzEypu7sqMNbql0d4DpAjH2SCGBx8c+RD1B
a6DwlhTWDRcdMu4iP8SPj9Q63oc9Z47pw/FXht27w16VePIqHNPU/UxYcTQw
uF4jzRIlkBVA/qsL5iCpXeHFtRLB1pXTigQlIJhq6ODod4G52bCYLdXZjBWB
vYhRjHTKQB2WAlQhqbc8mRdKjUj5ivlDjGcL1qNBO1OYP7q7BJgOJEUV/NMu
n1jwMbGjdRguDEfstEF56NumImBW3sl7fz9Dh/7Weefb8jyJRF8lpr1FtXXA
pFMlHXPSh2rmyrehQc4htsa5C7GWRb2aZPvpEezjzCKv+HiD+EQPF4DF4pRm
lj9PD5u7wuYhlAcvbhOUbI4iGdL84WDSZWMagAjnkZFjiv+fDMNIKI3Wm+sF
zpJlQRVOyzqtWntKcN94JCVeUhzCdGTtQWDaby/m5GN5RX4M4cy4yjYApKmM
cw7YQtdMpk7njRtCuag/QIp3q2c537TP/PvfK5UagmU6vzO9VuGi2hpj4sH3
CiPc6QUMvuZxrg0mjzUQtJdzN6uEF9wqWmJxYMltlp4CTXnMN7OtqWPKD4Z1
QOzRpM8kb2Ck0ckQna+IDdB4IzWnPJTJImfUh6XbpA7BcTAYUv+S/mu9N/4H
6JDdhxwYBVD/k2jPgOXMk1ag9DPL7bg5hHd9m/ktNzJZU4RnCC0U4SVlzu3K
M2kWaL6PmW7NFLQcuWKy3XokgyYLN22j7TBLUlm4zMiN3cN5A2/8MEhWI3iJ
l2fnAdvbtKx6VonusYce/kEPXAak3oeoeZAKzJOnXoNVuVKwJnZTMj4iwIVt
R+jaKmk2m4nrFEnKmPmpoX6zaTb4S+MQgLMq9r6JELGe/ylRnqabtdIpF0e3
gugEF4i1yK29pQjB3JijN+o5ppyGaefdf2rf0KbfOGC78XRQF69WLbEKmehJ
A8kTKj6jFfhaQDhSt5mRA9Us8utdQXcRFAOqnFFsFq9QoKVzaxnvrfGeahIl
WKhriLpNeGNa2Yggpk0wng8MxAPL3M/7wktDQfq+Shok/65Wu6KYA8mtVXxf
1gLIKVaXrPq245K7bNDRtcRXmYex3+cfGLP/UGyiZWkvXt74R/ee4fRCc4v3
Sd2ozAp3dPzFYqr7Ob2lZYDlYOuWsJbFQOYE6VgX659ElvMCLx2QTOSOHjbH
5pSRHF2+QsmCfwOxOfVY0K3cRiufkwXLQdPmLeXV8Oz4mrbHpw8o3pD1jKrA
qJitOXbatFaFs3M0ainLr0ckAB2v8bUpADKHi7o3q3OTDRDNNv9/wCR7ovm4
MEWqnCwyoSm4LcHHyf3zzag2pvf7oOAHp1Js0CpTQpxoMusR7JSbELnCsyPi
6CyI5Upa5rdjPqsmw6WxFLJEq7UcqvwM9Z+aJfo8Ix+PfL8/hZeWnAf6ZXLd
1t5FQIiQjGlqK1z0nwmEkQsLzopzz2QFL84R1nIF9AYgS5Cleil3GvYwmw/x
ZrgqqDXiyphuVNyImZ0+Crh6HYH22mu9Ou001pdZj60tlljYoTodnH0DrOcz
oZrM90Kw532ErNUIU5SPV4Ynj1MInh5wePfsQshwRQGlJVDOaZJ6iEdTHacf
/ywkA+D++Png83KZaJYeXrieDIYlT9EwmjXCpadqUZpZ8Z8cIay40ccmCS+s
PT3SAjr2WIz94kKgcsAG/uzSxmSZCJnpLPPqvTjC0s4n7kQiBMYk9T5wWQWq
CMxe02zLc/03wwtSykCdLdE0+mV+mpRTL1SIAaqzTQVJpWCDSWNGEWCP1mWR
vicpzgw8ZvI428zcHETxSNGqle2RpQzX2f9qskWe1aQZ/qQq9L9mqLHNxFe9
2Wa7fVZ9rnCzjB3fJIvVCOsjnfPCmb7k5qjBGl4td4NVbZxk6rrd36/X4Xdb
FHKJcfVXjFe5q2GQUKUYWtmDIiYl34iLb2DCsW7bm3Y3KzAiQ490BF8mw0mA
flt7Ohra369pMurzd/g5EuYTFXik/Gvdoz3dgGmZ9v/VIRDI0eleJXWNbCDI
Wjmd/nuIfnszHJooyLMkUeOlpPd452yOHi0cOLn3dvptdSu+qmOYnZ3DWtx0
b9IL5xRyiIEW47WLePRGgXYbufr1WPYf/cFrQdwJ04chpUBNlmDt5KXVw1Mz
7LhEIuFOvCrH4FFbAj5xBo1wGFxlR1j0XzYybDajV7GuU1r3CABhghOl5WYh
ODNo7VIDpRaZsOcg3PTGMxcxrmjJdkkdhdYQyE+pOGh5a3K1SPkrlai3EFHx
gmceG8lnXa66PsCMuK1OliFCSQtcH28sNgXf66wUJFskQd2Jzc1kONOKTbT2
LfeaTwi2ysPUIwiL9epCXh9JeWbDt3HTGmCZGhQB59K0NjqDrGwxmv0PbMHw
vDPdEAdWOa7of54DaNpj+qMb2P0OiwWYMQMhW+CNs9/MCmX3qGNQIAmgjeSF
EghlaSU1coUeyQN1f0mgFhUNAIz93yLVLaDraVhNr+QkUzc9yWBkGg3gffm8
8ARtzCuvKtiOmRsDxW0eIFQCFP3B6o7e+dF0xcdJepnUBamkYkm5hnT7UoVb
vzf002e+Wq+mPO3XxLBCjM62h4aDaaYNT4Ia+kr2Iif6so6zMg5duxW3SXj1
jnPVtu1PcFHn5CrHWnCoB1tYD2bKs+u/qH6rT00KbsR9hbfTxnvX8MCPos46
7QHs7Dlp8RKkzWAPldU3UD3vtiDkgG/UclbZSIedy6MgLCmkxj9iQQQLyyuq
YWN1/IeqC3RK9hmYzMIBYhslfTL8ni82DxddMo7IH0AzPxNJP/OzSyaXFy8v
vuyBZ0O2vYlhqe9dwuAb6qTohlyLTe4ssEGqDuZXQJft6uzxjHU4H3clXLjF
LJW6K5dqeP7+Yzqv4JjXpt7Fs7K65yx/iILc9qNDoScVj9wKZo0OJXVk3Og6
5TE8GoNY+FZPoYS5xBLsNg6+AcQlNopRzHwB3IS9AHjFTllBpGB9YFAKR22Y
Y4AyU9TNcaL00THYxocaAQqtjJmQUa4OaGAV2YtF/o9eEJLuc2dlliE7tFfl
ZYDxOQYGMwJpU1gIzv/0rOukuwzFYWwNBv2Un0lTlGY3bchwCBrreVe7LNRA
Z1QbhNFS3j1e5hv5i9xXJoLiYCvbkDjDDjM+LvR1VldMAeilpBy5SGl2R3+d
hGfRKJm5uCrq6UiqFfywLhFtPr6RZbj9USCdcpEHSFDg25qjV6ITUnvPk2T4
aVGr9tcjpdENyjpqFrHb4FDYKV7I9VtrSZ7LjVR5gRV04DlHoG9IvhHS2bKY
1+AE2rAM9TVTvUpkuKN7ENqmO3Gt35jsdAamZIwrIpbpY9ZvUfGTF6zyj/d5
t1pfzOkMQrE0u0ZegfS720XAIdgebAp4u+L87VfFOmmZwNTbK7Id1HcOvuf/
jcQmyjzPIPR6uGKTj54IjlTErYNsugZNtjveVd7H8e5kPxfGcGiFHo8AU7bm
oetC4uRvrorP5MmrLc+gTU152j+HL+2h8M1MdsvBUjA69p2pV2UYLActKq0m
cDLl+GSkNZyBCjEvZvvJDwPGsP9JsOUHdvgQ9E/UGE+11Vf0qcnb9j/bGSFy
tIKHxH38H4qjD41cavI1eYOLGESl3zeRKqI2llT6i195yvWfesYCQ/P72OV0
hNn6T5/15LUiM6B/Sm9TdqFhkW9S/RQtsxa/i+wuspQVhJKgxDbQzjA0ovfu
pkWOyImWSHd+8hkYrUL9DrjNXwSBjxk2vlNLDdHP1ILmctLbYPSlk8DIzTi5
87TD0J4yNeFI8b1CMEpjP6uVtwrTOa84DFVNDubTC+9HEYpepgod1xTHQVQp
Ib21e7mfrT7YqjMVftw/q+O51/p4HEoorf5WU5xAoRM1dvTeu4zNQgwMgqkT
t7Zccnvk0NPJ7fM7LZgC5iEAsGSSdh1bFjB83PNKF0/CsXap1khClwJymi/H
lqC8nZyDqGtIwndN4r9cA8DqeyO1yL9gaetUaLc2wtC85/pNI7uBytPxFvsH
IQaIJ4RyOWXrBGSPEZaqNUM1JJkyIsn8O1qFNSUQoo3+vdnH+dDedJ1CT6ZR
eSPfDKVlDFhgskvnndGtVS7aPqYBF8GZLH8utg/78IiZ0YQRR4PoDjkzl4q4
qI8di7moMyszbs4Oncyt5nJu9/Y6dyOt0tpEtJrTSe2ZaCzGaktHmbrLjQz9
PFlkKA572BKRpUdVa3aNOccnvsN/O2Zv6yCHXTzxVlKaCh2lKTnENeSluMTW
aT23rwNYK5q2xCyoz0p/3quufKrCQ1C/q66d8z/HaEVe2rDjHFYBz8gK/fvW
4aj0GI3MewWGD/now0b2ofUJ2xEJUAlQVOo0LVmngz1FJG0DbZu5C7sj2xzw
v+ToB6uZUp+YUT+8bs6qn6aiTmUBOus5oOquqyzTL2evTFXmXEftg71Xx2qQ
a7LamHK4USm1zqcy3WQNTnwdBiODrKseg0HcoxePE3VgYgo/JxpxnHKjvLgL
QEe47oNq8+ZXlIP/hXuoF4SDPtQmvX0YNe5b+KCo8FUw7q5DosWx3pn/5I7+
x/YgeOhz38VcBAjXmzllSS7TeQ4Oooxn9GApT2GszbqQC2uXptNK3gnLi3ZF
j6VQ9dfpQCB8AVTsKSnQC+PpVHRitXM7uqc5xL4LDwqCXARyoW9LWpW0bVA+
f47rLJ3GFi21aCF9ilnaB+0IVY5E6EAJxWcAFoAlI3e09AvAPkOFMvz2GIIT
6t19f/XP4JZ/zJDvA9VleDSeibzDEivMwY0zMHEG4GhXqTxkj8rGOkqZE5Lu
TsF+v9bHfBVhoPoGo7nbZ4X0wKjA4RBLM4X2w2o/ClG6Q07yNeFKi0GRbXyY
ZveCzZ8nEunpBjjaQEByDP2PwjgYpPKWl6KukgaYh9aBoSroNGrNzdiexlsl
OP+BCiMfMYWebp3LRVIP3RS7s9GzHkxjA4cr2l20VtRvXktMrz0uPUfIeb6O
Mj72AP5KeEJ02RgziLqhLCKhNFDQhrJ4p/CTAYOZgcGXy07D7tNMIh3Ml2HZ
geh3mrhAccgJz4TXGHTPGX3x+Jy84LUD3nU75pkvZELiemo7UsRiZ1dd9P1L
cir2Y40IrAfg8hxjRLd5Dpx32y2VLMgFgAX1x3FQOTnOz/kOe2LmLB7SOzXx
I1gI/BkaZwOgre9BsoMErsmr0NH18D6cNzYDJa4JChCZD8bO+J31UF8genkA
Zr97dmrnIxZZiX08/GwtYeqooWThi8G7fACSydQPxkAHJVu0v7B7HGJG5pcr
YznhaRo+SeCkiXJA27/DVxnKbedFakNBTFBX74B5E7XPP+klRSBhLNEm0tMf
r049DV1pYXq9zs2YJ8XAD/ol0vMDUBpGHsX+CXkH77RqsBFMh6ubSupY441b
E0/I4o351Nz1tvgd0TcVDC7mGu49HSNjr//gPGCR8kE7Zqj04d5qnZXO6kOL
qwz2C11J/aE+znRcZO9HJiY57FsFeSj2PVlr+syGAgOagZ3arrsn09N98xXn
ny8z9HQeh7u85phuWL2eEvk8b2WVZ1vP76ROVAeWQCp0bYHLo5JIQFcD9hMP
QJfmQe3jvIz75UO/ilb28T/cw7ySLkIRQgvkR8CWfIFy1wQ8jf9X3mLsseh5
t7kAWeFFBs7lO9h4GKL++ubAEpZExu0X4vwwVIir6TY41OFJYDzpkXfmAAEu
0RWoQ8J0JNvJ3vVDbl+c1QlQtIjulG82GAwnbvAeBxJtb2MIw+Hha/dnz+4w
lPQZg27xTwZ/KtcILqoDNirtEvTWjlzQr42he32UNfm+uSKT2CO0RPTpoLNB
JuLxQ4CmsvGdNQdgZM35rc+MrOrD0hiDZuIfar4XG5zqpIvjvOPtFN+v+PYh
35C14MoheQ6DLKCYlMMe587xInTQBz/80hLSoUSLPPv08Ms20xgv4Fhi1xfs
Byg1+VRm8W0oVGsCEvWL1m9p0kNOGYmcLfmPKqYKiAtUws9A7DUfOXZ9N7vb
HwdakTnCwDNj9Xj8wjNfzEU8Kwm17babN4lMe6ol0afLTyLReX5JsgezJOqH
SJcODl9+wCxPg/oFCwSy0LOmH5Xm8/wE95iUPcl76PhIxMsjMdLFZ9rVpZJQ
CLPXQpIvdSSw5D6arL/UI45UDXJ/bqh4LCO/mZdMb35kR7+CtDzPBqGbbQiz
k4oRn9itHYCKnJDc9HQ3/JO5KW3qXZXJpkBM+uDzXBtVkXXH1nLeXYnwPz0N
QzVn7jKXi+c0YSDTrd4St5rm1aIFdDgwbXFXlwW8LOTAbQWt06Lf9U64Z/6K
gl9oCnkhOgaI8qHBMkp9BWTWqSr0p7vT/w/MaSJiQOryuKm1CZxBjPHxq89m
QqTmxcn8r7ztwwHWxsxs8yPo9jxmninjyiDYQSipHXGyQxXb/+iaW+J3N5wd
9dHsd/s7OtUwh0tsgV4whzt7IoTUtIKmAkxRrTyb+rWcxb2YD/td1XYjCsoe
XeyBlZMacDqqQihhBTddi56+A1F9fLdrkyAoeMkpX/ERm3MyOVcWnl8O6zNg
3bWTdStMOpc4K+OqNW/IYXtw9aX+wqIhlE978+izkjh1JSNPzVwCf1Ntcm26
xDrtlK5sBA819lap9uT4tx1oE6stR6zA4TFy7muJ5NzRuKV9Rrps2jMHl1pH
GzhMAZ5/anFv4Ta/07XS8Etwwv1cBvirfJPxQ6aivRVrTXF9PtRKwMEBYnQW
i5yiJNNqYB/26gK6pcO7MuSU62tuQHevhvGqgOm6OozW1AAUP9Ix3NSgefQr
sV+q+5WEGAo5Vxbea/6p/3xBt0PBqZyHUbBi+YS3Cj8iIxmvW1VM3YOFxjgL
m+dCB75raIDSkCJ2KnT7iHsYKz1PGmd1QSagOWx+BDFxhy1bkH+olbP5WihK
+s+RHv4gQHTCguy/aCaDR2zgsP2Qf2RRsjcO+raF2zavppQa6MbOYGQZc1sd
eO9kLXUI099VqkA+0QKQZakZVWM2A551rX3J74wxtkMfVWEGjzuieMPjWfDw
965C1PAJqcML53/oFd7C581RjARmDyvLKBmYBqgb/iAaD9fjUZPE/rLhBQrC
XGqJrrLjBV4S/nRdj3G9EMBNvzp02IA9Nyfbkyyq8E2YJcAimt2Is0c2Pb9c
WKe17/zmsU2RAvAYRyaT+HwLWFGD6z8nLiVg5XOJt3qc7ZCkN5686gdza87p
AVe6SUjqMwpFARfBukP80paNoaNg2pYLV/lhWBe7N/ozoARvQpTn3Bc2B689
qqAt9s17padcwqT0SXzmDvxDfa+gNIWX4ycb3l/76XxQOZmBoyhy93wgdk/A
6lriLo5P3lTtPETJqpum57vzIPNB1Q7YmdQt09P+cCiBYpUKyt+8bx4aBRuL
pd6izFDtsM08RchQw+fMuYQQBEQWRzedS/YZD38QJnjhy02fpYvTLVWMuL9+
QCYuR9ZB6q9DSnnIf8UpFjLsuex9W8dRky/qEi10rOsz9w8RXXPdSgOefsqI
qi00EpLWHgISt0skOi4o9QmWVOfiTzBjiS/hulsxWiQvEqENDhjsNcrSRqbl
LakwOxY3Q3pt5L3tDc2oJdwrCTE4TezwgQhSoZ6vJEFqqOPVZivk7NaWtpQP
l9r47IIQn39RVUfdVW76u8Z6IpTYetPddLVMdE/BSkCAzSaJAevO3GPBnHiI
uSKJqHy02UMLSp7oZ+SkBDYnkATN5FZYOO3zJ/v4rafakwAfwnYBfRRhXpb+
uNWWoqalrY5rhGLbnECzC24XH7r+/pGG6/D48Uv3ClwR+8Ynlon+KdLXdCpd
y/sGqfyR5oRdKSbUxx/svJOZ7jFY0OaJiMkq4qlWbmib5NO6qTV+m5CE1cFs
jPebXOpQqAjabbiA/MMIMkD6ptMmDTMrzK7YxjrXaAWP/3CvlUnwgRCzl5Ts
H000wJhxTFziUSXfn4PRCKNFo6Tg1g7tgtEAX0MzIwOo/CJQcXIdObI1Pg98
lCsHH1RT2CaFD9h7lziAQ8Yzp7VmmMvVlCSzbEq9EBsVd7vS+Nu1Fiu4MqaE
2qO8T7iYdy+R5QmjNoYrvAsZR87F2TNe5VQOXR9NDkIEWHtMNcRXOfHMyshV
/cEwHfCKV0m/JiW1NrIkGxovsnWmCW9XtM7NXUjkbIsURsR9SWOfhp4NtM8A
YqI5hCStoBx2uN2Dl2OaD8Rm2hsauBkTWrZNYEPJePBFcTo1vs1cxWqEoPPj
XcwXKNGAlzbvnSJ7ixrGLMVDLHBHRdYwRwUk5BoaZOtAqqIlO5hN9XWZCxmr
skDES4q1f2oO4AYdP57qHg2aJGdTp31Avf/05vwzivK3I8pX0F7CAx9ZpSXw
YmvEI4En9cpWc4YrRw2OS+Q96fLIPho3WyjQhxZAWk+f40A5b9S+7jupjtpv
MiWu2GC1H94/fW99HtvkRBHkxCUCpUpSBVBy/PATMV+CUhMcQLRupmxFVVKd
3E2eYjwNf2KONi4BpogcJufEDqItbjfaMB1fxrp8pMy+9G2y5xodkcFQ5MYf
ppYln6e1KKflL/f9iT31MRZ30+5Kt4L1nLPqMBnadF7DyAC/qaKtevHzjpZQ
0M+sAgaZvvIfztMN86bpYQrJ4g5g7FnaoQid4kiQzu5bIlrCZq6zFGAm5aL1
wF+E/NGq4Z5IhVPQddRRzlS2xc7J+sZmG+GfHYkbMiaLEQGKVJXF2kptjbCF
lxHkhogL+RbJwYxwT4RwScG5EkJBBbJLhi26P7GdiFByY0TmLh18B/iVVfUV
kVgSfZsvbKzrLP/VzRed5fAe5J9/KluXRc6ExrOB60+5zQcmO88z822vBHih
B47wv6i79z8fNPCwyMcE90Iwavp4XfijQXGrhf58nvm9rbT6xQno9QEVBfxm
/QmLgrs2wXlMRfEh/bHwZW6zd65UqVA0Tm9xuT2tEA5kCGhil5ep/KJTy906
4CnvQIg920Mp77Fg8yXmOYiqGsk0c5SdKQVWKYa0n/rSZZPDoLqaom/PZavc
f6j7/bIC6t2toPuYD0Qf2k2HToy8OJPsrH6VOoaCMjCbyon18Brsf0g+a+Gd
4CyixdBpmSMwHgwlTW9Sy9MyiM1hqdkBQVCJcPKIr//vjkj9XmtEZoePE3NG
OvbSWwybUBuLDS2RNEH5DQDnhSO16BNlytWMzTxorScGIcNTSgY6YUqThYft
U4iK0ZXa/T/nKC/eLTqRvH+Tjrh315uq8ErOt+gTjCJpFta0o5ahowTPyzx6
OoABvVwMPGxrd6HVt682ZGsxIGPNN2EPApJgZzn+k2Q6tVQxzA0465cQ15YI
MRzs43nLUyuUSmvhxCCx9HK1CmzqNFbiQXIAGshBQ+Vp545ppTW7qnEoC96u
nQcBUjr1mRKZSpWG0tKmkEXYojO3kUm3vUlg3q5DuRBn2J9sZS+2oMPys7O4
BjI6DwiOHRbYC8POdCL1RgoPLn477XsfegohUa9qxJBJCZaUBDdPXuUQfmiI
iup0dl1BGwnBTbJQAgsJL4j/mc1FnDEsTo+BaR728LB0rD17PMFJcEn60Ika
ahsRkbl/9p5WQjPaPdAwe1CpOzVAi94oQzd8ZQ9Bjl6iQdmr3TEUijDBbjNY
LO68QuLIdvQENyY2ygFgq4iyQ2ARfoPzUxjhWCljK8XrOWMGBUZolrgRSKen
X0CdsZ0z8bQwsgstxv/hGkpfE0IA/fMQOgDPGhyOPkgp3axR9TLa1UZL1dkI
dXQwrKmyfNyn3azg5qE3S1xfBQICDHN1BYGczv41gqv3SsZP4gx85Fixe5BH
3tzBMacwmC2pB/7inUodsTRlT+GPenNRFaqzDIfeebGJAfu0h8SiFmeli4L9
4BAPDyaAKvNKVugkS3upe5n1s2mrpTr0/APKPQA14uCviGvsfuwpeSxAfh0G
SkZli5GBfqaEgsGRvzeQY+1sY9OcCW09B5EJb8F4eb1dHogVi2Mh5tNQXQhY
bO9wUTiPY8x4ZWcrnVCB8HYWACDaOTDxpbfApKOv4mXaf3Yyo7A46OahZ/Bv
z+9Klh6ui4+CQK3cfdEOD6Y9xflBkFHIVMTd63oT21AfLnRqsTvqDJrFs5Qk
jSGKF8Arvsc+V2YxU4bRYInAvquEBlYY6gbnz6IqLVWG/JNe1PeV9aoXr7l2
uq+CY37YtSGxTPP01y/Ak+6H9Y51ATIj351Ih0z3yf3EPd/bHMWBN0aXrGGC
ujNF1m2Upc7cFHY0tdaX976HiaEXJ+lT3b3jHCKeYOAVtieGfo16ZxT0y6YY
wxSBjn/NdfDUzZFjnC90oWHlJWFdtf+/cr8XBbKIkGvOE0sWJjZNkLiUVIh8
F0rmUVeFdDeN425JGyiJT4+4M/YUJvrWtGFEIMyFFMXyIw9zZJh87dZVgOJ8
CsznqX1d19/Qr4Vw6M5GTaDW3HTmijXy2sdN2Jp9BO7Kbqs2+6tBaQV7+leo
lgpj48EIUWgxq6KfEczCm/nZXxmnk9j7sni8Y3hMrzxUtOHzwZOKAA4EZDwm
Hl2XySAjmLgVh+eD6RjUExcoX9mlrcQuEZ0WrGUQ7pjWzCfURZZ5LDjmvL2I
Vao8Q8YXMraS7vd4mQnOT07F4jmkJIt1KkZhJ+8bLNccmSALhUgpDa1foxy1
FBklwN8RUJOtaiUwkKjgnbKAVfW5DhALuxwFlR48OWSNkpOaoi1JoA8Y93q9
nkSDZm44HMcuNHdgE1isXJ6/KIlCgqnMbNyqldiNJTrFhp4d5IX4MiFv3z8j
MgkNZAm78lo0P+43JxSZqrJJMiTbaCsUfZnv99a9KRlRyHCSbF2IsHTNa7ar
HchuoU3zg3OEKo5EiZUcWDFAAxifN8FvwEXGMwLqPR74XQNRdq3j+W2Mb0Er
u7KwP3akUvDG59NUmT54ll8x7OnNLgfJv6EUlS3zw0u/H9RJ19tAkiO3j1jT
4lxehO11jlpmXKYKffPNBU5Ns2p0wkI6Ri2WuXLFUN78L0Svcpzqj627XY51
mqN3TKBvVavw9lID7YuSAx0218QTljIEUEArHNhNAlBVU1pYJn0kabFLkFR8
FnR/mgp9DoYYM0ns9sSlGS5vkaadtoWnHuMRPQNb5Jo7esnYOxxOfhCja7Oo
NpggHmZ+KNXhlnOjo0Aj8Uhheg5fEv/xlCOR+/vTreo97I+emM61ZT1m8dal
Bk7Km8lte10TzaotFtWwjsrtVyobwMxtltswtpcWUwOJqanfwY7OCDn2LdT/
UhG8+R0UHHYrF6xSl+4TEz6uFBEz20RXIBHqbjrYI4xtOnyH6RCfVrAn7W7f
2rnMykdfioiANhSxObDnVcvDMzsoDBnO2S6tj//R3byv/nu79u1gBIQYl9sE
IfUR0wI4rYZQXFqfy48Cty1K3JM6QX94uVvgm6h/ORVCn7F0qkAcSdpYQxeA
+3KofCEYiy0su0yWwF4gZutqhgI2IbVXt7Mfkrff8E6l7zOhT7zwbwWQ+OPj
FvzzyPltY1fbv+onkhyPHEWYFZrl6V7AUU9mJq4dxnPD9Q9k+ErFyFBgQkzi
yhE1WfcQqsmu5VdSazEhM5Mgl/95rckVjuzffWWUtwCdQAv/7eKsrHFGSGa1
WbxeQ9f1tYHjTZC9AdUFPKlQhbPN3JfeKtM+/ceDMMifzboZJ4v4/qeow4iY
xxHSeu13CH2/w32d4gJKl9r1q5FPQzGANPdAyHnYeBxzRSs+SPp3Bquum7i1
c0cLuxRa+fGWeSnztVOkPP5mQcaEbzY8sj+Sep2UoJ+Gs1GmVG5BgGPjqkoP
gC5v+vCeD6G23SbFzTNt5lqb3HbjuvEYyiTEVg4vslAVJujxKIaJ7ZEUsVmY
XzCXbwbGr5hEm9sw9xgTjenJWV1ryfAdFsD5nv69xciNc6C3lQnxWPo1QXi9
E4EawLqmBfrkY0AkRQR0NFbhBWox5AmPgmLSvEG0bMPVjKrlkqEldYCPGmyF
uYNOP9kI9t7TNhVpvp4eHk4UyHa9JeFyP+RJMK9ce+Nc6dOaCA277OzXdp9/
17ApUzF4hnmt26PhzhRVdteKcDDLX4oeFuYiPPCqOavNWbSkpxYH40YXGeDi
12SLnCmy9dpSkaqSoa9p1+jZlllwuYTgxFI4+LRz8e/6CNA23WmZ9X6tkcaI
AO3dMhP2Ix7B10GphQxDWmYMnrJB4n4dOk51UoWYaztMxf+qS0RQ7OA5bvfL
KqPT3OZv8qYta34VnZmbM5UrSTtkDVzk18fixC25jFImA7UW10LlBbdr8qpU
wgKRqUAvGm/hdySTbwjOV4qrdDkQ2LO2j5ckOHvkQKkTA+klTpIs47ZdAcyy
vONVNKUbMES+HKc7tiDpNBbR3AqU7OoBhKPimHWI4duYql9UgTPHBhw5DMjb
3rn7f45YpblGGnaWoevYIBkWUEv2vIK1FrY0UZQHU6tQdOntyC4h7KDTatu9
QSE4xCT1oCXzaHbY7rp+wDmoTSAlas/EEWQuz737TsTxJU0188NV/eM5yv2G
8Mzor3pl42cIP52J0dHa/Wln6c3CTOXdPtAFqoppPOe8YMV7AFLJHl/x4lK1
RaSdb4SNyHtZTITkEuwmTgnClO8kN69AuEwoKT5XAk4bZT9sUJh3kz/kWjgc
ao9EwfVejge9096aw7ed52s7KDb+PEisE108ac9EN8PEuX1G7ozIin773DbP
/GaJwWTJN4qb9+zmnqxrXFk67pVtSbliT2+cK9fr99jtuz2GKgA9AyUrLS6/
Yfny/1rCj8LvviKa2PEDCyyiMZ+zN2JZB1NxXL5EHJ4fM1fg1cKochP+08mO
5Gv3LZyIr4rlDki3PSz4kQ38Fi2RQCzzTlnpsmEWki4vZ4NzKxQ+aPAmu8rH
UJWBrHrGjKVFjSnHkq3XdGwQDZqZHtVMmlmuucNkZJfSZwMPq/BeGjc09/Zp
nED0Co3AUZs/8tis3CQiYi4oVb7MqpPovqwsPfxmNmZbZowLMCc2NygpZwWS
ClwC6IJnUXWBTJG0e4t6oSZ8sU9n5kRKYVrhQrcg1OeXqG4Z0Y3sxqqv5hlR
R4W02a2vF/RQZgJNPTRl7Ok4meRIdsv6dfR+a6vQTCbyV1f0JgfX0SdDceHJ
pYbFwThY9gEhhHPGQfNCazbj9SW/HMeznqhs2PWmyLVO4KHtSWbH+xukqhH+
PkzA9QFi109c66ZVyb8Z+0VsG41BYsrkfvWB9WuhYUQfNix5X3kTzcL1xhoe
Cf4T6viIAMYQusrPjlMx8CIec7Ab9QZUZGws/Qh54dOIfFEAcPuEcKBYi9SZ
x4w78lBeJZgERjEWx+yOXeviWj+QNbg1QMa3/nFu0iGZYN0iZMXDUmnaWuFb
8Y/1U67gJtKS7jX6+2Ep2q7aqNsaMnbey34cJENfFrYloOiGLG2a68Z39Nm9
9hVAl/D1uUhG6jPnB/2LFVEPfqJgLEdrs8tl9KQ52mwudIuQdLRLbwle6JzR
dYIdO4C4zvzxqdkKUboNir0lk7bYV669OJZHfhjMmOeVVhShGU106mXL5ICG
MkmvYtPGfcr3Tihl/i9sDesW/b8P9N9x42M/v7FAD9Aq5JCPBRQBOVDHpffh
hpS9jifAfYOTY2Xp9FRLANofw2+cs1evUqgerd46CvpexEjrywx2ojk9yOtq
hs5EME3+EfIgg6iJw+VbQeeEyMDm9ZyYeQufBuhhobs5JVelWVNNn11W0SUQ
iCGl2t8/0OTo2MwpFMy6ywWMNLhD8Txf/mQatdh7HkiaWo9FXGtPiF0JuFQj
31ToRJ0VC88NcMgGZJrzPbD9Fwx545p6C+FqjFB5nrRO/tDKQW2COD+pSpXL
tOpfrT69tdaAKrAIU2QgWI5R6LyDOVrWBFnPuoReRV6bmB072K5VLORCM7/A
+UA56q7QWjYidleW9ChOv4nhHwaZr6BGg2KzCnhIOzfOecLYVLo95Xac4dOq
34fHYrA27+kFif0Rj0mJuyt7GQ2EO5UfDg21DE33/AtN/xu3JJZlP++TtXpE
xK5XWrffpiPSDc4ftqdpoWecZdl3R2ggtHKKSAyGapf88dN3PMEbZxGBoHHt
rIPfnA/aNCYttX3G2VPb8OQkLeSQDPzvt4OHbNbTr+ocaVHsEWfCn0H7ZuIe
fR8QNYvbiCzSZkba5FUAYGRHdxBNAPPyzoNZCatvcLIR+9JVMux8Ju5gICJs
cIImzeRi8bPJ0B0enWky/fOHu7Orcyc3ZnSIoOzowOmyrpj+n0TPTVp/JTE/
iJuZDN9XFTJWEtaK6X53DaBlIw3iDmgI7yzFgWgwU/5ADoHhLjeuKd+EqJFO
ckGrmwk3C1CZOFzc0h/NSfZ+cEDvnf/Vwa/T6IKhnhyDHwPwGdVEkLxRxNrM
qHk8ZT7kZFInU1erFBdHAU/FaYS/dFfdeML3b8gAc6fyDTel6ZbL9N8ySULG
HJlvmEmAXfXdjt3Dwc72eG9nf/SoiMdb8biMy/5wgTimuArXbHg064gDYl9I
W8NUBODX81CJ3zdALfHW+ay1en/k1ld1IRubJjfv9blcvRJcAjzOanAsgBZ+
+BvFH9An60MIxAMha54cIGRbKra1U6QKwqHPW4QtyZrdHMOh2lvbAsIYWEcr
cwXeX59goBiFps0uVCeErIuYyThNPO6dbpJfz5bG5qJYnDZ488ZNQJ/7aV5F
SjUB+p/Db4GXlCiWpg8IEZyIaHtm0pfMM5l4vZo73jP6iWu4mcUugSW1TU+s
1dTzn0VmWwlGmTfoYua0Jmha5wIOIVi1fmHOOLgKPgKnwKf062SshhRIheGx
xp8urX1d35qHc8F9elVGxMRheKQoN7Kx7aeCNwePdrftYjNSZNPXe2z+tU7a
3+6c1mu6457aDcl6UgGJaFs2UEPC7CVwBPa7wA4pvg8nMlUigeDE2zeLv+Z7
munV2V1A9sMSqAUYSEg3sqrI2qDmCLYoxQYp6pLOsuEI2oHi1A3m3Uvc2CNy
Y2WuFZUhlpBW9h6Rv/hC4widJUJNWRhqwXKIhgRC+rzNWGc1KplBxZl8F4Kq
t+mj5cub7IYqR6HbzYROz2jcH0b0LfGW7JLSudgm/2pzxAFKF0u4Oq71BgE5
L0u0La2AT1VIaHkXNuASII4k/mYrHlkQuZ2EPRbEhNbBe0Z+zBiW5yXYwzzE
mrwBetyGgBUxr/iOXc93GLiAqEvco0y8FTefimVRJPrOrpz5CUEEryfyR1ls
IiamTbzcOM1+O/duS7J0i+m6p7MrAhGLyfd4I/epzTVn9k4rrR/bxYWa1QFt
EhGSI0rpbHh3Q1HdYA437qsaMssNjFVgBVBmwRphJR6ZTHE1ZeSB9TYEhOTE
OQE1HHzxN55yrj18oEc/6izE64D5At2DPdy7iv5F7Rjbiow4gEtKL/2wRJ3s
84Cus+/01rrUaLB5OHEEo9tdudMTnplZ4E9ZFiSo5i8NXWDKl5nzATLHmrp/
VrLvxm4mF/7zRyET/QQvyVT6QLBmIkDBHXfxUoF4apMDfuLlyh6NSq4dO6uS
9lSofK46muyUiEj8XuyFsM+7CFHe76OvZ7HfPi1wp09+F2sq28oU8wsTM7kr
2/Jw4niKnG42G7CDRnAGO26CD8d/R+6UobjRpxPvpHV49cOp+G1w8YKdxnT1
yGAJgW9fCN8UAmYwqXRbwGxNe4XEmupgYS65HV+lLeHfrHz4L9I8DMfUxQwZ
AURFuOqyHq8gg4xuCGcvqHPo9fO0ZGkn+i3hC5kVPJrx1w6cr+/TXO6xZg5R
RqQWHdeRu4UHeVrgAFqnr3j8f4sS/jd6/PpvYmCHCLPbke+N2zKVQIQlasMr
lgOO6MuU3BlcBWPV+uSioiv3VdZLYuJSYvSFpJKpaMpL/6qP4eJteqjY9MLQ
O6zUuNBkbkSyLqgLeqQVCeNkkzVGuMmbu9AAUMVh3WVCrRoPMTsPWiUBizzk
VedChk0vXOywkmNmWCzYI12ajGdu/Vt4xmhysM8muRwxa0/+LIpAI/dbWNrZ
4uJhxyO16R+SGW3NBOB7EJAURqQ+Oo3LZb6JSkhoCeDWSqRwsByTVfVZr0UQ
IzTE0SlAjLNOtaVpj4MfLqCAFYXunxjgAXsdEQEFSfi0bC1MozMU7mf7/OQ9
LJEdjRf2ibnGS7ToMj6FjOMPwsGkBot2aOvM8cQikuoToDQsK/jSnqu29DGV
bb1nccFf1hhJJuHhRJj34RJHW+LgYIQ6dNs6vAi1olgfM8Oakfi2J5gwnUG+
iH0sk8cXtO93hzRt40rfB2maXJQ/MfPfX/5wTlETfSXKcposmDSVBhHVE60H
m59FZNOEsp887lhSCBIJKtUuAsM3LhWAMZYktENbH/SD5UrhfdyShycFjtqB
DsjyMwVGwv5+Xauz9JqeG+g7/4AJBoRj+WlB74rRYiXoWXzhtlcq1ThKfq9C
orSt+eyv1waSRlx+VyHkgk0WNpUFtf0BxOYNfwZJazsckhZ9nNeI2yvQgSBC
5lBrLev75xZTbfuTC8a1TIDfsuM9xHs/oHFfMwzSW2sBrtJ+lzHq6dAcRdGC
ggLVIM7pjORETXyTE1eaznHHUlhULtNQlnBKcWM0AVkWQDnZvf3tn0KTNk0V
niLgAN/1E7DxWPBu56vhq89zs1ZXVijNUH1ONaaO70ehFvp/Gislmgor4D29
rDV/dqw9ykEYuzQ63EdgVz9Kclps/8f4hYVgEo69Ro1AXOETMxaofbc/YmBB
0belgkXuNWhkHgDT1LHJctu9tdAm9oytEY5avyIzP1k/RzfKj0pwHHuZ6En5
w/SQ3FGTqzVd58FwE+N/06DQ3bbcEd5pz87f136Gw54ndY94LMcLgpW7brSM
0LRBfeqJm0TdA6e3x74r/6U/dsq78ThwcS9unD+v/Xcws8xbmLSGCLWatluK
kUN9mado7BXFwOYDxDu//LQTDYB+lNhitP4hgKStxNvpmHRrwgG5U1WbExWO
UZZS6/WiphoK+/VMCWMLLxpOEK+Ll2T0jekRaSlSwcZYPxt7G30Ffo0kBzgG
9cKGDb6YGPWWWXj4nnVpakNOK2x/VYHsu9x8UHGpfgmN3hQfX0IeuH4Tl0ci
9JIw91onsRZNRQptmkd3THmZapa1XTSXoMXLAipX0cdYkvyr2hT8mfju04oh
s1wUOw4t5apRyJ0qfuFDf7Y8PB1ogGRl4uLFI2NspxXgIuGEt1AizUPE5dXI
Aa2lQ+sK/zQIffusssOb5ySlyuOiTMeqbEhhD0qoM6DMcMSy+SlVze1lV01J
fKhPYW/2pfJO9ouW/uDfi7i62tH5L0S1nMroHE7Nr+xjup7gFTq1PhOsCM13
/W227QmLTXvYeVxUdsaJmFN5JOV1HzMbJd/FPQ6T3RewEcxMvOACSO4iqP0H
jVc5HF/woAYe358y8ENlpCFSSWDZn6NmR/s7oSmAFZoJCEVtHPXoj2kggKkl
hEynmeoh1FE5UsIkUhTtvXu0bSYw6kVm01QHIJSuT6I1E3sySdpZEkQJe0hp
/cvR9nQitLHHRa1wev0wVui+8ssftsapgR20vCfFpcvRDHlWIHXEq145GE1t
FcBqw3MXKqT7M+fLbVQSzRhk4xUacLhCzn+dN/FkCw6V74Q2GygjHO8goctv
WLiF3May3LUlwkYULUoBYwxNneL84Lw3VZK0m9GfC2S2RKcWgjoyyKf+WtWe
qFlPlExGl6aH+0Bud3D/zPW7AwBy+HpmmCcKuOqzKV+3DvM3g/VrBRDEypEo
4ZmxaeRrs4/Uu0uQCoVRWvy/yhlq5uzrQHObfgJQ+uSLqGBDTrbXXwuhFFqX
QoRm2g8UjZKJTM1iqtgrczxgeZRVDE7k31QOBv+w2cBs5Ufg5euo3dh1g1yV
PUxS8Dl7zm6WqYCav13pnIZk4mYfk2Ffr8kOMh7joziKGl7m4XNdNNxCZxvb
P+6Pn3FRc/WHEbPc4o+WuxxH0W2jk5GC5C2+Ni+wT6P65pP1RyrAi2pf/ntK
1eDFS7QthOdrV29uvW9P/G6Rii9K8n/wkXfK6DfjWv9h6jCTV3sjm8ecjUX/
wNVxIqkIuM5nORnBtkc8hfj0Cv0tndT6htJD9edoq3cTVWpdv7U4CibI40mk
IkTMNk+bXfOeb9VtB7n+SaijfDIR75bEhI7rfvbw14343WeQ2WWz5MVvpWVa
V7xQ0jrfVa5c2/ZbaHWZl71PAkuj7+UfNnJsIlq/s2+tekJ2V7Cbkk6EN21t
vnsA7svGbuFyarPZirZ8Okh1sRnyBRRYGYIyrEMTOYwDYioDfnHN8VLBTacR
0PSv7TtHKho31VabxBt4ci2Y9e/VaBPi7vIO/jzU6Lc+Rpi1FGiSo2wXSWtb
+Z5y8kJ3QmXW+YPrcvYs4U48snELPe2YcqXL45bkuY/VXNm1Q0rC//wu/55g
Lk1GMK1j15KSOGUFMEwgvwNleI46/CiwuIsK7kC99qgw+tdyqizZn0YKb8Oy
fh3YAoBCM4qPCrC/9n7OBf1Fa5WS8gIF3z/YHmR4Be+FJY1XVu4mh4N8kt56
fybFnIsiy1jD+oNYw56JHBZo2rmRnAL/K5cyvCH8GQH8erk9edrfExHQndzH
LZdan0CUfYZxMADftD77pxEnJ2aAxb0+P9X1BiavyXytMFE9ofg2l1/P60ho
BIk0Ar9MnG5U2+9Kw7lCIxdVhLE8Ue4fZC6mU46WUrpsXeFIs/j1HXIGIha1
2ZJNggRWdHQoYbpi8k8EnvwO5DBJeEoH122TqmvPskWmvypS5dF4FaSGmZTw
6++9zCrE7bIvnqScv/eqFDqiRk7n7CFGZdj6QGZs/OiFGaUsEWEnfXsDP3PP
Knq2Ws6c29xPjIa8wFEYIwWHN92UYyWpeSNkjujrzfoKE4a3nq8/esKnc4aD
wPPcuh1JTPdB9OFZPuzRnnxbjn0DfU1qC3rqQri04I3J5E+ycNu+/XuOLsIY
mgU4XKhiEjBvtQWtuDGW0HKiTzmVEDkoUf47nBSJyX3gX06PVOSYEzux5E68
p778DcX+MIJFhuazyc4iCiFwafGX2y0+qYUIqyGS8TksjPk8yfUlbuyM7ycc
wtzM/veK+c8Hznjwm71i2n1czQPaRLErVir0m6nkB+VaZRw62iRFxz9Ndr++
J+0o+blmRa8tr6qRkyaNnRAqh8+bZt9nPNcRbTdC7RIEPCWpOk9CUlpew7kB
EZnUr73dIsmlHQKOiQh6LHrYLdOadGPyNzP2i+294LnZ7LzZAAQl+fJxNM/h
jfS1xX8H2jAEMG8Dhq5hijg/E7DCS7KmSz3qNTQBwD/N3s4z+OJZ3+IkBixB
GOVgTE6HaFpuIRsnecnVCVavQXL2b46yJumAu/P+ypsxlXnQFnliGzocPHHP
qPVOwBVNPs7AZH9r4Ram+b7RuLbWz8e+Hr/08P7rqjEQTlRbAh28IZ5zO3OP
G0cLofkGDLpMTCh2SUz9LkDYIyvsDKy6T5RDpuRRoyF+4rlbK7YuOmpWosFC
WA/sQrkBrPl03FOKsejPkbLEpubVHpeLXbPHrXMBKx8ApLkpH8JiSbWChcs9
wHXBDRHxloqFDXZTb5SnqmPmludxP7qmTXGLpD5ssOQWhSzOJmzVNtQMwCws
ssT8wXHUk4jB1/wD3+dfdiqDkZRggLU7y9wN5BviVdal+qn3/QIjre86fmnJ
66GnxMu9xmg1kCkrUkq42TzNi7yn2IvnRZmDTFRfPm7f0p8KiQ+yCHe5Y1DK
6rWeoba+4kKQWWpAAs32bst1KUkOY/fjJGuO8nf0AC+31M2mA2vbH7/ntztk
jTDFn8tKKXD/wtcO/Y60GriWhMnXWuH8Ve18U4yJb1MhOPQS3Bj8BpVOWtEh
k3777ju8NO+Lro45iXdCUPI+yWdAOKMSjB1uAkF6668+rm8IQI8P+/wVKJzh
XYFJjhC9lSDEa8P8fugEVjrUuJviGDnBTuEeRAQMDznFVOFasBQhC3od9Fs2
LleRbi18SpRVap3NjZ1JvO2Uh5txYT4dbwCZ5SAonAil7HGbcTlYenzk6gyk
1rv5RDH6/T0dulYfUakc8WBNl1dqLxVEjhNjA5ryA4Wj1mUK3DeoT1i/SszE
kMD28d8SVgtV8RWX8Q3nLgHFD0GQk+hYdvwZ/AyQAgdYFvwbHydwSXniADT2
tkib8Ncs0Fifvg3nnaIpGEm4xWW/Hx+MrRWdaDI4VOS4stzdnNXJ7GbwNZSS
8oIfdozWESe1Lo6XbuPUQM3f7WFBHmOl5R0jy/TdVeTEu8WYY+Y3zJxpYuE/
J0fOj8aTEdyZJVeUVJvDZcE8A+IqwZTnSuk26CFgN4Gl65npT2nRM9ONO5t8
MCtyGVCPe6wS9pgpL/8UkZy4qw7hv3iAh15xAqzInkmRl7B1adeG/vJuEohV
1Tzgiwg5frB6nUJjGd3A+oYzZNNUAbawXtPomEd+asgtCFJLtJwYusie5uoN
69nRs+zOIraoKUFeRUzBhL8IYhC43lGVdu/HJF0IL6zyCBBd4JKyYXbTtDri
cOfG0YAtv0gj/fVbtPZmPquGtJzfrc5pg5vDHVSBYfkJqYZHiNFU38jg+vmZ
U/hsfOGHASN/VIRF9W0pH/fCDXU2UgFMXfzNH9uqcqFuSJKU9izJlX17g1Cb
aH/5wlkeX6DRUd7WwikjSj9IYOQPSAVlOm15z9kJnsbUnqkMoawIM2bBzAys
3sTQKHplUPrWwiS4iJHoyp4CbRE88z/0PRBWjtvkUHDl1l7YRcaEgK0g349q
JpUBZzu9RmT7FFLnuGmv9OT1WX6zMft9Vp92d5MAFleEw1i9BSg6HWTbxB6e
lgEOblPq2AaQWHlu/qPNH790dAVvAiWDLC3SPu2jTiREmEiO517HAYRfxh1Q
65ClLBFc6PB05mpjJevo20nmIKXouhdnW3Opx2++a5ScpH36elXecrj5GXOT
uWAORgbyyoTM7ArF42syPqHIOUZaFqYrbttoFw0XG7DEsXmS+xA9bP9kr8u9
/1Vx5cjsGMhImGi+yItbjWfaPOWt2odcyW0puy0tTc73FxAg9uGD4f9iNnny
TCXrAKsfNCBEPG6t6WNnt4d15emE+LvbDix30T5Mldcs7mGQDUBOiJLOUzUk
v4ah039t0DlUR1yP0vhNQLzeZhPQlWnFssEyTlezRHsx+1u0NppPk07uG2WS
g2iU+qCLMd5R0EQmNBRxx+Nqhhyc2FoJYarZlSrk6FnZLZ1LCSLzeSJYwuz+
jqBa6U0SloX0p1zTv1scNfyKpsuJvlavaJ0/7BS0eTFy9YZt0rAlQ8V8OW0k
Bx8T2K4Jzk9pPbZ87c1JphDo767bZTDO9ITCAShJ9cZqATmGU/jo1GwtO9kq
eqtc/+a2MKCU5OezXrtpemF70eohON8be7tJ3f3XCzegl12uWLt0GtuoXCUY
yR9l8m6H6lxwM/rJpnUw8s4L2jauuM+gS6GlVgtPCywVcwJf1Hyp7lKmD6HG
MqSjVMIAnG9FZ40b0x7DJ+mhiw1C6oqlvfLDCiWbdJQmZKGdgcoiwiHhl4ef
jJ9lLW3FJuxljyVF16gug2iqmDyqwlvQohca8YAm+whI2u+C5+ao1nAL7fFX
r7V6t1EXEBmvcmrsrMKuzFd+oYi8gXlslKrS5geYWtzdUU2+1neHjKOmyWaz
KPfgDPG567iuRyYeSeIl1m6FARWXKbBpGGvhn7pZnIIMBRccKQ7ispmD8GhL
vADzexDtpC2ZniAxqNXIiB8S/9XyNIMPkbtVo4eDeUHZx3bj2FWsGi2XjZLr
JMGmcKV+ZiXJejJVszWA9e0Mn9jA3aXd21GcB1qp7aDSyKvEsUvDvmswj9Et
8x8ZuWoCR4/HkLq18Lo144o3yP24miFSo+y9xSqssQAYqeSwDnwZkt+dwYn1
6Kph+XVrcEr1oALcMMPHtDlVBrbuTWaDLGW7TYcfETTV7c0tspmEEAPJElPH
29Rz/3tlx4XBV1SatH6uThVTIy3k2Kfgf73q7pyVU7mzX/E2uBtcINIaKjsl
MSODjGqK2lvfTEWa/ZOIJt4XEmcWuck52zY7rDHTvv3xXr8EGPD2yGty1fAA
Z1Gu/Qc5oARr/cP+pSblPEGWy07h1wU+3kk15DWpYK+0YJDmpMAoAl4+Eg2P
fE0v5PF9Na6izVGJp82/H9UTAda9bjpKVojwa9K6twr3vmaDwRD57SJjZn1A
qGdd668LY9dzUQ1DXSfS+OmmG/L902M7nKiHHyOJQEyX9b4yjYEBSgR9pjTj
pcDvkVJuKT+V1e6m8cgkbccLAJtY5niBMz5x6cnHpKOExITJt9aYyYAYWqee
IpoAwO/N78FpqYycZifwSy3jQu79MwAdI7+aa9TndyouCuvrwTkcgGlU+3hS
CreTgH0NmfpikPXyZkz5eR7Y9ks24PnyF7nB43eCc5rnfouqRSZ2tYlQEv1K
wXu6a2lpfnl+iNRQ/4gUcj8m7tDNX1a29dQ1cceT1qbXFzALv5pM8w8PfRs3
8XLE0hG4S6jtOAbtlcAANOKDgim+eFuZ9D84+euC7Viz8FzalP70h2p+TEz4
a8yNSjKlENDixA5lH/zlXjFKGT6a2NB+wq9aGvDMDoOLYIvJlSmW1V0u+G3G
a8w8A97uR2Kye+dlm+WcIzCGjNRcX/YSQyjTn01f4NGc84E7K3NCTbuEv4zU
Vd0Efa/1b23Q88IA4Q43HQTF3JP2mhhMLmGeqSK64R5/pEUI/2MLht1OlwqP
iJeqHi6oS3s/DsWWKc6bE1oTHmc00WBb5CJ0ykPvbpgCki+/wFDNpwZUp7aL
/YH8vvsbXI+YydELNoajg9Kw6l114eDEkWBxdg1SfGhC3kPZQep6SCt/7B0K
bgzNpHff/jkBzK3x5wJWuNF684aQbHSeh7Hx45WXsX5rT3Ve/FFiwjgzsTVr
Ejwm7sDQCfmIjIf10uLgpqfqiI9lr8Vap1DoPStI1qsSwxpIM+jv6dJ4IskQ
Licaa4kCfCGYkFFR+AgC12VKro7IKPoFkNtc3b+8hxG850uGQUNYLzZCgeFs
mSbrwLmU8YFUleX+k3E5ofoXVUBDNo38F1CBri03HMZ4ZazFMYFmGHug+d+/
x5kjUt0H+O1K0XOYAJNfnmZMuQC0EL1SaPI9SCmfMvggalCPYNvLE7AVikjr
Hk8l/ANYKyw0e3Ozs3F1aqpfJtlwUeaYrXHO+uQHSpQ21vvtrvSoXGVk+xKm
eNERx+vym4AEAX2JPkU//a4TdKXrmd6Mra8rKi1Z3k+J7SEiI/X5yTZvLA/k
8FC+Su31FXMqrs6T6cXws/sL0TCUTuz11aSVLnW0q+JB013wHtTGxkE5sU39
SFqha+njeGlKYR+rv8uOzMPAmd/MabPuL1SqmEryogYw8fuUP8AD+2c9ynz+
aQvxI+ef9PxVndL3tvE9rDOwFay2ZjweuIvSSneA7/Gj3ZkPbKih/UGVlhp/
3O9B00/A3tPXWqHO3rOw0fvachKd/h8toopc6Mx06bTKZFFbwfr5iBDK9MFG
jKmmPZmgDNBy+wv0xaznjOqHqFjae88s6yl90xep14C9PG1P5+8UKtduoBV7
CgY5Ia2zSBXjovOkAEYAhjoG+AtnzYZCN18hQViLXzNW5TB2sinV4jDjC+wb
C8C/hIa5l6a0iwBQ8C2TDQ6pFQtSqh90tte9r0bdiSgEo51ktR1Cm/U+wCwJ
uhakjk/zRRDjkCUEmllYeErwRQL3YjUG1dDHejm2nnyb7UQO4d1uhW7S8v21
zXqBhewuL5NZlSFARZzWOrRoX2cYzgj3te/W2CGvipgu6gYxy9BpIFd0Qrco
y2pGk1XMlCPGVKb83GcZ9/l96Qy7Xw94Tb2/YHPIyeV01tpaWOmo9wU5S7xh
7rIgDwbsOigv0JtWmKghTiq1lwy71fopUrm9zlRGZt2O9wWphwRt5owprywR
ZHsLiw3SBZKkc4Hyq0u587oc7lyBcdtRn2P3/CbH8p87+BXO1aXAr/fi9LGU
Tv2kqF6gNXicCFHsaM/FSihRCb1nHHopbXE6lUN8uVDepk2pwNKmh0RP5V5y
7xybNjVPmIbxNyprGXLo8CYdAcLMfLpm8I+P5lBAHhC56r+SSpa+XNyfQKnQ
M0gCOv+izCnjDzovgbLO1SsiOiJYdbkEohNJI4V7x5wI5eSQO2CWBiBmrR/o
TegJ6I6RS26BWlQfksfqOtDJgVZkWHedrlg9eVQcqb8/P2OpPafd/fue8i4m
kjCls4oxXcBqgGOgJZJF3Yz3BHsu+ZvKjGBkJTGOCATbj4uS1QoreqhQK+pH
OpBl4dYLHkBqCJZ/FPLdMO0Y4RNGPX4AmRIs6m21NQTFLjmF6Pv1FNXVOIAL
IfWBFllKt2RLXosoi3UEewSSQJPSypoYc+YVd9m7MliNZgoz2/dGGWsYrFiZ
lnF698bv08uN7zs0fG6zoDLT6OHatNZE8MausPmGIl3ULkbBtWogk/JbUbYN
WaIScCIaG2gNI4bV+uZAKVIzSiL6by8U7uMlZXxND8ZRHDCAHi4gJIYZi4xr
hCUvCKG7xhZaw1sb6qisUt8xVIQe1RzpWFJDQNDduBDJhUWzL/QdY1FOs0w2
74tA8Yk7BytDIBDTiLvHcgoAS/xfsH/H2bIwvA2/d2nZ1EDLvr+lIaLELLQH
Xjx/A18xVA7MJLK7Au9FWdpsoyVpacopgw1xEdNobetnaLta3oc80o0HdVlU
hmJ0EERBbUe8EdioO/+nWYOOTZCHsvYQ6Rrg3QRGbxogRGMiFN5EgS/7TsDS
Ewnd1wLWbelv5wMPrgGpxqXHlFsKonKXd19BQzWSZPVD33q5bqZ0aKcXuhtz
7o3WX4byM2qpby3CpyMK6Zr7/1JkCzN/7TQvD8J0bRZKJ83vFiTW43jWYkJC
58inhPWpCqM7Mun36bp7qztETy7WDAh7nzezMVztXIFaDEWALbzOC1elo9eo
8ThRlt/Yi/KES6V6YjzZU1diEKIrJagItTWrAGt1FkU5EwJhzt7wxGqEK+OY
9Ieq3oMbCMaNsG1R49CkniydaIYsX8oHCF5kF6Ny1hA7A1IluAH++D1EDVVY
nUYNJvhJepMpB03xyB/EaFbx4yAOGB981rXCUYl+krJoxlQyjr5UEP7bqoZS
Ux37QyiRCf/YimuGE1hjfSrSG0te8wVw+EU8+xwVRsTCjBGEwDa4fgtCKMX5
JK8Bnvjr5cGpQCfof50TQ5l4L1NuXcoZBbqE3bzqVmKY3qW3Rc2BeJIPIJwM
Z4pp9wb5W6AXDexDSEYTyB6hQTb+wgGhQzdPnclPoc7gp7gQVtxyDlC+mQ6g
AHxOWsorMJFcWqLddlxFXIeIy8CxLYq8FUyOCqzZpr6PpLR0+cLFyWabePF6
nOcLutgwWjqJC1US5hfAzqM+DD0kQU6khh+s9vkDxwnjfowx6r8dUfgh3pNO
8/9/r6iKlz5lTE8nIJ2IAdwKEv81mSUirNt2NHZMHt1r+995AUpQgKi5fnd0
v5RTZJaOt36QMjkNorr8SV7wNp6osuALLm8pdN9wDyGrj4VrJT2e+oBY7zhu
bCyFOIDXYYG/eLtSPWxNrhUYegZlZomqM+nnoETKw77+x0XaXqWwyOEpeU41
VWKFLo1xjUT3hVZ8T7OyWA6nBgMlydlyMDCCZQduOZLe41WTDgUfzUDcCvqK
IDYX/4LaUnl0exC3IW9TBqmfzbU3hlhnOE1vLiDZIft3KcOKyR2vVjGtjZ8/
ZT2luzjXT3DqPOh7TJu6/XNzkYPSefQfymbsFlcOw6yBRlua+umFCuhmip2K
URc1/maN26LK6CPxAaDn9FHaucYpKPtkQVfkqejlVFqV1SDEe1S8oxR+mieu
P5pjoKKMjyE39ypdp30ZAaxNQrCgtmYQK0Ry48/J8ANOSDacVE10/PFQ5XfK
QnNu+13FYeWCsFeYu3rdP4v7oSYjNG+NmIhe/Ug3yIhUoMwduDNLWmeOvAVT
IEcGthM5djUCd8leelCCH+H1RRJ+rH0JkvU4W2gUa7DEJBg8fxBscRhIq7JP
N6vn03MJS/BoOFw9LlQwbIZxhKTQWM7Smg1F/33S7ki7P+qUJBBufR0GXzYr
UzjPS9GJ6R8WCK+RA9XDi2KryWDQUE74Jz73fJtJnjCwdxsoY5VVmPNzrayV
ghnSZPQ1bXFtcPe+nsO4Nii47mG+PbSFLi/CGeJsfc4kRAwd7GRgLNbXwJxV
tA9uOKQQo7ygindkmLPezikXG3wU8V8EEQVArckyITcnX5CmYK4/HK/bJTkz
rMD4CkGmcstw119jzDOVW/X8BUImhoEiKNQBrFpXvOT5fsWSQQqXORLJ+ESJ
ghddXEGbAajMmw9peFZ+6xMkD+lizh4VVqIXTiCTUHj2UfZMLYwML7SqxUm4
Jky4brTJjsGgEma7wrlzSCOqkiCIG8/eOtpc9OS5iZrU3LQyDKRXbYmpWA9E
9jsTi1YoPUo6suMgs28Hcif3roZ8L3rmrYb2CpddYXL+F5gpvLOGuAGzgyUv
TqtkGNbAKH8eVgJDf8jUxBebswhO1yX7uiaCDsUYWo4Ge1VvEbnvf1SxbU1d
bg7OcHfLzGe97KWTsIJhqL1dTbFFt+wkm2TV5moyvYeKfN88dVTRaTVVUmrQ
+vFBBs0fkyxXKerxthzm82cB+hBgtnrUQSObyqnBOmKweiEZTcA58IH/c4va
CMcHEkB4KOvplnV9s/Ku4TAAdK/NsKhGE8NQLUHcgRphLbnzUkuRmspaNVzQ
setwNIki4m9K24QIu7u18xl72FGIvBTCU0n2mFOPvM/S78DnNrborJDFC9WT
ysEJ9LPE5VIA9VjOdC7lj0QMvAy+quVczn61qUmAWPCV6XGfFeQq/EtxYEP4
945idOOwZ32gTE2RMLBQlkifkqrMNFUK7iFbiILeHAOItQWm/B1iY+CXlCmR
Q7AY0bzGK7K+CM8FK7rNgcwzyb6Qqk51GC5K3VGNRXbzo8Yjcusd4QnY7Nv9
xPOjx9RkKH6TBFqLiz5NLVe+r3NHDmTUD8tjKT2UrdTWDYH/qRflxHvNcrY0
Ak7IyuT33SWAahhVKjatAL9NgEY+EAaWcNsRtTSXa2mAKj5VEGDpyTcexfiT
FF7djA6vewx+kneXCauhRRBaI/WnBDvJOfEqiL8FYYWU7JJdhS1Xxropn9W5
HpjE9kow5nbI8CQr3TrvU/nIOcqYiWasJt/iJP/anHIXwpIrPOy4AA3fdgOO
oiVwL7tXJRxRLd0U1ZPq/RqruaVaLYeCtJGuYFup2ZeVY3O3oU5tMZnyJJno
9+Gx9VwjfJbMWWYHMaBAAgrp/Ps0dY2RbUHm0/zzJEYI8zZym0OmFs0nPMJV
GKp4IDssTB6jjksrqcKjJSIFJImLMOwcCQAFYqx8JmsoAoremuLmSFTirBWv
NMtNv4y6MqbzaBR/EWQ3TwDT8HXKQk8VgPMmucZgb8dh5Df8Ikef6TkCVopG
CGS22XnGENCI2vbx57l9ePjFPHVEzibHKtdSvJvv7TiXJn8uuEzuXa+ZsXdF
ahpm4+3wIN/P64525lrkle4DD563TH36QaEtjZX7sDTJi4bO+GsWP2jQzJPg
kgZoZemnF9onYgFSafeR6+3u8YP6xmmIOW7FwQ/pqW/xLDdAUk85XH0aVg+a
o+qcwUeWzA+g48XUjjBRuZmUl6ni+Lgf5JYZGSxvgGhoidJrbLe6OBMUCJwx
1b0bh56RZ1uvpJVMVT2+WmuMR9ZVjC4vCxMOrLC1DnPqKCGanqj0BWR5cyPR
2fNViwbFAF21MRCzXZSKo1niTMibvjIsN0a9n4Cy/qCF5sT5bUIrVADYHNaj
hK4dmuF5Woyo0bk65HoPwnw0da+6UsURbEia0CQPdoztHjCMg27wXveCPuSP
m1UZy3SJI29Xz4LRuWpcxwuRmPNLn3rKlHd+QsIBn24azuWDeJLTohLyC2pI
dwecpMnmc0WqjEUtA8P69Wf3ytq8Ivqt/3amQ2eS1RRaKyQ5t4fI82jjPt5z
XpEJVeBLexJ0FEXHKE8XljvET/5pi8ERiSe6vRmHSKoifLurO+CF0P4w48Nf
Wb2DK78Psu9m4J0Y9WIGWdv9KwuyuuyeS7gGYyTXAi1xC3GIbJAmgurg8++J
XS4ynxHMIsq+F8l3CCCmJLOyIOgpiYJLPYn2hHtwVRH1NRnQnpJh7kQWl2uE
it/fjs6DQiiH5VJxS4iwKv7aUPmnde1hSG/PgleQ6v5N7T97BJA5kjzx4+0U
Uc+0ebrJ5ApZpofNn1raCXOEONnHWFruM2fGvDKi2ubAiidF6DI34aVMPA3G
ZRGAXi9fIUWdNT49IOWUI7m3Uu4x9WBclybHjad5d+FQUX1Xl/fVpB3kmUIr
yUG5+SVq0x2jnYVoff02eVH2c+Mwq0Rx1UbdrWbOZ1fgVYo3yJhOaTZ0hCiN
K8yd/j6mScT8mhHAS7rme48CzJSCZkHya6N2gBMZyB8n3Kd1nun7al6KgIHh
Kwul8NGcqOcvVtVD/R7P/LeP65flMvCiov+rIL5062kq8T/o1v4rDE6GaJCv
QyfUoJlfInxKTXJKFFlsELR/BiSk1DbX//lD/ZQ8lFN14s1o+49poG7iQagn
oidLukt1FzWnhw8Bnf2Or90M/eJrVQLQFjqO0A0/zgai38QAEO8wvh0qOPJ+
OJ8bvHZAE5YXjbha+4NnqW4Rbof2BDVdVG1iG9j/xoYegQvWeaRf2L3MtXYY
bqWaNf/xUeq3PuUhw27g9ZnV6tgQjT5cOhHj1s//tt0HKSIyGAT1ao+7Vdfh
7GhOCU2elsKJPTpxqWP5F9biVXc/QMQV1BD/haN1CJL3F3mjvPzt4KzIBr5H
KXimayHqVMj7A8r1AJUCmorkqUkf99dK/oFK8HJgzFJfB/ALZrxhR+cApWFx
5Xbpcw4TMjTSEQd9Ov85kL9lejNUcn6uGXSfXFlR6+yQJwpv11umPNau+v90
mMmgVQiITjkhOUUdhW14KuR9wGmHc0MMZBpPlVxHkcPWlI9oQNcKaAFtiQ09
OSro6LHYfd4xYlsaG7lojGXU8GrrCpHUJiHiVP4INTgenk3o05yNBo/ciCwU
3s84TFB71vM/PAMHitbEThVxFECpoW6BZhrg7/fELiX1oNVUueaDV0bpZYcN
uKbAbjx5ZWA2EYTADiX50s5vbPWSDvxr/smCK45yxezUemyVX5xkfXTFDTJb
wNaroHmOH3mIpc4VbDUfFgr8CU+nsCxk7tsDZyNJi/Q9QvExB21xW70pQjuE
rY/rMjdQbnhLwQ7YPSg7ebStBzmWKIMk7wFDZcObcDPTkEW1vjI/GcOqf4/u
IbBWyioKyks8jBRKgf2mCiosljIp3U8fa6oodIMVHPTogrDADz62UrClThHT
LCwq0NqHFxKHVCrRTIRbzWZRCgNxGKilbtISnppzOoVv/Vu3A9xHRFBJrnMD
3eTgA254mU63kYsb8PEutu7HOce50hQ7HYC5QwnNi/3Mf2sdzK96Fy9VUkQa
xSEImppdjqZ+9hlzXuTMztoH4V97KVv4wBMOaAK3Y1l7nhToDkJ4KKKiSWs+
OQKsD9rxjR8XlVzBFUr4A6bTYnC81u15jQ8ZUei6oAh+pt9hjzu3w6kxVoQp
qAhosY1JOJ+OVC92V1D2860OBPWw1UryAXgbyvz3FDZyHn7/nfC0uIHn5e9Y
F3LVzsnnQdF7kD9EpXGqrQ+lkjCOEgN8q20J+gLINdaz0YyD/6LAmBkeXF5U
z2j2qZs7Gnm2AGQMgsvBkhfmjDFID8YQw9/XMqndlUCeGVNvE/IODS2w9BaS
gwxYLdod0r7W0UVJymzg4CPzfvMo9BTWWwG4E07VX17WkeuffYDsUtDnh7lx
evjnj33ZmtnIMhO3z9VL+jWjtyhsLhplhfZy5BagnOMrJSAQIHLqOwhmGvRU
mw2uvrQYpWoXpvk0NOXbLSBQ/O7g7zg6unBORIq752pFCA52IEZAQmlgyZUl
hNxsTwOxUQFHAPtYM5qLztaT4rgxMVNi+ZwNAbiMy0kdmwIXUFNr763wGOGn
Nl89lbda5Of5XbT/cgygjv4ZLVu6vdHpkZE9w/QqhSmPfiMDW0IE2eMgvXKw
TY9Fj5EIDK2o8mAo2ujUjOfLEd09upZY9bjm55cPPA6zPPJcnbmQ6LvVwYGV
rsvu2pcmKXwPZTBZw3C9rz1Tyo/j/15GClr+Gw9G80n1X2spprhq04LVHjjo
N29Ii7J8IwhJQlfuKo1eQCHP94RMKsdWGOTsuVRmP4q3366LPBkd9ElJkVkO
hznJplO4NOMI3U2mdBs63+p6Qkg2vRrMmNM2kSQW0iUfz2epW/mSA9xCLG8X
yn68ZF5VKRPb/VQVRfgZSjwIshEM7U2pGmxn9P3x8PuznoC48DQSeqPD0C0l
F4sjOsYrrWA+gQtc2Fxe1IuupF2e8WfzujZTjqGZMbtMbIlQOsmauClqyzae
7s9tXfHmZvzj+u531D48Re4HP4j/octaRxROjZ/wnVAQMSFKpbaflGbzjgE/
cno9yyBvPXGQCrED4yAUHGPPQMIcbYqGKA9PM/5RdJ8G8eFG7gQINwamOZim
Nj3LXyOiZRE7/l9D5se/dhQfWaBCkyNYlWcK9lc7pi+mzLWS3AmU7HcbpZp9
hr3cW1/MSOGSFCz8uzjU5nelqD3JOQ/0tKMG6x1IyYokxI2bvCPpvZBprVbD
z6kWhinNakYVmS9+HTPOmKNMyCRPuJPw5N5QfLNkijKCa99a+5B0qAVy9Ao1
Ho0iIU56Z8XnGmeJ2g9xBMQY+H+MRcTEYXYG7gAD2YcwnVV786ILoZig0nqf
Hfpn7iuHq600vuhjXO6rrQEW17dAs4ifAXsjwWqRSXI3CHAWJ67iqai25HjG
ugsIAqxhuKgLjNwWovE7j+t4P53NkjMWj8oJyCytpHiLpxUl9LLyCSOop+Ri
WBgxpU7MjKqXCGbtvqznop438mh2ZJ60WjKokOwNImO4bGwuzI138uYzylDe
4n4lTiDfLiOxLXU067KIPxM1Q5oWH3PK5KQxc7TtgADiKH9woN89+7RQVm3t
bWdA9S6xlMoe0ZBq1/wY6q7ZkjOJRxs5kUJYk/An3z9BBT+kaM31f9tD82oM
92FL0Z560FVpm7mMqnpIJ1kTccrK72GX2BM2rsriB1qADSXn6cey/++JtyOl
6BXinTySB0dRWM9zeBiKylF3YkG16GcJAtsT3ViS8EFhJ64NwIrTztiCvVLR
i9WcmAgd96ncoTl6cL4m6+cdSFig4eqZoECnGVobQNdEiEHRZI7SL18tsozD
JQM7D7O7886lyz4PiHbgqpfapj9q3cDvKVGcXlsHpcfnyxI1Vq8E3mH5mUwi
RRthAjbezZ/BTxjludwPiUb4ocMN22pNsg7kppYHOuVYOe0DT605ZytUeaZk
Bvk6RAcVo7YcXp7kR+RDvNgUajcBVx/Y+lR+MIqJ6C/LWOvWBJHc1qHRbJg0
pYLnnONMG3goCxMTl+xgHrK14jRdGDxaIS1/7S7Rt7Ka+wcDIUcic13njidF
+QnrtQJWAX/f7Tf7/q3i//a0JIc1pQRgw5lqe5dSFZanIjcmtuYsuaBLsYmC
E+5vUCRydUo7nZGGJFwO8UqFCvJPV2hoaGhaPp7X3E7kvgyrxtzek1/LcMRc
6d68e0g11cQKjSI31/lsePaogpAkDo7IiMKR3D2FhSEzAYEozsOD8fe6/F7n
v3U7lBMXXo7ETdLTgbmW6jzmJDHHhOkRHjqrgaF9ou9IxOD4Tc0XG3lm9SVj
252Qc9KUo3qvfLVcv2tzzDPzwQyX+/+jRbSlqybLdVMgBFJ+RlZSyeM8gZj6
Y33oT7qn+W8EZAOmCj7sKMc0CAq1qybqr2qrgnaoODwDxTq25VebYbhLjbyM
8m5RfgVLb3G/htU9Uvvy9waCyXCD7t5SoQoUQ8xKT89vC28I1MnBZ0EfXjiF
WfuleluUIN//OeB8k8s5Es1ClYGqUIPDi97g0LjthdNrPjmoLiHWrssdeR6E
Az//loRG5gw0AGFKLW9UHXH+BU3wIcU/dIdcTNPkgZrq+y/WYzlE6qtTa/tT
dV+7Ni/nkngF/jB5oCPB8hx8g4R1tbFWnHJ1r3BKwIyIXarcbt1NRVdmF2b1
EJbO+TVDB6ptFsblJq9NJrZjbDlbpsnqw3KQtua0zMtKYrhST7d5r0EIP44T
6tCdaI72VEJ6V3uACNO75nX/lU3bHCIVCbQNBVvNGTJFmuW6Vq9VXFjgOjqG
kGVAhWrGGPhAHS8ASAkHwGolu3Qh2reWV3rwIfM8CnBpZW/alpfdQwX9z/qJ
+eQBOC0YOxQxVJpwizb7QtH2qcxbvBS7KZ39/GVQrkONBHswqjoJsEK8C/u0
JW5KL9dwUCwY1AmO8QwqfxZG7zj0AySYjpXItzYwzVDt1IxJtNd0zK7mfJg8
VHyaIu2wtAML/fJYC0qeq8wU+AiUevjMrqpanDTyZS80NbCwygUTQAPokGNz
QT/NlB3Jgb7cUy+4YNQI9RK+28qM1Bsm4A975biS/mgpBxpyo+cqhhjRgxhn
yRLBSBPVHN1QBiEesPI46tHbh7KvrYozSRiEPj0pfl3FVO0I/Von7h+WcGsc
3gEhYh++nmy+hE4Ls8pt4xJEEi8Z+SBT+fCLykAGCd37fCmAzK2tON4w+FE6
GsyWudNssAhmy/C10Or+rasNruxDbmMZND41ZDMO0dh9pT2vNWAr8NPbF441
UfWjnkO88xdeENeAbWRyQ64DWsGNE5pc+gQm+9kP8wSsAgXN9maqJvELWKf9
Hb+SzQy0j6wnt9xld2uL96E0lnao+RJlk5NRgG1xM4l8LiQ6EPiX8wrzh1vO
5yfRz+7xHQvFVtfBZPSOqmKCbcEqfZWb0GY3Xx7vTCvknmzD9o35Lcc/sv/d
9UucQWwGtnHikS5N2JgKZ4ZTABuk0WsPYHlTg7yp+YxlseNGtP5oYf9aIRTM
runVGn6LnBn2idwbOKPGveAJz5dweB6SfOgdx3RQQUqXro62a7UqlWQAEvOJ
n1nuDD1STO/mslpqrMr3OrCCO1buzsczjvcKNJ7nI1yP0pmIBKuzRwLPHbrs
fI3ZPGNM4J2NWPULnPOIWdOZ3JudINRDHiOw/+jbDL254g2U145cDfmSwxif
Na8yjxjco8Dxb/zNznuYgSj8WNkaXTSkSoibl0Kmk1oAMXhCHHMgmzqjAWy/
7yzqxIKo3hjjYd3Xx2foE2SZs5ibeMIRneq9qrsHY3h+E7xiWFkHKaDqX7dv
vOV4bkBXRNP4YLlZBBJ+fNNzrLpMAVr0lb9cnC5TXbt4Uj61OO2OURr0ByPe
XemSSRiG76UK3iglcItrbGA/du4dUz2tsYBkwQtpowMS4Ci6d0ROmXegLBwH
bG7iZfs3z3v4aO0LFInSPPJgmH0Kp+bg+jIIeqGLyD9/6c/LhQ2Pxe4qXW7h
MyNvIQDvcsLgs7BeeepdugSgiw7V6ZKxtyGBN/oteEERG+PNm1pp7/2ndhpC
QzPDimllyQKpaDTwuROt99iwIjFHCumnNo/QWvZnnT4U0jN/5ZmwQpacqDCx
mF+m9d8d0EYGlbTujdwFrTcLBIz0P3T2EnP/Q520swq98s5LMgbxzppa/4l+
Msa7AMlfV+JEHe3PdIB99lk2pItE/umRP+wP0KBZpM7+0bkYOOca5aTaBTTF
98MTYPonZ7u0P6Jq30VDGIqRS5zugNuTPlN/ERzCQ2Dt7e3bqOEOFKDy0ofU
JOkRGfq4cdDOzlkjV/Ipjk1yPCRhJXfWUYz0UhXzFPPICSLu7qukvYOqtsJt
ZplK5y1J9+FVMH2dWeX2z6FV3aVLiNZ+jMD2BKaf2FyL1/0qVzH+LGd3iHBd
59NJ31chPhd7ZtsrvX3JKUOm/oWB3MMKG4ctX4X3G+K3yDqTYvj8k4yCj41J
V7sBhlctIzjfamBxH6J5ebhIDUV3QKE0McFalekLA9DrcSiuqpVDnF6M2P5f
CD3HHBDqwuS+0eGBkXCo7CzJfrAKq2WvtmCNvPvZ7IKsLfdyxYxqFkVvVZDx
IKuqAwK3NpjGEjKAN8Sreb9YLrMW8dV7kswp1k64mpxElvkLBBdfJhX1q/MC
vIdv+oBebILj8WgfmSz0DFqzB4VqqEh6pZ6a9OExJs9HKAFsZCyTuj14RyUT
qy94+3UNPalnsKXDrmnZzs/LMaclADbt2iAZ4hCYStwkPm1KorqhrJK0mn0A
GB/HGyg1jtyRQMdDWS1YxdCkNST6tU2Eqdi4NOdGiQvvrC5z5KmXrBGLoGXr
ztdMTh7LME0VMswlipalCTq1t2FczZ6fOALt9G2XbiuDtKBiNdTKzm2xN93d
XXoD71/vQYDuiTydpw3GfNfRgOLE1LpiMVHB+wVNCL6rkV2VbVzk7boWuTyG
05fNUG9xRVfUGVkdoqjR19uUutPdgnW7RVbLdgbm4kD1g/QM34w4mlT5Patb
flBXJNDRm7xsWNgNDtfg+E0Z/a1g90jQJcqjnrekxPlq7MVl0KPBS6Q2rIHd
uEiphHZQKhJ3zRFodlqMJ5RpYnsBfkCpvK8qB0MMQsI85PouTDycyv2umK1j
HswMet506r03Abu7iitC46eU+PisivvXo400BG8A2Y6F8An+gXqxKYw+konz
iO5n/wTQcpBXkMYsWhFQBQpof1UMrt0iGOeAVG1iUF4+9FryVxRNW/tlEdRQ
w8KA3M/NsNMGaS2iG0Fl2ELEKEYVMNAUB2b+1riv6FAGf3d15aj0RE6CkZvA
RFNFyuVVjYfbS+fZ71lE1AdoizmGC0Ps2eXcAG0p9Lnmigd6oaPxcn7wF1pV
O7DCYiY0Uare3PoDZClP9kGZrkm6MNn91bmYnJvhqXKojc5CEwCsopCgN1E6
vjG0QoAlpDkpyp8qKLjUQRBj+S5jmVhdVCC6cDH3Ppf3uI5mRgsuoyv3YTAO
DT1mgx9UirI/HQtrwU1mAE4LvP/Jl/qv/ulHkE9jP4zj+3TAR2iyLLbgIjSM
Zua7K83DyK5ctVcwDg43vf2lL7/DWWaSIYgZ/nZiWYYPlfNPj/Ol8+i04H5P
j1NPtqPauJwjYS72Sw5mtimzGOI77LaemKo9HO5TeSjuwMNg9IaOzrLBf5eF
FhvsfiaIcx+S6512P0j5g1Y1TWWwCb6xuq+mKkRYQm43yJjvpaa/SSZQPJS7
IC3bOZAV0/zNeU7oeVkoZzH+o5MA1UsEY/apXwyhL7cUCOPsfyvD1Bq/oTsn
uhCq/gnub8oEwdMgiQf9fFr7XXdUPl2H/h5ESCTSWchpLnlYPXBBFb6HUDKJ
R3UncKbiA06w6oMwGY6z6Hqhn6LZfffL3Kr0Oxu7oy4X/F0QHDytBs+rrXuY
44eqYqWSM9wjcM/+UU7g7dkWWb4lxi0kikJyao500QBBpxIjZcVzrxlCtAbx
Lib2qjZSEbncqfbPKzU6swhtncB5xJQTyxrYP78s4eRNQaSTYNs6W7MI4aru
/Drk412hLh3f5ZLOVBCGVT7SgWivl+Aw2JGQcRNEHvium/OfH6sTGN2Pysvv
fAKlqFOezbjtMPT4Sxs6fTAMM4alS1iGDDnkFbBgflTcHlj6ZuAz6cqUcXaW
2tS1k0s54D0Q82LRqaShfkoXPe3f+dvrAwjoSfNrQoQ6eYfn4WWw22nHFLpv
Ov0Oyg2Ou8AWnX2XZqsmr0tvwf5jFWqBXb8VHOKXdES7xDMvo/02TSiTnGVS
EVp/y8Sl0CY4yb+GfqWER9bPWj301aoQoUOE6Jbw+WJa7yyqEMiI2iBPU0NJ
+1JWZfwvTJ6ccHp6MTgb76ZZFuT3hyWxKsJx5ukq0tnhoeU+/KczmL2jo+A2
pVqECAinYRxLJDVuQcCOD+kl9grWtWDMTtnTgH9FVORqn8ZawgPaDAfq4Jku
cGYlYHSi3dOVFaLMT2ZKZ6v5L8ebB06OCYdWj4S6h0RoxBoocTp/WmPSUB17
LWa3kFDPTcxXJK+HKT5IUyBhyyU8HGmwtkz8nd9CFJG7xwS5MKF7VPJH1Jxs
E0XdqG+fhblz1ucJHICtWQa+6BJ5ttnan4Kl+Y8hWBvN/rDH6w7a/4e2xZqO
esqroAZ0r75XyBb+Wvo4JmzxI2EQR+haH55JBcqC/hin2k1PUaEUo4Dsax8Y
ltGSL6wrx73Ef36anUsmRKNarO575Ri8rM6vx/7f4p/wKkByWcTnz09V2Zgj
eklfxKnBuZPWMjpasMxmP0MEGqtPUU3xw2nV7N5a5uT7ikVHZWaDdx6TwEtN
GLtayqY5Drxo8lRLgFpggCMVaRBQDlPi3IDyQfn5Cg9dau+68ndaYI7qxR5x
I+tUiWcAyINuj50bLxFRx3NaAOZnnYrFzc5KKXpd5zv28owZd6lx4hO8GqmL
BhJWFQzOA0fcyXM0KI6PYgCh9QAVHa+nnyC4T+3YvhaAge4J/n/pYL71S8XX
+OuZ49T6OCcJgDgqSaMxiTCAkBVRuVtpyRp1r3Id4mDByGOimTfPpaJ4ZXnd
To6hX/QG0weWEPtQIwTvPyYC/7992+9NyaWT+ygY8rYXg44KysFQdLXyrtQ3
GzJu4TEe8TmBU+vybvJcXuWrrW1CzJW7JlHxAch3CpGC+ydvSb+hJt/Q0rQV
2G4wOTDh+Q684jpU8yMibtXHKsBOj2MUfdXtSMBJHx+cd4oONTPI3xbjQBDD
4rSGQwYzPHaHii1pCLdfPPcVbWkFjjnc0Kf5kXnxXJuaZgjUYbI5Gw/l2zrb
gDeUzReIYWQ5Et382Lq4ts2+dp58yH7uqKkdoK9zngI3vh5Rz23brsfpVuvg
orL3wWCQqiX9N41s4TqDnekYFYinBZ2vKH1sB6kjwcx/skrhYEd3gPEXtwUk
/AS1m4Lw1E0fkqqTVuc9d5Z3HHx/dAg6wdq/pS409B4PS8B7t8R2SRLimQwh
xDzdV5Tb/m41XlXGncusuhzL3H/GFOty66Al1XJOx7F4rfyYG8S2ZzOmXPI9
4+zUAhgGeklvG2VXzwy0YVhMrker5nAlTZNrS1dFazN+qkhCQIj5cOZEmSh3
NcG55JEGxApcFkl/eiFois/pvPVN63ekx2ny8d+aFlXGpaJyzVDLicjIRf69
SvKvT15u2O1bhemOal0Mf4YWEgqloU8CEjVPlYkCYU0ItGRKQpRdE5iet2EL
a2eoedp77+lNbDiLJjuamPhqZPO5ynF5IB5ur6qDxMWcTtmLEW4C0N1dILQh
WA1yr652cIdXYNQmxC5HfUMadP7v2/6WHbBkkQFErRebHUVSM6QuGKZ5G4QA
jB7HXAkKWnlSJ9q4bgMxIKZdh6gd4c0KLnF+TTkMYFcbvlWmiOR4Zq/Oyzqi
tfwLMnlS8Y0e+JvAHDI7OqS4cL+lMqkUIGZAyVgPO5IZs68fXHcUBkP+p0fj
RkbH5OgBqZMmeseyYWuNO+km+kz7HqeMN5/YTIt0DghW36H0H0fSZHzHxCCA
56cVcgekzuqi7x2eT8uj43sUb7mN4UBYK01+dE+aSw5z5lWlKAqAk8hMkZ9p
uxs/OarerZW6aWfPmtuZmJTcYIbUI4aZ9vgrEu3N0BwtVXEmfBCimrJRbaeT
QNe0DkkE77BCAtJq++WECHfyvZpMwTsH++FU4sGQ278Dlh+JKsuNhH2OfEV3
umFeYl4njWE4pkXnbD9Z+KlECv/5B3mGhVFvTB7Q4K++0ewG3jTOHXm+o44Q
lrF4xlQP42CYwtyYVCirxDQ9b2FDdUYD4OvofZuKxbXouacdPasM6Yv949T0
4IAY82FF/jnjq/ergs7ZnXpqkODX2y4jSh3EP5vygkLa6iy2GMYrADm/7oTn
OKtK1g4qlHp0oUQncE2XKU4rYDSvfeMYle+337z5Ppa1kBkeVDFg8xQiG5Rn
rdO2RGjKPatSX85GlWz0b/59uEG5f9dO2IwNUNLq2paM7CesEelqAN9SlEZa
5WXIj6XCxL47xNGSPPMkWTCTqM0WbK4a3JqLKSvxaLf8ai+cEXbBhRpauFE5
1746vScq/qJ/sjCxbwWHCfuZRPPbD3vE2/Wp3tMz5bvDPUbcINa8RiqOZ5bU
Nj0AkmWNOOCRuP7Ko0GI79qbKtpcvClwOMvfQii/ttx+/NbevY/xMWL9KyYD
1OBywlgjooNk7u+8s/i4jK47PWI9yVZ1ibT0w+k98LTGn1EWISre7qRwUHwW
bmE5cZLjPSv0Jya4QrGMY1Iwa1OWePIa/ln2fZvXsF6WQQZCMRltP1tbPuRB
PlTK1f3xw1GAj9j4KpyITZ3ZSZ9hmMSeNQl5SmOGYXBd2AfXefsOGC8e2JS4
TwJOpllv869wk4S7pFJFIxJqEXGvlyMsAizFT4sQ8j786TqPdqbW8WiOe5hx
paCMoFRWJxz9BLB/354iLZNHH7b38LuLFaj+qNOluKKXD1chrtnPtLKXQI8G
PFbOKwtpQdw7CPpAT9GfGsXam+R6ELlbz/RNJreualJK9UJfQaVpAdw4EQ4c
z5LNqd0IRwq23aZB2zjE+1rqfNqrtKyyis38/izSJZhu+CKgflj6eTuUw5md
cRnGL2xAn4SlgSVFLus2jkS5c2xhOTRxzRdPdGtf1GCQSDO29XwLFtsUwGfW
oeAPh3XqmBvKz49cT7g9xmLMqsoF4LLoJd6udok3AMp4jViE64AewNDT1Cxh
+OBxLPqP5DVPyz1WAKOLPdIZfcAeNBQb6H/kDFeHtv5E0Ye6U81QNio1Ygk5
Pwa+qY2Gkk7jHCTjghSjEw5DkFwI3vf79fzn1WzvkxPA/bof9qzt93UVFA7T
7w0x8bm3J40SNVXFMG9xTDk4HP3K615mtZ6PlslbrkSfl0gIDg6uQ2TUDT2U
r7k7BFyyc7CYxUpfQsZlJd0jn6ij3H9A0ARenzOy+f4/8U0kq//hGaJQIPGf
gnfqbwR7IGamkW1m7nhTV2rTc7AL4r5mRGtQ5FqiBHvg4jzVY+G1naGqatSz
3Q8du3UEzZi8+2qA8oXNPjdc0Cfs+dM9iEodqsEqx9ojGt+WqBy3Ss2kjcnN
NHeuuY2tXE8Lb8R9Cp0CrzzgSKyKE0jwtTT/V5Z5ubo5U5qzpgKWCCPiDEVT
SBB2tyvMVDHDvppsuIcxkGk5/fl4BzqLGzai9FRFXC5NgmyRNOSQxs2MouB0
3PlrqiSzxE1TIXrk/l76kDPihQLaV0rssubVzYiraV4SJkcX9DtPDU+UJ38j
Ez7+ZxuuAWT0P8lUHScooxHmgZ0r9xlMTQYZcnBb+HaXXXMnLhD8ZnihX/B6
SGlrzFhr/ZUMhZU8U7cI4Rk51eL6MU8hy1NBGXAUMufXHvH+esQCmM+mNVuk
XO5t79psA4YoUM/znO8VUfPtGwKsOX6qHxhTnw9wvADKB9VpjunQZTgOLkhJ
AkycLYuth+n7f1P6b4M6kN8S8RaRL56W9dig/flg7lSaFemNGysXZweLwg3r
vebUhuYWSh8YoW84GkynBFejaOdTy4M7XBanulfRxk3JcPHC5OHApYuXRK76
kmgQjFtp+lheg1/piwiqpR8BuiCFIljf1aNt59ZR2VQxlPaVtp1rnID0DDp8
xzySwNBMwAxxHQVZJTxKQwUEHL16YNUf2wuEwuWlISdktEQVUAxSq8AS0Xm1
KazvCpkBO73YQPIvlPsriTFUR1AlLmYv/7HKCk9IWf5KFUcAc9woIe/oO+gU
J6VlBn884jPggzsVeLgd6qqQlPzfW6NIFYqYIXMDSNdeWn9z7dMN8fsz/Nsb
IsOlQJ4kpNma0AP+LNJESHpUF9sT8rfe7EDXQkvSGr6aCLrxaEH7pIzVxP7m
m+ZDV2hXCmrfHTQjHtsdjCt3mjD5zGuxVX55xbaWgJfKZFEmGSdU9mhW9ofj
BaAESIQgWyCcafLJ5KEKLKV3TpLx+Mpul8SO1Tto7s56BPekbDMsYH7tmQlh
pH2oav+Vnw/XsVfQTh6GjusIUCBuf13+i9+xhz4PFvDCLBw9ebgPPAN5U02Z
1z3l1oXk+BTXoIcWcZqcM9x6jZeNUAE70k9YdVWs6JUrL6opoGuu93n1qoiC
Mx6bf3J6T1D1xGU+rB1pYlkAMFwa3lZt17e0IW4zWNJ2xxHPNPL/P40dGUhX
xO5GQpfpJaakvabb1gI7Xes6+0dWsScK8XMJeXCQyvFIvf3NnHqTNHq6Qsqa
SQCkXaOWHXdYqrewtPzvIUb7eg6wM1sIHPc5bunvoJBF471kFCttkSFfbePf
4mR7mvkUMQdubiKMgmcqOJIrWYeaMLsPfH7Qn4S0l8A2RiKqF7Q83hBCrHDp
Y+O0xn4ajeXpEDy0dytjlpZs6h70fncYaTLL9U/pnHSfcmzTsC7paSUabIFO
w4LQK4w0cgerb4wJCD1vlSuKYrEPBDsDJSOVObRYGf3gVXQgKz/Fj/tkEaHc
BVxTwy+RSrtnYKqVQW/5nHC8GCZ44eiFRb6YnYjdXG7oJ1SDv8/YlYUH0kRS
+x0VIQjyIqq8o5tpf7Yb0eBPt+JG1J+Obk7r03FDxWM2PikDqaWOcEVx/hij
lU42RFkCdXtUpCvOqXwXiwvwZFcoYIalcD0umM/jqmLdccGax1oFt91Wc1Nn
j30dlL4o2PpIHpktTRGo8fMv2q+s1IDO3YjZqAXF+K8uypUwhNQ8zsBdH/eP
7vMW1glPgnfsIHtBH8MXE9h2b0tl4wrhO1/+b5ezaC594dk0Oud7VZCCD4X5
ajS1fN3InYxsCdx2aZOIi4Hd4N4ODl5wf4S/7Hz1Hctq8gULF0Bx1TILsj1W
8Dp7Bo+xz7FVdwgpc3gCxAazeIQ0Z4bQlmeeVSG29+z57stCVeNClHjcgEUi
EVjLn9i3HhPb4/rEPZz5RMwAPNcxKSHgS3uT8EuqlE/8IO7SXdL8ANcyFgHk
4Qmn+ZuRx55/AH9W0w8vAKe+kfC/pKqBeJpbNaRrKa2xZTov9esV4s+eZHye
BflF38V69Gmcu+HOZRGnOvjt0vgzqQW8LDjeoaeBMrAlgBQC7VmM+eorFGqJ
guzXRwqzjlqEU/qt/fqQKkm+uzNFqvpdmTdECU5hrGX8bWldkb1aX1Zd56j1
jsFbKl/HEjQIHy1eogXonRwLHN/RwECKcaOiHR4R8qzmEjfZbp8G2tWLo9PG
+c8v0lyCExV23tn+u9UZ6wElyAeorkIcc1QEJENNgH5c1VrmknkM8jUHT0E1
wMmhg+KapcpJEZIuFxVC0sHaTkagokVeBZJDFIK9pj/3aWv4pKL0MW9+Q4mn
NrS93qEkdYcA0PXoaoqApgo8IHcYxD5nZJXmBZoDik+a50ZVTrcM4awiXYSd
0pAmafCHzKxzy3fu0xsj+VyIbXGtfjFlC0ZsJ/xh7SqIe7NZCQ8jgkIDPkRR
JyKtksqI5tDoEl9G89UkQIYwKAQLvyXTr+Dd94TaPrB4nPLSqFcifYHgyxwH
GYf4KlNGFBDwKRfAG0Zrt3SUZ70GabYLVHgCFMh8hfYMwj6k+OHjIae+dSrf
y3LpIBcvnlrY4B95bCFcfmwewjCDyw+VNhpECwZEM/4LU3WWAmhE77NiZ33/
awGVqkvZ+zgaVD1Q/zWNtYBzL5hnTdh5Gqq+IPrXDBTiAVjb20xBkx3Fbfqa
1oramDjmO8OQhgmVXAZLXk/6wMCCJvUdfzHFgQY5TQ5KNhxY9E1jE8YJTWn1
lt8S4osZSR1/sVyGfglXNqrhrFUk2NxnrNyW0l7dZXu3f4VtTBFsvVeRNvC2
nL+Ub6ibfTEf74kd6bWpoMvN0SgY5fzw+bCoWF+3Gdvz4WObfeKVH0pQizUy
gpg+CguWoi1L99jwlSKE+WTnbE2Rw4FsPJqgunfcnz9NTSY3Shr33J1kHL8G
bsYlPdwqcO2q6p7rqDnt5YqbSay6tapgeKtl4WULEpq9v6u9x3Mtn9IOdngk
aqj5s6ScqpiX8XaeLP6qy2ONZOCzugYgDrpoBtFHFptCZeQlLuwSL7XWnOBB
04HfJfM1z8PPoxoP1q+EbRLRw++J0ARxCLhbZgnYBDa6giaby/nLdcmJ7XlY
wen+bezt36XxChgW7U/NcQsZMXjeKaO4NH1GBuMQiE93/ppmCeD9MQRZnanb
igw1rbEVTgT1Uou2tn8/l/ukscJyY72+JUKsAaxX8CGEJhhT2uilAd77UR0z
jocxHLUKOS5nEng5JrHPYgA19cUrPWzcwCcHjGEQoW1td3QRHvqAlP+fdI4j
8ef/m1VBfRPJxGrUUdpjk4XdjnViHHlzuc1N/QEnglWMj+6m/JyW8jl+xMgW
3PFh1CTx6A2iBMahaWl5OW4B4tlAWqW0yOM6dgAB0LES/4UIgUFvSUb4rlzs
VU5AjISb3M/jgmdVfwSRzNSDq2QmzCQF/f833cK88IpMuPk9GQCOQf7RREQA
k/m6N54fELgg17smf4WQeQtBAmSmP2UoaRw2Mk/cES+NA1bsNe594w1D7Z68
mTjoIrUKwEAROZ6lpL0I6tMOylAi2TB4m6aOaPwyTPWuZAXLa08nA/jT6oec
nd2KKOJD9Mg4gIXvNCvtZYkaLjsRFSiWaKcBDJj3rDXC+/zQmdJi5VLjx39u
mdHqI4jShd6nwEnnAIlAJJTgUyETflLtPwrNnVywO0Z1xz4S0N+XjFnKKUyQ
RGxC8H8pEOsSA1NojBfXIYDIozDQSS2mUdmfnzMw+iRHHNDRDkZxOFvMb47G
NrL17A+3gLKpep7t6J6M38T0XxGve1H2uiM9tKX/7EpqaTfkyrv4Q1rK92wv
QxnVrue11d5OtZTNDrgpfhyHyx5Dj6uuTB5fWOcJBwycvrZEQekKeXZfMGok
M/yvsUJBoonbWmcTuduyrgy6MJHhBs3ZGkEqCuxMi1CZoYd6Xxc25DKPNKYx
wKnvIJ51o9qlXmjvx5xkg2AzrzB5O7jDpBxR5BFo1U+rlCSyN3y8cyh9Q3p4
MShj+b8ZVqWGqCs0qk9HFCE3OD577HfbbPG3QmD6xUV7xA9JZ55l7BTxSQme
okCSosta/DTIN8YJW9SAgqGALlYMMCasclryAHk59tL0auclMxkOo3wuRTcD
yAy2YaV/lUj4flmHK0I7QU/kSt9jJjP4W5hHhCa5kog3wW32Q9L8oFjmGyz5
SiUt+JbgtDBMqrgsnu8R4NP88WCT2uT/vLGTVddoMn5piL39YGoyMKFXHQc9
CPDOdp20XAMaSPaF8mcykq2PGwTa/KKaqQVPz7YdjWIuo/2G8/P7c91FCo/B
f5FfNiTcqfzcISbnn6Ekpsjd482BE2pNUNkmDJs8HEEX46pzQPt+/MAxPbFq
tXCdHz+Kj7Efxz/zmNUg3eXCOe5L2v5SiYf17vKd5hK1lSZRiNilEDl88u6Q
4bjU7Il73oQIV2fY4ihkr888qedVf5xH0la3xyCRrAf0INV1wPxOwWq5FsJ0
wZs3K4pHKtjaIybuEv5VU5TalSTAe9HTmd6yiI892U+IEcanllwtPtKm3mTh
JV7HWwScDDQaK9hE7sDcR5lUfEhqcMmCKS40u2PQMtg39SWRxf4uYo+Xk8ma
Snqp9S9+m46KpVnrBFq2ajK1/bzyCgo7B4sZV2jf8qt6OnSzTPCIijrAVG7e
IA1VnhlbeKIgi/GA05a1k+ihIdomzEMmkuS7LLMqc3lagxDXRPPlKIAVTf1M
oxGhpT80cGZue5CqtDNLF+l3IVIrPIlFxl7/uFjz61j8hDBvGi2PfKEDVpsm
1i6DiC3muhE5gUDMPj7RVdFiTjUULhbBe/NBTyjRZC5svW/M/7Rx6C1VTthR
JF08c6m7d8LUmgVzRvhBVl850XKmBYVktZraD+ot92O47U1RAxihDs/TLqQI
BsBdNtRGQIJxJYAPmP/0PGxFZEM2RAXBCcnYw4dMaGVQn1apg7aiCJXKnHaz
KiVT/9JfIuNfDvcE+la+f5cxaTqrd9R92QIaWgHtYui/XIgWoTawlc3YlxgJ
Eno3tqHJmzevHOY3ebvbX+LpaOj+SgWEP+j7n3wYgEX8R3pCUku1hNCYMWZE
gdGgw/mglnyOh2a6LN5faFWXS4uctollbZzffAT5crxREpp8DZ8WccgR+P7b
+3y5wY6ANvI8eYwe5/BSMIqB+0bLBVmcinl3jSksl+gl7WxvbeVgrLUb5tsp
R+bCb5qQhYqb1w29Q/cvVfiY98f9I7OpnShVn0C/+/Mh+CcJL/inIth1MvPp
SpxToSiEoq9aF3alhBxc5ZTs1YcznJCgdsIOyDfqrw8MnugR+FCw4rnd3v+f
ZWg5w7boF1ll27wQ6Nj+wI7DzQEUIWREqWqr2jh7O2vJvv8knNZAobj3Zu6v
4dQdo6zU6js3AsYGSNpoT+tEztPep38eCx0BNJtFEzcymUyrm7hdgfWCG7+V
Y1GsXUYY2MgKuaQ2fR4OZ/c5jkQYNGBsISFnsC1mnedOEFwYwzs/XtB5Eir6
uqoRXZH47oeKlemgIHfenCgnKQVFp5pqFZmdOo4cJl1RYtpjasQxXkayvMSD
BKT3+EaTcSWGjEinhM7xqniRkZwoL7OxvgFLGXzZ/aUCLRUXH2zLB9coaNZ2
kVGKVXFxkrOiapOJ60CK1NkisVbY5fVUzPQfY5UKQbX4RM9k3uaBVATbuRDT
6mNgb9momlXqgW2aD7YXwkNb82MqWeO2Du9OUoCNR3v6lNArOPeZioQ0LpvH
Dn/gweSXgczzCP/78vNHxjsZivYbvLOewkDTZF3uZhq98xS4ZR18WI1V4yPd
PoQ/UBfUNUN7feHLEIvcx6+y5dnFLe7nlMmQ2aRQjR/c5X+0eSPELpiQ5x8H
YNQYT++yplXWaF11zQd/FSxc/xQtSzs6Ljrt/ggPtiQgrtk12eRX+9FwEvBa
TGD8LHabttmDEkyZmeqRbkwP5tw56Dwm9FpqeSAggCUs7XOEi6JKsIMTperp
5JhA725zyJQgANzujQpgkT+kp+BuKqOpZ6eCXwu/4e7V3b5HkJMn0Ey+AsLJ
KyLlqk76/z0g5eE0WtvhC/jvbEny2C/Kkd6JaV/DK+aW4SR2MqTlkZUNkSiO
t0TIJEiowVhqUkA02cuNWNrZj/WxXCgyzIAuN2NVNlMg2SpDfOSn000SMMti
6mCbRRC/JghNIc1lSGo6VMRosZ2Kq/d383ubNMb7EanIyj/1IQBk428bw2ey
4WmnG/agz08AxLYR9ZAxPkQ3fH1dEJjxDCY9/zdGVL8SX7bZlOBgGFhfIijg
TqpcIPPoHtYfMNT0XaGBgW8pmpgptDHrROtmNLi9WFxMMNa0nv4XI0W3SKo5
TJIy/vfdq266B88hRrdEFawLhTbcj1Vux7+7MOZ0H/0aoHu0W2O3osE+u/2g
HC/iuAiZ3t5StEV5l4EctT43Xav4GEJzIHPGjrdIxCpaXr1vXWIFXuUjxETE
0dgdFZXMxI2kblu3cBphsIk0fhnZc0qXx/36RWacYUA57vFhQIwo1AxLN8ZT
5SgkzeY5/wzpSTKce7cRbTr/IxWxegEfxByhCpYbVi2Ir1G1Myh4OuQbA0zr
BNK894wcAoCXY/kGCZDzFW1SPJcc37LZeAP/LlYvOhjVw8uKNAO/1e8Ff7sh
1fZs9hxxEWXHZzshQ0zLfOHvkAXUAH5wNWN2oC78Z7FV5yZTai8ajrlXRzpv
nIRTByX6ayg/pyudxmhPIZDN1zC0W7PDCESW7yfURiidDdE65tUzwc+/vk87
dTjuohgtl7BoHbbZ/Mrr7Gbhz+bsyvxjKmprBaWDEcjwQrEUmN3+6HgDPEeW
mHXtF6q/Su42wQ82rWy5xfGqMfnNSgqzZdZgWTVSkLbsudGzlXMTSanj3sjM
sa02iqyVoVfZClw5Y1VO+PNEzXJQsJGG4v9K0gMmggMci/uAh1+0c0AGU5oT
QOknK+c7n9/q2iWU3GrWFFXD/amrfRlqU4Vu9iGgOOYSnT3T406Y57CscwtW
IS3ixfxlY5VAHeuvDhy3aDYv34mnCYF73GV4EV1LIA8YkqaONnvLq7uHRxkF
q98yNA2EylGMVl64TYBF3gHBs/DOictksx+hBub+ZPC8yuqcn7n/xCMSFOMG
TcG4MW7iM0HbHukPFiZOc21v7FI7H2UtPov7u9fMpiPht5cTVAzTohiAiKga
ctxAOcbeyBh6kCyFVCHiEtpTMpFb/KUbYeywWDv+dnjnkBv0udSVUAKgc+nJ
LSL4FDnJp6lbwHCN6cRyUUe51ykC0fuS+4Yk5S7lorgWCjMarUVX/BLNsTDV
CilhJEDHNdfWBPJcI7oOTohFcoF0V3Hesb2vgopdtauk6SF19IjlmFh3VGHe
Qxc+INFxef4VEThBlZPqwc36Q+HNNo/ZS82FNJ0Tea5+8V1+GW3g4HObM0Y7
lPHXHxtY93pbNSP3y7TSiDI+RePLyH4PCaV1WkYA6dkMDC99WNkTw4Jublr9
2ivv4cMeb6AlOJq/E5Ntiv9w+1JeDWpC5OgD6LPsjbbaT+cOVomLpUAMJ/vp
YHfCVEYy9OuTY7u+9LF/7VBA+IgSKbg/eMplqY4sXylcbCWsXEod0QDrDjGX
kGp4O4xaLwlGYlTtmAN4n9Khyzx26vtzlFnqo0DSme2wPuC6Ps90g9WhuaBM
06RnmS9LA8jjqyDo5WwRjRse+0ypWzXHA1JvtU98BJ1Ge8PTmnLx+Jn4sl6B
9qG3R565rQ1GafxoG8babWpEoVhNqxcsFY8af+V4hFIe5ZQZf4gr68P0gXmc
fAJz6h/PKiEa2GB32+FGGUKOdNheVIrd58A5CWneAku4kteZdVHmToSVaFU0
YSvwJ5J5xqJCMSZXfcQsT0EWAFe8SSyXRxPpfDpEM8NrqGRMs9JJCxk+Pbr0
0YzUoitLBIfuZyqB9/nXO50SaI2RkiyyfIi8Wf9pDMZT0k7Vj6eMP/58CLmX
EMmg2es9XwC3MulP2GpcUZ1xMixHpZeWRyawUiqlS8nfs7wA3hVWQw2tlkG2
tijtCHGGks6+EZwAPEaimvoGg3DByseWvv+q0FQsLqvCARfuC8sUtQOOAOlN
i1GiokDOsFpXCRcKwDuYHXCJ55OygK8iTbFdTOBjC2Dvx3023AA+e5peey6Y
QpPbkCNgKr4d9wVYzTVSNyZsvdGWlvQT1XPmD5R6BBepQOFtjkq4TL3wC+dt
CARARJl/rOKfwKk+W6IZHAyIKeDBdukwr1A6JbG+rg439ErqdEV4i+h8aShJ
7eLULQIj1xPVXTi1sFLBdLn7wBHuqHE7g6+KWgSBAV7PegGUATHwoSWhZVqr
/s7pVpmxKcgh5641F0F/L9WqQiNnHhCG01WSr6z7Sz7uS0qzPD4mJhB5HtFZ
hU3hDVX9HanFPksc2LJi5l3XdvxiKqhqRKlEWmmAcm9k/uulQ55QuaqB1Bmc
4CU5mLgwtWh54h+6KIgnq02pUVcp1GIaoMV50o3F9iW7OS+2tVvczESJfuiA
3jyeUXnKQFV+yXTL6n6pYy29+ZO4xmgjQ93QYGCkWo1HEf7chQA5b8bOnhqw
9fkmVs4MKINCWzAMtSh8QsEb7/cphG6Y+DRCGoiqYprBt1a7qmERPGKTYlTd
BC1sUZShu3tlr9iuE4hH638eXX+NmWcc0VBcX92YTP6GiGaSO46ag7F5PY2o
wxFhnPruZw5tsoWn4Xdm1qBPZ6EsiOpqi6+PAooS61/qyXG1qUPz5Ka0rOeI
1d8dmlbJ5LTD7GQsvLJXNHNIyXrte192wv+0bcTN6b5jXecunmyUFLVYflO6
/mhja74Wthtvwe1iIBcKgI1FtwPywdfQhjvDlqSfC/uOB4KVyw89zo1xI1m9
soJqj0KK9KDGo7Ole8tJsoF2IND+Pnt/PAAqfR3gpqZEKIu7qI70QQnCTEvl
Lvi+uIyWF4qTXIZtUMYUj1H4cj/1y3cffitQeiBhQOxJE+/wlZ8Fr5IOASg4
AmdWc74OZCN9y0CCq3PzPjLXJG+KlqxLa+UMSNW1S0fTMQwbzijLAlrbzQuN
a0y2W8AEJ6qf8ealHMjd4UgLJHYs7D8qAoHJ1SK5MO2Uie8ljBtWd3QD0ln2
fTgLKrFu0z5cFqeedTUgTIkMlTLuAWS99qvjPiz4vnKt/SKPaDYy9eJHy/yz
BM5aegdXmQj36im+XY8fZOzGLzrE0vqN9Tm79vaZi04O+DNW8mcG15s/oECJ
27t1pnmFFtYLADAJ3oE9iyF7fII+INDvdwMoqf+wUW/7SDX3yu46r1rfhsrS
o1m+2efu3MguNsVNscFRxCKzUj0JXyYK3Fl1kquibSigZLc7uxghCC5hQd4i
TVAC1248RrzKvm51GQALUW86IRygq9eC3tDNwgQhGYLO/8h8rv4D+24v33yf
hnK0mr0CAhPnIZSd0BYUeVqNFJKxbbDFellQpYufzM8J+n9Lbti9FKGfCCCT
IFlPTxVpcX/8vafmfoOwPM8uhBB0cBvFcJTQG8/EWvyXnX1CY1VMcFobJfmd
DBdgBbvmzngne+6LxxJ50fCocJiIzo/ZORKppLJS7FQktofcgumKLMjtyHbH
/kHfHO/MSrFC2s1/BPqcOYvG3laMeeOaXS7RJXqZZgVVCViXbab9GVmnsRM9
s4rVZ265vT+QvVInakGUwPy6IHnAPL4+ru7NvIbYob4pWM2tx/PWhs9Xghlw
gU8IQRKkynXitNlgPcxMojNwfNG7FfGfbVlONVzwy5d/gCRAGjzaqkkaysSA
fX2IzC1RGn4+4KRwWEA7OFQ4o+x0bBnAfcwxnwe0r1RAZDATATKgIaY04QEB
X9XzR6ZPPfLx9dwhfQ47LxQGSrLG67860DfYo1xR9WsweWRbheg/LK8mDCBM
iHZuLKtR5wnSy4FFEM7XR+uvwT9QWznPAxLcXLe67yjKEH1pF3HDKg39RR2F
bRLi6kMqT+CFp3qxDBPbjg4qxBWWtez6Q4mnduKm1/gkuglfsDQ0f8Ht3DAc
OHTT4zMcETEQve7lnOgJOV8Qp0e+x2St5G1dPI7tQCBXLQ+wcrA0aNg9bcpG
HqCgur8BoXBrPICJq4XjWxyq4an+RzpsTcSrMbwOamvz4XQ0/2HkWAEJDHhO
yGBNI6WGskMi/VSZ4H+d7ddXyOwRibcwve5PoOrV1pnV2LsIVJUdy3Jcd2EY
bGoTg6IoWHOAjh60gsviQ8E33M5THFJLdJMTfWacd4tAHO6KdF8siYDLFti5
gV9V6ge7Luh/L3EhKlJrZZEdWqSoUegrNJxn2k7yjj9TL//ypCAUXasIx/Mc
73Eto/JA5pkstWk50NQ+QG05R9b1RrnGtIrgcEfub8/VNTTatVLAMXtlHLsS
xc12UsZ9HnFAYQ4WSe1aOWWryooRxPwl3fO1TX0+d8Y/bvvMr3xwQQST58A5
8cJz+tDME2bsplyQZ5R3iULz5/kgDq4knd3Nfebup6WfDyl5T+7b94cR2rR0
z/o7+PLoUgVkS5PRQ3trllWPU1TcwC4qo9i8lqnSyXxm6hid3LJcebZN2ud9
scAaT/y7SLFImz4J6ED3YrhvD9Uy6XuxLVYTxSNG2Zb0u+aR6/L7igyr5K7w
ZaOtQoWiOsJBO9dqGmhMURueDCFAU2Z0PnIaVOyoMwyGnqVgoNmSEoSNYPQp
13jzuXGq0irlv+N3Mc4S+JDo3sz3dAoKz1Nlge/1LpF5bVcchhp92trSFhJA
J1BjXuNcLH8mWza9NVUqhwJ6Z+PXhTUyXFcdsS1sPR7KKQBeVS7W40UbyLw4
843kHPvYIQ2Y/3B/SMQvdrlNsQFunei2fwbPIllZpcKF+zAd42wDtpX2m/sA
Tmv0wo6n5jx0g0jhKM5sAVOJYd4mxYaI+yV23S3+VIXDe0a1ZAijbYgzxGQ7
Ws1b2BpjYftc3f+kc2eZ1L1ud3IJIxjJfUjviWxfePrpRZQWnoJXAuSCWEKk
XQGdnwn5Gikc51SwvRh7QL1WVAxJWuxITLDQqyB6rnAET0P6O2LSayZ3SeKw
HHdatg6F4wHvfHZuXeUbHoVPZ+LvFLXcRuxHdfZaYFYlglyPK+EIO7rAnnqA
pERrVr+723Kezu0rCNamb5cbhEIF65vk2wsTNJPePVwPl1CCv8933rlwhHM0
pOzZEUrHLv/HwoYdIsYaillbmfj9ZfuQTbmTOqUMAvF08tmciao6Bp2C++Wt
vQuWwmUy/zthfmVH+3tdNVG6m6Jk+GBGPOhR3ky/s5S3Ga0vf+YKuDha30GY
Jv3tlqNS/XLaup98jz8rA2JwOCaRnQJVP1cXSzsGagKmvmB94NSm1Cv1Qd9p
hCqneQ6driFGe6GVanRBTTLAnZZeScBsjvr+5bCPFmXlXLCBPR1izA9WkzDe
M20oY+zCKgnRtNryLoTEECdciBzl2H3JZgh32gaL7Xge3laVDAimrfTr7xdo
FkIJbn2a1Q2103uCjVVU66p1Q6SykH5VZza2Mca7CNHitN4bEPgEi4MFL3xb
N4/AEBHDi/duiOHW+X7ECq/emgI22q4kBDovKp+TPDZVpEt1ESwjc/bzj20S
6FLWnxIfGxE67K2d1QeQlspVRnzzYCzGZK+CM7eYngDjiEgvuhy/JiEddU+c
w8WT6gP6COoGSSWqqLoVM5vrFOej763CHhUdOr17X2AiTQ3Gkxy/XREfE2ei
Tkaz7qWudbU1/cwQ8OuhM8pW8R8M/W3Fnpf4qJboQyw14t1VSoe8WTZ8XRGk
6K1lh66aE1fVCB+SgXIVvw+Pmp9ng8QbladTVtu+jniWpZ/UB1G6g33J2wTm
Mn0aCW0obPC414OWxJTqRKgrBBcRUia86+E7/UPNszbKpzfPrrvJQkmphpUk
iEvGGwjS/adoO0Vg9qDJZWdKyBVnpyHoE8CKpF577IggYy2cPDfRkMiQ+97K
viENHqXa6IYYCklxp8dbfkPHXVpDLlCSyFS3RKc+a/a89Hh0nJB3LtJtB7Bh
5X7QdDeTKT4Nu7xHkLvnmmx8r9ksQWw/CZ3wZ5HrPQoFiqxNqhmf/07k5rC5
pP0zrPXnQvqkxCMKSQ57mHg3yl+H3ZAsIBJEByWoS+A94LUwm3SO+wP5rLOH
+Y3843n0yjBbD2TzkJ2CW0uvP+kbu7Q7V67K5xmBqCRdQh6cSm3C5VbNr1yN
5Iq7uE5NqXopwH3S4L9ad4GGUUvSkcgoi9n05oDn+ybSGfIiYFJuHKpi03oi
Vdp3KwaFSXw2S3yTDX2sWviX9W1+1f9ZYMjKICmdflOp3tFrBYMUDfBQhPUx
yYxyb4fIqKQgzojA9UOqvkBshpnWbEx+I0vxTj2f01g7OG1MqfTxHy9FQZIO
11o/PZx2YOJCymZi2KEhFHAtlGlw2Is8LY7H4W2xLwPfoQSicKDnUyyc2EBu
iXX5RmqVmv87bU6N9KqU8VL1TpjC2WdDATljMUPsFZENl5mtgBRutMkS+RPm
SxB68FtgTtChFv+7WrxvQSR/NRCqlHYMcrDLvpM0eOYzYqLx9KHo/RLv1DYe
Vc3hja5G2Puh3DDJP88hWOFCS7lpcLF9J7Cz/4bgmcnwB7LW35Vt8JKzZOGv
97YFbySo1dcrzUdbUI6slSj92SYXwAWS63SY2atn4WhBf55y5NZNaqgWMWKm
hhzsOTzkxzDm4pQMwPRKA+Mz6AjkDK/ox7KerIXvtW6XmlLedgllq6+2MBOD
9ntv3j5J+Xxya6gZKmsLmVyOC2QO0VMNs+/etHEDy0hk2U9kLV4JMiDKT1WS
LWnyVOEXJhne7u4+1BA+ipSfclLOB66M9FXVmr4PnSNvxBoGbsCE78d+FLCK
tkAVN3PpyWE0Wu/9qcYABGu3dw7/Npbp68HOYIhuPStngz4oQ9Z7kklejPJY
U2fUBEaStO+goAXUFW97Oxpeuqgyd5FWvochlj16pwQkxHFdD0tCp+zKQwkN
OTzqdAhSvQtRaw79hqAs6Bp6y8k3aLp9Cg0yHb/XF2GHgqnzjd2wxRxNvUMi
O0mrRh4q6RfJqzzFGMwvT6WFzlAE5t3o5ihXR0YyQFEyhM69fjqWG+uCh2UV
8eXyDnNfnozkscRQ+nnzIr3yG+IUDFFxmsTeSXZqCEHNwJFmOBp6Kxlf2oEx
RNxLMmo6wUUnmlEylA+Y3mTZoPNMhsuGyrekA8bizmBOvK2nb2Hly08jIJrB
6EvD+8rmrvM4M2pt3jamFGcSQt+2h94Zbag/0qktyQO3bhXU+RRfltAo8+Ky
xDTn0Ul7W4bx2U9C+FsUAK5j7OZXa/Nm05yCaTNfwQzc9ecoO5cufYXofUZ3
kRC/OY4TM3rHNRm034cThvJo+FFMWoLlSS2EcXnL00muhVA7ANRWYGGTeaT9
WVNsbZpRvOJvxm0Tq1GjxJiFoQ/vbH4mSmLUdXxR0l80KD9eIQ/Dv9Mx1Cwy
6KDdYNspC6m1f7OBit0DZQvZdDJ+kVNCHUEGE+/V0gCxs3X7MjbFR/Q9Od4V
9+8f2jQSbArVwqRc/kMeRSfHh9Admb1yqkKSV7YS4hnrrtHB6qlT0LhYco4C
G+DiQy+IMtXdYyQV8tMZxWFEB6ICOfqRhhm3cZkxKh2FHiEEDpIzVe+gvY5N
o9AHg91rfJP01cH+JEG9C+2Tt/YKR20GCuve8jA/tKVhcoaf47HuE5a7sEgm
f7B+82sUfFd0dPEvz1amhuSN/7OBee4G9MuWfwaUGv7SM+DOdoZr9EpgUvYc
zT6bBKcjfqRQNDNv4Y1X/to+odFi3Vn1sBeYxK3sZpOesjmeXdrz4v4Rfbo9
RYg4B1LWSwYy9eBc5xAwOWT1rRLoaSIyivC9cZeiz9+GLOb1UacGmUa0xv3m
faj6tn961FbFTSnCOOLF5M5McqiYk/GEV99QLVPn39fte8xCpmsLCkKnojy/
9nwFL/zK8UzLSuT9bGD2/2+TsYyDBA0PxYRzQZ2mBh+kciNu/oN02t8Y2lb/
wrlFGpfMaCpfwAkd9ID/FD8TlrJJVP+QTxv4aJAkMN+NNMalT9PUQ6KyDzTB
EYNjQZaFLPausa0Qy3/dv1e+5V71Y37b2nfx9uXA277twngJlSbLiREtn0Gs
L22y4AAAz5ZiMIF4OJTwPn751ADFVUw8B8Xe8tF65XJ5JLOytyqEGEdcRAgM
LGuF7hR+2hD+i0qDib1fVKlra5VAW6UYLJzx2bfbqMtFgOqdm+cefyjofedN
ygBWu9FwwkLY0+wxaUcEhNoS/LYxvTHz2KKdQ04CM2LxjCIFubFCR/9kBB0i
iWbjOccXRHE/6O8ujhoDp9drfuSRGBJ6LVfPRihBL02iMjub4kSKU/VpIuP6
OsoDxCyW/lrvgt3xYbsJM1Ey02Dwu2uBc+8lM5ZZ15WT2ITbQbTZkv7ezP39
o4ADCNOG6ilCmZzU2INgEBiFt8lYVPLW/e/2sKE4A77vFWwqThvcNzfPMXXf
eUy8AwPzaxXdDD06UtHNT8pinIAySk0khGqHNmD7QCQIeuBRui/LPKcch61e
7mdz/kcPKs07Msb5HAjphMshTchrcSzt3aaduhc6oWqDfJXq94nfo4jWsisA
+H4QNnn4C8UQdHHIGZqlc7AYuBUbaVWJmdH7AEilDb4yERmrAbye7UOXVEwP
/ZzE1YLP+yvhWWIf0p7/UgR/6Lh5LOSzUoaqt55Zpgl4MtoJCS33ozCmFFmM
SYjMRN1fpLqWeSuHSVX98DJCyZPoAuu8pF+2xNLxSky9Fl6sH27oKGFIU9IO
aZvbajW7v3mD9PCLfzxb8Gb41jyW2cLwUZPZwcqx6OzA695JZiXv1dKX2XNt
fwXsYVOBPmKiThytW1yOERihKNmTcsrkKyvj0zAB89NkE33R6UwsgOLZAGS+
4su/ETP8BP6ZH9NYk6KwRdG5FzJdfDbS0RU06D5af5NnUnVjYGYwzZNGl9oM
CNdi7n9HIoRxxYnLnkFiJIGevz7H9Ub5VKtpbZGIZ5tCeuyedWXkPvytkOlR
NPZiQgD+xsZ5FKGgut9D7pfVE9QmaFodEqVOfzlYeBQ49UzD7X2KaQtLD/MP
k9ZrIZ8SU9J87S7UJ14K1BuBZV4xa1O680nNhJBBo9W1iA9k3UOjQ5EkdSs5
Pg0gsjCSK6vketxKCV6/CCNtg5ALpZ1M/tkzBCHt8cYELyrN8bkyDhAwrU9/
vl1rf3UkFQMtgWKhfUpSx8Co6IPVzWG1Dmxt21YdWl2nTknKvd5TPb3/OLI3
0Yrmm31PpZljQIYFobMiNHHXE+vSx3s/PxcMf32KJLK1zlHjy6G+vTFOIFJ+
P1Civ9W/c4sYJrF/x/AjOnnV1vv1J8Ebktn7kxhN/4p/+MuzEVQ7v8jBcY0K
TF54gQK0vxw4yaD1ooARBhr6OqzUF8sSl0C0w7TwM2GhKWrwcix18Bifg09W
p8zv5pE9ylK3z/9a7DhvlCQBzb6bONw1mv75pYY3tefxJdac8iavwCvnEoMs
xQMc6eVdMFU5kPCtE3+fiQe35rQ9LgtV/b0q17zi/Dwi7jLPjM6gWftr0jJL
TxisvdpdXXSFN+eeEBA7/WTigQU4b2Tm0GaWI4ivVIAWC+BVT9EukXQY1Gec
F3yP4hOSxuPA4qarn89cO1jkrQYPSnBtJ+a9uc+1kL+IrWIkF6af6X+w93fg
L57+wFtEVDG12Cc1vWfnZFsu8eXEZd7Bx3LazN8fL3TQfRmE6O4Ohf6x11O0
CHM9tSBvvWXUfG+Vt1I06YG8t91i1J9LPcfZ4pAga6CJO78fLJMi93OJ90Jz
Ww4K5lYSSBReYgN6/hPScqRJ81sqNJwc2YMzB9RnzVZCim66VUth2BiILqJk
37+YbtxbnMPquWT04Godhmyqn5z3a9JGt3oRlh/SdVJOXdckiUqeEISd+6JI
H3wO9c5/ms1OcJR9pTB/HOc0X3W5aXJoPlozBSVFs2YO8mYo/DPlCG905URq
oG/XK+WROYG/xhXCpC+MA+DdFcLq63uan2tYzpk+elZV7v9lZRs35irEFZXB
lRxBZWQKx6953NHfkG+PgmItOrmTfD1PAQmDNpbEjcsQ5S7fqzzMnpcPOa6v
DyuCFs4sEYjcgQsoybEpjM0gY8M3UavxF/e21C2aUzrHy3Ls0imgLZ4A5n7D
YCV853FPwsdGfIJQWg1OH48xzB3BHngCm/F/FFa3TCOMOTGJqmsfqfZpeQy2
KE0aq6joRr1nQ7cgqlWnCyPYQQbP8zPqqs6Fnz3XwdRmzIn5ziJ3dOYBmMsI
MEMuX/gZaFTpyfGBVvbqw5z4XCvXqEFg9d1gOz7csjOPgItPX53GCVHByojW
NwLz5LWP3wxAkNSWe4VQqey70RrA73JBkD1Qk+Yx4HafYKOsAwNsY5OkfyfX
/ZGWR32NUvquL08sWGcd3j8idJawpi430FJeAw5i7JsaTGfV9XFQpUZy7kqk
xI4BqxpOJFw4i/s9AQjjVxQTGeanGnK300A2Z0OMyck6yy+2iveUjPnNQGk6
3tsbX2xUSsXviWsusSobj8phuDYEVGbWgPQs40CA27TumcaSHnwcN0GPKgUm
DRagBJdntA5ppNzH9CDVGaohcMYdun4IgeynZA6rnCh+U48/9yheh24cD8oD
P7USY2Knr3fRvvEBlLgt+3SKVqhMJfkXQ3EA9GP3uozCbENH05Lpas5kqykn
r7leseeAjojdtj4IQwmWQTOOuUxhaqaZfFeirsIua+QhAf7dinMrKktUTnpV
UW2cVcE/juLZ9oIi+Yjd8XbqGF77Yt6QNrwG5m/E1BooP006ZDUSbGfx9a4q
PL+XPkZC8FloW8zM2nvVIHx3qGA6C/QoPoQ4Y8RIBF5CHME04cIoPx8VuA+0
K40RBYqBSFHKB8qsxsd6/pvhMlAO+kDkMklTMiUooX1dOyM0vEWtteIF4utu
NBMrUZBQDB0+0nF7gU7ISqzxXz88heOYPGwVLKH85qRHapQtBBrkZ4OzAlQ3
zQdrMUk2yC9SrPYP+KeF2DJra2/goSWv7Rj1DuW155PNJGZl1LiEwNIRus/s
YkNKoG/IDAI1IYep4/AVgq4FGC3/eVJ1OVjT54K2O5Lyb1s30VXVO0/DJ0QQ
/cBjvFuIwa03hCCO9+TAvGSyGSqoVHQBbz1wUiyumGZl9d+xhxuz6bVh3g0S
BZ/c2H/W8cO13V0M58TneGw8645Ung4hQCnp2eVCDbzsUGD13piEzzUaPol7
CQvv+whAaRgSObK4fdqovKHxkmY4xfptYh2AY2MGK/7t38Vw4u2LEVOjJO1Z
QALzFRdOtd2lSt0GIJ7vzk1CDtctgsKxMRPsspDX1oaweKTlrOobmrA2akvP
1aOya71D1ciJ6bGqw6HhXxTZeTfL8zBb2X0AAMZUULb+dsHHQdqUXuwJ8QI0
5cl5d2k0dcXMWFqiHYLwIZ3bOwLzpocDF0cOYON3jF+48SlKtjUU0+QUw0wR
MFGzn4KIHIQrxweOT3kGsGQiV4Mjs2tyv9aNL5nWLNNewDjiWJtfNuQgFkgD
02gkPn5YiWmuXHQ1u7QyWx4aPA5X/j49iCSsOGhhvEEn/P2nh8HScz1QEIRi
+2IwYErc0n95xrWR6EuMmS2yGR7bS2c4iQ7cKAbqjZz9C6E6QDhKw4kDELST
KW7kJFaUbLIYi+72BiRJqZeibRGjbsvfYP2D4TR4J2GFt/bBUIvIqk5qclAO
H6+NwIbCVTWSH0IfSbTSF+aA3pbi04PnfG4M4FWvxNazGaAJXt/t79vpwaFn
wfKun7ihD7yhEMS2UusmIpCgUMn254dz6+0Y3SK1B42pO0jjxMDUCJaYdJQG
JekmeiSQc4aSg61yEdTRf4h2yDchbLVg5FbYBxiMyE0XbWgZnuf0cNUMr9re
nedcO8uiOs5AGt21v1tGsvRrH8r1CrdyUBJ1jXJ+R26RcxyS9PO2SgqAo30r
5ABzFf0XD8rEam5r8wywzl7asuXzZIBPFmZ2zwrw0OoUODkzaZRs9eg0hW0q
YuxegqRKZf8i0gvtCaXevCg8XkH15/SEoBXLwIM3SZUg8rLgQSkBgu0QoRSO
JHvZaVMdeMQnuHBpvsTLJUyGB1mgtDrLe6GXpLZ+uRGjEcmJWVCc5ekFGHrD
S3paF/vUSu7orkc3sQVoOTtYP+z2RtoZzLeYhmJ/9aOFOuuh/XPuWKbl0uRu
oIVWypLiVZEhPK91KoH44eF0oyosp51E9/8laEfmsCqSn8vqZb4VQzZRj8DC
c+V5rio5VG74pmZwINDEMv3kme4VQR9n3R3KjFl7uaf8MH+X0k8KzjrvRtHv
wBfIx9Fw5VKAwZuhFWmGL6Cro2fd7HPgFMieJZqP00UFwTNJLu8ZILOLeEpv
WqtQVywXK5igGt+FjtoUHoMsPAkMUqLFqnvZ+Jz4+mql3hfDS5EuH5hTmUDC
VG4lXt7U+3Ex0oPpshIRtKaHWyoMn9R4aL3yL7vzYFisIqLj7ll+yF12ldYy
FBfgR7S+UepDOAKri0+GhuFmopfBWM+sxEv4yMmVIIbKIC+VydchgQVMfeeM
HHcMhnNhQAt75f3i6pVnbhbjmMn8z+DAlX26nf17GXbXuk+lXK0KNRhsPskU
Eip8s1JSEaNn0VLYTE0NMeST8dEstfWLKmLNB6IR0WgDeIXFzfObJMCip7D3
ZZ1O10OXDQYrWz1fUD12taLdZK3eQnJhqMle2rpUQsEp6Femu7YqAdHTvhHI
FlpXhSRwzN57L6UFW8K8JkZNVkhLg2IuOVcA7TEHufVUvW/4ys8Hn9X8iu8G
2F63O0/Yrzyflasz7ST7/eCV/QNXR4ywhbm9kAWQ8fxOQKtF7ydfG2A1/Xy8
b7jcPjh3KWeaR1LxMju6qpbqo1TedWxiT0hsaRDezREozBOKkAE9P+hiYuIK
xNgXl5AQ5zfQ99EBSbeWxOjPm5eZyp/lV5yprubcmzTIAwnEzKtKVWtnas73
AQIN0jax1pb+W6Ul0o3mjQ/4SspvQierpTPSADkqiNL70AtzPJXicOnFsFTG
ieS0WVytiUAMfgJE+0GHpli3amEc0IO003VMAoxzVoOq31E+mEC300v1aLZH
wrmoS1T1ucRGlQRSOpxIkqYzkTCHLvx4rMZFLl9pc3HOjGTbWzYmXRpMZtly
fIVPdAnbpRQ1ObCY15slylg4GVKqDbaNIEL8FJ1zQfO8zqvro+TlgjPYIdPs
oMGc2pkT9rW5qGbaQ1kqgHynAIIGby4gLEPFLgN9b852Tlq39VwrlVHcKRRa
bQz1Qn3bhRjjdC0t/eeGsAfKN+IIj/b2stYher7bOQxNJJ5+RGbgAhdG07SW
QQYKAJevLD92MpH7Bdspu7b2+VeOAjhjjVwmmDqMAaCimZ7pAUSyR4En/O7d
PJN38rHgNSvjsTDaE3h9gCrc8ON0bbXzjeDvUhxmIPoUqZLUJMdzXTjqLlRc
mNxnIgXOiMUIEn52pc+1u/ji/+iEWounAa2OxBR9nDj0X1KbKFw0teE+0FJ3
CkZ0gVy8Klf9pFpsjk2xQgbKVJFdGMU7tRgb4wVl1AgXEC/x3AOcFazwRo/9
G1NDk6+ftwBUy1QO/1/I/UO+SW2//FNzJ0XJoBDzpyMr6wRaQ0H88j43s6/4
2RGw1btxBxFDEGWDgAIe/yTglA4lIlecrji1OAe4WaUzAYcY2iE300ppwUQV
Cs0Uwog/l1a121ptW+sQ8Kxj0a7dOg0DU+MQztyuTVof90aH5+8TS0dAK6X1
xCTWTkYHtvY1PYGhUM2hl43/3P70oAbhb/ICMqbfQjH9z3RWwZSDGZpmedPJ
+cPuZkX4y+4lOUizr3JV84gg7KOPp67sqXKgKEFsRz9qXtPVzEkaKoRF6z5f
DHmX9DnyK4D8rERfDQRUc5ff6hJwDYt77GS9QzMizSoO6zmX3fcRC/Y3MZZB
RG7Jw2GXsELw4wisVugiavdn64Jts3xdP+JXicn5+RPsZ9BLtei+/7r+NxmK
PZMtPk9EHJNd9zoinoMjY5j4aJgHnsj9CV4eqJraGGMVG/DXBwtNaiySDUCc
mezGr6TamvnyX3/WxTWSHaMBtxt+fzbmKPdUm9LLk8ejKq6ngbkcruHhkUeP
PmRxzEr2tqDcc8Y8Nk/jaF6EjHOZiGFk90S3Lnd6q+wFwv30Gxa01z9aidYy
vS12Klk31D2zayI6iXZX5yxSkj1CT6AgRqdmIaPINgU8WkwmtrBhwtTT2H9Y
XfOfp70Gv13tdQ7c0ipRGggDvn2mr+LX/y6SbRBJtDVgmVxUgYlPsB3U5LtQ
KglwhSup3+C/5w7N3RKv+zHJbqhauPpvTP3ksFSrkdwPCQhhM8N3sLyIvAOp
rdIKIByuowVNqO85CE/pwZPRmaU6TItS8HyMe2dlYfub+lGPL7e+hyrO/xgz
/4/1wq3BRBQoAhTDMNOjhAKgtNor32kcl0tkZcA3L29mnyNMUmMPunkE66oW
kj8OKNgi98NXiP6GaumwsEHCqelaybGP8J290nXNciMpCKkolHZJi/R/icjI
Lu7yZfvnsJs06iwxIClPNHmAbT5Czjvh+kzXS2rKjdU/omlixCHro/GUQcvu
FFxACVMqQArTKmDjmLLr+T/TsWmAF0eTlqIDWL8VGv0iWEKyo7TPLzPu90HP
aACpCv9M75+IzfZ/xOR/AYURKLKaFRbqvdoJVwhHVHSKxRnKn81gBa9WTHvX
sEi1U7QX2csNmi6/02vJ7C96xNxlvnTxnORZ28MKzw+vqLtVFLBtMqsqmXgh
xByYR5MzYupdT54iZHfhfMu9qr9cFNPau7Xx/pC+Z1rEtc8yUDJhS3I0soet
LouvZS25Ib9/c1HjEb2xE5D6PQ/X4mr7LeLpa11Xh6H3I3aNnVCWdXQfmK5p
rSj+p1RKvvo6SSm52uZTvdLwYdNRQnW3CiRLeOLA6V/orZm23zJGczgKKMa8
d7hpkwEeU54aDVETEfWAWWj+5XX3p/hIJR1/7kc8pvhnZtD5xPFy4uTE2x0r
Xn44usf5Vj0o0Kt+TZAe1dBII4EMN8qxm97I66J+F/yJZxRuW23gNHOnfP6I
mALu1t6349Ee7QP0x0Mjy0+O6LwMAvOvBTPHOC/HLhFnQUYKEhfReB85U6dv
Bzlzk5/ZDByd73XTvA+ERgauL7+nJl035/LqkbvyYaTk8GAfKF3eCXHpjZ6K
z/VLBfDhW+6pHz/kxBptgJBHbWZQhHskQdMc8LOE5c0+2scwu6TK+Fihkq/B
agVymn5IlxIgnivSVLim55JbrjkbN/bYFPwIHPaA/wuXwURo01qILMCZStKD
7moIEWmQeW9rEgP72dq5OMH2QiOd1SfdYpC1k2rinjffSjiSSH+Sa/141HUb
SinA6CHsOiLQUiiRKwcAoJC1ZDINg7dL3BlNpu9toQ6HmPuigjCFWqeYzttV
Rn8whyywtflSdag+cFI1w9WqsViYNDkWrYLmQ3prrewB5m14eniJ2Dpovd1R
PoQeB9apePpEt6+X/edKKszho8M4UJlemwCWjf7jVMSl4LhdgbQ0bCsztlQx
YAF2bfCxQc4eIdPMDX4YGprsCVfeyVVHxt8ccSAexECukHes2ygSMEwE8wX5
KVH2arQQNZ1rcaf9tPpWOqRJ3GkoElfM0PIFt4xdwF08/two0BZT9Lcp0+mE
stB65qIPwa3XlZxS0DwCSQ6J1YCO9Rdjrd5re5SGNIQmk1x3SPlUH5zohAUF
6ZyvH9e/8uJYGsGOo3osJSj8fMllusL38Ibq7l8Pj2f9tY5Goj1zi5IdXW7Y
cbYbWs9h5aG/Ohij7900+LJJRelevEuDq2WfmkXF06ePNF79RcfqE49qKzl1
GVE0ixaAT5HG/CC7MWDWCNU46a1QzbUY+6Dn4QetXOqUXjGxgXr7Jpvq3jcD
9GxRf7Fe9niUlDcPox1jhyd/1D6YaszeoUJJ5acFI8+rnstrfahVTrvN47GJ
XeJTSSMGMfwrK4Y4SCJGb+J1NSzhZxN5Qvhb2Fdpi2CpcNEFEpHQJnNpOiaV
r70ytWvdS39hrQNlm92i0v7pg5uaBsHUHAyrQxUb03slksh8K3jisquHHsup
yw5RUZkx1zbxUl+hsNEdenIa+1vRDBS3uXWK7tUy1ar6uPpRsm9XCX53iMBn
BrESbd8p3WRiLPWszIWbkNxG5WMCw05nQFNiiDU5b3DOBV+j7fK9tur3BY+5
XOXDCbMGFvHjEdisu/wESYBrH4BXBiXRuQA+/MqbQVpcsny/C2T1Tov0dAvC
EKY+sTdHk9h+tYXZhvdhChYUCBeg0msTNEGk04PUUI5U0+c0jIsF81ybR9Rx
BidLFsXFg8xOeAZEo+ABioHd0YK/BrmwcS1DUvwj4h/AghvWUQFppKEWjyd8
5ZVeirUUpSv1C/JVLlwnJ9SCbSmJGa+eL3cXd7/ptmFv9x2BCbpF9DMNodTD
9e9ED9RfuMP/ej+5rArsniiYLF4Wo0OsLRlCiieBjcvOLKdo6BrZYOgsR4/w
KynNgSWEp928a5aXV7H8W7XIo3Ymz26MzBA+y6cr6FLE8lUVxNz0K9NAcUNE
ucsMpNk229Ern2w6B/1mvcmXc9DFnoSM8sfpiI4KP7Gv9deVta1wlvbjLIGl
kwYyeTD8cphY/WSuKJuFj0AC+dZWFIsaX7440NhSlMZh2yqL1fpYrCqdRcP5
NCESBDOBls+98DPiQqTHwUjKfPtmEgOQ1u/toqVGqRScLi+CdbiCBp9GOALz
O+2tkKjQzAH3TpXY2LDLrDfObuZtT3rC33pYofUfZwvJyvBhYHi6h48inaAy
xZDbocnfV5ac2iHuMUGu9hZx77Qs5TTr+wAxn6uoJqPHSIt8doc1CItxqMjB
vso78FcnIES0s4SX6+KnCmnsogYPoiCaX66ipBlS6pJCbM2uw0dBNyWJGfWw
b+gP/PXXwoxkM790GLSEkDu7Bl0p826uLDg5aTewTCwb8TEsN0QV5/fsP5Vr
eXPwsej6SeF0NIwyoAPQaPJORRDqL+53lDnUsYUJN3x0m5mqeWDGtru4XhDP
lQxhiSYW5fUecObZ47xMIRpLffIv4UrEbNpgQ4sLbkraCbLcBUBKpvuH+Okp
UYbKW0VYgVW5k0+su/K2nxx2LKSrCDQaZjJ5/0FoWAWzW1eBVzOx2ysWOjgW
RuEG7k99Bme7waQAx/nastqNlUcfjHl5pj0rSKJaUrun6c1cW8KRJEJIbDTE
9NSB4lbWLlZAA8PZZ57Le9rxZO+CSurY/WI+OTjEUMjj3q5Q5b9FkErys7Fe
MmKp49Sj8UqYLX/a6a8XlfF9QltYENNR8Wx+/D8z/cY4Al3SyT6QSAZ5msil
fuvpBkaT1Ki1vGnZsLgfHM7FKA0rn4RM+aBocC/eZ3jf9Lkc6AfXslfvx0hG
vCNA6xW1rwfok0FMfpHtQm+pBz8LB0yZeNQrB3DZeoj3+5EXMffelzTYR0R5
xjIsqXZ8HIOKNcJN8hskGIsBWdhXKA1upfv0Zw1pD1f9wsny+YWHzs/Hlb7Y
e2bSQPv1oq13GIS2bWttYIJY58GRiLHDeUKwj6n52Qu2vBb9QPAberS7ZeIY
F5R2zjhTjZKN4avtn1iXcetnRmkEQ4/0heF1BaZDR0SYCbuGzn4oCaA9LDGI
mxgrbO8mLvbhEnmsKkRi9ZVrW/ltpKGA0JzuJmx56vA0kbdAluJVIEBM6uTy
yqk1hVH+/Q4B5jPJTGhRQJ2kedSH8ZdsNSdZ/4iwq0woABT9trSbS4WMktvN
ZtANFu+ad/vsmlqCoPR1PWGi3n6Alk3Yw7xpiZ4je1b5NLoRnhn5nbSvECDi
mUudAxIRH8tK0cshFji9tfsW7ZU2D62npf3C5N6zVYhbT0wryCIjWBGfCSss
zgbiZYYFRVhfMjLvha+UFm4l8J4Jq2KaZcmFnLRu4E2j3B3+l8/emxCutX1k
ieay4N5mcb3iLTjl+MC+gRNKsM8x8X6tXWqAtatPlo1Pm30xK/63A+A9pQw8
vbYrHk4Hk930JyLc5NeYXj3TpcDXeqlra9MAhyERfkJXY6+5ITzUavOrpf7d
RgQJIpzBx/XvGRh2wGE2n1h5wDfmLEbGrUPmOMNHYaqRClZCcdT5PZzxEMc4
MnnADE08f+hcrMxm6HKPqol7q3wzaNbBCbY/LrgPxkNFezrqGVlSD4B7cuZV
16b/067NRq+0flKdp0pJn3Z1XdVCEsGVVez0qGWyF+B65Qk6UJn3jZAe2NWe
eYkUrPTe3hqSfwhwtXiLgOCyh+LIuZCUaP6ZnhM5/Zv5oj/Ga7REnMUT0wCJ
P/8MkW8kLTKMOFJYbWHM5Bywj4lYK8fMS/NtN1q/giKQA9LoC75PRLQCLHW+
+HWlQQwXDRexiHC3M3PrJLujNy4CrLm9dPa8Utk8fmaoHB4pDKKrjHSC4EzG
tsqJSVauUUVCRtmo8aZoLmwdWXuYxA+AF2sO//dY0jKHGihzbYC5sNA5CPag
YqCkrxDIH8tsmTBeBhR7A1vCbw63lLbM5igGbkXhnkiO8726rYnsjUPT58pr
nXyaUep+Dl/BUdiwQFQcBiJ6IBF2OyRLXA+6DU4DeWA/LYcr7HACVuyHkO0b
RkyKit1xtyHBAozqZJcf8yyjHeWYYr11JXoxYdowGhjqIQ3oTMEZ4irLfJ7P
dorLF913PFINe/+8PIhunYlCYSkj7q9XEo9ruMSuXPt6Xe2MsPhOwRLxxh49
XqI+mcCq/0OcbYD9Aq8IdeNvTQJrgXBJXfuVHgM/bQHcOJSyHUKeg/IBNvl9
tK2WVtAIanq30aMEZNhJVKR4vZqxaqGgSBuUldSB/iYA5REyIV70x/Eo8ijd
ePBroJZzOP3VUi3NVM6ReyxJfz0jQuUWJ8EpFZFmKnCHYahWlF0ghBjBFTjV
jK0C2KLOQpymRsipvmaf4EzIvV/ZRg2AdLO/MvUdrnIg2JX3eixZ/ScPbVYA
RGIZpwtQ0y/x0WHqGSO+l2i75Xx2/sL5uiN3XBx8dEK9d9cJ4tRA9mL3XpEc
bHOsAQm8yob9C8lSJjKp1C+hXDB8bvc/CzszjH6Hp5LPMUguwBA4bXTAf2lB
USX9HcJHbii85lSMBOmO7zuLSThlPQXWm0nYsqc07/z4UJg35asSvFWJJGDW
7uz9vVgd9/xaJwcVisaEKI2gPVGxXuNJXplyd1uw9CXaaIA+mDqNf02gKG5B
8COUkAQbCr/Xw9g6ErHkvVLzCTID24/gZ6C8HzejUA+Pnj7kxDky4hUDY7KA
eJBm6icrYgnW5AgJSewOeQwO+pSLRa1C+M0r3zfxZEE1e9dFp+p/1QIQGBb+
weuhjKeenvqUQo0N8eIqnAbauRjXStpj0OSjCPQTlH74+0BmJD5mzWC5aFet
8DLD1XkdzFwTnJAcdqIvHtCiVfOkR14VkWwL9ZVVJ1fIlfmcawkrvUvlY+IU
twWassMi55lDot0YhJ+XV2bKMlhN4asSfvnS0aNbNh3FY+pW+yMlFDggDEPY
a6W2iYekzDytqkN88ywV7bdzQIT3z49jbuZE6bf/PK+a/GA5C81Xmn+EB/xQ
WQaWb6i3MxvRNb3j01ZzZozyKplN9QSkRzygq7GH8BLlboDsCCJBZlSpuXfL
oumFNkKmcri7QIKGLvo2hotvsJ9zEUutWQTl6e59aWUW28IqnDPuxR1ujXER
amfLUSyEXDLPeDg9IUPGH8OW9ngWObE6CXA36RAtn5bj4a7y4AxhudZeSmCD
nNAzZXyoIRNbK9zxYfAqI1c9fc2OHREFKQSl8pM9L31s+yZKiRvui3u4yxmU
I40YwYsk59UTLjWCpHqaM0B3WDVabPn0ws1qFUQ3pxW+3ZxyWUzFPd4wsWwc
8xRYpkpRg9CYadH7+92Xhsv3pq/dZhwrY7Kurm91Tr7vTeBHrdeul8AeCfvU
y1STA9j50no2C/rY1LfmdySv7nW0oU9LR/r0DsmPQvdS7serRp+vzwWeOezi
8H2b74fFCOAVOgRXSCOg8T3vwVYxVG0nTh717ghTTCBV+IN6VyyjD9tUivVB
VOafYG93Xy46iW/LFLW2tuy0BZ3bWGiBe0Z9Oy7tn/5nQPyG/P3fNvSruC/U
9GtA7pggxTMAlFUE6Xy9ut1vZ+272vGbGmYnML3bWXOPZ/nw5qQMFmXQmbwQ
mt9xH+JkKOLqL+SukHc4m6vmmzdOfpMoAIkTa908X4Qhi67p+aJQvS5oP1hU
ykWVCoFUUgMxWziEzUXqXyx1QKt1CGCjGsKJRBv2KV4+as8QrZ/V4m5x78IQ
TVqff6BgyGHmbd3TWUr3BRs2slfgB+3G/mk6EmP7mHqXZVGnSv+3UjgnWDxM
Z+2BzOWSBzXyisTR2w1rp59x0qyUNw5LOdFYC05zDjhDz5eaKUDmtC/0a2Q5
/CoYmhCc6LpIBeob4TdkfTOhmUWyyJQIaBe4RBihXgHBTt8gFrlvw1F9z7lu
69tRwaKuXeB2x0xNCR6iJkvTAYMtpR5izFNIRFHEBvovQ79v38XI/91wwnFk
tPFfp4/WGXDOW3VIuJZ9pFgYDv6Cr+tTt4ha0IMKmu/R/tPPngZf08zZ68BW
cl3mGIbzxU7ehUrUA5J1kGe8+GitTCW0z7jjNuiHRihD8uK2TmSJz/ypNy1a
pMnRl2SyvVot6dFWeRi8gexuadJmE/7srGp5kq9Tit0ICDUnOR2N8/Fv6ZGp
lJySTjNZwrjxZpY3/osTwB7Rd+DGI4NYwrWCZZjV/TUD0IxgJe9QFaR7NcBj
ipWAoQH0817+ZAC1tuV9DsytQ2FPfOqjdoyrTGxaH4V3g1+5rUzvynooxB3W
GzAKO3BmJQRZUaDfIUsUtUyBFNpdOEZxtbrhUITMFrB3Z8XXTdB2PEcPABVD
Za4vxte7tw08FEt9oFCHH8Pi7PY/cA6da6u+kHn5lgzFn7iSPZa9QhrVvvSc
sSGEdfoyz7cCMxErZzAyGviQ2Ot8kPKpMtX/z4K7ezJFVvqCk8YsPHR/DXWC
UVetaVRtpEIrKLnKtEnPuytjos4UO1lU/w+knXO8rc/UfCIHpR0Evf+6Y84p
ll7FDsuqkxrY5DtgVsO749ea/aaOm75piCIRJpfJUkRS3StkskHUTsIdtRwI
hlP0KKVL3eEIwZnZtQ9TEkMOEanbZsVWEx8Wt4EOX+9vKxdP7r96R+W7C6Q7
zSwtBenS06sZHjY3tB5wVzl3L/gLMuUw+KMU2a+TUw7gH5Osq6g5aG1/An/E
8myCjFsz0xkWadpdpNTgSMXeyAT09YUzvQuHBP9IiarX80h+aTStSqta9Hnp
mgXW56zuw+If6ENbYQecSLk6PaeyoYR40EC0lL4b2p+TyizNJXFDPzVV4wLp
j5vlpSWkrGGqu5d/F5LyMXGE4pqOqdTn13Yjg9iBqiiaC9oru4tiinCpyBSN
kw1OfiYXj9pWn+BJKD4dw0/SJn6uTWg6nEhtO0Z0kSn3hMlVTwdlMjsiViAx
ftbD1Wlb4faczen9XpVViTh507TdouF9gUnDtzMgnX+lipy7KKKPiHbDCeYW
TXkWikyF0kxGcaPxk/YHI+k1hh6fQ9m0mCd0eIdV0SmcZ2oKDIy6hMUr3dW/
s0Ltqg5zOnKwC1NYq8z+IVl5WEQ+3glWIrqrsR+WlvJrTwpTGu68SkLr+npK
5ByMlWyW2PuQO0fNpsoB5Jgc5H5l+eMMdQymxywNItifUpc4bNIHgM0O+7an
iJavXYeto7Kmbap5NE7XmOHXrYWb1GANe6dkHtKAp8bdVPMLTLjO89MU1dx/
1gu+JQLLtz8G4yXuu6uM+ZLBVqOhxyyidgjYp7C6p9bSTKl6SRdMmCm/Gla5
hAQ7IwIMQ9MxQcKKIz9pW4Pfr0uZV09XTjbsULm5ryYLomkvXkBWPzJT8jVe
Xu12vZauFtn2ShU35F7n20cX49X9zDdtNnu8aPgccPeT4D1QzCWd9JOxMecB
mMckKzi56WQ1naIsrczEqAne64XOXSjOsTqbZc6WCnHbfwQdUzYtgVkxr34O
ur0sdFzO0WnxUH6SCj7aNyBqawknzr0J6dWqNUFKyvAcjOVnIwsiWGA5MkXA
LePOBk9S4RkFTWnf9xFtI5hn1ywO+v/z0OFyXWoO7LeKOKIEv4QQa9eNgETJ
RJRlUnn77bZ1e+ZLYbz5j9uccDBRE/bTHzx9E8h71+QTeupYpQ4ZwK7haale
9yqfkv0Xnh8LqCd4YbufRLL/wrsXOTbaVO/gERRWwqn7OtOCKL05Bn9W7jkc
V6SyThLqS6H3ngTns3tAxKA9Ptd0YaKLVdkj7T2bhJEhj6hAXoBlyaZ5SVxf
rcckU76h9IYti+/o80TYlfrC4BdCEI5GjNYQz+O/youGLDkrJW31xy1t5jLW
sl6m0kFRym0bp74NqrR81lBYVtgQ368Lsowp18qJgFE+4sAG+2YY4SF/stXk
inxov71191Ybl+ifg8d/zwDLWKNqRapXrAoo8zwcj7lFBbr4K4dEKYXExzXm
oUAG3Yy7zTu3Ngxdr3DmYsocp4UzFcS4kFQNgzZk1K3LFZvIbmBLtgY+R9nr
HVU0kwiskuZh92+8oBtg5YjG5TcXmO1uDglCwMJbgAJIQFvhr4fKmj24y7ik
8n1tHTibn2dmnaoC+bXtWyS0UDA+A0VfP4RLuuIvTaSgw43SjeZpTC1J4l84
fciYFm+TeWS7w+KQXRdgWK1LHghl17nJ2kcjx3bXDj+6+BUYoiFaVtlEoH8M
BuHRSLgWe2baEeO5wgVzDBDmitanlbCJTuWPQ/3jTMjjanj9r0M3oS0MAKvx
SpbdO2GiNZ6moWhZjzq3cUc06HYDIx3MIMq5kcsxjU5lgi3UdrEX6O/jcsvF
02pt0KC1+118Fne6MxACjUhKaTA+j+YV9A2FVudjQpJzF7R8JQtV7r3ktYBq
ZMa4krCeQNUPDsuOTGAQLQtatpi85mh5kfO50N8yU1QbJi9vKhOgzmv/Lj2O
0JrEIwlnxAPIQrmQ0NUpeJB/plG86ZO2hmr5Lz6cEdCa+GL0JImVO6Fd2Gc6
jwBtXn7FlQm/SlX+xy0lDf2zgJE4NSeV1mfr5L913dAxHZjSLTsakqtEcX8f
s9ZJZ88Ot/FhcL7Ue+wJ2UnZygqUOZ42/7VIFZEU0MT3kQucbdwIHTaJRmdg
IvP+0liNc/nidm6PJt4AcFQffAML0NiDH22ifmodDi4SJWLEvLp5PHxi6uV+
t0OX0Hsh6P57lbk9cSQUShF6hsWikNilA06mMuOwp1TbRyEXIIliQu2DTNyw
mrXVwfKCS3qA9g56LG+YyzeztQihmXT7MdO4DWhe9Xdysqe8kKTKyAXIIsg1
ygGHVvPUhhkb3tRMZLydJHQbDwKXe0+uPcC/clXao92lLcmLNQInu8L7b1jP
dwv79z+6lobSL3JKXk63zzG6X1sNzWaTiZM5UotqHcCHqGSoEpFEcL5W2Hut
VDaWvbACLShHqVjo0MeTAf8KBoUAhDvYWHtf4RqPV3BcUZq7hbBFvZ4o1sXP
yNuO6g4bcD2YOwKSe4ZA60+F23/3WnZo1pbifWSLgaim6wbiLUaYzWfM0/tI
LLE/PapHVqCYUKhBs2/Lr+aHl4oXNaHm3G0edE6cuDOlMzxuWTigwxnia63z
ej22/9Xksdw15a2vpwyIbyaHbmyC9EgzRCOPSyaacaA4vjY95jdcP8jBXj5Y
hklKVIUGpPAGXLCtADIaypSLvt2BQQ+/9P+oynODGypKo7d4jXp5HeGyfN6X
V8eiosJyblc66RAcNF7ZGYHrQxvzGkZv2Ph7hlP2n/52FV4RlynlLO3DA8nx
UA/vFIQfSofsoERGOzGG0byDjexfy9nWrZ1136LB9+JtoPCJ/7emGAxxU7Y0
X2dlaNcnx22QxaWn14Fhq7qj6ykQVpKAaZwcg8aHWZP1UBqX89rFiq4Q3XmG
bCCIjmf4+3xOn2ZzURrMOnATNGMVuOxstbCGWl/G5FIlY5vdiwJlHThkMCNw
kVX9xg6vriAzbpHkXaBQjmKM1FmPE69tt/6BPXWuE1uxO1l38ZNtyZ5kSBvx
EYy+wl2buG/yMR5xqUgtkk4NpDTsQpmLR9I5K+DHHZNjArkQHB76Y1P66p2v
4hcgPPxGuOGVieYKJDImmf6MFzJNfoSEULvL45ujqQa2/CifA5v/gwKYX7DM
69t+jqo9w90oqjZmlVWtMas6XKRFn/9Hd53+doGIIUW30azEgl4wangHnTKY
KoWTtePmkIyN++BIXk0AwtfEkvbj7QzcNsvVDl/7TGr26zX339lq/0K/7uWN
wuypUa4CWwMPo6RPN1W7vqZluaj17c0I1Au2KiXIRUeQmnYKNz2SdqVdKfz4
3DgFlcecmZT0TRxGCfUk2n8BGg4j4e7QWR1SS+xjYsEQt4SS0nHidVST9tIE
GBFsMH6jcG+p3d+diGb2XJRuhWTOs5KyNvkjuelvB5sXqHrYZi83n3Krm3HF
ACQ+sSeuKfjmaswfaRzBxSM+4PUA/YxhjfQLBkKRQs37n6q378IR40BS9jqD
xeIc9qmevrxOcm77pu2R1GgmOIZ68V3J/f5BZTC2nKrL0ZxqrFosbGuZHs/o
56ofmOaSFrhVeKT9XtmXFlrPxTxjKhOD6z2GpgPZZaPUdpnbZ/m+Y4xzEEUc
ac/JL7qVbgyZPm6OcBZc5Nn9pimcXbQJPbz7wf1obi6wV5VJLlXxrcHyDvD9
3qslGvB7vpJGqtwetF3mH9+jz30mDaypxbVvbeg9NGIgjdFswi+me8dEfCgY
sgkJ+zbJOahHvrnJP7ODGGOI+RKnoyPa6qNtdBNDQ323RJo4CAggUmgqtHZI
lNqX4ait5+U+e2f6DC4QaEBG7aQGUD3osfZzY6hCvt7Qpp15R+G34wsWINNx
h1UmNf535voVx4C6xKuhlNwZP3hoWLkoyyd4tlEorjspSV8inRuDEVaXVH2t
VlPnCvj1bk83OrdLTkkDb7laquZhiJJcE8UfJniG7SLkp5ZVZpEaGKW9douk
BG+bC7jvZlfbvnwRSuM6M4Xf6Drl6lZxKtLKzOGs1zZ8hqm1LaQS0x4Sn+l7
ztu17Ze5JoUkarTHhz6jnGs5GrLpIHqlTJtdmA9Tz1JbROhlGsIQln3+BGnx
agDXKybhr6VrtBnQMOw+HNFEMlfAVPHYUUJgPeud/afJ8wVspCiWU8wQ7ykg
AdNItqmNUbO33BbfBX90MTJiuOfpAjkPK3WC1IMEg4wP2UrkZ/yTtL98G8YP
lmkr8MfgdoUitFQ99NNLNrbIVcquwQ+rd2DZdt3p+juencC1aficmT5wKBem
iF4JfOEGG4dLsz7bZxKR4tQFVU/BnJr7auiffsa5jgw2h0M/dEjwNgafhE8A
+6Ip0PWwNJMdkOcBLCpBf0pJ2ZiKoskPZ3Z6DrCND0CqLpefm+ck9PEkfNRp
q6Y0Tvpryj55+3ITC34Q5z96wfCOWENx5RVUbMKOc+ztS5xJnYGJD/Ta0MsC
lLbqpOfHCdCNfH008dad2xUuMAn+U9Yfyf5JOZ9cbMZ7PZP1XN95aVVc7Ywi
LTLxreq3it0RWk2JuZLarcO60P1IeChoXEnmFhnwVdoHflDfh4g0vssPxDhE
yuKVIoI+69i1b3OlhA7Kyb82MJq6shzO4NK9/jgpXE+3nB2+Pyo3oJDANEXS
E57RXp/rq1yJjZmV2agHdug9dXh6gjbPNWDtNgwoMNQkTTi0RgxQvrMh0yJk
nFdJABkk7EV2uFCOgcfg1spSkTJTdFdqKyaYUr/rFo49oIjFNMivYNoob5q1
qV+pF3WmMEF8+BgGuDvA2yD1F3xIWBsbM1vOTboTPl0fvhAitX3NDz0ShZZ7
mmuiYEiQFtYQZ0fJgk/c4hiHLj3pnMnmMRkis3zGvl3V1mQ/alYc2R/rEUm6
Uzc05+HprZQGQL7A3QJzU91+vz9/s4WJ51dGIP5ZZLkDrB3oDvplNwXyGDS9
st4IjrYKzx0wBnfQQbJLKQ2b/zSLCM38znizxfjNFJGvdM6T5xVzjjsZ2AKb
FelIWF4kNg+bRtthNxGyjI2/DDJi4U1XL+cTMkBORKGBwxdMxvqSClH0yOPi
oGy/F/izH7cSLkj2IzKCdPBv+A9gA741IIIgFCyGlMjNkpnw+8BmZ8qDwgVD
y9OO4N+x7UY/qfEmBlMKKaSozu76wWfXb7bczImIPYWe+2htu356pLicTQQT
ZIAncVUmfnFdKKhpagZ8Boc3ii27cEBPPYhXNDeKIHjILz4gEqKWLZFXBokS
P5zNfvtuStgtHioiV0CcsNrDYHbnINM75U+frnK+F9wo0hOslbi/vQTne1m9
8jVEaTq/bII3+cs1HU45QyAaE2yIXbbQM5y9aRSJYy+oNips1Wlxtk48Ej58
7LuEmM1l140z+8nlB8BBgwTu/BxhHCemFJKfwC/KH82mJuv+xe5zC67NUaIk
hxttYiRmgP3mODWpaU1h33j99kbOOJlIIcZiN7uDjjgRV60IFL1glu1fBmcg
HlVw7RUE0GNDQiHozcBC16fRN3Rx9VPnholGWT8fcdChWXRZWr3iUyCVNE6j
se9p+kIiJOfvVquGQq0Fl+9WPqAnDF0CwIswOsKYOLEMpmfxPIWWKEsWlAT7
FzwUcxHbBxxDPxEbyek1I+pWPXXsYqsyE8z7JjgWpeVXr96GLTsiEiaXTXt/
Gku4xpIlR/jiZUBXiyYKdI/o7+/5UHizRyulAWTQAiXFALZiNZvu8Z0ctNCy
R4n7c22CDsc3hSFdJlDDZv2MZ1h2a7ndw00BeyyGvuiuvKwj5n00GhK3rxhZ
x55vQ3XXBbV9Zf3L7PEdQU3rhT1gCek9aIa8Bu1lya1WUvGt+7iUkf46maiN
MZPlB8ulx4JBvBwHJ+ZZDQYP/cbgrdTYo0Q5vXdk+si4ot90wnT37aHPGu4J
1komAIwidZQHL5WI1CJ5kmHirK2eSEOadRhVW17fWuF8mZdya7BMDm4AcDYN
baAGktwtTaLMV41KkpeackxN4yQD56LBZEcvcnkngr0bsKB0cCpfmIMZ44Ck
0mm0zAp+cLyNJqWuN+SaBlSBVT32fPvWWVuiDUAbTHbsUEvEzGeE6jucOO9O
3rKvk3oeuTVxUOjpYzHB5tAvZrqED830AuNCmRjBPUVRAgktUarAR7lajZ7A
IHviZLQkXonhb2TOEYrB3Xi335Z5M98qWg8QMMC6dKZIHgisd0hZm/PBO3rz
Mu4hZ4rb27mQCAQcyCjmopjZbOtMFtZmfH+g0MLk7v691j1/UGdvP8ohVTqx
WButzd/g2cp2/e01UvV0NhF+PvSedn8Pj6YdWHTuY83v5eiCzDxakX5QDkvm
kpBqqTacyPHqV3pInFpi6CBLewXePy/iKIHdB6eI6WnUfrLkr21lcCYgc4Mb
T/OkAimChSq6jvSBzhJPfGYGny7U8QwKozIWXM35eW/C1nw3LAOiIHtoz1Pd
FgZwTrKJamYyp0tLdSurKqzQUKpF6Qs6lJftjayrIrYEFOQ4Ryk3cLfSlHvY
pPHFvhUjjyuJkPZoYXNmTWeIegROKmoy57QnJ720sfpO/Pf9718+zym9KvIC
CCaserIP6+F/Y6eWWoIUnBtASVizCXLDqvkna6KRuJbFjcSrahIExq/Z8BOX
Tdpc0jkKD+MoRs2aeJ8bON9nCS8am2xncuCuWPEb+Rw+gtFkXXkIR5Ifr52G
CnSYnaomplYo0plc4HzhHuNJ9s4HKMot6DA084218L5+SJGeosxPlPtMwU9E
5RBGbKvuDJ36ltWhr5W2wCqnZoGJObwC7cdZEhimbij9rhUu3FL2n3IYmz+Q
3JmtzaYokNyy4mkYDJeBRx6owVDpj+bEoGNEn/1hg6Uh479UnBYCRI1qyvcy
AdN3ZXaNSRed7bmx9qAPMtY6YRKBQzMDBvlBG4xSCg7rsNgmdOAmGV4GOV3Y
np8LtXKTL8niAOpTIUrn36D7m7mKgq8K1arLLs8winOGbtana5DhhJrZ5qWX
VWkIdGZc3yd19LbZzioVnjUG/3QUzquy2Mqc/1I0iRrIohWKuVhT+zm5/cNV
PjTvUwwfk2SMEAss5AgszbZ9Ay1Xt6NQtmCU8DaE157XMeE3YJhbhFYeQI8N
+wCDb7ugN66c5E7N3+dRkEKc7XqhAIZy16LHLIZITbetcdd2Efwbio3feldS
q3iSP16W1NxXSYqG6emwiivy0/6WWkUoQ4jswF0D+VH/7X55pOX/7VSd/ko2
B3CDGjCun5emXsHW1fGDKqsRatWP3ir1vVXgTKG7lGIOIX6BiVgRPcCQGnlg
Cts7Sben9zT1mpTtEi25yJGigR5yRTSbeRGawwPM1tzoxQXs3mce4xRnpUmd
ZbkiMu60vaFgnU7Rjls0/5iKy3c5z6io+87ounoYu/MU14mBIgrtbWBCINud
ORmYoWOcsUUSo0jgKibYaTxZvOLoJteLYAtrpUuRKIq2oKZQgUf437Nf2EyQ
bJ+WRQ8enosRZK+FWIOYtEIwuW7LSjlLiNJs3Fco//rR2SqhmCOJGmKkxVbR
vy6znTDcqrt5cwV6YoQb5Xm6q3zj0AZdHXQN+GeWX+R2CR0FJbEjsDp6LC3+
TQB2ju+zrm7tLNo5uTB966r58KMwVaxptjyX4i/7Kxdv2sZCHToLgCq3hZ51
4bz5NsUDidPw/rzcC+MyLhVT6xyzox7WNXZFTpiUdVgmIlX1LBR+jqeey9kG
heM9P2udAmbKzrJoOlxwc9bOivF3gISTMh3eCrAf3+cELMLnDrUkb1xOY3bT
SdCuYr7yMstvzN4d+iNVqC+McCSEmFvoWcMflEvC16M094YFaP55uugSQ3Pg
QzqMKrT++EfJ8bcqwGUIhjYgqIu3c8E+rjMrghtUXGoDMOpkxuF41BsyeJsW
16R2m5KqiMT5n4ZTeIIIQ3lY2Sxa6U0ZCpiqrZzMXVRmyEdjlO9YfAQNSzg3
siXhCAW8UuHR3qu/r+Uiisr9ik5soYx7y5gJZRhd0tS/O8YTZTDmGHBXmSY8
kpoEDJXdl/KgljbrbS9nQGfTHBRBTRA3XA94dIKhETjHk3Hav4F8oJm7L8TK
+b/UXfmCCRCqzh8WoFl2bVgVLsYrpB0uYrYmkfZJlWbSFHcmwh8eNvp2Leiq
KzwkxDIiqqsQGuMD6M8loeDhL1pFBcsKp4znIoaiBMLQoY46wlSEktgp224W
K8S/gC0JznHkM6vEQ5tc6Z6TCWNmCOl+pqDCrMJQ4DE8OYGnAllXjvsMRv8o
Stn9ol+qPhbkXeviJKx38zcLn6/raNZLyKV/6SBZOsALEZhY9Ufmv6kPnm4q
DfLQbPyzgDE8rxv1qHQ8TIzUbKb553XSjAwLPTAt7jCy/fRfUgYTkrthpMm6
5umR5IFtVZ1T6l90PuolXIhhPk/52guoo0xYMzbpyBu4RN+Q+7eObvHrGo02
f6rbUhB2pENwhL7LK1mBi6KBDWFcfoe0RmaUZvLVeSNjTmtNyGmn8CB38wMw
z8MJ6fwlXWNkx9lBI2Zou6CJxwI3NGUIixin9WEgYzr8JbJVGNQYxD46oJzh
eY2oDk9EC09ZFOwAVlYa0tHY7wjVcMnrC4fTAnC7cJico9L5VKrCknxBEvkH
k7FhsePFxIVMXmnWLbq/eTzYDpVoQijyEEtBTbvII5pk+zY2gpeelwenVG51
T9lJYQXJxjojzKpqrDeRRbP783JOYy18FVKb7eZ/67taMPwG/aFvWEpOo9NF
ceEWMM2R3FKLqS2VLA94cEzcnDArhr2pNwuwf0T6Wq6qeSG2yZo38mM1QcHY
ZvF0HdZNpESekcXgb7S/YFiCiBno0TD5qGlW9no/6bzrZrThP1lHDJ+ZLDZo
qYRc2Q6QmtBoBVTXnVrBh50b3IOXpa8FnIrvEsk+59rS1kmr51hPWIEer9Dr
dtVSC8UKDaYHAguKQJNlViPPrKyB0TDK9DHWjXVaq2ZUZSvadu0PrXQuxpw6
HRITRvBts72hFCyKyrwgup46lwKFjmu07lW4LN4vF6hMabI6qWgERpxdCSYF
oKQEIBmA9DUForUC1MDgIKwLuVKBeLcm+A3smyEpT/4k8Fvkdzt/7g45Rw8f
5aD8BFXu65jY8FuGumtGJEoyqBx5pTm/gHnnMoO4Qpx3UJJwuqoL4FQiWuu6
e3JckTucrbfj4LFwHIVMb4kI6i/9cVxj/BaGGQESkhLs4vLOwb2iobSYDcrA
v/9YL9F7HceE8551tSu9AF/5/PGNB6dnU/sb5KQvTaf483MwieFERuNYIcuj
SJpYGzPvSvi+V5K2q8uTa33NwgjkwCZz3QCd6kZWsDOdMj+J4Xfbx8ucN9p1
T+BwTEzAr7H+aHEuccvRT3PU+uaosl/BXzeHYIbQc7EutRH1TDEyiEYOJ1wr
+H0yhPTRggbtpm4YinXUFTTyni9ePDPmyZGTAJAednKSusViAGyiqoExXw4v
kHY7TPrfrcdX5/aH/2qzPhMGyqWEkTXmDYnzSs1z10Y9ehrJItxFJOIhxoFp
hvjM3VHLDmlnNFq7iaZ7g0lWdEw/72KeYxNNqRfiQ5tQXA7Aw36R5rkMhnWW
oVcl3sEa8Qub1PyhNrZi7aM09keZEav0/1/Lk2LbN0OqzpUPQO0x34clRdBJ
B2yYXi0yBjCLBnebUbUNJyjNGKwCTA8A8kARoOZ68H+eq53rXHF8wP7OUHTr
fjF7LsvzFWvFULfLLxk58y8fC6F8B70HWt/mJFJcx45KoK9jSV/WD+2c+n7M
6TEtL74NIlDyyEnBa4qInFuhxrv8gyghLTc87k2ZzmhzGOGofVkT0xz64cIE
NTEQDWbn/4iEGFrdg4BVPCiVe1kJSZF3kGejPE6wqfUdM8WhPOTuuL37z913
E9ybhZsiE9O5h7XlqdEGOGUBDhtWG+KkuhTzcwWe3uZDhlaQN/idD5gk14R7
kbdkR/QPnkS6XlvFb3ZIh2bpLPl+7i9/UcIea8id9NBw0bgDwlU3OC/tABD+
Ix2FIKtMrHAvbIfaiU/4jM9ScSQDHFw/Xlio0g6pRdFG7C9PdRWcsMdvyaEa
2SBacWgwtNYGbJpRTvI/8V7j1iAvdjx2RwsGsun0ZDa33frrzfiXGL2F+WOS
9Oh+Er9zNofCGi0SfIhyg6fZ3kFGvYFgruFxg8DM+nJus2+I9i9rqtLUrtau
Ct4ytjX7ltOuwrAyya/ic2qUDMSOmuzNyyt7iJBSwBnpxOAsWQLZ19eqzfxl
7NA9brWJzTt+rjP5lLVpMlR69p+zov2NREx+h4d3nK1QuKz0PtiKp0il+ick
Ws1XE9ouRt4z1DfvvU14SfrXazjSz5wSG4DEn+aZiUBnA/6JUGWGB0k48pAo
071JCvw0fVsLV2Sj0FUeBw7FyIj4NvY7tTzl133x2KToLFHUZ6tSYglBqBoG
/UVVYiQ83tv9lReIvCkkEj9TFMOjNEGg6VLwgVVebt+9UeCSGXu28WfMo3rM
CSCEaisgcxVqAV/0Wr2GrT+tZXah6dr7MnG1fkbqwoenYHwpxvS2lhtUJxwz
yk5nzN9wOxwgBVmLe22Qt0OGAEONLmju9tIqQU6QMxiF3lUzh0rF1/MlDgd/
AYKfPkuo5/6mb8rRtMTE97ZTHfOPsBssju27mjJLzGFTZGPrVYLJLhqBoUJ9
Z9b2YzqVE3lytVubPwlJHSUJoLfFo2nvF9qxyn61wGWbCKeB9GK5NRPb1GRC
Ag4UA+WhVmHqLooVzqYJ5ZTYukRnk5rduvN7mR+MOO22AQ6sv2cudZcu+X1O
ZWlLdz1GHSMH9f2ibEv/pHYRRIIl14Ip09utBOmElS1GL/RlIWgYYF0g976d
gwVouO1hxNuF90NA4MBQCasbeTE7YMiZkNVkDEF2wXGFhXFGbno6y3YNUOoK
CsxP6hAx27/0hXmExeEa7xNekSGhztpn5F3y1ZH3BbtzLnt5MY8bVwxbgGfH
8BI5BitVrF0Tjll3SYgJySkxPWEgdMhCX7HkMGbk1DhmLQO+y1vk3hVG/IIE
VsLmPQnHjA3W16FmhgIYBoD9dWkFrHLz+XHCKdbLwFWrRspPiPjntOIVtGKP
oRMwMb3lNzqKjsOB1+gRmS5hECZwSCYd4Uf9WM88uwIU281qAuqlmaE33Tsn
6C4BW5hQ3s0ed55kHtwGr58+9TnDJXDYL8xyFIjYD1WwCV1Z0jjEkdkxfOAV
5lUfZNK/+2L6aV0lZgYvwVHw38hm3B8CfWWycEjuLW9BRDLa8eyPTrUuuQmz
BdVeGrUW/jVFowHLWOEFGAKud9ynXR8ecZXTCS8lGe/Ap+nWYFYXgr9RfBc9
pmSGjzH/8Iu+RLzRpCYATwQzbiMHM2WNx1IGdfxBVNSJi+imq75hGf1+kK6S
MRuR/izg/10h/CmOAV4FdWnwcSYWfP13qzn3VE2GyowWBlF58ttsS4gafEJV
Syk510nm8N9c52bnCz+J/nvMDXuOEDAMs69PkjjQ6XSzdMILxmYoYWDvBqQs
MBLfbFNL7riunaH3zYbXaoj96vFYSjhJh9Eri2vKC8V/sZtVd4Li8+MpfS/V
RQ6d83g1QXwo46TkHXfRyX1OaV/DogCDBokQuib5W5mp/hxsE5rq29gHyMU1
lsehES0f75LK3F3NP99zjT/jAp6/RrXS7D/vfYWehE0GUgGAUqr9cQQVeXoq
eAkDibG8brYxmL3yeWNVJClDUoe4Qr6k7mACTHgAzsh4WQohLSr37EQm4W33
cUcZET/Wa424LimtE+Qw5/dSC6B6mDGitfB8JhExu+HbN7/Gcx/rl6TqcOSO
8tUHMSZ9Hgf4L6imRH/P3cQJJlqCixp0dgO/zHZqti/38uzGDKvVfbB28TV7
j95EUH0nETTLWuJ3c8x/uxu65MFXthBY2Ny+oE24xRkHweKVMwcTI7FpY/vb
DKFYJ+kDn95+EAcaJFgxBT8z8E0Mhs4ZNmuBHXBknW79DbWKxioWdgaJZzJM
usOjT1tUrVr3srI7lbRk0RJ9dmmMLhQdIOAPlGfFNsJ/XVSM3/6UQofdt1iy
yHZqOMIvLSqUtXL/JLaPplacOo7nH/p13MKzb3N7Bd8zXuwk2aEBH/Zw7rJ+
J9JMj9k8G7K+qhbLUKt/82rFpEnEB5ujid33r4wWd+mYHLp59aJCUDywGi5S
2+PpF9fEaqb6EKQ0Y4hMrKZmm+i8izkihWlbY6AJon9EvNLEHPCD0jZ9QghL
TBLnpsElhLqm9OvYveX5sEhxXRYU+AI9Ey9JZnatYDoz/6H/uwCnD1DPDs+q
nmj1C/wUZtgLHFrwnVF4cmHo8B7+P/jeiXDlzlnQ58yKVFg+CYPd0FtXf0sf
cNBD+hMQ2w43HrUpLtPF75CYGY7SGTPP1ZNmDcNJw2lNsiePn5C1exS8C+dZ
NqVOxtiPQ9inejQXlVqN6kpEtPsUBn/pmEUYUOGOB/Fx7E403XzdCZgEwleQ
+Nz/FGw14R5bIri5qdmX91aKLzVvO5vwPo234oVM0IYBBTPpn4Bsy25kOE7d
MjByJzykICZEYzdCvOpcWpVBSbnQyNieXc8uIWmPKKXNsD6jdFfdAVHUeB4O
An3SIQoUb61q1sDkLSgbHYHs+nIqjGHGdJU2MSlwzQHkJwnL0SQmSiZnOu1Z
7LXDk31A3JyAmDXwJEuD/5QhLlRWWgZpQNDfaymTZYFEqvJATMatLxS21Oiu
siapqM03J4apc++Kf6xHuKWteG1gWUK2GHcy0hZcFLZZsh8aqJbX8ZWF6KMW
9RgzZ2nR/IKpEKint4pKfYA5jzYZqoBsXMXUX4igzA9+xSDpTqrF1KDf2akV
+hfLaVzCEMXWBwRczyZ6r/9hJkkPHgNA5eSxS1wY27cLruqhJorVjJDNan3I
GJnDPMsWotv31yCUGYw5Rwk49OCw6fy3dAbrrXW61xweHRs+TSSGTaTciqc1
5uKSquwwTA8YU+Qj7no8XTFKU43KaTnLnyTA/T4nqvp9nnbY2hjKjVCKNXje
sToMRljZXmPXAkxGO8kkRffmWJB6/mGplbYldQuyBKeTfHVowttDUMEGsxvh
lQSGdb+q1ers1ndCeEuX+saE+CkXMUhJPEBISBw5vKDWiej1G8i1rgoBzIS+
oW6I2ApLC+z1no7nurzxXx6ITNnav+9erjOpvL7xXIYKvsYYl3lA1UZmSHJz
DznxM49rMd7LOtVPmEFlFo73S9Y05c92QJCMi7QreVWYcLqTro6ECWnRhXA8
DvnEhDF3XAgscVZHcW5l2Zaeh4+U51d4hUwAih9hW8ouS9hS1BjW+YRyiXx8
3wxwfgZAInnjF31ErgogyT7rb8i4332Y+oezs6sdvMDDlk3B6Qe5ypULP9FX
mb2ZX18JuBSTy/AixptKdqfnmTtFdsPP517cKIRWfidy8hGEhQZkpv3A7cHM
e60C+aJA3Kilh03/Mg31/JvGoLTlJrR64DMFxt22hxHhTJDAhK6uv+C95jtq
f19UchvdxDyX0TvZ5Xhn1fRAqP1v1rXBrIKWcXzdHWqprbK1l1+Ij5IkMhDL
pOgNRw/QirW9fIxbOCoIY8HWGjMpK+i5v5UOwuV01Oex23b9EsXMDxVWECmo
3Rt6m6Odmy0YKN30V+WfJDxPGR9ZAJcdDvy00ZFD/HP3/d0zBKcKtnc6lnUs
LkqkQcEBk7cYNpCRYpIxM7D50vU/8OQOfHohNNPHxi+rDfB3fe27uyAKpt91
bgE7psPfSsONB8i5zUJKaymHAlZAJyflspHtmsMOFxTGAdi2tOsERavtLqK5
TAP8SDNrLTS9r3z5VaBoQdIjx/POr28BSFnECr9tROXrQB6t9mkyy5wY6uRR
w79bfQkFTT53LP48ITmnja/NsSEWaY919/SgKCAmX0Kte+9PVycYLbn18laH
R+gwIXymGTTbxir7muJ5bqzLkA8kJ7TwhbeTjR3gyaRgb3gU6HeeXy37iOzV
eKNtG3gKUPOoFoeOkgU+AHWCCSX33PKHB2hcVBwCZT1i8FL/weIoow+JQGsU
Smup1fiKJSwOkGy+tvAa/RBHw3YPtKvP9/cs6HFymHTT4S2JNPLVg+RUKa62
XA/xblZPRri5BufBk33WEhOFY6k23In0urrDUWDjX+IMXQX7dEXKMxmLJ7ad
kX8LlDiLaFt3rcTd67zAp4W3Wd6BbYOZcfydijGhgPy2RT/B5R18JDMAJZqP
/QSGsRbHLTyYvJqrTgY0KuMvns7smMfnF0IbGr7kCthTErFLHE0VsNm+WXqj
YiJHnNSWSLT15Scdpo5VQeCNUE5RL8OvquV/P2rFIX88XSsuVVhanCM6O2m3
F6taFFPZ422V/2rU3x6de2dvg/smIKHIJaFZLhz429jer9j2gkbSFo0tDVI1
I4UfCV75WG911aWiDIibeJoFoo7yEChmhXqhWiq5WTGdejvlOrOty0n3PobP
TYqFHoeP7PgskCSBR9tGWHPCq/LfPIXKKRrEZ/KHa6u6sBqJD2X29mCwQKNs
FZ86jUIvGJjvqfQSGzFCIVjX6XsgTGSn0VDY6wROA/l9LXuvW3BJm1ywJ/qL
hhEAaRebfxhZCbSuPonIUh3kx0cVxIyeTLZ1m4Jdzfe45qTJSQ/JSkGNBpN4
MGnikgLko7hdBVxJI8kScbO5cmd4TabV8ajUhy6IFGmORd8lVAK84sURBd1n
6FjAKhPBytfbIJvQfcqUwZXleP0Nlo/HEYaO23f+pgc1dKXI4ZWZJteA1Kzz
oaR75rrvbhMn2gTvtqpv9lCPbRYUCbj4MrURzkUbGEHyQ8vAUoVPpHC2uybQ
W3RTs3eZCFHC0RoSA/CSWsthH99QknCRqKtd8tYEiB4SWJWWsRVBq1DzHjkk
0jgEg6B6VLOeBBAk84lt9u3ApmL4PLGWGtJJ5SdEdpcqb78Klt4YkpaazX8S
2m/eolXF1/LddE6CUX7tN/ehRCDHydyLtcVAVRBImW81xRygGjPYEnJKGQTb
U0cwiFa0wGOCoktZZIvTI7J/Bz/32VPDiR8fxPca+mrfxPtshXLVXo3Dqamr
RFdAsJjORIcumkXSaSGR8MPhcw2UgQV36+K/2NaKvKiKnpT57n0DwKfdGbaP
DshCGsC3usXZZPX70MbjVVREVttbdsK0potXA/NGneYabBVfFWtx8VneL2BC
GTnNOQ+3vHJcYoJf1DzHOdKaBVtOSqIGvVzWbeqwgT1FcGCDa2QKSmJdfPZv
1NHzZ9XFIVXhCaC21jZb9OC379HY0KFSAN77Hs6HMOP5X24Vw8XqjSl1wd1x
NDubm1j+xQfX9GrjfpT2Vv2HS/R1ROP4qKobVGjeAWzxWrSHk11LNdrNIF4C
jTlouFrA2yNd3YlLL6loCh+dberIy+B2+uQRPMnGNrmW6Fh3WGronpLjphR+
8J5CIOHJDhKP/kMmBoDm5iLMJWHoWImCL7R27GGSIkoxibnioNriRe8F1PJ+
/d+0mZXzmPPJZzoC6QrLadYgUeX26VkGdL3dd86KPt/W8M0ShapoHMEImOOv
x5NxeVMJp8MLwTX9jV12Z5NfClY0KZQ6//t4o0/r2ZkDfOoanYFng1sNLy+h
K6I9+Ptw/ljuPbPzCO+aQdVXh2Goc6KQRkkzjXgoeIb+6hdmNqu4L91ILM2V
qJj6Mw/FDQ+dzJ58w9VbAOO4gCMCUNgf3EkcNE+XTThHWY28XJhowhewJdZq
xt/yy7O8UyxEmSCyQwhg0hZG3E+n3QCEtt42cF2BM1VzQzbgj5tdGPaKKEBY
YN45s/yjNfLPPuqFpSGT2t4GOmcxzRLIv+pFqahPPgVLBfxMPZAHsnZqwQHQ
k32gC+hGW0GNAlmOvJdvx80gAmFsolnhyxPJ2PJpfvsRiu3DqzOLaGaYoG8J
+r/tHZRl+XsESsmt8AkdMb8xsGsyKC35JWZzWw+DEzkDypkvL/4x+o0Brfan
9VXrFcyVGNLs0brP9D28g/7v8bU/jx9qhRdZykP9Vkh3WCKWC9k0ocGPYQkk
hz+yrvjLuP1akK+lUFTc01lXUfsxq9eOAxyrleBTs+s7qP/+jAP58NQ3TGYa
sT0RZKSvOfKfJWyiH99QaIp4Z2WNVrgwwQsYRsDGlpuehHV2nCiQM5APKlnH
HXs1Y3KE0PHR+3ggFlt7rtU3qk0pcqZZ8Pjo6bNKxK+/JfeZPE5EDmCuYdWT
xkuWE4ohlNcLpE39fYzhV3s7fmXlBpS3Q62sTcaKEkBTBAIXXq0prD2xeMk/
p13RBDjU/iE86bGDBxuWQWdJiKDsbI7cFPXpVrqCelpVGm4WIlBxpqySHKNL
8LDQH5bc/iyrEFlbVKfFRHjZHPOj7dseq3oehGs0hTgUhLrEZa2EpB+AB33R
QXafFSgDCumbouocZZZ1vSShFTMhaA5TQk1TuMQPVXavzJj+TEU3XUHRh2nZ
P+G2jrhXZ1lvSf/e/Oz7QmDg26KIaAkcINQvMlGxg7zD6IN/2WG9znY52y1t
qYpEzwoMf1/gO5sVIVJ+Jt72K91vB88h7YMWoT//FxeL3jKdnkKMms+WIcCz
IiidAjP9qXJOfL1MRi8hq2mfHrcX03x0TZV1DMrz8ULfcMG7EDhJhNnzno4w
3x/SOIhVpcSPZvUf6mzW3nMmqFt3zpm+nVDiLMnKnd7gvs0zu+dX3B7a2C8w
kJGfpAyPCu3FUP0pJy2jAmFPeLHzpgsdcjEAAtlbBBDoddwDJQCIIlZfQotq
P1agyMbeUrI24lAvA26BCeF+oC7dz2x11hEflFN4dceCSglgJAVGigx1qYEG
bzz+jLlqzx5GruXsQOGBAKnbTp82+BfcTMfIMTTR30u7lo7vFFLKpTyaiNSr
BS7bT/slgcnQv8bBOmUV5vOPLT1hrwmirbZJ9eQGYSMAdpXaC6HsWaKtuxfw
eBnL+JbNYuPYW0ec9eR5ke14FnXdymGofxiRJzkymKMIMKPn2n0zcJCmLCaQ
oRcXkRTma0FYE/Tz5y9Z64BwzTpiVqmk2Orw1RpoToTRShNFP9DNTwsDRhQj
cdK8jVFIVTFdUPsdEGSY+kg00CUOzHGgzoPqCJH91xZO6zJ9tzk17XCXMfh8
IX0wfG2tmybV0tGqC5NlBz0SBth/PNG8nhAiYN1W8mE9HuCCsAAR3CaIurUM
kfJfLr4PvIbXpufJ2KvJyoaJ0RK81pQQ5RGJ50QrKribX+pqfLQiYJ5/oRve
oxTtk8Rb+LqN8VlNlqEmgnf/ojRj+S0BU7JAbYlxeuKbW3tLRa+WtR6QcDHu
QDEPNXRM5O45u33ukHOw3SlxCrCF83nynwD4Zt/ItkHouKzQfypystvO/dpp
VMME1RZ2HZpOpbbjP0k12zzUbvY4zZ/NWVQp11zPbfr8OHdm2C+sezqxSXKF
G0l16PiDQLcL6+gs53nNeGvRD2ILzFp2MtqQV1Ph05kVlnJqnIIZ6QMnVVqZ
lKm7xBlJSTEftnNBqAMpif96idq+2C/hNlPnItfAbs77XhwVj74B0EMXufde
NjjQydzy5bxEg9zwoFqb5HrId1A5xpmhuiKIuycSrNYF5P4tzuzYejSy2EsE
sNBzp2t1JxRwxyzakxnyqmWYTRK2sOkf0+Jo0HKLaWvRPAPA0R53F/gm47XH
lRxfqrAbxe4IkZghT43adZBdU1tMrbWS0tz+27s+n6suQWr79cWHfBWnWbXP
JTBhygLk9Cv1hjAN3+IWIhKpCibzBIsLkZoFXO79VWVl3L88pU85Uf8eoprP
Wf6PeVGMOsojzX/5aVe7025HhFqxRJsZtreXefe3Nb+f4rIEMcdAuUoaWyar
RuNoqEZLjZg7ihwyb6VVziT322sWbfGgh27PoaGCj9Nqd1PjpV2k0VPaiVAo
j1IxiwH5BOtIWP7D1NYzH7BAZqRjG+tYb+wREpRXvYIU5Y8pxdNLmmoTS+nP
BGZn3rcKX7vLaS4BPBo36NBEZHqQYeAFaj7rOxEtJBKLgZgNhOrU14u/5jwe
Jgt7m5D0V6DWBAM3KaJYVKECzyZicGUe03NvPJStQqiizZQC9hsjPCwjTEL4
Dmk65xs1wvtbKzs1TcOZpeWP96E+RvQyt4rTdbDydkjTBxpglbsrinaG9mbB
hdRPCDAVCwdNEH0gXTSmDenTZFSDt0FMknEcbSm+9UNEUhnPOwhtF1CcAwow
U7gyS5AruaAYpKT9NLQ5pgVDwCFCcY0cKHgsTUZ6QIb8jemluw+/kw/8FQG3
Wzt4vNXsX92zLKzggCsup0rIMIBHJLSw3/QI9mHV1oZNk4DFZQk3BPxwPIi8
LaJzNouUMAIvKPjLZz9zx66RSuxauBcLC68e7vsrvhfPzWS+hEz9OUSUBIaM
ABbXgNfX9RCr1UbxMV2o648AJR+tQe+W086+XVpxZPtyvP+0fZ5eEqDEasZD
Qs4qBhCWE4JVG2AF4cYpisujiIh+DBpz/+gvLshHUTES7N6F/OXI+wyUrVK8
AS78eDObBdPyHhpXZT8nKzMyYf93mryStnSXOnBvGXsK8flZthhAN3TxpOd7
OM+U/Lc+yn+VU2W7PWEIMnDBUEyZitFQjBnT4oXi9lTWLjlj1KBb3gpo3+oa
OBVkXOYmUhGEx/pocM8p46gETSeU/3U7TmbTh3dKk9kYdz2xAzk5rHUglui1
75VciU6LyHgmn52DJhCdfB4hJF9kNul3FGPR0XLgMCYajoSydA2iGfq4fcwd
xPMOe6vcivj+Dxn1tVlpsnwqgKAy8Ykc345w/f14jfFzo2L8aQRHjdPR9C76
ZA3WyCrMNuJqISK9tsiIOTYXTIXB4YO1eHSFON+HzZFSRoPfhcyvELVQkYSF
18RDA1dnIDKDhgT8dZwx3hEpYhtSkbcIjcF+vP9lIF96ZI87w3Bx4AnP/f3t
X/c51LUSJCltzUSHVIaWnHQ9yjFK0Jc7yYIxVEQm3TJz9YF84RCorY+1X9LT
MQM6wT2GY5eD5MJEqHUV2G01Q/VegltmdVS+p5NTUWAjhpf7MFf6Zk5wDk1K
3yEIKosTDF+50oJhDaZjS+0FlRXPFJOtpvCCTmdG74zDq1R8vGx7HfJEXd5I
u0wFue1ldrHQ72chuDozOYxWOV3FK5ik3zzq1w8p6NegVJ7x8e+RLczPpJ8B
2ZschAlgUKn1J2LCYy1Lug8KWYrbYD2Xb+EDVmD6KLAU4/PoNTUlpz5f+kfC
JgnuRuslKiwDxGuqJy+wxC40y6MSb9VICajC74LkjrelPk7JO51VpEmx1NmE
3jS9O2RwxeffPU30wg59usVdY18LUyubw0rbOBNtRijTtcmjJNh+nL1CE740
0ubATuihOQvMbsdSy2f9jdmnZM5lp+qlgdsT2IqAS0O44ytuL2qqvTSiG+hO
sQtIV6zvuzN4qxXiyAbPEkcQPeB6jaGufDkhc5lDb7o9C5Kh2w5ZI8Wx1u0j
ViWbB/gWzXSn+Xi2PPYsUPnxjxdpBtX2l/TLeRRRDAPZdmE8jmnvD7yeR0j8
WCz3bAbNPbWPY5bjB1jS4DJvnheAUrKyXX3cm4D5eamTchrqF0GLC6uHtTwy
oNNmVzFOPvXrIJmxE4O94/EoXhjLaS0yVdDa5QXRxywwXHkN8bsiMiRe1LWK
wvDe5RbfXNiXDLEveiKS5B24aiG6krIJEJs60DsfktebfUL+rNZonfn4DeOw
1j79eT2vwM64apoE2h/S6LsB3a0NCXAO8PJR8hF9Gj0Ts0ik3tmwltBxNeYL
VxFN5g+TdmaUlWsIxsLv5FuwLkzaZR8TTrv4IBNTJNawPw4ZoxA+/82cqhLY
WUGxo883eLuksZHGRLeEeMXMyWCXbWvqogwSkVNvUA8LZ4ae1rJhchKXbIJ9
oweUkvMTLZlpuBGjl+M000WWUefuozJZsr5pH+FkyiCf/6nFu1yZdy5ycHp2
6TTr0D+rVDKNfvMWoFLYkNqSNdxTsqJhW5KY73Fm8DSN0i7tr3iSP2c4c969
YBBHlMOWUhcqUB+kccRGxfC6NcqRG7tzy75OCV1r/ahw07EI6/1exEqAmOax
EI9yxefv806i6NwOZk/aNOT8jJP/Dn6pE5aM+d8QhKrXf2goLmcPKFH1795J
dzMdCdG2SczmQfSuGgTPJaiPrLVEc8PzJcbiO0RAegnto08a/Uon7KwRi03Z
xZqBg2o9Sk5bR+FXxmnJIV4uVX3TLtHgK/Dl6PvLyJu2gyZ8kw31AV8Akso+
i6H8r7xIwdaeqLe7n7pdESdvViJzWuPSwxdXDHptqa9/JYCk5xPKFTo29zip
rB5Lw3V1ozcbxFctyjjr1Amzw+gQZyRs/H2Wh4DEuSsOpHXVa00GlLe89hq/
15ec5BJn1gsAxElrCm5QW8WgWWsUdRb6kFiwk0C9So7wyz9gSe+93vo3tFvZ
o3dMS5KYnLbxnumWc6gCmncbvMcGN20bjZ3sWrlSD1OL+6YyKfXSjHfa/GxE
vDgrbemfVHAzvLuM7iF6G3axySX4396FN/rlEX3W50EeWPP89D8R8tkQFa2+
eS6tmqqaH+OalOwnieccphHTuAJG7KhnWI+7hb2UZN9QmKF9hgUk3CNwJ80b
9wExtleWoURkqPKddk7AVLo3+SNYxR02VteTipojcezh683VfWJqIgHXF30n
kiLPK0dh73B4aXFNFhJNt0ByFb2bfR81LuHQL5a5jG+SKuNyQZ8zW4LlGhbY
ekmRDS1J3UcEYpVYK9WoEgMQJ+y7VdHgVq0GNlZXfd3nslFtp/2CEANT+tbd
NCBlgE0bgEH6QV5r+LQYGojcVPLLzqgJWRKACEz5xP9Y2wIetTWjfENX4CpS
iT3QGD20qvdV+njOVp7kikb43fDKKAe+Mk4uYyCvzu7QiaNd934VLvnCE6wi
U8k/6oZyoo1CdL/jUlKfcDpC47Ij6wWTWuz3soe5jt6l8gxQIV92S9Y8P9l/
ZmdIiGrCkRFiNqTzdgRNdXyrWHPCBRltPk60lJQ07JN+6pGrezOJeESmAV4p
M9ts2iq3g3hJmXNuvOhmtqUUEu1cJ7ansEb7eg4kG2UA0zokkgNmIdoNuzzc
oJ/2PWfi1R28Hr9q96ALMMxQ7e+Bp4w8WLxNTQFMNcflpiM1KOwQ4kwW7fp8
qn7P1b1yj2rO3opaNBnEN+gaXUBmTzEZwrsrUML+Tz2FGDNuUABEdGgLgYu9
k74QQ0F3VYqAoboYw2/4nsr0n6bsi/AMa8eFTALUSC8mH/hhTvYkCLPOTl7D
3okG10F0WGQakjmHHf8CKboru9gzrrCMNIHmhUNYg2lhObDmxM8Fgk6SlDgZ
YtzaD89bkRPsi3yAiv6z4rPkrwVhujvGtKTRIhUeVtzRxK2RKjbpz/4Yf0Om
8QKwNkdeCWZkq27a6fLG8r6EDdBLl2YGEVQHxPjqI3Dt+6Sga85kveoA/ct0
wRxKY/M9+L5oRsiTmDIiiat5wtU4/B+SFvJA0RjgdqNh4Hd7ymuS4AlaDykp
7+GJWieYa/Qg2097Hm4WlI93AZF82t0VYguKPr8InmOzwbZrYebir0j5gWtD
m1uF1BQH0a4v6Vy2QHjg09Pcji3SXYcK+y/TJTwjj+MwfDoXA4ObdlOgV7fd
/KaJE7U3e8aVNv2olt7dFFcd6QQB1LFEqKngzee1oeQ9bcMZFaAzVeqr6ooX
hor1dYNV46jUPNDc6olyifUz0jidvmL8D5RIYArxoSsv2KmWkqMsbqVJyZqO
zbfRxyG2v2cCZoSG5rqrSB7CH55omX1NEF3iJkfdo0bQR8o5jtb6h3o7BjS+
mzkYBQkbR4wuvh5MlxEjuxzFnzWA915vc6cdnHarpgkqo+ETqllshVh7+aba
E6ipRUdsLwlPGypbl2Y9eNn2SgBZTPwDGJI6gpw5jPcbVNT+ZGN0TDK5uecb
DaYm0WDxBds/ttuIXM64/j3SL/6xBR23gKO2zfdB4SCyw9RLVtX+YzKE+vDw
NXUnmWOcB40qMuS/1pMYbGFjimwdw5TroNMm/FjPOh9qwMeudOjolbkqP5bE
+Qa1KqWO2nZ1dJjgzj8Q0gTUyDlRfKeC57MkIoDVhuhs35uwVZaV4BWepPjH
AyQTPUOLILZ+oJ77B57chm3jJRueMdFcp6Gw8DzOVzNaI724AazfYMe63e6i
BpoRVtH5uu42X8ApS11vjabaXpffdH0jSQlUGZ0hkegMAgwj3tLLy9SiIEzP
mUP8HL1zp3WwSYOC/kLcm6kkekUcHNCnh6WP13ulDadigneI8TWrrcBzACo6
BVyVKj93jSJwA/APJp+zCzg3+IOII6B+e4Zo1QoFLu2Tm11uNXoMEQhGVoYr
sQ/AkH2G4u9OK+Q2C2QC4bEqrXna5xdACA8qzEQOB2wttNMAE1esBFeEX55r
YrlGZVnvoqRJOX+UYuq6liiEfTf/SmLamGNOh1Bp6kximJbkC8RIy+csoLxK
J8JUuqF0bRKEKsyoyNlWAshg1/bcuuHjXPj3BJIXENt0Yob7oFiqo2dDZ4NJ
UkBbZ1RAC6lBUkt02+Mj3lcRuXYtzUyxMvSsQckEYu4Bw5wkgPS7V6gd/nA5
S6HDNSygcBTGzY1DxTDuusJAWOgau1MbJh0PbYyQW3WyI7dSUSjZHHDeKliM
jAi4NPH8wPMs9Pjagjc6Zis6E1N93Y/BGtxyBPsosVbishgQq7SGhM25c2Gj
j2ZzJKJe4/SJKTtowTaHbufYwHGW9B+WsJKhhbV9W6wmA8Irp3fiES2vvQCA
gRqrrWUtxbftawZxLV78YORviORrfskC00jTik5gg+TaDn739SpCZKKhfMlS
hur6G7Quf6bCWCDRUgmzLyL2yTUeGUwom1eUtMz4HTT6Gh1AEddQ12zjePzl
mB4qtGQM9PPTSI8FSEAszP9a5tHKmk0WXOAxfjV7aTzkPChQjpwwK8VLO5uM
qLnlAQ4Yj8Tvv18mMS3juNJC6PXZL7A8cnUYY1sniN0W9IxyXEaiJf7syKoM
MqfNft1Bi6uTknm5jQiQCc/FKzIzcpGIaRAbwzehe8t9HVUfzKiJJcIrA5Kt
qHkDYzfK9KRcUoCyeNZ/UtJskjYt5bu8JGqMJUAmMveCZ8vyorD4m8KHurmw
aunHyc7MyUhgjo7NO2yMelkwxMOItr/psaALUchFgHZzb+NXCvU9IiJH9gHn
puDCTT/G3zk4qT84fQ9lzaBcmVMHkv1tI5w+ojqluWLr4AgZ369ZeyzvmO20
AiqLkeYi6cATTj6k2ElRB8PdbMxuKqSvb4LSYb31siqp5oCaHuHw8XVnXy5/
+r87Aqjm1yr3g+QTeLFmoVdBNTkBY+fpvyJone7LxDlPN2ZF9d0zdmw8c0Be
rgSiuaSSsTDngQEKyi6rBk89SC1Kb8TD5ZhsiBrAv5UNHTxIuNr6VFnkUYvh
3Kywt9U7DvzUXBJGHc5z1mJpwfcd5mrmQwLknVLQ/qlUdPRJWavb5S83dHSy
bX10rzCEXXiLWAKFcIx4wfCWURhuu3getnvjlEfHF0zY3OER8JUwHm1LJRC2
dZF4jyx1nXRMOwtQSImnG66dbPlMJmaY9/Lwq2yPsocGlyRS3DOgaf+wVvMc
TLG7lqlsLkqZ0Nqpo2RTxUbePY9vZsBbAPdNfsiySMi00XVKHj5ThtVZGyDC
9Bd2i73h/FstQtL/dqSd0eLgLFmn+dTp2JPjv/BYQNuBKNJo29Ks9jB+So2Y
wiF2XYUJl6rVKFccl5cdxk6Az8ljwO8nQCm6JXMALOTOq2TEFrDlMLBydaKF
UwkmTspyYXaYWQTyU1lWACYD8mcqETaGqT/NpAlnD6rEt1OmevviEnOhQKom
VB3PBRYx38NmHWoZykLQdtN5sZ40DW7p737RtUGNz7UNS7D4WiY8+6aa27NC
l364Qmkub6znjXlt1tx/yCFiDUxkshnhVE7LF9XjLSLZlJTfoWnPrpgo5Deh
5oRb8P8j0H99Ae9AbTtEAbzuCCLvzvx8sj3Gbt2ZFQ7GnMVGPuSrSv5y+OBB
MIFTeLcFJtIOJjGiJSADAeq9mH/oHtN+ngu/WIZ3tWcK6Kq/xFkXqD7NGx+W
NoGXTl1e17lKXAulxpafny7242Of+n0NhPLihtOIZRRbV7X5KTn9ArGpRNL6
dQm7wIYJisqUWIO25j8X4UghF+XylVb8hii7K5zqx/R31jDjl9rpAmdF5g4W
hzvRwhfk8L8Kx3PvoBlPqQvEu13cy9+bUAlP3CuBHYcLbFo4Ss6JDQ1tXWdL
/2Mh5pREn/nATOBkMrtxKMc9hRqQMJyfvlIOvGYKEFaUgZUA9HapzUWEqkbT
zmlNMoWnHQjeyBDG0IW/16vYBKiHMFoOlL29CjpIsJ7H+9kVVlYCCEmzqMxV
LaGuuAivFqemNa0lVazIT64tW1MxsVJN8z0t1FKCtSZBywnXcuRgiwuCxRZ4
5oG3cAk13YDjgM9fvTfCFiH2OpYQPgCu6q95glKTEEYNdq1TGeuciF0rCrh1
HT15OKD0HoGLW/Wd9ATB1j9lY6v2NQ1PKu5kanF1M4KCopRCJHQEiNt6CESW
zBcsM5SQsRutLZp7dziIe9SoyYJgxE2jkQOFYTjwGd3GPT13VbwaJUx8tfjp
3pwXrKMrClDn7mKvOVqBWcIOr9q+jmBG8zdeIKW18bCTFl2PIq70jl9aRa7s
5zmdGWwwZyftL8l9VoiVXhcjgeBCOGj0MjDjLmIQYLZuHuWOwAoYhHvCvNdl
dhPuAvkz80bjvGDbG70vUhAGyonP7GVkeWjWJ4hUUgTe9ocZyR8e3OlA4r7Z
ZVMGtszSp92Do93aJAdwK+jQ/fsvWqBL8V080tQ2SIgU7qa5yEiDO9Qwf9V9
XzsVUCUH8BD4z24EecUSC+Ew9mY0jHiNhB6jl8ev54XMW7oa+AoRi7PW1gix
8xzYJnG+2Vog79TPWgx9BPC7opP1mnEsxIm6uu6VmZRL+bXjZ5LDZ9uvSVta
soTvX22dbFMMSquXveDsRRCf+JYdDnybW41lt4lGO+gQSB1BLWGDL8znVYL0
/S4ZAhzMUuR4JrXrTfqgKNgkbAFPBQuVbhncdjB546RDNTW151+AyXTgsGAJ
MwIDELlYX3AMUKuu3MeAFNYjGPG4G4knm2PzTgUXfpANU/EOXF3CCposdpIC
a5KeM+Yb84dNbndoNCgjldWOrQ4yc342qCqGM/2JgVbgw8HT6Ozga+9Ji/4u
puKTDZctVGFHwHP7qtQGITLLsfMdUmwNV+E+8mb2kd8BkSTyehzMkXhwCTTX
8PXtWwcuj59JXBo9BzqC7sfGT9T0aWodw6Hm/1bfVKWKGh+eXUMK6Vldpfvb
Sb/RZyiaTE3OT/PWJzinKi7fD4sMkMZ1VqwmtJ/wUjX/kiDzvrCoc0py5keB
bvBjEUkDYIwp/NLwQJLFqUsycK8xxEZrMovTYTHVkvLUNTBV/38Fiek6t06e
C2loTBFhbyM5eAaHKMdU/U6dxTDTOTa6gjW+gs+1bbgNsNqUa3gq2tBhiGhQ
P0A2rtsSM6lx6SvCWJsQJoDtzDNjnMXwxVBzXLtg4y0JJfn56251qa63yNmJ
njKm6Ka1caswiWNRxZbY1D5trQQ+W0PyqXDn6YY02ALMFIzh1M0T2aSOnV5i
DPvs7362DpwWEDh7b/FHsFLCNGZHqTd/Jw2EIHu6eI7V7owEpj4NhhdkW+ew
0gLmscSqFqewfYvvETMvvrek8afwcIZNrhyrtBzvVz9nyPBuHo8NUot+fkqy
4IgyexJboq98xOiqRsMjwBsng6kKoQMTZsI3OKOVLYDhEJ4/hmQWohS18XjI
6H6dJtEHhbMn0AzjnSBS9TsR2dgaRWKV+6zG8p3WxAegrF3BUBF2QdfC/DiG
Lx1WByK0yymREBaVNy9+OYq8kqE62JQUin8RfsNAAwmHxtfssB6U9QP6SGtf
LdGAH9fdMu8liKKcZmWTGtdkp6YR+5VHFeu5c49d6B4wZSkHttmI2uWLayIb
RwP6BgrRIWTrxiiHwlrKaDbj87WJGpN7pV+Zh7lOc40sI0BHcWArmjBvKLZ1
42aWzgMmfuh5ToWJfkoqvuDMmMzlmuKk7MTixSkFfRzwXbePqDbg9iN7Gtko
Us6DPJivvu0P945/jEq5k6UMeJy+eaekQsCBxx5VxYdQzYcj5NNZyhWFWI1l
wNU58xeGOjtpRsedrJVZfpglPr2bWoOetcTCwOYBYX/uWdx/h0Hb2wZbNirq
svjMS5YSOSRkilV7gxlbJrMxAymSByKuTmuALEIoNJHnkfyisnUWWmQBaFW4
47jkUyze74v8S6s5xINigOYpkxGuNN6X5yQwRCmIjnfoBAY+ksAtS2ht2ntR
jtlxcjZucv/ZfWYb0JH0w2OItHeyqv0vXeB6jyVt0xwafepdjX9iQvEx0h72
3cIkJg50457wxS8FuX6KriCBpp0LpYkD8jAIs3REBRltGHgNsmE5SmOOpceM
p9Ixtf7saW0TnYY/jifeoMujoGYT+Pm3iN3xsCIb/n3DgtNXKh4HV/fbKVtu
jkIdl9gd8nQq6axtB1IqbsX7OSInK49GpesxZl1IGVdAcFUULYrS6QhEZMxV
RWubhxQ9xX6xWURs1gwsZZsLcXqOfN0vggIrYKZCpcHBSF1qjnX6uB42jgjF
WBSOuj0U1Ud5vdbfwJK70p9Hz/R//Q1+OYUx0kfQLBnWATMdykwWtdh7Jp+H
dLLjO6b81JqDMjede2bC5R1KCTK2IV2OBB7Xj+LwQHQVkeOfyO5SH46qJHkZ
E1kQlzTSEq5s6dHeouiaMDOfCUT5/A/QmyeR85nBMbCER12PZq1A+hmCgLxr
LQglEhOg+AkOgBowcIfdXZiYzsuiWqkZBBVi/Q48wa4u4hGtUbdiw9Ab4TLA
oPMjGlfBlDRbCM2A2zKVnMAMUOAA5xZbj1BXlJ+C8DRPDR1s5TNcP15HhLDp
VBeno496VnalwUkEG1AEywbpQsNtvtO3D1/R5JB8b6QD6q9NqZ4dB4pWY7wV
EjpHdwXjyD+ifuQRKVZBzQxHAYWdRO1oLW3zOivoTYbwuBfuilPFgSR12Dch
sttuhhkOsvzOpmr3fA7cVD7+N/XgROzd0exCD0syh9cQBz6SteuHZsxdrnQ2
RJ5oEpMqP1deNDvtVP51OOnTbRRHHqsSszhQsuCxLMY1DhNI2H+MBwWIQLPY
if5VCiY8Zde7nAwqQ9/RA7wTe7YXO9PdO9ok+s1+cFQo4E+/E0gV9GBcAjQs
pe2RG4MGNaAG3VDRWyPixfvsqS7hn9uoc6cfZE61Nb9onXgv0h2+6cLnEbmj
yWLUD9MzgDOBx4S7kyz17g4f/Zd2+X9KIC3n8/gzVLd4/usbyFxMmseaKqO0
h2QiN4GDua3Ax+JUNzJpl4IpwWGDYT8cpIiTQK1y8DucJaYL+awRs/eHpB8L
XJJadwzNl8IrmNsQAW84X4oUGB9rJMpO/6USikljUDsx1OWXQiviU0sea2v4
D6ZY4l4UNkKnoogmQZe5hSv3sG7R6eIn6oWR0GUly/8zXahO5b8xp9ADPRwN
U3Imjx3UYP11NKiqZzRWhv9P+ta1w5TKEPWY/OHffevgw8c7tncPTqGV1d4e
g058D0gw41Wff2+BEkiSdk9vDAQ0L3pOrx3V1socA+DU+IJCEaXIoSYwTlU7
4k3ZUn++DIyhsZbXYhfKHqeA3dxrji6dGmCqEAd0MIBFFWjzUo0mxt1FgxSA
tx3imTcNllKUvTD+/Tpo1s+MZ7WeFLlJKQu8apYdbOzBO4iRCZW7BnTFQysB
6YGsawXfOz1+VzaTmItCzjHNLJoS9mnZG8ZJFcOZL8iT0IFVsHlsozkgCLX3
6FlEsdmP/LPwMkKTSGDzlBYsGdduqDdWDGDMd/M1OuNnSm0aqN+xb6T9BElb
c70TjZWp7wlI4CaxCYmws7rI4PBZm2sWErWWUJBTcjQZ6e5uQqI8lV5qV5LI
1wedS6+c7c6ESDOyYfIphuirlP0I6JzE/fDofLDHy2yZjdLPuA9MenIj5fsA
CIBomijAFQY/+gafpBduKKERxKuLHdAdqqRuYoJk4w0cJkjt+PPn3Vb2d8nu
eDvRMB/6XWfa2o5mXn16tAgngY7LaMes/uGjUs6eP5HLmFsijFDx9FUIsleU
X+AChisOEvU7ELlFFF2zukhML2Di3DhTxwlPbgKTF3L77YaAFbJwnJz/eduu
FqzeKyec6yV5uSg0HfByl7ow4hJTIwueMAxaC9aArTmR0PnjI3Ry1XN6blay
ziL805x4TsXetZvcO/InOnkZ2zqemUqfUHVvfyg8N0KJGzuTAvCh3XNfr7Fk
LZnyIkhBHEA7wNwLhp0emFVCHyq5SuUBzW3DN1/i2e75o5+CjK7jsfnYAMEF
LaCl2ZeUjFznpGktbruA47NQFevB2KxqitKDeb2QLktPmZdDD1gzdgkXpB0r
xCVXS0gP+RGyK9GN72HO7BeCbSj9Wl667Zj5ELJqG/2qtUCII+sZn+Vj3887
/m3ImGk2po+FJcmZyE3+V8RIU6TX6cz7i4rhkjepdc6EyEhkv7ZbDysK+IWG
XhDwKVrY4Rvvpf/ObVKKiv95EeiWUCa5s9xrFmSzSWILFIUqeqwUq9lld23R
awd3Nt83gqb4WciEOBXCfN910jYEBxsMClTqDqalzUuYCyMA/AeGelKU8yBg
DXsfyb/QdacLZQSrUlnif2uzY4KoGYL3swGI3gPU8o12OhhLdWlUbhe9Jnud
rPz1KSKwKM3qilGRGvpcQRrdDXm3+TCwS8Rklz/G3Bs834n242zTWWO4mAEf
AQzuVtnVKFEzxJPKPGRJzHIDMHFZew0n2M8XyHtu0qt4n/ROTYpF0ZqY+1Af
RWTqxwuHnW4VpY3pEQrNzvZzwMrFtRyTtYZogZytZpUpwUVaEdEU+TwjrIyB
sz37PXHcIvPWUbnOcAYSJ8yAut7OVhOTAjujlXzACqR21MKjB2te90SYmsLE
ZFtgxFtDTwHcrJMfiQbWWlSZdIi5+ELDUU+5grv/unF9HexpLk6lI/CDTgaU
oYVOAKNhg1M/9/tNEwxfnNGS4GygE90LoAfhdFU4c3tNeDLyJfEUh5OhpVkF
THx9nalmZy1V53vBgik3/oaT4Ep+0u1TM4lzbjM5MjGt+BxFkt6baeE3BFFy
44zzYi1SF9/qf50hu50HAnknxiMm357EKc7HsEAy7zhOg0zgyQ1Yh5/uC+0R
1uemkRwH47YgHYh3nL8qi7GxEYuhYGVB7+H8sQeNUoRoRsTk7YQLxEgetsfB
oL9sE5Y5fnJ1PP9ySyDuSku2luu08tafymz11zU4ctD+V9ttINhaMonV9fqE
gVi6DX6pKn/DagGjBLcoYlnQjn4layxtMwOWEXuMsLwMRTD97yLmdrxWZdz9
AWuUJ4BJcDI7qBJeAIQzztYkOL8JSFUojuXAQkBZdLZ/OmI25gvo1piXktaR
u5AGtBQ8P2+5NGeiSH3Rg1DBA1HaBfPElNqZTHzriEgytl/yiOlrysH6QQ+w
6etQjV/1jmkuU0zjoUjiVfqL1PQn32ciSUazABXWnQmd1VB83AXgvMD510ck
6uCq9R/Kl6ege7Q2JkL0xREEXWIvOHi4jVGdEehIVp0iAwH2l3oYVOJMfnx1
Zzc3rA2u9x4AvPG3/sH0KBND2eazdTpnLkc1KBijIAXRRHNCqk/VDQWlZFdq
sssaBM++VTdBodD0z6waXMUM5enrRJf9rORU2ODKnzNLgQ2p0alMdm6u4btD
J/iQd8SUUCDzXUYsIpmdzYHALIos6uySI7vclxbGqJr3aushrZ1Gwqz90Zp/
6XRLFnjSM9wDBag4lVHGrTF8J/eRxXrR9omvMyqIcHjFE8P99RHexV8EkXfy
fQu9HUqZC2/L+E7MKpzke2vWReG68MgA+776kmD/x89QbuuOCdj61JR0OKua
Cfv0MhUame5IHf4Ht7FFShwZUVo3Iz9ETNX+ELdCI43/3tZPZ7J32GkQ7vkS
QVMWPnGt0/tI7isCqZgVocN5Fs8CrILqFNkfJC3Rqc5ebsBH7wwK+3uf8MDf
GvQwgY31sI2b2DVCfuwuw5BRvGJEmIR0TubURhyFS1ykxDdGKJPb5Sw+zLNH
r906FHnrjr0EX2wUNBQqgEHKe+47vkaTFfeHEtLKjxdeE6/P+gUVYcDH/bVW
mktYQbwDojlra2IBPp/YGqafEamJS9UQxNOQEE4S5TM57URrdTRN1Wth+3gr
wwBPabKb+QaDuNtYpvFWKrDmDkscUuN3sm0zTO/5XkA4zBQ9Nb1q6f3vauJ/
YyyuwnmqaS08ei4kYDpiLrsoTK+1FQEiHFHqkqfik8Dtuh8w+RQQHMwzmzl3
8GjEB1dhNuuNyN1IkUcFeUxinhd3ArpAE41+FxV4wZCgxqT9HNzVLrzLRmBv
WeppZ0qyU8zlQ7ocrJ/cXK5WhMZoqgMm3kulArB4NwwmzFKIo1DyZc9vol5+
iXMWsqUXRrbTB3YOCBjsMnvd5pCepohRcvw9YNfvp6UXezSCsTDsuWErSiDz
uMC9x18pMG/WIRy+7fyjsiTwXlOAjFxnAGY0GEhF2L3Yq0TWbAlbkbI09h7H
B7SktD/DNUyPQ25fytuPK8hWqDe1uiT4ffNRjVsrs7iisfP8Nmhh5DTw2x8c
QG0Xs/k6Oc3z3ccRK+CLmcxggzQNnBuPOAufWepmAb2cAYr1yTO2GKFFAKcF
uLLCDRq+aGryncTzlzTo8m6xAuyExKiU4dVc/8KV4Tkc5Ua2xXZAmc+9Gziz
vjz2DwERRqSZm2bHYU4N23CfVpYEmWxjtfVIycfO5KrDnPg75JiMyrm0OwSn
LKVECtft2dMxxvR5a07AsbfZic3NODx5SPuAdXiIfyZ9yLgFjFNzL4IPiV3d
68W1VxpnKxBcFXhwf0hUumQGb4mic+orvQ0lwWVwSwMjgzR6JXFrbJKur53a
sHB9rRTIcrtRTbB1338zPXoz9b5tTZQp84Uv0dVS8pVYvmdC/epcEVYRo0VU
/jqGmlXLVbL1ve7w/py5ZJG18yVnvuZ9lKvaAREPY68GBIWYYYpK4+nRA+aj
NhL9UFluLGgVMEsea0jjuV4xf/eb+Eu8z1N4Hvpx7aItqqfiBX9/gOv5Arn2
4r9TKw9gER1pEA8x2MWx3boF04MN4rMEt+s+CqcsdAHZD907jQmDcACo9ktU
TV0kVJth/a80g1O60QnFack4dGSY5Sfn5RfUaDgXFp0gZtanBgq6AceRdM37
HGllCLma3EFalu45ns++DMpCE98qVo3vFcYxiXFqPkxV6/4HjNYAO0rGXfy8
QKhXCTEfALbTqsvZFqzojX8cOLMzTPTWtgYVN+bdMnNthygoPMenw6OFpNat
uU8W1GP5IYwWvZXdGqT7d+qIekJtnJaXwzdQiVgKd1oh6OC964Ks2AgFAAWz
bjC9JVxvC0E7RFTyDBmDLuASnpgozPwhmw2xl50JBzFxH1FvJ4iGpT8JHkN2
5Nu90xS94Xhdc8b0G4pBch5Ccdgnvfq9/ewErNRdq03uiDiYJrVqDSjTfJ2t
SMag+Dhafdo95jSlqGRwqfcL3vWmJcAMudWn3Sb10eJPJynJKlW/BQAJUwxs
uuJpqRwvNBHXdcWaBJop+BXQa9j/yX6/bPFekuFnACm2Fnj7qJJX4X0Cpyab
wLdE6cypTIcGu8QgD2VPKdjd1X+/S0zdG53oY5hr6+aMzHPEQhbSqMFKwC0w
aFjwXmvCaQeGiHiS/11RQELfkpT1rGTKefGW21nRbCXZr/r4IWndYW46JdAE
wDjpo82VsH6z27yJ7gAFVBgOd9qspvZF7i/5s8Y4ATXbooa2iSEQJPuvppMj
TqY+dd7aomdZg7cXL75Eyuin/TPZmt11lrlyVu+FOCxv1jN2bAis3FjIlyVR
a6Iln0o0xWX7/RyiuLHIIvFFyojWT/7QTv6sDugww+RMyveyaHnnCea1bJDa
iYqynWt4kJ54t5o6pBZkDVN4avJW6QF/ScZFSX7kE6MPxmTRJ4nROSOJ6Iil
fLZwATR/JvKh9BnUqltkE3HKCISmzQrZ/oDlizNQ+HT/dUXzkSYELJcF5oJC
sG4K3Vr9r1ln/KdgOQMn3j5Ab/sDVP3u7J87IIldCSf9eFY/V06Ek6KABP4i
mXHkcyRwvdOfitiP1HM6/N9W6EjDC0CWeoqnFb02bnhoPNZnQHN1bM94GKJ+
860purG1gXW/XyWw59E36sDr14JDC17idu/ybBQxvylLSuYYIdtycBuLfbWl
r5yxioduRgo6qYXVISDP/umEhjdYdaDaFZGevitqfxS7ncVGc20ntsmgeg5p
q2/loA/8lMlkkQ5RcFiwRfq/8hvYt6fP2EUBi1O4XVBQCeL9X5l9MjBfMxmC
ZMO71Sp1tXTbN27MWQWo4HuciE9LHEDFuDIYaUNx84lXGVR6MYgCKTsOFsJ1
iQrZ6fs1vBC23uUBxnRmLXlbllnfm8puaboZXO/4W+qvGuY9mS8Kh5sGiOFk
NPb7YKxgkY+OCRyS54XArAiRWc/OmNz91Df//6O3m9+Ak0bD5OQ8JDPa6CWU
eCQ8b7lmNqcgNLp01OIS7WlF02JZyZWVMITqD530EdL6pNz5VSmsLvgAZzMP
njlG4uBZuSNWFlgTomxmM2V8uuCocVUQH59e4GbWFkhWFuB/vf6rDQACwUzd
v+kcn+6MlESe+PXJwV/37vVhqL7141fVzI4CS/lwkJD+elB09J2sKFiALSxt
bY1wpm3AcvZEzEEXTv/thr6YUnwJAMB7dWl+9RxNzBGUXFliuWsalCLQtGBK
mts/2PhLbROkUzkleL0tDfuuy0zCekGy3sOSw4guT64fdrTDDpFHBHjFp05K
ztmvi77y/aquYZxwHYoYorQoZ8LrUSxh46RmRDFJFiSpwMDkh+5UvIcSpSWT
HFToeocOdkKolqIVBUIsR9pqGsZsffXMZxrJ7af7Oa/FS4YexP61g0FwMWSH
32womCD8U6d2kC7cQ8p4SmMx1558WdkhKhyBDQ2xVuVA32u6XalydA2j2pTf
O/qzcSCiwrbb4BJWzswFzsIK1QMB71h6M+kiJwA6qpViLP15GBXTsWE+KO1L
luzwTrG9tBW071U6iIT+v82MRiPOdoNQ/1vMgskfR5eD0KnnKoOhqiYW42Fg
zAFktghZY0KupEY8R6/C4s4Bxy5SX5BNIT4bo0AYFlDcIKuBS1LMI++p29xT
VRqL4xHniZuJsQzaROwvms4NEY/wqDkqPumcXRzRNK+cctAwtCGgMooQonOH
TrTAFk3U7c+HojR2kswA5XQX6ORb7B1oz6f1sVWxZ1MB3f4b/03q1uW0QK+L
xuaei/D0tiW/1p2pIdox01JIYKOyhsxKqkNOCMCk6DHLzxyDJzhK65C5GpOs
A6yK60NcTzBqEhiMWnNEvOzfz4wQVn6kVCeUtCmwhI+hIF32ZJiuJED3U/q2
1wuJRwxqu5JuKhEZThU6b9EuVlKcR5BewKgG5GyO92KmTnNy9JKMxEbqG0YL
gYFbly5BisRdfbWgsWh4yWz8Z86k9MN+Lq/uQMZ+UrTRpn9W4q07rng2wrG1
RwVlohptO+aI8aD3du0uWYmlDBAbxQ8ikYcIX97V4tpJ1D86+KM7gWLyMKX6
qPChDgKMvvj9GU0T/7m2o+nfXTThGvBUrC3Re8k3H1p2IgFU+DvIo0gnEURD
w++U2H1PlxrJx9bsh0F1g6uCuGE868sa2jLU+3yekEnhrKp0LxZfw1fOvb8v
Vx1uhxYRhelrfwaiOOuFM5PZXxGXEMdoEls5eODHsdkgtja7MqhZnHcSOqpn
sXGd7J3hUh5a+FwUFuNf4gGWqu3q7Vt+I8R5U4/sZpOS9Gdi2Ms4ErAZkyka
WJjLFt5Q4Ku4krP3l+hoiFD3izI2BdnpvVi3vbvuiQ+vVtVlf7TpPw+KK7fE
3g0m5aSngr1HQZe9q9JY8Vmf77/nzhIoEDL4GSS0CuMWCozmgyQQqGy1vLmt
qdNWMu6c+lB1N7+oo84LuyqfhjWZBkU8DMAg7sZnkT43jhFhor/K0BiElzgN
+9XQlhCg0OB3fBx7e8KpIEs0MIkV0g2cD5N9MXD8m8JEtjKuqrlfoEHHYgHn
6cOgrQp96A9uNjnwT6Oeyb8ruRZZ8xmxVcQPdQ+0zqKTYDRKSIpkaMA8bL6A
sUFC/IoZEz8cBEg/H2U0OH6391YGWjieryjBr5IyZ2tUVpGIR9LrcderdWKs
3EWUCEiEWuU0kIUqySrT3qTHXMWM6K6hMZu+Y/H5KDytf5m7OWgzeDPrF8rs
65tXHTvsSTpg0yZdpNt8xAU6VCIUnEDy8XOLNjHS87tZ3/jt4A/ldEOglJrA
QlRVXsO+F/GrD+3eJ4Hq/ipotol/az3/Q/J0yaUgVHwXRTo+srZkmb1KThQr
r5g/24yy6G1LHrwXjwT9TGkb+A8EjDxhn2IcpRFq/PVtbfczyZ2UUtz3cSTc
abTxO6jWs8P3CB/Nk0vmZFuZmPiuMLdk13mSL7WXfHpRbkSGzNz3Bt5sUKMm
aOyx3HWNM/Lw9V+T8x7GDgsmyRk14HbrCHBWUMIcBnxtppJ3TYPAH4fs2Z+e
xPXZw/QWcqLYoc/A8/Id3blF+xz2gUBNcu+MwMBPLVc2ierF2TmB2CccQMw/
fGEkgQVei5SOdbvrd8Q9vLCnijn1rAwhMpavoIrWdl5HzzjOue7AA8NxWSAW
nftMNrACS/t4Ss2L55doHod8y4pHW2WzLBeCNzFklfErOifSkq8e1zPrGsdk
xyIJDyvPLm+Yk6uai4b5gX69PrOtfcerDwFtsbUsJ5CdQfbMJLOIeY6XMCXz
8ILMYmUsvAVYumIcASFjcaMcf7+JhVu7/n7xDGN7gsRjeYXEiO8a1LYQnTuI
dpM1o3t5pDrBmqn0jkLa60h/+J1ZyUHOopF+uRjwPuWUoQ+xmmnZAt32qzUY
c8r8XcIbCOGqd+zJtauLBmriyr4AZ67pUv1CxytZsi2MkZ8jSMrZvylMOqfB
Y50jxiDhagwvV5HwSqaqx8AuMACF40YmRiC8M7sEw5XRxpHsDBGYY27TT7Pz
VqVIvMr/u930VAm9Kc+yrDtIhgcWtAjKovP89cz9SaptalNjL1pkuQ8/yqE1
/fgEQuqzKHXpYfyeCSiRITOhUelQekg1PlQnvPtgAtw7mnmQQvESTLTTmTAP
B7aY7rd3jyROR/1MYZXr2XHhmcutG9FvmDEAbqfFiJqhMd3h+3vRMccq+LAq
DuEpwntJ83hHj7xDpM3H6C5O49W1jgacK1+oU6KIwzG1N2dfzy360Z+8l9qm
9wFerzdyYGbJc6ufxcrvPrbk2kDiKJtlux7Cfn0nBuK6+o0z7XyGhFAMgVPZ
t5LJf9bZlLpAvnOX1xJikgKT8PsaAJ1y/V2Xj+Ha4YJ8VEMwSBNImMEyICZP
wmENDO3iAjCGQynhlfd5DAvKnoOGgGSM/E+d4TvGMC+gvFHgV/60RQJh9EnZ
4lFinrxiGvhluyL6Ox2NA9+K9rOPe9MhRrBDvmd6qls1kll6VLi3VKJ+P/wB
6HUMch0E91iRNTvwUQJ6LI+mnD5+jpl69vIKf3mPXZtpCJIPTjm6zHa84DIj
hyA8b0mL0edolINXE+UWLZbRjC8tHY36REvBwf5nSrSPIFOtAlAdR8ZM/8gM
E6ru/gEmJrY/EvJWZg3criYOyM3pMCFlAYCkVsIRc5rq02XmcDsl5k4JYu3D
A9885O/rsMmFRsMfKAa5ZfxkX8VrRLISAEKu3VbYWEfQ23nuEGV2XcWzzGnR
D/ktgNXiOXdoH2B/EPxatjSICxWFn0cBDCD3zaKZhJoVrExXYFtwG5ssyxLh
FQ9ikjGhmYyHkoLx/DXoxrZeHZ0VU+pDhW2X67xim2zS3cW4jt86gEbfYXtt
oBthZGkRsaj9ymCEkhDT4HIwjHhBgOzXthxRrCDqsRThejCJ+ty5qBFDIv6m
7d9wfhqrFoAniy/QObNK3JncCSWv1t39UL/acv5j5fp9w5K6NfyDRbPSRYBS
Hejo6oegFz+6jlO7ARUiW6VmCjVX5/EP+2esRhzTL/vPNer3v4kJYJukRFUR
afL0ZG/RrBzwLkGPmdpCXn7Km/rNzhuX5YPLFeUyuouBa2DRUkN0Haea0aNP
ZJLtqB37KPdet85UfFrVCHJZTtNcmc2wCR2RiWKMTloRa4Gr9roxPX4xl1jL
oJ791fTnZxcvyMQKNzEI1Gw09+QzfKG//8larkqiZY6ZTQ/H4WiiXMCnIqXF
9Jr/IMsAkLc9efm6TX+/OUjZAbkLpP4+13H4TNxSnjfxKC4i+vf7SgP4kyt9
lYo3wwiHFW4P/rsBYcIhQbneIdPfdWGzVlHt2HXFWraD/U7XKamEK7UAyNrp
l1vXjCwJYRdnO02puuKw/sRmnIyk8ghmu0seI+SrPMuhcSY7r2O2devw2vGO
j7Oh67mVFPzrPL59RyJvtitPZlnPVWvbkkFLhSPpSwIqhKy5g0C4Ruf6jGln
lw+BNnwiIoue/y/7Ec/V+1FxrTd0MxfBDx9ZdvgWiviG3sZAIKfTzaGW0nB5
kI4yHZh2AGTYhJExj0i+QEOXrt9Mi28tCG0Zuw9kWrL4QGcgFh4w93610A64
IaVfKoWOrT58u48jO/7C/CsSs8nVoG6bB1B0fSMzwEZkfxJhXVJlUP8qQ7CB
+pZSxYWXDofd7WaioiL9j/GAiidsZ54tgKcc6KcSWbtqk5rBs2oDBdlVnFIw
oqaePQmhvbG0eMh6TzF/MFFCsYYjiIzoZo/7mrbZf05a8VqkWwIi9uTR+w2n
BM1K7YXhAeZsIahAIHs3FeyjCAGnZsyd3vrA853yjpN1FANoI6LEWPcfehvL
rQyAVp1wSQxwYSBLvFeob/SOPy61DUFKZBi7oNXVMR6OU0nm5K4qlwqv97RI
wFowA1w2JR5jjzA101ATwpLkW6kX5kuj5wwFE/mpkxYdN3r6cpDWubcgRYRk
9x31RIgBSwAzduiT7ZK0pEbjonIz5oGpAB41N95esMQ9Yjiu1yzgnwhhmfIs
hIpRiFMH6fjhz9xGQvt+TmTfKmcGhEicuyemcdlYzD7/qUTTSpe1suA6wuU1
igf4PPuVDRD33kFe5X1QnZOS2UEeYJVB014/q89E7nfy2ByhhONATh1tBras
pzyEfo2lp7wmV0qUfyoIQdSr6WBxxYWKk5yO4KieXy+nd16af3g4F2h+p/HU
M9Zha+lmSpd1RPmUxh958LZo06gzTeDbnGdbeKa9UFQ8e+kguU324v2vW00a
QknGiRFBdDXU9gWr6oOcvHNc7UHDY0ZKJp2nd6ibi9QDEEXKdAez5lJLvNdg
MEY6+OEadUYrPUqorhDSRISRIViXopwxC6uX5zb00OUXCyu/VahAEruMDamE
nRTBJupm7zQ5A89pN1VidutvMgq/UBx1RaCdZFHQsfth//vnbqgMU1o3sYZ0
h9uRVj3VKUun2ppTWklCej2oICkFEBw0xzq5VGZDaDHr7R/bCCVvA1ElU0r0
1h1DYC41XABA1D3AADDFNihrk5rXAvlbTqeWNJt0jPRI3haYHJxvffsc3Y8j
XN6INZXM4eQyPHtsusea56ANKjKY2Mwa4+N/KXbNk8OZjjIltW5VudscvXVs
rI38hFTZ4Lk4qQqtK3hIAyUrt9WW1Qiw8W9cSVW0ZcBiqLCOnSVFqt12UlKH
FOewf07GDgTiIdMytPTusrVGhrB+N69tGbfBWp52+5smyJpqlLhqc9VSAcGX
het0qgaZ1aRZ7e9MV1ifluoJmcVZNNkVVDxWYE4OITscvC6TrfaU6b0zR8zK
sCpjvWSjwBSGVm7syC4sSIiepakdYsJLIOaSnBl0RE5Sw5f4fGz/L3JgZxWB
5OBd+B95ZkfnbmwbFh5i9/tzqvn76YfPC8oEkAuqe4nuerdOZRIAVAyALVpx
Dlt+G/owOUNEnnpmaLoR3zHm5NDFMBvgvEisGRzL7mOV62o9L5w6tImpTvHg
qHnFdFGC1UCoQcrDDdSfhrzBp3cmYiyDHXS9DEaL2tyfC+s8OdnvGnbXseoV
FnRI2KM8efYplUPpwVg4Jq6/2ytKOaLbvYvxGEDve99fQ3oILDFN48fBa6Z3
pa29c64JH6obDq2E5lzE4+tV2Bv4R0BGQBDxDUSrID+Bv0CsDIj3KXZgoKX1
Mb2Q0IadYd1P4BQyMpWfu9UN4DleA7lScU1ci1t7Gfx8wauaVCH+mEbKc/mi
TIysyQf7InhjV8nBQnfcfAazMKjLw/6ozLN2kb80FsA471SWUQQs64UhqQca
N8/Fo7vtaP3UPp2N5EO0PFvZZyfkZOGZrcc5o+g6vKQVjuTDRGj8BmX7829Z
+6kJZqsZbTyaV7EorRMy+DXcVsvtqNVlb4VMSZXqUWHlEMKWUC7dj838ldfC
DiBvZeNFYqC3rYLI8pVseWmSS/PClR1iD2UHFaiNqOlVPfuHoukHlMblL1R/
cdPyfRk15YU7Oj3RKiFWi2ER8ftm5D9mlo2M3LPt0Td6fnMjL3wQbDHOCTnV
ADfee2y70JAJuFqDez71+ECXcc32S7OOIycFnA3lpTOrNl99U+0vjbVUHtOJ
qGdxzI4cWGmQE4yd96BpumP1qY3dBCttSikqt4SBGh86I300kUAPUxct3V+f
CDob3RriTJJ5pZbiQhy9q2uPxXki8sIV5EjBiwzliCgyoEt5R9Wz2CKZXzJR
uaUsHAkq1F53hZEPclbqh+HsQpss0U2ylxob2gUwqNOrZRNAGdfvi9Hk7xPq
fYRnv9bLMx5KgFBqMZxvVdPbyUEpoMt93Ai81v8p8LAAf2LFSSBM7rbWlWBd
ROCBR4HSvdpwwfetDXvQK7o/jobL+Im1JW7afrK4xjRq75Ij110vCv3NjF57
RZ8bHISRv1ebYriAROZ6OxHEk9mpWbL/HmWg5x8LwAnjeplbMUL/+Q5xvjwT
mBZOoT9HiR6lb2mYwB0YyAdX4AyCsq15WrZVI0BHg/HH5eEIk0CULkeDQVwG
s7ev79Hhboe0d18Cc4HOoh6Xyd9OmpGzTUQ7u7rzq9eI7c75XwAivWew2bWz
cKpMDJkOS4c8fNUi4SN9XTJqBQ3Ip06oc7kf2j+8PZ2XjEIuiGp57qm77TvX
lJxzknyqcVG/Os5yy0yAOq5roatwHghPTdZ+aK6wJTEttKhQExaFT4d6OSAL
VrljuB8Ii3TmNQIFMk93vwwDcVbzrPS3sgMFTXgtl/O9rxy6grGyfoAjXu3W
y1oEtd9GhPFSuw5Gwx8NuwbMIKWEZeqPaarrkJO8MaIr41lNoOROKqB37kEA
d2zOvQUiZj5lh1gpeHnxswJp0m+k89NLh3B51wc3Ukin6SFTNAzJKdBUII9P
qbxxfVI5fhcdi3JV3EvTaGrmrKGzoERh+XRSA7ELemWYAlz48RTyom8GhlsR
e0tycRPRKFWqUOcZJnP/Q1MMfkDfHvl45d9Z0Eoq0RHfpbptPGmpZ6OxjeyD
sZxXEHBBDelkoHVdWuc61dl8WC8Y8uWb6dO+I2GQSB/+7kLTXZxNU8hk++7L
QKJrHbevZtTIXpvjTEGF00gDjyQTQOnsrJbFfUA+kcvWuHuHB0djHZxAf+3w
XVhUF1bYiXQ3WNEZObV0RZxF0p7eabM+vzarwpDq2HB+U8R56DqjtqWhVGRo
biFXdZockv8V5cqSrStxegxYOuKjAGikaz0L43YY7cphyYcQcVRvIQTUVkpe
lZPOkxcHmV2Cv2gUDmI1B5Fnnopoj+4T+EcUHUifAW3ACyIRIpHQ8xsKGMjt
ApVR+uI+xLIQUJTgvjdaqXC5YFXxUZ7G8dZUQLyKhsrSCmV0FMGWVTq8BaQO
KAA7RQIjpcavxw1yruMi7YRnrETimFquLQfYWUg1pnnO4fb7k5HKIDxcyFXV
Q2+uxvSOOwWgTIuYh8hasS+H6lPCbEYD6Z69TmHya5gMyQfIiXVaW60VNfBL
oftkBJ6TIA9tV9NWSXIL3XqzsXKDJlWmwMoJG+k3wqHpJ2URCqAOU/ZnMiCp
kRd1zDo0Ukh5AuHrqY3sVz7AVE2D1QSExZPnl4HXp97Hs+nEJbLcEOkIBUzX
vQn4gVuG9U8g1HBYcCAtwQR1R7bcH/srBcCFUyudXmGxn49cY82UsB+OAOBh
HD7UI/gDvKo/Djo3KTxDHWf75aNGFAtd2pmuOm9PWRH/w3AR6TG5uDzr7FiG
3t+GKcd5pWDT6lVSG2Jvtfh6AL7OagU4WtZZiE0YXN8VOSN6H+mqpWN0QZ0p
rBs4/30qWfZ0IAz0RRhDZrm07iWeYKnQNKo2S6qYC+qzxEiCUyEkBdAqQS3S
c1dfzjRlLEUhS5KzC1IXG4yYaCFBLY78ydXZKUOpSVp6yIYkcmOS1lDXE4bK
ODMgeUxyI8ylT0h/UcZJYqTG/t6jqJS+JbUWemOHJSuzO+7zOsQHknUTl0T9
Jbpj+njBU0cNDMO+nAQyUNCDcLjFoFLdK6GSW7SxZMUtFlc6LI/F+lfsOlj4
fwQZo9ykzAJTEUZ1F3xY1/uMM0hQ5kXq/xtWTPWryjaPTqlgHVx+j22BpxqC
m5gavHsGmF/zkt3v1shwP/D8VeYdz0EdyBYOEcP4tQJb+GW6HnjOOL1Ff3dd
szf5MB3LYhw7OUB3OItr5mrEaTwEwZmBqb5MJ90n3M2QzPpUjKNNRenKaW0Q
jM4j+xqSsVvJaGGXOtcXuSh+mN0FPDUcohGnhRHC0KqsFJ2Bv8CTmKwiZ/fI
HgJkROJ1oiq/ymSvHPLNE/mcFo8x2OjA8w0qqcNfgPi9TqW/yTQbqqCZaCG9
eOZ1HXGV29n162cJ0Lwt1l2GFXyQTCDTYX+D8ySs1XV7xpbMuhsPMck7iAWs
DwAw7X5zILrkDgylXf+l2eNSIVmOeMWPE0EyCZz5pcJhfQYFmAh/WALASXnJ
8RFpI4dQ5wkEY2IJkoGVaQUXAAXUPeRAUiNNumY0/+XGS3pyZibgQ22Guv/h
oUWEvoEW388rFTJVJmsa/8GnPRMK5NpR6zyyAgzWI/KWU3FABGQtoUE1bh9x
U8qttK/hjMno4FLtpY3q0e6dv/uMzlMBR443MmpJ1ux5VHWwqpmqYP3vJ0oM
iQZbJUZ1QTafJt/cud0I74NwHs6iacjp+aYgnDqtpJi+ldunzeRgnT/XmN7F
1ZSMNGp5jzogXKkFy6sSWd7BESBXk7Dlen/z8296Y1182JSsCNFRnEK9jnfx
caXzkD3KZWeH4thtkKnvipYWDoI+LP3q80nbhZr8BdTHWYSt/m3QzPZ7+lBr
1E4egdVwt+Om5hwld992FMf18juNPpcfq7GBwA5+rEY7OwPwT0aRRp+8rRAp
lbHl65OOXis4xjJdCBFW1efa2unvzTzWXhzJ5S3IL5o9M51RD9nU0Ldx2Goh
kdgiWCyvTM/CIBho/8O7XpJpTVDAr5L7crY9xTft0FES+nGYDp59yBZnF/wv
5np0HYbyHfPkeD3jjCgd/fEuqsJND+Q8/rRq6HaB+5er2cReNOzCTK9BORRV
2w4YoyCTXtBUoTXoScMaKjbHyCJ7F8CImpSWNxAv3p8hcKWSW59snKr9QC1c
dzN45Qhza+40Uc/SEQxO28wTiGfJIauo40dql4ltBqtZ+XzChUfnKuZWSN2H
hKf79uu3Gt/uL3LNRYHpArcO1c+oPE4ngByN/+8LGDqFxLFo4x6Xs2jFcLU2
Xk3HyIthIvTDqSgD4/n8sSiAvVP8g/Fr1v5Egk5dyoeKegVDbuLHqcKL05lS
6xlZIHzxz+2SqWOy+14VpZKQBSAT/Z6Kj3LLCCeLmH3dvqWEbI7DD/Ea+cnt
8BFFrY983A1xVbU4sgNa3Sz7dybLYQzmG0cbgMH9X6i7lhs3WJn6jF9cs01N
JjfnCT/xPFrtovg87tn7jictLS54vfRQ2WGUEL0TxpFWfk6umv8NpRs3hYJY
ghb6WvLAQ7zXwVkoFZGZAL/4Su7KLbQgytZMcC4dKn14N+0j5GQkaknFPDaK
CiWPWUGub+QbKNF5KepAwf3dCVmmWtVHvgtq6FfGbBDh707TwB4uiSu1IeQ3
aCe2bSZwFAyrCbTBj69IwbeYIht2bbL/OIgsGIxPOjYQqe5Zx/NT9ZjXBko8
qouhhwPCQh5/OUBzCLRuFS9xZGEhULJiD/PLguKaMGOjMFizMeU3pj2i+LGB
wTuheuWUkddpILJtjd1k9ycdVSztrlDFzPe8Ux1NWT1VWMP33T0X/4usBn4J
g75HkzIiM/YqrY6NNg6/69E986sjUwfJ0ZZnArxs6ANjO1Recp4ioCan93ca
YhpHyXUcgPlLmh/pSCdsGe4NVHpoDlJWGzlt7cGWCTMRbybeDm8c54DVGFZm
9upzUneK5ixvMwdewnSZMQ6wAx95XBt/ZgdFEUWXfyvbTdEg0QatBeaBEOdA
0B5FLMhX95aO6x5pQHy/ih9fUENGUS3WfWre6uN9cMXk/FlHd8WOkPtl62Wm
y5uhmuBsAqVZw86CmK6Hf7QhZqnBVDTexcyzhDwNY1sw35vjsG8RDmCteJlG
pu2JXS/ZYwDR2Wro9rIjxDNA0200L0cabl1VQs8zYiqEaM+1YpLFMQQGjJMI
kzEnfwSNbB63F5S30LBh+x3O0aw6bhhO0I7cfLNRI92Sancm6FackjlsIrZz
jbWoeNE41ugZaCPRiVoLJCcdlmVRhfC6dxtidX9rNz5qweAljpYalvjjQ9wo
6713PcJ2yfiW3iL7MFowGqk9c3zoUc0OcMCJFJmroreLysh5tM7BqjR8Z4a2
KTfZKuFzqvlDhDdrb+u7OHxdWiWg/wJn8eNcCnuAANKgpAKHjPMJ9QncVmYu
WW/91CwkAMp07PF1aQrzU6NQtyj9Jt8NwDL/K1UNTPxm1v53QCGe5aABvHQs
fxWdJRv3Aig38I3SOUmSwvBzjVeUFMMfLn6UcwRY7r+cHcu55jjYsAYLcO8W
vBtbvP1aRPqEdh/d7bv1ePl24mdEof+qfSwYjpNdHQZQWyj7cs7CtwXIQ5uj
cc8UJpIgKdxSP9vxCTU/iIFjXy2uV/lILadsb3X03pLtlOiepeMn4ae5eb9P
n+wG7vKZ+vaBIfcFsGzcL4785G18VEmzp2nefena/3URWdVRLZWcYai7ces+
UQHCHiW1Bk7x+abhfH5VxTi1e+PpdVco/4tSIuJpb/7I0jFcKgteNITFrC11
Bw3V7NPC1W1PWArlo+Wgfx7APzpxoGDxMCaYtfwZahgRR24Hwn00t43rRJf6
8imza4mWCydaRxLFnsS3Sk03DAD+k4L43I8tpNEpvliFmYaCpux90QiHrUZ5
Ll0COuJGUMyEKI7ra9eh5oFKNS5jXii2o6HJ1k/FOIUuNgAdvwHOEXSpWKsL
N5t/DIzsCY051xHCxL8kVeTTnpke49IGZsSmOTbbCjKwISIJDciQX1WoTfi1
xiW+pJS+q0wpddGJqmmjjid67FFukYKrl22cLuHElc3UYaBzCglALNGZ1fsB
e2xs71m8iQG9LAG+wGYSLm80+6nR6jk+QYCTp3LnuPW+/KDB2aBdayIPYejZ
Hz3w/UTZ1/uCpEcjkn9M25hOvo8LIwWAzdn7THQ7n+XrfsKpobEZi3jAe0or
r28KNDahZ53RPAAZjI6hvjNXjY6+ERTvRAvk2sXKv/kuqBvD9I3wQDxxqwnq
/gjN9nxyZ7+T0c7K1NIYI1ttU/hDWHRcPK1BasCTDrlLKiH9NJiiILiAkC0N
ainV6APadudUiF3fDoVVSBG9gZBCHlL2sQnpcoDgnt0cbV0hfkVRqHSXMQ5Q
DvGrN+aLEfPvDCaG2Q9gYrQCIti/WbO7XzHQb99uhDFWwYs0D48TfotMK1Ut
NurncaSATfxeQwD5WrKop+SOnRk8SQIOL/pujVshstwJx/hhoXHTnBNwVmCn
s8dSuX3lfjfnKxcRitL1DrYF++YHX3cBI28roFCPNQGSr9B7d2pjr9dfjE3R
DYAI+aanBNPiPVXCuhDxvlQLDbLk1Ku03EpYBygmiSKKdEf1v1c03Cf5Yh4L
y5clR/PVgv4pLKPeBmbMsafeyXhsKB/FbRhjNMcG8xKRVmNKuUocsPSba/F1
Vu//YsxWzTnXB6zJZbsZ2A5rJfhGwiPXMxANMrSrRdtJyCdBVdLDs7yUxK4P
Ey3Q+RhpMKfy94UYE9g9D9AJfzjy7d6sWoOipsswaWp/VgpOvuujBm6Hg+oC
tz+ubpT5xEnWiS05MU3iFbNkUh58iw3uN5TzmxVXUxocvOii7GVfbKoMiHtk
f/SCCJWmbl4mXzisCzv3XHG+YIEN1vkDtMHqLOhpF618PasJw1ouiN/oR79q
jP0aDJuVV1Nye8kYzt7Xh8a4klv6ALVRqnmRq9iQIB8wwvbGQ75/o30xdluS
gK9mKA5kYBJk/U7h0v4IjUR9ddo/fHfoQjl1z5fxRXG8ycfFuTLaaYQlzIll
Xews3u4yRV4iMMzZ68VF5wyDG7biDsqU5QU2D7TyUi85P+awXq3Yl2waX0T7
cjbeJBY4eDdRWPKLcwq1/xiUq2kFb3XWq0hXzlej2xnm1JKgcE1ZN3aQZhdC
8QRNCXkDDs5QkDmakEqX4GazWy8ulLexrdkElTUjI3n8OiNMJJlQwAYKttCM
UGx2EeQu4EDKbNRgBkSQmW8k71GyIjwhE5QLBfEsQ/lk0ARVV4jNa18Fc6YL
K4rFr8cFCwO9uIN5aKc5X35MehCpBKFFseAqN3WpglgNy0GPCZX2x1Qks/KO
QzwUzfc++RWiUj3B1g7S2aai0hslJypRLHe3h3KagKGZ7sNPAiMO3i4i6qvv
Vf7N/lY5QeZVM4KhtKXRhnR5/kY1pch43fcjHFpn028ZeAZrlZ+JlOrijBLB
CyWYls8KWhTy9vRN67W/poAUlg/m/df+CKHW4A16k/UDD/kIzoi8I4wfFE4X
mhl+F0OA9NXLmkBRJiNRqnzD94wH5qMZTC6+DEEez7sdIhgImDlahcIJvNIw
/6muz/pO8pbUc0D9BLZhGHH9TbI7wHyq5VeXBA+rWaGlZFQ8AINjWF4/H4Eb
FKw8bH72XzC56metUXLYJXM7G/njqRlCPqRLnN2GvD7pYmyXVg+nH1B+1J0C
yoy4ncLP6HR5u3odYHhKZn/91dOEhT+D5GuynJw6F62T5Gl4FmDu6roMoUgc
gwnRIGlyyQUs0i2G8tPlUkzyTlHG8s1AfRmuXTL4CwInqHHXdk0jCfL3qfWR
4d92PEpoVeFHSmVrRyb+4daGJOESZ30Gt6VHuEggBCGcewCJ4UYg+ygFG26b
mtA6cwjfUntepzUzE8T7gH8mPOoNQWyUxb+gJgY60ww3jFIdwmuI+HfXlfTf
eqcD7y890EJr55kQkTh2flGDKsYF1RMXv3Ez0R0X4LOdtKP+3hevLB0KJ/Rb
mFzbPBvZhWMrTDZj/HbEYna90fyk9ZdsOJwkFP7dbqQsDQ6NZSR0GSTx6v7G
SLK61DtQyIQ3EC7eUw/lhnEqq2CGplePBqMv4QlA5KBRF24DzwYBt9VxnDet
v0AUShNxHK5HR6SqV5H3uOFHurQIQ91pdniQMd16YtGldn1ni5DVBK/eV4J+
DKDWtgiR6jzp32s/QhXHpxCkQtq0MMEYCQuq/+vQSFYf1MJjd9Mply6+FDXG
yfecXIORRs/l+t71HZpEq1kqjmOFAfildhC0Otf5HJ3YJefsGPG326m3wCPX
JzVQMaYuTW9f0zJbLc04TC4lAUW4Rx9Sz9u7jS23Q34gr4XG+omgmkLPfDR7
DnsVpn3KP2DNFA/lUSsFY8dUgvdUWzWyE7T59JXoeJifSDv6iwjGmnViEq/P
LO6S5/qGGCgeAiIECsZprpuVar6uGONSWZlN96uzJoeIsLcPEDvYO/qT/4vq
k5ItTyQLtw5pluAqv0aHngeojDAVEeVZOpPwtSkemHq0kXN/cNQwKW2TZ8I0
q70Qw1ljs1EqC+ScMW8FTxS8pJ/BHy70USWuA8HEHVhuHglWZICqN8zlTL/1
1bi8TjCxSnTYw5NnVvnocQ45yUapGnThKuDw6ZuCBzJI0hP8P/IQYHelRPGv
njnU+cYVnBqB/mAAZFhDguQpY/jRfVIE+YebETmLPNOZGHPQRtmf119eZhGk
c3ds1+kYxEX9JuLQfcm/J103zseNaRpXaMSZtbaPLhKPiwNpXPL0FB6Zgsen
oAYpLmQ/tp1IQrw7oRTBsT/R0lHhBpjaEjgQafpk8Msdx1uXxtRd4drmzaoh
Ld/xSi8hcNBng00ze0K+15fihH88gqeEyYoQS4MlTtOeYxdwhynZiS/Ry3FE
eT/b2l0wbHMTzg3ZEL0ww6vPOClF8gB3U/XLtbetuG/uvSxUp//lRUdR01Vj
u04OuCWGu9YVSE3Usa1nagL+XWnBL6vhszdsoUxgHgTxP3GpG++U992rScNA
zQ8uQIJJGfQAIhf6cGoShSs+2bgcRuWUXoAJ6eRoIZ24H69UBrvrvq79DxGU
oqfvbVyGyrREyooIcEm9GxWKy3weck/TfWc1tMOsSavcGu36VP9xHibVvPrc
0gHYQq+rHqFNodrG7XFpIPPTqtqG45zYwqMljWjyQo9GJhst9qPoMNJnvYe2
D38/2VIYp67IBho6iZ55mrQt2QiOkelSIc37XXnGyS73Q9jV67BzUhmr6ayq
B12BlHHcsfsIRJ8SjhmfFLRXzy6AUceqtYVVRE3vVFAaIekd8lEv8lKFfjSJ
F6ytllTsKzYMtcl/PjyCfOyQ+uRezwzBMN2KzuW+P9ZCEgNqn0FcNxjqSY9Y
Sp8wi7uiAykQ9dDibxzKiJFhro/kHb89S/6yKZIVwkfPmyObl6UDPO+EjyPj
HOoww7EvzNQjQUqGmUysy6BTxRfPSf3/HlKQFMnpzaQ4r7+vyX5wrkmDL3KZ
11IBIg6LAd8DIWn0aPDme6/bV31/vypytDQ/GT8FtCr1DZCoqvlHew9IXqub
3g5QB4pngkDKZGG1LnIBQe7VYiWU9KvRoqheceMBxrna03RMMU/DHuu2j4xu
Y9sUvA+ezInp1PNo9xXbx7X+2+LWuQxop3BAUin98+DM8p2ahMwDk8pzJsjL
nkygabaQ5FYEXVDCb5K4qKsPKN+16LGfZPxiJ2LYJhdlF+rhfOpyZsJl+rw7
E3gWUF2+W+QU7TiNBuzBMV4edqR7kYTjiOlKPMnkPxFyFqx4ySw5gzJHSZKq
PCjMjdPIGP1RYEgPml7sWi8QDUy+qbETOUYmf1oJRT7rYHyLLG2ozNjMnlOO
KYw2+5/50AL3+eBcu8xi/lnws0b3rXTKegCNTnvQH0WxgSLpL1kKgHulY+wl
GxgcnucFARD33ALXB8F3Fn1S0xTtQ8IekzKrm/r9OuO//a6hwBCCkqWR5bNd
Rp39fwI5Yl6VuARmRbi5GGGdvmDNU/UXK42ZeH57nn/v8LFGEKF399Kdr5tR
qVcSb78Lpwqa16keSGLMk5Ral8qua2NbDdBpKQCYwruRRJ1GLAFu65jKx58B
c9ep0F/fBdhaI/aRrUnEIZ4jFMGAjjMRO4LK+tNBNJaB7otR3a+IvehIDbsD
tAUgKXRmRqoFfGuie7RbIeD+JDFzA28gPUBuLq9j/0o8MxH20I7NZKnL4vdf
0LhhIbl72e93TEJjnsaZBlXmur6ANT2yn7TYJeaTxyW6pCRy7s2uROAKnnM3
2QEnrfX7Vann8H/24owKIu7mr/bgQQo0XcWnHiZdjPnazLlvQBFsbdmYJenh
Xn9XzgcY0uBC16pUUbNokjmX9IqBhud0EZmjOeDto8Zu9xJ8DOpZBAwMAL1Z
Fza1bgVb2Izjj2FXcF1Cj8+A0ilG9qpp2CMx2Xgr6Fuh7o+R/34YFIpHZN0I
/NBofwqN0gHy8WpeirKq9jvRcLHnDRjJUzGw4cIlPt6z/vj30I3LynrLePc1
lrk4UzkAt47j9aV852hk8TfbrgXiVSEzW4HPZBgmlq31cn1DKternyh66z/j
ahxlUMOKkM3GEvuoscxFa2JABTzaA9RvgNndtyz47dAQw6joQohBU6O1dysJ
kh0VUjzPM0KpFDtOtrk6ugA9JjInhgE+SYTEmaU6yVUw/qRpOAXdG0akfQiR
/PUFHuZF6tabjUSmaUTyvcmFpuHX5NTj7L3VulQ4CmQRjBEM1sfNfYi38eMR
crKn28Hj1T963JPA+clRje7Mzc+KwrNOcc6zpxNlVkXU8hhAyXoQM30SHR8y
9KEuEQnXhE0O4bCcOrF1eGIOqeebDeqiqVicUcumoMFgYF4nDn/yUW0dyUEx
dS/a93744jhvClTTa8jNJLD6GmVloNrv0Qmn23qUjjeeeb8trPaBDfvYZkYA
91lTTB9OvKrc3cBDUxnVR5UfboJFX680SKlTw04lmUgqPtIEiWhfbsQBdxWu
32DeASYyWxBJ+gnMWp+X/vrGAk3JbwPOtXbK68jaZ5m5xzafKEIHI1GBZopt
lGHN2PYFrvM+ZHo8dhMcr1rTZetnpRNs4YXonXxDyGqkxJMW+u/0zO8A+wj9
iLOq/zkRv/qaLZczraS3D13nnbCAJzNYWNW53JUbkwu6WxkP03kq3bKuSt5M
GHQ0tS3bEQpxCmvkxdfp+US7FKtAXfZ4N+4Z6n8nYU+vLfDlL46tv/ruiuyi
yzKVsmvE6sdNsneY1Yh5/OqZIooYEZkCSHA6lxnqriC3fERuZuzt07SDe2YM
mn9A6/msVZCDkiREeIKtW2yob/SN3EZScEn0ohMXnTX+3eoOz2kk/jpxfTli
qBEzj1viI6B5Nw/db4rraGBuaqDsg68hoSO0SjegOoMeISp6nUirrCU3l2+D
Ceu4z2MqlilzolLXtrvzwmSQXZLJeUsKzO6hA8FfFHzVBlDyv0lQEb+sM2Bw
Ae6O7lFt3bPOSCaMb9v/EhG2hRoWIaPgpVL170djGfAdGQtVR+ieWxjGZCXk
5dpV5EfDG/kQ84wqC0dWJWefzIcpPrNgG1ib6TFNJxG5DkfIcOrphDRuFLHe
oZWCEKqn2NMEw3MBxgiFhyWZxsbJhSqcfWRaViD54oi+btgqUrU0MHJjSOif
Gfbknr4+7/N4YHhqvfNExxyQ2GAQaZBObYkj5Ipe05aueDz41gjvYf/5miym
hWrDMAanbTPeI2tpiyZU8ylHwm61WVPoJmBe3Dce4MLQfLvWJuDv975q2+My
ZcJHgFNj4CKKUJkSIuoWNqWoCMz7BkOri6QCbJDZmReyRfQJ+c0QqJyW4IZN
T9UhYZ+MqU/jABVoLNaMzq1esj4gPjab+WPur4ogZRBXPGe3rPt0u6CGJ0d3
KxxMFa966Ucyjv8nbFtLeCQMVKLpAAKDh7r6WVvGdqBoHYFvdHCMfiM5DwB4
zPqF+8hcbXg9i0Bb1Svpf9AEEyUllnqKwkAQ5wophI7uvUj4QwiSpBLO1E6Z
Lntnob7f5mEb4K1Os0a1+muQ5eMU4N+4GUQsFTahg2xyMQbyMb9Rx9RUmuOz
3vGBrfsxJCE32aJifp/rxtEUYrLdj+lqIB1zVidd7wy/X0LMw0ylskuZz9TU
uD0JYy3hMZtikTIQVp8niSozxdfObjvfbqeeU1DjsOSeiHncLeZGKxjSeR6f
UmK98vN7slJ4iyuftE1G/lgXRlnYCMW2vpt2W5mQLb+MHcoKXfy/nKgcmrYo
N/VUPtb2prmbksbDTprp1bGxL8CZt1DsFVHmF4kBj+/ZWkocNBnf+LWLRfEg
0VpRMsiq+a2PrTGjgTPHRD2oZyCg++A8sA4PMNF/cVUljIDJbj3oX89k/EXg
r+s9voN1h8GVWzQD+LuuIen7j7L2omPN8NnQeljaiCFnVDqHyM45a3lDBkxu
zokkt1zQVrZoiEncdegefAWr+L+UwBiDCxHovtHT0oU5+zR6v63VNfFDgnSm
1bsJGaHH13czt+Zfo2VBKruNk9gLbGn6YS9UZo4jh6QcNSgzFq0tsnPRFheN
3Qz28ig/99Xzx8W+4bSxu4XwKT65aK360thJ9jgolMNzHgetOlHIeYI1vMz9
ysZui82PiQy5+wd8/GhLjiYamMypromUiDl/VyHmgHTHr/bF9vRRwMDS4Fzw
5Gr/YRUgki9BizzSebOuQbEoFvYwH29+Z9b96Ig9IzA+hJk8UA0rtypk3Emy
QoYvrJFRRuvogK4dE41kZyrgLqp8mTk+flZsIrCOnRZDB40EMcfIpRQCaj7b
9jPeUj5yelavIQ+2mEY1mqcIDy5c6PDnwz56waPWyiem+sIIXAC+ib9tL/j3
RlMU95Ayi+mRpiVljVvpch6wq4gmJiwbVblKE6q/m9QH49wwTa3wyuHq+nUV
dzHLX8YvJVrxX/MN3QfjALxBUzzNiD/Wsb754nMZh+ddMeP9/OLKIygCCYOr
FxP/673KEfk4MBfvb+xIFWJyctA+KHq2unl6SSn3wMvY/l/HoiJ4P6kpPwAA
jGm0fC36kxYB5U4gMyLR96/ZUGV+u8UDcG/z9xLtk2xwjwFmwmjsbJWJ2VDf
8QbSqdRZBykCECQyxdwkBE9ZopT9tPQee5VU/ai73VAeQ17zeSQAgg5R4dKd
nCAbSNTEy79AqGC3f1vNnBCtqbobYT6Tr7zLcFxI1HozP0SOdb3/6NssIwbI
cMrIq7P5qVftYP05kxPzzVsQ9JtPuh7/ajdBvLYYsuGGdPTqyDi7FNiWxqrf
unBmRhAH1J4UYv4YmE0pftSd4uqvdLRuhQlr67+/bXCGVgbVNdmyNPPoxeeI
k4gcZc635joRtj+Pa6OhYituJ6BYpJEs8gGtSRPJNNleNbx9HrSiatz+zRce
4PUcU2AW0bdGJQ/anAmzgxHbNkbObYhxLKScrygQpKYBhWewmgNmv6TYFnpe
SvFr4xbq09mXeamDN2KXefrqbDkkdmin5a0qM1gEvxsBaT8sPBvJb/kwHCRg
fVQXEx9lpNu9EL+ZIlWJQCv/76vzQvpEv3GwUw+1TtT5QvBEbJU6aWDva6VL
njVQRexuDmgstezPpgzsK7S5tvadetXdARJUteojPGpZ7DqP7h/qJmyUu4t3
+/NqRjMNBrpT5RcN6V4F3BZMAX4FUfYjPC/txBFe8HbJQkZwcc5mGZyAn92D
F46PwmIQ3X5pXq1q+zfVTfJj3xH4AA7BDn1sON7x1a6zpgNl/aIf8K4Un5+Q
P5pSDxc+PI1FXhHfY1H8eYe2Y4FSPh3C0KVEfhcz1GWRrcwOEXcEeFT6Hz1m
7DWj3lFWCmafzX/zv5OtdU/MB71QpEqfkAq4F43oU5GMgcq6QN0wAMy0h3wX
6QjJk947eIXLZ1rbpH+KHx0ZLiKnKA+eov7GXlpdEMJjc1Hkh72mLWGY7yAE
B4dD+bjuH+tX7tRfXK8Y4IwcyxVTqNE1U0tD31ZJSQixQm7rfvxJEXsD4Sd9
8pFzLMbedvvfk/Lz/PI5U/LS8p7T0vlcbl/ZpIvZN+fPpauEva2yyNdCy95x
J5XRqA9Q5IgzBg9STGWJ55q9KWqR5iEffRr86FVj9DaAWHwj2+hBAjNIvl7i
NgJpSTluIYk3sSNEVAcOyiUvAAoHyZ6TiGq/MwRiUQgozrBuRfLwnhWcqXhL
uDY8zEX9V5vD6qsty4VmeyArBLFOLiaw6967vPTCtQSSMl0g1FQaBH93syNj
FlvqfeWYgWcR1ZGRsfwyfsoeONRl73gXYHF+KfvJxkbjK/pNOBtxW2iY70AS
R0h0bizCZUx0NX+Y5kvr4hXgGCk8qSKn1bDe5Xwl3eL0CUMxUHMod4vj4HZW
LxE+v6ZSoCQQ91yzIX4UVezCfTKJ8lDs6wcO1VqZXIta6ysIZKnXlkVisrat
OAcFDsEy1FoRKVcG/3LLt4Z8k+JzPs+1SmbPb+KuHoYWeUJdJ4zP/ld1UwQL
SHriZHv1UuhRpK8+jeI1XFTPyV+Axe8LLeZEtnijNNr032MO4ab6j5vDkm+n
4jhyxywWCFzcNtBk/ut9pdr3JxyFCasdmYsjxsdUrvgIwq4wED/nSqykqwLp
SjHqq7c72PS2NFLFoGoWQbKUpNbthTdKsKR6+HTba+jY0TvK8KIA1OxDGx/i
jNkpj83JIIMcbS1i69ZHgynTWDoPapEc8MQkUOYrVp2h9/cS0twSONPAryOU
qTbsrqRbQ4V3UzG68005OfC1lGx4aqKl2Q/fIvstlK/8FsEZwZ5JreiUUzvu
2Ttoxrh0cR82SHF8GvrzJmwpKIJ43Pwzl0NXWbFW9m8DCzfoYjJb7GQaQK34
yryGauDldaRacwKW/npS5g24pgpMBv/uLRENYQF/5XxvvBeqAUGvP1pv0nch
d3A4LYw8Qa91tecG1Vjn7+fA1w9aRBm1pjS0LcGhymVe4g9AZG0vc9bTa1QA
v4LX6j0vk7oDh8RuHp8O16LwwUh/hgODEI3CBRtfFJFwqutZfdqVlAqBXm7Q
UmSFOL61uKQPUZLh+n+tuA3wn37628NsmR2oqZLp5+rBe8uCfu4n7I97+/t4
v7rd1KFmS03XfvgOy0QVrciJfHOCJBaqzWEPCSYWMTmH0Ee/Vg6x8EEE5TOd
Fa2X8pjLW2Ihp2TX8PvFhQUx13jgrEMxgi7sVTX//3ysCE3enM4ccgs9IpYK
9e0NWurMU5de2dLHDP/XSBDp7pils9rw8MQA54Vl0aMZ+suM6UXH7lJMc2sC
yhO0gjKbyMNvQXgXvmfHZPpNC05IeQUMM6h+QJwQL1r+LA7qeOnNdby8MZH7
Rr/GtcOt6vT/BpYPGE+9sJAkoGitNJgB4hCdxUpHEVLblwtI3WZyskoaWWV/
0JVFxBL9jzJfMg3wBi9ndI02gT1uCV3l0G0C+PR6+fnzzzvfna5wRRtKAvvG
9eMRL4kMtGc9LDnGPe566rATXOWhSKlNbbMoKueLtiODfLooPPPh5J8x6R76
wKgwf6WZJLFsDMYA0BUXIZu9kkoziqp1nOD6Q05est8WCgvka9yW+Xi+B22P
RGz84URjhWK32QBk3TrkgJNIDy7M1ipM6Zu8KWtdFEwbCi/BiW8xSC1iDqtH
3Ghu4FYfW9qJVJ0osM2PCKbvJK8PI+uXM0Oafw5F14K8XiwYVbU6EKEaM1YS
xuVPZoaSMJUrghjIvajE0lJUsJ1rHYk+3XoF2mhRURpuxqXObwagqMLCfB7o
vyGNC/RM3MguPQbwCWWGQxcBogirmmol1VXOQkqWe+uGu627uTQFEIUr6hKh
3iALt5l9pJyR99lotxm6vbferKoLMJjRc0VnpZbEUCEeh7fWLhMkokCDl6Av
GGUD6IC2rNCEi96wtHN3QZJsXsaxFIxbTrnxFY6x74mt0glXsyWwUYOu3w6h
1NjRmkRzuWvCw9sSADJhqLiiQjqt8Us2ZqyTig9yzjp6tWcQ44dX5JC0y7+M
zOnfyHDXK37Wu4Wk2DSEFj4rMPiTm1ni2LAH21tWwaDUs+qlAyVP5WqHkhrb
1awlPjzJ4zM5oMvMJI5ItdL4klWvZEbvmQ/TdwxIBX+2gO9tjljidilFm67W
VWZZrk5KEqMm3xUEaXj9OrtD8ZSitSGKeQTusrJRm28zFpb9svm3DopPpWQ+
kIsSwPfkzaWK+76oQPly6EJnWKb6B8YCNSeXfuQ3HA7TaXikJgBIkZXNck0I
ZFkXKSMza08eNOrYTsmYLi15IEJGjqHcCQra9TeJ0m+bi9qPcq1Kg6ctxea9
HRogG8vfSj3Y8In4dkNcuV4QlUgZpYLLESquxsH4F6VCOzOAGojZSTIQptbI
av0R+tQ3HgOWvKaL/LEKFDXANJae8I8rNZ49/cY5P55vCXo6pfYsOgzyGtC0
ss0JREKtbZcLqMBNYfGCeA5O4GzcJ7M5HmbTQainLK/hiVLoFMvDnc4fsH2Q
CFBqHQQKPXU54L/eb2/Kudag6bTnaebhwfXDu8uMLi1YqsY7XiwqME260AUE
jHj5vuussR1RmMqA0mKi0/UiIAa2r53HuNeAmlT2MfKdHSbpLBCT59QbE4xR
arEBmJqQeuvs05bNgeF7yvzwiKlB83pJgC1D9KiB4moy+cux94lJdtF9y4IL
iFTBfZkVsKzILGsYDXNdBrbKKDFlK5LYwSAfF+vFk4dVdgZJMKUWoau47WYf
in8eQkXjrbg/Wfve0lzlX4ngtOlawrxIIIow/9IcW/QogjflZQWXqn4Jdao1
/n6cRx/HjC1zeukd7Tcex1YXRExGJnSE7WLOaPzmDqV067pJ2Y64zgGsC+Hq
CqeqnPQTnZrbsLGD/0AQH6dtGbwWxpNOIQpQKiKKF9FDm2EGzvk0B38YBt/A
X6al3OHVF2/D80oLtsVOnzlzWJcFWlVTpS3Iv2SPTvkj2k0vBzhw9h/GT5b+
GgzMpnWrq88CdCScdgZDiLdHGkEbpm6Mg0i15KDIRgp2+80cekDoMJYNxwZm
P3ZAUSKa2NSFrOZcVtKpIjJ4UMBdm28855kQphaRHrNZQHVx3nIH8QGN/W2M
c1S/brc/O8ZzJlhIyrkoAooSGyXq8BfJzt+hIcn+1gg09l7miK2/HVHfLpWh
lTA4470sfin758IVY/OZM5COATqYPRiQN3X+B5GihkHYxGZ8HtD7Kg/6jVUv
0JD4HeDjlpIdRzJaddJqxcFiQXf+6X0660Ct9mBQQPugko45xSpIYaM0nLBM
27pOWaosAo7l9uY6rVJlVeGeoq3baJtgpko5t3M+of8HrwrWSAWiwVr3VMKd
Hms1y3aNW5jU7pxCfYmwD5D7qtmaSURM1E6s2Tjo6WSXuKakCViQTuFGCaTg
NBHEDgjJCWuTK9z1k6+H9mTvY0OMrlUqTUitiwHeoHYm1MhjFIsyLXf2PyM9
D7k6vo3pAQoL8vNjdQBMhZViJf0oTZmTwCgzq6a9pCxtZXE7tSZtrLWgCF+F
bZPhh0m4OFnHGHW4GAc43svlEgvCfusBbu7VAMtYaegAMPHY/Jopm9NCZ8z6
o/eriw1U/SrcJQSNUdquLX3edkLgd6t3Y4SUIkSeFLYuRfouYa3kq5AlFdW/
hwkzRDnY2gBngmOuSzAthgh89/zzccBxIPBMTGH8iQRC5LhaGXnswkyLjyfj
lZLB5KFstAnMEUKELwHUOmaLZGb7uTeg4PggtWvwEdqrpp2v4JbgMqEUaQgi
KklNvx7i6NKWBRdX+BwD1BNXry63cvKehoh7dxNFLia3ujPYiJRzjLcVYzZ0
nc1L2K9UU7FrhNq4nJPznqtW3aYVrD9ERaqcwijjHbnLnnJaqsNO9oONC48Z
uuKfQXuE6b5VfV+tezLlkLzEuPJ2/t18PuUoSoNoS1jFmdBsmGmuLbaqfck/
McAQ7j/OnK97qlXOAdnW/AJaEjmDn7KQGOTwVNmkvXbM5+lPol2zL8b0YS9b
zXNztZ65UcrssaaZnZfTA3vEfKpa+xlpMXL50GsPFyca9bKqRAELzhn99gCR
7he9Bq1+PDGbmV475lRwKBN9NFZ73fKSFtzgAtvau5TCFSO7nrRoJtbErSrq
9vP/pDy0qVnOLrFJZADqowhDLZQmKJUGYlihbuuluNR5c+Rzub7LgP7Lqm6G
4ee/Y3MSo0+J8NPDO6yhhxTXs/Ja6tXgWlEMV6/++dfC5P5LlxbGrNSa4bEY
W/IuSD/OR2Uzk6cBffnQgYgMLunXbZ0v+lrEpXWunWJu5CjC3MZf0a/xqoDP
qHvlArD+ZW4aCHjjYT0Ur63fWKco83vPxEPA60xpKT9qk6FWLrtaUyWdzXPL
j3NzboX94KZOX10LHsQAFuEpKCOBy2dGQzJIs3cf1pQrq8R8HIcQOe2lsvwB
yYUm8cZX0ToXyf4dYkz4beA1CAvLHF/CK3slUubvuec6OwcO+vwWfXTB5A65
lUcHtvZGEKc9J1ecjX5g6P1pXDJLuFVme/Cd84Z28npf69JoQOx/qpjoE5ux
N8xqO4qwCjgfeJXLE/RE3E5WNVP7Q6bRULE0Y+2OILzWfciVimXRKrrQ8MMj
0S+tn60qgL6I0+GFyJ5EURl5+COQ7VAKtzZfHALMNmJSGvCvGTwUMoOTQTWO
0NuBP+m+4HCtSVBXrjdALwEoQCXdCshTQBdFYKxmkExXsx6OybxyfoG2IrPF
MFeco6ygU7201OzpXxA2J11/Kl21ev7/tOE/SrFBi9ls7w5KVrUN4GBhluLG
CruMLKFFkyqQWXsQW1ur8sCVUoRJrc7GBH7ydqygWdIKokgcMVY5VsFU3dJg
Imt8Vnn1Uh0UwJmeB570UxEmKsCMGKlmu30W537J4jNd7q3XAz0aTRqwyzOv
3K0BIiES20Kk8zvo3CDAEGWkDk35c24AuhzewY+cfaepwMigJ3gGjypxKTLk
k9lh74nOc77dXSgG2kqwUY6SJ4VmuXbOYDEZs5AFW5yLfbRxJQdJNGLXWUMd
ITrKo31tomJxZHQg+FG+BEM8XU2FcLfng5/F/wFix0CwKi41/HnW9ThEG53S
KcL+RV2wygpcNnLZFsrz6JXORB02NAwNdXjDnnak/wvm1MS3USfxlZkQMOuB
xZFAyj5b1aQnvS+Rt3nrJOSAHUgYOhaPd6ChsV8ms9TfYv/lIrKbV9BtU5gS
Q/JKxXbByR3rDfX09zpIxEom9lHYz9FcpY0qxPjKVtKiLdgZZmmzYfNg6VOB
e+/eWDJDRYUeDrychtTxXY664nu8ZSubx1R9CU9wZ+QTt+xfcEf4YwCivVv9
5yjJlZk8I2HC/2v4TfJBvNB0TbjzLlL6tH9nJljal+QCqLA27deCocBOhA3h
CGA0xGLalY5x89TZRfSACe3MtleGGJnrpvXD5PPko0eiiv1NXDDXN0fJzFUV
T73ulhClWaewvGySsdcpyPpv4Rty9YPLyLKaDYzD8TK+0ZNBBquKMhySxdoB
cNyOvEbHy7O5yWAHUr2QIvtxNG5RJsyiuln3cPZg69CIUASnxTg0DCkLlFbO
3WQl+ubxyufcPbezitoaOthAmhDhh2Zq4q8zYeUudMK73b2xPmPuEPGyEKEG
g3mMuHA8QHyw9Ko518COdpN3yf6cA3TwAAt19H8rf9uxxIJgo8HItEKyOVTg
4QSNIg7aV+/QMSJQhRPsza3fIYkqAM0zQL7BSbqPUbcDiEU0ejM45OX2Y+Uf
jpag4icSs8w6LbH07KN/Gwbtm3pnTAEDlqlvxuk0ocYbxSOcGsJXB7AW4F40
mf0vJCOSuS71gkScUh1tmdhBL+YKMVdZ/Zs3uvP7l58iyfZj+KM4BF9WGNbC
dG8w+hydqeRXn9i/1V9wRWMpvW2lrJpxSJ7OGgv9hk7PQiHWxZJHFE4vh7Hu
cXOqE3v7BMcWC/iHN6vELa0AjyhHyfMkmG4rsXFY6/Dw05atGxMn24RigfoM
O55C3nkuG2C6nwVZa/y7VcuRAZeNwdAgMnY0NsIzJt83yI8OZVx2Jhji9K9i
2MB/hMw5Fbmrqh95SNiNc+tx2k6NrqAZJQayeCDjnp7fDZcbQpYGHclauvhd
yw/juelBdMYhHi/apznqUsD3M/uRRwJd9uhuo3NdGI0yf4bmHnQN6l1HBcPV
05BdoeylzesIYZSujZQsdRAyLihQ4S4Fhd39Ma899ixApLx5an2XXMYHS9vD
LuuQ77YFt95GJBAGUpkd11Csb1q3To2fG3N2ICg8OFjVc6Wwtc9HYnnUgJ1x
O6pAM0A9zzRXUYoe33DRvSYbUQBKrg+qrAw5UzkvNgiF5JfWaxCnV03JRamJ
8i1w8ApXoKzNLrUsANCPbodWskRp4kPN/k/35DJZvfonaK3QasJPAbU2DtYC
zEPSwHwAzgyeUWsbNXDo7ial5rz3Xc3cY2BiRNxtBLkKsAkj4I5yNp7YV1Rf
gS2QGgDUVqff4CI8agGoBIrK+9bG3MKVNBFKuWDyAS9NkT6vbg8d7jWkcYlG
qrsu45r3iw1czPJvmU283AarO+e68ru2XCh/QLNNEagM3bQGk0OilDjvSdQ+
mrp9VjU15qIcaXV6Uj+euptYr2YAN6Pvdcaqc97r7ao1WIVkpf9jUpRcCu5v
A0JpiTp2KFhSrP4g4vqfaRkGjGRx85utOMczWw+kPmsvknVPyX1UxSbKNiCu
CgSybi8AIcSmBhODd4g3hQYN04SIob/fC9+Ei4coEDQDL4ezVEpLci1EvBUE
QHEo1FmemjBUeKWw3uJ7mSCsWqtJIO1n6E+9vnZacGVk1qMNYHhb0qgQ7/Rj
0AVpnW8CxPaqYrvh/snuUD2b38sJtr0+EYYtqOel7qjyGClgcodTpP+FYcZP
oNWOE7N+iO4OJzW3DOnGwL0YOfUKHAZkqbepIvxccp7OsAclzovn5HNtnnUx
4nqOSdzRGepQ8sx74GGeOSW4/ykyoA+Py8L6cAU4byJT+CxEuP2CUHgVxzvc
qIPk03uB1WjmiKMJ2OYJRge8M7r6crVVcMk6

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5Mpegc4aI+TaSnqUelefM7IJRp4yna0xvypnkZ4efu1essq8cJAfJ688wwcUVymuN9BRJNmu0OHfhoPdP0JRwHGUJ6vEY4kpFUNLdctQ4q4cp4ePOt2BQMzpRBg5KDhDw6E4Qt5+pYmPVhej7UYiF6dGViLrrFhWqe6LivZxDRMw60YVsrB5izqqhBLw4GvpNTlAxA0+jK4SFHD+PaLIbzjxYEOFc7D0OtGm4LjeLy8u271Q1M3KIqlsI55lPJ3OgEwmc5Jk7Jp7Okt8EDR49MfFiW0Y1S71FIELSMg9VpQ5qEP/RS0v/BOsFKNdgP8MwBm0iscdT0eSomnAPqFw9dwWi1eE7IYlJNeeJpHOMPpqVNFYTXM6d4McLKppcDa57Pz7y2WC92SQTioWM0vuevu2oUQVePwaAA70efpsdc4kLWbNpBkt3/715X0i5ZYhwcxAQBkwMKgQLOGSSmWnGdze6G5lCs+7tMjb3ttfqB1ycdOCeB1OIW6jOqS7d0QspTlc4tSOV3YlQpXF4lffdXt/1brzYV9cTy0bOiu6dsuO+1gUc00m/U3bzZzt6aByE5b0stjFnYsg1LkZk6F0KWkohNk6SD5fTPCV8G7WZ5kCEMUtHnMM9EI3DL7RDiqtG1JpTLgpJyZ/mLtkxX/blMW9TbO6gE099ZhHtelhpEahbYWKJBVV9I8u0U32gRZZMejmT1NSh0nvy2XHb7Pu9UqK31Ss0DswoK0SuzBB4YmXtGYtBP4GIH1NH0hOSoXhQdNYxucIyQR5IDow9fkHn1cKDR"
`endif