// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ePyb2ELajdqPo9GnU+hEq407QWwGlcDRDAUfGWdGRJYHEIPlfg5KqmMNjo30
ACvzQdya8mEibg2KKTCR55i0MHncLuF+q1F/3tiTo7YrF+P4nzA5K6KqoTK9
xfNrM4oKsM7siQq23aVGTDNehgWUnxVKEiHuwi8bywqb4NpAcfPMjsoyD6r2
UHWLRxRU+RluOgrFF8mpvqBrYo44lOnfzlRpFoBvcZKdNBtayQpBYTuHStNV
Zcs12b3qj9oqjG+tKpZTGzoYaIWd9slPeeys7asU0wJKdoLKYjGk1BjCg7qW
s1CCT4WRDqe4UoFVpsXSwHbskezLvcPps3DpvXX/7g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
anOWA0RmzsBt1B3k+rA13gbMmye/xjQMaBCS3jgG5fxibX1YJl8wGXUP8MEi
2ZTDYrtL8t/gkXihX8sW/G5TkpLmgi6SOfiIGDdQhwRv7wyapCgZRRfal97+
v8YtTo5OkIqFg5T1ZOzSGdtQ/r3Sbq8yvqy2RPbLdieDfeBkvvZ+3usMNEBq
CV6Kq0xJw0yn6/ydtA5Shec/zJPZQhrnXj4PpLS4JFTXSMaCwZBe8U1l1/29
o9Y2hmT1NGkDve5AAjzx+ooeum/x6Ep4FikZ6E1+UWVdBV+uUX/QwTgHM5SK
fm0bYucby/5heMb9HNSLLM6Q7WGzd54EKPdwkb44EA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eTo+1XuI5CkTrnpQ6TJj6YVlI5JW3tJW38uGwvLraj6xtJKkiPRtOPr20PEW
R9NqeDudc37RZbcwsfPn/ZotOZGeIDpbXitTTElw0sVPbr9Y3KHE6w6HDtTt
xUI2cpG7/dMfoe5g3Y/JQkyNUGBHzWxgOzevRxaSEh5BrIvtYeo2Li8yTEdB
+rVd8wMESY7Wj/UNDZ7QFhEdH3cBkbuPoO/wrbFcPB7ffQkP5gPjgkgwjlsm
L6WUIX4dqjnH8zWVimLONqbZrEctSaDviUyM/dB5Q/fyRpNh8fsdejltj6CR
BW/yV8SKfzNpAJtGIb4VAgXN2N35gk6BJoXM3Nv1RA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QdqnKB5pVSIWpT53aH52UISI1IsD2/nc7LPaAjm3uW6AoLZ7w1d54HhHsUYB
ahsuJ5wch3JTE2X3qik8mvvUeDIpRevVGEQRIHhadfoYvX1dUXPhwo0BlQ8R
2nNO32MaU4m3BefMqT+LcClntoGFNZbtzuOXN2UVi77Leix2zL7TGMWuFs13
WLes5Wecmc4QtHHoIq2cMZVWAqp6EMuNnUFVxuoJngwLk3XS0bvLRAzZ4FdU
SqDdV8AeJi31GbHiTVZL2/oVuDf2QOEmJBxqdVVJG66GYwWmYvqle67DP8pn
q5Z6EslxISWR+aWj2z/eyYjOGhKvzHIlMU7aMFrqKQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
K3mhNfBEErCmOcnl9Maz1Gt424+uLuLqc+TM8V6pVYVbu561B5kTU9NEt9q3
aZ1YEwJp50iZeCJics+I8d2N659i89kup6BS23Ekd72fkTE8q+TjTtVMyF1v
C7b3cGZps3f4w+It7QTRFr2sHl4Im246UX8D4xruoQteUD37+yk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
OkkdnHnMe9RpPoPZ9SetFxr8OZjqgixSTKrH2d3KF6r+F+pB82zeBe+EB3DF
A1VJ/01CzJSoEynD41Sabji59nDSwYXnxcwiwev+XlqT1XODcVnc7ubEvBH5
OJ9ew0pff3H6kRXFHDXv7dvTIfRkzorW6jwgq/VtYSb1KYT4DAxVmai/anRW
Msu7tlZq/W9Knv1Q8MPCymE+Gs6N8ShfKAYsmOG0T1KQZa6H1jgqWJCzZZoN
x5JJzXlJUU7Qihknini4ffOthPgZsQkz+G/bD8smD8Ts+1vfFCXEnPzJjZsM
49sP79JSWS/8KCZk2NUmh0hhO68leHs5izg5P7x3K0Cpn1G7hEczsUeUQWS9
kfpUJ1qzmCOzQgrEVoPLZKMiQk4NWrS1vmnQzy5cg07/HWzIP4iO/qjDIWSj
+5gZl4fR//fVK3Wbm+UWvdecpjMhMkkX1ZtuxDamlZAm0bP8RJrGypAcbY+s
vZvI9uM2XD/PTHBGFwpfnbhSqli5DsAu


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qYZcIqW+KhcWz0sD6iiAPQWukP9kh9sJKXiB9QqBMTw89kdEf0Ign/O/4/bj
/hhcMS5Pz/3KIJs9qrwA26DHPILK81blj1L6CCb5FE3vOBscFa0Pcbboz2rh
VTw9DbfGqhBJEV226Fqb4Lrq9ZImrWhTlMv0uj1B87R4sqKWqmQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tG+8ZJWpv1fwKSHCM1jBnq4B5luhrYdrQjDpV1pbOiiHbB4rR6rbOly33cyP
8m+q/pUZKiivK+Rbdp9IEgbL01v7o/Cil/hJkQwKc3+CcyplBrgCsm6muA+v
lJgafaf2NuFC9p/QOzX9csRAl67RPPRn1aeAVMHw+j+KlJWe8pQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 50208)
`pragma protect data_block
QzK84MqqsVMr2y3U2lWquFefFa6pyE2/Ri9Vwo8FDzMw3MQh7nJZ0/4uLBvF
Op7KOXgE3IGHFUvobSsxWvPeaHfMgTGtfTfh/9Xs+jO+aSU7Z7yZfjNyQI+q
5CwKm3H0oyaJiBX2FzdEvrDS0skuD7ULjjaBDpthovizVlyc8Qj6Q1hiRMdU
OMlItRrJPU5iJm+0es8YCfTYMT5eLL4dAIg7Hjgnbd2O+/SgTAPgKS+9CZqw
rsovZ6nIxJBQD3PXI27RMPwBROeqi2tgcJCreW/+pOUJNXxNQv1/4mJg6dmx
tea5BXwmDxuIDAazAhNadGMEGfV1d9CulBFAMxIb7ieAaUDJsf9wqauvwjeK
1GkOsIOjmSI5QXSJ/vj11Bdn/ifaXuO7UcjQ6H21hmnqheno9wupk0JQQgo5
ebzram+qNN9AMc7UZysdGJFRQBClX4S9f/8hzEROr0mshlCqfL5QtKPBWzx8
2pvMHBqB8LZ2Hu14+VmHiAGwQw7z0k6R2E+alR7+mGXa3YojFIBfbxjF1Mjt
dF8hPxe5GKVihiOd0waLA0I7kjzBMry01fnpSmV1GCBZq5pz3ZvBVeQvKH5d
d9BpsBWzM3lF/dh/4l9khOASNcDeluoEnVsVWRtCPgxQXSR/qC5Q536sZOJ6
Qr3pyJoxXT0JF/M8qXTg/Ah+vgLBZ+lpgDNITg4oqZ2LakJkXDRMdYQx5dh9
ACE8Vb8GGl0OtG8zijd+hNKFQyHQeZeM1BwWp3XHe2zgpkxlH2DjM6juD2sg
x9+fIvyAi/T9kCOlsw3Dw4CGSxdrpY3+dvONsyPqGJ64VoyCxw/iKOzguTff
UAU8VVozsjyAEe9FhxhPtPQp0Hi9prs+zXlNpuPELY/86Mzew4MkPLK/PFYo
q9g4pIZ59v+0I/DeSKk/IsSmu+uK0m8NI/qa57ZjCXiJBSWMaYXW9lUXSLVn
cVwWFOGnN/lgU//58DNNSwlA9KQolZX6e6W2chhgwQ9Omp7CRAQcAbIDoqS7
+KTg68KpkUGx/N3nBKTT/4rsatyDEIxH+4acChqNR7xjTRqyyVWMyrVqftwi
f+XkWvOPkF8YrpxLKpGzAlmSdg/rOG9dnjCHhy3ZRwkTvmWRDoyCgAWfJSQn
7aaIFiPXeCj1HoiZLlw+9nnJG+prneQCjhWS5OZ//FQqghqWMfM6xvRajUXw
zxQJ0g+ikt4cg/vwM7KEPVB5eAxVVIB47ja+Nnyhf0rz75nPJsEpJdn4je1+
e0pwpuWFQee047k2Ige/Hvtf5yBqDp2Qci/rmpT0Rzhxd4aUQCg6CivDyK2p
cRtBY8YH5SoW9zE7BMlahMI4t+EyDQCfOpL41/69tmYybkG4ODr7Lajc+r4e
8Vby1hibDi8bjqE1mDTycjWA8IaMJSGnfBTrEWaMXXZGoetflL5q1NfNzrqA
e1LA9VQnAZpXa3BF2paa2cvjQ4GTO9a0j4Y2pw/nq3vmHmBJp7oTsfDKBSce
1A8mzs3Xo+1nCtjBAnKsxD0HM7Q//vx2o6RsX4/B66k/3EOBZ/ZfHeJ5FQeo
DH0AHYA9e3PBNs4wUruENg/r9eU73MrVNUGaa2IkqMNJEOhFtvOO9Ov2dJKW
CqemL+fJpQC4xI0mP5UJO5Z93db6itGiiTuzjMbFYL43AwAipbelv6NpRd7x
KWIpViMkFDstvXudV0ze/KT8BVsaZMPtCB5rXbagq6YpFd6hlb4CVLd1XzB5
yYhWCMxRG+wsmUovc6eLxQF2/vgaNvy/RJQkqS1LkSPkY1VMe5sChiZte5uV
NHmFzdwYVEfE3351YFe1OksHVWueZhQvYKZZkJKrv9tN/aDb2zjuxnwPnkAb
EDcoAcMtQ/65C40F2miW9/3tJ5N5HFmQATcKvtmmSpGVRtaNOR2kScIfd21q
uMsxDhAFFCp9blseTVZoPfORDmZUXysRmMcqMgevSxmd1kS411wHHcjHvqFO
1rj0tZjr4BRNOs6nLxWpPv+cLQs3PHpJ1Xlw9U/H7SbhbquOQP/S1LnNkunE
ITjtBfcM2JXzLfwi/PEfb354m0Njx2lcEhsgcLRc0f7sbw1nw1M4Z1rSkB84
dFXfAF5YPY4bFkc5L+96IkI54o4bReZ7HXd1HXaMHZteNOMYFEXzRWhJSyvy
5l+ZmZsfjh6FbK4OZAtstrDarV9UKq8iGhDTRo/Xd93lp1IjmK30Rf/rcRnO
B+dIG+Ktfj0sOQxTWSY9ciky8CaPrvXMLUBmMbVRhPU059Nn2scHoOgG5i+b
1jzCJ7lHYGDL2EAQ5I3b/Jt73dRRLuVDFgOCl8gZK6FR3FjZsWcL5yDPHgT3
CRg14auY6K7Q4lxAD0sjee8a6r9zabM7IDP19NZcavsuhzkfC25ZFjsoXSRk
Zdv/5tMKZM7i3UAklr9R+8e0qCbQSOVjP7u3bWcxgzatX63utSEBIM3EgyJj
s4RwsbrvPQBmxSYhtqoa0FDT/S4PdaOmNqqYSKTaZZ2fLf8l8eGB2cy/oXV3
GSWanOIX7fmBk6udNF0TQ9XBZTIN1S8+PpU6hs9iH0prcWGIoQ62D8C6RZZl
t0/CUzVf8jaXDcugXpwY4ULz6+ILAcp8q2IagOKYJC75ZkwDqoIJJYKtyCHr
zgJPHIIuLMuHf79UhvQHpQhRdp3i5kjzxpA5qyaX6pQHFDNkDdqE7YRs0v3n
ZOiIzfxGKXR5hTcpqehQfLmY4ihSkcKqxeROzJw3NZohcm1f+bPngT5kAvS2
4QuiGsdNiFb5YMQ7JhXm/MNsfBhvGdMvIyowtgKZTDb9wa8uZVGmkVEC+2Yz
5f2/OEKgTiaWAht+FnYY+fb/OkJnRH1VVaKB24vVlX690k5oJhdruSAa0etw
6zUVJuJVcRDSLp54LbrnAwHvZdsyqa9Cg7HB0KdN4ZCjyFAWDT/KyqZ2ovEt
9RkOlMYGU9Po7Wml3jhr//g/3HJeXFoaenGRzcOWanQSqX/huskhk74UYvdI
QHo7UUiHda9FgUzlDXXz11FIi0w2FU++SVYOgISKKH+ope60eHMpoegZZP6Q
tcKiYwDRtUpxqF/aIbB4SeDWABenEGOvwiYdZXKTSuAxqkUpD7QxbpybdmSx
ubr9zbaNn2kI+V4SiwQBZiDC2dUg1zoTUOk/XWdjekuJeV+0YXcdYtbzQyn6
eNA/ByqCqCM3nTz+NXHBe3pC/jA6VHV0CSgFyB6577IVrlZzS/VI/CxEs214
MMbvUhCf5h3LVby+S+p0i/y1jZnMyl8Oe3kTKx6oWAKBupUQg292rz5r81rY
5tsnxHfgAiz5uSfQoB9wn7gCbPXIPs2kfHg2HAMx5THlsg/OZZh3I0CQXdjp
dee5+yxSzzSG1CplKsi1LdXXDZbtq8N4ddhuv6lnFRiX2VrdPyshLiFe3aW/
FtTEdrbfWFMHAccazpzBO8kWaGGiyRrGNCilAW4tl3jCsfCXMcQt1ID3ywhO
W+wcYsnGJRsSYbiUJAeP/aToxvLBjxFq+A1dvEH/h1CSGdWaUOBpEJAu1u9N
I0Dc5aTahbouHzOMe9n7BFKI297ZNmK+XL5G0L08gslcbfDNu7aK6ihwyFUp
laZZ4E89NySveOF2ERinRh/xXmH8HgiqVQddzts52/Wy0hcNHprTBOxrEP48
Rs74eQBRPdlqXotFtBJ5zsAbdo+QCyXnx7FlkUeHoJApnqMFkCy5eUhZ+m8D
0jSbXnSWlG6QqDq+DiFVT88j4VQEis9mr4FrJRGcUGL7viTbwgrtoMKUgFlA
hI99R+mKu8AMrq4PSuBTqTGP+b5BLoyX8Rc/eFOrXjcQIWHSwFKHpOlGmUHy
UgcZbWL4CGI5vudVL7KVDAafLLNAJsXyBXzpR4xfIPhYhNFWjU+k5xarr3Om
lY6tKO6cxygQ5Guccpi4g1mqTUDHR2R8kwKKtMTYzDInNRPQ0bLKS/HN8xN6
9gdlkF80ZfpA0KpTQ1Afu5C+N5i/HcFEchmf963J9PP2yEjDlIUMcNranrQf
MQJrkbJ2UF8lDlAOfFKLJL1U/9dMSnKR8E3d5RHcMPVzKLCwg9cKG6+6e5VK
2nc0a4khhg8q2PnLh+2oGUunck05SBkK7f6kcrA5TEu8d+1N3Cp2xISSpJ6c
G66l0R3xlHhWK85iDp7VemoVId+r+c+0Nl84+3C1xHM+yRT3KV8vMKYx7P9z
feU/werPnU/jbr27r5Lm9cLjBPVxLNp080uHb68lGHZ4LHDoygt+AstWUEi5
gzeLKByNaPIjfxtTAajzFKbXJ7Jjau4TalegI3vuru3K9zezXCl0BqCY3Tp/
XmwZl4p5Civ4rgSVbzNHnjy/Vu44tiDmUBEsaM/cv3SAOz+ynFVGDoiL9XDe
4TMDWUZXcb8po2ErIroeLrv/Lgq4izNGjWI4eDsTF9lwNbQs13YHx6mxaSAU
/NwgaklCD030UFfb6i3ECHtrkH3fbQmQaBSwaMxeG08vf5RRLOcmH263GrGJ
Tr5KRzOQvLH7ABTwBUwPKDfMyH/8VHyRN8ljtTj2BuknytmKwm+vYNnQmZk1
FIo6TW+sBN/Z52AegYXeAil54udoT8W4hCdQxyl+VwSt5oToKaaf8InVxeaS
3oL9/NuxFLzg6XnmC+hvHIkRjKwYc2ZAPRQefd7+yviU+aLJbwaIWtMTRHoN
LTMQ8nutynRhHgc5xMyPVgU7yr989KRqMq85SJ+y+t8S1yr3ffwZVMPyx7Be
hbYgEc+6JvyQEmBrHiFTv5vaKUjBFGtu+QC078SVY/nKMICa3qoS+is8muBl
xu/bdPRxrt+iwd3Nmf78Tm0qbT8wFlQjfGxPTZS+BsR486OxNaPukODV2Scr
WZCrEjKXD4K+mqBWJxLChaB7dLh7Xr5KfuX0SnIRH5UQh7l/jkuAUGyOG38u
xBkDVVishiLYJBbTQW5YQuWH3l3YVq9f/eVYdbnOfbUV5Wsv5fKOlzuPRv7x
KIhbHr+nO5Mjuk/JsKsTuRPMqplA5anx8vUNjSjXd1goGvzbdTZb32XYrHz9
3KDRSKJUc/hbQzJKF7RoKcDaJInAFHNtqFI4C7vtNyFqwD9ukHyylesyBH5h
HaurYjC6bZ0F23M5md5fLgcwxulUfAAqcOBiAPBXP795Y45b+wl8ZPGlmplx
CCMX2RcP2/mGnOUDghGAYMBJTyITYDkB7LSjdhEPIheKLGitrkMllYZYkxYB
wgNXX2g/8UrO6UKFjOXAPzfGkEw5l3ZNZTvbOoJj/aJObx2EstJY9IjGjmA/
2nVGOCt6tf0t8Ujb/NXmUDN/bS3KfiaXaQ6q9q29SzxC9GqRjYPcn8vDhPzg
7r6L+TwVLs8bU6RVerlC4HKx9raBpTZiEDhmkdxRNy95C5zfb5MXPLBph9gW
ZCCLHE0ZLCygCTbf/lPZuXEnpD0NXWvJAHkab+6h0S1U1+Vap9JgGWiEp8el
75anzwy9plqprVvSN3FxKU2DlIdul2YWGuepdRfKo/Ufsn2Nrvr/4DBUXV5j
myrAMldX693cK7lWvTK+xClp/w/H/JPYDQopfSJCO8Nw/uBroeIRfW64Ycz+
+780g3q7ulWjRyN9HAGe1GYPUytBUmK/IGii9clVFBpvXlIPI/HxNO6MqdKY
JONCxAbuPr/f5UnMHuUBZvuFFFSwXGlIHpE0suXw3hBEu1RcSKPz2iMq6YnS
zXg2dhGVa7AZiYOt0RyomfFThFgjXGgIoOeqwd74RXLq9qzTLCwmjWLvot0B
PcjmaHXDwhjrI5buqpaovwOMeQmb3AKHGcfPclDUstGi+fjA1QC915XhtTrG
ectyTO8Q+DZ3Z7MvZsreoL3OIvTWrw1i50vM+V8uuzZEr04gGdf9i3KHfzXG
R/+Lir/Uvb6t7zADl+QAo2ENNjY1uZkXsecJXDL45eP++6TlSfsU6B+d/d7K
zbvBSVp8faoBkt012xLMsSjb8O0JTD7jm9ZP16alpnB8d1LHKkvaSYJNSyGQ
63lLLW+0ihJXhcwpP49TlQ2Po9z5wjwJX23n1G0kmOcbboW7QY88JTWGi7WM
PF4919CeTggmesA4812+HZv4BLHEGagbvmzrNzDeoAOUlAgXPSzKPIlpbEah
aoMhFZVelWjzhmuelJn5eP91EimpqyMi70+EIi3YsF+qID1wZjIKwpr+1Uy/
C2xbxVkEJ0uGuIg42PdHuPLwsp5jePY99rLi2zXerHZSsfPv3jAZ6LW/U7hu
qSpJTXo77mLlvPcrIF0dqTqA5Ll0utDkU4W8BUcfjHm0pyl2HBXZwWwXhjS7
aNGY/EShxgHZrfEGnGSSwirKe0TT6X1816oH42efvg5HYiFAS6AGQO23jBrc
hJdPmLoqrhaqjDfXHrCkbQKKNyN+/ej6zoStkR5M4/U/AaABPfC8x7Qsq4yl
XTsf1flL71XsddQGLzKWkfdmJU0cmJFBOIkal6hVUIarAQbVo3qNi/WFIrHD
P7oKs7ySBUWaaniIfWVZL3t0nZteTdGCjiOJ3dxxrlqpeMFWIQSshe9NIfFI
nuVOJ2HBQxOSbsAkss0+6XVFs9p2veRKJY6vUq4jgFSF31poO6C4et/vO+WW
ptZzg1KRtys7lpOhObon1FG1lRxPREetlSr9KVpwBEcIDlZAUvQV/XwxJQ4p
ZblkNFYqb36tbYcX0Q1Pspk7i6e1RkvC6IXUlLEa+l69JuZErJnbZzaXzfk0
dEmupYbiVIghf9UinDqyDqAUnBtUrK1yJYmVXrJ+Be6nRA5LL7mto1jzdp1K
t9V78rsXzz4FN1JiPbMntkrAO/KZNxgOBDzvAgt3bOen3B/xR7FdTVqXekyJ
/DIalLBNfuv+HbbBkf5zpwK7/R3fQUHWvCJmcYSAeNtgvzvm67d04/4jxUti
TnpprN+RmfX5mr4ck5FgEbYL1A76mFeNDXETYCoRcVV2MihnREQD9APFdiSB
EcCVzLSc3RhWlSm+VBvUJG2q3SyRnCPesfadamF/UJLrFQblNhScFn1A7DjO
xkHWdm+qccauYfZ5I1zCB+lKUddp/vcblIb8h16CNIzBUMjrhrDskrR4Cyd2
8T/q94AlYGcImdoa11BdP8w2wJF97WgglQJOoQ9Saa22u8LOXssBTIEMyczC
TLB3m7ek0ZjmPrYgxwQUStjHvnj9akPlVshREa5rN0m2J8nbOzilaWM9Aulg
4PpgIpO3OazG5ZejclL1GCenWx6SUa3uYM1W185ZAdUUJoyEFvgXmxMe3LHN
YBBFAnG+iUkxxsyBpVc3U55hNZ5zwZ8FIskrll3jOy2xuacUL+yh6S+BTvFe
1Lkwo1lmygwdPxwCE2pNITm4HLK9C1AJ5GOWko9l04GJjcgrG50g2IzvQqbN
SgVTsn4y09jLosfrDTaOY7MkyCYkVlnR+cIHGML2AZgP6BzDwt8llLJ5eNHg
Zkldz5q9c/7IBEJPUSr84YXN5bDyd+bDF4Rn3RECt1+uTDH30o7QJHaSBxjq
s76rsQGp3JGVKhJ1bmGXv7t4cMOHde1OHuQiKM2JwFaaI0qQKTNmdds7x4gW
+T1zmCZ0l5r4OytIbWNhr9axu1vA21DvFA3o6Rl7QDKXP5X4TZ0FbJW7VlfM
0pEj2Njqf3iVFDt1gWNJrIXrYziLi/pHEfmE0jpV/tbu2L4lqd2n25BaAVDk
/Wr66EtecVWRtAxCr4OHFpfg1w97PlgBv6drt8LQl1yPP3ajAB0DdGbG0QYY
eVGRZYPcaNAW/j4LUwHwqNuMy4/8KZ9YSyGYicY5xiL5zL/OxGnrdjm6YgcD
5PsMFq8wWmihy953HgRKXypDKClrMh/7iKbOz0yQeK5VPKlGh0ZKwOtg6J9c
gl2HOhY+7+x4rj0bjUsTrvWYurE3YBFPeoaL2+nqrc/0Y4oeK1v2SzMVneM+
1q/biuaxbDcSQgCYndjdmAluDa18GD+0IJX24UGnwoPzX92lfiuAT5IBfXs5
J0QirF8GKa+E2fopzO9zyOoH6VMbW2lkx8sumstJ0TS3und1YTJG5j93LvJI
oXYg0u4NVA+9/4xfXA0UXggn2AOU7o3UXCr07AavC/8ghZ4njmtnSGdPUZ4l
ZR/4r48LTdZI3fvtP3vsWUofusjWowzBKSkHmX0DdRGjt9uCzPcQvuyoVaey
6bJWxfZbQMwx3UVyMFYavGnt8MPgkaV458YuJ7Qsb8mz/Ju8uzhrCGqIQ0wd
gys3CoNh9rJzdBM8hWEj2bjLs4AOH1x+lPXC55L7+Ap75Aawe+strrfOiS3V
mjZvU4s5s+x1a52cJ+bHakswsSPVuKTNZ3oX80e4/fLVuljyNYBR+rg6iyOV
Sx7BVvu6cPz9nqLab83FoReraCheQODZ7/E6Bjsa3bnA8I0Asqvgg0Q7f+er
ozabd0QyVSNZ1odJRH0B8eR+/cbAOSrxWk/xo0CLgXYms9lTanFZo9scExE0
RKLsX6ezTHIg1eWCTiwlyVMiIb5FA6bkRoW9C5De0MInmzA45LC93t06sEcL
nTKJch+hS2o97EA25eQ41I+WVic5H/gonBHCUlBL5VwMZuodmCMeV+asWZQx
p81rijbuTK78Ggx2Lal5hJfHrglWz+c7ugCZ92lDA7hnEY5xk3o3hxClTyb7
oBw58C/S7TdiuDJLpsXYqNplm9Nk2KMgGSsgiz0Q4ICyD/Y7dB9BrUzf1+yx
LVwwh71ARAXOyIp5kLgMs+zbjTG1uAKgbKrU3uWP3dvaQe7gv5J60kswWJvx
kfHJpFF0GI4NuQLPNw9OyL7cqhFWw98rkpWv3oTVf5IcZRXUQdplkGseJ7HJ
kDHoHYPInY5oy/vugwoA7nO4eeBIxNZ7I++7twN3WSZCqMx3FkKVMPteGoDD
IzHBpdab6kfANgB8ocOqjl68G+OGsvFd9gUhePOK4eJczUGZ6Wa8dLZoNXOa
B2DY9BKd52Ag+4GqswQhALU0yXxExe6fZKo0UzAeAlNIr56XJUCCucSu98ms
nVLxh2Mr4VVd1K+M0v5sWNb9kj+1DJC9GKNx3jbXa/hDvirLdqJjjjDDX/g8
QNN8AnvCbhE9LB9Y8OKWTUL7TLJngeT3DgUPb2s9sjjbcL0BQjnH6WDmj3Ug
5khDcVJkMSy5sN0W2plOnVgP781iFjahnKLUlzMTRMAOaWA/cHYHI9xcw3G8
0+ewa5yIYxlHYs09k5FHxEDSleeheLxkGzXPY/+Fqql+mzD/OKxztwvW6Y8d
mNkrkTC20A0VHZK89qJbYiGR8n44o681OQVmpkZ2j5G8jUnqSFeI560NNnp4
fieUGyEK/9OTqI55/DQvzvXel8QIStTS6I5u4v6Bw2/vmfJoTME9mAzSY7RR
SSCQJIBaUyLRwSfB811iejbmg3s4D4LPnWTns+66n5ELZr28s38hiDwTyx+v
7IiBTtcxgM+ne486rkY2u8V5uzwNoQN78zd1pUzz1glHyT0PrNk231FMdacI
BC9QhuT3dHd/H+Hh+qmMeL3aznI6LQ4TjvsWY/NyFZnfByDayV48vTnxvz37
TVPFRzDQTdB6jVdADgiur7axTh36H6EHI3aBwB3mdLBc1xmFHtf/d/Z2ck/p
dapB6nY4JgydKoyHKNwlSXGFH2a2+fw+y/+xJ0M8Qow90TxyOt80z5kBgYhd
DKW2rJR+bFSUR7apIHDYyIb4UkMzWoHeWezsooSG+d9B9X/cDZuJU3GVEFO1
bSmEVqrMuWyV5R211L5ef2n9sP4MLWAzkysNYw2d8x8zVujyAeiDBE5OR7ps
ajNP5/fnkAxOTp69fWvv9j/DWuamSYX4zXb/WVV22IhfX7XpElma1Gq8TNCL
XDgDcjNLDjJgZ+CDOn1xia4CGf1n2NyWXIVs2IQpFEslYvcZlSBNSY6YEsGo
vzoOwI98GnXmvnoiIsOQhIZPrfA+cLSNH4R78oJ9Hl8XLFYv5qHfsdri3sTm
e73OmeqNCUaHlPMc1siU+/LULMXiH5hfEpCPfJiY3crsqe2aUjgQcykdF6+T
jL4bTjNJij9/3Ps8+sovMzJK1gv0lSckIa0P+L14c+Y2ZH89jkKJ2VlBpv5z
cboeoR8t++DM9IcQqCihJa8U5gtWzyHkhA2AqpOKJLEH33bvkQVin0FE3RP3
4r+gbNoFYEzpf8w+zfX2X5H3m2p87ZaYVZDR1FwdHhG16US2Ant6GQ64qZa0
KcmxDPJlCfG20pEkh42N/gCIPwZ5c6au3b7Uxlzo61CfORCihhzyBcH/eh06
MD1hyJtNPpEIPZ6ztdZZrfb5l9d0YiJ4+euF86HCT273fVYDETldvwiUZhDy
qfwwcF3LW9tIDCiDzOiNLt19DIyKERaOfRj7MtrNDSAVqqoNreBC/1d2IbYz
Ay6FfUp/EuXkSec0ccRDuIV4b34YkJ1t7A4Jtsz5rp8rG+PtYGBZhy0w1XDg
tp2OY5TC4gsaglcHsI2YBQLTPtoVR0NByxtxB4RuodyMLOJlaKYWMkCR1VPY
+Te9qzPaMum+YDNZOz/eOadmJwx72mWvTyanWBtcvYBwmP4/vr7TPy6+Vkhg
Gxy1oj80l8Hdtmdgb1kOABdSFvjUBEdASbWmeNZzl0Dj/veEVyR7+pmax833
aeDs2SvptbNFdRpsQXw1nmkqQ7QH4FkjLEYkcp5KFJDw2OFlN7t0Bni4oEjh
CnAlwS6vGgERaJtaZkKDFcHU1MdWXtiF1UmxqBmKe1AnkirrK3ZNBcb5PjZ6
BnFFttq1qUzRlvRmN94NgcYJau1v9u7TVTxCIJ7XQBuybSCJB+9rD2or0tXQ
DLD0nIoREug7qEAF9Hs+BjnJaYv9SAdI4VsLyLWKQO411NwQH51Y1XrYLxUw
fQ7a1ImxO40A+vQ147PGG45bKBk9bfp/bC51qx0Buu8NyA1XZ1+4YlBbFwX2
7/Mv5WmRh5xRy1FMSRQrYnm7U3nFb9ljuMU6h9UNGPufPxcaAoOBCdvBGw4E
rgKpNXwAZlUR3qTrZ/ZvLI4vHs6SD7QXeCfU0XrNlz/VyQWPWvC45H7Setk9
766teaQbQM1dhHPJ64WLZP4J64idbNcSdpXXagD3OEk2M9mRdNx4uGOgxXIY
lAcSSzmVHSLiWJPsh6eeH1MZS3YDlV/AqCNq5nUBsqn+BHdUedy4fT6sqb9v
K/We7rzscII+QukZJ2qGO9TrKKPAE9QCsAY9D3c3gti9wg+N8cPSabmZ3qU8
ty39jw/busMxmz/Exh6ZPJTNrBG2ZRNURocJXnO0bVafOz2UtEd3ItpxpPIF
iYeKU0goZDYC//t++HRwkpy8jRLwfXxZDaEclYr3MvnTG6WdXD1ggf7h70x5
vuesI8InRqAl/CukzT5IZgouRJME4K0ajoRqZvI5039Z8DDqUqaN+8HER2vR
Mkwi4a9qYA/VwgwfdZ8i1gZdmwUpUEJrssZLZsAqO6/1AiwGo+VDxCHvGHzC
CpoqTAIYuB16QhNCl6PM4s5loYGGW6YxT0wwR39WlL9HPeZGTOKrJsxE9jQs
mf3/BWCA1LKs2vVbgNNV60a4qDN6IoFqi4FccvaQJpycb4wfu5Ebvj6md+I4
HDpo8pZo70W30JnutStMVVhrQwwrMvec0GrrfQMTCW9nRVbLg0uoJ5VWyObT
AMi4Gq+VYG0p2N4g7DSbYWKAxLQWys3wPJykWSNVWB+M7UEwQP46g31jGuNR
2193IIEJM5Av9GqM6+qoVErz5FboijUYXpix+BH+GFXHo+car09r5dsxSjNR
I6hnAYGdVJoIuC5xpRkVdza8lv0/Kc4QxLvxNCs8u0VMkGY9KDHJIiQvR+gl
8HfLeZG2LQ7txorgU4/OKrvDRDFv31C0C2D9yasN53Zvi+z1VBSU88XOKZ15
KSNo+dkQm91nInLMYK06lDw6b9nL2GmGW2/qE45CJU5Tho8t44oJDOPb2/Dw
LMrvqYVlIHKqvZZlMHVtiO+zNrJSiuNDfDrAO1PyGda7Ty34dFcf6XXV3jZI
FqFwstyWUgeQiVOb/Mp5QkPBYwBh98fAo5DZPKLIh1CB7mXo5NTxCI9jPM07
oxax/2HkVOuMu+hsTAp4WGPD5K+SUNtTucVt4KCBS+8uHNuRqu0qtHZcGnvq
ZaGba0OK1Q+GT780r3ZEIuMlbOSROi4BJQ6/T79eBSKjNzoyP51teU87b9ll
Lr0YQ59eWJb8jefNM4igPRyjNNy0cNe79BVMSNk6fcN68YZ277buMP0T6j8R
Ei4Kt/Uv+GhgjvOoMFfTpOsdC6hVa0zkgOdlh0TUPL6yo40S8fWitlNlD4f5
12SeDLwLEgPRRitomuVA9zA0lEXXR4q2oBQeNxR6TMBiBkg0/yzDzSwkWmWx
wUnIyIvmz4+RkEA6hk81qzVWNLreMayEVWiRmiaZP1RnFWokskcDVFp1k3M1
iicJg1WU2PhoTP8zyuUBiK7X/MACncQ+RJNsTejqya3O73bRBqS2O0VIkymx
X6j/0Hf0LdbSG/THOJ9F8A7sRSoKQKW5fhozl2bzl5aLaqxrGbdLBUyYCyXh
A02ae9AUEJz10y/kh6+SOANs6cMW2gu5lb3npinsSkvztzbIFloaxaRCQmc1
+UQwA7laTU1jnOPNFtc2oXM/ZLg7pODj+N+Qd5b0slZWbaNSZ+0wNLtXfnQ5
yS/YrPNkRJUb8r5NQ/oJWZgt0WR+io25FbMKZNtrC3TcILI8oXuFyEgrFMBs
PYvJymHg4eQ96xgfW/UzDz+7NjVKx3Hrw2hVhcc/99PDeIZhHJIBmGG9vfFs
NCxsm/4A9iWUSJVNYhxzMiTSUy0DdFYDCsuAmkpF+q6zipYYX3kzNGnm3+U8
dQ9CvL/KSdlUa5fRxq9y5YFLp4uK/M/xMBsQNl0GAqgFyYxCxCAnYv+52Lee
/wgR0i9u1cPYvM/8BKXmdkhbbYo5SkOJdbO73dWVKBuP9wnctaJffgch/M9q
SPAKPirSQtALF0RmYgXRp2djzlQZEgJH1+cBIY4FigyA6IAsC5Bcsz4SQq2V
wNjoiXBLYUlQ+5rvlFgyjTZGuFQ/mKsU5aT4qsVKtKV4HFJpug3GbbK/gPNs
GSJEm98O9Z1Ut0C9ufQrDbLYLP2Gf8iimMULAx0wXyqZ2YKsNIVQWULmjigI
Hgw5PVNOdKabRQPCsBV2Yjfn4oIE0EA2OApf/3hwnaPckNblTMrTNA3MWUD1
sMYjEMdvsVTvMeJr2DQOIEHpgu1JH9YKbszXs98sn3Xt3uKDKn/czPMj5eKU
clQKRhjdUVPVOC/hJAa3vQJfCrtcU8emVwQsPMEdAMmiT+W5C4BrbIPOU/Kj
nPGjJ8x4aZuuO028/CMVtBXZyNnrsduJ9TaKpKlVoyBjh7VW2Z3tC6GCh/pn
+6Cb51efXjQHEH43fV7MgeSDLG0WvXqkjbzjsodfWdx9p+LHaRDRUC/Q1Cwz
khlJNUraRBo5eMWYrrypksciirP9zSySaj7yl7DgksawtB9MlNoSRE0+QMZE
OTaoqETac1nzE0ycnoLtVYaO2zlzgGdQ8kWpeZp9uD0iAGcIyp5CzSZ5xZ10
bcu6rP90wIkLfR6Akw3rsIFiZ9WbbhkW8CZfl/kKW8+qonl+PblRxJ327D6K
3cGf1t84O2xSRSi+nR8vUMlmJs9D3CV/FE0lubwpA7Gr4A9cBaJV0fFQuUV8
UAAUWCvZaCwACA4EAFeQvuQONc+PW61Za3PoXJvz1ze3FTYQ/VNLepd+JCQM
3xcso5OBWd+04lEuXPAXbCkPtYqKp2CF/ctXCtC4Fhs00uiN6825Niv9M8m9
22qYEjmagjVl1dZ350TCB1ahybL33vBpbHErZDQAsUqF9nnzNJHlUGRZVY3E
vwsuvwyU8HMtdXQAbEIzqzvKTcgNg6nG69FtsiH7B/1y9aOSdM8SFpuL3B9B
sjDZSEOld1r/lHM08lsyy2yF6m0yDvDS4oTs61cUPPwKq3rJwgquXSFCyS2W
2cbz6c9dTazpO35Q1kYXvm8ZZFjvl461uk83c/ASyfkgBidsFCddzhb0tWO3
fANkHMPL1iihpl9hXBKXSc5/2Q8xelsaEqkoWjYHBDYIxtJkjin+cqrJdL78
SR2zAaKFps+IsqkAivyZE+hb5kM5QJ88ZjNWg5fk/aM6n2XlC6i6ihl3exVj
sFHl3oJ3gA7wJtVsQ8tBfxOcjOiLpWew8KNlwo8ZT/8xdcwnDKrFI7UoeEFD
S+rnPdWJojHGb3Zn2M1KECkjNhXBygtG87u8cG9ubk3iKNrmiwHPc23a4/9u
R9HE7IYVyiPo4UftwkVQR9Uok8QF2MM/gfCA5In4T9tX8aDH6/CERyKVCVWM
8KjaTW/Sxi8304Fqk+Eh2C/kA1tXTrbfwUJCtMjEUulluz0u653jcUGnNAWZ
Qah7Tc72VacBHEMfH0yds21q5Q6UI5+92BZD4fkmtYXjKcwBqxpGnLL7Pz8l
CadkFDVb+EIYdPhH8HjSoK2PMN9/qIV7NNP5uqYRAmKDpnx5lONcet2wzgr8
IJnFXF3pM5t/Svgg2TZcMsCgzgU3gCmGdOaXN9hDLT69NzHHoLO1nVigWOLa
da8ax2f7toUTpje+NFJsF45Ni2lu8lkWL2GUiRQBUCUxHc9xkI0UZDr7upmz
za+XJM3Fc2Cv+oyD79l8C+K25R90GlF65APkmrU4VgUMqaOL2tOHw0yrcmEc
CRnNL5ZHec4gJuFHI6ZnZet8sliJTsIX8ID0e+1OZGbWqYEv7jjHwHapUQup
ITBvzB22H0BHnoBWwz1D1xq/UpxBYb/I3XJKpmZK6X3ThKAeFOmx7K6s7Ec/
f1AhYo1FP2E/FvkypFvoHEy0pTfyXfRzELYXprRx8Zl5fy7nOO/+qlhei1IQ
WhdtEpxwq7/zPDMyidmwiJIcpeWCRr+hzD5dIDhEuXfeLGIPJQvvFq5fxyM/
EvIO8mn+CYBCK8hyUUxEhskVtsjX9SQokrvlfU26BGE3wRnEFEUpMHPaDiW9
dHwQFs4PRbdWKtVNw61GdOnYlJCjx/VrWPkz+LzqEnbWAYXY/TYk6N++ia1Q
E+w3isGXzQdM0R8FijZyMIBpufqjPj3MTk5XUJyup/arHk0QGeVhut66fNF+
or0+paUvcww0Y3ow9hFQQ6qxbEKqmAc2PmH4c2pTOJxgMcnlKNca0KGpY+K4
g5QBj7aRvv5emWXUxBRL+PJ1J33pi/lZVf1cOHeLXCnc6Ty5gXH3SvFLJOCD
AvLtdV/+fITSIzf6IAf8MlHPdvE2d6Qem8++f1qNzWf8bOD1TuKQ+0WInaUQ
NJaN3xkHGfnD5XgCoPrJUetOHrSAaDijrOLKHtgECUUdPgSeqhF3usUgAK7o
AXPBFgqOWVGnRjdB6GnMNNm6z5KI9Tdayfi/8Xf4PXpFXdBUroy8oxVKIiJY
0vB7+fX2X1v9xDw/AULO5CkLGr1MGo6DJSRDYVfa8MXWDrKQhpdOEQFfyDDP
aKcTIikdbSzumfgLosrNuFOO6vforFsSxrNY14H6IJiasVJCUhKfxCKzDwAr
SAwwMzIeUhltbv+HJYua/KN8JooTw0ZaeJqu4MUt9pP392kLHhcor9OsM2aA
wRaxpu0ISqQImYen6KjgCWpBSotxO+K9yyMQy6oUrypgg1vONOsP5Ebd1EUJ
RH/KNX6gwvhHwrUlsvZUHS2PJwjMVVy7CfL/OgpJjQJM97nVkB5C+xJ3c8Zw
3AHgKOrNbY/T+AmRANCiow5pQDsC7yfiGRTbpmqq3O7oU8wj2DPjrk0UEmu4
dUfMCWImgkQdpUmL36fmuwGESqkKVMzgPe9s9VhOVatcLDR7F4hiS5A+mVSd
i1I/Iho/WyH3pD6qvtYlEsbWdVvVe6+g9fJuOCoeCY2x3ptgTxHSpb8MxgPo
zmwkhi1FDtHIIATGEt161h4lRHFpxGg+bMp95vXuHZsAfEJwUjyzSt7hmJRd
P82UCe9pnB87XkDiVcHwRME+95nRgUX4vMuxbhc05sfArY5ou8iBZR6UaQOx
qmkgCe83CyjGzvrLUByPblKjNMJBokleZs+SkQPJ4XBg9cl/eCziqzWDz2Oa
phSHnbauKaRx5Nu3mlXnt5yb0EOz53Pe3G8wAYjjYSdS+gg11J2ucoeexnKI
hlsfqRv3VTP8EDyJ3mT+z4l6iDxr0PRqp3JUGrbcoiofHqH+dlK1feStR21/
ZUV7j2fRXMVdfcBfB+TZ7aog9tVm6OIX8aGCrBL4d/WZGmuxAatY0lZHxRKt
B9l7WjLBxSHZfFpzejLyfthxuNqYzhTNT8vD7W6wrKH9pnEPCfuz2+/dWoJ/
LvrC24MQNJQAqGMtaloKczSRjlgTBcsdtYg4e+1MDNuxx5Gp4gUL9sKg1aVh
2Pdjq2BegEOwHxuUOLj3DVOn6fLgxVl+cF1Iq6pcOpyEhuJNoq1FurmUWkQl
krZCkxg2mUzRWk9QoFVeBBPOb/UJSI2crTMhGi0IwXWbdJz1I5atBOJBfaX9
obbq4IQtEwOPsglwWeJvwowMjr+r87/vARXWfEgmdb35ncVA3nj8739QwmUQ
6/x4S5Gq8o7enWweDe0qGNn8qgDnR96lk2+RW2uwVXFh7n1yrzpOpb11CO5p
BPmq8yhl361TIZg6gtzzEL3Xr54WbH13QhE3GwOvEWuM1gvhXV1RD5Q0wCf4
Md+1UGARcJ6LAyxBIUJ/KmPJrsLCWCcDawS0GM5Zo52OTWNSQ0JzDUtX5wzJ
dUPQNCRiQoIsYUmQOKwIl6Ha5lriyn0XAsCJ9Ma1ERpKlvke5YWWvMMmQJHM
8kETSNTyqocwkX96vKTASeYtYruLkQgJNfIIlm5zW+HQHYlb1ay7jt8yI9oz
EW+rj1egZy8j6ImK3qp5OX5pI4Blc1QidUyXNGyWu8RJuRmXVBksu8nTFSdZ
MVaxO1RVxqXhlediMZ1vSYqLR7ovTveqtGIPayFseWELfJLJ5FPY1sOwgckY
Qv40Z7tI46sNMM0atmVsg8JYeiHZZwjOfywocQaj3eoVU3NaPLCJXlfKFQX2
szGikan7FJU7CGGENJqKYYAP4w1v317FGNgPcDJjkP6zJ/zGdBvueeoDOZ1/
vtko2F8GDB1TvWOiP8nJN6aP24ag9Sw54EiW+I0ZkKuCe4obP3aWAkN4n2Ec
+EY0dyNSOHwc11MxzopHTqEgqanET9Bet0mclQnnX8J+6orN8tyUOVN1tSkV
DCBnVdTXM66ckyKhipSye90eFxXpgDUashr3jxrnsxjWz5nrucM/gvL5lk/P
9r6wzlV/415UelyHUqY9x+7JXRSjbT0XK2hDx0qQCYgDbAPkuRUepEROKqrR
1A0dCGxhdmNO7x3927miP4h7z9kTFXFVIbsmDYrSW4H93YoCTIRGeVsxV+/U
J/XMdlcNrb4kszjKPMIW4RE2rFbMMJn7wzHg8rgdw3JwiTBpQ4tGPyL++uiL
hPKLnJu+5EBtlgS6Ngmtwen50dZhqxkEPNNcXq7XxCHVtN/CTuMVzb4yASp/
3Junm9/iH2+R4tCZQz5fDteNCUg7g1KPBv6rcZa2wWb4rgj09Q4iajTkeQlt
/+HgRgVY6L1qS+L5br43Nl7U6Pt95OQqaZ8C6t3ZgorLP8Atvw186fQP/dWe
fj8+XUz8eIXVU9ISrByn2dq/uJDoVLL+wBTtckX3GyO/tnZ05FGuqPZNbfKo
y1ZZhudXmNnH3BsF8+k3m1kO1Fej9Lz99MaJFiCc5Adc5r8q27M5Q6PSgOiX
AhpSfpgNH6qmB3V2UWvYo5KRxCx8hBHgXJjIbJDdy8XgxvkR2yxc7D76BQNS
588odzaCGMpzBBJiPJcuciDX3K5j9VrtDTL71YEOH6FxQRtb/s/srArMWPF2
yoMoP4436P/1G1ewjgKcessAQgwBB3BhviSL6asgU/XwqRsxkY8tFABlhP28
8kEOJuTbCJWYU4TIgZwwByujPQhl39N+olgRqGxrvGIESW+fw8COlqQSfKey
pAiHxw/UcWA6+BwHM/B75ZARo52sU4PZaPGUM1rrIFvwbqrtlJcvYGeuS0FE
Nj371xZSD+g8IWJAJkYyWY+SSAD1mO5E5VBG+BUpU0fqcegK3gT0qjb3CDWZ
OIAatY2PaOALIpcJTpjthn0Gw3xdTgpeGhDI5C/WXD3aH1GbKBIZy2ame9CD
65LjDmME73O+yYQfQ7PaLBwFdI4lPiYN+C3jYheYuwGYsh9wSR+69AjUgboQ
GwxHGWoew95wWWbWxxODDy4mdiD2ynV1oJgwGJejcEXF/c/NiovGtvJro8hI
pH4U8KxjEB/6EVC3Ip6DHSUoFXbcY7iDVVcgCa43ANzjORQtxNnCbi130F0T
wOZjzC8UjqILuII2gzS5iuqoxTgf7Iw/sJe4DXWAN42nLRK6qzR7QUAARGTp
S/kIHYhGXMPwOo9FSUOgjmWQmdBJNEGhR7kl+rhftirDfnD3LTZII0gbCTZU
J7pvmKklgdSSyfNMEBSMXwsrpsk2MVMjqThVfOuiheJelNsKtJ6P6lZsmih8
WgM8ag2HyR3NsAFcICfqDqxAFtiMaokP5JaUijX6J6/iGNEEpUYmkEfvFMDH
SH7c0/GxU7gyY4gmmKanvjNw+AHIzBsGRpWZgb3ARmqqN+8T/lkD/QX9WzrK
L0JPNMtOXdiwt/O/6Mun1Xaypzo9/wHLlvyY/y+3QruCouefAKGjN6rlaAIv
YJRDSQhzHMyBcZGFDdgGTktfK2RgeUNFbrrN9Tf1mjLbCPyMVmbBe7ARpwc+
JUUmg3CyVSbQXiu4+51qK2oUt41Ev10GSgbkuBaZfMLmugXR31jpCokMToI4
obfMX83ckcs7e41YYIrRxJolBisrj2osLYlabFMAQfEETB8IjlTEIzdANeRf
/NyxGOlns5pcnTuFDn6N4X4lAcN+9lk7LlECKg7QvJw+EdaVD6n3LNCS73tC
sI3uornM+z6vNcui8O3gS4ExDw/BaMMisPPiI5hod9CCZY6AwOxi4OzvWdg/
97j21MeBfw9MhueRVKxbAfIkatv9oylyasPRmWD6w5NH0kJ4uwEIt6gnX0ih
BGBRxoDFRJlEJiZC2nPv5XtvSAiheEQ4G89Guz7KfDBXECYh8/EduWitPXIG
ib7ipXgYdghoO+jxLC+o/mI7Or2y5s/ACnsrGjyIsTm2TpoGVKe9QzvwH2g0
7nScTkiz6KCwGpoWQrU83z86i69T7dA97cJ7GaRPEgNFKFaO23zkawTak9Py
hWI9GsuhSunD4mMeDIh+vWJAt+zdYUCYyxqby3CaIv7LrU8gxbmCSkLqS/WE
A6hNYTQdvHSnNtavey1yJj6qNBp1xNiZbx1d+zQiQqZGDHR0RxhIFgLrdjq5
JO6WEvvulMLdVGyMRIOdNOmcxBcmask7kq0Y7ZRMtnrY4ryapQcupq2zHL4a
4z2Y4dQPjqqbBGDMMOFnCSVyThrmcMGPRFIv7wRAdGk8cWWA5SrKzluP400h
ULHeNMUhelTkPgD26WJow6eARdNFp0G2HE1NO78bZ0CkswnOo+9gzwJl3RLF
6CPZib6ArtvLJDWdcom99pD2LBPI0obFbaNhjmCTTNbXiyxZYSu11ABYZNYe
bWes5LfTvdNCK59x/sPMfDy0bH61z15zEjjkBILRnpLiYAfkywrhdjqW0SOv
+FhBfsH9SoLGZrsTod265qma+7YUwRKPkqlFLsOf8uJHOZ5kiRSBNZDF8prr
yYes0REN0PLVzpOLx8tLLV4S8BBuLaP36SullR2rFrFAzRY58MBX2k9KBoxS
egEpsLTouheRMZ9BXqnCXQHlkY7VxXovS1al7s+YUX/AuTuSmUo0quPFKCE3
ZCt0y8kHrVhxNeoUVk4FQkQforgWomDNpPROG+y0the8uerOanzcxYHhQbqR
2FGmOxuAsBqY/jK+3yKcqAtE1cXi26D8BNZqayqYXarQHyw/x2+cKq5+cGex
6H/cYlXmfLfPW5tu8oYALsYJ7hL1TQD67opsiHe83ocGmKNv+RPS4ftRaWVt
oj5xaBaPhL2aY62KQ+WUEFisG8Ln7tJATE85HWO6p9EXhTifjDb8uLwu/qTi
cwvR3932jxtWLjZwyk4fR0GIIgAdHZpHfhEX+QcFSwLGssEFu6DL4s6GAkRD
20BiN8xeaWyMex0BxJl/Aa6pwqqIXWkKVWhsv0ZSl5x4wq/qI3C+QECVxtKm
3z2FRfF3Mwf6joUKwA/3OiCwi1SRgQLNJ7jYA1Lmh2yGcKUTQUj3EFiNIH3R
b6JQtx0JVG0c3wg1QbnuUcLNo0Tbp+yQvPygKYVd/Yr1EhUZDsj2Zv8w1fEP
1y1KbgWHcC2tC/ZAe4oSIcUDEDabcQSbZeZ9b5jXa9Me6JeLYpMoZ7GkAZhL
YEdELIe4bWnplOy1qqvdfzTryGVY5eC7BYphPAd7vr0cFbVxRRYyxQ0aoFq8
SnX+Xmqn4GCMIliXRUtZA5mOHz5V2Xcz0CNkb5lT4V1fAADjMy8jHLf/S2BR
0qHAUVY/iBd/pZzcRyr6JJv5TURiefi73vLyqbVwjxqbWsVLtarizGQozpjs
Cz/BOPBM8HAGF6BKKYDhWvmdGt2GfU/s8LJGAp+ez929BKWaU1Gbq23vNsyY
sl7tNZ5Sr6RBGELibrknboy0YHltuiUeKuBFw96Db7mUpHEkgESCPiyIxtYe
fn1+d6d+xRJRw7A18m7/jKNQC+0G89P4LMhbcSUq9+ZZpRM3ujzl9KFGZRaz
BMNrS3Kr0IShDznmaMmiAuDRiiCo944uWQgClAEnGI9FjoXu/DcHS1Hl0SXd
Oi5RxOEv0+T5TVE3Mxq2tZ96omxXkrwE/xTurpQIlS4Y3vacoBxu34DOtMBj
Ikt6M0YHfcXlj+zzqDpFjQ2b32wyd8YDBzObj7BCHi/G3m/Iv+8XVIGF7BY9
rFdqWBMltbJ0o1g9G+/geOj8LjyBAo8az6di7mUyywig3haRDSrcYr8TBD6r
RRRiVvbkotka3IMV++B8udv0wkpO4AUcJ+xZbyCYibaXcPQW1XILtAnASgbL
tk2T4uWVWBwTKpL5I9sSiAIsPp2lALj80c0ryqCR7/afpbiWFgzQchCGrsnB
xrhTYL0dLZVBnUD7rZW6phld/j9iGBQbzbuV4Uf5BsLJ0745rGqbmFAU2XIN
IKX+AxUM6gXnKJN6kXWWCySLiboyTOCzbMehorco0jqzhZrFihVqCv2mMl/1
2M90nzFk7KS2NCiQuVrZFR4SU+k1+NsE1ByLFoDIzGtEm9cDmlZC0SnLTSTt
OmJFQ2Nj+HttUITY9znumXE3a1iMumWbMb8zU3BHEcwU8jEQT8i/vbK6qur9
AUVh4FoP2eVweHefVNQZ3F8RYP5DJi5pvTCgwS5DnjYiy4N/eY0mBVWwMJM7
dDS1iDMJ/69pFXI3NFjA2Zy9QUo2/yqBnsh9HlgjPENnBF+udWvwbgBjgVcE
z/Sy+RcYK/uqMT3sQjRcpC2htOyCA/mL/geLIiixhAAmiC9hqBt0z+uXPUyN
HAoQZSE9g3ZWpLE1lqj8ZDc4xuotYUWY4lTqBq6iQipdL0c3u8znwaCNgS3k
ch2f3WB3ejC7XO8+K9gaT8LM3bWN+JiYvQ+beyfNQgmGVMCo0167auKcipzh
grPO/ISPkIUZc4/9/ppNJDgPH+LWqTp04k/Y0Tfg/MfY/giRREUBpPa8Cm+9
W9GWWVzNL5BAR6PhfakrCNsaB8o8n4BCIVgmHBMtybocQ8VNcoEdn3Ozdc1h
HPn5daYOk+S1AL16OiOSxDWyKMou6gFl0xE8Lj9WfqaLRr+jy2A2+4kUVsnf
EniW2ak9TufUtTmJhq9MVOjaGmQOS1kjbPlHuUz16pYCQHPb2oJDo1i5sjoN
5SlL/SXiwi1i93QkqvqoOisy8rWOyNDSCNG9Bj2kAje/nUbFy9pZWtmYHr6Z
RQLWos7UFM1fodWaC19Z+wsVpeJWp4JyBkMgZFAmnv1YyY+kenfLGIdcjpe1
2kd3yjdxooy8DaXM2Oi1ZLjnkGOVxJAeYvAGVUYS03Ecq/zGTv9XdudSPgjd
6TeBytRcluENRj5+LRXxDV4ksrMCoHmuXRGfULmeqfYZRyhdz4hHXdv6H8gT
zUvhm6LUzvtMG8TnD6o9zzWWED3YpVhbKyr4p/l9pXtu+V2aWidU1OSmeJTp
eUrOBQT0X6dNPgaUWGO7Bba1ZbvG8P09KROtVQtMnfTuzV2a8cmZ447pCjCs
IjZFaPzICM1saf4CTMhQ+k/mH4WJMciAcxdCIbLvIJi/ZDJ+UGAGPxIdXtdH
/maw758MhHqJTWVYLoKcwVDI3+e/nerFEIbW2nAsS+OUVrTNAqs/lsnlWl0q
pl813SjTrDluMKSVo/POHjb7DsvGZ10zNtmbFXVpp8amjwEUhQAKYGvWHZ6G
aUpFJHekT6KDvIpUjgqpdZVp2QXdS8i+HhWsypfpaEA0Q+WbSWb4yEWx+63T
6roUot1roWoi5/e/NigF6a7tU0lAqLus6DbltyxathNVrQdhfMmehFUH0EBv
OLxuDmklrqK6K27OtH2cZQ1Y22QhnEUQHMDnAsJc0NEn50JvDKmjqsY0gele
mAmdZNsS1kfy4+YMTxX+F82mgK90rX+qvK9LRmoWtIuH8wG36NH+Mib2QCB9
Jr+jbH1YIXTLqJagh4kuXrQzGVEWyBWaPtHqkqH8W4nQDYFGylgNxld9u4mQ
ILwF8UvZweUySuwrkQaSTa7BbNKZc8RHacHONIN6plui1ukwwLsvwxUuVPK/
offGdHoyCRu7HCqVvNJ7+R+/qzqTvtiS1/ulXvgWM2YQRFXUxTlPpH1mnI6A
AOnIBHetRFl1Y/qSrcSzAohWYO4Iw0BT7lW6h/o+RZW1Qv+rI1rKCKctRUKl
GoIC4orruptzVw7MubchlRRiSEKu7wPqzzQifYLtuLQGapkGcsW1tUPP6Rak
PIzp7+ghYmJEVRkgCzSZZ6VmMKYsVDO+Boe4JFb4oBUwPMi9Bz0YBcXWI3OE
Wuc+umKx1rUGKzv2zfA3FzcoUWdaYfkbq69uZ6VaBbxdO0EvyUFeN1+ymovS
q+isJoiTb5wD9LQD+4XJj42COJL/+JdXUqqy1+7ZNbawkljuVBRwTXUphMUt
FPkbx+2uAEVOXob4HF0hFFu/gqf+uvp7M4hfLnqHEpSCrcMDpte7WYpuvb7V
Q7lPR7gAdChjTDkQ1+xhvTR7Loo9nnNIH28QFGnH6+ar6Duawytg9x20okod
o34CzX9Ek+xMmqrYKEFqw6RLoHcHnv7UjAhebSRy7KvOC3S5mwzBpNmI0y4M
6DWw8wnIWKYSBaLbQT15zFvMHWMecqS0qBJVy3t1eJdSeOkKMOQ5u9BENaff
KmBlzqEl6t4zg3RyRo5MPsYNfLHNLbrw4YTmhWP/j2yxUOwZEqOu4FQZu9IG
Pco0OhYazcD60VA4GwLOBDasEUsyvh6fdumruEIX+JtLTsi8Siag1Bd9nSJ+
CtJXaYp/gW+bS4SEcf8j6LxkKkCELPWFn8YxIIBPkOsxw0Pv2svzVNwCuiTq
Mt8LFRlAYdtwMVWEzcS7DxI2xL5xOGU1llOugvS64Qf6UcfQ4QObvDc4HN9L
No7V23lbuflzG8G/cANVfANOC4na8oUfT1O69daCucG43U+d44Aj4vgRkvZK
8xnN5KeUMT8/82ds5K9/vjByR0ihblviw/lCRao/lGi/qkClCXGRjUiodBOQ
Y17waRyFc81S7fdglqnAecCNSLQ/Gb4woq49S0vZKyRge279I/45Ab/1e05J
QZCs4uejfuud0ciHFmI1ZqQLrgQiPRxfqO8iZ6Lo1fpC72KKnIcuT57hQemj
M+F0vF37uL7cFmtPXQlBBXOgwX1luUvZZWIkFIN9kd+s3B/2CCS3hOZk6meL
HgStUwJCtktDAKKRUT8zRvyWraBw/8quLBvBVYOkaKxUEVcRsBZg96XGTdLz
ir6OPYA7ROjFRt3Fw+FuThuQ23I9s6+dPwmJcbrwQvDbS0IL1J0xR/iZ06kz
lxtiACtIbgxQmVQJ0HVrANm1PMwhDwSvSrBEphVdBsFxSUPvXhrZIlCeR8wC
nOlP0oNbR49e6atkbXuss5OJLPAro03evz1T+iW5HOdgv/ItVPwdNXPkkUol
zxKAOgzfzMvdinjOEieUfWVm3cerPlsMYB+Ruq7kM+sVFS0f7zB4D6MqjlXG
HVST7YPbUglTY7xrh/izHeQx8MI4rjh18ytMUdeSPIAwnfcE0zLRLgWqWz/m
T5Gnf31UzamdlZIXpaibk91SJT2RQbRm9oQwRMcwh68QaGiGn7QN5ZZJVeSi
3pEL9RjszSI5dat1AG0ftCgJgfxYGwTo+pCZRmPokvFTZ7D+yQ6J7wm8YPm0
r+8JHVHkQXL7UrvSXehevh3TDqUWYRt3JExQr++qlUbKBsQOFFYw+6DWhnZu
L+l1Ndn2T5K5oeulq6vSX+m0Brq10WgDVpT+uNZO8d62ay43e9K/b14fmjBz
KXiCfKZNE/JCJFg6r91EFsL//i+oPHuj8pHyY3cly60L2z15PNL3QAsw6yYb
XB6hmjfKAGqb7doUHLvmnWIMAQs7QhvG7q5aIXwR9ITRxeAGuhTVCsnEaRgD
GBDmP370m75melu4vZGYJFwuaWMb+vBqXcYCrl3Ngw7NmMihZKHSabVLVZ8a
BYZNa4hLjIFHZyR3nqhkb9DtpZw4QQpTDofT9fnsIceZdtBJ+8MI8SHT0cMJ
kTlaYqP2+zG/QouGBD6qxJvrT9lcBZAAQ+Ufpedt5tjBDDY1ujzn+B/0HlFb
gJ6CX6QyZgdlU+MzsdPjB9kiQSG2QPuo0mnU+VKbZ3H1yihGg45YnOKrcWzd
xogCkZ0+rcWlU6Q/VV3doAhLH58+elb44oa2qLxa0lRpnpsCB2uutfijNsX3
4KIEWHBFERBLnDkmHJIEuO0HvfZEK3tGzq/okmOytZNm61ELjzKvMTFAZoRA
7xO9scXIXJqkbZ9Cu1T0h2UwJpmAPQI8u6oQVh3FV6hBOHMrblO0+ZW45xbF
LV6wqVgiyLa/XIUwHKCsUREZFnxTZrMba6duXMEgr6hXObIw09rtf02c84CF
rFZBRXuh1R1Mw6KfdSluj4vVcIN5ngyd4wDOCO+HxocOoWUKFZ+8hxzr7Km8
RHIcW1BlYSFCLJwO+7CRKZgnJlZL84VCm4PrMSfuuoDJ8jq1vsIkhSC0L9AN
XGcMSb2N5d0DIcYdyhS56Uq6XPXGNCGH17JWjwIXeWda6Jw3ejoP8QxZ0yVm
OlF8TposWvIRvoMpFxTiR/YBWvcNQRmArCaPkmwvMHc2Wdn/XThB41F9QBHN
AMiXwHRkluprD90rhq37BBS3ZM0jvlljsxXX5GmajGWKdjrfTMdy8tROouy8
YmY5GZzx5db0Xlj99aPgrzokN5ZN0JdnRkwfHrkE10C0U7eC7nQzo2Z3scvA
XdSyFGJwax+muwBcifNZfDbkryENf+ZQTwuvU6wDSiCoUEtuClONTKHU/FAL
5o2eYaZM+CUpvHSyyYaE05EZb7PEEDJSG4aAoFM2BIOQwLr3vZ5AveO5bVuK
gvaRU8rNm40Gq5a8rfGqwaeE6tss9Cu4UORaU4GOxm2IWnAKHp+j4s+ppp6+
aBX9SKfsl00Y/lNiUE0fdm/ss54wyZWwCy9ISrIiXsMXGNRFvXZ4ei5NNqvq
TByLighgtIYT4dWouLsLcDUc6hYOhy5MVECMxVGgGrpECjOaiTlUPeqlPd+U
ELqEbdXKRJKJMtarklYr5hRtMwW1LSd956m6it9xh6N57InFobDllOjRGXwt
cqV+NWj1MWYaVBFMx+wLYA8ss0wTG/mHTUqd88KhUZcBW7xuBRLlrAisqzJ0
UHmKjGD6Wioc1xNKxTnNkJTqtIDjzpmx0I4xpfuVzOAUvwR3THRUHoMWSCnp
P3XK1OFr3BIEPrCrr2ZGNv90mmcZtP6q7kQF7XxOC278aYMiG2q3817RcZgb
cT7BMSWky1nbFcrBncCEwqCksmiLGpPedNp0SfrYHX2AZsYbS4gxFc2tYhsI
gpIyNfq24BdUQdX3CBFWRAI/vrQY+WX7LHwnbt4QzTw/pNhDkzereVQu9THB
Y4GBwNFPbkuCQUi72h2abN69zYViwQEqqZ+uI5BffAe3DkCy8HPxeRKoDV+P
LJgaHvf96szy7y0T4iIaKfHEumYcLWYOdDJvMOfBGcFwkovULLBB1MlL9H1o
5/cRjoEVTLOfvJOrZ4YHVV3dFZVa8zRLpOyvkx6MXdXQo/zyLKXNEsTXC8dF
hMi/YLk4TParokWOWcLvUZj0baPrVZ9PIvc5guehJCRoSC72Oh+xYh3tcUBZ
ZvnHIuLr1+wSV7mjziMZU34203/9YGBi1iepRSvYx8qX5jVaCdTJTLJf8Xm7
2Ew+DG0X09vOIoyD3VgLFIXQPUQLn+CjrF/+O9tZXLadjSNAynK1+jgrO8NG
O94qk2b2bNg6VU9y1CTdj4np+CPNasyb1OYxwqWXoMritLM+Ug57Z34Eyhg/
Mn0ZBdODqZWG5oNfziy7OfAlfvy2uX4kAi+4zaZtayZqwKZwHh6UwrCQ8aw5
/RFRs5KwsTfzcCX+baU48x5vh2g4vedwegi1RdR7jGDLEtQkwJfrOlKXqD/l
CId/Tr38B1z04yLTr9VEJou1DkP2tgmRo1aoKEhRc2sBXmjoquVLZpcHI7kO
xI5LB8EJIoDCAvLNpsk1+PVOz0FIRfXK1NvuQPjbmxuvgbPs0Sts6yt+D94M
SpC/EYgsqg9ZWskOoUtVpaQ16moe7VcnRvABpsvBNW0AMMKVd9Y3lU/xFwXA
enyXYMLvTJegRKt6DllUMx0d8JnHBu/Sr+YHpWhajl8ZBrVkRZlrpKrjVpwT
87KWBdQmAEZIzUF8qpHEKjvo18YzM7CkvUe8OK9yrU4UpHWBQhf5nbbNWg8+
ziEIQGp7Tb5TloPBrjcH0RqjGv5sj/rRB8CtSgfZy7wG9GN6MCGtCUncZwJ3
77WIeAYp2yTQT6Il5AtlGOIaTSSlYhZsztxmfarqiqHtJAnAfuQ4P1a9TPBN
mB9a75dvqySqnl/uPK27zHl1L1D3sEziDSlzCm8ZJFAaXpu0mVn1htp+lLh/
OVqb0CSqeImndT3xBrNCPOoQdCGASEYZ5g/++uIlGNlDZWX2sFJFXa5d03Kz
tzbXbHejV0m/DQGw4GMqARO/8E37mrZ/XLO0lCG9G09/Grd+mS4X6rur6dYq
5YHh7t1P7l+ztjYsy/Wa3VhgQDRLtuPVJe/LjEhP4zdyLt9bllw8lMEqamQR
5+4RqOox+VRPDeDm29okirhO4nU/EFnded2c3rtlIOV8m6Y1F1+1Kg3H7zuA
aM+Anrg4qhgZsVP1GxSgrnUq2cjW8lErp6WRV0kWZwzZh7XZ/di/DuY2t8Gx
MipCY4itfFUb6DteCJiiAQP4f9J0RqzEz0I+PETB22/NY7esAVchl8N5zrVl
0cCbo7lUFj92enzrwkv5Kt6DwjfxzBrxl29D4YajZKnYVUUY4ZYnFQBjsCCD
ZIfAMEV5nPuHGtuY/Fo4x9lPZOR7vWwUc373kVIbmGAZu24ItiGEIfO5bIsp
cxD14Bo60aZFrgPxeC90FpOXIti3DfNXJ8M3xcGUOYtD0L13CfVNcR5iLqG/
qafQZG/u7Vs8tFkuioZ9EaXGx19LJBn2cMDWdZvPTL5cXUJ3egSCXLzypjpe
VhNbHJZqIjCnbL1Byp/xs371Fc9+HzDVTDfgxqLM3RLliciKdwHYKhTFDBaJ
Cq6Ta5bVUaa3/+cqaryedul+elZO7qMTCCeqMyXtaF2d3TgyqfTnFOiHMtTC
LNuKw2i8Gt8GDtQ3LCZT7ubRJ/asHuDNtPvxEhG1XG3HXZO+tvcyWUWV2zW7
guiPAWvAK7Q4oX1CIoRnlecsLIV46/U7am2oBzoYVXtT4R9IVvCo1zmERqVq
ps5SgjkwVuDi3X6RVwBQ+kv+V7JeoL+7n5nPaXY/OGRThaOCaJcvhBpuZlvr
XO/7vp88AHBxJAyyqhz9ekgslyn7Rxa7sH6zo8mk+Y35FA3iBg/UPpdEb53n
04ur02lcAdnCItLV/yBEQeBgROU2K/BJUXkbNMXyxJHGQtRywCelREy9ypFF
kL8TtRTFMjkDpmPeoy+HyPFFgGA4MYsqLhE6M4EmRg8L89FyIR72FhTscdE0
EK2Z9ktgXQlF8wglGPkWPbwfQBMxYNkm/UERE21pCWkYgjqaEc0OgLBugMsN
TONaY44fN1f7nNvzh8Pg+bpQ9Ypq8A6xv/+FXWTSBqwubPNsiM+VpGcYSk1/
TKxU1tyS6EOpZqX5DLUh1RBcxy9jAYjDZU7h0o+kOle8KE+ILMhPHN+PLya1
M+C8sKUwaNOsbwmExZL2tf9tDQjmqgR9+pYivQgb3ag8MCmAmjwrgjleudEi
HVFWSd3aapBExHVBCP/JgPVUOi4heu9vs7i5zrwSdmM17wZcQ2kcjbWtGYD4
q1LdxVmgX41gpY4o6fjuY4IMeRODLj6e+5jd7Q6OvYp61hm/0Dd6LkJ+TLAJ
2DKMXpr0oX0HqTFysz7Li450YOj7CEx3mZ3qjnUaUw5r0feEkMzvyVIRGsyW
/klPy39AcC83b8OE4rl5QXjfMnnNfgBcObPrskuqs8ZaIC8y0/pkiCRw5bLt
kDLPhVRmaDplzgjwz8dg7Z5gfzVm8LZoFMNNrzBuzzU8Y8RrEteMfb/H07kS
IURBxRpOgjasmqP4tSbRUkE2sTbYdf/zm3/JJt0cc0lTgymzRjg50q04TXQU
fmt/HdoWYu4pp8DSBiC4Er83sCRATP6N3dHqFGEULaTsOdbKlS/uCmompqM3
G2/ke4UzaIyuOHVD6lP1qsR/3k7KzaP4N6lwR4yJQJiksnTn6Nd4cT3j9UUB
mdAGR7ETEVXFQOeX2qzn322AESmxo07rQNCp/XkcM64EAIW5gEdD+HNrLAor
ppr4pIvBy3ZeMkgEcJuyGOfGkRC3QjgNjdnWwKrOxQ4cp07Z2TovcAepgmiS
pTdiMQwZuEC2TFw76qqMYJa8/JpY++jzhR4YSggLL2WGWtfAF7k7UNWwYlda
aluMC8qbBBvlsQLkAv8EkwvmBC9i3sCKM8zq1Nm6yfgydxjfqXW2CFlBi1Z7
mA0M6TQKT7SKv3QossmIHydip9s2kOdArYqTbmkenzG/HSr7YscS4tpCbl/H
mWxGdzXJxMsASclyNeHmqpjG4aENdl5auO1G8DoHZzvPs8jjj//ureXLVaYt
v8ome82J5fjSrcYMkbZqoF97LKKAEAyKtMWJBtU+XOFAd9tgmtbHn8U0APbT
EmsMKSjPAKjY78hI8XJBqB3kv7Z/2Pw0A8l138MbapROqUbdgc+dJnFt1BW6
Df1IaDmbUosYavRwjLpCgy1J1fnfMV6HO3Fa3Mndr6maAjfu3iDQ2YMK9AgA
dkt383goFqCiF3lk927Oo6hgDhaMVBBbtiane7z8IE5+P7tpvHE2cout8L+d
nt5JyhILDHP0R2XX4c3KREHtcR8EeN0kxEKfw6PGTduLCEYs0nvvhadlRb7d
8qpaD4y68UcxEwTnZqcCmojWD/GqcsFxyoOvEh5FH/B5LvAdUfh65WF7KTl0
9lypbmUgxhn7xlvJYlKZLGus6bEoRauv6oqpOd8ctA10ifPGlFG9mcy3/ZD2
J+CkTNd70DZYcw5ryjHSZwQMuP3+8HZRBT43YsApWqVmXPnaS147KmyUFuR6
WR5npK7TkVFimaHPyGbdq0TCk3BVubkXCIM709uNeYUzHfJynk2FQBsq4PhF
3YzuBJ8tApW2QzZTRyAteQGLb87Y+sowEgTK1WM4gsMT1tN8HOxuv4FX022j
vouTHGQW2LHIyCnj7mfJFU+jteO65gpg3di9ND4unEt1uzIGXboZFv0IOxnx
ySrCf088RverbFz/3UO4v7dweHWj3eUQLiso0vuH5Q8o44D43y8YGyNerJCU
qNWnlNDbWH4UStOu8rMPTxx2uQ7ePOxE8SxSpRRpJdbn2kltSYgtgf+AA5Ai
YKuVBBXwNN5ZFPxi2TwQDqMdwOYtSx+W/xIBycNulSGkJyvUm82CqhGk9Hdo
wCuyHAwKNIsvQPKz5Is8P7VwOmL0DmqJgPwC8E9tE4gJuRIQv/WsI24BGbrp
BkVFU0ntaIAZZ2dgUZ8IepDFQw1xrtPCl42SoSi+XiZJ102iDFY35C0A8mrE
qf0HRgWEuEhUrI5zbbw/xis14SQpOz160H+P8Y3Oy3mOTVspdmJsNiOtlQ9W
LPe3Pzd7dJAADUBgC4JqWA/kYQS3l545uy/OiBVmQawNxf9lU8ivYcDTswby
D6Myhfw7PfCie5OK+riIh4e+ZrbudnoawVreLCjZj1a0W5mNu5RJgXPRXq2d
EC4L6K2PD9JKYfrDwRdGYC+nmhKS3ln7hr9OyMnTDRTZ5id20u6b71BIMEiF
nGPI8zE8W/VOd4ZkreqZ2NBB3xRKDYmVbQ3OWSDJPm9Wy7ETy73Yqy/eixfS
8B86TYCTcW6MYxzK8GbdZhO95+mXfcb+ZRxMLtSi2a9/j/xK8O8rN8cvhjQX
lECUgg+h7E1DmwDatwx+88/zKreKdD3fBV1QOiQb580G2Af40taGQCVbWo/v
akOaJlnkSL8EtPvUOXbegpgUy8R+SBIRrnoFcXkylQBaEMN5rm8T8LBDU05X
UP44FH+sLwgF8toelD0+VAdPS6AqRw/u8AV1j2lnZ1zkwI0V/wMsVl4ZKMT5
8y2inwy7X2yd9PN7b0n2s1MUYZOsZT8/F4ioDXyNPDTc4FnI4brfHdMcpfdd
EHe6XBSyiPis5ylatuhO/CwUxjbzh73/rK8t8hi+kEe84j7cdv9Wf8kuy6bv
4aSsKnXv2HQ+7lVsKmdiFQ4/O+IlsOTMrIVtYbpIQkFsqONpTWzDq7jdlpOA
NJj/yhsdR6F+KxhZEJ5QfGg1eJzpR9d7xu+q+dBvJwGwsVMoVh12BWa6HL4l
G+hjE+xVnRTL8GVgbWUO/NBrtMC8Wbc7+6k23w1AmQqm9FazXMfTU058lRdu
1h42PKhgGCDfNkLSTovHlOiuoNsdV/U960cY1b3C5A1xh09fbqqKTvt4G+4a
A7B60EOjReq9TyvX4jtsK19cryXDbFTqL7nEcsedKZ+Ia2KUSY6cF1BoelT0
FkqixjXf5wRgLwJq5w/Brj/KFj8G6tM2gsm9AfVQygee7/WinnGLLSfYj7kK
Tsa84VlTqntSRA8eVWWDxH5oFI6xMKfuMx19amPD01EaQRn7HC31P21AWRrB
3Oj9owl8IN1bT8w0XpfDUu7DPHaNwzjm/Q9/Uz/x4Qjan9HY3aNHvz8ATUpm
JWMtfGQCBzGN7MB8yqSUm0mrFhtub4xaXxMP0QL9amLP6hyjko1pAotZH1tc
ZSoI4h8JEGpuIb/0/FeqSzISZbTH+8xFDnoGpSjYLCEyYIv9/bhAxnkxC91m
Ul13npbyyUe36miEy4DqxDR2XNsG28PxZ3bd6GuwcaXMP9f+5L6qpqC6Oaig
swT2ohNQu3vYRg0U/RGfhDrenxaeiaHD4yq9YIvMQyY3632eqsktMQztk6Ja
Jl6cojb28lnwAhzwHOFN8Qt9oyNcTery/WOHLVQm253Oj1z15IU1f6ldc00/
6IYI2zY2CyY/yty2RP3kYGekTADAyc180YjOZIpWIQuZSmbmJwZS7l16PkVS
c89nQPIiVaIFt9YcFfL9cCa7+99t3hQzgRvmWCFIMAJgvwJ+K8gROGVHwQHc
5WscUTqBeulKn1hYe5n3rOA2mKdw2ApyJXynjDerlL3FYayxulkwBCGWXYS4
2VBjBdKQKNiEINf8bF1uvUUEjT9X+3bHhxHWCB0//n02yP9SoImY9Fku13p7
ot73g8bOEj5RYaJzHFmZiZVji3S3Jr2U2LIzc7dIzWaFuZ0sp0TtgMVTZ0pF
f18QUpJ4LCN4CFFuJJFNMFukfsy7FoYLjhGIe+IMmnF9PYuUUnew+ca0hZpG
Z9LYvof/B5PkFk9z9VXcgQ/AeirQdZadsSCFWcK/wrhC+5EN7lcXhvFpbD3p
LUw2u0mFUc3AQO9gI+1277jwPHzXNinBRZOo93vjo7Vh2df0/2Foj300EpPZ
x8ybIYHWIIZaPCRBI8TwvaR8YU8bVjbyWqY7Zl6cyK1uDq4Ni3Jpy2EB02C1
l2VmXtjT00ZVHNJPpsdZcK0mXLQJ4FeMf78Bjx9O+PH+TswPDGL/p1KEJGXy
dG9gx3eHPpFhioHsq+ACV+Gls92fdnglgPc+x2oc+b7HeuGQ1om+gKgiRrr9
+yggftnHxdePsgGIwCmwTcXQCE80BjLzfQdWF9CNRipxU/d+ChchGQepRkow
5jeb7I08vr8lqRoPlf4FHW2eHr8BgTrKEsJNl7VcYY+PtaC0Lv37V6ECKt4w
hZIZB6GB6gS/xqnqUQcqUQl5mXBLNgevKgDCO4CkQj/flL/meIKiBVDG7BP2
f6PNy40TzLilHoHEjAzNFW/d3Ruf4eFi7FAJG7kKz56UGb8wOqO++X8uUYmF
TZIU0GlWrxI27Q7WVT0i9OyqJgH4oxFfp8gvrHP71l48CW6sOMVCzmTsdnZ3
IPl2EveX2jU4HNGdjr/hpPqIWX8I/DfUR+o31jFOYfYkD4TKcfx55h+Oui2S
49LmihHUHpkIf7bfcqfAnhtR3ICOlL5ExgBYznR4zCas+XRGZ8zLR15cRSlu
8RBleQ5HST+xsDP0IuCIOgtMo4GlsBepIpX85DFg7oaX2OaYFlokClRBx2+X
EZkgk21zYNp6nfgsSXe5ZZRdtTHYS5n/ex+pZ2KVc4+wte5FO+sTqDvslU6C
7I+L07YniG091dpOalxL8SDqE9b8KqEMD5xWeKLJs86WQcxKzYn+qI9ul6Xc
wkPKBaJP0HWOhaMT2j4hF1XOeX7RKZYRlWHOAhLvvCLbyDY0Sv+4Uu/49Xdd
dAlI1oZWVVYPhSZLbH1u8yBBM5vJWS5ZXElB7uaEjekkdEPRBE/QqG8TeLSt
n1vQv2WoiS6PJVnDXHQPEH9HtUMTYaB+cjydZyHJ2bQkm1Jrmkx3zaSYglUC
eaGMtRNXi7FOcc8DxQ+pSVJuZdGQflptj8Mw2/1EnIhElTvF5vYKIBzaDntC
Y+b7nx4vEt4zXYm+Pl38khilvmCmeDhNi9FZqIiEVH0RTUftoiszCpoaF75S
yiqWrY0dPD7fYQWaFyyaItzEFB8lQbIl/5IyiKnRD/TUx9OqMn+hWG9MFVP7
+oFiAErUsxU3Y4nFuOpMMWwNiXHlWXpge3a6XUN7g9hAc2awAqGvvuXyiphp
LIkzrnZQA6PMIAgZMCLTju/1vhTpHcNUC9ObLJdOikBfWQEdWrcvnnbYTa/V
xRl1qOJKi9OAl4/wvjKPa8sDlnUnZPIBT6nrOX5mjmMbvLU1iw/eews2lASk
xszx+GYqUDTgO/hy1ZaVypjeKKfeCJK6Qbe0K5HZQwLDt9MA8KIfzIq/p0u/
yKzOvJwoA00IBU9hcw/vKVYpuXRolxTV6TxO4g2mWizoQjTwAej5C3zmcXF3
ChPIamYr/e+U4e6ghkz3W8AXV6uwpn4NFxO8p7iRbm63IUpQ5ASOqEg/d9uW
E+01St8NgRtMqcPRNUNf5brB5u2VFXbexNheBCQUcD+tc2vZW1//Gw4ltO7q
8AvqSmlnMtW0WR6dUybVnujU+BGx6PSFupcu0x5ZQeEt+XAxm4s/uVY0TkUP
oezU6S/gRT2Nhq1xog8mJTEBjvN2ywfrWTnWYvJTPXB9Zfc7ZzYdpRs8XXa2
AiulWFdnhzxpyqkt+5q7qIMznSkQYorbLscPMPHj6HcwbWdpXaqgNu0L5DKc
509+1OaXIqI1/36+dLDDXZlJI2j13kzZJ5InK7tIUh7+WciFkxQ7opsLKZPc
wNmuaVeeK40xbRxz4FeM5Qr+IItjbEqwfgXFWc8ARKaHPDVAo0u1od7r+Try
c+JctMc57rEcvMN0JWT0NVrtySxjpH2KS5WhpvMCr7WkFos1RieBK5WkQHjf
1VufefLmnwBB3AJv7H2blCLVF4nSw1apkAtrDDGWznSX4B+yE7cQGjok/7Ar
E6A44F9F6fqB8E2r289DbQ4WgB2RQfSzLN3cazeTaU0OOpTO2dBV/vGFJPAC
zeX+bESod/AYTpeWFhUmOSSFw+aGAVglHKG1SrnjVs5/ZWF4S4qoi1kOz9aG
HIdvZDP5T0XsKw9fRgOR3H1zqAOlW8tuM2K4v5ENq0vs6FbSa6yZ1vPZOLgK
Bsq8NjBohagCJPsDXxSk1uQ7V9TKEBQ59g3F8k+1mlPWkh+DHe0jWmM6Tkt/
hHoCypU9d8kPGnTZCLBBay5jgjXB6eGZwLy63oEFcY080LcFc20qtIwjXyC8
PWIKDXyd0lU8oZIWQriq7YkvGsmPq2ZSKGlR5i95Zldy1gEy2TnBTkCZPPMc
3JIizrV06FNILSuVG09KArDhzH2+pIzRtETG4eg1xhxlyX1tymMnuGXTExlZ
xOIuFtdFbb6TepERKGc+EKzOtETQshnbEIlPSJgPahPIgowQpdujXJYpRbG4
9Rrg8OK3USoGJTC8K5a8aMiUBi8to6DXdPrmYHJJcXMq4YNNumntJ+teOgo/
00qZlTL5kmLRyxWQZ0EEbA07ydnp6HumEMZWndBPEk+2RfedszTNP8fJD04O
79oaNxRn9X/9W2tt8ek2Gb9ODmy5V5oXmMuT0xWFmi6TBUaOMBdVjEDw3O2V
MNvjY5ZrX32XJUmZiQJewvAXnZyM8/nZo/7w7awFP8ogUZqZqIafObnzR/tP
5EMsDNg3CR9F+4SYGV+30fhBVwqwQTk0a4eHqAN8ng7QzJEFGxtx5uiAaNNT
vP+x8r246/YWX/akYrohW5qv+Dqi4I7h+LKGbMVqp66K4Z7VL15wjS7YSWeF
XrfaUfDgZAW5+R+GJ5XeSRKmG8YOOEBfvFu27J3BSbcG4BMR54SX1PGye0Id
oIJthERY0l1VcmSzE/lZG5nUn/HMtjb6XpLSYj8SD6bmiCrwb+FCn7jIelM/
OGdo1G8ZgeSsqnyx+cYCxJfUhzZPPKEjRbB0bfe3cXEg+5WLdd/v4gb3IZ9Y
az8Vy7Q9cMlmFuWrczuhXwWzpc86alb+VIXYLXqmyfkg7XkoNigF/xyX4bCC
jQHhidmphwiZ8JDDueBZLyIMznj9U50CZkYP5z7qGUCGb0dlok8KKBw6JiGf
9N/tznEsNOZrq2Zy7t18PPk1ibjej7VFZ9i++RDE2UEpbkZ0NTOpx+43I9wi
3d5uz9BloK/o+RB02INX/NqDZN/IC58CZe0KhISUzUJlEMQfngxy3jduvSrq
6c9Y2P1Iz+mPktl/XhVgRFwocYcMrpqexSSQZ4nmeP2UbJQgBBkAp7yRA7ny
A9KcNkSs2wDFhRbX1jQ2++xCtwCvftxTItF7QN20I5pEFqiWOkkAJ6OtjmNN
G+xTshThWldxugoPhjNDBlfoFyLy95MtLwtcUJ/F39ET6fw2CNU91QPEuFhX
3D4ZUEstW7Md1t5SHjo6ovy3zQIoL2JBKhXXqGXKyf9hHjYbSrUjYbEe+eYb
+/oSz7C50B0Aep2QqA5DivvZ3Dgh4L2uJWTsxmB4YGaNCfnWrd9eZeeI5QjK
aWpkiKiNhPh8phKa8iiCXAFCt/4oLCIf2uTlbOv4WZ94ncoG6RW9QrskASAd
qeEdQNJgFsUEXgGyFzlNaTC82ZlJGi5kpA1LO2VknM8DCgXZ+ReUj1n6B/Uq
XkvRQe5IMYnzR/NOropKGQpVdRSf30p4P0J8MRf8C0khm51N28BomxdhCyAv
cV5Ao5o9djgqYESqFtrDXg0J/a8R2dteT4VlxkzJ85AdwBjStEP/4NCvsfcV
Iw0zExXrgjU3hPyt7IqxFosQLrzoVEsgA/k1zPaEberXFKhL36cZlHnSU1Nk
fZMSByZyLWOrUVujO+L/7T0t+aRFJ8scP1d6M8FCRV1RVbeT7s5iu+DeNOYU
ePghvRzmnbtTe9HzPHghyDsObUTWU5vGE8IsB4AeIjfXXx5N0QJnoPNwua8i
4sDoDje8ISz8EavD+gTTZ1vo7uPFRChD8gNAxNzK+XoaDIENAN8XSbq9UbUJ
wRKXVz2I/gtt6QDp0T2taopmhnBNvIberK1NOoG4Vn0SVl3lRd3tYxmzR2fo
bezEj6EXdlTd2514TSopy752IY7cGrrYBdbFpT5jCP7eHFfmAtu8C1Pv0VCV
nqktwSbeuDAwktW5j6Yz21pyY/+dtsZQOX5sVH3cJFQ3naqdNmpj8GoRJbvf
ArQGJqzbeTHnUCySHWZMqJVGPIfzExmArXbdwnLYIVUvVONfLF4JbJfFZVPG
/WHsRXnRV2srimoe1LhJbaUCQ2km0xA2AE6mQNwXqOhmKnadwD9xPZirHAB5
dJAEFK84/OvSV73ZursF0qYYCG6WewpUXPNr1jYql20/RdxUNRVqxrpEcsj5
Mom9PvjMdSM1q9HUwxqcNsR2D0rXWo4HVLANbdRKpHRKSV5/o+2PdXcCl8qh
LrkYesMAFXJqO2QATFItUCBIZMtnXZCdYQ0cMgjTMZjVZktfsACoDQL46tD0
RB6gHlCdIRmFiF63POGWsTC6E/CrsiMfVQAzDMVOx5oAqI2QKDzBsi5QeT8E
NcraOdXJmTYw3Ad91nduf+tGI2L+n0/kMiJmvY5i0vUS548HaloSBpUKvwft
ZuiBXFPeKRPmPMJLCzv1Xsn4JLWGqVh8RnQGq2O/80V4GDwd3bR/LDQhcvwY
8F6go7eZnp8QB4jR13lYanGj8agngDHGaiaSaXSe4KSQHyG4HqLE8bTXHqCl
QW3GEAURPS2J0hc7Qze7DxhfxMRVhLTNCq+5pQ9KLCatuxInC7il4k1GiG1G
mYq4p5hAambsRKvvs8L9Kt6rjcoxJCmS4oyCcvBw81kP0daEECJzieKVhBo3
w7Og9qIyYs8TCv1GaiGSo3oRebYYIsvZoMw5LG3MrxLCs/X0lmjrtWPW/lRb
mEheX0n+ROOB+uAStT/9iYXrBuy2Smb1FUeH9lJJzlNCDHkAp+hWCI7sOsfw
s9+KJdK5DDaYviA5zzTclmLVEaBlJuUg/iKKwxGfCA/7n6QtJccL1OyLP8pP
gf2QNjtUav1Xh8XeFy191OAEhKrt7Umk5uLOzi4ztEYZENzwlmjJ8schwlgw
HB8NHJY3BVvsQ84P+6tUA6E4jqFVAOYHusiInyCKqX6s40+kIBBiYT9/8QrA
VtziV8vazCzR49dEa0H1Q8VU6jknIgVCwNEzGTnP54w8WdqXjCvBWU++VLxQ
xcPMPXyGDU1ld+zXzzVqpJealKQYClhYrTzFo3Pprieru+MBnoAyY8BcXwLA
FNJ+0APqcsPjRXdPw71hq3X91Vubaf6s6nsU+yhrDmaTzyiKNsNu+uAxpocN
knjtDrIwyf88d4l5J8zg/dgXYezcVu599FnMsbkfHTZ9alW1WNUM7dkVoTwM
ofCRCYrmJG+BwiHJffnWe1deLDX7bMASL7K1co8mRGsbdRGJlQ9RDeDeqx1n
qfNdWyaE1NuxAeN6O+GxYVqu+c/Yj9yYONdF6Q5ajyl6LIOEU2jgJRjYOjYO
T4LkG/w5VPbGmx6qMDQkJG0IJY/6a31NLanNRUNuSlxmJeOI3pdZfWzXFbP/
rJGJuUryEdubq2MmFjP1ToLdb4e77u+TFpgYoICTwESrO9eK6rV/imDLTjRQ
jDAaLMMDd5cJdyEC5mXIyLa/4AtcQOvNFfpE/u7qG2CQkkxEpgVUSC2zhBQE
zNgFqHmauxwz4L2tj5B97S75heA1T1s4ZtZ2keeCJXRdOVTJeOMPDzDfotO2
XSsqopNbfSVVc/yAB9KtHLmGmp/oxk+GruMebijsmXZ5IwhrW2LUCf+jfpfV
EDklnM2turs76bfkCPU1EV7Vq/SJ/qPJdPps4KK6zZsSz0z3IGpek0g39PQ3
jYiZGCTpyqnigsekhlJwR1OScijD+7Sx7qs6H2zfRjENYqPL+e+UkbMl7n/s
99mNVEZynwACY6W6fVRlSrP7vKWWynYl7IYyax7lC3XL08Rsyyfd4DpOenKC
hGa0ahTqWOe0SR6K0q6rMSHi3MK63nmGgJTPkzZ+2gncwYl29HDZKNq2XDC/
oSwFzvWkxjXg7dK1Oe37cTdbsaRqT0d9IQGhMAsjEWvBuQqYMhV+cuVYOPnu
9aUGPOurfn82a1FUipy+8jnvVvJddbO6gxOv4w+1CiZbPXGpcCZB+aaR/Pyp
YJaeOIvXzlgYppsVytFdSgLZsi/F6z64U8zPRm+yyWJhf3LWeNRCniBdEqgZ
NEAZCwDZF2U/55qwzpSvU1G/977CkKFPjMHJgcm796X6XggyuQoDmLYL03hh
QteG7t/ktz1OKod3412HwKRKkYCnNIFA9vGVdB9w04d5+U4Qrn4r9DV9nTVO
L5ELKcjhE4fe8mbGJaWmb8PM5SPmRTw1c0rIMitmv9pD8s+Hk7Im7/9QRVds
tog8mK5lIVd+wdsw+lYNPyro/6JnAjV9YjyszPgu+lp5ixQ8nB17BxWWSc0k
7GSXtxd6pd07Wcgr/8N5Y24vNazU/kR9/q1O+/WCpJ1Kvta1LqW0GA+S3wJW
4F1LpiIC/pLJ8IiE6jFvWrd5EZIkdUh67q4WwnsTS8q4RaQPddvGpwjWiKBt
LQx7FRFNY54CEvTojFnxBaPZlxzTjtvhp+Yw4QX1L7iNW5pdfi2IbA0nh2+f
w+Apr7rowcOpa4m7VhVhBTkBkmlR4P6UgWho61YO+n3v4rTn7RbCvNzkAXNS
yLJ96YgdU/ebU8mOuY50yO8iweIIgCX1wsQOZdnJTiGr+lzsI9XcxPC+H2Yu
BkwUSwTApuopTfNzoPrbHqr1OHR+ENiyVkOsPOl/Jl8AG+LFWoLq+d8N2mkR
LfY3uL1j763KBPdLn71OOpMyiriEQEx+Wb5IG5jpg4D6RhWUytKbJ0Sb3t4p
VkgHcC2QM5dJUAN0hWObplmWQYrgthp9kHAsiAkLcVxS+CvEeqIUhvwqiHqJ
n7mdGT0QMVoT7/qC3m5tPWzdDLA7S0FvSCYDE9Mlt2uoECSkfGIl93kOyzgq
aWeY1g4ip08IA3MMv106Dk1sQLzXuuxSUrrvNn0l+Rka9KgMRCeE2atUF6Ex
qD0DsdWbcn1tC71nCGHW/NyJYzyypJCVDdbD/g+zPNE50Kf3DQIWl86TVeW0
3JzqPGtAl8zS/oy/PP5+81fg8tjQM/8q0CpVFUIj49FsrktcCikrq4y/iVch
4DbmShwENwjGPLpWl3/vbiC+HEJBtrjMNmjDR2BK+NOf52aXE7ruOMiAG2Q5
rjPtd31VenuZaAohhze9Kc/h95ibLbtNXt+hBBynAH5eW17YDYEYUHErfIDn
qKcFy+NOf03clKbx3Aj9viObFHsOUJh3s8CVaZwyfGJRxdh46G0fAjXhVCIl
aw0YbkQmJ5Ix/IqOAabd3Le2u47qNA0WlkSVRzjT74zUsl2lOa7R4Q6ZSXpi
/eO4BGuGdAk3rIt+Wzy7iIfxFPzFYTPR9ZftRPHd9UfKxWYEyg7DuVlaqkpc
Lror+7AxcBqpVk/sgCNfdB+6rJIzM4Bdy/YFGKM+CHzvvWs9EV74Is+zNmRL
C7Fc+o47cAR+nz7NJHgF9WBsIVnDrjqWDwoBb8NYmtq6cXXPx5PXw946cRAA
d42L5LvR1SFw8cy4KblKrhpYbCfiQi/LdWnINrb2qqhg9SCZEBnUWAHqFRqt
ImMc1w7MMyuFkwNKNqC1b3dz6QyYaCqogKtOJ/3uvTZ2p1Q/kKLNAT4a71x2
ZjiGCQQfNMyCD18YrLZi6GXGF+CUQ/NuE6ose/xb/yP2hKY0WoNf+WO8RWu6
0L1JrkdG3S455+AarmJoMDV8Ie62aOe3/MLx45ZV1vPNEsa7PjLaT6kqDa+l
Ab5ydD4PD/b97WehHtxXlv6akJC+FJ+YMUvRrCX6FlbTChrPLdZgUHanBC8V
cZdzUqIbZqs7gs51Umhc7Exz4Oho0ET666szwmPNf6dl3i7Mg8BxstBwA3Po
wkHxGFxApwi3tQS+cwGP65ehrIDpZ7Qgzu7zF4fkMmuKc4aYvNO2lVJN2BUX
wk1+xsiTFO/R0eWe760Gef0rhkirFNVkfK20OWjMti7wej4QqtaFohpOt4sP
QP5Y7x9L+61pu2PPQhQSZExoWt6D9RJFG9j3aN0E9nEeWrDFqfgfqGpL3PTL
u75uLrRepDtIePOe6JqMoUw8PRn4ZLE052azbY4AO2WqxapgBFiNuOFfZYYm
WXtfkqAhDHasxX1wjo2keJhUcjgViQrS71kujuH5s58RwVxoucEutJyAjO2R
aoJZRSdNrwf/mjkd4yY6kt2IijNMIXLb1zZ1wU8JQL3gOy4R8sAwsS89ahsu
Kl/4f1J37E9l0S7L56IlxbkeL+bWlBMZsH2Dmd/KtspjVX6DgbnbWhv7SyW7
PlK1hj/wojQL+5GHjE4pei7TazA3vgFUzX/wr8N70o9NtxqHwTvZVKDxjtbu
33BO0KzvNHBIztukJGUs08AkTTweGm8LkCK8frnUlNy/mm1Gx6lwg0QDzntE
h/IVBxPDhjNiGYxmg8h30qhsRjmTxtgn7C+dqnBPsUJz5bdTM+NW3A0ZxhoU
q/UqBOXTe7xaFwAb9RUizRC7tkBcfMUxNk7+Bd/BXWfsacdoJiDJj952+maU
Jazdu5DhGRky8xwC+TH1e2UcneDhTbFvXaUF/tYpGR0rx5211Im/Pw9t/Qez
1+/4xMF/s+ggSOfD1+DbbEZEAQnDlCHmuA0EFqtLSMiL+Qd/grGe9rkVa7d8
V5NOdpviHj+c3zC+6VlIxpGuM0r7BimCvnhXhhzB6FRJO5JFvYuOaOpalMhj
uzxkJPdl4V64gELuTv0czV7UomEKtmNbEFY9wV4eHqqKNKNcpuJnRsqg97zr
AF1nKxrsMyNVUQHmYBEbUSMv0dwFZdnmc0bV00TbjU8lSFL9aKr+JP77lecH
Bc/W8bKJJP16+KG7MkQlXumZ/ZUPWZ3nAt4H1mh4x19zR7RljCs2jEZ80Ttm
RtHhrjiL+RPagv/BZroKS++K1BJyahzGWzJLKXL6wm6ikosD/P0R4QlLF52z
53t9HGqDGGXP8OFJ+mWiRpa/qYv6pMiLuJ9SvdqixuwIBq3kwfhHxlq6CS1n
F0jp4x0nIAFRUA9Pvf+aFEOwV6igxZ4ZEROSoq80rUn3ULKIeAAMz8F9sBc1
DVywOaTXacNk0KdHH9GWC1iR2AIMVKSlDP2fhEB88IdkTxwfyCUD9rQF1qyi
2LCn64/YkcpS+Z8d5ben9rQCZ1xQifhidpRLWvF7wlxe9A6He3u9LstG/LTi
6CRw7UAzvHFojGrQa4InKNkd9ihTkarzenb8B5krf0yQtUkpefHke4x8YjkS
bguYeu/u4xaimi8hvb/RlAfjtTlhgy1cJVP2NRrMSPo16KybeFi8qSRqkrxh
p/2E5u5DzHfuk7i5x3vQ1J35pb5vlJythwJVSwVykwTwwLGgut7SAf5fA/Sb
aVUPzo2NYAMFMxt9TjBTpm88tNX3SUuzxrQLBiVhKB1MyKETHpdaP4+uFW3J
8hqZZBHvTQHnJV/Ylr9vKetIoEHXVv2MZvmf6xD952THGpfI66QR8HsvOl1F
y6UPgfvL42Cgsqz76DmOriLHTf7bE4txbgIEu7gaobZm9ST4VFEvkCrYgrUL
6aM1H0LyhrEfEXVlMrNAmendwDKhseVpuHI8bhaJBYCkX3IP8Yk6eHiaqXLI
0AhB8ySC+1XJn7xyZpZbezrhpSEna1YNF56GL+82qQkcIZNJVbYBPE+nGHkS
bV1mL9qLS0PvA+0lKleaOizrMwwH7rap8F7yFTTYTLluVKAAEf/3K4M8EQaD
yuQfxDD+XMY0UhbLNvcx9DzEoQoccq/LetiAZ7IRc8QfwDLBvmhx4v/JK5qh
klklMJv5k4mXFe+1KpBa0k/+JnOGhkLsfPBIw2yL/BDddO1Evuum0ilIRYJl
Ws0K7W6kif4yoEZFAqfK1bjlI1sZ35we05plSIZYODY6DcPUh7CQGelh0SNW
JZq3SkQwhWgjGTiBopE/zmZ+0yuK0OJJ1+ozdO1FL7Gv7SxAe7DphRdbSn8H
CvWOeEc6WJT1NKWAjf98iTJrF1fu71QYifk+rgGqb7Nmnl04dHyfSpKXN2/n
kUt7gSRTHHjWqY4GT4fyfDTT6x0FuTvgS0gGLFSBopfKL59yjUCC13Te/NX2
gok2rJ9JGD31He3OAi/EAcDUDdF4g8c7sf6a78uE0wu6JEqeC/qmgbsY6S42
meT6CU9cqVjqJdczba2UM76c3UbS663A+/IpSmkDtJrvPE56UZjg8ywE46sn
LeU5Yi1tJ7BIY7Jc2EVTKFjkw9u2vVfwK/CkQjybZiix/os/nCNb+5r8huzM
dcwGrbhgkkYoQiLAAmfIvdCOdgWdA6Xn1K+4ub9d4nXQL+ESUpiZuq1I+yUz
VE0QTYLy3hqYqU4kg0O8QitNB2g70P10mjSGs8X1bJuexQj9v7DdKtP7h+AF
3R5H0A4ntPCSGFDT4H3BxozoyIUWIEzmVD7zQFjwxE4CV9XY5RWdnCxrvEyl
YurNV9yFqG5WpDh+jrXH/IXoQczeUDanavInXTLxn/qEJoaDydyiZdTzdMui
HAFJt+gtyIeyDBCKK9M2luqlkgU7jsWFfZzdPO65Zcz8kVkSCvApiW8JNS1+
MWzIRaz1f/mJk+hEhEYIIG7WI38DUhgkz5q4ay32dVovCt9Uzu09JoFnXC1P
U8gHEnIFajJEXUrQc0IRdyoDNkWAaUkwOzSvgSBNKhM8yo/Lp4A624FrmVGx
941lQa5QdflDtXWbEDovAkyz0FA2W74pM52lGGOE0cn13plOUElZrsfv5uyW
3WZWO9A7drcvKgrw/MwLMiG8DQN9EiHDWDRa5+hZc6IL6UrKXzXDTdQCYU9J
0l90znNNoaZJXEKExCYHLl7qecZL8PFmFCMMEUZ5ld3CrUvwop3sGt6Z+fjp
GOOCRz4IQxAbJOuv8a9o0c+M4Ke6DHZmm0TpGam9T6HSTh53LLNsXRjlX97X
N3xjrzAMsdNIA/jvPlwczk6A5JN1fMIJg5ySEPLlzW5fkIRV7N8oEfcSxnX2
PZ8Th5B1J9NKtmCHlT2sT27SRGk+i0180KhDfzP4cz6vCBzoBpMll2Etapqb
Vx2wyukmoX5+eCLNYtb7RFCfrY6+lHGxlhljsXh0x3miyLGB/9zDNB7hCvLY
lhQWaU41OMhGDIdBBUiuCHL1TCoMGExPoUZHRL7w9PMXX84LPlZhGJ3jYJr6
IPZtxYx23l1P0u/5cjBxwhxXILG2VR+weuwl27JKuhlEk8+vrVinlt5CZfdr
DvzyMD6KvagOnXHmNr+KNo3ocoWKoBpIVBP/Sc6gDqpp3SXT9Kpjvxp7wjce
kNcjY2IOVrmHm+/6BXkvpUKhCphzg0rpHHkM7jhCR40/fhop3Msk59EALPWa
Tki/9LqsD6TTYe1sXqVimEfKUfNPkQZsielYhyTXqAbQ4AIZw/a3BvZU5oxl
wxGkzHerngPfKKVEyNLW22Ialg6/Fey4FPM8bIYXuD3FwZFjg5gJI8/RZ38h
NbOpk4tXrgP9u2vWKT1WCu50Ifn2aDftnALUab1j3wyxNZnZLCDtPaxIzN2q
uU4/OU4tw9Bwh7cMjXGwP4POP70C2C1NYoD9q99wsrFcysV4lXV/LG2l2ekg
zvcR2p5uRDCy/ZI7j1pnAoBsHvvV2cvFUTP17PYZ5pDBYR9KoleiZbHIhSsa
VaJIniRNN2YBsFwMn7GMqhabLMrosjkJuD1yf0eyNbvM0v195KQw4oMhN6Mn
mM15TrIM4Jcvi1H9/8SjpIz+Kuusf/GRd8erPPQKMoG6lYFueDqHjmF3Zfct
Yt0Q2kGFip+IqyiQoXdQG89l5VFwe4HOZUQ+5t/2CIGrC/+A5+iFFELr/sKp
PQkuGLs37BuUEXqOBLA6a+5BN/T93llqAKdI2ncdJp4+/UvitoSi3joAjvCQ
nk8Kn8xHTy36Nz9lLWx0DlwfqhrbGieBPTHVMR529B+jGlnIXH3+biOqqIbx
2W6lWmucPHCCkT++MxtB4BddV9H98p7U8Q7iwKhLwxf3zcdMBMHPGqEuPpqQ
NOusJVpn8XZqTcSZy/e+lQk3yqxpuSKIpEvPFZ69IM0LqWdkZyZitx8d9/Gn
iBM0ITVp+RlxVlrh5x9xphsjnmeoqXwyG3azW6/c2QH/Zr35WyOB0XYaphpf
w5DX2woBXkq7BYiKIWEHHWtJVq0VhofIz8Qefz7CsacHCDBlo9BjN/L1z0i8
kelV1ssB7O6aXM/mNDiQbAAKgBcItIoydP510zBYMtiP6r0LY+ktBmo7foRO
JFdxMJBloTpKkXsdGsE9wvs5IfapEa5MhM+VFhwJSYVIbzI8PD5wqXrX3Duu
6BDHpWDT3P+Ao0k6ry1XFabX4zqNIpg8Pkg9PpIdEAYkUSGDOxfbedb63Juh
OUnuaxu+VOescCoUb61uf1MpZCuL0hGqa7mJuKHJqmHO9s/9w89rJgV317XG
Kr0jxmqswm0z2M/IQjJ1XHPRhktOnAczLQbW9QVEvOu32jh6yFEJwKiUHmgk
cMVqpvUcoKHhHw+TxFv4XcgHaxvj7OlWnAkLb3x3hB71eaSAx2ROkXIfP0k2
PeFqtdMi6ZmwslN4pDx7WldpluBl9jOzM9aBX/odxJub5/bYLtMKCSa4UeLy
NqB7eda/irsbZiVb/AI029kqJyvwDwqIJzNESKFxLqgBa8U9HNVd4iI9990x
JGf3ZSD3SPcHdt97HxE0mV6UtqrWW1q4OAWoVcjmi+wNbtQ6YX+goIUMgEqp
EpShMXanx9ZL5ItRzZBFHPf+PPujUC0zZBSff/M7n61mg0klshEkWQKvvyXo
HtIjm9s20VnxS8nmMTs/BNDUWVOYU1TwZ6LtOplzpD5rpIb1fQX2Clqfchmf
LLS7cw7EZ2PLOzwzq1BfCM9LM39zMXhnY/HjPVWTFDwpQFAn5iAlEx7l2heG
BJGiyNV/pgUMmbik4OGwcsaspA9l+yGK4kolNcfH7zQ6cgfSvI3Cv+ShTlCp
5o2ibFO1LPDr+LxRLaSnm4jPsh7X6rciI/Yc9G59gZR/RH5/0uV6k1adDmni
1AFOpGjDo4sDl8iKLnnJQWN4opfVqyEdBUJdxF0NwvmUj2AQ+536u/61st1W
mTJJfkdEBowlynvtaC8nsmD12l+Cp0eoXTmXoirh7is0f9FJ6e05R3W0mOGl
hneys6s3VqfpsW5SKogd4INIPl0sEccPgIEq2D3qvHnofKUgZ7vJh0YcLHib
+ZwgT+Ts/GPUi8rylIHP7MdXvQIf/spIO1pL9EszpAQ7VnbnUMoQYsQIPvr9
wD5KNz6Va2tAwj6f+H+Hi/rgOxCekltx852yZjwFwsaxITmipwzIhmW2AHy0
OkvMpbg36Lb5PiHCHaWI97TovwyHyhQsfQ9Xo7ZuuN+0o2SpvAA0yf70T5qJ
BwMJ87nWb/Cnac+gTT5VcPkpDDzY96rOm8WQyfYRhWScYa5Krhrvep+IGzxl
aVc2/RKmhviCmjKinlZzyAXr8pg2igEe+Rn9lViR16QlnayTIC5XvWmpuFFK
nPi6ryD1TPLOw9Nx00VRDsj6u3WFg4l33RZd1Sc+GFAp6lxcK//sn2bvyhX8
XsGCRV2KtTARLOrkWydKO7j/EkeY4PF0TQYnePksIv5OXp8/E7U3+BUwB+WC
ABokuuh7FaGkN7VoKBR/RxOHk5yaYf+0Os9DwT6J1XPUj/dHgkw7r1JynUoW
UoQHXQ/9gF9FekAYpqLFhaSx8Urv1QaSxGftXP30wro4lQQTYIWpAroGVT41
4AfG+UwCVEnap+oLL0Xufc6CikI2er9bEDg5m8rwjC7JhcKyqpCs/bB3Vkh7
aigAq/TUSXU14Vt7GrfVONERzjxRizMSot2sGaDnnF0G+QE2dsHhNrbedJ9t
jfkBu2YHwQdWgeSfiVU60Xp+CXTV/4Q6UryJ5zuUfHlTrT+C2UJh/vzU2Y7Q
f0O4J/hBnapHhilHE+c8GZJB++twLl+KcrnQ017HhX8th7VSwHfdg/T1bViZ
O/Qov4g2iQ7rfc/nZZuBm7xrUzQyaOoWxrariU1X27alOZ0n9z9woOMcN1Tu
p4eGsaOHu5m0b+EVCpHmSm0Oid1490JYre3SZK9qSlgM0OyqMEESHV8+eQ15
Td3gpY2PDiKw0MUhdYaCOrcrSkh8p1GD5FRgcqCDYmaeNC+pxH/M0Y4SZ9c5
a/hQWivulW/Jo3F08JWvS14nyX7obnpd2uuGW2YFDQlvxc+c0E3v41lYwby1
MG00Fcf+/sbR0PBHOP4z5IN9eB/UjrrEH4L+zUT45imY7ZOlsQyiR3unN7Dy
2iGr5TjDwXgBEn39vKZGgVbf5/ejiP0jOW3UUUDFjQim5MR9ErnarBYrkrYQ
oejmZ5v4+2KwCyHxtiH2MMdeTIshHyUThICgX6Cej3WqCdrf7CosIWSQ12kW
8FdlhHhYvP8WnQS7yUYQ0rleatho0xUiewU4x5HygNFkENnnPQXrILgBLKFl
QU6m8afERkQisAiECjZtcgOpO03HDt/YqN4JwNSWWC0WaduxI8oqG2sruNAw
5ETls/O+NY2JLJmKH9gkrraAdfhdnAhxclOT2xFHi6CZvySiUdiNv83Igbnq
rQrNPBdwOP02k4NelyB/4HHKda/U96KxW5LNjF9U49Psuigdw4qTqmJbA++/
sA/+E1NMwcSHmHKJUTHMBOlxoLhv8y2nBcdJl4lMnYWIAlwa2wUZ3ePfhOPU
f1Ml4RRSt1pbyocSQmsk41YVnMQK1bH8Oqwaw6qFJN605XDb7KvEvtrNcq7W
1jt+69006FldFAXOuO9Hb+YUw5ltM5MGV4uxaaFr8KihfI6GRAQh/3alnXC1
jVxgSsZb4yR0jYb2fmmEVjjgnC5CVdW+FQ7I0aEgQ4Z7/HMGO7+7qZnlUojk
9LEa3alwh2CD3UkB95OZ/OEi8iTXBkINKQYy430CDVOsXHwx+Y0Qqdfn1gy4
5culgNRmDye3um1g+iuXAtQ9wfs21a6R5C+hqIAlqkp8qD6H0PUx4+q7YXvO
ltVciZxaEeTPUFeyogzMfTARPIOeBPU88qob8la4EHd1YBg79idW5i3ncRb2
qCBAvWGvtnANC5DYfps0uKYUIjk3M4DaLa/1bCyNiIv75T7pFPeKF4lm/Zso
j/2/chaLikeYk75ByqwPwQiVNtSL37poSexpgEcHT5ojxbT4cE4fiwHE5VXS
NqFblv0YMkLk8qT8vfcSuCjwNWp53ipQL/47EG5Pp+SkTWkzQh5UuAFdGOYs
wsFU+MBlxj7XMcXN9V3DOQFSc3JrHXjQE4n7ogfijVUPghQq233owM3LYt0U
Tn7hecWw+zAnLgF+gTOkDXFXbB8xOalIEi09nVNY1eoJ0rgVDhvC4b+9XAA/
KcN1GFH0L/W+SulNYy4KvMNhzy2XbmKwp+3vzVXd0BFpbDa2oyODfjNa+9tw
DxAoeidOPEoLHKu1sx/bbNdIOkENCl7LWwexCAzjEFImJztRDn5uhae3aQuQ
gYR84jWfkFlk96Sm0c8Ql10g4r6cB75WdxadCLQULmzG78HFHCxXghwSEkmf
m1URQCI2tKlLBOM6eKKAtc68JNAJUxtSqR7jU4TsZ69PBFEzI09Fz9GW2a/P
CnCYJcaROJDhHYw5vYzW+c29Ii8uqUEPuheoFTEQQT5ya9Q+TpJWOw0Qqn1k
30Z9yUjOwCP3cG+K7D9sqnjojKGFxozOxVgNh9EZVITnamqfpAzC7Vf2li8t
m8gQtSvCJgjiB+otdkCgbg25ZUvGH6tJ+YvkvcvvzElPLdJzY6nTjaIsqpen
Y1k8n9yCiQZ01EqE7IsILktcy7MwgObM+v81xf0kfzA2Gk8ye1rqd9NSkwxR
5lkgTPedyCd2KEORBhic6jiXRgKUgYFXzdCBa/4673eENAL/S82L3ArnObFt
CRj5mDBdmPD/FEeAQgU98BqIKE8/AvqbPbffmBv2nSpgFL8usfTvT5xf7/k1
miOxy/ZlcsUgJp8wA/KvEQVpTsYIMHrp13O/y6RC9GG99sWU+J/E41c25u09
NISK7HCYK/YuwSOu9XQlf3BhCQ5KvtQMa+ZSV+8NUhmIpFmmzE6tRcEt2+D6
ALG09hbThXAMxZ8iDyDPUTxZHrOK052F7SWa4Dc3nJpVnXp9OciuofDmesTX
JnZZx0M1n5upgVPEZXlAGELA5OeKZ8fyx3I5n20zC4x8pKLxcFGEsqUyK874
+mjwVd8Tc2ROESNDO9Sbc6t/7BgpM+kCF8bKDGrVb6yJPn3bv5a/UU2xM7jq
nynUAuuW5HGHSc0dye9RtxkhntjLCYfjQeLUmmyWFklTPL9ccQ9My1hm92Pp
r7ssreeO5mJbXURO897IdgGtsfWUlJzLoD2SiJ5Kt6wgzZaoj7wjHO1euvxX
qS8JDTb3FpjDotTC6whKxJN8hmrm8EcUozJU+fDdBwRsKTrQXNg1tR0ahwud
fkbl3M/464WFs+1HTOqPYSpqdBIgMWIBLamuRPZInudBH7BscXcgxJPaHUWt
68y8X/9z62KqgHCxjGZgq3iclwlbE2mkQ0Gx9sHqtY10o7eVwVviRn9hFZBg
wyAtciKfcoQGnsvA4WlyyGXEyyOWf2nQPfvlTaLvH2H+3nu3OWaB48ehy1zt
nDB6ylRQIxmFMmTUmaqu13102rX171c1iyn9J+v5mmTV8IFVHDsnFGyn9mLb
spSBKxYhIKPfh4kInhjdsqfutF8IUu98gjajCObF5d/Oj3YbTDikJ/5TLK+L
654qQoWbdzqAgpOsk8HYIAOxy4K/QEDtJAwzwSU6TOfAY6G9ONn6RBQDb/HN
USRbDRXy7t8uZM8nXpdvl5StEtb/t6u2gLeryL+ucLpy7+J/VN3vrHhvPTIo
CoPBNd/7ktPbUu6cqNcm405jURdpLV+REw/3pHTp+1H/TAwcWxYrcbxek1TZ
70waeInNgbpkOxnsOXa9UReTQdvt54wveElU+oH09yVegAyyQRTywZhj4QRY
e0bnzQDYPsL0/pPcTnlqc6EGTdQe1C5f6FuzSclZd8zlTjVwgPg2heWXGqEH
GMiootX39dxJnUUjR25JTv3gRYQyxkgJgLFsQVENlG7r6opVGsNso35+pUGy
C60UEduvbhf7rSpx/0/nj/ybBc7XZiAKeEd0T1ADuC36oGE6euIElYN/KubW
VRb75RP79AWMFKW1gkVvHdlq8KjBAnKNoaDldc8+MNFhs1NvIF5W+vEt0PFl
e6QJ38/GRa8yjm0owWTO0YhjUepmHx2KIseVF8Af0rNRu6bAhsZpM/ZzOTyF
f2e0g52yVGndFrGGvInwsi660ARnYy4iHlTJ57yTFzQFt12SrPCAtXn1+gda
vSx7jinIcWeGuT0H+ubkQChP0aN88KiAzF4n1OLV9cBWcdIiJd6NJ1mXtVwC
E+Wj+PT+4x3AKwLXDMz+/t2HzM4Xtfa+sm9n3DMbI5wMSAq0rEPWbubSh8L4
l98SfrwX9GWNEinPHUpXbUK3p8RSPmLRYd8/P/XlLc7mbZ4ROTo3Jp0lBCl+
z2Isx/gvudYmGEnrHTp9IIGZPYaiBxsRaHAm2zGWyFNHQy8Zp2eOYpWPhyBg
+v5bPGOczSBfGFX6ulRXNpJvwBOocmTnfnpBACVMUvpuH87SXQ/vDZ9JsQJ7
Xxhq9Yr55hCs0IP88anIS2BtqGgfWaI6HbYPKlqCHbE3hCqXRbJ+GrVDLriT
3NZgGPb30kOuQ+MpIk2+L/0tYr1MePP0SNYsr0ERzQ6XOfrBpaGQY5DWoDg8
T05p0cI2H7oP0RulrHwHJppgx78nFttTfKRbBd7MaBdlnYEQ+nKG2vuIGwpE
zdMSVC2J5VwX3DGds70WJgsQgXT4M5V7C8+rHRKNaO3F4UqcghYnc7JxqkaS
nMpCB93B/kf8AJ9V7x07nkivpz7r7MbycVrqG2wSGhlLlGrmqF3wRYLDAnf+
ECyoDk2nm0lS/pBIVxNJSME9ZxdnV7AFq6EMEMj6VP1WfPwPu/7bXwpGe9Y2
PcnvPCPE20HaR2cLchoRnWEjlNYt9mlhN4U7JxzHUgldl3ehSwiQSkRbaoaz
aEVateNrle4ehPFp9J5HoJDoIiZCrgbGiza9NkI7Uin2YMgol2QrVyMwBPAl
wIXhkuO1c4kKnO0Wo3Jscm8ivXNM0NXJMpW8uaPAzJY/Crqug/GGgwSFHdmN
lEc1mm1pT79LsTJIZG4CIRHXUc0LWGj5SBmTsuPvSOe3j/TVvBYxhBbyhSuw
CnsfnPen/yiNt6nSz7wuaTuvxO/LWf5bxhjNUTwI7js5obRnqi/IiwVL6BN8
1cyCC0yzodBAmOil/7q4bUOMwD+4jAdAeVGmc81xxkd67N+rynJ9G/De/ZL4
Lp5Jpjpb0/NKPUuu7p6HRX1VcBOSObufxR1PuJSiy5sr8/qcThNPNxMMX76k
CwrtGBQIsR3vHynC+k7/VzYo4HhGW/wo5VCAlU9g2fN0gRwN2vjTMvy1hpjl
UJfz/PYXQ1YVvuqdj6TgjVXIgeXzBVnek4XmpZUOhdrqW+x0P8mLyjFZ8Er+
OwVdnr0WsiV7P3mxKFou3SQ0Z9FqYXeSmvsG/SqgqBnkOw32eAB8zcePQZn8
uefGZFOFIwHEOH6pdwbe7RpyepTwIVu906gmj7DNP0dZeVVpgRCmhnxBDiBy
0rFpC3HtUID6Exc440KFulgQ1AURzuf7ZGy+dSiAHlQWjPMwQP402TXzW+PS
oTxoGtNsdLZJ6yqN7lhR3NzhnIIi/P8Zt0bmQnBjS7BkhbD7cHFU5HhAE9Yl
VSePKZSYWu9iaGFeQCIoCx1+Amuaoo8zoFD9uASTTqUS/OXjcpJXQzkm+5zi
cmShOuxXusYf3xoJqeQrs7J+geDNrYwq2+M3qAhV8X8HsG5eB+lzI1Jh3Erw
7G2C4OrLssdVFc5Yz6fEQtGKrMbxpR+q8LAgXUGxKj1bN8sd21sheEoeUxAC
dzNobr4X3+8EwEa5RhMIdyDN+xXXyf6Om4Zvm8RuhpyspsI2STH9m7QVDEiw
vp0Mf8QtWTXDzzYU1NLd4WdMMkcJF1v3YyJvFdH3g19+L/DadX6g8Q9pvUai
ZgWhwumwQ33Hznf8+Ypg7nXLf/lRYLC37cYt23eeo9pWnd1Equ11BKncc+z5
Lu7HUrb4E8aWCDdO/RxHCKA0/4Ga6SdJjYsL6ZYIbUz0zH49fCsHcprfm4iE
nPP2Wfv/K1kgZN9ghD9osHlnE64GI2I+Opg3nDCubTax18M1MK2BKi3EBmhG
yxFUHS1LmV9RjWVNF+4QpykMxq4hW3c4Dl0j6aJfy/b+FWzqJEcnLBJIzAA3
wQp7rfGylbR6PSMUj3BOAAtNSXua4x3D8jybyKFUZh/ca69Vm4ISWBNRlP/p
BBqbLfMPIL4SQCeCdiYK5+/tWNZWtLpLEWUobNbRVUo91LIG2WkIU1tLNbK7
gu36Exze8AfSMoFzlinMY8vkv/Q+I9wtZyV+Ghf66u0UevQfpZtLb8751L/g
lJzWnf4ATDZTQrmkam/Sgvf7rIa28QR3Z67EudUBbwPzZ+rz5y+1bITEdNcn
OM3SnNBYeluFybtgrtiL8Wv6fcUp+N5Rh8bf7IxcGtocXuZr2X/E6rBDwEjs
WcKmjNPSPPLH+I89BJ2yQvsOvK8lbDTNBsNl8QNYrmYpOCovDSiVfbKUg3Fj
LyDY5+2UfOvOoWBdqRV6J7p739eLlVt/gYphH1D67L0cPEUqe/N6vx15QHht
GUuqYS1pWDQvjSjHglGhht+kN2QzRPHzhhucc6A8wkIa+o4FX6B1yQ7S909O
dhzOZUK0p7zywDKQvOs6AE2ub5ibSRYbfe6vptXhuYq3Bysrc7hi9HiNvRb6
QQMhgP8sK2MBL9Q8xJ5dot5p8BOv07HSX0ZHRZVgDh7FXSQUBbZILpZAiqip
LTk9m1bS6CmN9vmV3ARispPCLCh55fxsQn+luJ5p93owpDHn8QlKm//7Ldqz
g+jU2VFDzJZky3RT9t7j3us/mAwbgm6EaHtv+qvoWMtF1UeCAdI0+l8SM+eN
TO7z5mvb4kC18rlcmQwfWM2EDrhdfnbCkEmIU7PGuni+HptBVMFxo6FJZ7bc
QsOmFLXl061hMmcDXH2Jxq3uOuTBsgrNYAb5qm97HvqyCEydLGZavXVsYTOL
9QAl1Mh9evLCx7UaY2s308mSdy6MXd6n9Zk/lYG+G+8sHfXn4ZpIxjWIZDtK
nR4YX0i9EJeBsUVOfQ2QoDJZWxb0UKmaPfuma/9vdFeuOehQ3m9ksJzWGnUx
WrkF/H5oWYBzsL346QNayeuLLdTTXC/4e0D+mRpVOMgylTUNXEKctSDPc7Mc
oVfo2UnV8mpSK4pMEQXns8F4Vx6cOlYVr5ekXrTSltQj/gNRX6bqrvjFy1fO
juNG8tvm3IRBnxrMdnOkTpOHHvOpwi8vMyLNgZNtzSZ5jpHgeWQZaIWIsIpI
yx+kQ5OJwKsCg+/mIj7zMmyTyztIeEOV5i/Knb8MdeFwsdgSC46qhyHGEx6J
yMv98pP7r9T5Cv3jDX9rInaARPAuGCjCKiT2uHBGMD286fuUXKPCW5KpAWGb
xsWQV52P/j7IfTysEEc+erz2cEjjKbXSnR+7IYEMcVidiOQp36ugrPF5P73d
Yro5/Y6lZObAcOLU6ZyckSBfi9GaZ8mQy5OyXJpspeKrFaahNEvg25F31UCz
zYQGZXht8xDVr8AorJQKr6hivfXIboJmzxy5iBydwdUnXeMyXFbKcBzv0fbR
0CswJflANhr6YPgBQP+FL+SjrUKpfvCvJvwcrahlLf2NQHKFeU3/a2nqKSPD
Y1RlSJef0nO1Vgs5YuVwTJiIanLGgXMlV0Mx7lW/hGnnroI/Nn61v+CuiVud
0pvEOppBFsPDnaxdIjKHdTrcEpFYZ/3ntPcHQKSnorwo/57JKn9R7p0gXNrW
7mZHdek8hSRQy8dRsjHHHTTHMgDlF64tXKZaPgAOlNS8HpPviE8SO1qSQQM/
Rb+dXKkDGpnHwPn1EKS5T/+maJ1yN5Mus7hmHXH4rMLeMqjrDBH5DuFcgHpW
zb/lWG8mGg1v19M4ovTO/R4jwJw1Dwfp8/K1mcik5S698Z/K5GDnhRSRmqGk
9TzcrwoNON8EPST8dstX+u/MZhUp/TaRndG5khrgm61sT1XCf7F6XVWZP3vt
dxuZhUbDOZa4k55UIx2C0SLQpo6svYXJ54HpChLmqThqPnMPYsl0GuAqEV+M
3pWfMIQrTpvZktGSQgw6W+/4YYZH7ceAc1PYihFMQQ6Dsiv7uPqBX++LIF2i
l+rcwSPs/FRfjWl7HCgNudDe2hJEuhgKaC3by7KFyj06kbAOf6/hCtYrT8mt
S4+vuMhcaiINK2EjfEag1HCTUIKSqqjiiJ2dTdj9FwmGFMfOaZGBqIwt61Tb
DU73liT886gjv1xP47Tm5wCNYKHxlJMSNL6azuKHkccOAQ+szU6IKo0K3p2z
x5FN7biv4T7EiWPj1/I+C2qANoyjOiFOdugPAFryFckIIitgW7E/pMIBDp4/
C7xhe1aEptOlqqbEbQBDoKaukI0VmMHGIeYVA2jYPGMECVNqRDEWrP9HAEjB
SFJuo51t+/Y8Zf6QDmuJaw2v1G6w9xDODarkSVZul6690FnPBJcj3UycaEQR
DbS2gvSQcp5B0oKUppeMqr6HcMLTVlT2qkGJZQ2eSNy1FifbIvoc7oCA7lh9
fPQs8bzt9Kxwj0gwthLVD5wfLSFZdaDeh9h9vm1HOaCcJIYtgc/W8EMXxG8B
F0tM8BeAapNFcV4tolqE0zbPfizUBu9bwBgy75BKlUfcj0V3S6KURg5xqGel
mQRsXf+9hrcWwu4s5djob0Byy2FKlen7n6KY9qBMX/Ht1OvsqzjQ99m1b84K
VIYDh/4LWZPzW4s5GsIF5R3nLjcN+mN8Yk94D9whDqFS/mb/BTcVP4yFIi9v
+rnOlsdgtMY1NVxZytKObGUagj+B/tQ0vSL308Jq44ohZeuEZSnxHc9PEH9C
97jHPPP/adjtHSuq94VPrhoxs6V2X+/i7s/P1wQ1Gm5PtCQorexpVm0vEseG
Lv6DoAkaCpF44wFxJ95+wWDwONZJAGz+LJP4atczHQQRnRjd4VtdatoWpOsJ
kUUzFd12TwCXKwneSqbPWbgWzZppWMi49NSguIi3ulN5XJK4vmFmqryhA02v
EDE20bj6r/yGo+dd3wB7nsrcchjCOSSopFYHgwdR19tACRSjO35fgFHN5pR7
kgFx1JUZa5LkmGJmIjA/RWLB1cL+nK2I8c0XVGaHXpwd65HQehHFrPcFkWav
xhORnh9tjRd7SMpLI9PO/06BgonmhSAoLovECmIfgKQp1KLbOPpwO3WZFB5/
OwWjh2NkRhxR0yQjuzp7JYqpJw6wpNrpFqmX20uQpNsOYRQdoZholOHgwzeJ
WJZ0I2iNKcwjFCwftuzw8KOkS2SXn3MvwBDRkZ4BO4FJ3tnjBjmMjFfPBZnr
Ku1ppWjGuIjkHFFYXmmodjPnyRYWT5UyEwXSBX+hICUcREgKgkfvzfaKtboA
DUt0lDwKbGzXZJVHCdB1QBnGj8Y8eyeg8vqJyCnIqaybwykQyokkj09Oo/5i
ndZqcFtIZ2Oyf8EDgMCpeYPtBpPYFzBnUl02vYGgCpVCRyiYDLfULiEJYYeF
BPSvDbYZnYBzMfXQyIYjlTnpo1OWKpL6sKrtayjlA6kPN/fzblpH0aXwiM01
vqjLMQjbym5Tnc2EemdUO/tHTj1tn6sWUJXTomiBaMTUXR3Q6cGFJnjINop3
/OjIax2XQFuA/sVatbEJzIqlWEMt2AD5huISWVNwrK+LRAFVylkJTjcbtMVh
MQ16CRun4MaLlCRXBWadygSWXGB2Kn4+33cJ97WOgBygwy4uPbBt2voyrkNi
bcTDIp7I9FmRTRxLbLZu2lccZzjlJAOuLMo5+BagB0xPK5zY6zAxlyzpSQP9
hGh+3jGBSg/vM316Ep60idSHZ9iUBmi3qFbfNeU0QpiC07kCurlmjT0XRaNG
S83dUdT97efE9quHiwVNOfcGjNuPCLstLZog3ULWBJhu6xn37dDJV6iIsi7p
DTRzdfR0PPcVb3RRbBLtvbDjZUibpFULa9yJ/m5xogi0kqUaNwcw/DNyvZOv
SzZzIjFyhbmlsIsxy1jqTVLFwYVoTyxL3VQw42CGp/fqK/9zUFKrkQumcB5S
kZmlFr4Wi1vSlB9OZRDGRct+m9qrrWBXsmPecCaRx+m6G1YrdqO0cT1smp1i
Gdc4mmXx4NVRnen/NhLbqGq9i3kTugMFOdiqEau01G2vRJkg+qxvYcAKwPr/
pvhNKQR8Z2aRRY/3SM+PwLjngTlexeM3FkPETYiAfXhaxMrUCg2vMWsvSczu
OC/uehBbBOIZymzzS/rwGLKZtRGhH68aUIDHUw+S3jgf9hqU1/YLmyDjQ/vZ
Mm/VnPr/HlUtHYE77jU8KKD3hWqSk4AeetK3Yg+NjmcyCCBIzTosy6zfW9Z1
/Mxm4J6MuQSexteqyfhk87gFgYwqsQ1ls1BTjfQJcK3iaCxESJHgXWxvOtdk
Jntgr7L/NkwmEZMKWnqr7c8sCgAKb2y6ST6yDy3e5wdYRLJsePrHuBhZRZvs
2ktYvUVW2yFdFS1nVRfDw8XyP/2pwQTG88SjIThEgRq3mxe82XBfrTW5bbSv
3CnIsotvIqKOkcewjNd2rRg+wXYz/Xwi2+olsii1yFunTlRpifEH6Kq3F5mL
UZaPEeTAwLMt2PX9CcSSWRfIQS18Z3OpWqBoRfEUwpDCtDvhjPlwR+UQdlHf
voEVYpj1D09fJaDhZbBY3EKjXKE44qcus0keCByH+mE3piQWofuAvoxlnfOO
2pPF9RTifnDWj5L+UedNCH6hBhFXWfFwX3Tc5E6ZyKG14YMx4INoDGfFjrJI
aLoN0Z07klVsBl84fgKge0Za+Nf4S/NtJhYxyBsPUg1GJSKKkRk/DoH7ydtL
ounB/Y2TnyC4765Cg3AZty0nprUd3fq3bKPTfySZyWqBDD3QLZfRkM8uhUYm
1bZQiM4Dpe8lTaahf45ibk8HKCLVZwhioiC9g8j0EeQCLGfODUO3kbV1mVS+
WuVd5BwdGn5onyzioNCaVF13t/VrXuFBtHfzJLIAIXZwMonNbqbraA9spTkI
PIpcWj0G8vREFqCFLpEbGa+0xvqtKb2aFDcpSsulMo5Va1qFmDX1hs0iX3BT
w8O0OWlMF2ge2koA6tZ8o1Ag4eKuaxr7mEf8/Ks3MCNR9QjxVhUUQPjtR+3c
mcmrSggeeONgBSOpxttL2QaPmreZm69ww/Qsk1zJXPzcMVOmeP3Ro0WV6N7Q
07sM76Bhgrn8sAa5ZYJCtmoLtGboLsNVy2l2hDh6F8WCLmAZxeTLncmBVpI1
fIb7EblCZpIuzv5CXjRrazzYtN171WIiP7FhvHR9oHSMzbFu1wRCxHvJThy7
exNXSDChoC2jfXG1IzOAz7HLeFWSiELyaWaE5NVgXT10l0aMXm0FLxqZUdMN
azf3e+PQ0yYFZoz6PmbErewDi/2J/Mvk/hOrspWmONdfKBmjGG7ZpOdylvr4
gmugsmYBncc8MlM33HcQr4Ttv0nS2/NTpSHOcf1Ngfx7Bpr0qdzrmWUVxcsj
zR9CAdYiqEaNzmtAgN1e9jPxRJEZ2EM/q2FqLXOJI7UXcqCFNJKltV/Ar3Q4
ON1mUyPgRHC36IIxD0xnzyFf8NphSuqrCjsn9QCXOb4/417SEBVi06XTwWnW
FmLTzgFZI+TnTm7b0/mwILvO+dZtiyF55BJUEIZccVE8YhJD4xShqByHkdcJ
ccn09r1pL+kaXfeW3PTrzAZHzanfIG/b1IyqV53vSyO1ezvAtYVZW7T2KmLI
GlDRHNV1DbYbnaPYgJic6si7yTKu3K6FdRPYn0KB9ZG9HjXMLJtHtHDo25dg
7aPa4wD95w73BJoWfrqYJfDAjRQc/2DBkwKOjEz5TNbaGtJBl3QQhiy3/zdj
3zJfITiezjvM8/rUBkwJDFqmLdphkD0PKHDX7lPj4/DITmCKzdx7DcHEg92N
B3Hbjm5NKUXD7eoTrAHNIQHK8kWfYzA3f6bd6PfgRWvF9/FkOGjjipkUyHhE
CMIleqJyKfMbK9MbHT8YB7HUKPKJv0DdZ4cDIgOK0JgyQeLVdlCk8FqW1FPJ
IAMucQxOZ86JPuIEky4eBEUJ6PCdVVRGHtBImWjSQJosEAK/FDOQ5+3BcQj6
/EKsydvB4fiOHbdozzBnpYED6HxD0j471R4TYtPuYIUnhyw8RQHedIouxi9j
AX8tY/fiNMbwayozJLQAjIpCt/X+NZucEwNOz6pO2HVI40PjZR9L92bnQFdp
f/9qqBN11XkEfZrqvopeGsjOWtxFf8d+ANKPYLNagK/PpLIZh+LtHCWNz280
r17nI8P1u9qC2BthGo9catxrT1eY4CztfZL3yxFPu7DHr5piHEYD1dydLtaR
g3tDDaOKBV1AgcGMGBO9uYeCKuh3/9j2BMFAs6Ivl8XTl4A6C2tl1ycomwv+
iryDxo/tS+ganO5iI/VIDoSacIKzHNdf5wqjOz6Qp5MOGkem8MN3Gq3j1Ogq
LSPydWhayAtpLYjGyNHnTfRdJHiJQS+dRtoU93HNhu94W29NaNxFLaJMsVhx
IhRtXGcB0qKEufPEmlmLhOT0o5gDGoUCI/pRQUMenenSFwGiGtlH7fMJbRfj
bRG+rtxmp/zwDy2eaU5/0aqJ00J7vh5El6V1XP3+cOAKWXeHRG12NeB+KkhB
cVuZtHAis+6PdWU22MLooh8jxBG2CgIrDmia4vt6O+q5nGAVyeej2a/g3en4
ojIZlAhcP0sb7L+siC5mnC5ecJdriYIP22Cbbmh9A/hn9bmQZbAiBbhpXbnp
VE3Vlj955bPm9+oTNEUc7+kd6CUMmjrpGF8+HdaiNHY/4rkmyRqxBjEHWStI
UtIoLnOJp9+f7NKqp6ToRSTAgUyQU6nFuqr6jnWwGLobPoRd/kAZJtQwHnj3
/t1UMy8UKEiWUk9roUugKPAQLsp/LnFHhyBw8PQSkQnu/iouOXiIe12/9a5y
y28kWPWvcOrf2koCOd+h06h97yGorRqvIAjpJx+VVUHDqPhOuxsCtio/nxKx
Bs+jJr/tUXK1dgbEafZi1bQKL/xLtdG+YYD2jJkd4rKHdJLwszQ0YhrSsRhl
94RU5vfw2Cx47fyWr2Q7Hb0FZ8TBovOPRlE1KFIzGzWzlzUFBYNluSyxXzuO
q2w7nmCPfXmBK0Si82YMEMsv/0VpIscHtkTpTxJrllzl/HTBkuhLRFaXd6CQ
6aIRhYoOS32IxPPGLlDznajW3HrkPTZQR7ylJqwQPk+J9qPDaUI+tQ1xaOtZ
9v7aRlm4prTSQtmtL1dB/AFiVuxFjeDjQi/xuH0zKVC6TnFC5cKuCgNlOl7C
b96xu+qtgHn7A9u5QVto1Q4P94TvasXY+MgQ+3NlvXp4k3fdeQ1zRaNBHMvG
hSDbX0txQrpP/W0oi9dhEjFimlrk0waKJdKCMLHPSev72ARthW95qaLokQXI
UPO74XUI/2aN9ggCSXIm6uoPXdOKNDyPoN3UsC3aEdnZag1WVXvZc+y3K+Tz
dMY9Po9vxu6ykVxJJPL0ZLcp5rBTbSV+9FH5WFUXYXrFYN/SGhWM8eD4RunX
wgypMEofFCKfEMRRPHXx8wbAMulnwMZrXG21qTTqOz071+KSpalSO8WDYcDq
NsoDSmjXF1lmMGAHyUC+Ceof2GNqT27gCzYqXZhES62fVZjjExZEXW79D8lK
YWkARm1H9ULEV/sWmQe3JTwbwyE6r8B92fM/XX2kiF9kLNQdZVu/oRsQhK0x
8YqonRLVFuXcbE5gQccTIqz2UXscf77cvfGTC1wNrsFr4qamdXdH35fcBgxp
pUQI4ptQcCA0xqAuuwBvxZna3JDtHk0ZCijs5/muikmwFYyd6nrr9bTBMrmr
AlgUW9HO2V8XN0bt6p8UIT2U8Bh6EovczJOc9Qkc29liBiZD4XvDyV0I6slf
ZlAc7dnZ0zHZWwO2tMkvXPk+cXEkkfYFMyMRHuPJm0D/hBo6oBv2Zyo4Tqju
osQ9wfFBMUUWkx9i3OTZY6SqNINgkh73/0vDP4LT3K0Pj2bW9yY86f295P2B
Lkf020fJaf6fM3ZJX8PwN7d2cjqAeKsdKfbJmx7hrpbpjIpv+BvKb+SaTTte
fZyCwr4cl+lnUQK6w9YfzoE4ChDNlAU3BlDzMkB0JTbGbKlUcwu6WO4nFLfB
ugfDdv6NtdVLl3LdNqZwM1dyyvVW1wT/s0d9VZE9hqWgsu2+a1N9ULoQoXHU
KWVW59lcOFVxCCOI9bERWfYdDPsDs/t0veBqMXQmmNBuN/xttinZQkIuUIKk
JZXc2w53X319EFggxAEjGMZ4L39FqiU/4td4N0Gsnwg9d9Esx0B/S4kEzCSz
6puuoOa1w+3t7xSc6VOV8P4vKdrCW3ImIYLO/VmsftIL0PQ6jhmHzkk6VAly
TEHztxTOVyGZ5EjRXNC0pnfBibo+LPC9kY1o05iZRYl9BDmC+oArNBGk/xBu
i7/8F5gZC33GyLdVXH0KZgRH1CGkLvTfpFFEkYOC15SgvkQEOUmGon9lsBgx
Fc9+mW9WOx8WUh+furiDhS2KVQggJNoFyTXF8CLsiHmcKG80BKAbxbpnWpT1
cfKs07MP22m2Wl0X5otSPV+Mna10bH/lhUJMTSlj4o0yA+rQv7dKJaNRyOct
efPjtkfQ+IPL91ufmMkQ0TIfFc9iV0J6KWwsSrwouEhbuAuy6bqMbUeurhUu
6vtqqHd6TlgKsoVsvAAs067emSjoDw4gmpeWhWA3xRGhIJectK7IroOMYppk
3lZUD1z5PxGEkMZUT7Utw1EIXjyK7Lli2JFVWPktwMhG0HXIoGeDmR/mCKjU
jfOyrnfyctGHPvwLTWOiJFbI7Yel+8MxId0YhOZrguBqDVvslPNH3O/fDMFc
JCD8agshJnmsqletQnmqFhKdaJfklZ2ipOTWtHln3Nupa9UYWB4yIGzfRVsM
VG1fsGLX+jbESD97Kul4kAgdrKJBV8g5Awr1rGBXSckOsizP34a2IMakLEzX
YtXtfW828oXeLegmS/DNSp8kvyCejUf17OB5mXCgLnPRAXGD9f4opOT6/zvA
9DNTv+DiSj0LoFrfjMuRoFiEHCl8O0Qg2lUaXztlfRK1nMVPaoJ2c3y4zYsc
ResglcDYy7cRYwhwGVkBBJ+skJ6DNLVeDlPDZHgC4i0qrtnQgdq5SPOcPywp
8QoqgvP5qdsfVr9es2r5L+GuaNl0n7Rdf6Qp2Qp1TekhTQeu/M6x0ydwaftu
T4TNYcF3T/lgUkYRE3ggqrJflWG5xzc2XmjplXUOHIf+26zABvOUlnyRjdfT
wyqvw9GJ57DJQigtRN6jtvUR6l9RwyPyauUbPp/9TA4UQaeEOGij2PGm9nfb
hl2Ta2sBYrIrZvj9Z9CmWERV6QsvNZIIZbM3vYTVBCJjCiGSah8H1ltY1QyK
ccIqwdHCGWTOJpDelNW6a2GYgvtfibPF5GhxL7y9urUZsVprFLvwt3Y8/zHe
yRWb9KTMqW22EzVkEdLP0/CCNeTBTzHipL1h1M4Mz0JSMl5xxOd72aMAQSZ+
3O9hg2xG2t1Uvf2ByyVnhsi0lRZ+fEI2kFxkKOhJTu2I6poSklolB6jRkIAV
BTSlJoycbYoLz1in+jyvrau1aSCcdB37tI4YqSHPSst0FSsktTgnYytF2B1D
cTHKqVOc1Oh9xZGbavp0MMTSZGyPip7FXj+fhDuoxJPHM7QxICMqELYWr/wR
BUo0Fw4bSkNR6bYCCwamjPDXaJp2e7tqyTc3o0YdCh1JUNgj2Stf87K8wnhI
+Qhkmkbsja1QlBg5QUcDrmfUHYits8q98Ky2YxD6W3aKhndWyxRHZ1VsYi75
2Wio0WND0+g8PHjnWWeFNIQh12LGWGjnzHihlfw52VGstO/8MfjR38nUrtMY
ZkvJN4jBYGGsLbdfvFZI1zp+Q2BX2mZSAQpmAv5z8EvrBQRM+ma2mjTlL1mT
cGYcULPvJlyHn8c66kWlmU/Sfa5DRVswZ4r7t5oDd5Jlq8U+q5DU6CQJbF19
mVewMaB69uRlnM/2KOJr0W41kc4YUr8P3rp3PvaA/C+08WehbEH4PCssKMwT
kUejkZzd+02NqTeqRNXa7+0l/OYNM9Z47oLlI7IkcW25AH+i1MfL1Oks/z5U
7eMm3ocp+brLO/eMv/iGOKp4adLuqC6Rx3dffAgHoW1UFbJpGCxVym8XDBIQ
hiFNiiL8kAzgZEXOztRpj2L87V31IfpQj/JRz9u0YAI8JL5k0i1XHMXbCPBG
7TrnNT8t4wY2UUXjXCQJU1hKl8X/kCEVdH16kjWEjn7IhScfq3A65KO0b8Dm
SaLsK3Wysd5j1Nt6ZL7m7VI5Mg6LOv8TLUpZ+IsY70uSp3WdOsQ1PB3q1/3U
Yelq+pfkVzq3HvI735AsyC1g1oGPrEn12FI3xhZ+dspnQ6JTjKuW4lkq8rCo
b+eA9HsIPr9D4kSaKCZYU2LaP18PfqPHG5qVLyspvVkFwsjKIULD4dcbDwrH
YGT92mQdPXJxE9BrZoMubQG5YLr+xeBuXeDbDMiTr4LEZvGG7owZQLPPhAZC
HNLmTad0YgrXN3MiFISVkGsrs/ed7f/QIv0xaNbeM3gWJFLcrbtyXqrL0t79
wYLOoIPWO1/pCghuedtKTTRErOPYOkswWBQW5VCxNnZ+NdDsHNnI0kirjUkj
/HxqKohjSKrlJsDqk3oY12YpT9LN/PBbsmyUZEtzU7cCPK5BAxLez5B/LuLs
H5Z2miR0N29wWJzleBl1tE+cP4BCEe2RjhEnRAmSp2rK0hx0igG6NTb6pNQq
W2RvTir3qMsFR+HU29MFIv/NF1qrO42Os8NZtxBRnPC1tAE+A3u8IWl2VRp3
Ld4J0qOlgR6ssbxwbWLvw91k3MOQNjBXAMSKF6lPfEpTXk0U7JyN7qMmAB9n
4F/sWIjzrhnjuI8SJG3AztpODz76nlyR4JSgekqjIs0vSv1Sb2wSzj72Z2UE
2JfAuf3/hG61phNkpJ0PPoQnsly/CQqyaxqmM6G4NKkHInzcyoInOPI4Dq+t
VcAwzZxjy0ksb2lysab+BPWY7riJ++8gzozm+cjIHsaqI6Qa90iqD7onIoph
nMoa1/5wmUSEZYkpy4MvW/oYez6S2wx00UucQGKwDx+txtDS8N8oxgwjORLD
wiPzD7olww0zR45p3jTS9R0lrM32NFbuNQWtEKQNBxV42S4aYg0PaqK4LuEK
+FTRhIKuhj0hG0WZDm4dnU5iYlmvEcalBKD6FD3Xi29pmo21HiGkJk0juXYA
xPfO3raFuq+uS958EMDBPmx4xt0mPnQVJR+8nBpifH8MJTV5SoBvQP/17nPq
YhmwkyOd68cyW1DWK4C+tYJ/ZX0s+s69Q52ioDQpTyGKhQI8pbQRrx0uCHsT
u6tRUu9tg6Elu9FMJ/S+A3zzsSaniSXFuGXMr33j5dlhjmMXX8gwFT21jFcT
X3xbhNJgUe7tMl427PhmsAVap3mpzplPYN5Cs2gH3JB5G1/uMZWP1Zd5olQP
CU6uO8aiDpcwFUIqyD3PeQ+1FC1SVlFlekMvZ9eZpXB8J2eORnvcSE6sIZo5
CpwIHAFrYHR17gO4dQ4R+HJS1AMvYBaGLU98WF7Ync13H8H9InWKoxuHGZnk
VsCGW2PJUUJLwtcGC7hJJkfD0WioxRhlWVNXR0s0Bxa99BA9jcT9RUlcBOrF
/RV1CBWRgG/KzebhdqyppfEtDY5gzJzSU0N1xJ7T0s8JXLhMfMDYtrY1eUFs
yiWUvW+kX6F0yCFOlm2o4mwT+GpzY6CRJocyLLSrbJXxTLpjcJEk2dL46Z0/
NL8PFuifN9AsDvrZjTbEiah8f6km+DgRQNzG1G6N5xGkscj4WHtGH+quLBGe
LuK5yLnyoZqGZFeCJmSIdZCoY+8UI0vBcaErpbA3cGDKbyM32IbutBvDYfQZ
/ZGar8qkFW8Xg61Crl8GypICw52yRjIxiRoTXdYhXuNpu/chIXlf3GhibHDw
JtkJ7ATWuRSN9V+ylIYYcKT/caXVzrEKgAPzkt0/OaeZ/69ESwM+AiN1MmKq
5y9p3FbekV4mSMbDMu0MLOoT5TcQTONcawKWPL23rYYJaq8WTgAYnpo0HF79
ydcSry2uPf01wOFE4TolwG+ZG25dOyWfPKw/YqVnFbbMCbzW3z/hJX4kj6xQ
MgoomZyvD8r6ASYQ1FtU1TNTFK1lKFas18JxFoze9VDkyAvaZiDJaC5dfNS6
+NarkJ9ZpiS76GVkCwKgvg3Y4SKO4JnrifebLEOS4g0V+zKqE3HjHgXm5KaN
q6BmB0QWQKuMK6YPOC7Z4OYYFLKRKBoESLfjWYxXb3hAuW+rHSYfWI7A8wEi
9r3HU1yYZ5KcY2tlSWMc/ZoG1tCUCEGqRjgfyNwsAuedhOuZIFsTsxf8qjbT
xfta0Hcr7w5RqOFudwLDeV/8SQ8u+XhDBrmlZ1q8GutaHsVXTWuYxQNtTJu/
6p9QbddU6fbqj9nZoMS1IPoRTIFQCwGnVWJOn5Bw75VRqtA9wsxdUuNBxni8
oDesWwIRhvTmxiOJk8VFwmRjeRQo/klBZRP9BpICNKIczKau/onmqB4bqHn6
tSLNTfqWG8cUjFbeg+kHOBjLPQPN2s1CSXGWNvWhPerAN7N1rKDUkXj8nKkk
9o6KXlJJeAuvlrendg2FdgU4rmx8Wagos6IABYzKYr1nlmg07Vgd7C+EppSJ
wIEBwcUnJ+GdeaStHiXkV4irxlaBQz2gP+xcyGF25r+Xottx7FjntGvw8KTz
gg7VY6aFT8mxCjdEodu5dKgWlD4+PRkPsj98nwT9Zmsa2DGNqRseBpO2geXl
N3P7BPeGyUg1lR8y/Vk7ziZNSaDKkMs478kBrL3Ke12EvcdA+9WH1ae47LF2
5sBpLNP4onjHSHGQyhSwbbSsETQZ/A8nQWLA0ECiJi0WjWT/Ytk7JaU6bkls
VAm+tU4qodtPtt6UwyWMcAi7/A4byWumB6bFVdATTE8wpiy2YYEUAWcn1nhs
aklqJ9tHAbTFElgHFWzXan2u3gy22OObUmt+i44bm00/+tOPjzd/2ROH6zTQ
extfU7N3KD/XurXrOk036NIChrAlebNyfXCs6TB2xSNj+lBaIuFomt06+pUR
YfP8VFvnWFnxYrVXiXt3MyVHu+1AeDgpoq3dEmvS7K9tIBQToGKU3O+PoMHo
QHCGnc+9gGN6jbPg/lkGdTbdRQGa25+/gVes1oFIvuwMGNTwan3PgBUWIRFx
W2HMCQTrAcaQJKjPSLUiK1mFVZGHhZE7ohqY2dWtI3TFqvkb2VWzmgjqW2SK
McNZ9Ji4gN0g0sLIGn10yxJMdplgliDgsR568gc0BV8nEZcUL9qdP5l29sbH
tHDG7YNDVkm/F6mgK0dUsz2wzQeloGFdDxq0XJBoJtuq0eNEuWNbI5AMEmR9
V2l+4pFt/AZF6+XQajHSh3pFy2jl6jiE/AnFeAItArRUz4J3IKP00Ejkm8LH
zZmYaPc4UBzqt6BwpBEFZNszkGliRSHuA7FjbYq38+eFnhTNJkx+q3JNjNSj
n1GZa5l/t1CLFOE5dPBJGTx9ZMbRm6twlN7cwV2Xht6930EvyRvklRrhbe/i
uO1+uL73JerMr4N6LJWjjimhgsRPz/7Yre3s+LwL5qMxftPb09zmKGFWL76N
qOX6790V3utgfdIN2VL2csYt7Br7ex8aoU9LLDofLrdo4b4Rs4I+vcEm+5iB
f7F2mffDY6M6/GMHdJxSu2va9vnSO4Ew2nW7wPPJGhlf6BTnM49j8uZIL+8p
2PNmYIRx8KLWiNH75CYSHRDycIkURoEomwuIx46FZSJua7CygeyI+IqDRy3b
0JEIUXywIym18KgKKUsVdugXOM2NpTcv5VUPPR6IADIz1cH9hIYBel5kXF3X
pu4yQ/undEvsyKRPXtSxCte4T07G/U7YDwvUovhtot4jHmHT2ZGs8/jkhwKU
gREkTlhn4ON9M/bSjisp6CcRg38GFyjoTQ5TIY5qnbATX8ztV6jiFwiX93p+
lHXQPpWtjNUkJGNsZ9ejuqzQJJ7IdwEqTt8CqlGsrHgZ2kQanhrtaPHOYx3c
W+xs9wHsVU22NB15nopo9O1ZlBAsVuwdPEfD+QyWGuMVOxjDXn00CLGPk9vd
jAspv5afCtClaO2u/fxlc0C8Cq+4EEjqntSyKzI1I3eSEDWkOlT3a/+23Nwi
jA+yxwBowqCQK9gdQ4SkmkRw4BDlxOAGFuVJfzLqmL+EgXMQAo/Fx/si+MSI
3tbgP4M8pRNdFgvIPwMTJ93yqSkh6S3Rah82shoLgXcwDHY9lKsGGXaloZik
0w1393qrgZH5GZeH4R3CDmy/rr7kfPHS25bcjK8e5RQLDlVcBbBvaoe/xu2E
xGUihPZUBi1Xs3MJKLx7JFfOt5f6nh6oubn7TBExtY+Evf238Wj+MexvEx+a
AmokL2Grm9VBW2M1eM6wE90OMJiwGSmONHRwFPT/mBko5i1PILcILithmo/V
XbEEABdMsRUm9+R1HuRIRsWyMEmU+E+Ry3/dggHdJYwrT80yIJyE2WxjwMxJ
I71yQphhgayT8a370St2T4TJmbRqnTu5kK2+H+UPFVEUMHqFWsp4ETu8R+Zo
AgDGP+VLkH4FNSnupX6XHeK9YGkf3gDC+yxNcXCPAQkvC14YoobgfxOo1d6O
MTw60lmGbczrllI7iPcWPNIKWNTx2zXW60jsHLp/zn/PMJM5oXiH2WZWWqXy
bhReKfihx8ZbjwQRlOSEDiDNqsOa5/UNRmOWFzLSE245fposTN2OWvDc865c
HeoPs5pNaNFD5pYa9GQ0+QIKadt9KpnzzIcsxsegA3rgg4bxF989yw10hEZK
mrJe+7L4k7ae8rr5iCRhq+sv55bXynEGghyZqfwVm6m+OkN+BAUW91G9tL6v
5zb5JB4jMnQx4K8KDPj0PuXeltTMMP80IzWyGaXvscVmRTms23Tc/bLPisWq
jgfEPdN/gx2zdlRhbIKOri3dhQoZqdGSgS8dEOQYWG9XIkIYerEPtpsgte6G
osRb5bCk66z9dcehfY0g11TrIlh5782liwVqd26p4cGtgaQP/IlLcGK5snvw
m7Ni2b3HJREt4749lWtePGeFocDJ1NojPGQlgHw8W9rCnATb8zOwt068Z4Lg
LoIPpWaqB253rNhIX+Ctu6lmVROssiTCcpMOv9peq7Zt4EpvocO6lnYyWv8v
VEn7HBsoHH7dkb8GxN0tsqhQoyL9lenMCypsWVnvxzpM5tnu5Y3M37whSySY
PTPh7XukiYt1oc3NYacEERSDNiyrytHCQqFWYlAPBbFwn3jVKACME82i1jh4
CdvLRgOuJ6jgmuNrj4xYZjfT1C8ydZnXp8dimQO7yJWuiUG+VW9XQb0pBULh
zzLwqEXdDIqsUhLOHlZQauuJOd0ghCsdK7IuEcC+UZZ/

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "B40jvh7ud/ahkCWXo8CJP0S9JYnc5+J2pwOdONjrEnmjRzb1YpxBEP/gM90XdEQFf8e+9j+GJABVN1VA/EUgHmy986oXHU6n9uJJjaeBsR8h22iSaiy//95eH4kKFakRZgkZDqWp0dX7AUTwRg4vZKk0rom9cx0xsiuc1Ki6fTzxDmmuuNW+yyxk/luKJogixDl7f05H1PhFx3JTfD9y6cRFGovJ+RtyYHOBbLpk0whcgaMhukuPpX5/W0z7h2n7DBj93Pz5XhD0Dr+pi5p9WXWfKHzRddcohLyBMKk31/My0zT70wyL8x8GZelXM4z5T1jQzlzTvYASL/ahk12lXbz11H5sCD6W4Aj+uqiREvssNM2UUtP71CmEFS7vEUPwkg19Jqnb/5bEtQE3Nz3R7pEXHCceZ7h/324jaUfyCeQyPudWMvFuBwhuwl3njIHdTeJnsY5LL4CQsEfxi692MhBSY2XV+rd5unxkYmyAzPE4hB2WEbTaoG1mFwEHNEEUomMtkoCUYAVNH6+cmlEsfhhWboFKksNcKiiQROCXYZGczbMXRbNT4ozIhPM4wGSnL1W+E3Vwrr0MVfOM0t93kxf92sqBUOIUhTH0k6+odUg7OYr/AwV2wSCkcbYeQw5sJoSaTllzyjHdM2MIwuKqMaXdc5ecLLWrjd+/DV2nGw/OdxM2mgLFnzowuwvsIxkkmYugjLJ6I82szwmMVHoaoQddc0xlEvkSC9iHjawT8tKIFdaL2Lczb2rB4Dv2XIIZ9V9mGTq+hKhVev/dHrQe2T34WDY6nF5kq+EQdwmyWDziM5v8m9yDSopTO8IsQ1oTCZ3rONkO4cz/q+5HLy4OA+EKzHoJ4LU9+ZyUkQnNXQRusUGJ1mnhn3/9UckYokyn1Rw/pgAv6M9+zKnUFRhbLyVXkaiSCWeJBJ63HL726RUULD/Vi3fa3YKpXlibEU4Wjt7IPWaxVl8LdXPqK9NfNeBiGUA7nJ9MtQtjW4V6moCku5fB2B81VBr98LUG6jrl"
`endif