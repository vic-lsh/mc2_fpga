// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JhmFoLbfeUi0MR9TG0DJjQ8eoB2mB4+ytjhe9JXh9aczGiS9gMBjPQjeu6Xx
alkSl63cGS4ibCFdCFCqHY7pG8d2l8q1EYN9ZCkS2MOHSzFyz0WYlWbCmVaf
6RrSwC7Tt2+ifmwlavJ96NXF004DyAgjk1qwWGeFs+qwzqIXatIGqwxQn9c3
pvJoDBGzbDi/968fGaoh5d2g9bBQz+M8inK59lR97PuqSqpDcBHvnMItOKBY
mmO29MMRA8+qRO9rVupLWcviFAtfUELIW2T1iFW4stIE1WbjumtwNwq0K4zL
PiXUPjKAgQ/G78Dvcsxs+7avUtNfSoWMj6uR90a9HQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UUxuUWdT7NVg9of2A19D+VIIqbeCJkIhUDc/rahEhcj71DWHCf00qQYjSmJr
YcoHgVnzMjGNu9mXdg1AgmJSzxYR5Pqb6aoPteNN/SEbgPLs27ov2GLgHHJI
NmKX15us+KN+64bP0jWzfO7Ge8nt4jUBbXD/Z7wFvNj+1dHoE50kpzjydKXC
45/cgjDYztXe1SU4gflslJ3+blwOvmDqeFhAP/MtaWlpfgQTJgnmFviCyIqc
7gEqO14nZ/q8VjbBf5ekTCSib7wHb/fZXKWwvNKNSsebG+1/AnGKdtXxb/S/
3pAmb5M+vL5mZfOji0rO9Ef5S4QdUi9dcZsbNWHt4A==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
k0k+Bi5Buc6Pqj6pueI1xMe99wHZytCq0Wg9AhLZVefct9V13fzEDZ/DrqTv
2KK9xmoA46+C4m3gom/Jh5A9Run0s1RXDy5fjSEiU5dPd5nhq1hPTyO2lkfz
iVpq8Bi4DH2b+a0EiRqWS1bCX7HT17xn/9Pf69paKWy+9qpy28LNZzbFytGe
+HGRhEH50oiTVKrNYCEu0iGpr014F6T8uHArqiYnKlgoZzq3Y8JJ6S9HPxul
wXhbsnzf5hri7bThq2HQx7hFBPd3AH2q+SKKbjuVpN+NugVNNKi/4SEog7Qt
Ajs0k7DhTM56lNyrxb728JcDp7DscZXl6KVf8qmCtg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TVxrOuI+MmFlHVXOM85PqXdJPtcIBXvkO1hfW/Ma9GrA1/q5udmCLbJ9Y26H
oheOQaGU9WhswPvvOoON8kg83tb+wzGkQlpEgFFyoosdl0cnH8tlDtp3AxVS
6UVNrkf57r1oH+IyCTTtvjrxrDmearnkKthbowZ646HhQGGMmmf2RM8A4UNR
f2Ibh3JLgn/fCnPUAc+N9+7cHfmxcVo164xYsXwRng9Ahxr/n64c4z/JL+LJ
o19VvlDzMTmoFoN03AVTJe2cbK7WzkjGfyZwy8Y0ZrauFdvSrPPRWIqkn7hX
OKXD4EQQtSA2FbSbH1mX6Z8sjtYi5WgB3HIj1Vhsxg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EJxEIoO0HuzvaIveoO76UFflZIRpL/7VpnbTJSaMDaEWKbky6y7ZsAkXyX80
jRqkZ2pdnJrZXQb5LL4nD74kmeRYa+s6rlmc0iBOFNebho+jcrNCiEIfFXpQ
dqRbsfxccSg6I4/nHQmILWcEc9qo2Uu4jszZ5JdICZzzjBEf0OM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ZRSL6oJf9LHqAEaO2fV8XXdFD6ssDmjyXfAva7eBY10uS9eJSqO1TzNEcqJk
F+MPq9DOyqXp+KxfOTbc3WD7FrIr2moVxz/2u3xBcTZOSfX3/g3pSH4lZLmI
nZ6qVaK8MGLjYGE29qh6HombOJOr6s9k+ArgHrnoUsQC9S8ozI/6HkpmIpot
pr5T86PXza/fEWcQoiwYyrB8RaQNxeezAhLoQdF51Aq/67yC93XFSO0SOWAX
cpUb5YFjynmn5/wOZh3s1vkhxUWthCmJorflbAyfAsM2xe6OBckCsUc2zuWX
TDiV9JN3IA5mVU2IQ+H2NVSXRXRmXr+tN5H7ua/Lk/o51xLtg9yriAeoCUxy
bmhd+DzTQ9EfnVaDUcB5yqDVkwNOdq3suVCB10wRjrJcAr4HKpo3kBLHqp07
1WRNCcJS61dTxbc028g33bLu6LI8Kh8rxO44W2uRcZjvQYkH5S7qUsOSbTAd
hyR2OHLjcAlbirBQD4zHgkmi1Mv3zl7H


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JTHttdU26dUpn/MsZkt9Z6wuaXOnzTR3Immp7UzXDhVsUHo9zxecriFgFSp+
68M7kFbbCNePxjWxUM7Zd8s35PUN5LnIF6z8/DMYV8i1rzv7gpQJZFhPgEOM
KSzfGfQNrPWsVS9KkmDAYjXGuLzdHVlukwsIuwjtpfVFlon3F/A=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nDzAU5EUQa4BHu2PkZDsM6jfrphbLvoqQMlP5bRb7KDHB/piU2b+0tuunQfH
GPasMSPAmGD4p4/2kO3nskwEvS0q7RAEu7rU1O5oM1lAbzIYs2yRMUXsm3d3
ldGuC5HUoXdAQcWE54QeVgVD4eAGe0ugOFqJ8q841E7itT8oLE0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 80960)
`pragma protect data_block
Vw4H4AEXF4yYFLtF+TZEjyPosFRjxRXPFTS7XmutEfhAVabjCfF+eOalcEif
bgCNzWhbFSrYt9w8YmXz3T1KTgdOkyBcClED2/WTYeYYz4nAjgMCgEggMIiQ
2rx5ud4meACTnOkUnx1drDojEAOlq3QuNZJLGo8Vi5mG7iTthyRr2ZPbQya6
HXYizEpZJU+8JEyjpeCKG3PujkkWiGnuzmiW7nRhLuCTDDE5/7EA9elGjcpf
Nk6C900KF+gy8H4guudNm+iBfdiz5PRLIfSzEq0tz3Wb99CSQ00HN9LglBlJ
N37Al41r4NYfyg7+QR8bWwhSvJtQJ3Fs3fY2NsHx9rkXwWdCY90kI+dfOU8N
KrC0mJWick02e+pJRauJczrhguq+PPbPMvYlB6R1ampFK466gj0G1EO703U9
xz3z6nA67CLfl9sBFHLvHy/RJSTewuHATl2avyzzcXECdI2EQzYc42hU15zN
1LoAdSK1J4MBjp6KHZM3wWG1wbOd3c3G6S4Wi9irvl/nbPBjm3LFwSIaG95o
c9rrhr77SEi3fOGDcuELqzVcuoj+c0PYklUTTZut/6z7xKTRCK3iqEY4Xq5m
GWluYb4G5dw19ZViOkJr6etBNRMmbmezviEQXqgqxgkZm3ViCiI6YTjQT5Q1
PmpKEiHGOJk3W+jZSJKCxC4eLT69ciDme+EprVO1yK8dl0TYWReFCY3T5KPH
ty3K73tgc89ZVpD4BipOs2j1joU8vSSJQyoun43ppKc+2xO65b0ae/lkFVCp
wboSyQ9R0ThmVDu3PIkputSUB35ykEvClyaTtNJKfal2fO4ROgGxsKeTHxNo
oiQiz2wfSqmDLY2RQ/ItLQeHCeo7PYOhmEwMG9cYIg6Vxxs4On6aV6ryMywd
C6QDoV83yoFs56wv4l+A2mWGpLHQ2r6qEsk3eLGnBBAFY1pYGEPzRWwMk71F
LqRq8f5hRuT5OO0+svEY/QkjN/RFhQZI5fhNm6QaKa+BUPrSNbCCUjye0u/O
n24QwoCSQhzozPipeP2xn3eFZI9ib7ntrN+UyD8nvUPrV/XU1/ptntAMuU3v
kUFe+sgVTdI/prsFzmoGP4mTB0X8RtAQFW4I27qbufrkapFoMO6HX72mtNtv
xlIPJBzDTXouHojT/uNv4p79OIJYxwPLVNdNBUkJBjCoHAjU6h9J4PAXnNet
1qf4kNEl59gMQt21rRgbyJPJUjZCIUeDbipu6Wuzm6U0WH0xZJ+uw1sozlto
/7sAooGy2TNhsVaG6i+7Kg7eFjZ/S6jnNRgA7bl6AvVzgsysd0N5y5Hwkifr
i40vjXfxYKgFB7lCBNIkNL2+QpIlmB/jwzbt5bQaED5rhUNP+kWCMVvru5jf
lOVCkqjPD2+0XJtIB5dWSwx3Y8Fs+585IjxZcdcfzBldK4uba6keTVzr+iUh
L/OCm/OWVuBQTiIaPydd4/9ubQvbygO+UgZKCTBM/34xGezR8cWZjCYRhWUz
8wOVYTpqXUeEr56T/jYIuVQDnqlds4M47t/BI+mUKsrvlC6o6u3Y4FgDPgiz
IvgOQNrE8qSVww0/pwc+LjCeo+hjP+gB7FMpCx5w4BHNuVgpAOAiH9z+kLHx
P69JY6vf+lqHSrwome4ObrD10+gM4I5Rh5+nnyLIkILyoGupgJCzIBwFxA8y
hC1mi16/k6b+VP5zempLWlEGo8Q09FRmmCHTEn66pR8JWgl5nI2rmz10oeWL
YqedRBYb8JtA9ZzBLWQZSdLAqa9Kg8zoZzjZyc8eiRD+jhS0l9jzxKdYjay8
9ENmngBfCt9s+vqtlMIuvxphh8Nh41MgA1lCWzF5TS46j9sPWQeM59SoIpsu
JdVqZfcXtG8CKXY4Kknpo9i6T27EazfHgPhKQ58m+O3t6/M8Vgpkz+oIMMEj
xAmQ1y17upCaIq1vywBwTsDA4eCgZMrXtdD7tev5gXaqfNpO5wJDs44EFexJ
KKGOl3rtGACYTHnultKHWCFJBQSPNMn1KWSrPVaEcsZKIHhYgfpGYWtC5Lr5
yrNsN3n21FImF4xd/hVDGFe+5CIOwfMnNAQKbzkqCKx2ekb44lx/mmzFdAt2
QcWak/JvjfdgHMFhPNuChuCVG0yPXZKBjuCwOn57vGlbftWdVieXZ8b3k2Um
/5ZGrkBqCNHOd4M6jPENQWvrYmGx8x01otYhxz9aWzs8hYIqGblKzSOqW9Wv
G/ciNp66I8VwnyzPP9lukYq7U3H9PTrSfL0XqsrLojEz4424q4jZ6j3s6iZp
ExXZW+/ZGq153qwJDvymEiOFWm2A4xKUvx10ezcB3J1aKt62hSdykVFPHFl5
/DVNidgvofR6vfwXgWopeni9y/PApvrFITSSDJvWu8tVy8IqJOeSoU9aodDA
VrS4x86WuKCHrC5Gk2R2rKyT8mepbzrVUFrTuLFGZZdr+geyeQtj4LNu3BnD
co1ZP9AEvIyzMESgUIWksZ8eM10YGnjXDaHrlH/isHPHgOIwE17sUln+DRl+
v4UEwMPnan3nprYZOKImvOe/CdH+r5SqR0m+zX5zwp8jjJgV0kqL1iSrQCFk
WxBOvmjNGg0BBkdJ6FXvKqhn971iW5EIqI7TdvyGHyEmMbpuoFnBZD6IPoHp
F7H9scUF4+LMro4oDZns8rbbxY9VXGm1XbpUjF/wKe3gQxx7w2LyCaih+4eb
DEAOvkxRcF44RTb1qUD0QABYdciGqmO3odlyNwdIXZe4Zb8mLqx4NXqyCpvS
+5RLlogWQsaIXlCGNW8c8TM9FVss44u/2+NLvSV/XtSkmNnQiKTetzLDUl3e
ikgYPlNftx9O4TiyCsf+ENGuP2epyFbI+WzYDHrNTuY/jnL4w10KJHmv/pmm
OdL67y/6qb2gndh5kTHOfY2ZVkF8v3t9DoSzo4cMGwnm4K6tpmsD/x3nJzBH
dGPjd0q4oCvjzdewiGgdut6AgEwLG0eohpxgbp76Dp0PI6K20P710JA3IBw2
//dGvzdC3tuv3Vvk1TsDNmEIyP8L0EKusj3TScFsboWnbEy7S4Yr3tfV7Zl8
YLiuuSEnGsjGJGClaMKao3I6LotYCulSKb3DbXR/kxKYUemAzywrn8sEMtPU
N9PbqaF692oIAQw04pF3MvfinGPrhEAUX/SiGmQnEIgA5v0O5Sgh4+p7/I8s
U6paXsd0NoWHpG+Iz9pqDSPdpduOB1Ld+4Zp1cZCv+//Qk1e46rAXd0D1JiG
FHo4v5SMB1EN9SaXsoMA1/jzPjgqqjqv04ls2zNSggb0dzHopzymdBx6Mziq
mGbhOMAM5HvO3OrB3UX80JxkAy1D8fssftW2G7+No3c4G/KcGEogn6Tn5FVo
IO4tHjA35v7e0G76Lf9YIU0R3SOxNUicA73wmjF2eH30zpm6d4moGd4URfEK
LNGu8lmVveXLnuJLYPUqX03vXRETQ77duBcQVYHdUVfYeSIL1MUHKpelPLYf
CAHp1b6gW4Vx6iX98RKcS6BFZzG8kJI/78X7yPpCZQrr0V7Ws7RU2xnnO3/r
os/3+kq2tCnEslhhnPqPMDQ+7cXKbuZXTM56SWvOCyCdiHxvCr8aHoazb5GW
M0lz0BoeWPFXE65Uy/ZMdCxm67TQQ+hwouOveiD5F1rV2G3mmZzfonwFgfVe
hcI/J435LFSDr59tnuBIf4M+YDVDF3haby8TYQeI7NbI4J1WOzyjoXrvLp1i
bJog63xEocjGQHEUq2ySZnzd5Y0S7pMqNJ9EJFMKIXtzxlY2VlDpxIpT3UrF
ZSNHJuyFrFbfEMp4ItvcHigveZxRqdBotP1CC2136blIBAgqjWCTzIYtptF+
7aoBsqv2R3bmH2FDXoTC/eya2QkUdKtLb1UAt1d9whXxcb/K94yAD4eYYG+0
uCSAvzdDjVMbmxsGPG08ENZ+B+EmwzZI84BuFubrIm36g/kMlgAXIc6n1/BY
uoRCSOxu53kwxpmqMDEnP0IvoQrewxfQ7G/eYEcSWjgLOVzVq4a1mZz55Mrt
/+gDoMSxafYuRKuCnIGUz1svkQnwt4sXRNX0DF4s9bNI3ap59ppzdV/FmtzM
Syubf/AmfpM6vc1gnuCqjLVoKVmIFSO92lgCZvhSqTxsc+I+eIffhfhz4TCw
L2sAG+geemwisdHs9l/SPAdrj1dGMaaC2pbif8lGy2aZYCVUw3lxcNH78/tp
x6ZIkG9M/ZAhthW35ji5KnS2MtTDeMOaqGiI8eD02vCiJMCXlsFAx8bd+mdE
lsU++tNwt4GKQNvidZiv/Fxar2mkKOXTlnItvj1pvWCoOJ1soZarE2AXWnQy
G1MTsqhljjyLmTjkpwio4VzQ25ijM5BREiJ4Rk/BT9YVXQFTHWwK6zuPh2is
xEE7FNIYcFLFCUEbpktBQdEcyocnmsUjmyNziafEZPwWaY/m9wKklk2AHo8O
iLOJ9RbvM+MYD6b+Wqx4avE4/KHzNcF+Yvtwwfuo4abjr5TnmKd/HDc8nd5W
ZF2sG82vreViSDaEe3XeKWjvVCA5V6M2uaHQtlUmA96HQhG6JGs0VAqed9wk
xPPkY+npvC4kQfAOR7i76irtuijrmbsgVUEWjBWHfz4kFqcRlPv5APK+Rh9O
7lTjvZTGFlJkG34sXKgdj5N1cTasUBmzQxFPuAyNirOdNCr9cgJpzNkfiGPo
BJeCQJqvYjJyB8kXY1gDOIptQs47Ve48NhkSbN7uItZhGUTnoj8loc8MITt+
9AZ4RtAlgQikWOSvpW2175/MQc4yRDibpmI9+mrPldb6qKJWAqy/LyBxm3bG
V1+syVm7ov3EwZ5VvlYu5RYD8w/pcCbvPcDY+q8RzWJzJI67bXcqscAjzsHm
88QOdslmXWM9cn9HPPl5Ukwe2Ndzg228O4mRX3bCwY1oWAtWkWFKcwh6p4e2
SkFc4uguWmlV9twW08o+OTdAmzT4mxePM1i9u3DKv7puwNFTSdJHA3cmPipM
1BjiW5u86GGBPo1XUtgCwy9qB5NBkvbEvDP3YpAS6xRj4jAFQfW5GhxQGqUA
FtNVfpxO+0xDDAEyN0haCFuWEyio8ckfuJmhkaEGbacv5/GyU/sgLU08xE4U
bK7wgdsYrIUU6KWT5nehxLnki0BPn0RPDAExm/8v14c36A9A1oCTEdaWGEmk
o2gEXIT92nBxmL1Th3xHiihb+7PYzBnX0L7X9uJ5zNo5VoX7kyX/SKWOPA+j
Jt2J0PqJWYe1rstnblstnOr+Dk/BRmynoULtI7lxTZj4vTNpQsT370QEtVew
La6FR+YqA84L/QXzkMSEQjO41m+qdij22wawhJnG1mrQN5zT2FPy9no3TWw/
ahyoSrVz3j2lPh9RyqsO9an9bMvExbWCBzHNdTf6ZYW0xdVY4RKWieFJCfgS
pdCBawb+mk6xJas61noNsKBHhARSEhlVPaKj/+4NNHF1eZgUEX8sWwaCXhon
tPGYfiEHHfS/Y3Bb/cziurTXDHh2wrQLrncEPQ9prbQ6xHzs4Bq40bjuc8jq
sQ/3BKa/6Hq/szhjV/2X1cRO3npVIu9mWQpy1HkPTpGqe//cS8kB3eFmZCmE
pUgD8WKtsNIX4SWP22cGd3XUsnw3/qzkfuwNMwWDH1JU8PKDfj7FBgFhubAO
H+NFI5TELlXg0QPJeg6ak/0ItkeZrSU92+jKKbtztN9sP1IRqku9TjbNLFrI
vA/ZlFukTdCrnF0fprrBQzGkLOgPiwnQC1xLcu3E8CVjHbOR0eUcJm/jvAvU
k6LpqfyWKLgADVmTJBwlHnsmXxmpKf3J1uY6fSj4yGy1comci925w7M9E0iK
YV5ON+lizM56k6fhInmcEKwhIFWCEBj34qiO2E19rTthuKe6LiOnZvS/+RDC
09/6tilh9e2tO39Iz2gB/XGjsMwpwJp0kUpKPiNL3v2GvcpJeOnmADyTgYKn
5AkqVJuvfNpUhWnI+uHhgs9I6l5zMosoWifJI/t626zpnc+ygJz+BFtblgHq
8yd5x53380JYIJ2DHjHoE1FEye4NrMP8jUDqlvtG1jDtYnFndq+tHv4moeGS
hbwhG0oV7LPGiDkAGdvsFBK/Vaqh+VAd0iVIPnZN/wFAxqyPkawBbFHYPT7f
cBvYEWqUJeNfr4M1WBBGtRnSn8YpCeejuHJCEKxx8doDThj/4s3On8qrQ9I3
EMCb+KzUoIvzD/fxoYZT4zmfQPhsNI9SnLh8DYrmDUBSGKFrD9yw7nxQwYG1
jQzu33nFWpJoKzxFxTK8opLJSDoWUb76t+WCRwMBrU2l2HNmIwYX5L1lc/7Q
c2TUfSFDNLBFUmaIAQ6/zZX7n9brYEGqzikizEwbzQDFOxvmUv/OCYey1TgE
1cPzc4tdzm07iFMq1x1ppMC9M1k9jxuQSC+2+mIELaLgdmJGzS8sIrFviHbO
L0KznWn/XSGOyXO+RL1RVmIKVxRbYZLF0WinrFXaXX9M/951k7UmikueP6XN
FfzYEvzozHT1QnJ76knim8fKyPRuDIzcQ600A+J64vw7Lnt8DIVe4AoQ3iLY
oZcx1MbXzBoXyc2ikifx1Bv40XBHdFC8h81NiP7TxDhZvRQtGqFgyrmsmQHN
KQcJBFzxVMih9nqq3blVL4+ZqAZIQa5wsditIGvxjtF13iXtjK0GCIKbCGAt
88eQLzCQFrWpoabhgQvIGivKJI2HmBgoJ3SMc4d08weKNJeg1cCRkS7iPcIE
afyPXgAFwiW4mE79hWS+Nivc1fgY8rqi5H1drNdXEoBYin2WkgD/0i8U4BwV
fX5sKDrW73tq0/M1T78BgPxfgN9s9NDo5nZXTLQzXZwU1O610rmPDpTMfo34
/0wK0La4esuELad430s+BsQVF299sN+SriV6Nd73amcctb4zmsvLbmE1CkPW
AYdqS/1axZjyl+shY+fMUEIZGeXqgSv7A+4PsY0+WDCULNxGGH69EBWn+0ex
y/79cKUTm7RFTdzXgevfKRJb8WE59BHbnT8sqA723T61nrCtBUaigny6P+Hk
oeuzap+pdgVVaGQr7yutnpOre6DQDMB9jSZBYyyz2EWrLCncR6oziJ/oO9l/
2WtHH6uBXf51liGylBP0np7OWubl0ibwq/ARzgCf4ZRbauFz6h2PWBp0TJAe
wEv2k+GA6La7KF7lg9y9LdRtEYtEBSfU8aFJ+GbjC42QjC1a0+3rj7yFH8bU
OUJBFK/Cu6NAatPMko5H2eS4YYDSwZuLdm1+fsI34J7LsxU9rGWZ9DlCjic7
2TmmFlz9enr4xwYIf6P1yXHzL6hR7PhBHPJFztbSOkWftCGjILJpsHtAsPGI
EKzphlUylWghe3tSrtTc0vrhhZ9Z4JJYXh1Xc9A/Fp9vegaxJjwgrLv81P++
nrG9rJ22e+a5CEfgbKWNHbbzDjuldLzeL+1l+BgmP7HlRxz3bL5ClJvYQJQG
45OUWK/NtuMT52MHySPJXQ6VTChnbHIVwpLjsZgypJ0pk+5Bet/kjTrlUCj5
yb56uLN7SetY84gwejAXS+urgcBZoP+5AMLmH6UchLxH4gN2ZCgtNe7bi0qx
I+eZCXCD7sPYJquJ0f05hKiSpYlBPiJYwDnA+8dG9ItsOfdNjrGQIceaJT6t
9geQFdpC61ofuqP+XSPOw4Ta8k9KCfxG/k8v+tB+4bWXLOP4RxvvaUv/rMWj
pn0eVMWTQwOJfn8S6QuGSMFeLcjJVg8Uehrk8FwVGxWWmVh+rAYgYvkX/Fyz
PSgUA4V/nc5x0Uak1APw+0oicmzmOeCKt6i1/4tTCg7ICh5Xdw/P1qSo5p8y
G+HmsUbY9KKbu1/PDZdsjvD/hWhTLKhRn8s9e9PWNRtHRr8Ggr8MbXXX4WsC
NYdzhKdS3rqzdJ0/ifPpeIBa1vU8ukOiCy0NPBvCw7xQWWTYA6mGUSUaHdE5
jRDzYDUmWEIi/K8QjpDs4PYhdIiE1pXf3Ou+oxyNJpsiWvjXj/eGyoW8PWqK
MzqGe2TwQufTaHEmJULczQ5Fa418xW0hck0DtJwJMmW9tmBlUTJ6+qZS/cfK
HP+WB2CDi+oOF7PS6qBGuL8evX/2BrNneHnwZdEgqiiZkRaF3IulqxxCcKCk
zXgQUmbJHYjJ6D/wmyhmzvV0RZD+Iopn5zbc4nWGp009y7huKHy9uaBzIkic
ppNm0s1qgEQlE4T0lpxS01AjgsBohn+7366N2f9C3HHepsbSiWq/Ih/idVwD
hJLD60iq0+l5uISixQBTM3fzuiq/p6j3noYQ90gP3yfbI23Yx/tU2r0Ueeb5
6I/qCVnEqrFo3VVz3n1tzx6JipjZ8Hx2KK4bqhwXmDnpoqxcY6WPNw6vxNKR
R/HJfobKdiLd9mVDw7ir240DLkMZmguHM2Hf0+dUAfJU0Nznhiwa2Xkuvst3
WYuhyd5j6+4SRjuEb4z1xHlbENa6f/J7nEH32hJJgQaNQL+r+FXlnNEelaps
HpMqLfCZPCWYvwrLiORlEdMlzsGbNMPLnBiRuMTz6GCyMrQGkR7UzeYfRzpV
HjipVK1rPjTndqSSGBDkOO4nWQQFYTI+I5bx0MpcaS3SLKN/hfEJDZ9es9ae
GwlEVTBrlG5FxfATqzu+0nh5lAqzBJDXXT/GgrYA2qiYfqYowoQnK9ScDkCI
AnSgSaIGtVNBT9d05uHUIBldxV3XzJcCDRRYiVJtlONmOyU3z3tTYt8MDJKi
w03wockyyztO0hiEeSaKy0F0AAWJZDO45sFkqGaQb5XcgS+k6Z8zo9xt76wx
+Tb3ebVUvpybEADbkvTbb3HeYNSACClFx+41Z0Er2vMs9y/KlHd+rKRRThVR
/GjzT3UzenXJJOtKEcZjImb2ohPqI/oOsH2DD+YJ2ZZIG/W0wE9a7YS38Edy
mqNHtJZWLz9GoTkMBjMlWQkCTCUajwNRo4kjtCTDaebH1wU4pXCMj7Uf3dLt
ra9ykIe+iX9agEGuM1coMqGawK7Reng6FpuBW5wwcwPEC7OV1L1TSmM8HRvf
PlCZUV9vjgcGvBW8gO22TPqUPMgt6gcfVfFGnIW2llj22V/NwE0ecK0UpbVZ
bNcR+nUGahjxSuDvq0yl0dYXT8ma9y1e60M3OxfhvGEIpHG57JHvj6IBb1I7
hoyJG9aI1dPZUhUf1d3uT3GwLaOIpTOsd+JRJaaHVIXUvE2cISAa5yC/0+n2
xpRC4v0iciq36FSZTBfmskkTN08IcSpELsZTYtFfbNmaFgLu4kQnK6BW7sIC
xq33BzYY4Y7kYPHRDk8XbiZT2rcCxqY1opjhCIcqAuNj2IMY//+yv60qCQz3
IUmqy2r8VizI0wq8kC4+UNLq4w9PnCDniZkYcgHG0UDY8INnI8VtSBhFGZQ5
Wt/xiB+ya1XdKTMMZtSDfyuxXnPmTNgH9+j9mr16uz75VPbnRvgMLpc2wtXH
LKPhVppZYQ8kqB014/oM+FNvCmBlaRyCWW0s+zM3tledvp9k3QScYXshEwTB
A3amHZt4MOuauZBF22K1uO2kLiC6G8KaKZW8+DUBe3lBPSVZQuacrBJcVO+t
5NBi8/qAxaMTlna6iLESoKchy/AVcQCWhGiP38hn8t7I28pMzkSZzebYLEtX
vrBhmmYd37R/Xb6qM740Iu4qKa8cTb8UGiQtZvzmYOZmlbPTZ28skxpiG8H2
dqUhbIVpY0HeRlf3lU4/gf8MkTU0qrFQPk2ktf8u3km77oMqyFHYrUlD9rfy
BBZA0GGRX1txy3zNEpRVCIrrxBs5jvXPjiNixLyueNl9ChZHQAYdY3qkyX7E
dvZa9fBFi2mVp2mt8/YvzOPQhxtq2SSCQcWV+noeF9fAm/Q6ZE11Ke5FItla
89xMz56EcTzMbxoPMiJH0fO+RgUDWEbpQKWE+sBF4dUvZO2XaUgoTOr22CIl
2L4OOJ4J4WMXYPQZUBgantdzd56yaVSdXqZUKXUbZJhDWmyolWZmJc4aFKdc
LzU47CEMzvP/Ql+4CqoAM/5Ulpp8zcXSgV2ko8E81Ztf+C4bcPGwHB7JehXf
rKgzYumOkQNWJEmh54RzlR4bYJWZZwtqpEe/A9Zo9AiNV1AiR1T+yUjtMp0A
iZRijCTWcSMSJ6eMYDC3B0X3lxQ8aYXf2kw0cofnbp2nG066JujRAE0okYEc
fre+KyTiQzez5+VXKMErJJm5BN3A6z9cnhOBnKanUqP87hil7CuR9W8Gh+s6
u00J0euNr41PR30YK5fGczhju0lLWvpQZs9ui0kWCU46wxYXI2im4UicpQRU
LuXCQ6O12f5N7MA/zeUBTRFfUDA8l+PrehvnhwnRcQjxPW9h8FMTXP04UlHZ
Kx6+1d8akCOLsXTJ8KXNUxXitAEK8ZMFYE9Lr0NB0TFWckC3SKAlNaiCTH0M
33UIm6hS/ca1+1WEy+URmZptfgpFwuqM/5xLq1skk9KmQoaAiNUJKblnutLN
6SCj86I/Wa8MBOflfKaDgEYlruQipJ2h6716msWjhsXfQw7Ad+d8Ye+k4snb
MNOb0x0EUfa9BXg8x4Px7CNSiwJnAmKZM65tgOYxyYmnsKzDR5iV4mRJ/r83
BLqJrx9BG8tbB3gLKYqGqYu+CfVtJq5EMiqhpSZrBpexsmYrKDS2vr5Z3FQt
BxkuNg88rW9qAglk+cIkwCpq/89a7KetHX4yjAM1TjHzizthK9T86NfOOFmq
XCwpyrXbAUCVPM3duAsNGG/XyMSX9tr5UukAaSyFGCJgy26dve3hTtY5uSiU
eq//AN+Zw95uVL3S0o9YcMJVzqR6Ts8/4FSjVfr3W1adMpHyr8uF8DfJIsMR
UrhIS1Uv4WYjgh2RxE8EKGvozm9mG+ObwAWjaJFosg+dxlcrTOPF9oNhOyEC
FQxEfSUFS3Uu1Etrij0dxoodGdXd6QYQX8CEGnFR+dtXT8/KXraJQ+Nfr7I7
VH3Nh8BawhiQoy6hVQC7CRq2VKvLfqqEQx+bnWp0JRPrTsOAHino5C2hBGrq
J9fZ1UPmK+AQAOzVYTfdaYJ4pVCAaJZzKKj8fsw8YFiVuAGkfSdZSWylrklu
O3s0NwZBCcNcBt7Iw3s5Y7NLZ5exeootsjbfEQnYYgpn0tPl6/srOdUyaMXU
HqSZ6hD/c9YZaDgr+4InTFASgd5MQRqhv+YiCZ3JJdDfoscsa5ViQH+4p2Kx
tQ8lrL2huXXyZ40OOh6/J1TOpmyzyRmlRgfxzbHu7x6lv3ZsG7TTmlYmCXTR
Vnjljuhj9nuwV8cXrhjY9ycVKSwIL/ow2R/mZvYpEqBgKUFkg6BrLYwJoTzK
CsYGoZ4vJ51Sy4WTEO2pKCMspdnINSmMJYyT6O6WM6mWGNDzo8+ipgffFN3s
iyDj57SOLQJl5mpoQ306lUky+lqXMFBOX8eqAI1xOMe2VXEWuLdt5Gnd6O9R
Ro6qERSu8dQ2wRETqUW/jA1ZS6J2HqlL1BXM0LZYuRIQiIkj7KE3W6OmdQWq
fA6iOG3CzDsCCeAvBOFkr0DG1MSv6zxoAa+UwnMMXqN8rgUfg65VxY33Md+k
kcAlDVOEqVkjmVe3Pg0OjfpPQwcNATY/2uLNzf0xoWYhoC8gzi+SrBLd3R4F
VQC+gmJxH+G3MHHeCE679XsJhuX1v73GEvJD5sEdQ2z3eCI9kzEOv/NPqUMj
4iCBsgjelyECDVIdbv9MGVnJ7LN62dr9B8qiD8GfR790j4xWNriVy/MJ/Xe/
1yHb2jPVAfo10F8kXc7BvpwOg+hhUTRy4W9Yd0ODozb426xKq38l2rRRA43b
XykPYcwGBA/cWpdRdrdaMsXzoJIsgfIt+ECOzrCW3KINJNxScG+MWnwYCA1o
VnUDvORUiaUSZoHELE02t/gshjpl0A69DqjhnZ7ZhiyyDbMIdIeFbAlMWtbX
uWeJmUbyFvLL8y6iFXUiblLlxbocEq59809zIwvjMKARyKrjl/Xp/ZUscuv5
V7YsGNHgWKb6nC9XRlFcEmMzM1FXTp5JDjZ0tMYHi79Pt6hMMwoUzb9SmRTh
ds/HKFe2Mxow3dG687tn0fF85CwQWg5PsvuZE4TIrtlTCnZAceS3ruYhgPzl
+0sR7CTK2dWPX0VJi2SqbFgP4rFwUam6Ar7YXK1bwGbMbdQNfgFygu+9hup0
LBZ5SsazenMd867MY542sAzDiK9jtlZO2SVPhqJ3sKo6VV4s8YXRiEgIsAxM
q7cWgbSPxhDB32/BWWGmnhPXVAYlEaW0gn5tkvRWheM7lrA2iRbPLeuwEDSB
JoMazNdtd0lKiWhnGoZHPqqyy72AdrrWXpOPquVCdRu7DhPu1BKO96PbNz0b
+eQcky8pFyaZNQ2MHCmz3joIiMFMG6RSPQakc/B4RtNNuYGHRIgrTX1VQROW
zC6kSegOtBEZW2yxjw8ClnR4QgBmds6h4vrS4hG4IHjJtVKTX3OfDhONkYnH
151arObxbtdhWaeibJQlfLc9dhHtL7pli6ev/afgF0lAOrEE2/zmZbHg+9e8
fXXqr7wwT57YbObJGJAg/cVbdlEDSpLrBLPIft3kc+gvhz2BP8ezTa4/VgjT
lQxwMY4KEqDzfFEwr1+b9NeFZm/UvS2SQDqNgbfz7WSVVmNaNecFX36bk+Io
mBd+e3e7+Or6P2lkrcpfOW+0y6QLxHSnQrAm7y21VxAlbkK6EtRPEnI4ZqMh
N5f+pw6DNuhpZ4Ti+07Aj/Hw/TFXxFNVTJNqV9qS4YjJykA3o0eqZRDy8aEh
mzSQcHke/i2PcYgQSAHyhNKHcEwUhVdCpt5WIz/PtfXVOIl/Fp4pcQS3FQjo
Ah61o+J4+ZND0+gcClF4KzMW2n0c6F+02bVDvgzJO1B1RYK+mZHFG+8bZ0j2
CrlLUZfubOmlUTzueUEuUZyPPQo7CFpBd+RQhLhzUj9IX2E9oQSJng63Tr9U
4jsE2nafnBrpwEz3eejwqV1e0qvHuCLHLxKbBUchbZVqsvq8CiogTmCfXrrk
t3qMgX1wyfnf78cGKdzpAI4fPjcDbIQWXZRcRVul5CL6Ab5mmGVbP1KO1S3s
eN18QY1wpsxotNClPOtnOUlDcs93X7Zq4qRdjQWL1WWK1fnMrTLHbXPEJPwq
uDcq2EtReno/H79ymtzvF6Ay+VRJa5bA6zFY2nQHVmj7d0VS5kDutt7Rwp0U
m8koPzfVBNu/TKi7KukfDCmTr/SjWHG6mSvjU0qx/bzpKP1T4PjWnXY9z+g7
zUwxwUFOa7AjVQu2h4twdo5UcSBfs6u2CGFfrdPWKOSMPRZutFWulKt9JEmP
USslQKWcqpswtbzingpHouxe2xakEw0VXtZWfqiQmi1XHNSw+Is4glHGZKzW
kHVVQzJS/TD0bfUpKiv40s5kAlOJHgwnqjvJDDaAql5Wz2ibHjCfO6cZa78a
3i03ZTgoq1GqLiq/oSab8hWXitC5hswh34cE99YuXQEa5axPqb0R4uKLjlfC
ZY+eQ2IBbHr45yGA1mLL1AmK+SHKjhtrV9ihNA8ukTy1ziym6d0/9CdT4Bb0
RekYrH0sfzdEnAeYdoExiXpvCtRYqnu7KYxGYr+dOC/qY9VPAmst33yt25kA
lqWQ0/gV2YY9leFz+3I4Asm6fN0pwM1sHEhLDhB9jLqpOi81tXtg54Mf/TrH
3ZP3YxYpgnUSzKq4zRnYdISlFPrT/EHNLpQsAbxXnWrVPrhqgMiF5tS3CU0Z
yMSQqLpCO0sSMgYlgJCsG8N8H5LbSTAYxz5KGzgCQvyCKnmYNmmzkgYzNJSj
oSyOVJ6KwnAGC/rfa6GuAVdDVbJXBPw3P8p8sNaG9hVZbb1TJ86T5M6WASFH
pooCBkY4efZGL4DyfESW/h/kqJv1ykZ0BgOjUXKgBPnm2jR4/kXZ+jYbart3
Rtvk+8IYOvVSli1XBqofbPg4L6rpLgBX/yvFiHHoBxfhwLQ9bZhUDFiIE/Gb
o95IWkKG27Tag88Onn/yX2n7afAu8HOWRorpv72+LC5hFSR6oW/NuwVmoOR2
V9NGMxxB0RWeYdv68e7HZl//L+AsiLRUXG5N1aQi1odRby6C9L+Y+I2WjFqV
Yv8gwd0yz5lJqrUM6CuiGsvNGMp5xNMD3o283++6AzEQwXxXMBSTd+dxKZDp
04XDmIn3eveBf7aobandSMUhyWrQycj8Na0zPGG39sJDhAlTIx4PxVwt0GbF
TzAD3HQksO/8o6+HQvW1rybv/x3h33xDPw22oG43Jo8BJL1lfl/Y8JrGwbhm
3WS3842sfGahqPIBJ0GC5+k+juS+ixHFLXnR4MldGnAOlqXKsRClAKIImrSw
FWmbXaxysGpzLvS2ApBCudCz+iyJ76+KOX1UraIBDcY4Rdf0vIB4iw+vvzNI
kPPzq1YxOGdH2Gti9dsv/fUQmDGKJzxA3bUFM50fl94AGNt5wvgvPAhbngNX
t+XstqeMcA0GjG/80bNd/bGAkmrNkxVm7iWl/xqjBPPMLA6v8Fr3GzYnTneo
l/6lK8Ahdm8HO0EOYq+qs3ot9cIiNDbKqITspC3ahoeMUSRendb33eFtgl5f
8JoQRt6Wb0L2aiTqRCnkqGOQAkRtwTH0M9dGos/pAbxRKcPW1pNB7rUG/+sX
XOHEqGMwGS4D8sqokoi5lKckq5weH0Y7rdoORKNRyrDV9i3tSPasqAFZ9Koc
rj5ZgWEJeFu5NZuIj2z2dnnia0DIct0eatWLkPWHOtAP7vvK7F2Jt6XJ/Zlb
eWLsS1KiF+7OG94vvumhGwvZ8+/UeWHt2GQ4DBgnqjQ+OmbKd+jU2wzbiSsd
FN4nVwrNxD8JpcS379m2LsZSDvKjdfvLFksMQWrtQJdEtfkeWOV+IGpgL6AP
NGw9HeigC6FwZ5jAVSBLtdSyySTJXXwIaeLMHCaswp9SE0J7XB4JWF5zDcQO
U6/dyIPmh/rTEbIvBc8ayY68aZRpZ+j0tD348TRunJlW9FCwgFbrAVzV0M5G
2EnzNU0PFIKos3kBgCe/thCgb2zReAAGs6lwl3QivelKy2/xBAhZg4FeNnaA
Bt7AWeD0HfqAkICjuF3n1RPKIm4FM1nxktqWh/GDMh0G2YqywiVygLkla/2C
mRVnn4KiwgzaDBq7kq8JFYwEdevCXxNZofZeKroMzcof6xbndnTZjBCYXAlX
NDnLorz/jb07Dnyy5cyvuFx3wvdUYCCA8Us26UUGVsjx7KV17IIXsn5HVADf
mQM0n5gf5spv4are1/IRrsGtUfmQZYsCiX51/tB9DxXv92qhMgH8or/6MBkJ
mk4fC3nhpq3Wfkm2ffgGo+QR0oZT8ipAUeqFq6PsoaIiwKPYYebuSiZ6Q6VM
jbuN+n9pOMZN2uE96oqLx6Sx3Do8ODUJvVQQ1avL51ywyIzi/0J9mT3FMPm9
zK7ZhVRGgGOJhcP9G3dJ/nF+yGOW4mNRQc4vPkZiXAd2TqZDQ9qcuU9XUqMP
5imvDaHjDaubUsZLYQHzQ/BqctQLWLAKvmkF9YdUpyNTnevEp0c03fTRSWiR
4PufLgk36btPhUy9awuCrKTSHfQql13HbIMfjZSQiGziqizcXrRhsvztRkIv
+2pkSj+g2XzPbbTt5xR+f0h0U8Lu6oSY7nHoB5AT79kTUIONuofE0QNbeOA8
8wuAVgDk2H5vjesCbP06GK/T/P4iZR9m9LdrYdLAYXprySIlibm0XgRTaxXk
YKgj9V1xslZXnuUgaSPrekdjA6Jc74OBDj51fR1dz3hpRv2/yI+ypahxxAYA
F+g/o+cPyLESYH7V7SOIcZkktl0AgCmC9ID2/jYLo/3Cl7MBR9DKLfTcmEtq
atmCbT2AYnohGWYjecToluK2SF6DqnTyf0DWtftr2sfDm2kvoRp+5G6laVg0
vcQxY7Y5sfXBIV9f92i8QiQI/VQm7eQFNWk/iVO+vnDYHSZBkNCJWiB52UDM
/p4R2/vyBHwhbQ5uypwAPj9JHmVWokJi3JZ4HeT7txvJTebXRRuReOopkiW6
OmEfvMeqDQjGrgxFRhcoYQJbbP5SsBXRYth1LS8qJM8bKd1i1iWTtm4I/KTP
l2ldnDmRFctjwbXATJe+j2IuG8O/JWZfLvPYxjxED9XQNbGDnzMWYO+Nr+N8
c4RXCyvnsk+e4k6grZm/I/zP3inEBluXeLGC/XdLNI+dzW4YkzIW9FkzRAv6
PQS+1AaF/+lOM1ygPWN/VGa7uCfxChP5bn/YbUhVptpdX9AvrZCbF2xtj3tb
crQndCO0yWOgmnVBy5bnkUpRW/7hElvETPCih7wPbXBufeFKajXPrxcGFlS/
N5D7Sb4ip1MS9KBaVVecwbeiwp8u01VtYx/EInelPKeL0ukXzkYBCs6vGbt1
3vN19FfnnkqBpzmAndPqx5jYiOZS556NI7VYyu+ILFBxhlyZW/5qHqQPlT9y
NVDq6hZ7fCuYsUrxXHITtbKj7I8pnyfH3CPqM3W9Q/0gF13N1xBCUk1lH2/y
7W98aY46TKiNFblLFLSDsC8hcxMxb8EvbePODCQDO2Pizzcqmil56TY0G6mi
E6UEmsBsVYkEDsrdk85ypKV2uSBt0cvYFFbVYG2sijZ2qVC2YdIvSM5Yeh8u
uSpNJLUk9OK0zvNXcfxYFdPDhMaHWzF0zsjMshmGxFUe+ZPjRwxxZ8B+oBpQ
cBEv8p5M4Wn4WemCedvf/K/88+Ou+A32v9vidouLxqalnCKUuoOg+4R79IKY
sOdC/8lzqTPpelPJQIlk7VVbepxG/UjwsJW0hwwyyv5xGXD+4nNpeoKwd8CV
+tLyvbz06GawxaJyt06auDoaFAZjAKpbNZTD58Utgplam5Nzd3Sa4hwW1UWL
qQekSPvY/Zg26c2U0cKHYllxaLLijI6zJxXVD/xaMNSw/bsIcwpS42WE5Ifm
ppmo2X9KCwg4gtWCldxACgXQ4E2gBJ2XhmFUGdo2I0YPyliADRuG9sS1Fa2E
QxyZFFaUYWZTsz4QZdirTqZWYGMw5yVQMkBenfZ9DG5MR8e1laLlWY+q1so9
/WaDhRF2euMHvHXbZCf/ziojr2qXZ1gsTqI8OXEIqL6qDk3tMmdo6rcAz6Zt
YVunWJRMC9NaZMMWEeVuWrnAoXzD7x81CdBb8dKdyNuSM+1mLGThimlx6Czh
U3kytt67W8kn0u2V8zY+djoJPpzparPY7A+4KFEzei/q0Y89IVu2hTLU4vjU
XNIn0EZSotukK7TBDKfXGnQUduWSefyK6Sf2J6LI5iMMmOuPhAnUCA70ZaAi
7nXbZ9PEzjoN/MzYKjQxVfc7HoekJXAxoAfP8xslMqC1EUk7099olVYY+Cge
yhJvMp6Gf5osNzPuRWSZqbTwm7p/tyctJQggwo37yAokUmUq3DRtThfX4a91
ZIB0dg4MmyCY7yCEV1QG/UbMIfy3wVkOFbnoZze1w6hDONcF0AZsNRo9smnl
faDpLbKgyJcp+snkl+QOmli9/jJs9YziKvZyD7dguXxTHUi42K6Q6f+eN+fS
Z4uLfPy86tgFv054k5ya9RYMoQ83Jmtf3B0T2OOL1o17dVxOm8Xgpk/TFcGw
NdIROZN6FlbdcTENfqWrBmKYfquUk730pvpuJXHeTctgT3gN1AI8hPDSfLpB
mX1UwVqRfJcUa8nNQ2TD72jPUPZgU0OHlhr/y3+VD3t5Ry55rUW2p4FXWOJf
EaKvDT+cgvp1MWDbsXpEDd2yxZzVDdf08KtLTRh+9Du/Lgux29v9jxhSN641
ZXViZAkH6t63zoblXL07Y4+6lw0obR63h6omtOP48U9e3cEn6Y+oakUEht7X
xn+WQ/WxV91Os4Vvd+we2P87w8veuV/sjdgKG0gXCRp9qxruFfbTZtCtPuQw
3A9FH8dFOrAUX8G74D2VilANHLIT0/hMvBTI4yW0GfeZLIIH9d1YfnzeLS5i
WS0Qt0SeGnD54zaEQPg9hfGkG1CuTk/M5NYWpSffa/DnUUZ/Ng6V5iaBcYGc
25WrLXyZ7bYKK6bkTUfUNxT1TYMZV+7Nvc7SeDLultx7n2uUXV2MuTpLepZW
VJ1sqmQO262o9azvi0h6beGw+d9OELA14aFqKs1pirB+52reqRQdLACQk9vP
Mogf+wTqaAgt0E6CSIfmAbEK/vk52FVijNIOCe4kiaxedAO3svHIFaWwh+a8
erzqyknq1KRAS+sBcVPC/02CgM4GJzAryNSDoDtmoC9D/RUI5PsnSnOaZ9yw
hThir89JkZfUgsRcYMw1IVg33O70Ga8TiKpjgATxNZEqUlktUKLdqazl2ScU
dEM6+tLJey3kLBrOBkQR6NfR5hzGHWRW9P+ekMkV/h7ognOw953pNJx5Alb0
N1cMsQdgkv3mfhwwHKIDe4zPc46AvB5P6IcP3Ny92SqrWf6xsGXbhwCu1DXn
nLdiWb1qHYmQVBlGvNQACKnnt0bRheaGD71iJNjDimoflnuAnjdI6pV1CGQx
lCzTgwAUsaBJwfic/07K3d+SiRf+zm5/am4OHBdoSZcmSoArbFg37/y2QkYg
sI0f2UkMCEGEHpxkbGrPaa7X/Sl+2VH8DcwQiDI0zUi4foF6zX5iXrEI79Uh
OQquWGZT5MGVfJWslFLhCjQOcoCE5GXuvxPcOLsnGErgf2UQ4OPoWkksrRyV
SFAkDMLhr+RgONzcQWmyskD0AVEsqDcN9IQZcLwSP4LCZ55lU9cEDffd86O7
yQkudehKvGxJKT2FfKBBq6l6+TRUGpDj5aLuLGEE/pnULku1BjsNonw15O6H
QYWkD8GZI1wzoDJIeLQ57d8D1wmj7goXmsqZB08uCvVkoJylZhA3IuYikvrk
imUO7xy/MB0xZwSdSvNPMqHppkp/IjaEx4weE6jJBwgeTqi9LNNjsiLhLYqA
9XCgx2NpbHyJKubEGRBLhdQymGl+helllFJicl6j9626UHdoK2t7bzJ/53wW
kAR4BmMQPEnWM+wR21CoQcz+bADfameLyMIjq3G/8yWYUoZX8797PzjQEK89
nP2NaK8eRT4PvyI3sgzO4tutAIQWjrH+I1KCFG6T2JWrt67fpNqCp4LBq7M3
VjabA9+g9OBTg74IpXoo1fqnfXsGixRNQMe3gca4Vrrfs+P4Kn4DZZeVpOQ9
r8E415zwXOzF3X33knKP9G4Sa3NFY8HLx6UatMItWOPJjmKsm2blUNbHhGhN
mTg8G+n/rOE0QB4uUVTlmmKlhqBJZQTIqdwozNYTz8N9gROZZ6kmC1bdph+V
GNWB4JBvMcLfUp0m9xSc2+NL8Nbt2hBuSBGWhUcPCOPtxqYbJVoz4oNEeDrZ
AbNhI8LfsMkcUMgw4Is/nlMxyvExGjxIdLXZs1qd0WNp5jLo5VatgjP0a11S
lIR4ORf3yuj3Md6zdhTwQ8QHr4QFqcbhXQ++hvJcnoVNqeiAUhA8+LruzTv1
f2rn4E5EZm29UfNm3rNotKSk8Q5h1ZDv54wsZ447YtxH6XGQxYxjtgBAO2Ol
GT30b11MqyysH+L9ScGYT+g4H4x4k2XgVVL6z6zkRApHgjT+BRH5qdw1VccN
6dU8ryYEg7LqM0/mAGO7MgLQka75gkEKJy57OVh+x9TkkbYaVhAslhuAxm5E
qMSMNqyjMSS9YXn8eu3ApINzU8Oq2PyK0pQARKL2gT0Lrm3ptNlHk5UwPZY+
eiLZxtfXnltorDTCsCggRgJMEDLTw5fP2VmNMoUiqK7mR9BMo9BOe5+QDaD7
YrJ0lY5xJMUHEaHeQ1aLNKiQt0oFsslniVTI1a19dMysvYALji/8mGR0T6Bs
coW6uMntBt3xXjyBQkv9AT/JBaEWULJkWivUIIy0yqjUl7X4ATloj3hB0uY4
Er3SZ62Bq6HhkaEK533C73Ai46PoO+9HXvCXYX1FFdDRxNA/70oXiCs1jPl/
RNfQ8a40JvwbWKtiZDWcwp+RQ1yW/1XgRNL/jiXDRGz9kaREMPYv8HqpxkIj
K4j8yPFHYzD+DZUuH+PC+QtFBg2V0csmB5pxC+64pybD4TE+iolZmddvR627
8DUv37O/+VQl8lRraBmBrNNZ/VPErj4FpSvFPE63r80l9XLEROCICewaVAEo
oCTeV4akxfVoECctuqz0/BD2hk1hc8b1MrEiKGytXZWnKHtpZuLG6lNW5WHS
tB75+zn02zO2inx7B1gpHmQQ8o99a/cf5R/Tj68nIjQRUe5e1YRgfOQeg57x
2s4ACN245K6xxh7csfFVj95LaW/RpwsxMQdWvPOkl+h9nQjn6+QbMctiKonZ
NFcaMLfbNlca2fSyBR4itqnfg1mWxhHApxGxJiTVoYOsSAFRu40oKD0+XMSX
/a0BhVoK3OLL+fIMKMInalgpsI6cK4SM4e48i9o9A85PAoZkOoSXbG7F0FF9
5SMILjXoI2kDw6ATT5XG3+0Ck7g1ZiqywpheXrRtPYv4ofJ0W5hGTc2dDGZa
4sbr4v+BlIC29inuNebPEo54b9mBAgCNbnfPHllZy6f+x19osyZmxO/LUZj1
4Q41JWCo874Bt5HLO0oAOLoGD/zuEGb7WJ2JPbvdEcFzfDXInwjjH9wPQE/5
7lWuQNzHlG8xmtbq5LFAiSf6wvWdIPKE1Mg3zcgF1Sm2vp9sJ5ueBlhz1rUL
a2q5RgHBoK9jiuNgnEzwBaDCKFb6bwbAGbG2/7ztmMBFl3y9CCIPEos6rst1
ovjJC7bryOraxA364fvpG8RQxCwKLE7bD1SWU7vO3tMOGzEd8s2QP2ttllpJ
cpLnxvvneHZ682Weh88LlmPeiZyRMlpp3FQRw5CwVDsy8iEqXSIqQD8Per0z
oQRz/UHx2acHZ8ZpJEw3eFtNtX3PX1l26FP1PJOyQ9ETnFHMbG2LeOg2hgFc
QkFzxpPj457EGQSvhAvXjri6mLuS1qGCTebg3qx+PG7Fbi14BnyXhCZpMUJ3
iy0AEjBNXa3TGONgoNYpLzkERlmprOZt0OQyuyLwtSySvQFNcvmI4mYqw6su
SQStdO/FReswR6y7rpACOyRJ+sUhQI35TefG1yZRu57biS0JS3LUJCUBqQq+
qBtPLJjmvMiE9zR7/A3898tBM1D16P4LhszJuLQke+mNT3Kl5Mtl1t9hOAI3
mlRh6rZl0kK2lR7iKT497kOEHeaM19ugG14yeR3BXLaLIwArJ+Vl7E7C6ifJ
OxO1QXED0ziQQ4S/KQGkJXUVJ5nFr2CPLGxH069y6UdB21Q0HjIPgWV673mD
Dan7GoUC5Zrbg3bR/QvS5EkDXrBw3V2nABOMyQHnN9DNJlRJ36grdBzHq9Pa
fhSfzbdjOHRqdY74CjqGsP0RxVqKv8OpuSvvh1l0LkMjaWbRgWG1U2BlMLhJ
vkQ0QerzFZKIMAe8GY1r24DIJuueiJqXkw6c6WU+Lwm7ydI1YNfhUK7qnxk5
mg2/xYPUF5uvjsk0ATrPwRGG4Ejp++wF2HXkc7mp6Anwr7xIDBIHQUrX/lPy
awQmHbDr3XGAkraVSJVFOyg4AsopgOZeMK6yg+fbLTAyrHJXFAxRuMqbl6Q7
GiDXIQ2WcqKnjcUXvkLZzn5/cwam118o6j0y+cha6CR17dmDi+Ay/OFd2Kqj
S47vcrz7NJ7JFhnCpkkkyVM/9JS6yCfbbELpEJaNX7OTSaa2fQ7VNLDHIVW2
m//lVOCf+JF6GyZt7o/Ha3gx/n4KbIxmc6TlkMKFgycjFdbSL8xV0No9ol5C
/Z+f86RnOrud+GhTutvUCh1oVlOzJuyLzZXbOC8F/IiYz9VfbFc8qWDpH4a9
P9Yyni62o+YcijpIt60yHB6bC48QOEqnhYvNJF7te+2IXmosOR5bgEyGewoY
WYIRwCEO0JcJ2ZoRxoXr/7G1C0tHv7FXxlJ371HUuQtF5rlokdavoLnoJBwv
LWhzfFGylLktj0Cg3/dp1g91OubS5eEEbSJGgfgmNBovXT9xayRFAtqWl74o
PLbIHGOTxyA0NosXM1VrDsOKzgtB99O/qLLI8uxFWQetkSasY2mNKr96eLnr
VEYxV3Yb2+oSjL8h5OdDOP99boFw463GdhsZZD+lmC0aOON9WpwSHBBrm1Wi
Kw9XaQdNed0iAqK0MmIKVAl2rU3ZcTjmXdAzNP2KlhiqXwFwb1isRjvIOL/H
VYug03R3cyvUHTR4rG/aogQPiUD1dk4/1pbXi0IXpkeSljcu2hSmAGKtf7KF
IMVitWaEUG3YnH5Y2StJMMpuBoI+FmPfqVXwDdjnY2BKfke+XyGkAMPN03Zu
7rrIotlbeufkO5BpiWhba8akuiFkTYskiD5fKEyfxgpFSBMPNT25ii6Dr3to
rSl0IKuENH30hjY8M6soacuUNTvsEKhQBpKBlCcXnjh5BZ93A2M0wSCZf/qA
wVJliN+b1bxBEFUaCkCuF9BvjA7hWh9NC6J380i5FNzpnsyBnrk8UZp8OXNg
lHYGljcyGro4LQzAp67wiEjGq0csGlkeFwVidhFKJhqLL9NbLpXh8d92zcOw
hwoBUC7IRtWspi5mxalsf89F+aDaQ/1QpBqdmnItjUmFI3J5D5DVs2me8ScT
TFz4zaEh+5qnMDFj1DGwUNJJaHpccLdoSjfbIRVb5GTBlVsK7E2CxW6n6qRD
cl1dpvMGcPOJrfIILAtlTegi3ZZlVIJwE051qIeHi94ZwUd58hepsovZ4SEo
QKKtHuR6njXHS3W7AwhUgkOACDnKo0WO4hNWGI8A7Fqmx9ZqCfurIohqir32
ZAupAm0KIwmS2M56Mda1bY3wl8hVqd0od6UYNz0vf+thMI17YDYNwEbQcIqf
idH1YzMfPK3FMuKrNPIivz1oIWfjvZr6CfTurrYZIZzzwk+LAroxGTw2W9yL
bNa/H14yB02moKxkUsrA8h+UeUsBn5/04NHCO00H/vdKFZEsD4nzavirbpA8
vcs2NkIkzawQ3dgQ87qqna1gxc3Khsfz8eIQn9TE1XFsgx+ugBTZKyHM+D3r
HPsFXAtpwvcsMpv2Zh1qw1YOvpAkc5SE9y3zeRp6lY6n/tk7gawBvB2zKGQk
RiNgLVPAiTUbmoXDSLT9paoj/C5+ykGRVCev6ZeU4lPATh9qHmsGY3bcLmsG
wlFl3p3HgZOk2q0ytvQay1TiasphtvP7fXohFBJmKF+rPLFvRJ+q3DmEgfQJ
KLcaggmLusxMRQh0rH4//ZbXt+YssatbRHMP4QCRbj397cD+6GvEdjK8eoP6
jDrNWZ7VXW5umeu+rngvXimxhepFSmTlO1ySBc/iDIEvGVHqeWT2Y5LzwmhG
7NcfWh/fQAEOcCtaTI0GGZflywbAURGuQz8MDon9Pe6H7jyCZlccoE20oZW/
UpoElfActFAKgmmZW0PYilQzuhvsDggvxQPmNUR/VfTylONVEOwNoyY1/S8C
2xhNRcoX+kYM9umLgEksuUVtIo2lPAHUtTz8Zp3TTt18NdttZ79aT+oJoEyj
V8h1YXj/Xw+rzfeqL+FNhSKXw3paTkqI3aze6uPyUxcFT1H+pogESdJ/BCzS
JnvSyXfXm/26qCl2RDII6M+ZtSmqObu7u2Q7q4wKuXQZG+Gq1Bp/M2tlpIRc
zcd9ewP6YOz2AtD9yoaP+EYiCZ0woqiatYghxU5LK6c07tsj1nlPumne1VRf
v/w150YsoleP8mftvUwQVKOdGxeqcm+bzLehXS+NJWc8zGcrOlyNPVE8rGtS
I5US5kBJMo5N2eJXuSTdj2+4P50Wg/ZTCfuamloqkbpsB7xl2q5MvYBqVi/I
/SFzdumGLXOcUH7X/8ZLQUKntIC3CF1WHgOj76YxApT9Q1ee0PYmujL75diz
P1V39wsBUfP2Re5aqx4VOocugMbGGIREcm0MyUKiUaZSy4LQwswjK7qbvk2a
O8UWwgHWfWz7ThX0NQbOP9dhITxTJK73rNTNLtdi2n2Gqi8dHjo+U5YQ4SHv
0rcv8ArHm2CbbgvEl/gvA64bPFuHOxmG4b5PXU9QOqmF8zyyOa7T7LczmxZs
Vt3rk4idff5gPuYbjDUyExgWtoOw3kUlnliqZlfRmRO759UpfddBDDSPcHRr
ZaKLW1s6Octp3nZc67Mlj0dPH6Mn0KhYWueAc4bvCKry8OOyQ7QOHa9w2sAX
UR7b/MzyIyq9oOwCJU7rXUdPILdUXP/F0q8o7q895Lm6QDiipbrRwIKTUJb8
DXJmK+mNmaMvBzDN6LLvdcffxw/cLwd5CBWpMQh0ynwREEU0dUuTPNO8GrUz
RDFqq4nDtIbbg1iaBdevW0iF4RYinjwyY7q9kXhkQxO4H/7FaLUXxZ6VO/VX
ybhkEkjekGqgtZJ4EciouLSLBuFcDjvzlGAaO3odudONokGRObXpKCW5Jua1
WHplfCN2QyC0nie5eY0IEnycSpDMyoZuQV+H375u7kuuZ8QJ5MIOqZHLiDVy
hJmIPkfJ/f1y5kYXgzneXe2UXv5+qKx8jhBYlZTpsJQTE6kl0xnupxrktPfZ
zKnNJp4PRGL6JPwWrRUp+8l+ixm+GeuKWMtaUdKRx+MPMxe42csXTAAHI4Pc
ZV0NHJ1/8GFBaD9ndNFubBrnwdyR10kcwDJohUv8DIVQ0uZ9OZgyBblJCDbh
Ljo5xR+z1R5x+LrmhIgmWmce4PcSzUOyNtr96a0jVuxtzp3MTA2E4NYoZ/3y
SdHl5EpaHKbwQrZHw/yL304OwrEhRox5pghT+Iec28iXggVhFB2OgcTCzoHk
u3ypmURngUyKZG4MGICP/+euL9jxkWjJl1G/VT+AXho0sAIajhwVKpxT9YjJ
7a9ODMf9aC+shwHwQFm5mtxrR1gj1/lJ0q+07ce+XDQ2hEj5HP2RliCJl1Sc
vD4m0YkP/E1eHGievkY9DJYK7WBpalRxsN1nRGDSwlcYvNr0E0kCZUP/jPpv
fO8VRULB8cyJhz67CL2rWma/MZ4GCZjJvHfBv1tHCAbwvhl29FT8kPdQqltd
eJt2t3LOXGJpYH/eFqKX4IQtfWre3eVf25SjzLobRvjv4R3ZL2tyILS1DI1h
K7dnxz4dwirV0vqaiKsGxLheA2HhPvilk0nd3qj6xRa0xtcCx5utVJSiPcLU
8MMc0Ah0drQJ/4s1VvARvJHnq+fCEDuJS3Sv39XgnkbMXrkwjvAZTLGYY6fe
yFPb8P2DYo6u4txWMdS9UwfVParcnh8p3P35bzq3HmVv6WZnnYN3a6+K48yP
ztfZLFxxn6imVO6mVzlzt315pAk8riyu8tN3Hp84Y/hGfeICgNtgT5pf2ykD
urlx8ONuW80i4qiutik7a9PQ/QrIjPDbuCaNM9cXJipedbo3BJhRQAXBr8MB
SJkTvnlFbRQnGo/vlBtZpixuUf1xXzna44aZOjjl+Cc+gGXDyLcWSfjBK2pX
XP3bKfOfMGF7DQzwZfSu04/8F/oShruxaHvKlXx0bmuoEo4roT2vy+5COa4n
eSsKnsWrRccbFmf3H2Mnv1BAb0m5tH/krEUBUok02gkck2niHnxlHn72/uC/
zlcQsIcUqioNfL1EbgvNvZVC61aID0mMYNVo+wyDpp17ui/sh0g5myCxmhY+
su9nhGmURzJeHlhAvVWVf+yDiKX8Nsfa1f1KyWvDqe1jDIV4kP2ix/+aM/nE
uTmgWqdja/aOPqsQ+5hQ+g91M52qD9aJQHdwNG6RWbSBMDDzE3/1IymeFzF3
vRjHfTVFnSH/BQ60AQv1vJ7y/9bUvc3WeJlsy3rXpExAXXBTrCiG14G0WYKX
WtlI+/F0LL3cGGzlXcuV1dZMGM7TZiuHcobd7NR4Rm3LF4P06K/zMaRXs9wO
hKM0/i7YSQhND8lyVHYJ3SjXu5g4P+l2UOs6QVWxBWx8ee00uIMuuABq5YSS
4J6/FkyIVj7oL1dJw6KGVUa4IKKgbUWYNefGnr5Qslj4O6yV87v+Mg1cbmbW
ymzmgsajQhzPlHJMV3mD04/nQhb6K7qzy5JGJAkK8aC+4Q8yb76NfPNr+L00
9tcucR1AEO+r29CikakLzZ29JwkEAfyph6BWEf55CEvi+izztizegwcN0CxZ
1hkVCMtye3I6rw0+NeNxCrFBMECVc1IPoMlICZSnXMB8dmwHteNRGGhXJs87
FNpB47hgr3+pHTTA22lWopATKVL+9szBA/XtX7ODbJNWSB5zGLuKgUokYryw
lTeCyAYTUbDU3+/fpqZIHkOfCMACnOArFep/aNHGwaYRDAUmf/VBXjjsewmD
BUhG9GDSlfOYGPnliFquW3x/NGalImeHGjMWUXxraBLIt5vri7le61hKwPOn
43LTBUBmGZyTqGkirGSgvqtbaMth7XWBufdcSoVMegFPxWPFy2UViqtxFA82
QCPSrmZm3ixqmsKDZxXkMNXw/m9S5VAx2Qmx+El8sCCj0gjPlvfyTtCydP0j
oQim/5ZzPrquMRJE04w0JzyxoWxZyUpq/AlAXWpDSibMYJ3TEWUNAwhRCkhw
Wg7ouDKzST+YgGVyuEiMeIftgJeHyhXkBmzNVWX/nni/ey20jUDOHOaplf7G
sOyCTuMQjg8FHzw4Yt/4/TuX9QMFSUdU4nkSSlDBmShkvraAkl+oL/pKlYg2
X7FH+/qpiFEuxZ57dgnybjX5ACDNe2o97yIIsFvY/yC5WZo0QUIoTHUCdKwA
eUXpshfx7vwQH8J2TKLqWuQ/eAvF6m8K2jVLoJIQyRDDtXWrNOAwPrvD9MCW
Zo8+0DCJsCnhtdoRL0/fhMi6h2vHUqQnnn+cytw22P5LxGfTGXrZu2zxp6mF
Re2Os6YzY+D6Xy/LpbuJWar6ccRGqwgAwQvo3TO2/VTvVnUK0lg4dVEiHYb8
zdT19aUBskqb4n5amecbzioVCwJ6QhmS4cyPPUZIWDw2XwOa1ePC/ku+Kk9r
Dp0D9+zEruIHL62shgRFJnKOx/3r1stgophg2B4LmHyRbNnawPYsYX/OKFLp
8BSAnc/iBzmwdDYh+Jfvh+jgvxOvO/vHjNEkca9ynVZeNSqeMYYOhwjAaiNa
ZKQMxCUq8F28p9u0c95NweUXjSckXViXMw8fxreLIuc2Eh9yOm1FGfGf3FKV
zWjJ8ngSNnw8SsdGnyU+JJfl0lCWdhLGgE2LEdpyXgG0wibVRv193cTK4YjO
0u7WkBP0NBuSDUQl8AJrRuE6ks2eixrh/K1x3Xp7cEmwuJK+vplCP0PstlWc
DDu1dkr8jo1RJhINab2geEk/iwF1eyypZPZLjFIiLwDjlg4hwaEeOpZScR+8
UYELJmbG7y2y3+Bx2d1/HnFe9HuNz6R7IsSzu21fF1+RipMGMo7mP30QegEJ
N7hH62ZIBoDapot/UsWGYQDiJ2S8PjRy1IcfAkmxe5kexlZ5w1CnDv3+cKVs
tyWsx95XtKRxorAS2P+arryk1ZMTyDircGlIyUnXnfQ9st4jPWfm8sSJqKMC
+3iXXSK+UAUp/u1inq9q8zcQ18PZt4EjVgzH6pVRMJnaJK+SJzICXdg+Z5xp
Z6XNuyDq/cuvR3te/edPLfjrs0HEirIh+fR0Jz/5jScPpeuecIfr2TC96Jei
jG1OSJBKMB2OvRl8g6ltWw73/53IcyxRRJFZsX9wq66IuMDOXZyG34V4hDFd
TSEBp6KHfKDysFaGN0+xb8Zr3HzEFLZB5yTNetDDeJU11OtFjpYmgdV2GAc2
+weMq1YEV5Rq9jy80hixYSVyxd/x6Sk9HftZWFAmz5kRAhdzQKbwEEPTH9Dl
vzc7LLLZdMFhPb0G4qOBy7uGinVIg+cI+mt2cS6URar1Y64nzFdab42aWa2k
7AOR3EDZUCb3UkCRTmZbiQaXW0rNPuTbtGR5/4vA6TmgrLnc9SIONfgI0pNU
VrcFb8jx5uGD9uE30mwCT6ddnd1vOOkAD8FLyzKVxQxGb9fmNLNZ4E6nBPAm
frqjXduuw4qAjINrvRw7izohZXwq1YjQmwJzWsB9OwV8Dq1XJLkDSDRwXLbX
PPXoVRJOn5mcNjxQjd/zPhUiOg3xc11vRGpkwS/138MplfflaE0nmLel1r7e
2g8QnOBv683gCsOAEi0+jaAS/zRJCyVxqx5EuByR80GZiqGEieH5IaE+/LGp
dVtl57guQgs/vKrprkTOpASfBjj1HTgEX0fsVUEAamLGYd/s8NHKAsKNRKVy
tLwMmyI5JTe/q2yzpsizl/1vHBp83SLwU8gG85PKvD1fxZR8oztwDfafl/DK
f9YujT7zkI6/p9AizwgqbgifZXza8OD/w6qhoVk+mkTTrDafvlqYYGsWlOr7
7/rQ14dp2ye59CqvN+68nW1p6PVOKlDe7d3E//ibFZcuJ1TCFsyzwcPMl2+3
Re3fTptrueOtgeg6ZK71seskAj31uvumUzuW9qlo5acXrb/d/GATXKWk0MAA
+kMPoiLfwgPklkyXEACayPXmJXHIiqmOxVclerJRQvN+12iQElxwqPf5iX+H
f6RaAoAJVZSy6DjCmdDBvbGjSbUekupSZCQFcPt1wrgh5kYqUKFp7b2urHMS
CGANqAvTDoFFpGXJMGDdo4z/CLJC4LwhR+fI2bjIBUoYqIDKmW52H/EmIJcV
Dw6s3j91Ae6+HKKt8FhQFopvFhtnD7mUloazBEtGES0O3WAy3CbiKphMBEox
WN8j3zPwBUqm/eWuRoEyZDHyDrz1sLwoGca1DkARGLcKuMVtqtq7rdJ25MBw
riwg+fF4rcHlsblkaNTkXwiizwaZClYWVr0M31kf9hMEVJ1XmfZ/SpyHHN90
6kz1ACiwoLVAoiq2YVb1Y9QInENZoFXAegAMTQEC7/tinUoRyz63eZSbtAvN
Sh69AFDJ1lDrOB3R82ILviOqg5JWB1gAnyohqxc+0FhLgnU/UZ9JEk8MEjtp
LGm5uCYA4AvEdFXfAfYREOD2Ui9jGLGwFs/DwQZor1lnr+TowSEpcT54Wuib
kUafjp8+6BIxMzQkirdc1RrR+ieBqD0LKuJ6ob9ooOqtx1w8DAMfh6oXR+MO
cWsJvgeR6NhJAJMoP0Vk0XWNWWVWFcWxlLdfO0LqMZwgQVb9FJA2FSt7pnSA
Uy6EjBoVfcTBiUsvchrkel9psyhgHwfp0EQRPrMdWEQtEV9SfM8vwQqmXWSe
Xf05jGZyZ243EOv1pnN2vSnEUhXLpUk4+7oHV22ZeNMqA+AUt5RAAoGCaHM/
GULeDmAoFmenU2nqFumhKLUoH298jvcO77gFRM/UQ8zwAMH7H8bHSREV/rMh
zhe4VCXFSoU3oYsbunFyKOAVZ5d+fcVhg9OK5lam1tQwZruEXBKEC93UCKJ/
OnLS34S4xJXaVipE4JRLJKrU2qOSPr461RaHSWdnHmxU7/tNupiZtoW3i0yI
+0UVZTw5Ekgdpod+oS5MF7y8j0QQHk3Ua0gnuZivw3abrCQtm1GKr0I2pUfy
0KMo+uBsdUhBOsGj3TuGPNIq/wDBMt1BHVa5bTggnYf+K8RZKUJ2rXLE1VcV
5uROgL9cBcxe5eVeoVjKpKVWrIqsA7eCmf08gjCrtmMrNtAvngIgEntCgJ++
QunLJD1T4vPKi0jT04iogbJZaKChD8GIqvXjiPflEyKdR7GLaK3iD0BVgcho
2OY1kHUnYR7UJ4g1LHKLvTS/O+AvqnF4X/qtSVqpqO1g8ACOMvpeDb1JeztD
V8eR83NZ/3206hlL46ne0zlpnqckg1jTct0Umw6C7fqRgB/CPSDXN3VcN5oY
hWoFBfugAQTXqe+gaWYmnnHjd242OcHr+PL6caPmYe5HD9g2Q5fBaHvARJtN
rW+VSRwiGbrCtiWP8ziZ1nBBbxivOQ/lse7xqW4OV5GZUywIpCxb6i1EuL9W
pY9pHNPDgoOSxNcnsXMEqE81cZNdSIkh8GyZrTfza6c6O4pycNqxgMjNsHXE
s62Uv1ekkuGD2lEivOtDN9JN8gZep3h8VMMA9bI7K20bnbyCTlke8IKpI6t1
bESvZBUfzeCY7AS0HpWOkEGJCQxL/bDPlz0icHSHDc7Urf8Pf3lvvMKbuRKN
j73Gd7Bpy3lypqoSVElm17k3Pd9opBTE6zo1qV6VQ5vDhxpuR0dwJg1AQJL0
vNr5EFDSSiFsNeaHKLgDadniwNz24SeGA4gLWh6SiPvnXJ7mWVCUszqV+vkh
PAdea6+LlHcRG5t0IiLASrwTotAF64DBQSifEJTb3Ar483pN2nP74gQmp1Ut
ZFAZlry632/yUZdCbMzlmbcxU6KUKegP42qHv4d/0e05fqZfbZqCFRIgrvIj
p30DbtdyDO0Ru5joGJqTeQ3ktk2cgtdi4T94p/OLpjrt4S1jbbMOmr4FZL0S
DgeDTvfL2og3NYVCSvPCgZMKPeo9EpcVS7ewQOF3WwYYB3jyFOZePfsaN3MW
cJwBfQiMfUX8+BY/UVFDTC87+diKbBlMJzSDyPQJEVk/H1wRGtaukUbWR0pE
KC5F6BFRdYQVmiPi5AUqYecnXBnUUd2wHlkmZU0crGmiJa3XjJgSF7bqfL8u
dOsnDubDxx2NaAo7b7GtagVods0EbFKvecu85qvzQEi6yOlh8PaMaVJWTcOB
DJmMxP7183qZhW1YG5jteEqeBAgCRjoJQ95mrZia8TThMBCnCx2XxKh9njig
dE/jae/P1+L7wrmz9cyJbdLNHSw28OuenFPHxqj5R8P1YkHffxPQAJFXmhv1
RgQPfm7aD7eJzvQU16tJjbdeKs6QrwHLM7JILM//NdeitNUUeX/dHD8YdDKF
CuKKTofxvS9m3+focj8Z/0ur/8jBGmdHLy6QnmAn7Agl6m4/y0RxB2z1srJ9
Oda7MN1JcVzNci7iMsoc2iS/OpurrSTWRmwTzjb80K1loa4V2Co4v93JFqrk
Q+TzNHii/CudTA6Es0CWX+qBvrrobWEyT3Gw1kpsz0iOs/GVWIRtaXQsWrrY
w36FB3EcQYWC9ArGob6AUME3liPerprAQ7DF51Sn00P8gnwppBu9euRC3a7j
2oym2i6kaVUZmQkAMpF0ujKjWZU4myQA9kUrvC/AXlxxcRazRr5L7R07/wLA
+gO3Jbo6VPB1ohOPOOjmp3z+6cEgVuXU3yKXdBGHwYUtJgDth8G9vMx+qr/a
C4Nq5LNTssz6BhQLUnf7uKAEoza/dFECQfOk8e5G5Gy1jtdqaJPW1BmsxtuW
T+0WNqmjIHTOpOGYf4pL0YdSPNcD9GgShYvMHuZhmJB9imt0jy/U7spVJ3E+
3rka9aAieGeDQdj+PpHlXUtjMaAYMKzZee17XYXp1vatD5uCHkNKsKDGc3Tt
/DH6/EAbefmBOCyN86l9hmiO5nIaF8cBzokIZ92gUZvyOpT4s66FjeQVPuAA
eRKKLAg3cDZvKYweyk35ggKdll6CQsNKY1T3HlSNtggAjDS48yNNxgmJU16i
wJciYTPdtctAUryVdZcRwOOwGKl4EenOgi64/URXOtwDUpUQkScNfQUfyi3s
mO+VpBFEDLA6A4SGDeYHeACU67jzC1enB2jofWLrYQ0rEhGTy/20WVImvkGz
5hSYSvAyW3qK0ZzBpJusnySOdUEEJvxsOA6wRS1Uk3dAOt9Uj1yL/A3+RX/k
ejQt78/FrRIVTSRXwRgvVFNy+npEj0d4RsIoQswugYKbDSz9kXIZUGWWz5Ci
4+zp9eFBLgLZ4W1zqNFk2TxuBV5QxfutPhPcHDKzY3z6D7yB30l5Hdps2VLd
AiZMZAGqWgze9olRNGcrdmH1j243MC6jkXS44BYtVMTwF3pe8+PbnbhYg8ay
jpLJipnKqGDhfNcNmJ+4oIrrUWlDg2WfM8h4zSrCdXWUA/8iVvPoJxhgUKa9
wyg/xboLswsBXVc+L4bnW/WgsWd32DpMg6Lpo/7pCz+zxuVuaGwrJTizmtCX
oR2ahBvNC7aIz2whC89Y8XtrT7NudUGamuT+LDJ8e6fOSaV61SlejmbCbMr8
EMzY39YbHUCoEVlG+1/+y3v39BR2KP7unc1+pqeMCql4a2J8ztIWrZ/Ik1Sb
pc3P/gUA39Tbgp3revyNTEIK2XBozkGdDhK8i85lfV9nJaxQ8R56Q/gkcAD6
4tX163VvLohCBNWfao4cBsZsACxsmUq8KkndslSVxZxHDDRfMHTTb6vxFodq
mePd3Vf7xN82GG/n9ODYEWzUqSCzpnJHIBsfg33nAr2C6lSL4xuN/iP6wZcC
BnRi6je3tDvSb8YKfoHYjWrLqUmflL1JU9pdEQRFMJ2HQvaCmWU0vBSlp6ae
Ap0Ilw15xZaIm4HqCvbhlVxSprFH5r4u8pajgWCbA953lC5LksdfkgYynE1D
mzjlfgOkSsbdo+DPhclmnuT6VQjV2BaWztOpm6mqGQ30A2OqoKLWgnWnICuU
wJ78OLJL4noPrF9elJMK1Z983iWQFLY8J5xfbcNfJZqRD85VSqI+VPxAdtgu
0AkXcm8oi5ckY8lfDaFWw6eFE4r4CIVp3jcJ3fsbQSdG+vs1qZ7kvkngFjoj
G5RZuKe0IxDmkkB13WL2w32wRaRW8OPWcipJmdqpaEKT+gNUswLYTQnGQLzC
kpm5OTPv4IyvrkAd37c4t9bLOTLbOsVv45+MWUo76pzarGKJhFfS4JlbMK6o
RDDDM5vm7pz3Fni+02iQOnOyM4r+AdE9BZEGn6a230lFNQNGh4pl+db/+gWR
kKV5G7kH7xIQif2GUrSWLe1ScV42B3+4dwTg8FeJXWkiouMSvxs0e+e33rl+
MiJdspEY0ISK+R3BPotsINZ4p8PHlceOTu41Gksck5qFht+9W3g00pmG+u8D
A30prz5hR2UxOO/xnG++Vvwg+oJoILifPeqKXifPNZsR2ftpNrYCQaXdpYYx
E+zdrMaEdqFhmsumqnKE1kUOv9YSSle2hA2Rvcrv4GGfyMKJoXeYTap6lQcc
W1dVxzPYiCvQrfVsGCF6thT/yPXvTNc0P/mG7aa5OuTju+jXTibZoMq68dbo
34402bKWeJUf1nn0pzVT8JMMRcgKqbdIxh8i4QcHFM8/KVV/P8azpxzbBXIS
xAchbasJu0DNBwb2PLMgagpPIf7lKkS/abEooh+IZbSLscuZ0AlBv00dLZBa
tzEFM8Q6OyitECA+q9gOH2x2Sezs07CVI2ySeJ1pelWQHwdzfGw1K86FoFKh
WZ/yr17TLoRovmL0zDcLY1/4Omj4Q52hLMbQ8Tciu7rUW7lBmqaF8uUtyKfp
+6LNJIpAx2ttzEdTpyCc5S2SqC5GjOyUF23iDpQRVGIPiKFJNEYq9dy4j7WG
9yMcdAzpEFcfWschvcFxv+KwAec4+vibT5Wu88+mKuPaIRsBOCKymdZi4gBH
UpqfOySVScIYEDYsvRExLOOGDjxltWH3RqR97K8Soa5Bx4k4swEH5EKU5SAS
pUNJuB0Fs+yy2dhFgOkMdif9l3no6MZ2Sw0puLo8gucsQkwdKNW6hutr4R/6
D/TIuzimiglkpD9MbDinEGUX5IRkOqPaMYOCUUEYKvhyXFNBY+2R5ZHgLqCa
b+ecNCAgb1j2mgeYfb/P1YwuNq3aLYCyKfsrcL6srz+Xi8cnmKXSjzuMcsAu
CiTgSCtwK3qWkx2c98hd+brxQmxYH3Gb9jGZS/o45WLTeIiv+NimWm30GUwV
WYfFxZ1pzewrheiIzMZ+hFPllBN7U4KvpWALyysW5HBpfO6b3TgaYCtlCEDr
jc1HczNBIOJ82tQ8dqBGH6TXgqtDxSQ0WxjFz4I0kiDZJV56jhTDodmP4CZX
O5LEHZZiMWBdqfyF6BGEGouCaHKkLIn1Gf9PICzwmPQcSP0n+OE1eXfzNbGl
IcD096Oi2KLU3LhPEPVI3ZqDPEcadSdWBEb46IE+NKm0n85Wb+Z9EIm6vO6u
yvFLZ92nve3gXX0UaBHDZRuIKccYS0mB/gQGPiOEqk6NfLJO2nVTp82q9YS4
QwuB50OcQuOsWXXwgmo/c+h1YRf57DRDBKEHEFMDd9RBKACBBHolDK1cac2x
ZB+ZvZZ54rADyxOSXMjB1pKC3bkwdWLx2JCcg8RejHy99ZamGxzHvg3y2zK9
RXDoE9DrWEuWmZa64PgZr/U26/vKDXXORsIzEzVDeC7aEuJOuAqvquzImLl8
kt1BvPy+JyhwEqaCkOlg/TANsHC88EHxKAqNI6c7+BPUaKBCbiafPjrANB1K
MOFg8K6PpngDdPpEHeiGU9eyl3xKArJiASR6AcZMhskswMUES3TdqX3LmaOQ
I/MVld54aCX1izvp6hy68XmLNM00wyOgg1tgqXCZheaVopn+nNWbD1+JzTLQ
umweZ3+B7IG8lCBlrg16qjjDICqf5NM1D9zOUiDAuqCNtmvaMYbNA5+24ACc
o7XJLK4z7dBvtFqkUm05jSXnKWvSV/wKW5DU+Mb/aq25jQvbob+EgTKLEV9z
Iwt80PO5seUY5OGMH/3mGBVHYDq5h69w5NSdS7nt/CWWJFKXR6dkxPMdT7Sr
0QmIICnJ3nC894ZYWGLwTG5bvhMCWgic+Kusr4botTtEcBvFhpbuSp9frmSm
/zWYeMcDbR+txAyghX5vTJyqY4MISpIWD8QHreU1qsTK1LKmUcDcyNq03mQA
BdJOpe7gAoBAhY88Js96WgJruuQRaV/1fkg4/G92lrLtumwI0vZQLVxdSKuo
RTd2FE7PH2r3xQyHA0jBlqLcpQFn/uMx+wftQYWkdlJg45NqlVOGm2M3vOvD
TWewS7zYBbmIMVCA7sLI5aW3B1gx5wHXZrEIPSIqRzqWyb1IVeIIubitDxQo
fPc771j/zHAkYoLWNVxh6JAXmY2jwXf8PmQL4vhrzqd8FDpcLORbOGGEELkP
C09S/sDrCZuOe+TRi7VMxSI33rgYI2WsDBz2s3s41y/c0AzLJsqGpOz8Kguw
1wG4FrMi54xn56EvIbsfpEGa80VUwF00KjzcMdjUrl+wDkMu8OET3ryBbPLs
QdI4bSrNc7P3iGps6xftQByrEUtu3xBis/TG0v5eeE7n9EmHP8HWR05b3hUB
oz1WxiE00+aCtjNOme9F3ViAVuUYAUetlBGlMJKRklTF6OMulZ/FU92FDnPc
qCoYHIo5o9awMLDNNZ1gIH6R3R44yrc536RUNXmXAcdzxKBJSneKsnYny8oT
eyKSPMlSysrN7IALSKVrsI3AkFlm7xgMN+vIv7ikcgzqNaNrZHFQ9Ucs9p7k
bkv3a4neIj/pELDTVr5GWKKcaNX8btDtcc+dhmbiY3Sr/vG7QXz7ImSPP95R
NeDAR8OIqGQga2OqXeLgP5RJXKbEgmzOtQmJb7hfGqxC/GNuuqYuU11dh3EP
SFPGO0yobvaHMuOVIIFlE8jU+tw6goqzBiUYpd6QdoOnaRdd26aw19E890I4
JAFX+KPIeMvaACNO/F31lZdqE+mTOkCPFIiflzE/uaQu4d+J+4lj7pdrNo3L
QqtWQWiECG52ZjT0KSANzaCLZdm6tvpMfXJUnhOCcoRJ+LTz9nseKkHSbbgW
fjokj5p5iR8SDGqMEAiArn85D5grg5XrxDOfzenJL1G7PnGWZuxj12GKRaAV
G3Aru1aubTYqhTyDfFIAvAnWdSJOU5irBHtglLe35sw0pUe6syAscJVJMrX8
gysUuzP8be1+Zu2OsVjnSFiQTveWBqQggGKl4/aD/TNJWrfaDPzQzebF+giw
z2CafHLnmgjsUGH7H0DIFR00inmv5C7InFpglM69I1cg8qmSrsVzX/Bv7w+9
hOrhUAenNg9MZOCQOHFQDvM010NM9iVU9+a5kQxExLJm0C9jeMPMWe6rQSfO
/vTRfg2DqZ2Z9Qwtrmwzk+4GumlS0XhoRR7MIJBfRGssCwl/kRboR38Rnn4J
a4fZg3p2jEab6OQ31vxCet1M/R1n1tz+1KM87NsSvovHqbkKJTC0Vla/FVhc
cxKO9b3R8Z9yKo+GRKzRiAauDLVuFX0dgTcbIBCByFg9Jxwl/wG3b5mVA3UB
mwyvjN9GJ/DpwSLMaV7GcOopHJxiroY+XiNExhTJp1EuvUpCWvlQNn+oUm+C
bh2ovSGAxoPfOV2DSOOmwbLyfEpKJvAowjs6FP84xGdNtEsqfBNfdozJJQJH
2Qgkntlh0dphebmpnYcTj+BR68cPNWbi40XgnkJlzc3eixvVO5jRONbYEaYv
egx4fqSoUbV4RHmAElXER1C1RrRs2k+7qqaYTSkvZlZicPsf4Ss+XGUmVL3e
XKQUvnDahj8vuoR4qpC3xckQec//YgPKPgoYWaP0swllBWReElD5RaBOqnQa
C2MXeDdXmvF+mntvZQr17ITUffFAfBAEAiIIwS14CkHd1e6DYquk08Ch1pWp
NmukpIQVXJdIRJUxqZFeAvQPuROZyHppbcLnYhDzNyd0r//wCFTRU3x/u++t
IUfi8GCVdAKAzRyMvFjZ2DTpEFxz21Pk+udjXcdeQRAN+N3K4FobEMZrb91P
sl41fmvkOoIudIcjjU8dYhepOzuQ8CB1WU07Y2Fw9K4Im8fpsh5IeYtQ5rMM
A47dqHwD1rfQeXENvl+sxFNZA+OVxrCccE4nN+jHPqI3rKbiUrYenFWExr8p
H0DYh34XsbjMHV34NokNW+GCGVXPPRQ7NmjhajpTSZbxOmpuz5B2368Ew4Q3
cs20XQO93X5H97JlCS8+Co5urfvdo47q/8dGAiKjQjpbxcvCV7UiKLbvFhlC
TLyShfjsyKac46MgSl1Mp4C444yCi4ez/hdNlpowR7viL+rUahLOa8p35KP6
Z7lBCEgd4Vqx9S6uUwyKDXM9n53kfFG+/w3CWYKknuvZfMrqhfO17TckJ//T
CotzFP6wqjTOheYLw3GzQxJ59K98oXnxFw9eX2s1c4j3QCEmkUfYvlz5zMOn
4lifDkQ8iYl3Usd0GVGZaELkM4fDfK8upx0KLCpphMUYfqRQaPrAnmXboTa4
7foHQq3msDvcJjpKyGjjrNc8i50+rYlRTz/TmMe7GP7NC4a4G6Gb3ge8K0fJ
0sCOfK1Dtag6JYUucFXk+AaHdPHrTYVkpcgcgS1t7B3jQkBzrOzHZ625sc4p
7IOehl5qOfJrUTo6Ol9oKA81oKQpp+cUgiCDp3bAf8bGFZBbJydl9jxxzSQA
CNo/jQbZkHZfTnEAPGCIJs/Xrdmk5kKyV/emrrwhWMZdexVJIXmJhIoTsQKk
Vbf1yRcLc0k2zA+OAxXBC20QwhgWs8ymrKpyGL9lT3uO3pxlrjwJUk84NWbe
LvR0yZxJB50Su1FuOdrR79i2DTeGL0khb12ZbU7cekiiVrJMFnK2ZiSyGbky
GMiertnj5dTokGe0+9YW8qdWB5AzQa6dvAjUR7Are85tapBTMj2pe9oKiD4H
5eVY6J7DKQWT/ZaGa4lReSA1wEkXwZpkFIwYQhPBkshjQdZpo3+IoCwisuA4
oNypY4XZtu0Ydj1E2rzo06FttZhEvMLc3V9nt5TnHs4xexC+tgxphK4c0zst
L3nAUgKqHu973Y24yDtGVbtJc7XQZdAEjs+HZITgcul6K03MFkloLrZztOTX
XRBP5LdSBFNQYx6AEykeFvyVqhtvh0v6Tcq/U6uEU2NgcbDL3HBOgQojLpEJ
zf5ps8VlgVCQWIyMb+/Sa65cmGnn78OBcC8fYUJiHT88SxA1jyiyNXx0Vzv3
NiIGIaevQ3A+aHuQffxlhXa8LbsZPxe+MA3LtQKTBf8Gt3Xe0NZVn8+TEHLR
8iWkBlb7/bjRCE4sFk9JXWNIxlTCSptlf8Cf0QK3DsfktRToIoI2cxFex8+y
lhObNg98FjmDKJXn3G0W8n6ZGyUA7Qw+06Rek4iqjcAeeU9UBkq7yE/RT5eX
Is4rX40JMCHtM0/tfSu3GZPdcG6NObPd7RLTT3bxQi5Dfj3MtdtnFk/Tk8RZ
blTO6aAoDsPx4/Seb16WMIH7T3RLekCXGi9mANnAyVdsonxIAmO22FurCjWU
KsvMDcWJjgNGbxcDSz3I/CT1LPLX+993sigJ4Br3FLzfjU+yi5KgXIKfsT9/
rrgmfMmhGP0KMGxfh0l995wvQZTZGBYFtOhd+cbPMVIJqadlBlqoUTAO0dnp
Ljh7CqXa1xRE+jeoUo1mcYl1VgE97KVFGRgrITv52M8Hz0iNsSX7bC2BEQJR
efjgIKA/imVh9p8xiG+CSic+iKT/9hahGxZbbHv8joeRfzlGup1Gy+lCS8GS
JCKZzvJ6E4pjWhQNwQw4JHTEmsOkhAUQfFYwrCrhYP/eeZknHxG47a2RVzzM
pSkp8alA9zXoc0xfvBjd0EC7RVh1Lzut1e5FXQlT/0P89o6/l3CkR8xt8U4H
nn4hYTxM+yWUAuxEdQ5rBihKC/B+a4bQLSX7/GsNrufKUo/bsW9s+oxN5kc5
rJ58q7z8Y4irxW7ZYtDXbp0ZCQ+H6JGLUFB1e2YEsbC73Byl6bdSiYypljpM
BBG5bbqtCdO8iHSp0QZBr4UPlpC1b+/rWD+aHCqBG5C4sJ3IjvYsfwswno/R
y2Ev8sLcZVgAynKs8kejSNYm/ewrbbbmYCP4CKJSVjELq99nhgIXzirh2+qB
poUGKBS31pJeFypwy4XA4mJt9sOvZucN3VIKZfELTY7JIkdypjKOn6Jzwc/P
bwQJ7l6NtvcpfTkft468XV5b+ZlDVbi3Yzp3/G8I8blPnx8AmjZF7E3TqcCG
xXmL68jJUcwGLaGV6wnZ7UpgOGQE/8pkZJnk0tW0b7xk2fR3IcPknfpKQ6IX
RQfWNMn0BJj0Ywjo6SH1Uw8CY2cnE+4XPDa682/BxFbz/F/oOZ5AHtbvMWul
nCEzM5MFD1gW6i79fzYvYTQ5xZO6Ia1j7O7ZTD+PMLpefmKw0fJi6VLGyUJn
iBepQtPpxhqG199HTEwo/dcZw+x103Gf1AS5opMHvkE0ii5b8E8T1QzMO/86
99ZmcqJFlNyYMAAJvxrtzYd2JvmPAJ94kgq3UABauHbU5z/sTyZJtLyWjMJj
mnx1YdHNZBreHsz1JGtIF+0OrArZlARu2ReQF3fuTijgB2qyVCZQrMttzohk
NMZ8grOjww1AkOZk+5HPs2vJtXfOoKouLhkxO39W6iEN+OAAjAdP2oftqqU7
1YPIau2Sb+DmjJUSn2MXP2Pu5/AbMW462s0LJRF0/qSNGrTSFtqRdDGDorTh
//3Y37zVkTh1is8m3SgcJN3uJVYU/UOJZ7KX1BLC3OWzgM/To4PTHGhhhDxz
HbnugVycdYSJzhcbbRVWvJ+fz7uuHsxFy09dggd9Xu7k3NPM+8CeV/6kCZR7
wz6LcUsg0tCczgk6pcbWjF4cTJONcbHi5cC399kWqyT/ne7e41KssvkOgI7u
AgxbABhIGsQNLBF1iAnU0WfabbqJCYAd2sO/u3s4U0b+kYDrFhLSLH1Z4p0G
t/lbpwOFl9D2NZa65ZONbk+5AinIAPKBGffDe/NrargIZEUkp4noxSVH2EJT
49JE03qOQKdnUj1Un10rwOC2Ye4UDOoXCCeRRm26LUMeD4ErkcIf21bH3Vsl
IVxWZl3HfFAxtghABISJptATMgKgCmG4aXgXOHXy3EQ6RoTiLMz8MWoBflXQ
ZuTnJV2VWpY4OfDDrtqdi1TOxv4ubp8RONiRSwNlogMBR04D73fGWpf9xgXZ
NUsvWbfqa0eyplox+j2tAjLIDqrU7qtFWH/DqEDJc+hBbccrQQlaf+PWmkWa
JTgA02CM9N1mOX4v15nylRiUu8i4vUYgq52fjiEuyemGQ6BynqtIVSve9uVO
WoMYPbOtD9Exef1FdWVh5ASAGxJg6ZyrOp/3bLoEafUUuVDdXr1v+YoCVSmj
7+EVdf9p4RgA69zOGDEOKZjGbYxw1qWSf2xlrZkP1743Km7xt5W40pM15sjL
hnkWUrbylnP8fcs2vpFcbYuet5ffw1upkM7IDs/Nbz8ONnhpj3SKxw0Guv9I
gaYAtlJwRZWutJiqbBBiTVL7rxUYBog8mLt0gWxs9BiLmArilkH0OP8ro92F
41yWLokaPQZwmkIjCc91x0v1vwZyQqDjEpmqjW4JEhJhWtnW/gSB3FFsVYOZ
lw0ho3EBcciGRnoUQl4X+raAOsVfbvwkpqQfngGKJRGDuMCo0Gdjpnn8yFub
mEH2S98g+wNhSFjSUlHLqIxsTYXY8hL++Kb6UfD1Mi/8+58d8flpp84rR/Tu
Z1Q+fzGmP4o6IJHJ/lVGxySfJ+1IqfHoxTp4z6k5QWB+y/9sLf474byNwbJ7
8PV0CKdC4qkamtelY7Gp6KF5+4BhuIzdB7cNyQea5wElU4Q5RvWzlREeNlVz
ZjqbupZigi8IoaitTjVCFEJHDupc2MEm+j+aSiWv868XHL/x2rBHC0n1a4BV
FXnDgIblyDhC3dBB8NvgDcN46BFc7zdlMSPR1WcXI1646bKU/2QKOAZJalix
XuhuZ4FAPS77q0O5tfolmrTOVihrAadcZYzh80bFdidaHser3IdhXFpH/Z1/
aDAC56reaJ923AkBUmAuWdD39EW87j3Lbq9BZ0Jq5QmePl4yjCX49ux1qahL
HPPCIOd5sTo5WFKB9q+qrUO89Eq6KrjmuDJhtnYiQtGHVFr+X1edvTPa+ZKl
o18l9WREkxd/LAe3ARyznLPKJl9w0380w11wLAIZYhCRMHRa6qsn5Bh8lLH2
3XmpxUE7Dwbdo6yFHV8GBjRhP/3UQrsvON2+OoJYu1jU5n3T2fHyjE7H4eRm
7Ch9F4SqML3vLFNPisHH2NCArxd0mKXnj5Eyxi0HHqlZ+a3NI5Myti4zduvs
RpXvhy+qvyjMmAasOKn2NPeWHO7XSCn9qixf8ENxQ0Oxg9qwrL7i93LwYvva
ur6Aysl4flRb97h4X/DrEcIvca4Acu6khoNmHy4LA5oP35KGX9Kb0z1Y+zBi
sM40AtLP9B+7qUSDK1WXg/3/1/IuMlcRLB2gcCN6eZOu6Sk1PqVXHF9zesIB
sxmd1Idl+dRqYFLzO85uDif0Q5mSWBxpJ8Wlx/ccgGNdAg3YLX9IiNSifpde
H2IAgYQ3VphKRlMoDkuBf583xKj/314NSErNnpuVR0aOzvaOXW2nl+3p8EKX
Nm9+Q9d4RihcRnYejgFabRs1icsh/DhFOHYigeVaVa+Ib2sIud1WQQa6J/yl
AU1+3XtAC7S6RfQaHQFZ3sdHwaFzmIU/nqFj8mHePC7AO1oaEKKu0M6Y+eme
4na9Wuq1+ltTK+ms55GwztNAPHSBQaZ7Vhpg+94Omrp2xxUvoeYPIBZuAetN
XDJIOfzSSSyoavWZTd40hvio1b0Vpu08OmgqelkvtbpI3CbHZ4q1h5J+IA5T
OSPMxghmL4YxVpqAOIm7gP4ZzeS3I2zrX9E9HPOok5B/BQI2vH/A1Mmbh8Xf
wFMeEd3yygxmS3YWEryLJejELhwULWpi+wA97ojIPHzhbwN28Pvn6TtNRK4H
DaglAcvdsAUcl9VxPSCZf2ezR8XgR1425JKnA3spZ9knzKyClyYt/lQ+35EF
KPcfNOIyTofYeQjCwyDjyrzCQI02beFe+ByadXMzRS5YKCHlNgabf0LAnZmw
GseUsGZ8Mf8IvllWnZmYm6L8uro1v5IzHD6iOwU7IwRtBlX0AFigN0YRXJgL
BQ/ECOj+I8CniAVFizr88I426eaMuShw44N4kJVHV6IVBzVDt1d8EvMEXrL+
Ky1ASmlL5+QVmrhW+Sk5cMhXLqkvsohOV7JYOuX9lz6pBV8tg1m9+OahzRGp
msOO2uB67/Jk7/07Dyc4VjgS+XlhNVESRHImOmse7szbJ06TExmPDoOT1vtT
y9on4T2/7VB1W45OFO9EdXLsi/DyKuc+FotNQQtn9vYxbbdxzLV/lIDgg2sq
NQhOlDM+zwSV+3lIwmEOyZRwNTeOo9nVxpWSS81bMN9kdjg1FSru/b+yX8X5
m2GCkJiVQN9W/eOOte+ZxWhgBK5uoGLtAE470CIbCl91UlH3twfjkb7RXz4C
BfS+jPkrexEGQRhG7iAnEUl8iFr7caxRGZkS5y5ru2V2w/Zdt4+CUwg1IMPf
P1CaG91vYdGynvVNRl11mAvdtK5m6DlGphrq3eJ4QmcYIFyCO8+3ge/LABYk
bRLaKw8P57jvLkd85ivQEWhUN9s9yW9scr9TanbfTl7GMdy58VtN9lAXj+tp
DCpEofBUwgFUGS2oL8x9CtOsBKSCuiYI0Q2N8L/GZy7SjndHA47xUVScs1eW
d0opmGxWO3sY6R4eyNz+XrGr07yelIngNInejDvczbOLyFQ/FcgvjFMUoLjf
v3NgJ7ZxEXWfyJtXCoDXhlLev1M+YeRQr5rXTBDf2vJeax/BLRpWZIg2xAGO
Rt/nhlCRrmSBeJHTDVmLLiICIbTRLVL8r44rY/+H36tnB3a7FtYLIxfiFz82
2yU09k2TZ+5tISDJ9e19i5eVwhs26rio9csxi9O+aaTWlM8VuuiO5XmEfe9z
uEvuVM+ukk74hwXStMl1d2ZDQR7QK5S1CYZoCcIl6HQLAIdBfqi8vIpxbVHL
2eK2T9VwN3KQHSLIP1IKC/SzehbFd1G5/T044YUhLqFtjkTAP+Hh+oUnKdvM
XE75uzp1M7o3aOPrbWiDG7FULqOtZ66+gvroPWgH88at/83LkJogZuoiEfPz
2QWvaVIBnW1ZeQItNa6xMzyWana1bvz+JL9rVOfb16vlaMH4wKYynM5xqVO2
oCum2mbOtKGC7YvwiHNnAPibqaHw3Hgd7IjpEpreZ4DGOYaxsrSP2p9S/lOS
n/fPK2yVXggODthOfFjlIbg4puHU4NIIPXYWPhNpi1d+pMUCTZgBVMsNe8hp
TH5rhL5YJFfXlnC63gw0CbJja45TsYicZsoHZ5SRXcGGNq8NgcxRlh3CaaB8
Ee2WrUA7VeiHRRvtSYOgkgLkz+nNo+6/m7c71Xdo7y/dKmePb+a2Wnilc6mJ
UjB44QY33o/Y7hbQwm+iMivoUSEZGJL2XnqdblB4Tmp8i9IH0yA0ovOfamA6
ODe+uXiI0GUeeRfC8IDYiLuJY68JPZxW+C1n1i72RpsJUwYLCBunW2ucyHuV
owak6WcIfaPhOe5c8Q24TMD6TH+/OCpuI0bUpgKTZonu1ITL68CFnk3XCe7n
0PZ3V5BkE0ngFHRaWg58wHEaOkO6peA7PQqhAyJGHt2z+0umMs8Morq2AB93
rKWza5tB0ClLqNja1Q2ZVYDanDR4P9BlCW1LzIe1ka220Tc+CKbeoBe0ESre
3cR2aeUmkbWO/mK2G5TeAZlqMXc8ZpPEHWpGp16kL9+Jao1xqAQS4Tq+xd2F
+E5fap4mvGZzjCeMD+dvxxgqid5iE+rvKrtBsidgzD1emlQf47LPDSZHLVTR
OwQCILr97FYNfb8kc5OmYnsf7pCVsQ8+nUIZm6FjaaLRdiHi8g3MYXDILQJ1
xJ8jQAjByetAlb52nxWsX8yi9ow3h+7vJ7+vH2+QRCERAH0vs8g41neix0j/
dGX8IIBzspRKH+70lNJk5U82QVnjuw8TX0A4ISFjgqURPPvpa8/FRanNNmsY
YCZgWYZUlvkI91BpFB4VSYnayNRTyfASgpj+h73st/0DO2tpCfcoG7wAzM+p
Buy2b7xWlAjhXE9Ejd5ly4NalODUmbn9TgMDVvD49ZDWD9Q9ni2RctkD2ppz
M6welklwsUq5eo/2/LTWWVWG0sd/ooUonAUrvWjHKu86DpZZyu8PuH6ruDkO
Bfq5c+D0KgVmGeFgy9H5sZIYizHvd+ohMqf4AYub9CeOeMdLoTFQWlKxYI0C
+SYYMU9TAXhvh6KK4GQjx4Z4fYyvnMvGCrhQT5O4C0zMCGqXeA3hYcR1gNeJ
aPo3HXUUb7Dn9M3rjl/DfWeGFnXIlWoRnsEDyBB5BpbQTSgAb7Z9EHe5p+Ew
lrRAmmSNn2s1CRy4s6PEjHSRpzutPcRbcF7RBC7YXR6jf/xfgSxMnH72saHp
JvpVtPHkVB1JJbBqKBAucZkHuwQYs6dKn7uKSZV/JDXsR4/zvXgFhrSwpRT7
0bZe3Tux42vqIzaKt4kCNzp5MApyYtvyDsZDnzv99s3q7vwaiGfAQjNTn1OJ
5EXdFz65q7chVKDlmuQMV5sUaadZplEC348M5f2nm7a7aI9oyGOLZbv+rhrr
ALHDP4KctZrrKFx1BEi60E1K08VLP8mukQ8oZd5tvEQOCGG/3wTCl+zqGXEV
E8VRaXNf6+Wl8xu7uQBHajF+CJ6wf6KUyJ6P7byAhl2SCZTMkRI9MuZ+vOzu
Pb82+TIwzwVkHYtC6oGOTnBqtg4Qin2KaYO/HUypYJRcFEz7gDdEAtui2GX/
3PaXsjbh04eNWdWs8/v8CN+mR8TI72Htz7SGA4A94Au8U/kJbsPFSFHAgJ2i
2/Mmnz6PoFkUMGTQxLByb+zuMb6RhKmRJ6c6vM4IC4hieQiIanhk/8NOb8P7
0CZhsq5TxFHsmBQ699TXr2psNevIcEl+SwBrSV6pc0tHFvDucV0v/5Ek2oJc
IkR95QCSinRuF6y+Mxiv5FdVk0XzTx51xazu2KY6vYc13B6nv/vgkfHfLUEK
fKvpWf84wUh/qORHOueI3G/xeGeV5dobDTZGoA4f1kgVDzx9l9a7PcfC5e4Q
zICvrD7tteqXL/gfWmvoijChKj+uAt23wOoGUK0ZkY+EGAqJtnmDnPBz5XCi
Nhu2SSmS/43Wp4njtTrlR6r4/hMGYmRqp0CL2hUKRqtPnd0Q9AMKjSQyTQS2
C/EJSwMfHrO6A1iGlyNzW3dYRf8Gd46VHpim78Ys8vS0ZXgeglPPh0O0Ja6V
NPJr+7e8kewXqT1FyQX19KSwtVJuqHid5cRZfTbnaClnvY2HKqXktSUNH3sz
MHwGpADqDgJvs4RU5TSjxmSBxyaVIeCZ29O3Z0oQ3y3r7k+I1aLAx7uQJKHB
flksKNNqO72yWQdzWPKK3I4XtTnqWy7xs4Dva526cwvX/zjerrQ9R3go3LLq
TmiWjEKrlhrAC8XNQ/CyudC7QzjIs6dEyc9FM6Ym5p68qyhd1tqAcAbLUfwg
wYGtf4s1Bf8esnYZWyDif7hUAVsjqxvZkHjyIJJ7/XWXxl05QPLK96ozPr3Q
XcQS1lcRxK8NVuTA2lj6PVEoq2Icwumh8PKjyNj9U3467W50idRr99J3T7ei
6PgkLJAD4cm0EaiDXxULpQOxMVpoVK0Uv8wMvfa6IiTwIvWtsqws5OGZBlGI
J0XDRIqksZ1dhE4uqskA2lfmNTAOyfp72k6GNdQEtY/nGLdDULDb89uU2QE8
ZvKOaDctn9OTVIpL29j0mok9GMWAClxD3Mdb8WTNMRIqG8obtD6VowH2dyEb
PEWctWQxZGXUOgySFaZ5eVdM7mK5/jsBExI9N4T+bO0AMfka6Lg0N4Mkz2WR
YoLI2vpX9ZAYsKOHwqIXWb/fUvsawMMqI2vDx2OoiuI4HwzGlPN7FRhMUC2Y
i8bnbVJo2pWQjyzxr9amnEhfD94tZO/z1BvqEq4fDXlLqQi3zvqRM9YLfUll
djpRfvb84EKFzGLm1T8kMx7FWsoweg0kFXW3wtTPqtoAMaDMMUV/MujmxUsW
6VGjz8gK3gVVo2m6yVnHTvcnJDAqzErauIsJQCJG3o4dDFQ6tktBQ7Jos/Oq
c13smPCQ0moK0XmOxw+jGcXvRltApCjglGrXO0U6YxVL6Ut6bwB2brWCEqlq
l0IFfo/QAh219QEPBlAX2Qzx4+NPTIgrAQAgTAJ53gE6Jsz6PT8Vu7oLYrPM
uRZ+GOF0b28eka+yFakRmbzjct24mHiRk40h6K4hIYkac9XUDrRlw4JlsGHK
ramztyHlbhRE+LJq+M7kYChL9sClHYfd+DfSTk7cM3CiDl/gMi4Ky8IEiVKs
MqvoIEkhT2M7ov8zM6qwgX9re/9ze+En4b5f1rONof3TO8mSXFhR9kDZuWuN
Q/p+hCs4qiLaSlc8NAkJ/rdXy3t/vZoY9Zui+uek4XaJdaygQJh6R5p56E35
vBt8duZC+N5ChA+imkA0KwhoEARnNkbJXipN08EhLjDUS5qYI3yclIsc7CZG
7X1F+o9bJjUzm1dGTtNGouz888O9Q0mRRLf3Ru6NfOTeXk39nyydVlXRyaCK
1ot/atUioVGIh5DfnJ1eh2vS5UAn8tP0amWciuvVM7JrbsuOw5+VyalbS/T1
SBCKQDBRIsgzcOG5gBTLK8YwO4mQeCQk8rKppcwQbHy7AEtD/vywt/IFzJYs
d/BvhhxYZ8+vG99zpUzx1MVhm1qaRvShs+EUuXYC00MdzjhgYw5Av7b5vyYN
LMUSMJ19LjSh6TRpxzkraQiJi8bYjrQcF8sGJHN/MSR9sbhqKMCmaCA9Y0jR
96YaugNDo3OnH7gfBR7Be9REBLtPi1b7MgLFR+ABw3QlI0RxZuJ46pvRpyLG
JPApc9lwT/uFjkD+nHN538o2iP7b/czb+aE34ZrjbFy8EOH7fWcD4trJNJAx
6H2IZCayiOZ/aSo/ND5aCswu3VvaJnleauoWv8lGwR2B9YBdI9edH1AQlQGZ
r06uvQJ99WJ6JI03IQG4+QnOodQDWQympL+b1NQQDU/IlNcLXjnAygHes5LS
rxQDzxiT40NQ4mLyS+T+m5MMZF58NrCBIxdLsREWPRC+hCf/ou/mjQ8MrmHv
6E/1OdO5GdkFDXOZ/2ZgugwQxQIZmer32C6iJjv8J2yCYoruQsrBktSW7fVv
zanFWmS9YnEaEKAeac4Xo8mfvd25pOnZD8pX0dAPlcV3xfcqh86pmqIumMut
qyHeRukxRB39mLgc8nuu6CvmAVxdNJPYHwlnkHe+Mzg2QR07pQ1HTpqureXH
y1jNXLde1fSHmoA+foWhxhlpYiNAHBAdy+bTA8BRQ2lfJY1/TkABkg2EUaEM
h2cR1/DApzimHpwsaUlG3dXr0OjmZ6jsrejItme9pAGYKVxxBZeH/NNROubQ
4oRfLPoCFZhTIXj/Ulb6P8VUtH/XRIXXPqfherSO3VZSb0c8xEQqfpeKq3nw
XzyOakrADzoEfOzXrXRJhAU6cTuxlGBwkwkoyooIN9Qbyx9arsbCxvZHd6CQ
fyGlptvLrWDdT9iJf3hYPeB7IbmoH1farCEpFqNle4XeH7CIe8i2FSRgicyo
2/9m8bZqkfvAFmA8l/gmLbJBQaLUQX/u5gBxcIj6ntizXdAt3DmawBXFLH2r
EJUG2aNEOS5aP3gG+zVvVZ5Oa/gEaVVdWCX2TwNI+86Dafws9i3KzCEsxZl7
b2cAM2b43GuVG/nZTVZAfNzy7QNiPvLWWspa37ZF0XC/yL4iTN830QjcqpA+
32eP1tJj8WdBFePGvbmpDoVki4sDlyvUM0XBFdueW6ELDxOvCi7akcxDTs4E
F2F7cYBsxtYxdEplzYD3LxAaZe0d8HiMdZsBnB4altMtPIsFQx1IX+mKanWh
R4ZZEfJvtWuRlMJKd6m238FKYq3KGS+gqRcDNMPOndPes2YOIq+yq5EtomzY
uaiPxehAZAvxITsuobxI5K30/IaBj234YMaC/HQZGZfiJdKIEnjkDSxZDHh+
TSPJ1P2LUCyCg08jOClwSmq/1akd6dgPFtT+5lF4qKyimxE8kPzld6CpdD0m
99NGeod6YI8D0hI/5yXf8gnqGOalgHhMzliYn9B/1nlgqGA4i9u/J5X/8rzv
Wra43RSgIVgyLM8OuCOOPQpis/gJZ03EZXdvxgTN4E9VtN0hI0xjzoczj6ps
zeoCwZRY//W982vqxAtQ4c9PuUkvSVWEMqvYTj88J3pNqICm9BUzLRWxykAp
fnHXR6mvy7lr4QEJwaqEMhSfP1NB2J0vUl+tES1+JATj5ObHTh3M9prdq4rH
EIaifsAiCeYvUNHGEZVl8M8htLYB6vMge3ZVL4cxlYID4ISGPJttGS/fIdho
eAXlyFvHI4opFHPCzgSn6MGNRRg4mZebu174jgTM7W7oDrK0QTBY91b8co8N
M28Lb1Dk4G8xa7cUA7/9cmgJ2MmPoC+3oK3+SAA6XQ6oI6PD0sXgBbz57W6Z
ZRg+oQmzE8pjKy+MIyBdZgYOS72Z8/z2YGO54ipFnDrOEU9suSkYPo94Z2Jx
hOyVcmGgnho5uKLJBlFFymiznRMqZI/LZGgCNLr21CbewbXlYDiPM+QQYgdH
rCNAqapG0C5Soxzw9VjwQ9jvz8C+QIr+xGJJ+gZCcAwMjS5qCM+SPdkVvULT
qhGh9JcalxhVeAL85FOeEZMG1EHSsOvKVUp5AORL8uF7OD7diqBd2fn2NTNf
0ZSW92NDTDSbz3nTDYgusD4JOhvWciDrfdV2k2oF6Aiw3yfAwnR7AvU0R1Zb
qDYTdoxYGuX2v7rW8Daw7AWthRzaxvJP2/xgt5hYmaen8Glbt0t5E8kQ2X79
95HC61V8vdn8uYam+EpOyialyLhoHf+J5JTgVnG0W6Fa7gfBO1bRGOUZHNGq
j7v2qovfdw1e1U+vOY9Kx829gkRWVrNYTZ0Yk0ns/Y8USsNs+ZV5KOUq/NKo
UoijRtQmOA/sNy59Fv0EWGdAHllDABnnsLG1KjPVjFiGJvIxcgMmPQeMeUeO
n7Ymj/i+L3CthlezefDGyMkW2AApWw8PtSzagr+CDUXBhwlFgHe4ES75GmhY
Gw+9ANsvvSepXWuhZHa5kfWLkvzU5kRcNpTG54ntdclCHrhBhqdF0GuNQ+vd
semxlAuQE4D4/+cfjDX6ybd2LutrfI7bMnMsmplw3+bAYw/vEPDiVnwrOWP6
/JNjpH6Xr6PAXk6hY4rzCu0q+OTxrQVcJ0OD+v5oFRu5xTzk0pTrBF9/g4tO
dN2RbujBEHimhVHJBD9rIzP0n7ZWNMhmHVhzR8ZAJQbFOoITH2yK4goqnvV1
uzIiEk4eb3LFRjsCdmF6NV7waGHVkw0prh2Yt6D3TfH0Jb9/xQmyoD8cv/CQ
1LkKezR3qY4eJ8ooJuFh18gszsECBf/obHPC0xhTFP6bwhognpRT60YArx7U
1mvBSa4z/PGKPiig9KG0JaH6cG4ZYxLWwBr2ZAVH9ocmOqa5pqIT7QtykTqd
S40QGvmpSivIu+NQBMU5yaI5NkLW7ZGa0OVRsOJmglZ1N2CpXyqj1vndBjxv
2tFQDqOy3FD2ugNjuP2YYYR06ToV5qLEG8+e1uOnoh5i/pyXnuzQd/smesWz
vSqOOfbA/v/fhpdSG6/ewPfgg2aHxBC00Vu6M5Smf9OYZz94Rhg+23vxPUVR
m0T3aWzB3UMQi1VIeNHvrIS+UW6J0kB/svmhxq38YJxxc8htSxFqm6waMpEq
b5+mzQ9EAtvvnD5RVHB92S8pimcC5RFECLi7Oi7aZL2uE4i3t0mOlYQeldwy
QEXnARqKVrcqrdBlC6d6wkT5HgRcwUZw+rQTWFmCaH7pRDSgeeboRWGyB3v4
OKs8Mh2TIPoACmcnpGg4eyQeZJJdy6/mcaHkGxEEGgFbrhYSmwaJDv4TZuTF
HmKr8HKqA11HotVuc6jm6HYSaQ2XpGGf/4n5splj4Awf7WNKGTbLTUnEyHMI
niqXBIo97nPQgH9kqE/zJpfvX3LzQ8DIJgRm6m02D7KfXS9X+8/AMAcnLv9B
uk8OKxKX7Dp1pg/VU1O/ZaLPVrOSmfpLWKddxR2h3GU5wblCc3bxzABFMUET
49n5o7op48moLGTmaKZ+WQkG3+B0EtqZxyDRY7DWL8R2S1JE5hEV7SW6ajqJ
1hqwiedWnGJKKofqGBVQWnuNqcibVHvleE3/NMbRu5HBSgSGx5dYgYMfRhyW
7jSfHZsbrZQQPk55un3bBMBTiBD6X1Im1J3TcKPnryZl22EDFAO+K7PCnNlw
e5yy7lIT8mjOPL58mZDxA7G05D2Fcji4Rlejli1vWw3nZnPD8jAPEwv4rcZh
+LJpNXzjxLR6/XpDMmp/XkvlGuHx0XzxHhHa8szB7MHCSI4kkxPyGOZ5E7CG
yNJtDq/QVeOf+rOaNXUBtqTh6dcD8J2rQw7bzr3rY+7uzvxTdMhJ6EXTSb5I
mQorAv/v+zeyEfb7z1GSiHVe8xEmgV5yaV4p8vEl5x8HKGmXAsD1Wdd1mzZp
xUj8RbDM7YfRtmfxn2xByhx5Tz9577I8hWEEE1VEFiNb+eaUa5KDKe8Qu5/S
TkXD38DE9G2TwJtGpO19sxIHeUrDRBBxfhAectCxahQz3F2MNp4syi6+xTwt
hO6uSnhJMxFaWeA9LM6M6d/TruMeqoKxVNFTR2wI2aLw44UVLqu8/OnuwNlb
NC2i5tDGRGwmuSZToPYO0CNNDtCYklRq5aqfzqwlysk1y7bxSTsF+n/9b3QR
p+uQEMK0jKT1uieE2r8J4w37bvuCmYUw1BTTw6gJneYqpGgXUezu/8XZN/CB
BzUoev9pAZcGavabFNE3vpYHIoYtKM497cRvU5sjoR2AVmTrnJTZmn1EFwF/
/cJx3jEvIDz97zVpnsXNlKdb7c/cJNaRz5+RJZHQ9LKel/pPLIIfqllv2zob
+odET7YZPJ6rhuhFyXMkEIgTilXi0r09cw2i2OTSGnWFs2ekLhLw6olgy3dj
gxpQvwykI4zmXI17dKWr9pPB/DLH/DePIegscAiAHFTDeKV3Vx9O0oQMlCOp
6L6l0VXfiuZQeIJMBDE0UM/5C5f2nSrX1QEnQUC0kotbiVTR+fENLBs66a8h
7qQhFtHr/h5ujl9l1XBoc//YgZCkJyShaHTIySpvZp6aAqrKAOZ4R8sjQ1nv
eFdR8mOlpCDzrc57GtIBOyZQCYmuiSHVVveqMD0KHmG18m+0YMm2WmxBAvVa
zZ8vnkGY+rZpEgKavApZeAiYtpG1UCy1RSANYClwtJLuh+KtfbwkglElHoNq
27hyHRScrn5Avr79uMsj1zEiDqKxeUZTfj7yvQwM7pKtgiyWNwC+ceMd2Iwj
xuRoP+NrEWsV4pBkmxvYoswhI0jLm6dSGc/Ql+gRZNCCNIaev0k5uOKnDbE7
OiAQZTgef7mVofmFXepsSgvs8wP/2x223mKMi7sWEG5dJYcRKc0zUmbtI9w4
g/bPjCezk4CDiW0p81YM+evTCM/kTQ2IiIRt0GvDSq3FNeAoUYYiwdGhj+Ku
S9G7MyNWiZOoR3k8nGYQyogMdGksWlVQwa6aajzMe1RgaIfmnfGSCSsUP2C4
xtxmy/igl8mtL+pGBpGctxd8sGKer0xjFldGa8X+TuGT+OkH0uZkoEGKBMI2
Id9JKEkzycGDYBzbfSFgRIKpLzBZsWn6irmr9yNJUiGFZ+JB+DaPwevh4Jr5
GoH3kpkUeGWl4lCAWBEahbzqTW+LuPAFg9JlrvW17ReyTDB3/oEboAYgUOF/
WITCSli3aweNsAFUxLMLRBX2RaqA/8+r1skaDWd63O5U7Uct0CRXSekIV2YG
raxFlAvAEBKNuW1zih8I7iADA5m/Ep+HmX1fAtX63c4qUVFaVO165Jb8jBAa
lrQg48D/ijdQn1NCft8VgxiEhB94jE5eL+nBEZ0NxcZl7AeuU1HET79v0zPD
4lRZ4Rp8RAfh/dk/nilZDnG4VuSSXqEbPQ2hykDhUgaiHQM7D3Dle2r+2Wz4
MPW/glReLad6Uf4HV1Gdc+Mz0NdprUs42wbwHWr01Of0zV/qMqG46+AnjDv5
ZnEr5ioUqc5Mo0hF9+u5Ehxth1UymaIuMAvBwotz9s3sWUO4TJay5yd5613C
6Upw2/M2+tqf5Fam0jce5oAEmY3nqi9Dn/Cj9tc+aTS6Xn/tZWwXsf4g9lLW
qF43gJpWx8YYv0tT8xP/h6LkZd86BgF5FX3DoV8ezRfe4Od8vNrO+VM2+UMd
hqaZSmn2/q0v/vyNK9QLtocfRFVCJyJR8CougndVbhFkRTzKFzkCm6gNiatX
ji9qj7aXgNC3zRkxfX1EFTuDZOv/wYIV1fmeS7Pk2l1zYnrLQkyx4fkR7TIj
n/gGZ/Jk/xe/J5E/wnXqkGpuDCV7TQDd3KfNzi82NHZQOA90ErHaC8VUqLCc
bY/bQOCoTxQG/+wUOj3S34/VYkRjf1UQpnRuhFHhhLZl0lxhekcd5zdePIxz
EjDhIQ8xyA993UeGOPAy2rALP+COiOnbVh3QAPKWpyrY9gnyWTQPPh5sq19m
G2x/9+/brb83pC61s1Ha8dYtiZsDiasCBbZ5dG70/t9QqjHj59XFt2JDgvLd
GvGd3cTJ9Mm+sJ+77gBjUkfc87m1ore58uZS224J1ZfvFvbYFz0tF0p2mFHl
90CEbMHIGG+4tP5463diFDBMAuuGySXY/g29BR2gp8JL9KHrjuTefJHS7GD0
2fmVW5msvw2nc8uCXlkYJWYPqBJnUxUYTRXEglPHVzly4kzIwwxfBWHsGpn2
zwpj4GvVvB2/IuQ4aW5Dgd7yBK2/v9MtlFYVH6bejjTP76cVNb8m5stAuio2
WoL/Y+ahIuduudwDWsNu3zJoKP2l7PXrW7+W20VKX3XjPDS42oHrBpTZRPbC
+GA5wOebCc+aThV/HyNuYXHKD3n15pRUYrfbc/uKtHYmxmq6blNrYQYVPkUc
0I0jzLt5+6vB50prRgq1DMz9NXD8Dqll7VgxJ6lSZ0b6bGLZVkPO6zZtJ04n
S5xMbKmzwkZhQT6VPPNPhv1sT5rHDMhhplnCHzdL9gXEwDlrlOOQXvNV7E5W
YPC8AfBUOVppqiRd7vEIerrKSz9cux4BUjjY6eEllrRQqbTmNkfsrWzc+LBk
JJO3JudywhjAhU8SYuYLoCtRGktlGTWaNz9q6Jj8xcF9JesKUJqm7lC6zMbB
+LQ2U49s4IE2qomtUgyn/CLysS5YnbEai8D6p2b9zrxjVzaA6yshp+V3FQiQ
dXg7+jdXa+1x2vhDETcP53hj5bsfm/5z7fSxeGJ8/D13itNh+O2PGqqRz7gR
JFpXXXKgpnVuxVlvw/YK2J6hm2ZBDkJckBweR9ypxwoRN6i8rzqAfWVe3VKR
QUmLc+OJFWyYPyMI4x7nG8tDoXje0a4LAb0uy4QELeBb40t7iNWTESqRU7il
PiyLnAg7BqHwUOnQwg/5rJ4ygJFlA0D+Rxv8bArWsampIHW/Ae3GNBX2vP1H
5GUvcDWYncahvD23yAHIYNtxt5bUJKEYlkLZUC82oxaBat2tZoWExw6rP3ql
3XzVYYw7rIiZ2/WZgVWSctWpKWvrozOYW15hc4FM0T5HZV0nVXt520AaN7rU
8dIrKJ7tq67zc/fFKZPmva+kp2YUWEQn2Ccvzk2wWnbMzRgZzIcrTWt6Ek5V
7RvCpbeRjtlT0X1NUbZ6lbZk2javelJSd3ItsbVknvswi6n0J8L/wHlea9p1
BoBJZHGcMHNbEe6pRlGssF1ZQFzWpsLwbnO+bNgiwsta1SWd9VSrDGQl8Twm
mKEDVP8bL0FZTaPCNnKrye1nk5EYMJ9t3G58e96oLlx4IU8cmitzq3eTP83H
He9VrI14XPOXFWDDSuHu3GsJdxJOBY9HcMJAFuumyckYOv2MTw1WDjBrE+ji
NHZ0DysSZnZR+ouIOR1W3vW7zcQ/yMwp4+1usqjBtmqz/KZLnKKWv3D/qwYV
F+rTVdoZr07nUn+r8N4NDguWyZQydGxqRQaFTFImiOr94L4Ow21Xa8mA3zan
3SNxu3HOZ4lVD2HoU3aFcoTw5jsjhpBAyP8kXPX7xmC9nfXBksEsYDDaLF8J
Pd4Cz9ruUCp7Ye0RXaRUwejqinjL4+qOC/dUYiaswvMbgzGyar1Im5mTnt6n
uPS1AddxLr1CpmCdkfZW3Stp5BuBLBKIOTRMMM1QsL6yx/YPzqzcT49ONiZV
9PIKo2o/RvGx60txrLFqxEenkEyY+krtE7EiWgrzoG7KNO6Nt/bS6vd6G9Xg
JUs2ypRwSrOFIMk+BGYP5wyHT4OcMQ3ntlBrABw7D5iTh9fCejSX6+zQaUO+
B6ZT61CBDrk88zPGZpZeubPDDnS+N4zo4sbnJSSioSACSMtJwyXqECAEMONY
rfnBmu8h7jir2ydH/ZLIyj36O0aCGfzmnBl25l4aSTfvZ3nqZrU5U9uXuVfR
qXAVlLmdqUbFbuMLhjk4T2wi1APaS62t5056DtB4V21T1HagUq0KlQqeAqLE
Qy+DBOKCWi5nOzX8Gbz11XjugSbAqZcKJyLG8PdmoyOAAnk9LNRlnXPfpfH+
Qj20wmeIwiWKI2k/TvH1b7pwKPO3p6J8DncyPchj4ET89qmwi3ZtaSgfcCsR
LDxZggiiYcmkJyxe+eEmX+Zg4atF/cIPmO8L9qYWy0mYoXna1rhnMf+EYKzW
IicDVDf1rE/+bgvBefgkqjuV7SQwTwciVfDqB6kCL3FVS+7fah+hJVEFa9hR
KSwCwrLCNJV/DbOoSQeHNbiCzJnrBtWPGHfGLRQpcnjLNDbSKxyy09tS1Vy4
H5PJDcuUNCrjh0mQaoy0YtnMRoI9Y6+k0Por4x9q9WxfpTj7+gECT7dx30q+
eYS9hcgKu+p/rgnN0yx+hLTnkKRsNPnfq87rOY6abpF7WZ2HyciMo8OtuhR2
iJZRhAbA0ANu7jepZ0tBS6A38SWSTq+y41unLp75LjH4ms8twY4PF+xjW8st
Ysif51BguH1yiFVxCT7ufq7cyXyWlqUnxJ8Q0f4JJPySSJFWl8HoTjylCntG
LnDrKLceQh2y3pJS2gqgk/VUspIVC57t0TdCfS89BD7iKVkEBLAo/a5RiXVV
G5HB1O8JWMDSwZZ+K2l+SzZyOA9lhtlk1Ti/FQa413t632+BLuu8xW6FBg+E
ZdgBVw8wfGR+/sLu2qX1qmjYlq2Dx+175pmdqrXGTfx9zOn7DQorbUnFfZeU
tzLbDhOlpZfGzb0fJYjX2/bdI5a0NtyzRCFNB78d5wlSrRTP6WpaEQ0DVIjB
sucVQtfDVwJFSaLrhWXyUKw549SauEHmDw9snFLGycdusqWGh0jOSKKTBS+D
khYM4WyvWa1LTCMvtZ15HYDYNyMLpSPtzumeQjBRNEpHKb+flNrEXDvzOUZp
epIubFnQD9+wdU6pHUh5zC1uGUaWJPB+9GnJdWy3JS9iVeH+Qpl+tyrH5G6S
vKzZQ6oXk4BTde4C+O+tl1htziz88Y6O13BYN2GICcAUw1/yge4XQK+9JGMk
545U87mWi9jbZzxeRgJkofgiWGauZoCQOG3cI4sO6DRRXDzIFRAJoPiosCIz
XT4aEsCZsrtVc74d9b/IxhJRJEe8ruvh0NaT8nxn8xxC3JC93mkqx8ZvaIC2
LatSTOu7m9mpyxU4+rCxOuvrCW0PBY66J61VxZzTGesBr4w/7sH6jhFToeKY
zNsVGR/+COuM3kzBZB2SxyKfe9IjTsgo+NcpKwwZgqJiZwS36Z+zag+KsBYz
v40tUD0PXpK5wimRP4w1bA6dBiiivCJfg59Sn8An1qPKgPEkkuSvGhqEqkOy
pRvQ+NHyQ2CuP4XE+XFNzPAB8X4XUEzijt9aNvzTMIrv9BAotHw42VhwrXfc
S3Cbrsjj8H+AyLZltIrUCJGEsuKUmY1JyOs60SqbHUPXQxxbh8lwlUu+1HyG
SX0cx5Xj9ISFRugddnBbyI5+2qLbv3EXY2EIK8Q9orGMd2v6BpiZ6SlzpwxW
Fkzapa49IVdBmL5KySRxtUdyVkBL3HS7p9mttsxFicnkLdwzDL2W2r2m2dYD
TqL/8OyqN5hvsl/1Piyl7ntKd52hnjcpk0SRSnLHghNjxzDIXlSA8OIUIeHW
b/4OIPUGZOHGTFeolkI7chld9UGaWHd4EcOlctHaB/e7w+TD4eFJVjQ65cFn
PqveAHMMNge5ig7P3HAl5Z27B9/4/xuNMyTFD7D3OIlci7/9OieRF9ShRWbW
lv/wZ73LXT46GDtPezGOxh1lPS85j9TXCAwi6gjgYlqvAFOZenykJsvDUOkD
GTy3qoXdmBWAY2aFlq2tWiiDWLxN5sGL1k8HAat+V54iU0Pi8YiWWUK41FUi
jsNcl5inDzORDvDf4CyjcCSagLS6UPpDxc55te6e03SBJleSeQyzoOb0/HPy
Dza0DV+zwOqwxL0UdB5fgPG/clU+RhzPEN3zP8yjv6Q2u6OKagZqpDSBYl1L
uE32rVFM7S7V/yRjTMojX7P/QsCkRFQKyPxXlDppiA41GMO0mhGlyzw3f4gq
zkIksXt6KQzh54Vgl65MjhMG61X7a0c4onfAB3zhdo/mwzTbVDv+Yb8BB90s
isF+vc+qwu0lfVQhx/t2MtL1yLQp1auvYgvfKV+5RLR3u4iaNOZtxUmj/bHf
eQOkM3Wjxdy9mX+7iQExs+iydV4BZ0Ht1Afw3jYEXmeXe4h8lIMdfa4h4QUP
SDcbl0jCQaJNJpNfuUtatCezzw5O9nwYUVDrD1Y5KNQnfqCnYNJ6GGWdc81x
EYSICnz6AyFqjT1Qvlsm/JiU54vwGdwMUjrvE3If1+gW7Xw0oQeL3LvuHEYc
8A25AtiB7vjayjKsEM0EXy0lcxnmdhNLxitDUhWpWtlnrkJs7geQLj5iEs29
hrUClPiQok2xlJbl+X0qB/NKG7yGxdzXfBT7EUFSiYpo/JYDHuZOClVlu4On
9DpHBiCqjl/jfEFjfxhIrRXNSCEB17ZtLNGfD7ZYsAMQ1tJLIYsWRJ+BOioU
zIweQlDTMs5axJ9asTURkqjlHEwHDA5RtX4eDObfDXCqO9eK2LOEs/rBeRoA
Hc8shV0oV4JPhlj4VKG4Yqxnm37stWhNCP3Dn0PB8ZqmVsWSHGpeBDPLPL5P
im3pBcTNqGESzFPPlSPf7qx9wDgAFy8iNYLxkeCjldzgvu2+8TycvCU/reIG
Vn4/9Wu6RNcE7Tr7EL+Hlo9X7nb825KDSLbr7OxCFzi5uzb5fF1R/iyLzu90
ilKbZ+7SPPWPqOh1YV1hsqHxp10a03xXY8AwzC0nB3/0p3kTGSgRnlE4Vk1M
VHIVLUxBiLo+a50rzuywBKhSerQN4eHYuu/ahqGhewisKwLtz5pth4UOUk+x
X5hyznpGrHS9JxG9tcbGUardLhdkliVlsQrA89rsqk3iYf+y8D0FaQPRZiq+
F8Z+3uNtXsmm4jXIWUg9fMfFDP712r/TVn5xbofAP42yQm63BRQU3wi7v9CB
6IxKPc4OFhWzwle6Ew6sZAMJH5H126PFDcr6d8Ng71dNGsm7N7LAjAZ4qSNd
7BqZeNrOrG9e3J/g8u5Fm/rKhM0XB5KUzoqIfxBQex+sNhUhq0ecr0yXfrMc
X/ddbsURStC5KhRSWkEIxLHZY43a+rIEKqfgpkpvTzOTsOO/dmQUxeJ1Kpg5
qi5U85Zbn+H5l53vJ4ea3eltxFrlMZTR4vNCDvfmRwpxU+eH9vMpJIzHoONA
O5BU3Vc8F0w5Zkr+7oI5A0DdrmSfP0JYQFBM63chjMCXTy0ab+WDOBHVADEs
r0ViFJ4SHTCya+TjlXCtRP6xisN08383EDPfnA7uPGP+ZYUVZl/1xnAcylFb
PWuqSgk86Hptmm3Hkkp2T9RVxvE0D2RBhNT3XTTpnxLZN1oIJiePK4JCRlgv
X8dhlG7InMvbSeqC+HDUvFxI5T/b6ai0pqovclCrB/+mvmLmX9fwvGc9BM9i
RNlexeMYVZcpzi8/0XAaVDNVfjCu+X+JWZSj11k/X4d90MXyspcLf85fMz0K
ChUvZA5170gf8Mxl64Q41YLQ5A5EpHGwT9o4/W+fQ2Mzc7BNcWNzNF4k0P6Z
LRiHLgmOltwid58AN8Dj52SnyeYubV6kgq+FSqLBTsc3IZWwSFp07iWx+p7x
V7m93u4YqvljX+Riv8UP0bOenIvE1yYXXifK5SwRQo0USeIJ+He7ELBTukPg
fPWZbsLi1aqgQ08TOZSdlkcF3o7MKK2p10WdgL0ba7D3VKNKXsOMIgwz7hob
1kNZlpu6irzF47AF9tJbPJOIswjQorkHhcLqMCg7Ah8C0CMnePytkmQPDNWF
l9SsJI1imZ3r97FBmCDFK8rY0guFgr3WnFpbRjwuMUFP/PMRgXEfQFN5BCQk
d91Pv0MktelbQs0Ig1h18KrOm1tdC4hoEC7W+O3Hy+kudqT01EPDDmIXVhyC
GuZ0mjz3pZqP2+v+wC9jvCCelmj7H5CNsC69u6KS3KlJmV9WdlxVFH1kcqf+
EgC5meO/jSEEiufRMJJioTHB5RQlPZ9wmlc9HX2iPs6B0+OMznJ1SMfY2LVW
Sa/fUokJSm1Uds1EJt98xQN9C3cxckkncm4NW74xH6/y6sKsma89D0APQUJq
5jKqwVKn297z2I8GFZ1pIqVN7QQNLDuVETnkUdPDB9jZdxQnyQ6eoeaMKb/I
cV8Oa57VrE4zUpkIZYRpZMDX/70+CUzeoE3alyvKY56ic7gKU6G9cp3lULar
Bksp7fVo0bE6M5WbBs2uxlKo3EC0o/2teAWAeJ3Cd9HLQk5hZW/IFhbO4Zs9
PwEPPv0rSuKfvEt11FylCn+6cMTvlMwgtR/CjV9/MTcY7i8bePI2qZWus9vP
00/7XKtuVsyb62NWiRNsJAM/8f5rHU6PYETEygn2IpFfzd4l7508Uz3RhEqG
CbkUDugXpabYzI68qbMMOkNIEola9/zRKwAHTc9fJil18jDCanKV2Ak9fz3f
Gxub/DW8hejW6CsZpUT4mHd+KucpDvi+wCW7+RzELzJsTiFgabO/kc/vJReC
qATQ2tXXAhHBnFj+U2KxfqwtgpA79zz39qNU8kWeReWYc8n0/6/8TbO6d9J8
SH/Q5HPMOS4uE7t3WAZRUxAYo3P1ZM5gboNtaXlbYyhYirfzvhvbRnJ1NPgR
Du2QiP9xHXFDrVZpq/2D8xUjlkTxQ3EhsiZ4pZ8ZHO7L6AKWgn+lVFWVQsjP
3ilSgzWTbJ7Ih7T57ZKpTeQEm3LeQjRC5YTVWmsZ4n4HSDh5QiFbjUfywSrV
10WZ3Par4be+bKkSudDs37yfgTZ26FrctnT3f9Qd4Fh7rj6pqxoMEwOXt8Ec
1OXSjp64JYu0F8VMQffhck3JSvQgcbyIA15ZT7NLtPmyQl1ONyPyfdxvj5zU
dFTh/DWhQqpI/I6r5b/ktPWT1xd9I0884BBJRgz8btjHGr1Es71j4QRAkOcY
eWYKdWk++ZEah0hV2aRSTfUNqk4r10aYPiWMUhlqAloo5nN4fnnpY/RicCng
qjXK3cTLKp9KkOO9ugVwB6oWQxOpwy7MHYkC828INCWwWnhy9uxMMG3GrsEY
ZqR4/iYqc4mHjNShBJ1Fo4w5CBiW1nyKM5CB/yL35Klyu+ILWpNtQZAFWTAb
QdnM5fdVFwXPrlCZpE3HSSh2Cur1N/2vTELARNQzNHUmJcE8Y51qP/2fI2NN
WCJKOryiOerAUV4NnywMfOH2BdoadfFUi4fT54v7MP/hT/JgEAwI2VK5LZl/
8rWdI/fWq/9WmoCaVHMMufN59H7jUpHHQuOaAh088M8myL4rj4zSKMJvc5am
9uqUXliqDH/m9w6TNCJS/41Z9sE64+7mF5elx+0WAFfb2FrPELD1TTqpFsxf
WLHeFz2pN3fyvK24fqFFydky/5tMqHDZfVnR6DRke1XaxpHRXW7CibFT3p4d
+L2TlT8975Z2FAEg7RCCG1l/tXxzyVL+dualyIBn/PBBwGCv0KljXEmGbqnI
z9wqZhaYQmlMy4Yb5hYxifB7K3p2Lk1+lyM/Jzl7r4QhO9nal20D4JT4gxCY
aQdz7dyRZQOkVmcacAKddDpRH65yxoGhfK3eay0sTyPLQUYWruce8Al5323j
qJO0ThS/K9RuzyjV7lFUZUwvtMmZw7AJh2i8hVxcgJIrpjGxhdLXH14sd3D9
DIyJEQQ+7RmkviQE5TO/1dGy+co+LKsmr+zmY6vmM70cnqqnaLLnwxe8Lbru
jO7ws7PnSlwzoA33GT85ADXNB0E2wVpHEPQb0ORqhtyPMIzMrO8zWTV2LXHz
i2BCGdCMa8p8jg7mu2MMvP9BfmQ1lTStsLj4WdmHY22A2b1XoietQLj6pVzE
ozjI2OpdZNpIRgUWe/bbKCToTPsFLijMk5TI3lY1Io47tyrTFqye240f5d7q
4F3eIhPynhUNEIUBMIXsRzCG8hn/zU72NVqrFsL6Uk9/WmM0GbMV+MBQapSL
vsynVgmLmdy5FEN+JBxcTcBDSJLmkwZn4kw4ACeHwD6DLslFJIO/tX1BJwsU
kPSj6do47aAGqBWcWZtwESFbtM9DcBQJ/7oUesAsoamgU84GgmI9zNoCT1MZ
dFDBo6UIaHiph/CcRqNowAuad2Upc2pp7EC+U0ouSNTZH0zISK21gxQtz13a
/5O5tEzNlHoS3cZ1sHPWuzfsoBtsrWiqJysvNOUJbEBz3PipYYQ8kC4IZYaV
9xM/ehzHZY9CwG8O1CGwhWWsb4niMjPfuP/FH3OpPtoS7qD/etVvW5/SD7qI
xrpBoHo5bjRoF+qiAGV35X19Xb2yQ38iOeHSwca+zvkYwTFfT/bRxYkO8CkX
hnWwgQJaOysrTFz9idqpiOw039CIALoA1ep3WP5WWOG/spIHAVcb6TXE+7Dd
ZH+jq45+AgF0Zt1ah9Obwi6V7weBZyjVmv4dXd+IKlfsmRY5vXYCH9aBVbE4
0nJNhuiQleZ0JUpBXftVCFKFHuMm7byaOkQ8HlFs95dVLHsNeVFH3cPK5fwG
mHR5saspsZ6Sz4V2fhDixnaD5APy9uJSgqTCLLWhXEXdDz+AldXxf72P1+n8
rTvjnjBFLrxlIYSRpipMSMv8nCnSdVBdMv5ssmrBrHe97vWoWeuxwQA/AzOm
l3WH99/Tf4lki9Hh5O7Z6WWKCGIl8Y+LZyEDRWv65Rd66p/3T26MXHh+9VEZ
hbcm3sy75dwtdGCiPfXamZyUd9cNdbeKxPxJZIbKJusKJnT/4S/qhNlopzwF
a8oAeeZDTWI6zKWDReygXrtjeq4V0WYRrTmEVqVt9/3rvdkH0IH4PAyagfyD
/tQjr4wigLs2NJXKb3bEMs1IUlwWYu08aWNh3PSpS17cC0NwKVpONRaKkX35
lR1bsIJqhA4lBQfSWAIAGtY+S+2UMb0FB9MYhFkVBTArNOJuJTomaOfUf+vb
BY3rppErI3mSVRztxrjq74bRW/CB0qI7E98vtB60brxVm8+LMdo6479cTqXa
0IO+O2Wem6ive5Dt5fS9l/O0b2crUCOtRXyy0ZCZ9EjOF4tj9o0RtKR7tpVl
JRsTLWt1qnqBQem9YVCosXjH+Fz4tLvzsNhnRAnTU5Yl1zpck4k0z4G71qvy
hSx1LsrYi7Q62xkh84NQmL015RpBnyMc8eAU8kObBDxA2sg8OzDxuTpOQM9m
kuMgfipNlt2/fEHNAVJJtLgHU8Wi7DU9il9d6/DRiYWLL7oKEa5tpSK89R1w
NdgWoy3X+GxS30/7adnnwqnQwujaQytnb0guydYF9EGv99vxDAlMc8LXaIfO
MwQJxzI/Y6M1ysu138C2hlt9L5bg76+yUsyVi8akxyXzweV+UhE2wKNhQIZa
dM3WFYdrx5sg8n7xsJtzbIXXGN93HIX/DnhHbGsfVRDS7qYu5h3WGnLdRS3/
QOxRH3j7yK6cvtEixVy88u0F8UYFPWLip4MQxat/qk3WIj7E9D0a5itumHHh
xWdZ0tNjybgjmt9G/wNhUbrWBQRQYRyS1cfQhngDPflgvrso4uWf0eLDR5u3
a7JmtyrwpESjBWVFfr2WMocTNjgyB27IMWXFsXICpj5I28WY2FKYJQgJJ2Tx
hMvtvNnLMrScINNVBsx7htCtIxHnghB/FmOrng2Axwx/A9Sel6tLQkWEzQVR
41dAvyhsrHLksSyd1gMTkEA3HIKHLmK8+3r0GieWI6/xK2t2BY91MfWpOsWL
PI1+KcsuhoWCmuIxt53dfwf1aCfL2Ab+b0M8wQKncSQ/NwZlcVhnHm+Rp2at
1Zbtzz3s+i5+QJ7NzJyecYtxjlGmsWM7+3ZwJKotwqD9TP7O5UTU+4aXatKt
FSv2lL2OtaIu/Y3cLtDOdxtJ2ZHWO2Wf2Pj0j4Q0kNdFeCRATxTHPHi+pJ//
m0DRuiiqK6NqHAuawYa5560WHQdcEgPkWVQNSUYjEdG8GUxcYqNRPN216aZ/
gO+fajH51XJTrVCalet4tNs4ClUMCentEtrYwnMh4KsVuX4Hr21LfxbBR+4u
adBJjumKz0mHBC92IDTJuVmlD3Evsd+1xkCBedCWN5HS5tevbPy5+xfCrqmp
CKR4kc5v5OZT2VJqbCHJqbdz4rWHvH2Tq1i5U8u5A/txScR2vLUCHvKbaI7B
0G6EvS5Y1nk5gwJF1mAQC+cTbZDO/iNyuE8qYw9pF4RNDrNXjBkpefN8pVj4
FeYxUUB41KoRWnVqmTKp08j0acAk1T10aQU9zdOpgM2l+bmwqJdbr5VJ/3AJ
UQV8NxPKsH5oy9PmKhO6fCjvZDdFaUXkZofGimW/i5OMLv7iIilz6sfty4lG
ihYL4W3sGu2P9mOQg9GCJ69fmLB16vYQ9xJsuRpEuQJplMHDq+OyF3qj417h
vgsDO2MUqBHFCZ0I0PrQVzR9fsEijH5Uyq7XFcsNVJK+Tk2Uq+b3h+Td68n7
1JbMIphdFAdcy0KlB5j4eBYmzaEHQFT4HYbxx/bFrtEcVz/5pIW9rAGqdcSs
wc0y0OP29NBQZDdUnOOB3aE7ZUqTXnt8sPQLrQwgqZa6RWqrrNTkH4sjnxC6
+MDfuUF3lqpnX19t0VE+2xYgrcfrh1HyBJXjYFjvDEAhpOAQSzXmIk+rvS0I
AaPin4/50bDnbob2E5w/Fep1XcQhgIsfhFo/GRUeDDjt5cDhboo3pXSSZNj6
QSozvz7+rzb0Kw5cNEas7dSIwMDl+3fy/eDG3/jnXocWPYXaBalUPFjcE5nF
AE7d2MalokTPpt6Srzp6biwW1xlD12xOpq8H1NLOkLeSik6J47KRlWZWbr88
hwRSGNPeGw/8jsfI8DdHQee4Dsd2y/pbXMVk06cegCN3cfIHiB+JTQ9mmNlD
63vOrn2sqOCLt6UWFRXJAgeCkPs2qmzLRWzD87CP2oMoaSNRm1tZ3XzyL3fx
LPNDuvw5BRhNpqG3TAVn8w40vIBm2da1tRaMbbQrl+Q7ixopbMDmJk3dTFwY
AeVSLM/vSy5418PRWX9AUbaJbucN7l9mTSlM6oMkksBCZN5EqToPJ1Bx5azK
oOYIl/IDHHrWqVcy/EU1IUabG9fxf6rVWyqpLmEcxxaEnATcHKDhdPypbGcH
iRr4QufpH1ymCiDM43bP5vn/TCCbxGqcXB3l/6e+gQNmKPmp56wT8XtWpdv5
n3lzJM6KwtOGqCxoY0Mky1SXYAaKmGPRbhM+v1De6l2JCp2O/LVzAvvbCOz3
gYdJ5KzT+39mYvxip1YN7qBJnu0wF54Pf2h31XD1ZbqeZBOlCitOWTwJ6XvV
teUTV6d7tsHD9xiFJyV0BDHwQ+GF9tHBrUdWsDvLda0R6d2pjQ2zf6i+bftN
zrf++m1ngp2prbkFif6dN8bUX7sH7XSvVkPaL1cS5xB1akAtAI6KRI6Ymov8
/TlePZcHM6HPp67tPYSOc4H69XQggVD0aqJskSsUs/8UjKXXABfyUDdVz9Vu
EIoZFZeGqJkopPePSB6tdFyt89wq0k4ILl2pu0WCErodlFX4TTCtxkn1p8pd
Vnbt91tP6A9S1+5sqK9kULj2S74NYAKWHhz6bO8JOcReg4fMHvN5rG9XsBOA
inR4sHLRriAq9XZli/d7rPW8/c3v9c8uQ1NT6x5J7EP8d1aLLFVbfy4ORD/6
mjshR54isM26s7g0n0r8t4W8h3k6fqW5V3n4A4CVL/pKjovMIAN33uAFpOZ1
cdAPl2MXVhh3MUoKVxCX5FIpeypz2x1NuyOlfowm4QQt7Kgul3CzC70T0Hdk
NQm8r9DNE4OfI/XjMtm+uBZjBC0FWLozb0bFHTRmzi0RvN72DZHAa5uuODsh
L2xS70vToHn6ZV3N51KxhPDWcAaSSloNxf+GYPegKNheRgW+vzlUr/VhWa9I
9u2SoPDjS4K995LgbG0t1atS5naS4RB8Q5o5ERGnjRnaZaBSfsXVGxxTM+pj
oAYixfnJfcGaZtlKIy5Fio+N+Xt8JRZvfcNC0oJmxgRv3QWNoBw8a4z79bFM
JcM56D0NtdqTwSplwZpXtWAb1lw6l6CXwj88iMDtn6Gs5fRAP+O48IO7BDRx
fIoD+vrrCJV0tA9uQavtFGDZ9qelaWr6s05HR9g0wzxmMWvl24ArAa2am1tB
AJovUwL9YRxynszuFbN7zKMelL6Vb3zdjjcqqUqtNDf7ge422rabdOMbG0P4
OMQkWVB5zt8ECpLK/FbGN8ylcUUwbYvrX/QPbm5pJmfNmSx1r/XPvj3oxUvl
cfZzxb99MLoJ+pxjzxqsjFvBEwEEuHsZMzouhVv2c9ul+U2MSwPyNSkY84ul
V3On8YZdl/HfvqJkARjDmhscMuYGeznL4kz33Dd2FDAQetRF3Kl/jOL7BQiS
iNsi8xfnnJpIHTJWrIAg6eTaGIj1F2BwWS/pWcU59GcJSy/h1lrdozEZZlTS
1S4okonzu6S40NaCxd2qBe/JTMY08XdYXXhAG2dg698vo1YlwrJoWNSH5z4k
M8RocEwYATzCcKrUfz8nBqxko57q0W/mzkDY8pRWIKK3cI3E2Uj8O4Ul4Von
AOErYl2KN1hEWBku48s4oc2hPYunVLVQo24LVyGOQHAUcmo9qlOhEnBSet2A
WBXXN+p3ukJZF1xoL4uaAujTODW+z1E3NfsfZcxYIPA+BDCV60ba3apjNu/2
a3lqEquDTB73YxNUSNQKyyBPOeKjXb3slmA68J6R+z8i2+kQOLj0IAPoHS8U
IyOEetJKB0iwuogKdzKtKdrxp6VsM3hPla4w1MQzNYITCqh3E+QaIU0/R0EG
ShHuK4psWHJcjz6bpKefWzJRoagR7EYv6FfTIBIt1d1CMC4DCfgaVYjLuHt7
W++ZHtoMP9tz2sk59Gzn5oUfLVUKPY906Kjz5OdE5D6vF2t1/SGOqFJH9x+e
DQh/s7D5SXTTVpy5RDl00+iZdrp/4SnRARzlRFBRmULDTPtOV1TW1WsXhDAT
x4Pv01X164HTa0vySx9gNgLixQHCF6L2Mj38yHDnvlW6eIWRVmSRlb6v3Gcl
F2T4HmvPkvV6rLI4U0niXiUoroRFxPqtehmcCePwadvwQFNstLy/LbKNV30U
Ny8HzjrIAURcgOGbJAZqNuzzGxIB9ZFUKkGBYDNRl56DvA1b5EnyY/VPHR71
NKKs+1AHytyBDKNPLVWQNWRRuLhTjpUlzkIqSyzAndCXlSi85HqHFBJ1kRoF
qxG9jWaKcPfybG8v4gCfqdWw4Zjj37yJw1Q6313GOLpK2Jha/jw7jUW8t2TI
P+ocvX02RCOJvr/JDmlHxi0Pg7LLxAflhcLaPWi+BnvtyY14RS9FwuSiKJHg
rCIqylyCc7YVEb2Ta36G4yR4x0z+vB1nshLSgtkc80Y/bgpAxljAFHfgpBXD
MeNYeE0+YRpEdA8zmAVtfcd9HrXu5URgFMjxfHNtjOmF/ElfEnh0erflklXv
zwf3lfuVpbdIf9/VFIeXzIiOSQvEmCWuPSFHgUupzEkDkBeps725RI6OEjFG
6QSjEpeN+r3k9o1qSxKGtgabj3HAvfDF/FU1pSdiKqp1Q7G56BCo6TFIsM0w
ctbgoMYfESkq/Zt4m2oFUkEwvIgQ8EySnR2elesZFEglm7aOWGlLPD4pa84f
qVXf5lYcp4j5ENmQ74MPjLAXZeWpnfwreXRNGvUo/RzHRL/xwqY+oduoU3gs
Otn1Di0BYaTcEXkayc4xpxbmgOgBCTv141SVQcBCrfnTDmYPCvT0aG4VsBYJ
yuSpY9eNkfmWyUu6GnqyI/pdkzEv8Z+145Ub7kSBB8tLsA/qYmC0uVaMJs47
zMY/GbZDX91oZEjgXUUiRh9rBf9iaSLSON/XMwb/HNg/w0UvrcWRXb2Y8m1i
y0/wEXEbPG8Ri/FZHtBb85qJhLYVcGUHu+QBRmRasuS2rXGEqK+f2gIPIK/n
xtlwNgVKxSHUCf32WaUxmwvMxnyXyLfFwAQ0IDDvTfPtxbRz1eUPGcmiBBOx
BMMkoPm3HqzRjIWTm3plFsbM2Dd6jZ+DuIspynfJxv5XuCL/BRmUeLDwCcRR
BTtsn6/EIMLNAWlcwrO9u0vE97n/A29noeDFhmZC582R8zKA21aPqU8YvMYM
bsVTUdzFzMlIgNx583S2NSXnPyf6ggv3h5UeHpBqujDM8/5d9mERwRLPkzUc
xFoGGvJ2E65eAmtEmqB+ABWAfUw5B+zBWVuOGsXhTLozIOzUO04X5y5zCw9z
/JciAauUzXVCJElrK8QH3U92Jf0qToXc+I3zU+CCed0e3IuWjRe8VVNPQeth
2m7AIv3RwPbtgm+uJvDLPB2hzHfnR3TBt30agOoxP/p6LGBzPxUYXL7KpvCu
JEbHP9/OsYQw7plaWOygoYpWwhkYWWNV9oUGfeBW8HiOeR7K7zwhafLqgFKc
KMqsc975v/V5q2BcbsjVrtl7QjhYj+fIxF/b+1AKj1i3KtnUSPlXvugSEVXf
QxGKdtxocpoFkV0AX712CW+inZlmf+4YHPCjV0AFe3bp3FRbdtil2xOymvLN
Mj23AmB17NslMIYvIpcv3qUXG2zUhmamUc8KpIIDzFn/GWHL1Ityi8VAx7X+
aD8v/OoIdolqLFJ96JW+3Kl7J5D0lvjTGInEc69HN/FaIeP0p+09YvA9iXB4
wUmPQyQawKp1sZyS/DA58lkh//fDnve0XXryrZ/qCE8CJWeI9vWp0JustDwb
tYdHQ4Ec9/40tiNGDXXEKXRMVfh99k8sqvN5fzHuqsMzUZkz2nrDs1YMJkf9
C1VNqn2fvfrKd8a61cOWTLc4KyKDV1HVXkjTiWLNBWUeU9uqxhAsONSH1tft
47b3mHPxGVqeeVYtdjbjQmx9KrN/AQJZ3U1Ds5NMQNYu3ByMWMDLoydetTw2
i5sXw2xHxKUrY70jWPukhiI4rWRFwDlV/lspKFXvkVI/cUbng5wNOTLGXZs0
WaTXoKz2NVSDVQCgr2mUxmFfeb54L1Lv2ehtWxNlIKuUkl/0CCpOrWrKX5Xy
Ikjf4tdKgK6IfTPtJOtA5l7DCjJYPg6uVJtGwAM+1xTcfJ1EIySZZdGY6MUz
f8bZBr1z3H+0IR4QgyMdvIhxIP3+URkacgzLG237Ddqgb7r50R/6gM62r13t
LywPFQz/t+OpN76zjvhAIPV+Idn1sAZ0cTQF/r5Bl+RHULq+NCY3YsJ04hRk
TdBXulzNOBtmsjZQFvPyYkBdTpt5CJV9dYMTqB844C98qWoDUuegm864vBYe
lLYTgRRSm5tGH0T7hAzxbao88K178TY7iEsNY4OGv2S9BxjFnKEbYtSPBbu9
4aLpLPDtk6N4e7hIvKmR5G/jraS+S3KC0u16riTmIBmBIJagKfBCrTFSPqCE
TQZhXPCXmzodJuac987laj54OfiJgrxUWiNZaUXbrb4Uws2YMN/wJmzE+poy
FfHOXN7TEVFsSlZn+4M9RksGwZXQItQ3A7Bn9PiGgwPFYYMTzZYkm8D3LxyL
KlwF3Eeinvs+E3Jj24syGDVsyFacN6J1ggwzqy+JALzUJ3ttAc1U1GxlqE8o
ddrHdwE9kbgajJeRiEPRixcm0qJr73TwFH6WBNLgl2aQn6ff8gB5YMVPocRu
9d7B1agm57kFxq6C2YM95226CMSMmi9jCJPtSxIDvhFGPH99KAo5blU3mHb1
wzlzlLjPfHffKgLSLYqxZ3ep9B8/udrrjHa4gPbKZevx9LBzmVsBt2pjYYgg
0PsolMJyTSzmr8WzhXI5CzSNRhq2u5mUehFG+FeWbuXy08cTCMUnux3vPo20
DSaWJ+g9iNGs1OtUf3QGB8bJanapuh0E1jTjpM/JR338pSJ6PIRUl+Ql28/v
FLPu6BqS6fI05K4UvrbSV15mmrVDAGQxIiqErn8Z1G98yhb/2X3PAtewTDXU
yNSGZAw0eRJ8C4ffTB8F9+31a5zuuzwCA4fvJ/pW6KD26dXDi387FAAj4VqM
asqd8VXbtsL557fzkKvPhXq7X5+zGWJc28hnQysLqqHvy2Nsn/S7Jv6lbIRW
S3pLo0WALhXmZJ+DPr838LRqO8fLWX9utVmrW2+Xx2iA8mGlOrPeiellwzYQ
vVQ/czGrmsNBGpppQOe3rtfTlhX8qFbEv5FDLZDIbjHaFkaXPcLDBvBw1JzB
Gr+0WZy4Z1A+Eh8zZy2OOwm3qlHk7eTU+DHCWS6D9OczuplzOiOW3mEh7WOT
tNdSRc/UsaEE68f7eXeEyRbCHvZGJTEhMzOpD0x0ffd22wdLNGLdRRNSsQuj
Trz+GTsSa+Pv6MhctQoBc5oEvaVvljha+uRQEg9BiIFBLRwLs+xXBxaalmsB
Nk3Y+AEzwkiuE92/Cesq63xxu+7Xgt2YAEBBRS1k8nZUkQnenTeqMfjvJY5x
J/gSMcOi+N4jLatVg+1A0zYXRIXGg/4qxbWng6pl0HOozuLYy8YGii2l1wL7
3ZD8DA9eKmkx8SDsweFUVxjQRxuG4Pcprt+uQkwDv+YJaKsfpOj2hF+ihC5n
Xz/dd7H0hXcXLWZtQky/zVqqDocJoQX/Jhl7JpzglvZhHR9qkiwqA5bHTGrZ
x+23m9wH8hxd/MPDC+pu32Bp8ZZhjs5/ezmM9gAcktPHiH8ZYg/4aZfcLAyB
8n+wFDRhzUGTDaZqghmS5icggquEygLdbBIZXSMF2FQJfnt+85pQj8QMZeiL
RSb4nAm1fXCt3RlY9zcTL4eyAtrpmB7qc+AKf38S8qm2ylsvRhlv3schJH2c
PxFVY52qy0Z4b4q0eENv2651lXi2O/wCI6jvzUK7/agjH6tvz96CqFAg94v3
WtsWEvut16ksfyoT9sdhZb1QQ0KHhwsGmjCIQSTGLpPtwphuTWzbFK6ndxVW
xhkCDbDpD4HWqSNn5D7/DA/rjkQcqRvnJLYlanWtlWla6ft2PuN6/vrwcdn6
zcZiC/OX0p3J/ZXOoMlHKnwM0DDFIattgEpNIcALI4W5CvrUxdPdtaBDw6RY
a9liKI1eLAzd6eY696N4F741mReMiclpBuNiUPG9ozyd2ReBiEwEElfXCfOT
U+28ynDFA8TNxViIEGsLUtMcmFf0yNV4+DoZ7mQsxlEafvUZLK3mcKC0Bvuj
QmeNNOTLSeFC82uCtOzPu16J1lp+g16xUpIftT3fvASQagSdA9QG8lb+KqRv
dTKWxDYgQ9YGQaM2+3yxeVkmplT3oTshnYm8Pcn8m7FCsw3U+ZZnwMLuAz3l
3NwG6HziMkQifn3ERZIQbpxaJc1VEOAQKQbtwdJvZjxc0phrwRyzWgCbVmkG
D3tNuVlnHpNmuRYiTTQ7GkEj8a8A1XRSroQW87/WhzceeLGcxzxi/v8tzh/b
M3S32OAIo/A0Y4iZK++1W1iztrrI2S5FYViA+Cv+iHqniZV+I8TjB06OqT2J
X9g2pt7v0wfhs8/kpspouhUnjMYyHW/RDsLnFph4KEKs0UqXq572KxLYQs7Y
DOR312HfpcHAMwesqNWpikj6+XE1FEX1JEs4euWFvaXDGJT+QDyw6mHFjytv
6nT2Bf3YcPY+RT0nIOlvNW1XwTpIV39xA6ay40kMPy2eXads3C2SPLlVZk0Q
U6wsLCvJfeqKj62BSzvUM6RJ84oRk0a8xjxuR4SSvDy+Gm6kFC082KzNWhH0
i1QSm7cnd2IbLy7JmrhhUM2iQYsfTNRuehiaEoebrQKaM99Apr13ti8rX0WH
VsrLopWFdjVK2B1ZgAzgkfuQz+g8oEI3cUm48hRQjJCALSH1GKWabav0tPlE
lvl7KeUQqqvjiPzdadohnqyKpDu7Mc9a0F80kstLbbnZ67t28mhoeA59YlSz
OPC7F7OAazHqD81mwb8xbcoPf/498ErYxmN8cAAdl7vJBIIEB+eXHiHFbKjM
+0JiJZf4auEbJrQfHBHL4bzHkOS/cqec1mqrumYtPnDB+XjtlA7DBtmjt2vg
ykA7vDWIRt8wHa3AxOJ1X4Z+lyFni893eACVNps00arX8ck4yDc6cC4hUk2E
LF/KFFaau5hlEaq5LFKsV0AtLE530q7Rve5reMWDp7FWmKgJUXO6hhsFQ9HP
jUxJX1/mqqxzciPFeIXlV2W53MMNywLaw3NeIJC9gzLTvMDyox2ZpE+jMUSJ
FB5RDZRWnDzY3ICmGjILMYmimWetm4VkTkWzGCn4LAkZlp/fR+njHtf7Nj2M
9dXKqHpC00gOTGwI/X7iJsswjlM/BswFw9MrmREmRuKTVXd9vsAkAH5JTFaQ
oW7CJP6lbwPER3vTWhPwrNBzFXxidmlpER3BhqIRTuqzGB2SeSUbmNT/r6mA
zFXQkGtV8a5IuFzQrcAbpOPoEXSmiOZbFb6h1bQIjTIeoS1eBhk//TPauw1o
GfGDFxhcY5iAxqRjZasNHITBN94Qo5sll5DKJ1UrdEqElXs+j+ezRGTn2ll9
0htvmeIdmDyNN3+VfEogJydsjqX8om37UXT6GjW0O5RoFotX0kkR1IhfFdGH
9xSy0a7fKvRnCGGSFQmGYY04puit1juulqlF/bR8zv47fIXmnhgvoJRYQScK
oGT+1o/OHmRK76jlG1d9H1Fk4oV4AJl8hiCTKlDrjMYxCqRapTfCPae1FMSZ
Pu5fXXkUs8Vni8yEZanPEK45pJAZvOmVfxNFym5c3TAVNUmQbzgEGV+dCpl3
1ppV1RovydkxiJaLl+kxiGiiSdhgvU4GZO8ZNeAYzs+hEAdrkriZKsgOrn1o
sygzR7pv4p398hBqXLiR3whW7Ol7M4/bfAnvb696Z0XwCAVc8lWuPF2DKmmu
xtFTCLqGVzv2Ca4gNuwB05tJx6qrJQ/IBDoinaJBJOngNDV+60Lu/tNexJB4
9xE9DtfPrbI2EtqpZIqnI4U3Yz1oZBrUEuLDKmYmsjb3tRvY1vMEgVzO4c8Q
EnBxbvr5v5SSlAuAPocAEjpmZ8Pq7NuuToT8qG72hEfgB3kP1BFXp7cy2mBv
Ilupy31fC1qx922TmSRvbMAdfW22RFP0ji63MoaubxesSJNlZzwYYrF6AF39
IrhF8RZpgwSXQnU7qziCrqmieQqc4EnuFzndbyccDyHM05CDsUJt2sOv+S7F
FklQ8il1cQX2w91W+MkojVp0Ohphsg1gtt8YFbywl+Lr9/mYlk2SmbnSwdo3
LXavpqaXfvuEVFCxSI6gqj7GRFr7CbMAYjpuFU/nJ8HOmGB3CYR0Gf3nh1Ry
ecIgZNbTGPvCZGBWy2R2n61yikWT52TAUceddcSJasq5DSDcw6LydsN27Vv8
sLsrku4AoC9WqT8zz3aSbEdNmnJ3Q/CedNDjlYIGTd2MMljVh3XFmfxYP7WC
gcboAZew+a1RVudefqMviKY9nEqclZRbFUqEyrqh66kuOC2s/Jn4wxkMPoZ1
NMOl2iBcoGRzm3ItwLJ3wMFuALSWTuaX0olKLNEHvVSm4+Y1g/cKvYhWpP4h
bdw5VO8OXXGYDBnXyrriG1KuUuBdz74dtpwEtJNBYFS66fpywjBEEAOjqXs6
j7Nc/p5j9uN/xObgJbPfGHW91Aja0XiAWirVLgwwwPX1Ls8c8ctBa9S4fVMC
bu2+bmuKA5Mt1SotWPkq+2boAl1SclCIGX9BAjNIzw94+FcVfVp6pafSEaoI
Ud7K+/zl7/63+u3u6v/VzFPFhAZ/iMiOnIgF0Y1CAIrH0eTPVVJvNZ04LM7b
KA/OVjkvevmbVavqwoafUCfSoIj67EX+q4AnFMKgJmhvKr6WrXU2NxLXd1ak
jjti59lUZSxpdT7Jb1SyDPT3lowSe649J/bMJE4EEiE6YJqsGiV9e2LFe5Mw
ZUg6N8W7KA46hLmcOwiZgKZzkeny9J8xwWWGplcPYiSPFpkPYkj8P4E41hEt
ZOBRN/8I6Ss+rog6Egz+xBZgijzB/Wwg1abU8gb+7WRLm9ti5qViJjKo99EN
fyPjmgTDcDHLFARMnbOxhv8VoETHrbz7RFRzJiX4Gg3w/kpsB705nZsGbR8O
99bc7eWNuDC1GNXGS3Hugq/v0OszolhHOtIeJGjmDDaGnLseisFI7IATeuqV
HZDU4MMmEgmrPIoMPQjOIsh2HBzxwEhVE9v4dalnnHPSnkf5gFY5L4Q/vrum
OFHhVRZZrOa0f+MSmQVXqKOzWupRlEi6tWM1ZPz48ps5CTWExLWfQ4WUa11j
jLAVBqTpMlxk2bK+ByM3G8X/RgXt6BX7f2ahlEeYpameryrbDykE2+J02rZT
bNioOd20gSfyqOcGLAgaIJIOIWgLXhOD/YhFaCCEYe/VKx5//98FPgNhx93L
f4/oEMvcu5iHfV0gdNCGDYKI5CG2GwxPS5I+GrKJa4Zes+Hv80O++f8n0npq
wJ3hEnF6HjY9ptwDFJmTs9YJ66Q08GM7DgCG0GBucs1MI4zs4jAqbayIYrpR
0KV9pQqE2NLVCzHqfEBFPuBBHJA2BCjS/b/xW8J+111cOEOQl0veRxhIZDM4
ewQtM5pudvrUyqflFR1c2ncIaxCq4E9+FirLISLZoLwH2EcI6eapl1b5P4Jf
1ccC6vFuxJ254Fb4sD9wK5F8i8o7J5ry2XMkfKsXT7DJ7bnLoasKNXui19/b
lzY9S63zdW3/BUEpxlYzoClM4AX2JQVOFqTCXqROBKcWaFberTbd3chom87T
SoROAR2GcuGmTSzYU1CYczQDoXj033kQOLF9ZhXd2cls+ucUDrbvqnwkNaeT
MmjvaiqxxD0qVvTJHgkr8yp7fbJU1AfP+DUFeoEZyxDmkp+vJrTi5FWhkF+C
Z5hnvmJ2Jk3y0AFS2UO2NYuKtHbB+CqAtuy4x5+oiof0bmRg887b7FfWd3lr
HvHPvSgupzy6JRN0NlRQ+rcZ6ay+/TS7jYU5TiKW3CqfGTk03Gp7fktAMIW9
BaoLqrTdOa4r4IohEQePCHWOTFxq6zqNPXIsaC0CBWtc1wmbMwi+GPmev9fj
sYxFd75RIAgCwj+jSY1c4iYhLfkZVGJXlZHKE6H7/EaT82nrPA1WYk4s6GXy
Y2e8QazQsSxz75lIM8t5oS7FL1iUmx1QS48FiLluqcxNqGNzkl2psHk/aNn+
fcpQwBskwsSdgTcwr4/8o9YsBWKwNvJqXChqYEJdiMmY82MdbLClyrT+9UrK
CX6RH7II0BQLJSR9UClOk3g0ZDkCKCWjDUpYdsVaZ0Do7iNPhye5LSbNlpg3
thSnFL7MNkZ3Y4XmO9MVtANMjVjuHbStx6bq/R46MQmn8V361iOEfszOknlI
iLvSwM5dUEK1bzsR0F1pWg2Bk3ZX458fFX/xcGFUt8y/gll8SuzNyyA0H0bs
DyGNxdR5rJOIwa6MB6jJKMs7/w+wMSVclDMzp7Qnrku9W5aXHvU6OjVrb0Pc
+KdxDP3BxRGSrB0/HcBp/80o5P5Z0yazXfWtU2yzIHBJKXCgvJFYfpQaJSpu
G4pd7qFn9rY0MuOUsSXV7dYu+7B2ur+3aNIItZgCDkJ4HHYvRES0smmp+I2d
m5BAt6/vhq6SyBvfhnqom2mfGR0nbaSWUcR1Xzh7Kv3bRbCDiw9Uq+HMbkLQ
BX2mICGuLYo5/1lKFW2fJdvudK4+uoaItGj0+C7qwTFDbk0h5mo0FUmlQQ5d
ocYtWdR/DB/Qfkmjw6CVu1DQY2HucNr9ZTl6sCylZGSPiAUtn936nJF8mblv
7D2S2G4PCOVpN8PIM7xgcf4rcbnHgpfs+AMNP1wiTUv85vBSVKSybzzgt1xt
WCnjmI9GaoZZCpslJXgcgp7VBK8AwScE1dDq1iXvsKFZm/x+xm1TrPBhPzIV
P/Vb49zT/VOwVacC6uUpM/ZZHMh48kuXdSMYCZxWbTNzY7xjAF9Bauyn8oEw
UGKgSzQbGMlMclmqKF9YOY8DEC6E687HoZmg8lFHYJ/yvEtY7y+/QfaqlrJE
YRjUustSBZB/ONotWDu/nO7eTW60DiEECEaYcRRYUgXx54PV4PqsJkQiQcGH
1OJE+Y8XxBc+WsmhL5c1wEuMPMhrVetWqFUlqyaiqAxCYZkhKNn/B84KxQvm
TRa7kg6B7qSghY4VpxBQz7LpSsbsmNjhsHejo/yHzz4sYi7Q1cVSbgW0qCGW
ME5NsQpGNpfT/egf2RJYexqEVWw8II8jq+PulrCfbxFlg8ezK040fHBC87bu
11urFNJeAgAv/k1mKwU0sIKQN0/Fp32rmEcTXJ5ONtOkRx23iJlHKidEbVmn
yIbzIfYSmZC+/fZy4UeyAgV/dgaVc0NWNnkmnR+0ve6OE1RqPbTQ2s9C2Htj
ZnFqe3nbUY/0SToOqwczp+CT6GMHT3CjIe/FBN+1umLsl19SMuLxaEDdbO8i
xKXllfcdSkZNJjODPRsTQ9XVMHguJPJJBZ76QWVRpfh0fyMnmd1B142umzvW
U/RFT4KbH/4VvXFTCk5kv/gmV5pt35eWlJwyEh0C+tvKah3d7vRnuEu/Ub/M
duzEbsxHXnqtc2RU9Axhi49RVNt+kX7zQn2Vab2KXP4cVpAONEuVvfwZ4YI2
hPy/ynuKb8+byzR86BKeRR1fUuwU/0WEEobUwB7zU0QivtOgwJvuWa8G2qBv
uvVIWr9AWc17qzp3QBSyp0BQ+PFVgof4DQ6z8lu4FV3hH+XUSU/3kEvXDlCB
Eotwcu30R3GGuXXgko44kXhZ5L/8o9gC0eVbZs/jTpjCHuGC18pA3lxfowPL
HxstfiCrDpw/SZkHkWe0yYAZYMWrlKGtRaN62X3by/z+M1p83Ij74SJFztQv
G1ZhGQaEPwqvCdPSxF7Lvgc7OaxSSnwmVB428QNARufTupkg8Dy3rErU/tFO
XDGDHPdBmmuN75UAhtoo0INlgRyFgxJvxaOORzl3K9lPwuP1vosl6OytHB3D
JAMV8ynUsHUtF3sHQ1zE66PC+N5uaoJSR3Nq7lMxmEPmAg52LVgvbDL+SfNY
S1xth6aHjdEz/Et+iSjOuKpDib4R9rJezNRFogoTmu2R/a7fdYkOx5FqHxg9
4mIleXO/Xv2aBbpdaiF+UwNqpsmqCHmPCPjhn9IQ6vSQaaU5+GKTENoSIYK9
xX0pyHp9bNu4sPBXJ87GK/dUfJM4Bue3Aa0RjFZbSg9BX1RE8epA+ttWkDUj
YgTWbtLGmnJJlh6IIksxl3lnpkz0QKA1QBBIRi4oUvxyVYMee40ctiaAM1YG
lb/9QfS35SylvzDbcc/27d4Dlz46uIhOM1XtOlvZI4mlScoXPhtxOCjiI3xf
980+dpENcfnGrLxnxMe914R9NWUCf7HEpKJLA6r7TKSRLc6c96vAchmekVJR
Mw1MPyanxwY2BZOOisSbwxyec4KmDzCZglcNYV5ITiBKNCfLjawLok/fD6T8
4vRp+PYjsmTqpBg0A3YLYn928gExcVsUI/pBe/s9rSOgnsDPLsymHN8hjIk8
RSY1lAvMJm3kv+KOq6HDvqqew/X6X6tyWncqby7yzZzG3d3WaZsTt+xq97uz
X1eeGjehvwaiS0oVmNNI3DM08aqV0uhxpP4OyewNzA6QXqMRARyV7DptWPeP
Z4EQ/Eu1wau1Z9uLN/Y4/eQBucCVojrS1+7jPXcvocO0ZgyzQX8GlE4GID4O
WAVGj5H3d3AGkqeJ71D1eazAUH/SD4nIjDxXAoTNbpmi/d3rQtn4F5W1QU8W
r0+BhpC4uJ4v1FfSFzHsVTQ8+dtmw0hBn5Ol11cBHrNr3cR26gPaJQjFvycn
sbNXOI6NePstTBj3ytPnahwCsXvC9QJvo7yefFD8a8q7C0yVzER0mw0poqev
55noYTq9dR0pEHGCMqGxI+UoBi3z2HA8TbCh2IEL2qBBnWQnieOA1kee8eF8
jAjVYzVbF/yHQP3x0mm8ooSemVRSIs52KhRzugXmNQg5jYg7QZ6sWhcurLIQ
sNsGYQr33rz1lyJ6LyFESKerDDQNOYxVKY5RhhPauuu3fz0nygzNHp66BkMx
M8R/Irk8Z3NGI79H/CJ3f99xaVl8IWXJtE8r3xeij3IQziLLVf/oLo2EXUJ7
kuIcLWX0C3EMq7YAe1qAFTLqFOaI71p3FxS4qZa0Go9iEuKLZv7mqyPwYzdS
Wy4vHcZ8bhHWO1XWEDWhj12tfNFYlZFH+lKfK2A0o/tJcrDDuWVpdbdUQRwL
Vi3iTeh9Nj6YWtydBwPjg499Ae5+K1fD7gWTtTvFYxl4hTl04MOND6/vy/kQ
7TjsrKvhMykunPDpy24piLJq/GWZxojIEhPFdYq/kI2ls7XTxfHhr95xHJCM
BwY1SeLhqalunEBr3jcmYJTMSxyeiIU6Vglr4zMjvOnwnQG5w3c25RwqDuVX
UkR0W6Ho/MYBKjtdQ/X6u52hUw5S+BgpbOnzFKLLwhPN2KWSsxlq+9n40C1b
NdXJuv+qSDeKnRypzVNTIaZVIkkX6vysGCpfQQtzvkRCwnRbjkBw/+jcFmTH
WPWPLqt1b/nuM37vDBoacJI2M7xKaO0Qo0CaBUHtnctUvNd1tqdwx03tS6Xz
ZmfKNhzSeV/9gXotTljyDkBo0HHyHLl7F6aMjIYP29T2DIVlcXkhXhXcbjfB
+F81INTtzbGksoikpt9epl7vMkX9cq1CTLd4eeawxRxmWye0bv9dz/AuSyPb
URpo5MRZFiWJR7onvfOlU1NqHV2PpdxQAghFpAR7E6PmwCYR93V7Qxprybz4
nZkeyVK1nZNeqgt0tXFl1vS3Y/04SLx5rw+t6aivHUc0gsDm8gZI6da0yZHv
rhBE6TN+P7QDWknnUMmGhDmi0uIgat3daE1xfB2Nk09EyC8uIgAPvou4kPTj
pFjSfk0jWiJipemw/gzxQ1j7nx2EQi4ksUaYQ90v4Y0FJyl0JQYJn4Ik1Y9/
xqEYJp09HIu4tXRuAofPscpxzRQBreCFhZoU7m5MhZvi2bV3ppG8Ks79a+gT
SVFYBMf2M+ausW+36ZNPt/b53gwIAmwZuYjfL9nVR2i/X8FxuoLLu92Ab7Fh
skv9xE7346LnGRtqE56tnTkdJgPLc+JvN8VPm5fIJSgs+qgjwGdMg4LHYNmo
1E2mzxJreyEgNcnemHq562TZ+caR7tSIBWLvf6zspB2djuBakF4k77vjAmq4
8UHwNnkSpFKaMd63PQtKrBHBM03vCmKLA+xGXGMGnvQ5moFIgXXM3Mc0Fx1U
cEZ0rg1b4nUKDO9ZDA77KxjZLNfStCwWNvBRpZUlcGTTOZpq7YWxJsbKzwPz
cfPD1UA9m8yNQeN2tnZl7GszLlpZIXpCjyTF9KpuWvChrxmzwBT15euW9poO
QEtQ+7ZzDytmJUIQNSc2sMKO8m03o+lumUumVoe0IFv2/ragkTXmbhJ4m5Wp
RHrnwdNc2n/H4P3rwNt4TZqI1COiBM2JshhTceFjjoWkxPvSZwWe5JpmqrEr
LxKYM8+gKUltKk3uPEiFVqREZlqNsooRFoKtmpUFzdsgTB7PEip8p/xxXTNg
l+PHHP07W8IXP4rVJycYAZ2SNSmZ7tgcI6pNTY454b2LsJKDD7eTBkmIFUmL
y/+TyEvqe6u2jns3k4Cv9vGoxKfULH6aXQl/PZshENI8plySXyFBtwP1mFEa
47ObLM50urXMUI1SKdXKbz7McoY+s22dB1s4zXksXIfZof6UXTXn24V3J7QP
Wio26msvimSi+rqmvvOdGPlaiInQsrfUYfrwUPIp7PvesYf30QXx5hHMBUm7
lRMASanvu2CcurwRfOjONWK8ZMoDKHJ3f4KL7dkXkyHk9rVSkHhk2HP0Bi7g
nZ/lqOrlGIfhBUUrja1W3o+zKWaduBpSEudBI2nWEYnvM3OUXgUjFBsNBMwV
AU3CtjQz5WqJLa2VGtiqKM0wkKeJf23h3buxP4vtgDEgZ4JzDzQVr75D6v/a
fQKDZeWxYzikL+w9ku8Im5xTxz1qbQn2YG0ZL68nwlcuBswc/CJVpGJywmki
o/JzB7NPq6ZuquaMYMIuUdMVxbpwAgsU4DZo7krlMRL48ihFMXCcWS9RzeYC
+151P/0ISgdhxznocpDC9Dxz+YKydiqvTxJuIUhC1NAiT8bXmfS09TUo2se3
q0UMfqz7EW9LSrEKIWK02h/M9DMYzIdUGgCb8j++ExaatL56kV+C92CxxwN+
P/zxHjZsHFlubum601GvzsYan/8haawLGMUUS1pXTcD4aSQV5UBAghXTHtEX
jm9+d63+d0JY8iNHpPaTczaiStOyBDVBgN/bh9LBFT8FwSCdxdfc3gzDoLwi
vm7vKOCXe/almZS3RbF+G2i4N4sDwDcCGNI5DwUyK06pBNmbAob7DK9uFiTA
P0cgodkE2h9oIKCwxj/WazXMVRLOPwt5R0sGb9pJLjQnpHaN2Edb50T1ETet
ZkS3PphoyMNz+jSKGLT3/1dXvpiUQHtKkQm7CV36TJkBh1lnwLLlynxZvtdH
D6epU6js5aFAR6HWqm0y6NAKtfIwQ2q/hioInDO5f/wzN0zkrhvc4iMRQ9U+
WHYTjrm2PumHJ8UnpFnrWJZcTH/2XeuE1zEGxLhRXqbyrk10fdd21jGVuLJM
gE0rdoxyn/V6Qf5WhCRyok1rFz0dNe/LKTu1Q5AQ2kLsU8Uxkkq/FXF0FWMt
gKEConreSncbqc+FHUU3cKB66p1sEJt0jUpk9l7uWbJ/84oiA1l0v4uSH31G
g1zmfbwJtyvqxDl/EywwPWVFQktbjeQgzvQFjEfNTUlYBSFv8Rq6I+nhdTym
P6dPtSQDALqs9+1WdaAn3OsixA4cWpXSzsJLkbgtAHlB0DH+S5B+631aBh/v
c4sLO5N7OxWTxdJR5M4Hi0D3vU3a+3gBNCUdehKUwwvm/ltIn05FzJ3vEEkd
gmnH1Sp46XBEGAYV96+IWYErRunEemq3BSyoo75SQMi5xes5AfK80bKcW/7D
Ln68BztSh2vdeDbOUBNMhxcOviOit/wqD175ixxPLliXSuTPyguJPLbFQfzc
seWnKDjX4VWyHqtv0YLH/9vXd/ePMsMlCqiUNbhHC7xk/Bi1Hp9854jRlCyX
kZXsAjDAfXP0t7fgZSHX9eMaxHxILk3Hbbfaoyagfht+Sf9FvtHve6nv8C3r
kvd7NZR5TOHVxohf7I8wRutck5TJb5p6C2heSDVfHHDrmBxof9r2T+GWdJPz
DrHzWrPD3C+aHN3sRx6UBajzanHndpAaLJltZXOI8T7mnPzN21rXagKhte9c
GUZ75s/vaBs4OLi+5t74cCswSqJvxMsiY+mnUFVI/UfVE49ohg9dHmatT/Zk
2HJKj7xhp2rvjCSCq1AMQcAr4jymCStHcmo22bd64CJ/4QO3Z4Badpb4+N6C
h3oIDeo+QtHUxuE5kla8QeAGos7AolK+9LAwikY3f0e9LmgS9X7RszEvOWQh
o8JI6h4rWy35tKwCoTeijGqHOIlrSJXeR3TVaf2f/y45TIs4llc5e0whGEt8
WAXy27/H3KX/6SlxZu3gXlHBsvHquaER9OZgWeZQ42e3ma0Ud+BSHuQmF8Li
OCLwHKSD5ghoFJTxA+HQKAkkABJr+o6SqVMq8/EZtiLXo3F8ayYDZ2pmDDk1
jrBmGeopCeXGDkGkfsBLMkJZK44FNaifz3qP+foBGgW20uPHQLbXJnqE8VJ6
vOLBsriXSxd55gdw26ODjxAlndt5G+wU+tbWdgW5YvwNECak2+ZPnbdUMtdx
iCWSox3dARSSUVihR8umUiUqumAbKkidQMK7WmJT7+zXnh2p+UCtUyYqthxD
BeepWHFjtIfeSZJW/18K1zqfu6lFHFz6xYuJXjIPk/rDd633p6X7PjWc3FcE
VSLveoVl/6SXYui7JYAtP/71+Vb6/ISyYz3pUvqpNUcxkA2QvtaCrNsARJ1o
HxUxNHM27wEsllcuTEmpcEh7vI8bVOFiY42jEp/iqzJdh7yE5Yid5oqSZDPh
r9scPHPMhcaMdG6zZhIV4JeckAUgZ5NiDVN2gI/w4SEbsx1SskYjIg04kj5f
0ndfWvanFyCRs3X/R3FivrAqlMyYKzzCejuZ2YEBXDN8EGlbigbQLXbCqLCZ
wZagXSxyeDgYolvHwQNIdb/XaBB70y4Eb+0mbpFKHnrMxtPP4J7h15wnhn+I
R/i/qn0Qp1/fs5UbGQC5SgUyDmN5iEP08zwRU3ZOMJwgbAhAwYVWY1P5oTYR
/8Mi2fmbNrIehkYj7tAas0ILZXZbDkQgUx7tGEYO7adm2Rkuto6J5yTqNLbU
GTesm/jM559atBOeBkoxCmbwmhd+6cZZx/qDOSNHMukyCIXNZqPvo2YsUY7c
gd90Zmr+ERnM4cvY4e4ZwljJdbaA/cneEAPVSWs8SIoWmZWnZtbJsrULbVnT
tMiaLCm2E/q9GfS8qf8gAQ/+SAJFH8ZQz0S6fWqEsYW3RvVpZM9ZHZvKr6t+
ZQLX/7TQnDgLcMrZci7JL7IJFdGxxrTDbavwHTSH3P/2ADGwAyiXZsbhs52y
MrGGiQcKwYq/bGoQtnL+ecGDOvkiD4mbWbZDmVBINTjR7rmFiQzkI8Fsj6dL
8Y3Ditpt/Mycefwmei7dAy9Sp7ZO1ff1WJz4HU4Oy9zy3EBq9lhCMpfIGehS
aLW5H/i387/GsoffpF3sYFUnLXUnww0Ff5Bs7OSBLDIOsOit4reTxxoJboOE
UZvSPj/5RKtGyL52JL9pKDpqVTIZFuaSzBo0s3yCTy61G2QUukvEUVXZLKUA
RlqKsjUCiiQu0ej3Z5k9FqnFYrxCT34eLc8idoq3MRICJByUzeCm7SHRVfNt
KwWmnYnR8rJw5+3kuZw9epe3SE4idtqjFkeaCkT5+ITp8zKs2kzocGw2EnFS
2hpGR4eyCUrquQkpxfR3LIWK5kI+znlYN1JcQFLNJ4EvgAX8tPy3e8eHbSIB
e/KZNbFyUWNLYYvPr901wdhxH4ocVnNQWyiloVe+lv4MGasQUuGNkwlP+eMD
LO3c+nHVCYf0th7zc9htJZiihPLrvwr2UbKqsYOPExk9gn4uhzTccYeth3YE
cY6K4Nk1v66ZQnxf0LCjPucCfjfjNB+ZHnq7DfAomxqnuEu3TWTqa8T2Cmjx
hSpqw3OIVenf9SW0RvDj5Y2W/hlstBC8W2Tf3FFiRyf45eqAeOch82tZLLax
kdGicW5lKqWI3nVaAgipEXy8lxtIkERv7E2qGOL25NaB+9jBbT1sELvCUHCr
a0apc3DqaHaT/f7A/Ay1723jQGP+q2G95U6z4iwWryKaAr4vfdEZGhDy1oDK
gFRbm/ttQFCH3LiLuHcDvfAjyOH9qZIANkLJ4rWu8wetRBvhphT8dw3e/x6W
5j3i3CI1b7tptEzxoIH3mEkbAwX7xI74lTwPxP1esGi2mtpXuPFGL2D3ZLFe
4/ZKLIegmyIYRn/Mb/1+McZJuP3kjxijnbstoHLaMTe4clpRc/txCmeEodgh
+acQty+I+DNNLrLhfkwCSl8lDLWwHS+3Y6jh1otCRWKThpMMiTByHFbpWUKm
xEue3ieR498PBdgqwIjdnvY6B+nmcHpNuss1kcHJOeeowNP0lRu0bTaxHZBb
LfohqHrxp4nLBsG1UKCcjYLfEc7V2Fn+zQ365lLhOVSxrT3YrX85yvm1jsEr
blOrUK5u4VgMnrDE4qzgyOGQg2VJkgW7JktTYqR79ySiZD1FYOWsot3QkODC
FlY2DR9sIRNHihP2CzbbdQi7Ru4xQkah09lGXapMcLTiXjPqNUgSAOxwDl6a
FoG/yA2e8JDGOxgJqdGWGNjEDL7qvKFRuAyFubsUvFMyakJY9RXc+2XwZLHO
AjI3TAcFnRvV8hKcElXaYEsCMqd8djEzT5YB28k2sbKSgpVNqEV8AI6/nSZW
Kubr8xgN8QIeqMj/ivuNU4JH/DhgseRnz9Bes2SalTJ/tnrY8bVfSC+jFUOO
3zRvTricK3yy6Ym+c6bMNoJx/jAVYwYVJKS9vQnkAv9jyenuiBIvFsJKNbyd
f+Kw35BPGm1Si3A5oWojmSG/rSX7AzTczvjLhQ0K4XwCuke21Xye+vMaLQai
NnGd+TP/3BkjrQCMUPPb7527pYpeB3AR+69Cfy1oRaZUe9YomzYbycUk1CYu
E99az7fClourESaZPQOpJAwY3I8PiNePR9SEY+qnJzYmykpFPqhfFsuSP1ae
ebdjZ5izE+Fu0gZBCgRUZf5XweZnGb4pzI7++shJZCaR3gZR4AWBHHhaXo1/
YxAnc2dOFVzEYI1fATnAdCBHabbxt1+Foa/GkuDi9TFOfIVvJ1OTPiPws1IH
TB/JWWPCwUscJAcyrbclep8nf2E/YSFxHklcDdXeZ3N2oWcYsVrw0xXUUH7d
QiRxhyvFeVlePi6UdnIHwiaclx1rqtripDOZt8nWJQLY/chF+bQbBlJR27sO
2EcN7YZmuHHblpzq8Q4T2ov4xKUH/j2lzt1KpQXqN66Oq4j49+LG99BXmUeC
IPbDLBms+55rZVKhhuuY6wkLab7+W0Qvpsq056rgbzPAyo1ZW6hC4UxdG7za
Zvl8SnN/X+epPP3k3TQDr3iCT1uCh+mlofMnzL/yRRjXUBhdiF+MCS3YztQS
pEbHalFLbbZ62E8vgl3ql/AmkbFOL5ASTttC1/CU95N3kMmRm5qd6YJeLcm1
9nxyCRG+u4zK30zg1LqpT8mDY21g8JgRxfhQGECI3qRyloFrr9PyDSrDOQfn
O45iF5Tgwb8LAJDgeDhxwxuHZjo/yjtgQji5JZ9PC6aSUXV2kgGaYfBHJ/P9
ak8AZE7ccx+ow7qEn1YreVJU5S4s+prh4Nc+tNTfhYov4U8gE9u5V0I/exhX
GKPlEKrVPGU+Zp1HuPezU/RiriSoRpcfE47qKKm0xCo4f+8IxaIZdvI4eleJ
UtDLgkx+TrF++AyEO79/pN30+uevhDwqrrOEbFIkUJEwu1MKN9yEvd2CqiDe
EDX0+iXhZ8G4i9ezEH2LcH3h1jik4XX14zj0S2/e+3D3AQTTgG2CE+RO4+0q
tYVGc2AcOapzBiY3hhhfFtoVvxt5VTTCUMP9/1jo0KKHvJ0TxftYizcw+r3A
q9FjLbXY0HbA/brBZFJA3b9uDPNQ1VR9THYrRkZQyJtCZwk2otgj0EIwIa0a
uz9PvwDFMWbDUmPhLqeTO3TTZ2TIsq6WiXwz31QFY/hEu/40z4pXP+Dwi1VN
LKjx8WNvJmwE4pDAKDGDVYVPh2rlJ+qIdwQT2Bi3agdD++E+02etIxEptrqo
lYaBhY2VkBvuWg5LsYjpdY5j2UHKXlXZ6zUP23fgl228weFVwzy0j436lBHy
+d9N1oR+WZPuqGR3nzxBRuL4ySsXVFWj/tGvTuy/GzkQsyAIO2UbcZcN+KW7
aq/zIdKS4P7AUBXRP49oqUAJsolwNnL6MBPcQvR4c22O7yWVL71qXCxXHHlw
+D0pfMK4ExEfKljef8QH0Gcqql8PkxAjAdW3Ox1eAsYOw7uT3GD7rhahPwJe
BQmEn9wkFq7LN42kHSZ7Ubd6JL/LhxACEPD7TN04qRISeGPGL1D3puxcUQ+f
nZGwvBjdlKMBMqQBwGMH9iWyoAg83XRH4q//0NobniGFDHEd+VvyzK3c5znm
e/pEyTjLN2FwCUDXHCrOo/cXYTerfGsRKSFR5c3B1knSx8eE15pjyz4+gb58
8QlsxKTGlQdnUZENp0Dtqc4WVROx3rcY20ey360kp0jJPVzLE9pKV4VGXsZT
xjHCfFZAtktSS6omnhCQ6gNSWGTNCx+ip5RzKdFl56sSENWCY3xFqg3rHwp3
Ux44qFKi+xwWFQbcDSV2FagqcsD4tnzycgHJ5rKISq0fTLM31TZpI9kFYVJU
nGSbbGYn4annSzVt08kl6Tispjul/3Z/QcbY8i7ZP4mw5v/R2A29Wgo6WUWG
af+PQRmX9jSaHGPRYpKMtGSdx3xcMRdRh8Pek345kZ+DM86Cvrzj9KMLoojo
iDZS3/BSpwXEoNMxLru0lncaeJxPFfk8tlNRmxcBEdj7cCyj4mDkIMpQbNw3
RKC7eC47wB7l25Tj3EAwzQpyXCPQvZO4jsHIwr/giLZwEnZ9iXgi0LMsoQlO
ZEe3TPPO9CZQWIT3OemRLc3FGgcELcQbaY+0TPu8rf7366OS8FZbISFrwt/e
TRwFPJdcmAHCv6fQQ231B7zIKIVPgNewIblRGZcpNZOJViPEEnVTipZVvMpf
+aJx96NAeBa0wglXusOTzfKH5Qp1XkjaUCTX41GOmV0DifXXd4Q7CeQfvYgH
PbYUQjkap5G4oZkgrYs4y7DWBkau5gT3pnYSEbHTL9gYVRjnRc4RzP/22IHq
9PVhryBLAa9um5xwMsz2MTjfxSwl+W8gmh/L1eudIjFGlHMZd5cYnhUhG6he
5vTn7E4w/iktyUzGH8AEN75BfZ4HRZ4ALXPmRfZ/vhR08RX36UfX2vpf6bx/
dVFm0I75GlQo8FAPE6KXJYFFlPEgED4uzrOHu9Qz5PxaJxjhFp05dvByJgcS
1aQp+hVk2G4PCaUsFNBvoANGWz40CumWsg68ezVEjl6RzlpTjp/mM/F0MNx8
TZwd5D6PO/lJRtvfhrQSUr8LKyGUFUAYYkINBPdIvZVzFGZod1yD8ZgJ8/mC
jSRHv4N0y5RA5VW/bPTJAsdyh8yXDu5Yn1+qSq5m99RsbNCYFLs8mMkvOX5D
QugM93EvdjkFTU/mBWMtVWSvkuipUSArMtMdo0UWBf9qWav57XNgHEtdwomt
KgjrPbraCNOa+UJ4zOU8XCiT/Mjni4AWoWy3RE0nW4kQylYHzsgFsUxAuYKG
VrqE4YnDp+gSbH39+pbe9Fsnq40943T7kyNFF0oy9GxuuZ56X3ItIjzfQWZD
lXFEM7bBFKruoxGP36Cm7IP1uSTEXGdvmRN8Mm99pxkq6rzYY5YFGHisPIaA
SyMENv9Li4z1ZfCRlS75n7Sz5mgolDnNQ9m1RW8189Bv0VWuNt1CIsFLPR+n
SZd5WnYJfj2YRYZNOFO4LWj20nzX17Td3J4VDmSI76rahRajv2pSgmy0WoDD
dw+lqvNZDAGFfi9KUX4i74LsnnkGoBzPSe8hLQwvYQ385tMJ6DgTLAOFAvzf
GCGtIC3y8iuRTU4ljWwfi6Lbj05gTAK5sC5pugpU3aSAs13BYkogaMu0gdAL
D/wyEh+CTtLzQESIMcN7Z6A5LMg7+LYQqMEGAMjcLek26tanMKd90rs8shaI
5dG/M/JKoOVruasGSCwFdoF2uB1daVjO2UFY7Dpj1RhMHwrSyXg+i8nafqML
sRWw1pYQiYZaGZ7VggtQUKvIty0rjqxSZn9XD2mmEppZ6SCnoVFZxjjvuoWk
H60qsylT2jKUKk3E1akWM9ocsKUcCPYW/5uVQ7sMzAEV8qswe+cdEwSBVHH1
eemiO+gaX2SGXFhDGJjoE8ryR+yEcgOyp1T3I67VJRYc2ALwIEn7YogWbEyh
feGVhQDgYhTO5Pif/CLDKHl0JEPniHPivtbo6/Af2zCR0PWPBhFvQnjG5GW+
kMoUJ/wmXRIgnNgKIPZwCUmBQS/z1O0uLq29ORx3cbQOo+u97ucGYEulIRbh
WE+jETqL2kJVIPkaGtKVbedd1rGMPOE+ewd/LJB7g6OfumXfxpFqsT8YC1Vf
MV4Q4oMHLwdQYyyOwxvPm3tvLiY49rw4jj6wJf0oMDwDMzZvijGAxjxLUFIo
9duomEJa4GMZW/ix4qDYbIzrd6DoOBSs7tcDAoP6x2MUXi6FDS2/IgTQhTzM
JvRMgkhRB93NFcMEfQ7iQv5aM1oTFoiwovD2Onf2BUpJXaGdTW/4kIZa2EhX
DPNGnd3Io/s0dmHwgi4fF31nN6ORuejiJtUs9dmrGnN19wwPTaYhPdFI57xP
wx0xd4mMGYkA4WtGronvvtSmINO7qnSSYCCBfIhqmcdLTP6L41Llq3PWEuMM
JpCplDviemdEeC7N1SqhYmsyd54QIu3A2ungurx9rjuQmgeOYBYyv3y4tZhU
ZtT1jTwY8Y93Y2hL+9YpNrsBVnk70aZkZAtVr9jutVIPvy1irMd6VhCrAo39
uw6STY9fl3YgTqtCoMZdGqldFk/F2KyG1XLb/1PC59IOZ0kslp4bkU2S7hTY
OnrCthZslsIZzPXI1YA1Zpc31DEeJTuuLXBI3HEbYohi4+K081Wz6tpHCSqU
q9nus5VeQZjpet+8yPhsscBdpQt+Bh+6OKN/AYFKdJQcMUdCBQYG7pihYwps
Q5F2OFtLOPMoX4w3YNunz9+IhRH1YRyF1aOyIqI3LslIHEY0myAQQnv/Zn6W
0KcMv246WisT3Yhzmto4xxKG7ft9hQ6WmeXa/RdUFC2vJ9wrGCVtQ5yvO9OT
4JQO37MiDsfCvyz9cdDHExrVT+S3DsPVnp9V/PyS3eg2E4c4Narp8ppYKomq
kjrsJzuL326JlIdPq8sSD5HAUevLIt0lqaH9s1TH4FSpyREA83lKNYrLdkEB
noCD6baPUD7wl6HRMvsSLh3roh1HY04HRMwAWneSFG2PK448DUrdlMSCeOpu
qhtXdn+d84P2crlhFlNQBYAZCL3vE03eqrJymwc3hhvMQ18KMyDcXkh0lvR6
PqQOdHiLedmI/JR2VDKMeaxonr9Na7azKhGtsGuZKK9YU11VMKPQQ5zNbAjg
MBwBP4GTMhPDLTlCz/ZGJSPyoJpVA62Uu4G6G34dCatA7wcIbZITrPZK7m5M
Pb41beQXs0rYDB/u3L1xo/bJXcL9wssPa37KaBjtBqQI/bApAoGKovohoxI9
L0Ot/Y2dtNPHuJ5kT56T8kqEuEaD8rfAX2f4ysS/Zl5R6IL3K0wYBo+UA6Wb
3aiU+gNMVcC3kk8wquwGdkm68C9RMylogc1ejJDz322sfY8nDdgd99X8vSH4
k6KObtX42mB0v3czXMavO8K/rx+44LCTLTux+Gtw0wr9tCIghOjwoyZjHZjs
fl79lCFjyazVsY+B/OuR79hqjQm07GW6xXKqCKHcosukbxK3HON8sLTVOi3x
KMlUxuSWb2mCobfxhv2ErFHn1P79329ffUJFJ6sz4SWjS6MMp/N/KBTOvgDS
VCtcuZhakNEZnKBbawCJ241ATjhoQZtgGKH4BtD9REiOTKarZs/k3uCN6HaG
nS/rVFIs/X/7OE6J44IqDCW+B6+G3Cs3x9/HWOjvPpDDrU/8JyT9FLTO5kp5
zzI1k8y4UIKCYGiyV2qUGPMEYgNsFFWWGbjuRy/SdsZd+k+X74+QlxyA4jnV
jgTskRfITXhIIOn5W0cjHhiwdLHUoXa7esZgub68lXGGCABIHEXk4SnwNNi6
00C1+ffgHPbi4UeFLUTxkvKWjzAl56N3WDYjZulznVPEJLE0LFk1QHXQud/9
QQM4PhE/l0Ig8K8OXUF1DMgjyqiHpf6qOeR3ia3rIWbbE67xaCqL3iMITQ3+
iZoQuczlWqmxHo8+F6Av1FIijZxjHe88R+mGnZZQabhsJjRngbV3izRjuXED
F69ldlEVXxtpfUp5aftOpUYebeOo8Ho+L4kx3gdftigVGgIMTngwz5dgEuiZ
gAlJDEductF5oMQ7NJsQDRCgu7j1wtYRUihB/7Ud5Vpvrvnqonw3XW1inm0b
1VMbApkT2a4ekm/1tNRzKzulHfhCnBdpnaJ81cYahuv2dLor6VwUvHGBYLXt
RvA16Wq4MsWlgyPL1A8LZK6fzhnUbDBuvxYojz7/pl/v5YKpmIUhL1FSOh4N
R3uZNODkNDVuNWkHzPf2TMuqzQID/158ptJiXvEIXfJF2dKpbEXFBMkyNcw0
90Ea43hOhGbDTlvthFrzZV3tcopIPLNEIM7eXeRVooR0vv3Widl5NoUy0u3M
4cdNEON/6GO0hYT5dAEktjNdjp8VUE4VJ14QYS6GvJMoKVyBNhNA37FRj6NF
rBZ64NJC1z5cD2O3IyCm3c5dfpwlbarcIHs0wn3JjHYwviPKdsnAazvzj55/
Uz5ztxr1WG8nMqUM5n+X9bcp/d53WVWcjna/zdGaAx3P/fwsXPnP16CbQbRR
qs5vEOfxkuHuWBbJ2aQNhohvbwosKgcypAEp3WyvmdaQOszCmPF+YpEmEsz4
rvCYTr7d+YtlJDi5hLLwajzQZKJuzQM14OFAiV+z5XgxChM61lVwwGPNkhJ5
sahX/Rvt4Jr3y6PQ2yk68MeojDISH341Usiy2IzVyScrB/XS1ss2dsCcFm+L
ufV7RJ5r4Y1p13STwBmiM0W5f28xNgxTDNumIoCVcBn7hD3O9Utx93Fjz6qp
pllfsQKZOXsu9QtzNssClk+SfJH2d/8GgHkkTFWFAGfTWjHhWf2lHdG7aJzo
LvXMBcwnWegStKrubzUE4ocJCppzccDzeOlUwPVHzuQluAIGpvWkvTUrQbD/
q8a8cSm5qIHv1A/bcz7bT4je2PDqE00FoFlrg37mpRNU+3h7lnUl3Ba4ngQN
i6RjNBJ0C+aW4WVvN2G2HOGmROsKzqHFvtneMm0aOz+/TA6xyn3u1J2qIzbz
X4e5WgrUJOduJvPTyFNQ0/YhicZg1F1XH17oEltehB9DpLa1PhVIMtFpbc7d
5hSwYRo9fJ2/gDkgEzzFgBScYED/RCnPEYc2JA2WMTkAp9bQ/zEJjtVvBDw3
A9ppt+QMiDMlfrOmCRt++aOp4/Em8BY4qEw3OaTf0zSZ60BiEckeEFWbrlNQ
gpqmo+allxS9HEnhe8lq45E5w8q//6PLLYBd7JF4uBopyxUa6SN4g2fHoT7i
baWegmGt3k7jXv8vz3dAMESB0Nz3NtaEGcsCL8Tu3yGffmcP0F5/gwuYZ0qM
MqEW3DBOXu4NTneRMaeIszOHUJIhIxG00Bdd708qXIQUw7uNKrg5Cf/avwS2
15NTBPhGxFTu6Fd+RsgQc9Z2il4USuBGkK8oKZazi3EEFs4pUW07n1Ho/81S
NZ6Rg8JLl/TBzRFftsPb3cPe2tIrHAYKEjjVa4V4mmtQxtOGb3RwvMn1+xYD
FX9BQ8omjpHiKR8XU4vfIgDoxJjAUgvpC2FOnuw7rh8mSVMMUiVg0lg28aJK
Hm2kEY81QI21DhSxUkSygRk/lA7wov6ZkuGGOXEIE1cc3ZJ6xd8z/3CpouHP
Q6tI5NspVGJdvobCU8L8XOkMcuaM09CptwUqqtk8S4PgUNjUl0+YsX0gk8ZB
ED2ESS2yAlKPrJhev/xXi+Moe2PGank490AHEDoeMcGpgkjcScrgfNdcdiMU
IgCxoonssta0xJaHrlFZBPD1Kxgkl+5WLJ5qh9Za3OXfNJuWDQlEBP29XEoS
+ugtHlXV1CJsT6WsIFgyQQjNnywSC76lrR+GXFCzy3jZaARBZp8E/gQ7CaYb
ig6PDnHQhHpACYtQS9bNmNDTMBPyxUFo2Oc/4DmKWr13eQwC6SvW2DSYjub4
B3t2yRhvp2KiAUYSL9H5Qvvg/hMzbFmAdDt75Dr/MewiedAePnTX6om6goTb
V3V1cYhGapucLZIYG5EiKNYQPfX4Ita7LJF5iyyBXSqfTm2zPjCH4mPxz8xP
OGBmYcNdus4wu+gLT5cW5q0BhEM3VkNrB4ZwfxySaI6+tdUublxGQwneleQr
b6kIEkQc00vsufYyG2q+DcjJx2qEqpQ4skFdyy8uruwyl4l9mpJfF7eX1JJ2
MLR5M7Lc7KLBQ2u4Ph1JvpaS16CXkiLjz6yelSms2CFkNU79EIQKhvE0wmIN
1Q/hwr5bGBpPof7zXuFouQrWpEm8WI/uT1MeGEiRTvJgo8zuWxJU5s2hWY74
QKYtdzC/Ih14SvpBNYYO3XOc7HyzwGx2QfJJ9VDdLJLs7eK8vWgSvkgBEZn6
TK346Kn1bEKkvhAw5Es5UhIPWcDxalbDqrP9GiIcFiD4sNdy/tbQ7LAdZkNs
/gIoI7f2G58F0upNZMarFGYlM/3ACW76CH+oowVqBJcfCyw58sLahSaygRu9
PagezZSH59pGtV2fdpVMinusMhGdWL5LEFe7GH6/BhbdyixnxDWRFYj6zANA
uRhP6Rzn00xlgOPNGJdO5kmLvIVfhJ/zU0qz60d+Vtr5OVe1H5mSEHsZcsIN
pQ9rGAFO5ncRlkTqb8KV432svQ0pj4eLKHrxU2qX3u5JPqJ0WAF9dJprw4p7
HcboYIJiLP2v+mKAWStkxstpI18EcgWoBCwPThp/ARglFBS2k15ooZPpcnSx
QgKamg3desz42eeb6oCuk3EPIioW0mUUUX05DaqhBT8k4AcbOnumxZfn8NB/
CywQePqXlzKRKyNs05U5X3iGZ5XdiBVUp+tB3o3LM4mvJvQiyjiMH50ZJ0/V
HCxWjcm2bLXFK8gN/7yMDuNPtIZOluzGY+EUyJH8tjb9E8GIlDSxhX205u1+
T2enL81q2xhwein5dpqXhGEsx7dHXZov9mICQu0vCWjV/Hekmk3dR6GJ2RCE
+/lj5rjyIyEuYmB4cCva8DKmhiuKHxPXExPOKPYVuYSzEolNUj8WKiGyFfMi
NynKG6vWkvKV9nr/HrzGtZ+gaQuOx3PyASJgvB3K3h2sT5ibWKZibQ4VpogX
Myxt9XgUQopS/uG48d7EdSWJ0kDYDgoRdS62IE0oW6YmoBssRFYiFDsqj5Z1
UWcnHkG+qta6Iwo+PYmVQIv3joX+hBospFlLbA23D9Cf/xcE3Exr4Lib/82/
8RywW1ed3RCufYnPUJy/aisPA4gMunUVo1I2HPiN5alR/3Jwqhl/hJls8f9+
FvG7f/s7ZJ98RXlhnMPAA86OPVWpVqBjJngD4/U3CD4URZZDRDMUosi3PdRj
5enfSZ1aKMrIxaoQ/PfhOSto4BogXA2ZMBbWYDmEWjEXYTMk/jLlkt/aJU1r
g/tB/gPmZ4agUhw6A8oc++qrZsfZfTzJvODOVspSOj+dzLmHvnv9F0MuOKzt
x0ZFFpylMI80s+iAJkyE2QTFmaMIE57aZaoGZ2oW2ZjUY55wfxeildnJkwn1
lbMuW2B4ZrIEDLV5k+27yvUh5obvr5SeBL3i5BOxvApJ2GJOWN0ykFsJMVar
c7zBrpUjbHxQyUT66G34MXrRw1ZykNb8YvlNigzS3uBMtuw80H91J8E8ruA8
Jcvw+HN3B/NJppO8HGV5uRgc1OzLpHHCaDVrUwgT+gTmQjUWJvAyuDGaZzE+
HgzDHx2bqQPHF7uyxfdqoXvSfwScjsJCpb3fPnUjjTAW/KHKrldzcrEU8BMD
dbc6QlXiXc4w9L6yJtyypmGhZjqW8E4c8K2CPse4Kse0pyqOhSlv03ajHKrs
hrdBu3pOBxlnbLrRtfXV5gv7915sW/Yu7dZ3lEcmRClvkZ7Dsx4lQrdSY0lL
8AiT1mSAdlgrKuBCjV5+xEkizZj/DbcRhiwi/h3XWpPnsMTK4juMbWEj97YM
E+LEM1Jq4hgY4phdDbRye9DDXsMzJE3qPlW2G27JQ+M3/S5Aj4ti8Y6ylTg8
0BdNZhicvRQFO/zy61UwCl2rOEG2nttUXuPQzbcQfygkCBgiD8jW0Lb1F11J
x9t324S+YUbAHeZ0rqKStF0rQfJimIXKJidcWqYiLzK1mVuKukdQRsZ1w3YW
UEXEjHX3aM4oSx+IEb/arVcT+2W/heR1tcjWJNn5StjjOtSul2jSKF+tcAi+
TeiZEclvbhR+k7Z4rY8eh01bT3LEf1UjrUv5jFHiV9Ha2b9IYLwhAP7h+RuH
p8/ceZynjyu38rKQWh9tBD/IywKK3DFDjK7eg7b9vi9U8WrfyuFuhxM+MXPu
UA4og76P6pKhRt2vDW9YyxYMlc9Ks7XmDLPwTob+v8JxbNgxBAiYNWuU8CT6
Ilw8dPqPOcuUKHGuF88lX6AzKumynJI4UE37KYueSUpFxbsL9T+u4lOI4vQq
clq3qyJ+Y0bPKWUC1b0DQSIwzxjLOnEbg018UWF5EzrHff9gjLmh1eJgCfc4
/qqyyPDk73gaPymifl8MsY6MhlR0utOJWibYmSaRt5yEL7zsnsunDSlOyaiT
FWCw5RXl62D0rreauP+FgYo52/JU3/mDlN0/5YGeqsgzZR7IrY3gkLljMqws
b2Oew0v5VSKUIwXj724Je9Dd/xYb3UdeqtBu6/0Ey07lCKZUMyR1WRi3meP2
3uU9fe1Y2DKlmtFFP+e6I0beT/RKxYXuerIado4S0yMIzQvJUGSmvpU8B7rM
hrWIPPcYajxyBF5VjAhWcvPiTgEOnKyztQEqLATHvoHHbFeET/8PmsHt/ZQo
l0SS3nGFpYTP0WC7SyFEcijSptYZ72xsZyWhR2liEXSHSPo+NZb9NpK9x1t8
xSYmKq3JQzkkWUuMXDtDHTuTK8xQtujhLxs2pkxsIXpszCdVAisG6ukAi4ab
3doEM8lfIYOcOjGJBkHP07SPCQtbkKPpaxlPce6IsOoISNvErSWrA13h1+w8
dUHXHhntkeZyQaeHTL7opvFoSCbU3/eA4oeSMWPE/dt9I+3t66YNR6oeVSEP
/8O2VvbgyE+sIHlXIV1ok9CwT6wx+/S2Q0LZFIPtHfrl9PPVGHBt4BQcG+0O
r3CuYE+yC2JQolB3R9SL2OKv1RwhHpQvi5AIOSKnf7FJ1Hu3wyLaenP8UfmN
5zaZKqNbnlENp6nzQwhvwv6yn5gcE8LtSl+t7pXwN1fSLAKjOnooHcAS/fjw
lK0SA9wdU2b4xaeNbZiJIXfERlUVI1qSJ/K/pH8emXEmpo0BvaiWlQRlrvR0
E8JbukWV4/Rkj5o+p1GitxNLW2+tPYvJ/a9O+h3XMwj2WagKBm1zn2j1Ffob
gONvrbW/VnB1XdutMFEHLgirh7MDNxZOG9np9BDaF9gnRUiwaJVZkoLirKT+
lfLqAIPx3toXPbIE3ID2TdNRY4a0+thjL/pn1iD51RjIMV+ATWCE2WNk7TcH
Etsux7ziXC27AbhhZd/nTSeyePVR+tC/akIOzdHG8A6yGXLqbIXAgYP0HH2J
tcoBEBRWdH0dGtferIiRdaM81roJRahWJKZlLOeiJHLmZtsL5TWj/Y8vfiZA
22i04/Vxt0fZuuP5bg/Yld2PsvxiO3jn4rJWLPFZpDRRIM51dW2dGqE0Z37q
GU1+b+vqYnqMy4FNAySENNqryz14yGSGcgZ1LekKOCj/XphDXwuNikArKQ9J
gIEIYYi+ziCpSh4yihduUzeXcfyoHX/2asH5uZW/6s7MyeFoZt8rn6mnXQ8q
mcMtmzwL0kfgPg0R0co/EHIfZDzV71kJFLEqH9l2orfXmBQ/eq3W5lQB0V9I
YB5xGuebHffBuBehY62Q5L7Ps2aDnEs5J6zA3/ndBKGlcq/pOq08paAjM41u
XdZ/hSaAo43jw8CZeyH8Inh7UALeyeH7L7uKwk37Bvakci2i/OusXJML+WDG
QmWIxwgH4F0JQocxGXV/DvpjTSfzt9n7vRwGkMNNL5Dfrb/TEFvGBHeHZavV
e4cF2wCpY0mKp+iIRNBORBXBeQqNWBSusXoY7j3UnmMXyRPtNXjOYNqsIMYQ
1CBuDNBzX6nuSk6ksCFh/00BvdLDdmfb11qQ09QY67/Y1F0b6XrToX8nYRRq
otWPtXKnHKb54QPimx8AJ4XTvaMvGoi+TY+/kbbSPSjvcgKftz+Q/VSceVM7
sESywkXXrJrTu1cR93bBOGMeNwnOEr7B8Eda7TcosRuT2oLAgirKC1Hmh5L3
31jb3cPCQv3azAHxp8sGWFOku2cnAIJEdmGj/3GPw0qqqRA9fZFOlrSzLWex
8Tzy+XVXwxiAoKVMpkKnQ2rELsL2NlMXXnhUUqOvui1nxW8wehCkIxq58euA
ouJlyNoSnU46wLG6Gv7XKLugaWAGCSh/xqKKUbNZLB+3ME4jfH4yOVfBfel5
OmCqilnCedeMjxRrYP8KihexfNG4IAnbvKsFOimRVjbtGvveg9bEOgMfnYKV
6iv4vAsXMbBPSu6exztYmdbVrjJhR9IR58bpzOuK9LxXIu3nj4QgFci1N7mo
2KtBP3f1nkNd4B2ZlRLZhU8hPMfxly9jidRi1U1eXjgYQfg2BQ4sxaPIR7H5
mOPFIpedterWBhQz0vvQVsujbFNEVRZsyp9lMHJfhBVsfywqM9G59lzr6HJ/
6a5y0PgNXcJ69rnUx8M2pWVNU85WYdjC/G7VTsP8KlezfUmbvIw/JRvHCxzQ
Z20EFHJl7SdWDknIks9yFrOQf40YIui0VlNatqhN6Dp6Lk2ABhwox8IgL9WK
ZSLfjGxILoIQO54E8u7slilqPUc8rsZeFn15DN9rsqMbJNa5D837XV1Z76hw
3htV+TIZfAhRS70vzYI3aKY8gigdTpWji3Og+EdlZQ2gqfbm2k7uOhOxcKEI
TvH5gNjeK68kqAruMtMfc+RIJut/YG8C1MoPeeS5P3qI6lTYCCBpfWF0Ik9J
UdkrR1dO9HdXuICc8jGxrV8DnuaJAod3mNQaGM+5Es5KClrzExV94kv+CmTS
ftrJbxNgN2iEd1Gtvdxe93zYgAclrt2Pt2dGXq9TOLfotTOGwyf9jCv0MaWF
4nxUvkdYlE2t0FNeTI+vJc2tJ5k87UZZNiPBMbtF2NSp+LovlSLNe/bXmQ3J
d6/3eyi/qT8nohEv3BP2cOvn5Z/wG/t5k8nwruW9KfHFSvIj+d8xolGM1mfx
Je3w+hUUZbrcq3SRDQ2OvHLtVFYK03y+E645nqIh222ikKoyJpixnFXli93J
BpwmnviUSw0CL/hjTRlU5xRrOrrhconxIQsI2snkho44/pTu4Aypze/lfNFd
43a4NCSbPW/YG+E/FNdLfqDh6npOHC1AEvaltRrTC0EOW4NOHQaoRofzLAms
h4DQtD40Ts+er86XfxSfwSFeyH9tbG3D+rriCqo6uV3xUSt1dmvtEVjah+fb
ue4UPiBnhHyg6ZfpQnQoOZ0KlB2stCx9gx+YLnUlEEuxERl5I3tqrxOkuG2f
YD0PhoppX0vrEseYLDE6RchLQuycIowMvduU+h2o9KpMPyBo0ImEosUBhkRd
UtFhkuCY2Y2xNV2sxyTfCJXGzgEwUTm9ZKWpMo+ufYWHL3UgFLzOcPm7WL1k
ljxrTFHOYkY5+/zFC6FPTcH37FhrlEJPBw9ps5xs8fRHmLRWBC4xNJE+0rIA
8njx8SS7BA9mH9THctbPIePTei835wH4X+viPqtw22qQhkKowRly712F13fn
w6pnBE1Hh8grgf3RcT9gAkbKHD3/RzQ+4thWMnvCJ2O+ueJoFu4KukJYVwfy
rQlleF/zB3OZfGKC1td1YJ2W57GwQv94efBWvVutdTbNzOb4vSWknsMY9wQz
RRqWJqb9zNUyLJ+h7Eo2NE336mohG2kDiBa3Qkc++xksuw64sYVKFs99lJ9+
1OCk/dACN5sPQ5DOnM+kO1I0VHqv3V5ettEuw0VNI1JA7m95s9i7Wym17IiE
wd7FJBPozLiKscDOSoxGBtS33UQIbox7w3bn4xfGQnwuyGTamM607xj6FLNR
OZYvGzFCU1NX+d/gVldScM5QVIN8qpJK3iioiQtu/Hz+CpfzGheTBSMk79ew
PrioKsLh5+MQnij595bUycC6kG3OZtY+F7z+/BCgcbwtxyHrwZ1pPKVOwdDZ
dyEjNs4ak+4qRwAhwSaW5pNpLKq6qfp4aCfT7G6SbeC4qgPtbjvYX/iR5azM
DZckKkH/3QGDD7vuTXwTNfO7WwnX/9l9UN0bUbtlp63Lb/0TXBfHlmT+N0Fa
7WA8EBfFozFjOL50G7GYqbC0wGmH+CzhMWy89JPPFMI/oBcL2jc9qjcV4dGz
qav4ln695bK7SVM1hqNjjyFoajEioJpPTWmil8oR3/yomEqA+hWjo7tfCpgi
aYx6b6EBIgnksf9zjlfr+Tkm86F4sU0nXszsiIw59BSO2n4KBOAl1BEehkFL
El3dJkJ1TxrzY6dlMqPSNO9fTZXOW5qiobFgXre52GOsKiaBgJyIjRp4v1Ie
uVjBYJR33YZEDmXGEQ6wKEBMC8RmH77D+6K+QlQ/H/eU+0LACEsFuZ7Uj9SM
FX697Ken3YFr09tTg5b8szg5j5K2I/LuNR2r5TzHAogZi+PZmuFyuM4to3Df
Hmv+Rkm/XZTE8dBJ5jjvyXnfzhXK08kMOJzZlxCaodX+xiYPqt5Jj4ifSSnR
qTgzJsqgusaZ+J0hng0T/urFWiYdVw2R4/PRl53X9Hff+8hoRGBlQ1/aqJnH
TkX1zOkAZDLSc2fHZHfu20DUwZmVIS7lJLoyOsow2OIft02kaEjXcjfJ8vkX
+GdGi/PLf/FKpIJWcP+PJf/A/2yagQKxIq/7QcCVKmKMJT2adKCoJAqJjFXA
B9RgtYZXR3sJu+we8SG90Ck3xBoWIMgMQq/+di3YcjYOLKd9MB4/MKB1SOp2
J5oc65k9XaJkGivC2xjzCUmkC+zmzeDlUrPWsu12TXQMSz4XHlms+xyQz6PH
+0L/TCftk+lZSvZkLskCk2Uk25lzo4N16sU0MuIUmkCSB2hNjJMLdXuT7O0m
2jJmKj7rdcEZw0i9TYQtrYU8lGc6x5uo+z3vAI3kz8Lt/kA4ldRvTVczcaoA
e18AORzYeDVArioe5KG4M9BBDR3OQ2Pj9ZpgUgGZB7orBJ/yjFhTBLjy967M
+TZdDA2mEgCrUZz4aGHbkjIanrjw3pcEfSn5xGGSCagDS06ZmSI0U7pgzao3
sbMPijwYK1uAofAvq0lZTCqhpcunWxBlHF8Hqki6kVEQ5U6EisW1qBveYweK
pnrHKBh+fHOCWbw+xxyQSDOlY4Uk+EXJMz+liSH+8JpbVgLI8/C90Ny2CqOW
+17/SLjCKttfwegdD1MnfFF9aUP9OXwekRmxsQAIkWAP9YbjhLNgDj9p4/ny
bqVix8c2EYzf0agq/zJTQeezewtmfhvnMluDSDGupNr2yQcv8UAUFVBqhhKe
mmAXxpgs4I8FnF2S7rOcKT2QTkQtVtuFbb1sk1invtD0CupiO/ZY8da0BDWI
u60B4bE6PWr/Dzo4JLZr3ZHV/u5sLEMyGM7O5eJTiQ2mLL4+7zTIjbI+uugE
1JZ3SLX1mmeF+Av4uw4F/1haif0ZZE5o1rhFpEIrptEkJX6o+kEyf2R0VseP
wE2lNwmQuJQPiCttBw4G4El0Vx4LMaspRb7CqwTI0iFGvNQPJO9/QmI0g+QY
qGnybi6ZdmQnFmKZgItnVWaH1qiduBShdYv7/CrLWO559xc5jCTOJfMUhGAT
mTnBBnpdUmAKcyHgtTiQNAUKftEm25rWBpWkUhU6zGlazq0WzUpLHN06ecab
F0ynJHXLAwbrQwMatazjL6/gAFXXRRzSeZCPXq8VKbFVCEvKL0JdvVG71sS2
DapOVkLUK2HI61s62VIb5nC5ASe+5o97qh9GoNNETkAC009w/KYPGHmShc6q
eosWdt0wcEIdpYRX+uZ4cE8f5GoQ9UmVZHK4S2pXDQL9D39DB6PVMGEnk16v
w4uncyVCR/sAG7O552yIQNt9wZHV8g06Yzjs39alHWd91vXrN6WtaQHSs7Tf
n4e3KeG/gN9azwHHi134wVLlD6ROwb/IuyZ3HcbbqxlkEU4Qp+tkIaCuEvii
W6YOiwTpwifzdj3Hk3YckNCKJxwLT+cZoFNMekawrb2Ee9pxUdlBJrKIR1t7
sQWrSP8MRbxJLDEiy0zAU3l/mUh9G4fZy7+ntc7uif58plwqrG6Wood+g/45
2GWrWAkui0dWCZPzSMuPd6IJDkgjSFamzHlaZIEh1h/XXPlE9rmZqpINbhxH
91qsWN/HqJcwsWlR/2dr+1dwVHVc7ynmg/M905f4jMj1pM4zkkiXIfXmxsuQ
TVNxFlkcYSnNLVqrMtkw4Xyvv9m2qOxgUbl85U90acRbTfL8xTc+E8Mnjzre
lVFkxbBaHdp66aiTJ0ewkdQWUI4sORNbhyV50QD0OEkfvOY42mMMZhAShfua
EnnxIFWUb+4n5vOZlLGaa0h9EPvCXRjgmtu0Yaqle5s3R8Ngw4bBa7ZaJsvD
eR5AEjxc8SSqEsnfSSw0gEKH6nzTL+PxVnZF4jlawqm7lZJEzoZUXf7xH68l
PSRpSuLG51mKGQVr5oOKG85AY/MJB8Rxlj/hC1Cj7uP8hlI5lK0OSniwX3Sg
PUpKT+c7OGYLnvJcBWMHKN8mt6GxNwGrBN05mCw064esSeGkrj5kOW37cRLE
64g9EFYIm2J4VtYMaIn7Qd/vi36N5jKAkOaptc6Ujoxt3Q67cibLCKmmPRjY
OGEFHFsoWHX4oJClE3EJPMnj15jnpgSUcWRavhV54D8ph7y1txMq4e5LLgdE
FYupMAXKNl71yL4uqPeBymr6/xl29nynlWep9/VdvQaW9dtJ9kAMLJ0vLPIy
heq2BFT1UbyTakdJXm9RRbBiQTulos85envwJQopPbT7pf2O+jBK+Vfii9cc
OppAFc26INXcY2G/s+1hORpPpwAb3lCZ6p/SDyQ/zsZ1Ytop9LR8V1Em1Yhb
l1UMRj8hRO87ZunJkJ/HGa3Vg4g3n6oG+fGGK877eflYlbMzz+7xRC1c+mIK
U/AzvLUgs8AE+sbGODLNAXvPkS7oTmSZYEL0/RJfMADXVYllFACTUMqXIbl4
+0WJM5pP0mlT7t2Z3JZcDJSdzG+d7tr411K2OT05NXUGWU1krGQ4ZKx4RjrB
3sI+/+Xjf7zXzgdUF5s7t31MOxvXK3oBxMBj5COT/u3Sx2y4Nh9JS9wdLc9y
b7omR/rddGb7/fxhaQBVW9gY3a3OWDK7tfsTI8YxHmecEGc/tyCDeQyhH+Kx
aF57SFzhnT7Dw+s0woE5TahHo9KLhHz0e0SI6MqD6zWFL2rovRbSzjbECxJ9
JIOIOjmYZcMK8om38dCA8LzaQWVVAs/Sd7jfhLrKQ7fmeZjl/6qzOSvXMwJ+
BphsNfcjukm2hGPO22u7OUZIK4J7v1JnL2TKRSZeb+oTOgCMsmwDwpbIe5lm
rxs8YIixVj6jAY40G0/LNZ+dX3vh4bkvwMicW7l35+jpd4MH1DYyhW05hO9t
jtG6qArCwjzadIR5GpbUMilMkX7RnJgEo495pHoIj0W/bZYSBiMqRrqGXECN
vjJe++0BdslXTB/14DoGya81y0JFGp8Ai6qgqP9mevZ2yIWxG0Ddm0ZG9bzn
KltvTSWIUy2RAxjgP4VHT53RXSNvrbPyxrRqE4IKCgcMj6hKpP9wLVhCIH/D
dXLIv+8MNJZakjl3FcBdveRObCu8ynVaK+cr9npmaXwrMNOYiLZbTZSTXPtK
qONXsoHOTLpKekWxDrX4MrvLqU6sCbAQIPodGRPMVPNdf/UeephC4xv90/ug
M84bbIOSh0LJYXDUe4lQ/ot9e39weHwl+jNYuZzUDxvw9PLiT1neiq5hQl8q
eVK1uzYcvqSJzVLtoX0mv6wfmkBlBps4o3IsV+0w4ze1A0/CDsoFr0DG46lC
SEDY3TPp35LdT7bc1XCoAjWPbLiSrmXnrxaqqYwzSqvOb94VFvZ/4JicK94m
VJV3F2P5NuEF15D1boece0OtxeMLzkTajBeWu6Coy1r6RFQrFsuLFOfWfBtA
KAOUVxRMuX8UGCsL7LBsPaHnpANIjmY5uKrA4gTOR3rcBcPurRmFjWhpWwPa
y9VFjGCz48WULo/PPtCQtgYRvxSHI4HPCn+joHWNy7YVxxOB+egyg+mMbTq3
KZV56D0+3gctEaMuwmr+PvyO5PHXJMIpBpFqvg8Ho7ro1lTws12BR6CFXcsT
e5klb4twpnh1sJGIgJHpZvENTQB/ob7Z8uy+YmpC9kIRpLeTuqyNCbAhLkew
1wKvSLUHmvHfZU8TBHXq+o6SgTuqnXRwp5bHayjO7Vz93z/6vCP66RIwcC05
wQntwyOA5hIbjGt/ViFy3WhydKCtq56A6UPos9yNniRgBo4JE5is/+fkajNk
ErJyMshbB8V/BX5cyyuKKWGeh1p0bAKeLrIt5J9D5miDSJZFpmHKAMahmVLL
KN+wv6ehfwSTzzGUqwwWwFE3ibE22b80JIVROWbMLscR8thtElvWEwdhh1AA
V02kjo5EhGfgX4Ukv4+CIxoB3N/ySqjzAhPQRb8RqodJpNYHY+b/lrMOF0cW
u/b3DQuhl2AyyYGeOQDX84gZiV30KpCsbpmyx5SZM6TD7pjJqqqHmDihBJTS
8KIkBTTKYzZOjWmX8ETsAYnCO3Thx1ifZR0mLkxoXYAP6VLZzypCQekHSgNW
1E//ADo148b2fcqGmOu2tzEW8GZloW0QFvzUWrGIahvXzi1rEQ4p7WYcfE57
qaeU6/RsdQum3Be0N6T6IThhW/RLk/bVw7nZ1qqPhPs/CfF7N03g+A4JMVFw
eOpXE/0456j//BLI2ZngCi0H67j3XrJqHXsrxHa7TTK+6Au+3Ll37pjiDFrs
djbJ1MHdIF25Qh5NA7R+8qlUfOQ/Pt4Kcq3oZ04UkiCqwjWokev5x+GnAZFJ
WwylJIFRB7vXGZjbAumOCIu7d4QlsWqabMnjzWRctPke+Fn1JGMwxOkGAwoV
e17vAk8BYDIoYDfolUWTt5+m/ON7DZ285dIcQEwN0gRIxc44F0evSuRidl3Y
3PLz1vY8fh00e1+kTegt+27ZE7u5VQ7mZWjBI32ZeuT8ujbWWGg8Y3LmZMa5
mQd0LgGJZdFz5VmyX7P7bg6l3G97x2NzHGTz3dvEG81IKdBWico+WKUP5maG
grlg2HZnGLZ8nsgD+0nF4XN7pSMm9b77yQXK2wDDqXbaAew6ToG3QbWpbkOM
iixe0IL9N9iNIlUTmrdFBT6xgtiA6CnPPP8spjEO9UpLgo8/Ngg693oCfvOS
k6QDuCVmDtVzz+CB5La7GrGU/UB5D+u9YzntO6gLvsnt0CAmYzi7imouvaln
lYxqhLcThUBP4Ppbq9wpS0N5jb4hkNxy/bR/IA0hSVyyUWOQ7D7pD0GLqLOY
rTfj8r/Ad5wNg7BGPFt5bTUMsinLhUZNzfwqs40FTP2WxdLFL07eQw0bYx1+
gWRyAGiGDp/irJ3bMsfbjYnSXv3sA2UvGTCU+Udui7aD/jcAJ+PzAeerq96j
PSmQq32QE2tQlu9/HcspPHW6fsa6EiJ7ZwRhRqwD5UZTevuAF4u2tWP+GZQf
qvLAIKkJ6E2j2xmshlcxQ6mQkvLcwV9jBPGhSTiZUKEFi4yqCadPrXZuXp/K
fbhWjpJScNeE5ly0z36uhsGqtJ5quaNTKFcqXzRuj3+DLl/vHqIKVk3dWnwF
K2OCqoygv4t9N3/KzClEitW3BDOzQH6+3NnUHqlakFgBOdlKNoiTmcZigf8/
LJGRguNBPXgEcTTympkkCYRE8TUHpgioeRhNE3Mp/I3rjo76zvSI5q3F0sz0
YCPnlTbHPoUm2laSBiX2ZbsqTnGdGZchDyYDO49RF/w1pNYOdKf4eRAzRycl
ri7PRVWAR8beJ+uRLPq1RgAcEIgHnA/2EIwzRqkaN5p+3xSr3BTI/qZ0nXEy
wuvCGmegxVDWrCEW6VgEA26vC3wZK6q2YZyfD5B4q5Fdz2khmLzkmTIgN0Cg
v4NEMJQeiGCyFqIzFExund6jnp0JNuVzDWDAimbaJQEPgxp/zkkiCr8F+D+n
85ivzRynACwnrEVqro6UtjvEWyqhGvYq1bfW6nefO1d0Q9qujTN5sP+0M0v/
OtBymLxDASPnigqMmp/55U8OC0DawGGKnuPDBb+j86+LVQ96/FAlPIm599ZF
OA6vK/gO9ggdhzzw/hARzY+khcrvdVmCiHTEQg46d8T0bqKpcTkuMEqvV6Tk
mvMTSuJzsGoXAvR87yt0q6yOxoYhFinlxlPh0JknWHFAVWaIBu54aUi9o98k
RtFB9D9Pq+csEC3YO6aA5184E5vpXrqs94kt1pODwhq/eXW77PH/NWn05vTm
kJCA6+/pbbHe3nB7UEGc1nV/5ayFBsGJcX9SlrdIpfOFaS7QZ4jwB691nD+E
Iyvq6kpPj9kPXEQL7M4E6J5nSiAULUehu8v6r8A9cWmN6aA0YHiAuoGaqLLx
9QD5pS8+A84Y5OfJ2AeUJN+J/IxnYOvSwxpO8WxYD/HBoo3E4Wyqd73Q1EG/
xXMg+eKBRnXTurO/vLjR5vCzKqHIwSluZf8tiCjyUK3rUi2NQRh3qdgaespE
X6FfEKeUMssPq2CTWWS2NDbdK6gE8HmZcz8dlXO2OihXbLu+pq/k8L6L3/76
lyEPkXyBdAV0hJOIVIu63eumOjSOafjl0BE3PhlByYqwaNecLKnuFrjn6zaZ
EtrI5wylruq1rzyTztM1PK/LwEMf9sSSk65zSRA7vPT0TTk5lVRUG2UA4OI+
beHrWfeDgNFIIpvFSsHiVtE91kUBnvh2UeLGKU1eFtJNk9kQPzDGh4DLjyV1
ddDYdeATNxGV6mqZWzlyYNE7j05YFbshJu4G9BDNLgygxa5qg5K4lBxW1C6o
0Nh+56iNv93Z50lrfNDzPDuntldvpbTn3KvQa3DcVgjJZdYP1d9dmXYBbAnm
QEydOn2jB4VFHKP8QcvPwkYcRl1rV+bdo8wZBEmCi9z5B3deHO0GazEzXB3j
xy3vyXgjqq50HGlUKaTEZLsJcQXnx5czzxi378fZyaQVHyNoKpwPNPkW5nVK
lA/XmkmkstS1ZAzkXVMlNB8yIhpmBvJPk3NaD6BFru1zSY0GX7kD1bzx5lnx
3F8qVkbSTmsTbH0tYIC2m15A0YWAQhjNxG8v2mLrrRanGWf4IusAqmIXggZw
7lSRtfLu866EFKPv/lj8vg2phIciVukCiTULGxuzPmqKJU1qjXFEYpfFd195
YAF4TAaiaj4AQYJdLGgIqNIhA3CaermVLypIoePd69VnxacyO0FbZFeAUBQs
v7laYwTla+DzRuQMVtx3iCUZUzjkxb5EWIiolG9bnuE44hmhTE33A/oA9yj7
bdYYqR+Gecz5fVGk7R5LxSo8XkCFV60rexU/mflN3Nb+XCurH1ilJRNlfTi5
w131JuO2n/wUaA5Al+qGgub5sbda0EniXag1/6CrFLOM3NsxZPQF666hgLPb
7bKrHUzuBRDgB6cZV6aLF3Obkbm8jIUSFdsr9RUSIYM6RDNnkJu9bJAuYpE8
54tP7tv/drYbYD91Ivh/YBXCaT6mNn/vidVIn6HahdQk6+KA2+Gk9IOubG6v
k9KCiD3EHojJ8TLO4wTTYN1h8wlD/qjE+PLWoOx59cqdVr0qFtUGEry4BslJ
iSm5Dz1dy7I4nDdiCSSxw8aKswzU4Ifq+p091iTD16xSZS+KUvxc0YKXxD4I
/6voVJ/y7tVLktqr2Qq5MwVhqGLqWT1qfFTTDsLPaH+9a18ujXIUOGqwW9pP
7NCkvtN/TNKpeMep/VemFjLHWzg29oaXLCZXOjyWj2IvSBV9MKL4CCU0H32I
aKnGaaNwm2csBylgKu3SzXtachflgoSGcSLvbtJIJydwsCAeWafDNUo3ncKN
ZGKHkw9N27pQ1tNqt5ZnaviSdPFnfA0OzXKmh8lZp79oDdZPkfKX9jNKEcic
l6oxfA3qn5682SeQfeD65mvR7zDlkE8UGKQRpLBdFRZPG8UbLCpXxr6bUbdj
JQ31W+PTLMt27BphDG+Ju2zG652zreZ4vIdaZm/o6UACNlSMNrYe9Tl73EKF
mpTWjAOp1nxXin0tWkcdpc8S9G1VAamAVw7A1L6A/iqi3BLm/aaoxHp5e2bR
+WuDbR0FE0nMFbaV3MZiMZr5+Wl1JiZSnJAcA5kL38z5yhR0V8qk1MVdDC3D
j2/c+EALt9D846KX8CFHihZnzGAnlRln/pzEEoGwCVxgJCopslGfJP6XSHRd
nXPjuQmzAXhH3gw7dnLyvMRhPZ2jAv9xeAnE/L7PZMWBOXT1QB/lYISai2rt
rssC4e5ms0lmkr6qROTx+ZLn7lAqEDYkZwxviXG/Lz8WgfVR0iOXaFuf9BLW
9Q0qPzyy3/GL9BF7Ve6Ek2mwH86PTFdZJ/k7zsmeTK1QFci5vijvoAtfqZDV
4uZP944xXMQRljkU7HB0RjNr5jgOirqLLWt3Glt+qXDfpcVXLGvZrBdompU1
wZ0FdHEboIeLo1q0Dh0EQ8yjlbrRLX9CunFONwJ0Fy1g4Nb9SlJCJv4E5NhT
LHfLxUzQkZ7mArMT8lZbQKoJoz8cbeCyPpYO4d8ekM6VI+IrSIOIF+/sqGt2
m44ZP/1EXhxtt7j0lkb7dSeh/je47fFRkkezsBtXASpVckN1T6NbfYwjjFbI
AJj7MMbqQZwVlTE9R+uojRtTm0+1jvR0AlPGmmR/WlWncJNY1vrmlJdgy4lh
NvHNVNHh0dTLY2gvTBZWcOyPSSIo0QBsLLVv53FpUndzYQ5aZoMrAm5Sr2jM
PCK2pa4rMb6O0tOWB/iZn/mUe8V9MqU80HZTsKd8RS+N3P0vi6IdqkGBYTlB
UCKTVkY0K8k8NPjqOFuNVR4fCP8DlbDX2GOkgFDLH/5RJb26OXKe8FclhVWn
of+kK+290u9wB5+Q4HSIDJeNhMmYRvwIj25O3J41NVb/cmGRO0Y/LJcXrBHs
pGYK4gFvJVy/3dVvk7Kp0h1bzgVySRYRaWfMPpNYsWzm+rkIVLxpSE5NL0ef
4R1SP9I3AiwBboJF0/RBa30yphWrmVT/z/uhmuQkuVIDFw/PXG4/JkJ89zXp
RaMUM0cZ+tvU37mzQJxUuX3YXbF1sbcCuTpzesSE8L/enixe6II/UIl1iyWO
mt+rJPFT/Rw6wN4l15Is07v29kX+i3IYjay3hEgV1bE1TkDBshHiQEAOrTOn
ZzZNYcQW7GOCzeb+SQAqV2ACuTBuaB5TsfR5lYMm1H3qqvIClz3+jgGpJVWu
i+mSK+E8UHOSPaweAW8h/2ZEHA69rDrdYAvTse0bx4o3KZZyBEjDbW0h0pXb
NNqhI8PMzM7ZYWATiEAbgt44vm9SAbRVP/3jmZ4WxHn6mwLCCLBZE9Dy8Ch5
R51ISyJSp8AKXZOrFaGBvPegyrkFpinsGQo/nPzHOG9WTvgXDjpt3jLf+L8a
lgyTMwm7u+oIUeXLjLxDIoz7GtgDIdSGV+frcBNEU+d6AnpTtCF3IeIT7hIp
yunDmqKqnk7Josy94n/QlTdVatYz8+T0Zv1cwglQyktEXH+M4mKr0Dmli1T8
QK3cmnc0exBbLQRjBP/5WgspHzOTw6OjHy2/w5LwBmtL4cc4h90ikta6B5HC
unQ+epV5fyi/RgQ7V0/4T1Nj8XnwNKl7mbSF6xlLn/AICATFYYI/YxRzwhmW
PlTon6JXLNsd7UgxllTC3OI8Uuk0niz25BYoweG2/hfCA9Y2w7pjUTquQ4LD
huUWh9ufgUXy2pqgrM0QT91TUpOzwoVNDA/tkb+70cWh0XZO9U+1e60UweR6
iZPGyfHaoRvU0ICeut8q/v8EOg/i9QDlHHnsfbdaN4YHnStDw3y5N09pWt3F
829ly8KQXyWTD3z/t85jorWmhLrQKg4Sy0qCgRtOCFWeZRVmF0ThVpNWViVx
i0+0zATNgDq1IR6v5mmiUWZ3RvmgUPHDB/ti4SvIDnHFmpT4UwohClZXBrqt
qEuFO/u2Bq5lP6kPKx1IeJHV8xxA2Qyl9pk6XbPaOk575TIklTcCQZBIW0oV
aKcSTpTkZGscKufR24cTP2z+vFjvi3rbR0xhKk1fyGxyroLYoP3yDhwv8KRl
DDRiViv0SWV50510YPVqpwuuc/bHFDsOyzdPSF1lty3FlEC+GUdUOY5k+Mm4
XYTcf/4ERnWUc+AaSOpIj4XXHXDK0BN1SJHzGgkzllwuSDRjQlhZX9Xw2/g6
2acOxsY19T5tkRxf1IWZ+YO0ZUy0QEFROC5PY1t0HsUUxQZCijYNA0mZoDPX
A7puO3J/QH/EbRvyH564bHqziwqFHsqELvCjaNfu/wzCwZULmDtZKRMirRPv
rxihiHe/NoO2AsvzSlsHSohZfDGRavNTnosMfCgaVcv2UwDEsGwXj6AlksJe
hFf883yNi2nHq5VHzq9Ju2wLgzy+LAfytvET07YiSLV9Pq0S3dHwS2ZtVkpT
wev+ziroDedGd1Ew5WoZ1N3IJoyxwJg1ubsoifmu7SsA6oDLMcDDNER8is3N
Z0Pd9CY8pGtgSje9AGmlFA+ebWMJEJMbbVdRLPTkD41stK04aw+EgmqGqpSz
mPzpNpejDy+ILIF0WPOCwVj0qCXm/JkUYzMcIfMnXJ+A4UDptjn+O9++A/3r
RZDm6gt/uqvxNDR1yPYFJkU9qXbzbPKB5Fy3WI7N3Vd9QqxxnuD+XcU1msrs
dWTSxm+eDgwtiJbieI2DL2O6ThWlFSTllGsxwrYUfvIbJm883cUG+LIFU7SX
ctqSIsSpsslBpTNhPxU61rSNrE5EZS8vRveE1pkbfU5Wh0J2JoIM/zHRaJ8e
sDnFUKRIjPCHS3j/tQzJOBvqR36DFRTW19jN7a1ReYoaeXw82AehbsaSXuxB
NOR9PbbmgYWKY957ZbO4oW8CaXoIGcSZ5TstKIXDSMpDV6KTQvDaC5D6H41P
ZV40osjhSFpkpKhcX4XNIaxP/N/YP5iCR/gxDp5Zff/Dq3i72hxDrIq56cvh
IqzEGOBIdkS2frdzpja7hcTbX8rSRUkwVnLFKKWUDCHf5t6Jf0TCbV9bFiXj
bJCs83gWHaEQhePfr/WFOltL5wv3gynpFEJ0/lSvx/FaVvBbmiA+jCvu6xre
u/89cqZPleQ61Rx+sBm8ZJVUYe6KIcFL1qtL167CLFZOu+zZYUBbQyoDcC4P
jWnzY/jEgh3rBn8i5UpWOlZ9anvleDERgmNom6oSwukHOOrcU+jDsIfbw9Le
7QlT+6jFScjFK/Jhs6LtoUra+R/TgpInezrkV6bTTiLizKXp44lgBPMboNl9
JkWRtsgMdKca5hXRpiUru4xl4SNU+3zp3szCYBA1vtikAr/WsS/VGFD3wPf/
aK/BYdtrV1rwwPhkWzw/Fz3uHzSV4u2KromM1oOzcRZG2zhNzmAmXzoYxZZU
8KZKEKU9SpC8JskX7d/o8kHX8J06WwS7cwrIxg1/QLRtG4ye8pmRUQL+QxfX
tZcSdiqYxJV+lfhXLBKoh4RJEXhNDsbTV9kskAZ32Nw6Rikza0RF0UF3WnyT
wo3PZ8tHMqm6qj+FmsDfwT52HvHj+GdlQ+BX4XrjazPkeR48A9lAmYrir7XE
WV2vnM0487cuerc66Y7im1bGa9Wil0wP3T3BIzQuyDFVvxnt4IvNrLvFt0z8
jmIVZN/dAkq/VKS6+NFP+DX9xIQdXsSrc9j/Q/L6ZFDyiNxQRngUQwu8U1v0
ifJY4cZpBDW09SDTsv2ewyBcc3MamgPtOymz8MjOjXPYfYUma3uFmvD5PfIl
RWBfF1EsdLJYqfyFz3CuWmmPM93Q03V4MsK6xj/giaBvZDOo6OIvllUepuj0
ojcSWwJwk3PQlyqaoAbtQ3aA2SsCkOA7Da0JcLCBY783rSGFxUdk+ZEIHLDA
seJltsjlTsVEd9ZCT0vXMJ/I5oo4xY8i+ZLiC8mD5v9wIlCI6+T7ZRovyztQ
DhBJ02ctZmfKAdgcKO5txUTARauz8hxzCsW8bbD8QP1tN4IfFwiSQEICr0A3
VaLRyQhnft5Rgm6+DL8pbfVbvnjmkAlqMRvhObqSCW7Yv2Y/t5J5XVKGGCDY
VIAEw6EYtGQvy4/FnMED40bjbbKo1SFOPoCbq2DG0wTIYD0/cHZDq0YfU2BM
aF34HBFWk0by2r4vFMYXIcYbcMDzGUBfMUTDKvIhFkYLIVhcXGrqk8WZzeci
TGyGCpoIj7IWm39FQnlU+Y7k8VSRs/kVTocCxKgyVAVvlTx6J4hlPjUonOGb
JFCFkiheaYnTc56B2WNMRenVZkh4VomQcwWj8OvMyMxO6aggc/Ib0TAaEshp
HaxO3EzjCXWYSmF5yA1Dp5AkT+q9dpOkfy51xyQ3TVcAFL4z5mfLtB/vCVgw
XYghrpc=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AHFS8uhOzEEv0qANUjCa5shxFe8bemKFNhQTqRGtC4pjovR6jkEwCgEM+HVx2+RETJ81jdGctIsI8rtsCu4TOBbfINYgMfPtAhYoq0pIwXzpBYW/Jwh89yYqmQ/8qwf+UZ/RCUPZ9uTW2DZjLM/8DQwcPSaWPn4uluTziVOYaXqZBjqnFFKudtGOgi9fUYcdgmgi1Cr8qg3AFyDXZaw0JPfMHv+sI1tXM9FJgZxRxGOGBKmldWS+iPjtq0SAvoUjx3YsxV1aCqNZygxNfguFZVImXZtRmvgNFevSZOOraV04qAQYaIWTb+ZWVDyiucFUpfW+4Zr3/B5rS3rO31ArSXh+i4B/NK0PrpXuFt5QqtB5UqK0eFR9eKEPx4VB/UyPqcSdyVmeRj7504fz+0nruMacbprE66E8RJfiMhMpUsa6220Ur1Izc0Oxu1unGLUSl9vq2GHZNWEnGl65rw4Y6yhyNLNzNbdid2LkGIg17Dps9H2JNOWeGzukx+Vcptk5CnFg/nxvvPUQLzz1bimvMNDpM+X6SCbOWam3dGSv2aRCAZyWDoJJdi9NdKP1kbKD5JAZ9OCpRSdLOfB1tK5E1v26cH41N7HIjKauZE3ugvCOfcjU0XlLhJdUzksbYRFlNc2arzGiEh4ldBmFhX7s7/cgdGoT6LrCS5VVovTgP0J48AgK3QtLp+AKNz1zzwaxbZ6uCLpHeEQBOwCgKYoZfGj2hAOvakI6CeQNofbX3hQ+f08zZ2pJnGOtR8Z/eXdakP8QQg90j9oK7m9ZpXf0ciWRU9g7UjJBj++KdUZxW56DqcrDwwelXxRpbFjZLd5JSQD72MOlqbnbEoEcUbnikPYdOfeM8Yq7M7D77674GETPVCU1aAfpN18jiTsjctJqkWqg49l6HxxzHV60vWeZcJQLUzd7vmCOK/aet+208rlJUrTRFCel1ZK7vYbBur3xjdi8dou8CbqnpIflL2nZL6ZKsgBsiAGbVq88x1R9Vvm3Z4WlPSWxDmGH3WpNB5PA"
`endif