// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Pwpmqc7x0fbeBkTch54R4eEHZPjnsQi26dGrPzP+2Ia/Gk3ixzD4rq1Gxoo2
h0VGMw3dYYNM8547dOnEjfmmCEkJN6ljYkXCo0sYVaSt1WJnEF/bCyAh/htI
fVnnW0BLIip58Z5wEaSeOgT3HXxEihWTR3lSltrd8gIID4ZMDKINCZMk99Ws
CId69T0S46iQxiK2XgsWmBAwOWIXet+B7hHZn8EoygSHv+5eR8ns13qJUk1o
jz9S7kmmlMdOokbTPWKkudhrh72luOBdbCroSgB2LFjf+ZLu5LhHRpUf6W0H
FxVf/czz1nUKiJi4bXGkUukKN0hZUNzNOyJ63+Jxkw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KwxkFW8RBr9i7D6weU67s2Zf+qoRu/YIZmu+pWFSVWD/ozRDipWsaAvlwNMC
NzDtOvYSIwL4nnTzaRSIvw3YbrSdzK/meckxY3UzQXC6YtH7RoXhJWcIcmWp
/vWj5TQJLFWGHSiUay8Lwfp/unOvVkuN77PjfOo+ekuFMlh8HzpXAdbgf/te
we4xurT63fvMuFVMTFkNuwwYfFiz1E1EoKZj2omcuu2JlqmCiJ1UiaSuHcC6
DsUjIrVpkTEVw1zrwxwI2SPRwd9F9DsrLKCPQhpZEC9B1mumSWb1JYgUxfsJ
crVS7Ey1+KAS2RRR1qqdpRRnx9HAB2lxUpGTJ328WQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CwPKVd45a8XERpApb1YHd1H67ARalTNOn4UgbzO0k0gWL93mFPyVx/rVGoBC
V6uq1OoUe9AB1miaraTR6zatNRfIGDqEMnlwoUnDKRSwhemqCQWVFc6sdyJ9
L2zXIHSddSsUxFEfk7FinvwUlu+HLGXFYvQPAejZRszgzNv2PtrFLLXlk/gs
t9hbq1jX7xn0iE4XLgMcdcKVH0SdqRm3UhZ624AqnOK9i9NxPdjaNSpCsovg
WtOBpsPFNmlEPhrygk37tTHl3+DotKuCzyd9aaG8Czu3csAS8XnlxEnHdtrA
VhoLhGGJjzSajzl4Y043tjXzcjq1HAwx3FWXvbd4ow==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BNwe2BMzvXuwL+h5BTei08Csdk9VaoO98s7ZDHp7+gJ+w5ievWox8r9gdDbw
gsfFwKMfpnUh4/9/jJsN0gVyqEf2YmYrUQsMnySqa2E1t9GOtS9tBrRlJE0G
ONqZrxJH1MNGZJgtOEuVQZ8wG5g64afFeex7DF4HgXpGcHO6eo/qeIJT9pdZ
uI/3aVaBhRnVv8K91t+FVKQRdZ2+cjWGBEEf9DbNtD/nZI6/YI1dJEJuS93U
4uCJZbXn3io6AYw5xiNEkCH5ZCxiJ+y2YDhHNIaoUSFdXSe+mU0rQbPoM36l
oaKC3m7nIYqWfREtpeD/v8N+H2nTxtCk1OX3G7kXsA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YITqaCM7pISmAqzAqyhM2Y2Gl3uObt2VbAZSAnv/h2HP8t5SnjJn4Nac9mVy
wAaGqvm7Jd3QzE1hBVuHcEobi7nM+Hxjwu4EpofKBNdMn1c+1p7eUt0TKRCr
ufL2CheEm6R3yxqi1Y9HlB7JrQRb76z20v4ONS1R9C0OtDqKDmA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
mNhwLX+GBAIkba15hRiUNn/l/dmXYVOvAo8heZELJYzzUStdeaZrvas28zO7
iNrIpq+uIrW4sB85KTIsq7KZP7Bxl2/s3lY2WoaU+tbPQiOsihv8ugJZzl+L
ITb90pXRNMaN1uoGTk7nDqsnoGQCqa46ZDkLh95aemRxc4ZW9WiyDWN4CFkj
IwiQKHP+n+2hslcpABtJmvVU9j3n9wz4spMXqtEodlu/6HLSKfZsa9Y1IeKr
1/qTrwjR7LN6ynXlm5bNH1+Fg7ilsx0d+Q8cP8+ZP9AUSYQyCZ4lG9joE/ey
Brin7/bCXLWVArUMeegUuU4pe6yp1YZUm1H3i9VdQXlSMVOwtbkQzQULyE2o
pasOa11SjbvVdFNxE99KMKQN+p3NToo7Fbp4+QwV0/CGzHxmQPdobl7nJ1f6
sZju+fCxksjWGCzU7JXjJ3tApBxgIYdNQGOB4ZzCLKfj0cqf9kHCQlfrt5TS
OY+dBVbNSZmTAUvNOv8fgYuyX2bUZIrC


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
euIe1vLFD2utW8e+RmCq+HOv1cP0OxZSwWVG3+6oyUCNeWyt4JxWE9Ipw6LC
ILLtHxyKh9Elku173HEqeHU7QXyhSBBtlgLnwb6SgrZveBRPDLlWWaj5BmjP
7j5QT/FcHgDdeAlsuZDG/za0CEYaUmMLVZ5P5zc/54BBxctX+Zg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FRhDnqIo20OMy3H8SqvSz31ViEIV7Y/8Q5fRWc/n0w8VO3kCo9vdJtvvEBsB
8Uzs+qCVD1Ta10W70XrSq9RIY0WZif5smXEGyNIjM+58FkORb+dJI6sFiXwi
ENkn9g2oloGfkPSFCwZS387tyumNadb5AQA59jdrz3URzpbEin8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 31408)
`pragma protect data_block
nGidHqyZ1t8VFt1KnubXbrbR1z9wBCDPE9DYRzr1TRbERDRXuMfipxbO+KqW
ogG+JKohrZBQqIl5DVTREiBMMBSB5UM4O27wE2gLkQuoWJR3cS6owEU5r2oc
iHGpGK0eT5h5997snTem3oGzypNhc2guZXklXHOoBEhjlPE1pj7MfFqBhToD
fFtdkg51JrH4AuIpqj6TPByrf2yMeJr7eC6/5uxbjZdjxeJZVN9mFVwYaVEO
/fdIH32VTD8tZp2vx0h7DSrzB54hpLKAuoWImzgzOoEXDV3z1Q1ul8UDGAXP
R/BfrWEL0a2Xjin4FOExdt2HAIiATDLp8cNKL3O0NAZzRCIA0xeQz3ENQDn9
TjXQXneoOhw7QXzh2M9LEn69VGuiwp5Pa7hJ21wmrmCpkFgDyVcWj5UV4COB
3mAvrx8NQ1WHS+PUhXTo99OTVb6NdLEuRBKeL73pxdlIPSWWW5a93CO6vsyY
IM4UdJLGPp8ZutORXB1pU1x8MqzgCB2IvEivwZXEli6Md20MTJyWQAdgMnN6
T7Vbea1hZq65QVvbM6rqYujFBb24vTjAYFQyJJOYxiNtaHp3ezn9UjVHguCr
Nt315cYFFQ4BA7jXyo9Q7OW/U0JG+8j8d43xp6r98wOcrEMvGeBfSEOToshI
OejbFJ5a1/Tnky6yoy95kGr/om5zBHIYOYaHlwEWkSKNgzFWl5Ixu3NKe4g+
vrm6XEMv++3rGZXqmfTCXMNYhwlWVSgQDxzCnsANCtmtJez6ZBx5uh+9fDNg
ImOcLnnlfLuUBcT7owSrpi6Q/X+kEV6kOT7kEa4qAcsgDCnHIzxXE1lkB0IL
tr/cRoippVWAorfCGXj6Lhi6aakbc5wTD/DNIVyBSqKAI0FpAIKiOmaR8VIg
CD5HIvpwtVGZPirAMqqjIx1S1s98dqsRH/LcqpOxR5di2Cx+HdcGty5X9+DP
odYU0kpxc8zI8FpKC6B7cEDxxlUELdBsseRrx+ur/PuYC0pEyVOO8UOr8MPD
79G/vpqTw/3DoTkIQLX/srJLvpfDTIHXP0jfBeFiQs17lnmAzD0tExZMQSrN
A9QF/RLJp8gdzRLz+RpD1BMlMlqYZb5TCROCnt2/2NccrtxZbTjTXfmzGJNY
kTLV0mLDJ6jNSxW1XVrCiO/37TYqdRPfkb7B+1WsU2nmdM+rw5+8bMCDlSXB
w88Fltd9tEZJGGN+2RcQxOlSN06BWd9/PSTuOrz8MgEGPdUAcaJRrKKu83qn
tghjlxOjwntLQYu71lVMk7K0nKf9EVbyiAjX99vsmqnhydAu23rcsfNHGvpf
OV3HV6kQrZ1Pp3tIrk3sFmFJA/D2rVhuF80HmyxdTAJ9Mufrh7qOqMgUTUJv
6xJTwHNG/iiJPhM49zEqVHctqqh7XIRxKYR2QOnlx76681LybRukOboH2RXt
4kis7Hhl8/O31RmzA/7qYrmO04Ov0aXwMcelx97gq4sFygfdRBKfqyV3QvAY
iTf4qvMLeQWg9WQk34l2EPeLa7irwfY9OPX/znwEE85qHJ8h5wDe/NQR4VUs
0NNVLMRn5WqB5z90EAc4G5mOrYv3iD/rKfmS7R2Aw2bod0aO6Q8/ht2RzSqS
jRbEzqbA5DUUUlpGiLp+DFmlCL4rN1StkKGPZ1Ui7M1vZSd/worfPo/EDwmS
7gjkRwx4NKiC6B0UEhhHxbXj1uq0hJVkyiuK9KiCEbT97jnXAVBQTkLQEWdC
n0+hjey+kdJJGph/+fUbNiRNyTJ4SrOqxv+ofIx8LA822UM8OMaLpvAJNR00
Zbzh1f8vUO6NsT8Gb5nKdzPm1obnFK1IzcaUz4Q87Q1wTozqVSRqTJE2RvGf
OtsvtIuzkEKQw9RHEU6v+5Em/Q9lHCfh4/drfGq2xMb4/Fz298bUB7FMK73f
uzGlHPksCY+s87odHBgT6Y/hOPlyWQvwBDW8FFFfFVkrCFVRxtgbwcfWIdqS
6NNLvq+he5VJ6ZHrnpvxsSSxaH9Vy3s3tw4mjcG0DuND6+v8wkYTdUy3XxoS
hNY+MxlZaJyaTGHJpiCFIaQCb4eiBU7Ct2h3lGIQJlWW7Q6DZFVeOIFzg0Fo
JAUhWTfhyhk30Hy3S7cnA7tG4vR76zMeJxjBGueYoDks1iFV0DAiDIAhURF0
4ihPogfHLkT1h1HwiiXbwuWiw0J8Ar5B/qPlo/6hxWEMH/NUsmN/0riWPrD8
YBRibr6gArGivhCeI2EJF9cifyi93ZeUFqB5RtK5xfB1exb9sm196YO94F0d
hVFWU7C0JFty6y5NK6qn4wBumM2LLBGjx1/g6YJ+J4ed9UQ1G45W1bylzG5i
fYEc5/0qOVac44eClQwdmKepjy1OrVemiZapPRaFnqBHMN+S2brI8WWtutzb
fu7Wu2nwfRPK6QisrCBbfI+EB2yHtWy2Upm+WJx2IQ+l4/XafdQ+QQPrdisp
I8YL2LbJ4UCnX9+MdnWD15RU/8lUuO9bpRhgfyh0/ZmO0GkDVwdnBVOT+FC3
nPZXQvCxgbpx08dDXmiTiFzrCqYavhVkCdrl4PEzA/yB8Bfnew/Mn9U7KaI7
ntr2cpAjdxDpNfkuTlwj+06H7ElQ3HH1fzlq+86O5XV9jxv3HPCgQd1fBVYj
yX0SQzlcRid7Flur35iNOlikTwtqUfJKgAVw89j8yEo5mPSWh2qhVJvBlWSa
n06FAjq6l8GlN8WjOONSMSwzwy52yRtscfui4jiMOYrxIR6RbAsD+OH3DvDm
Fn2wYMdFr+SLUto2rPPC/w9kD/+cYAVbPDrmTYVZ4qEQxrIx4j03tMOD+daP
MttJRgh5qz2+xFhC5QE6SqhIhtnUgWCPVFwDM6QzOLoPjFQUsGAkJ4Jkpy//
HAw/bp13+qhNeBIH3cvxXQiu8GdogJ51agMDKdg3CeYmus1M/opgvfefedmZ
o3M3fDMBQTE1BTgRHMH9fQLrYMjoRBdnptaF2xOBqT8qt9TJn7VhC1fkvkr2
3jxRoz/NLgZRntS/Esjjasy7XlhcOqditO33FeEnd3N++BA/vCgXh+VXts68
FbfcYUNTCtu6oTHyD8L5NpJrmKX1BRyxHuSDBW8lny7xYvpus3PsTNbRWMsq
HojXDTbqGzjasHfF4hfcgDOSqE6wDwGk2cR4hduaDuHSjboKN4vGjWn+Zfp3
ZbSp3btp8C3VBLnQ7DKIrk7eJl/kShyePP63MkGH5M6sPLd8kovkuNmVAnac
Q+df3tX53pSWyMKjkvg6OM5G3bKu4kkj0VmhMAXy7R6lNJJz2UV9L7pro8Uw
c6RbB5SN6SmNlHWcDDuWVpqBauahheZo2yvHBPna/aNEgfYSOqzl2s2hnhdD
PxQ2+WrYvGHoVyP3X4EQrIzN3qLNqjnuo9dSfsHMVKG5s1Yy0V8LzvfcW3+/
8m1uKwzjUK+4rtHAxvvhoPDkBIJ6MjUqACaoDUDJtq0BcsQ8EQKO1NHcgAH8
TsE11bakn/TfTr/MwIq76cTqoEOZxFiAjesYOCpqL+iw9njTDo0aD2cmTOf5
JM/BMyRYAVHAdbR4f4GOfuPzVl0R8fE7NiUuRPDxTSwV33XVqXVvk+OqMrFZ
0z7ThjIE0vaGxa/ACSX+1DF08xuG3fsLdS660YSh5fhPoLF0HYfdPd6bOITl
J7Vrn+zPQgboqBKvuGhY0eHsA3Xynb5F8/6zLlDq3diZOdG4npVFs7DQ9xIY
4MpwLewJb21C+jI4goj0cWYi2Ma9HizqXcc4mwNWcC8wfncnXdl+4cfB4Q5R
6G7IyMm8QNGxiGTfM3zkW5c0yLBHUmXOqAdnIg67ZUdxq1rumdBHEaEcZYFC
08SvnTBv/CNCLFUg761ZafoKKn/Utb14wOvqHJSRZ/8HncmRISVDKlmhshBG
1r4L5wBnutY6lk/Wq6MMrKl6iDubqWWk6S6Iy8ERMRXaAhAgt8fUrSoYj/Oz
w5V6Y9dzsD91mNI4EZi4RCSOIfTm0hZuLyCRvCtCkm9yHXkUmCmfpMhM7GXe
YPmUbUwSw9YWqpmpINDj471ZC3RcHe6+pyq0FGawkX7JmG0jmvIhuO2FJUjt
RKW+i4xEnYPnPD8MtiRahHqem4mJ6npjmbYBUlLYlisacC89ppaesk48mn7d
N3JvFezh2Ay1ZGiSfR7BcddSiW/YNOIDs7WJeGblK/gox5rMB6MQgnLzCK1T
VyXopVFaf1iBQrDuPG30B0zamCprloMVDaYZt6SlCRofKhSIqg0L6jF5/meK
UPKa9Bp6ML0BPHfJ6ZK/uLrVvFGvUrnafTFgNINmQijz6JL6M80Th0iEaxvD
tcFReDuF/JIegwnRHDb1ZqvpOejolOOmymzE3wOy3JxgC5BDuqgkaMcAO6oS
X2WCwT4rzDhSWjjAKcZW05ANRvpJqqUsKfeAQtySoWR6ncn9mmdfGuWQgE7i
5FhlUJydJaaL/aq3XVvl1YbYTEAqRgSHJ8XQUTVkj9uRTTlelWbk/0bXcl0V
N8P63MC559njW7Omvlzd2c+L3TM0XloiKCx3UESikL74MMSt91FWdFyvddLM
iIZD+ICx+e7BRwxJ9V5aN8AWIa9p+Nx5j5ajbi5AVKWVco29n7KTsIuK3LO2
b5tG5MqxMOGseHcFWtsxArB0XHfNXSOltCVz8JS9k8AkB6Xv8O1g0xHlgbnC
vA37qEE841AoFxRon2C1r1WU5Ju9Qs/FyKQ7O5onA7ZH5/mgHA5Lno882yVB
jXoPway3An0oxdlsNruPPd+OL1nNeZQHZRcBy07LW/OeypzKbGGBCambLDcy
4/jXHdaaO6/VXHG/Oel5gtRbpYt5BKxN8A25eRIZY/DkIhyxE54LHhwjAwb5
fb8dGQyCUuponn5shy5rxFiZepOtF7o6u/WgAVKdYQ50e3dN9ZbFCLjaL9M3
FGlxz1CJVCGOf9cN1cQtwM2OVfV7tY23LohgtEKuHXFu14YHMJ4z6QRin3DL
Uh9+8QUkZXx2XFPPqwMFpi8XPxk68PnR2CHRxYurQCugb+Mqz3VbHoBjTwQD
fjtpyv6Axkd+h7kq3QWYfbSNVDZUQYHq/1KLndXwicZ/tbUmYbbmM+WSem4p
1Z/MKCEksiSwskNrZ5LROMJeKwJzsCA0xVtJgmY9ACtf5bnNdvj+acTwd8WF
bPsekYyki51q+DINCem25gqxJ5NdxbX2Cu/ePCah2gshGVZ8GBGbMp8StUeS
k+8tGWeCPTAYRS2+HAI7NbcBf/IUOjBd3MB7tqblY3fpKSRPD6rPtvGGpNHc
W93ONBr/IBfBrudYzfz6u64XFOw59V9duWyAuYrcP7MnkanA4wFAc8n/y2lF
BkJZDSNO91rsdGl/BGJejqipj8zjzuCJ2j7PAwNl4kxb3J8xY1WPVxCF9JcD
9JicYfEEclFbL3r7xOkAqlgrXlNxIo1M3Ni2P1MCbnbNOfCs+8sFRpbjpUHx
JpSj0x7cTUzxTV7LPjdI4hokrDY/mOtK84szIgoE15lRMthsNUv9SS7xmY4D
8nsGbbmf7tvImXtwjY076pKt0wUwGJOMV8e5aSKoidXc7PNsd4bZ+SEV4MDY
a5ZnFDDZ7GLH0M8rsa0wUZFP9bEkxlBnH9plx61xnNK7DiJqJ7PfgVQF6jdB
I2FbJW3DLx7j7vDBBBbFH9tom1dn7kg0lFwItaxGP5c5ED6aKNET+QFsLaHk
HtKsOhDEVYEq5AIvlBiO20D1IGGY+3cF5rH+5OEVrXe73psHVPPTUBtW3r/m
AYO3N4piB5RSwWanXZNZEddZ7RaLbJGGYR7FufPxhMjAV1mqQ3v84hSAEh7Y
VWZecbJNa1Rvh2qaTuenErIsLpA9Z45WpskV3tOC0AgVy8CIF0yamtpnkHlH
UPMAOOhvF5MK9Xrfk8LvJ7m2MeVn0vhJspltPftJtLe7YlP8y+8QQowvgFQf
LzackKXPVMPEOVbUo7yr10ihvSqfH7fdDnIpErzSRBOhfJr3cMJ5W9P501j5
HO1zl8e+NmMooB/S9UhkiEPWGThBKlOCfC0Jofi/1dqoTLi4o/v/f5ezKCQi
YB0LQCdw48PoVrQ+2XOXBCtlzeaarxCRBXK9d+8hijWI8iY6smDCezpBaedB
jFaheUTh8xYmaEnqZMVTbqKEHZmZiw5qg1BwUBW5sXriX3P8W2HeEUXETr9h
8tL9/oataa+0TuTjfymfPnymzeaBiyGlRQUNvJRc+chSvIbirh8xnhyJkWVB
BjsVnTMuMOVT9bqhLfhD4/Se8lhYgRD5v0tSIBcumnDnAMLaVaQ5zJHynEKk
mFNOPRlbmVs/W+lv1uQ64rZXVbbSyHEcRXubXxU6IdwiLrilBpLVytzTYIdU
EahAf9PuYLbJCnX6rEPD+lW0TKKL6Si4pkxyDpSMOT417w6h6bULO1fzBzFu
G96S8Ap1gZ+fFy6t62c7CXN8N6K7EemXGBguFuKCjL65YhRuWEqS1uH/Yxt9
f8sLTyJP4Av+GwE17TTE8aH0oaLa7kv/RfbpHnQfhHgxKthWQ7x8tYcE5hMh
DrPktdAyUNDC9a63LBfuNNuczQWk/ak5F9311q2ARUf8E4gwjoXIxu1x+Fev
8JC4rQpNYW5W/kLXs99hP/vw0pjfRUka2lhhq7GnzDj5p/lTL6n9qedWqg5w
7/kJD2ZPdhJTqqzFEjb58Bb+5jJbP3RySFbTxe8uR6BnSo5JMzaD6vKGLR/p
ZJrppMhJJQIiBgaO1kiDWwFcT7aFSTOiuA7VQqP5C0vQqIdL1UUJPzR56enS
ChsI6BGbgQVjWmkPDcZIelaEgR5TzIV6SmGV04aiz1olVKplcjx2oViEEo90
Pw9Ri43dTF5ptyfoj+CFuhGKcKbRcNu6RV4zcMkxRS2saVHxwytCBrFt6BGX
rhKA/4RIRKnVpJzGCbWeH+29GqLJmQUmAYgFGdcwqVJNfxnbpyK0agabeicn
YTMboIaXCTAUirpVy/78xoNMHliRhymrSuWXaBuUzeECCudLN/mEtYYl7Emv
j9j1hn96I3pYWEKDgQFrxAURhHoVx5irNZiDud17O0iiz4ifUbdnOk73ItiG
OajiL0UU+1lAWkSincw9IMkYgwywpDxw6E0J/Ej1+nETTncaR7TB3wT+JaNm
MNsKK278Ka2Z6/wBpEJJ5Wmc5nsMmqySYIIwfbQtpB5XnnVsaTH1JrZ14rL2
HPG4SIiRTkN4RDwagifed8cpgj4+//K2hRYq5sMibADWgWvfgrLpf5bheKFC
EaO1yFrEXfyvPCNkgGWkjDPHRsNaM6pUhrel5V/TBt8hvmg7+EWFks0impzd
cKwIjCPMLOJeCWr62XgEcDOBCyms56qI0sGJU7ZEMfgqlbFElBzCJWROtX8L
+YjERoYzRwdl6yf5qzf3/K0N2OHJBn8usodJ13DdbdX3Cus7ii4iUw2UXWcL
WIGX2VUVzDwe3iccT5DjuM16utuRr2BOe6lHen7Msg9cmPUbvLomQrmUqxnm
p9HKXUelQ6Dqna9exiaEnOK//OePo4YcJNXOnapTrV7+Nm9l99Ox+UqqB+eX
dHBTpZiGjlPT4L2BhtrOQmUR6KKznUsjujhvLDDXC6pNhdGFMWbKT3KtNCGw
Zs3d2nV+QTmvACx0qz46eGQXFbB1B9Zx5QF1WoB4rIfV4OG/7AScjSOjHzVS
xaMaqAdCoYCgJNJg1Ailx9JWj9HUSa/T4tWkL4XO2M1+fxhVehkGZG3T17A0
G0rqd8muOxZDJqwh3041sTFo1FfbGgpXbGZa5cpT53pKyxikkBK0eFxgU60y
bPWGCIpZvzH3YAszHeLOabthZq2q/fndoi88SEEMaFJMCx2TEqMtIdHkQyyq
bIZDtsH8c4FksHM2v8gicQcM2iRDeSRIN5koHNUIPb/tjYLs18u9c+D3GP4d
rlHfO7DyGg5X22Fd73J1k0MTrmVvU5mSoo/y9AiXd6e+M+gCSdTIhk4hFqTY
vyH6rpapPjizQD9S7DTKDSvjLDLjPL5HfFlA7zO+tpbXf4da9/Sqdff087SW
k0QA9P23t909pW752ODT9fcDnYr8BBHIujVkvNaJU6e1RHf6qvylxnZTBrs9
98+nJN1ZBVbC+7nHnVHsBtwQGaOYerHdaPWTStjHjMO2z/0u1Py7u3g4dSNH
XEdJgYt/ucbWrgJk28mxZzT5jw+07P2BvRvn1UeeB0vmdMo9OMtB823Yjq2M
CbWzudCJnHpP9RrjWXiRgKZX4nLXsOvF49wlmuL9ISqBePu8OPvpAHWeTHh2
SLsk1SuSQqcEg9pRUUB1bYETP/l8+uAQbxL20yNB3WoY0wniP0WWtvZmv2/9
TTK+LtvFllfpogGePmhADFVAhwgKdSDocq6eh0P8qo1dvSRXi6laAlfqTwXu
z5dlco2KsWzQNLNJRlzfc4a0A06YDj4GjSGTK/J7bVGn2HinlyQrYt+e46PW
sY1QArKxLLOsbYuN/rAuys/SHn+xxIfVz+CvFhY8l8DTcTCupt9ZRfA4Pv6k
uvPXAQEqynn0RJ8GHw1U9TGOgTMp4h7RgxnGRlnX+YhAWDwE/C+lxqVirem/
6kdcKbL8ZNz7ix7yHSJQksDxECodrzJkcbBlqAu2swQ8zVmn1a50zAHbqFhM
9g4E2PmA3K6T2Tq4PXDqsrEGcWvvpZpCf/JxLnLkd4yByv5mRSlBAWC6PK7e
UI7jyE8CAPbW5/KiRvmqlPQqFH/57EAjqAxKNgqvoaI6Thi25BqjrSrtwe3G
k0tnFWrWfEHpG8UWJQh+UbjY1y1J1ThPF0LDaudlRPRwouWhuWTbkT0xkOOQ
e8uZzlUJGxPTZdWW5nI1zz1pEIsbljsJWk3zVL8B6TSm0eSwSMGVRNJBR6bj
kF8y42NYX91zvOL5xUDu4siZlSfTmfJI6Qq4D+j8YvxI/SFA0bFB/UuT3r0c
FXROex6HZZ+enauh66/F4Nt28iPcIQGrjQxq1RCixl8B9OX9TMHOHqJNp++O
yUG7TNn3Ej3uusqVM4iJDeaXrLLZZ7rMMzrGhdh1tNVR/XejqYF+1ugZT3l5
LfHBB3JVztq8Zsjk2AzY/t6qSfP1jsDJT8/wbyoVQ9adN53WShKRfmwGLHMW
nlV8N26aVwOBJ9VOZR4TTDsoAbsM0yrtWWUHiL8Qyl5cdL5vME6HeDYLwWFV
5DDbpueT9qHpEU3Fq8f5uJNk/3KSkH3xJDm1cx+R7MIgb0rVRWKXlEFfJmuq
dCsaL9cfbagUHFunyeP3d3mOCU4dhHXyLkJ3T7MzJrgtrrpYBSvlTZeaJjgu
jT8VIbWjyMnYRxfQVzkcbDGPr48Lp1JtmlJpDINDiDwz+WQ33lYs8Tdy5SvT
4cCQ3qu8SEgi+HX+35ooCtTvDwT8/KcyynMtObvJ6cwO0XQu9hXMQBPpz9nP
jqj60lLkJa4WDtPNt9kj9UhK0s7yznHWe05eQcwPzud+iPVu+8SjRjuzQrF3
ZqcqvLB4gG3j0GMjVztV45bFMAHTCKyRQAEiNSRhiiBEuMpE1De9A2HW1L02
BJW5kBz9LdjzqgmvcQPFSr7zNLLzKhUYa9X/qS7xVarpON0HXVnOVF9E4U4Q
rmoMtGsYJNMx2VdvUjGP5Amo63k2rTAJbDTSknd6XTwiHqxBWBXhOPnZb128
Ex3ITSzs/XAPdKHi68mrFuVw/Ipn8xZzwKU/Y7ujHwr66NDC6qBgaPUmShLS
qLCCvXbecnOpplPLHas93Dvq3GcQ9nU04LaS1LeDgYnLxNyCHen8FxUQc+aG
gHFLaJxhpukaDepBE/lwJxVK/dP6J/+uN+kjfL2oXzqnrltvCPo29QD53P0Z
XBEDb+Oykx0WrHYlL5H/ro20lsJH3hUOqwsNV3DducIQlUXwO1nZd4TaNyiJ
R+1QWFCQ2tqHA0KXt6/GhDxqaVBFQta1oOwS/+CoIRhf4/FOxOWWcge+a7/x
mPW+V56lTyjUb15EmfKnjXvmiYTRApll9GSLnuX3RVT3quK/5hhg507TlgKD
HdpX5u1DU8J4xGs8YM7wwHNQ0RQDndCTrBeCouQHaIhdaMKJrNZ3L6A+a26R
9PgcMl9tSLNmC8I/dmeACiC+g8zxjBRftmQo6Ucjmk7L8VbLmmrPKBRf2adk
EqPoX90bBHblJ4fMwoTptYE72K9wp2Y5Wm1+GAKGwvpX2drj4AnI+HBGz66d
yayymXLZdqN85EV4h96JxrviO7OzQ4qOMA4QP/plFWMGFIk6OIgAQAFV/f/K
Jsp6mAVGvJV94MBpinoyhjf0wByXpbBLhENv0P/KYf/SIMTxma53rUTqi29P
dGJARqvmaItMj3sv/SLms38OfSL/M7Ebs0SMLvB43jEqEhVKvZ4p975NiVOI
mxUpLq9LFhHM0MyitZczqCOEZMeA4MEbLcl3Mpp2LLrTn0yhsBF8o9NrD2gJ
VYPA5zJNk8CpOy5LZelzDQAskGyGX3kIxSEiaoWAiNSemoz9oLmQN01k1s2w
93dv1BS1LQ8j7K+4tKnRBUxzF+LVcxrsFeDkaQXtu07cjtdCM8Q89nEzkwly
IFND090BvCXrfaY3vWQirY1ZE7M1mTxidH3hOtoywiz/HCVhrUibqo7lvMl4
I8dJAPOHJHLiALGRF2oaKf2t6SpmHovxEKDK/sr0AwYOmTKnK8pWYFsPDTQz
rjiNSHyIf6ApbvcMgzczz0zHf4fUXtMIhuJ4S1W26sEhuQakOPaZGhZW3Y21
gDK8+ubgD4FA+KKGtnVYjwth8JfolKWcVnJ9PnmXN5ctmdSPE1OPv9aH5DgL
BSbU/BLqI6x5UdIemOjIt1eTlEZIjJ9NJU/tpHjnE+nNCf/oyAOE83WkadGA
PFgVKVAUe1x/v2a4+hRbXUrocPQHSFnHrQAHYc/kAYOt5neM3xIHrWSjjk/h
50SGlYOSB5sy6WgrR35JkXxHYsUcrcCkQddFJJAMhWmkXRFVD6pppw4wM2WH
3xx1TYzEU3hBnDN8goU4ZH6EzPsTv8EDi3tYaA06mpuIQLSvB7FdIf4/KWzZ
nCnStVOyn7l77Nq3k9xaKjVA4sgO7EmY4nsqxieHiA0v2nIAeNSg0KDRbO/s
0NAp0V9QTtxk0hIrkA0v44TWyJMfn8MYOi/10EbW+dVZlwEb4DCwd2Qh8P6f
GJ/J9MqPLWduAICm2ienFr1UpiRg0kFNgnXjdKSShVSkZxCg4k4huVdgqDXR
3mlXIT2tEL77G5HyymzK6SzCsT9Y+IZCS9B0itj4ba9hIw9O66nlRlKtvaVV
FcPIef+f0uRLxgnJ4OEfZEfqRPtvzCcI7a/6VjlMsYbWRzt2RIYQplThHc72
cCIeh0A66i2vU8yydTo1amAj/jRHKHqZXB6BnBpBtMqIQ8jDgMPBf7YXJgxE
ZiqwV7i1lJ0Cmlj3SuFeFVhpwOznmTYmzCekz08n5M1SNpYZZD98eK8QId+R
Au+eND4aJYx8Q1/soyYOfhcbnsZkhrRVmeDFncD+pXXiHOFA+cc+2pWlq53N
w9iN8xs0yHp5wt2oMfoXUEEJ0a3zez4x4ljIv1RIN4HzAKkHk0XAbKuBAVBE
j9rY/fhaegktZnB1vMnqrNVCnOo/Sm+KGGyt+9L5xol+mLYad6mYlZwwPKqF
DMkiPuqOyUtVKQhR4cQVvRMEco8nV6pxM5c6eanQUMHmS/jvhmRjw9EZx+cI
AbaWa8ARib9o55ZfVrNUfnmS8jH49UTkT2H+S+yUWPgyCSSutJ1JlC333Flj
JFs0eSlwz2+6j+yJwrgP0Qkf8hQRKLBcqwZA81C5dOxk9S9fVC8nkQhenxI6
HcR/z6LVEq8RNOCTaIFhUq5M5ZMDfRh70YyX/Va2iP+xHXWB6v9BUmTRDwMq
BS/dOZWOMvBzfm0jz2vAOLCdTGfOV5baJp8dwkrfhPH0oD1ngFFh2DdgLutQ
nVZvcRTVP7B17KkrMX6Ikxp0RKM6u+lmSKbgj2CtamgC8Zs0Tg37AhjxPCh9
9+sO3FoDXX5gNt2dJkg7svqb3ynqxOTDyHp4SmxJIjM2w9YtNaFA/cNQoQdg
rtMgyaadzgyrSEGCgl1y7xzpRyW2K/QNEdB3sq2Nn7P0l13lOQVYLeqNl1Fc
NX27L86agH8rPkiXt63BZalrMdRFpR7bIKxZj2Utt7WoOZywCICnSAElhBCl
fpQJzZcSheDzDRXczp2IyNrsCvLniTYtOnmXpYdcoNVbTuJVkWzHoxH8/AnL
mwNj+DZ2sezxkXBIw8ZqjpbRPQOwLTnS4+jyi9TN0UuCS9j8+XnL1q36CUgy
qobIaHNlbBqEhxfXvbfRvOpmim7T6FXh5LhVSA3jqvnd1b7/xk4Gw0GeCoT1
FS0hNPw8xOTLdvuTrP4WC7TlIst56Y7Gy+aiFValkcer9HcfTCkVWF0z3AQO
Nqr93u/rGDllMQpRK3JLXtDc5tQrfStBrzlh03JK6ykY8UWmY8xjSTx2syOp
y3wytvWoiR4q2VPTeoNLa8Pydh0l+dbuhuFb65FcxRd7bOpdbDbdgD4JTLvB
fQMRUDUqNqfIKdTGL2E34PtUUMatD9q2XjWt5002IB3pxm+v9YuJtUULOiDb
A1/JX1qy6MElKbjlpD7lFSJS1wdlUpEmkt0IV7T0e49+pUWd/ugIR2jOZEr4
vPc+Kjc/JGDNOmFzQAS4jMUofb9O5gpeLQ3gDSM2yx0M7UrWfBdCRNGEnc1c
7ylNW8/EWj+d1hYVsq9r9sqzoDmFPBw8cYvh1N4IZT3zZqcC0YKIbRXLFTPe
Y+qlt6vTStjCQ5nIeXzJ5pDBb8tyzG1O0+nUGy++ZeVbdbjV27Cc8g/LFj4H
2isH27ij+Rh3IrSWjKFZrH3aQHZSaB7DQc2OLDIfsK8nOI+mi+dJIXR5xO4E
POMhhnAme+0SLvr6DWeYSQk8wfbfohH/zTMCU4bbhFJOX25PQZDemztMTdEd
lT7vptU9bdSti16Q5s9yzeCWWD9GjPSRvDrKnp6jHIYbh5wJ44RnDf/XLoNL
m9UZt9NPxMNONqas6wuXXMVtbIN4CeNljAhAnGlzU+qIzFN7E8ux6LXJ70Y5
Yk6h0zBGOs3ZfQbY9ID7xMu8vGp7JYmX9aoKfNtMLSGtJV/vtMKJbpEqt4A+
pdKRP1jDH1f/TSWNveLc1ek1w/Vvo4xUtdeaWOvMnWsav+Ad4RgyPG4MMHT8
Zw9IzFI93lpDDYOxw521t2EDcjYlWffqhCrdEERDg6I/2g6S1xT3e5WZFXOn
P113XZ76Q2YmKZ5h+Aut2OBxhdICh8MshcXLqNhY618LxtaJf+Ql2YDkgZmG
ntflTqY7glp5ehGRL0tw2+m0YsfZRFrfCcQGVsB2KROGn54/gd1j8IwMwH0I
0Gf2a1UMuE1gVWNVs9sxt+5PlarnbL/1TwFDo3oBq5vhpK2nznxFTeEQ4rMa
FFpydQnzYXXBim8yb5HxP9r5I5O3xSQeUgjO63uSeFwuj1YvzfGGk7uxpHzM
zi1WbVC2fdhpu5o+oVTemNDron+WimdTMKw4pM3e3A8Wq+CL+ENnRdZCFPjX
ivQxtN9AkTqXFAGB5evVjeM4VMRUah8qoW6xUuzHwhgWKmuhJYaby9WITySs
Mt4WbSW/d92Gotze+TH114am2JQLZz/2OVFphp8XSEBkFYF+sgCFWTbtOCSe
q4kQ7u5V2/uXNVP8c9Y2HiX0DS1h1c7Vi8anexWxGD3BWoUm+zLV7vTrlZww
mV2JyD2U8NeoRvQ3vE8l9RM78QjEPi99mh2TaqIAPm1mMMxEAePOOzr57zyH
ym805YAl70rksqP1/gYD81nYgMr8IrYaVLYVJoZx6pWjFjBzWNNeXIHOMwfu
ed8gMK3IWnGU92k76iR4IGB+i3UB3wH0zo9R3BndMh9jNXanJ1lP5+Pj+8LM
ODl6p9MsanqL2VOpmhvMm5jkoPrPboshwThom0u2fS6qompqz+dkUJ9pjnJ0
dkAdqcSQyvQzhd6TnrmsANJvwPwNGvRFBHZslVduqwrSRLELYze/2dJakO8c
of3T9KvVVZUP99n2zVUF+wt/xZV/4Gv3e+24ay/TdfNNybr6pdY7hdd7omfj
rtdeT+dBgd7Ob6JdgQEsQw/+FRvFUJwKAm9ZInPbd6oYSJzFxGc7W+GND6yX
ybMStIlB1fn6/9KOaEy8ntRCJig8BGfGLatdft0Jz5LAAIgzJfbde+s3EJsL
CdumAqpirzkRZaJrttkinXgefpg5uSxlhoILCjzxLaMm1q0sVuHYH1zgPhxq
Ezn0sHSfJOBcuxLoHNAwviH6zF49Br/vTRuZ/7dzK42OrD1gUbJ44razI1pD
fJphPfEBmB81W149F7lPIkfKY7WQQbN2988Q/KB4yGdMH3bQKeshr6wc7IBr
7YzvLQ3Xm6HCIVeLYnDSFsBaNqr6YMEiBtRxPRGMvKaYcPXEdncTgCkhk7SR
/zsvYescS6xwNz7aLPZwfjZ/kxUs5Dt1bhyE0Lxfu5hoi4qkB49RCTQaVgfH
Y4weFNCMSmcvz98TsjgHiKx7ZbSCaD8z4TeGfxbqBgHMjXszrCvmKH69VPrW
IP5r8VAfHvEvnt7hAjIviw2U6i4iNZoEldKwsaRU6e+/FXkks346hFFAJysL
gyRu8afI8K1GUiPn0JZ0ZDhwILexS4ySt3ZLxttz//Piok3ZB/jcbmgTWpn1
pKhj0hMbE3MHWUrGtu8x8BH4+lhmqbnZ2+fOOEeD6HrraEa60Ae1hYdLDG5C
2k7HLsrOkdZth4gAdidHb5ASlYgevX5yUpZ+lXZmXiU1nyp/6gBYoDexS/5S
iqUvMzBXPkJ6hS2oW547ILKwl3xzDf+GoyxIuvNA1D1bOyAZuvpdaJ/HEHfk
VQzha7vjB8qyUlp+2ulzWFsnlhw9symER/371ggytdUPiC751DLhO/v3Es6N
0juTbyK/PFWQzCmVF7r+Im/0uFJ66zFO8JMWNrEb8t1voTFPE+Lw0PGbEte7
MQLdujOc0CicXxcbyEEX+YZ0ZzZC4SFKuQbFGhZmLZmEnZlUMcJCwReU7yt7
OXKab36X0FwvSgiw7ByvTP1T2bFQC1HymncO7K/EnEpk0GZ1ryO010LLfzzc
S3TiluvBoShplDG0Fds8l7eWZ7S5Vkh+PhxbyDBPSyFtzTCRFVxBsozFk8eo
5POBAwXpbb58IX1oVFmEBo3xZLjhWn0+v9Cdv2BpZXgcuQ8MSx2HNMrDWPB/
BaJ+JdJMaTDaT333jE6mfS/DG7nFHLKycDKyK4r+FMuDSkwBRtsoOklqlDff
agt8A2Yzl1MrvALPuRhnq5s/G4XawAnxdwXTdiYDrHintY5mRbWB97I7v1ej
lpY2d1GpFz34gXCxUk6BqdeOxKeZB/7cG2phN8FRV52iNBTJx7UQo9KnhCcU
16Qvhr+4ctwoDDcXOLl9IWjwIDFhmhSb50EuGASWl8rE9Tkh53oFqomIHSL6
eKKdVPlrcilEOQTrRG3FCAWMxOvym6gPXi1kC3UYlFLe8UHMLDdDf2EfKFzp
EirsVe5PkmXSi2f1LqoXTgyXuHsGMl5WrkSt3mtouDFVUvgt9Ni9BGPqtUwv
owzJmYekCkGWZM/ahjbRcEn7JFSF/1MTuTw3N+6N/CMUPGu66u28Wk2q26Ds
kXf+BCp5WJKvA2IZ8NJPb67m6h2gqZwS+1VnYkWOW97mu6S521QPBI6RVO58
dUfj0y1ulvpLFq8f5Ou3k4ngSISq7/VZIfZTDJ/tnja9Hp7wHFWdoPCFaeDw
kAc7kxfdmCXhgJmLAIrAGGCUqkHQ0BfwAIt0JsF1Y7zoe7xS6AvefSi12G0c
rA8nmDn0bkt8vuMiZnTCc3ZKxgh085+dGXWnca7N4urjwWMO9ZY5CqdJK9TV
rKP98EkNbWXQqrZmV8Yo7ZZqD+qiru48atCvkd1Dvxbh12IasAlNV7e0Hpkz
d3wc677E/6s90IfnwRPuNxc/7m1AQ1r79FGI2IVV+li6N9pEIQwY5QhddPRK
3FJOa08uQTI6v0q+CzREKjRkrmgOTyTtc7bwqCJv9sDQb5m+E86zaGxI4UHV
8/yW0qFHF+1CKmfHgU9Eihlx9VRSQZS9Asnt0ZCJTqkcJD7dDX9CcS4B7pmL
6I2j3Q1FE4wp7py1EuivT159t7eOO3hVazVMvxylSQkysxizHXBgfVSGrJX7
B/ajbv8Fr/U/u9Mn3kpvIeapibAYTGOB8kDLTj6AUv1v22iPBGKFSrkG9wV/
l9pEF4YeRLHP18MJP+wVUHVZ1CSI9ElWuS4FrR+L8v5Io4xzGJhsKujPubTE
o/v5AtqLvzXR7vrgS3pp3Ge4DWkm1/aYjDxnukxAbZXfmoIV6wnwdav6UwlP
+Hon7oGIq6IrT+i7ZZnBsFDZ4rPUu4RsEMK2a4jGdjtCtr/YG9o/hiQPs3rc
dL/Y1Atr7SIrbW1RvQ9jPoM60TbGn9TELzgRDMJQpqbPYh9tigUaRM3YdJcl
dvNLnJqfQOpnS8ugJMD+6xxCxQxSI+poyB33gNVMjiY3LR5AsYVGv408mYjZ
fmxTcGb7fTP+ke5y05WtKW6t/0dI9Hl/zCzDP+N9jNQ+NEvLEJlb4L4h7wJi
OaqGFoqJe6M/KM0oHNfK1SfLa2dSBqOCKpHPdnVmPVDoizq7KTaXBtEiWJmI
uM/Uq3VPJ6hCK8rVo7rOpDs43u1Q7s3ed+broVYS9Ze5xzfIgORpDRN/JeDd
MObEam4sN7/mewbOoWV1FAVA5ywvvAL1nqmsxBOiTfBfsvPDGgtGbIi7jW/G
LVdZjo1CpE8z8pjObk8y4RjoA/aJtQ6qPaiHU7sk2XekQAnVQroGOr2EPRTJ
ASiR58FKM01OFiw7wYj8Uqbhz3IERGp5QNMzOgZOeZ+NFtC0D+XgN6sqhWNH
WJM4Qqhv5cAQh6Y7O3Ohfy7cfgKNxr7IkOnSLmRa7wZVIgak9xR1Lws1jvWw
qQ7Pqk7byWe0exl2IbIdyQ+M4qC55fZBoel8I3UBcgyETYoFM9hGHcY5Am9O
RtRGfT8EOj1y19A2VyoP2X7KarQToi4snfN2k02H8BoY0nUoSSLwoscNPrSm
mCDwGwVRY6euh/7cQIGJ0q9pDvJKCmC7KrU/3sim/bUyY9elV2JRdO8hVVa8
67yoKoiB2mjr6V4wTwPybkpodNBHY1sSMmltuNte0XlzEr/kqBt8spiYC7qL
xwvJ55Y/B5Sjcd8sCZghl6IXxFcFJNnZxBCj4AVRxuwss4gq+oeki6fzRH7Z
vMfaZTsnsKBP+CnrmvwaX+YdrxDcKx9SzGbgNUA5lEE4NWfw28w1/mf89JNw
Tq1Ex1kA7ruH0PTw358/f4JopkxuT5roLpWu77DrlsLwr+d3g2KbZatpqz/J
IZo9NwRFGxQkl1CM4Du0l83z77M+cKQoV5nh3k8G87dFFn0frvhbsgwrhnB+
wFNRyPbaH7FJnTi0JRN+nZJit80SGtVJ3rZ119XVqOY9Q2WqxhJk7I6nbtKd
xUVUq5XH697wILjVBCH17Jy/lpP2gDQPnng4i8B8gzlS8ex2mM55g29oxZtT
hgq7agUe+nlhN8Is1Go4YRWcpHXbz/o2co4TtbPlcqO1S11Dgfduhu57ADE2
EyVMzF1qS02qanjVi7EA7A2B7mBtxPB+X8orR2EV11KBFX9ZEI/fEWtTMxDD
XhkAb7F6V3s1DCztA2OFL0wzblSNEsWmH4NJjX6L2k7y1zJ6vb0qj/DnKQp4
5OEGIVj8Q9kITIy0+ulS9eYxmXEPTaM4BaaGo09F4q7VXogZ3Vtd1a7Pzajg
ighnwYOQzprbLOoEDEqpCJ5M7xfkU03kl/43A0BwVyE12puiOGUupuTXImud
OI8pFpvAPHvtxaZQCxz5269IunSPLDbdA4XYZUbXCSI3wyWG4DxeI6ACziBF
PKbuMWINHDQwkVZeqzkX05SLMmfVMwBzKUr6US7kV24hniR8MNGq6K+Ez4p7
nXMC4+jhLl7nhtQ/4z4d28cZo3ZUjyTP4rOqDr0TFRbRgu/tZllOdNTDKb9U
jsCSk1XGJdWLqSSuJpkf9JLkSxuijHVDEkde2HJC1udsf5RXdB9T17CEwodx
rjSEyLJ3hbK9K3QNVV7YOQwZypc6++5L15tXo6Sfpf25xNSxJwpp7tQjze3e
f26I5CgVA2YKcrj7vdSz+9iUHtUiBS8xI+6NTZYq+u3fcS8+8MyeBcrLiHZs
8jv/t6AT3OcUjO6dvEAKJZgMzIgUL7sIjZnbzuWgjTu5Yx18HJr19v3LgiEG
5ajSnvMmIbCCw4eKIh0sj4Vx+zZdXkSYU7Wt30s1ZwJiL08HJldtqAFceuje
ruqi1wXdAtYEl79JbbvlGonkmNp5l85qgZB8B9oqU1T5Z5CIkhJ1BAMtvRMc
/d93PLkKi/2t6bfamzu5U1MBlmVErQU22vlYWklxOczUea06tm2Xq66mRZyY
kHcRm912d+PHuiD+l3a9l97LWJhbZTYNTEk3jpqCroQ+VQxKYZMr3qxn6wLx
EhYlq/UqkDCJkHWmdpMwVQSV7mzOFeUgz7Mor1+iSCq5DwbHrWazXbSAfpJi
UoMwOBHk8D3yOgrQGrBke5dpIBS9uqNQzjEYSWsEH9+C5WpvjUXsNPM4M/9R
C9Yzsyt5uKBJIuZ8wf9dPuC+Y1nEvMELjWxLmEPx6Eb/V7vNZyCFiy6qMX8U
VQ3oZkphjxE467JrgT/eu+jJVQ8ToGTg99bA0PHaiVvLS95Vu2431/9eXfS8
pvNyAG8wdMcbNKDHK6Deuw/8aMZuTlZPsIT5Qw89kfR79U+WCPTwFvSYn4YJ
u61BiIOMHhKsDERB+Zvs7rSO1G9+you9HLHryhy2rv9H3DfsU6wgzfti6+lO
AA6ABt7xb5V5un+0vG5YzVzuxrWKD9ge4z14Dfyx6zJjdvLUvPsRmKLpEy14
kLk7zgDf1OmDQhO2NxBXvWlSFAg5eSHGp2IWixK+5iKG4OZ75yfLeXi/8NSp
rZTtgG+f44vxFKSEOuwJX8IR60gDd5yrymKKtPVaa4dO149xq+L228jheKxR
7PFUvQexH9P3zpwSV29rLiAbXxBhzn8uWnStf2hjSVBxQYlb7o7TzpDo3E0z
6qGZt5cYBKb/qWzYuBk8k2Py0CtGduJ5KzfztDWT4MRuny9pUqwKXpQaB7JU
R5a2vct+VQcWck756a5s6zRznBc/D3NBcm3fM6YJnSxbxmS76s+Df76zj1uI
kb3KBz6bMW+j3FYYz8soQaloxgsJsWHlz0ZeYbb3lxJVBc+y1bc71vp90Hzn
vl62Lj2yurh+jNW/lc6qxpFdu8boM7aIw8xCwEbt4m3XzRW0txaHwJr8JPnS
ZdQdO7B3muH9pwg7QvKVc0LyZ+0H1TI0l6XroD+ClylAYlXJOeIxBmwuFboj
GL1S4Y5F6zbS3ksIn8wSRI5GcZ6G4/ThYeV3DuiyvJ9iREZ+ME02JlZJXg9j
J5gTE/fhopYmnNOE4tSYE3uhZBdy07b5jmySQUv7dZn5IGIwRT9u/pzxGTqy
uQbHRLSFtEBRvgXQybOuaZBX7xkMkPAtUrCitBrYKmnnKrvhUtbagjG3rleU
guRFaHgWQQ8R++yy+qM/xBs9mu0M84zL3GFjglWE/vCWrmmbNsTen9c0xkRZ
SYq0z/9rtHBOunar3MtV2GGgK+Huu+vMgwmkLi8Dpx/BnPr/2rf5C6zyhNj2
V1yuekp1AumT1CdOtebKoUDRI8RkYYB64z/PfDCBdCPZBIWWh4mdQWhG7Dz1
8Gd5B0biaprpII5BtCXZtWtCD+pRpx5X6ctVe1gP7jRt10vYapk09uUSVT5N
p0TfHjOBBVPO0ibncOdHvpimc8cZOIWEDpILD+evV6hZwhS3p5SFzRPFm/gb
cl3FkKqlkbnezBGl1ucIiYV41ks3Z18MUUWIH56C2pWHeUdkaTckIaiu7Aol
VIbEfJbW56A/DPYajaZxHn/1QieJu29Uy3lSmlnb1kOC94faFVQ4ST3NsuLl
6sElptgxOrIUlyj2tHwOFgScBZFZEqjvvp1Qnf14pp2quqs7n/hhSO7ERwCk
jcLEXyBmAdsGdJ6qFbl2dl0QzYKWlqVeHDWoPKtvDLMlPegdwuvRLp3s/RmA
R23+k96m8thSH/tz8nxrjo7fRIF820iq/CoGt1JR0xHrM0p2w9+K+xFzrz9q
O6x7n5e9Rpda7ogVEE1cCjkO53nZ/EKOU3w0UFkTq7tMWMqCkgM+FxkQn4Jz
+mOBMJmXZLOQ72Rw8Dp9xYJ1Os4Wg1hy9QeP7O34KTSLjYLoWm5e5dSxVi6P
fmsAQpJSL6F66lxDyIprramP1SMTgoKiZ6N9E206dCLdt1gU/C6NA41hA4o1
AT2TsOtv4Np4GDYLQt6Zw8VriPMZu9tKb75pxpgchqoT+C2K1Ab+O8AYXvDU
t86rMLRTFSChRN1Fi+T6GDQosqOPtQZP6h44W/uy3UCWC8M302Kt2cDagFlW
trfp/ny+eIjFpaFq/0CsfGeDUI2rudyWP+Q2zDUPH7m03au/2NAmVcl6VjiS
muCKNHRnSWIWiR5SAAIlJO9wgQMkDqjg3hiLOCCs0z0UzEyMsF9ifYJTdHuz
q74KLNieZcfoP5xqQuALcRjcHmWuRpvVKfRBzjKv0WjJN9buXLaX6OdDVgpZ
p7zo9yYKKHbYPlfhYXS81qTcR9XpTNYd4mk7E0iqwrPN6Yi3d0ByizUsv0pb
ktVESVCKQwCJxvopixmo6H+lLC5K7NLX7Qjb0WCQI/En9DBtEvTAGGXI6gQz
a2JEsDwrfgGocw6+tI+4GwlyJ8N+Lk379bljVlapTviHPaL6jF/DsbiETThq
5YmXhf/A0UEMwZnvBWINGPwbFaubCTobIMAQwNkzkq4LY7jCCVZGT8OkzHV8
KSkCpq4ZOMzM9WgXDphyAlH0gxV5mPM66zJ99Tke8yPz+GLMn1b9S0merM44
C+/XPL8cfi0JogORI5J8D5hdfyM3uTb8ADT7kBvmUWHpIgld97CUBVDAT51X
43tFfe5frLvsL1iM0xFauD3PIHAqKi1tvmbm5N979b9LADPqRFozjbzRdpzY
ANAngmz5r5s93tTHdUNJ+j3Ehns3ofIDBgjVACi9NskBHDSQ9z/OJULvXO/H
qA5oLfnDvFL07vu55GZ/0qz02iHDHlKM997Dt24jn2/NJgRPNfx8zmGHCLsD
IHZ02LlHdBtOp/ltddfTDkZDkNpLxrXWaEx2WXFFRmrjBxs4ZRuqYzmaIgCN
tfrQRhRCDYk7FumoGSIYFlk2lg4fC7nARp4wFhS4O5PBuEvDnx4JBRAAClHg
dzh8waQAHuEVs+YpzU2/BcyqAkVCk28fXc73CnQukvGEeZQJOUCq+LRspu7S
+aPiO86N3/R9qAZABkzn89Y0Hv2eUH64WhtHw7C+9ON343UH4S5dsqdkVeSY
N5TYZ38ZpyqnedALBYbIzaFfzi5kHi4roLYNVKZHaGg4uD4TsvKZ9l2pPJ/F
+XhqSc6XOo+ozaIkk8435ammiVn+cdcVBUGk3sGeCGb04zyEen+yrHUDoNRK
TSJ2NkIHNvCLhTlluxdLLxRW9U2fw02KPYa++nYd6sYYVR1EjWCyjqsmafDT
44D0vcEzhI5S/bMFHXbuQ4rkuAOxmmrex1Vm5bLqDE18GVNaYYHwJUD7cexL
5smRqeS/l3d5ZLivJzLBK3Ic5NuoPhezF/5iwrdCNRvPlOVQHgnqT8warLOH
uUmBeLmcQjCY+8CW5plRwG7A4z2Wjv55GBQeDh1Tth2NbzApsO5UWbpbpinr
t5CaDRDxSqmFthvDgVTTFwGDzltbt3VsEoywpwRzVeoyxQ7gWyGX4bMOR24T
MoTlkb/FYYer3Dcb+BdtsNtPyHcafJcyY1917MSi0v6uNqOtG3ZIFZl+saWk
P9cpqik+b8hL3OgpILM5eU9jgWSb02HIpWflolMHxmp+E4cp0cVTghdEGLVE
nLbI+raoo3l/t6iuw5H/JArYE0v2TaH7+BAh39E4rZGy+ONKA2OBrOW+RghZ
whrvOU7/Wn8aEWzcrdSNLdNgMOHQNaM4xXz+Dnpbcm/oudKNbYCsvhT31SVb
pG6GVumTH0hugp31a1KAcGeNNjW4CDlq3dLesKcHi8HtAamxlyJYnOxy30Q/
XTndETc7m1sD8f5vfOOiW8GNaNhowkweG1CsBY8R+2KjSY+RR1KeHSa39FCP
PEROHbCcS9ZfP8WkbBF982XTi0W7C8wCV7J5ED8DGxtDJQo1Eg21kqmMEex6
R7T/a9F9R+0/nfBCeaC+56m8wCia+fDkHuWB0rcM4h5AhMARB/wFmAUAp/t4
jc+QIb0vXW1KZjke7sTarETjb1MHiqNKHGvX1BPVUGEpoR5rB54jLUK6eSca
YKbR73BuDfUt8TX/H23H7nENMSzy4E1eeSCshPjSRO9Ohe+5ExQ4FVFsc2gJ
bFWyAqBaKMCjiSt7GimzuHPVdXdfi/x0mLKl/HCGwK1LcY4cAwwbutctemyh
jJbYCm/QaAVvj6IyrDOGYZsIHm9mIEsm/E9AFpmEIbgy8+phkFPDDdJrOFGU
hdh4sU9GyI06BKn9uc3hQbHmJs4hfP4yFYILReXgzowiIQLcHFIjBjlAHF+G
J7UmfDbcmWxG4/Y1NxDFb2eo4k0ufK0avQmvL7e6wAyEhxUB6SaeYuc1cWAv
pxMhLCjfMbbarHRq/B1hwAoSUu6rmSM23Hw+8TEo5Nk51aQ03Lz0PJltI+ud
CoZ6fhlujimJWzLBW5wrU80YqkBKppVMUl6qo1/tvf+wO7u3l6GbwNB31deE
Y2A55SIH8xoEtumhM3/MDFQ895Cf6OZdpn0Pr5RTtwx9rvyFJ3Ov9h2Nqqo2
qMEB+Ifgdq8XcDD5F+RpkDlv/2fwL2gOFRd+T47TR/VYRP9p0yOzcq9hhGjG
sDEYwv9WjhL/mffK4XXQCgskLQilTDp/5DmVo0cg3zbzNrL6gyDwo1fdv1Zs
hyKP4lJ3bkebx22b8HueVd1asg2nnn7kJR8w0bXW+3BCkydtLcyYa2uVDjE7
2YRUCCOecCPvgWSvl7MJQUd4ZaeoQWAvtTfV/lsCM1dR307devpO2MrMGRpW
NLiXqA4Tb09d9Ixn9jgVO9v4czZEkLWJYYrLl1yt+PGnk46s7cd05mYMm18N
+c8W9gmlCbSLIDiMdRG6K+jPcKnfLNQ/JwF6HjW8e94rjXPT77CZe++y4boS
qhCB8lvLQbryGXO5SQ/3po5iGM434g7GVtldJQceVXec3Xh6fSnd9XW5FSQv
uVHiwjX2xvbFP4ULZ2d98GAr6quNEzA/ZyVb2uDD0th7kVOf8NbIb9iylCtc
54xsU9cpVCEisf5Qn7wWIBSsicVSbpNXPPC3LD4h1W0V0HJNJ6ZbzZUvrFTR
rtrtyk+mx7MBkL4L6koCCOM+CMMqV2lpwhNnXOgL+ZkilmGaavik1nG0ixeA
A4I3pM9uVZSErhmn333cwvcNSCKDCQJ0fxRREQby5c6djmrqkCe+1Vs4cLb6
M+tRAMODVDepQuXLKtr7KacS8cWSHnj9BV1fjmEFQh0VhOp4h4pt/KxYYxla
UHJkbIOlHVBimDDerAwbgWeh0oBLzyIJumpd5JDkJNojfK0SUo3lJz/Es8hX
xGC3oCgpVnlXDXUWtJqKaLr0sNQPgaySLT5Ou352cqmOlJeGp79QqFYsisS7
AUL6MRjwm/S+N6smfwxp71p5Z2aowEDw5IwNyVD6NrYA9rIva8IMDixibzZP
uPoOuwVQ5TaM/es3A7PCFX+LtEmDLIYPMMcCeD9Of3BROlaN3ZVgyRYUUYXK
P2DUzF6kAIVOXMALT8Pl63QbNI7L0hahbheMLnPPYC4VJYViTsg53K5myUqH
tUbz9qh+0RdW7VCqRaNA+Pwx/+QrM31TDUBFqTtpHa80x1MrvRLyex/t3oHi
oUSvzdfs2olE3uP+1TePD7bz0RaRQn7ogEO+/yRYrfELU+HuAAUmajyItBK0
pqEziALpFNoXGN2R8uOA5CwZISE+Dwo8cC4AlzsS2Ix7bmohYZN9o6yhdZHY
rG/ul0yH8C3CzmYkQYs437S0t1oTnaJhBId9sRTEJEhDUmm0m0/X4F/WjiPL
ArREIW7Tk4+az6ZXikgC/42gmTDc4FjR2jJZHQ484gAI99o28/AZm/lND6oY
woklKg1FDNdIWeoaXm21ncV3Xqy7bgn2A5yjGbncuvI6sBNA9vSJ52NDLHS2
cZAvrKDuKa0b/tRrOvwhQMmHH8PgIcITknmTYSaLQuLv98lH8mCcU5G9HIjy
Lq58wI9jTxdI4jP0Asc1v+NCiAq84iy32hPLjrM4llL3eArwDivgeAA5llgI
ehP5LbXDLDZOOhl8HUW/X5QP8G3/Y8IL8sKg0h7we9/U9xpmeod8KICVtwZ+
HOt9r21C8wsukxRhkzAJT4riyGBBArEowDd2OFxEHD8rkGVRIh/DAZCgaLiA
kM87dQdtnRroFbGpdaNLSJivq3Jn7XP9CUTdGdoNBgZbaC0LBBkpW6aPPZCk
OBeedZMdhhHh4QxEhlX8fXMRXEUWrkYF8iUg9Tg7tIDiCc9aJ/t2ZtNsWxaG
LRwaR51RhVDUXHqwQLWF7pLOVjFk4UhlRPZARzCsdVyuhPlPPyg8JOwi8evb
Qd3dT6t3JMFo/XcmYD2rEM5MZgSLiHM8OHCwmLwawYKlDCZnPJ2RXmVx34Nf
gslwEURJ+sjcN4PdWl7w4WPi8MxLu5K6NIAe8Il4KWX9lfTwe0CE8EXH5Wfw
er26sQihMkgtWpjn2F2f/n8k/TVMdihSTGjdtWzg9OvQi45A24QdhKdT/Y1/
3VD8KgAukGZfnjI17PxOeAjxlyifzRulCmMLA0W8+/W9m8aC04QXtkUN+I5v
tWsWjCUO2Su/NaTzWvdZtSddmcS7kh2VhHIWJC8lEDdWj+N1jWfT4Jt/fKlL
dVEDUVanSPIg4rY/6Dd6snpc1g1RoM4DI0S14sFza7g/qByCaPfa5KBm9dyN
yH9zDFaMTa6zzv9KSu1Pu0XgCzFpMzaM6JlrTcisnFzubOhJpwJccZ/AN89O
qTJcZJgjR0WVzaCb8PcgfU4ffJV5xEbH0gZ71tfvKxfMUxflg0zs+3NuaSp8
1YuPWa0RRVADl5/YrHv3uVcrMXd44Hb97NkhnZiv1r+ERrQFu7/Hv+jraCJu
CdE3sQy/dNbHfFQIW1ULWkaptzna4JfuFX53nRvKF4qHV2S1uMo3bf3ubgCq
OOwtLlKIVaT/CQKo2ZNm6pnSbaRkbgcd3DcSuVqgvJuEHWGkYWL+gmxNvb/G
YzQKZwRNIv3YTBA95MyWtW02Q0+kpVifkRBRPDj4lZWKGqbP0jEAGZAYMQ+C
T4rvEdDlh/EFz9ICF1uD5N4W2TbnmZ7yObS1AtNV6pXdpEFCJbTe5mbS/bVH
xm2b+h4lTffNVrpEZZdGWsLRFTXoVvZ/gZzYyVRZ2cMkxT5mmjr8hnUvw77r
y5iOtsFBBxMY4L1iUoCXDTWrOR6hnQMs5o20m+nVSGUupYpdZZsJkhgou+ve
pHn8/osLe+yEaNsihG7auHYIAyVlNEKJFJ4si6NTuWfO9Apd3DsuXlKX7DeQ
BWMYleGpk8uf4PnFxfG9rcpCOaY/WJLxykGxXN5pEXJCl9b1TA5dJN6rcg+X
SglOCn6dYmintiVmefgAb6Imqok033SWcbN3IdEzJE0/6fdjYNNqeqr9SSes
Sn1TEszDsguEYdnKLPlSiP6CVkZKMmkIH3Ck9NT69WWIVeq2SBHLNAOyFUBf
H1tLA3hBBN6U2wSrJZcOsQ40rLVonWpATcOoIR2QmxDKo/SKhMPTAh5lE14n
jYgO0KmmczSuvFe+u9q5c0NJDujhKKzsaHh4HFTPm3XNrsOW12WG2o4E1ci1
H+lP2uhMy5AKpNgFnuqSdNth6XDxDV0NyDWskJrAI2hakQXUTFCAbkUzqT4/
4ao7OdOFZ3ex47aU4c6oknT2caYhwi9SZU1jZNq1TRVL8oGxQKtKQ0nq4MIB
SRnsuU7qVYAcZvfEAsbVIIMiv7sL6DvLSEdxIwEEokgPUjm68crqHaWxxDt7
9iAQruuFXvMCmKdtgjQZ7MZIuxAQhemLEKINAwqykjMm9fO5Cpi/CZ86OxK8
lu6JR2oeYocAK7nX72G2iz5Ug2qAb1NSi5WdzPJi5LnRhMyyTA1JqB/guCwO
CfAQFlzIINyem4hHuR+jk2GiZn8W6DosLiGEWCz8bQ25rAx3DMf+fZ3Mr2En
xKMe+eIPnkNLk/mm/E5vv23D2r+4OxS9u1CSTeOEv+aMUdizdqZ0EYZpYHH/
JOlSAZphETnm1qZZhgTmQr1UmDlWi5CVHXdWVBUxvLg4jZSfdXHjmq/ivPJc
j1qDVDZmSHug8K+Mgb8G/Cue1w8YWrjt96B9MI27El2ETaN9C9qnbu4KYCyK
jiuaLx4l0GxeiBkPoLzDN2ognHwyzrnrIdby5L3glHUgyWXCqsl2Wh6jvlQx
7/CREkTgqssNM2rq7DUuUPhqe2yNBZxfwZtK73UCtXdgiDoZC2kGWqg5ydVz
FZEW+2N331aIhDDpp0yGHVu6QN8wlPCwnl2cKWW0axvgzGCGAqTl6lwCU/5S
Y+0kbaO5CaAwFIhoKTxwN7JsUxLyJ+9dmzcKuozmBLF8QVIJOgIqmuHABwcL
MwV0H+TbNo8U5NwWlQqdwKeAXuEuCrCVLNePKQi1H9hH4fSJQzI0hFGLD97N
4pb66L5QdxGouk05SMxYZvi87oYljtHeKH05D7htx8VH0kcVUluQOVDnMxUb
Z782XHgM1v+jyWTmQW3vvfAmsBzFuc3MUGeKN0KvarGNR0Mbnnw76q2hCsMO
5KPhS9KorU5/68kuyPVayzeZCX/b9aXgBgznHE4XxkrebOqsRky6iAS7txMy
bwjbwoAA3+P0b/Z/bI5cnoNcFZbxIjCupfulB1ujUK47/z7SqDpRfi3tp/hm
3fk7H+p3+JKR8/mMG/1hviFhjOxuAtmK0DXadyf2+53BT/vU6cEXggilLDQ0
q8+KleMMdpmJiqKEwHGgKgePmUqniAg4pBuRuJB4BytEiDDI8qEm4FEKPCNg
/uMWjhAP2eLGbKis573PEnIKyQBvMO3JmDcUuYfntb0P8avXhscOBsAZ0pRi
HuTSnXNEXrNwjxpo2SHGOq5OH5pGXUhQs5Mb3A6lFWyWyXjGtdYeBRu+Fr25
9wpfaYOj6edUILQAUB95LBzViO9zLpRC6qWp3jP0RaYOgSIs20evJa27KVzm
tKl43X5JbhNZ/5fCosFrf+mZTP70K/TCZ5Peo1jN988uuT7KtwxGLDVuhSvi
2d0Aheu3SzlhJboRCJltTcV1FBx1bqZLfyhMt2ZfFQDVDbse02e8q2jofATb
wiVsFN/zNPGr0dux4EZvJkZw4RW3jGJX00PqCvPAn92kF0tziwFvwYRwcWms
8jibYqaTTAsezF4XiBw+urHfEvuEB2xM52RJwEv7fWfB7oZ78NbrnS1FrCoz
LzTp7I0VIWa7TzdmgxvzQD6xnYu/yQKrkTyb0zDtL6XJbAMiRwqXyOItDq+o
tGacA98Q+b9d7TrL9ToWfhijlB1zivuikI1W6nqFzovlx0T3mUWp/gsYGytc
kmxRIduLUbpBy2DhsgAymMByuFRQj0ShveWphdITncbYnUsWoaqznHw7bd9O
3w/I+bqjv3poHtPL1znRnIv5/Vv7PwqIGdyUwgz3uGVZ854IImRlWYIYp+S+
FuKhWnJg34tVSu9x6WuGfpKK2KnbcudrGGXe9tKBVNudIn+JkTU8Y4NCtgqW
cBpMCNsXIoogoHd90wBvG/OGtGGpZiTP528mnTnECPNu3pTLDs+1yTwgMCM2
fwyf1Ht9N+kw9eXF2KDvleuDnndiCAkdydtPBqwVPdxJES3TC+MVykighAZG
0tY44ULdtpATQCIV3zBcygGNpBVqpup/nr7ELoa01SLz9tD/3GbwrJRbbZAd
yJnsbvd+5nPIQFMvIF4AwE56DmxJc3h1oMwARo6445xyxKLlBLPTstFJYiQ3
DWp8SrN4c5HCyS5Ky/IzrmTymtbjPX4vJE2KqUAwD2HU8DV4kTOjusC3QrBb
9u8/hAO+8/4e3MHUcweBhTKE/0mWIpm/e7q/prdMkIwFpHSOEXyzUSfIQ0TU
iOIOgakQdOtKKLs7ati9HxovOkuD72MnVtjlWkCQDW0cRia+nZFKEdteJSnH
Zv7KrfUf/XqPlPT9sAr7DMyUYBY19zCWZBHk2m8u/a2y/9U5efMRxl6kTVZd
JT8A5MU6SVbBrxufe2RTzPs2obvbd4vTmv6Gv0eEUSZmOglLFlGYWWW2phDC
TJGRND8Me5UGfovnPXF9Y4rAK43vj9cGOJ2bmhymG33zJ5sMbtkESBTAMOHo
lTwXcTuH0o0PJpxtqHWpXB6WA1eW3hhhlzaTDZ8Q8FcL028w9tMZ+3BY/qZ4
S4LfJtS3kow4GwZNBG6/+buSkVBfXrriP45IoZqziKOUy9pnU8DPLq3t9/T2
x8JlwsohsF8OFePg7nl0TXrt+HL90HPrsC3DKDgfZOOo3H/ZbVWrUZE7ales
HJY7khxLJ2wp5crHym/tatMjfG6+4Q6DW/usATNE1yVjMDlA04HrOrRq9dT6
0M6aaSQhoUUOQZEZ7zhNL5GbI8UYeXE69JgcVGbHCj+np881WL5YUQqmg3U6
h4Z63LB9psuzLRfKON6jg76cr7fLpBxD5Vm5PqHuQBut0MQj0mu14At/kHHj
4mCaELFAMQEsU8kDaAqh3ggRAoQHhW3vOL/ikRvHY3hMyHR8FCeb6nQ8wfX1
SwlKH2vfxs19cNqgoTxNsrlnXNNdmGCD2zUYT7lDmhPyI//xnj0YV/XfzO1+
uZrn+yFUd3OoNRHNOW0TdEz/A7DVZXqDRcdbIsmvApWp9n7kMRkSna7jZkvN
0diavJezEaUGZhWwvH/1T/qE7AjKLF5ZS2v/dT+FlKgUHjrIU5uiOqPoQ3dA
5n31fFOE0KeurOOBdTjhR5ohDR8MSRV/ELH1Hb6NrrE3gSSSRA1/0M6gc7BD
w4uK86PlO5XXdEvMhj5fzpdUxPQ0UDStVChofIAPXd6YpvHZoNx+1+si3MlU
CScgQJ2fyYWKbUK2o0eMw0hLQnrbGVu7iP87Dd5anFKE8yhnQhHaVHm5hHly
2CZdyZ+1RST9092gbG4xiWt+CvXiOHHjGRhCbJe7t7gS93FoqEzse5D5KEOy
xwwasEgd1MkJEBjsSzJ3Cao4yhrSX5WFs+aAWpnTBD45RByziXm/+ezS8dY1
341Y8WROuPDzB/W+maitwaDKrzy5mltvtv6EKm7t3XpXUZuZ7rUZG8gmdps4
vP8JqPtB/KheRB0ugXzKV8w+/UY0CjqNem9g4r+S//0sO3UAqtc8TyVKt3ny
6dAPkKoRImSN4ATVv+lZeTauEJAit0Rm3L57xIO5080OfknnHrlBQ5jwvOdL
pXH9gTzgp1fP43yrXvzsDKgPwYocXL8PDypQJ9lS3nfxlijsdtKGMH1i9xC+
4qEj/MJZJhjabKepDrD3aox4dbkTdds/EmOGhs13TOu1GqAN5DUIvsuGcRA9
4ZwsCCeAxuSZgEatLFJ0p+ENjS/EexDIYdxDFlT9EcJzsHbNSRtjeFAC3asg
gecKFiLKy+66Q8CMvICh7/JvCsyHi/jgFqFK4V73YsRhWX4Exgs/htJwlDDn
n7ooDYSdmH23/ja3zUyQkjiOj4jLq62P5ck67yS6/kA6ZxSa/sf6e+bAD+gp
Saj0Eb5YkZnnOrVKKmjq1uvK5KMjoyIOB8fdo3L7txvx8Ong7mYovZ0i3lhi
UT07XSslaiXtiwtQQhEBR9m+7OLZhNYroP1vtpkaA7s8WU5EetxWaUQ51R+r
VdN5gCnEhrsI2eSJjpncDt1sfyhhnaG3E58N0HEsWoQ94luVgsKeMsIjenFO
OQd1PUmR74k9FYIHQgTpNfzoS5flEWYN52HQVz2wTNqLirPVcuPE1idyoQDK
s84Wf5nQGKfMGZ829aavob5Fy06hdAiS37Ck+q4pqJ9VcEpEfCq6Ih4Pr5Js
IiMgAYJSmmxM9EVgrVvWQNtKdmZZ4g/PxKE0avcRq945cpIPxmpingkmJ4Go
mEgZgZygQ5NDeC6vcEZ+ba0JcHKKcdg0S1JkBaamQBp8bShbJgo159tWtAyB
Qu8IyThnBPiKvZLwFtLHsL8OgL7BwswVei23Yz20zIjWu+lQAYz3dCsrX7cP
xElR30N9/UQiiUmmcpYfPWrSwSr2sDZR8dBMlBVXPqjXJNPfOaZ4+oIdlIlH
R4gwNCdqSEaaPtQYSJrW6d8/YwyWSODOjIqZK1ispkwmanvPmLIqSx8Y3xBQ
VRwWxWf8FhtFqdXGv+QYH1RQoufpsdo3lhWaV/avRkOMndAeYExIgrcxttL/
Pyx43eMGFowKzdH+3Rngf+py/uODg2CBR6NtcWAnr76AdRVOnfVv26EubH8L
QC2VRZ1doWrpXZk8ajQYYuh8oyUiSAtcrl4IgIdKj6qM2SMsOVZYnZYO2LEX
IE3oJIYP9eqw15TxAyNYTS02IFTehbli/+c/XRTh+wDdPr5NtxGxnku8b/um
vWtshK7Mcu2dBK4TXxBlRWFXuFGDB/G1bsonBQHnOqH89U1fCBLKL8ocgtb9
+8G4G9oNyA1VBt/OGfsKpFYgxnBfL01Q13wC4kfkPO/3toddjRWvuHGhBc6K
Ko2wWQ+RClKkpN//c+10/rHFNXYXXj48gBQGFAd4z5o7A7FVdQ10Dvu+yHOu
cPvXSCvTirgE4+c+qjszZ7mqSERSClEJ36IXtxZniyn4XCaesZoLeAtRczAI
Kamx0/kFc9ZCMi51MtHlBRdgH4n4wOBbl3HEcF+HUqCTQcb9HCQ2E0R/+hOP
OZRS0AcIKpR8IydPaefQbGFuWV1BPgydPBIZD4iK6WPd0SzQ3c+3xx7A8CBA
vSflDuwWqRNwHmLI5HQy2oKdZGYgLM7Kj+jj1EBfbK8yxMHJp+S/rDwQfPVk
SYMxsWg2r2xPcy9JXqFCKWJ8OyJzlcxSAbztSOiaJ1oychUvhSXwM0bjkxs0
3GU4m7XWKMkWzH5ehyDiuXm6E1skOjuw0woLK0L3kJRXpOfQpf5JW1ZqXDNi
2jEJWcRjj1MqBniQNUQrzLtcHj1/rier3FH7rxKq1OGFh3dK0h/hqY4MU6e2
8WPLfR+idkqjZt5Nn3w9EPoI1vQ7Wr/tBz8p85TmaG10WamcOyfRdFyCYr57
IQ12mEQmpnRUsPRpEPJlrYXe098lobd1J2J5xMC8PSKG8/CUM6YLZAmE0LJ2
SA6DUbWTeCA0RGP41kgd6iyoNcAg2ere+gycKKG30LDFvSgwkhx3qtOfQXxc
FEJ6AGcjmRLgkNR550m8vWKbeh9uF0cX7KMViUYO/DrN2okfYZAfvy7NHy91
qzXBYpSvVdLhZDwLUcKs3Rtvo9FKqO5R7qF6AVk4j5eWMpoFjfLcUcG7JEqs
n73i6NREJkck0kMb7/uCJBTG1nYi7GLvT/1sj+4wWINYN/s0/qFqcUKWmby5
MTxuuzvouHry2eoETPcnJMH1F7F2McMh1pKICVvRc+rFESckp1eO1Rq+u0S+
WFaLDxRDUarA8Qa5nGM6HCmTlHYjzYqie6M6v3KvTX+zdmiauSpxsloL7qre
wso0wHZ8Q2uGQxm0tASZdbi2C+dVuC2BH/ysHHCu8SrIMvkpKMZmrKZHzN3T
HYsQey1qRHXT0oTPlfaVLA3jE4ShI7CwkyHED+N91bFs5lWw8r+nqGMIG2n5
SgmWpOLGdusYRKFgRAfeOEEuCvNWAjFrXNeXO0vzXriK7JmIryQ+GxwuevcO
LRsfk5N7iSVFiDxmXHqrxRk73SYDmHbZ1COzBL2amweI6qOIVp/hG2T/gM+J
s+ulHJwzX3A6PPCNyX+9zHg+SBLZa7xjCgc43s1OOEax2bHAtqsE9MkOaAoR
vd1M5hG3tQ9Z/tE1QQqSYvEeCHbPGuqdKEGzMz0hsVwQMz87sOPFzEpth+F3
gdI/LEvvUlhNJB44dsp8W3iiMgkZy1TYIJbNf0ZOlOCoH5QlfxZcog9E9zHS
xvC2Fm++V/VKrxoSO7VcgJKi4Pxy5YYCOj3nnJ9lVkrHrlIaQAsnkFI9gp8o
7rSm6V02Wh3HvSESv+ywTTC/nfmViIpwvNJ/1aFzBiZ1TeQCSTO0fUXzCuq/
Vpq7tG1d3qARxrB/m7v7jfIa7dKKBXUuIszEBF0bPs1RGw6xjFi2Va+wqLw8
iJzd6UQhhmlKozmcOjfYzxHNQqJ6ZLz8KqqIRcYeqjfvGx/x/AXKHNNaxSZG
xG/OwzwgusFyIn/8DygHCui9ME1SoauPU/0ge5QyzmfnUjyyNEfNn6Tu8DZK
NyU4a8rqiOL74XWeCkTWJDcD5Fo37x4ODdWAQ4oLXA+sQLEX+HuOpXAqhGTH
pJgPwr1yp/0Ht9zpIWWa/1GzDkP5mD4GCDfYNhmypAnN5MvAPf3hDfP3dWd7
Cpf7B/iwC+xoSU+kJk4Zs7E2IUv0+k+MhyWsxwG0YmzBnMgbAHPk5LDd2lR5
2lOAAlMZKEJ4q8Tx4ys/b4mIdIw5WsNKfVFfDacOsqlgwUJGgEnapBW5dcwQ
FJgOpQ1P19p4Ds+nvHUfYSQ+q0m6+UcsWfyxogPkTK/DyHzkN/irnrc2Bc9T
C6ahAfq4QkEEpXRcoMf6nC0G3Upbe6i1cw+BeE4/mVIzrktbujNfYJMJzoVz
EZeCgguG3lZgF1ppiCQ+MX+BHQW+RXmHWlMYBxJzVflxz/3OGOH6Vs18gjjh
lDPZToHnUqpC9kMnFc15bedhj4fNxebFVIMjquQ8Pi6VuiTEEl4ff1iKZ8I8
tRFubF4rejQ62B4RA9mC3VziRSwnOe4b4brV2kHP/02Pyd2Gh2OLZsej04Io
1mEhDLypCsIEeCfvzgiMiXgf/i8gcbOmskD7TcStcmEOwZjpYIJe0sY+FLEt
3wDbZfibbqKhCD9zACGJTSbNdTvMa0kDZnjSS2w/lhZIO8jNJ6QJ3lESJGHE
V9xooYWUcW1wKedd/BLjoR0SzeNbP9fsXxZ3egv/dCBd77dZ/Hw8CX3cFym4
9py/zalaHqJ4WWJ1Ni9YiWo7Z+ZTzf8dzVKpnRYrc2yKlRiL0L+X7DqOaOKc
jbCBP9sM2zom3LY+9cEg8Tyinb8NQxGwQzJsm3qqIU2GTgt1ZqyavtqpgHpc
VpMxTt8aMiP2C21u4zpe4VP5p093vJbtQIED0Uoj6HauMMFrf8c8wUiddlPA
16y47ixBxF5BshYc9mEZ4FLVICTxa1J7rEmKryBZWXo8rcSYHy84KH/oCrWD
aVGi+mrz8QhVfXJJ7OPC603kWeYBpOmJalslX55Cmf964/Lfaxpq8qMEmV/9
eLby2TOOC7haoLikFKj112EzZHJ50DBadj0E7hHEQK/pOVu7QFDwCHbsQ1KS
7/RpBOoLrapKbEqR8WGvBDKlxpB5k3HtoY3fqRGqg3lQwC1S6WyPwL02Ryss
nlWBD1YRenIT5bq0FPq/29LvXklYMQQIbJrw1gmjUqqpDfVhHIjrb3z68JIF
ZtFAEKwQV3qOH7DrliJihNfhvZyoJWfKvbHndjAlRYjtdYSdyTVFxXuvER7j
CJMx49Vk1fugueRWggNalhx39O8E2bwNe9N5+gfDxIeZXseaMZigp0ajald0
9noTNfQUkk/7X7MA14FzGKd5ElTDC8RhxqXlT3FdfBDUfXCYWy+UY+jFOfCp
7B9qNUcx83di+pezrRtkv7pxJyelrXE74WgnS2M3PRv/8+uRCM8iQGQay2ol
+684I6yBRWo1tEeQrzmeXfIPnsoGrwrA51Z9rNej61hjTVkGfa2Fybj/NK6e
SR8V71LNlC8KlU3f1krZUFMJ4uGqerRn9Wzzdf++eZxl/+vVHE1OsP+g9lrC
1VGrZc3KT+DSiqUwYh7WGa79aBMaXNqUAP1rHo64YabgSIErGE2gqkXbVQ3A
Xp8VnadP1ygLkMuEEV42H3P1i/NzwnvfdWmLLFus9oEarg7QaYVFvAm42/wO
bLDIMKLWCxPQEGSMFzA+r5Kbc+JVXjqVd4gVf4YvoxiP5Gc24cpVXTwKQQyt
0bwWv0FT4Ik+Cp581vV4nAZkozBAaUTR3oUz2B/ickN/zWMMJ4rBXzRFrG0n
xT48oXTXRRolI7nIHDZ27nPGYGLXsSdINhhFGVXmcKLXN0mZboln1Bbe+Bot
TJ1evURnBd3tQLcJSaE/35F+vl+wBM7jO/YdK7DpYWNVZAMdIP0JLvLg+uEF
ThwQIMvjAr+HJpm/S0ASNPzat+TvUC95RgMQo4Nt2Q3Q9JMbUORpazIO80k9
KIarf5qW2ckj6S1YKgqb+jj88bi2CMSNANI85GyyeU4yFCHLbFjjuU5/G17E
motBxVj6hz57BNSnpeWffk+XgcwSRfIk/4ay3JIA7OiA62mAErcMFBIH2y5b
xHUfllXb7omzx3J6wP1TAFfko7KYcalolUckBZzlT2ZgMScVfU9vqO2TfdjE
1CLaIc05y0VH7R7wRTFsl7JJOFLoCqCwSAY/5BqMlbXPhJ7xMbjQ4aEiYwnG
LAglU66QrvbbjwlXpgM9aSDk8+i73G2Q71HNtYp0ZFEwcIirYiVLvFa5sTbO
V2IB+vrDy+8ioS0oIFjZLxYZQWtMozmW0gNFZxH+v1v/+C/gSVQLTVER/pji
4lutI2ctxfDdZgYBJKgvPB3038DeS8saebjEOCJCAgFZAbyaKk67MMHG8FsW
920bItT9ISaIztL+nwrylH/NDePkCalMl5Eacxz12BKWVsS2ytD8fXNMVzp3
V6CSqn4izVeHUXL8P0tsCkBVzb+c3vTKa2eZCrM65ZmdMzXbhq35wlFNe8hI
aHDNIUfHrPL56/+bO9zo+gZEhr7CKUztgW8eGn+fzohV10BBLQvvGvXfyBQZ
aIoq3X+7SxIF9ZaXm5ijmRx83RZYVR8TL+C9V2VCNeOOSXk8KD/zj+0btgjy
nsDRH/FpeOMjfWAs704F6yKj+HW5J0Qcab+Ag+88Ag3W6pBjITz2Q1faeW80
xDYTjonELj7Lx3h8yqUuwd1mc8NlR/v8TxMwVaD6mCZBv6w4NGGextZ0YptQ
UH8yOLCkQCTi49sXasXk5mdMQRyTq3KKNfJBkwLGv+quObxpMtlYapAoY+ad
gzAZr8acggnXNlxx3rLGdio4we9X/k6Mp+TuGyYYxfsXxVkN2CfbGAN7sXez
m/VT6/7jQsF09T1xHC5oZF7U0dvRbnonT3SBCTFMuK5QzC2fPLb32dCvPWDR
jMZJ48vZnqniB18ikIJ10dR/6zg1R0FWQ9vG/LBTs4VNnmdrHuZAD5nwKuQN
VVP6l1Kr7fsfcudc0/cIjbu2OR9UC+PgT/it4bshFlRWBVi3qbztihpCoycX
VnPyRsfLn+KvQf+T/QI0iAPkF9BvW50BOSFcRR6LyeAVC16LEBc7GrmerniZ
z+Q7+IQHzG2qAnVZ6z6L+nSuZ0Z7e2+n0zpmn8bLKByWCvM2KXEikTqn1C8C
F8bmVDnRCHXn/uhmEfF2hF5HOkKxNVWH5CIHnhL2FspRq2HyVsj4LrGIOdaH
RWXHGZduGWCi45vdTJKLgdXmISBRJL7OlEJ7u04teBNGdFVNDj5/Pat9eUKa
Sk5c5NaNOvBj1NZBEtn024M97exGyPl9ftdXvhfBkSclwK0RrvKtpuBBkgaR
seBb9MVjyMpbbdT04orBp79Ru52w4HxVgSy3SY8M3p1EbwebHUfTvBxUsV6H
KCkzPtrNeBKUwwMPrzNV8A4nunxI56vZG2LshqBU1MrokfqfMiAR8sbJtPjX
PxsRibYaiw3EKf6ILEptIU8sLGHkaIyL9R0S27FZS76JTnatJrCTN8cbmz1w
OuT1H1VM2038KatEyyAMY+lRgpSUUOETeY4oi5ZnIv0qNxlFIwIrgIrGvK4V
O2w6ckWiHuk6bDcSF64HCvCU16lHBvuIEusrQ7CxanI+JgeltzclgJ6JLnaO
0+FVXLo5uWy7CCKTSQOxxDXUGGWZ3g2Z94tW6iLovzFV7mUtBFtcEaFdPPBd
gAB5xKuBPqlOHWbBgAQPYFbP0ue00G0rJX/hpW8reJn9t53kqbuusK1d3E1T
Z+1tqxx4BbYQ6jtDDt0/aJSope0UpivR6E/RA8p79eFWg23a3j1g8AOFLPUt
dTDvlOAM9aLFSyPMqrpbhvNfwl2UV5NlbDNVbjFJMiAAdz7cSnTZ7ujBImKQ
TCtT0APRzdI0nAKf60/MHlD/xG6gViKNxvnns31ghM/rSdkhZqJailMgbapU
sxc0bpTl9RfpUf1NosSkGBUbbE1sEYds1nVor4HxNvsugwKymWXylx+Cp9qj
7gndO5BuCi7YJDm+ju1moDiIOqNnw1fMp4ozkiLIBvY0ZTny9b+0sDJ+MBy8
mdpwKixhHeSRn5RPrpthlBDnaX8gWIZ5BdKDaGluLch8FeNGgEELWY05QAEI
x+ueFnR8iV/cAFrrMGQ2zqbIlyaA73p6KIUmQRzk0PCPosCnd+SoRucI3XYB
uJr6+Us/hKZxpKpPVsxOJednV3B8gdzNzD5sgmYU5V6wI5x+8NS/ZZHwMv0C
Ak9Dwv3wCLOX2gkLy1I/JVLi3utrB6H1L6L0X8GQhCvgZR2PlA8bgVf/s3MV
KfGhpe8FVqe7tjqFejBdFL21MrjDYGE4of/e5JgGD5LtKImplJdCKS0MbUKt
+ci5hZmG2R+ru8eVXCm4i4KlGDlej3wJ0VS8l2/k70rBhC/pMMHBMWwYC8P3
bz4bOTO2DTFcuL5kazKiOSA5rY8RRU6L2sReUXn+v/2k+lJ3rd3vKfakMlht
km0OAezAk4WG7wf0GWlgHPj8p4mzODf6rUVcz/uPenJ5bv2f88BF3rs1duS+
9629rSaXco//FIVwnwj06B713lqdLbeTpysRCz7hHhO9Dxuur880QHovvtwq
sJdtJlflwSy9IBeCekcx0GCyEd3GFQg8cAEFIuDeMSsIi8+dsO1lzjW0UMnF
NV/VzAn9Fpsehltlp7Zu0Vd2QWIThXvNEd7Nvv5YrQZEws4YVtQyk3buraXy
un5c+J+e9EEfCrLQFdAyh9VWl8ALZ8Bbs1yi6vc4eWmE0kAldHa4FgLfAUap
ZrY0aPeYGZMv0kCcyn9gvVZGXNUh+l/lAsORXW6v9Yy4PeJoqBGdNlEOLG4S
3drztkiXkRCM653slmtmYwU1O6hbzmEDIZVoIy8+NeDguW4ctcn0pSQqioHT
8pvbhWIVraHyQWWa8zbwvw1G2+Svn7CDZwPuUtPFzJpvQYN5O2VxRLl35MFY
mYlmzywabdcv3vPwqr+0qdgT38oWGdpWtd9TPbOIXZOSPiGn5iZ/xNVPBxNp
MHyxc3yHW1hpCgovUDp/+033t0bsMCIy7HttXR+TSqm6CLjvGzAt0GgZgvbq
jIeH25AxtlgAIMxYaTqrEmNmEXDvbnuTotKoCa6d2+/FuKKtVcN+18f0YCZ8
rQyJzCqw4LPgcn18FIKjJs1oo9q54CqdSuftNS6NQM1UZrg2ysuj+mOHtfeg
54qCKe3bFD7r03bZAeR8J/HQlV/2dT+NDtbV+xB6KZJzJ/VNPV6+mNKt97HC
xwClxox2q5NhDxCOeDsCSeifvSyGma9F02lGGQPy6VN3bYltXLIg7OQHCfmT
zWqaAErOBGdR4Ig0rcuFl1uFdTZbD80Za7YESYE2bwV/Y/i7ezXy/5dnNrpI
cQsXvWluaRJWimXTcF4rlh2WHMSlD1HDEkIdSWktVwQR9TG3E9EnoislMJX8
Zq0GuNvbNTP0mRqumONei2/y+6XREDgt/WqYcGImzVbg9m3mzuqS8SLLRD3P
ppS/cxnmvdC737zW1Xs5VKpESU8oNzsCC239s5Kzp8MMQyNI0k9YlRJlMiGz
j9bVrvvN9UwUn/Piqy8G8jfibuzEG2gLsQbnDZr0TyJk3YjnL1wBzuwHvr/z
oO3gnXizPpGJxbFOnXyUdPAVFgIsQw7ud0r0icxTeaFX+e2fCXEch53YW/af
X/SU7CVTX2Q91hAc6PxgkCfaJhKrk4sTUen7TcSEaVUmc19IGa4He+OjVQ1O
zqhSV3gF2l7JcIQilFJTa12cxaDGLB/mX9vYYZPqXTRR5LGXj0O+yqT2AGKX
rTztvlAmyAzJh0coEbvfoUlSxFMNx+pZtKP3ObOyy09Jt+O4+nlyjNjHqsHE
Odkfk4D2DVCkRWuLp9zr0M4afOtp6sHEWvNSwrCvpDWopSoUkEU3iCx0dM8O
2MDMR4ruMEwvEsw8rtV1+IlTWTeVflHC0BxZyy3IIeKZIkhiRSV1/Ag24WHA
RrO7rZTen3eiwERplNrDxApoiLGh7GchPgVurau3e5IPrYco567OPrSPY34/
6pIXjxZvQMVUNSOBG5+DW/sAgKWS5ao1+rPZcp15M/6RsWjl7UrLiS8yAqPF
wQZ7mCfVn54fsAj7AZV15rHJZrsio4QTuyR+5Z1HdpyuPmLvFWuhLHZebu2x
EpQKKQNdjVWMBI9G0uVpz5RTTpZbDqbXgYyI0+tgFjTYfGEBjABiJOBHexNP
vlyr0bZqXOpy/TeE1IAoTF/a6ZUF4yhFZdRvFNZEtI7mdxUbGfFAaU0tXGjI
fBf0xPIBFjjit6WA6Hb7H+NiSK0tjtvslP8tioXa7wDx194IxESITQaCPsOf
Fn6D/cPHh3/OYxKxt8bn/bCNz7c22hhBkj2JLWg8ONdeLJtUzrPDPeeCPjWE
2ruywr85CAbFTx38HcXFp+n8EoLTSQGe9LI91qEwuiUsxAkoPyf5tvYP0c3E
ueHKb++SCW24Q0Yr3noDohFDz1olQJB7WfHsMN8T4crw5VR6aqXrIJ4xSloT
zYRbpCmemw8l4elArK/DZqhzfK0gfN4Isg80EAROK6LiWqlZx4Jte/MX+01C
e70PRZrtf2eengRIzRB99fPk3PqhuFz0c8zxAYVGBKnN2LkLGyX1a4mlziWh
Q4OlLmuXTttAe4UD9F/AGHGN4ZbLwgxBtO8fGbmJvJSXYsKF3XeKdWGB30gq
Cr9eIhMYeFgPmFc9JVcopdFc3mEoImlppsBBV/q9ubsv+nk8ttwyd0OfTEvZ
mOxu1itZpiVlfsfLz/BHdsYJhPiBnYbYKNfjqQALe+d0/2yDeTICn6cKDYQ6
DSeqkUdpWpCif1gaRQRvLvds3ZOmpbbdt040aUtOOf2YTVFwPypC+dWk/TEd
GRyLNMbFOHwt2Fuh7Hsd5z9zR84cAty/fJDzEkFUtnreMn2ChgGnPa5O5GUz
55decAFPsug4mO7gOO4j/ig+LpyX693o279Om5Qj1hR1BzDS6vivS9L0+/pB
cW5PUoSEH7oJkJanyrKx9Wi5JePS1UI+2MA71lqz/Cpolb75PCF2wU+auXMM
v9P0iVQdqs6U2Ajo5+GdjfB+CVcDSIYRz6KBr3csGpvO49liehrTfdLESpqZ
qg8uQj7x/+3o4ZyChHlxFOlxQXJ/PmGw7qz+zLbr2tfi/FpeI/CdEOYzMK18
nZSXfwnOR4ORJOoBDE64Usa8wQ6q3MqH8enoczrMPTzqb0I06LfMEn5hBC9N
3AhxjF8OrsOq9J45hd394vu4ennIe61ctaKglnRP8ARmpNSLQmiQZZbf7v9d
e3sYrUPKe4Im6c5YIP/Kq4S17eIFG6Yys2Nlu0EjiArHDeE3YT1D9kLT3PIr
676tPA2/u1nhiFjwNhwvzTT1rgBUZmvhlfKFLE4QOnQ83grsde+BRCuQL7ms
qjmcftNyEu4LtLNi4K9HiFbNkwR0ojp+xMP3TQQz6EOhiG9yhdBA9n6OzRbn
4qiu/dVWWwX7WEosJgHmbbRpigWiEGdPlIfpOTUFXGjZEFc3DnDI31wfT5ud
aka+HTMiSVXkRriE3c5Mup/d3onaxLtR5jMLBU7KVvleL+C6q8wjCJMcAhXz
acVYjnvw9yaAFYiP4GUIqdvgFuxMN0T48MnygaFmUYF1STesshX+/p6Na9pN
UwhqOv0/HTuKRDjFhv8s4Orq3OpklWKguicAFr5RaAFDzye5TWtLQ3fgqhV9
FyMBqLdM3n568fBrTndfNgS0XHMloc2bKQIW5Pid5/PXqC7kqSeVBtrHNkZ2
DhbSNNS6rgFwTXVoWbMTXIUUH67tYtkA64eUmN7Cdlr2Jive/G/9ZMICg2X1
FXw2CaDpYRqHZKfrjHk0PB+fMoyCSslcsNZCCKPJerdMr6HyafSpv24ntanX
2LrM2OH4lHoiesWB/iY+SJ9S3G1ngq0CEZMdr60mE6I1uPU78svUFPYuomXu
a/EKjmJuoInLd2ZL23srEP8oBHZ7IMHzExeMOX7Ue5A3A9bzxSVLJwalN+UY
7S+GPf5ssqzv/EDYsPMCLvRh4ADEA/ssTlncOf4e5pTaM1Nt/6zTZ5IV9HOq
UR6rhpcYo0WeRycAE3Xfw2SNuhbYFk+Ugt2yF8tgo0itb6lAKhx4R1KmdhEG
Jxa7ybU4jtsFPi7T/Vav3VGUakSLalW4xRMl67hlUETAC7ah3zRvS45/K7x5
/29KIn8N1gCx/9V7MIs23afHskGcUmvkZt8yudOPGfz3r/dXzjECdWEyc/Y2
ejTneccnrN1Y/YAOX5J3JavvUX9GgmOz/4FU3myDFsWiwGxVvzaivO6AywdY
kFES792209v8zo6+IL9QQP+nejHqKs+EQLvFwvAfVYaDAsu8g3GP1Nug0k8y
kLgdLLSy4FJl3X0uVJaOqCRgDJnArv+RhVZykhlO7HAr1nt/EA855xSPz9Jg
u04mXgHP3qRECKH7QVwVzNJ8PVggwZmWf/mzGw9rU6B+WBPCwopb+BI5nePA
RRj+JyzdcqfG58wfCC9h6hfumwkfBR08y3cohB9GimMzGKwmBP5iLC3Ia7gv
nqMNM4MUYieKgcnVipPcns4uAG2pnhD3w+/cSE5abops1ilHpeTlQny3KolM
qElgP+ynZe38121aLXFaLtjKKSmB7qBLsimGPB8ydT3/hQB932Y2D/5bF9M5
rLZZZ9WWJk57bHJwtzOdTPuMjk5h4W5diUIMuZXzPocPEQhed7H8uEZSYxsI
1plvdD7IwBvO6fTvrmow6hMlh0Uncu2iZgpN77WblFSRSX4+kdEBw1Q5n9/4
pSRl8+pCT/dILXfEzOmkumk4J20JKj5omYk46FDRn8IZOD+FrsSMQZCz+VnD
wOicLSKh4PoFIvnQi3YR/BCpatEb7yws5vVQcNrOK4nSpgsaT+H7BgOelds4
LGUWItNWxToB8okuPW+o1BqyXRGynmUVgy15MiyHP6dcBIci+1dw8uQS18zK
pNPSCOeXXSdiNJZHPCz19FuRbfCu+2RHci96nvuE8G15JfI4XGs+rqjHo219
OEtopH5wUSmipThD/QTVFts56kIDCjuZduT/FRDYBUOE5CbC4ZWQ1Woj5HSl
EXCkfpPvbTBUAw0CEdYN1EVU/5R1O5vTSpnYvY/KrGsKHAtLthvEE7vPtN32
yJpAqH0BRmU7KJCV+Vbazo5d91xX7S+xaieJdmr4efT9JYs8icTGKu1yPv3u
R2Bk8PzKdnbm94kTXwo3MHbYaqIC9zhpbIz+Rimv9gb45JD8Dh799qapp4C+
6WYgIvPIWBwH06vs3itrjdfKxDsIXFmh9+gt2BfvKBIsbMbSKIUWNX56oA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "B40jvh7ud/ahkCWXo8CJP0S9JYnc5+J2pwOdONjrEnmjRzb1YpxBEP/gM90XdEQFf8e+9j+GJABVN1VA/EUgHmy986oXHU6n9uJJjaeBsR8h22iSaiy//95eH4kKFakRZgkZDqWp0dX7AUTwRg4vZKk0rom9cx0xsiuc1Ki6fTzxDmmuuNW+yyxk/luKJogixDl7f05H1PhFx3JTfD9y6cRFGovJ+RtyYHOBbLpk0whgtxG+DMVB5ShGXliJgGgQgtS/OcqyiVstP0PFPU96Fxfw8TkMYRV5IKCsgU7H8WOWoE/I+MsHE8XZM3u2ZhlaNbBInXs5EemLEvAX1bJ3Hl8ZbYURbrxUfBRSbq0EBRmvIIF6Xx3/Vp3UEc0f07FBHPzU4YfVMjzLhjQiXwljndwyL4jPci67opTlmr2SDh8HOE8cw9R++PqF3pNxhcSKwJ/RWtQuPILDBI7PXyo61Zknc5oml0BDllhEYwfRxxAnMB6UPLk79P8zc+qH7/oADMZfXuM0Gy9z9SUX2JajYnyzeE/PzFOWLKa6BJj9VWhJNyPkwrF96fNFFXif2fLc+PGIFKRyorjeWEfTfiD1ZDjLZRhx1fQAGvF+ye9X6P0sExjzayjZhM/VhxL5vR7EhdB8xKn6+zPU0bNcOIePTfZw+hYjTFFOsZNiPWSGw8WasWwYtjZ7Hnzb2DJ87PiIg+SYZBMdgy9Oihn7ZHodFI5f9++P2KyWOIXQrw7trA3QlgxuQTIvCPzEe/jSYxHoYMR9cA4rgYm0uZHRAlOZ11KaZzx1NsOsPR64VgHjiyuz+bfSNzE6heqBAyLxBzyP3xyhaELg+6NCwS+cUGAHan8shQ+lm5JTUjIfNJXj+HmyCzaMUTVY8Gx6LPC4blfxI6ARSdyjj/ocmhW77vynNVxeqCkLuFaoZKhKlLnordIgBIAHEjHF2LvvZ6QJHERsJEiZQldsOdJ2edeENb0wahBdO8EZVfzotMz+4sGvwdftoPpoGqbeElyZ7tlInQfH"
`endif