// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SKwUcD7pN4hGqLjQBgg1KgQ9z92D5mLTKCAfrXkq7mjPbfFLVeAlQGrkWIM+
pV7DbN4rJXnUuaq5WSjcxNEertIfGg1T52Bh8Rn6SFfNHTxceoBCW/5kTFt9
2ah2FILA+OYlaXsMRdyzhqaHLtQRfZGxiBsU9MHn/lT5mfsHmtC9JVU5l7K5
q9E05TlDnOQd4t5pDmghRPmsZsXlCOEN+o6QhQjdz0V3l/PWWnCPkiYVYIhm
dtMgh30lSvc4ChoDJWdIENzc/Llz+NEIEWP0N478eBOfFBS/LlWTRx6t+Rer
5bTXn+4K+8VRVe9vzmfmlc0JsBwFqOpyYiE4CWPThg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
k6jctTtInQMRxRflnysrMExqqUuvZ8HflWfvtL4cYFL1Qg1r3SnlZlwj3J2G
nunBiK23NKwxhl4AHWAk+yPN5KvUeSzLk755gDbJnJCxNYXAl627bXpE5jha
rQOPYa8474OWIH47/UE9BiZsTdrXzkHS56mFSmFdjCH/2QTRgdA7s1H88z+F
L8XCbZsrRRlv3hzih3iXFw7GOx0g251WahuNowmomrwwpZCOeC0sfSfgMiX+
r3tdCJOiWKjGdsluYFrtXdMRU1f2qnpun4o6Zr3Q0UU8Qngz/b6rmNzgbFuF
AGYcDBlcnFYhq2rWI/kwRRnFgtMpJkFiFGg6B+PaYQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Pbma+aUvOf6rD+9fKXk90s4te3hHqbtXINCvpVmuwm644HONb6SCV918LbJW
l5YRZ4Opcoc4SJhveR1f8dcaWA+y4veLm2gWCy8EHxJEYE6U3ehNW8ezS7xg
wEvoPYahDM6uEnih560LUzYvn++iwTQOQQGm3ozKR9x3udHDRRzNV6F6Zl17
IaJVNRsgJTUokHdxgJGnviG6I1RVZ4nImPPdanncWKm0YK9tN4UGxrBKl6e5
WwDS90rcFPSvCAY1GEweJA64CQy60Bva/0ZsHZe9FIHu6Mki4hNa2Plx16oH
bN3PjsBcB1brNBEx1WvqszogOYDBxVlFIgKvdx99LA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ggx3Q1wYCbeIz0lxLpyrdLBiYZ/NuTrQNREsf9BYgM7d8kxCw35YCmd7WMvE
p4wnKp1nSKo1+mURSsY2SKu+7MhUhPhIskC0x2MIqS/aDz+niyqqDh1K1G77
8xcznwK8rwxlXVB2NAqfsmVglCrFqjcVl48KU4Jmu4r72E3ahOKwes4Yoewl
Cv7Nz7HE1JT3fUxbLc7hjh/21lmp6swVtdzJULQ0UcnUCoCaYrPxxfgcOVUq
HFafGFaco6Otm+85NWjSu3i0S3IPII4DUiWHzwvI9XRbG9U6WJRZDgl01oMC
gJ+8BbMUezEjJBJKBmWdDwMsgXls1BHSNppwXmz3Ow==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dK6xZcp/Zml/19nlOt6YfU212/O6KmOTCCAswx8coEPYsoTq7YOz93W7XFVh
4u+QhmAoi+hyiEyQUeFdruhjTnqIK3G7Je2Kg50ICa+KKcTf8V+vj3/Og8mf
Q3GpBuv4HoJw2jJoellww0RbXXIuKst+Xw/r4DZRIHJVZaRI/Ec=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
SR7n5gpUQw3kazVoCJ1IcDfidGsb8XWgN3IvirE+uLAdhoy1LzvTT2GGFS5f
SzgxO7ae+LBSMi3X8gNl2/E65Umg8S5A53E7Hm7ipk583jmbbUwiqC4yNLje
1KgRACuXly53AlUdXaWgmGIFtKZf4jnGgV04lHipJAE5Nz1A+CF+Il3ph5ml
zkMK8Sc2Ib00jwpeQWQPolkK//v6c01m8uGbKL3pYNB83spDvM8UmZPP6SgH
swHAQukUfAqjvoAOlj8pHVhGB15J0PML2AzDVWw36BQUC4l0Iba10JSPw++O
cUxsiOJJyGyRCj1I4lBeha4UHWtasR72z00sA9r2ySeZ/aY07JkP+UzL3yeU
Obzp3kVxnnKbYc+J5jztPyD79Uz+Vuw87wPH/1H15ygeaIlQN71kCLiYq9Ga
2a1DFlEXVErKixTd1iBX3aINLgDI8FfQvbl+T7K1rQhJ4XkKMH2kMc/du6Bh
zfLPflPcQD4ixwYV7pH0mz+bY/nk7x+M


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gnRq7avTfdths6Y5vSk5pwIhqXSIu//vusT6jcRn4Cn17RwFtIvojEWm9yn7
m746Oy1ThDyvi2EXNcw7RRPYkSc9uL9cxl8Sz7wH70FfObVEcjKne8gZ0NGS
2e0/qNYR2h5a44YT0DmydUTG5ebcd0ST9u6AdPN+8UFOuHZVH/M=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
k/pYeBEYdMZcqV//tvtMyH3HCf8FnFXMGMaiFGbcg14FigDSnizzZpegwwnz
+nHLTTZ3PFX1ibMU/RdiTP/olcwBUcBCCQI+zmZa3v5mFkHLuaF99nyWKyuh
ccc9Rkn88cH89LrcfjlDIKuhSb+DP90rsKJU+17QcfyPmY/NRQw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9280)
`pragma protect data_block
GzwB9Wbim0OMGbzvhaDnArszyruokDQxKL37hc9XYKJtiDkfW2x8lSLjoM5I
7GUgAPp7qjfvQkmTYZVwOvkHjC+R6u5Kbm7EsGh6mJjoPTzMeJPHYlBfOk75
m7/HUoglUQQynERauTMwTwtoNQroPyitiVSkeiEpq6/BzDZqu/cCg/BSVz+C
vB+hcZvT50qkHNshDrA+SxI2N5alhX3pfmcg64MYKw4qOH4c9IMECHkMj5vn
ZnAgXz7uJfjRsV8ehNmNyi7K9xXmhgAm9R/M7TmhuLgY1mtU70qdUBLibPjJ
BQSs98H2j8JBkX3F+IvB8OYy49AaF2Wb2TbXDabcLIys8D4MM/QfLailzyzl
jIIXm9Ml2N1/Pxa2OryqpV9rR93P5oGClg3tmqGJr5XaW8Xnw/B583j/WFG1
nUdjebVt0raEeYgF7G6qanAfHd+aD6vmLEnTahQai76HO5uO0/lAuIQ3QWcZ
m/sXowa9IpETMrkUMvvEhQu/tZqWp+Ah8DlOSNW4GDLctGxxZn03hDJCrZdd
lyRoXaI91hmYMoJNsX2j6mHWHXH1PgOx1NBJIlumbONH+aR+nCAZeSqfCD7P
7/JgwFnP3IhHbYFLa2RGmLpDkca8s2B87HN7twTFRJscVdkidIvVUbCKuYSK
bhf6i5CiXiNFvdV/KSXq69tHTCXSxX0uBjbBJBiGQdXWGih/blUmAPCaeJhx
eBkJzBsDMsIwiKPFcYEIjIc28OpRHlVx1ipNW9W62B3M0gu0mvMfZD829OUu
QJjq9LOtZoBmqc9vKwCXCa1y/qfFpRS9OD3a+Y8kBBu8qPW1x374+CFVZHUw
ZBa6hRm35XUQnvqVgL+41xJWz4FxzMdBjfTUuWI3MhVt3mpMrzVgQ0QM4M0B
VIOO3LXGnTao7J1cY7Q2LdTktQzj9qCl1gsPjKOucUqEEK5LpDliXsUPzcH7
5fq75Dilg87anZICsEVSwalvv0bJ2DNUC2CIiz2G2/19CmKvopaw+5oeA4/T
yq5w8hGaXABfA1oM401HjIzSuqED+LHh4v9fJEpG/5VD4UWzw4OcdABWTCrm
B/HkJK6Vo7IvPWZhq7MdfpvgOxUFC6kp8EERGk3lzIE/+mCgQOoita5MVcFk
e9mBuraek6736bWYVpjvdMGtq+kkHbtjTuCDRqKljn1AcFrKfmU7cyvQcyQh
vlEqMtPDqSAGcbaoefF+1TA7OYGPIdnraMPPU9nSUA4WQE9XWntEbPHzL011
nzLM2N/L+M+9WavpHFWUxXArC7fX4uzLkkCM1HtdvbQuJIQRvKgw4OtUefCC
LhqqydBtctWwIE7lmkwLXU+68JI//Lh96oq/Az9nFNtHLQHk5l51ll9ayWN1
TZ8EXIzI8ipKg53wyfOnDyfMyELyrT3g7wsAaBLlh+7vii2YU0WSLFU7JzFj
U8KGY8tP0P5PBGZAE0Ck2h2YNIGVDPqtv5RYE2B4R/MfIyxjeK9HSqt7XtZx
7ijiapOujSyS9YUu20fohSa7NeIqWnxoICz7sXeHsAz0yToNiCrVS9n3j3lF
FYNz5b3urH6hiz56BfirPda9KrIS93oEeTAd425OGtENNqOBAi7PMimZKZkM
PCRcCgzcvATtAQyTCXUp4IdhNuE/8bAqAmzf4tg8vsrxlYkNOmf5lPlq8+2Y
nZi2agiS57mBc1fg8H0MduR71g6uDgsIuH/EJiUnb+N4iNP+LdFdrvC4ES0j
A+K73T/FN4sJ1HWRVZaeCnINFQ5lloxg1qpARF4uvfjC0LMeQfpVB95C8gIV
HFAgZLJ4JIK91bJmUfzp/89LC9nwtVM5MVEAbl+Cif+ls15u7cyKfv5dDtCQ
NlPV+gSqFiMKpuRZOC1PV5eHPFYtk8xkEkIuU+hlxe6FeKp9knktqwCm0Vb1
GkAuQBVtj1XIjVB1aO3YUpZjD0naQH3VpI0idCcriNKxQXYZR9bFS0MbD0yh
889VtaSS5CfV9JvOmGxWg1X/b34thu5BA0BYLm/j39xvUzQ/umZYBNdDSc/Z
F4pavOVq7VGlnnhnKJ8kTtLVTYq1sVXIvgwGGKHenlbXy5kJ9tRNUW+G1han
hmAQ/vnvQZl/d2jNxgzvwLDcvpWeeuvp0zjON4BfbDSoaJNPy0bbzIx5XPWs
u1iPQsQ691Uw1iXhqncDIbgzx25oAYc051sfePi8AtsN8+UUeesvq+w/+Y6a
anG7GiEsdqp54jLlH0SN9pwg35JTCJOCr1eKbzkMxLBRDg/uHDeoLN0t0Fdo
sVSrRQ8ZILdB3YXXq2Z2PwLjUFvAjn1zNNk4gjjPkSbI6v8kYLFCDqdGt9Y7
cZqQqyHkIB2D5QPwNUFRymAjrGhTWVI2wWw/6qJbLlOPz5JI/i5h4UHQByHa
yQ0E1IjANBwxgM0EGD9nQALXvfr605A6M+D3PBHPGmB22fiLjYNv1aIblaOe
Jc48vIlEjQUweP4GX/8FrP83ph1Ae6SExVSsFAkng4gXXUT2l5WZ4UzEPHLO
J0DDljhoUT3jQH9GIVaKYy1bj8ygtgERczgumAh1UcLQ4cNCzs/U6tdTWyF+
pFrSWq6xvxUklGrcQBRKNjPeYWwaFSxQATtGyTCG7puw1E1BbzK8p6D53Xtu
gryt8KuGhqMTllSsczwGCARTeJUyG5ckxZHZg1Kk+W/J17BmdROt/02lKVbp
q88W9ubg0R4pHgHWntMdLCMxz+PQ5hKFCH8XwsIg0qcNChsKS+qRVWeB2O1m
qfPArNQpvcxiT+Ze1Gg+/jc3zHSKPlpTVM6ioV6HtcTLom/o78dk+J+k2FEk
IQ6WptLl8Nb4EHgWMuwcY2mUs72g7UM5IxC0LiDpWRMHw3++tEWGE2Mepvh5
TXVWT6h5YGrCUnn2cYt7Jhcxt0zmJFXt5mXkY4vsQh70WGC5E86iNwbJoadf
l4EJc2fBtrBZWY9wTcQis9yXxkFv1WtMB/c12cYVLNL5sRRzwqaBnlBii90A
PyNyU41X11hbrrdLHWcgy9CmPs8/DKvLOdOTqOmT/ci/3RU4FhwDggptQIbT
1rBDi73LVvVtLOlv7evB+gRLHwGFZO9dXSP3VvSuyzFo0zEA9dgbhks5/CLh
ekjlBpJn0x+kVeriQddOS7pvg3W5EbyOKs4or6PsclpPTPqjPg7KAuJ4EvoS
wcWCQLvPWD8kAh2QkmXMs6mJMM/ITWfRxDAzELHS2RQIiFFjAX1gWpr75d+M
LkE0tvzEvU4T6zUsWHxQp6Fc7KAg05pvQL6XccYOX8f/KFwJFYOBDQkCKCAz
PKaTFE/4PxQG3qe84cnDqNUleXjlmvN2yIjLTBitsNpB96mlqxM93sR0mzBQ
/1WiI0QgKhMpfcnpKYSkKyKcNNLCeZIIX6E9k1eqBxGbaMvUlwEmOGh2Rwch
wW7hf0ZSSf92Mp0TWyXZd6YtZS58sCIF/CBTT7GE1KtWcX82F0bktf2StaYK
DD5AAItZcM/hFCwoM033XIWfSgbeD++Yr4aZRuRgooFFmgA61iG9eBH+JCWs
f261DR/r054RE+EL8MJ7mcSPClAvGOhrhSSCGXWaPeYRdI7191+6nr1e4qo0
I49SsV9Pfxkk2wfD5w9NXEhyy9YG3yMwKuQ99ndiXjk7xavoqRjP8UggL6Zl
2WcgnDFeZ1LM837G+uCii3blJmFubcWzX6BVgvRKCvN9qEdGmLMFIOMPCdzV
PYkNXwwQkDM4D3iWkHggcVx3OQ9CI7b2dPNLkJ045QsqPVHTaP7eANYf2JWe
EfaVFMZkc0sncwzGFb0gFOVnJMZhEHGiUWVkD/IuLZtYxGFnhjcK77IolBYT
Kfh0EDZ7kWAaYvwZPCq12pfZYZTdHmZ+sihdib2FlLkKQLiR4aIhYETmwhdZ
DDiF0O3uUxwsXfuq6rdjJsIsWXq6OFm72NyGUyaMteBgMrLlqKgIgfCEKRmk
kJP22PY5y3aVPCnjaXKh3K3dvea7MDqcj16kEUjaxBn6PS6y4YIDUPCuqMlI
nFS/v10AuDviDINF5dV7bsiSGExQ1guFZMn57zljaJd2VXbFfwAoCYTZK6n6
kNpuvcMCRDBRyx+AZ4ktR9CIBzxoqaax+da1eVJV0BUFIs3zG4EJIjVOhpJs
bMX0+Qas2a6FVnEGDlvMQkd4+1ivJ3W7yjgXbRr6CaOLyX7W59vi671h3xe4
m+svx1xOBBTkSnRC0U0XxHFXAR9Sx1W6QYRv2jFZt/ykXxkVmzxeBORjox7N
BVhDrKkX6ht3NZhoxiAahUGve2lYd94Xed1dzAAGwgG/44sj7s9ORKeGIael
Cw0AY9QcmBEznHjiNLaZYgFgQPY7T5Z9H4vi0cgo/U4zHp1snCK3zTVIE75v
ITU/b2sx8KvauagAZzjR/1GO3vnGZ24BIOSGFLGzUOYm1Un3ic1r+jED28nK
GcwgBxzk0lf8w9uLifLPEgC07i5DKDhATHvn6Zht4HTNAIMD11+/vjiggbkL
1YNZbhCElf6GFm0Ct3tAnQ7W8w0Loh1lCgd46fvIc7Qtp2S8iqwVvaYYy1Tw
GdzvTNeabZuJtsqtrkjOaC+iN2uJoZ3/OWptWYllAvQUmj17O/AuQLYOnwed
QARmuLIT1JxcMOgNIPUfokdUQuPezDKns2rTSYbEyKInDg0svMGWMH7s9dMs
gC1MJRHvUnijMHtz1uCDxphum7uQYDji/414ZjvBBAKEoGqk84LvLh0u3I2K
RM5VItTFPu6XDZ6uekcWP7OaBG2p5Rr2eQbBsbnnXfh0Lk/Einj0Xm2eBBsn
IykardnkgIOyMWqIMwd4zZwMw9lmP2lkfoU1H0UY3rLKVLP+I6ZlochdeVzi
AaZNo7Tk4PohZfJJgyhOe21ON4wtd7KZkXTBGkV3QWdAH7JQqjGSk6NZVQ0b
lhr7R6lVzSuvfPJs6OEflruPx10Tge569AYYyfbQn9uGGt07qAK5lylx5sfo
QrYOkCUp1otCxuPM5jM0vJYVP0SjJyVG5U+K4G1nnipG7RC0AkCcp5DdvwFh
GPrLWcUbNVODp8DFB1ussp0dQmjtE1W04VqrtVdgVGKxtHFCshQrriHqbFq+
QM5j+T2HxQ9AUNqw8n+5Qq4p5FxYvA+54GxrhsWT+ZE6rHBGdL21aoZdUjtC
UoKjYvaP9KG5qZaAugMqmW5I18ufEpzIWtKgqdwwV7h8XHKoar7kiemOFZur
mZ4ij+cFrHl1bj8QTpSpVzh0qoyMVC3ZvbeBfeibi3Rt3MQu5cFkJUt12akY
P70Auos3NImWDB5l9KBHO8HobNStJeJol0CVhXwuM7nx2e4BFD3nIdcrGS7A
jmsIo4LRzG0KibM0ezJ5xZWIRl3qhRVmDzuJBpYQWEmtewSo/YYtAf219lV9
aVxu5NxlCXr0NpY+5qBemYhpnK2Ig4kYoRKDavFSApX8X4Uo6wgpBqy5M/9N
jXxb3a0sUswiKIXek148cLz65qbxq1seVaASEXbPNeJJyzbTs+/Fnio6UFzX
hXo3apfCLMU427bNDPHa9n6uwXTiZaVnrfP2cTJV7L8TOCA71A/BtilSMc2m
WSkQp8LL3xneLz8wlEaTXj1frnLvkFEIvpE/MFsWHNWNNp4t8hUfXLmyox14
fh+kderSEONJgyM0UVPYYKrM9+1L0cViR22DdaXeHs6N2Gh1tf7EneEuMBEB
cSIa0NKDMU5DlmUNMY6I2znYQ/HO4gXjeNzDZYp2C48IjbEJbxJ9BTWBkSRE
D58+QQ8sm6OPLlW7SVP1NYK1Di0efmuv7LgBTw7OJiLscjtb3VybGjO59W8F
UWDpJtAs+r+EEEnl3Hb7BbsjAAR3v1yc49RyAKbga9eOzothZx0AB4IaSAsb
oJNOU7qzFgLF8BIq6y/eJNGf/IYZKOqHlk2vlt6p1OKGCAfAx8RUxsVAsd/s
O1eKbNFqup860gV4YM+TcTsQdHiCndNvkyjMmkU7WSMuyEX5SHpMjnsyzj74
getsNsMrrYP2u50NDkiYsI9Ad1H41P+SYVy2Q+VUF1zBpSK8qllqr8Lq3gEG
i0Er6VYaOhrHiU1k6Swcq3M1iBjP5mfN1Kq0xghx5my2ta6CsG01TO/OxU7v
26LnF+YcMayvwOFOdYzpVwagUTMYKUhCEslkhZhDMGQ3kQYMJkB6tDPwE5Y1
99mz3NRU/ggoW7SAMWA5o+fOIkRBz0CCIsxNLAELflJT4te5UTHHzl4xcXlw
derjw3saxdXlUwXwgkGEnlPJH+69RTV7XzWUFnpXwlgAEAlCVsuwGKZ0zBID
MLvk8f4NzoNcgLeRS1UVSy7egg/fVcVJiLk5Y/YkIX9ewTOA+GckAWnl1qCI
DRCZSv3JkAXFRLEdWpGmyqFNd5zczu2RrFw3YkUln+nqd2eaip3cjlP8AKVJ
ZyQj05hcngmlNYedQ/qg476+kj8alNzSEut9pPyuReJN120IEHIG0b9gfZ5b
KIySMoh32wQVC/7d9umwkCKr9muW6IN2trUCDT1nzjKNjT+6rbhT65PhnApg
k8FyXuMw3PflBrCLFwOd4S9mpGuWABi28gUriNfLaZrphWGhfNG5y8C07E3p
wnHtSLnBomW9wpbs1WZWJ+vG1GtrfjJFwE0wNx5kF3CNYjjwnxCVzDYTWLRM
Su8rM7sVECK3vu3/ofqC52kCVZjYWvGzO46dAio8xJ77m5x/o97vgfwKi4D/
o16eJV/HlfYY14oNCBQc4BEw6zVqewhQ6sJO7HrVDlQVJJ2WCNV+41bBdUBI
gVkbpQAZt8hSY3C8uL68BM7t4M/T4yY+cUVwqFw1fhQFHNFBNCBZ8Odtmzrn
i5CWS7H75WB7C81bDs4GcPvKhc9n3fkpv6QyCXAKmlFgzjYEizKmrAjvFQSV
I5QxDhKY57HB7TXuxjrWIU37vOs9vvXdQprOEN5Cy5aLWcofk+8ZdrS4TFq+
RdVyoCo1iCwgTDOOI8IA2CgkO6AkgH+0XLTx6xuwUbjEYjR61ppwrHghEnEQ
kbMw5GSpf1pokw/zl3p235BzQVTom0NxjAmhJFcsR7/dee3GZDgNw0H7Shb1
LBUvtKtn3NrYvSUQfINtJx64/1Syh9uV1Wpr13/m9lqnpb3350m5Q7X3CDXN
OUudrFG7lZDmApg4KNteMnLRUiCRG4l5T47AblRt741qP0BGFHvJHj6JPI4/
gkSZnc7X/Nr/jOQmHUUgTrYtVdou9+rczdyna8epZjDEgnwVywut3zOPV5MW
HnadeYXBxM/Dkb6KtaJKjCn1uUt7B3TWQkVmyGToU6ha3Z0RiTgjlOkQfP+s
BCgApJ9P+IrRyRpe69oYAslb9EvGQKVuqSiC7PHvCmbk6OLSu7ZtJuL/GR0P
iR+i2IcF9PiQkiqBXfomukggnN9aCa+XMgw7OFPLNKjfmIYesB8XkSu7V/Dq
xSyMehKaisNA8SSJ8MGORHOC5kx6iBAA81XHqStf7moNhZJUL2IHp4la6c21
EooZmyYFIahmjIYxV3qzPxEPk60QDBSz5jBhILPY6221/VAHoIe8fE41nOZp
mMmdqtOkDhvArB9rrsZFmSCsyLoWJcq/MrxOfhbrJDuJ7Q5MLis2PNX02Wut
gIOg2ABDAyVKtr1q9S8lGpP0hQJXZltB1kQklBvLPFJ4F/mFqXtasDu5/Uai
1uokeUf+stMh0QX91h5B8u+9Pe9QRaxdWEgyMJg3riQ+viq34ArLzxk9iQAf
lxsYSvJ4PFVgui9+N2Hw3RcJNi6CBve6dJ8YVtrq7WUYVcTZZhr5LM0u1eHU
fCK3QGnQIpQZXlE7dFVuE/X3qvfTHfdLhQ0I/Jgi8op6659prL0FsPwclNPW
ENjnH3t7STrjPoAmI5ZscOXFKM/fhNZw2iXF973TchtSf+yDDoWTqBnl/nmB
jS/Y+2mQjGlsrOhgn7XC71qYHoL0TBMrWJTjB3eeNG375dNH8Vox4P6z9Blv
Tfk+QtLEH0MT4G/EZqdfEth8mhINlgWT4nprYE9a07LPv6/G9u/yIeW06Al/
XdCDfOamyCKzFdB0v4XgDI3zAQ3OIfw18OE9x8hSR2QRkzohPAbalhJ9txKP
j3xVx7Q2OrYfKqRNZWj1HuL5Pa2m8AuMq2J/MCsUPQRSQfs7EcIXCDlhTsr8
exMox1ZI4GxqJpsQkn/vlxHepNk1o9R+lVMhHTotDLbWuVH3TF1Kh8kINb6Z
7EcqkyGYKeG5cwohruBVCLD4LPhcvm2vkYJtvrWz89EsRAY/v70IMC4pTXBK
+//U70/tmo7w9TqhxOQsDVwt+k4T2tJosae9TnPnC4hDMB7/wk2mhIS8c4OI
+IzDNQhmdC1+Uahkha2rGZofA3ZJQM+6+Dqm5NBYhCueROTkVhc8G6Cqxfqx
yz+9c33UL1Ckb6NU1GGHBvcXOozcF6iezcCLE8dDZsto5QgSfkvm33S5RwUA
ZX6EAE2scFHf+51UEKalg1mDos7tSruBc2fA2UOKBifdn62SkwhwtEbvdczT
T/2TC7NB15u24GzgJENWxRjUJ7CNtXxJw2BupeS9YYwQRyOLAgc5YgMvOSO4
6YZcDYTAGf50UhIk7RY+Qeawp6l/q0QKG6x1268T8DPEcuiDrCWTSNWO6tqw
r1JjwKS0IMhqNEmzS99viFpOyI+KybwvHDvPiZ8074jZ7K/bvplrmvlDAa6a
KHUkybNSgoTPCy23ltEVF/sHt+KkcDs8udjkCZDm9mlNk8uo8weNQsY8qODF
6pAljm5SQp4hQTmHMU8oIFftmmLWpN3nkgpOhZCQvcBlW46KlzV2G40BJwWA
6d7UXkT0goIQP1fDBO0ba0SFwhyLHXUF3IaU2ym7KJQ3WyEML0bH43jOdUU2
bX5ppK/U1IUuHynor45HjAZFSz1hA8PN4W3tAYyfvVSwn46twK8A3IDtOTiU
4iXItQ+CVkw9rkM3ZQc3geLqyfM5wxdxpwvgvWbeYyt4/hnCaDLCQcjYTWG/
vCFLuBKGO51wTr9XXuJ07tyukOxDHnKuAS/SHIcpBw8koK4haNrSEOPVDOoU
AmoyQ6P9nej5oqz+Ovg684cIV+JnvVJPXqPzJ9mH5uoir9+GSygpAo15jcE7
RBFFlIXOJ0El6YjMBOv9IR5uzMnujMuWmNzI/Q/YoaBvjqyiiRkjh0ohADwr
RCMIZRfoNLJ79INQ+ZOMZTwP2bRFIltQHMHsssvWC3++2G6v792prHvIEtNh
Z7070+YxspYhCZ3tt/ISyP6JjuauD7FxNvfrqfGBZhRx4TSGMfUkvPKDY57F
1ZXrmWI08cC2GpAVJHZx2kkAbAhvwgJexVrtE2PF8E31f1BakFnBmCS0CjjY
+QxNUrVnEKm3PXcWCeicky0h50PomlVw3O4X3Y9tRjcwIzzLS03Bv8ykd3t8
/6E7aSLTxiLxX9KmUh+K25bUv3o1I5iyIwdrsxJoD5rtJSygFDjLdAd4/2n8
LBL+w5kQF6EmHH6Nc8NPTX2a8UzgBf5pFFLwIUt3DUE3VitcsEKcKxBFj9gB
wZecekJ4aHzTvGwKhYclZrnqd9Zm/j/BpHPyhgjbbXPLq6HHYPhkYyhe+DYo
3lw7Sy1HE6Fny82GUERlBymBn87aTnFnCBrDqPAWSNdLC7D3gtls2RgF1xM9
pwUyRjYH+laq6OSP4q0OSfkeCktRA/1/Rv4IhF+LabBiqKmPHriF9nHvnh2j
ufarGFX3mUcuPw/CgFi+7+tFNzyJ43eHu+8hOLIKhDijBeLlSpqQ+fub5XpF
1U0NoqVAuZswiEpbBs3MKW2lJ1LA9I8+yU5YWB/RwdzYw4QUljWd9Iu9AQpJ
muoLIyIBgg71yKi/34NnAdiLROApvqIIZoIcqd2ma8qvCsZ1CK6+03KArOvG
FCuWl1NRaknTIiqo3Gjtck+z56f0Zw58a28wlBELDWW+wd4q/XV4kIe4OGOQ
zAsWDw36Zw0wjFF0JUdi7ImfsSayVPeL5inyye1i+2aPgdyY5lquvB47RCSD
Fql/9Ql/wFN/xC8wB7mZ2WX7o0GfH2ax+vl+E6p2IkfRtLD8ROxoY3b1ih8r
4AW1dYw5pS1UmKvXriDxese41vR9mKdi+/JGlWTjXu3aLozKNroayN4VDSZa
OHge3wGlHVNImnZ0tvqJTLnLSuneo777QkpfPRcWNqsHeMwh+98jBM/AEKHx
EIe2l3stlLF0CyC7wyOHikZQnDYVbNXYBvvAh95d76aBJOdbF+YfNO83LxPJ
x5YTkGrUddbXho7XsPHHZg6wUzcuQmcjwllhxFrQf6P3Hbf8C6L9OrIbhBiy
+/AtObdDKHMhd9uSO6J5fPEyvLsDR1ErCaMs3MOZ1ZB2AhsEDE9dl5ye2S+z
gviKC7HtsXO3JZSK0RnX0A6wd+qvbUEbKeKE4BJ7k0NK0SUsnCOs7w+ABAhU
a2o4EuX5HwaCS15tJA4m18jxz977q3sXHIgAQ89XRC0DOVvZtlUwtnkUC1aU
3uqZ7YSqPQvYc18nTl8KHNAz3IRFRi27sq88mZ/QptNS/3DocUjxlm86/ACa
8ZuCciJSZ0ljF+2lIYRKgMjD7t0B9cJaSUKwL1QrRbDZvu4gVQ3xw6pfYDDH
6gsDYeJpTe5thQ9j8oHT+vA1arEOCrvbASehkcoB4glXsBNvuxXXPARcj0/J
aUAZ3SvBUtiOtdNJfEXJ4tsi/5goM0mq4DDPnItkVen0kp8XDLJMw6FGK4Lt
8z5qmRq1URY7f21HdpX4+XpLi+jDgBxBUpJXGaCHC4y5t3OA8fYUjuHmbjpY
BsL0mbAVrzoCXNQIz8TvYlcYfxm0XWJJ/UY57bEdlc0UqwlPJohPfG5tiQZI
NjM3cJi/VmdYvpo0df2wAMksTdockXPgykxrUdAkLf8jrTHundZoSGOP/k+D
kyju0amC8SoK7B6+kkBETpUbZ0sJ/VU2dhC1/MsKnZXztw6wHPh5lROp7EmA
xAAb7jUc9ypoMHT3axtAx1h/264cAYe86pfKqQBFdkpaKnIaxW1jUCgcbpWN
7daynUyQdwI488ydlC/PT3V2VULgOibDl7gkzVHjIsW0ixGEF8e2Us2XgGIK
PSG90L02hncxdLJxLPJ7T2WY10jNkI85X6JVQnvNY1oiEScm1QlXCkDDj0sT
XbOCWghuy+rot1GjQVo1pz/nQ2hv3QEX/23FB6Vi6ZR/1gK7YA59eGxZApY1
kE41NjJrK+YSPvJKfexSIow3ObInQFSU51lPohPemEosSCUvqt/4bJcICZ66
meLDTQ78JLI422iAhlehfAr+8oERS1jGROTzSjgfdKtZIfb8Oz+UpzK20O6h
3NviAEo0TZCDFM2qzhVVJH+iRH95KwhrXG5hAzVHLIqwPQ3msyRmJ/swSgCu
3EXPzuVE13B+8kzdmrzsupi6oai3XF5LFThRh/3JZYI4gTNvQ4sDnpuYmnCK
EyqnJYA1aNAh27cNMtdp9mpJBdLsjzriWW3C44XAc2AHlBATqiPus7eC7O3G
F+efamOki5DJEHaofx98GdxIC1e1YXEINANTZ/lqEt2rIxp/hW1yti+hlkrp
vJ4H25Aht4L6quqkQNChx+/VYwbPsahZ/W5vvR/NjGFSpjSREjrRpiljp7k4
WaW5XzTF6vCXIWGP6Wd3w7yW6Dw4bTMGlgv3zTF2/ciyUBo3FxFF04RK3IEa
d+T/q+VIPInm3AbJdr96mwCLxXZ6tfoZ/Nq11nZMNfZJPht/cb59OS+nhPUk
XG4XAX2pZknS0yhEgTamHUNJrOs8cMl/5+UI1nD0oTMMg7C5lkxkNPzw3YBq
AARhyIs5+PWNX2o7c7asym6dqtO1nlUXfIbGO7Bbi5EUSOZ8ydMqxZ1T6bzG
LHr+m0TwWJ0AROgA/eWdiQfQDca6AMP6NDkhWVbpoIfmVV62jdWBuFwV+V32
ppj8BDBiuPgDIfQQE5m5V6XPV2YjLnCY1EDP9tOJBLxQk5Rk2zvKKSwSk8QC
6VLahORMWiJpmdBBL/UfOq84AUIlhm+MfEELzQzDPPdc6qE2rsFDqn1pbw+Z
wvzhhLmNShqfk45zz7IEQY46tKFvNgwAmJ+e0Uht+Bp1ML6Mk1Txidgid4Yt
fga6PkzhhUlNZodf2OciYXBZ2ExD/fQc/ajXP6rwGzoUu1LYMA7KeNDafdRx
e2aCBvGjopblapYdpMgVL1Bvl+P8e/O8Uu5piy/beOoOSPZsn6cz1NmsA9gM
gHux4yCsEoe5uJEy63yOWxKY+lv1TK5pXuyrSd5CD0v0VWpDfSqNP9ijlAhp
bF7o1VGy75QOIe1Q/PujVtb51vIBpYITvmFQp6ljIT8/u+C5CZu2i/I3i+XT
ttozE3qXMMa8Zw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpeibK65tHG4deYstdWtSTgcZQys+G464Ot5h59RjNuouxz9U6WoXAm8TZmY2hlouJn6K13tK3V2TAKQsZuIaaQ+biJQiQUSktxjV/+bwB2UY00ynfuiFFh/khDaumHkfp8un6XE9jaKdOQGkgzYQ0WI7udJ324Stf/VkyOpIjNVJoP7wGGVU8r0sL0vzro5aCPV/PbUyDfwKDXK58Y01qanHT+AJcQluA3ZXULhVd6pRw92b3JNs8icGhOpdquA1AH2rvzdYQvAH1nrCv916dS3S/LDhrtJRA4hCumGfQdq9l79Uk6w/a7RSgxg94Ye/D0GRCEvxgApOYd/km6SqijBdcM3eeRrBYGwqkYwd1f3P1vjxkZZUva+vF0OJJQFmyxPYhbrweDjb7CBMjQrNm+TMG80zAmiGp+/JxfR6dGsWIj3bqRXzgf9Kp0NVbJ+Al6/l1/q6Gb5LokfIO4TCczHgjdUiw7rJ1KnP0EdDMqwJAtNIs5J2toHxsELE6rI4Fo1JRUpnQ3vUCTtpPLTAaCU+OwGXDG8UWeMXn5OH4lAeCGfu98W/YYq95mBlySRMyUz7bx51ZnHg0+GbQK5A9YGLJi7sF+i7kGn+9iNL9/M3ykaaUijWb1eij7XyxB3ZZbZ2j6tdtYCVps9Y0usZZeMbbzDpKEojZbkAVBIeTdh10/pmp/ctYa0RWAFTtsw6qHLVLzuoKlsiM5aeQnUJrys1CfABTipbgQBtJ+BBHacHkMdIrWa/xdY54/Kune0mi5mxK69gezy6sYFpnIDy7SEV"
`endif