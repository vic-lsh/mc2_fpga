// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
xbv9kwAPaq+Vkk7rbjm3rQXQELbMGlP/qy395r0HbNUcaGyQYp7cd7BofMFH
E5HTs0cBcBNGF3JIn4NxWyCZcBltsnEY6ghoe/nMmAE3CUQrnqPG3nIm6yIK
3yDJGZ0rqXon1yP0F3ozwdGtvnQ0fdYGQkb3mT8mab/vd9CUiNrFdVWGmCnM
NBdJ9UxJIkEsSsrFok5fXW3hT3101THsnRHAKv+Wh5qUr7AcHY5zD/0TU5tP
yTkGnM74xnXUHu2XP7gw5azFGT7CIabEKXW+wHuh+Bx4gv9OiiaOCGBzrwvG
hIJWOesLL+qc1v8WwSzLu+v7G1GlKcadbD+5mZu6tw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Aj+AaRzzZdaiJdota0XYJ23PaEtMTZqTNpPDStlhPbx66ZZVv8sJICin44ef
g8ki9rXgMWJUU6/oUxHVcN8F80xk5PlMSd3l08/vaJnc5M/2+p/lbKkkyU14
QAuvfbI9xidxuQXUPHZaqHo+SjKZyyIwz7ujQfhM8JZRCtA9fHcM+69IdxFh
whINBRHqAUfR5v7xJ+T7psCfws2GjalBTJsqwKODUvqpwxQmz3M6gPZyKvdn
p6IbInX6sxZ9/rMUngLtTlAAe6fVJgOYisbob2kgqKj6OoQyWwC4zuInpiN/
B61vdHnQlu5XP/UiW9YiHvLTU0PCBtGp1ozqUWai4Q==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aV8n94cV4QIifRTOh9M2+44l129YWSf7i0TVnPRPiGVO7wxAjhmTmxGqbnhU
t7SCBUml1l9m5Lrr7R8bWGRzqzBLDOiJ89yF5WtWQl0ipVpRV0778fSkAFmI
sTAyta662i097deYoLwebdi+ZnpvMPHbCN+pBEm/rUhldrl3K8pTsfYdJ6oB
SQbS56tk5XRUhWeHUaTEIhAXZfQCzZ0bRs/aLGQjVNClbt41LJTJag+Xm4mO
I9lVCQE7pbC+w+fD1x6dMmXPQmSklNyeomWuWEb+KgvE6EkeOEtNXlGbmFjM
d1GveCSYoQ23KM6Jbs7vf+vFW1sZGHtl3zszP0XwCw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WgbC1UwOSnMO2FwvXDxvTxjeshCRnqD+pFjz60sskGJfp9GRIXvVpTpX/UQ3
uB344nXlNvhyWiMUVLHcG+7D3OLYHGvQ5bm1RYuuIZnMwv5RRMgPoPTOfdos
1MpN/pwW6Pwq+rcldO7O5X32KuPgDe8a7h6Fbq3Rssbhv3e2v5F8HvATbRMI
ioZmd62nQuIzDqQjrTlpcxG0WnB5LdMxnI/cOFvGQxJkdSm1PnjvH9Ywc2t6
MmU2nQjWgLiTZ66bRDlx4fYTkol2LxPOy45SaTNwgVCQz9naNot9IFcBZyuX
8v32BUGhTIO+h2SCuVr2vX1McKddDiCm7rijv4rVhg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bIVrHxPTgnEiQ6wMRB+eRpHUYGXvMIBjkBc1vxo5k3CXiRBLtJ9i6nRaduSA
zjpq8wymA5RX0mgsG8j8jwqwjMfYooMxR6Efzw53ct86feRfC6t8Qbo/18wy
wk1HeTZV58yTXy67F2Hg5BR2+6JlbGuQfPqDCaDMouHZ6nYFFpw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
pChl5mX0jyGmTUFifp9aF2y3XNoFQIjFjL1NywAGyjEGDX0g2y8fxXj05dBe
/L4zV/PMHgVpSscx1zgcggl1wbYIkeYQRxufr8XF6xT+gni1ZJXmGxG/m8Uj
69fz+l1l40LqFBDekJ3jQxKyIp5SCK6XM2vtknTRiNcKsiKSkIZjB2+Xrj1S
spFzc9YFfkRlaCEqShWslWfyi2Y+K30EDA6UoyxKipomypoFIgbcoy4XGyEm
D5w83kmDI9AlSBi5frJt0S2gqk+ozexbqJcOOssnEA/EGj37K1xUfCJiGF+9
OLhuTmzCmcmh0iI0Cmgid3XBLrqO86Nt3Ui0PULM2xwXfzJgdytdmpPI2cch
402bdQzymF5t8mtg6GLjAtF85eoRi/CX7ZyL0//Dt/GhHNJ8poorYwUkojJV
9p+K+kkp66nw5t5uZwrVXSEQkoYwO4m5dT+900yVJp1AQBeXJ8X9IFe8kKn/
bUtV3baF3Q5lk43EQAfvrpEjMJc/1s41


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ny/fnbdxk7jTElKBe1OtmSqOB8nPhI6TutEwrry0HObCPo6R0O/AQ81fWP6j
xB3SjiwD4eXqeYS1reR2ZImkSpqaFqUCjdxO5UMfUx6vYXqxolywLkMuPckE
t+EEufbST+FnJXpLKPW3yYOtNjM7oa2KjcEeLm8SogWuUm8cfhg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HETG5E1iRwIjxzg17fwYlzpk1JXcwoeBwH95V1RO59zzmQlhsvdq9n4kFH9b
0bwex5uMXwaDxsD+XoJqeotU9EWvvqWiwoQMhtTdxihUGyMeMVKTcNieNnwC
+bhS7OdWh9dtfE0OxWgvjp9nA/t2JGVK3X4b6gvU2EwSIBptmbs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 976)
`pragma protect data_block
FCUK/VMltxoXpu4wUEs62Und3wPIEekbpA9/wsF0s83UnGQD3yJrJckUqUKl
voZb+iq0UCm+AloCiWGRSPbAORLAXA4et+98P4y8GL4tgXEf1y9PLOYo5QXv
5sqGnvZr0kP6+IV+eEb5viZZGorZmw4c6xT4gzFXO1gWkKsJ9gtZ3Y9juJbL
AqgKjpJ+xmQBkCTq7ovIwQZNNogzfSuyIhMipIozgAsVYAsApvVv/7lTxAnW
3XDPvNY1kkVZcktk4ZA2UexMfEHK16jq9SwpkEJ+0wnSlColMBAwneyU8HlQ
M6w/8rdAfUWDp2zl+JTu7e2n4yWZzd60ppxOiKK7YF0YXeWIAk5+QfceNmKw
M9xAIFzRSLFQzBAFu3BNCUVn1SY3NFWfZLNW2v+Y7dmAzO3MqtYezpJqvwrs
xfAwOJ95ZNKM0JMryo09HlelL3wlwNH9xuQXMaszAKSsKpOVOgzpLzPgg+18
H0pfE5dK4nZknQlHiQktlMDIsFIqrsxWAwDrm/2RHNqlP2hhCmrwMcaxCi0G
xjzAWbPbrkTu+zdsKSt+hFOdiOxe3F+12i0DQ+2De32bveDb+WRFOeO+cOhZ
I1D0rrkRnnGeYuFAnMskJ97VNWtutOpqdmN/YMmvO+WH64A39O5RtWjdnr0h
B8x1TmdtyrvlkCxwxCD+UlvVhQ8kMYK5JeJJ/as9wXE2XxA0Oqc9GXZ89PhE
slNeE7PB+HANuy67UPosQgHI2bKlZMj+/8QaI1XnzuX3M0goRJALOR5m+Nx5
O26pQXy48/Be3k8w6XXEIhobY6cFJACvp96CC5xBHkmsH4xGkootTO1kfFyR
qf23VCzWHEIf12QRhupDZ+8RMZOirSpWPVr73/xB2oeKOBEvbwxI8NDgWnOL
/hEqfs/LflR54y5OVtR7q+tJoWkJz4XZvaIwAKx0e1VWyH6Vd6K0taaJ+uZX
ylOplLjnYzYruersWAOm+h5L3V3Ru6greBcgjpKE07VOmUCC3RxzROA0OgUW
/fCkiXFXO0u3pYFs5SeUkkq3dtUzf91PbagYzkSW+bQwZvbhWwL5RvQPR8nQ
/k3oEjQX6dN8qR0sVwuHYULbEMFeYF/zcr4hl+BBUYhEwCUmiYNmgWNJ39BR
lghZx5e0iN90pGdEwQD5A/np4+YXn6ZLa5ukRUG2oAgXegVj7VUCUefA84NK
pU7/iPyVasV5Qv8WX9gQMu9zFimFbJJ8pRXRdT1zYOOdTFIxpKcA7FzVySis
B/xOzhPrWp6pTMqPUBYRhlaR90c0KWUcUUCZcH3RkQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqdjlHbg3H9fsvtskHaKnxIgSZjvXIEAU+h+6WiIcoEdKymLLAjHkqcgrygAHcYEdAH1+va2fNLbbCVfKSjl2tMABVzr9/b6QwH3jEfUKfYIkKDP+P6GUvoa69dfZ9HII+i9N8mPfxqTodh5jCtmOau+Pgg3qy3B9202aDo7eEAlo4o6KeC8GEiPc4q/vYcNsCziDS8UabITPhMKgB/Ih7GHgJSUHFuvxzjjeiiMg3iZKl68tlHNEHlqgWNtcChfZmQiOhCw1OUIY359ujpK0deVlD92Ozv7lpzXUcsjMUyxadXDyDd+DStOQHNaWsxhyckutg1LjmNpnbLBW6dPs3/H+545ZfzLCgAEz5K6NsidOyI7+t5SAkTJKk55yd/6QfSiFloA0W+JKvwLCWRid8n0EXJnKcCf0Uwt9z1JTnJ4Hcd8Pr3PjC2lpTdiLcL5wAUPBdIIp1AJXQNC8yEULbA7WJXMaiuE5biLtknAmKmBIyUos5A5hkhnCfmPht9CRC3WyyjHXgfmSibeLop1/hX+ptxjsgDA1pT6zKxN5VaEN0Stp33Nru+N4wipdjs4azeAC/V/pl6RKBZxciAoA0nxJnGHz433AyH9CQqGQUSy5U11tv5ML3oroLKiGhU49KdgdLxjS7LrYKTcHp+hhBgZMZ1Dfx0ZVfDj4x6r95dxPHXp9ClpX+TDiGYPTooTU26HGkv6IVLfxoJwofwfOnPpurE1bUieEvWOMNLLmsJBxEVUzc88Vw0tSAFe+bSsL+WLuuRrWmO4zZf5cfILS7V0"
`endif