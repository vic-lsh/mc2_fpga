// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
og4RL5OpbazMDTSigHByv3VXOdn4Zj/4UngoA3S/ktQcWT9xw9nm/zt4Wn+B
HkNGjif7XQ4bjv+3VgukKNYIanyulTjxYQ+v3SYuvy3Lx3V+l9akOeHnexvj
MyAy5Q/ST5r+SLOnHNfw+NEHqkpmVyTRWqxAVtDY7GcyHeB76rGnY5DPuq8H
zwuhe9wqmq/WF20j035CYGJJXfrwuZ+HXUjXRBWVI1z16ddfEoGW62j1g+eg
TlwIaKKp7cg3LWmpyNElz52RJ+kS82665CLaaNrxIoZmdOYk7PF6BRLyJ7MX
NDeRY8pNf2MK9PWrvsacKnYcUCVg0VoA63G6YvXwkg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
a3y02VYeW4IYCqV5fL2bTeVx7SyvnwKhsnMh4Uyul7IFbMOwrB/KYtcjyKUq
hHjoLcN6SqPCkDIMqkIAlzTxXmtX6hflDagabqDoKYxl/zhewRzcmPFlRXq7
Cd0MVcoSNdwj4gDAjyt+WLLMiU8h8lGpTgZxtO3d1kWYSs+o+V3Bj6AX/ZjW
lUHTLnHLa5T/LeWo0P5NXs8c/M6MgWFBtPqtsLyhYW57jmRKBXg6NxFM+Tue
gteTIb0D1HXEj5DWB+xQCkBfPAnZihsIWJZCLXdH3swh0HvenUx9k4Lhc3Sa
3x29bAUoi7gQF5JHMEK5JvHKly2xJGkTH9UyM+5bdQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UtcHXs7FiGqTtmkHIpKKugFzPB8aNhnBCUFt6Y4JFfY9xZzqYet3UgFV2A1b
Fv2Y2Xa5CQ9Q///5ffWXymEW6BI10gwlc+l1u1XPpIG+SBZC68j8JQpn5Hg1
QoN9xhjk4aTmPxSrluUZNMYM4bKE+5XYqO4I3InJ4zs8/MKIIt/HdqtNVKKz
mmmKJF0QvoohZynhr6zzRo9+pTqj0aY/AD35ezpn6BjGIDdDO/kyvH/ADA58
mfxM4huP7Nvz29UOAldlnr0YRXLF2B0wWxerWK1n3yF76vc0/iY035MahcRQ
vyZBYvEqJlg1ACgGOtM21FAPgr5jNEIEznakcGo7cQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
n+qn2XjaXSS83CA7tUGgpdbcttV6QMRR20/BvgGZrjBf8wIQ/ao544diKzZE
Xunzf3vXS1AoA/7Z2YFoB9IROtNchn0vWuMAdP/ZO3LvC0nW7AQ7hR11DX6m
qgbqVOssT2nYGx6JoRFYb1eXaI5n1AioLAgTqlI28YrrlUhCbiV2sZ2i/Vw4
rXMbCJJ6esgOA7fLShUU9ShJoo6SVL4a1iP7q3WBii2FNpsMEuSkFw+VebUT
swirC2dzomPSGZ6bPY1wapyrp3EKcLhCjblbh7EpRPFnSnfqSzKf1t/3doJ0
drs1T8Uc+EWOJ2TF8LVrqziEKUskhc6lNTO77uAGxQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
E5qXxwkpaRiw4jq7aaDkeDoHdsxdYeaMZDJETYfrXD+JCRj8SdttNfkuLIOm
Qcf/Ilg29/g8wlHqQi9/3jyzKwTcF1vl8AI5DG8J2GFGSHrcb+81DoLcM+d7
XeGHnwLcFRPH29anWQh77hIBpIXDGUB/MtzFyPpuWTvu1TPn9zk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
FrnZjYoG412B2GVpuZf+mn5MmQfT0GJByCzljurDtHb/RFdKtunWqUuxck1s
i7IbzhEOApNeeUurSfmdy5fnN5cIlu1w36QLyCZeP4fjr+Qi4BPny8Kc6mi6
Qr8jL4pYytJ3lZZ76sTAYkMh8JXORtF+kN5z88d8wqPxXVcDKE7SbN6ajGh0
7O4XaI1QErehqCoqJOITGTsZPHwu5XwpmM90l4617ixA7wx6AhtacD3NHNE5
t5NG271oWnukA0luiFLVDoayCUCDcy9FkHn4EkcFQivSMAwlGpMshwSr4OTf
9I6wAxjRpmkVrWPYpaMTiDWaSlx9un0rP/nNPaYgi+6zPsnCUXQxrJ6QBHH3
shSFR2t6MrO08cMu0JtrRT3ZFFrVUvZ8F5Fk+d+gf1LtTcnUZYeRG4bk9C2k
yxpzFrq5lseyjDHlYt8E6DADR6p9m08MIBQ96M/p4WfaKsZ0WVXG6PHqxynU
XtoQYByyWZL00NHki+YjW2bvL+RZGRyG


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nlE52O+sszIhOkcxmGcOnPjUJDSWL/mgO/hOodzq/WEfIjwqslwnQQEsR0Tn
QncWLMAaTQeZ2nEClR2RXcEjxWXl4trR6JuKIezlj1wNZY6CRQAWaXmDpabN
3HcNEvyn3YsQgH472MKREYDjWK9FAqv/Sua5vNdwEZOvAtIJxuc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KR/S2LFxdcLi/WEgnv5CcY8jM4d+jh+jAE6x8jiWEWkr8KWEKKck4ops24Wx
hrrlih+MRcOYwmRJFm7KoZoDNXKR3LFFscaYFoHutwFsd7nyrA9NPUea1DgA
84N/2sQ/06SdctXamgQcEXY6OJmBMq8xS1t5WXfZIP+EhJDK0KY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2470064)
`pragma protect data_block
6htIuj5QZXVAyNcJ2fKXVB6SHe2tfvZO8+LD5g8F7cDC6DzXJQyhoQcvLhEg
tX2ICJNW6dGXbSqpWhg+vufYj8OurbZFIF4mKlNxnogOauiJcJaIa4gauO8U
me4C0SIta0hBtsrkmZbhKRICflF84CXzhKXT6HSQR8EqnkBl7uZt8Gr6VPKY
BfF6W+fLHjuVjSyfmvEgbm7tDHWVQF6EImwzeXOsG0TFjDKboEXjtM9boWBu
nEKMHL70bh/fYUhfNPbXqQ5+u2US1JkyGyPGz8F8alJuFgKWbZ0QiCCNlcp9
TpmQEQd06CUJLKja06kbDitpIZyDXXPSYxLnpqwFg8rVwoYKNocaFiXCA2L6
1GpSYUspNYUxNKMFlG4C0RNz3onGrQ27bGmz/tL35pVbmH7Y3qKhMPTEl0VM
D8TeSdOTZuHa051DxPcvePWn83wWTMURPIcYJReh0HUX5pexE6xNeaeEuBgk
FbJuQ241QuKFHs6sC/Z1i7AUT9FeGB1XCPhT3zUWr7wm5/IBrGOABUtgDm+7
xgH783s3KFI0Co/8vBZV/g68qp7kDKZHGj2hk0HhYpM3s7T/MhwX7L4h/iI7
1ZteCuK/sGGYIkcVt6ETuaitwYo8P/N12Ygz5bUG1K9XOSRZ0alHqumI3z04
gqZXQs1VhK9Xv+NZk99wf908yghYgiSTHNUXYwJbtvSVrwCp2r3YU1MFmvYk
lyHJnv/OzmLT1QNCi5ZlgJp/V9b+RY+f+UO2EYapMpeFQBaXg7XG3aooF1bz
GA/VSKNcLBDSFc1dSmuLUbUzonsY1IYdQL7YHkcb5OPriAWBKXPmSWDfjaml
Y3j58piy/VBP174CObBYsklf8/fy5xwgUhgHwXTucLudxNUjFRYzhzTF3mMH
ZePi+d7Gbhf1000PPllUZ2SxjAJ02/NG4eLt5h6F8r1AxiUDKfIlYQBMASJI
JYrLk4QKtW6tLNqRJip4HZ8ZgS5SIBlLrtsbcYOaYmh+0cCkO0Axpf8Gkqxy
NESjrMehSNwzWbx+EjirUyV3mEG7HPuBQmVDlAEH81JuvqMyYFqOWMs9b3Te
HctCGImY6PjINjTztA4sCvRdFxLMeDzHoAe35jk/qon2Y4Kr9bB2S8wFgmHn
NO6TUf26AxeeL1ZepVyVNsd9zFZaMEwutAG2Zd6hHznK0mjLYIeuPU6nGbxP
Uq/3fnUzPg9/Qo4Ve7Dcbge17nUuTn3OcQrK5lfz3DDXlhDgIfsZsHjFP6gy
idjJhZt/C/8GWPxZOuOVlEp+iI6jSH20TdP7C8zWlCAIL2FBtWnyclmyKcWt
9dv9spAft8xz5Etrg3v8pvCkLxzVHhr/29SAFofNxyvVnymY+J+CAyWeaiD4
vG7KV+H1mG87Vjf9ulgh9NpIXG8xSL1dGbIN5DNhRi3K63iyaVx9Rv20x01V
peQstWmOqRQZg2mvRbFYKhY+P7APvivl4/JfHD1ihWXs3vxcMgjRrlN277nx
Z0TeVJh5RLpp8W0Z2WnzZLNWkj5h0cLPD4zQDwCVrUG8fD67UOw4L3Ti0gDI
Aly4yoseVrqcg6tQV//RR/v6ofmOTy8XcVD52NAy61X6qDGD+lk/iWdm936S
GQUhUbR8cY2TlTZhEhXlb3gafw50HXN36aKCXXn++jHUaQmGmidLkVwmx7HA
XBQBDBCDImazmf8e5zJZoKqyaeJQ0703lrEig4goQNhCUDjUCSZAK26yVIVw
yQcNMBMAWxBEVQqJHLKWh51oaeE+TLMSVXV1HEIkUqgZmr4Ns9KQ5SUd5bBX
Jjjr36YTIvY75oq/3UHqXeNv0ya9A8jn+azCNVmNRySy4IiD1qj07KRrrROq
8O0DYSNtkBZY0mDaqFPeLj3WxfCfn2taavqooK2jlEFVy5CI9hMgrufaDQi0
sJakHvPKi+kTLvJ02/YcNXNhu4qTZpnj583OFC5u9UIoJXOAiInKe9IGqpOo
H11v2owSRVMejeHzCOlfGYxm2Uhzddjvckl5LMdQi7lPbLhGb7ZkpAzPcaG4
znqdcF+oFDcx1u2GyohsmOgsdt4SW8bOBY53Ge6Wz8aA7R9ppPleMkNUOeBW
X1B6DJJXq0ZXiOAmYL9nfIiuj2RNu0BujT6tGJLOvpRUJqEfqBPuJV9bEGt9
lhRyWeZGliD+bc4T50pr5kkNp1I7hPbia9OlpD2PrmzL5i4p2W2zVnEi/KCy
rwYd59I6z9pvBzvN00hc6eLqrvYe8bzVNZp9IaNgT1zJi3mbK1AF8ZTQZ+oi
uc606Ox21Mgoretg34fLrVH8e2A6BKi/7HkaSxd9qRmH5qKqk/GMXe0SuTfk
YicTWjZzZ+0nRA6oSOuCIfATixXgxLoBwcXzcUBQkAo8mbn8OnaTrsU5OcTA
AjdusdmFlYxx2smFOpjnMAEjzZh5zhZtFUKR48eedxM8l0A9tmcIHeDZ175d
XPo6QQNdrIhUOXBX1AJ8JJ1jUSQx8T45/RDrgW0cENRRPFY5XYWwplNbj4vI
PPTKFjO81t4l9bivpg2hQ71UKl5/xVAq5dcvxkhSAq9/LrISqr2D6LIP3AKG
PcbHyq6bgU6yaNhFij+4igBPDeFF1ZgUdgiTRsQZFk8d9ZNDuI/O2NcSBs6O
Cis1828ROUOr+w8zyOPE9xQMX61C2mLjJftYIWh1Vf0UStGMSkprudiuHYKa
be5s9dIHTmZLJ70vO4DyV8misLpjcJnJKt0gP/YkQ1RT2dUEYqao8svOAtPc
53aBdvJp7/0EuNxYjRmDZM5Q2kr+QUaLlqvywscPzX777A53MzdwjwftqPFx
L1T6aGoAELXG+od9ViiA52KZh+mkJx8CsK3THN4orXgwbxp4/yiMq7UzkD7B
uaZNlkGIlrqdeR30cYqRA27c7wzksfhHib/cI77he2S+rg/sQfvPx6YYqWLr
gkPL82kpRsguNCi3A+q5QMxE0Wx8vJYHxKfqs2Usj6iBS3VYcYwE6clmbrSX
srFRgBv4Y7LruW+Hu9b6pKtG4CnsUeMyD8cLGM2Evs6kxvSyIAbkHRq4dLfr
Kg7n4N3PdHratyA68ICHO+otT8Vx5ge3Jg34KZlQXw1C9/KHHob9GhLNXlfB
/EuLgd0LfOOrXM3A7qQFWj2u3kdyAxte9hQ37eiMAKgmM4e/J6fUF5CdP6Cb
qOvC05QUShcxwof8ptS1PeYm6vZZKYsZERCwZckSopECbfnQiVP8s2ahhFdQ
V82aDAHh3YOD0x74TBx9clpki1MFopisZo+gZCYfvqm8NdUICqAFf52RDlHj
CaU16Ka+gQneWLVrHHRgVln1MGeKRsdR6sxfQrn37xvCDDfDpn3TpfVomc1p
XzMFbyDD1gTklRxJ3kULo4lDOUmVmXGJ0WuCGcJcP/gn7cOL9ZbmJ+h+qDss
Mr1s55p1KBpAB59OBawvop2vrpvrI4kyaDO2Tf/owm/kdXs8PeKvYOHJJm86
vazgpUy+OBjf5u8xv2fg8LtMA1hBx7RnJRGBDB6X88fKQB0FJMH/3QPzlaqL
5uXPo5h++LHk9VdnjBdydjaA4HQLYOYBx8gkl0Jw2vZqRyyuKj7CSbKuOxbR
Dm/kV3LqWF6/VMo5ZPY9dz95kN/4rqE8iAuoHO1bsCZt0fsMAdwu1vsjKa2l
1LxhKtVRzSvCM1apzWbbFdQvb0kCh4bLMU4ZaqLzufzdplh00RJ5YlSPGFS+
/yVVzWh4wikSL/M6oiLfg6f1vCt/JksGiWft7mRYI+/3RmBLVNXgsDcsLdvJ
Xl+wdrqNpQ12tinmCxyNndkVeHtQAWjUgBJfU9C77lhzKvetfRHSZkChKo8b
K30Jpmp4hj5AoYybSjBpJqj0lMB7hV7O3YOiLAjFqmXiIc+lFmureZzVgwed
fHfoKnIcBacnlU7CV+95RJmLTNE7OmAjX5hc7sDup0nbdBaI6fgBO0P38lEd
mZtz+QOTwY3pgECnmhU2u7Jly1ux134SWkKFkV2Tg8bJMcLw+HDdFqMZ0aqv
/3RiWTE8cT8Xhsk2tSxJMtKQMToUWTXf6I0O1i3COZraSlLGVcaaN8DtzReo
4QIqI7g8jpKod1O0aFlRAjxhn4EF5E9Lpo4V9tkN0pT5tfZGJMfr7TgbHpR9
VL2/9R9Jg2c+4V9VEv2eglZbjTtsj4tzi7/KveRtX/PbkujUS63HS1jOamDb
zyOUDvE7vPU+S5aM+ZiMW7vXspLiiacBMwYCr5lFFP3ygURK6VX0C5vjIDsn
mYu0EvFp4IhfSfcmL8m0mPgo4KyGd679Z9ldmPfi3wvF1BelkHOSTFO0/yH2
IiFCDl5yHAio1hlZj9ydl7qaIc1KDXUCUnOb6axEdrCCkig33Axckfh6F4zp
Jx2XwBy5M70WxRLWrPYt/bYpNgGAHUYiv7Iz6+YfTwzCcP4RG1JE3bf1Gh3z
1DsfczSey4WSkGvytzY5rUzIs+za5qUmRtT+shKiXPaXVXSHky9dsnOvjhsi
ZtfyDS8G27OObAgRAE/A7VXQb8BeQS58RwhlP6aWB7zjfwy49A+/cvs6jL6R
xLotiQOAOu6vwZWjhSX7atlEl8Zqwmy2N9bJPsMyA5EVlBH9BoxmMb7O1zWn
pXb+Xi1W9rrqFwpB3Kb9c4ffCZjp6Pv4sg+f744dc9W2Em41s8IF4/OUiCOj
8uNjgMxUklyCmp+Q4SYwIm/V/zdozg/ljNzeKNEP03dsPLFC9GdiuZ10YYs+
ji2mSaQQsTvTBnREnptNnYKTsMpEA80+xRZZmnpggoY1wuSrM62uGIMPYfDW
ybU1L67n5yKmtZlaUKiWPuoXIM4U5dWX2KsCCL8UTz9B7xWPGnJG+TO1xtym
dn8AN6lNGnS7MyMIoFzt64tPkT5AzeGm8bfw9ZqMh2ljC4h4x0U50SlIDUdQ
LGRwmAk8/IsVHJKERs6p/f6sIxToFN3ycHnrVKl9j6brLzzcPzweviyy2bI1
rkxwgRAzJz94/7t+pKtpfPxAh/Tr3vaq1530va/Y2kSCjcvHZyclF18dAwkD
B2gkMDTOU+jrzb59vTU+m8c1roIlXE/1uJ+67CyVOtg70BGxBQVyVMpTSJb2
KDQNXqz+mV+EygwScA6I69aLqrWYFenzCX83Whez+C205WuDJe836/Fx2WIh
ZLnWFUk1UGjF/N0Kajj8G3j/4X4IRqLTRGOMCZ46TKqL2lNcwYAEIaiAVzwG
ifrdEXe+5k/3iw56+v4sO79cktW5QKODq7ZIfKXytNMjQnT/mX6lkSst/yQE
LsKVGIC/18mxjwmCmcgVOyuo+4CNus1SFyKcD2ym1zy/Xnu+Gcrq/Vn0nv23
CwCLHRpS6eUb6Om2H4x4h+qdbT/VxvikfPqXG8SOFpsUlIi4PivFUKxmVDub
69KN8CcgAq1h5w4JJurSFrJQuBJk/pqHuKKidRHyoNUf97zDfc09K2X7DVaC
6ovjLXKUojk5LR9Iwy5p9E72/nXrQ8Pb4gtG5NKFB2a6qwmhqC69HuVpyo32
8MEfMOk6sPcSeq1uDyPPGL27L5soX5UYZFL1U3ejELHNs2rsSNFCQ3+P7Z5E
8KOEvjgwAiTh/nXKYCXD06FSpeUYYtA6jLw02iPrB6jgETDhF/OgfycdCwQv
KC07N2a2e23pvjeVizkcR8V6n0a76/Y00dK4MBZwzk+C7tXfF5bXGzMLvDUG
0LyxRjI5FcrI5W6yoilF679/r6D0C3cDKCy/URY7xIQgA9I3NUU5+0iiba7K
8h32/+kENaEGMkbH6rN4KYsO/Fu9rlyQTJLGBE8+DaCmbACbCtFMFCWE/2Ek
w8utZ3wW+yPDqk/yKaZUZjgAQz28mkI1a3gAU+CD8GcZ3X9Ufd8IghoNk4Kc
hwGIN6OtWZPpXmXaNYIq4/DMZmUt2Lt7fV5eKf0We3qRe72CKRoLzQa8IPIe
cEqIlCLMDr2+YHnAO9zv6mRkyiF+g6ElcOICD3HqeZNSu2Jc5PF1mugMOk6P
4bkGtDyHAuFaWg06ot28IOrLegMM0ZoWMXkrCZziTyeyTVXhJ7NFOEX7ZVWT
0nMc6LYVeuucHSrOzboPft9LkO+G2l3Ps9KfHd+jD9nyxzpO1ViVxHBccULu
1WWR4UyvVn0w+0fkWWNhCAddC4VswFdFb+Ek15iBHiijeKnEDDt/sGHgDlfm
igmM8zlJrLFbyOhqIcUbRF2GmKTU4STs8r6AH3WLRU+Z+U7LFX5h5EucA8NO
k/ZMaJe76eoUic2HLcRJd06+ziS9UEieBXRxDONw6S/Rm5r7rFcI4gyNtvLy
QRyiqbID+bxhifkOzTCYP4blMNVJhHKpe7UpWYK9g6s+P3CoymDHZ7OjG+tO
ZYG6T591hygsaef+3GqmPj/7KJq6du/oEujMxjrGW+SAmZ0LpgJz9ofDbCmm
+rKWY3NiH+KUSxhY5C7UhIpLQZcl2o+Y2HnPF6dbGBCdRDCwH7+Ey58BNDZ+
n4cJV9WpkThoEf6Kcfm8nohWqVV4QlGQ9d4K4+xBFolP84g2z2ZPKD+ZeArI
s7o0PXB0qK9AcRCMN/Xf/LLnM5r+B5F/jM2li18ETxDX3+yg2WwnSk5+Notp
MfIzki9YnKlpZ54Suif9D28aJmOzquZKzYkQVK9KhnIBorPKPyuI91riQyov
CCgPwBSMxPqVgEGoXF3PLKzfcjn6e5nMvc36YiZwHSjhcbGXTqoSCPqUUZSK
TyIzpgA52IW1KTaLaVHq6le9ShpKADRBhQp+RG3pxTXcAjY6IXPfZeIsu0JS
xBLLzrIUcGkGFPacSZoWR9uqQc5spXX7tutgD+8A9+tXYquN/oM8BOQvDVnG
HOKz0T9ObzNPyQYZdJDfM4FKgnTp2IvJkmnotg5L1mpgJcVltrW+glOITbOu
6dMn8o03P1HqCGVGF0L7EHFFn4j/SqmkXEA3zenW0tJCDM+2UlgW5/HnGOJR
7ubiw5dOQDS5EJaOgdYRCX+HrxOMVBPtlrUiOmy/xFO2/11m2eeIOm4KnZkg
iUEsweQgP2YjAv5qE1ZK1Twd4jTSIvn4rdcgY3+v2GqBueXLR3YykQzcbZZX
Q8YcYaIMCX5lJ3OxkUWdmBMtv869VYeD+Q0wTbDFevHignI+NdP17anKN24a
rjLSC+6GAG/9Jz28Mz+p1UetRd+Yj/FbPfuOC/fUXZYjV2q6SKwaCM/5oIF+
N1g6QdWUiivJmF+gWBCEZz3RogAt3zQvTF4B8r9Ok905HU+6ELwnIek7NlTS
zdsZhC1OYNAfQFxcsjJoHv4VgzWREEEgVpW2Erwe7ExAb+xxWVG4qUIJFJoZ
b3rFZS7sxqU25o1IjP9zp7FvBaY+m5usVrjU0T5VpSG/iOXYHZJ+3z1MtO4X
tz8jnocv3sLISHJ6UwjiMs2jHoJ7U3CjLDMftkqOl/nphO1cqB8BtFc3fpOS
eEzfUM80feOn02vSYZ8OPWL9ggvW3dyvD39lOULcclsYECQIl7IjgFDJwTQr
0DwspFbDZ68eeDKmgYQua4D88UY6CJPDO2SKtJk63u4uqmh5gSd9JnnOPNn7
HUvtcpOkkgbbHK3vVLhWAd4yHGHAWAZbx6YBKOaBpz68tU14mbwZXSCbqW8H
XAaFpaeP3efCiBBZOsqOSpmUUbcUzvOCuxfgi5XZRvJqfMKl4VXKdLTAWkkc
0NdI74MPB5JzIa0365m3jnp6n/GjpxOuqU96rreDHneRk4Jsmctq404Lskby
Js2tWrOYRPf72N4J8uohIW4GvwjtWUpXZXqKQ2YuMnSacN3CnQ1aIrilEdCf
GqzawgBxJ6qjpjiKhMvVmbNcPQVdn0WIPlG5hSpDNfxwodPiuR1o+5I5nQ0Z
704/NkZC/heLD8DAdpmp+Jip55Nifsk1buMMSv0WEAtkw1+3DRr78HowXCKA
XjA28IHzWk2+lnhVwxP59W3KbT4HrZQbdHlDne+JWj9BaAfBaXvygEl9w0RL
D3VhINeQXCfCl5YwCmIZ1E0H4DKpG7g2/ooPe7fIiRhq6TgslwujvXhGqEzL
e2T6uwXwRUjn1t80whRBJSd9F1gTHqlThuM/oH107Wjaz9uv1zlyEYHyFX3k
oZ3lpwDovV17c8f7m2qkRdoelC81umEqBJ3tEnRWP8xFYHhERIaKWTn+4Ny2
InBwJOEo4gnd2jl/iQ57cVyPz5XeKe5E5b+7mf6hLdtjsj/lfXw/dHmSf1VN
aYf5EF8/sbwZ5Ar3BBYNkuh2jXtvzGqH4UITe6X9DZH07l3k2DsxSGoJ7+JY
o14LKzczTGP+ABUW/VEyAkts/AdlSWBUZd1/OUM4KzZ483Kbv2t5GD/2P7zE
VwhHZFTagUo6R0wypIaoGPQ3lHok4eG9D1ljLal+/Pw7KtdjBzkGkjQ/lWe8
TljWDCW8UByzpaB4pjYjBdDTLjLqQhv4U1QQkUEMPweGzb+/GVwWWANZ086O
OHRUkuZxH+hcxPCoCV+P1eEwe2/gx6mBSkafGXnPvqOZLLhrr8lKHj2K+WA5
oTWNJ29zAN3iVcurqdL1WVFeOnDuNWounbhdm5SE67fWhidaF6alEh0t1gSz
usk+e+tkKg69MqZZh/rB2NISesrbeehhzVFO9xj60d7F+pEQrUNvaTjDt5Z0
bpu15JF/a3F2eOFerKCYEh5TPlBVXxAktfqxjj2/nIcpUxCahtZIVcmZVhmM
pyq3vu/CAZoY5wpWlAI136zjwr/HFdPFBW2FuiQSOaJG5vq3m/P7eTx40QXQ
x38rE1y3reqXfbokDDFjadAOaURhiGl5fkQtp/ysFAYXzPMw1bbSI6jL+R1y
0mFpelnLFcu/9AmsjcWVQaO3Dly5RuuqnJDACHwVi8hsVWM9rdZOnWJ8rgxu
d6qihbOSVGP9gPTPmrx/JvBhsdZ0wvaU8npu4kMiA4SuruMhIC/9/ypaobVp
a9puRGfy/UB2t+6HCKCjynYAI4Gp9Tm4XCCabMi+EBjjjuY1kdX6eI7TkdSj
TDdsOK/8huIXyETESn2X2x7DGUMxzRk7MAsv+v5sq3NCpGr8oZ1tmoswUb0Y
h3Yrx0wGVcDZYwc9jcsbvzpNexl+kURZwXWRYocMfAW2Z4Uxb5Qt+D3dQM/h
Sejs+UCAS4rzA6oQs5OrVTgyQo+lOE9ZWjIyRV7D60xwiXU4K1qt34y5eiPR
f0LtNJv1T2RRq5GFZ9lyEbaig41/CuI1hRiHX3V4Azqbr08EztCcWIzi48yd
g5V3Duala7UelOYBFJ9qDr1fU247Ef/tVaDfzHRtPSfKLoeF5s4VX5PnE5mO
I9ZEUH/ywgQRUMhvqFBPQcR5VyvzMLql4FsKvbHCUFdB0WbJhTc1dRlyE1Co
UD6pV0jTDnjDn2t+eybLjefqc/cEt2c8iw6yaCFf8LGj7zvaspY3yhx7+pmD
x3Ek++XB4A42kqzvrODGQaVxRL4ZXm16t+sO8Uqpec1fYCAycy8MQzEsIelF
tSc+LjmqUGWO2Jlcc3oJRUQFAcy99HEGNauddJdSsgXmuASWqDfutHzbJZ2N
l9xSmIStjYWw2JFPUo+eEpB6t6p6LtttE0VHqWKX43CtFT9uO1Yut9tu8KLY
ppJTqSOqqCNTaEJxv5LiBY2WO4+nFp7QSub8Yp4QZurauhBL3BAh8/b1Jqsy
jjVjYIQEBNXflb+gNJYNJn5GkjHkDz5nVyWYbbjHliUvJXi/Ya066GiXoUZm
B9e0iWbNtQPymQUcbDAu4SGkCSmLNILOTeWdh+Uu5IYLqM15QDEHFjDSrA4w
hzibE7aZTcxUfo6UW4xN/bIWJcJcsiO8RQj/DgjNsc7aAOsMuAPMPG8TjVNT
qpHeV5FGYpBboc7KcolOq54dsl398GXvdbR02IA7DWw0W/XP/7PdvLAzxkf7
wIDGZDGPADb4zhO8/oWBx+hrXm1V3gyA362p/mCWWiA7FJ+Y7GSrEnjsT93E
BpZX3TZl7Ck4TPQII6XxhHXc3mVe5l8SHq1WGujT3K2JTkMv4U8UIszsB+lu
t87lEu4V8S3G3WSSo5IoxbgZWmZ2ItsxuwfJTCGkm/gQkws0OVzmIeTGktb5
VAKqyAWtGDvyGYEfZFBfuEzihQPgT3ys7WwZaUXYp0P81nvyndTz5zDhV/Dr
/NtIvfqkklriTAH2QZvu09Ri1/lCwgxajQoal8JPGrJt6tx+N07+WgqfrBTl
q+mhlvtNfW70dpA3vgYAGD009NfCb1asGcaE0qTqGKUiAJ4UE9Z8XoeFOz5D
7xmcYzScbCk+V/E2CYVnaN0pQBhO9p1Q/O8CMCifRLbDyR4SVnRkzRs5F47W
krJgs2i4Z1iLWRpbdIdCv54nBMr3LBQQwR67MAYBxhyxWTQnrqTXg36hd+WA
ltE9a9DzTCkMogvHmZ+8k2Dd2yf03+g+1a7tiGeFxKBIP0SLKavT01FDURMD
itJ9V8+c7/moYAze33qfBSZC/wiQDuR/tTmiUcJyp25FMDo0KR9zQb67y78a
9HTLU50OtrNeqr9R5W5LVdv4dHXzgogmrZLLyk0u+bdF44AbLcTuW6vtVK1y
7FOTnb4XXnNvffFBDgvRVv3Ium6U2Hrslsj9uW+EFkVCaD6QJY98+SE+D/da
KJwHtVzSG5aqgNtW01hsjdZux+TvXHiGORDKHsgYbgPNYLTWomJqJDJdY63V
RGGg6lA1lPfeaxn3R90X42VPepQcr+CNjv39eMiu53skOQWgMKndQcZ7pDoc
k2E0sk8Lffg7EGSQ6AdgS3JrG8O2KKp3gGoniL2SveU/SB9IZLzOB9Xv+62X
1vFNyXcZjZDtmzfw8ogrEnlrcjcJz3XbO5HhPSLtaGZss5shjS2IYmEVVYTh
Taxjr74YzPS3uFWM6scIsbObVBMy0tY+DbSXb+R4TEb4AnuSShBQs09dgHFV
/le89wL/cnOhxEjkhLfTxhDDHxPpl8Z3WB65ji0BMgCxjU+1svuKWGXH9AdT
UDWMD1VXmVALyBa89uwnZW3397vj4FDlGVwPMeP1NuS4cD3e99UgRhn0bCkJ
HoS1e+yWprQD2/tHFT92N1ycoCapMGta13tPMWstYmFZSoVTEVzLEu03uk5B
4Ft9J9DsDgrZ5suoABBhRIhKBqWBJpHrIXB401BHWVdZ0Y/0YVbMqhd7ZnWE
sPldaAwtrb1A1kXA0MSZozdod7Y6eb5Zqs6AFatp1uBDKe4fKr1X45fUx7/K
Ak1MGIJjkTxSrI3NW3m37kT7sI4OPGjXh72WeH65eOQJyzxbi2NvS2IEBCQ4
kO31e9VNU1es+9F31o1ZLUhqshqr74LHvSJEA6CI3t0+8kXGk/LY+O6cTj6h
dDOaCCWdLXU7Muuf/YGzkBFOyxBrahQoCj/AtjnLRUM0hQxgWB7WlwNhQLuc
34f7ksjmUWPJYuM7ZuPXgk8B2pGI4ttKF06PrHGh76H1nIidj7x0CVHlAhOM
q+LkHM33DhTkPNQKvM+65mHYSIpRq1iCo033RAwP1QJryNVUsukPNny2Xjtw
SZpk+GvctZ+xuX+/CEGsvffTEUdcL3CG6rU4OyeKfpn4X8cmvR5miIkIWmiY
fXNJ0kRJT1VXd71+rrvjrOTGuaHosJCMN7mLE3k5YMe9Lo9zPa/vIl1VLfEa
WMzE8HHBJROjgl3UsgVEAGR3d7XKbRJUqrMFIGQ0M7QnI98GjqZ5jjFIPEQz
2kzZVW6xq9ivAGXeltH6irXxYy4jSjKgbGDGGGQ4FAPHXjlkARtFVxvdIdQy
fbPVEWGgbAZSRhJYBMHI3WDnARs73GrbHc9+PlwFCOQ8aBnrQcK66HzCS7Hr
68VDXRA8ntMeDxyYC0e++F3KtAoosE6jcyWT+XHJHmQ9u6e5IMENPbPexpIw
cBybtQMF0mpesOH/KS9LmYpMQi+bEz5kABh0wZxewGqirREFIn3mx8+BE4Hr
KH628yLCIbzyIxJPDni4sD3HLrI0CRvk0bYTcdARl+rwKpXr8wRhW3JXyuJX
pgQ5S3RsJ03sJL7wOCHzGxgpaRNZdW0c7MCTbLC0hbx4a6JY8dElwCFo8nnk
GXvPixEoHTiqEE/SmZHoKeU9ukQWgcJO6ywz3DFgrpI0TxrPVAcGW2uo0PBe
M73igpT+Fhj6CLQTbX5NnQYvB3zPYKXSQakEV2Ii7nabmy6PeorHF4PU7bh5
SVQVri2T5HXXtOLi1qXHogcbdAJi/abviHzRJ+MiwtuNwXuV9E5w7klyVCSv
Yq8uept31PZ9jx3A8FBZLRhTbJKq3bUMgwovOTTq8+dATt1KLgt2XSF5x/nZ
BXSB04N+Xo7Wz2NE+RLLhVDrala1MInnR+6PIwBzwnmjHg2axh/nUObM1KD0
RJ2vjkEGbG06qHlpoaXRZfZt/ofbRUDBxiRVtRivsRnwF9E/REBckTBsUlMi
kFI1pbOZVySXYLwRzDwHameNUJyqNLHsQzkq/jYzJB64tPR7kMjz2tPsKWjW
cjgx2KYDOm3U5X/IaNd9zXousi+V/gXZQWaU4D80Ex1l1r1k4VoUUZrnos4K
lc2A67Ji9CHrVIXy5IYmOtWz8igI7zlPF35CXrEu2xcfqlC4J2mDd/Xr+O1P
LBHlRxmEQBPsBBFQvQiFUvsAFgO/fZXJa53ogrUTB97O4rM9/NY3jUO4hkof
LgYDIZesDbOSOQz2LQqlg8EUCM4p3YgACprKFs5aOuO/x3Tm7Vm5WCvFobmi
ao9zZCGai5mnM6nzl05QZki3qdj3SgP/GxXyXXpYgVdT4sc6spy0/kquCRxn
vSndPw3fzqF1TVB7+RJrFREJvr4g2EioHoG5OgCNJJI3hY3v0vF83cPVm5t8
JjfEUqipsj+n8Blp1ryQxX01hQ2HNTtfCwX/Gl8C7++pDAkzxQMOMLDpTZG0
/aBe+LuSh0qqQKzeynpNMta1OqqNORsHTfPLbFtT7KshPV5fpE7gJNSOtK7A
aWy1HICQ8V67a0D/uz6/qTMTxMRNg1ef2NNfppvcEKzEhD9ucHdzCIJe1Snu
l9zvrRO7Vnmc78psri+CfLGAlLvCKjwtCT43xM3gB6lrcuYCLMg6BAWaKpn6
S/uRlr6ABimSG6Q4Q2AasuNhxif7jP3m82q0tPsTU+sKLhCXksrflY2/t7GS
ocSFJswDgaK9gmtnWd2I1nearbreq9nGbKiP0WQxB5v5rnJs/C5U07PmQ6Qu
/KzCPKV/lMXTWWPBE1U01QegM07Klwu46QAkV+gYegZEQWdTgDPuUnrBUfxQ
63/RthyG7KcNJm4pc/U6UeH3nk4XeVTLSJ4eZyxkRmwVNPzSilpghZ/hgX5r
UE94NhKjbg8HLxhx9FMzKgZpB7FbIe3bDt9GGdoGyEM3Soi9YMy8qxED4iM4
MN3KtYhxvd0XaW4q+ZkUQ2bCnBp4V8xkN50mytPOo0cFpZNzOwOA58/xyoHf
69ed0HV6AYUrUxXCT1UJ6NKSvGeOh3wcLrhHCrHVCs4rw0zEcm2D8KiVKkDj
sQJn6KtNZhk93CtBD/NpXEo5XFSyByg7UaA+WP9Y/8rbSwLSX1s2WTK4+hHc
JdMNQkymCMJaXbOOyneFOBriHN80wvRUc0ismip1RPwU56z0ZKBu2Tx+tcmW
zw7XixZjQei1cdOiOzgk0JT0ht1xnnXVORIU5dm5jajTPPJQ1MWuGbOzWidq
eZ1xeYYf1aF1/q5vuuzh19b7plTSeSN+HIf/PXB2VZznNnfcewYqzxaYl5kk
6oVQdEtkGpZE1lg4zV62B9RVwz2K1bBhjJTOOvfWdqYLZrGh/G1eieGHj49G
L3AAG34YdE7ab8kXeUEnhLDQoaQYS+thCbRPlLrZw77HtGmhi7F+9SGNpqh4
7IIVbNoPtWTFJ3YicI26bf2M9lAmxtT/do3XQLhO9+vNzM2ZGqrFoJxhxJMh
9OYoQVleeI3mwZMXcjU60a3/DZyklxb+ZQa2+xs8nm1XMTP8lyfrOKDPAeHF
mcTbsKXSfPhTtXzsY1W2eetyQEhkmj9oG4TG4M8N3F/MW6wyXPZ/pNGZaErt
XWshqksQo/59JlWXn2cwhZe5qDNQnREZiuF1lHCr0UBi1YuDbZfSM90VvIxn
MCJlh8HDHyp/WPdVe3T62GGUbsoUHmJTj09+hGIGLP0mOVjAyaW/5pHYyYYT
MXiAQ8BcsdnGTnb0oMCm1VrmsfhjbTS6vlN8kKiDJV8RskRSLfu4xjPcpcoi
oMuLSgHKLRgRAvTA1qgBH1pPBjwLvijRoQqFyHk5snXEQiaR1tazp8c9iu1M
MH0dy5LY/dS4JLChg4Piup1AFgGdpKj/W3C+mn2n+3EijL/Sss1ecR6is1fG
yG7fhJhjMAbsMgGzE+D05IVTLrlrqlpPf0QfEUeVqzhswQZCr/+pYZ0UrXn2
iyPzxkSayByUMujFxv+r8o9+45K5wf3wNe2r90u8OdcEWS8riPQ7HNVKuV2X
8YhdrVz5e8KyB4FqtOk5wFVGPScEsQ4qycFDWo0iNCn5f6jCASCgUfHsw88i
zBPFAYv251E6uass8XBOzvZqze6SAQcRCdDD3+cqvAgjDfsnQdreGL7ig+SK
xbJD53SuWuhlvI8fQeBQXuiXGSv5VbCTU/dTQ7QMt+NMkncPwE+rxLDsZd6r
/Pf6CSllpvyW71fwKeZ3455XaxsZBiFPk/JvLwRd+bqyF0LBV0AeQIGzk6P4
CcqUyISI1eGJABZeWKnO9bygcGdK6WGHAO5fjTt4XBSbsqRWmQrtG7FIONt1
FfP6d1WaRsEJPjuSHN77Jj5Swc8kn7ZXAeqVrdPN2srU6f4WPjHIaOkyEV3a
fsBjld7L2aklb36cdN6N9qH1kcyV/v1WlQjo1FtDYzyMuGII+5lmgw61poxH
Zp92MduIcE3Klcmkxpdb5CnzuikkpxRLqRkbHJoARW1je5csS0sIbY/zvOd6
9WcRFi2JZRAYFIKK6PgC/igFuqwtYyqidQpTD10Hw3SEvwVZcUEqSDS7Zt6h
EF3T18VOSdlpFGPbKMkZceD/cnz/o/wLlhleJqHwTw7Ywz6luTaHhDsCyVC4
GAyuwDosuKWjdUXMZj04+NxPD6HDiAuGbyX7AlZ09ppTyoqFH5AoPoQ80qDy
pWr6dEtSpTXAQBfNspv/mxUiG01oQSm0WtGcv85dkKSE3Nswuq1jzwLiWPVY
IazuTTcqZtLc3wMXEOQwqwkkvd5GQ87xykp7NFFEuwx7DYtSyCWpTuxr5ARd
Q0GZPcav5i9Xdwbhvt3bsOXgNksmx/iQ3uwCbtgY5hkGBdP8EaIt1UABN6KY
oNKh6gNZhI7DiaI++1NjRSVPLh/mmPLqFn/T8tyemDyuBIbDK6lTs/bJMY08
zadYXl/2Xc4/mr3QhePmsdGWOyOL/VxIA+YE3YBDuIwz1JilBTr2b7uQZ/HX
hfhzv1PswQcMl/ezGP9TJinuQlVDcxcxSI7RZXDF5saHqTf/a5q86Sflh1zO
66pTbYKPynmr1G8DcdQ0bQI+W/FnhLLtNS8C1SpUMyZ0iD4QtlW33oyf3zOY
wO3pX7rMrVnN3kloM7E3Ky6cZoKmZixHnTT6+ioYxFuwInWEfc11fvTgNxiy
GM1LB1DusRo2sjBmyhqNu0BEzgNjJ3Dgf8+tcnb0K9ZoQg4MRoBkL52BlNep
J7EUUN/43Sh6yHQq4V5ogvRuPVScT6ztGbf5UfWUV3MQ2amnJ4AZEG2Wpcfa
y/cMCM/Ir3xXsg+X7z2a0cWWSjV7F1d2vqwcPtEfo2fwC95owjnzPGI1qz1i
AxFGZ5BIKvgRLC5GJ0IylseQ9+ym289FB7/yQMvur0nsBUZ2aIorEnEK+uw8
6FqE2hcZkWBjvp94XexUEHCTvaUFMPiJhst5DZYI5nlbhnheMouDIsmYF8wh
60k36TaaKcLqUCJSvyKp5eAtK6h8/2SCtztUy9S/n5ROMpmoRpX+P8uFDHVw
n0ErBLaqwqAm0nLpqH+67mVzTZgS800A6ffx0EyLtw1/QViqcz1SIPq0Qni3
/77S0j5/trXEozyqKnnVkXVkS9LPP3BkWVh+reeYkL4jdVGxAdGMOv7ZL5Sy
TsRFUuk2vQw36cfLfXTqB9V9HxuUgZkFvMrpv1+DhRdHIfftJixVcxF61jZo
DCo12VKMHVuHWKEOXFk4WtZz9l7EZVahsDMAH+n0yBc/Vr2C9OUUVJQ9q50w
QtVhamowHINZAAgUc73RViJgiAZRG6JL/BiAZqE1ORnZ3JS003QdeG+WzkLN
UG/Bg1XN96F2Up8A7xqKfm6xat7Zx9iWY1gxEDdPbOmE0lzligieKMgO6ABy
8cDuoshK0ifeZm6NO7tr0jOgLBAophf5nVadr7q1bBvehhwhUGQqRzrcOFcI
IK2IK/lvbuXflApC8WIH2D2IaY2oH7yxD+Rp+EUBOeR8moc/eoByA7RQsOji
ennc91l7AtvIhbhF1b1ToidmJ256yIBSAcTbqtpnuAuVD1YuaXUuw46IKlH2
4bjpBF+nz5IpIdlsXsyZNwFVb9h0dJZfXBOYzjrBlfmi0vYPJ4xNM0BvURBm
yo8PGwVgm4DDYif0Ti0BYPz+0OwEgolUGSJk1FGMvtn1JFeKNj2Zv9r8791o
uJ8KcsWvtCcUJusHjw9m30KnhWgJpVZUKrcfPvHAjLfVKvbbHS6lLwFPh9+Z
jUHbyBDd5Io98IPdWqSbgnP5ICny00YT2thw5cOQ/E1U6hTp30TkIamKVDOm
EAjSZP2cIcRkEWOIzpKWhLJ281KSkiJwfokMLo9mmrdvJXD7H8xjwg2TW25K
144aikZwnx5QKKIZyrJ/dQEMToVLyVqphzyMuaFpJlW8+KlT1+EZfFdlpe5u
vdCqWLexPPFtH07SvWrO/AEBYxfuywmhuCM2lhbFm2Fz3HVfzjhhmnOoyFf5
bgvWpGgBXhHhnkQUwG/fLe2qIs+1ReSMTKutV8/giZfQ6K2gtPEq5aC4g9LO
hXoJfudol7FCxtyOrGE0e9TZkUVlysijqFrjUBXou8ZJTY6zxKKmkr9pEtkX
LxZFBkyXr9UGA1+s9jyJ7rtGR1ArmjlIEoKQTmCl/HLMHPQqQD7jga+yEhtK
wLFcwOT1x1PoRolsuAPBY4lPghwybeXdUFS3IPapt5RDnh9Bz6sJ8KE3pBHw
nTmCoVl5gvymiwWkWAsHBWT/oLZaaWjW12XnegrRd9j50oWcRhf3MSD7hGf3
8mcAaB8qteubATl/vRxFl4AHfCt3qhDT/P4tZE7CmZ1/8cGG5hHZTXK4FKak
YOCbacaxZAS9dp+IgRC2oSqULaUBXq7Gu5cjIeJ3Y57Dy4fL8EkTnENoPvgQ
qe76tfrYAqGTOyFltqo/qcWNr4iLyIWDBtUS56t+89o4eier6Haha7ys7gB7
U1voK4lUcDkc8q5wgS/5txJgFDs4rcRPef5b4hc+8IJZxISCUSb8rzh8y6yn
HxUyEkRfGrMOEs578wO5kmWDmtJUZqSgbuHdDMunMjy81JlqJPH2N59/lOUI
Z41p9cuVfxtdV4cSVYaexvIppfvKmFW0XSCLVfZsxGIoY5kxuDq9VkyuHAC6
Qslh6pEByv5hSP1m3VYGuGq9Jho7/rRJLfglCdjLzhxtsKLzr2mezFhzbXDj
PNrASZ/H7EISWpozUjy4wdISC2JBXp5VcaXiIT1Bt7uKWr9AjRDzgPrvbeu6
YGST/1vUFY51TQ/ZqTx5xIcXndjism9MnBggKc6HMBYmVagSmZPlq8ovnjZJ
3QBnl2RWlcgblDYob4cHExry3oN1KrtsxL6Mvcxc0Q+FvM9xJEPt1sq2N2yu
CEOd9aQfCtzw6CcE0uipBFp2ym/4VqoNVs2rOHm+JxSCpaRvcoenchU/sCfm
KNRnTcX2QDteZ3eNVNne8zwZg43cqy0OjuT5UUfCKoABylaarqbRLgyq0bJo
VBEhqUgG27aNPyPVCsSxFOroAjCWzEgbAAdNmkeVPeQqMgXK4iQR8loW6RXG
cYmOCFSlG/qVnNYkxsdMgjbBZP8iFrG0tGVUddcSEy8jfpcRuPTuUsESpzuB
BaD/awlThlFlprSIsTqKRWRKQG1yii/GWtrJ/PrZH4rMnGqgDa66AezhyjJk
kVSXGgsn+99NHrRlqRRMI5SPu4t6rcW+PYEkAcAZXuI/JufE2hKJG+6FqKdX
CBYDYNTnrdLSKW2JQQHWzoNqHD9FtTjHlG6gelR/TC+7qN1ZrygKyNoqNiTl
9pBUiegGTtH/tptiVCdhwjZoCk6/PdG6eXaWi2sJ0Y8wiMWoRKDobyzaNc9A
W8mnd2Q8kdPPp/6Q7W5jTiTYZCiDLmjOCXSjE36y2mG3R2BRrhAK9nm6L52m
3Q41T2hvm+hQwLFIS73MKGHoxW5w54eqDwnd2sLb9/LsRvIfw4FtgfW7syrL
8jHob5SWCyDLUcG4HEB6JlroJmztlk+jvgbTyI32+iXv2IQHTAYPPJvmuUHp
6PmsF8fEsL6MYTvJhbZBd9fuYRDAiUBN5wIKiX/xL5dWIbNB5vx3WStidXaE
u2CxBxlJjiS6Zp/2cNvWO9Wp6+49zLsu9wDv8UMKdKWVjXuTNRmJlK1RwOvv
ogF7PiVUS9V8hDenpQsdw73P6hpclqGaSrH8hVA9gB9S2ofQKiWLKx4Czmts
oi4bY89x6n7DGtAiCl3UuD5WSYGZMlspHm17xbdLGeDkOcPwXqxpVAz+Fb6l
YJRUE4zNitQboY6xHsfvddvUVNxzYridThDp8i09OqT5f0XIy2thyPLJXWVJ
A4zWFPQ7UL04N2nKICQvwxYPsEkWErApAjkzsPTYuiyvpTQjpSFHutiIX2sa
+5LhG45+3KfO2j1zDorSoVJkDVMzBGxDGd2jjbuLJl8TdxO9pt9dKfSjaNbH
xpJfEPgC5tDO9yAVmJ8RMYEfBWHYSSyDoy1wqFLfx887u5fheNZ6U6IvxcUE
AShk1KHa5rmvNvyeXEuh6JyXarbcVSr4fs6axKPaDcz4F1jXeJ5FbdBFfKpx
kxudDJhXMezLgkZAGAhGDyDgWseHzgj+M5BkyRVSTV9pcf5+Jpzmg94v+vqt
2+WS3nopcN9mz0KJ19HpYG7MGxGPdjhkXQXht1KWjULsVAeEDYeM1gRnWi+d
1tL4EXBho5DUGcYYvj2lQY3ZTWH0+os9eHOsk5Z7sMwpXakGIdDlXX7hLHKi
t8HQyWgxNujJM9welVosvOPPrpJ3PjSucFzmY2TC0+KeBtefwpAHS4l4MrBD
JfF+7aMiS4Klt21An0X/Wia9+foHKpQ/iHwSXbDnG1DlKc54UXlxg6nZl0pi
A3zWS6BxB7t7PkHvlWhOUkEyATrTcrwSZylHNoru9wvDVxrSXu9BZppbAMI1
H/k4qV+n86tpa5HV3Ua3CD2Ewi5MarWV/RidUjMdtZkhtrJREXNi5BrUpTRO
E3jveiH0s+0RciVI+flKVTg9qh3V7Uwjn/SA8ZCIzBDrjjAHWJceeQPizMN+
UEdzrIgL6p+6ktzF3LuijMcSbKGOdrmA6N2OQN/iIcCI55DZVjy6JfC1g5FK
I616/pxq1e4jdjxHEiA4DNcVQ3DIHWDHo+7RFQGpgm5W/Akr/h+2qHGPNNC5
F3+sN7WeWJ/HBgA4HJ8azUAwRvFvl69kfgl9j/ZbUMcMqKO/OkjblRxleuRo
4XYLwsqvDo91o4NlZT+enee1GpfM3y/b8qJ7dBHThcMMXBwGnpMpJJULz87n
XD3OEHf6ElsbD4BdiKtDYJ1LJba5g/QGjeqZtxp5J6XEzDWbQYD9SRQMCVAQ
6bDWuGMt2m8h6p+cVhZavMt8N9mX1WcIz+kCpsglN68WBEZ/Vf0Uq5P7awK5
ssw2rX8TzPPjNSWLb5KF94D+YMfm1jIcox6lWM1nEeYLlXcLpP5lfEid1qzi
YuEoN4j0FG0XKBA+Ahh6ltLqRH0494c9b3vcQ/dsur7g31Lz19ZRnUFntgwj
u6GuTetdaYa1pnrkA+y+rMz9NyAHlaP1Qvl0977+YDW9uKFXR6YAfU5pQvr9
WvXq9HZb9o6LvF4lyZQI4mtTpywzdDlANnWQf6cH/S2JrNUOhbq7zhqoROTb
VgvBWM1yeeRk8ddhR1iYjfoT8SVm+op7EjtId/uiPpPcA5e1WaS2PtCAXWe7
hMzdGtlt+ScQTHfynjhN6emiCzq6WRI0a8TFKCNW7ZO7e/udKIByDyfR49UX
4NL8XChNdFBVe1YjapdnezzEjdgYcD3wvWdvkm0xr7/rjQOQ8wthr18BAke1
gxLUfyEIqO+ChcfdjHVbG503oJb/tSBfyn5NAYEjwYO4h0Xq4+XlEoVfBAzX
zTcTnWIBINVyGxCuyyVTUiNrO9YoDdYHo+Eq577+rl7oWdSte+n/QCn4sD0F
S4esi8Mj4VWIfnDnkx7YaDd+c6eJzL2Z+Dt8Mhe/YOeSYrah7xcuy+PPm6og
0bWPlYw6REofRYf20oLd+FAuE93XtsetPzHV+2lQ6iYmMvbyMA9XRJcXcVRB
xTeU37f5PnZ0hgw0+mp3QLikjaGER5U/qalRXkFMmQwObzPj1uBsR4XXlf/V
pF/0LWhoQsiQu3JoYpkZTI5EFr506YWyrxHE3tPtZW/wJFRyD476mya4zU6g
CTe02AGv9EOhcJx8Y9NUMb/XyoZ66riohx01I4V4wl7mgklOF0g1eXrKSZJU
Ft1Ip9lh1Z6ek9XJAxDcqJgiD6P0mfLLeJWjlWkNzr3sPdLFpOmOXPibRkAv
IcCVJGbe/IXsHdgDSoWfkDF0nNDcGKfJslWrl1S/ssk8XgyEhX9giKsl6KRd
Hlf9IQUcocTz+Zsu0TqL9STo3YOubUW3DtBeYF+NqTc+UIKwampVDzx5CLAK
0cBvIoriPWWRomfxL246ds6ehUaQaNFQRY3rTavIICkAEXhVTozl8penJavV
QUTrXswq/hyUOsVB4ZzS/vEc9dc5uWVww2w+v/Lt/hYiX1i+fT9pR4fPrDk8
yOxaQcewC5F1afdaDhE3hIWwbPkCqVecoQk9Jv+0+rbUOOh1KMu1QJQz4c3i
2HnjWJPoKufllazJTCiWWYRz9M4Lb9oah6fd3bGTz1CCuxTl/KoqD/AVXWqT
6n58TgLIHzJfN3b6qKU1JjsqNin6Elg9/6Cf3ZJZ8/1QgDCZ7UIgqnY5RLJe
SSd25ibXkxzuiBEesL3IW8pCqIRaxB1aqFrTk05zbS5dEKJuNg67Q3bgarQ9
HJSLO1VL6JIAkSUMkCo2/p3N+J2ofXKIGTRq5z0W8laoAeIJ3/0GkM6RfTYq
tXY6WVVvxRVnSAEO0bG90JVEd79Quox/DgOfB8oNkLdfHZop6+Ew8GPR1RjU
XLhEB3cQKD3ndQ20/veFBh8l/U4thGZudJXFaeNxgyQbb6WEuWIPlaiUCXbj
Pky13zZNj2aGuvG36Iq5sZ73sdbUKbNI7TtOINFWr6rCRYGPxokIu6KwTvuC
BiAahZBP4hbgZE/VGf0yeMjhiSsFN1/MVi2nsfEKAmxZiCR1H1RsSh0zMZdC
Tx1R23qrCoyklljDIKZThsTxA9QGMUb6mpZplW9LJZYLgbA340qAznGMdvp+
sQrDg9dVV4WRanU+AfTf+jb6tkJlIZO80atNo6nCRkG8NcUVLYMeQDX3hpO2
WAY/p1v6+pPQ0xTDbLuwj7fi6p2V01xKwj9KjUAC1+8mH/Dsn3bQCdvkB7cJ
bhc5gXgGcVQdr7BoKhgeuLJxwY0C6VexY0TERfxs3hnCYK91DA8Nb7R60Ibl
/j7TykFEhZqi7qCwxFU1JYWkkW3sR79JkXXD9AdvV1gjQjWPpEFHqt5S4rYP
5pMu7cJb7cn0c9tDfoBoK0K8HDmdkhE8UCZZXJFBqvFNozUG1rFn9Ez/aEPA
Mmtz4IVi7xC1uwmv/UWLTedFZAayvN96ajignWmjwnbuYqNig6lwibc7WHqS
zxq55kXohX4ajUjszd9Ekaym5AEcllTjIHWcnZuvGn73i4k3MyShtCCj6gZZ
BPppoeGO/GXL3Txvn64qYGEt590maxwnJdssWxFWkUgqgLeXMTjdAhQTiubs
oBAZm4y78YI7SJOUzCNElCYKRElwq9lYW67VCJbXsRh3F+8r/j/TwmcWJpfR
VcIWlHEPpJZGYypl3PCkn3VkjI2V/Rj6UITqY16XlXScL84Ixr33M3kyCevY
Nd2ldm1H/7R/RuBeyX6UcwSwY5faeMvue9UV1HpYi5tlFMhzxyNt9OgeLXOH
rXM9MbdIvJ6BOYfD6WwYRpvxemkFlr3OSgxHVIVGfBANzg6QG39Y9pnLUnGj
d77tJB3IhKoueVTQU7zHAEBZe3e0WO5hkeL/9D/Eg/7ql1/oJWi80Hv/cmNf
tINlauEcngsesg4lHf71kmGPxQA+do/8Fpb/E/m8EyTxbkZOg62LpndKq6JA
KZImXLdSng8nyimT18AMBe9oDXcD7IngcosnUUZ72O4BCoDVvk+1G95GCxGK
7uhnehGsXPOTV8tsjOz+ANxM2RqM2efTif/Mpej74ST0ruoUm4fbUphCwRTg
nKL4xOmgQ9PmklM6YDuW7rDwys8yf9auRhEG1EXVAauOXfqRU9ZzsTdj2jGs
u2Ud0UeJAfeAFM5Eq0EZHh1sFTTgjYRoBi25LkmGXM87OvhS7CbuOFDSbL97
r7RPJBQrKajLMqErIpujDoG9Nf8gdyo0egpV59LLkwi0tjw7yh7Nh6TexMZa
HeAFpY3ju5/05qzG/sVBYNmU2yHfs1a3/CClcMKmSZ649/SQUGP8HBjAunwb
LCvWeOaoxG0+cvRVDkcwClVxQAd0Ans3dAP9XOSNsC/M2VlqelUrUXzFwGEK
o3qF7CGf6FNE5q5HDXZ86DR5goMOOseON6lZ9IR/s9p3xeZvaPg8nq7oQl0J
yvFzWK7PKZVpexbnD7f2Zpk3hKNNDW1LZW+++dNs9GqCYAOLRESwNsPl9aN2
fKi8WKLHAm7PdKnST/eMmDjyTEJKJCbN1/l/2zbzMTuYgtMMjTtZfWHYzxxv
zHwJLRd/MApR0AgvTSwH7g86RgFMp1Js1oDKTd/AkYj6W00vrwe0db6qJ3fR
BSLPENUUUfZocwqB9WGyV2F3jxZUuos6eZ06nwdBU4kuyf20Pa6xyzWP+3mg
AuOErKvTnSolrWHisYR8h5Wi9qazDn4dOONUdxw6yCHXohphCAZ12Yuwd6ou
9Qlta+8kYIh2ggpt8xdhTBqarc7UE9HsQdjbmWZgIFkTSgZBg/+gqJHXb0ej
HwvMYpHW+FuLkz5qTX2zMTfbjyYy9fv9kzp2c4AsANWUOTOHn//W1zlK/6Rk
OzUYaUErr+6Z8/m0K9P3FLEn7Uea9133yOr8N2FdG5DHngSCdkKqDhQNJDGe
UbY0/nKUq0yryVl7OvtXFbxhXkO1s/5SdPquTU4lViRD5r2QBD3Zn89KqTop
UYi8LAlDW/2CfVhBbPdO1z47e2cHeBNQj71mlJ4xZY+VG+icmVnm98E0uvfF
n5jotmi2gZjPh6I8c4m0PIAn7xjztrWh8GJi1w1hNyhRbNMGfHbS4eNqM8fd
1682o9cSaEKMsClFUXzk5bo/0Y7AjNb2ZpvV++IFg0Ru23O4mHBVjiNwr/Yb
V0EpXXe5riG8j1AMyFOujPWyG81nRJX1OFNhr5ko0LrxFN6br0gA4gyvVvw1
UtHRDwOJNKwa4nRyKYzpsdxjCqPVbxlu3ShKEf+U0A0puoemOWM2XTqqrs/c
2PHS/eM4bPtPZgckt+GgUTq5Rd8jQYDAN2tjBKvW7h3JtE7qw+ahdms+pqes
Mjt3HYA+MuftzayCb1j8+1CP/OcsOVWc/roeuV9R7MeyCntHl9IA2VePkiyq
DubAzb0v37qmSIKOfDP/Q6ZZCX6dfVj6dVUQGed1RaHDZ1TVHWFdf+f4895w
J9rBMoD90k8H/HBeHp02jVujgjRkPd7ZTiESNfBu7XD1tZEpWjU0aFay/4E9
pXQxGOeAc2XUdfB+gXhNTqNsky7mx6PZo5yioPbK6F8TrlDQq6kJ52MYAVsK
nLaznG4NLE+a13ccM8+WeScaKsW8Xnc9oRsYO+G3wGaBXQ749wXUnZYD3eGe
tFhZKLjWNLeOj09b2fQMqWXpLQeN1/GhVtb/sKLp9cvQcWq3+6XMFq/O5SLl
LXPmlI6TJOTqsW54dlz0xw/VFQPLI+Q6s2huftiiGPuRrF46JYyvkAe/JEAC
LYV+O54o0pF52+6SikL3bs4sksbXKH/jnVSF1RprKUjRoGawu0c4WN7Pl8zw
/iTjUPPTkPm0B3NYzp8zwWokWgBlSa9tOXrlVFJLTo97Qs/Hig9hwxY+vtWq
wzCmZOWArpi5bgUAUBZDxZL8+2hz6NyfPaROJUe1uq5LnLzuVrrc/jQ2BkVp
CJQ8e46YqUz5Z+xxvd7XutTe7nJxHh8P+Ea82Gbi/dnKQkolkDszNT5QGk+d
ydId6fwUZ3md7OvfA8d8koWNZVyQmxYpNIaHfSIYEZLEBDqbYS9U6jcRUS2l
ARSBiU7OPXk9SiKukLtKAObYgA61YM2bay1SIYGnXhA5OLEK/njJtM0EfPNv
eQIVxi6WD805W4B2OdSpFIl3VSVrsdX1zKuzAW4GT4L8joxxplyMJEiMgqWZ
VpzyvvNW8y0JkLRHDJicmvfR6LZ6k7JBUba8b9+mLMZMGVvwxcw17L2rT9IE
eyjB2iW9wno//uFtgHWuB9/k8XDZ53xY4MHGFq5oMlGqTLJrgcLFY56OuikG
kKFf2WA6Sz0Ud7UMFIltyh1TXaf9Z/T0HHY1azAWFJj8EwVfiH6vdr4SNldj
O7QYIMZtqy18joIYEoGhxhhb9+pRzSZvrIt3EiGg4weGPmcQlCOp0hzKulJU
YCCGo3UfpuHLDCoLXxdVxfmA6/ZxhBM9zOAFgRoeR8eq+IdlKrk0us4GG/Ul
VIH4HDhwpWp7w3FSM5VE1Jz7fTjbsch0d+bF4QJ0xFyv7P3ZMD9yJs4cai5s
KLK8QLbz4F529uTxNFegG1fmbk2USsk1aceh+1Yj94733lc3SQdtGyOJGduB
O3SZhK9DckqVXjHHHqL1de9qR0dVF03yOnurqSt3RcqZbAEnWTmtnWkl+49U
NXx+z4KQA5CX4lhxzNadljJVGJ8pk4T9LLHllbQZgd/GzdOFppBDnbJPqe9a
F9nAq/iyQ9N/QU1Z2qBZwGCVv6aOSfU7M4KFnryFJaotTtSNeqrwrEzSHqvd
r1B1P+5H2GgWLXkeLbcIp+6O3qTuMmLLTwiBzsDzWqXebTFBtdyeOg1dDZSI
+6cfcSYeENz7MVt4NNK1A1FdgLvyDCCgcGC9QyZmvYMVbPwJk1JfgFFnszzm
Lc4DWbVG+Q6QHIkSapELtoM9M8dlbPRIA6a8zCJ8bTLdeYwkeEKJtT0OQU4i
tMBJIfym6aOhHc/2rQXZ27yoWbfJJt3NPhB75+K0/Oa7QqHBwwrp91N/oZTn
eI20meWeayT1VjHN37DbUrenlaJWC5+dWcTl2Jhc6X77pI3eE6BcFalJ5d7U
gEUEttPANvTGDs0/O+z/fvG94B7UUmK7VD4Ro8/V25iKAGtYOd1q6gKYLe3s
AsCWwA7rWXCuPG1R3IGO7Bmz+t61DBiM6N/4yqjDVpqyrJYm7VcZtSNns5TC
tmEJtqDqDtX+B2JTEtmnq3pCHFXKreTmnt42KLmVmRUEz82SvQ+JEJWeufrZ
X6q2peIVVk/jIgltGL4/kqbeTu84RcVe5C/pUWS7wYv4itq8ZRDir3Dl1AgF
ogun9tHU6srUWnKS4nd47CYZcezpQTQ5Lq9lHTS3PsLSWvcLBW95TclcqDQp
0WdpZJkKZu2mIQcc17qfAkN3sqGgSuOl7JZFCB/XUpPOgCmslPj9IM7FcXQW
LJiM/sUtqrgrAG7qUAmUwIGHsmsNF5DdC6sp0pkiC2BSU9x8YDmv2p9XnWcP
mi8CjW+20Dkmuv5fmq9hOnmXlxn8vbvOPEnNILFCYwr/9+fO9xgxRfKGZwVK
SAglBTeX7LDnGDixZ/0fmrjs4xrHfktXA1jw/I8agyRNAvAqT0oizZg9bS0X
L46BeEe+HMMhLsCOgAocJh4K/6Q7o5/XJ64DQaqKBCRfJpYp+kBoYMJ8ez7x
3XgZBKSMkDaiarzTaorKLJdloni3Z5NoMgyg5DOfAkMM1wXc8EmkJXQFEh5D
5mx9KdkHP+dr7u85+x4i0EVwClvYTxpOmwGxKKjosfCCE017iDr4vldJLI8V
CRlPdOgbq7Ueh4eAe1Dru166TD4BueELapnlViZevjhH7kC13YEsMJvgAcm9
mkgnBbgR16I/SfCAcPiqfGz7JEuyPeuqPAzJz6AMB7bzW3CJPmvu4fhJRf7i
s5XradGAatLjHSHlBmcwmGak3Ttkgl9UYtKzRjP4NbJsRY+jU4VO+7KllC9m
5Jmx26A3jLgPrG/ljJ2Us4Zji1bCgo/g0ZZ4zILEO33nRXIw4cfwwfw8T2dR
eKyRFK1E5K6O+ba4XruUSgIG5Q4v53WEnvdurGo58VdjXVD7z90XEvYRxcAr
jonQc+9ID+D4XDL9VWnsAf8apHGYrW942YR8aSkMOf5Fy1Ab7qL/aF0lZqzm
Rl06rk3y1LCjin7uit2JwQxafUTSipbQpFtWJDizcSSaY890ZwfVx8JExN64
d1Q9Fps4M/d4Ih8vI/QeiiryCa44SeHvzKdYjVdVAVB4dqWgPTJI6yK8wjJw
FUj1AyShRgp4Nmvkye0hXDVVWSBdPi/nDL3Nm/iqAoz05OU2Ki8YNoDVo893
BTXpNpgHeTBJ0yn7zyJmnnKu5FHXWhfjx3kvwdBuvX4r3pi9B7NlF6RKeZI8
RC6lPZUcONTAvGxvr9PCefVNJ3vhb+D1yushq5CsxlUVCUxhD3eXS1FCAW0d
zaW2N0No6wjZneR3rkjb64Qhd1gujoFUdLGYMA0Or6uQquKX+n1Dn08fsUEe
PcI86rFJ5nb4LWan9NWGiVxNbeDvaCQMjKRKD/bm73N5z3lGJJDhcELNIzHx
1+iYLlSd857wsAsWUxITRF3WrUDd41Y1/RvJbdG8n0g37nFfNPFaN17dvdGv
FETNiMwAsc1svyy6OswWyKXEYc2t2z/W8TK/gP2R01p6rGGXdBCTFzhLrYh9
jVem6bFulPNURhLbzkisciv28f547qzVaSSEtwcv9XRa5N96S15U5G0UKYAr
fx1L3DbFggu2hR6FOHWlgwhYD8cnO9MdexEN4QefFJg77oJ21zwoNxw85zBE
dkAtncHUjwkHhFA6h57BPMwqk2t6NS+yUKNOIq4cV3HjGaW5kx7phAVxJlpY
+HQ8/vNkxBVE0xEjao75g4bW9XP1X6lnJlM1guLq+3hbAE3O3G7dxc+P0jdn
oGgi0VKyGNz3S5c+N8fZZnecG6d5P68gw4NueHt2aA7H36gHpqdDgCKHuhBk
WoPhDJnAdbiEmEdeNMMnClsbWS43MDgEI5pQOqTxd9G0W5Ea66FtaV11XNV2
BkTOJiFd1UGmLSrddplJyWAFCNYQ4kg+88UfQ1LidwAHURe18YsN6zbUO/Ef
HHiGjY7Rc+uuabbO71MrEaVre3+LeCxMYi0bZ86u/3kPr5+hvPSUMiIcmgZo
xYZDNzVNYJXQeQKN+PZGsdMKFokk03Rk0rVwk7m5JbLZprKVpx8te3sgyYU8
yRpeNQi0j7e1alOqNfr1deINsjat/HLe8E0Rgkt9ligSQfdW0s1UmivyLoYu
tB00zxr8TJOXqIdi8TosaZnH2Onc2MMibkY38J3HGAQwSMIvfXkWKP94iaKG
Upzn6ILJ/Fl+oGi480tdwGZJwRREEOfhw5+c+MV7gRqZ69dVdW5yv3VSyVof
kjzpr9UCUsh/C3lo9bfR4B3SCtWu3WALnJqZml5G7jeseCszneX7rSSdezD/
QOUlTCgBWeiwqqU3vwuJAhzOpDRwoO5jxAIQ0lBGla5N64H5Lr3+DmWdHjfm
o4/W1sZ2/CuJpiDDtff0iqgXO7nCknQCtPQ/9i8Xj9HpWCUoZPgjPHJPzqdp
GfwbHWq7+0xnta+dOEw14TwY7qkT2hEbcIRVzRWSoGpuri4WAT0496Af8fQE
LjK5LZmgT2m+LcNdOJpmEG7s/LyJZ6xYxnGxhCYRgcfwLay7F7Pnj0nTIEAR
bORKhEpsndFy8UESMOl1ebGBvNai4qNd/xxxDJSf7cq5NFzm0ESn7wWFyXVC
OD8uZP/fOrRv+LR5YFngM9lq6ABJvIloTA59Tm8tSSaJke0xsEcttxD5/kCX
85Q/ITysOpTEQCjLh588RPi5zDs1RpCDIZKEIQm4bUEKk2h49RtbaHSjHKZC
dfrUvKXlkwDyauKc6Sioy5tgOWYdyZtDuFMh4QsOiNN4m3H4fmiHJyP1/1pm
vuggpSJT5/J6rA4FMWdCDr1akqn4TryWoetFWI7AnKoimXk270GXNgi/Hgjj
AlYIbbxI+PUnevHjfCZCpLkdQ0Hc7+u0rfrrDzyFNHMKJ2CmCogBL80CYug6
YGPkp8bUVCAQA+rZTMUXt2/IM1bYjEutWz1ti/SO3xXRZU01YxeqaOc77fbk
BVrRHvXyNMAP2nwLmFrpa+ibRpy0UL2HBqyLXDHrawsfm9Yvhqh5v8yCHF95
+Y+tdI2aOaM9i3bUDFD4hf7rANGQb2j43SAnEzBEFqeb/XsdkWGYDsPU9QSj
vG38P3u1zAIBM7ka3Lei/rCXWdn8f1XpgA1kotEr6jKUJQewyQOHrdCR3I6J
qT7dQtO17R3jrTuVnqtw5x66mvt7vCrj96iCn1kjmfTcChK4s3Yvwf5UJ7vJ
KvBzjzl7OVs+0rH8/UnIWFVWUs6KXhu3ITTOm+lg5+ArqMYXH93awOq9pKDb
BnaLkw8+Z4loTZLXZ8kNUAEJrZrFSV7ZCY3qRl3lpnlyaAZnxjwVj1xKB2LP
d6IoqevrQci/VvEXj6JklCYc/8aXrzoJPZSA0+fwcr6V/k/EHR/tqkWl3SeR
9oH1H8TnUVrrvS/i5hpXwvsuUZxu/DB7uQEiZSo+A7YS+q6AbVGQMC+w8cCz
DK+/gpKP4ZazWAroynKY0AwbZvQSOANFjyxOcx/TJth2UCOesfUsqZK0KqXC
NPnmid8xFpsSoPTN+H6FmJRb21jwgJsGkUVx5QIBqhpXj7XF+XFwlTIncDic
qi+sfSESK/zEcHaIGOKSP+SpshCxt2iWxHjCkVTaGPEW/Bej20mbjBobAP6t
oJIRBxWptrPi4IK3dDXbFDZps3lAiC7ifXxmT4BLtQtXR7BvOGkIHiLLICTI
hXEpsfloNuUndqRnlI8thdUkGfgwv8fgTO75QY8sf0P6iIyAypS+bmZ9QcWa
QkVzcTZDNJVauHYOOX6T2qeGDRvrFZpk8fZoqkPX6QG4pyhfeCoSmu6VEyL3
xQfFgVmU3iegRW7CNExeOWDhixKFGphW9UQbMsXthK0MD6MepKLNOQ4VyvpT
kWcbiJSxfEZo8y7DPP9yUUDcYOZ8SC1UmsPBfQfLiGZVS8vlajwqzW/aaQ/G
CEwfcG6BOp1mGVQnGH9SZEJm4FLcYmfbLufhiQ8OZBZ/Bt3lH5iM/NN3/yAR
DKr/jWGkwwcA00C0DYVTREngvKMSfLIGKGnZgDXG/MX8XqCRnee0ltFNuJyd
AU5QBtpTlOWsG6evS4W+ag6HgE2vBwWFGVEyDHctD8L7wAg1HjAJuSEx+fc8
ztpcmAH7KF3Gkv1MnLm1uEhvY4CkgcbV6pqhSftGLamsMGbt6E9ebsD+vwLN
DK4GC+mzPpzY4gUpHIfnEQ8VKWU7Wz49UH8qPVdp53BItPlkRfuaAsYfMb8q
MJqo2c3B8X+ZJdTsIUF71w9FWkAZPSta74FQrei4zhDKSX7mBYmuDpXY9JYa
OgpM1mIGBl1RRZP87a+wlgVFvInLeYGqvD4YoXrUnUtlXKYusJt3ZtDiK32f
zRdMoBuo1SyfbqVOR2TIREZNj4cYZktvj1GnWiLkto0NAUZaSXKNQewBVdhw
mMq5/XmVcErW9gx1bwfnLY0r1Bf2Vuso9Ab09vat+6q88Dx7Q5VMRsRNTnYY
M/6A9eHueasWlN07eAs0ea6lU/bkLk6vqspvCtwmwCGWW+tYx51Q8G51M8Gb
WTkfo7mPmj17Z6J39BdXYwj35U2jlqoFWr/FeDhl1qNgLD/RJVneCTesLzoQ
6JY6NLrxgA2R8razME8ur+6YHY6S6vvwx1CyOGeH8nTN2gWi7n7d8ijt9ETk
N65PMluvZII4OOPhTw5bYjvW6IvosAo678VCyeU1/g/vjjdJbo/Ff8snlO+T
FUOKQe89CRMtY/ldUyhijMXpe8WpxN76Lysx5czdWBElNpAdehvgrZbrTPfr
utwH6QhWlnZ6fKlFfO7s4sroQk2ZIMXuhlRs8+4vYKz9UPEY0hzp5EQ2XWbT
VKcJkoNHGP+Ph44TkNMhnIbdwOJU6oomLR7x8NsRAZSSSpZOEkIqnS3cyVR8
u0NDcsXIqW5qs9t8nQmBwoli0R7KAG3ONZo1JP7Z/HSpg7MC5W/HPbtJqOdR
aX0kMnt1eWLub9NFDlQCNX5PHqQJsGgZpVEKSIqNsj9Br2Bn5hOrxXaIYbRc
VYH9xJnyYDZklSM+QFHRRy4a1wU7NX7Ts6e+g9kEftQWhUU94eeLjgWN+ed5
yaxVFX5G7i+drIqZBXhQi0LVVHpO772UOlhud58PgHNrEWTLspymLupypWpW
BjPGVk5azZvvrrcK+R8R2TB7FEiiI9eYlnu0Ik48UzsNrT5zYL0mQ1jtFBz3
mbkWgh6lumCbkHmWTsvDSWQRq7Z6hcfY5EKnoYZ/2iLL1Z59sMlv9jB/5l8L
/qc7MDOZQxgL6Iy1IcyTlZEcYnNYExke/jvDR3xLfx3pKtAKPqj5wUzEdASl
eCFfv5Q+Geecsj8Hc42l4G9c8dN8D3xADxjh/OKULgC+W18fe91LG8QCZBiA
//pPEYKTyKbAXU4gq66ScFoGLtkgBTVlSMPTDe+Kpbj4hN+QwKxn3EnQXoTd
z0kiyRQHd6daRx2atw9XvaCkcYi9BBOzKva24XQNmF4BOdMUHNIzqby5chxL
ZixKcrzfdHMviX0nj6AkG/19JNUUFS4NANEQZcDUZuoSNZTq4zzJykrp2YBY
Q6KXXZOEVjAKUgbH3QUgoIdyBDrFLBWhIHSpXYhYDRDDl/rPYW0AeSazrrrT
3C6hcE7UG0gZTe7GOYpSyKA1yYU5gpclUzd9cnuuANODkEWq2FKOdsMOEVor
j7U9ITqL9WjEQi5fAKG+rvjoFCJxjFQ2JhDUwMV4SGzbZrzDDsLZZM/s5ACu
DL7KU6ZR/mvYsnBxuRCR1OBfmjpaHLomf2fAIPur/Pi8Ojs+YYUTFv+H0X3I
vmSsAtjjQRkG6dibfxQbOKf2Xpj1D018z+HUKXyXxZFi54rrUW8ApYC7LQz9
UzT93mI5TWtnSveyeMBgKzR7s7QCCP9lPpSKSNgyI52cHSHN5OboI9ukFdo+
V4/XhNGOgkQ40oKmvFp3ZOMZ5k1stL8oadlJmVbSKQ3HK0KAuQpFJRZ/KBAa
z/vYHishUBpH3iu4ARFyVrb57kjL1lbbVvptQBaVLRJuigi/lvMFcNqQD+a5
fw5/oWTi0uwh63w/30c09Q1I/tGXQ41uTjdFF2ia+Y6ye6iPeXSKqPGbhLRg
VShLStZgp4yr0zbPFdR3mRkgEqT+OiJu8EsqWy2nx3tB1ai5qG3O2uqv+W7Q
f4F66OsZIa0PF1EUTfxfaK69arK/wgMe9FlwpKS45dpHGzYfzuY22pdCRtxD
sPM46wC39M3QdAfI8/YB/ufqweywZpPZqvHktssuo42+y/efLyURWpZSleEn
3MnuwWTU7Yrf+f0KNWd445NsiAav1wjyGIIUAegSEciZNrYCKdliac6HRHWj
bm8bgEz7q1O6/jvYF7PwpZeZBFYp5JVL4DVfal8MeSuBXeuvtR1QEbz2HROw
ueoDkv6ci5GYV6A4b4o4u8T+elhJ4CvgercbXEgmBt6XhL5+sxX6zazEoRc3
X9l0y8/Fk49TVGd0r3z4eVhi7zuD4tm+YEObm6JNEQQQw5LPlJBSk0jljYdq
vNHBJP8Auj/TiUSQPiyt85B/fiKG1kLow+5mNzQD9VSUxao+cfdTinp777ds
SybHqBVspZuL88lLWf2dRjH/N8gfvJfUu8JPObZuSc66mWiJTgHEriMDZ2bf
MrNhrF9CYiEMgdR7KNbKkplB16AxdIcfKbDmpcKs8di2DUhXhk7ULvMKnDrU
aiYwKBkSSXg3SYBTGnGMMl0TNmcL/cWPoNbJCi5PLPV3SM9z9GfrXF5rCrv3
JvnqWD81YMfWJQ7j2p+EBNUInVcuBT3jzYzyiFZ6B0VenxzRu1Byg821Ul9W
GOBUb3zbTASdxHE8FtWuYu79u6odX1zi/dJJYsB48W5pzH7H8bTG7lSDHHy8
aRUeilWhshp8XLNKFVKN8ZGWypat3QTBYQ1JEiF9bJ1i0LnmTfhSbd/XpG7f
aQ3KBEQhlFgYR22xc70OgfpIwh59bQOXA/NoAlid+XWcBitASnTqULps2M0L
mFGpDh4Nxv8C2TofXRf/sCW1qSfziZVIWkfotDdwhHzmESeXX8cismteUydk
WUXshMOyiHAbfOxiBf7GyJQ2tAO5xkodOIfCfZa3rhTqrgDCqdCsFrk5MynM
HUEJhAuISRUW9RciMxrkrD0k3qN3m8bTOOQwQJjHwGW5sbRH2Nr9OajweHnx
gRWAUqmjqMg6sP7qbHuRqA1ar5ffQaYI1Tqdscb1NnAUYTa6h1bpDIjTvOVx
X9ROoaGLJt5ob4ZssWhtQhaPAnxC8LP+FSpKuAyP72uFUh8wqPXSnrtoGJ1U
U479ypyDzOzt3PfjqGVR/iU1X9GE0pcy+1El3m8WY+hi1Q5AjKAtq67yLymD
SiBRyyXMi2z+CYtt0HVMJESyHL+nIlER8KPcP69975cKLK8DQzV5OtVXAvI/
/DfM5XKvNtfnN9CBSnO6HaGBVtPN5MgZ8YWIzIB/NYwtXeE/N/kJXCf2qoFH
hW+mCXthhMDqQT0U6FAi6N/gCV1QqD5EYeuqpKDGnwp7CuLrcqVXfhkMbFL3
znGh5xoPc4IM51RVCwJwZ7wQTQQH+QGte2z/ROJkmPcDwMjmjkJA5FV4RJD6
boXr/T1BfIFYkkQQsTCmVEDuheVF3PFVib9JC7rZC3AV/AmUe/yuUVZC2p9Q
n7YQ30/aqnM6pGavJgGL+wr6qw7QlGlVkC1YFL+CUr6PFmnc0IcjEuIZ0/Vo
iazJqpWq2P6aCLLKNyH3Yy7ZB3jSoPDWzvH0EvyLJKEMD88DF1svMZCVSlbY
VeysMJru1o7HM76ibb2OGgykRzhJtnE77mmPIpQt0f58P9JWvPDDGlkc5vdA
C/xTA5mntwvjDdykwvVj7a0lbZ4WOA1FfAFpuG9438bRMKng51KpK/dAgdhl
9NSFdQsno6eQUzF2RNy/Cdz7AOIWHQXhaXMmVXLqFFT632OwVQX1adFksiP7
Q0TVRDTGB6it15qB9tkUkP9kXbnwE4LYZCg/DVSYO2SzWahchhZ91e0MIFIo
/oWUM4D9XHTdgJQKsUuPPCoogzrxZ5L+n7ReC6EpwPNuwLpwlnNqp3k3NIk2
BKRS84RcGSAIt2H+aI2pRHue3pO6NOsJhPJNW8/XtF8RoonNJAznYaY7U3fl
XqiSY5nCer0bZUIhT8xT/tN0c3c8GsnnAzZk2ja1ukb4UOUvd32OPEQHI0W+
dwqGgE4dLfphJp17qJsdQnoF7wDOVlsY5WdhVsZuv2x4S3OwHzB1UUiySHlO
B8w4WQAGLIiivrifA8aroMo9p6WfcG7O0VD3JSNdD18bOirT6Ku16f82W6V6
FaVVhXOTdtzetkBwZPUmKBN6LLWqxpyQPUQwGdMdUyE8oq/FkN5blFWUF3Cy
S6959u8JXguz+T7VoWtV99GRhMym2SQ4gP5VV6J76J6Or+Jqs3eZSV7xMReA
AnS6me8lf2K6l10nx2iRyYko9JhoxpoJGqxz3suEYaXv7CCds+pCusytqHhP
aJKG8nAWyqu1INrbkqK+INGnozv3aApMauzkOCkDwyK3QE7sBQvA20n/m4yq
wCJyGMNuyFPSOKf7IX3iFdeNcOZHtiABqTJex+WyoDR/NDWSBJyC7ZrGHvZG
2p7aUJktw5DtplAjIONqnwsMAKfRKC5Mq1PpOrKTpmFQbB+IV5URwR7FQkNW
n+rDoUWNJcYXt70Ta2ZSbn0WnlZ3jl6MA0vajX5j94Me07a1GZ9iUmlmOBMd
uKbKj9llhxS6ntjN/Oy+IpxN1lhWRd9p60Bnl1GfLpbFL0PHxFmUxphQ9Y4R
fDhI3DZTIX+g4uwwIGjOedhDd0fZc2BsipUl7agkcRGyTTBMdnsHtezWEaVz
S44YkSspA2wTcLEEns5GPmVVD7UJ+wxPifDCDDxXC9qny21AlaYIOjLcNiRS
Yl1NwayEGYhHp29Gb/XMiMTPfpAtgWkZ+Ysnd/poBM2ssdP+Dm27zrmHuSzt
6TJrCDv/i/pI8ewBjwUhmUjZjUeZrw1PAaawtXglDxg+OVT+AAJaEdDBEOFw
lG1BX3JvUAJm13SwKU/P/c8RgR+wM6Ca8Yp1lTml96nLY8LiGb6RP2jwU8pD
mPYreYzUTZvOFC0JNj4g9vU0zU+UXX8YB5Hz121gkR/i5dLez5KDolw0Wgcw
na+rOUvaUEroqtXQ1UrajKGybgfm535np835ffDkyJOKdd3L7nza26grrg5g
16hV7tk3QbHyQBXtBOr9dGKkFfzASBOtXSvUyPufuVZufhew8bgNg9uohsD5
BGtkh2cMhJPU5oXpqYPFSW2xNg8+R6O1K597y08kvpLvNA4Gc+waPg+AAe08
r1gle5lEHAhZKtxGx2PF8/uoIHXcCRlhkq5B4wi5451hE0eETi0GUiZ5zB93
Iqx4Guu3IBWlVaP9wGG35LMKl6UsqJEFiib+m8DsYoUFZt3lxtae2jmwzSE+
vMIuofHnncYHJTFSTkUABqRQed0wZetxJry1WHlrRKwbGBffpbWk5LokeqaZ
hpA7o1zKA+I+mgB92jeJMCAMwYLh8D/fMTzc6r0YaOiqH9sUlvwu9VIy3auo
i0KKUhcC75oJNbiiCIXXcftEj2G5mvNuEFMHRG6uQ2E0nvz5v96JAOeJXv/f
rWdlNMyFxIxTkUE3YR0/GEKpHokb3jh+ZANx+x8nJW2tULR0Ni5MsEjlGokk
zJfHqz7sa9UOE64LTxlk42smtUEbHf/deXM2apocKbjkQ3Q92pza/YSJ86kK
rynD3YewOkNtqs+jgwkEOfQ7bqIMALaGTOCeZBFeiecEKRbjCuhc/yXqZtgQ
wjm63TDKxavREPQe2vjnKlUr4qwMrIISKdvrxY0q2tCmAPsrxH+k0znEEbdJ
pUz9aZnmcHNJRgfCgOMVVSfn+S8ZVvzHBQnqPqUqY2zNrxBivOhaMRZadnGm
KyDFRo9iXeHLu6D/AOUKq2cVeAc6615bJlGeyzhn+HyNItE5bmwQJAM8hdpm
PFvavdT0yQeL8PRlFBXbymoGlXkGReXtR5Ym/MlQh7c8sCI/pZmdQjWxVLfn
7nj1vyUcZS6iqIalNtQiRvjtGkkrn4PAz/llw6kLVbYpHhRSFU06sLqCj7Vd
VT2yCET/qXcxEe5q6OAG6B4/ilcrcbaeZLgnZ8If2GGViGLo6MNDE5xijxQJ
HJF0waoxn7KQ3VgLhGzc5fznM6VyqxnohDfboZFC+M9f0TbjRpXo/rYkHhT2
flenr2u7XDA3h5Q43AtWw7MJObO0AGMEl/gfSTP7QJO4klSReXnbvrhWDl80
WR1rCnqwUhreKKFxZrg9N9Os4t45swNExW9Wq/aaLS5+FKRruyBwqm6W6KI4
BSWRBe2FzWFpa1ooyMxKVi+vTR1tnYGfPWtXUu+rG7o4Qzd189uVKATDLt1b
vpxyqCIzlVQiI1tjmu38H5rFs9szmYn9TmLUEs08D0D4QnLOC1fkywzFkL4P
VmvwtOy39stH7b9NQY9liyq6RDdKmNwC6cH7nFPjEmyzSqsPlB8tcGcQ3CtW
ozxDWkdHHLGLrrG/9v85Va0TkP6rkfxyBhfUarcptalOp0nch3aweO7YowA5
1q+tg3Dt1Ds7FgXWgEt2ZeufagKlWt3gX/NYJVhLGKXxQTJSVz50P6uZhFsI
0TH3035Sw3PPyzSWM1yS3rzp6N1AwMI7Lw67z7Xb8tRMyCxOPFVzGMjXVo5h
1p3fJiJi7kFTumHIp+LbiSx/5HPMuvjQjE0l4yIFeBfAySH9V6OvFfWuVBTT
55beYZwSGhJwJeOWmv9YVAH7QM7SlBM0QeO0AvGTV+sKCgJrsElB/sq5ymfG
3ZFzvLUA1rrVVf/lcQNA/oRXPCLzrmlsK4Cds1iDK62hLq8UfAlbmGjvOUMm
5SRcKicn7czwR6U6Tqyx3HFJO1BzDQdyJXPAATGTgQqSjRnOH3NRhBdm+kEG
t/0F98JUL/kiS6HDC73+1FqVkzC40RJh9uu5B0Hu+189X3l4kFlr95Fs6oUx
CQ7iYd9hWnWMhp8FBsy3N7Itksf3Iq+7E+Vu/a4CikhU0cwC2e3uaZiQFtoX
GJ3W44kbTtQEGkep21Ml9c/DlJ6fTP0E68nX0QAZwTzSl85pAP5Uqc8Tx3gU
qpVPaFQ8XRoWGAi67vCVpa4JawRiCfBnlVI1eEYYO89Y5V2lTt45h6YEwh5Q
ASobYu0UR0KPq8wYzCHwwj8dNDPpCNHE9WU7cPokeZq4g+tsSCU95aAsvaTM
OnkyHtE311iHjXgWABlp3mV1+oe22Wx3eMBZA1lsd+Iww06IAFm5JuU6Cqvp
Kb6NgVBJIbRdwl/FxR2IM0mM1JjsxZZnAa+5DshtJM9lMYa8SCU+/fi7Fluq
u4UmADPHUPBRfoQOh3j2WADwGvX7niWZqkawlIqQmBRuZ1FT9MXCsta7EF5c
RiftYrF20fAMGIWURPJOJ27T4FsJQh0Uv5YJIqhbDFIEaaJTDWbgffMGRNkI
+oL33E+HFgCla2iaFrtrNN7whwgvVhQqPHMnxhUvQ14VOFfv4gvyzAeJOhpF
Sh3hYltj6HNMW3d5xVu+1RUysw1E7wqUb1EqKrzFtvqqPw2Ufvf4TcLbYkD9
0IkrD4iKPb45lySAextF1GZS/4A9qC0N+YCd/dBBfyxnoTqRl5rxnPKZB0VJ
3eOgteqCCa93m97EY6JG4RrmsYvrPjSuQsKrDLz48BzgvpPGucWUQ65xAF5u
1Tdd1Mg7N7qlLq4GY7gUSJ3eisWWMqq1T0bwTvgc0mPsU0U1vgjwr8ss8DFG
BvQyLbMwlk+5urZ6WlflxqK14aTASQrhApZXXWZOyk9+/a4LkSPReCFyYQZh
FNAKrjIzVGWdBM7UH9QDbam+G3jlz70RfpSvX0kuxB/LlF5EpV8NnA/xMdvT
YY6vNipqXRi/UzcEiH2AZZ/26JZ54dINvMxSnusSWS331DjhILli/3PJ+htj
PYCXxxMP8kxkCrF1fr2/2tQu0pnbleECZJjVh+hQcqEMxSawejYAPeD2jcm4
9fty26ZIF5ymWgyTX6NuqrYj1ebEAiPC+e4bNVMO60Q9GBMYg8oHM32yZ3fF
1Q2LFA2ineAafDcKO/tj+Wk1LWcQ9tn6wnoK2oo9fF+r2GfFSIOq+U8nbqmv
0YFAiux90nWhMolJHhOFTbyO0hvjHXXADqGFOSOaUAl03B/WEgJkoaKcYz4F
Da8MpuhcOcmmipIPnbLBjTIqPIN93g7OFno/PA4iekqZZgbmm7bkr5Sd3nAz
rJOsSVPYsqwbDPiGZYJi1Nq+pWCg6lTjUFN/X1l6URAB57DO9Rg6Eh46+YUL
R6t6IrJ4+ygqdnfQHB5InHu15fvlDXLxqp+SaKZsfoo8cjcOKIhlztXCNuLV
lF5IO3UAT5aP2itFFDJwhYRs3FL0hSzVXRDKSb9pFPrPmXuF+hxssqBGpUzs
LAtZ2hmkR6tehTvaDzsjAceliOmlaE38DBfgvL7+RuyhpRUTNZS6oyONw0Tj
IQDRKQUCL3iueUSeZnx+6hHZvIzgV+a055pKztlvJV396ob3vSQIxN38hrK9
bcy2GvZ9/MYCqtVpnmNzMh77jBfQQMf9lJ5+K27pM2V0m6UOXb4417j6dK27
jkhnpAnpiZMsquDrVotiHjvNjtG1eywelMsVCybnHoPvHMuL1de3v6OdR0Nh
NvE+pumD1qWD6zKg3WW3sSGC6WAtW/jOvZxTLFnOILeeEQogQ1FZHFJ8ohQ5
DXL6PBK/xsdY8DbXYE8z+OhpeDEYM5PYMy5TyjOp072vYGoVkAldWnWSIPI/
Pc1rwr8xFwmzll6mFmQvQy70XWcPWF61nVZtolBbiYvGvg5CypROHXs6/2Xr
TY7txMApMOFqxJjWbMI5JGTyZgmQRNyPh4+1iVhBsMWseFMOh3TSkaJShIO5
hRCYpQVEwv1GQTkGwQ4lQKKSYPPHDkBCiLqLILTXDmSqV0rMFRSMX2GUXIEP
4apC2Yh5pLPYo9/uFZXQg8klKAXR8+r8z61HZt1srsqgl2YhOpoM0LUr1TaB
dYm0qCKjWIOCZp9DjPkN360f2qVVUnDX2W96X0L7cnQHNO5fqVgMGamq5Jq7
SY61Az1E7MhIaJv1n/Rmfw3c/ufKa/tDYc4JCS+DvG8gW13wNEw1YhPWgpmy
ShXuKKnPO2qv6/EcrMdiPilkGoRAk/ZOLuQBEMhQnCpUjX8u2Jc5I4edQCCy
suY85GQUeI1Yi0ldUqO5gRJVJkCTxACluulcHKUrmii3D7GUgjKz5uVlM+Pr
CQSM/lH7fyGlb+dqfL+Mj1w1tA+g64wNz0y7DW46/qXjIBUsl8fFvXO3W0hJ
dGJlJFFjaVbs6uZ40tuxHTlyUC+vDtcWtxC0mqCXoSnTsB6F56x1+RMKvwJg
IaiOfof46IgVpu1f/SO29zjGk1aCYIm7paJsTvI/PqCmV/83pw4U35uK0blK
5/AkyjWypOO8akTix/6VQplQ6y+GHhBwgieSyMwd6WKzUGeyVIkICklGoJrJ
8avYH1oKxbfoIA0xt+oyO1PF5NrzYT2CCwE13WiP34GYbx0zit7tjKlrLjH4
73sIOBABG85B8f3iKc1oSbjaBUMWajBX82wpZMK0cu8vTpeie975JEVIX8GI
nSBCHWuXslRgq1yrpxx5BFse3nySF8a7tG4en5ahIE08eLsGFEF90uKTI8QF
vE+NoSF+06k+WxivIFVIkt953TqUxTp8wf+vJDtatxaQraiT954tXsq5xKZt
mIF74Ga3wirnJ1ViRvG8x578Kb3Xv2O1sQv8FNdGdZL/jptNu8UV9VAp1epB
YeJUD8OCD1JFAdbsG6kwu4OUhaMI/CcSImJyMsZKOVsytQ0vq0QD88Jbai8g
fjVo2Z1/1/V2IB5LR4siRRw+ATavMUrSwl0vZi+yMtOMtOT7J5Z7tQe41Lac
0DelxP6Nm/FkCaQZzaXQLmT2+Ot6nb5m+J1LEW55vtKnhZ3qSb716idgI/zY
EqmTjdFmy1UkzqJG32KhOXfZtHstRdQMCUh3xOE43xfLFv4aitgv67we3Lwl
ro8CaWKhGMSw1PsupMtb5XLNIMh858RQ79A25xpFBCO6kZLrV7iKB4hRIiKo
zFBKIdcy3Pm2dLMGbBFbQ10Csx651S7P1kshHQ/hsdQjzufr0ZCoBsu8ot8N
bhZ5LZkt0kTNl+2A0z0s5UrBqN/KHJEPcsUpMfJ2ua7fOQ7ymt7UEpjlcRDD
X1Qv4GkFLfhSw+BKhFeBLr/Brh5AObHn1L3F8MtHI93lbJgUw9ncRz+BVH6v
cWp9yFVg66pxz28J0FzSC2j120xWTHSdVNesAPPjEzWP7V5YjLwVNokz/Tfo
1pCkjGkAVPyb62/pivHWeHVUowWy6cUrunPkvkQAzX9hnjFbL5mb79FOX+Vm
7dXpgGpzlyjAq2fAFs5hlKChaNKgSHftRsys5AXXayCbzi7gevHuQfeuItLs
/F1G4zCxAdzjE00Db8m4IxuX3M23b5gx3d8XkfbaS7lpRj1RM4oyKSjWzCHg
Z6+EO68n9eOS9AQ5O6C0BzTpy4ohrr3cxFlLOzZfPFPL+U3tqB8VSbP3rgs+
QiyDxwsdo3s/lXheVt9KF/mRTmbmA7htkuh2WYhv3ZM6TKGSxyl8NsoWVkCP
JW9q15ZAA0kjF8DOdYvoouJlgGZ7zp5/1Dj9C8P55x6ibu4uszcuqUt02yIw
rxPyQ3tCLfa8nBvXH7aWifyAF+1GInN74vXsMDL4dK0YOTeLdKrL1ZkRSkiP
VBOy6WWUEGgzPOVddTcYbdnMg9aOEdTRzTDRXrfQcYDk65G/nHVesh1+76++
kWQOwTnpnLiccyyWV0/rA20nP8Y5YiRuAotjBi1Vke1nCueYVyVLYu/k3OSx
LTWoP/w8XdS58XFGBFtpQHO2JVB3MEuWDpRkWXSNBxx/na9D/DYCLGoCFRp9
SZQNSeq8ePp+DKb59GoswcVYcry80sfRdYQAGj6DH86C8Gq4moPAdma6uvT1
lDvLcrLXzspT9Sh3diBcCEZCRbQ7CT0fic9aQqi+D+kkIPZnbAsLMbp0vke7
6RVnGvjWWUPiZQuk21FbUfY2jfVaaxoqWema9Um6Yk9mqK+Wwk9n03ZeCDz0
zu8akjVVYVOGs1p41TB3g0rOOWMXmw7AGzeK7lX6sI8g/4uUZPCV9+81Ghga
8Rf2ZKGeh+2udMuHBuSOT8RZeQx9ptEdTyrvobHIw4FJbg077wPu9lyJgkZ8
wHN5OaTaGKAJXT4AIGVyFH8Ph5aK5YNlx6aYqVRZFwMq1F0d6MwxZu2QaMvh
dgNNz2F7RRSjE0PeaEMsHLmXct04Na/4E8XvEBIckODOW16O0i+dJjIZeV4y
9yvf0GhtlizP+ZAKnKt/QoH8+Z1I/bEAIrk0wpfeiul87jCDEQ/eYGUnZORI
uDvrZ4EWMiSKXBz0FfYiK6+qa5gT0Zb4tS2dWwkOcVjc7MpVLcVLM4SnlXNn
0gspPnDCWxXWi8sAQFDQZ/L6C24IfR1XuV0RoX3mphnJJlHrtgRCDvf52e9y
OOoRD0RRO+QVcYEiiDWCFmA3+vD5IPqpVAWpkBtyYwxKA8X8ziTtUDBnI22E
zSoVtbK/6KYSOS/x1Xuhh73eLs96AxgCt5yfzJY4C92K3GwkQFp/C/jLixHg
KH6A6Jl7cw0kZt9lj46G1T9mhA9v8OXzunqDLkjWu097pM5mFHpyXisLonsz
i8e3xIxsAvY7RUqGl365/aBj1ADkvoY1xVuwtylzcQ6mcj+3FaWyOZzjZfHa
6xPUBq/0QFR3VOSOoUXiZlAmvGdDRTXAuGoqpOuQOyevAAIU/Q/uT7GJxxyp
4kKw8WlBOu/9hD4jo8wWbFuPWDypv0P31WIMezbsEXha14o55y75yfLI6g/I
n/D75+/3WUr1i0l5Zm2Z0Rpjc+v6soPMt/CMKHXs14mIUVb43bwMybARhOY1
su4ZRwuQA3+8zDpme84MIasdGLO1nfIVHhExR9i1sEsaD/CrWf0YLv3cjONh
twsrKL4x3s2UVQZ1P35fjr8mALMFJplC4nUjjlEan93FQRWHlgAtCXKjohyA
KsnlUocJbJh3hhtl+HEPDVUdCuyPSFXK8RvP3Qi/w2k5GQXYZIudtzUQFu2B
q54/lyfcm4reuqp35bfvnjAli0Qkhsx3nddYFr9yOVpHmETGqf8l+vx+kVuw
KCqw2SkKICai4TTp3k3mXF0YIwNxBJ59iNH4YNXJJ79SCW1m5D9ihBJZpMh+
OM1MgO9BOU2P9hC7TewQuDJ8rtQiPPg/8qqd14O45HAcxs6BhHBBQPcr51hN
zfViBny7lUxjO5V14t7swrWQ8wnl8CGYRcrx4xGpNvQFCfqpQRQzaP65y9T8
0yn9QHJ7dswQhgkWSFfPK3RdJ59e8VPUiJKcYRxhVzUWc7URT108u1lZ+rgO
zgb1cPL8XACbXqfNWncUD7ZIxqc7Wzt8sRB87jfihJHHQm1s6dLhnTD+qt+Y
I6iC+F/gydnPDcU4sxQw3tlXBu+OF0FPIhCLHCc5QyXxo42wlHT8hg67Yjy1
8tqfmpuonZW4ZnoYiZNxh8bEKI7Irb4YNG2xBZJHQcIEeDhbpQ4wKU0SytVQ
DDmizGenqKmTQgTvhC3BZEAAOgyaQys0fj8Qp0k0OC0F/xp5zIZuE434XS04
FpXilZIddmsLT9puaMwGpWn72ppaYFXKzPazpDzP9w9ZnSX3GtDZaEVtdR52
yXbLUSdyNz8qe4C80MVNTFl0QBV/6qlc1SnrtIFfVZVBRseZDw5zqS21XYcH
8ars+PVJohUEyp4MRiOz1hBNNs6F+DK5rSNnPsLHo2/JU4UDqoR9Z7kpzrTN
C5jAnw+XNVtP0opf7j2JNSYik0a1HKcxpyLeUDhouchMfvNOVGrnO2b7qDGB
1QwJGySnI3uI7KnOPJPvErJQthrSMHjfbomxJ+I/Gj4jCPCIWMg/I1xywvm2
aFApy53CVpN4KtIwxRw/1ZL4VYp/YOQEwpBVnoiaauBxsWwvW9KVNrJ3/rQM
WVhpRAIF+spygVIPjefcVMqqzz6DO/ADAKkjm052vhZ8/KW6fnXhJD6WAiT3
nyM8PJ1Ul62ltQtOnm7ONIVQL2OGaNPnP9RRHTJhtGrreKPoSGSv8SHmWTQA
PjdQm8z64IwQKmGaV4VHFr1SLEDNL8UVIkxBYoq5KXU/Dll1+znf9pXm5JVU
zud0myy4qi501OtcWM79pYKoQpMqv91guyu+bFlj0bRiUk+J1hiksKRD95x3
qpw0WoAs6DlbzTudG04f+5M5ALHVXCzmq5ST5RGK0RpOerXXrxopk5182zjv
rb3c2l0XwlMVrHX4TGwSVvzba5tbYLs3Xr0QjN4ly2HPbZQWIz69o9fVc33v
jm5jNBEfvD+Fltcw2aLkO6DQ9aiL1QUA5JMqWfyvFh6YKcv1YEpnXGmt9kt8
Yl8Qp9pbw1f5yhBz+8vYFRep82Fyh1LO0Fx6B8tP7cfcjkuIf0yHxXpJGZKE
7txE6r84f8JdcuOvKaSQxFjMkMkZ9pZPoeFfi3o8na2FPQGxuAjnCuYDWlyM
I2TXFPDCNR4T5K3kDXM/AE6QfwDlKxelGG8wb+YymuyCwnX5mQ4+5a8rAGtO
k0L43aJR4Sg6hjAQEImfR4QbevwtHBq6yCr0bNA32Hw7nWx3plXSfMHWQu9w
YEyBQSSiliNNbaS9651HPSoVLMqYq+Iow26EwRxws+WSJ/iix1nR79M0cA5E
G1SxMJ8DcTcmFqtxkUpIysqIjfnZW1QbD/qPqqRWz/yfmF8QSgCUqatUt3nO
2oVQzCahU+kLiQeEN+6/uxCOeWqq9fkcouiuiWPn7kwNCqYLpu6eTI1cbOhu
KCKPuwQ5qXalnOS6hFz7AWvfkRLO/h8KOPhwQUpoRw19dbup1QNkCko9KEa7
/wqHa966Qf8crxR6W+9GfCzaF4QVlZygMbvTGT2LaWPjaFlcqL471TF/6UmA
/2nzQn1XfWU80uSbH3OThqmgmXvogSis7W0htiuaLA+lHdtmCPkR3srRNS5A
3dj0D17HoCpBZVWscPKJT2L4g23sESdM7MC4WMaiDISY6H7bIR8+/fdIzn67
MhcJoRIqJdA0aETU7pJ2nZYdYytVKPHxHa0gK+0EhUgH/P1JGN1z5fej3Xop
caT4jl+XU0QCM9oxywTTZWpMNYOP18AicxR3yUoMr0iTSprC3dv6Jty6TmfF
gen/qef34uICli9BHt7YA25gEnZWkGHFAdy3MUoiMzHqTDtvsUqBbOXeVAAo
QmX3Af3Icqu7ivw6+O0k/ryWhhWSeKEhgebOT5nu9gLeeeKvMWSa1CSpm9Ur
v1OdgBFAiahobjzzIGK79MVXOCUvEMva6iFHn0lrEQgwGLXnyN4R7cajBpPZ
IhNUs/lef4Nm2+UQRd2JirvMF2gVn+n9Vnu4IHUaAoCXyp7iO7CwdJCeAQ3J
zZVizr896E3WAYgXGMj0Vvy6TeJmKXPfTl0D3qfStkmgtSr6mIkxt+Mo6JHu
0EuOIR9MhAgEQz5cBqRUX6/SrrFgG0IsYEZMwsWVNSwJsFNsqtrfGTgDdoPf
0mA5Q2d4ptb2Tr1goitK4D3gH+VKCsMPQhJApV1NW01chiyoN8JGiHyGQs/c
ZxLiNHlMLhHW6qDHBselTOHAY1kOmFWwYdOlveWITlvp5QL5NqKjTV0GdLW3
eXZlN7KQ0Z+Znn0eVjz3tPcIeo9FRVPxcG4XpfZjPQMH2pFkfgHiQuDdoWzM
dnFiYZl/Lv7r0ZgTbHrplQVwHWKhb40JU76FxBDQJ0xNvpfoQDeHI2akLtRQ
EicqXnbiiiZNizDOvNrAd5G2LtaeIN3nivOxkfz2W0NQF9eN2elqm4DvggLK
X0R4VLrnqwRvJ3w7n3RnRLCOZmavCYSAZReDefZYsL2FoVH+hXkTj8Clcoad
ShLQY0GeKIC1+EG1RUhHxNpw1jEACtv+MaicZC7f03wVlbo5nNBjAF9x3rzH
9T4B9z3WB2pOcATIcHIK8fFK5vWzD9fPeqhZJcMJAnbonBIhblm1ayJNvWFr
JrDB/UcLjDd9UtwzzgDRtZOl8AAzjpuR1y2hxL1sB3sZYjL1b+YVyDNPCip8
gcTBhOn98HdmICEWNjZqgDFQKLSSagnVcnuFfEdNIbra4XkRzT2sod7WbDQn
zagYi3D/QPXKDhBwhzFXvnFWpNEUH6IJN+iidOSJFp0p/aoQxM2HCTqve2Y3
GOwL33dVczQHvmOi67fsrbcGdBkJz6LjO4O0ntAqVd4Wwbq+pM60YdD8zM9P
dGr0dv7rR+FsU0hqXgQKL0+FBWsEBpTyA0aLs1CIPpPJHW5a3g4m8bPQrW6M
8sjdb4eNi+q19bJHKWGXc1DPFuLzdOLULeInaxSWI2aIPpPdSwwXBCO5moh2
GxzAtZQeNu0YfBYZbqQUXUKvsirH/5vGsqYpvamHiJF9ELQFCbrDOAT/5TLf
qQuqOEvjD7bx08kBv0ARUsM5Ug7Uc7Ban/VP9OGjNEFvZK2IYUwJHcG8iepE
eT7mP4rXLtiw9mq4F4VXogpM0l6O/o9huY3vvZ7qTkYDzs7QQ0pKCXDKIv2D
U6Jqm/O9wvnX7/tsL18IrrNGaatK1GZJzVgA0/1qAnMiBnYvfy7LGs8L/enQ
o1eFFWYYVSWWBwS5gbVJR44828uyktY5KjAL8PEnB5uTz3wcHwlNeZXx+BnX
756O4ydBdzaX5JCdhAVD//SJ//6kn0zNkYpbeR/tbrqOa7B9Gw4mLaafJStV
pVcrfNCMjuoWHjWdzpni1/vVBwowv0drJdfbkovAKD0g/Aobq+DFWjX76r2J
LROjFy0aL96587amBojpcbo+Unbov0nmwVTtTWlfMKqIW3zwhWxojjaA+utm
gZHYo847UmbJHQ9QP6FYizFP/zWcwNEwZcYujN3u1E/OXIILzNZbd6avSuPE
fJUSyr3vqtQrouyAIDnLVzucqQwFsTHrOEOPh/mjN1mLwtz9Jy1/J6pA1dHk
r54NGUvmYGk/5bLfqI+Cgh2lv7K/4jcPZBGPFkK8e7LS5Gs1sJ9ioOKfWhFM
7KrkL3yxdbENfLj/Uuw30T4i2om3priqYv6BT8NLFWeumzreusZjzRTl/sbP
M8Ra3cqLSwrUO317Y4WuRJHhACmgiyiC0lt6JfQJkmFn7dEZyznPirivGXkt
GM/Jff+5v9KNEC6dSVblKHMDhG/6S6jVSrvULuss1po5QEFyfmaB3B4HL9Y8
ihs4tBMfpwC+zp3EyR40NDhfGJyffD9h+p+UNMNd7gKjBkHUnK4XwuRnAVfj
zJWOP6Ociki1nU482cKnhu2vXqoSIEGVfpun4CDCo9MWZHi/ETFjwohgjzFR
0SgPO5DNHiHoIEgMkW50SleAcbSATqp6DgrKTi+p2jKaPz1kV/ueMPGR9eA+
51DH3p6OFPk6Yvn1u+RiyABmx2JUijtLv9ZFQIqJZvjodCkLZhwf9HGSUYrM
B7Z6eULdI7slCzka+2nj9KD9YPdYDJaxQIkTxZKD9OIaKFExaAa5X6wS0Ktw
naZLETvi/SrdeUhKUz13vIO0/UFgNwGyk5bbOqYwtq+OqolhHEy7QCa6BnBI
k8Bl4xvBDp7EThO3m8sAlWulvMVbp8uHEkulnWkCXgVAZS39sWQuHWMxJYCd
WIkjlSTHXVMg9a/pgLfyVJNJH5t+jISfn5XKnOy8EutvEs0SbXiPKeJ+WX6k
9J0qf5VDALEyhhLKWbdd3UJhssMfgQCLWZ0myTSo9LBM4ssPekCH/P2nhenC
V9IPRSOidlex8pfisT3+T2iQt9qUDAjlIYv1RlvNCvfdUzpnlpY8TI9wU965
ncNGiXeuNClZFjlal7RCzfPoYZ6dra2eR4iR9Xz8HwZxeOtr5hkcZyKLCIXn
ELwuFL7u8Gn9zcBcZzjgP8KJRDj6UP/Ybuk9zur3wEoAbJJRQ/9b+qm2XOsd
5K6yjD+p7KRMGex8w6kuIPiOAKDAFTBBSi5IWtG/eYHCOXOgb3mhiIMgSDlh
RAufche0xeQhrVpapy5ztKiLEvhkNYTtIGvzQuaMctVrqZ2CSYbc4+RzMtrI
Mmk+mGykb/Db+GwMWhmd+j5u7+R4Jq4z3u8PtEpH9qjC+kfEdK6bEqgUXZxv
PrDai+SBh+bzwiZfVoZRT+4oDFxMoJSPrhA/S4+pnLcONfICotwSiAm2xnSm
Fskh+P0BlKsmTQBBiyVu8jwe9ee3CLe70yTv0smwJvsOFisw4Lm3N8f/Nqs0
egkfbATHs4U55l22iU2CaPCkgjE4/ktyIlVku0X60WhZemK0LHWcbn/baQeK
njIxatLT6De6js0BIvy4SL+q1l7iPWEzU3+nA801EI3bNaMAPBs0eFmcGCK7
Sqan5foiW8rPssL+m8TWght1t7ye9g2UNuJS4con2ek0G0gJT659JnfdPxUz
9PY9K9eMYzcnbfVwS/WDpPyLZAhuIcF0V/unPzwOVw208+wRJ0Ubfdsbj7O7
vHPlGZqfut/45og5vVupGVDR+h0ya7CL65kyi8GF+Eh4aTUx//P3qruu44rZ
CwnZ/7mtyv0yv1oaGTGccSkay2ChAF6JkXCsIHvbr7WiP2UlN32Lp7ztOpij
EXlIalylx8q8K5QmfIBeqzOsl9/yZLX0FsEd1oJucw4cYXLCPQ8+v/cSklEp
IF1m2RFqgSMfsb9VlpMZ6Qx24GLaH+9v41ef694UQI5qhXuJhqccVKUpl0Cz
8kfCdvqn94bdGzFVO82xwtqMZpeCpRyl4DJTWpoCJiv9T61F/5D7ZcLlkFSt
Iiizyl0Ed+iNwZiX7OlJkr0LlugRR4FJNO/KdqwdzKmaAorWVV/UPpGyU6UH
7xFsJd9wEylUBeNhytKMK2WiZsZK5etgf4S7mUo4OCYVHHOkIK1PIVZFp+vg
2I8G+LeQndoPzhX6I+7pgJwua8wTTUxKoZcSs1UId2kF1uFixsiyFKVCez7B
2fWcwpXaRORO8VOrhpV0WB4hojCYW9FNZ7dbgfzqpFdrM8YUOdsHvg79ra8r
x5v23KlaAsaMynsiII2AwOj8shl3i5naGX/D2FaAYym4a9TIKlbk29ZCjvoi
YUjvDRFODdv1CsVW/NwQJp31agbAie96ZC8b4iWZx41186URZLPe2TZ7xYii
ivI9M/eWri5imu1f1LrCdZFk8WVf+/U+1mdNO/deXedPct/AMJUc9lPuqTDn
ftjJJ7GqOIM+By7yzx2Cn0f92CAShf5G4kfwr5qQ3KMm6yHA/sc4xYCh/Xx4
xPXYYf2+GH+yHHWzKss4lucXcZ+VBE+W/6LsXp2ebPVp40UKYVmh2AD7+hfM
TzquxUuiZ2nJ8Cn11ScBRHPUY3P53+818TKz0h2pZ7DEquVq12rCjSFdOsTi
IWPNigogDA4K8Cav1xpKQvHleoS0y9F00imFnwkBiQ9OfXplK0bvolwDxSVq
KmUoJ+5Qu/cm3u9Aqi0LAkEIqfzfI680tbGvu/0JgzWkt5Uz+wA4CvHiwFkk
zsUJjCbu90cqU0W27rL9Rd09KsUYfM638fGVodCWgfJ7YFORL6Pqr6OcVZy/
zyrKlm8x/SAgLv3DBILdLrY1CNK2j4lvksf5d6FzZi3LdtyKCwUUOVoLFhfw
UK4KqN8GlOtyItknyvm5E4GMhbwBszpXzWCRAgqKWmq50n0KYB5YrHfjQlF0
pSokzB73silZld8/FPyBBGOLH5ML8QktyVbcIh9xHxgtCDEP9GGI9uA8x5bg
xeX07xvqsYOYUJaMD21mNiYNZFrO6vTYqtFHFKxYkJ/82CahqZg+LWrkhnaU
crWATj6FOmCHwgx0C6UOa+AzQQc5OB/0wzUTOW/jH8pLuZrugKTxeCtweohX
h9mGyEPMmz12HDyG6fjCr7fZqJXJVUtK8QNUN8NUBCuTdSjukVMvGeQiusso
/n1BjL+1I5JZwJDkJTpI0SojZ/T+pPpOqrSSrKPdsfLyv/TzNxL1eN+dGQv3
nGiqkaRWVkcG/K85PWoHn9WOpTWudW7rD2KMjtBM7hhios2tnv04nlvV90e8
UjC+QkL/8F5y3woL+gJQlHY8ypSsy+xC8uY2V4fB87utDZV6G7YDgIOtV5y8
jAQdowSUruBkhniMMzqsQ5jV/eY/UNbY/AbcyaiTT8dr01tqfuuq4hu/lSq1
/T6HoMS4ijR0eiV2DEkZuL6xxnZJzIBMCWrfKp9SeIm4Ab2IM/jvZ7ywoaY4
6FsVC/OckEtoipSZP53I23Xod19Qd1QTCepFvewsT8R4/s1cU4hJI4uAvrrR
/EpGcTChpwLmVxdUwD3CVL+PWbcpEdmIIFZ1RsgxjJ8xL67FhvEr0FLltRNx
fNN7QIhMws42/mcx5WkzBxh1XsdOYgG5NaNY/T525W3hHMhwGGZNtgJfiESy
KS6IbV8fyiQ8SFvzWxwh6tI2Q3bDWvF7dsGblaLqhKLPcZtcAo691WFOvJrB
yO0SV68dELGRLKU45yzbBc8nBrgdiqd2gWH5T4oQZAu4eT4AS69bk6M1dvgG
suosdGT3Q00y9BBH14e+4XWvg0RlrmnCQaglLAGjG3yyULeoQh1wUrHF71NO
qTWzECMmktgoILXKeY4Q2dpjQ9+/KzOdt9bhWrPtCkFrlZ4C0b8V9/MEPSQS
y9DXijHInytMW9xpak4otFtKbTsa+H9jKto8iEFuEDZL27z4CPJBuUCPMF3D
nplZuYCG3+x3T+B3Ab1UpF265eJ4l/Hz7iZzbfBLhQ+i022p5VdFj7/arVgP
Z2TJSPfEs4g9kpDYj8+q6mgzeUfbsuBwTAaHBdbR2rxHxHIw/q/CRA+PZK4b
1o0WE5KmgHoTkNKplSryzpLdtRsQSZXUdsXAwBdFQY2cApR0Z6GkAvB01k3n
rRKlOxabTS0pCBedxCTFd3XXAiH1CKrBHe85kXvkfG/gmlctiBFBBQpwP9WF
dllmVhUww54RjmJUWCWiaKmBE4ocX7GI53UP14KizmQ8K8ZVQNk3UxTnWPlX
Jn9IWzS3k32hWqzl3ivtkmFcP8HHJVYA8m9VaVV2iZADG5KwdqY0lnRQKTfr
fyhfMaiiSeIKZle+2s5b8oGSxnH2XjU2qEQz1iN77gPePcv+xq84/ytsoQlS
UBHnVk+dX5TYfMMKPlDotaeqjTZGCWqhOQKkrJkV1Yr6XFf47kgbdUNwc41r
RoaHgyZy8BsNVrL4IffaI1ssdxLNQ2Li6tg4AG3RqdZ3yZLR6vWxBWXy52rL
NkuGa8GgHunamEMPprSIx8nJL3ZFjQUJpAI18kewjekoDvqzZRt/ODQbWzo0
6Ruv/67AJembRb2AV3sw0u5j7BhVKXxBnoH1MzWSLdWAmLpjz9y/bLhBHy52
uyJSoeCkfgmkK3o7eFL1/82DfUmO6ME68vuKpxeyoe5cyV1QNbEMhZ2f8wlY
qsxW8u2D8PFEc5ggmpXsrRnkxinACCkrjWCaNiLL78sYKMOWmS/QvvPk+6J0
x1nY4CIwhmFOlu4gDmw/Pc/F9uVl65vlY1xyq8Q9A+/Wd4awBlwv1dsTHW3y
fdytWAB/p1Qcj7WDf62dQLzlgLzv3z/fniSQBubzLdIEUca7eh9HJmO7wb5U
Nb91GVtC4LFdznBMwP0f9WDd3DzEHdFIdQ344e4T7f0idq+bL3S2VFQ33Fxa
uVMtHcXGO0CeGMqotRqBUflAIAKF8G1TzWAyZ8w5hkqgWaY3cjfzrkZc1Hz5
kHQUjPCigS6zJuSYPunLl+hv5KfN0+0qFbTngUxxu+vwDVn1ueMwd2kMtE7Z
+NDR6ZSS1mifypfcpwZlizcJUrl6tNTgWAaKBzbK4yUPcpuj/wHmluNVBRCv
Gl9MELJ6UMTbZ9xLdgQRVNLeDp9K//GPkthj7O3ghWmibXgvYENRFc8kwNFu
H1vf1ODTCP+g+MR4WOxiXV3CCCIWn/QTJ5i+Bio10Otx0CJjYdxYUevFWoAk
QiCV+MhDqtk1vSZ/07CsWzwkZQDelU3sv9/08t0dxc8Pp2sU0NOAB+T83N39
ABLtVJk8R9dmPsrJUZG3an8RIU18f2ntOk6gFZeESQRb7pf6SHg4pAyac5Nx
zZKYXTlAfQzRbTapL8RHazKG+t17zvJ7KDNpheLrl2cD9Z5lsDogVU+NRlQq
lXdwP71ta4YlWIP76UXLxIK5NYAqsHUnaXsd/kr9+GuHgNJKyUsCUFTilSWw
ok4YwZfXfQZXwUmrT370CewHHlCniXofnEie9JI6hSubDrqNN6fbRz9q8ixH
uCjckbPSNDalkQJtQ4r2ic9f49OZcxABsA7+m2lLgMn6RxxTNTnCK15SLeer
M8YlaQKDpvZ4X1iWy+eLQI/yqIHY9GVUyxvmvNg3wZWL0BAzc6rzR5GKoc8A
YQ/fHg657RC9u22b7NCUYrsZC/Q93hi4OIaYglTQOJWEn6RU2UJj2JwgvL2U
8Grd5L3IHqABbaTuLCRErBardI1BLUa3oqt1ObdYTfwJF5LSpoBmJfIf5a1k
1dgv48YWtHKHwjeVp0GAGcUs8QPfoqdX/Rs4zYXAXw4uat7KpzyHyczRv1GO
b2oqdB+qF0gN3Qt+DzGqhL5SiGww3m6zIEobAiL9RqqTQ80SoLUc91PR/9/T
IezZfVCnvPyBG+yqDcHyipIXE/xSJ9uiJtxxqoI/BxpHTeuHZrDvSXFhqtdW
XmbjCW+h7AJZfFvojEf6euV5+3L6QP6XRbWjDcF0ee8u/eU8SgKG7VB7CyHr
VlDbfRinvYsGD1VvPsdftf4TyBH+lmzh4qbLZ0BemZ1Nq+YV/he361DK2gCq
ll6i1KSc6dhJmJ2AGzIKUa4gqOggh1nYP0abYA/Z4c36vprZYrKNoDlCa+XK
GeN+15jxJFykfeNl7+CpUbWIU8O7s/N//AGrsoEybdAbn5TTeNtpqa41t6Ig
LufBoWaKdSia77ixvbdYmEbE2J46k5UavO5HxmlA/yV+FGL1pRM/e5WlVwIn
cpJmy8imGiKIvSBylz4kStRsuGWZ5oqHkGcJ8bgUm+EEuE9nxmPuY4RBGd5G
ykkCo3rpjENYLqtQL29GKn77S6gl11H14jH64AQOQHXQMyQS2HhttObcukzF
XqA9gTiaBPgV5QubMem18bUXBYwKPo5Hb0YKPCoV1YbwlwoMaP+xoR9uaD8D
7aXV7ziL3JFK2Ves8q7prdigdD+R4wXU8Iflwhnl2uoWumZ2Lj6ayYoaMED3
/bQ2YISJv7J8cE4rxKVr5XTmQ0lA98nFwLp0Z1ErvyyqFqWr0bgJsyhDes9V
JpctKv/LM0XCS3rw2Y8FPdO8oKzRhBWtV3l0zw7SThouu38y3urCxz36NLgI
HQWeKhc2l0wMJqYvrilEcbTRFoFMyS2vIckM+lKLau75ZbQHbOyHvRQ6Sz23
gMOYf/1Ww4ndK34BD1oJ77xBefO2Tqv2CxfcoeKr/75D9aN9cTQHs/pLAFA6
XdfBOcoI5kcHv1BwzSJJBGUDVMa6eIdzBXdTPdnLLIuAw3COFPVdz2QW5UkN
9h93tR5Jfw6tIfenLuRovwhdz3ZX1SAU3y30bw3JdTfw7UPV0alxiQOzuXb7
fFyzQ/3KQTWxKR93ByQzUTun8XXmKimmIH0IixnaT7F44QUR2U8f9XEoE88u
B2zaQgQ1B9C2MC51xMHVvOD8cOLosKKc1R0sS9GTPc1Ema0LijptwDMTv3Yy
838AInJ5Bd5qzDnBvB/GwZllNBYnSQnXganQvXhQvXTAWBF1a/mG9pwjBCOO
3S9RUTgyICaEwEqnrZq2b/V4SXFJz2MQFZUUD+ehGokhEeuBfDxWZrAc3PJ6
gaxsCPMGeGaveG7f18rqgVFjuLx+F9a+Uw72lK6dPOUMv98a5G6GTyKI4gzw
DvTNJgm+MyjvNPH4U1jqceFtfM4MdyxUv6lhFjM1Cl4BjnniUpf/ZC/T2SoS
wtqTsY0SDgi7FPSwj8h/+JNiQ+9TvKUD9DQoqfQb/PrI7RpxlbjgCUle/SNR
PY0wGgaj90uVlM4/5gRmohJCxvn5tnbHtJVqySSVq6xNTmVQH6r+7FfRDC/W
NqAfz+9PZDor7/k0jWYRIpGNO0B1zrAtTz745PZSgj0H2ZRMewiLOnPbDJ9s
qGx4ot6BMxBzN3HZnsKMKs4J0eZ5KMyj5GqXHxYK21y3uUADIsh/Abwz0zeP
cS7FgEP4wnGBbMPtm8FvRFg3Cbm4Pru7qYiatNaTqPKfxqYKZpGfxZpP878V
9wgruh8B1GElPH4k3mnJqys9YPYEPHxLd7WUAGm2R0q+L/29f0x4HD1FwBml
JHAVrmMtVDft17V1HvbrfL68mXV/2k0xlLDNYTAL1Ix6X3mukDFgbMEE5fZg
IFFQhlK6WyJ7tAfIP6ZPkp2PY5nymc6JtA9qfGtvKD1P1BPcL0lsc8MayVe1
F+qJ1FBkD8hKD8Ldq++ssaqlQQRqXOZjozwz3JrBHWTefuOiTGEAkcTBf5uo
r6sDNUbQOqoQwUZa0i2DK28iuQvMj3V71A1j7rP0Jgg559RVwEjoFXXJ90RG
XVqSIlZhff3n0q+aH3VP5ot7ZhGPTes0w+vF6h7sUjpzPxiKZXl2YMuMANyC
GD4LJ5UCJtrL2tHZ90iy1PaCjU0EmveI7fFjkbtNwYHgvCH0S7NPZAziibqI
Sqo8QLWE79NC/RIX5rJfAb/bL+EGQVtSuFgo5EqklKEJ+2v92XWJdczAW/GQ
CmQu3O2hpxxCNAyCxv8Mw9PLQrvFfStDe1qOgvIXjOt717u4Bo+rOPp7p8nK
sHscqSjLCEIzIw8PGxqaxmslCB+UaTM9Anp9ByASB+bsymmC3BIceka/yjv7
ZhdWj1GCAup3i4hsEuWhdCz1heUBPGxTnk9KwAjUi/yhpOt+Mjc0olH15/u3
h4jM95fDHeXNR+tdTCHUmLDepQdtjDF6SrAL2a6ZhhN9Ft2jZXV2AGUfXAH2
EVViJ624m+5ZsjrLatoTCSOh+DqjotKwRFJDFw4up2qWmLw7Hh4GW8oKfB5j
bGZoKcUBv53Fj+UaRWhWjeqJE7oNw/yMlyc1bql7UJveOrbiDq/ELTreGXOj
t4sKDRgpKIiTwa9Phj08t2y/SUS/MxBjt32NI3r2t+Pp+N3mQrHKcvD/aL4m
XwxB2Gur8C747lIjrqPTlFeL3KSXkg1aZesxu/FouMQh3iJvBqlG55K8uonk
Kg9mooWVU/0IS1tJfw2V8LLLd5NrmnRjM/483Askd4LoXDwBy1Iy2sN0K2e1
hELyT/ruTVIXorr0PRZ4Mugf+BXetimXjsoi163DLDsvq3FVY67/xWsCuPPf
FL1XzVqTMjb0qg03fWNbJHesK1vOmM6RFs2pwEfru0Sw/lTmsAbIMpwpwXoi
WmeaL4pIz9SaflGeDTmMBX9xaWyzaYDgjLmPNY7XPzlbT2gvFXOEjT9pGH1g
9gDg6Luv/fPpSELKShqVPWtt2cYLB9gDLjY8rOr/j1mOxhsYMKVy+9K1zrEl
+wgX34fbYvgnG7GaCorROCLGAcCZaA7gHb9VioyfKvZ2unoZAWcGpuhwHTDB
WZWzP5OnrXYnKl7CsIfHUKvPBva582+d6H/tAsa3XK/FHxjmlFODuk2HKFRv
F7M8YVqBHsNO54Hg3Eo+oPnBYy9LtXvTZsWjcCe5tysojuO+y01FE75JLVl7
BHMhQfoBU/v2Nt0ls/QkvBRQfPoNNoGAA26i78kbO14WIN9HocWLCYvXDvXI
Cf9UmJl9qfvurx1V2DEGCNptd8w1sr891pRIOhbSWCyRi0/W9yR4M78URbhN
R5DntyTg/pzhFk/VNMAnnUmnDKiGW1XMUF5ue8euVJGiQKdiSZ2KJhmsSGYO
XZ1VVjllN1K+Fm8j2zsFusrMdDUGi6FtgQuTAv6i9uJP+b1/rlzt5Umb4nDn
AGKfU0XU4tRTwxrKWw/mykL3gC2gtuBCJwGxKRueieRLHRBrDoXfz4Qk1XGj
ZLXg7jZVwCF2V1rQr5pHpHKQUqcvmMBzZzeDNXvE40JV7O5o9HkqGBkL5Dh5
oonPFj2qsGzjtHbNe2qx6uSkNVDCZiTJG606JFsSjYJHGw1euSth2f8wRAUt
7vdAmOeFmzwBH/2JpCEhTfkGiUJu/HAm+p4r/VrlGuyLJM1BYThu1vogQvCg
tXP97vX4kIAo6cgkN0xYg0UgWfyDNT88A0HHKgggYiq+uxU1ajxpQITFxe7N
SlimW349ol/tdjlOn2E71rN4zOF4+RfGBtpJ1JWOV1114d7UCG9c7pI0rNsU
kPnXMcvsGEQ7I6jOa90FuiCi9XrQTme9Zvr9tJnSCyQ+ii3ah8hek+G2rXPk
xOjxM9tsC9MazLLVX4X9lm1kH4VaGz+hQ0ibs5ZOC3qmynQmh7rD3BRs/vxr
bSK9xx5VuCIq9cK+KsAtZPvvDpvSK85rVsARqaaTZKKadLe/HPKMd4YyDMw8
5SoJZpoSgJkVV/P3YARZGedVX1guZZ+yijUbf9TB63aBVF3wEjHJbuLh1xKI
Y8OfnPVUEhEqWsNqfm2t5Jh16y5G789cY6hG5Tm2q9jve1Yfo0CtDTE1FC6L
5S5nRBHmMLnW+h/V4b1Piy8F2BmdXR+dlMJm3TlzGszHjox9cGCDfgWFAiOq
JZPBh33m6oHXO5QqxV4Pk38nkwG0FwMQEJxxxHXy2vtmb+HVLdUa1lbiCRTI
qmQqzUQha+P9gac4goE21vsRuccAxzGdOas/PZwhB/S1V0Hgqr8yEJd5jEUQ
rkmuhUGapsKwHDwiBFmyXtvys0/3TER3FJSB0e62Bp9XeU2Fc2obC4sx84vj
yd9BpVvEq2fQSnuPuMCGWSGuxSJCquRYf4PyWBUQf71WyZFcpJWRHjEtaemi
cDxnZTuF75X6ROqSYL9eX3M6R7WdSPIRFWt2OHmsAE906A5FB1/K+unpzE4w
5S+R6KlisLqZW/hRO3TolcYwPQNZdx9pjG2kc+i1MmrCd3NIDeUtavq3b88x
NCk+dZ6Y23doNIKHu4YcZBG9jOdBR1IIeRyhIUuSehxU36N/Hom6xXp7gkXU
5NeKpLiwJic/u1LKYNu1G1dRVJZwObERXQKe29LxcJL13nNCZQSZXeXRZ3Yq
V029NZqtrkLzjt9IUW3nq8sS4RrJu7SE8NHRvt13Jx7TMzMYKz9PAPNTtZNg
vxuKyag29zJEvUrR6Aha9jUQCqUIJl2Zo4GSrTMxvAk1hnBo54EELMnrymfO
IR++O+Aynp2C+IAjuygfjrNJUgF9ge7kmsWx2e/Sy2us2nrn3BCNLcI+jZ90
KypZrPrJNLA1k0iTTv9zvwQKtbC/cRkwuj0TgtkjKNJHF5H9nQGsSlFVpFqJ
gIokk0u+8bIYn9IYCkHyA6VJ25GdI3zZaojW1KQlDBMDbON3CT2QgL0CyHNA
NCT3iDHioTU0zkD20yH1On5RHow8V3r38mSZJaYs2rk5sVuiiLMJjR9GT469
RmqGhacmLPcmw7iBrmNm2mjoLvlZulXkv6MIAQUMzsDkDUatGD8oetLXdpaj
UFrBVWIMLg4DrCn4IOzC8PS1Fsfg6kj2q+fvJlcFQtTKEgRjsy2ks1ACK9q8
FjaZxAyL0h4NM3qG68PaBukEEegNSSAR0QF0aEaJCf9nHW/FTHontn805cnY
VmSfpsCRd90o7XrbMq4XTVg9/vH15OsCrMbwfb7WJNt2Y8XTnsVh2uMQArzj
mpAjbipOilJNoqKSUHb3OIUNsi2riwkrZ/6k6IKChyq5XU2cm/X0ICbXX6YA
F614DCl3T8441fSlG61zimZ30IuV17BxwWkzANeUJ8K504RsQvqNOgctmMIp
cLCNcjGLT1WERXJOKlGiTcoa3LfbBJXgliS04MyBLWZzzieo+UHH6eYqp/CJ
G5hCzWzcgEvmhXxafhx5H9gqQiyrPk/lo1rMWQGNEHMSiF+G2Dn4Ewh8/OM8
7LujfaXZadcKMhdDnD/eTH5tX69+X4De8njifFlm5jbWXe+fzjIfaUSDp9/d
sFj58YKt8tlO2JfhyFR7JnmiArDxNWtUaAXWi1bOqNsg2zsO5pvaYRF/MRu7
jc56arfx9UmGalyLlqwamuvES65TXoN3/w7EO4F13WxpufCnl6WfOtZ7vxAH
/sMSlrGnFsG85WTgSQUev5FKZ8Tmb1EObGl+QRi76xI9QHydFTVrdnHdO+5g
upWggiuts/lRd2Qk5trNvq4kTK7ZhrOXf81R0UGyWo01g6z3Ir2Yc2tOmlRu
TZ0o2KLKfn64l4VgtYH8ugPScTdZ2fAKxpr79HcJV4vaH3lPlfvHMdNH19l9
+0T0YQiGBqCoH09bKE9afIohdII2o+F/20vp1FhxbLLE7NM3Sw/JmMTfhLqb
+EZh7obWXBXHQTfNfWL7jJ4zWhiAt8oiKeMcq3dywfiAN61lD5BJxPZ/+Gn2
CsLGBkipWg/gOAwWhsfrZr3necT3zvUUyDWZqSQGrGU+ecE6TrGWRLVFGCaY
mp1gHewpYGuBlMk0dicjK2qRH0+03gHZxWGa5v0DFVWrFj8vIDm3kMLx5fZs
sFNAJnCWKZ+Wpdgb2rMohl0hYK5j9nCA4FbLwUKxPL47p7a5l+Av+hGPd/dP
oxoI5UeNz3eVN3gJf3ijJ5cSnPVKsm4uBdM1z2tws0CFZWhTdWV/cdKVeAQy
yjrB1M2RQ8O12GgDb17aGAgTFpjQes9GCBqXvJs1zXurUkZn6DxRihncW0lA
R5UI48lo7iZ9ONAO88r8QOYzr2D6XXI/SQBEZIue/QrqwsQFnER4jIJKSFjK
ZWd3tZBOldGsXPxtu4ybKF8cN4X/BqF+GK8D8BzqiaIt+2QqwUwOqJSIFujF
y+c4iiQs/XPijx8bFxsqdpFgCfOECCoo82TtolkjHdizWNUMaAoLoBTYxLKc
HWyQzg/1C9ROVcv00DkaLb9qP/Vvs3aHv+7zoCgXLnqAeHiDQIXRt+H1PaeG
BkagBM9AtE+bp6JgueAXDEuSzcc8e+0yFxDTMRhn7ObfUJI8SjRw1v+43px/
L1l5dFPcCLqT0j2QalF9YIkTh/SL69LP/DSqcNT1QSosW5uCL9yPpDA/nEhd
f9jxzks7Y9dHZoIh8Jtz/JjiDW/IZpIiJ+icqOFikXu0ue3YEfTj2FUqLEzE
0pKbkg7+PJAIUfOQddwBYJ1wEldrbwX7Gfs0aXB0vr0//MKWZHzvJXY6K+Cp
Md+JbBINw26YG2ZflxQUabwtBs2kEdXGq+HooLluNY28cQZQlclUnAgrj3/N
VF5ylvNsL1e2I9U4DttrlGb/Y6Eie7QcNqvGQMd1LU3qro9Z2BeHMDlz2Kro
6c2iBaM0Gt1cdhnmKciOIHPedTwxMP2So5/3PThhii1qa4SaigrDzqL83c+V
mRXrm2Qtj83y0bPBYrs5V3lAdvl45yV9G6G1boyOEqDN/iJWOzH37wb1E6si
D69JUneFi6NTmGK8MHCc6W/xnBfxys1h8eZfYJJbd2BYsEVzoBZrnS6+k4v4
7kyI+ETV97ytMfui5GWu3i3tPl/CAiD1rqC9+544m9KRxByX6g0bF+QehSDE
Z62wjciwZsxMX1fzJplzxLmO6JPGTX6BnqW7raXr82LvGV645SIFmgy+s3Zu
rHNAgIwcf421ayxjkGYJ6Voh5xik46dMaIUvOL05915PjwAEabAsHYSXg2WY
MlF1Kby9W5lB6rsNr3pXZeKl8UXouAel6aliJUPknwbzjXhxNhn0yA3hAlms
yyC40rXjzI+jjWAuLYYNEDRsg7spS93gx+DhFWmBPAM7nNiJeyJut2W96Jxf
Hz5NiQ/T51CZbAO+Ayw9ykR97zYyiRSEWMaXf3CPJ0rnDTa5A2ryXVOnY4FB
2iCsXRjw1Cp1Evyq1/0Vg7xw6Sp33iF+6DA4ifEjEuvBgMuXZlda2ZzNx+87
Yg0fHpXuCdShRbwcsSsboewMME1HX4J5sK/Tqw18lLUrWBGArKts8TK50bnZ
jwErGTpk9RyHY58n6Ha+9XTKGQ4oaSQGea0mqLW3k95NL26D5dwL0PrifHYx
2xcp1YrsXE757y8q3/Wk6EdZDJJeI/RKYDD7QIQLkrM5DBMYNXUZB6VmNmwg
qDX2t7XvMhBiBFV+Rdw5BKSMnjXVLODWR46lH0ev5CCWJwZa0Jhryv02uIBU
ODKp+Dc3+LWed45ErUaPf/Ytg1s2Wp39lt9OzQJIkTRzDQCYqsqo3CuwBdVE
5ovRdmjx9YEg986t56VyGM0iTdDqKHpSCte1iFwKidFivE4r1+WFdRC6XsPA
MbJagO+Y1eUoTSJ9sCgIf0jcZh4lXz1ZN8xNuaEZ9HS6OKk/rIyZkeTh8Vml
R1MXFzKlE0fTBhdSEsmFlZlZL8k4VoUFVStBoyV2Up7rmn+Lby6G4y2dwXQJ
jmhG7M3HQ1QKbIKBh1e9RJ8HUy/o1mByUcwtINXOiHA+A8P58HbyKJsVdWwK
owhUhifGowqUpgbXZ0E50m6niFHrDDPUdrimZOlSHRVfHpVIlVMgvnNz3e+6
ca2TMHkFyCqZQNk4tIvgm6y6hAC3OUM4+SUTUmJb0UcU+7klF0Pw2TdRBdS2
UQD48+Pel1Er94K2q5Ie44528xBaqHQfPsb84dDrjYWsMIlT+y9Yqp9zZPFj
ekBiZ53Le8lLlciJapFb0PcpJbfthz696UV2csjLQI8QXjAzlBcFp2P1xJF/
dwqm9VXUHruK9b2bHEhBvyMWI2/0hOdBexWiShi1w4zg9i+MG7TenDVo9pEE
v7noqpL2eoSHgL+rcI8d07X2TNVOkuX9SZ5pDTt27wuoPkuA/yI5GtrNC8Pb
AX97NdRMU6WWs6s3aZsFt9pBFzua95NPNK0P0ettTGNLZ6JqaobcDIKUGIIz
1SiXab4RkD47h4vMznbLuzuvOAbM/S3COJ4mzULE/8FfhqpCpSCd/fXiH4Ob
z4ANVFpkCOGWNuSrOg6LYDbMd4uFHl4oHlaX6l2bO/Chi42EPQoyJxIK8zOq
I/yD5tpJOyG+g6zphYg7DUKGdz2ejIn2d+s03ZKSWQVGOUgz6+7L0ioRQ1Eh
TmsjgDuCqPxxXvw4Fwi3MKM3s9IgS+qvAhILZAymKxmCu4JpLtDM4sQpsLIy
XyQK9a+iAprPtC5zSHZYnXvlWc/6j4dcwdEQIg52lg5STYifABTL6c7yBors
s44kzBkv9CnmThHwOJs1jeuHe/+lV6mBaXaKDMCIX598HIpOHqkkRPJNkFke
VhYJKvwxr0YVnFFt9WIWwhHhD4nfuV3dsBLDDvfEYhJ8gIUT81ruvu+a0F5L
nEzC6KU59qy+DYDuTTUeiFjK2YP0NOv54KEvMqKuR7iFbkh+04mi7/XvWX0m
eA+EeptHsAI6h9aSVBbo5abk25CDbJDMt9wFj3n6AlL9lBzMNnv0rHVhxx8V
mgbd8/tTRJ0OkdWNFWrh8/2wrXRbNCZG+E+Pfxw4c+mquHxVUike9gy7d8TM
j94ZMqT3lbYA0cRX5DGnRxF7QU44Tg6tAJeq/IhaSdYPisUn5XZx6z/uT8XB
HmTJ6nuVd5/9KOAzq/4IWXSavbW0hYUloOsxJXj+hQdvuYAVq1JwIj7iQjgL
CL3tirjD/zhee7YUfXGKX6tlcbpF/85Gyk5grrOaMyqSoxeFQhF6f93ekJvO
eSRLcX+t/nVCSMnp6d8P187DU/I1Dpd6LVyN00XgtFKNyOAKRmLEJfuVLnn3
2eMizMbHB8gQMsLuqz9Lb6BT2RRx1kbxlvAPE2CB9Ht961DOcWjw1r0XaG/b
Y5jrQoQOYF39xmjdf/tJSaQEB6s0pyLA6TBCpSgiH7C/dc24mTRy+qxKcp8t
p6ttRwxpamB5k+m6WdTOzcUm91zt1XQkBSs76++nb5oFNA2jcPPkxXRbaNTF
6btLY3c06TPEA/2Cc9H1P1cVFqvHW9qJWsGlT1VoZ6Ov5oJpmHPGIzKq8Hts
AsZx7O+H+2qhG9jBytDyQWr3ZIV62PQu62z24v0ODWnFhU4uRE7mJNNr2JtI
1K/kmJxrD6kKNydZnPlA0n738qcmr5Ite2o3fT+TUoUPS1cRYBl/k+OK3Hhy
+F6rECLvfquhYgxphzBgYXm/HhP+BvbX7D492bYICjHmb0F0WA7brbs8Pj6R
NNZ/6qeEFxKrxYY+5y2XSMrBD6/4AhU1Tw2pAcVeCwkS3qB5C+ZC8V2ogBQU
xFPFLV4WR59t3T7atw9+vmRZn7zStcHy1jHKfBiz1EZGA+L0H7Y9SpUzGqsK
QKTInryCaADChJETjBDXoSjwf+assV8YLpsRC4LBZ5PhDCb5LuMXz8XhgneA
SW68fpuMUPO+t7AMyRoIFkjz3exZrD8mrONf0P9X6Hd1dyUc8HtlzZDZPClt
oa/cxI3td08dTobITDVVtgM1JQg8GS+k/0eDzjbvV+yDnDKC7f4zcFLQYZA6
IuMRp61kzoDaRPc6hQaugct3gm51LSsT6N4wwzrOJx2CDcm40Xf8uumrtUzK
+o5tIPnXtrnzDDWRZnnDoDMgNl74laUA/0kTEYWnxkG166UdyLa64avpdCrp
tGxjzDm7dFXFd5s3KCHLn5ZA7RRFD0TC236OZzwv8xu3cLNlsc7t2ERGAdJ4
B6Q+YiRlyzjbbokThCH6518E+t1zgBQLyYGkplDnSr6tnZq9S0s6m88yOYSb
9fG5afFGpqpVRqMNeHTKO6Kj4XRJZAlLEVaV/T4FZyfW1LWL4T9nKD7htfQN
RRzUdKVr0bZW/E+rr5h8TOkIO4RRjpyIMSbfPmibP/G7Z/k08KXKbQA43Z/9
vrUPnwKP2FluuzdNCENYre6fpyS7x3kHwjQqB98qAacM67kH3N/7OwWHbynh
AYnchxOkoFTiD7oElWnGCm9U7tcn2rFX1wtSW9oG7WcZo5CWExsEUAaREb8r
tpUHsKghYKJHO5SRfnStseGEP2g6GZ5dscgqv2gtZWx5ASyMk0ACtNy1+HuC
40E3HBXH9RHbFTKR3dtrJ/GPUMTGv6hFvD4L2nCc2h7OFY9/4s8IFOVVd/fq
gM/soNYsBfCCEAE5gRRbiv3pHwkRHsFhx4j+jv3KeHtygy/Sw+H+gfibwsFP
cJFbhIY9nMHGMfG/rUJAXKZvK+peF85P4bfGxqzKPgVCA+haX1oAZyX+x1Qm
Vy+SFGqUuDiTuGqGeN3tdaDu9ePWFvmphb9933wZgv1pC9m1/5YwSZfteVX1
Mn+0vLoXKeKDhDOkUhYqT4kFOwU41Q7S20K8MBPl8zebnF2Me6lbNibjWPfD
b17M1phdDqR01Hq1lcCRuDWy7jjZyCooYgXhUCCWYdUBCVOWWNGYP7TWvTAh
E6RnM+pAasZrk8xvguOe8pyWbvkDwCRzzjZpaoW0gdALNCXrZf8bIHwx5Jvp
457jc0DDpCcNH75A6/Fl6iDvhriPz6Kh9x0dMLoEslkMVkf1RPhBNAyxLo5s
Qq4IPJ+bjlxTeDWioxMn+yuJJ/O57gDydZMmfF3Qq7ZeR6Zi0zJXxAX8C0qV
3KMtGH1hbttVwNv+KxXTuKpyHSN198J9ZpFM51jDJUSQsyWGUfd0ngqSKUqp
gMvRPPaU3Y/6kbrZBsjdD803ARJz7E+B2gudeWdacsvTKT2H4wb+brj42Isf
Ia1XlPlpOJRofGjzOs+6sCOxSHe7zChq6K00lI1y+GcsvSfirwsQQMOrYwF3
MV9iakMbBvga2Fnf28mnStt8+sa/C9ORPGat7eP9BWYhOCW+gRaG/7ZYe41o
iBcgNX77xKCvugQ6nw1Pmrsrefx1G0bYPIEvdlBiErCGMLaSIWvakBSCp9nK
jlR7DWxzLPt3hZvsn9lG/37Rvq9zB0a99C+av3FhFS7I5OdOAkiuiGd1qaIa
BWNFMeje2ButsBo1jjzY+aStwyX1r/NgjjBEFSf/2JW4JYDhp4tIPL+JqyJJ
dEvOj7/8jQ+5jJSMz24s0+7cFCX+OjH0/XRCgH5EJ7qsfTDufDF//7YUN/8w
B4mZhVmJ9BBOY6UPtZolLLCaZJhu55Yc/MQ93c8HVNBf7vTZBMzHDOMzjIP0
6D1xF3T55AB1ah+VTDsPdEWSrzgvve4DhvAv50hjv0cCHNbvnqqgms47REw1
rSjFxPwji5EG3KP/Q7wwVZSCc98S2q9/+YAbEXoSM9dkpEo8EkzDPUq4tqSk
njq0u+BL2HWSo1OjlfoFc4c7D9rWmVmCmTzEt6P6Zx9ZjPmRxWAyVxZSfMxU
3ro+OVmA/ORow5k6RYTofy/qsWsGCDMPTUAxxt4BU6JCkG6cocnZ5rzGlRei
NezPwKVEJocsXuXw98zPbSrtanm0j+bWn4MCM0ux0spS6cRA50TXSr4h3aOP
J+hUF6n+fn9yda1Njiomz3upC2yO4rwbs9yC/F+txxcSesMVV0VCwtHrWqgc
w/RZHtWvuk3bmxnuWDq8B8GSXKo/NMT0UL7PMH2FDO4bDWeBFam/lvnnSXpX
h1cxPnX1J1su6crfp33A7J/t+im2Jz0g6+44JDZaHmiY7mNN2QyecyVMauV1
h0YZ6tN5ObSPdUduvskvDonEfS47yJPZ6tVhswv0fXkEcOp5M2VF2pTv0ykl
xOn0noPBNncf5xpg/FqUNJnAGFFEAv1zPyaofzfXp0r1feTl6+MpuZjV21Ck
JgheaBGJJ+0ZCp1nUcEtSjRELF9Y6WLtLioNl4OlIUNO7PkcbTfmIA6O8FOF
dyinZFS79CrSd/gfww6I3BEtTmUeZkHCr7yw8gl0tdJjWrOjbcq8DA0jQu8b
mSG+kWzrokXrIqt2r99dALygLDvJThuzsmqpWkhwVQtAUVWqTykv95EQyhDr
ESfNoK7MO2qm7ynyUefpLrsWd+zoxeXnBobl3U1EEiIN2wvjh8sivgLg6TBm
MPhvL3fGHHa67w4iXuB4Q6U3tvrcBqPvztSpQm1nHQ6Zi+W0XAHupod+Xw9l
jOYfojvpa7wtxmeDk2gIzDnqAWFAT/KlCwpxy15rpdzz5FXdMM9vLTjjA2oZ
z6UMqgHklFIblr7rdWXFiCR5wBwtR9Ts3cKSjgZ9WtZ61GdERBONVX0mJJC/
kL+JVqS/x7VBMm7DNLbvzQfqgvbORujVzOBDA/fo+pfhZy1MlxdqeuCyOQJV
DI1+3XxNh2uM4zs+pnXeT8d7o1iDAsWxRrv7yLuYtHCrR/F91zWPmtifKUW9
5Yo4vZiUHVOyFBzurASNZ5y7071D+KnEiPtRUdvjimsOQvmuYpTSM7pMIrxu
+lyLo8uK16XPTvf+JrTCxq0Cud2GXujsvn8LoD0ClOc51BwNLRoFS5AURxEj
rx2rTnurNCGD+LpoXehTOxvrfHax5baqPl26QkP1rJs3wlFWPFmjy5rUQ3k/
HvB2QhpYEee+2Szg92SeT63AwpBgP5bQm3kWEeEssa/+isMjuKX7LPfgStCs
ee1pfmhmqJOtwPhZErNJy/JoTcex1Hojq/3rgN/79diVpk23mhIKUmTcvBm9
iFHbfaVIb8Ig7WFF/elIBKPfIkE9ZphXetiQt2d/KGTxRK6P5KTCaAQiCko+
95tMp8crOcLKnMIhNKR02aVaABnmepzHjQzcK61OmlbRwGe5lZXiU6rjfZtz
wrAEGttxgbiJv9JENU4fervufpsMatlcfTWFnfExMsEuc12x+OuWxdg3sgKw
aQM0iiRHAoouzcgtRghUR1mP6vJLgQcFoP86ZeePVQ7hwIw3sCdp0EdLt2KN
4CMYJTlBGy7/vuGKr+3QscetSJ+vspPk5/iViUDbUGoIaAJc8l5kT8EwJuW3
5cJuf3qbrz01tu6EkVqMvItKcZY77pU07wL6qBoQsyK1AGmbiB1E0R7ypxyh
z0ayMgXEuSMi722L34n3QeBjJlPUm4WGB/pnWVGOG3+pKh0ttB/AlIERcJXo
oqlOZLnHJDD7ZYSWIA+LXy7UG4ZNNJjoUSMUkIe1rVz1L+aOgQq+XXXAYtu5
nwnS+6ngOoxk26FRc59j+q2ZVXFBRCVLxgzoFIi1rZH6kO/UUFhb4UoL4sGK
aDbkyv+55szuoevTBVSX3p+4JdUz60J/cXry7A4h8gjSd2VsPBSiluLvTQaO
+di3fbqmC4lRTNM9EUvDT3cN7tMx+Ld1lntOuMh96Jen3jMcbVpB3AG7pRGo
z65TTPK3/4wCwUO/06rjkdVjOp9WrQuJU+ysHLqVdKB62w4jnxT4uWknzWD/
WZfBdNcMBt0PV5fkVjqkT6z2MVH1NoWmQYCQHnSgeIuu/MdcB60s+1B/JHF2
oWSYzULki/CRH0o+J1aXFAfR924XzPWi5YrpdrFcjWgwvtJf/XLxyUxwx+xc
CAqM5Wj6JUWbsgo9/MZnbvE0n2Za7RCsY6UpAZ+UZ4dtijzHmcl9DfWf+geB
bMn8+UGp7j8vvqYSDk/tU1+0dWWGIvSIqhHnTLNjZAsY+/X47jBO3p1dsYwe
F84RdBO764JoC25i6944byPAnJmY7EfOcxjaMF3TfFK7uCsN9eoFArryxB4M
3wAgMi1IwgvEp3PXEv5B2aIG7aBjaVrQJRJPrda9cSJrRSJ/IOGxtBKUj0Rl
RF7iGdG5A2eZrfF6J+wLhuOLzy7+4B05BZts+VIe/4dDEmB4I6nrYOgJiven
DL517eYSECCzf90q4gsp57qSBEsD7z/ZRBom8M1Ena7sAadYn2qUPl5X4cFk
1sVhQxBtWSLZEAHwkfxDO6M9Aj3IkCUkjo7gdAt17XpPnQ4Y2mYjUYuN/qKZ
palCHfDhWZAnAe8mGZsc7KQjajpdN8GmXCC6Gr5J18tPmfNQvJniad4Wwtpw
5mJo3RBV1ZbeY9HDpROEotPfTfgU0veCB3YRxlsvLLwzgE3pV7Flkqq4PTm5
BblxwFLnz3fZ4dO8rql46EUs4dUjbLJ0oNRH1pB7dAZnJmVrQ4RnydGeUtXq
iIW6gJFX3G4kI+vxOVti8ua+2Wu+OBJ0w9swTCCHIybWoGPoIrVjl/Zli73f
wsosQHFrk98WGladLjOZqezKG1WeOlEm+l1m0QOjyx5i3eVzK8f4400x1W0m
UWIt3CM/pWvTN0dSWAeVkPcwLSB7rgn2jLVx5xLZBkuZdfIYkth3JZOrI0Y9
Dm/SPg3giQEXhrXQJHG9Ww+owwYzF0HLddN0nj66dilBq7KNAiImKEKhJFrL
mw+UU6GIFzyBGoOpFrRv8NOosLT8kJY27S8tXy9KMnlsZIyIHvoorhJxfmhJ
h9XIedjA+RjHV7hU7iM8HM7sFsvEjU9VCYhLl5/EgoGFZKehdDZLvTYXnN/x
UdaOOo6A27pd+LizEY6m45eOdmjHDlFVyIRyqdxGvN93f031GBefP/TJ6yPs
E0bMx12KQyGi+9zHVZJQEQ7CPoSm3IwLO4HieCxy3aHt2Bjr735O0nFlrp3f
OibAKPgI6LcFeK8YsB3EzGb6BbFUemya0am0QErWC5twE/wlXWU5B4NRveJh
UKV76ODeeucJwrUc0bscamzDqh8saEiy0H3f0eFbyZHf4jTKlYLQ5tV0C/N9
KNt5uIhUeIu+nUiwBhZOBf/uoNnsDiHyC9jFcdjmuAtrlvJoLtPrsEQn5XCs
EUEAOCcwpWiFjw8/ZrfLiBttfMZSmPPoNvLsBRXJo0ftxvxaKZujuDBSJp6S
NM1mJ/XSMyUSxCrzI8VGfjKornBZEwXKWUihx2iApUDRmNXrD/GwGdm/nu8M
dIIzPKQm7JQXwHyOwT8LR8Oh+XqR3f6iiDynshU3dYuV2odetJhziweG/CPW
tQjYb8JyZsEv/65Q7oiC0H3NIciFqknUONE0EfGdxySPzz1aNhHLToZUncBd
7MWCvoqVwOyj0ZUEBBzqaun9NFj7mCbBlYZWuJxt9+B48DzcjHmmK0JYn+Gu
f+6rkFYSw/BvoKqutuXoW/y1robcvSEllEG0uBXEW21d2tIiaDo0xksN9O+Y
VDrrQNQsnUss/T7MiRLSOc6MzEKb7DChKeNfPo0plfo5SUCX+tfEsZjwZVSF
NJtX9Lv9JnvRLY2wkbSfAzvmgLeoqaMGa6S2wP9KB+FCDBdvEsH/5OLHOKRt
JV/GFXByDT0G6Ov5PIuwACY//PjzdpSNM3ZTAx1hdr2VLqh6fTqY7Ur4ecWS
sJcZXNMaGUp/3cLYj3/ILYtWPwIuuYSh7Gg52t75SCcyrwhiSnsBeAFyYveR
g3Bpgovw822K9lgBuWEXMdhCq09K/kCmC2kUVhmEcu7t/a7hHWpwzhzNGQZI
Yh/5Gs/I/83Zlrn2blmFcoYTc6x3gsPywnIRZUlBvxbIj9md0xB7MTYAQKCB
HSQmU8aPxCGSlksggBBYMSkPjk60rzWbBa50AAtDD6/kPZAjZfRl+AxEUZcQ
iRZtkzHPzTNkCnJDmeNfmJ37W1XYdPQ2wAYiCJucu+Bqnf8G/iem2M0GUwkj
zjP1TO8r5jper6QC3SJ9R/psXWrCtYkaB4Lr3/CJJSTlAViVIyPosgQefHdN
ZhqvUFQ9IP5iKq2JfLH7EMeIgu4/lYnTMrxYA9gQC7sQO/V5Tlnn5MzELtyR
kjWu86LHdcmrWUI9UxWVYiLCRQJsGAATNylik2xYAmS2PKJrtKDIYFJFP5Xa
jtzCcK29+Uzp8Iyqv8/kVJtxpcTCqNR2tYBC2p6cjX+JXEFVQS2wk3MRTUzk
AjSN+ZyUP1+O/CAOL4qrRrOQ4IaxrTR3Htc2H/AGC/m+mCeRhypr+ypFnWjU
xjlxCZFKXZN7iQCnxWZ6UocVALzcWuav4FfMGDz4t2hxVPCc/mdusHv1hZNo
BouxTd6cNCE41qSMcIQ7FKAZIctnigsopoPcnNzGg3uDY50/LcX1lxBlHnFl
s/+6cP9V48XZaBNJSreyYwUf27zY2aGdYE1NmKduhkF7Pep+BCR6FZWMK1LO
6t7H4XDVKnpLxmM2mE4CH+/2oMKuwtntmTtVoobM+mKXpw8pzRhzKAbyUFVV
TWqgdjPXKoU3CnHeMF0QJxvE9qRxHzWjbM82Dp/rnAQ1KnD7mZ6iUrT537K4
G2WhKtFCUzdc3B1ejdzsxz/hqnxk+beclOPUr1JVJOIEPKe9E9XDgiBbSz5H
6CNaYL5x4pd28HwHDiz/qMdbUM7nx1jJdjhsVHEafgx85rNKVNI24kEAYcg0
Le3agg/6nRtITop/iFV2PRNI5ukTjVu2sof1QIkVBfMr8T4rv4x5g14UGevS
lrj2pkoodPiw6inwnNSinlAQK+bwEyIVcE4GKIeZSOyydhfm6AvtFhNnrCGt
P5Imsdna2oKa5vX6YgFM/tGjlzDGBwfzXmnHyBvgY01Q2dOBetvvVknR6BjN
Ij9drwJdIjFe/J903TnMj0nRjMy9lCLeYrNqtjh4LrqyC77KcTKyWN8XAa5P
HJzxiVe7l78I+3NT5k86yzkq45axyOi4U56wwPwed41wympuc4p00qc6N0np
x9OReji9c+5trj4yXLdhc8+XTufjVYdAhp2xh5J8s/dKmzLryO06dYDD7hk8
AsrLTjr931NRsqm7zHSZ2ddmcamFn2XkZP34f+whmlguYAlh0c/r0OSxzuan
63n1UJWLNFuWxmUGsiiSSGZc5ydpu/18m3uINemmBTzuIp6LDPRxTcM0WYES
KLcU8I+OyNrZ9GGTsBsWoh9zdW5kaHVwo6mrpNBEs3RCJ4ms+TSfclROPWRi
3kWuseQvntUFx9Z2ajk0pp9hJH/CqWpAKClU4R0HDkBHXXe1Xeo7iPQsGEIX
E65Wv5sv+fvOtsuodsFrnNWFzpZI1n0QeGHiRyrUiCuJfm7QE+rTWpHeU627
OZJ4Y/BOMGD2EIiFiG+fPGCRStzwAVlWHwFNlLgEcHhJeK39PWoM4GjDUzVd
BXsjPEf2BD1xJtjZ0qSI5iSz3N+Ud5tbr4m/TSwou5m4DpCfKPcHZWC1wib9
ULLFR83wDEZCikkkigjImXRBf2/yCl8KQIGzBG8WfjFtZVqzHotKv6lFYRb1
U5ZHac9eX+18pbS9IBBhis6538OzTE8EHQDbP3zCTi28qs1yJXW915QG+YSv
KqPlV9w8hfIwrEMRbj70KBPmhnr19QZ39ZM27noP2d8WhV09kdoNdzBEgM5F
RPsT9gDo5rrWaxntpcBnVZ3R4aY0N3KgQw7ai2I4MA+/ip+T6WPvzwVJGZTX
eGoOOk+yPHtxfhbkmagAWrkQXiB4o+HeV4WNVfVGe/rib+U4/gjsdXk4yNyz
yXSIQSMmFpf2iaxRPxUfpC81ABRp1QF/HtA7ThmklGwWbwuDv2kDRO/cfG2t
wL5d5SpxnoN8jY88ICelezQq03YmUd4GeKPj4Ak6qDjyB+TdpaanYFdYQLFH
07j9tJQlMy1Ou+8mktuNLeW90ga9gmXsomrkoG6NSdFdiPnwX1T0x7bQ/l0a
OGjobr0gK3g7EZ5XCj9oxSfVH1uAaGmxyX6kDdSfDst+1Qg7qq9FUUg+5eSJ
qVhHkUdECUdvRvKygALHdKdnRmcSRDOB8n9/AN/0TmBQFkiJOXbUA0dXdioc
+YRIM9KRnmF5g2+2c4VZ8uy8rJgW11oKxRT+ZVjVyA4TyKmmEIcVOPRMuhhR
8NMz/fpyLBMJblE0O7XhH4zP+ciXjx5yjkca1Qor8L/87THR44AhqNRuidnM
avdxA3TlOqWlMILyAnSdpkJWeUy7lrh/hfR0bU4IYJyYX6EpvIevN607teby
OUuDdZL2TjVd7ZMpRpE0FdKuazD8DUS1PcNx/5llS8MHGv0AFbf8ud0E/JeM
210Ouj4d1iDCxp/7kwXKwygikGIVMpmvkIT7/NXD5acc17relBL8m4WwKkWW
nxm27oVapfUxJM84pcJO/Z29oFlc21WA5uaopqa+zU0eVloh4epf5718CnZd
ADyMhz2E6JkNKor2nicMRSwmH9dpjgpG0IIoH0aSK5zbx0oBgArJxBY4FUrI
g99XkrD0ow6/ofoDOQyb3pXIMTwjbmHsEOylvgW5Q33zw6IcUCruvG6qcLEo
/JhvSkRTxeAU4R6v+OttRrJGYzNp4sobKrJHX3B8cb5u0aCEWQ8Q9+rwUnF2
rZ7UjkswBWG6Ecxh9qAx1AG/vxedYsHdQbn0c+lSn3+YLcnOseGSoDUof6ky
ZograpNFEyKH7BFgYuF0/ZvRFyx9SZVA26psRKwOUhjKQvwmjEhk3R3+yQ5N
q6ab4Sy1RsSS00SMd9GRv+ZpdKnS/YSOQzfuD6kcMjwwDb153ffHMorDafrx
BuJePX1DniAIwQJeu9IamgDqbrRgOGMwt+0hsPhgTzTxFyUiDbUt9neZmdx8
i47FYIdneS7ajtMYg8Jr+MgtenIigkiXHQy+3DCk+/ANFg6dDXKrSn/lauQf
tBLi6KKIFtTVJ9uM5q8bXczCPgNNHcljRwb4HuNS+PgPEJ/gxv07ANB53uUS
jEabiOF42I6DzTf2+ILHFuZ0vXDBNCjFtzHNAWOB+qHrm86gJ936bDf2YntT
81OWj80L0H4LrkNWvXHtcEMRPXvt6Q8r/ICw9QuK8ilzzrHKijOs2Jvh5uv1
K46ckX+I7fN5wROuJ8VlFTDUnX0jnlqV4LmHILGo3epo6Tlq9HcFNjQYXmow
z4bYqgn8eKnqfal0Rua03YGzyvP+r9nxUZmQ4n4B166a4Xmqa+TDcms64Qwc
RyTOiwrve4uv759kttpa/CBepxhb9+UYB2Tbt/ivIDMYNkde6boyn1ryAiXK
Zu1gQayYtC8GqaoVu0TAVi4Cdt/GH1HKkPER4UDFbz6X6SRI+D9GZPz/nwWQ
4FDvUFaxPeeRaClKIhnuGZdfnTIgd/9shOOYip+wX3R+BbkkRlzPZaVFpxXE
axonYmAXvZYYN64PQXZOPKy3WlNH+D+LeJlzDzzB+wdm8wD6sfGTZUu9cE5f
2pnPbvX2Hb31vqN3w2Oid7uhS+iiniW68C+r0VSjA04EkFRAJsU+TpnTUyCl
vWuKaBFych1ZuPtLA5irEPzT583fPyfdqqouUx/ZptK2hhIXN1aL449Gp3Z+
AYln0Uc6bQhmZz4xq2KYVC+zXhFS6RK0t8EPfWJclcueH0LI+fClTnCi/bEn
vXdKmFh8j9fTmE6NgLMTCvXoyGiTM5HHzEulYH0RtwTuHU/tlQL8oKbHOL84
wwClT75sC+d+jqwkwXdSyu5beYY12rGBMQTfGlyBHeMB117T9+Y6SpsNIbk0
yqGlGFh9grWPkUcYzYNImTuqFKhcHKfV0eMfUFW8ZPaogOk4LNrRm2KnsqrR
lRtRSc9RuSGbSqpV/DEemth3crxRoBiq6VDCGOwA/6YBa18kS1zTwocvb6FE
JaGA1XQbOOUxaH930EQUhLiZ5Waq2Fc4a2JQdWhQB9RgjPvnIqlRImy7iAo8
9EA9/vW9w9glUBFPym81cP0B0gJGoXi5leWOzu94avQsCGNmqLKUKim433mo
8HQo98NTIDCq+XWLlRtT8XOwDWu7Fa7EvfAGOzDToyZYBkdV1TCLRY4qPjiP
acwmXYscNtQbZAnrJds9mxnc+iAq8QDFRr7SoNdhf7XRhh3aQZIcz5K8vAPd
K3kvfk2pP7XUilm06aAf4rEuCGbox5VglbENjjMkl/yf1+rIrim6KkywCvVn
drtdxqSzjyja9A0f85VhGFqwEFiJTSba8K9BMamFHbYXRkKijdupxdeRrs/i
pu/pabxYFIi0ZWlcfkn+MBuG4p0gQ7QRVG89UcXUBIcD1gDmM/vusD0vRaWU
DqYeSO+2YSqD/6T+qb5KAzz/edduSaSnhdfZByG/GHyXQy0AHqvbRNSJTcEg
14gFdESosNzK677pFQvniOpzTkNpro8Z9p1dX7uctKqCJC/CBxNzyQ9rJY1J
rQyqzOcP+/YOnyNkkYLfw0A4mznwSto2nS/Fbe5Fbfx4JAwSgUG/dfyWIkiD
TEFqZW/fYxoSLIFr/GKIvsVxXZTaHsSInXurPBJhEzYaRMcQCMtV5zMhIL0i
gQSw1V1SqdBPoq8l+uHrCWxCmcDHp714Ei2MThvNyLuODXZ3qGiIeLgrGkaL
KosUyPfrF42M0HVI8nBlLYtkq4sdbACHNe1BRTHGSU35YlHxgyMECo2QHfoj
+mw8bK1vxOgAKrwGr40IkVXd/EJmzr6cU/meb2aBuNMjJ1mgRH/OzZ/3EO5P
Czu9Ux4l7RZB84S1bodjDGG1ferOjf+u2iJtFCeVRJrXWEbop4b+Mr2Bdmgz
1UR/b19mfYhtSmfpiImqfnBPFJkhL3XcfJBnfZ9o2gBeOpJ45QsoA2UU+tyX
kTD9uVmgLxrocP7rEf6EM4Xp6JLUUdDsIQIzO53eGsjOSPiRvZ7owchTw8vL
Mzo/YtpNjT4YtIrJhXzMghxStnf+z6Jp7I78e7OPubSGO9k4ijjK77GaBFhD
WRARlM8OiJWsBR5sB6uF+vduaDKr5lbhBX4uirn1wZOTD4Ee5E/up9Sf9Jqr
si8Yx35eLNNcqlZy5lhHX+vdbb3GsDsfvCYXZ+e84+SLsxgritKsPpXTUHVr
iwzfKT9n4a3BlhRmSxCuINJ8sFeVh1MaWy/onbaUPkMSue4vLm5hCTcv7Zuo
MkXaZ+b/7Vnzh/bYQk/AlA0Adoy4tAf4T51zTPzKzw5bRmcuCfKpZ4gadep4
rU7jxV6exfGmeNY3G+QbThdxuIrZI7BPS43pJ6KtWmbkeFqQiXo5JJ47Ap8i
+Z3d1D5+7IfbOmzPnBX+Vxx/7FGzOGuVVmsbyt3F5/eEbQQ1s5CiKF+34NRc
FXzFsIKOObexikccEN0ckoGy1kET89r+GccMB8KrywEpA5GvMz7h69IkS0AA
ZsvCJPIf1RlkC8G05ziNHrbRgXWUUJL32uR7oMY1vC20s/suj4HsW/Eyl7Fd
1NCJG9hCDbryJcDKvQao7ZnQyH2dzfhz02inkJHnincR38eBGFIBBihWTw1V
vgXVD9qnyAaR5gp8M3TuGobvTZ2ZcTmKB+niUEsTndBxQBFRDksNu3JFr4YL
9v3KmSZ1J0tfkMAFjevhne2pnYdaBqJGDb9dqvb9+hkSoL1AKYO21ktHH1LV
VfiaPFgW3tMJQ/AdQw4kFmP7E+YU16bKB6RIOyKGQ0l4UwVegJwQaZhHZ+hY
iuED7wApcw7m+KvosNO0uw4atysgaEGs05J0652WiT5n1WVyMrlEGMnEPHZw
LoWPH4N98on4UD0FADrR3MXm5seAw2FKAqESCBTH6d+5f5PHJDyK+s2mAhj9
nsQOmgoT9LFM1PL5piBLXeLWZXV9cHov6i/lJ6WLjM3Faudrq7wxjV9BV7Pm
oDdp8XPxh8NiuAlQzkA0elrVElnD0mP1tqkZheqqiNMdezB9KbHIhRPfEzDC
WEOFyxCtnwd+IRXVFWlEa+mHseKgiP7gwsstYkx3+A64bwWZw+iUYcLVIxE7
E3/OH8HtVPqo4AbwS6vqkA0G/NQimWwowjpI5bwWucfsTg5VrRNi9BbligUo
GVtRycMMNeNj0xibsnoExhBajptD046DPdXo+9nQGSzktAccLlvBJWcbcedF
ywCjYrdf8Slr4P2ryTsLltluqAq5XF0jA40SKNqYJ3hkBZ1zKn9WlsJ7w0Xw
NzjosF3uiSbvTnSCCP8I8+1UV95OvU8Qkm40IIMLK0xHLfdsz+cBWCmgG4pV
mFvx92U+Byhs1hiOBwV0c0Dlm//oCz9Lj9xQoi7ZMhT8BA3h/xOVv9bdT/Yz
M2TTjAxc/E0FzbILTuq9KuLryWE1yLwosVzyS4uCSX2+F2lEDnsSvP+YkwLf
kukSdOnIB20n3EDOMDqUlh5G0UaK8KvOUoIWW5nuM5+rya84I/Ffw8m9PWH1
bKRkk7fg3eeFTn/8nWftIv8BWuOxUO5ZKEK6hpLwV5tDzKYV4svRP8e7ZOBw
0nVDCqlB5vy2d1UAk6Q3OiOfGW/DLCMw+T1JmhTTBLmVLwarJqKe1G/Sh6NR
hD3/QMIA7AVAOfEuweQJP6TXbmuIA0wcPBnmoD5qCnLWnsPRA30o5LFwIQvl
RaZMit5EhffSbvhwtD+NB0fMnaopjDJDlQ96vOxKqDr4TihobPhdL02CR5Oi
14+Z+aFYrWjCMgr9YxCO9pBayhLw2AaPvOmjNGi5ilUnaDu0ON3OGpbgonu0
LeSRTcY++6wcjTmY3ekHfxaAPm5u13kf5N6PZpiVbrYBlAosOlTGzndCaXuj
62W3a0D9C6hhEsXl9qRBqhvWTpYU5gEna6RljHflZ8BoxZSOM+Tt4TZFRk+6
roLcA4H4GuEvIZ0dYE/OBhHinPoE3wGIlN9KIZcHwt9Pu//zShA/HVz9xBa0
8KwrZfzT5K8RXCeAXYkEfibcL1DVf/0Y8PAyPafu8Qxqx72+FI7tPJ9ny7H/
a9+evjR5ya7FeV9P2QzrSmzwHiAw/gMB7FyZBvhFbKOzzjww1Bos/8IkBiFp
mEIQ+qC6QBUbfdqneCCNot8AhSGI06GugyMcnJB6Yg1Sv4hHp02wmab1sJhk
SDa3zvrkx9Q/EashUtSjy4mH3VS5ygOJPTeNRuJStwE92BULX+WilEzFLYpi
aBCMWNhY64MC6cpnVfPGjPTGwD8qxjIci0ezoUmI41n700d0yWSTQ9PGkQVY
clAhetOHvtalkXef20js68U7XvX3p3XJwdZkNF2MaiI8KCaJ8F9W+/ybVIz+
P5RDK0m+NwHQ2P3Hg5mBl1dhXa+xhSrBHI23JlpGlJjW0QBYgFG2Tjgvj3wJ
1LnOur9RNaVZALQ+nlG0sFKwjvhseXYeIn5aRFJWelJeAycQk9/u8cS2/V7r
TnbM4kOhzDZfh2cCTwW1Q8cB/os/fpf8CpfzAT75+O9wOM8IZalDE1Qp7Snb
PGKlQeojc8A8iedZQ3ZaZh0cXR4phc75jsuL62UTLt9hZV8RrNsSNwnApOES
3tG+bR6cy99AZV0QqU83UIFQ+FwILtf0dTumMAJUlmn9iDhwywLbt+nvjN2z
qIL+KnejfCBErmv7K88nzzXJpb8J3C4BZ0o0JWHx1waD/XN+dt/yMy5dou/c
myKZ49E2KjXnb2ipBLqprH+xA/yhchIE8rBMSPNTE2rg/dWyVDbrS2qGh2lx
5DkS3JhvzovW3m3HkrwAae6cFx3F1AB92Zd4HLeybaMT3kZk1CYGpVVP3BKE
HX64wnHqBPL1jnQ4FidROSoiRkWt+/kvb8U4cI1idosSsqjt1j1fovU5IibL
qdSKb/00kPe6fMotkAHiin2cjBc8Y8A8rKIViro4QRpjXCI5dbofx6zl+2z6
pWPgXUKBD5SyS34oW/p8irPkMwLTC9dzmeRnFB/ImNW9D5TOwAmbxKm5PuRW
twoFUQDx6iBm/ygBA9DxscV6dwqh9cvNX2XowsbBpYccgc4rIo8Q8Xc2X81V
+p3OvB5812Gj7z9mRIjKt211P3JijxBEJK9j5oFFvc3MLxkTXba7EvmJ5bnJ
64E38dQjC+muZ8HiDHpAOUFqbZM8u30pvHf/offCGmtu33959hfU7cS+kAUG
o68yMjfgUbJ+nOI/iF+kK7vEyVUoc+I78ESzLRKMHHtZCrE5bMAGu0SlJhLU
VwzHJbkkzbQPyNrTbg/C1gWoQffJ7tuo/wHfwwcYHZapMmDgSs1pa/FL/63V
EswnEPo7gYXXTFIueby7HT4hbvxuPkoprJVWVyVZB2KBz80TArcYkHr0ZSKf
BNcg7JK98YiwaEaVxvuQjuOYU9sn4S1WUrmmnM17U2Hxt/hZu2SWx9i8mRO2
aecTlZQxLWqI6eUBoLLDOiDzh1gqLQQo4wg6j/A1YIj/t/0x04jLukG6BXg1
iCjIRYKwQPYsU+riCLHKXmzwaD+GTiPVHWbVp9RXuRmZuTXP0CKv9M7LlkL2
JlBNHizUlC/dVEu0ZizGyVBiydzPzzdaIKCSC+J1OeOeBzJm34P7Y5i1aDEx
u27XnagFaoBB0TqvovfhJzqoW2FfRuSD3M+djg2K0n9TSjfpmEZ9IHs7ngFb
A7H0C6UHCaJHnGDb8qDB2G8A9bH9SUdNN9uU2J9oaBP7j6kJKGpQg6Mcg/Nm
Y5c2gGUcqqlNoM9n3orhjAlQbZBNapv/y2zHiyWQN+XEwtoGkkZHJMW8hevf
UtFTVv/hQ3nsjkYEyycUQ0/LHpODggVCrePjeeqTbpEpDT1WCftB8BWlmNyL
ovd+KpkFgEGQz8FT80mMVfUfC6udWUS2SATMMCWAfVJHfhQ/MLkgv8F4BxiQ
FTgJYojjHUesQfQeuOYChVlwhpky3D3rR4S+clQUg2UJMja1CjlKrXsNhXQf
GeWPp3r4TRPTKl+pSgFdyiDPu/YxLk+YBUsi4KlxyeYib6oFYyYIK4Re4r6i
ulipW1Fv6jZzqn34hjzvktc2Mn5GNhVzrg3oe6N5wvIHcxocYfLyVrgDZM2p
sdyKsCs2/D243W25ijW4sR3Wi9o2kJVS3ggd0etd1FsDhCvEWsXxWnuyqyLk
3Fiv0baG0inQWJU9UXN1kA6sYRUW16qqLN5Y7IwlUlXSf3se/M5AZOt3AeTO
fsJOtyBbSED/J0Ip7XF/ZQ6IEDQG2yzMB3JsLBosu9vqBB7Bht9JsCkspFDR
iv5llIy+NyUhwWkV5lDhm5piLYUx2qJ7imi6k7HVWYzNN27n6e7XfR382em0
KWf7guSi4NwmKDUiEdgGNYpS7tdG/U4doPuIqPGbF9BJilXC09voYBvEGeV2
KiHW28HodtSItY0QeKA9+Wf+Q/w82Mc8NZRWajdT+qgfby8NlGVOn32YZCkq
oTlmD8tNYLtwhx/nNNByg2W7J1SkMcYE/bqaxC0mbt8kyNomFPOpeTuwxVcx
+5tn6VSPl4FQezx2yCI3ghyLburJAx98ZnirRrfVuRseIYjOalMrIu/vd9kn
8maBnHLyTbMQT1MiE2Vh7rgRzCYoVpy1s6g3kvnPdVaEGYeRcPY8cBL0XOml
FPcsQhNPWoFqQgiUZ9IONte40HU4HVyBG/AI5u05qUbsbfr5gYGwiNGC9Q6q
/X8yW+YgxTJCpYcximKn72CysKrETkPVgCWCvXtQE4WFnq0g7CDxWNZ6IgQz
iIDaS0zUIBLOX4zePn5AWFv5p8P1zXbZGHZJmhHNdg6SAb7ISkzgQ8H0Wu7u
wBA6aO+nN9v5xMr8lK8JHKasRSrCmoj95Gpx6SB/RkwztENoY7YBezzZky0N
oYYeFSejAJy1m3zF50gP/GRiAeRuiVUxiNm9pXo3M8DIN1kPTEh1DFDVQkJf
lazSKdh2lOoGEo/t/7BgZosW4dDMBLkmACw4kWCLtc1b7xbq5TZtC0CTE23M
urSoXcXKBIIihQXIxINdyoIVf5rMZ8+LwA8fCYBJr+ZH9v5YvYOzzEc4wRC0
OBoh6h7XJ4jfINQw4OYbxkgFHV6q5EapgeopKoS49TmvGza6cNqG/CXW2WOz
qKAXndiJlnVCVySJwwcHwlXaCQZFFuyV1KLtLQCPZiecDVJpocP+GLfdbVzC
4c9m+pLjLd4gQxo71ls+MOARKPW/gBdJCExrEvlqUAerol1IeqcJTavE4UHa
3B8Mc2AKttyB+OUb3pk6l7Oj3KUF21zAAkg6NCUpt3t5VQuhBhoCfW5MRGyF
edv62Bw+Y0pfhDxMBoyJ2jYpt6z/ZH1uU1yZBh7GXzAJ8TfqXJ47IVths/IO
5COPrNgnCSLR++55z9KzN978ZcWDJzpGBgfnZXX6OsA0mERYTlsUiGwpkSdR
ascO1QhHURmTiGr3Zc8TTlMYUvL8Bhr8rQpx+Ci596ly1gFrs+bb7r74FjfN
z1wHdfzpCvEHqznTUhhNYQpvV5jH6+56Lp2n7u8YQxmwSFS0iAWgWaAg2olv
338vCWCjE31xQ+OLLAO66wcV+8B7DLSl278D/esU+fJMtqZ/fcCfmg+mQ0hV
D+c0c9Zk8tdxGKqGk1DGLCNQ/JmyYEO3yxLAJhTaksjY2JCb+A0O36slFoVB
8F/ZYmXk/AKv3RzMYnzquAfZDsigGluMBTv35Mz7DeI4P9JEMunA6sK0fKNA
fKSugarRa+W2w/zbWCV+Irkb66DdrtZKb3iPKHxqpTtOh586V+rZiRHa//wJ
MaSjEhDgKMFTUYeGHUCWlymeN6E/Wzgq6Iy42J4wm4vygBkzncqwasOpZ+Ud
dXe+7KVeXx8oBvVjf1Pi6U6BA3sOVgT842/8M+mhEf0MydLyj9ebDNFzEtN+
c/NMDPuOY35AykAEMfQC7qn9ZAkk3Ev+Drt67ozwhKiL3M3058RGqRuBZhCw
7O+NidMwQQ7gVn3D8Cf9KFStKZ22ioXc4W1UQDCLVG4tQcJ7WpW5shj0oTbN
DaTL5jzTjAO2wKtws7mewI/3jImswSoPYoE3nyTfgjMfK1Dghm9hLu0qK68e
C/DDfyulLFjDoH2bXWHnxW0hPgfZW4rJTYm0ry0ztm5eyW3revm2ZYSD58iv
4dMExtTJuqB5MGE5hgBS3MU2bJdPR7z279Nh4rFMoE9JMHusx6C+kXynTx+D
5jTtHTimrm9h+tgJH9QMF/NQGAWPBLSo+9pqhY4gScPz56ez8sK24w0vPyTl
PJtOEHTx3/r4JK+LQ5pxwari+MFeG7gsU67AzEmmmovHT9QaTU5pT9NgrPcd
N0Qu2+3cx2mzc3k9veDk+5mjB5yBWJl2e2HO50FYqD3dDGRpvi8s/8x4VdzJ
drB/q0jASrPAtPR/Ry1dSmzSm0iELSJw8HhvjmJCPeltQ/yCb604B+NdNd/c
U3X1xmNgOykYj0aFTNExKAzU+l0bVRNFLYL7UGMKuAcrLxDE+YOIubPWldrd
by3+SiRaUlI4jqFqx9jq659HMx08ExaEjFcNfVk8rV/MH2iTGkJ2bKJ8M52y
2OdcCQafmTISHAvIGdWNGSYCEug3JoyHjsIbqXVB3jt/d7XFIq6jBU90K/pQ
71ypFaZ/iKmEPKL7zr3feGIS/FjBtvCrwPoNQ60dermE7+wCc7kH0Kie70ke
Nywz5HwBPe9poAuh12TkPCmaw3ZRAqC69ghmwWH263rnwPjnaeIBjUqnJOUE
PudeHBwxn+sOl3itguBwqj7fV+Qs2V0obR1Fk6vVyPxDAuDXvnH9XcIgd/N5
+i6TSe2mZnyoy71tvQuFwoAz0tAOFHdAWY436zSZ8X6s6lstVbWENBfsYhsF
yyYG4W7djyqW6ERahy2ER86mTnbGkvCkKoTPt9b/wDMilSa5vucDys3XPnyc
aGaRgxBJSpCfhkMO2hESdLgN9ZecahE+ZlkgEAO+6Nq1ZbcprariSwXiemjE
1+so1pnBKGiymAcQnVQ5tK6LALWW+7dPYZkHAapMRgyTcIouysp3WdWaXl4e
2OfnDQFOH1Xxhfewn1EeI42kJNpbSqdX7tdQpX54xe4DC8QIzFum/ek3t4IM
0zOSdt71N4lukZf09cr1/7pwfbQlinxhbHsKcMYDryJTlESZjWmMlT6xjXJr
JBPYrQ+vLWyRosO16Sko54EkV2V4AEYTJxAF4gkXOa/TwUoTNy3BcktgTACL
ObeY1hPjG53V22M9qza3NSshQ2NWURWqkrChgKVbzIt4hsKoIE7HuQvImm1n
G4ijcTPp+3APRjnkmLK+gBiAFUKLgkrXP9NnWCUsq3CE0oHrlymBH4QEx7w0
qG27FE5bEj1HUCW7X5sUp238gFPFUuen8mj9QJeMAhgx2yM73NFaX/lqzZTj
5ZbjKKbxQenGiWXX/yguVxy5vabW2s3ZaNozL3HO0CdU2WHbjgclo9PQp9tR
aD1tsXgpwu14NSHdClxCmXXslfPwSCTddtF5VzbT5Ta/hpdznHzGEgr3ojCi
fvhS8ZY6b4lcUS+Uj4WDnx4yAbYvF4jo6bZyJ41wLcOdxlhyf3iAwKruRXjh
2fIBPzftnYybir/HA6/cFvG/tfXckRopHA0gdZjHQvyW3+QVltlqR9meHhs1
qwKKli5GTv9bj2tZJzKrWhhLtswcFyMsM2r59U5iwCgYiw01tI/53q7Zv8Y/
77zFsn45wNONJ4zQjTdVHmu/jwzpGIuC2fIpJXbkI4ID7lrZxJRAQGoHZlpN
8kexc3PTkDozxrqBO/8BfPuQmL3ZrDigpnVyajHrYEYmEa1U/UR3BLDBNrs/
xAlBWp/5mm7bBjMUFTFLwT2DU61A+eeio587uR6lIS8PvTOthLMI1obFqH76
oIeUNRjrBGVe8WKxsSGZqERTb9JTreJapxP+nYFV25OxNU86EoXkZUQeDppr
PkuD3oMkOxZI0fq9Ek18NsTNqBkVYkXJC71XDhub9H9JRC+6CXJ0gvanizOp
H+GJAPTf0CaYmt+m00MB8vLhnHztWqiVnE7/VGwefEzYBmqSF0YgZz3o2yHE
DarrK/ll3lAtS22j94pBe9RSc39NlXPptH9+ET1sdb7xVxh3foeg3Mol5MO5
wuBlS/yR/aUvn+RuJwKg0gXipo9mwqRaz8ImCFA95GuXFhxzuhluaNzYGpfP
mbS89DWn9YN7GBAY7kfgh2u2elbRiYZmMStKfWclpTm/LStBZhGBeoTONIsv
050yZXUyVVKeob0REm9CQVrckD3jYmDALUwqz3bJiDgst/lTVRvNXxpfNdgU
RQKii1NjIJtPEpBr+QB+UtQVlyyhNZIkVxtgBm12wVwLTgHBdX1U9gddTlXN
lL09MUqSPq+Sj8AtcvewLHlnuFBCVcRiWtWB1qoIr89T2zS/gF3JGTIUdjSo
zZZQbR7eme9lokVcivbMrXBx8W3kpdypglgyqj8CzA6WceIqvID3kO4He1e3
/L+WYK76iuWkbSGHwMIVVXDrqm0lh+l2vtnr+Q2YiFze40y+PbbF3xu0q8k4
l7xA+GcBB5EPTOb5JTGjNt5wYfr6MCPek03mxTjRI7hHtPmHvdpHdvewBA8o
PeRbjOY6UB/pQiYRusw72ftJNuLaX6aSowSNmqoLKq/y20ybLc1+1v6r2gSn
97xw4HdPoV4SGZjCKtYuvtghyFNThBD/0aHPMOlNJ6iwt54bjUneZ/tuUN8j
SdaHt7PJUTYJp1w46Hr1j9qQFPxJO3dksfzUg/84kpdQ5l8km9B+yjU7TSPl
4GP2XUFninrnM6Iuf03VTzRy0N3Au1S4uLmedzAZZjNgTVbS3Yl1oaogNJCs
gPj6OTVxoKjJHa/zve99cp21jFwPqZeQ037tZ14bGY6DFtPT/o+rmAhfMb/4
WMWRpcFRQiPWC8I3Cc48DC7JZ/MSV6YYp8AJ6+N2i+6lNDzbZYkjLpED1RsF
SmYkw5j6TphlDtyaqaLmG82C+bnZ0nHwkQVvesr4BCTqt1zuP4gY4HbkzXNZ
wT116NmrcNU1Xx6YpVvIk9j4oQjKtwa2hN3KdqfJRtqoqwch3prZvi44Cqez
7ECoW1RFPkUQEgkGXdEViEVg0bPiVS1aJot95u8wqXGI1NbV3FLeyMdPA4ZK
b6gE7OF1t4PtkwotRxWMkRf98kxsUoa7Ivz4/SFaeWIE59wrI027kZF2/EW4
w38R/DS36h/EEkr+gYqTPu3M47bLls1gjID1b5yiuBVkF0bQF1zzeoZ8ft1h
nWdnhD5rPokNXvuv0pHILNfSDSj5LYxNthgIwyEP/H24vf9p0xOvW1QCsXsE
qWrngThIoGTjCcCijlBgBYThy2jwWAmhuqaoB+f61281pZBGiZatjIN9RTCG
vK1wTBMIm6d7SwUL6BmPmhPKwocUwJPcKLtFaOJiBefcDPr8NWKD7Qg8kZ0z
LXpXVUogwYfFWxWj9f9CWG2/qOy0WpqdCkd2cb71HL3BOWTyJqQ4MrszWcg9
kngL4xxeEVCTTYpuB1/duNHZuitID2UJhWnfr2lyEeFwOb+Svhc1Yl4E4Hf2
QcnA2AgUt6rxgZlgEQnHHJcguUkcbm5EaKM/0q0JXof1+C2bAN+UuNv63dzh
cqdhzK+Ch5aoWDnKJ8HHVYiY4T/okSKitj3souuem9fCsc3d9ILt/LBkcG5e
Se5e5/p9NkcV6wlhS1dSieF7YT93VS6JUutqaCLneMViqJ0vqJc1IONDl30Z
gFJXh+Oh8dBvSP58ztqeC3Pas9WHy5IPZp5w2TqJ74O/9lfJmj63LzhwwTHm
XV2BflSBlCT2U8Ecf5P+EVsSex1r7MfRFZWqlrz+gTouLQxgt7xbH/vKKVxD
+PnjrSV7VWfs/L70z2ALQ4CNEh+kPLR6ezazHT03Tuw6eKIXoxkFIUqEAjFo
MscSCQ7gotx088BDcFAOIG45rbeLBXKiaqZiolD61lax39iyEYun3gWNNAEQ
UshupcZTzAuA+eQToM+rz3Wt/MgfQZpdt3rYInq6t3mbXuHydxszvgs62N0Z
KKB3Og1Z3/1VQkBbVa1RzdcYQq292xU5AkQDaKBeoh5pFQuLlDLr5kMJj2rQ
oDUIFS5IuDieXJqDCY01aCbvV20JQjXqkYR5IsEnA6BjfZjxfsUXt1yYCrZJ
0AW+n/L0asefA9WWO/1Tsf1riQpYaAxtBVVvKelPeiD9BbDfH4IjbfgKYxO3
HfkBKpVHceFf9OnnRRhFeKZOcrd3fYuBMVW2y9YGldhLYl4q9PG9bxFvJaOi
xUF0hcZOWuAOdX1zylBJa6LAJgIkklvinwoYFH4vrufy62LMBcmf82XEnM9p
Yh9H8QI1sHjQ3M37Rn8uGZUHJ3rhXa5EnV6pyiX8PR7vrtOgy8WQCxMaGAUC
Nfr6BZOTTmbdIGOgfryCfTY3ykAUephcbOg8Zo593Rj/nMinT8RuaOEvPUWX
tI6o2MnzpLaZJhp+snPz4F5eUIXwndv/3Nozj8c8qdIIUtptRszPNp+gSAF9
VV2j7us9CnOu/XrnMA8crKdmB/5e12VGBn7VTGJN60NsrQrBKrd4oEzYABMG
eO2ET8Dz2I8I9FKNub8NHpO9L52H37UxQoTZjN9u0ARIQBxA/SyanSiF9uQj
kYsdcRLqlAjfo/16GjCUyarHynOYCshtQErS6L4aVqe0WFkcN6NxJieisArh
MaZ9IjZKb9WQ6BlvuRBUJJ8rmL4/iEhRliS5HFnZV/dH+nYrlV3TLoWeZSR6
bUZ6btVRU02WSTy5i9iI0ynahq9V53kiN3A08uVVNpSYRBleF2w/oq31bnFN
v90BvMr0bn/Ppm7oLcZQ34tW5JbEmFjmocME1zBNsNz06SL2x4JoyNHA7Y3e
eVZKpsIhIVSsG2Rh+IYqDzP1bMjx06dul5zkAONOe23yFXpaNije72PWEYSI
0Pe1PHcYS7aFCnT7GSCzJKM6aqBbX82ZGUZAdH6h46qNyE0XV7X/DsDLR8L7
PAO84Wz/cKB7bh/QwdBWUrITUmIZmRDQAmjpRBZrXsQ/PiXkn+0sLHXZiUb3
Xo3L2o2BVyIiyzZ3IEr5Mvqni8ll/PNzm3TT4Uk7v73sM5gMmYC0PG2LT/8J
+SdK1Uvuoz/eOGD++qQ9ElmoGGH6HAvz6ONFQZLNkMBBIt9blcBx7y8PuvqJ
fMFBe7jnYe40QonRepDKeooO/jxoj6pF2iaFhzNJSY1Wvlf3fzZ8/1SO1PJl
fKu9gLnLxFT+ZIhEUnlu7CD8j4npJqPq248DFCr8ylQZWhV1wnZ0DD+zXLfw
T5HS5w9wBTAhRSDOHyvoXhAk5XUa9MgNJ3h4BPqzauA5M7qcPWLICx6/iXWs
iKkdNlpnHFK5RtADZV3VRAFtkNUIfmWIoyI+ZUVgaL+wGsLDJ7s4LJpSCe1l
KGk++EH3HZ7b5U49GHA5w1xbmE9gJlSVyIwVy+T/7VjnugHhY8K3mhY7DNXf
4jTmhEt39iD70frWpJDJ6CL84fgYhJ7mT9HtdODfjXdzenoh/9l0urT0duxl
sIHGRkJPyHY9a/bHvxi1E3NEfylUNdKvqAo49T3uUiLlk2IRRTWb74aMKBGj
k1QUS96feOs+XYxSa26WuRtxMyxYTlazwEfSu3MufYc8HCXzVfTPLf0mAnPM
BrhBImNwE6hZE2FzXVBLCI+iig2+TXrqaEbJQLkFroNxP6+iU+lpKU/J626o
teylq8YNBfQqTH6c58fARggXipdvyfSsOXGyImi+sPqELkph5lBReOEw7wxz
XSaCFEGreYWVlAfrurtuKhg8KkLdTNttQ6+/FnzMWgyuHTsB/vhDiaEN2TOa
2ciaIfOAptreNzaYvgWN1jc6ZiDJg3LR2YR45nH+yNXz7b5RUWmbp/dj1tYh
kV9+h4TChb8KFAXm5HOtnEmk2hjt60osdoDm3uSevunn0grLLuK6LC2Ex1HI
xT9RpeGEetJLmAyYsEGjEnjtkKllBfLhOGsREjsHJBsImMdPRp/WJY1heUqT
pov+6UPFLWcfRgHpUrSasEKbtjslJ8n9XSJ0FWLTaeVBZDpH5qWT+pRRLkMV
8mfUaTj/3Z/p134OGFUwc4gTycJ5l3VC3ItxCO1It4qpAzhrsb93RMQNvM9a
jx3a2+Z9iELuUZrPXK1CzZX/ibuDrkYODF/2tXvH2aJpi6JTguW2MqoMxMdW
CDAYjRchSV7OZ0tCQiszV6d8YTmroHp8MPFceImZfW2l8b8k6A4FfB9CnG3c
uz7Mk8UD1PMH3ZErhq6nE5KYXgz8OJHnH1sDlh2SpvmnFILTciWqsac2KvZn
orsfQD+ENGKMhayqkg4eU0L8LSSkqKjhWqM8sbgDPcNGlHvzx12WJMC5owVE
wf9E0/TCZRsUs0N2ZETyLnyxyCbUbyvsumagfQ6ORlgsdJSHMDumomA3+HdO
wiHgGJ941USZbnl1TIuzFQXjmJcWe0J0GUmpPIOofxrAtvwvJfWxY+uLOWfy
ECs2EIetzMhd/VgSU/ZZCgcGpYvv5BkQ0J3dTvkqWv5m3749K+xkbo4QKknX
Srr3vbyeJiiODecczSj1I0+K52HtnGPLDVHY0N8GsSZ7hLZGmnlNXZdMweV3
DEsogn84rP0ho9Y0OPIV8tVZZaIpxNDGWyW0Fr/d2VaLnOkLbo66E0FGHKfk
mdWINS4elqom8f2VHfBCUeuJjHT6SkdoYWNpcDnLml91dZ/5KbJUYOage9im
uakydkEx4FlJhln4gS8EDZWMM/r9utK2SFos90fMvaCfs+yfn9EsXTkGqt2L
6zWCoU274z7e4YmxH7Jl/UXeq6N21SXmJRuqSRLV+nOQIwiew5F/FpFnBfa4
Klu+abgtrRaM/YeAu0OYWAzxwvQZTF1CT/0LOfUEtXAjxxpiuj0N55/BMVXY
wgjj5BHvKm6GoiqlwdtrdZ01EGhOfn/+SOwpU4gDsvCyVAsg2sTxwk3x9u+q
lKMUZBIobd8NlvXo3QHSZ6KN/xaLhCSZUmXUQdXsCGBo5W4W20cGJ9GkejjN
tsd90lcFpMCHZOT9YVVRVPkS+S/h14Vi2jlny+75X3RTH5jXEu3eQHVmqfCj
at+OucC18J4DkGVoq6/WuKdoorQ1ngmcji+QO/vVftuS3Y495tSTAr1gzIvz
SGZY2e6U+7bpULzESsuTfXYxd4niMY7uGemD9/yXIC+CzcBVLwo/Bki1pezN
PzdXpipO0pTY3xikln+yr7+qEEFSbM2Jt6KdSNkvOVH8i+YGDJv4UZ11NWOJ
BqzManvm8jV2umrtPa46A+VpqlV6NMZwXVVoBwyvoVTgBn234BNTVkXeV2d6
VGBbgzg5tGwpPUoPi0qHJrU0XFIfFSEGX1KgURxhH5AwpMDl12BX9UZa6CxD
HbwUiw3tLW5Tz8E+8CG8bYVa2DTio001suZCKh8jPjWmUdZG8xmTukx5RZO+
FltjckX0nDeaCpXxauRbup5zJMpqv2Xtqqur0sDaUHbmsZ9k7xUG7OYD8btD
Ep8FuKilY3T2y3oAXMWUOFbl2vBaknIdVwxGLYP9RutQKhdWMGEZ8h7lx333
W1CoTMhQeXW1Q3m8T9uHJex0SwFr+ig07KAaBwrrKQL2zBHRTMb/BDdbhDqK
FZtxoDxtvxgJ77wLfp0ClttiA627EfpACeouynxjPtaK2px4RzMjYKrrmw6b
qrPm/yxVW4cty362Hra4SSftcSzIvh4QeOYkPDpHFq6qIbSoU0XTNAEixkM+
Zvp/Nady9hCdQ/E+ccTGiRJJaKkIhDYtIg730ZJr/EULmCAlqkBDL0zBLaa/
4OJdUigCGOV2Yqa6X7/0kfEQTX0wYFrmDe6BJXzT4LpKh4Pz70elVCS498e1
edqLGLjdUYBJ6A0acbmy9PU/dMuqpNsM5NTzDTGtIs/+pkInTKzwnvtkC3xr
GeC0VnEthZlBJqvIY/os95YtQUMhJuTenA1IapZEY36fBySxU0jVeNvtSmPC
y4t+VM0p+z0ZlGRP41bD4+IGwZA5Vbhnp6DN2MvaFgrmLgdh3uRRdJ/WTO2E
BlHVl6qjfP75ogxrU1AFpmNVCVZmg5S5nnR78a1OcKV7FuEqC0jksjoVoH5d
TDZQuIU/mcD/0IwXIeCw4WOFH9QsNMEgt+UHxyr1RfXD9THGf7mPJ9rT1173
gz+h0bzqLQ49MBD/AZRkQ5An74SATkYC6brTjzyXZJaZ5DFimim1CNUJABxM
ZhVbQrGiti0xiqyr1Zh8J2JDi4JVZchAobs5VkWoJ4Kkp+qCoM1pBlU6rPTU
luz5ABnoa4M4woyHzqoa4whuQork1R+GFRmHKIp6eyfoV7rSCwPRtFlN2JCQ
CD+/iUihQL6LUl9Bp6j/PID1AE25PfhDRflzwoBN2TZyZlJm7aw/0ddHFpJU
xjkwUWtw9nhYWuIkeeD/YetTMEAZbc4f44/64w52ZdnDw7ZWvJ/NJpgODY0a
vxYWwocNf/HF3ppf8fIX7s2ylzIzTZ06THT8Sd8u9Sn8Ns2wCR4tZHmf0WZX
/tF9GS9p6WSUchH84fuDKCPr8xc23S7sie4mlflZv9Txi1VOz1qvfFZVqjD6
g8lMZawsQAtd1rS4T4wUSP3Lw1LaYqWab1fDAzqbZInR4FFUsVv2AxUW3eYc
xMlpY8wxInHX+A7vcSPVCdnhM0IXYvAHd8OHrK3mkBm6+8bNlXXkUKO7C0Sd
iQs16a9fipSj+Alc2rbVAV9PmcOBzb9vd6xijPj6J8mG18BalgvdN0I99PBU
vlLt3FuGUgv/ktYbTEAkTXz5lvK+lSAjuB6Ke2f9TpDoxKn0bZ8QOpm1f4+q
WecJlzTjjBSOS+8KYWHDtIwoQ19MqjYZ/W0aLstR6lI8P7TI5KKdFae8OOq8
syA4qtuxdq/RLgBOxdkdQ2+5ACxfGfdi6ftA920oVAoWyTr/3layHYljU84t
F5jYWPAhwcrvG96Dl5222Vxu+2+9frHIIg7tJyJJG0XC2kTvFHFiP6z+Rs9E
V+QsV39Nite8FWg1BwbpGrmmSieyUV7OPoYLmP5B0gB3cDJspy5XMMUoU+41
VnNM3sHhGAjg5gParDdmOz4N3BLfhB+TakDAL+74YYumkBEEUJ9FOq9yFpPv
BZnlkIrnU1i1W6ZAYKZi1pp73K8WuOSGE7JbVsHipfeXGeFUww43luy4X6yS
wLztdhEC3TKVZWZ9IF8wUfDGfx+Jf/Km8S/wto0HUw/wmhA/yvXXDysmPGOP
y1ETNweD0oR8LwZSF0aduvMDAxxZYbzbwaXE95vJxky15zIShsndX2UIMMBX
NYdZaLHWRe6zSm/7za+vxJBjUHSmZ0cayfigR6aRHjYXFKSR9aBs3EhnVq5s
drKeCn+ccYea52snf7+Rc9BVGcwtjSB4h6PgZKHZY5ib3Vo+gDCttAlLHDLO
bu2h2vDrydqEuXsbzqG6CFIJfbWmqX0//AiGmU8cHIWdfxX2plsMyR4fRW7L
AdXyKUWxRaMTJL2J32h8y9XzDyW6lKmZH0EyaQinZd9vxUvgHp0NPMUlUCWt
Nd6SvSuG+KOkbIGpQxkWMP1Ulmbu3F/X/ehig3NDGkiD+5BXQ0JsyOG9NRdS
dP+1ljRtrDrMLHq4fmi/cP12v41Ms4EXpHREBoYmLMlidG/7BNrYemoen3cc
5C5e5VbztuMc8WrZRJfYMhPmoEZZwfytTfONP+Vn0CFW0ELt9adT/IjtUNC5
7/KvplNlJSaJMDPRbu9/FifL19icD0R6LhQIezGNyPcFKbyhygvZw5htbfy8
jHEsdRcpaq0XMqFB4zJC0sx4s/UK2/FjBz0mdzKa7g8/WFdW0gl4dMyL4mE+
X4ih1rtxcQ6A1BicIYdu5tvcWw69dhMO/Kjuqt5h+tBkZ6TKAaHMt2e82tVN
H9pv/18GBO937l191i1Bf7S8wFEFZ6cMAZ+YlUuZ07ffKeY0IjMtNG/plIea
akyunO+Ij0H55Vl5+TVnhJMcbojTIOBv0okPE/KCvnFUOGkF0cskgnK53XAX
Sx6WyUlQLgWCr14baKCNPxnB4YNJSUm2T0f0t5x8sRCz7dL1Lrj1S3y6BeH5
+FoPmKtt3udozy/NwAPuNOgAURhyWZ9TFTTRUeRsJ7noGrbeCu3yGPzadUKX
yRc5diIMOAVt4+vBE9deB0qkk5WipjgCuj83GyMTDFGMCc2ljhG05sV9+CSh
CJQf5CM8S2aKHkk8z+lPsthFx3Txdm2/iJR9b6ZaR02NexD+os5BUjc/TvlI
VKH7zTevyjfD2GBWiRponm7Vi3LSk2zw60l+NL03BturyQtZXNQN62gjuDh9
RC/4gPXeqEsZx04cpxysO3enddwSmYdZH2XsHB2BCD/K65sXGWDuyWCTeZaI
LXJSPZMEfXQTawzUFwsyIcQtLbPjl55fhJ54CIyjjZLkCp/C2F6gVLLDPPti
s0lImj3JRASS8TPadm8TdCBzyCMj5bpXXkScTSfn+i3bKNSN1GRgPdpprEKE
1WfPxYGtOKFLnLZ5LpsMPxPaGJmpSdYDULzcM1RmUetOC1BKdXFj+/Xmwf3t
hF/CfJTXw2yf9fg7JccPulW9IjLpkYrTH6oM1LflIK9TAUrogX3wyaF5DkX6
1EchnoU4P4MVMTxhIKWvZqdPoDk/OzGEjCMvOohVmTwkWrr6/ClV2rai1ZtX
1riYhrP9DUhEx708TcrzatNV106IxaPRn1+0v+Nq2bCkvcrZDtsEC6TdKYuQ
gzLwLKu8vATpyq3cH/M5wbUEEEZgMJb/myq2+xSEY90gyXqjafegvJrKWeWz
9HPKynZ31oSUIeUh9UY79ZCdgL4d6YZtPXtE2QG5RvJ5Dv4a338B00Q6ZIGj
TqIHiHGMkjYHIzG2IWwcDWb4HS4qxzOcoy6UXaYdr1/2mVPUPrsAd6X45QJH
MnuN+Zab6t7+H43fLNxHkRizf9KiFFT9eB13jnvHlaDBLEUdprBp7pvdtKvY
+5Rj9yY88w4qVE3TqvnkV7J6Xh9qtrc4tMK38baYmclMuKqed8L8xalJorKb
+jtlIcD4IEFsbZfBoOiEYa89rmfyAOLee3+hLMl6UTOwwHKfuf8ydW3f5V4O
qsiInaWJZBIRhfToQYd2JdCC61LGr2C0fuIf+j5qymT/4a8FsMMbZ2eZhuQR
VH3cdTOYrXiOKJCTT4GmpSk8FBivNQ7q5HNMGukAvr/s6O41SuGwNFftWxJb
HJI/kSNhkYy5DLWTTdfWsNa58Z+P6GfosT1+lNxw8RAjmdaGj+MKveCvmk+g
uFSWR7kUXBTPw1wqQ6roHH7pVBZ13SgOmcutqVMbczb07qn9Yy8ij/mbQUBV
QLx2B9BF8sc5U3W44c3AkEzWNkMQQedzw4cG6msnTR1ECFEQZad3YczIvknA
N+VaRTHR6pnqL7rcjYipB9nx4VX3pDnG1lVfs3RwO4pSG6zBak9cFwpzOq0O
BwNgQ1zqlzhQGMnu51uAqNXN6kpdUK1fCo7ofsQ2ZiQvPZswwQuf9rCdhDAU
/J/S2epxIHdnbnBXCc9ajN8Seg+nHd+qX3PDZR1Hk8z1ZKXoXstNSCHK03Lu
sIeYvc1qQBz6pJoBsYwm82h9tprKQHYpm0/6SR7cf63H0l50v6k+lvgmDsdd
6lEMcFmmQWJNSPh3XJzL82RbyXfN3MGE4foNQP/6U9RBBW6/hv8DRLZnEZs2
OQB3QXCi+goRCyCiTfnHBTMYkPUJKx+hRxFqZvFlRroHuVCwAf3XKTI3Fs03
I4/WXkRDOs04eleCdSxCGxFthrz9k9hS1vB2ojZTdk2OYIy9RQuLeFKl699O
VAat7TybVgJyRK8u4Sor/o1CPZlUG8yQap1bsv7x3lA0lUVG/Kr5h4KUim1x
+hcewwXNEMjxyeF031IYMPImFlWclyxfJPoazxukcZWo2jMK3Yabkcec+eba
16T+zMxz62qBAfeE/j5UnBVCm7yryNcDLW+L791g5pRBcZSnkHgZnpbVEDoc
mJ4PE0/axQMMK7YZvYTsPpovb94VpCnzdnjFTvxdyWH1LdLVqhIWJeqKYjIe
hwWZrxDMcCjKEN9tZmatWe11RxKIL7EeCP8AicjMgCHsmN60yIQQbiQGAG9x
D2E2sDQ5TIva+Kgs01NDpxzAfLEkfu0QfgeB+kYXNFIeL1KPC9hPHckrEtOZ
ixuYepmq2GohMXmo1Gaqh19HnBxFYu11hZj6u15JABM4e17VMldU1p0csVFL
N1O0ewCN0Rtxt8gAKegnnL2pT/B8e207/wZILg0D/7G2VnvFw2uAWIEIBfMJ
LjTo5HlA4VfDgApam2l4TG5FpbxruLaiSE0SEWfqdttPjtjORwvtrLHm/bnh
7Nw2rjaboJ95ziaPldXMuS4KAlR4EwzH6cjt8ELAC0vEkKrKXE49tux8+sdE
X0QXZj9z9Ir2Il/0Alg7HmOnUJc9U91Fz69uoWfT0kcQXvshaDmwDnai3HuJ
oeymKNgaDYwREo+yihQ9ZquufiGJs6+PsUlYPBBK3XGtXJge/IZWThQWC/uM
4hn7kI4XpX/h1nn3G9VEfPsg7xodl9Cbw64zJ/eDBjzQGRUu9d2724k4ejip
AtzvuhjldvndTqN5MG4GTEyfz3VikqMWqj3wAc6wsVYHC6q04ZCm/etWcB+n
1DVL/HpN9ZYb5r5zFfddVn8/bDvCM/33R49/1IPGle6LKJdd5Yok4V9pjn/V
MMa8Bhmuo+pPhq+OWS5zxCn3YubRgAGLNpvQOJ8oYw0w7gxFAbiHzRdcPAbr
zZvntoFp7URdtXRZvR5YgpL8+Utdgzmus8HhWz2h+RW95iui+hEXVcmoHPBS
JCQRdk4iu/UX3RiZhWEQJ06J7RTdw+G7oVWh2eX6tn8mEWLOe5CtewHoBIBG
rhsw5D1zwLo+TJ52Vm7aLY7wmo15dI0+CRN5unlqgozK/YKbnRnH8+Gpgd5V
0eoQ+LHhvocjCdvmtFN+6bUhx0Hq+XyZEB3dSGa6rwa7qC4J23VJMMDXJOIF
+NI3piQ6sJZ0eAbYrIXCuf3EO1+KUkuurkYQxA72mRYXSPwekLr37OF1Zigx
aZwHav3O+ilpGHowciCxyHlgPh/fGbq0KEMSQMUtZTZE1p1a6Nlx57S8Mzz8
s+3uunOvFd6vtJ3ft2IKbqARnjNJq9ujl/jvfG6H0VMffT8cdqVvfTCsuaP4
o8LskRrelHuoDt2pKsGH9vOZaUZDmeOyQ6O784bQoh54jm9+UXWlGMubqygR
WL5QoC6o6vFngzCEQSXQ0F13iSzJ02M5T8kGBRoco7OgszSOxcvknivMzjVF
u195rK9WUFokxRQS/76sie8ZdHm4ld9fyuFBdDw8iH+5x/1C32PdNMJxIR4v
CrXsfgp3GcaTWs8rgNze40/F5rNKaaaZLlfMvh73NLIkOcjQyQBfyZgr7Dlx
wmYrJXgL0UxMmWPmMLA4tax7TfBtoOwW71prNMe24/lHCg93//TVRi2f+6jw
rNoJawzoZ7/eGPlGAIQ+NpL/HIL9FPOwMTVrf66KX1Z/mw7F5+ZcIwRgeZQK
P5kdh+/3P8agtmqizGvbI4COpgldc1j0J+pPDcLsh6uhSLvizukTMwSRc9yz
xC/roiyKS4obqvobLzaItHWZZKvVBsNLAoiR8xRa/eLPsRYNTcp39qyTgXYZ
WEZeqbhoBwA9s3b0mWST8SFlaOzcVWmPxQ+YDgNiNwwOgC7tIqSDEl37bTfE
UuEdSYnw4UoIm8WlNBqR02YdJGrw9XVJnnz+JeL8hpqorU5627GbhEL/QCDb
pHCZJ6Cgn00wh3yFYJhYRspiaf/y23PN7Yt5TtUQkTntknEbUb9PqYdRa2sm
UPATXTyQo+r+fOxJ69j23qHd6h+qTNAWv9wtcPp2tSi36lKy2SisPDkV/1yZ
NFDNYMAYD5wMmczE3Fcg5ofwWIEGLZNR3t/FVaqZD9yBOtUW7+mLImu0Tjo/
G9OQt5kA8+/5iUaogy1Kucu1NfIesoXknOL4TUO0MZAzayxYZO+VXgSkfQwL
JUkc8nnS4V63Ifr7yb4bHJG5NjO7CNNE9g3nd6dtPBfLcswdjIYz2VWn5MSZ
GohKaZ4cWW1jNLRMTGkvwhwSlK6W4MWqObN1Bit76yE57EgujuyA5PulMy/N
1NvT6Cn+C7aotwHSv48iNzGA8y5jEncl6hPMMTqi13WLDrHzTfb5mVi3EOGc
b62UuBIN8WEFtcQWHZMUEBZVqp251VefG8w/HYgmrT/iNbPQcDiLJIbvTJ3L
Q8IvH1Mwbym4EU0hF/8zqYinFRFRpTr8dwCugZ6TCpWjKkMKWkQEDNj4ShTv
7x0sCAzegZQPBIdVuTkmh/wKPOCHm8BdGZj7yNwCdtGwAVBtRwrmmOEeHDCR
GVz1yuQur75EwPUyZxKVmzgzJ3bvdBbdAsQ2Hl+DmaQinxLEd+pSz8GEtNM/
z3Wn4rPRYQGVlMPJfmYxVJcS/5nHOZDOJaysaW13RLz66LElytGExZyw06Ye
YAMd4YuDhH3V8ghb5aw4FLIPdboPP7vB9YF7Awhtu4OK9tiHwbZgZQ5VS9m7
qfGEUmTqRSGgFUN3thOXyw9gE/aml9MYM2Ds3bXzMU3YmPH/DEFtNTRHqOeI
1YjnU5n9bRObWTqmwu7ymx0Z5ehg4S4KbfsY8yK+OaFsSNR7kSziHg6P8gD9
PGDIqj9hLNexAxxFlNwN9d3NXTng/gX/wYQWui+GJA9AWaBy836/f+8rFjju
BoiCRGFVF92dQGpBvtxXXxRZyl0VzOlf5y9jVf5EwwHSK8y4RzAamXlUgEt3
tUdeJNweKgWUmXoS7zdLZLUtgMNUozTRJdKSQ0qVwWYbQBY2hg9APBlzYzQG
/n5WqSdA+nIltB1VAp2sN0OEQy80xRojNW7ZmKWHAlhW2vaghGC0R7ii3/Yx
D3ZMSOC2xa3/KFCI/Go8ktwWYNTM8+ZjwHVzRIHCAZgIRPEnUH+3hKutrhxC
WhRMz+rvpOZUll4dzJZcKXoabvKKgHmzyu733gTFXBuARAIFW0r3PVsqssqC
UkXa8ptWQACxM75eUy3a7XjtSAeIvBUHu+6eQgMpvNMK97Zj3FjR1JV/mLry
0w3Lyp8TxWLK0mo6ECSuVAqc8ftVDgow/3G/bJsg6fPw2ax+Ki0JhD3+gE3h
DpVMjcJD4aT9LIZW8L07kpkJKKA1sqhZjmMxHOEr5UeWt1sfm7PGYYy5RP2A
Kux6IHOaU2eKL7vUm4HXNUik4ABBpym9SVBjbDIRrzwpGra0vo7y5RpxriZG
JIdzE/oGq+kLwCjwOuwConRiN9mJxtcFXX2KW+gTG5dj7Zw/2Dp6O1wMctkp
tI3wmaeofO6UeLtUVHkswdBxtTxjH+Bl1Gnze2yjVQghZZiR6G1lAghPfrcf
HAgQERdVrfkln0J6iKVlOgXvlUiatVsEY429eMS65DeaMi3BWxXz+BGQ6/pJ
/03HEAz5kXxlrFIrlCzu5WXSNRKB3MMJ8BU2E0YzpCmz1ZTX9ldlIlTA1Udp
rAR07vGM27IcMT2FvkRoqEtJ33lQ5h5m41jERRZb5b9I/W78jg/lwB3Q++3U
dRVuWR10N225hf8RS3apfosxaws3LBQv/mdfXZosBbLOMbLCLqpjo68WquUQ
6AEma2PhFc+VyzlxAVTiAraiEXpd/fPjJog5Y52rpfeJQCJxPyru5WqQMvY2
tX9YhCUEDUaD3RtRqIFUPCp9AWpEGQrugkvkb8tuU/amI067Y3qAww5pHOtp
3Dd4ZhAs5+4l7yjeh4WE5CpHRA3A5cB23D2SCoFXcbdBYQ8AfZcVBEuRYSU1
ss6GNeLI/717AAOlPKOMCNObSr/CU327sThJesByzMpxAOdsDWeqvYsbldFI
45XHj5+EHOlYIwDowXe1naCVf4Ryp/PQyDvvvhdAoO8kehw3KvFrXJ+tkKno
ty6YHBxqcI3b6UmwwVb+VdCAP9s8Vw69XEWAFiAhNHzsLNnxiQ2VN/Tzd66o
zsc0WPittKviodYCIPeHaaRNokGAbJNItmeZX+776HHybY8I4/wgjUcJzDoB
XLpXft1KVY0LOi34ag97ESlq+RD+d0oQXzV0YpGfD800RbL3CJSVCuqMho4E
5amW8b6IEZXQgjtKsuIPhMr7YZrb/Z6P1aY4kn4LXIJvAD9kd/u1p3u4Aot6
Lh6pzHgBlG1lemsQ+NA1ItLHTqwJlG5WQWkwuO2xoFslnnz0VnMCukZddRUy
FlsINmx2BkQbF0oNX2gG4sStLe8AXouj5/rATablTea/c5kx5SUNkjAD8+TU
s0KssSkTo8JCqI/BwWOu44TO4or1h/GHgS6fY3OT7lzm9BvqL7EYcSOwKUMU
xvMjzKWkCz+9Y5OwfMBUSEiIOSKnC1JeVTyHJMBvWnPfXHRAIKBsHnyKPSkB
LMzo3G8PtN/jes2Sw/mX6PJRgW7PIC8+S+wp2BeUp4xWvfi1jTG3dl83r4gf
1b+i76xH5CaXXJS5Gr6gSjM1MCdB8I/xSSfA9Hf6K7wxopgYLJDzaVCrVEZX
nt0kWS6aJctOFk96onY+xyPtjDDfXEKUy7J6rDjvwZiChlkTfuHWDRjZkTxq
YZKw+HakmpBgXu6uE/vg5qcaXgRRv5CmEgHYheae+xsMKgcIRJKVA6Gcu4hw
ILoAWj/xfXWbhcuHj0UG0Q5KaJi+3fu5BypqmpszZkMLUXN5Rg65TUFnjM9J
DEcIJlknaHZgTBjNmwLpsafmH/uQEYaiC34kq5xucQIusE5sZ7oRyf0WhcCW
fgVtR3trjbEJTs+ZzA5GIF2Xh2nraf8AopvMJCUX7+Wzz6C9Tl+BA3vkGsxf
fTLGS5JRO+jWWu/P4F4Za3AsUv2TXozCBYbdAIWwJEK1Khsml5f2PLB2+Qxp
PG9eBo7rmMW6CxjPwAkIo3lqomNanZ5mFIoHsVaDWVg1VEkWlkEzwD2m+fW0
p6eI3/UALE+UHFnas2jcD2/zUcOUTgN2nHYbh9/9Eo8Kk/uSV7oc2Z4pK4GP
clEFCBfSpEQunQZJepAgZcXXfl13jz1Au3ms5HgidOgcGTGKWqEFDAbw4vw3
4wZ5wrQmMfOVNROvgnfGE6P8ihTEHBFq6TzIjbT+DYTQSfhXj3EqXCapn3S1
9ZwdudogSvIgUTWGFO67i1a54Z1YN6ub10BCD5NIeR8vg43SdGEG+7FTgkkI
xIIwy0RO82TbX5z4uXM2IexySDxxG27YJ5DucLa2wb72WcU360aWcGU0dY7s
iejjVeeAteLinKhZwrbY9ZFN9IbLKKSvkIK7+rEtr/c05hYEoa3gWR5OWFkl
2WUTwF1ekxbKHzREUVdxO65FQmPm3YWZvc7B9tNetKLvLsKDsTAZNhUIvcrG
xGrAk4EUzIlvefuoyzNrJj6adEz3+DeRoRWnPtrr0o0eLreE8J3gbplK2i+6
vxKER9NHMt1YyopAmHkVgITVGY3DNiYTu9T4wQ9YJAOnYSkG68KUOwG4suiB
OYh0LRsSD7o9mMpz6tRlNrHk6quE5luc5l8HucZhKGNHH6jXNht58EgYTlma
697QqC+5CgV/Gg71EQOgatVihUEJ9qVuAyM0rZi7HbEIkDPfq3ksQ5uueFLO
KrEPO6NYFSnjT726oMdcQl850slOTgYkvZ3c4qbW0MwOKcMEph3tZoXhe/33
XajdgzKSodebesAjJig2rE4obLHqMrSNQV6Ur76msCqqlCQmD9ikHD3Lcdw7
2qlrdiYT816fQ/JUew9Tpmz/EM9UhyPt4ksrA2oBBbRA0mVOFJDx5EO0gPsd
RBqACDisijYvjcrrjyiDi6fAI7m1ObN/aBmZfWUQaEHAKDN05qn2XnjrRPV1
MseCF4F8sVF29YPOx3QNicYX/d3TvL5wQJ8vQ7hW2OW5G1ajt2UReATtaQeM
VkWz/jA9y20r40GTE0vISU1Hnu6gS+m1oc6yUWgPAi29no/Kv+rX5RZlE8Cb
E9eBt2TcJHvdhdFoUx1QRCFpo7PNj2kJA1vjJnntWZh1cNyezMp7XMWghlhD
C2YpOudTS5SgPVP3+jlvpkRdO/6pmBnfFi0AzcEGvgwyQHQ+kWoXUM+R8OTX
hkjTIKTiFT+Bthaf0dqs5WbzGqGgRB+JHjqHqEnLirlPvNHTRYEZQhiV2VHb
8ihgOje+niAPGQf+MyRsFsIlH7D1+ItFBIOfTR7tnQHbh7kzM9fRdmE6yCPf
dcdZfODnuc57qG4j1uOCGYQ/h1ZWgL0mPFIjfla0e1gRXBeBpQCNzfIA4Kcn
IBj9CPlgARV3+A8LR+rFYk7ZeLCBSr+CS8O53Ko2/9X9boQTB2aHLPlnItTj
B6t2j3eEeXR4RXGKhNV8RHk0VQmO45y1bsnq/tbXSlwIiHSlZivn8CY9F99w
mA1HOh+URIZeBbXVM3xfsoJx4RnJPcnnO7FzcgFwkiYtBf5AAGyJEIx/vrFc
DvARp4/eyOUxmLsZ+3TLlqKWE4ezRO7xRdFBCe0pEgw5S54ddnmyZu+dWgzd
S/H7X7T+Et+Y0eeqqS9dn+aV6u5SXmjNrrpgJBhXdfnwr3tafi1M+6FQTlXt
PPFwYk1UhF3/YPCO6gzJiW/iGuLkGs9HbS5cYzq1xXEjc8TavOpnzW/wFMSg
7SsYXtqXhN+L+2jboLIus843nciPeTkF74PP5GA7rK/EQjXFB7gIOxhEGqiz
dn275OmeQX/OfqRsa6S2lc+CSE7emC0zDxGoY8C7P49/QGUp/YIMW2vSOsbG
TnZFrOUtC//JSWaktmXx1TUEN5UwPdzZTuTpNIjAmvfsTY1qb/lSJL/ZBXN1
78VAjFjtdD7pyAs18gzaaSf5pT1vtIbl04wIaH4WiT5y+aUINrI1u7MR++ku
y+EAJu2wFhpiww8n5tgNm3pFMZoJbfSeLpWVWYjHBtkurnHXke1vKZGikJha
PtTHZsCD+fDl6CUJZ/ogfxpyADPcE20Jp7SL8jZJRlqdxoow3GgTnBihnobf
vcoPQCX/jw7AlCwRBmdGfs8WFVdGkP0tY38oqY75Yjj18PHl4jhQRgAELWRB
D9N8ntRJkh2wmCC7joZpRVirB88aIpOYbTckkYIMNbELWbPqaWAmyBLxAyuP
TpBqm1E/Y6PCeaVfAkdNmvDv8nukc36OpIGHyYQheohbnTb/imQtg3b2jfAL
frCx7m93Y4AGOj4joED7ti8kLHzNdne9uOHczGeSRy+RV0HgEctWH2pgQpLd
gXnFmESf9S9qixMXXZfLzVXBz9KkFxYOChS9wKYY18yZPL0TdBK+0RoPgbx/
ypCTM9bba6IQBT4gyLKpbyuBGxWyB0zNnNVHOGxkoeraQCoCee/6GNSgIqIg
aQ1eSWzhnM6Z5jL7S5om7ZVEKb2/jxGbq/WYBL+Bax+6Icy3FheqQfjbPPqJ
h/iBrTvqJS5bBZKymAPJe1aDJjhqaa1UaZrmX1cRJ4apTRLF8kztSoKXrERj
IUIXpJ6gUtqvYS/lH//8yc31ASWhSlNSEr2+swT6vH5mgJAolEeHx5aCFFKu
YjXSbHoaJKIHPJMt73ZV26bjtEEqCjr+vk+gKg0/MB0HOloBMnwiUk8Rg5Cn
bZK4k9jvEAu8LxsGZcsGMj3TCjXDjhccECZfwV9u0lLCppg24zDXaF7zeDXg
5UASYr5Ll4x4b1uSya1o6dP23J+3+tbnOYK4Snmd6Zb8bQaEhAH36P14CxRx
GqeqkrVaOU/Ol9nZMnOQR7RQ5+YhE0qo0f9i+qYbDFYes+mXizxAeR49pt3e
bEqUMsyshKWUEpoyCKAEf9Cl/xzHQgYsZd48lW7F/beWWY0f3EXVJd1V99nb
dX9abkqCgFWdHTEZR/DLr8o6DDBnW0sdiyNyWPTTCoGQmW/EYgR3n/ROPX30
V1Zmx47ET4zWWo1cYpsxrCgO3F6soDX/+GTeNLVJ1o1aMc3+I06m0opuFvOV
skKME4AuPpZO3CHzEPqGHO9inmnNKU9+tEx9Kg9WF78Alb3ZUwq1Afq/tbXR
VwoxNIMmJuAX2IZfVudy1aosmCtCIo7lnD4ud1+F2DwlXqC0LLyIVCNZU1vG
RsFFRE1XCcazRXx61QKZP6skxVJ7v/u56uk6JODj7J21x0VIbq4OLJr64Ys2
TyFAsEyVeCoxUP3j17H1JFRVNFWOsg5Al93YGk/+J/78saUjq7Y6RmFrrTT1
S2aAy122/kBigReWxau+HFs5AaH8ZYYtJfxF0F3OZhGE9Otz8wnsoCziHhUP
vYtLTXdfAEcBfUsyftbFoAe5NdBiVnRbW/679HGxitUkraEYLgv7b1D1nXwp
YoAIZViNpk2FQAfkTNE06j57P/gNGMZjyVgcKMfsNES/x54agHDb5NhBv1ax
HW+CdFWei6Y5kbgcxTFBQ1cGMoEo+1pBNpDTp/xxB4pZUaX+jpFyw+96+jF4
dqWxpP4YUYaHtUAqaortRTqi3uMCJZHpIfbg+3LarG68er76K5PxzE8SDmky
RrtB4o0eVvcg1/Z5oPX/VTSt6meZ8IlD5PjTd0YwiyZ1ZolICCo8PXdX+kaI
4SqtStf/FwoIYIPHhw3TDCYxE0bqqPgo2PM3yptfWLl4MOgc/jGPRRmqO70C
ecerXILhwL5bf6wHQUI4JPAtg8S6leFWiP8u0qwHZNksVuA7QXOBiYN6nhsM
c7BVOTu6fRKk6UcA5BOHuj8n5AEdFATunTSR7GrwlyXd2FtCkcx0f8IMTVe5
xGy9798TswmvPGp3lhFfwfalERl1m5cge3HVGvJ/NZjuUeVCn7rAUc3hFJEU
V+rKtkkPMcwlpfk6mHJezx+YIqj6WIAmJnOGrePwVCJSTotQ3Ei0m97H6WUW
08R+zAsM+lIrIaRFIVBdjVIQ39JAsy4tdyktlVlX9DX7a1pubNNEP2I0VGn7
oZAjRvsAh+RGE4FPNJ3YkYmEXbBzP6MxnxswaQfIGNFDetHiCSR6H+lLssgE
2jH3tPPhdbI8MLkwwm4OuEq7U2i0Csduecx2nDQpGaxLf/vDlsR7uJYEZNV4
0eyVqba1Z4Lwkxu4WnGRe3c2ag5QWmhVSQLrkzdAfKoTYTL42GPiADj42/ms
amU2novptZmQ4AG3CU3Myo+fT7rYpaSfSopZADqBhFYhxeC1EHOnJQs8Y5ht
qEBxK8itQYmxHXi/XeKJ1cZqn+Le1FREsFd2a7WbPwlx+q+mTC4c0NGrtyrT
keto6proqO48hyoA4nbQ8U2Ag3jvE8R2Xpp5Yz0rG+aMlNUDAI+yoJ8CRe0Z
KZIjC87lzBgoGGrXnlJ6/qoEL/VqCvqIBdO4+/ljIP2NXHTfUwj0QI7s9wn7
gsgVWXf0wM9Hs02Q8r9NOeuKTa1Q4Z7D7zCmAAwD7hdVf1uTr1OUc05IS/Tc
FE2v+wsOeRadX+kAit0ca7hMWv3O55cP+Jj4R1YJ/ohhC9rjcLD4XhV1ouQR
YvHxp1Bsox6q7SuoEEqxseWX2L16W5xvOph6dLg1hnU8N8gCIbf3A6wsmZp4
zi8a4jwpIqJB4micWWO6puYIWmd09+TXSQiIVgbsRrTyo095oX4m767XXOPQ
IUigZPqYlUvWdWB3pFTOctEkwBdjFQ7v+o4iJPLeD5PamhYKBto6Oi/HJgYB
Mx3BGNF7OmisgZcPONlygvmFOnRB9SfSSml24YnsAuyhmBGrMyZbfRY4+la0
976UEWFLajLqZhAEiOQiQil9bjiSXO6B8A9fJ1vXO7OkDHPRcZ/rdEn7G1rh
XsJPi0EOistBh0YVb/TjGkuCw+LySXuvUW0AwecWZrjTfSv5Sb6McCSBEy1+
Wq+iN92vEXROHV96GTi4cZO5oyyrM72F3pV1M4uSUqLcd6aSOcNbmfKhhZCX
6y00CXnwvaFHcytG5KQFK9z97HIgDB1SLe1FkodSTy7JQhL2eYAuRdk1Cg3s
XKC3ZEWbH95S7urabGkkPlZ7O31lupX9WpipA5CBzfnIvenTc29U1yO8Qkka
82xmzgYw4R2H32w9YskJx8CPqGFfKf1mb/iOSSetQ/98t69c+3Oq+LH7lPgi
mkihDjnCiN250idU1qE3PkBzBWEaCRPMrjPEhUlm2yBVMa4WFfmRjkx5ts8t
kantrPtYBYzUTMaFRoTKtPlK9ety0Up36w5xXoa649RJBDYwDm3vqLw0rAlV
6TkiO4NSUO6wNlDEUTPnUxsXGqmZLb1c7nvy39jke5oskgie5HsCJnwbdhbt
nbe5TEbFDs1GMVshy9IlrJbWAusTVQDuI6FW1/+P2zMQVRTod6lKLPnUnku/
zx1SbPmCutddzueYVHR06JeCjsXWD8JZessB/9vOul5/9CEliHY/vntS8kla
YqCric2OR3W7D52/hRXQcjWFjyXP+RTqXAkq9ussvYVNmZNeSIlZCRUcKGvc
3Yg/HM5c4DTtlzmaHOHPMpcY/WEl8aCDa8WkKl+Fw0C0ndTdECEFVpGPCCOX
+vbNTaID4xKMo/6zvcuwzjOiPs55MiUXtLBzE+BdTcXMRZat+tyq1l6I+fb0
V0epXruZgE3X3wP75RxTyXvASDPdAgDEMRJY1QF2TxTbTRaWfpIZcFLwIcho
nGAuX9g5eNj7iDXdvuHC40FRuprAorMyghYB79yeyVYym6KvLc6FcQpM09ml
NXJopyXzZlvkS4ZM/KGlVxhPJkRTwTjaTeaa9jn63ZsvU9VkT8FGeOSUJWDY
3Zpr0ATE4/N5Hw53OgQj9pSRUPM0VAfYzIkIkuqFsBoY+KLvwU+VmHkAQl3S
z58kO5xyoPmrozAh0Z2Tdor82b5l5g0R7ctLpyPdehRUA5XjyzJx0SbAX9aX
HIPHRVof8cknakqOCfe9QgfvMxwOz468BPaiGBQOBgMyMxtgcM5Z8+2588bO
uNFqDvGlOECiI+D3IXxSkiTYT1i7/vJQpJNXF2jBWU1Lqc5TxWuODTYR32CD
F3u81BTBwqDW5iuKhuPmn5s11039vTgX7gXB8Cl22UB0yk3uT4259Hdy/s2s
IsOoNNi2LkOxXBuBC7VE+f8HKGz0dd8rcS5dcRbgVd6PgnNusffBF+AndPlQ
qh/si3nhR6GEmy5uIEztIB6oBCVG9fRiCgeUU6s5RksffvvoIrcQSjChdv9N
cEPx4JU4MDhWZ4eh0mTdi/nSX5pXiTkfSMPHGNHMgjXsm/6CU4weAhvAjLWT
50BPJwFhTlMAtoaXVMmcegXS1ulGxUR4ZjBUubiS+O5G2xVdrBquxwfrmWLo
ol4AUXO+rpijx3y2x44ksAuyB7Xl14ektvfRB5KraMbaL17ro1KPT7KmOQcp
IbKTv4L3ABug8D/xwW4hFKeFsnGTlYNrcRF7vdnBuTiF4GXVO/fbmiR9snpQ
993K4nWqLYV4Xc9Jfc6VUKwIMKu7/C4u9Ap9lg4wuMox77OBqn8XdCpr09L+
tK6rnh26mfINC72f2XC9rlhZ6JJKzQ89wFe/Z1EgyuJhDp2ERFXuaXxoDTJW
YrhV23NbB6tP03N1in53GmZ1DaO14YcGZcrQGTLLcK4w7Diz711RQN74ViQM
W7MoHgBbLbqiYBScCAYlBiVosGY1t6nN5oQQp9tE+4L4Cv4iWF4sk/+F2eDH
PvtdFLjQ2uIj7YSugq0XXaXYN0KTzAFduxSqduyCGFmQi4QuaPDnHkMpozId
Wf1GBbH9nQG+ziRqdUYtth4LfUVf5ZfVogZHcKhvd8ybgtAKmxvKsANNne5m
0PLIyHeOO6zhk8NQFQzIF8v9t9yY7CwKeFCEceUrcFw4pZ/9T1jK6yunVk4s
3yAcg0SQ2bI+ZUuaiayscEXnabCqZM2xfEnSubNFJaR12A/s8bA8/J8L09A3
u1HlR8IpYu0Jvu1C/XowHOcWMxizlKq9SKmRQpvTzrbDSQkfS6Zmalf0VF2Q
LWdUGvdhQnyUMa97YTtO+s9U5z8hqEdwcMkhsqpuNoI9+wzvi/pMFLbKxapD
rAsKUSMipIye+T03qXJ6OZkdyUIjyGCtNHtIIkixQwYGYZuajaLciU/vfAmb
S5BkH4tIPpzEXKMS6FSzOxOcoq8FrCyLMvadEMuSGjqFM12jW5PBJWVa58L5
XjTa1dSfMRVNepFpxYjk34tKydZHqRjjgUUUm8mt0Q/cJvPi82cVdxTdwpbW
6839laYMuOx8pvs/mbVbl+RYKScvsmf4WS9ZH5lnZbYez6EXtJcGhxb6Lf9U
X+lfLR3dQ2jsmgglKHCpupRMIVUTK0x2iacxrYt8oSDneAvZBB5J4bJ6EWe/
uKX230bUQa3e5sp8kwEaL2dQR9UNqHFHeb6E6eqWzHIPVU1IF937uZIZlL+p
m7cjIlwa4C25uq+fsrfJnDmk7bKnWJN+0NIQsgkzPhmZXEyPOfZ9wmfc3iFm
KFjNZzvkhgEUeEqFEfHBjszAUTjOXo8t97ZT7055Wv9pOflmyJXyXgXGNt1M
FkXCyODZdxVODK47tDflL1uLDKgHCdFuvD1VO1byGUrBgSQwye3+8gkXuA6I
rqB8f2S8L2lLpAhOKWs3mR0q2ZVDpRs7bLhPfR1A2cU5s1gBTmSbbS4AelAc
rU3rTdXKJHlr7pTxdtqUt5jR5Ybyx+dhBkXgOzEnW8D7QmrHe0CDV2W8I96d
cMePe55E84/uriqfVuY4pDRXS+lwQ7keABcE3ka3VcZCAsAsrkxv9Wdqfj/D
b7Amc11kV+36q3d0JO8DgpH0onYzQ7hZAiIh/y9RoqT748lUtZSHmfTCmBzB
PPBThNTinxpbg7yunA7DwmfD/ktwlPcMnz3p5bC6Tyg88kfBegOx7dRecUFj
8Bmy0fDvc7Mlmla56mExeGx9sziHKsK0MLF1ODa3Vk9JhJNES+U8n0qkb+Gk
D7S7drxq48s4+L2m27BK/x8VZQhZH3Uzc6TwpeBVlD1PopGeLRXw73gJ3RBW
l4TsHLEwRJOd8HkcZYzAWQPv4x+5/yUnIVGOQ8VcSJuPtLF8K05mm5AH5S7U
gE+XFvNjKDMqCr6HIdPOrcP/IC3BdSwKQyn+UkYutTYb9/T77QYb/cELMMer
326Mnyn/0VHpWLp2AbARRZuX+1zcD76jsm9aFBOcCDQoQvLRvxNrOgwsCWQE
XBA1z+EeaQ1N1ThZNMFlLFvcIXAkMKXFs8fkbg8zyZgyy/4PGAhZcY4RJ5yf
usedvBjll5ewDdth2RSCkZOnKhEUs3RdVxup+mU052H5dyJwi8fK39zorBDW
euMD62qwfL8IFKw8E90tyeLYNbH4FwCZ4BthqNI+Ui/iITa+Js7AosnuqxGX
IPTCksfjEjLMn6diTBz77gznWYr1eJnqMoNcUQE17/29NkGkPkvT2QlwxOj6
KM2Wok5U5J0e068NclDEmS+xyvz8Y6Q8tsdcp5Z7JJkaTF1VigQNbwyGSlza
qcuBdkTrb0u8JisQEGfKx7M8tkgcHNk2nYb18aMMfPIk4XuDvSyAG/saNOnN
9AK07zk1Yw15hVFK9rU4F6OzAlg1WBqgJhbnpqCHND39YpU8SVX88onBU7v3
ggoxPz8RYTPlSBjKYuQA6d9Jtjite2YAOLOrb8K+aRvpV9H2Y4O71EklySZ2
LoVpFgOxVjNblnjf7v5EjwisoQ5/Ft3Vog8JMvtBYV0KZlBgF8pcAD/hFa3Z
s+b0m5sbi7/NBaR4HUi4fXmn7GOzvs+iaG4nIFxJbBv/xWs4zjrwlg1vPu6p
38kiiTaJ9xsMmeGIB6eiDOC4zKBnN0MbCygP5LlPH6CJuZVHlE097ILerYri
gwcU0QFfwLnqmuIgHsPzRPhE6zJSKybs+Vguu92XLPPagw2KxdJ44wZz9sk6
rdEJfXAtLPBWgdgYBkySZoVO+FculE2Fhb8CCRdSXNRRi06vcskdS7E8LB+H
OVWZFDeUX1Gz3rOyKijgwdgj9RK73BR1WsNosqYR7fZt3ImIwfprJSlyIhud
WB1GtSNN1PcOZb4DzHoY9MAcqN6bR7U9PMjQwwQ9dZmNqTVy9dBcynC8ymIe
akNC57l3hnYXIi2pX1fVCzfOwP7dbQc5JG5XYcIy5U3ppxEylC7mPit8UGLn
k3j0/b/juWfuJVMjV/2fZ0bypb2vV5aSJsh14uD5GcLki/bcVhttutITEBDG
YdlredEWvopkir/I1kE0RQ25aLxTCwPzpvrOy+xR9vF8lXqNBTCak8R8Ipjk
Bes9bXO2/QkJAqSgWt+JQyFH97HWY2yP3Sy9LiD38PvOjT/LeWzS3QGou0mR
85mUVqwge6pgEbj/45iaFuY8d/UztsmEzAFsca5WkgTUECLj00kw2L2FH9fp
q7vL/Kql31BwGwXQ8LuD59b8e0H95m08hWjlmzdG3VHPMwMdRgf/DdOWepw1
SQREzSnVRumsx7G5Wj1OeYFPfSqbOo63adV2zeBJh/Ln5Kc5JnY7EXay7Xlb
wlFiJMntIZyGnNbwW6T2/y5Jn9p7cqm/9SAFdCCJQkdsH4d7eR9qFhJepHC2
r03gkWSw5aa7xPAYh1hHPC9m0ca57NeD7Oixa+IiiTyOHSYN33aQZb4pFgiK
0HlLmQoyQeNF+9+xZbTsQucbhqCtIiYmPtCFk0/FuUFy0G9xxIk/dSelmfId
4GCuMFPI+GQd7Sqcezo+S91Asn0/zu0e5fQjqJ7YdxWvtNPQo2xi8QAwYEMj
BpaRhTYoTfrVDRQMZHw7E2ruz7XpNRTxoLYBgj9VWv19IpOzQlSU5HgPMGHr
BXMCqwg1UN99UcB3Czy3IzFwbAla1vz1LybCv48pkFsKkEJo9iT1m2OEz4yo
i7ZzoMnUAmaQuR2tUlw61S7TY+LSeF+tCvSEJo9J4lsimLvz4CMVCfq2yuoc
WIf6HlJrrjDu4S2fGT+xTpnHi6GxDxWnJQ9kGOnEDeTT0RectySEIwOrR0RF
ovzeRbw7oTxiu2MnkSaOHUj4/kuZMbgIiaQ84UEqmrwLLUA8NQQnDRXJXjbZ
nywBBwCoVH2/QCwD/jv6jwCSELwWTjOzEPTyZZTxmSbmtfXuSN4i0rXvcLZp
7pva5n2qlmKA+Mzm2LmrYGbkGZ3OKnHR+L4Y1K0/gzOpGC2XrE/d4dgZ2f8Y
a7+NARzo/b+SYn4NjHkqho4r5USovbT2N8gOUylk5CselY4gNqxmyL9ahpOj
3xEc0AK4mtksAys0NKTfrp/LQODbm0vB2TP9RUz/8znOOtLoFvvm0q1AIfHz
PTetNQZ2LRsZuzBR6Rt3RNFDqH2LHDzQM3l487ZHx01W4Lr0rQFEbATTB3Aw
/TdNal5hxxG1OfDCdcVSYXIWPqTXvRUlyraxRyFciW7XEBkME/nAT10OpsTo
7PB51VMuYPAd1zxq59hABtLeR4VlgYsqa3BzzlpUKh2eo3z3Lmx49ZJHIDXp
CP4rPJegzXG8Ok+y3KEzxWx/HF4o1fhQkMmkOJZa2pXIAZ41zlsdKqiVzFTO
annd2OD6dWA9YxzfcxONGBot95JDtF6R/CObSua7HBn3a9azUZtROL0Lop6z
n78E9CuJ/+pi3NT/RZZB0CoiP3anvnt++8rld3BF+icfvYMi2ERIBMuqFuUX
J/RJn7UpQUIU2YBf6jNp/Pq2dmaJvNVZnOh8H60O4PhVNZqMWybl/XLn51X6
Z+MajOw9s7pSMI8KL3AfNaO5M9maOtdjpPHD4RHfWtzCfazHTOc97hXvCi16
TMgdcODVGa9zSwbVF6aoAOYdZQkQdB/Gam5/I29qshyyxS3CwNz/Td003KL6
AmHjZniXSoXY/5waZ9cNVTnnzB53+pd0rMx3cgl/McIxu5LddGhiOgRrVBJI
hH0lup4MD8nl0AY3zqWnAugu784OoHIOILRVcH/g2N7xVt/mOBTl6oLnqdBW
HSShYa58/OO+wz899jqIvK1paBdDixDo8me5F6mSB38Nkr2ia3ec/OnDSeH8
2avsCsUwEU3I4oSTTjIdtmlHVwuAVQ0ZtGLEouidH6a8FbPrmoGMVjGzZ1Lf
brp6K5BFDmUYpYLf0E1jTBA64GPUETo1ehRELoqbyNChQl2DKFoFUMrrBVfl
XPmOEb5TUfL0Mkwii0Vubh0I0N+t9cRb8ujn4f7yo0zQTw+97LnDuWXwuW4u
4MQTBQXKVEtnbT5XeS1WN0i7aPHQc+K6D5oIYM453spGkkYcTCZcRN3A1PoG
5fsc19ov1OMmZAHx9UGoOS0pNHvL4MuaQFY5L5ZbhCcYp5sre7YiGgaxEO4f
lLwB2Ma/HDmrz18Yza5vA/mgVl+/t8ocI1kpTir1rC32CbWr+EytNdyKIu7F
P/XFKxznkXcOtNEE9DM+AwV/HzF8AXc6FcbVlGMKeIPuIkebUyXwejeGNB4M
kZTrSHEhRWWA8oRD37Fq7FRkV+vRf9zRz6yb7qDdhTbPDrtzGFWXG/ooY/GB
X1Pi5OqmOK3/95Eby4myYd5WXcOGu23sBFvx2M/XCBoyNioI2kJs6vQlqkVr
+c4BELCiDYv6NdrUDyuIgws71y+9ujxgNdRkfYrLz35nE2pRt/qtnv4y0zDS
uHetznz4BZSCD72SZFhrLkEvq7dl/YbGVQHae+9soIxZnUm3t3iddFdUgAWQ
Ble03gXTLQZ52zQLsrRL6TjGNRzx6A452UZyGmW3Fdpxuu13x6/xLYOE3gjH
MIY8fmrAPyJgCWLmXeoaJk8c8FiHr7NUS50jpnFpFOPG61CdXYQxCxJ593W/
Qt9M7vEPR+5W/jEhZwac/bx7xgheIlrYvojCuqpGnpPx9mhqBArQv161S2KM
RdTv5KHwfX2VKCPfBRvDD1A61M0v4DgX1q8dykBTVH2tlKIe6aiHGtt4Irwf
uC+EY46ohtCumVg8tUJ0KRr1J3FPPCK9Nla5yrp975526cg7YtrPQmrLkDJa
tyS9dF/duX8Xpx22xy/K8p4z+sL1NpDAdaz7Cd9409hlTTOE6H74wooBXgmV
1BQUzCD+4xgNYdhNDChv4ucfIYl5l/afmkysDd7VyKPI0kkCxodLCTmZgxNZ
1UPP11FVbrn51vZn9GWbuK9FVF262rF/m2uE0k9/vteZhGB34kTZFmcOPZgr
z+dHE2cWQ5qJAJit5EA+rTjjKTJBm3zqgHUR/6TkNC8te3vzBAoghu4+l0zd
o0S6jeTsS/uXWN+pqvEk//CISDEX5KglnjmDn+/NU5Be/xdGILgalVsS2Jvi
6YUXML7kwVDuhhUXmrqIc+toEUDnPkuUDi6yKdS7Kj1i5E7FpKOzF3oujQO9
W9zsr6bezdiNl6RwT3IBPr4MjfuJxHIpTqRwpHgTrmtI+4jBJpBe5U6Aw2tA
3076i6g5fbyVqUm9sPaE7az8kY9CbJNk1W43uIpe5JkLvrEjjWsB0XdpgJC7
sP9pL9ai07wpCtZAwCu1F3hGXv8JnaAB2Wfn2eOdL1XQdLGWXKjhSGc9eqEG
GfPeu82VZU8A36wN5u2iUMwm6FToZBIv9bs0IICTMOvk6RcTrLhBOQAFr03R
MvAYtkr1hkYDNx/ByzVzFvcTySkt8tdFB/Yk7+BlADKNurflGcKsRT7uIIkL
OqzCXKWrhuZFxMAzizKn9Gjfkxxm9XsrDPptpD1SRoaG+5BzmMrjtKCauOrS
40O4IYGSO7RjCk4CKdosvevTWGbqgxmdFNz+svpN7jlDKKGqFNMdt4vjLFnC
8g+3U5U5cb+tuyAi9Mh8iGv7wJSK4ItTmqouHnaM3AZhvOC0MY3hZigEDEbN
4FZOPEdqVwCNyMqQtmu+pYAhcsty/aVdGMoyea1I6uEe5Ylu9+3KMINWKrBd
m2nCzsDJzLGbHCmEGqOOipLR7rH/e6JWCnVkg18UtZvQ2er4DkdvWw6DE2Q9
0mv28bv80x2uPos5UFH1EicQ7U6ALkVPNhFkArt3190qX/+iFhuM3kEV+HPz
KSi5euPZmrhHlX/p2NkfXi//EjuBKUtI6YgSgojblmjN+InQmzb0vQsTBolU
8UHn3xRneI3f1jVPEXp22vCjWBxpwR6zXnrGCrTp2IgwJLcZcQaET0qhWpfQ
qKw4LjiWgwBOu+ODpiHflsVjKrlIS6hBQoQ0c+9zTNt5HRoIug42pYRFiNOF
XD9JdawvgE+4xMkLhghlmn9pyLOF3HxjKouEMC7nhqpvyHO7UqYTSVd2hA2r
Lb1A8kWoIfC8uNTxVXbtJrs4Sj9VdNrcNkirICJ+vq6wdivEbCjnuRpt7GBz
MtIMiCCgV2kLF5fZHDK5RkgVuyN4AhzBEVivaeBuMa4pYW8y943fcSyLhHtW
2M+1vth/8Kju2eG7vYzDqtO+IHYpAeVgw/5+qopjevtvNVYkuCMkX2wr8zzJ
3zJ/FP8kKmx7UlruakN8sB+dY4bQ3dTf6hFA+yrZiGMF3FtyoliEsfXRzvMe
ZBJGuVPEWLdgF/Es4t3ARFYeirVAOYO/a++VFtKHSSXSmoctffwAoGUZoSLE
/QtrnYVWf1oiLvBDNV8U6V3t+XgE+DVTb9CzhDdV/F3p3HnK+5l6IspQBAGJ
EgPLOq2ejvtEJWy0CfnpQBvI5Ik5tOxD+GVjbN3099tK88poOkdGqsyTc1DY
dHRCv8EE7redhfVdcVvh7c1ADKRB8qxhpHxvrr6Lfn6FgrGU5ViBqx0hA4aX
cDGrjlVaWZWm1fLqsx/XembwqTdhEQmqFKI02XyeokbO6NlVen9f2RLERlJs
9hbFodBJWF7EjlxUsKs6QPCUfemVp2m8EijgjOpVG23AzmFc17uvZil4vWSw
gCxFvjZtXPxKGIii6H1leSGtlYeEXojV0rDC/N89g3cbzBjAotASjEogVRKr
os7HzKsqgS+AsmHJVciy+WthDUDoNo8i8xL7rVlfvgS9ttBZDmNeCyoZOnji
0nGzEgK8RIL1hYVHzdogN+RPE3WAjEdHeSkqgAvy6R2ExPOvjzwUBp97hOYw
VXFiRoO8xE8qI9AaJi1niU8mwMg7nVhb3hvgcPKn1bsvE6L0XihVU6p5cL3F
Yx88uSRu5jlqGm+rzto/NQ6hOiGYhh+DTq0EVRDgMPHeYOxeNwgUTxUwlVAf
wOkG1i7hGtGMOlb3VmK4yqOgPvYeyJ3R78VM6TNbz4EnQcLMHevomfk680eU
TZDOs/suMlkM4diegyetAFtSF3M4OS4dV452nzd768oK3udD74thYUTlKD6c
W91Qd2UU8slN3lpadlCN3FQDen9t8KdTq+WBUMIIQq5fN3CX8HEAYHJXUaxP
m9cX+/aVTb4Xo59cCVh35jRsG1sRIJBXDeJm2ocRki20JlECkktcFSFC4YrX
Cl2UyudW6ShATBTikoFV6v/6wYmgVTSjVDcljZpgnWZSwYVhDrHs7KxQird8
Ebfqu6cW076nVWKQBg1W9EX/JbWrM1ZKU2mbtLjDDY7jVDk76yIMEiX49ppo
ACq2kNuszcxWUeKqVyTLQhCinbIRzQhYSnstAvtwoB5Ucgo6jsR+E5y9IKIT
gMRBVAvjfPSuVD4JzjhGKRPn4JqgkWEWFRgUiS6ZdHHsLYdnEZjty5kPKD23
LYcTNPWBevRR7c3K6qN9Tb6g9lPS1RUvnjKVMvm1jD2ihBdia1FvOWIPY3Pe
KGeU2alPoNMpQCGYowjmHJG3xXjbde2kpiNbfc7n1HHhnM1Bd1a9QxL9Uoyl
tmfnbzhD9U2d/BEfWztVVhJMR7Phdxc/NP7zLIntvsUGBswsSRYOGZ88veCi
qI1wpBX/S2m35f1c9xdnpMcIANy6BdPVGY623uj3WWtazKPx4tStr9+/uMX7
CjsBXnMN189sdrhgXhn18wMw6GcBJbnO1Re4ALCmgSLlwpzlZatcyPWTEaJr
zRm5Kszb6INov/ZTSk40RRThn4T9clTrlvaR0i5aJ2PhaBjN8MqmYt535stY
lFvgHPIJa6tZpUya25S/vKEoRgmnl2xoW/Dqnt1Pj/Lah4G1YwZtK1XeIuw8
rlAF3SafJ3gabXdrmDMx11zWDuURtLut/LxPBPnT48n73JkjM5PZuHA+aS2N
ZIeCR8ExI+CcpzwSb8pobC0eb2uC9H/zML+Ad8q71egosx9PYI//zi858c/5
NstbrFbYeFbTwvIXYk60v9mjhxwsOiba4cgAmycLmU/ACTv+hl2mELUUm/Yd
ser0l+8Q6c+GV0VcKASKshezY4Dnlul5dHjW7NR6YvRxmcKnEsDbxFmmLM8k
SdNM95Z8JpHRGGb10VZloc17rL4c+IToW8gkxQKlI+u+4xxUrmq7feOo2tJD
zn6QxhecmuDiK0xzgJWxzoiCkiJqay4YEOo/Nq14BUfXOTycoOsjwteU6C3F
qxMZS2f1TENo+MVeCqrlVas91gCw+uF8EFiaujyR2geJc5KSVwY1jBsFMeu5
edLV9HEENrVPd0IvlrLqvQwfQmdmLWhpZ+lhf2EyCE8lOHn/eyIOq6n3Z/c8
0P74Eid2XmVGVWXO1LHkvM/2vmtYQakYDmviVRf/38WzK80LG3bDDFpXuXhw
3u7vLxnRG60eMy4OIH0YOG3kXZLIkPvWE15jb44aQu3oVDqh2TJA//+wB/k3
MjoLOD5wjqgrvY/OQNodELs30oEmhC6outsAkFOVb0BSpmJj2iBTt1fmVqsK
UzTRZLd+iiWgmb2m6xyWPCHfyvsuiQkm2twLR18sV/Awskm+k5YDq2mVR856
c5WiWW1N+KRZLeflLtFkYaXbfcrA+xN/eg6qRsz10Q63pffEHlAL8gzno/b7
cMelcaIFZHkBGqevs28FMGqxEvSyirG5LAyuPU4fzhnstjZD8+3G27N59Dii
IbofyX5DfBW/X7R88OrWkY+S9HW8LQFeP7E/CnYLRdPzPbPYyjehmTDGVpFh
h+j33izBSNBuJ0X2+bRTY2GU0EK4VyGWth9Bqz4s30E6a8dx5sxoDip0W+ib
nEfnJQzl21wElVB2C4RF4kVZsfqxAo+gTha7R5X/9NUsmhFqKJqsuSNZzBYk
AJCmzeyOpb5KwwV6pfgu1CK+3smOyBBS2yk7Bqa3znX7erQppEZv/w4vnVTH
0+R+Xmr1N87K4LR0/LpomdYBEUFlABJM+Jx/XX3QwyC4Ymv8hKZx7CcxIHnF
iTbASl0G5zRHsgII8UFz4n0uVi+7UxSt3a0xNaUmd6yjLjRW/OuI9TQBxoPu
WdfyyBdFDjIyNk0m7Y6Kklm8DxmXg6e/piLBW0on1uqIVDy2617umt11OM91
9eumO2YyCA9L606fxqhjTKZfLtYct5tjldqBTxreOcXR7JcKrLZcvixfZ/yU
S9p+G/VjTVThMO8eymBylXVQwE8I3bmV05im+RBqC9Fjtziv5rsXGTF3qnJn
AM1Xw3FfF5lQaLOnCGAcsyUHADpMQBcPIkK18H8ERdAYs3P3ECK9YUy5ZqvJ
gO5g3xR8eQh3ky/+hHEfqXmsxR3tnVMaaDLV0gCk2hmt036yzaUilB4bpOlK
8YGZe1f6l05HmbJluQrTquOcSAXl1moTouNGNDc5QS0I7qXMbyoZFBxNnEuM
7hQaT2xSvMAeMa+CAr15513S72c+6me2AeBX6xTpdwAWhj61apmDtAp8/9St
UCnNbgCfXD1HOTlKq85jK1rXbBYcRYc+xCrKjmMBTaVnmfZeuMwVuNh100GV
IHK+E1/dV1l1Rj5HlIWv2BNRGlf55zqFRLv/KvJvcB+V34h9Qi4lL4YzQk0x
OGAkT+jq7w6yOl1rk4pshQJJa90FVIzJIq2SC3F0jiluj1SQofhTWZ+5OuBo
uRPSq0j4HfP3LGMaLvzyIdjSdwWCONhQZmrgAwtgBk9nda4Yz8oqNKttLa2n
6xMM0TQsFiNaTi3hDOjPSIETr6giHdUdrEEQtuEqOqw+60XwSmsAGcZ2fdaE
6kzuzxBILJ49HQ6KdMXnI7Dm4sJ0IJ9Kb77EmWZAbcR49RgUu2ZJgUBIjNhf
Wd74Rq5ef2ZIgc3pjzU6NIPHY191FroksjelniWmNVGe/4zneX4ZtXGMWVxk
gdf00YSrGwE0HwWuH6gPhPqe9hqmYjWQnzmAkTdRf0I3AaEvHXzpygxDSr/Q
t9OxcOxAK2moKrAFSFe+7Pp3cvIqUPT9pzV/5v66kK1FCxJ4u/uurU/vd3zc
4ctC/cGVAd/yx/hQNiRVHiWCwF4CUjm1EX/yITSUwd223N3x/y7S+8yFLxHA
5/a4/lpcHMwoJQqvwxLWUsknQApiQiAV6coyAZ9ltSrZL8jD9vSl8Y8gdwho
36j2zZwdVIDvd4t3T+uSZh+4XWZvf+gVrMOjgFgQkGVrDMgjLTu7sGNHMFUb
37+RsKzYbb/apFF4hTU1Tq/l1zT3p2KYVklmIO/mGhVX1J5tp85GjA1Rp6HZ
CXllSeAx+NJI4spVocpank3NWyfQS1EKv7c3Ne6lEi9zqjBCSIQx97F7iYK1
PY5LWNLb5vhJYdXSf8SG8ocAK8FG8CwW4KVWY7ekBcOA4xzImjvG/cwmE1By
xUCc6ZOVJoYVuOdaNpetJ5DcSztOtAwspq7jBPe1xcXWjn1fgYsxsjUZNIsu
3YrRO6OT78yMA3Bji6D7iiByHdvvQXId+QBpcoK7BSb/BL10qvJHUBDGtpKh
T0iZq7Zb0sZQDpmUWQM2hD5qyVYnu+Z0TFVXLOinEFi+uWH+IaeKZQZpTX/I
7NnrYuIFZIPiMB97y5AnvbenIjumFbjTcPKbJELaC2TT5dxVLhfym3s0wVBu
6Z4MsFpKhuBd5zbWbysGzznZYyec+oPm+yE9jPWEB6ugk1wHCUypU0X+B9yq
ntslH6vFvBIiYoIe/8TqzfkHj/IA7EEfIAH6ssz7zRjN+ycbJDJc8xlPMidc
UIeLahiPqLv+RJlyVqRUwJIdhy9l1R69WtY2k/NS2iCvGfLR6PxM0oFvW8rn
0vZhJSnHR0sKvX5EC6+OiAHotSO+GB0qILHOv2k3rXW+kC0ADSniLT5MjLto
BuDMTrIQ8+RyDefCTOCiu42OJNLdE2akQi/u98hKVr3jU8dMJBzmYZiuefxQ
S+jvt7xRTu+exCOOmXfjpJznFa3mgyPqSmUZmFr7EHkRaKZ+TUDns5LIwF2q
zZU6Cco/BTQ4cHJOkhL/SpNIYHz0IqiI5fJbkEk7QOek6g5lAWwbvS7pPOHz
rzWMZuAaWsjxGTs5YyhlC6hrhu1QZE0BPBBvggOzYX5G6Y+aYELEIddeaYoe
HXbjAxWXYTsln0tqMPAIzwVXBBr0XVnOSd7r9iVizpmEZtUaM4m3rVFmyKmd
VGnqmyZPrZMp8ytnNEmHuwV5IQ3ImrkYMC4sHRLa6sgp5aYAeYb+T5kmH6BO
KAEBiNTf52DHuEDsC5zz2XgV/h/aE0YeBJRC9DfmVX2nsRSu2gpp8KhVl1hW
Rv384OBGeGfSQ7EJZ4tnAeXrhP97bmWhuEpgcOTgxUgAxtVHnLSAEvRltegN
dWBx+Ag6efnHAgdDbcRYbIfGp58D8hd06v1dzpiC+ttNfBDnjZv0e6gZw89c
sDx3BT0ev8reN5joJ5PnFacwz7RKxli9j9Xmu1xNZd1lt3JCEHpirbfcMmXN
zAlKVXpvRKLoIm087ADtw4xJyDwagzzy9Kdu0uZUJMj7i57M7bDQTnxIZh8O
w6dx/hFVf2WBYWU3c2u5i5iXfqqcFViYXj94W+7tK6DFHvzY5rwrljCOrC1x
5wxaCSVmpdlS7AZzi07Q76op8C657FV/kTD3HZkRq1cTSVW4zYschgsipfTZ
wHH/fEy8FKzbbul0yt9P59Cv3dRIYqwBnDWo0vCzTkGcqCFTELjIC24Se1qG
E+R/GDPU3ZrjLlb2Q3Q6djDgXqZ/PLy8028kvneTfdU8XFXB8mHBZhDdI5v4
9DfZbUMPjU6rjegyPHJcfzsANzq/lpTX+hgKxqxvcxA+x0IoTxSMXYtW6tcO
oHJtjvXYWDDjHytPG1TK9PLVgdeq2STWsm91UIZldsQSQa4vulUYhpJEzQdI
uUUxl+CQ3v0gS2jxnruhYbBCKAndUGiB4wXsqo93jyUCYNIKvIqaV7z5oYoF
CU4luDwbDusIxxq+Bvl07blulCKlXDQVONY3wcmwwwe0Eauz9Wv+sZDyxXHI
6X08XQ8RDYEliit4vj7SVedUgiOxIYoeMj48LkKaGFvaYid9yhQsfK5SEKc7
+ZiGRSfszs6ju0eC/xlzWaTEpm5zxDzhLz1XolCe8sc9NqAL87iOVIrsBxqQ
/EU3caSoCeKZfAgrAJ5SAYSuPZLc3lV85XKE75bqqlcfLi6IKJENymPzwxac
VZRK16e1TrOwoqrt/rAuki3aLag4FQEtJv5YrMot9MWxns4H5igmbnbIQUXb
hE6sl71x//PwcfTa2RTCyaN7P4rllpAIBulSOD01JgsMWZ/4GMCynnFV52FP
nr8wy2PNkmdobRQuxWf6ghHEkSwJ01nUyaHsQ5SyOVw9kk6ZTfIuu0dKNoZj
IQGgOprJTNKZASlBjMhOXVlj4nUXBxyP/muNXgAxHZAoFTbaDfGMtVpCMePu
CadJmTRE7hmxab6Xp1sH4EmHVdM8qqsA1TKT5rZS26sLCZtRobUV2zUTACYH
jOYRnmJqpDfkTS1qnsooB6jS8DR0ZJBgtvqzuysopQNi2rvw7G18xfgfDtDF
/NpUhflP6ViJS20VtoPPcVBsOEMt8n05LZ5/bCkrqNnZJLTiZ4AfWMSV7yHs
DpFJb+XHvuGS0KgAPQilo1UwDyGU1ROzfc+qLYhsU3aB3eG2AEsNPgA8/DFP
JZALBi6mVMRt3dVEKV+X8+Cbwb2jlImQCCiCSA4OIP/VqRhsO6pVRTO+pC7n
a/ZcBRk94vZ5YpQk8gSEZeLRjtWzNpf7ZHNUk5LXab5ncdRlHDDUi9uH+52T
IUuyL/E0cTaxA7mrVYPyIugGwgMmzytshkrteVSZTvTJMlEyMoO5yQ6/vBaV
kPYkhJUmFi5btpMSLU8j1To4CotyzPQ7UBhSPWbZCkJLa9LErG1DExHpDZ3Z
wabMSTLjD+d+Xe2+hUCUVrmfvh94UJyM1SE9QRmYoV1knm/sqxT+oV57Vkja
ecM4r/XQYmUEJefb4OGxoCMkhQE4btaixLkdGwW2DZQ9MbhJX6uXqLkkggTF
nFrwFZ9+UP0rG2sqmcVK2KT387K7BXCDfDnc+lkHmyTH7Z51WdKGiRnBxKsB
kGfwdNNVSnIjXolD+Rzv7tI9msdeDEnfikOMiGffNh2l5slMAg0ajll/QfwH
XXy9Zmnh2YJwC4CwVrxtxsTYP99oQ/GtqlDOPYaoo0RQZqcPQtVbImnEf6Dt
gqdNCugICfIMvdxriSelVpSVGO+zEPssTWTLVYAUkhkldPTTbmnCm9UpO536
wQ/n93HNIa00Nfc/XuFuLyi/JlebgB4xVUH73Bw3zD3J2CMyZBcWkXkzCMPY
ru9Ebw4irQculW+7F0enhAxKCBHGld756DBBYyDbwNfDFJmfW+7I6fOIwTw2
Z2RZwg+PxLjrXICOzNI9LXOvaGM2j3IPc5yaNPCsXsYpwXr+SsGS0O6dDQGT
KJN7eY0ukaWMhAfTFXqWMWVGqK0Asthi7cfmt5hd6PA38YG9Q+3VNLrmolBz
00Axy3PLxviA9DbBTIG7dJc9KIb/4XKP3qY6UdF33lyNUBF81oMGHy6hLSaW
CYvIq8CflRrv0SaVHMef9FGLL3cz6pcyoxnnqMECNcJZYIsrz0Msfeef4vfW
2wW03mfXdY3tfStQCCvFZf7N1QdRTsEOXKXw+ezrcnarSGJF4gi7OPqAAVog
zN0MMUClnXfwR/rxLWGR/efW6bcWBBxDvYNuSvj1HjOwr9UDsvQbKHA2ya9O
XeK+SmRBsDgb2pBexCkZ14ieXir82RB5vyfIjc16V0g5I42jnchTJRx49Alf
u85/X2JlW99fV3XqW1GbFX1XtYFUzy+Eihqltg2O8JWMEOqvhru53RFN1hq/
CxlfKCXad/6cjUCP9TmfcZRzSFozN3kSbOZRR3CdhfgslNNxYR9+IowWBT2w
PSS6EmXkD8vIEEDVO93K93VU3KNgGIabNHzz3cfQSnbsyoLPA4LoyECSm4Kr
6Ml93tSHSFzrdzN463bFL0vbfTpJ8UTN9WFqYdRs2wLrSvFMBVFAqd1sakoO
poK0cMWR38a6fQvTEUV1A8DWddV9/geeJjKIl7Nn/QLin5f0ktTpswWZCTmF
RCSdtz/m0q2ZiAQYj1k+Rm2tH3VTgJTqavY9TCM92PIsptRVr8PSPKszMxeq
DGEoPHC923IPgWt3vYMfQb9jKJi8aWydSFaqodBKjI60LZhtClV0mQNyzc4h
ycJc14MOqRJDPa1MczdvMXpio9E55aDGpLBSJ9+ixZg3qbfG8plRWA8DI4X9
BUD8P+6Gl1kCeVJupC1JX7NyLPROZHsScbUUMcDH/6NwJvCxs9qHRUmKTs3m
ZOIIVSp2ZyCilXXoUsSJtSzqkrpFeuWRgYOnTMQltdYVWdG9zi9gpoekZbHn
0/+kHQtQ/L9qbGN3z8EY2L4QPtATRHPlzk7zsyambyrdpBF1fQA93lKg1axp
RF0t8xxIs/2guwzaqCBY/OuLdqPtTUuPF3vrNJVKl4YatDyZPKZOoh83ppUf
Nzz2mbElyaKkUR3KHp+KxiJiv3YO9DeSaM8GoMAgEBE3jIOcfbgdt6Vk2RzZ
hcQ7BzxndBXCaCxCf+lbtQkZVZAHjosSETcls8Xhwwv4iuHDOmJ66zKvEZD/
5YZdkgl1XKWRHfv5VibEK7gEcFvZ2G7HwN6oxuRZyFs42SrEs6CpisHAc7VM
INpjUGswyqtaRvVpjUb9waERHuOmx/K/XVUGmXHGba3nwqapJY7URgL4D70U
ngYvgh7dvCaaYVeXaDceMTos3rSchVxh+fUOl7/cG2OuesIPW7h7GJ2t5D55
EQFtvTxPsrCbd/Dvw/JeWR3DcYbkhVF1xNypiQHcBtPb2fc9BW/EaUz5C0Fs
0KDA2yfZlyNvesl/joEtUwBOsv8+LAy/eHSCs6Is4v2m5dmnq53sLUwnkyYd
xOA5VMxWWUSE/OamEezBqWQfhxEnoe5TBuwtLAqs6HUPa7gJv+BHy0doJvEx
W2fw2Ip6UZdAd9j7VFdsvnBT6zvrk7ui+/l0qXhXXSq0+agMg0xJM0pDMo5E
Dp9tex5gEknXIiEHbRJ87xR7OXupaIrLggvd4s7L+pr6IIYZbuVZcmMXtzjA
46J4EOcuezqQ7IPD7QnDTSl6JMVxHjcDKcPza09gjX9LnC9yT3TuLld3v1iw
Ptm48zAsUFAsFqXVGh6bTyTeJS9NDsxD1DXINxdNabfmAK9WlWfRbaRmA8ox
fmUD0MDqy/3P7OWk05+zkHNUeg4Jb+F/PitGG7p1342VnGaBci+yeSPqHorx
dwWtfa6MQ96ygzu9a4YhZrPwV++jDBuKEDYc7o28skupdyq/gKYm3DhKRVjV
3LGTwWPEbgYXGRZaJhhBbb8Yek3bs/sUE7nojJ+qL5bvNqDaFSHOH4MQ7L9E
jii8SPbZjuyjTHT6KZJ9tbpd2bWiYo91Pll09XMC4qhW3hKttq4cooOyUubB
ejCoTVBpd4LdLCg5uHs4+Pxe2DADrj3kDECCiVQJ7znd198FnnSeaZJYu2yD
9/nICceQDlFs3boV0396/reUQtAor02BBTQRXEN2l2tWIUv2ocG8urqBIWPd
HOWBhVq8Vk6ZxsJ/M7NnH+r23ch4jRHpsBOjkx2wWTYaziaGl6/mo0JFjnQz
7bolZz1ooVoHVjH7ro07iZGzl0r+ug2du7YLJW0w0uddyvetaTUaBDE15qvB
T+3bGssaCXJ2nYJUCabAJWz8gOX6DcB4QphIHT54wCJOapwnc+fjZu1OeDpm
GhW4nFOKVJg3Zelpwk8XdVfZ9BoFGNOFXOrrX+2TFC+BJ9BQpDl5EOb4u8K5
BE85EMd9lWmwfsAHdG2hV2W+A3GBu4AKyY6b3+CcKI8d7O+Uf2/PjYhDmuRh
i08Q6HaZxFCWPru3lWIOifRCI7CbFqwzOeNGTYWCp5r7nN5FcLdB2DEL13YD
JDGSC8vOe99rC81HfV/+b/R3pfvuFak3fFBjzCTrR5VAG4S1yLZj5ZWdW2Gj
hpgR0lD2YXh6pcqar+u9eO46JSM2bHuqvlyfbwGKIY5Ox5gFMdYP/CWrQdRC
SYTe42g1B+SaF9cPaUpuziWJ0y1DkWil1/UXWstkQSs5b7xIHj7cGZzdgp3/
ZGjgWNPGLD+0+pW9B24OoGkE/UN8W6OijaMhomaKIkrcFin5KmdSVWhOp+BT
kjFMS+LHOmzpk7h9K59CzwshsBQEAnqh6Rf9r4l3/iXq2hzGgX0hiO7Gl33i
aDTE6ADh4/nsCXCtZlzw+R/SiL5DHaWkbTKV5qGkeGGKD049DHFggWHWLrjj
1acN6iHOev+5WyzNa8rIw3eN6V5Xyc1bgWUzJfhnT313NkfrwDcqUrNqWZL0
DfCIUS1Ysu5nd2j5tKMA5w/mVCPHKGdccNRDK80Yx0Z+DTZHCWTa5dgghVQo
EzPzC9tIaiVarvtSrFOo229YRhv5SUMzNcBMEjbomLqRB/LOzL4cy9UcKKhX
LxX/PEO+xDn8GLGEBY7h4tVVD9IS/cy9S+LqW6T6n56UvOP8zOCkybdAlVEV
g/t75uUnC4KVA5TDX9w9oFIek5Hrwq326oddgQHfCLl6zaJ++L2HeT9F29ux
aPr3k0rQG6zRzQARHO1Y5vGQjdJBXwoBMJKNOxhM17gWRVpxSU4gPitJqevp
InBZCYWM+bjXEd4v08Xz6DskHu/IGf92KAe77t3k/JVJqtHJZ9ETtuCAHpnG
tog5ShX+Gj0fbxiHFs41nfBBNA6SoOCd+k4lYG9kYZau8I6ZaYUm1FpddVY6
n1BoLiPNYXe33tTgCvAyWBh040O0kSgtzhKkNWQPap/PNn4S1rdYWweEXjiN
9aYIu4Iy7PbFu5EfyZKafSG+CjPXQU+Zvk1qnvQut/WPIDr44KDYUZUnbJ0o
WyOoYdfqLQaSVX6YF9kmHwC5ApBqNc98YzJm0rY3quasnuBXC/E2+Y+t2R/f
hGldAnMLHfvEWROXMlL5fYZeHtNBtKYg73YhWThvDDsxXjo/xBTg+jTxeWnA
8fpxM1fXm1ipV1YOomm7rNhK218H/Ay0h0Ab0QZ4IpV7rT5WEko5TY++44cV
ayWl+cJ3kKBPWaOViVaaVM1wpXor2CbElOAAF66r4q7ezXUJHCx3yjb6rseR
l+KCSn80A0ew1atpFKdNb4zivbFaJ2V68jJD8WTFBo12iF1ScQ5VqoZ7g4Hq
fOYdvsFX/3L7j1wNarfUA1CFhehCbQnP8jCqYCYI+7gEIIkdS01sFvaJ6WHO
7lHx9Sp6WfDPj/o8DGn2Ov8+3xyCYtXkbqqnBKMunhUAKa8IorInrU+AURIA
9UO7XRxYlIus/AHV/qLQ5yBvhtj7PRmpX6j65impDNbwjZDqGzuEswVQxJFi
1EN3emGGGJ17XzuMcd9XRJN9P/CRFz0W6bkX2J2XgD9DV0wWEeGpaUUaR4ZC
GohjsWyIV2j0YX0rN3S0bVfXFte7aj95YHna6sNdcUJHBigPHu9zUOo3m2Tb
Ir7czJF+FHIi+X6zwMLcWGcF8UjQC2JmZjIrwwzF6veM/DRBeWq7tZpGiJzh
TD+GHb2Wcth7FMQP4CcwwT3tCeZCYfHdxo/B7aX+Xd3Fd/91N1XjDpo9Kf41
qViXPIVkbjzPLxRJN0asd1ywR0MGZgLvO6WsrnPiLCOb/wO2UcK8tCrYyILp
P8g2zTnMub0LQAOOxtMFV7409FURSGAZUaCsxDS934lIHOuiQnhSk2mlQbSm
L5GoWlAnAYun72X7ZwAR1GMI38DbMELlPJtZD5enThPp4+S4J9bWZeU8cB7d
SUKqFXMMf/pnuDXDL7vkgCItQufEaNe+CVxjDw/MGOx+0KTy/w2ogTN4vl9N
uJ4/VuaZCzX94jZ29WenO/lrXiaFLfxWTmFOHdPJCy0HtUMzguUDLSImUs9e
e6C2lnIdayqghevmlwd7uTeLZ6kdXb9nvd0bi1+elFHk4DFYRtI/Gmn5JM5A
xuPxHIhH8WgCKI9co3SjvkpOS67NJGF5wEWP/wCIn+0CM2mKWgk85m79KH7b
1gIqWwZeaciumf0YLfpPIEYkk+BUz/pd8wt1Sw6ATHcnxdQkMR7grgkBSr6s
7tG3KSVhgtwTwruyrar6yLPyWQ9J3FkYc4Ep+pGOZaojj/yAfuna/4Aghsaf
e7L1m8rc13+mIm+QKE+6Gvw1nMbUFMoJ/Jm3qm9PLoT1k+OG14bc40q6FGoN
h6IwiY9zQUYYe5J70NYqIYNrhdRcOm5xp08KFy8EouDWkrDs3zEp3vCOKyDa
xAqLSFsDH6ghgqs/LteadVMcTlA8X/GxINdL3+oSxN7qP6T+gb6Ui2G6EN1A
7KO2IIIt4LYVGEBGxWCBBEfCB2DSMupWCYdVW8bAdbq54ih67RIKegMb9oAh
HhU36NBl72lsDrB17Tg+PS08Yv0vYcYAtqPQFhyuMIdTS/mdJtdhx3YpBKYb
WgNwbGYPW0FuCOcEMFoAofgA17cR9cqlQk9pC+TzmDtAVa71OG5rhrJ0ogZx
i4ryFBYqE0lpqV3iwiqtnpjV/IY3iLSdinVzD+qlkxojnPqCma2zMnf+SH31
z1qZ0XpzRdf7ouNMTYgpYIOXYs/ElWbO1AGZ8bNl9GbZqvIPeq6l4cBbH6oq
UyWCLFjcwEnxXOet6VIS1gHZriwn6N/r0sCbaVRycOR1doB6t0An9Ori3bFV
iLS+MKwKMB+7meUFtY4agxJ3C50tU7NeDnq/KHxrD4T3zxFRePrXVt09G5+t
NiHtjWfRQVN9QLRh6LUxoX5kBsYmQhrZpblVhLl+UamXeiymKBiu/txclUm4
JlR4qLk9cF7zVkekT6HuIvWFnqUhNVaehCnOW5RsExg2wZhhzFhjuOVstL/j
QhMEk/oSGYhtx5JTD5KMSGo+XVr+2bH39k60VhkqVEcQysHKrd8PU+wHdBFA
qo4FTKLXpkZV1iqHOJrx0uPqFomuMiqokhNGeCGqepEXK9KkpwYgC1nw+Ehk
Z9FgHX4Ar5rsQB5Y4+iIhGn7nhuy9Gv21q0RugIqYS8oIpkkUWpHjKfQtDEu
V2M+It1z0j1s48hIkS8b1ZmMs+KaXTZmcGvxZ1+0+ysy39GuErtn15R1ossp
1kgsI8AbDOEj69FWKPYyMVTZbF6fnTs9DWIUwP6l00zyAls18ERTRhBlnlXr
mLNKj9L4WM5M6xRKI72Wbi3kQgz+BslB4kAby3XQjMF0tmOIL3n76tay1ny3
a7XvWW21HLjRrIZGtKf1+HFdmUJJiUj5iEIGmYLB86JSxcG+5jhjwu7yEves
+tzy6q21EMZW4erljTxKR3+j3elVQSc1UZeOzS6hvCPwk5bT0tYdVrhj6b1e
HzEKCfUy0BBZKZOlYC+DcGO45uY6oD2kgcumzOLMTm0JweyBMUyxymc0v6Jh
C83aDYDo5YGMkfnJ0YLZVdehzImAwQXqP63SRzuRYI0COMQ17js3b+TFhAj6
fKlRvM9CddFZypDykALnolIlAB4QKNyAD+Jl/8Y8V6BanIY/BlzAx2uxEq4S
UJnpZOXnO0oKkRIRhyUENSfNOoGpL4bKwLhkp8VrdGFCnxeyybxoTUFBcVJd
M2zxsGMaTopnGCsJ3C8yEQnVMIF9D48I5UdbvbQyqW3XNuJIcSt/Dc/1QDFA
mIE2GCCg0aYjUMi58af6SWnElHvLmmSPrG8YSZNzbSsYgw9tLZIi9kntU1rN
o9BVq/xE030bWk2Kcae/O4xcZHNf8IpdbU2vH8A23uygHjbLRkNMttg7PxBQ
pFOp1hqr3Uf9kWjBAudO2tUPbOUG79WuLKkes3ZqiBVYnNTrw3BBWBZgE1e9
r8n9in30VzUNziEicqN2V9C9qU5XEDCYc8bDfaIsBH7rw0FOzL7X/YANGx51
wRH4XLmsgOeM8Hiy/2eKk3l2mxilhaakfCeFx2B8aTPI35bejXQCD1WT09XM
XgYIuT3m6oYmLaTNEZdbECRE2f75G5Rr2tPENEJxWI9e+Cf6jjyHXUq2nTzg
5MIPVVMhTY7Q3hsyJ3mve2tkKmyqLmhS4OhZhK7J2PdNYFzgOfl2IvvqJ9us
Ml7Wi9G9jR2TURVFdTIHxGYwdTaQMWcMw3m//n8Bp4YPHo4yfpTEFlhfOLpJ
lW+F+rvYAk4LA6U5tsGQk5cZvAY6MrQnizeZYmTT6gny5JztrdbYnL/MKq/E
Cmffk9KY5PWXPgpEmDvgEbYZ97C7sUCqlEuw1h1c6rOauaRZzvpN5Kw5duwJ
3McA9Kcuz3naDTO7C3mOaK0uZW97ftEedb6tDRiM1fhOEr7VbmOjheyt78bP
LnVHryqdSDCjdtS8fjD36erA5Ij/CjtZlwF5KrKMTzraZ/f77EENxK9w9T29
NlZhZ54xMc5d2qkV2Q0Vmv5Dm2OTzktJuebRGm77VaTuczmAD/Mm6u64U9OC
X6qUETUU2Rvugvr+DToiqeclhATeZ+QI0KvM4ba2QYIe7/n1ZcRjytaMwIK3
QidVFMtbVuwPqMpHlKM9s/0wXaeRjjPGus7s2KTkXVp35gR6ILF8hu1S+Lq0
dYvdDe4IPaj2cdFg/LiRFJ+hHvUdFNWTfUWW6LV9SOMqZoSpYeHtZtVNGXJ0
XEkdGzvelJayaw3LmbfpUNBXKjU9Dd6uhsLNnw3b7BeUouE+yBMIB8TUfKan
z7xF0Frl/me2M/+tFTGTnqWuvVj2geqGWAEBAULF9Oyqb5W3rN6BS81FeUBn
+WYnahIfR3d1SV9LkR7lGMpJZ8v+L00y1nSdJ6HYI/R4YRX/WhJjbBbSrRXr
iAsR3RPR9rKwJGlEvkUMiVxon4qAvhwt2rl5zB12+3FJRktKw42GhVwmayZZ
ykb04SFBIhIhfWXdRSXh1poK92zFS7HxRoM2qppugxsMSHUPVr0yyzKL/Yta
eL/CmAhUEEu2DX+jJMBa82LgB865GaSb5rk8hpznupLcLsC/3iWZ3etgATDI
eXUmUlPnD2xd+lPLYtdnmziVmva8INYsn+unnejrnKIoWtKoR3G7QSBvPt3b
Ht7Tu0sNtQgbdSEeQWufb0GKyKrh22W2JU8LBhrFXwL1kvZSZ4HJiT+7gSNN
1do60o2+qbI6tjnFSvOx9uNjsYtsKudFTeXpqN700MDAe5IAA/7adTEIxb6P
jr5FOJRI5gFdtSiDMIqUx48ieiyNLkCHRxvMXlLPIQK7/xFJWKbn+iTn5Dra
IY3kFt/2bFaGulVdWcc02SvyiEoxna7j+EYTtQmb3yWUyI/DKu/Q4MLR/NW9
rDeFr3I587M/juWAz4S4NLFI3We8h3XJPczPV0p9XyV2WwZrFjr5aw13Yn/S
i7N4+1C7OA1JrfjtsO87CQvaxXYz9W/j2V7bjP3Hk6rzJxtmSjYJPoEPr82f
8Jy6Qmnawy/KU3/OTckq4om91G+zODfVYwHGYOj3p8vu4Z/++d0f9+dKALAF
gicx9IJZqMsUMr4tHk6xqfIlTyboJtDbsHR5YoLfJjnRlqfHalxa33rJOp/6
xmWFs1/090r5VpmQV1F+RmCOfLM8m+jA+c4i/PUWa3QdMcR3K7uHgNSnd0Wf
lwSuJMyiTDv5FsrLLwQW+dPa0PiUQ7HGqn/72eT3YUlPqsGe8Z5ctMC3Q38p
LeRgub3QU3xPZO6KEtizc+cc7mqFBRHq6OFQLrDeSGdvAAELGu1SchV25zEx
BVbgKHWJviGuGBm+gBpXA5hVsKNn8/Us4/+/o+HdxFjF0BOXpN2zi2NN0mJs
9qVL1iIhlGsHhxnpvdUkz/a7Lp9iRJmNfx1eCgVnmeV9Q1RrJoVnuB+Q4BQ8
G083HSODIBQUtwWS8oMiTjg+tkDmOEihGa4DMg3Fk/wmq/TaO15sIEICl/hS
N0pbiszXlanJ6XVzOxpFurSsmn98Stps9cVrEggsuoowfzpz6npKc9uqIsha
RrBiqScyakiQnoKyXJQUPGnN86k3II/NdTaUTkkLW+icsW0wWrD6VtsulpA1
126WZGOGyrYyb+bWlNWUmChabbc8xib7GnX07qtm5DbfGwuj/zXBQfrt2V7q
23IeljJ1cpQOJ7Jn7dkgR/lg9AZGPZg7HS7XeVWt+zER/Hupj3hu/ihBxAOv
n1joxJS/7SqouGBJSz/iIX533CqDwcBfvbYmplgpTLvF5tyrPek4h3Fj4efg
bkFuzWwS+EUoGhlegfS2RXKZs2p9IHS3mazpfjo8lDqiwtKShtRn9Flf1wOq
RDLq+adCbhGssFDf0hdQo136SH4mIKP1ES7gSr0feZBqmPA7WE8j/ZHIBuVC
pjIn2MLVtTazs3HYDXJeDbnJmQiEU2uKD7pLyV1pSsNbYjbQ8v7XHOOTB5uF
iBu2rtnr31L6zHTlIVQBRfdgPdRwO18F/M4IrYJn9kTC/73b2ZMFYRkRotf/
rzNCO52bVpMktZSgXZOkqazkuBP5dXCduKOboF0KzXCqF2hb6NfG9xngJVsp
EUEoZLWxoKYJcxGnKGhRiO1KAoskSdMAbc/IjAvywMXDxMmzDWV1qQ6Mlbgq
cd8itGBatxI3gzkd7u7VbFYHxYUm9AQQHfNvZ/tiQ/vzHQKq8s7W5HgwVC4I
NaGHKJEZCE60OJtoyc7+P50hve9t2YBm+KkeybWIFyp9S5Yxb6IvGryvZAgL
i8Wx8HMNVAKuy4DnKRSAAqPcPiafmZPVbgKHjVb64HNXC6vz8sdtmlYlRoFK
Vf0fv69Qti19fdDGB4SZQdgg4mwr84rP/8nXATDMPH9BLkNbvqjsiAwx2pio
mRJrLr4jkSwV91PTkzqj6sx1GRf1tkcChvv7hz7Ttbw1TpZyWxfwuITOXavj
PumBNC0mh2rDbusqR0NmvU34yw5Wed0QTYZ4m+vVCUHDgWvmp2Pp3tGlcR0G
R8AiTKdCkFjW1ZSdhUP7UL+5zmNv3hdjL2Nwbu6BhBcd0Zb2v0NwQr79oSTm
GdKQdiPIUFFcjXf8X3yeFD3BZXoI5PBfcchimoAbPn80A6CdjjA+6+fFY0Om
YPc0nFORzyajTvVFFAu5rdk3ivBn9XGlSFvxskgFIRIE3BHdQCeQxl4J/76A
IhChXcRidjZY9L6fF1DZzVtBJzb50qRB0z8z8Wnlcbq5GgLFRSD0y4XSoZ43
5HSyzGF81PoEkguwz/d8q3CrRc1CikJtFJayUvDND5FFdYw6vVJuvJr1tIFE
wK9HBDlPqgA8rrHRQ/rXHN62ZypasH+dlT8OwWYTQ+CroqY0bLP69FbocXHv
GTOxxCXHTrelrDEy2TG8iH07h/fTQpY6vL1D0FZT4FjPm1Mr9Nnz6pRtIBaK
G+y4ppsJDtKC5POjOioXa8khf94HGkijMVoI4qe9DRuH0hwI9Lfe/ZJVkgvB
30podXMY1WrWyFUeY/G9yYvhThMN3iUbuXNsOAgOyEkW5q12UNuE4JtvFj0U
aoABk6XQxkoBCD5qEjmv8EB7iHHVZhkIPCPCyNPNQssn3vzNbCTJFOX7uzng
YyzXsVV/6hk19Mlz98RQ8MG/uZrgHLQwfRAELCxsvdrh2BvLhhaEnTp+q0qx
kqj2DX1TEkuWqfcljsYRvs9oCMxzJmY71gmSHB7z06mKCYn31MEziOcydImL
dc46YoUBr5bzOgJKgpEBbqbQJ79O8skfQ1SPmm8Aft5Mot4laEeVqOzHg7BF
QyUZ7iC+QLK6E9W+M+tmzvDklTe8LZqtMufrxlHBbgDDaWC9S3Yox+/cmerW
uvOUI+S2Ro3NN8tzLW8U4GNHClyhO4SVPEanHwqiCBZXwlVBGPs2H8l++K0l
QjlwlG/RCWUtfE5fkkIYhny2QFgrwKkeC7B9uNd1KFXH00njYaVmNLutK0km
2VLq6m0b63hmN5pwluSWGIg4inAB3RJKD5ECDZgER5F7matCgPRvEEY1PjNR
KgYt44HTM6J4fP97m6Qf3LJEkdQV1uJFzPLsLBzz5Qi+1OiLWsOXoXHYg+y+
UyFl2Dkdl8c7vI9EfbCUvhlFBbOQP/518ClP2krl9EMjbKx6A1YlrOOc97RL
NyGaQ+/NPwcwpbNViLUExBJk0CygaafPBE5cTbEjunc/QCbUTP3LodAfQLzT
p+9UP0HtUauir0+SWZ0V5LAtwoNciWQrjTarseYoajDodD0bXMym6x/NebKu
sed7ymSm6bfia35730xSJXf5T22OZ0faw/3M8J97r/Um9mJ+K5X595ma2qt8
XfxgpAy2rfWWH5iUpNo3E4q8+1WLVBwJzEc5przytFp5QiUBo7sgRPFqbn5k
TSSPPt3zLRO6WrN1XnxnUMqq9odd32mySr82CKvrVvd6XOuiSAc+WpuLBTX1
LxvkST0RvD2bej6WaP3ZzCLEIHhV/Z6dRffdfARSe4dna56Uk/8w4ngsLJxz
6KQNBPwrQJwQkfGj54lYdQjLoflC9fyHT+VDFyWsli/62JQ/ltU4a2zCr7fP
yPH4tv9JMRz7JFyXrWFMLKzdUUMi15SvibE9e57kgB1pAQnALYVDP5kIyAuS
lkA81V0FWZVu0HE7WlWG2KTcj2srXy5g+c+Hui1kmzQCRTTY3UR5gCzjUuLP
9g1sHORDjPDFLQI6EhmTv8VXFAmUDGhpkyiDC3juCCaJ2bKQ3FFBU7c+sSt5
o8hCmLa731gCscll7vkC/ZMOFPBwM/p9veE8UYD7prUBV6osD50lZvQBOYgw
H0JaDBGKtRX+gKTfyPXaTv3YMlziIj6Kf9p56YwX0k8qVCGV9RuOy2Sf1/BD
d69xfzRBBODGePdjDtHIsAh3wlayLwaMJNzw/meHok16hOpDUcw1itfDMmyp
q9Jxal7c2t4moBWrm3EebNmdGdzqdjP7/WvMDfRwUecn6lPmmYBPQm45Vx/s
XN1JgoryVpTY+UBIFJpgAsL9slBetNj863XClSGF7Z6klpqHFnB4xIDRpwvu
Lj7aiLhX+qdwKeQkIlOBOE4Wm+b6puGakWUa/MFwht8x4gsfmAwwMx980dQS
rFDb/Z2BRVmsOBw+26JFEPqvgXuOecM+ECsvOHrQntrK/M1pMFUtrXJmyFK2
yuVj+KNCb97ZiAkQkPidVlfeE22VyMYXH2Rj8fA1KcPDV6PPbehIKO+7AvaN
cW9oB1qAiFZU6JQ7yLuYk1jMfT2n544N0+joVV2dfFM/NUr6RyflIlrti/Fl
Ck5wfrQgf4fyUidr9FZ/Vg2Y4RmtvdrR5hFIjWphaK6zN7hF6Wg7GFGQXpZx
VjCFRBaBggmoFJ70/coJSLyo3XBbSs1wZxejskcBP8fQIWhHemze7nEiaaFk
Ud+tHeYcpefvrTqrk1BHhXl9ANjTZ0wRpo1yTEuRVEowS3rDjk27to9m5z9w
sRB0rV/uPTWPWIPo42pPMlfFa17M4HVUlRhKZ7a7RyVaNfHboTLp+P2O6i2t
HIpeWr1DEKAg0DMTAthVtAy/zEvpco90R49LmQouqwU97BtJW2ikdyxGbUMT
GSSSoPEeGGEIdykbGmoFbq7OUT2Nj9UmOqAJtn6YJWkMX7diazr3cGmiVKqh
evY6jLdgeSayy3LElo8/TIC4916gsWzIsmIF4RuNsPcwbfFTbDbqStBIuftn
CWx70IQLEQ39Dtg+6xphh6XEJB3hhCXax44I0Lj3/L1y8JqtPTs8nBqEHTL9
3ogIqcGma3tKhjGj7QkEAP+DjxMe8xRNtS4Wo47HBCRpPZCSJHEB6zPqcsS4
4VEAoA0jHiVaPI8gWZnmPzZyW/RzAO7cOEN9h7tP0Gb/zR74TOHC2DiYMFxL
Z5eYBROdSffgnwLE3IG4EzEAujPI1ePegkhtyAPGi8RSrFUKlUsF1dKutYv4
hb2+ic8IZakcqMIHTaiHiYyd2JFFeiKvJZLPhr2TSLvmUYNkZ0ISW0KjFu+u
xRv/AihQaTOHrwkXH+AiJwDWWjaviHfXPEckLK5Uogjn0Pb+yc5BHDVd0FSa
rRbn2mnOh2ktu3ifWycgJs3vYlq1lJHjQw8bS/dcZhGwhPdRUbNlE7B8hKCB
VE7QfxyfPPLSejZxjU9aIQVhUi3UfRc29l0Oc9jB/rpL3Yrgzqan5dU1rETi
h1JE5gtxf+6/a5UufrRDzYHyclv5Tg30K6GwpJLWkDGBrEkqppFcizHOcdZq
J4tEw1N3QEuxh3rvhJY15QX5Y9ja7qnYvnWdPlO+EPTgoihCKVUWqUo+DLOB
+IxvCEimLMVMKe5DrwYNVAZJOUZNHELm8Qw24At+h78/5AGrdFAbfgUwUPM9
kuddUu6cehlmB94orsK0y15nNzJ1wVKcH9nPHw7nazp0IY8MuqU9zD+l3blV
IQFW4qiwciNw8Nb/cf+xnP0wR9My6v8QJFlqRrxwrV7C0hOkGzAAou7VYwbk
Nnyuem+1AH1+WMCEWUVQmbRRXYGc/Cu7jyqmif0nt0Keu7tmzwo4XFoq19Tn
IBzuNBXS11QBlEmWQ5Kf0M+T9KlzmgtXno90zwdi0pxCtPpT7/4yGgv6JwWc
wTVX6Hruq+oYQo2xU6bHegpSdbE5ekAUS6xgr8okZZ0LOaChyxycoaZGGkn1
0UuZQNf8NkuaxIGwZCe2F7DExao3i2j4Ut0SvOZZPRLwxT3dnTkb0U1LvfIf
IOgfzV+oBi2CB9Zx4qj0nM+AG+KtaoVpYLn2fUGj4i7XLR8lgU04xDvYtb2+
dDNHo4idXkj7liHIkjdAtSYbpavmt3c66iUvMZhxsQSdEXGvur0DsoI+EqFt
ALu7Ivk/BN0LHZg8wo3sx1rEYdht75J6E2mSkowaXl3cjsZ9+R2c8S6SAClb
Q5Qy8NCypb3uT0z7tfasSdH/iwR/RnD7XksuMTY8NuV1feJaL/ia35cTLWYj
9DfAs3b4fvrtYLwU389QrUEafqX7r+vmO+2w7S2Iwjgxf+PLlFgwY8KYmA93
4Yh4M19qlLzjULC56rkOZkorQIqUtWaoE8g3R1uULvGNAaQ6mCRo1PdeNvnC
6IYeUu3gQ2vU47NHhKFnknlTbiX/ck/IvLf39mr5WRMnVViqnS5BZ8HF9BSf
8EORGX7Gwo+pCaQG3IKB9Bjl+03mcbB3c52agEwM04G+147z+R4K4BJD61TL
T7tMQT0v4BQ5FE1y2UZYLB98uaPEoGnklmYLv7r6d19U2aDHvR1VVUalyVfu
Z38kSmPsIBcN066xro24LNsP+d9c1KQMArSxKOa4Hwtw0wsq+tlQmDo9cFqW
atWL3p8rhm6OrghSBZ/PhkRSoYileYgyI95cx6wr6/zktEBzMcgP/bsSD0rI
TXsSNULchOwW2nRJbhr9lBYxf5e85BFcD5NTF7S7dOqlu1jzLM/aeXqE90On
6f+xalQ+uE8Us1sm69IiSihSZvTM2Cc2h2vcD2YfK9422H5cg/xp59JohKtD
lUxpg3f2tg+9FvbF++dC90M9e2e7PwontT0ymc92jYt2XyHa+axXHWHeSkpF
V1qwUmSqUWVPP68qhBa/4yA7cVu/hX27Q6Kiks8dOdl+LBEo7rHyG4Qe3I92
vKbWcMF/5cMB9NqfNUDLrypmigP4o7gI9DLOCcx1pjnZUA+nxcA2V0ccsd3+
joPJTkizAbVHgoT4NJ6YQFBgRC9tNDey1IjAEwSNHbhHPbE7KNdI2qSi7JZn
HesVOM99tX/PnS/e/reV4NgVg9gbcfYP4TPnD2i+mO4mPleIdMzvn/EgTzeN
9TeHh4zRtFDYx5VXO3SaLrSo9J5sark2AtjCUUz91Jn22s6D0br8JpRMARDF
F2Y0zNvKeEFWlt5jgxA2XZuAXP4BFU1U6J7/7DmvQjisUvC1R8vdwIOgno4P
IHxuJbjdiz/dIoEfj70OBkTk8Fud9zz4wI5XdlEQIkk4GEZjG1V42PblRLSy
86ldNJEiW9XXyhVR11Pmyl8cj9N4xNa/jfsXRSBRKn18wbjU3HpPuLsFzNsm
HkUqQnhx2SoIUzRwRJv6iM6QVgWCtj8t/bcEy33r33YW+Q/72cktcTkzm+X9
MySwQXH6vTorq2EFOhqs8FY5W4ybsU4Wd3BOLP6seySsdd/vG1saGSSjdLe2
1VZktIhzrSfMGHS76He4nQmC+ORnXtcPILypjLDsNubEZ46gE1Aoke1L76il
zKjxW+U9sulC41wVoZ5ZwbcAJSemjQgkG38hBGgdfe/ojH0/j2rXUHZLGCfr
CpwdWjxNPaBrSAv3ujAZjHGRy2pxMR1+11MsjeZC8OqnuCmQFYAqT/fjYQAy
F9eVnCQ9vvtFWCSB3v91jbo5HqrD7PRzXtJM/yjCimPshIMRq3ev4sw3oGwW
kBGkYOpWB/XzJhytxCNFdMTd76FRg5lofJlZBexmGI3kXplxWGeGY6NUZ76w
viKJfglEmAD1NCT2vGJUoZFnrXCG202guwkoCaqhom/AOyhHiNY4QHHYY6rY
DaeUmTvpigyvq1DS9h17KDUzMCyJrnU6YvZPxJ44GPaugVb/6yVcPBS4hheb
/DQFS/9WrKVRrBTJDeWcRtG/PRT3QJG44Xl9SHLmdToV00eorMsiLjANxMVW
GNFW4fuTVp6pf+agNhH5itDOgVoHM+FZ62zBFsKn4p5vxJ+3dLtu4M0fuRLy
u3d+ud97TXH/IHvfTisPG/dZ3MkbJwFAxGfBZ5cY3vFWn/O+4ZvUyE/DiJ+I
+IN8MLBq13WHKsl7LDIavNxwzfZQ7DtlJX3uQ3avnYm9LvTbRWQ7Syc7L8yW
t7MqddzHstHgAHAd8lps3KOm9N4A5vXKp4TjCGX78/NHDa9NA47+zGh2KpwC
1SH/ZVok/jFe/eKW2Y3EdYKnWNRyDwlfoF/LsjS4KMPfYDbGN/b0Q1RnyQ/j
qrNXXLoiQvo9TxkoL54XhvajFUlG+w+DdhV/ZLlB/9FuxioKZL60yZW3O+q/
WHRZnfhd3OTsGanQ2h7k0SEeCy/pTT6DFc0xfIYJPMdLQZnt+RxAICIlbBEz
KwXhei7IPyaHeUzLhBlC+SASRazGBoip0tCjWN7s4A5FFggRR5f6GIU47B0X
yFQOVwnzVjqEIVWUfKi2KnfxTrZK8XMUGF2K+WPvk5+YSFUqs4o4PdQ/6Nty
VGYoDG+jNXzYbZVY6I1gyGgDw/CtaXjzgdoEam2znCx1cHlhIkIm2tvdk9xi
gbaBufEzNXB4oYJ9PI9q1q8i7b2Rur1BirmBcBoxoXZ8ZEcuch/2FBVHSLXL
kBV+4zxO3zD7CNA0NuPQNxvSGKSoYDmxwdvCgxwp8bZhAEoQPKSC4mrlgcny
mf+5kROo0F0cWvwlM8FUPcBiXWVrQTsPXcOeEg8qQKQMoow38IyV4K0nblS3
2oT7ELuCFHCE+iHMK90D5ofTWHCyDLXkE1Bv8nvzVrmsvkgACUXwA7niXU6W
bWs64ZuMi+QAoTAmxLgJ2pk3e3n29bT2xwdwdRC5s32Oy9mpvdEBlR0+ANl4
i1ek24pgb93b3qfKnG/r+zB8CkUTZ5C8sSpiSzFOKK15mLfhDhjG5S/H5Y9f
m1uO2N+deyZPqAYd915SGgfU7e2CSh3BpDgU04c1sCc+HSN3aTd9c8MWe/tM
kOrsgpkf2Oh+7txtiURbYcZuA9f9hivXTYGnqXIlOlDY3HZA1WZ/mXNdXrP1
9Ezo73VutXb/84/9NoujDYe2HDNg9f6ohj6cGSSiV1PsYHQNlS81RWjgh+uG
WOg20zkeeOQ6EfplAnEwMpbUCwYAGGA40Dy2mTQFdVVB2irzRCL7WOwF70kn
UO+DwskNiPHICJOq4g3mlXQetcRlh9bFaVtfu01OUMftQduoVuVu6y1J0/WT
A+G3MB1BpdLp+owAg+ShZMz+uwAYMVv0iLk4aPueM9b1k8YHH51nMnglCcEl
PuowNKgMtVVtzHxKKXg3pwUvyUQNfIHhukACC+LqfHEkOh0FoJJDSIP58uNq
6JQRVIcZ7xFsqd+4xv+uZNrtf3IH/04wgyLZgm4OwUNtSKUzJPdruY1noU5h
CdqShQL8Q79onXMm+VQxgJXZSlgh+Q+x1mW4jRBI4dZ35hNNLiPmjIkxj581
9dbo0MzVzebhtGV4Ygr/0rnrQKIR1kfx+s+Ks+I3fFtb8f/bSF2Xnsx6kbhB
E39UiPkdfAjFZ4AVb9sHsQOJn2gZlpHcuLZJZwtrmoqvqrmUZ0RS691tzk4S
pmPAI/tYO5VBGOnQs1ihidzGtTlB6hZpbdpsyujUINJQbPQwaJX28bV2g7UK
EbE3IrLq77G4mKJwFUp65ykRzyiuDv8OGdZmgylvXRGoJJ38v3lY81uFDvM+
rtat4jLnYGC1GSoLK7hedyyIrYEm5MeocgUyt6F63K6lZ4EVFP4nkCoLedmi
hDXG+k9FfkduSR8rvmNPJDTSHGPUjv+tnbIGHY8SkZ5XZCpyK26+8tE8QFX+
yAIBAYVv/PrA2Vyb8lcOuV7nsRbLzd64H4t9AXMDqhETIe39Ufq8/iAMXI8k
Ity782WgR7un5lsit56ZYd1nY/kPqeHr67dmpOzUJhOfFfompI2LbJ5iJPKh
tHsuTC/GfRrarGCytg7z+Pn6qTazHil0rmwzejCNeJtTtO7AfYic+m9e37Ng
gN8fzyPSlsMofMMW5jCAKNoHX4sNJc2WqMQReqeTi2ziJFjYabXeHwLPtuQn
3eyt6iQ4n4GSjNDnhsa815BtF9gRgO+rCViyqzr3ZhvgkAfFC3ykwqvqRrB+
8C6LABbQo/0XQcvcExktjGztGoPSTGDhQQ1kCeVd98G8eQcpehLsRiYApxut
4R9ldmj6euHZR0t6ikUhIfrGCW1sDwQLK12n/PrdHlhgIErJ/lwXR0AMqssK
jaI2DAY2IcHpexIAiQkxrU+y+5uZhVEAdHQ235SoQ2sZvMFZNO/5iL72Kh76
eDQDbWHyQVoSdC00Jcig9xdEu4kz9vIoxo+cQN9tXUC2IMeum4Sp1GroCGWP
Vw1nTBp+AJIsuF262GFE6wcSOKIsgefYtgNf8rKGXlggf/05PBq7BnJdg8lo
f2MbVavesQUxd8+e8MPmdDhHYNrN52uPPSYDnLrPU0vHkIRFFLcdd9jlTEbf
aLNTY4okXwQ2Zi18gFLlMN0iw+LMfaf4EICnn6gZti6gEA1mxCvZ8oZQzYQv
1wVUR+MPUIkUPHi/HtULCCtGChO4Q068PROU6qTFKUjbti5Wi/KPTP2TfBw/
CDxf0lYIruau+Gty+9Ig/MLXtH1qJnZnznX46AGCobR8T/Os9qI3lq+R/Ir3
4o0icF5ajR40JA3wqM/u61boIdDckI3yrGs8EelFn5UQfwqNRRrqL7h8rSXg
2lSZqFHhFuwiq/Hqqur6lIBl6CFLHwzC5FvqMrs9LEiuVpsAZxjUF/rmJVpF
lH9whh+WCwXVfZieCkbxQJbTG6djOEKt/UpGhb0biTqBEq+xISX0ZrJU/VSl
BJ49Yqjtf97Gy594UOThS8WW8HLKnvtHx5/5MYAAvS52KJc+TWYqpY77oGaW
gNHdiDfA0j1U1LNEbibLaZoYWPdkuwYdVPvuzkRLtQ6qZ+2t2qeprH3VxoA8
lXR1Yf8I+XLMzrEF9iUKUpjuynQb+/PawiTkgAOkHE4sHDH+ROqJAO2RboF2
yOXZs8nD5cApMmNexW8Kq3iy9t8uwn/djPdUgTd7EL4UgTUJ3N9VSeDli3L/
j3zDnIGhLQ5BV5PHSDEGeN2YlJ487xK/9D5NJeJ8DVrsq69639xfuwJujaZz
ue3M0jLuLjyEjMoR0oMU825yzxQ+6SBa5KKZVfrv7sEfK+rDZhi7mOa2eEzl
8e93qS8hSLATkYShTJ+gAg2H/OsLENJ5k12h/ftnDs94Rhgkts3J8WY/27uV
pwelmef8T8inaxY4FGccsKgEWDc6HagNmThLkdajgcJ4uQIN1DNJduek/Y/q
MWJSjA8ycxDXFlYfV7yAe5NV5EaVdfUW9pTqEvhWoaLKThyI3Vz9KKroMJjm
vik52o7ATIyql+aKxESQRtdj8NMISIKl6GsgHcTqoyNodfpcR4dZdFy6hgM6
jKTPdFim/8Vxz/EZHc1ZuxK8CUrmunOMPU5Z8fKVfDv+Xy2z1MXzRfgb2E8L
vIN20bw5G3G4rZVQFxuPVGncQa+ZWtcqW8ZGulmmNiLPr5fiMzdC4jRgtbb/
Ua8BJtqIibbJsQS8j00oRiDV9fC6CFSnlqT8jmS4TW0IaedkvHW5tvPpo5ot
N9SE/21iE0J/g8lk/z7Fjd4QlBiu2nXDQUsxevUDr0/tLDv640ZSh+gXcbdU
Jrw6DKFr6VIOuX+HOXWQssygvvSQFGkQW/qU2SBM0r8a4VXjjWEAC6dyuH4b
maTWq2q+NpaYZKGtzl1ndZd1oFVKPWkQceQdOA+/KJZ7ZW8s5scJJbyQvz3p
IcHMPLdx98tdGfsIQ4cRq6Eh09dnOfazYdAO/tdzVTBjPnOZ2rpU0dRkUiDm
RqcDSmcm8ZglL/RAQHonURI/Fg3S9GNCWB4rBEqgUg39PGphht+ah2zdGhy3
6N2F7gBYIIdeQB7Oi39pn80NMKWMiVdlc+nxVwNX817heaat5RniAtALISvr
Co/97MNSk8VCHW6elV9FlIGUJXg4Iz8F+EehuR9uER84+y5Lu60xvJ6lS1kp
ZwcVt+Vn3LFeIO9NxmIFMm8laW+nxLp8sceQR5tGj7phcfc3+/rjg3/PO4Gn
/RvbjxbDFSmawnzmWLBIl+G6t1crHJlyxzH83yAcXuzja8tgyNSUw64baHxi
+aJKK0xMwTf3bxpKD2ootdDBxDgESN6Zsu1zlPNy9aimM1bM8rbdH/ccWBrF
QAaBoWpm0BlbaWdQ0kA5P7PzYM7a/qcraLTJWRsb5ct3ED/a/5QNPdcLaTN2
VWKrkGYzWEfNmOEsFVfY2Es1QhjHrJLxFwDgrm4JU29hT7sMTGUWKbi1WH7v
dnlz/QQhKZEZcqZ82FVndBnmGuZaL8hOfSTXr6RfWIc67hG33mO/kUKHJI81
iwAlaWayBdLwp4ELXzWtJd5iNwG6Kj8eVSM2zal356qZpyy+DqIsl4pnuALp
FQzlKq2l2XxsKHSabtgjFYfHVYf7JRPjprlVTtpynXnT7lPs/7D1uAXUIW8+
JxMpTX5Gip8D4ibF9MqEM6+KiRUNV69a5SSwk3buLykDOAHY70eFCVCuDsjF
cTN8E9HXhiAEi3SIi25YJtqohcnx/aenAyalOpSsD00fP320nRpx5s1lvR8q
IR7FhgODiNNLot50aEU336ZSeMiZS/VRvDeOHL/oGQqiaa6p7scKgd9gDG0w
yfoq1cjBrM1DJZe+vvdbGTtq01NGpr08qjixtET/il6r0Rqp9bHQIOwdjSmx
3JG7pcxvdjOg8AD+cnD1UY6mbY25Yxbfqvemkb5+Gr5hzEy5YswLuDaHbVRA
B6yYA2H03iGluDlneehEvKY6UaMgHPl+x04lYW5RdRgqBW1CeCk26seva5/k
KGYb0pr2Ww7epak3CM4eHwuXk4k5/XB4GZVX9a+jdN0cKpSM0X2WUfbBhHbE
8gL7c33zPoZF/tmtpbrOFXbChHtL82xK2XyoBPenuIvz6GmQPqqQjmBX7m3y
+f1mCQPXDLzA6ahKGq0+qRfoO4FtZho37mRJfLcam5blWj7nwQklGsg6RkXe
gkFOYlWcT8MhJcL7tP6Sl703bLI/NccNRKOGhuvFjQJ+iVyu09TFzlZKeCrm
zYHzV1JO4rlEc7MYYa9QitUnWN6b08DDuJu4C8nHRPWFEpu2rDIOxTWUwMb9
jA0Lnv4zjycr6yl3SR+igFXtRucrkOC4gPBq82lrtiRM8ua/z9zsEdL97SOa
o4fY3gDdd8XjhJEG5sEK09D7WiMDJwIoJCWxa3EJBRRwe58qdSgGWk9rR4h4
6fVvKCxAjjHm6ujs7eAAdtGAM3fLmufPkyYdNz5g6vm+gT5oneQRNufWjByE
1IFsDUoV17WgSU0Q9m0Lk/tFy4pHBEw17NiisBf0QpfHcPiL9kQni70aAGAN
VH02Y3WwWF4d1VfuZtVObEsOb2GaoTIt4bNyBWunGM37aUoVoSMQaciSY6sa
y1J6C7lHN55pWrF4TIGSUivVOCkrLnfOsjdDnCVDNFU/dVI696+bQb+EZX+8
Upy6dOrTN/o4VVQIWMWn/ssVHGry2siPr6vwA2lJwuxFAHdbQ+T/ZbcW83nY
IZDGKkxBSVpxri3jDRqHuzP46FA3bWwad6mdQRxaRkQQ+LG4DdsYdHhSJKzC
dEQ/iSIhTPWRHime3sMex3irM7fFY8wQDWow/hIZov69W9osEgzPH+prOr1i
aMurweXdapgImR5GYSSYACtNyeInKVR0PYilA9jiYkK9bjNx0wO7rydJf3zw
biXoGMb6FRlEW7ogWgrrOTQEVeiXnwnZsxhkV+18hNJrfHL7sh3r+BqNVf4B
tkOh39/Q3+YmPZrzwJo0b/0ZeJ9ljwwiJhkTyMcOPlcRCMU6FfVg6EsUMY8M
9Iigf0Hv2SQ3/OGC9XwgVmxlvGK+2q486HwkqegTeVRqqQT9p3v5np/xGytQ
kT+X0QeREzvQx93uwi/g0eK5JtmGJqdDihO2dOBg3g0nOg3+PA48m1SH5VF8
bx1I0bFSl5l/Ovoyj/vT+dJ1QMxpsyXIQROz2bDkB0olAcQYWgDw03WI9/WY
WptJfS5RqCcQh+795SJN/pEvXmm0fdzFo7pnOZmvWz2pVqk89FDzVwLmuU+g
BQzkwFife2d1r9aPNJFrwBBgrD2tb7n7h0epKzuMbx/vWn2ePTdcgrclc0Xe
pjE5wg84x+FvKy/To2uCGgp7Ut/i9MQC91aac8Cff/aHk3Ays4NEjF31z8Xk
C1LqrZVL+PZaL/acQ5Qo5sgLCJU0IUsacMjAH6hw0CKNm97I6GGjSB6LLKqj
pantVtfrSyqXW8+YklhykenkegOnpT8SnkGe8JbsQoXTh8b+MtM04W7EMdJf
uMG0wd7z88AqWDNYUIU0AEeIG9ICyn0i0GBEIHXsUpCJrA2IxBDtYayJbKib
+eVj0DV6yeUdtmsNIbS4qN1tUTdZrq7oqc1kKkcRfljPcrbPMhChgWeTEH5C
G2VGOmlTXviJwynHOa4SmpOjsl7Dd1fSwzy1zSOZjFEAzPODC61zi6Mr4v7H
bnWF9T3oaY2AuU/GigIDZFpfz6cxf+CENcEca4hMToC0Kujivh/y9c7Qp14V
daahtsPy283dCXvBfhcgLX93kItlFfBIphfb9trOCkC+DRieYf3dDocFVuBG
S9G/0jkqS9hlcc6BEig7Ua0+zX4WnXak39kJN5ksBG5KpTSRGww2DWWIEWmc
+Wlakwf1wRBUApsMyoNwnvMA4yeD1vo2kTUb+zINa1e0eQJcO5tixeHqr60S
tzHqhDYXgYwECWfp3ysTTuGL2okKRo//OvdhBL9/AF04ltuTaT7/BoZ9zcTC
S71jKy5BVTp1Ue8Z09JT3Ad8Elh/toZdO86X6IAdbLwvuitMti+XwB7p1Hw7
O0ZwayLMf5FldYcki8giVwbNtBwXbTGOm/jV/aUkS1m7PNxDQ9ArA6dlea0M
RDvMT28mSeP0CeTHzvYiWDlmKn4ezayvQ6jTxOrEr4H0d/BGyU9kcw3A2q2D
qu4ZvGC7Y1RlRgMrOGAoUMWlBfR19ua0Ejq1Fu31CW+OGXFyVT5/IdYwiB8C
kUS+Vzyas3qmd6UNBi6DPbC7d/FSu70KIK1PILMr6s5JRHlODS1PBGDz8Hpu
81JtnZKYRbNea2+Uf3p7g4+Kwkyyt5lY/Hf1rBmlarS3j1d/JhVeUJ6s1SFT
qgxQvMpfy2uTky/P/W3wPPQVc9kjIOLRTBZrLH/OacxHMe+5HjY1gekYaTct
BIuvyx9qymdW7k5ucLUcs/wVFeNSY3o1yrbYqNZFL6l6RTdgeIvtmXA0bDk6
rnSq8xG0zUy2S8PoyNd2fQfPcuApZIDRqG1rN6s5IO5hL85OAqPjOxPscfqy
/jSme5Ebv5asp4pF6HaxbqV0TT9N+aPwdPcUMX36uqQSqwAozGPijgBnD7CR
GAem1M2rS5LnbEte9JROkOsVQ2hH28+8KY1nZ4OMLL4vIkbqWxvNqGmzGH8q
rOj2de5m0QNW6N/f21x1U4Js7dQTz5PFXlT7pzHo/wVs/708LREc9je0LPJz
ng0iA4qNuF8XF+bnDCkaN4cXvLVVT5NhGfP1gN1Gb9zmDLULHK5CANITzktJ
R2IA3ZGJiF1UB5OlpIafPLCJF/3h/y5dS2Y8Q8cGMhkWMNkzgrwaRv/5Bz2a
Efc756yz+sKz2QzWBsRLKJtsjj+O5zpBzkLOOU3ylHrYj3DXbLlYTqSZumgV
J6JJ8ZWbFGUcE3ySYM/4R1Uy8M5XuD+Pz2ki1UuZ5/phCcZVF0w5/+kHDNF7
1AoFE2nF4J52/usSxJdtJO0+LWlwQifcsyVJZ9AFrVZuZscs1TpkHJcLSIwH
JiZTJo020CjgLaFDqxmbWjMA79Q6jf4SHFTWAhXiQQhQc4MReBPP7UHwJ7YW
8hjFGSLdIicTMGeydSrhkH7jt7ufiDzLLMWzCrYlHKZfc2ViDmZIo7Ats1bZ
UsE8IfPXXhg2kfSo6z5MQEgklf+2AjXia1kcSttO15L/K+Tc5ub3fMB8oZ25
H4C4Hn8uKrhpTIka3l9fnnjWMyK9cvV4K/QaNiY0e9ctRC1kStOIcrWrEf0P
l5wPARJliIxZpXy9yPbdImqKxWst8raeDfIn+S1uSJ5ygso3VvdpWqoICOZm
t3VPXt/xOPqwTQ7gJZM/9IkR5W2TrevocmgCOqNkSi4hMnC8CrsrvlornDth
kZ5bVvaeLJK7jCWQvWnZKwIYAwswuh1Fq6fecwL5p/ELknP5/J/mLVL+MLbO
LBVzB4V7VuYANYNfN/SWq0ETcxenZyPGlK2W9vRGZLXkjnvQYHiEIvZIN1y0
xpz3oS3pOzNbFMiua6vW+sc6DWZtjIfAXrm4wDi4ChTNi31u2LOXGgTfle8l
HkCi1Elq2i1qS1kuszrrwipaYUqwVbAHD+cCaGbKuCHybHrI2QLZvVgNtw5w
YIIroleMMqQ3FtJNsnadgramLlsvAeSp+lyEY2OXloIIv6cwrGhc9zfPAqBs
BQistei/pnfMDLLHguh4FpdGuoux630hUccBaoxurKPmfSJKnktOpO0an80K
kIbjXwrTqdIN4+eo+TwLX3cK5rr35LKPXr1jbekc2Gc8qMv5PM3Y5sjlZjsR
efRWK5088EWlm7rykTPWqwuC/Cle0v5demGuQgPpFLj1owMF7YLDBMm163ha
1fK9qwGsZGj7UWY+JUEjDkkBFIyObdAJ3gLZ/B6qGtisDttcIutSwmX4tHXY
L+37bWBTTfBRiRF8o0yoKcBrGvZX3pYUVWLXXsbN3PRjksAtLqrWNSnHmsug
XVpbJQ+VaDZ5VuZe+rYlU70aQgcurQNlY0lzt733BajIScGf4zB9889adXLm
Z1AsgnZPinaA4AujZymnmmXkGld7+CVUrUGqWNQMgxvjYysJzCpX5HVFnxZ8
3T9jbsdGMs/HaReexfmAHfGI+Makw0j7AA/M7OEx7/eFLea1681qcYzVY/mX
Qr4CnLq27QFIuSx9s7676zvOoMACl58nM6R/TfKUvWRhUVvvZgm97AvEoVdc
ClVmou30eAhjJ00FDoewntOpmFEuTBOGUaX6wijJGdldaUhrNstOGw2qiE+m
rWMaj5lOFM5FTe//TUJXd2/JYtM2IKqeKvofbuNYS+3wFRh4zeLjYv9eyR67
mlyfiFxxyBAJ+nLEth9VveNaOFCXb25R9nqpFM6sUgaqbp60kWCrtheourLe
bH4VtkWF6ravUhVvr1x5ymkFdJAfdVWpcaRbzaN2gjtriN9Hmq60I9Moe4dW
tDSsxTzRms/bmjsGGFZoIgezhhe+ZtSutqWpUdgnfrl8hIiWgri+KcmNJ+qO
j0MixOj0Hm43EcJ+oYBuayhfr5k2eKy1Vf5+IVz8g5ECi//ttHmmbd+IZUDI
pOeAq4IyncYzXAVnuSDzqlsOViqQoLyPDOAlLSG2c10+xB9dg/+JXDMfkSNh
dvmABETH4LDqwrx+oFAIzuDEmDwYMaTQZ+THJHg+w+m/DmI7Cnt65pCNekXs
LSWjPhiD2o2WwuhvEV9aArCU/ga+IzoauQHtwgUPG5wARtB96ae19wJNtHmL
gWjnOwKni6By6f2qu6sU+Z76QzUs3/95E2QfrIT9R7NM7imgrZ7rwEhp9uIg
I34aFcQxqYQOEIQ/GRRLpGUsAIm3h1bsv+wrDfEA9hxsoYe4ESV0zTbmCxBn
hspKPlrOAhjrbRSbvqC6MJZkj5jcxT+e0rqmNPx62KOPSLMMbnAflHUAw9Bl
uFr01dZQ1w2ETatqQvWXlq5/MadReeEGnfsrGbqixNXKSIZMQIm/VNX+ErPl
M94imtqQ+6/aGvt3kt1YFiWref67qKORjZnwcHVWmLIDDYHQejNS+bi4Zeze
EjZ7aHjrJ5jdp8iq+creeaGF1GN9neMPWpMsJe970/wabYuuYCYs2XSUJU8l
o2IML28EdHhTs6pMX5pe54GWK7oUA9AcppnfU2Ztzpgi1KwVNblqcm4yLQK+
ruzihWfSUBCArsH02s8/6X1DG7rdUJy/pAunZKptcIAm11JVkYLv+LF83prZ
Qlcyi3Ey5NNWXRH9olzCsRXVUCoFM7uaWzu1cBzn94nM/TgZZK1S3sAtGCTO
P7IQJy3fccHqiYa5r7fY5aBUmdzXYchjRus9HD5ttm5ca72pMK8TF/6EI1l9
0IhzaKJjP1ZoDmE4/fywPACYUYyouTgDKfQmfDC0IxZDjbxn15FvIns8Y/7a
HRN92sxxVvAXKXqvv/TfVOawEysWcTwyyCzVYpw+UfLim8aF57y0D/GNnLMY
SK0s+dKwJXfem7MrYQUNKfjA+yJhrzgfV3iwHoMDg7TF8mp9qhpTEMEqZkmW
ER+dzfmAgTbJexj6qqtFUFefcaMDq3N6fPLb+O7fQ9SBXqImQq1P0JGrtrY+
dBwgDo7GIKhindtvEE8fEAei9a1BhmzLhVDYpMN3AKd70VHoRCEbW4OlFMuC
w4IHabFZZK3XuXGLe2fgff0HFEWPajVHCqykTM/huLPvQNLyQdAPUo8oyENw
GYNL5lxT1oqDeIERDrGckfj5+Jwly7v1AN7AOF67fPXBzdaJFz1UD/xwkH0/
jAMp5pAaEL4Xuzzs27LVJq6M5UvShz5J3D4lTD9EtAUNyRwnR8+hKMKFutDX
euLWk1YN+feARXlLZe5bJ8gHvI3Xzy2pdKABSb4rf5NW81dOVIh6PaIRcGlM
jxDW26UjUyqU7I0VHo7QNdOijPZ5AWiZHFFujvuq2adhv0Slj3qyFRfpYL4h
WophrYKvGooBeWubZt113ywG5h2BJS7g6v6lZkZoU7SH1vNmBNUaAzsUmnOX
Zr9/J7uPf8Os+lTqNIzrpKzkgHlkdHdKPn0xD+uKRVVOM0OYSqA/76AG7xp/
32uMZQPAsWYzCIS1/sfVmiXvOT1ELA4TNnIdg4n2cKxh/odCIwLizNEy8dHk
RF6xnlQvhUWEYnecdTrE75Bg2xKXiRCfvOn4p5c2nDAMmJEKoHqJJa0kwCzX
M1JZfdqbS8Tr3u59SHZdwaOYoqxCEjAfg4qxhisyUPoGtLaLySCLE8nAZPLN
lCif+7yhSFiSfEaE2WW2Z/N1NgMIVm9c7b4Z5VYD9k/ho3Lge+JEnPNgMgqg
iIGR1GQd8nPl26hcCS1TbObC5K1pR51gbsV7xiPJ77N7/3XxIe3GRBgKfZ0n
088XmJVEuN7sEUbpJ5E8Uy7mzkbsS6v3X4rhKDA53L5ngck8VrwUeheGtbuP
TcmQ8eNq4HSiP6VDAL++h2lYhu7ApY5kxmIQ9lnGIlzbrTCEs9Tubq+lzMJC
ywL7KKa3knzQRZMIeCTepI7ctEvWYxL95UApJwHFJV7FHVzdOjNaX2GjaxXh
0jWZNpW9p6aFYuIfIVU8LeuIgzM9emOyHJvcj+xFTtM04A7ZNe3fhUd6kC3p
k8fkEDQ3gnRWR0kJU0/FTXkm+sZrhwFHgwV2BAA9rt0wigHJaP0vXBERCieK
tbl4Vbubd7JpBOsWlkIQ1TtHUUFU+hlEt9jFe17Q79c6rKPv/Cwdhwk9Ta/d
PMjRUkvqjhxT8X93AjHGfhJsf47XXpY85ij7ITkbr66x8ldcXwvjm9Ssj8oV
n5QOxJ342dEQJ21nwXRbbTBIvZNBlgh0/RLND2PHwJj90d3QpB1TktnYOcyM
xRZ38C/HOHbo6/eIkjWzvB0yPTpApKBWelCTWujFkthDXRtDQhnaDXoCpnQg
Kh6cY17wOUnIpBv72SvBN7GBATYuArtZezeKuf4n66mDbRyYMP4zfFORSdmA
KVw3bk092kH6kwXDviXKO8MAblqvppXWUzBfH69XAbXdcZ/3vUfMlHSi7zYM
Ssmj5Rvo99GjoqjBwfKOwqo4r0CWz9yBaav/GuFgf7CAE6vvKlbmseo1Rihm
QmKlBG9U51C6ZeFoSl40VnW/fSLIkdewDk86HneYYxFwS9xHWsClsDsf0Dpb
Khwp2vKeTXTbRitRA6ZJCMsi4gMWwbxzAMHXbNXQvoqC2YbJ6OGgON7Gid5T
w6bzBuYkVHDkjK+ocCHyJ1CXqqiZzdbZvACLjFrnxyYkYndw8QBnh2GRG1wg
cDF3SfM6amWstMUcDF9bsltfzJWaGdpqoymA9bDS+GGt5sZdxDgpFsi+VZgO
hRO+ZsxdJtPwp2j3FVyvacL1cnXQ60A8lafpoiZPR6Xvmj1Ar8Km92nypVLB
Xe/Evt8rf//+WJhhJwD+6XcqL5fJhB1NgNA/kIqYUSw3yEjtAUsf9FFh9zk+
+uiz2GQ/9ANdLQS7ZalY+D5hPGk0Wriyq71CeXPSaWa4/5xIUDjAUBiswkE5
v57faGzhBRbqYk8kSvDB2iN8R9akancdDKR8bSUFYYiGUxT/imXjwLzQU5K9
/Eq3QaCZZ+0zxB4+DegQbZkSWZ4zfDRx0kF3vE3p6aG+kG18xqFJJttuXExI
rqwdHn0NGnUDhZYd8X4jmR7K38J2ADY+Y0mIgy1DjDtaih6rsU7r4DPH/cRh
iI+4FjSYs1dXTv5i0dUFF45g2Rh4aAIv2zeC85CnyAfmi+xfv1RNCpJsrwhT
mF9gNHtxfZHLbY7P32QAA5F2ZQ8ciVjcQQQnQJIJw1ooftZ1+TEIw5y09btf
iITHuohRzJqJHTiVWRTgcT+PbRYs3PacGbvYOeNhg49bqXDl+WbussgkVXZO
LzW9/5RUdCKWRC5v23tOJcudz3SWKJ7irQebZuw0nbIQdRiJnPhS7OMqdOL9
vvoW+zPEGFQwh+fOMGkw1HSWrzDsr2UDYzVWV/fZsWWXl7woJA0txxRxIrcV
0AhyHYwv8WCXz8bUy/xiD8DtJh1BuuGDEOi3cnueN94VGa5a9BDq2hcKLLkA
+0ut0QK+pmDy87/GJW4F6gsxzSP86zdbd3W6ysSAr6hmiiGpqBfoLS1T4kJs
9fI0EUxrXVmn2r8GdfzH8ie78isn1IyGzeJk5pdknSHlV1fMDBxBOkbvr7Ps
rZIRz+p31XUOOTw1pHoJCt5Map2YMOFW4zhTuhUxg+uUMVj/iRL/9PAk0n4d
bMYGdDusBDVBzb0bTEC3kxfZDHsmvLALUKCT03az7KiNIJgFgm2vGRPhdcTn
5h5z/xU4wFky0og2RBiDnFxcO8hgMlh2LDcTBJMvQZ+MUztQrv6U5Fbe1bqy
KR9rsPKQjr5X4FeF21QCXWtKSSW5DGQ9+MdRmsVmbLOkvR/JBifPTyRPPuli
clb+c1BD6Ht0LfK1XHNi/zM2TuEzt3EToRnZY9oSFlFN1mwi5XZuEzb24ZEO
CFFrN2FZckH804cTMR/W/fzYoavdoCo102IeqgQD5+zy7+AvSHYlF34JCiPS
f1dI1cveOA3RWQIXx4rHzHJODzDuTpwPc3He9TE5rUaI/DOJwr5GJPV+3eWo
aagSGPviY69g4XWPPkkUCNVLHoYz+e/tMDUIcGjfwb8RN546GrmJMWT4xVI4
TwSoC+u9iH3OYh7T0QAVwt/ig97CN32C88OXHHCRGcrXpMboxR4r4Yxv3iSn
zxtNrNqFRxJGIYJmXeYo0gpweamOIJn08QorvKwvwgYLxY4eZ6UL9QhwLz0E
+gnX9TN8WeIjYInrhKkwQG9cqqNlSDAi26EsRKCfIc+TZRTfrR0KB/IdDplQ
iaPiBzguw2a0rJvcnEV9EwTmVBs2kiOI6vN+eSdqrC/dRIIHNZ3OA7N/Gmix
zth7Da2J+TRncaSxX2OpCQXyjQX0jwptBJ/8Y/k4TGPJGVqTt4DuduX7dHEv
QnDV3I00sBkRVVhpnjHNytItp49xg8en2byYgXwUE9toJoXh+sAB5ZkzRwWl
6SG+l+MEyzgC4TezqAozWxYiCkWhPTUH34ezDf5crWQ9OBCOwcJS3+Zm7Av6
E9XFNT+OyDnzAInHEdG43SLwkNO1lrTxseND+AIKFNnNVQAOc4pfqXDRc6/9
e6uPuA3SvEhKrvdoVt/0fZyGk9aP2+UkR6tcmaJCbuFXxsm+sg0ULUL4wlat
m8fAqLMSoZeti/UL7WtxE+REndVToijDVIbrDmHKD7K1hh7aUUsHEC38CXrM
dgX4haw+b1canB0xuiFaD8LaC/YkcAILF/XFRMl6gBK66zb7snDV83dS5l7W
ufPAFLRgRVJcs/3g9wzxvr3lucfya2HTV8fZKBpjCrJiLbDE4s00d6QLqkwU
4nL482Yx8NslH3Pe+977f1Y64S9gL3LdmCJAjlEbQwQiJL/iGKlNQIrbsYfp
ctGF8WLmI3BuX+VN+KaECDQAGUf9nHwfAW07B6E+Qtbe+ZleG+4T0woLK1iL
bA0qEKM8y80vgl/VcrQXQlUqy3me1QBE9+4ToG5zgCruGojJYLQMNIzLrCdN
WTDPo3ZV5r7bP16X5FL3c3a0yhnG5CszSlA8I1W1m3ZoRWi6lioelUseaFUv
3Ypw81hIVTngyKYkx+OU1Gn4hbdINJO97ouWVECgX41dYQI3aPdn/2dwNBlb
4R6mKlgmtYIQFr7GPOsX5jQGE2luHNBxulMTcG8UFzXOTlo2pjGVxZmjztI0
kuqFJFhC7CWrEzdsvPqQZZGtsfr/lnRVZ+oK5mcF72qyDuCKqxsHCW5f+2BU
9fffWYrOenUbMAs4CHS5UivN6s4y5CZVjx6oHpK7BA0TvaOJbaI3r3abTYy6
2dewk2+JD4KPg3Nsy3KQ37Fe6Hz91n38jVOThPwBivkqxp/KkgEnI6etxwcu
ZCx4k5W/jYgsTLkCXQEN9NUxifBNb1mEnGADxDBfVvAydk/fzHIa9zLzycLE
pCIhEHNebe4BqFCVrBScdPLzILUQAqI+ZjDbSQsafX03v+uSsUP7X/RraqbZ
usMXGM4SpEzafIoJj0+PYtEczX55q6ymyPs3F0EmNgDZgorseOSx+Zbh+O/W
y2/ZC5OF60mL2WqPQiZld+N3Qez8a166IVwENwVO5vjQAv18DukGEQecdNsB
yiXj/rCJDLAgC7wNZ/BKOzw14xS4rC6D44/ZSM5ToTMFfznGURzDf1ClZAa6
FiRGbe76SuIpbXyeCQfMW4rMuvXUZ0m8kFZZ/tGU/6wIX2rmVV3l7Kf+CfOk
D+kUiPa0XroSZHTJZoY7GfJECZOq39/57XtnNEglnDzRxZ3/x0K4e2kT3TtR
TYNNLRU3C5CZ1jlamBBKe8TKcyrFV2g02kQGjc+u77zUteQ9/oS5YmX7HGgr
xfou4CFTrdyGEe5lmT1gRJJUkgZxFvHqtAFg0lUO1TSQ/+N6xrfm7uZnzHWv
8SoMcewIya5px/+2zGg+3mmvApvu1wY7YeFa9eBlFp562lSy5PEQ79fP/u9x
mTIsZwDEInNyGPHMWUDPLqmi33UuuksIUogfuwjTd41bUvTkhXaH6T25TheQ
582qxSdeOHsqhi9hpAS/VoKsj3+Y5+Nf8fkx2EcMrPMygUvi4jvBtTAXQGrL
PLoydVvS8nKP30LWWTCDy+uVlimT31BrcF+QkUzPl5pN/otIrVdjKYXXyM2K
i/FZibAx+o8O91L52L82lOslh7OIcAbCle+q7LEL32d6KyvOPozhPegzasj1
r5+2p9TKS+tgShx0woen5JWNQnq09GpTYBp4H7Z+yVXzwfDjTdAWPK6hWpeN
FrgWGsbqXLWLCbUtp15RivgPceWkLQMwP2gDEC9B43j7D3tMWud8fpkyugAq
Ljkc4F3djBX3dzM0m0IihpCjKcQ/9+Lif5LFPUiZ9PAtUoxp1xQYHTjH/BCz
2b+yoI099YvzNJ2jZEGQYu6bByn/GQfQHzqr0x9zB/wmlTAnUcZBmcNwjflg
7Q+THdVdIUBJMGXaEDiQBsb76Fx0loESzF+nflfIUwaf2IJyBxFy1KSdvsXb
UI3T8YCvzs3qmyb1RDlhjcy1T7mSWNgNWcCqtxQ0JDStAEQ3bJubmiCCY5ON
A60g6pbWkDA3iRoXO5FjDJZcc4vF5z214JmIQr1TP/onlA7s0+3Z4CtirWod
iZYrt65/Z55pVloD2g85gRBtq69TMmeLKpETIjvXiUF9sg8QDQf2TWXFBUq5
wUMKO34HDHRvKnEdG7dsdA8TKgJLbqWBUewjdkblhl+Aap9kIWVlOvba4t81
+3+5B+bdvte40JcxegSDodPyAUs/ADDkeKwwC4kJzadJvn1uZcYJyLPHvJPK
0y3un/R1AEHHm0Y9xYrOOrsLZIEb4NSJYpW8SM6i+LazIkp0/xVcXdzGyh50
3ENsmjrvqrhuOCjVa5+jdNmUgmm8a6Sscb9wrX85LfdvAwkY9ckdbbiBYLrH
HB5FZRxsfLapiVS4TNgtEboBMOY08XQyoeqnJyzJ08u84QR/GMeCJ9mK34EL
tgdeiMJjXaVYXoO7iomXpoYXSs56VqzZPdHXpLvFDq71IdFV61VN9nWWKusV
4NO15jl7+sdowhW7JPBouDkjtQxH5+Y0XGqGin7sEJjTnSMnTjBZtAibfe/m
fwAwke7MAoRtkEw2ua+Vn+qrc0cPvkhxeO66TOPX0IMGGWLQs685lKz4qB2R
R8eppvHNnbZgFd+pFyRsDgf4WuKo7MPGz0PtxC8xdVqkUu1F7QcBUyhwrA2p
+l25mQfRLONRUfJxPIcbbd8ECTHOE4cPswQjgesRh6zfz/7V7PcCfHebfm/Y
gRh/yGW+wKWKF8yBDvQo+0nf6jjEM/dnxebcaXxzsVBLWxVk5OgNE12NaauV
CxtJhWfIFpwxJxGwf6O82M0LPwNsoOFbtnrXROg8CN2LqejeTjWCGEYFpY9m
8sWuscIZeSyBRZoN9CVAaiEl4GEzscPIy500ZKEkTIqfrLtARTSAfoGK9QF6
8QrV43nELCpSJP/0f4JL8wncJW7+CymoDMHmaFL+t/W511j+Lp1Nn58kwgEG
9hAB6RmqsexzX2bZZO9DQvDnEg3Wc+cRRBx/PdCK+qch+73WguIlwBG8QCPq
r19R4ZxGOP2RPtSs+HNC+xvmj91fYxlZd23mxVC8S9BEbqgO3pjul1Z8H043
P+uXsS+5/c7tjeHE/z05tDuwxNd+Ip2950Dgxe04EcQDHc5ill+8Adyu37rx
K4ZKgBNZPRpuiOzpt/qjxLw4+NDWhQlk5WftVLk7+YHyv/1Rtzi9Xz/seM7Z
lyZz08990IKJXU4G5ebcHheTdUwIE8YujMwEo7+iEvml2ufSvDT0aKXYnC3G
/84I0Of0thlWeIclNBcZA5ZHAnbReIT1YgTgW1jxq6ftEqxFHOq1IQXwYWV8
BxPEop94BtDIp/cnwAB3Xj7y4V8uxnNJQkkaXPxou1mfaUWDW/FUd2pPQ+Ut
ZqvFJWXhxqgVgzIQGit30S0IfKAZ9eYW+M2Qi1RAAfxFgRPM3XsKAbv2uBxm
jv0BLJbmnYsCpr9JaSisbsj+TdksMQiSQMiYbt+eWFcvM7M1hUfozo0m5dNX
GBTDkKjkKWDlj6Oe7nrcanc+9Riipnw/R1S7f7d+6/EMR7WTus7Wwi7r8roO
rD7EKxI4QeBMjAFnp6nUl+uPayZk6Z8IKGirky0977kcG819xNnD7IuUe8lk
Hstapf/ZiR3izGfwntMky9mUJ4nkzzx7O8NekfVpZMZug3pJ7Yqh+ofaEB+9
I7FcH9eFAJD0yYF9poqNDQXufKo/UREF1YTPMCq93UjKh7hdZCw1mb1Ma7Oc
mGlKDrNX59QNXjrwbYLNTvGiXiHfu3mZr9990+sDqSE08sgJjTM1QxuZOBzX
ubL2YHQ6vnD1Thh2ChN00BRnNWBcJJAW0AuayBomwSTjzpLUafSQjzIDUVwm
eclNx7SiBX+9FbLdAR6oBsUgQlaWJNdYjA56FgpaPQ/JDghg8F9E7l0Pow4U
CxsJIp6hfwnkdVzFvN+q29O9idvG5L1JK7V/oD6evR9vWdctHut/V1Q9tulg
Wg3hlTpZyi7CuegfQ+e18v6sSD5uSPaGDNG1EppWnaFEdRRRDD7WoVJ9nm8K
iOCLWYFFAVQUffkjaB196PB0NELLMXdvbFTrXCdT1SxaXpwLrX09mCCus0CU
1hnvByMa8uwjU4j35bJH1xhdHCkbSEez421LFBRgyQYoYTdhYUMl8kbxA0dd
GaCCmjekYZfF+lZBCwRMjYB4PGHwswBecFTYcCPBSF7e7ShJLaQhTONYxKDK
X2mFR05jOBMfC1IhIbXH09sN6BNapujYZN9VxeBXjqzTELwrhSaGYqPIBk5o
Om28VroPg/b6RnqUBO5/0VCfvXG0bgo4oE9H7gUkYIguTKPbQS0cY2kbmOYE
NfXGBr43RZT09nec3g2xq0c8YXcuMUEhbhFikbhIIaQ29CTn9rtE6vnKEgtq
9Um9ex8Joep/8MYFv2R/br+yx+1tM23BQerWtsUJN3K08h/Z98hpH9MdNH/2
4SvPcxijyPlsDpgtqskOWm9dtyU4N6FYnImc5PXFlVF0/+/eZlgL9OIRSBDL
l7RH6JTf03yTnS6wHQjG7Gx4AmYKwop3ZzqPaydJERz7Mza+XHP94tt+yC4y
mhcJIGsZFDqNOt2VuX/dUHb/ds65nI18PJAdilqEBh+WhNCS6MDkc0y9n6Sb
Rvft5/TPFyRZniwXT3vYp5I9l7HiYXSxWt4dwLScUukhtyklDtptVzDWld8O
tqICM+lC8mJKsKqCJR/whu13a5sCrfPrS7f/y/2ypa1rIo30ng/y9onlTxOO
KCXVI5HQQzkDYlCwdqNcLK4d2FPLj4+EgOQyT0zK+kixY2Yc7KXhQu4zA08E
EW8vuomxGANEw3wh7SySBehXLQ0nkbOms7VXaHQIAeJEpJsedkWikB8t/X9K
DHuWJVMJRCijUh1CEpTSZ9yZnXUyiRqeXQEcek2codewR2gp1TeYFd+qoxWi
KxpEK7HfFnK1lZmPKw19Jc6u6EuzI6mbnJVW84uYn+Sqz2TI2zdOx8o6cvzp
SyTSNk2Y1VBRh+YuQ8CSxUiKkU2R5vIEX/LoRWqUf5fpzeO7WBwNEkozIG9T
AuPJJ0BHx9GN76Uk0YySFe2szHL8brCXpF8CgTZEh2GZPPsH1MAmmHr6//VG
8W3++BLa3FbcMDA7N1zU8U9Dlk5AqyBBGCLg/ExMLyPZHY/w/MJkbAbsVO3x
yelkphEHedLDixyn65OXUgnib7nXnBRL/oLd4y/8xk9vgLTSgV8IOIRBdLZk
z+l6GA8W9TLQzDUl4hDV/wQZ2a4xGcDLh7AGxVqEYd0zAh+1Yd8AuYVVTjfu
ITTAKn84z6TOT3iDyE2QGUP5yl3UzClB8Zg/oVGpEFDFDSbQxUN4Z0iyzwn4
mOldJb9NwxvlRKKe6bbaWqD+R1bpfBW58ABjVODQt16/22cg29qycBggaycg
zyFgmG2gslXetNMXMMeD00rmQzkVSWtSrlwP8syvEKe7L/Mwce6zGQrCCbpp
JX5+sHb1jRaxjsnXDM27sRw3S+7vuPme8zyhQKAPl5f0ggC6VTElr8z0uE+U
3V/9aCMLh9cBuejLrHNhvB2QpGj9JXt7qE5/vwoLHBbQ8k25OfEa8+Zu6Y83
qPnfM75f2Zjenns3h/ExWDNSTwMyUrJy9L4qUQregXt/DN5sN81pF4J3PNPw
/Kaa7+kmqFSPie8jxsbIbfGF8tdk9/b4hBhOoadaO8W1N8vrCZz3Lk+Cju/8
5Yp43FdA0VznlAVlCdSmzTV4JtNPl/JMTQ8irpBbnPBJug3cevfKnxoEsZJt
YRmC3T0DbOnRI175ByQ5IGkGH8bD+Se4ZBIC1aVvExdf68hGP4uQ505NwvWg
+cZchWpHKpryg20VjtorUXJnjCxb6NQrgQEzHZ/eLjfp2QhGy6FiHwdrv2KK
HUApOaWD9Sf8y32Md97siNleaHAAxtH1lqsko8QGRRyNgjLzxkYcaUSteQSa
38f+gNc3w2Yp6jyOVsBPXiOQB7UK0Xjzqo7/oymq8ueIu4Rlo+B7RZtv+knb
xj+hKF0XuHChZ11dA73LORl2k+Ojo/lQyYnklF3DspEwZAcTJM1u12O7N72j
1uxmrF/Ns65yEmfyeznMxhNo+PtA9EXHu9oGVx5oOMXmadxHpscCWuQDcIG2
N50439y2BKcksfxncFMsr9QD63bHypvaaNxDaEoNuMkWh7wamn8j3670+nUH
y1BkzfsK8aY5Jwzjc4KRPK0BdCO9f0rkJfhJ11mImfKJ05xhjQenL1C/Vwkc
Bld2AfdW8Z8ndueuZr0cVmPsgOIUPAZ9w7uT13l8wBpCANf2G1txp2yXOSIw
40Nl8Uox/fqMH2CCd/BLrLY+f1P5MHaqQHSCooUC2l/nRBsbaOOxF1sjn3Tk
6LAellVR/BuW9j0x/EzMBWp8JGnvCsdlf9A/e0GHtq0eE362iALuz2gcV5Yb
HUwe7+32X0MRMckRDTXgvi++9mmuRWA2AnljofkBgTca2BryzBC4NY58LAEg
sAzJTXDuloIfop4VPRu4BlW69VcdZ+0yx5HfjjumjMc3kiqdncJJUoByhnIG
PFFxtRPzbRGKGT//7FUm2jlqOIw/glfxFHnhZEhZZZhuSgx6MkywMBpg4EEz
AlbYOxbIs4wr+v6jgOFRpNuZ6UOGoylssfJYDGQm4JOEAVYYQ3Xjkgg9BB3U
cJeRp0NA0aa8EfsEhOlHr+8GztALdDjAdXpLCm6u+ojAyQnkQ1Rwme190f//
m5AoSyQhHNdioW6Qkas6P2ynR/ZNXIaX27nnEvWASm8jaAq8xXCvDFn/WnyG
XKcSdrLFcJrSmeCuEnoeQBr6qHPJ7CAXXAjGQuhH+xOdtsS5dn4ah14eEnxP
aFu+jRSHIkjknrez4lpsxSe9EUlVlPGi/nUI8z1JH8n3UOfRn1fIFDZcQPsZ
5kHO6GbQ6tE6L9wccQEvYQJFN6bv5FxzcaOdKKYx+elmR/Xa97Zxo39g+kRj
2LJ9+2ujJZRep2Z/NeYs+wzCexH0Ah88XAEIF2ReD2LuAoUeOeHl09Q0HrUM
HQJLREkKxRGjPtjUQO8RO7EswvU5fIJZu1dp2xREEmwi3cNlsXsTJy3/iMt5
7TFC5iGfMH+d3vJEnb7EirC08lunm5EmFuUMnD8pp0SERTQVU+Wqmq7+cdYd
4zjKCAJyxoPq3yIEAhUMq0njn2YvTt5OCA1A1q7TUp02jn0lyMmuilsMXdnA
cWbXepPWWyGo2nJr1nMfp/z0jplctoeOl1OBPphGXfiCVPBM82y9pIGKKskP
XeeBADdF05SdwXPaCC5v0uIu+pkl24UD5qOXMJVk1FpKOv1601oiQIVD8vwL
o3RO4IDOzcZwtGU1nf98q/WIFYBmdr8F2bPqJgKfIBGfrAIxGMEk3/l7xLP1
8iq+LrQDtQHiyORj34bcwlwf9GNd2rh3vpgKyyt0Y8XFeRWY7+SQmH7sHTij
ZRk0/ynwRfRbZyXqiH0jLt0JqoT4DH8z08Htt65fNFKtCAsawxzLXaKytsvC
+I8I4XdPWhmAiyKgQvYupwbHm2RWfcvCQ/CENwMfRt3V7XNkSyRVAQ+z1KT9
7LcVzb1SUlLJ7cVDjaC9aXW7wV847KMaL1+mqQ1p7aEgG2DwearjBcGCOJH7
GUH0gdzvMT08JOmIuxKzEd5uh4r82YuV/EU58MOnzSBFq5d/6UvoW7fTNaO1
jxU/X2J4ElmDKVPg5KN4WScNPgJQxj5tdtRaMjdwxfwFUsGFj9+TYM9PDJxk
TgJLOybdfSR1Z8S9CqVQ6bloIst09Lc9+mM7qxZ1hgAdrccrgx2Uq0rO1/kM
bC+ftgh/tB1BgP/JPEA+IrFsLs+ReyzS1JirQJ9n09wWu7vTMZYKDIVFXilt
vmuMxTfeVvWpvFDWzDsCBns7WgR+7tKrvG/0laSBbCLgcLxJk6hcuH22RprG
hN3OiWTYTgEQ0B9oDyizs3izQS14BIoprWT248ZBch8n4VyOW3p9PuhKXnHM
BINsd5p8BBGMPxtL+Sqx9PvD48XVsYs/Tz16WIkHuvn8mw6pxqHjGoyurzGs
8t5EREON3CEa1lfUzoK8vQRx/BXoXMQnoqMemXBrtJr6jUWbxEtXoNganP5M
lMlr4Cb/ZR7ZP0I0CW/UBI7RevaXdcay5aq3tAaGll8UK7P5V5qVK1gJ2qWt
5ymWm51IZycfxILHsaU/T7nVy4+LRSfyUjmh35yrRnfOpZDYhSBayvCgZPem
p6lROinFKlAod97P88EysJSQ0u2pynGT65bp3MLYL4NiaI98HAJXMLlmmFAK
axuFugcd1BPYqMnzIeWbH7v3Vj+7r//O5Jv7REOqa83tt977r33dKJVwdc7x
8tDRpB17IYbTsgOJhI/K/qjDroy87mjCJ6hEBK5C9mn0ckM7JHUDr4lJrCw3
4vLCPpluzCKYFboKaLhpJnjPM4ASV4b2yVookA84oR3kl0iOyRIjJdpPcOkZ
ctDB4zJUkUXC3wfk/fNmUb3r4cUgy/mo2aQCfsjIaoGUn3JZMSPtvSVB54lG
Dq3Bi+JWQf2AXjaFchXwMDjRfM5D56GxAnby5wZE+XDjlwhukxq8SgnIDcd9
FBVSR/J3urX5jQ+73iX1NQqWUUzWoQt4DzhoPlKf2+ZQ4u9dDihlkPiZJtRS
hxBkG9c1w4gwrGgfmZdFufo/PQliVa0Z4bPMPx+YX2iba9n922ELl5Yt9caX
0rlArHLulW4bWGkEx/Oh3HzMSeoYYZtMptkZoWvNAoFrM1l/VZjYG2csHFh2
149VyLqmOvayXOBinWaufMgPkc33k/y5RE/kfhMzS+o9AByp9Zocrv5qtK3Y
W3saiOKHBWYnRny9xjMqtUWsjXE23Z7WrbfrLHssard5vmzEZZ0wb+yNyZis
+djHNlS0zPq/wkIu1qT7awpAE72TJw/y031pM3W/7KhBe+Z6wZQ6vZ79iRDu
1wgKLTHHPwmzV/zFusjzjNshzo0YuQoWr2sIRjs81YqUgOPRF1yL4ekvZZSK
1HHbo3AwSzGxYbkhY9sHftCDJQvtgua9PlSNZwVBU1DkQqLvdWlh+7UM9cuo
3Rk1/fx2bicFIsmxhUW6nKbVLP+pz76Byj333Yl8iFCXA+qUeLTBS+GHYqX7
RYEHDCLKolGMUcZmI2orUb4irvWtgGzMDm1eqMyhT7x9z/IApHBBv5kUqKTP
b1jHUWS5WLzxD5AMtZo3pHWcls5mk//OF+LJDrpkYmDW2o5dUYp5XbUUAkXf
PlvdCrjbDMEQnpdrxjd8cZS1mhet7JSUqM0iuwt6FFzfi9ZReH8r2hxxnwac
3u/rs0S6KwRSzdUSoVn1KK5cmwBhS55LPtRVC4QKc4D4cndXhfBg0eJ+765w
FJ++lKa+uahmIKE7YEZWwZnFGnORz9FcCrLooIYOEcaercXupR9mG9sU/ru1
axoP3XiC8pGgCSrKNCW+wCbnvGjscrq8ec6D85SJVFgpjvUQE4xDTBUtQLln
DJXM1Qq73NEZLRwopGJJuSXdstu/zFkLAvk/vFE22lMHTZwYrdcbjexf8eqU
PuLx99J6wKXV6KmS3e2FmVIUISjIptCbQZb5FuZZaztRbgdUeZzqzY1Kj15Q
S/Yw1RkRmn9ACGqfXnoDEJqyTVTNfN+o+nkRitbqkMyGVOqTY+RPpKpQRNoA
TAbLbtp1q8Wqv0AlsLh5+DB3NsCbwO46+kCrllV2gxlbuW5tw6uytdaU3bCc
qczSvZ9HY6w59S1T8su3vryj2TeuX2tT1H4OKWIDzIdTPevPJYeKAXA3iFhG
jGKSAYgcoiu70DOANMO3bp7Dv80gqj4roW6wiuuw2RO/HXU9QFneg2qg/zmE
cdT2KSgdGxQ/0otSYS11uhl23bfJ5wvVOcpGVAtAPCad8WPo6hOMFR8eeO/2
mmtVhKDc1x/G+9mJZQaOvn6EYCyBolpC4TouGxSQW+F6BuFVn8mPaHqWuXi3
tyhfKD63JFEI6tUn/ltea+2qrzvPBIYdMV4U6W8PH7t/YCsgwCtHCb+Pwj0L
/grcrrN08wF6Y7vdwa7qV1/m/rb4TqpeKzz0hdHjxZPkRH0Udj33b3/hz3dx
9/Hzb1vL+AIyCs84GhVcu5IMFtmandX1nFlSWHiMTkRHJHVgC5OMjBTi02dy
cYPYoLPu74udgAL/qomJJ1R6C+/zeK/sIe5xQFrWunzqK5F3cbTFOUG2oYO2
Ru6ieLM0YsoSesROo2dTWyeo67+a0meEIQScWYKoQb8gAytUGA2F05RlpMGC
BcB0Cqaj25iLh8pXN53r62+KcC3McWTrVuRT6A8rVO2r0OmlIkazZdNWl76F
6sXUgJuCiGb7BEiR0zzxjghGV5toIPKQsu9LH8fcy5vx/5yTc7Etl9u/nzeq
tGbeNVESYYZruw9JdBWRWURIOwetHEzW2ZdH3kq2ZBsdRqqfMpKWzbcQncSk
G6F5sve3xajzK9tUtnzvAwy5RrgpOhHKDXQDHOStDX7rznrXOFSKRcAcEKfE
A07uakLjmJZ6I5gxNwtdr47LBIPQwm2cEeuUSf1sultmhtz8wFsIwaiAs3V9
abTiXDZBYmGZeVYXc3ySpMGh2aNhmQPvMH9n3zXlXXEkTuwSYt9j+3thRPQd
WBczQeQXmoty6TnnlQu0Pefe7xcT3AjhEciNAvfmzIZpcK844HRM5wYvRhQP
hkrX1qOJJ8vwIppxCdKUet+seZOExkq82ndGE1DxADVnA3C8uJ9Y24bA8t1o
lLwX6s/s+377H6sgQpmGSaWIDaGX0VqwtMqpMU8dP1hXo8AxG1QOKv/PSZXc
jaHwb5Vj2mCQZ6ulnIBMP8XUJAttVqCD/IT0IgDu/VXnfsv61EsMkR7+pRJE
Aay4cbxX2QNH/q7qz2k5J4ZiEhuDHM+iNkIQsYaWlYsf99koeuWFYS9VLbNy
uJk2qCbS57+ADhl7vgiGc9TAb0uUQOc1xB8DJCb4/3Hsonfsbv1K7WrEGAQ5
Ur/4UZBHKWSeOe8oNBt15GT7b7TLNG7ntJDUDobJp/Tg9fUikZLkhtBOcdwT
84ow9Zbro1eUFC92f635mfUb6dL9yMl8e760hhGYsWvUDMTwcRUPcqYuj7Z9
T0kPlnh+aQHged/mJhvp/g6mZdYn1hy9KEcQzxw3pKlXNqjrvRXn+FXalH8S
N7wauaGJmwUzeTn44xS0iUkNeXXOlxPZIAauJg4oP8pKw6EtXb7ym4Yp2VJt
HjyzsJ8B74R16JjRCU48k+dqAsw8QSv9aXnI7iJDAFV1B4Xo1cuNjB1e85Qc
JY72fz3FVrbxWhCkFTB0SCKEYlmTzVIIfnWCPogip4ctcTI9uPvavrvWqUmL
c5VwWbsuCe+fRdpiYsSEqUONJHO7tx0VNxXQfgBtfrjuLWnrpp6HMeqx0PrM
p75bCtNfQTHVG/LdtaX0JC+/Rdlb1cSy6Oz1S+GH8Q+ebnH0Vp032NOiJrmH
tVU2zOs+FDuX+FcK/IbGWN1rysS+ut7swyk2BVKs+CT8jrxv5s6GfQIfKuSa
u8Ykv2fKQ/aZfCsrBAJSadcX+6Te0bB45vuPiJWNur57dwNJ4G3znlQbZ0cU
vzLtw80mae7AS8GCXezwSFYNhBHkJ8zzWwlE+MVJL3IzIO8+mi660iH3E+/+
I/Jeto9fJNNzEYakxWsX8kFVDuR999mcNaDwCifndCuLtl/I0Gt4C1UqqGmi
PCjdun0gxOX72P438cvf7z+3drA+lYrz/dDk66OpgeYM/wfbPjnFlxB+qDqb
hjj5/6JLNIbiOqr9QlTO2kEWB4EWC+X5rYEOFQdK3FS1XMfqj5u/aSsCGUEp
Y10moigxMtfWwZUaZdOtnaABvEiirMbSKyIznCA5A+K+Bls4vadjZmczSSHY
BcYloBdm3GAjw/0TjLQ5wT3XCxNO8eIy4RA/L7mjHHOjplN4b7io0pBcTSp9
j4bI76Io1s001nFuNnJgGxiG1uAVupq8snrtZXsW/evgtYE58YhRha6TxqHA
7g/25swQGxEZ39Qttpzuf2mK2NLuLzQQYEW4G4HcgXW9+02lxRkzHY+XoUs/
chtMMqTdCyo3Qx8WecJ1sXhj++CSCJa0LApGCXjGfVJCCVXlEz/I8ywedU2G
mIhObUdahTIOIv4erx53dANayOAUFymnQBcqfP1q6vf4wNZEuZNtBjwpiwXI
lPR6QcpmV0qpr+jBYJ2O2vMrmmmJKHbYdv/2xZIUCijc5tI88+ss9V3e/1ZT
GG4VY3nHisvkas9+ApWfm2oMGVRMVlYnDCm24VPKwE+B0ZOlhasZlX+Jhm6D
9ww69cJcN6fz56s4gV9STrHw1Jr9BNEScGvHuJ+GmQuxXLbCgVapGb+f+6HN
qkPRgl2A6QMisoIQ4jxlWPWNK9QgH1iLrUS6EUYfn4l/MTeo4Z8gei3c6I6p
IG1b7nuvSM2SwIn+zGHllvWa2RvXgu4KFr+xSBcddD5rfxq55clh6HMpQ5ex
QHZItTgEylOaByDWpyt4S8KIzR3C5/ChRQFQ0IMKJ3fYk1jISE+zfmuqkov2
4owv3FYVGIA+okz8eVaoIld3QMrgeefMoQBEDiuJDo3gKTpr6aHowR0qx453
FFLehcp4dtFAJpN9e95sGUoVMPDdjgWu6TvhM3cpjloWPlLV7IYei4aS9uM5
FvccjmQDd8Z8CXl4RFlgm+IM3btzLo2xVwyJbrMJFPIQ3gmvzQ4z3YsPK+Oe
iGKKlkfLeUViQlRJoq5oylvWXlG9esCucfk8qvjHEAPrNCiVntCPvldQyxs9
nd37bZG306jXnsQScs0RoEJk6szYFx/egnBlyisoO5CQ12s8srOV4LbnR+cv
iltRwTBFUaSfxTv7cHe2cl35nL0mrow90XsylQ6k/hhTtHIzWITbh593rXOR
YCIqRnCy1L5TQAbFv/LYEKgiT/dlQFnoJN6lw0WS04HWbuB+ipLhXdeN300k
u+vmUNIBPy6lH4oVa9lh8P7u7TY5bB8YjD/I9BFSZpQ1zbngc2ZWkQzd5/sl
yP3aNzBMWUaI+LsTWLZD3qefM6G0N8GdDKv+hQY+PkBTz4g6/fti/GYsE70M
8EZmjzkjAsFfNBmv7D8NANKFr/WENeEAS0tbJsyohjLGe22lHdbiFOB8nUmz
vD0OmHKzMTpqU9537x3qH8wMmLpprJUkGCzxjv1AM6ax+kMknb6cIlWvUkpW
jX2My8Fe0YBmGOwf6Ij4I99eKMy3Zn+iPQUfM/q+g/PlOH/Gqat626+H3zDx
pmQYs+ZI5uPphYcYwhr4R0ZjWDRkV9a113Yrfj7BteuhpfZfHMzH1AYfPIWk
bOaALSWhv6NobKBYFuf0UPyQ16Mgj3IE42U/FeH7wHqZ3lxIgCk1PM6hqrnV
IH58XXjRENQGvw4BtI83T4B1Y7PLeABy9ClMHIe6LmnL/98wxQQ+giorDrN4
W3q2BRQY6dDIEs/GDbLbWhsCLcBjjsdZkTg/ua4EoQGUAcp+qZ+ppSrI7Ya6
J0DK9ZwHWLAh/vaRasLp252kcG4zNHyN0wuHsmUWfJMIVGy6+8DMotQa2O52
SuBmoHBUoBrYvcAC0hp+CujiosAuFxD1VTvn8G3si3KEmlqj33zhvqKB/LC+
S/kT/Z0pGfpQjYsfF18ouwknyZ0DN3cKutZhZXNlMAgD1HEKSvY5QFfeV/Na
4pMwS4QAWOuv97UqThWThJK0yuDKIn0yIsxKLqp0kJhmpRDConsJVQpKEIOz
3i0tDo+lvxN096YBNwR85WFRxpIhe/4TP3wCdxtkNvTdPkvkWmw448a7pU8V
3C+6SNLnExdMOiFdedizh/dQNZoX5lqUt4ksEXeNS7hPj0FyI9GgrBw3hHVE
Wibro6hD0+/LuEBXmGSka9tKK7j6LcU204hFUY5lX9FkJ1qbpRl3JXBmAvnP
SYAzb3HDjtkqHhrrWD8zvIdTNlA5e9ponsxL+kIplgctsIjCdv2rq/5XgKO9
C/lWt18JOar2ERdR8IPY+WzIFlcGRgUiR1U6AbkTqz2bY2KKMR4KEbWsfLSF
Q90X6QW7ETmT21RGOI4c8bbNHJY8L1HQeny+OLIDDbEikCuDDcdcUjmhX6jy
vJck8No1C4jffn4yYsJ++DRXO+2mihpHZJMH9oF/X+l9RjiXngKjMRCHs0vN
XtCdGndwf6y2KWxqosMixzcSxsYRFtTgyPjYCf9lWu4QKvXzA6SnaweJvn7r
yoULUhkAkaqEhoac93Ca3QmT5fO7JtiWQj/m0IHqJBq+0e+XJ+sR5p7635O/
5QWjI8GGwhexbzfeCsxPbRUf6YW89yl4e3Oll6k0YckuwT4TecHKWxwSYcwc
Ed4n6sKskqZC10AiT1iwaejW7ZtrtdgH0IToFyw+M6GU9NsNDKnoabTflEod
tEEdgcDj8uakurts3uKufiFFcV5N/vKOETfk2ynNpTAzwItFC9v5agttkAKg
qmw85R8GrFQbAk9KV3uR9emxfBXaMsUtvtu9Tq1FEVHaUjdeeoliuOCJwNr9
Fcy5Z3qQXiTb/rPe0pB2FS1fNSwTqB9ua9nM0Ug2uqI3lc7/23utQ9k3hQ7A
+QomOftqkzDUZ645T8Sgw0VdPF3SitxraUSOWvVYHGd7tHB0WFrFku7rAlcz
v3283YLiyeyxDczY5Z2lcwOK5CTYJfluhN0KwMyuU1ce+kK2+4eTeheck+NK
uex7AF7dDqgeH+t2PII+Uh5/nJjQ2PZkyav14jMQmpq86rd6Mgwrk/IQE97d
jl+ldr0IL9tKYWOT12Juzg1+4V3Cz4KOWqwn9Makl3JD3Qs659QNwgKc0fJw
AsvGK5t/2tRWVwqjV9lWboZqscqMqHbO1vsnAeTrZ5HJ6+0Cmqg0DGFk85o3
4QNUBUp2X6eCk72r7N1bm/NMhTU+1C6RXvH+0t1mC1kGemZ7hOxzlTsIf4GE
qSKuRymT+iyoQdfvVilRYqldqrNc/fGKi0yfyIFZef1WF0lvyjltOfaLSULg
FVrctA13GtccFZMQ4ftrZn3ocYyf4jtLRlTtYeBKmZp4q+MElNoMPXPZd8Mr
Pw41z862vhGdQL+UU0Oq23ikGl8tnDc5YwNzl9up+faLRobkoJq+A0wFS2qt
iuWXqlPw8NlGyEc82QWSKZsQiJNQY6QMllxSMEsdRLrJQ9LCR+AvfOcVfnhH
qwTt2AXWEkgjtWGDHNyuakibs9NEbeu+c4/pjkCYOqCx8NUB6TyBgXt/KCoT
RjzgQwFSY4YVhc/OwavI6LYwS4psgfp5e0kRjFAp8VTYDMxf5lnwdsAWEeMJ
PDjpodCGmvhWDMkZW/BvRNZMSmMcp+wm5gDGRLHPQVvkWPEpjxFgjuDlRHJl
YAFx70QUOt8CxY1EjgiVC9kNvsMiYLuBAeq+JhXpJ4mOq4Ywjgw/8oFu0jtM
XiXq7cMwtEJtAmTshe+AH+dyXeHtFnfLddCjbZBMc7UaoOzO3SMAMW1NqKFy
LF0/nVABK/rkwObElcj3/6Pcq+Ac7bUY/5tn6uYTGpRzbseWiU3LMbsSgCKC
9ogHjV7lcoiyE0QEY5bR1o+aE4ikfeq1zFiX7c04ZLDZzkfhZljc37Jh5BDn
hfm4f2nC1yN1wW3CR9+hCxsEzsMe1jaABfi8wcWIcLQiP3541OxaidKBFmIv
sh95Rjk/ZDcam6HvXpT6uhLyRqoGDocPxxWollXIpcdqtalIH2H1VVP/TMQR
ha0LSgpMvFBKkR9iMmwBRDQfqH228DZdfzGImVLKcPWp4fct3EwfDoosnSyC
XwHOL4AoEsrSvzrXQJn1BrU+wGnPuaJo2ICblpCsQcSl7cNXMEtVeH2a5+1H
eddMSFeeAAUzpoJ3QFrV785iiTooIe7fBpSpI79Qm6ouxI/E9bHBhxgQRg1F
bm8eoMj9dqsRdoI6z6+TZxp0fpIyw+bOkcHkSbGxYBWDJUJE0yIo0hbAPEK2
Flr574rguTndAlRHsFzjBlhWdRAgVG2rt3/seefXdtz7lYjmL02SZNYdL2lc
zVO9UkdobuPu2V5oCxDNcdEe7515ttUXnTMIGtEquOSmpeEXYPW+PMy8A+RC
V7ba7kAJRRWhINyGlQgUdtfJK5bTEGzkayRoAA+KTSsEViVQIT6bPg5/sHgX
ArqtB7ma9yajVc/Dg6tB8f8IbPGmLqwKYMU3S4oCbeLKM4F6OSL2Ja/k68G2
h4rxhuL0rdSjrwDKjHYi4vTQAo60XXBgQdwFCwEUBz9Wxv5o6Jg0wgCm90zv
7WNe71rp2+OOPuo0/TmoSZ9jS0GLf33jlPomiV7ZU2EjWw7Hn0apzTTknaAv
cGM7BVZ0+D0GHhXqr3Hi+qrpwVTuD87ODa+Sz/PR9xWonkcs4zUznFel2YOq
Mt6a9auYUmEn7WI3wnWwrUWy8363Q3cBKByYYQ3ELqhyMmqlashqD/pEHBKL
pPoTkVQ3QBVCVsh4ypvqrYya+Rr6th4awJ11iW3UcdrbisaZGK4o4q+2ImoP
qPJqv+7sekqfk3gLeDTGDOMYvU8wJSSkozsiJBi4fPzR+SYyjrKWFQ18cfvb
y7IM5xNDoZ/pKQKx+9N/Q/sbnYSYFs0CvQ+HfS/ptcsnmkCAVDcnCNyR633y
UQIFk42Ue4MR9U/65DK4CBzs7P83kGijanEQsiXrfhSkwmrwL2GP8cVYElS2
GzrbjRfwJIdf+o6ZNdh58MaDtS2QSyZhRBMAKojfgambpnTqXrrYEM8X81A4
Qulqn8Hm5zpub635PlKWu9yKSIunpCKq3WJ5P2Hg8gqV7fdvasIjeNZxyTWp
OP/YlyVHOXjVqmztbaDLSOu4p4UfrS+a5RTk7lDKfByQjHFKYa+xWyxDZv8A
k5QnbjOjPoRbwpfs1+spIWVd6q6e2wR7SKrHXFR/hj5ze2BZfih9Jdh4FinR
a4JeOpMbNxr4H1MMx6RfVUbL8gjNY3KNP3q6uIbr2fazlhVU1xd8WFUdXpx/
4KlgwtDxOzk751aYNfEN0TIJT2wq/kufA0w4opt7UADeipBwpFeJJZ1alym+
70jfiz75YiU8id+3Ys+WzNSAQv8pJJ1RbCFRu4e+VXEfS3Z1Uptx13Ku0cRU
8M2TYcpQgFLeFZlv1LmzP/eFeYOv5Y4MCRAiXS+BID7NsqsPqIn9tuS6NLvh
tHWGw7vfBdtxAH0FKfheyMCJyWrlZjTgQEFmhVLEb6S/FiFD+qwvRr2r9Ouo
9RIG6zueDOuCJxylKUvFfSFROvhNv6r9RQZ9YgAZLWA3WhvJyIL6rucTKMpu
8B9uD+g3OKNugKfeDWaaU5+apRPqf0wl9pXr07ni9SCEiEgpIibr9fsoA61i
fHxKanxDWbFxWvpl/esho73FX5rQDmpJWNUsEsw7c0wH/kHj/PTKGCT3L55c
4V8XdooVICn3V65475DyzCMhRFPiEWqOm6AuEEcNbnq1KG3kgyeGUboP53hO
GTmP4ES7jt584i0rEXnV/0ZY0tDj7Y14NRQYDMWdSOek/7Gf+MJKAm4wdxN3
4QGA5lpgQspNrSwklu4gtYVYMq6QaBLmkT72g7pG7jNEVSSjSTAe9DY5B5Cz
Xsrk1isvpajXFgDARIx37M281fGUKKfqYOM2PI7O8kWKiwiukukYMNDXUPmW
eKTJqMAecgnSuhopVHYicZ7oTj4tAOeja5XmkBxrluSmSvPXlMXzKBaasCVA
CBOfYl8h+huYm94bNVEKC4H/0LBkrUFdhxlOaJTvKJT911TLLUt79Q0U7Qxg
uDDIfeoAVqkqKry9KtLw9XyP1qkzCSGC44flQYaYVjhfry6EPqjrdbP2ueOA
0jOgD6bbWbEcJpN6slVPKxGUQNHBEBSaXjQIF6Z4HpQWtUXRxz1q4v5hzXRP
cXKFkW3Bk+McNd0KE/tLJoUvsyK9ouOroiKuZL9FnGK7JEdHqXAk2E25O2JT
kdIoH4oQrp92OdpnO3y0XEZn2PdSiOhETtJwTNSKA3JD6EKwdvHvLmRS5aNk
y+wjeOMab9dOm6YcjFCpkFn4+3NARKQptV03Z2F04SSazv/QsCdfScPv74Qb
HWXdDf5DowezrPhsMMgrUJ6R3CVPq89vAXeQHWxwJRS83/yKsutJzCSvSEBL
gF4Eg5xG53N20okOdDiP8uxJRUxdMOHOzyHXGSIBmjYOALeJQVfPClLrMK9p
CURDHEWxxrs8AXq4Up0enGJkEcbe7plIx778fgzddZmdlUgJ3w/u3XLhqhN1
H+eoG+MrDnY4O+YdB50JpXx9p2sIHTicn+3xncJvP8PP0hgR8j7lApqq/Pqf
2WuepoTVUCQGzd0TAoqjLzEK98ZPGphcm2FsJGWDn8lp3bK9BzmTo0D+I8ca
VxNQlu7QWfka+a81cOgmigBQ3vv8YBTG817ug540Y2kUNnFDjMf8GHhqFOnu
zpvmYe6lWnIWfse5BFwZzegzlkjPWHxMq4VqO7Okliiw8m5GFnIPMx1RHHdz
k0qIFaM+PXx7UpTb6CgnwTYUpcAPx1SAZP+4wnyf1MP6btTdODuvytWpjm+k
edKZjYrXtEVgEkKSPBUFh2MRbf/cq7jtbTZp4lND+CFSiKiQiXkDJuKxn0c8
32OiG9yaNjVYzz2Qxkj5xUAkSM1MM8w7eoMUK+n/lXqqoXFCqouS5Zbb0+LO
nWi2i0EHnyKvAlJeDldUf73bfBVu4+RfVm5obm2lJXyYXEnlVlHnnThEcVAR
2pPBg8AMK/qUsvfneHzcXFDkdNuH7UKRCxYjA3bLs3x2dVjT4K/pXBOg24pg
y4J0/VenSgO7n83QOjt1B06dSkb8W+EjYHpTq4AtAXiuC+9zE/81CQ6ZEq+6
hahyi0/El/V2ukXcj4s1ujsmaiGISMAmLQPvnaCKvHu5iDNxItU1LYp1jp0n
RYFoN5CZuIQs2dTsWvqIh214vcbiPK/bCaSsZE4ere+CjC1A7X8vnru7Oku6
QzB1lja50SWII/Srdljk/di3OjRb+9ayx38hCheRKvT1QwkF5Igm1OiKFROG
HekR9YiLHBtQB2e+iFKp/2K+dDIZrOPr06tjvi1QHP3ci+ZOnbHQw0CxNqQA
LEaeZK4boFzytHPh55Yu1RM2e2ogkT2VQm5uUlYIDHnIGSRvIoJYyanwkrEp
v9dtr8upXBJ3dN2t7ZFL0IWXCWmsNXksakP/UhSJ+QIVZhLDwJVZgRWf5ric
jGq5Bx9HI3PTvONkSmC7fCO5jalOIzAjMt44inYIF0sRytmjXDOEv84+EXx7
2w2DCAXmiYRFUgYHvTLTPB99iQgw9pgJlYI2XzszSP3MzJX17C+pid/CLny2
Ums0pDqKNHvz5cq433YGsPyJ2xHb5+pIqKjxzFxxkG3VWVCIt+TcdQZm7cGc
F7xXc+85oTFZPrLe62oK/OOwJsdoIgNtewMRqXbXppmf/Kxxhte9v7Atzua+
8czWAbmTFBb7OV8FSXgxNJndFGDm8tc9qVrpltW1ijVS7E7peLCgq9/tj3Eu
dkPcJUMi3HaMq9D9fcyb3i6Zsz/Br0PPJbsYFA/Tw76edGOZfLpYBcG8zGwa
gk+0ovwJPnUKAXpPB5U2ymNyqwOHKmiu8E1J17zhxQ1zzefZlnFdaGO26SA9
FoOfALg3VkZKPtXNHZ7HRzaIxqfJ2CK24hPl51Bj+nBhatE25f6N9ds5n53m
ieJbUpc/VwyAP9n2EEdFRjsX5EVSg6p4KVCQyiZpq9hpzsN/H0YDrrDJlXBk
C2ZjMWicJz5m7lssS52SHN0RaywIucsNy4O9gaYMGCW3xb3579rjGF4nShvU
JYpv9h87hY/tJSDSWedKRqPio4hnHXDimRlsH/yDdEk9dwbosAXBJHnhv8Dz
8RqdfPCD0OGbUm3rNkc2RmFMPnCxMCYiqFKF/wun+IM/dB5IlKqBxgeLvN58
CNxJiBzWg8ru83RK94fovrAwl3V3yfz6ZYF9s/Ct7AjjOhp0ZEIx2TKVbiy+
F5fcAPJzxMRhdp2XGJda3ecw/+n0cliO89P74MK7qAglsjHZLkZY7Q2pvOT8
4dNrmVaR51tQS/i4Pm2wYx6zmcOtDqPXdzot9DQcKCqHVo/iYrHjxGWEHnAA
dj3jPBhLTBi6Bf9RpbbKJHX5y50+uYGLVgaV09Pk3i57hwo+MEPlcWPvdKa8
MqooRmIOZ6qBDUvoOYFzTXY+gv4MxtoBNFehg6EVQIPUSGVXNFu2eAC/mjfs
EC7nK8G6i3BbBb/UhC+5bloAnIl2ji0uqXJbwHmleyqSnxO15BG720VfcTix
ID23mUEAE2LZ3ghxYHJ8KYuLOv/TA8MvA6pZqHIEsEVhiepbg3M3Fnbo+Xu9
g8bsya40YEWYtCQFs6xQi0Vpx0XaalWmEEheW0P0X6ErdvlsAloWSGt+JcFU
is8x8hL6uRaeV/qbXU0UndA+QVPHftwiWZULknTSuBhW+NQbP3lSy3qSMaRx
2OVPgjYB8p2yzUy5mkV5XbETQPHn+VQCLoFTlW3lbbO+rM5NxvW82/Q4vu/M
WJNEC9RCz5KYHniY/b+jDedPJAXemiN6e2o+JA2TVEbXKtK4PT5jtX67wRdB
k8jwI+rJQfWLq89wofjPQuuRAKoa4iLxr4REXuAhOc2FMI8iFVnltR5d0DkF
VYOTpQix+7lX3wdOEDLqA5A3gQB0tQd1R1xDadnwME1o2TxPMTatUs9Ryvjs
MG47ut8XYsGpT2teKvsMJS4lcyerDBRez2jOWX7UZu4uonuHvcrHvQpWd8Pf
r2PpGQFxrKASzuvU3U44UvF+BKuUVwsg9oYS5mDEBwVXR8hhQ/ThLjv14i47
FpU5UhsaAIEkFeaL9di1RfmO/dHnOLRA8HQHVQ7dpYioVNp2fAB+KJbsQfob
2JzgxhU799+AVDvXEetcNHTtW3/+yvzJJchzQXmZOwNpGtxyJTpYIFex57Oo
cEC9hL/kWrd1FsxP6uT2oy3g/dLj/bFWP2cvm2ojUTc99tMW6n7/ZS//s8Dz
m2GImGKn/9HG9usZ7e5qWtlXkBxwP9PQVlkxSyM7BNV+4ASVOKUu+aCv3MM0
AMFiEDlqcNdzadk9fBpCKpC3BxGwnMNgTY8vOicv5X9YVRLYNCBmKPtAOiXL
JRL0H7/han5Zsz++criJp6RnJ7K+FLW2gG6N1ZnmISaJpZvxGiJ+nt2jrA7X
BUx+HUMTtNbk4TV1F0s4I8zsKZpk3XA+9asWg7sVsxZOUmowB9ncOv7oh1QS
e173rxzjdvGHcxrLYP/Q7E/AerYtmBLzWBoU7Skf1IqVEGQgR1rDfsDhLlfM
Im/a5w1ox7wQxmWFF2sM71bg3gCECAr6z362b/vJS7kIpC4jGZ74x99rwDaf
2IqZNrKgZOG3NydXk480RgzgAvmAjZePmeG7LoW9NypFxq43Fer9M/x96R5t
Z1I7JbyTaEjzL1sX3JsYLJsd/kvrbwB1+N8Abo9hvm5CPdvYdEDHH3K6Ac/m
VoJO7FLjYBLCRThdF0PCdS7nviZTiI3iafKX0yVjHJwXQYRyuOgAAmrc5NC9
2qxW7kybmTIObdotG4CXEyKtPGFwUmxUAt1CZA+dzqLp3vWdwG2Zt4yUYxl/
rc2lKRmGK5JmzGttEWxEd0MnENm89uk2am6wJyXoIHy58i267UAilBaDPZQA
rV9j+ZLleJC8M0ziMbFse1TUWZTCSYRiexDA1KyVnYRVwC+q9mA/XYLE48Sv
UJ/SSN/EJYHz4McMTfoCKfLi0efpR99dapvGakoAyslTjiykYGOJR69MGF9a
ahJwC2WWq1oBvN79k9IpVUj7tDcPy0byy7r4TMcvsTIMPS/nTDZjY3gzzudq
heWFi7tVV4Mp8KrIJTA+eixREjijz2qTws6T0fUMrrkCVr7TGyOnRdaBuHyM
Ta5R5szqpC0XGTmQCzK0Os7Wj0tS+VRwJyTSv3a656+H5C/JMEQqsQgX1aZ4
+RsJdV/niWXIbzbESnnFzMgSLxG1orouvbNnGV8F8/he3Mo5teaE1pIXc/Un
n4PHzKVJtRin4A1HFoPAkGz3h6BgHvNOQkVKH7BvE9sxYC4d4Gm3/pflV9EO
Duk4OpApYR7XRdymXyrpGYRqYZoDAL6Pd7eg+vr3PXz2IZfz4wzDI9jfh9Ba
BWFxVNibhkNBT8R/2e0iFvAttq6+0TOCGPc9xE9xo+WL3pejiGzbtopyEJkb
rZsoVN16OJwfa8zEpEaOzDzuHOkJInRvjvS2+IZz2UkDgsdT1kS23RXaRmQ6
CVZ5CetnCClJnhlCCn91XS/SR/kydIQZZkLxDJdmslskXF1xqDRduyHCwuY/
CVgFVowcg53y5M7oBhGKxt99U3wUcsnXR4rtDtleMF9+5eHydxsmFYcR2Tni
yQ4aiNSA3OPcG1Hxk/2MxeKN/EoN9ONTMosQy/bwC2aVgk7p9kpEzHoyX7bU
cGIV/aBZxifg1M8+EPFkTWyQZHVddE327fQdtwCyolLqNXFsJUFIHA6Ejjaa
Q2vN27TKVWs7ctX2pnMfwOeF4pGf2ctAWr9QPW9qoCnbFEA2WNGlGQZsUtQ0
1LvtpAv5tzuhPgvYmGySh/sbI0u/r67QqBfv+lARHI8EwMAMrKpb0KJEUUeK
P/VE7RVO2lD4jxMigW4tiA6lZGLkBp+MtepAxsRvli8AaPo5pPUyB6m59nnP
1nWNBquo5fW+6QPj29d8jW6+vYwCmkAlV87xaVIfvZzkZZBaJIyv266L2E5Z
d5B6fhykiwqKbYH/lmMuTHvRJp1RuV32c0umrgSYr+Ygk8gm1EHdJepCxmfV
GRt4L4ZvVfDmUSBIdHhFZZ37agYek8rrn7OZ5cklMuXIXMI+p4k5cMR+ZkqI
bn7DRUxrtgVKAnCfCHMIdN8GQIKiM2sOQG32nLPFYOGRGzoYeiZ7pwtNkp43
hjPJZxiWtYa10Xj3q4BCAbnp2VlzHJz9K/w8w8as9dNIXe/OGzfxmUIprkNV
M6r0a13zGkiZ6mbV48N89TSap4nIw6XgKeXZALS/GcLbJfAy9fm6I03ec0zG
16c26AJ/A9UHqZm9fVX72H546p9QtcrNrMYL4uhwSlMQ5WqQ+Ru33nbIJKm6
vM19oRrKpT8PhQIUVIVqbSbndgWdUE5ojj/KKknpJ4DSmmptuaktCoAKl6TB
v4FtGdEdU0g1V7wiFKGA4iBE9DTzx7nmBKi3fqw6cdrDC8W85odXIdVvuU2B
NgMuuEPqARKpbfD0hDeHBzIXGUSmM9s0LOPboh7pqGj/dBvwxiT5yu36DxrW
SZiH3UVT2ffuGEktWAtZZwnrkmZsSQY11rP9f4wi7WMdUsIuZTVV+/vZExG8
uK8I+d9D7nqOP0+wJDJZP/nfJvwSq9MBNczU+mEoWUI7UlDgG7u65w3mKWQf
roHv/lAGt8fQDmRtXzykSxZM3M/5jbhshbs/8H+BI0RYs8vRjn8mbZ1U65Uz
DC6he36WRz1opDn92h1eWxiyIQxJN3hK968Etz8FsOHfvPylkM8XnRoaUjgf
5NaXhs+zBw+giLpfbEqeNYVXHiX3ucWJCE4zDGmf3Txm8sOEg5w8ucPTRZAz
gPxl8Lo1BUnjYIhQn3yyQyu4m1mkCJVQKwuIX1UHhzZ5wgqqt1qTsnM0toiq
j/hBXUS4vrL2cdPix7EKQuWFBuqgXSnHtv0vJkJOFe1svC6RmgfAzz5e9XiO
fTYYWCtLTzCnsJDwKFtbFOx1CZbzq3gARfEUedaiIetrVqNjWIxYaLbF7I3k
1/vvN+c5f5mKqn+VeBEpMjS44Drn0H835JSg8LPMU6n05IUXR2QM35tQzVey
M5dd2lM99HwNq7PNonCHwhwXgNUIl94V0qx72l4wUPC5B5g7VNNwyrvOim9l
YH5EMQ/+ylVlQT//ZZqIv/VEoQM+ERIbYyBAYrwDiIS7rd09fzBnnmaVfo6X
ssPd6ktxKrSSPnlzx0tsQrPC1NDWCwNDSUlOWnGQ43ZtVAaTOg+RcEwxBxtV
zotDjMa1mELFLfDxbkClghtOT9EhohwQHQCH5vvrzljOb+4ChsVOi9MrWxw0
5yfaR0/c2g6v/U08KLOyON/SLM86QS09F0KfZh7c2Rhn5SGVtpsHmu1psBqX
DtOgJ9kgYyupfa5sdqciHvEBIEqXPDjzwaw2guJ+jgzwH7NpXpa8AZs1eG7E
7KWw2eliOuplAuZvSx/ZgXXXQ58HOJJ5IszAwPyY8sGDtONWHMNYfz+hItSp
tFslzyP7E2YgWLcLEI5u01wScF8yz97ANXcw+JV/odZZg6nhYtJVfOQMDypx
DPBfiINPjMkpfx1TzdcDlhWNJa85TFHCPnTLDc8oasez1vCb7Ln22lPnbiX2
kr4wEkLE5Pi8OvuHUnBK/XZpD6fLLnw3B6EJhvTI82/FZxWRXSK1QyyISxBO
BbCGHMArOzSIjpe2h4l6T/xMhb7+4c47PjXbdKplP8y5hN/zZyoEB4k7Uc0C
mD0koad7c8fUs5fGpG79SAnAJ4BRBx/2Fi5ZrsLpD2bQhrOUdnqv8xeg5/O3
h/F+1EHjHBtnLD0Y+Wuz1GSQNB3J36YnwqEYYMMWio3N+mk0wLkFJPVIQYHP
g7Y7NbJ02YRXJQodA0c1bJZbu1XWIbgJbK383qc8boXI9T+lrI58erfe4wCf
fEBOKicDHsvkVi6ewUrAx2bHbVbEzQglZ+b/3CFYsEk2be8wIz2QWgRmcB1t
L+Zh6QBa8PZETm5OQtLI7dfGn9Aux8oqwDQT9p/WSf/mB7wKhrj9cbF5ZBTO
HCmJT6XnmDcQNpUozXwL0d7NXcrUpzTTVtHiZ2qsfWlewPkZAe0JwGLCqKX9
4a99teMnscUd7MAMMtUdCAatFCJa+9rbd/5q/fmtqpS8F+r3DyoCCIW7+0NB
LQtU5t82YbDdRtFGmbJ2vVYTeqAY+jPBrGOA5h/CZI4qV0Ko384nsojZbVMS
jYdmJOIqaXGztMWH2LPhYiep1VMEk+Z35GhWa840y5kTnKl26oqlLbOD+1eJ
AGJiajXw+CFed5lqUfrGneJxz89gw1gQu1btJRgBSDYMCFzVtppzW3xT8zEa
lW5s36xXgLEH0lEdy8/2qDpvuVcZ0UgC8GDL5jiCeXiBEZgFt3S86FSQP4Xk
z1Uma0jIUKRNnTxUwHs3baWb8HlyHhhoprRazCeuKLhMa2uTFvmeLP/2YEM2
B5fiYA4aUWnyZYOfbltkMel83PyYlctzi1dsDl+2McESSAohwxDKM5/spLhx
xWWP9sMEjLDpbX5kw/Fq6wAjkARcAB8s973/GF8neJYD5nB0+DCSYOH40sUU
mC47Oti9obAn+Z3NsIhkgWuwy/TDxdJNGb8tOv258gmjmhhvEFeS+sLkJKYn
sft5o7Ib/bv/hkOQNEdxEqNAOT+mDZKitIabxOzGIl79aYt67Y8lI+bkCeqJ
0VJxDn7oAznz6wBgFpnMZpUyJL/faBttGJmVgEeT5QsKlhpb4tFdUcf4zCxc
7b2St9qCXm+tghd7bQsbtbw++F8kgp4AinnjyMYk7qx2CR94m9GFYlc2GPw1
lzFTBm9z7OkVtU3wn+VunuzFb14jHQWBPAdpklIhaEDpiVe2wMVs77YThMt2
a/UoNnPY+ID4Fn9MkMkXenzWpNyr08lteZEJcP1ndjT63gsHd8Q9DalrjcA4
Yl2S2EPqkbX7PHkYS6T+Y+aMaAu2ievSlY3Vu5xkrri3//fqScoIkk7keVlD
63qcNTk8w+v7odcMTHDBBXJrYHdOP+bWbH4LBWyIMWULPYGLtDqPEVyea2fl
gvYXMTTHyw/DPUnR7FIutAZk03Sbm+cLx/cwVTg9Rj2mf9eHarzS1/wi4Yhi
X91jcigUaNNRC3O+XXzY/uulgix4CcW8pPFUoHK3FfuvdtJU3f/xw+mAn8nr
6+6Qbz/6RO+Qbd4dai0r64CIfAEx9wlIBELgn+SeriyQ9XhEBhmG/ocqG+QO
Ye0q8JssvPfccSZe4GGTY4tuYs/9sPOOulYPOGSSETxNGtDS1CXYFOIOZtXC
DLBRL0XfYEtByes27C1o+YfaSdZBUrFxZ/6RlccbOloqR6EDjggfynvq6eEw
vs0SAIl/jCb8Mx1T+wSiB64q4MUG9k1CItQcx5+/09qH3pLptUQMEgsRpqvj
fBR/JK/aeiyNwxSFS23AZqpg3F+7LJZUMFsxfa5R/Dhh6OJjg1SBPNc+lgma
Q6m9Dgndlfh/KKH81FsLDRYyLHkKl2Eq81ISHYCpFp+R8+rNXMMMK8tBLSpd
k7fbcRIiPc+b+mdRbJJAJC1FHFddmB4pMACGasDB8FZmYqgf/mSAfIATaa7p
Hwfo/HVBhXB6Myi8M9dmxroHX71WWCxpAS3OEEtt3K8p/1DdrB+ssNZNYl0g
80UAxLHgjYTRGPUpONJv9dulfgbCFVpwJtWCpNF8PtMl/ASCOcASbi2FMs2Y
G9cklv0YMKRU1dbILVJvUZuSLagzFbzX4edOnxtqLezV3Z2R82QpA1nMYl+R
bgvD1mOH9KMWkzs+w9R/kEZOcCVd9aYdY72jyPvd4I348yOxFASDFPJD5lul
GZa1zewYnuwpQULZ9tOzwgzZwz4gdvlXv5uC9ASIyWtAJhM93lfVfEK90M2e
OabgEwTXAETinlm4fa26Xvh8X7N7hjNcEw90B13kTw8Elt248+XSd7/8YZUY
0wFYvi0ZGfQjAJgv+lXScD0wAFU71XgRAGkZkxF27AXeQjYqiVyd/JzAR6Ey
HpD1Cl3A5J4jXRNYJz1zBkjFkKFmoA8ajUz1hbjvPolZxAztn1Ew4dRi9lfy
zkHWIXLtvjeDfC3KB5bB8nwswtDOXo3YBubYxL5PyluXwv2ZHnOI7R9N8tOY
Uyh/GOMx35WO2uHbT+b0sSnI3yJhbHxKnDhQezw6wdNSHWV+m5+zFItwAV9S
7Z3EXWrafa0hY5aBO6/DGTI3TcSL8zBmlSef6XgmpKqGtil3K21NNM55Faa4
deDC4ipvSV/eT8xH70nE82WUPHhkHL9BBreVSiRFcy1Sh6CJfd0ILxteaFaN
Nf/F4Ds7o4wHhvExaDIjKkfB/cK8r/tVkBSEt0fwdwCIpLn5m+9izxMyOryt
Ih0yLMo4PfChkc+YH3JPac5HAPSKAV2Gco2p1IGJPZaYt2YegDxH4Ni1mpmf
6ccHY7DaHwGhw2qVTVD2+jlV1OihxBYMSoOUF/pcIbPo5Wvx30723u55nTs0
G4ZN97aI3Pwl0mvebfwOC3TD7XAifKEWPmaSoGhnzanJ8YmjE/SASpIWPasa
Q4GTkMoAF4t4XMjLvxsSnPRk7+g8pg1k/m4jpKfd8YUTxLbMI++bJ2FJP1QC
j7lBFuyOCD2+8iiQ3HMGduTQY/T9+HYP6d2ONB2ed1WOgYKXYxlqH5s1Tq+S
iXNkBIXbVI3IU8eeIGFdGy0VlRWOArDrapURQK3JUzbxxoyoC/g3qNJb+gEA
hLK6XE7/+3c0d2DZXHulg28oIWLBS1PM+obC9xsPkgVnyOBxv+1WL7aBocFA
qpwTgVl6YfQs6EL5PLTYi4cK7RsotkbOv/9J3FGksVbb4Po3SurbYObR4SMY
RVzim5mlSpOBOk7BtbK9eF9WY7EClp294vU9piBaNMf5ENZT64UP/RjfDJ5j
8xwb2U782Gx7pCqyarZTcEplGovXklJupSdgadr6HhFhPkTzSfjSHgrsZ7Xh
VNGXrTSBq0dmYm9v+AINKKo7UCV98DQ60St1Vflq3gFhjBJa0/64WIrrOnhz
N773kVgjeHLwTH+XuMPP/CWWN2G9wa3UiY7D+55VCGmo8DFHiiI+4aUQxVEz
C1nXnv/YQgVOE7eHlkKRT1YeaJ80E8QV+waW3drH8tCH43F1jKFD3vvwRd2Z
Rqb2l2Z8zzdFy+mZDErrnjYXbo8SlqqxiaVJwy+WYv40VJqkoMm2c8cH8nmr
XtGf4LlJQfUrYvkJCzx8Juk8GB24BF3JrkBfMdXKCSnrHg/I/regf9HtYSdU
HU3N7sWQY8xJY4U5kv8uFBtqc/m1lyG+nRT7AmWFB+Wo3/H18EFWS4vF+2Eh
vxeqpDUABg/rUDCr4s8acHSefnYvUEV0gXIb38sq8nbl0QdQ0alo0/66qBXz
cihyz4SdNSEv0Zv0g7By6u8ow2/ipXw15SsQyfWEQoJLUeS9g2bMKArCgrW/
RYpQ+Z9oLR1Yeb7gW9qszT34X6atMAiRkCiN2PAkkFjO7rrwPqUn35O7eeKp
WB8xxkb4pRgKN4XWmqUv3yqz2nFXx1syv8Vn6oG0LfcfLEpVO7gRRFXblfJg
yR0yoiZNvE+x5q4XieIRmZ9/LyFCvDau+9rYNSEDGn6Xak94rR4xwNVdZPsa
fxpYenD0rMOiQbm73v9iYt7OdjEZrSViOzJQEV6X2kZMrCCkHnW4xkRAF8Na
USYh3TmFGiG1j1K9cg5hpteltruySNLrgFw8WbRMjgtXHl/F5tgXYUJz3gQK
MecuMw6+HL+liqZ9jAaj/pD5WNVFZoGLwc7CWVeuHXONyIE2KuGzZT8Ppjxm
O4yimlumgoCsh1T6sA41u7ChS3z93QftDiBST4DjPU9Eu80aJoLULjZb8w0D
KkHj2OCwarUPVgh3xbOX/Bq507CTF1oBqxJSBzPncOwfSTfEKyoBPIk+KwfA
A/3o23+3+sA197nfAl7XNL9BeagNhQM0WVoqwRU05VHlCn85+uViIlwBv+Hx
XXETcTDVWS1Yk+YPKiKg+mEssDLI7iyeuDImVyfmP6mCbWypECDXkT4ZUtvf
Hi5FctnYAUv/Mw649KWdkh/SSE+hxo83dprvK8ly77/r17lW0x/5unho7NHK
IsiJhd7yy5jP2lj6hVmhvFTLEmMG3TC/Zgx1bZ3vC+L4EgY3S1dke4iplraP
GGHIpb4lkT+a6/LFHf0kZ3UQSQgvt4K5q/nnoDlCKrNXZLGkXHOxjdTLg3JX
LAkhBk1HNBqxdrUYUY6IqlCw7xU6BiH7bKaggZG1gV05y9v3TzYxv9UIIeo6
jOSrnMjCqTPiY9A9c+pByTfoqjzi6Gob8UQ50/Wwn3Zyfw6+QUytnZZXLAo+
er4o+KP7dcd5swwgFk7ouJZabAiEY9AktW0zwL+2uKRm6sT8E2yo+snQ+EHQ
VuakaoinfJXIWdtQb0i8/WQOfmyWeQLZ7PacsdcLq9mekeE1mcOKzTe9g8My
ZRmIAx98ThD7K99lqqbY1+ZoW0qXMsxn0IICXBkw/6zDRrzCBByiL+Wvb5gK
kt38iJQ0amtHB/d7DW2gAMOo4PSvqC29Oxk6PXGylqxhhTyL30H1ENqZuqDt
jggEqU8Nxny5mnMZCNFfHeOy5QZ5PBNUGYQPk6ywSphqgzN/nM//NxBhro0u
HcFIpfK50RTrcotSacb+vxibJJSWXZujHSBMHqwYErLQOAvmCwqQ7U7t0I87
SkCjS+U1E7CpObrxyxhIpg9Nj26VJTUF0+2Jda1IpyXQE+D7z+zFYK2mXg6r
dgsMOa0kN0C4Q3Fju1Lixa0XUDFCpWzOIWceWHZLQ0HKjxA8efqX/O+kY0Vx
6M1HqZTKpH/oahU016NQMNZylyuvuR+GVSvqGp0t6ybY0hqcsMYH5tZtkvxw
qojy3ohE4bJkmLpaOFDwWqTa+9CIGHwr4mb5F8z31cVKPEXrm+XWH/sXXHxM
PtwfDitCsPblXUy+fQlBy/INE94d1kOlLUUret5Jwph6QDKf95QhUBRLSjST
o3sOjPF7xwQ0QT4EbAd+WuN+xn76iCXf+UFMh5q9PXkimOVMsMs09ohHijGi
7NBVaG0t4Ttff5msHa7j5Zzju8DWGtzHXpGcPDr4K5bLdX1cdIHdeHxSCk9O
bepfOpdj/OhlHbM/Jjgo28YkhKXkHQo07ZuLdX+bdwvRFG8EikuzLbJvwGgN
hr4nCdPaW0kNf4lZ6JoJjjzEtL8ezYsoxk9k+67OY/c8D6rpxVYtvqXxvcwy
fQ23fNbmQmZzimIp9nwRKZXIU9ABweMB9Cyni5OEgfgDNA1fXaNtlJnahe/f
XM1GdPEZilOkMjMUjhyZ2GOEKiquFbuIqmszkDWwSyHhLn+Xz1H5xqHlYXs2
5QyAiQfcQoZHi10k1nCj4mEQwn6MUo0orOW8SpD7AaUKBaqO9hneZnpWW3cA
fjDfjLETURgiew7hqB44m1HQGSOaI3EwYJq0F3LGeMyZSZ5R7xIC97iDYCDH
mPRCXZswIMmeSDBFy9dj/8k4ezCpTyRSj9jcQZWZYwO4gS8cjjlodW8MCKOg
S6UUzXA7ZVUV4bVjUHZ7A9UxCfLIwKbBb4q+U4Jho0x3Y/giYFHJqeR/mUuu
9XTfHJVll3KK1JFJz9Vvw29wyHmGciLjYDiv6bozKHgD5pyXjLI4my7hEkAm
m3hF+fUeNF3r0qCboZOxoC4zHyeWuTzXrhYE7pJEaM2xo8kAjd8Z2jx38wyP
cIVreN2NakmtJpblYhlHoJDswpGIRPugn4GYvSikCQi7DeCPwr57+oRM8QCD
dAdsxgDSxNTn5WMwF82M37p3WdJnxDvSNKiKnulUm9eMDBmrqAyEs1PtbE3S
hPZ/ZS11tdZBbjOzaybYGq9pNqDp5MxXYmvvzwbgcioeRnHBbQOL386QkcSI
6QTs6TE2HswFfvCyEUZ4LkUEw5HvcubifX1QBtjHOfoxdBdVbOYAJkZV9IWH
rhYRJmFQ+rCaQCoGp/QVQPcHl+qt+pYVBYfiseC76qcuwzguyKFLsphylN92
FBb4bieXdKAd0U+s78Qyy93h2z+pCnciUThD2FKrQ1NMHnhprH9jfushm5jB
6vLMoWffyY8cT5Ay+ENIcoVbSK/NEJBTwuFXxRS4xrkjfrCa58MKZzxD2A7Q
Pelopnxc9TzBbQDL6KdsM7GBAB6PiFB61Mv9v5I8DJ6AsCxsna6h2D/9BPbl
1bj5duuHU7rMXqwB8QxmT7Lofx3HWrkWgVZVDUnKEWwoo++zF+uh4SNa4TsK
q3qTJ1WPpTC+lNq93D89aKVPnDP3EAXlngODQoJ0OfcIjXf6spzl/XGYwiQ8
DEpo07YPY808K/awjT/vCTx12sgQE/eUU09OdZz7rnZANbKOAb5u8FlcopAT
Y8OZO2s6ZpqIKqbz3afY7Z5PW+qPOhH9bTj7FfiZpXoDhse0KLMOGe+01MHU
vAqc9Ob7YvWUE203gO7n+nsY/LdfHjDQ+oz3QMPnfUeMUdoybIXGqUdsIcMt
AuHVKSUzXq08x5fKD0TXz3Kk5QPzAlgoy1KyVhkNYTaTfJP1a4c+mO5sexC2
rAysJ5N3TEMT1RHwuIatwWGCiWOladMzKyLWB3zKIwlt1iFo0G9ajaisJEWS
ER/uq174jSVIhC3mHuFj28eX0tCv037eXYI02XCkar9dEv6cHrRqxw6BgKZx
+yEIU4sCtKuK/0KjiyueFrRBxryPf4aOrP4Y5bwRnKav0/MlG1Qtwkqg/UNZ
svA4v61Lku5mf0KoGlXiPW+/wA4MU0IgpnvNyA6dGp1Ew6CKPwBDKxb7OoU7
ehfxS88Ifnk1G4vzWCZHw+7emjNw/e/PPvIC0WZWdqeK9och8L0kNWGtSOK9
NuBJ2h4q41ObmHYeRFCY3i4nxFsZrxrbaH+WwaIRX2OnDw8ymG6JX/GYGV/3
qUWC1HO/jJ1XWNYsrpGRFHMCHblAP4enO04ENLpGrbovIvmT8wtEKa8qChLs
EaBuVIn6dQarvXxf9+pU5Yh7XJeComSviQx7SheRyEw3ovFZQ31T8giF9BfI
s6cEHLRGvnXE+OShAD5AEO+CpCHRODZnW6ciHFq7Cdr7GmYNCslcQeEsMPWL
z1L6LEOigLz1tNCXLOPOt44gG5MR0qLyLmMj25g1yqeCyL47MKR/sqox1H5F
VP9jffnoTx4AM++6MVPPohVXHJQKfI1YtKxoFxSXlkvFxfq41DNWuwq1ww1h
CsZadAU+EQyXL/XROs1JuUKFQqUJEpG4sMV+mz3VuHZii6MJ4vHcPT57X7lP
uJG9FHv63reqnen2xTcV0M2oWk1ICjGZhpopyhNwuXF+2PPs/Wvk5SQ4HWe8
jzdJIYW4+eQhJB4JrLSBfmIgZXfOQb+p+VJHBUE93lbbe1E2RK4GBkwdwnLY
oz4UFDPB9tTdHnrrQBnoBXRNr+R89AhmWPRYQC366KF106MiGrwhW27oBf1w
32tAdjFHn+14oMcCIJlGiPE65rMIk4q/Orky45inc2ObcdXl+LL3acZECL8y
QW174h5tN7L1DkxdAOj1/D21f/czm49ofL1TGMPK6qu0zYQDhq9HZRQhvZQ9
2iNywbUcEM8uhbVTD5R/fGPsECs0k45fjZdkIrDAXt7HvVuejpnPiJCVusbL
yNNlNilmWW3XCxCX/9aaOAMoHtxdfHOGZY6aXFglhUo4C63q52XWI8WmU6gO
8XMRnx9ooSDvrQe/lUAcGUG846ZN8jnlsRzwC0e5ijVz5VkhiZ4EDqX5gjQ2
N7MGSBxkGBYtky8fdXwQEGO39yrDhNQ3q+AZyMZqMfy02aPpjNQgpco4rR5h
BV8UgZaP7EPBZsuoavNpnXsVwlUmR4DLeFa1LexY4Ve6pvAenna8nxKGmSP4
/KADEaTZom0sqLfwVZIUOmFmkqn6mgdpdxO7Z6EZU8K3HF/VCKoKApRhKxma
NyXlMkb5nI+d77VdYABO9exUWz6kGio4H6yISNyJ5bj7r3MUy+eE6X84ScS1
SDwwX+GWMagAK7ianzw8w9p0nZpoI1VS8+GMO6pR/e9pE8LvJyk5ScM8R1dF
WKWI5H2q/4Z1p41doV6XIC8Fg2defRtgLdIXsO981zfJmzUiWgDtFnTP1pyq
oUya1CBx/6CDJDyNHVcAz1IvmvVxBpo2WYqP1HV/n+vW8L7R7densyzAE3dw
fmY0j/NhDo69dx+mrHserR4815qaeXbO9QQ1slBtHgrWxZd4N2RX0Bk919YN
GK1SraOwDLaOrGeS3QPZzyT3mFaFAgSqRRxhcQ78b/OIIwBCimLEVGjuFZOT
uT3H5QZrjDxAmfgR1eaOSTXMXQ+dVyU2p7QWgeCOnwqoTGYBwZasD5FzNesS
W2Nlt9BgyFtOnQmJjmm18beBRbj1wlDhvjVSXi2Bv/4OXSX49pXMEFkzfc8m
LF2gFsqnDQvFrbwvzUDufRQfLFgBBT8WwByGrme5FCnjBbKMrMi4Cm6rjA48
RwPI8hd1ZtWMy8mZOgAXSugJnp0t3RzxA18F9q25dHxpzlY4BglH7bGlKZAt
93XTCNvbqHYdkUxWmd1WXBpZfs1yEA8vywGFOUyceK6U/1mDoqUN+4dCXecb
zotYjBo84+XHPsNL6EABaCELDDf595P0TkYd4bQ9g/FMX4THRiu6Cp7izlXo
1CB82GMlkyNORWOYE4H1+VLTu51Tn7YBzZ+TGWYITLBa/4+Mp8JtcxwRWNHl
zCJfj7DiqwNCgyKIEtgMLzQhSbuGrLAudGZkpsKRk5vjnmL6tX0xMIMF7laM
xLxX7a0DWjDG4ISg+Km2g8sTiN4YwJZEJuEuf6a7YRfTKZh3UIuj4l2ZWjjX
pYqDcTSf3sMk14C6rzSj0e7ks02Fm3ibw+2g3jgNxSRnQ6Vu1ZmuW7bXgJnF
0JRcW4bFGsE8qGk8fqVpmBJGJ3z4VQlifk/zTTs/5zdy0tjLES0Kp0Us7xc7
w2fjEvQda5OJO+jLwaxbfqDig1HkMWsmn/KrRyo8w1cvuTURZ7KY9hMXP6RY
U0/DrXOJxBmj5Y2gR4z15xw/Ty0TyYlOf6wPGsrF0vVz7JueFwYKdgahiTCr
puRMHepXOemN1iNr2+DTFp733Sf1s+LfPXR/1GH470W5VX6zVFF2XkeaJlm+
4ocRqvRPSH8ByNAp3iG/O4Gftj00jYETGKiw7m0BDzoNmq8geENkI9oOYHQ2
2BkvFLy7+/SFSoI6wlnmGZ94TpRcGG0mp4ntobH/ex6Xu3BFrQYBaMIrjhuP
OfoVQ4K4qn58qc5w3KqJkmjzYXRPzJ7pY4F5r5N0wXm2kAxlX1w9jSMIzfkg
PUGT4EIBJ6B4sUmYPcQQjUQCLz3LoUrPRMfp4S9I7e4m4rUb60Ggnd3UGu2p
kHp0zhdLXJ/HqTcsZxY/GZUGiKgkaXKZe2j/F/KQF/yAGo/P6jGlNRRzWVQI
9FijzJyuNSSr7t4/uRYZBKq37ZKh33S7zool+47gVLDSE6infDpltUIw6Smo
0bWYNS4Lh5DTI+1eIjh23pEwbVaCbDbTtupCiAAcBsnpuCZi3FEdc/6WezNC
XboDE3sM39CxHebpwamapuTLeTnHWDpVCD37FBw8npYXC/636HQ4dpLyrMcU
PWTdoEuJcwukrsf5E9yX+TdaeveLj16IIxYXnIMCjywvjDQJWYYFVU80FMdR
NJlErgdfsYM/3vpFeIR9AYu5gzIElMAGoqUPAYugsMic8Im1ANXuUdmIo90S
Xa+73a4rR2ke90vrVW6tPjkKP1UZNXTgf1Ag/IZKyvm81Bs9PySrP0E6f7jb
WpgWTtXveoIyHUQPYDUgLj1XjwmDBTgE9YIudwnlMPicP32+t4oLMWjE7sl4
dh+F4ocutR8RYkPGB972z5L5Dr5b42xNxxtWpukIOgnpfgPmPMZHCPQvMaAl
YIPfaRme8wwdsO0fFyTf6O6WH/kc7M4hC/+abyl9rzKsBlMwYiPWF7Id61A4
iXdEiN9SPzvymgXcF/E+Z7xGrvc3RaNUKfA4SSAWaNjVPt3dsFQrZZgUAfus
AiGWdTw3uCXm1uznYy96SAB8eRVVjqnXxk0cZZUu2TWQnRHnbBRlDmqwdh92
7ZF41TcAKJtEzifVtcFX7c7qvePoXfcxkXHSt81QEmeRutDR5Ee7F6Z+LYBx
5G7YdlvgidFxHOB6T4X6YIJUO1nMVUOUaNNH1Wxk/IVRw92kKmjUhJGFVfNY
uzwUrJAYtShV+i3cUU/wlH5PmAqot1Sl8R2s+dAB6zrOF5b8kWOuUiiOLqrU
b7VsQ4MTxO29WANRV1Kpo1Uj3egp8guYJhpatcUEz8bO/Rd0uvI/WLTypT8V
kpEEkeYlgqSGVsTfhTp7d3xfI+yteNIhslb41VZKBaIK6Q+NJULDBCdchSWB
hYEvCa2o+avo+uglrYGbSj4RAXZKNm4JJozW6b0STHTjk69fcDofz5G5Hymq
F8739wxqV5OaVLtNGQUcvfA1deR5h5BiGc18O3a+f9ET5SVhWnO5hSuTumDd
FR2ozpERlE7ljc7zlNGjd9BQTss+J8UsncMbvafGAMrlJarYcXg9bmbpwacg
qiGzzDz5MgFOUG64uj+ljdrYS07R948tCkbC9GJhaRHKGPEZK2sZAcTRPlyy
eWwC5jvJwGVzJFveI09JgQNXaE8gnLwxKoBZ8fcD0YmpdewstFo0dZ8atx9x
0CpNCYflD8VfG+bPrrIDlnxb6VU3CV1Zko61yRP8+6qcrr1nLrhNtfuLCcvy
V9wL2hoFsqqa9OCE+x3FVe/QnY5egCiHYCXfi8rtHEq8woNqdVevNO9Devjc
5sikvjCpH8WEuA61eK9QHnRAdnOgVbnTAvlrK2lJknqcud1iozblaHBZ7UJy
VyuUrJctJLWx5v6oOHKtzvXF8GKOdwUw2bKC+6k433spE35cktceHzhjm3bC
10YHV6qa+5UDQQ+M+Ze+/lmzVtmPTR8aIgXMWz0yVHs4i8e1w0Z04nDz8lzL
kJ2ULCOO8cDLbPM5PX5yjzMe3sBVrvGt7OR8yKJXlo+TNvZL7ogrUarS4QTz
RSJfHRnnNLOu3R0xRxJxsff23XVmZc41YxaDTJ0mKDCyNhJNpEj5OC9Q5NCv
NaVbBxL4fF2KSSF3hgGftUk9euosCZ4mjG7yECs2Xx2m23pChhSspJR7/vRR
VVH/3QOi30tfctiFhlR01gG3Am9CRJ+W7slSkEsO/FxL/pqv+WWe5D5mESgE
rtolL8ucui57Mr+5aIXNjiVVc+/kEDOQ01JHW2zB35NtashVW8jvQ4+HkpkQ
0Xnxnwk4ePWx4JLjJBhezj09xIfBzlHYWsbPQATVQb+EhmOGz16qCTcd1npq
2hldeblYPnNlu5r819Xi5gcvE2lFWFd8yT5Lgls3PY6aOKGEpFRrVJXPrU54
Z/H9pBZhaaCY738dUdsi4EAT0j79ATZYIeGmCGbXljelIrf47uSzc5qYgCd0
6/yIHw18oJokMkoDnH6hmivulmuw73mucFdWXLQlWV+q4++NRVuQHAbsX493
xO9suFCfZtilMwFfD4AznMn9sp/1latg7voyw026ZNkkkECp0AQS9R7NZWbd
rMypCo4J0HJ9pSh+aZ29XvAINJydzNsZ6Su8rTjHXaxGTcAzccP5njuJgCLC
cNWxAc+QZAnAceAC7/FPwkqSKzCbPhHDpGJOlxWY5leDIJ7Vn5ioU0XpRe4k
RbZ+J9Rp8TElLsm7lYYGbxUdaYCRrZqJKYVi3r8bmZNi0NhAfODidz9haNg6
yBuDQcjVWutuspK1nbgIGbjAr4s1JZxXFTRbanBljnAplxCoOe5/ygFuvug4
NB9sC/1cAUdX/RRvAyWvfU87rlQz7Wwnifl9segODYZcsxR02P0QBT/KULTr
bWJb/+92ws5fmtQgvSje4sokqZb63Kfohw9LIAwR8Fh/VbWkl5IptqlTtxN9
jjYj/pSzpOzUQWw+7Ti26Uij01yfD96/BTshLlBEYmIjVLBEXyIMDkvroccV
sYrYfZ2wzDiZieiKt6NwnH2SnA0Ty+if8j6E/EaZ4NO6KpYOiERw2asPK++1
HHkrt85eiQ6Da8ntgeZdub8k/Ulyhta+znRe1cei4MjzQQPm2cDq1nzX8EY6
TbR1QQxO/+xKRpY5wqramxduxCKyTrgipq/5O1gxJrXyhRStPXsk3lECZsIt
EaMAUYqioNDQw9AltRfcp7DxF0rlByILYpcw7xI6oSoNyvzpu1ucyUKGoJB9
/1dX9g4En008ARAYoo8JKDkTrSrhCsIB0DLudltkHxcpZMUmTG7yzV+u0cYE
rwGEZmS5FxsNzD9gOQRMj4W659nQu4UfJVtiVB+vqgaHQjK2gvqw6RfXgg7P
44Eyx4NVGDhASealxFTLo/CSenuEYziNhQAl05plmRsB/RZ9ac4ka0yMzO/a
3oRtNjPKgHp/vopWlqhK6wEWB8t0IwU8AvFaYqm9ghDrn7yWbfq8997xxacm
DgiZJwubbgVPvLN4l2Gllvyf/M+P6POuhXO4FL5hdVZk3wUW8rOFBAhicD2r
3yr1ZSILmqQLM37ivbsovA7Y5/SOep9DUwt3AogUllmDHA0LvOzTDZqDEjsz
WY038ftyECWRIuy6nkGGiJqh45CR0TlSD8hiZclf8yZr0mr2CidmolRRnsIs
UIyrRyTrl6DhycU2JYF4KYqHTRz6cXSDqu0lyhrl6neyfX+7vNiUWZyRLt+p
Aur5qro090PGcUg5mt4aeTs8uWMS7PuN8NKTyIJXYhaBEcTQ/jV9vmVebifk
QqxWh4MdXEGIoy8g3XaMaj8XVUwM2NdJy2Sn4mUnl5wUllKhOoU9mkT8f29U
NSCF1MUomiHgL3IqfKIAlczsNKj8wOU3zHGr5PC+v95BmJJvbHwD5py5e8TU
72npOetm0c3EJ5xaC5WMNr7KkP+3jmvcLcms3rPv6wED0AbP/b1DMLRpVz9V
FttHpkX8kTEzK1DBkjQRQG2B6VHDzKp+RSjRd9Ak3JjfNoEYXi4m4B8sLWui
Von9nA0KycrkmuJK4BfWJSjl3bI75NFRdeSCjvm10pIuAw/bKQ6nn5+y+/ZR
F0gXIMXwPXUJ6zim7EiObN8f53HYgATm1m+TvSwt7R7mdegjW5HgLQUH1Ec/
5+05Yb75XucFkVwDUlHJ0vcggNXmK34V2Jh55wH5WEToJ0FrvuPyuHIEB38l
8zAzfBeSj3hAirasYwA9+uAEcegkhzt7mexroB/mrQn0xw112CW9rLZa8Ng7
SOwT8nKB60LZl1EFqINVnVYLXCKyvBExd9o0fK9gODYJsPHujkjwP8G3KjCf
0UVqjby1183avt9Jidnpt2v0MQW6wP8itfq4VPfImPgmCbsA++TJsULuquKa
IH/Yn42PnnoZ/w/Regu9j84O59teusPRRLssD0TPj4PFwJZYaiISeTcHcUsO
duU4ycaFkij5kCaP9CN3yBsPfTfVTtsVhPFTNDf8DHglGx4FkS1cFvcwseiw
wg4j99Flj5BFchNBuz21/AcKD7oCHIWpcdsIFVcT6fyD1zWLp6kNBDGTvLkJ
FnjjI07Jg3BhH/wxcsxuqL5zCjyOcuTPFZqKztiPF/7tqnzODS4of4WWXK/i
wQkfAynF8JJ309KYPSjOs8f4WSCYpf+2pGoM58Ft3b8cL9vWZOdYkLHWmxWN
LXUNX+PGMLf9huQN4uxBBxydjGHT4JJOdn+ANpFuDJD7Dxu/KidTsFd4RuTi
avN0D2yCwjW0vsqT458KEgZ6OMmIq3S1vbWMpndRmiU/zg4HDywQfu/+zaq7
6VZKucJA116M0NFRojzDRsBmUa4MK7vsjdapslifSXaJajwlmTbmZzzvwbaJ
R8mLy0uD0cRfp1obbFYW//W7CIVzsUZp5FkDre0KxO9BhJgthbi4FGVeEYdO
V4a/iAFAMeDBN9sxTEKLoa6H7ESwXnQvX87ZQyumLe5VNAJwcXobNXPOs+ux
AsRnuyZhiPe3Yj4BC7jPY0O5FhgQgI3CyTjUo6JL/lH8RXl2JgG9KrsPSM2w
D3dfe9FcIxJlVB8ccZbMe/ajAWWWaSVedZDlIQSmPDxaSdYawtoaP4joT6ni
k6vBQcCgP/Us+KT6jU6xOy77pw0Nw8i1WSHS9mKDYyibJZnrWJ6gQ4Y79inO
U3a0j7OLjfrKvkanqQfGoMtHyQkTuJPQ+6VnqAQkbRk/oYD5b0kRv85UGASZ
FsZVuL3ycBR0Zxs8UeiptT/fXeGEYF0tYaM8FErJ6nUd1dmgiSN+ro4gtH1k
lfN06l6sgyTiwD0e6dLsAkI6nDJsjRemIMvuqlIQbGu2+b7uEbNbQufylDS2
ADT8PTq/HXWlz/6jALV1sgJb9f8Zup7Cg/KFUxeJ+ET9OnGqdae6Hz87GCr9
dyPDJHw5FhQID/haRs6W1Q4csuFeZEXPUiUTKbpdroZXBkozK9O0WgWk9mtx
JBuDix9cp8GWgASDfwQ8V9Eif4IbhCzePP2dLi3H/jsVgSTQaZPPYxmXsXqk
fL/lM3bsr5pTG8Q5AZlXbXmKeD/LSuKX4aZgBb6bQ6Tc8XI2EAQhIAOUVXU7
zewI9cD9qGSw6zK0gEBrinrEjd6IT9wklulnJUx4ihqdnyEgoHoELaIYYtrt
yHsZHPyZCNMYehd4LMJdx1fe+nEhsPX7K8QBNCrMTBcBbNyfW09dK++AX5EN
YmHGUVnLPTwI9hiEgPKjsCLwndxuI2yP37bvCbogayeBB8lerZuTOuzyIrGU
5jOwDRdwd3SXr/xaD92g+EmI/jmljihxzYRVbJ0bMs6QDxrbcEf6E7mBBna+
JG+i5rRAiksu9mIm2P8VIyh9iyEyv1za50ewEFIiFzE1wTdixzSGZ2+/YdNe
bjEtpjmJJeoINMZaEJZz9wMII8bNIiAAA/MR6xTPI2Qvrb50X2nESCWKsq+q
Zru4duIQI7rLrEbXxADX3Z2EtCdjbzYcI5nAky5VI/CmpUYQu+TwOf13wEGN
kjjc/oMwD+2HS3BFmGu6ziaejVpOeLFSM0QiTkeJZPuspkxd0Dxs9ADMmbLX
aY6DCi6SOwk5YgMFSHj9V6seSWqIcc1Ti29gWg0udSbSEfjnHFd4ka09Udm6
0nk8PFoh6nExA5JGh0XpItdOKC731NkSEiOsgY6hpxFB3nNzmkw0WD8/SMqT
lSuDn9inyS3JCD1HnDVE5TWSS7tuuo/IM9IRQxVYBQWtjVnBRPd8SrfRmrfk
Gw1FF7Ieg9JuMmE5RX6LDRoDFNuetI+bNTP+8HySpA0qtJsFMsfwTTLib7dl
se/hh4s6TGYMh0UB72xQatdGysSJrgh7QL8XkP2AmPr429n1FQbAIiogDfwf
z6GPN7dMSm6X7RuozQact1V4kvYLS3oTnG+mHXNLweg6LRokOPDzlRJUFGUb
CGkEjG4UJ593mbY+SMvdeDiJMd8UDnazPG6HG+BGHdT/eNO+JDyqR7xEENJl
VwR1iPTiDJu5apczoycBjAKw+hK8yHd6eAwdTAYLNu7270NCcWizkaQxqxLT
Mh/BWQhdVQbYC6bd1CpOm0WOxbNkOq+p+SfWilmSg5K8pRChor94okSSKSl8
ZarVAOhhY1gddiCAnMWVJP/0IgccC2AFoFWdElHo9dZ6CEqOote4P23Q3Qw3
cK27uuYg11gA/K8zCD0EHecZ9n87pQ1batuxSMe1QMO8REDfgrCmVUZM+iAl
N80dqMh7zqIPVx35YJpjEo+db6wqj9luaOBzp2e8u3a7rBAHByzw5RJgPuXp
gzVNDtF3F0hhz1pLWSNuXUMpEqQQ/Kwy2O8bJvY1sBIblXt03lW01kuGruv5
Ahl+LcoxgABNxsDL5ReQ/TpZp3qsrK8qdRVJUq6eU3JaxxJf6MXQYlqXzPR1
DVjVz3b2INzjPjPx9THby6Dup8oqcJzqTjWJiYJzijR1771BbZOBOPkMguKW
i9EOe4wWzVt0fRhNuC4l27qPV39s4Wyt0DCrOg1n+the4jYdmF2SRsh1OB6J
Q6na1d5MFGpJCW5NznEv4QJLp6B6DFDjb9lHRtzpby3SwnWiN+XEk5pOt/aE
C7TdPNk3cO8mRU0ZuiJkE439K8wfEZKxWqOvcBUI5mvfwkOioMEyRvKgWEEe
Tu2SCxBOo/xyNirkAbz+qlFiuaQ0UZagbZX6wHW9ehSUTi6sYHAADdlTW2cU
ltHEV9uolK8E7m3MWXtE77gtR5/TacOhmiAmho3c67xmdCAuo8KTkOQPavXT
OTK7moZDllGfRz/kR69AajGfROgNey6nm2zpQYxti5XaFz3HEo2dwqCaadxk
SaMpM19iu/2QxX5T9TG+8DNnWTNcHku1gR2FwWTD4U3BHONjYfgBJGDluQea
+NO+3c1spx4Vr9j6GBRhLOvN1mDI3NQFahcVyVFVPLyCgG3QNF5fr2L1es6J
3WCaXWpgPfbXDY1s8jYYlzUp3fK/f/2SRpxiW0qGIzr70PG9A8/yofxPNPAi
6N3+5triDkfHzgCLe6kz6uqujFnYFrg4eVxzN7sXx4G79TTKcXUIKI6cCgAQ
8KJo9/PH8rgUe93P+RHQazfJPyO6rZvjok0aOzsbGBwfkoxz/qnkwYtJw2Vd
WRUdBLzfOuaRfKt4uO9HiQdMZ7cGqaHx86Qyv7IpcHU0ObGioKyUZ1kV+a/y
9tfYGp7QnQay/TkoF3Jey+wMzgAxW5CtKDmjzLsuuR2wzR9ULEIT4YMRNFcD
JAmyZqpLjxd/UnFCKFL+wZstgijGXBlhlsNw62+khk5wyAHY1A4sronmQE/G
zIqUF0Yh2EyAGpZVEpB1PNLdWCqEyIO3LcxH5cCjciMR9GRxRLhK00BPqwuD
qpIkow+AwExQVd3TPs/bIZrQEXd7kjeqiC+4PnToJtfb8nQ1cZPof/Q7F/3w
Zv2s/yF7pJXZNSQ9QV8TedYx3+ghMkWym5WiNfHdXSFg3MW6LmKZdAiwP0fq
XL510Ia7bjlfSPm6PmhR7TEzCKafTLDCnfVXOD+5Z5FD+UpC9ztpPtqi9AM6
0UcxBcBk977u9ybUvovlhHyGZqDM/iCG2mdzrpyp8JvNXi5cVOBWGijnJAyD
c9WOT5FxU9Wp3RnBZInrFiYGtqUawm0vcSw1jWMzO62GRzuIsjztSXe7Cv7O
qXdaXlVWGhxEsEPvDnEAA9zbDgLkV1bcikhyh2RS2UaHx9PxLWyTCH+IQxMf
zGI/niCuvzjG01CiFVVcryWLQjl8pDVQ04D7xoVqYsg/kM+ATVPmBYN0Dn4k
HiT7884Q9Wcr3MAIp6D+1SqgsFw1wcCdxIWONN2NdLDNIf4OeAD0fKu06eQB
izqDa8YnC4zq+gY7ykgWgMa03fcTUd4RLFZsXp1+HoqtMhU1QRrYv+nwuiWV
eVuNgMIbnNZsDVPBTx8GTd0LuojfFMLKe1vE48yqTJYRNHOzB34wavpwVIvo
PlMwwxPcdr7bEEtQZ5LVXfCt/yAppQgveYcqpkOTa/k/GIVtbo9CGv02MOiK
IKPLqbYOEO5Pds+AY9Jd+/a+ujirlTpcmboZE5HQ5lQqAdUrZDHQ7DcRtEsk
pHiqCuJMbsEiFkED636Fci07Db/qmzjvKcUjkKZurD0EtFpDSJ37RYAwdPsP
jOw/vVAuaQ47utndtFWiQeEYjLsRNKzy0qT7Enu7PXimJF/AIxDZNpv7+w0s
gVCGT4fIt3AASsYBdj2R5745Dzwa42HfBnlwab8zIZnOYcCTtyX8HB3lFE4C
xBt3YEjELRsV2cog1YAyUUmASwtAzVdzCz3+4gzNUafflO5KwtMtY0/midSr
ZBdgR4UoD3SihQXnUm5fQ5J5vbcQTFXBbPYCWf3zmuSzgWD735nDw+2+5Dpj
+VKMaZBhH8bv0ddk3zyUKSVjEz143l4RlE+WmiuK/2mBNmkGIxg+004ZzUAi
dMexQMImf7rm8axeJLAX+YK37+U4BONQtPijtd0Fzz7Lh1o379RK8Rjb4/vh
MZQGnulMGiR6Aa3t+TT04mrB2fJ7DRTFLXD5GXTG1cchO7P0OSWtcVt/VYYj
J3RBnyyeLbulFFyuClu0q4z1MXUc2zYJq17OnoNWI1bIYM/xZQhQkJoTb5ip
CFsq9bR9rDIhOG4ye0XhX2gggBXpeb5KabL264vkIfG81P5hXnoK8wHBmrF1
n52jyNeGinK1PQG24jkdIFyKzGfymC88AcDswKnH1BQZiHvXHE2QfHp+r9pL
6ZDtfDu3lfVutGQH3OTYwep/vLJGGi7XxhI6LToc6rT+zsEigK/krxgmdozY
or5kclXwSZN7u0iqafDp43pgQNAJn9+2OSYtdudD2Y2zCSydbu4DHvlxuAN3
V1w1pN6ed2EwfJXT1wAXph5Sc+VXUyoIaz0TLWLok+BOTPJFFgf4ZtpWIOML
HhxhTs7FHk2iThAsxusPe4QiBUeWuOCKbCzu/zATLEFghJoBVmNSfBgeTp7Y
Oa/6/Y1NUAe4o9poAvXQS1/tWRgpgshWnFLkfgicCXwzYbb3mFjsaVHIlC9F
MrmInMzVJw53gaKy28bhKZURxyzX0azcxAv6NovwBlykSqTxtQDJfO5Uh4b2
1ovFHn+f6SHSQo/tHKbCoh8MpcibtMdELDxwyJK9k5A8txk2gnBYzgM+QY47
pgnIzQY0c9240lNSLlWsET5gV22TQUFkIfeqzor/2RJv1cqpJDRJOJTbFQnQ
5U7mGyQ2Hsm7NghGuvWvJKf2Tpukt7UF0hss6CRWquvSUgjc6ZVbGQD9u78y
9a7u1OwoQlwpKBvRL4wKNHXJx8WxhuBma06jwcf2FQi4NSD8m3TBtba8aTdA
PN18jAgd6Ts6UAxPKUZTQLovSSPSAhiC+XOJuh8L2u+QPhBLbRj8zkCBKOrz
yauuOJzqI6EC+yK9tmXO5SKwLNQAPrR847uH1xiJsoOqKw6lPAGzxLWIbtd3
RJwgSRvcV7RAwnbo7G1xGSiZrvUI+Q/tnkgJoLXgd+ZCcPaupP2Uo73SiQaC
kfNN7EkqDK4icmsJQ7zVuzRYY2Xqr7vnAhSdiHP/bSURAd0jwOr1S14kC+FC
kALjB/hw1AwdktAd1SYRiWcsdFpytpr8ko+CXrpyh6bl5kMjjdcgTr0h89mQ
NFyoicOphHzf145QUBqdAP+fxr88uqnROzkZFZa6eC699lEnWXhSKuTD6AnO
m8VTv4EW9AKi1v4tWuUzWCqBbrAy8tPlxp096GtOeYZX3DFLBjwJXt9+jms7
Z3jiEmpEYeNjM3X/C2Gpy5zXN3+9RgS8AIkWKf4sDoOKBKqd4feW5+7NCfwZ
F5sQmeVQgE+5AN9s/bqR6/xFMyYrD2cy1i0vWWTomVIh+Cg8YwRcGAZbPU7f
3hhCDOsgXjiDkbghlgBdDN6mDX++84IyiEVFzdAdvMdRjb/yISlSEQu+8b1o
UeWbIh6Ovp534k+sLQm6VaNkHF+6Jrumei7Wz/Qeve9GJn5Xrp0SDFAYedDV
pWra6L9UjWIa9Vfmhc4UqgxjxET4oNC9m4gAd451G03Dx2SJOlPdnh3uTPv2
N4UtTthvC4N3AMIlM6hPD3srgGsAC5tmkBLq3C/POVTQKSG2wsu4TVsKpoeH
8wwpsJzBJQ4WHZO8oXMkeTKGmAWR5RXtZTIxI6KLjMigzcg4Nc6Xgf4fKzAO
K1Cs6ruUghGpK4WGxYiH9BMy3/TmNtJXeLusolloNBHsizm1gvq7YExQsecz
atm4DW1leZ7/X3+vFiXyc+QvpUY47b0+vvWq9YW+g7ogJkskZI+08SXSthiX
7otxExuBVPt+aCBeyMINqXyqN3yI53owaKRmrD9gIUrQ42f2xWKeM3WiSt8l
pn9E5t9wcC2pU5SXEaDlm2Vmn0U4MpUP0ByrplxQJQO9PewyRpSn2csMQm6H
V3PEmxcLUUBmnQxRbQgxczJFHP0QF4Bruy0JmW2YlRy9Cw+usSQabjYE9nKf
GOP5JDNpBc9IzgwsmOPkVO9NxxWeg7wCMINNbMay0rtn17kLOT/qTbS2jl7D
1F/+DP1P0nhNMOzRa2vmVr6992gfUoUi1BZTCN9JU2qBZYs3ImXHUbjaV5YZ
QxgARaFEt9fCyxKRlR2Mwxq0mBVfk5EkBrljr2SQbLHOETlHYIuxThNqNRBo
3tmG7qYmoGY/wm4gHnvWBtpWNI96XiuZqmUSP/Y/PBuAi2GlOZT4TkG6QfIy
rkPXWCebSCE6Uq93LDGlyfu8jyFJsHPdoI/mGy3/ajsPGOosPQ9CoA9izOLK
oJ26h53m9ds+35DE8oHiGVXNtdkMoiDlEMf2AoO4h/WhO0AjjoaGuiZoz+rL
95TGTiCOUyVREpZxH40Wj2S2eBwvKXvcJMi6HM7KbiZIMxk71WKxrNQnN/s2
jq9xzkiTzw+Fc6+Wq9ineC04niiToF5srQCbjalG107DXFIVsEWWOa3pujXy
tRgwvOpIqXVkev7ZOxHrCiHMZVNYvvWXX2XRD1oarmXiDL/BoIyrx+WIk5UT
84V2GqaW5R3vn9duFa2ZCBzfxvW2tauGjJ6WrwTEzUhEyJCAJuypnenWx/fZ
U+sb2NKWzC/NrebnZGERmLpdua2N+8arKYee363Bn8OrPcLwpu1zxdWMDwzj
w6nVMYeAbTXo6bzs8RINFWuZYtzLB68n7iIvnl2so8hnS3juxWTtqxazd8Cu
TITZascPFKfCCkWbkJ3sGJFJ3VmeWL3mzRtIKMtX6teGEO3KpYHRL/4f+6lq
XFi4IJoNqGjzZ80v8JLuWdHAzY3OE24VAkh9FYkoc4PoMksFgWWPkSv0JoSo
2xwXmXwekhlcliXqzjd02BTeXsY4eebBDkdRPZhopyEDXo7gPqc77OeM6LGv
QVSvCfUZPko7IpT95JzkhmTAAc6K8V+HPsB6gkjlVebaHDcWt/N+0dDqnO1f
mjQUTPDF/qI3bdUZ+QiV9NxwNI9wz9QkNPCZUpsueC/3x2L2xR3vgtvU6ZlN
Q6FqVCuJtNu26d9rJtNdi/kThWXOpR0NtcB2oMSqLssRXd6WdApawjpY7rko
WDMkDyon5JJVHY738Z6pH/Frj0ONEQbT+qefLJp/UYpyzLfcAMi2RuBGwZ6b
d0aqCSQ0x11Jp+hEqI/S4umDJlJAYHOwNpoQMziJeg9UzSmUUVntOv0pVp+9
09c4VCKX/Lv6PmNFbpFNLEX+6CyzjPPzJc3v8J9qGPQYx0HHevz3xBI569VV
P4ac6+orc51hByOErcm7y9UyERQQc1N/7Z3vshutWLxziQDEBW33O9O9Vl6V
gDAqMbjDCjSrWNk3yBOsYzu65EASWCJCq8/PN6rASeaLCziompbCjQ7iWBQs
kNRLK8l24LFJHwgN8AxUa6xBDI64+MateBnrKr7tJdW83SKGX8kAU/Y76m1y
Vu37xMNgw/n9J1HCfVPrlvc9cx5EptQeMa2fqg+ZHFqThAdW8F4cPVBDzY3W
DiUA+h7q09J2wDcifbzOyfIjBJz0WEJ1zhwTpLeOaPgxh3u9fqyeYUpNgi26
7+WK/GNB+UmuNl7TxrSQ1Z51thSJgDl4iI8X8KJ5o9/UPly+O3QTEuB+vF7I
XzlESCBwBuooMU3R8OHa2kiXUjSP+RhNUVzActXvEfVIMl00fTgaT+LcZwRu
aNllf4n4DC3PK7EJXnj/4BIgFco6vqgIpT4LuVNkx/F1pAHZK8JYCwPxvenD
2+FYJnpXE4H6VyqXolA555qOpPyhxpSxYacLJYiaYKKq+1/BfwFHQZp8Chpx
WDPI0xGYqJMETg4hUGyAPUXlhX+vwPYoJbBSTMtKQqZ8q7lpEfQnjIFJ8OXO
I+Y1D0UzaOcD6tYubqwd5Pc6AhOs++Rl1iM3iI1AqtoShvweNEVIfIvgjl67
xAEeAvkyvE/+412mozem1h9smBHgobJDquChB+n/ViIF60A96TmfJ/M4e9VY
d2g6mnH6D3JjGGSFA+Ewr/41M/DAPO8pd0NlNl6OlOok6MvfzJBsagtx+NDG
L5aEc2+XpAPGfXgZV9TSdIcIidGiA3PAuTSf1H7Tf8t+JOP40RlF3htF4dKR
OW5yej6sMRuKa6R9eio947BDWJYF444n9KxNaeGqPjMHRHdSMAvgFDQ9QwDj
/uvZ/aS/mgLLu79pKkiANMv4wr4eBUb4bG8wdL3ywia+omNXDyFbveRPC9MP
6+2XbDyn5FFUsWa233MbMX+xb9wKP6oyFgOt3mremqLPINfHl+Le/6YuhfK1
URYg76PaubhHdloKfZEJqURNo4MBJ2IzLBNAoFeVU9j7+X0bDCqi32Z9dGTA
+tu5thQitoJXdR9sf4bRT/7slYJIonaSH5soeLsFYlAzSBMy/QQWPSB4+Vb4
NWhiB14nf9DOk6LBju8upspTw3JsZsezI1EJmzIfYv/nFJOVf3ncacqWeFVU
OvWpjsI9ZdOGVvipC/KhXV4XZT3xnzHbae5w5VS6kTYXRKsaKj2F5Ifl3XKU
S75mOXTrbMfEAidS3Q6m08Sh3YKNNXblv61s0OYyF/4CHuGgE5hQWpyDxYHt
j+6octVEEF0fy48RXXieBcDCz9YZfqWjh8E1RqxyQK+bG7IQN5EZFnHPCpDq
lmB27yT1bv4sE22ud0hRctMgBWgnK5Ox8qwhPQ6b2rBR8z7DO3zsVara6Yfd
imPiJkXrAWhex7DU8au5ahrlegjbr8DwtmPMtLnLorlCXk8NfYprnVhCcAzM
DSmXlta+RX1k36mNL0778HyShws/djl/6Igu5T80Jf76neTynFJejiGbJvX4
s5ipRBuTyKAgXd8OFArjAP/FTz8XMzA4wrH4EcDq8xhTX6tsyAArR4QxzMmi
MpWc7mg0MCKqDX8zfYpbSBPPutHAJDWEWPkzXHnjzF4WsdYRPIAWexS/s/Xa
LMM/YMviXThpMm+7L+OV4osncaRJUhOmsQ6HXHuBV7kimZI0wqzNu4wyzNdk
CxChEKUew6nvMK1xbsuN36sIx6YvI5HD4KmLPfvml9qMLGz4NQLe5sX3AYnZ
+7mOyMELF1dVaEJQbuAGmM4R2JrKFlIvnobYJWPh0ZrKGBgbyS7CfySyb5QJ
DBKQa7dClJzrUF29vwqJneo0/o/dFEnTA6uy2GJ1FtRhdM24o1+eZS4pZ9iS
c5LjPfevNngzNVfW+WIl+OJo1ayT4ADm2e2c49lbiFPYH/+T8DCAYqyvbsBE
PA7dhKD3ZDmKlpsQqOiN6WHDjqpIIbrrqIW7GMqFqMI6aARKkoGEmikL8DlF
PeUz8Rip9qOTtPVbcVnYZNwubq/+WosA8C34HXhf4r7j5qesJ4NB8K6QXGyX
Evk4iW+LSQeflXZ4/vGrKCSfW8/Nf31XtFag0hZ1OheHtXZe8ddz9V5WcNti
2GwElOfRBdUrP8d/ePWjx3vbE6PMzO5j2+40ZeLC1l1uDGTRp5qPCE2GZY5v
emI5k30dbpaH/sOyUSEeqO4+pjMCAWaoQDuXDENFJIiJA7wFJ6XSo6irhbma
MwIHGI6aDCp1cFw4kFZq2ju0j2qc4Jfbvup1GII4RPmAq4Oh39mIDLhxJ2rK
8iEEAYKSnSFgdFn3UXexHrSEIDWa53yxcVHm0wZdmlG4jj3clBPXERxh4a4d
Ak8DtIbVurB5Bd1hlWcQQpLCahtT093YDSm56WzOQTBJWGWMHEffkNmuIF4O
dw7EUULGmjyl0U0/huAM66gH2beAifjZTyJ9/QDcBMBjI39iK7UcyfiL/bym
9QsFowkVFA2gBLSRKUwE2LltBpTqygaXu4A21TyyAq10A7QdGF3oZbLPez/5
qP/PfmTXXk0L0tdDcmH0HBqX1UayfJf95t1vuWO6dHv4F7jImiDBV1BKUIyl
EfvRWHGfkYJizc4xNh91gAQt2zElA6Lbze12/Msw0tidBCiOJMEzecg4P7Ee
eG8xPRswM1KglW6OW/4+fK7j9+s6OVKMTWHAefev8RHt4nj66qU7eQzq83EU
BtWkUpyXLx+tDz/r9rr/ejUIfNUqz45GCg2KIDpKoPLjmSgVefZkUNaMotu3
kYCVJwxdoOUdl+wv7zNjbNhkhU3rJ5EUr4TCbsACh19yWoj8USwy3AdyGKWM
adol0eSdAYHB0HLQxJ53aEUyIPUNCYqodYVhnomemgeq/gBGmH/cKNKQzqIl
+WjGuUAsUgXb2UjalyOhaHWUywcpJuy4eHg8XdvVZR+chtY7rpMt4NELChyA
pXbZfD2e9EkacZDHRhGWdkDyvWbEdILq25xVFpgS6noXmH6sBPiq2eova4TA
cPyBGqYRE1pIfyBa0z66+/PTD4lCsEMu0AQL1bE3ocEAZzsAj/HKQwc4g32P
FlF3vp2fBOl/1DT14CbXczkZN3V+bqUmr9fyvURRQHpX5eba1JLwyc7pMdDB
mub+fTff/NQ6f4KrlJK+U5a7OKT7DSnzlhUPvon5XkjCa7pol/8B4G5l5xiV
Wf9xr5LD7l2N43KJMXd8N/gwNaxQiHiVMaoasYzO3HkQQ5I+2UEQZMjCDoxS
Rn2JXEzXPSAnxEFbVdQTjLwqx1VjU1XevF0Uajmf8Pr1TwpmBNZk9MU8Nv0J
0OU5SEM7ugOqip6z4EOtsUcCb1WYUEOoblCaeWStdCIdJ9XDOyqOsWyZVdYD
FLGGcIj2dC8MYmsTaqeZ0qKkP0kYtgS6BnQsuIQzDIc1qM9VEs+TA8gNMqxL
QG9u0vhAZJdLjUnUPiJ4PqTBByJAU/8uPjrJRb1ZENrkyxDXCkxxJagmj1PT
WbT/4zv2/QjjXcZc0IVGGKxKImVEMkERWzIoAjm9Hq4K2iBTOnMly6QKC2YA
QaCIBnX8juu/pFRdYlxO1SHw08w5ze45NpNh3HMvijpSyuneBN5qAIk71mVT
AzVD1eUr1jKtfbgrIKdg5AkfHtaC8czZwlb24xBjsMO1ti19zAw8TgninGrx
63jIF6YkhFqN0kUSXdw3cuLcgNxCqokgJ5Ajnpr49s13EGox4LnZY2NvybE4
EFMOy10RLeYmVCeIfeF3DsH51zXmb1rmILGIsICjeL8UuLSuzkdjSR/luezZ
ZfAugEDqpERuZ3pU/T+EKO4ONjR4RW8HU0LakQ4evKaSpQrc3px509hZ6Gx/
N4z2C+5tLsQ3WEcrpVj2KfAYEeOLXYN853nuJg7EJWcrA1KWqauLjUBztq/A
6J6dlWstXtxiN9c328Ob9GmtHmTwxh9ZwVGJB9zD2qfxkbh2zDlTW41UZNw2
TbUTve2j/gP9GlMZ0k3X/wrFF9dj/zGYEsTa4HfwWa1JHN3OORHUkBdXJE5Q
1MImNXB5HZxPj8/Luwok55kUrqL4NUVxtgB34RIWaC8Xi/GXE/Ij7CugW9aC
ErXilfnvqyd8zpPjf7OEnWdvPi2mIHM4YDbWir2jK+H5QmWLKxXdzxm9E34u
bZqXbHUw3HIwvDNUIhLfIEyAj6ISGXWlvXOK0QwbTvj9riEZSDAdSSKSW9U+
ZBaF+YvfOKHed6mfOF1WYKsFNGNi20IPDA4OE2S3WgcBVxjZ6N/oMHO+ebrG
npUXVVqsTBiQt+LTs2pSW4IHRVFlCfYpPRXyR1cpZ4tehiTNN5IOHuX0Vec8
K9qQ1YryMLUt88KPeyB6O2dU1Q+s2L+tYaXB7qSKgTg2OMOrepHVb/mscCRZ
PRYUeTE8DC9lOFPHn2po0tdh/U+xCWIOrHBQBhqUwOF+2FMdDWBc8/r+vRkW
/Bao7S3RQR69GqUt9PfHvesDd5/hmyRfRU6CqN4D8ZOR6mGxIJI4xaCu5rjQ
QTDeXIvWVpTnAZTBIvVMIDQtHNq3QYS245p5NFci5N2UjyVwZQen80q36vYX
yR8ResjzSnZ4DV9Gw5ikkZc9zj2PUWKqWFXwnx7HmHl6CNwF+aaDHIQoQ6Zs
dgICvGgzAu1Dwg7zvwxjM4rCsrDGAC7kSruOnIaXCh1q+MnwyGDqDAKv5Xfb
q2Z6l3mptskeT+zzBwQ5XFW74EM6N5VsTjFvT4IBLTBsxY484+Xln4Pepi66
m8ka1VmK1D28k9AAgreVJa2MyLH3GMZ8+OJa9HSYB9cOPQol86U6xIFzgV03
2sl6v9xZw3tTlT7a+bQ/SCHGuBg6eko7zyojz1ahYGbh7SGSFPJw1C1BYbYt
QCU/CV1SBRTJ0CCBX0Fd6z5cy7E1giGN9t0Zgzq3eUCe2Tt2OniEQL8MUclD
1suUkqrc8Xt7ZS4I0aGGrpDaYLM4wqyjAh/at9IBfZ3NyK78UuHI+BW3QjPQ
CXoA5R0ceOgQjcp0wUJSCxyTf3t9htnLvK6/L3CII1mBv/qx9fFamQKAtSuh
pVD8qepOCSDPjSltEX04nvOPLertJK6b/8VO2NJhqgOo3I1yETkCLJnci7di
m8fagXg+NlKnhOxyroGtiBOUdWSa4MFZ84KokMFcMVpMTRjJg/+lUgR/n55J
qC+0IZD+QXwur8xQJz+y1owxFCfsX/74vzka6qtq8nfNfAgPFnY2X80lN0ut
l+IeYwowyJGSrbQl34nZTcyi0OzJ/oJdL2ls/4fZ4u1aDDdgmzaFUkxweMWa
nNzOChuyQuLew1JiFxyuebDtkgT98nDjt8VjxRl9YjhcHlQdzCWnsXT0cFiS
wHZDfDLX6E2u+7cuw44LFJwhScDdF0A9QLLVZk8qwrZlR0+7MP85hzhJsEeB
J1y75OnMqEy0PwWhHojvlYSMqhSQAps4qZd+730KsGrkRot3iL95qrt42p/j
Xwd/9l0eH3p2iBvhm+BRmTKBwXseTowc00hbkZ4Jyu/3NoLrYoEuI5G6NG8J
UjJrfXL/AM6kRQgi//nAIt9PEXpeOquPBNII3s2pZQp+FPPfZm6eQriVrRS8
CsiYk6Nmw3x0S0u8BUVQcnj+AJpEBEtmvT5kem3MU8mH51RtvJqq+SMu00RK
800gaGTbhNIzRD5nubdXAcvnGItCDifmHDvdIl6tBTJ7qhLWdFHoTec+aJMu
/lIQRiOGd2WWpUGDSxGeiTIXqzM3SJ9JNb14bDfw8WaiaJkKFI1rEjmZcmJo
XF1VCHPrAY780PBwJ3FyqRG5XxCJlzqAAId3STea48xEPRhIxfvFZiWu87SZ
tNQXhBkHCx7QLUJ7yprt4XzLcHuFRSYO43EbrjfU2eirC8BDgOZ6MrmfArcJ
/BfoEJX9RVOpgengey0TEA240JXm028s+49fEPhwndL/OW5+1fjx6pNwGyAm
C46URhrJsaJwRQdX87Vb4Ngv24bu8pncltO8cpHFGs4DlBt+uUj7ycyZZ44a
MFWcmYGzruO2p6vQ7ixLtrPCDpJM1Dr3pude6VXptk0tv5amcc6DUpk8McTo
DaMzFsv80KWXTK61NQzVixTlx8gd2jGX5Xum5ewZqE/yGdC/K2TkjK0IsgDh
jQt7l0YpIOkooiOwMyXlf/bCGmd4KWg6+X1RDS7asf6NDMqgKn28I8a7PSmD
ZQcPF+Kj5h6NIZYMvLboObf2Qv7XKao2SLbagePtdvWTQu0DpectBEy7wMTj
QEHecAilIdL1JwnW9jW88CLYd5RjBX8WPQt5S7R39rA1x4dnC/fwVEdR5oZG
FzeQ8A5Yj2Rxe/kj2LANB5PjtK3/vGWWz7m7b5lA+gcN5dNg/uls7VLQMdhC
/F3NqOdzrg32/24SpdQpY5aHFxR2XfpN81/RhSEtzRJSemIGAVZ289RBUOvC
PWT3LJ6eo5C5gyA7ytSeOlcTmfxuRHRanUQAcfdGqoklTZMFtp3ExOGIuGuW
DawzJ4ILIelyy+NWw6HFjCI+rvobWrBuDXEQ5Wie45KRuaO0FbGBox++Ngoq
SW2oSOBhmscGfCcqQCE4Ok9ntU0SGAgBlb61MJizxge+cw94fMi5VcTCxBbM
Jo3YnkDxIRYkHkCYpOIs3DixgADw7T+Ef7/csriErJX7T6bBjn8yhfYLzdKb
hZaenuEbZjAaCCImHTO4KQJ3ac4CrU8Pjxe3/IgCBijMndjFL0GYiYxyBaOV
e/djXV2BludxA0walS/IL4mZFvYYEKy4P09ZB8k/OnnDjiRDA30XDY8Qkm5g
us6G2YPOpfKydpXa9CmmVlkzhiY183TD8BFE6yE04Gkp3Hv9fC6AeT6GpgP1
vUesOgXkZ0pUVcM07WxTm35+5L6GCVu1IHXO1//yWV1HF5kzCWGa7+7eRhc3
VBFZ88j1+/VhgEw2AQCdkNnIzZPuJ18uu+5YXQDNsacqgZDg9R4vF/jojSEP
f5KuYzKNw8d9NuB1k7EkwM0597COGVeYpVliePtQbqcJXrCD/hDKIF8+LNSN
uYEjDFIOYgklXQ8v5irANO+Nnx3GoMAhKIASRbrP5OZPRDIm0v7JNFLk1EW2
VoOVObF5YFqrNlaMMLqNB/dN6qOedCGvQgCUboeEanLBnXfNsMfvya8cMX3I
6JpVqCbKKybqZYLa3zDjy1qRzIfMU6OYENEQgH5vL7jwAhCkDqIHw/pqLoGs
NHFYxHoMgd0o5c5vzcVlUoKmiY6/xqwkEg2G+wu+k2msR1Qngn3i0JJzLeSA
Ud4DUHBR2WsLm2P1VmT3p99CJE4Nj5DzMfGWWjCMJmYXfQ7zQ1JBasjNe0/K
FBvIyiy4c4G0OMVMr6lEot/YrkABXPjlD/+wjg4E60klfaH12+LzYmZMM1m4
lmhGi053jl/rzy8O3FZpwy8vp/RGrQ7e/gG8u1da39n2Ct6hkiyfQctj7IoU
7I5Dro3TuZZx03dtJwpbT9FRovnWxpe04eTI1nuZsjg+cEwxA7uECKRt//+j
I0lvmroT/oLyfBp0Hniykm8RzOLqz/JRgarpmI3bPk+ZVLZY/iqy9iTznYKn
l4rOvGNS4dyIYjY+TssgHbwpnMfm3sFN4IlVi3XFeJsegnGUp0LQAKH9NKyz
AbYsgOYoAGdaoK6twK9QFBcU3KIKpBcDgn0QqHgcGS3w22SVL7bRuIe5JBRI
2UWGk/tV7DdV6bBL9u0+UlnVEyi/0kLQ8GujgU3dWsWvXYs0MvcBsc4Xl7ly
PkY4ZkGF15STtPUo8aSXzP8/cZc5Xk9y6wsolOxiARTiK8BWA5y3Ww6JDk+J
l1WD2cKcoBJoPvO+xoOCnrwYVqNgS108CyLvGmGd73+DBP2Ef4YZL2r57yKb
VwfsCQyr+lxnuIFcYzzx6tMdn6cVnPM4SDQC9aYkX0qKdEQjLkAkTGS87A14
oj/PeHYs+G8jvBco4TVkQcEy8YAu08AmJkPdVabQM5SwX+QO6Z7Z/EnyPMuq
ucnoGu8eM1cg2tbwznv21ra3I6uIrtMLTZm0jV6cufCwcY/T8VpELHtc8kWr
NUUogafJT+zFtK/q38zADKsjLUPAfpPQJ1cdbY28XAP3fzPiMZ0ZJzph0weo
Xm5KhIaBKVe5/uFhf4Q5Rmmw0FURN24svfZIIAsyZNEjuws6Eve8vpXlw2hP
YiYiZ9GwIfBS6z/0CEWggnrOYn+kS0G0hN5SZ7nE566ts8NdE62Lk6FDEooz
DqqGWLKHQVTDMgOVEXfpO6vayF8Io7jRve2JBtyUM+ErZcM3KvjGavMZKMj3
6eD6uQoreqaWU7N6EllLUBqZx0sjk7tmyYLSvgFCOsh3sXCsD+63oX0qBoWX
3sF7ns85O+WXqFBRCP0VUADpgz1GnXR6LiEOPDdod0YzbItGn2P5FZ5JG4K+
A4DooJjBo7Q66SE8iqgwZY4OZmgz10NeDXfHOKwqOeLs6swQ14pN5SE+wOZt
YnOGKuqkoLrE377skZ5oAEKaMPDR4Qyk1vfpn++1z2p32O6VTWO4921IcLkR
7yNnqTbBcL+w7Fz4JK5T36S38yrDxR2Yncfsa1PGp51CGTNTatjdk8k1mq1s
FavSQL/vKp/JSUCxRT8LDYeUMDZ/e5Vw9DOfhnK0InUBySOyAxD+SMI1g4IV
tMNdbyg5X9VmR573CS2+ZPaBTDJmj09hnGriMq4Y7sm1SH6EdIs6uf68QtaD
0EAVRrfOBCBj/c2e+X/oLheUji97XDSA50uuBCfwQ8dbyJuexMnEOr/ZyEQa
hIduQos4SRjbtZGvRqpK/sNHKvsGdYC5Jwt4/mqJjI7Re77aqPo89YQ6mf00
3vvDKLzSmuOaptwMPJM2eZyS2fJyMwtVC05ML/iFgqhDCHs2UmRME60uNwsl
47mb2geFqi73RWYNZ56AT0hLmksgjN4hFQXGziHHIP3m0bmJYtiCkr5Wt80a
cY15XVQQmWai1/nO/xkNNR/wHV1IgNrWIezU27Vcf0ECgOaBAhTj5DO5/pTB
Up216bYyIjCXkKeKCPvWc4Xw8qr9Fm2Sp9t5lYWxIoBBxd0ReuGTZzrjAFoP
oWNFn59Iw6HrQ0IQaW+cbzJ0OGzUrE1bGN/ZYCt/K6YvWrF35ZwjwN0Xbhib
i+9p5V1EUoQbWz4+tZ5elhxH/M22Fur52zgjyFL8AJj43ihXFhdiWyBWRFGJ
evcb9RYsuKdHuBfpxS8e8uGfryUCamX0HMznH1lUhfAQkH2nKyl0dX+MgHPz
ZFpBT56YHBzUsEcBCgxkVMdOHIHOrJlyxVqquHBNv4CwwYW/oD6HjbF0XH2l
Ck8YstaNyyIaXXAPNnufR8Q4PrM3GgBQuCVSHCkK70MYrt2DEliAK7xEmfYM
nhgJe6LjSszG7A+JeIHs7DtNag8dKNWhi2ROXnaD+cvCF5QU/GkE2dRGhW1l
mam2dP6PeCAm7BniZ9/kM7UarqwyEsyhoPA9mbAvTpzA4hSRUn7N5Srs4aA1
wSdg61lt0x6lTk9mRUQxvueBUX+L+C09StCnJu24m5u/K72yZsLmCJDvR97f
68j14CS36c9qxxU4lyfPQhRP5L6+rPs2ha34yycl6o2pbSDpahUwToEgG8jY
gZ9+3VgnOsh8BdBWJhpaqc27XWegLLFqrW9CTqSnwlkwtAgDamjiU7NCGXjS
uwZLQb6FaC5IlQ7GlDZ2kgdj9uvL2qh4HDTPdCZyRc+1ZoORO4W6PZF/cbtV
KqEV5UNYFBu8hE6M88Cn5XodM50aIWBj5MDTWEl749T2z3aQ728K7QMX6kU3
zUI3XfWVNFNM6zsxkEM19KReszlYqXAa5RqXbZwRmZ7TO0vRPwN2iwss3A2/
JyAbvCln6Jy7D8efOQnRsuI1xrpkb6EWDmKxFdnZdmTR4k0kxY6v1vd1oRoN
ytiX28GgorOyvfz2DiS5DrA2qKqBeimW5sK4ZzGnkC5wvAdBZF0BXjigUzYR
c0YcQgrbbqszxRrGxsjTfkz8+eT8DQZk6naGqXAdetgqvwYG/U/aNnVp7jQ0
hWtgCOn1DRGhdPFTWaZYRQ74CLPiOtSjr9qku68fPlfwEzOfSkfwIrbwuIkg
ls9b1l20t0+YoRVJwRVU1M45dqTg9NlFz/PM30YsUXZQoXZYuJY8jgPEz66m
dD/LGNvGrTLVnH/82s1iayrUKVCDRhaguxTZkTyPL/vAOtAntYKBhZb7hY3v
x8PZUzuCtEcgRiInORrcnVJm9JOIsl6XkqN64hwhJKLlR6XiLpAa//CTXnP1
PogzmkN3OLerhrxOcHvvAKlNsg8Tr7LtmuJguQcRPzqfkmqGBtpybZMC3nxH
mz/jjHndts/VA4oChJK/Q77EJSzZML3oFM6+2eJCijE1ibabPaDSVU/K4MQq
fc2fclzbQ0EOKnRwxyVwcwpPOFrj4YIGTaC2/OfV9ivZypCCIU/gb0DQ1jc9
t388teOyncFufE0WzaWgjDmGkmx95wmcRZwBnghqZuKltc2Zly4uueqKepBA
YwHPZh+MLxYOYej1B+xYtzUAOsUSoqJ3wPlvoOsdhWxKtpcaCe6ObLR65G57
ccwdKAe2m6OcSOUfA9i5vpzw5kR6vntQ5b+EQdFpUYSGL5KTBzKJCErKVL77
qi5rIqWutflJ3C0DHLnACXIVqAWVNMOQ2ushspCwq2FvbmhiRNbglCtaYgSC
3id77hP5vVBlZyBSEs7hRTf/oyyhfcSYPC+KydP/6PheEq0lv2lWOrozcd5I
BwjMVLhfR2tfMb/hGtY7Mzgk7JrjJH5/lrb2AIcs9pn/TZFNHunTZkpSRb1R
tCWHSQ0rUFfAouNUovQHDCmYJibeFLN7XiZC6C20f86upw+qnQBH8jg57Y3F
UFRQwhTAXjjLJizoDs2MuL5lJfM6hpwIuY9eirqLClw1M4hxFJmllRaPIG2Q
anyw/PK0eacs8SjuRYZt8OfbLLQEfGPoYymOqfWdG73sfc+NXlCsGoMXhnRa
zATTX59NzuiN/gOaBI10DuKMfRwXRIfEfTGmfetDBQMZO0bZAT0MLdvFQnLq
SsFPFB/ZYBYbcUgKx0t6v11cbU1lZ06MymlMPXentBblOuVk7fQNMuh4qb11
bgoOklgpthkshKVnck4uyyRe7eaOpXD7BAAoOdNM2/NZI0m8Ju5A2VzwUSeU
J3/owvwqvMkx4UobqZABTkleZ3QwR3q3aOL4rjlQA+LlBqNUxGnBLjkrw2yD
l1xUBm70Mxav1QhBjKBL+gGKWhxlqV74Vo2+B/FhD7wKLhJFBW/b/NP08QzU
0EqDInV+X22o4vSuilZ824XIffxQ0JP+0a6a7vfFZ/Lj2h4DudzFBs2uB3H8
dWtMgppWLS4zl21mBOMSznRkuAH6V1Ilr+rdGBM4DoTjLeHzcauJNiCMTcBx
VOz9JKNa3NYQ9GbLteMfX0oD2o+O2AzRajSHo2jo+Haojhfp/NMRboGy7DkE
ls1egLElLrL7L8yTrj5jfLYYJ3hwzJ+bQviyHiyC3j9NgDz/23qiMRxxSBxf
ce+8WLekp6QBGhUnghy+cVmc+WdpszHCSDdv/yZk9HczEB8SevkhC4fyzw9q
Nwm3qGw+bdANDNalpYn6SUo4eA7d7cSJzjFN8RQU+Zd1PLo44uUUGPpvBGep
+pstjXq78baijgZKPnxIsT8PzhjVmlqAx9oSajAM4tRIxHWclgnXc90lIQOi
r/qRd2s4imbXDrmGGOkyamAKW1SFdU/mp861uf/0LlgXsgsvLQRmixie+AHE
0QUiTziD0rDBUkXv6AYkGkdZHurkOkDSLQkZVYFMF0sfEav1enrEI0X4x/Vv
jGbR8zWrJMTV1N5Id7BHTuSOsgXZM47rjsfADxSzRcNIRXe9prVkGAbi9lZA
G+gLD0+Timyy2jTI96bvzqTblO6vqKu7AeVRRo5BQv/De6TSGHn4Vw8d1Loi
LOe1x4fHtox/4IUD0uF84tMiG56da4BuXSaUj6mU+1k4qkvMRE5+KMX1MaEL
rD5hODi6dYv9wMLChZ5Cz0vJi3LdvO8OsMleQ4T5/68sMFxHe8hPrGlQ7dYT
r8Ra3BzlOZCOOv9almD8rPEd1qSmOx8WpX3hiZ1bAIyKgPHc+4JSKtbgKbux
qPSwVIrWyc5KtH5HRw0wsGf1csJo0OeD1BIq1tur1r6fYrnKWejPLTrpfv0D
KG3ijx9DbLI3tWXXb8ROUUpBbiXg+t/1vCnL2LEvao18FjOmk5Ru1Vhj06Yr
FyIToWCQZpT28eDt4YC2yB0b3xVtB8mo/QEIVQM9r74BXBQA2vrTfZM+YYkg
PVqTCZSdc3S9Hc73xw1Umlj1t1qCX5PqKWiYBLwEZ7MyL/v2ecLkLlYs/cXC
3u/bhEYrZtNtqJ4D/qdNNRZ95tWx/4IXU8nRjQzEsRHO0ILjWxtJtKoI2U/8
vh/3x2bwfIiSa/M1qcQ0EbzM2QZ9mfvijCAlMce/w9Bj/FgKoOrzv9R9Qu8E
jbRf5L+hJZ5XsZTkkQ8y05VQL1IS9TBJwjKYB9gNBaKMvNQtCdfJoEqfcq4G
pIE8Yelz89E2Ffge7asrjEMVkx7/Yo8y+X2IIxAxUMgMmDS3YMtvGqErGIVJ
TRNGRYojX06x1Kd+ytZWG/rOiH6fvfEDBlgE3p/qrkGkfhx4MRRmKdV8Bz9S
Dlf8EAfa6FzegKzxbHt8o3g+uatKL8lYVROlCTLgPv+WHpteHf4pqjbfDbC8
jRT53x2lMYvpyTllPvTSQXfkzz1GlP9YZ2CDwrE+xugOwhUzJhN095VhrDVO
iy7RYHLOatjL+5HpvGYT3BfwknkuzNWhJ0eOd69BA/upJVskJNPnvqGDugV3
sraX61/mD6NdDN6s9FFSM+9FW+q2aibFMsi4HbQujmalSUYhD6eOyFG98B4m
ZcO7bwfHjo8RIG94vVYJhHjmyBm5O+btUiVvA2yfIlspt5EJvNqLJiEgmonp
ZNpFMBbJcIp485bP+Eo80YyQbDh+nwJweTDQXpC0hSfl1v0f1eVNTw22Li7+
/3gpTdTGxJZCY5Rxy31SROQjSrXyevEt8NFb5034nqDZNBMBynE+KwLjTY4U
SfZTDa5vxYybhZtX8kI2dLiehxKAKW/YEXS+56dl/iAAgPpaXvvKZw9hSYlE
gzXD3OJgcI4YaKF9QEkRVBLi+mkWF66IlUJ3CadsMtSpOT7m4yJ6yw1rwzyE
OZepZCknpS2EtsH3ThmJU8EGTr07x6VvIYMfy+gaLw+iNngwFMNPmPqs4kwa
AN/pFwJuMF0RaNhUMynjk+/88cEWQG+5g4PPw+qeEnDLvHV3726f5q113Scw
PDNd5ZANL5IusoONjFpGvq7ymYUI62jd1bjckbrA/DSwmHL92Z3jL90+O4U5
07+EKRqzl2m8MrvbP5yyXAZasQl3A2J5uBysiFTo8RHPKFhw0p+hVEJ8DY+E
KxcSChG9SUc5pPkhzp9nh2SbzYSHHLj1g7n19UU4Va/WdC6e+2e2Qeo1dIl/
JIjslkprkQKHMnmZ9+3umsW4gin6uu+i0r/FSR46cl8Ns8o80k/KdxAUXV/Y
IX1kpU2YM+OMbp+yiBWLejMAWR79MdpE2jKc5yKHkuum3yLoT3TRGr5KTDtT
IU0VBk3lY75vUwL2Q6VEo7ZEyCNa9HclNXgcnelQo/BAUuvqdl0xu0ZhJemL
ni6txEpaVlvw3eDh0ub46mqLVvh0jDpzn65zEYE2Fy/2x1D3zcIubKm1jg77
S3mbZg9XQanvOtDtWVSO+WMI3wWfj4l0PSFHU+RDwMRMybo5qtFT//S9em9q
5gabyoAUttCYAMxrgkEe6qthlWdSr9ly/v6J1pahkaMeDEzsdt/cv0RPzyOb
ON7ZXzgf8FzQZMBe03JlmAZUJl0KkhTu/SHybafMdMIvq5gDlRQXGtZAPhfi
HvrM+NZwOMwFvYcrUcWUxoqEjoelySxwmvD0jI3g27tKi15U5eepcTGDoLRi
paUjsKjq/96ZIJkLRLhggcIWkUuWDizlw6Hu50w8nAHgZwmf4FEIcTP6f9kj
2BMC/DLR4liJ2AnqjSGNHEK59C6wFgSnNbx3aML1Fy4Ht3tN3fYpyiePGUUa
gXxUmcDDLYTSu6waeNX2nHvdkJe8K/20SrruhIX2d6g8L05ISrsNM4Sw1nnI
N2tV1cGeOW/OyO2q93gzXMrlYRecg1b1pqB6fYZRcgH/OjcZ2Ti+Efoy9T1f
K0Gu5V7nvjT9zniRBcS4DntWeRf7Z7mzLzOOvTSYXmMKyZ+AgyvmVAk34iva
K0ljL8TyGYlCywhR8fPDBbFdSQDCCuogmL/g7vfhxi/zG9i0TZradGm1ErkP
UHgUZCozOblB5J3VTNP9eU0hixBVUxjc1IK/dPMeZ8d/oLj4tMV/w0LIY4w6
kIFkc6yM4JlqJso9k/jFJGdZvDWi2hlbyi2O+7qYA33I8kupXDywhDCmtVUi
b8AztBasDkKj9eJovrVtRnZPi9eoSSpW6+qU63hdlCSOLa/NqE5epvIyh/II
5LCWIDlkrVvyz68Yj/m5d3SMxlDb/c3Y2fnsbZGVsi3aIufSWfF9LOfKwUoo
Ulf74j3b/j3u6gPa9RtJdsrfOR+hw29RDcqcZ2e/k76uSB7QY8EEC5Acd6no
SP3pl6p7Vnr+OWfFulLrhBao9iiqNZfwVLFRUkrQ/9tU0TvKCoKZ6TL7/E12
owzffJbaXTBzzKASzdCyH+yvTKXrSMXhGr6I+rI+f3YkTxBj28gXYJm6s42Y
tMcdQLk698SScNsVb250821szc2z6SRXM8/gcFW50VDfVpLf3hUD2MohQy60
rJT3Gt4ZMoZPJVweTYBz/5qD7B1zkFtwJm3Jl8bc1JlqrC8tksRRk+wCCVxP
7UwZ834TKlhUipGJw2hF3QU6wMr6hfQhriv6dxQd+8V5TSqYnUk92f1265AG
ybFvRS8uVC4G+jIF4IR10iRT+CSNDeluXfjU9TAU9Amtdbj07CsL2jmI7m/S
wKM7prDfO4dsvNScV3LoFk8Dq0dGQ2lwuyz0Jju4znU7atDjO89zdJzpcom5
u4nVABL7Ou266QV4NKq6Fn+l60GkmDGGXqyXHWSa7X9Ijjv5SkGYY32WSaj7
CETDk0fM9niF2ccuP4bbcYbYzIkOcmBfIhea7EtYUAD0upG+t8dgCSUmndwX
+DxAA6doYxzHwnAOugCa1gRsno2l7siQCSc+14SkxbQA0O49AzpL9lmiOk6Q
LwmMJh1CCFfpMlgn7xaf8GVCj5qSghjwzaVBWqGZ/5HoMC4YtAJfb01qg6Yd
RdTQmbYPulue8KsNrBmIpWNXLRB2d2TNwXKTXEAwbIDVs2+clYpLblHEt31+
CUfO728p570dPZIZBFwQxFuKgA8ODnYfEwjU8v010M+pmiPR7My79H+oeDBV
dcNrpzTOt+AMHzz2rS6M27qY+ULe2i27hh8i/Ar9piLprSqaRazlc+yJGDPg
ofhyvrPfF9CDDYkT8YaHo4JyPzQyTna30iQbx/cSKoDtV7mLEiAFLrRluGmB
CseenCfQfraozBKBmgvBYqVX+TFRTpjPMGOiZOXO8wHrIrpTyqa7G057/0Jv
eXmC/iA9H127nR+J/oCbrLs1IeBI84w7I1YCGlrGyaUoupdJ5p+VHh0y3wA9
gKURgA16RiJqfAcMFJalYYMWtmTPS9pJxFfE2hLXPkfr7ws9oSSIzvsq8Plj
HQ65X08LgBMfZYFqCLjrBJsXEHthM76NBmsljTY3r1XxQaf4AsxiHCGNJLwP
tCBsx5AB99oqBrPbrmkdkwZZP8f+8znaHae11SSBOgmYl5HDAzbAaqt7e333
m0D187DmhIOgXBwMnrx12QsPo0hWZhqb9em51UMKXPqf/b9BxEzDY/yxAAXh
jX0rR/5xDoftZgMH48xo68kKE5xgyWVnXRZfi+TxAYTWnby4pUGQqVPQFhhl
3gFgEsGojxcYbBg1V57I/B2w8uVDPBZRj8hIKZ/H3UPf5F1EmXhprc8oKsSh
JbrYwjW12vLCEH+hjglKVtpYtbAWcghQptjFWxxJACJ1R73tRXRqEb4Pr7sb
0ubwqk+2lZZtIWxBBEswTtaEVNHG93rp3DISWlQTi9gsX0aq+ZQ/iX6JUdrI
XrHo3im86+cBQ+OOomSjrmuyP6ou7JQgdNKTK/KYd7UPZp4YG9JzpVI9R9Mt
rWl9XaRe79V2AhQ1gE8GTOFR9ZQ4Pqpmn9VA7wv2z72U7n40KU8vj1zO65cS
KLWr/exaiLVmAC6vWUpgjn/TGMPmQT17z6yjA0YxFxyw8tF82UqaMTMWGctc
agi0h3f3pikM2lEZE/ft8qOFxv/1vShl0oCc+QHbcb7ApD+cUpq9zZC98F1X
DoiHVbgPAXhx4RNQIgZZR8Uj0WW8Tdk9efmIytR9MKlmP6y/btUX0La6jeCO
3Qk3kxVlrZfX749yXCrorw5u1j5pTiGsJsTZFGL4Lihbyiv7iBWSqIIFLHx6
KN9QbsZR26qKQLadyr0vsXWFvR/JIceKfjf0GdebOUseDxkvEN4gUd1ZdmV+
4Aodg1QPvr+sg8TP3hBQ5CGxYGbFJKUdMRaEvx06hH9GD21t6RfqhfFvWSBo
FF2j+AasEKQjQzfp7myvO87ZuYaSaAhTkprzHpEvUPCU1ukMV1eLswnqF/6Z
yYpWufoVsPF2TF57kGYwN9l9mdqpN2A6Qk22FV08f7cQPbCoSOAbrYdA+r7F
na82Nzxp6DhYjBJ5bjaWv1OhcAwpn7V+VK/PPm/wxnCfyBIdOhIbKkpLl+AX
xmWj0a654rIlW99wgK9jkZcQV/AQzqAfmm3d9ZlXVnsz5PKaAZsZGyX57IuL
5S4gdAIFLRW+6VKhqvr7/jw+UiheikJgAZdnSSn1MqE6Z6Qf0NNjObttbO5a
NAcMtFZvjFwWxyrtDaw883IZy0gzrVGQLuWVZQ02vwDjkTRdXrIHCivtAI/W
XJC+HxVc5fqJmzcvAvFExcefM9AKnePoaeNxyxOQTcAtS6zrLCMOiwG/mm+4
XebT8Tk/Y5MzyIIkHuwAh3M3XP3kcBDkoLpiclf8IKSyVN1UnT+xb+uKbeSi
YaO6MepKWRJPlcIi7Qhz8aCQe025GrLRi+B36sP4mtsjUL7WPX7HpHfTJyLF
XyqDHjQPxyQPIjAyNQQSQ2JN0wfy5H0yNj1lcxLKBvNi4CFKJubvWySifL/Z
YjEANPPQSsSqLn4EHRYlpt+FBJ04m1VMt15F7SuGa9Lale3FXzxxnYUlrAke
3U3Lpav9f1y+Yo46a9+D1I9wibC5qtRRucBmtnco0mjMCIoqgzFAYQyaOIgL
NryEFcL24c6vLvPfyhV+b8hu0MCtVUcNkenyryPhLv/Dm1PibJZ9QWZbHMP+
o743MQkPDLXphfS/kJI1w9Wh7W55xxi3YhLPrJDElEV17rHNUKsJPaLi6/E5
MmuSCCSdqEn5j424yLetUMT1qcNIqkJdeCKCos+pzX1J8L/oDbFeXKDnfnxF
HGSgiND5Wej/P7ROD8gMpPijSkTcHQFdh/VpwMd+73kX7Un5NOZIsLOvSawF
CcSJI/oW6PxK+E4N3Kt97NJPxgSvC/6CkAwjb62ashhGd6fzW45JPYyk+rHD
y3h/VR5f7dt6jy9vmGjMUEiBGidGQPUWlrTPYpeBd/dnffUaTeaBxwKNetFw
CyZd8Psq6HxP8tEoykFPBr8hQXjM563ETlpW5B5/JRBwOUM8DCWbwSlbtBOX
slNqOSMVuYgKz/HaBRXFT62YsIp9/whbT914oGP0SNXTyvOvweXX2kGBiM6L
o9esZO3F3Inoxg0r0AoNrRUzab87HplClBzxxj9vRMYHUS7JipBmqUb9XOsC
bD0/rgNNyEu6MaXdpjjfMVXFZVwF7DnmRcjd9KxKTiR1PLtc24kyhByxAhi5
dYcbyAyBOlZ7zHiNhmASVf5iTNIM38DTYkbYZHWN5utwV5q4wP/rNauQSIsU
QPYaBt6IDeqHytE/9hRdxoBoJ+mbQEJhl+89naPwVw2ISMCNXJloyNuZWmt/
fC9hQdRu4MRrpWO/SYF2dmUCefCWMfaSfV6YXraDgnaG2f7y9zGSs0XsZrPr
2A2iWHBSDqHO/aTtSZXaiPYl3LLaq8VrSZYT6YNhyj/X42WuJnzzVWZc0i9q
dMPcLZdsE5MfqzchfeHfV2ef4VxxIkpp3iAj3lLXD3rr/yvxt0SSRCWmr4LH
p1DVp5ANrZE8sp6IgHcQxvm/ehLXO1AVT00TzBSU8HYYkoLy9DGqQSeiGwuf
idMHKGblaWoDyuUMcO0JU3r7jAqZ3rcc2mbthOqqAQICJ7CQA62B6hRSPFc7
ILyba98k2LoP16DjKwfeylrdxogdSmyWyevGDfX3RDIBjlYf2yw4IMt+fb1v
4x7AHdZ2j6bAS+TAI4Jkfkx8fjdv4bK1C1fB0fl1A9fHE77lVaSpMhiI7/+T
mPQ6skfG3m9GDBH2Ewhqds/UjHPQw/Kizc0eRo7fXpjSPH4b6LABMgrv4Qli
BE1E/cMO2ym91tCMHXzbWwnFTZEo6cNgurOzjvbWI95DBJn4V156dGmNlwZ4
vpIVtf47kFhziqVSuEvsIYWAqqsOdPdT25po7YuYo9QnyCkhi0tMACyu9ZlM
ztpDSF0fq0vnMQy/1GU5uXsStomAn+Jq+fzQm2gajjVBbLndswvkTFvhtKwR
FLecZwJUW+Ay9N9rNG1eT0le9i1NJdqsaxz0yeSXGdSxTHDOW7cIIIM0Kj+L
JCfk7gun/ocz2Eai3QiqwOkJWPaL8B6WOFemlqRl07MOYL8tYjIHJ9Ws8Ckv
SmmBfUsXmxYiKrCLyw5kGEUD43AJX+ssHNKY5PzJeiyuH0i3q0GFxVgCo1QH
APK3sSWmtN7MjY5YqpcaB/Ez6BujVczarwfy/KrJn5pGfirIw2nunv3Jr4nf
X/ctteXCqLVIT8t7L7repRGCvOZOd1gRgQwCrH3TdN2+6+wMVdPhqswjJ1xe
cLfx+Azg96SojuoT6oemFKiw6oXMAVGG7fzfN2E66JssfzhUTFukyCoAazGq
8DI68glYX43z+Cd/BfPs7hRLTo39zoSzlkBUqm2z8ATuSbBXoXQm6f5URrnM
jWmk77Q34Hj1uapXevHkqW5vZgIjH8j3a4rrL8DMp3YSGxmXwzr3F/f5sbbl
jUUD8NnIbuJ/1JrZEgI/8hJn+H8v7Ht2sZAkiMjNRNEVpRlHHf2ppHCaodag
CpaSyObNWHYUfOpXyJoBmAd2XPmYsPNbXuyybBhP/AdDmHfyWRas61oGHrWI
iD1UAsC+j7ma1y4zzqKLhyYurUw4SPGPyl9uTn0Gz4dibrSgqH4RREORxlHL
0dyWBPl9UefUTQbXGN4I4eqjTBl2z92CUK86pYCEsRxuIQODAB2dAhEbxf5/
dWejJIwSTpv8ONkHNLIbPoYtywCUM01vDFTcxbt84OfwNgx/D0X2twpxCAG8
40prxwANIjDjEMiFqTLNEEF0PuX8eHci36fyrSoauzOsloEwWA6OPyFFHQ7i
J1NcF9U16T1hgBFQFdaCTRQR7U7UebsYMQCLFLewgZIVZ0hPJv3szwSxMBKi
z1d59VGc88ahIBX/l23zT7DXVnbXDGD8foSjlf0O828yvkGXlVduWk1W1qVJ
5ylnj41j+cH1OGPQyG2kUuCliXVaHTlccV9cPh5G2eY7pImm31BkdcFmPUZx
NFeae/Db03xjStYN6RIWsUOo+/FZKUnHHKiyJ+Zqz2kaGPbbMFZ0ctVG4xaK
xo8TooMryKiQwedinbikXG1CrL+g8TyO4lTv4j+m0XmPPtrukmrYiwv5ivBm
lN5FvpvukM0UEM6rfHQZpUR7TiZGA5cGMFRA6JC7GXIKlpzuZKRqwdEPB3Pr
GVCs9PiLjlXw9S4RI5tZhmM6pn6UoZZzTWcW2KiRSpaXIE3cyBc6KYE6uFYd
6KkxqVP6NW/BVtZVXIeQUHGtL7jEViRAj1rir4xXsjrgBspXePyQMKAqZmy6
nO0HkOJ55eG1aSNYYZ2yf1eLyRDGDxQyH09MLa7P9OnpGpq1mRrTIJ+hzlQY
zcQriO3JB0lhxqjq2veEY/1/8cvu6bmTvbKJ2eYhyL5KEkNEloI7VvtNoiNI
BVILWnGXn5W6pVkKgmlnEyUXsA8hHX9fo9U61hbHkI8yzmS+FvQH6f7LW+ZJ
uKhLpFthhEqpB0aqtaTpRn47O74g7vo9Rehmqm9qLqinl/QbP/PxuWeO1Qqo
Oujv23uN4GTQmmBuATYk+GB/d6+SQpNnCFcKRPDNaSFmcKHmAklpTOGcUmPz
+i4gaTasFtpESz/ryoqRWcJmdqFjxJXaEs3NtNavphhtLexKUVBTdqmFQmrb
E2VU6nPxm7CcGzajnI9bK90KqIZAW4nSeZgWUY7+9BD8xgFfIUC1Yasb6Vir
jbOYYEBpCKNgMqUh8164aIdTJCl6hfUHhgDxSpyJRg/xvIgGCbbPZ+uNKOvD
NbqNqxUbHfvZEkG5VeMgYswe2ZmZMzFBm4KgLKmJ/fn+dJosFYI/Nw2YJKEi
3eEi0vfYWrXa6I2FdsfGlmGfVtf78sJiDA6w7Q81on4w0y/uJj8rYT1RYztE
wZ8GXP52NG8KT8Kle3UjSJAR5XuQ1myNdCQkIH4hC0GFUmZE9ri73LQtVrar
pJ7YMLXvO4GwTcn7R00jRCJXcNQrmi11iIUuOJ/BejFPoS3rn2j4j8rT8HoM
ACvyVICen9+kggf+DombPiAIWDjQ4lOE2uk3+3eTkS/kRZAml/KbD4+ZNp9O
kjGo/UJz2LRFG9dTDS2vRumpF6tKNDkamqV6CwIUJSZq+r8ebgvou0ZPWLSQ
ag81mjZlKVrrj3wWZrFmdzd5tW14XzTUhfiIOf70jTaEu3YcF8Mh7gb0xBmp
tAN/G3qvjwKXPOZMmahpvdfmLLfB7L6DcMmJz8mKNzHxq67cgaB8RxsIcQ46
LkjUOBLa15QUX1lyTPkKdf7+WwQUMDAFW22jHfmYRSTc3g5AsfSQu6oAye3U
LOgNuC2CGs7jG1wGFCUgMxopvSx45kdbkMROGBTfMTulf8DWF2097utCM4yC
AN+ico96vb+DUwY79pZXnLOmhrRkSONkC3LHFOxW5AAUjFi9rL7qCcP9mC0R
M2xP74vrpKtc7ghSDT3Hb48V2Er1fwyiIdatFbxQ4m33BpmYQXAotxZKdvYc
QlKXDrPCYgFep4GNknEKpM2/khDkgL91FEP4gjzru3q+HLkPTZrMR4ul8hQm
vrn+hWhM5iixjlv9UffELeDY+5lhLsj5SJgst2Vac/fNLQ3liDzs/t1bqB+0
c6iRh6L4EqRgZa+hjBpfJq/jPr6v1hAQaV4wGzEZTZlQrM1eoQ0yWnZ+BD99
NzJz7efbivXP1DPuNsF2RpONDp+Xt+9/FXNKHvbhdM+LP4rjOcO6WVOfySYO
wVKHig+ZtlCC4zCjGQ+cdrGD+tGo0lJv0thLwKkLVg3QODnkQzdwOr++FRSg
hxhArGW4QFLvMbwaXQKUb7fcAEt3PjXTHDH7dpN1sFzTbM0njOspCmffMGuT
ylwbspsCGHHQ4TzcYfVm08mrFkIdoZ0xcW0uLBuD+cO4za7KHXzXL3rh5Pgz
uOYYejepunBFme+ev9rLnsUktpnbJkNxf0yE8LuoVZHd8+yfFeHk22zYkI2g
j6i5QPSdjc5I+zkdQ8fsQd7cXc7ObXtQbhiHOE1ppjBmL2dLSPaihwvMj2B3
9it8d4LSSCOiB2aBdNgGPhloLFSB6EqKnhjdx3BuHS8gJPSOs3MuRgTbfG5z
S8E8147siw94ykUAzeXQhYDhV4ztRQlRF51lJZgmasaRzyorJmjWXO4gn4p4
UY8FT6jZiaWeM3Fej51qYNvmhQGkN4wFGXuatNygyE+oSf1U2XjmROvkLYBQ
XeV3C7+8W1RPM9R2XveRytS+9TiissuGvDCy0UjIW4Wp2uzFLAftko7mvlXe
KraTl873p0JpwZZjuVmtwpsPGdwl4zbvANKujCj7U4VtoLFvVW/IaEnWB+1X
VruG4MXZE5ZBvt9lAv5fdywDx1Qs3OWl8djB7TdvSddIo2aNFFIMct9jmmwi
Mng/QYxxfuu+678bo3W2uAD/icDVJOKQdLxhg9m6d45q8XuLR7unpBZYtATU
ixzDR+wNWs0FnhFdI9OKHJYrcAk+csaPv6GN5fOFvJqVqQfuwbWJE+4tISXb
CgjXatGVO2odI8dzffRr43ftp3CHE117BpHKWxv5teI6l98Qi6YVISC70QPY
4CreHZnfaN0mOKvNfmEhvL+dUI/B+mAcUafRVOSLO2Eu12pqs+uS3OGebpvw
m6IPKA1OU5++cMp6KA0k1HQXh2LLAd7l03BGFzGvNeRxVEhPTrfZd6vwvsAJ
Y/RyXskJaUj85yrbmSIG0ycffBYzGw5PaJ1qDQWyfx6/kE1VrNpIHC3PPGMM
e+oeI0JBujJ30vQaGCLIJ2NWUNc5Y9knUAfAP/hFE+sIBkncHuiJzRusb9X0
jKLc6w3zOS0BDOzRwmH47zdQpRDAGixkewZpEwa+EoKoJQ2VIsOBAMqf+zu6
XLPpr3dMIrJH1qli/9BWY/UhD3BGgaLmP9XUER7NLNFO7xWJvsPoew3irHFJ
0MJtPg+/krFriiRFJvJ+QGDjzLbm557bJQ/mlXwJoBissmZHmT7yFRtXH/zk
X1rOe8wWdgDmKaxXYFdHTzJgpkdYbw3WUxLy0Qhbx31oNgCMm3DxPxoOilQH
BJjN9UK2Jmhyq5x+9rIloZTWS+3rlsuotYSdreRJUDmKHo/eEQJHdzxkR2B1
e8PGungEZkureg4U9JIA6ZHzBDP8GiItQRwLab+fxsAuVjkhoL0qa9YyvxEA
ryoT21/FjAl5U3A+djiu6yljxafv9cYbrDm6s9BOJtBiY39b2SbOcTq5WPa1
53rb9yvdHKgnCQxnvzszZcQQSc3NSNEzvhsofAl22jZDEtCJ5kOcEKFzZz6o
2faR+pm4Yxe6iNCrgPp66Pj/7WU7KmnS1Y4vbU889sJd8w6I4eeOWCui6SvF
0GaXRhuKHOyK181zxTmxFuEuoeivwE3X3bYSTlX2fTi9Qru2xS/L9go0fSkg
xV8rdErf7rVIlLUlIU7+3uKOHFIkfDdheivUCG0u46sTLDb/XGl/LtYaTjQy
So+/r32Y29bvOlHJXJJMuqrP4RKY9rPHt5dszdReKhItE+Oss54ZjdsLh2aq
8muweztVtMiHR+d0nf0i6/AzPHJFWCb/AAxNwfiJVagD0nbf5YLj3RuHZAvB
xUALTwY1vKBlGFbV3V1/Jj8Ak+R3hFZoE1G9ZrJemtoD3Q3pDvWeIXIwVWE+
yNNLJlQETNp7MaT7mp2wHOdo47HEoDigSpOZzf5JiJTMYThxc7HelYm3Evs9
tGMAgAdknUqW/Ds8rKRR0vVdymM73KvvItJl26Dg49o0vP63dKz1O57+jnLY
dIxzzYDF546lBFEqYqchoyLWk/RN1PyqwMreOxmZxm7nShzQqWkNCebFriKY
KbKyd7fyHU0vwF/OU5bG/BCw+JGx5Mwg5EKzHm9JC/AcZFpl2npv3rUDeMAU
w+keqhfcQ+ADHhf/+/ff1j2km/7D8z1UJosw1sfyshKnXLU2+FBdtjiG7NBf
+Tzt3SKTn9zyMvxB+RjUxJKD+0feJglC9OdHbgGzzYsZvUDJ71/a8B/sHulO
jKXaPIKlxfydEg/Da1fxoq6qE5M4BQDkI5Kgk63ZMOUuwCErU5WpJtaZg4ZN
vzMrpr1Y5SdqdpRWPvpRCmik9vspDPzO4dH4laZKb30ryuFxRAIlaKg6OplD
mEOYExyaWSCZOW52qjirmHzC7OYmJ8HC1dB6BSieRv1adnXwYLwc6PMwsBio
5EjUROfQT2q+MsASue/U6iYoyefTHVgaWGRXdGvFl6/b2OTzuM+3jiauWPuq
6eY6ILhtl22mb28CgP9sav7he8BZKzOZpA2uEC8HEyj7mH2NqzoMbmubOjg+
dPsPUosG62GwWCa2TKpaBxUAmdJdz3W1ZWIGID4CjWBptLqjwVVa+BrbQxNv
2UKu/Fsntvp1r9Fxp9KP+i39SnO+7NMxtEkJq1najYiMQ3iGjmLOh1vqektW
mgq2gqgfuGCUWYdDCsrT4lBVaE+K/x7Q2y/r2zsMxSmIE33RE/vZ2E+6ecsO
fhq9//poMivKqrVyuQftW75lUdDdedSFMbMaSxHQ4t++M0QadRxjxlnFxNnw
1fsxroVMyc5JS4TOS7ISsRsdt7T/0e1uMDCJRFqS7oH/QIklxvED+CHeuqa2
feX3zkskv1DmEN3WlWgldB1cAyyI0eysC2PYou7X1Mt1GpnjdDojvgG/5w+3
XYq7o51qMCgEk0jqL8GxxacaEJXAReK/l+Izax7eBqLX6s18BWJmovYHy2YF
GdVuGSucFTtmbPQvemRf7T/fN4g4t55AtTjKszYnupej0Fepg2KXvfpGFedT
mLJqQbiyXmWY15EHuCe4pV/RPSxwzyrma6ei/4HbDvuPGk3DtI4ejR/Shhs9
Tg2kVpNFJts4Db4z+LfLrlxAJIRLIvNNZ2vdXDCATNAOHdMxmemV8mss6kyr
1d2C7yr9420xANS/K6mTafGCuNOEtjWyiNMvKoR1KIgBJYszpoN7Qo7thAyX
+wC0M0keG9or2C9xsu1xpo/wQntKOEzw7nD8+Ul2pzSFYJIW8oW++A7FqREn
26ltvZVi5ebXsvzsWaXbl+bzrfAYZ98OZl1ZBQiqCKhwF26zSO+cLWoViF4y
DCB4XN/SstNowndEY3yvV1lTtASb+5WR8Emd9wEsNygNHPW2eYIUd3vm2NSI
oB5T9ler44C1RwJ2D0DJDXhHdYktjGavFJvCuFT/HQm8tsg7EiDKLrOEh5Xd
+O+LHYF7zhCVMDIccf3Ww1NJ/g0W9pTdiwAeS60iEKSXgW0JfslX71t3nWar
YuWAlWVUTXaei4mH4qNKxiMIMQ8hOfBNkXlYWOqgM9QqI+X8XpoPy6PFjFNZ
m1edyKONL5gQB+ngrGeUtAd1sYHrEWG57LsDQTIsqk6I5pd8+QKA1ZT2iyIH
s5F/9trfgmvVdGF1Z4WF7Xxw5Uw593fu1rAZKZ8jj/ui2YCK+jdbBzouE/F9
p8h0OMZLzWloUI9QBCynfnaRUPvkTglEc9ZfiMcPz6Dw509n3FIzOVVdiyi5
sVfxotT3txECWqjNIIdUBuOQh4/tKM40onNXqxnbBX70sQqLChKCUMLbTwIg
XnV2L/fX5d7BKSfQc3+3hh20Fqm2GswWA8YYR40eMBj9/n8geZ+ZB7EnetYF
dbMRWzwAtFlBjBnM/Nm4RIuytZTW7MQ2ylVxbT3UBbJlyKWTEVWR/RWrF/qz
O1hzmp2s6uQNYYjTYfn3gRuHG4U6sIB1X0pT9PBoXZoLejW+rVbb8IiiJJy4
FGDIj+NjhFt5t2m3PiFCFvfhRUowrt39eWRUlfq5MRuvpFtAIvkc/edWMFvg
H6UxtqxjOmY45/olEMMlT2ULFNB4BCfm5mdzHRMaFJ0I3oEne7YgihSUT29g
R18GRYJNxHB+dR5vWib13iVFDanEfncgDBiauJtJFtm2wq4E1z8X6RJMQA92
rI4h/aB8lLsWgCUrERvLS/C5v1cw6WcljubewaOltcdCKpDA8tdlIGtzdO5H
BY9QWwH85dmJZnx7JRAxQ11rjriT26qUcVdDAW2pactybBx71Mgt5rcFXY/M
SVfnm0/7gcNvf0CfyMTxIqKU6U4LMD0eglMCwcX9/uKFSNc6chWKRejlo+Hu
uQRtUvY9TKqDR5AOAj9mMjkymtJt9RBjCpF5ZVP3YPMexyL9Y9iBGGbCaMR8
EhkFhXvkkTAzLSJWS1Zg5yhoumMi+5ulYWoJsqnsDGRxcaDVggFCygWIUpCO
MBWLBawttQhmuWt9ZaQc3FH3Rh0QwFgD/FCfkJgPd/Lqls+3mSkS7v2EmmBN
5zhlC0DjOLWOhTFPs4KV+JEZXRIaTfsTw6zbVFxn2iPplh9yvJa9vvg8AOhi
rqnhzpdsxtUA4VwEfS12ORxe/Ty31affH60DXooU2F1UbCfWIk6IdqrAU5GP
1Xmm0XNmNv/Lio6r0xmQGwOQbO49kD5uKa4LCpBb98jmVve8iquwTuEv6Iqc
w0pJw3mKl5CSvmIaH/B/Ol/ZrsE6XCRkRdIirnH7Fi1y1cps+kYhxbSp7oJV
Ils4NNUwdpT3EwktvXCW6w3Dps/+xvTRzLaviqlXG5i5AHN71d8I6crwe0yi
8GnSoLlMEUSjco5uDOsexE9s+9K7eFjfw/iCjLd0gMqkf5hro5HLl5Gf/k8P
0nsZJBp0HtxctfkCcCE9v7Q9Ie5wVgJw6NkgLBDWQYkLOpiG9MWU6wZGsF8Q
VO8AKBmSSmcHLman6DgJMU0e7F5zN77ntjes+jETP64AjSKny5s4I1+KGQhB
CkW8WUjKphJ2wokub8VYqX+2ceOkniugaAEX07Ifa1q1lLvqytaHwkM9/LnZ
DauqN6weQgnovLg5T5PeeXkQ3a9Vioqx0M1cCGcvxqWl0ar2gjM0/zxk8s+M
lDCMcGEQOEYG100UEOlpc+LXRaw090Ee6hmkCYxvW3oz/Xghm0vB55GRqJpc
PDg+fU7SBbnnUk+9CvGTCrGGwfGpNdelK+YiTkTLZ6/RMQqcB0vV0wtGrLeN
FED6mh2wzq+N007mWN42RK6aN0hKt/t8aqFWsxQ3/DW4l09RpZe9jgHqcmVN
P+nma4QtVaaRRhMXiqEvOPgSjokfLlil5AQNbsQA3IiLhsjKJvIuCKDO7RGh
Q5Gm3ahk751fEzdyFjr5uhgnOqMa5RfNQW4y0XOdkPkjeW2vYaQ3QIhqeVni
Kjqyp6iMbzLPjKk166CkTohdzKWiDArCj5/s/Yh0icza5K2+capdQzT0dzRM
Z7tSqaRiOel2bpjj4SNDvcXo53d5G79hUluPfDoa4Mgsyzgh2AOdOy5tm9YD
1/houYr255XTjomMbMssVDbzM5rD7pDWqNy2euAiSF6UCFMchlZ2FudJ8n0V
cmydTNt93YrOpjaGO3Alz9/p5GpQ9I5JAJd/Q+YLIVOZmLEtfaU7+jvrMqFP
RRYtDxrB0/BrpecJRLYcDK/0uGjOdn7SM73VRMTNbp2XIVkeq6s97HkEbw0e
INM4/RvzAaCMigNLklTxlxHJDUYBscGcU+65I1q0Q6Dh1s+BUXiMpqlMSz+m
BMOjl889+lzn/KZYj+X0gX44pwQHRrbwW8ubsgxBqjzWOVDmolRIj2oDtmAj
tLdNHAlc8yKkhdhvyLmLYxgJhROBoXeaGvEov0yX/riSY4tYp7IQOHaOARr1
qfkP+cqFOf+GEkI0fHF/R+fWrjzyQqzEIYcGpcmLKXmwn0aV6EPpLBeNt2I6
OlFDCMtqB2HD7TB3A4xftzPjXsDnsRR6s/gAvaQMv1iRtfZ3G3fukHJk410a
3HOYazmixwVSDT4LVE0nrCBuzHqNFN27m6/zmgEuWyqbaylqFo/9v+xc702A
sfjI9T1w6b5Ezy06zeJkUxmQCLywa4BHQEzv/ZuwNCdEwuxtr2w8cMKC7pLG
zWIL/ECIKnGQl+cmvMSGMhGvyo9F84ZnY1iEnDhThBGCdeETm20jDI439MQ7
5cFcxmkVdgb/Hx3dawjYwm4zfIAgL6urdO1fhwabs3PK7hDy/EIhDEClzmg5
7NlWEn4xGnQ6xt+It7MAqp2XFVJ3VeFonwfbBHl8Fmw1OAXvLbU2oGzBYmna
kl6xZYLNH8x2oLIE/JW8HfFJ16ji83NO9P+qD+L39yuJ/Ml6t85ahQ4xQ1Xm
R1xv0xXSWMRwi76XbgAg9AMBBqINvwWYdc+v5IRiTwgi1kf56fJ3irNUntOg
5DsbvQJ7WTJPU2oMdgKweindWtNFwcFunjlGYWGzAokNxt1NfLZQEkKNac7i
uwZdbCktzrQYc7EwK3KwDC85Fzso5pkAxuivJJTa2lUFelQc/Jfk3GTqVdtj
8KH7U+PlbuHCHW+1M6mQmVwyUVHo3N7N/0d2/u2hZoM2PoTBgwCnC+MLWvRI
8gzM8X91ZdlgOdcHxBoalo+IVM4KweDbrzs7PjOZ36ulwyvvhvMA4rexovaE
C32kUfXUAYafcJmld94/vl8jBMhauNdQtzvhTXq7LPiI1wxl1VH2RYHe3x3d
pq3tRDNQGyE7WK70il+3g3I44cK8j2cPF7UFAiokbGkPNTSZ2bCNQ2Rhmb3O
rERKJvkoAF8hn3t2q8BoypAPrybbMwNJMpvM3GjkC05OiL6focD6PeD7VXIG
xb7JSZykP39JELuVh58WJv/6HsYscGkPIYku+yRga1DajNbiteKgH62ytYG2
4d5U6RgPKza22uM3cYR/96R+YHLDlhvmQe1U+JiAyQ+q3nBUVwROodgXqJKv
msQ0Je+jKnebDMjuS6/Aw7CJRJi+ZrTfPpc0bUPZS37ZhlTDdyyYV4Bg16J0
p73IBOwCQs2udnyo9jCIrSeowChzRoIfj+31ZBGgyJPHT5VmDgst/yQZezN/
kBE+7Iq2X7kHnmHfSha1nPBNwixydfA09LVjbGqZWeKYm8z3Q0qjzJZ7Outh
zusLmuQgdWwdCkKblQfKiyj0i7Rb4cU4XtodJdGB8v49pUG31bKohT4vOTZj
7Vo5J2BmCo8n1gq+DYdiQ3m8Nw72oprc47Cx++u9RE3mGygd00Q4x+QQMgpI
3AIQAo0qxh4eGVMZO/YwrMB9qkp2n/r5tgyC1lkG33P79MxnUU4hTWYe+zKK
QZ0tjEjfhtIlHDaJHP3pUKaU1fDSJgyGkfgPhRoSgUdpUdUZEL2o1kStxM/Y
uwl6QvZPLqFeZtY3fEJO4jHclLyo5qTVHvLRysehuHfh9AtVIGNo1GKWyFpK
2wQJxhYoYqOSYfbhdzMmbBpS5zlnJBQTiivpkTdmiErV3QUVXAmXHMjKEtq8
Qjp0skwcIRX+E9V0j2347XePYC+iLlKKGhrzGHznL/ifIlkBORtZrqLyNqSJ
JoymQEA8fOaZ3LDk6wZEcSItT1iH2RSF606LijTDmpSGM95NM/DkFlzh8KZd
x6uwzezmOg5UcBkHqUaZi76wl7UGdwktiDyukVNJWlTDoPvEb2N5AaLgFCp1
r68xAzz0w2L/OCXDH2b7QGuydXfCD7M/eGyL1hPpBwbMnM1OSxaq83t8tRhL
+Q/cwzTIsLJJdCxJLLCw3YoDyZD8WIEl6Hm6vudowwSDVKdQK9zGm31ztGMl
OQ9ZGJYr0KI66SQKtA5dlxoz3Llz/1W0Xe/YCPq8jEcoNm3eK5ImhQ+RLiqs
n/SdPm0mXRjpTJ7WFUpi/d73qByuItHcMrl8LAkvFowNigd1eyGSc4qrU3tt
MXyNiq/dH9xtOWx38nqo11o+Jvqwm6wKd1ORbxl3L8nElH9nMwmXV7yQzQQ9
mIuIrKEOztGoVPj9QSrz7wijA+at2ZSJ5ENhJd8YAKjjVZJ9l9vwqCVMwXPL
VpIrk6KnOy1i+9HZFDgZFDU+HKuBSRLVampyGse+c35QtMa29CAMEuwvWp7s
IlIa1B0xZGJYFVo4gcmtWsLCqLaPP0zGxJR87C3Z9AjiAvJNMyLsqW+riFFi
nfkAn2wNzD6l3cMQ4JjYxF1RFwO6G8j5HdPTC6DtxRgd8nSCJDAVrn3Dardr
deN55SuYb5QwLJbtZIcNWUIl9S7n7hQlz+qVaP77L+8wFAUe1GkFLKyA6f+E
KnzhOLRN30zd5llCQwaOKqBOgvxCj22Car5uvtM8/LE/0EJ4KCdfv53KarIQ
u1VnwtGByMVar9p2/6VQJS4gJOdT8ribnwmOCxFOuBFM5cKKqssLOvvl1m2P
sjyGVJcF720/aqS8dxpmXkKy7SPOUEPpCUMOSiF6XPVtqCU6YOiV+KBBUd6y
nPy7Lmk4tvX8yHH+mxG0XKZxfxjcfl2F7KG//HUNfVArCtd1Q+Vrcqji36HU
8MI3oNbCb4BmJNPGbPxS4EbX8PIZePKmk5zxNcYh2JGBvWr5qztWZXghINSC
fcpNQwIITTsXuDS6iEPRg7ZxIkYu4snP6UAybzuCIyK7+T2cX1nRFNiAO9Af
xEDInk3OXVE/sYwTUWt3arcmxQF4h7salspZWrbPXPfEm5rK9OsvoqRrOflM
BwfnlszOKDPhVSGJGv+koCa8nqux0yY9T1v9mDW2ZUu0m6UOzEzISep4X27d
Pv51meYCdHeCtBgt5d7lBQ2QkJ1yoacz3yNn8MUd4yA7n8rZ2oIENPjeUWCh
0+87pKl8oSYJajJo2OXNotl9hEByjjT9IoXG8XJUVMoOAsBe45obJDQzJMK4
nfgcmy3J0sSOUQgWU5XyXQ3RLtJu4H7GuzFswlpDHdk+1HkRgGUkCImMezk6
fGqDE3D6dtRCWY6rU97uIG9WtFTuYPUSO9OUb/rgbzAB8hzwRbQU6h+BkfeF
fruskISwiGMovOdKbKH6oD9HSwl0hKu0xWhFklZ9WepK+JXW/FG4E+SdW0ee
/JkHKEun9Ff/amoG8SxyJFJyEwjGpNGz1mqSUjIrgB4QMtWCpnA1LKZQiQ/p
SrHMkHhEXuKLrE0np4n7+eaMMr1DagIUIHqKurONLjjQNZVYW7J6WfyMoyYh
58vfHrHS9Jiucr7spG8/fYVb3/ZgoVCWHE1DLuef0nzzaoDnG+TpNUGe1pyj
v1ABjFHiwxVDM7DQw0VXETZkNQjwq4lV6bjFGwBUwZk4v6QB0+6RW3VpFJH3
u5um/ZpTvujCsbxr7wZ1oW1OJCz065RcvDtWYizjRzXUItUHRarIACPRlOsp
SSbWOB4C9lpmE9a3hoEzI8Tct5DLKlJfaCMXCT78QaRC40dqfx8w7vgblPnK
lgelPPTYgdOGQHi1v5/Re1NCHZ2PiCDdNwSWvV6p0SsvV87P7jNgFZD+xgrn
WaJZ3uCnMP/uO1EYku804+0cOU1gUfuaDfL18LcEnXK/ZVQziI48WbXyvDJ+
+uihDDGYO/zx5syuFeGmkS810TMLfrREH9lL1MKKPe/aLRdvYfM8JD0q7nDZ
bh2UdMzs74c/VYLZD8Mxii4jiNLu7kaWVVCgOvaJt4qRpHlizS9ypfy7fCEO
MzuPHfcyLKBLcN2h+XUS3sKFPJZav/RNdzYWvX0JWgo1K5wygXEb3LfhEmRe
SaFmi8lLQM5EjMN9KOyWGMHkMfNjEsLKSiCGJVmVTcKkIVMtgNn2wJM3F1zu
yjruo1vPzD/Cy3i9dqrzwt89RejglMmHI6ZXdCGXJn2qPJs+uqSitNAe/ZqZ
pDQ+/JwhFB5tpaA0CWsHWnnRBXdyA30fK6z2xdb4rAvS4KlKe3nAvpemcDsS
jVjvukOFKnL7bBwR+Mo3qzWU/1LiKZRtIxGdNGNdjaHOGtHNR/uumAeiVB5G
PF7xkKlNKbBjkbDsoqRdKOjc4i7/Q5gALR3i0Cp+tN80HTPuuQnenHsHTWCt
HGyYpWuK9qNybPf1b80L+OU/AXJ8xGK6cPD8uT4KtQnnZGr/P4qPqZ4QphPH
mqX82e9S7ut7z2TtaGdtBmt4dsQJgdT9JyxRuBAY7t0ESq+DrLi6PBvyjijY
2RBcRRxENwbqccLI9vsQP5F7RHu4jUgF4WNAujA72B3iI3ODM7ScvQS/JhPR
J+sb4yi7SctrdS+c5p0NbmeZt+LA/j5BUJ1yoIWkROE9YOnUSGoP9vfaqgjO
xmhG7DPVi/eTplwkgw1ocSLc7pV3dG7qlIjje+jevOYNNx1tIRR4w5DMPT8M
cWK3eSq5T760dQWyxf+MTMuf0Hif7QVEXB6stCRINokEUNtOQ3I16lvs4iZa
z4fu6c7gzB7VGBffl1zy9bcoE99azf0oaJKnb/uQqTiqgCF46eY0ECvAfZ2C
fpwx8Z2fVz5LDbH+vGCPC/7/2KR2xmg53Kn1/CgsQXrGVvjomRU7DiEBMl92
GGLXbXsDP5XH7PRjSw05gYBzdaw3wT3STGlAwz8YZgXoJz8vT+z7OPc4otEj
QfZ7CittefqkasiNgVBiSRoYIpWPpxSlG0pXNBQUi2nPAMTXZ5dVZRAci5SV
CQvrLoXgrqoNPpFkfMKIMOcoCllIbQVKPK3+SzzI44p+k/HMTE42rRtOCZBt
OuVpn1lAG7V3Q0HXm2K29ycb3BRWt1AIelYYTXkTwQ7i570mn54uqcjlMhF+
VAFjmhyGB9nkEkjohcpywEH/GKORGc2BGPGAIP9nUmrVU0yzVE0IcdBXpC3W
fE0QnPUXL9gzsd2620XReEEdMALtSvNZtzmRap3VdlUQr7H6nW0f+Ti4HeKU
zQsVNtyqtYHDRXzNzY6mN514+163/l/YdpbW49q6Uc4nz/92ORMGmdn36CjN
CjWQNBz4QgM+ZRGhILxfHb4pcRqebaWXlFDLEhANG09PVawdDFcm7+48wiBu
wiywpHexc9USK9d9zS47hbrP7W5QTA6oKVS97G/7R3kQsyVdESL9Zm3AG8lP
rNeJm0DXPvqK1LIfi2JNBjGb8WtMntYh9Gz6v4lU57rIfV6mLvrFzX7yMSVj
SRNl/DwS4iqumqQsrfYTc3lMErvKHfSzGIvBOXvOq4tdScqzNE87lIWHp3W8
7HiE9499vEKDthHSeI0qogpM5n7aVc9ouKKK5/TXuBfESutlA/49eRPm67pL
RGtodPvDaTmNyxqrax39gsijkF5ETj9vyPGlQvamNKgeQkDzWgjrt/OHWTXJ
FV+7zDc6z8i0MHob1wWIrzR5HcQdsnkqwSlNQtgIvpe98zViAEeYZFc8B+vF
4leiogTAt+wLJSS8KhpvNjKlV6ur8Jum9ZuylUY88reyqZhvjE7GRgGTCT5h
DCnGgiHXnqjcp9DOHhZK5UA5WGbV9j8CEhs8CrvjDrUGY09ou1romDwF4mzn
mlCNNy1PrWZa+VJvEn+JEz1LQnnvfYZ/dCdBs7oIbvjv7hYuN1EEZbkCKH24
84nsORkZuuCWbSwdu1gsjvfQIdHqJ6OZs+1vp3PGNNTi/SNJDNheeuTNVK4K
ntKWgyUYc1Kg8waoje6xssjgL76rwPep/Ead8oWhYsnJiWJ+45qpcbXMJoWZ
D8SMT1H4gZ/7zbbo7grq1oLxJr+ULLGkl3uZT5gS6p4B1eticAsKpegael8v
7855gpJDsu2pw4tKRoUnqJISvm3aIxDgMXiLiMFXPsKi7NpH26kUZxsSn80C
Mg0+EEwhbzKBPMxVgQRWEZc9w9gioatNxhv87GvF8WXPqG6HVYr/LKMpy2hS
oRiZxClv8i5aew6zpCLSOx3KhkeQwP4MkMnQ3r48JzdNFGs6agu6lkXoyGZ0
jfc61tQhlM3WNncM6EpQuvLdfHNG6mpSMMi1BHS9yySElyFBQSE8TeU+nCAk
OSR8rs3/HW6Jg1O622PT9n49nyTS15youEjBSykhZf2cvBN4GzbvhV2ybbJW
59zKeHDmuijrohxRaco1jNWa6+M1Hlnax8wvqtoFW6iJkbDK/RuboFfqb6TS
3d5Pr4HT1m18m9X9oQgzhCNLXXpABP1+r4YJ2t+fiv5yCci1AfAaqT9c/8BX
NwIFpWINYLAVImNB+2BhPxDoGzSf7tQ/QRZxNsu9dWfSZthbzQCG6IKdM9Cl
Y1DQHh9YxP6cvea5fwEOejTTn0dEot7DPpDtidRUGGmkEroAdDS2sbMCQ71O
FcUeGL8yxytg/yQOPNN0e0o8ayN3eEBe7c3aDVMThR18z9IEOdFYVEvkAp2j
ez1Ka0nbLEQGLC5vKGlsOZO13PBjkbLBgAiy7oInJ65waJ4K9QgfjaddzC53
uVKnQD7WVxM89cDPRBk1HFzzJuhUdEMWcQbliEe5R2F0RrfWsw1ypbWOoKAw
YmLoszIFmb1OocyGgW1nDZKnAMYjdgDOxAGw+SxKhfhbQZYt87s0wNIS6kHC
T79qFFRGhIWjYuUNZ6uLa3oIlAIH1C2VvGpL89kMFbxzjFKKWrmDlmjLMKV0
7KOFPVEyqTa3OG/2jwEiF6QBONzm5B/O6emNi5mhSEdrJ5qRmYbVmf/pKIiz
oWZ804j8kdSEReQ/yLCgJGDMKIrxDFcwugcPwux1KB2zdmDOEWu/hVmAprHF
MEO4XUSTkjO7YPcqE7Ij1kDOtjAgpUVocUHq/DkyeELQ+XWdbtwkmo25W5jY
Xcu5BQwBKrAFl/NVUF9obYRizQ/s7QSKCmEgEim2aMFdYxeMYpQlvvaEhq4Z
syyXlNQIfvXZOA2QtKH/g/Zkk588h4YdTIkG/+0ZHtoQ7Yvb3Mmw0rqsatRj
dDHdXwfeMggt+sQIrsIOuY9snP6dQN+NwsBe6GKpJV3iGa4yy7EPdup46QFG
3AuUu9WgthiEFVWFN5ToKnlxfQtn/KJf1csRYXhX6f7Tv4MkTJyol8JEr5VA
B3Q7/vXX58s4almdO8ZV0FjYPm63dYJO+2/OHdgJz/6UluqmRLWwZHrh17fk
Okai2+nfbr1npfuXD4y81h7DngS3LOGmIIbpQaoswNb3dmeFZRNHokqyW/+r
z4YVXjWymQktOlklbmnvD4UrMcLxx+F1aubmDZJp6Fvh9mjsl9vUBPcloG9E
PvfkC1pppQOSWtn3jW0BE2ZEdJN6DAGvQtTMgsMwx7Smb+ewrPlD7JCOTDxB
5SRURerdLDPRRWGrxaExrv8vl2sED9BbHbBvgJxJsXPPy4GvQF3Vrm2Sq5HT
f6AxS7YBt9omAqrTtPbdxIGmFt8qBZ5Ziim9JOLjizmOF6BiOgUlPwo8ldS1
zu5tmZeUGCgqJe9HTm63UlLAbYGxs+605gu0IEb8xUtPVswnDUhn/Hs0RcPs
SVpPhCne/2zjrIT8vkNgKB5dRlr56UbNtt9k7DNWImkklYbiXeL1ccDXfBNw
oBr9QSMuMdJrk3vmOU4CHABgeIKyuScIFTUfaCModhZdkQwlouM1tBGa6udC
GA3ODZWiuEXlCsbBpRNV9I76JCWZCtYnIGn2g+2K0a2EE/CUQoWyWF54AFc8
E9X9M/Z7lyIQ2MwSKuMJ8AyhqaWvzCqHgdbMUGW3+tVs+FDxjt3laMMyExAp
6zD5+XfD9TUqAQplQTYbMoJfq0gxm6vETgZVpvdOJ5lD+0y51xFw/CFYDSWy
d6itne2H6gqp5kJ1+IpsGTnnRZsE0U/whtJMwunyUbCCttHd2nBm8fhXhlil
3jYanEJ1yfOQzJNWYOB/w7hXh80xwBNvmayEPKdzYcX3WRKp6oxZhnwOpRQ+
TxONLSmmO8LazC5ALSTmW9jT4PRSYaYmVLq8y5bXSYTSWxqH/97TCWPFeD4d
+WGPEflZ5pPuQFAhJInWsMq0sPFB7cxtHSK4Qgk376Ed2/78C2Gi1id91IZK
OLJdsJN606vcEHG5zeu8FXqb729cq//IhjItFsAVYXB1Eeq7f/R2rQVfVqV6
0fiP3354YwVUXvvx9bb7C+L+tBXjYZRMj5jy7ql93UV3JA/n/4H0ZFRwjZut
KombsqeZ6ZiYbT9wq8a7D4HWhFCY6kA33BXWq/WoQG9upDoQB+NOYygWKPC1
ZJiPn5lAxeFarBKugvODqUYVgp/xy8NLMzXOM7S+4YE6Q4T1k/LyxaWpmhoC
ZTyJCYUKC0S+nGeqgqEr0an3GVUOYS3B9Q3lvOjJNYCLbLNbXWS4d+eZHt7G
ElWIkgoDeMRUadhvxPLesI9CJNlQ4CiBgqi4TD2rN559Q0kRem7rEL0SU0vM
40rN0mqCW+wKzOypRYR/pIx68sFB8D4i9+/1od0gWkjcVqZ6CPjDEBXc4WdY
W2YIEM2KRhYBIXei59YCfcohuGyyjBoHGyNW2eQi75lGYmg0JPQI150qDoYd
d6t/mPWBk+BmizWd325pZZDDfPAbAcj4qD7csy0L5/O/M4RIY2BRqvoNDGww
SmzNBZ27GGnkLofA7YfYnX482hEgSaZZlA+bcrYZo9pWMn+FkqPRjer45ObO
M/UU1ZcPZ17VWex1Mu6j3uNkbTPEl3QAvXq/ubpxelTOab88S3SqH6wdTWCG
KiTrH1rOmPC7ZOhxk93gOke42HKPjT/yD3OALMQZx8S/P9NZUt6F0tjpxQ2h
6gAYlMyHusFvxWxxs3ftFiKh2KhY1HwRMN+Ned25BxrDQeXgiaHs3ffBwhdb
a70t89bNcPsP1ga97gaPSZYVGPhLjO/ty6yhe0M+Le5PJTAfDZhTYMbdWNLe
A9rMc4Er2gyCi+LO/QYsLZt1k9QighBFXC140cDphmIxf3xqn1MpZf0CidSF
mkh8PShtcbnCtv77k2vgiqjtNOvd2DJWZLjGHjh+prmRmTSPVHop136tEeR2
xBooiTkdEu0MutrWKUG5gP4zcgfRSSMnimt9HGeeAZ3PdvJxsB5oCdaXtSur
GWWvFaMUSy+hfQIqdqRG/z8F3kYgpCR5FRIQdVHkkxBPoJujC58P2Ym/1t4K
hIzbPYQA/UeIQ2FePPRmqxGwDDRrosPIRTuiixT0klgrtO5vxcqe0vnjIXAE
PGBeFKPcztlARDEDgtR/g1uY90jZDMkPEMiSnTTfM1cOVfKdAlhRzEzrhpqQ
vFf9rcS5j76HGgf0fid9APDjTBIf+WJodi4mflmBhGB2ekURJKhcJQpj77bI
25aByAG+P00dz8BeExHl0wQ2+cEjzH3Hjrdcg6zxQZTd9v8MB3kLD65/4leN
vMNuTwKpTDJEmdQyN5JKvCv9vtW8DePE8pZZTEHa2xAXrJYDyCUHJb6CuzBm
uVTwyhzXY7wb6d+V13TK9Do9C29DzZHBFgk9+m3It5c/xtT5+U5f0Xn4fD1b
AvS3yPcyblVCEHQrlZFbLDo2I6Wbkueel6TcQLwys7vLE/SaltJvirXcLl0n
0bvfCNhBMtcu+4ZGQtNSylnpZXNKduDE+NEJ2Xx4AcmGNW/mCzVoU6WL1TxL
ialz86UFcXUezlyxTrZg1T0nQ4VprqwCJWWphGrWxBXr5GXs876InKIFwxDA
+Hj6aY0Xnl9KSzrDhupO3u/pb5hlFKOllzttSKAROUhFasUQYB4rUl+/5QTo
r9tMEBXKOasqr6IC7t7DgsvxYb09J98IqPCGr4FF8HAfaKO2TqAvZdQfDKd6
rfDwVDYVWpXpa9ENWF2SbloGn11jr+dQXZ4ARsRYFjsPyY0rI/QLAZ6Q8Lro
AwhnVPqaG5koMfopoU8E5AQnycqRYcoNkZKM4M6aenXdwHXK4cHV/S+wf5Rq
moTmGge2+7eBy5PLEcVF02574VllTOaxfh74kTw2SR5bw9f6h7iCTsqVGLBB
MdFtzrAV40v2UIQKtp6JpcUicRpgcUbcZYa6l2ojn3oAdfPiHxgUratdQV9W
LEizRAiT0D3ImiaHqsZ65ry6BEmJaSXAvSFm/nBKNo3yY+UnNoi+LqoN6gp3
/yketJ/9zwLdZrd0LQWxpsSAt4nD3VAZhG+uMrGMAiaUYbNSGMnyYudP0hxj
uD4hthGCRoXvkjIMpSEbM4dHpKRf2OLF/1Qb9ekSWxYnHOkRiEgsob/BbOsM
5GDEa7ioc7KBsaM146wvZqDv9ZssAJAPjRwX8dJZ4+Dv9TEnYx19AqMhK/wQ
O2i0iMic8uGW9ClKCe55amYcB71Qeqez+QAKrTrkUbGHEpxWqjCTwkederq5
JHFqoBVN4NIFW9Cw8jG0Hl4VFTbDdXtcsgTP6eEE5NylFSL9hl9zMALwNTV1
CN1QnGK/J297oeBTRB+QgYpduVyrfsEdq82pAvVVuJAlJb/ggfwFEVLr8QGs
S2wH8RDNQ4XWbUrO9y2ZoPTYkfi6H6pAFYhzTmUlkgolABgG3IGG+1IG6Zv9
4IDbcWQzj/7ZcjS9kw5CPP8H7KjzaYCJcLwUEebqIWREr4QAmIAdhi9o1be7
qMQKFff4CFLRFGagGxCsW/Nm2MABNsWV2LBRfZDDy0NZJIreFFRmhFerKapq
n0pwNX1z2p55RN++BOZTJfL987TtNNuLHG1x3nFlANhxcrP0Nu1g7qUYXi6D
m3SfoHUZQnxlyfUzA4S0Bcz7hAH5rsiXxEHN76I9fbQ8+2T2yvkOyd/8/X7r
c871qK39XPw4zJ8rR0KvfIzu7EmbnxZinsAHs10hAppCYQjrHD3efQQMb8+X
AEloW5ZlJPlL3b1sswCi6h2wL1K1d7kv5yr3Vqc4p0VL1gJUdIUo+g/6zGuj
gt+3szrd+NZbMcRQMLWnKImNflbHs8m/hnHUoVMEZRyMzTnwmoqhr0MFa9aQ
PEj5BFPxPTf/VCByVy2t/YhIRIq1Gl2cvl83W6za8+E/7h8McL86/ypcGOim
5uIggtpkRXG0qngWVFMUuiHmFkCTC4G+bKXDQo9cZ5qV6OYjjVw6zAP55BEP
WQCY2Jg6eEf1dRTwnpczQ7x0D4JarlmKxn30HqrPu0VrLC55w6Z9N58rXM4P
eDjmyYTOR7OyWuNVA/Kt8RUlMnAxLM94WMKe72RHg3ygHA5aVY2yqXE6DZA7
IaBsKF3o4dLmhRd1Rh9QNVykgQvmj7+3jacjxLHsrVz+tMp5kawJ2b8PlkTm
y4ILeYWeHdaKkMGFrIFK7ktq9uApxipWs0cyPLVVJv8Kf9UoHPMkFTj6O3K0
a0T4AFgctWb54LZtA+KqWIbfCxlb17YVbM+Ku7Qa3idCeDMPVAEuShdrnTeD
S9VmYPKm/dd/LfWPYys7Nd66ssMwlW/U6o0MzuRSM2CHatMuCtRrhnhMgt//
OWYIGEPef+10fNRu4dDOfBBUuHmr9ASMb/uBR0Lw59VtoFYDrqEaSBWSNIoZ
6lseex/YJ/jygNJUtj3XsV6huAwVEGfT0oxa/5Iw/zEYf+Bi+awhMj+GO6vQ
bo/vbaJnb47AoF9TWe1cKen8YPz2BtJFYjWAulagudNbhAsfhDigFkEK1sPQ
brn/6haqk2+eSyW3nL7O4wkTCWlhKbdH5ay1jWBPbnNJW2JR2uiwpbsMetGi
vWoFzChMM1ZZHCEbCkliVIeZ7NQeEK/Ac1D2kYh0fHccx7eeTNBjmGi5/hyO
kggnu0+6IW8zBEev3IrpIY654VsFk16I/SD0W/0w2YRBBCMnLWutArKq862i
0nHVpvOIS6EQYWbjcgNK3spyqrdi8O9cZAiyNhEJHxy4w7y3EcILrlihJv9b
vsY5quIlphG4HuJVQKk9p0uGOvSwHSorAdCaA7rNnl+FMdVv7xOc3MFMRRGe
dTlOW9bS2PJnfd/RjLGMwO4Y6fEAUhmMNPfo5PzcAfYtv5qCKUpTJqrGka7+
/DzmZaofZE8c3SvJ2tm1jUe3hqnob8LUmR04bGBDOq2wgc/kT72t3L3pkvrh
y4/iZ9Rj2FGsaJLRUT5cPaUduROZqyEqcGjeLPHQZMkhj4s4fjzk3BBojp9E
YpHVZb15NvhHqsEpMea8XWWCsQf+cJFHIXvieZjFgc3eR27n47kWXL6DwNtl
s10ZULcHcQIeYsarG8y3tdQsu4ZO2wCgZWcmLeNAWOt5L6uM08BTZO/kref0
P3fmlREMDMB/qZSXJV60iYMqQeDuQpQKxs5J1KZlZgLDAf8aAL0UFL5enXRd
XHeS6eFe1OU+8cXqfHSrfm3NAfYzAayrvGX8tozmhXTmyM3Y7cnYiB/xgBJc
xWnRaShhHe1OSxUPdqMTxpDAMBpehwjo6crpWvqvm9GNKX/7ImCdTxTjymcR
9lv9raoENQ3V6wdMyq0Nj6LJiHxST7z7N80EXjkSxFJHXKo8IIzV9lZFevt7
JFsSVe0yrJNEbm/YqNyODdho3wIcaEJdZEHitneUh+GCEXph/A81P+XQL179
9re+DTgtEB5YIXJCESe20YONdc3WyxFZJmNysxYyP8GsWcuBXdF6fuh2qc3U
cVZLx4mD8pzTDBG0oNmzuJ+p+H7mMFJ1hmbcsUmxi3Fcq3OuuMNlBJiQC1dm
vmc8Y0OzS+dWNNYME88J8o8M4UuXye/r4T/QCwA7wKkIe3Iha/YqhLjJi9Ef
VCCotYVVbiKKzLvVUiNENrjNd2xNt4fSti4dgd/WBZChE0LWOIavOiaKPmmX
XpAoAMc6KR2fyvBRUVwonjrLHgeewJuBq1OIvDGaDU00Oi7eJJK4P2c0xWtT
CTyK8c48EuXMGq88O8kljAOuenanE7mVhsdN4Ob/e4vtBiT+5G7HI/IF1001
K8DcQFY5Rq8hFQ/aqYGu6SoGJp+0/MpRFHVA7S53ZwGcs5P7dS9hGjAx7ak4
5lWk2e9MJycDnETGD+CG3heukZYtcAzXxOgyd6OesmSkaDkduZMOIZO4whgG
dX3De4ecIeU9dPzP51pwfGF0HJOLk8hKJRARTZMVmtC42u0Y508R24R1PmhM
XRwbtnzrC59jONrna5/M6f7uUf62QGXRDN/CKF3jWWJXvS/6DDygfSj44dIg
pDCVRbFXe3RxpLJnbPOTDDe5YriViNRrSj5lXOKqhN+UcMWf2FH1+C+H9r0C
bVb46UYWd5eKFUpUlfZ/WPTefmAe1nN7y0R01si+RkHp1SfHyiIj1vdDOpI1
5CwstsaTv0pR8FjYD2Zu/sXgtahEcJBobP408eTP7I62fQ5tQ4ppKMn/QwOW
gwVop4VkCbmxS0CZRwp7Shyfbp5xhAoBQXHZsYOPgLg9tANmxpNKtHIZ6cWQ
KwV7sUciEb46Db5Nx5PUWGfjvwtRxE3YitLyIlGElWkr73HdIFRdE3K5So9J
k+phVezCeG9QoORK1bdxDzaDOkTW0mOeY2B0CZKEbYbfN4PR5qMF10e3bPw/
gFjEJOl/ZyWmXX/fTMUwyJR+FN96wHSTLBfu49i13McRrk7k1oD0zRBh7yVL
/g3oAylT5S28/GH5J0kW3a39/51h9CVi56qPV5KCkac1J7EfIdJiCoZ3yOrn
w8c6OyD7fIJPWq8eCG66TibZkMMPPnYwlHdB0w45QIcuY8pqditYrFLZ72e5
rhtWL+WP4PveIsVeWyFhUcE0k/Q5o8PTAhBLkLrTG38lZodOgE9UBsP7MsDy
bPG57HOHrqytKjMpBfHeEYgh8LYJfVuDD7SxmyU+BU0wBbEYWJnOl529Eyta
snvMPMnRPxk5jtM6NbZY6hPpnLm8VySi0IgFjbydthmT6R8gboAvciYxSFWo
4kgZe2QlBgp8QYp6kT/ovftO3CiwOuId2wt5TKC5jqKkyB2xGq/zLnqe1izI
d6F1hKUswt490kGqWLqOXNFvbxaW1M0cCdc5RdaKWb8UAcHrH6h9/QGTNWN7
JPG4tHETp4JI7CRj7nfTlQf3Fv2d+lqe4r+cxX/r+zGiosYBRHZuH2/S/pE8
pcXwbgM7rUF181IpyV/1j18Tt123Jj1am92Pau4DPxsW4hDXFzog4RawtgYj
bydlPtuXMUCFFI4DsdRamBefkJtNPF4Z3Qp7f8sLWMhsMJG2GPVSH9PJKxgr
QPsDbw5bLjT9RNr9qmS8M6q0IOj38Xl3FDNJ17zYcSiG+CsbmcNOm6G1IYke
yuKwcxlaZGy+rBRocqPY7da7OuZo7GdVf907SNMRZqbRKHnW6TTKytd/MEea
u9iPnkm0nosnlCoVWX84EfVFL+5jD/JVXIRtVdW0Y5Jv58giHk5sKvCKbd43
0BlvqKBcFZawqR0FIhRQF0+JGBM1UfRJycU/3CkKlPhPawpKlDAppAjQtmuh
GSAM0wAy8qsFC+D03fXoEtNWPOr+3ZOI8x7T0i6blg1nZrWan9T0SaqhQyJe
QnmbT8PsGWglZOl0rzA6idgpxjVXOdL8uY59VRsCGCbwUgd86aC9jrlhk2Pp
0Mzmb8KMLcky7BSyibj68viC+PXq6JiRaQbVEMgImQLgPehHhl46sDJQsk2A
sA0m0Kn72/9ip+4Z/bDrc6ZqEi7VQKjOLC5V8A/CnqqCiRkhRE6gcO/DjP3L
lQkaKK+LovUz8i0YgRuCoAS7a1b2MUItLCPseNK84Q8cYlmhjLwJ4bS3G6QZ
/gAkaOUnUc3+//ZRQ1QuxhkYuuHTqRnnOrTgeX3qz0qftsd2mSbb/c/BQfbt
1l0JghCDOE6AQnM8fBH1GQOoNZoZVvVPYexcFOWEBsw575NL6MpJih+gAF0s
oTeeML2WWGw2gWTTRs6DjbveX1vOT7JrFZjPePdWLBffV3/D1iyCBnp1UUYo
rSGzptR24YGQ63mnugRDwH4hfpkMNO1aaDI6yshz6DZ3Caw8STG8UUIS/5r+
/CdERSXTz95hNkyHjh12Yrl+o/dAaNsv+Xno1boh8pyrbiOUzZZ9jP72PEbX
jQNsRd3MMQ8zW2AckwL8Zj4yaNoLwnSghWK7FKdkhL81vrn2B4OXHl40gYlF
bbE22eBtcAREsuDi87EzAbiP/uNFdyCDUyppdYEN4LscUXmRwEUVk3WhDrZH
12GZ4yWctjdf/59JE+FKMGU/4Jfqu3j3ixk6NEnv5oZzRqQ7T86GgNcHf+u0
Rx0+UjkvH6PxuYEIvPcqCQQcGLO0iXr1v/5uOGiPPkfODhDpI546j38U3ZXd
k0sqklwlyu9s4TVeAn5FdGOIpBDj1WaXosohCFIXx39SNNCwbp6p/tK/N0Hd
bknmdoTX6KoN0C+6Z30R6UalyHL99AzTBsR7udWlAV9kjtif6DAy7ULCs9u/
8WHHFITaA0ESgko+ogHKyEuk5tZ47Nj9edP+yCav3+s8g9y6/vmkXmk3hehq
9/jKXnWsl0HL513erRhRX7rBosg0dyith5c2uTxNT1PfjUra15AKVD445k1P
V0GQhXpc1l2zCFvVn4zyAhpZ2UOxlC1/oToMcNQAripe+vT6br5MHkeUIaah
K+Vx3nC4JsoE1UqBStFEMr/JLlg3Wsgz3duQS4oq0NdJT0JsiW7gDBIotW0u
FH4GdllmeQa68NQvDyPmM1YpCdS5SO9hh+rzSCIk3Ynn695TZ9nmRoy6EsQU
Tx6FubY0k89h9g8wvQ0r7WnuU/eGqgof3F8SMOH6VV6N6KCdvzW607tJR0e4
8HGAEnzT6YpKN3R7dMsjCSgR+/wZBfD6XNtKrmotMKr4Hl+Xj43qX4aOmq0k
NNyuVTX78xAmBiWkfTlfEoTfjIeI9R8kIQ4urKlv/LqlnWrY/23BjGEYdBNa
mDebax3PPBtZR/UfVwg8PCxVBD3l46WgkckUOLFQtUwfLufTgglhe/alFaxt
NqISskJ/vqsiVy6oMrozh4xI+r1sd6lqjT4n84e1mzfjhBjyCc+NgaKUd1ds
65l0Z2/SBcAlkjO8Ekds7QSHeFQS3JhvZAmHWNLCEOdEAuL4UPuvSz0PJ4eJ
zqvba5CwF1qdg/qxkv9naPdgKo0Px7p67qf9XgMXnlaqGlPWCibD/3oov08j
Tff3xlz+xOy68gTmxu/B7si87Zq3dUGG5Xd7/lE4qsgzt7RNFC2xz4ge2QSx
kqq0ec3z5us2sZU/mJqiuKdUKJzlcNrvWSSDe1mfNaI8z6q8Rk4DEiWAX57S
SIX7qkpo23FhMUI0BIlrGMJeL/qfo4UY9S0f3es9qsr4k+zDjmDvGF2BhUcd
NDc/xOW2c9tynUy//0p2p99XBMdwlkP18EYMrTNdIwV3294Wo9gV03izA2Hz
aqvtSyECMgk/fIUTEVqZ/Mbp9GREmEozL5K7wCBP1b8ZF1aS4nWo/zpMWny5
jlLGOIL9lJd0Epix0DzDLk+FI7FzukhVu5w2ps3ok0wygewzi7JiT8+98mO4
G0Yu/3ErBGNs2gKktoGKGkRVq4psM2Lj1J3dZFnTk01ID07EbRQ5ZxMXJnwy
ReGw65BzgoDQLmKmPTt4Ht0pVeaj8pVTeTlqxs4wJvWXmSvOZNLZrR9EKDbf
3lgSBztHNtijiuig/sHUEcMcEqVDaa1heUltgKRBmNnd+21lR/y7hyqnoXY+
tzpPhjP01lO76cz0JaI68dINli+ycDWHH5lxP3vj7LiQ+6D9EIAt7UkHFek4
gg/QHPIH0pg2QD2u93xcafRmv3JK3+zoP4sY7IA79VBgyL8fCfb2SOfunmWJ
YLZJj8YGzH9tinQWhQfPgJkt3PMTtN5TW3VcJNL3DX2paAzusZwJbgBQlaWC
9NSiq0TdIXCMaGtFGkxJJKae0jnH2KPU8ugDeh3k49USHEtBk9zZrkDE2fwF
5kxQnoa7PRvw4oBVDoudv/a/hczkH/04qnqBOLdUJDhpUfBU/3Z8KJxYNIKZ
wapkSLkBWsnP51JVGX2LvAV6SCc2RZwvAlLr4OyP7W2kB48I2vqQvU3Icsvc
QwqDQTKP4a5J/D0CGdYhNTvOh5AD062pdF1m1YK1rZqk/9zNPL4a3cBPmfdl
Nm34ZA5//hfqQVhPD+kMUZQ3epR1KUk7imnOH1GjAh4NPEf6nTKFpM22/cPu
dySL7A40b+6aZwN29Yz+SiMKWcx+5LJtX/826cOJrcHfwgVWHnVYJDKAMeNO
jy8od52AHWmMNUjW8r+rU2TkurLOKGkAk3Ko6QxBmitZEcBmXyqBoDRTCJF5
5sVnhc/wCcJlmvu/hGjrAjNNy2zEQV8UsS8AaPB/yWT+lhaQhhUCeC3vI8Zc
Jkg0fv6mqVOpr3LwtzRpFXCw7xwWLTrmHcVIXXUlT0g7sLK9iBBAJW2Qq+E7
nA1cAKZwWpq/4PnDunvAxrloHlMNh1BcIWISzthbVbVfQMkg89LTpWDD8vqy
XCVoo/+xPMZ9JC7aCYpSEHfJPFvUMrtuMv857jvE2Y+Gu2BRuTxd63v75J57
NZhJHZPP4jRQugjqQFONkNuiST+lVDm6+dxUNHpif2rg/4Gee3bjHN3qLTh+
Whu7S0He1DcPd6v2Svqsrhq9Ih6Xio6hzrKZ4QZCcL34JC29HLxvu/DPmx6b
Rh8ezp1rc/GjsNnxQViC6Py8GG6M7qyOodTG3gTpZXbuDxBrOFi8Bvl85zYg
h48+q9A1hREzRdjzc0Yhv12ImMKknlYSBDZxG7ck4EX8lxnTsed7FArt7ZK6
v5ft4lUSiw3d7/PGiDW6XTxcISdZ++SUmnTuxbktnDfBMIbPEyqAY54eF6do
JpQRfIDQ+kjpycd1+eEkF4ZvFQQbhhMTjPm4ZdvwyqZNi/bIzbg/l7/aBcB3
YLIcYeprbQzpWKnW4yQRSR1Ejt2iWtP8ShqyxO7Bd4Bs+oFbQDLCUccDygNZ
8RR9+C6vE54YMKIab/Ah5Dg1oBFKe1GxaaseqvwdbGx1Epaimm0qHCI6jVk/
yDdZXu0hLxX5rfZWIhs+E5zSOT4NfxGZIWhK8tBsxxplONkVu4NT8MXlB1Hg
zPr0rdB/Hhoti3qnGmuFuEf4XNeBFalD3Jx0BUHV8j0NJciyoaSxC+dUAaoZ
ArhpDsOCcTqQa3vQdPxdZ7Eh07xa8v16cVXiPZhddjrZOlkzIyGN3k2amQxe
Z72PS5wJcjWUxQ3pvFeVfvjn9gqyajR40mnZg2rgVFDPTZFV7G4eiFIHajV4
6rV/9hz0lyCplm7s9J3FA34IWqvdQoktAyh2wFmCKOlLcxfg0Brfbf5NwOoB
FpWkx/spS++IM2ISgpmrIJv384EryEPNtsPlDxJ9iyHQhs8h4CcLXLO04rBQ
RjMJ+GTTfcAQRiz4dcbngjLnJAIu6TD/+kQIQGOy3y73aocTyTVNDmH5ZS2f
Rf5GWWE1l1ukUiDNAdW/rJVjx0od3r+zK4tbW9w1y8l/NBdAhsBxGmnk+Ssu
s8UwLXejTvifXYlKb+5/0zs8Msa97y2hOoHD2buiaZ8w3mEnFP096cN4RmjB
CRaYlhBBRj5LoSoz4RjBmjCtHrMO1pCLR4eTO7/qQnVDn1QXFbEoppYPQh7m
AYKVghq4MCYi6mn/hvyLXl3PNvKp/0LYf6/aDxL9lJBrOjl3TepruODM//jF
lggwAJU2thUPTm4Ku9oftRdqT5Wmmic2Z4BJWMuV77KKqZW2dtH45m2Pj/Ez
hzsDMnGGB/+zE8H38Z59UuKF1rLm/BXhl2P7oWg9dIg3MU3/z2obHNOI2A00
swBB347/wTRSMNVdGNxTUPtsSRSALUwcOJgbZxttTLXBYxWBLvyeqTXScn2V
j5JXb5M0SWjQHmlxwWo/qKeLgzbM+vB/TzM5zC0e1LlP8xZfSUmiomTC0uj8
pzaAFt6zUM/zwxUdxgG1iRMkSu/8gEVsGRIDtboR9tLD2D95jYsD5bEPA/r4
FII73XK3zkTslA6zZNqAVD+j0J5fE2E9/BAXx1rOtX3ap/uGTbSTLj9Kx1pA
IBUCO+bOyBL72Xfe6xlIxe99aIjPV6y6/VT/2AOUdo2Gw+8lJl0Kw2yMYhOe
m86OYBYAik0StYbUMZXoSQMgD7AOrL7MO9RwGkwFeOEuBa4kXkB1NalSEaLY
1HSPtUbCav0rdMOb7ZH+qizAcPd2ZkkzbukkTSbc28uB2LPbJHdjJiFZLXx+
F95jSp3VV8E61QATlMUAe8XzAN/rzf7WfqL9rEI9ERAWABzTxVxrmou4gbJZ
rDUhIjactPSnKPd///YCDOl9lpb4+pv4MfHE1/df16Gt+03VHtAuLjsF7l7s
x/o59gUJnpb3CUVeDrr52exYKPYELWO953zwUZMT4GtCgkX+UsPFTl4XK3f7
8A9XxxbhPyy8ATO2kyUu6K+9VzSZ3GCurQ1dXliRCP2+uiFEObaLX8nS73i0
Fzo4+s2Tiu7ZSwhWTt1GyhXpvKyeXvNKMf1Dmlf4xT55IFLuRMMKtzakVPOl
3S//fkxJfscl3WDzUEahSzaEwmjAAw5vlzvZHJ7YUAFoPa43Q0Go/ksmqbPg
B3AXuaCsO9hLF+GEnhImV1uAJHLIbbF3zM/nQdlud1msCDaeRD23UtH0wbIC
hVfo9t0Jjghiaew8aOb7ul1O7mSzFbBTP97xiJ0HRmBqFmB5LkFWhvTLSyaN
hBSQJAMzSf1KDqz/V0C3po5SR4sh/7W0Deyj/KS47HTVgFibRZdACHGpwF5l
NIDPkUPw+27Ah5ENWc8h1IYmsLk8OV6VEbJrLYvKkfM5Y8IXN917jXZFz4p0
aa4HoBnzyZLi2uYd+QCIA0keV/12HiHZLXzyDKBWWBMYM7mWr2akUbp9be+E
7kx7D505/wPDaeZ7uy+U5o85qnqTgTzozwLM27ygchg9uEuVvuFdsjjHJQ4f
mFku4Cq2ydcFJS1wa0FdTLjl6OTgUmGN8MQpSaEb0r1vdJ97tDmfnvdcPAYa
oIMC/aumorVwYBA6br967myLYW3viF7aM2Fsyr57ue520o/XCMueKAEwvFA1
w3SNU5lll0NqqvFgPeSBp7TTwR29KLYK4hew+LMdhnlLGwIvGyK/goqMH3b3
ANJSHKDrcivSMUfhNRliLIuWw11lMFjNMdj0fKdme/HmnM5mT2+dVhosBJ4y
VgdblKRO0DIKEBMkOavTRkzR1RBuRJdGdyoWZ6GmqP0IsqVcuf6Y9ImU+WQT
A0PyKos10D9sIL0VRq/Yr/KEjCgpQth2WlTqlZkG3vC4veOHOnYWesc96494
QtZIDobgwwCclDbVXva7qnIvOlvhNW4Q/1u5VA6OZzvzSesqajz1Wzzp0dma
uMhMC7p/rhgYQtJTT/jxKKgEQqYTEY0F7UIbYNm7IYYeTBEJLIIkEC0Fi05f
HOX6nEBebYdI1tvCwwS0B9bxawSfBkzIMxJAn4/mGq2HU5aagayev0z0dc15
HwFB+s03jifik+qo/7Gph+8blPUFNynxz0RTnJCLlhqWx9l+Yqnb/GjzxgYw
bUmRASDu9RtiTMMNqs/b0igMzWsKiswLID6dLk1Nz+ggqWam+bkxSpuRkXjG
50yd3r0xr7yAB21i3dPCiwKgPoIOnmoMtVlsvsVuMBZmplj+rVDJywyE9tHi
3jnsBFuq0X76/XnCBmUOxQwvX57IjSNDi62TUBhOaQU4xG1NeK+vaLzhKv8a
qvegU1CC5q177kwhcvoQQtQ3Oj1ZpdSFZoo3GnALGQNzRPJ7YHB7ETyionyF
3DrCfUEZpjZ3lpUFxMgBcLxDHAiW5hotjzrHPnVJmJyLISW7QiEtloAP17u8
nik8IAYX+Z6BHtT+ChbjwrXb7Uc1b7BVlUqhuYhigZ+U9JOVlsVEgrMRfBHe
lvxDfDJXLD1nZpgmESZhLnLlTYE0oS6AM8Lm6YABsFcXKlJDiPsElNtsnnCW
D9n3TtzriWGRloCDkEXu5Fxfkuffy7VqocVHEAb7w7J4PCkAzwBUfjrJZnYE
fQllpdZapYdchBg31mbvv40qpCq7uelZqVOCy+swvkvIkgcjQeWCvOk8Ma9G
XhaR47p9JMZgCNTgc3g18aL3gkFgrncHW7aZHUOzJL5e9befll6SByTBOUdT
l8WowZwnPtg5XMGv4Kpl7yFKDGDVYznihaOi2WAlF47T4hM3aEyojv7MUL6P
T4zPdnVMSCrhwC5CbkIUBIdona1dLvqIam16c0+kiVBsyYuaKKlGtgCSiz57
xulKKnsUqZGm1Ix3GPeonS4HN3JjpaJU3G+tehyki/3qfDteiEwYr2+tixRk
9BYDos5eU0AIgYc53aAKUrK69GaG17QRDiEnSDEFkyV0cm8wY9mhPKFAukAY
GVNFvL/81sNimReGPtgWTdgRbmZiG7EinY+gMOAMtsWfvhECEDArNN6OPqSm
L3dyEmqQOgY+ubvhTyBU0s17q4/slB9UzfBGDN4+TKD5YXoQi83MbkDG6sW0
fGQrsPoeF381/2oZLjITA/Yx/vDivHdYkIHerI5V3G+nZp/aWaLhROC/bxDW
THoHGlIZqssbhqq/Oq/xClNKYF0se21pBzu+xci6SFSEAzWrPgtmuAFVkJTC
+qPabNjw29CsxzIcr+4DUVj538PiDT61aSGRlq7Q27s1Xw70nddfoHAtsSku
gPood+Fd0X9NheLEq49eK4F2xBeFLM3bjqW8EMFQmwd109M5SFauiB467zJY
b3yA4YliMseo5fLensLUE6+DCDxbxtmAInixHa7nkU3POc01b63U3wLj4br5
i5B0cwzp1r88iP5vn6sEQAeMbFNly0qt1FtcTgQv78eN/lQFfanuzjWCF6G+
7FEX+jctWmKpQ6zwEmymD+eQiWoFYs8kfiVXC5chD51+Qv+91gaHRxkd/3WO
rYt0/AdFExZ1vd9pW/rPVntrFcSrRL9DCn4tvj7dJQWJdE0cs9Tq8dtH9qVc
cBXyPopESYSENMPLjMYSz1761/uSZMU2KlQJx4vEpToxwWgmULAcucg/A8wp
0tYzZwWnMZ5OAExDcSwYK3FOaNMZVSUp4TnFAiXpJScPiwPk2Dx7XJiDBO7E
CWEP4cNYk9yawOZGP607/G7LUCSwf3th1/UcI+9VLxXwaID98ItnAk74TCOo
wiRcra8hoYJ4POQE1FEN8yGE+VntwTeVNGoVc4JeG4NgGJ84W/VKAkWF3G0E
IdXwnHavAP4b5ClsljfZX3mEpZlKf3PpgpNxL9AtcKEfMP1+6e5nBgZgwDic
7wrDTy2JaMX+u4eGbWsA+N/rDgqPzJOxLng7rFv1BwGZx7iHDEec/8aJPTj9
mmpjUijPjm7Kp39g+wZoFHyAJW6RziO1R+wHrm43xiCPMnXlaNKVOUEctR+z
NsoqEwkgIC7bjUek1gmD5F5FrVOfoj2ZfZuiMB1OCJUOoBPTBpul4ibgSiuX
umhrFB76I8sRnWjapcOu4FiRuL+dsZTrOsc+StA53uuIebqydGturvON0yit
jCf2eErDFAz0Auyr9GNDqQLW5O0G91i91duaigJ1blKauoMN5c9NQgRAsnCK
LsJ1ltsattl3dSQiTnjds3W1gyfGj0MNJZ3cMV7L6VQuCbArEZE2CdYBFvdJ
N+yrFCRsf9W8UJvHoFewuQtbbMJSX0/avaq9yiMvKYXaZX67d0YLcsl5Wl2A
BgjV9IyqBagBJkeSsWy3k7HFO86Bvy+UzKJtJ01SERXajlPW1pDCAag13T+0
gqXk1e4EqMf3fejPoUW35oss64qvKUx0LttaeJqyoI7ObimxM/+QwpMQGnyd
xRSvhdIXWDq1+rcjIV5toU+AENap1yBLkSURE7A6x+OxxyNpuheIKBZn+QCa
KdFKi+4eA7zd7H3ojXCHOxGD08IaN7M367CjDlPpKKLX/eeMXHEom7q5AFWN
ob5318lFEELLRUNj8znCNz5cOuCFj64J4pmCp2fAKfzZcBTwz4eiijk7/mu3
VsdXvsPNLxherJBBDHZIowTDix+23YItc1fN1eJmcqgu+kvHXPFvY/DOE1M8
cuah7LaIFPrLNLcY4CF8LBzPSTNceXomVF+IsFJ26ZI/1u1CpTxeMOXd9gjp
np15JlBJgMdk5N+Po71m/cRxtbhMJX3thhNhLE5LFItzq+CwtQ5t2HZgojO3
fb8k0GNLh3YMSY+QgfQXM8VTXPqKX9oRD0kI3uEfVOHEmemM5gR0OxHK37Xm
Ny3N37Y5YGiJjrh7izDU2RVxnrZG+Jx3VMGSjLmVv9iyE6pKpNwbiy4Svzru
mfptzL5QjFlHeGgcbIaXzQpPBov6FYtP/920Mn6ndYNYmzyVsxmv/8+nP0HL
4Ki11Rg45xxBRWbyZZzZUjJocofJ9gJovuMfM+1KQz6wbJjWjV7ZZcon4MB1
GcBOgStpcEopEb0j78aJaFQYdH1xbltoWMA0YdwSjti16v+sVR8qjBCGvrqo
I0fJA9miqTSQFyaBmJq/EDSGg7MbHjaHVcMkxYAMz5XLRHfEmuTW371meNQp
i2dyoKAo+MfZgfGL3r/SyIwEkGABCwUYhpD6CPPbZGxTt0djgfZnt+YNlRCU
pwEKBlaQVLz6pYv1ghzBhiA+gu+EJERbjtd0mvDiDr3HarMAkoizMbHi4O/g
9v6lGj/CZoREEqMEsTsu5LPRCu0eaeLWsTRhXLDgRt0sBKcfM2U7Lwmo10TW
tJ0VMcyI6CjAAkpQ2pUf6XrBQsPxerE8nSx5IV9pMM3AH3qGCKRoO5kxk7lu
SusQE14p89z7wKgS6N7ZP5IpPdYi9uRpS4GUJlS8IR/4JIdrTcDJK9BWpkU6
e/uZYLMST70mjMMtDXDuA7gh0dz8mrLcw46ISYG9zWHTYbJE03phek/QT7yA
8Cm4kQPazZl3E9Vd0DU85mmrov69/fK5lNdhRMxoL5vofyoR3xvu1iYBITrm
oddpH8ETbRrK+qdgBwE7y+QSW1oFamsK+XlCZBkbTKOR4sRNvnxssoR99QwF
LSLxI7pGdWFFZB3LiwGhzQOObSIdxxmLOcuAgOqdyiO+Cq5IWg3zr77VwI5h
nMxMVJtsIz+hUFL/Z3hTxCdcmFcWqT4w8ENPN8Kvs0AIb98h+9IGZtU/GEX9
TN6zblEUWVVkxb6Eu7pHIdGkwc1oyE47I7xWar82RjdvCrUTWRtHzuEtRzTb
N2Gk7fAZ0pHofEujtWSI3dLNJQ2YyvNq8/IHzsHhLPJAqtRLOxNJuwsTuFSF
e5eJ0EGU/1/DQCIZbPkEhH4MDKZWsMFoIrjPDzf+YTlOZxtzb3QsDsg1Iha8
P26yu7arNh7IWIMjUZM0RwIXb/KafoQ4SQ0zXL3hzEj/u3q3TQwOrk9LtwB+
fNwNPFN2Q7yxhTFkUvW6TppJNMx8imqFmhxachoJozgpV/iFTzPuhY7iRuta
SAAw+g2DHG3VwkMMAXWmq5y8b212gKAirgveTnKSQCHet7pM9ssofn/JMKel
8C9V4wAdH6jde4VCs7i85Mm1DUCcDxQdmyH8DUGDcbv0XMix1mys1cd98lnC
sTLV4L9kOtzjdhrZQqZY9+wX7Q5h7JurnxdrfF6yb4R5nWWCwS3S171uhOmC
Q8wPoxARUKI/DDM0M8fq5gxpJqxLisnCabJmAkr7zXbxFMTMyHza+UFclpmm
+Pb2W1Mx4281IQ4aIo2asaFNrndyyXd7E6v+vVE+c5liMNHSamhd17MWfrB0
wR0OpvrJJZVkULEDmhK4h/CKeHPZNP9xvb1RIQJkuIRe2qegWI1Ih9CeX471
HyTJBR3MO9AZs0clfsnCqsVD9iatUriUYQcSGDpawYlAumPCvShkBFTBRpBk
pOBYScE/Y3WrDR297UTloM9f2FEIvgcXTSDpjnCOTtk9/qTgu7wI0+rkJz6b
vZg4duhvXp8ZXwW8bFwnwfq5NV4NMzk5FgdXtoQodXY9YZ5UsHwhabJiex3k
xyy2BZ5WNylEvyBSgdcqyQQ7jm2JpE/6Ts42tTe5bMQVvaHCFwlCwtCA6rXk
mFHmyiTl/I/QjrSEHWtbjsc+C5yx0nGqOJrPvh+HvAmWB7WX4AqQbhWdudCu
2zuK52xU1ylfxqBV8bk85SxykfuzGrwxHL7If2KAw8JJ7VY0dXykcT4Dx1tk
BeWQBHKvKR7iaQC8sDdUqCKYQV4psgguvPZfygeOrRBgicK1NvJE0C+2hR7e
WFg6WUbec982egOJFHSuVnVlE0oeojumwRwnodnD0LbSMkDRyNUfdjIBpHkU
jyH9vuBryfHMMz8EvW2ky6rnkzU2/T/2t/XRxFsRA1WoPbSI9xEhLbj6hBv8
PLRCaFA7oswQETxOjO9Q2Lcm0fb0GxyiK7jMuGHvgy1093um5u7dK8IOsSIg
1eK4wI5CZewXBlpPB5lRSDGEjAXVKC48GjmMUL4EkISN6wNo5wDj6SVPIFNH
Xld4lr87dE8di7fmeUfu8DegE2DnZ+id3JKm6vKbUsu7hNXdu/kVQtZ9cwRd
QtUyZYUjJKRT9Rbt7+h7ajR0vuBvyu25YzESAchA/m2bHZihKz3DM379QMZ+
4amwaKh1HOAescJuIBUsO/eRMNmVHcG1MgpigMmBwPCCdVJDa3coE17WG+F/
L3TerGEEIUv7l+Q2f3u9NmUEkpUg7wNvyURWqxD5kx+w2QT6lj/f1h4bqWma
MZSz4uYWq5T87E+0naS6cc2CdohQNPe3LyMEx4MLXmLjt0/N8zO1/ZMCsBUj
C0FLoOaVPC6qs8nmUfogg/FrN7h0X03oybod5nPmjh/uIcA6WeGn1e9467N9
Fe/9ua839+rrk8dVe097JAW79wD7O7ti6b3Zk+oFsJIs0y6rTp82ZxAqKCf5
S5CZyOJ/ekNpc6CVU8B3G4ZYQzn/QOBEocC3IfMvAFoeie2Xgc6hMEBQ/IiY
V2V3oMXSU3KrOQ+3p7fGnGLLVMBxQkTx75XeMGvDTskoe+4D9FRnCkW/e9L+
T8q3UpFyOfka4g2MxBzsOQR0bhzRFavKZHUnz1PcY62d4d2Dog68qq1Lsh3L
QR2mYA4b4Z6Q4eBY/na8VAhvKad4wbzDWxokCE86FrjWbGi4ekhRKoUmsOOF
Dwohd6+Fx/bj5fh9mLHTMPQ50yXhJB6kZH6QnuycheLT2tkkxcZ3mLvVo/wW
QqD9j525ffZRtYP0cmsxh9BckQJHM17GhPI5W4Q9Ti0AJhyxCfBbLNRhzV2T
69X76DeiOgma8ZG9QGfezfuOQrWLs1b6gKdeeRVYA8Bik3SMFQn1O38SBpEe
zmiWITnsne7ihHrp4DYkRVcKwHjsfkGzeVKzuwMGSWH3ErYL8xaEVhro8WHH
tlCtQLSzrnREC8/PqXtOcMriYzpO7pqs2iuZJCC9t6hybriSlWFEdAl2tP4h
s9+2bFixDnhJcewc19vFePrlfXGoIZRo5fPtcPH8fUD0FNjZY+dDUvVMnV7V
h68lAbQm5rBZFwJa4WKnSqmG4yLEuY/LQ0IBZsjYwtq0kT8L0aEpHCzAkN7y
+930rZAllZ2NxpxRcLw56qD79VVRg/TJAL7zXAwq/XaliHKPL6fHcSwAxnET
9OWKBmt53z3ZFMKGvNtdsKae2tnuzaSPLVhRgn597bLa0k1GEuh1Yj3FhFEV
f3N7dCucNOY7IWtVaz9a6XFL5xmhMCpQDM8ZX1mPkOnCpv62K2u8ejELcr3H
1EDCehCPLsCeQm2nCevhm/upqA0Do6i9xCqgHVNsvFI4H4GbDmKD+Vjqs+n+
LZX81Fbln6nzxr9z0KP3IxkNiOjAhvX6Kg/PSGcAcWW+yc+bKWzq/DIquGfl
J6j9JftqhB+B/cDdp0LfB3BHPbKqnCwwUpPdElP74aKJBVKnZObdlf5xSZrm
+3uMcuJDo1Pft7a8trVHdSzS4BFkS+qGC5sJC3ZB+z5GSc5vD/CRIuTeBgpo
6FNlTGKXttfmih2NpEsYCwoJjQ4+SQQHIKr9onpDSVDz+ys+8Kn9XJvA3pO8
biS+7v2mnumPY8H/qbPhVosQeVFONL7phS7A62FGY4M7j0oIC5wjgBaE1wfL
b06/3CBr7hyrAj86HP6T3PF+Y2sv76mf3PKA78CfgRNIP/kQ6ic7+sMcbN4b
WyswQ34RQXKrFpO1HfIjMgq5UwgOjNWJJoQRvoNagAaiBuCuSBJRtIls27pG
h/d9cKr4qsIELNlQiovQKyoOQoi2rtCDmhW1d4NtPOrXb2BkZCRubIlBQhTc
SATng6cYWCOPU+knToBLNeTgLpqA4PKkzTcv22YUCt1Tp9CdRLA5CtSlRmZ0
iM3clCflgfByoR9lHOmClrZ5j5+9C/VjRpDTMc4Kzvm6cXBrQW5gVlMVoUdp
GDM4NtdfDu8+MWrc2zjlBOlHF4MOnB6uS58P1nFJ8bN0y4uVuldfIqgjg/qs
QGENT4LOXYNj3vFGMnajzgu7TXX1EUCSbfER1aFpJ41NJGpPhExymETC1uNE
7LMgOJiw8A3lXP4fwFp+Lrwhhmq+8hxOb1ERWyzPGZMbmEFlEZ9UKkUoA2VP
g1zjKXGpmi6PEj6siFXU7Kd5qnp7eDV3pxEvHvvEFXksmh4IUPPWoxGu0+p1
n5HPG3NCzdwWbWkTgkMTHk/qzExnQvm7ag2+2QQdcfwvGlKmuXWunl/8Zxx+
ZC92A/t7h79+nV8NhzC7nyziCthcV9NmTJUzbVR/KB6wL3BmFnA5zk5YR2qv
M0SO0+EJ/32UhARoyeDmm12gHWFqFOMfC4W8VrrcjACSXtZUf7gK2P+ldjbM
1A34j0tPb2oZnhS/84FQ3HzfZS/U+zwe2TNaWHbwqLix05FkmdgvY8VFdEAW
f4WN59KhxQlSL/M4C7D8gxt7jtwc69NTx+wNemUnMsDv0F+XkdoY02Q0yR/c
zJHdHdWxIx69srcbkY54LNhkjZuy9t3g2xgCm2uG9nj8CkhnsalOlWh0o9u/
MDxmzMGpq0IN39Ps8M+aWKg0tZmbURBnc+EOyhGFxVdXeYOpmiG8DF/XHp8j
BR1vayWjYYbCV8DU79l2zvO1IkXKN3reNGiYolLkL66vFzebmCwJrkARZ08k
E37z72uW5E2Vj5h1Elt/FukVJwGAMUC/kp6b8opMFpEurB+W0lq380s58qHW
RlEKc9vDYPrWb4EzhpEdgk1uMLgXdkBK9Y1v5MErJyfTCuW6xpR3CoVocyiy
rJ6PQAGjqzScdxsnb+9t+0g/tin1We2W8OUXdgtCf97W5XmGGeOJbSposx/b
LJUrEeFnUx/b4eoDZFgIeWOtfdaZGY1ykeR/8SM4SJ6XV3zHa3/nQEFgRXbW
edxp/LPDWP9jub0GiT5uMlG+yZXmE7NruZxNB8KvCxxkVUNNr5pwbfK4jEAU
j45S2XlMENbJCv26e2pv08PmgunlaqHJdfHt+cQTe6eIyiXOMBGNejGEjvy1
plJKuYySsDpyR7horKVGoe748AMPojJvzSkZP8AATav7gUlnsVlpmVklp21X
FwaRRTVGLAe67Sj/nWPIXJDvqD0jmPTShVLzcsdKaFfnJDmDRHRhgk4l63Qp
awMnTyc16C4WVTmsLZWVtJ8EseDxf88a/276ZejQg5Y2t/HFbFz4H4s3oRXZ
HR82k3qdBNwPzPNVJQLomAqmyIfLRVLN/pB3soC36Ig1pO0wbReQX8w9xaJD
VABHcqU3MO8sYgBB/0rES96Kx8Z+Nb5hbS6K5I+opJfiTZ43LkLORT9H2+dy
cE6NHcXWsy3f5mT1LGOf8zyjTajSKsb51TXcSSKj0382bnvf8DG8Gn8+lUDP
pZVDLoPpIh06DObXDgJnvYghYwt+B+NliHXOMuXXadXpUU62Bztoz+4mUfPw
OK648aQ8Tj/5IIVZGiY6POwwo7aC6dY+Fw3hFpcs8P1DPvXV5L59rKVFzwWu
ETN38KUZ6g6dM/e+S2G08azRoxtKo2sd3tbWK5gWDU5N++NzPFR3wFa0T0za
ulUkNiXBXYXD+6CYJXaQoebTjAllrvfYhthyvRSy+IQpmFgumgE6yT/W/GoA
tr88jSU73hfu22dtCmVF3eBl00dwUYg7VvUHE5l4d8+IrMZJZXdigPnb3PKU
XH+Gnrau+aAHmcMCjD9gGp6SDrZ6xFGQ7cbS1CKgsQn1ryYCKvv/6wit6GAc
w/+HHvc2LUMG/ZaxAmTAN4+ih0EUeVlavedoQw7am7mc/douZOhvT5Va/QxI
cQS4DEjRzfY7K4MKUZUOXLqj/OQU4jJd0ZPiVR6d6+23Dwu+30CGjJZATtxA
dqgSz2pLjuPOH+60422zKUnV06BqU6DnAg0YLLOVMf6eiAyjYWyWnse8pqGl
34WfTM87ynmD6NdCt5SHm0zWHL3pn4IZc5UYN8bF6HnfboBbexmYsXNNiHhk
8LBZeEtbjVnzriV/g7IgVlF+wThPnhYNIqc7CZb8P1ZiygLYJ5uFP5VwldLG
MaDb3GDAwSHwWsmCtoI02CKEX9o50wSWERfB03tra3b8iU+FkIJ2vD9NCAPd
mj/+XkTPzKMz7ypNYcxtbIc4dzXrf19z0kBhfbwAzUoQxDHU+WCt5XSTDJlK
bLPw5R7VZSgzc2QLcPCV9P+usEqr8FDDjC1SbO51rwgqqKdZ9SyyHDxRoGEr
5cAqNaYsugTD5L6qqkcbc5aj7uQQl7XytQqsJ9HuTL0HljX9uMM99VRVQHDb
PEDAzxnhyZgA9IZOhl7ZKY5e3ozx0GDhzwJtHARCLGM1FawfUka/qLrj6t45
Ve5RBeorM9ZFNeOU44yyjHTHhoyy2bRRHdvnDmgVaO2f8fa+y9YpPCaCiULG
KlOo9jDvsphFK1blzJf48i8FevyDn1emQrf7vsFg4sGzymyFvHZ6Q830Ey+Z
f4LIiHa94iuzWn2I5UPXGiro8sWZHX6PPwfUVVEakdcN7zYfd4JnmqbtobC6
nPLU1KeZ+QI9cjmTk8F5I/itI8HqVOZ54kCN/LztQFETAd479EDUOKtBRHDI
7CED3qB47Z58k4uUDdM+vJmxoMLi1x6MIR0ofJ3kbPscCT1kLaA30OmgGXI7
o5a9rwB82enmVX1DgGHQrKPsXjhvrRknB3HimCBdmOUDEmqYCY7wp+CKEQ6g
G0K9mp1J9FNTeXaUPSUTHgBlOZYqFw8neu2DV9lqbAM7oo8S6OVfBJ2zXEw/
bW0sfG6DDvof6O7Yb5LUbCxnKHAaWCamPYqbq+WAYmZIOJ2Xg1LFHB3mM78t
aFWs+gPKY4dZsoQ1Jx6JWzDT1vVRyOvrAe4MWJDNxVA5/xor5Zf2q45GIMiE
dpyNBy+e6QSHlTegXGGAs2pJkNDiNZhsB/7YNVgpqVQPVfKeugTh3n04flrd
X1Ll8DpuXdGWX8qLTjS9TRUSj8kE346RQeqITcB1cgzk53+leLK5mHBBZFxx
XxdMqFHYcXVDrZhFO4TU5CN6Hj4pKLRGEExSQlseBf9EHqNOqmZ4wsb3hA3w
4xCzguUOYtf/TjE2ohx/lv02gqNsoi6cBe5+a9gaNvDgqG4g7Pxr6XXUXA60
l9hiXHSTKKjB1ve0OE1aOGEycEszwXpKStbyQbXkFzEQ9Ag+FPkDoeZpUHcX
UBdYeOirjqqBeX6aIXjqSlS3BKWWUSioH7N2KlGJfg7uG3TOCKpn4mU+vus7
CnF7sQ5zrEdiY8yyTho+8owacEq5hHr8Czb1LIgU2uj5UCnuYQ0xcr/2GUie
bGmBCqdfv5DfKOZHLKOSEaGu07rknp4IYz3l6m5vPv0Fs+4gdm5Yy1k0XGjp
o0NRwS5Vc2Eoz2WVZ5GWxVnAJ/vwNnrAa7N/Npy6LY2Z79o73+v6EN13Ji6x
mp7j3hS2LidCXeFpaGtrF6TlgX5EVvKZYh7gV4J0BQ47Watuosrr4jTbuMWF
lTAPBI9z0B59KPNXu5Wwua/3JCbdB1Y+eZgJf3nS5Ctw0Cmek/JiS5goxBhY
kO/9vDDahym5BUDhHETeNxOOqLxU31fPmNuOaiNLALMv03dWN4oH+MspwvQZ
rh8QWGh+WWuXv9zmRcc/YGtdLpk6uwoWdzdyzCwj65uy0aX7JIcjrb2GMPpA
uKaBnfp60DxoaMAD0/1r4LEI+dQmx+woChJcUjaOMoCR61yPEFrtku5k+KSw
bF4FQP5YppqYwbPcUnMTmGMGHnvlYttBmHsIBcnkpk4neGkFJrK7ygt2LksS
3UBVpDOy6OxI1dvT7DfFbzkrZ0JfQv2ay1EczYBs/clRGjeHtWzcQu9SgcdN
TnP+LwZQ5wQT2mNdWE+nRY3jqwm7qdQr85H650vtL1JkC6DKrPslSaWlhE65
AvJPWHgRIyZslmjSXVWhx+1cqE/sglJEbIu03az8Szs6sMKwRjKEAKiCNGmK
A8x3vrvhuguiX23z16peP6h/aN6uKJil0uqqjnVzcD9pgafNoTvA2FUa3kQu
RvFqTlxSCEBG/JSg3MiMn/+odFl93gshw2irBCUiR/GNQyHZrCG/AkNZ0pn0
sTVjqd85UhJw9h3FOmFYN36xTIGFdNEw3Cqf0xmhIht0SET6ov/IOid5aeQt
WxfYV+v1fkOJJl431YuqyXq3psSPREkI6Mh/lrGq/BAKQBMXMG52N6GdKfvG
bqH1ds4MlyoL+cU8xFG59q9tB5pN2L+kgtfuOQXeeTNWVFGNpU4Isnc61wm2
Ifa9RGRUDCMzODsFJTbLmQ2ymmxIk4kGCR6mAsGvv5DWGClwwnBtPEYuN6kj
DCSpxh3ZliyaFg6JAFiqcz78lsjnAR6bKbrHmtMayez+jaca2LyiDrqDFsLb
RLr4n4xAgapEshzSG6EYGDn0FZ4c4E1kcP/5oVgkrTKJZT6hwd8ivItQNccq
Gh5ugg4O5b4/5NhXtFGjEuPpdtEN0E1WLx/n1B1MonL7tN1/Brtv3bGOeBC1
NDP+tQ0yIreOj7Kpru4h2erZ1ueou/G5T7DESeoqZ6wCTMBHfwF4YdI2RoAk
dL9o56R/ihLuegA9YpOXrBzx/9DJwwzWxUBHi9D9BT5jSpcn922wU67n4ePT
a2S7v8PMcqCbRN7IBfBeINF2rpdXDlGv2F4gmKOtCbRQA3UPMz0Xgg6Z8tWT
u1Q1BkYxdcqZKPfBlRdedves9Jmv5D1DGQ227Dsfza2vd+jbabNbClcg5RqA
c/QLMOt86IMt7gYg3T01O2Y8au/+rZZhCSVYXumOrbjjGt14NdPD7FKmemeR
aOcabPbrbsGc+CLwWnfAWWxiE9OhbsDT5Y3wAjhdfVqqDgwXw14MkoYGxpId
ptwrfe0IcnUaq/WZXrfsBUvb950AG3KgjIULZK9wNjb3fqiehi+FGwbmW6he
igTFAurCf1T8Ddals44FmOrd5nb0J2OsdGwKP2B/i636POxq2KyC8bjIhvZG
iSzdJ+mzr9pyXlmuZ/w2/HkagMpZDzRHmPX7rg9A3SvoiP3XtjxhFMCBTicm
h74C/QiXSKZcGjXzzDWjY21Ce5q0D46sWmjmz2Qze1sC2Z6hBlx1KjdN9BzV
LK4bAOP9o2njhT2/rblIRr95B/1HeOTXoPfVI+ledXdltHyfdgwpXXNySqfJ
siQDVlIdYFD5Sygd5E490GLd5hShkC7MeaWnqA35qrudbpIMaHpl3TIvgUGX
vPCtObhfOkTgZQ6L8cKGDuQEimLUpxgsvuVWG+0U11Kk9luM1w134QecKZKB
hqo88JvqQBOewpsxYxwdu28w7TQabMtrLnnpLThVFrYcalnzC8LPJ2Up72zt
QVm9BW4L2ioZryptzaDN4q+MyN+ylHNiJAGJUteArLg8tmHBPGuScLwFVRKV
Dc85kHfoPcVzEeaADMxLAfeFPd227V1cN6ojrgxm6DFX8Ig0CzBB+ChNv1jV
vwutFzu34rYk5puyB/hWm2VN0c3dqI1upF2JTdXczH6YzGyS08gPo91txUxE
vHS03/aB9Ur0cjj2pA1SDQrbyF56tPHUMSF7OPDWjsr1auv7rTkqytsth5C5
TDSKlBEDenUCfpwXQb4jtAZKrAYgunbYiVaBC7TQZmUKP4//JfGDthaTs5MW
4pIdeY0LVYA5KiUY4FCMt9OqI2FG0ETzbYCLo6rUuGEFk1e73Qh0vh7a9/Nl
7fBtzYgzWyMIthBBeeGT9+HYU5bgrY040rL4anHbaSM2gGzG1RzsRR2v6vsU
71GyUvlPTtRkxOuaufcDS5SvjAanLp/TqFOCNbmQYvQWVuepCZKgGOXF8iCo
FyXj98TdGfv78owGHBfQFxJxSYaZCycdhhI/3ITL1cVMO7H/rzY+UMR5wEZp
LneyMsxsHP1vQacOwg1tczmXmQRI8XQcVuNLEfEAvtbT+ZhfO5HY4FG7bq5q
StY6KJxNJsQHP4j9avNmAHSa7OSnEHwsYutgqA4Yo/H4EEdqLbAl4bcM4O6o
PQn8ddAcQ4Djm2jZISyHPSWsNi3P51WpgX0IaLWGXUqQHUz+nyyRLIRda7ma
+Eq/QkhTRcdylQOuZwTmhqk0QuH2ettkGPPeSei5JyosHJAgyc+GiO6f9yxR
KjMRC5oIAngWc6zRaQoETeUuF64+TxmSC98MgVh6Y4I9zYe7c0Gr2jptU9Hg
JyzY0RMvtyM4oYO1/pzIQHiSYhPprbOWxOlcOZkxP0Rw5Ql9LBz762jNBcRn
EegbmK6UWJpvH3SfntH5WIr1hZKMwhPcbmjuMY7rJiQNuBt+kQFQshnKcLi5
QM+jVWIvfATq84iRPInhwzncJZcuRdLZGXZfd9DB6YjOmxfZmAzL0nHm7+j2
rm/KfpiXjo6WahjSBoKGcLv8eGnXPG6yC2/64HrxHt/GPABKT7IrCW8dO4Q3
rlyOcpdpJRBU4faerIFn59qS4wwuUppAOoaCwqGZ/wbsaqh658tUfFanSleE
+daf4CYPdplBJcsTKs2v/CTK1mAyMhy0i/36xZG8dG9EI3uFvUbY3D/WYKqm
1KlM77fQ0ItMFEbNFyJ2i2RtFnb7WZzpBifri9jMqIf8ldrS/R/zsvEUD314
YlV0DzV22wSgHgzr3temd0bCfT0XH/sPedUJofx1K3SsJWB0hZmFZfzoHric
Ah0ldLJw97qHhVg4eZB+5OdyAO6HvO18PPqvdVAPxuOJc+x1M2pYDAUAG/IU
LnrbIx0+a6txLRBEpD3DGGHowgZGvvwek4UmQOL37fvOwkdjJHfMouB7K0lw
MYqG5tf22SXYd3gmmMLeR2UWwfr1Ib31bOFm0ZRVZeCMbikT1cV55CUchwGw
tKfVtqWiluZF6Sxtjg9gnJ80lZ6P4torlrj+lWK0O/yFfBvWR88NzkFPhZBr
XqUUp9orVLzMQuIbWhQfnCQlwkJEUotEpqmATKI+wM3Gj6/OsjmG+Lx7iFeK
O5J9v8eZnibYWbQ73vSIuw9uW9QpkAi2yaUCPPLkgZdWhmHw+aHVCeMb9W9S
t1ox9gqCf28PLu4nDxn8RdptINitRaU8OgIU/Xk2Kb53ParczJfcCLv63gbm
QkgQxQja7hSr3m+nYlbsbCju0olUutEwTMCFuRYc8UrSjotWAztqQ5VcYLBo
5N5hCHkPzSkSbyC8B/ukMjqnFxup1qdqX8T+TrcBgW29rwTkbP8qhnhOdN/A
h381OgTm0k/psaIltdZqHMXfRwHWne5GLJeKxrnfi1kJ5vRVdtImETQ+8ZF5
5+1gafb/YfGENGpRxCfwxQ++GTITqXNILdI+a1t5yyH7AcYUBMd2Im/MiH/F
bWUxA8u8+8qIgqD42DqmlSwjdATX0czdUyp1/7hoEgfrQvUR+Fk2QSOm8TP3
tK52UXTvFCwUMQV0N82Hc6L/yGPgjD0y0oOjq0UfwGQdhh1gCVQvIB5jmVTM
9MijElWAC/e87jtgPnzPt4NisfhaOkNQ7DsiwvEDcaezv9nq3PP/MfSFdP4L
tOjHNwESlwnVKg/JfOoVLI2eg6dXaXoVR3zhbfN0H9TupqCQDBxHjIJbpJ45
LhLSlqYg6TaXLv/AxaW7Zp53bziRV0TdQOFV/c4mUnOtchRskBiR7yYMtkjL
dsgkx8gah6pNfpsVLw+gGfbUZ06xJthuCHVP1f2ONnzanXbB2BCrPlUwm5H3
RohVv4zAuDOIcOBn4uykRSv7gOXGGz8hHp1OQmTKcLKz9t8IIpUwCn7OrS1E
tZAKF+oKox57uJsx4IatDXt3tbnj5e/woaOG24BolluViUmu9uPqxR0VrvQj
EbQfiRDP/nIPOPapkIya/H7WmwbEQ3WPvOI039gVyOixNdyOz8/ZODQkde1S
ArGdS2QveOmnG5PEmBSrqjRSQ3h+QIVo/O14auJcIMhaupbkXwZItOYxXCz5
quGM3/RFFeK3pOuA0woZKrH3erX7u2GpVcoR+yNGCuflgMtxRLy38MklZSE2
JO6mNDTaMEWIlYLEbVE2NkOckIsjyPCCYNDbjmmYslXpLVarPHRFFiwsWELD
gprKketOCYe6Odypgcr0V1DVLXQBx+pUQs9FWOQS94vTqpMR9uhTNBPK0wiw
F/R1i/KIzoJHYACnvUaFIDdPPhqJczB1JzwSFVwAxCMU/YzIs5HmOkYoy5m6
7LV/Q3qGpc/8kDMWamsBeT/2mkE5XGbx4QeeqDJaLY3o4dkD2y6XwFUM7OHY
niCmC5X5wBpjwbBDaYF+gQwvKm3kuOXL7VyxzSGmicU/sLEW2ayOvqqgnWAD
8RvhIBy04cwlXFcAD3ImqyC8Ws0IeNqQ/s1BOQyjeugqUwyJW8Z0MMBnZleB
HK8aEHKobsoUhrO6rhWIJuDxX0ZMqvLwElxjwMH/uTmth/+SNkqTdUbTVU4O
ORC5HHMuCjPzat+JawDTvhnNTo2OVARqmNs+lGTzyNGX5Q3IQ4D6Mj0rnDBw
tJ3aP0LjqJp3o6vOYk513i9ENNHtQAbTnWycUCJh4zVSCkxfPd6G8LioTAE+
8fq4+53uQjGtaKl7MSK+fG5Ho+aD499D613bddObEIiuRJ19LhMYnNmKDRFC
BhXEeKJharpXvqaTQyygi6lqSS79U8eIoybNSOOX0Zrd5mRotMqvipQHUzxI
UEfLFbXLB4RVAcOiakfo5q1HyAMgr6gkOwBcfWh6FKNd4jrc8St6BEbZ2dld
RNql8vn+SK9NE81ZKDeZghLwukt+NsmPwQNbiNpMC4Oja2rcBOUAeebCxoHv
XXOd1EODzOCbCpC5bW5pg7w9nK609BYzDmsXTW08ezKkzRWJaAXUr+8Znnn+
FPnyx5SER9Hhk9oR6C6COSmbaavGbqWFXYe0+bPe19bWU3R06ZQUFz9n0uGc
/tg0W/GF5J/fgeYPITTA8tjo51BRRT5CSyJZc+7oLa+8X0o2+UxbUZ2XGAAV
ngVfqBLIE5DTh8+YJEhAaaY3+HN6TSpoZ73abZYo6ODLH5SCO2TPuRwSp/4z
LsJVY5SeWXoEBjdIBGjDuFdJMjIgV9qWZTgXM5VTHbbLA6N96eEO4P0MsdFh
oN7A9EUCFKqIovVfDjjT9g3B7h5TmZTae0uUN8FDb4GbnGXFQGnjLbmymOmp
qPKXmRuz50F2loG2g7DrvSofA8pxMyy1jEwc73IDcSds0hwjmwpdYzaXI7Wy
Eiw9MV67I9zjb4feUPB652GgAlekn07Zz9r+54SwddgEKY2oHF1cG1E0TWX6
pUUKXuGXGnr60UzWJxTLxT6F6VjPIrIHdSlv98gNMlY+XHLg2ClcR5HT8M5o
zf9WTarnDEohSV64e1/4RVHG8jLQf0HYHJrhezUVjIs6gOVS46yWYcGVuQFP
QXng4YkM/S6HN4ALyDvljyGaCzeaonhWNweDsWO+a7JseMIEwCRZjMjF71I9
7CPU+d3WGV0n5W+o81wmDBNOo1+wmbq2LuGfrB5QQKJSNLQQ1KnkbAvWhpE5
aew8l6H96qwIZbmSmn3HkP5GKyzPjEIMkleDKDuYPifh90taD4A70u/csqgH
vUr+DawMavmWrQ5BYQpwdWmek4/utBReYzPfkbFQAWLa5zLksODsmTOiNL+L
TBwik7Nk/Lf5raUB/CVTU2V0InTc6vI3jUdhtQnfgJTiwHpriy2Zpveh8uR9
Pbp2YUJVJ5gnlJ45MMFXPA7WdBNTgbr96TAv4c++fW90pLlMwl5oc8nIc588
t1NrRY/ORBh5heWW2WuSK2VxfoyU8TfD2+KaAOgkq6hiiIU3P4G8aqciBFyJ
Z1fLxpRqvhVFXOJRMW5+1bukMyycOBqz/DpfUGybTE5HublJpwXn2cZNyWRA
qC9MiXc6+RBN/W8hovXAGjiDEQ8+AxYh/UwoKYpYIrW1YMuO1yWbrN0by46c
b3HdMRlkLpfhC5uhwEaQHyWm8jMt2G0VgCChjLIdb5bZDkq7Fjnc5MCLKMVM
mFqC48I3c3ntotiXni2mOM/7Q5qY4aN9+hBoqIYsTE8x4Khz5Eo73eFZhmmg
PF9/Py0+J63PYmXUp6re/1hzekzMr9M7JgUJ4uL6HHQVN8sj6LQq9MwqHvbL
DR8nKI00zTGGo5Au5dhbcAozNSSKH8v5HGh/veeaVH5vVluKOLyfFZDvUNdZ
0JwroGAnE3m0YLhVJWfYFOeJ8vT4djD0J9WdFMK/MO7TD55Zm7ozgpMuNHrj
ZvAJ36ZtBZia6XTi49ZnHuZXPr40DPnSLZFnAze0tHCLkZ0LRxPV8DXg/pRh
em4MH0ey2j6ZlXOOBjZm+Zf9O+2njyOcGiOWx/dJt75FI1qfFN5zGKFKrVuZ
gteW7/2w09U9NedoJxBMDMLFlz9ie4unxzEMAE/RCsAwtwT/C8hD9MENUjc6
YlNx0LQD802AP+SBdvqeoduI//CZukvxLyld+v1/DjBaC8fdqWUIElEbgnWq
r+g/MlOa4tFoXyzI64iEctxvB7R5vFamEltaNX1jL+8KPWqkzer1fbSnhsAO
NBFvbjHtPF1gQJJKApjr+3Vt/sl26zE034U5EhFm66E9Bl5ijSfkZbNW3AyL
8Tac+hh5flvHY0UWgDTTOcquYDGf4/fw/ehAXWMKZUVPOfgvxOtLTb1eFJMr
Mooomc5/FVcFrtohglPyzGi1YHb5Q0ZQPz6IEuUTOBsTpNShu742TZc4kIpO
MvPtQU0ruLDWQxn9nuLHg2QwJz5vLuk9RfgSAqSX7QM92ZEJzojO1Ey0RTAt
bxblaWZUHxTTDN2cq5QbTUMRkv452Qj42C9NTpiPC4xQH2adVDCQFI2mp3QS
bZv+XAhQJRuaD3+FCJADIAhJiH3yDxMOpFyGUD4J0aV47Ec6LkWhwfptPbjc
FOeedOTj50qpnMcUy//iekhKzr41CyKa/UnYTrBTuPdYqbnijiGNMqBRi1JN
CiZy24vGAMt954DfBbb+nb/M3+GB/kEzqbZrN2Ubh6gFAm/oTevUt02Q4OAo
cHau+sNL3RhiiZjxPXgsWwcYyWAQApaOnBZpcR/rFuFLi3XmWzSZhSHhFwTS
rJoNjTEccWbHarC05yuw9p/GCZdnRSrrav8wXRnqcBgCVi5BP05f5CAEzcYy
a7ogGuO+0yjbsOdwdkyFbkFMwhteNS3z5GCW8ozu3ggBGF1DlC0CjEg4IgMp
LPwE1zYEMIdWFYhP3To74vfiVF48K1QQd5FjI2SNeVt6KmOZtjyOGeIk6Ehs
s4ul0z/qMJebXIjkf7O+jVXyGubck2oTqiJP3IMs8rKY1BRJsZksfupAPyEt
YJh2NtQQebmOJ2XFvSHutt4cAtyb9Xo37CrY/uk0wW2LEYNe19b4Lhlu3WZA
NSh7kuU8Kwrov3yqBi5thnLXKoz+gxDIbWUlkYFWgUA8yzErEHyTRes8HMWF
N5yZlLZVQYmCRpXO9c7bX4EMiXw2gJl++q9Ug77ub0PvhiHU42dUd9o/OeJa
FUFNXQ3W8JOOTn1bd52cXz0qykUlttv5Cvc/Q9NUYWxFlR6y43vEPcmhgeFM
PCLBE/MCE5XdrAYRIaHAcLW0C+n8sC8IAaDgEmqvlN0EjV289CAQfYdg8vFx
GqPYd29wTTfZHdjzT5PvgZQhsnWmfNurgOY/73E7YYoSyrpzN/ZXAOr/WT0/
stZZSFwWSOabC4QiRW1AJQNlat1j7Xw5gAXr+wCYRSzg1w4HmThDP2vbKMs6
j8ebOHoaL2UUILkvzs19C26qt+59sO7wTicQoWsMLU5pCJ6sTUcSrBYwxOUH
FnlLhvfnrGJaT2sCxaB3Vn2rQCu99mVzWPtKimq/mOAC+py1UHcWlqehPeom
nEQOez8pd/dbQXDswEr1z+ayu76chuq4l24JMHHeG2AiRDH1ezKZTNIHE3A2
j/uPCXjMuzR+0WdKwUkmCKZ2ebq5n76/Bc5R1D5iFwOEim3Oomvv2FlWHDAQ
yUBfSIziQ1nrw5Wv6QvDGb5MWFeUwC8kIDOdJHHPKfAL0B82iaOWptS+a1G4
oy9Vv6FDidVtzZPaOEl0oEFrl0wMStzSP6DZHVQvbj8+9jDWwIoT1JgkhnQX
EPGTYpFoluTSbwvTw3FHpWTpUGNB7rmD98x8NJIxA3tEhpx8SZ67XNhSDj5m
qvfMQVMMMRECS6Ah8lfSNEJXz5g0oYNwWA4Iff2+lIQs6+cUFohk4XB5XSiz
jSHulaWP3uevqurouDqctSCGQ1E6YG8MeUO8hoIL/kxEUUTHtP9Akp8o1DDG
7vO5uqpnlBhDagrqdjKjC7DNY11BAetcgCI94AGtSySjQE78j4/Vt0SIO27V
+r0Zi/uXYFwF5Gr/qb0KgIJIXCO59qIR2BixNQJgLNuIpVFuj3VAQWbmjh3H
o+Z5lMUOQQsn+vUBzFeyfriIiB+GYFzrv7iOuRy4LRuXD+9veD7S+Axuir0n
8nF7rKksrxErxwI6EPw1a2C6yjorIHIImpBmu64goUA0hgKU0/VtfCqeUa69
hxwtSc+j8ZP5x+D0Yo62jaYA6n/GQEPJBHRKeufQ7CgbfR2aNuq4CyP2/LFW
bPb14axQLcBJeuToH/JgEFA0M1ps89GVoYeCgkldfle/453KqFwjiChVDhRA
VsnEQmkLjGppDXHYc0h5iP+AemWCOCrbJLjThwNlmqlbhgXkpqrCvREdQi7w
tWijH5DB0w/xZ015fbXcvoqRhGvmoPwZKqRsxNQB8hGlMp5FKCvt5Openzoa
q6+Y6fPFq2DQLbUJSegJxqK80VCnUiPFO37WJuW11vDd6r5Fuf+UTl2dLJoY
FE/0mi2Rri0pCAWp+DakHOVM9Q87kSvv3+5xf4DdgDB+BF/AVbYB3zAnZdJi
6saoCqNI3yl4u+AbYi8HoS3iZdZRS2lbUb50LkPtAo5Jf8jgLRvAcFN3cGx+
XjBHpBre2iyini6+gBKpi+//VKwWjUyVJ1mh7qvMtdMe9M+I447Im2OI+hm4
1FtPVcqff/e82Q2Rk6C8XL/JKBCp/16rJmV/rbsgR4gfOQDqrsX+IxuNTBkb
AJUQXUzJPs6TupyPYbOvym81cFyfI04AARaZ/H0W5B0BA10stJm1RELuNyrc
TxBKhn65/6SXoXqWIpqWAE/yoKuPetHdDxJHGtVGTALIgoj70h9JyJsODgSQ
ZZ5GlXnnvN+bOvaYzLwicXxldhBUVWvDcSW2di2BAtPeFa9RITlYYngST6Z0
1YaM+6G/tVsuu/LtRvI2WiaX8ClfzZWSbHZPdds0WMK7hkahh9GGEC0+rNGk
rBxnayMIHmDqebVYZyX8vQGs5uC0Pe8zmwOb1ABN3smvwjkZAnLTZdZYJQkr
ngW3kqRN3YFc4tv/OjcHTiOG6xHSbRckvyOWXYaIZs4jQcWJNvUnVoaVOOaW
qQhKan726jN1oDvH8KhwxIMYMfRmua28ZEBGePQ3u9N8hN2j0Np/hCA2F4Zh
NUrN2iV6KpsnzAcWFo/55Au9qaXhLvK3tQveBYisnRMTe0v2K6k85gb6PEdL
dYvya5oL9K8+9jiDTgEVuGx980XlX2ltUaZ/m1W8knCJmpJHW5ouAZTJ3LzR
VWLT1CLu1/tK57ARFPRevJ5OgyCWipsdsaQBvoXCawoufC7eKmdbee2jXANg
iFvKtE5Wh//WGia9TjqpsoCWEy7ZsYxWjZzYgsBSQIPGv7AHvxSbQwLbRooh
0w/1OAjOYKNgGKh9g+HH+bkxxxyFzHBkCV17Df6tn/5WhAwY1ANBCXdL4wxh
DVdb366G8lJU1edXxtvPkm04RaWjOoH1NgE3IkBuoEF3DZzY0SrRNS5MvVin
OALJBM5cVehO8hIVlCpyz7wyctCP+H90OuXRotzsGc46fKbhchutGQfb1ZC5
psHuiJ8A07qt4IaDd6aVWcZ26oCNUrqVdS7is47zHv7K8XzwxZci4q+dIs9O
Bwa7PPdPaneX8DLsORMwzPq/Ig7SzjrjCWdUUX7CGEGuz6p9lbW5cV7tJVWo
t/DvlsU9sgJ9nUzOH2gqv1UKMjnYjJWQvPf14dIkidIi6sKbaQIfA7wDSdGC
xLlc2FI3EfMo3+XWPnG0xIJf7LWlFvUePj85tB4HYcy4RoTvkE/H74Pg4TB2
lmO1APy3+miK2PVE5pojEr6Fj38MTtxtSsiiX+kdrMBUq43B3v7iHSe0gjyg
9CCEGIMmTYUYgKwDbGBMtgW8nfIA9ugcWeCHkk46LJkq1F4X3KehkHSHemZA
tsBi8yTayj5GlrfCuc84A7Ls935khGPEPwSYvzwQW0JbDTTD5b5rtJjOSE/w
K+GYBhpQjYdsyZxmbef/MhMJ1i247ZLLZYlUPgffzq/mjPLw+5RLQzqGVF5g
vLJ3zFV62OVHim9cKXQxJk/Trs5JR+FQYwQ2PoHGw/5wlB0flZS9RSNBwKdk
Qu+yDeNUnbwKn/xqvhxruDrUrdvqhdx9Hvf/yfwCRqUol7xKrpA7qK9mBAy2
Bn1rm/cRfRNkCP+bVfkjXyBRZXm+Y7nTIX4vfWRZT15es30C9y8lXrWt1Xz7
Y5r50jog4FPpzChqNqEBXWyHBIPxfZqr6QeT1qwurBqzkNHxR2Fu/eI6nLaJ
BvPQf4+VTesR2adj0Zqs8JvCsIfzlIOoYbQPNjj9cKnWyFNRt/s9bnlJHnjA
wK8WMl95YRJTKPs0pmE0Edw/iaDY3E8jyRU/2zmIlGQzgTQhJHpd84Btgdoz
ZKCP/9TQfb8VDCy/fgILCBMMmT7R3e40Ty69WrGxOnHbFQrNYB2awcvSY2RB
X7YoWlJX2fK47/nPZf+0JruL7rzhXgw9bdkSjkAKHdZcgoiefv/wnDZS/7c/
ySgdghdwb7Hnu6yTVNDYSZbJbYizm+/0AddZel4c6NLiKjqYfvNfpNEueLAb
+vwml1rrrWx/QUWIWEooME2yky5gO+QHxqh5zVSsn5p7R0stqHCoExkjR7CX
PVgQgX0KppWZVxvKRNX5bsjljPc9us0dCnFezyDkz6vHkQnu9jPE9/zhdi9e
KJ++ToOzu0kBwh0lkyQ/FvfwfBUGyvkkmX46Y+IsMmk6oSbYSAWv3Lgh+jrr
ON4k2TJiIrF9DyD9xWmB4cduH5yW57uo3RBqCl2N8xbzRP0ywnITcKUkgtzb
9xqUY7+FD0f2013Ow39jMdbRvqbIBvYHSNib/yy7Phmp8j4Ena8x3/gnKq07
TMEXgRk4gtMAPx+tE662V76Nnoe0i/XyejbozS+GFgRNy1vtgbeM8MN6gZ6j
r95ixaqUYywBpCbvXqbthruKIpdZj8V8gVdFZTGwkSWUnMeHh4/p8zohf/Xw
7NGtLcqW2uaRmqIsh9TXAyKb9SuuUke34JCzykAbS8brY+68wG4fp9Qh2v1M
w7Hoz9tpcn/D2SFz1F+nuwighkPxpQU28XyDdDjQci38NA1d8JZX7/pyClP0
mfnFGSaL71BLSXEML7KrlCTaVyrYv3gy7fW9tEFTBqhsyOY3nS8/vjcLQTgU
Qz+IVBMqJlqjxRAhIVRSxOq859NLBQ6aexXM1mzgoEsqHkmTlcDN27z9Zptg
qkltAWPr9v8LLzxAAs6cwYY+9Rbq6qYyeteYHWbYz0P15qJeEG1Uqe/c4rdS
Iuu4y0+86d6TNT+XXyfQKVVMpN7LaNV6OaQNwXMgG85eZ6ur7trcEPynmx+d
es8t643lHapNzIh6M+zjAjhDBwVDNUMr7gfZPUBCXrV6s7G1EjbN96MlZmyi
My8jdiq414yIwL87NkB4s7ODrIQFlckqIH6AR/1Ztxd0crzfyMK4pBdyvYXB
1KIfnxryt7zrYxhIp/piu8Eq/eEX/8ojBWJwQdlOSq3R48rSie5disy+a8Zb
Tjial2Apbhd2KFH6azFVGw8enRo/K0z/6UNKVxj3oJ9YEkIIMQNeaaUIWEhL
ewuHaMOWWhhciVJ30A+ILgVeHA+UPSxvqXUPtMq6CBWDU07d7P4Mrm7YS9M3
Y2S0eY0U8qlnWK7W5jv1pq43hHAyrN4XKn8/jIxKy5Z1zioOUAOPovx1tAZY
y8uzLzHOU0dQnPssJZXTSx3PD/Ck6fJqXsRrDl3bMmNPPk3/my/bKDdEimo0
daFkWTHC/qTiZGgu2KIKvbUqnGOogUsV01UuPAd2r1RVPAneRUxes/vNIv1T
ylQDbsO7GD2PeqDwEu5EbEUpiNDZB469EQzM18wrABgShDcLOFqxyLsy7fdl
nRcSg1p63CLgGrHN7GPT9ogLudx9a/SS094a2AWHjadxhpn6ssg8R6gNeWhd
mPD3pfaxSLwQPDKbXu6FbOcXHksqkkMCHAu+gipb9Y7XSPGgnQ/hxhrtj/6T
Xv4909tq2IzkQhlAIj+Ik5VYIvmb/vZnzZE7b538u/lTo4oGt4srDixhhsTj
XPJprWVDqRLQhNsMJ5zc6RSqZDXl6tA1y4R89chpwiJv2NXuWc+kdPgzNuRf
c7r35eEnpGoPYzDgQEnaFAVDdg4jVMy4Dt/daTP6GablYYA/Vmr64Xwmg3t6
9ev5MtacmDTSjhEjbcbedfdIqi/3AvcVxTh8Q7oRYbUsXvgqw2k0MlpAXQhf
/x43FD2GnAFPYuV59xKUravix5cAA8hPKGFqOIwCq11dpfFRJFsogbWNPQsr
CmJogc7a9a2K7keD4mvGc1CmtLazqK18CwFwkFCDC98QsgZvDpqIQipgFsR6
OkW+S8SumrLJTUJSjgsMdsz9YjeWBOYye4Q7+qTQG9Yj4UPrTBMx6hGWJcC7
O76t9ydshJHGQDqzADU9CbjtfqpaSFG8xTJv5aPeH6ucQgXGIFH6YGWduywT
UEnIQ2lnd8+tYdON0s7+4tukJt5DKHiBqpiFvAEiMSv0g3xLt3T8oNd+PrU9
8om0UbWICizOfqtpp5QeF8Two/Dl0Pc5VDNvwMZTVyef/RyoNmloOZmv+vVZ
wUg8JIi0G9JKKephc6jvqnH+PerDJ3m+8m4xQRix/fVcsJfZBP5E24spf6Ve
f//gD3ne/Kv5dmouYpZRF9eF85bIOrdcbiJpllpo7XzreqRP1kFwIlBWRMcS
0nId+7u4mbDnOSQiVX5XRc8RjIxz+F564wINZ7RQczgnw+S74XBiLcIaFVbG
ehU0+II85cv9u9KN4KE/cdCx9caXe4GaVeDW3NE2t3B+/1nY35PZj5GNmMfk
Wu5T2ixbBAAHt/NHZE4aq2fSMWCf0fXpaYRb3J07FGnXycca/CsE6QiEDhxv
9oqv1CD65YmUmeLOyg4pw5aArXBldMxRJs/6KVEzxkMlhA3zJgg8LiF/mT74
amCspAn+ktJNN1vV3ofOKZEUhQohGUWDhKFHxZkiPPNGKvPQp5fy3UbK7QS9
fr9lBrPXTJqXE2EAc4PkXzGlBTKVzGJ8iQNsA6wp3hDY4gx44z0pdETNDijo
1mh9U5SdU4TBh+53IAWCwYq/I/wndBIBHElhqgjEm4BsWVXaYcz5UOgUV8Az
YiEGfzkDJI4cOZvyDNu9SxWNxDoOs8o/E37UbyZq0JWWZoIXenr9tCHw6OoY
PD4nUE53BMa35ZN9g/uYOmzvEVJfx9Qc6fH7vD3YACJ18AKNQSAqD+JHRcMk
y92kmT8eHuehJcI2XWa5U2joTLgoDybjxaQj3nlxl6YDJbdQ7P99ug5sWZ9g
SzEp4JwlfLLEiKbXNzqczVp9eJd+e1/VgWVH0oRc8udnaddtPMFVlj2kUVFv
op1oIyzf0rQHfIEVTm9HH9339KCxddHom69EnxfuqPepFqw8QZUWwhKR+5qM
IWiYaBZwEVwEYDO4QPmDWo5Ki6XuDtrkHAVO3EMVcGe/QcA8eF8atQQCECP0
g5Rk1eIODhZucHxkMdxyH/fT5FQWfXCAvW4M0WsnihDgi4ETwkvXsM0S3/sS
6Fu532PL5gvIT5LRhlG7opkRkiGvRSoi22exLA1UHauxno0JxEwWq+G/s9Hs
rqGuQZg7sYmd8fFF6OETmOjgVC44nqSrYK47N8j/lBpe6VEF0SsHtVQSvxg3
2MjFjfs/DLu3pOw1rfExZTh1x3ENQ/gkC8lx5b/pUWt2hhqexgCUTLA3Q9E0
Y8JWnTWVG7E99P6WAYsBSDiS5oB5O0fxRA6iP5HT6pkUHPbi+41U4B7utbj4
y5g0XW8+FXu3+KRpYQs+3tFNcDeT5YNtaI/qCVOigfvFomW8y6cgCUxAjz7L
qL/gbv1YRnijpYKfi7Osp/FoD9vRtOgHsOC1U+WByNuMPsm7gIqw/o+ZrKUN
CGthfIZB2PhUUlldkqpAQ2nfZqxk1hjQsg5w8h+aCIUglBWNv/0vdAONufXG
u+s6NOSnUH4WVapDni42Di96LxB8s8NxmvKrs+SS/rJo6ZmqyTfkK+zTcMXY
nMPe/xY5yfmm5QOJQ/QfwmPWNQeibiV73huqXId1eyI1XcTmDZzRasgn4rXM
0CgUVcbzVb1RiEuKgo7GaYjdXdXClwFW5oFLrmBJxbK4Sb7QGnztB1oWK7fw
M90mrylL3oJ7LknX2XXxa4DYZm7SCyJ3dLvZs9IiyqeksVHCNVfLbzUG0HaE
fS+t8JoZ7Uc4CVFeIGLnzXJNjiE6oDUuDrR4f526mjZ4cR0euZpY0oPO02zt
QrPSHJZoxB/XQ47tPjI8qxHahufdMK3jdXL/M+gp40VArLomXOUyF11eOn1W
PuhWISnuZB1iYsOztkTOhdqm6bHhNnKqEgqY1q8b08sk9nIto1MUgA/kdh5e
dFdOYsGqoVl3K9u0OQR1zq0l4+hmudqalZo/MO0Y1xHss0clJBQKFT2at17J
9fY0k1OhneYDcjeYgaUfBukLOk+B6qlG1kAeyB+CkTzwI79tlVKFcBBSmsHG
COBn45zj/+RTgF2VG9Pl+ojvPidQRc7wz5uo88drCN6e/CnolUV8O05RWfwc
7kYxEblKZHW7MCO9xix1BII9E2lDn2ZU1iv+BsgBAhzmZ/FVKlU+dcV7EBFm
vHMjKLUvSiNFy5dw3xV3C5G+nkjd2jRaNQYZjRkIhkO0FBO1c0zOATcvz1Z5
vm0BU7mTMp6rENsflYdiK9Sj4jSW3RDekKn0XSCNxB+6WFtv/30Nu7b2mqJy
gFJbT5gZ6wUx0BRDzAt3J1weTCzRSiDtVwge9XYn8QHViCj9h7xx5qoACDuv
BhwV4gPtoPnH4VEmC+XwSE0M2tyE7/kEjJENmj+NuzZ7Wq7XI06WIKW6/Mw9
F98vRIQ+nWp2+PMmuH73TvxGRMtt6vtMnsC1K/v8oaLEnjrmlBVLt7cuRd9u
XcacTPDqW0VHTLZBBPQddpZwLxp61tG68kjVbb0Jx5X/XmKdF/YdGjJxfU1A
+1rrLakbAO4oo7dS56AuEIVC1E66jB1sIQFqqcq4AClUKxejLsJzfu6UaIFr
wcVXYWRkxEsyKljWcITe+K1tFlp/TScLMf32FuM3o9yCJ3Ikjv4AnVX22cM8
pF2RCDR5ZDVUNUoSb/AyjAIdEOTZ9yvLYgsrqXE6VveXhp8D/O0riiFK9oSP
k/aRljukFyRGJhfqkYz24+MmVyuu5B6HR2583TjwIWUYSNNfV2bfz/JO+kcG
bN6uZHqGcnQXvVZYnJfcT8p29p1aDD/y9L9mIU8FQVEuK9EYdrVMJjw2IaTL
hnDooZ/dW6wIQDQBsYxjkAEkpC1yMLGrGeJ+bjIZt2BP1miQTGGegHmFb3sb
reY8YqfV+Xuh45TIrtqFzleQZi/jPbNvuUfVuRuIfdMq/pvVx6qTVQSC6PD9
9451cqPXP1Nn3jX7vLtfLD7qs/Qh7oGKc3ErsPlZ8Ld6r5sfpcEG1ZcG5pAy
2fxcVWtF7TZ9QmJdjOwy8xM+URGl0eZ8mUa/60lJFs28AK3RDHIoeJgZ4CdB
LVbsjfZz3Xemq3I6yWokIwpQFiHrvr5hYTshsBIHEZLnRbRwaRLKNvnwSGYs
YDtMNf074b0o7BIpeEkRFnQOvR6FNNkuM8cZ8u60Hqu3mLqgQEAkSlnwvBIM
g9XkPNluOoZyZDUoMQjpFXjhco70nzTmgcSBW+GqHjA2vqm1hT62IMHt1LzM
6+6T5I+WeM4D1p7EuKeXClkDhcfvmxOrpsv+fn75/CJlsA7Wr4ncN/igOoUp
gG/hliIkNM5+BGsGWhQL0+Qa8/53nBWJ/p51TfT9RxSUwhuAWrWhrLDczqw/
w54eM1mJypkojgKvQvCyjYSTHA2HfuDZ3UeFTcczBWMgbzj3D38+ym7X+EOL
0mhF+eFM2j0wmHy5mRUYl4LQCyRPbAVgtLXqMC+IpCToQhl1FRZSuxTlLTwx
morQLHyBmtPvz7GyexJOLtv9LlYkFLx8iWXc08rmGoK9MZEB+3TJqik7tkTF
+7w5HKGh4g1Ao6zympEYtSZ3P0S0Lj//v/gvdL4yoVPelhohGtPTAKrGVY1L
uVNXLsRjFRMB+hnSG1RGw66chQmGoQpjuIOyKwG+mwqYjfj0PIyNx7806dae
/OMqGmnGr1LpXOcjXix6hOggOveERHWXu1vOREKE0tDtEJlbEj0btZaf+/Df
jtjBLWzfZ8SkatVtwxyrKxsB/bRA7vulZN7blBWMB7ia7B/4t64aocrpmLGs
Fg8ZtR6zIquoyDSEG5NfdAxzJB/Xt38Gr4DINIosdVBCCaLtMZVhYwqoIEut
r7yC+TRFbK4HNaA7R5N8JySRUan6CUs35JkA6Cv4aO3rQAP6jYZqR/NXFKNo
5EKiGmxepLCW2Lkls8Wrd6rP6gwqLXvOlBeAPAtxbT5lgXUEAywkNecRwThC
2vf4qLd19+UOyfWsJ7PGMqCUxOpR/5XmDR8Hw/UEp+BAwvRfyH1ub3Hw/YAL
EoquKtI1MHsqLshJeKw1DL8KvBpfeuVLY2TFKx6xve8wr589Tk0Ks6QULtE3
sFDfEZomoRvuNdQX2X1ld3mFhNu+//0ug7TH5rRqbLasuoc88CYX144bDqjv
y+TJKfTqZvWT8hmRm0/dGaFHFYu0IhAEcbGyCBFMWUggNkqhPoyZ5+dNgTRF
sc30ykjFy8F9Fi40D41v6R57+ur8ONl+8TlQtwrcEF+x8NG34TxUruUDlf5H
sqAvpbWHEUYEdtvMvzUQd1+qz8xeWVDM2FYVSHfzMQ7/bfmXIGsFz+BMZGbo
PLCzpj089JdmvBVlShWxJiUiS7iNXdUX2rUmDBt2CHKbyazfur/TaWvVT4Bc
xRq9DBY9sSiVs2rynIuwAQB/tp6vgdQBwoOafyti79Y+tBtHDTaAWwyHTw9L
xo82ygUXZ8cAwJU1NVeJNEOtIvSdjgB4mqWDEqGhFerqSLJEV3Pbw/MLgc8B
CtEnUf2A8dT9J69fw6Y0ktXlnTMDZQHsgJIFILeq6fKaAdzpFVr4Jnrb1geI
yL6RTCYBlQhWhe2Vp/078/DLk4742kRzfvfFaqKpqEB8weMNVZWlgcEbNcmg
RruPkEAX2/rMGqdJHKGBhrJl2EzmWgpBgEJFAbPuFScXRrYszcs4xbruy7mD
hrPB7jE16nuCS2t1o9rYiUvl0kqRHmP+QNCkFWKXJVV2Gamz4q/3NGrgbvCG
8T0W6yYlNCOcxeMyN5MjcTNq6m6dXvUEjqCiayDOZME3TwID+Q/VTPSypOzl
SFYr+XYaoQs7VhoBye+hNlPkhH9Ob6fvjfBa1J7u5Dyt/sGWWQSOiJRfLyUF
qPEHZandy9fx1NvH2QDPAWssdL/yp9lfD7DXIaihcUZFtSS84SOoimkIThlZ
R7RgOI+XrKvoJhzIfYPHH7Ndc5JinyjMt7zCX0S1H0j+XTuxeKdTo8RFWZ3a
9MLsNJezHajrVhz0r2B8+O5Cm8nCqeUdxG91Q/1U4Bl5mxKc2C09qWxguzUO
BW0wqdK5kM7Iew2ItrozpTpV6VGxFeguSHFlD3uvtysNzLD9sE7fqNx80qbr
6zK3hdsZqTUSsYEJ1j8NRxdJ6nlVVKyD/AVrtu1kwF7DCp/X7n34e6glInEZ
C96GgqRcAUG1I3o1uKVunwcCWOgWz5ngWSh1503XdcyoSGvRzgZuJo1fydmH
rnZmQZQBms0/JQ/Ptht4ANYBDXU7sBMzM0I4NEdVgQnWAs5ozZk2ZBJoCn8Z
W2KYaC5RVRx1RmxoixbvZuYPn9lbe7q/JC4KkijSgiOg7F/qa2nmRRRGOOIa
imJWRFnuu2aYG4nP33r4ghfLHZK8FynU3gm8az43AbTBaXg20+tTCbejqtN9
kDuUuY2jAWw35OVevKWHXxtkn5N9Hd3vqdCGhUrrBveiHYL505M7nu+l21Xj
YSALmeQfi0z2VZvnqWBMT3VIfAb7e61OQiyBf1U/Lff/a1+J7jSodkHK5zau
v1G8iokwnUqdqAnIsaur08t24+7EegEwPM67D2SSGHx4H5jxnzEXY+gRVZrY
fzGvOOXF1F3oAoO1uF5zAw9+3Ch2U1p6GLD+70c75tEM33HT75MPG7K97VgO
U7djYA2+nA/g25hST8BHF+HlYLyyAvg23mkPSGCfj8k0vlOmyBlit9VRUggm
27FWalCH1FcU/CRmJ2avRGQ8Xdx3z8M+47envWldGHPjx/ZS9zN0H3xYcZEd
DueTyzizpNerMIyGv8qvrf2gqGT+Uj61bHoYrllO3Bp8vfwQCSn5s4K+c98x
Q2XMnVJiTuJ2bVtd2zuCNdr2qlFcEX/iqSN7quFYWbWRjeKhZL+LV0ZuHjP4
WPLeCQYUeeAll5zPs04HuKBLT/OqzG1oCNtOyiCgo0nYu+RzW3uwlTyO/79Z
2JKRTIx4i6ATLOKQxnnXopUcCR2DsA3rDIq16b0hKxd7Ju7StCaK6Nn+592I
SJQqJUwWHtQisdoxhTwWQLp/Q+CQoZfta5tjdENX+ilLw1W9mi2SxOShYh4j
RtprSOvVklxgXMJehOmdCUVUuMG6uU8BpHGdklGi4DCNiQXFGJbBmtRWKWPT
la/sLBzVmoUnOLr+EEg1cuRE+t0CHIBMPZUxZzaeUiX5A0vlrNfItMz2Phw4
LHu1SFiaK249ATj42x9KYbpwMi5q3gFOFFIcb0tmZS7P1cBjb/5PfoLlMwRo
k5tA/PZhAN09HwYONSN7bJTRby87wn4MDSWGDGCzP9MZIP+tuWHVy6yqWt8x
M67nO/INhfShZWUMThER7ECiZylVjZeMMs3ZmovVj83QAiey2RSMOwjwqKtB
Ealh4jivJnc3/3fWEdK3pmJi2loO3i+m1Uw/HL75z5BdOHrgAoG0Om/jdION
KZHcBks83KA7F0gtY8t01LAFNEfGvb9Wd4+Ae8BQYebewReqNttWSUU6MPLS
hn9AI5OFjTcoYvoQHI1m2h0xmYfK8Np3nE7h81GZSXFdVo+CXcxY2sSsA40Y
vjpeIqwoIgHfZIZ5jwhW+bY1QS1lFJH5ejP100pdWCcwwVVaTqtwD9+4HOKs
rcHlnfi3GXfBwFXuVIhgyhCyl2LSc4p7l6VSzW9rONYj0ZU5SQAAZ/rf497K
Z1Jfhj9sWTGvbBJbR9IyjmjqPOIWsp+iyf96zQV2x2GzffqHBEWtm/2MfE+h
arV2dfY4HecB5/4mgkLWoq02DZL8OdpLg+MUt589LXEYvg6o0jvBHA/qwULw
rRhz+Z6O0rHqh+7w3pYPvM8//N/uH0wpXjEl07rxNzLYHPoIf879vAKtbK7+
7Q6cjHO7bH07MwCxy5ILbRzkCpDVmWQVtejkO88OBTu5812X0nBDX/2kpZgs
VOjtBKDGs5iM1jsNiFx04SdAx06czKewq/01/ORVRZCyIHGO0NftHaKZ2nqw
t3wH+87t4xBfD8VOHoR14vS/r6puPquY4PXUP2EdYZ09T0/42QxQUAefQjZB
Mlo8WTcTX/+DWUwXtNqYB23oIVvqfSGCVzS7MeibQqVYarKtyMWYFE3FxRm6
B0uEAoE9aPwIPWr9c3hihQRkTGFb190T7bxwWC8d1maAQi2x7TQHDV7LuDyv
8dtTi55xkMsI9IxJUYQ+6+SwjYN2kr0rnYq/EMkqZtOGWFJHDAOT2BptJTns
sRUmjUx523gdIqZScUcoH/Cxx4yyWM4u8eq/nsZRMqKetmB3BcRFmKOio5e4
RbFaUDwE1jJSmqWJg8p1xHTBcsc4t5d6cp5ewyOxhArpbnhUKmUajdzL4ada
aqYMn9bI0Grwr6qoSbcc/ZZQqBpgCpzbuAywDkv8EcTElDsFrDVpeYjy2k7f
lR/fQvXH1WCtT6Yjh26lsxGSTvYsv/ePIeQ9sRcuLakTHY1nOjhmAM0xgqDP
W90PQTW/3oVamE9bXykDyP3hk4UYjajvr7B9CiEyyQojNrH0+QXN14YKpkNX
rdOgJUcVqNak+2evivrVPpdIG/L2Ac8pmO7lZnInCzdIfG10wnUEzvzCysla
mNBaHuGA7aDxpNzzjNULczcUYLnzEmsJNFwrPsueLwflQqSv8NO+yTKlWaO4
zKvnLUkt5DdfaCzecLpQkFmS1CszETnyYy+KKpHVjydgPsp6qZhLFlDcjiby
xcrwmRqh0B7VLMr0ZFS8/W+IOKYtMIaSIdJrK1/nh8LmpAUolYmwjzYMb1SD
4Um6iGeSid4a/87TQImEo3PgeqOmGq89+TbiESCXhXsU9m5p+rGp9txOYQyR
GSviuPvm3e/94d+CqESGNRJlNMlfT01jgAX7rFnOwcOWT60X+QeA2BNCGmTU
7jQ/wxN39d6FYAhXOc8qRF3+RIvXMQGNAkb7nbNMazQDHmEjNYX7anf5vbCl
YRw6cKYonVAA9ZSE868qEFfqMJoky63RfFNOWtwoVo/+1tZTMcDRf4nQI4Ya
NESiKRvvGSAMdsu6O7J5RFwhOXdYsEZPTBphGWzW6WiF8s9kR4Ze2CSdWa0S
8HGh6SnXoiAKEUdAOFmCMNBDGQbG9yny/cZGDeu3y/o8wXvy4sMxaX7uYZ6P
WtQyhrU+EASoaIQb9LgEEmyBPx3X8IbOCjqtTJkq/LoK8UY7kc7m6Jl8d8D4
OlDdaiWLKNGFVNdMul/lnlpNT67CdYsmHDvuICLxe8D1CkWatcKINZPZTYBk
E7v8J/xZAUylnmj0l24cm8TRCDf3MtKLYcFyd6PWIzEmuJfh4oeLRmUj51MT
C2xdpJkAs7sL2jBoxyECLLIlBE8sL+GaRFJIun7vXlpzNCtuMT4AekSxlM9y
TS+EIqsTNoPgUqkI4Jsjt4bsJNDJ5mgcQeqSnz6TT3hRshYrPpsLYyvtMVpT
Fuxe7Bdsk2R+LJzDvDt9V/auABExmlhwIuuiFXxJNbyAeC5fW7FPgaCMkE9g
MnWNapQpeZInpU8HwAH1neFC/fEGUDhAczgrJQVl6maJIXRIqMSm2unPo5nE
yyj8WQbTVFJKa+RAnU8Q/w4A/2Qbos5+toNy8YsFiDn/h9+m+Aql708L6jvt
7T0UmZfXyyUGO2QTwK5ZxhO5QIghfcfO7jOAPkbJzbhRdAUQ7O1Wi9ss6whX
eG7KiiYbwxnWXqjmXV5k+O2eHPc8WZxXzybYr3IWyahT34vDWr+maE4BVGI9
65cpp89h8oMNu3uyPoQkjCC/HXULFg2kaJVIrwaSBrO7mb7MJ3+rGMgoa8Tj
P2gHFXhdzouhVs76hDwE31Pzg9uFmagsoT2RxuisMaq4kX5wh5kAWKW3uSUh
dEJ67LjFARwu4kzvMQrQ8ReaDVeIY0J0Ma9jFEDkvJgVyPqGSozcfqdktRmW
bz+pGNXHUHC3urKNVd2FuijaqZ/8ltoq+DnB74/lmsY7yBjr82nTUDXSIoAg
fcSmYYu7kDy6KKhINMgoAzGfhO5WyUSnZ/8WBV0bLwe3lyfqmh5liuvVl1xG
tWUrAG0qVdBnrsiUtc3uMrXBABOI6fWdKQWyUJ3a9EdnNiMLPlnCsoHgfWOO
cfptoLcQevg50037lhvoSR76qfJrUGV1wdHKmdXFnrnz2c44OPLPM/nQ09tU
81sLLlIccBQUgcPGlCCofi2BT7YXYgKrR/+VjG6vPTMlnoKgGi8fINpXu7YL
b3vkkuNVlK4JNmBNoWc/5J9BLM6fNjIDnAopzL0e+w+SnG+L3xK4hNCgj9av
LCRamt5H4p/yrS5zdOYaKUrg0azArC7khZ0qb0LUcBzABcJIizTfS478giXP
gOTj3UjcIZOxdmgMfta91TET2rAJb6NRry0hrJhTevRM0/SRbzx79d3xwfcY
mBUIZ64e032Epeg12d4hKnmqCaMq2YGwwBsfIvpymqa8cpJc5Rs2hXdx+sjy
yPGNQJYqqyz0+XUv2jOwQbutOHV8KO/uwfWhh8QO7j/0RhhIht24HXrZkOJQ
mzPVsLobF44h7/kgyEkIyuLnytL9QCD7ww/9BY9z/d8x+Bq1EiRxA7MklLLk
OR+vUeaU43VyxQYZqlEaBY+/H00oj2w4ai6QkLi7epv/C52PBegLW46vLaqU
DicyCggfqWFJozInmyxPZ6NP4GIKrem+b3EvK5uGRLrukmDtQiSlgu7AeO08
NrX8k6z1fOzYKze4cYVNA3XuklID0IjcPPOTWJ3gw40Svq0rTedapZyt8Dzn
vHE6Ri0lvqOzSSn5jeLhx+1Ebarmlf9VToT7YMgMWJfkiQWGVwIyx/e0EefR
cQ/zIz9F70HZ+UeRB93oxQkHh/IC5z967GwcCxPEk9V/7LQ9F+pyI9+sJ4uz
CSTI2PWBwqHDZQnLiqQ/vRqcuX3gkyKRmSDURsmMSskrQU04EUYlpmszOz/L
qUt44qNBxfKBPTSEWd3mvUpkRQFCRHA0aNSfW74J0TMyRN0cmZ3enDFqI/6P
TmHZC6hhWl1hIkopoy423nIE2S0vaOpGPWp+gBJ5fzIsjgBpmdXZBgmyxIaX
ifiDPAJByA4ZLBXbzjd+sAGPIDYZpqM+4IwIJtiZj3zkNmUEho818SYLNBUD
EhD6T1rTThu9DtqWWrzjvnzx++dYFwGsfGcPCf0uuhmjvRQxE7xs8jM3Y+Nb
bZSTqvW2vd924IOJ7mEzXJhMo8+4ImbaN3ybtbPiHtOwtz7LYMz5ezQszz20
7vKqz444mO4/dEk1rpWA6Meh6/KcPSMnm5DQ6ZahgwVgi3xXqI9xav+5GK6I
AE5MyaPanCEZ0n7Q2qVOgb3xlNyfF0kVyBgGuT68/RqNhzy6fTf3hARSTYGA
5c/AP0ZCWZlJ7YmFv4aw6j4PQnZdhuzD1KiXmntEiEVqrIY5yjXeqAZ/zHhB
9WwtJDSrlGZV5X9suju+Jf11wdFE4fM22sbVAp5oy+OFtItgqnBjK/PZ06Uz
80iaqSAW81L7TgXKsBByeMbek5qe+47eE19e0AvfEfP2MklZ/kuDjj7fXq1Z
s4YKD8lMWLtidTHvGuvprBJ5G9J9x2DLEsEgXqu7CArlOLl/dUdqypzfX4cu
/E2JwWfguJG/2UZm3XtiggqPLTdh2zFH9RALj6/DIO9xlbvRkmQs2tUaSYKM
LwWJshWJob0hpD6zon07d+lqaS1Io1gW4IrwuiidBI1O2Jw0rajn/l0H8BQm
irSUlMMnUOv822a5w+HBoWcXYEijCUuYRt4K78lg6WzX4iAx4HF4oekjSf+o
QuO/Odz2GOP6cXrsB8aUvKY5dLrJ6W4o+dj2l31QMK6/rqRfOrnyQMCn7QTD
rkmV9yfxTqe6Li1ayW7XU/fTJYHnZNJm69gGDNH5H0LhtMOd0inkmsx22C5o
t8pm9PvUb2EYtM/TOFyk4QMIcknJYFWV9gkkpl7yao4RpgN5gmr9Wf6hgrRM
35+pW58kyFlXtJegLUgdPxFIeGqPvhGAyCFIjj8qDA7KzVTG/tvEXRt5qJah
C6wSAhfWMzI0955krb+ihU4UcQlsxzKwdT1NoI0SMAYjoXklI0GiXSO1Zn71
8CbXI8Ntz/9WYBcs5+XeNMj6ZDM9wyG2WrsSKbUvQ1Xp79B0TQqKWSE5lGJI
/MRJH/1bpE7DsYj+DsADdL2MCrfRdoVxVKuBEiXgElODW9/gufiHryGqoVCc
VjYpL+lP2SSm089MryxGZq4cLYhL7jV6J8On789Emdh849sTsOFuIMf5T8aO
IvsWGHlB3Kr9COpcaQSHagLYFV01AaRkuUZ8D5KJa3xskxknDGGs7iUBPNvw
hOZNX9yPznpdXF7PEPTcIADhe/eKz3FQ0F9aTCrCa55hvexaJ3NSz7opNWz5
6eWdxF2M7ke58mzsqHW2Fn/HXcUb7T/BJpdByMEtoLNGAuMSNldi/Zz2mGmM
ee+ye9U7S1ovOpHhVJLtSTD9KgL1Xcln0duO87GBet2q/vhAaSA7mkzFgvBg
x99bpIbs2/YxXNNJvKkOplrZV8jldyw2pWrvZvB3WpY/+QsX50eB06e+am8e
2Cj0gW4R9ij8++cLmSLQmpaI3HkM/9OH3YBhUVEQMJD+Ww9tP8ZvT2FlBo1R
0KF2eisrhOmjusBl0bmboJskiw+Yvn8QAaoTIWLJMDhtcUZ9xPy+o0exoYId
uQn+O9ltFihYRDcHkLHoGXZv3xbjk9snR1mgH2a6svTWh+WBe2kUu/a/TTFs
X7bQXgep93WsNKsKQXyQ+2NRITjcGCCfZu+9I7AI54ybWlz30zpgzXV4PF+A
iGMOsTiTCooUppn4BRC+hS88EKKjK4NrmiTtwCbMaIPE8EGyERQEzLN8HGka
O08Ibvs/bMODYGojOonwkT5QudoH/5vKUxGLgm1R2jo7uvm4dQ5661CN8O0Y
Yg9EuU7a73RkqVq7NEhTh+f8WgbrOdTZDVFcg3zQzQrQThSRGw7bD0CXut6s
P6MzbKGaN4I7qxParTMfHxvhmRMtttYjj59V7gNSVI820FLipp5aDQ/eqG0n
FgEijAHmQJXVhIPdzhgiD3YBvRFH3hQui5aJ0Dc6Znq3fFltauf7vlbASlmP
/v7O8a7Ju8y0BzPHvAbYxwDnWEa6vtnEWvJMwqk2fWmLT4R7aVIosUV2O4DS
DdXB/+flwEP/v2F7nw9GBK1KSqMC8r5QQIQtL+mPK06aHZHq7YAil2bx/nrO
bPjqUyGDeNEIsOznJ/4y72YH8pJnJk8AFwPp7bz3tnMGaq3xMLUX0vc8ewxq
/XVo7psfAk/moOO4ph/iuCvGauEUSPsiwXoMSuBQFazObSKDxTEFurnfMslR
PxU2ylA/I3Q89Kb/laKCYVJgz7q1diuXdPKI4IrCxKv5P7V6txGjL1dhOauo
6NMiOQ2zbjxOmUkKyyyYDyPGo1G8ZknK8JvB9vtJi7ijW4v1qcex/uniJmrD
GmO0X8HTr1hQQvLF1dvSO8rCTdU0cgYDd0Ht8kfO+e5W+8UiyeybRrgLk2fT
iN+WVAyqwDe7RputuL2SmIWmiyZ8Z6ncbikKOIYxxpPVd3HJ0ZhFVMnuzERg
RDDsC052uweedzd1nsX76ruLHaL4Znz4sx0PmcLPe2UDRw3BFfD7vleqcev0
M+RksndcuYmgGCbUNsb9lW5N5pX5nktJUK0XW6CstbCS9Ecvhd71wp6yw6VF
G5rQWmnsPNt9JV4f8pd7pLXHSaNdxPv4pkH5ojc/Cr441M8Wy9X7eZgsaDw+
H9Sn7TNz/+5TvxiTQBP5tn0JMgj+l+guhr1XAGmXaLW4SZS0W3ZH+6jeYn3O
eL4tl9STWv9Jx/YV236O5G1tAy1uVV0oN+HoXjH4GoMQKufnYb6LpMVKh6qE
+7Is/Fo38Rmrzf4Lbhx2wELweDCr6WutR0C5Hu3E7Ujs8oBCB6sVD86jArtF
I8gT93CKK6qfXoE+U5nReNx8T8rqQCdU9i4CsZ0Tka4ZSumQlO3lJsXXTwfQ
MVoYkekgl4CThnp+11ck1e2HP5uKH6e7llZ+5hS23slIUp/XtSoHKoILLZiL
HWqpLLaIHYg13aR2ptrnZcjt+I1fc9/xUYQ9W5eO7et1ERNNLkVRYChIZAVH
d0QCI6xjf2YcG9zpL0iVDFO6o0cFWFG8u2dyOcAnGh1qDqvfBEwcP1saqPCC
eavjKKUZsEiFg+eSdJO0X4863LFdsiFD0ao8LyLOXAvD7Jw30Tp+TbSQM7Iq
nCvntLeAKRBhdDySWXJASc3ooKXWsKeITSN5rmDFQ0S8u7fBK4K7Qz9uV/6j
ynSBVJAicswDUgziflt50s+fUfTwSsC7aBIfB9aVAz+sIC1AI9lfpgMVF/sB
l/ObPLIQ3ZjV92+19xJnC/7TkHq8e49ctQBXuCPXtQD6h5Q0V2XZkGLeh7MW
uevXnti38TwJ2HRL34Dq0FQxMNeqoYyoIHSqoDClRUCLAIbHXkZ6uTvL8Sec
ZdZokVk6c5mMycGct5BQPp9U64xdRlp/DWRkYAm5Ts0pq+MrTU4v7a8PPe1R
tIyTQiaYyvPahgQQ+B0qh9G0/4LKmJiow2WNKO+ms93C0P0eg3kMeG3ggdi/
0LM98D4jEYzWsR7398auGLkuvtNnN9JKeoYY0B/rR08Wy5P+z55zKFQILiHl
I3EjjIVUkS/hIXivqP5qbdzDI9c1df0jh0Kju3DKoE4BGrX5sU+iASOSMXPn
u0OKqsj1lsuV//Mze4LvU/bP/uFVYlThW30/iV0SC2Rh3jSuQzwPSa4NVAxc
kUYuGOqa7wRgDQSQDQw6cYMdFAiEcUNckSMEuwq335ESZ8fGyeZRnZhzc/Ai
lZZB1UlCqkOvxLwNFc86ai3Tkqmxzl7ecFTf012XNCennskoO05g9eO+6ddk
nPWbziqqcrg67T4UKontBOphpSAvneOaCIDiPeMh+0YRCK7chvOzEP/wg4+d
ZEapaVd7B+XiWNNUoQCexp7AHD6knhPhFoZkRsTgvv8wRBm9F1kb7WMOjQfX
BFECgCw8cRXhQUHflD8TBxD9Xe31Dt0yGDYEj+Hbvj2+26y9bQtnJngzQqj8
pgvq0iJqjdoGL/ZfnO2I2kYq3PmZRlBZnz3kcxdozbK9g5eJZk1i9jx+P2jS
UdvwLBoPC27Now7mW5oTMqQ3+JQXAzfiIp5qBWytxuoRP9riHd/8KQnEIxfK
5LExKVnmLK0HITDHcmIk665OnL2S54ctIyoU08tdfYy53IFIPG3fq4faExCo
w0+UWB36j1TSaOroUQnYOSjNVmNlMFfmyygBILPKSHy5FzgkJjxOVqB7v8fO
ViIAid1wn/mHrIEPRp45mBnPho74JuEGEaOx2uOM8/R+0PE8litGmzptykqR
G0zpYmANOL4EsZw6GbrDiu5ictqrSqUqhtKyYuRkrombXljeZmIN51CGk2PK
JM7R7OeqtdEN4t7Gq7rr8DSqtZMGA+oS1OhIxTJmuWKnDohiX+xOhN3jq5F4
4pYAkMxAmH1RXNvPYQn971Ih2MlMTiv9bsFFYPpeno3OlIQxFFMVG1phHqgN
tyUeZ/2+cPIm1UTgHKPmIaDeomZtmifqLE4AqVgLA8IPHCAo+FHyYYbGGlnP
GnVtz+CEcRPAdnfeWKQcz2QJgnUnOGvxt1p7x3cEZ5hgm1ShBly75/Zb//RB
mv6dvKmsR9kItXZSzh/8+IwVCh7Q3+z8EkfrrZlcZ9qinoBrS4fJ250HfPav
0Xiv0hSSbttZtQmY9cJLTb/X8F3BrXYELyC79CJFT+QQo+OtBHWIOtH54/bp
bOlolQXhgnIy6p0HdzVCKLHynjEGLN9cPSG4GjdjtAFBvtnL1p59VjWCS2Dm
zDj8Gh/rTwrXu3BgidR3gx02WPr06NsmAmN0luYh+e4wk+FGQd2RyqsazGRy
ukO0oQqiGAOkCuS1pH9G8EaZlZRWPRxvgdNI96cNuGnglVFLOMPzSxiTcMyg
LYj8U6hukYU4oCx5Af2LeQe6KEEEUxw9mfi7l9icIN1qKZkOuzi0vc9CEBo+
zubP94RMBdWho4xgsLZajR9bLsj/dj2DKoqX6SSYIA4EzBPvTf3c2eKr0Tqf
YiVxdKDF+5anrUrzuQQBfnZp8rHCGqU9vEOiiaGBOAgd7WWysbKWVaISh2zK
r17x762NDEfGd5L8zCH1uS8vrw8k+ZKI/c05GTraZpW5hz8I4m+6sEH41KVD
zs9riD7oo5t3YfKz9JEJQJ+/ZlaaR0Uh9kMQdwH+eHhvcoev+XDkSNIjrZqJ
t4qPL8f7774EwkpWWzfchD4uOl/0zRQYI8AjQGroj8vyJ4im7DDXhPL21Kzs
pyEdp8WIxHRly/fglgUhUUwUbmAuDh36bAh1feJxHAI3fxzwSypeJsKICZGV
02izADLjvBaH+YV+GQfvNtA+G3RqmG0Dx1vwYyZM5PPuofX5/krAfsJKJDdO
VUHVrSyPA+Bdyd/fXF6mhK/cOUZy26DymAExNwt4axKLO1VRa6H41bF+pPL/
Kvr8esaWm3eRk4shFsMVUAF55/GpYe9ogsQU4fqoaoW+zq9AFYoY3N90eh5W
AomSDceXkXMPCNbUHVr2/cde5kusFbRMthrL10JlDaY900/4TCp2efBLcYnE
D2iteRLEC0pTT0imUpnGrHdtTCKucSB/vnF09K36E67woLXuglNS1yz+3iCE
qLV+QyHSqV4PMgPhu4Q6a4xMWPAvtnl+z3Lhw3HJ0/kUdAdCMy83QlVQgQt3
Hhf8I1eDh5fdX8cwzPAjuvKErUM+ZBU8orkAUrv8mLfD4xNxijAgpIiDLIOR
c78Pjkd68V+00NHe8OAfELPtOCABm84PnA8cvhWJKlcfzfVBCuoUfnsxWvju
d6paxmHloughhEvlQcBRFqxWHGS3rFllZhrX7+72WnA98TKVEwIrvFkBAtMW
doEK8X1ExP1xq6So7rAg8cve6gsZcbKy9DDWPnWjS6ZC7NDPSYdTdfSGIlsY
AtAIlt0Qn3mY43/sBIWjjXfK+qK0EbeAzdr0opUxAsA1H2kqbxPSXPeUTF0G
YDeWMn/d6IJBinE3Mq1/rJMLN3/7xnWHavBQwCnXevcOWuO9JK4YzSZw9CAK
MDsSBZfuNzJ3ZnrFxqYmW0ZSKPniEj2mvczOJid4ZFQF12z2VkGnUZEaxkge
0uSCdmHZ7VYE5pL7moqj53+veEjFJFmpTD/tp+puGvGxeIZCjBQM7B2eU36R
j01cTvPaPtzkQsKh5G0qU4T0bGFbfJwN1OXONil5u7NeQNEW+1zi1arIMl66
lL5ydUnr35MjMYreK2h43zSmY5f5AkZ23I03vN75Pf0unaKddj66Ay7K2V3F
1kOeiryEqrMCmKinFewFWlG6nV+4qApFo9EuHaLGZj4ZC6QspSqnoy+4gAI2
q9fpZ+lLDr3gYgTi624RWBLeM7eWcf90EC4SClfY77Fa80RSBmuHu7tSQaqw
pTiYe0bOy03Rcod2G59onT62o64QVk08jn06rr9ZvHhQtjdvfilVk+m2+tZv
MMtcufQIfm/kUPzs0Aood4MSac5h34KETCOTvKQf6tFPdK3FgyhDEzxL8dTD
BPSt7jGEC0PpklRXXRSCLFOZ7k9nfFWR5vq1vjfsAbXR7eIgV3B4e+s1Gc5q
R+jwHpp4vFy18ppb+fX6QfTOWEPEtKrfAuq6nijA+kPM4nEYz0z5xlMtfohO
s+Mj1LcuBI+BoNA9Y6zMRVi+n3w/yIvWu57phNg1B2HghKZKeZSqMQxUvP58
tquuwMM82fnhe5I86U3rxgnm06I4RPLFHI2XeM0yRanX/oVHSeTB2/+aYwj2
dt0atqvolc1jyjH309AT78fZLQ3BLaCyqn0lMpNZtzV6ZaOFEzvXRBrvn8AU
JCKEqXiZUv/vVvfyUFbOZxMzq5PmwyLcR+WDKdrHlWel9WXFWNajZXlTzhfx
6gAVmOODNXw0+6GVdUe9dCEQ1zdVahL4JHSCL7p/LiVnbQxX9ZmsfZSW30Bf
bck4ySTLOpIX1RC5zupz9rldWGhzq/ogsohw3C/M4Rz0IxXfvUBobz3JZA9L
eo9iQM6yDEUnMbXKXkms047xATiOkJ70afV6LVDdfakcu4C+2RA3b1EaYGe0
8ZomKqCZ94MEQPy+0K+TxQNjWlYCUHCOnpnLiHYnbKEGe2pB16egUdi+EOmy
plx/f4x9gHfWQEhf7mAXo1jFBgYrjEZKb3Ek056oMEQFQseg0xq6Uo43y4TH
BUNia3yd+8arzJTuD5ozY7CV33iX3lDUHQceyBhop9fZaPQKYY/2lxwhmRqs
mFl31fCm544ZhIWiXh5evorukx/NQ654PTstqPYgWSyyDLT4Jy+ov82fyOWX
ele7VjbMizp6FqoiU1qMiJL0ogNHkKu01vtNykRsb2QA2Vr98/DagXiw05WP
G16mif0rieu3utZuZEH4qVZ8N/w9gxZuHoRUK6dNt+rkcNoJjDrXd2NV5INB
kpqjGVpvrdbOWpgajwh4VAbtDZYPNyLA4UXnp4k3cfdZb2ZvnztPFbVqgo9Y
Oif6RaHqNH1/ZrdwiUbwdhDgA5AB6j8yXBi8i+YaB+QFF/sFONeDaqxVGhtY
YyThBWfeC3k0jckhhKAuVahVVdR7AfVde8+VtSolUrQNZhYfybEAMpDtjslX
Bt/aI4/Zw3+jVutBThbU0qfHqitDpuhYiv676Kqeshgplyz2A7nNqJUwvATd
+cbfErylFKtyyi0V7AjDlz79n1L0Mus5jp4V7ri1mRBC682AfQ+Yca9y1sKf
ppHvp2V4jNgnZ6QKRQn0dFMAgCzNlWricvrxHWoU+Ux3w05L+IQpGzKfGnOF
SnJS/+Jgw6hzB1WK7/oWlKqgR0rzWSfrO76qI7vhOSrfdwpbhbWAu7sRli1t
9lYn/XNt6amCFh4i3bZNGZk5OVL6IZhYu/Ea1XESQ7RYVK/vEDJnhr6QiIfV
pCewMAE/biVebRWZDIR1sdiqJloncvcIYEJbmDOuJqgBAUO01LDbzhTDbn87
g+3ThVnnTSg0JN6kfJYkiJFPg0ugbPt0Zp15W6F/Hz6Xlm171iV6lSUCme/U
fX5kDailI4lWPA9hqed+HCkpnFDJWTyLMIEQK4ib6QrVuNeLe4raDL9LMcIC
7+zMJsfmCS+MjfarUSjNN8AUd0wK0sccskR0f56w2/9BlikbYhN0OzqGZpre
7+BSyjgqc4sFt7RIje1Cgf9htzHXOyvqXHw9S+jT0I+bmy/20MmM9c8bOsXZ
bJDZbXksYqgtMZWVbob9XcvyG35LZIKQqsst7P//AnwJznkDsKvl4IGZMvJm
S2aLuWr9V+PFVYv0FNb233aY0R+Wfxn9ckrdr5DneK4Kq6c/VEeyxu3oFNo4
TJE/4ADWswPpgDT9087PiMBn3afpq2ItdNliHx9eExhlz9wcwdXfaU/FAStq
yQYjF74rbgNVuMmY6WTP9RxiXO4icf7a+Lagam/pygZNc0/QhbuRAFUW5JY8
g8/Iqjzpnxu+0R2r/ShOsITSzq/m/ePgXkMTSgJM8c9NGOfwgqbxKIeB0YJw
fgXIxRHsyDUlS2ZXd/W0t+U8qE0OCsPxczqD4qGfWwhrcCU/HxH612VFfr8E
UghvbvW3nHtD49Gj4alO9/41uC2hC+eNsBaD3tJFh001fao6yL8Aq0ahSN2f
KTGmVZ2rCJNv90x1uRTCNiqt82wIxxZ4zRBszLPuqqk4QitXkL1Hh7pnkiMO
b1kGq+J6+H4o7AZDFyQS/9ehEwI/rURPVO/JQRgnCz3ZdFqnSQLCtLkRnLE4
ot5vVVpjcliB7kzzqxhU5dqNN+t954YDZAsySaBFxW+PF+RNoa+DmMDI4XXL
iFrlnpvB/ctaNJ4LwUvRvJoqY1DQTvVGyr4UYnxHh6DNhU+dVRULdYrWCMlV
YDW2JVycwq0CA+4RqP9twTtAejlb79MS3evUszLQqzFrSAedIdD61O2eE73m
6Q4mXtvzH53NriCdeH0TJKtoCyPtLqxscBIjdyQO10c3Uqf5mSCZu+FfhahU
VYZYpjE77bZJxfgMMvYdaOGzj07wxV01qRvZiRlbFdy3Rq/7Uob8DIHnVozD
fKGR4/yAp8v9pagPA4daryb8PxLs3TNVj2ER2kTf6LYmQZcN5NOPZTmVmUQ9
bdAxQi50UkDwzY3b4aCzv7ozrvHlCXi0s9ontjHJeZrfgeh+L4+Dfqq9KzUQ
HLs2MJlqGKb4GMLcwVS9Jq1hDMHmYw0VPg2L1ChZbdlBfd3AEaRNXS8rxO4y
Z99JPq5EWf5PaACtH1JXdAIa+sJ/c42xljTKz9nzzLuWB7J/3NWG7B3VgTy/
8iBXTKKpErL01p6crekXnVHJEnNatTmI6Y99lMkARtk0uBzzN6cilsgumHtE
NYNrACYKqHJMgEVjpd3lCxIK+XWAUFOWg37nO+Lmob1C1tgORFI/T6mSPmE3
Ys6qfpflMhGLouZlQQBOvyEK0OQLLZNuEwKQDtRRS0NEPC+R5RSd20Br/LnP
fbqg0o7EdpanZ+jNymMdKGO0x86FoFJOnEC/jDueAyHyywDXyVrltur/KFjr
uggslaogjj4tMcNoCOvcmyUWjPg6g2/zsEjTJoLgDlnEBjArWpEUFKaJQ5Lz
RHJd0bp1RJURHroWyy4a5pBScmP8Z/QIoRftuOj1io1ocTNAHpOrXXGmVcN1
pIZJ8PmCDnWQV0J5/g6nj3BB59VSHsX2xA1A44jn7Dt+FXMpkkpxvLFNrORn
tbVANKjO3pYhw0/b5SycnaalnImmtnTaYm/sO3z0uNgMCAysHp9PVD94HL6W
7dZ1O6gT+PsIkuOYOtN6UNSi+sX6HeZ1tNOE/Pom5c2aOP/7tVQ4oZz/m3Yr
Sx83ePBNNszRk91rWJJrpF79k73RFZhPGvMioEoX7a1jI255vOecLR0NBavS
MiTXOAaC/BjdFkbkRV+koMpm/SsiKp3wci1Da2Hgd48b2pPSKhqUNi9LrEZ9
UPk/ClpwoYwaG7CG7/+hVdeQHE+OeKMFWyqK5im+PpjbZ/L3d/G1n8Sozmvq
Kj2cuGHgbUriyIMeTLBn/yDZDfmXaHJQ3I4D+FmxumNoqAJ3K6/A547TYWBE
x3WWx3M8lEm5lYf1VppZO2C9UWKeJYfDwOaVpOZtbhRR9JvxxY2NBmKZjBVQ
+CY5pc5i8WOoh2mLkhJUi5t5tlfxHPMrHvnAcItK1iwypgOB8vrVXzGS0Vrd
6fygDPZkXgLVhc1WzJrKwrn5I6VOZe0+NE9ScmkaztF8+dVpZaLOEKwVw3KA
BUVv5TX9CuhRhi4cg94EMl7WOWrj3H5yA23+mTUlgQpyc7kIN5OEtykNTI7Q
Gah/h1IyS9Miqx9FYeCNc1/TIRpHBLAjD2BalO/lBbzSfctUfdbYR/s2dOVr
fQnFCpWAWU1HTptcKA+4QUTGg0q2B0Y7lG0DE5UqYQ0wBYVpZa/cQPZ0e+mF
Ud1y+ggkWo3lDEuPPaONn5TjhnbV282fmdSW5sRR5WKyX3XKJK5meh5c1KZe
0SQgnM/Y1UkmH3wdXj9XMwSE0qEwVSXtUaqaZkbE125Hr9z4cYD6k6N/DJHu
Fz60tQYoFPckVa/I8uY1gVO0SmCEQAC912bn/P3E9kUuX1mWva23XpAL/e7l
0TG43JiVLjECPxgX53mqh9Vt3pFvb92TjyXW/01EYiScMCI/FL6mxNRL4X88
fsBoG+ZUx9Yc5X7PKXytFrVkUpaRXdQdUhC61logP/63e1wUTvPqaIgnP5r7
j8TgjgffkNNrKz9+CEddEChgU0tIKUdt1jYUs8jBN/v1UH9yvpy2SETBMPr9
Riov1S+yVKcGwLqzxA0LAwiEyoZ3aUREN2EO2NNeGGHKdvG1fV+6xFoVeoIB
M0KLoYux0evA3oUfU8dk12pPPGd0XozRj61k/55THIe+LA9pPsetTBndgwcB
XwF0nUsHa7ACnxysa9OBmbpYy0QFsm+2GStFb7aREXCJ5dYlqQ8cfkyIlLnG
bCKn1tnSizHBnZG1eVJzvlmDtQaop+q7+kUgK8cl+6umCIa+nZc8K6rfI4w2
hq47zLSRuZza974GQ5JxNlSef+osbr8jFcdIDLu+jrauG6dslZ27W1vqZfPf
hMLhof3bpADcNfQuaCW6nbksiDjLIIsNsOIwoiHe6g0fnQU9u+L7IW2jhyy6
SmxkViMi89YwrSOzabT6X7XKEsaKoFp7Db7totiq57rZvNCcNhUVDjSt0M2X
aVItkQQHmflvekFzRddlHREhyzSNZH1LaXiCQyCCGqa6ZTbcz2Vn+S8QE0UA
Hd8gjTNoGFIAIFuBZZFxWBaTaubzLHbK8eY6v5oduHaDSy4t8wUs0kL1u5ss
sUaQ3HIPrCe0t4gNmWj5yNEA0rOw/Ieyx+/iOOq3Zv2p3gKseSDcEs+sRaif
MJAVNNhg77egpma2azD8HG/R3qGwF19u78dszz4ATLKuc6GCy6xg5iGvVQM3
GK9euayeGpD4KuxuJUT/5SUGwtSQp2OnZMopPjdTYWARalxtntCx1skf5zo7
JViwtmJwnU5YbXkMCPqhMW7MQ7ZBTGNI+EGEeEt8z6sJQDscwhA14+LRkXr/
gUdj8tp2880afjy3QmEedOYtx6C+bDC+d4gOsMwKHZL0NXWG36FDahjQ5Ms4
Txkv5rjdFpM3UYAELSdjWSL7tIFCyleEXPqEis7kL+FM+3ozMzHiWlqnyeYz
h2ZUM7xmXDfi5kYnSPpEc+mKu+NDNvM70lbc6yGkqfRYjAIbnBs2F8AfdZZA
ZvDy9ReHurYMd4MQJE1U8rKKxLW/3JBsqA1xUD9r6GVTVSOknY4vGflJ1oWT
o0Z1DxvkcKYo7TUpruKhKoC2MMRlfs5sE2WkCdNJ7GlCxWaYtaFYBgSwPwhj
dZlqliHAa0kGvUnHU0pQD/gjhagU5w+bOF+MUJYNTQ35Oxw7jdZjrMhFZGR9
WqTOswNJuSCchQQpoHzMl/AN2MQUrGfY1CV2UbWubGfBg26UIYRkThlwmV+a
Z6SzYQyPEoAsFmlLOWjhAz32km7JjyOdIP6FxNMiMksXVnbmg6azsOKyTOL1
hRGQsVhD1GbbvWRz0FUcagVRHjVCc4m9q1QHixRAHn8wYQMvS4ezDKNZU/Vm
ghoQVhfxZPygRZ0VAkcLiAtVWR1gzojXcW0JzyYIKrhbVbq+xoaYBdFWHIm9
dnktrdG5AJvtDfGmLpPrwVxleTfIK7bg+YN6wfErCM5bds/EKyosZrgFS3Uo
p4YwKQyZ35f+NAEXWZYwVbBv/e+lrHYKZ4VaoYp12MbeghwPLRHkQiLow9xg
9nr7po43qg6lc6XxLQKFg8wNM9PwaABsdqjNTLm2c2ZQvH8PCQ0+8x5jWTJb
tXDP4fs1zgUAYHwHRtEHLwoD2jE8gl3O9RIaiREb1o4QkGblC989GqDEazC7
FgflXy+iZbVYkqjMzfvLv1byJ9XVdLSffxrilpcm+RK29YkdZwT/ol3RXDAu
D5DfkH1/AhXsypIhvjf/xOiuZJU5+tkArYf6qqjc6yvPzi4AgqVeYbXlVs9h
lORHSgbBjKuSrCz5Pm2mcGXWz0KGoSrhkFqQ54YTetIs0EYf2UiIfvyqs+lA
RuCdsuKrSbgsqkMs48suGgrXoSse7cH+rEwVETF5p0nJegMlkX12hwA1j0yq
A7Hfxb9ro/ZmGzk74CUBbSEFpDQ2h0rjFhOnlGH0GmimZRgu0BhGBZgJk6jD
WIs456kg5064Qi6R2gTNU8KpUda/ORJjP9lIQaXfdOlBlqNbwpyHZkk5exY6
Qs2zeRuqfTGKjsuUwxijVV60KxfyImih4w/XBWxQtBmz1YPYyqscDOFnkSMg
CygvD1dBcrAyGj3TqKoVPusBGopbFB/oI8c63riaKfFQxDaS2wdt3mbTljg/
LCEvJgnW0w2L3d+g/rp94txtxkT3qp/7QJeWCS5+ZkEYLPo5tNE+diMJZfRy
TR5S77zW5apcsAQe2n6P4JT3tUeVMrPX27cqxY/wm7dedZPi2F0JmXZiFtav
TqIHslQ4OO8g3orGoGg0PMkkRcsR5QW28gjI2BucADoGWPP2kG9HaDSUOtZJ
309qqKfwPOwFMIhjwP+KNc1pg64HjItE817NKguhNmA/8hQzF4yhAA8fGs74
tvTiFycI6iaNPw/mqx7W00jUJUNq25MrlNCOFRTQgfFBJbUBvtXTbVUcsdGB
tVboWmMfwFDZ0wcTKjZ5X/0UNQeEKB1W89TB9x0MTrYWB7hABFEnrWs12/Rc
VWtV0ThkzJwo/fifGI1ZEr24c/8JD3ubsTeW3COHOA3WfWJ3hIziEcpOR1Vu
P947YOKvt6+HQwGyATJzBXMuu0Y/jj+B4lTkpfQ4fEpFy1C+HhIckAD0XhTi
dXbAa0KaSPJm2QpJDmNNwPJSeBxFMgoIwdCsCCKQ+7Wr8fT1aX3PGjQb7lDL
KzvSUdV48baR4vxEZQdJfm0+MuLgEInoxD4Ds2EvZObTYRA2RWVtbOpko9Vl
egzuNHLGCCXE6Q1KOHGiphu48cyG9dIGLDfVQpq7nd4kLnPf9bmKpfQ7bCaI
G6GKXxqiOGoiZGuQPfgzdkp7vcVwsRGWDvCAGgWCsAZ3KYcDs2fb6McZdDOj
+xmOiOFo4VGkY55BJCOgxHCAKXFzwwoohHH/ZnBfvKhwXzBjvllN1JqFqLV8
pjA8JJ2TsrF7+m8a4zO85MfAxSXv9k8jbGsRxjHRBnawtGZ2Ww/Z2h+BHff6
/ZQ3irUX20pFrC/K6G/NX32NN5u+yU91MkUUY8TfDKT6SPwRwRtRXJEzSB8M
HLCLIZGpyuAac2ijiVpk748xvTXnC6BX4xtfOnqEoZxvokSwjUhl264m06r3
sSYS2Qxzj2FMIVVVwv5BILmPhMvSpRLSfDUyloIST7ayaKWKwOCM0XAbEaUC
LPP+57O6TCc5A50Hnf2PdeDrt+vQcl+slgo4+pZUD5qfwX3otlrHoq+aKe1d
beLJgRBA63NMm4I6MLoty35fsUpx18yu9cmqjZV9nWIkZOs5sBDH+JjN7qrd
rAoVIXG9D/VuzDk7KTMNUi0SlTLRQdKTHTiPEOJ9s6zXQ5/83lZYvWYRMyIS
8jegkEwchOGp9x73t66yipyrnJ4Z8G3Ja9ucc0YzMQOhs72aeHvh8jFCpdg/
COjq7qwE9VWkSs4jm57Wf61+VPVMwb5g+3bN3Wwn5G1HIMPdGrJMaXjN3Jaw
qjxfkcXN4xlXc3RRFxaSvRwXng2Yrs8cmdwVnehib+FUISBQWv3N3LE10kl2
XScBhifnjjuyv9QyV2PVwpQx8Dezx4kxemms2BFnt+Zbg76rBAby72xgkt+w
3oI6pnGqHx3946K6q7aAkYWvXw+J430uKtWmoXsggrb4sTA8AaRJUn1/+b/V
vRDcEPMEMq8bleB0iXbE9HGqcl8CANMRwNmzZwUoPMenF6bEEuG+DtRo0Zh+
4LNbbCU7K250VeGWbHRFg1vvRzybRFk8LJr2G4/MCSWstwrQmYDm8QMi/L0y
iQ+YZQn99+0f0M4R8BMfnozPYVY7SHgOHUU0mPTe/NAsOOubu46K3CzYRCu0
czs0/0CxEOxPnPyJ97v+xnhhayGRNDeb3tlwOSe11ENkuwYmiJ5prmvu0fXV
y8nhhyXOSSzqb2Spa/OY5Xjsv7qCdzjKqxmrh7nEYxI6miBVNh8XuCPcBOj+
TALSMJmB7OrYnu9u0X8d+xxmSgXulc0cerg7ynsBBjXFPbyA4l/JeJXI9XUk
pW12xa7GHMeGPpwjyWTuJDS43Pkbc1d98QxYkTIT31asAQbbqjbsSiB3v3ab
2zkDHZb1AvFYMLZPgyKhQejLlNtgCIED8dQZHzZyhj8MwuC4Rk/vHYdJpADe
TDO/nsfq34LK7dSpkicq9q13z1eR9KEsyrq4RzysDaMlkOkGoSBz+X1jANe3
kXpMQA+wcffJir/wNSAuzwtMQz3tj9BDnr9K8ZDCNUTPFhkMDI7D6e3Jm6U+
C315SVaY2EOUucJiJOeN2DCaKZ/O1qPT9EwZyP+5GzPdeYnMWqhMEbE9fqMc
g5VKEz4L2dUWOT5nLyHbj3RVWnJE9PX4kxUm5aSxme2bQMrEMa82/iY4Lqs3
SdhehPmiMtT6b8rtbCUG/dVImdFHECQgUOcBQuwTGatMbt+nNKEIgsMBzfm5
BE7dIXe3YgRDt8WuE3QtPZOPV3bhKnEOW9TLTuduNKUjRNCGIybgJzsXArd2
MND5plcjN3VHJo0ziafE2SBjpmLHw2AqzEVJsBqwCRP2YbUoVIjLGfVs2OYE
5kZUGjzk7ZHUvUpccDmOnSixi0F5GxK32yAK+Te2gKZPYorN0vDlg1Emm7zC
YWrKWZCaHpRsIOnq5kex01cLhp9aUQei9nENymKUR/Sg+N7TXPDXrEMagKzW
Kit4rYtuUz0LeISMzaVc9AyFwhq9F/a/UJqiymi8TsqTbCfWKifHjTXYw0tw
OnvEe4vGDo0UMtQwCPy3FfxPJknQ98mkyjENBtZg2pwLwkZ4DXrlh8D1wl+o
ceOQikUSydURQG7J7Ce5phNapEulmErQycYuyRzzcD8Cbi9w6Oib5J16yek8
TrqywLj/RemAV7FZVJRJbUlRjekYAGSeKgDRqa2w0am2bA0aOWlUgZTzjbYV
VYvWpZ1jGvZ2wdaJlX0GjaZURZedObOjd8G7MnfZahLKTeMsGee3RGz4dia5
BP3LgO9HUM6SlwbiwI0E3Q1c1tmEeo3VTarl/KTJxwDmNHXcdY3WxgO71oCC
65hpEAztrvpQxLDGsa6jCh0anETVgFGMyyMI07wNj2foERcz0eTaSHn3uJlG
wtDJpAt69DyE0s6+XBhWo3VCQnwklXKvUxVDKE5OFEqxYSaqq1XILtlJVJar
jqbInXiR3qdcqqjxkWxS9Dy61Z8XmEgBWSc41nkJdjwOhKdPZpkvFVAym4OK
WpuchGlf+ul/41VeaIoRD2Vocc6OO6dn2FOWYr5GjiKFyNjAheJr/4/46I/S
d1k3KyA5l2J7Bt8WS80QBVuj9RuGV8k3ARQaXpIVDXp7CqarnE/sK7EGMWFN
t7WzymUWtXgD4jP22d+VtT6vETH7907Yeb7sAIq/MhskReonp07fwCmuXWt7
qesTdBiojhF/zPf2DJ0XomuD65QHavjBK3r7Ypf0P0zGuu2FLSwsWh+GTIL4
4AUUeYOo715PhqvWwMSXgQtBa0OqG8stumEeGShnw3DudcpuGJbIBks5vGP4
ZHWBxbZKYcwN/7yftSMVoY4UT+GLSOdfhHv4MA1tis7cywJH7jRecSPK+Pg6
KN7/LInryUzlaP7R3p8vPRwxDAPjw0rM9q2Xvqjjmc03few12iMk9gEpyyOS
bFYaOb6Qtp5MZxZjIr6j8yeKe4mQ3X2xGzKcs//uyF3hqpmIUTz4OnwJrzie
SM6tu4Mrpp2HYDEQa+1/tG0XXWBIgvDPAuQA12fdOs75ikWX65pEOAE8yb62
bdJ6GIwc/VMix5UlNFLTZjv9/3t2qtOkAmdy+w3UvOI/TAQmvZ3Bd6A3yu1k
cNCSWa+O85AVoWeAIDZrYpuyV3XxFkGYGr6GJoi7izh9tbWyV9bZPcR2zeZ1
fyiHdDtskTYHlvTOmQUvwXS3wI3lHyfXrmONpbqMQUDM6419Qkvp+4O9j1YL
1T7YaFuTHoJmVNGG7lafbYwwJhR/md6Mcg4WBPBJtT9WHY6sGiZOlMarQGzS
alfJDqKvBqS8ptQx4O2yTpKMI4uByjf101Y0tNOPRvYdo0oq4dkzjQi7NQ47
cuuocgs3L+IBzTJRdRHFwaChvsGcfbMp6eTDrTdFSIacyGqTrlPZGbjCNKsj
tzgxoXWbJ4oNRufiVceKf9hObiBMWEvFFaKh2j06uiTEWLbHk8o7BMQDauCO
qMShUvw8UdeHdDEDZuua+WvWmi74WoypHLLyoqBz+wU6Zj51Oj05Wjv2BeQT
XQbtAe9CX4p/F69sakXwvCBpZhSNXvRmIRA13nvpK71eOdFel46/jZmcFOMs
25PtmdjapHVql4sPFAiDM62dDTDcurtFZulwIyI+qXMlu9CMmmi1d+g5tVni
LY3WpioxKXKVKvLYtiR6fbLZgDXBqChcTRqtoc7ngg9w5U186CVYoFEricmO
z6ja+/vhQnp5/dXqU8ROsdZV1zXbE1j3r5/eeZvU5wIMgoRYWX5cmvn4NmuA
4RUf2w4v7Og21+OK66liZm16FFSD4KsrXtieJyfnwwe8FrqJmbvdHSNwmV+c
9QIv2wjht8KAHsVNHcuSlmoKoTFRsGNJeS0NYIJT4WUGOiGNDWRGeVLQ9PAc
FDE03zmHO56D2IljfsWPArDmUjjFqZKK5YaXl8W+p5bdXZnQVFP+oZ8YanWP
NciOL6q0JlG75Q79XGKfspx37RecLmb5iGFw/6gDnck1EiZM3rL5xmDx/xqO
RE7e+VUHG9BZ5OxpKFYs+dbpe2kaealF8d1xLcgGIZWeZ50HxozKoRT4CzU9
4YyfG08JYomMnD7/oC+e/PkHhcIRNf4OzyGzSBDBwyn3mnyxn7HLhfEZ0+jW
rBCveOL9n7TS56qWxYvumVh7zfuOTLOpSTv7ByCWFt9x75W5ZzHbiYvOhjnr
f3J+j4Ulld55PdshXi7kC2Id4PkST0Plr+hLWyipVqEI7C6apc9j0txEBnmk
mYXuasPYpJ+8v6ciCOJagcs6CVZkkmdpV036ydC+iIvZU0fCJLrgSU7acGkn
RHiDImbV+w7UBpvuV6eXYrHPzttH+un9bYjhfIAiRWsanvh5gDFR94POJE0b
TE4Ez9co1KRKV55wVWlaY9G/uFESaAx81LIUXAxoioD6sxzCZI6bsWbIwO2t
TlWOQOT/GCgDuPLHJ054n4kiHIcrb9jvKdeX4q1rixzBqfKQp3RER3AFPJzv
ehrizjfHTs4CgxAJ2AVkmh2w+31s6dZ5XkiKErRBn2DUYJq9H48KJJTN7Xou
xT7GH4h4bucCZVF3CWs+s6vmFjED7pPwHsZGLFjOxpdul1t3Y+3eQZTF3KHJ
07IvrMLCRRLCmH4IEvqM3wyxu11F33VHwk4oMd9sGtcLvyPuynTVkWx0gyto
XNRDey2ob/JWdsAR6f3I2uaRLFmd5mxqkUrNBz7CLf+sncE0NWg7dvwYjN6o
r3ONohz9eoDGFiS1yxNSpYcik0DuHlS5tch/Yks5G/g++IuNl6GIVciE5K8m
wTSFzZ34jqV0BK5C2wQ5ujaS810vhfkRf0IN2DzBRDPvjL70lJg4MxvKg5xZ
12QPvvPHILn6oxqpenm8Rd9B06f+9+/541TMALX5nUEyO2BBv8JAPDvsDG94
pKwoUJhw7QFXNylrz336QQ68aYKHz3beb2L+y5RlEnyAOOCM2ZZL4GRGGXhV
CIravH+rMctZVnfhBWPlmouPI6kwNw3JZRBFlKDa+iJ3uVsUObgkVGDNSmST
oR//3+8uriN4H3r2j3VQXJaN2fhKip0d2PYZmwynOqycjasr5yJJsUacOMB0
yV1Urm3DwNCTqvlN0fHFkbB4Xj066NOmVeIB6hN+Oz3S2lnmr443Pq7qZk/O
5at/gLX1yvs9h0+RG6Dc7IGc9MlZa/q2DYHM8lXN2OrdIc0TmxNPm6WPQ4tL
5f/X4+VrKw5qYuk14kHhx1OGeAbmMLcquFM7h+zjyiVq/MRZyCwQrfKwBC9o
FFYfUkETZ6kfM5VGvQI98jhfEs5SF9um3rjj4aNICPl+d5UGNVRHsM8OLSZq
/chi6X1wsVVgrxWo6+U52Hc3HOJOi2zuPUMslCn36BCECdZF7vO20gb5s5qX
Aaglo8dCHdlt6IQ1CM6VwHrf8rFOm8ORg91iNWEWCENBdGac8xGekkoBIvqP
FLU84wuhSBCmBGZfINqoZp7H+zmAakxbse1UOrr4rG4B1EZjWE3w0x/KHNr7
f0qzFjf0Xi3WIPavT6lbD2UkWsSyFYQRGMjZcClBpRO7wIe75cq/xfmeLsXh
za4G3LeKjNRZpTiTA3jUKPEOMXIX8MMllaoPRwi9lGAUvOeAXwH2oI8xbV/B
8/MhoNep194Fm5nFZ+9iwMJ9gzuekH9mDB7XrRdbrfdPxPe0qLZdR8+1lunz
je0WGtiErCZMysESuK2ViS5fIKoDgoskyjFW1kX/DyrOr7EgYgTwGhBNRNj/
OQIghjqbvoSCM/EBouOXOJjZ4IKy61R4oLOFUMND1HP37bBe9GqTNeedgWzP
n3IVUYkwxcyoFqE7sWuCkSs0z9/ANoOUxo8fq3eBwt2DJW89rjaWh3REePV1
X0+VxwPyI6Ttm+7KB5YnVaXyyPB01afpln5maj5BdwfgAb1uHb5t5Xgqxe5Y
6ilFrlcuCNLtmfaPJkKnx3gZ1Snsv8EUQu9RBqLXt6h/s/rCqflkCfouYhwW
pLDynMRpXaUrIFwXRaDPLZdk+3oYx6P7IbmQc7OZSy53Lrj+iKJ7SMd8Hh5e
nvFzSwofIrCJGnghLMDYBGbqBPCwImsWUU1+shDH90/Eo9HG73jTYgpBK247
xIWjs4GEMv+NUfuGVX3pBWL9NfDymFX7CZTcEsRXuS8ZDcnVb6OTND/miw82
26nVvmoDgSbo8PCDHqL+UaLy+GABcOYtCYpjp58MtPryNjo3xR8gxHoYyJAc
CKzkIuyEiXRf8RLtQDvD97IGJ4C9rOX5bK1xqcqqqktfPuWo8Rx7C10FWMr6
OP2ujk2wadus3IU20sVpkm3mQ+T5zKnKM6GoVquU7qZbOEzcaBH+yPNMaZx2
ePvV9OkkLWW/szTu1x98iQtBxT1a8cthvEHmyn8TtAmjtJXaaAdGZcBkQdWV
Q7Q8wrVUsjFVVFxbR9BHzQvTfqIpjZXOKf8ZAGMm2OLM7yvxSjeVn1ioD8h4
2lU1I9ZvyyqJnMxJcYHckIQ+JtxnTvl9SDJYd55759aX9UM5nu+Yjg21rpRZ
PcHXd4ccBvb6pLzL20Vro1AB3BKnsfP3o/Qek/3Vg2nQ7y2FyI+LBc8ki554
nfHTP5kVsqZX0lPloy7prKKgtnQBMyMnMYk8FSJBP/nt+2ANyR5WHxmk7QRg
D/V9KJrmYbj9pjUwVr6NcuY4GQM7b9eu6PtEKK3TDwe3pUnN110DGT2b+8Yt
m77KoFQXL+7Cej7DPFz6c6wjtlXpiBYmK9iaF+t22I8NMUNZ8ERgfvQutzmk
e99v860CqvorCS7Xw6On32sY79opNrb9KQexpKQ5/Wzyn3b+bUI6rQigUI2L
ulgvr0dY92gMtytqrHRepX2wUYjUjASZEnDnhYEoiOo5rIZ9EDaV1zKk6dIe
uhp9cGax6T2B0Pbd9+Dr87CHMX0r/dIaM5o6E38GiM98QQAZAegMqfZloGqd
4LzmbIhJiWLGYUTHoykx8TFYVly8zGiYX2LztYj+YZOvMR/kIYkVBIOHSJF2
QHsX+jUJb0ogHZQtKFcISnV+uCpHhh+o2U4Zx4AAdChprQBPuc0BzUXYfiLa
M/6g/wnxlpJi2R0OycyM9YBgb8uqGQOuNW6zgqUaXZ86StcItvBG/UY9pdio
5E478d65WMFjMtJ0ciIMg8Xr1b+T8X/5Bhd7XHkstJCAJutfyxPoIz+hEH9v
DPq50i+wc4LmITkX6ZgQtMMvDteajjN0k69+rgglY9afCTVIuCHx9HjIrbV3
aqytNZxdVKbcTkD8mUX5KCwIWZ9jcX8imLDCjRt7G+ZAQ/PK2W/PEIsSTXsn
B+imXB6SAxFDDjfCi4/fTBTW8ONFaiPDNVaMizOQzE+srWs4Gsz5QpGfa9dt
hOFWu3AUpHiE/xj3a30tTCQFVPjp5LfHl7y7OzVhQXidIin02GbNhtC3AESt
FO7O40u/GNeDHN8gU2xUbmK+vaa/4ni4quFKYRt1moGKCs7YVe2JXtF9M+ER
fUNRhiS6KPh6dwZUoDlFW/5lHIhyY0kqYS3fZkp7LvCd+kjWmAks3L2l6i/w
7wEUBRgilxqMBiUMPbO0FeE/CTmVvd1/H8CTtfiRi9C3r/l9XCTm1WUi2dlw
hnjFyI84ZNpI0OPREcIMAQduq2TDU7AI22nsttyyeR7nq8Q1GVuj42s7yfXO
WorE0hAgPLrrATQvdLxPpuh/iqUG5oWCd1oWW6jYPW6fAfttN/bDhnFWkn01
E+jcrv444kH26+XiJnGqC7ogkrljguvji7UJ14fy0EP1i0ssSP2+15EO9B0x
wUdsrPqjSOqvQLmEf+tJTMWkPYr9yKzRUJ3Q7EpHafqCeVYrIlLygYAM97ML
o279Prnt5kuNxWWyB5BNPawacP+3Tv//y+wFiBc3gv3Lz8xTTrTvsyeD43Kl
XsiQHD+zGy7NKwd8PWaQHGdcs6BeKVYJVE5/+mDEhdPl4R8xklfq1ZfU7ECs
IPNec2/BZKN97/8Jpck6YKOiKOSTyVXyARly8DNn7esoPksos/Z4t7XIPkL2
4ySTWpr6TPz1mTLU4hJMeDEjTLygHVborDdy6tcPZ22D0jJ87lJyg+Ippl6f
WWIrjhB9ay2IGh4+SpOcq6O93o5McFfpb5mWu0wLcHyozhQBPbjQjcFZOvYs
CcM7Xu+PbLE5tioVebI1B2majvdRn3g0aCvGLud7RnT3HWFlmH6/CM4+s5zh
2qo2R+bA2MhMgrzzuhOZdCbvOQ9jlWFsDjCiXRPbOUBxx/y5gAcCPZKmZ3Wf
rtbqVxorEjhZlDVHGHntKxnWx4X6ywrTirn2MNtlEYayFQYOEcSUBDxjXPKH
E7f1T9fDFO1JXDHrIJgNgiftpbwPHE4nm37MbYzOBXCD+OZo6Foj+ktSB25Z
CQV3kHf7A0qnAj0HDFKnlM/Pwhos5wPsO+x+qjoKlED1AxRpT+dPhza3pRRS
JE3WCmGP22CgBpyM4HgIAU+kBKCuB3kz9GnjSGR/zne4IGlLVspT1wH5y3X/
QWfZAe3YLEs4JWmImVf6dWfuoJcqZ1wMZRaPf6iLqkBzsExf76ZKalOGAeeo
ijHbt01KP9dYHaNT3lP4Tlv4IvGFR6TmwP6++yI/n/nfPhK6iHXe7FP/kVXe
qogCaVXW2fXyn7ofSTvfIA9JhWbBIb7W7oJxqDNdxwBwYpCnd04TA20okGeo
8orwx99TIPIW7LytmoZie4MnwzyQvBRhSi2WBPY2a85rnf5xIv4vuVMZcq+j
I4s3lX80xBX5R0cYhNx+5yOUsq2ttakkuVNjtxubJ/gjypQ+8szAc44eZtq/
8wpzyXGC0v7sB8a/wrzWksshH1kKf3FWHG+Pi/DJn01zPfB+OE2ig1wV8jzL
WkgD24L1gXOiMEi6FTMsQrXTaEsbOw2DmMlS8+ycHP9JGhFuuA0oQkFUIYwO
9BNTcDY0GTHRUlKUMO6o7AukMzkGu3cEu3vjba7u10HJsXbIbCqt7u08JkQh
U6XFJsVRmysq7IT1deopv7iqPeNc7fh2xuj0/LpPiz3IpvcRFtNKtODGJW3n
XU56gFTD9XnueBh0hv0qgibxTWZFzfczenGYmWZei2cJsdgX2aEN0DydMoKG
jrDDdVBd1PcdEUYEPSBZ7sTpeYNzFDz/CY8Kb6n7KAYQPptEy9WE6hVc/J+c
/j1zeBwPj1jQS1RSc9r2hDOcVLx3Cq4T03872RlD/h+H6Yv2+jgAIAqh7lAg
Kfuyrd0m+Vc0y7vrUSg66Sfoosv6an+3liIiIR7IOZsumkHCy2rj6oOjqtWo
tiY63tjs1LH8jhTF8kg0zslkLW2HiY1O2tEJgeEZMyyLcLwYVtNNsIkg9+Wy
O9nUrJp6iQ2jKC56GHtlXAu+rTLaBRNJmPZtwoi/hBO5ZMs6KWwSWFGOn88M
GELawNC9g60NPfw7T0iKXh+pclcU5FqQfZOLCyVv9JC50s24xebjAXJpwm+H
8fxR0LrSjuv2fBNsnP5T5T8/I3YDY/ikLlOmHrAUjSRiSuFURrHII+oL+WJI
nPI6ljMzfywqxzFQ2wPrbVv4YUES08FUtNlHRLlC5eV1Vt8ubkbUjJL55REi
mUce0MCAqWUJtB7adsjs22/YlS0k1xAR8RlS8zpS2Se3peSkLS1gEAQPqL4S
ImKH7eT4o4oakybciQoxac//73EF0qhnXhOQKmUU67OUlVExIzuViv3xiLJh
uPrJ7s94kKsCiqcU4l8Z+QcxDXWU2gsE0H5gS2ppfAJKKi4Zto4mz50eWs6h
6ZbNbFPaX0KTPlAAiHWczfVp8yj5SXpmGf27vrBQsdnQjY+zpgXzLF/p3+7h
68NKp3Kqf53f8AJltTJbbe63MoLf4uIebGxllDw1+yNo2av3Ju+NAk32o56e
vnHy+geCvI9vEqp1WL1razMjAUWCyux2OMK0/yeh9we6kcv8NZ0KyFtG0/TU
0bcZkb2TSwWg0ontqO4C0wtfx55MJXpBc/9z7CTE8ElurDqs8bW33zyD1NRE
mhy3oY0oG97SWYn5TQSRTypCBLmepLpSDUB9J81E8f4+gJJv14gqToRnq98d
aZMnhugdbIQzEjiHw5EMafNqqIX39I09K11nMbxq/O6vyX4Ho3gSQzKRZLtN
qDQkKgbCsltjpidwSo2WvsonxOZXPMbH23TowiLVi3pj0+AtFYfHRrlGrwb2
ZG7Zvx4uh1+D0MH2TL6OXSpZG1jKDOa/NmEcfS6rBaOPbHFR1h549/GAW/Iz
psksc2rgmuKjuE7PvWZD6FAvkv2cDrbDLVIB1ap4WkBNUVSlsb9Oeo3ySg64
CadERCqs3ibSc9UT9Ks7t8rc5ovfiUOwPTULX8tjxArcS3OZBle0sZ9Oaots
ru5g73OG+MdEkTqWKwCaPXu7xUnNlhCLflcLTMpf8KRx/piD708it+090kHn
cTFg+b3Lodhd18Zi5PEok6Pz09DZgutkMiAyBcdQT7D8vyZCqgMA+IUUxFtK
0viidEq+yw2Hp1TwuUjJIig2ftQzi3R3v0nAk5z6U3Wk+YAyrJgH4G+qxGBN
5I3tEa/nJklHVc0kFmlUj3Qiitv0EWDDiA8ifKAjoTkCXOVIg0VpxEL21yxg
+MV/kyGX9riccsYKAL4xYu8m36E1QkmK7rv0LWAk8y2LormlWtQhClEdfW6f
vMLLAsR7ibOnW5GDnFxl/wbJs2oeyxP3KmJU7+yNjEiDY2ubrFYQy81L4rVO
ILhNgI8M85Ag03mmlwIY5RpXzR9ooBrddHL/4JeUxWz/MJWFVG/+1hUELT8T
AQJvYwGwpbeuXufz5vYKVQBT3N/d4oBXt65cBsuEpsTJ/UQyA+V0qIfBErvv
6DW3RbQO1i+Ew/ZbT/Ot81ewKMO2h3cqMZPFMKaUujW3sy/WcyWA5QhsYJeB
T31QOYfH2sUpZDr7Mh1SgFIsKC/fH8GbdYLGFGl9rysd/klqn1KYZD0QoNFK
LQjJ7eeJdRc29QCcGyQrdIM4m9z2JasCTIeuMbugKmK7RX55B1H2ZU/X9evF
YVN+uCRopWPWf/b3TSrr/+vFZ96qxVGqvGMVVEwwoq4pctt1tE5BlxH82qU3
ml8YlfGYqmJSNjEnebtymQ1vr4ReSUaK8wB0t9jRx3hdlrZXLyod0seSBrt2
ET9MizqkIhc0cF0rxwRs/K0euCXiF8aUGFIusS+uulUFxPtDfgXFhN1EI1Pc
teBQ1ITUQ7rlmWxV40w4CC7jiGjEHLNmNdH6LX1I5UBuFey5bGHSSMsrVPcL
uGI6g4k0+1Iy30EYh/FBL0d15BXs54iVVhnfeoE7n66D5SRQtnrntjJVu3EV
hXWJJGv4UAO0Sv0NuvSHMkgb46L196t5tQD5nFsPQbZanLYpt4moad4UV8K3
0E8tRfBFH3xbxtzFb4ij7xNfGEG0PuV2Gm5m30DN6i4E95QrWl6BuA8vyysW
I0DyEZyMFZ1H7SDpAlAKlPLbyQFxdEJ4dHUpVKD/o/mL3d0JDikqNNwLYGAz
xnz0vCM0KpiSqlN0lpnX/bjIDrz+6bTxTXngWgZMQ7gBe/Tpyvhfr9wXhLpd
MxvPtmw0nYssVOLpcqxrjjvExtROTNcbPukKuM3DDIf4FQNaaHLLSu4KPgvy
+a46Asf7MHNB+kbnPpwVzuEykfPamodVXHFY0CEDSU7+auVZbSIrQvfL6IKw
53NkQSuqnB2rTCsR0ZeOhfO95/NxOfPNG7MwmYZudjj7EMMHv52H9eQc2DL7
yfEkpD1A49Wovtqy0MVc+VvZLXDHJW/M6GQUDP3O3onVbLDEMBWRsVFeqWSp
T8NC6ZxLC7n6b768f6cC9FJR1psd/w4G+rQjiX7BwpEk8PTK8lCbSELp/3K/
fKYbQ0KQ2q0UNnBegpBws6TP97tYS1/Asaw8xkUnNzcMDgIl2blxrm0YSyVV
tXWvAs4PxqYfaZG7oghZxvdwsa5dSFcUfy7waI9u0Sn3caaN+L5lRRZtU9co
Iz2Ci24IpfV67X9LJYViIoq3zIbrSpTPg6o/lpGN/Gvny4fxnPGmk2NS5N1K
5eh9WJ3dTYJQ1teIbd9BDwwZ1dzuS7rTmbVayxoRvk7W2ivQN+9hhYroLX+o
BMpTaChhW/URsQOPXVSFa8mWMpzrkt/rPcXlo2JUeG/zc5kBB/7qa6q9WQcE
YQrV6D3iZxFmkZa4dvOWomnBjX22skSIcsKnKcOCR5JXEoHNVfBsFuhZqdy6
5i+zazgfjDq9S+go0BXfFDMtrfylXjXIzpr1cthLfG+qGWhveBRSw2zla8Mn
FjlPvvcYHT3f2m+VLveT1WMEZ9DH7drJAtlxF5yw81QdLBOiv2SqVbfUFozv
3G/AEAf5bvpjRH475wRZeNmhthuhGY65SKHfuKmOK8uitbPTa02vkGYtKVBo
GWot3dxG4jQP+cFGSX0Klj222lV+ZAugtRdiFVjY6OsVIIDY9bOtmEKlvPQL
hhLEgA2UbADugFyLqHKhAiouxYfodjlzcReg7IdmgXP7Pc+oNj/GfUeICMsv
L2nf0Fe/tIxTFQAzF1OAp8OwaozBhPNpTSr8Kwge2EHUaTYT8qG2lRNfIH9k
e+CgMJdWeekSeBoaa69B2Dc5p1+CjDCAeoNfclfq9zW7G2a70sE1gsz0EFEB
US/1+wuRXIp9oNDqcWTatYWZFLyICL+pCHiAfW8nFbdLt1xnHpxEfJCKlxRO
8up3inU/d7UhOITCID99m5lvvRaxkB3advS29o9u7GwR/ZddnTdgcGJUEav/
ppRnqQSPeJUZP6G+9JWJPZhB1c03qRkRnnD6yuynrZVzayYXaMxU542HmqSn
DeaUZ2+Ss+Mtt2RR5vveyGKEQZgZje3k6VUDfPl4xW+0dcgTCnzHzuFtD/ix
NjUssOOq7DWKvPavA5YFWwvhnijN+ha3NXMp+3XrtmJQ7I5y6oMeV2R4lK31
SezS269oCALr+ovcnuO1wQtn+KRElDYI75Bs7rBjJpOKAKbKZ1g+NWc9uQjf
0cUALhF+Tm03nSK0JBfd9ZJSJvi7uzeHY6dC9QVMwvXpXRtdlBgClDKAjVdA
JfsTB3VIBq5OBl9+ZgeU7Utw3d0aYhHMb/G+ILg5mFYlnJk0grX/dg+ZtT52
QJNRQVmXvbanXRmQG3pLMMFY8Mmg6v9PqcrGBUUkqJz+BCwU9ADt5N74PU4O
EHuUGBTvbQ+s5lFnQMmba6TZs80sMy0oRLXf5QYyiwM4+G1dn8Gv6/erdyBV
ZaqB71Dx/Nvy3mgpO87mqWuGpRXSRzSrfuDYeDRn/SXaz99HbNmCUof+aYtG
59NGc/bdoMZqKtJFhsK/4hff1zZfJyhnKRRh9bMgbTBxjemvKykI68SMoTah
HieVn+ZeBu/o0NOuBtWBMXyTiNd4uEVqDSHnGkWDuAfZK/VsQk4u6D0AOOY0
qUFfNfo3pztJZgKE5mxpfEupdKkLZuEV10twa2GTjnaoG15b0pbuStSlPUuS
uPEdFgheCPkvhTg1buVONY8mnVFslKunOOn1qY15ybatasrJARN+6nqmaESv
hMA/cbbWDBle3f1izoqITTmJBeukksq+IIPk4UcVrZD4pxK4hCmLk1vCdSaw
k1SpDAQNack6BQ+vZVS7gcLRnaPM43EB3I13lJReot3lq39fleSPLq1MiGKI
FjQLOc8wIDZG0G4OIM8zh1ZDKAgxqKmNO2kZWoSzovxLvmQWLsPANcLFwyIm
NxvIgyFjU08IdoifA+kDtZL8WxH+TwUAIzjB0b63Yf4YBeRxpFZJjWDpHLg3
UEkv23ib+Yr8aKfKo0aQb+6F0P93ugtnMYNeLhnZMBrfCg3r2sBfCd5Pyxs6
PoRURC3bFWtKyQz1Ii8++GjN920MtLXSJwnlXepVCaops5ii6ew1iIFzmJsw
8ppVpDMrPcPY+MZDDTrmGFyHN9W7Ab/nZb9vXswhY3rAo41PfbB9pgl8U1Wm
h3lxhF26gWn3Y7l9TJq9wbgw10Ea/UivVMJO19uDB792ychOiW35500DQ2VJ
ZW9ealJ+vy2tw96BkN3AhrNItot7DdykvjUEOWLaxsrq3k8I6BZa8bAiPbDH
PuYaZrSDdsfr3NdoqRuEJLZvkX/UoWTqmJm9SuqlqdMW68Woq/h5RL6gE3ET
bp3Egxd6y6HkI06t14Omr1EDt5+nFY+7Ww4LgODM3Sht84HWEDmG2iVbFwOe
pc7zBnZS5EvSfZcPECWbwStPG2dZeURCsJZPmVV6mZG8C1k8hCprEu40RNkE
R/pvOIzjgMbLxkMX8BodcsrR08HUFyz29C2XbtkN88ik6JSfcoSjZjHvCixP
RqeutfbHPd9qEprK6bqfznUt4W+6lWbTia4Mpk1J11GIrsk75fojEbBEaatj
v0uVSDaD5/+I+qWZ0VSYtPk0Az3wNgRzRbO4EIuA9YyVBWtZ9s3wK3QvyEn3
DcGtKSZgzDFTLFOphh4LQYqjiTL6KbT6jH7+Afk1G2wmsbtdsRuZ+dteXKO9
lIj2ZdD9QxXoB2s663TYSKtenjPdHDg/DFrZfWX9zx6JL9cQ2sd/EENf4bdV
h4uap+6rfcBNClBnliuQIbMY73hOuPfSTVE4l54HyQv3TaHOVoLbW1xHmwRR
f5Qp5f/U+dBbpDSFfbicgy41UGEapJYplLA7uBvIKz+B3/qmRYI+M+ujfTNG
YUePeXQIJwcmvCMi4GOnmolcLhv7Wf/87OxosbFkjMPUNE0/FuISkYMkMD64
RIkJTzaYjrderqU3WCpyD14pyBDy1ugpR8ep1b2SAaOgcSVYOd6TxwUYekeh
mvWh6nufulhcs49gn2GV/ZSTVm7VuWqVUVdWf1FCi5iTkWm0rxlQaVkZD+Jv
NXvY7Ip60uTKEWvDh4dsnu4jHF0wUhrcY4T/tjjjgA3vPWujCPBDS2qDObKR
wlqrvgNkeP0t+H6UhM8AJNTg+bTKUjCvzZFkKuUqmZ3Vt/M2yS5hH3WxZKsw
E9AjTd8vKwoReTnmKv2cwLtCXWPDmtb4QQRWLLMtX1dTdvDlPW50IlLOdqxx
G7uNuHcQlrP4Dx5uafbEZb4Fc9DsYDzTZBoZ9uHAJ9qkD/NvuH0JDvFWiEbn
qNiScYJvdHI1qRjgdSulKHfXZieO/rVwtOJuPBARiq8QEMcV7QDHupKO/LE1
cl0j/91jPY2aklTfuzZGcNZA/Z8jNT3OjXJrQ7afFy2LsXv2fYEA/wtPcIns
9HutAlAdAHkfZ9bRHTWPt0WhWeQpk1wKV+EZeqvaPbDU6UNyvXhaNqBbt6B4
rmlrYe85cCgd8RnQtVJtjGK+GH5T+CzdrmZFzD6Vl10o6BmVxWInzOLCFmYd
Q955xRay0CAr0YDMQLN8/lqPS6ph+aXGbbiJHwWThQPLtAnIDQqKotRsgWg5
ZA2JCLZzdEJLfuXOPRjlZKBvelgCR2ST6sgjNtKcaQiST+XZaFemX9PVByMX
Unu3hs0rnGnvNVx9F9JvqC6c0upbaxrWvGY7TgFO6Z2rK6UpwSVVnSs3uCPn
u9MMg4z23iU340nDCG8mtU33Je7JrhBBbbJf7x6cPaUDHDJVmgeaULOaN294
APp0uRJ5kPoeppoiep+ksoTvBSiyW9G9tnsetluIFUtRNK2hTC6wWYRvfiRR
FYLkqNnGGr6CNKKBXIKkqCYKEAmqiarCivtuyApP8mobYBBIh2GA5C3EgB5q
jZdvVqrkaPMJt7lbXnbR2SXj7LE6TIrgm6tm7RNbaVmWAnbsQrG5Ig9fnvUL
aZ/ztsLNlaczpezcVmLyIz6Lj7hVuL49MhFIbYlyImPNIrbaCHNhqFaPNj/t
R/JiJ3olHxhS64FcVZRtlHQ/YLZN33I5oJfC9NBiP39qyJ30bsQWXzrqcUYZ
UFjwzR9YRvH4bCxJ9rnLnFj9Rel6dgM56XqbdjTtXgMV8cZLr4M4zcWJTdry
a49+PV15Vaxpi9ZqhH5Tm8vQahB/rxE/q+uyXr1pwIepiKbpzDiZJkiR8yib
h5O47WQJpe6GCITa7LG7gYOdUsYzF7f+QTcNNmnjPIwudr9XI4CCH4M1imrc
7YKIKfGRIIn0mt69kijmYhNIc4lCUW3eQCg+cokd4XywGmSnQVaLZ5w2oCOz
M0tdOsZoO6tP6uPZdEAtiQoWkM1MJcWnIC2MUQBz1XEtW+rFoQ4bIOJpouLZ
d0zyYld8+G1NdMft+Xp0aZ1nf59439TkMeSDjOdogtoeDIhKUt9UPw+viLzE
3fl+Y8bJ3PVJgeF2iBddYyX8C79F8Wv1WEVxQ4fbiPwYPuIS0n6sR0qjiUw6
Aet7TQTfWfOS/mrktpNrxVr+/GMir2lCDLjJb1Udi8342vCq1jjZ5tE8Cq0b
RpvNAzm/Y5vtQLSz1H3uPZwCWHCA+gXPf6+hGpKwsR8Cr23hectued22a5SF
nfLySVqxaWHVuEBkCzpGrJAWU3NF9DAGtB3X5OuQVrof5tZJzclB5u3yKaQO
lB6XgzuzO/exL7L46Z7NZ91q0nec75TF9qaps8iksnij+pRRsLkcViyKydZy
eTdyDgTQVjWwOh2Qsadsbiv4i+J5gKnvgXXsdqjYeq8N1uUuc62d4AzpSJ2N
yBIN4/6AFT1mbAmt/Kn1WD5wzTO+yCxL7l2rR5gT7mBvk0QJrxy15GYMmBkU
/C7hjW3GYzUBQJ7c95fYeIoQ8AaRb4WaxMimb8EQUqWjPfDYVJWHOgERXHxj
r+hJsX6EF5rXjFRwr03MVz3whP9arrhIJdujmAx7vKwU1fH6ebYCHTqu85Ui
cphmwC9RDx4xsVFiv6zL62CGgBh9Ei8m38ZKBut+MYrFcKevhiCq5UD+3Wly
r8x+Whml2fCQLSKj024TNHeC0AYBDjp/ATNEIe8IHbDbOnhHjDvbB70cJS1k
2UtX60JV2iScGWDYTMnjuEUsxQ9bCkYHHGZliufLGkhw2vWpBBbOzkTc+05q
ZPOObqv9vayhOBmIoekpTC1uacOI/HXHsZyjsQ+BMjaonxNyQOpINVzrarNj
QcRHGysO+7vfdocXnYhnktCvcud4HMsSWaIGwVzL4Z7+ZUVrtSqQrlpxOGRn
8skXZKRZrWWdA0RVRBzVBvBO8+UTrF9O2OUlRyGgwhpAE/CJIDQtFyIReV+h
y7Fbf37G/nvyTJGDCi/f18Gq2jk94iVTcO8UO6fxL0801m+E+9vp1G7gHmJR
EN5MYu1n+JTfj5XB0+34FK6HKH0xCCqhOSWyr9W1EX8X6pr+AfuQ68WjUXYg
az2p9Mz9PLxdyLZ80GxM/SJFjE8QU72r7EYj0u7o+tc7TNkjDEbO739qHeKk
g86IIyahpYL8ED5dqOzivEQ7H8NuXlH1nLRhGl6bTWsiBnhM8MSVseolFUVY
d1kqefWAEaw0Sqx+CugUiL9UQfD08Q4/l25LuEBXiHw5jSxMRtdmSRluauoP
53lAQIrcMZV/MyHl4vK334HzyrZu6s2Q+YuThzM1H7siLpw0tW6B9Pwc9pon
8/SlhA97X1KMPY1iWcHnv09B53M9wo5Fx7uR8oD9CRi9K2huPbDgCKhCRSMy
sWypl5L4YK2u4Rw/Xk177hJBta5EROc4Iu+zAUL0dp9cgy24S9B7EMWL9oWv
IBkmgQZ9L9dZHHxWOFYqo+xoDk0QsJLlmid4+zFrxy63vSMYqT8Mh9xgatar
KyyclOeI5frTyPrFxZeOZhhtBx8BMSIqWW7ZT7G5Sww11lZIL4RljKHYkFXd
lZ+8qG+t2txb1PYt0BKaKkRLiW+ec95/f8uIXIUVPy+cS02VplUHckPr/jCn
+fpbAU+PQXnoPBoHkWt2RQMZ5qQFg0gxOPg5RzltG0S2YNFXEcKUnz3CKzlj
QyntOateS8/dOnhmXeIYglzrxUfFct92oxHg8+KZmx0xFORjZqX+ObbtT+g6
5JdMt71Lic6QSi1//5q/6zIcCest5cbPh48jQEir1FVqaznlmQ4JKhP4k3CT
AN+gJmELXjjlmwJShArWW2ceYYbFRpEGPysmhrh5OS7yGwPDoRCHoyRYrAQY
CCHvgaSAZW6z2EXpDRhECxRsGIZWcymhA9aDL6h6I7EFn8eEndAvBRVJkee7
iILMsCzE+w1/Z7lnmZjtNj1vNpEGu1oYLOYxHoEVVGe66TCImhKKGIF+Z8bh
munceNTfkIlBKppt5asYXwsC8RHrlNU/dFlgqumrDGJ4R8LmIbYKCINk61kb
cWVSM4JOQXwI6WFjFCaQK82A4B+IxefLgXuZ9GEqlu4s54skTDGmE5Wt0fWn
Uzx6J6GXrglmqRKyA91FxoaC2cfukNHtIGNNY8luf1GSTT59Fwu/xggorTLu
9Ajt3OvhJu8myP3RsPRFi76Uj9jkxNFSdUMUm8V5NIthi8lqMCG5IvDAb44n
Rcg5XiT8LmCwsTUwTcqBjnHZqM0TpPydC6zmdTFqFmVsfw8TNIYo5N/5DeZ2
6YnAi4q5oxNKn8I5pgd9ZyDFp5RhrIXSvzxrceo3ZE7bxoxXFRVrh3Vxs8WQ
KK4JTUDAf/sYh1fkjKxfGjH843IeUjn4yGe5iurVPGA6R8sH/M524qxouQCj
L+xEXjFBbRRCxjBU7ovYSMjzocmvQOqvXdNRtbMCFg3clTh+WkgeJ7CeIpl8
sBoS2+1+X2Qdil9RLzwm5V48Zpfb8myy1DLCV2jO2XHsAZWwjguHWFDiym9o
TZ/MqlVJUwZ+mgoI+ZsdgpZX9CVNv1+tDzOsUsBIqC2TwKsPMlssNzBRo2CL
FUgcFKb5blW5t8XlIgp99Vo9UWngqBf9LVK9UAZcee19WLa6bSSEnEHvdxuA
ReID9jdGG9YV6ASfLP4gIvsIolI3aVXj/fBPCbylrubsqFk23S8pQ2QOIvMN
korQZfX0useXyXjjbmYtm0LfmYx8ofuaxSAHeX3n3QAelUXnZt4R7ajgr7G0
rvBYDqTsCNJ0X4Me3M50/DXeuO9cxUj24LWO/RYrJ1U73PxcVrWIKgnpB6zX
Xnlhyv3v/ZiQ7/BcvIYNpWxPfpaD9Kmyd/iq+ggABN6juxq0+XXZG7retF0W
+HL5sPn8gVZ7MzZIB3mz/KhOLLwzyoW0UqBdNj2Nm0BSRERJX4RTIPgPGHm+
OaCwM5pq1kQy3COZwXGfqHL2myL1khPsaA3soLBYC6nUCC88dYxBzdeDswN4
UKx6bDLOI2X8Daa6Cf54j71yXCWniCDgkiOefQEjD9f7hX4WnxDOIZKDHKnw
PxkkLeuUlOTSNXf9Ld7NQaynX77u9Z35A2Z3QzxE5tN/C39QFxF9kVtNkorU
6tFZd8bUXD2sga+QL6qp308DUmqpotLhHlyll2VHRNKt90+q89oRNllvy4mS
0eWcFRCyaWuE5EBZJAdtVJKlxR+cju1L3/W3mSv5IriaR6EEqL2Z73r30HTN
RI6v7BcWeCqLE+pb7d7yIBDsSQ+TdIZTAgBKKqSwR713WoXPnggIfItpvpoP
EokZoOGaxJzj3AlgwdMMvsGb9A8B/1BW+zsCxo5jX5LulRktMaeFX8Qywdn+
z/MrP4ay5WLHexeeS6ef0/y2lkoPucMYYUuziiNe/7wqsRK0CZN1AT9MWXyh
jJrCqqz9rjac3AQAjWNj9nQrf1kx6VUjdhL2eSwtalDh79lPd5PumtW+Pj6G
PTg9uGhws6tlBXfUUBmb0hIjP6zUZEHmIsYeU4KH0kZE8NL1Eg8iUrfDGMRD
x16NP61f5Ym0sDH9UXx/8ndAfA1M6xmXC8gzqmjjw2AuNOcM3+EAtwAb3gRP
LAcbacS30ehYOT/Gmh6yo/iX1s1RGL4zJpuflUxAfd0AP7TyIcF8dBz3YFV1
5kaWj28docCwKY2fvigYMLZFI9cVlkp5BsgNanY8zRDI43lpkul3J8QsAzYn
Ld+vgqY8+Lt4WHwMGeZ3lCELIFSScLytFyDr504HFJZsQYNC7he+sVAHjznJ
08v3K9Ehj/RBJ5Zlg4yCkgbyrD03iVz4uNbC0eQ/uZLSCTCVrl8MN+IYrqZr
qJvfjXAiTX59MSk20HaGsz+XqwFgctDO9hE1256JzIsqHkhQaDPckPdLYFUV
qEUb/rsWks/r/z7gGF0j4eaolLFoSSt9XiCS29FIfIW+jN7euLXChqGkZA4P
LVHPeF8iH7oz/7K34HvcWCXqVmJL+d7urep+IODPL5It349N+p4bHzWCWPeb
gqN2m8bhjmT8tkXpMHMeCeG9FObso7JWqVzg22eThPsyLg3GI+OM7ZL59y3Y
EvUzSHGUMh/6otInNfHuad1QSTN8sl19RD0uA/Xgsz9ujy3mLma9dJgMs1pb
rauNa7qmRn0b59udpiQVsMBYjxn0W9W3Dvduqf1Uc/KtwCc4b3/atngud+Qs
yBh50tIccILpRTLlWSGhwNHO4XB0tOdF3kuRdiwXJGT7wUKokgGRJy9vo/5Z
ygOvxcD/Jwj31tyi+64pNJjTTmaHksZYMWUiYofIkNZ1j7jGImMbsHQQPLFv
jU0ISaLIhZ+2CCWMY0l4asynfpK0AAjgEskYaT4J82+vfm+3Cs4BmplPKZKc
kkWWOAqtTAx7aE9sNAx2YwDDCebbk7Z7SEGqcg4bTS02APdvx7VSODvzpttO
buMcZRbKQn3UsuujvdnxdQzKNk2nvO7T+8g65Kpi9rz41ckqPLIMJAyuzyZf
MPzbcgoVg7U/gC5IGLP8G1dxVc8443E0gRWHH6406f2yOtQ33T8OeDbNj7jp
VPY2rKkArKHPJWJGSzD5LqzXgTEdlJ06ExIQxO3yUfKB/MxP9y5d2sMtqV7k
zKmPDc2HXbKMw7MqTVwJPm3c4FchvZ1SndPfoC5aDNKH5xab9sn3/fIWJgkZ
dcJ1kla4LLRBiEVFNb1Lx31IZZxEkmKgMrbXToIYV3yrLXsqs0mJKUfJUoSm
5cexAwGsabb1rHzz+VNp6BJmWrp4488F9HcPaQ/eRTgGBiel7d6H1rLlfEua
B4k63IZ03QqO1CAYuGGvBvBCYVDwIEIAC2TfWOXe0/h3GMYVweYlhGuo+F0J
KlLdDXqvhyS/mqk+y7XQ14u83ovAgReF6lAY1YoqJ05NvYX8aBmfjrJ7FVSK
WU+KrX5lG0techONZPJ9BuwZ++QIAYqvIRiYO6OD3UDZDd0R9X4bGT8wE4S3
QZHnFa4WFQ8GTW2CCmfGY+6MHppfeNMFgvz4t5krX6XZhKKnHcUi/lwGMlUT
piw8WGsI/J/IRx0ck3Y2kOurqwmVT/pBrACx23Yu5cSiHjhsxrrMcs2P8Hyc
/UjzPiJHyD/4bnGieSpng9ppq3ultcJuK2F62C4/emCZFCfw4cSxcK9guveF
oGkQFfsJ3wRbqx2nsdOWnl8GOpGsRQrjz3j6IIfGhW06ce7XAC86R+8YA506
G22nZiUhkz0u4ccLnS3ddpWwRhzehesQKdWNekaGneZ/xBDSW15VRXq9r2oC
p6VsvLlfFZDUfnWayMkHUJ1j0ewEblK8yMgA/pxgtwC7dNAAFW6Rjr/Lo5JI
QS2FTMVnyzKtHR6lTmQD8hPM22Zc3TwMPQUoaJXrKHZCMiKobUyYR6WNZKA1
cpLnAV4mLifayRCEFwz78ednUODBdxs0FbkKWHmgG6vNZ9MfOMl+BIXlvdtK
cF5Y33MiAiyNzwgc8torJVniFho0UD97IdzbzZaBkggNbxvUog7TQvJN9nOK
N3pBNKgwShCfQPcoc+ir9/YoPXrMzgO5hX6Lgtnmhf4d6kcTHYZExRpXKhdo
Ll4TK680ks450DcVmsHRau+QWL4jGqm+2DAGItdj9Y/6VN3WlNhgprYbTLh5
ih7574PLVtGWRS+EIAxgj6hi6rk6BlfH4xBWzFzc6I8UjCpt8HpMPrW1pizX
RjhyooMX3mimxMam9MUMQbBZBXzoD61joThx9bW31rRVniSwDxKI+odh3o4K
XoZ2pvucWcIFgnC9nEpf5kTiTYu1OyHOA+UdcOJhsrnpM7AvnVbLvTWWCKV/
8PBCR4l9bww+TJzPha8locxwwEYMvbk0LH7s4v4EueMiFSNLAeSFyh91EEX2
mG50ptYBaENglgsW/ugVK7fkmriYqtBsKklq31Y+0EhE8nNQ8dwxp1Q+kXLJ
XVqxBnzZE5iE0mXgzagy2H0tkJtGuhJrco6BdQNW3PosL6/8Z8IVwv1tCsZ2
89Fn/6AjxADsBp6QPqbiY+/zyF3nX8CAz4gLcXZD4cbdiqOdh2Hc0apKX0ns
4Qq6EPVeFDMwA8GmmVuSnhN1BUO3QxSaVxWwFP5WhjAnUSRsOckBAcyz/JBi
OWdic1R21/1D2k/wAx+SYB7pq1i4cvbtzelzQ6xhVdD5nF4R1Fm3f9Jd8Iz4
JYfJ6pUC/wzDDVhRKoegSoByBv2d55LYIwLVdki20HCn6HdIEzvpk06NhPm/
+QpaXFW9XSdg0nbb4ZjsyXyBD9wmppz7lLzbWOq25QBImpx4tzABHO6x/tB5
KjmBx1nKs8U3NRh6xxLSfGND6jOjYwSNytlED3sCzsFp3SrOefm4+VWZJSgw
QhUn4QLv1xECmbMe2zimqOdkpknj56Nfigaf1nxVFnWVDIJbORoBouql35gI
tjqdYhDYEbl4SfjT+Swo9nGa1sgV21/7usxXv2tJDaCWBW+/M9zty7GjFlf7
N43RAYH6jyucvphWPzEfI109N/E5BLuPChdrmrhZW2eAcO10VowNverpJKMI
K3vw8MJe9bjdXdqL8h12ng+xFIUMxtnF4G57ALTdNL832x40nkea1dVyB3K/
UnvSEkFU7mM10dxCe4q8C2emJFuNhoVrVzpJAnfCoQ7cgyk6iP64G0YJ5iPz
XZmZHghbAjR1fDd/n89ch2h0/PQOT5yDhChJ9aJw8BKZoHerjaIHAzIAeNIn
opAPFrlZnPCA4FgavnRd/NY03K13vaMCN59ezjh1Ow0ZFmq5ryYmQ7bCvnfZ
tWh+3fq88dHAOVHeDAK6Vi9NJ1eFU04qvIW2G8rOzG544fDf9v+YVaJsFbUp
DI7TP9ZCPz0kJzMguV19lSrAv8nkUkcHlsiFkjfFj5f31XCQl3KRBwJJmT6h
FMLAYzJsfHLi3YbQPUYJAwc1ClhK0gq6vNr6OWXh2Z4OHDhm6tStXa+jDYkK
DQL5tWWOmzeJT/NeI05Na2HulDBFkuIvRxlB9h8D4JZKCVU5W5d4OkdWcF61
PeW8Wm1QvFJsQkumt1uQvnNwCtZ68XlLkSvVgvzknTy0iPXApb85Vyz6XPPJ
FzlXeYKTQ1Tg8NTo4vDXg51lHBxu6uwAqHXzQBX0CF2X5zIMJE9HFWjvdEVz
byO9QTQMXYh8v6xr4IW16LekDIotIp0Ek9WfBeSU4YOBv9BvBb8hggkFnxFI
1M4pMJNuwxp7MspOOz6x4M6m9PJaNbzHZQGBUcbDp4DHw68fgGHuPyp6hkaX
T8Wb1AFu83IKo+VBOCIzahzgBcMyjHWo4JrZcyU8L+K9I3JR7lItPNhrdjdx
8b4Sq6t0tluRgCYgafIyxVTH81AhAwQ0weGviGUZLy4yfYTvWbiwhX5HzGzy
x33B+psbiLleqbD9Lc0luoa5gqdODjlwNUwOnC+Mib5anmzoudZkMu3Y9J+S
N5UH+S/PnJedfrvcIS3ZXeGg/DoksKVXzaoTkLUzrd1o5O6b++7WKqWRZntw
R9Ldqz45MJQPtRgPDHYWTd6DeywfRx6GtNRpwTe+sGOoSmgp2r8/Pd6txcRa
7lMahaLihL5vdg93PaJIpYQw7yrK1JHAxqoo6sNaieVpffM2MUzR6kcGfywg
4UBEYfrSAerPxmux2i6tjbudz26Eo9KJ2KcfLRl0dvKs3s8C67fcWi0KG5fl
/fE5fQQDya5I6sYNo32xoNtAXItNKYw/+rYnFL7cdyjoRM/pFTvSTKs8qAhy
Sdd7aO++9plApbWOV0j2IVY1YabyliS2mT9vyCW0jduej8c6+C3MSJ9kf7HL
1x8NQFgHO7P+WcJYGtmqLdC0/1n2HL5yL1DlIdZozGtcdXr9g5XHZxNrCDEF
qzXX3h+CrfnidXHlql7WXwYu5RqKlco/KzAEvO2VVMeknnVfBpy/PIoP8Y++
/sutVplHgwFP6QwkxDJffqY+O3OaZXsMakb0ywsGoBMK+EZueEmD+LGA6Lmx
MyDYaZUWwiOolX2U6iILquS2FmlpdOSntns9Mic9hFpoaMYfjZ1ORCqPzc6E
H+VXdh4GcmtXvpjCuNSEl+mE1SmYbhtrptAcEKaBWxpmL3cKx4dVQX46wP1o
S01TYkd8gPI2OP1Mq4BZ9ooAV1LSwQAm6jrwCelqY1O9MBXmV1azt/Ijvf8h
DUQnFCJeoe1xkFxU9AcbBS14m8sDX4LolYXyf0gI6n7vM4/B+g+vfjz4xanA
XCZpaAG6+hzckF/3l/ZMv9GauZ7UdQLmDPzzyzCrb7YzV+z/O+E0xnO9p5Wb
4EFQjSAUxEKQNkhCDv0n3i51iRV763bRsqG5V9ct6M/cWIrvRjhypskZ8kK4
xx3CW8l3x6dfEeuDi1rsIvDdVPkYNtJTEC+ZFyf4O/0pz4LlxjWcutIfLyOR
t+Y8rpdtSc+bGko1RlnPq4y4SI5xfU/lO6xt1Du7CPh6NcytkXap8y8MUtI9
St6SMRF2bSx0ISb91mkd9KHSDt3XWRxY3nDDc8GtgYrYFUacTntDn/9py+t5
qmwovg59fBnIhC74S4rQ5c3u5iQd3yTAVLdP1iOVxEKnZQQGki5X3Aqu3Y+K
lQDOvTuY0P89HEbbUSXATko24dngquRxlpQn3LxSShIJIx/9vFB7U2AR3eWV
jXGWDYH87blfsDv7+ZikmldPN36fuw0/TgiWQuSbqBsyqz7Pm0qiUjrRaelb
wFNNhOyra5QTtj9mg1iw2+/FoUT5xKTRu8NxlVyhkuadmGxuB6wPiNQe0la8
0ZpHbRJbOaJQrTYMNkL2ncJjazACes4If+Y8iSUyamG/yP82rVMIMM49IW8x
GGDGjheKXGlFbiordNRC7zxuspF3MBoOn3GvT+piwGjZupg4/ErsJ0OIyce8
Kz4Z/sAWDHcc/0EwyT791HtLAC/Az4ltWO/KzeCJOkBun6c/PTOoFF/HNAcg
72qkQjEK60MkuH+Il8PdcbieCr/nzlOuJ+HdJzW4ZD6RcD0l3dEAABWv6uvs
1ylGQARo9RNrO/BbTiKJELGRf7Yo4HvSPS8404/D9d9DbOFxTqVLnbKb5HYm
8yPn9RhMa8dIlpEAfKCV5BkcLWdYiVT10wlyyEMd5MOD3dSV09Ga+m9GATsL
EUmu8ySw9YBlH6IcanQbldO69a6hmX3iq/l1qV2Pe7pjvomyr4VC9EthXdsc
AKeE1r7lwPuLcf3roSRey/oG0CxZka1TiIkaqVt7H+qbMVqNE41Hsif+5DJF
SKuUrQqrQ6cHnY3Z8NekC3v0ZX2n0xTNd9s8Q245piqA9E2fH43Djv2fEzKk
XCypusLfKUX2L4ct5+pJcOsm/p4Q0Qw0W0s8UcxafWIBBoDoK/yM3nL6wehP
doL5XPwUdPEgaQWo71cOzuc6FEv3M2FOyNfMRc983RLpud70JPPlwh2Dd19d
tIMdHUsBAW86MAFf96ygPzQ6P2MrIJ4RnU7I+cJT4Bpb4F1rgzTyz6jI4gia
CRZF2uwA9TYhKd6MC3UunDohpkfyNO+mdwl4wVSxY5aSy58W9jsxS0z3rRJd
uv9eK6TVc1ZyD9SeLXaCTB6nQgwBYz0+RdrJei76U6rj2y2JjcAvAAmrlR08
zo6B28hB/Hb4LVK9j71+l27pV9vzLAFVyxpf5S6bK3fBq5YVw+/55dHoqbl1
PQrrsyW245x5PORSnQp5h7Ev3yLZV+DBnHr7FyKNLhdUAe4Sen2b/juX6ogn
7wc1c9uwC7sTPHZeUqrf1jtSx9LdviyA8UejPLlqqaIAZh/KzzlsP4RXogeo
k34miP3WAJxbal7rcjeB7XqdWyOc76kySYnZ3OUyfXHk2L1hnqqtBdLyMuXs
jfoyIFWP+gLGDVeFTKTftBqafrr0u2i9xxfnyPmWVZYawWiiw29EIYgB3iGa
jKkSL/8W6dBjkvQCD+ScuJERqOM8zsJWvULpEG3r7p/N4PD0X95D2FYOuZFy
2A+ilH+NRLRR8R4rXRFs+TULNHHgdPvyYlfNUMRTUZ2iy1lpL5p4lZFCKfBB
A6v4yH+LqXdhlCQaaiU1NSaIvC4zf2t6d00YJcVM/rM3XqgTzmXIqtHAGBjZ
jYaRadgKZ0K+6jC340R6GFyHLpUZIlZWd/mUKpnIwskMRaO0f85+0NHZSe7P
063/NbSX5ziBCsNgVpnn9nfdsjU/C4G+mRoE2CYp8bRSIgO5Od9LomjWxA11
QKXj45TQsO2qcdE3UBRf1RSaylCaD5IEg3NRojF9BF9zbcIQNiifEEzLPYKk
7upg/S5Z+NOzpvyAVpnxQpW99+8X9vhDLcXgdgl0xW1LCFynAWbX9HxC/eGr
/ACevRD+VTcTiT5z8NlBmYLz3SzWcmRK8lGynKBNjGjUNT2dbGBF64tLI+x4
KSnLi+2uUNARG2H5R+G9d3q+auGmfShqnJpXqDw3zf51WbKyjKgmwjyRc8pb
cSBP3jC3y3cAHgavOOa19gtd2vhAAJTuuCUAKfvQWx66Btz5F3OQN9rCtH+x
LjyIdeQTFs6D/pvoGCRD8zWnN7p8B6iV63/7vdIs75zksaOwbdlTC/njR/fH
WMHZIkMdBeJwtVvUc0FNMm9CZ7L3cJtClIFl7rnSIft0zqgHmVDejuGfNr2q
ixRSkmnSRK34IRr3hrJ9n0oBzrp0fEGT7oQSKxOltoib9dgSH0ol1PZRL9Eu
lyh9rlXZw8VkZZZkTWxy92BvPZoz8DeQg/aAaEBQd4bxdbh4/VvbuCI0MYZQ
u9obNYA9FKxeSx3vDPUm0l39Zj3ngLxGgTljGPj9TnAlfxUGNl7DbX9ez75a
W3BI0g7jTavdaI9PaXlOwJUHW6IWZZEFvpuMcSqdR/I+3vPTZ5zLpWUPBMN+
YRqDSnRlOL8XlUMG6mhGb0zCUWDfy0yyiwuDy06Ju/6MMsRSHCUEKvDbur2e
IeuQl2yHb5d2B9f0qCZ1K8xZtAj5hSnu6GQPrbKXnUmfF7RpRxoa26eJZwCj
M6Z5B6GXZUdrGl7K4LMWleyPJFrFexORtG2AvxqnOSrsz8uoRpuNut6nsU+2
CLx8+EHTKb6F16k3CP/9ZdjjNowLFdyPGYO5cfBYaOkuzYjAQ/E5SGbv7ZR5
TUtIm//eCSaVrbTJB0zc0+JeQl+FrDX8fxu9HIkrRL5wzM9Ig0Z6959n30Lj
yYHEYEQqU1GvzCNbq3OHBDWOBywX2xlC4EjqzrjFWCEAY2ZtvHQAyWjV/KVx
pKCsuyUulAqxv6h+HtwnFisk0Q/N7heJETjwFBjbbwRjm8LT4wo57ikdJHvV
cRuoN0sct9QzrhafaJjkzRWNsH6UWIYQ6UFjZ3BK6rEy2DGHTGiIo1C6SxZ/
c9xqHP70gBUWpfKrKPVafRHr+7Enp+Ap7WMs2t8nqDdfBdyXfc45kP3eM14M
ORYISLSDXPi/v0a0tFX5WxeCeJ8DtNrdzpf9wKuKeksPSHgLcEd+ZbO04lUH
Wx14nweSRu5q6hn89Bkz7Mz9qlsswQ66jp7IXjX/hGQ7pYV2f9A5YUIPWzSY
arYyL4ErmU+IzW7A/7rK71zlCUn6xLt/yh8wiN5iOouikyq3NuxPK/tY6Mhy
UhwWV+jRrskL03Zd6NO5vePwdelAKqrjOf+m9FJLXx5Q7tmmXYDt86FocJc6
rJgHJkHnJZCHtbJ3TJlVTnOdPPYcLbqAmpDSfcMmYTeTHVsA9LCPdNtgvp0T
BxXMEw/3J6PEggs1QQga5+Okz/3avm5y21TpEfMNMMCjJwSIkIWQ8UrSAoOq
6Ubijvp2KvJANy9Aw8z50T7w8+vUjUBqLq6+7+3yxYtBlmiuN5b+a8+wviSw
sqsrY5vxvC83MaDUjnNm8zRXkUc1DLieJR/mQfOxM5xn7a4Y0J6CLudve4Id
eVLIQEjRbJcLdlCEcJEY5AfB34cogLgxutWcOn2Iw9r9XgJUmhwKc25+M6ov
B+Ts3QLx0mjYe7YwkMd5aq+RKdyno9z9yV3c3iilrxzaIVNTqL5k2xUJ/7Wf
xNIHQ5VlR4Hv+9TA2QcCQVaDv9I6QWJ69RpV/47oul6XYwrROCtEnetGG4yb
6F1bUT0Hxp3rTMSaa2OlvWvaGI8muT72DByJcsope/ARAt8qoRB5yE0ZWGax
6Qolh428HmU/92wfjMRJw8CVMMHpYh0R/1uJ9RP6exuA7WbCN98vjFR8wwlP
9cYJ/QvMN0eu6lSD6EfwhFsfxHtCd8UJAXMuNTStplU32jKmApOj80DrJD/T
ihjK8UYyRO74Q+h3qwUq/M1fVa4+RZqJspQ4qSV6h/ChlYPMn1ieMbH8BvSx
HSG0lPhIsrWji94Ov3cosC6PRmVrRcOMLPtGiwD3hT5Tr0vRfDL0edIzqO/O
CqvKzuHkKKabKALlWPH4grtxvImk4kC56fGZ4w2lRwDmVhopgVgW2OVhRXhs
I9hW0L5Z1/v8wGNEyNE1wnZroUdwre306Ezbch/lvBnSTobeKbRaS5bnhkaP
2EaO9J+wXMZahJASh3YxOCahKZgoBZKEwsQQQaJOS7ExoCGE7s0aIlppKx7O
KpvxesTpWwRIpP4S1mfXtLYCbdB/icNn3c2f6Di7x83KInF2ZQrEPoWCN50G
rQvcQvBAjMUMSojz56+qC38ni8eWW9HP5jXs7eLVf8y7cdhwDgOdSqXbzuQj
EY7s9CrbN25P9WHKRKa32IldUV6Sgs3NfcYgKUzO5iSE9Beb1cXlk4hTr9W1
9OBMXCTt77GyAgSlYaJLUEWrMFvtwjpbF8vBJmNFIX5HWxmwEPTPrUenkAVQ
oZ1unQ9WFTFX33iuAc4x+TmsmTZcQK+CYhmKFYoaKGkZxDpjupHi/x5/O/Xj
0F7GX02qcyvG274DszpAw/Jx3zZiyrrMrU/KNEc5SQYxegmji5pUw7BuKLQf
2KO3dq//CJ7O5Y2sNBR6xF9+kXFcnExUaZC/sVOca3nxKs0eW2UBeOjQZfyO
Oqw/s4j4wJB07d0yL5RBCZ6GsJ4UnswC1XuqrolAIWGcB8ktxSyKgeGi+HMF
TDth+wlYkdE3AVtNoc2J0bZJbbq2VNK1xW30WhVJJw4xQNztQ1g+I/EZ/75B
UH4+lPJTi5a45jmmCAxbnsqI+v/aRJisE1cnI2311jI3D6Au/lXCIV0yl3+V
8E98F49ER/pamhbmOpv/DxPQ5nOmqtuyNCodBaGttJYzS6P2yiXBFWwRSS2J
IJUlxrsX9nxqj1XVMaAj7UkQacfBMq+Z2Edw1x7wL5e9Tk/2NDfnGBBC/RZb
hRquSKMeHwJwdOwOg2tqNlbmF+nfRl7FK+rIjudkBlt7foZtsmFkctn1AjCH
PgboLninUiwOlLfmRhjdzBFUiwTbh4duwi2IFpjY5NwSxpc+gZJ1ihJjm3mP
CJ+ZH/QqeTFy7Rew+A8OavIPdliTCC9SRrrwgP6usKN1kKSL/dwKXJ0wBFVY
EemHUvMHAQal538vni9FBKvhpdJiqmYaIz1Fz9Od1QZm9k3GSaro33unFZw7
9gwiv6Wlzirdz3O2ToNWGNWmcmpFM35EEvwD+Z9pDbYWz5OXzfhTbYss7Nkq
SLqnkPWaME5OwUym3cBPeBiO/keSPgrnsHs4oSORsp3K8O3lbRRyFZXv/rti
efIB/ojeD8SvK6A7eDVywp9Z8HJsM4RpTxRw+noqJ6nwOsVOqozW1zVBpXay
30iODGUMsGwGTEXomOjaObJZrmpRHdOom+1GK2OAcxgGSO9z/H+KVhfsacBR
ur+BvTjxxthZtb3PHO2yry2XcD1Z5A+5YLSWaLXPCAAagUbStqTNdxmmAyg9
osepG/C72JBy2LdZhvZ86BrK0ufYQSKGQLZ1XMwR3ZXoBPRlvourNw+EP1ut
X8OrGC0tySWYxjHDNasTbbhUREquchBpwvrOmivwfMuyfVE632XqU4mTaRwZ
RGtBrmHR+f8yuj8Bb5+rrGGe8AkGBpC81jGEbq0eVkVUyu9mecrEBQ+wJv6A
s13HrbJOPFlyZtR9VsDpAFTpo3XOi1sSryfXd1V2npcWayZBKyzXN71RA3ng
PpL8jdwTdSGb1ZGQNrNFVdB12NKx5HNnG3k1umR8ESOJjMUV24QVlzTl/4iR
7YymnIxg0tDuY+X3hwb6k3xdMFf6Vwst4X8aziM/028zrCVxScWT0fWSRJqD
bm7//wSfA+g1r4G48D1dXPRtPwCLH3z8ZbBpQHXGYP4mwqBXls+w1jNe7vtF
fbTt5M+PjcyQVCTWhxXDDxkB4USCRUZJUVl1+AZKkLfpWgN4gg2ECteVDOxP
knvrlwIG0wsJgcHjU9w6lZPsXAB6Je4yr/18IliFufGxp/6zugbMQkU7BtaY
oJ9ob/ZCaoTitBcaS+CyMS0b2AzGSbvZblSC5ZXOCfAs3Z+FDC9Mtzl5137q
3JlpmIEgfg3I00Ac5/CopZ87gtaoqfOFJmD9AgNH4e8aNS5iZBuLHISi4mer
cHC/SRybNCpqStf2vBDBxsr6k0597YQhO1TvJIkYSehbXVi+AheYX4nH+SbE
8yOACTjIe0sbLv2mdUBGBPbqClp6Wa1Gtpf6EKsGYD5Uzvc1SF1/ElL0r2sP
vJVEmrKzobfaABNxZKo4BwpwGFWLuBzy0HnHWW9xMXDnaD1mcCenhS5cGP56
KCPY1fv4e7287CLF1uKGnJ0Qrc3eUcm6BfRG1yoiCrm9AqlYrffaBFvwjwBO
U2j68m1xJfClXGwEVoG79hftx+pHvPegiao9+K0kh0ZCN3Jo2bIiERBNqvEF
UuCkL4oyE6XK/k7fxws7ZOqaCUaUbN2zUaJQD//GBP/HBq0Tv+2izOH24QEr
0tL5FE0/80AVOe+HJaNj0qJwRkpo7OWPk4A6/ItmCwc19W6eETJ+4kaMPr5D
x5hxYE/bOo81aGtQjoF433ILsB3aH+67zwZdiH3SmBDzK016NNt5aWZ7DqG/
Ud1OPufKg60Ob+oTammpnVU+flkJSzX7cuobl/GSTh2hdoV9ykEaMsF0sZaC
prWMzxr5uEIj5U4bwFpDwQJzzImMBb3P/8C1+9NTGZ875pX2D4G3emG5p6Um
9i7u8DAqhD2l/ZwboFZ2vskAxOL1tRCEyn/KvbQi83JqOlg04w0lk9JOsVyz
dtO2psLBbMWPad0v4F7o14SbzrtY1xc/mDt2WDSRzFizONfRxra+qQ/ULl0O
rdpk7FU5DpopXtvnPoi4hM193ytgIX7TxOG66Tf0VKvru5yyKtJRJt/jQ/Fm
+D4kAenvZYJLlWfmJnVn3v7NmqKCjeVtti0Wcpiuz4JqmmKzQFVJXofLY1y2
V0w8GFklarX9Sl2L9rPXe2AGc+8HXxvfJW+rTiPhIBoskWhbjzQ/nu5/FOfc
x027lCaC4Frdo154YO/VlvbBEepspzB5w9SFLc63ZI53Z14UBQ650UdhClDW
H7JfK6pn3H3/ll3TDATtnU+RE58ap20h5Ony0rQXS80nclEiRFrDf0kGJNNt
DVgrbnkqV3YE2lj8go80diu4H1+IM93HGVsbMqeLg9F9QMkWnHvgnWO6BDoW
loDPT6i/f/NjPjXPHjMDZHjiBkFabJz93SXkqptFcFIcDttb733nxERtUHhy
y/ZZUPEqzWQWlv9xakeehCYCHximtUQYut7hqvmgU7crecN9/i+qKAy+Z+WU
GLCGGn4pIsgU7xbX6Nu1K5I6brEjziI2si3h3l6BKxgKMD11efMlXT4DXdhH
8g+iP7MijFPOfS4VVkPp4fWEMiggXmlPSoq9XymTXQ5kTHvtNPNp+Lt8lv7M
O7QDDueoE8dD2oceRVaRIbO9TZWsRvCZj3y8wCiClO9X08S/H+py6d69WO+b
MaO0kT6u42fQgHU/QuaRRCWyRuu9EqJm+b1mPnD2neaf5DHm3aKFquSs+yln
zHgnTYGe2nuOnkNJbXcgvDIIhIlh49PEH7Cqd6D1X4VI26mtyn13fpxlOBAr
pdnEI1fYZs6ML/lo7kXPErzy9YYAqknbixWHnkwwq0ohrrKe/eF9LIiAVLKW
G+sX8dpTl5mKyhwGj7mikS36dmjI60jfIFSt5tZCXwUgyeR8r33Wn9l2HBb9
MpaDtqWqzBD4Xk1Islk7e28lVKeHt6QtTD/w69ndXT2wkeFgIEoJe2iEAOyt
hT70W6qw+ehh1Ne7LFopk62280n19hSkElDzKb1JuiRhCb8VAhSorUl+DAzZ
/8wXzXV0DnPosaDyIHp/46roGZGVIjF3Sv9Zt+8jo/6Y/P35AE498HNV17yk
Bx7Dc5IVtIfflw5KqqtdzzhTDqT2RD1b6WEvr4uKiZM/3OJox4ljJ5PiPBw9
Kefcb64ojAhYFuJZFHG0hoX/YIO/BavjLWZkyaV5NUCx/XnYISLxG/xszEhg
1qSPXHYGxZWFIp8BJ4zgSe99Ta3OnySlvvRYMKzAhjg7mwjSTaONfPezD2YX
4b25J/B/zxD8w9MZWZt9Nzw2Sxe8AjKh/3GtFqvoewBIiOMtYrUdFFxXpNTF
Pafl2u2Lvr6ocSyndLo/G+fLq/bB6chJTezV+6OIHH1EIUDTZrAyg0YZQvMa
I+pr+780nZ9ZupESVs1YArXqFyZPEI7ZZ/RnIsNIO3p7pMHRUafSnjNA6ABG
00Aw7vFYyg5TVT8/EC039GsX4RKUJfQdNcv8qZjrUg1EqSVlLvcSp+z5BY4a
K/eVAlnO1V1XDV4ItFPy1jAkdenL/OyLNiAKpd9ojHzhMHp40QueNljw+Yur
1yQvELmS4QHXTU+6zDrF0vj7hFQPAiCg4iZD89+1dQKPcxS2GLUzeAbuB0zZ
RrbPtrZoCmtiztoJCNy5EG923Q6gndFDOWI6uzC3qNAQ/q4ELu4pxlsLrM2I
FnC0vmDJKGEPYpqq1EP7E5PL5zSD2CktOgMnxYw2e1BMOdZlnxVkXLLgHsjK
IU4P823FrtY0HB2+HKOk49fO2Du6Y4gxLoittwddznPXoXSyadFmwLTW5RhQ
TYOxVnI9HX0VoBgoVzPqdlzBNrpBdI0zBuQHdAAxKFNnmbniOcI2UGXXP+BR
IX1gF0g9gxEtBNXqDdGaQZ9aexwIVZD7XXMRaDzf75VKaMX1iLFXkS6l6303
pMETmsDefv9AOyjBc/TyOvC0y9yCBq0aiYFNEkPk7SDPofaGnmdQA8NuJkSM
9/8H1yEFJoWJLlawPgEC/X/jv9pp/2TkJPUAa4t/WeC3OACF8t9rgPaSNbZJ
Fidm5RtZ8QFfvInyHfnOGICx+g1ocD8x7ICJ/Eka/91bQzWS6mZTc0y8JkRM
UZXJJY3XGC1eQg1OBNwua6IOKJuUqcrNmYDpvv+pyZmQfSdvkdWJI8IntW8l
NUN6ErF5wcNK3PVm+6hOHn2165fZ1c18lxtmtdLsNi7L5brijcMF7lFvM6nE
FGQI17vJVT+gb2p7ruRdvvIqKgzbXtHZ9MSZvlwKNngT450nRMUeAICHw9m8
/oD9GLn9Ew8Wlim9gaTeNCOUzMkFrpp91RT6S4N9tX0YtXJAsScWuuRv1S+Z
k6fPPx6p+urUAklLkJpsVvu78TRQY5Nlh0ThpobRin3X5D0CkAAQr6+3o4mG
x6ee8qp1ro0x3eWaR0ETsHvRwAwNR4gqmkfSbn9IgPD4dClvyRTrMs8OfG50
lS1wBqV8JYDkrxr+LBfrJt6mwdp7/Q6F4I/eYM2ppQZR4Mm97QFDupFIMbWv
82LbMaRphFuobwGqIKMRhXhBM57OmuxshWHN50iUTsHeq8wfqP+p1FNPKCAs
wjJzsLHUmJUGvYlkkpnc+2lW38u1194f21YdrqG27KQVmoX2ua6Jp9CsgvL+
ozxft1YGVFBgUxFJcI4hlcpiNu9F3wPSLTNTk0mw2SH4ABpD6DML0O70NKYo
UJoPBdmdW47KI+Lqv4jb9bemu5tXKlPRVth0eWTvfMVj6jqE1JaLPEjtK9jL
qjWt1C16AYPYW748f1cK49hm8yYWy5/23tyIuitZi6s5NEuPofHpnJIuRg9z
V2nZmBea1LVanqqBH6BcfOIryQbpMXQrMsXxKlpCK8ZtnB+oY9EU8TR+NW4G
APlBBbRkGL0wGwVlsu1t9TQMxOGOMiCbjwgOkBbPvcdfX4FVPOq2SU7J0Ztx
oVK/6BzDU+7VmHg2BAbqaYYWtC3wyDEzBXHy1Asg7QAkMAeQacAB/Bp7xa1z
txzfssH+lrINOCnG2kBYTjepsrjjfy5GSpQC2AQr2RZJV7zEpwj5Ud1jGp58
2jn8ljHFUTwfcsCT6qxBunL2BythtFiuBtV7WIPyaEeT3VR8GH+9nBAeU7B4
xku4eRzSUZcde1YQy/eBZ53tJcjYVqNXVVUqiSXF6dolkwsKsLgz3ORgF8E9
dEhQ58qih61oo/3kM6gUOnNBu5DT1xYCWvlKlADZYZZZGHo2wj8kIU8kxbLr
Fb1sVbF0ABwf/ELclmOrMmzOaHlBR2IaxQVvx8Jyjd7XLkMbQhOZ4q6RoiHG
e2t4f/FN8f5co3uAiv81hApF0PcSbPYed6Np9R0oCMAIvTMb8SSvWxDORh5q
hE42eWHPwfB2LGBXXdGurlGMYegfjuEhRT3fzMyIn/LGBqnTB0Vl9TRKenZG
Zi8Etv3fca1qAAH1lAJ0sMhxBeyQYx2bLej4Cm92kHx+RXHL8ROCyMqfrCMM
HdEh/7T9Xt2Pydgt7eTBT7wHTsG/aYAnAJgXGA7sY1H4pfl748gR5tPG/tVw
TzZ9BfNTQKecVTS4puOlM/zGu9Oan4QqBpcR5VL10rn2xGCDhvOTa72sAIIi
ccRO4+2vjntXEkitb1kK8yeDaNYrTnFJOFU1xlK8kL/ogBXFoPQYxPoImtRa
EEWYroqC8IJnq0bgmMnAZPr8NziLsdvYTSC4KQGk+lbtf316GLclTHByI0jA
ZbvuhnSNgwKKLPNhHIey0+RGLzKNpx7AvnSvA7m5N1SgCOjjNBtK/FwHocqJ
6+HGXhaO4jI5Y3YJbh3sX2kl2oSuOJsCqsFVEIwsHOjzhrgObDaHLx8pdPmK
++b3aGlUo5DoN1tTYVqxDqJ9rFamigSIujciCozi/130dD93MtdaF3rotlMY
lawgbQPJwgI0MKIkeodwS4uwsez5kbD+3VuYSEiy05fFhR8VbzcqejxuiOuE
DclAil5mlilA56NWqK7ZY3N201Bwae9BIdF4NvYmJb1Uf3SozgceEmcQuYbS
KFtpsOTBmbVGfbFqT2245F8SPWGWjf3eVedu35AAYk7/Xgm89a3gr7IifZxX
9J7NOKYk3zr8G0Cgu+Rs+4VNcOMjVmsDxN9eLCUXNLdOqGz9N5xf2AfXyytf
d2n726FlhnpKhJS/nurRNlZZKTFr4uaFro1y1mFTRLXd3BS23l6UlKTX/QPC
e7QxP9c9wjAJqwCMNRYa4FKpzEGOO4vZlGSVa7D/htvE4jRfsMt1qzzlY1WU
tYyc1TOHKot/a6I6He26GUPLyZcw2Nz5Pk/6jMAKxS957bbQQgS0iysNxoBQ
W9QNyU/NPgZb57i/KgJuQumYLySI61O44UpxhJioEmjqTTJez3X9YPH/3u/L
nOKZvFjDF61+rlB6pneVKMGuVDyFpWUMIRMtDGdv1825G5utjvn5qS/fByxY
01uh1kyehTag1eG74XJB1JhLz+TrkSSmOE9bvsA270NIBXofWhyEBmiczElR
VevEYEhIbsilMxtbzlKLeCMggDzS6S/F1dmTomMQbJRpe2T/oVl1BrVeuevs
I8hHsMoQE75svR1zQEC0fgJ0i+EL0ppn1bZDR4YMEQ+tQ9oO17JVFnQRr4aF
mASriJZ2pmyM0mEnSF6k6GI8t1f0icoi+O3IfenmaV/pJE6RdEJH4XHo75yZ
cKwvA+6zD5tr9L9SKt5MSbCgj4RguwOBrYwYAkO1GcbNp7x9TtrJ12pA0pyl
SJZ9LQDjxg6LJfjceWd0JFSUBPAuTCGhCFzgH8qzQlDZLDsNkr3ajXjbgPcL
YueXW9y1RUFu4YM2BV4GTnxuAMSGSa40dXhU9OWuxyMDe5j3ifuoACrKc3FN
/rytc9rUsWOUfELIeyJONBgTzgNApOaRfafTSfIkoBVXK7o+wPZELRgO6hUh
udSnPMBn/L84murQRuYuNsQr8IHZ4m5ry08+m6NdgwKjxSGxrnsu+NXfVC4P
s/NWGZ3xfni66mSS9JAKO9OU59b4K762ljaNaP13/faIB77v9NXlmSDUQMB5
yYz8EBUx7Vj7wUTUqx5eZDodJ01vuEBBtAKb4suas7aXf1UYOxIfUj4Q9dPS
aJGZVahTBIuFVk2HQPwEfjXmumwVL0e5KaXphopItju1YRYuBaaf1pabxHd7
/ZHXuDogmyHPdHuveRBaXTjDwC5evPEScSz2/PHM/tVXymyoztnd2+vfraJY
PhaXxYJCEaE5Koe27H/2/hLDbR8gS7PmydnR1UjkMs7vyoeKkUYvnq854aGd
OB7VJsB9JnFlkFwFrVCf0YmcN+Z8OU1GoSJoSxH3W5zPRI22Ku5/FnUSY1l4
KNnppPwnGiV5cdrwTyxeRFIxg+HzWlwfaacL2nEqKGGuWoZysr8Wwhabfg3x
y+0ifedoOZX6D8fxfYD0Ziq0nDW0hblwMrcyD++b+pkxbI6jHHd62BgdTOar
79tGhqYIDOelwFv5TcdIkmGsXR/XEBOHSuP/ZMvS2KyHtgcoI2PjwXxcY2xi
hl9tMN/1KeFEHS1S4pthODIzKJmKTreZgRaGoElhNqgCi1NLVHLoLCIeSODT
3AEJW2Feu/ViDBKQczT82mfJXIyzFz3pYTuBtACpUcXN6uP3q5rU6JWFtkwp
658Rj2g9rM4OqgkVvnbVMMTR1YUoaE/nlKW1v0Efun0PNOwFYWbUzPacgzzl
WfEF7iBt8XpB7Z46dro3UToVH3jhacLNjTJ8l8NueS+Cn6e99Zm8rro74asn
Mu90Enq/81RjpsoJO7mHzh+WjiH1insRfLjNgK5zvUGxGqT8QIeGDHYFaCbq
2ml2q0Mo4RnSHS47W79QhoK77duab0aGaQzbGd8FBGoFIKEFEJj81UCl3Uzx
9CdwVNXMohM2gtCjidkIdS92oa6owmPH4O0pswYKzOEVV1tv97BJwvHb4rzx
KdPlaVDUOrpNJ6cLcVsP4O0O9/x/T/2PO9+cidEjz0cL7YrmF8efObTGCswv
KhSq5f2d3uRz6x0tPrgb3WF0VXr3jw2dMO6FVQVWxsmLgwebR9sA8rPHrQqY
cFg3GVejWuxs30mLyJYQlea2bCYdnEoO3YfV2df4ToEZomKjqwAVxBbhgzha
2it42aFbVcapcdr1r1d5R86S08hzVudNZ+YjYs4Ic8NYhcKv6h/eir4xoqFd
3uTI6MeYZXDqMnrJecwyb5r7nPObvH1C71x8z+RMBz0+9+G0L3eGbN9fV8Ot
Y+Qg9yLlrQzKrnzIXv/CnIq3wZFi/9rFsQV1ai0TbdMQs/Db8232AhDwQZYy
dqgt/apQlxRZ8p00txrOIiTdoQ5kQ9zCR93+fjOz+M+slp9qgBs3m4BTzPfG
5LuYN5RG5t/7K32tozGhP3OB9MSgSIl5pvPbtj5issFaJRXPDiU253ADFhks
u52FWyYMEGO7WFxm9zAooRmv4o0nvYH1Kmh7unAqAU6xVOtvWHAfyWRNSKMu
j0lNh2SGEuu+HHOBWr2ZfpacNeUnuk9+0MCulFAQN+dqT9/jAAmDhVXSbBma
sDRsOxYkjvoQ9DRNEyPHaSLiqhjPRI5myqIUOpuZC7kc8RfBRs/fWKYPh47n
Z7LMnOPd0dxAYkxXIrQMNSDIa/q+K0UrS0V7cROChe+PygXBEP00A8BJElPM
4AZxBCKW2eNjJX1RaKiQZQZNs7TXUZubAFnAM/7Q2hV4Woc9xr5ayYG6dfOR
mEb0Dr1xeRLRz7B98/tC1R8STlhK8W9SILqo6J437ltjwq8fEs0Q82hEfbX+
+QO2cKaPXM9jlLqpVmn7MnF44F1EMjx6S5OLqjlddb+U7AXGFmzCgGUu+LDr
3BQx13AZ2xW56SmefvIpQ7yjH0fYLPPL0DJpsfDKT6aZR49bP29BBZZ8tNz0
WmeeE+pEb4NU4qJHyZX3lgI7hRtx9N8Azc6LHA/C4/KpPDiPxsOYzTUN9cx4
E/g9bUGPx/6tZqD5n48OgUVQI1RTbSHJxTctCfl3unuRJQwuKGd5Yj16NSKk
gIY0A+cOlJXWVTEMMa1hdRKh/m0MowU+h/FbrgAr8HWCOmRysMormQWArvKE
cFXJgV9Ge4T49TXJ9pYY4WNcTnDuVsKHCTGDwJhHKz1BqSY50EfPoA+BCfrC
ojtqDxZixwdcPYaZR9/n+kuCqwmyVjzs30u3FbtTywXmnJfrHKKew0ins4mq
dwfqAQ1AMa1rUyLOXWrod1UObBIOUkAMsGXSNnItrLCjyCPBsB4rPHXDrw+V
gwSMTuRQS065bYLp+g7uVnTV/Da4yAT4g7v5Rp8e6C0qbRzj+p2uq8Uel6Yw
UD4Sef2rJFdhHBgZgpClB5OeduPw71UqeXyWgqQv2RESkpZC4fPWMSw3wHxU
2uD+ySLD5FhXD9sUmWFwxyT+MaQ55KNAkZHF4Xyw1gjMB51lPVxndqxQ8v51
tX1TgqKKY/SQSry7QT21IO6PS0UMRCmlievxxGjltfLYmqGVgoQkcmL8JeT8
jZAu0LpwhSt25qg70NBodybQjXX7u8bs1JvQ8qHR48Ndsf6sWrp5zb0GHk8+
wPbZloVWQNsXjWllypxVdGRYlE3ikpowg5VFr27/BGWqWb3QO8rI8GPIL67i
PbzuYlg0EhDC4VaSKZ7MLLRw8FEjjb3vMcri8pyv95ODKEmpLHLI7Cw+xa2b
T/VHrRaEwtZjmpore9zS1i4UkNW7cuXL05uaKQbb/KDwuOw6VUzpcrwkiyqN
IzjhAsz6QIjDYUj9QM1ZLTRk7lxEvISq1gu2BLAU0QcKWLTU7kNIGycK5QsO
fKFzLq9ku47Y7VOnJ7GtiWAnS6TTZPtHMVJLvejwzYvD/d5Q9f1s/QxabF/x
q1sj911BgXQqXo4Ha0D4r/0R5BzoCMSgClkaU0O+LpQQTr+7VotDEs7+uQsK
gC4ygyjOVuDZgo59TJz2UX4Pd47tJaRdDvS9qhzmf8SxWGC1dIbUqQrBs/y3
R15tXNXUgRtjNcvtMRd9l7P8+8bcqFzPqeefzwlxcZ0vvld/zNzWgw3Bvuke
kkRikhKxjNABQmhLQIhz4BBCOn0E/SWfMNUCmWkInzcey9b4/Afd+/S3bstY
JeW+Q2oRr4rX9RQ5oWSYM44CkyRNdqRDhMvq/WckBsYOVFBVxtSHOHF2hXV2
VXxYaEG32wnTi/dbYnXBkFJY8xLMPLqNobtnS7LDDYdyrDwZHVBWiRj7iyb0
a83atBlV70UJnj1mYRAWbSPv8uEhO3dVTieSNd20WpzdkQp6POO6WQjc4NQz
7sW/GNKXPXV9xUzjOyMporqXYuEOyXE8WYpAvYvDne5vGR2iw2MAW+XpGeOA
cTlVH4Dx/3N8lVlku1lCW0lx+yKSDzKg4AGGf6L0bY0iprpVnejUOpCRh9z7
KgnEi4M/7+v5d5AANNBgj5SDKHBcDsZvltYbovyqGZIYEN+CfV3cgyJD3lko
tEQGFGsa4lNxNZKMlcnW05Ozg4bnMKS8ltHZzWB3ffQ6kqJgrkLKBieBwSi7
6d+1LCpoqaqKF6jDNzmMRVjNjX21mGikv/nLFvYf8czSxrbiX3VMNkCjmRbR
UmVxhZVopns/iUWXOuwQC49px7WcsJG65zYhPbCadxzFpVMWpyMxNZbXZY3E
s2vr8Bc+JEEoPiiHpUb3KrC2evOkMwZ0Rw1r/yIZK20OQtKI8Ad25lMTMIFl
vPNnQoWJ75BqXTF3WPu6mHi02O0b5HK8Nw3gfli7LlZOgbT5+MSt3xTxwlp7
pXNIZ1KI4FlQ8ck5OYAhDvJfRkjt21wE2m0CKbMKPo26/Lhp+diq1qLBjaqg
78qGDnhjoo2OE/O5WJQ4qOAdgdMDIlXGdiPvTXcby/Khyv98qc7PGjflU7fE
Rkt0+WTrgZFE/VY1h/48VlBi98rAt2+RiqRdwAl1tyqvmrNSkMEByYivD+N3
OI4FQADI6AwF55NCsmFOuh5xc5nz9gBMa7XjOlo8Efj3hPqD7oT3dRGKk7YS
L/qj5gq4Cnnl2/5J2LAGZ2yM8qTPqzuWM2Yrh6cqJj89fUrKGrWdRMPKDm15
0xLBDh6N5FhFpMWw2Ut0xWjJZPVdFYCxaur5LO9ljQS6AaJEA+RAXGEfoAy7
7f6C8+n2jjeTbiAgQw1tpjG5eQeRj9mwPfAbGNKyO1u1IX8Ws49y7xed+cSH
+rNAk1f6y5RIWaoOP5ZjZAYQ2lXkaN60zOeBtqfnnzRwsppiUhQ4VzKGdvR/
p2ngUzgydNKUZ7dzSCwdtaucGFzYemuEEu2nI5dvlet+SPDp14r+aaHgFSWA
ZSj0HnJpkvpHbOkw0iYO1eFm5dkVAGwpEr243Xslj6C+c+/jJRPqBUkDqr45
8epLpyBgbaQTC8trnkKBI6ja/TlbMoDn4BGQ0MBSQsYqfnNiUXhXzNO7j2yV
UtHVwD+Ubbgkc5/Gukcl6d0fyKY7QS7YwtyoihJv+VVHcGAmmrD0tzSgnb1x
lfF2EjbHxvkao8INqyJS4mGd7MsXF861WHIOxf0koYqCTkVn1eb4c/Kl0om+
cvKAj+IH1yHM6qsTQI5vb0OB2pkeb9ge3h0MpDeWDCv1NFQAJkkawX2mHdyK
iVriQ3qpW+jn1/iKjRK8XR/YqlabOeE4xMqr4+PSqWLvS2gMSq0HH9D29rzb
12IvimlBvh34ei/Czp4vevbYoQxHwhj4X5b+qYS7/8B5J5YIb5x5w2cHQ/TY
LLjRqqJCANh0N/QNrhRhzAhC4fqoyYWVb6PZHo607v7DASFEE2cR4VP8sM40
hWo1zKkGCdhC2OtjgsntiZ4bdMqdzgWiVeql2oGWAn7yRIDugX8i2p6/fX1N
hzboGpdjMLnAhXw6CocSYrFDbRQFLs9OyEje3qMQno/nRBt/8fCTlI5Y0uyi
AUGlZKuwsmS5L6sYTLKMc0ddU24Bs9XSdVhw9iLUyko/q24deactIvcjUeDV
K4yXkAA7lD3ZIFGqctJ/CA2VVQWuj6k3ER/64gNMvbAl67cjCw51fw4fIV1z
t4cU6jAgHEPTjE8EBLxB2izOt/NaHmc015pZEzqxchvPqdB2juXqdP9PGyws
7i2fze6e3Jt325vfPFDeIRYd9AIySGJmR+OWJZgPg0jXcqSvL5CLJM/gIMOX
kpwvXhQ/yON6dqp6wDppKRG+wYUTuxMzE8vEQi3jtkhT4ybzjbSJiVcEnpJ0
Ct2LLijO8pPb3VxDJ9ula5DfEPtkHG2NM//DdgdbZdzV8wpsBqgGzrAZWOLC
ISgqeNPL+f9muOgbMZy/Ez2epK/foTr8Pni7TvCeYRoHDbOEL4j/rddUAQ4l
cJR6qcLPDBTCyNrJAFtw9XgHpJ1Ft+oyst572Pv4354ANTGeH6+wgBBSFCTT
mlpJXshlGxCsVqeEzxTeF4M999RVJOr1N5VTcrFZOFF5Tl0nfNcR+rz8hBvx
0K+y/zgg9VWiLojqvXCKVK/zjl/W+cHjdDlGFsnwR3xHH+gLNdiyppa3lETA
PUWzZFFwlBe1vo/7l99kq37nyCJmCQmfLrZIdx/RkDyY/cD0tBSWlD4DqeJ8
/oehqvzQ78rAkihyEsR/uOSEJ8HAqrAEy+Vc9xpC6AAv7IJJ3kEGAFnF7rZ6
dF4AzSJoQLSAnPjjy/RoJxUtWJJuXEcLvww28gZ1BjjtWpgMTGz1YKdBYd3w
56CmhqF1HLZUcEb7J4ujGkCk62am3qG+0fZXb6fffzvXJT31TeyiOUxoBVg4
SPGu5kJAZXpTzfkWWpGvQLz2yhOz9BQg5HECpuD9llfNNsgjOPnSBdSNbNWc
+Wanm6/wfH8puKxxom6OGmSHVxDnq2Yr3peWA9hvMC+34eZASCDMZ1zgYyVA
LzztkiqzFFmYf7KAgeiUqPVebctkhTEbBgN12uSctO1ZsTY+AkEI8JfpL8jT
3MhD9/ZgHBTRetfHbmpWnJwIKcEw/osNBjU6NKkd3pe1qLAo95Qt5ckInUF6
U7wGwLVcPB/UtbSwHTOBJ38JBMb90U5nUqRp+X/54w1PacIqLsqTmB7JmdDb
AEhSY8Iu8EEJlxaUcImjxsSvyv6QkK9VzUDCzJDun2Q/RgJBD8cytAhmIjXK
7Bup3dqqNpYmVn4TWKKGUdyTLo0/+vUa7eKQm90Tc4EAi8cm/3TdTvLf9D/q
QWRghTdpx7ja+1OJIBKBXwGL8+IzuGiTJXkcRy+YIs7Y6AlVKdSiogGVzJ8L
+IVXJgircrTk8iPoC+F8EHklcCWHp8eGCXN6dMSBq2QoPBh2KgQYjxTjnMbu
Ro4kj1d6Bx0/dDttSSbWoPMchOWcG9EinSBhMQa/BnNJfrTuhLBR/kD8iP9B
N0Wf7EEkxad8THWzzq70LmoYJhV4gvbzuZ0rtUEe3Yy9k33NmJ8CvQPWTLx4
yQO91fHoBi8hUW62aH25zN4diGOdorfFbqaK6VO7kuwzS190XZPTTzqeG2XI
4FUdmVKbtIIkdlotNCRqDELa/qGsjh4OnWEws2K4AgC0t/elU+uhTrbNWnMM
RErF0tOSeNz+V4znv/F0s+b91szXE2RNWZKzF8JIc0xKbkyXNJjyI1UT4k+g
LXNGy/B3xLO+fdF1GM12FOigAf7fmzhHEcHYUf5sPopKeITH9/ibcxJfk+sM
ujss5PwZpQjBLOW2imebFTb7/m7Ppmq8fV/X3hWmVB/C5PDhGbuoe6vmt/YH
RR8fvLhkUvFMOdO2CEKegoLUeGRE1UVmuQHEyKdLXZvtoJ8GuFFxpb8MoK0H
KtLk+0Bg2TpYVPfMVNuSshhYhrE0lBPQDJ4t/UiFNB8+3vY0Xstv2cpvCsur
7zn6UZRDw5+MC38TmDqz6Bgh/P60AiGnO2A1QgAFAMqnuZaJjdZte9uADZu7
pVLIGTWn47y/7sJr66G0X8a9KnWpOPZum8oZXvfZowPObvygUd9tXP3/twUC
YW+LtwIdhrCosx11qE+fYCEW/dItmlcbcsfHskDhFsEtEuz5id73p8qzeRo4
KzUhDF54lJOuClH/gg/nu1XaR/vZEmCQoHlcRHKf6lqf/1JEcQSIvR/UuuoD
7OwxQkRZRC4uaETo6NHooSaIe/gw1de8F6sC65yUc8T5I1Spdy1iHvRlvZfU
YbU+IDUPdj67jYnn4NZPNCcrisJKIr5wyK5xASdaqrUme9ImBvVbgWpEOFJq
wyOt/h4HHGMyq3adispLJaMExopjeHuW9TXFdHVISoUfCtYXlk9TBw13kbld
MUw9ygtbo4fjSwEe6x27Xqp5sLtRrP4PjfnTleW1S2j898b4mHwMJR3on8VE
Gx0UJ3hkol/urnVtaC/asXOdKCSzCBMyFTENdF1R9LihDG/xSh7UJSYcVLkY
qL3IceKcWBdBMg6/yimkuECtWSq9KnwiwjGXRw3eaiP1Pm45wfY8BcLjTTVZ
v0BN1QkTow1oDNcQKAVjo9/eLE3xAaZSSU88ZKCmgMLhS+ujHCKnY1sOukZ5
F9mJu074aoUf6+x3oNdOkA3vdXoP1TW5WFYN7x/Jf8l3ur17GCAUGdlDPrGI
AfYb/1Qq4T3cqqxQK+Q33manE8iBMtqL8aBXLJD6onZa3WNb0N86HYN6FjfA
4ca/2SahSCb/8In6V4N019+/+GmgTR5hDqpTplqLdS67MjjkghGc1v14xpTJ
+z89KcZDza0u5rf6YwbEUCCyU/qtaq1UA6q9IFk1XF2kNpoHa7CytNQtNxqN
yXBfcSCYG+eKhZ5p388i4OyYTYK7oToG8MD3d6uL7Yprc0MlZAaovkfOUa3U
cOLdJPqzM6nHDLlTgG8JEHggSl9Y3SqwdaF2ZbvsPJSC/FeSTL7cY4Ye/G58
gsbI+VPG6xBbR6Nrm0FziOW2+99WUgybG+ixybJ02e28EqgflgGrTmMtcsGP
elXelWRxV5Bf4t1+JWqLUB9mD2jULYASeO9s1AuLPcXj+avN3pyTkD0qUdyR
vaa9Igz843ZEVZ/AjoOAvvvew3XxKvHv49U2NNkjQEd+qeuDkAuHw0h7zCfR
nGM6qNEfyPZDA3nFfUpQ3ORHrPd6DnGKzwwZi4xDlRp01KAezyahNlffCvIZ
z1UXyvB0TJjAZa5Yg4QNevUbs4EwvPmcCRJD9MSdC2dCYJPEWyXik7HTpyR6
16GJs2X7KQGDb8L6RWZoBmS5FvQT9Pt6JuUESL7l49pXwJIhAz3yg/pId07x
2hw1SPnzjbT4SCd10Oal0B9sQIMTo1E7gIa56MSVgFK34EUeeV6tuDirPzkX
x7KjyZVv1/sC49JoCCowRPjQV2EIvZO0LZzgQfC+xKp3c/w284Xw4Yxezk7C
qRTllQlQTmQ9l50goaz8OBhoFjR/Xny+JdcUeCDhOcI2MjP+64x8DXfRvnfe
kh5ymaZBxF+qk4FsJXjTZO047/hYGVNqukTDC2rTHGelj6E6seaIasTtmsfW
SExGlUoy5h1osx33kaOZhavZ/fuuAXPVHo4m4P3a7/9e6GtAlvy+piewpCkn
psnh8IssosatNvtucBzGxQtMplud7eQPdIfptGPsOVJQZQOvlJ5rj6fubgDa
h6seSkh+ailH9rmEAk1ypo3P0HPboZInXYZiok7Oz6x28aJfjp7+YpnHes/4
G6S2l1aBmrx+ISkbW0fWf7auN8A86N3Q+DF5uOwfebpSZumdNprDMZEkm8Ht
89BodbQYBrayi7RzDoJFhddQ43nVyPqhm87jRIr0Z3AaxpoAM8rp2P9QrayR
QWf5gAcBmR5vraXt1aNc7MfRDdJHw/oTmaScatZbvmgGlQOLKP2g9f3R2DB+
9m71AwlPUsGgiuT3/MRG6FeRsHx9XXtCwkCNwckYHGaynXnqKvHcxnCgBbIl
mlBXe2i+p4CnVtkHJB0cxLouoImbqZKcBGdiL/gKvdR1GebP/b4ReIUbWX7k
cnlTNHxuWr9LCjefYsmBoq22/zsQ+70QuXxgfDzY9hYYfUMO3YNBl/fTgS49
dCKj8CMXXYmitGfMk2TKHJgu5Jn8sMo1PGRfBrTBs0mLnX7xB3OlRWZI5TXg
Qd+j3M9HhAudWGnrPpGy/JddLS8JR2uXH4715I6lYYUapOaJEiryZS98eAEH
tQEIqsjMvXt39NmYvoJjl63kYku81S4dOQKDRNLZ47Fk4kxV04T4csc5yy6z
0+iWtz/Zkl1/dHklgEbsLVzVE2VYjWfrDD310KCrXWUZDAAVWDApE1kzzQE2
ziOUU7wtBf9Bau+m9eXhwWcowrDahMOh493+tf1qwALHmN8NjjAWt6Y+ri54
GBe7YF6LaMWujCYHLnooZUpH3ivHCe26LEQFBf43tRAyUb21f6ren2YVOEtC
IAkVGJJgWJSmruk5JL/jqh9h+q/l7JfOMOpSl7/NwFiKGaD1War2q6d30c2s
/MZ70OBFwJUI3JZ4Dwc8iXqnr+6X9GPOpSbdw7MSFJecKyK3tRmIYwyu15Tf
NjTG8C9F890gabGGGOJd3wJkO+p7whs0wvg8WxCGLbZRtziRzsuWY2D7ybap
ityoP1eLcrL8zgYfZltYMGzP6bev2rurGaaj9tdmjC+YwApkVCKPu12Ve7/f
Po+AY+BaEu2rirLGaW+SvhCmXtvvnf7xKDzGtalXuTi165juEH6sbmyERUsV
E5zoPq13ip6+xV00A3pQXBp4/eNp5rZzTVgJ2IuNPE5qhTW0MOeGdVtp7VN4
uCgdYpMUKZtiO1iqIIDTsCsxA8dCr22ZG4RkNx+TbgJUfZrwrVgLpYiil+vl
QI3RooFe1FBBNegyRH7CE7V0uBEMC8mFF+xNsFR8Y9YeH81h59OkP/u6OipD
b1fLry7tAwmokwcV44+rR31cBuxZoRGRLuPCKjICPCdkvfW/qtn7svwt/cvf
nHLIwLKv76AJEUUpC8WcyGRkxgCfLeGcRRiqu3/UlwScXRR4w+63ejAhZNcT
qLv7LnXaawbu52Yr2yBtmtfXQTtsLbJn6hKwsVJcyae0T/h2igUGXfnHXQ1V
vbOAUuGn7Me3TiLmYtEs2NFUyLqlHoHNIMjX2sMXYDWrazHyUYWxz8s41LYY
LnR3T/Kpts+MpOLIm+baD7uSbXCcKj/5OfyF6BzoBJYZ3pbgXc1niqC9x/KR
LYacB9eVUmMZPF/XXaH50+24jl6pq48z8Y9RyyHT13KmoabzqO8YLAO8u5Wg
1vjZNoqIk2Rmh9GME4+uQ5x1wmZ8wtTWJu9lNZvdz6IbUw/PmbFXKvO0D+pq
ptp4ZnNS1wMsK+SRym5lBBgogjTtk/CNzdMImAOZj4pDJv2C0M1zWs+q0hr/
jteBBr98DNvNvDHtMYPCVva9uoKPiaZQrKbzPWz6NBWjuqEUraT3PpfjWEYY
2Ce2oCWjxOBzqc791FgL/JT8FzVBYx2qyJ+wfTJutBPtSkLDvO/LhWBPAA7q
9Fn+V7L1+GHww3ODC9cCjq2swIN+bzYWl/uW95Hst4+N/LHgcW9nHCRrUsU4
d/nYSEh+CLtxfUzFQGVLr/D+4fvkDYGhJ6JktPVdcKbNhGUOeiLNX9hD2ZI+
dAuKt4EvncnHOSy6jyKK8jqQEGyGh5+YAsLRO96vMdBW2dHzQLTS0/Pqn3MX
ewwtmWtKyXcJf2lGWv/TeBXzQgwfraqOjMugZc4nusamfg/2FrCuwime6wNy
gi1ZIT9D3Pv+bdfUhVnhGivf2tWU9XEUL6jdLNIAmNXSKVXyu4z6lxcyzXZF
/CUroklWH35m7FyAD7obAmETtHIjgFp9ddw46dCcPJBfxTF2vwrsw5FujR7y
StFzHFFxlEo4PN48NJTUO1rePqIaPsvKsNIacdQQv48PsZrhbK/HDLjZ4/CI
VDjCiHuHRiwosmopEFyLJ1LO5/PmxL01sU05kcQH80NdI0UKsmxwGQukO0MR
8EYZDmC3Zzzx21PGfoKRWgc+S5y9OmVN8rtN9s7tcLouwEj8x0ej1gLL68oi
ylW7evGjYn3QHY0AbCjEI0s4FYzIVN3+g1X/PQPRN+XEeveOSngI81noAT5H
OQjajYf/bPmYZeH0m84tKehjHsMEKWtuXpP7SaUW8Jk604a/DFHzGrYEQX/e
uWVUqb+ZrRZ98rZOv5Bv/Kx26jPQXNeIRAPgSF6sxeqQGnISNXzMG/oSptAS
Q17yMCQ18yGYRqdYvC8OeqZTwSgnN03Is4k8X04eJ85XX3dSeupsNjYDOi88
DrTeH04F6aBNmAXrcetEPY2wXuep6kGFAWiAYo3HKqCBWfxPmm/uJqnw5VpT
f7iwNcVso+Pe+UEDA8ehktvdVshgOlgtp4sdoCvNTDQrhIxjFnvtLqSWJ9xF
tBchynQ/8rbFDEfi1UyIkg8LO6WeOz70Lpggtfd8lFYNqMSFclT4hOuKpQdo
9HSpiDRM2sqLtLw1n5xpCZQxYeaXAWxW34r2S9zOlBEHWolp11a9zoJokRUV
PlRuejEBWIi0iGRFaVPceWUaFbYjaieMHp2lLHt4E+DCKInwrMZxi4F/kten
VcuCzMayU0CSJzR4Kty+MnxYxsaAcSgJ2wX+GYivr4LqQrJYS1IzMxXje1Zl
hXZI8p6NFkD8VmGKaeZivsJUTNJFWwIEcf7Z8WFcqTcVdoNqDp7X9aOcFNiZ
IzJB+PVp7uXjJw3sn/5hspJbWdWgTg2+fF68+K1HstYZIb5rhSrz3HLNa0iL
WkhFXOCMDnd/KdJ9WjNti4UdaupG3Zp5VHS0rKY+1PZ+gUZ55R5TDtuMNLLq
j5nzFkjogsrR1tZVg68wVJ4PPlWbM09INWKzRlxCujgi6AtlPm7IxNr/md/g
vamRG1c/PWGzzNe/JqO5k4O+CSvkwQvFO7TJKsd/C+RBrV6gOZ0YeNXNeRCY
SHWbsrZOt6tslSuJC8txy7RSyT882rz6FoNvz0IipF6lOlg02ZUlP7HNCTRS
lQ7Zq9A46LP/dT6QPf2pdNfwZ4RTIQuM6FwnzdmAVtIygmrBki7baeg1Ym+h
Yhbol3L3yrYIxcMQGOEjGTBBN0GxoGajPyvkGFLVTn2VMx2vjyexfcpd1mOD
V2AvD/qY3pYqJUMd9PTEAdF4lLnuhsiAEsEKX0ET9irL5nY5oOpC+6bjBT6f
OdZ/pMbedej10s9WZYVbSblCcNVj3bksfkASl78rIIfjmL+r01BXnLcxfl7i
wdMjk1KAbo8CZU61YA9Ukv9kRJRbfLaOvqUZpJmHHvgRyXVAGrAnv2jkbrYb
GT00At48oXHPDxcrG2gjWQZjHnRv1Bu2oJmYHemPSBoDlsUyp+pLe14YIwv0
g9yK5T/HZTUYOpwHecoPLCmPfTASpz4LlkcF87YMVtIrQwxr7A9oL5EgC2Fe
zAf1CZgpSHE1B2YSKDJNuwExYiuw1NUr3i4NW2G7TA67Z61h3WjHpZtQU4xt
CtkQbaJKxPaZ5/0rqgVnS9YwQXRXbbW+9yPNqjh798qTUNoKkd4P5C3gh7eD
bDSn5UIOq7+PNhVezkfR1B9plcpACDjrITJXTh4s9AhOUcJbrzuLiE1HXdeW
6Z8mycVxSZbgCDM+u4Cc2oicXfgfft4rVrOF7B4k40JO/dRpNlT1C46chjJF
FVRIxH26PshZSR9x8pWri19VgVG0+zJZLgvDepy9K1OQnwyzrOuJ/j0KW3Hu
FDRP2dM5WezI/DNv89miAbcgswbwmUW7vF4RiaZyxmHgOtc/ixAX8/2v+59C
ES8ovMP5EWYZ8A5tcN0u727E7lVMitUKURJCRaCWLxiCaejgK26C8t9patAJ
fY2AKFw1sNXqccbnuOqfJ+389lCWyaRFefml0Ua/sk+EiiNlQTg0pum5hagX
EFfvz1VKG/7M9faoDkQKYNWdbshvMt5Fz+iBG/BvLe1IH9OO1MxIBxGCyQQU
cSWf5E9WbZ67fu68Jmvf8kqwVx6IpjXbP09suxjlY/oAJE0+k659sVQrQzxn
ywcNCkaYzgw1SuCd69AFaf2cYCyWdOJ1bkXF7x8B3m1Hdbxthp1ofnF84+2F
ml9fL8MGAwIDnxvqT6VDHgm4hH+mku/qPDE9M1uxE2JISe+CVk+HnoMi1/Ca
O1Ms8wBJrxJpA0cQ3nuF+CXSYh+sanJuq2T+qrek8W7pbdXSYroDNr+QSG0a
sLQynqHXy06kKUCc+5SBb3Uq5JD+e037Oo+NtGQx4PTdVzB8scBHE9rBYXsh
n3dAXaD0aFsj1Zi4hrWh24EyRPYsAwMBy8rFR3EN7AWO0TRweeCG1d1GEXBE
aQmCx+tVgoXhOCRvXHC546K642jyDrSGYwzkeLx5A6H1gAAtshZzqliFUgVR
0EfvPiawzHeDUvWLwbjaqvnw6+CuzGa3+dinDtGbX6rlSOsTTwNm+tWfGp0X
DiLwa2/5cWIuNhC2RQvD87aeIQIOuGPs2s2WE4xUhHsebmXwzGHsv8MSTnN/
bA7F3eb2rlHcrtoUCSmKzHA7LLsizzUcvKjIDL31caMG8XS2joCyUC3/3pvc
L3DVUCdQLOq60ozJgOreuIaC8FV+wk7x33d1M6Yxa3xnML6y1KptnxtM8C2D
JeO8Mw6BY7ZS+zvINmqLH09KR8O10R6byFu45kxONd+Q1DWbarAiIRzykVJZ
olwjYvxnBtLOIt/yjqWO2mWEggY/8xwDx2wHdWj9/fLBK4IEvdXAO54m3bhY
ldHnjSleZXyYo9hbVWcEcPYlxCUl9avEhS8yQheiYsMW6VX+iWLOekapvKCb
4VbxfqG9rvxwp3QbGiWOKupGc8qcsGMgAWsH0BrkkOFTdszCMfALZYAOUeIz
fLaPJ+A2TQqUaSOXegM85WgejDCZ9MNbBonmY1vOYC9uIpT/L6diwhnGHIOA
XunST5KSNEAQgnEmJ19RrVK+ykimFus03ZGAlZh1vGGaC0ZNt1/gh9RdFIhE
90TinkbO7tSzfdsZTvijnwXaXxQMiVWSnXdDHnhQynJqaC9/lmj5ZQAHy0OZ
8x4T4wGIXWVFeC14riCwOx3P+EB5RQ7Irqk96s5sYnhBDBSF3DvSyzaiDhT0
mjlQnMZlZs0qAWw+z6oEI1yuBVtV1xIn12BK/HFHSzpDM52VkiA2Z7HoLmxl
DebT+Si3nCdF0SzMGmfcWPyJLpnsIzVEY6XCVyeLslZzEhiqTAJAsl3tNa15
iXpmrIV2iNI7YwV4jZEf3uePuL+JoPYnr/BcvZh06J2adN1yTyvzP1sXdEa2
uQ2bnNTPapuBThPaJCOmgrWkcsQ882okPZTBdjvv98TaK/Lch3pthe7xlwZh
GCZ9AUFGdB0UhPvx6xyh8T+ELm2KjpKmEOL6PeUvmr+UtWhNnRVTpTIUuYSz
rNhQVICOAm157Pk49NQAOn1AyoGNxcrucEkVbz+/pq/u197B4mDTYUKD2dVq
1T8F6sL3hm8T0DWizkBMMfj4r1aMu3Nj9884IEim0jzb700hDsEqpvfF/ciS
coxzhRNzuMQv+HfDAVLJ3i/9wiRd6zc7IfI+JQdreI/A2U9wN1DaMNb5E3yq
vyGwG45JD+bac4tg8xb5Ro32w9lmJrXaXr5WURJdc5hArRDM0aAGHsPErGn2
RuJC5LEPoTlTjLBJcr5te+rczXcMmBHfvCPu1yVUpjclhgGHuZJyHMb9WeiX
Us5mZHvaQm0kyLW6UaQSc0OxNooZWKwdTI4RViu0Dk9sOFSc+gGPwxl7HSTx
33FXRcJmPL/ceMsC0BEO1GfNvBpK2XCyRPIjJ6nZBU6V14cVTB9UatI/qHje
x+kG6AOFqOO6v2maym/lfH1kwguZfCs5C2ReQJtI/PKAkiv9XSU6RhCIbd9u
LffTK3yl3VVkOfdUeZ8G/mMNCCQbC8AoGvcQ+DOXKFD7lTeLV/FV7MZyOuGu
MyDEW52iuMpNEFJJoh9pBjjs88VTz/tpAlgkjHvatcDivbmdoz8ypoc5TZjT
MnqvTfpY1RNSUWbrl/rQ2Pvw4Il+aI9Y4NfPpRnDLt7nWdtxRcW9DHXmG+UZ
bQo3veHJTv0kk1xaqUWV3+yZO7rtMkd5kq8QGD5btjMBLbDTEMUazjwY3FSN
vOfwVwD82AiZGciPGGW3vzeXoHStpv3y6mQ7ygfbPKXBzZiCQIvF/ABP2Ol+
x1vSdZQ0xC9iPZ5VEr+/uDEVRb/ZpDaE9wcSCbNgHfn6qJRvqNXYzPAjsQI4
U5ZhttYiBojxBER6A688sM7+5CZ1maBXujgvSDetwKp1WkjjdxWenW+w8vb6
sI33TViif7E1BoesR8E70SyHrUqs9DyL7B0P61uILFU8EWX4dY8+YyP0Z/Sh
s4HyJx77ABAc/G2xFvXJIftWv+/qCjyLJY2ZMLvI3a+MGqM6kHjVh7NKYwTS
tCE1S1Q7fCqlyIsAtGFr5EMUHUtTrVLn0J9t0RS18mD4I8hFh0v+giK37oPc
6BiZ1C+jTtL8S+oXtJeGBRsxTunK19ATEM/3udzeBEh+AxSWQYWMTFgGrd/U
U/+LgtGvX2ObbAXWuofgxncwMUdDGnS2U3d23xnkN632gq3vopFW4cDAhIQv
RNyLc11m4mb94VJi/tVeErtxms6wEZScLd5E5Xv02olyR7po/3k6ILD5EBnQ
BO7tOCpECatEHHCKFVRxrWtDTd2svdgX7xs3fCbrpm//jANvYRJCiiVg7oky
mWVyf/QecrvFfu1dNPDyXckw/6a+XhZQtJO1NndwP96YcQ21IxM/oHg0429T
1e46vIR+o7ab3rutJYkG6ypW+TNI+Ky7SkjpJ3nfur/aN0sVJ/bIamBzEkgG
P/PTIzwaBrUw7oAxlh+5u69KDkMe86on5vn6A6jPjlTDP1LyaA8ywoh2QyWV
jivHRn9CwQGpLQHMasLpEcWeYJ5wg5gZs5LhPKULA3xTwSoWcoyCv4yvH+J0
0yM1fAbh2ewI5Njq8ups2Wskf494ZODqStcMiKJChjS/pF0F9OPEMjHVrnxP
SoVdgLNh7XoT4LN1zgigRlAVOJhfqfLHLQYRxjPx1LiOdaujgY2wC2PkVMIM
Upjb0bYZKrOAZnT+VWvdWcm35RAVV/hpIDSRw/YYeCJi7QQhaD6npzlfwqEk
71tjOiDsGxkqHbhn6jqURPvSgJxoSYTtcjVOkEYpp75j3nu8IkVOxkxb6sFG
ln4pPw1QHzdBbHO1RHWkU3xwxZ7jFrI37+tAgcepcowHiO4leYlPMMGChpbp
uXt+vmzn/leECrAj5n/5N7SxBZ4yINJ3iRUzVzF1M0lu1vIW4pr0SN2ooDwK
i/vNf1GG0e6xjgj6P9iA3LdnH2zErq/Ki3KRz4x7FTmmAeGqB3ig6gVOOmm9
dCufIUK2Y4wb3mtFM6aqmuPjOksRLUM5p+TueQiYRIx1Dz1OC412o6n+ZvCE
Z5wWMoQy0MStOAvgKiJRL2q8FBpT4LRcARr6NcgosnLXgOTm5ukOOq5/hByx
HljBdaOUdwTFeMWwCbpvos+hF+hw3jQs7LxzDLZGz0gcBDfJPQEPd0+jMa6+
iIfCGyKnRVy7zriYxf5xCSPnrGHlTCtN5iKga0XxX8Phq0T8+kCO/NgrWXc8
+Smcp6XYMkwf2caBKJc6gfJTs3TwIcpWdt0RaV4g3rH7tizBz/GpYnaktR2f
a8nCtQd9Km0PY3/k5rjrDs+ObkjCLI4F2Ca+J8RxLQBJRHX12m7FMwRc4Yfi
70Hr+kzl+ixZ3e/vQJUcpJC9Ydt67So6ykTUS5SGVWZ1UXTtKeU7+uSWqE4v
7HX7ImvuGLsZFgs4uEoEAuaskld2J2FZ3h9xFnMOhcHx7He46JL3aGfixQfr
Kw7axsXhiVTUZ1vHwiN7w4W11SssOsogEZg+nm5IQnyOnlJnu+lY9Wt2c1BN
wGStKx7IlEhId1WOPI4F+gvc+lzF9mjcDy/v5ocsJkuM6OWFKbLn/mAWKTsa
zzKdyoSWnzQtk0M+JETWuwlZUi+ZIhSeycGFEDVbi8rdeLePiafhOLjP0Qy4
3R8DHBmN+PpAbvyyjuanS7Moq9B+4qL99C1pTO56rPMvyZPnD8gUPiChin//
aN2fvgz4yZfBQA9RpIHAWQD+4GT6sj3t2RsidxvinxeNfBeV5Cn3hkdvYW3r
VbpbiirEX8TOLr/kZps4zH0nC/aaFvN0WBbPtLnVgvt714ug2zKDiP+ajCkg
hLd3/yu2dRBHLUT02kW3M5yiyEpAf7a3t/fliEBG1afWQYZgx0a+S5ySZiqT
VelZWdQOp+kWejYUCUpvkCt3YVot6UUn3sTdYYhzX0vJ6cO5t3C0/kGo7uyb
7ozD+eXEfK/AoHrxpabu6huC7GLJW/apuoAubwNBGM8pwDv8HrahQbWzh5Mz
j+gFwx1P19Rzxb3ZG+fWFFHFdg03IndghK0eycN7xy6Dd96D7Mv5Z28QAZUf
aaBAfzQkLltrTXitoz+ZaWwVgIiGzQt6gWd3jl5e0JMXHPB2iJwiFN5QajGB
qSWSxQ/zLLw8E49BY4OUamgTkWas90vzVxjb7O4GuP4KZ+MQtjUoYO4Ohbvf
n5Oqpy8hL/saMcX6ZDc/wsBm4KtwLfTAodqaMV8maL+W9WOncJhJ5MKorrNl
6je6yXktu41uIRSZXFGOyPbu83pjmPsgDL2yC5ULxn7KL450iJnYIJbD913d
8R5UnsmMAEkYz8uP/9YthlnE0nhC6EfG/c40x42hwmfI7IcFZubl2bJVYHOK
dxpazbBtGJtCh6j18jVkCzPuL5xoqlfwWqwF6TF8+U3s6qXHF69qAlxZ5Dim
ss6z/aehXMj5Vx9Ncn7q65dFvYrypKk82G3Deth5uTILjW3s9dFyV8Zby/2e
rherlphGmYuR7DZ9sgdN0dDs3MQAwCrdTBg4UaAYwarITs8MZvnz8Gna6C52
XNxbeqUAnJAIN8dvqfaoYEXziydeRh0Zv3bgTTCzYRZinIT5xRyBW+2Z0EZ5
aZeC8bbxdbr6Sb/0SKjAELt+/pZsWdbF1qq+oZ/SAAvXCm2yIrQWroBPh+tu
dP1+a17D86m2pDOHTjRjdBQIYtzL5TiXmSvrb9t69zEYxbx5tRth8/CNsMN7
cHjac2UozGVj61+Pz6i944aLFljNt1CU9qXLPieH0PdnTbt7c/a68ic4quXI
9dTNkoxxJ7FO8tNWljnmwvuKU/f7dYXHSkiuu3PGeyv2mNWLLvl/XWWox7GZ
swQBCDMBlq9UfiGOhSEwTKC4YNMEOe4bIgyFuL8c6YyZVHeFRELLFcI20jL2
3N75AXLWL1ek/9bQBgpzgzukwKMtPN/A5yT9AhcijDmuRy0+lwnRCT6fSeKj
bEYzTEoP2oFqIWB1OvABhOcWk2VMqVNy1CU4jOKyMAd0Q8Eu5CWG8ReVen+V
sADFXKKRjlmmaNEfsGfknfWEHkLmJam054h6Lxjr1hRuUzw8/8+56n5rQzIM
SrVbC4+kUtFHaAhVBVTjI46FHtDdxcfPHVDovaGjBGl57bzVP0IdD/zO9VVR
AgSDByVkHRVrhW70KvijZjVyfGjFkei59KWbRzGwZh+PhKEwCcHZ+77/vm7G
+JTPOD6Pykdhr164Qgf+6/UuOg12udgGBFpprgzq5o1IklLC1L3ZgdkeT1/V
K1P6W2XLLdfE+X5R9Tm5W2OFevo2fYSJoK0K83WbyNiFS4SBrhaaHJgTlW4u
m6zk25M6HykY3Kvav1DI/vRFdoUny+o+aHODP1E0DSmqD2ORPrMvgzAcDZJ0
QScI5zKsVTMHtd9dtO8JLZowbF6FdsyxUO/8BuJPzCz2bLPIKm5AZePt5juV
zY1VWWlHILnpvPZr32+Q1YbtMxe9ShLeRQTcDH21CEfp4wQNtzGzTZQxKaVP
qZ5rLbwNXUX3iPdUJ8OuXz569B3lElYgt+vy4fzxNgmPJleulmDE+l+d9r2G
go2PHcmKxRHmvf3qV1e3dlWgKBlSr8ldH0td2jj58VzwOvPnh0mC7aCfTmA9
G0VrZZ1896oMta5yvV8Hf1gp3xJe1VOjPQj/l9w35xDHsUtfnZNsNAlqmEOX
lvmGvVQuqYDwn/noG6w806USDTIGxsd/+7aWT1f6heuNn7xPtnXFiBH89XYG
pz/2/+pQMpop+T3iZXORDEsco2xfhV0HgrkY0lW30r3nddIJvApkSf+iprIo
yZTuVLjx6bWkyDC0BZRnKEu1HzBPUjX3oLWyM/XulShkPlBLh2nmz8D0cYEz
J5vP2Gb853fbuqUxenh4BTlpgIPka2FwEKs72LZgcUOcpc3YJnkbFwpkmgNk
CWuPjqcQQ8WNn1Z4qap6pSb7em8hO5GK2dq5TfSKS9o+en4fYWXw+C4oA/KZ
j8ZEJ68L0eow3YrzcPXEKLJ057ENIuXGipo9PwJIH5F7UGwCQ2IVfNcXDup3
C/BwgQz3/1Zgk0jwGxRONG1zLCR8/DM2S19f+esXOIhsJl2XBIPoVaXsyJmk
t1SfO8bVAo6JZEuoQWzZuCwwMkKhzA/qF0eyRQ0seebAecvCBLLcgUOECEXa
lnMlqQLWMo0+1gQYmncqaMCGeeQqJijIAJetsKbxTecvEBy3FfFMvIaf2L8i
Y67Au5+NpZHo+TDFW+zGNnwFHcsF3U1URjIfOjSYhRc08+EyAeILnV4Pqkav
OFbGkG9orAY3xXF28/b0ClSN2RMHThXGZYDWylpQRJm1fL6PJUdU99oeOerP
1+ReQT7YOOP/eQTJs9cfyIuOOrC9hlGf4PxnNzH+vEMWnwyyVBw+wziK6EOl
Om+DT1U2VSTQKtRREQk1qdAbpiVysil6tQD5PXMn3cWlfNscNnutUDBNLbDm
1ZHfXUnHyvwRltDk9Ft8N4fJUhchoaqzVoM+EdUWCXEklGQPAGd79dHN5eJq
We8/ORtMj4PIYg5Pv6ZuNSq9ZzIqnOgQDEXEpMPT+nMkuZ2sgeRf+mUgz2Z3
YG4h4q+hgRm4dPvBHDh2X+PQSM26bdSgUkcFozC2bU2TvDAYclaxExHV+sdO
ztz5Gf8BH0uR0cQM1HaSFs3LOkWE9YPtgG5pR5bkiLvZKQa95q9D9Bi43x/s
Dz39oXSd9kBHFAL/21E1Els612z+zwE54Q2ThnofPy+lSPXPPnsQJsnthllM
RcGgChMKqrRCR9GqpS8M59IQWScOQRVwlc9fXU5m5uUsem2RFRBwIs3avcHN
WeVhg8Qb83sXl9Qiik8BEJO/+4/+nqk+pD6JHrPNrGDQwqjK7rZ4FA2BD1Ax
puhQhUehFJizUAnEio3G6TSQKvzfF80B4PFjXRH4v1bjR6gi9vx3uRL77+Iu
p9JKeNakzHYamcigLBvGEo+ebf0wKqrt+lPaiSa6GCOnJe2C+xDw3MJBID9u
GLjdDVDIwpkUPdnl3fON47hw1yoUN0JADWOY4n3kQ17wxJHG3hHD+KE+wOFX
8gwNxYm3uUgKuC59cHVaaOp0rGCfMDktmSXYl04vFV+Hrn109vcSqJFGdcZU
23ye3Xb6rfgRnUeW2yfTIV7/kiRCLZ5Xp1fkTxNxKLQhYodKnRiVNKYrqCYS
LkugCoVNntI4/hVEkFdtIhr1bYpzTsbAVGEgW+CxUnR5M2X9WXtXAmvlAZKW
xSLXRkZcxOi6oivoqnJz0v41ZlDGe8IpRDi5TM+Ky27AVt/YZlMJMhdjSD5J
dDJKj9oagHaZTOv/fMTIXYoqnAssI3ELk1WE8FF9Fi+FY7B9OWCgAnX7sqEf
ZvMZXZyxb65waYeR0mMa2QQSWPOT3pMmPdv+JtXWe5ABChR0gk2JRiTxIzeC
6Tx+jdpV5hHP7Na0kPVYzLYpPVNyupusj8AZUqmsrekyacRN3wGXv0rZqevg
JWyMtLmGtkCuYaIHkKzQuix2TNAsXs29H53vOPhA6oSuEm2LN0aFcNGhFw7D
+GW6Uq5x42eIvYuL2Na6XAWFRBhVTJa2g0AOSKKLBgalxNGvCy4SslacqyVE
9cFqeFj25pPPIMDaoKEwAthTd9eIFip8jaExbdXmV3l50DsGAip3wr1lACE7
moZTr73szaQ5/CQODU8QY/Zuhy2QUVENzkgo/IJbPY7Gejvm9GWPT39xSHSq
t00feIaG7aIxVEBYBz8nwMofGjjnkFVSAWPOmcKbkttzyDY8NRvNSRjSRNYF
VnWMJQJosW+NtccqLG64PkcMvo6X55J8XDQVdEc8vUBKVV82/K4kkn3DzvtL
gz69IoNu3U+ebpUd8dFr7d9Wc2E/g2Mh1CY2C7gSOm3Z9RrHQ+J1QcoDKE7w
DQmr9p2rNwZjXShjur8+FHZAjo8Lf641yijr1FzemDSirYLurgYIdRZVLdJ3
AWt6bqeoxS0o6j9aIPmh2SvrUQ8Pz46+mU7D3x6Si8PljrTacP2Y92gluyC6
ohJvlDMYhCxF0lL2J+doxg9zvvFNMHftd5tkWBklFVXtSiE66LaG/f+1cKjF
YZdmk6M5W+/biskIMPQxFIBqMeb+T4kcAXC1uSM9ms/tZYfgOVsk9nqoCtcy
NaomD7qFKCRMQSYfuvruGNjYNSqSkfksA3fWF8+0KAp4DKIIeMBZsTApzw2a
i38HLMkBH/Sd8cWRfWnFu8yKpc1RhO0Re6EXpAIPY5/TsIvJ7Yfa8678Xklm
djNjPJMFqAUTUPeqB3pLpWNdz4+Hdkm25SspIJlFVUMAquz9HsvldUYsQHRg
e7v1vx6/Ym6j+ZD/R4Cg0Apj3SpvoXi0M8/vszyaInCAJISOgcAydRFzlGss
Wu58vw59+NfoFt0myJVN/6JJtNCBbkIy/r6EXyfI23d7B3pKngme/8cS7sVN
SP/iUnlFn5OwsgT9rCFku7GgrW6KoK1ttrubqYG4EPgWexofWbPHn+wlOJt6
WO4loueYPdRiQB+QVzgbd+i/saxOwXTGwqaZFRkH2F2cxQOJiKNkbd0m2NG+
Sdx7xVh5U7TOPQfZuzbXsCQ7/G+X41gFdRY1kOLdXvRnAkRGGLBCKICBByw9
mfVjPx7fwuBAp8gVF8gh7CXVwOUaWNsWQHF8XlTfbivZqnI467CKN2xawdn8
YBWWcqoFeDSX8ndgFeUR3gq4Fk5CApm3fkOz4zEz+tpbLRDBQYZxYaxLFqmG
LYrUi3CMbbbcOq174j2sineMQEs1/hUXYqmY5/WHZsToHfcuyAc2YhXLP4ie
88Ne9zN5EfHX6Gt3jzAHrHdltEy6IYvvME0IlpdOaksQepQ0OycfJpDce+eH
9MxYQGujiW5y4tlKp2T2YPDknsFnPYTqmMiIEnfEwR/tVo7xm/+VndbgtcDU
aIww0cwloMzY5G8RxI6gD1qo1HSrvAKbSGRHdu+cLfGC84xQtup8ouTXjGC8
9xPLTOd+oBQ0Dfw+mjANAWE2oRUdJWUgP2WDZHsk6ABUAEorekqGx3r6rZm2
7KPT5OKCJFC/eFXi6MJjl16hyFGyqNCMHcOJFWnx9NoyAG24M3dj0zpRvKrs
jWAXNObrrcK55cX3fiK5w72e42MUgvVOoyYcMwWbTP6dHQp0pYuGlNHmGNZJ
sAaPcRe4tyEIIog+9tsrRy6uRlww07XRPyAd61PFgyMnrqoBKDio7RdxVONf
pT9SkQcFtcVwFuUJvkA6tmTxLNefDR+3zBoq0NjSfM297tBV0J4O4YtCELfx
x87OdJ6FK8uJTsONuT7QaTWR0iEHVoAM8d832b6kALZtqgw/q86AnZBOwCiK
Z4PAz8GhkrkgO39Pzi8CqyAYTNAETE/Qdrwhm4qP9QqdAUslp+vzIO+pIkjS
n+7ZsHVVWnpNSQB3XmD6xOfuGEC0dxYLr4VXFlNQzz2Q2moCEYswQLiJ0fhn
A2udzMYh1BzxG591cSfhStd8lDomdAnyfGEAMhKuSTY1Bd+9989Li53SIIX9
3ML/B55JMG/rjcPNJRHEBZTka6gd1nrs3W9Pw8z9/nIqI6b0AKSknKGkt3xu
tgpphBX8yISbv+jsAnJwraGvDDn1pQgB/wnYlNhtvZ1wcGKQdtidHbu26fAJ
e65RwgQp0prFH1063+5E4ZJIQZ2rvjX1kqtXGMV03DnWyzH/ELs5Zag6gJqD
TT3ANqTGXIvOR/IS2tkZTAMyqIw/mbOzEZaP6v9QYOmmqwg8o/4g3Zr1z0al
CGxNkkIsExLE1P7SNxoILCEuiIa1WUvCe+HSzRT4XrXU4KwlKGWtdZ1T2ZZg
TDoAXYLf1hJgEZXf9Zhw2qCBjG/jJ+c5YdcAg6yklrahfCKvAXDFeWEtey/3
JE5hrCulwLIsNPcbaeVfqerkLgeFAG5r/MOVV/AFe+Gb+TLA8XG9JNtHK4cg
W1CKhbKkdkJIwWzdmvjg9NRJAqTvYNegP6ztXa9ayqteVrj8q7movJfx5PPA
hg19hl/pWoa8ZZKJlFrzBdyPCJB0sy086c58X6w8ykfuMkA2nQZmMsNsRSwG
9DYp+lFgheDc0Y5Q7V6f67rgoVSrnOzbh20MIgfZ+1GK4dS/a2Rajezw2t1M
2vW2x009AkBNA2+luLNXBVltIr78PSANDkiX5WvEgsGLYFGrvxV3tZeiarKX
SdinOjxIW3AsfQ22oF0VdTyoiNjeNaHUDlN4VPVukz2WiWss2bDeSOTy7R3l
HgodlI4aF9EoBkslhK8l5TJc/3nVA8z7NYGnNkMMwBKIrBjVnsjpihx+aiXT
4RZtQ+oNqcMUt58HnsCeiDNcgBH129eaRGlb/SQ20P+XwzDXlcvGWNYA9Qtr
TrejkerowUvAQCg8B0CuP6Fngov2XWuOfpupaCmAADlx5WtTPku2dqnu5i1E
eYSPxRE/KeodGf0TVR8P8PThVAK4eTHGrzNKvyXv5ojsoJCQZ9W5KUxs8p48
2rg/jbJ5E2WhV6bL0QDJ1IN+ZW46UCGNH0CHr3FS6shKd51LKxAnRgEXvhw4
uNkGvO1WHIEpmFxZVqqpNfWnkm/YO0vf/iogWdDQDtLU8OolXtNB5/DVhEaB
bNTye6OmcISm2WfWFl+hBoslh/Ju8qcdNeX21rNIelEYvYvGRS0pEAKaDkMv
5eiNUvZ6bBW0z2fPG6cy0K5BkrNwRAG7tj4vRgGWk11xItIRUyTQShllR7/p
IgukhQGIiHgNW9wa0VVZxyCQMS207iE8yqG7gCrWUfV9lbid6Je2yzqoYHlz
orZrhRX8SInZVO5oeqUHkFu4SWWoSfkMrY9S71RY0ZtKGQxqBgqbEn8dbNqF
j1rMB2BB7V7jiah4PKwp467w/r93q4pt2GIr6uGaGq7WKFRy8yans6vk27eE
2rn+uIupnFgBwKrYcqFrglaMGXNyfNOeGqztEXnBIcCOaO6alRBYKA25ssq9
o3pWwQDJ0ub72FGKHH3/y9hR/i2kFPFm3ZAR+TcaQgpJXRwDCag9IHcaq+Do
Ofl0F4k/EN3TBBFmjcnNLSQw32r3qln+WCwZ+3eZuqKSp7J5rXvVf/ipBigQ
a/I8oWk8e9Gwk2xJsFEKOOCrKxks/ohiyAZ0NIyH/A6hArI4CCUnHpVuuXJ5
Zar7pIw3w50yCownkFVD3j076PgxjyU4jxKtoBNF9HP7Con6SF+euqxMCAoV
9rqJ7EkQAdk9omLJpO93BxOvIn1E1psNGEL1XIvg08M/T+7enfphajjGJtmS
wGE7sEn/QykLD55uKarQdwov6UHFABkJbRswXsQbIUkZu55PuYNjyA95eGOH
ciVbpJZ0MKmF9rLxPoSXmcTxMGi1KBbZrJosXlQyFqtGYgCpasRcyuyCLNKF
g/HB5BbUIhG020gUMflO1b3XkpAIpNaA82XQF4a17qRsA6Z9EvevKsX8s1Hu
r5jFfjcFK33aZSK/z/OPl+5+uXzWtwGS+5zmlxILQ2WCfeBs7+qs3Q1+WMTi
f8gm8LFjNaENNV6DA0hl2PTWhDzQj0fckA1j4TdGIgpexVb7vJmJ1Bg+LbPW
wXzcXfHUDihSr5Lo6CPC0PScF1mTNBPUu9EJIHtFHAyYFtVNDrW7/AtmRvzf
y93IDPcQgqr7UxcOAmR7iz69EJkWshk6QYWYG+1IZtGhGzPcFiF/kB5yEtZH
FQxkLzoL7BL1u631l0E9xkP32B+XwYDHr2p3NoQvfYRDEvWB/UQm2ctIomjs
4kdvgpu1AhldORVK+ifkT4t4hK1WfgOOyhODttToxBNVCEOj+fAByGUZ8XYe
dqL1qRdgl0E7aMSt42jXOvh538Ls/qBaEvVnST7WdlpKKI5gbTfhmQxrygFg
vrrR0Rsd4lJueXWHarBH3Mv+IAYTveDMoHG7dz0XbPGY2+CQ/elVm0m/tOSl
pLut/MbGMXdkxkF2TpMpwRrbCCMA3yEUv2oA15MKAnUCdM7TiK7Jaf+UsDXO
6PaxA5jTq8mequN40wEee0MmQ8peo/6eOb8xdiDsFj5NxvNZRqVcZc/N9XoP
HF8LYnst/gxfMU1h5LWn8WD1qTgoPNTNwzcslEYJjf0KQRO2+INBdL2fHTOX
BCJZ8aJeX5j3eSpkQSG/WRi3xtc82S1+cgUgzrOS5a6AUNFx9cUX6SFfXv0U
m5OxNIKDh1N6QL1COCzJ4nFl9czSm/Z8BZq+MSgEJRcefaq0wF7ALCEZAN88
PWsGup5IV1CkQhreDmfMuOLAieVYoE3h8w3qW4+32CXtN9dkxd7ASPPsjC/N
sFmOc8/nQoZXguVF2eiEMAHlW/K067ruIzh/paf1K7LTGKuoehdXT1FzutsP
HEN5LWog2xkMszZ3weuJXhoKrT6fQzVcY4mHnKGmQPyAQL1YKHKRibL7zTvA
b9unVDvUf+yh5/gx4z2u6ZIF80bzClFjR31uXOWvxx9xwcVLStKIWQsHxM/Z
pNtM0ZFGJbojSOg5C/lnvZVvw+QGdtHJELAMibkLpwSVqNCHdqhhgsXddIA0
4AiqeMYUVxtfCQtIFb51ptZ9sSJZP+D4QMDKVKrMUs8rtzaEAWLH7od+kZpP
AKLUHead4TecIoLb3/OAdr7aH9iLsHuj37KW7gUeVRlboSfG0I/quEPEnxZx
+3FjXgmFrBKPAH+/Pp3RnIfUgmWMWlaOp5RsNR0/rLlHUt8SyMhEM+m3tQBF
kl67og9j2TEiuUrbt1lp0Q2KFxg3/8bvPMC06WM97CNJxLEIRQ0H+cFaEvRv
9ETqEJ7KTRvToe3IHcR7jtrTAy7LT+H9k+nzZGw0wgi4Kl5BgeRmI4Ii/oI1
+mqoCINwzVrs5f+11KG/i4o9zLzqnQVYC+09+kjdfrsJqHtWQBCF6wkZpy6/
ECVWvS7CD+9g8l8ZPocjROeYNtkcPYUbBZChRJqVpx9c6Wu2tPFTnePp2q4Z
Q3IpQ46X1HD/mEgv+4uy5zCTHrvfv3i6Cz1SdQVRhI/gpsRJTyS7ubveUN3H
P2eHirTeQaptr9jvhdm0EF+9m78Ve/PTmzSIh1I2UoAf3c6Z1bFdl/GmtFU+
2JddEUaDQdAdidc/4Ck3wohoJOwhxTcEN5GzyPyHSWZf/l6OcFGmWxJVDQ2X
LLKu3GoFMd4sYKQVJ2aVYWuOl7uRHAwo7g++6qwq3aieYL3LA4+PZWtBrRCH
YeY5d8VYn1mQ5EkcfJxnO7poY/RAjBbWdh2Y6PYhT1TubIMsJ60ZXo/3gAJw
EFFChjoQm37ANDi8vR0Ouw3yJ7RDSWhpV/qB9jBqoslO8a9H9va8Ovj0LzdQ
ISlPs6TvEQOW+pLw2sQfkAo9bpqCYhfx16CtNMZcm0+tv22pqCJUgFu8gq+C
prIvIIa7gyvBioAtVbZYmZnXvttjr+02SlN2X/8dZ37oT1WHpwDufZ5984ZC
MFoDDyyXqZcJM7Gxi0TXWO3kqpa1FTAKm4uXgXlDkva4pvr6XGESJHN4KMlL
6fgDnK/dGAFdQGnbtiqvyIfYGZ2v95MZUFl1GGWqkm+5gX7yHY9irUBrxDE0
FnZDbIhcLz927iT6EbPuvLQ2m5oTHwQgiwXCSutfVohnaYD5Apj5Kpvz58S/
9Y8704SdlkIdjvhWD2+2rm1Or8T40lGMvoVOhpy96fNu7fR9Yooh1BDFzl4w
miDLPBaTPsnQ+B1mXSoGOXvu56J42POCc3EhoaQ+SUuIgggZfLXgsfAonCW0
DWulnY00KxeVwupingZOljbMUjWSazCajIwhCZsdoJ/eyRHraa2ILCWE7Oma
zTNOJu8tHiG0eSyVsxBn7zUBZU63JuiQ31S7hPSmYlcGhyxBpESRGr7LqU5r
cBN723omGolVCv0hhNB/VV3ia5gxKH6Akm8ZvB80RJYZTJa0w3/vZSCdCLnU
+AeRgci/o13J3WyX6VshT/6tkidaL8JyyozY6UWf0Fgm4xgRuroO0w3vIFTD
GGOueay1B8JJjai+LNzXhF7gb6lci41O9FLYzTBbW8QEyprpWEIZMsrIGi+y
AUhd5OzAvYxTjkQxUWTq8mI6nDZwDFLYek3z39Q0YTYXtGTpi58IxCXo5IIH
Akhfo4pmteowdX7wcjJHbpnNT1oJ/OxPvQyf0sTL/4e8b6UX7cOjoC+vxDDw
D47IpHzuX/BanWbaMW5TEBptQXsqGAazDMVX24dLc43ZpwsScYEJdLk7/g1e
LYPnj9lXbeF6cyrrLif28cndB6EK9JxwslyaoRuRzERGYMzR6uAqHLBnF0K+
/TXkTEwbu0RXsHEqDPUPVPoxXsi+EXaWUmpKvZTZzqt8x8aTeuC4NunB1rtv
g6C2tA2HDhO7Oixlz9XmI77GawrnKgY0DgONONMg+G7CCLrJ5ikZH5kX4Vhk
8ihRuzx3z5uW/VUKKtmF/DOA4Bhl8g4S+3vELLBm4f7EvxLKryyWZyHCm5C5
JdI1J2zLc0wp5RyJ36K0KEi79PqRJImg08PGQfLX1l/hj3hl5VTGHApiMcTU
IolY0CLPNUFg2kER6zX8jgvITUu0REuVi9QFvlR9y6gOJH44ISPSy0Kyz0od
ibBXVKMevcyNCQAetFwGXFjWRrvthvkGQijQ4RiJL12IfutWMjomYAxWT+c1
iimY4PJ01X4cXQU91edJ5NEgo4SEhxRW8QiUeJ4ae/Y9SwYyCGILsJXx9Kvb
9SxSMeHYZ70vwWNZCh8DwyEScCQvChP+9eju0E+Z+L8qgQ50qTDj8jVb+0Hq
MV1mb9iXLM0C5KVMlW++H+Az8haxjDCjGzUtncCJJeKS950wV4cBqUskkwQ1
E+N/8NBCHJ6+hInbEAnGQQ+FNeTCHxuae17sc3M7tn7Nj53UkpcgUAa8iys9
E7zounUKug9B2bSoV+MgryBIEfN+VVWjY0UzWLQYGqtUbuk8fJUudYz1J5F7
K1rPuLr3tIGnWuyCzDl5xvV9puAzG/Ae0ZKdSsEWVh5UPIWwtg9oQ2xExta/
8XzDYQpPflm6rMrkUB+vNNERCCBUi65Gx8y7r9UeMrzs192gnDzyH13fb0Tt
8FeCcp0sTjhqM8W2IOl5zItPH9pd713JurWHRUwVYDV5xILg7c+HFRzLDvOg
u1BpJZcBg2VIv0o/c27b9h+GyR/JtVuVKKtzgc1iTd2o7n1OU4fKYtyzmNcP
rICD7Drb2fHutgIHtTRSS9zltP9Ss9MtMgjusdZTA5f0mn+0JBrc5weSB9BU
o3MTuUm5NyBTsQPDQAjHNI/NuNpuhMpc5UbWlPY4iYygzI/GodXdsQOYOJ8f
NEdEiPGZI+3YdrZslK3pfif+PXrmUqtM8lrqCdxUDmg2vuLElGgQmAuCzYGE
XOq4n93RNH7bgRvbXhbCCzIk1eLu0HzER3gv7JBfsy64yHYwK+XZkK1zBD+H
7b90Ubx6jm4CTy2Mjgw+e5tI9vvQ8j9rgzwRqOUDaXMeh0IZ0l0aGrn+a/O8
WwlbjHyf0aigJL6s4BcR0XxnPBPs9paF30EQ5gSPaboYmP01Y3LcNAoZryKl
/9UcWN1xIBxXN+AXlyPsRGDHnPHlmUV4N5rFkF7cUAsYTKRjxNZMz0UMdYjp
HOTk1aNcntQOEC7SJcJyKAVmbWOsS5rAdhj8F9nFxe3VBwMtAwaU7OYULXbw
1lLUU4THk2q56DrfXAcivraKM+3uuFk5SC5ftUUTB+UY18eR0BfxQR1zOQGc
lmw6BKpzAFsCOACCsMZa8IM6I5U7zYIcLSt/GCbfDPvf4afXAksUgDin14Xf
f/uerMnTZuYjl47T467DeM4xCb6N2az72aeToCMuMSVD8Z9Qq4nHet+8RVVi
zXYlCcmaNnSZte/EW1SrF10iLQlPuJUCp5i6kbioswe6yHvFJZMu88unO7F7
AqvfMg71aHTb5oH/OuwfuGiodBTz8pDBKWpJsP1WVOnE7/eWpNaoxoR6mq4j
EBMSuwFMoG8lucDyDw/GC/nsqlP2WAqiZtZFfs3OnN9k6it2cdFcllXdnmOd
MSiHXoYfbvKI6eI/3xRwXw6YBdPiDylx6hQcnPlIY+gqYWMXqAE1hIHpeQ+l
y/hmWcnF4WlXT3v5yI7TbaRvQyD1xc2a7vSMmQc7+zHJqQr+wN4XgsEWyizS
mWF5xJIqQmal5pG/RKDuVJk3T6ob+O5KVfJjrASAnUleMH5jKpPeRbjPdA3m
JCo19MU8FfC+fOvOON9LTpl0DPmhiZEs4Sy5eWPiaKFmSfaRFSP32cLf0VEx
62JNPqG9EyfoyFrNNAeO2KaIOMcXQSekfbFuzS7GuQtHZjQsUfeyeFh7LUSH
Fjy/G9ajBDqwOqHPdNp2korMcybIT4q8YjoAvT7r/kR3x2wgAgyioMQoh8QW
fqkE3rasnzVK5RrNT2A61fq4gxitPGVWBQo383xIRoF6gaOv/D/fLA78MLuN
zywSWlUZr/0QUFkzXHzrP8CW/58zHclZt3oJYakym1r64Iz9z5dOzYXbGBnW
JqugbV97xGiebQA5+JqhEyZpxREqJn7BtAJyH6GFUMfcjH4S7FFpvplvZxSZ
wtbkGeoGmBTO4FB8gfAU3wE2Q/kFUdaGwJXVe88OJF0pjLwJGSsp5O1/bjd9
+P1FR5w/M3sFlwCmzpdKL4Q1CaXeKrDKXFmanUxWR8MmzKbscYefN0kchyML
2gRd8PK5NjrW6uRFfQqiznk4mBHGjnPzqsy5bULNIKNAlkMy6a+lwAJ3+k6+
Y/hlWCnvJc2AIx90QfseEHeL+vH4I00x7EEzKx3fdcZfgBgTJvDAJWtENlrR
sHspo9kB18cT0qFc0woA0/Y2ZzrDBKMPGl5FQ0Msf7M4bk1ZFxDugeWVcOX5
2VLaeaciiwySy0xps4KIwj+MfJU1vym+XFaKrk2yYYHtBUgE8u1bYGHclXRU
YQYXNrBwXCkp4IM2+Mbbg6mdzwsbAzTUovk1l43BNKFTWt5/C+cN2LWUdYLT
E7DPHuvz2Qb5N8xp7KxUS9PAbOG9oGBl7WtzodV+QUp9mLXRJthbLADbZ3cm
RrzGbVennmM6wsMK7TCHodCly0b1APk+c0ZkitnEv0uEOSSzJqgW92LhkVZS
Tm73n+wp/4Mo2fR5DjfTYCUQ8BUoO5K274fKBGQL1K4d0hLueFZAFk+JKVQy
4QvKs2odw959HZJYWj7m4jLWfrdWMABUg+shdlo77OqnTi+Ays0iFFh2Ys3h
Ul121MXTE72qDq8M4XrnqKdmaQ8yRPBIGpbydWLN9yTLplC5LatTWM5j8bBh
yX7W/ueXQvkXXxlEQ2pIwmUo0n2E7bFdHUcLZDmte1Nh4AuZGvIpZP2ddUOD
YxsfDl/p0Y3YzSbbh1/BtWz5E683jjuRrpXkD2DTuYIthyYuhtRujtiiFAkW
OZ79aHL86YeefOTs/wwR9xGthgsCOOcRXvefYbG7k0gWpV/VaTUMiVblpcO0
ezKhUWJ8e8CYIcnereTOEAtNwe59B2ii660/gAGIV8tnIg8A1LG7wmtdvtCg
9xfR11VnPPb4D70FzIFkHLn7TjX8FU+xfz/TMzwgHjR7chWim9AemoDJND8Q
kMd+W6FkgXCUmZTMQB7hjKZ/urHXzdOSeYt9ix0RhgLBctgMlhyFab0MMDJW
LgHJHWsbyXKzAGxKwivxT24NwNPREz8c3wWxbeNz9ET7Px9zxlBsUu9OXP+S
j4es8hTrLO6lSlJ71cSD3muq0Kieh6ia3778a1lq2mRjXHI+u5AxW35+E6pf
Cad+5iVDY9DbThihuac/qn8MmeduRrBprCZTjXBFUktjgTHbvlypOo61uhcW
qsCiNjWZLxEOkuKrIJ/rkek0YWDM3VHf3jM+/uw2cYWU/SlFfJWz4dcFDuH3
kMc21uVvNK1BMD6QeQcq6w/3V0Of3p69YxQaf6MH9hnFCZGWALrp3+6i+gye
dGtLDn9GcPLHUu2uGUPnz15DBYkzFeP+0tRW/7+keWQN2U+NY03Rp64PI0Gd
AKO+9gNXdLVQONIMBw9PgQtfWGC+olk9CtAYUHbxf0T9o5ozt32Fa9kb1yMG
YIE4Q1cgjtmRVM6LStg3ZcgsNxRyVY0bK7Kf+rLbHhLDaQmJz3ts+nuTrBjj
JZCR9t4BQ8MsuQVs2UbD+m8eHebr4vB/Ie3cWiJTnC/z2QAz7ov2uZGhB12m
OD1CxLU53R3hbJ20vRK3ibrHP8WJYSzO8WNgiZUbj/OO5Rb0646ZhB2Vxx1R
NM5nOiQkA5X5hIkNtOq6n0MVNVN/n+PFxsttY3S/AlRotSnehM+HU+xQb2ee
9wwRbhY0uT7kNZIaDenA8Xe6e3JEI98RmCi18Qlv6ZkCFpd1Wvb6ToZGDseD
YD29PbaJE44+xVxvOI+Xo8lQUybWj6ffxzELPhWtMTFll66Ek8XuG/Rt1HVf
p/VnKtI4R4AF3FlxiCTQgqH22x9Bm8J/ajD8Qmk0x7Le/vUfr7jyXgkhJpya
ykOaLBVpd8+zPIpa5zoFbvfXGMFqRrLY5ilXo7Oy5xe99THtBamKAUdM8me6
vPwslAM4R68WiExVavuXJZMrYYkQtqSrOpiVte7VvHUTv9VLb8tiRpORtO9h
two0bvRIqDi3qV1/Zhp8h01jIwAs8/gMXsFNNM0VJvQqnzKhu3ZA2CFHjqho
snK2EA53Sii7kTG7u2q1nB0ZlaRwCm8EpNJEEX/c0XsKZQiKh+H34edfto/v
F+UfB/hhRzS6kgDjQKwiO8Mwb7t6MvFNcvrse5FXqf8ocLPTewhAmLZZ9JYx
dzXrMJCFVsH6o7HanrU89LVgdCtwGDFNTD3xPzKoiZ8+RkE0dU1xWZqJeaLn
rdZjMl9dxosbLXx0y3azfY9LxT/GEU4fGbkg0qnGBsleQvkSiHMUUSSVs2/z
eApH2qx2YMscbMGSVHgsX+L39TD4nfMWFwLZeVN5s9VmK2v7ajT3Hn3TRQgs
muH15MgYYbf15pN7c1H9+X0BysZbogl16gG8wRA6MKelLOdH4vMkn6zCiQY7
OEvdJ8HWx9of+T27/jgJx5aX2CE4u0pOrf5jjlOOp+D0nK4AjAxV+PPj9QK6
uVXwM3+niDK30nl974zkwE0JX9RjIXaW/voOy3Z2RZIYXGzzV12kV8iErOmh
L2S38IuJ7r1HAmwff483jxABndE7IzYhf7rOjrUZlsyrlXIP+e8hRqC1k4nN
NsjHogu7kgcJxhAe/g1OQ8koSfuIQRvvS427hoJG+7Pd0CML9BdYoE1HZDtO
KkbAOZCmSNnDGTqurgrPuMIQYPMBFtZMBy/woCLCbaz1YX/2cZhNtl199aB7
xUIPO3W3YUGiZh/wPO0BcT+jkWxSPkAU3QnhSgSflXSuPccIiiYpfhP7Bjru
7JZIsM2Ye9WdCiSAX0x1gLpvXuJfMxDMHo+TwZWopB2iV1CnZz+p+IE2YquA
CP78SUHlOo8483mhkdNqtihuTA19E1maAz1Ko2GVUdTJf99EpjYK32zNyNQa
weJ66qRIc+lz9p6fLo2kZUw6UD0A8Pkik5pToTyHO642iEhmkE6omf28LMEr
eoec3f1eqCXw+Do+mjv20fGl9eoM2tKq8q0Nw6E4xZpyMpbe+bYI54VauZoe
b9YmAkfEhHVt6TXIW72jkhID0GOXGcdc5rtmk86NTE69Sqjan/GbO+rjwVaY
C94q/y5f3P/xmax5Zn1vfGsEtdcGzF+ngzOM0w5HzIBeQA3Q95MVcGxtCalr
OuNscDK5RTcT0VYBaUVytI15CwmEJT1otKEwE6bYj+IgWo1cZ5d8jtux6+2N
38iuMgY3AGvoXFlwuAOBANpYN29TzP0z2doIqqbziHjEhp2siyO7veM1cO5H
qwAbYsxz5yxRTF6AZ8jeLCIIdm8eaAAaAs570LV5ddrijWc8toYyspTRWkOX
uQbT1gb99mCHWDm7+GhmO53aRy0yY8H0ptOCxa6ohRB4Rba6AasyQZ/SZZOc
gMXrYcyLZLByK33Aoyi3u7/KLPJVlyl3hz48hcurZJELHrIsNmRa5vK9XReR
qJD13e8px7MB7ZR9x+P/xeWEczJrK8XEoR8fAg0HAfqnFvLBn9qVhp4LLRw7
SNQtLTiM9858VTN9ULiQZiPOdV7Rpgww48roICxxnyrgPmj9qhuqCa8FD4rB
coyvY+UQkUURDSl+pwIaOKAnTuzZcMsrCLLfESIDsND4poS9XVkyn4LuiALX
OnDfgqylODnJfyZhOjCzQG3wg5xh7M6tKaBT6RMJe+AjVVOkua4kfItjDVz9
4TS0nLl7OLxP+4h0+kApv793zMXB4dhk/XfAMRAX0sK5T1hrxA5cntFL6Sg3
ZMHRZwqwvSULZuxhbbUcsNF6PfTkWU0f8qBN7/AzMPaTfXQP3Cztp7BB+zOK
vDmF7/Ye9FvfWsuvnlbAIaXso7BsOkmeboE6DaQd0mXMjIXBMih54j1MGdGA
nEEUJVnuH/syHNR+I5+Tk/6asNQfQKwcQ0mtuQKH/VaHyNP5TdQ1Iv4/7ner
32+BZOopt144s49u0mfaGzWASzN5EW+3P+UNbMsPc4f++bGaSs0jblYdl3ot
X0HyFUEFPqj9dqdRfdwsXUfHSLw6Lbm+etb4uGObpDSsca3Eb3w7wP7URss/
wSqyWcvwNiqsU2BBzUBomUZIkBGTludy9pMfJZhZRpf7NGosMTczjJuziMB4
sXnyyF+7eSLUBlRfQzeBx4RUFutloBQfhF4cPr9ywN8VvwXdYFAqowOnTg/p
QMXx+b+DjcpJJunMHLXmE6eeMuoLPOiZbvRgKZWWylXvCbehFYKomJp3GhYo
lOfuYjubSEys9tDgWxZhBYHI9nEjzTigCB2y721njdY761kjy5ZEWg/ZCrF+
zgO4MqK1dyB74R9CfcrBrdMiA6uCyb6tZxF+2Tl9UlwW56R0KkqcXl68D1ia
yPVgnBW83nRUNzA2PClAepJsAUKvg2fsHS2+csrlMtwrooYB3a43+xLLSPKZ
K7K90FPU/ESnK+GXgSiJ1o6Am5yiAqNkU1YRQGFsS05TW67kbgHgqamuWR0T
Xh9SH3+sNDK71AxnCrqMhbM8JSwRDHwhVfMl6r/frSlXI4vpaNAwMdy5HAIM
cb44JTiU5VZi4qZp8wvxtKDfTVFf7M9YL4NzNzzKukwAWk2GHAsVq0u/QV3z
GSzDV3B6m4xi1nOCWEMVUdK9HEwh1tAyIgcFJA+68CdCpQxa5TK4T2co9vmz
pvlLz4hK62tk7WlnhEmSavQRN60uQNzyeHFNyGU4c4FuHRNyXy7BNvTilYiq
o4br0XeRrnZRFXuoyX3Q6x5pEVcrRcfEd6TO/UdpJhOHemlNDm9oWCttmjwi
48cNKzqQBnjjGve7N5HsYa5B/gSXrMe7Xq/cfsZqJOhKN5nShQYjaHoa7RWA
heqP8gEoBSb52Io32KXkBS0di+g6PeKHv4HtJRNX55bRODVsHMilb6S9SrsS
zdPWgv207NOzOaLD60i8Q4ldMM6AhnV4tdP/YWvlspOHydSC4RN2h+tO3dPf
+OPjNZjC8FyfBNqmc94gxe8MrZzLmfmEzAdCkTvGdeNCoKKEnbVLgWo7wXmx
cGC18UfeH7XUacFVk3eXwSOdUhMVc9UAS3iSZ2uGonmo8QBgO6ciZAy0et8m
nVg6RTjZEf8mPS6diWQE7X20TjPQI/5kQFeaHWWP0X0ApfaSoSdjvkpu8UD9
yPj54p97RNEb+O6/FwFfkfe4a36pNZRM2wuUyMycGJws10MwbBGK4h3obtwM
JYrd6fJFyxEA/QtrSv8dbxG5gc6q8YRpXrfb6Tt4ZgjS2x9+kG6vWYUbOihV
fkx4e6D9q8GvIiToC26BT6NRRjmXiiP1T1E7+PtwWLRyYSixdlCVRTBheQ4E
30+VeUrHRLG5KFzkce4oIuvwHbWCwGcpDDs+AKUmgSUJqtgRLx75oRUHOARk
c65xdDGNU3nlWc7Ngxgai38bRqdPttbgzzcPkICK3uddBGxWuVZ0XZm3lWzm
J1Mq1/d42PFxeuCknJnBuz7YsE/OikNvQ1mU2t1ixhzEKm5DPlofQhEMFX4+
l78J1NjnDjft42zFno4PDrnhWRNIDzBJkQs5LLxLjZ1VIjRkdIw/Vo0yb3TT
122/jHHripNOvvYGJUgiffLZDZyJadXKYVUKjlbwwlsT7CJdArt226nAnio+
a3splPzYJFYOWY3n2/cp+duVLTwj+YWKDY6o1hW4l+iaGxDHvJ1lnh566sdB
K9EA5QOrxvUhmQWWP+UJzD7JCS6axIvdNPk7wb2xcTlo8qbIqzz/YCh+2pmV
rrKWPAjFRSP46ZQ9Ol0GvkWEcKntkaB+kcKMm8Jkzm4ALm25mx/jAs+bhHXU
hckifDw/RJ3KAkCAzM0kmhqJpGS7dI1E1EgBIp/5156PkH0jliRyodL+4O14
wFdpiHJ9JL2F5eCPZAGMD84PteZQXO42AZFn51HNHWCjka0Na7PuJ1TGye/E
h4OXB1tPKJoRB/M5QCgRpYLXRIxaMNEVQ9lFvrqfvUQpcwTNnvxDdAZSau7R
ShgN4gqDAMfEFJMFQd3tUrpri57lBiwdGYhIDsBOhXo7/WFdXFHrk3j+DR1A
orOYp/lJmC6S6cTchx48bHxEcn6vMptxR50lAmkxEZuIG6J090aCKjSWGQb+
akpVLtAt9sQni26i7aNPzSphOZD23MzWBNXXHbcY7Y1jM0EzmjF5ppnWge7r
LlyyjkpGf3e8DZL+lH6BGfu9KKKKIDiLOSvDNmONAP6a2hNN48/1oMAs6CWv
FweBldOC3AOdUraYBO3jE9GgpWvHsHhmsv2sovANbj1evDX1lsBaRwC6QB5i
3voQkxrV8ynyIm5mqtWBSwVS72Vr78zgAQzDSgrc4cx/Q5Izi8woyH+ta6UA
7AKyMbnSASY8HTCO4uakT7DCk2CZxJnCDzIUgYazQxc6BmYARiwc/DzdeiH/
Rv6cA9UPV33IdOvUX0oYodGH82papAe6bARHRDTF9R10KfUPjLmRu2qxX/tI
QCF6pUjcWylTFGvk7pRn96dURE+n6LEtwACABFS69rfInO2kjoo4GzWKlwIh
Jb4XCUazvOukCtPetU13aFp7WjQh5wbYEGqObdSdcldf9x+H7nJPJdn9vEGY
l4NwOkVjkeoG8CmSdtgdTCYn4xHAgqpvnnzlpDYc27e15RmoUArPrVw4m0Bb
BHS0hvtPeyUmJIJnDzYL60JHiaC50j+PHgGpycP0XgB9HpeYYHtl6r8B6H8s
iwn5x0aKfhvvMbRJDC/1ptakftRmYiEQFhAuZGuaURRtwV7q2WVJEOlvwzVb
I1lNH9IVqwyglfWe53n+nFhhMl7G0cJkuEap09cMFJN4YWkrN/w6umWfV8zu
3h4Q7sV6oxPm5gIBDq0MMTvL+uVBReW8TEiCyiuH8mExI/OBqiDYmsShE54z
2WfUrlUP8I3NbEWIbR9/HrEv+Kj7R7ScWwL+U9pBPSkZ13ZYpKDhZsm6iDTV
qHbJ65lLcgU+ulv4nZlh1dAOeqy7G9dDm07VLBwoeZExvSfEc3scUwsGu0q5
4mQzjoqQFUWLuVLl0qR5a/GqVwP1Urr5tVjh+rABxnUcup5yG+cU/eJEVG/6
+4joLqfb2Uvsfi9rWh/g+nGWmk7OOCStT6H4R7GKr4o/PYOQKwGrvXAK1EgH
AoJ+mbFc2gHsKUtDT0MRrgItpYnFiKiRjoaSCTWVhyTwxzmaRMviP4bXp07N
/7XfrzZyDOt1GAI1R+aUslaBPZJuhb+CLAzT9v2m/O0sUjkzbtFofdcT2Ppk
7+DwLTMQJPwZbfCnpebFWIlN0EDxFTNuy3MM+dBuPaRaVNFnRj3ZmX9VzlLw
5Gn/3DojcCeP7DI3K3esZmzXqeUvMIy16TwdVhu/OBryufiX1cgA8KaQ4Ho0
DYqz9t8+QPctpItg9ycvhmsnTcO6MgvSxRCGPD52fkomAJovU1tm0IRPuQrN
uB+znjhgk7rMMZWkHwFCWZIGI59RwWUYBcRi/fxBm9Ab06xkYOrNyq1dnlK+
RF0c2LIkBHW6sES4gvhu5chlVcQTQb3BlN9Ca8pWMmRXLcLMlkPnDP7rDgjg
Q1lD58bkbiSBsjGgs6UzB9dQM97gOgX6GvAgT7Fv2lo9uprF4LBQURHS2fKf
MaBtJZzqONv3JIwrwfe+eJarx4Qmrch3k3jVn9f0qoE7ql3fmsmmvFIJPfMN
6fjSNU/eW5xQEqi/M4MIbS7R9Li0PX2KwF1asZ9pI62m2NQ/mjgRsdbSK0Y/
6F89VjEDGb8F/cbVmSoPmec8p48EY8wML/dZ0bNqLdpM5UhQ+iz7P76nep/v
ttG33/TWI29AyQqrBRIjKpl8G8EU8fIggvlO0nR7eBs0Vv1kmw1dDrn3QDj+
cJEmKc0gvtvFYkSXIL3b5X11J/YdMZS5+l6kv+XDWG6R6SgOTEKeNvhVsH6/
19nyx39u0fgg7QpDKKs07kkoyrtVkVeAQrvX7YG8VTUufrwasCeVU8AN4Fpe
HrpSPdmN+uc83urNmBHdD2BFyzGn1fV3IIgbetyVsDFO+R/F++LI14cwggjV
fMchWeeshZakA6GzLkNMuWg4G8l1no4cAsttSgCvhb8eo9ZXrKtRXwvFV0Hi
Ki9dFTwHS+phyOEpV1pNznJKHh11uUAP0gE+r18MfJSNexJFtjgE7iKz9e8X
rEaHk4iJDIDrd9/aTeZNy8/2ZhVePbKDpcvbavNV5M9d5QxWsUdfky/hijT1
ff21wEEpgDoxGFLMSJND21e5I48Iu/Jmq/OebLgl097JzM4H90lRFbcK3btC
O1bQNlOTqwBHpfThwiNXOJ8wnB1G2aJmZPeJNGQjWUAQakcllQFSaqfNQUjQ
q9ItPF8Zvhju4esdhZTZx2cVJALvGJjvGSwWUDzAdhbLT2fK/MsLq1pHfc72
r5ZTw5GCMknbuH3LKjIn5XQPF/9QmkFpALMZnGkpTPf+yOlsPaU7bINePo3J
n195FLR4G4JPlMyE+x8ujEmUGJSItZXxD2wDDSwWoJK1ckTWVm8/Fta9aPMj
37g3AjiRXKq0SvWbrKmPNxs0ku6gH08A7nv3R54LuEDOt0ehCnJRotyz2OM8
L+gZfMsXLki5eKpGBxAM9YwH7VB66nAkH8ResJeAd5d95qzgkUMZUlNiKIQL
JnxyZatlLjNMNDthjnRJcSJpEZ+pIIO3B0GWmWrKUEa30pcJDV+sT0J88qae
Zh1LkSnPInDeL5RQerRc9+Nt/hSLKIgl70HCnDz3u/ZhFx1akQN1UGyYIQGG
zjYVD7HoDCurabeORvlIw3yz4fZIK92UORmn5emRwq8hhYhug4ikc0PF5VgD
OGxktrGm+2FrBhQuTEMM7GBVnx7opY19CqXrCuXTEWmRroi/eexYAh69OS2v
JChDplf/MqmfsUfAYk89MeqlXYoGWfGkoTE8HvQWlaEMMxA/J/2JtJmlbzQ7
3xrjNTGQV61CFnx1JkThLyMYwg6vXjQlNBzh5W2o+cfhPt0HofyChF8Hbw5/
/7hib+avklyqde8CcuT/qVYX0usu1H/jNQDVD5MktNw6r1EkAgczsNSErmGd
kwg3C+EztfYFAj836yPzg2HrzlOT1VtVAvg+9ffa8Z/Xld6RbtjHhisdXsq9
zIrYUI4ov5p4nrhsOwebnGPWk0oBF7oWUqYim1QnTKBxT0cR2stnYmDhHjAA
v/VnOcrcwYYt8Skw5jGOMIp5r9JtPOg+BKORKu8mmvNjOYr78eVDZl41+UrY
JFpiawMO+xp3EpoS1K9sn2ZfsrPFe8Tb9yr7ZcBUhNhh/gZvSn863vv6FMz3
rdaKlxOdH2FrkO7Tx49OqN5nRYt+vNFMDXSGwbsJl3iwhAcyb7Gw5hugbWZd
P/LWO7z0hG8RhkE/zO+Dh3QlEddxvuv76ow7uyZ4q895cHb4igcC11zHerPv
WMUWQHL/czKM3/XLK0sU2RW/iJfuiTA0X7JoJfLcuO07pM77X6OAZIbfrvFb
zXCF56NGurqA1sqg4DIY2njf3lIDjhjIPoNuh/M267F2MKXKzsstRFjDEsrd
G5qaAAOsBpNyCYS64G4kIsy7Guew+2XYlOiibsUNwior/VswWou4wx69xCRt
hMpkQdHxWrXgXXpieVuYdqAh/8kWFpKFIaa88JSbOHwQjAg7EMN8zpl+1WcO
LU1ykJ9eYhrvpjc4TJ0MQ+H9fJ1GZgGtmAQuXlb4VgS0BMoUey9j8ymjwwci
LgZvgcUCkk6jWY/f5OSSoyRIBQ3tjU2NftfyYgCV2GZ64LOUXDy0c4e43gTE
586vZ1RAjWgNwcGZc2uPiVqv9J+LEpeBgzN9bNNrvLnkSncY/jraR76Jj8w/
3um5L48GqPVXbQIN1tS2d4Iw37fdKD5UrRRqwgtZ3i/IyvJXkKQAtvMlYJvQ
Kmf+2dtuicIYQzOUzj98Mo7lewbGXWRnUJY2e3Kl/ttxF+QpPhtUhFGVy50A
QpNLAsTCshTHxFgRDH9+c02Bkr1rFrfZavChBohCunAB6t3HRP/H41NZzs/g
6MU91D+az6eGTvKUSkc1aFFLIgdihMFp9adS68ynrJUm381Kip/U2Ni/r53g
2zIldfjDRxcyzRlZZBIOE6t0ox73SxFKlLXZ0m92vKIVIFM7NTK1EAhvUd+a
rHjynQP91ux2Cj16/5EpeJSOnV5nF1v6GJ4So48aVMjzd0KjxYzxyAJ6ijgd
e4xLD100+rauQHathKMmzE+8gfm59yRuuMdRu3eeyyu6vaRb+lPb1OxqB3DC
tLJWs9ftShn3mk2mQ4IeBSIvKr0zd95RbqGQhuUApKKWFQQLz3R1bVlJzFen
TK7HLxYc6chhyjgmw0ogQySI0dwaovUoFHDeY/oBr2wzQIg9x5tS08kmkBTd
wmgotfAjeHOGY9p3oWy4uoMDgEiTWcL6wb15COPmCZOnrwnifgrJaTi8VZuz
GvjACXcTLfwn4usr75BCeHTsEVR6iGv0gqbBr73suBqsvKz5uJK0FuIkdWm0
XgmCrjmClHVfcQdAxpphGgOCDcvTqFqac3aCm5Y2kuXLC8onu0lFL+gk6xU8
+MJny+jvej54iRxOhSLbx1BzMWX18jM16pWyx7+HI/n36b17zfDOfTmBXpPj
X7JJbyyWYnLSzbZ3BwQqoGcB2puX78rHcMsqweXbSWl1s5q4H79W+11d5wK9
5asnpfNY08MeX9BFEH/fBTOjhFT6iBOmlGDEzWmKTxYnAw509VV0vPnVUuo3
7PrTs5OlaN1PJveKMHnjGRY1t/SliLOEiE+326SXozVyaOs+Xi+gjKwPpe2d
7wrJaszH58ZB3P51DzkiBA2p6jaB1tEPFc2GbGgOtyki6/khKwzP9a7c1Nnv
5rja227l0OyuE8/zseJOEoDtMgePDM3mxgN+6y5Ihs6x2mOxYJZ8+ZvLwp0w
c8rg3kVRwCKjl8/c2NuWBUaE2NppJMPEip5EuEcREgyW1SN2hr5ERr26bHl/
UtzQZYqBE2MXSROcWA44Qx7C0i0jXnFMpRTJ6o06GFy2fLdvyp3H72CB6njJ
tbMIcQ0xGqT6wfShefb4bT0HKq2Dr216iwCZSUyKMAWrSH902xq+G4L4Ik7O
21ML1BqIkTfHc7seAn0sGTXczpiVOGr31r4tMsH3YKDQzYB2vxpFTnfD4FnH
TKsd8CH2mSbYwiC8GOq9zbOJeF3SQKhqPb1XcaZtDQelv+ur+0+1Ewbls3/3
nFtRuDWgEybtCYkJYAMpYimkpWQxaVgjHHx+T01QqXeyLekYxpPszLD095hN
8MrAjn+D0vBtHD+nLV3B0vm/swwYjdqGj09knu2Cz239i/XL+68C0k/Y5An4
NeEaASwbmI9LAc0E83pnkZwnvz/GTtfRQDNdZfzM27IKmQD2ApTIjMCpGRkh
dyGgf9GMwtjsOJryYSCxFdru0aORx5/8CV29Yn+/oXbO3GsD8btgseYGZU+w
U64KflMJzfpn4QIoAej0y53Yse6waJvMIMbCcDlAWtPYIa0hj4naRl8qnNW4
YSpVViR4x6b9bTlvq/2fsZEyDtt/MhTPQJNdg5EqbwuTsvTvSvUDpO+uEXQw
3PqurCeTzAUwB2sCRAHk3/njgz6UyXN4wmK+Kl03AlzEuO9dpEeBNBItYyM+
AfDOAZ5+DtuhWE3FX6g6WTLbo+dHxlK/6oSnYkG7CcgTnAI/jNq6FnhWNgKf
pI1lbMFPDMx/1JqbGjX3FE2vUgTq/fPZGXlI8EyOctlpoEIRc4W4Dbh6SuY0
VltuE0ebWg92F3A/XNG0q4JW9+/JvmLgeTSpyf2i2xo5oER7bueq+xaYS1ZE
N7FvhNChm+7ym7sl3ZL7EwUN1GUUsMNtLZn4VTVcseP8y1h8Qe1CH7Ut9Eqi
sGKmFeUTyMXUSe/j0t98dyVO+ifN0xN+9Hou5fztceX/p6AcSJwIfw+iFt1x
1kuCbWDq7EIVaTi3ElP2l/jyVIve1fwxPGFegkkC0vjF6Dfw4snRlSLHUArv
DuHd3rNMKYeTYSMNxxlvV5QECmNgHRG1vKYgKv9thS2n+pn7AFxcEMpvcX8M
xTdHKOcPTDjozI+Q26bITcg4aNTOXho7pcuZmJTt7t8JXhTw+X3qw7okx1rB
wGx1NW1gW7ODoh1p7v+CQgavhzuR7dgtLyyhSTClcGB+0SW0FjyA1BeLZ0IW
Ad8nRsZLsSIooUL0HzPKD4HS2kuz0UAWqyRxN7HHXxhxKTVTE+XtzmsekhXq
Tp8P6meGM1sHo5ZGMjs+rQrZ4jtL+GHZ8lpU7DSpBhvqwo7IXHeUyL0gaMFS
CJLC1wxP8vrG06TJIPZEPKSwVukIKRD0aEljTC0HmPOg3BVyzNjbmpLUGA4/
Xkl3ZUKiFMvSoWjUkjzjc+gxyfF8XC0b0lFExZCYt/GzA6nd4VWv0oZpXcQG
nFH9+HIu23pBDIpZa6YekdZXyVGhb+fBa8H2IJjMwOBWBokvITk/Lu8zD+z1
qwlX8WS8O0gsKWqJsxDCs05eE/Mh8TXM+Z/pWSx/44SIw+5X7xqN3/4egHfm
GcytPwzwK3QIM+UIjg3A5jxH/YhzcNDyP/V/LONnRObp37NLf9jC9JBM7XOp
WMSuf+hSglmm17bnsMXfiKBk07x1ZcgGt+5MUY1U8KGn1WhZCxqqo1EfJA3p
2NIUYZRfcBwkXIP66T8KnMaBOsckg/M/pZMwQErm+kiGZxsAq5GzVutcbt3O
y+uTUlVSjZzy8LRyehzBxZATxOc1bhXc7VgR5s7gOVH2HQ7/ht7et/Ay6Lu6
Z63boArOulpoVrAC4O1BQj7DZVJBt52i0WttDwQmJSvSGy6WFvUyDA+ZjGVQ
Nk8uUH2LEYdJg9e5hcmGkMgIu2Fic2uYlVBwcSa/+L8RyXdL3SuQcO6AGOOk
T1QE5jX/CvfWFKn9pbtUHDA8U4YPrApGLCjcxE9GiqrhvFnwehmAOcfJ4uDp
ChcCyzWB3mPW1qlbafJ2yjIJypGq0S/rvgLhRZztGlVxSGPnFgi7U+A0NfIA
txvzkXAD/K5I7aLkxcl5o0+dTBr6mTLsm74BwzUs6a/Q4wIR7tESxqsl/dbo
gJ/OHnJMag6jTe+rqHScbK60BEUMuLtcvLxR5M9P/adUF2LniRuK+Q7wYkyM
Qz8E/q518EI8ZvmQPeZWJXqc8T+++UjBYBn+yykRspETg8Jx+Cr0Sq6e1svX
DUfCDWUN2LxhjTAscBA5bcbSjAZqUA6gEHr8AYO0eFs06i7w8in8SGcyP7KH
eot8+XssRSLckTQx+zmWQW9ABKPogF3wm3LMoKe9HsP+3npTFy09upHAr3/4
gG/XDt2yndsb2fX7QJeWJ4yRVAmM58ynRi4PJC/O21sOWtmkuQRVxpKSwY4/
nxTwkWHb2die67eGROOXaF7SiiS4OnfARXx+I0I4Lq+hNqb9AQmkXkMzq1qD
pIUHOau2lFgm5YTPUjmi3JteC2vb+NvlhVJghkFwScKLGBoNGFcOWVoJ0e0Z
TpUAvYx/h4muncUkbYng8ytn60fuTSOyXN1d5JGC7QaOzSdDSlPciVzrilyJ
qrsTnL2+TxtOZggtEyvkmDwxWN6i6fU4WjiaIQMNU12S9fMZ87AGovBe8RWK
VDKYGIGZ58mRToy/vuQJcI8jGNHm8hjeqnBUq+rbmLph9GVWqEXTmrURvZZn
oE8fro2HgMquZJOt83II3qYfDG5mfRSx6Rq7Y1SEULD1FZ4+x4RUVassAwjP
GHz9Cau3edn5JOa/DMkvsmHazWxPzeeqYjMKGXNnh40ERHVhQWJ2X+NW9h3C
MW23N+/vL23WkxTgiNKc5Jjdqp7o20f8SCOqf72D0JnQMkT04yVRtzKaUH9A
KO2gCOpwczRMetZtwdJIIm/sF/U16c+ke0BeYtEaSn2DiW7lwl+QcMp65nsy
qXl10Rx6MsFSsvtwDYjev9fodbHoRJQexwTca1u9MGG8jI/xzuPvXArZBYTm
gs/d/Oxuk+J2aW5PtEt2udbzCwyJwLb19l3IAgRkzfyvlMI9Pdk/grSEp69D
0puf78LjPcafRkscc8FrB7V1CRg9WHV6ps7+RqhZv6TJozI7zdirPnU1vWSL
fH0d1m1KuPk/pZtfAkVQjUlVyuGy7Jq8DzogN8vDmEVFGLZ+GmH5Nd+9/zE9
hoM6ZkW+ymtltaXkna4LRLG0qCKxv1skWKITH63fZEme1sioO/KYQi/C9bCC
KnvLb65IShd0hjEXl3C/fCmdeNN/ShiS5IDb56MJE2hjuEn66PuWHWU7W93l
zXb3nYWqwHAcYj+pRcXbKioda22B+jBmBR8RjcnEHIUa0VHbz6fSYV36i22s
/uVzxcJTi0Ppn2/XwMPwUQEI23LdvsYmueSehnp06bhiMktt9c3AlSWhJttO
cIbnUQmwHW39zoVP91c2MVqTMsGp4QxUiz4NAAvUDH+BOX5uK/nz1KQOER1s
h71Sh8KuQclwhpIK4/UgrgZbBKnqbIr5e1R3EQn8NaXiT9PU0mDXIuA/Tayl
myIcaW/1hki/r3CDRDMmI18mm0Rlls1PoaoAYcKqmR3CQxW7aVbYX0pChG5a
yfWcytyC5BMagQaFkLL64yUqwAWj+BzJVbslGxEPEwhaepdbyMc4vVhx8bb8
qZwAPhxdHZrfOPpIV7uu7uCWUBSvcKbUs0c9vCNK7fO4qnVdlxds9dZK4ipn
k60dZXYW9FVB5VChzS7oosVDFZ1dY22n/P+UUrrM9djBNXDEwQ+bkuYSifDh
Mlr9qrmQUyb/s+wDXLXuaxv+z7w/kmYex+5cHqVisrb2iGnizF69pEAMQRaT
LTyh5nBBGelmZ6mGk1P0NTxcy55wG04AY2i7xRR4ww4BMzzj9QLAtIXiIFhd
vgwKmKfeVqXqi7WRyafw91pQV9Uk3Kt8cwPB52HpH4gOlbV3OOuMh6Tww6LR
LMYDAohJaKPhKWYj7iNjnXNy0UX0JQw0l1MznZRIEuxXBwGQelgPNa7V+1iF
OplHv6HpU2cQH4hua2L9CE/z9KeycP3YZbEOpY7bLf5967A6P4u9rPz6yOzB
qpDmuyHj6Yxsl+iS38BopduKxpBjb+Un3PDpJxeCq72Is9HzCHgPs+FWVy1I
Soyw5qiRRSYddGEs8kn98uZAv+bOT1uxlMGy5xkLmeXwsS/BC6dVYtnXf5wf
yix0txL34ndvWlFOZ2+X1ygIOb2FiqlOtsUi678vMZUyIT7Mzx2tFja+4zHG
uAEjXK9AlWY3wONkoL2Iz39WNYPYOInnrsTL6LsW2QygeyPxyXCU/tYOAuDk
nEH808OZhoQqaztv3npwEWOM3d5SaoTkyYAIExjYhlRZNZae46Vr/hL1ojBE
7YSUAJYhsn1DOIAzSfpZxbHRGKfE0Rv5ZQKAcz3eJ+h+f5ImgtMMnZToL2JO
pdNC7zdOcmYApexxag0R04YE8vnvqz8wFsBwYaqCwn0kNjCk1/oyINvQtyEK
qp6WW/KW6bYsME4WJFAJR78sdto7HEyKVFlnBicX8Q24i1pa8k8Qcad0zKMN
e15aUm8mcxZjyTp5c0tojPzYM+SqMChkWnNpZoYONsSLpdIpYVQEeiVuRtx1
IRNu+gcXYNeapasaovoAb1q03/7Zu74cwi9fdgw54m07Hm0kqLkOaaP09NC+
Eb05K83O2avem4l3tq3yU4QEus/aih3c1II7uaC551lNKW02gVWDiH8XFM7D
F11fP+WFA0SWH+OZcCVrlsn3uBnxVCa3Laleu0z5uH6mBnnFqVk6jcIh3aUx
389sQx78EsouFQJ7saC5dIBcb+uKcfcmPyVqXo+vnE3Thmb4S6IAJP4NmT6X
/I+QSbQsDNiLJ5pGut1QXY4wzXui4TyQ1cFKjUm68UZe68clOkOG6Dz+smvv
31noR4GwNZiLKqWjvn9EVY5d53e8+OAoLcw+lM9YiGUNwzUq4PsSqcNlUKlm
IGahyDEPeZUfreWH8VGlvYok+gBjIO5P3SBlE1uSioNQyPP5fWlK4odgj6ob
UOroOfLgl92qsUauw4K8uMokyGd/R2vnAq7XP/xKLKS8LATbb3MU+kKg8rFn
vzICWm59FFS3OVdRctZYAMpvKLf+iXvSCY42h6eh08+W0LjRdGSEDQEd+SSL
pZEd+4KZM07sxEKIXFvI5WU1EYVrVZniHzpqDA6d9U2TaNHHKTe/XNLkfDi8
kymE4BbIILl1ucrVNObqcHr4JtWBJJm5OwZ5K/LyW+ngFIP4AwE/J/DAJLb8
hIOhWEWNyX+1HrlbhF8jrgXf4qIZW4Q4G3zO3tW4MBT1L1vATCdvsdZw7IKw
NYGndzFT/jkIueyUig9pkioqv0P2AU4nGyLPIbO/4mbe2+7rdd0iDwQmj1hM
nRPZG8szsI+K8rNsmx9im2ay38etUccYhQTbQPDAfj9HM7ow8puT8dzHqIin
LSroK1Dll/c/M1z+7I7pG4wEPdQ24jPB4wtacE+LNsVyKZYOY275OEkEh8sk
F1K//di9g4GwtZO1/O9cWO+YvhK0OzhpsGUQM4Co6QR1QhH5eVSuDwELvmTX
Bd7B8QHnrP2tjUVbsnZ3K9kuL0ZlLT23Ta/YNGm2IINlwg28j7Qnp2ayCAPd
CUVEzXVswD3PIHu20oeSTveNM9MN19XF5S8fn2AMf01bOvjq0qw0M8dVgeBj
ATnl5pJaFh6Zm8p1QZGI8bRpcGZmiizdZyT/zTKHjhJtvZvqLaOmG/WM4QCE
YJ9wQiAS7hGPkyfg0DwwyoUA4WaxeVppwzPn+GBjljAIepm+TTOhTX+vTf/W
NgQsMRRW+0JBdzL54VFlZRsgf/ni07MTQxUWWTMPlcaAiia4gf3eDBG6dXB5
EH0oyEqIGfPMUFbCi8f+SShDh7ijgEES628pT088SzLRvAOhWcwjIOv8VHDO
T2R3MysYEV7rhg3R2WVFIHMjo2SbJE4DSVjIF81soOg/W9m9xWkNFkn54BCj
vlUiqW744Sa4r0qqCcWfL1Nj+UT61rihZKUb8B2OZzxJL0sRHdFIMUGrKew6
XMqm4WITNWFOcdHmCnMW/CREUAenzLxACtVDxuBXJzsxUsoHhK9RsUPuumeJ
gdiCX8T/R6xTwdO4ye7u7H6r5mbDxom2ogU2IkOOULXXUhcOeFjft/ZrX6i3
PM+PVltIFyaGIho9QvJQZNLfdruJb0t9WTG8PBsajvzh1GJhyZhsrgvkRVa1
0VkLimmcyJQuUcPzs/FJZ/hoZ7ZDQ7fBVnpM1sVrpnfw87VkoNjs/51D7WGV
wezGnuT5G+3AuX5ZI25MFYd5DzjMJURwrmI4Csmcihhf5RGUCLrWGP/lZsOY
RBab6zxb2eCiUZ2w/JyTJPWCd4szZDfJa9ZK+ujuAO5z4xgAZpJjTVxWfTrv
aeMBPIA8z+o0gEgWqm5nRFOsafw9w4adWZw6Kg8K5soAMvrsNYQJAJyplV1e
9NCsI133SbY6VYy/30R9PkqoZiuog5nhr+p2RvpYGL0/+p6rROo+4n3myUP1
xZLFHYlpN0H3+bIX7iS/xBVDR9TqL8GVawJ566QLU3tOYJQSVqvMVFpNClnZ
mmXDMecjnOVJFq0rKc67Iuo2fQQvWKAhoTTZMy9xwoes9S6PiVvH4iXTFIoJ
dWpYBrfBM8G1VdZCOn9z5oOu9dx60gmuoAkjxM8JZrZy7vcDXJqW++Hnal5p
sDPn5vcQqaIz37vq/FvvlWsz33XVkE2p3O5MDs2CZSqR9tsK8d94z7wrbi3F
2dFZ/uVgMX6ub7gDIKQoKA2ipMXYEu5EsYAG0Q4SV5A3fzVkN7lolgnYMyU2
DtRNltZH2kfnznGAT+bw+prtBac6JzEGd2VxXvW0TvnGhXxz2lLtdivyKCjT
D6yIV6ekJj2vKGJwEZz6Bg6m2Eahl5tN4LP5VeJq96LL1wg7luWSm42rVvLL
QJlwfKnFsyQorKS4tsJL+V6NiZfNUDsF7AVJIKJvZ5OIiU1Tp8UrAQE99xMN
mcZGpHLdh6a6AatOZibz7bCGxf5m5FHIdj2bA1ItpznyfDZsyqEVbsM7vVE6
yopzY4XAY1rsO3P73taxVS35qeuavSeC2Ea7kPcFlTUSlED1ZOHrD/6+bQ9/
EUYtP7btCsDpFnkfgPighSerYCr/DRXTDza3xuhnRXWZ4dQcZfYr/QL4G4Be
Le+eqd4Nq7TPwQPwWAWYZUaKqxQG7RhFztQbbsojrMSozvUpGpqRq2ku5Dwe
3ZqNoX+FytB2cmKgJRyzVrawLZdjPjPDZckgO32vWwxu8OqbNcZg1DcLYuYa
oJz1G/JuC5wPBqWA6hxmIzkKp+uJJPZY8GOE9afIcvz1psujZFruSB7c9aSJ
slgg6OdIJcZ1CfO5XjfEwvtYVELZzvRurd6v6T0vkccTcHkb6vFr/qjWVSdJ
azw037j6pl0s/EhXVCswGknYk/TAQe8JjJ9DWNgPyvSJsn9tiJ/a92FobOgD
sSc84BddU+8lO35NiZ9iWnxCVF+1KPuRCAyoTDjlNVFembkSV27p4/0hf+yy
MxKw70qs3synWsCAMk9P39UM6XQyRUpGBU4PedR4Tf+rxZ7EpGXOiab03LDS
a4Gm/WGaINKaY6A2VANa18MHQCUNG84GyLCY+FIo9tZiSzgC8jikTrGsUxCz
4sLeMHqDwe5uzaVUMM3gNmQgyvhwFf82AKE9RSv9BpwFml9fDZ83+h5qdX0a
tKj8lrO6+PBQC1r7c4iVizy9TrHVysPdFye7c1XcB/BPrQnzoEUJZ+1O4fte
K+2F5josioLTJSygHQht3SAjFXQ3FsQwReQGU3gpYVxZrPgFA83hnAXXvByR
1JnSj1gFtzgwokzzB8J50d7Q/2Wd2Gc8ETgqbkNTC3hfN4NsvjAmI3U0i2OQ
e8WRCdjiQ+kkUNr/ty6nC+4FKh+5vkqlsnlZBbFgYYS9cr0q8xs6hRpcK+2o
bNCCh9q/Hij3sOe1sF8w9XiV0lZGboqQSlmOuYnWVumC9s1dZeS7qz15hJi+
6+/OKFtcN5IltgBPe+HQoi3INGzGSVJhTistqGOZeBFwwuSb89DLd9JGD1J0
UAeDyE4D72Ycx0zIFX7jEM/fsnfuFmwroMGhRGSDKudpoTEV51D+VY1H442Y
i57IP6LZ/39uHaQ/sRmWe4rYu028z5qfcEQsmN4d/GJfs2ptIIMLNY53Hsjx
sOso5jprvbHJA7Z9cZkBXfi6vqzYS+mqyDS581rHGslsJtSdZ7vSOvoaBlZI
etQRkAXaho506T0CFh70WVoBOQNvhy4PwcimaPsmjMWTykvAhsduWeWw5saE
LOKbpp1M9MxUbH/q85q51cCHqGE/z+rYcVHnYm7ay4Ybj9LXLnSmH5o/lUCK
1eqyMlJnaEYF55yPHabb143vmqt+2AhXmwQcj6ViIFZNpDWcweMS2D4Wy7RA
k63zdgfRZvLvFEioRkwmOQ2JmR2jvW9vyX/0aKiXLkGgwRKb/V0xGnPHxLf6
MlpdzQFLiRFQuEeG4kXQ7yMdwBXqmzZLLN06Proyw8WEOyvAqzNT9GjYOtK1
OnF52ZBb/IbAj4QP32+hLK1qZKiXK1janNORLqJO9rIZZRPJrnLnUeWd7tL0
pWuIr5gEeVmMMKlNZnB+CbWydf6tZ4HMK9N5JdyLlwv5zD1UG+W3wk9LTm8W
taT0QAK3Y46ht+7Q+K3d49QazjBI6jpr5MvnaDRyzO6BZajLFDrbSK9aPmD3
PbEqoNoNEWsK+Ov46dIXNG2+9krbqEJQ5gJrXym3dwdv/EqxJfCHQNmJdNvP
WB5KSUcHLYemW/BIBQBEYNV+qQ3+Vs5P8BE8AbSe1vr+etdtKGfopBSStiDO
I/643y/ZnOkD8mbaB0csl+JTmIV5dS4ZpL/RD2MjF6tG9uHY1xE+cgKPvbJV
+L9dA0GqJ/jftRJIOKvyp1rHRyiEzVDoAVZukPoXFGDmpHjeGjH9f3EPq+MA
D9qro1E4x61TBM8+pE322q0r5T+rHCe5HxSIfaT+mREaOLheTnlQSCDzrz3A
MLTDa5tb6Pn/g8GmUkpw99WYZpbPwAHD55TSFpj3e/HiZa4sWXfas5kEFThm
JhS+C5W36rXBbU5XZcYQOnoQTAghstsiJ2CSLFqak9EbGVaBwmC1JrtoGZG9
khle9De6LYb8ZLhD4uMxlk3f1QHKYPDL4qH26ch6aHFBaBwy0wUUhEyzq9Ij
5a2eHcAQa38wKpk59a8ZJhraeF3+cieqdOtW05YqasrHYd3KNRBTonqut5TX
6dQ+R+SMXFa2yj1WuAP4qNINFARaGtfcG/w03aKh2QVF3qil43Oh7rXmCLsk
GxGSziicnHc2qF/5dND7YYFBkH07TmpboKNKE96bPBwh5Wo5hkg6UBTEs+b8
FMlYWygC+Hj0i8U6B8W/0PvmNtd4lTWWQ/jDvNzgaCRkLQsavJ3aP5pvKqUj
9AvVPZ7QovHweCXt9jJzSqzQ7BHaZelPD3abeYqm2hPWFApTOICqMB4f8Q/t
i6dwQdKjnLLEgvnkiyEsOTPpKUfUwGnP7E2PJrSQWrFPSsB5HIxnq78FIJwH
RAXtKDJOkAeYx4a6jHgtgWJdVtxQhyxbqssx5bYWl5VfR3feYjI4yQkCkgkL
LPFEUKRN7KFd1cp3fRdQTdC1gg37h8P89UfxI90gbsKcdOB8smM73XaHi+NX
/ZrKPlC6Ak9jmveH5QawjsYN26Ql7WSxMm5CEcA6rJyb8dD6dIiqLYq5Xkal
65h6zLL7Q6ded5x2VendDeyn8la5G3f+Bc9XEkE3YPLtmMTKEqqwx2v+dfcN
tbv/hq5cz3fKQfiJGMLS5P0dwAmJaYXg6cPh4o49k1WPNMEe0csGEj1SlqV7
c38Iu8I2tetNy0hbafdt3G1yzotJvnRz0dJpFklbB5OrcCA/KaammBXc2Xlv
bo4EAF6m/VKZgfqS5nW2P8h5Idmbfw3oUmyBzRztgyjIr6SNYU6DmOdI3Ynq
ZjMn4QWq/ZXAZi+4mwJ0hDawgs2LivmA58QLu6C1naMQSYuHrKY2ZwUHx/BV
1uqCQb93jmncNhVfdcbSVmnTyHhB20hzcWu6I9w7WmVGJ5N+m7QhiIDthLAz
u//hweQUm/9XGSXXffifpBGdv9Up+LmCi7+qE9is19G3nkKhsakmpHrISS+4
Dw1ZHEbb5ZApPPCNCR6XPMUKllQHWF1TXCjT3cr0+Mk1IVICS+jRsgNwISzF
pjvDFFNYuJvc9QC25kJNiz/+oLLtWiNqzdJeYqbyzBuVH+knA1D1rJg3t+gq
nfmm3924o488w3CtGjmiJw+ASwU17xdw8tDqwUMF8KUDdbx9VKYeAngfJtGu
ff9v90yegsfy4ISlTXp666EDeMDGOSbcqfWdKHiRXZ/TYEDSUR5Q1fmg5t9n
iYYpNPRUaG65lhaNXmbe2oLFLN7yxVBZ7qXRSQVRB7RQROwDT2fD4NeVl7zu
P7kIggFwYaeIYogCkh0NCuy/b1zynIAxSxvhjvfkK3PVPl29PqDZeuU+iyV8
Gm5I/iZraEbeZfQtDO5AjvqPgMLTvogi2vkvC6m04xDrvekJtspY4zEFdPfN
7TZgkWSLuMxNCsxxpSb+C+9RnGpTxaPJoTKPPdv9dwyRqs7l2BUBMaWsxw/g
v+4ks+LrfeNl4LNyJKQKaUvu34AwI6D1LNkmYLhoGbsdAvwaipyfTe+jSh4J
uWjLROBXCnFyLrbWfAO+j3I+YpOvihO2BAvGycrWus3/Mrh01oMVOAIVEHb6
CrECrpNMzkKovynJgL6Xy5CmmBAZnERQ4WZqbZXIdFMrtHAkBaiTpTWv8G7Q
H2isL6ghCNTuk7mOFZf+8nl5gYK2ykKP/chNJ2pccoqbs5WFgsdxQI21tjnm
aT9cswFClTtn/aw2AO6XR8qZST8EmJxehZ+DWSMelGDUKGyfOkUTKtXJjove
H6cgCWdnWG/05J7lsIXLN6n2RVzrdlnp9IL8zpQJhgbFNml7J+d6NL+hQGGI
o4Te2MFbtO7vFnEz03AWcV2UQJJpkqU7Nvefi/TpxyaQ4XyHCHfVv70T/cX+
ummFYhOhfIt0vJvhq/TCcM7eUeA5qsL3EfzxnSj9m/rGQPo9veZRO1xPq2uD
NaMho+qrj5ZG0HiGG6nXc6yt2+YV58wCOFC3YLmSOYZSIUrdsviw08SNwTRe
R6F8MeJiLmJjdHgbw0bGrplHw5mrklbvbknhUMbgfCFIdcuTfE70RtFotl7O
7DmueepeAyxRlnFszNPW1YftTSaeSJ3NO3opH9potRkPgWtFWh8ZNcLi2y2v
mgVX0RfwyPuO5bOS6Qf8PPwzntIC0H1jBqyIIhkL3rCux20IJ1ukGpo7FQB1
z2Zgpzdd5JGU3mH8j0gZcZoEmIJ13JKzxJr4lq3HDYoJupF74F5sOfj+DqYy
+uaOjEQtv+XifccTYihSSgnmvUFv1YBucltypc//1+kKEk1rjv3fUD+jlpi6
Skjvuk9K28404UkdhCudBdOmSUSSmfjVWMKvq5JZ2SWXLPHSjvwyURQDYX+x
fHN7uDromDdiQuQG4hQ+1MglG/9q1Rv3cZiJ1XiKWCbkZw/zLTSZNuk5Cstf
3ng76XSbIszzr+wGqo5qifMnGKpPefRP9bt9z8fbpErMI3KM00ICppt3nf4O
x1omL6R20e4uS72OrBSQBaME8p3STiTKO6LLUCrOFTJihjmub+QnJ5iEFpG1
gyO7DEWv+LuHEEoZQOukNydntfv5rqTRpv3Nz6EMqAhgGOFopzwZDCLlFMA4
N10mozWV2Mi+2MZR0tpiNzEBIIFkbYKN4eUbQaDuZY9v/RVYhfsMLpxPHsbb
hvdGodhyrJHtqWrlmCmvptGsiLvuM0TQ5Ob2X26FxsxdfAnd+j1CASlDe7xR
qyNp9piIaI4k/wtjaRL3Xq/2B9d2KlffN3ij16hs89EO5Rb9eAJEykpxLESp
DUjVchjYAb+HXGbKtpB2MFBV9VpN5XI/qo/AkEyJFOzhRwPpK5xAMQ5nWbEs
ihw8uwx0VOhqDl8i2V/XNYrYBn06Vm1M0KWABX6d9zZN+R2RJdVSUbcgYpAB
umVA7VBUCF2vBme9AZX55v0I2zs1uuyWTCMxNP/a7KbqK47NHsKlPAZUW8L5
ivgqmUu5BRCLlcgqIaeY5y6x8s9cE4KxXm/mmRs4OyXlMgQ6VEAUASfWP0Lz
Q3pmIB9TeU/ACCTyLMPCjxU96BvNbxlHY5Q/XXOsXDV30P7AAfMBBKC2nL7Y
rrQy51qID72jaKNRA08EaaASzDHii/7Pg7sGAmaaQoMUuBq7A3lyg0AxDH4S
Uz25V+9qiWrYv5k+3UpTablctXi3GUSdXS5eHYCp1FZAcZb71ejKJBLd0fZY
FuMCISWxu1d8BkbQyWlcOadQkw3qUt7r/JPrplHZ+n4L2DXeTmbu0Qd1NEOq
rfq9MAhWmXp7u4VpwU/TkQ6EUZueB2iEz0FJ6+wsmXLlYHA64eEot4Xj014n
yNW1h/CN2VTnhRsNPzYx0/WC7/I4y/9e5ktM7LsOKeBaHrlCUYfkm/iVsASd
KIcEOWXUBoNih5cYX867GSZRTnaRy9nkh9JRBtDOwzHwpF8tzJaoybtyNkVM
G4A2TVkMuO2b8xx02sCvM9vbs4bF2ZKT943hRcF2JAtZ4RwOFJAdYHhrGobD
S4+zR/jpKpm6O+xLRJiqP6XoPbgtFT6otSh4IjcNthfORRZqG+Wv/Jf9ks/A
0jupKNo/0lO6L4BD5a30WILXRDpnrSWKsdJnxN6NFwEI/mbEeLD3S2Cd+Kqe
8xr96K/fDGJ0wNcqZPcYLdacRnobTvARuECUlKmyRTk5NbN96q8Yo98ZhYuc
gZ1NiiIyIcWs/++UTaYShLbsG95Py342xc1G5PKF44nhGjhFbPr+IvsrfDge
IAry2wzmHvQYek47wYUhgenbt3vbNkpp8B/EtOVZv1inXyTepQom3shD8zh1
jl9skIY8mKCz6YXVY2pcX+33gaxIfaDGPu51rYKmbZfH40jSzk2fPscFXa4Y
u7431Sg7rL4zgveuD/xBfbTY0Dm/F5WDS7pMVDUl8vVEa9qjdM1bk+VhljSN
1XI3haL8SZZT2X05XApdGWJTf3xtUvVF3z7Kaea/gnpUhGNT98zcLxUkJtWI
MyXRJv4Ih00qkC/oCX+GP2EFo7WPo15fBz3d9knut3opvcSyG3zME/UNS3Zp
NlTBQKHa4G6Gz1yRb6F1Fpaf9uau1IruQX2dWQi76UNnGr+h0WUlIl9aFck8
DoXm9rr1LnAS2G1zir+t4MFzuGTW/9wXWdBGb0FZSfV418ZNvOIuLP5KfSEs
+/GIVwTLHwutHfmyHrW2Z8tRL4HOLU+WzJgBXXHmPErFl3wz6kPDga6NdS4d
KBSpLX6byHnZLb1NUvKw2A/V3blhHAW8FPDt9MluX/bksvYiSs9pEbXf0/Ov
0HJPhWJnbH59jqS8EoKYPQwoW64EFvwcASpDYf8+Jiy5UnSeSV5V625dw/JH
6V/957irSHBvsIoAQDaRuctLMqacrnlQiA2VzgciWKMW3kw56tEAfalH3MZD
/R4bVZnwQsTYSPh89ZVO3i42O+wrwo2uno62zYHPbENWfi9p0mdrGZkNiEzn
tsbd5JPywKD4HemqlcKdSq52kwIBr7a+Km8XXHAyqp+UateYzq1EaQyoXe99
biVCdELt0ISjqk+Fy/mkdi2k58vgkLG4U+quKb1NPJXo7ywqO8WEpf+ZqNHO
JdT2KyI0aM1pgL2chQSBRIQhuvqww0SWxFlvHnTbTYKngrhQMA2iypUcHY84
7SEM8oaMZXlg+if6dxVkkRttQ6GxIUav2RCUH+HsqIftFtrj1S5EO1jJdGHf
KN+uhCScd4I6RH2SX6v8UMTSB9/rWoTpTCpaapSqwK04Jidq/a3DtcpChuhE
V3DM9lxO1qo9nZQZOd41KlZjfE45UCAPHTVZ+NfDQOrch5AlgtV8MlNJvECQ
e41C7eU8ZBv8YeZHw4dWIjD887Pu0Hfj3jsjWOsuP9tHqt7G/N+jvJE7IIH3
7k00elGKiGjscPvuBASbjarx6bwii7TjALEjmS/x3q541COfqBZzdyaZgvUd
Gcfel2cDsAz/f3PEXGiM4JpoS77xDgysXoi7oxFZ+s8rZGfv2qv6hKOR3Lpx
aRPyHszZjBmnX+UjmdjpD04u6coeof+Fp9GOPGPm1F1Q2ZKBdF1e8o+6aT58
g3qoAfIJmOaQtncLoLcCV2wUDOdUgV6lxkGJQG9Cc684A2te8tc0ouR8gHnP
f6d5tVxVC+OejoqSpRaShx7TgYBENf0P83pn0QVnRvxWp0NhH3Z+mWEAQEHM
oBJ2cy16OVUeGGxHKaxHV+YDHKw5TLdMGbdEoItwkTZ8tl7IwYUYwkXLcMhs
guXTAdELua05ElWQQLbU/NnvfgW4YIRDnnnGUwNyBtkBML5z5CY0x+p30SL7
LA0ahg0l9+xbnZ8moI6o+PznGVWQSA7UkiKvcicn2K72hdBNgu8QFzKYwJY/
fegcLdvOwMI0P264MHOGT9M3uLTBK9cFTP3+md8WVqpzGibLUyudzb8gpgGk
Bc4sg8bC+MYR60OkWnU8bKpKeAgGkEdU5ksa3sI91TlUqp8FZ4XBAoUiNcdK
jko+2FQaAKFszmT7c7tt9YDiHXariMWldETFZaaA6+wSWkpEvciuUn+rkIhr
b65mhdgMLmMQSgfIJ4RsyqzAgsBQOdq4g0FeWs5PjPq18SovNyS6kAUw5EJM
Mo/kWz7Ygrvsf/eYxYhcGFeaQZzM9jE8UNNC5UXcwkthRnUaq+V7xHEIWl9N
Y3hnhaFeEiFncdZwGK85q1dj/6ACDRycAPMZtoKDqrRoxmmb5q3oFGVP3hC7
KVWq3WtcHQ5ZPN21H4fFRxV+2yx8I5JpHJ4/YqoicuYp6xD2YPGG3f4k9QGp
ao4QPrspuiBvtU1IY93tc4x16q1+XSuH0tl7tG34YidmAYhfuit69VUxPFiR
EuPA5d+wEFIAWhCH5u51gHkhDZhK/Nltlvf9i7bLV/acMIdAIBhISQSZqcbR
go7funL4/Flh6MEnqdHyMVJoKH30Fi0k7YkeeNo1f5W8zANBp8iypzoWes9v
zWTZpFjRCpSWjEHJvhwpQd3CQGjNDDR2RUUor81C9NDwYc+jvA+ctxMw0n/t
q6TTnnplC/6zA/tk6jry/VVis1pGxpo/h+tHemTOPM1NfvyJLN/aSGKx+W33
HgQwHLPDhE6qgTjtNwNFPFRNUB35CrxIVjlqy9ueZ6gjRskeQE0E6X2+rlKZ
cC3ryKGL0G4tvTsgCbcHYDpwyw1B1Ay7Of8eiEyFYV1wgA5osnKWcBSWPAUT
mPeUbOrplzlt335YB76ZL2o1T24ZGQ3vIYhZCzqzs12RadSiJxq+N3M0JD19
fEGzzddvCx/AYKGkqY9WL2ynhKKMk16u+dcoYJptenBUB9aBPE+zCRnVJ/iZ
Nuf6QK33obv6nYTh6U4C4HpvpVYdhKF3nlS+XTNXJ5wY0vdUboNQAYlKRGN4
AV9xWVSgR6OfU9E1X4mTdsld8eRp1z8SWvJVJS4UR9Xr0Vc+uSUn64S6Oye1
GuHfBsnH+eS++O5eUCKwpCWOi9mWRdBnUYakLk+bxtdkszuO1oyqKUXvUnIQ
igAVR5uvl1J+McnBi0fArOoq2Pf56apefIv3/ddnXSYjir89qixJgS9GH9BU
OLKag4ULVzJQbYKUlIv5EaPESxHE3wB8c3paC+55XHvurosq+Fdh69nn8gW0
I1YLtUQgXsJbBPwmiSwravxus1cTb3VszxD+nd3nfVBtCwaYqII9lX8qserq
bfB+1tkxHK7r8sVcMzWZnb4uI/2PJE3gaA04m9f0PIJBLeZ/k1Lnjex+iAqN
aChT2+cBYdLlajeM7QwWHPPRKcPYJl54OxH7BiecEWqq5WGx5ZCzyyEO30Ag
B5NMzKs+IdtQzRX1OVBz8GY2DgleTkr5mKk774XODH3V7R7HmklZ82sMRiGE
T7yjYHjWoFiE+zBnpn2GqUcNcjgILpeZQMreVckT1x9jubPqHQxBDgNEJTW2
Pir8mf65/YEoEinE9CmYRGRX7fuiIWJHE14oPMWLYVGcte76mM5nbRfC1MRa
OE5YPKoYIH7ww8gC7qBodCqDivJOCtLNToU/87iBiRCyxP5PbfMHtd3OEkmX
PrRG84ia/RKkS6EotETZsIJz7HUkzH4G5qiiyl78MVyZviJq8GKTcwMgcbJ5
liBGCqim9Cc1WEENXACOyI7QMC2CgVAxErXcE9gowZk25pHW5uxjEOsOQdK+
d1zWiTJZamS/c8v9fdHp7c6iSXnQXGeAQ4Zk4V+40szfpqWBMkERtJ1yHC0Y
Nm2g0j6qcrqO9XCrDMsNz1+gVQIueALk9QnRLimbFszvJY1izpwwo09Czxev
TYud8AJdvsnDXXo86PgkQItOqmSi9r2BMJ6LfzzDF6r62L7r1LkgKzzfxujy
F73+i+KdCGfZ+nRc9GJNIV9Q7OaBAoPTPWRA0f4zlqaOllLGcqt2cNl1JnFs
QOq92ZoZznS/kg618vN+F3YUqP35rsf9FdiXXqaWu7NHWcQumuY8WWs8FuKh
pIlTpHbsQnBVfX4vxw3KG6y9sl46zGzkzKHoKdypHNJoTm29kDTfUStrdsWq
fzNTfjpl+zbt0XMpSKlG5vVdLfdlYL8wbgavCBTjL/34EY+zfB/PdA8EtYjm
66KlZtDrcvmbFlBm22OQ0o1o3buW8YY9qm3QJXR+5aH4HYKSxJ5oVQ8WJPA7
tnPK7YK3yUJb/W+3YuSHlv9J3ILwN23LynDlXqmWS9/zRSTKCK+Lj2yOt1VI
gHKbCSiWgpddZiedCoKLeL58iE/wwUeLIeh7BwIAghUmSQjAa+epDGSKxCnH
Nz0U6p7darKiGCIcbQDT4v/NRx71nObMMIokJkr92145yuMOypMxVKtTiRHw
F7jdred256zOQhEkM8LVmc0SMRudyFfAqp1unCZgn8+TOozOrv+++PZoY2yh
Fo7vFOQ6VJ9xpK2cMl+Fb4rpLm0ZsNL6ayNFfQ/i/QZKIGSL3RTlTSDuh0On
6ISpLccDTeuKfErruIT2v/O66JxsIcdkjpckWTtUoVkM+xt/laCvSq8qv4/S
ydjhF0Ux3HNeH0rwA9raxilkAhreScbW8EbEMlqMsT+ndKm9KBW4qtHDBD55
4ROStmRQBEbvZLpbb7hhS4qPez9xDijAisnTmZbts8x7o5UUscp21+bkaBs5
oFi/ZghtiZbjxVjJ1utC5HOwbh+LZwLA91EPDcfq80vg1Lbc6jDfgoWYgb9K
jCANBCaxBpPT61IXYNWydT84ZBVP9U9j9/Vix0FHPUGU1gJVBp7VjdClYcj6
oo/0SszNCDqo2gsQzKz8HSfjbY03qffObRqSE8oTjn1eHxALRTdQrp8X/dB/
sLlC4n4BgjA14+XxFcHkUA702zCNStcaHlxUUgXyAudyjn0BWn3xtgn3TOkJ
C4YOcDlscwAg4OffSKnGZDtj58sFNFJMttyNppn+56Qz+AIoUDMHe+Ub13ce
DRZMb694i4KrkMeYahhA7yUB82xhKTdrATI+2Ue0wf+iA6uArEKM6Wsm5s8a
+Dn0FNZ7G5AtPBCFS85npIzY0NHhzyUvYXbSwqeO1T0vTQozP8hlvckUd3Np
NMFP7Cj4IFRzUY7ZWRBLXy743EA1337yeEIW7RepIO2O+Nnk7yEvnLNGkwpq
x/daZsld5uY+TLvONh7OFuq0YEyVQAnVcQ7ysRB2Meug+vZi3w7Ps2wGZQXe
VFtmMxQOu8RAsfXi11bn51KRuPJIpmFnkL8o7JqS/mbJN/PArEJZHCJdalCh
r9DlAsSgRPTqQ39jdRyQ99LwplTnX5aLN7CA0d+oP6wPRRT8HVKyP8m9YqWB
L1AMtig+HLeNO64Alo1Fmx3VJBx/7s6av3QBoGWKHZ6pOrgj8ZLE+AN7GrvO
pK+GQX5ztuk8MzmjBq0kvIxyN1JxS37AVRU4It6WaCvMJvFIztLt5W8Nnzq4
ZXx+AF9MRRywDumwWHF7wwIFNTtBzUuBMvhW7+KhEuYgpNt8CASZ1Gn5vk4v
uLJCyANZVfNbcMZieE83L2jqHw1N5icYhjdRWQHmS+xxrDSd7rN32L7uccxB
Clw5ZHWFYtWfrLFvH5peFkJkarg5OSYhf8kx16VO93Zg2r5zDbHZ+Si3QD+7
0oBtha0zxPrniMGEO8WJ2TxNU3I9PFETF4tFtxCwT8v2wNHW6rcejM2iCAoC
cYQcsDJp83D0jhc6POj6SEcj5wI+NE3xUJR7cKux+n9aF1vJmJXzXzQB2Rms
iyYChQ6rCC7aFvphj0tAhsu7gmONsTQIS8h7Jk3MXfw48RxfGhzW5jN6kIHw
fZ4ReTmDuWlRXMjt07xg4n+kq9Fs5+HCgXyahpd2pocHBt5dbEnQ59s0eJMg
aM1ZhQEznUmpf/nbApCPojb3FyHZYE5FS2H9Soc4b29fuJkt0a0g8/5gE79f
k0y9BdvF2gD0MQujqYOd0qrFQFgRVGFhHUtSML0GQytO33FYf0wOPxB1Z1Qz
E3JZ7utrtlbjBrZQUpSdTARGgYcj1n3XmB77nfP7s31tVVN1vguVaVs1mSvl
PS1Ru6aBfP7s+pSTzt9mg9Zoi1gh3jV/Lf96z1p/6rxiMqaMSUyg3AxtP9W5
S3aIqYpsOZPD/6SRRTbLJH55TzJ2TK2Vi2YH+7JZkxmBvBJMnaT1XZJTi6E2
nQp9o2LvoBeht7mE6/DYgIIaJaVrCSf5isjL9fUHuxcyOWnGDRDJSwALN50M
4FUEjiFeq49Y/bdCEJJTahHKYcCqmg81QzbSeKnTRoD8M9FpW2WbLkSCLE8u
OcUGKZ7OSFx9faIncxKvwutSenMxEOod5hY0pSpW5DTT4ihhOIvcAxXrmPeO
984+3dcHw3EImwq6zpRDwx4NPSg4K5KtSZ9lsRGt7Xjlnmaj/P6qoYp4xeAe
EFVGlSOZQT82L6Pucs/G6x7ePOzE/+lgLjRqenCLERrZ6a8pcWhWoUtKYmfb
9FR4xyoILmSiV5BiR1Jn2B+De32RWV8S1h5wFsq2r6F7j4YtbkYlHEaz+FZj
W3hOm/OQQisN2iOLHid5SSLC4fNi1qGYf/aK60Yv2fp3xP3ZMW27O96wlfu3
ZtJ5SIYVXMBCZpn+xGOLcFrL8VH5Fek5WbJoJ3WdrAMWc2SC4GZuH2o59ybc
vTSeM8taBi19h554pAEYuq2wOiX2vaw73L9hGkYXaQ+7C8pCKK/hgT/1pSwP
ORlzfPlCzHY8oDjwoJk44L8jbPuRYhz6HxYgRgYhgjvO7KD41wpJRr3mGe2v
H/9VKY/5x1w6iri0zYrGpslW1BCaz+PwElObu6rA9M6pmaZ82zMC9HihSI4N
TyrrfYhDu3qTvwIaVGuBlYvzRr18QUa2UnjAgxuFI8ky6ACPQfEan0bWw5rX
RooLY0gq5TyS5ai+7zdI8yeTAnl+j8AWpucuDFUJaWKQRCtDT70FS+d1OQnm
39/2gFquSryAy6LkRR/d/mTYU00+eyGivLbZwxhCccOtxGz7eUU2d5wyWiig
t/Uflke18P35+hc/RMZtd2c5JHa4xxjJsvGycdSIbdnHBVTV02pYNNOAhbXp
xqOyqr8U/MjPJ1TCm9d9QxhYK8crb6BvBcChVXyAZncMfSI4+isdkmwsmF25
dLFGdaz2kyGivYarlDMMA8UL4yYUldeuWBgYmENaaIP//RLHDOubWYwtp0Cv
rF+9hnyop4yWTAhInrPLGwkaRbjY6qcp8OaVVgWJifIT/dzIXeVBs+LzajDZ
bjQaDOcgeMdUCflV8RQV7rrExO41yud4GxfyySVSt//p4jrHzHNP2/QXYkZ9
s3hKBDGaitR0RdROzb5Vb7F9ekzhvd/aIGIRrnf8yUYpu5aYNGcRUCNzmJlm
14FVpIcUAuxk3zd4Rzx8vr4+u3hgIIKAklF3TY6Jc6MAsEYp37aYmRz1x7Dc
MmwaF17xcq+BlPbQFhFw0aUoWbXLPH8ICwggvMS0CyogRhEFjT4ji56BHgtN
e9ir8CybAiI0Sn8rfEvWTwd/NRKL8L/Z5G3revb9pQFbzPDuDxtxL6mTCLf9
0adnS8hQef8zSMTxvHTHMAPUT+DzxOxSfR4ZqqLkqELJDhZ7FPM/R2vqo2iz
hvJC3rFxGA9wDRu/DobxhgYaqBZYx8+GyyyxSEggxIDmlIxBnxU8wuDgHRYB
ta/4XAaASEe0i+1Onx350Lyre3OxM5d3I1kRF4/fOGhWEegKpHiH7APVb3X+
tKTi4BfXCWAB4QN8KIv3EjJtvDAawIGXyXWN746cmp3RO5NpVR/yOXnYwYSx
0FXawoWhiTPeKgWNaIacbOZcbER/s9tEUCW64iVmtEvmHuD3dWJ9Osr0jqhO
WnW73uguPTlGXExrpDT81ME8nPXEJBvt2eUtuBNmD4UYggC3eDn2yHlZhDhn
czR/BIMtq//Ul0p0+oaMDkhKHNwGLw5KFLWcm5GecVe+XPdc2VyNhDFyB/0r
+XAGMXFVwQ68MmaucYYW5JfyCbyHTICVU0CF2rWwnu6fCbHJFmjwlJossyHC
blXCeZRg9Tt9E3qOJ7Yv/nN0X9MkEOyiuK4gulCgolZWGaeNVOg+ZWT2rQs7
rc8WExiy04VJxI0EMz16RakADNnCe5a8CKuKv6NU+uf7HieSKxY9lRhqXvpy
7N6KZwj+HgLekLymSUNRrkl6BIdJGIa3tfZEtI2DPMy/UW48DsPALFjm5edO
nPjVF19QEzy5+L0c1oFxvvuxmZ96hCtxy8vrdau8GkHvFD9zdkHReRfDZVwQ
Kqpt55GkHOoZCqt+IAMdqYrDy2x9YbH1CWI7GeGLOJarO27U8s3MR0FkK8WR
cPIV9cCh/oOigtSbfTxpBojSY+w9HINOiNUceLZjMMAFtEMoWiN3oP1v4uhe
Qh58LZfBY+S37gUDfaUeRFBxdPHAKVv4t9A6oGe7h6BtkJx6nNjqA5YuwBUP
y7fwIipn4eWl8iJsnPH1m3thSZ9LR5yxRfqIy4+AvmWyIUFeBAJqSyTJ18pN
04D6smWUiM4JBS29TiYNxdnnagZxxzzSg5mNls3UZcptnX0o2Rpw9EQYuvxN
tRpTXP0p6z8r8xvujsw9y3wMvxRvTLUl/jHMg3gPMCILVMhccIzUcVxAaj/a
cqLOAA6j2AkNZSS5UOc4D6vuB+aGeXFO800cTvXgL34qjIXbRc+fLnK/nqQM
kb7snNl8vZmfGUMpxFpM0OTEP9XU2MkllS3VEAyNWox8Qk+vydIavOla3Cl5
tKrYQxnAkZT4fdrrys43/BSYoI6BZkZupt7FeK3N43YCy4QMwC77z4IeHEM6
wInImpRXg++wJhpF9OBNqHPiS15RvS8NzmFmEx/3tCEHb+fSSNjbztoHdoId
+VPil6LS7+OIXhJ4ybunEEskE6wdlEwzYgn3u13d4tVdr6QKJognAo28dAGq
I4UKLyvIMfKTsdR2ZkLiyaVFVnx+NGAI+nsDqEngi3LyuqPcFL6kl6+HpaMW
bDbcWS9FHz1fRgKREqxdFfpZ934rGZQF6doJC1OutdEKe8ajD6+P+j2ZBNl0
AAAuIi1YrswBwvUlrAnIvjmQ3QP6FOz35JF/Eulxrr2XK58OPL5KH8ie+zTG
PIiyq6WvoUYqvbfeAKMxdRPQIwrXVkZ4JTd+EoE19hsabAbDuSOz3TQFdygO
9gP87UtB/Zp4rM3l+gUJ76ttgsX2N0M+m5nHdO06eSwa60+olG4qEIZyEUAL
DbKrmJAXPPhjWKeat2ir1L3cv0jc9+F10GyFznaGstpQ887dJ6c0WVJlm3+N
WuCSdXCoIMtTXlprMC/awRTPjxvfamYnM5KfXWLfQX7t093KyiSwlksurAZn
s/ArjE1HI6AzDIrFrPnQ1Se+hyCysVSzb5U42IqNZXr9JBG6a41UbXb59Kw9
07r++OCf5adAUEpJuR1cOTsn5eAg8Pr4//dk6Sm89YWtNiarFOaklBhdmRjK
2wSPo3jKul8s0W0ems2xh2yE1xXH3726hFt7uUm9RG35XfzZxioyTo1Bhh5z
p88T4RjiEnZ8bp1OOJwGwAIkbOhgpUkVNzMBSipNSeVPorfeanx9wzVBb5Eg
ARLH3ZYZ378XlRzbYR7r6alC5XLeHAWw6f/oHCI8d6s67Rw17p+RDfbvFqoP
igeZPr9pCq5xa0bBa2+VwPfRMmzAtyzDS4FiRhezn97OoLeB7fMCQgwxxABE
F9QwYnKNXAEE3hjAqXuOcKVdmLTuNNYVjjUmH0d8bHnEn0sj9eVpn3QoIgAJ
B0FXCEln0zJMj/phNI2NtyyjIbXcoVk7rNjXQH1vPoJyBXFbYk0M8xo3V26M
v+WkI/S4c4YFrSCdkDbePaVMEoKNZyWGksnE3AT6RphGutPkVDqA2NlbwSiS
8M5/bMfYjijCp21PcU5dh3hL9wqFPgtHTpvjRKqyTdV/xAccCUjzFahUN4Q+
hQauLsR6Kio6Ah6io0korNwwzbGhIOq4kB05WH2SxMw7anoYtpM6ZekmBQ3D
BIqQ8nj/Wy3bITLV1GMpe7e63xQO+3KYPtCPduU7tcOXMJsV2TNw7olYqbm3
ndIb2qk3EZKqqGrR0B93juMMg0B8kjK+r+RHdvj/0p3aIB3aT9stoBwIYm6t
AVJNWlcohJ3OtKBOcjpQVrn1Lyg/OLR8W4+UF998hNIU4W1AQ56FjM6PJ54h
xCywa9vSe76m6HjZHjyCDeoMnCsbMde8O0H9nen8ggJ4hCl0M3cPz2yoHgBz
O/0FWmotYcTYHQMM8CSN5b6wL/d2pwrU21O9cxb18Wtl0CWKzTcMnqg9yQcw
QdD/8SI+yYh8wi8rq1a3rQxpuy2ZLr0yMeuPqVTYvb0DGvajg8LmcrrVd4+r
e68/5a4OT7dxWMAtW4Ak8dB+p/RCYm19d/3sG6GqmDgrLt/fRhJYCzr7sal2
DtLw4nrYBLZHjjfQVurGCZmP9q5LX7UzepftV/FCS76V9cftaZA0kdiYGMAH
kQ4WuIYx6Mlx/0m+0Nke7GQfTbAFACu4xXT7Jur4RA96hl68TRqXvE+IV9PR
HqN7FeT1bYGpTKuIB3EgNXbtIgXOdO48R7J1B0YcleStZKhZ+VeBjFSI9sDl
8/apG7M6wJuw7zz8CoVlsaAiALKdmnScQY+TkNLP2T6HSph/GYniPBlKxlb7
cRoUgV4lCnMQH6rynUcFPzvbQ8cLcQLVEcqSmwrcqx4/+kRXzyX+bIuNT3CY
sOT+xGHQSGUs8e1vvBB2Hk+PkTGs2e4msAU4f+l1yj/SrCQN8JLNk9bw/3lf
mOBCOI2L+FUP1T/ZV8dKIax3B98sDdWqKZ/uP5ZtN5R81Rk2N/S+xZj5gfl/
TY9CRWHsUU6ChozO9SStL4SWoX5TqQYCMYMxv5sEjvTtwRFGtnsIW60qhjRM
Sz6nykSAtXCJGjSNa0LLIHNAYahWXDi+Cm9j9zEQyxHCXFObWq+9LsQp77xs
04LvpQLuAozy3C98IbMUdu/UD5q9HMkalglWTYBxw2TZ/JsQOfISyWVjcd3f
mixa1/NR+HQ02UwH14P/rpfznj6HV4FoA0++Tgbom+7RYp+fvYdgDFITp82a
D4JjaYB31Iv6CGkH7oviyLvPnElQX3FFFXg45ciEpAy9wffyCTEDuVLKyJRt
XD8xz0/pco4EVsO0wxEjskIllbLrCoEiOR0S4NJGXiyj620aiVPBBeDk6JS1
U6ZImzO4DuGBipAEzzllopar55OpSa1g5yIx9Un+YcOHBiKah8v/egtaz8jM
HbmzDLIf3XisQuTibr+o7aiDlgxbMtTUJeHiLCtSdTFLGrtbjkgl9FMvGHyo
O/BQYUTP+cqXRNgHay/aTuG6x4m7d1Clg0zfpa6u8QLOxDVMFMHgT3Icps6x
3QCCMuY+d7zoMDdl7UFfUoN8AgOdgM5CkARlL3gEpAQFtiF8miztjbTHufZm
JkaQUt1RxIWwSuF/u0FmFoWHSitdpXC5OyRS3kbwj7nWawpWiUA+FaEuP+Ok
1KhMT+CHj/pWhPrkix0iWc9HMqbxbl3bQWFzpU2HqlC+ejDYlXPJhTRbe8Bx
arkrxKsFJURSDnu/jhSDSJtu0qGzzDzS4BQLAvP807KN4dUQpoFYLoGM0tw6
mrlevxFMVlPIKGqEYMIIn7rA892eLHuZLHsv5OhPeWjwFxhnJYg5NVEX2ZFq
0Ac41T6/cMY26tvxtia9teLPk3LwSKj87sS61JqgjRHgGbWzk/C9vNErUWmX
p3rc6VNdqGjOl32C640QUXW79bMwW4QnZrqe7GchMy0NacIo85xR8kqhTyAQ
nV4VDjuwoVLMVD5Z1Z65FgkixTd9r8BnBnMBpr6guoVRHgcVzsbWCpXSASmy
4Pr5NSrtPM+lCET5fGyxd6xQpJEv83yF4XG0bVq9ccaf8rM+pyPYzwW5FGxv
KaQyxWnKvFsgja73Jt7qOaj79ItlksT9e3sRx9L7ad0QfKA51oj09FF2nuZp
E/a3Fe7EXTUwGbuYaC3EoOAA9Pdnz2IsOaLjyM+xDPP5CHVk62HUGMXrnIVl
cNN0nHNIPHIYPP1KhV9XZPpqm2/r84VN0OYE5qiDhXoI/nqGhnsXoYtX4cag
jRuqTO9UfTiHq/YRDXGXM8Th0tP/uH9d7wLLzIupDz6EqW53/25Cuon5KstN
IlFDzsDnRlGpTQHmjPO1jJdqzC9wH2nSnrv5NpPl6VsZH8DovPF3bcAmGsFP
Qx7nLxDcAGhn3tvRUSzadyAVmEeyk44Gnr8x0hwvpdq94y11zXfa0H9tpCIW
FuIg9peX7V1bv46fG2BHti8TARIgsnBtOnS9to0WzojHghU3LJ77J0emPQEc
totnomfQxAwrh2o+P2t4s8k1g5FuaUr8ietxuAEpLRKEQgAPVbDDGbQhfQTZ
z7Qwt3NqGJNQb7Ud+nfbXoCspDz9gFCH6yfw114eU27YYuPlYvuaaZRXe4Xq
pgGstvDSzb+hQpQzh8Qj7n5towdDuhYTiaFVOOboYjTk18Sgyjj+A37bGERd
ATYa2UezPQBpagPcHjMpkZ+xvPoTsiualnG6xZyU+s06T7TW0aq79ktoMQgq
Q0Q1kX32ajf9f3I0L8N5YqF2mE8qhTdeB95pRUMiHEaQJAFHMi5ow8WlzSzg
CawcNcDiq4SfpHYKe310SEwx12Pe83FTRgR3zgmIMos6BA4cBVpY7vvycUeL
Med2Jzajyj8aPeP80fN7LyHtsKIledPOq/EH3yk2YREy2aAzCOrh1vorghkm
EpsmAWfHlnv5l6snr244wAG1RmxRZbJXjgD0rkPzo8ZggobnFs5ECfP/b6uI
WwJJRo+dJhl66RkmDbPS3t38gQzLWwu2wpCZT3WFLcWJvjYmoyrQoLZE2dt0
/lyM/Afb3aLjY+gtZWHeBuMhgA8C1WqU6sVmmLuBgXLsmsYyJuza85+v30Si
X0WFsn6ASHHzpDzNtHAxo9XEGTzlxft6dfmjeIC3jUg36KeTYfOoJWWuPA97
ZDmR+Q1Tvx5HhBIs2S35qpOyR/BakjNDMMEHKvHJpVq4YQiRxu3f04Eyj7vc
tzjEnKgGUL3D/Li1/CVLjYbUFEZLL18oSlAQts8NovY1xxg+i6CUb+Sx7tqP
TnIXdAX1/Ergx1MltO5cNgOsDHyRrt+cgkmu09wrXgd+ssTtgBPpvNq5vT1v
64wqDngRLcnBEjXMJaJBDM0fbo683TAFOdISQlEeGG1/hUyhq6xzqudJEW9X
PcdwBC0a+OpSvPTuljKT5U/Oytthhzp4bgdOE13jToWNEAt0fYgEXp6GwU3Z
NgyfW2GVf2GbSzykVdhG3cb4lsplK1FAAOygtE249sPKd/gCEwckfWFbYMrR
aysAUglbTWQhB9vMG8nCS1g3bK6IN67H2giQ0ErcDV96Pm5Bk2xZQBAlbdNr
30rUmHgQoY2hnMzTa71bnztmvbUMcDKzk1O6gJRaC+elRsi9CTLe8pABxq7j
DaXCdFKPJudwLJnURkoiyprOI7TKkRVq2n4bL3t1uPy5T+mUgX6KqwortJar
ZPlKt1D6v1wmSH3L4qoWXS02sXXRDfOegxsgULrB5votMjgkCzWouavnSCW3
YSyQn7ABrOcHwRwiYDH+NI139SnKfCQuH0TyGo8zXeNL9k36QpuW7Bzaj4e8
JXZYiQKc3JmsQ/D8OhCU+Wm7R3443ehHET5pPzpUGd5Qn+s7pkaVpDPKe0dS
9RFoNajtS/+1w6DqIwTtF9D+To90rYqVZTFyHa0mf3Q7+cbKNz46QjV2FBla
bRnprHSFXrMQpTCQwPDNyGLQgJE+Bft1asl5q+zNeLFMMszMVMEioxR9TAKl
S+s6rMTkTXX9gHqCP1Ul8xuC7l6Dp+dmvWGYJPRhF1CRHfpfOLShbIXct3Uw
NI54ju/OnGRRmD1brl4TsjKAtzPjKunY68zhnfxrP5TYUPY3J6LCPv5mV+tH
ED6cfDk5RLNmQlu8F3+8JIGu1lQLvXb3/kvsfvVMwM9x94wGdOMi0PIa2GK5
yKyBpyXL5hbQfAheurVuwM+ZYwbQqbHWmlbfixyWGHXNGPoAMP84EgWgDd98
cBJEzFZJrrbVLm5EQflo5KZC2zyOSfppIapv5t5T0oh33ue14YsmBvKJNooh
k3Pg8LHaBEQymdwmUjSUfCHKSwloQmv80l3Z64ZN8ZgJ7U6OUz0ArlKfn/q4
k2FxVFpotQDWCCOUObkRTrxl6OcvZeQMdOV9nyXQsHV9AGOUCbbW0ZN0k5Lu
OQJFbFyryBKnfCN1SL82l2L7HyOp7dXoUfnNCaq8dGZYecBc77zjqL6Viq9K
i5xPI8dJN0xJrPrkVwxLXuWS5yXsTZ1qBPOqjK4SZd5LgSTtehwE/ve7uDNi
sw+1uMm/Lc6mkwhVmYZyprvsJsr03LuVvZ7YNBKLiFq0RkDfU2kIJMqC0GFe
tWV3/1K8KjMMO/jtrE6tssCTiIp5PasTGVqwY5fZGObqEVAAB755E8otd4i8
U6z5550h1+81dxA0PQhp3f92vVDTFyrtL1HPygCONegFz/zq9dl9gxcbLAWq
VQawIml9rABJVVxBPlQZo0OV57oz6LFsClyy9gUvd0sjj/OytGsKKE0bDUN4
7qAIM08vIeut5v422gNJgxIq0tjPqdkABBxiJktfOQz/MUhfyDkgCaK8dMGv
QVVkSQmsJxmvNWhnPWUXwTBmcrNPNc5dbEluwCVFiBHJwyHOXBouEDqUJKXq
HS6Af5etC6ZO7F8Q150zzIyBKsL0RaXj3+W5Chdj7oN5Qy7VhZK5F8XkW0+M
4MmjMv+RUT1t4XUsPVH2njXU/SUFp7A81OH0ZI7vAEBMsJsQIRmGRROeiOv4
RvbGVSvUHXrdnS6FDiaZPIqD1KHWod+rKhzB8FrLYNtVbZOhF4KeUqux5dJS
PrTVopCnZpNs8RSXdipmZKXa9hj+UigMPJw445CATWfz0tptvJ6BfblZnX5U
wafChgXMZXAQBpogdXGCb3SA33/Q11wlj3SzD4a+bFDkHxyART7WGBp8teBf
QELmgigTrQO6h9mnwPUKwCKQnUljdNNrnF/7wpyGGBL01pAQY+/7Yy6pxVEj
+4KbF7ssK6CHIqNjwku/Lj6WTW25K8V+t4pVGfDHCHkVred7FHSDEbizWe5o
QVhQ8BArab+H3PjWa5dNwDK28VkDaPVlhsXdURiUzZrwLUeTu7Tn3k11/J3B
YRl9yIReln09k/YnPt6v0alF0tTSoHzDhDEYJngnvjSePbhrOmmzQAXiTtS0
ElxeybIBP6t+UwqY73E8/WdkER3tzcuIX40/filjrADsJ48eZD9Ej9OoGJ7I
SXKN4byCAtgHC3Y+rJap1hstfU150SJmAt9Qbd30Vm+OTX7NkOAlmuhh746K
YjtmK5iUaJvmFSDyjyffcSsbV9kq0TztIQpB3i2GfRJ+tRFddoMu1bNgoozp
WrNB8p+UThzWclU1wzbqFRtmrcbrpX+iTc35TBAPsqMwzkp10x9FNuSa1uLk
xq7vnq6qdlAszfthuHvpeQBmLeWXpw7XZGEPYRmVXu538BmXNI3C49HBiBWV
h4YZWlnTw6jdVLje3G7JEuOCOX4G1KSqJV8HoXVuFpg+xzTOH0yPiTNB/ZHk
Sl2gO4htF7BDcMrRPWL8EBeTBLrBWpTr2J8jaS1fOxH4MAqPMbwlfc8fXnxp
+OKqOJ7FAOgxRynjF+TGg7HFffdhSexBviUpNi26r1NOUNwlyWBLkOHULpds
VW5UHhpjpcYA7bhQSdcm4zJgjRMYbmfb7a7xS92QZdkzD+K43WQMvyMiXEU1
OWTWCl81smaJe4eDAQfKNPpmhSel4k5NWlvlW2X8xof2YCzKzxulppAj1e4S
nbOoYdPiZH2VDRn1aeVTrJ/p0l6cmVridWfeicckPXcM0Q5iZSuohlMWFK1C
iV7iUHTO2epjH3DZUpJ1UlNIHvcwgJ568GqBT8cplYMqHrordNUaopQJEeRv
7AmDgBMLTJ56g9+vn5UvuAhkKTign1lgPNJvg/uoLp0y7thrde02j9zk+1kG
dmiy3EqlfsDah8HYXcReFDaCLq7VlCe93BWF9RKa8uC5+sDrLErKdqPHH1zl
tBqteM+mgFZgadgguAocny8CoVzAFvyDDAigOgFDWiwHGl7MXy+XVEawpxBl
EfzpfsCM4aFZ6hfMN1KT3zuzcafGDCS76a5Y2Fkq8HJieLTgVNtMFhJMUSvG
frrnJKUZ/Y+76LZL7/hW6gpZfGkz1D2QbejaytTvK9lIYpBoME9TmgNAY5QE
8bG8o/WyLZZRPCjCCSAbb56PtRx/zrjUz4hEJU9MaDWqcKyer1Rm+JkSIBMO
JmUDd+kkuCzSGGDKXjLkFsFtdqI4B9qB1f9yCDXiq9q+YkRHpb+oN57qLcZh
9ukdPwSNOJSXLXpFoqVQdjycTgeg9fm2+tOxrK5446N8E44h0LRPlyr7HjAm
VHB5pitGEVqqfZnm6H4sFPB+UkeLTaZ2LF1/FFHZ3OXdJerVvguulic63+PJ
rIK61wdRTl5Pm+MuByFt7gfaXSMR3nrjzxToxaJWdIy444bNcObR001Uu+pS
BDcm2rSmltUdoprJEvM8KPRZMJw5ixowaEwA/ONNPGwTWq+AbbpJYvr8I475
lY0IZ8vp7siNdU4S2kRcSdzmDBvit62zMzoav+TqJJqEPKTMBMPqsKWBvjiy
EQn9opJHoIOTHI9tWZMQSa8/OElCXBaFzpbCQ6vxFBkJEEhXFw4dh9PrwcR2
eqmmWlSxyFvOpfnktnlGq5G1FG3Btmidd1h/8hpAs/ilrNPjZ+vo3ZhKuFlO
KMr+CWTNkZA9yzOxxAIMcaF9f6zGGS4Iaga9SI0gLGh0NcLLzbSEzPuCNnKR
rEsQTzB+ME5h0Xdy+cye8OkTSHXuJKgVjsLTP/l7K5iOgsuB/WcIxA34nSjo
gXHdWGRqGuGKtXgfiZ6mfStHFj6SAj33em0E7z9FukI0rWwMKX/VmIUDKe3X
HBNeIPeh8X6K8KPnJ8ca4OQGskEL/9DVveZ4H6YrZXIiMMa3ixbfU+WtOT2a
8OMiqX7fXOwsXLggXR/tnCIPQEqHDDXGLdiehGpugxwa1wu+MrlNnXeroafp
nnnBQHfCXkw79Eo4An3Mws2WYTrLJs8sN4izTaF8ojS4lCN+73bpekshYJ+m
mGUdb1xKbAxGQ1Y5pqtH6uIe8ROEdn7cpt7WR6LBx5/szGlI+yJOutuO94Jv
jUKF2z9v50pB1Yp+Acfh5j+WLoAcWEW6DnMaoT81v5M5xmneLKFxkxh2bULr
CTsM4s52ywDiHzckNaZhPK4mYEF3kPPKuLcEKaBSeBeuswQ8+3eAJEuiQ7Ro
wV0xfg4MESzwOvLAPUM2HaHV2bh7vOPpFJYV8pI1yqDC9Y79Y/aaz5PUfkuG
IFFU+KoPcuzoDoF0UGuX73/rKMxQCPqe3uCpGYgQJmlgFPUmejUDzJxjATci
JJTsm6a2IpqXQNesKD+I4JGr3XvshgyFdTcl+iFXR8mBJrYR8TWcXLU+Fj/H
SBS0UxlUbwR6APoyaoI5jfH7s8h4rrlmq7lsDTK59hjwr37cGRlBxah6gsVI
Fy3xZpx35CxCyX+gv+s9MvsswiTlUv8CaT/qLyf1WJCPH8pqalcavYDNcfdC
Z8Xt/cS+w7TcW861g+b250aqegRvRxWKDBPlUM9NQk8+OWA+Mlm/AVCS2eAa
OkC0F7pUGQmR4oe17lx2ouJIJGYS387o0vx/eHx0wvcN6qet+9ghZDnQ6BbS
fOVGN12j2A5ZCRWmMOpGXydVU1Tok/hx7XSN+moTVxByTGfEeFZB8wQWDxWs
Z8lsfBmwjvCLqaSLezF54LqJHrX9QGjNh2y6tV/kuW+tHXo6+E1SuYeuEP7Y
RjgQLzku9Cv2K3Bd+/F9200UzXzdkJaLEsKixo4qBW2LtKF8RUNtfROZ0DF5
D6s7r8oF7saTLNQkfBnG/W4cgFBbcjMDPnf+rZWcCLRwft+uMQ7kk2aCkvCW
htd7rj1tUw6CGvAiAaGaM0Cr8kabiY7CiCWVN+9tNklWQrtnKAZSAqwY8IKT
g/5P49Udqq+hgWZd1y2ki4eZnw1XU+JaoEFd5StY1mwIKYjeHMvK/uPVoWxA
TilFbCUfUEddv4gshaqgdCQmairgQddX9kzsUO1IwhJ97vUNIiYtLMuVd44R
5jJF3o+yJrxJl3YU1w2JLiDt7lib2c5T/d5x06Ep+CVoZ9vELH0bcCP7Jyqt
Dg0ekSo2WTdy23V/uqsqUKJKHQm6Tc7/9v7BsRGKwdlIc3OtHZgyof/jF0uU
IrbgcjfTscet1QxjE9YRytI1zPuXzOo4DAtfRqbKG9op5m8Fe1DCawjRZe0f
w67mKUBs6XoNR+gzbw5oYy1DR39V+SyMUJzWcsHcj5lflgJuhzj4cH6sSLLz
m/DXqGC6MsDZ/G+Xcbnyy/7XffgFdBBS7LPSM4P+UQdi+LznZyJMlpXAxanf
P92yiaM/wgox+SBgUO7mQOMtRNA+M2Chf9NWe+GNxMXcLVho8DXIUwgWaz9z
xHdqZff7mPAWF2+bUerDMV+9iHcTVlCdvoXD30hychllkfitZKfU/nKE/Dy/
0cFqoWwCrogKEUeY9P/2jHQWa8Mjgen8+HllUPAYpeWpRxaJC7HGAZM1/6cl
4S8o/RCBMXsAoKmM5WgeMTwXz49Nry1SU/y2faP/1ayXaKujaH2Ibs82aPab
ucVEQ19MeAL0cTZAhVZ0p5Uf7/Zb/HeUoqzfP66TQJ96e5xmiR23DKMZ3lBq
hlY77TG7U92lxL1YkrI3TkAn22wfbKiYJ0jC0dAPC1TBfyqOxk5vK7JcDRZ7
fx4tmOd9q2F1gyOnKuvvqIqyVSWnnJKMXgurbsudRBYA/NjjaWXhwDCImHUN
+Nn7lgLKfy64G4djavkY1TmvTywsfuZlJWA2PMAs37rJf1rPs0D21YBeiH+Z
z9WDjJwVrai/XBM95M27jE5ee+U9ukto9Y5NnsPJHCW0QZlEkoTnx3F64H3+
FTaNLYzoG5OEK/TJwlx7f9gU3lSEEPUhvx4CyuS3uCx7iiicKXi8pJ0e8idc
o0QpO/QwILvTzTsbgbcNVdihAB9NhT95pP1TbV1Wl1cWZ1YOE7k9s9WUlRxx
Uam8TYoi9tHu+NSQK4f6kWNUWOJGIletDfmmPLHXdD139Emtv91U5wEfTIJe
GCxIgBYV8jtSbmJScdxPwI7aWTdnKNEmIlOhVEpJInYqNKmpId8EiyHU5v/g
rs3XUusCPP5UW3qTQqKC5MfKniDLTVJNrt40xDhw/utMkziEWfsLV4hSm0AS
BoJipKOKKkpWvXe9ijJn4xp5s2LveWgqtDBhHRRgih5XW8PhO0KFK6qlmncn
zT0qICOZmlcRxbQ8oPK+GwDmTBUM/xFYJd3odv/HfcCEV25z4ylwpKJ2+LYy
0YZurV0TK1poCwdGgdgferYWbdRF3tP/UUENZLLW7ywcyD7XpKAdmwhzSz+0
E0ZjI0H34p4th8iobBKmPM0ceooQqLDo/cZi42UABWygF31LxPvERNkFuj+F
rfy6C7z47XNaWwCygcKRIQaNzr+RuBT/RMvvh7f3fJfLsJORCNAglX8rDXAz
4V5eGi+7MSC1zNR/7gDXmrPcoQx1lGkjpA99+/HEfFDSCP8YT9mmSEhREOdL
OcB0o9+K4CtdN4Xxc3K1BH9fG9GyscpdSrplBahd/IKIP8K+0nYZTmCcUErH
TI9fEu5wPj8pQ3OdEXMJ6t1m4bxhftOgXT8LjRY6vMPMkLRezprBQI60LOLu
ALe7Rw4GpHnPV87VFRzNNk8MSy3aW81SzLogcrWscXmWyNGlA0jxwD//E0Xm
Yetdz+bmVQNnF+WPK7VqECGeNI+HTLF5akFMC12b7ZRJ5CULQdHS3CyqY/31
t94h4vN0HFIMRYdefnR+R8PSDU9O+oKAP/WNcYNFPDUWFNkCUeNwjwmj9ULN
Y1w9kXBS399Gxc/FpIbXW/IMr2zUqh01ZAzKK8Ul1lbTdn89eFzIYl9fklFs
ZpqCVzHJ/gotJD1yPH6Lw8vAIb/ufgeX3vhTmu5EziiOudzfrnQQmD5y2ty6
JiSOSMzDwCG1+i299R8dClqc9+A+LQPIggbXJ4qCligKlig1PXYhjTASsGpI
XicWni2CVkHXvMaGFbEEWKRYzB7rVx0rPQXezj35Qkkjs6iTla/iTZ9XZ0CB
icjvAQ1NSX0kIVu3vbxNwg43ZW7LhrzDOVXeODTzGDW7MdlHY/p0X7pHbz3s
lbjvg3LgE0ACbXHtORbzSFW/tXWBW79j6HK6CNQ6XVgsQflBXhtn57km533C
oTXa2TcHuJQcUbWGhir7wczmPr0nszYofuEofvm02F0aj3SgGlMeJjCK+G1E
OKm5KsFMD3FB82d1c6k0Mciit9tD/PrOBzNUdS8gx29fPOYiQcQfJFUOHdIV
zMCCHzlCUZslxviEDaeyvguQKk24mFBy3sFagqmtU8rw2ePycaSroy7/gXdB
2FE43WgE0PTpFyyWEu0FvZaYUwPyHn+IQMmTIfbyecr23Mh1gzA1GMPFrbeB
k89JZCznLYoKyKdeZQgfu/IlykhPkZ1uoXCte8FGHRr5jHS63yU2KXO0m0Gs
tTV/g+/Z9BcNU2FeYU+LhuPbgyAtHRlJvyBa9vL6qMx+EGWCSvsnN2kdS2EN
V3o7iawJqbojPJYf/aSOMAwHY/dh99sW3j9sXTzZxNERHekVbnd6ZTkHwK2C
WvcwMgkzkkV1KnMZ+vTwpCMKsXab7XZASO/5jlcCJZbBx4S4w7TJK8BRUg56
JsLCDfH3AEQmCn9tAVcxqvZfs1/8tdiN6qlNdBG4Y3pDW8AWc/X/wplLg8jE
mvPs5vG4Y1d3Wk83duLIIsaTSgv6F74vkGPQRq4yV5AaXBfTfMbF67QalNWA
karvqqo2BHPLG60afzWk+vqaJEB8MMdPUtCHCBKf+pH75xwGUPx5zVOVHNla
7DK8gDzoFLhF9cTSi+XKV+4h6PxBWo7EpJDfBrySdTB239Dc3ynYhTPUnB0y
Uc1IyuWgDsbKu0GpiLyb32uTO61wx+AF9ByztAIFohtN80K8A5UGEY9BxTGj
i4Ef/DCAbfAdDhyTTf6KnGwwCfJWrgCQBQae+SS2vGXK7H+86ZcZtfQjhTVn
ooeKGhWqNkbgsB/EjtJEmJ8JYBB/e3OZWdmH4Du9YHeuw3MdDVLuSthtt4E6
hVNX/xSrHxiRhGifJ3yREgd3tkLqlc+NKUuwhabLJElPPJn4Dso8Y080O4Oa
9zBvrkGbI/F3ZEvH5majMBI4HzlWf/IFLsV3rtIJ09uNyrP3TB3Qndj2P/DU
F5QLkTJWgOYCRpU8EOjwz7XkbMHDT6NnJhohX9r7idKzOWl7CYlLwuFip36+
/1AqXsn4bJKxluXgYp61pMgPqQ2SsfldzImgAeBRf/GJas5RLA3T7Nw0YRE1
KASbxhY4tItCfa2W6I0BaofV9LckCWL8rnO8sDcs4yiOPV25uIEfdJrvH5HJ
2+gAv+z7R60y/8ukqPFzlE/uvzTmv7n5kegNa+v4mFuNXJFSYO5OzH78IBw/
2xJhqWM14vRiBIukjRonZXY6HYeIqi4Lu3xjihVT9cjeqZrdf+yMaUqapA6d
/UXU1poKwnV486Y9pY/u3Qig4rMsPIRPmJtROnE32mVHarmssaVx/eb38sqo
Ej2cGbzgfLc1bC/2GcTqxNVIN4MA1cNg6dFDfxadYsY0Gq9aSzVzLxWDNSkk
HudYs0GENhZi/yarH/zLATin2V7IOm/ipR/ml0GBSSmQg/ZiKwDP/Wfi+M6S
oY/BqnCa5nFlplsZiFoNUEYff+yOkTEKSj3/gn4xE+WeWefY5+LgLXttJIhF
tm6/oys6YK3qNrSKA1i6Hxf4ea1DmkWND/B+lsqIgDx/prwMj/KGXxHaD4Ry
4AQkCUs7MaQNVLPvlDDLmOySypDW5xg5QneNsoTdgDrsRWzMZ/YdXUAvvvKK
RqiBdnjCwXfKKZQfl+6rXDpo42wLzDO2mnxDvy+RL/liyTqXFS4Fb/GHchKK
HmkqeorQrX6XlNlQvsKd+ycWjg4mJD7bLqKI9XsfaojfyLvBaYBqHTVpWumD
AoIWVvuCpr5Ez1xrQxbPqykr+XBN6fiIjvJBt8iwtwzVTeEYOsFJhMiyaP0X
juqPnRGgNZoAsyFGl0o6Uv5frD9iEbFWJFEfjzRafQk2VvMiLeLBg9FANcGy
9//EFVvTNKBocUhXskVSCOtFYsqEkGw33ubkSFlOwrlnBWIB4D/KBUfZ8kL0
jGZppN74++wo4yqMboIh1Soee6QSjpIqtwm58omyT79rto+aq8xhWQIBjGyp
fwCfrMXPPk90OI3eODIz7YwB+XnrCDaQNIsUsCjCSTUADMT+P0f+zN3C+Cyg
+c4K+lizSc3wvskuC/Vzd5okvapyBakADGWj8dcSphoe11k0p2P9+RbSxsK8
vq/Oo7Bsr5072XqBMVmILQmhpGk2qG6xL19Cuo/pAQ4l6qWGH3fbrdr94nHJ
ASY07WYloXkS7zSpm4HbvCDda0fXCQTGI+C1mOZa6A3Ddz/HPIeVuWiUb1BE
b+W5ui8TgO1P96bGrkEdOBfFyECPyPCznNAUhZWhhqOWcsgf5voc/d+xz8vq
2sxGtpIWrbrbS9DOzrqsHJTPeJ4mLkpvad2HUhMq8CUnDMZn10qNAm7r/B3T
NxDyJfYGKsU7/YT3NinWAZT1SiS1iHRhEFbDI4vkQcwBQ20QyJTLz0jZ5y//
kJyfPwEz419bkk+74W66Tro9/ogQfC/VyWgrw5ZdgVJCZzdcE0HtJe0+OZVl
raREDFAfUz14JrYRt1Jv/f9GyH81W5dEr10DfwHiiVEMvRJPaazuQzv+pIDJ
+6ySsQwAkC9Ym/NOmwrUPNwlHw4xA6k3BYY43qBufg0qpbqkQOD12bPyd7tC
P+yk6gUEr5FXTW2i6P9RnffxRvVsuxdNf0wL9vm9y6lDT1B3KDKsWSK7KoqP
N8v769Sz6aJSD5xO4JNn7F56f7BxlejqWHLKhW/x0QM5wKWnVBoXiowe5wwr
Z1Up4gTdSrIQOMgrq+4phLBKvBkZQWfjUvOsmxus74tbBXXK5HeEHkrDurhx
qTiINXVxVYGbqhvGdsN/ArC16Tpx94Dr0cN3P4LX3ME/zf5kE9TIsYfwf9oo
3wDGkjzb2HdHBCzu8eXwPOpkr0hWtkH3I8Ef+YUuW1MsKvqQKqi00f755GTS
oa7xtuwq1pvH4gseP7t5IL2dDXrgmXHALFgbUUpze4xeyxQgkgt3nFfj9Sfz
qjN4iyW2/D8zkKT0Tp8XJhFaLQXcUQzkK/QL9E9md+UkfIW9my0Dcf6nGIub
vUAkTSVEudp4dFx0dt/baGhQAe7K3pq/UoZk3icV8ZKBvENAhKdYM4m91t5a
r1X9qpTjX5RFaqINdZTZbxwjp8oDIjRnAmeEu6c6/hqVN2EoMBwMQslf4748
EwVObGobct9E6Qk/Wj5ULLHfKITvicQfLoiCUZvdfSvaQiWiC/Eu5HcwF21Q
K7tkJVlqCu/lTf7mjQfGe9KLKoRbwoYtKxiPy63xV13F7L89YmWVKVRMZI0B
YYpIU3KQNCT5WOBaWHSqGTkYJaKLkMhUMA9iN/TymACirX60XRm58VCXfLxJ
OcaRcWTc3w7rT+MmdINkkyKTYO4xG+AuThtSL9l3Xmuz2mZ+d8GdrI6dm67v
QUfN28P2xtIY2C+ZysQhE7JeGRIYVQPdzvwsIEwjf6lexCGhM0rshBeY1ruR
j9pPy0TDypyaoEvRJzr3opxpl6F3Ol78fNMnmHtU689Vd5qXULXnoibuZOrP
Nv/ith/r/VFqb1g0yedIAXGHSAcRANQjuP2zQmGpTV8cvhtzClIru7/M2Dbj
kgvmkZkjIb+GhrzEDtweWf756atWiLwGxUvdXK0JcGG83OOqjMWoAN/1+jN3
i46lX45849qEMwpL2p9XO2I6pWEm6V2tx0YV5C8F9nDVGzkVRtt0hNADRRzx
4n4y80u21uWQV0Vi9iXzkp4GfI/uDCIv9Kpak0uQ/5W+rccSRM9dLpoJ3AyT
w/kRS4i3W2o5wcZISPpoPPI4fjiaiWPnoBAbsfOPi1KXoNOMzu+MRD0AFFV1
aNqNSPMqQmbbEKMqIAzEyGwNt8eWGpiLUw+kx25sDV5B4+tkHXgYrrnZwz/Q
VuciV3csztDryYf4MCdu/dSIurXPl8IK+8/yvWtRu0W4dSKS3fYM2l/HpW5e
tx8UjS1htnem6oCz6xJyLc2tA93wyqLe5qsu13ncricPJIJbJwr45+l8nKEi
jbC+ney0c4wlFRBQuEkAOswPH9/qm4K/L1NUsqvSFvqIXHuMIatg9AVmiHrd
osG+jjJpOHDi18hT7rCyM6SuUppyfCR1hjGy0/inL4/YBPgo5/tjf12aMhvn
X7vupdJ5IZC28yDEO9OzTU8Hv3/HmGAoCOLzyJcpx6ZtiJLiCnvOUrIM19Ka
6D46Q9qMiovckF1Z/nQANhtISKnVOO+TkLmpLO2gpmpT9WlWIxCKIGCEFvEH
TgkGDNzTjujIbLiYaGDJ+W1sYYUEk/N4/eyrmnIBMUk3NPQVe3cBjnf0UTiV
GFLWp8KqoUm9iAU/bC1uaYj+NWG0BxHEZK3cEs9wqxeqJRRRU8O4OIsZ/egP
cWjNOp2p4dVOBhiFkl5D+N45qK+AOspBC+Q+SEJ36GbRbW6eI/9WU2Fh7atB
W+GVVrgGs5dIj5wkXgMjRGyyRuyVLZmwXxT3ANHLZl6unJCXPA9qE02j3oDX
xSCB2oxGessORqTp5sHfsVGlMqPmty/OOZ1UkeMe1rpJnjR7SWLdSU4NbPQL
iUK36O8LZ7wsQ7B9rPu+kSD4PE2duAhaDZYFOkm4wPY1qwA4ThGPrvhnxGRN
a5ovedWoekSwwton1VcXqVVBtKr5nAu8bupsArHkODte3JcRcx8PTfsTPLen
AKhPivDhIFKGtS++urPPLCw8jdnl+1X9THsHtTAb8+r1szoI+rZKSU81dH6G
azBANMy1roJOq4mY9tZvwtYUqC5ffz7TWQdMFuaAMPBn7eVo7ptm8qCMDNN5
yyfDCYt0w5mmO4I5aqsvdp/ujgQVUUWuj9HnnSxCCk3rTsElSO/Hm+PUCbyc
JIKhdU6lunjTcJXEcxpLIhKlBo+T0o3pDtl/XV1x/pNy4r4JFI6OcNnIMUqf
GB90pejEgiDoFXCXarmdBypIoB6EhEPx7UIj0LW/4pwlkSqtZTv3IMrQBU0r
jgNkloLX9M4MeALDtAG43lfjSqX8X01MMQuTSpUPXnr0HCY9E6IpHyNvBqGQ
0PzIq6OboSnGgpBNDOgSUuLl/pHWSy8JLm7Sh9O70Ymr0LuFAo3ycPZSWK9P
f5wafurKy5+qWzzTLb9usTTWTeJekFO5T9NVvoPKRhG/kePsleKrD0xKNnOj
PlSFolcnzi6eHmqV3aUXl8bHgCogmc8uIHOLmXYev+2eYrqiLEVn4VLCpjRT
wBGnpRlwnC3FtTDzWMU8AaG19ImhLSnpoQKNp+jDAjL5Fj6lwFHe7rc30hMm
hq8jZFteYd2QtHJQqGPAqH99M+htios8mw3Hq/YJrrxq/R2oyXEt59MdfnoY
uMdRmFVdzrM92rWSPyc/IpcVWYJpiqcvmw405CyrCnt5X1irOnkZE7BLI2YK
7FK1KHqdF4i///cxBXB4UH5M4S/ffxWBmI8b1Pvu4cagfDx/0WepHu7NGzcx
baE576VcVilx7POq+tTHrZRKal7oroHtthGggFCNWRy+3xwEDNNib+bI2qwH
k1N2m+FKksrQhrAA2yvicfgNQuGusAbbAdGhrXWv/OG0dykas4a7ZsQO3deH
xko2r8NkBR54wIvc85ldxBvI+DqOFd2xXVE6s3I53oC8czNkDcpmtiZRQmCw
DLjWxBi4M89YXpdrSi/5Jl7a0pJbvGBIhRr71odHJcZx05va7PQ3ebUagCoM
5KaiPhIkWYzLxaXtn4uwh6HMlT2yOh8OXtofP7kotdGYmc0oTv98crR4rpLD
SPB5atGNy97YB3skdXY581Hs9dGydgJa+YwXeXYGrgHE2IShRboq9XzJNPuW
I2RHMJl7R168u7hjyHXJPrp9cNLeaGEpwd6NY3fypxdlosDXBRC03+/9NuRF
UVMoM77hQAeucBZYSFfMlVy6LVilE3IhC45sJIMixQ3bRBHovJ23GkrDyOpm
FuhAVUGTM/xmbvNaLTo06ykqlYAVM09/puq3OpB+jooI+ohU5AUVdENlmyce
r5TbBBinpLi1gO8Jxm92zsDhDL363t5YPZ2umlo1U2bg4Wbpdixg1KS4G2r1
5qB9OkTiKlDkZ1M+hlNmhtgu723Nd/B+kg1/w8QBBjtVUo1h4OR62QqzjP3r
gRg6lu1BtGzndWI+GoCv/wt8x7BQqPQQDuJPXGWE72sJtavlzuCNEk9h2ADq
ZQrMRy0pFEywIt42EHEqeH5SHprMK9wYP/m7Tbb4bV2nlLQsJB+HRqgyScZy
AyfMTrULu8PmKh9EIQCknmoULB+5h9PE8DZPSKqVzd2XBsGzFjX+VmueH8M7
KidMedcvhgDOKOBRL1ZOI1vTwhv4lErbO4NWXBGsfYRcbn+tkj+QkP9Dsk82
1V11zeHKUZaCVEkpODO5tPBtM+1ZUQeCADC3fU2Ycr7zU4SxcQ6k5BpOr2Kr
5EY/XGCGdORGyvAPzciQiYU3Lhii9b7RJM7gVWCDJk+KsFk9XgyLEAnc0Vun
1fk4kH1j1uwb6jJwPzY+I0UpjPfo550Iw4YwVAerWOyEhmaI8i7byGDOdAwB
+NDQWBlRi78Z2lYr5A+jaJ5NQUa6AmjOBFGFJ7pkcqtlmRywf3D/pfxxNZTg
KuB9PE0ktc9xk8IFKla/2uxn58uZRvOwvr2g/eM1UFH/UpAquKFa+MnY69zl
v0xFDTzwvk1mBkODNPlftENja4KDL3rpBd0vyeDLORXwWCjeGHYdzW7gKNQd
DNL/k6BgKJUp0mAcVnyuqzVithy3U+dyvREtW+d4s20YjEjY7pKKfML2Fkzq
My/GyrAqlI3LoXD5DNvs0Bm0yhJVUKyQM0Gv/h4D2Y6di+oEIy7cAFv/cih8
Sq9Vpi/EM4MTItlpU5lq031xDwTvZx2LYbOwNGYCsEfvpNxkcnHBmsohmros
5eR4b0iC2SyoJkKlrwpt5mJ1PbFNmXqaHlE/CCkGjo0+hAR3itUKdu/GVyQY
jZP4wSqgVgqvvuu5XEB6ID0HEJg53ESBm6mcPZlVbR2DT0vWrRKguOAe0IcZ
j84IouMHg60BKuAHe/PVw7zLC4b8I3KZnF8aVHmbBHXdaPLnoKdn4iVOCC5f
R83uogOQdgHFMRgIFXVMZuxiiC7LE8Wolf/Z9YyxvK2QZ0mvjqHDS4ExZ8zh
SdXNoPDxvwnfZXQ/GJLM16waTChnJgC86QPWd/y1jfTxZ3c581GdcqBh+ru/
GgivkjSURvEOkmUis/pHXqhnTQSLY9crJG5scpV3f7JPj39MYrx4jkpoUspj
WwwjtgnRj4g04pmgDitBENZEn1ax5Kx38/YsxMWMH2ScPBkBE7YraKZsw76p
n1LaeOr2mV0ixFDxFuuKN934D0k1Nw7HEzDxnfSGcl5r89dj4nyQlLxvZAHa
C7v9RjO60Tly3ANW80iw79Jw78ErwVwQY+lVm0h9szreTrM0RqHExqoxcS9U
0o4cVc+jHoUHYp+Qjo1AREnjZjt1nMIYFutZnGrLA1q3mSledqF9PAk98im8
BFzEmUcsBZNBtk9mzwivE2jbE1ilhA6IYufkwBlQVPjLc26g5bRr/R7+HEYr
7AiT3FgSO9t77FPms07l/SAfBiugAQcAwVtej0++5hsO96ykEiKFhk1MyuO5
jCjqOoVExjl968yPmUWe4gwO5njYNlujUQmzIYSNmRN3D46f7rhoMKhf1tm7
9RZURycwNK2pfKquE3ye/hs1HoqSrVcxUnZM24Y8nybLnuaEqGt0pinQ/UqT
1I+4+v59NjytyPf0p5v5FtnoovzWuCRdzpNxTVPFUJ+VJ2m5GJ5gUg2rrVsT
vE3MfEe2tZTsy6VGNoS1wcUPNvtvjq+UQxrBKFc6ZUB/UcA73YbjptBg40Fa
S6iJOWc53qASw9DrxPxiI1OjWY6SsKBx+pJgXeQrm5KijeaTlQy90FQH3gPd
kkR3biKbz3VJl3nrMWDsXq8nrtbj+eWdjij1foscftczhbfwSpzZ8d6i6g2b
32UZy3J0eJqjSBagPalFCmtpKa0kwlCGBSX+oiTX7Nz6uox0vhW66c+MkODe
P2gFAzkHZusMbrI7MHwkg5eDt9S+Zh7455gCBGO7H8VS7s4iuxh53+ms6XHy
F4+VszIgD4nyNRRjBAGcwCz6aOiw1Ok+iOYdcuSi+Lo39hdB89P1d+plf82h
hVFJfUUiH9LsG/U4jpJOLDSVEcelDX/iUbbqLe1II7frGOI5Wce4Pg0mmCn4
Qt9iHWg3XdTOfC6dhiNkuOSE3Thf7zDFF3nYRJBPWSgBuRmYLdd+TQzeXnNe
/T2ce9Aa4UQCI4Ak+UkWAOJSZPk5XEooIEPLFIc7QCQ9plU/iT74j+OSDoWs
al6VyRoTToALfJe/rXO947QGK1naFYWN1y3SCYAmnb66mgIjfxU2auaVzkQI
4PK/DxjhUa3jOioa+2kvI0GOrRvToEY1UVGqc2x4A3PuSLGI+xOCIxj3i/Xj
K4ZhJa8QrgPrzS9FCJHP5tinAYKcANLqJYh49nuDUP1lLjktcITF8vw69qib
fhZs/gsIxZEKzZ/WENAiM6qX8yhPbXCv9NVvpWGAd9UsAhoYO+FN1TXoYfSe
ey8txNSSz8NweCuBNJHCIidYyGnArFsWN8v6DLLK/8ogwDOXhTmWgmyYQbDq
PD+5A3WC3ESfGsfwGV1f18rJxM1BMXLefa28bVbHFpF3720NCJDe61CQ2KUB
hmyqW5TyBBuwmRLEcaODAvMEoh2sQNJq6qai7qaXUG3xFP9ekTDg26nXFgJU
Tq0CZmliUjHh8Kepe1AgpIMhsVaTZgC7jHZCB55r9MrKVFF9+la+w2iPisIs
LojNlm9DxQOjhzWe7vLPPqA79u3HbBji5ql+HvWxKV3JEj+6tysMQVdTasmf
0+WLZT7sJ6FiKIBrIblpJe3UktulUx8YMWwshE6VQ7q4GtpJx9Hqz90+mwhb
WtPJh5A1uB3qkOL0X4aw47h9jqvRbVVM49JjnX521qRLncBoEc2UyH4JlY6I
3/8gQ/C2PvFVxBZJC+AcQwrTwhB4MkJ/eGTBAIDPgrUomHfwgzCxTOnPip/y
BJ1G15zMZgolWNAi/gYI3vQDo/e9jPZjs5KsuN/b0eVlk91CAO0G66iRR2+5
jjKSr1Rym5mo26Ss3SJGLdYH/rIZ5BWc3fg2QF+aLk8tHqhToSZ+rb98d9Ap
SddNe99hWOhrEHbZjYCSlxPSdEeA6p3ov6MH81XU9aytiwy6G2nBM/dyMm+f
m8oE6IYVl4W91mszjfyoVSWE+W+ItvGjfIZyGuRxWCeOf9hH594ERjt5MSnp
wSi8bfDxroyYhK5Xap6IVhDwDm+ypzmWGLhGZQMxZLsFJ6G18l08qdFqPjL0
x7lWJfultdueerXY7eIxZSoFSYhk5mOl6Nd8h3fnXA5WRDeniT9uYUCFU/tu
FKz9UQLLL5QCH3tmtljnD1J3jElcnWYlhCn1u6M3GX4z+Bp16ox3lD3oM60H
MNBMZs1E+0Ma5j/m5aou5y/yygDvta8sqmMkRm+yrpiiXEaN7Kce2i9w+f8S
LFAnL17KyataCOzjc8VHb8h/JBAYP3Z3A6EcOqJkCvhrQZfIRvTl1Oobjmsj
JxZK7+kcilxqd7QbAaehfDah+FOZLG+0pqEKU3hO/TDR68NlarOeG2qryYPD
CVrpq8whJEsCqpq9eBVSAgubVJovdur+6fakm6fE6NOaPzb+PkcnsLq1BCRl
fCmp9C43RI0EnP2LXeU+J1PhRAo8M0/ldnRRrEOL79x+KRNzTawFv3+Xx+nO
vqwB40uMwsnV64Nw8vhQo8BwuDqLOEVCD4eoaIxa8jSZF+GiasOqtVWdubhN
6FxDBdae32eMeKUSQ7OC/3vLkm0NnkUs38dSP2n1EtfZfAQSzngwZL2NyGOY
qjjwHc9Hoi8/qXfkeOUkwzjEJThyq3VIn+F6LAbonYeTE4L35sAcWctJo6vc
JEOafo+Gf7TTZgRfmaj6JcEXE8sN5JdBsaKB0CLfoMeeGJ5J1KOdPsAD9Dg2
yk3l+LAv1SOtqATVOHRc/2WhFdQSTQfP2Eu+A72f9iiWSRsSmST4TPWrXWwc
txxHwW3e8FtWyWqV6HKwF+nWx0cfqkDXiUpSq/wUDLQve/RZkS20+lD5P1pa
yneKvLPZba5APbMxEW+Uqx+nlgHBxd/kVWzIUwK4+lIyRD24/kspkvT/s2CP
zxdmd4RemZtb1hOuS6jTxEqaPZTqoQmKKbDG/q1/GsnoRMbBSe2IDzVrLU+H
qfFOqUbZ/dGdqIFKIzVDydM5lav/Lxwp0q7AKhdVG0bCuypVTqCquJ8NVagh
l4HfscyzRxOLzF1dJ7MTNs4AEqk5fT22hAgDJIuKIWvEN0Qq+k8qT1fiNfl3
RfrgjQUgOScl2LSg+kHHXF0HzFL6J1qAGqFMAzD9NEGSKBnB6e2zZ2M7Hchf
xl2S5tSLuVfQuy8GZihmkmlECzhy0xfxwcJIXLG2aPQXPXCGOUDV79Tz/SLi
fLjeqvMRYjh57CPkQ2dFAA2TfnSmvESjoAp2ClUCreyJEY/rAR0Jq7mHRGwv
+D/MOhkU3T6xTzTMwjrh7/JJM2uadJRfiPUOinkbivnSN8DIuy8JYuR0RZB0
eS0TEb6Pl+zlMKrvqxnzXewKU9Ca4X6q5OxIcw1HaxR+Y0dNH2GnVy5zJr6V
lfe7FMsc/MBNuSs34SHcUdjsQmntRIl/3KvXNWU6njqoC+ZEwzh18VQNWZbp
45F1IkFj+qdqfmqdAFCpydG9Thnq085QV5LZEky8G0yuzuFAf/5FF9bMxHoF
d9iOketKD/d1HlA6dS8J1ECm5AFPzy+bggetdTmaPuwvbjT435I6GtPBhxh7
3Y+Tvd7dtnvqbEQkyoYo5q7Vhqx/b9OgHck7pdPW5mamLLPTuTwKkzpepFF/
guRGO+gn2++96rlbnYghnKh2WxlwaCcfSrJOTq0hePXAR3W9rj0of9ByadRV
6QhlA6Gcg6em5CoI/O/GcYIdoAwwLauxPR8muh5gxcStU+NzMLRff/gbkHT3
1asQ2Tk+dE+GBe6vBnqM5gGwTjN26uH1vvQua9mrLeSKkW/Nls3WiePCMUJQ
lslhldydE5G6u6hCjuB+6scc11RGQTDZPmndviqXO+zp3QjycANWdKaCPr+s
FN6IKxhUW8laN4t/gqYRHhPsROhU+IZwBb7/vpONmWsKjdgFnRsXOvOXt8Ja
tLggUtYxdHpVtMKTmiyTM4DrJx5M2STH8eM62daKFoGwXpB7vYyZZ/FJdCW9
c3O5wLGc4yG9R4F+rQIM3+VPwLThyHGf6Mx7EV84Lba3IYqTIYY+PA0A+jrH
XvwcFJ+NsUr7ZAyWk6xjKA9R2S3N8kI/kfyXFb0aU0kFSgCyrTVLNoO+PVmx
f4QfWqVYQ2/ayc6x33ulnTHfmY3nXR7NV12rFyjZ8ZbZLf8uIsusiORvovNp
1D96peCIACRwWGIPhPhFIP92c5dr6CWKk9fbRw9bQINku+td5uuWSCdwRsCG
+pFXNl3jUR/c3ZKQImMHVzlT5fmNISbOt+8qU8NS8cfL6p8Dp2tTvVW1GuIE
etNt2XSYhGwHgxPmrUv4O29/qo8OJnu56MbxpP/KdFPPsIAwae3NOUCEbLXh
cTNEP0tBkwkk2d7XQLDTrja0FwbW6GtaGtchQDdsQrymrtpRxjm5Ya9baKDm
s+FEY1tim6uSDSLH0xixKL0Ye5R1xFpAwYcoUyq2wwRyfusBldVeMWC+jEOW
xnJ+i2+mtDZyGqI9se47BpDo7e1xbdKsY0xQCb2qfBqooR367EFdANN50fDO
1ETHogIRuCbn9kKjnIrclZlf+FsOZ98gH30AVeat44zBDd7aECPmaSX3Y5wE
8trX/RSEHRdS1s5POkAkeN+YhtCIZigdyRSJt0CI0Cx/K+Hgv5UV+S4ZUys9
1B3aEQ6YRkG9gk5kt2AY/1I9IbUUt9OB4eJKFAxirheyGoWDVndwtXwV24rM
Ft5hhYe0uSXwTK3tSTiWmUqHPm9WjAAXKL1mNpcB2T3e7ksck0n21rTISgQ8
/JD9YHMdKML7KC50YV8MoUjizoI45aj9gk04tte4rT5dsBlBLOAyPtYuiPQz
B8Pk/dUn5lXCIu7o/2ghe7gytJ6/UlaMFBoTCUL4GXrwAAKaLmJb9y16k2Mw
+aKU3s0QINfLkiWZpYwXCHXBlq/TpI58XsuO4PEcFUZTkYsRgxxMgtwVyrcm
weA5T4QS+RAwjMXWF3NTn2dVadudmy394LNETH1sNPmwQBEmgDEOP2eAbAAo
+YXMj8VoRyesUVH+iEZ/Ug+BgpRBgo/9QKMCX4NfR4zjB4e7YiTpTKXyZy78
dHoUljLYwSTVhWyLfIVbWvs3qIFhc2WBdt01Xvq5Gw2ADtsevS4YvVx9PglQ
iHsxqECuChacg+owUzRW1vDeLvEpmQ86HEntxomHJdsBSeqYOodI8rTDhRO0
AdpjniQm28egyR3KDIOkx07C734ir3TQpCBq79bLs0mSV3UW8c4IQ2fq9a/B
XZ6IkhgBXcMG9KvyIbP6ISn+xiY6a3Pipg6jCDUVF0HeHxB/gQh6ltEKYprX
s2s2v1uW9SPDeF2QIHtq5XqCcT8Q0ctwld6xHsONlUirq81qA7dXbtWx3Cl0
A2mMO5WkBVE9OdByhRqZ0JK1JTpRtGs5PQ7uwilTY5Z08z8brxfnnKkUXAgY
5T4b8a1SsicDWxsfJQlkWLK/VzUkBV7Yy9sRJrbvqpZtYVnoYJUySWwujyJr
UVzpCmHSw0m1NhspSzugEmVdT83aD12zEFtO2BDDxCpQ+r6mVunInNirehL6
gZYZ86t6x9sIwsqOcvGZrfvzlicJCzyrFlknjTZ1MaTlN8ZXlbrtrkwurCO7
YPSiqFE/n7rN9Ue48JniUY4/HXtwoGPEfTkpu1WevWl7pyuoHpy+eECfBeoA
BOFmLbSm21uTYLFCIotOlruwMJ2UVZtnyeCLDk09Qt0iBb0PYPoFDcK87RmC
J6iAKH8mvYPKH2qzP8uN/hME062jIwzgzk2/uh9ajVbdC90usGrD0qT17UYI
5OGnJPCMEZ6g78CK7YA8EwFC9CfTJFn4vewKNZ1kVIhCvRDuIKM6UE9qY1Kj
U7LZRQyognn633vYKpN+mufksaWvahjxvjQj4D/sTyUxYY9PKJukj9VP0ZZC
WNaPFhbuoK/hxrVem75nU/iiQE0RJdLojR8yC0pHpASCvaMZK/ZiiKRcc2wc
vjcPFBap/Pg0sQppX7kNADkgSh6qexAuCVKAys1K9MVpK7e4BgH2nUyLaPuW
EyUu0llTPBhpeY+aaHa9AO7Mx0b8QEUOX59s7DMjXubwt5ARYpImL2+b2d/g
3L41Vs5tiVocN+14C5zCJXF1C26l37gT5ChbqVjotATKV1gntVQhMjVpjjFU
WfyGRJjEJEAre3TXIb/FiYKb8HmxzFggxeTFfsBL+8bKBGsTpxfPW4AeE1MB
8IMU3VMbzm/2Piy925rbmYvpJ6a8XPHXO5i+jC/2Bi3ya14G1qEeiqinFBQH
SQ01b/01QAK4RDkOVhY2pcUZSKVsfXHvhriqME1tTehDwvqQXZ0Mu/CdgmKL
Y0Z4tzqJfFLI6KeJK97F4X3lAZFhdTlwbGT/NfGgBp4Ju7VBuDFLOUIgXeIl
PUUEz8AVreyd4PA6BD3DZJB3gBFOdwzYw2D1qI/FBDgDpiH/r+s/5gLZ2xgC
Dqq1+MA5MSmTkcL98LfBw9eqRJaOe2EZ32nA9nJaKdznfhTswgSfbuLJWEwT
Q/txBHvgM9X9pc84ePOwIPgLN+FRnMh4YOGIBEvIB8i5ZO33tB5IBruTI4Bs
hMriNXFWeeWMmSJosU/+soiA1V2VqjtMqtsp9sZmowIQTzjMV9OsJuXvmFRA
5XChxpQ6vRrMKdTGnSEWEyStXXbVE0fcJQL8PmPqmAcL9eeSCAu7kCT3mtnS
bvmbUPk1WFKZwvjFdGW7aXu+f6q2LvH260dnlAqynZ2aJs+UO9SLC4/u+Yfq
IOgTZ6ffs3Q3v+He+dvX9LB28uqo/KPFwTZ1nokx/1fXT6y28/lJF6wthJ3V
jU8pGU+13JqBCfFB1Pyi7hUNhsYBltNzEu5+g37cjy651a+L37juVvRCIRSU
Zl71XPBuBX0XjtU0WNDC9BhT22V5cLLaoKg58JT63kmuqdGg5XQyjC4ULr0l
e2sxd3TWj4e2ypZuciIJkQ+C0M+4VVzAj3UMd+UVrmkU6ZE1O4iNY8vLXE7U
qc/HCZGhbYZnSl7OgvgU2t4+xWG/rBDcvi0FzdZxOE7sgYs4dpmveD2hB9no
1KtDFDMNkP3itMNFM5frvtqwvYhUcaPU4IdcpfHI4RfBDFaRjk3LPkO9Q5WC
IuhBBNIEAd1iH6lyvNkhYWFyOVmfEpTNwn7/s8jEZwNRsM3D8MxYha/Zn4li
qXcxUwhsE2ah1BCi5d4uQvg6+2/29Re7eTu9HqWZrjfK2WNqeNXmv4gKFYa3
C+sK15i/TKQ9o5KIo47MshysWtlHgITGz264kUagM1pBXqtm2NXYLD5OfmMs
wvV37rdfEAZbMZQ7baC7azdSqrqFGIh+KWgqRE9UYMO5G8RQnulfn+tQ0prU
Znxp1qV4nGE3UBE1nMuFhON7xY0uKgtTAOGJ4tTG6VWlBA3b2EnVxJpTet0k
GZbmBTZBmOFdKnlKdnOxQ1EgRN0n5A/Idky+nIHL4KZv8PmflWVXJEHLKJu7
OY3aJllLiX1gAUgxrax+74yMrxOVNA1dDvZuzZG0RVVr3/8j+6GUujlWv3X/
K3dAFacGX3vQ9e8nBocUHT+D5puGskZtlXarEs5s3iXw/D0qo1J62TZfP1+9
WPz9+XiF34aShUfYD0RLXDi9pn11x8d19ItYFbOTlWUCs/dEREHtaPySrNQ9
SqaMwUMxy2MmhtMJcoTP5hp+JLy+4nGJVS0Jfw9v5LrxFzfWIFaD5C94YP2y
AzwM+p+Uy/CRNo84Ck5usilLBcp/LBvzDp0eaYhQgRVQXxLzY8QAwF76wd88
z3nSwbzlyBo2g7yLMIu2/WjbgZqzhT4NaaECGurpGuoVv/iI0HajMjdF5hPv
Fz3dwZ+TxGIIDeDKZFs1BC8BpV3SUogq/8SMaLskguycOtWWFBUNEdplC2l5
mjqwDvkf0h9I9jNFgcaFBkAizF1kvQYVyDkoAAf14XReaoFGmA0eijprJQ//
4br+F+COGG0sVzREb4XRjYefwYxK8Lksb1hqRFVzVCH3if9fwvsGUmYgmdeV
AUf7m5gX3rbIcxhLOuu2o5A5NTU9oHxInJyJ2g8XkYW66KpbPXu2t38PPJMP
9LsKKVEQBC+rJtGvVg/Q5ytsbUDMqXSJW2yRS1xptObrVGGIRMHS9Q1DnpOM
OCWGTxf/PMOa6hVF8XvnyWcO71bJhF2lXoiOhfJ6UzowzhDbKT37N92Sbs1c
T2PvbXY5L+h3p0I7g9M2D5oW3jyBASJbA8B8+XgmIu3OmeAvzC2QOOktLyXg
8RGbWCOanxTjC35q4zCb+3ss6nTIw9cS0jiYq3gRU6Kvpl5e9InlEoWdBu1u
mqMbdtdC4CWZTyVYpa7st25tW1aSJqrtGuSkYtXwrO2LMZh+NdTw+8anZZRV
h98KIN07u3Ru/AcAywSlNbOhbjpw8wMZWxQa1bWMDXxUuIDWP2bBAhSs9Xur
mXj/DZ++tFvIHxzakcuFTWEfWSB/2CNEJGm5iIbEM1T9ziyoTpTIVZ3fQ5ZW
Wz/P4Vt5/u8kyZGjjjQIN9H1HWvzqhspXpfVpHnnJT7KGtsRD0RwPtvNAPSU
hNITZb9WSCnTochk2xtgORXWDh6W8mCvnj5wO6y/HnGCicz13hvfYZw+XDMy
9PwxqRI34fl9lMWTUcTXkp7SrPwRiOznj9/Iq4jU0eMDit24oESkplGDKGY+
RZ21w6zhSPtS0VJC1XIRNpZwdilJ3RuB1ApUWiv/JmUdM9lfdXUceSj+aycZ
brCWYR4R8m2vf1pERN22SIklFdBnJP3L14YFiR4d69OsfQmpHqDKUxbXy01P
27VbgMDEiEl4rxCqQnJil8b33B+dPb9LqqvQK4rfKPdKjVIWGkzwOcQh72Cf
5aBOM4K3UNhrKsEV1eZvxU+Oc+JSpBYlecKSq9K1hOptCE0R01j7/EZ8BqSh
kBVPmr5RAecxLE9Lv0izFzQRaw9orwhA+JvBtpeKQJJdxPAqlWVhGtIrWGMU
GSeTcCjwPyide+nntHa+1+sj3GeR8MEVE1EVoqJJdw9Zd9TvbdVhijHptcTf
PPkNHMkBe/GRdSoJTTXxZvDS2nkDHjkf+pzwBSrtYNAbmNEgGuETDDLs4veC
lO+hd1RD3iTZq4xQPbQO00jZVXZp77+U1+dB3yW4h7e8VJvoz7yv0XdPmJEx
w0cLhTrkmHmGbhWF7OKjHkSLZf6nb6b4E7ZQXsf/tO6gRdkarsFjAUtbgfpP
yYIbRmXZqsQwCPCI6EyheJLEB5fR//2GTVO079LuIa00f8zvhEdLWfR4XYLd
o7hIEPaDZnZck1cSQw18GFLVCaOJPEZ3rJ35rRnRNZHJ9+pY7po+idESOqnA
V9Eh6Hfy5MFggRHW9z/GHjLtw4zIToQyYWK7IC7IXV15T5eNKXm5eOt59Zfx
ZKuF/AYxnqjpJNg2yztA+z7rHBy83dhPHFJ4R9lwxEMqKdg7lrC83ecwkzOP
lSA/8d1lTCnjSdDTklHdCaVG0QZVF0avBsiHAHXnFzhl8+kgoMhf2I6jXBhi
RoRTlFNd1DRUXnY6mYui4MPaT81gPs7GhszXuCdVWXme52kefMVwA1b/ZXzd
irgtlUe7LE+Vx7IP/8Xz/wwCjEwvWC1BN1gbdud1jNbfb252a30ql4zLFN/i
dCY8/uH3d0XAxy0V43c6ehFygaf2sRTYsF0agx2ibvcnWEti3grT+LVPF8d4
5s2bw3zU420S58tr4RKwPzJhn3kVUtbk+wdZXAg1KuuKapBlLBOKxBfat2yT
TM/9qzDJTZTFCUJduVGuH5MppbP4LyvmPiJbTlgEoSby0/m2BQwZ4mhAATbH
HCmD7pVIEiHjbqnvruecg/xSORfxLsYew46u798KpEtlLbkJqEagkPY6eglL
nm6Pe4c+gNLVFqHjAT9JYBuE86OYhkErmQO1rmKlMlf6JRXDOGgSGzRPLu2o
gkX/hJ2edvlb/Fwf7ne5UDqCyXEmFXGM6CXKgJi32v9S1/jrLSK+xRNktkQM
g+0/W4Dq4p/OZfFKv5hEoXbzdnufs16A0ssblWeQzQAgw39j1EX4ockQo9yz
socDBMb0ck8hv6fGLeS18JeuLYVl5qS3z1ZLnRmRbMm7Ya9zGH8JTVEYtAJF
xQIMM7yfR9TC3hNUyLqXC38//UilIh59AfX6TdYDxx8maKkq/P9hHzQQMZjO
lHli6PMYuee93DguGFmm46o1184Pwb+b+MRBi/ugFTVCCoUl/las1+9ooRFy
F5SCwjterQKxC+4vD0QvDCBprtiyZ/Cc4IdJxn4Zu1tVftUR5tOdHH2nkr41
54VBHA9C0EjkaXco+gNZw5ypyY7i7p0XjLxfZvRkLR2Nrak11ILzRbtyePWW
V2pNXBw0zNKsh7CwiWo4zU8urCZyvPxprG+hjgqU7FABcS/kZHNM0Ahv48iS
wUVFsp/2oaN6lGLnR1zRhpLE9ciSYr3y1JajkhUkYNmGtg0abdtKOZ/ykHmY
zO2FJkOvmYTFON9ufh7Fs/jHq5xIq0CvmZoQDpK1hvqtL28RpTUW57pmxk5Z
z8cplp22GW9XyK39/QhM78KbMIB5xqy3N5+YCSpntsgQYmiGd0YqgAYX3xW0
7tQHBe7NSdSQIhh/j49hlEOyFNpHwJNMS3TPcCYPYNuZ04hV7UmOYBMHgDip
Cw9z31JxqSESY97u9NYkbmTzoXVBrALEvwfRI4yxpgwkje17eveDJttwvYxP
iwXICB95bk5fJGvPhxkNi1eZEtIY2pBKr2E6VNXLZVO3KwoOYuwKtIJH/0SC
6IOMzhVOfGUJQ/jeQ5becBxXoke0uwyf8c96iEVczhj0SWfJsT0LKJ/11j0O
rs/e6wd0q8T5OC+YVWLJ8pVUjXt63rw8piBlpwSC/kmf30l2PO/o6HfG6/8u
lFIKYU5Svzs9ObCW2RAPYQfUDY+Ge7RpYpp/h7j4SRMIWe61NIsRYXQqa650
ufbKsCbpx+dGZ+jz4DFaWCGlcWiMaHnXCxF0m+PIlNe6rvhYJXDexBqKYpzR
kp71xzR+0TxRXQALrsUoD/atQPbKVJQMdkF8F6RjOPGzqaVUx1pORzS7ttev
Mf2h0D2zzL413HDCfwL4OphX3NBCnilrvnI+LilA9+hFL3V/oXEuMx5WOPfx
gPCD1nErq+3+V2O3kv9wdyoGxrQZ5Q3pgE0SOE/s8nWUsB4Kftp9JGQjt7z9
d6EsT8qm5VNhsY+IwlHLkFg3Rp96fqhTeybQL8xvHWxrcrdKwgLv8QWYVXhg
PGJJdkW9U+3euucduoNPbf+Oo7WGt9zOb6m7VgXnc+P6DFUt0hCf+FFFN1a3
21XhykdLUUFlqJcJOMT44iOJ2a8aM+DTRkzHnDYjtEe3w0qTKfEwa5JZ9jzH
RRQRb3bbdhV5spO2UCnA7npr3F1AII9fO/KrSXuOQZfoqS0X7ARqvwj2Ckel
x0Tz9AtYA1MGG1EF9+nb12xdiSQGCIRp5Bm/J+xTT2FXJ84WTdC4K8wLtr22
dWhjxj+UpwDCXxWD64lwd+YlofhWUOgvI6oL+13KZ+yz1hCYwuSgc38lZZAl
ofVnGkhSGCo8+BILbhiYEVLiFCDg3BA9RaGrG38LuCagc8yIz1H2NM0GVjrp
QTkxhNC3dwr1qBC3YQGIguy14D/d2CL4R+kSRyd3vo4IuKX+GOfm4jyKX2kM
ZiV/zy1Ch94Rq9Os6tnI1DbwiQQFEwtUI93TlMsCqaQfQJFoPuWAyFq9X27E
0j/WEOZRIdsj3IgrN6G/dHP99LjyhnxAoKMSOjO8db0ZrqLZNRFXzLbhtZyz
L9yhKAQS/hqG6jvCogUCz3T0S+nCNoV1lFVviRut4HRaERy6aVL7a18KlWpN
p1COJmEUwb4Nz0GcjQrYHpcGhXg6kUiFRvukl+wY6OQsHYVqinocAq6Fu4Ne
dXrgHcn6kqjSxwfdO5qDEZI1mvrvvGHEvB9Mqr5qqzseReli8ZIdFsSNLen+
ZSLA3aBQuaoE8i98VVgWqcPJFZSUNG6gB173nhgPKgT3JW4PvsPP31ITY/K+
CaFMQwny8JmZ7YbmjBJImtDYTQO5SmPMUlRLEftptjIYyVlOolu+wY1RiS0i
xzAzmxSu8e0eo+0y0Fbw6QbFCvRfsCj7WCy3q9oucCN1N+9Bv9CeagwnEmZt
4a4P/SkOxBa7+tzFQ/ThH/Nxf1aUvW1EBCm6zYgAa0HKY9KqgCBXSzD4+AKY
IW2HztP2afOxvNTVq85H+jedNFtfobHcA3clEALqXL7D6DxIisN39oyRI/+o
yTguR/+82f5Qf5pc+bO/QXUrNliJFMALvxMcnZk567QKy1hMFkGtPoTTBU8u
Y6hteW5mpEidkc2GPZwLTpEVhRQ64lVjWzAbgqM85AMf8EOR5Md6DpYLGB3o
dkFgvFfvDWj4uutsUAWEN2dzlPCPcwV36rN3Fdp4bMxKxpPGIafW8FA1MDpM
7NPlZZzPgGBMojv8x9vAjYepG4bdWBPEC9yYMutRw/rtamyz1dstF7tPxfWL
hSZisDQvIWOUo+vsxgnFDjzJmGPMrtybPkfWNeBt3fnK1/cTCq/bQtn71ppe
IvBzPh7YpHMFqTAjd7beekn2EGMZJQiwBhluLyDfwwrNauSi0r+xFKcZOiUw
jpZdGhucLwHibeeokpDb6uOt/pBCItwQ5TPD1UHM7EqkTg27zAopcJEmTk9D
4fh11mbTEZZtUE4O4AC0RemmIKeBJ4m+1V7PUIiFYYAvabXRbBTUOjbR4L1N
Y0/DJDaX5gDpvOw6vjMuY59X4K92SVCPIyaRCczSy/qy7XUnMuq9uYE5QBsi
AP3DMdBxmAorA8rwUpTx5i9WUodIa2RmWKQjIWj4/6+JiVj1zZU4Echur8S9
oLvUGA4J4ynkuv4noxYpesWUHYws6byVM7tbxAhSgCFQ1b1FR9knMm10mlZG
R11cQMQc2H4fOo2lDgPMa17xMQcnH/AESBkF2Gz2k07E/+NM5OgRWipQSD4h
65mKwk3pcQi03k+B1c1O7fVr0oFws29cBQGfkS//Tn9A79C3bZUdWmW/2nLc
wtroBi3lELHm3xPsqC8uZF5LOHhMfkkFzKAMwOzOa1yYG0lvc6KE62Hf3uV+
i0Fuc1u3gVVCyP/NmOCZvyWXmTLnb61j5IMNjsJyH6JQTmVJAWj6mEgtVgkf
mZjxv9E/nIjaIMcPlx3fLDOWxYvbDGVXgb/oj2tsjqTIVaR2tgaR7+Vyg8Ld
Pnk+h7Q1hcX63IeaCho8cRsp+ApzeyD1vIHo++VX/f1E6fCLAy/Kp572zgJp
wqOCpMiq/9rUy6rtmNGt19/v1qYQQwqLuftnFajmisnnuxCqztlOtdUDWPxX
uB0QBqLjQvOKzEQRkBuAa01yFRN/68+HZ5EIIKQb4maPi2oZzUL4rLISNgcD
ghQVG2imEuYNipOmeN79+qYlsp2eyLI5CAY3zCnJPl5em2Zq54ise8h6UlYh
WugJUZJU/Wlt7GiTZUZ649paLjxh/up1W2Zc+sBtHpK+ovXfk1h/SOkGDEXE
MXYy/Xp8xjCh85oRtUwCSFh8sJJNXbQyotEINTaRjItXmN/RdlmDTTEKY6pW
Fc7+aCAbiCsIJbXqrxxiQ8/0+RZtSjXnTTGfSGj1o+v3xGhPfmT2MHaKtIKx
H/0XrQkRtCkCUadU5qTMXBRz9nb2RsRb3ZxWHRNhB0MfAGFfXjqEcMqysCXh
WIUJaTbi+G66dIAwY8n6baD2O4wikavg7/CyUCndbPOFrrVVt9bauQgQAGdh
9vPg25s8NX+OKSexT72LgfBsSJxALyxwj4QLO4cmsaY6624V2LffqvB6GiDk
CaGdzV7om8uCP9u7gS58sNJYQBV8pkfnzYzIuIrlpOpLsV/EV/1mBBs1rhUL
Zp5BjwFsyZDwNPsLsGEGOKKbswpBhO5My7IWbzieC5NKzMsYDk9tsr/L3tq7
WvgnQVqqw5u7YXtUV4GiY/q1GR6b+xUwgdUChUb5BbrDVY+Qrm7W7uWsgl8p
ggnZftlCbtRjvrhhZY8sgznPOZrBRn6okUZR85b+C9IqZPhfIdoNNi+aWlKr
CNRZd+pa0thn28S/l7qtAM29x/kifrllDThHPMW8+5dk8cNbra7Urf4J5k5a
G4jskZEpMtmQUDOYArykku4zAgxsvtjQQltd0ZYIo7JlzXHTu1gof+O5Pv3t
zLlMSqIlMmDW4xUPk1OC6Su0sOP19eaGCrRKZ9sHxGeKqdZ3T56LZrQ6s5hq
1D6r6njclxK/McTLmHhQIPfJoeLgePI6MgfVC2N3g4iISH9lXyeu9V0uvqGb
1vcDPHOsnqcb2Hszfx/SR8KUVHMYhkoLMIyYepCl2gr8n/ADgUqhzVC6Ssbb
/CXDDSXHI2TMiyVyIx1ddHCZbj1EHQMG+Zpr0cDrZjH2GvW5olbwzDZG+uoW
mVmdP1vWDUGFmO1ShU+CIDAH/fg6gAW4rpwUsCocRXQ5lte1eHRPL5e2bFqL
Q0WeIgfeOmMexuEMB+LUBoqkSbK3xo2ewx0jnNhm0isI0rctPtDv/rRnth9Q
Rt36GP7fGxgUJYyW8UqcT1WC5LBoqGI0v6LFF1dpZIPkGNEpWoSqssfLbCvj
Bapxu68mniCDnaCar1juqFqrg/5jc5DPid9nkX2fF54s7O4+3NVvcY7tCJpG
+rQRjTPegII226O7WpthEU3+qHvzBbzJJAhbO6FZabscEaUeMA09uhqrSjnZ
cZF8gRIQ0YNenVQCRBbgbBkl7qIjWLuvlfE3icxBV47PCN+MwUe25odkcsoK
2G5hUlsFM7WbQgi23qfHTN4wYPAPNLztpHuejJkiM0YspWBztqX9m5ECY9nK
/HfLoxMsmWevi/LacAfvrNSESPE5u6oObCO3HQp5+yaOYW59NY1pc6FawxIh
fJQmnONCjxRHgn88N7sJZXizGc9UnajiAKsA3NW+CAFzFZjw0Wv5z4olTbEJ
8hlGJUa+5iFKaBJO/MBBYezJ6sv7r54pznevaENoURtbQE3a1hAGqI1cYD96
ZVrvltWNUccPI3eLTLqA7xxuNVQZ38VHADdiXGcsRa2MxhxQxDviiDvq9+i3
jfCrZWarDxVtMolzSxN2gHPgEc9Yn1Od/Yw8snEsygykgfKJF61pDzNHj6tm
Rn7NqL9a/l5jhyckPLSlaxhwDwL0AlwUXHokuyZb4ZATqfLymzPTj+eVzwq0
jzoDYfDn9l30y6SNfgrF9+UTGCxHzFrzoHJxfcA1+xqKo1NQ1z6b3L43ifFn
0jciMk8450Id47BsGa4lx9tlQujCKcO0OBnpChn3jOa9XiU9md2ZzsIL+YHH
mRG0fKzchrtQGkcy4q2Wm7cLOmjZLqMHKP6Ph7lTvP98wo5Bh04g7KpGfaQ1
jjpXPm4kpZYkdAoZNYn2FBmTbjADanpS46hM892NnwDah7DoUiP3YKHvGwxc
Q3QzjQeqacL0t8j567EkDUAKEgXS/TfxKZlfSCDdp97g/tcP4F4zby4DtuDD
WtWJreMkLE9YkqkjSvpllDf3hG4YEkKhi24B2EXtRH+1pa2P5E8wiU39Acqo
F29v0nKZ2NRg8UmVuBwrrvUwsgorEKqznX1LEDZUmerEvV7VJfMl+TaPGQg8
5qM0ZSuMHsY+yS201QQ9B0cRQjLcXD+2ALo3dKZ3myT7cKspyCvaA7hH0Lzu
W5WTB0RRgnBfxDHBreYGMdpdLmuaZC7au9xI30atLpgYtEcKieA/CJTtWleg
yh1modf0bfavViBEWO4GEiY/XczGdvONwSVZux7+zvG+NHJoPZ62xPQY33V+
NRZidINDT+hNSAn3F5exHtNCwr2yuq6DtS0XDfhfKSW1/M+n1HqRB7lIEKMc
idzrDgDOg1bshT5FCjrOzEb9gvwnqCg6c4R3mTysj2dxebpPdUq+VqP78zHZ
/5xzOWv4FPZTp5R+YIa01MrujojRsPZK08WjGTsxLjK0q1kwW4b7p4Vpjuni
qwKgemnpa5nW84lQxxDq+nNjdxWDemyat3E9q2sHNuNaUxnZ4MpSGAj6K/Vu
CqFuc20CANAzmFReATUCUKlvDI8h1ULeCwxoiUu3Kkfn1rleHkAWDkPI4qPP
5VWRDqMXudbQgJtXLN2THwEhtKp7pdQYPJ2QuPsZCKmMBFY8715rMsPS0cqD
0BXaFAqmfQUPSeyLDIwVDWi7l+I2QCy25ait4XqCkgelirb6tIwpgYvF3VC3
b1us4bkQSvvhYJN6zRkBZBKjQ+qEEBPVQd8UtZ2Kc9qtLTgUfiNl9kIkp0gE
mnh1Gue30lhwVhWoL8dbvo+PAbOA6Z1I0oWMni7MoQv8ZS2j/SKZoJEyn2UM
wFZawUv3nwJfzzS/cUGkC9KFXeOJHQDR4RS0TNS56b1FAgu1E4j2QmAKw9QG
ET7kcWs0GJHCQKYg8hTMw87zz+G7cDmrIVmS67Ph2kZXu1YJhzFLDyUn2wCX
Rx7brJX3qdRPxzd1MrC9kPgR727Z7NObEixuQZgDurrYQTnYOobanINyU5ZU
SEbAk27//47qoUfPTafLLzqLgwfHLH1HraqlEDSS8xJRCfVgzVveuk9+srpx
6G4WadvyxW4NepYrjw9WBCXDZ9Ini+tHdwC8Fd2OAsig7aQvj/KiNYIh6fR9
IBnGsA+e84NuddXRoOlm9tfRfBx9Kpfh1KtOTbk+Es0eAj/WRiQFNkJ4dN9X
7ZdwU8ErBEdUYx0epNep103j/BvU12Flj1DLFgY0tmDcMwnPJ2xXZ5kJXstn
dXBDqgGElRllSv35KzbI2NxpukLJ95hPsi8skmYVINOumXPYVmcl0cPVg9Gy
AkglVYdSYbjN6NwcIZJQBA7iiyJfFXAFQUPWxbWGAtvswWdwgL9zep4jbxpA
ZguwIYwH6o9n0XBFgRe2nATvUco5kx82cfTS0A8HokKVIiQkP+i7NW9ZBIN9
MueXyA2k0f/WvVS2MHd4In9x9kzzCqnz72NupOj+czfnYJ5QoJczX/M7Gj4T
D6x3C6hZUnNWQxhFJIs9t/8m4PeCi/ptt/DJYNM2yUmYgloy69IVhuxfeAgn
FpJgoEuXnMbncKsjn0VUj/QeHEfoDbE5aVDdK47GlBn+PjItPvlq4ChSxBO1
p3RXUXSei0PPPCylO57pEa6JNtXvRBoV1dmLGGSwJFSH0patK3xdnaE8DZk5
4KUxJAYf3Y8oJTFnZ7avy5osa8vly4BkYHVNyPZFoInijBgDRAd+MidZerTq
sqraeM80TmfAV7DqLbBhcS4kdKvck7Xv4kGpUStxbSWKbx8NXADKlnRDGOWk
TmSWqMA0m73YKf7kF7q7MYH3obvZZP9oFikvE+v3E92FAWQKvOvTCJRSQwgs
xGVqUiDIdoso3Iao8PRrV+/Kz2J/OPXhreXtakiw/2Uor+8GDcC4PWqxUXNT
hVV5Ri2IY+Q829dUqzs3BOYi/56XhNDVurjM0eRLcSYbELZ0e4p+lUL2VK35
9A1H2E1gYc1fRr2fFH68uan5FNS8UkAdLSt+M00hq7fZzj42Fn61F77AwAOf
Wmf30OWugneCkfi3zgiIbRCY3bpE2bHIX1DIue2O5HJSFRLskxElTRiEELYh
lT1dz5uXPytkz3k8VVusTLYLFTGdvWHKslYb+jwUtxJJEVcYQ4X4r2NNoChV
mTZakrp+I9iXddY3aghG63Av/5/6oc7QQbu006BerNegRF441h7Fusvyw4y1
C+6b3kOh7B2GyQljnidFhia5iq9hl4rvpfirVNUuCzTRBc20SmQo/gIh3F0o
02oH3n+Np9L9WVZEzLSEVllEEbehkgB629ITtfATfVxgpKU+Zh5grfqg9hkq
KG431AoCq9LSQZBvxA5inmcTAhugtyKrT1Vj6879+HQjWmj2RKj8K6Zs+1h3
liTIdegE7uON9rZ9KM1KcUAZIr+98TeTwBye+Gq48WCijHq9l4ksbMFjS3qF
kaTG1aymt+ptTNi2VTR+7Y4GIdH9bmhiTnX3wqzMfwgVXLdz9vLsplknNsIh
VwzCv397dSaXBSAcGhEf+4dZYt3UWQrAry+1b6EUiXHWMI5KX21PMnzDPTjJ
BEvpz+FsCevRwb/dmNIAkSpkHU2DfYkyxW2n6kc065LOP+KYY9WkOGwEoDQK
dWQEPHZrwtiTSKC1PC7XObKobOVNTmkpNbyNHCR7b+gIUzRFgs7ZV91cnbFd
FYOemy2vZsO1rL6McSSmPyc+fuNGI4oxjlGta4vp+J0071mTDMPhbd1O4Tnd
wFPl8hPpLTv2iYLZBVC/JaElWIQUOsGN0WExkIK63LSKI+gTS5Ay8S69Xj2p
YF021+gFBSlz25L5pAtjoQ21twQifM2DRp9GUlCOee5pm2UMZWG0AMjruEzA
6Hlaz05/zlAJiN6GpSPabyrETYoPOpK+QK3iUepYG2k+kT4pT9eV591feBNP
7fpnARHmOxZR4r4Pjvc65pBlClZuGPbeSR2abNOY5UYU2PXlKE4Qg5LOmD87
tvGqV4m9OHsxvNu6ayNq1bbwUmlx9sYyWj1BkyEgnOHSIfAo8l7rWnYZCFTt
6/BBGOaxfUGIiE7Di7Ov8Vpdpqs7WJBPgA/FfKRK5fsvAoGvbBzz08EDkYeD
zNovoA+vsM0l79uAmmT2lDxf2UU7k00Zsx7wEtEpygsEpAEqgqpXfyLwtuQn
bhzsu4Lx/EDbSZvtCHSyypABQtndJa11sDZZA+5R8u5VMkdU1ggHRVh8/Zz1
q72NiquUR90SnIGuiqi3D7Jw3JOs6eiqWAu1v712x1GDNN12Ey2I4cGXy7sA
I6RgCK+h4ZGjvFQgHSpVs8bscAqwtdFfgilCQeXETozirFRGyF8YJmvSzY3p
g0qBnv3r4bnOruwJ6gaFuh0zP0Sjt0OsAMUBGPPmJna2ETnkorUrQL/OojoO
HwBD74l7/Szh2vczNmXcn4rwcMiXSupLl7suQEROdSm379GckBI/7BQwWHm0
A99oc8UY0wBxt9p5hNczVWmY6nJaQmPIY9MnmkunpDGQ9c27JG9E1Czz9Hu/
Z/00QGEy1gg/k/GxcTHlyZx8hQ8G2s2r7NEa40hJr/ZNPe4RDBCukRkv8K+0
Tz0aqY6i23APiZ1LoWrgIgVfvtMKOTkyZRK7dHu8X8mb0LOd7xAYUIetItGA
0ZYDAjFqB+Nc1NpE9qXXdlW3MvA8sfZNFyUfWJA8N/ac6tVpCJyEwgj6LrYf
7YSKMmbI2cIZeKSQitsbGSpl0oB9N+FQio4owNv5J6FhF7SnSguWpAQ6SykM
geMfp7vNRC+DS1/4XWccz8n9ks+kFCwMWUKAn8Mh5XrxIDG4u7E23dT8JXid
cXB+vaTLcQWcuT1yBnh2Ip/V4FKFHYE7VwQ2znVsBpPw1Uw2ay9ysskQKO8p
6//j80ag5ndnbBE3bbFlpVqW4NsbnqNd4uFidosoa1MtCgPHI9dRxRnlt8hl
goByc45LlOmZ3k+yL+4q7IC1VkL/JHuw/FF+V30d9rMMGSrwTaR/yqz0dmvN
MlsmZYR2qxOntB6eE+PhWhu1Fb7kb4GvIcyWvvHMj+v/4k29aC+O5vNWJKn8
97rraFro4DZzOZDXNhUd3hYDY5lGog5xG0Qm/k3p2z5Atu5YwFVgsjLAu175
jn9Rhj7BwxL54fYUvZVPwkoYVJ7r2Dv4peWKqafHOPwZtyfKT0tMg4zSpFnk
2GSTfISjxeW+NOtBQ4L0Ezvq1HX7Qa0Ch9yHNx7fzpMMPms2Y7j52LnFpdBH
FDp4S2QcagGicLYx4q6Piu5JHZare9xqa9nYB853GRtkkkPHQlNTd3hETybg
BC4aur5g1rXhbnmwEKQLGUAan1ClZUXG1L/uBXTcXY1kpP85pLMGszSv9SGe
YGPxavmxMOEj0OJz2vbkAkbj1aKM44jYBGohv1tVbDOyXpcI69WXeoRnWlj5
DZyph9ihirx2i4QsCpDFqKTan50TiNMDbEQy2iwYv+vgkzymCQcXnS4/pUkk
Y/p0qlcsUl/Ffs1B8C7MZA0T1zc2ybPJgW/ajjyb82XhhmU1BvtYevTVUvuT
hAXYbGAfe2zVS+rQpYpIj5iSniGhrmRNJdeN8RXRw3ISrA/5GMMFLACsjfJA
IkyO++mmbAZxGkN7iwTjtkTuDMLCVYQDNOs9/og2AtZNSkfSaDLqdPpQn/vn
xsTz5QWZmhjuoPbEEkWhZ8+1URM4cVc+/TXiQQx7fuiMk9RQVioQsw7e5hWf
z6GTaAdfE+ytuohXuv4q9+PQM2LD9nRClaYKZOiHM0STszfq0dmu7tbyQSEz
u6JKdQWo5AhnM7/Q4zK3I3mWEwTITKwxXE3zYG2Ci7BWit8TQ0wVD2ou2Lhd
wUVPbba71gbV9Y0MoWGOEYm0MoHPvPXjO7CNdpcjLlTHf7hGdURUjk7htjgA
XlL/adYGhlgfmNfCk3fMCw4MrVVIFH7w5sVkgf5V63C40t/Rt1gucKGUJkis
7NEC6HMI/XlA3vjRD327r2mQQv3nwE50Q6icOwGGkyezSepNxqS7doXsOY7K
cwD++YK+/PIzAHJQYF6rTAA72O1nhC2+um0ARdkBSV0xBwgS+sZuo4qBvxg4
UHcaaoILArUbRj2pOWvp/vWFdVNlwHp+sB1MMm9l9jCaM83zqoxoRXrU39QW
93p9AJHH2sM9/YtiTioQ5oj23DLYwOOiqLpDlweGcuoo49TyOEDTMbk5D1e5
XCOPlP3pVFDstUGwhfOfb6ZQ09+yuZGuGFoUk1O3Md01CtUs85NUiRjvhfGl
S/9SpFM3QxPsYqS2rQP8NTiVYC3IK2c25DuVPfKPEHQeC6rEtmmIMhd+1Gnd
VqDjrOZXdKDwC3FLcHDZ10tRQwUhIe5c6rXTIZ+EjqgcQ+DqZfwQL9SQ9oyz
oFq5++Wgl+lOBPXzYWBOjuh84WOsBXSOPkQali+c6BSf7aRhgRcB1gQF8IIV
1qATmaAsSrr55s3Y9iua/KvC5UBprBawmDuC+kXDX/C9TvZBXpxniqxj9Fxw
AhaEzoc+xsRY8R/GZCNck+RucXBP1KbBnNO+1io4pmMNdGJJablBa260lRtq
j5BTGg+7bn12UjdzHfERAg8djEf//Q9Sr7G4SNX7ay/tvTKGCHmBtIL6VJKx
fDLafv+xOoxE5Y+D7h02qqpBNvOe7SGiKPx+Hh7DHG+9Ap3q0xyi78WLEgex
HVC8jpmT01OeIPIA947APxv9/i3unhCtYk6G/CFtIgKPNHv7XopV6VP0NWFm
tjck30H9GCGcDLjqXhliGIV/MF4a5SBzuxGknkdrN+yB0BYWtKmaGmoC3EEu
vIGGFrh3st5HE6A4vWN9id47KyMYCoXtoqISQabJ5jbLMPr5GvNOnaOojp0d
IuPnBNXLRgsjK3GQ5c/Hv+a7kCsBmjp1cj2O+pTxite79XbzzS3vu+DWct8T
2UBL2uYf3LdywkdQkin+ZDxQnP79dusJnEDSghWuATCN0qUcTSmQGJShCb5C
QXz1VzYrEVOouXzcXvY9U3MgLUxGmJ2SuLLfRw+RXt2dXBl57QHpqNO0wWzy
deU51C+3v8ocFxikjhOWrUV/ahTnc1MvJ8cH+EjIkQFiVHyPjpuKBerph32D
u+dTXTLnV2GvCp1ykM0t8frdS+VEXkev5+72pVP5g7ujoHO9JIkdo0qFH/tc
qjs44gd07nUK0qzLW9gNgEabhQMWvG5P9zHmwpPZCQiJiv750qkGGcUXPWBe
QsfgEAVZqqNkLiSE4BFimwEnpcVDyzsac8EY6MEz44CySIP7kIQ8va7Itonn
hNljkuo5WI8ckC+pgO2rJ2IH25YMXN4fojIEyBnabgoLy8QQMtwwr7C8XV7T
zt7X4Zgbp3h0zCYomAmkpV9Ih9wjJO/zVrdaBBEjZJ6YqKQnLhSCE8fE64PK
NmEhkq1icxySE4UmNoLpLy4xi4zoCT5A9cXYPg9SszMNc3kUyzH2pmLl0yCS
BdFpNG6gGF66dLOEhwtw9j+xvAmzONcM+FETGUBnH4COxgTyJxQ+lvgTepW1
QnWzorHty6qfAsg4+aWiV1gaxkbSNovMgGynF2usL3PXFvM6QahU9V+z8DNQ
KtvOlxn+oc4CJGo1ZkAoG9sdTlgNM90d9rAmkd5nQB2mEs8N3eD/pahYNNVG
ZJDn6ZrvtX5q/Xm/qVKMFERgejgtWj3ww08knuD+a0E2CikY6r+V8+m3KVrX
vk/J/Ok2GKRZwAyXOt5toIuG5NMnh7lseFpcoYZErrOnU7rdQiclDsHBfarP
ZYM+67sGJZ7t47sehTvCfTohJMjQxB0/Htr30vbPG3l/Neekk80vkJu35Zvy
Tu9OMPt3a32USA8zoY1Udg2wlaDuKwPcVL/x3L3PkU/s8aO++rNOdX8Jqp/b
IEcpiKAJCmcT8qqCgP+pirx1dzzbYpVn8tJ+o1D2zaWpeQ+9dCkspdaHv0Ir
t0aqCF/kQOOEZSTolr3h2XJ+9ar6W/tf3iJ7uK5DxgMHSZapMzCZoiocifHQ
6lKGZiUBUf4CQtVcLcn4pHwXQvgLvPJK1Bvf5WFFVfYB8V1wOcvmYYO9jtgH
NgQWnwXW7klFvLa647H7iUnNMeyuAEd2SMI8gIMLl27s/w7z8tSRodKhTiKt
dGUtlLCdDaJngL++1rpfPwMHIR9v46vaN41ztLpp8Q3jlcJBOhzsy9A3m6Ff
iyhfrwXR0zPybVg9YlN94ZlB7SfaUUnSwU127jNmnzU/E3AxN8WsoX974i7y
wQUHBcEROZH3h7dGatwd8r5vvDqb6Ik2wd+G49P4ZdqPH9NHLFTZcL0y/jac
DEd60tuHBqXA6qNjJtLnzIhG/brbzuSUw/PCy5lQS7kFkEImwbN+1emT5V+w
PGrazIqaBHi3ZodtxdhIdcQJD7xBYPDa+JXKQDu1OjXdR71r/np5bzoB25j1
4EheN71KAJaW84OXxVRbkrL1mV/oKrzuxYc964HO+rVh6yt/m4BdBR2tDvif
DMCjO9u4Yc11Y/Mo+sC0l89m2gJiSCCSczoZNz8fMpAe3gF8TSA5H6EtsHY8
oSckfXN07VFzYnTk7UpEhwYsXQwI35aPx1fGmhUTX28YTcKM0Kq+QIW+42ra
iAW7jcRkKtt5HMi7qaGBUxioUO5JFSoUF0n4+J6HHJncmv4+5C5hh8PaBk2S
ssegDSG6Tdio5iX1N2FNUqKZunxLdqLlu6ULO0RHqeR+D3vA4rgsZ0B+5CNZ
zFM9oMl3aOxSuP0Xh/ySbppGmic3h7lxdkeZh8YQBhqUT1jZb1fUpV2LAl4d
Zf6+wSvtEx+R2xPtiPU8/3W+99YOKSgN9eTJaLqbB12kIdHRSWMP3oDFJbof
KzxeKRcq27ax67IsU/loMqUj/Z0E9+k+KBJr4dfsfl3TTEu6cttx39tkuNFn
lPFk6sUHDRVIevTD/iwQHXULqfxhIIG6pSCnjavydZ0kXTNLtTuqDYEM9glG
tum+tNkXJfN9Q56aOZ8sK3pOz5o+EKqminOeRhIzAusZ5djML9aLnXLmcPRF
5XEQ+DI70C/HL1P9fwEs2yWMNqmx7+3V4c6aOCu7nVCBqYoiTVM+Qn9hknpf
aj9ZznFJf5yUAJw6inIQMUD88haq0g16mg78OidKXPWpENgFsvr2HZGCHNyU
pETCaouxIOgdOqXqqerEH3L5ShKL3haaGwJmfXXhRMsUMjfEJUBze1tgTwBZ
ZCuMeW0J62pc6YyNUieoybvFqhaGEDsOMVqOtWn7KNXnkL40UlnR3+wC8q4C
lwG2OQYlmFrt0uYyls63C8D6PkSKkN60nMi7oYR/s1Oug++DMLaQtx9WZSNU
2UTKccjxhmnMOUSk+Ia4YNwxl70W5RssYmv+lpS30XAxhJr2Mtp5kX9jsrEQ
8/V3R7SBF+m/HOEszE6kW77dXGl15hEzrYvbyRcQvXogvCx1h4HFgQpludlA
syreAxehKiL5dan8veao0bbSODrXJfL1y8H76NHXX7cgJoXc0p4pSRKcOwxf
Q/RYh+pL/FMy1FQUrBCgcv759CFdvDG1qEXhoPhh1jsNMRQl55eQ3/MRVhNN
3YPinRhJVVeeV9zqqeFTAGN42eXtZ0KIL34+01c21eM6U6W647XMsrWJlFTw
b6JH8nspmIbOJX1QX5tDAkJY8Jff5DuEBWvAjqhI8+qUobGh56Ms/sBzqY/f
8hDgkI3xArjEc0MZJZ81L6tumpPK5KMYVm+/7IoFlVspNireiAjN/ePx2jbF
pgqFMB42bRA3aqrh+2SwoO5GNYcrizbNgWd0z0Nig75Uwh27B1/vgN6UXFOJ
Y2IhY0YylIGlzob1SDUpnwnDTmYM+3NzbdydTRvpnnnhHLfT6QaoZ8sRwGjX
30CX0KXuAtmhc0yl1X/2FVXgs1eUM6qE4iTe23RO1A7YdN22zEQAga/78kpt
f367pqZbzARtv0P0tmyi9zs/jKPlK0BXyS4o+GKYmZQA+uRIxViZOqdoVyB4
ZdEznWW4Ig7NpfGDhvZnZ8REcPKXHEtv+CspEA12OPsVkchKXg+aW10hPYwM
AvJoE/SfqvakpmAFNbV/IpeXZYqQhm5Ila3rwEjMuZJj6sT7SbHiOfb657H3
NpnZZU67vjVF7bWDmuOxb7fN03kiTPfAXUC+LU6PlUwU2VyGbD0Wa3pm5bzh
uFNMKEI0q6AvWTrCP4lUaU0TDZopEs4NUHALpiH0LyQI7Bapm0YWZ2cqjyY4
M0wMeLp0StYgFqJ3gPPtB+4xa3mxgcAAHFg8Mho/XMrUDzlz1AF1zv4PqcjS
gMDk32t5vRj0rYwC/uaI6IkqcKaR5RfGmRDlLaHglaa41RoVrT78TZXNTRxS
iRzXIdxkjP7jMmFRsUuEL+r1iFN6v4wCIwgOhPUcqq1iRSNG2r+EvKjwKrnO
EMQ6Ih4VMgDlv26oziR24bETyvNvjrw0tilB6HPxYP5i1nu2ftj+xs2hAqYA
OyXR+NM+I38wzBNWGY7Ly6NqNW7A/wc5+/De1DNaZoSq8++jvqGwaiql5+k0
wat1CoFHK+syGgeCjUfOr9RVNxWONvHfIOzG//sSTH2/tBuQYRAbF6V44myp
Hze5foxcrvw3XmNWZnDXqgcuVVo73sCEdoD4Lf3DSpTChX3KyzaTmvnrnOre
7Nmgr5QJQRv3DFJAzbUEE3pkI/9OlLyD4eeRXLTmz3+22Al48Lnzs6HVA4Bf
/ycUrCh8qo4thz3ZvKJi8jYucNwlLnCcYEsO1dQfF9QQSfOCg7MIVPgB5Wvu
XMMsPFzYa/GFKsWaHb34lNYuD4aIbE/RoCPPdtJxtDTPAmBYNlz1b4d+1UVL
emfsfU/PR5R0m32NHmAksVjOBtq8HxvBJLn5F7ep+yyYm9s0+hQwN2TrrZeI
s0X4QtzDLJ9iyYTReHce1/NGMAHUVppKCv+1UtYv19cjqh9T5JubMvLKCGS4
0XFrcKsOwfC1IiD7f6uVVil1RMPSLl0AqDgEOJ3+4EqZt9iL3Fgro+nCElDe
3QGMpOXsljdWgyvvfRTcLOGqSQLINDf5zLb8pieJrGYisuanNC0KpxkivTkv
cMGfwcFEilo7TpxBI32xzE+J9Ns6O/5uCFrynnRtqAAKZIjkGVlq8qT5HG0x
bK0ZBoNbIKEr7hXyzbyu9ZmV7kSrwDxNrpccZG59UjtfFv4VmCnC+5e2zRLy
dQsTff7Fw8pNmI0Bsr0kSOPZq+t7TxwQw9AC3EDqa9b+zrTALBEMACNnfeqX
GjqKBJoaFwOK39b6JTliQyY9Nfjxw8UM5dapjJBROXzTdB/muH1Y2xd/8jRj
fFbGkh8X58D31jQb3z5k7dmTxo2sn9c/DeOQE45S+iTYrSgZZqB0HYFVpnNz
ti3BQ/RT01YrWcc0rWshT7ZTuLwPgcxbLE9rgvQHQwf1q4/ZP26uun92Qurb
XgRsBuV2uf4GuCLgfDtJDFt9+8dlw/IYkPKPtyEXScDMxVQ0IsMezDviQTyn
WUQzbO5L8UxmzifAHAZjm499X/HdhF7cYyhAe9R/js6n21kHlAlToVQyr1B1
v4c6oerdffDuK5zJpaq6jt0ilKtgsujgDrEnCWXM6mlrjj/iG4OeXYHDAsYc
V0SBSAhPhI+FdijeXi4GGlRvRi4f2VG7cztN1kM6wCREOnIY3QbiPDdyx/Np
VsQREja0vxFvPm1xgvgT00rNr9CfzDMzeYoqeWjxnEGU6q/unGpU5d9jswlw
kqFfis3/lW6ouea9Aoermkz2PkXtZVf42t3+C81eFNnagiinpj+qhBpzw4dO
otDBzPrLVwCBz6CHAbKY5qcJ9u+nsqNIjMhTLw3xSNrfaXQyYhqRgKwbpssl
u7bvlyarnJog9cofnXZqC8jaKTO7hQo+iPrjrfwJLPXtGId7v3/8t0WdNvy2
sN4kRul8CbIwGeLvXOjwI43L74HsNwbnExb0q06sI6mS3P8/zXNNmN18mZ3O
JAMeIOd23l3wXNT3Bh9bE+rplWbjJ+9AAfynEGsGE7oZZDlZe/hRLS3J0jEL
jbN6deOZ2Nk2VYW1uknmuErpxtyd9bjuaHf/acPGcZQOHICVZC5aBtL+NfhD
LRqJDJXKkbzbFgi8S2vhgbWskcsGlUqY7+cV/slbNmWuSmHl+qf//7nz8Gx7
21/2VXVLN0nCxStVjmLUgVAZr24bJGZpPcdRKfBfDA2SiW87MsKiUa+NOwRZ
mLCm4RSwszrp5uGGsT831RMnPqQUO3Gk1/V6x8QpgGecRDdGk0DSXkzEb25E
COMMSTw7b30doMxARPhz+fLT++yG+itqSYyifLqHJtzyaVQX12G9Ei1LbhFE
6YYbC7Viu93Opg2wDgYYlfhUpJ9ByuwiM5DcyoMQqurQxhHBpGnGBWlTmEDB
wCD6FgnNFBXFEakLQacjsbRHmEyGUdMVtzEF+S7KGSCpBiJ13H6bSkKSt0/O
OQsPou25RdqDOaIiE1vf8DhJTDWecNDzkfWdzQ8hKqNTx8V2a5e1a77O0iik
0vSjqrbPlj7SzRPk32QyYhz4zD5m2B+k3NziCYMICub4vDJk30fsTgQtrgzk
/SAO0ZPCQ4AZ/XFp4dHW85pADI2PSxOX9pMHUpeBUT8D4YJrFiT1mCG7/n1F
AEGqrExUG2dNQreDpnf3Kvk+XKN33mTaBcGWpkhzJ6PXlK80hqBrERDbD2nN
Y80VVnILpeRhvnSbu8ryWlGpskqEbpG7rJB6LEx/NmWkZtjGvKdSvtlNdZMe
7+OHscRWx7c0hMtmdLRq540NTgt+QQLz1jDSNLFgryjSMPyoKVGFiMj2m9Y3
lP2RkOdfBa/KH5yWLkosZ8LDxTQauIgyLkWnZIx8kv0NBByuNtYjxktbthCv
ukpIZ8yovbNNUKZ3ECXmIbY/7GIjKYuCx3vO7BE2tIydNPn3zDvV16MgKr5A
ke2YcuE7+lOvcdV2F3+ePXf0B5/17B3dem39vFOaf89gi1c3E9rFu4iOoWQq
b2h/4N6le5dKYX5JwDARr2ba2XCS5lfXJSje3Pz11BF0x055EOVJKiWslVjK
3RQS90ymptGWtedurGeVE/PmgOLQndKUgbhZmSnrlz47RsE/XnYjfM9g8upQ
PJvi1ne21XaYPa/IdPdF7EdeNTU/yAFTN3DhX/GmDN0FTBITqAPo0HLOs9o0
lx4eHPlOoa8Wp7OqeP66y1ftrrc9DkuVLy5jwtlbynubw+isdaE6OemnUgtD
Ee/wt8Uyz55D25H+G/BLHSkbQR2lf/2/y63skhGO2TafF2SMcq0eW/WAGQkv
apyENa87eAgF8lEG/dfP+qfvGNAEMWUIfIyo9OwuI8/vm18J0wWMNotCo5wL
t2fucSNOKFtpQ2AVHFtfuaUlnAhr4LLi0IHwKpD74NTNKWe2eGx2Fok/AOao
LKhztvVtvizJsrGmIeCJ96Qyp3QDsXoohzcz52gKcguFhCbURV4Q2arnI+oO
UBMSJsf2h+/gH0mfYqsXnCwVNnUnQwvk28cKQf+FjH7nGmYvt5fPMMEjenBT
G8Hm9+6Ej1aDzE2VtK1AHhb6OvYZIWiTRW8cFqOTJN96aej7eDq1WaWDlG7H
QOXBCANcHtp7hkjndJYO757JSn7xhCOusWu7v+v+D2U/FtdCyNubB1YkPmdL
tkXIiArufyi4SWDK0tuqNsuGSoOiGFP34LQDFlFLbSncT4ZEug2jKhtreXBB
jbvrPOX1oEI46wYa3CfrMrxhGbNTFAV2zqR7U3UXCbzt7oT83WI+J95/UYOW
QMG7Nq8OscCg6iZrU8Ec/DD8R8Gz5XKCDI4dvn2HMz2NJPrItoyR+kLtra5Z
OPnUrNM0j+Hxrn8ZXobC8aEp1D01/Qb1zO8kPEbgc1VP1zP3qPeVKcn/fhr8
Ps0BgUuZsn+irIyYoP7b3pIuTb2t6kvrdYwCbpv61Fl2u40iEp6IIi2KWx/J
6+qrzgACHoOZg7NpPYrgbq7mnNt7fRXfNin7SxFC6HHq/EShlveBAED48OPx
XYsNpy+LvCAnY5M5MHf8zTOMmXEM6U05qkMJ0+qZ1024fbIzO42Vd+Mi77uK
JjnDYWHgN89FO4FAuIe/2oFS40401blSVcgKHxIwxFeVyzju4KO91rgCr/7l
OqQpRIsWAdwQBwviCQyZQW1GqPvbVK9j1/5mwAxnYwn41M3wBEn9IkRfRTAf
9N1VmmU0oWgyqY/o0Jlqo/lHCkFUiZ+FnaqNC2dB7Vd/ppK/SdMsZPQ7V+In
HoVKavPSdTMgVS4qwDv139zBO8C+xiGVCVvMRsF4aVnKX3emBznnf5N2LUdt
v9WUJy5uMz5tTsgNJ/Wv+0AFVO7RiQXEjnSWdPY7nx8LEfdwaRX/mdhOzvjs
Mam222P1eqWOm/36IVp3hypWvN5NMaMvnblre7RafIGhIa8u61NLXJeGQJns
rajLIG9KfzRl+5rFr1nlp38mAae/0oKrudzDR6eoJ0v1SF+Sv2P6b5XMWc6c
90Ij0hNjujXiBaMYTddEUGrW7itYNDBIXEbU9mbiVav+CYJzE/XyelP6YtLY
3TvW7N+cTkAH+wK3r+UHJGKGzN41JYBEnchBne/dRLf0kZOGrwc5sJODrfNy
QlbeCuCWh0OiNm8a6M66A6iFb8O04qVUGwF435CGOkbOpueK0DWPjQr3eOw0
hORwQKbwQnl9FKlmuxo+ij8x8yjj/7tvxAAs0OASD+fEnXnWB2Scv5QxRu/f
wMfznGHVNYW4rZbWmo0v16JIFrXi4aJjK5nf7e5b+e0aiR/aT+V86SDtKSQH
A8bgz3WDypaMOOjaMVHGOzwwi9Bm4w0jA7jtKxAhN0mhrjh0H/jYBBxE3oPE
hnJAZgZn7X3q2lmNoeAjkuC0M9mYK3YDp3AgsJGONCLtOvBgdtFa7zuW9w+M
5LB1db2Ux7slzYZGwHvZkF5L9x+p0IdD8+7shXmtY7FVshhdiw7l9Sttjf7S
oAj3VUAMGon/DrG5h8qua25FWWOVRuLUeCIjzwRpTfaO0nCnoUl4r78erqNy
lDQN/HMorUF8aVP2PiXZAEV8YhE5MB3qpnAD6ZaKufXeK2VYpo73ndy0lOvl
LSazzA+Nu25+75GWDwYtFTJt9z3NAo39eaF4j39zxnB8eToDUYXqvfJr2LeJ
kUxnIMPr+0ZSFw/w7UPY0d6to3nUxTVc8nMPnXr+HL0NJv3+6dQ2z4NAvJpV
N/PTTmWz71l8Sn/6bk7boIjatc9Silg+Av2TkVChOB83J46GFmBC35D+cdF8
YLLMe/+BdnSK2S/FZ/n9OkKBr647PdnqGuRSMUWV9WK8pOS9eTEfJpsFtZGF
gw5Ewq+yydP7ZUKj8/gdGMf3uo0lLF4KwuXaM1bPbMerTJvaxt0ximWbgulc
cW7F8s4suxq/XuqqzvSZXLAbl5+KzfP+XMWvhxLluUhbUUGuqFncXBIKM0bL
c82UaE8Xavtdm7pYP/CoS7dkaGZB46hjR+Gqi34DFDRkoK/1StCrZDgTimjq
htS3guJ2HAlX9YHS/h8pEIaF/Yz3mzz7XZonLX1KNdVBRGXBcmepQXPKKWsB
brDo/R0Ga3Mn26wSSuRgSYgANJ4htalubm2hPphX9FN9ffhsna+Ce7YQgBny
lO3YOfQPywizy/6Apx2e9YVPBB0sra5pCrYoOb1jKHmjI6AJl/VxSwG1UdeQ
sgMPGAgKq6+TYODdTO7rbDpTWJ4ZfWO7Dfami0FkgM/E10anroZuzTuDZf+j
NmFu/FgtqKkhlzwqSmRWYn/popiJAX04JB8wIKOoUlCmZalWyH4G3LEWRsmI
vVbeBMSTBXibRfLAC3tj5T2ESsEfclWhu0fow6DdYUPwkBPZebIiGK7R22de
kuaEvIoz2O53mpheSpd8cmljyBW7fT6JIiPVn4sLM18OQp3Za3/yp7KjAcT5
HPg1mSRUL0ViO4WfZukP5fXZhv431RoXrBzENewRjdBpkAGqWhLKsvBB6hB9
0SCkvDmYC7VJuFJrq6Egmbq+uUiVP7sDc/49A5mMVV2eYYYOGIqyzZD3X+Jv
tfi+BoMiyBE1yMazfdeHkEAvD4AelwNNf0eciSN7PJ5N5QXa5j9Y3nxuWv0X
ktuN/NMxxkIwGYi/RIkptAhIrLuOE4yOLHchQzMtzWii9KBGqbk1qfKo0X8j
qqM5QQmPuMMiHac6vLpcquvmFmif7pKBpRLY7HBvq9wD4lE1miBSMIi9WNJK
2yw1HibarlODU18Hs7GiziA5Zuo+wKvxPXIlasej4CvLbIjRmYncZR6LODVV
SLyiEwJjbNAmd1dnrygXTgyRC+of8yc6ynofDDxldIA0gxinuhGtoddC5yd/
Ul6N4d1SRnhhGma74T94Jh6xkH/TUvQKD/5m/E5KuA33wzpmiIF5+pjVWx3b
PCfHYWgkNEtg4fUUcfzX7ofNnvYeVdzeh+gMgIZeTJehy6gZUtbpUuB8IzC2
ZTKB4yR/wsnG8unUDew32XGQ9Mr72cacw8EZ0rDgSaE+ibWamFS8rD6at25h
MGRIj6YwS6o/+KnsywCutO47KGpAQuBe5l27/jXuWN48MwjfndK56CZCIMzt
eCdrVxuG/mTmM5cEC22RVe6m2rN34UZuqheA3Mg0qumlUVNUZNYtFHqkhZbr
INxXGnnN6vzgCtVJwFCstDPTT7rYrlAVH8EaKTaQzoDFxxE/rqyC2oElqo6p
+bmezBQfn88GscOnTLBppvwfiDvWacVauM0itej3LGAF1Q5AV/fbwt9hbiDu
wna9nqqwI/1kgP3zEyiuhgzAjz+Pmxkyk8VB45EqH1lKvYx53vHzZpF8V0lm
+2BSqsNuZclUkvKr4n75T4npZTivVIlf64nPzPyLW0lHrH9J8uUYxLIZGhfS
S9ys/lo8x+J0Ry+AU2NXDzXGEWy8Nlo6YUvUjP+8ox3b0ywoFmIWRKaRx05z
4Dy2g2b0KOvVtzqP/91AWFzHVexRp6y7/wts0cXhoO5mna6EpDQC9vW22/10
64qLuvLeIcgNRhyVFmjgijx/NiF6tvyesFnUqcA1hday3kwiYBxLH0atjbOb
jrJBHEhf5mw/DMPA6BTVZ+NPPj+pDgUgIQDICwMxcMOz4LdeGPRzFMenpgcT
U+UI0UR3wDQKB8XMYi/l0eIXOHF7tn2HCw46KB5go6hyOzwVgopsIF6OMP8k
um2YJJnrBHf3sMrRW9tRcEsRfQTpKjK1zDfg2V4dpZq11T+Mtxv27d1hQcSH
p2NbkYwVjJCmElOSmisjx/r3m7anrzjBvcQYqzF+IkvzTDUg6ofC4q7xTW0I
lSIhy+7AQOcQMXCMhMXIhRB0TJrG/b5TE37txGSJNyf9A5JjIjCrf/AMRMr8
Fu2dHnppyp05aZ6zRnboUkOUvaW0LN1PPOXS92kfHY1kQ05ty4NU0dyShtJN
9goC5bs08fV2bEUMk49gN1hSzgvTV9uaUEZtjvgZzBQA5+Tl6IMGSzwBAaCH
j3QoFVj5ZYwlMI8LpuPr3/yTpy02PNRkLRnxw5dPd2w9elyKbaJYFE3pEG8b
hZHE535T21YBOUhXniwn9eXiF9Faz/J0L1DLe6KKZAbkhqzcYbvaCQ7VCwrK
BLM6CTE6RaHOyH5XCNnG0I/XWjCRvP6iRRydMrHKmZto6jZ8wntsCirB5TgC
XLviT40YHpudvwZsR9vNE99e+Bm5o+hVSe+t2W2aOl99F0qQFImtNh9VhUld
DlH3PrZSJTg205bTKUbAgDjONHe9dIVKPPmcA05Tj0QqUBG36ZEilRAFjCOx
i4FOmCmE0UteYFoahmHILNSAnk1UxxymA/P5Pbp9O+Q8idN0hCZbg6C4p1Tq
F/BL4Iazol7IqhCJxoCAuxZZhhGDDx3ZaSZwMsaIkZiid+oGDcqxIP1ZOY0w
7IfHiUHHFdJB1qAjXhL4BA3n+mP496QmZ+bTn8YQapyEVwDUQv9pNgmq/GEc
SYhNjiSow+u9r3QNuwYijfE4fzTQ7MHnDV64uQCaTcwTKxCrNa7isbpgm0kB
dClL0O6zwOBwF5bgQGKWFiPR+z5QOde1YFtYlRT4pQ4i/j+n7Iv3BzrtZwJm
fGBPWtIhFgbYJCRW4Mkgk7vGhOFjfnK/+Elc4teSTmQv86etx49rMHkMoUOf
Nl2+/7V96v44XmFnnP7d2yIBGNAiAcck0Vpw+G426BINB/yndZ9SIb4KV6px
EWJX/PHXrqdtKprzmch131/yv+T2qBaZCyAe5xuV8Q27VSPShUEF2BYKZzbJ
2ANP9XBfchCcTB5tYJYvuP3UBQJUME585bQYruc5Cxuw93FhY6kJf5cPH+b4
q++rzHlY4lI9l64xG0M47+1QtQI/QRZ/dgIacTqLglbnHTsTe/C7EjtreL9I
bw/6Fbp/mUAms2HXIZ33WYvwtOy02vOZQWg7IgOs8m/l/AgatNZIys/Pm7xD
nsL0T8B5amoBmUTX5Y07HFVSqYu05iHL5+nMl5waOIUrH33oN5VC1FVGB1p/
dSW4eE8WQ6V+jiTmYmbPnNBFdn14goW7YvnGfaxAuHpiDXsOGfJ2unZ98tuY
xwIJysMN9tsfrVvOBjbux26052juMqQiT6Nw6j16MEJG+ZLuFgaA9dySrtmY
m4yjgpbYmpi+QQQvpIV6ZZ+ReV5WKJSvlpqVVrdWIoVry5mbb5adNhvVmMpS
tDWNSpe40++kZ6NgfSE/cQKb03RsKQpEW2DAAFBiiwA39yLE3X17auBqaci1
H8LC4mHgwxPbjD+36raFdRJXm9Sa+onEFhfZZCCRiJb2e/HsCym1Tz57/xZs
FCzwOO/OOf4+sDb6v0EgUa0Q0stV1GXh7YmDvE2n49YbLCmhYRbZx+phYPSe
PXoi4mDb+jAABgqAUBuIegvRovN+ZFvflVf5LJKVrf3pggVqf2QUBeXMhzUx
i/yp9p3XC5uAjyOe/TkpUcHSOoedFA8HEYlCvdTzNeJnntAqg8tm8HzkHahL
WJ/oNMXqUs7hq3Az6F24FEz3C0DhbIxuxIBfU/BNnydglL46eKf8qt8n4ZpI
SH9S3u5elL8H4gaNz8Dzu3/RiPrvXTbNvPdaZJjVyPKU00CqKLzvLbluZg8P
QorJXr4Gk+QxF8HHCKY3JXFNmX/PGNLYlaT4DFk8tyDCozfJGcm+p3fSQHqG
Udot2+At7T1rNiHnG3qMNWm3Cxd5EfxyR7CLV4B1huX3hlV+Ip20yOldoCVz
uwh7DM/qWKD63UvwUnsKRQmwrD4JxVGlDzweo3GgMQzYlxZmR3BuMNZMqp/y
WGmEDMOAt5di7iMT9LpxrmpACCYTZG1ONorpc6rQaDyh4qv1oCdhGkLpSl3G
2yvP865Rzf12rsAHqr471nWelZx/GUA6WhZ2fhxQSCN8YDqAdvd05MeXhxOj
xrAkP+amtYGnt+zQJMx1ZbkLi82FJBwQRe+GMaa2l1G7LoC4MbnkXP+908cL
jISc6Jwku+co+2pdb0edTdMl7Bka2F5RftmaIKeMtAGy9054nNg5rpXRy7GO
4C5S7c3qklLRCg4uLdqC2S4SVQYPz9btlNC5kFNBGcsjvwq7jLaljEYQEJq4
GovxF+cz3YUMe8Qd5YctJeJ0s3ESzY9yzT21pIjChH879035qvK0zmJVwBkc
+WKNvJ8Bi+eaZMm9c/P89RATBisWYfC2G/rU0HxB9D65P0M9Y2SAo2rAFXSi
Zf0QDRzUqxCdp7NefiEH0BXAXi2v6fdm/rE5hFMzgGIb5qcfRvu25p/u1Mfk
b6ukGJ41LeXvmDPsqiUhyYRC6s7XkzAWHTyn0H2NPWiaUDq1th9bdVv/Qs7p
r8Heetwn3R8R9Jog1LOtF5gRwOgwKnYRdAN7NDOJayl3oRH3dwxX7FzQ6WGt
LA1ccZ7VW5DWx2DakbR/207gj/RpwGLCkaA1EjUx5Wm9G1R71lHTENL7kgLa
2ONa55F3CrW9N8GVvn20L5fIJexz/XECCoLPGVBuP4lJVC7pES+R7IU1dMpw
EZCnfJindJFCJ2hVZJTtJziHpfBo1RlscHafsFsINs9qaQ4vsdo0iaSWo3dW
gclgzpa/V3qC15+2q3B1peWb7nvByr+oyVN5Tr64Y1KLnSj9UuwP3GVBCIX8
3up3Ly8axL/a4a0RxanY8+5Uzz5BuUo9HN3ze8NZqWhkp5Md1vnCqY3z6Lkv
X+SqIX5y/zA55plIoWK4nzPcz9J7fa3rCdj75/R1/UcHJt+D7Ix8AwTBfeey
4/t36VQXdKGD9h5G5/azhfUTp8QDaJ/CAWkaTAKZGcqny9wP588BD04jcQZu
KqEdFuDJ69UDbqWNXArtWCMJ9XmCY86qrl6hcCGU0nnu0GxJBSiSmSW7wWvn
tu+jbmrsUWBfNlDNJf+qjRkJW35gFftb5MsYVO7LscwV3EcwsU1WlEjKlzWT
SAheX5rQx8zhwQ9UeoKDiImeMTeBkjqU8AsRkTgo6X4eNCsTrEmEnpBA1mh8
vuGJn1Es8uL8Q+JY09jwqzb72DrGGbB9XrhvmKgd3wDHroyswOKP/OF4aLl9
J1iYNEuwNF+9vz9oJcyz/T2D6pWwWebZd8W+0GhikefBaHrruSL4IGQ6z65Z
pu9nHpCo3lU/ryy7uAf1bQxwXDgbYA0dZ+JcQfugFNl41ZYhwSUKWh6OI/fN
JyCVYRm4ITgbp9OELtmFYl/r+2padktI7UbW5kgGhbCuqLgaL9BD1cq4uHmV
Dr8SGMbh0vZ3jm5nP0AOH9x5Ane4c+PXe0cStctj9QZ3EXQRSf7xTh7jCCS9
/kkEX7N/VhHl5GTgsOHIRxTNz6qTbqtZ4/hUMnt5y9S3JeRRRFLLRx19NTvc
Ym0S8ovydPTXb6krwWs89rIYUkHJZK3BSndQNNWnQolhQYiWBnJ5+GFpFWQZ
RhjY2l0i++c4qP5/XO70aDQa4NhK2ZbH6Fs/qjI6+KeNVvnTPW7fLuOAfGPc
MYYmIbYVLlAqjJ6UBBGyNZnNRFeuiOcmeORDPW0p9aUX7Tt+71Dpo7+/jpN+
WxvnPccN+NESGv9sFQxeUwKEaXYYX3yIB/fW5JKV5lhg5zVLt5xe7AqDqDsq
c1mwizoAGGqtS+Fty8gu1Qx/MGYGvCbQAzp85cOi1gE7qQCx5xC2RgpVU+Xy
JzXeL9EwRL00OWTkl+gD9mQ0FY1xCJP8hSsRWNazwuMk+Lubr80qt9ARyKg0
HfJALi2aqJe14nFZVxmJfs+dmQAXwNxjzZd5qksbO5jw6ZbqWxFDnpda6T35
ofYtjKCZQjtctitDPBrBEDPRFOeo3xRd6BPfgZsAkvAqH/vFje8lmdDlo7mr
26IZsHUn4y/T9+Ud+quIcQ4iE0snx6F9oQarFYU/AMxyVz+C10WhGV+NNdQB
4qF4feXHLCkJTZzqh45r+L3E/Hnki7tM83/gZwq30I2mB41ubUuesApnpohE
M2ghVh4+2oFpAz+Rt8MN8HkPaSEYsG5T86secYSCiIoblkkBVJhMM/Amr/ti
X8uD7fitxd4CvTgLPn1EYyXPtUe5J5mZtUCCTNLXaq4QNiWCD73NbfTDJSMN
dQm/CzhRrT1na5HRtT2CQgJIAVWp2Lctrp1DH9p4BenlrsGq75XYR9ViKom7
7I/UQ9QLd3R9bA2GSNOZ2TTDh8+MHU4xT8K5vxTkoN3SFYRzA5XVvSbUlFVr
g6etR8oJ39R/TZvfM+m1swxsSCf8SyXrxmFrEbr1PqfEGUD6jMFuRz5jNpWb
qaV+C9jIKmQJifPfk8+8bcO0FixWmCEYzrjxQtVEkwN5gM0uyOR4Yyg2spCJ
h2hc/KNXuf+sHixkUiC6WLLeo4zl+G49pYQMVgOupm8LdTUlqhh9m/EkTK3G
IMA0pDOjLTKSKr5PypyzqI/FGBoG94itKfBF1h4M+PqLkeQEk910rQKs57KO
3xkuZ2pdQUWVuw1pU9EYlznrS8hbFSzj9h1D1ZulTL52Liyoptfxp+6rbQFE
F9PaDkE03kB9FXMYu6fBxGna72tU0X0TZdqOe/TdM822oY++2xlvJrEmP7V9
pkrfSFQj5eMywGqblml+TOnMo6OFJCpb7IedG5pwShXy5k05aa1QcnEUpHUv
o+riJn4DgTI8NYglNV7o/J6WqCW5TjttUUcScv8Yba13yoiTUfLrn6JrFNWS
lxJw6HSB9nqgP4SF5UqEhGakQyDgv47YoNX8gDH8zBYe/d/p/4nwiv2wdeVW
sP6Q9C6YTIcbwrSjTILIXcDx1aCDVatiTjp371f01B+xJ+eAst2fetopgkgl
vzjqaWYQUr66g9epF71yESJEAQBgrg4yZrLyoklnydmBlvc8x4LUlbn3bRrb
LfLyhWuqbbu0WKYgizzSUlqpQqfOQFx3UhfByvyvys+NQGlDKfhvEkfkL7ZU
jKXyTVuaxXE+iDB77YBpXuo9zKgLLgwwu00tq6SOOop2riK4xkyVOpmkerwa
epHo8sAfWFfTq+z6Doxx/C6nlZXsj4eLArkFtUYnCdZjZ48SIkhxprRnxdQR
64W4ycbSg7goerJxmuoAxmmy0QHDAujZ8A0ZbnvZJ2vTqYksk14vVJFasHkK
t4aYYOhncdGSY5Ee4U4mxWStJdliBhthK+xMjRY27EgcpEG84eLeqeZ5IVe+
HzNIcocr0VOBfxFVqaQIf+Ar6qkYZuuv40eg3isb9M08MRJi5oQjrATcvXxU
b2QK92WETiK4O/7LztzTyP1gxzUV16ETtjoJUxvYVeem6iP3TzKp7rhFt4L/
mYzxPLx9OOAqzaq53TOrpR5T6drsmlXThGhZ4V9sowSUXKRjlN9TfFtVQSjA
xwH2msX1+HX8Gvvkbl2aCn7DmoY/xU2U17fglAmFOuU/8qglZASeXnqsTOXh
lR2U7rOr2XmpvoSDWPuYEaEywNCS97ryTgTA09Wt6i3RfiOwJ0FT9A8Fj8Vp
ww2d0+/nTpJTnP7ugmODC0GpevEN2hC62gIY9D4mDdh4MnTLLAoFvqi40fmC
z+tCjZ5ZgpDgubvvXV+eyeep6l7KIyLW9CG/i/3jBJZTGkx25YTv+hRV8nHa
Goirm5EKI8LF28//IBuDSyY2Pxz3mLo2gC8zt7hSUNjar1l6EvCAWwagUlvK
nKstdyYzLoPifBlhTlQCG1JNbdKSXGMl4hDzedG0e2xTjRu5ulYx2I7nEJxs
ckUOim2lSicHCuEuA953iCfUTTDl1/hcl6oF20L1lzGoXdpcprZnGj8mNbYA
f3tVXTEIeXcOaTWpIqwvJKZOElVMfwDWCUo+jBsvUDXvTgAuIzC3/kvT1aev
/djg/3rHfWj06LFL2m9epLqYZ6K1zfybHgDLk5sYNCjEVc2YDiyTtaDltMUX
3nyl1NWWSOcfEOMRoQmGTq9UZ1getY7Kh5AE8ECGpEslaZscZ1S4rxKoFoGb
bfWxazuTpk/pVvlQfgWeJgG2FVSSpLIZnLmkTo1lSUKCL4rgpolHxhKDSJ8Z
gv6tZnS769RG17eo4IFzJR6wV0B8Gd1DzBtrCImP6H9OwH4XkPQQRzOgfIiO
/mDUQ8BRIYvxxUIXWSGQ3lAQMJfiGvxqD9JTIWGQkuJ+mE7GsLYzlFIkPSKq
sH6pGvepHDg1k1wlNbRTDDX4JnjfTFJqD6MdvewAcDOr8F3COl5Pwo3vuke6
D8Jd5P3UGUXiWh7e94/Ku4BYa4pBpvp0ngOy1eO7VWLsl0Gptl2A0WKhfBvi
AiScxBIrAQjJuG84DfuAir9paZYlmurcosmtusMGaA6KG308dksQXRs+kfdy
7lYXtxv0I4EQW7mZWCXZlrbYybOmY/b9GQqgfaw/tMqSUYw/b4/bXIpHF0/M
WQwDEL5ZUe0RJ3u3+FXU1SgZqdl8THBuJkZQIHuXw0bXYPhLxzXLmVJ+Wcvl
e3kZ4iSfHVkLRAePTWOBCkNosywOhF+tgvZn0FD2GrpGAHdwMZSKRUpNYie3
owLDau3Ojt3VMxT8XJNHxNFIPrtmfYQvwFKpdpI9Ay3tUU22QA51TBke5itD
IuzHZHpf+PuV51zlTqvMY7np2ZDm0A7Qx/bHSXFCpDmUw48+hlaeEc82x1sy
1YFQVlkN49Gl6whtWf2MOI2r5vKys8nhh9xLsgMfFv0KAZSgaY6pf08t1Xus
HgABEIBMjBjvrY45bldeDLwCnSJeLFHCkeJCmnc+3OaZOzUMH1msW2aZp0GC
J+NbxR9ZjvtxNo+hc7Y212G6Da3jHZCFXJ63ImYf4BQ3K4iENr0GGlRR7yc3
fA+wJ3QF0eB53fw2p4naS5YQ0AFfOJUD9+wsacd/qOW4lfT0tMVVa2bKn5GU
EoIrvrwGbbujziTh1OuQzzSujNcnf4PIMgN/FrkQS6F4WVP7PHAYY/RuEYT0
efVinptYgE2CY1hngZlY4tXnZWyQIsHIpfIyP+3Q7cR1H4WfVMuCL6pSwTvv
E18a/ql9zYDNoYo+ZYdI5SK+hI5wY/V/0mxjRvrUOl+K7jp9OjaEiQl9o862
yBrWVZKWewoJVn8CmIkSbT6yTAek2DfQB8EH669hZGwfDhrSV4I59urIXU9M
6mW3t3I//p5wloCopknKcBxn6NdvMAtWkgj27ilD4syYDmmyIZVvieoe5l2Z
dnLHSOHoO3X8iT29MgNU6Go+KFP+KUb3G9YfcqCi4dd5LhuD8DjnxprCmFZL
4/i8vQakqkLWDsC+KcOAi62Tqvr2U8SO1g4+t1uZB/7dN0wYtt8oFduMYAUq
FzAf/hzCWzf7IS7kwi0dz4pPiVayL6K+XrIf7GVAB1tjWhKrVhlY2rO78l3Q
+SjA+7ba+ZuB04jeHpCH6j5R7FlJ7pB8Plhwu2nPka+cWU3JB6I7pg6JQ/VG
baA8/TUSdkamS5YaVFseHqNpKPiKb/cXBpfvCHk3npH64VS/qBiq25DPnYJZ
qF4X17hJhVBwdrTkQPWj/WwPFZrrmLCnm27JtNTvQJvrZ1mPL9f1x1530T0r
vQZSHtNXY2Rbm5uZp4EjaNCvb0hF0vECK0wvwXpAMOli0Z23nZ3dVE/KnxFg
EXZvIz4bh2b84Gy76valNe32c6LtSnv5/7kJUn+oKPr16DM4ypE0mxwirJN1
M9F+KfndXYANqzf3dHA5+Kos80YYsD+Cr35zPGKQJ3a2tcM2TJUU6nlqBfe3
M9hLZKQme1K9CBuaQZwPLdFqUDg86E7doIGqZMbZBBloYqlPLYlLRz5pfIur
99htWs7YSaZfdN85u6YIQOt1jo3eLarWTR8l/FLfCaEvQknrS8DXG4r8Zwb7
EKFOAk1fBX5HmyoqQPQyjm+XoGACvk7BAmJoSAfHxy4hNJI4hNmHq5ARalHE
xM3E/0Jm+ShL9WCbxXxKioFyisbEQr0gdq7RwpFXGnfmt2/xCHJBzJranvwW
1eH/cOjpYfk1dBZwgqxiPmqnL5PAkaEW5QclrEpEQJCpKg78kDXxcIZzsVz5
5c6Zb/2YUnrlopzDkmWQRsGrONphXvO8RIcm8Qc+3znOJnc28vjGKngwnbEr
RqYpINiKUxiIrL7IvppA1FGcmQrVKb16GCaTxFD1WvIwjohMdUERSrvACsnS
PI5mMF/7Z5S42zihSGAisek2M3bGncOh5OGgRMZaOeJ69mGDKb5L6B6n5yy3
NRIbp3v4HNYqEg1A0UTj+FwGBCPmawGgwTI6faL8iMmsWgoFsKbLa+TMxMD8
sCmuSD3JV8gjAfMYeupuVMr9QTKF89Tg+3A+e+BXu4DKf1y1lt8Vc5b5NM+d
GnQgfTD6fjZ7Yoa4YoOjPGuRFDdVmhaIQ9TEMDmLoGr1amYtklCuzHX1TB1T
v6ytdfllhOsqoRbWQbG1w5eY7vxVgO1Xx4eTa7Z2872+dby2hhWQQ22Eq75P
NwCkLkJimykKWdtmvmCi9/Lx4dc5Oicb7nsF2bVo61a+PloGxHx15h/t5OPG
++Zhpjzy6ht1mYQn9fjblqTF3oJPnKIBD7EI4vpmZYmDRII5ub55e/D2MrOA
uS3ONgnw6FNFBx63BzWcE9UunHifFBpXxRa6yRVaQ77HYM5rbxKrujU6ko2A
dQBZi8m9TVX/ia/qCIgHFYKuznzIYXKSO2xmQyBWCbgBY+R/yuJ+0WeZLrHZ
gc2xtTYS3kYgLmCL+VMkRq5br/q6Uhjtr0Txsz9Zf/TOz1t8iTgCRxJCMeuL
ga7D6Q+px6XOrWTNhnPlGdgTmu32s6qzyunoSWCXgborcVZSuBuQawt346K9
slgACr9RlD2IUputUxzBzWEZoKiFjLZVjRs+0Fqlo5wX4/Z5OurZgmRz0d2t
hZ9fGMLWk4MBYqiI+PPHQdYZUovG2lBMN25V5M7IrEEk1tmcaYHRv1IzzrH3
C3f8Z/R8nHKKCwEozrD2cR3o9feVjuV1MwhPh+tLLp4adB6Rd2+vS5tCSQCy
7YlaJLQbmFqy8L8978Jk4Kr/vHNZygIzRV6nmlNEBRDJT40AcKk5Ip6VcbBE
yJ0wooozRdGGcFrdxmqR/XGU2L6dcMNWUSaQ4BoJI04OkzLJvYrZBsH0mzEZ
D4Co9qAKcuS5UKX4U8pnROCPLkojLiJYv/e4JQQozGMg9cg23N38VKb9t+bZ
3atRw4E/bFmf0DIxF3Buz1wXQn2cb6Y2BVucf+uvtPUvI8mV83Sjtxh4jRSQ
ET8GFImcOOcje3gG9rmQVecqEGl50KZGqYMyccjRIKeZ/JofmMXYUgFIp9h5
7oLNLR/DMcX1CuC6Oyf82qEc0WzOz7GXi3Eir7Sb0rzbn/KA+i39JqrIIRT/
4lcDCRWV4KAePxofVqDPxgGMtcXIN9xX+zECz4bbfvKN8Z9e6D7K9iGcCFMo
LC9j+lxs0/5zcH/T1ttjolVu321kxjmobEaVnCyl6v0FYllgRlXLzRZJkoat
kiGp0fYqvJKuMP/mx3gcKYhHeyDzRclFsdmPzd+BMUrRzN4Jk1n/tERDv/w5
iPigbonS4HS10tOzOdfez8bZ3K8pyxrpMYbSa2/SfA3gcwEgQnl6GN8TUEBq
HF201cHkbvHyHA+5+l6VjWRmm7kYvzfajT1nQV8WlZnVr1+9h0LNMX/jank8
ymyrMlW5J1+80KvYhoAq/Avo/rJR4LIi8euNDM4t6OnpB1r7GdSADHvu79NU
v25owD1LMEHbBlwVOBdm9UicW1zJEoIoKBxKYpt21yNO1XgYBjrCemYxy0RE
o2TtpKLs8eeD6FnafgaYlCkHh59lTgiA26+Bqks9vLSVu15eV96ZoOYWEEU5
5y3c30mB5v+Hkk9p5jLErNLW36YZ3ySjIhi+SZ6S2C9n07YFZ0VdB1XQrUgb
quHlyKPkVkm5maLN5zKCKU6us2RsHjzbMSK6Jc4Dkd9QgijDvQQvs1A919vk
7mN2nmD7nw5h/65eenCCm8aPged+lKDbOB0NVAUZAT1++4VDSNrQOCxV+EMV
sprCpPKMTQA6sgf55UNbOMG6Fm0vvOzSZCIvCfvHDU0YziZvIf+RX7QUb+dW
2q6LMxXhhMw1O6ZhdAajQB1Q/539CkTwXO+Alph7NhwPu2ilQj6MGGTPxY+d
JIEQcELUVHbVNiVJHSh1LpcplGjmw6X7ZiYOlFIJf4conaFv65/rGQ2Hx5vn
FA/ZQcoplEJFmbvxsKQOwQlUgLVR5wKxnp1Y7HO78pVhZr0G+1NrqElgiDZI
5KgPlN6BombB1C8HXjMC7UndGjBi7AxF+gIis8Htg/86NHiC0zcyEw33t27l
6QoYrAOyOOzQRnYmdYIvazUkYyl3CMH3W+gIv8cwI+U2YfNA54vKX345r/cH
02bfo/buIYMZVBd5xFgFuaVCs8HO8GSfJGO/957slBAmongLjIoNyDoJ9Z8l
y3m/yrS/0uYyCdCMXXPi4Uycnx5MVecC+MTEbtjOns5RJQQWF90rzzxv+cg5
qIDsWx76TAZTYOqmZLSodCS2AWyCy+LAFJ2BJx4EKJ+ccCBT+fuGvzopzwyS
puNwrZpNJFI4AJ6G4K4QDvJGK3kr8orGPdJjjLRT+VEcFu4SHCgTV0NFAi2d
hWPQROfB7YS28ldC6kTi99kdJ/wXp5IbMW/Phm2b+E87/jJb8MlBPi3RJcBo
UpdcweYo3qAuDghc1OhYl00QCCABHbPWwz2aqK/cdsFJ61iON7iALab4OY/C
4R72ySLNjzKX7HkLjNB//o6lZrlcJoyMrHkvBBGzYDUnLOaWEI1NrcJpFU3z
cMHlXrguIuBnPipNYZOL1EX+v724l1fbiEVJJ55FAGxAUvbWGDgZHy8HPXRT
l4X/KYatgRU8tqLppvEFxBxAOcwI5S0UlJpJvbEPF5u8XIMqRSWCRzQf91+g
ubH77B/3RZWRDcioaCHcANtKHhaVuxr5p7HanRjLEObWPAenN4sY0bgO3IOK
gv6vgO/qfSd85X54wAlBsplCGmJBF+E53YAcSs8NRQMqhMu3KC4P6lRVZyAE
M24EnZeWNz5LOf0U2fWsH4T9Dhk80dO1/JGZUxAfHYg9WU+H3JFte6hJlhoJ
wVXKolJaORzKS+dkyvui8xTMlIvE8u8K2Rkgd6w+F3Dk9oLLpF2cF8F6xamF
UPTPs7KqxEm7dPDPmQHvDCc+gYnjJkuXBBBSzw5VdTTnYyLfdBSRYxf4+cpV
v2os9jCmjHiM217iCa1te6Oa02Cx7SsBz8x3bTndjau097+LZ3C3fF4AbL/f
5srmWi9atAH0LTx0R7iNnzT+8h3hpa8AQL5OPc2yAUeIFixkELUXk6aQr6ls
KtdMDc3g3AwdgAhFKDcG6qlL8VxsTPCRljnxXFm2D2f2lNguQxSHPcP7WugM
04g1TLmjxXnLZFIfnTOUEcuhakixHS+PqZCc5YCixR3/jm9UKZ9tHwmqiSMR
G8x6gyDc+5zwYjhSStNpgg2Lb/z8OeKMxUBcDJbd+k2Q/FTVYbRzHVcSmNHb
8x7I1prZNhsm9JNPXLdnDJNhi6eeVapEWsBMkBWpgLRZVPdzL/z5lDtXoWlq
K0K/imV3Sz90NwvNKIQXfrSakOAq+g3e7hunqkfhZlvr3+55kzQdUgWDKIjH
3twQ2GfZqxLFcyUxE/XQ3iR860kp77ERU+tjLm9lE1oN97GcCKGOpgP6B3OO
Dg2yTwmWIdUWJw5BUhRHx0bxuTUGVhbksE8pqAT6C9y9J3stQV2OaD7nRFO3
ovFoaw6VpiA1KIJqUkuxH9MsrtwU261a/rPhOeiQ8AHDarrCju6kbbRck7Zr
/bpfX+YhI7MVyLqcYLPizWG2TUij7kaDNO6o85ps2QyM3vCZaO88+9ash/an
9i+WJMgDBGfDXVKIBSXZv7zyliGwsYesdAgnLv/uy6nL9xEPh1GBZ9brJAvv
R0C1+fe4ROdyhYF7gPyLFf3/AENu1pjjr0fBf9odi4E/MqaMdhkILwQxVxWF
UwIGYX2TEtNryRudUlUm9OP/ZBd7aGkQa7RWZymQTl2gGmkYRSQVkhP3wTlj
0OMZK+etQHJZId2lICAicykaPDcDBV+jbS63UhdHH2QD1ud8TaIG/7YP/7P7
UrSUuDT5M0kiE2GlpYsPSjQYFPgGyO8fOrewTtOx6lyVLdL6Obz0kBuZ+ktZ
V9BIiFlvRHau/qCb/3+hbev/r7hclOts5YPTDRiopJiao38Td0FgDJJsj8zL
RbqEDYKjuuxjYY4tDREJHKnA/ldJDpwq0ohEA0EL4kMK9CP0Ybk7LeO0NVtD
IlbyT9ydWIAtiKyAsQ0KD/fyA4PYA+sBIsq5Unj4CjFf5eVRdEjmCXifVTy4
EggIbkRQ9IsssTkLPiCILbrHyvqykM2ixdcQ+vvTUINYxfifSxoewY9iNLO9
gaBCAkAr2n7OjP67BX5EuX6GszXpcSDqjSIHb6QYPV9N0RRgt7/Np5Putn52
qkdHTexEX/e4ph+IOAeDJRdWV5H/Ly5xUHh1wJqA2e+heVmy2UJZzFXMq9pa
FqDPCLyYeiZdCXublOquNNmBenlOuM6DWiwCW3qpnLia63Z29+0AynWfIGs4
f6ZD4v3o+RndQm9m/Jh4IJPqq+ziBWtbaS+mR6/81uYhKNGNoa0cWuayPs+Y
pfLW+ADizF8hpX19fYoLfvl5H7Ysa3q9dnuGG/tydyln0Cke1mOAwridBa00
T35VyQeEt0YcmMsQJf0FcbjKglbqLtnJigJeWsnIINKpAmVCcemo6QfBObJ6
/pqvFfLFfjgyv0qypZvIan0HhYmuFxC2i+9774kd7HKoCNeKBdEUFK8ZRU/e
drR/mOo2R3AS5Kh2EA/FeXlZ7nEhBfBlEJhO6I2z/FqFv4dkvzR/QvDh1We+
doJpkUfaKmtWk/v/tPXuURjbufWwLOytrv3JvNkMXS11xIaCbeo8XRJlJEkW
Hsm8gulCCM3ma1DywxZV2h0HcF9gOhhDJXz+lvCMEZZBk0W5F3nWxqNn9ZjX
TLnN3EIveKKmg38zSIo7AphYC6UTx7flHnmv4RLCEe7rLbqG9XzFDn4X64N3
u3PejIDpHeAZo5zj+LJ7eoUXGCurGYy04gXqeMdA2NA2dOP5VZObTn7Z4e3w
kbfuJiBle6FuwaQncvDHQ5vToEb1vxaSE+fVd+Pj8JdEFR08yVr/vbWC/r2n
FsvaCV8hZ3wi9E7NGxDfOIj+ort0LjWErK7ACZE5lEDXgI81lg4YeNxiBOgi
jDe/Fbcj+QgTjQQsUx83h+4XTlqCsjItYko6FMhBT4CqPH3FDWrTEroUG0Vh
07B/XZ5vNorXRaS1Aw+x8fF/KJlMINVYru5d/8RAsOn5+pSQUjgMjflT3Jpu
W3ptydOQKWJgOsBLLdmToeTkcVxwsaFnY5G7WO0CXDSVmmUEwNTtDBVOiZzu
WXNhRPpUcejM8fqUS/6SOypB8HwUD7THJ96ySnTMvUgvDytsAzmbBa9iV48Q
Z7TbuvxB7EbBQRpPXlbvLQcXlZrExirh2GMKKxJrOo6zpGGJPVphBG7+CCCE
1BT2xaFT6BgXlWcKV5Wvb0EFDmQjemn/D2y6SMW8QW9fQzCdm6RW4H8BjIMU
bOaA8pbNNQj429rhnP32qcf3h8i68OmvawlQjIE6DS82dHwH55u0IZGg0TT0
xHQRJi073acpiZhd50KAB2vTiWCs326Dtej+/hJfqja3gsUxf+aqqbsqvGDn
EFLtEZ143uBf7HGYQuyiE3Ywre2m6s9cAiFC/ziV+lAbZizErcVOf4gns9BE
t81+MyAKP02z0Zt7Pp/x0R5X937ZLmLSAQGLzvBQPjgG+w1ImVOnNUe7n89Z
AHZn6shRaDL1ZXXo2lJX5Hbxe1lFZY2zdRtIpYcz5ns3T0jDI7jCe9+7AaUZ
fei75W9qEgylk3bakhvHSYWjbmBqKKkC1rdI3hlm5VQ9GhQKEUH3pH+/ZpyS
bMMI3l9mnstWIFK6D+77KuQlJRKWT19mgWL9IlOEVUPcJGzjgAyCpiiVqj9J
awhUEkeslfs47TDQyJcs5zGTcRLKbWti8Sa6OXGwNzQboXWTRaY873p1amlQ
A8kuQE3nDFbnMdkWr5/J/k4YQhzHpHKX7ZwTu4rnLmSt2c09aDfDh5VK2Urk
/Nl8gy5ZriHHf1NDSO3QuWdAs9Aq0jVwLd+9WpoOIpJr+8g8DhRPYPGlfT+C
Tc7EIUAALh5Bm1abxRtB2rCVN+gorLgi9QjzB3iSi1nrx2vn8PAEvfd/zjFu
1MFC41le6q1HWZezJYsMagy4y1sxzNS7SC2Is3Y2r1znUEHlBBjFcgvhz8xb
2NfgNNzqiHXXmNB6EhrG/y1rflkBoX+CTAhOkXs0Sh898N/Ra2fRf219v/pm
fB4dHkgQepJhCZpcQcTwE7b4x1ARAJAki7ftJl1VPJb7JBAAPzbSml2GPJNS
E/xx6F2tUIBhnQOCmnnAksSIZ8tj5qVNJd9tit0C31/6yH2QJliyX0SejOd7
OBPmpm0hrDfQaKycVVP1+XG7vVKhGSuVqVRCV2+GqhT3N0/YkXfhEY3rPtPA
2Pwg9Ux1vhkfcptMAnkmJ2ZT1MPfBrRbv4LVsNPtcjUPOUh37HZTE3ngkwKv
uXt4rpwIw1Mb0MoZ7iZV5YZ8SWsCrvfT1nK6w41caZ+F1A9DjcFVOoaBV3dr
2IHY1kRvRD5oHiWfHGzdp6JcjfvbrOJAbgf0Ro7LdfgJ5SEgXUY9zX5RTTQb
VnWp/CLr9hm/xWG0gWWfS9NQYUheyq7nhOaNXzhWXwGVBcCl9rg/M2ZHKmVe
5UnZo7+cFy3SjbZ1a1iiDDJ15FPuSdCeM0KhoTSloES93j0tuTjcIi0ReST0
W0qx/iih+qnupXr4z83lNb9DhSs+LjDVY+mgRaBs5mqjnt4mrRuZ1jrysiVx
MAVXgxK8Hky/zgS4VjnpApThkccGrBvw1We3+tlya2r6apljmSX+rXMB2sOa
OpD3+g1Cr8QKaWJq6jviXY9Sr373XcgoO/nxagJT/EmQjz55rYiDpmGfwoqY
lz6CI/TWq45GtUz9ssjT7wGrWN6ZFak6Hnpv6BjQEde/A2GwwASuB7zNTx1X
k6DthPt71ivmxvuAAtaTBlmLJ9CfzTEdJ1xaINzPkt5Y+N15mOJGqpRhKpuW
XkHFkm/DS6hdKcZUjgXFAwNRkxXjGIAHXaONkd7u69pYCcSTfIyyvs6/Tr2d
EyvytaENcQLXj2b0KMwfpvutRr6+HfJ1G4fJJ3pJnK2PPozY7lQfV/Ll5h5o
wgd+jqbIAbMyQp00UFXnMI7snHVwrlFt27/pmvSpDovpSy3fc60JH/8RQk8x
RbPM0a5QZ6e7MZM32qEcUv15MOHzSywopRCjZKfRGI6ONoKi/Eqhi2znh55+
tZWkM3Sp5x/UJYEjsosNkluJ1yXvLLasygmLNIAMxj11Z+e624zqubmObyFh
gFyZiNlQygiKfzRuoSIow1LTiEGWMpmyfglsxLVsMrGXNZGx02mM+X4WEn02
B6ahiOKU48ba1paMIvN2iVLtrhv/2ppvQKxclK6J2Vh1x2fnC/Vm53fKotLY
1DeZ3dMgia2PK0/UUhw9XIH9X37ohBex3A5LCbRJbbenCBRgmaU+JuZP7ojE
vDx9Voh+2vid7IjQ2OJCT7Gg4cdk6hASJnvVC36dIokgGjWiCQ9WFF1MZx/Q
0sSCTUmozarKhsmeqIyCFiXd0nCyN1MVzgb3GWqrzOikshEgg67gLD8AR65q
mnJnPSekzEI5uN24szhPyo6Lurhjgdce83cs9bmayAQUnQn3gg7kcTGPjNyq
uSKLTy2Bf1gU5/q9nc3LNJELA/kSvgbFbtDvXAS2w8lfl2TvYWmX2FijAfZ8
qAuqwYOnta6zliNGTAy0Zy4hpzVmsIfuh/Rz+JuuOH6lc2tAToQCj213N5qL
KKz06YIubEV+Y3lPXec2Oaa6hnyDMaAKWb19AGD2uplpiNSpg4mBEP8em7YV
tk0B+sk8SlUFDvbvgP5ihjE18b8JVX6gXPWHmdBHqMoV1p4h3Tzq+emWTL7H
MB8XrjaNbjb6Bo4c8uLNU9yCZDcphV1iS4CJYef8XHJnwtgoPWkis8NJdNmz
b0ZGzmFSD6j1//+GG7QV6mZS0aIPVI5M6TqGX+l1Ug8XSv5ZE9yt/foEr1r9
5l15YnYft12ef6FFr6ljc213QLuf+45OKuzJ2Y5sBBwDP0bHEa3n9R5wIBcs
f6jAA7X/WxGaUwbxtfp+hjSbGvD5WA4MzPrxGFQHTAyuWJGDMqUmThFxCYyn
bPmNdGCgRc4wQRvJuqtIQ0j/71bATOLBRGPYhH7ErOa6/BjSZyL1GwjjbQTl
hQzEacymSgeqtIoRgsf9+4QAGPpFIVFAA/QxsezqT6m8UvvVn42PZGaRxdYA
fKTleLt98RA1zuJR4c7a/g6DgjD65ver3lENjka7VjOiPBlhamaSNy1gp/Z0
EQubHkaBf36TMdSmy35Gk3AfvjQWMpDaPJ56ypcrCZpzijC15LtvRdppY7x/
jgguiYZli4Jh1bz5yHpds4ydm3wIp+6Kuf81zqe5gLWkvgAsJX5e6d5A1ecP
NEzVeQQGVrAiTlRlJErZgc7NOk4MAI2rAAk2K+L1YkjIKBaVMrGYJ+7XKzjw
m8JC7iPYsFSxWlvgVE94IwPVdRa5yV2ES2xDSxGhxB9iX/ZxKPEzHqFeIZEr
+xYMJ9zmz+pSTyRGHkB7maiP8CkBkZYX/5y96ckUkZ8ewgCo+qMVwbgnWkZS
ryzh0JQ55EG0RhbpHXAqRoQ8mfXaW16Zlo9P03vs87Wp2wZfGvmcq033nLwj
1PcDvpANcsTOwuWWF4+lBxEW9JuHk34zdk3O2uEk2pu2ra9GztWpnUEHdTJw
HKrFaYHo9VMraQ7FFdt4QlMK/PVfUSwDRvxUDcl4OVopFEoGaBVG5HkH8J6H
FjMbC49uyK0VqhEU226tuzLb3CtfKQcvCbY27tcUb5yZNE5uUp7adNFt8ntf
5mQ2ePaQixscwfzHXQ1QntWCwDcc1wIfp1mxcNiUVsQjyCDq2P6riB7YZhkL
tnNN6ciQt6DwWdiuVKh05L0WkowBgo5XkxQs26rs1yOoQanTk0GvvaWA+Ps8
Qj4H10x284ip3BeAgvVsR1br6KQ/Ux9DLWHtyy1xoHmdsgtDmApCqxXUQXFq
8I3TCoMoW6+apArNhylTpXJaiDlgqoPinzI8u7JcqgQ67Nm4aYR79nsyIddn
8gZ2Lf/sbpPixE8KbbfNWVceWqJkCboaY6wOuIwYJM2+d+hY7C0jmLKNrI1T
W+9dTTa5LKrbM5uQxSgZ6J2gHYO0iNFNDJmeI2knL0DdqP9yFAASLnj6+n4I
7JgE9/pv4MhA91x+8JNoPK4D/a66UE4MCl8SL0PHM2oR+zmLzmlHEWWZ4+M3
1PM8JonBoeburqA8LaR5hDwDb3eIWBE3X02+JbHL5DB9XhX1zSUtRrG3ZZOn
i9l5i+111+iERYTi6c0tq7YQUrOUUSAlcS2JC6YUcWoCubFEFK3YEp291Twe
5yMW3pECOKjxu8plPInXjS+oiZ1tFCzeSn6LrMi/ImFGrNiuM/mFc9Pnf6vt
uIN3MMVwM2eH9QFWFNb/FVJVynU3DCiO3xJG04MdGsWgwVpgpv5+I/0qLvod
27YFqop2S06a6fKXAII//wXUmyQiZx0WSTkFFpHIjTizXtoXDrHcn55Nw5rW
MmkbJNQs+som6DDYy4JchLWKvfBb71gN/kLJvOJR8xDCgm7efpNyoYFrytT7
CL2Bf7N1DD+ZGWiClRS7kUs6JesIEYqu/8YyDakIuG0RAMzT9jQWg4SUPCgg
srIeg+2l0/j+xueaLB986w/3rYz9CJGGbShJmLkQjSSUfseSCxHz3LAydtM7
ZMJWxuKY5NZ4I43cvQXLARhWV0l3feAItNiS7S689PgIrwDZwVwdVHj4w+sd
niYBAWUlcYWE/V7eH7pVQ38aSivr/Y/g4QprJ5oDocC63EcUyjK1+2coaWk2
5YGB8q7pzlW6SDKmiHuPeYOrCA+arjYmW+iOw2W4EKNilsSwMZItHmurnNX7
F8hWIn7BMv+JTt2w2sFf0gn5RZfoF9/dbftiLfrQhlIsQnHsbIPpqh/AOi7u
0Qqs0I9e6sRWZX/sNljyeaodLvI9iStwvH0kGR0ovvX3UMLz3itZX6IRVCKQ
jfVZjIk6UFu7xJ0VO9mYLgV66jUxA8/laDP250rdTUMIjKdFzQV3iBtqzYaO
SBgxv1xslnKBIdwgxI8+cvPPViGhz4dhUig2LeMZF1DvJ1Eq3r47WAbx3jI1
y17eYUFd31HhNGrRWJksj/HOg/GTvYb10cOSexZuBGq7MglNtOV9c1QJVgdu
/iUDctjeHXuVSFvQsHOS+LfL7VfS169xEpBEsMWmyNjJtG1FVDwgbPHfZB25
2bCxhaqxSnj9P0lC2KeVKFfZ+2ecX7q5SQN8MMtJsjNNknFMxEnLCPP77wQJ
38fWEicHiqkF+T0UsbEbd6kOk3eOvp9YBIbMVRiw6597KFPLCWHCHOciqbJz
Apxgh+IaAeZSaAAEy3ctoHTDyp6Q++WV5Sf3guvPJeH3YeBkqY2TFr6ujHZc
/SqvaQKhX2HYrO7zG3vSJEuhCa97dt0QT3l6ys1cfwXPkoQU6c1diCKieKI3
xg1BVD/M6BLwnU5eK1JnMP/TK5gyPiEyaPPAQ7Wq5jRDMcBWgpIzCjSXGvzM
m4CPNUBEaGzOGVLFM8aQFCCSJtlFmAzd776HPbfVuMiTsqbD61rylFfvQw5k
IbDle/L4j6Lya5+lR9uWXsY5shrMI8NytC1Gv9dyZm8b0eM6wEiIBEZjJQr1
35i/J9TCnNOPCUocSDUZ5+q/Q5mmZiZXRXtiWxvhNaPUaQpFHPG6ECnzx6HQ
VPLqC32ybnOM0Z5ZR+jvYCMh1HAuqwrHAVuhMK4JLgX5EDoe43PoB4fY9gYQ
no7bUFCnPoEv7y9C8uTtc/cdkt9KCcFlDDEv/XxQ34ul+tYegcRv/J/S+xrn
ptLccnPVtY2TmzRyyANpKGZaqkGeCvC6X1MCT0i0cRGxH4Wvkc/DH+7baZLM
uU2k9tji0mEmXe/GhmoWtMxaMikIVHN4EjTcktXuRyyr/BEuaxbESJXk8fUn
p9qmoYv8DqEVAY34eONgQSP59353qW5eoI4bpMmnnIC0jVmYuLdl672PCMP4
5jCcQyU94TgiMCQodurwH+U8PqNB5FrBRJboqY6RQNKxoxuDMzfS8ROSwNIh
H9H1TERvivTwz7eJp1dhIjVcEFehBPBaqKXdIxnytu+rJwfIHgmNSczpWfvI
jf30D1Icmi0JK0Ujv1myopu9AxGd/Aq3HzG0HEgkK5cqhoFuKfZ8jNUakI7h
jSbE120aJjSTAeq2lJFZdDEG6BVF69zH0kJQD5i9b5c4ouZ0tFuFdvVJzx5g
uJgXWLiknpnYYkBRbCzVbTo5++S+qMZ3mJJzrv36pEyDhdsgjsQbdkr/1jqV
wjX7/JH1Idx6ThCDUmAGbHtnUjbXMVqjnj8CoPgnM9i7NXTwFm9WbYpXVarx
rKCDmtD8/RaSwBr68Qa1NCqr8aCZaYPxHyRuuoqsuit9TApYAMjy+BPIoLFJ
GOHQd8IbRz8jvjLgm+vie0Gy5zPw5FkEUMfc4+E5ZUtjkCO9X+bYLcSfI/z4
tE/aiKOLvA6wRTLGDqiX1xxYvyB43wNPmzr/55dlHDn2xFCgPNHrMbhhCOYo
UW26KbO+T+rcqXQSR4bqYxXixGbU0h1V+YvfWwuRCPsgfunqx7IXpNNKOipW
tii8klc0CFBRmyTrXFmxIblr+zzXSHGejKMNIJVugaCoZL8qKhnpVqXMiKwq
N1XSx7DOI2eYzeScsutVvF+t04NyCRQb8rZlrmReqQ5IPhfNWXY1f2p/TQJ4
vn0rhm4GrqklqzEOm43k4sGvNu4nlFFMrmOX76W17Tq7Zf1HZ0uvpxru+xOU
V9wvZ8CAnopJjdotMz2R8JL2ezjpLRZuOl1eL0LUpCs1dKwZHRVpgvEw5LYX
IIvTHQYMobV3zOBgup11VIyGxl+xi2Ct/aJ3QFQxghcwi2ZqPOUXHzEveHLc
NTPoH9Sqndk8SqHvau3d0/ZVqxDCzbc9BN9OpH6JGUouNrM3wvRwTRrURjfS
acBzGXrPx4cbiBfnLZkpDdLE+pwDcUf/G6Ab2BqKBsltqzjzvOHg5PauazTD
E0qBD//b7ajG7drEmjgVtCiKIcQLBVq8547T94zE8CcVibzXaIfmV+wd59py
eJvQGHo3t2m5oxctGtUXExqxG90TVNffT/DOmeAkOv05yz/e1mFBBGn+oP2b
3jZ54zvhFYDMWE2PIkaRxyYMR/DxGLI081BXZbihc8BY3o+p/00v76tr9ZZx
20n4IgWhqohhQqgmH8og7DjNsvbn3jXuHblQgyR8tlsW/TKU+ynmAxtbrMgT
qJ/UdBJoxYXdTRcE9/0zNQicFeUlQ4rgNDASkbv9Ifeju/DqmkR/c+Y6/QmN
jx6nwmQFu7oLksPe/FQ7Ch31M+tMuwUX1y+5orG3ewDa+G8hc/f4Slgwf0/b
z2zKqOlBvetBIpIEn5/jfFfg0NQEziMAOsAmjw+TT5bqeJFchBi1GILgq0Mx
FO0HdZj4jRP3A1br3YCpb3NjIjphs+i4GhQaj12/K0iBrpKIa8JlQlO49Xux
uZqkiF8JoSgUpNxZARsOD2tVsn4pvqeSt8Q18E7XavW9YjwWQOcjmehktmva
xQjAVlqwDwXJvZUsgIaKcQ2ZROBKsd3KlZXzM46wP6tM8Vn19Ybvjxz1CLLO
vnzv6TEahpLDULwyAr44yK5kmIUfbEQUCk32GdPkAx43V3A7MZ4jIFwrsBa2
HlBdF8o6dbeqq+0K3NycykH/wdxpaXR5GvnleCsdgtz+vjGUgR7EC86q7HGU
vMMwy76htTFtsrWAIvDZk3uf2/85cklwXCjtpELeI/n7ymGUbOOh1DL+hEO5
ckW7G4SjNS2eKMuac6DjXvjxImTgO5DvBunDKUSU95LwN/iaObngAwWQhU7m
0phIHUWakMxM/2AldwK7FVEmc62HuGyHiRNHTgF0phggkuT8cO05qS24zNNm
TiL+N0v9AuOLDv7hGfq9AzENZpnBGaa4FJvCCBBTsquPke++zsOiTCLviEOv
LroP2AmQubNQ818q88ACsINQ4ByaX53QEGzFmSdtson4wBwf6MxuPfz6xo8b
rFQOzZzLyG6uTB1G2vRZhoN7ZBwFJ2upZW/teB6Zhzs9G+uagL2S0g1scw6v
SYEzft6RuCrJ/A8pZ5kAbtwEHIzKbVn0tfLfOaXrvcR+IGtuPunvX9nHY/Or
zsoKiX4xnyg4UZxLBVPg9c+5om+4fjJ1yUpXZEDZcZdjIpkyayq8tTZAmdkj
YQ6/YuBXxMnjKy4RPYkZ2eWZ6Hjsqkx3I5q3T2DzvwpFoF1ntcrOigAsUXzc
jsWGqFk7FwGQ8MIF4hAxWIpOZqmums2k4OntVBl9vUw9ssu7YSQbUsCP8Rs6
OCwTZ/T729s1+FXVpiCL9n/9GhbfsEEhRtKgzf6/tnq3z6Kk73Zm298JXqJk
UpSpr7LYvd0GG7tYjdZZidbVe+gjXauIXfWxiF/OeIUOmBgohyKrvAnVoJex
8hOfvZCy8C8yQpqgXMDdPg8OjoxVMioU6coNIUAcE47sYkshB/L3gMdNF168
JBdwK7a9ZwHi9vjzAvYHVQrycEucxOZKuYLo8DExyp7fYvU5EqENmruz30pN
+SMTQNGMCyETkXnw7QerrBWqHIvx8+xaiIgWdrWrL8CU/YasbKwj7dCU/2lq
02n/81dvT6FiFVLr5S27tEItor+kcyef764y2kl59KXil383vHR0lfBExHlB
g9E6U9inGWMibm1cx+eoCew7YgiM5/10tzRXTGC4ncII7gkArYM/FZFN9f5+
TVb8qBKvVkfnzVUodQyda6zSitw6hRSafP02A7lPe2RWQYbbUinDPzgkyzFc
x1X1ns5QueZN0nvgVteBH/wzQhiXGi0uQbnL1TQKDYU+ia2p9gnCttuTBvzz
hNYf/E2ZVpKtkJtb7KBPgJRvqbfLg9Uu5Dspbc3P3OyvDjC+IrRAXwXxWUai
VdJkksJ5Mt9riqx/GMAxeTXZON0nJ7Tk6ZeMGZ48yLrT9Xc07XFzqj/x95ec
lsiFQhLQhX4NZCu/8/9AGi9u5xrO789GRmCnjNEwDdsPGyjHpJbIYSXoRYaK
auOddCPwN/iMr0KswzzjaRsHnSFNfllPRbfdvW0NwlTbRDfkwHp4nEAKAKU8
T3htg/B9eOaYzS4PgR8SCgBZsm9gEzo+5UKriBzuReodHPHX13U9vlU2dUde
BzpYNLpdivMukK35bYBmuIBA5FhVWXfK+GKizR+9nvrYubfkFCT2LU8VWTwC
S2+unziLeoL9vGNw/Y/Bw8mbyEaQvuemNw7/mLxMCU7Iy3cDbTKMTq7ZADt/
K9QzgKpD0M+YgK4Qg9ul3zx385Kkw/y6q+/23IInjpgHlEKViHQ4cuSUi6EO
S8HLhjEuGkxfDPcgexzHs/D322C5DYnnZxH6+6h/zGu4OeG5VtRSuijpzPK2
jeh6LQWqLRQ+jIlTFyUB3ODJsBdflypuWkw1zcLZY2mAqUts/2YbOXzJrDRG
Dpxxetj5PZ1ZsIRkOdjaiz/t+vat80wJJ8/9tXw+WGEfnVTqZM7h6bLXkuKu
WMMijlBPSVT0kRnPTtMdYW1FCkUPsygXblqlbSuWAymgxwQydEpl4c4t9mLV
CUnRdQiuRTg4YVj+p+AMSAPFrjJMr3H3/rO8vp0HirPu8hUbg7H86d9mOXTb
BcHBgFSch7vEN67dSLrb+LnQnXOHAlveWsQIkDoAdto1yJ/btPiQm3W6Wj+5
hqoqq+4FsppJtlNQNeRnhd6isDTm9G9AzKUH506zGhggPlgjvozDj4kZk2Qr
CnURi3DjmZPFvheXKtPzKLJ5msRcZgOKekA4obG/gmVyml2OCzJd1aACjR3m
kPTy4O1I+qbLRyRwz9LFvzLjkEicfFin2105+/MN+LXmkDJTCd+CPqnQlQtu
TTXDo56q54mcSZeDasduoE5s8hURonwSBN5E6KtGeguDLQq+uxEpaz6mlbzr
rsKQZvFHy8M3+fO6dKgj9+ZDNw1DQATtI8D00mk63eg9aNFaguuk1jrh+W7A
0ruwis9Y8eRX7wSVlzzJN+OHHGwyQHxSrwTK4E/euD2bCFqRtmqSrggbiltX
KBD8oGZzPby0C/zfBvuTjyiaOFf747AWWFEhE44scBditrnjn2/1HT8/fG35
HMrH5eNgW2IgXbtAAUW/8r0dTJu2dLTxzAMNylnJJAaKAiliE1wmWQuiCr8I
nDDhgrgFNopVXbtWbzvC8NbQmejaUXf58NTFkoPkf0jYyW0ZiUYZn4bYyK74
mij5//zu2JUp+ZZqDzRDTpWPofgBZ3BL8K7IQRlvK1B1IDLNLC+g6kdlbfnt
ZVk3X0NBTv5wJyOq1wwlfhfzsmAD5XyZz6xK6aaeMu6UXyRKSg7KIIZBay3L
K6yjq3A5Iwdv7LYCuQhSMtrvoMhqTv2/Pm49j09HABYVvOFKvgR2cdbllN8h
MF8vvUiKrEERmeyTS3nZgUola5quQ1kbZKG7F2/YJCMaSiDT0c7gg1BnRuVX
4wZ9Oir8h/GrXoc2fMR8xPsYcaGFLqmGcDar7zK10sXzUCGHd9yH8z+pe/2B
MmBhwXK2jVWkrtdTTmON5ee7T/MXrpUXs89IeUTyvH1c1njZtlcY4nGmHP3J
UXqKX6duaF/X7WwnER6sCsdBmp6gwQsELZ01I/tU+LUk/Pjd4PdLBbusXG6/
QkyNTMy52X/5Yolgyfy6KZ6z10s1L+VMvzIK8lRI5nz3vTOJTq9t6ifDASVB
tZvoz/IliY6bq5o7CdTnA4EHhpmjl5P8yYiusfxhfThdazTp8k0mEypouzO5
B+boTjSWJ69lw7rO/hHQFVhO4Qy/VFCiqZKX7wH9eyYmmOByHG/muRT3ScoF
ogmhKAM9udraZXO6RNe3ndWaWyRg+45pei9xlobwkSwJiJhg6+52ieKTfTXr
Vf5xjItQlwODaAa385EE6nx44G0OrDW1XzCmxPtqSxhVaM50umxNw5NiDnjI
ZQV7rbSqaWt7lIgcAPQ/QCb3Wq/fV0C9ee+YcY6qpSz5EJFaQ/R2rZsHopFI
/8PFYXeItZOZglAUj7ZRGeefL7FvuQXAoScqLMxE+lfRGDE8Tw0HMZh+hz0g
QyluwZSoYktWSa83mmzFJLp0luHSLF/9+vwkOuKwsJo724O5N3aMb8ADiGMj
37ApqyKLSWi53IgU5Gld6J1uBMmCSr9EkDQ9evCxMryhO2UVnbgQfj7v0q9H
LyHDKQD9yLpVOVvDnYyB8wkvMEivJy8Rk69/Xvc0QxL2STWnAXQWnrDYfbMW
aWhFOZd1TSF/V8gmgHXsxMWM9IV+J6EznMS9kHfNRK8bfYkKGE5OXAo+oW/O
5yO3PVbatpQIuxpncXrC1D9wH2oE72s2GCPh5BejoYKxEr7uwYjDFb4IxjNo
F6Q88pmx41JKdhgWuCWQOXjEMSQW6no6MPlKYoAq4zeZhRrmB5CHb9V4FcGV
wODG7QQtG8g+4fFx4B047dZpvNrUIw71LVIMr2hyqSxebFwhRaX4XQ1L7QA8
XhwMDTo0xUmZH3AFvr2lXaxEwOz4ROgJZ+455lwO/1Qu8bYt5qGCmftOtdaN
HGT5E6I4SfVE63vRSNO4NEc+TKiEk324qSfejTDd9jcaqIHC5+F29m8fsrzQ
Nm0RAdrJdBE62ybIPTytm4vmCsIh1aVhz3bRRSLTflslGrSV5xmJExsKtMuZ
D4W6NUWvAPx/aRenIh/BAy1p9HRCpNHjW7O3HUBD7QpaaX146Ue3WrU5+6db
WudOuOA1XO8Lj1X+y6sg1OQwNdlZgaVT2Z42drt/nWtw129MvFqA97x00vA3
aD2fCeXsR0clABWAd2fF2e8xwdT9VtDaNyZAcuayLG0On62X4TW5oGPkt5l1
7b6bhJ1hL3K91sMgl+eZG3FGg8wPYLVDU/vnoNH3NTwyCpoIqKKmstWtAC0R
0okyfIQ968G5/JduYtUc18zE2iHDLUbyLjisgImXqLtoFoq8Qj4BLJPYKhRB
iMph7jh9jHLa0ACyRzJsEbgIoTPqaUWIjsfntB594Y45RxKjQmyi7Xil8o/k
b0EV/jMff25SBGmtKhC2mZlTJGvYQTLpkVKYh8a1Fv0QU38JbwNzaSD9QS+d
WsuiS582gwwlrdr8nPAxvpriVt0sWfZG8p7KYtqwDmLiMr/ttJOJTEHQiOli
jDI9jGKkI1n0SZVJiaT3Cpa0fVj8uR3SbCdtpzo2WGj3BBQ7+dvvSxY4F+RX
xzR0sGJkGlggQM6N/pYw70nO8lpmqTTUUxmwJF6HcriqivZOeZvGXIS7K1HN
GnAuGHrFgep/g6Xi5yOIRjIxm9Dp04hTu3BK1DQpS0NCL5ntErLqQqj0QRVe
fTKm6t/lCbFVYnG+xYa8OxJc0JJKpuqEEjkeUPeqAn07kbgyyZstFHeJF2H/
Qd3LQGHvrswkkbA3GaVo8aILwd1HGSHAPiqblgKGO/OmIN2/RXUX8BjZ88Qn
fGbTs/yCFQhde/CpWHB6rkRkGE4tvPNsdjTEoCjuC8JjRSTUsKWeYw0waO5i
fGtMO6u4nuYwb75PBkVSYgrG8B1V6s1Sz+I7yoaSLuR/i6GDNoutZTowYEtC
IpuWSr2549sVXM/GPCT/rNIWyftIIoWeBkJ/05corapitQxirojHSuPoDPXG
Y87j+TPjXh62pQLy9IEbhQ9jOuj9tqnu+q6Xo1uB64J5pm2uJseWzS2l6mex
BuRK+0z8ubwOMCNOpjNfQtBGJNoJF3IDv5ZjGcsvIkVwmWlTn5mBmaiB/8mC
60NpsxtQrLqTztDwulz3of0G1lpkJXweQAtW2tK5it/+DrCC0oU/y4EJ9fMj
7ts+26xJZ9ILXQYA+LPRivwnOp3l7QKR1OWfZ8+l7AqelpQGPWG9tZspkp/8
hdloo3jx+Bd/E1OBBOcdtpMvSPHZOejl9QCXx0ZKE5L+UEwWDnJyOE7pLSPu
ohxUfx+bPnQgS7xaAMlcxMQ6U9ASs4Qixkw94zt2Sf+fEan6iLXxZqg6zd2Z
jZYB2nfxAC/c+bl1AY/au8FX8sVnOvZKHNZvKRah8TKhAJeFTETd0zKsq53R
YO9OP7oANcFC5avEsnHCxWIihCRFtN8D5TBh1skuU0nktPRwdpZkql/16jxW
JexpnDyt+wp93x9NTgPho6f71Kb9KAwSV6THmt8kHUHLlBvwsJVljABa1VSG
qaT70fFtzT/DOR34zJ0Z3WZcit2dt6zQNL7/ELdKUr4yhuZdvbbFHLjk7V7O
95OTbOgi1fHFP47i7boqZ+Pq+BBpRZm3aV11Lfe2orwN4jK6vxZ4sbn7rTwg
TlvzZ4mRnWxlG2f2lk/NMl6yrh7dF9QY8h/x7giljC1xfpJetRfu9FM0cjpx
22aHpNqLIR1McfC/kWIW3DCxGB8FcTx8gbwx32mPQU8Hnuzy8YoZkFljKBRJ
USwHyS8aIcTOCBYbJtMh3vywzsU+aEwxswq5HJHEfF5DxRO3B98Dw/e6JsdF
j63j4/3GWZ75plKbiTBiBUyqipf/+cT0aGQFaNAwiYIuNGI4Tc9DylIXkSuk
8dP6Iu6efz0rKbjnuJyLEhuvwN5xof91QtPOc4j2k9XznqG7XSJ8LoPGzBsK
UuXNuShdgjA/Jklivdo9S8AcAMTXBmnSnyCIXgPtD+iSYDe2g5R0A6LvK8Vs
F5qwG4kPrw9Ucv+GDSjPbdmU3MeeY+OrnTPO9iTVRuIHcpgbaYvMNaWX+unB
3/DkiCmOoOVAvxza/08QTr1Ag8f2Vl6cC2r29K3jYUXxko4pV6zqZGLaKQzo
Hfnu7P1jnHZ1E+ONS2pQyhIHb1ym2GD1LkR+yedSpAk+8O1uLqYiZbqJBdrS
o14GsSJTk7eDKMurJ57AbfD134AlT9OAV7sY3CHHF5IdXJGCHON+dO/KYoW9
ETaS+jc6bNM2NLTb8aofYnaPklfBHpjvd02nNkSBZN5AWcMwajD6RO/zfLGG
yu3bEa2uosO5vWS/3Z827sh+QAvWxPvPl2XCk4SO8OnPnKpY68UFCmPCDKoy
gXFdWMyHYxipCxJlswQK5isgETnfYQV2+ybzc40A7CRh9NOSRWSyC2SDmXho
RHGPXsTyGBU/7fXRX6diJodt7Vzk18JDO1tLsBjlHn4xMy7278mFggcySGh6
48P5LycoY2M24dfB/C5Kpk+hyhUKyX86qztburOSqjbryzZ5hGBVS83hl9jI
GT9SyCsqV1gklVbG837XlZvqg7HVIgC5Au3OtbYQdF1WW9+pkU0memBKUnu1
tIi5C0s6vwy2cyhRJK3O7N3F8zYiB36dHqruR6vMxZ/O5CRkyRq/3WN5J1Xa
eSDRs2UzwAVV4/bvXNj7ssAz2c3sPl7XKUEt7ie/ct9T+hEBX2ZG2qRuigHo
sQAgNx/VBPHEuSDIJdquis3nLPU7qeci7nFI/xb7/StLz2BHAwGFvLWWlAhk
zgDk35D4DShfeEPvh90S4Nc0pbmczl42M//K2yKTmFJRo14rFakinab//gRO
Exg/qlIb1sqx8OvOhpI/BOHJmHFmjrguvhPGAsJFgvXSQUESohG9Rw+sXBHT
c4hDb/L4Mogf9fQ3e3x1BNBEow65snaBgmRVuNtgZEyiSVKIkUdGek4kPBsp
RsvW1NBh+27nZIhiyHDDdRWVE0SshnRsPFXFj/eRj2hieyrDZsgctqzd3Q/x
PkyDC/b89SwogSJ66eMzv+S4zqcQ8mubfgxeqgH+hk1X6NX50mF2azDE/uUb
ryD77S9V+CFQnZvvEdsiCJsR2Opxrn7rFFOV1R14Tu2KJJcxjPgzIdHThOj3
inWiBzSuQlqQ/rgRxIsJnins2Ao1iej3WUeJWzqfThxKiV3pvTyP9FaDB2O1
DvrStPDTQVx2WEy0EPcWQsKmAIXcsKn1IibkDRXiIF4NACxisQ8JADiVKa4o
G9X5aa2Xzkml6XHCxE4Yo+SpBSm30+hAvtPjrrAr8oXbkTd9yJzOQSD+pmkA
/IpDgiLL8XPx0Iifs0Vjn97dL65r6mrGn1Z6xChKXXiqkbhoGFtkcRgEm71B
BcvHQPxUDFwSC8Ugu1vLJBeOJ2Q0WdtRTc8pUiAf5B7CY1PQ+9FEPt9XeSkE
MPKMuVs+iW45lbUF5826LnIhPa9cFkHeZXfIA0BEyhme1/QEEAA+fqcwQ7xC
yvUyQtb1gRIX7jMUfdr/B1KUaLpfJQNzPdfTzSBPwIZxec/py5qDTX7/MNlO
oevnCZtjp2NbTlgGrQJAZ74kMmZVneT8evsd8rTZXzaWF18Y0TrmTVVhYFnr
2th+epgVC7S1gT9X2YXVJFB3H+gkuZ3GpzpDSnAd2AF/r6XyoyGNeUgrBAug
puAvj46aT2AoN9nQFq2Q3OEEo1bd52/pBrSIoXucRb2RgY5GmJf2STsBeh/p
/qOJBn0NO9I8S5AYA1oICKpwKjWuzCOjUBqPlYfkAWjTHuAgHYN4A3fP61iT
qw0B0lJqjMQT5y9TbRXD33HaWSKXThcIqG+4A5o0m9z35/sYS3X/jV3D/HR1
7pOdxP4+Su7G0eNjRFZXqk/Pujhbp0r/cBefFa8MswdUf3qecL5MZ6bdRBxk
Fv3U0K16VKWyF3Qti3Lm+jFOuEQHSexVVrwaM++7xlMqZadtzNmV6DOeDPfy
1fjZiy0Y3V2GM8foDm/bd3NK9Cx9riAGJD7SP9a7nMbcGsNnTxZTo6q7pylf
XT81rXPpBbP0pB6J+HnlPiqTUiJ2uT4NhCeVzDCxWJQ26Z/Pp9HfI5LUPf0M
KTUuspXEHSVk79mOomzuuRwE3OmUNioX7AckLXTS96fJpGTdTE9IsdGe3ikY
uC2fDNd30IIyyDgLUshoXZcrx0A9RltMbtVNjlNP5tGFItlMYO5tW1PHkrIY
nHWeulMeZkeUsh1E1GSh042c0LwM0YJ6Ldj3TXW2J1GIZH5k61vKR0xdMIQh
Z/oPKOz7mBtrG9pbAVN6ZuIBMJu8O7+ZxB4k/kihILOzt+D2ft6ute6rVO3t
RMru/m/ArXDqUO7ALJJfrOhKhkEn335pu3iNbUQiNVTSkvNBzrWectR5ZAEi
NJZ54Cn7Skq0otDJGur/fqAF69xlWuvpjIUZLWfPHsznyFXQg66B+UsgJL+/
GGAMgU+RSokCiIguEbPbP6bBrvrL5PE6BHGpJBbtmzxae04V0WcPbN2We++1
gP5kK0/b3WbhDThzJraTlxbQ888ysuDCVk7vmopTa7yVgdVjeEZ0rWNHiGdx
9u7EKZygMhoC7VjwMWtiqhI6vR2bN6hCefykaOA4daeVxlmdn62FBfK01ebE
Es2v2Skv0cP83DD/nl9levOTGI9wOKfz/0DPWvq/RYcgpGSokNIZwQXXyKbg
3FXNMiUHMmvL0dUC0AEuSk4lrH37NjPqwzzewWmcBv1QNSHNhgAxYj2F0M2E
IFTSGhVCdfKqxpzdyPEbGGh5c9Ib7LQzcmABJEXJ6PdeCAnR91UcAg0iqMYe
BkXPqnR1NO+hHvafx4yB/rg0MnvaOofWUebFwKWePWcP4eUpl7ofs/5JNt8H
STOQJtLu6ooVwz9mpikf2DxCTG3MXD8fzDcVnhTbq4WD6l0715iPV0RMZwfb
jgva5tA09YCCVMkM4xc/zCOyWXleuQBMhOWOPSCYBIFhaI8jY0Vx5xzDZNEE
XBuvkpc+2bhoL+/LW1qoILWdlgzazG3V8bE8NbYETI5aKa7aLjy9xr6/r9V1
9Q/T0GGMZKsZFbIKhXJpfRgmPE9Q92pixqstBe12dvICWtuSRttsHUgdhzXu
UrmWs4D51d2eBoJwbD3A6oMT9saGM4ZzudC+3dI1fyyMaBGNZJH6/wNhhtAE
Sv4mgTqsa4LaZ++LoPC9JZSe57qK+3Lap5j0iNRzdv7/S3XvV/BjJQiwzPCY
ZMK2KlGI2JLAsBhgAtDJ7B8qdXPIStXCd0X9bxgZ3ms9kvGwFBRVgVdWDiR7
hreXlpyJpNt+nHAw0Jwrt8Pkgvpi352rtd8+BgRapMQes4czyzgI+qBFE5/g
bqM3lbw760GXSzWA7LQ8Hs1iXQsa647Uqd/SQi2ogwuE9Cs+13CAs01P/DDd
r4U7oSBD/RIM+P1PVIZ2g6E+y67MCvfriGbj8V7u6SS8FWBlwV3Hq5hsfX1q
/yjBXbaNekOUvm6Cz8JakdzB1kAKlkt+Jmvo1ZYGLV5vMtVG1Jrzh93QegEn
JTZstxHtyO0vwLVptsXhf3kRW/c3FCF72YM9ona3hTgoGKK928nAUpSAL3lH
fnJ+1CCUjNxWao577GJlsq91ReVZYXBQRSLKkwUmiSR2Ma2u1UJxIrlv/Qso
tKiolNF7E2Kh3nHCEEQgM7klwMBxXFeVJlUws+/g7+mx6sSPj+RQD5UDwlbE
S0x0sgi2hI6KrZthdV6EcR0qdlxEFX2YEVxhw5mjXIqp4xB23e00fYw/Efgs
jYhURyzL0z6IGtwHIrH8EjmEDyIjAhoZ7MoKB3b9L595ZVMVzs+J2qOyTUFl
AXnV12cub0M5F1wYguyqRmTDyQIFj1qryOF482GBSwULcjxQc8gwgT5Dh9DZ
xaL9ToGANgKFfrb0lhGs+0opOtmrEEkDgTuYXxikF/+XswN9xBoleAabyhV0
uolmfXM56zLZtqMXDz7KYy7Pu6idKHloOkGiWdIPkCaNpgyQRraBu1GDAj9i
/5I7zqLVcbGQhyrcJjmbnemyiZFQoLd++vvoRoTzoARTIFHxOMsTUNgEM6tJ
wn/Wr0q+Gyrp09A9ihQRlHKXf1OWibMRS830t0ohcTX8IpSI1PRwNgHVKd0C
E/bmu9zsqEGVsjPbex1+wA8A35m2ASB4b7ERA2zL68NNENQByfHKYtfdX9pG
LZFOpjCHXAp/aqVgoh4PcCQtBPOlNBevxFWkaZ1V6oadsl5G+dbwyR+cQcaU
dQJxrgS6MXn90e36Fs3mqwmKMPCVrRUdr9DQSDRo7bCQPOPoOTF2zzOXaa85
7KjHY+QbayejaTNbX21t0kcbGFgbHr6bSMDeAjdMMIcQ/qVIKw9Y72umicVK
bYUi5P6tpWKTSyAptNLA4XCE3KQJjK5VZ9sdWVYXq6rcGaw7GNW7ofWZ3rqB
TJ0D6iDgtrzsd/AhbIirhsGkvCKf+NalDc3dvbxFd04CAv77OcnY/GaibnBR
3MzAtBldjcN33ir4oso/O8vSFCnl9W9KNeK3DH6cViWpHHt3H0isyyJQWE66
Gthhua6kqkWWOegwU6VPpjzeaYMEya76x26nVDtAqN7n6H87kmJkSY1hcqq3
Zh7lVY94GPrEP9Nu3nHbDxWRikL23zhFwaR+Rp2Xg/N2bJGX8l9cLWs8CPTR
vve8zbtos45GFSpmAOLTwjlpeK5aF8aW35h4QLju7J79z5NZ6yNGzF9Sq+V8
7oSqyN0aZYpomwqAipFrlYUqamHnVITQua8dF5YP6mBktYluMRuN4KCzKhJG
5DJJELaMrxuaZ+bpobGqUd5KUNxuMueeHVnLOqC7DwebUzR2mZYZvUVPONU1
C1GlQLqm3/m0puJoW+wMn2nzgESu/UojlT8jJ1+jDIhfcqNHq9mlM3Ni6+OO
EUxJ6kQScVGgla3C5mpiCSLSHsxWzjWjWRUTZbXB56vHVS1lywmuqS7DUCSh
43XUOXVtixPMzwKnehzeFYodxd+U+Yt4CEtZ12Brps0pm1Swz4bVPhC8GasJ
vb3p5r7X0pjk0GGQgYkaEr5tX7w73tvh0EP31aTvy9KXSYxk/iQ5B/vHso0t
/SuWtysYWGM4CuPrn8Wuvpe2x0blwN+Py0Sft8WOJ9/FpTmqPg3uYyIrvs7u
XjIkQukNB1CRsBdt0z35+GwxRwS9nLnCxV7O8oYkqoMUOfOnJMOru0/q6B87
WTValOuzlrda9AnZJkDeQS+bmJCUnJaauhSGR5pZ35dw9yhjcQGTx9LPl9Ki
JDEXFQnzLaHTy9kDPdjW3woXGD34EmSMuXYaSspt9jylUtipO2OLnWp1Viuy
4blIFMgIgbiH0+6mqkApihaxx1cnBIl2to1UqhfJcX5whRdyCt3FIwc+A7NG
D9OZbAmsdeP0lJY4w47Dub0+7EQUzIZdp3AkBj+MqNP65fgu6e3PQtc6muJG
GRsooD3tcUNhYxAIacW0wjZTjMZYrkwZBrEZ4JMwz8GiuSHsC/mtFeBvxQNd
/+lRJ6ZXsligecOU0KVnHN7sDnCoQb1M9XlHWy7pFrR3+GPViXK0IrjpMD1d
zQgqMKDDgxbJ9NMnFr3wCCDnnelpjUIXyPnETYnNl9rCituS++aecZBdAPyK
EjxGLNdFTuXpwtZW64BUW1fXsd3MNagBBQEZ7aTRwgS53Y0nmPBnrRYwuolx
TEsH0IM3vev1XSyD8j/6XE3nG9iVGEpmTaGB2oiX04VrG17SXRY/LoODmQR6
UrkfGA3/UeKyEAekh8hOeQNRuFBJ1v1QDhjKkzd2DEZu1Sj4JXLHjN8pE2Gw
WZM0kW6NfTDcKzUq+foxh90XxSFwsv1/5ALo+skBszJFZleIBJn0TeWvIqwU
DBf763pQCI/fjH0xl1e19yL8GJpyqrqudPqCqAWAMJkPBrBggd0HMIjWfTIJ
PFtKmIQubvgbw0TzvB0cvnj212sK3kgSJmdd090eCdw2lEL45Qeu6KFt7UGu
87E0EpbW0G1hN1Ts1Y6zH8Q784/nFDqb6KpEw2v/IFTw2025a+i2kK6exM5h
jEqyuKap8C0eBRMqaSFHonz1uqFVmkoji75PO1DUUEoZgSDvNbYOp+qcYnNX
TsXPCxd3GiDC5sGS4sUM/Rec3VOLZtx/8oPMUoXxh5MHsX/lrqJvcsJckBjr
xpqZqhdiNfKpznACMkkEGMeZ5BwmFH2fq0/icDwKQoOZz/3ed0DH75efsONd
AboZPZokKrzShheYlO14en0aKOWU0SLvCP+uma5olyasA8j3EEHs/HHArySX
TGm+8sNmxZwZrRTc0//AY4TnlLd+EvXGqIKnLpwd/WmlQPSLoF+ZdIJUZsyE
jjCzhSCBD6RRIxOzY83T3+8ZWeDNxc/4o31uRy1GOF7/D2u+Deva7Ib3I1TV
LodM5Y5y3DMjxWt3av+aNscSvkMtkEc71ycDcuyzczdaXq6G8UOXbma3S2+p
nNU4x6kPAwwA/DzCwhWqPuYNmRh0ZP7xRB7XnKz5nkG2y804rqGsapYA5h29
Gvb+0x7go/indq6dviWomiBuFxxiohDCXccsoOe9CH2dj3dI3QZzCnBbYVfp
A6/V5GHA4TGcNPNg37p4Eb5UqdonK1hC+vZkhG/l09yJgUG/87T7RNfNGk/M
IQR5CqlmjoPAcmWbInaxLLmZV01HoSg1dmLP27uPyaXCtiIP1nc9RIfhjeDt
3mo662fyADBSl5Qpsf5VjYVAn6IZ60H8tEzaUyuLZvPGj6qgFpFPrInzRvvK
/K13Fdx6RVsFI6r5O3Oox2TOL1uulHBUo0h/3L/OSzkknPdYX6LY/f/GslG0
R1cHeUlYU2/IoBczfCCCugGpxnC+BRihP4CExs7uW9nGRGW3k1xUNCmTeIAi
XDa9Vqw67X4GWIriNhcV+NSp69CP/dB4H1AyOME2pSNk+ZOqIqjkrDSR9hqp
I7IEbw/XPIciw4OsY6ZOEFZ2GjF0f6OLsGGppCWISrWvggJSeFcccmxf7nyn
MszGU70rgO203MWbHEVDQPuSeXOgM4W0lZN7w+2YCrLEo66+aj+kkvJMf/Ag
8l6TgMSIl3k+S2EdF/ovl0OZLa4QTwQak/Bvm3Oy0LdpsHxvSuT5VCLcUBQg
dfw5ywe+cjwy2BklW++8fiUPukz+GhK/g2F4XyqsXaXccCUjbvxc0bkCkvhh
TtgwwikA4Xr4Lm6Hy2688Yj1qYRjSTalTDolqZgLJxtxI/SJD3eqRq/qi2E+
rlanFj5fhONlejbXBSMWI2NwJMxudArGC+NEwuEUwg2yfF//lEHM452NlDSP
cVpKUeHa9oKWafhOYm+fKbkmerXG+CHa8KpLJvk4sOP3A+b94jHrIJiMaCKt
oEzOI3h9YafNHcTI8Ir5agtCGfbtPr8drjjsiu6X40bL3AG9AZan3rushp56
ExR72a0WGwGFpdQucy+L8pMNYQz4D3rqQ8Ui5n4CkmKfWEm7rQm2P45OsOkQ
m7nFWXbBxqHgmIjEm131XWW+KDGoXRHplb9UCF5PPrpJM2exSnyK5sLikmsl
8QdbnO7wkxgcKx9W8epClO9RisIswtJaQFCFBePv4n6ZYfVaneB/F6cyCKWE
ghg0EVgbWQ6ugnQ8B4da0tPz/hSjzN2JB5grSW5iLAC1Vgj0zPlzVWOMud9K
iNsDyBGVa97oojEkQ0Y7WSOtWOt2YpaWOnk7IFzfv9Wxz9kP6sZHKM77WYJN
umUOllQJfwVx7JGtilV22wbReIXxTtVY/LKc2pBw8uin3dqjsKh5ZP+tqSDy
bsytKa+IborZZkzGJUcNrrOGuxnIh90pDTvncgpUHwABEhHhP1hUnA8uDgtp
ytSldgefIElx/dPsCQV5oycgah6xd49vS5WplfEM2Q4q2xLjOGl7FOBk5oh+
Tftnh9eyFKrsJ4JVPNqL0ZW4Hq9iTd37IoUbqKCCjAHrLbkkkH2vu0BrtVyi
KLNHoPe/wUOD4VwFnOFa03QvzQzhjWF/RbeXdt0/jNYv/nYDeizz21ZFPof0
0u+J2gvwxWKzQgsa10etZpkfXa2VOMELE4hoiKpJCcjkG2nNAnqyfuAI/4Yr
g/U4ZFqwr7U2am0tHEEYwCFoZhU+zTgL3YFX39+bxyupayLtc5+dnGmjK0I3
dZvzf7VqcnxeqVZ64MwfCiZqeiqsAtgRsK9RFkWlgw1kf2gfXp8w5KEYmY9I
xAvpmE/qewGncrTdZHsoJq8wGuFEfDORjlNx4vsAxRt8OSJfM5X8+wtk0DKl
3mEIHEo7tvw1H19YWq5u3MP/fTBrAXn+zcrd2yE/bibf+zFI15+bG9OYdjbU
Xrnl9UOtUIXjv90QQTTl5Pfjlf7NCdFme1RXysKOj1ho/1Nu6NJgxaDEkhc6
hbrV8pnMNFtPQ1dnRnV6jfMFjuTAJuOa8uVMGC5APGvWLmtHvmq2ya0XjrPA
r6AqOFiBIuHml2TLFibr2c0MWT8msL0Ex5EH+m11b+VrXpGbpoUx9o+gMwnS
lNE7gPsCvLq+yhJpzGiOohMmbcyTDITtSXmZI3+9rBJq6OCEjw+3/nxROU1X
dB+97h0X95nEm0B4vBUkomC7DS/HcxYZGVBDCoG9I9gTU+IKYmy6U5Gs+NUo
vPi1DxZwgTMC1SzdJGcQDjjWIZ2a4HuenSRqRVK0yLIVdEgNaSYxmhK/TeOW
oesVB2ySmCSaTA2X2w2T+wXklzivf6/+yDGLbkT+WtD68qTB2VNPvLKe4XEr
2+4VZZTEjrE0EJGHo4sbEgt3NfIGfPpogEr8YVSh9LGYwVtvEEkcAbM3EkHX
dkkWRCqSnY7wrpY09erFn2Op3UYYtvTDljhUucAqvBQ4WEdb94k1aUvBfG3p
e08e5XmVt62HqaDUQB9T6/48fAHq7lZyoyg3TkWc8jOjSkTpc+04FpV9HF8p
gTDZbx3RVlfFkApnQMAA0jz49Kf5RhACfyCBtBGAO7UFpCXS26U++WRJR5du
lJu+y80mmwE5ezUg/veLEYqu0nbGGYJtbRyC4REFbpLgn1pZcHQG/AgtE4oX
1WQvt918n8RX8BkVzmHBsTtn6l8Ptr6Q3Fpd/ufajjN9R+7iti7nUnfnjEqY
AFpdL6nZswSazEFvA8+fk7QZTId5KXVSwqfMCdojyf5w2+fl+TCDYfV6S39M
zHglIr0R6A6M6kX47El3ajx6ku/PmyYjph4nGdvuZDJfA15DE4F3IutT9//b
k9Tb+EXRAcBfCpVRA+tQNABOHY+llqlY9YILr1GqJ3Rs0y5NTVp+HQ54Aoe+
pUtezW7TpCajA5oQcZVVJFls9BAq4REvEnZQNLyrhGrdJsZuTlkOGuge8etx
Qg3Ym/fXVUHDYqRiKJeJ8ldLEISFds8GYeBRq3gv1EUs3lKqZFxXeuQIBzpA
Wq7prcp8+W4U4SdATarNMpgckgFwpSkkyVNcsmAlbM/TX426ujozWV6CgVWs
lFIHfHpUhqgNP49/YN5SPjacK31JbgjbGAvSGrBVK8DGtHUhMOvgNxnU4NkG
Wms26nkUiduq/5Pjjil558308xFsgOZWLlUsYOLIWrxW0oq29eHwIgb2iC/t
J/Xa4W7fUCxCoOof/CoRLGokOHgdhkDqS+ZSc/fSK69oxFTI82zybVyDDHxg
/lL1RFeo2EbJP/s06lc6Ckvk23j4o5YA9fDEkPWxYMJXWIMVnj00AA8+U8aJ
0oxkfyEFWauDMH36bUtUgWE0rbp/qweTVx3kZxm5arud+9QquSEdEMEWfA1V
4Emmqv0Ya0PK7Up8kdtUErDcxK65eTN08U2Yy1Nem2Efce0f3P6aOE2C2Ffu
HVZoBC4Xgk06MhLNyE42DVgJe8qcP/1GTRnuypKrt7Vv3VhpCDExkC20i104
egwvI2d64xwYaWXPVe741D8uu9n3cpqoHeoqjXbWe0X9GuxJhJauQdxlfaQR
h/xb+scQbb5tEaRHAqjh333HeRZd9XtSuOumna7uvZ8phajwvdb59MjP8AWT
QbNv6n7HahCyjVFrOn0vVfRcOyTrVpIWPP+QE7iW7Pk+G9R/dO43GSTjB8wH
v/6YnCsGHej2FQzmwD2K3d1Jx1hq4SHCDnuF5pZ5L+sYvkDJ4gsFIbGlHOk6
WB17A45iKInaUK1hw1+JDACEO62NcBxYhwBWqtFoQk25uxy3DT1SjZ04vFuF
Oj4qwgTW4+zbi8wlsLf9AZqpfv7wLi/m2297cwXZK5FXl6SAqy3arno9KqzY
H07SShSTD5EcK5Lke29g0ZDczVcqjBnMzOBdwev0Ogl4ky0kPOsnWBmQVTZg
jyQvFdhpqlka+nbIPWccGQqkKEgjdJ6NVEhQ7pCJib+KVvydHMKHp5Gm5Xgs
fynIS0L0bD6YyhlflkEuT1SAtc5heTJx63V/RYw9Kvf2cQPCmI3GiAnoGv7O
gRoLfxej0YE9vZkUO3zz7SB30Gk6vS2a0hfi8sd1aYPR8wpGou/zf6LlGoy/
q3saT8LI0j+36Hve+EZoFpdXdZJ1bIY/bvwV7De16J5cD5CBYh+Ll3qBKClG
hEcxMcT8O/Tr+yFerN7zSnOeEvbVlIX4A6yjU630eXnfmA+v9nMmV54H/WVC
b20tHT8WJrqfrkqzdQ6IwOPx+tNh4or22Ft2Qft+pxWT3vX1rBW0p3X4O95q
M2YCwRI1ulm61UXjzkhOakYvF9orabdKJCvuyz//QtH+bbvUvN1D0YpFZJ15
OCRqxtMlhWOl3CTCy2tdcYp9t+4JeDtNiivLQ+fN6YyKCnyZxChl/S/Q58A2
Km2AUdkuEsrKNcJIy2eQystwbx3daswNqlkTYK/Sq9yc70it5QDY5vy6bV7H
P5F1ZJVh+z4sZxkp5DEAwBLnYeEkPcxiywh9oVwbq91TGax0X9C9utMrCbg7
3UnWJ8jgwtuLV6tCQAVxqnLITTZsG9cg9hP1y/1O+m4U2bAuniWgOqCexPMv
hzTBWCnym3s1DYmECPzugj8QZ7r+SYufTStKBBGapYhoywg/Bv2zqPOakddI
AkG5KIVxSoAoi67Xaz6ZJRW/2unhHytyEAjIGnMUu0HumWe9bqBBsi9gvmNp
/dxkRpCnzaCMAqQ6ZW11Y+oap6holiKA8Ly0z8WCF1EMp4aPIRGxZnEFxEUr
i/NgS5WuydWaPQgimnHnnleVskoJQNaetzFKHIUzcEyQ89KwmcCUJ0T3S9+k
qyGI0EldFGyNBXfWivNgWoj3jg6a6Un4sjNXYI+0WQT8GU9OkiUTh4g6Sc0l
juk9jx1S3bQi52W5iRIdQ4oEJfxcaf1j4z0QrvLhIP0/fiOLkXmSMoBDVCIN
qTO22RaTE0lBl7JBWZFpgYSh7i/tPhEBZIgYnmwsyWkdRwRjp5NaxBIHR0N6
lapCZ2Q/4Jrd13YcuUewNHcMMxHu6YGT2MTYbAS+AtUDfcXWkENXMhjsSFBo
cBLcT/vg0VU231NEfUqhBpRrflj7oe5iwstofuBK4qW4ws54RGuFemJD4k5+
FSMtSMbMWypF4MT2ubFIOgrJZhkGDGIxr+XS/tAg01f2Gf6jGziIUT+lex0e
6ULZS/HzyiTk0WpE43g5uxnjSRATucaKo49fnJkfmes06Jfj/3xr0ZzDDi6O
WLfRg6uhZealjTPkenTo/OMwtAO4Te2OvGThtVt9gR5MW4O6QSTQKk6QoqEs
8YYsPS6h5YWz3m1jWwoRtmH8CVH49xHSHzQow0jjdEPz5ahfqVPm/xdd2OaZ
qrr0+iseUUJhIZNvC8tof89KBiwKECWvQ5xmnUyxVhxJS58gaU0jThyJe6Dg
1JghfvBsroSFC/mjjBB8/s6fJaMRGkZWIVcq2vOq+pizl7GhAem7reQ3KCuR
TGCeJHj78+Nz4pmdIsxi+p1A4zqJzY6bJi2im8xgGmYQaZLwKNh043Ybq4qb
P6qmprRYy1pPfuwI6K52qcSRtCc8KgLfzrSJqVlBlqfXJhF24/1TEsv6gxLW
FcB4r8pS1hxb6kyOTdu3u/xORCtGxqKsr0+oeaogu6I8Twa9yDgFxKfOA4oi
OeLoSCbFyp8c4ibR6hMxPOOwNd0GxgSaYRI87TKsQpEFF8OawQU8YCF0vPFx
RSCkfkdMkfo6XnrUieOEnxRe+zrU3ZqKA9u+CZMLRJqy9xpg+OqKSI0mJPNT
gTfj3+1nyM1SKzWX1jnAqJ9mZw7OMhJn+sQ+6a/jYn6zfnGqf7Gq9hZ2UflM
4TnGySwAHFURNwf0StIv3OQqfkM9TyCTpPXJj3vtoLAaxS8Os9HJGDOwX+Sj
XVOT7G79E2g0NdFgJV4SRGEEFe16/s0rb5B4VvkdADMcSCnEnGcTfafR6ucT
FniX5bhdS0VBNzZQxxcZWlU4HTybMxBZcNvd5WTwNmQQRoTBtJpMWpHZxYZ/
YtoGB4AKBBO/WRQxmeI0y9m8O9Ra7cNr2vk99QF5mvclYcudQ3kSDb4OTIwW
2kuYHVnGiptRAaW6Wm8EMG6u35Mx/HXTBn1HyFcOdSizoOXryaCvrqEUTHqh
mfyVe+3lDeLbM2SFkqYKjLpNfUdSpj3CaAOzrLWgalMwdhE6w/0GxX5mmqIA
PES+ZHyb76bodPQ2RHQXmiaiOEbKTObJ450DcP2Iv7SfevIMywf7RkOP5X4z
9SKIHwuPqb61ul7byXGLBRrKA2WkzxR1LvHYjlVw3qKrKxD74vfq+DoE/uC9
Xi7w/cN5xRv1uHGJfqLPs58N6lUuhjHb8Ij/9IOVeudfFrWtsuk4JNXVCxRU
4vYAvM6c5ggL6gZ34svOsTf3abKbsafJvZP8XpGZXGjRKwdnWYJQqS9hW0D3
B0AFqWWECExjPnlAq+qbH0iOF7/exffVE/tgxHndAVNYoPaZMZcGfZQYWk8i
VdjBUmTzMlJP6fA+AJnohHEwp9k6l0gE5r2LypraracjwT5fMnOmNMAZcsPj
t6/NxoteeIlNEcyEkS7FZuGpM6zDSey3E0Kda//C0gk07IeSf2m26YW0wzwd
Cp6Jvut8RvPQQ7QBmaKlUbxlva3I/fuXkGmtaA9MZHFWVpNZvh6ZR8f3TFjm
bcb0SL80ElvJ9u632LPEILsUUaWySicl3oCoLt90vhLRu4839+xXXJ2qnfCf
1AEuIWbFXKXT/RG/X0Jsy6285BqYewrEJRjtnR4083Xmgwh/tCnYJWKdw6o0
4ez7rm2UTCnxv8dMLEQf0N6yVujpuf92ELxg+rwZvquhMeEpgFyDZDTWSsBe
gexEF/7xbufAlVeSRLWDiREcGf3pH4P4wnhOU/J30bIGOfdbaUl1Nv9ogklU
Ppl9J/ZenpMmM3XrIRRvt/wXMADBkgcJBX/eLPBodqG7JRRM+hiPDnipc4Om
0L5srXWzR57AKQfyr4EEPRSvU6gaMmC+a1iCLOw3MJHU5F+/VnBi6Ib1eTK4
PSovdQj4/pnwFSg8qCg15wMJrdSIn+n4q1/ofxplWFUPd2DXf+A9I9st0rIl
E3EYesn4n/oEmBojAd+DFyEF0IxaKu1U6clebJYIpU7GUpgZoLGD71HrsGp+
Iz0EeJMsMrHvFF+PeKsKcxnoxqdcb2lCJTOsdlSEC4x2bFloNHOCaIZayVsT
8N5oXmtTHq64Or094MlLt0+cIPoHiiV9IOpE2FbCgyyXF/zPf+UdoV+jZ7La
s1/R8Zoj9WGYP9vL0uzSleIbmE8Xltwb59OyAwYD21KNKHSl4BBpRk7AwH5h
H5lMNu+hScS8XORL+s8xuzaF+Ca1eUaKDg5NI4YJFyr7RW57eI5vBwBAdI4I
OFKYCAwwAHssVigqcj7koFWLRtYEC9W7OLJwGOnd8I9CaA/BFLMYggspw6Qz
feh31t2nt/ImnBRCTKDBdDzoF8pIItV5HgvdD06KGD3QV4CdiLyV1g8jOtdq
dbXSDtRXu4vnlpiKftu4xixuJ55icy8wuJNzLFh8LbIv2MrwsOFLslbg3ee/
G4Cq6XgWwwRG6++NWfyYjuLjy6aNLcy5u4LnFWOYdRFGh0mJWNc71Qtz3kWX
mnVAJoIhehviuV1joCb9rBhkhs+qZsIDrAZbUrJ0hn26+VP+A7l2YMU9BcoN
VlbuYiYPJr+Vbp3klam6mn7C+D2mvtK8WfFctMWBqklaWRqb7hAjYk5brGcy
1zKhfOYsd45s8eO3/0AvDdCK28P4G0R8mBHSzH/AWjkbXXqSeEHxeC0aMrht
aDPQG095gc8yzp8B323LImcjryNoGxUg+g0iK6zyQvxFA3Yc2R3+bftfD7kh
7rQeXVukZ5mIHa046XtwoeHTC4FAd7I4NxALI4soOR7TXfnV2Yvs1LwCCxwx
5//r9Nkcoq1CLGvD9aDmHoUoPJTi6Qw1w1Rn1dBRsOlVsfQD/nubnhorr9hv
uytWRRyl+x+4dapXD7saICr9iXr20VwGnwgo1SpiJ7CPrvs//lEPf6qr580Q
Zv8usiFmrbLVXsjhPa5VjLD7IS3w9ixdgzPbXRA2/ZcQUKhxXlVqDEvFSfvn
fzarRxF+qvMOFR4mAF7D9J0VrtAPeIyJLiLbNw0tFIjoLBZR3QDm4Zbrh8/d
msRtKPO4e0WwaH4JnmDLBLRHOKInnXz8GtCVwRoik5WYdbC+lzT3Jd0at2jX
R6TUzW9Es9IiNs579zTsae7zC6tQ9Ik8zU9/iMVd4ewTMXiU6eFjpcKprqQS
IrG8rORFQw4iPDcnjk9UCWFIWq8pU272vZhvAuLj0QfaCpzDyCDNLT45LmEo
JbYO4Q/4Te1uI1uarna3s/3V4skl+jlm86s9YRyqkbVz7lxDsUwPt8dXj7x6
40ChCKbFsoiR7jXAg9PBDiiB1KdY/CVzOSg/OTn6v5BGeuwgJVipUwEalaDV
zgiOIYXG+Zct4rPJxq4kX1U47npr79tJnqwd6wZdtulROaboEDIuwj8yzwXS
HmRfODOKzCOMm80sGGz9vkPraTQBiGGnqFckcc+AFA4OAHCoBFOWLkAxQiSm
U3kYZE2KWNZa3zeplw2FzmWmFRq0s6hBwmON1TTjjr3Jgq15r7f6Q6Ej8/Be
CgsW5eOG7yF2mMsmS7qk6WixEApn7+ZCpaaOXKO/J4anrwNyu/Uc4yEg0EOp
7Ie1kSHooEp2eRrgsOi095Z2a3QkXQXKhKke27QWmmLe160YDpzp8BrdfhfK
2BV+mV2lRFmmmK4hU0muTgU4ejUyfX3OoNBRutyMDyrygLi53ohIVxHNfVaD
7HP5BrS6TASg20p6vFsU7L+CCF36XHfd/NOyTdyy3yg8lD0N2Wp8hJjzCalT
P+ea114d5KwgUE3pamKIeOGYJqQiCavWseSRZ95TjpF1wSNoPt84nY222haq
sPT5XHvYfOOOgoMKPblii44g2LJlwvzWIRzlKNbU8Xqk0xGe1laHELHBSXws
39AIEN9sUy+QFKTL2P8lRMzumKQnvJfSKC28hUgCyKpZl7jPI4rLBNujgZl+
7gqr7kG9ALDJ5dY3Xx7faBkrUd1Fk88ta6/+D7ylI4/Ia9KBqzAqO0R+NTaH
EdJp3qx4TBskccuK7Pyeh3garGJKGtn3tentbvB03S2xd1CpXredt6445WZH
Op2SaIi2arg4fd7MOhLMlUcMWUiKN3vNvifYqrszl24XYhRoedSnzxi72qLa
rTBTbNH07aGkNVkWvqHKxtNhYOsokAulXGnyq4ZPQIg4hgIyKpXhPfMMgf0H
E4ZMOjPz0XSkNqYFCJfKRTkEEDrHIP+2uADh1L9F2u5gArwtK7gg+7C2w0kA
zISdmm9c6eVYz9obsKKCa6EM/0NHwSPzpVr+b/C3hyT2b2x2IGoqcvUYNufn
xxXHYGVtbYd4tDw+VAlWfBju2GseifVqS+fKCp9WzemIxGMGVU2aw0FJA3cb
zZeScpWAZy3I0fIE0cavst84JkQaakMOXhkcTPaSMUxOWnEPkN7iCdbU25xJ
vvLWW5J0pQONzjbhpzJuagLNULbhLW1dioPVkQA8gdMtd4b/5zbSUhbb3rS3
h87qTbB6ETf/la4pNlc8TwQygkcXSG3QspjHzr39VCn0D7VG5gMxBTnUuFvU
czr/Hl9irl4yywkLSY0bdP/MqmX/VbnlTavNjWbdR3Eh6EDT3NtqsxYp561n
7ECUE8LlVPN+4EqjLWdqDw5MnWWq12RQwjrT2LSl41TUp/pEhPxNmrnHpIMM
ioP+D+t0kddgFEKjjgJwNuqRtSI6P7+Y4JJInOQpiS4euP5QFLoHBoICGK/U
1KyNCQFoXl4Wnc4uQdcishC2MEKHQT74jkt8e+fbrPQaQ2Ow+exqp4IN7mAl
L2pjXkrNZ7T1VZDcdVWw4ibOoTB6VmmQxZzd2Jw2BDJEtzG4pCFxBpbdMnIy
ZO+4PDB8heH0y8bnyXpz/2nc3g03bcfQJmpruplobPeP1adIIph5D3/bM20v
jpXP3kkQyz5sdRBZx9lGI9d0sq4fgBgD/549JkquQvC5Iy1UaQPlYggdm3YM
uzmlKMotShYwM9qKAtIa+X+QTdYSX7SxvEWONOKXe41CFFLJrIA/CrqaZLuQ
8CDzi1dEqfPuRW2Ns/S+XQzEaKDXy0WNG+EctOInSd7iKv/n+R/OdgZPmOMI
aQ1UDgjRcBT8/V6VClXRS82Fjq6wWf3uUo3Hvog8jbJIYUMyI5OYrdAY2oDk
CPUZlwDQ9ysraEQghmUG9LueT92CGEiLQH7qMHQ+viOD3/eqOUfvcviIeCGE
97Hia2C2N05lRfwTclhwRaGOlQfFQhNptJu7YwB2SOUE6+LNMHbdHYPsOQEb
N7b55x0jp4Qq2pZXB1lNhTW08LmzCzGL1RogZuQY9FHgUQImsI69QR0RqKNz
mq8N/Y4724o6wc/NetJOybHVdaG789vyTt9rB5B0uTBM2RQepyK7sqhmVuzP
UucU7+xJcbukOTfKjoSfFYcUR36s228MV6RJrFivde37dfXurFcGdWJk9P/o
u+loJ8Q+XMMtQpuqV9pAWjAIa8z7FnmykaBEnzQsi/mUB8nh01xYcR3DswXT
YjtwL9aSYel5k4ILpd7BjjUYe8UBFtjS/D0hFGfNXazNlaP8+Li2W8uRVNQC
PgVri+6rY/e+s6Q+us3l/GTl/jGY5rbfcnggBZ/RCj8J1ys56yhGRjaQjrG+
P8xNPOEKhuKOIt/VIgQT5CXDog5Rwx54gThNAa2H4tx3EgfRHf2xlrcRC9vl
7LU/ASSRmm9DOjrwbRteja+0GvN9G0viXdV1iJlXXau394DpMrOgotYf+EkJ
ArGxG3VQ18IKXTHrYBIaxFb4WfNDj6CX7HES/7Ou0ivp4BZ/76W/B/rCIsIQ
CI0CkzsR6zAOIq7ammpZwjnIPaUngyLyoASZFPj683sC4YQ6gInVhPlgQ5Zg
+QtqZ8LF+IlTl9Z8nCf+3BMaKZ675AUj+pShx6ZclA6eM1yaz+S/aC5zyDeF
6kSYBfBp/z2EuIGX39zkZ9jZQUN+TQlzgAIJLFREVWkh46B0S+o9TSI67NH3
a9O5+dnooGT1/sT5Vud1tOxipIisfzLVFcADYqI+3Qgubrf0D3ZiYSXPCwHV
mg5+32RfaYiSBt/CtzyWDUcrdDpp670ZLcGvzyxGQDZZjeh1Xl5mJcHpqYNR
5bvblPL9slMjrbUMop+/yr6ldF0p2wEoZbRB37PDOPSuBx0F9zB1o7lYaerz
MJM9Z9OYSuAUcqcfZDWGLa+DyycMQyXhyX5H6iThjO9lkvLQy6CfkLoUO6gn
PUECnnYzYnDQGSUAvU5C+Yzx00ug63OmZp1JdLnXPnElxTAzXi1AxAMDmZ6R
CiHxSP9P240a9rM0wehyxUdyUQkKTY5HcJ/DHn8PcRlR49Fv/xf1IFJ5i9kb
Zw3V3O3Nwgu8r2RZkYZHm/G77AUGmrhrobQ2w03HqoN79NlyjI1ZAHeflJ/v
LSGehHrGoR/kumeMMIhuqdWo/SJXSAYungp0IclbkuHOEvdlmRYuCEkXbFhS
1BBHt6YW4aG1RhR8HFdqLD7+/jS0h7BagTejUfbJsZWqFRAjalYZRZRSXS4o
nefuOnls+3/kC4T+RSrRQwVHqkOhdnuagY2T65PgrI5BGEpsEzdC9bGhyoK2
IpcCudey9fc6w0ePLJwRHPnqP5Z0XHZO2m5fmxmurRJ88DlJOpldHqO0PsKx
GiOihZEIzBEGGK79RDWDc2pORGmshSwxUk0TbS33u6ICQPR5ghcKxiVeej+u
L3DncIyeF1CcUn0P4z7vanOxlkB5UHwBI50jZpEQMSSpOfQNVEudEwCHkFZf
KrYDZnknCMgxe2yWrAp2aPedw3SDzNfsNVzC5aSp7kTuIrZnFZz7KmhHsOa6
HC7HAi/jN1Hgqj6KhUhEhdeFXFo+2uO7zVTNkl5HRiZXZzg9F5x9eGHpe9aj
QVVDjlFZiybOo3w476PxAoTXmg5WUckerlwz0V9QXBJL4+25iMZd0K872oQg
wUxgnXc7Sz8woZ/3wxj0ql0uiY+nwYOeWWXNlxsP/VIKtQcMn6TyTnRzL0Fs
B3NhEnfSZw+GZ5wPqwPfSDl6c1dKf2KE9vpsBgoko18rxQ8V0shYaS20f5Um
Z0+sVNqXMwjGkt5/LulJpSt++1ccfftBF8fnJuzwguE7zHqCOt5i7+dou6ao
se84sFC75dXxJ5IMS5N4jrCg+Sl0E+4OQMHC0AICiQUYhd1gK297GW6JNISz
/QhT3ndja8kAvoXV/2h0yCFsrtQ8mAVDx3DzFmbAwH9IXD+aEJZXTAJUVL+A
4eWHMu0vsZ3+Z8DmZKyecA4nvcgWPQDlb+JJrMz+fOct9Os/cy6nIrqrS25X
o1IIfNkvxtJ3CJOXl8v7+7yjSj0dbMnFshbypref9kquP35oattevHZzLAMu
b+zBNaUjOOJkq8nmGPKJOkoVxQ6V7+JKnNxFYWZlbbr0Fw7JgC0s1dF54kIR
f8RQrrWJIbsSAJitjs7V2FJq3Y2xyeu1UL3xui0Nr0y9If9pIeNh91izRoSC
rD3cGL6rTHQKsnsZMA+yhH59PD9+KGGRxYrKLWz/D1UvNc6Zuo48R+KQWHhR
yVfJRQpJjsFrS89lLtqKnNftd4/TWfjpUy1w8++zH1K4HxsDE3GV9zu0Amuy
gOX3ep/mpfb2iPM+F1iEwRbSmR8Wi86E4lQeND0SBdrpyFXe9IRqrOuqsjjy
6KcdCszPaBHWEadwGVbr0Moxw7C5pgZigLRe31tG2E/U0QS6KYOlf4sT+cKL
51WOz+NZWzqMMkOv8H76rIgC+ZDaIdqE9sgUECbHnAj+O3eWO+9mq9h9Si9f
7We3SZmS71Z6QkgMdLK4/iFYtHNOuCxoPmkA/q4emmsooJboY6PHlYdMKbNj
cSmUDrisQjR5TMZ8t7tDyidDRc1JfsM+U6IEojN68x+66czJ61RmwSSsVl4S
oYvtgaf/Wd4Q/imItQzBvO0ylpyKppNAI1E1rIE7qCOKv23//J7frloqB8W3
7cqpTc1ia7DOxzHxfQHxGvlnjP+b2Mnq9p9tdGZM3iufke8FVKnU85Mf4g2t
xnu4kv4dl6rjLMoI1GDTm63+1gwsZtGWyq+LDTBeY8yUBX6e0CX+GFFcYm3h
ibbTZFSdJDLPm1y0xAm+I/RUd8R3/+9tR00CuIkz9uRoUFohJIvflgiQg2So
2I9AdFir3wT8/+1CQtO8u2/mEYWkke2Xj41SI1ih5X9gpitaps90kfAMIHPw
bflfd/eislH+x9yleDxd3YA9TdYiAtoPhZ1tR5TglYL2zWrWbbr4rwKpzG5/
UfWaHxM16OmLWiHZwzvyYwlHsfVvuuXKaHXAF1P761tAmxG2Csi3bMZCPLXZ
rSFG4WoKZp3ZaX2svSHehs6Os2ZeAEX/wyWkEiCoMAx7p0oYCTAl2SpiAM8h
M5JNSYB6bwl+4Nt0+8VhRsi5wV3IUyW1EwSDZR2JDPvkZCkK0Z5+ua2Vu7UA
OjerWjTy2wbOT1tdIjWP1E5qc+5NLoxwqdiibi1PrmN5wgNv2+s77hJxXEUL
NEuAEB2so7PZG7mQNl3Vn6iEYnHSKuwfXX+10zQNN18YjGAod2ZT4cff8bzr
KHx80soE5A2PY9IA6hkRjbeP/GvyO9wIQOYGYq51ajYlOZYUA8bmN5WqNLTy
9r6I6L6yK9nEduFrZzkGrQZkqWo8yqc5wrW8eZ7AKh2wgTHY6NarZwQP93cI
7yKNqH3Ta8/52Xy9uWNlpu38ou9NNuUleuJQSAtUbqgVCctNvW9MDzosrQs+
FjNmiXVk3WWwWQF5ok91cu0/YDZdn7/qwAbkFBXouyMQWj4ZFlJQosfdGXGI
UsA7PmQH4mdf12d3ySwsLHvLhtYpCO8/f3D0AEojPp8fUdMn1Zynre38NrCz
tQz/xmENu8rey/jI6z7khRGalXCAz0xa6XzEJyoxTn1JtZ7d6BZLsfViTC6a
jcLFkxkUl4iiKeqEAFBbPRte43zZ8HYGkoy3Oy34f92gBb0QeJjiRgyABrH+
x1HFkczwiv0H5qQPtvsh0VYqqQX3yvpW4J2hXIjCQev2PmIn9xe8t5CBIfPT
cq4RDTE4eb2mAbBlOq1O2+JycNpb7FEed5/2VXlz0vCM2xb5vPa12Go+yY5w
ttkQNe5k/naYJl1zNtvsd112ODRYacPLvQhgnlK1lwLa6ZOsYLxP0oY6inEu
YqueFPmtSkf2MOpsySLkK15MPMv0yIdkBXc7bfK46vWvSV4WMWkktv9iHEWZ
bfhsw20YdEg47s93WpSU4YzNmKHTHp30EEqNnvqNCohyKWrp87zpSwO+eBMg
oe1kXsdFFCnsLWDDoq0+JqhcDWmJvscP6qLxQrY7BzDCYR24I6uEMDwFCbGM
5ANO7WP9LkIfzITjDkFf/v9vMsCTulL7q2+aONclhsra+A91xaunnZrPJaJp
dwT4XTekDX3lVK/Jhj5rIQiVW7WDcqla62mxg0+hgUhPcyt+6IZZxYNcXceM
LO9faBIIfdYY1+gMXdRtdiUW70uDxK0ilhOaLKSBfzlF5rzl3Oi2HjZbcAKC
dcN/Nv/ZXK4M4BNdjoHOv34PIhji4KGaP4p3NyfgRgaIMjDeFisvzLp85nCu
Y5Wv3fikUlQ5Rlx3CAGk/oG0XMP84i34My9utZenWWLL047Py+BH6No9vLZU
PfKRBQ/fV45mFai8GrogPlbu3s972SfvnceqJp6G1j/EEvzLaD4fmJkHqKn3
IMtBQunQvyJ++yOP8yJn09qksdtl9yi4ewFdMUtIKYWKeDfPKLZWIRMzvVAp
8udSuusaaIYWqZpfY/IkcfbcGTD9SX2R1jkvZkQdqTKFUHqgylts9tO/CHsZ
+yAcqjrbcZNOTbwwxEhpjzjCLaX6lYnMGRwDBI+Fz8uJp3WAeSRI7ZeaGrE9
IZaucFdoTHbU/cGcSJlkXWRWwVNR7codmRiQC31cDd3fi8M/1vZ2/4wflqgA
pcwLC1OAZGWlhvIaVl9tATIB5/gxk8lQ8kIGTEkXvhrAPwQliFuaK7KSKEf2
xpNondFrR0r13CnO6u3qVDlAs5MlpUg3Zu/ex6rAzMfCDPbZlnmICSchqPk0
GnDM8dqbUJYBTs5BSfDdenLYiOl+EGHLztaRXMYtDpc3nulHRkzx8Ip/MTdC
EFCltt2+xtl1OstmS34YFDFxjqmVK+sRxfndgBf0FNnU7Mb9P0aEhZRLGNd+
JVmsjXKmesmNJz6u6dMY/64VAOkv24vrEhyLoOmIjV9dtERc+JHr7CuIsUYr
5rFQYP0kpxsySKlWULGwGOWUIHt28FY6NFcArbD1PilR9zIblwV8kvtxf14m
Ru7yGMo4X4dAWuogdNz8e+0GjrzTCnIRMJe3ti4M9gfQ0YFXBuBfZ7EDbsfx
LEjJ4T4zvbCUaLlKLGuuVA5tWAx8OHhfZYK6NFovR6xVPnnooQLVkcKHAohB
b9B7i3syNzX1UuSmvNgfy8hmfUQTt1MadYU4LV5asJTVBo8G4qV2dZBbozuw
NyIvp5I8uQ4VctD7ARWG4I48nLqTvysQf2PTgdFw2LRsaPygPjCKx2YjzE2A
JVWrUj+2txCDxzOMX3WkoCFBzmAFf3SETLIg5ToALG3wn0HS581rFTN/jZhJ
WdE9KMieui1IpdhVmX7bnXKMZjV1cnbBmvptbpEk50CHsaqPP+x1bEiWr0H7
6hZBdH/eYZ5na1zKitQsGawHOi+BQPSEpldgv0ZrgdmxsjCwaHQWYvUs38vI
I+br5FmZwV58grL71kQlwiHIXHa11JYamZnRICBnL1rXX1lf/bQ/HwwKq9Pk
iibGCRIXLq7TDNtVNn1SNYLQP/6cFThtTLPDzuLnAs5RuY5JLNZZ6kJHA+cO
CSSTF9GNxeyckShC/HiY8k4MptBB13kGn6tSq42t10jMktLIVgpAkpM91ZnC
h4EJhcMPi6yQWmqht+KDtbnybx+PoVq5Bg6hHrfCVOuhazoSRlGwDaDjoiN6
G6oUdgu0MTOlqy1xqEsoGQUJxz/gIOs+kDFpL6AVEdZcajpvkiBj71rc+D/l
PiktY317v1KhioJSMUD/YGbSaL/2Jv970OZwvy71R6CnjaGAsf9yU128AQ66
7L+FdVy2zCXmVMw8jHabp2bjt9bNiDsn5NSEAVer3ZXvNSixvnAKmDgKGvuw
QT76pwd1Lo5gZaBZZ4gz9Z1K/FNCWVlPlJaQrmxgz4yKMOagy1jSgkUB4Ps8
MzS4JH3i6At6a0uN+sFwPQz/YUxi2BmsD+W+4TlBGKnThJoQiYYLgBVKkHh6
u9fQ1JCa7UC3SA5GLm/yLjUUz7V54+xgSNklAZ81vauTiWlpeWelUCUyWM7c
shHLsS4TgWfCLP8+xqwBbEF5UidAQbnbHKrpID/Y3Pw9BfQC8BXfmbNrq+Sk
HCYRyXSMPHimhplNe9xlO1XfhZcRRZ5Zbxe6lfNt13S8lE1b4NUtd9g3WFWs
Ye/Zah/xyrp1azAVgTn+Q/ywgsDXp7+7pc28WJnz3m3UN0qQKwo0oGRtGu32
7hCf8r+rneSk7nH/2JVrMrSua7NYXlBdqr9aaWrzbEfbgLCHB9m9GF52EuTS
Y2TmXIbO2BlZknqAC8ZdODzuODh4yw93EFi9t051y5QXyoJdJFfIp49ubHvj
h9k7z4VtDvtXsP5onSCmOfYWXr4pePd8Usc1cQ+XRgrONb1kPGk1zg4MF9u4
9TyLVteLATWuQ4aNb0JueBes/UWoclBgIaW0VLUnkgtTysHRmI5eO4pEw8bG
AFiG7+8ebuPbU27YIr1tj9ZQL3kY9+oeWj3/81mE6JXKIW0NkcrEjGoBlIPB
Hnf+FsRTbD0SPGVfFNeh6neYHZ3kKjianYFVQNL9DfJwB0oPTF4FHVxWD9+h
rsnzmGuKZu7ONnsk0yHMSWq+//gWcoU5B8bmr0zh3WD6bgNeD198MjH9Lpbs
0xNpukiSjDRn95mbj67Mwd4eksdZGwNRoyK8on2bQfkLCNa2SPp+lXmX9KFR
0lepW01cszRs1ZnSJA5jCc45AYhZmBuDICLBm5c49RWjqeY6/2VB6L3Zegl8
tl6A5FOG+zjUYQJeING732hrV3TmwvsGP8FrRhrLkVEFh5eDLgOTGvtOLbfK
UlS8ndYf8LrEruAOAnlQfCMHf1gN2chFERTtELUmiFew3IpEjLWP/CJmaYC5
OsnOpafE6QN9wOS2XbJHS9gOMd7dlBH4v3WOkg/yMsHZWKv/LQZB5ZVK0qjT
eN1hEyW98ZbO3wLcwd96MtAREAd726YjxJwse5+C21VT23nfr6Qh+UNsRMPT
ixz8dmUIue1ESVdy4T/D85PmL6VcqCTfFBU8Dn7TTru3n57HsNcwYnoDMoJi
uebPwXCSbtb8gMxNkEUfqpfLDSi8Op2WNNPUhZT396upnRi/ndbkXvHPT9LE
+eUDUUX9S2ag8rGqhlCTEArW62s1z1ebGiFLTBH1yKUEIfq9eCzuYNh4xTGB
OnXnc0ePJPS4asd0JzwVdDa/4bifcjpNDVzMoWK/uaUMxIZFht8qIwAWQytr
4yn/q0Sc35YanbP9Km5IJsLLpW8Ljef/7UVDM9B/p/OgD5WYjY7P8e4GOCIn
qQaR7rMLCTB1yn/ZK+dAxLa6KkSgmBcCnT6KUcFdUpl+43gN6Vga2YHEayB5
IwArcxv0hBDsMPQ/0U45Yy0DqT+E1SJaY6BrtCtpSs/AS+HJhmnLEPJtJk2F
qRZu8iKm/eVxhJYO9i+EHiIuTn0F4+mOuzpnfs3ZYCRvCMwLKPPdNSRPeuA3
5PldaREhs+GzX6dznL0DTddGzjgqvsw7jlhpajiYmSrd+MofSf+wWuxY691F
JWqUvTEw03bq/SmR29dG5voWISdooUGcP37oEokye4Q8FXnBCtpSNMsddbjQ
iIdvv1YhMmACynkKIL9xKmmyw734fF9IYeGaLmjoJMEz+ShqSgP0YvEQqTaZ
pIrdzJuLQ2jOhWbFyljhE4v3Lvmd1dY7I6zYilF879lBDugCBziiXOSNkGM0
C7oMN3gI/XqLEYKZSq6Jg94MwFHnBiUcpp0PxjAqg1QqYoS8PkucvegiU6dT
IU7L0XE23AUhPc4+kuSlPNk63+8wCm/nen1oniOFYaLk5+QeUySLMHSa/PqZ
vZ/oYBFZf636uSpSHnTuCSRVTChc2Zu5dfQHIcUOgre2r/g0NXvx6pa4kYXX
QSF+m4qelSqx86mS5bQ9Qy6+qE7Lkf43Gio5h/cAr5wv38dyeuMKtgvqxeyU
MvIylZfg6qaFSkOAaOy4b/Nuj9P0Cv9hnMwnJUqaPds+CozaZcOMN3AGDh9h
Fdojm17PJuBuShCg3UG1/dLF13Xa0WHNZt/4s5Svz4PTHYh2+zS3mLU1sYS5
zpvnYxtdYZu1t+s7lsLeFzgkS2qlEZ0EWhtzaZOmrxfUNyXR91/c4tj/I4Qj
XbORqv6XHnfAmjgf1hednXEj7e74xISRJCmWFsIkmxhfGJCXAdIB6tcaKczQ
PUmQHbkTrh3GjlBZPFRVbBQqaq+eqvJMU2g27Dq5+DdknYTtrd3eGnRc6VJ6
UTgV+HUxmyvpagKo1SPzLexNQZLDfzu9gOWDyRysjU7Bi7FdM2jq3JD/hB4D
DRKVr3VMaXv7k22rMRhGbHzytt8zL1SsQxeP+hvDLRD8symaUAyIndDzP26P
SnrvrJ6ebx5hRZ8OXP7jQ9N0UJaHf5k2cEXvQOKkHL3sVcKxyQ+BG0h5i6lc
+gReoifBgeavGmYzZUWr9xPYwwBl7ItPOg1FvymcPdJ5BDGQHT+RN/WfR5WB
DrHdFF0jubEe5GeM3WoDvo1L1tR8XQcXWbe9H9uDXdmgBj55nWtgNcSMQ0WN
clKdeXdJ2HE6vDxCILsBsBW7GCX8e9nyD9DlHZa40tDt0GJGnA3igl2Ex6Is
6l5pqdIVaVGxXNnAaIm3V3p8/Pk3Letx025YotUJoJk4icBRVzV/kT0x595Z
MTCcTgWz1LrknLqR14Cb+jRAMaSKKkUk1oJUH/Tps+4c/d+aCaxs5WiiDuQn
OXgnxyRHGpPilWAtFcRWGeo+wdAsiF3a5drtcPuB/VYkXhTVpMoHmdg29eKc
G/1trqxjqrX1FFHaeBL9sWku8GblCjLLWvO0+XVL9eCLVlFAxyMsnq2ZbXdQ
WzK8zbORX1SOtmxdCXlw3gXGZzBZYHbf4+BliqLhSstKApZpIJj9C5wfOFRF
wMZzf4IovwvgJjX8rEqqOJ3a6zE3RQMO0d/577Pgh6+fPcU+XZbPXbev68Zx
wm/LttSV7mYvR4FkDFqLOuBWxM0uYdEGUdvxoHCmu+2bfjPIMDqj3/mHqkq9
56etTMJZofJJSIBu9m+9+UY07WaVkPZu4Iz1DDEXgB07KPxK1YoXHAY/IABc
zveV6waHbOZw4vs0RlihpDrTYTXa6Z+KaM/Edt2z0oZH378uCteFlX+tNDuk
bpBU1JociWAIfQV8P4o5r2LkH6Dl0mKaoGqgU+V3DgPn12l5AQ2a/RqAybQy
tabacPkHzQjD/jjlvMy4h0XsJHI4yPG9zNNDRRqkBaUqDOQQUQlnRi5gXmBQ
Ux9IKslfFKbkHiq+hRqJjv9CPavj9X2XEwj+5RVQ739At2vY0fnkQCrXOgc3
VMQcXHwJLYAxeqwEqtnl0wg+MaJg8WvDF0KHtHrYS6NFvpD4pT6i5FX38fjv
Evk8Y2/hA/GIBzM0MBcrCXyDpq6FUilQojP4ECzEklnzJratgNYvnGT3YFc1
jYtzis3PTZ1f8XZ+c/SrMEX05tlVfoK+FE4/QIP+BcinF9xSvhZGxzXeDroK
JlpQaGGBltQVf8HLwkfgVcECDOhkpVuSZv2JEg3rxI0LMXvwHnVuUBexcDnL
2LxXTWioCyFCwcBlnMhh9j3tEgKZVYjzM9TXex0z+z2HoLhXePlUQ2CarmtG
+jkQ/bcJ3PB6XWxishtMN5yFWsFUjNgKt3Z35U+zxEaSkKf9mN44J7ip78Fl
2Yzi7nkIQEkd+/lLBeA+FeTWLCgZR1/NWUmSWbHxc8dCt2fR3aph9eMbhaQv
IZio12rHhIwrNbt3JxbUdNJGZTyL6yDU33bqO1aMlCluZodO/88wP7ojD7vW
12a/mEcY0cwx2e0CexuJOkDOHyRL88Ps23qmOOgwLYvYh1UuYzD2XjrBCCOy
dvmDaNg7RcQmL6RPW4KTyDmo+MnoKd/hHDnjkFzLsRFksEH6uJjb9cXG5Q0B
O93VF326ChLntCCdLOIpQ5I4nChyblBSiXJ/IF2xnE2yApRbdpR6R/C36Qcq
ypwz8qCRzMFQyQBqq7Z+U5fYI0lrPneL4BKZOmmbIKR2Pc7reRRM/HwhdiHr
bahI5ZhqCEsTRgLT/QBtwdks97OQahgVc91k73NsfyI7B/Ke2XH8tDzBrtDA
F7tCDBr+a1oLMutwyEsEPL2xBahK8bfSaIWPfbYmNqdGkt58JGo3l29SMgDb
L9CHJ/HStc0+LnQMNwMNN/Zcm1YN1C7mvMAraWmnAKhZUnf8vfSkkv0n3fnH
aNMT1oVSEMp9o9pksLJM3glDLY75TBT06GRfmZO/CC2PGORQz7DjJgj6XkIJ
sJ+WYraotQvkk7PMqRxOomxO8c2wPTjF7RR8iQNx1kkWGhp607k8bxSpKVmp
cZENbqVaqpLbZyj5LNCn5j0BXveyjD0L1Cb2eJQJmxp9/lTnp45taIVpc37j
ao87I79SNlAo4LFiO89/nP6Z8FaLf7KunmtTyqfjRn9ElQ+QDt/O20ir6loA
gKz9tFCvpJ53A290z27A3+UVWltQ/utVAmT1MrwCdORRUL8+tQwAeXu1nuEy
loR/S8+xYRA9ZRaUKE9sB1YJPn1cxfVAX72F2Yba+PNG47ZVvNDiv/ty+iss
LWOqsjOUY03hy+CKABJNod+MOp+Awe0xZRNR4UO7y+GyQqj2KPkTPdTvDkgD
+GWrLbRw+J9kOwT2chKM+qYLqSCZWQX3d28xEp3WGM3Ahp8MMZKapfIktksX
CiVdPIZCyrqVqHsn1JdZAgv/IGZkDC3/1/u7YI5i95epIdqOdLo0wYKmzlKw
CsjLI3KR5Pv3fKG2xmhQBWIf6YSh2vK5S6f3TY1E01JLKcNIjeEk6MoXkZEs
yHuou2hxSVhuhhxjlYoGCEyN0USEEDmbByTVY0S+vlZ0z1exKVwONGN1jGhE
JiAkxP14IsRdedPQmQmBji//id9XDJjCymFD6AS2LgTYZyZiyI7INzcStvLS
UjkYyjjLoWafjuc4e+EL+p1h6MmSuGTfbrZNeVtTMnHPD15Nh93f1Et930kY
Nw2abGxdQDtP5PApAJQk+Unl4hOzgMeqC9z11OAgzMqIg1Z5j1+LxrTAyWRs
SmkXHFW+cgzU4BziIrcy/dVD+m8WSKrta06pemkGfH0UmloEH07XxFW1SuPd
mDZ2JjlMccsRHIbFcAcULJgm3cNcGBUsprx1HizVAci5x8r/6POezQ0T86Ii
PSYUhF8YKSLKR6C7LMyeK/zGaFsadO+ckdT/VJ2zi1xFHpc77mkJr9UjXuUl
M8qhs8fVG5FEYJQGIb+X/n3Ez1AmF61rshU8eceJW3+DEFQF2R1UOW4aYRU6
9eY7u3kQHfCHFcYUgq4l2yPojVHF8cfJ3qc6fpZuTS72FkPuHmd5diLzF1m9
ilYNs0evf4pup2rzg4/G/rxLvVCbR5Rw2t0DwECWYb12FxE79yysOQ7FExKV
9pl58/UXLlMDVGQwRxgg3sLTsyZbrLPiPPYgG9QLdDYd+qNUTT/VnZSfLKIw
AMVh9xATIgTkp36hkwJpU1XYJmvflF/0pSnzROlvD1kDPpiB5O8YjtdOsU3i
Ijr0POTYSX41H94vz87dIY75c2ND248PwtixpcOGgO6CZuuNJZ+6+YW1rgCr
G2rOvnfw6Np7ISdk/V+AZlp0MEOttcDuAwMLRC/lfAHZp1Kd+rphon9pQDqx
GMiy7jPzMima/RCWhEE7mWK/sQAVGQ8iuteNxxcONEPZr5/EciH6J4yK/qjg
HVCk/Y/N6cnVMFSAslbXI5yvYW5TG8SR8X1MzAs/T2dObddD/2ZnWa3rvozT
plOZlyn3vNZ8P2fVuqU5OmSbFPXax2RCDss/+aaJdGYcazOG3paVaRHNC0uy
7aIrepGcc6NgDAzZ4s+ScgeVPJSM8w1L3ey1uLuzXofhf1SG3v7S3OdaUbUc
cB6hfBEDdRPvCPYCSZl1RfL1sP8l06fcdd/tky9ygXIkpkiMiOS5u3GX0UzF
bBULfDCcDHezVPtyphfxFaCpHKpY76tDTX+gmGnYhDGXtv9bstE4IFQLGbyq
gSBdA4Dl06gJ2+ZDix3dK8Ootmcl1gV6VKR4a/x6qgKbJ3M+Qmcgc6HKkoDS
BnrU+YQOROOKVwmPfws5vp/dNOeY7Rkvn0NvzOTjhI5f41S3S0V7Ox64RfHl
CkS8iHq8o1rERA+0uPAkfU0upzhzANxTVmmhtNTqGVir+Zpz8LK7R1dj7zFF
/VqLn0du0b+noWqhqF6y7myc/81NyfCAdtkbBPyNrK+HTVW57jPEbDQG9J3b
OKitRR6K2Zc9M6TfpNkSASQ8NUkQ+/Q7J9V+qeHTar2CW12f7ylxXuVJcndi
bcVSpM2FXVl+HKJKv3v0La4w6ApJTfgudC9nMR5teuZDIqtEK9BCdbZ2YP4w
8me/mDBqLLTL35QF2usIUEMmngcbjxwgRku1dKner4lVVeDt1/aMkvmI5919
y/BQGvIrHnJfKgpyB/tqCcP/ldaRFPiEkADaplS865YppM0e9gZzkZmvamTF
LrQziVuuj8ozaapg03n6toirgf+STJwzgo0xyITTQd+dn1iGCssxNqLNm/n1
fOZZtnevWHS+eYnNplY9zIILHEwaijwL9Q/WEcUelVYdtDOekP2yQl5OoH8i
AACj8QNwm5d4SqO38O8KrOOZg+eBPJqR2zk1DjZJur/VVpZokDy72T6VboZv
qmZAXF19h7G9pGMSHcDqIdvch7nPhMQBbDijp5+mqVnCeEZW4bQ7PR4JiK1u
ZNWH6vbybxTNjmCQNbw6FPZu6yHoQtPFYQd3FKbHwGUweLDqZJTU4sdX71PD
wSCR06s3d9qDB8d9M5QLtmxmANeFX7fjA0eGAVtEA+HINWdu1ewNU388aUre
w0oZpT6BqNYwaDNKngLwz8UHDp0Qc3EAl/MxaD3pVETlf5kvPRkYHefscAXT
vzV9fiYf8/cQwWumaE8qEl0g44pKmt/K3QbVas5f/QUzcQEVKv6UM24kvJNs
O2bj1sZ78pDeoNH+NO+RVWJgdECM2IMGVCIm4+m305k1EsRg1vQEBh+c3LvO
I029K7xSZe70xbwCIf0fb0by7R7rOnYDGfDwbLYdXS/G1NXLy/3s2eOM8ylJ
85g4gAPaiXHupTqFQTBxtGBc2YQ+u1G+nikZ9a7TuA4PLLjolqkOPu1NvN13
TSNxT6+hPmM6inOh3enFZvBPlSxp/ZuhShcodDXic2gPOZMpNo6R4X9Y4zjx
N91uKUf3TR5f1Ia6fTU+V/sufc1LCGcfO0tEyQh0TKSUb59klUIZUHxZ6WX6
Gz3J8tIItKF2tJv/sZ88BlAXuqP+HrOroRfIH3Vmw8fcatVSC6xtBhU7vY6U
9XBT/HG1hI6nr7cjU6SNirujAruVsXjv9O5Uc1DaS3e8favLz1sgIdr5EAHq
bAJXtaYvBzv+PwmtoyClS2V4vBBAb+c02i8q+XYA5W1sYyN8Lfpp6qjrp3tZ
t8qomO7XDHlbXgjfULiqNU23FXk6lUGjlCCTcKUgMCoI2ShL93KOuMBfHxFl
/WKe48fkTs/7LkgSAhIj8HHxhzj39lTOnSgfynRpaHHiYZIUD3GCxGjwTDb2
hDNLMkvLAr0mNBHeLq6nxs69P0Lx3TFLS365TiZJ1UFVYS1VODzQULOCrwZt
d/h9dHbiuFvsNXPXHjdjf5LIolI1RyZz9bw0BZ6nXzlUpgljeQjGaVmLl97b
4BC/VvrAqxOAeQmu8PUh+iiAT1kwzIS46/Rr7Be4honadQrrwkLSM4lXL/+Z
ADBpEDmBQ7hoJdt1KhBA2EiY03Pcs+lbREr7Lscqo696T8qdA5i7ZwrgxEcJ
W881VIuTVXWgfVFelImsZ143PNvjXYoJW6W/2zR0iTmPNcNB9a/Si1guw3ke
pFg9PtNQ0bjZPg0mLt8YgKiW0cgzqKMALM3WxhQxKfRqwy9ZWeHSOr79cEfh
XVwiP5V5TfUU5/g/KRSxqfxy/dOVGu1ZghaAI2CGB1jlg92mEBcbY8PLX279
91kRVhtGK7w3RY+3eLp1EpQlcTBFyAsHeL6L+02ozbo3td5+85vMmoBeqsre
sLtoYQ3AIYeOGqRIzMyCChL3o/I12cCXV9DxUwXSXXOxtNM1Y0pO8eM4Ju03
mhb99lnTLujI3svrUf9NZCp9SDoDkZsDlPnFocDZXHRbusB/0UsvmIE6O71x
cnIqLhZ0yZlsH2z9/o4qlqMQfc+7EcE2WQSs2IBdQ2pDpB7lIH8TF8X8+l7r
NT5d15ijttC68oNa4yZebS8NwhF6onmDHZe6FpGrSEwSab820YmdOgFb775A
oPUXnlmR9vvZ2/+U27xwRG4CKVLlRlIBm5DhrS5KcCKtPbzf1fXinVCmgboU
iLrahz8hgdDRmRts287uQaGxBP2BXKZ5x7bxg1lIEptcjtqCutV1sif8P7Nt
IMALANmD9N/uzA/HKBZGacSFGcsgqsvXxeSxGq6g9F8xmmbc+uB9XyFpnpWu
xyaV6I/0NgPAk879bbxOH755tOn2fm4dUn3fyZQzlq0MzxOwdAmJ69JD7Dqa
I8uCQWYUU0c0U3pMaFzp923TuRZo/oZfVcpP6zFEDiharZMVhRODFMgipCXb
E0e9VgRUhSIFA4LhkzyOJ/X0l3Q9ssN2cMTJHDn5CZOacVpU+6XUjpMCfBN7
TEBkASAuLBIU7S3KKvtMBhfzRCbKPabu/nqXDJuaekCErxlvK/FEQ8LRdSpg
e/JD2arRk2VMXFrHdJdZXVjWBQfUPChdkyuhpnOYCmIcv2NzsjYdSdsVtUFX
mGtReLRKb+6gnXRGJrELUld41bL7S6+zth1IzDFeI5KJF4e1kGkn8mOxGFRR
p7yZmm9RpF3zn3XM+ZUWCY9tc81XMV0c5uJshpyDFYI/ymHQarc0ZhZOg2/H
7y3vf/jr6xn6iug+CQ30n3XNSOm31WTQwdR2Fx5owxizX6PXhZ9zIWkO6Y2T
NwrNDy+F4zqoKQXSVhhb/E4ZGHnKj9NQ5lJOf6RoYeg9wK5brfj/VBmMQIxr
eRvs1SjMP0pA+g/glb+QDIKAZ4VlLECXv+696c0gx7UcWk5nj5AkbQUirJue
w5qlYm+ZCxgDVRg82SJVq824OH5rrP6IMjnWep3eGDeCRuyY46biKdnhT/El
WD6xjz3pLYt2sThuamosRclS9+rLaRtdnKhn0KabuXyFBv7hLB3j6czrqW+P
YZs6CSQLf4OcuZUBHN6f3+EFbWYRcV6jtzRkq4pSOETe8MU6+niqCgl+Iw4X
l1tVJbYc5suNkd0KMYM8kQczP5QZhxuvbUOuS35iDwo8oYCFaqIsQjeG510V
Kl/8j4zaTgmuHP4vMYaXE1/dizLwQaMHC+KIHmEYwNuMaMMwDS8SRIHsCqzX
wFqSQDnV6Of8/vyLgrANQa0f18BM1ZS98ozFOQMrWuUeXoY9Vx0/fq/pXvCR
glnY7K3pjD57d7820ZzWJ588WXyyRgn/T8BeVm4jWQJCtFNq1/a7IkRiCs1r
/FrmDVcmznr5ToIm7e86TLZFVwQVoH0/go8WicEsyJESwg8C+VkGxiBuq6Hf
l/FC1IawrWtp65iXYSzeO8TMnfpYQjIctUmXZnluDhFy3wyEMvhcs7bER6/T
hfYyeaEH9BL11pLQ298IHyIKIXWBfdnyyTyR+/QeKN5tf6b/ENB2y0vSsSG3
dTtpKAghM6+wWcwYN4bBBN6pEgN878SkqANHFoXtDzV7zVjDQptaC4GWEn+p
HRqkgbhmOxDD7XUFU8hHnSWMm5PCxHw/jM0btITj4F36/bZQIV4pv5HKr/pq
ckkkoifnUc+ClPe24p1ElaCQGdSCcdKGhTImtMtiNSMj8GN6no6RxqN1ogZy
341dDzrNusfLMYOjcF4zXqExwEYCyoe82Mb1aa9OzfKo/wBPZZDrNxS3lR1l
pxDEfNF/7s8xSMlfQ82vOv+wTZKCKl2dkRwaWNnQGjyubJavx8NggH7wkdx9
N1OpZ6NLZpO5/gtiBIVHLAhD3LLFs4gct9BI5MXAoWqEmYgvQiF8skY+cVu4
x5WiIBk0H99WZEXqdXphED5txcAanivctX60LurywLM53BwjxLLGM123gKmK
n4KhyUalK9DSZqm4JyWWUuXXRT1ELS/SGpWkPI3aNg2z+Cwzt6uUA5l1aRTG
6AFhtmHMHO3ADmJti6qvaPXvzVljxxgez9Tdj7NvodKB15X5h1GraJ0TP+7x
5vST1Gl2vvFFFgEUHaG0L5FClLOE7opvwg18/6W331QMQM2hLkvH3vcpJpwW
XNxqwyQAOUu49X5+dPOfni6lX5y6HVQTdTQDYJVbukut/ruXZXXPq7oVyHip
hUioaTAO2Mzlnk7Fhk5zlqQoe+TZj14eQIpzNcaDPilxM3mjkrjBoBIhnjpH
vSIKsv+zt3koibbCLTSS95iidLO2ji284ZVNrxy5gohAZG0nTkFZir0ZZAN/
+WS+7s+2JzVMSncnIj0TqIq3E0PkRdepC2nEic3M3dNyoMbqYZ5O2OLoWOgS
NnsxJNndrxcYstQsxn3uYnomTwSh44rhrFdEXscfjU37WyzLIaigSFRkb8ME
CnsDZdcICFfuNH479Ej10OK6iZnviDkIrvwRNmcpg1HO8ofcmWKkq8iGdktn
YuL1O3xPpG0UKB65v8HeG8OOuc6UHoW7ZDhiR+RWofo82rJY5Q2W/Evw7NcO
jkIEqw7Xi0+EWmuPqR/tBQVqqQh4HYI6AoXuO7PXqeuFQ3edV1IWQ8HLHYuS
eYdnKtonrJ97kt2JJfBJEivRU0/ZHZueGI2HYNHruxvJ8IIZV6Jnsb7Cpcn4
Sux4svjXnEvK7rag0VUIrlJQAT5Cs0mVpaHqwgWns5gnd2UVLNQ/Q7vvUHLz
O4l9SS24aRbXVCehw4TbNdEdrnZiRihbkhD1AxFjCi0p1Rg6Rf/KpcjPwv15
WbdzH8bQTfW2o+Cwvt6Yw7qwBrDg+kjSg5TA8MQYgmOcSITbxy+tirVJesLs
PFrhlIz9qvcFziWgj7S5RPm5mbyOWrcG4B1Q941rVNXF/2fU9931ZA0SylNn
qgKH1DS/h0utRJXI5ETZkd+dnQVmAeolZI+Iouj34H00gCRaaoy/YCrD+t4s
IDUqn/DIp9f1YQ1A+Xslt2hJuQHgSDi2x1WMFbfRoRICvLjqLshfRJxVniUj
oXmWt4xHsjzYXVehc1fChglG0A225MOhZajOoUFrF1c90zOQDV+km0QliLCF
NBoPnJ/QlYiOYVZG3FGFpl3fAD+JL8/QCYBSGK615mfKWwa9piB8PEgu2jxW
cRFIkC8vwmsbRL8T2iTY4IJnDotr7o9FX/C0Tr/Sab//ZY4MSG3VW4mcfcqA
yqafDJjM9Hq4HELUeh/3CI7j1xsvyf0lE/bgVVOBJ+xg6t/8oUg4TlONt5tY
f3UOdyEAPbi/4/Zeq4Gj/Sg3st39n2aX0m5G+lvK7Z2nJHJsnXbbq9D4DRsu
C2HQl1RGxpxrVK4mkDLfkFerxcirg4en2dcT7wj5athuFSnZoZ9CBSiZG+Pu
MMmxVVEi0RU02y3UHznNK4WT9xt+sqHiGdKDyxfHHIqvZbV3CbPogKjj5VJB
T9LH1vZ+ZySd3fQOTF3oBHWfmT5eja9eWcBhM7CKsr2fBcb11hmCwkZKWt/X
1X5r2jav1xowdH7x26VtP/6iNXUuruQvJUxnEFePFIwQATe7xFnAarC6BC37
DIXpXatxz5D05rbLTXk/2uofpF5No+WmTebTjuRS2ba1dLDJs+Ah9x9VyV8A
DdSsERwbxH2t8CdNQ5vVTCwMocRg3mXAyyu/XCBUvO4Wz8M//p6ZyhCpXFZU
pVlBlsR2i9sUmuJGDBfrLBYgyQl3L1OcyRGMwyOSYTV/7sbdltYt3b85nTLK
VNIrSO9KJZUJGrGj1PkevdNuq/PvX9cPpUzoTTehL5cZeeFyL/sQx1TIByo4
rAwLFbT5YXrDYFuyre906VO+XFfbblDqdADDHG8XsLlZgsoVceI2km1kasa3
Mo8JML+oKyZblTh8YTzGxJq463W2XokJubAU197aMFsS6EuKCyftsO01apMw
hi2wRN40X6OUYy/ZxyN1mGIgwopuqIgAPh9t5O7WaWig+5PkwI/ZX2DN8uyY
3S1sqg+EepEVkmXSfAu0LoloQh1Xn3DmpT4FXGI3vFT/m1I0MNS13Z5rhl2U
YLYIWW6Tu7cYos/3H6fbmv7ixfZoz0J4buz2LMXr8I0hCHMZvpPaKYeF333L
OAvkRwnU3gg0xbAUnwmSnUL1NRsHvxLz3vPzuY44FqwqNV0X/4aEkuJL41sI
ULhWNh28AEWB4gHvxxpzZMnI5ifJrqMmC5BcTjxNlWzpSin0PBtRUUQpJWSH
jVkvFRpAikmG3lbg/tk8HqoN6C454+icrJbUnE6QnCN7VneNTRDAE63zX5cz
ZUyKX7NgafPAgYSJkXye0BQTjp/xfTwQXNvSB+GWIwt5c+0Ron4RzF/2SPyq
aT1wFOOyh5aoqYHIjsLnN5ckQjImIHJSXUcJgd2nOmBFF5C29KkGgIFRE3Lf
2PVt2e4n4diL+nB94w7O+E+7a/ocKTOrz50jEggZ9rD3Da6iDcnrbuuaYBbz
GXaUHGIZPfOgL5BbIo18pq08tkq8KXkWykeR0xQVSMph2L/1xlpADCt5IwOn
vDwdiV8PfTYreAi8t1wNDoL2ST4WybUBjJkDUDYLrVrUfVNOrrbyq5Bciy+0
ctlhHxQiVeXaRzRfhxVNAnFjvkdPqFBBGDfnO1aukXMsYoYtSdRG/1d9aYvb
Gy/z7kmOP45Z6P8wSutq/NXW/K86CEH/zVJdIek+4fz22jojT1dVu0ynh7eF
Z1uVTEDepjsK+arP28VmkN+9/205OwBdkoV4OJBXw+XCNUBlSIsSoee85pqa
Iin08eqeqcMoKZIzkdFiWpYHMsPDv94g8q1lF/H11bI1JCseYzq6SuXuR7SY
0UNluF1Uwelfluqps0KSTA5tNaVpIuSrZ9c5ltVtq65jzbGWzsJKrpPZPnzI
LVNKML4df671cR2d2HC6/qBRmdVEMWHgG2au3SpHCFjGmfnDSdnTIaTuC/+2
R2RyRZtZt4crZ2K1EUaIf+l2u9X/mQ/ipfCr35gkdyqXg3KbQ0FwYvzsCrTB
9DjGrtv3oKWRPpkRxaB0KMpi7J+gQVu7xDIWu8X7N46EPMFRNiMzQzMluUg1
lVY4a69n5EtOpO5HlMvmGNEGl3olC7Xym9Pa8FHGjNo1rrqr/o4lSVRkR174
SmQI2evOY3ZZPbroNiwoJtbXS1WoIHqwASHF6ZLR89fPOyZcJkgBTvqC39fG
lBb6fMcI4w5Eti2PBxPrerzUXWX/j5R/XWIeZZ8bx06oJYbfWhkWUYiFyWro
lQAmJ1xeDapRTYi+HtK5nuGksUEnnaiSp2T57SgFK0KXY20LCpZThoDjyt3l
zVq9ZVV3Bkt9/bGStNoYrOt/039ASKMZmnzJlqj85gOhQl8y3tZbXGsQv/nL
WtyZhbMxGOcMOG+f8aCwnWcwfPNKALbu5CZy2w9N3+0pVkzJ6wKBKUa7Oavf
x+Frg0cemky0MIMrUfvl1hbCGy+Kw7Ipw4saQTqO5qu96MSxyNVic/ZCtlf9
q8MJeGLlVa/76A2qaiCScAH6+AXzxnhVcbGC8oc0rI4MHek3/ILqPeH0gdW+
9sAVib2wNRNT+zJ2y6V3tTqmEkKP3pNYRsQaO0rhUgJk617j/GRLfSs/LS2k
14ihO9o+jsO9DGe0RTo1r5y/+j5+gQtFeLChbecadrmkaLpbkkD7WOVROtgy
73BLi4Z+t5+wcbCGQsnMFj2wxr4QaLIo4DGu49Qro0Tc1W9Y4vQyY68Ks8xt
yiOdRgmT5MmMCEebZnfRNFY18Y4ypiVCpyW9tv48revpEwnOI9Ryfa+TP+rS
XcQ9K09oaaV3ovLPSOgyZZ4DUOphuT5jKXRUhhm+6gncjBJzYmcoKo/bvVwd
3l+fV9wY220DkTRDAcoqkQRoZKRoHKWKnVjku7Jk075feUgGnbIq6tRoMGtK
HMJvDNJyjIP0nGNbNP26O9CmVIjrlwYP45OP//aArwpMpPii1U7h081H/3x+
43d1tSyN2jpm5E5Ev0t0FcafopM/27SJ71zr/bPUO3DcsNpyQPDORmr0tBq7
xjEtqd8Itcc9+2Zl5B6QL6pNi7ze1S3RKSJEZM+WDixTQS4aIJ9BYjOF/4Ku
ONP/CYy/7L6Gndkcf9qUQsNpvyUhhb2T784GEBVKhsIQizTwF9CX5OFjUs6x
0n69nr0QSE5HFcLvJGrci2Y+WX851Ub+Ws8Yf86meDLw1GMKjZKrr9BYgg6o
w4YAo4EatUmXoDuhnY3B/cuRblZl6/5Pk24CYitFtzZ5Feeq0V/ajfVQOxtj
+hy9bL+GWdWvWSwK00dQcM3ETB2nm508mxDELbVXfxZ4RJ3atqAuDgOtaO3/
lY609G/7d4IhyZhL5vRJNGstVCzZKMRWO8stXgNA/IXAhpsfCDh6AKUAvHd/
ptmKL0iDYExUt6rj1ppq748qsy7qZwKRHLSWu3rsIMJVgnO7dem00mEQAH2U
AG2YaIps8vgJTN1NIqWIQZmNvk0ny4A2yM9WCk8D697nFT2NoP3pgvIgldka
xNMCjJQUZbvZtyx1hdD1hmQXgjOfN+4aDmHMh6O26+tSA1GMqcvL49GnPDaf
Vwi/Q0tETXCOlYeinIinr7hiOaF2fEZxqz7TXB6A5nhj8QTi6COHnQ345auJ
boeZjx643PGWojvXcNNswbj1EzjgZtcPQ8tX+8MXUFjc7EUxiu19hZjieMSy
oV7Z8cWv0ai0ch855jUPZEM0n4U6XYLtB2U6h+HvGhifp1CIfDeADG8abAXf
chYe0zYFkvHZXGtOv1Fo24e7W3hVpu4Vi30sG/M60Bj7v06Wy1U6PyM0Sdre
+qLTlTrGQf9JYKGZ5saVSuU91FTvPjAqiYumbsOSuUbBlr5Xk+SpK0ea8luX
d4xrinlJG4T8FJkM5y01yE8JsATrnZeTtrunznbaIBClYcWKFiRqMp7dLlTe
8BbYMRaOkYxxQlASJnHNdSZJrlPxnE/Y2apFMTGDElvBXLZ1XvbNdUGtMe9y
11A0HeITCS2uRQQXLI5QAdDVdHQMgpac6vSEs4X/SdlShDnvkMoh9JnJzf8R
6C2Kh1rAa3rsnMtsnVVGgfLsSdT2JsOH0oQiOovdADvsO8S0zwWmO5DiRP95
i9VF1Grciba4+TDWlHZBrQQCG6Zf60caU8Tn/8NB3eRymE0VVZfWqyn4fjqC
RQgMLs++sU+y6CfG3UrSAqqNZdonPavxdREzV+CMbtNj51gsVeJEtcr6zQTn
2h4OyAJIRk9ZyZpoMrmtqRfwybtWYQSyHw6yUG3/tbgqGBl13GEQkx7R+Nce
TEDVyhdOpABMIn1yl8fZZIQ/PtYTYuVM4vtqhyPn4yqo+SwY/FIJxTZM59k9
hldZOXbhO8IqELyJIVdPZq79Z12rGlVPy+NoNOdDv0c2kqrLK3Ihggct3i5d
1wQ1qM7SvBzukrD2aqLuGVOk6v6VZs2PyBW3W3pgKJuhCkJekqIybCSZGWYd
QKCeYq9qLDhEdIX123mU0Wo6+sdRkIL7eD3hCAOafQWcGOaMthVR/T3qhvpJ
WEPUwNq1rfedLoRiRHJ3GgGSkPCPZ3EXthcPZQC8Zsv5MfCMuAQrISxeN7Bf
ZlYXI+poineuppIylhTAKhUMvwrc4EZ7qVSsi2VmLPcUXl9tM39tTpFHhx/b
axupVPcHNcxOYdlZ5mT+FedPFVixuZmclcUMkw8isb4OdNAUacRIfYChU0iD
/vEPyUusptNvnLNeQ3UdKv8ZMsqolADZ9NplJuHwICpjm62AbyO0sFLxMTsh
EUtexmqXAvomg88taTGlmmYIoSotGFk/JkQtRSvfYhBOaGxqipDJk37TXMGo
ito4MBO+bYUOqFlOZbhETgzAoen6a2kKoclxveoM59/VA7Fae6YyRtdrecwr
CAqZGEQQtSoDvOSIrl5/rrYLvV1x2CpzcXRvyOg6Pwf/BuVhcPTW9XBGIzPx
6IVoYeBiBWhv5C5+DXA7vErmXVpijzEV7xET/aG+ld7uyCK1jB8xmYXXVPwD
wEA2HL5CEcEEsg+5ecoCdUrclPkbaBESpW4gndVpmc2TSYkEiDMnICl/IdQo
FvNzKew64W6kPrMuRNyCuuf9SZc5obeXtGXmCdgqwVdaltuVnud8bjFuVf3o
cVTSQYeC2a9KUw92VCReHEAegSwhRbrDe8rRGLCquWMPXIsUIwdQIjX0PMhE
LeiHTpz4MAYOhZjWjnsw6GgdkNV01Nror32OY6v3p2Z19ugKmT7RSMgV6NpK
g1HvHzmRN77cO7BhVamZBZEEJFiY9vfNimJUfwPakX1LkNOHOPP+F2LLA5NJ
pnsaepqVQzMKr5RodL2ShesVynsFksgfwFtPEuhXPBfgHum4YR+zlwf0+7Rh
EAHnpqF1jtkEKgawjWfmRbdvQe3fFCmumHMtcW+2FucNsfNmsNPoIKFLYPsA
NBkTa+gBxOfcqp8fclPB/rPVuC1nf0iEs9WkhkR4l7SFttgw45cd+4d1BPnQ
IjjepcTmtIUtBPbu4BpR3/Fv435pugVZLWN9Fj91vJBhgJS8NijBMNLnIOR4
3b4yjZrmsgxkTenu97XgYnf0mOzOwsM0SzkRAw5Di34MCkat9XETvFK3sM0p
e+egbaq9dKY/tzP20gjfudY/cC/kUNd6X50b/8a+ssew4TwnT4eJ60hBOIWF
L1Sgswj1BNTnFv6boBuc/R567R5X8rC1Di16mrRpw+XjtJuxRN+At4XeluEj
LZ/yT+C+hOohNzjr9qJ0rmqA8bcAKJ8xFMx8Vv4AL/gJ+SJTeGHNQ9rfNUBF
j50QAbfyuq2ixU6kJlkVW4zOJhs5oaeA+wJNimeuo82yG+Ayz/CBCclGAe8C
qLiVilyGcj9jjeP5aIiWjnioPda9HSrNNbYUXEl2AI9SSU4oXskwjGk8ENyW
x66O2W4y2Nt5duIJN+4q30BpHcrkkRiM1SHyawNtt7TBi+z6vp7HsSKDTYr4
M5I1rOKkPFwZjgmn0ig6MarYkSZmQ0fynvt5wFXzeFUm6Ex4cR0u+006V8nP
OQWoM1J3KOyhLc/zji2+Z8ARt3sFPeuPUDCRFwKlfYP2HpckQbNvyeHaKvT7
QXJfKRjd+DHPWoZNb8pJZzKUD+Qjly2uQu5KD1RezN0UdQpy2oCyDpajRIGh
YkaozISxXJ9Pzjjh5Mi0wlGz8t423JLORUfMS/H5N4GiaCKbW0LjXWlYJjT/
IgSO/RfQkkEYcobPOofKzbyi0n+EZEKOzG7D0Tb4ULnNivBJl5vUYStbN99p
bgUv2KJkbFXnPG+fKadDe+ZJGMfoPrKiPMJN+gTR4oQcr8nFqo4GKuziSaOu
MirwHDtIV3Nj8rb0MibwJ/7pwruW2dv2855wKEAfmADuUrTZDR9FQLz0uIbL
5lWaoJJI/ei5xQpAL9VZhI0rlRP8Q1OUi6wvdnqCZeClJPOCMcNT4AzROFIa
Kidv8b89QYmJYkzOJ78WiOFVmG6cSz/Mz4HJFvc+LF+FIY5xoeLbp9A7X1gO
dVYj7rHhTbXsUckY9wkxBdNqwXTOhoigoLHo39XXX3zBiIllgW6aJLeDod4p
N3xcbFb5wXcbQuGuEjFfOOEMiS2QwUvwrVHkbVAOBdFdS2gfKYIEXdPmH+pp
xqD1eXDvUBxMMAI0yqW88hPbOVy+neDt2RpPcNmmBaToXqKoVBzicwUIVfg7
vmr+CIgykP9+45HZVWmf4OzaXGDg0T9oeC9KuDjKtj+RxKIXE/9llJ+kGgwA
JTpvor+Y7ri5B7zLDKxkLPyJs07KnC2zJNZcd2Gm78gXJuOLujJPq3t3ldio
AJCfreFouIeo+apZcJbXCfKJa9MUvX31egWVd2PXEwAqKbzMrGO/bSAJZAsQ
q9u58cmXPajHpVnMTyNkbC3Q4tAFGb+Qq0HBwyE88QLDa+PKH2kEmsi1ch7r
QKWCAnBKqbJ1vQ+HKoEHrifkyHlrFv4ozDGzKh1a/MhyBor9VmDkVYuxP65l
hdDudGoYZoDDLTwmfh3FsQpnGAnn78KPNDxCSc6mZ/XKy1ZdHpuNwyNU+4GB
XVCyYAKmYTb8Hc7sSzBhfPV++M6e8uCL2fwdV1aO+h2momZM7wCTBGZ4kTsz
9XaiJucPfMLyl8S2/PN4oS4rAl4Z8XZ1zcRnwa7/7YQPJgy6ElPZqFoPYGdD
DDLWyl2Wd5knRyXnCIB2xpcEqQOVkCQ+MLJFWgQueVt0Hn2RjM1CzKB7DCoX
rQhWSKeqBd+56zJiokBJDKzHdiien4BAIuzGgbe1asAgbd5DFtp8Zi0pK9N3
0t89AsnIcirg+KCexBpH04SEzF0JdTYaxpd4OjVmDvy5U8wVwr0z9xvBYkR8
5zxLCKjnIuobj0cFizA0c/Uqq1rjYPsg80w3P3ZnN3uCnZS8WnYdI2E+SHhI
jIG8ithQn/NCjXiklHp/zDyJsSdPYETi2T8PItAuY6pHTsqpLmyTdHiloB2X
MJwt8eF3qfg1qxJ9GOHxRz6y4GeYKxqKze2HQrDo0MKX4Bmqes/pShHKOTj9
QR0R65F0QFOFQ+dIXIyfqbzcKdP6mubCswZQOWxk9GkGXuw7aLSCeP84MYSt
o/Q2TOX4oi+mdmqitqRR9JprNQZrQHQq5k6AG98Wrssz82LhtAnnryLlKcA0
pwh1bBJiwldoAsCJbeX4uAqd2Wl8gA9ad2YY2dAham14/rZo34LcEO33zVP2
IzPjWDAYYa2LOw9ETcnl30qjURcQuI0NBnYsYH5mF/rlRAx/KtMR8ZwFucBU
u/E92SxkTvR2Yn7PEZ83ehq4oJmsLUdVFqgokrh7j9JRiXBgxjMDQ6Otcadc
KsIUVbpT15ZEs9Q68YEKfgPrqPH8dAUB5qN7w+rd7MRyyNY/YKiRZXzHNMFm
Itp3qJma5mnJdASmnq2WUP+unqXr3hzEa9wOMgZBNYA8XtHLLJwupnyFTs3H
6gPbzWBYfTygjTZML2C9GhWdvpefOs6NYEgQUTemV4ZnUncjNG/hZISR+NsS
Xqr/Bn/8Rj3braX144v5+1Z90SCBy9G18Fk1KyINcOMMjOpGd73W9KEDERCX
iKUxUSDmALmdwiSLK0ibPBep7vKHYyRtNsO7xIqoA77cHoKKk7tYFk2ejeMU
0DOY/S3j4lGrC53xhk4bES8ylpHRaWR5181KYvdf8d2EDnIB5SO515Y2HUbX
LAZjx1WpQy0pK6GBf7jpx8+SXhG3NHJMJETqSt2T0kHH+OUNqRZxrjNXFueu
7YDIp68e96yN7hvSqztuOOSs+iEc/c+xjKykvavSv8InX7wo/cP8NNUvsuXJ
uO4hG9e36/HE/2fxLwNZuGaMH7IK7qBgwkAPa5UxpjK6M9npXVvWgZnNLsHt
xAyvUAq/eV4BcQz9ao3dwGb0jbPj00fjfcJ0vMQZiCJxm3G7V3HKjrJp0h+4
KZJhV9UhXaxW5yszBBR3dDo9ceh6Q7u05ag6VqXN3yHTG5g8gTyrSk+2sx8h
VYIZzZQCGL/H74r2gNhpmd/Dg0eiBKVEucU3ppNIEQEYb0H/BiRJya/5paHz
WQDj8nxzjhF2YfytegJR6xFtu7Qmw74HgtY4dcCeDkcKEz9Ho283Rp4++a+S
O0oS9sXITUAvAr00SJ2Of9TbMG5HrfUe54DgjV8K/qaaB4cUt9hah4Zl79JB
mWqBCBkS043/boXVsi4W9AFCU7vC+yIoJcS8ZnnO4DQi3uEG8mVlOQ+/AucF
63YV5sDJBIEAgAtlqIZqsTeWKZNT6e+cbx8DkqGEuNhXu1iZ+q/MwPFXbGab
nfUdqoa+RlTKC8G5CaCSIM8Fg9CldSif81FOPyP3cDjF/fOLaCVE+ilx7O/J
JodwP2KCmZnhm6UvNam9d6obOeHBYKM+mlAyPhkujk3AVwVm0leJdPo3vTz2
PrCIs8H3NnioUg1Cd06x5LH716Rj4TPAiUgXjsDwPxpc5ch/45saApsdl29B
elT9pBQAyek/+6r5xhWoF2riRiBjZF97XN2pwQgt2s3nzQbvNhMbpoe7/wVC
WgXNCEQF8C8BnsWRw18g1CilAlSd4Bup+VFv5f8XTkobsLahBaXRPbbTYe7l
SlvAYrvJHvVPvAzBZ0h//w72VDhuJ0C+vlg0jXeNOEQrFMs8dX25PXrOcJX6
sXImxdv9Z68c5KEA/VWwSfDj62OP4Ab6jXCFEAFSDVx6B/q7Ard3He+bbDUf
Rnytnbn1s5D/eBuzS1xNSeB1T/GoiL3YahYf5vN7Vv3NdiJ09TxtO8e38nb3
uodll484f+GwN7fiG75s8xiV3Ve1UIt2+BGzGZxUoYfzSt9zjTn81n1vn90j
MDJy73GGuhegGp1aQF3Nt2nmfMVm9qO8gVkZW7S9+QS6owExLE+OhlaCIv+X
COP/69vxzK6Bo1nzkIYed8MalimwL4Z8q40tLe774QP9b23rQxl14o67svOr
1e7ZZ5eje3rozCo8aQogarGne5qmKmVfFzDIoWOPsclCQhfSbmhYFfemLzXu
HiUe4yf4KoHoC7AgHmGCcFT41qxZsogKRvKlbVZPmURWjCb0jHZ3iQLyWIVG
2BNVTlMUgWsYAaRNT5Csp+ixJTwaoCSAh6qJkjLyXXBlQB/YNEYp/LaG567I
L1FnQRv5pyOQvjaJlZljIsqSwViKlm9qFrqxHCXEEox6frApYngKQBgQJt0U
yFGgJWcoHL0nVC9+lTmGBZaX+RgBl9582Us+o9eJTFNhDtUrN7ZxFnb43xPO
+8TbdaAwaJ4XneGC1yOpu2iZstZxQcp/Iw6vaN3K4z3NAe7aQZZTB9vPo0h7
QgyHom7ZrKBgMHVTLhWs+exq6JBmZSGwZhuPA2V5EHe1U3V6UUq1qVY0Qe5U
AYqezpShnd4zg++EwhiRxsfOXOqaWfZEn2+EpL2oDvd9X4qtTeGPYempLytQ
71sDqWqjKP0OxGybwjDTuoByax2FMRGECHoOnz1KV+6Xg+qaukP/iNQ7yxP2
B5FJomXyp5SEl+so6ws8BDK4p57TozqEVx65desdRtCcOW2O9evbYmSwAiGZ
MypJolLbq+g9GXskRDAITb2N5cNe2/LvFHxGBDhYQUHTAGCgGThOeWVSgxSV
t4LubgOW2fFrXdF/fnbHOL/9cJNj/Tl2DRB624+PE0Hr624jS571a3x0Tk2c
4RFuIDIwydkvK0bIdIW7SzztC+UoS2RqShjdR91Oy40Gmxqdz+/KxeRcLuUz
gjluR2wGW3759qsI3DzcQiIvAP8aOW8d1smd8e7vLvhbMXt0ab9/7CrKGGd8
KEiJwVXu+1lsR5nM/8iFTkd+xl+kDkz/C50G2uPnu1j+qGm465vSswmbMBS8
zL5CqSkxXdMuymO//emd+gx29Y8wO/StXouUX6U03MXNI3rR/AvXNoOWg2pG
AiEsFYRjbT2fV2CMrtkbr4wS1ABs/apRzc3h9AW5ELiO7F+Hclu9lCiEpwLj
hEt4cYoKknwQGe3Fh+p2wOeDd5fxyrkG3ZIFokdlnzp3N5EMtNra/9uq1rme
v6cRAHOAXnlfy08lTqiZuSzHm0Hf12gg1bPaRJ2O5vTkvzpASddnxel41+be
sJ9leaHCP+TM/PCMnxMceeFa3X3+ViKcovHJuWRqLvPPCg676HXpM+HIeeY3
GjquYgbFELffwIrwZ8LqNot+1axW3CE7fXSJ29h9tRvg7tp05M5CNuU1dcxa
U+qw9s1W0E4CeNctIwDzh8h3RL+1ftlWNK2RtrMrUD/IUN1q5LrzeylueBWm
r6qnLW7Hxc7VILAoLDfsPx+uLZ1l2kS7cQfnsZ5xdTWSz/c70vp4a7teguSa
nIAeYrNB6jIXcCJwmaA7g8WzcN0CVlweQn2+YOWwXwYFoJA6jzg0PDfmEMFd
r6fMjln6yeJx9xkulHTNsWz3xcm2POt6cJXQluedR6kF+v8egjbKyaGKr4YE
UyVjXBgSXx+U98+w170QFscKi+X30P2BwwwZjc5Gpc8P18PBqELSOymwy/fv
UIXOfBRM6n4xW/LV44zZHsbuqnldOpyW251pwFjaJlTHf2msfmH106z49PYt
CeGCfmE369UtPQZ4UMhglBx89qhTeoIxlgx66JK9bjIDXDwDU/XTrhFaGtH9
KgU1TQZ3KrCpJR7zyyJ032nKGr0EBeTGi6TLK+42VY0gsL86j6jIqrB6fmLf
A8cZDswz2KbqLUryiM8dHp33lzpZCE4vCz5ca0kcio9GCf586+AvW/SH3r7n
LXt2jH0dtVAgzuNJarVek16+aA45vZoViqnSRBQdTwzaRwMPnA+z4MgskKy+
WYNX6/SSPvc0qt0e5Wy0QnzAyyfKa87PnkGOyAuf+WEQ5TeaZz4KvAAXc1zL
FGbb3zbZFpcPFY5nk81V3TeXlmu8emyO54p5JHxExhUAGqhWZ0fb5hi8G/k1
mqhycv1FYDLdkZ0gBD2NIma8m5ZfNMrafTQdQF/FbloMtnF8Q2LGYos9u4T2
xOVRL0FyB2+WCopPBn38BT95BYAxrTHOzCRf+jr9KAB4RTK7YsSR3YdmBD8c
I8lSJCNvZDMe4XQCHTgyUbzQhBiF5CZgoICmyw1VVyRS2uVzC/ivnIKOf+Ds
Sd+rlsCqQk8Wj3PXTGltvFr0I5iBSRARoocHodIumhKlkKkaB7KHHJ/Prh/E
ckHGxyBHOp4PwHWuo0LxJONit/nSpO4DzSUFdlW1UuQd/NBBFJK2XfanwZa+
AD5n1oUlf/3GEHG6dmvlvIzp2MmjLuMgmV3Ut2IxYfwoE49lsT2gFcbTFEKe
W/J+lCCpLBYX0SMYDu2Hq0xq42jcGyEQ6QN3g+0JMTOC2yoWnbQBRPvhA6FS
ZMvsoCo2ck4HLup0jikLCxwwRwMX4xjDv5jsqa/q711nXByvHQcXgmHb0IP9
eWFyESXw6kDIx2dw7Vu13Cf+HRd0k75Eg+HeRsfhOlzWz+4c1kzjA6hRWrpK
+WJacLU7lsJrWNtLN7zRXmxiBuwXCz9QLqLw5gVah/VMycKZrXcqOVlQJjZB
x3SwPdYnMi0P/z9j3cD1/G8cd8dRoeVeURnlV+RUe15vmzWM3QuqTqYEUHeU
CQ4V58/sPPbxjXWiPl9fUh4l2/NKFTra9hPQSn1EHGtxlFUihb1595PLpyz1
pkd7vi/KgEnx17iDs8N7Q+ZcH2Ql3q+IieHcWqa8QDRadFO7PorkOOrGWStl
OnnYpz0SmmL2wEWd3iZax6j7mJTwA+orG8crEovqMmMSFS8ExeGw/LpYuAP8
Qj/7CUvdN8kKhARhvN2LH6vbMaknRP8+E63yU/CFEmTFBXD/DRnLJTWSIW16
EZlfhL8zgid40Je7NfDBqBt4/Odfnxfe9aICmXfGwI/2Dk8hLXgLZoJRv5og
WYLP5wGRB6/Eey4cN9NDXeYp5DsK7y+r2dVTSR+kf1YpLQgP2EeSs3xnh6B2
72s1BdL0O1Njv3LmwDDZrxXCa+VnF6eJMXpYX/9M8JhVTpgWR9U6zimTuv8p
StQYKKk9nyt1rKOV7Nxp8a4LeQcVkx9dblqUYx1kp9p+9yXVE17HkIpuCsoF
Ok86nUjuffXdjYndalDyTRWyCQrgiXw/mU0Q0MArXQ5pwRadizGeoC0edQvo
4hVOQ3WAPM4xLy0JTxAma8yJFubaD8zqskNCkDI+GpioP3aJXKBXIszvSWb5
dqs33Ic8v1bdPmi3u9FFSI9ZKkqNKwFOWea4lCPRJM3AcwFSNH6Zz5ltvbgg
w5NvIciPIgzt23ShiTB05sWaC/J0UoIoA8+l6RTITcBWriTZNhx/0RR7I16h
w+obBO5KRLlJS802o88o2+MM4Q38My/4/A4Zj9kpA9Vx4+HqFADaguqF1zNT
dQP2crI1G96bcmfBG+ZkLICiATHaeO92sRvNTuO1ADZMdQeEdhJI+9lV1qi3
aNtItMYZ7EMQHD57Y9iHWJwalqxIcM8x9SL+tFIj1+aj7nzq825ha4UXUQ8s
IxS3SL2AnsI17wdaSowZmuqFmdL+AqvfB2JxVf96G8AyiSmJU27ymCVQzdJ8
kLpR1aZetIGjzKh+8+OoTD7XeULIXJ0XnPs4eEmhaAt8UupFF8RZtLwWjmN6
YjXhsQ4OyvQwZ10PUQOHtjVVmP1z7Yd1NmvZIG1ub94elICPgUhy5Xg5FLBQ
w0oidnmjKXvfrbn9MDPx0RveRCWJArck0OevhRx7bdiC74bNTEy/RJgD+xNP
aaqQXX7w//YKvsYx1kbCpPVZoH2z/IEcH52BpXlWn8IDKPKGQO4UtpQcVhgj
XIK3IDR4vyPftsRxyfkO/Q3aV/bRt7E+M3a/IGQ+Wf9GiU6FIfAXJ9UASjt1
CtHHg2pluCjIArGclGeymg0sAuvGc6Opy9gyPd5h/9lZVQT+OqR5DGiapfjl
wMARuPDA978hMBYboiU4U/QmLpgqlXfHp4SItDbqEUYeQ1T9GTVbVk+5/ZjJ
rh/xEWJ56ebhRipKZr+15iplT9ArrkG05gCRs454BPbPCRQjfQEcCQ/a7Pmu
ceTzpjPb+5wJgHkYtVWHcg6VL9e+a3nwG1+mgEpwL4YHefG5Br2ch6OoCxgs
Dou8q/4dwXl4OI93PpHU6lnGp1vh7C09wilrq5+zER6PFyrgf2nqraziSJca
huHUidrh5niyjlxS3Bk29Mox1+4JR+L3sTigeRmJQuEk4EkPuEcYRNpL0K3G
HyRlk8kSF4PiMU7VJpMFvfWGT5o2/FUIVKWYUyWCi9bZGjkzVsuKrzyEDOM0
nX8xC9xQhXlw4nQ4bLsbF3szaS3ITpCHMFfmVnVbj2uHzeiSxurOXhRfvVIc
LeRp1KaEXASbfcZjpF1XXWFIeAVMzs84imgbBl9koP/UWoXRwdB4eE453ahI
b8MWZs2JTP1xnfMCf3ThDZHv8gSqVjsHCbrbpqdGCPfGKM4oIYtoZkVyPUIc
cA4xfpMCMUKdp8F/7vrQy5/lL2iHvg3K7/tVfAO6OwWLvo4CofC1yn9ArYz1
jzk0VwNzabeNSMso3Ae0ZHZprzqNdeu5Jp4vvzQteW0vKfc8oTLWBsKYR0KT
xgDVRYfqCaZF+UgmpC5xElTtxpbzf3HP56n1aeE7TPkEn2E6vra7/dhzRqd2
OIZawSbmCRBjcFhfR7YvrRgP5R9nV3ZX4fIVVv1d3mJVc0XV3U14e/c0Qvib
Mbb1rE+enXTNlnuipdKYTC44d+LxeCE+9cJ2tfMz63fF+dnrnPxWjVSzMLsd
6H2kAdPHkdfW9ynkveab6/TcKC8g7h2DoySDBp1xS40VDP81vpRpq3Svp2dh
p2qraSGxYUbKxkzWOjCkTR0wX7aoNvpGMTr6XJkzcIMaBVS/2Ge4QIu0Fwvv
BDc5QzVpBtmmGQGZCZxoQm0okpFYC5rUcT/RchSJxuJCX8T8hyLzIPfLjkXF
rFyPgVV4Yncy3FaeDlVvnEzkcWVgeUjELMwPVUVnKCuAcuG325HaEd/0Ik/u
l4/BIetcOQKLu80NQ4Hr70hdqQ+LVsZTL4OxKagGpxKqLg5k5G/17dXNeK91
5Eu9arDCLhoRaHnxZUugB7xJCX52T89TJsThdR0N3g/m0nnwRAwSAT3Qxfib
S/hQ5QoGiYebQ89j5SN4/owjrBvcOXLxwZRT7t5aMAPhJHC/IYNMuuy2/IV6
tBnAI2rzzpWmHI/wRpOTrogJN48EutFcZxtOSop3dXO9/qN+tSipCzR79sDZ
FQCtBM8oM7VNuZKGrBq6bmA/pYYE6vlNRhhD3R/KJf/Y/YJjmsdAtsBqMhHG
sFpbIZ02FxIugp4rJSjoNKjIFPh84PluDRFbPY5eeBDOcFm6SSsgewts3HKz
6As0BTLuCIxIS6w7wwVEF2nMeDTwUTUt+wWiJikWaez1X8qwM1nUC4QsNm0s
GfQxW6EIYNDX0hiMDc4Anps90WN0a1D0eSotDTY0l+cYLOlc1ou7ASifATF4
M90usken1oRy+Bq6Kp0H7viGYiy72t73pZckuDuQGSt00eS9kMHZKlKoSEuf
B6KtJxa3fKb4vk+zyVzq4Siz0x+anfJWXHwtA9JR6ezahHFIux9rs34/dSnB
Scd427zmXs7zpL6IpSPjNBko2IHFPhdfY896hwaNF9pEqKn88t1rgSfhAIDE
yKYyQx8AwAaGbdpBDB25Ukaknm/RW3QY6rXMTi5hBdy75Kr0vUhfuynYxr0L
qdtung7dFeMjp9zVm9vVP9Nt3hJl2QHJ3i4/uHZ/edty7IFYW7oYYDuvlqF3
9lqW+B9WRdUPorHxll/nidLw3YDM6bzAHYA6146EarNxI2VZWaMMNQGJwx0p
0GICS7WqX53owa63BEP0wQaTkIjImEl0vkK6QjNZbpshMXNGt2P4wzPPIefk
YOs8Sxq51+dxAsOB4xIf8aosUy7KWqdoIIHJUks/UKCNugTghe80bZ9ZdpJZ
jtS+YVAYvCiZj8Xt5P1vCOJWRjV3i0urq75rXOQDv4xLWTpDk3f71JIaG3u1
McEPOGYJb39W6aqqAjSFGKMtujeThx3XuiidZ1FDwV4QCldQm0WwZs2zAq8G
S0+PDvkGEPEhD3DX7gUI3LxQS341Sdk7sLfEFNIWloMtX57zPvtnVq34JkWt
EtcyjH+R+3Zo+EhERrpeES3f5Q1vGLNZNQ81Xh+c93+bGGKcLzJFw7LSq4QC
IliwsM5YjdczXYbvih6Wkm/Itlp7kgO+aRJaw3Td7SEGaq9PHXBBP5esALfy
fSDyKj4sOfrsdEM20WVI7WU9OmdIIsoZCo2YEu/XlCC+1Dqw/Y0sMxld18uq
Kdc7uaJweLS4ck4tkNgc9RkGx8Zp3mbLt+DV0R7Gwb4ny/fWEjZ9hQVgYswL
YKn+WszCTljBWP/mI2GGJmuwVaFWyt47ALNPycl1cqSzC43CbsaKdBgbfajH
bNZJpMnUGDRKnRlt2AI82oH7wuJztEapyBx/IwBNHQTQXYrRz5z2BiKGaaDa
1UY6gcwJya1d+hU/5uWcsjPPPnHRjXWgi7HOcpqF1qvkNg+pj0okgBoLo06q
rS6gj2tthCkJTMCNKeDnnqyQdrVlvW9pQrqfPjtBcd/KShOPMkb2KImTESBB
P37A8uRXlqi7KXvRVV3S/cT3Zq/ML2eZCYj1YbP1+COtWLebAqUT7GYrSIt/
kOAPw25oYkpL6uC+v7LjZlMiw7BPO4UZVpQCztfVIqPGDyNjkISryTdi7ukR
bpxpzSrV3yavTdL3UU7w/jFJMHOyVsYUtUXgNIOYAmYLxfJBpMnBebE866lG
dSPO+jbmTcM33Re2UA5VXv8iZ7W8X3BOaAUoNW+W+9E8FPZZDICkPYJTSYN4
S77y+PUhZfwSHGr4aUFEeVOPVU5DR55mGQATyDXmcQ+3+fTxkQujxUN9ynY8
Ewg70gI7ZgzfnGgjhe6Y6yici8IZGIg+IFhxE7hdlLRnqZaf1RF0Lp7AMBoF
dJiKj2pS/QbTcyWDREfnfsR+uwwhaaVp6RVRcKVvXpZqk5yT1xbOCv9gH3Kr
YExQLBUpC99wz6szsztX85jUZtZJJCye7OrvjM19KUDymlqulpSHHG+polCt
kC66RNAOFemt/s0cnWSd6zSGpsXOlLrcxOaoHpoRrDzL8ZjnoR80OYnzor98
AocD21XYRsv/gKqVPo88XC7XJLDNUQRddlDsl6k4CrirhTQ4+k/uL1VaosNZ
xzylK8ff8Kt/bwdUr86zYJPB3U6+ZFiszlzxmdj/VoEI659GgvLioRoFGvav
cv5SfEth8gR4aXzLpb2JFwbj7Nbj7kP3h+3EEELLqv2eR8ZKAyc79222K+zJ
y0MaoqOYNfCqP0XPgl1i0Cj0zjliguji3XvEBOnzOy6ksaSgzcsrOIQQCsM4
ikVi4P6JbVHkL9LO4vLICKk5+LGON072QEID+xmlUDKiG+82I3NZj/fVUnfp
3h4ewRtzJjRYW305VozhUE4iWJTaTsb3pYr2sH+ZGnj7kEQNJP008sjW9YOf
IKfRTRSvf5WGSRLbmpCm3i9zmUtxnEMJlim2YiZXtJc6K6jRXB5ccdmk1Tx6
mBkCp5mMEX6TCvJ0N6PHGLa7gJE0pBTReCFX+Wr5BPYOolnjl2KmzZHHtxRj
nBq+l1GxMZd+8Ufjkgn7F5VGZdk7qjH2zXysnX2UWieOdcP/7hIjtxzgEn6K
T3LLeQUV+tYPnydGV2Y4GJusY3fx3f9NcAaeEy2AkjSezx8tRDnJK1rN9D2W
CgXhb1cs9e/q7UGvfLG+GhcJkig+6keB2FwZ2qHjiRauq8mW3Uyk/qCam+Pl
BQzhyWELtVr7RwBIcqH/U61V2+s1kJdqtNOlIcidxR0qt4FghgjSl6PQ1x42
Uz648vODV867hBdChte1EvzVYzYC38Uwah+PfphJFVUZoEMfG3++6H/6K36s
rmbjvW2lguTQcfc5P19cT+eK7e6IGMSR9i+uWjY5hiOSxe8JrJHU9kqIeD/J
X95dKSlk4dF/EH3/HgOIO62ZoSMcvVW9/7ZSl5YjrYxRl/PpJTBRzrLu3V1E
ZJoBpE/UghGVX/LjxVf+KZG1sAC62eZzR4DCFcCNpChGV6QWyx9jxWqh8+kU
6qpDSdqXJ2PfP5EzhM4EnzTD80Xtwae7JqX8cmxrmbvhk6e6TZzlWR1c6t02
pcm8AaSCefLA73+EY9qXdjYTu7vidCFIRc6Fmx0V2GeeYOP6D49nAyhhNGlR
z0mVQ1oVdVB2d1vzG65ulo8B4zXBK9kyiftC0HiYe1PI4IzrJzKQsBmbn1P7
euJRquU1S+9NfXEOYyKLl27bQscFlfn/fxpq/OStUhrno9iquv2kBMifWEYx
sYbpDeilzlx8NXl9AAVEpRGZKkGDbQj6/GhMXFKQLMD4elDLsuuOSJNl2lyR
8xhQiW97QaQWztpBeK7jT7bz4GMWPCVxOftgtCry+KUXKBIEPMLeytkeCDP/
/vYEOpF5QSXkR8v8FdO0HimqAyiLVhM1ZZu8Rq0vPP/A5RtJiPRC6baokD0R
zETke8jdyXfQXAh5lMmWiG/S+KV/+/R9QT/VPAVgRnYzKrmuvUQl9xhSSaz5
sXLL9iNCx2Z/U46tOSoOAbXGGU6HRuxYb4+457I/f6NT/da0P9MAXpgZChgh
yFGwtiaC96HQtSuwc9qIUnwKR7c6UQ8V5LRdwk3fgyKDdGjjH2w5zJXgrsgJ
MchkoHyVsMPBZ5JTFG0ZpmyHycOip9JEpioFBzDfrl761sIJAmNPBxMMHw+e
5Z7NPhYXxrg4eVFdZrCG3N1Jle18R0jfKsmbigO9thwtMk0qkCMzvnLEw/Hz
HSQ/ykfDN+k06ge62J8yuojB1h0H3kYlhW0FPIZET/617o6YVZWC5eH6Bnqr
admw6tm5mgtLE7lNS2vvDAg7RAPNSOmIgBzPg22I4LdOV00Znbfr7ANNvUN0
MKyPYhDqWNwhj689wQr3WZ0baGp64i8Qu2h2+YVwVlMeHQPWl9CnDkc0PcLk
ehvnN952CBlOUiDWAo3AmktdmcUrS94osFMncfaMeeS6JVgWKXSCU4y/gHQc
Y1NABHYRHnW7jiw4whpwb5i7cbPDtS53CMWifL/Z4lyUt0j9n8/qCeNjc+e1
f1QjBnBw+hPW8vXwTrtAAaBzTybYZzoMT2bZm2G7wkXe1z3laCMUHULSGb8t
/lIS0kw9IhPyJHyc3hufmm1s1ct4vQH5EghH88xsC4Vx7uXpkSazf7gIBc0K
1E5+L8yVRIMkqNTjI/ctpts6nIJ9byDm/K+sJvWk3qrvAGsU/Q4zp1opVSEJ
mgtdnRTHGMokkfrrsDUTuy2pTt8M5LM7qhSjQE9+jw2X69Ik13/2N49C+udZ
n5m2WBsRoShZqLCKjjHiglr8jUO2OgT1jt83rOi93HCUr2XqJya2Jftktwfp
RQwslxRAnIhEWimiEZ8f/0p/pR6LPqRMHwqA9msxllJ+Cfy4J2YbjwWPI0FC
P5FKunuGjVYpue0dLWHD/w2ReGbKBtlUK73O9NRUOn7O7UHLh2xF4yEmp2Ag
oHji+6DN+2Any3cOlEcwdSYrrLgNgTIm7GWzhe2hAyTpFjZG5hDzzrAUnYWa
kVrNu2OmPKyb5yHSriIOP2LBB6Eym5OZZ13wllZhCGBmO60FYz6lT50RPBdD
oIDrhBkbFkI1mB+/B+U1eWsn+UDT5ViA1+J0zxYmrImYTvPHKrWX1LPmirVk
gl4EmZ/klOEHUY9SPPRYVOCAHv1g++KJmdo5tXgazm5yvIdc8h7aSxYbwull
kjr3mR+wGdYqQpw1xvp74IIf23DSSl4F2O2W854FoK9jNma0dtHVpD5ucbwO
XdX/DKTcyg6dkWjZBULKrAgVdI2KsxWEMzRDeFlkhInLcnDaXeJiqz95H1B/
COA6QvSTfSW7M0ijOTOQvHChUxA6ajSbO/BjIRWHYG7HNeu+1+yKHKAbtmiQ
Z6qXF783n8OkS07kQaEwb9UeKxkyaRUzo7ArPkh7oChnsocawPTQn1es1D+3
01+oGAoAMoQax7GTTXiIbamUuQMqHv9WGqlp3/jC0Yn1r55H9QTb0eNCYCJ6
j4D3JzotIXPMxno7A+NO2gAklx2Fvn8448B2480QNEb72Ufrot3BO+qU0nbw
5mmSBNpR9A9vgYhq1Jb15j6qX9nkekDkh/T4e4xKJhqgkzmpwsS6XW0cxd1d
1JV+BZylHpHQxIf5Vfsoj1Z8T0uhlFFW9F5MuYJT/T0eM/maPuQGvMbjrHLW
4eHezDp2vR+PmN86eWiXpV/l2EKyCg/7mIccmb0wIPRGKijo3k58u9MOwDds
e8KWzJdBK5KeFjXzRb3ObTD1i3VL7y/YdYBFCrqM+xisy52tz6ft/eq/BKk1
7kk6P6HIzdFksFyaCO5NMwndsuH7ACJvN1opDQfKsxOBcZQVj6Vf1ItL7RqT
Hk8VRbMFHn++pNThWxe7v3kMUuYVhdjrq2VL1R6GcIaDWn+Anu4cehXLhH/y
cQd4Wp6J4eB282v9sI7QkSCL8FRMPYR+Flnk6zkx2WAnLe4ysdbVCvqp6hVu
dgFpEPHozpwV7BItpIeHK+tSCPz95FM2PTIodDMZsgpeoJn1J5DJMCjD8Wdz
Ln5xmiBAWHWP99AJKgG4NmI4QhZmO90K6zy1cKudgE06WnoQ9pAVUxiM0THa
e+r1+oQ0ImaWBZbzztSrZVTfiPa7w4t6IwAYdwhZ6+7MI8umeqeuYDiN0sni
2iAkT9mSBWufGmVn8SVbEDS898P2Pi3QWhzJX8Gf0G1UAqPxuiw7wGKfgQgI
gA4SA7CBGAHLLIY1rfnBJG9lgBqFSi0ayvadXJhxRR+4oXNVY0mY40uxLNvw
rC18zlMvcPRNEqbkUAN6qf6HzR0fs43JZN2ALEDO+KrRwLNjsuvM5S/sNkYz
7mw92mm/8Zw7xul5cKw12Ja/z9IKuwcMqCdHRQ04a7O+UM99nKO1ko3VOmSD
rGY5H0YVdKbi4Hn9+sQWVLaFKLmNJOvxGyjeo6tlDaQanJQNmAIp9b+V07Vo
VTMyoiOeFA9SuNs7X5umNbVFmX3ViAQQte2vYnL0H9+QbBvNyLcyAI1aTNpC
4qdC4V6qGb98r8tNI3CRNgQJ08vww30XZwdwGd162artQtLjSVAQdVmZ6KEx
Kdh/CXwTwyAZscR/d+mjSQdqkUU6nSRVozc370ASr0JrZ+nSA0eEwj8uEfgg
jB94JmYU/8m0utCDN2qeRJbQHz84nhJ0RMDv6+CtMk+SDxaY5Xt7YMOPwClU
jYkuCwqdpokQ6a9dQ38fbNpsaO/9P1EWJ9LMxf8oFFewQNlKQuVsBTe3nfIo
sNY5y7ZtKewTuvQWB/ftPuv1WOTnX90yOaOgPbvsuEPnt4436RsKQfFJ6tUq
FUS9FVwHnpOcLryQDlhchAHSoJ4lOqtom5DqMGRxvQLnnDgKZa9v1TR4UaD4
C6XQYgxXcq6ts5+qkEpiAngJteXNoFrXdLdKvwa2zpvoSifen5UuY3LFipJ2
TtzsEFZ81VFftpH0TOwrWt3Mi5FcQIS6J8uVZQKE+Ww/9HnEDWQns8rK3hD1
pf8u2SqTAwn62+Y0Uy/iwraJUuALfcrubC1rVxOmUZpx7S0mZV5DJmmH9eFX
p+HfMR6EOcMa2OCpVTr72klp41ZYN9ZdeOba3wZk7Pa6dAdSeTpkOPt3VYVh
2MAxSNHKSkUCELKYGCTuDmMlPZkkscCcP8GNCU7kmD9YFYaj+ztTrsA62OPw
1Qnmq0aEb/3c+eniSWjfF68QnCpPpjjPbSMqIVxKiD8lOAweykU9od61P7dx
jV+W//xCfoliYlt/Or3nfyVBnmzdNsiy49QVK3+22ACX6qPGawqkQ2ONMk3X
TK0vejhC85gPnKOY/DYPeiQYPMnzgA+EXk56p1o4YYoFmtQ9KJJMWix7KLei
/0JEU2XS5kwDS5ObZ6a32beRdGYgt74gf1Rlx4ArqUwrz+mtoesw02tXURbh
sQXh5h1GsNSrXRfgJWWXK+35m67V6QrKsZ91df6Qa3fjSdlPelhCTkoJ4QCd
21ev4eA2Nem2U24jYtgU6AbRpqWhoB2lfifWQ6/Tq/xYx2MjLWTOaNFtjlUs
bSanIITngKqjun1KMmjInvGxvL0VEgtzID7VH4Nl9QnkuJf0yMSwsccI3WWB
LmxdvUsAe6eAOm4i/kNBqMDi/vszv+S8hpr68gLfnOFDYYtWoHeVo98cnGrA
IuZM9HJODIrDv/7uEGYT8yHHE1ZmvzSYwdRHI5URFt7d0DwfIKZ3BcXslsyL
B8TsGsX/HmS8oqKnewss28Cx3ikJw/gh6LMafuH+YyWdvwhggsPl0n2ZYtxH
WF9jRL6FUh1Gl3TciNDDr2pXvJmYjktusAh+cDtruu1bZXrKhYeo5DG4yOTM
Czc2fnX5zDQxq/0jzhKvawsn79r3G6NOACwx4FU2j4KZ1+ZnU7SDAMAdqFj2
j6L8oi3acvRhZN00/FlAp8XjdCGUTDmLm72sW/JmR13ixxKttXOEVoCOj9EX
UEur339AOsvFJphD3PoALD63wjeTjKOHFDGTMRuezj5LsyL/vc21m3NiDJzx
wPWICnFrDG52dTuowlopGjIJhKdPuP/lEoJKphar25SnKtgnjPE4RXRRSuE+
u0fFHMFxeiE7wmkLDXFcbRrdCMWJ/cqI9Pvxh8BG/3g39OGH8i5F9L02tgPd
X7noUr4Bh8OmCs75Cwi9191w4iQ/LdODYuY0dH+wsIacjfeW0+BkvnMLtRQW
HiHy3xYZ0i2CB4n39O/dLYFW2q66Xk2izakugGC9Tyr4WchiZiVNnnN9Ai0m
EwnbjLdzmSgQBBO3c9G9ML+PA9e+WYQi/Q3Rdu9O9OmXk/pDg0CwG/ohna6i
zCr0Y2E45dshN2zz20iOywIKF5XdoPh5fqF2czsTlsVv1lfQjItg5hx28u23
30C6t2IEyHBy/IKbmdlVES/CTzC4ef9xLLalI1bCKe4AI2GE57Sj/LIVHNvi
YxZMEEgMJ0gaEUV9tZLL+el1u5lCdmOQ1Qc6nw9NH+WJQTPfRKfzMn8Tnarn
DRYCVOgWJTU6/veeWivnV7hACuNrrqbsCvFImVW1MTkjA3pzr0E4k5zUOMJb
bfgRPbgoIG42ome9jixOTz1vfU8BnP8XV/WIOs6m0f9Q8z6+cYqwmKXEuACT
yLATSXztTJcZCNRpTpvSxeA401VVRkQ6vMjp3maxpE9tNJGEL7sQAk2JT59X
79syurXOE53skhiWvu3bihnHsh44SOtksBmORrknHtXFZoHl26RbcKbbVCbE
Nau5yqs15U6VOzVhs6IDiptZAZgTutX9MrNmugZd60SfeVSQvA94hUKdUnsp
YqokstmzQ9p4eoDzcdP5Y5xU2oX2kQyO1tOogNr1ldee9BaJ8KQbuHDZaCMU
3HlU+qcg8r6LYLjMOKyciaFJ39fhbUDQWZM/uMnexiJy0GmyPswOIpf9TxTv
5/2/0hXqpOj6Qeg58cuAnkMkTXmb0WXfUTZJvlOJaw5W6m5ypCCI5Bdz/H/B
rPJCE8sqZQy/a6A76+sa5sfCiC4tbBfV2auNYmL0UZsul7hmNPN3D6sFNjY0
wffaNQa47F0GURC2s1Bh+cSkgVDlUmq9lIMhWYB333+PFEk+dryry4A5SbRV
+09EYkvyGMFZSlHMy9j8S0bYJvxuJT8w+2lpboPGpHsDvrm5OVgbB4eS4tav
GLbAFE/PtTCM4BWDX7HWXB+5tcHmQKTc9N8W9cN5AOLRmmRwGUWLADxVF+tW
QYtkZuIDLmlqaMKb9dzSvW19TzzR9HdvQJZtMrSqjqNuwk0Pq2jcNs4I39bX
3ZruoDYvMGjX4UvtQkSB5LdpXTw7mja5waNP12dXtQVM8dxgZCPyT0y5ZYhM
mOw1yXcO51oSxQBVx+PCMxsCtgYVMRu6ufHE3L7slLC3caCKjtRM+TVe3eQF
gUjFgOz3Lpwakn33O4BTOUKxiwBJfsc22cqfRwscALKouVyDoC0LOtAYzjqE
soWr8RTcREn/CJTBooNU1euu3eab67GidxhQzaVuKMCrTydu/69cZZizp38a
zR4vdCODLK7V5vdeoKdbBLMz+hsvlZy/Apx5YvF+VpSgrOV7U9SbsDgUuoJe
rjzdS9uMUsLVYw+Z3ZLTpchECed/opJzrb76E4athK/NH2RTkxFCZcvIfVSL
GNJKL6DBF3Hl0uOOMeS6+9m/if5rl7PDPl20frSDr9A6MfNybip6fTJ5pF4D
JkiS0mysDNwmRTMoOXhqh0Z4HN/GEhlCi08bcriLtxhM5IHPmx18yfC7vntC
+cd49NEqFGMBx5f+7ZGE/5azJVUWvvQoYQbEoStUXXDd3cd6qvZJPuoHkoeY
v8SLkQkyznB1V8xBXS37CyajtPvr3lQ9aGzVp9Ylh2C3T4l0lMmUClImrGOI
hH8lW/oMurLtfrfaUaIHyNngFJ0TvjdXq/OHrEoIvpQrB4CtENdassjG3Hsi
yE1v7FOHNcp+AepjB6NR3LptYn4cMhp0XTEFcRPeMhmdCc8UFFiektvfEmOH
QWz/Y/WTZDkErZyIbzbbf5YJPGgSir2LxU/kpZmQofnXWn4FfVV6EIUv+ES5
d5rr23qxdW8nnY+QC8lBFfcvw6vx+89YeuDAn+/KThg9p+YoHvcCcTwr21ZJ
R2c6V12A12Q6ECwEJi0zdHBY0HF1NSnLBpJmgwDVS/+33o+Dq+nWu7US5AK9
FXBneGIOOqGIP+6LCcG0ekEZBk0QAMnGhWK1kxNqvDqtRH0/7dTOH/t6YVv/
7tIcBJZgOC2z21QvcoayVHAHBgPHtxJN8kpwgt+DML3TyE23zSPPmj3oYZhd
8WC8aSzEVz/5cebTVtoz557pw2Bn/fRIXEaaKuVRa6gKiK+ujEjN0C3vcIZu
2j0A3trVdzH5pK56irQeOhirSLWcFb6+uLfgIIq/OjvUY8JMUD04RGDw7aj6
ZpCBwqZa7qrqzS2RnQPXkmETBGGZibzk4ZYeAKX8KOUyHOHlzLIbwVvPAqsZ
wRv4e8TO2Z85BnE44aniZr7DQqXgg0lsRQePt27ldJXhe2xkEO2NBV0CuxmF
YT3F9j8kQnGrXoqeU7OKfUJEcmcZOia59Vek49fkmkAhuPfnyRjo+Ncd7mbC
9yAzzphDPE6jWjVzylL+RZc3+zv/HrtPr91H37yG7MrtMijkmuBKinrPmjVV
6zfsrHjS9TgEnJk0zuw7g7sjLHQrIl16o3KwRV0Jc/tmyLzy+Ne5zfXWjlFQ
XG6szK2TrDk7P/+48v0phf1NpaIjRKke/euDupeMkvOE/6ppITVJRaDaNw45
Uo80bGKw65wqgti8Sblrvz0CZLlibW4uILNf5yPI8onqFCE2PUzXn0uI2tT8
ppPDirbtSMRt9VZQ48l3E70U2Hv9mQS8HtMALJxAMUE849Ad5TJ9Y8SqZZ8V
h8zPrGA1nSnWsTUGGdGcWe2n0GiC/wUff2krFir1xgSecp80DrD2Ef9KshiW
jqsq9p71dxIBtzcnE84dpsFT/FoYD8ZOa43JkES87E15KCiuKVAc7LbLqLM9
G5pQtiFHf1awojHouq4KRouLaabb0wq5oWgkZQF3I0xpLfxOiyZC/2+Juae2
kqlypevoguvWmwGuDFi+lrh4ztMR5kv/Wa4GCX9dah7cqLWgIfSJfdUEnbcQ
7/LryHXN6AogKChlTA6+In41UPriAeyWO4IcJp0p0tmaCYxw/u4AggxNnTZB
BxCsJsqDo7Dol8ob4CVPQHzL/KI/3mWkyiFbOoxIrsVbKj4AP15e9kbcX8fo
y7ctg/Uk9RIm6FhUckZAQ6jrzDjqtBlGE36jTo7M8NWeoOYSDd4TnHTz5UUQ
WUqd+DHTdWd3sKD+nTYtajJBIctw4m2gB/aJRhKJdqU1Cs1oHxQpctT/DH72
IfP4sYcKfpkUT5TCyElWczLLQgPbkX+OBkaWkftvZHhUpZfL0MWjNr/9ovjQ
fmcAhybLGM6Azi4XpEZgtfuagf7A49NpJ2j1EbkzGyd6rXVJegXdNuNYkBIT
ZxFIJaPNwXqyVCt4U4tUnt90mgjhI9vsjKm2gxh+/RqtlfEGQ0dBrqWBFg2U
OVdHpFHOmqlO9dZ1u0x/9jjYqB1x8xuumN3YgZqAn0RHCbq67fb46xUFbzUq
e9BncWlTFIU5pTgNgAyNLtDotw+S4ou7rT/AAeXsU3edG/2MwyIQDBHKYqmA
zW4JacsmH5wuyLN7zbDYy5eNJUdr0VV9wJg0a6cHR9DZCL1ubb1v3THZHKRE
F5STipwZ97uwh6WTHwoxg7k/YYhfJPB6MvM0UZGMiY7NPhtNEl69UsRWCupf
RY8euiL2j20BpNSgzl1IJEeqBne4tvu2OL7u4yAL3DPCCVIdZyXGKILADSaD
HIhDrYO4pHIN9swYpN9qfIKcbMX5kVA7tZFv5PgZBRWkq/TNBaCnB+3temC3
ZQn2ytqZBRCb0DMjfjzRqwFZg44exZYCKmehAq9BuEysFDdiSq9LoMLCBFOm
ufr40u9oXYf/AKpkcndItoe57U3wVzC7o/Z9Sv+Apqo5nBFlIUn29pY/WgOq
C6981w/VGyAYX1IUTfz6HtDWJ4H9WgJvu/zWGYS5/U3lJaFrt/hc2jwo4Qjg
h3yOnueWkizgjP1K7CFPZ3mNSFVQSNitCyGKmBJz48R8vDlTDs+pVnE0E7pc
pNGwau7Ex2zCu5y3L2qZIRkDUJyJXgQ5yuAOqpXYTGXuZMFrmoIKcgTsKU72
DGTsSdruzrOpnJDeqqf/pwtKLVWpQwBp5B1AGjrvAIaL0z8WDG2gqyWrnXTo
gkzJb5V1R5lcXvvKI5sTjJRyS9kBqm7khrOyfeLRtL+mgQnvGJdHHzNFbofk
NP+V67YEaa1MQNBPYN3iIh11cezDc8II755CVPhYR6n3Hu0m8u5Tsqwp3voV
bZT9qALbsgaK5/BNfg5nDY5vB9KCTFuguvUAvF2P+fT2i2BoNskfEYa7woJV
9w2hiqREncF2c6fIYSpAmi9LCShza6C6vTlU7IBci2PfWIzC2gpY0l3vq4Kt
RyMcqvFK+xAujhAODAMUBU25kianwPj4F53RyZcRIkH9TJiUjSaH8L+3OLYm
Z29dfB0vnhPXowBapHsyMURBlV6JqDjtYsCpbc+zzx31cDih23ZTaSvWrfOg
jiLEWBAJ3uRHKQoZQIKgBrPWQEk+4wWgg8F7sWpwiXc1aL/xwA1GRL6PnUgl
GCjgUlFZz3eIv/fiDOrjPbmI0AY8oqLF6o7iLkz9lt+huWdR+eseSer4cx0t
o8BPeRADxobVw+AoLOgwOBKcwj71DflcjPYcW3hA6oBohAvrDD5LoBXTrGh7
lp61fZ5vJ+g83PYc7bIHaHblozw4i+xZgqUvxkVPMH4Px7isaKrntb5pLIFY
7AoARGgrxUoIPXkzYO4UoA0rM3lkONJBr3FH5MvBdqecy+YdJQYxOS7t2/H5
yRxfsRChVdLLw01jyu0fMmAue4Rryb4lUxLx7tYbgJnWRT11H9rGs7v3HdkU
RSgVZSVri8ruTP79vb+j0fXT9ADru6hin8CdqaPzpSE8yKPh0myfJoqSsxe5
yH84FF2p334x/NfPOR41pySp9YgzcoxUb6npzKkE+1e/bZ53vvu17F38MSyG
PfCxrmzNIP560qoKA3yegQcLWLE7Io0eJ0UPn6dxt4AItdymACQ6ZzwXc8xN
+gJ7aRpUQV3ShAg/ofphIN+19dHKizeIodBZcEKwmZx5W7HwupiwE/cdOT39
Aor/j8umuTX/nlRSkjMsAkBjKQw1m1qJ+bvcn5tgQatIC2bmanq0Vyr1MBL9
NgPVuFXjFpTYS5A029ew5/BFl/4YDmvZ1nnsoXld6sOYJsk6Qbj/QqR/niFc
DbJt6pvyVjFYHIaULy6binwIw/yRAE4MsTWIk2+4gy0YWmWvZCqdqmoorwBV
S6m+gWL09JAdtLeMNNIzkyodBjfgg5RGCKhzjFqWsyW+1NEh1ZXNs03cnW7R
uI1MbvThTLHNJxub5EUXiwxA1DW4BTzWt+1O8WzzNeOrMpYvoQOj2dyAOjfI
zWOyciq2SE2sHweRa8uaWMurI2GkwrCMwus7YebN1tLNHeYyDP/UDmQ/hOE2
33Ndk7XabGdwkcXccRE/BjVTAea6GSn9MMbii3lE0BnRwVV/qKOj3Wh4p5dS
7wnj52no9SxCAv8L3ilo0JS8RJqKP9Cv6ItBoz4WD/rWDZeb1RI92QfnaSm9
nH+1Mj61HvNpQHSDoJ1FbB0KgtYjteDT4M0vrqQ9Luw67l0xxylN7UzPU/Ip
Gr8pgS9/GdlPtWGwRXunEHnNhLnqWjOaX0YjsT0Cr1YTgapPrlxK9IPb/cTY
Xe30OBoM1WdGWL+1UEfb/w2USkqZzHT9HgR/s6cqB4WkS84RW6mpz+VudgT1
hLyM8cz9Gei9/5G3zQtABhc+5oE8OFboLutylS13POztji6/f725SHlmfoIM
lwVqM1YMe97LzsrfV9P1r/Z4jhC0cJzh1Z2K/57iCB6SZmY8bqOqYSxtEL3X
Njdq1BKNATcvtkvrVeAlC7a+wTQdB4O0nBIzribI2NgDMNhjkdwQC4zbifZn
SRX59ZZKIuzMnOUS9/IF51Wctz8P95KqjkIdaGwznbRyZt3fCp5ulI2umTJ0
3dalDhXEMAHVfvYSULkmHZrE/iAwm6R6Zw57obhNdJUlaO3m2ws3JHhDQCPn
Eh/VysvUvoBoOmiroZdz+IZH6NwVYNQemoxEMlSTs8Cnjwb30ioGFm1NC1/e
tUeeCK+m/vr0edKHGRT4EMAz4vOWMqnuuzNbp2csWv9nJM8Xq7+qrndx4zuo
E23Wpafhhol+c3YsdxLhP57FkOkvCHKWLY9JSRCinkcewcSm/HmgDCF5tqK7
2qZyMoUU2UKre2C4uRkpcvwn5Y7XXIGYbBgzXkxQ97S8Gw0ex7T86DAUsNAv
EosuvNdChaT6z198Vnq957VegD+xrbM4D2366ubNI4uAZSd0yVuMxdQYj8Ka
XxzZluvK2tPmdRbjJUZ8B3E9ZFDtqKJfWC2vQV4lQW2UC/74R9AMxQJPoZHG
nWXsLJl2Gr53FmUqlTKJZgsXI8qIVcI+Yz2kW/hzTwKelvGX+9IjB10z7FSI
1YvcQbHUm2klZtTPljlzPBiteDn6DPQMCULOJa1xDtCnAUOUTQoHwwV04ok5
YUuAlzXmPRx8OjqeYALFV7ltzX2DK+EW5i3eLR9sEXqKr5EW+/ZgJYCN99h9
N3I1ECr6jWFqAdcsSNjcGcOd1DJv/PXUz6mpjHq70eSF3UimEJwoRWxLb/Yd
86lgxsvlf1MC+ZdhInpVZG9hdvviSsnlzfrQ/N7oNtwTdNY4Kh2roTw4Tkuf
Y2af34zrek9Rryysfm8Ki8LAYtViB2dhCJRaLgFuekD8YloGKnYnjz8qslrd
oqFS4z4B7pdc65TTYOb20BKKUo8koiaIOuE4pOhMVrGqzbBFIPzMpNhio0+G
jPgGgVMG6LeQYLHJ/riawILNdPjU3OB1PQ6g4ezSGfgXbbFxawWOFol5GryO
gKIi0tUmnrkwvRyLtWgjRJ1k0Jp+X35JyvMbFdH8kuxK5ftntKjOgDxNPtWx
EcnRNsBSiniVH8ByvEImK/AZAzTOppSF8inctG29eMaaBp6Zry8YyH/9nt75
hvgnuaWqPWeXusMI2ASaR2nrlfnbLeeZi2gZsbat4699A7IVakrWjFq9Ghpq
WPGrnBPuOhx29D3UtkXruGpcSmdF7QTpms+y384CUfsGBrNfg7japQUIDjTV
tKz1mRrfOuF2AaXQYHqaYuQ+BtKSaz0a8QokrsnncyJ7LNFEuTf2Q5ofG0VO
O7Rtyj/C88LGu5tL+aSipOCvYtiXVBnk697ixiwCzTkuiPLkIJpMSnlhki7P
qbYb3nLKQTkDyISIoDDyp4C95XZn8xYNYYOVXMudZkZRKIT2j/8DL0PHPGrd
rkYF9UPkrqV66lGagU9g7xgBsYpG7jyVSMhz1MSZEiUZgKn6DycXvZdNA6S2
ww8DjM6AAanALLK0qasjWGbGBIKGU2RFq8nNdzsPO1coLb64J/08RPjiZVXM
vFxeh5an4W8Jy2r/IcfVQ0UQCydq7eO0Z5FxpRlozu+lu0FJo1ysQ5MEuvW6
AMmcdnetuh+DLf5HjV3h4xY5CSBvSJroD+BB3k396rdDTL+YD4ccSyVA49L5
n5OOS59fQhSIsunVV0DGjQ1qgumOOuqxvPJXl1lX6x0wejs2vCQm2sDw4nZj
CGuM2OfxErXfvh7lKXyREtyJVskT5CJWt0o8H2iDwWdaJ9Y9pm/o9GZ07ECn
I4sQGWP4553lFbyJDhVmozNxwAU8PxNuGvcyeDs7WBShmBsOqFw0kNSVmG7Q
21c96sHq2z7UyI/+a0BJezk+O+4wb9CvgO0+r0vo+rsLYVg1/FQyRZWV1Mch
7I+yNbSccL0Uj4ZLHJSjGDNYbIGag3SUOQjcvBbL52ox7/nWp+HwHRg+fcKA
l10owv1kBb49x34FDp614RzznxWjYFdMqRyXvgjYFSiqHm0EpEqXYOzd0Fgf
wSwg6SbAYZInfbO7p2goqH4txxPqShDDmU/jxmbyN4x17vIq0ltj4y48ZuYr
T6FADPnAe/D4o84gkPXhAfnM8WEL+5yKxhr6rk5qGgl3RuIB1jV6qIzlr9TT
ceONRQLh7lFOIu0LEDuCdSu1RmTXzy8F+xtiHGpYerujX693XcEXTzBecvfK
GbDn+F/Ev/btimgNTCEr1uDeH9x1gsXhKaTQV69QclRJKwkbHes/sjnR8pBo
j7tpI2smycH2I6JQYEpPPQCjTt+5bVUujFGHawpVHLyja0gLH+SM79l3s+bT
7wryS7+kmgAuilbB2IInNeL7cxiUowYVS9X0yBK5L3ix4tIG41CQWfyujdht
w4OFvRPwYs8iAjkp5kIuj/1hvli7ideMFxBwAxVYuvg1KQm04yz6MebrptGX
1xloIa+P0D9p2zFq28eCZmcS2t7MWGaoZItsgoCc5YjbBk74dcWG4MxpYAX2
nMj02oZl+pRuQW1Pze7HA7H3J8WRL7s5LlLtgZattnWDgwUO8JXYOewLbRe7
d28hOCRaZlpNOD19+MgkwH+fFeuCqq+aj84SXG8d3rMp+GuWH+IFkAB/Dblw
kM9tsmb8vA7xqHdOAw0K3NAw8Nxjcjh86GEO1DD58mZIOZ7SaxPQez07Gj+u
nB/KUUPvCYUgGkUZk7Yb6VDNNO4RBiRcZLYlOPZMs36KTEDiXd8OLu2/U20m
NXexzcds9aGyAg9EGYQqh4x68DjC24Agyo07FeBsI00xc4xpk05k914YzEEG
TcRhGSRxOBg3MP4HindiwPVjMOdQeywD0ztMH5LyCn5krCjtGD2qYVI3Bgru
iSXgn9Hje9KPlcLHNJsrJRApVRAgCQ1MQlX742G7QY0sE37XxTrtbm0d87mR
VhiP0qmfk2AZPhwMCwVq/oqfJHjRGJJwyKF6DoMGHdo2Sm0oBrYR5P+Bo/+9
KLxyh/FwrHcs8FL7uQShXRrR1MgbP9/1k8JEjMDpn/KoRESZ2yWtW/X2U19+
Qhe+kCbeEXG93yeKc+NvIDCfKpnhNzgBZFBzF4gPppg8l9isGMCWRWQskff1
P+xEdE2X9SCXsV+7i6dgq0dqozA8xa/lekW8NQ5HVVajOMY4cv9U4AXCkNCc
jSj+Nt6K+OELZvtjj16iWO9+vNNIoxRocwr0U3GOa9WlKWob9k46gdUBcgKk
0jo6bUFfGTAp/hhoX1kfftbyJueSQW/b7+4fWmtua5UEHpkhl+Sc0DZcnlJk
GB0HWeUnVh6vb18OiQuDRnHeYyTJO9y+50FB5/AKv0XcvTLHKe3OE3xbp+PT
DW0AdMh/2EzUqrfY8GH1jKGnGDSBlD72CA525OrXiTY8W6Butl7XbGZkxmV6
H2VGuVs3YUJjnV2XCdGhBHg2Ozg3HHo++dVTrvDjFn0iH7gRUf8MW+KXiljS
3vZaQsfEbnrM1btqyabWh7fqLlmzaMNcSoj2FcnmKvN8qYy63v0hNR5mfJRf
hf3hLEpEMWKVvzls4Wn9wHe/uyrBHLeLPf384cxEtbk5NZzxDeH7gswFl7ON
mfO3/YVG/bsw6CtYqYFAwmSrOXXaGoySSt7Vbp1KbU6ENb1Mv8SzZiPsDN8f
TnH9XJ/9M4wLk8wuccE7WoidLSWfiuWJZZCbgpmegm8qbb3F79Rv37BgwemX
0w5a7cGbIt5iFiunbrn0errvWW0fIvXaKtarvRM/qOWGUsZNaKB4ml8w1A0P
oxhPBgEDlkh9nKykVMZ7vcFfaAKY9OCVdQeSeEJwncIZOiaHSKSDKBVA2sK0
AhgfgvsfX+PT9FQ+AuZjausqrIJ9GkqxqGETt+Oym81avAm/mN4KDxAR/MPb
cXkdhPTfY9Yd9+C1QrRPksREkjHGV2gelrw0x1clkPeXVCTNfMntDHpTYPmS
GqRaEamaz7oIMlDsl4s/5DXDxRtm+ZUzO1s+dko66vb239J+P1yyevSqIqBP
CJ0ES5VuDlIA7GuIFWFIDlDWRg2ydzTPyGKxYgUD/7WtP3FpGAUpwzXSXLEA
FZ2uA+wozacr/mlMoQ3+agcHQuTQ9Rnpyv6g7eZYDb4xi7ddz3Ah2kRHtQsb
BxhMsoAV/d6im7mVqH+L8nvOl2XXurtc+152IByrIeM/QJZf0N62vh+nKXI4
xEM/RO9+baUW955kLQKMak0ChgXrzdNxOFloXMZftidZ3NQMftKGIvICh8ZV
EeB1g0Z3KA43IeyT1DsVjwt97KuE60zNmc+Vax1Uc92OAIFjsG03re8qCEEX
f7px6Y7UiaDZu7sPfSJ5Flg8QJuVumLlpjgOYNaevpy7NrAmKbGYr8SlZ5CU
t2agX0VPZSFaNG/nQvK2Ko452f/rBJYiBFYm0oYYVfw7Iip5AyneTktNLo60
DVtQgyfqwk8v/zCBrGKqFlM6Ter2ZTj8Sm0jlOCtpZOfJYnyzfnzfxg5BnfK
ztaZkgHJ6wvu0lCoR58OZ8Cwn2pMGA+dMveklXhYobVmDHYGqC5EuCSv/uQi
6qJquMik1qHILpfexvhh/eSeSLBaKZVgZHNZfbt/fUBLa8dDoGMDCNjahBFF
GFIWDNoYYMWaZZH8lKHTwoWtZ6DEwuKprl2IEHX3vjX7maXoGHW09Qmn0q/k
ROS/+3dRl0l84uaCIvFchoVIQka6V2SuuTQOLREtakMS2cAKD27FI/0rs7Jp
P7GCtKahfco/Lt5cJHGPDLFs1RDl1TQ/KXeUMiEK8lbs5+nBX5myJL9zsQfw
5/nV2uUENm6lQaFSgbQijxA/uurqK7p5VQzWDW1y/2vyt+J7wtY2YH0pYxGn
GHbDG20fRDwzIwQKKdgl8nGQ0HgoKzYdC1kcxAubNh19ALCVgB3FrwzbgfbT
R148FhYP9U9Y9yTRrXQoRV4/j99kNEAJpjI3UKn5AI5Oy+owBN0XsIwirSQD
vkN8SgyI8yJa5ZTSKoBgq3y+enVGRusYEsT9yzLBjuR/rLKBGsipbZ68emzP
7iWrOUYhikvWWEKkhDFELJFmMhCQc1N/mFuljySa+Ng9OJWzh9CkYZ73oDYU
tM622ID+zuIUzmpMeYpHQy+QSY1oAbq6U4iKNXjKh6BT5gSqfSZSUDHezI3D
jqFqJygrUHdqxiFfRHhqrJHDZxR4/zmd7vrHYC75RXIsr9BWm6iFIF0ksBf+
MxA+FLHrdbgxobdfoQgo6l8gMXNjWgKY7mTArVNOudD7r5WTF/EZMgtG9B+a
M9plRXR5H+jic+lEFQlUTU+9HIX9vRli/QoMWQ3PR+8fsWH1jKTSiqlKzBjB
kgr5NrckYv4MemTVcYUYYsI8ftp2Y4FbLV0cOdAr8MVVzpy1XDwo0rRs6K+q
F7qYkNAauchfNthAP1I5kl2BsMe/K7NyPZR+/JmULm+W6WspjXMzKE+x0sv5
b9xtBDOtPZwq5OqJdOnemqbGzGjIR8s1uZuQ/2QNYEneZgSursAVJYkNX1N3
piuF4FFnBd4wB4AHpJ5pkE8GRSxduSBS10mYZWOnJL2BxGEg5gYLBJAFk7zX
9gh4bWf9p38e9o5L7rPZEQI56pikNs1w4tZdKCdGItN70+t8dasVo8l8krlN
NXZmzuRFSugDfPkVPdN9pP42O54/0578WcGPAE1TJ2oOznXtjtSaBWjX0Vw9
ll5T+liRW/jRxyPmSPHydiU3BM1z26H7/7RR+uw+MK8GZTIMIXTJwlY/O3nV
xqGUiel02Wv7TCv2PMNFliXmVZSn0uDz/aYCHfdmU/YrvtkmUhU5nkf+RMGg
IWKwFTyvKUIRhZzm6VFupqrOSbFZ6ptzwravzF4eqozAP6AzJmwjjtCZvh38
qFzgHEDaCbaw2SuGrHhQawhevviKRjE2Ko2FMqlI8Z4r2Su5TTF5kF7Dr0Jk
tI00f7g8yLtevYmWcLxXVcJG2VoZiCDSoDblKK3N7b88YwZsH/n2R1vcP9Yy
Vn6bY8hOJt8jdbSWv97wBpPFbCjDkCXyVPgDdOiJRBI+cblyaP2pJ1E1HAO/
K3qLIWTgETKTIhj9gOm3fmI5rrLX/nfk/AII27QqDNKl7EhJVq3Ff49z5tgi
rvvHcXBbWJ4vpJjhmCcPQxrbuB8rThGLMS1n57TB31JxUE64PAeytrKGMETt
vbu7beemWiPpVJag5QAbc/kJBVf+rFDhllNgOKdjFFln9PyN49qFmEbrr2ZL
b1o40UHeJFiTpNyCGVBt4LR4wf/WeBL+rPOwvMCfogknorguZO+7uiykCkon
qKGccGBRcArjcegLppY4M6XgDXE+Eb3K9ePC6+9qb81R1br5od+NajZgMqI2
MeR7ahoEoNBkPN23B81he1RG99FLi+4IBkC0MZ2F6dTVwG2Kc5Jc2X1a/hey
dBuyHC4fimEXyTfqDJi2XuI7lsQ88065bLlTpQOeJHNlfNTEizoG/YvHLGBz
2Lb+WgRO8rpk0YNCi8OWpVRupl+MSX6jlEG2L9DBbKL0TJGfWC6DjEqR+KvH
4E5f91/dPAn4zBRFa4Op4muUejVlf+4n6BAwfofRjOU53B6NeTX00rsgoQyo
P686L+Z3lkHga+1zjDfnKKsAGy0cumzAUBOLKQTeeMGaW5yHDnzcmjgr8IC1
wCPP3oKsLSaXZPRUY555lS01fL2Lv8QYt10ax2jgG+h1rzC8RkA54hFxAO3L
y6SRpycMexN/xDOr8ENnp+FyaKY8BX82nPFZKeOLjHHFXBriFrL5WanU1Bty
GdlR2lHwcpnRcyHCe1fYZ11EpGoCzcctRk3B8XHtiwE1g6H9mjqjRV8LPPZr
WTOr5pV4Rxz1g3hKVZwayvCLN1Nd+JrfeqUhD+sVyq4bBKBwfkkDTxScyiNQ
jyXICxdyuc4OBhWbjz2yNRZyicm/JyuVJ5M1FDAiNR7nlfYWaTXtErcCLA5b
nWk8QE2rZ99KVxFozKzHWQ/ORtKLNUwI2RDRf/+1plHTSbyWTTpe4rVyATjT
hRAtXxWoquQN2crLgS0+iBv9vqJ18D0J53XpUKhY81VGfJaUs/5O/mviSZRm
S6eNX82pra9lyJlfhfR0u20Or4q1vZxo/gCcpNPSmi8fDalaN3jlmR5IH/Fo
bPIIiTlxdDUJCu29KeuPBnB058xuNfy8nk1VJKgxPHUc9w4Qj1vqSwaqXRVS
3dOxkLiiAtQI3wY2zksbtCeLJXb9B751foWZs6o5Gefjhwa1t+Mt/49zLgDA
0hKLf1HJvV5eGIxyXkZp+7A+Qh/wu9cngwKAC7Epu3Ik9bn8LXYsjMyPvA4t
UPByx38mq2BG8O5mHI/+aJcPfyFqcSFQjJ5I7ri63Bpn8jnHh95TjSN/pOXZ
JHu3urRvU1I4Qt4s/YD6q1LZ5fyEZ/X5NWX9YTmTKV+YfaL6FNcMN9GPip9Y
8oS3ZhG+KANB+I3PPZRP3dQxP63sO2Ti+C3TR7dybh8+DRx5FXtzAU2mdfxd
+ws7lwomPRlOb9kigr1VNeTWXZlmiVujIK0zS/wFFvMETqMna1Ex31jSOaY7
AKyKvoVCW4IhxsBh8t1CrSQYrV88To+t20qx0Wo2nT14WEnTsqni0M5/bY1S
FV5BwHsw7ajHL6OSiM2y9IBtl9xGxa8KBL6zY5QuOSLkLGTW6YUumDKqvyNY
chUcqWDHIGOJalaPgdCGuDtvt6po7MaOODZb/OMvQ29pEdKPAJvd7K6n4Qo6
cr6IBgBsdcg1iycTdT1W/INf2Fj4O/G0sUy7QGWQDR1R3A7juCuetWGzaYMu
j8RozA5woeNKLyo6y378swwkSKdMA8gFhk1yuKXfCfOKyRd1dIbZ2K8uVX/o
n5/MzhU74BgL9O4KDGlUjKlVsLfvkBNjfckaVo3vHFWeJe8k7AXwpHXFAWmB
B3sUh+CpSSDcgJR2HP1K9JqQpTlFKMDVTvt1AnzvaDlsl+CobYM0KVcNK7L/
JLd72MA1+QAZcGUL9zHtbuVHjeV4e0nUkl7ZM1VbUtfh9FGpI6pVdcJoalE4
Pq85y4+QF8AeRtR49e8wIjVaknNRg+ECrIxlbYeXNBIBFUPeo7h4ncQiI0un
qrRHznFTuFmUYJjD3YgsFZRpxx7XgQEeXqF3fyXZRLQPtMe7qCgYm9tggQTI
NLScSKbrQeEUHWJxMUiseUfb0/aXo0tqsBePkKnpVILU/NyBt9Nh4qF50q+K
6hHtLjGB3qQYOeqrQOyQiTHC36hc4FLqBmAkSs8H5/NcCKi9jtqjaWo17vyJ
GKMOXwBwZ4fQkPBGqjnQToKJY7N/py393irKjEPwEcFHRvb1cqGpo2vvHLwC
CjpxfmgXDIgE1pQCxuQJaDCqOEN3KXJR2mSb5xkYSOhDXvp40wTgnq2+kYqY
5q8l+j0VtIcAUzWa4hbqKX8rNXxPqs+mm0tQE0M44g8ZBpeZdXgZgZbf6Jo7
yfMG/NuaGzV5tCQ82rR0DiyJCrf/Sh0ez0XobLD2nY1M9swFL7sUjoRYvlWA
1tsJ0WwHO8TuvpyMJZdb6QuUQBb36+slnFD6/rwQ1CK2q2fpw3iBljTx3xWT
GL6CnmrGHP/581JgEv512WfX5Rp3eXfHLn8qYX5z0LHTgsNOund5AZUx4Rrt
8RmfICn0X3THDvSlxwbLXlXcUk+IEpRjj5bZovz7Nrq1S68zJiPZfjhyO3m5
fHRYccr7kMVoEOmjt6UH3XquV8qNzLgYlHlL8BXNwEeQEtmNY5aWiao7Hw7s
32SfXO7AwD/azkxgbygPjU6K+oYWOLGUYEyA/hLZ6qeUuvu95R3cx/CsNWOd
NHJd2N849eucacYnB9m4DqGowVHQ2rQpVAk+filAWLtJnuUouTESxp8JYJ1h
1zpPILwaFD3ATbkHhax4cP9iY876PBUmnNR2+Jjm7v1kXkj/wew8HJM/XBPl
2jD2rEyQD4ij6Wedy9jCxunfMCtTJiStAfoaQO0g6UN/EBdDMKjPMkYH6nRm
sFkOoZUcadp47Pf8dI6+3Z/uxdsz6o54R4UMD/oTzoZT/GeXHnTZq5cFGD7Q
+NgvoIVNwKcfg/WYF1/b6fFT8TxPZv6JS6il/tEAgCZjFpp7zi4iJ15dWHoa
3NIQpkKOVVZqwSMEONs0M6ZNBUlOSZa6jrLOX5A1RzD78cm7OdO5TGW8WTOO
hC4Oo9g2ZN0wsIn6veysjDqwBiiHCDR2t8TKdzLNgqAGNdISnKHBzXZQFCwV
TMINFFOGNTcO+6xc1Zp+gLaCeHn7aFFH7pvud/1J20y0F7XHrsqYBBTfmqDg
eVKzTHlu2oiJxfjMKDWUoZhP02WiqDPZRBvxHHPmN1ebr6xi030iGrZB+rNl
WvRdv/P2hrMotYONz0FX0i/598YT/t5xOuYtDKUvAuN4a0xXpSk4PNy1Xi7k
ExevKJUn+L0u6h++ZKiKZYdEIli/7CfkIzvTzEzbdHlUo1GpPK9u8IS1ZiIz
sgFyOSNtB/C9oCt6+u/1UegGhyGwK8k1SMdys8vjxPoGYTUaeeVb9gyr4dXv
2kkxCc9dwSQzUicGYLYkzL6PkmbORl0blughYFyYk9qnTR0DOAgFRmN/fVC5
Hh4rzw3XUVAuYm4J2Hprqd0SvJ5VJobO7m0EA15DtkXi7LLxu8pnScX4KtoL
kFM+3EAppJiRrhODDUyrBW2aW4CPKaHbVsofyoDtts0nv/dAHnXuLIt6EqPe
5qBIHt/5I7gZEYL4Y8hKDvRF6jx3tmXVKWNpO8Qmkov2Jv3pMxpglI5yofM4
v4UIw/QS61lbkU+LczZa6+8rTMX0tx15y7K2xz7svq3CB08UzC0+HSe3kzem
mElMV34DuOVNkRvbzeToepqYARvrR2KpS1ZArZBtiexO7791bEc5XKaG3ZWk
u38sdnUw6/A5upKPoocDtQFL14cWGvCfo6eMozMCxJeBE77+VDGasmhEg0i8
nGao4PCQZ4bQSfhY8My7BjmPeA70b6+zZeiZFWvX6NKKRgtGkAR6b7tFZwoF
E5BOft4goZUvUP0L1XSJrr3RzKNe8MhT8LrBrNLRtoVCacbeYpZ1ArkdTumA
jadZ1Vzaw1VxGqM5IUl20+dWNU6TQs1kG0DaWUDXcUN4Di/my9nh695ary/6
anOd+KQngveXaIEwcfSvYWTUpJvU2CYXo2K/le8QlOAxKfevj19ksq+DkLr6
ilAJXCz4pcb6+n8xEQazKE8HiJoqo2F4NwalJCLatJw1WnQ4XzgEjVQKbh08
O2/8Am8hX5D7dTYQzahiiYdDbdGviXfHIGNDLk9PZiX3ItHE3T4/I+U6klp5
z7owXuei9+xvthma2LYjQh5YA/pcQ75aYsxENp+WTKCr5/HjXVXRXGQvzpeT
YHzb5kyOOiyHhoy81Ghd27iT0vD6c7vVQRXMhqbeMux1GGoosP3UtRdVLb/F
Lg4MJmiLWOYGRky3FhHsg4ohEvbRcOMTw+RMcj+9+KbqvOBYFA2YVBS0AUwp
IKAWe4Y0KA5MgVRef2USZdIsuVfpzeI82eR1qxmqOJShvcwZNlSH4kYJIVGF
zWBOqR4/XCk3Uu9iMR38XaUSj58KKh5lvxDjeIViyB+3SHJUCsT5C+DwZm/6
UXrp+VDNyWx/HLv9q3VXmQMzVmA5SJWvzZ6XNyDSA2yffw8Y5C5QgUhyyEg0
mn5qitrl2de3eoRD736zKfEm6VOWZjzkOWXBudlT+onElrd8bZLbNE4KRNuZ
P96ZpKqLnIaV3pr0vO9zN67T8K2/sajyj/oIIDk2arVCtDjxu6i3EEPEVA6G
hjeaafSHGAGCDzrivkQL7eq1QZTJIh9gOGFSW8oyQx35b3GsxE53s/2dnjzl
7J5CDDr5Moz7VqUigapyBLtsxX9NVAvELq8xQrZsBBRKFdN69P4wTSMziLrl
Jnb2IyUrHRvfwAjdf0cfzV2IvStgnUo+59HCzMnDjiI2zlv6WA65aHmuaYYH
Ir3TEEDOXpVRF0RAHpHZheObzeixk6YVW5BGjG5Q2gFI0S6Czdl7FerOuXto
8LtDN4LPrJg4oS0DZ3BFwL0EsFMDWow1xhtVsEfCaddb9ZCVF0PKCZjS/YQl
J3OMSATkM9jfWXdgdJBis6KTuDzo/h+267N9QDFwDK04ufyEJTK1Ja1qjiV/
nzrOcZX3qr4xTLbOYjc1G4ugjJPNZ1IZaqhAMn3wk9IqOZomI/rj/3dq4FBl
u11OpX5j4GfM0IDmTUQY1/TbyaTzuzxORX3kht3yOBw6P3BQyRgtk5K/PbC2
ZKnOu1HDvepiOVsl7qcHQSkrBZWAN5jz6h+QOEmVDK2vKFZkivRSxMdPSsv8
JHNdxGfnz6iK8eh0YnAwd2Jdv7+mzhbZrSbpSRXD4TsTyUIOcOGtNDK18mCI
F2Pe677d/BZtd48VFLzBNEbCeKANoRHSIF62t9MXQTIUuJ+PzA4Ju0EYCKIE
F0BKDSrH7bE8YXBzXTe5uQ5Q5k7PjnB+gNRWWqbdEfSNYkE8tpxkqLjr7gXo
RtJDV4hyVWoJ3kqPLtOr0Hl3mx5qQTJvGnZOZZMC+AZkCcL9BRz0ZeI1F9pN
lYQpuJDo05uQQl41KsfrxA6N6144kWf/3KzyUjtYI/ni3WBXPMEtoKuyE8GL
wvmpje93z8vtXgvEddRxwCYeg2Mjry7Qfz7YNeC8RGrt2nbpEFtjFwng3EOC
dWtfDB3CTWNnWArM2dqouKFpfLUH20E1ljv5nuDXStW2t6O5fOJBsnoRGZka
KxyJ/qyQfr2E7d4b1HJbHShiWkBr9LglYNI/PrnSJ6YL40C2HC3J3I76GXCG
AdeupLzE1UizE1IqycpbHY0MNHwemCKfaDIwo9/JleQRtR1eWXENB3XVOXWq
sFUfx71g9Y/tJwkTY8LHB5cpOC6mzI5wOySOe7Pqzm5bYahx39j4QJ/fw2uT
RPktW1rI+dnsGvUWuzpO0Rw/hs5EdgynGECdlQCG8qvr5XkM3RVdct32iWIL
meqtgOq2b64n739TqH0iuV9joy3ELwCKKejTLGE6ZnaFhMWwGGUo4VkCitGP
5hKcvyn3bUeaXsscHwj20N9njYoF3UmW+1ZnH++OWOksHT8KkiX17y12Q5SC
xuCEYgXQOGXFqVjP7dGhJLTF1nNsU5HzRtJLna/3VRXXp4/XsxwuTLy+JD3i
57d1tOJ66iwsYBuRXi2xbPsjFIoy+M/iclfIUSmR8VV/k1cGbjAf3RqO5ZDG
rtZPZPAwfVFA4p1XtlQHObH51p32DfLeL9EIiIhSA2g/AXd70Lm7d6JrOJxT
kulmkbAx+mtIZaR0PEmPrJ3CKeJA9NJZVulecjYpJgsc3IBwHg1ujvJfauqa
dFUDZKCLDIAAiuonHoVXpnP/subGzRrQhF+bkNvX/G4YBcUulpGr9Y/ee0eI
4I6q2LePLWaJwTFmqowCeqcUuoAmHuhCWmYt7tCXdSKM5SEvH82AOhMFfYyE
rySfSF7jvXNnEbDlu+1Kh7h1EhntmRyA5odAPDYfx0TgEZa7sb2RRPpJUpQq
E3edU2IWcCafVJLYjHKygotbyGrH7unto1I31imouqObZNJVhppyAkn3DJo+
N5f1KBy2tNqXOjmf4VSV8CTgl5GF7kNDUa7s7sN7yLP32+6BzrJvn9lv3rVL
7bCywbliysW+aVatwcAiLW8Ywn1V0kKbpGtYMwMAKr8GXhXjdR+gNQ5ErH1s
Y41KxtjSoLnIN/iPB2AYQApCRp8ONMWaP1Q2WvXAWhD/VS+grbzqBQ+Tf8ga
Cpy7yABrO+W5xV1TwhTihdj/GYb6BGECJNYPJ9McWM3algx1yFLcrYigR4hm
Zia5cHbRlbgtHpVPTFbu1OFhASa/J3PYR8H8PcfTi8IaOp9iMSgQnYCs5bIm
8sQr18wkF0wS0ru7oFJnuRYSbsrvSbQPtcyiMu1TvwcThRfGnisdpvXJb15p
GEdKG+tr2Lp7rJg4f73hZOWQUD7ohUg2DCi0CvwrKzbHyr9am89I/ssZfsAk
ZoQefqn1yQcHupPWYUQTcYhm8Rz3WaRVErRWkJ8Ruu6uZ6UEvixJZHVPb6Lj
RPE5lJ6Tic+3R9MJxdP+J5eDGL6HmqP4reF2wErFiLtCD+5AwwxJjVvoin9+
8AMTPPshRfdYHBGZmnh+FA6ozuSLjwebRuU/6o3ErdhHoNNXAPdlWIUtuKZK
9BqoRWbe/yLZKswwlm5T9Gr/lq5EPqDcFADYYWjz38KzDypEp7HFa2atCh6P
llXG7I2NmeIwgw83EfhSiv7DcwYybbyUrQQr5EtTuWn77bZkZzdAJ0NAkHlj
LpiSioU9x1b2aRXVv7fOdIBWuh/tIVvjS8n0qUkbyCD+pVk0LYHhaSLAVA0e
90hBdktITkWIhn8XtspqGVMhub6YNehyAFPUJt+Q2/Qe4F/2O09oFUTo7r4a
RF06hj5C0Rau06imZ2V9bJMJqrz1zTzo1eMctgpwxvmze8tbiR1OWfcJpZqc
NnMmDPKOYIwtZs1NVkT+pEVFydVTL1xbvMavBmNzSpnd4pYs8t0sMmT8lgm2
CvgYtCK8wro21q5PU5J1XMKzkSSgUaUl9GTaBC/bZoTjKHeOoY+KjZDqqpe/
dXZ6BLK45iz2+YABbTvUGGkOmCyMGHf+jTtWR5piEjZzH/1mxi1c993GFFiU
9sCyH7oNer+Qfag8eppMDliPMcYNDW0wFEJAtA+ak9KwKhMUNsuzPTaaWF6U
Cnqm0NibnbyuDUl3KzaCtntdav/Nn5CN9n47XV0GYMkmgrlnhIkeFbfm1pHQ
AxYNumQKb2h7bmaNrLBmkYTBG3EL5sF3w3WCMj49KY/BRNpTAs756oiHS3Sw
x6kIrlWfRlCPTDKk5G4crrtUNPw9cg8ZSdJ8RGRfMOTZfOne4G5O5pyYoPu6
5nKJemo/1XYZ7E1uioTaifWkbC+aD4GDJeJ+o2Ac/FkbmlwuH7M3+C2oK/6P
oDNV/514C9XFI/fZe1JIrYYN5uET8DDTWFuG9gwlNEMDk+yQopWPim5CgTIN
j3yIYGsKlUypIRM2w3KMwTN8pv4pnDx7Q2TJV0MCB/edLcIT477vHjydW2V5
5BkA8K6LMYDutQ6H3/eQaoZ/h5vxO+ILcuKryxrLGNRk522NStpQRIwDWItw
3FZyJq6yz6WjHMJUTbqjm9OSVJr/whqaSjpF2V92rzX/epiJSLvKBGTJ4rFY
YVTTeFwUNucYwVuQ1LykWyTzenQErwcqDhpx0OYWgczkOm6tO5jiUj+0hqEa
eQabTPU6iRrIPQpI45JJNP6bS2z5/1Jz6bMQScjyYzgZWbe5WDc1bIxLyyZc
2ymozbIS7K0OhCIKatGRBqzofOOr3tmr5nZlW7e1bRNxN1bNsRxqQiBz+Tul
tZfLtWM0jpNLHsgYTxzKqw52ayEiItkhDCvu7UszJaqh+Vg7uHLnbI0UZDPV
6w5/8VYjx/tNjGLfWLYb885E76/8+NjWIOu1omHnK2sayOyp+61Rqz/ILz7c
MdVwg1THNcPHfZjnp8wZ0es0GHf6TjS3YeMezUf0LyHnComWRPeb5bJdm376
jh1Qna2dlScdF38KzBA2ruITg9JnFi20iVx+zBqe+RTEO0gtEvkoQ1GIYqQV
Ntta8FCJzNxbn4uMkxBn+GhsHkUeqHX9TQTPTlvSr58ho1XUD1GJvIzFcEQ/
YJjwvRaWmJhVRHrPgbXImBz2Z85o8JEPrf8p5vOupcLlah48T24XpJjonAFc
d5nrcRrpKFsCsXp+8ayqFAXasI6HmL83gQqIzcSGYUs+MKW0nK/CEXGI+QEe
rtRVUTNpDW/xkJuRCpQsQwkkU75YYXm5S2NbaFGQe1QTAYh94Sc7B85RzVUi
8+ABoPN/X3yMala0fZVecnebzQX34Kl+DB1+8YLOcbHFGwPXhQ79aYnGgisQ
gFPIS9gX7bIlJiZiWU+hQvphqfJA73bYJ8mP4V9f2SIZC6teCFgqQbkjpTZO
fV9fkETQZ6AELJTKyt8vmsv3LGh1Ju4psP7+Qo/jref7jxvTm29kq7b17vBV
kDEEhGvFMK/PbzblHR52u3/XF3u7Oj9mgsGxiVBAT5nd5yiHwFFFeCppxddv
8XZrHu47KcQmcOWb2VPP87cuquGMZu53Fl7P8Rttxxh5E8e3MSbcj/yIrPE1
bOsMNocE3UgQFhp9foMSXqsl2XNQi6scpDcK/1Rt/M5chpcBz/+d/hROn/UH
t6qh67RDmzg2FWtDN3ni9bB6niI5GavStPMcR+1i5RAVmuooDI9CwLd69ggZ
mJzcgos8kS9YZ6vxQ46sHeek0PG/TOMAxMlwEF7POyXCAokU1bIaqnXRj52h
sBdoJJSxVvNC6cV0kgmyIq/R9QalxAkx8nKhwd4mBNfC9iWnfSfQQe8P+xdk
nzAFG2npUHsqgI/W2FcLMZ/wkzvb9Zp6dSIqKjWybWb65BQjn+9hwbdUC0Bk
DZACzTZRXVJhX/7W7aEy9X4EOeJo2QQHJ4mepgqYREPjbqu1hfCxV3E/sQZo
RJ0EKU9h43Nsq5hHm7v4xhOyAK0TomyjFCgpg61C0ApMqgl+WtACTNIYoG0d
WyuIdWAv+E4CW/uGcc3mnvEgIEs3VEEfi56NCHfbRy47CTeoM5uh3OhEg3rZ
BBp5c1V21UUUryw77I2rvBgXxa7spt5e5HxwLXB0+gZXI1WwFp8GK6JBFmG3
t+y2tFXUB6+L3REX72Pbs96N/1BCNlSLgs0gM5X3ImBzDjLfY6K8P5mtPU8/
1NSGYpZoGCkAzwIBr+QLizLRYTM1wibb4o/jaXz5p5iGRkET9UR1aua2znQE
IUgq4JtY4ggKt6bZBM2ZqUalMts62mRzTiIsEe6rCOIvHWH8JapGDrSytXmO
OowniN153q1wkgmeaxLiRL5aHiNClf+xbxYEasiPO3x6kUMqFvZ9gx6frKyM
HZi39Xj1hHfsQ4DU00oIcbErsh2x7PPd/FNPg7/O0dx1iofhiUwS4KOlslxo
5zdxuJrWmvHy8r3Kh25/+6QtdP3+9OGDha6zq/Mc/llBM85l1CpxQ8Pz3OXF
eeN1LYV9c6ectVx+11phrQx/g+Yx5Ihs1S9OqmjAAH1syVf2QdLUozjk7bLJ
lwplatlFPEIr96pLk6iDOJWN2lA4jWImZbEPCQSl7Tz6McR3c8VvyyQE0Ycj
Ecbmpp5Z9+JQJyT1WKNvj6+Jl/9LFowNRMA9XSlsno/Iu5y1jFPSVu2tJjmm
L4b7Vh+hZ3vShdI3KBW91GoYroQfi7tt+3OAqdMz1sNdhbX6DIreJgspU0j9
C9scmWCi6gADOH0dsZmPaDPrHr/CD33cm+K/MPBb6B75eeK1+msRKTVzW4CP
+F1NrARrZt4rF8DJRxosyc9Jb3PNLZJkzQymCHO0EKtyFpAToNlRnKYP5l3s
1XKxLCxZF4OnqoMu5gba9e4lGoL7NfBvt5ijNss1vw440DjbQzaaAYYoztdm
+uGcDo7c0wKNW5IHLnNokIQ0L/Kv1a542qEFz3/JuaZEgg81TDCQ+M2PhfqH
blcAIhLM1iqN4kBYGGJgoJSkb5y3weZiJP5Dwvd4WoHDEYEpFwuwLqyf4siR
XJD9rCquBfuOc83lebVYG2jxCduIYrjBVV2jj55VjiaLdmVdE64jaJtVYcHt
nR+bnOpB3RheugjscxlZscEWYV3F3kUdQag5hWlss4v3prm5QL1Nb3W8mqqr
cGC0Jurxw7t1b7QxbilSn6kwP5sKwyc44pF97F6c/mA/Fs8sYmOA/Pqc9NHH
NcHfMTpnEos0KhtmS4ZCeNVi91hes9lamG0tsIqV3QnAWTEhW1f3dc89ctP/
NQYBfaw2hQZQf8ft8p2Gud1kk5i+9LUyNIV/e5AInRUfhUrHRO+GSo+e4PX2
w9p3yLsl5utvim4f2fD7iE09nBKsUfEybGXrOZEgKsvSYUZGbRCq8544yeh5
8mqr77brHvau+5ZyJ1bgqaUmthJvV/vEpfCLstVmvx2ueE98Jj5tB0nbsdA2
FvwtGULj6sdCnsmIsFlpbmVwWpTbVRyhYXEWryto1XaFihfVAqViePYmj51V
3yJOyrrolOnCyaCgWQH25IvY9IyDRlcdpIm45pTHjDPt1oLsuo9r91TEF7wU
tfoLYsUWO6ObjDDRQbZbUrD5u9TOL8ap4K6YW6wImMeGDU3JCoyBUvMUHdpS
8pa4VCyb8NDNqKj4/aceHKUfK032q4wCueURmIzz+O1aJHO0dGiWkB6x3EHE
TqG8SOsCtoiUMfhcD4rDcWvWxMJDV8ss881DSPssb8Cj5HjPprnm/GUXpkQO
8OdMJw9ZIqER83iA0Bzd5fAS98tNvNmJvirmI8HP+6Fvdolg7h0YCaWjzwSN
lnHkuy2Qd+uvw85QNMW/uq/lOw6+rJLof02ptjZx7uGOj3Q7XdOHRDAocopg
+jgeJGq3qN30tIXV7lbKzJnOoXZ3Fz0yjxHggeTxMny8kfzMEAbblf1OvYYI
zNIYpSVRv9vu6Q1fQ/Nsm5Ljj+VKPY96/qmw2+W6LflBMarVCEUq/cbGb4JE
bu3NsGRxW6wq/GYKW0Ap+lfV18+dINaEpBzHgNLko/9+YUs6tHwkEILa8bQf
ubY4o99dWT5GHj/KlTYBu9aHkSqG/xvLGCjq+c/9pL2DLuGuOAg0eTOo7R1l
kKTuYoAWMqjD6Fxsf7K0KWZQRtzRXleiWpMhlxiPGPTKdGwKBFe0v7Bcxva7
lDrG2Cpa93opl62H7osby7SbQeY2CsS12RT5dVdoanHnVv+CUO+CgxfIGIIg
vY9DUiDeO9xxenPbeBdKHE32a8TuGL66vwKgjeKGZA96FeXXg6ZrUjR4FoXg
TY73drKfzP8JbMpr/+ut/bmvZ1WwEWSbh6Gys0g30adyBvVFtrTDPDZjzvR1
hTpBVEDywFmpwB6g9IGwWzxJO40hD0lYKMTmTbEm3UFJoo7aVKGNcKOx882i
YW/LkqxmTqfRZFySeXLR4rZpLhLfB53Oid+cjihSq7HFQaBk8iMIa30OF1TY
l4sRwhrMWewMw3pNeIFs3LqcqrnvtdoUgkYIJIv04wNiAzilZjSYHGQ0ykwc
/xlRKIOtl6knbMItt9RJGxua+xcdqwNyNFHRb3VJE7TTo+xL3PmDvhEYpdhf
28TAad74qdsIvx4pRY/HmIqUf9zcOi83cgSIFUxeCu2PPpL53RJU8MvQBHos
cttwKr5eJzI9i26oZxxs6VnKK0pKM4161eBIFke5p41InF19seUPIkZlkTAj
rJFbUsPWCvvHyX2Dv5Twwnav5GLVAueD69+8gGXhuDOscpDU+vYz+/tnCGj2
5zDk7bH4QXvq/QbgVJIPV53cidHr6bbdGbDYY7YOtVtFlVt10tItFS5eYJZJ
44FFwzICYJzIPwgUjEyHz5kdm+qeub8SZD94UA/cJbDl0LseSLCtlns67cHD
D3OHpIsSVDxHbf2NCDW5b8umyhkhMUGMHuqW/ttm6HZlsxFDRNcyyMJZSXz3
C2aSFdkVRWz/M1YRMJDS3ic9mjah2m8UrNIVVypPj4cnXJYDJeDiLrRHiuvK
QpYlv5v5wlkrZnPnhZoK+Jbklpfx+ZOF9hQ/a5C2tg3E8lbWNTCnsVcea5i5
Ls4Ea/6TymBr5Y8McFdUr0G2/CsATJIseQT6dDsDcKXXhoSo72MkZuhAcuFZ
RQUXVvoU5xl3/NFt29Cpn3ycmOGMrQNQYkU9oOBnDj9dW4mDuLjbZcAz/1fL
05qZqK9e/3PDEPdlmtv+ut2774KY3bwlVhsVpaO/JFnqFVo3o1NPsu9bd7xg
VAjPmw6vjiiPK/6iPxPmqx2SMtVMk/aG2nDEuKk4wvsIBy8yuzMLqKPwW9Bt
HhdeDK6JEjcMSvCriUJWtCmN1JXyVpNvWWmuDA0Rcdmyhdv/KuIYWvTzvMyc
k+PDIJKRwSAWzbXTFgpwkK4OIMGC9aFnxrvJxQPmEsvkEkDkZ1ZHuyxWn1IJ
/D01YHldXuPEoSUL+B4Oevp01dmXfhYxyQMG/t3AYMwqGmsjBiV9K48y5Yrb
kjOWzukKHq3PnPACBDoiyGoqAP6eRV8bb/ET1QgzyzAdPQAuCOlFlgYkzoQS
QBR053KPWoPRf6UxHbeWo8xQPkkFyW0kb35Fcx7g1bTSFhptBv8F7wzKfoO+
QAfYz4f6nvmupE9npmixbwNPOJCrJpxIvgTCHp76hzibyd8VuKu862NC1g8P
w8b+iz/gxLvW6matQbaZmDRSBJt34qoMYgAQqad6KTp5MUmdiry3ukPwoV5o
W5wG4pp0VMMGDtWuOh/HqTmFu+Qgq6GuJ1eecmojxJN6UBdQPPu2DHz059Xd
w3Tdj75Jdp0MyjxLzIpHsZeJtjqjHGO99OK4ZwTtCki1sv6iyJz3e8PsUvPW
KS0yjcEANA9xKDUEue6Y0MUyOSy+G4rJ35YRYV9wPxIpcy+2BuzL81mgAEUx
JqrKk0Zx+vD2vdS8uOVs33aaEI5FdR5pdi9X7YZxIBMV1joJ3LNIlwlXLhgU
PkfKMGLet0/5QWGVNgCmLIrCUFDgpFdVOpQfdpgyFHzUIJH1IJH9f7cIj5Rh
K7X9QivR6gsrn+C4bMw+FJ2mXev19i2x7/Njx0VEznvTtv0uAsYidciW5a5Q
e1GBbF15KJoB/+EO3wYi2+m0nxQ6+ajOtLYrrM496vzzlWpFupCMLNQSSLgL
DA9lShK5vFoCBC71X5VR5GABwcIt4G0xdS3LLurUpjMWFPL4fhyJ23oEb5sj
2xJzROwJQtXKdMshdTdyBEf+BFCl8w8plOoBThyHyZh4n4XpDBm/fmCSjgql
PiHPg1QHf8F/qY0Eq3uREROYJHOBFM4ocmAkhXkDA93x+FJnC/vbRAg6FmmR
uZfQJsg4994bXucXkyJq6+YHuUzIN4FnKv0e/fBGbahO+J6YGzv2iB2bjDsa
pLEfKdEySNIrKoLEH16rx3qToIfU/08dVPzr/XP6g12XkwUhi0io3NvueLlv
r5Rr4a+DyoSyqh6jgHqJhouS0qfduSDgEQYnsJfF40ASQhlqBFnDvAc4AIo9
hnL1q9ujYlq/d9t5UUk6NG64DgOM5DhjaFVHtD+HbnUVy8+KVg9YFLjFplWy
/vlmhBRjaLTKMcELUZjDpQM4XanktA1btBks3EqVHLivWOoXypVVI60BSsWe
M/HUmixWdit2pYxeF3ysQtRqGUrhokqzOdIXfNTjGUkkxAA9VCQoKL0qwoaD
9K6VzMsalZSemSP7BaiEAZR42qEV4GFhE3BgdN3EDnSXohIWRZNYvFDTbeG9
Hd0DGbsXGob81YXd/FpazIJlXq7YGD7P1q98SVaChzBG21DUEVNds1DJz0zV
FPFeHjP9zYXHGF4EDlUkG6x0nPYp+tf3r3DwIuRTWIWjOsJqs2B3j9TZKen3
Fluf3BzimQm66Pi47pdgG98h0ItUOD/auKHsPWvkirvzJkWgMgyDU+CxFsPD
RLUyRzwikTYVZJTwOlVPW7GvqGsPFcqmst67yf/CQx9wxEpuhQJztIqUklDg
YuxKeS4GnkeEkYao7gkxYYs4ARuifbcwj1eMJB8oWwQS/hYzg9yEtiOsYdUt
gdsJEoUqTRYsnqhAwb3Btga7O1Pk07bvbxGP4EqJi7Mz57SnyQvICC4qJ2Dp
mEHsF6P3rFq5qoem54otPHPNrGIJpGfkaNLyDuFGXEO2QqXfuEp4dWAnt31k
daA+KsfBhonorWUkCV1J4yxZuWCyo0I8SJ2m9TSCukaXvZkPzVwWqsLdF7lm
LaUYmLNQd9/gcdKpPH+tP6+gHNmjg2J/eu/ueIocy5+pi3YWxziKYFskaXd9
leUSNPXTZS+Rts3itNSd2AXtilVEiKqyp91PQ41OQAyzS5o/kVJI9J7Ybyd8
M/NqtMUhqB+F3zrO213P+YQ/WI1m0Y5/hAPNfYPCW4M+AOpQGiGGUVspmQQ6
JfqOhKH60rLZScjapsxQpMosFFpT3c5FTGKNhTEv2wf5CJhWaO9Olb/xTKjJ
SfzmESCKsUj9yh60V25c7lrtgBI424f1h22ouykZT8U1qDnQz+1kviitcmKK
MXhxidNRIOS+GcUa0kScY6ZB0EqgMt86/+lToC+j3dhyxvIBAtoBhJN8xiZm
n+RYsy0cfR0eKbg3DvvWhQqtQVjVu1UXU01fKe8W8I1YHD1Tfl8YC5JNvbY9
nFyTVXuzwG7HbxtMhAzjgZ0d0LLMyDoTr3dLhxQcgRS1tIo2OqBnJFJmv3St
7tZfOsn1EWSu53wyNiesxDDkFJIbDJOa4IQzxQROp6JGQS0DiMjWSHpdsZ1F
Ro5/GG/3B1O/vNtlm8DnEiVchnpRnDf/aW3jazEoLka5MZ9aBUjpNQtB5WpP
lW2q4ZBdvUNlCBIWqdGjhqNz6K1BQeTOD3JW8EufdZsLLqrFfHY2NvsaYjnx
hA1qenSQ1SUvlKJ6zVEvJDizwHFjL7GbKgvcvWsgza5ncDSYMbcfH14wSuON
LmqsnL/P49G+L+eYW9PJeAaE3NZWa0cBmI1XJnciHBAs6ar0APVWxbEVawaH
T1WqIQ+ZRs8eOf9FFU1O5w30YSMPeJiGYF2eLaH0/AQ86zuy7Lwsx2N7v7AR
IhAHpplivu1ZToG6EQqoxvi9ot6d2q1AhrsvcovharnkxWDMOUE/fvERURrw
CDjt1cdHP8zmx7Y6q6KXTJv9Dx6cBH8h2Wmcrw/4wfRGvIJeZUshvgDPrPLm
WwrG/RXVZmH9c4P1A50FlTivwzGjAoTLWa1LAxx4/l0c2P/qvdRXZvzvvoui
04x8k8ecKBF2abBJreO36am8gEeBG4hi06Man1/ivEiCx0y9/3t3v0QR+GoH
/fuZGMwvAW8c+YoiiGhwqYRF8aARCfFH4BcOyL+uNPi/LlQ7PWtJc72JbKWk
cxmPeZeONhbXCzsZPFp+EgVFoEbyCyqx+8HF2yiJG9hlN246MSUt7hI/wL6L
FthEryFYWWkTgawhe8H1X0mUnQ95LACZCKcC4gY6KG4Q+EusYNCdWx5vMfH1
VdcHrx/84w9fmnsT68u2tJoYUBs971oy5KRIVh09OumY35ThXGtYydVcoyYQ
WhqGz9KlQWALlDkmNb82HpE0/mF9TDPfCza9Bn3O9LWrSm2Ppz2mYMDNxnWH
oGlWHhq2RGazol1xQPYieNU5z1Aej/AvuwtnkiQdk1O4tVf7LpfSAgK62J3Q
6QB6I0LGhdcPN97k+fJYPM8Gj5dKi6FkLtuv+aZuS329IVc04eX1h1SUUJqa
+SDu+8uJj1T4Ozcy9JAJN0xmaCxrh6X/dnmT80nxyNUQ6zFY2YxaWPXnyrPa
fAuoTIiUElcvS/NNmOW/o9YUmXcwZpnAqCfYkQGDMAAYmAOK+TT2gAqyNpzD
dXOaZKon5yO5AYGuZupG5O5P/wHorfTgtujlVfoMkIeNDO9tkDADZRIa615W
8p8MFNvG+XcNzs5oxEiXlBoxDVdV3zEp5Hop/MwA3mLNuaP40aHHLI0EPkM8
WEFZTFOezsaYAhZXFJ8zb/J0SBPmrLlgfRpymi11JUUWA+EHzSi2dL/8xBfq
6tsc/u4G9HzpWbiJUZgT9AK9N74NOQNSos2jqGqcnLEBR6ERQgwnpHhCP0ir
Xqi5BNLa0neixi9bqD9BbiQc4CfkWVytjkb3hdZB7xJcXQ5za/g8K4wAYHDs
22s3fFLDoRgfcVCMlWTIeYXseZo2fcPrUyKYy0rPUo+Ko7IftI7udemJE9wD
sdD2U2U/l+8rAQijPY3v1rgTG55071ZQIpUI0lASUF8ywCqILhAyRSL+eIC1
QaXop3nff0Z23nFkT21o8pRdQD8EUOuFKp2Nb6VgKA6uTCH8RZmOnsOb1NMi
0BSv1qXLrbP+xXyAQ6W6s6+IXUusUQer6DOngElVuypHHt7Wjt0qVbXJYWG2
oeBxshBPsg0LPeKiNSpHolNXzCmTYvSAK6GL0OQC1YVPo0R4KWjzfTwl2koW
NVs/KWBzqKcwPlfnRhtIrcofeEysXUDRcIoT+bU4QomJuTmYaX9CV+dwLbdE
HKSjd3tjx4Zunu6qdRdHdPSsp5YboSYp3XokG+hzkAiA9nPPlrvqCVAhap7h
c3cg9YGe9cZbJJ2pdS0nq3w0di3Sc4xuSG3z1UvoZBW1a1RnrpaL4qgVpGic
MOoVjzKqqGcEB3goW+KYhMamBsLMOhvFs+hXbDJQtXGfQZbFXqByUhWyNmmM
VCjOfonPm26SEPDC20aAncJvel8veB47CbgSvPrK2lQJkob3gTwRVf6VV4jW
yfsiOEDFOaWTYs3ldqA/YToVoFvC/6+/0NFNmAk2SAkN89R0P3QDKlfv7Z2Q
aH4/1Z3suZfr10PpMecVJsf9LKiEoVisjpEHJkUPqIT4pB3EqIll6RFJyNbm
ssv+WSLBnO+QQZYyGYhq+eAUPD70gPLGZEEaJX9GCTkSaj30frTK13rEQJCX
gKPhOIasZSjhjr0rwqmD5Q4LwkBD7pkIolBYPrLbOpPIlV+RGB+AhX0auKMW
E9TdMHJfOmKsBqwMdrNjYayCyGZ39fGIvGaSss5w4N1sJCws1YZonQRptIL/
YhZysbsfkDatbFgdDeIU9GayAI0als28uw5C5cGnCASfY3Eq6SlwX3DVgMWT
ok46tvB0P99Ot6ZI1sDOO0sVlrN8POzzkJPKia5B1MrdByA2JAHFGwwsJof2
5IDf5nxm9NPUlt9wWnmvad9e3djraVUA+00Zz0EKW/V4SYm57lX1LF1eQPXM
zswMUZbRPY3uPuNa/lNEAqWzVsOmINd/y+tQZlH7xxOQC31/1s3BeChDEtp3
thFiAkohKyLMItpAOnHhQP3LRWT2k6lxAdaFuilQ1XL5Kuuw4h7fkg0OuVRb
OKjqm3302U7MGqtyA0CSq19nKjYi7LqhcadXcURBjfTh34oF0AkheHPu2cE+
wTQPqSZP6lbV5by2KCb1VG7Ia/+gO9U0hxD7k8evPZl/Srlu9srYVoqYZ9vh
jgB+CVVbLLm/XcNeyNh+K1fPiGcAfxN8rg7W6tRfS8ICF3H7ragdpO2/AJBG
Th6e28FXgEeFe6rT/Cj+skiIkYzVghK46EZGeLpizojYRLZLzRcE9w3NDJWT
rwBhqGgerK2w7X8xKEMaVS80XGEYrQu8pPt6MhplDs9UzZK/0Q+FHYi5kKMU
r0234CNTjB+vEcuEeB9jwtZFAHqNk0NGqDVcvX58XqY5A2wk9Gyi3GsIlue5
+Yck6owVRN5My4bIzJiD6MJiZGZvgldAjV+2BqrfXh33V400AzjgJ2nbLd8E
F1IrdGCDXEF5dcm/7KTeK17APEoAqQXFq1MeBcs33dQmvzH44S4CHn0u00BE
HxeeILR2xDZ9vphvVOS24S3EXkyCLxCSPyQjAmLTwHptNZ8w6hac0oBHy/2q
jb5mdqV6vdg7o2JeKN9ybX23kto7ndr6D8A8um+8HOvlNf2ZgDpL+nCV9BgN
ING5yMojChPeMPQMqQDzXwu0RB4AJbp8ZXKSA1c5MzhW6IBp15LnV+gx4HOt
VT8S5MtS4cNtrWTG9B1bAC8lJb0FIzUE54Rco1BiUGsKeXweHQ5CmBoJUryL
tmLIeI3y2RONukZmXQIqgWd1+GzqmwTtK/L+rgCH/duSFH2lYh77zgPZXK3d
5y0/rv95jIngq6Za98qgm1+YeovDAf9WfVTjaacJDN3XVIGDnXss6cMSARVO
N2+VMoEhLsQ1O5ul1UbaM+1w2vlhrgLCLX2XxMOPHi8uECrhhZf8KH2s5Jbz
wRJtLC680gq4u+sRYunOicQoRcTAbIlw6sCFlnNPqE+zTtk4/1eT17UW/M2X
14Q/UE45TMC4uvF7irjAj+4DdBT79POipDg2yuo03QwlfciSw/zvViFWIo1R
N8vm/BlT4yZiJdQ0T4f1Cm32xwfG5zYn+I41fF3OgcnhdfoozZGtw3iv4CiG
BN7FAW1T+BAuPoxvQtsmfjP0Q2DnFG8UyPH/Y+xwz4qkh/kFMs05C92XFoUR
zgRxFfElYOXfbqnAMcHAJjdOaWdAqGnhte9VRZjeK4N/hgQ9kP2szkHzA+yk
hvyKFveyBlJlQ2j9H7+a8Dznxm/vjbdicZqMNHtG/1iSYEHFf6gBG1mBCq3O
3JSR3KILl1a8q7CohQ13L2eo7ZuBLdwh5Z6pIeDiCUP8Aq8pazzDuiVpsr/r
jrAjW8wsqy8UcoCNxavO/64dIlClyHtBmKuZtxre8VjUPLXICC/rDU1PExgN
Rx2JB79SvOm1ymn3xA0rk1LY8rdkjMMUw/RJJ/lgBH9HKXaER/rHDGT06I66
6kloOzNf7+gNKMmU3z1A666cMJThj+XAkbrFJhRUKOXwNWNu9DB+EMT/uO/L
YabXE2pVa/7BVupYykZif5OQAyaPUbFFTGTI+ToGAUkWKTTJcXu4aXgkcZnP
3iPR1731p8P5rVcqV6y5OCbm6gapaREGYupz5vVZUgRi9i4cZa/mLHWMKQRg
bs19g52KrkLlfg9i6D95TCmtt0RYfXDmjON+hLUTuSOCLFhkAckJMyZkcH0W
+2USSMDS7qb3/TWWMRVtH4bZmRUefytB+56UYlrnv2Y95LJVB4t+lAvc6CJ0
Z2FuSpoI2GmG2pPhxAiRyBru6qTW7CHCoMI+ZUUUrZ3ChxwZT9Yu8i+CPP3j
BlLVISUf0EYRPLu6OZDAKjxzgUfxh1uFF/O8U9LVwV4k/IcNpJGsvQW+w3ZV
1MtQasXI/qp5VCocn/X/z1DX5TktiN9nxeFYNzYQf8QmKIikaZlVT2teDfA5
Y3nmzDpw5K4+VkNvkNirXpoSXn1EwpUir1ps+WZKCnM/SKnFya1xtxfN7xdF
9SrRjjKTeoBPpEyDwUzhXWCmGz6WojhJk2ddePkTiwvEUFJLSG+T44Ncz0MB
HS9GsWyX29+8rjpz3P4DjKXqEVn9I7ecrgf8TTcTJ/lpSTzGvi643s/UBnKE
GH24AJVQiICPrAZXW3hIu146maj4inAztXjdUDXsOM2NvhjAL5UnLEa2IXUl
VAc76CelKHoBPNMJJmIsdexNFWpi1eeaniJeahxCfYwWxhD7Nmekt76hm3F+
IFTFIRwIUKNc+RkOTCtx7CZkC7ZznBRZf6lKzNiQ9CD0ts+KAPDbM4eHiE0J
D2yy+8r1fsg74j20cly/RzY1HEnhDSr+sJAiQHAesoUUUVD8AmrcwpFgpxq9
MNKzg/F7HRoLmvMSvqU3lwqeYbkb9GLkV2ADT9JGEG7Lui10TC5V5fuGBjnc
okFvvjhMStkNoAzS78rYjr5PqLiILhNVdM+OGqcp4AUSH9Kztp/7zJxjnkhW
FW6VSRIpS5WU/FtE010hW+CTRxN5qBl/gttnVvpE78QRoIPKcgzNlxg2YgWZ
Qr9Fx2H8KwR3rvgwvrh2GHbcudUNexWowcQnNEdTs9G85MvAvpSr007X2T7l
iSSyDmmFrDs8jwfdjWgOo+FtMMWHLMZGYrE9py/HJYhTn66Y3OhgZYpJ3HkB
EZ/PzriigvI6w8IPVl15npsH6rUIH8j5aH5fmhdzYo9AHjVtokKVciEzk135
sKCZXdcaE3zKXP01ehceeG138cevmiuIN/P1+hpyGXdYjk14MRs0/YQnVX6U
TfpOXuq9/XZerrQDyd8wVDFYNtmTT7g9/2URzWPaAPujrVVB6wQcwkM3AN9Y
mUe/JqMK2v4q2q8w0d1apkdNPOHXfb6eXx4hxvVOOMLbdHQwe/8/q7kXRVwh
zn0EHqBL+hgfNVUvZt/u6BFZk7Kfg2ZNKSeS1sX2OP2dYuJhT45gR2IpkGXp
KceZxwmJeq/859uIQ2KS98dDLBzAAL9hLuIcMGOFsssUxC30J3BiJrkKcl8O
qM/cedHMRMWcItDPCE0OafKo9DMTMHG4myvebN/wws0k4gVeMu9qNxRH+aO6
0NgXKeVQQkN0ORDYLTEmKyOPo4uP3wogJQS2QJA+SpptBRrI5UJCZ+24CY15
AjLg6iBgmmCoNraYIf3Mv9DuY7qzqjPl82VKsyPJ6ojymYwK6W4jMN+I9p5b
sU8BAirc+lDn1QZVb8Q+P+cbwF2kkL6+dE2SDE5KM+M1ITNFKNXoaXRNzb55
2f6SjvFEiIWHMhUcngZahX09SmEKogij5TyCpjQA+kCTxF/pFI2HJzAORzTx
WPcL30mnPnbEnE4nn2jyjaeHYWRDWmgWB+BUFPJHrRqYpyla7sBJBGpjnlQE
eiKN0fqgROEfyEUcPSNUxCGAmNgJhc92ZAoCm96KUnXxgMiHQwcRf6P/UgOv
jHDz5wo0vr74BXo19pp2xn89KydWA2ghFCx9zWml3toGeif1nnAGLdxd9p7k
Vn0HyqekOMIWs4j77d3LtrmC3f1XGSC4Q93YjYMs664D0EF8j5uQuODKRzZm
DpEvuGhuoZj+blMDbS1J2RJ1D06lG2Irx1QxlDfIwZDLSoC92i3NjjCa6Qgc
uTYmd7J2fkQkJRC9feh1eJLDWYc2WL9KTyCeZ4w1JZYi3wCTURvGePYOCHoW
8A4xwkqypJcsbfaUiIiypfxBj8oiz3Yktx2JJJQlrespP/5wpth7OgPqxnKo
mD/+pNAASjLixUjdIAwxI30CCPOUzPg30nOUlJRJNb6QwTz9udAzqorDmRTq
yyzZ4cs7vZrMgOultHzUZUPYq2XdmSSBc8He9TQpnSYYcb9dvLOOMPX2ih7G
/Ynp65Ty4esUMAz6G/Bwx+xpAlMAFZi6QGNxlrtmmrlc0+CXJ8o5h+YaMNRH
5KCPxzHJTka+/+lAUT5ClqspJCUXUOmD9TgeqPTsmtga1MMo5rEsVlYhgyoB
z+q352c0AAC3aelig3sxmGhXp1hbMgW0hkb1+Ms4Y/UVxuj7LN7i3WvFjrCR
DDSfT83I5NKYmdyJWifrweNuK4lOX4NjrSdiDBRITr3F4YtQiRm28OWC6Wnn
oyehFSnd79fbL8oSnHPcPyqyQvF2T6z7TsJBZq2bZtgAYZ4WBpzzA73kiy8a
pVLScGsMtuO5TKvATuLVaKUZ7bwbZ4jNtgtW4lYDCg7pfjpNOYhnsJIPomHu
PVNKCVKF61GN5P1fXypYcPpRu56vITMNyhvnvp+Fuyg4JI+QZ0kemO1gFXe1
LiRaN/6noXJBjEzurDbdRcUQgqnKXL7ZPhtAkdI8owSrQb21g49SH1eAhfjI
8sBcv6MfKUjmm4O7hXtREH4qbxUq2T5qN7235vYQDud8F/y20JOZOhbmWgAh
EKf690/6jFgDo2YW0O1VW+Qy8Q1PA5mN7DUAaQvuKBOd/WLJzLj84aL01T+e
RgdfApsk6uRV3DfDSyyXf2Zq30L9hwabh7b/HfgXRVGjJSogTYVKrJLmDSCk
qw9mDLMPcBtwa0vCijfhtVbGFvVFBy61ed3ymKO5UgNJTZsoDjy6IcVzQZkS
OBEdgJy0ZIIghmzO0YBo6TNMp4V3q1Wz1WvnSl0mfrvL7xTQ9XB5PBiUi7RG
SJ2xRpXRG4nE0covhFAYnHOl5bGVmF2w4X09+JhRa9aKuKTwftbrLOZ8LaXo
MTZenpZXHoNo9GsxtrtJS7aPng2Yx5vgOi4IsdSmRS/oEepv8AcaxcgiEfzh
W5ZBsWR4F+yPDL8AidZilrEHXbiy4aqEUzIAtmP/oGWdzIlJVEE41K3FlWR3
YXyvfj53WH4GVuqjnifJMT2sRvitpR1syNyONiSwB+/ZQrAvjAOb78tDn1gk
NpCi7W8umky23ZmYS0KqmqfwDRMrj72nhMI+xHhiRKaohOdsQmloyQbV+Iam
AcH4mC35pbsg14s3XG7c4YPcvCqLi98SVNdWb3AW9Kym7VaRAj+25P5pBF2L
zjMsPe6LtXp5zxqy1UU8C5eo/c1GHw+eQVrvy/eDysbvHEOpmpNz4d5zFmh+
HGsb55mceDTpKFP31tjg7NW0Qh880hOyADX3Jjdw4ByE7CUL3MUY8DXicyzq
rk1DGSXilSKGZrLXPUPA7og/XyAxuyRcBTA/RqZ6vYZ6nOV52eazhZmEatfj
Xx5upzz1bRqK+n0P51uQ6B9JU6r0UpG2h3MhLkUDqTwv5p849P2cB3Nouog6
w/YwjE5TPcDZcKg0plpGSxAvqastVgyHzv2uEK3MgQwouWlMJaa1UCGl4iuw
HyV4yfsyZ1migdXXUkqp/suCygkWb1R8q0B8AfHA7TuG4J963M0vha5/81Rj
7LuSQzHYoKTPxG4BLg4WwlNcnvmkj2W7108ZWNus1p0ZPuGK+YBFj4eV1wE2
PPwWE+PrOi47c1x7sIDMjPc2O6mG8ijDqMhfmJ8QXRal6EvN8ZXwk5AV5VGS
i/gu4B4gj7vADzZ6b9L1dPBg7ALuQxYKyoOtr9cLtuOcoRhWoIR6zVuaKK2F
DREIv8xeIifhC/a0mTnivyt8AOw76LJAA6hWj9cjGTu6MsjJ1y+B9CjCcSDR
7C9yh9GcA5bMsfziNbU/aJ7T4EEJJe29ORxDmxUb6rjugJrQ2u6lSKbsvyZb
27Ls2ffVGPy4dJ2RxM4gJT2SQsSpJrBtsU/2jxEBwwsw0u3G5laRy6ogRudP
hqY1IyIIj7TzpQutBS8q0+6EPvygDok327AYDXHHMIDIPAWe2Fch19dFWdhD
YoMcG02XaD7wGFBdXxyXa0PGPwG8NE6TiBV5d+9iKtO7YZ2hfHcHJgL/G+JG
05KAeUxlwcPPIC53E3VOjB2d9uHUPP9rOAj6JojP3EX+Pkwf6ZL+1gevv1vv
qPayCpHwmiweXboTZk3wm1uJTI5c5X0UhSC41X7UKWGfabfw60VtdHWLIRQZ
HIVwTvVzZbCE3ogVf0f8e1ijZRDZQWPbsaMD9USwVRXFC6Y/kVob0Qv50atm
Tr/MAp/gb13lYtaG6u3jLSuwGsTDnKFteUjrRN/Bm1hPP+eT9aNrwHLJ3qkV
sSYFWG2DLrt6FO17duGaTtkrJ452VxrMbj09jn77RRr5pSMkAUl44MFMsmPq
Ek5KqcpWPKjlBoUjVStMM3U9EB1M/TpSVWuVFCuSqEGE2Tps/sHaZoMQVulc
W6lK8LtZF4aYqZZn4sCC2mGBl/mfNl2B5VcSrgz1U1jK8q5mg8gCDBtmnxdE
R8OcifGAb/u0xg/iERk+7P7UCS4yCmE1SIv0Iea4U/arzOEQtnv3ZT2xBSaE
FrRFWkgrtFHme6gCr6wU+eQUo+njoUpTOQSEtVQhrLbXqNr2riRXKNR7crp0
iXDKZ+5updMZqxAeB1AhMkg4EjAAbg6V3zWSbttDNwdP8Cz7qkKVMmc9uTz/
xzNRVp5OPAuCYhQas9ayZMR41yFdk6AIOe0XT6eY7kZwxmjcdqRtsixs4Crn
s9W3TF5AjtWhSXjUYJCXOgg1Ky6/hafAv8n05ndSWx/vOBi98ad84HLlhi9j
oWyh2/GNYc+Bh1d8aGqkW6fzS9GJUPw3Jp54zhP9OdIm6HgD6E5xpnwSKwp2
1u9mr8e3W00VyjpMd7kMmQfO9LrxEFkEzRcFixS7fqmNGj0T7m6QI/6Hi1VE
Yd/TG0m3F7P3Ty5avBmw8h/twNrOMUBHDmx3xZnttMDlmfkos1h8Wd15GNbU
wWGTPo++UXOH7gg6kqk6QyjNUWAdgru1GOK1qfm9qvP+SuMqWSRosrmwOic8
AOgo6t2ub0sf8oIXggR2PQPSZvSdvkvJt01gdA/6fPhcaeh60niAFSgPneTe
uFzJ0/H2ZRWFq2saVP4DiItjPIqpVSxBzXTe3s3rKGlAdFnBgZgvDDKJ+BLX
Gaxapytwia8AK9A8ZycrIysZemYNI7Tk4rJmGveG7Onze6a5Nu4F/OcyCGz5
slpc5VO28N08DDoM1YY8BcB6DagbAdXZssgrSRgQyjAn9uIxEwMAoSnZ9hYi
zOTpfRH4DzjZxxmpqykM0ijQAOE0qomPIdtm6hVtLOtEkLgbPb9qINIjs6kI
F9C42PjaWzOQoucbz4WRbeyWPcEjsfI/aaOJUcWf2Z9nEKFuqJBYbow1vTtH
UvcWgwMN+MXaTjEeeRradPg99aazaAIsU/77LBCBa6EHM+mCFCwDTtbWU6BT
w8jZ2+KWT+u/pIXx6uV/4og54GrLyDl0RioVZ65LNfOdKgdxMll19bUAj1ii
745q28y1nvyk4q/xAJDNu6qILJ8ZmzRUXVVSDWMJSvWms+uziHZcx0PH3R+F
uljsAovamaKIApPcPm/+oY/aRsxggO/q7LIW2/xU3+a5YPT/m+VmDWP1OIPq
opLAObxzdvFchfq0X5ZrH0xQiKTKF5cKkUBkz36RCpHifdX84IXFYaT4m5Rr
FXhH+nPmRj8pGHQBjxIR4qmiC5CrbaAgtKziDIQ+Ub5CGN1LftsKA56FngpU
rnRfmVPvRSkO4n2QzXE/BUCbfmYrRMQmqTZSjTwr59B1ih7Q5scrUtrysaJn
1vdbj5/xzULz5uhVaaLbsUF280t+NvXyM5s1XmvYSHYDxEiis2+1Z3+i86uH
m5ZcV8PnegkrPeGwpuK9R6qsHw7ANwWNFFcBaPGxWK1qdVKz96k00wnYCFkU
CiesaMajkYdlkSYYrnbS/syRjzpXpoKUnE/KaE0bFJ5El5qWRXndAFXCsS6D
8/CkHW6PI7NXyg8gaHJXYSfm/X+EWPgRtl/oNejB8cFxJSpVdIpWZQOtCnff
5nwE3Glk0xyiFtu/tWTvFQx5WiCZHOOYVEozk7iwvNLjH5MDuSkJjta/v6eP
IYHSiUprNdHDORuHQaHWFOvSqFZBaEqu/YK9CP7up8U/Rnca2tS9dsw8zBtN
BCHyYhsqxKmeETri0DZczN5FJxua8Azw6iTzmIlyx9GJbSQLc63AzOY5hgwY
bs2Ozy22YO6sGVNJJoxcrfiXRTCVxa0nh43aRRYH7nPPtbwq9WBZ4bdTj1Rf
QFzJJqdDIReBOM/gZ9+Id3GesOKKG4ZWUS0mQ+zNtI5GGTLYrg5xEDYywcid
r7irnJ1cC3SWptCBqOLcETw0QYzhRU2MMdai9l0a6zPF7V/s2KxNDNNxrMvb
Ta4XK6oDUAflQ/yIfX9CxWDzOUr2VrQf3BGj8Ny8F2mBuw/sOBJEB1+ap40G
8ozZ/DLudaWAlz5Tab1cAvtA1UBIj6EnS7bPtkV0OamGz9MCb58wyMbacwGp
TpUe4H7LLNXAJX8fgXnRiSo6bZ5NQssysTslLT1hyTvo3fVI8Deoz0n1qFef
JXhq4DFfDKCNVR0ZY4nuPZXzuMQ3A3BXcdR1Tul+FVrE6ci09Hl3MLlCq8zz
KgIhDVeq8/nM+Rq5O0HbgQLXI9QQh8J9A8UoOCSzlFuW2dNXossOLNYIelpF
tOIJvmC8v5deppfVhFAIB3/mydcy/N5GL2lruy1hqGmPdapVHe+bukxdZyGT
3Zucj2IsGRLuhxmjl1iRJQiDY02Yij00nKm77S+WaaWRl4Yw5nxQKyiBJT4P
lCYsv7TgP6/gVLAYcADF/YE0XOK74T79xpVBD8NK+0uj4G0ANWlc+kScoBOG
llypMFN9q5DStqPTe+0sAHCMRnVNwtr29SuM0Ejxgk0+9z4p7c5TI5bWbVAl
rDxByy3IDeHa/Q6ENufWwuCfJu6E+pgLWGHXxHgvxo8Shwbb7pcOHebaNWl9
0mJm+3zGnAiVh7BcfCF6RNsHggVr/Ru0XhqMFWd6oqyPWEEjt4unCVdrfPFH
a0VV6z0jaGn/QPxOEjyq6OrmlMECcR5G1owTvCkhQ6iYuwwAgt0EJ6ZZ0SEo
0VWlXqi7Y5c6ClKFzq8+8+m9HdGfFMc/2TrV+hETIKnYfP/OwKFgRpSfEWNy
TBM7beEaTI+Cimi6+jyddNL3KWljxyG0Q2Duq5sKIzTdBaLYQBGqmr1iCdUT
NmQ/9bMShqtcMKBa+uNR6aCoDAD0LXJoRveecTo5bpFHCZzAcmObvKpAER9x
SheGPQKK/ES63ikb99u+3r86SAezJGpPvjBFEt02/UcYn/RP5Zc3dEOPYtUL
4GGzSHB9lOPIy2eJk7msSjQTu+lA49+l25flquefe5Oaesxh7KWwZPCMqZvc
41stYxqFHpTC1yrzNKxxC//tf0xwBHnWCSDTCOgcIxUBs51UP8rryEviJx9N
lRrZ9VfEnmn8VCEDYbqPq6wQmhYUsle8+l73Rfj5R6IHiKjayLyJXU/+wo+2
CCnBXecamZXqyN/f+DRpj9rXGJct1tJQd/AbrlAEU3svMVNNbHjRoeDqXSWa
vtFHSfh8RmnKNQ/VZllp6M+T35f5T0HBLU4JHkXzcFGF30J4VoCjJbOSMOaC
rA4VarGaEHz+VEkEN6znKTamBYjcaFeDoNtCpZlQU/SKd/kUIMN49k5PWyry
KZCN3dufo3MK1X3rKYJBFRDe7RkykWoaqpz5iOUpCxxV1AhM4hikUPRGkt51
sU0llLryBlAyGvGHVqPZxX9eoT2SCVYyUCTrkroivEvKCzOPmMOxoZhyHpNA
X+QotPRAXdj7OeTwoT9CADnt43uHouNgRwVJvoLx3YR7L0IpeD/6hfl9yfFU
UriAqEfoiQ8BqIaYdcV/rhJ976K4pKHX3MQDyf6sBIFwhwb68u8qpECvrol+
vqdT1+UUSlJ4jjCs/KF7wwL4cL/zYdhMBIn7j/TAj/F4GxUlwUW5IV8hRKBr
I88BJ5DEPkLjbRiLALv9EGbUCIM2AtKNPqVIeSywpOKbdtZj9DkVCKnbSykl
PG6xk6LXMAZxC6f2KBkiTCjk3Sri7v7CHpUMUhrNEbur3635eMynIl7/JQYe
L5OF1a/JyF+SSsKiJds8JPRTPVGe56WcNfXrySVTr7PximNiWvXIXq4naqo+
oZRluZ1ito92D/KihRmDtlRWiWALiIyGKWToNz3fA+p3f3N+Y79uJEC4yiMA
A0mhW2LqMtFetEX50n8w+uw34qlZvmNIEfEBrlmiFSpXqBsXhMpM2pbKalpt
xhkd1IpbLxfdH8bELNCNb9kXaLZoG3mOos3ZYWlBKk2dnVFlb5466ER5r6XV
550cHpoHYYOoxJv8AlSrEYHRMEZCcxku3DgWtsxpQN+Lzt+lcmOuTcF2LsK0
ldaMqXOmjnHAH0Mo8c8oiAaOzKkL8hBF193U8ZkvFSfAIVfmUilAZQfphjai
skEMCc6E4S8BjTNOPGt/y2tiBhWHES14HsYLYDtZGt3Lk6HV8ytHity8bdQg
eGnv9Xqcj704rlRic0TRFnaIjL0bZ1m7a6UxWvsFqwURiRFieIN+heKOhSfT
A5KpwYY9wrfM8zhBOEHKjKmQazCjyX3iPhdi2FMeL0vWQW6GkGFnqCrs3Xt3
dN6YhKhY3mK2LUDbwmPmtTSBtsWEFKF7vhp6Qon5E5demr63DJ8u5REVQshZ
Xq9DFJgwROQ+/eCeeYSTltFtBElPwU9fvqGJ5n/DiSpqiS6NkAnHVFJL7HRd
8w08kHsBtqcoB0aaleWAh9xMfKSt9p7AZped36hrfjDxzkZqitAQxUT/FSSs
LxmH9REO58B+4Ir1IGuUU2UpQ0E8u6SFR/flc0uAjGex2C6S8cN9a7LWy7pL
EHdcWU3Nf5SzzXCzzcI3mkTFon5eUjjASHdD+r32CBvKJO+yxLo7jGgjDO7l
Duiu/gZPSWu/enTYMrYI0f2NpP8yJdceIKOY9DM51jf0e1kj7WCy2Y7YO6ji
iiGAoygXcNL/tyyqIfCUIJroQYYoRDCliSHa4ZqEurc6jhmg4ff5AC5mfRVV
+iry3UjHvF55a7RTOhTs24GMVRnPMtKnmH/T66rjKPeYz8p6T0fLvweOTBVF
ExGDQbFj59Zatajbj+OTmDweFdtkNZF2IvJLbBJWoGu+VwwxvCpBY0Gb3wXR
WvHKm9om/Z1BJFTUqPRlSVOVOtCRtf1+bgt+NOPh5Y4P/0OlPdTD4ahI/Yfl
rRTonazWlG/omotFHDBfWoDm0lwwj2nxbGuHejmtdyUXRV2RWDF7XoXukd4D
SO7gvN/HHSw0XJRm/UA0nQf+ZEraZG8XOq7hRMDWroPy0tuzfIrL5yI99wg7
AceyRprIKbCl5A93zcjiSWZHSDVcn0Pcm8qLQ2G9KVUm2/7BaACSIP9XlIZw
mpmepPT2jLoMZj5nl+BxzYy3aKx/g1U9FsF73Brf07gK7qhhtZ0gYyG9uuHx
VaLK05QQdTyxCnWST86R3TVuDc4b7dpy+9509Qogd4kKdOQgbAPMyQ7AtTmK
mu823bRTbv0g/0lnA93wacRRR2Yd8U1GjLrHZbv513nAamq5xKcVW0lCxHwD
ipnAiXUy3rlaLF1OB5fjtKx/vilIy9HoYC2Dftau3Lwbiv/M/r9UtiKyCWf4
od7QIfbjb4ySS4sUB+NKjsuvlDldxSJ/RutiInzL0e1hS1eZ/+W8TXOFILfu
1RQcEWJWWkvBXsK9hMm/grMETEbLDiXiYiCrogbP9Wm8YlyL12Ms/gcJKtFY
KsNlQRZo6oq+DI7vC7CchkI9OiTN2lMwR98pUbh6z6NuR4eMv6BlW6b4G0Aq
zgHSEcZKgo1VHJmNzSWP5Jx5uxVcFgXy5fiNFOFF2OSxrCHc5LijE8yEWrw4
r8e85RuLWFDQeSgUEkEij7CsBz+Av+NcaM78b3do+OkPSP2Im5575KjVHR3J
EuQI9ayx+0i1iN90uZjKyQcRVa2dgDCgqF3HIjFFy80a5k7sARSloHZCq0V0
V8inqZ31J2zWisM3rVmYRHKULJEdzsiFpZdi7gLPYgdbr8hMsQqpu9SImzTN
jRlRy2EU+IaOZ4MXBgu60qj78glqar44ygyXTg4nKFsRIXh4u8T6kGQtojzh
8Jx1tDDMB9tFjgUeAJYx+hpGDDJLsKePZwBURSCI3O+CwYnELiITlYBQ1FsG
Fk4tyGrECPUaehXZGCy6HNNbOA0O3jMh2xSRWGCXrsCx0uwoEalYvfKllqFi
1jt+4TOpHSgrEOCuAReGQybaDHF01sSxYlwPuNDAx/aL73PGqKsezuTzp2Cm
detCEQ2GUxWVYd2n8Rd9AE/EJsTEo5SpzV4ROe8xj2q9WUhm046QLHrZ6wFm
DcXmdW2vt0x02Ckv77R5azbYly6oaxi4pBC5feEYgfX8PIBVB0Jt2EtA8stl
cOHxonVUy9UxlW0NL8XfHd7VbsKGkJtPR9t9ol11KOfWNkjGxGDvDgv27ER2
SmFKxNonMjYrnYd3tmtjaJIiSyrPrOc19iPspCzMGnhWIZ4cwRn7bL2mgAcr
/fifgBRNSD9YLUKwMfKWDsEhmEP6etYOFF+JtujU6mDsmQrhuWUb0m9hVidy
V8zn2dFPE/trPJujPjsh6X27va33YLq1ukOTnzV20xEoNPP+Xd/m3HKgmHWc
bpl9tNAKYVAu6e9MZAgTiRMmPHQPa/5pCxAaDxpQGz6LOSpm5UhG1OoZdTZC
cJFp8k45BchJDUie1KKun2PGRsBnrahbkAZnmyn5tFxCHrJjw4QgGLxg0/7N
WkQdxz6vk77XrsZ183iX5rKqtPu/YioPgCgUql+CiLnB/VptVQ5Ei1J/Roi5
JphlxgZTI1rKyKHt4jr9cEhREOCvUk+2QKCLtIsqXVnHC0itcxSVniZs1+d8
pqEMb+bZQzZsrVFX9w2L6Z2zcTjIZZSmmnYinRfTCCFeBZSIhMEeg+fuRyiX
JVdfqmURExJUvWrjSIa//fm13SEM2YZjIjBU8FJ8BR/lBo8OqmqTy4AhDbVS
ngCKWPQ4JTJaVFG85HaUNqKQUc/k8uslcLr1pwdHG2eNY/6yr+BjW3X+WZRD
7cvzwzkTRod708rf0+xhRf9El02TaQiaxwHpX1bRKOqnrQiTINj0E+UvlyHN
jFFMD0gP+EIsS63RcadQo5aAXSrPnXW4hPzI4Fzg5m3+xKtUKd0LZ5NA0xjy
ZeQlk12JgcJnhalYG2C48tnU6VYI1SXg8yJLpMxIzh50Wok/Lj8qLpNsu7eN
eh4RrH3KIRlKPb5coQN82vx9SC5T36o/ZSH8biq45HMQs6EoZWNBXAnpfXc1
PHJtiONyx6tFCEzujfM/Q/h/BZXjSVd4U0NrYj4zEuBSpDzQ1KE0HZU7ihDs
YNcMbwvZrAPUgTyAuXl0mqTjyxuJ7MDqqmK9ZhDpV6ULx5b+Q8+s9T/6VPN/
2wbS7/BW5/GnTwfwZghNxvdKT/eqIpp4yPRDOufOBZ2XCMgW2EWtxgO1bcr4
cqRgwNrhp3Jf/S0W68XqCNQalqS1v5JNXp72iQkibekKUUYS6hkISBRihxam
g8kU3oc5Oo4q9zykJrhoAJ29+W90x3uzsiuIBvevCiv4QCGE5SUsvBYBHFqo
UxJAgD9UQPNo0EEyU/tVn3UmgNP99GkGDMmLmx01/7aE1lJHsSRZR/fOfY2P
T/ZW/wG4Ql3d+JAsZ2XluSgR895KF6eNpx3OM7cYFDPlqwKVVL6WiFGhXPeZ
YLT/+UzMzCbjluh9kq4XI7rhLWJVEKBWtdWhE9Fju6EBOOxJTkXk399bZuUD
VDQmNSgvZ6oXhhyi2DwztQ4N1bTUY4X429q8sEN+Lm77kZdNu/Qi/PTNiNrG
j1UdamyszDUtLxMHAAfTrnAnlxsEKZLupE0qmuXGCcukmIvg2Oedu7dez5Ri
ZOkw/8ThOEz74Ryji/OoFyd4gZWVwKFz6FKJ8kzhB0EwKpCG8si/4cUqhWnk
Y87ufCIHMz2dz4E/vG2/M9dgtBAex+hFLKtCHiN6zXw+7H5gx33Ysnlkyhrd
lDbTPAsfIa7/8Yi5tQjow6P61As5TnO7T8ZCo9OpLFuXNNGfy0T83gzEiA6o
HV7Znqazcrelgi+9zaYGf2R/6TjrKaL36fy92Byf3YA46ZCaRjhwM9UodRDL
WsC7GBMfD9sApcl+1p1+SHSSQivoMzRsB3SwKKUfWSLJzE7P27LVDOikDb+X
e0ni1AtyeE9SDN3pYgL7eTfDTHTnFxaEnlXcVt72sZulgepi7ren8ZaKEjjX
07DhiZEePGgcDnmiPeMeDibpQIjA7e2Rd1N2nK9SsjHc0g5oyTjEY6vr7bws
59skq0prj8xc78fq0grBH9sE5//oxL4Hmgfcj3VmreExvdUYgitFYNDLgAS9
3GeW8TJLs03cxkr8uWSPsT0D4WWq27f85r49AB5QkIPncxsA7NqlOAtq+AUG
aXZ+k3lgTyPT9tNgsqMlJgxPXSsDuwsDlSbcxBNu6G0rBYD06xRNS+F3jE2w
fOJiFtj5lchBIOWa4fWRcgVJ8PYEa6SxmpxKznPncRmW5lFjJoUqp5btiJAO
k9lqpTud66N51vz/p2Kf3pvk9GfFKOU8DOtE+9mYrxNO7k8FZ0JxlOk6G2IF
pZBJkcVq/aj+9hXL2UwttTuxjcBYt6FyIJ9jPzIoNYxpQxRZsws/kNVRoV/N
5lcfkUyslkHxl56bMoMOCOsmbt9XeSklF0ixG2MeLPZEq+lAmgBmrq9BotB8
L3Y1wCygFqnrp1uAMb/Ny/RRkyCgeCcazBKI/B4acVLzdXBJ7TwKX92t4CZl
Kb5PT52xcZUNnUEAkXItGd7hl+0wVXEjSxmmJ7C5E6h4ykd7nvCzFVfvT70s
d7tJwbWEJDo+lXBzP98fsT7VHAGavKgCOagEp4xcPS1ZNlq4dw6rnqPA6O7z
YQG4rAFxJkwGigbhyJF45eJFMJ0ZfeZD5P5f9JzeYfVTONwMIKbpORGEqkW0
QbaXCMhIIBrQ7waXpuHVrnQ1KvTZqR3W3tP8i9p6EgkFcXo36kwwca/doqJV
5OeP5L+WcLb1ty0tLDAQxclu7JLqJjfD9XIA45brXDdqFir77c3pi57LgKpp
nZxjzbkNx3tWMfDMcP/ywcO05dWInX65EJQ952ZfsJbN8PJ+1gmtBi7mzIAS
tK9GU9OujvJVj/nPKk/73RvnBYZHhYuAj7kkDuK3+dUHZ73n69I8u6hQ0DhS
8+piSeG7HaQXGk7saLGTJWm9JgPDaQ73w6huA+EjxaMi5q66/9uBJFbMGRz0
K3HNHohIljqvvQINZlQBxvqbhjdO9/UJJlY8VX5yiQr9YymF5buBVNA/pC24
kzjGVMcrbNwMF6yzfljekrie5+mpPcpJoerihCCEfiZ7Tc7d92fWHnKwNmG4
qrZgcn/UwSlinYbrrjxWEXkFF1zc5lUocD6tcU4rs8rpeg7UC3qsU13riRNT
duaqcIeC/YIKaotk2on0w+H+8fYQJcP3CvX4Zqv+pHixXes86yqEDU4WXasY
ZsOsxcFEC2aLTHCkIEJn/iDUzI8n8FQXaxCh9ecqaDymgmJ0ICbnqtuwGFzf
qbDlErhzJ8CG6y8uY4uAFd2YmpC/swRluz86mBhikCYvtfrvTp7IOmjjZK+p
ZgkytzT1VhGCMzXTcZkYON5QBgKGFEyp3oeOuhjm5AdTps2K0WNZ+CUZSyG/
3XG3GOm/bzZnwqWdWt7Ypv/dXR667gxfsis2X8jNtO7Ue1lot1AZX2fZVmWg
on7PV5ErUDmWiVcNw+v4vbKPlxMAmwgB+8xImNogorVEkrc4BYYtzr851Ag+
7PxIj2oCaHGBSf4MySiS3KRZKLX+QYqzdTqdEYPO/E/JC33briL4t3bIhRkk
5IzDes8yX9kVo85sPe3IzAxSFhylcALP9TA4vHJeGPQ5Cl4Jh/67JA5jAh6U
cnr8hXD987mdJTWpL8CugBVJgsbmXEQVkxdTfPWb9J6VLOt8U/z21yPK4QBs
ElTp/3JJDPpurtJtbd43Bi6B99nVuBWtfXSV0ExI+BorDaoOyWfw4EHf1P4q
Kb3foYmLIOTFUmz3sMM+Z0pGWd6pV/ent0VajeiAODjUivGWUsNAcTUkBjCU
eRiv/KHoQdEhgUtVue0DfRhY7eSLa3TE460N0REcXVjl6pMkKiNcCP+Z3WCl
0XeWnwSwIwIN9wltcPMFSo7tmNqcE2zys6Cjhe27wizBr+sVVIfd1IGSEVvP
KKKp99Z95xIf7geapLXlMf5gHh5v5by+hB46vkghmEKUrDtW0UTCESEOCCgV
QSV91Gq3eSoUGpszUwnJhEBGnfJRLoDRxVwEIE3J6CIFDOY0ZU3RWUosxeUI
K6ZgIZy0Q4U7oGPnTOf15iLcFgccqE206KcB+Nupx5XLRVrq33vhtT39skHf
4mhi7zUc6UkrNBBMcW6L9CFgyhSrUyyFOpNcqAu8tYJzVPt1v2DCdz4Y310g
adU+N+9In0WsQQWS7PXmEvFpscB4p+Pus0+8zUSoFVjZcvu7E5ebIoRpcuzC
demtsF8wLH2VcjfQH+GGqTecqMQCroSprzDpBUezLsbZyOrTuNWd+r/wWDrg
OUi4E/BR0eRhKjdoRbfQDLlUQ69xBmWyrLFwrRW52qyC2WbeHMo5LeYuQC79
zp/pU6aQepqTDH5lxzxXwa6aH/C/cz8Y5EXTVlXwPgyPIU7xPJyBa/NDMbVI
s3ROJI3/hAhlKhz0/VpirdfTNflYfksmjtEMfecqKytr70ou1TPaE1yZiIkx
eLRpqbL8DdErq1G3XNtTDrfyd/aoVXH89VXjSQYZKTFG5NRV4dqkFi9ImkOo
H5vmzsopAFDXrNLjK0+jenyKGeZ1Y/66gJPHjGmTLXgL2E7aQ8/LFZLQHvre
moLiLDwWxRMnKMh3btXrxAThuEeVYv/giQGkri+cL+iXgywPjdoSxoR9/IdL
6bRfl8vUhIsBDqzbhn3T8nlm/EhIsBe1tY1M5ukOAx5acQf3yWYUX2rlxqK2
L7Y0ysd8iuDvgGlEr0niYWwqgLCEdSTmFczCOxGz6Tlpp1Ni32rsEWQFEDK/
W3bd1aVU8LOYIvcvNci4M/x0xPYcj236uAQnSezuf1pqHdZPzclgB6k9CPJB
OoutnTHtS8E354fxnHxrmrUX6keKgktpfY7wLk7+ZuPo7VSZExmPufzjjLWd
yCw8hGSZBWMJ7YVSv1mACI5/IMKX5IVnOwZNqle9tZFld/KFisYUt9x0Fmqi
INcEMmmqssacuW1MCzpwRqCwK0sHFST3ouyFjhzK9uYpvdxFdaSE9EtUIEx5
F0kUKq0jphs5Gqgf6+1lRU3nY5pADZ8zsYMP134B5nRp3uQXKccqDabBKZkU
bm5I+zf9xwWlfzQdet3Eea6r8HsaHzdiBgjDmc8vGwNuoEy4STKO+gLYb9/j
j9iqaLbdSxzJKehJbVba1KGWyryNHKIqsfJwpHRIABuBXu0hzBs6XX9FVrQr
i0j5EKLBK1ozHKZkjxGI/EQEjV5XN9Yaa2l32bnH969kKrDmYkBw3nVVaeQI
cgiTJOCg4Lqr4o0lzFhsM/SL99n6WObHqiP+Tky3NMqEi7h5lEp8dGHhhvPp
wdf/mLpbyriKdM//4LBwViQMsrJZUQJlbVVNTSsU4YtpiSxmi5cidrp+4N16
lNm6apjl+YxhrD+pqmh+8Bc/ob5XQja/t5K4GjZdYd/oeeHHXbX158RqxEU3
T0UX+Juj9Tv85USPFsWfTWjQzLhoF13SK46IrIxPFbfNBJZOB6IQnzXLpi+t
uyQSG/nHuNVTa7dylu7WCQT+AHKhZ8i0+xEu0vEzbGXGX4Io6sePzKOXCK6j
OX0GMCJH4Iw+TJlZ6bPKl8wWOVaqm689Mkhp9LcLqmwInJ001fmXsV7BxNIQ
1IuPtWXqDz8Hcl3i3N9LCHk0NAA1YkTpSNqVejDilWjLILd6eVOnw/5tjGbh
ogP/sn+yN+dxZczENbUAYRMV992uVAVSpVGMlW4MBlLRUfaPN4XsOjL4fSpt
kjgrRdic4IHUrvOb+k+suRusTQSjC5TzYfyIisEBUOTas1sLwks1XtrzdbcR
HTW5zsPjP4QNG4CYrm2jR1o/4NF7ADOgruYB2eTy9XyQbIIYuYXpEvf5RSRi
Hu/r3OoCdcpRr6qx24SEWCXEqYkOCkyqfV6KCIY9GC2uM+cy5egJTsgdv02t
imWEK5bDMzOxEBE5GFzgaYfAhOgQb3FlKyf+aZy8J2GMhPusyG3ZBfDIpHbZ
zmvDE2aUfV8Ki9BMog7ubFniyR48OFPl0zcqLs8Bt+SQ+QAP8T25umQY4dNC
tm6ea8uzBwqM32N1H6neaNFzTIX4V4SOjKO8QMTQBR6SuX4uSQuF6kc9maWB
C9NF+GBkgLwp8NRVwH49vrXp6bJYbOpw69DgfWhJCjnbLY4XAxmzkkwoFb1q
d8A4hDr35rvAu0f6+aHgtBqNiIXk7Tx/0zqLyLOtoWBo5Vl29KfbVWyg7+m4
63gJ5nypMrmi4gRKLZM0Q/Hqw43a3IOlOsLvq71BElPMF+EQ+tBfC+7+9cmq
tSRmaJj+WfUtCXbF55uCLYvG1wm0kq9nIpaZWoX+cGAQmyoZewVobaK7v6/L
s7TbXQ8zao9sBcU2T7AZfPJGFUKXAzXrEeu9+bU3xA0OPYd5Emr/3s7Jtawu
CaXmUx5QcjqLCQW5T6Mj6VOu+noIJwZTkW9/zN26OHJrdFlvJbNfLkdDbGDz
SXQNX4rNWKWrnA+0+50t/hN1uF6BFNOhKBuar2qB2gRjZ2oN4YbemSoMAMHq
JcwolHvZBUC9cp1/geYYC+yNlCDhsbeqv+HdocAJN+Ac3/jD4EL+rl1vbTqv
Vi8E6nk0gjOfLtFarLHoHfXh/a1d+tGzS1MLQwhI/gF1veB2KCg4RTDvFsG1
nSZKPRD058JH9b/GtjPa/roi6c1tF67by2iuyQhk/56ddkdu70bJHBmTJ15V
O7L5WeE0hZe5cJdx4tMSxpTCy0RGDGhpv1sNrLhDtEwiDH6eY4n9RMxi73Zm
H1uq0vs5non3glb96lUTNoaAJweTW4XRmjz37owKIhSS0Y6Kp4QC4z7JtCZe
qBsAVzbQs1/E10lqUcgCF+MuHQkmBa0gM9wWC4dwMQL8rFBQianwxLFT/0Pc
Riu3kbcFfyfg81mRFyRCGfPht3UbejKvJsY/AxI/Cs3+SFlc8krtCbAYY98L
DGFbhjgylwvprShIu20Evxkyp91euJp7qy8ogGGAAnySPJHOmE2F99oHUOIz
iqKIt/FB92wPjNT1LnEaxQD6Li1rMzZtxp0vo08HZG7XmY/h9JQhnxa1RFQr
JwMNBgwcrzw0n3/mjdD5I8KT5Yw7ZCD3IvEt0jsFsEFoF0pVvBdLFHZKqO7K
FFlRTQJwxgNVjGNSyp0BsL2vJYpaT48Xf/Bm4EGQR6r9eFKQvfr4WrqMNiq/
z6vADd4wae4r/ZsNIZnVp6F/opJeoMsNmOYtAUDiWzyMN9f6XjZliI64Zpoh
CLr9rAUdHypMhIqE4oQ6OnOsg7R6WaiONoei7FipcEsjVZbKPCxgX1O4zbAP
ICEbmtJD77zqIpWERX1XcPU7n17hkus2inKDTByIo3so7ALLyBiuBY6serLs
SPnQ/jw2gXrEt5i7780z4gVemnuPsYTM4XoLHmm7J/TAS62Z3G4WPb4rCa/Y
oj/XQmL43qSa6RMRdjig1xZsWsJ2EkxKtxn43Hj967E+uJiqSCK2mUfFFKGu
YwEStFUEdPDBWJd9nhwgqhuH0YRuguZaQXK0VRHab9CEWRnPIz5SJIvHRlb7
MXtTTwgVEZCavhexpeU1VZPGdUG3ooOzHY43vK7N0liLzChxGVdcgeIaHIR7
aKi8/RfaWInXLL8mVDi8WKKHWCmnCaRcGUY20k7vuATwuHX2DZgdfq2satqL
316z4Yy3+Pg4Mak95rgy5hMUxjAYVnLoiaw4SYwi+LlMSBeXy+l5mNrMN66E
Tm/UnM7CW+gVv+lOWl1GgycqjfH538zK6DzjdaOKtX8me9VERcibxq60BfCq
XKV1GvZOIj8kQvfKGa977Vn5ZMfKCZfTChlCierDlO+VYrHaMmctASiuK7sF
Z85Z5W+RUINa6YcZfS00A9eDBFJrHVuPxuBsIawsbQHAH/HZduFDtkLIDCqG
NJvunZNzDmQTlSA0OQuasMbYBL8SJKT5VgAnfe1nbRd/3Tgl1svuuYhpnyJ8
fi4cibPCAdpKcFACkLvt3nU7tQrZj6u9Hatgbub6EosiwC6GF4LIEi1+0Qmc
VhSemNQpIFPysKIaYVgYk7tfBaVvYVeeRoK+pXQJ4GADzPXGdE+NQGmWA+PK
3IUaD6u/85wQplEsP2wEyhVc958N+1EgQ4esTMTwOHN0vDDHFLUFF03n8p1L
RF4y1isvxat+ROxR6ohXwuqoWeNWf4a+xXQPq1qahBAIjOTPE7Uhh31lO8ll
YVDilUhc1/8irwKUlWgro24gVV4T4DeTrrABEJfcggiZpzGsk9MgnnyalPwB
OihhGWRXgAfP7cmvNfPzbsUxn5R9/+u5P2gx0HveNqGdOR0Bfv1tubNZBGA7
lHnKjkHDPqtUpOUVCUuTkLiSLCSZvxhvd6cJppaCh+u7hpPT9E5CJYDH7e7g
A4W3rLlksm52h2rWXbDr2qhS1m8WAt+jFa2R4Zmr5IzZxpOjtGhPrbZkuArk
vQUrjf0wTX3Lv1tQTX6ZwvRk5eFVfEkPFTQ9tOrw0a3SSN0HeSFOBqn1lbmt
QI3PJ3h5o+1V1on+AT5ii6fEOhAX+rXqYSEEHcutYgM823ouBnGLaPGbkwB8
FuhISNJYzm6fXOu1sUaylXTwxZGQgLqEKc2g781x1M3fmEOXgXBfZdmB/Yec
ijSHnZ2XiocLNk8vAuvzFjEkBqGAiBvs/8gkqhfBy+K5vWX/UuQPwQnEulnE
u23H1wOnEql9R9Z/m8ydaP6FZNmLUu8/zfdLruMG/+tCIf/el2+b0OJIA8sB
gKzTjj9JNDFwBzyB0Eosl7dSuQQR3TbtHTFqhzl5sfg4wHqHg+fXEPfzUvaT
H7DQxh4nE0c25VC3Rye8ppbbrzgoyWbMaLof2uvPOQS53rtxjo1sBtHnhMkq
lbaadOS1f69DJU1aqDc27o0yct6RK8rzgSCQVfthjexmhKKF5TGMSGd3Ijvi
dRNr9jYeRoPMZon7Q2zuYpS2OTGVS+E/O1RVXl6QJ6e1eIoqoDkdFgjTubin
RJrE0mEtyT2WjJJW09+TJt6h4W9NWItnCSDnQN4WioNWDa7DyQfjg/gRc/Kh
zH4Nl1G7CawwXYLl4lm2N8jxcpZ9wKJC3xIfFVeAbdrLZz2eGVIQr1STuF+B
vXRQrhkfKL6gCBz5yKUFJXar7h8mSb/rAgkbBGAjrlZCPccXgLgzNooRPwQF
lqCuZgKezy8GTPkqI2eH4NLNl+l7jHk+CxQK09uAzzXox133WmZLWCX5GaKe
PNvWBSEkAsfnwzFp3Odb34c0/YOn1q/apWWAvu6nkI4TelDl1vdwLrk2PoU1
EloTSi2ZUlJkP3BFn7+jTkHNo1OUkQDPgZXNkd8CLX8dIktuTfskPc3wjP88
gC6yHs2fkiEQTs2hzI7CS+5TZaAnldIUS6Qy2bAgxukJtQb5dSSlcB/rYjn/
hS/8L6CAvd/umL97H1Qz6F9BS5xjLgIgO16aDh4ZPe9vPSyl9YRVPrZU7nQF
SHkJqGeh9o/waPBczeXZuwsUNHWon2ollzMkZtOY+WY6XOsSeRxV1UqiNoOs
EyGW5JO2dfn8SwqF5TTx2BNYOdcrsglTPgk2Plr8B28Vr/bAQlekgWUOmDpb
5oo7kNi/a8IUdK0EQONbtmGOKOqZq6ku71bPUdHOsCi1czTiGAJ8qqtTH1ZR
hK4nbiIVcy5Q7u8IhvC5OKv1zb2Era9GZrcwjuYt9lAt/rFF+mmRtblGN3Ka
TGJ10MdQ09BtEzmjQcEq+9o2niv8FLJOEfLUFWAQtL94/LP2FEqg6dTI7YRj
ksDhGdpQ8eMJeO+5mOMIqwVISKoBnYxkam1YjgxCiMQ9u6ucljwgIAkEIh+N
GJrZ4Y8XPv4PsROm/Vcoz+SDJGXVtrt70JUYxK69ZksPKA2WAvV7POCfDlLu
qwF97RVLMDW6gXVgoVfLcwKfz4A0YttmqzUBShMPUfDXRDEn9lz6+oju/dLm
inDFhZtI/3i1Sb0ASz6GEKPv0TG2Db9ttCEFF9dfMGWmm4d6hMwDmDMg15nZ
SrKPm5EYbmGFyVJCFw4TnSZaAG3DEIHy4OlYELeZqvij/CgyKYTzAWPOgjOg
uVtkJx3Vtc9vDhyj1yI+77KOBCGzgBDq6EC7lAOA9oKGmhsclu+IcnHqF+Lp
BXO9c19BUy8MnilanD/GCpWoJ9g+r71D9PwsULqDLqChGRMe9n4VBSf1M5lQ
Vqmn0c3FC9ktHkx4EqPeyuOvOHdQeWFZ9m3RGvo/wn0Huh5U1iM6JDlRgm6G
QP0cvI7FGbS3FNChW/Ioc62pajAq76naKbQbm0fJcwmznusBe8bBYMJs2OUI
l9YdYqqP7w5yUJ0zs09d15fsKy6vrL89yz3r/NKqsBT9D1wp6RYErbMBSSsy
5lsFc/Fw5UJ7cV4cAqWJrDVT0BcgSZVKcATgk0sI2VLnNQSSaAj4hUIT1c/Y
Qi+JPzlVAMKCzhqnyVnx2IF5wJ+H5qApCjle3JRuGlppaccplcrOLbNSTVi5
UEg10WulgvRH38GOXYqGQDQ9CBfdXgD9Du4OlAYeLs8IZHSPG22qWZU9qqFs
bOiP4uLix2+VQ77Op2uiN8OKXBEhzP9JH8gvtn2I8xAGg7Htwjckz3IfCZsP
STuZ3kH9XkM0l+t20JjdYQVlpzL1JcCoX/VimrvJQSvGjtAn98orov1TWUgM
PZyzzUHmHIUEhbvWQQQgV2QKk24A34078/Pv+GKXFoQV7vJdi6ZVArpVxJCl
TNeviFgazlYoQbpV+bS3n4fN0YeeVH870rQP5o9GIzFgfZ+tezPn/GbagRAN
XQI82FBOa3/poykCbsUdldrBlX/NIrV/c9BNMFQ7I80pLtXCoQrkfxhmxahs
/GLJSvJey9v10I8RgMySM3LhLrSlTXDEyn7LdnxAwiElMKq2i1KvHz1T4Gn8
Cj187Iv9MB6TlpGHmxeq0H2N+I/LS5rPqNtAHdFsdYHVXujrYp8F8J3iM7sp
v1TnwoN4ETYw3IDhxp3esnH6Mm4JnatzfGEYMTIROEB5F0moxr8LZm2Q6j7B
Z/LLxHu/g9CQDewrJ1on3GKPpqPxwbW90xhjL3o1Z/lXf9lkgBE0eSNOYLHU
unkJWct4aptvz0Vkk8WyJWeTT8UeOBfMFiBdyHvmzDD+xeNIN8mQyNrFrsvK
DfgLpFQEzKr3+auMzUUwX8fKpPinTwg0XMQdmnxtsNFCvxYF5I7RzjxwP/DW
D0a2cFDRA+m0yJSKo05DSIWQmHGS11Znf/IztnWnSQKJytKD+inBECJJxswU
933EiRt2r5WLA41q5Qd+sbSHw5iHCdDLUeds0vJFegYJm3qTyCpIVNcBYwIU
3TXaW9Rr5eEYT2TURX9KEEmbN9yuI2EnOLAgSvV5y2ueWZpVw9QvOZlwUIsP
OH0vywbONaTPtmWB0wDOB6I+4VEVAW9OkQj2vYSr32QpcRWnFFlSCTWzE0XO
KLSonSliTdB296G6ou8N/a7trd87v2JcVYYhKfz3VEVhvnD/63TtPWEGnWlH
2x/d1Hz4haw0LAM6yTs3hTQpPUckP1JOoOOy4fR7ogAK0kWmFWXtUoDXcl4r
URbtxNuBuVvUiaRy6AgwgP63gEA7JpanY1OGAr1tMxaG/b/2cWZaipMlSkya
eZtV447IYRnrzYFLfdvJckGE3bmuKUzOLtw60a6qODtnrvObBmSqYH8zJoYP
5svDHG5EbBVhYOfIW2zrZ9T+SN5L+1sErSPNVwTUVfsuoL1ZyOFciqCVfxio
F6pyXsoI+8xw9gDsNVFh2MsUGwFLHIIOtjA/rZw6oS35gCfZ3z47ePrhvJii
rzSjtlU9jwyxi2Ak8Jgvb/sq5lil2Hz+9GPE9xjUMaCIOZIFcAuXuDotfiYf
cZ/oTcZjSLIk+a0/7/b9/8gdjwPb5gqdwErCFdFHM5XQDNVylhFZWyzbMaWd
8niSm83dSmB6jYQDDjFn1desEuDc8feE0q+FlYK56Wf2FDdXsWeB4HhluWJm
PIpU10VRKiOU00bcHD74Sz5UloYnahNZsEiG+GOKw1d7eMkZxVOdpfKFkhPA
NQxia230oxm0xBicS2DA0NLCUBXBi1LaMIoBJuZbR6ca7U8ptpMQjLkzQnr5
HDwprzhZNYeXPE2luP4neZsP+hcCB0M9ozrBxlUePq7fjPycVRIKzrhpwaYD
FBYKGHvIKMoxyAU6qOpQS0WrGwO7GSdUaRf3JlCN/frd3WFWo1fig+ywxXEn
vgdxf+6LLt9tbK9veJvm3xW/FclNlkZv7Udf4Y7d8sLSvTgR8DFe12oVJxmU
VcAetZ35sidgKX0MPjFMP45Xhl4bxq0VinncpyzqB+igTT6bC4Bs9BNR5tqC
gsW4fG7QNFGyP6dgkVsT3MjmEuwuQtjjSMgTLt5RLZ1ktcjkGkErR/i4oEA9
QWdXsXZE70ZSiRAxzGbWoRx/63vm0ifRPLFzoPvH4gnCz535miAJ7tfurOlC
+1PTtrE9Phy3LAFXew6njI4HGTr1g3g+Ft5jwaR0mElwAEA3PVvXLvhuuXfL
iVOf9npN5mTh97kIqPV58mUEGlpBigPsX3g0osYDyLhbzOBegG9N8cZ8EEes
igPkVmpkzrq254679OQvmKT8y1RsxTotLE0bW0H1e8Pqz87Q150J6nq6aOUR
GdoUU3bpU8ZYK9dIF9CyQJVqTyx5LGwaW3IZypF/S+AfZP9U30ulNgHq2XeA
MQhYKeklCZF4QlXVJFy7ZnYyZPpbdA1dKZJGTc/be5yw+S9oZgyBhb1DoMeL
28D1w/Fuil8VB+gLgOa75Z7E0qAJW0WzHxviG8kthi4ZnslyCjn1W2+DzC9p
4Td1cphIJCjaQk7PzPHhe4FPwvZIK5+poigVk4VIXWIJ4rEC9OoV7Op10ZDD
wPlsSCtEg8Q2/qyLYHwrDu+u6xTLfJyYfr1quubxvt/1TFGU2osmLnqqbWHP
ovJmCYzk/9x9Zk81Jipd9WRQVvkCRksIGPxRPL7pd9zs9OtciPKlaZzP3qt2
PUKBSyysYPTDAaT+9Ts40ikEpv1NB1VZV/f3/h8V4P0Dk1swauvOfUZml4vM
48ymle1gzQZkVjr7ggpzr6E1tsorJKnjKvsGrjajwZiHeYSM34QTg0szggMc
J+kU4UQyuRlLgIeiGqCXicSPXr0lLPrrVRnQk5jDVJdsFrHqWX16emv3SN+U
Hi44mRKpL7Kva6j7pnemguBSp3OWRpjppRvsCNtu0yJbGqAq5EEdSVPimlDC
Fr5rRiTVyUzZ6WhOdNP0Qz4EZE1t1N0JWHWmMHlRX7owd0AkitasjQM/8sVU
UKQrM6eWp/bs5YJitBLb2oqyJTqDupOwfuBrpsQp3FoZx71zmMzkYgBwvBVl
1mJhTlT/ziGq2NEvyJvpaFfksT7BkU8jXmy/ph5yczFkcCr3UvGTCaKTszjL
Hv/mK3Z9psKUur0aUjFQS3oYXlA7zD4Z5FQmgiUt5Byymkv6V7InpsatV91P
UHAXqMwyUVERRwlcj+mVqdy77wRDz4i3pXfavcNev1sHSvo30eGjeU+Acb77
zDDkxoiK2VhK2sFUHU2aSxLbXnqX8pahCdA77eSAQk4ViZQRIftniizcnNw6
eMAP67kuniO+rniaR0UvBpKS98tNetuFdYMFQIcvkeG3fJv3nyt7AXFylAvt
WypCrAfQidGwie7IT/dD02ziSTdFAv9zaIE0nRj+7IOsi5QabGXXeWGHRQPd
BNC0C+aYWlYlYH5jhTYhh/BY/KHjSHV9USE5Yy9UFpWJpIzRO3cQv2HVK81t
uXcpWJDivx2RlHL/VazaTv6J1pyu7LJnkRWQwoOuWvdiQ1v8dpUBtAynac/P
ostM3UF9shR2CwXLEDQvs9helsdVEXPQPa8ijP46VW/1vt+Jg+RjG0T3bQbX
VldOWfXCr16zuYK6+mxamtHfBn+aSnyTnpNqMCawzVRy6OnwErD7Z5WmVV+Q
in3WI6rf/HwXSE2ye+7Boba5pyuRqFr+POaI7tAlpZjqxeHEZC5i6qm9ngwj
n8zGgtVI02YFfDtud/ODxOWw7jLvY8HPEMLUmpm6mMXbNML7hooJXq38mDuI
68mf70khztR1BZ6ZrNagG4ZlYUm1AjPxQTZoJBEE5uyCSQrR7Qera/HJ3pOE
eAdtgJtjskW47WEuLW/yX0PgLx4fZmfaMYqyFz1OsTB459fl15CffkgbDo1j
BGCz2nHlICaRwyNiPfYwlHCL2xTpccmS/hVajw1zD7ezNkXMvN9YxEE8nilK
IXNVpWD5Uor1gIA0ms/ootg9NTzog57C9F53aUztpdJeTHUYA/rgrhyMTngm
wn1foBSeK7q2Dntaj8HCsuEJS0A10Ewtkkfs/LK0DnzTGgT1de76poO6qM9h
okRTsWU6CruJk8N2nAA5ugLqQz3Lp0k7nXyQzOnQ4L3D8pn1MxBQRU9Wwd1C
LuApms1AroTcV2NeFHHNa9fs60Qz21TKZbSaI8/RnMA82XbqYiAPM6bWRG1c
AEdlCwPoqE28azN7SHH/AaWGAe5fssJxbgiovH3lSTs92ONpJj7hWImyff2i
CXhNlhVDs7xszwMHfAFmTq8iX6YtaoxKxtolD6QLthZl5/q3mTjOHMSNGv5y
fF9Ux3AMdJcrye6hzws2i6TEE2K0VWY6WzJQtvi2LbO6a2MirYwfGJHhleEQ
zLnKrgYKU9DATeEO3NUG5PjgDZx36XJnekJgMhBA5+2+9FyD1aa0RIiYlW0w
+G61C75qWfvhBU1xGdNei++JusUSKw7ZLQElmaBrV5awwqQu9VtKScdegc4A
bQBrduvwhwKoBCIMPIfTGI9BNA6S54mknRUrn9IiYQ8xP0khvDmIucq47Uqp
txX5fEzX7i6N7SiZbvr4+Y7BBscYuk/KosiZHv92FhX7pSuSNw+mfJWfnHkp
/fTEVoBWhbUOLgB8mdcZrIi8g73HSRy3AOmboMQqQXw32nhMYHsP0+/QiVUG
60fbQcW8tcbMWuF5cyxvHOQ6QiT7e5vUhRsrsr0zKVxZZVgyk6OTUpxeI/N5
If8QrQEYGNR5oGOpi8ZJKvIYMYNsLV63XntddGVnXyxEeF+kHf/0/1psOeGS
r5I2tnnpTNvg+wI50noLinPerRrQ3t+AHNStAkAAWc+llxF3FY61BYTKi72d
a4Y+qmc7h4wR+LXlFpaNUjH1KsMlOH3UeXmsghFRJqbSDIzlWY2xUysvvrxl
hZJVoqAFhJ7L7k0tJlCiz6zi+NYvddBtuDvhsMVKzMTSNYne+4kLsf9qfT0K
cM7kGW6VEbrqy9HaUTWymdUwuAxixrs7QVvnFFQb4gv7b8k2SNbX9QUWSnhX
cHLi30ZKGb0G5IE0I0XAVk5zzzEIoai+o+4aiY7IXCL4SDpCHERzEfxSEs1H
6T3RQXGmSTWjQkVSFieZByPVvihq3vsJVsJct2Q6EvF9mFrWZkgmXokju3+1
QIBFl7uE6Ogke4gjjbrOcefUG1BdsMFpZRozVZ7sYXKcs3fBK+dblELYW9XQ
jWpQGZM5Z+XvjeZCdjbm1yo5UQ2TyoeowbaHH7w8HYVM3nRQdAlPEf3+dmoJ
do6+XF4h6i8V9WOafJtRwc9612xrE8QvZmHqofcson1dPVaF6Y7xLqZwVODV
oUuNpAXc5PUgJczgoJ40l5GxzfqSqPizoN7NEzb7g+ShpB2ZIPxgI9Y5kAhT
Huxv32Cb0IA3gn2vo8mtf8k93Frtex5zux/x/e2btwTZb6C6Gvs6mk2Hof4z
5UeMpwjJ4lrWs+YpbpE8U2NkfEgvjPmNzO6IMu5jbjmzIm4C6Ms3Qu9UsX+7
/bU56D8Feo552X3ZMufjSiRi+kdJcWr+n1bS9oRxRwGFY+Q3xtZkyqJ4JHu9
apnwhRy0mni8M4MpBs4kbM0FFt4bvlqaa6xOSxo6ufBCW956TuKRO/NDMhDV
ejhV9/g34sAIW9lOVuhxcnUqfiEPfVr0iYk58wCqUwK9KPEPFn1sAQSEntbA
Bq8rrzqDmbz+zocVI0mjux1qDPMKQ+4s5J969DmrZned0qiygMwO1jVd/bgs
ZVL4ore3L7xqSMSwJOml1ejChYQLc0zOk/MbFkjTIzOTNdYAXQ7JYk/SuK12
H36sXeEv8IGAdOBYt1ZJ9Ajm0YtdgaKxeE3fIDeIAXibq28eFsOLC0EGI3vp
8eOXpIVBT1VqIjjmfgxjjMHp2O+FAY0BxBe5DLcV9ftYLjcVZnD4Z4ufqFws
5R5VDzO390iuleWKFP+6MOPL2XX/7d5yrSSZsGc3urXBEg6mM8MK93TknvRy
P+XADedeS7/kvloiifthSDiU1us8NG3v+n0XDpRI/PGPJTPnUJRbDzcpQAFi
wvDerapwUBJOOW3SxSxhvdzrRFMjp0RX5vUyxC6kQt2u+dYFw0TKgUlPjhkC
ycnhlItckAzMitKplWY01iM2HTE+KzjziM8Rfdm00wXPiGsYryWYerBgJhiW
cIYK7ZNeFBStBgHl773g8C0vY1nYS1Jef6tgfnAzyOq8oQORt3CMEWm4FcrR
ysSdT9+JmSrRJchQhNQrB5RRA370eAgV+WSS/qyU+hwIWqIpZYgjVENnDHdc
uhOey9B02/4vdzCgnQ14emYjVd0LnzFiNccgNE0IlbpRBrHRSRmvY5UlXOrE
MJIA6NDaY1oSzp9LG3HDigeAwVhHaKBaNJqUXOfG2tmi4R9qUSR0w79VGaaV
wOMbIM2+njAwlTIsxiMEQ/T3TCx6arsLwZCjt7QDSpk3MsvcnNIxH3L9kITK
Vtx/Nf/EwiOjBBJUja55dkE3wJC9cFug886Bk2fRf7VTw5KlSfmOucRAvZ9+
ITJ6ZcZ8nAhDNfrAstd7BKv58S0tli83NY7hqRLquFzxjleHY38M6zbpdSKh
rC3UrsD//ri4AvF1Y9jqgWiLsUKaVgGmg1TWfCPVsyR0/5xhkUuH3Z13J9Lk
/wJVH7WGsIwsa/bbKUF114Uma6/Qz61oW/HDHVYj/lN2at2tlTL3srHAexak
jmFBQsKbkZl4YbgVPrdZ6htN/yAxHoWk2C7xsSWnpTK1Zs0W7tbgo0UBcWFE
akOxE3xwUZWcktfj1mYdpWFuizdLVtEMVDmSRHsJBiDKiLYJ97DagUhe5TF+
qAc/Ge2XiNl6x/pgnMZY2HXLO6hvSCCGSW903XlKmhd/5NDCMLV6pzCxwSvW
4diOf7Eu4dXNTOhih+uFwaaQYyWUc81uQEfL6q8SmeSmyH4qIbn4fSON9Et0
5xgl5rN4sUDdgvIiO+y5zC8p+3ItHowC8ZC9Dq6DgA9VN75A+pCoFp8FdbxE
2lzLox5wZJ9AbiJA7NFh9OjrWGEHFbJpcIF1O5TWI6C/axizDinv3S2Af1lF
mwOWLnqfsbnI3i9SdczgKZlKeIh3O0s6tR6LM/FUjrG7IxXXhTR0hjcE1/DA
E4xsfx/XUphm10fIQhJQ96brajpoowVsBvUit5vCic5d4nZriaudwFHFUdj2
arxt3TMM6aOeZPpmJzefWN2UzwDSw3Z0sgWOtkX89pYd0bbyRl4qFT4sp/sp
yPOxK9gbHMZEAV0G72it6xqVKJE8p7h7joeR6z3Y4kHaSDllO/5fmpRS6nT6
sbxCu4vi4F/jgTmSRc82z2hndxsE+r2w//mgVvGT/gYjBpJS1AQddnFNZs+8
qj5lKPkXebEoIZCO7X5bbKJi3zqLawV9ZRuXOxDpWY5IiNSrkUXk1NIn4l+E
+5CbV2rrOomrbJ/gxA2N8TS1KrCIspogbr0WWk7mLKUcLiyZGfnrnXgBRDfl
Eq26RP/cU/aBoD9MAwL4y8aoYI7/5Bmg3tqIGZgTkTpOFkbwgYYAMea2fPHB
hmOoUzushDLzooYDSd4PSVaYJTpnZs+W4tE1beyFbiCAWnNrKSE7+jPXeuR+
d6jemN4a55rjmAghOV76m2l9wqnFBd5HDcA7/vNs6tREr7TARlbAMyapwdww
i7MJSINxLaNlXojLhzbO0OkW/hcQf+ZWCnpWnMFFtsAMr6fTKYvR1LfgFktc
CttmGKcdzz72kvzL6c/7vJhMWejiTgFL6VoezKV1lwsBuBW+QwIohICCd39S
G/DUiUojdDNXDm6sTlxqaHi2jQQM5FGhhTyj41eIA0gactMNhyGBXBmcdrpb
vqFDJKgO94O2r7YkP5Ozvm+MO6xZTEnvckDPWbu8Hmt25qgl5RpjA+qsp1kf
BIgcaPRxvASewVVFEg8JmoYUX0XYkDCbTOxkLBGVf1xnkfR0VE9xaqCmIGN7
5OfLqtF7n+IoqELbyeNfDULEC3txK+i2bf0sVcK+Lxp7CKZcJ4eAlK8HzFuv
YQh9ca8JMlkoodPgDJVX9QYztgxx8TMkp5G1toRiZsWk0w+fOXJdHmB4b4IX
NFTXsG0PcFA4gkYpXRi+WyFtXd22+IoEZg0R8NP3w6snFAk/dri+i+3hgAqH
CyCydcdvDi3zx+yZGRoLRh2uDuPWv1B1lKDo5dVfOC8ktpJg129ZsT1xxEo/
/57Kbp4yWn1bG5ozISlwk+9WJnQkTCj7/DEZyaLEyYaHcHE52fwfaMgHljXM
l6yFHRgki+y4A90DE2G7lzNkhOcUHIIhyk44aVHHeBB3cNR9DzdfhtgLY7eE
n8fcZ70rjmi2L5YtEGWmHa4+6L8m8Rzao/LGBEFZlY9QN3+KCWLYblLQ3Lxr
Ky++igs7JErBFgsjNQJSjRoVe778vgOqJVq48uQivsU7K+YEiXdN3g4HjA0i
yDq13xPrbVjcPz/Avcg66+ojLVBCtfJAFNoUzTj53kzjpdVUfkZbigs1b+g1
kfIZu6XyJ/SAeNRFFBTKmCX9zpFUDJeTPklUzMmDxoWyQgXA8SMdB4xi3ech
qawIiCtaVwUFgKrUjqPQWmqpLzEC3Qne3yosNk5OaoEC3iKeB5xQDR/M8897
ytEGSSxvJVEt77ijA0bzvCOqj02cf0rY6h23vMuNujK0kNnPQy6p2+10sG5q
+nvCYJdTiWoLkWNwHHdzEAhKecIkEXXH1sssWo+tJGsJMaOWxlchV3+YOMMq
6JpFdFLmu/mnmjNEwkcAjcPGWeGZIl1srpo/5RZ43b1VpO7Fm+s34BloXtyK
EVgFXJanxnz9fLcuTRbqtBA5nlMxS43XK6GyGdVit64u/BGhVzqP7QT916e8
TVBURq1hdiaP434xk0+WZokcS++W2FMZsXw2tuieH60hAIIc2d6THQiRrgZN
rfK2Dv5IdNzeqtZIgZ2EjqvNJXaAkNfJaW4cDGOa6gouZdSyDZJ3e3Nj3Ac4
kCU+iFSO4pyNu77HPhw/FEnKt16j9RD0auLb4elNgeEL1BzmDvu+LUY9PsZL
674Q4/gagDvL5NVXRpeLYb8XvYv5VfI9J6WHd0w4Tb+eZ/y0UeayAnKGKH+j
cYEgGQaeeahmw88ciZc1O9OrHsVxnfYL16kAi9kc7a5rq7XYies1AydERtZ0
86q6FCNBJC6UV7CulK0R0ItxsbtxXJaHgjXrDF9Z51rnqTN76GVwUSayd7yh
YfxUO7dxMrSRVMjgfSIIvLsj99QXjg+AfnLEbYfB5Yq5TE5uFVQ9r3WGowAi
N8QNkTpFNeP9h3Qv+h+cqLSbuVkROJMQ0roqnj1KUa60uawxLDOieEj19UPd
97lXdJ2j1FBI8ynooH3/JYK64Un0o/mf8wgxCORhtddD/8JT+eSGeBq3u0N9
zxCIzKLWASaAINDj1wk6mhHj9NEhX9UdapqHbp9auQG3Iy9/BrPf91qfxDTT
aLd8lI/84oR4zHjniF+9RjkWoz5HuVLXVLVDCoxxoVqYxye+QVWrhkrJGGxX
PW+CfNJyJPZIgaiFRcxkJEMFZyZQ7bNEg8aR/uFXv1x6qOPQa770tcDbneAH
q4nyembeAXDZPFO3j7WrDbMNt4xaqTinws3ObDsQ9YI0L/gUEYD6PbGtlBdS
hKDtaGJLvvHEaDoZb2yi/i5vpPpEfiB6PD58Acd/QjlHWA4NiHFlTfdt3mWa
wOIa3ciyav7vzMfKqgczU5PSo7KXeIE5Q9BHCYA6UsJknfGS4vAb3apQss0M
u5OeQdYQxlaAbM9K2Ej2yn0pYR6q5M+3If5s7S0HxjJhkcyFM/WzqfaymIZj
g9J+4MZ/Ru3aVtW6zkLywiTdIgoV2ARq6E1I8mMNVJmIlLEIlnzGAIYFlvCH
Ifp2VwMxRVVv4Wk/3vD38l3Vp89IuBNYebl5vsv9vxQRjTn/o/OL/dN8v43p
S6NOz694ItYng4bYkLYXfrwwm+lviWaa3DouIQApwVCGMWnfA9jSm1TRRdWX
v+zUhEanal6Xb/tzx8Z1BRScRiaqBNtIsVMUgvPMsTklyKnnSZyixFi2O5ex
usYNHdIAXTXsW6T8RhBA9R7JpWV1FEuPSjGzzLHxM8KfIaNAlK8FnkWG4h8z
ezp0CHd7HqYarSw9tUP+aMccNag7ab08efDehzHy3TP+l3/qUjjROsHO4eij
YT+n1X0QXG83ZTvccF0PNkaokOIRRCnoPp8sxOPRb6z1OCAQrcRWHTjNahT6
NJlw2mgVQNmalAkH2G8YGGEufoldgqmgWQgJSMEQXFmCS58pka6TbFejqE64
pIbPsA129ipAi+w4TeMe5brVfkei+x4mrJtDp6RP6b/BVqdEZ6NCPwdR6Jxy
WaLi3Ksrnqh0+pvSUbg5M9cX5rCMCKik+aia/RsYa7i6N3YRvY9PogK4TasK
rwspE3hyD8jrN57h25VsDiPV176uav8qL6NA3FFcdrHuDhzNQ/FCLeTFMYxq
67SUFIvRK3UwILJYHehjf/RoX7ioqKsN3sem1hP4hVmzIhQk8I/9ln5J+gOT
mbSa1eOZUuVkAvZXa+sE/8CbaT9Nr/JfTn0HCD6lNBJkCyRDyR3CAYPN178F
BvVIAFoqeNURlarszlf4FqDz4uXlPm0ReVUcP8CDMdFJRxGHwxru+ilD6HaE
viIcVYpd9YQ42iVFFhBGznFzNB9VkAcYUz2gfgtAgcavlE2VINQQz6F495SW
QWKUE8DSoiSbdcjhA1fNe3ERaDZDsUkt5iMQYMqgDVsS2HUnEvdSj6yX0Ibs
pu4vcwi4EtJXHDdG/PRv6rxaDFeJxSQ4f4S5MoWOW+zwYIr2u8sPsNTWRp4y
yYKIqvJkDWgW6meEOwi4B3c26deMUrStwE/1k9X5mLGeMfWfTt4/19DW4/UF
lzyk/HNQoioBwPNyHDl9Gaewhu/kH1JbW9FzIE7Gq6Wb74p61+t70iueP4no
77/UvdbGWuYGbiH1JD89/r4POw3ddhSQHthwMvqkRE4eK+kVY4dKlWek16ve
cqMpH0DY9qKL+Ns2uKeVbiueXVbw9Qf2a9vnhhsMhUk+LMgxCVBVxLi2KI4+
QRneWw2ZHOjUYGLBKux7NS/pD7UjyUyVzROzuuipHyxv5Mam+vzOWn563B1Y
M6d+CH2WVNC36BlKw1EafuZjIrblEs4o6ncxyp/SK8Bbw6bVHBBN8/5qP/Up
9myEFwxOQuXYWVbWvp/mLhCmwETyO5h26kfxVWRl6fBCU+iGwMaU4xatedpq
3H6qB219ME2+kZKmXxXXwvxail07eOt97yIysjg1EoArm9V42f2gbF0k3Tf1
88L0+UIAApEElwrEOTYkUCXmccTiyjihH/PuNltSUud0aXBo7AOXEVCqSf5H
AgE3UdxXawSX91aKc56gIBrtIXrAMn4ag5PQyF1OS8F6sjSe4kab6AguBWOL
zsYg9jn77+e8BlQ9iz/STbjmrjt98kQJDBHrZCX3UGRKjeUEdQJxuvSC9cdv
M0il+TYjmQ4xR2rekpwobafK0YUCvDqsyTw1ipESYikDwrmww05UfISRyaSg
tbxm8WCtZsep9bZN7IEesGeCpQoiHUuCoPBROOO2j1T16jRmMNijnifXHRCE
3kAhfrHTrA7qD2kM6f9neTOaW6Qtjndugt8/Lj/zgDPxAINxH3mv2RaCh13g
U2r5+PAIKWiSoaETyfAYLEZAkY5/vlkzHwDKHvO8BqhSHssCBjpdqRJDInoD
2IOw/xmBOA3H/u0Jq2c7pbk5ZI5d0o4nuiE2oISf1mptlZ29EkbWDTFB+xye
7azkqLsfDElhK3AfN0ZeEQTVW+OY6LKfNOFP483eO/Mb8uqiYgdywN0dAouB
HhcFV7Ol7lXohZ7HfmtOAXsoMl5oc5+bobBQKGlpxUrbzwUexk3gThY2iWem
87cF4K4m5kjpKhm5TE41jWeT6RkRbQRETsr0aN2M+c7XM5eS7C+mRy0COBea
mzqypGTFIe/jEUZwJjYh2CbeDAXzVv8s0bx2a5PQYAHCs77iE1cLAKgtuYua
sp6DnwjIhim2bzgRlby93VeAks+7q/H7KZCygw8ih4B6UVzuz+QqRSkk8Hwb
CLxPRACR2k4526cVHcUrUCNGjTk7QXzjQRwd3KUAxjDQ7+2iThUcYiGLlnTd
EOa13qTPFUiUXgAQ64f8DQnQa8v8DVU/+4vJpYWZpfjorZzC2ZQ1VNazSPvZ
oOwl7WvnsnpI4xv+H/jJEyx8Mrq+cyN8wxOXuWVptzO45NL79cxwyUduv/d0
CFLjbOKIYS76re5fTiczCwcx38sl629Ej4EaNgW1U19EoMsPPHx5UkaC/9sK
KzsfaXiDhw0ai1z/CKSAiraVY6b0bWalfKDJvBNFx/PeBBQ3P4M/fXavLqrt
+8J4HjLECysjHWurH6J+zX8OkANqFB9/OoiTpcCgXJ4v24S6kLwQ+Chj1X6S
daY+LHm+jNexRZ4DbBKwi0cdADi3RAb0jPSrLLaZqC20C7nO7eliQuwW10Cx
lFDmKkNhTEsEyFgm841yAifBNCymDcxnSL9hP9yn3gCYq8qH8Hn0KeZolkEv
ys4esId1CemZ0wiJ4kZq0D3D19QQiexEm51WXWsumhzmt2Wetkrv365/DToo
o/bvM7TtIoMLL7cs2AV9GyYRESjruZ2WL35G4tfdrfR0pwgA8we1Jdgnt69v
7/YcqOw8jdHnzayr1rUI7ssHJbtJ6Rq7H0M7sZ4iU6nsd2hfnG1hKgCnIjgX
8X8OgK7IFC2Ns2q/gbXN0IWzsD1GraKQJB7n8lQcasUQGXOjHk7DcA7D2vKR
5jwtGPc82Q2e5fhwat6SvPGRF4snnMyb33rpw7WOiw3wfqj+aPWf/9BtSNsq
s+9sqytHR7AuNOrvXpVMNLPUyKoryanmW+FCFP/9lT2BhFWa+Jd1ivRYaRVA
ZLyBDbxB/1QbcAJAtPPmfYOOCXJZJ1Be0S5UyQ/PZh3+q+jqfZoGGOH32baB
+cg/jEHtjNAG2W+1G0z7llNdZ+UFcLOIDiXDpCvHG9WnB+cak5drvSGXoTXS
ZRiyJos19j344lCfy6/EDaOO/dtjMhueJNqZO7ym6W3tMNZ3WfFmHu2wIL44
goXxc+h2pCT2n4SZgxC7hPM9OcguxP1x3Gj2ve8mm6mX329EA/FFv5PxAO59
HIPjhScsf0b4ic/GXyYu7NhkMLBh4fdz00R9HGyla5av87RS+QXuzHfPhGFB
fJtXimaVKAwFoM32GaVtifDAuOqyNJBn9WPml17HCXSBdUMR1orU/HE4EMJt
ACOtA1dOI/HT5erL4/bz3gCcADl7l3smSKZSxeGxzg3+GgLszML/ShXQuFz+
pIvMDp/jPLWWm5mRr07K965AMy/xz7T+1b+Tc0yiQ13S9JK2THo+jGhZqk+h
nuLw7wsDe5u6xrwGGgTm3IrLzrkQM0t+99Ai6tFr3CJXcmoyOnTR8a9qRvno
fYIxwP0h/Si6AhXFIeRYKdHco+JZjObG3zqfukfmTjX3KWh7Zsyzyeag7+hh
A13EbrR12f1CeoomfnLzZ6U+DGS8/2VR/o5o+Ki6Ojlu8RVh/AL+jl6QW5D6
Ac09aFjRVG4C4XSqzpc4Br/WlhN2GGqQkbkMwPt92eFBuhTKB4jduoK4xafy
RkILknJjaUE8Njiw+8vdsomCwBYQRSSLd//yctLiWEVkiO5p3Q2R3XgS8jI7
YPJBBsFXMmMklX2a6D44O3QSl8qIPX5DHRGefViP/JW5Rz/Lc99ReX+v5cbd
HQlo+I1fj2gQap9/PEAZ2xJ2ArzMTwBooBAOh+zeu06ewyx+SQr0m1a6do/c
ZKB9njp3IrMs5w0l4/rJSPMI4dqMq/KxhrZk09kQU7/Wh1KtCL0JvRsBRrIl
/5s8k9X0EywtYiLVjT8Gd+69Dv3/JbsQcZYW7Os01SunT10Bp2G6QsaP+kVE
YzWngfgLS52stlPAeLMtZM6h7MjtoerMh+DZV0i2PZkkvW29GWio2chL3D0m
UnnsMLkcAEzfKgvulK6qIjWKEuuidMdhodiUsCJS29Fnd9YbPVFeEEKvyG/A
kXUfAiZCwScfU+F+aCkQX9iawVKCeD+JPriN+itkBa0goprNH7sMtLm8zuur
GlXD8UUPmNIwpi1cEIHqaIHhzPQEAP4VlZb842zuLgCX/0LIQEf0KOi4jSOG
twwzi3gGfshOol16VkIkhK5eixZWrF24oBsK+x+ab20YfzzWJ477P3LwYHi+
EkeXWjLhyNFU5uI7ryoRLWKbTntd5pw+rgLTWA7zVSd0NMfALHYFp1tEQs5S
qQcDgNuePUhVtlyOg7ElJVGiFpneTEgZXz9PMBkALApKDtFOg5D0+ar+mLG0
tUySZTo82Jt55bboKUPzeHEE4k4jAziFJDs3KOS+vfeCM46Ba69Ou/KS3YRV
MheOH4gzZbciI6JMZMFxPtzA+ijHXy9nvZK3R/49qjOW5uJArz0f/9ViJp/l
ycrM648UdwJPwRtFBJt+DENF9eq1Cx+MmJNlG3s6EiByx/Av340mwxlNvvpJ
cyXv5kmJCiMRMo49H7yIzC8qfnJSrc6khJrD0t5Vq9nu1ofS66TFjD9cSby3
tvRC9hU3LPM6YXGsAb3/D0XQ32TpTno8Og5xj2ERqyeTGYj8NAojY/jdtVjm
APVf0QBQhuSLIk+srZEshfq7Qni1SpWIBQ1H9DYwAck4F1jEtE23iKY3WXaT
3SIsyEZ/HdYNSl/uCPHLV2ucqpdiSgqiDterNJrFEi20GDYqDFdE4CE/OBiZ
hkUKWUjoj6BxkzjejrAk/8XeWzZ16Tk9ciS+PTLzdLL6FGLjo44y9adzAH1c
15T4NpOfaVNTcRoyppcgCFMRuBqkEgBdZ8dQfNi7y9B/slBXftnsuAXSqLSx
bDQk7OVmSCT78vRlJSyIFdcqOSBWrqUbDIsrYho+bih8A8vHuI0LjDvAAkEv
NRFyc4xOGwqWNu7XtF3aHMo8nBtaQgKFeYxgzWw6D56aitgdo0Pa+e2jRtNK
OBV9fxHZ+XQTRDq0r4txpDaCfgtWRN6ZHT4spGDmCVMph3EFC2NUkL6C1+HL
j+WnPyfEaf2/wESLIjBY+csoV5L6fsrHZQn1v4lv44YRfZ/APj44mr3o4yiI
IOmDXkxGxvpP6Tv2lJW05sAUQbHYq19KVivt+L6+30QJwUp082WFzyTd6wW1
qtHny/ZP+i0HCFhh4JuWmf8Vt8St5gtUfLdDt7ksF3moU5juq/YRRpFdj9VL
fjrkYIDBPgDrwvP9NfIfigbmkk6WsJpmk0tCPiHYwkfO8xOG1pfSD0QZLCMV
ZIU7rxVBBb1klUzzCewsnjwqKkLmw7jhTvvN/jYXib+ygNsSopsIZPAmW2SC
zBXwwTbCPva6fOYobcRFentmCC8CBoCROC2G37nSJRq1pEj+sm3U7tbwiqUM
HQxO+VWF5GJNf3hD831xLwQMC0ngytuRoGuGLFDeMHCksKsamYa9mP9GxCUd
QApIwPHBZG9tSwgPIkJkFftfIqk+Inr6RVnewluSBuOEsYUGMxLPGMzX3Mnf
BpS+FjxCseMvIINzAKfETdeiXhMkSLqvqZ/A7uUuTUS7OBmmfK61Y0HqzTO+
KoDNw6PBOAK6kNje7G+7PbT3S9Jkt7Jx8kc85mVk2xpLt6tLZ9fxrwE5CBFs
IwtbscEBgfqvAtkPuHsedhvXH1d/8hjujLw3t2lUGjAK+oqXe/iU5HB0KXqN
DzKcqSx+gb7S177i+hCnRJntwgihXvX2GIkRPA9LXAM4rnh/L28ds/OgvH9p
yFPYSpGoX8WRmlNGz6mdG8WNleoR/PisnclMflYYYak/YAAFwN/NTDZ69e7C
N6jfJGae8fje+ZSPNUf9fNWdyN89EZdWg052kd+ye9i/JlB4Yh8fs6eHtP5M
iipgBl0SvHCDalZk8mqegYSxl5wSSzZQsw8EcYe3x1vJ+W3oQnY+nMHMf8pa
YWw8wZ9t6TN+6MHRJBO+Dy+GQkMc8HQh37oEwdTxjGdpflomfjRITw3drePN
TpNYl8o4afMN0sgIMAB8Tye6VcxRUtLS4wZJcVW5We2oRb9XNj5oOg23uC+l
7akHzJyAYveA/f8OKtXWDrVZBfPL3dJa8WPJksJfopELImkiEwBjN92WWe77
v5KZSj5HPxahxMozsQYnl0A0Ku8jLce7+ZkcXL9lSu43LGnRFkHryjohiizY
4/9COJQSL/CiaeaIsvLP5JXGqO+xD/t7Xc1yem/6YD2LS9V3FImG0HRMqmlE
KBUFVaDGRJYStYWkFynySQ7Nf+2YWBOcw4ylf3CIae9xbq1R9BO39zC4jYKI
xSWR0f6KyafKypkM3qCcEbdC3Ai9nwXQNia/dWwEBsx1y+2YwcDFitpCddS7
KsLQFwqo0YCDQ7gPBd3rvCOqbdfajnJ3r8GX7UjQZikiXSRi4Wdyfctf3y7q
SlP0hWlB6JchpJz6wjJhkeO+zwvxorTK25cNPubQgQYTx2aVzsN8WT8mF/a2
Y0o1zIcP/ClA+/6hCP47Ypg8vpjs4AXsJWwiuF41skthY2/jgOSdTOfRlBzV
NTPYqEpxfL15YeZqxGcsRbmlrLhN6Q/Y38ZjDFTMTR8F6zWh1p3TFsdGMMwF
RoaI53MtkQ9H4MLQMdH0WpQshue9Qi7nk0oDsDSge4mUTBvY1gdHbNdNg0Zc
zHi9X0J/diSoFtN0hfRHAUpoDTBjg6NXWEI3mRG/HqyNBljM5LJ8jnAQYSNB
JyGoP0GJJVRFWZcDmTUhfag3uS/gAHJr6loBdxqmXwIRFhXQdhslkURoUIvv
SOkjSBKPAHNq3CvQzqCCXxAi1TUAsXDX2Hxgc7kGPzDu5aQa88/BZYy5eS6a
wJ+eBXTNwafbawZETfACPdFFbOR9jxyJ6BtCxLMQQMH0lAyh/iznRFAZjJ76
XdjkpNLcaVxIZliiSh9aHZMM+OQvlmBdCEnMh33RFQOn5WnB2/uvwqZFO62u
2SPuIwqSFRA96DDMYxG8pk+a2nub8VyOyCCKp+X2l5pwY+iUJqC/+Es2PEOw
tRJoR5SEMVznt8NowtCZsqFFUWQzEKDtHDN/C5C7Krj7j3QqxMEfZqEc5jPk
D6+H9D0PQfJIRKCfreVffFyh7SRNzbrpssBg8WSn0/y5JcV5EyGVZGwburLa
ZJp3ULC2WEepZVOhqdinSzy1flSA2g9LrG/lCXbpeFAphiAt4PCzPDbe85jN
F3mC9aNbuvMgKIByCajFLl9E1iy0DV4vPrV0L5KWMzQmIJ1C2GB7gV0PITxm
IX7ojvSIpU8UJaaDddnEruM4flaAlgf+ErhXEKD/gt4sJdK3Wv3CkPQFFp+j
V62DiHgDurvT4g7fNJoiJaEwbB+ACI4TIBincHEGL6hHYVXvlbdP3/FZF4la
LCnD/my7Ve1gKhjDSlbN/87Ut4CTok0O4X9cztcYeRM3E10rFHDOZ7VFJ5h5
owbxFRy4YkLJYDGWxbqqfmaWhFhtjzew5RyTk/WeXks4wWnVtJyLiUdqgh1Y
fHcgESZgOV72mUpSsIn0EQtDENRDxurOKKrx+2vcJL34CXecXhXkqZzSdjb5
ypSNnGfUO4PKoks9qhsdntu4YQmI4bBFzSwQDP2+vO6G0NNmeG5vu0qaITSA
XOGxwb4aXSutIg+yafEYqU50fO2kbQWyxxtrs/ohi2TM8nsItJs515rugHx0
jrGkc0HtO1L1D9+sQYQqFWTmqwEW1v3XnDCq5GWwCh4Vy+nHwjAbz/bA/sxf
HTk1WRmAuM4D1U7uCRrfEJK4npgtey1xVmzKq3TcngwbLgSBiDN4djQmJJsH
FKKd7n2+cbKitP92RQ6qxZld/R2xnrJbQg17SDssT60VHgfZ+laJqFfOQ0eV
1Rna/E2EUOGMapwpUDom88N3AMtbPN/3Rgy3nQXPnt17hQeB6uAGrmQOASji
mUWLOeOGdfkGLuLcvOoDS4hG6cwrUCIIMyhdfmW661NLis8mTjGOC0YLTXLX
D5hmitVPRDt8bEmJfcEo8V3BZypwg0ec8SWnFRH6oRZl6/UWzYW6ZWTftJuc
99Dx8qWi5apw67ks7hgRclpvh+n5BY3PEHq+oekUciK/H+KRyo36PYHc59Fx
imNBR8UHNimNi/Za+7FZM90IF2ieEWzwN7UozCB0nyAk8nDHlp1pNh7OwCUl
lIYjgqIV7Tu2EgXE0F3K4FOrGEO9zPuLVUR7GIQTgPYRCqjuPY93LihuGkUG
GNeGIpoYnNIVIYG8avedSDgxiGlSp2sxwmsMHhP4ROsVGg+w2UMCUtpjPNZw
56awzd5vsUImmCqVgI/K/bQhCiVp6tqmeCs4Q43Ej2yRwNL3dtBcViD2phOj
4tvGL4l+hqjg/0AIVjReV6tolV19yY/q99LFG4BKyZa9XdFYg2+/1dYD60zt
MejwAJZrN4Ep0PM4UoMIswPhECeX/TaDEqiapCGmNvNi7n2C+Cx+WoObKoNH
JKZ/e6tq4DOaaG7QdNFxojYd5qzHnxVLkngWtYHSUwrKMbhPQCvqaITsRSBn
oICxrQm39bjKOhWfhQze7EY+wUyNUs/m/2PQYLv5uK82/qoytd59giHXJ1SF
VX9VbCFcrbbMTUiRCW3MrttpQlRMSlToVxdEd5XxHmN7oS7ZgHmv7ZOJ/dQ3
uzBVwd1GF4oDvjmHWdGL8r/bvrCNKzz7MIKIxOYman0Btly7lcLklvdj8HCQ
YtoIeElcvhNFEX9HsgiC6Crxwm6G5vqxMVc56G7KlR6+cjhyxipQ9gTpz0Ob
GezHnHZqq1hWZkbjVRlLD1Bja17w0DNU/jmEE4Wj3RV45gkQD2Rav0dseBGa
XvbUwxk7YSZyMsrs/mttIPwGmjt9Xe6gsXnO7Qs5Ih4QqH5h6CGmQMgvUX52
Sy5lJm7pFaPVjBLtbQhMtX+091AH2lERgEgF0soBlo4m8cLT3mDqUwULhSNe
Qektk2H9z2j37+0K8RaSocmGYuGLYImcSjbCx5nEsPqbRakNqCdqMCXmJFTm
gzqwOJVlfxM7layFqciJAbWZVfH3XM4JmBQZwcBhnVSAtS/rPUafs3LDF1/8
7ra9fZADIXOYgX0PbpomSP7vVc0gBrNK1yclqXjpDVTr5gmCfHITEeDa+ic2
IX3+eHAgvjcVOiUQlDMd484HO0WcrhbDXIcawVporhgdGtIiRhAkd20vWTMV
0mcwPZGmV4ftggvN7B5Dm4pPFxt7fxjxJURqMv/rPkM8xqzEwlnSLnWoXRZs
Kuk5SoHmyooDb8XjNoreTgU1Yz2F0CpJTUkQVqmRo6BuKls7s+jcbE15u36T
CSZ67MXdBj0f5QOEcYs6goYTGc7kxqAzvBZo5sNRvClDBVQgC1gQ4ySik0mB
uACVyrn1BaVL6J4pR/uM5GlFAwfZcAANWx0v5fl+b3kIYpwLCzQqri1sbuRO
va+5GaaBQ3+p8FnWqvRAF+y9qWCG9qwGPWqjnrWBLGM/5b10F3bCcNPbW1at
lfaFaHUoFPTr4QecV8iDplBQoOqBbEsOkCDI8Lx3rPmUKAZKFZjIdJnt6Jgk
cz7LWtfShYkHIx8uXv61ubo/FZlLkMNi3SxSB+LdzaMEROmjkHjGCCs1frjB
IsdxefcsBGgjUXlbJFwtSVcSTERxZelzJw4HLzx0QWxET+6ZE1leVE31xIjA
wS/Tj3bh1S3Er0Ybw63x8V4RiHAkn1MIC800RtSAQErW0E58Rl2r4hSSkqh/
O4e2KJvVZLnjKgTICfh/mhYdEev9kUkcGMeh3azf8o62Pdi3kGRArJGzve/b
SwM/Mfi9ExfBMBneWRdrjleQ2g/ZbWOcrFttdTDs7xQopQWcuXUpg9nEyaUm
JvzopEqkqTu4T6t6hjUV9uROlm5pY/7GQWnnauQVe5Mf5WlLFlKaAW6/5d+N
IR31mUpyUUK8KJPgZN3xZAnotJ5FNTKJgpGxkdllOohiS+YKRcqUTbehPPw/
MYGURHVZIq0bLo7TY0CYGo2OwAWyzssCJcdqxKizjHajzLIpBTfm713ZoDOp
12bu5kjIWFFoWryeAwfpYRPWurM9Ge8i/GiE9gPrnvLdO4v+ML9+PJW2L9Km
HL7zTzSDfkk5loz1FLNTVlvoRf56U8DcESmFcVvntlct3kqYfGAJg6bKntHh
jSBmt6xp7E0SCbjBMoUlDaIGhVPEaioLzq2LevkhxYeP1DBv0HYF2QCXmVcm
xJFCCTSdvX8J48c4HzM9HZNfCuh3JFB0aVi6Q2DNpZMAA8cpzNOvhiDGWyTu
mRRU7vlx8XU3Etc6bfMbhGtFDyPta+XtYt33+RKcAsEn2aWT3oUHU0JLiIbj
lJ45jntXXmIlKt1smhsCD2edqF+cx+Cv2+3xhn2RH65Ko90BlPdiPY6lr1KY
oo9QtT7C6izPDjnmvx29fCcq+kWJOWmoeMR9R4N/jNNYnEGNIOAXyUBivKEw
bho+BB4k+1PDZQJJz2CoO7krAlstA1GccXnFhUa9SRq8uA4h5MOWOD/dwkv+
S2fGM4SXhAj9C2Q//BZNEWIgQMp12tHzsEavrgUDja+v8+xwQE0M74v3ImYd
j8qG+bFH7LsLQmqG0/0QA1TAhwMfIXHWAEdlupoSPtnuN2+JncWGu2Vin8Pr
ta6KpMiO1GNnC6L7EGG60UnrghHaVbpXcpOehld//w4J3ArUlDTz1uoxImYI
mP9ZtfFc0RyVKdIph0jdUFuWHaV2Ha3Z0Xp2Mkf0Z98w90PZrGMw+NtcgpyH
UZaaxXv5ERIaNWNX+xWG8x1HfHo8Gt2agE9Av7dkCLDvDAYRSwXNabAyAnfF
OqvJ1z/xM9mG0/Y+ziPy8WpHZxxlOqAHhltKzHoXMet2bJP0kleL8Xa7YARl
o0mYEtR5GZQyqjpU6XOILE4LHS6YVMdbBFpXUakT0BDsDAp/sVd/YNKW5wEs
xg4Bl9O9pw1gUpkS2Y9Y0Ob+OTogoGZdurZbaWsZCwOOpGE1A0t6ZE0kTeUA
t1llw1EYMEaBW8izptcTDmYM2RMo7lsZNW+7Y+Tl+MyQUv2UL+eTIKoNyHZ9
xUBgIQkLNmx0avFOCS9DoFezFyvNC70RGw8LFMXrSkXAOpp5tIkyRGY7r4cG
IcuM2n1f6ws0U+EQTkEJUGf09qnVdkhF5E79L0DLgy/FVh5pPgC6/JNJG4iw
NBje6EouRenXE4fqhKEIVgy0Ar31dzMN4t0pA1kSg6tsbXSI1+NH1FMLla/u
1tGGvw/paIwOXKUxFw8Lv0n2EclKT61wz3ImLYfIA6zp1nvKR8u9yPqUtHja
Wqhm2VV+bAhK4JSidmJKpQ0pHuQi2OiBqE0dEp8utKnSUkiqpEsu3id4AvqM
nrQHR8IcTKcAV6SfL22YkZmTTiYQfy9vI8SHZSh6DacjcU2DVUBPX+1hDt7r
9FR4U2rVLyc/LPZQUCNovCn84oySLqfFbAWr6kO6CZP8aLhgx9JKNlHCI2y3
jEPU24kQSVDolwMHfZhXOAnZB2GQDvxY07/n4+8dG0P2BbJ0gcBiNBi/R9ke
r8H+eV5u9MNbOjnP57dVRV/9FbxKvnRfKsYpdXcCLv7HXMK/OOloOQ+Zu52i
0gZ0wSo/SXRJ/T9czF23vRRVdsWH5VjOiX+3Tzh0g/ti+rgh45eWLggCL7nC
d142UI9s9iwAv++cP7k6O3r1nqc6kJnCLWs8O3nBruKd9ng3M+BYMmFNl7NN
pWJw/qlausUf5GII6AaK3wB8OkMoYmpSos0qzUmZ4lvfjxtmBLq/jVMPZ46Y
Y1l/ZlwF5OHU8byo1PAQIHU4l7PYBtU2V9+CGFNVKl3gQl1Ju1ITuEKHZqIy
aK/2oi60CPVLsk65nuroeDIwyXoSAs0GQtLFeGWQ7p0Ew2NryW+30GuhU5+n
UJiML48SSXo17/dtcs6SCrt1ZO8+XTOnbObOlpAw3GYlJlAnAInrJvtBMLxE
tSE8URPjUELfqrhkRIi2g6ju0k+xXA+o4oZVV8h6qMVPbrKUgznBkKtYjAwP
tuyNW2zbF4JvKe95Nu6g8WU1Lg8kU3Kxd3mmhGdKQ1KyQ2n25XfLLo2d3zui
JxN9jr+/Tj/SZFSBt0qPsxFNQSxP1caKW/QICoRIiXXH7Pd9UIa9UmRO+aim
ZEzSMeLlhZDlPPui2+Y5FOvJZ/gvd1piAIxcBNx6KPku9rO9td31HNkJGMvH
cuRF3CBtoyipLVl1sJYx6fqkz6HdjyPZ0JmnvB0XBJXEB9ZbBQSKqZcIk1Sv
JUiIEUweNOLmiKy0VsMQ3OpY8P7Q9I3jLLHddZFUXhM4Of6DBDOKrbFKl+Dg
RP6DoQlohZFBOwKXjNVudeKSc1u7xaH/lN2QlysBk3XzlI8hh7DZ5MWTGQcX
udjvWBqcbiEMrVvdduQV5xzOlQSL+uDber2/+oOfIOUCBrW1AlWo6e4XZpGU
AQ/pOaGBPUPhQZ4MB+0GtuUhD5oVL8Fkq+4P5q+Y1QMANUPFSVSK0G+Dwqw2
E22ZNTopjO0qgsfjPya5Wz131PNRmrHR34+ZFeRntc1vbtJSh0DVWmLS1DqT
GRF4fOJtTsXN3eYtdwgBaJyuROwzYN/ZwWcD+dJ94OztMCxG+izpBNHIHgUf
qw8YCp/ZJUUqgZzfU5gYa9ppdfR7+McQiEdZbOATP7CslQ6KWh48w162FZBK
+2ST87G7xTBO8VB4jqw7YVqrI8rUIzsHdLHIeYwTsL1tKmSjQizJcYAoL6aO
UwO6Qv9f39IV+EfX6NG8EyBsC9qC5WzZy+/XtnLFahTRtswcCYvNSln3sjQv
Eb++lMd6tqAsgrb33IMP2nz0H45bw1/mdRo2/7ohljxBKjKMhg9Y3i3gTjZ9
Vt+iHMV/1ksTfj6I/IBcnbV0xuyOUwSGOu5mJyHkjRyMN/s0q/LtHaKsiLRo
Ju38KGcgSqmh20xgNJ84riwo/FgkN8a/2zEOuhaeacV+zM1zGPlR6q1xaGbP
NErfvitzej4LuWIqSmrmbQmQlxfEuCRhqrADHZVhb4Zdlyw895XPrYbcJrvp
Hfq6mshXuvgDMDIpBrlpR7Ljeg9/ZFO+g3WsgtoJFESvoGv4sMYkpFj4IWQq
FUU4WCXRPQUKscPs+9Mz2Sjse+h+zyWjTbag8czO9iGQpBvsm5gLyPZUvBDR
GGw1Oj7lbamCYTH6U2ZDJXFLJkr8eV6eh3XDU3TnvIq41e37wVmUbWr+AeBT
T61eBLRaHVWGcBktAvYbSTSGtvBa+ZIPYF1D7IGLWaUf516vFKMUESmJVYBw
aX0CgozlpHcDUTJ+BPhFDQZnPtEL7GUWFOGfwqBJ20P4+Qk5yj2FogaE+Puz
h62WxufYboSlz6lkV30Gx3PhpIZdN4rVRwyZUeq7wLr6gEWoZ/MCXphAzEdJ
NjDc2LIcJcLEypZPbFpvCbBCf56NXXfbl23/B5Itp89uJf7oYZF2OKGEckOW
jcmKMcqv8TSIeFtCOU5IJV3+TN4PEaR7bzv9G5Vb0FYUhyqOzO62Oaoqp/OM
2hF0FlxUeQM2euSFpfbdMJCmF5V/ZQfMnMCviV3O+HJUCVvoGUc2EJgfDSAo
mmK1inmbjYzLsmL59/5NOQT483OibVxHhPOf1HygfAcJvI0gweRhtf7DxevG
nq+eG8Gj1ngGC4p7ewFyEAQYdT7lKzn7jMeolVv4TELZIcrXLMxWEoOt2FHs
Z3rGajjEDUcuYdx8x98xI1nFu2ReN+91Ftub2tYSAPhcwFKDbOWX24jcilCQ
yxi81tm7OG4ukKlxRlyX8EsrrxXkmaK+SfqoqtgEvAxXWttATpqUd9sIHQp3
klVFFCt/w+Fh9py0qqkoh6bZMPXP72TPDgpSrxFraP2mUuAhiQUbcmeMqi37
fGZkfvVCjcFhpyATBKdMStBEBXjeMjtqV7OxNQ/6xpqzw1HW0kkYpr2cjLOy
EOhuCMuV2MMZETXFdj4say0pCgnLrqYJfiSRzxQFYTe3jMlTtw7RyTMrx3Dl
N2wZojd7ohTqJK3mciOioxXpfKJaqiJawv8ATiMNKe4sGIpu7vqN5bVWOEPF
63plhGmZPtNg5VB/MEY+uz1K/T+oo2vv1ViIh/lt2zz6rXCAK/ctfPQbBkwL
CJyF9ZpHhBOQN79Q/4fxQQuiKI8NCFIEikCZPjssj8OE+L7mwb1q5VExW65K
Luq/W55SfydGeh6OO5kk2No3GPIfSPxGUsqWC8sSwBZU5tmhO5LJt1yWJyqO
ky4DzGplSVzyhOXi56jHkLoVUkJt/kumnoHd7AzqEZ2WTMA4E5jpZYkvKeIf
j4e0zkmjddYujjvQ8hAUGFb51uO5aKQTsJ7sCwqV/IgZBuQ1s0xWzU/0Oo6W
CUgPEiHWiHdfWMImpB2KMCP57ocdc2YdagAff1Ndy1ZaYdnnXCtTQ7u3eG0Y
vRmtf3JmNNmAOVt6pBS9Tbb4Lu+T3odlQb+D3SZp54myqo+bqJbLZBv+N41P
aqQml3WRqSpMOL9F5UdyoUkVs9BEbNnte5ZUFv/Zr0lHhRZz1w7uOCQGey5W
GiXBVZ3OCuEv77cFpqIPrJR47ZjdUPm8S07cQvt7qIpXMWIdorOtDq1h2s5A
zLz4Da9WpFGhOya+RaCirX+ekiFfG5LiTYUvj7g/gWsOIAqZxvZcRwh7irCY
bKRxwoDENjopzSBSWDk678x3ffFz9/F7fNW3YMH21zQBbDXfE7oua5ZBbV9h
JCz4MR3Ee+2qSjlSdRUa8ZFTHiwX+IUcNSSxsS5Sc4Ff6mq+lSsZUJ6p2P0k
6zqkgcUkF4z/bmG8Slj2zoKHop3hYPZzpawYgrb6/3BBQnFJipy8GMVS7e4g
YpLXneGDGP0MRsavtlfMJNkDkYuWJid/n6ukXHLDAkWdud19ewa/ql4eq5i1
TKcKTqXLCqqgGU1UgcLKksg2K7ouUnmUH5nhr9YwMwjoHwhEQFGZY/0NUHCv
o3k5j9fRZ5XiDvo+25niCcMu0wkteMLIljUIQ/HDWAr/QH/HUoDfNh+p5tF6
uO1A5knxjz8l4tN4DrN+hzVLTrNYX9HQYjvgpI+bW13Olp7ko6KDwXuOAFSx
eA+PVSyOK70FkxTH6bmFCY7nAKZyQdQMKXm4tV5XtoD2qbIWTQgPGMQ51xU3
8WhbTcrOFlF8DkVsUGNuxjzVi9NqXmVfjFXJ4ltyXgBpqzNxdvyrXagASeId
g7OFqz09jFW2/XEjnfU2zvIc5BBDqJ/LuaVgu7xKVcRAHI76Xd/OPU7maouJ
VGeoZOIvjJ3EIj35OXZ3uCzx0rwz3blqp9Ivv4JYkEIZtGoxJqg40NAvP5aE
4JxPeHA4u/ZYvwOxFDv14JwbsTnzgy8uhOQozQyrplhvTlru5ymQ+z0EZBIQ
GJWreTQ4lZNHjFooV0ukpa0T1UNjjk+mnzKQuggqpuikWmHSCoUIfktahcUJ
nedzhZI/miZmFGQFW4GRcrOmAOLNippnFt24HZE9A+S1iKj7dBhYGzcD7Yzr
17Fcmc+cBxZCHADjBNWXq6vKcete5D97L27aCUxpEeMmJ/rPzWEBEEEJKw3k
wuHLqoCyGUPHrgWrnOGOdmqvfR4cfAA53VTOQ6NiWBfopFywQcjRno71tBHL
TDDZaksqD3tib2CgYX4c3evjK71HvDWYWBW66KUFmDWthJLctjJpZ7n0LyKu
ObxkD9MZ1uDhPmyVe+mUqjHbjwoNQqwuOdGnG0v768t/fMIfEL2J1kIqhB81
vnMC3eqxTLRCFZ2O/qbatlZLTHi9CuUbMbDaah5N8GbEdOSvkNnxQryMWW/C
eHYq3L1a23YzidGwU/9+bz/AMxl+jK9LucSQvLfTmotdk6y4VIBSkAew3/yE
1ykWY0AYYmGFI48l9aDRz+okjjtNdNH2rxme1o19yAsnhB37Ao26NTyW5ZQ3
HI6YmadRSol1Dwbdd0LhDt9u59UN3qfwQrA1NGcFPZjQwZwYDoLju597ofey
WfQEnVhROPa0gkeH3IvoEjVeasYOzmVvL6LfhiDDosCe4em4qLTRB3lZSxlo
hRuaaJfDpf9ZSzLJmzAR9GmEAD7ClwW1Mjf8wKKuZvycitebcyZp7ncTRBof
/QWq2c9pPQ3lonAIbnHU1CyZ0L3l0xAtzCOg+u/35j2bTS278pMpLqeIkrWM
hM0R8REu4LGQdx9ScGLVZ1s0QdRGCwZc40wmH5S28iqhCh427jV0fUi1glis
RE5U3T3B+bGsGEPh8Dm51rn8a7ga5arFNQHLi0ZoZd1JV/h2DqsROXaZdzML
sV1scKaeLsNMTiu+POCsVyqkfuFkOW1wiGdd8JRiM53Z2OvxkS4eyn16wZYe
KZ/xm9psdv0Ft0LnpLkcZB2F+AQYcx43DT3pbWQ0/81Qe6BHEh62iLsv0LKn
pz07188WodyXfXSdUWYu2o2TVReOlSEMmtuGnEbfjTGbpJcjcJr/P80o0zHi
0/UrFFdWMYir5EBdIkSJ6RS9YIe8wMQ3/K36rivsb/H8xDdhgQanVq+DWnNm
+IotDKYI6pwya32xYbVEuqa6T8WUuh3qOUoKV9hH92d0lH7BUAlORFq5aiT8
+wQNQ/jeivt9+PWZW4wYyQSNb1DvrvrM2VmJR83YXhbxZH0tDFqE6kzA4iLy
wVK83w0MQLJL5wgI0Xf6u4Uyous0wHufL1GHw8/pB8AX4wVM7fnfbKOS1Gy8
OgkNLKYXJXhe4xkGCrSH4WbZLqe2XEdFGXGElp9IcV0Ro/+vaXzEyF80JW6H
gxSveDL0liqdUsJTBGeGXnqUolXDiUvG7Hd2cEaWDI4cGd32nxoe4D11jTjr
SCaKeSxEAx4o4554/Twr1roqo2ExGAU2ntuUKOs2DOdtNPXW3F/nukaSvezA
iLfUboF7p5FaDqLqORt81E6OPeCNko7jriu4RkgO47a2kTs9+0e9HJNFVFDS
kNa+xWT7fdtv57rlUa8FTU9+sIbWT2/nV3bp8Jd8B+TwHO2Ac2hE49cEHoIU
le7hy50KPKhkE2t2Ku/QfrCtzSrDOqcGV4A02nUDJJp0fDFMZwxMnLyDipp6
9ITb04gb7oU8u5N6mamozwVT/FuUD98SwO9oQgR2GFb2N8OgCNfZyGJhXhFR
wcMsjzIYvZU8EiB0S+v8NLKNnKmmT9CCDlJkJFZLyaRWR4R1SpmQfuPtqp9T
iUUNxg2INNRfGXvpR/jD77QmADRILZyUIG9QwHXEdoCWEhq/UokP9+AgM0sZ
AJWkUqwemYCtkfU4xD3mN1Ux7TzM58tK9JZ690CS3yenEY7LutcIbatHnOj4
4iivrKWjGzXeImsiUnMZYs6jK3kRtsyPL6XnRrzUXAky+oUeNRKNKOP0bgUR
/2J40EX9WAl/fY0CC23tEXVkkuZrk7iayoyADnTrIjV8oLQxGDnhIKmU5IQq
n9DOEeyoB/8wf3Lc1hIpQr4Ul9RMyJz/R9rnysdm3Ahq3FvyAIqAgZQkBJrd
HG/1N99ffgyRu3R575/ZkiKQ3caH/35i45yqEI6ELjdJ8zKb/LitOefKzIRH
dAbN9iG7W3m1xiU04nGQgZ/8tSrwmwS62JAryn1dezNla1jXfoBmlUdtAKP7
bFIqzgRqBDrY2E6tfEaF3Dw58ELOhFTmsBKJQg/g8snB/ZXhYIuS47VQCXzM
nQ70eYEmD7JZAh4EltDJFxGngdVm7wMqX7UtmWRw85gFwayqXPYc4i519GGJ
E6GOqnMOQZLl9rXuA7vwk9hOSJV0QxDJ2qS3wPGJRt2J+QrveC+TYT55/qXF
szek9Lca6kka67IGsYcFNt18gA3TkyceyicvzwYx4sKEe0JYy0EJBkR2TH7/
KpMAX5tFe0XSb3kuiCqF383d+8GmeKvdqboF0oPcPKhTntpR4BDw453DXSHQ
YbIgEybxug26FlbXJ6ifx9SPLFDLncYJrxrsvNvrYsRe18haAgGCG3gstnln
cVI2BGQuEY/JNLIxHiD325Hem8w+rjPdxHh+mu8HQhhxV8e5K1eUjXk8cCaM
vIfwyib+9Y9HTzEBt1qFy22eflNp3dJ8cFG8XQXI4E488tHrwk5XpkkzgbeC
mYcZr/VsYJEAw5LzdmFpcYtP/60hbYhhvyYWfjo8Dn/FMiGDdweTojgczhRr
x4xWnKKPJajdPsVOyenQDn3SXAaD3iEkAYir37DRqJSJKNkaQw3OI0cc4bsH
3+zEy0kf58Zf790RA4UIk3yYCcaBDGcQp0FQQoIUxN+CdMW2SbkOPFOPRk/4
kTrMW8IpNawuoZLE88qD9GmG3n6Il4Dr5OdLj9xUNvc/EegK0XYSwQZx3IBO
F/xB5POEA64BoiqIPQYonft3iEZORrO8ngcJm/L/FXM9cO2dzfy/epz9w1QV
KectMtRSoIbB8ag1iMBzlxKWId1YxL6YYasHsCAjunsw3iktPywyxJqiJe9W
ZKeetO8bM94fWYr+g8xORtIXEnNPA7FB/LHnJqHXFqqUGzgoyiZ4QcGU5BKl
ad3t6nRhb/jJ6vrzKC4wWoEy8B/tD85tfJstZA5bST+1C9t9HktiU3+p1jdo
0+wFYMEUVHr9wSduDMP++EJClLjOEgwDq/tDYNvqZz9YBslqjoFPEbebW+lJ
cQDvfBRT+TaC1wjrY1UzTVCCx6iluzsjPQL3aOConPqSRlXEfxlgyKXIkAs3
9hUY+/DKLqFsSoJkXHezA39xQ96TddqH6sfsPnG7chi00Gy8/MOwN1uPptN/
oPBfb9CEaEFOH+MPWSjiVxgx2P1HVrl4MfZlbbeAe1FWBFGFSVSa05ZaYOQv
16v2IQpxKlnWVpiO0oqs4yAWleosnfTcMm8AdCNpUiLYePz2/G0M/EjvK/9T
qs/FuU/eeJz6yvwPl/UJrGuohQfZtug3OL0HIpK6h7PJmzuzLv0prE0DOg6j
uU2GIiKHuDs0mgyAo8zB4+37wGqq5lb1gx3qjlAacJc9k5F34m0OQB3KDJzd
CjUmsGXneqnYEowOawhVYiPQcCiofg8zySRnnQuzPQgJrnj+HynycNfNZN61
+k337y9ecbDtITE1NwWeUcRL9alle6v0G8SoGPV0I7dPFRuV2Kx0uPFGnV5p
Tj3bCJkQVrlPasrjOKl+L3JoA5LTolY9szD0iZmcNLnZ5hzINJoFPx/YIQ4L
6RongmB5fVbryWI5D+IOdF2XLBhdqAjnH/GDeb/5wYVxRw+cmkK5j7cTWeAi
N1pnWMt+/dUiUz4LrNumKO1qs+YYYk/gvPhONGzkTLzNa2K+ZNVAZxquluTt
sxCE2jv8FcaVd/JDnV50oVWwtdPP/QGOQDo2tRia5HrXDaMyvwfmjr85HdDt
IKxP/lAw4pjXroddcHEP8h8WnIlFD4OZ9TZmOJoDFbUdZGFDSGO7T3rkOKhT
M6Wbqt3C8U2UhW7vvx3Kb4NAyZOXUFCRV4lVHbNB4TX1laLKYBsLXrSl7Rto
4I60MSwQdAemBePGqdbz25UDxwm6zOk/cqlVYIxtrmU6l13IQOyUNDiRXstj
aj83VcejLcJcrvqIqh5eF9hlTIhsqx9qb40BhPRqlV4ipMQmFt0HHo3+nkOE
mMp65dg1yq30ynCVrxi2/32ruiz4JGkuoHyQqr9XLXDtp936ArNZ32nHz47J
uGoKItrqCpFK5mKRN8z4IqqWDuNJVsTsyZaIjcXk2cxVo3reC8vi+iSN+ZDA
6brrn/vVajYZLEdSlHU0q3fivp+rLxTPZS8TZyo3KfGfPErF0dUqaO4Fq9YF
0KQY63wlTL5pBmWi1izpJOamNFmqe0SkZl2K5zMyGQl4/YNln+WEtIb5I+/7
nfeWbp0V1qXDF0pjwwNRLyh04z1T8e3geaHuF+Z/6bJBuuARgk47P7MAUA/x
KiuBYYde10ihoSg1OSkC2FopmiA/sJCWLpI/rFj7m5DAj7PYsYpPhT5VwNO9
hcbKcIqq0Fcug20tEVrioI4paBczWO43VPBJVZ64fuvmqQ18XkS37pS5yL5g
BGWJklJs+H1IjBqKrn/l2ORYMhpancq7RrvcMB6hRdO9HRXZmGBO2Ma0d57R
xNswIoRyLgitFzrOv83JB2+FHFvyMw2Q3D2iFC9rjFzpyZEFZjOy4xV9wNGm
VYsc0NxDsq+JsgcQVA4BGThzrJCCwLjrV4sDOhj2WE9qpHMnvaarUyR9V37z
HXzTQyAWD6U8Ik+YAvCAVbLLVH1hI0tVRUizILm/7M88JDUd5/oTXkHS1K5H
42juLzdSJJ3vaI93LXWSgfwaMP/GJB8WR8GMTi5K/R441yiUtadz45tGG+kz
7d4QlRFc3zdl8Sc8Ftj7hlxyoAkpLXM1K+BgXR9bpPN8xa4pWHz0Y3wOkLgB
pS/by8PJjhTutms5H6JD5Tg3NonbmpBQgDK4CTzTnqEePTA/oiJ7Hk0CLkx2
XzLLtjQqAnHYWwfWRE2+4soFT6bqmmOebqdWHg9it9Tk466sczoXVN5PC9wH
ONcODBp+9qJ54Cvz8eTyAkK2A9s72ACI5eWxp9hQR1jBcOmlSpTSnMzpodhq
N31t/EuYBW5mxfI6X4jrXiPmfXsmD/S/IIY1kUy4osEcZdr+R58jWBzqlYuD
QrYx1KR6DuVm+WdOyAcTeSMIl3U3QUDp7Rky448FwWm2sLBG6ZYSHnQwoYo/
6frVi5Dk+vOBk7N2QMvhwS/stP4ws95mycl7U9Vef32/gTysiciCRzuQzl7g
WTtwOByI02k16BfgH5eqxqRLGyR2Kk2/lT6AaJsMCtLu2Aov+Iq/XKOPH0tg
SchBoyzHnCU1EojqqASOFxSBA9p5Zt1WejWvIrQdc8Q5I3KwnAdgY+XTr6uB
7+IC6iD49JXurE/RO15fkhoGcP8ugfUHH61qmmv41rV88sGfXnRlzTobH9Av
BKCscmrgk+J1N8U6iMfEdhA2z1o04VFQTMH6+68cd/swkBlpxuGyNlqP/rhn
XKrSzBJEk4c8XhyGHskZuQK6w8HwujyOwaUDT12v4DHz2iMfTRFcEvSKaLMb
5+mjNT3C3trGbU0eh0t80b8SmhueeyFPr4AJEoALaXdg5cXwW8BFVR52UcZc
G8gbacNheOc3djP9gdh2MnCRBpmTITWN9eDFSK2Jz2+8NOzFTmuQzJaUEvKn
o3yT9FaKSISY1ivXY3anKLVpYQ/nk/Rl+E8AW1l7thwT72g1RzdepKpxqExg
PLFY9r9VJ2rQuoHMZcxzx5Lf2QLrOuGc6aDMmm474wvgFUCETUcKZqwoGuer
hCiWjQL2+BPtgUgftrDb5z0BtksL029ziiXyKFCB6y3THabO/AJYOlMKp7I4
5TBpG0wdZBKnEwTdmHeLqvFnMlAiacjQfWV6UMmvKkY/VnpbX+SrM7NoCWZO
H9V+a8nvBHJDWJgH7u6/hC3s5Da9yHnzYskNSg+33PwzFmIbMHq/M4uo2FmO
dkk+r4iYy7059EfBvJrebjyHYf/FD4p40I5wp7Y4f87CfKFp1Ip4Q7hwhUyg
4KFL3onFbAXnvvvdxhjU6VcJboTdR5HXmtugyeFmZ224NTUqNHCL25mfMpuv
bylJr1fXkaQmPuO7yASC/x2QdXIBWA2ZfbPMButrp1w35BgQuhVAU1kPt7Wa
29doAG2njygTF4+To2x8hePiBpT2rpSJXI8FmE1ITgEc9u4pATGafjiOjf11
kQo0LRF0BICWZFgxdIFJrsmef3MsQ03dF7LZdM1R+4FyBV6l2loutpqrcbbg
G6f3XeZ8NrFKLcJeFTnqAqRUR57djiuWgD15NOjNSGqaMITezwaZQKZJYY1/
qHnO8zKZiFSSz/7DdYPXArAyzYbHJmv5uFn2jHf30Fx2AXybjxGQWNOfNTpM
JC1PKxeRzZEwVUsd+cznp0AYwMMej+ACH3KM2YB2ahVGERoJlRQwJTuETfbl
vwjhSgVR+ey8ih6z3lE+Y36TkjaWG/N62joR2NErefkFFF3pGq26VCCeQqHE
9pveBGTozlhHRt2eVgctkU5DZHKAgkTs15rjONg86q4uYZNpkbit5Ee/AjnM
ZjuArRba7eQJI7kFV+9A3JR2XuHZ7uw11t9UHpSdkilP/k5pnnZ4aOxLtcUn
tj4XhLmC6MKwO3308hYR/tGOFvTqXdBN73wwlQVEHIl9g9jA0Uuc/F9e9GKw
kH5xk6jJAL/g4Dom5lK0hJr3pByzLfcb0NWQ28MbPEi1XwVC/kqONC+Zyyrt
kxTtuLVFJ8vqtQ84jnpIb16PCTqpX5fIGXK0HU2nkME2YP/tYFBiwzacCVqr
2Pl85uA7yzjFe+VeIcLQj7UhOS1GfVlfeDyfmQ5cpkmm4NjJ2yUMv2jEUhoy
AuPnA8tIsYO1QjAGCVSShCwl5+yVwmSdR/AUJdCe6tHl5McVk0+DIh6UUz4D
Oxh/zEA8DdfxNECodg26Mok146ONk8BpNXNgQd68IYxayo/B/jN3KZZvmLHV
EPRDpMW5j3m9lSqd0DxvrHI7+R0Xpb2hKkMIv1lt6qec6om3O9+gWCy6AAdK
6RuCn0LYyh6J2njTeMXraHYvkfR2vvZ8ALWTUwM4MViBewA/Qg274tIjrIiG
3VIRUVFFLQnAPsQ5hnqGIW0TEgkGVNZi7L7aT8MIVDTUTMYZP8iyfX4Ed0FY
o7uvCNW502Gi4UGTRyFuD88gecdJTt2DM05qYJJNpZhQIl2/sbB3P+lJXFIW
XCpz4uUDDMaZmJNFLQfJF99wEoOvTyJ5Hx1NZx0qhNVVgMZ4af3QeT1ZeS5L
GVKgeNgKEAeQKm4Nqa8ULM4i9rlqvNJ7/31WHzXFLwa5REATkoOm5qrWuaIj
rFuYnJW9dPPXdpqpZQLev/fC2v5an1iH64VLhfGZCfDmZ7BlfUIlpGL7eSOq
dbnI+MHjxlUFeUCms8ZYopbPalfXPXsC/be97utk+6u/9le0IJ0tSahqeyuD
7D1DM83Z9K94p8MVWWVdpR5tD4oiZuVRrBkXhNI72ykJ+MvNQw9CvadjbbM3
47pOjHq1DQKeNl0DMHhm7JncMO4NX9kvB2YlB20eKbnoLlIEXYmRqSx9n1yK
vPZjGilTzvAUOwfmp828KZE3/pyPClZg/UKAR/gEzKhh/U1ISCLSzNcXKhzp
OIQfp0VuBlBTmSUn64gTVAvJxqBKdj/xhDSqHnWOiKXC1/wCD0l/QkyuVHrl
JSyn0vSkK626OuVt8zPPKu9j0hnh9gZ09N/5E0XMtvNH8xiBQYIem19HGwq2
X+i9HaMj+MnMcN4l6kGnCMTB3XE93RDdjPklQPzN/g/EoZ2D4WKSEr/J8M2l
vmNpdO1o9MbQLFpxmoE7FD4jiEjusBJ4Jcqc5Q/XXJxnhU4OGslLB1vdDUyQ
ZwLa760WhNi6tLGM31wf/rbWO0bFU/0VbxzoI/1Xgdb1IUBf4CVDrzqegXIo
d2JGDdIid6OjzbzmIG7jH51TngWXQH/uCwWjKe60Y9H2enUnTuAex7oEUn+q
NnGOeU75FGj8YSmy/KbYkTWGHP4Yl6/D1BQi+zrRHDb6PyM6i/fQn5xWBOn4
Px4nGWBnG4b8Rbri6GjTo4ZxdW0LtQjBaVlx8ajD+uOQp/XIfWud63ACEyf8
x+sPINaFHqbzlX7J9UdYme2TrNUnJtJJbkSGpennO5BGva/BAGRohCzaRz8J
eZVnf1M47v0q6I4rsyzMZOBDFbNrsmx26hrsXAdSis56C6LAOTooqDprjrdl
S+BOXIOHe6RzGMJAodEGv+BgzJt4NvDxMjF1/1//Apo3rsIY6ojdx3UZQPYj
Nyy2XaSKd1ofeW/sCt96z6xYF9U32pY3h6VvotpogFcpVQLb6IWSRJvpmTDn
UXvjxXKWM17zGfVArCSekPd9do7H0sZQqwyO0+c5k4AQ0D6sI7oJlBJvBvOf
Fmd7OuM/V70ZUSo6SB8AsZu/w37llT92K/PeNWlwM0Mh5HK4KLDiadxsexxY
JQ+3eSOnHKdKL7q6zbzHYmVaTzg3aqxKaxr+F48RZ9dl0gJ/GHrxXSYRWBfQ
/LZawCSwhCngS3BWey909T/R99RtM68RVPTVYlec8ltA7ohRNsPa73DiVy84
1kFdbggTxFE3l1ox51edIN1Zucy/lVevkHQqPcKifRbLzPja8bTgybOcRomO
QMtwKJkmYPN9ALKtwQngEwZDshsFMKNQZwXrXbNBJlmrRi+b8fHbCxPmmYEN
XQVbfYU4u5GDmyKafxJ+FrgYnc8+uVkVYoI1/5BOBJ878Fe3p8KciR+VyIhP
FMluHCOIltnIGgFu/8aWCbtfYQPw+SSMUCLOTi2duFxN+5IV4zgMve4bXgHQ
bGrHfBh/1X10G55WrfM42JLKJXQgyuogaK18AgNwruk6Wxk7dp/Uz9jeiINw
fyJeJnheY44mbouLaAAySmyoH2r6cG6OR4OU8IZzLkncOTkYINpYjXEbs1bi
CjHCWLJHYWxKRL8yDADUzOJnFckX5VqEnzKAs7aUWQttsLZbx6kK//pQF8Ox
Aaea/4gb6/ccZsY/g7jQonWh2TVxEE31H1Qmro6PKhZRbaawHNcy8Iq8YDo3
ax+dTaFLdLszHhhLvVmK6+IDj1fiyl6sM4+2nOVgLluAJeX3Dy8kc5VALvBd
LWlEHKivu1vcpu84F69D8V/rLdOYGnv2NCtnc2+iSPx7FlcLxfEpSbrCU8v5
m2Z/kTId2JDn1dNKS+ijkojQok2INNFADi589CwORoOdnQggDOf40j4n4hna
fM9bmAKNLBPZ2+rtLFXvgQIXBgzVmSe+uXDnt7C+IAGS+be7Xk1YR/Ruh5S+
S++6/gmRRK+ctZYYeX48+jdn4kAdqOM+xO4KT5ldKQH/i5rcRaC6ItaCbrUd
xp1N53bebXnBtKEk55mz6RUFtbuno3yJmMmSDi62WdNZHqBcdhqsJ/x9pU8D
PRW1F4JH9c8FXPTqb6p9jFLePPR56OuiPF/iZWnOrsc+BybzK+cWU9r6kxnn
uUiGqtsVtGh5oNPA8Awft/3USMLJmZkHJtqot6rjyyqJfwrTMwV6gkrIaxzu
J/V7y6T6Z0KTwisBUBxF6cjPwJZWjt1gRXHaKP45GENoTUZHvwyvdiKxGjWR
hfPZsVT6Cp5tuocEFbLZCNg0yCpxuPlPLVSDEmbfaitC9DvZZr+4uNrZq1Gi
sixSiFdQ6mI0H56NpcWKdZ3uXHKrKC54D+DLzce2ysyDsGQ4JikpgcM7S+n9
+fqOIZ5fFgTRuzHwuD5W6MJb4AfAIPSCIA/q5fqDkDqCc+QPkTIo+U9JLGWz
TGewV9vb3a2tWdZPqmSP8kA75WjEnAJlYCd6zSiX1ZyrXQxCol4nM5aovf3R
l9U1vZBMpLTE2hOY2OEAHwZFdBnKNg/2d8w+deIt9m5tlLMxyUbjUiP77ASc
hsNbxsmP5OT0qypu600S8kVLfVec8CaUi8JK50E0VEwQMc8tPPUhZmX/l61G
T6eItOje1KO+nEE4uVYAsw9RI9kXhFIelhnz8G53Or5wwNnVfT6wnC1gIN/Z
rhDXUzdnXq/oki/2H8mTL1PhTInUierZcQIY3bXP96+7MRWMWROo73+sHzIb
10sFKh47/97mUz7pKSofk5WaSZnR69WWr7f+1jjzCNbE3QDFO1ygcHR6S6J6
y+WG/wUkeGoOz9ZHA68FrfFq010bcp2UPNn176xIoQrp93vGLTykDbogeXlX
temVdf0SqK+t0B2G7mgkVjYwwrUNSgSrOAaoJMGSuZkMiA2JeQ+TJTIUGXze
PfN23qW6hTr/Kus7elzcxI8tE7qsyXBkKLYKDAM+LjKXmLuaQMmfZOy20at4
fjvRh+wMJEmQt4sEUKGUSvC73krAGX3e94QjJ9PtrnrNEBjqf2tDgWj0a2mY
nbZ1eBaqnLXkZkrCb5/toLsAYFC/AqYlGeYdoykfcgimTByZF3G3mOOmRNub
HtMn1Vtcj9oCyuMhN9baTrOUEidre4vqWw9QcPIJ871DC2mQzWv0Mu/6pXA6
bZq5+UNYjaFw96DEHTqF6nuU9m25K9VFVWnip7uHj3HqxJQr0Jyr8mH98ujP
hmFlsBWiqFyRcTUH7oLKa0kC9gdh2ifPen931HhjAV2vcN/xuNoGzUSw+q3U
6wlylbY3N+iwJtkOEQbofsDpNXPnLDWEA/yWlPBiosO1Yeiauxx1VorQwkXj
G4ZxxV8/D2xPm3CbMA7XTfPRcjrlrSnWhS5Hgb6pQDj7PR5vE6yeXINkO2UN
nNtLGgGOPEKhlxfJtgSjI1t3GzF1kktDeTiCG2yUWpmTB+WZTuDTR1GlVLq0
DuqeaYPqZtccVfbUnTs1EMLH+YjdTkczQ8zosgAk2SE68unrfLG5u72mEXGt
q7Nm2GcrVoXf7vlvl0TA/tYxQsf+dM9FGVGvMH2qaJhEqoEQJNTulWHB1+mN
w1XmIBrhp65dNGiqrwcE12Sow2tPrrRhi7cUAfQTwlldx3N4crhpGqKZIV5h
txW9WCjFOovdrT8XinLjakOhw52nJpQO9C8BgKPFXd1FmoT3aU7WdaQQmZtm
8m6chtwa8n7TiFTFa3Gj1CPsgOt0jsoLPaRlAh/QwEHV01gdd8LwXIoSXJFu
PdS8NFYWcqwdIqLiPaZdfz6Mvo89P0Xg5ZYqMQOkSTdrwOqHsBtds456A9iy
ufuKQgGthVhdxnHpHvuajMpUVvbRG2bxvi+XDV6pNRhHOuRBsRAQG7MbCflp
XF5AcL+bpD8Z5NzxB3gb+KnXEQDBe+PXKSqemYEsu0RYJRu78Cy7J1p8PWaw
+g/nLACYidH9gWGrykMjkOVsom2dD1gbqKN3YkB3/WExYomMGdsHrL57YFYy
Wh2MjFiDOyiGk52+D+K0boPLKMmO4kSI7nos60A/mX2qi3BVJCoYvDcE4RU9
ax9nhMsr5prhyF1f5pWN7HgOecoI2Q1j6TsqPZqS+Dl9If0YBpRUO1+w/Bif
qBPBhF0ITfApXEfq+mylRhUlHIaI4Q+3YaAti2fnxV6NNyBVQ8XgTy1IMYBn
ElNvpWuD3Im4QWTccJt8FAvpQNpCye5oNkAxnMxWPHqUaqUL3MNAourlyZzp
rWg/6u3i6mwkmYyc4v5+yduTnnDr4mTzYc0MhSX++prJZIhIcxIEls1/r2p9
5pCqTWzPxUb3Am6gJo+rTu4uEnF1uM9vpRiI1evIhXhmerJIu/ngcsMj7OiZ
J+IsTyvQn/mxTuGAoA/MwEdwK4GNAoFU4LdBK0bmtksfnqsMcu/EA6RZkcTH
8iTEX0LmjzQfyt5RwCUZioR/1g17Sg8MOcL2wPwiXNoL43LY6GpFSkqbA+1T
Ll7B2L5oYjfxBbhddIM0c20orvq7ePdLF6meY/vV84MVMwg9MDrvVPVgcimH
7SjV6SR5uSjab3hFunLukwTvqgoLY+8885bdxu219ubziTyIZO/x/x+y219L
esSRynO61Qi9YZA4MAOq+GQxzLVg/oDvdg7juJM6EY+stUpczziyqeakdulu
LsVwxe9dB6bNAOwf1cJip1mdFnmou6OWrvax3pjsfti/3IENrYmypsQQCpqG
3hw1PGuKVm0IbyqQZ5zKE5cfy0kPa4sV5y9QQl/uMADzKiXI2DiXRh7JGtmA
kIQGKGEHsfgcfUNKHW1q2CPGzs6wyx6JIr88WRfawOids5k3GBrBYlb2kv1m
PPYcw9cIWydm9HGb4FJF/HaUzn4bbDPjWCnZ2GA9nVBiKWFqHQd71/AIv6QJ
/uM/5AhFkeqQfflGhzlWnG05aA+GZGkjIMZEnDQROpkcyFcWfoJD+0383Rki
T5DC7ADekn1TGMPfBCL6YzliaHP9MuAUrewKHSRRSZrEPmWbHs+PxoXb+aJN
I4QCebkQFIncfP+9oIovQo+862h8vvYFOIyJL/TngAzVEwqLSQ9SySrsjw9l
hSpDtGZXjna0EwU74VIkBic+zO73B29wrm6wTOTNyB3MnCbX7W7NEDHnz1rS
DILW14BxXqApzXwMgfZYkhn+OgvpZPHFFWO7gLtThnPzjNSbwc0wWHIF91Jq
W5cLZGZSLv8TxYsYbjyLQpYrbHZT0f17qNcK2oU2nIDvvK8KhBdX6Dbvsrrl
Rpk7yOGiRN5pFzaWnfz83LrNrr4QZdU3Lps+fIo/1QiYpVsvEAwvbr9raysM
0UOubEbg57O4s54mMQyNVQorXRoXRPRmswjQHKQkMRlWJGjwkbUuA8aMYRfN
XEtN4p6jrM2Clus6Xbs8216RMyXY11zMxcZ7aGXcwty+WFyvjTW6TxEn5xfW
2E3Ucb60ARhBO1BOLK3eytoPMFwZM6rxnrSmdN2zRd8kqE9SEIQ8s3wosE6W
zUNuMC8GbivGu1poSgdMPWJMWBwRYuM5D9zJksI5fmBr4Jl0S1+Pin3gkbLp
2CJv3yUO3KbJZw+Ld338TVkOPtLVqW+eV3Wd7+iNrC71DzgWf6kjR56LnPKw
8TlL6MPpqhaQFxCVPm67Uw8AkRrH/24QLJ6BFPIizuxRzOWrvjgD2xaU+x/y
Oi7Z98HWZmKQJ46LJcT5uLuYb3MYBQdU9txGc0h7DgYnZHgpMMgw5Op8M6oq
qsdCKi+GNz9GBDSibziZpeAn9ZwsUMd7d+F6TYBAKO2/8c7Mb3htMUhPo/3Z
ucWR+9KFm404xTrBbTwbCYV85qgKSpiS/qONrRdce/WEuIP1d3LivFnbWEvt
j2iquOBzACG6EV//du6zmHSf+Bp1frermVI9Z6mgVHqyC+EUssywIRjeYD+S
XozRUlf5W198CaqKZJ4nhlEBUsCiTah+VE9j8cW5Ky2eJSgGtHiGoaqYUJk4
7h3Wx/cHvzWjGt7KLFfo7f/0QziRxNIbC5ZP0DCHVISvtrr/qir65OV0sp1h
q2knsAtBUBXsKTjzHpPLcLVIE9xY0PACOKusmucnmu2VMiT4+FhgqioljSCI
9pX3UlX5uq20ZayfYFbyqvw+H1IGFyKQJofcIXOtaxAzQTVfxPpurVY+yJs7
EARr7AM9zX5Jygzt7RS08bJ9UKBWlHG08LNJE3IJUMhmAGFhBGJBaW/SSH4m
jOo0opZ0Nhef1Zo1nD25x3NR9zqBLA76CyKSm8zP3vYqDQt50R3aLkW6bOem
q0vx/u5K1kUv63w8y+0PrVHcKnEhTH4NliK35isvBw0WPgy4UUwTUwsQdDi2
DVpZXsh+Dxp8QdskD3Z+QIYkNA6xbW8oFGzObCurgU7vAPzvVAMfKSw59SE+
Qb1f0atQFyu33tUf4//hLPPxmaclFzWw/sqjn3HDRoQ5BOyEpIpN9Iu+vIMJ
0E6O6rlfCLpT2NLQLKTzcEHRr7eM4i8QOQ5sEqR7hp1maHM/sbc2n8e4rVVh
GLIj+u4j9aKRyV7xk+xqs9BbtHKgxTvQrzt0ur54kemftv3GZRe7ZmMpjsF3
Ah2M+Wwsnsh9fBTva50lwXdQoVipnOlUi/Qt1fg7lKZ+cSLRsKzKRMUIgKet
N4XfrXF0ef1YJO8hOXOg6sBRBUUQ0LVBY/7U4lVndmranQKoEfNH6c+Cww/k
cV1d+96ChqifzRGtxxFHhzEswwLlbF4ePt9tMe2N76h6ozb2D2M5/wf1ItPx
CkcusIpaX569OsyodiWkl/id9PWwvYW9vhCG2J5+AAGPJZcGgqkgMi5m9m27
gYwt6loiPFfH6vOZIimQbM9dyynn4mJkvzhGPnDNUgdNQ5BNKQvCihWZRHhR
FyRL4Ch1dIlqE4bPOhTeRcMFDK16fe9z85Nt+Ydhdh17rzeZBDsFO3GLIykg
Su/Hg9s4LaR/0wfdUjgd5+lzYDVT+1lVBHAumuyJ79KnJxF9GQ2B6uVmhkRf
57Ex2kj9fl+UEpqSUlJ6iohKLe+lRA930FYAk3W8pX5WEFp4o8nuCUa/05ie
G63BgxjhmD/aAg4evHlApvhbwzX9rZFIqzVmAh5fZk3aaydEq8PNNg+tDkUY
D1FAHe2brsiZlpHCY/JMiuGfxIdjBT/P/KyrfIs5nWXIiBCAxO6xOVQBOx3X
hB5EtzvCa7gFki5zn8xcHsp1mLbxhE43ucnUTVFWmvocaqX1Plz7YpFDdmA6
rUVegkOwWnYTSC2KqaZPgStdJ6QcTC0iM5LfEYrowe7pERuv9D+Ck8EnIDEu
VlFk0h+6ej/z4yCRIDCJfP5mufOpUnwPPoUOONtapLmssoCC6aPLFfMFjIon
bNnbtmTwPCjnF9cCi2kSP1r63qmmEFdx73DuIqZkXCj1fgZqzxr1Sb2rOh1p
9oQLpZ1XoXhJd+SETkEgOVzOq3tC+eWON1bBc6KMDm32EmUNHNSUSvE4OK/g
i7exZ64H8tN1+B0/LaVnP5qkxsFmsRTsVQbomo6tAF3lfj1snSNQd2zLbN/R
UHQWHarRMbLE+cQfz+itEvHYbdSbMAuhAkk5Mc4NO/J1zlSLwRQt7Xom2DaQ
IUg4epdKqV5/VEWAFAF5Q90igRzTESq5/QsVuAf9SjNWnDN1Bs6P5vutpTSk
SypKhOzO4hyHZIOQjH5g/uAcypssBN7EFJtFPftWLY4an5PJyXJkSDLTpCV5
rHgtnahnbabOUTAZSMz6dVCFyHLsf2f7McTXC5DK9MyT4B3ytUoSfGCU4LuJ
Ynczd5/jinGqFJA4Y1D67iaZo1zElHzYN48h7bm6M2nt4wYH9lSmbZA0L3YD
0Ldajw7bsSzEG4gv0xQcitZDlffkKwYvcVaXlP7MiFXRKZx6vl5dhe/Kozkh
gwpNG8825/fhiT0Mg0Y87ALKpvm18/eM/2W9GSPvubTMydy4XPPBnFZiZIC5
iG3JipPIZRfCpY02CbeK6Lf93CilQ/smzm4o6bcXTccKzqE6wahhjvRVOO9+
5uB1h39jTSUTX+x6dNGdd2i0xAOhTvD3YvptEaQ34O2IKy5B1V0S6/NJXb6V
PW0cIecQRVO1mA9vMAjcfJWc4lJG4bOGExpGKLCVtY8CX6Tk0m8EHe+twY+q
bMbg57gpcmhuWTcExsG/HfNEOlOO3OdkISUJ3fVws9KPfhM7wEf1rtORMRCV
V8awBQdtRB+t/0Mh6E9wMUe60Xep3EneRi/K2YN9ojiT7mkH9jXGNAPtnevR
fL8D+D/sHhLlYJm7INCxEaJO3aR98XJxkmMLFAJ6mNZgRq2ZbE2WcLIfdBh7
jSwYIFxUDjwsjrUNIQLIWy+aPgwwmJL0FvFGV3i8IMqsjOyIZNPb7d8IHBSp
1V3vb2dec23oIL8VkT1PTrx/bSD0d2rAc5Crhq1UKsFvZC+wSBRygiK7tX+i
B6w3MQ/UpNsjq3ih58iuksLP/XLyyALnV32zk17Bv1zzr+fHtXJHVGf/vwZS
JukcLrLiKEw/2iXYzcaZVIxUN0e8EadY5tqMdshIIa7Og34c4hNB4keNscWU
HQb/8ngKKia0hB7N66HcprpMqDtakM49EUN6YJQnagvOsQYqGQv9X5r2fgCR
MSQVGvTreKrYKFnX/QsrHhzcLD0ZkA4gqUNJcjIEnTAGDcj5E+NiUxglY1gK
sALxiWfbTsXIRurJC/yTKjAt9dHoLk9R6b9VtWnVdmnNJi4K9YzUSUVZYt+O
IypE6YaxNuue46FqUvw7j7ZzXw4ZUSCLt2hXI8PFbpHW7SfbQULIPtVTzm7t
Nh3s9h/M0E6ZizoEMOKapof+3nUrHMOsIo57g4rUJ+FIZBg2+72T6xutsA/P
/XBdKf/ayxhDh74h52+wuGZfUHl2XYbkwKBzqXWRH9LGLPLCJ9P3Ky9q8C0b
O/iscT/+IGk/1acLJ6kDdRKveMJaOYnGM0wkzdPu+tbfRWDgVOT/OUynhL0d
oVLZD4Hlh/pEn4xWfYZI2nu4Mw0PILm5KeqFKMO3Lkx1Ny92aLYUvffW/qUe
xtsy8VdyMjrGkBGO0d50l3EgphBGG1imVbsRMtUyyFxt4gkoVK8TQ2otIDz/
q0OYysNEeTylxRT4Hp0t5BGEL7nN4uguZWKJd6CIE9rJn+aozAGaIpRoxi+n
61QNQNoe6tJOLpc3sqgKy3atZ6di3JOa2jFbwtCFemymfuYxp0isVjM8romE
7jbJjmIKrcvfZH6pJRngSvMuB17/2f//wPLa9qg8YOygUKzkkSxD7zYoet+Y
ArIcQVIgA1NCb5ZSpk8O+euezbMWjCxVJ6+xdIWBGoVz9jIiJ7PiylWPYL+J
CGQcZH28JSmDOT5OfbqRw/Dwl0ahspw53fLwkHJP8Z8i88flBiWKYmpjomRP
nErxfMZNqFkb6NdvkzfCG6BDQFx2kVcykELACkDkkMOiQL1myMaKfVSA5YKR
HlT3lYd+kv68H+JEMX8SzFIZB/gqR+kipOsu/blwYqMHcCVJgxcb3RKDJr2w
fnYbuSzMgICj/UTjn4mE2Yrz2PPa5ovX+K2kWhssOct7vAvXdFx3R1behbkO
cYUj+VDIXHASbny9h5Mpm2fYs32F4xTJZSBbGp65BZPgmI7goYoYAC9omewT
Reg8yYjzRX/lI3glQEMIRUpTdUDLaTE1Z61I/Bzu5CA/Yk+YR7LzBnDMA25Q
dnTyqsxtp79s6KUhVj/5bnEDlncE+P1tK/+Fxs8+/F+BiY4oBm7EzuHizTDv
igbYX5pVN3GsGZOEBgJ86gb3YMvzXE8D5FNvKgiIXUBNgL/Pp1Z9AR1dHzoQ
dnzoJ9+ZJkqB+85X6IZeZxIOR3P9fScIDYsZihBnkuLNAW3jJPonCXbWnash
atP++juyYbjtoZmE5wXdgxy5BpKY23ofQe4kGMgJOHwg2dWjJdcuC+N6HqVz
MLB1aG6YeFvOlzYLzEG32jhaZkbrGftvlJ4Pbjhrj9M15wWLv/49snhhbyz/
58bP7936+zINk36nHrJGQOVXZ3Vyh0sWZErUh2HnRPixMbn7CyPinTTsaYKs
hweXfJKwzkkQAJk+Rm+tmUIW+s9o9280kUqmgQWi6IcRHO5bZY3Qkl93pWHk
HkHUrkSz9OdbSbNwGnBKi3mO4B/mmpa0Vy5ovG/Qa7dS8HFdp7qvYQ7bbcW5
G4kJ4P5UZoPKXe6mw7zrfP9LuKUcjvX7a2Jw+PJrK/R7JOc5n78VHTcPkfrv
oGdb2BqNDWh5a1zgFpcBH0sTzu/aTEVnwUUF6R/ozVkER3J6d5ZIy6nK37xB
aOJ6UX8+fXgFi4F2MRTfRVv4T/zYZn3+APdTgViZeEqi/5ChTXX1WFFoZ1Rp
Qp0MU7NBqtwuw6zNWr/zoM/36sdHbz1OngEg4Kpt19hE3d/TTAtJ/5Xr2k54
vl1J0A0W+CoU6mm7ikGFQ8SyDenP6/NYZ/LC9+YzUxb17p2sb7FnaBr4x9fm
6JFRfGE7UIa0eCcFe6ngredqom/Ih2hQEZjJa4PIP2auoBA3CMvBiJWBoJYD
yWBeeOYQ7YQwgYgIV+hMQXpK3zCHV0tQoN2t6P+mXCN5hnnoYj4HYxVyPF3w
9gTqe/PgUsOr692IYNGRPkNLskL0n1p7rBDkNtgWks/bjkX+5nwtV9qcijEU
PHDuTC+8gF2MSY1d3prG0z5olF/Jx8oXOonmKMMfJvuwX6YbW5ESWoU0HIGk
wUOvnapgANiZK3v1rf8Ka16D2uy77oWNTyBFfTLcRPynrYtiCd7jD0D+2j0a
TmhL+yXSj4Mj7Vo9PtX3lzBDGz611DSgxkaxJYNrCt2vVJSf/0RvGcVBI4o0
d25q2lD6X0JurMukdBaVJb1F/dF4TKm93llqwwPxoJLwq6bo1784teWOwU7p
g1u1ICZkhAPXM65d1Msa3FzKXFvzxDMFkO1z/2rSdKUpnHXDR6YWIbVv87Wu
vCL44txn67ig4cI8qZNFu1L0P3nBaseDrhkC+eVMYEDDNSfeAvBfnZWmPZ55
2wbGcSW1DxELznjuwDUSnVJ2q7vZreOkoHhIOxp036EGYsRaDq6UIcd7AvyW
wCPrIoTWoKj8iZWzfK6q/SVK3MkWgnQhLFZHTuMj5XwH66JPSTaBRbGKObM4
6tbd3ZZjLAD28/uncnMMqSvkeB/c1W+LMP0ct42S/gSnVLuFGa+Aj3wO8fhn
rwFwGte89kEj8QtN0vY9CDRSxwEUszj/MH4iAV2Y/ytN8paFixFc7DWtVafj
R5mR2CpJgIJ44Cm2gl2MKwPROSAaY6SohltT/zSY05VdsHZHxEVHnSJg/DzO
V44Bb6g4sBwTmvfDmRLSR5xzojtBNWBtXxBaMciLvdWR4oBtj4Guj7OU0tCZ
lqOlSuefKeKuJfVyyEh5swZxuPETKaW7yBxY33l1eTBQMbfB9QJRmKGtvdUx
d+lybG3JOM6IWArGbkBnas2hl9S7J+7eTFxclxniaOSbxoUiCcV6x6/LKGfg
h1FLUZy17aDjsPXDsx5KSXWHNnZhl0+pl1/mEFz5B9xkr/A2P//9PTg1odvD
OvC8SHvbRrX2OvgXYtbady2YMcAkVJ+7vYJOqnbvv4AIFnkiNSWOccMvmLKa
9BfuoogwLhTume8hz7EpvRXB2S+Ey7mHXmZ2zwmX/T1sVHuw/DNWKN5cu/Uk
D/Tx5/hfzXjF/Tbdk3JoW7ygT/1FVJzlZ0+HRLFb9SNPNjRgI4WzzZw68FMf
U7YZDGfwRBtTXD4sEDHvtpn/v3kQJ822Z8eBiJfiFZeqtMWP3hu2YhbEHsAM
UKb5NxHwpPPyjBjlePMtNhLtNMdzO3rQy+1yVPdrySUZuT9vaVWyuftJ7J1T
qKpLbvlgV6pxS06AlEQQe71TICREnVVtPrkMRuIUM+2HAkr6yZ6L9t3dwvLb
Adub/etu06Vpf94kIFk85YqCPIipRi2pXQzq59JwHx96fHdh6Zi1AhcoxWxj
bw1vUl+hxF/rBWRDK6n4i1Vo4AuCj/iMZjZdpyRtQ1fJq9RPvdRO9DNJNgb9
ItJ+uPffbA9y0gLWtoOzopYhUCdUnCNQubtFE3NUGFKQCMq8vh26MVY/fZ2f
8FHzFmFdF7EawxoxhgA1ioY93ixAvSqzut6Fw1LuUlG23G3kJhawAjfnZZke
Fh94IQSr+BOnEsXc2f4xoslhxffE3Wanr50xm1OU6j+tdsGfdzIx9Bv8flXG
fKH0ZozDe482CIDq7WwtLMnUWoD2RVVNlMeceKRyi8TZzUu0djw05C9LbApR
+hsol9wFGwqKWofrB24d7ZTKy2s2BAX0rcQnF39GqdQ9yq+gy/lVVz7KZ+7/
RR1AvQRR81RtZ+Av4LJKbG7/Q8oPn+k6EMprUcm6RFCecY+dXHiLQxOXWu+9
ZNU/WmE+TwaVrZAEt/gVFxS79YXjFzT8/OEIb/nJiK2EnURPS6aODR7h/myT
oklvSViAl4KnIUvxbM/TUAuQcQQAB3zznkC2QHY/FubU95+sEHYgsWPgeAIM
d71lHW891smwjBjwcdcwUTCL+ie3wBrrLRpTNvoq42rFKq42amwjPE0R84Oy
oPwYiVIvb7n6vvRqGZH/oOTopZRb2ZWye6KVxTQ062Bk0vf9vlTq1TO/lr71
U8/DQjFKO0IHRKTE2aZZnYLCDp3niJFv61ApoX08FP3Ea/yyGEgHtkOx9vMQ
6wqlIhfOtgqDc850WVLDchawu5OQ91GjaGOqEi4C+U+KegAPh5qF1aF8JyyA
iKVNuVE0FT0AyKk5+mqs4xvZTKDpjxYgbtAPMHHLG2DelPkWBx9luHeYMFdx
svWtbthh7uKeAo7ZaQP4ultJo0yYYtZ+Q5piyRx1YIXeQwT/ykLf/12yArmU
Rk3XmNJNvF8vrj7aksPEfBUtYnXMQW3cKUCJPrZwzIkkvaYG1AA8KxBZBBj/
TQsp2kgzCo8hP9EFLZZh5YC18YUwPVCQ4KxHyc4quJ9mFtOqgdEMJeF61/2H
sWXUt1SouDoNhX5NKKcyQbFPaX73qOAXj1DDsKUMKroSX0IKVy7olX3klZmi
xX+zWVIGviMgHHyLD0Kl+oQANLveAxO/jUhpQOSj1c8l+HU9zsHGC6YOmToK
+UkUJsdINfsT3DSbnZlNhF+Vq+TPLsA5B66LDNwzNcrSuN2iNxY7dl5mVZzV
mgpVefYHElhu+rpmJ6rP2nB6MZPnHsIvOeMd/FuKyuOxyguWEe57jCqOrbZs
Rti2xx0746UKh1eGcV/E9pQ/gPM4EmqyKSP2AIM9W2XK3/J5fINu9WDwMNhR
rJnNDa37qdyGxUE+W5+vAIZyOZOkRmGa+M8e/+VnCtv+6NaasSCMk2ZKH1md
YtoKX+2NK/M+tAEiTtAvWKA/b1cDzBFuwdF/3f99Sc1wefytQ0hBJ/UWrtWq
rTWr+sgrmwAAYA6JqnoNpETs5X1EjE0LskLxCaaUHL/Leh16yCCNo4bgn4XE
2iVLYJEUKHJqxelW10TQ9u1IOpXP2ZTzJ6mc7pVbMEkwoFFK8/cUgWRls/0d
lN4azT4kazanviC/n9/EmFnJ2CRCqfeZlo+KHNq5e8XSI02yKnrdMEX8Far1
oVJl2Tz1iz+mdZGOwxfd05/Fa1JXmF2V5OGmLMVKhSThciD5vpnzMSI7yM+r
eqXcsSLi2hyJGN8bzCDJ5NoyFHf/HWJn/69bIz9cchuDGtREqEtK7hpiYfDk
QHts2ztxPXnuyNSyk/WGuouctZ9AqAfAYud5Idk5t8eUhhJ9LpKKjGhTEOsS
2GIpfE5z6rLV95NMwhipz1DW3dUmNs7Hk4xNs7YCzp6pdVmukqOrjHY6Dynq
A9dpfcezlGPoSk9PM2BtAHV4K4k7zVJjxiK+UrFbjQ/M3KQVRvGctg/W2oTM
IBdBjNneIbFH8sR8py4PNdPu0IuCkMz34PjNNb4BdELby0paLMCC5ipHkvvV
FQ4UvMNokw1KqzWfRguRE6VsrfGlncHi3C1sGuWezatFXFhvDltc4CvCU6nu
OXVqg05/akPaiuDSr5Nj9Vfw8+l3xjmOpy9rG1sZT9kdbHKywiZvsYiUJLxV
5MhXJKWWF7RODfpZeGyxROHjXV75Zytjz9njubjQrF3nUQ/klsrtbaOiRTfh
nU/RFmaJFlCcfBLSW00ieajB58xZSH8z0v9cI9tDqwpshkQRkwTz1rhPiJRv
dL6L5QwqUEdPzSHhDYiq4rEQBfV5HeBymUXv3Ps2pwbClUahShXYvMa7LomG
68gIVcin8kN2I44N2ZnY36oro6J3hiu3uxOtjj71jqVYaAOcY32bDelzyPq4
Az9+HxYnOGRecIWw1Iept0TtJakcxG8rkpZQU05NnRH30vi+uZ3kbyug5faT
0R7joMSS7+nOshvev7N2SVwSrDiGs5gonqJfBZicJQQ/1Iwz9WMfKC8Kn7bO
yNgOMseyagH6acmr7lGnAfksw25pBwf8M4X7o7uvgoKuGlh8YevxSpLNZ1fp
dk4L58PZjqDRZFs3G41BUuPe8rKQtJe+oC809sO0TFiYDxwJLL8y83tFKGjf
l9d9hP94oTSli83aKSGyLdKPqjEysY4/V2jJRC28bfeX/6NsUfmsRPaR4Dwk
vFABTrKLTEZE41mhn+8jBHOpSAdDdglBPDuH8VdXScDV/g2iZcHAT+i+HQ2D
W2KIedTu0eu9MR4LUiy0zpQehBnQenoHltSQLGXB2cywuL270hJUrsMV8GyJ
4XJXkQBlrOmNSf8ZLtio6BJq3APz1TJPiew1Lnspl47sb5doxnf+l81VA6Ob
mtngQNji1bsd2LtrS7r9ZpoBmtSlu50yxwfwSts0jcN2cYBWhgPKERNJJr7l
sj+Kf2UAiHPSqUznqc1bONJVxQEYpwhlBnCy3FuAFS4Gjr8buWOCQMP2MlgY
LcPfEwBuOXf9zABFHYlWHCuGdipgjRlPnBOhQxvLoVsFVRJJDVksz0EdX2b2
BxTck9whS2yQnpkGFxqskSHvrmVH0BtUtzduMFxp4iF3dPAZACQMkTaqK2Eq
5zxnRm6Aev7y3IhnpYbZuOSAbp2trcjt9SMbmEjsd1jk4V2xE69HQJM8d+e+
zgFDcIGXO4Uqer2IihlfD2VIr5TGYmJ128jjiUqVH49RR48RbFIs7Yhw3BBl
Jjj9k1htCwfDljwGgHoefzF8+gdZZL0A0RzKjf7xkdAUWMAy3hNs1ISx3S7u
5mCN9djnyoy4g0QsJPzFqTZXUcuz/rVSZK2EUA8y/93R6VlGMa4/BoYKGU0v
hn+0I6m6gGtr0LsKdk4zPKz82tEFqXLPpROLjO9ptLigBUFm0yq20hiLC2P+
e0lM40BQr1d59IxnqidYeBBz33KuvYn8IBt0yJQ5ED8tDUndvtRiiLibp9K0
iSc8NEuv+ZwLzgdaDkyCDVDPXdT9OUN7h0xN00IskMK0A+KhItL3EDKjtwxz
xyMS7o1EFE52vIQnu9h7vyNsUnlYeQ1KVsWWsXpO/DEm7vd462c7xXzOZNvZ
vy8rms2/N0L2xVDtaKJC0j1gvgkP8r6b4R1cGRNO2lxZZWsJqxfKwD9SdQkP
KKqE4EUyo95nS5JHnafLS2LIBWSG9SYFr479nYtkseyOmvTl8kCtWelzY2NU
IFUU63zdz5rCPODehXDc4B0uXIyaF47j47yKazWTWoH5LiplPJPxBydgRqD5
akLk3PzMiB6ag6TiIxRcMVNpWmD/iD0C6uOy+ZZQ/IcZ64JsBri7uvz7GSJS
/ldmNYpxdCid2omh/xeV3UhB/KY7XSYKA08xnj9Zl7iHSFYx+CQGH/X37NVI
+FSXsZKkl24Xndu2/AIEs/yfv3xSHeEmNseYZrWFqLwTngVnQ2Mp2vN1LGcS
XR6O31kBrdDggxctHd0UxgoJbrdM5ivVOm8E8tCnIRpYC2gy+5zlWfKPVEeH
ImrI0qDFJhInLdKMKKruXemZo943YiLJeYWaj3qmoqDqqxMyG3l3DXWZ1l6m
U48de25ituROCN1MqjnbHY3d+Pdfm1VoS82xKTxKRMOphTI7MdVEDHWt7OLv
xmHIO4oLkKb5ndQRRZggDjuMwRz/1Ms5JAQZGZG+HsU2PjdWwuGub/IzZo9s
YFX5IT841X0zqZ75xzhg72ugo3GgPu1LF7g/lfgOnJ3MrMqtMsgk37atYrYe
bV2y5P0yL/RjlzJE03CqXk/91SxCSQHj4WeA4yfDJ04NpPZZclB2HExmdJh6
7D5cMA4d8Baabr+xJuwgQnQbwceoiodvFJL2wtsftBwv4Jv3f1+xlAhA6paX
LSNNyZxOS+GgtbPGqF5MD1QnYM3Xjfh2v0CYBa5exWrQltsu/lzmWHBbmUp7
sJYOG7VnjjQEroD9dsRMZQsdkLWUNOibw/BL76iZuxzKDqX7Be+ZuFAp7r1+
5KKM+7erpUlMx6YQp37i2I1Hlgc4JhmSB++8FQ2sODaq4YrX/EVmKgOuBkO9
okDiX357tSnR3HxgjtVv2lbAQBgWL/BwRsCzBFRJADja6HhVVMha14rY+ZCA
NuRdMAHI8oHhGXYyooB7X7adRJwUo66BV38xEXQWLLyvcOETr93bJR8CMEMZ
YzDE78iuNAT2lPuV49YrpANF55aEWV5AX+EyDodBloNpidAJiYDd3wxH1edN
b2T3ZmECj8hHxToPITpo/iRfW09/oiX/pCk7h32+wlSNYcTW1dI59ahlFyxF
DsCmt2C3g0xHf85rrCC0wJ+1hELmm+MICLQStgDmZdVrAoJkEjr9PH0X/G7m
QXlPx+dw/Yd8mb2U0LkLmZ7y07Jk8b2UWSPNMG0rcskdB421RXImu7P8qz3V
E5H7/VqMLMvc7J4D1aWKRdE6pc2eOdVVFzigDOkSDpPejq1iipjH1RoIFwBx
+QE2Bcd9KaiuxQmfkrDb6dMIcxkfOPYiY1IrcQRszARMhVldgy1R3byaz1Y9
x81d0u3o7cttL3zMvhl2DV4PuUdvj2fkx82pkI/XYBMKBuxGj7l6zvjjZKSi
/VmfYsIu8uRyxacl8Xw4DeKl31LcVqW9Jp/QYr/0XW8Gtao6BJV/c/GA3ZVu
j6xzWb4vi7te/3cPs/p5XK2e8SI52hTMg05ZvZ3h2I5dpXnz1H7IaAM136/5
PtpNvHjUMvduqJU/LjWjvIoUxVG518lkW15V/Qx1PtsJJ/crAZyKAs0y9YHZ
YgXiBXnIXJ2ahwkoafUALHSrb8anELfzHdKRUb7VJK+pRgcFlUQgOckBvuSZ
7XqeMSkCQGtLfSgu+YX85y1YE7vDVfmB9ve3c7ucOUMXAiH4aaxsVJrjkyZu
NKiazqHVcHTMops/dUiXRuHh2Rs5NiPGiPp/1AVvcqVAQlfOYwD+iDz7RJpI
y/pF2cnx/2RHPxHNBiByrNbFstS7Owz+1nFZRbZ9RaIJ6EzbBTkS3/pNyNmF
7wGR6URoWPS8jS5vcNXLJJenIBecJcX9aqJMDXQA1OdVcjkfjeeC6gr+pFhi
0F845ApRupGXc+efPW0n+6UuMKoGC3LbNCI+3GaS6etdLZRzWv7A5nGDefkd
qhTV42tPzMIOdVjYESY/2dWtaTCUkgV1tFQILwG8QrZiJwmFJEqd0tduBpv3
fbeqEk5fIPUh6iNTqHGOkKH7Pz3TfYleaWK1OPke7xMcdBNsTETuJLFisIOt
3B1yZqbdE859Ycb3U5LZIe7LIUVMi6LueyFonvaCC95qQB1XjSIFQ/AJTZlq
wl4sc9m1CrObT1zJ6HYYmbFd41aH3KoujlIdKFao2PSzXR9O98pcZT+9R7Dm
n+6vMDgMSngdJ4B4LgVqEtptgOOqDAypxOu3+B6nOTFkGGJPiwjIQBuv73tj
zfGbjG/haZseIuR4oqyN8sJjppiVd7Tp6ISmfc8n4RjvLHlElXwobnlZ+zt+
KXSMwsre2fw30d6W+eu9yi4pnX1eXlEOZFj6Oy5ugQVVLljpYRXetLiyCxXy
H/VD0I3NBVPeu5fGK+kVgnDwsmjgoZrhtVVEeysw1DX0vH9jx29+w5MqIbKM
KyNwT42TT7IXl/DY3Y6BZ+FCdnyZK/G/1Q09kTFbRBIu+G+rci21il98gaGf
DCJIwPApVDsMP3sKct/8i7AoiXEmbOcPG8/BYh3Fr3jnjMCivDTLWKFhKBlE
h+3cWQhkr9jYgZyoeGCfB4/LsnHPE77MhSZSzLhk32rIRzTK1KWrO+ZDFQH1
Uyc5ZNQPmbkZWzZdKwKm9pvNWORiylkAZMbS+us+sO5yus2gAZa63huWPXc9
Q98HiyiAek3ONOMWM/4VLqPqVXkiVk5ASAxcHTXFXgr0LohpfpxZVRde6TDy
91ascEq0SmHsm9NvHV7uX/ulbLyi2cVzgymuCLYcMCAD0CMTyTIPTBzkSuy3
7mO8rcAadovSCVGZSuNATtT8Y+6rSoHp8x2S0Q3ghfIzknbHHaAOFyAuMMiF
r5qES6JjFAKdB/E8GlAwRqOPqUur4YP1Zhc65MskPzBQS0UvAidonrXm6lxY
jmhdOonOZbJwhAvmVqbFD324htJ3ORQvWjNG2BvRqFdPg6qBQkV5EMtrcG2h
teUSbm1FUBS7DcboVKd86E4tAhqdYSEoYakHpcNDnr/LNcctYtH+1nRFaEE0
gmOiFQuNqukMipreCFPf8a1Yj77oMkU4skRwQ62Zx0bYjnt8HPCTdH04n7eA
xd/AIWdik1dGm0LwREZ5fSxraSlC/3ROTe2i+KehC8Fo/QI3FPTvT53q2Uyn
7Sr0PHNNu6agSJ2cMmoIk2BsXOAasjbTpuB4i7017uOAussM7aj8PXigbZC4
Hx4qV1NlDzsmlhLIgYnAnPP7QvlTimioJOQ1rLjIGUth25uzS9WkMOmycToD
a1SPBMZ8xiLZoOWEp3pGHvMhXCFGiAiwGsoZCQSKzGHbWMJIUncWw67BXNOS
b4ahfTddjodwMKY5LO/iHoOZaCpxqAoqj/3sLW1upCm7RboCE5TYf3NCUb7C
zRzlvQc99bhWPILxx7zzyrHxAMpRDmy7QK6WOJJurgkk5ZpB7zKPbAHlvQv9
DJiYDxBAixGIecs93P5UCuB0LejJzlamtf9pNlwlOYDLO2SfwqhuvdfY7S5M
YkLipnhgblBD9oP0PmiXE5a+xG7TdG8qLE2Oezbsn9PoqbqFzeibCXaR1Nuz
sFcJi6FNg0bCyeXzrnhS2O3P9Zbf5darEuxFRb/dnv7Ymzfz2yEthgBUfrOL
2vgYohIx7CX3v7qUbkUfOjsP3Iir05wLZLDk3ARGSEetoG3cQr0g72ULYAhu
wePTvl20uPGM9VvSY/dFWWPOxADP/a2Sl8glzFVkPmay6HnQPX4eFrX2FJyJ
5PI0AEfYMz+f1KE9KRtDskhgC9ukWU8Z3J3eL2bPXGllIaQPDP2f2GLPAmhW
qzSICZouSne6BcWlDeghjm9n8pbVNcQJkGZn82t/iZYedcZzow2x5ri8Ky/U
Bw+PiapUZuc2//rPU9uzHre+/1fqSFI12oK+KziPjHlRo9s1R0wwbrinM9pW
qczRwyzUSMnaMOY0bqWjKx4IytLkojzofRUQewLTp1JqTR/ogys6Z5Hn9dqT
Wrc8cNWH22Yvy8LqzH5bbdINnDvkXvVjJOzqyKAqXNG0ijwQrR7nyJ6I/8af
smGYCfEymbHaCvb0JJQ6+AVdccMmdhs6B8Zz5H9x8MH+64pxG7b1oaZhIlLQ
TUE24LwfprK9OsTuNKKQ+sHeE0GX8SLOG72xHPm2JGrnfLiZBOXPyDy2CzM/
Y9HYDjLd3wG0u9PUFSePls8Fn2xSAzH+gCJI3ulBYmA9i/s8xcJ2Ioad1vFN
iKMvJoex4Vq+TnaPOGyNrRNnGqxY1jnxrFqfIbxhLWOU+Ej9y4UQLGhW+85l
VthldIYQVrRonn1J2njsdexyP4A5M2LFV1IkTzM0kUPb8XMQLDcOs55zL3ze
J11sbSQ0cGuUargfxMYSuVIX4Loo+N5TLh+6+GKKoHoVDv+m1/0cMv1tVwsW
dOMysWlvXSS4qsYRKPqRPZJOCnbp6/kLicfs3xfpUbLkUg1iEvBnJ1sOntnu
XUpEqIHS4wpelSC4SuT08RVzPIl1w0o9xSJJXWSwVShmVodITy+EBrp5MgBz
yO4cWVeR5/VBaARyyObNazyk8GRSg53ijsFOdayzjkiG1TpjE6qa8QAQ7g8N
Hs2FMxukU7kIuXLlfnKeIX+qR2BaE8HZJvhMGnWA2NHBfuHMff/K7sq38WVC
BdJmmoF3sR8M/lc8BU/kIS8a/NWBcuzvkdgdRdsDVw1KV2frfC91icx+wdWP
enhIm6quQMW4gIvMv01pXH9Zg/umatlTPykc6LrEQINKx4Be+dRj+l1COSXV
MlrOfK4Qsd4nbm6FYzIiGdBEpokP6UOPrBbd2tm27TvcaCbn8Q9dTXF86roc
mTcVsahoVgwOuVd6vVauWkvLGFZbL+MxOgTPNw2DSgSL5QT5snvUt6vITI8D
gl/S4fRCE7IlbzMPeI7+L1tn9Kp3zem23jcGJ0TdM3TGN4RkVJE2o1uCQLp2
iyb7vdD5dTC/B08XVWGtiVV7MHYnh6do+NXyqnXq8MyCQiHoedQIliXtHJzi
+yr+8dPH8UwjkzmIZ7gKIe5YSraJay9Upy6/UAab57+dkyJD+MFTYhP0xlsn
GSQ4Vn7hPmsPW0uyefHlw7Z18Ra7+UvPnnYfO6yNsc+TaMZTOZFj18SvjaeA
1kt8QEEsEWUrk0d8LyvRu1ercNfJBE9dddCRGUFsbDRi2P5pcXvShJJSLdJf
tPUyZrvPWDvZ52xveHtHDLpAVlPB+4oEtXAYHLurEnOwxwkUgBBscUhuFtNf
qYNwylU+LsUGe22hNg2ZOq7YKaup62zVZK2Q/2Dw3NrxSeFO8xbHcPG7RNLj
/qvKilyjnh6kQX1I/reWak+sxHXJBep4nREcCJrzcPamsCtxpGOGd9BJmS19
S1JBzEdYnratPqUb8dzzkbnLgNSpxD2e7yymL7kzA8iDyhOwEkP4jdg4QsrB
t9tzKyQYqRL9llmKsgkXEgGqDv2+zvCevSgpJEFvGN3ovL9cKcu8LPlSDyG4
WjIDNGEYwgHLikZhFSReB0VjlJo+19f7AMg/2h5pzoOnfxfpMMQGsxliWdnJ
fStrr8lzIU2fEHvyUqOE67DOiA2uBEU3hrp1/jeIQ1A5zXryRAX9YyaLRUOe
4a9WWqTfKnT3RZKgqLh1RjGJmDbeLZ+yGJVW+2Vl7P/KOTbE3btQ+EQcWojV
dgIXjgmNJTW1/78QeiK6X8WkR72w56QjGp+c9gSGFmwx0cZCx+hRe0sWuLTr
RBd3aJIxj69KN2W+9Gwsfq6alhpu9/TrYF61URuJ+0rutVuVxBatB886N8y2
MjqQoOHuhoH4wLRi+34jvbWd4UBRNA8ypAK/cq9N+YG+bEXGU1yyAB95Rli9
y911BcMQfk2GOyOrEZpTYvd+aBvyyKuykOOJm6u8FO+E7S9wvV9LFYvaoAR+
0fvRs7GXbDMOuS+mMDsHPj23iZX2zVRDl3UrKRD5IfBy6P8N8zuO/3kNRFka
xCq5ey8ckSjPfnr0RynbkCPhoavH6NCNruScV+7ikiruWSgobwS8ZbGqPhzo
n6nemsAwkZ2v8LBF46Wxk+2an0G2CgLYvZT3ImkHwz0G85rDEaaa49Hp2dBe
DRCUJ4nRE0PvaseYQvW40GA/H9MzAIpX3hkS1hLGr9TVYkafGEf5Vk9A6+8l
y8+SMdELVdQ4zv6Q/Xj6qyLoEQjgEVqgIe/WHFSmmBL5ilxS5MSd+9033N/2
bnk4WPPjs+rN7b3l0eHJimQCAl0hESgLNywOhADoUHDGm+N9GIEZFac3CdxJ
VcR27SRYBrfeYSj6A5PbanQUwoIrAobcGlAYvei17D2X1J3zdvT+Cbt2BsUI
zV16z65UcaSPeOIQmBO7pOSMEoussBUL36R28dSkAaYn/rOvM/ANp/9v097C
GwgoY3BuMS8TwKrZnOE+H/ZJGZCkTJGlEWVnMcOFzzk3l4W9p/+p2deIAzGq
o0oM+djPz7BUJtA9IkUm0pNRxjgQWFV6Q0G0XK/d4pVxYKTHxWsNaGqDuEmf
StrkJJgtykjvf8ASP9XItMBw+vgcQdiPv6IRiIN+86iPS81QFGUWQ2aV0mvG
Sy/p8ekRZQGohd1iEnDiddDPzxHAQpE402EOjFVZbgAjhz/f6xxKNTg7xM5D
gFnPDYFZUSNBaUe4FQvQ+qsw5LfqVXhBxrd4Vim2yNTLqFdnqThd7e3RsNKm
hxWYQ1eY9ULQdLE74UwFQSKjggvl0grSnfX8KrRYrDdzHNfh4LNX0DIIMjj7
bTY12aYB+eHe7LmbG8sv7KaBIb/6cxhNiFtIT/yhaUZHEBRBKrkZ5gB4k0++
qFzD/Qd+Ega/IZ1/QWDlbMhmoB+uLdNPNhQH30iQFNkKOMnAWi2JjqypR1Ak
vDgGdCRWkfYF9lPk0uLqlSlm8iNIWW8SfzgolSndlJKVWI0VDz8VLy3zcPEu
1zAmpYbpc2g0Us/nvkKm2lvxH+UTi5wrk1KxPiXJ8upIgFRDQs8vE5GeWZT7
ED4Vp5HGR2w7l+UkvFmIAyfEuDPFa4yTKOK7I/X5bbJObPHzRCGeYfr9buI/
K0fdXwZuBw0aSPU98wYI6dCirF2ZrRHxXfaVkrBWDC1pUkWzUl7mqnorBEGV
C22K3vSpDropS2v3N9b+sJ3021mItguPAomrc+LkfUuaOdWQlyPgSrnpptPU
kyCQ45ssdtOG4ltnYc09e+RmneB3AiLVm9JpvMuyudQS6KZnZBcV3z8ydpb9
v1Nr3kHbfkZmnkSuMRQ5MkXcgqVayTgcoQPo0KdqsfUCsVPffS6igXIH6k9O
MSYeEMnDF2ABlPuxwCg1zTwjzXB2nee/ngFKtDt6yp+2rwHfvLFKTvTlfMq/
AnrYSxivVmoMPr9rlFDroUR7/eFZe/YHiZ4BAJMt9dUdmGyp5Ks+6ncGdPpi
Xegqufh/lH/wffpHwdvAjw7PwxKxO4Dn3fJyTmZ8y7UTdyPNFOcOZkuk0TX3
3/rWOAfvvKaBXPx4gaplsM7eeA4N1x0/uc+KMOHNFmjIWo521DRDdY+ABiQR
E7jv5Gyd/W6FBxbeRGt3e/ohe9RmoqGMkENjAC4RAyu9IlJXmPLza/ngVBJQ
pxQskhQAM+yI6mBffa8sZtyw+fmGEiQRSxkhJ0wT4za3NWdz4vrtZjDgTbp6
S28IWIZMFA6c+lqWu3PSDNH/tpgnURl9X2g1HDb/6HVS/QsLxzBVG+TT3ocM
cfT1YSX4q0uPkBC1mz/TytcUYhwzZfIcv7CRCvxtH0Jxrc5bhd9Wmz3bO6R+
6z8RRadW9PZVkBCmfxBE5ToSTWsnnYpRBB9VcbX1U2dq3fnmAoMFXbAkONFW
6ENPJQW68avbjcPPwJFpbNv1er3r/tkQuswu74FfbclVtVMPPZl/vMwuks0v
NifWHNb3WWXp9ytX/hxJrvjyc0oZo/uysY3iNecZjfJqPsS0/Z/AALl0Jkx+
PsQGjYdkpY9pI9D4AD4vSj+4ABn2hZByC5XWNxsZpRbkYX1nR06/YONb4eRv
1mfHWc2WLdj95Y7GXQQhhdeZc6ibDc+WXbVPjz895ZkSW51VAPg9hgk9q6Ye
csRATTwTjv+etMqyNOgVcAgPpXoLgXhhfkHJQfI7hVVYRvDXzkDVx9zFXyl/
ctSbjs8PUthg3beQ+EMRss0RE3Ncpx/nWTZ+nST9M9P+yh4vERMUAyIjLw3N
vr+Cme5TLHa7zjlElLoSaU+efa1AWZqMmaB8fk2HkFOBZH3DCOHZBgTuE40v
K4FPVHfKldfpPenvnZmKcWJnbdeUzwDYFiqmJB3cN+hkHt69dVSawiCsRdi7
N7q4OucLjrOuBBOzm19D67JNxbT4WVcrEPz9RBbpatPtJPsb4A34+nuryfVR
j89pVim2iB0HjDR70WBPEZ2FyCWeFfVXFb3fI4nKNk3QBRxh3pUBQZzEcKCf
ZOvrlRnmMD2HpKRRb3gf6WJYuJ1qYynhIAGZt7wO0D/ZZgFZZviS0AKprXXZ
HlOK51CgRt0exHwNWWfM9iuhrCvhxzhLr/P54i4wp5U1ygNc6KS6wUkQ3QF5
Y2Gj83EvI5yBRoXsy1QT+HfLlqbSy8XZCiqUo3aWIvPiq1NsFDZF9Ixkc9Vl
0+eCsozbvmXIV4Pfu+JbZBO/EkK7AnkO4D/b1bkCppcn6vZQ4xP9GMzXI2O2
zSZuGvraDqMu4MoczsY9H4WW/B5+837h+JYbeWqqbmOtOjiog6HlC82VEXnu
hvddz/lhr9/s+P9+yvBiSkXmrWwdLsoCsqfNpBa4L2q21vP2UNEPD7JRRywv
paCBJFyYYXQ245fyF0zCDTmE3uKvmbzRG2ZJN1c9iJnteg7IZyBYosEf3lHr
9crXwjQ1Geq1DE0jfPcTUDRaZHhB6Mq/mY2d6OpkBOo+jkwLBVr6NlYSDWvD
ypyCy3BH4RJggl8VOq4IyvSPgfxQx60bnffV8HZRL8yfBC4nMM8SJOnl/gPG
yqFogYmAGxhmhevjBpxvJf9SN95Zdt9mNLKFO6gqe9DPtHJvHg0DoqKIvquz
GJccLmOoAFq0voMInob7zRJGeqgNTYyQ/bpGLZFmnu5hpW20RnXgpJJSD5VV
KXdicdvnrMUgZJ4QdEj6sBPqfR/YZ50owtJXH3Ojf88WCV4CBoTsMdGYJfRe
ALzBI8T3Mz4ra2p6nzDk2SCXs2GzZm5M/1mM1lwC6vVgQAZq62K2tIcHFzSR
s3HhpHaHa0KCI2UNHNk8BzqbOk6BYtLijuG6uK1974xWtfJirktgftLjRcW7
5/uLdBJlE/5sLJ2Spw/AhzhaBacl6Kcc0gQO9p82wTTTxfRVzYBG2+vTq2v6
2O+zDeVz3SuHkQ+frE9hM6Gp0MWYboQeFPjg8MMkCTLThYf2vhjPPCKesaOS
HqfFiiJLGBWpel1Je2huC1/fYb4JyLgcRpV4NscCukPkQC4olhQ4H7J63fe1
vNxSo3/xA5I4+BK+yVSlWxNbEI13I0VX2+DJyvvoqvQNxCQRYFUXiFfx3K8M
yRcAKJ8ju+nx1mr8z5/hPMh3ygSodXtnQEBisjiZ01CYBsT6P+1kAWboxerK
BjcCjN3KBvahh67S9BGsbcdYyQqHOvrX761cJHKTJ9CcqjUEAU5gqMjCMzex
JR8FFa/gLF2K3KjjOQq0/ngY4VWhYO7TeQaeBou9AN2EvxW/raYgse/hePqz
q2hT6fq5B3ChK067IMZ9nJL4ek3cf3gtMKfL530jKgjyewQ/QSJARSn6syxb
ZqKRJFCVPolEDMe52Q99ZJciZ42GDQUyGO5DaMpYC+MuLOfKf7M2YFYpyslS
M6eeLtiTW7nyloZHX1A+kTFwY38jzz0XQI21vf/sAETYQiFZs67mpOf/j4rU
SoRsOVcrAmbig9OILkGpJoLOz9PUk1VjkoAYe9kWcqRbFn7nZnr7dtwqWkOK
lJql2vH+R4gA7fC1OATrhm+Dvp58Fs2QE//An509NVJHP2xnhFM51OwyVad4
vxsCnnKYFvGOCLNse9UXQiZOWfUvttOk3AhhQDD0QRe8oyJzUK2GDjF3wPs4
l+r3Qaxy5pxrRd/YfqANKiGYoS81GWUrBjkHenTIcj8nZLiikrIczOD5FJxq
RNyuvyoUUx7aUdNc7XrzgVmPHMOEieQL8RX48hSqOCSGAgO/sozFLtmqy+T2
U7M7/QAr0c9XasIU9Nla7Q+ldh45tw8HSwtikTPnrovJBxGpvwSNXYk6bBG4
NEYmkapBR22whO/6RF2fDQ6/4jfJHA9V2CsUvUoWuBFtVq5v8CGI5x4yE7Hr
Nf4TG2As8lGT7fJynaPSYgF4eL8rpN2QpvzeYKYYrjZEQ1h7/eV/YJWlOSQh
enAvz8bXWlSQ3jCeMJXCvyKeVv5FGzBDmu69npNii6IfkaUDxrH1WmLxW6e0
L7XeARD2/isrGEnSKh0MaazbSRwJ/sA61/oqw5L5iu2U8cBAq+Ue4JBzCVaB
hEnp8S3MOb0HUxPKfTiyLi8a/AbIVX+1JCSUWW6lVrB1T8i453V9dx8J2kva
JYLIh5Mg+VX4ht+IChcnNJlcXErkz5bA6+4O8WI3faMvdtTcyVKPc2x5Sen2
s+C2w9d6R2/j83tjuf2+ewR/IHanhLZGwYk8e9DopT0g7roCS6Dmcvg1F+ru
f6HdM6K+kW2Uw0pQpIflYiNwVkzSajYPkLvO+dgSuM5RJDTZpceMTqgOC4Vy
u088TNmopieRYbe1rDcALIhU0QRu+w4BNcAQdCHU0aJXzvqJdSklFyYuzKP3
7N5668d6/twulMIUJQ5FXsiutBsUPo4aVTgG+nt6Q3k9EymKWvERpK/NuG36
RyEJEoGRcTjal7xmlOgb6NzVWidLHD+eoNKGU59FiH2rPjGw4mtg4bP8WLvK
jjFFmhjTqlHf2nVjZCDioskv/Uxs0WHf16ya6hwqAvFUSBN56fwqqj6ctjvs
vjNFX1opusltH1sTykeVomJUN7/Puus+4oVACauzJ3nXB+RBO16jGdT0YZFx
ca2+MqTJ5E7bnmYoY57gkU6Hz1ZdzkyXOnRrvvRK6Bo+orpsY8YKS+69Z0xh
FaPHP/v+V9JIzsLBHmpHNXi52o4SIXS8uBF9j5kyddK2vbAhVJrjE7pjYwkx
UNVFcD57yXWCyeZ0eNRt2Wj+oF3YN0sZBywfv7+k7j2RDX2UpiQmnXfH2lex
YHw0qgwtvli/3nIUhoXQR//jS31DdfU/fi8M4WxxU3sUGl97qfgLWEtk37ru
jPJTQzAgp02WMXj5GhXPIddw2rZfvI6/SSF+V1NHKvtgVnimqGhrqC2TA3Vt
3OZyY348Py5yHJAkesT/mMQ9+Sam2zCm0TRn52tvmguXzYzcxACmzTBpwUit
dKpjrxfFcDT+3mIzcsq5anfNeci7zzvoZK6RKiBGdMy4zl30L0jptGlg7aDK
6+wgmqxdpGcyl1k+PQS1yrz43mrluFyuLUvdI4a8IHfYAAI66PpkhahiqxE6
HnQsdXA4BKXp+toyxL+MhxT+xJKzQYxM59z3dJRWh8u1Oz3det6iygY4s0Ll
Wi9BE7xZMbPAbFjhFpCPHlTpadyFz7HD2Li5tGagHHPTPWyfMu1Eo7uVB2F1
zz+bVxVTeORE1jKClKkliQPiW/zw7Dh/hq8QByBqKlrmJGmg1sCD/hJqZXw3
wSvCzqNMi2hLOe35UgInq/HUjzmp6UtP6JZ2SAEnRE7dApDKJ4nLIqIq6P5a
z+rT1A0BD0QpwigrBfBIEXb6hWwLksCTVJiQtU/jwQltowuKYZgFuD8iCGMb
hJxKB+nuhqJ5vlSTzu4ILRyY8d6wB4jrr29A5YQfTRaLZAu3OLNH5BDts5ki
lJn63lkzZrc6Pt6v7wipx6o1Uy41M9TCVIns39tIWC1bnEvSj+/E4H7SBVZ0
EjB0qd3Z/meRXdLVbN+BnTBFBncnGK1o7rzVAXGSNaagvdPH/pyPHxVLtbAK
UBu7ri4XigaowgXPJhmmDGso6SX2ehePvLMEK2l551+zND7deHlCrzLb+PnJ
SQi+nUxI8qJrmfiJdvxV8pZFbXUGXqbry4oWa5Sn1FO7eMumtKVxhOr39NNQ
/SHPcM8KQJ5OLPq9Av9XJUSV+MPqW8xlJ43NYdLNoSo7vhYCnVuYLQNVGCzt
mqvEOYC1BdHTwoYLjd2Qibf0pZRynJ9Xvp7SzvJrJyTTWdJSkkO/hVmQBCWm
CYsXEojyofLmCNRLHBji05PoK7IToBtxKz0U2xlNx0qYxHiJguOLwbn8pUja
FwwKMf9wuk98FXD9WOi6te+REDhoiEmvt7JrnbDJe3ovVuRKNRZhdwJ0sgyu
Ym41ZDb9otV48HRPoGgQsWHhdlnvGwTpfO2Ao5w8LN9uHPX1XJ7Oijg1AgmK
vMAjlOU81b2dKHBBXqMay8g0vK2/6+Iz+1t3kXINxxg0wzJSqq3/IKRpcLml
HBQgN3MeSeiWdet78WNFW84NtLIH5jpN0wax8vBaoLIMXe0NKYvOtp+YIe7q
3ZRI/ReM2xBcGwB58cKg7yC63rXEJvkAPoIuN6G2R8oCkYtBFRBvYNfONZSP
kcXytoYu9H1C3o6if0rTYPwLK6azcKS4gjJY0yTlTIQsaShpj+yqqcRlnSQT
zMlTIMmemsbZtT99RLhB5otSeuJDQmdq/B4rZQYldADMDOlxeucEhmFzCwBd
yXGxiQfspfvwn3oKW4pH2fGKFnjJx+dz9yxCTuhPeo/Di6Ta/oHkbaDjMiYF
/cA46izSYfMsbanl55c8NKa98h168hTX2YqXgxdzmPkVfNYdn0SNsZFja8kO
a0MZw4JuospPdemx/9VErEFN4En1t/xzpcYpY/9SLjo5ZK1JYDruiAUP6m+5
z7yIiZ2eqPe0z8/28phMcBTU56m2dDBd3oI1tkgtrGOUG2T4zwQ830Wb1YnC
Hr4kIU0nn3x+gIoasGmhJso2PlJbFQY+DF6GbHkCJZzE0mxNmswDY43Adbk3
eo6zOTTPamkFYyOP1+ucdAuX2s6Y4ztlJ3CLxtHQh7aOt1ZnpUMz9QQcRAPp
OLoo0Ws6Q6tfvaYYkOy6/2nmxLHDrgNuLb5FNGmfr6A5PlbSPsxtIToDirJl
kTcwWK3QAOrVYKtLy3Xwcgl2CyOgCbD8Hsnhj1ev9d8A0l4OAAU5m2BAPCMC
Q/jxjO5/rdZCA/B9Oq8HmCI8m/0XV6FJYXsXeFkIgcZ9Dy+iyWgKx1uCZZjs
q4b2ZE6Q28pVPT5D/OG7ZL2UpCZLSFXQa7yVwFBZBJ4/vW45QshKcsr6Zf6N
j5M+T40TISI+JW6p2tcvgZYm8CeX0uJYSCycvak2TkazANju1Yh8G3mHrw/U
hjItvpDioWsDOIYcIipFJjp/w5v3aBn/ZEfLz6g26e+DFAGgBfUMglNQpnEx
rN+9LI7hXYCx/kYRuv4vjG9nj5zWvcQO6/M7Ox2T7DO/Xm3YLeTCSRXvJcW0
4SRM80CZ4hnwcoO28kc7VYpY35ituY/Acc2quErIZHNHXQ8suL2KMO46pxBH
aMTQeNJM7iGs3C9zSStvtIRb9P8uzlcgC3n0+vK+qi7e1ek+TullfbOMmdFZ
xnod+uANiLdM5uKjTq8fz20smP9TnHkwOEoW91yiqqqdcxMgxaHEmgCQYp0W
QwxwVOk88e/UtPFRXckjVtxVzWGlvIRBpXgsPZNB/ecz8ZPH/0z7OUrtVnx1
SHJYIra2yQ+7kzwVh94nxF5/DUxGjnX+a6iZaZcScDIqEpuOhI7vIug2r+QA
IIS1tBOl/fN1gzTCmA0RZF8FJpW8TX1NBQbvK/T8OMOOw6FJsZ1jA3Gh7Icl
4tkfoEXXVpwboQY7a+CVFYyBI4xG6qhrGzq+kjOrhH1T74fgvQiU8HL79C6u
SIQvMSj5pAnK+nQmuCgPoP7OMWnMc+Nc8x6aBc7JPIhQxYZsW3x8L9XFXxDg
ycHWDYz4pfCMTjRiO54cxSx8BB0AA/Q6AKO66zh+/8kEKCW7Ta/XCZ12PIqj
X2/xk837F5noaHi4JR9pPuC8L8TkAo+FUuVFPKhZrpVkZgHHGk3ZwRJjcuyL
jySByorNKaWR5dQWRZrE116SmjPLrATkxyy2dJQRC82SLvGM2uC1K0mUWGN5
wq2VTFmYmOz13pFPsle5b9qGhoNxjkxxlUYULNYCtwzChle82Odukxu04kxU
pDibmsq0YMwjLwsy1Tu8xxZrIGqFDoF1qteDV5VgPAI4yN6h3cX84HHr/ljO
rUqC2WL85KHzQsJ6QwqS4T6qtD8YsmT73S84M25w69ZGbZFvR4GQhQYukayP
BPoyLqZWY+/0DSYYjw1tH9cyOfQ0L/2z+ArVMWpTPCLQnErcw8hj49UIn+Hp
T+joeOAIrFmDls4Dn2f73Rmfj4gg05+PGXLV/28wbwOQGxexbpTgmyAa/4s2
I7dzfpjsa5cijgVOLMtlzKf6tceea0++GZVXDQUzYiGbLPmVlUkZtiUSV5eN
J7nnzdGZMsP7Z+vFTWCDAl54asdQyuysDW/BAR/Xrd8sDe373LHdKFixBAz8
i1oSds2+UPk3f3gDkjqgoLFii9O9gISGlVufVfc8k+X2Ir19GLnVcJvHkk7r
wG1S4T6LcY0PZ28xFeCtzkQtkMOTYHQSUjlWU9fFFhI017tCpKuM03bDBRLU
eZHjVUuZJwpevPTuaVlwKn7QCMv06jOtuWchkVmyKwxZ3cYktTVJ9DTQysUO
eNiBQ44S+ytUPkdbwBbbPtw9iMQosn6llBPMaXSJjpKiLigW+1sYKrgeL+41
/Z6YCtwjPkhe75+v2awlV22jMiUkgSHfOVcoMdMd8KEAtjccGu7shly2lyPr
4b7MaJtfi4b45wB9hvtDwa7pDDxYymbmqtTkfNsFoqjM8Dr59PFbFhDo0srs
b44g59Btwv2owIZdVpO/aFoAH8DX/qXcyadLyZywJt/Hnut+ylg7F1lSq39X
5MByGUQeUK/P9gD/8SvrIQBOGmzf1I6unYAxmWWxy6fNN7ckDSQo43GmMhH3
enV5wQKp9W6Kh7CS8UYJ++UWsG8D+9xd0VWh4Q+CoKGU4derLt5GKkc/myXg
3DZEy5MGBnnOfGDxREuw9uEcHPX6vP/QagUfEPI4ZCJS96RFkLBSJNGyIXFu
bkW8+/SIVHgsyskN1A1QRE8IjD3Ee3ytJa8NmnAOOOO051XUUyDFmF+7LfJr
OUQigC4dvc0mGEnssEOmIKueXNd0MRf/OgCmkT8/Vm66+AsIpCpw38Oqreas
RZouqCZZ7mI3VMRN1bQ1YFCpm82FeLbgt5Rrr7gCV9OnAdAVAeZCNbanvTY+
HBnOX/xJtVrGhqD6EG377kI+ODySVuBTzqVMlArenuUwWr+4onp+RSwwAJkw
ip9ZxdYE1AZhGST67X2foa9EZ/3JvcWMCpTwwU9bNQbfaHj0Mgvz7XqVdJhc
8yO8D5H4OoChNi4lcNdUDL/wNGQKXWPQMiHRsxoFtUIHmMj2yb8a/bC7pNM8
eeXuawKutcZGXmgpT06FqVjc8T5SXq8VsDSSQBkwYhagebDLAB7kl+NZgSpB
bXO8NJAl96fnnuiwuiYgB5KmGUx8pdbaRp9sNl4VuyxMirOSmznKgmi1N5zd
N3tGyYC1cv22v1+2JcQF/yIlguk879q+l5yO9Wy3s87DmF5Eae14BYJJKfX6
DaYE2YthZrIzhQCX4tHVPL6vGKtTr3BiLIMUQr6Z2BGu5SlMDzTlTVpPCpG6
IEbIbt27nJ4TDNiAZgfnSry/zTTAmShQxO/xLbl7OZs2AwBBwCNt37dn4HB/
6A5gG0aSO2dUtinvM+uSrCk7g+w8TjD10AipzHQo9bNR91SeRF+8fqTbbg2c
tadTnG/7rvL+aX2WysfdroawDR6FwLBYPl+eT5TsoCRJI1/n7tEBdr4RmwFT
byhw6T4nWHD+1LmsdygfbBrynT+t90xng2dnl/SdHoBAq3poDyOq2nYCSXeE
zCM+6FvldG8TSdjRJsER2BNyrr8FCIBKrPza4CLJNTpBq8pQzw9MucupUurP
fEPHVA/DlCSI1F1erBBgGSrn3F376UL5fSAq5XGpX5CTp6GDNL0UCq+YN9yH
2VtsD04E8+M+cP+JsZOjF/5GcJSsWxdTbed3t2yYAxuegZrX4U8TtQN2klpN
k0YQ//M093gu/mgjfI7Rg+MD1VWy0qHulaSazybO6FxWh+JdduzfXIdRyyCK
bzyMu0MtPw7cru0DYxWv+fUu0yaYIC2zRlJfCai/3LkMHkknWqGvhmFBDz15
TvbKG1Kq7PjHPWVFTUlkLEoyMmPhSJt+fr45XZYA79vMT2iCjlFCfiSeWH4H
28XFmyWaXXjZXP6m7NPxuSBSabJR9WUv3Hg3eb1wykzeRqEjEAUxrnrmqOT0
YkUqQXFr1gpvJy5jlV989XGi9TgmqY+thkJiv+H8gY8bzXmKlNByhGexVPLX
RkGB+iiQWl3WBGfOIJPWV7x7ml2iKY8FdSV8R/RyPFCy7YxoMSt+tacvKmG/
E/zYQbeQ0hEiOQS/5UoY3vK5tEpvctEicq7qY8OORxMSTIavo7IdKYM8X5p3
65ME+paQk0ewiCTNgMPQLyjgAn0A87sEQgewGa1PccyHjGJ+I4KVhfyWcsWU
ArnrLa3mn3z4CJrSv7tnyzXvpnD2+Dc0XoHQUk2LO6dp1HLjGpOmn+orT6yt
71VKhC4R8fsdalHTQpD4hDcI8ZU4wmdsfdXYwrQ5sNXYcOC7GTC1hnftJ8lq
9wSFnzfM/jBh1P7X/586alQvoLW8YR1UZ5bCvUFSGC777agHHtWC4oWLqtBk
bQ/1VP9oxIDBErKcwXNNJ5P+Q78i5+6ce652IrgHY3CrtTqiE4avv+/dGGDn
uG9HntE4Df7PvXMhqsXOgRU6/JmOeHU2KcBqjAFxjrQxvPxWpTnpuaO8DpyI
h3yF6RbrrlrXmNOGFnxZ0nhktT1wgdV8GY+ooSh9QY0V8HZJlZ+1uU+ORLpp
TnFYnejc0QnV2kK++EOET19gnWRw6Ac1YffkXZt1Xght3iOkPm2VZGI2sKLl
Za0DEOz5OnWJL9ahfMbF9Te/PPtYxCdkqhXDNjqqQsMDClot23rx4EMReT9s
F0L2fr4N8K02LTvCqVklkOGJnXbueizvMxVOg5r53yrrbc2iJM/q/mbvjzJr
thUDqvhLpTFjJ1xrDibm3kfJvinL2yWSFZxpXbaCM7DcDYjqOZG7R3DsT1UU
OhzXi7QpxF/OXJK4PofRfyizeYaX7CTJZrCqHVTHpXaSNCA0GXsEXgUQSJv+
UG7xgw20IfE8NCNSYRbFSNgbFi1VRlz85ZWFV2PX6o0ecAOVzO65RFgOqYhN
2M6vuueYqT7j+kdmn+MdmAN6guEbItXWZgqBUMKdr33K5/fEX3Rw1PTcrvDI
jpmnzfjDitlxkuJjd1nsgb6O9aYBeWX1QlYCOtUvoBurF+indVOF1+T4wr7W
fu8zyLDUqJ5H0aNh+V2EkVV4j1B//+TKpbfy9XZIiQZlWBxhV1+sexM7szm9
PoBVoOA7Xs5Qj7buCOGRy1d61LYJJwuQHJf2FuxLjQU6QAh7HPsC0nW6e0yx
5FmSK7N7wv9op4lPalcafI+OeJfcJe8Twz/VhMJODLM3wEvEvd6wdp3c3Dce
bIoEREeahUN11kQOGchymZyvv2QtuqxSfUt8Ka8Ldh03t2UhwPZiXyuFq/wP
1Tsz155FSw32Q85H7khN5dvZ24Wj9HwGtwH6yAMX6cagqzmkWXMdAAcfhau7
bL3e8sT0MUShyapYot0dUB87hOdtib+Jt3mwxoT5IgMzQ3+ww96NJ6JgV37C
xIulaGR9X3LFrhnnRIm8HtKFJks1hE3LC096JNXgDpnTIgvmBt6wB/PnpMFw
556OrT+ZVOF/E3dFh5lCz4HKwq1WDgP3IAmRgpmVQEu0tgHjUmybhPKgtUbO
NRA5LpwjL4iuJ8qH/8g7R4ObbmDnUzoy94GU0oNbJxQbgEg4pTD4ohN7WuMV
dIM2aQ80y/IxQsTZQhksZmOQHkQJS0F7cKXSdKV3EU+ZaGQFOcOW1Gz7lfqF
e+KpXFaeKwFgTuXgc6IHpXh02tcBfHHvk5Q8M+qDyT3B1mYzpLXtBjmyQKMY
EWvL0I8E+ZB4DcCEQzHv9BueJ+kw3vvUtjXUoR69PWUEz5J9splwrNvKBKP3
2CprhQFNqTUJ3P4e9GZG0RsJHYE8vAhBf15YtrplwMn40gm1ezANSgju+f94
zEcubc0iRzlrVATGkZ5VGVQTU1TBdBSGPRbvlfGFKP2F01A6uoxg3oA8Vy4K
YhHd2e0ypQY05/UsdqXRQOEPklqbcjanJ9tqiFU6utELZ6iXO94f6sW3yXiz
ZwN/a0Tq8DPDaLZ+n/FYyWR8EzWh4ABRJODqIn2xAfT0MtH9nBTn3JrFjKvc
uRLPMNUaPbOmdy785X00tcNw/NJVnRrCmPZ/F/nei1RLEOYg0q+uWHyH3iZE
iq8ykbVILK39oCl00icWHO1NwqQ6vQVj8bu4E9yA+CoZGhU7JEEEWuch7ZFu
qJ+D+dvSjext/+uguZO2auH4T8fnq+BKGuMNxTelvdoQgxevzMLWLTYQA5du
t+ldQ97PHYMsLimyMZtJho+oIyRu6mNLwzckqfPTaoZCJ88EMJTyYtXbGEOJ
pWxnOX22uFIChilA+uVyw0ICCIWkr+96p/hSXUo6P0iWszTWNWgdjcbxZioa
kSKFG/Won5XJU63IdYGQcKYE+78jrk4tH7JfyQ2LRAohY3PH0cei5mB4GiXV
7bxllVBzChuRoR2PItYgc6G3yxf/KHZmD3inCBexP/8mR9xt/7ocnkAXIm9L
woxmL6IGvBFi3ZGrGWqffHu02YO2oMdqEwKGFFygBQsgA5mnBEnZT1GOFbW4
iNpkcv77PbOZeoOqLJMSUjB4poiNleHx23+ax4VNW5WW7ajabsUgIE0rFaEP
QdOiLdXfkDCig+sK6V4Z5+uPnEMXOZuxYcoNhixuCEXabzzdXDwoS8DluGDs
He2QV1J4Is55PI46DyYSXUilM0sxF97hBs/BDjT0THRii/FweoN9vlRQ3Uk1
fVWehzIKTFIZzQKA0pieUhjeYfgmJ/laBLNAQVryZ/w0b/DQldXncvl6KIdr
yHKqoloHrF1PtF1dJnj6sJgpi2eMka8fNlyuN0erk24IFgqXkYDYEUAuJlmT
cBhS0Yoz358CEZWTgZpedpFgZGAJ+Kw61oPhw1GD3/GScZ3v9pUEgNz0Ob/S
IRMZcJbw+MQ3u9NqlLx09Cr2OoFCKLujLfc5K62Mez5P0RFcBLXdQwQQiLT+
uEL66OxRVv0rcZ3VfZLucFnG+eC3O8LMRlnXVmBnk5hGtN25nDb9lpT06K08
ZyvZ5r3TSQ22U2tt1Y9ti+QEp1GdAOSSra6xD2bOAfsTfWxWlGew83NmyEP8
Eu0aBgsONLPYQ5A8lv5mlHmZtehZqeydFEQUZ+uINLoVHsGrh8zhvS30OaKn
ZNWBKOx1niJbh4JoylSC58M2fDNyVYOI2nxYMSGPgy2Kxc+/jwj4mzsVxuA8
95mhtP69RZLkEUBUQrXWAyVJT7kZRwQzD7JEgYCWeCvy7nE2/7ZoXcMJmamX
Pq43RdZe32b4dyxxvdfKkjQpRHIv81Dpfz2l+v31OjiJ/hI8TNWMtLuUK1UP
Ig+x17jnmODE4IZJNsz29/bAFePymKTyjkX7DC3kYQ9XEQh2GTN1jHMJu7xi
3wy3+ZHjfCUP0BmGzJ+ycQBkTRpoFy5Ncbrt/xVReVf6FQCd+XsOevc07xRa
L+e6DJp22SKbuMos/OXM/Xj6Euvr5D4CGu4AfRYe6nGatAw9gf5L4htOVTEp
4hTcMSWXFR20uLaFHisyL3LtpSif7WBW7GZ7FpypT4GQHqDFkS/JRoqDxxkj
aD5uCiSR68RW0ayxmmgaiGzb2MCWlEg/zK24A5RgidQ0Hj+QzB9J/ELYVL6G
R0VBY7Jn71JxJppCQJIXocZkX+1IRNXVWUMH50amxALCpeaThFjderUtB8wG
igBLr3QC19PtpXrcDBGbv5KTeBSb0Z80dYQxb4/72m/aT8Ipf+fbwwf2gQeU
nzy5hppYFiljMxvmq1fCt8ugYxvlL1OyCejiHijSK8C/wFATKippXp5CPAVC
jxj3GKNLu1ceUKqqEX1iCY7ByLhhZ+ox6Qr9kqdGN0iOfz2nNOiiuKURRsG8
HgjM0CSXZAQSFzp50M7n4cIHwRP/jz98Up20bKFrR+xZOvQbYr1+3JB1t6OH
W1NUCVfwN3EHNUaBRhqswwyUo5CBDD0u4LyfBOniM3DF3co2irZqWNRxf6sa
Tz4iH6SE/gb0jxPAD4yrSnPPpMvs5fBtnUUqCy+qpRjbo9tPTo3p1GMJJEuw
Ob0rC3DVfbqsQ5drpsuQZCxN6mR2wDc+6BWFrxV6cX/x2A363T3QkznwEoXy
BP6du19fHXuoxtZqb52BcdbCd7NOrH0Wm9vHaIayqlZ1kJvDYcKgLc5QQ+lT
0VJsc12dSXfItAQ53BmwDelGdXpD/MIIVqbozdoKYipjf7/leYbsVL2/sFWd
aTGUWFHmZJXz722YUBMYZgI25u5j/Au9rjOe/CgPJduJ1DciuosEd117vBR3
eLshzxWWHBYKKBLbufrBdUbgH9hZ25X1xdLmo0y/sPYD3S5TA4KfUnZEz+Lw
m2eMqQ+rDNIr8Tij/9K//U16ohKag9j7biGksiTwiru400VSKkZkVQKxxehC
HnMqqhRxlVqXEY79qC8VJ/8hqRc1zTHO3XOxZvVT3KG7I9hCiHqys7XG9UhQ
CDolO93wXUxpYE8dRbSL1/8uplzqPjqvzPjy9/yPm2boilmO4vBtc8KaMkvr
ScpN1/5qEtmq9WzG0Q8W1WzH05NoAvmFfIfdkzj7ui/z/a6yFN2TIdpTsbWu
CCuRnCp/3vvnMz0F5EMZk/VzIjPdxGWYLCPdytdA/k0x/Y0HgYhoVJh1Whkc
MkEvGL4omAvs2O5H8O5syMi+WIVQ9aVy2o84CzwmiQRYxhKpBV+4g/V/HwUS
+CPhGCjgYZIkgPxTB3Ep6xiVLVXrOpsCkM8PFPX+7yGJkZoK8Ckmdrzxzho6
+w4aBktvnKdUcbzE850gJlu3U1TKNFYOqSA2+ZfeeEIXJjvlD/ltSvfMgeCN
lsCs6XbU2IMOCp7Wu2OEW1hceB1soBgpz8X2PTigb1XksGOAcsyz7bcXOESM
tL1SeSdHRNkn+y0haIS6uUZdm7wrmApgZCq+fDXZCCTxFpXLF/uYSWbdl7KB
2oSSaacYrLs8a6xo2FB4j3q2CuuaxynuWHBTqwoWnZYIZmzhHxk1AwDIyR+N
9OCGRsGGm9LZJbJs5++asthaKjYrVdKaRzuKhbTcUi2+HqjKeoWMtpXQikUV
xhDQanQjTyLgHjbB9AU4O33mVUvzXSN7Q+zjn8C/3tE3TfmrMe08XPJ9U8Zq
2eqRskaa+WS74uxfeMmseIG1IQ7ocViR2kNjUmMd6sQjyyzo5duL0sS/hNXA
Rx8bO4nUPhrZLHsjt2c+5ALZFi7g9b2zXapimedqAPfaHP19FuYRsA+vKhlN
sfN1G6TTqhwGVEhe94BIH+QV7/MiuISuW2ZVy6YsYxfWPl1I5NrExEu96GHw
am+2Ao5g1folkdkchcvYIq7h7f1lqqNkaMRGTbrfBnhg2FhGtU2X/WVwR+12
oZTPMAA0EWBUwCupr3ouzsb5cntRiQr18H8CCMtdh5Ev4SfYyPhTWU8g6mmy
1uY0NrMppgEbOD2ut9L6bCizttO9afxHejpXBNM/nNHU/Yt/DfiAfUBjtg4K
oKONKWXw6r7/4DKTBVgE08kG5d1RjKYF357Ay/GT9rM2LEsITY5HXj0xt22o
T6neUr8WTSPXEQkFN0b2o5Y3Qvr/k8MyLA9cwr20GogCKjjCKS9f8QlbvQ+q
TB9gvLh0SzPsY50UjSpp/YmHB8R8pWb0a6IRDxpaugHpIUXmsAtTIMAnqw8N
HvtgORJVE9fck9NIJnjX2tn8ny36oBQD8Z4ER3/8Intd1Rwz4M9Vt8tFB0kD
ZyA3XjaAN7fuAMPRFwg0/5Hj7RwnPI/YboE4zW6Q7cISWOTiyCEVaCEk3xlW
7odng2BeS3o2g9+w8RCkh22CYF34qEqT8jbDj5lGfVpyZpAScRtL0DEIUHAT
TLS9cDrzg9jPMIrJAa+BHCly8b0kXggAEP6KF/bBa1HGsh667XKVLactTTm8
iKOCAH95ehuD2lYyI9meVsS3LuHGDOFYvltd91V0iUixUU4nP39nga0o0qMa
aZq4nFAfi8YdELWf1o9peI2kk2DsftIi+MIECcQU6ewJKlI7gNdD2VJRj2YV
a9TW8nZoLeivAmvQQ8RyGbirX9pA4j2HmdDVOBfeMC13/c2KtHW+9B0lTLTe
8WCfmVgbgg1Lx8f6e4vxeLSifWsjQk+Z1ExoKN0KKPnjKqE1kNPgCONq++Hh
041AAoENXj5P6fHeyD1Tgn7UxfIbzpy2PXU/F20yttnJCLalyT6ggR9pahQ4
LBlCIZFJymvQpwGSS9XIiZJ5Ook505MpNoBMsW3co4sC2bRaCu7i7wdqsEQB
91uYy7Qh8SWN6nIRyxF1lrbI6+kgrQKtnrXQQbHiw2hC+bioq0Q8ApjHw/Di
93rDxXwDqlYDi1Tw2Vkf/2RCFt02/6JIqMbxYl13Boya4RvoifrZTqBtb8UW
Pwhs8y59pCZSppTl6ANiIV1Xn4M5u23uvTZO7p91bDok1Gly99KFuc8VLYCO
AyRMyoSaeKJHMX0CTCiXzgwx35GCoKaEhd62X/mo8SkJgebdleR6dYsG1jXB
Tit5A5tL1fBipKuQ3WsUZ3u9wxQMlqX5FxcuWJXn8lejEajwcmPSQZGFWTGv
XO2wHr8vUfsZkERpeWKRbbdOqRhvuJyD/XfxsAVYj8JF7T/LldygE37KhjGu
O/5Zoc21XEdEK7OmuAuBlpmTJPRykYxNSPky4EgscQtOWWZ+Qz/ppbMHQ16b
lCqoaOmH+8p6PHiCZKj38DIrS4FnFL6VnsPcX+qKs7eiU5LVqRm293JrCZ+k
qkbUnd1ITdnqK+iyGdHKTswcTKrIfoTPmV+I5WNY1IucnnOmHSNMFVJ5oW7b
nqLUqp9eZAfT+8mJQGq/G0F5tXpDrJ83z0PDpWDRH9Alaa0rjQwQRbICGZwN
jlxE5HpzOvXQu00xERAzFkcuuqgPuHFy3U/PwmpJXu5CjvBP2w4Oa0Q+Tlxk
y1xYRIPqv9XsxlXD6bockrHM0aA1X/6Msv11vmEH5EOPgomGwbEUxcqHuiVn
baEtltmaO4kxBXPM4/LpVIkqAIFH4Ih5+/lWCgHEFrCspGWbtWWvJGmfavxf
K5Q3sa2vsxnfjGFxERO02U0azdqvS5QWgChfOs+dCpGGBggdRfzJHoE7OBYD
udVsNXBmeLlKL0oxW7vBUw5kkJjVIjoQmKvFoD4ScH9D4ZyD9zoEXVIzE9s4
4F2/wzXBpoJCvW9rX5gIUvqe2uvUiwj7YvOtDZOAgTn6IEFXNu3MK0OD1vUh
1ol8oBviFc+ogVE8+rBvMiv/bH7MZr7TywSzMPl35sWkjNgxVDpIcaroq2Cu
8rnoL+MFvzF31szwq2D+Hw9dSXgDDpQlBgi2YdFsK2lKV/gxNdZCvm67LY+j
ggnR/5BDo1k6sHVYuJjvaweyeOuQOi7EThKI9B8aq3VJduaWClTahPIidSLa
xS7L3cfb6O7u7CAOGe+YH2ZEdxWYDQnGRBkLvK59FUyvAtaZiVPmpIiN3M2b
DBT6EH/zBKQQCWoazen0aVN2TRZ9Qis+yd8zNnwas28Hd1cl7L+98S2q8ctp
unHbO5M6mI0gGZptCbiSRDUUDdVUkc2WUyR4HXmO7N/YzOX7DrN3sA9H1GzS
Go8+c4f6m2VCepncCK8RTanXJYdBhlQYnmyPhfuT5YF6L/vAQR0xE3o2MeTk
0Q7w5IwCXFBGvKfn5/PQcxixN25ZNNfK7Sl2ZRb7bKAOCF+cSpZ/qcOZPWp5
rPnOdHKHvKI+v16akL6pHurhqL8I54fq11cqqER9Kzw1LeH8e4zXJJ8W6Er0
krx4KeKVGBJXfugp1vdpgmqNVm73eqvzaLUtLO6Hc+1DIBXb2UvBnpnwawj/
AR6LMj/3m93oawqs37migVVGgAbhHsN1Hmlisj/K3ELWfri1X37gcomWg1vi
8OhxxO2Ht0zz8vuW0e9yCliye0OoaCzc0pxldW4UvZtegsZ18FQNc6gvLczn
hQWwxptwUsLIsfI6tW0kH1s4taJqBZoH4IMpQyqx+387YM+qK7hC5UJTzIJ/
tkQ0RXpw+k6bCwRQLLZ8SwSEB7NFU/5zmOBe/WHQaKrcMcNwUCq5UROPZyAn
imc3E2HVFrN5TzqGUfFBekEkbR6v/uRZHNetl7x9Zpq5vgaoPXqnEA/328uh
XCl54qTdJQf0JfINF3siEEhx048TFzwYZDkoHX6sNIKULxufM1JqEf7p1vUJ
NsWU5zbSg3nAIPndvjM7Zgx/QlTCRKvdocIjK67kgJgmGBhiwvViRIEof1fg
fJKTNNigcYbNQ19wu+01/uab3GaLj93mO72+/4faT8PcN5CleGbvVh8Rcd3U
FOUfwEYJQrd0hNYk3JkffE6UOSCYgq8enftbVrC89OWvx6hSGSTKRGRbqwLb
4RWDX/zHEkG3mxSpYZQQZJq957lhj65vc1ekmJrIWF8lo+cApA/QtW1MI0Ys
IFFng9+05JZRd/ialQ0gxYs+817oM+t2JuMB1d8tD+veeW7huXSNtLNjART7
qZWH3UlTUd8iBzezHEyVACbHmR3jO20fuvINjuk8hLL5a88CB9+DrpzlI6Zz
J6m3XOr4s5EYSCZWi/efBDVUHWLyHc+xdbNylfmSbevbbIlRulN1m2v/wjrH
vLF+qJuHZrXJ64H5+/RZIq4wlxXkffsFatP+MShWZkn7AxNCOEYnerhYetJf
95oHLK2llf/7oCjTZxBu+FQpq0iVNtGJhs7YVw2LnVuCZ1CUdHUIBrPCptzI
bP2nSezzwzkcqtS8WqC+dx80sngnDZTLEqiJoAuWAqyIQFqKqQYHKF+HCUzz
JjTr7ZUPcxjhcpvA52AsDxBjXEppRH9MlWJPtpvmxJnli+qlwY81DUxFAMN1
0ek4RLCW9r+qsF+bR6n54ulXx1i2rkgSJ8q1zhy1OqmsTC2HS9thm4i8ma1F
ifDi+R9EukC/lWb2qmPZF6srY1Q9rRgeOwWyuYkTh5PxauaWplKEPyutUkoF
NsRW59UBGQ9BZyY4TbS0VSomjPGM0jKwn9SZYh3VHni5D6SyWOSA7sIDqYW5
cswfvGhXj+4pn8pmg2cnzD9ic6RLsWO0SnwayohMZj61NR6V7PqERvaGclxh
vT4+y57ipY8lCKE+QiRje71jtPeGvYG1qW2StWbU++U7N+531Cp2+BwoFx8n
PjSHixMVr67RVidpoOtIsi8KGs8hs48XPNScCvMEWnQq4uRoqe1mRsrDKRIa
fBiVfvmQD+OYCzBWLsWtJR5uK3O0bf2cyy872PbFTKNQjkPIcSNcHkp5LSCt
wVXRqAzeewNpwWFpKLUhqUXkW8pMnx1MWbnY+rf2cFcMVAIjGcvqWOypH4vM
b9oINP2zAyJ9eAS/oKHyUr9Tf6i3Vxm401EEISWxfstKdQsNhqr6Vm8k3gmp
lNORbb048GNpu3cTr1RDtpueCfmm8k6OIUwtFZT8iDt3WlEWD8o4Mr5a1hg4
tDpRroSax+UZST6kZKDYeIwLpGlnVZpe0fi1RUh1vwSOiGmuYjaLA/bUHb7+
8sG/+MGlVBUhrE8IA8aj/abEgKKZlpLlYSfkpR8lWYVbl8BIiaHZx1rWZd9h
M7XP1J+hTU3xSXsfieA3VM5zs5HuswaglDMsEhufZeqDWFkR+yWjIxlJBwUs
/UIOiqSonNZ31BdXFU3tfe3P1mzShrF1eFJ+7xD7AebRTe2dcUVfrOL8Ah90
YRXoiR4g1L+9YltQf41n4Ea6HazttlxeItrD7CAbfxRZ+ASK/c4P2+ovFsIe
dMARbSV+O1dakCxnqMqTiwCZOVaRxccs3y3RNUjkzK1+ICE+tM91P43Uje9u
6+lSkUcblIEJi2PJ+VsliY3JJiZMCIQ6MfqrE4GF5mrNYyTFDgDeMK1FG5DE
6tZpI/i/DGsc28i7gzYc4L8/aCTdVl/EhGunKm2WjgzlyOt5x2R1XtcukHfj
CDxQEI+YYcCbxSRgtjq4kCjh9zTAOtNqIcBtY2ad1rAVIyoIcu0qd6sFP2Ia
R/j4pbtzsP2F1qaFHjsRDpm5zEgAKa7vrSOU8M3T/ElUg1H57qvvOMk+4vH9
acpEyTfkmkMKGK/br+d3/Kperwuh8zdBsnpwegxDRaM6QI8+L4aowyAD6nu1
+kNrU12mPjYAwSqDlcb5DYov14k/vNMNq4Giatb39LWeNbtVp2zUPk7JtbAL
G71h6d21+3+wa3zLn2WEm/tt+cXE6sUAeNJXTjV2cou9oZQgvRql+IW1E4XB
DzVuYOmBVSP/2DxW0ybSG7Zv32hj6NsAvo8uqaONClgtwdfvaCiD3BYxsi1w
MO7lYKxoHOxSdbYtI0F1kTI8cm+AWdTXwMOK3Pj8ghMlpYlZeiCE8WTupAuk
lVVDzmrDfr/lIEWrfLskzY1Ao6gSJUuxVDUzuDZ+ORUY2eAEl3eGzE4dHgkH
4ey84F1pWq4vMa2VCqNv3UgTd1/qqSRQVmXO7Vd2OgDbC5NX20zSaiKdR7Hq
lXoPI30Yexouz/iSYTX5MtgqYK8RSr16/dJCaPz77Irn219oz7l1iPTBt9iz
P/zv08unaOXRULfKdnLd3MbSm2kJO9K30MehrIsp1ladZPX3fOYUNL8g8J0z
dwcOBjJirXvfihB3JzujeFjb7Y4f/BQuzrO+KwDWUof8B2DJM8dL6vatdonP
1wfpVImJ11YIPxRVY+MGSo85g1JNVNOm71bjscJ+LslWjt1uSsHP1NZ319Y1
tgbIA83nly+J+Nw1eCgaUj70W8p9VbMQB394FAs3qCSGwjbHyAA6qmv1IuNQ
dbFT5vw6NvuOfUgQvSGzR9CYBfcPhxiOpWl23uJeNpU7wiVB8pzyDpOkP5ZG
m9DFz+1aJQaeAKgf8C3fA0u8Mo9B4+rBmezq+0zMjzLytLMq9IceG/A8GJPU
2VXuRQSLl6m5ao2RVYbi1mmx+/SYSUFyaga0FACd5BCJG8Rgsl7AOz/Awpre
FdGMKLUGoH/ehOOVTaSJBkVSC8zcsWFTqiJqLlLKahhm8008kWyah2NURqvq
AafcSbPIVF7KFtu7FwvIz9/JodNCEWrya66NzUqMzOcYSuEb01FoLbWMpe+A
oa34319/mjLFM7ME0VPXABdXk36suUyX79qdE7J6comB/iiEvu3arleA38Jn
2o3eDMMraaaNKeZ3oqFkZuTv/epTYhBaPFjlbC5p0wKFXaOjjolUZUdfw494
TQvUgfujFCwVlgZ0IB8pHtqnXstQvQ34UXli+Zwib+RjplyW/0Qn2vVdF8FH
gs/HBfQRAFNQGzEG5dQMYxJIuR6JI9JO7n0GZyl1gYV3Lfj28+eUXS1Anyl1
9KNK1QY0tbirtn0HUx7PCOKBxZXNDUK6GJeDWEukpOiBofOOSlMNGgmtihKO
DxWdVOOSdap0J2LtCfWC5J50LcMNL+hTTs2W6tJAMRFs7vnlCKEtjY+jBTIW
PqTs/aDPYj1DzxKi5C9Lz/LPzXIs2GsrYnvRZxNkzKczjAPvKXs1ztgRUYKi
QQH1xHS5W4HQz+Dm7Yhsp3WRNODzWxlfXNRbmgutzYg2O3GY2oyXxkNnUurh
W2FKDZrPXeTGNXx/7B7bTY41vDxgp4ndFQrrpCNUjYJ507oRUDyDKiltFb2m
+0YPFzx5vHLY9gGcXXtQ1+6YVnoNIgRHnkhh91m2Nu4FEymtesGEgklaCEDM
cZMQP2SuKSbi253TX/wbEPhRsK9gNSkCloRKfWjYxDNrQP11tZNsCafvNetk
gZMFGdBSjVAdpZuZCS1mq/+xaOtTabgWsHPhbMqM8gZjnhKfZYuW/7QaWtQV
3norz44aPm1xPUWFLYWkYNBdiXOYyVnvNsO0RcrdP3w39AiJqXl8sn3RUmjO
PmQdQ38U/kTd9mTqOl+Q3CLhZ/VWO2Xgn8MW/kqIDT7X+jkurPZ3GjoGF2MT
BhquUDLoZ7nbHsre/n4DvBcoZ3fGMxOVRqTTnykYrljvIVe8+CXIjGUY/6fq
l1379I4ZDVXg1nNpZfoEgzGrXr/XPL2N5w4cQKq8jp0QG8oqovO1j/WIHX7q
jEdCjM6hOQ+xQkvXTmQXgy0bTPzlJvDDCzfpR4rKGglN6ucMOV+1kkbf/vs2
FPSDIXzCVpnSLMps18A/xvfes9aMpP9VkddbxzOL8oV12hcgzDl5IPwPmGre
jNsH5KN2zDZeKADRUulncmZdoCFsNUDYi3HdlPN+6f5PgSFMrVZohit+1MhR
lwrqp3RyxxToBQtomc7offcuQtZXd34AR5hdxQbJyqxUKh3XDR2yKFMnAVlP
+AYNGVFHVxnb+gWpcTbjho+u2ekbkM7hPHf4XFfF4iw5gpJzC+aoXu2m+w85
3Yz2SDD9ZUHn8nelJr6IRuHMgYvnsv8PHFBWR+u1YiVclb8MhDnpqvSxIvPV
6W1socaGWGw+/sLBrP8LipJeK9eVXcIeF0wXtUKGAPV3NskvKa24FsAuGnyw
AX4AymFRD2hz+kPfQfJoLUV2qLlt5FztuqAdGpH9A3BuSep716SP0Iqqns5I
tweJRnyXBKRBaWuhdWaiAX5RNvalg2aL0xzZRWCE/AAxgCj6RctsDvgg9seP
Cw2YCXXpiZEh2hn9IOLKvKK3BPW1D6fNPRf17OtG9EXCrGRv2y1tJ/Xk3tr9
knq+lkkzBr1INJ9HKmSTlWSrBcKBFJxgP56RumNDuXtu9Tk3WkTj6i0o3zHm
Z8YxYAPmPSM1AjTcYmMnUTpSKSdUiclApmPHnRD+ZBMFP6mukzygsVu/tYPo
UMKPIuG9m229JCWmkAoi/vtd19/OoxTmBBHXd5fxNBr2SFdK86WDpPtSqtPl
HSHGwyS2yTh0Q3v4fyxRkUfjNPXrmUCDS0R3f/PmopTIiAip9SXW1dFM61gl
t/00egKb6NqChGbU9chX2PVhoQ7lp+NX7ZqHcuaLuITVkigSiS9cTETS+Cns
KYmPHpEnYSbdfH5Pq2V+8Ltraz/9C55qw6YVQKERdDqQ+ZmdKKr6m0MxEX2f
V4Lt65mJ+yUz1lAhwIUuCM9DnvQ8zt1wiRnfW0xzQ0JRSFqDhXLRgISAtW+b
/bFqvxIHcooXHG5JcvZnKWwsHv/ml2wJBxNeE+oM++ti3LECLvFp+2cQwA22
S2mCjfkPCtaJLUwRXnszvPw+/o+J/ZSjqdo73ORXH2FdNBha8sSN6yHxQTPn
w4XHOTC53xCd0JIyk1H9fXzx2+ZIfqfQnAde+rPJW5cDlhFwNkMFXPiM2VCd
uCF1T9qHpi46cJor+FIzO8cIwxpovTznslOF8oIGQ5ISCUMDwFCruV5z0CLH
FMcjb3mwxxUrPdDSYeRz+VPJBXgyhXhWnF14nt/Tw6U5glspS7St/zenYPtJ
yWIS0RBG+bOXIgNH2M/o/4phizTck9MPRvwmqCFXqJHbPGJYcC3XSPRk8iOA
aqMkZcUdZF7LM5EFhS6IYdldnRfYSOlZPGy1rzAomrnEmpFUGGLsytmUJjwY
hH7KQL4AScisqwK/g6MOWQ29ExG5ObSWA9Msmzz2mIHZcxns5fIpxTjZwIA4
CG2q16mzcU6+S9GdChe4HxLwFvM8x+ndZRn9o8ipY51KtN3izNUB5G6MLvXO
2qSPURRzj0CB2s7/uQqic09mY1WnSTXJ8raqmDMqHN5xfPhhRGeP2SWSJy9N
8WqPE3ESO+pKetkKTMtUSCRzt1xKDvxkA3vQBt9H9+qwo48/auefMXEpmyDo
3JNVebb1nP9cYa9uoBE1QeHqxxLR9m193YgAPJHPEzUhwmbQp/SesOQYpZCk
6QFcgwalUqp17ZvQYAvwKn46HxAEuIHsBVLtYtREyhaFdkEbTkyrwuFD/zSs
o07FSdU9FhU0Z/C9F/TNgDqNHG4Pg7v1RQFQbnI1okczjFbLawehm6vco4D6
edB1xqoIcmeSjzrWIGGAUwJYtgV9BjW5mAeNCBqzZC7rdBUxV4Bsur6VgNr1
ddfQNek7I4bSMjszy1HVKUmqEEX+oaCC/Gl5TTzuHncSjnwPW3rJYvOCh5MK
plkM0xvskoi7aW20KV+u9Qv3Mpqch0resvjmDU3xlTOUSHmAw/P/vDOYiZjE
TQjI8llSZGIbHP9Nrx8iHEPJk8cG/ZM2pGq6L3pqjrfflRm9/ZO6tcxahT3s
bAeDf7BYnk4LOrRgH+C7G7c+nLeDAkIK3/F3i/SJaZUP86m7XFbMcZqox4+h
ioD7rFX8H7wuamaOD+SS2erxbuOZFKkwW8tnrlV5aHKRo8qeGm2cKYp6lrU2
qHrBSfY01lNVEwUOALQ+tx11sMNeL8kAhaB1CFZrIBLNnwnNUYhlwMDkmjle
LM+Y19Qhz14i1IzHBHktNU95bsM/obYe4NGL6hmwA76DagSYeyW9QMjrRfWY
iNVYWzqLvLvNRYRMq/sej04nxIEnyZvr0rnWB2nxXHVbQm70g4Xv3ky/fhD4
y3FwGnR993BjCkvTHSez2Pc9q2JYvmFDOe+iqbiU1grCTnKCNQLktSx5rxQb
+xL5HW2IzAEErRPVdhkPxvkFVoPkyAxf291r3+ybOK3G5XsrfzRuqNHbgAMV
8tbmv8JJPLFLqwHFWOtzfk/NtgW0XLU2QFlRVZ4pRbF4pw/C8Ml4I/alueDp
H3WFpTDrj2zo9UMD8o5ntwjjomzgah6RmBs2Aba70kJFNz7SCki8FQtEnD0l
HY9m1sLVq7H+aNw2v/CvuG54fLtmAPcDl5xS3gkN5UzLWPvItNs2E9xqrPCE
/HQWW7hwAXPKEL7wFaPb0FzR0Gumdeaea/zGDTjNTgL3YCWOMr238kWCR2Fr
Z5i8KXjUWetetIfMHsI8nobh5OkLGfbx4aW6rY9esH8AD89P79F6xyV4x2Bp
BTJp9/qJBgpVSWdL4OjJ7R/WDVTJqIs5Hnvq9wreJfimkohFflyjEOC79CNr
lxWH2BSIx+qx1urTstNKTZZ80VLtquXDMw+T/86bX/SR+7bQqv43NxSEb6Z0
JKGrRjbP3G0S3wvJzkNwon+rdxNmwLgc9AqgEzmsDkteifzc2xAVszezUIGo
8VWbnqFL/MKpnMEMyxq0SwT1M9/moafxOanTvhV6WRXKdqxMcLzZoE7Li7Hu
YFzhGKZ4gcEd7vrJqAY5WdsaW3U4N+tawG9IdYxLX8cqLNFN9KljLAfzLhef
vMy9vtI+5RHocE3piC7eSE3uSLxOlmkNMN46EFBba9oEi10ZICYy0s8ARCZl
wla2KzIq6OC2L5TbP5brBU8eLqdgPo/SfmGh7C4ahyS8DotURtnCF6Q5vQeX
8znt/ITj8MLPm8ecvX4SnAdAm8YbsEDrR1mNLtQsqHWPZdhWixWwin9Q7JjU
JWcYiB22ZBUAYyQAqNVsHBaVEJMemw+UAsQ+hkg5PGSJl0e9GSfvlfHjV5wp
6sSWdQl0wEg/+LEw1zbgEfxq8RHAzIuXRrGQP8SwlrkB4GzOrB40gsuL5d7+
mKvW4RJhx5nRxcmzjItp+q1e0FxnDIZLrccJyR7Ie6KdIzWvUc02YvdFv0vK
E6ibAUgV6ofLa8R7by+FMZY41g3rqEut9AE+/DUwna0br8ES11et6wMqchXY
w72ByEOgmGABLF/TJ5FKDHn4SyuWfiuVPx1Q67QoGmSgLhwv5En0gN2E3+eH
OAgo4WS4BPXItT3Fo8H9s01zDYz6cXh515Cf9JIPvyW0fUb9CHS9fBY2hdmC
oHH1ENZTBwBO1ziYu2XjGgcDwAu7a0yPure8ke88asA9zS8Iu1hFoqIanC2+
ORbrUvbJTkiPcsZmJxRIgeupGNV06cVOE/Zx/i3xZIcbI6e98QwemR20KvHF
7zYcCzqwEYFnyslBOVM30KehnmSBhVyHivoF8Y6+SFo4SN9hKbePArhiYuuf
KzCepem28YavTZkHr1c7HmdsU93BdZDK8MqnabIAvBUZzJYTHftbrfc95R+E
uHgdiaBHjVmpNkG5DrZCFg6etBa4vB/PCg8uGaoBYDmHcObE3U/R947Fq3qU
RvuXd76jd6PZGyxaqfvu1DG5pCsmkwf7P39oHfR2j2KCki2R260W/P75nkIG
kGDfYizOSqocAAxUupvuwXc2ac23uSBk4dwflNrcBoOqltpL9PJnntxu2W5n
oUKkJlufXEWBj1RGF2Zs4SzR/d7+WncoXoR26iWY3nMchqz0gwSjiUskbCGg
q7/obfR/ZbwmRVGthl2l/Bw4U+ZyJyCAuRVS2HTcZuuUVaUx2C7tRi+yl62E
oXlDWkbPnVj5Jg1AZ9Eo9amXGCSg7nvG/lq7M+Swj8tNz96ASjucooyGSku1
3pXdGj/zJaHh0c8JWQHh3dYjuKtUBgf1yrp7zQn5+2WlIHa8SIjA+wYFtHQ5
ORGid8YWxZSr1iTAT7KTJXRBpbkuMTc9lWbzc6t1GUNW/0muDCODvPWNcWy/
o3Oy2zT/KJGWY/Lg+T7BIoMhts5fhLV5CM1GP7nAT6sNdjg8ukIUkHsR3aCq
Fqgtx4nUvts82Bvr1PSxPtELnOUEh1/TCExOlZMkTS+qFQf6jeTtnLhD37IK
sVT6RU40ABgnUSnndiAJig2SZ2YmSQy+D6syoIEtR4PhLdHXK3Su8SQ/WhGd
wfUfaggHFYgYXfskX0b5NLa8c3xceqYvV1GOtsnG7WrgeF/c4+nAMW5nsV17
9JmdpygnmjKrHQeeHdxzigOCEiNOvfaPEWcMoMOXl7fH7tXhSCWBUSR1defF
v5EDNYnNk8bCrbizIm1CNUtnwFv/Vjz7uTyC64SUV1DKT+UGewesiaBGZg9w
75FuFgufWVF8Nhvf8upM8whnN/ncDqxy4+3+0X1WLQuX0j4qU7LZBC5fDdo0
Xk8Aj6X4Ph5+q52AoTe4LmgSg8pIXHJ2DKeRRLQaE3yLLai1wIP2liYavqpr
kISmoK02g+xFih+EHjUc6VrAnMcDgo+Vz0n91TEJjgx4fla9Fpjc4ajyyfc/
cV3QdpbynEGCH777c8DDWiEnCKh5pG+ZVt+EeTJL2NyDEQSECx9XiyEWV0ov
T1pfr1bbPX4FtS4o70kWpqSJu6DXWY8tWYB2PcpItJQeEuodmjxZS3B5kN7A
t0NpznvwFInTqO4iyZcEd+YD0NlOUxiTDXtTPEiB0gws21U5OHuWtJE0F/EH
bT/F3x60IiBsxIuUk0+rKYBaS/mEdN6sJ4Te3enqkNEufORQHV2NFzCyrJ9x
eveOdPPhTawgHObyo4GVZR6QtkAv6xysboJ5ncs8yWvALeRldpNPnFXPpnd5
rH3MN0QwtTLJ5CwsTiQ/m2MKin5S7OIe/tqNCZB/qy1/DXflVUyOhcb+W2Dm
lDQfJPmDJW2ZwX48sWq96fFQufoNvqfjeWaXktB12ltfC0kQacRi26dyK4QW
FQAr8JAV3/ZvO7NjueTsM5kzzz6cWXPdZURa5YexK+vLSVSNyyVgzkZ/bTCk
prxoQeVwOg4uf7JvchbF/ui8R+48EvE6aV6zVynuZQaiOzdZvwWt0dpboePe
G+W37GpL7IFhgiTuzHqL/QqGoTOI4te3KgazTi3pmddBwQryaMu1/4jbIUqw
6wcm/PDwphHZJ0MQ09gWwE9sqUFhiAcqdESuAwG++etiG1shT/rzXL4iNR3k
YHw+McuGllJMWgh/55tnYPBT0D/ur7GwXdsXiSMXJjWxZV9mwDeT9cfXfyfO
5QbZj3jKTlBa2bJdrEScLX7730nyfmZFMpzAhONyfbM6GdufYnQeOH4MAU3k
X6PO9zTaVAk6ZvA+JAZdgEXOd0KMCfJ48oMqnICjolf0gwA7x9jfLvt124kq
ErRG3XCjR2PsSti9rn48CGG66TKExBljdqU1wxgNIaLFjXWN2sA4TWJ0C9b8
wpd9dVdUdSoAht70bsTZZgj8GFHiSLr71lnHptA8fEmMDHqCd2lzUaYL5FMb
I97/7gdTEYYKe2amCEeTtwHDK2LF+kf7DsiIm/ZW+xPTFwkFSfiuOmNyh9GJ
WBKcOqYL/Az+uSrR/ofQAi9Z2IPjwkvmro26uvV2f5GQVUUUZOP8r9OPAFZx
ZbMefd3pF0d68qVkyLou9WlZDTu3tkddlOi5Kky65KweXVv1qLD8Hs0LjwFG
2dFqX6K4FRFbjxTa2YTYXI35hXMT1L33Ngrwpyz6NW1Jm4jXgR/Hq6TNdnu2
kAlaHOq+Hw63/e0Yvemi6pavrL9N5XBjjgDcwa4oOYmFQzmUtey8tGb0/j7F
FZpp96ajMpU7eu02L59SY26iLmzyID9CzvsoPYbjU+wt2Kclf4aggsc1OT0u
GscA2bV6qSu5DFObvV1tvWqnhZibEsLxA2ALxGICDQfE/XEN4kJg9prx8KHj
vdOTeHgwmDxhdtFzDNhdFrZtni/jHelyHtXzGot9/a4eQHxPTlBb1rbowW7r
No38nAOrhT5Ebq10vYd2F3PcY5NKUlPMy8gUlc/cd2esNx97RYe4rnlmfu0A
SDj4GlKoQK2O+x2vVzZ3KGRanmL7o2rUunSncgmBggZfautGZEVXTOaNjURB
5mYg8qrkxw8Z6ZsYAc1IsP8896mQ99pwFSsP7xf5ZHmJigZrKsdJU7UkvtCA
KlCPiW7pJ5YA7TV97QMGOA9NO6nDR6gWD6o+Ke8Qj61MiTnoNqsqKU8LOfkh
G/iDib5kVxLWjqHU0CjtY8GgPyAmBRKzaFfPFMYYM7fAY48fh30VwI8+EgYs
LkekEMqQAUaynJ0okEEtVX8g7UtyElicJLbVxKLQofpDxGRycceZjWTfvyWk
+VJUARE9xqPSlk/rU9dSquvR6/I9jzchZmx6msSciKXjw6xYYTn1r7ngFWPL
i4s5itgoz6YyMw/nfw0A86/FiI4i3AO8pXfpXT8JyhHjHKMNsOLgBk6q85NA
fFgd9TokM+m/Cl3R3YrEuSiyDVNCIT7wS0T8kaAPsb178DlSECayqgdd/YCp
Opu2TuKvIYvO/k5/KoNtoJyaH2UVVriSQyZohTqeONaev/JS1Yi7sPLa5uAx
ghNStTTpOWPRzB52OQQvVmVQH1QVA0kgNMRnF8u31g05lNpgOEplbI8Bs6HJ
DEhujTJz31myYfy6sqQmYV4szwRzygh4YWY5SMcPkQyHPMhme94iW7OgUo3C
utMDm5HKgXdVUWXiaMURwvDpEPOjpLM0Hpx/MV235DwlbDssZRqbO25kMUR2
idectf74cyhNMc3OxQosmqudIGlNaJ+hjzJ92bM0xIc6juNP5PqVvJNwxmZ4
2RVu57Y4kLgYlbQDDqfdK5IRmtsD1p5d0uypH0lLpDPHZsuxbrYEszVKLFuX
aLPrmJgLS5BKFYnLyjHA4/2iKKgjbf0Jj22MJa2dqAIidB4kSd5rXGRDB1bg
JRpSL2Wy4X+UiRNBzGHRn6/MhzJ6HThnSPh7jQQxBFYOEOjEa8KJWgSd6ShN
ZgqY6qZstHYat6ZATDm7+BpByDSapotDcfSe9RqyYRA3Pr/NaxvZcr2emhdk
8DH9T9+XLVMu/b42eNbd+ZtqMzfewtX3HAtB/dwvPvHXCZ93S88IARMPXFEE
DCn2RQj1O77gSVmz1P5c52MT3pOB80OTEWkl+xXizVo3t1+rG4Ta1LkxVyam
P5dFqNSWhV+b1yiSKhee+ByUSzbPH5zxJMJCAGiDB2grqOWzClsbU7aDzMJ9
fNyI4kiKO2j38foKZ2ziwV7pGFPoFVJotCA269TBc2hOJIbhjP9bdrcwu031
FlTntn4q0LxnNLsOEZy9gYTuM1RB8ZWHui0M62YaT3CgE9CHeXMVa/mLQ1OK
TqplJtU4uLu+J7egMX29BoSVyQuDngP7hC5TEmTIYrYt8VB8edVC4fGbskbp
MKOmwRdsI8PGq8aGC4O4HhOIIBJC9LIUN7x1WVT7Xg5Fr8PmLuN3LDxK7myY
vdJHwnZ2J4KBKIb4+ScsDp8vpUm6k7FL6O0SO3Sv4qiTppxbQuCpa2N8AUs0
W8INN+mUm01lNR2cXh3FM3iPHOvEuldhMjIQgm6So3aLNjzj5MWhd2LcMH8a
JBuNIwX3Z4Vm2d83LAOGpcmiBtppBEEOabADcEDK+jv6k8p8UdN5WZKJyemq
1G9j8Dk8gTPwR4q5tTmUsToKIIbG28IfzhJkOHarqnKc+MotldXWDgTvx9nb
9AhwEs5w1ZEIUKKexDlDdqhMWjMJXoaLY9+OybExpBVsdohBtRQSMYWITi5l
1d8povvjvf7Th///qiyuo1hnTtDCzYN1h/gkyi9ArPuJWVDcT5tA0QD+7YGN
kyiCKiLSLkiJcnI5GdUs34hAw9wI7iuYtq2237MS4aaJc27GuZujQ+rWA65+
ghSNrCt9BGLwbxtZl27Y2Sidb0IjRkJjhkmuIPM2iQgEb4Ap25timz3hRGfu
YHb5NfvW++qz2Ty7mpqG6wbbSeWxM0G6JDDIKUhdEDncsO3zY3YDYztJKF6D
2iYGFJvHXPHxHmdPD9SNSyvlTr5LLuFdlPptU4b3+df/T0GWl2JDB+E8JyXx
IOflK72ds14pq+cAKEkucsx69z7ItVNB90eks9ior8AMQkr/jA5cpAWMLbFs
4SN71zpIy8tQTseeBXyvaCYahY1Og3hm5dR8OWov07ykuC+wvNkzaKPHTGJ2
ZNGerNik8h8oVnl1xtjIQrnK9td7lfwcfyD9wHXqGKJF3ex2DLBM9AMLm0nm
UgLvRB/gdDuM63D4kXsShQRZrOdUR6tl+FE/UboZvNVJYFMrBkS/SOzUKspr
0ERyuKUWyh1DNZYQXAU3ojCG5zG1+lDRT7AyJQZFJ68K+IDkPzhTIOT1PyLT
48w+dsdDo5fUSMJS4ayNTM1ogEQ1sso9hPz1O97cKlHx1ydTpDJ6tYBwpXw0
fBEeDEkyPhQ5JzboCylwAvTMZkKhIsVBt+uPsQXT8QSlrHeX5+qrFZP1Gnsn
0jhQ+VVGBeoCpMCWWXXDmogsMsslosGvZv7yscaenuyLTDdzUU8mDtbo3jdV
TqVsRGZ9iKo67Bi16CfH4DMnG1AhhbN1xoh6/LsVT7kHlX07qgXB9BszptgW
SZtc1+XAzxKhZTxgZnc3Sn2bL9uFEnY7l58MjXNtWLrH+mqMNH/LyCWf6JKz
pl5nykmr3JueuEFz9WLE+eSlWSwYA6MN43HPrKat10nHoTVGAYpHN2tDAKH5
Sti6sNTa8a38ItZvx6jUcorX7OHp+OxCAyE14pREMrkHTU+x5ZCKZ39q8Wub
YQj/qqA4hTzMup33jNcYc4Ll1Cm0Em5b/afZQ9InxhOF3Ifxwe6HkpsTIZjx
hvKIMSBwCcM/nFSRAth0VAUM8V/bm+JrimjXNdxzcWosaPSIQzWdjyJddDuF
s9xiBmbpxN6NHIH4TaWpNT5HdGhNVqzd8PQsqDVyNEfHh1P9fM6LFJfsRMB7
IMTQFOZzD6EiuOEkfxuFGSYi8Fl73YAQecPxMuEkhZDkd+yY/hod/AB+P/BO
7usjByhvC+EiIAFFDrQiOD4bK0LL2c/gCDEM/iQK7TipiIIDLTdkFln9N/d7
W+nF8QZKc/3WuNPxBiKkcHm1WzE5rsuEWwckQAXst/2P/bHZOKXeoaWmRPas
InTlBYDj5n2oobUoL4c4xp/+mFJV/LQfVLgP4x3yUitjpT5Y8RQbZWS2J1GD
VvyAg/7QAPoS4tvj1wTukLhBhSFFFxAT6LVSLTqvWQZMJP57iRjj1eCgmZaB
x6Tp8mLsPLkckqqsTw8IW5fOXWUUMmnzsLEHnWCx02Ij7RJv0ZVjiP4sEXxE
ZlfS/se1KOAScF137ZghRYM2X3T9+FjLXHyvLkwuEUzD0fOD+rcFfTk47bFH
KYkxowUsVH/jmzHer7FgzjCL0pCkA5PrsvEWsjbyzfCUCVd0fItuADQ2BIn3
ncnWL6JcxhqorZjmLXVZIS+FarC1wG8eQdiGfiWDVOEZaQJxfr6ozvdrYsqv
t/d3v+fLYj/ktcDUk+ptgkALsu0M73zIykkGcNHNXHUT6dNcW3KY9AkOVYwy
eKtxbCYtPlAg7/9JJUD3V4Yjzw+BkSKmIhi9BYoIrAzZkf30+xbTOAvzBZkI
XraG1pvi9T+yWf127jOAdT2r1tzMuxvmJxS0Q0U5tt2dnnHxTIr7jvhvr9t+
Ii8HNAA5Yj6MgEghEthTsVYFdBxrQcLETAcs18DsNMoRQrabyBydrtM5W/v0
4VSEz7n/jHVftxnNgzYoICEpBYZmzbBaEf6AO5UbiHyyov9njBQJP4/NjVDw
uKmNOZFI34Ao1AgBOP88d5YrWf6hGpRMbdoNGDzjQNJSAi9iRF8qerZSywSC
O0r6IDDFrIfdt0hEdq6j/lfhXSHpCQuhB3GUmZXDNkVbtaUxUYSxIEgTQz8s
UGmsqbHjK9iZj41ZI+og+0m5vahzT/P+BhCvdjVXrPzZiY3XQZQgGEKBSSKh
wam9BSLeRkaT7WW0brjwQlrbj52DA4OKbQXmbXrebzA0CYLYPzNnNwdk4bvO
+5Ull5BrL19LnTZKFvBgpXX63/m5dLWPD7gbm+JD8u6RJp0OlIExLL79xi3B
GyazWWAQ16bmZT6YltqbbOD7oXjsrAogMaIFPxsnEdTxZ61MjX0zf+JTxEot
rMIWQ8S6tEKkFfY7GADbJ8zo9BpMne0vK1ITfwUS9+ZO+kWKQBs4N4ovJZeU
2m3XTaC/EJ7ZDF0Xs5tnImn+R3Io6Y+TUwAIcMAO7HFZkUzAv1oCh4owlB6w
clY1dUrjUldBHGlA0h1vcRxBm+90txdM2rxFRUDpH5Z//p3kpDP7aNV/K99u
jI0ix+KRYarnivrzodlqjmPGpTDZv0EM/3FA9yntsc3BoZg/9CHNlBEgXDSF
M5J1+0he4xaPHhN/sWjLeXlL60u8lZLm2zC2tMaNIqnx0N3YuKSHgTRyJEJg
XhJGpF5hCTMwfj0FwMvj8KShLnuTrXx/tfIv4xh0qAjljAjHxLkqOu6oN+Li
ThU8Cjpw4DD1pJFrQLTm8uwM+wMJYJ6/9WC4S22XQAv5lPzPLXOREaIJG/3C
/ZZBlbEjwt+uNxHM4UNTG6ypoIJnDWgc8chZrtYvYa6SyiNP0rTuAnRXkY7u
+7l6NPLstFbYceKEplY3AJ0qGA/+3rNZ1fo5+fxupHlsJae59iaDWlPUxEFx
kNOffOiNjttUk6vQmM3YrZKn6PBVpKThXK+gY+3zRdqDKGrv/mvG5wHXK2B7
LJEfbZwQ82iJa4eGxlhAiBI8bMfAmIYxZ2FK9+hL+QX2gMu3lFDk/HmJ20pi
QHBZwuvYvZYBzskGy734dn9kdIDLIbHnpbN4hqP3DBU9S0vF4kWXJtzSF/td
BMPnCknfszwNZAyzOg/vN1tFGue1cH2uTt5gmpcRHsLAfoztt5QigFfvoXv7
ZxOOy0lqttJDen9PsNGpD74iCFe+MlMaONpogo53YlmKxOJtItYKOQfAX5Pg
u0iFfjQ33/0ozCr0XuLrxFs/06B1mYas23wt1s9pdhXa5NcpalewFq0LlBT1
219uumhM+Wd8zPZv/2b5vuIJ+q+ZPx3tQ6EVkb0l6RQn+npvd/mWd4kEAMlY
xZNX+fUc88rrN6Kp0zbGgi1KXNgWX+3OfZAbcVe6j6nnEmUTlOubBtMokKYg
EbNgfSpcjOAFYcM8o6dUxwrfAMMHrRrQ45y20kc5WBh7PXqL+EH32IzVEezb
tqp3RiAbSU/kDEEqrld9hShtCLQhotmKut+UnzaeyihDHKMDsVfAj/PbVClo
kl72u3vIA0fiz25TijzCvhUcEJG8IgCO6bb/k6+mrPuU4Sdiu5CtT8shfA+/
x+V+3eht40RoO4H8+9/300IlONkbdJZ1ayi8Lv/dheYtxyVzuODZET//GE7Y
2y0Z+TqSXT1EjUWz7nibASQqepOQ6be7oCtPDkUzEcmd9RtzT7at28ZKG71g
/DTf65eZ6Bov++zQ5VwEyBnFWmcc+2b8L1H7MTocAAkJsTu5b7ZU0+haEaj8
iv5P6nLrfLxtp4fcuUrIrFof3KsZGBenYEksa933NXOi4hQ5n4cA1Ny0mZ/R
0XxjIE2lwr9Uu3yXaqaL4BFNMTnlZVZ9pmaUN4gORBTqACBtctToO+x4VW/B
TZ40ywhDxTSupaiGuA/E84YfrjqQ8z2oh3WMktPJoCp2cC0eCZjD+itpLHpW
0HecxXrPVbSvZ+i2Ae3XlOtki63x7AdWaPAVBxlKXF4n4bNekzEn9VS7zsds
oZhVB5cssu4CKr6nsoBNfJRO51Km8Q4kwqCUdlLiRjzIwFxRltW75Ghmka4a
yFCCwfncF3zrdkx56tm9Rt1KJPlN7NjUE3SH0FBvd4zpiZEx387cfBuzRHLH
FML0n1u/9HBrJ1ttKCls7Rj5YphrpLCQQMw2FXPpfXXhp1QpBlVCA2P/x3yJ
1/Rp1lga1H+wxTHZwtYaOCI628xaPSAcdyizACWB7VlOViyQpr3wBUjMVD/u
t89MrZjEdRN7PhDbh9z28YnGBM8UCtn2kvtpQIz1TolHnLruMrBOuWeG3af6
KIv8X6lqvqN09RGXgOy0+ANWjCKR8M3/0fWdlkeEobHUSFN48BVkRWHK8pE1
oQ5zh2YY5APUJDZdudI00Nk+czMAVUNNjxbi7etpemgSSpZK+ndJHgD5cWkz
dCwONRROCrzy/E9vtKAMY2DGdSZlXD4WlHnhvINKUPkM2fK1RIBNPjJTka1V
IYB0YUP5jWPlD90fVq9V0Uoe05o0UXd3n7H42gLY1cDRhiYQSPHZoJhOHt5j
UbjphrWMADJrifBv+iU587oVQZ6SIkaVre5/9gajpvhCvIb9yHJ/+dJp5Hxk
mvlW71G0k8dohfKngrDoU8EJb8/mOH+Ytqc3vFfF+cbFx4xDdPZDWvzMRTwQ
px7iVj72aOyDQ3LoExEiaRNmarLlntqZ9Ajno8FUwyE0wnStGYHSfwt+NilL
OmVD7EsbwHTSZfgd9UTRENFqtwFvXU2/u2xgsB+agSnTeFzs9Pp45EdmRYcM
HQTwE1oIlaPpBaoWfnTb7bPGuabIx36vHvn8J6KSnBpjmiOuOXWiu4p2IURB
LyL8Nz6xDsYpaPnfar1WN2Zrr/F4VTlIdwufNW0C41JF7NjJq9xH4QSGnq/H
yEB42V1slAECals+rbEwP9jNzRIKsFZeW05euR442jnvDagzJ0hb5N+IuxPk
/O1LD8JtOHUTnMBSL71hUs1sBh50bTN1syJCWn/gI5P/en3oRt1UZfDXvFZw
fwB56WTxyPaRZthD8nL3VmIsGb5oHjn49vMCszDyR4Nw8D9ffRIRs0LfkggO
/cWLDo6OdjqshUHDO03ek0hZ3DTAo00873jxTi6AklfiSwQJhLG22KzIGS6M
ZN83ioigq9lKAnoMw5+PdhLFTcYzjONves6GZMF3wiij3Gh1DhcLjHmU/uhx
5h3ymHpwzaTVuhYAzLoDcANjznOlpCeiU+0JM2QrGjQpNfi9yxOx0d3kkPLL
abZYG/zLbLfvNXpkGlZ0dQ78Gg7gMb740Y1HZOzwGuuu+qUWxUuACzLB6JCx
UDdARbSI6+/I/zRRRw0yqUP2AphXlA1G7UIC/RMku1HhyvHav470v+vsh4uL
jSAn8lwhfE74BwYltGfDzMIKGn+wzibB23JVHeX/chM3NKxDOIMN+/SY0e44
YH1FGGUQXPwWdZC87VE+Wz2eaSNyyPsXLCqUMDjqsdMknZoqTB2k4SiQmjja
J+fXcC0gWpOLLhgAUyeIuIUlb7ESJ9iNAQmXJnk+WVKEl0lqK9IIDdBTfmKe
xrAfEbhOEYoFTd/jOmMLkErZIxGo23xBSg4Xdf5/Y2UnGwFKpfJ4wTxf1ud1
NxJXORZjfAZmKmxGizG1O/VHbgyBTXCFoRpk2Z9jrbRtMsXnSqSPdaE0HEoy
rmzYGSfsYJN0G7th77oigjyq/4kDiwClCwJoC0MHvXoXO2YAKRexmV2VZ00R
GZYVqywJkIwFl4+ze7FW+zeiananhmTXHL2S/w68jZjpVVJPkMUCKEGxZoHJ
s3b4JzLOQrHRp9FsSXlFb11C1sSidW7fApA7hWNRDqJwsprsebRAov8gKdBb
8Ng6OreziCy8ukknBiHqqp2BddRiYK4ey9QE9EYKvHhWeC76RDzSAgu+7CW4
4qVUs9t8oBUSo7z8p4U0YaHtGWxGnqWhNmQAo2WFDxEJk9YO3HtwCdVASuUf
umHcUjSKMKYTpq32vTJq3QFDwlmJ1UfjJNnVpTAX3yQKFyhVXIK+LKrmV99g
g+2e4pCnV3hvKgPDbTtkqgQk19CuwCxW752qcdZCVGuhIjOSl3iSqarbeeSh
bS2RIW4HGxWDG945HHuWsfURG1IwB8yG4yB3pWgdxgXlmqt7rywZlggeYblC
kpnWNZ3P9XphzEUsGjQ/hZK3He/mJbqwrBZ8/Z0R/OG/vPrMZjFimpJicbXD
vHVjoS7eu3Ebu5Q3WCw2lazTxOe6Z3npR9fNtmCrk4xZ4KYsaUO2/FYOkqF/
R1B35Tb/E3gOxFWYOB3rEqSZONxM7tdpNTFiA39xxjJwS+1gldeg9V57pPz0
UalYI+p8sckfwdPWpkLBMQgI4Molh8gCl5rZM5j7Ula7a6Ml0nynhhcB9Giv
xVOsCCyU+8QMvIznEW4vFjjVdBo+8/NUlbXcHoo3zgAssgKPWkvtURD51J4y
r5POFKTOnazrjoGw3b76cjihZ5r/KGi8JLodvHPY5dxf2QIAgzXrbhafEsht
SnbDUYwR0wwDVrghOEgRNiBA1zQkbTVZbgGo9PL8MTFWGP9tCxQFvJMLI7Kf
D+E7+MDRubnzL9nbqbOsJFn+ItYkTVrJY+D4eQw8rzqcIMQgpbxJf/FCuA5X
rIfDCx3y68h4DCIs74XsFiMLrJ2wrf2Fw4k8kqOq536+nrlDmvE4u5jPMChO
vC5xAX+GCbDTA31Zmo7hbafmf0tNAswsgFQ+kb3p/QvPs4Jb7S0X45tznEs9
iQP+lKBsHJodKwEwjcKgxJ6TA2fROVMF5i7yKgnXE0nDpq5lHvMFvlL+FZGZ
yvkUFbEBHub6ApweswYo8hwyO21X4T+DPaJZcREYQO29qkgRD4H8OhcDQmtd
1UtYNAJdjyRqt8VhgR7F5L+Z2WQ49CdGNp3Ogv7UH8z7LLgYsWFoUur3Xeez
EBReDirRgNpaxgPIGMNfH0pwa+sZpVPBf8AT6+sYy2d+/a+Cyio5QmUA0j0d
pLO+JX35RH1cHHPf5Y+c06Vlo7OzVYn3EQ2kW/XfWyMeozZYp5iHu6mxdUf3
qFo3CqirkVmEFeN97ahHJm/pb5RN8LiTybHinLbDro1ReWYEt8+23nJ3zZjz
zv/6Ih18Wlrt67JQZjssqW5Osx8+GkpFmHxAJQtLN7b1XPxGJH1vy661qWhC
EUPtYhX6Y/U/t+fthtzwObX+xuE56SFhQ21mQEkeJV0Vo2L3gwwhUC5jKvJ5
Xjv+KeG6whn7t32onK0spjPtBBYaCkK1eO6lAna674mHZz6wj6oVMT3/Yob4
qxwyLkof6VUE1X14gNzno4VMliN9XSz+TDS5MnjrMQIYJ2BJLJk/U9gmobOR
FvG5EcJt7DFH4ZZeK/OX0AIWPyRPO91dzQa2s3wFbJLqWsanLU9o+bgSsIeQ
tVO+fuT4XYAL+seOGPUS1akkmcGB+hzOKMXhGEluVwmQb1aTGw5q2yCp1IPA
gDg/GRzzRe5DE0Qgepv4C9YJ2uX6LlL5CpGQ1xY/UB7SjPvZvxG3HkQNkV/V
fqfInPlcdGw2NQmRv9LZkyPAGgsniN3EEkoVR7FAUFtBvTUnhA/JDuVU1zYq
uCKe4vs7Hu8/eJLbUf6gDwh6lFaS1FwkH/NFjIqM2uLJQiLRfxPMGBIVzZyh
K3dDPAOF9H9EVvwGUnswThCBhGNbB5BQ1L6JBG9sgIecjkSko0s/s8V8K9rY
/oB+J3HyX95Ea+xdRLNXepOPwNBDvoV5JOdjnhvOzs07PqAAxeSPtT1y5YQB
/i+Gm16US2+eMADzGYPfs/UuklMV+LAyeKZP/BtC9G7EJVkNn81vCohetxqe
sqXbpBKSfvYiRP0W9Z+HFm9hFqFs+eCMohnYfsXl7QQlxDIaNhbVzg7lv4R3
O7DsIznQk356cBSodHwzLGRf9V+JEXzObPt6x3mqZyF+HzCKtzwAOBe1ApYW
YcJxWjdWTgHKaa6apPhGd3vSOZs1Mj6gQc0S84N/nLX0njwaj2YlbnOVEGKn
pSq95hQNns6Q8tK9Tt00cZ89jX4mW7nSQr8W6iy78IzBJ0WdWaiWgGy7I1dS
luuFJt4PeBPdZLSyKY2Yn1JEMCIs4kNCtVXrwA9iQ19siB2BOb+Enh7yAzcw
d1TEVugZyxJBtlqXEez4vzKEjTS/10HQ6JlQvslKsmNQRjvg7gCjcZSrFmDb
i7nNM/pFH6CBMQj3YOTE7EWXvSkopWCjFZjeOBIGuhFHYUjrAUjj1wfV6O4a
leWIZ/bWQQDkcW9cqnpUGBTAvRK074D99EeslwvEyOTq0aV/lO4FT49n4tsa
FUB9ThlFAnAh+h1FiypSg94cHyonZCbhyNe07ce60SVXzXXdFDlU2Lb1jux0
I20frsKu//bcAZAe6IYtyS8cwQLalV+fgdjC/KDqmKdK8UZk9V+GX3BbED/N
L3oCgDCcJ2S243x7z55WtYcFDJLgw9AFy335AeRNlhzMp1W42jYTOJsxCv3U
PMwHNQ2WmiM85CPU6K3vfaG71idYz5+geZrqAhuIu5c2rewXRVUBEIiHiq51
1+JxBfU6Dpz74J73Ps3h1ykatxv8aWCrrpz1nvl0bvBtHE4yKzdiUR+r5RH6
VWNuPL9R9HqiGInzY+EYQ3USyRKXS1P6ias8Vtd/fRdkiNIPKxVcAdXuuHDP
fib8FvWeTyfJ4aZr8CVsmuxINmABiqVaRX+Qk7iEMcVGOVzyOmCuSAnC9jtj
sJOZStyUHO5kIhRlWW2bPcxFylxijbxrFTGBTwFjfurHuVyUQ20FFH4/IH2C
+Vi+LbSYJiqfxUvXzcWZTwmjtzTD0V/CdQU+bsmAW0mCG7XLEBPG9KHl9PYM
grGLeljjcFhztazlH94IRxqGiXKgPpr0QBbrujeZztrwafoaOvV6OMFIs18k
VwLYvZuP6GrWJ3Q+nBNTi+RQZPvKA6Ep6Pp0akxFHf8C2pVqWIpm5yfpfOjM
u41Ga/jKAJ31rCDr0y6zKiqVaWnNxqrswj//ITZiB+x/3ITdgI9h0TJU/FYW
AvTOZ3ulBRI9qRSV/jrc5WY2w75zvulfASD7eV4K1RsF1WF5Do7MkhteOoti
Byrgg6xWi1kREufpZINGtiudiueqaTAt7OnDMd/lOcRHvCAtZGNySKJT6tQM
Yjgk8PRj7G31Urs0b35V6tjGIQM6W+jG7mF1plJ7h3LC3EnKBV3/r/Csp9LJ
vRwIDFKFRYQYrq5IDbDSXmu4fdxfDDawMP5gJBCqm4Oenq+h5TLMjQYSHa6Y
yHE2SMfuaNr7A5KvxLa5IonySUyixFtgZxmTjHrQsuCz/DAISYD5tSWkikV5
pJieyCD80wpczcvq2oyITgt+y0LQBXimQaVUNMglpjbf2+unGpeKDSKPUxM6
GYSmbYOTNbJDDmuDP1NsRGVsqf3D4uVsKdODai3JmVd6WbV9F01BI1eENv8B
uWFGBh3x8L4XgU2Y1cNqaCp3ZJ5dpY3fmYLVc0x87GMK0MP7lUS28kSxSglL
TRx2DS6kIwhvXtyDZ3NcGCBjYf82I3vgB9GbzYjW8ZNw9g204S0mhOSDJkC+
2/xjyBhLQL2J/7F4oJuYeKe2U4vLFZNl6ElhMa6MWBYyWiDdHdFsxx7bq/kG
7W5gpEvRpXCNq0mbF7YGIHNQhiSdbQ5W6QlpaKlnGLYiA9/bU0XAUpyEKIM+
MHB3wyrqnOqYzDc8fe9JUgvTniFzFgxCT0tusUZM3mRXcNvDqwNuF9/ThcrA
HZWU+ZZqBO4GoZoA2kzEnT84s3pj34l9UJZjWpYVugS9LIyQyQZeSRfSkkiS
yNgtdrHlRmV4s3v9sss+Gw6JeXQkmQUF27JLvUp6RSO8dGb6ogqOwhUmrdcc
xyYE+hX4/ZwJVB0bn2WZ8JN1stYAXOQPuDqozcVrmzrBP2quXHMCe8ulVTMK
XYWi6e4cYXfIijgUksCGiyJY+6BJXbihWADyAm4kpTHcIax7iIJkptgur62m
Q0vN39tDXvTQFFZX+KEm+k2EaytW42A54g5sYAHZ8HonDlWKw7LfkdPpq0nv
scy/xom9MUTHrsTAPv/0+hnZR4kccPAoSwe1o4BhdWnlfMSZ+mA24J9dhQ5m
bQC6qeAJtQVDOqdxvpVbfwAIqx/hXC4BzMnwZGKOqvpT1XMOR+VGba2/EqjS
kqfmEgYehBU+pk+Kdiv5XV2XwIn0LXCQxmzshrUU9aKShYnoUytO3q5GDqOi
i34Y0roB7mC6CEXqdkoXvLCj1hJgqFBRAvHzVYduVEwKGqqMcS3H0odJIpxk
mhi8LPJSPQMhmeNzk/NN0pOklI7J7Zmk+lHcbM66sJgx2CzrNpqtyK92gdSn
mLJ1yj4llVgNBgNHQubOYVxPv81lnRecXXXUiFivSSBXGxtEZZbUZMvVDpVG
Nzjg34D6bK3EhxX/PmRs4UloAnfkQmLpMC92cVkU/wFuxMzJH6QPT6KQh+ed
s3g/8qwJsRI2p7W29d7KJqOkGHyfmFyij3bQLtFnO1RVDIn+wrKtVffcphwU
1nuTa0YLeVIlbdzVvXxH3IrHKIqkbblC9FT1AA9htFEb2q4t9qC7kaIkMxCu
CTZvyrjgyh25WYBom69N464vZgC9cTiFYsw6InC4g2gNWfMdH/0LS3VoFLKQ
iTpqKHDCzxt3b5ddPIunocz0etkB+qaxY26VJsbRYZzMHAPUoqXrVFHX4PIt
WuSVXwLkPAKKRh5J/DzSN8tNJwRkTt3LKpbjUKQiz93bzBA7wXgFNcns2sDP
ty4Lml9dxH/WLnsNv30MRG/XWw0aVlFHGSztpHBYR9NABiDSoWBGL96agjtV
xgR3l6pQK8NK2lbWJDpIxHeRR7g1amQwzsOOl4qVQ0k8PkV21d0AW6L6Wubs
OIPbKb2nXJ3AI+ED6QvyXismeUn7mKaigyUOqGJh88zbbmoO1fYT4p9mVJti
antT9qeEZL0p7efoGJ5WaVyvZ/LMw664wYqs7cQmFBUwuY47AWJBbcpNmo2o
ndghszO+/Eo0CFQ9P3dFbRSVQrGCWwgo20pAx7Ai2+X9tvP5Yl9R7uyweZ9m
Uf+ssqGYfT+ZiNb0YJAsd8kFGomWMgp9FXvQBG9ILawfR9Wxzx5e1trAjPAS
wNZLrI4wz5m3/iO0WPnOKdln/WIGegbg+eLpoEv3nDTpQdbhJ7HHqFu3+IUk
Cg6hkNFe3MdztJRgsvLa7Wsf0zXCKTttzmEwbUH6xECtLuyx8CuNj3ZOFlFC
ogtLvUGS5nY6so+wdBg8ZEcaAkOZ70xD0GuDYMzp1H+wZawCYF47+igVtDCJ
zsGpeJKjnQIi/eThC6fev+CeeVOmhrzP2yOZLr2KMRATkJFR7nwPVh00WOaX
f07JGaDERQnK0JWMJPCI3oenOHrhK9FP/5tf9u0jB0AA7O8Gm1PA5lagdlc7
1NaoSxDxFuuTVR4+ScZdGk35HcBLtSmo9bW1ENUx/IRKxJxD+6EwRQqEs6N7
sXS1UcHobL3leO8iWpev+i1YEG/XukKp14Ph7ewjFA36PcTxLlFEPfdCNpEA
Kj2KMu1zXDoU5mJmLFO5u48SL1WfzLuOUHmWmlVwXXM0EoDYvR6BjBYlS9qq
OtQwEbNPSZt7JJha0I46dAV4vHWLH+QXVMfIErFxCAZtwcU1izDtpHffOJEp
Q5v55aGaA0bNoIKt4Vy5HRShO8yBerdhCKanCXRCkN/zWUiaadMDWWPp61F6
hUPPniKzTV1/pjmerX/K7oMMCyLBvI8Fka27Z8xda53YIMP5nXi0P/39X9cF
0D4ij9wy3C0bnNssAZ0O8zdq0TlxNXP9Qlxha19Fm7G+YmiglrZl9+69W/n4
2jGhmv9QqIbzUVP5mII/IXWy3H7L3hXFimWRi9PZ/tvTSsEWHe4D1hSjPcu3
KApx11GtsPIRc4ycr0I0kb5Nuhl2xy9f5CiTTGTerprj9RxKhfALK3VBte1u
i5vmXAMDpr8KVp1SxlVMCd/o2Qk8WwRPOjPud+Qy23syrVOg7/YEpWQbZyXP
IrvFOFZXb1J9hJoVLVCvuQvhOq6h+27Ci78+vkL/amIfE28o6ZdH0pHIXwqo
keRn/XrQ1K2/5zhem4A4duHa6uTRxyJJ00HbQ3Sq9evvdNDznmCwuQD5xsMi
Ls17ENFAcGMKjY6e1w/rPSvtqOQduXTJ3ss7uTmbOzTmXtSTxOkMHULLOOxh
75ww8QTTD/KfWhMPynfCKQHgaueBExzg0/VfQGMjqvjxpoNkAUyi2NleYviz
TWOVKFRHC3MrmFeD9SJ7hex44KoicxXjvJHYWPz94qdfPqS1iRCsoSGU/0ia
hToPbuunc0gDGiM1aO6DOIjmDNehD2djpakrqqs8OTSus4KTqr7vgkzrmRqx
Ho3j2jM5IEt0XTyrYoYT9DB69F6k32NOYhgl0t3TN2tIGWf3o+Pe8a4H2Ffl
wB5qDcdsAW98QPrHwQBXNlmPPRQ6xGzcak2Q7zuWTMxGV9evBZd7JuEgoTDG
442mHQpFWgvld/bRv62xU32tLv1E53250xkhGGGh3cuu6K45nIBG1IwvD7dj
xIMYAJunU0J1vrfwyEcBrGWJFpUkSZOuohrMUM2riIQrk5MhT8Llst6F4EBh
DUBhiU9wdEiFBnGcn4y0XXIc+1f1v3CZRygxMjG2Q790eB9DHNk9jAVA7M3F
8KNhh+C45TmQB4RggRpJq987hF4mvuxXMQuZXgjO/OE3N+T3uYt3CBf3kxTi
TAh8j5Nm6gukfOmAbL6JtZ3YuVMYs2VpLzZs9vBbAFMq+SG2UF5/DQHb1yXl
0k0JVOT2CVI/WOYilptz4wvQCJzgmK+Qf9SkjMYTsfuuj6tEkn6dEXg4tAc1
Nn3Ax+LFvpoqIWRXQY0jozNsqzfkUpsmDb/vGyaqWWiYF1JnJqabsTmIsheL
MQRXPqlfMZXX1Hw/8aoyDfZzEYcHvr2qbyrmemv6NC284Tpeq5zJildgPQru
H9QykpNUgAdWK+8rivDGQt5DIvTz43ubZxez8IHi7mSBEPCtdHWFhiQvHy4z
qW758A+3SakWXJeEdaA4/Om8UrQ8/HgGl3JkGMtDEAxIMjJ5GSeUDrpPq8MN
XIMJIZ9PTMt6yNabmJEzc0IGCMEwBvcXVj0EUcbI4Vjm/0LqRCv1i2R9x4n2
g/b2uTkHr9QJnULx4Y3oQ6Q3ioo9uFKVH8YlvO95TZijaGg7fQA/nHQ9Zl4z
tK5DoCq8IKkkXtXS3sCFIF2Mn+2aCv4wmR5LnR9QiR21wksiawEsroyAnIsE
mYkb8U0CZk0GcX2bTGiI5UTZvR1mNriY5bN5qdRok1CY5WVmmDdwz3SGQ0aG
/4bRbxj7ydYPRsKrfZ6WMHZ3/OOLLMdYEgWYh81CkOQ79dWvq856AYo+SHX0
oRxMsiJG+XVpicrQvOPhnMyfdD0+fnbNuU7X5CfqFZObXxd+gm11ZdD9h7Kz
taXB6ozMU46SE/Y4knWDc0aToWuIDYvFn2kgDxkS4xoGJZ2rg0DpWOIgS0i1
fnqSD9Iikvek8CJ2i1QRTVvXWPDhTrWDyFU9Skdu4JQEetQhtl1Pw6kyWM1M
kAx8MC4WL4L/oeGVw6CXd/6Ay2VDj6tWG2nnUgMWaXHSG/Zgh4EILTtKcwjp
30iHpv/50eD5AMRNFB8rbXA44bBNG5zqfTFpZoyQsxELExVsZEXJTdE6XplS
A0V04fgtm7l4upvzk80IQJ3yFKSqoCSXS2nbDfkwLhsHCf0ZteXyGerC4E3h
+Kwy9e8cM2ZQkwRB2E5M3Uk7DM73ZjfS7Hfqx5f5a6SGexYvx7rU7xa6wpbj
ijIwcdSZdK+NhXzZ54U3XX1yF5KAFSLfJdT2vSpuuBlVNhjuHm9EmeKDR9+L
030ev3pEirQ6k+yjV8s/7Hrlc3zwYsAgd0SMu0tI9oGlZTvP6VmX9cPC1XWn
UAujM6uWx/SPBKMSRLMfqdqaF+SrvfwtG0Aj5up7yDBy+asH0nTtmolKYoCy
KlpOFyvycZ0GqhkhhV6E2AXmW8sXN/JjGELq7blbdQ9DCIYlNxE3fY4vl2B2
TMUoLywAWX/KH0MtXis4A9HpjfMEm5bcJipg6k23uGXFJ9Zxtg9WYvTdF85V
yBo7A4ijARBUyOlMMnEDEYL1GiEdAbDBqk/f+CnJdlSBtSdo0pQlx5to6deh
DPEYz8WQHN2FEIHm68sRFgw0kp+Gs++BTXdWnz7maf7wx+sVf+H7d6j1AGX7
SkvMsE+qSP4l+TA8QW7z7CNKIhTpbpWwH2M7Tk3B7kdNyAQPaBN3I0CULQ/2
sIB9kVCYrX1swfExvW5fd5wO5eudeRO+3H4GLOHXmQzijvYL3JBNhQRCCjIS
g6aVegqn8xXbAEyQ0mOa+gNikGtIa56dishSkc9UVy1RCQ/TFVmycRGRoceJ
Ju3cyrCXk9L1H9vNJ1ZF26LjrFyCg7HZpCbEYzdGZJgLDlPq0eKjdz/axq6l
A8tjttsuoUuBDZZ8bk9zd07WMN5yKKf8MZB7LfqQicrKaOGUpYk5SSVyCRhI
eM3Vy/M4gUFv+IRAwICkKeZ4RKFF3vXvGTxsMFPnTZJj1eB+r6OT7WFTQIfs
0geFsICOZl84dQB5v5aFZwK31wNo7kFMDq6ul3aE6XSQvK1L7jty4XM1ncrc
y4dmZMHQk1MwVLlkZS4UtkPCa21d/XeS6FrkBlFOBmdPZ9gr/is02C1wBAi8
05Ye0zHVd7gzw/Buu3eV6hICVaPixeIUyvF0Cgdihcd4gbmDMEfsmKyOHhPU
iZk2zBRwRDyquFywzNML4o5w4IEDxoWeRzkN4psowg8+xc3jkdr0eL7/vuAK
j7vJ9snv62Csu5KVi3/FVbWRWHAxIOx/ctAAMolva6YBXAwnsGmtcAVqe18R
yxSK54X87fo0Mueon1VC7xKUxrIl/V056wIHvxWokXjDXB7ylKBPPToOgyfo
ArQqnPWAhL5wtxe0n1XXDRNixVLSWosdzp5JRN3vypB01+z4txtqWrh9tr/j
o83es2faNKOjPoFQRY1AvaKCvR4belgScuiSS/sRxypXFiZ7Gv3C/0mqIKZW
0MTzWxDjOayoeUgkEE+jIxKX6gKXb3UwoO1a6Sq/6oRDPIb/KkLdZLJF2D6Q
40FFAChHGYyNs8AR6LzzU/Qf8fKJUNIdroh4xSzOoECAwiNonzmfNn5Q0MgV
VEbNRDdHs3ZAjjsOYhoJfI6LHg2wF3xuDbIms1GJeKbxnPCGs6U5ibMoey6r
BL36o0woGA5u57cH4XjxqQkRgE/nW3tzUIex6fh4LYv+iu0mvqCF2TwAmYNZ
05NZM/xhV1lDwKzMi6E9+DHzYO+2Lkbhw+Dw/fQI++v/4CYGQsZC8TuqXDhL
68r34m2u/rV/uIh8ozv6NT3CohD/WpkC2FwM6KLDwldwrzdYWQdAwr8iSlRb
HURw/D1m26xLY5VqsPyt7imH//w1L4RChd8c0j4SEKZRJIjlGDlRNiP1aQlg
b4c1ODqVQ+Q6UsiVN95SpE+wwYeSpjdSjL8ZO05Js6ABx+Q/ovQXrgagnPNI
MJfUd0LDUbG82ZX42nuEggz2An+84T3dmMPEcLqwCDZFhkVRODNVL6FSQBUG
C0EP0G2vFAPpQGhmNmtbO/O/d1FoWiOhAYPGy/I8sfYTVKEJlZ3vq7Db4tiy
nhC4gHtPdbpKfodYRI6tdL+rf72sa8RchZtku0kidUJSrgeGcwyC6tEzQmIu
nWEY8Ky8qPH1J8LBsJ9P3PJgB9zqexucoUgEQmmcZtFNBXFkYtjP09q0ATJd
Iwe+TLpjLlul929hAx5fYILF6j5TS00xstg8nOuIAd8OGMQ7Dwb2s4YXxCBF
wK4aMc88Rkzdtl5vfvoT7LZ6d+1XmtSk2ghfZXQJczJZM3MN9B5POF4dBLUw
EdyHetQDVJUgFUcT/KB1jRK4LG2BXikft5cB039fn8p4e+/Ir0SF8ZPtq0Ev
qhsOxFp+LjXyJP3m5lnDMY4TWZyJVD+sqKqcva3eKrVldOEabVRk6Yxgt4gr
Kjd7qh/XE7WD5r30kOSNkhFRLA2gYZx8IKdccBuX/gOpVDf6yRlhizvMTX6q
cxXAMQknu3KgVSGOb4xWvSZbxQn+xMIwJRHikhyduU1ECfpI/RwIDxA1QNWB
XehD0Eh5beraTjzPJ5bQjd66lu/eEL4fUyXQ5UKB8VMkUfyuCfg+Nq4bzzkN
WteGc1Byv0IjTVFBMkKaGcgS1kCHe5mkbSsf9p44xgfnBAaIYWqbjZeSRduK
WJbkSx2OmItGdY9CUlQY8AgPvh94dKAIRIaG1egKCCHBzveZ6oSFNEKRw62A
hbtiwQGrolb0/P5fcGu99lh3BlLmOWoMEkdnTZN8atTfqBNchwl7OtowvTU2
AeMOXJo5Uvc59DNAd9sKoiIAeG/r6uetlMlAGXSYO/SX1y/D5oHfamfBQG63
eRuUZ7gsf61HJH6i21Md07wbmHTE9UtykyjC42OIMn8E7n8m+oU6dLqh5K7G
uQm4BDcXIlHCeomeO53qrIjIzEO63z1lQ3E1wfSFIJt8ilEQhIJGzWb8rtIe
Ja69UwRaZ4b2k2D52O+ZIpBF8wRMMmzdLID7mQTDbgJ6oc2yUYlQcITYwmIR
NiVrQTkxIqhx86IPCzYo6VuT9w9F/BQXKU4zMG7nUDdQEOhkQfoowf1lkq/G
rcoIYL3O2VcqulM0dMsiwS9Q4zRc73MT9foMNYTjIsF3/d19U47U/xbyRoNk
P87rgQzaEUFITBEtDaVdpZdKJ1uwCPI6yB1pmQ/FVEnp4RNh3THyZqKMDP8S
1GyskRRas7M1N4f+YZE9mM2b46IUCapC/+15Po+UL3/YsCahk4xQ8hYcWh/T
jHCSP752x/xWew8PaCEW7UMxAXgwCJe7Pj6nFC9uQUszgKRYmXfaKd6fcJTI
cYu037Q58Va4bkND0z0gzgYFqTEKkFwskjAsF2xCWRVprcc/LXbm+8rzyU6Q
+9hi6u1ulOfZv3JUq9ZQzgl3R9uIDtF/sqtSFOC4iP6PB6HBFWs06ex1bQGH
Bt+ffP+xC+1ohpfk7JcXnV/keMIvfCY+g+W9KVlORFrKqZCOGt+rGzkfgwzo
HHNdAIGj1AtbHY7QMgRp31A6IOLnbG9RTpTH1cHicywwyM/AhsmKZ+GOUSuv
AfAoXnbKEYjH4QOpFASEHnpyq9Upo1s5modGYJgngXUz7vC5a4oLRsK10VAp
AwU94yemwm1rJZXnyo8adzj8g0rOLpEuIQdvdyF8s0EYmf3pPWMOPFO6hizP
21FIOUbkClEBFqcdCGWkC2BrK6IISP2ySy/ePaHIa4niu9xm5gnrMZqSiYsp
Ka1HBEHWmSwTwyaBH29njcIxAYSgl9eMEnnJiYs9b3jocuKYVnFAzHIa9scJ
aODL4fDDJfEC7YQaMmCfW+M1C7oya5YmtscCKAGo/E0wkPhkOcD7+2kWWBKE
C6Nr1drjWoB3lXz92n6fttctZ81chF/2HQHwirnsN1jq8pjI8luv4ceHB976
oyUtJ2B/xHviwlx4JKMPzg4hXPrG/mVEn8uiDeeAJEXWhZNjy4rWIJAd+O+k
WhNjfFbx+wO0Fa9Y7l7KH3pAD9ttdEd6HLTVEIKJi6XVZrbKHmu3WY13G0rw
vnN8ftIH4nbJydmYCRv0lMi99In81IGwxeyLIqJQX0C/uavUHe4fiKj8R2Wq
EVoT/94Vjx5cNsWv3lpbd0qsIwV1VDhX/oy01NElM73SrBFnBMHveTZVlufC
l0Opctqeo+L99TSKb//Tk00f+dOLoyE9MAEtz+aH3oJ6UWE1DHTq46ZzD1TW
R3wzhzDJYYzMGubAr0eI0xxZZr2qdwZuKlKKgq+UMnzHeL1TqYbbcRhBtbG+
ccbsSsFeG11rhNO1L9Az83v/OEbJPDIlTDIchBeuAjTAlWsohHeXlg77LB3V
b/g5iTAy12aI5wW5Jt81IVHpX79IvVCrITQs2oaBZv1H1XXLzIdQbgDaECwr
4Qo1ZMAZO/poJCgA7fDdtHMNSsKsGIiDuRyrNZ3wBWFDaZ99jt+y7LL+77G9
ta7tXl/6agvQtrvRxXroPePTZiGD24UxNRL9QtWGqzc4DD9OC4Rrz3IiWGR7
OlPl0KpTS7rTHs4Mbs7Ezj8o/dCAlvZSZP+681ivZjCFYR+fHrvO0+clcSm0
GBJvD2Sza8TvsqZL2hgnIEJo5YqAJwmw/eR61NL2VYYu2GEQmvSrP69kglCS
kPnpozlcVSLLACh9EntAcPy29Kf4Nmm6jJ/uVD3dEWb+1frhgsbF+kwRK7vJ
PX+gpsOxnuwN5/Z9YEasnA4rSnE+5YrwY3pWT1kHd0vvQKuYLLajX0+P8Rxd
clrRGZhF0XvqdH6rhk+Gg8dFePWNjWGcCf2RQX1EqQ6FB+IbPMb3K+CNKsZ3
FjGuO/BDNj+JR8r12b+NZa/+Bcvnb5ga1W2BHD5VRyPCRN3TVETTwupdtNsZ
TlkcaQ4jDcpn3EFI/QPSpfC/XrKpxOIS1YnoOsbeextcmzBTDP2KJuk80GYJ
kZ3i6GkWdFu1C1A23j6UJIoOHJCYj6YhWGceMwBcdmOFn6RD4JCTk2YVZ6lM
HUIDYqMcq1A2wd3UMUDB5sR9Qh3kpeFIQl901Jkxc9pP+ofbLT3QAiNuX0M0
YZsB8wNnw0Pz5DABngMG+p8gVFuU4mkq9b0goMf/Drdu5bhK2mRb/X57yc0s
yyio0gW/VXNKV/XZApy2otcGAInlE8FA5DSnEgKaIVMOvVexZcnWwaZL3eQT
KUzUHj2vuil3EOjryvV2ZNs916A5jBx015P+roNR43uHgDF1Idxylgt7iCIn
Py+DlerTXPqM4HAqedBYKb0bwDtDT4NBDdeybsToy6C4stIEql1UDqwMkKTi
5dPtpWgnCvSsHRs8WjyNrb6MqvbpYr07lv5jMCS/hCKzofn+wolyPv+aV1d4
LSNGAvT9dO1ajlT63tlocHV9V1zZk2O1aKZZRwwuq3zzRu4bjfe4mE6fZDp+
9Nwn6goEbR2xkfm1bFDc630fRKd2v1M6YR/wCHRDsXggkJJJZ681xS432+Tl
l7EMPZsroGHtAA1565GvL+xtHXE6rB3CQcgaHJeccR13pmv0f0Yd5xGxJuKE
19YXX5vqYs21aYeZmVEQ5r472ZkjK9AMOcWJXrK34WFk20uuNbvjcUTdeAGW
GXHINzwzsnPONYoEwPVttQz/1KihZWU65ZvzbK5W5Lt1BfGttAAAS6uYhqFS
SBAd0fGHpvU4yrihx35aZEnBeOKrqvJnnBFV3QqEbMt49xuVBS5WEYnWWZgy
WYGKVaXxlf1YOXSQE1YyWtQnCGelNkyOpt3hNVfbe1nJ4i29NTBSlj3VBhcQ
vdoswOl7Fvag/dKvV4cohHSvtCtqF8n9c5r3HEv+2ox5QcnEe144XpPC7xtB
Q93kreGVLRBlTc00KTfULu1YeuYXvPmBS90wjSrWeWNqnFnbyX5DpBVQWZSl
GuJJFxKMUvS0F9hOcm4VVTjvjlHifZk3ZnZD/S8mDwwH0bF7uxhGCxPbGfkN
EfENBjiAbiX3ckNxEL7d6ovwyKotn4qZE4JKXIQCCk6adAISR46a0nIhCH1a
AcGeLBaC9IABGnKXEALzXk0/5k0LJrvd0QnmMLB7E4OMQCCYkQgsj57+e/0G
Z2ZIPmjo1XQ72MShqmhwNQFfVrEo5OG71GBFAKPbnQYPSnPmTFYQxXqavpWA
0m8NtbB32dT2j2Ndn9PVaTCdNJNIONzideJDnw5Dg9YHwAdVXLiTe5vIse6Y
2FU76qh7ByfSpWq7JRuKmjA8cUlUwiGbmNtvHHzP6Rp1qCpAtCltCiXM0VjB
ukQamJfhoP365eQX6q+4iYB2qLhyWsAi/5Rib2hdBjeqAUQfmOUF5GgIjsIx
7L4IZuGg0/wtH8NzbKAcx9juoP0kMFpPMrcbuQIbpBwB4E0JE+oHhMXZqb4J
2LCGe7eCXoZvsXFxIS4sYXuXkvH43ONfQjft7YGC/8yzWxenvQbuM5oa9vK/
FVVKhUAI7qZ4vQbslD2wyy1DdXo0BXyXMFxHhAU7s9tj09nBuyTL91Ja/T5O
2n62Eb2ccXUuh55aotaLKuvNx5pNavXYtg/rvesjCojrTP4M4EPNd88SpLSI
PvxFYnlPV5A9oGZHFCTK9tHBqFqXt8EjzcfLM7UJVfSDgNZDxbbDu69Owepc
kpG90T9YvRwsyWFyWIObLPUT2iJK8A7lIv6hLCvkILajudzdyBAOTX72cmV7
Q984UoDCl59MQJXDVwcsXOs/MUowzJmavnH06ztuI0c0rvVq0Bv4wMrFCM8H
di5dnsMaY1RMWEBvC+PtF6C552aqqdrbipVbk31eNig+pqTR/hf5/qnRpAwI
9hb4vlwbB3/9w4pvq9ruwiklgGMjxMFPZhSbuHpm6ctlz9X4b+x46pAThGbf
9TgfhofR55qY+sLNsc/xOu2SX+Zc90r3mN8pb9cm5ok3jz/ltPS5JqlBxZRv
B4OqVjeMCdmsWSYLdpqd9GpdZYRfRZyVs31kKb19ocu4EJIzFhq69/HC7e2I
irSXDOuBgpIXYHMZRZtmXm4lyuifjtH33xWZ9xF/ht1BNkQlOCpzt3FyJtWg
qPZcyo5vN/2cljl1I/7Olax+ZqK27NYXfezU2nNwxdlhPMkOqAfj9sEDCrsu
qE8twt1kRyj4WVrUJMTtUpzYb8ttYtMmoML9W5GroLRVKyCtNPkmSkY0IGY5
yd9F5XbvXytokqY+hmYzkiy+h0o1Ap1ZCBOgMTMVYQGLnK6WnEEB9/sQMzYz
ja90+Z8p910gJU77nh9Rk9FTsN34u8HkhJTKtP7JlcFJ8QIwxyoEXohu1PW1
hlvK1RiRL1GLod61pXB4PSMx35IHMr7CAx+bTSfSKoLN1LSfrkkEfFKLo8wv
eWISKxNdhfeD2uF1iR63PDNNPucetIa6rZ6r7YHxaMnfJKmKhd3r5TvaaMS2
wVD483EHKcwwS5gq/zorxefxdPI5aLIrh0ju2mJ4yeDzlFvA70qcomj6611B
qMhLl1fcb0GUQdOqvybUyJeXvRTCEzJvAW0GXMmY2OIC5SLbWx4bS40tEdO7
nhkHbm/2HVDNImUubU/juxiAdBLTlj9BpSMxEkRHhfj782Uaqj/l8NIDUXpm
lqA5iD+Ccl1WHl+8gMK/J79/ZaZcVbN/kPabJEEe98QNZmtEbv7c3nU1Te/d
MDGeEyQqrrhRDGq0rEX14o56qLmAKVMdD6hF8x4l2s+Z6Sh2LkLBu2jWhakO
0PYA7qfqr465eJGWtg5Z26av7Xm6ZoAln53vNnb0j6QX9xMMK4b3CTYDdpQG
uGT1XAK7rt1i0iPHo2ZlYpp1upCtXvZfNe9tquSQ7iAWwaj4dWTBDYw63WCP
MtrajfuSOjjuZknAV3xVw3MkP8+ckavD450fqu6g3wlOHBwwiaoxFMC1CKcp
uSc2hmMVLIYRuuVd5//c7H9wSMuLh9E+pGFIh3fD22nQVjBXdKzVfn4QiWgV
lFhGKylzcxqUv0tBtS5/Fe0+/CRShMhLeYsVfVIXTli+Yl5ep/JqoWYzFCeh
N6Fr++8XfOEqZqSkZeLBXc1/jsOlk73GVsJu2FPPHQ0EQx/xIgFyOLsngXTn
L7PCQv4zK7xE4hdduPEfav65znoRDXiEqeJ21m/87lmM5tETFn3TmB0EwYXR
oKY6lVPLSPOgXyRoEWrYTvwbCkbRj5rYCE+4Q3OAvqtD5paXSmypz5w5GkFk
yRdFN2K6cWEJxHfhp+9lGj+FwvNOTbNyxL5yMzhDn003+Zih7hZglr/5rb4V
aFGu/1/oQFqxHAX0ODC8IhHK7x0UBzTVhCwn0o8pCREk+WBgf063atUG8H1d
BInasa+0M+G5ezjN9ity4F+Kj6KKVQ+p8kYHJlqtCUI+BdLA1iW3x/sxo5hG
3OJWuTAy1Ucj7PlUZ9XlI9xKVWzmLqB46vhk1WhcQpNw3rDBoqjcVHB2iFbz
cfvdOLNRtj9cV6lS+QSeTwWL1dDEntqLj4rwO1EjwJrsMS2knPnrfEABskz3
5TQMq6oFxWpzA3RqUATcxCVv6zQKdCJnTpZiwd+W3hUfKhoRcRjEp1BMEmRD
zhduPZ9kMgaLNy1NKU2zFEO/q9eb0dnUrtpYHgScfXyp3exNLNN/ywb0iILV
eLE0Ym3SvBfZvcewrpTjaN1UmAMhbsEZ1izyp1IJsj4yK+pOTcvzZQBFnYO3
6RL4QMbTcCjLYDRjhtZ6fBExJsDv5p02aRitK0X5ZJT7oMbG7CBbSQ3NpvRY
3lG4tvzH6B3sioMs9S1UGaQmK944mh97WEiFAu4BT4qHU2YizXHC2MGWuT6k
CMI4xA7PxP+O0t09DXVPWG4OAEWljII/IX6s1p6jaynnYHJleB+nZ0VF6bG3
nFsZniutshflZTQ10STptGP8ILQRUG4iOYRCkzyDClLcoELqpUteZ96m6zp6
ILvYaD16mk2MphlD6Rv1Qk7QtLRRtOULzfQmhjZhow/mPlTTly1HperVkw/y
vU4hjGQ4a7jXn0BN4SsbnW/GK/LH23BxtBF9WaesYfv1WR86mi6e8SIDtjSr
AcPT8cJ5YLQTRbfTWkq/omv7+QKez9rY9cq/2YsXEza9NvaKqHAao2zb3t3p
bD4sBxh6K/myyXhEyxTqx9WvcSb8Cyg3lGUPusdOkx7R/XHyvPpD/Mj5qR9W
ea27yeP/qZawOBBdkiMw5UQRSzUp/ffNT1qx3GPggqsL1YbsspnZ+d/FEteL
v6XsScZd3O/i/jz0LC1E9ZfEx2Jwb+79cSEoVFqCbWKAIa5SWJsIp3yrxeX7
Dw43cBHN47Bxd6WkBZ4ncLUgsQexXDCb55zoe50JRpXNJ6PUOutL951qqKD5
hJehnIWiLe9dZaOZVmLy8GOj2P8kOy0scm+mbhTEA7IBG5V0kq2ME3vm60F2
w2CQWEMpM9/rXCrNj/VtZrD8E9ujLIxIgP/VNJ9xBz/NZUGbdwuG9FhyzVFH
KatttKgUQ+39RQIiRWknPqJfhwN9Nh6Wze2yhbj6pFJf9sCktCw4oV4qstH2
jqaRXC3zJLT8FzwmkY/1DSjUeRwdYMHtNofz5x6zT/qFPsr9k1g6xPR8ULIx
E1A5Wbdg7Pd3FqMdojoNIRSeQUSLx/y0mNQV9As1DUyZVozGZZJrRWAV1wJs
u0/ZFow2H+g3EihwydPF6OO93aNzE7ILpuXFuF996qcpLGmI570kJwAjhzY1
aFvzvLGue6y1LoOxomrMP3mfnCv8BEH02WgAAhy0HDSgekuDWE39+UrJSaqT
bsoq6yMETVMgd09I41ocBGLKkf7DyDuvb4z3qTFPdqst1a56BrbSxHLv46N2
A+M97k7cwM9uZHoZm3xqEChyQhtGiscfH3NdfYNuUzLm+Pp/4a7I3RM+JGfQ
3DPv69b1DaF8Fr0xVXFqO6ho7Q299bYfojImbNkZ+XZPftyjYCkPILHX86wG
j2l+T1SR4mXaJuQkthsT89n4WG1wOvZao3VXuZE1QMBpN6KUO3fOPzOWMDz5
Z+VKyTTGKFarGuacCt3Li8juBRtCj0qqr95RPYMp7LZONN1eTuH1t3sq4Cro
XDPn4SxqiIvMxCoBcHTyHlSek1PPh3Dx2hwbevgWjaN9qhazEd4nljLZsjrE
q3bte/CLZtlp6i9GX3y3SB+t7k7Te7kA36QZuAO9gVwz0uZ/7ikREXxeA115
qZ5AI7L344KZ5hF55KgycR66Gmd4OcPNrKj2/Crhd1/mcAj8IC4m6QIwzkGQ
EqfdhnHnZcbG9Qgbj3zB8YJpumCk79zKjAhokXMFzjdnrGC4RknX+b0WLlfJ
YTOopQ4e0pHZ2WIajut9zdpBcrh4Hq3Sd/+d7/x52uA94YPOQy/SGGe8bHTs
ta3H9hCrovyRoue2ewkEPzR+DkRDF/GHmIRGU3qbpZ4oHCGJAcb9wv7WA8uM
Mx0cnh+tti+3AwZ6bzuyI18EwKb+YTQ5fCX55lhVhXK1HKZjTKGcHefRYmBN
Zo4nnJPIz6+J1E68toW5KIQDI5okqZlltWUGueaWbFIgY36cqy4GNQQNbQjL
qy22PHgRJC7FLwIXWPtvu9lmzWiJY4aDlSzcZXBarHWTv237Jagly5psqkh/
KZ7YBB6p+3WMEQbk2vJSuwID6cfkbkp3aKgT7B9H0lDWCtpzKDw1pR7w/vpw
ZNjPW4WCv+rPOps0mjNpRtg3XdEpdOPADA9plDjt1+92xDMH16V3RCfJlgqh
6Vib05CxtOlI9+rh4aoYgaXyr+qVCRhQNkRdvM+nXEuikQ3RjWXFEPH+srjE
mtKrSnI8me3DXWwEKcH5yBH07jvDu7DCXWZK3wnVz7Ore07IShqjUjnPnNJl
yrPnaKCWuhovYICLqAW6OYaK99e04ZZSZFtN+4jyIc3Bal6DOWSy6oWMARBK
+4Z6dAdYKPx2dZ9QbAac5QZ1KTCd46qMbC8A5N31+rGBNrHDzk4Qc9wecsJo
TtfSeysnmHmzpNdsRVQKrDtM0l+MCVH6hdESrlTgaGYJwCuU9QrgmEmU9RxY
j7fX9WZCAGUSUeHOgkCPgwUrJLkdg4y73GHLqdRkdJmKmbNYmSU5qRdW6Gk7
Px6wSc+G2mx7uebrynyBD9xFM4Qa8QVShso2Jq+il2jCOP3iddM7kChOl+7u
2WT6znzO/aCyPK0XF+B5o3xS8r7EyQdbbWxfd9l/chJCNW0jAQHOJSMt6vAH
89L3GVAd7/MmxGEALM/ETmuBG3JweeGWxgImrR2oBvx0OdqD8vdUqCtCgjVL
n6AtGLsKrt2nESX19cURCZAQt1XVG9fONg4J1T8YaozcnPF5qryVHh16Cbqw
3MRBLhFSgLQ1CPhEfvHkxY5XApbyh9bCbEshORv7YHuqOP1ZTbW6lut2AkxF
SQkB351ANQrHFIMCf542Sd3dDeMZGdHDUYCcH7E0ZJS5v3D+qUftau+suzCS
pVXxdmo3NhxTxpHsWBF2l74pVE1X0/AnWC9OvPazZ93E8NWUcwN7kVn8sous
T8qSJGyCXZt/r7V4LV9rUh2wnjHKDt3nkmLRxYjjyubo/3t/enGWKxQcHid7
W6ykKG3Tv4xkqfGV3+Q46oGcGj+0aXCZguU4dFI2Ny97OElRK8vOcVVlV4RY
2fTSo6lEMwrLNSi0Ap7NfyYSpQuzyA0nI+qpJ3foMKu0tFVQJzpzSnYMIyL8
+lH2NkkzrPSZ2huZbiPa+ERbEtMxZbPOiT7Cg9HfIg+GAPVr5zHOUyCvrZIa
6UrOTST8Ne0dZO+4gVC7atS6O07brkhg9kn5BVRDs74NBWmGVgrQmItWfnBV
jmPO3C/Hdv2/Si1wI+M1mc1XbqA2LQjTgYbP5hXPa4xgTMeyg0WLmjMYCh7D
/JCx4VHaojqU7ZkYTje5jf1hDD5MG4NANXUV9kMYx8S6KcGAqs6cUiV9bDx4
Y/WMqpYjGv8K2u2BC7peqRHg1xcItHGQOhTKpMw3XrmUO9wZRnZqRbc72meI
cNJpjBBbMnMTLmyXuFkt97SOcC69DDzcaMdiqWUA2XEbMUiGFK6+SS0TqSUf
qLAp7EyQCJE9sztVYLs9qWeF/Vwd3DtPMgx/vExhXuJfutlkp0uDKocpYa/C
JWWv1Zqqnnnt2yZX2YU2eFnxJNIR4fVrjm6ZJBfUwjvDXrVKeqQRT8HLmORS
Caqox/MXMRfcKWlpUHTlblUurS5cAhrNk4CBSEoDAR688tDQhIHM7X5YMM0b
9SY5D6I4RvLsOcyswWX8X5sEaNSsarifnGGEtctOJc+CpVTMqk8fvhswotZM
2wfaB0O0+SdnNwss8mA9ODIrtUEroGtcd/fkz4AWHhAahD7iPpfI/irshYnK
yj72cy1sD4QtdOOFQnMBYRJ2jAF+Bx+zwdHZ8gyolq18D6e7U2Xx4l0qy361
Ou0dhKHuVl+VCG3G9XUJH6YttOiQdVg5RyMGOsny9YQkdIAuINCm12bS4VJT
iOC7Zp5nOPxsj5gP+9GJ1k4LusjG2xxpSdqd9c2gPOl/ZBl2YL7RWhdjbf/8
OLVIn8Eics4QkNAOYjzavIRGZg0Qqso904Q9Q6ByC1qXU2fQm6UQEX0oE54x
ZkUjBdGTr16AkRtba4WgZzo3Tz8jJcgIS6nDfZcAY5izLmGmuvw1qO32Rg0b
UFryGrBO+80ah6F9FtS1eIs/psq105RXEHjF+WxL4U1DI+96HwVfI3Xn/sJx
FC1uq5aRwUfzQ0ANZ1//0lAusGWUURQRquZLyUWRWTzzptWgkuAUagzi5Jtr
X1ywFMvK9HkLFLAdYswVbRHkqhX+/T7vMTv33otnsJdkz5doTGvFcHYXQMxe
dP7gSaRk8tCRsxW4Gh96yGawth9S77gj8NYTrCIkbsyeM+2WU5SnmRllQolF
TY0IqTdaBp3i4bnMJlKu/anxKWOsINARsRNV+ACeKH1ej/cD+nha/49u0PuU
5cxHIbbsnyH7qi9ACOfNfJFsiCnHjsihnEKZkteXRAYWYYEpmEFxPEVKjcH5
NEqWuwtrL3ROpcsFS48AXNSgLoXsqg3f/X/1El19UbOaAWC/h59n2B6ts6h6
U3rFX89Rlr+a2KSk8T1X0Tdoxdde8tJ+nhR+TXYrMvQgTwYrzgRAoa/PrNZp
jkTeeiphGRPZ1VYXHIhm0j1V8aaf3EmSUkyFPtmpBrsjmGJHSP64z7fkzszx
r8b06C7h8vBAQKTgc02CJ9baqRapgHqRsbpa2wpcExSg8yh/m3FALlWxHF5v
Dspl/+YXFvhdhM9pp/RHsVYrqjuGDmen2q14KKhLsPYhFYisLryO2ZfJrjn2
9N1kyKifCGCqF5OkiYf4Zlg18uvszVTkO/8TTpnmSVFPOiSCY6xHzzCmAJqa
scR+8xeGTYKSwR54muZsnn3aWZ5MN0SIjYEA/EDVx6W3SDCD+5JZOipMEatX
1ZuMiwZZP2WW+R3bAOLnETlAjmbr263yvyEfRmWx59uOSRc5LeEYP1lIgF33
cruvO+9lkMBtA0OyekDf1mqpWeyErTNge9KkWCyFwMaAUv1bZtQVCdL7FDp5
FDmUhgeThGIKjeAdCRnbvcL2nSxANwdfgFKVLIttWvO6SDPinK7lFe+fiB5K
xCT0NvOkIbDu4hetvKB9rwU/ogdY/2XgTnKILjRtpCE54yaIA0FYUKIWqU33
VreA/zZcuUtWvV+oBElln6/306o41DvPlyth57ERJFM4WF8Siv0gFKlj8zhX
fhBlcKokZvuZjvaJB9VZk8FA9rCK/dvSD2+fF/SwDLbGRzycYAcBN6z2/hzv
/+FibK7CdGciHb2Gft15fxh7H84zBu2dLjXtegutKX3gBvV0ggWltx0ql1YD
k62C6WcsuQOVDAGdU81RxyOwXNTnmm4jeE2r5+0+IX9K9deSPmpX72Yd2wsE
er1hdH7aLPVjZJGas8Qm1k/2QnupgF/gO+uowieDhulldBOZSDmrAjn/0t1V
euPTKjvkM5TH/iLbxPQJiae+8Y2wDY6JZbABD4lAXZm86Xcdf37p1AH2gUxW
EX3l7gD0nJoaRwf3Kqj4ahj+VvaBtgWyI4SZeR958XUzzzrtSYVQvRN+hEty
7SQzrOZFqj+xL0ei0ftmRFNuZwXRdXWhk2AdYX6LYJginEcn5+K293073Snl
rqP9omNSoDcntoHZ0sFRNVHghw86qb4yvgfNKn7w/rFnT0rsFMln+AFgtBpX
Th1he9huIUGkyNOsfv5GsWqode22xs91Ao03enWRx+V7QEZOJQXTvPjN+35X
rCIRfb4Zv14GA/+WoYlPwUoNBTkZsP2C0qDz+LnCLw6sKCMGZF5M0hNgPy7+
QRzjxUZIIMfBeWeCn4Qaf5VOpFtLHZSm0LP1TmaNakKWHfW3emxlKDztIjH4
zMN37S+O36BCPavNY+mOlia12tnK7ixvHnzhLzygXxUTlqGw0aultUMfgpRE
/JTY7vxLjCJEA2v3NaGMLny0kRlOxn6ffEU+mAnysLLzkAOvzlc4dqBopir8
yDmvUFSGuyG/ttEdWNXneO7MyEzVHGqkQ3igLrSqi+XRhbvSzPUqyFr1/5rD
L5SPn6/15STLHVnHH35b2qUclPQlJnhfgzcrHf4ULYI8K7FJ9zFXfnhCVVaD
A0eP9jxCTEA2NSN+FAZ7C02D3uA0qKFeuHB9XOQtPrhw20rSoMApRDx43GLx
HkN8Re5FnD+k59e8U0ATa7o8MmSv1zug77B1+ZUjoI2a/vGuLcgqgHUQ8SjJ
uveGHX9EwHrOCJV8TcaQJi6iiATxEF39gC1+0R9l/Pwi3inSvo1f7BK2ESnk
GWbwWq91ZEtJCilDqa4LA9y/ran1CIWZi8RYkWCqxNaK7clWWTXI2wlTp5V6
EBTW8G4U4DSpQozRdi+1q/FFf+S2grBbdwkyAhU40R77uDrEj45CbtVeRy8P
bCczMzEua90dG8hrPHCS4ULpZgpWIfv8k92hywJlkQuLRsv5uqmU5DfZFQbX
HfZfKsWPcX3GYtPUG+Jl+vCD+mdy5xS2rAxGHR2kcK6jrxqQkfR43OP5orUH
W81q0N+H8Y8y9lib/PIQ6Ca0/IKKgUFUjBzOOXVzFZUerYDx1YXVD9Kl3xmb
EscXARrCPCKNw5e1kas5dVz9MXCroq5ToNHCjqxreVuSAa2OcRpOzSa6TsQ3
20wrumhiNCAuYkvDNAVQBW1Ikeqjnjx5TYlVhruVWqpbnlFPjn0bb+O+z7Sx
DxnWdXdHCnVaD2GMWGI2DPCMTTESGvwnksU0uAvobQ/SadXIj7bXLVLclj45
/8X8HuOAnMt2EIYdk/tTHa5LsZDZ1PWaK11NxmPIKrxlX0IhI1cm7+/hf1vh
ZPfs9omJ23UBvnTG5TW9k0KL4RRGBbaTatdRYw7OR+dSEyvDduaNEK+RJzGN
ZcEEY1d3TlAicMbTjGu8+AUGafpEk05QTP7GhWeE96GYE4VSWm+7BWkhQv3A
uePDPhr21cix9p8pnYetXi/WxQPWr86gbU0UqWO4j++5pVetLw6SXclkgtCU
ep9SiZvCMC85oyC9amoOLBGh1LpcQUUSB/MDdvNSHowaoMUMqFDcgtORW8qY
40DxTSI8KbRuIjNiGRKBYUe+p9TfzbgnS9qogTX6aGISVdXEwB0idpDcw8bq
CO8gvxbpHmTsbMDVc9T6cqSMHZi/RY/sojOgYFOOY8Xio+pK6ax4wIoOzcxu
IV8q7EumZwWfu5RHCR0/hwhB0/8+Yxx62HtCEelq/6hgOgzqjxgeeFbbd1SB
WyOtBFHf7kBPNdWA8o4Xg/bpIxZjlyO9Ryqy/x6ScGdFLNPudUkxFoMgASqj
zuvwHZ/KzkmbQ0Umx+67sN1oUn5rwyhG9fGM7YFOb18WeHW046PqEnzwFIOT
JyGHBNzHo+PHf0xO561Es8riho6WiQNobxnlWCCjxzb/J2HUCAt365vg43v2
Im+XTjQoaj4h1Jdh4kNdi497+4/614hJbkzqjmDXlXi1+2u4w3WK/k/VS2Rg
ZA8g5DXBP8AUSRqhVNuQu/j2IcnIeJPrF+dy2lEUZppaK0WQVo27tX70x/I1
XnpshxCvhw108ltuuTkeSA9AtSx836cx0TFIypLdpqsFOn7QE1O5mINyodMC
c7XR4CGVKnbQAFBw/e4vrsY3sT0FHr6yMtie9qUQXnAIAybfgvmaPrrElCvb
qKe3Y7nc5yIcVXyKWXYBOc4eu43g+LrVQb3UUCtJtuDHpMtxt6MwyeVBvIiH
lTzPdmACm+BPIBQHwr31chGTVPZsMV3hSVGVVyrRw7GAgIBcTilPg9mcKS9q
tb/yHPSfF7k6w/YpY7QZhKEotHskdDt7NP8SpEVsMtn5KFt4ShsHsEruhlsu
q2WiEfNosT8Gdy73oav5Pr4wZUqoiTU5/UnJj162o+k9IyrsFlOgJZwI3gIY
g0wPmK9EJqjMzxYS+BJMsw0cBZF2b76GHepqrSwbGftv2tZcVxahx9Nvj5xk
X1nB7rFCJqttFXJmsq+k1EIc7BgHwG2uEYMpdA8kKcl4bqxEt4CIIonY6kep
aGwfFv2ROKDjWxhXdWHC9xU3HyKLsYu7mnPJvhRn8G4nDhWV3bXN+XEfl/D6
lOtrnQMs3a1hg7h0INwBatE7U3AXpqqC8B8rMwwxTmr3aqP4Wkvm/KCP9HO9
bseHUvdIk9RSyn49Z7I4gq7O6WvKPeeFDyLnLd81VuvK7ko/PNIqOQxeVjW8
zDE/Jz0NolQMSD6oxpXcUFoh2xwvqM7qbC8zbc0FGGEeic4oxEBw4ZDUjKNd
FWExZi12QY1DhJ/cyBimo2BkKlq9iJhhCeR3YTnu+orIK2Gi3VFa+G/9YQz5
gE7Y88+LtdmV4HWCHPFcj/V/BNw4hXGpgs5Qt/C1VuNPm11Cw3Src9JueGtS
1/PmqoRlf4gY1FpUA3qtWGjV+vEZcfB5N5w11AsNokPbDIRNw3W6TJn9wma+
mtZPH4Pqdi4TEelKb2Prs24XR4t8iROrFWF8ac3lydUVi6bXH+gJLNWRwQIW
rBkFPMGIP922HqP4FVVcEgj1y1qO3dp3qfk9Wb2Gr7HpvfhRg4fqUr/YHqfK
+p7gggFUxt32BaQYZtApXxKnJpBiOyZL8xPz7L0QiI0XAdJeansIq524YEC3
0uaoXL1J+ANy4wFPn8DuYZgf4n/jHSDaqK9EfqE5tHjghIVs0nhzZQHkeIwk
xGKVnHeJvgBU671N8ENxrcfmyxYmY8HEWLswlB1g/7wY+l/SSrGmftIxF+2R
vBfV5M1oyJI2g6VibtnFMcWJ6hj6XYXIvYct18hPR7LGg24C5E7ReCcWsLRE
EPvf7sgXsA/c4k4d6ibf/Iqu7vwPqt3WaMAQYPavlKzL8Mevs7Z7JmRS4fAl
BFsaJT/YFvkX2Z/hhN8YOMeYVxjTGlhfHYP7+5FE+guOzdnAuJ2VXfgxl2J5
MzP+5m840UZTMoBUEbUw6N4RunsnuYhBYtNQ/OGEfDEENuGIcmOYYakdqRk7
f1f7eG1T4iaScSwUl+v/fiU1WpnFiJBZqUMTZobBfYgyv7Pmrv9DxO2+hBiz
KSGQP2ElQS5Femr/Ars0FOvG5TtNCaaEmCbt1ewnKcBuTjJqpCDa+YVSe9kJ
NQHOtpc9KRL/X+LSUCEVqPne8UG94HWlF6HN+8uD1hjGOyn7jYrhUnYkXO6l
nbipLcEgXyfxKHPS8Z2c0aPhG8fv/CIrZYpOoh46sROQ0xKGmM0AOICbpf+5
2NrK8o01NODm1fgEuI5cihH/XypK7NLrlAfw1m71FcE97sGJyv7Je3m2UNVg
bmAY3fqCLRNVCyWFpi2+C9Rm9C4qUmlH9+ZUvSh3i4AG7O0GYgpAG2BdMkcB
S+6YnTcGab/mRP1UmftYvdbWG/rd2AUq9Ix5n2bYykhDWidnGD5hfxFPY4WU
8IyA0vW7Nsxk65tSAlzj4sEJlg3ny1GjzAFCBXx462qwVLWrwBH4VMezt/Lg
nr2yM+L1KQ/BiONmklLs89iYO/gJx9OcORhNB9sQC004tpQwxaszAOKouHT/
dlR3mHBW3JMU+b2hQft36lt3PxT0eMOHhYGDBrh5cSbHDA3YkBn5MOkKYjwk
Jy1cib+BoNw60wJTHcbkjxGd/7VKGS+cPSeUXytac/OEzqmYr9d+Q3XC6613
CbgkaBQ7OozuaKoWzELCqyKAE8vfGKRTi804fP4xj4vN8+7BKewLLzEOVBoD
hGFDHhhEadJlHpHl2Fe1hh3uAnisoUnTvcfffS1dMSh2SGZVH0D9CDZf5LpU
Mq9M1nsws7XQKK2TOfyL/y/wT9/dsH1FM6r0y1GdRGZXUbM5aWP0k5olmZBK
ukjSFuTC8l0rvtBNGahnDhlz45Dv/1avCH43OVycH6xSCqLMHGXBzdft7Ttl
ph2bsbtYPILAK3mtF/G76W0XLcW7pbHSf0CRkmI4m1ClWejjTJz1DwWcQYhj
ttxcyuB7pqYLVgD1UoR2LTRPl/2Ien9rQRMOfcrSBh912mDcGXv0Pomtey7L
ela0io2Mx3y1W2VzsjHbpwZMYS6AU5NbA+jc5Ajk0mdCGOAERuuhLYza0wgu
NXxRreC3M3x+SnR+lGwyh0SOiGp+4YxHlmZRimUXgHU/aUkSTPU8bFzHpO+R
aelypyvJx1RpxkHCw3C4XilEWqGAgUFs6BrzpJAGRBFohxHuEEmwE+yFwaeN
ZnCUFNxEWqlrdpb6ssz9qSs69RulHYXtoIgCb+BovU92Gterak1gtIcW3ZF2
qr5cHg7m3EdTNRq/fQza8MN6aB1gpy/zV/CEiWRgA/2hY3uczl0Ac/GeM2lJ
tEq0kR3P1sElALpLhKyJlW9HQs//fCqDp0N4CkzOiyVBLC9/v4WL0g/Af2hr
2aeiD3VeHlyl14BDAI3VdoeU5c+6ypnHGlpLDXnk4duhTIgIq4b+DqYfLHaa
io2eqbJuSpX+YrDa8Se2u6dagHkYBkUzmaErNiMOqYQ54NuozSDiiOvJ7oH9
BebL/zStpTT45JTEQSm1EqlFrTuEDjQrNMrTXuc0jaYYEwQs/z2uO3LpApGZ
v6TGcQKcnG4y5eT5KucR3jnqG7qau+jnqhm2iFQE9ug72VkXGrc1IzL87PN2
Fx6SSY7EgYxNzDj4HMyj8QofDbkEfc07cyujXDAQ5QFgWMmExtaEgcX1Q1mT
xj2RmGX4ibB5ljpVMaA4rF1mu+kGFPyceLuD6p8HKUo5QiVfcVSoUWjNP66x
n8aoR9JLo2IAo03O7XVeEO+O4foZlZZ4MKwbWBSkvpXT++yFXjjdG5yWaWxZ
8TGK53S+Yc+t8fdsD79A3k2k2tNFRvgI1AmO7HQVlNFvi4AdQMjFkrLj81zC
ytrhB3SF6j1vWdlFzwvAKXjcJpXpwH18WIt5TqkmgtKpc0OLxvuk374bKPsZ
TJGRyLiYqxMD0FziE1ycY4TL7N+apSlfALgkIYGskGCRtG6lQsfbfi8OX6KX
ipiG3ljyCJPV8b+4erg56O/d+2hBJdnuw5qMMMn59i2juxm+wmq0rIcInjhP
WlN+DfuDyv+emYa3VwidrdDqsz5yBzmAj5mbmFPQLnswaIuIRPo3yfpdxVwF
SGqOI2rSW+zx3Hp89PGJV/8hhwSp5E86i/MQPZDcnDsm/d5oMvNbvS51TXD0
2LizFj+K5ZY9HFA84PBE/Uh/66mr73NOymki0wLY50Eb9/eGhOgZdqTVfnDs
dFp0e1Q1CDL3IJh3e/3+tV/c5r4m3Kl8nbOhPG4xnU6hIOqGSApoXJ18AJW5
sC34GwG2FLDXbWaW7Cr+nN7vm+zphXs4CFS3iAqYzlmB/0BBqIJlxmCT0tAh
NayU/K+C1cBGnHmpGbMGhvwf5b4jwdFsSQgh054XZCfurzDxecjunKJrSoLN
/efS+GnU+gcVqRhb7bAexOkzvXRLy+eC3x1I5tjln6R+vBKPKT/UkARkp8Rg
47aQWgKXjyk3fuigV/moBZPP7x0UQGREkvtszl16BTn14RX7oUWMo9EQZGhN
LTjlKDS32nqRqOtCX5x8kQVoPlBtVomg0TaF/Pe/J77Pif1+cy7FBFTOhzff
XXofvqxvVMTLFUunJ+2ATn2S2F7bgyMDZQQp1AhFoLn7/thF/Zk5rih1dTTB
SFnvJJfmDoN3U+GLF6j1s3oaFgXpQHyiqSdZjQvqUNzJIGRioq0FSvPEzRqY
dkYcFP9Iq0jCw6jMTfL1oK1rMJTT5SA7m/2i5jjJpUx1KXhR+kOKLhb7KUAh
uePDneDHvDoVM4YMk0yJN2XqvG1A1tf1YU7kMIbLymAtaBoFqMNmgzwQnG9o
3AzYetIoiwx3s3RR/PBUyE+8Oo4LLsVaVN177UoUx51XMCSYkeXMvNLRFUcM
1oroYYfLQZQjuLHs5LAzdrkrMBBsjkYLTnZb4couTRJrV5eJ3DvTAplI2zxb
X6D226AlJIx3XGWia9bsqcLbpecVar0uX/jKk5ZmNwrm67/VvRMQZ4cnntpY
cdh8Eb1a4OyAKgAn7hWyjJ3NaZ6iwMmBs35I0Kss8v9JNPzCrX2ey8wXj1Ut
CHYb3pOd1WRmm5yuciJltO1FystG5R3S0qMZnq1fxC3tYH7XBlMqeszySIK+
JnRkung+WKtv3w79+yuDtwhFpGIZ+QiPvukzWV1Ql+FD7jS7GWEVMzVRaFtL
XU7nKTp3+kJEPLDUcvOcFgOG/3EiAnboGolJIkfmeArxBTZd48KpkNCuk2GY
iKVz68nnevbHTf0c/tkMsUdVnPdQXmHsrIvamN6EUNqKVM6BdMdPdQEEdkR0
RO53AqdpoIjTuuHuAmV54C5T42kggO0nixvEHPyy4R5GCGoLRz/qp4U28rem
JY6MAHLL4Tw2JDAfh6zL1StzQC6wcDBF3v2wwuz96HhUcciuBcWgDI0am0LQ
q3VFvcppu//3pV2LCGYOa9BAG6ZEh3qG5uFBsznswsFuzDxcXeptPnob7ZBf
n669p1UVbVXWnZCfNusTPQ0cdKQmELWZt3yt+HIAkGGvAmIsXN2xG3rD5/Ey
Um7Uv7Mj8sz4NzczMRwBjIfnKOPUQ6qjenokT/rjri44YHR2dVNhNxY22Ci3
SIqtkAVBtAvwBETD320X8385YCIF5wRW9l20BmiPTFjwQr4Lg1sJvWL2FaxN
BylzuBnRqsB8NO9PDgsjcYzfNAbS2mpgKK7jPQGCV4/5cEn8CYeuSdhhq1ml
etglv6q4tF5jBhML67cxtwUOeUyK8RbPW1C+RxWZAYfR+ptJBJm5zWWKgWEI
05vwNAOHNIJuQLAy/2G67WnYlQXQPs1hRxNeAeP6vb0hQT49lRS0lyEAdrbw
kacRDvw7tQSwVxyZIKt0WQG0CDjmvGAuRlC23/UolzpN31ghNcDDJoMRuoDV
v35WC4BS6e/8MsGOf7BI9jsr/Wbkw9DFVdVJkaI05Bi1YIc5/FYMXv6aUzWS
TZZ9SObHjjtZ0jkauqrdVyh3brar9Hw9RKzFlmAtTgNL9ePMeJfXzH/oPxwE
8CGsPWyJvYgteIzASu8woCk7kboX3dKq0x4sk7egkoVHcQHNjTR+C+cXW9vK
N3MzQ90lrfnGQQSGYiQ131vnfwy33UKTc/xLCOAZGSA9jYvtHw8XOe7HYWsm
JROBaUXtPZhaLFtCNpvss1hsfrH0eYD7kMMiFWBKMfZg4WS0JAA34ZbqXw6v
LfD0gu0P9UgygQtaIGrTXil4L/SxE7EYcDxzkiuA6ZG4fxESCtXPtSHf/5NS
17bIWUh+J4AJDule0t8DqKOg+untwsfrTky0lmV9hEIqFgQmGYF2/V+hDGbW
3lDM5Rq94jUyf1s8+lTSpnPRmMmLQgBdmSuEGJ0hM7orVxNoaXLDRInNNZyB
+vNUvJMqAwZ698uFE3MzrpDgf38S/IV4v8KK9ixt+c4hlszwCe5pn6gbvApb
kP7o3jzyoLuLiURfctp/Iv6jS79FSB+8Jrid69QU1eDN60ppxYR/tlAa/4qv
6XkHP23dIZfGQWwLNx4QuV4sWvHnvPYGPve4a7RlCH/iw6KqUqA9XTqffese
CjzsUwMbX3GKtocdnA1ZQaEDalMrcHPUw+dRh07Ccp9HcQR0g03zTXmzW6Db
TdR1cdsp5Sz1T8j8aMhS9bsf3jwGygJXsmWyBeML6AMRrkI1HxugGxpoTp43
Ga1K6hmWXcDLdFVLfPDDCS0ml9qNmHNOs4PjHpPLaOBwKdBXWEf/S0gQRqsR
ul6lSIWyWYVqYytOqeoSnWERURFWo/QqeIni2ogbl//6fA81WfN0JjNkZk6U
W0DXBa7u7UUJOcHm9F8E5mNyhGcblzCEprhg8AIGDBK2Vk0p4CEAzaZ8z5eU
OIi9FxWgQqY8ThRquDk2CZ7pPb4TJ4lkoIHzr2DBASV/NmUnR0FQTo3s9COl
Ct9P2QwpvKxu8wUSq/HznLJiINuL3K1xKXWosugHe31BayIpB40XpgmXYnRY
K83evS4p7wrNnNxsWPH4TdeNGOP5Ja7gS5A9TdshMElI4V3oNr0+Y/iBSX+b
IIPRA8lwtbVjWTmB+sko4VboX1zdv0YhfViWGcOIEHSvgFwsYRa8gVkuL1/F
5H9AzcYpxsgH630UOg923vGkBJ+Uf89O6mK+tT5tOv1tT11TotyZuJN1vs05
zrjVoAoyifd1IUwJFpUca0pdq5y6Y2JDokPfWgKG574skkt8MmHfaoONJ7ZC
tF7BC/g7fuT3v/ThQtXozcLIvuU5V/cGnFVASVCMBvk4yqmA+R8P7R4ChQl6
tMOqkNtyv2BuUzDLDpgfSgXwPBld3Ny0XK4Xo8++RulKxoNAArPVf23ZiC12
kmyQAYCCtmhut1klAFVbsx7vQ1CRZk01EAFhAtLG9zaP6FLo3ed2AAtkWVQ9
vwtm1sn3rAI1Da+Co/yLbG8qYzN8tlhRZxgssDve60AxrW/jaEe9UgVG+Zze
xzXgavEuqEy33cZ8AtKad9E/CvKN4qj8h+5IwjGydKQmiLLJKGE5tYB2NpfT
HLxQfQdG3saNew3Ii8Tw2F2NbXyo4zUo8ujrUo2hEW/28eO+MgIQNtVR7rku
RGDd7BserS3ErzOmT//9DRij/szhQHZbD/XA/UOsPA8j/laPHOEKLpnIbXjT
ZmCvJcOzTOyqRUFOE+MtZ6IqiXAFPYA6V3ajjeQAo12pyiWxpsWdWBZar/jX
XrqSGha0KsZpwQBXgEvlXtWrwwZ1Y1V37ChoT8eVQSeWL8Yif1Nk4JP/uBBu
am/VpZGtPnPM8BdYeKc3Z/S6oX9eZ9+sy5xLE8+1ONAcekZbA/CaK8kkA4Ds
cgbgKbQhXMhQgSTQoC2//vAJhwzmyFt5jZXGKd848fW9PZmkoXh2Kzs7Tblh
3Q7SPkWKWD63HTjeCBHiZU2s3Dvd80qZLDbKpXCyy0DEVHDjBCBrD430YLAC
RaLSC93RfDHbsLvum2RjiYz9LUqaCLihVEWZyWcUYJ10WLRxMxgSqegeGRry
kk+4k4089CdtH/Wq74pSPKjksWMKY4zEEr/MPfcBgqAEOzY4IV7Lx7QehYia
iqBjaV2v2ORvcfuvkYvyUXXzVE/CKqvWn2bIBoDCnANuqZOZ7mK3f1EXFWpX
+9xeY9J67SQTLGhx/B2mZhE6PH4SRFbGEqod1h3SutJvIv+3d33cg3G3eBai
qD+TqncCy3r3pSt8yIPthXRXA6XE8Csi9NS0tOk1A4BGDPPLktoiyv9edGpG
GHDk0Pya223SKQw9GkMqP4hf/xEDDMiA4rys0vwwjGfahx08iwPeT7HJ4+0Y
m+Tn2sqjJ9/uSBJ0YgM7irjzXLvEQ1qSJkXB/WksdthtZ/mvdvi+5Jr0mFb5
1lm0P45SQevET8ikYzELWDG64G1YCnOf2Qgvccc2ML/q3TySjf3YqtYp6RtV
GXzP/0fQadnWKfTEsPoqTDxIxln9qAf7PmxXLWOsMfV1tlAAHy1974S6OFaA
Q9A3iyN0tfuLr4KCvJfxXHtiSRqHcnAAX2SDz2ZZI1t87K4+GPUSxdHS07ls
kA6Wt2I9mbH/1FhsNmzLXYbrJfdT7vVqbiogLkDNdPoHO3aXeLKzAzS1MQkW
2z69kDXlzJFWxIRTwMkNc/3RKxQAQ5n+QS+YRWVmOykTFZY1eGae9Ut6WTWQ
L0c1DamDTj/eV5lt3LXzlFXdeq1wygro0wv5jkfzGAGoJP3O2CGJFMWcQ8BH
H5fciqgPgkJVWxhYmTa1JXxMqMdQ1AeWr+G2ayiOkbDdBVtAux910FZRBgEF
oH1Tg8eSaLyR5IMfZ6r3qc9Rds5S5T+gScBMi8H61MunyvbqPpbeD3wDDDch
F+HOYWKwbhOV+umZrW+Evagt8ROnBn7KteARaDVbufgqdpbsSarcX6sN/wWQ
CfsftMBXGF/1aiVx6hLBimLVFp6MgKkvJ9q9XI/iQ6W6vcCNO+2fTS2bL1Sp
om8RZ5BSnAEPdNIrdmrTwo3gLCDypeN3R76Kr9mfvnzXJMLr38f6qzI3SP5O
qpBz4ptDtKlygR2f2/FP8A8zrqF9tekPKHDxON9sBbDumFPRJmiXK+SQQ+n/
mX8U+qt45OE9bkD9Z63ce6WJKZR0gBlHAF6v54TwVl9zJ6KdLnBRqnvN65Rn
5LSYwwVIUuJABZdUsbW+gIN3NR+D8oq9r9OQZEyJkIC7YA/BcTEwx7ohZgCI
suTPvL97Ikhxfxm7Op2oRwuFa4jFtJTWrvTIETFmaAJRYdRpsWaBLTzT6eT6
BV0T4MmE0l0CGdN4D/w/F5G/fgAzddSshxjxs/tK+Qelh/0QQI+pmEnPrVvP
yF/wwsveWo1cm8auGqWRfQgfPWGu/PrYAFzBEzeX2glcc7EunimAOYOy2mn8
VXkZC1A1aOMdV/wANviYJZ4pY1EZHWnyzXbMp+px3aFLGfvCPddd3KuFtcCo
qgLzCvPq2SNANVcUboOwjZAEDnLKrYcQBpn4Lb3kqjbR5p3pZEyhgvbpJ3ue
4mIijziajSf1DtMakbkorqycxoVX2MzBTjL8S7fHzDMkdNeuwnOrfAJ6oajt
Cfjzzv29Nr/Q6bkcV9EI9qm4OyMM019bwu7J7k4XHRrNd0g5wgJYhAdmRVRs
jFtYWB5bcIKUhEduo7d6ZjJYQDStHWQu1JH8FouR3/3KINe7s72K7mxioHbh
2VyRM+4lqUzyryGQEJytb+VWgeJjF9iuVvwzp+NBp49w1h/GoCoqQIYa5b8K
hrJJhuyEpmFhb/d8vv6Erup35JNAZhtUXplEA3eTMFRfwIjBGnwJGkBRoITJ
o142Fo++3i/TjlAqxrQRL4agNCNFxLU9U65JprIkosOCRmH0WcCzqDLduk4E
h1FsnunKH9YYzaPXqYKr2tLAmeIIVKADqmRXQvZUlBsV4fd8m4vYhRD++UpN
UePv/N48gArnW48jz3+aGCBwn7DbYSJQCs1bVtBcmg1FOry8fcQL+6pbTj5o
EUVMeaCD6yXTZHttdX+i+ifk68/fYalDUaPmX8vjlAXZoTlR5AifGBtGn+kH
IRrRhQrP71REJfB9YHpWihjykdW56Z8Ue0pMMcax/Gxv/9PIlZ2m64D6fDsa
1VtlO3VYjBIXmRnwGMcLaLl6+bauTcXzmNWV8rintVid13TlFnyqG23tq5QQ
9gG3JUnaQArsIw4QCjducoTBBz6GAutps/wHzh5hL10q+nlzMB5o6Vt1c4l3
A82gWmATOWmunVSfkUlWIqFnVxqW7rBM3t+hKg3twCe7fBVDTod+IPlM18+l
5ryKc5MrtV5cLRTl5cikOAYw3dhWB5NLY2ATJn8CoLrF8NcPafxHWuHABUdP
H2Zz3UJLrbY08UGlik0x7OBefEK4NK58G2DXKIvUsWLTDNGhY2EIbiH6omFK
nvJxZNBEPz3FQrlkGwxFgYERPHcCZgbSbgMa9i2l8ADH7qCtCjd73dBjG5pd
ODKHt+Uc9HqM4OeLLPoHTyvHr8zs+u3BBh8cju4KGJEBeZuL6C4Fg4B4L2eF
Gms6WRnHcVqrvb1ZGgXP2piNCbnffgDluLQaGJpyc8bGmrIJKiNcCp8JlX9g
wgVTuTZlSOLwiUAG1JVbu8yDiVDucs8uG05AN2tXGMufs8BMqFWQqcgJwQ2q
Pufwv9duH4t2nfedkuVs7eWVn6BtjKR9I9JjhuBeqXNTntsn0tK/dxlJ/Gst
jrU9tpbEKif/PmzhvI6YW6tPTJF7gzGw9Z7Tapy/tzpD1N2jLjrZtNbzk1WS
LhacNRAq37Ux3fxHCRAlbNcx633oJjmCn+bdTvqe/xvgIVRSZL7wiBbvFww/
hoatVh5uO6d+UtgvRfvgnr10NdtFJc4QCaZcTCHtsxFDIY2Y+gPaq39HcLYb
8rMi3D2uHG2Kho6laLRdy4h0oatnbGZOJWewLXGxwB2veOVCLqizOM9GXMRh
3A2zTn2gMYTaiz1nSOC2LfaZckd5/CQLMJ82DE88Xl7zBX1+hdNHhcB4NrPB
ncdIe45L98tX7IeWk0tB/XzAC3+QUa9tqdt2RthG7cP1xDSCirbXnlPaMR7G
pi2PEoWtjpmNaVUHgL0sPRpHwBMdsZQrIzhtwD6ZmNU8DUSyl53ioxY5uUPm
tqD+moOtU8s5dVOOnm36PX4FVsm6OEuFSdkiaWpfhnSYIyEQUjJcMKe6IWM4
yXm3w3JsGxoBZgfxE0DAzihesOawosd2ChVBztUYTmqL8iIijkzZwHGYcFFB
yNiAezODIMaAj7GrYPgBFTlgLdWmTZ6+N0Ktc22xV3eOXuFAwkNt7K3Ndz+l
LWtxcdZQAPc6pQ4RY9xbJI9AE+H0Wfz4/RrHm5gHEtjXZJl35tv8MDixztZ5
10EHGIJuzlQiY1TgUt3s0yIEv67GE+R+VCsD2dN6oNEZDgK6tjwBQqFfT1z+
cfaZrG7rh/S40r+kUHdV4+7RFaMI4Lz72tsYbO6q4Y8zECvGX4TicYzls+vR
d8ksDp21Q3bx97ZubO/269Kzpd6/PwcAvO/s0cLs7QOiCnLyJVFqd+tZuzBh
D2sG8qQVUpBRIGlth5wp49GJLWzfaPOLKlA247YWAl8Kit/bKuQ4aQk7Id3s
ydnmrsiKyp2gHe5fQ09BqXnXmqc+JVYUJKP0xVa77i5nuQIKU0jPHmPUrjJK
3gZrVQnmr/NkkO+iK9KV66XVIYev7w2mFo4uapcQj5LbPcxW/R/a4iHuVjhH
5bDTBeOwkHG06h4uQyPZAz3AHhgjYWBQ0T5oJci+1JRjQThUyRLk8jOmgITd
ygGfTfBG3FR0p0xrpc8I9zZMDhjnseGRcuSwXsgAEo3oqTkrQHf3HCyfg+k5
xuD2+ZV3BCfxKRhbOZu20VrEDVr7SXGAPXFjeaSly+T4zkXY4zEkyOv5esTh
wdkVIPoqs51wNXz5HoHFbqLvvXpMgrCQdjD3A8bD0XMrUXNIxglbw0izeX+L
Fyt2g5X9sZ+F10JozuK+SWPcI0RjHPt+iaBo3ec4Q2aCqKw160KUhgDrzqYv
TRscppb6TeeR+rgtSttiao958sExJPsNXDDPbZE0nMRXlWDxngsRWVAp+ZOb
lseloZm/vUlO7EY5ad0E1/+um7emCNj1/fgWSUuGPL8JuolgoR5+0RkFBsjF
wvbk6ZDzAmtLtq3XaNeGBj9NqrGzOflc/1cZ+uNG4dcbc57FYw+C15KVlRtY
8ouC53gdjnmFzkmMa63nirzRpWg2c0bNsdq4COhCfq1b58uSvzZQoRRTdDH8
zONDYG9eNvOjTyzlPN/sMCYtxDsG0vkbXlLJ7j0fAe6uolKRrMONFCsHbmAc
wwZB369IXn5a79MArF/T0ajyoB7ULnX5yYsLppa+hwExyDkj9FBgE+TbSQ/L
MO43VoZw9B5sa+LYmv7DP1AYXXsgd17JpjgqCp790WYH9pA4LHgClN8Cr3Pt
RWrt7YFL3WbtA7fjZi6NWjirt3++ljtc0wDvUTb6Vfz/+TZVah/xGPNnS+km
x3y/S50SMLkoWrjakAoJVRDyk2KrWXhTKb56lXAxfb/zWKnNG9R+d+/j/XqK
3le6Wq1lIwZ4ojb0b0zN+vZqHjSwx6b0YKEID5p1N/zaOFniFmGcGr4jjYdX
eltdkkE7FCU4VuxP5tS0bV1YCQTVDyg43NZk1B3DXSX6MiU3p2/bhGqcUSeo
fDNsgzLacMUdgkhzQLOK+JJv2YU8UjYBQ6K/1or29p+S5BhFLyHXi3yE5svR
j8Ilh1toX6JCkiW0UiqttmKhaMt4KnTj4r8MOvqEMsxcDT+zrEpS8Xmr3yNI
mpbjXb0uy0/7XELwPw2y8dtZjg3V3hgTQzdP57nYSDjKlLZyMWY5Qdc30r1+
DOLE4wqVpCboLsLA8vYDRMVPcjAYPkXmN+WwW+9DEp/WmWzXratgMeFAbjyb
ZmIMCQec5UubkrP7u1Q6OqhpYyHPCQU0f1xIwxlsmhzFBTq7ey4pQ8Qq6Pr+
lVqWdR3lah0/DsyNGzqw/+yAKVzC71dNAoVOzdDsxg3ADcNzCPTismte3EjN
fn2kC9nfsUKJH/QUGl5TGkX9QKiX8c2YsQf4u67M8q93cmR5WsczqkTEeel8
E8ve2kIknhtt6e9NhQgrlOFEkHZS0nGXwCyci1Ww1RS791Mw5CMbWE+pggmk
fJz+EiDhMOi/0DZ/HNwgACqTIIVgjPOlr5C55ubA1zgu/Ufhx54DjdaTSrPD
q7cZ5boIW7cnuY6W64GPc5bwfckcfHDft1d4WIkSvi43KqNTrVuNBsV/7678
W7RZHtKbNdvF6HPOYAqoC04o4fB9MrabggmMt5RrzS3ZLG2pwBjB9wJVn/5i
s0jJsIN3ZXy1bATXziGuMTw5ANNzMuJV2zUZKG7Yn5etlLecRMsaFsrpL/NS
/V/sUBY1j5CB5ec3goiEjOsVXhxxUZPXTDAjBATNhs3C8HXQ7cUjnXBs7nY7
yD63glvCvV0s8TIE+Rj+PpKPHRA0GZx8t2C97MsRCA5PrvL5sHAT36a6PEve
IQle4DMPkqD6yifRFTpOteXs1WCe+wVQYLNsNBQDGZaCmXKL4ODAT62YtnHC
r25/8lHKYNn/bM0Tf1itpfdVpocs00BnhL1rVqoW3NJAPLk0BJ5xfvaPmYD2
GLdaBt+YU28L9msBxpyr1cNjfS8+WT6lqe8kg317/iro9UnbtJk2GDGeAdY4
VyQ6NmHO+/ypW8oIfJV8U53T/rWctFqgYW7RKhxLVK0ruW0lR17dq8QyC13i
8at6RTzM5I4lSYarn5uCIJCOM3xDxdJIDxNIigbmhxuO8BaYSL4AM7Y5rXwr
FDxv4+pDWv86iOiEFRkuUBnPcZzaYrpm8qcjIz7SCP72iE1cJjURQW10KEyd
nJV+DMDI9u0EjP7g1o/urXAsu0IzlgL1+kIonNqNT6BYD4/t7KYgHBnwviUf
Sm5eo644DVM40BrgL36GNoOxLrfG4iKWWPwva67aZrt/9eTzLsvDDaHV4/wz
e7Yqhjd1Kpyvh2sQgF8ImEaLTJUuCE2wXWcikfrtDpBHTdIlNa/XtCpnKqR6
swOOFfATAoN5VVQJneiGF5tTBwz0/AsHZBbWBOGOyAJBXauQCv6gFn01VSbz
A01H6U294f5livHAPIQsRJQyBBTPo/x590UGl3k/uoXIwk2IcwxKt5VItGuI
b20eQuF7BvyMdGpJmUkuSYmiiY2lXUEYuIEeYGobDNTUxWWwS99VYkcNlyQn
CgGZJV6OLf1g/bNrmaCaBme66Ah241xK9/g5/541+PiFM2WUaPxM26rvk9gE
zDGvYQXo16FQAX+qx5jHPJpXtO852gvZkFlpiSYb1pB85ulPOgjk/mmOGJwm
mf4qqwoibYNINbN8BZbeIsv7IrpnjmJb6eaxlb68bwtrKVoLv8QmvDITE3K8
IViZRSD3uVbZi+glImo3Naupqwu8Hhq5EydxzsHAKGF2xOApkc0155mo+RBs
6INwNSxxlj36S5Jp+mFnWFeX0WJd5OgmKuQiOxTlnnkoNRdGvjjHbBVDcAq/
VnvoXAMZyhHGOh9lJw9xepvXBhq/3GlST99OceTtlrwJxQPbBU5cdGQtssOB
vkzQM0utlbzAARgPmgOB+5fjUToB/YppYajNf7osoLnXgDB4bYUZ2HmSddJv
PB8to6QxuRLwG/xbZu6rO2eTmlenFcDKZfqHSoClP/DgWRYk1kLn0U8S7+IC
Tgs3EToc70vn63gkRET0XmQ2kdM0KICDFlk0dfx7T8yuzWr91i1CD2Is2z96
p22zxOE7ecByQTDyHWX7+TEFc/yI644u8Xo+dhVhad08Aqgpn1lYEzbtcyO2
aCvBa2tXg26jr32T4+5LqYFQnkqpfMtpmOzN0rMdnJIBQKzYCETiMrH97K2d
TzP8cS5cLEHAqDyBd54sSOqbwztiWAX5/SNnvz5WF/CoHKVlYBmiQ41RGo2w
tLhr+1JIXlxOUk4bT7gvw0gYs4Ng8tRhqABVmSIkt0FTq2CNO7MH6V8dHQuR
hjuZDE1iVVuwuZK4pE1VIzYAAYh41ktgWIZKuZZ+70PYwLh3karFt7/TkUzH
kFLkAU+e+kkwg2Yg0l1Xj02yl4W4/2nlsLyM63Rt269IRmY1GZ97srwzvY7q
mKZNcqVnKaeJwz8liRfeJiD27CgTUkZZONTiGlWy8/AGUHtESK/NSwZggja2
/6qhIbc84BVOHtQTlSGtB80gHGxM4FSjzh7GmMsO1CmsTi5dovVKNmONJUfI
cw1ZlUUBCoqCqqtC1G/3pu0FpmmZ8wJs7qIGkp+XvCU/tmDcNR1GXhDXkxRs
Vg3UAquJYhDrkTBY+X01EKTOrkb7Gm+ZSYanZ/bzrTQLJ9FtZtcENuKEOBkE
egsXYksU+S2ujLaosY2uqRZmbk3ZCCT/aIU0zDfzmnrv6altiPP291+sWfY0
6/HyPhPTc+LDp9Z+zcrEzWDziQE5UKgI/X5m20RlRwnxBEz85vz8g3Uj5at8
c22cEp1gDJf0VSGV3bUvUXMn7JV5LeHQ7htCM+JXu59l5xhe9DXbS7mI2SlO
98JYmbjCRLwe4ZPCDz6J969H8CIhMRup9Y2NYbqDI6WwseGSKkBjETd+kqyp
uGlO649wsskZiNvv0GiatfFYLIS2YVYivPV5luLMdmX/O2Zw1XjrP6vhsUqR
kGuXiZ+Js+a5ERTr5x9HGBmeCcE8dVTquaqT70VCocVZ4Tsj29svA/gZyncF
U2Wl7Bb+S3hAa5ApBWV60v5BVGte4vVTZ/zGONhNxVVJSZSbU6ZprF2KM6dR
Il62mvd69GidTgEPBiAWPdr5MjHwAGmg/UTlb4ADue3YkboZDlVPFWxrt35K
ai6WxM7iwUNWahCwyPK2iYxAguZdplrYo9m/1eND0ge0lp2uCyZ137g4HnYA
sM1ypzV8kJHmI+0MYS+A7BJVi2kbhnqAECCkMFPFPa2eiVcXLQCT/CtzfYDK
RnUrjaLLyv4CXLrwSRhsvZSlO9x0rKoH0I7p0iMJ+upeJf+nguvdof6I6oxG
k2d7zFKcOs8Jz+/ov7sFpVXxa4aYHy5Ip2fvVCk4Ccl7vonH8UKIKi9hs+kQ
UT3O5aa6x4BZ7+b5Enj7NSFCzdHeBJZxh+42jTDSDxy8U1y9pvlHeWstsQme
3+jHEFE92nDOoraJx68uXz+rdb/EbMx6H1uXDyMFpSToE8cRqxyQGRkA0khD
JSW5SFbKexpMfv1J9rRIiAWJHlKtomdgr5oRIOLDTD4McAeg+wT8/lq4cguQ
tZuoID9X1MPvvMM4HzG6BcpsjRyn8lJuztyvfGcaNKXqzYgeFc2wSbZ5xsPc
Zs90qiCZ/7RjAlF07YFBPxhS7X4X446D78lsh39sw1WTsmmPt8Sw0ILzQFjz
gAWkO0SwM4d1nTij5f+ly6xGD8Fl9uyaxEOpuZ5zLzFjvZskEaErGILH23qn
17uhN8Wfrlkk59pSjhYXcV7x2HBqosCYp/xq8gKN6P6HZTqxbbvSoNoDDrwO
xIEoGCZUlHrw0q2yny5CiRieKuY4SdXzxF7ZPFNzt638fQT/oV9lLjeByL67
t22lhDX93xWCpxO6Wec+K4o4aHRSLOQn2hg1wHmuaXmTXYCi9rMN+XBVm9qo
Fb09Cg8pF+YW9NTnfJGmgooYgeE+SXhAzt4wxwREnQdf3tDpgkHuCfpL2qDE
FtKVxPqawLVx3Wc6AJwV4AqfMPZyar8B99S4XndgVV0T3bpBjUDZYp/1vXa9
cHOFO6AsbjtaEiyViLhSO53T0G7iv/k8j0Clt/4e5w1Wqe5HMDDIAt18QtR7
vb80zAgyJnsG/mGcbNYt1OE1vEQYqvuB/cqAf7+FuiNIs7RLmb3KGdixDYWf
06rDr5ZLbAirz7kEANQCX5ENcawuCQrFtEP+EueqV11ISA+QEXYwPyZTDfYb
4NC9EtJqMFBrsxPXxgc4ej/F63ZN/1oZ0nPaiHaGBtPuEDwbk6mU0OeqURlk
yGg7Kc2Q9m9i4vCn7LHIrZyXm9fPre0NclH9kz/Bl4iavabUSACgz5VYV7e2
WJylYnod7PLGgtJyDSTREqGQQCf0G3xBFrHs55a/JMghKjcuZvR5l+gE1CbP
Xk2awQ7SNLrMQLjujhDpeqB22/vUK7ur6NsGna598Rh2qyYsVAm0s6E1lZJs
nGg30AGdnEy3OQs7b3UaD0twSysAaujsqodNokHr0/5CAbM48gbSuvxPk4vO
5anj8GfFlC7u++o89bR9mW/cSdmTqGSs7OU68cjNoCzeRe0cV0ubTE6uZ+tX
b0Fm4qD2wFDJWZsxfBLSAADFSMvfKGQLRDbhB7Zf6JRt7OOMgsUjLXGPBs+H
hH0ebQc0oiXskZMm/oehw58n4GBJa91mTy3wRYdmeFZLopKsN+DBC3Vdtco+
efIKGIiVcdbCv0wfuvgXtrkPgehYKo2Yrl+GmOavxmKg0DERfnkn4Nxuo6gv
tvuF7HsrM8BNNSHAfqrkLbkeBxI/CitURvZcONmiVH7kR7v6LcotzFffG8Hk
Z6R8Zjg7McSSuzEK/Ftp4TOGAtAkQFG3xlWQl0PgQznEC5YvpkR1nQVy7uRg
ZtaSMColnLbuk8KYqMGs0I6liJro/AwE84hHkBteU6DvlMOQ06PzSL7CDVmE
INQuySfuElcMp5pdqWcXD6joC9ruX2r4VWqg49au4IxjOo54lXkgmDBqSpW6
vdvAMMQX0puTOPHwlm5BZFxLEIXXsN6PWhLfU1CezTXdm+0IfVG8QN/AfDAO
o9fqitZ1eF8qf410+po16Vwo2/tJ76pXlNY2k5NRglbWwhcsfigICcElGm4T
titXAZ8JzNi43afdG5n3J320weP8ePKveG7W43mHsOorEikNnQwRd+JZHSxz
A+NlS/HJrKV1jms0Vh4piauwz+d3H9jFdw6COTXmnuYFmCTXorRioT7q4Y46
KOyZlc0zDj7JJ/1fdDGMqt5i2iJVj8FrNc4Bfb9iEDQSKTHlsZFx8GsfFopq
hhth6y8LzNaM9BEUtMKPOXyJqpI5gY6n3kVFA8+FPqjmC+pNyqlNhSWyItS6
UEqo8c4CVoJWWfeijHbkzMcaCX5TGx1ADV1QcEx9QKrnsg5ecgNfQ0U4uYAi
0R9/edYYNEUPzWv4oQaMhLikXp+aF0OAzw/zpYvh9brw23+UteqTzyGAhvd2
gBrDswlw0KIweIMlbKAOB/oxKPA5iUYmI+kbJVPAiSccPZiHDE6cx7SE6eAJ
EBS+A8ZcGvQcC6bTCSyoffpsOpeUmOjViiPCDfJpFArVvAft0J4x7KqrINTe
ek2KcBGZG6FrWjEzbNJ10wQNB3mM5SXFUmoxPYclnT90QWUIu6qBrHJQVyC2
/jrCWRFw5S/3PpL3KrYfHd/NY4wibdNRqZsEi+sJJBvTyIn0Dm4R1KbeTvb5
JXoBxsPsVFduM+lokdNpNGxOzfF6xXmBxXNtfdjNxWPDsnTtTfBUqQ9Zr5ul
vCQcUBn8iE8oOW0isG6oVeQBCNVf+lREFADJyY2tPq9HM1Tint11jrLv3YY+
byuaeG7wc/x6/MQxJHLEFFzVuv8bdevKnOyzO8IHd7YbfT9MHUGaQsKlpzlR
SpLn+KkvoM0+3OrJjHXQ4pJTei5LOV9IYNNFJ98ihKGq5sy1x0ur0EwS3zby
hESHI55V+9l2+QEyhxMzrIZpYgdJCqOFrl54ZBVahTp0F2EyP7GbXP4mk65n
XtlYziZ/sZ3OhMzkUXPr04tUtDVXfGvGduPBiRFdzrIVQx1AlbHHjUKnX//E
ZMTLewKTiAqIs4lGQx79PJ72AegLHB5UtNnRm2p2cD6gwmEoIRP6mm9MSKaZ
c5ArEPdEbhYotQjt75xWxMs3XAN7uPQOdDy1XNjlVoqUQcMNlb3/N2pZaMn9
8OElMheOdecXs+H4KvWR3hUbgPnkGZDaSMxcz1LAolXDxlytkoR8pdohR/WJ
pzZl0SlehTWUlW9yTUvMoWW0qmDz0bl/qUNFxrTdB/8oXQUqB16+DMsAtO4q
lIXeTKaKVPgGtH2Fg3uGiXQiItRGr41soELDrzOhuLj+7vmk/X30MlC65DT5
SYMgORC+S/fIYM6rvancvriBkfzrYVkSEXfpQRN7EGTISK0w5ThbTyoQE70v
+X1Aa6qluBJ2n5ZkdUCZQvPbV6qNhC+VDCUgsM5uhY6bJnA3kDcthbOFdVYL
EQNV4Ab2c83ZLAkbWQk8JzmDes3aOS3HySKHzhMcG/BjI2xgjnvfGAX23cUY
S0L97yEf3i1wuG4sNC6+kv+LOWG+zL/iIRXAGyVuygQ6lNFfnBRt6hLY5u/4
J5TMz12l8KyrzwZiUQueIMLxT5zEUMkWAKSO7A0AYMkhjYspZFNnrD1c0J20
PvWBI5KGhMKgjVNrO05izZyUIucxUgQQHyuO1UF17+MsSc1Kj/uNu1QjD0F3
JYAQU6uMW4Ua3HoZZgKWp/YHZUy22xnFSLIFGCYqdGIKWAKXYIzJO5N/O7B5
iPBRjFZDdZJ0gGnkvrJ1rE6vZHT65Ihu0DRUr7XVCJDd1J4b/BkYdUtpPDBK
HwZi7sVu8DvdxfVbKJX1Boy9wKcj6UjQFJudYC4ku9mJs2F+n1LFgNhgmM6p
Xb58RamuxMQ6I8rFsVBtrshbKwtbGiETvvr0DC82BHHnMV5/Ib2YCHOWq8Ea
m5k6XbC2usLvAhyOtegvEXQFn+QYhyawpSGP+d1m5sx8wKSDOcgZ9oAt3t2H
KjuF7wc8+no6BgUs+yGnHHG9YpidLg7JTwFgnCMaGMI8G6MfGpHLF1VXcWLc
8SkkGmuhD/YKg2HpMYeh2L1GMRXeQzlDMv1qsxoaMIxlLUlM695QUII/JshN
eM7gEKI2h2fokeWqkMS7wkwMqWGXbXEXWCZPCQpYama8I9kw8crW9nSym0kG
8k146rq/OrXmscJxcklucWmnXnIiRlXdTQZ0hnG7x7slHGagwl1QL8VivKes
ab4vRgdiW9vGdqtZ8L2TXS/0Qh3iL1QbZ4NQOQF4BDHhj0UBvRPaHYK/2FG2
F/WM5mNAwI/XaU4WJAeiR038QWDOV6DW6x6yd7j3NJFyXjTF9fz881sDk8tB
ansxHgt9DqJnuahZR4eLKSZa3OrRUvY8Fj6c7bpzNfzRU5O4hjO3ykOFsRwV
FLsLhZzZ306Mz6QDStXKcoXyl3TzuMR/OiCijQ8GrpEFN6wfUy3pH4WmYTCe
VgxRbweafoRJJP2Chxzwo7KSK1giDfQpaYsySmmFchA+O67FKlo8JzEcJVtm
x6RfETFf8Gk1Wa58Lh+WLmkFlGFiqnx1lIHHMsIMkBLRh2YvfpVoWtcO9pBC
FvL/a72i06XjpdZ5tU+fQmPZtJaenn4inr8badC6NRFUc2GLKS93u/QEVA94
ZJG9xJ4beu1ojOgwsG/QYhjJw/kqMtShOTwhTIb2IbCu0e4e0rd73heXpX8r
F6I4RlW6oI/0xD36gW/52YXU42uLQq1hHboyE8JKN4w8djYkO2p1oOx0gVTV
xMgA6AxVFA7uk83u3etLjAnxbbX/EK2MW7vioihrxb9MnW7dMUrgQCScQcfl
U6sAu34+rXzCa2Dc8i9Ylg3U2H2Owe+3CqvqbDPsEJoE62oVMgY8t2LD248T
sL/nSDMnjkg/eEVc/rH17aJucXCwvsaUu6HRDJO3oME6hwPijslAaQMRHXsU
PrpctwThqD/4vrJTEbB7zXBftRpg7tTOE4QJ9klsFzNMjVrpcwO1rN6hv/B8
XN5kWTvEB0xQpD7Cz9Om3j9v274DWw5feSjuh5LFY1cwtGSkj2Z5pudokChh
7BZrwbJe9ACTr76ep2c8I5sAHX9qeoMMEXL0LFN90t9nqmwg65bGyeBT3XE6
RXCu1mh7+hlOJ0Cq1fsy7yfzS1mLcuwAQyknXZP2Mkt+PkBBU0mQiDdiK/Qb
JofKlLbfN4WtQ2CDAlb4TaU4c8U4DQPs82N4yCyK/DGaNk4EyMA+SK24DF6L
JSu5SFzilXZ5KwbevWMwV/1NRU4R3t/NJ7GjUu8gnwwn3hAorLWkfD1pmdcW
mbo1biAVKSTTX+CN7RATmqNm2bAkA2QrMN4r8R7mUk3B8L8NiNGZ2+NuD3ma
PRLdDPk3FSjcpXs0ZUL9TzQHTTm7MToGW5Nq7LJKqR1oukKpNvUfKqpeLJUG
GtzzOdfxKoEOpjcLBirX/KpxwGDTmLVvtOEGs3vWRguC4cqv25LnldNSj1aH
RFsOv0HQkVOnAT2IcmXuxHxB1UHACs2d49pZUw1v2YZySwhg6Yo3xKhZYFtl
pYnLTWxX09O1STbn9VitSy+Gz9LBSU7TAzJyd3y1BXfw+k8mjMtqLdhu5Ky7
owTTrTt40B67fiGTEonpDbbIO0pVc5DkEbhC2LVygrgtYUxrnPLOO3EYbLTI
NFK6jwCdhd8/pmWEuGo+xv8i996sL/eWc7mcuapLRukMe0nEnIn7N7qzgk/w
NGourtkjjuio77iZ8luzZENezyKBwNkgpJGS7EI3V8Zy3BHNhBX20i5Z2TfZ
znF5ayxzQd1Q92lPkENKK+sTvsEU5DlEeFYLRGBFkXb56PK9KS5fW8gURJDX
iM/fH8qjHfWS1JzXR97Z4svWG7u9t/gc2gYpWBYwQWHRUKPdj9CgHXy08AWO
hOafBupoTaz9uCb9ZE69oj7lAoZMoer7J9spyr3uhC41YlRDUJb0LHgai+DN
L9LdG4WUGz9nzm65ClaCOLzHb9KwqcAKlFlETTEXXUSP+5EN0OpcX1lgLBrM
cEfk/FyUYR/dDEe3VXoer4N/fhyCUz+lRpCNMtvPTJ01207N6XtqKK/OL0a8
HW4qQhEza2ZwAhgnAMVOZbZTNSyEJgAK6xn+Z97OdHyRkSPuvG24vOtqS9w1
MDVivco2LGY2VkMUIYbXTH8n5xoUuVgB162qmyIITBMsVI8rEZDdv7GrfdeP
K9Tsb+FOglArP71jh423s4YYJq0giOL+7h3rjZr+pnyNavpATx5FrQk0IXHZ
ogee6ECXty7AECZZqvPuqtDOr31GOu9QvJhEY/2l+8UkE6MlpUxa2Y0WoaHW
+G7hDtDQNyjAaSU+yAJ+VModCnuEiVCE0ue4EOP7CMu4z2A3xebTf9s/OMuo
aM9nrkKmsPT4kTRXnKWfOerbZvWnmRdNE6+xvhfWmkhk7LA6uZmE/1LHO5+l
5DIKSQExScnxiQV1gfj9hTEbQqqWJZ5cqNFF/HeOCL3M7MqcVKzN60Sma53h
7CJbPNrfMe133DYxLf5xYNacFzK16E0Aul9L5DXK/4DApBemN7hx0YvpWu7j
DuomxqxpcVQQZcD2AA/Fdni3fhieVcgtfPhXGB0f/ieHmeRJHEFr78rz3SDW
SOViPuJ9RDy7sWQlOJ+MMfZE0TSoUzjngotgSVUr09AW1I21lgmXoAp1HJjJ
/ihwJicm27LLHTOAuFiVbKyy/NGelXVIv5sg9YbcNLjl1EWfbtjVp36jprUL
W51UR9hd1btK0YjrHiXpam6F9kdFOo1tKKMJ0ba6Mg3DBniOOO6EgmPOuJ2f
dNnjYsif90oqf88mlyueMKd6zuFsJzjIsrg9kfzEM+IcJwqaKy+nYBL9d9NK
gzXmG7VAXwNIHvonHF4MVI6v9eEkILCqtwjvT+ikLPLFMZMPE0jfV116jYf+
CYaC6XglMZVlR6nGz6aY2JqNSC13w1C4FGE+SxGj1zN0Ter3i6AKMYNu09Oj
M60OTJC3OKmkXwXNN9K0AlT0ioNFNgrm8v+qWvOMfVzGJQNYj6wIkemEPw7M
jKuFWPpS3NQj9+sgJQfckw8mhjKr0fBOq/DMvyS+dSQDSLiZfTw0gf9fyLOj
7dMULNEzxCb+wQwoak9/L9hbuNGaKH5Nac4egAQNffcqteI3wf/EfRpHfaH3
eZMd3E6hchIEQGU5Bk95Y9IBVF9wgwt3rVQ4vXTTzjk5tGtH/xTErt1Vc2hR
AdW/aA0yonsvCWfAYYKQjXEECpX1U7UOUCMW32iaK3qcq7/iMBeXKwI+ugWO
lPzx8hnYTpF5YpHcJ+E5BzzcxivEEuXw9Z35Orl1HFqn34ryBmlp49DJGTYz
TOIwyAaYZAyyxV9TSNs2wiBhfhtQpX4irs3meWjokuqwXqpB7COWnDvWDhhj
0FJYZIwZmVKWGYnJeSrdUYnoRfNEK12H44+lrH8lpijRx4eZUDY7cH0ldUJG
+bbrjzrOOHlqr7Y6A8U+fqVq+k7aOhp6XqNQiYwlBPbM2P1CdVI9fFFL0kwy
ejHMLJvEHGlJO2dEAmsWKqE+9Ai7c9a9vwYzCHJrSNkk9FIsSOAV3+JgPRPd
b7bBgQ74fR8Qjzos2kKONfcd4NE8GTeWTrRptelao7VkLU+r4XanIS15+D2v
v29uROduWoGvzXYu142jYGOlUYlbv3y42B3+/2su+PG/CfsiXqnbAMO/MhwL
297rpU55MzuMJQd3YHSqjkjAXwgBwAksUyYC20q4PbJamUkcIh9BOaEDo7cB
schGlH1y7yPMuPSwqrsnLf+6j2nQ9V5/H55WspCeII9QCSl/jw20kyCXRwmj
GTnXBwfy9y3GwIvtl9L6J+DfW/WcRzXgSPwakhZJCJrj0UK2yXYVxR/4BhMD
5vtpYW+/NwIj7LGIf/t9izif78/O9I1ow7nfuuLoLnzAvU9bGtGn6uNnAArE
cHpWxk/7lOM7hFEM3gyK58ToCb4iYsBJV+359YjW16qyvWzi5RZg9++peNBM
0eytpMBWigM1KuOn0vHmGKJDh0X4IPJqBfpvmXoQVrZM8bGd9jHPqZWODPFS
V2C0MJ5A3mKIgEuS1ct5642hBBf7p9Apsv3PuutUNt3dI0bB25axuG6QVQ7E
HV17BxqF6loomSaUzk7ZjW4u1klTW/2xkhlaMrw/LAeX331BtB37iIJPUHUK
jmkAy+AOALO/IAEIXTNoAHC/FySDNKv5PjV08LmAlsWNLvkvrOlSLZNNq3ZX
qOVqPKb+X6i5CiRPOCK4O5sbwEtFiOCbUfV/nec+x2ZAAm7ou/HJ+qgJZp/7
NHhL65vfFupQ4venCmVwVXV28pEpGDCLqu8mQgaeLh4ucnrQOtFcw34hqXB1
xTxskzv6jXJLq6HsWbmZN6AUUKvTqSPqOYuOU9U5j17BVNR44NimsGXj3mUY
Cys2qbXvf1fGr21xDHhUv4E6PPZjizHuW33RYYkxfiBOflP4yfvefPlae0J4
7TiEkfL8Pm4PH4h9FztXNA2symwdrhjeVK47k9SJeQhnvU2HfNibzs6Qk4Yy
A/lZ5piFJnqUgJU+k0aSTgP+Cnqf43/53g+wP0N7aL0fGTMjaG2xISHmj0f1
5mXkybmiRzysjPdXFufIdOSGpBfxY6I+MptHkhUNLLR7cS7zfN1lbTlhtMfd
FrYRhVN5axC4J5ZzI5z1T0KofvKLw3HxOeKal4VmuoJKVIkIwMQwKej8gSlK
LR2isVU3zw6MA0TvvN6qpAc1MjvddaFAycUUVWQ/n+aj8tPszuMZy1sUUieG
511oY2iZO9pfA6XxaEnNGSy7dYjov481j2lX+ycVdOOeJoWBSCny011Zjn91
did9wLdrNgHfFpfNWClv4E1MXFIyxjdZ9OMKX73UdYdSLkRwyDUHFJgwbGlR
G3LQk40xyOlTcvHP9GkJm5aV0icHKNL6QB6dko/+ECPvBR/Xu0YSRKjRgiGI
pLWC3gl5gIXq7wYWbNRDxE6GiTTDd78g0hgda55ArhzRe54lYEpV1AWxpkma
F31wEzlipXP8qcpPOW/AaFvQN+9R3ynfWHZymHWv91duoq0aDUox4dplp3Z4
7qUPOUFum3bJ2CZQUgwFL/kuDg303c2ApGctQK/d4Vh2KcsNHeJDDDXgAooW
NQVdku5eQfW5CPMRghRH2yUtDXL8uwmIrj1ceknVfYgj8duM1H5pbQC4sNBJ
3iVI+Jqb282Pd/sXuCvRxmEMkOQ/C1kkRYGMRLJZeskOhoMBbFevDJZLVxJa
T+9hi9Cp4shb5yIp+CIvlGbTSuYqG72hQ993nWP/Yd4pKnUZrVHzAIpUh6i/
hptR/dWsV5HNntCsNTvc1Cp9L2urYUlXFbZC5daCtaaoaesrRMeDuIqgZbwS
nHenCjZ/y/Y7j+I7VtGRCbAySQGiLL+ZCvjicI8tScZCcUJlWDSMEPmkqlWL
D8/jCj6fjBupaug9y2R81ZPtMTvfhBqH6wGbkBNqtH8/zTWOflmg80AImpSk
nuDtrR7ZxfxfFCZvwwxixjqJX5a1LavMyXeEdspOZF11mSBf/TJOFZiYDaAQ
0J+1JOsJRVrjFMjUZsfmBBlyOQYLPNB3dLsT9tJE3GAa1+tAZ9ET3g0y98MI
5fwVjbiUKnaP8ZCF0upX7n37h21e4AESeUn2nR1z4dZ3wugl3Mj8ufBRfD2j
sUO537NVwT9tIFAr25e9EZ50eC7IGXw5iRe4nTUxJwrbFQSRxz2PpJZADkmb
3Qm6iXxxgODb4P8oLq+jmiYeQPfIeRzVCQ3qcaUHqn2J+HajgQeoHXsrCbGa
8A9HFX6hI7/YHhq0osi/dY8MBzxGXqrk5oBnKBqGTRb4L7Ji0EPkFobPWpBp
KqyK55eKzQpPLOpe/P5jE+M+O9M68wKdXj3/bQADLE55eE6HQUvtVCglrytQ
Ec2gI2Y1fpOslgBiXzDsWvSavpFeZ35c7+KlU2B7iQjH7Y8dORMw6w3k3apq
xVKlNBnhFHFPySJE0hmLn3BQPfbJcElwIZKsJLbx02sCZYAIyk6ZMeQ7AoEU
PgK9FfiHFyFesduvDRPha0JZxZ/gSO8ENgJMq8GY8nogGpiYxk7gMzcpi5Rm
LpOrDyXmvdMzd8C93pv4BQ7OP9EmxXIG9ibiKOfIygnmaxblVy3BXcAZicWI
dTI9j0k5JqGpmdgbDjzRnnSGcCWv5cCXY6WOjohmTjNeEmDr6sxJFEkfN+hS
euwUC45mq5xQg5fnIGNdDRwBhV2hC1Hq0u2nbCcfUVE2LwrUp90ybqxikIpQ
n/ceEY0paHPPvk2bLY34bI5HDwtbGq9mwlBmjkRYjWLx2zQlt9fLgZ85cmGT
DqCuDX4zV/OWit3w6NdmJNLzqNwCn1Ng7nji0dPmhMSzH+6dch+bjgRjvK8L
6Ytu0zwcAWLB+q2xfqS6Ox5325CUwLlabtXP8tvoUwjJzvWlTBsHW9uY8B0T
UXv+tAln49Y4Yloy4HQ+Y04SfIdz95aN0pulmnShkvmDe+s/N6+WsolTl9fV
38GKi8Y3OdwP9TDS8pZ3Szf1tj4/aG4fTiOkc0IFW8aazoHXyL0dDeJZGXXk
3vUB8rN7uk7/fkJGkc5fZbPU5RNxq+9zHzthl3VPXZtU2CNbxnAoVzLJ07Wu
SBs0ujXKxVDdLCd8OXokyTzdEWVcpKkPUooLdeYJIpfFHNfiEP7D+Sj7ECNL
AI+uKGTvsvvDbnH5Av9r+kEwdBuhPMl2ZA05HYDD/nLsoIGw63wkizZ6u6KU
8049NZgaiws4IagWhtTklMQnMwLfVi7dwbf6ADboXQRVRoL8BZhfsQY2Mu68
wU/HyonF3fY378mBJsoFcgBREOdBOGtGgux9OKp7qJ51FLfnsiKkg+FPrlvg
75culZN4/YSIslclnevQ6BXk+dmsWyr6frAAQmD2SvwIyP8Qjl/vl7aUetwv
AIEKea8o1Z9Kryamz4MsFkB17mhX0KAppEYsMztRgGZ+HVlZti1zjP0W221S
6Z4AK4zkah+1DucVVtNTqq1WFWpXhBXAQJXm0LUZI4NWM8cvLir+Fzce0TeM
kth4/9HZswYRWOHR46xtnS1lPYTQnadWqyayqYpxwQKdK9W3AYXYdVk+WLc/
gAxmTDkQQsUCHgTXhy6AfZsIWrhH2UzlyKxDz2bYr+w5Z752WJ7m7U5gquR1
BBoMLCQidMB7QJgY2YFUePVDYIzpZ2qYSCtyMWqJ3RVHKDKnM0frPmKw0nbV
t+xM2eI85u4v5gllsFd62VGi5rUA7PSu6fDSE6UsPprJubohECU0nA5OqVnN
eAI7lHRrKt3htclOf9isfb79u7W+gXKX2WRn6Fr6bj0CSJSEj8Ll0U5oYDRE
KovIWrOIWMzbT1ll29WMeJT+vq7t9rJSp4XblvrYrH6BVYDBh8CaOWc9gPPS
G1RIDidEPj3bFxF4dclhs91Z4WLl6nmaPCFiSG2ZzM9a5J3FZSdeMLstAyYI
+Retw1e2UM2OYbG/EE7L+/S8G+6r3gjjstWNTKy2u4rThi6kHe0ik0ZlA8xg
3GbgOJ964OoZmmetlK4YVP9CoIfMWyN/LhNA1gFiNd3PrzmWMxoJzrrlN0EF
fzKhITFT/h9xX0ANIYq7HhQe9YQPH9FmG/R/55FEIyFX2yAg0vlaPkGCV/Or
lmPrGqHKXIfmCIS/eNkuJ3k8GKeuq8gR9Oh443mi6vprD50GcEFZrpIElPRC
Qo4rOPuLKB+mXkn6Mqi1Gd/h0izrvNybEqvSAEQN4qB4xmO9DAr1Ovq4McaJ
x5SpQEvcNHwmIZp/JbiX1tKyFCaiMCqzgNfxG5SQXKl6ZLHrGouFMh6Gm8dN
tvNIpu9zypSD1g5izUKMDGypMcAYHeA695MYs+w1WtLx1AGwXnkhyRkRqj+k
2vnsFwB9StQFc62tyWFpv8ICPLRxHE+8oQu3bhSQgPzLo6VToPohjjHNYPzn
U6FQOX0h2YnZvYbGfuJ6muKx26Rw9K2GjzFGwhhE+TQ2WnqveG35Ljk9IXUZ
MGzzcvK9D03F65TFh8sSi23duxboX47YGF5EP2aFboistQ6WzjA7nMDwJgZz
0XbMVDs5UQigfOwZ2r4hr3H3EU7ORjWC7qCMltxBAgiOy+f0G6l6M/Yy+6DK
Y6q3rM6pNDht4gcX5fXmGbk9FK+judV67QE+atNHl5nvSPvwXgCB/+nuDXYb
0UtuqFOVMYuLNNc/dgilxtIfVNblwv098/b3Crc4dOc/KecsBhHoo2QYWnIf
Iz+b14DSKpSrWUpvbwF4Zc6MPi7fULpfk7q7vemFWt0kzmc863TH5lyI1z3a
/cdJbsvi0fGi0Cy9rRxu9EFPAZxq1jAhiwUdOLdrj/zlZ+6qOiUL8Ehts1xe
RuQoRvN+ML3p9SaAy6NKL1bqex+8M8zcVtsumoER6boyEaUfHIyMEZ/+cfyd
Q+TY4b8nTBHKeX7ipy1YM8koLM8MSO5Hm+6H/XNatEq+BVdnKx5znFROLtyL
SWLvjEcBO0O7JpkvbiKrMF3yuMkuxdeD3WkbwGLUNje/93SBwZ5ul1pC6rJF
kUaOlveYz5EV/7oGziukGUhcykhqGile3e0EI/T9lJf4S/C9LJyhNExhUWc1
brGhH+5+M/9v4UCH8OLIW8BDwhuZioEHvO7eRirHLMsK9Gl8nGhL0cnr12dk
CTxxbfpKah657xvw0XnN59SIlfPDye1jxQb2ug5NImBYfW3BB6A0l4/Totzt
SBDeLpFS+Vw45XQr32IEQQCEWjbUmLDP/L04YzylwkZia3jjLuZdjrcPHQuJ
8grS1dDIvlK0RnDQkU5M/8eskU7ysGFWpBiMaAoGdjRIDgZewql9kEtca9c/
3Bf7os948EymT0R9RGDsPamJyzF0eIq6noxmO9i3NRIEB2uMnzP8gIdYhdWw
XwBdDMtZX3mxypAd+KwLIamykfSAW8ZlXhhcozj8yy2HH0Wc0t79V5b/63EI
p4++8DCeaY9oTmH3tKm5MSUeCU/ZItsnPcPqncjXxXTP5C1SdCKOgZCHhoLb
bdj+sFHg/ZLLeA3mMTZ02RYnC6hoHeyWQFqjoIGQVuxn9BiMnJBZuo25kMMt
LcoxYHdF4UHsHjzaLw2MOeCRY6g4pi2pIWWPfCvW67z+8CfGQptu9snM2j9p
aNF7SzpG/HD9w0LmJZIpQBfyU00xUStgD4SBihTdOoz5qsou7467TK03sZTS
YHvm8lEjDg/EAtM+CtZGKHw3e4uDhmjuYru/hoPvSwV6/gHizZlDGvaNeLIN
MGe1l12uZwmpwPbZXLr7k+KcZqqtX5/7g87CkaOUfGs/d/xrvs98uxo2zJ5c
h69V8MeqOZs++MbWnwrnorWQtVwNTj5vZMLbW0NLpyHpZ6HaS0VX/XYzYXb0
0IZN/p1etKqXwAyEHWQXoDpp+h4ZIAfWK5J7bREC40BanD+QCc9NmRMHoRjq
SgUDIWHXyQXFavjaACMOfEC8gKiGVUdiuZM83g5c9pSPHI4kNYNQvDup5PnK
R6rxRxS4lifvPd0/b6PVU7Wvjtxqb/Pih67obJ/qAzrBZA7pWa2/YPm48VVx
tCSyvqaUECVXOFo0H9cGN3htEwnJYYqHZYod6NGGunWRuHaxbUa/P1o4/ZSu
oN6O/4AZyQuzWv/LSHtBBjYa50ezEhHPoIY7tYb/PbkkrKn4K9eQYroSEra2
y3CpucF3+XA4Z7kVIhF2v44oxDnZcABO0i+bAh27Ebplm8DizLYIMXLM6Cgv
gQCBXWx9rmPYEVgdXOut+T1GRfSnTp/UB+FfdZo9tlyaBBKz++cFLbAG+ZcM
rekpaZNrc+im3IxlLjdr5+UVVcDCqgk96T4aV2kmRfpAPTfU040hFswO3tNg
WEbu8arRnhTsdfQ/GXKOQhknPYSB9tc58G9gwYdBC1T0iJXEten+HN6lm8jk
vE+LcLsPmJEfJNgzj8fiW55mJQ0v68nxh77dSvlqRbSkjqTcYz9odi0mmaNb
mZzP9e6GgJ5zHp4lj4FLwT+S8dDMZ/0k5KMTfa+qYzNi8LXz+6n50WHAxLX6
P1KuRDNB6K4lYb7U/57KyMXe0ToN/XygmlVHYHZTVR/Nl0cfg6tFfyHGhhlp
sET23LcFu6WRY30sOqr3nX4ZBhr2o11smDh5FUO/KgFej6Fij3tLjo4hVAPM
aGY6+GPo+tact9OxMtVCDWHMyrML/VLY+TqQcv61oWxVc54Lwgp7iBDZllDJ
Epc7rb9vkTfAdUeZwCL9P0aYQRr8GaZ3WFscotrpXOR/aGmcWre9XqS9wl7d
pvlDA3U4dJefMeOXNqAH20E9REWSDtrBYoBU+DK2r+t3hWp7Vuv/7q0Iz/Iv
XNlHse9NG2OY/VoTAA3WjxtKLwj0UZzbJoD45Fq+TUg0nNiusj+4q5V5Un2t
KxrCMFHGolW5gzfoFy7XEptYgo+3fs4fLws2wr06eDVodMSBnH7DFVfghhCu
15YPInN2JIF8/qFBRhilpPcLC7wAonPgP2eEHgxYOXe46tiSdY5l5PwYw61u
yAqXjDLiFvEo3s/2v0k9/ywu63StLRGEoT2ZbducT2d05Eu3u4c+vgbQ++8J
junAimi7jb9HWQ1DMWnY6TN6Acmy7ZmzV75J/SvrKbOJoBg+pGtcOS/OV7Bc
53X5gOARRG/W6TiFK+sgDrtcRYdeJ+Xdbx1HijFyDqDy8r9c7Kq5LIwl8197
5TQgItC99EeCa5OZ4luL8BOp4mnsiXFDjn0jlew9JQ1so/XNe/4uI5xGvUHa
zs8jiRyL4NmW7bkEpvqkTjbP1Pulg8KJwN6/m9Jc4+4OSNJyhoTYTaDtq9gg
UoIii5tQVf1mj4Ubm42GJTpNp1p74zoa4WrEq64pM4s7L6cbwtRmRQWWEEVL
XDjQuI0+oSrAyYb3SCr66DqLRbNkQooqYCgtFbKyHS5BTN6yuJ50g2ey2TFB
6YJvDtSbZFSpzZeWgIG89rjbcZXCom+xRR7+7Afcx8jtl8GsnpgaIyZRtWZz
PWCEfGnu59wf5ZQaeJG1rAqDHBjJ0eCrsgFiHalTtlFyeIucemSvF9x0rmdH
lnjUCg4seA7lm+0B034Z6FWg+kyjmZjSFY4yg8n7oPsKfJgDS+K23UXCUzLz
QcxAI761M1db30Um4Wzkoi5PrTsP19AOlvhYeu8ulUkTM/iaVA2oldMPZ5bS
+j8I5Bs++n9bJIUPPwHIEtNBwHV/7U8UamLCKGrbRy10ZtwTaAJ1N5f8ANOa
G9xv/q4PT7Fr+lNFKTtnXWkxmn/iWwlSe0ol4ygTgpho4itLuqXKOvIbIO05
EQn6O6WOmMGYe00jqGeMVFg7s0hHOOC1LHdtnZHPJ434wBYTJ1jbxJFKmWdA
EVvGQnibWErCHR+Hu9oOvmoPIUneFhYIeQ2vr0CKQI9HtMUCEnB9OabTzxib
mZv0e0CQaQUhT/W8//xnTHbd1530J1SI6dueqHX2olDTPIsOZ4wMZerjdxr1
1KAAhLuuNyYmJ4ue//DG4BDY7lZpST7+0YsoD9xp8GnIxg6cBud2ECN4itAX
kx+EY31RCbITt/LjYlIOSLHXBKaWJpsi3AwPW2zFFyhvFZ9NmBXFpNBXjYro
LyF36jFAJWmAIeDM1iuPv5eq7x30mHLqvrxWLKIrpOu1Q3rVp/RpZOJOQzbg
8/wlF2IXVTHxXE27/ngrdZix2M2NeALqdt2jYpEI5bLwZ+fs4Zv49hrGZx38
IIEaOnz/z1u6Esqm/EB3TllS8nKZ7dLk42O+HgRU8+6O4XDPDKtHQe+OIW8+
gdOSo8fHat4VDrt35Np4WSmIcyWBp62SWeI8bAVTidizerY93RAwjZdPo5z2
EYi9n3s1vnWLynEuf2vr1HbKnPeqUSv1bGP/loj3xMnXTtWEHzCxnp8LF+LX
kRGxiGeREl6J08JJCuCohCeBOIeiR/1vRyt6MtNxdCtLrVXFWsJlfoouGLLB
iwfwMdf863WuoeWc8xE6/in3i/LOBkhIMbxsj0kf252e3GAlhpzlqe4+pDsl
fVb8L0lQZXxTK+9N9ivmpXve76rKKKw6TB3ICH8FvuA9i1/cKcKEHBmPjKXY
RNssf0sonPEDubUv3yiFIwPsHci5MPIuXCYN71pY8UYhmeRCkqKui9eMVAsq
x6rhf+Fj2duXGD2sCo9obBASOq1spIEiBi1RSuPmjJFQZVtm+CSmuhO+2bB/
LDlmrRh9rNtbYAyjnpwxUvZEFCxvey5ctu9r2rFNJTqcHXm+4JuhbJ6MO01L
gdT0eYoeJZJ7amJ22CXlnL1R5fuUxn9ydcHkrsh1UoKl/nmAdTeQ4fgkWIl+
tvA/Z1ZKO8DeH+TR2IsOM8UyyIPeNdYpDHrPG9hI4YdjVGwbt4ZGRk1zQHyB
aqEvBVv6dOfEwIwMlu7C/dJ+1MGnJFJlPFNqqx77Se4xLDRY6jQl0Rf3Khz7
OQW70GMot+d/YDjKA/dV+RlAMW4HCMIUs3mBHluXFzomLS1Cz6dO8dYKdPmS
Vvs2SNjn3px5fZ5SrjF8lip/kurcGgFxaz3V0gdBafQ82WK7ZrQFao9gzpKj
c7pHDl4UDYimqPzXxW4Cb4Ma2kvEZYfoL8hKhghDhw7J4YUx/rqsXxFTQsKu
lIusXKHhMzbo5o2OZxNqRglopZ8w8X95LGW5pFjPCSztD//mwj8+t1DkNi95
BBVZ5EvPvCrgZewBcTV3JzaiY7wze9oYu0VEAkkjl9I63dh9lGKJWaQWlgJD
NjDVRMyJ5L4pTtvo4fF4swDBdk0fzDes/2pJkhzyLzqXSxURglahgiG7JEma
alEl4xz65+JkV0AiZTu1bHGR/vifj2osIYjDAGGLahgknDhIktTlzQxePubk
xv8s/EHaj5HOd6D2bI/+ZfMbYLjp/3Mu7iMfzfwUVD62K5gqM67BpUptcl4x
hnvDmbvYeFuZadvCvUez1jxgpqbBbPTBpO6YIKPwxIuMmxHHo52cxCjAgezK
psi3ZLePX4W/ZIzPIfZNKjaNN59V8WcxknV63WXynsDZ3alAHBh3GKNl8fMo
BQx5Fy5xQGnvhs+4W+B7qu71WQoTrL5Xm/gFnWyAhpPL7QuziOPBLJ1O8VF4
aZT7Koi5S2K5amB53M22zsyP9+gV6q6Z67+GRwSpBz6T/MpYo+vakYMe4yM5
a5FKj7VeZqCjaFUEqhuELmHA6860i/tD2tsTE6NOlBQN/FbcTaUjKe/U33Dv
bh7myTCfZja/u0pHVKv0tj+Ir+ODBmm9ZRx06BJvYzAJXff3dK+ozzQ7CCMI
8DUNpSuOaysHo4bjTcWsRcvZHiHAdxrpYaBHRyehV88HF8T4FdrAkzajexG2
3tIz9/nGg7dbyhT2EuKsLhMzZCr1FC4dJ5+Nc2NQxM8zsdXZOpJPpAurIgHm
QIpPKjXXvS68dhPicxwuW1JHE3/A7TPe7ubFuz49jd8M7w/PxRKe9QNHXKJL
64wUkqd1JpQNzj5ESP58BRtFBWjfZbQmO3LiZp6yc1gqFPMb6rLAMf7+cf6n
HoO/F4o1xT5kLbFS2YKYxRp7p5vkfSS2QpVj3VTXPyFuS+g0Hqccl87gfStX
sRnq777CXfAZwtq/7qigO1ki69gS+HyQKbeXFaHv/mEbCIXP0I5gCoAjSh+J
ocYtF/r7zhhlIuY0915x8TPmqZ4lEc7O3jkGn9SvcqS6Y6T43+DfnN2lWxHY
9psfER+8TuldzzQ9dgYDG4y77I+C34pWOShviFjrTlYUTXc+AwJOy3OFODc+
LQeqj6qG/k9EiOlEREdizq2ONOIWxbp5AaR3vhL613q4znOyBJaTJoBbtiAE
snQ+Ss3rPIzfwifTGhxAMRygGwfCYRbSlHZvgXyj2B6PqdOYUzX1tmJRS7lT
GDrBtllKTi9AV2ap6tkNzoj24VijygxBPuGu/7WtSIIbYO+MGyQrU3PgFXPD
G5UWBTT/gJDcVLtGfsXzKY2qoV1QgXgD/abe3OK6ZJxyKr4usLKH+jxwV84+
lAp4es6fnPAaO+96dfFrVhleyC0O+Vcdl1PPYNIX1OKireLFESJR/v4NCkSZ
lu2M2/Y0jaYVXFMqJz32YJ+1GNqs30uRh+/RiIe0hBxOrYJesk4LuC/zc33s
wIVYqT8JXo1S7n+cTpMuRC7Y+pqyZLaKgAy8t7RDafUFm4EGyhfLqQBpZox/
LcfCpZ1FY1va7o3lvGFZKFsevZFaLf9KfdPsPtATbrkzXfYvbveYCHSDHhXZ
JEa/NDHbDong6CdonGxXmt7mlYjXsksNL5qfwHPXGiJKpvA8fI0QLxwK7J6R
9w2OfRJ/GOWE+WgqWHS95xCSxOmQaYjfqmYlEog0NT3ahV+Ax6R4IG8heMiM
BkAtLvGxv/WqOQaj1SXAdO37dkGmakig66dtUW2fb3kMZOUOORL633DBM6r9
MAEMMMrf8SgO0kttYRsmb9PwiEtelrHCpjDNh5qMaES8srVZCpZH0h54WnjF
lhOy4beh394OEHyb6VxKkpRsRrL4DjxfPlwFz5LUV/i+cK/F/GEEy4Cvv/Lm
b3Qsfnh1zY6FSbYr8aKJu9pGuRFD6cTnJMdS5mW5vc7jvEVs686zbZdXcO+t
u6cu5hnQ48MDG+xsk+ZS06/0UgXtwevhd2oOT/JlWNegN3PhylqBu5AhLK+c
bjagHTkduSQSQpZ7lPSWKGCdp5kNFEUu1OoXEWSCsWeb8ZRIRqIUrIT4+qme
6fwaiZxbD8x93UfSQ+nefjIDU7b1HIig0eYH4XeZpjVH0xc7LLJrQ/4qttCz
wDOwi1SG+pxdyTM3npGBIgBFhgUwyU8P03Zygv9C9eJn/YYbqrw7BfCYd+wC
OwPdQsHty1ijIdPw+7sTlUyZAibq4vGbzgCAF48Az39y0qRuoHrPgFTk7aJE
c2rcTrU2maly4HRm4ig5L+qasOjMXox6CmlFb84N1BSANnBKVEEUWVaZEkwC
V0KxokDoxBwWOi+ttdNNrbce4Q79Pa7Xphsq/0lsL/DoEc6lkBRJ4FrH1s7j
gn4ezoI1fJ58008d9LMgLlRD81Ce1PUC9T9H58Tha5Wq8UGL6YMGyPmWOWfY
foKosGrzhdRLZht9c5hxRiCgx5+5zU2N+XikZDhf0FhCMv+3e56PanTYnF0r
pwu5/gbAx+m1IccTzntDi0oNA/MFd90kbBbaJHJjUmzpisxG87nCGHlLuVTk
U/nfXoO+bs+dyx8XuDCESUYaHTrtkDhCrz9qzTO5sEOpP5rPbR2ckmISKWSV
OW0WZ8FCwkzY5qqQZ4P2xL6R82mCk0qERbD5CN5Xht/XYjs2wcZg3cfLAKWS
Aa+JJF1NmcCv8+23SgSXEwGoZhs6BORem28TooNY3VPq+bmv5nT2DOcem9xl
GaZgYDCQm0lgsN1En06R4r0m7AizfRmSx3VZcLRse+MBb1E8WeWQ1SEuUVD8
ogYcDZmMfFjs1/+uBmTD7cInyz9Kx/rg8Mnj4zE2hHViW95fga1xnSZl8aXZ
SScU9pSxvav4PYyNlqxgKAVR3/MmMWw0BAdZBI6RrX+lu1jXzqy3Y+y9UAUs
pI7bJsjdWI84kIiRc+iWdYZWhqoUphDIvbOXPqQojjfvTmjBw5F75N3gLFmq
yswsTmyE5N8oEu6ePTAcDXfOr+hS75aj6IEEJbumfTRoIRrV1xMPbnv2TODm
PRlF0spteOp/SWWWuH9shnsRn9R8gm4LtrHtpyMMKk+NQOY+jw/X5kIgMEyO
e/jvlEZcXBxy5j0Lgfx1MYlmwAhee7RfML3UXhm5Qsb6BHtors42mhMnj6gq
26Jsz722lOxxW8P5UBrhz9fEOnd++KW41zn9sEg4huqkl4l6RECP+YfvZ/Qi
F0DvbbA9MDwIWvgijWhXRokKtd2afT2PgTD8y6uUA1DM9B88Q+vmwyJBQ1Zz
zUZCmXaf6abnz4bmubbHDySrnZGpnw68gaIUchY6ewtOVT+h6e08fVyp/eda
1wHmPDOxJkOrkzBQ6UJgyr0muP818z/iA85XXwTiA97wt8VgSt6cX26jG2Qs
F6rvOkYCxoAGWFRbpicmCttsUf6ufFZP7lqiyyavgzDBfKewjSfZL2f+1bNH
KOV2xpXuxrWdF/Ts2F6p78IhH76ugUqUrxYe90x86E2f1DrIjoFrQlEnINpJ
5gHs7Wwk7jcw2ft3Dzid1FhnvhFgj2qsnM9W8DWujS0Oahez75VcdM4dcPJ9
18FHQfqdtL5SGVS/Tc2nXBSUMFQymaG/ui2eV9Zxad5kXiyq/ROOMxvmSXDd
tVnLxPhVsz/Ia4v7+zcLp/27NaawHNWU0NHElrjVkF2+6L8oWKF/V7KJtw7a
MFCyAo6FhfcpXgj61Vkoxa5/cMg6Xn0cFibFsqtXUo5A8Ve2IfcKbIixwEMx
KrRXMS4NGg66fTeaBq7kjq7e1Be+U7KiIIGrjbMdMS/UteRlOPcDYhLbsHj5
yR1q39UY5TpkbX5HT1JQTQHSFyxpy19i+iXu/q2911rJ3qqWck2wLBrs9AoQ
aON34wgjDjTVR21/wXKWHCOxYFHUfTGOeI2DZqnVOTQn+6oY8rz0BpqVBBO+
rxyPdpWJPLbcmEYZLUdV3wcm0+HylDEDdWEIyb4ZZzB9DPx5UEi78UE/6b2p
uRLuaNmR0+jGL6B8PxOYcCQLjTh9hw3Q5A3qHy7AGYMMIqmf6s8DIAP5z06B
J0TMXCDRLAbhliQw1Zg4fhNxp3VLsU7B2sbfn3k/P7PMvkcgyT2zbzv63ilw
405k3Yi8g/Rhbq2SKO2vrjBzg+nt2gc0Ke+qOZTJqQRm83CCSwdUXuP480Cr
rb+AcMdI6JU5y3yhMERGHqrWnHFusvMiCmbhTR5xul8B698He5qe9rd7Txb1
ly2/uEUhPl8QedpPMjYbbjDPwCoHKzL+tiwYP3ZJ9MMQ/07EPC58rSu1kBWc
6nuXatRGZweJURRG2RZEFu9cOiH0eO+tlunkiPX10nnLH6MwoD/Im1kHeyOL
HVHqrsfcEmZUDwlu+iJw2Haz+G+UkT9Mos7AuPZ76WdaHyQ7KEKZgi2xjWi4
LEaF8wv44ugR3heagE+sY4uxdm8kIMUzh5BYkslQ2j5PNRqwUM1McMSBhcD6
EV5d47rmu+G80A7+Gyf5Mmao8DPsQF1wj2J5F7SVrCnx7iPPUNu9nANL7EWR
Hkrjqrs/hPB3OJJwDX9nUncZmGNozynpUfU1DpCq+ADuWsjpIc6H4KoIg+El
zoGXaHBti7ynvg0eTja6MCaBG8k38dDcLRyqHxPlMf+Rx2NsNTiifclSFSqo
xNPJpcJcyxb/fJsro6uZo4XGO9uaDp0r2ZboFU/3Jgn5Phk4aNJiWRDR99pd
wSWeaDL0O/vsErd6WlK57Ug/KKbNev8jYacUwfAAafx8SJNob58xkvMIZk35
0EYNo5YqXZQanwTUqaL+PUQ6GZLU3/E8s1JYogJQL4pgu6lP1PkcWf1BjsGH
OfHvPwVHmbIIh9Q8DegpES9SyhVXlh+awoebZYxQHUGhuLNuxV3FAtR5b99K
L6qVF2OUEAyTT1KkAvb3Qu/JhQbq60ZSVN90cD8MrmCqJolIb7D34Lo7slrE
D1Q1FcgK4j5IpYAk2nUhN9ZJdBDRLqhUCi16NH9uIeckJixahxPLY9x9qg1U
UHGQAagnGN/r8LU6YE32PMdIyLfuZo80crwVd+7fp9EaBadlM8VuUsRjeNXp
P1dior4cdF53KXtWsXm2PywWWTMw9nX+Hyzx2TdPeaBayaq5R3Mcx8vo1B6V
or3yNiI0KSJsQTpfcLeUsE2yJhxeC4WZNQHQkf2Qe2BEzqA+zqKISCV2Lh1Q
MGVzjeLRGs2zlnPjdOQfXq76yFFnnDiY35xUjS9T1Djt4rAm1rvqLmCXNPLN
pTrVDZu3NsMhfcs2zOWAyMTNeO49XXyYRawt++xFvneJO0H/SO6uhN+iYZsL
ctYYFtCLUgi3IdkGzgIRIRwMvKfCl6qKTUA/S8ZJpWO1BuFovgFmPQCFzMsg
LMOxzSHZbeGaqN/xp6maUW8UATei0MYfdNlUAtcH+rNNmqJsx0yMOZQuTMkA
kVz8B7a8b44q8NJbARCm4qD6rN+SZEfZKYll0ptYit61X5MhyuVTyiLWpyeJ
mHTWq1+sAGK+Q/c85UbCoHPZeKKVDV8ytM6nmTxEYjToRzvWYQrR6qfhR6eJ
ctMUa0V5dRBpo0EbeV0ZmBnbEAXjBudhZ4e7KXefS7j4J2fZYmos5uC/N9SO
9MttkdEHyd8sTYBTtB27XhzBzA6g8vtV0FV6nGwG8W+/lu0UCahPKxDXa8jU
a9Gi+4rrWhh5VP6AGEPhHiHwaUuGeOtK4G1lST+MTxjrtloyqDGohvYDxxyJ
Lvbqz8QUj3ADLbeMxusnTAexM1+5/ErrGt/On83KNZ0LnWlefm6KaeX0KRCN
ER01ZncL0vZuJ93WMvFGYfB1NKgXdDE9DJ9e18QW01Kg5HZXgpdp3uKTgBiz
NjexMRaWlGpniWT/Z6Hyxgsn/mIJdKOW201/fFlbKjc7hS6sRcx192Tz+zdC
PDdgwzDSUEgYhlRIrTbbyqqu9EahKhFGfd1B7lA+jnNlVEmFtHryGRj09WQo
U331soq9U01W6Aspj5IU3vkoe1k7AJiF8kUVPiAbSFMfnUB/IBBFB2ZstT+F
L68N3LtWtq4kBbIFOWHkZ2WG5WxIbBIRVScNWcSA866krl1YNkgeMyIx3Oah
4GLWmzLjK5Wl9TgQB7EGGhUkbeIlcppIdQ5Nssjdnd/G3VqWr54UVWyW+pWp
uetc6s5gG68czvHpWZRr9PZI4hVYYwjoVXDLF7Vj8oAF9SMudnU78KIiRw7D
821NkT7AX9rO7bqhTl1tqAddU5ncpXPWBkJNwrCPRBWtYTOK3jlmINzAuhw9
ZCavoU4oHTNwFR2TED2IJdiFC8oynDOd5Ilg008Ak57faQR4nYCiDWiBhWRp
oRPh+3GGUFKHgtcYw4h6CLLAq9JC3J4V7zyG/DCvIQDgamCc334Byg0Zf0tC
3+FdbFo5m3oV2oPlunioysTrN/18YTOMsOpHcTD0a3FoDukUZpvHgwkiyEBM
9sRMC2lh8afRJz9SWTL8MK0kNL1oxAn7liqofZVCPy45IFWbhCiGYBJPTAWQ
8IyCcbxXkXX8GT1WYHuIRLDfeMpB1WmJkNhu+3C2nNqHBghHmj7vvkghY+rj
X6ZYcdX10wKyr58n2+S8ZIzfem0Q40XeSh9uscLYvINCGz/vxPffX7uXON+G
qu3jp3n9BzeGDzmclcjv4T3zZH/kBaC5bb13hJz95Cgoj5iSHr3mte6bCAoi
nUc9Jk7QUeCwZ03p6BXbJYcyR2FTCxRCMYuwvSyqdzI3zHr6X/4ALamqSeAy
XZ1kuBnjRkBDiW6oo79oQd/LHeh7zFknRRupAY+JOV1Ya3WCuDFHKbAGAnlq
RkFJ1HBowMAZaQEAwv3crakylzFGSzMJf0koNn8ZRhyfMJPXnXy/gxovSuSs
Iv5T3RmicoRouGeZInPX3ThK7UPEBhX0neSCfEWQm0DsGcppf7t85GuG3CCg
drnmt5fti3lWIxtCY4XQrNmuF8efyR3p08s7HgCTOsrQCcog9LJgm5/gOEhu
5eupwpemgeVFXzazdyZm6D+ERkJzW/54t/eVF7+MVpOtxRkC+nBL7pYjRttj
K9CnrNydIhOujkVgxr3Wuwo50eyilQHPraHdc3DTLCa8RiIL/JaRQ6XF22ej
wt/bDhsPA571e+8mdmMoxG92n57yJ7KP+kg8TyXvp3w5UpNw0AmPwzY1s5Be
3JZVbL8j9qrwjHwyj18P4PwXzcOkjLz8Ij1GCask+zMASO1VwdEKRneIRCHj
b3HnpMOWahHLvjsIU7vzU7ib+aQRdp5Oh3Qebqo0dvX/vQDqP5Vaf4xRSg/4
jVHz4X0z3X0qhRf4KAKRSNC0ux6+Vw9ggydCbN78pcYo3j5Y8r8WkjPM80+Y
kDgCt/B5F6rBa5aBSJXq+HPIq3TYSWCz6tveoHfq3lw7ApLTqAjOP0wt2bXu
MbhM0GxSe3f+FvYhvR9TKX9ys55rJzMsnM11TPun4Z11NdeL98jXpnEubknb
ei6KYjCcwZ8lXNqr75xHBW6oxqIbuZ0VdDffys+drSdgD8Thdjc4+xAkSi0o
zfKu4nvrTAHZ3GfFVi0gvr77oid+/teF9TYtyPb4J4xkrxe07kH8DSJ+zdr7
RBAQ3ZlJq4TEopvVwkXoodiZE1BiPFaXPx3ayJJoMgbCGhU8VIyiysoY2kRB
zYw3SEtD+ANsJmXxzBNfLJYKB1Tp5h4OLXx3Ig0UlFkFnyZyoMKH6YPCxbVp
A6SBxyYcwTT7alBGZTKik3YvnqHtkwhYHR+Y7rQo5bAfHYP14T2iz5QWaF5I
mrE/zURmX26wvUM3OrIVMjxqzBW1i/ARsBXzD8hJFv3H9I2gX09LEB6DBDAC
0PPaRsPaC7ra6oozn/UIxXnkQSDfuA6WbMDjP28wcYh95LTZQLaAE7BZbOgv
W8UwBKgOgZk8N1AkV/dW1RXrsS/prUQgO3jJWO6ggeaPAJZZBRoWJw4sxtyn
0ctqMGwEQmexbYLnn3mK7vB//QF0CmZcEpld15PfUB97gRBfuzip9M6Rzld/
MniIaEbdbswJY7vRNovJJYCjXyTzkj/H0HKr5SAKPhXlaOqG7J6WocuwSOYT
hOdhd9Rftcv/+8CeFp/0FEV5mmkjRinuvlfzzIe8inOOi41r5Oea+zfFXupB
7JOGDZAhMdguyEzR3MD4eSHEUGWupGBQvbX30h/hLr4ZWU6seedJTh0bgi6j
7ASYdc4ZCPf5NfM6yVxbTVrxKNIm0/RXge5gz3KZUKWqjDWQksaI801KddqP
gbWlaAe/uHfAx5Kgpzmqk2/0Al5GlpEyFh1LE830YXW4i2d8Mdhycypcg2io
gcg7lfH4InawMJtKkpyqZa9JCKYUoHwz4J8N8fWiJeIMryhPtZef+sgfy2As
u145yxR3NVWjZtLkiLqP3utZ/9r3kXy/27vneoAq7bEdbqC6Iu5NtW+PEM3x
DN4PSDrsv2wfEqbqEblE34cSVKiyRGrMAUgC/Jzd81vz3dKcZATIbvX6CGRG
KJfAUOQJ4eTFfWvo3vz77DZ/VibVqUIUD3UyrcQ403TgVO8R0eyjniDdojl8
e8n8gWotnCSuNIE1PuqZsv4d//QQMIb8iMcVcFmlZFvBeh71sgzAvE6RmoHF
ul5Ig1mjOyS/Zc6lWQkYPpXBz0iA8sIUGP+unC34JV12FQ5sN6FzmLY8rcXz
FU6Dtyu2hPQrjxm+EF80oEaMSwlcz8wiyfIPZNNqjZmlFy8Deez1H1gPhEQf
EPUDuWmurE9OjrvuDqDk1zVhf8AEspgCvhCP1QXh3+Jdxzp5zp1ioXy8Wiok
tTorAgHMi9DNHNggMSV2z7PovPkINuFAYq1BbXSiPf94jAhQKl7gmh4TN+yo
kHpeem6KZlWRT/aH/il2yNdaeOQI2OqKGtHKCFTnG0PVBhhNDUiiiTERc8Hb
D6d+OElwRpUeRvJLj4Od9i8P5QPKWqwdp1Uzz45cIWThJvG2bwnXw7yO/F1l
F5Ai6PDWd98r6quUmLvOj6WWyuMMaRuaY2L6WZWk7N6ktnCrA/2uKkblH+UI
K7f1WoNbB+JUZXds2jz0CW/4Cn1Xn4tNi4PO66JaLyE/DtZwr75EZ5+tMnl7
ytqcemXophzfCR3PFbW8uCEhus23cB2z2fWEr3gb6AXhutGfzypCbkC9Yg2q
/um7BKBQ4cRrK/IXTrtNXw9mxUgVn85JGHE2Jmf9rvgDMk7tiCPlnvJ2+/nN
4M/OvFCmGkemgt+eCrmVMUR6szhm9ZgQ2AUfM49OLCvn2Ulv7TDHF5PzvhLS
9UveEYPG7qSw52qqLLvGXzZV1kxpvSFZwnZYWcNWWFJCnU7DomRbs04iIVCp
28T3rba77ltDqrs6FL7jwfVu4ki7WQjYp4v++6JSWIVOPDbk+XHSLQR/vBjk
XGtBaVpR6AioL1l7Ax8m1S2V+t3EUlN25rG0C4frdGp44akdk2XEHLzM3jiF
Cm9ISVt0YTLMiOr8554WruCRMFTnc2NdbK8oah8T8FGvmUlOu+/mpJ69HSCi
6PFeEOfq1aL5i0xS0b2AskTLuLvZc+uTW0fZp0GlZYcZizh44bqQvyEnLTdQ
KzFrRCoqySbAbxgH7r6+yuGkOjEJaihvknhWQesb4jfBHW+VmqI9nZUdY7CU
peInYQRmnpxtBxNUeV5XeHRy/Biq3rmYCrHOgMaPVZms7qIYnqxLXQW7TASr
Aqrlq+e9sHTskP45naX8HY+awhKDym80ZP4kP3jjwvFACdvdsPn/IjqUDqR0
D0vPk6+Wm2gt+u8cHHqvjDxdUtn+zIxuF6fK7HEqIS+d6Ffb66QnKiB15VXa
imzrNQSnJeCCOAQeTRSVFmob6cXDBjucBP5PJNMNPrxvN0g7iS/VSQTl3m5q
e02p7em6VPvG2p368zpvHh6x/UG3oqumF2DUHANUfz6tVRT5DEk3NzL7FpC0
91jEMf2QIuHeVkqUMnbIr/UGmgGPYTDERgYjHATvJlygaf9dzTsXRByZnkf7
Wbder1UQIakK5GdMn+0ItngxFufE3p9i8QL7xV9FbxMKXuCOxeP2MY5hdKS1
iooDOh99L6ro5nQOkc28ScwX0rXvg0yu6iU5CZPYOMbt7dmFC+1o05uAnBo1
8lwu65vk00iQ/UzTKqsMpmhsihG/gbX/IJ8BKkmLMx9hE5bGtB9yweJjuLlO
kwTJ91D6uI2La5DUyUj1FcjvtJyzRL0QxCZBoEQ/PGd+NQnupqKYHFfuDqsy
gB5ve0sJxQSKT/GkORSeylD8XqjKxE0cul6DGmXNqvyXe6by9bfz9dCjWk3Q
7v17GfOJj4GHh3NJJxnZo/iBFDlGt263uc/LMX8avruwyUHU2KJixnM25B22
qfSqRzFd1WSdajB0oQnHE558EdSzsuLKUdsHAB9aTyqKYJAOLp33CutOzIsK
5s5qSUbs6BGj4YlgcuGOPb6qj0ibk6t48bSMEiGr+l86wdnH344bXiB30D++
lMYoA77kcOpU2G1eGb9pQUabtzykAhaV0uHiPN3vx9AIqF3G4cz8+u0mBnms
9An9vQ6Nx9k+4RJGXaLrNrRX5k92zhR2R+x1SKgQKNRTU/D4EEVOQzswC445
8z6pkAfTh27Hq80V7krJuCXtJuisJZucsNX2JFb7Kx0Ozy0WgaJ2+4HFi9oC
NexnQssrnHfU+1HArid7eamVyMSyPKbRRcIlEoTwHXoncxK0ucBdCIWnras+
8aS5Io0qQRQrnbB7bUqd46JTD73OSBtAEuqxiifn+gvZ0xwA+TeRxITBVZZA
2EHjgYXHn0MhxIIo1Po3CsGeQ0mQRPmNtMnqbFQx0xWATNTXCjl7HRgkwAWR
pfoJ+lhlWrpdr3lXdWGA1F/gUR+Z6MmVCY+tSGmgqbVU9rOcT3epZxk9fTM7
Pr1dUbWmslG/qpAFGof4pohuq6vjRTibSz597ADQcVOu4KVMtpTawdEsk4oh
V2O4vEL1n2BDzhKKEpE+7UFGR4G0Xl9ivQn74dbxJwwfdxOC9Z7tMWKGDSFv
oZIg1yns6tDlve8nAgLgVaXt4vRvhl0nkiucLuqsglLZqAGCAT6lsFY6Vydq
d5vTeXQ68PzVsKJffRO1YxCj5W3vVhs2qsDAIgFXLKnOkVst1vYsyd0uMB37
e5cCv7nwlUxzH7psNrk0udvcZyID+SXSpUqHLP70i/OO5hDpl8gX9s0/vfmz
ensRhUbGpJf6bS3rBrNsD+a6qx45YId+0FM4vL294Pl5psyiDYHqCzWdSwbM
RZYCkHaEj3GpGDqAu2rS/fBqZY67SzUwfjfIj7w3PIufn/lWRXW60yDMdsn2
L0R22hCXiU4bA0Vh1ho5DHY9a4og4f0YNcwdqXCd/gYlk39iGGV+nCSGFy/a
MPvwV5AWOssVv9ungoipu7Essc2mk15PU/ALpClC9bOOIY2IJWdO8GDBzyHp
rbjyhguiXrgptdYABVhQnq72TnR20oBYOaGX4gD//woZ4OuFP0AQ30UuMQUJ
wBgpJBKi1Klv3L573D2EFSgvEyFdR0MUDL7tSJRw7IkI7AsQh9VeYtLQWcAI
gZp7Zu8dEYDA1/803nGqPXfsypIH+wJlzSLAPvcQ7zqILdCAtALt0F13RJU3
2kh3iCv70Gli3Qtc/AYd6LrM/6sYKKd6c+86X5m4AuxDgyY33ViJidmtMaCp
2RxeMRzRH1kEEDi6D+lhg1ixlwwk95b3tg0FoUBYozVkaVeJbRZ2dp9WSVvF
Vs2GmXT5VLNV5DTWAyDvRWWKD1jEF/ll6EeiTi41cX5/VvI1NWfcKWwEG30F
lgIxFC0X3RgswtHJTTDwuFrq720u5sVn2zcYbbrjicvN+3eimTAUh2TQhIrO
SOv3vhFBXIdc3qm//iipb6NYBMgZQN0G8JWETHDw8VQwdgxpbep9+3h2r4Oh
NmzQ6F/LxrXUOriCzhcp8mGaM1FgCilUGJ/vSvEo6qlirLxyHePoW0KZtNeB
3MlPqSrDtb8fhtV6zsyGEvLSssxIzqmRCDgiApdYWY7iUP/rO0EjKbYaPPU6
3l7HuVFupwC9+35hwlzNZPLfFzV532Wbgk/7chj7ZyC1P3wEsnHpcNTDdM5K
Ex2M7VkaK+YvU+E1P6+shu6IREdiK8GbahrHBXpltGBOGz+BmibhCgRVIfpB
hQbKyJSHlg/0BnTWlAvF+EsGEpImd5SFj4TJ6YRFbie+tqPUXC7RUaiccKCP
ukbkrhkloiCDesjxD5hqk6sIU9MXC+m0McKZI6JxbI1t+sj0/91AuV7sgV1w
tLVIjR4WhaHXC8SVSbh8CoU5QD6leTX3tkBQy+2Fg5H+tglRxJQQ43dzEEbV
eM5LLzH8WI+5khOQp1zOboPNbXKjiAdrzw3Bja0auvCpyqUdcwfLVJgc3eZV
wcx/UrHUjJr1l7mWslOgDchh3Q9+qnnRbfQ+au4r/F95fGoQbHIvLe1YZ25L
bmhqsnvnNiaUU6uIFKDTERpFD2kFU8VIFOyk/DKdI+VEZQBK58B1MUlE3PqX
lQXHymu4ZAsBCujaRlfvgvnZZP8SVoyEO3I16D/z5uaG1qwWCkqUTL6trTNh
9Omb1a6hko0otRXPDXYBRn2+8cEVMLxGtVyqWNFxdMOcQQRRF9eFrL12DGcj
DkyULM/YkmbHR5jnb87YcIrMJIQX6hBjp0rAzdWnTsVs7dEjLC/GkCpfB6E+
bRJx1XWgH9imHt6fXlCV1oLxw2zY2VLoPHGSB1tP9ttWV59dvp3+ViRPmmu5
UdMlqX2mb0/53dAHATTuTqa823C3tP0ngCxLWWzwaKojox2v56IgTcTYEKJh
cm9ZGY76UAEYSW8efXHzWpwf9J3gnZ9OltviQfPGvTy89J2NBTH0+ZwL9xxZ
819f0scolJuK4fANLUp6J1s+T7/ecEtjfdBSyaGcamFUWdjDFFN8K91GwqSC
2cDoj939szj/c64WugYEAtQ3przsZvtZ5zTL+5BO4x6IyV5mcKMu5qgyPxXY
99jp7yziz6bLqmtsFXL85+KHinqzjrP4hs4hBvx+vdR/329npfARWALuxlXA
M5/ydyv6tAT8ogW6CTnKudzncmUwwcD0VEYNsLhHLScWdj/oJvztQQAkay7+
oNNgWhVqGancvCnghO37Hou0P9crHgyjayEN3aKJ838Rbl5ZLIf9rvbmH+JD
U28QpHJTuVwq7B5fcbps8puh+Tw5MtL/QeRqQo+huxftzNWWH4UMfK+p5CRA
kXe3L4d0UZu+Q2pbL8qLt0/bdKpYRghRe4yPHqqi8HOgC96IjjGpNNA685cW
7bvG+iDV/UmQlvOekJ7bFi0/T60MPW5SCXb/saLXX7zfHq9dp6JfqLEgbBeI
lq+HFF89e3/Jw7CGKqOQLiQHfRyb3kHWZVqaJJx4KQHncIUd3mNIhDbFEC8T
R2iLbBPgbE4lE9TiHaWmindsACd7ui9ZMNyD/Gr0EIcF5hy4OiHi4E5Lc26z
/u4bsFkhuxutX4s10MVBcRX2BMfnMqYbHykGuIGJOWUu/hnBNO/DIgSgi5vc
ajUQXIC7BUQ+tA2HSGWDzb+3kyNYjuEDC8Sm+Sj/PYSi83oIY0dIMSRDiByl
vkwswDm1vIW2bYfksdB2sFM6kRzX9NWsm5vz7/IT5CELM0oBJqiBHRsZNJOs
8YRWAcIIKF9zgkMVNRWZu1fxX8gESNJVoKTc67lmCISbWKoP6zR5CE9fuvUT
jrYteAz7jLLiHQ3msVJz8Xlu5SViLhu8eyDac5KGXUlQRLy7aChnIczqbCsk
e/IpEOws67WOgkTRn9dl9c1Ff94b9/qzFq12OQlmlKmMWLnN4/cHInR3DfP9
KCEC8Tzx47gT58Q3Y4w+Fua0zrGFMTyKJyR1tjJDIQnbeuS7SETcekuuUKJr
2y1HYOagBrhX6OeKC9C6YdsCDkMKJUtkx51HqhvqKANOI6fS3Cla1mNtYUSu
WRq1Ru+95vjy+eK2FZMlePpU2AyoC8mEvWJGY0tGC6luCt5OEg2+lnfzcBTf
kJS/q5CT4ZMs/PJLV/VOZZuQNyrDEX+RjqOp0kgU5JzCmegEFalgZ7ByhB/T
0S1nLAPyu406WbBCY4ELcpANKfcPMhKO2q+pvEMH0jACAX7gU818S23pC6xF
1eDgyv2kPoywJpudR4LMKr6xH4INHw8Q4b+iU8oModZRbmt8IXbtis1LWdP6
CT/u4Esbexfnb3GOsG7pBvjyOD4CEonS2Nz6ZSxTgjpMpXU5p72UUTNVaQwl
1BJauJVnN6tOHg8X3KT6E48RSjUczLCZUhyhW31lUqk2fovRi3AW05KI0OKT
dm4cEOBreeVJuwwi3aWiZ8BrTztXkbZTS9w7IkiuRgaD/MQ+R09jf72+uFKM
EoulzkwE5sau0SvWNAbFNCgNu9PlBWtM0uIGs4aZFkE2oS7ppkpq7QY06OLQ
mMSIkcw0HGngaDjdQPPOasjOi3nutFNMS6+PyTkfU/CfKv0UM2/6jv5oUkpE
3vct+YjqOwBpcMBO0zFNhhI+ymMInedgCxyLsbTNSa3wnQolROHF4nvXSoFv
KQnW+CqxBJ8YDJc0jGUu9uVKNaxyf6lL86RQT2FrKIHon/yzPkciPPnos+sG
EXzp4ANxlWzqrywjojt5NAVq/eFsjARULjvUtl4jIr7WA6ZouMsZvcI5Ys1c
hbN15g+29up2UA5QEvxd6s0dHCp6W/O3Yv3kOiAmFEJGA78zPqjaCqIKF4Xd
ze6rdoQqrmPxOpDpOMOsFuDvLZf7K65n3QJ8CQSRSWRvXB4K27JBB3Z8Xdh0
IN04w1TRcwSLuTr6fGMBheXtS84Gqo/CegpXDgVJGbGc3yOZsZMZskf9O6xT
byN+KFFkV00h/j81CDyqv3WDM7ymbSyoxyAr/k4QFVeLoMEgliAwh2kzAz+X
F+WOUW5IlUVQhia0GIeCw1WpcQYU4RMWVtiRFnVmzLs1sMrMyxqLEQQ9R17y
CO9XDgG+KO9/JrXVRwhyYbFSZ322AHW3JEwgg9HFMlbA4fFvZWhkdEZQjnda
QP3NmN/PH1n1Vz0mpS5esw9bq/CSwWV7q6QNMaPfdr4fHOAb5JaQAboMJm7W
qB+QO9nsCqpWcEuYaP/5z2VSTUOOOY4vQ2zi6bA/Hw2gTpfj4RnScjY37jlD
jqOQwKiRbWq9y2NO/YWOtpVX32B9KG0cUdXwwr21Nc/aPG6hMb0uzKdbyI3D
9HjwcIknKnajUK3IMale0RPBrtewYzkrh3Mp+pM3D8KTeQdHXqmnerl38vkA
D6gFz6ffuBYCVVKFCTKQFD7npIUl5CIRLBrGdRkCvoNCkqp1TPtc4UFL5Uzh
2zwtj2lp1eJObLpmRfkDbxzJzy+W8RdBJTQ5QMdOXnRGTB6CthUCSOtbJdxj
V5/7es4b1B4MFJ41gE6btw8Zyt1hnZLT4VZRFH9az+4MHlJR/3a4/Kpo2xc0
aBMST4qyPYNoEfLjy2Kisp5p++IK+VsMhVOhfr+DWCozErLPYYaK3oqIA6WQ
Z8C/TPqN4wxb0pEM+BtKG9nf4S/zm1a9SQB4MvtZL9W3wJEAZyirmGuugGzm
70rKWPKft73N1Nh6BRZENLBg7gjbSqn8I6zAsy+zKE3z6f8694b2LMRvf+wO
4oHuQqcjy39XdK1ptRoGnu1cs2MC6Zhk7HiaVLD0csTz6TMHfMIwWOs9FVOS
KLgNW6KvIx2RBOacaaPuOhWD52QL5lbvn/VhF+nKTYO6WN1hXeO4QCHf7ry/
+Vxu92MHdKILNu5/1gr1q8YSkCZW5VvOjn0c6B/e9R36erWdZVx/ejTzdXnC
sqBIimNVkWN9dAXGWONltNJfs3SzmLGnSWDGCkYjWX2D79xIk8A/vQgM0vk3
jkajGxL/cbm+fM8zWlOX9IoCTiC7SrD9cHarJkAiMdd+bbKWcdoEInQDvoha
nGS+9WpgCdy/+iNSg+OQiMMwUFCCdylzoypfx17TsYADuShdM4C110M7jVcC
XogUI+a0n/9Xyt/2a1AVv8Ix0snVmJZrmwbMbPprEAX3BPquEK0HRneypyVK
OGWmkjIMpdmI+nkHpKjZU6cUid17tx5fjeSGATF5Nt2hiJ8Qy2bGpIE0r54J
NPbINcO9uYFY5MXf5CaIil5iPixFFy4Ucj+4EOq/w+0q894T6g6Zk7yNMNJZ
yZfJyGRBFU0D3TyysoyjY41Qj+V6qItdlq8/OFv1GaHq6kWnVhKGXFtCZPPW
1/FzDxuH4iahafFsIc+SXScWImsqXdYR2GE4Y9r3mVp/g6JtXsWZ8RyUlHU5
LSWlxWQM+GYgWUv2VBhokOaIq5k6CdppbqmGxTFCogsU6ZtiZ48GM4f7WNNI
BVnVumEp1D261+MSsRHxP95f03itVJZFMLtt7Zq/k+ajql2SQEMnsDKyjZJ4
UKcPjhzF+hGX3aSFP1elqzaQR3PR22gI9Nz19ortNfd7GTf/1kk32gqwPFfU
NrVHUqd2Us6L1/MIY52BdE+8cVP1dmWinffnJ/VYkrmnsRhgoPFvmN33bc8O
ozc+YZ2C2Hmeb+jTmoqz3nqQCIIY0A242AqFIM2tiE1M+IeLifazd3P2pC8r
jlKBVE4LOf4mfIOsNhz67AHJS1t4W3kKjGFEi1+9KOID7rEeVW098zg7WjVu
tBoDHGMXLwmgkpqIAkZptmt11LhOZTrQ/sWAJBah5brI+92LxmjmhZWukz13
0t6m3lA3iyNx/TYu3Jeu0cB1LWhGG5Ct/TTOG9C8ufBR6iAC2vo8U6H7/S9U
28R+LKnsISpMT5YYxCs9A5PpH7HDoOMedLX+IaBDGZ6qhl7JAPHr4zvVvLTp
IOPwtgaudyIS4km0ZsOT0QeArfr9ggk3mDw0asnDENNE3khuJzUoF7xUBNS4
WeofCTHOKyka+HjHb/zZmTUb11a9/0k39OoIUbT22jbQ3I+J33aSQQ45Rqrd
gs4KGnd6cOgBQvcelUqMsH9jcMqpHEmKy0+FNpdZnbIFRUKSmoZYr8WSdH8d
eue3axfAgFETgtlAi7DAwcr0SgfTP/gYe+Xh5qdcoekWd14ef9JwKg57n/Tj
uTf2LC28kRsH4FpUF5zlazIkTgX1YmF5rRrSSSDZENCjp84tncIalc1NObs4
tPRoziu2PG9Uudy73wKzqMNLFlE/GmZeayGd+5LFUiei3sS9qogFldH4TvUa
9IEdUzlLekZ2vugRHShr9iWRWj2vOQ7C2TXouoK/4M8j5KLdD0TOXGWeE9C3
Wy5KaBLzJ4q2pSbtNKvf8j/YdJJlbPoVYEK8NyXgEdPJBfc/fidEZ5puxdSz
bggus4t04rykPzFKAmfSSr5RjxZZi6YZfCmPeN55bYhTG1KFQiGxfxFYwWUX
3fgygizFgdlqju/5RfxdmdLVIDzZzMFXBFH/JjSWupvUGp8mgrWYmvnzc2qx
NKfldqT8ukvjkrwyDJ7jk7seE/FSuwUN56FWG2s/58Q9w8DpHjq5/uER3L2E
c3lia1Iu8xudGb98iRZssPJcuiPCFL65mdpkn4pFcbTySJYyluhiRr122Tvz
I1hwCW1Q1W92U5sb7FYaL1ujgvA8LixW8AXD/setAh41b6b8vur8FwrVFNB+
m4gr6Unb3K0DznW9Kk3LnREmCCkjPLk02/TFiCfQGY08XKb5XzpGOclfnFkh
DaSFwWdiIZqVRb9v0LP+axzfoNwYZ6oWro1omMN97Vpd7ZzN2ui2apghjjZo
uc8G/cAmRx1HV0PsTQwzk3FUjFsywwd4Bs/GGJwagQ9pEKOcysY6eToKmSs5
/5pPbFtJzoZpRRpuPSrgTF2dpzmDV9a3QVCVws37aWZNQV7bOu+lEB+cyug1
FXRAXZwkrc3assRDTez0HjnBapFfluJwWVGDTFN/+rx30HN+7J/FO4ZBm0XU
u/OTvHfiB4YeqSn1pehXtZ4wTtvLWZI+HXdDHXlLhSORYLDozfsuqwT0NZup
yFFTpYFqevlVJFEFSPicObbk7Ghzs5AV8SYoxZKlm+pltnHckI8S8Gs8Mvsc
6n0oOxZmXs9OO2PQfqwdOYBtm8ixWwKnjlP9W+apX+mrgMD42wRI0LkDLukP
3d9CBweMh8Pvq5e5b6PJszZ3lJFUA1WOJxV1iMxuC5pQWEbHGMeLusc/ALQN
wgMVLaxXoJ5PM79FDsdE5pGcv9gidTYwUz0cRZWmGb56DaREZpZf35BTpb6+
fcbXrDJqgPxRuskSntcvAD8OZyqoroWXuIcdCSUpA8SwCY13jEaZQEg71jUF
nUOGmtlxy68JxBE6/NanZmXGeXKIDV7QEks8bORNkw/5Dsg3CN0d7tAdJvV6
4QovC1fIiFFGqq+akwK0kXDgzKKGEDedZAx50I5UzdutJpZR51d/a1mcjOlC
Lpu1g77vYJ/96kXgsFAM4bICsBRP0lFLwGEuyO6f7+t8CdaztEdg5TCQVv/l
5xencTdP4Cy3UQs4uedch9SewOdykQ5pLuWaq//8E6Xx0hDVje9oNFA0+W4i
+nmBZ4DUMVijcjzdMY7jiKI6Q7VRCkiI8+Um4VpILRhjvIYrYo7KyBYJnJ4F
tXnbvIYIJDXSpXz8aq43StZiqsWHSZ/PkL/3mqd8jQ5KzxfESQFjTPfVAlOQ
M6dB/2Tk2AqiWKIoM/q5cncfkj+Vo92AWX8KFcU7MjKncMuiDlMz33F3W9Uq
hkfn+PCCxxm1xMlrWjev5a086mECkE6ToQc/iFUh6zYrp5+ZmWEt8B/BxZsW
VipK65aUYRU+LBv5KIA6Fhp2N9z5JVUf5T29FG4XS8wN2qoEjMLtqogNvTdu
Nm1bDEpM1kco+nssW1pD2w9ZiF3khxfNmRTtWhTi5sNItDGGfeX4pNVcIXev
QHyS/cik0mVgjuGVMWu3eiBiVRI9PXELxCTFYLERLTPnPJe6OYBHcp/IXTzl
q/WD9dqIcLGfibLX0SF4HFLvq/Wj7cqbkvzvWqyqhEAROrywDG0fZXTS947R
R6aq8Eu0otQ1b6dFY4RQxJDF4QZl+m2rTM6yR9j3/dVsorabjdAoYS0AJ+h5
aIs4/Ye4hdfAdPD0ymVyuiGFUJi1nWwSPmhTd1H1e9KLGfglEnMOl5lApG5K
mtRrezLmL8BUyIOnopb6xk9WJhwncwoCm0O33JQgk24PCz4pC1giayZzrCa1
iOxugE0YCPpbhNDbrio+IZlxbVIpRoV5h0bf2V16IsHi3WX4vxD/nZlnbX75
3USBY/uFZKenmY5dIHNsD3xTatz/Nr6E86oPjmpuojedwoLOu4YYM+w360LY
n1c/f43z0JOfkBXgyFf6yUCMduyWIZVGa004gmxr2+1bOmgkxlebSa7ZSER5
MZBP8tuNf0R1o24O6l/vSj9vt461BBpRGgD08g6r/S8GbhRjYa4dem9ainas
8GxFUbXKMzUaAHFFa4f5lkB1AnYZqgMigcH3RyvN78pWYwfWbmcoVKHPp96l
d6EY0DGejjDyzfAtHHt1NglwtblV96M1qYGHVwIuXVY1x9agjvhzPMJu6HI9
3iEHg8DrWD26iTjWP4Y4ukUk9aM13PMU5f7/B7NgckPt5E3fTd950DOaaMib
W8My82YHh5zTi/PatAHy2oPxcGA4/x1QweXGKSLKcC8jn8i88Ps17AT9Pjad
YvdK0pEvsgjkrpCXht+P2VGCkF9br3MaWiZ9yce+hLia4KsS0hCmLd/VyOXf
OEXFuMDq5VlvljwS1ECJXv+4YGhPBabnHMsfw+8MLDJh8FnU3Yb2ryiL6D15
uu8xVz5ldWZCT2kWcP/0Nt2obgLT/idOGny8LTgNs2nvXZAqnekGxFqCWZhP
xX1RAIBFLb8JPNBrI3o5Zy5syO65n9pIA1s4iaM5Xw/wfqqS4iPkTHaO8sqY
MvN0nB35jmyFEzFUQMWrHP7btidlfaEOo1PtUAEx+x/BpxVJ6yXwSiUMLPNI
TKf0a2GRcXa60H6UupqQZaOBCywQaLzsEUDhwwM5AMxZqZln9sxYlvLcDuzV
Xo2H5tPi5dtcS3Cmkg6i4+IaBNB+iad/lP6+Xdf98p7QOaajW0AyhTRRohD3
5KhKNBbgv1VJAFyuZfL3oREUOglSjZ1qTUYFHhImhhaYSAXsR6PF/dKyggyn
Ca2FJS02VV11YwX7ANTiXoUKFlGfp6jav55YpqAVwdDExAQRRm7ob+oqD+S+
/Ip0HRbHa/EAnnCD+QTr2YdeGBzhTLWO3Xw55aSEH2RAq2f9LoAQ/4Nr/+L9
oxMX68x628aThUgLK3iGnTtlzs8lahFjDKV+i5wvmPdo2LvEQlDBDdcmeQCC
VCMgSCbd2a3/QowM0crcno+xXwBhoQiUvnuQwNy6PqcyPka4rPTV07U5ACr9
aZS39x8mTrjJquLq1/Js1xw0d02YeRCKajgJE2XuzpnQVuQBYnpFgRTmuBfc
GB7gejtiJWfD2eHVNU+7cv9LQuhW4lN/gYZtBVss6cowS6LZho+hGy9KUHA3
I4aNrnQl2+BtOK4vMF0qREqZTc30sX0/MmX4S64cpsuJrqTChFD/SgmR+Dre
Z/CBTXsNLUAxxbN9YHSZKyR0kqtFjJax2lV0ZocekALARgZ+fKJbPS8bHl35
kHlwKouxRvgHI4mcGITKlHJFYsK8YcZozv8yWTfzUSSKocjUd4bFNLXgCNCM
c8JkN1TV/1oJzqSq2UJGIapj8FAfiqHw9fflZ4/SIoWDGUeQyvMUVUB0sqbG
A3abJqwnkom1tNfM5MyT+L1w9C6fxvxDqtOjTZVTbhVQmMLuq81niq6bL64Y
WLUqbbUNMUWv/mEHyeoH/bQp4s23y3zn+180DkfXRj8lFkQ9QjTRkqMQX2RQ
dP0mAzI/R4Am3vMU8R7qmHi48WUiKp1o1fsLjcY6iImU72FLDBPPN5VnXOcI
SVTFcb7ji1h1lVh+s34gBBaK0JwtalB//o5YMDiIgZCe03Zf/WyIdFl4E9n3
RY1IErBFsmANAs5aSw8FFDMBCionfUvttxzvR5GjafwIqGNc+y50Um61eu2Q
efQ63CmUk9F/kBnvloTtMKp/w2YNSaZKWoYtJFIaertgWh9bqK3qaFqIsSnf
rAV/5F5MrwNMGf4XBpNVBnMxAx/dyRM0DVZbfm2DUuQC3CprGQFxGGOiVTAu
3jHOP2q3whpTQ3jnDRVokg0ZxMSZkuZOI4N0f551GnBRyRlSdnUOFn9rJ49X
vi8QSJQvK5wvxprhQLRZyJmkJ/PENxxp+oQ5T/+qjNDqvdSjcWaL6VDEvE8O
7rvTR+6NEKEFu1EAnKMXXR7RsKRoKMbPdR9pO4RM/nUjCCSRribk9JMF/I4H
hwFczYu+mLfdymjc6Ez83EgilZjbFdoog9pzwN9P70UuSbaFY6W2Fj7n4cYG
jLX18DlO+lMf4gKmluUhCbV7glimV3Qon2N0/d+remk2C5t6AXy4BC0Ng5KZ
NOZ04DqFSRLVN0ymcvxwH4p13r7DF+FHCBKaQFeSx5efBWXwb7OUwqisaLVs
QQPVKV0jUzFKuWXZShjJcb3hBiG6f53IC/LqldnQkzsXCGPj/sH20NSVkXCr
/tCtyEjpejUVFpEPIaT1GqKAWAIIn20pU+xfV33veI5Nx4tY0mMRaKkgAjcX
a7OhZ+ZjjOU+PcOWzH5jhqNUcU84CUs0q2Qx4VX+RXglw6dw7b1KAvvwIMzF
2eX74Lyv6t7RDv1icenwMIOKCY/sbTaggwbOWJ0rGnlql9kyLRAPRvyNsyUM
BOIGkr++yQSzLUVnXd6WunRXWLUiv7L4/j2r84d0DZLVFd3JgL3pQClNb7Nx
XMXFFwlnhWkfafbz8U1KJo4CeAQ1902XrQJ+oc5AfPjSBJilT9iPEW3d+Tvh
Rm3ShAyUsqk3zV9/SR9f/IF+o8+YbpaFM/NP8223yovbl7N1Q7q/pnedFZqV
wnrCBRho2cl73EBz2l2wub1aU05kj0CGet/DpN0R6ZiERTjUvdd/6I7q2IXP
E8JS2wqS42/bRptl6RZqk1SJcNP2njzTOjof9cVXb7vC+XEbTdueNkB4vjXU
+0iqScoUZbKjNn86QQuz7z86L+DesSlXY4CvNUzHifdkhvvUHXMGsp0PvbV9
B1CG2ahMk3RF9mDjNXEkdDmJ/cvoSjiKzVBRZR+PqWdRv1PQwGGvmtOfoxVa
Yqgcf9vZFSeHKsTssKFPfXHUsGr/xJGPUUvVOWmntHaAg6RA3GbAcmz+FtR3
LUNOtNxOL4a8ONUR19Um37EXMt2LWY+jYlZ9aXOAQbH2k5DUuzkBYqdWndAu
j7g1iHq7IPnxcgtRBnZT2Rg54W9383zd8WnfToPdcTvzuWSvuF/UGiQDr88F
29QILRfBQjEJQVHPWgBvcDWFpAKAeh4KxpyXzS0/ZKMJbUdfFzWW4Adbt/7a
cWreICKGObKdI5scSVe7gfepj/W3sJBQ9x2vguNtHSYbEiip3A8fy9FgnMuL
PsqbBVzJuAnTng+82+5TXLujBVDR8rGhh6ft1NbJltrJqeAngC8OJUpl3D1I
Sq3nmw6vfZOPqFBd+DrzL8wIkWqILaRjeQX5zikI2dULWOOo+6wEjET7sjAf
BeBhQQZNBX4ocVuKD0m5ZNwZ5eWwdncyTo3NMzOYCC1E/RktsrJMO2uduD0+
5t0DVD8B6sb9LOtcxQPaMzUfqwTAcfwvqMmBLumgvpgYI5g4aKnQJcPHR84F
UX0UffWv7ZdLWAS94u6p26VN+2tiKal9HydPuhj0GXFcyelTGtUOibmYxh+g
g/9lMPwcykcOVcrm8vlocPou7UB4Xnp4RspBpbxE9i18UI4+dM9zz+HaBnBM
eXjeFOg3zitvai+YlzwqVCaNVVNIvaaxwrrldqI6eZzF2QgK/tve0Iblp3jV
3r4Urf76/dsOolf07ptt4UeRPYbCbqdHOqqfIMnFUS8RoKo0lHVksT0Lv8Vc
vxKx9DYqnSNVVAF4yp0WzOnzfLx+EiLAtsjP+TGNEK8qr6rDLTHGefGGoar+
a40YS7WdEHHSDNldp9FwZTwl+xc3yh7poEv77rxzjPxOT3FEsWlKGzSl2aTL
FaFr00EDjL0/kkARnNwpkkc+WVEcuJOdtAP+Q/LutE3Xi4x3U+nhpZhwwryG
7L5YNJ/hrIhfrfnFlsaRWBmfkkdKYkhEXresOVFUV8YtK2uhj2KA4mtoUM3J
HXpeYOuLs7L0+PW8kirLjTT3wPAwJF2CPxJ7pvkFvNh8Tp1+g14yY3HwibvS
9gwKzbLpHnmZSTzLlQo+ZXOxUu9svstJxan5A5qlUa3VM35ZynwtHBp8tDZ7
YXufN5s12pQ6DEPLFwQ2xjph7U9nk8wdQQrVV0Qo2Gce2yXKj14DP4Oisjw0
0x8bPdr55woNMqZn/LLbRJm7VeRyiC4IKdnmXPY0POfNFHsO+n7fWrWQDXXM
73l/8xMoQRJx3ybbcXu7vPcU2r8g87KgQlfk7ZE+YRQP7kyZ3dLE4Q3jONus
EX9KrokHQ07dHxJxZY+Wo56OF1hudtDY/KPvQXT0b5bxiSlkONE4uaihwHer
rn1wd7BH41CPhm5JmBcdJ91idepUIGLNwNrmbCrjlGL/UGreDyN6LLg9EUmq
XeB+sfQ0fSJ8I9ZqQgbPcRLaADmc4XC1wx/LYr7s2Nt0hYFkS3gwV1zHkdlp
YIbgVeF7NAwP7yCWvpt5QmRpyt2xVTuajrbyJPiGCq17PcET36XqME0O3jmA
Vtn1VcJ2DDrYdzS82YdDBSSXT4gycpcpFxzg8R/Rmp2516hImqmHa5cYc82Y
dvE3dgAo5vePE72ZoC78TCHjeFFqvD1UViqZHaweTWW607vb99lmzEsMT4yf
mFHPEl+nZI9ExjD8eSvvPKGhINa/lPtmVI8uBhIAffBknE94WKaB3UhnMmck
ypJzvq0jlIg4arg2Q7s1B10ID1ha+iFL9vIkWFngLXm29TPIBrA7nTPWZGuR
YXPVVI4yxJhwN6fz9OCuk2V0u1XG7yPjzU+QexZo6IGP5+ca6oT2SAUkNQY7
mw5GaPIt6zXHR6QhhIH+8jzErpEjiLJ4vGc3qq+9kxkbQxBmGaouwuBSRwon
C0iYh40S0K2gLQq5Sh/R7yKd8p28BqE06F7RWt7UD/dSrjPND7sGs7NJB/gP
A+LTqmn4gq4s6VGPGmAv+U0phfDuBwJvcuP3P38OtqSWEGBfFHQqeZvePT8I
dpmePWSmQnZGFFQwBFZBapN1+amu2zNJaJI9k4mKZcfmo8snAk0UiLMzY5co
nc6u35DZZg5YmAuZWL1btQtUg7QfPHNCxzAzeRk4xamqObaNEkSdjznutN+5
66SWQpAETMQCsFW5k5f547Vf+EkSKiC6J0gu89XtJnkLU7Zjychcw5pAzV0x
TGzTCfDGRhjgXM3yB2/Y1cvLOVrU6UyzSsqmjjbwwpYLQnwyRmTc7YsP3R4W
X3QM8BOqFiVqq6lIpeXT0boxF7IcFQnp6zUnedohJ4TLRYlDM3XORs4GnDiz
x2lUScq8QYTTPOUlG9Ft6PrJHrmkXu3hbPQxwtLTQyRNdth9hnbSRK09c4iH
MH3iITnAU9l5g7V1RMnix2F7+gVxk9PgZ7a02GnM4k3bwMQ7ogfkEWxpL3cT
7PkJuyEYomwP7rwk6kjsubH6Nya0K64/v/68ulH+qcp78QgiLXlwvxfoVC5P
QAxdH7/owCR5CPkyVPRD+YpE/MiB4QCXSA6y4L6MbsPB5HF+EXQzlciL19MR
VNqRZU5ZPk4O1PpER35jZMu23LvGza8I5FJDVRhmRg0UzIoT0S+TO7gYsKw2
R3genBwLD4VN3kvoujqWQuXCjyf9+ZGQhgh+ImkVtQNElwFhF30q2DiYd115
+ouVa+M95g68z7EkBN3SPnSf2uKFlzXUH52JZL9nt7VVbE5bjjQSzyVvAqFo
3Ma0VomLNS4HHc2xyQ4aecrUDPCYnPp6LiWxyXmJYj/bYnalUurY88xLYcWO
S+8IOT1Zw8ivm8G9Zf+zqnw/7IGq52LsyyNWfZFv0LOYK/JecQvpN2JSFMli
gY6hFeocI7mzGlQkJtKBLP/S2v1ELVkhhQPv97k1w4RJJYOHrVMK8lkeealV
pII9WzvsJZ83NaWfJ26wH1CulXWuQ/pW2ErFJ/E2FxxMgPsU3nhF3nxpjYC1
oWUHEKcK8m6OtgrPpESfac16AREzAx5Va/WJCe8OKFW78RqPjs/EElTsR6FN
br+vZoqgev0bagks1E5AKtCtPXI18E8owkRfjeSrtinQBuY6APRCREtHIzyH
0Eru2ovJHW842sH9TDc7cWIQu3sFMQD84hsWQd2vWtaaUxz6306KVvGCG/bL
mkRcHK4+KBTt3OFDAk5omOcGdLfZOSI2o1bXymESnsMPLfL1lHcjVKCVZnFu
4V42Sd7Q1HLR/ybqwPaS17yqeiuzESp3yTxKoYpAJHS5Lzl3ek/ewg2et0h3
L1GFQ4aMZ1Lb2T9nHnSSjqyzYOxCstxVrnNYBYtpwmMIBAv7up+TImKiOTVw
fsA0CjbR2UPVMi/rcLV0E/qYk5C9jMcQtHRcH0+mF2AZ3bw8N7HdVMdHLFqU
KGrqVFnyIRTLJso8ncBDMk+LIz2LA7fssQV+A2sttBeV60aaZKAXM70LtrSL
COmBiipMzLyyTPB0r2q3M9qM58RT+prtVq+XrJXSR1QB7CWxYlzRvOF9EWob
f312QVWeETfBo+ZSlotF/IQkVs/It33aRaW8kQh6RQr9Cf+LuR5P/6pj1WS0
3BX4DY95yHWGaGq7klynjZttV/Er/q1YnRIfnBDFd+xomQlnzVAhDCrC3nH/
29e/ldYz39vB0oNleJIxFJW2f35pW2dJX5NPRofza+5WrOs82wJ5rBErB9cW
ZsROkZfa00qKMzqzChhBLsBzJA8AN+7GXSqei6Y14KKjcnpvlYM3UUM6LtU1
AbDo74SoRn4F6je3H8Zq8AUvJmIcZ4lm3OrB0qofCBkJwXnDgJVQ0OREDJDv
L+/KYyeGDJcPLV+2cb2hLC1DBrWKkTNyAhsEPwP7g0vF1IemVyDW7iAA7Slc
3x8+lgcBGky1oao2Tou/6clhDXGWqJ7k/8P9xtZBHK5PP49ldfRrpnKS1wze
6IELHNrEBpin8Q8WtwIAQ7X2PAdX1ip6SvjelkjZAUHWpymWUe1na0dTsPVn
JSyQoW5Iqhzkfb3k+q/tg2kf8IK+7PvZ0gYxgl/qVPA8gAJWuUpC/0OnsnaE
cFKAUzerOKEev5Z9tHmOmswe1wvXARPFSUtQQj7/N4U8CGu/4jMN4NqueXiJ
twjB2XqmIl2HUpQM0qmyduHA4Sr6sDR9IxzoBNGc/ISYeFI3derFoJ8bnKaa
/3B0ZWr92MkSe4Qnv8S3lVkPcQSt4RYq7dbrzwEI8MBJE5mIdkmiUqndT8I3
7SBULxh6etfEVGXVkreAaYfhVqqBaFmH84GhWwRkJ1x5HzMECmlS35dbCSJH
w3iw4V7pIu24AAoV3/G17+Tjt3rBDCISItNoaxawTj8BEXeRYNmiDqAD1CCk
myYivNNYV2jhBMqsrLHqMg0Z3iKvIYwfLwd/2jjH190HBnmaf6+0RDaX/RaP
y5TMf9rAwFAAMcbdaXYWDPWfoZ9Lp+mxE+SY2pjcNwWmMFiRBTBj0Ff+bboB
sRb6EFEENT5VE1JYAhhbk9fg6KSNQ4ts3/MzqVu9WqwQWzLnJ8VJsgE3F9ih
lpt8CLkZv6j3TDMeQ+JsBXdpXUSu0txX1NO3RGj0P9RmOzoG6cBkYXE6P5PV
m3XblAklJ4S2rCveK2ZF0HpN+0If6mCidqvlofmWX8J8iUdsZHZFgRWF7wMu
x1RDGUFo57hjfmEwH639Mr51tuYfSXaZnCqGhv539CFHWZR2K5UmQcMLEPih
o+iPVOJ/WCRcZdfm9HWL4a+AqKOOogw6Dr8J88TKn9WXfYBIY7pCWj0Czki8
lO+G2QAcTUeFalSFXcm2lF1SnN0whApTFXryIF4dzzTfCOw58gh5fOeTp0Gj
w7w7m2iIrfM69D+/j2l/ZdxdED0VSdMVL2P76DRfRpWnW9RE55CZgYXpnY5b
lEZzVSjRmbVEfa52uxYWpiw5AghI3Gi9uX33JSiSiasLqJyoC+p6S97d2mJV
rUddyg/drzIuHfeB87jNo25SLw72SAtaS7yNIAkQ0UO8kIdDV39IYmhAH7hL
Ql5j/BhrAqgbSN6sz6a8hiZORO8jOduYImELJQkNvhnIoV0M2gKCMb7lqhxG
ygkQkNAlX41saDx39NRuaXi6cLtw37RLqe2KPkrtDESSh7MmnRh6yPzy3JiF
ur9UtAvVeibCHu94KJcLcEFIo3KbAMLVfauR8Bc8bttCtNlNPz847h9GcR8Q
Y/dxdxa7tJgpP2OMlEdkgMU4GYp1PQSIq5j26SKv+UFXibvefhUhsiNLpNQx
w8i4g9Tt7gtQOqPHAkCZfBJRz3oQmGiplN0lfCNoYgY/vPrBjCE1Zpp1mBst
AwY7igaeobyYwwvbNSp9+VW9X4Y5lsQ3aERPZXy4QkM6ghtRe54xkEtIWMbQ
rXXDxyeI9Cg2vCpgax0C+hcTyH/RE436CUVwHLeJJyXX5WiROfsLC5JbW/Px
uooHGGP2Am8NGc7dDOmJYnDsojlrTJknHMw/UA3P77FAQ/YrNtOwdqoFCyV/
jeNBEGvieKKAMDJ7lK6hQfAZlsC445/Wa0D+nl0O/lWle7p+f4/LTXIAqIuQ
KB21g1vj8r7qy1nL98n5xICacZTph8KR336JBSlkm+xDDwt6HKpA4pZ1Ww8M
BY4Oui8cdf/nKssfUJTgdcD60YgEyy+yF9K+AczwRZE+ZUGgK7BON/OeCC9o
vFcYZzdo3Ar97aGgXWl0ddVy/mnosMlljNJTXZlP1XNifzApfnsit3giDjq2
+W+ybd/fusmZlH8PE7VgyROtv7hCT2hiwFkaKzbazMK4TWi0BvgiVDoXf/lV
0/yY3mj3snl+tsPAfuizU683M/uX+yVy7e6NLQjbQILQXLpXr2xr7DWTMxer
/DZSEw4aIw9nrA3QHhwilPBpgUMrofKlk8txe4Q4JDLJZtG3sAJJBAZMZZiU
5Gv/vTBLzhDn1Von8n7ws2VeY8AYTBVZwS/3NoWGB/f8GDT8uVHPV6lYvUI1
XtllWFGTLWs9oZYxoH5ypfv7c5oriRHtbJC+8qag/fd/Far2BUzrMpt8TAHE
Rv34nsBwVAxgqpf7nfUkgOezsNL1fRXKyglCpZN4lOCdyLqoTnJNLpZEwyEI
NnDPH35SYQrk4WL3KXCeQz+NPrYvr/qxZRErckR2A9RCs08+CuAwSPM3vyUA
CZrUd0SLukKWtiDdrRkfWVUGvR1wM2fCGOjwGaZhWJiFdCILJNM+9zJ/GScf
mk/eWdkiMtgXhJV1ndW+5CJ/yGrDKwVdQO5Ou9RBq7WtIIjxP9KURRWGzl2N
4+O1j6qtTfn4OLi9J5+I+6Urf4BpAKXQlfiYt0oAnMO26YxeT46qPqfrU6ZD
wP6Bw7a49WT00HhwPK8MoRINdMCc5lltH0Gvmm9dHpQAcYzJQtD2XMkE/EJB
j4QfpJoqz3JaFEyAxPmTvIV+uxW/zNZTNMdWXO/GaIcukcy9jCOvYljmRNAX
Bx8T3Izt9H62pgWAaG7jYmC71bKp8oQgVydoi4Lhkkp9QvA1o4tAVxNnapaY
LXmO72zVQ0S07W80UzhKMF9HhBoGkVIDGZVVZw2vgO8gV3ANSgBjljZL1o0+
LieFccFqrrLqVuhhwJO2KVAnzz1lNT0fag77HJRiI7Rwj0PbvAi3ttQicMf6
HgIrlLaOnTEDOlHYJ9xuIDMYSwDLRSSz7Q4kteEJ8ITgJAnuRuupeYJ0mOIP
A8AGEKCe+nkiZhsRqPLdM0ATrvwWqgiXpCShDheZNmO7cfu/t+WWtS7gs/xY
lPGX7M5u1qEnjul2QWdJ9xVbTcDDA8rNxwmcCf8Q08FdaIEFY7evBDyI3HAK
U2qLtdWgBt/lc1XHETXioKFYtCYL4gm+F0XRchGKDyaTFXDLkEV9XMKckKfE
pBPAOdCTH3GQkwQnCThRsW+QdY13/W4JzBqc3c7VDOxe4uUugXFYGfhTTT1q
lD1T2R40z60ShLKyuvrPZZPSY8989BhyFU1pKZYoYet1bFHzwacQCqWT60Sa
buACB3rCe9ItMv7HJP7CuH8VBude5pURIaWkB8+LAdX22FT+eVSI+Twm5bwD
TwIZyQvZYeyGHVCEtwr1G6uNwTHu/SDjZykAEGcwccF4PQ0myrnkz4eaRdwc
kGyb1sf+HWhPFlMmMl448kxw/zNiZtELEqqbmSNYNyDAT2CAkSyldr1iTQOX
acjOUvfY0A9HjheLzv5QABaBtGyQLoP6J6LI5iKBwI95tQEDxeNa1BhzFSX7
YXXWxtc7tlPgRwJIOhfW7ZVCQlgP6LkeWHsEssCpvg5QRKl9p5cCETvvdXNg
PvuIMbF1zfiz0LFHPLWejW1JPm5WVcEZdM6OL8UexdAM0G+imPyEYIs+v4dB
OVvQUeQ9+PNt6yzbc68dcu23RLdih6j7tiVJfG988i7+TuKaA4tk2tNpkZ2s
fW1Whu9lPbVS1d/aa7KsFAMJWgTZUvjxPZVdFO4m/OLfNTzTlddMZ1BSPHmp
V2NtjdCqpObVMpKrJh89TE5azxORAyy1+1YVqy0YzQsTeZB2GyNwkNUY1K/R
ADF60uDLhJfoUP2OjWI0JOZNp8v2guC6xr+Om36F7r9XAqBd4RUKZPa/BbNL
AhNcS5r5T+q/t98VBu5FBOIx8+TDjDbhJle2hUX83HcMyKnz4/xxU7xh9HUB
CidOw+iIlKa4xLs5gspbEZVxYvPTmfAgt6dd+JntIBG4LO4+2lT1C0Dho5K6
cJ6o3VQ1fFU8VFhf3RC2iPqKTQcsQ5+2SyoFWyaCQEQ04zLs739xOQ+5NyBi
Yz/GMRAlYZkKcLB5iYTZoiinOrngpeeofFW2guPORLYc1wE9qE3LVhVH9NFT
J/XbWIkuyOr8BXBEdkmbizi/+OCvEqmNfJ/Kno4ND83Ku/D0rfkZ+piC9rkK
dnE3eN6LPeVuAnhWASDvrzQ1I32MfPwWWuWBeVtNQzncik54bmAg7gjCKdyT
AkgS2HEbQnkG61UlAE/GcOr8lWnDiy2aI1E6/US6MbcQtsOBeuItvoC3jkPa
wubZyMWdjx9p57Vu8/rbWk+ub7L3W/Hhto3+2uVf6m6Vn3OW0x8F7NLGyD3o
MV379wiboA0Thg6GctAf/C3mP6l8iGYD36qr4GJNRY3AMYrkC4qYEoqf74c3
wASxbv1YI01A2QwtSj3k0zceC392qcu/4jOYUVdBenuCUQhuGIjeCIkYzoWP
YP64Y/90QyDMwMTvIzohzOyT1uusQQEjxggPXmJsdHEAm6zPulWCyHa/fwv6
X1L60HjB3Tu0rM/5b7er3cj+NICjIk9d5UY45zL9MYXORAo1XfKXVEwKhAub
8HfUVsiN+VeY3lAHaH9VYVmvoqkJ6FfwxMjJ1CN5X9OeIhJqYWsZZb+ezx5L
9qsKzQ5/srYzO5o2lkVlaFEoW9wqQBcfQ/9WL2RjN0swrZDeYhOesYZTckmR
QdyevXUAwt9qBebY5iFabppPikUYcbM8WhXr+DYsrhMylrhExvqYf1FFiiPd
AzXx3z8OVhH3/pxBwc5f627U60J2fKQE0XWzcjJO2hBeFdjbOAzZVWC1xm4E
1A8weC37ZSw9TE63Wb22iZZ+W/8lCYodW1m2JXdHlfQXELZd/ElyRh75SgER
pXbYDgjjQFUiCqZuZSUWgK+EL9HhYYk2YbGdrW5EnX2Vv6joPJRksH7AcDmz
ZMsQn6pxCVd9JxRzwsOCRE6yuRKSJHqH43THagLF/MSudJGz76R8GeFQT67J
W1xx1yUUuy8rMQ3dudJRCXcW8aJQYluc/Guput3iwXO6khQn1BfpbJ8gQYo7
zN+hWnIZS5sre1NWwr1D9HxTCYqbMHlH3Edfz3dGyJ3hsaP1FU2NlmoNruEZ
Bma6vodq8FMbuAKWvBxCfmUxpBiVVJqDqjodypWfoNqmKt7V+z6l1nOPJF42
NR9fOYphzb5X5LWufN2jyxEZwKzuNmfbCzJIb5mQj60aetWIOg8cpnlqrVGd
4rJw3SlFiYfe/oNt7XuHlu3XGTgc/pnwjL/pOtX1vvGuV2BkquViKSdwIbCg
b7BjbTI4iTp5dxyYe76tFqxNvpQinoH2bYWS4fIYJzr0nt7t08pafdkYPQKg
mveC6/sE03aDy3Z2UBDkubGKuxTFJh1tdJVYLn50qR8vm++lBhtU5vzuFuhY
99Sw6jvzigF6fuHGSCG29Uk82N/ZnWM219G/hcFL7OVhPETSmslnjiNXHAsY
KThKDbt9YkpVyzmvhUHhxo1n4hfhoBoepjGc1OAMcUcpejAIE30Ic13dZFU1
7dV1tyKeoHQj2GDRVwBAiUFuDHWEO4WH/eboKn3iziNgAL3tT6iYssziTeJm
ejXWo7tM6H5/6oKSr6UJh1kOp/5IVEEEXaSpM9htA0BDpPAw2RplmIQV0ltK
Zn1/zcAof567tZrhZ90NmMbWPx/tDFmTJgO4K7KlV6nu6oxm666HoM3656u4
Z+FLzSywVKaNwEkE7eJRrfvqFjM2jfUODBCbxUi8X4wYyH1aCeHASkdd7YFC
NgKwSG/6JjspKrNRgvgGFY79+0Ygs5mYh7v7T5BqtR5asGCwT6W5wZi9WmDN
d+vP28qhtxSWLkaX6VKSVdtajdqm8QMUaYrO81cPGemfqH7s5wceeHB8twOl
/N1HbIWsscUXGsfhqohHrat3U5c1n2if2UcMgv4SJEgLQuKCzMCj8Kg4ckzs
DYWq+QjtzpztzehNzfRJCtI+/KgpyNZ9CEk7sloLkiwqqpXXRuFy0FpwbCqh
rXHQ2YYi6HMhrGETP4avlUKTtpPpHQ6ySBYlpvhFOWRgcljb24q2rl6iEglE
5FRCmxybQPlopk6QcmN0vAgFbYGoLCrkQiHsjvHLgyEs9J3Jv7Mis2tRHkLO
Yweba3019zUtfU2qcCHByQLLhNZgMhFtH6zkHiqlzj2xHu/Jd5rq6tf+nUlT
Hw77IYrRaw6uKsmtogdqKG88CyiFB9u8PtD9KZc7H7Kdq8kfcFF5JCfvNHzx
uYawsEyruS39w+QkRR5t3c60VayRzzCtrenAasI1DolyE/GWF1xMheCzA/4F
Mo2oditGEXm7Cr61h8Msb3FkNvXsN4VSRwvhxyqFZci51p0NN1iTBCAwnQLB
XuyuTXVXpTW5/+egQwRc1lk3j/pR1C7GQbe7ilpRTHzyt5tCyrd7pb/MzkyS
NSI2JqSI5adVvn6N4+Ej6VsCfoHVfsZzTh6i2s4pkPRRXOgpu70GCllji33G
MTh9EzW9qBido78sjE18vp4J9FpqsLLdHVdDNmxQCAvl5bXDI21vj/I+H4lW
mcXqrjW/352wlu0ht1LF7o0H+M0hnhfQHuctMbvKJhK3dIud6Shkr+PT8Uf2
i3XhTNSOy3Rdu4KWtfudbybBVkdNDpewU7jlQnHVpU43XuqRLwucxMfzX9iZ
whu1ZA3VwQImm0Hek870Ls9Il5GokaKMjmYJ0DqmUO9SWXghlA6WnvhBzF6v
0GpMiDvrGxhs1dYUbqr0V8RdB/2fAqaW1HmCw3DkYLyzwTQhpAcBeArvN4Cc
Xy9wa7ElEmVIoRJfFg+MDKB4a0AGQR4VS/20mh9z4asHIRqBTYGpd1BVUhhU
xRibWzJMI5V2viLYpiwI3PaCnBij2sPtSl62IEqnbgsOzjelLg50anUB+eQm
pkJEEsCvRgTqV7zF9STMGRWE5yS0QTdeWsWJ+5agZD4fw8/xUumP1WJeoqah
tpG+zkSmPlVM4SA2zZ1Nh0U/I50TXncftV21j4y2JW6fv5KlxbqZGcV1irtT
DBbV9oINKOWK0++812EgQjzv0aYBXYYuGaL8mLbM0FR2rF+YRiiO9oACrCar
lx3j6amjdA/YdK60OOEaxuBlOe0vgfPwsiIl643XASo+PskxsoU6yJf8XbZP
Sxp3Ppk+clwQTstlDwR4u8vgTUaJWGjf2R3GBs6uRRXZrl7yWwqeViqgwICd
PJvHnlgxoDBULMJf28T4KCwXF7NtI0LRFWPvGgbyx/mVbGyXw9cFi/1t6CmS
8EGKom+lzkZIl6OrHWzgIHtjlHy7jFB6+7n0T3N3lLuePeDNjcdhu0vErY0c
RIcvi5UMyKc4TW2kWTAqqOms5iEVOq0eq9pms1EYciA04Xvusx2rx3I76+8o
++z4YSM/gXSALLB3Z+atXwQmu2lvHI5vhhDDRR4HXMdsTZCXUtgzEuoVc55/
jLxYEhY61AWhx2sNthIuGXZgKwoAAXqXR1zl3oNgjP2undBg60GDzbdtcnaW
YUvqryCalzh8/SINRbQbghxUwdT4WlF2wdiD9aKuSahYvDNaEgwp2txn0knC
8zCMlt57LptWiRIj4XLiegY27oonNcjTF0mIMqTZIMkVrbzgk/t1ggeOT6gP
zStVWMDHDlJra/EQTqmBS7Oe4MN2wMrGRwvTuD/FvbYWmtl4Nifv/ktxuSC1
NxyFgEOKwV1iuT+J7MemJZO+OPivJC9pM0COw/j47HBuNwuoSCrWVF5/fC8l
G0zuh6PacszK4DReZ4uv5JaUjexu8M+m4OwQ7B//3HczHPBl4elIWdJll43P
CTAgDyK51Q9o8uOM469lpKwznCDuTWn2E7y+e/ntEV1S22dveOg0jbiUpYAn
MJBc5XV6QYIHPkFajCK0XhtpxKiDVfrO8a5tpHj0CDM8d9QyB3DsWWKTDfKj
0mT0w/3AlWbrq3eF1IdgdeCibTIx5s/UI0ak8NvLQiN9mmxQncnofHmU8nUQ
4PPLGAUlS8IOxLnoxzc7qRUhpR8U8WhYSQU5iyIs7OIqJZop2oclw1TIr5Zy
FsHyKInqksqeaha/pCCgxTOVe/girjgrcKOx/7wI/PPOgBSX006rO2d0Dait
okDPYSNRVadPjQ2JtCgUYDvgJgBVbtJqmiRzz8YX10rFFAdzf/cuSwOLR8sB
A25ieJpejs2gsb4SFwk6reeJFzNxhA+4SEyMaO80JMNjtC1WgG/i5bYp5NsH
SaKq9y0bfW+S3TzArkx6Sgl8gj7BmlOGcskvc87ihX6hanlF5XWrYH/Kbjhl
uUwbUxGCce9KsMZYUUVLsV1HehWb2KdidAlV6rnS+WPi6RFHogO+XsjvlqQR
RdWaZcccKpg/M3QkJrxez2y+hdbLHxdqGt1YQLUZ+55fvydey6ySGs5r6drZ
FElf2Pvipx61guwAuzhrcMqKxaOezwU4/MnF3Vt3FpW0kXcx4uR2sGff3i02
XoeO+2g72DUiu3yI/6x6BJ4w2/Vem++AtdMJAgkMnAt6fvneAKNJQMH9KoWI
9CR+QlKSLIJiKy6VOIpg5ReAAgHtukW91+PQMGocQCQIDBTd65amq1+7HqpV
JT8vrClt/h2Y1h17C2Q/V2dK1cbBnHnUuARMycNkLAlp8vTuakSt5fo3v27c
uigHoEJ9cBgctGD9VUcWh/7c2vKNmiFNXakHWQsLKcZUHKUHIbfi59fE9JaQ
L0b6cfVcwxk/AaWEMpIvAryl8QqO/tdDq8mWw4BQus2iRxg+l4x6fq1AjFp7
3xj7TSZcY6tGWB6uK+lKmG2zK07AMzGPFpt+xJHeZt/smDcc0MV+XrwIO04H
E1iNqFUv7CUpC1XwFxasrkScekcLkqPAIE2D9xZwmOLxJ4DWYXPidtsHljkP
GGqZVVW2idOzixyTjUUukO0ptgz045lYybNuM4cSkF2YqORXDOKD1kMEAzxz
4WdhQaDkKVIiVg88lP9rlxKKrjCD5O6pyRBqdt/o2tT42aQ5jh4BEECDst6u
pYYJuKk3i7nJQgijKuhKq+5lY2rzlBs3LVVBWyR1ALgWi54nlXdah7BEUhdV
3KNol+TjS3reR94tLzJ1j646L/D2fDaYkBT5m7IXBqhz0kF4dGmu2H5gL1dT
g0eNWeOhCwHurPUO2QgK6dv/H1lTNWvuhVErbpWYnpJx0gAhElKDX/LriSeK
Sf5IgLysXiWibUJuXlY2g4Eo92YQ9HjKhs3wa1bldZcbYl9Zbep27K8SieSE
5Ntp9Caq/2IPoT4GsE3NHOdbAIBC5p8zN4GvC8DzbqUwJ5FeUv0KsE9f3Yc+
V/DcKWWOy91u3TGEaXTeUuEpclC3/6AceGOOvGG1Glk0pmGkVoHGrUsGlPUS
bWCe5z4Mq2VJf5xXb1iWeDZ3j6jvbQ4HVPVlwHqVGRphzO/UHxwi4lWABSyV
Tv6gCfErIhOfwgHl/auwoSC/g5eK6/9ltyAh74kdoRuDPiZ89ZLemBHqSUnB
sG1Yy0reQu541sk89xWJgOszY5j6Px2flP/6RQWDMNtjtlmoPd3poG/92YtV
K/3Vybg3Oav3O6KrBZN1+FxpSBpi5WnbvkbL48hu8wN4I/nxqYtbSOyAoP7R
7AKBAuT/uOTbaMcWJnNeB5A0tvspNniQwSwUpBiXV9ZGWvguBqlzMcjJSdLD
YdpUVY+4ezI5qtYLyG2ezJxyepvjz0npOtnZ4ZUDCmvQe4PwJz6cRwFX1rMK
IRanOTTUey3/Bfo6S9/08IwmZoZprwIFRkdrthG2SA0GAnltUiGDmoEkQZXF
+6M7LEBfKfscDfeI2tjXpCcfWQ9UTMv3KSqAzZr+qj+I9uWYvXz2JJsNBkdg
cLJiJ48F147HnBrM3jNFrrWI4EMSj6NSTNDdIDZ3NiUjycKE8FsYFBucpLmf
ocZhxNTDO93ObUVyH+SNEbR+WtllRvcmq8VL6kV/agxCiwiGbl17Chq9uLK+
2NbNNf5uf1y6hMudEkZqWCN7I/RPsqupuoB1E07ykviSeyHyVMb+//PBhION
KApTc/4RS3/6YJXs01fEzYFHOQm3qCQn52GKZwOXPDnyFIhTqbNftJVLx4tn
r/aE0OzLMwQJdddJDdh+iyVnVbL9F9/3w0kco/i0RRNZbXkseAdvc8nLDIzY
AkR91z0gZxvJjVwTEL7AHIih0vZb/825nRazct1PuOIVvYO5BcWvQJwxqrHv
9HhhVmp+vrfXKwaKByOSRWC8jiLd/gsHBWCCGVP+xpsM6TC8/KtkqO6GeQ+r
Jpfz3bIgANvd34h3LxgCHAm7TR3FSL/wSj2Uvi7bEsX4bnw7cmz1bVfTCD2O
JZWATV6dsdbM4v/jprhAZLGqOwqUQ6GD9OVWmjOvoh1iqfDpOsMlWrC0F7Zw
M52WDpg2QgmxFN2PCFVG0zZXrDb0uGFPBiZdesWXU5ady9rS87XToFvK6+U7
u+RB0/dQjFgIdglyHni0gQK5yu+VzUmNAz1ALDOhw4SItobOhNLjeoAJwC5D
lO4NdqGQQg/ar4hjD16A7NLtFiPYIuKWr7FYTs0YgPuk9HkiQav2caBDlFN6
OtsfMwq6XHjVPJaA9WCuAvCgDtzazm3cuftX/C8B2kDCR68lVn+X/WmRP9EX
oOyjW5+Wj5z+Ejco/adaEvGMvSIwhI1v2qdZwYfyodjXdWNVXU31FTklgHz6
Ly9ofR8hUyeQjQpa2symbVs7LNWKDk/d5H7zhnwHJpg9774f/GEi+nq8GI8z
ulHbeBsVkgasJEEVNA5hgmntEoDmintJ352bzOdo8K6B567Q7qYvvVRMJCOs
iYziBAY1Fq8ul2Vh9k3Yn4BSIM+oW/THHJ0eGp7tVd7QyseHVduvzDrqFuD6
99l8VpkyXLnavkn3LHI2vA1mtBIgy2gu7dzoIlwhbwHXXIMCpbQ13b39Jt+B
qwOU8QC6isHNJuAo7tfls6vRZGEEA17btAQQPaPtz7BKjpJVHudQ7JjEt42S
wYJn90Dp4b08CfR1cD83pJore9cSrDUDFLkPhhI8KQQCGD4HPoSLyVjkBUd/
vaKCwoq8wbY39iNV14QDo5NFloOGBe8rxnu/IcZPZ1VNkbwgEsPXY37oVvYR
LxubacHlNsuSMHYWaqB8z/k2NiMmrDKPmSCCU/HlWSAprrA9Pno1GPFZUzCO
+UnirKWcE2rpkmAig0U8iM54Lkdq7iNzm+g0ZpujmE0B1kpZhjAVDOSXxvhK
TYkuOMGlPyE1bQ63mqLyhMiMZrjj4ks3OTGGouWlF77bdMLp5Gy2E3HYJICM
LI6CB5CX3okvJ9kCal53Z0/BSVQLQ30vETD5BXLOkUIJNR37IINlW1euJX2B
wYpNXjd1qOpMBKiLsf3mOe1+PiSn7O05cl0nm4kd19/oc38jkbpEpXaE+ub+
OTBsJPE8He8F784rrX2O21C+z4bg8ZMo7TqvraRUc44FR7CKKkT2jfW2uKZs
QI7EHz8WjlSyWKiM3kbxEst5fqYDtkyUv2Xmj80IGSkSwq1+takyliQAYzjb
/EmHAWFJKLx2pHJ+uR7Lp4K5kUTzs7uhI0XBL0h4T0c5HV/iVQi0+e1vUSZI
/Dd+bvDl1KGaQtslFxzEfkWn28VtEd4Qk3a78L8NK+MfOzVuecm5VSLnJSMB
iE+FbTwn9Ex49v1R1qDzM1HPa+vCDJfiaJNp4OU5wunNwZIDy1dB62UV+qo3
PPz1ZTFv8VLRVfRvDN/yRjdjFLwprO8zNHlBWzRsmi1wzch45mryDKjj+QYm
R5gWnF2oMvrNmCQuZDZMLhPduZh4QXOfCgu2NsUT/X9KIRdCj6P9hLM0ckL6
ayuzPLWB9E0AF+BwC+6rG1eTzv4+YfslDju6ZRgYCLECKwMX38pYeOVkl7Mz
KDFnsYsAjasvrrOcu2i8ZuIiPWzmgB6pSFGZZliQF76vk4reMk3zIjrGEmDB
zI47e4sOTlKzYqLzfDKkddEwhiAIa3mAREx2PYoJ04cfdEPQjlz47xNEYgdx
ouZmG1WUavFpSZf87Lnn0qqN/FHFAmL9onPS1xuVKGtNJEqiud6jZwM7NCP6
JNvNqTp/XPRuAgotJVsEjQD9d7GZpldDxh/XTl4OJIekZmV+AI9Ha5x7A6Bb
ykH6n/LRUaMCM8+098OjNV2fjncjR6kxlmaFcBM1mVRd0huDY6aunxlw48Cd
SU1RmXSse/a9hGC+uHn6POQDIYTpA1Mq+gPB7emw2ajb0qCwFxPq/z1p88uD
OdgpXwg0BNTd7Pv+gcFSHh0UL8EqCp2/FFNStQPpKppjQZriKQF94Cp+tZrK
5gU7oe4Qw13wdP4nkiGYpyj4mOAfVHgguQabgDHsI+lmlYd9HLfvwa9qSIEX
N4CBaSpAu6mfCJT0XXj/nIGu+jBm0AKEU5U5t0u02YIX7AKBmxfyFQB7zXKl
qJ23grgG17TVXCjijc/7EyfYSc5kR3JAX+yPZHiICLEmTnFLXXoC9P04NiOB
JJZHiDrDAZBxUpyIBC5b6n6PDpjuLGiHybMLVzC/JNK5rf/xkYlSzMezjX5f
Y3B69urE4o+2SRdguQhb0dSIAz/29ci93FCO6mA/sKmqAE+U5L3Bdu2ojzJ1
aOmsOpVzxKwdZgO22vYY4Lz4P9k+P34b8UjX/R6gM37tlBRgSJGOd+fu9pn3
dwpC+Ns+0pxiuXsB78an1RDATsaijpbnBemW6UZUrbzj6Pl/mN3QmjmyXNxE
TJQY6dGTve2waHupU2zTDYtvUjYFU1nNM7kd2p7YSoM7T729TSlntWgKrOQW
+G6mCbig2Wbe5yFEQX/tIAD+Dtyh3EqzcagKY/QL3t4q7KQtVCQvBXN0oz8/
59KxoyyIuF29nKIvVMf5CZI5M4ElZ7/k3pjopTN5dW7FFOU2JyqaFBPuFT2k
e7wga3bLu4UKry0W39BwRnlDiEuqSXXq6wd6J/OyABKo8gGtKqgpjISK9Fif
Jg2OrZJPMOBHpBZmiiDuUjPgP/f4xmaz3di6PNO+LHnPrzlucvocHINIVsbF
4QbtGnIEM3AohjDnkxbHyjAbw5aP6MzB3+DAo6l7tTdLH4CBNWmsgffUqcNS
1dPe3QLed46B4hkm7WlWVTDNmDOWeRKLtxBOMwaoyA3gtgEHF4ECLSEE3Imm
JXjTxAxmK5QKmAcK4gTzMWLEhT21RrcveE/0cu1mYuBa7g+/EUZvchWwUpmS
U9n0TUPW0jZkRS1r9UgJwCJh0qVAbvnbx+R40EuVUr+/+Ra2NmEbs+ys+ZzF
VUtnJ7YijVyWzvafZKFR09mjX0TgnW1UV2FYfroaOv2qQlRnXutn9OdPhiwf
4JwOsis2ujDE0iqsUCyf3+gbGIbj1Mia3ly5s5mRtalxvLeZzps4PgALT1jt
5xO+X4R2tKT+3zOZf+PzSVMxeH1yKprPfHfiqDC4PxqK2MDLPaddKCtruGoz
KL58bPVJmjH4wWJugtv0W8EiSuz93XbYWOgYOxXKJYPzB8D1gRloUxu7o2HE
lu7IEoRFmHmOlDWIVQskpactgqTf4YV42bTxmpF/H+xD981pmB9bZWtls5Zl
yFrUh9jIpy78NJirR6gWAdUVn0FCn1ASHJBK+zSsQ/wSpLB0n1ZXBfGhL1Sk
Ka1kXPUFQvBuIC3ZPeZwilSRwqYjdoKy3vuTcwplhua3/Q98NKvN+NAu8GUU
PnSIKD+GbkmsfuGv0V8P6Iy4Wl/6QyUsVU3+g8jdpWijRaTj/s9tiyUTHGoo
3qo1DXfVx7nu3oPuUIu+XzJykwUesQ6gf5J5XeejXRK4v+UlGK4n6VrInlDr
DDraLR374HQXxM2LuL246xKfRQxHdec8tU9R4Zzs00kPsz9/TZ/3a8obLeOZ
LGpoVRLK2zOCd5E5OCTdUOa3zLcRj5Qbf64YmFd5k4OI95tuuCQFD5g/fky6
w7tZ8frPtKvATx1U0WKwE260VDI6azzAk7ju7vRWWnQK8SIRCPSyJy5F0FGR
ooxs4DB9CPb+GeTDw8+7+7S0JOQCU5sVnMxikBWCwf+g/Xx0uWBhCoaQLY0P
Nu66gMkqkIL2HVLvvFIfz9hLdXZ+E/BjsHD6ct5MC7WVgzRY4IUn/aBJpzvl
pfpQZLZ0mmTXjDHszQXyKC7tL+inP+JsZX6GmoqODkU+mPRXwVHsslvwSVqw
j3RpShoYXTahwLN2eCv/qeSjzdh6zWQf5cGrm7N8OJp9XS1tWRy2QhVMokfD
5ACxps4EBvJ0zNC+dgz9/f22bw6nbkiq7op9Mzp/N9Ts0eyP1vn/zAkF2znC
RezCBrTjLM9CEJbmiV3Iahh80s0OssQ8yalyNKGzJYwPSSOn8TrU2ajaLmHa
Vf7gF8Vy9expEXo74ZoQ6KPZPjjgXH1qtdlg+6IIR2mre9+DdI8zBaHKDOxP
J2GWow2iGcgG9hstBmGX/s49hfNWse1z0SklzoYaef8JtM8EEzpkk3TKWCiw
KW+RaNgdtdn6WdJ3uJwBdCZJSOJ+2BLrHTcr3xxj3NekMi18PPyZTy0mhHKf
/GlihbIrQ7LHrJ9V/XoM1XSkQdOfFcaQfIFeJSrR52QZi3NRyw0BmIjGtk57
Y4X0OT6hMTbCauLM/BPotzY+k5VXUU5BT0PTkvUzo8txKCeJmwcZpLwGTyJR
WZpdJ61p2ez4hk3jwAAnLs5cMeAC02YalWJX78Ek7nU1YZ5C8G9EPgCRKBj1
l0AfM2s3tCed2BqFaiROH741CLUe/yF2yVXOUKiEby4caiDv5l68W1yx6xc5
nOhiVURLm4LZ7+04sHbOY0+pjiU0ECefPpxd/VmR02TUhTyQYwfNfdKWqojF
x+9FmYoTeopE/L3l5I5k9dauq4+Eu54BTsT2ymySouzkkKXDGdmfTAn9BejL
YO1Fug8xi7kyS75sNi4EKS6RaFxuxMGQeiM3+rCzS6nkCPVmO38OiDgeu2CD
u0ymDtkngJCSNAHkrxQiUjgJq+IQ4H+wcj2Et5XTeU3fh3sOV1L4u9P2Xz0o
n2D/+2KXfVwodsx+5druIoAQw7cYfHgQDxVxjSDHlmcXbbDSV8vAWCKiCpea
wVFYPhreZ/r3e+K43Fjy89vfHGn0TNhK3oYuty30Pthlnh6xjIizeAkvW4Nn
8KdD1NUbuDcKNZFiMyUrFCXMy+STqD+XdQErqiTZo0MVufzdHqz2ufXaKd+m
COYOBvLu2CLL0xgzbT2onfb+LzWv73/jGdSvd6Qj3s3mtsInpdPrpDdT2+n8
0LUT5VZ7tMwKMn7t8JR9OKDvA8XOHBOOkXaTu3PUBtuars2x0pIx2AMIvqoC
BVDS7ZRVe0XPn0ojUPaXd9dw0Jc/bqKq88JirbKqJ36EV/j7lniWj9af5d8Q
sxVHL44Apl12mEB41Qkxhw6v8M4XjpqDEZwtQVH0Z84NLyl1w11eU6UFagz2
mlrrEgFGNS2SPE8gDz/XLntRF9Hgq3VaQjNmUHfVcJDBULvmK963LW6z34fD
9Za2iwCG+JQwzY9+w3mRYZnb0jsl3KJJ/gVQdnNH+cUc+iKqD0zlbZ34ez6M
/Vn5bREUmJeFk95T+U0WXzT9tqbAx+++VAR2hYWGr7Hx+SGXc6n29fZJCmak
0xo6p4/OlhibuUtM4nUcCZ6P7ui/1kGfHHPL0bCKS01qsWJvXHHLOCVd0Jgf
7UQ5OwSonYhTY1R36iX0s1sM4cybX4CwzCpYdLsMjEK3wpVwUbD2C7HjQJ69
NiA9V/Da1Z594CwI2fwS+ZTRwiZEjIRgtjZc8Fb7t3J2wlMfaJXlzHII1aKp
TCnjRTVoO64Qd3piig5hD2BvkoH+N7nKF334FMjkD0RXCf/TKybZ9nvXm9/T
Dh0FStTcGpKfJtUUJE6dXp05dfZJCIBvA7t0T1bT2uILPo122D5IQARcy++m
YwQSwVsE0GVySrBfMupLwULHDUjHYAs2qeqfiGqg15esiz1/RTCiW6YSZYUo
VkbwshB2vLiqFsydXMoZ2kz0Xe+6PHDbMoFz35ImDqJfJI7R2VZmZ5VAUlKM
Ii47ULjT5WR0HT+NaF7MXhpF4bM5bXHYpf9Ox1CpcqUE4338AQiYaL6gYG6u
OCQ1Hn7IvcfepAUxOdl4erOTvG3tomqbeK9ZrgodfQlfWLsndMbO+o4fjIHW
Do0NsGB5X9EE7rc2eZhQbVlCGCmuE+cbOqT9jZa3JWpKxAdMs1gYmKp5dFkv
rUVhh4CR7AeLkUo2f3UoAuDkNIszUWADMNP0Qw4vIaBHN1wbxNsrZdeCM0Fn
GFPwG+Q7af5GCja2lvEU3GYtPy06JZkbmhFKD+3W6r01QOt5wDHQl8c3dDOb
LsEcwI6Xhk/Phn5ufKue9GgpOBdj7vNJSaCNhnMHcgSqzgcq/qlLgj8MdKoj
iTI4OqlYi+mWvyll+C0wg/QmeSgi/PRASxlbUYRLQ9/IYL2X2mLLG+lB/Deg
6uabPdBvmfttF2zjQM7pdEWb08cwwSeodzOv1kQ3Fz4v4tt9QcjzL/9Gv4Zf
YFk0GWDqnDb1GudKHfVAEr0qTTVe4mau3252WZjL5mIBVO4xqALiC9LyI6UA
LpwOdet8SmhmprObcauy7uSbV/8rG9fK0uNSIufZxc3a4VCYc4qrRz0IpI6g
ownBlddY6FfZwSKC0Yk3KnA77AwzSFLUqtS7elGYKl40fbwW2usoD3LSwMvS
a00mvZTbdRnf6Gqlj5O9JG3hEoLAOO7KAi8mpjxv3G8wvRvQGBPqvTp0TPYt
2H7Q1zFJHrLnTwkvXVAlL2aBpRkDBhppPYJ76YfXIeQxaFkIEp2TIcnsDW8q
WiZDjUhcW+JjbUpNAaHSJA2QkjNsERJqD8ei1NZc5R6lt2Ch5VUTwzukty1k
NrB+9lXreEIYugrDGXfLOWRSXjvR0gvqTg5S+IuaNxMtVYiaVaG0YTrPwFML
9phDoyi+wkTsEcr7fRa7PnibtdrjJUZ17lIUaKARbttHSYTlhgOZ3jTJwF4e
uvgyMaA0g/+xB3PMRnqUC4XQcXaLYIgMGAhGfWd9ao+mx44v2wvNnbEdT/BA
OvDfvHZd6R6DM0GiQdEhlKDa3dfsrSO8Ko646oLt6Q33mdQJL7tnTRpnchs4
BLPcxTbUyt+iS29c9mROGMVa5dO841aNjB4zjo7fluEj32Uglg5zAVHOk2zw
yDCfhR1ZDPCU7HhggTSQGc78Xy1ak8xjvoaGUA7/WuZNdGcHdTbkrTmjIAtw
Ahimot8e7dEK2bUu2In0r4tGBmGN9fmjzM/uE89rs599F7eNIVAuwa5lM+/i
2uLdIscVjBT2r/kntC4WDv7KR8PD1ccOEaVfH3PpvQUth9nOQqVGPYYSNu20
VtNCkpNNVSWL504X3EMjvKs4cRyvW8nny2RvNJej2raIUhzy/gNP+4flAVNG
pg80ApFaJ8s6gSIzEYP6w//mjQGLXRRt02kdyibtbfHIKir78qfHPy2Rgfv2
1evRzo1ijUjDEAKGUSbbH+gBA6kyh+PAsYqsh9phFxIqBhMNAbGIxx8pLduj
aGy3GPhighxTRLuAt9TCqnx93qLLHkMfOQzei4ajaPl4dk4IY6Rv7Q32ndaz
5GRSIkhjdV3N66Un+JYRkE258x7MxoRvrudqbhaqfZOfgGnLrZ4b/hCAELeT
WAJZK45OqREcpWPsLvWXIHq6nGfwxTh8d0WoJ8byoPZSduMdlYEcPLjJjkQh
TfUiJxq81NSINt3G4jBVyUvjjaZ26XukbwXI2dTd9zmLUlM3KQyR4TpPAbT/
VPSQV9aqIBXVrnTGLfWKXFPM5vCTA5HATsISUJWThClB6Slgejvwl0V5DThU
ZdyX22Yb55wH7eIxnYEVnYj06LFbJGdmIUXfJkpx2gyJNoSu9rLjvF2+kTmk
AVw0fiM0t52n2jWtOMq0NGLhI7WzFDBKA51ynzBCOASAhTrCLkRYPSMpyH7/
26IjVmB9Zk+zLYK96gS/lbXvUbnQ7QV8TIs663JNBgXVrjU8uYqAfCAxUz6G
wE7wH0wf8elWR1yeYRM/n4fz/bxGxUzRuIyW7FRg9QryhcvCuwzyJLku4nWg
4W/OxROwqeFshl1z+9u1aOKPGQD/1O7N2NBtiNPQXgs8PAMXeU1WuLmJB0IQ
NuzwJwy+iDnVYMYUrP8Phxzp1fRWolLIR7t7MOReQtxOPSGfQuY4gDV0r9rr
Mimz2V+JO7OgbjD1NFaW3caZVLi6NKoXTOr+J2/+PWItrTDE2nwKt68spSiU
vrDAPpI5biIV7t+dTHrnqQ+5fHrhuhfAGtCOncAL2IBW/IrgIcOCNGpEjviG
nqYi5esApnx5s2wOGjpC6rGXHcWgurkTBG6ffdalbp38CEHwkO32siP0Fuu9
+oKqmu07hLWSlE5tDwJuB3sKeX7qOxnapeBKwOSNSYI4dfl0f5yXB0WnQ53Q
9cfIr1XybXS8x/OHP+sADF1v1TZd0oo/yZS8iyAfESXVpk+MYCrQEN2aKsYA
oNnCjJJO7Y9NuMi5SC8wnxm3iaIbohfRJygATYjbbFZ6e2M2bseImSYFHMVx
/fa29g9hRoZEHrri6C5xiiTEtPlA4jtSlGFijfM/HUbYJix2yePkJ+18U6qM
0ddcLX/mKhdLOr+J1Zv9RJmOIAcCUxYPDtX4B6RvoW+123BNuNpKypeY6a7r
cSe8o+YHBd/gb9L5EqCiGZXNpcChK0lWKfy10otq7dUTUUx46UJn3rk2l3XM
KtiUXYfml/YOiLEaAUB9CkOZXHj5jTXpcAZyj3DI+C4ceoHPu+B77Evk0ztq
aenUaIk2itbm/aOn1a365K7xI8JDu+gh2+vkXNwAhlEQduNe4kxcJwE1SR6h
NlBh3kJTQuESKSPfDzyMM157K0lXJ2EDctOmXtBw05q0idPFVH8IqYwXcdvB
70h7U/noOof7oBU3HX/KbARyky5eMXW3SY7Ur6A41Y+TG4XKVGJuIlG3oGy+
uI8PksiFgbKI9nopsAeF1XQQ1IQ3aI+jsbktbN4lz28OwED/q3+IoFCPx2A7
RvBA8HwJjP+fXxL/Aq6VuXJCzzO7rtFcTYonnitennK74Avu25J9Bm3i/WL+
aMlpLiT22QrpoVjqA3KFsSRzswiw05+mkZXbDgCQ3cuYZA7drFc1l65tE6V6
Gu3/f7u/jWbvpj0HdTt96TIlPLmXcFVaCavEbq4KubV+rBaYybdn09fxTWjC
tI23qAVjEi52/QpEnybo2PiX+Dy9LJaLYbQeoGNTX48gP+NOTQwCa7seAseX
mXhoyA2pH9hakENKme+zQMbWUeDpsz2EumN3nr/IzFtCrAuQ2Tz5NCO3l31r
Bntt+iD/8k3XvSFj+AfNIKdeNZoofgztg+hP+PjXu63dx/FeBXpJTvSJ4Ed6
cGFTZrOSsorh9r16UnqpjYqUT6jE+RAvSNKL1AOCon5qS5sK1pc9iCmwhCQ8
yIOQgY6Bku20uCEIM45NcysNGrUc2GpZy5mVY4gOzBSx5G1YrVBflRBI9r1t
4yGnCXBrfsUCBDU4iMsfDfa2GCQYB5AtgcJpChTSF5tNciiUx1cqkqEXdUfH
NQcHE5aSM8EvDU09t7KVEsmSMt2WR68rWdN0p+IED9yoGr/czbm2eryTgY6V
5LG/bnX0tGQKgXQuV/Bp1I8z2Ub8wLKSuXOOuX1uc30Q3SVHzwId4WdP1sRh
9Z8S9K+UvK+7/nJCFL2F/d/gjDPjgAITP8U4HamQdtf/GnjQlDxeAsNCy7D/
7uwcGzneVIeDujUrfBubxu/Ts5dvUQstFaWWiQ/KwMUoI5q/qxgqqtc3gD7E
JOASAsS0WkeQe6N0R1VgZ37XNDumEIjJJutD0NppTXeMkL3S8JLSvCmvoT2G
P35QXxKMIOcCCJLsy970X5gZDeovkgLH+nGyGzWFWrPo9x5RfyRyjYqngO25
qUiG6lw87cU89tkN1SLU/syO9Il/HSfH9MWIDfxgE7UOt3sSuaIFq6xYitRh
7xBWvxwWmBvOd0i2WsIma5ocaLszBssdPz1ijf+wCpjB8YWEXq60zQHVuR5I
IldaX14D5/gTb/YZ/nlNi7LW7OxOCZZMCdEKNhnH7kGuXtwVtT3lDywb8kCA
rArLO2EpGjJkR+hcCk60ryDKO/n8cPRkpavqYqmP9Kpn2hCBG53KAe53HPL5
6ypfiQ9qcEGHhg9QuEHLUOHETWF4dSFXQzP0nUnu5gjDugC0zSc6mcMkEmp+
8VaUUqcEIpYPkVbW4e/21tOQ6jCakRdREAFMnXWDRY0/eOQdaYZCCcYFMvXz
lQWJ7xHSrlk7Pap3H1en5lOsI4nFRIZDZiq0jnjQA4L0qgy0Y9FwhBRDMvzc
uJzO88KENdz7v2jVLSyUnTQGb7creSMGPgcA1OnSUuRotwwZ4tBuEf2Hj9mN
5XDAeebfrHTkOXVdsWom9Nf+DBG2c643KALXPFJny2dguTCQuM/xEBLTnveP
apbwkGgzt0Z1RA1VePb0QVHIStiKUAHY+WmD4dAOWc0j57y8NmgLHN/QPXSo
S7SJE1D13aIYnB7nZ7U42nhBkGoagYwZfBtndHB0DbEhblne/7ZVQSRB0iPt
Yet7LzgMXZEkCERMQc8KaSJq9xt6nrPZuJF51U2G9SSFlI0/2fyYdREJgEjc
cP7+nJ8S0kR+R2kt+dVvF9fgOb0xbeWL238XusSal/1ttU+4GfU+AnnbtLaH
PlL77wRg2M+qH3NTro53QUZG7EwzKlRdijinCC3kFBwmHmoj/v7hqEAF1lNb
JG0unhlMPjZn8b4HUYukLWJ7gHZibyIlYfhjXSBYmucRyCVO3VJ4VyI3aKfP
x1mWNKayP0MySh9owx+cn95iiW50qcmmtWMLNuXpfaC0pINJU3TfBndHEvRS
JdD0Vgdke51CNwqg4qzQtX1RcWEomy+GdAGAFoWRA5guk4B879fCwLhqwr80
F2bDxCgkTFKqrkxBUKmTt2xnani9DeQBx48WAO3eTJL2h78if9kJ3q+269xg
FRxyY/25T7zKXjYU596e6USptVl1/6F93kzEQl75yvOOeOgxF388rt/P/wJE
gCtPxltnKkxmLl4BIUNYafTZqGgIOqdAJOVawVinXg2h7NKMHSZxoJSpHDMR
w+CF5+ME0RyXisplAXKMTmeMaNGwbuRPb7m9bmhUqYToKxqSIHZ83Wai8SxZ
uPwJwj0oNR0vsEiLBD9+oDTZedyI6NLAWMsPLT5HFki7eUQ2Zc8+1JBsP3Dk
VrXKy+y0EWlm+aZ7vNYVXs/BsXs0yB/2wv2KBDeBnU++td+bpQTaNgLB3FyO
FWOtwF3SIWyY7hmxJ7JsUbxxM7HT05P8EkKnSC7jWoJcVewtOZ+4p70lM5YB
DIQlycXEiJFKEoMGqGEeFD7H5y6CoCLaM4d+73la6kIpu2V7HwyG09WlSWJH
QkPotCjAnQhR6rF7HmW5uvDRDj8Vl3O3BBtQOShQQQsaF4wTx//eBaATb+hF
B1XmK4uggxp4F2xdKkekCqPCQluqLCbaGZFQsed7Xe88wyGSIEPlXTMdU+Yx
KMXTWYThCzeunBH5BZhEbcbD1w8Xc5AiXY+k+zJUqb5hv/7e6xJhEYd3F8/G
G74vA7Ov5fZ5yNON/QrEv/cIBcAf+uojGetx7WxIdaFE4QsQXcx9+ywqjaqT
CeK2u56tr2ou9jDd26GQVOomRoQOyAWnGWpjp/JDlnYn+4fR4ecvqLUJiLQH
Go8J0KNZlbdlIOMUE+Sjomv65RS+5BKbCiZsjTUmJM9cl0fSoqHZFg3g6Xpe
yPEmh8xcgZdsopIHJ8I+/l004w9PgK4a8W9d+QlqgRfPzZzYilgR1xxy6frP
S+o/tXNo7hYLWvXlMuBYqFXycwJg70tMGKGtU0Ylnocis/VZKuKcNCzJRKF+
GTSYh4npc9tJHnLtj9rdLefaACSS1EutsdorRybikTH0qHvxKLnYFI3axu9g
A9FeR/mu1YZchkEPpMCTsC5pRin9rUPt0YXvRlgM1Qq7XUSwl8+f7YqNjBr8
G/5fRqJaYzH7ErC1vQ2mrvGLeczJIIRE8Z61vI9b2njAyeEDQoer922X0z60
Tp+hRL9lQuydZgZeKckx2FB19rSBEVDnJM/3XBTX3fTAojjOsyvAe+uJjTq2
MTmPVr1ac5ij1MRSq7S5Mt3ZI6N1cwftyLMst6US9g/Ymi3Gy1a/ma5NQrSt
Cey9bwv5PoQvbZjnPsgiGV9ApTrsy/cDo6aRl1hRN59/dzkK/bdUOhrl+3Ju
B3ZuzFuPljmFrwwqhd1zD12WOAlEZ7HuSdZV4JNT+fXScSqjNmBa995NYiHo
bJ7UesWIbPacyg84z4gBSVpPHIG/gZv33oQlTBgmuNxt6hjfCsT/N91ra9ch
llKMuj26KgA0DUPwFghYMFtiOsar9Zm+SX1tZ9orBqcftEhJADN6bU6YUF0B
70lxWCuPu9L+iZKpKl+s97L9YI2WHsPqVWc8mR+lgam6+9H0lQWK53kpKmUc
NIqys20K+ksZAfOAnoDTtmhgqbjTYaVMUfHdGtEVeAQ1TXoxUAhCF6SnqsgN
e9eGUx9PfWM24C8E/62jKbEeout0X4sT2Y3suXjeN5dknxBOnxBgQiqmfUrm
U5J19HBtvIS/EvR7hTfdS8Nt1vETtks70iKXUjopmoqoTB8+XQv4vOYs0B/h
S5mMfbbiivaTZvPMbhWgIRPanmVssljN4xejr/P8Oec3kAlQYFSpkTDcMI1i
7QnUdeARpgtmv+Lm9x2L1/kwwO6HyttT64Kub+z2O4dxGEg6dQhjLiCRUYT8
WgIdfn+anQgKD6Vno/wtcz4ltdlUReDWwJjwFtVM3aCP87RHLU0CA4ZL0RSM
J8d9F/MzQ2KLFSTRHZbqW5vjWiphG/c8SmPRH2Mf3ZP9IaYGDOu5IXU7pG6E
G+6jT3SCjvTKXqc+6Qzmz7+pJ0MY89X90HLSTDXDWAtFUmIGk/DRm748cYaK
7Ln+Cf2D6EZYy2Z5H2Xr3J0gBPJ/l4S6ln0eVdkhnfwbIXLBkzr5v8+TVbFw
Lo9/dKgh0b9HXRYsvJe6+b4srtrviR58j3faFKKr5qkvLtb+qZT1iYxMUn5E
wBC9veREYfiItCtFpaAic1YUjWCksnI90MIhWzlnCcN/m6Oc+vNBKoxDKD8Y
fnrFojZfxJcFc71WLHSatEOPRMJsGAj7QSoa0sKUMVfAwDJP1ggT6hNIc3Rp
qe6NQj2navNKIYHJnpk9t4ZuJd07sbQNW/Jd5eAUUJ931O5isnh5fltlGRJZ
6+zS6qG6itvbj48Jjj27XolpRBVecFiTIzqZpO8YfsjKcJq3eDrNM0a7yov3
9P3UTNfGQ9EJmiFqV6pqrtU4m+mqP8iWEPHmuESMjxtj4TojW2awU6TaXzmm
LK/CMKp6yI0OCGiH0ieon+7ZwaKjQeKxMfdLYNBZuJ3f26JFyGDYCYc/gUAg
CVMQJZFRh4+F+7mudRKB4z1w81Ew6RxxIwxvPUtPBWeaUYjJaUJu/5A9960i
/zMIKNyX46OIKjgT9lb2uxMC7vx8sUzifBHgAW+xSy1X/QIH+RzM3t/Hzb8W
XoCfdkjW3vAX8igK402nm9pqzQmErwf8q+l2o+K09l+7eLh9lLX+9VERi8RO
77e4B3cUpYlRYVvUjM7legHYZlGZBAZuUEqpmpZ2U4z3HVzOvapIlYn4zr3A
J4AR4NSHVNE1C8KXfVrkf7yZUcNPZZQpimuzXqSTl0IHQHbmCO86KHUjWXHr
4mbPpfNHzSqtuN7oG5ya+jIj1EmXoys+ax0099wkoXQMfxQk7nY/XfOtZqe9
lACZnwzOTiA3Yro7hL/PCENNFL6bzVsS3pTNiR+2laqIh3iPE1xSwlbX7jH8
EfhMb7qAYEcYF35bQG0PtOyTMtq5H3W8ifweVGG9aSTqtWd7qRwMxY4j9vi9
00cYmAj3LSsi7FZlj7vKGv8vKIqawHx0re2qwYlR4V87XwLevFfnLNhwo+WW
v09wlK/Pg/BGJwXzlvqYRRt0k5ImZwLrBinjSuMD70bNpXgiEI2DFG70hiGP
quYgCy0ze8blojdYvROh8gOyhDq0iHE2gtcdD4tvTnX7l60hluu3DTQKiowS
3d6XrCbaEdry+XR/PA6IAj/qWu9s5969klhT0urRMUGWnSTj7Pu4exVBfG0a
oOYnSUfVGOcCoqsUXH79FrZqOrnuYUqjfO2KbiLrULSgV9kHS1OEb/5MKoPi
D6xjiLbXhbTyaQLn/fJDH0YwAwgBMgSl7lsxWuKiV4sUixJgj4djf2DxYnTN
cxvicFyjpKfvCOokPVKSaZ525HnAz/CycsIf8nR0UURenthLMxchB0PuxbOD
f/q2RcaThpMAlxlEfgQ4SN0iTkoeF2T0T7cns8Kik90rnnxL1VZtLUSZf6+2
pmrJtkWhE8yTEnFx+ciEABM3+WFKUIw1BaP8FrkKIDZAQ5AMzAyiYbXbWMgT
x5NEN5YNtozc2t8CeUAF+dmY8LZxxr0ZFbCINipZ31SjeM3FAwDACbnpExPO
7fgE0yIiiqwJLqeciLxJoDrit7jXzhlcWTl/mfZxF+5sKcC/C5Q7M+4qlcUw
hWSUtS844sycxwd8nxyxtkvGLfcqtO1YLvEHXfRAgJCZJtCY2VC/uzul/DOY
LYTEo+lcymuFUFxcZpBb45W0Eee0ee+1Iak+O1qJ9XHyIbcICn9hdgnQCAfQ
hRFMGerJhaiTSdVX+aAxas4lJITFrY2rwN0Sh2O/03UxGUd0kaR69lPp8FA+
dYNDi/ZWa8jQYY7IagZ9FhoszvnCWSiUtVVTZFJKqGUyNcVPo1TquS/yEGbG
Mikd/0OTj5HpMFTxZxDYo7/C5ysNLVcrW8h7GU0uHUlIEllJezZJ59a/blwz
VSmHk97txGv0SzNQwV09M/bUNHIQjGN/TWqUCc7xDjmQ2GR8ZObzXA85XrWz
3bij0A+1MyVt63cKot3S4nhfYn+L0YjWZV5WTcExE+F3wcQgPPYMdyFFzz7g
Cerg8xsQpeZhrGpsymsVB5DlvcCcmyMQO1dEr02rGFedVakAE5Z2zWo1sbL+
FOJOka42rCPsDj6B+xWjICRxqkifDzUAU9oWVh/mVkdeLKcJ3lvPScw+FWZ+
UKXcYWt64APeGhdTVV7CXEz+72yubM/KxbVuFKftAEqBVFx5yaSeajDKqdWP
wivYYg4ALNpCV85RUmEfSH3jkA4ooHvLp/BiFG65N106xyDEgZVq82xev0sG
FzXTt71iVq0GhUXB65kWGUlza1T3JQs5TOEDqbskbwK7dKfnemAmIZMWnCTK
5X0vaiRbFVcYvRHLK4AgyEuQt3iJh+/6A/wxUgzklwHO/YSweoAClFKyQdzV
ueL4oKgXQiBaO6oR79gTbVImpWownVuVrCqPdI//tHPrKE7MnCMIAhpz7hOW
or5bOp1VbWGnjq+MRpQ1LKqCIdiTaoXt1OBeqpuGWi3MZTuNdePpQKiQohXu
qNZuR2PcBfZjqrtpRk331e+lfWRre/qy5A4/Q57U0ZSoguskEhB4RcofrNyB
m77jYBlamyV5MLc/PNbJeeAlnQieGeuJxnx1gdyeNaBOrJviR4fMFF7I5Q4Q
KKZ9oMP35JmpMNdtTQhemATYSvzLU7vRWdIL/ODOyS0aTZCfQPffstI4P3My
hgLOlQqbutrO3clE/5wVkbNcBx1KY03fEP90qPPD91C3Sjcbix0keJl5BxCq
Ij4EMxIF651zJOPe2TeX/MkJXpSyV7mh3DiW+jzBk3MoCWLSLWBhoCjfqZJh
QC6SO2ruvIV2mZRfNC7XJ+kyye4+9pbr9jJWwJF087dg2sluoDspm3hx2cb1
Bocv37UN87EWzmlypX8BaTSJIEkgsk2xmVPxF4C44WRA0XpjLrtUEw/mmxHq
rYxfE/79kRxzdAXhyJdeAovezXqyKSemgFtc5g1ndGkK+e3jQc3ZCgQEOuU8
TtyjltYJfG80zdZv1UpOTGY6sran/wbhAWA/gUviJssSHA3kkBfHBxnIPwUA
MPMIyQlyFT16MbWlUBZpP43yPpWw6Mtn2/1TF0GtXoOqh0k9b1tnD2cJOsJd
tyUPweb3q0+1dKFEaSKRUNRpnkhSlPMb/+FfpmRAPsThk/dsxVxIse06RTss
L0lcNoQ8vCzjNFb4PvziFu2Ed+pMWbahYbG5JU4ElVf7Fj5crAl65zNdusU9
+47MRxmNpMoDUc+HFtWquJKcLAuN/nHgwcQ78QM6PwP1thL1qxua0HECt2KB
cyT3fGeNvMFE3uvD+R1hb5TTVaZNNS0Me0JaUTQDmXloSDCXteYJ3/jIUtar
ITUeyxKVd7u0DMlKuOV/HF1+kuka2izvrxmNQ0puD2J7KQMS8zUa5DEvY50K
hvybWItPBQqaHszNzC6RFTEDrxk3k52hrMw9yZASA8Ud1VeEoE3W/2+sPpzk
cUkM6MPXO8kwyBaHHBSFPAMmr3hSe2lJTr/QnQJJOd+BrqXe/q27wt9p2ZrC
OeiBgBZxaBLoHCn03JhKd3Vb9b9QG8eOHIlxojBWmMjABRckJ/XrxcVaZOd7
fOSVD0eOFS9v7+OXQ1GESZ/5CvTEbuduXiNUcNE5Jd03EVlR308OAdjZzkgV
/FFkOP+GEMRxGeyVZIYQh1YH5FvinsLaQB3K1q8yYzcjGM7qTkaLt0LlTMLy
IQIQrHTCTTAAWpPmFHHNjm/AXvCcC+oVAGkGHhRELXZsZqQ8xKAHHL5mMzob
+a8mpxUGbLCQCibldQrCNZWZ0mxNJhTh1RbwqjzXMcEWmQczmJ5fvxh4kx7c
4sgRHebvpaRdn0bT2er/+U0M/cdzfBjlC7/xQSw0qwHDLt0qyLM31Ig9mVDH
RnhfWy879aDPuiH63BV//YJMm4D44uSQyDmXlWneJeD2HSWFvYJq1trhx/Ir
lM/GP/YkYmbii/5eqF/l7fAUzTOFRYuHIF9hrvZuEFqxP8V69Hwrbw6s/grV
snNaq9o+LtOQnLpTqoQOl3iJ92SDYptyK35YRZE1bm/Zw34tbZV4O7NJ4pO8
Kh98YKWa+Fk5nq3v1g4hyn1yIaeWkspuC9Bbi+H8U7F4usKKbRH+mDxBRXbN
BY8+oyPn1F49EiQMo3uc6eZexO/oR7wCzJ3YEYUkk+NWE/A3EL0kAoKj+ikU
+d6iCEBEb+eWDu+RB6thLirrhGt7kb1IfiWST6tCpiH9kyGtuNOi4ebDs//U
g298nGHy1XgIjV7YGNs6y/Jlp770A226fRKOF657fxdLrcWpDXOLeS4d8P2X
0ahLSgBtJXtB/bFJ1m8n1qE+rzyubP9HjD4RYCGdwOMpm1K/HuqxLPfEc9X7
DH9C3gqQ5gDMDOmD3q0F0R4cpBYXKzLJOsomi0rxlngs5xGE3Z2h0sMFy2du
9+GG6j6CzHxx8oxFglSXS02yQ4RNae7we5JkBXB5r6iOhfpwv02DDPZuFd1e
y/GvGF2TfonX3iA8KU/TRAedb13wBPQk36dq9FuRyn5vsZn37i6DVTJ2TBU2
KNzakCi5KAlBJcBbR8+oBfnOBG5n5EIwZlrd4W4gjJgUgxI97Wgf6vgLpkzB
07mLqn+gdrxoPmflOLhqlH6DRDFLJD9DLHiVQNFQccTn3yOjiKiG9AQM2QBz
QULVLUcW6Tk9UcYFwANjx8LHNQnMzv9KdxbdtzChoLZRWGd2VekB8l7RMzHZ
G58JBmI5hMukWZuEVfEbPblBDQaI2fgAaVGCGYgp2+wvUM2RlbzwRLzLD5nz
E/yHiM65ayiMo1ml1RGsuNXu5UBfPzrXNVBac5BWtvPW/4KO7/+hBn7eDmcX
XsYJ8hKRovNzNQugPnIrPkM2YEDFSNr3we4hJDNsmCleHVMASbFlcHZpaJl9
Sr0CYEl9dXi1c9P1/y9Q8O2v2mex3r56aWGhayUxVwPweXuazBnjOzOhgLDj
AfsrPC94HtuDrCW3zf0K85BEQUI/GRpDH1DKWzIIRf7R4x9mWXlm/NGvhTHS
GuzxxU6GjWRbq+Szj1kBlOxCu/0psFhNKdboIE0wYCa3qU/9jsyAyS++zJyL
SJ9tbSMjIfTR8axW7KCXBLncWnMZqtRtXDPLBBFp+hK8x4v/YFaO6hyQQDV/
DuNUWCPiyB+PZ8SNqCp8zdIiMY/znO6yyyfTL+kBxdqDluRqckz1LJWi26fZ
bkzIVL3xgu0bmUTyTn9Cbxrxkz8+PghmoyCdN6pw5jl3YaevypRhjNrZbBip
Edk6/1l2d2OUtr/QJi+2+RDsAycyn0kmhL9FqmniMWLerlYJ0BtnYJqNqyvT
yjjXSeSS/iD45+gRzQh6q8Gva+SC6tjMWrxbHVN2srv+/0506Ld6lLzstNqK
gCFCYZ1kbB4uwPCa93iFpCzfIUBu7DAji6+Sjk9TJi7+jji2h3d8sjHvjtg7
4FCzGtRcmbfYap5iVYuu6I/8D0tWzGQwKJLT5iZaNUBxLiwt9vuxgVfbodgH
emXW3o1mLap0ZM3/gixpV52wFXrB4XWRzZlh1MS4PWe3L4QNE2zQXyAat8B/
KFtkqnYe5xijqcGX2jKqQzdfheotb0jQbAKkBuwTdU5hI9TU89LKrlg9mtKd
rVoAeAz3PDY1TUA5yK6vqMmwpj4uEevyNlWhA2MJUfh3tUilSDuqpUDWjrnO
9mrLLP6q1jo6rbhG/lLOo5NTecDkqN/qY0uUah+giKy4ZqkKezz1WRNhubOQ
oJbeOqTN57g9vR3dTcxq7nB9bTJTBn/pHS5iULdyXazfi2oVHe/50exWM57M
uL+Otbrfyy9jCFYuE1qw5f98UIj60kcVV4zFM4mPVUo/swhT3bYVUd58Wxqv
DS1YL7QM2Fqq2RN5n3emuSl8Gk/5KrleATK6IPBUXOKWkzkC+TdN43ZdDRm9
vU+hqfr1i67rQfCXJO5Km+6iooZ+hOcdUJWZrUot22cQRKYIsZioq1MkkWUR
FICNZJjDtGfhWweP5mKs5mALKRZwagksSev24Uj1DDB/ARGhi6tEVasARN6W
qGHTZJniNCtorAmdb6adJXg6HdeV11wyQXNZfX12AUSmPNq3yy+FTAn+9r0B
Z4IGgYb1aAMUi5vALOvV8GpsauWnoPVrlV7LmKIxTrJfdDZ+UUrR3n3ec9GY
Uj+Lzmci3l9V/xk1Ge/HGtviFVJliSNy7poNUYFhhbKNYBlmelzWPUIkvyg8
k72ncaIhbJyGSNWnrH04+Dms+jGajnGsyuJT5VIq+eg+2LA71BPRnrLAaBYT
RRThq5P2ZaFUYkFJ7++yyYs1AsQHUsKqP5DB6++6XiYukBjrJtZSxHUJ9EM8
45d6rkt7j2QODZAHZFt4Mu5UVEb6dK3Cj99zcPxfLEqVdfpDIBItE6Y3BXgT
Yx4CFOc9NA5CmY8Wr6lOTsbvWflS9NCqeXv6nNEizeh7KvHgf7XiTGLRVOb4
uyZwy1ths+3eSM+GBLb9booWt50v1cJMfusqWjlM1q0QAVPyMUiBewYqIMlP
jXkszIVadBilWkfBfG6RwKJVIL9h1G+Lx+E317GefHSoE8BfLkUIJ9C06N0l
mhfrDGxq6XfhzcJiyKRPttFurvwn3Gk5aBkumx9wjg0lNhbvxssSCCG+uygS
NGGTJoXqjkLDG9aeOXB2x/LzbP90+mhRNsfMlJfG8ZwYOW4CCp84D/UfhzKW
LSfEWJVMokuYBZe6kG8fhLfz5HFnNm2rFzBcSVwTe7MZ+3/yQQzA4amcHMlB
rLZAfLhb9J97xxGJiBrqW5CDOap7bwrzLXk2Vt2UcoUR9SWWYW5LFdZdtyeK
s+K5LAyQcSz/IZEkCEcyibhmLJmFR+TfE/2mOiXR3uhKqzLjH3iN717rRyC5
0ClJTgg5/7w8wE4ZgO2zp8mbPVTryZeijSUFhXElHKCDTg5LY60aebIU2w+z
lXmtGlhNZGYXGTHJkn1p7TZM9xk5kTDHgWVlC2Hzo1+mthWXxjKYoOUPLM4Q
i9Ztr1RVZXtryu1//JL68bvP2UY+Gq8+qNwHB9+sqkFfrvG0amPspMkTxH1l
iKJrJUjB9QLHSqvCyhrnF8Jlpeetodukr26+AvOCoZOku1YlR1VN4fe1XlxB
5G4sfxqAV0+f91TU0Yb3yGIj2aYva9pCfL9w0EHhOgiV+56R0D4HxrAAA16r
C3ZrnRyJCpkJXQhnA8uWZ2tr1037cCGw9J+lv17P7Tn9BKBC0Zbt2NrDAz12
V9IP9rpy1bwpaEg2yQXrg6a8rqoSm4tNcBXDy/fO8YBKH3W9DDqmdmAp6DZq
Xpu6I/04bZsureps6eliK37QKAZn3DN9lO63wgSqEEZatisXLNW/IxTIyo8c
PONj7IrHAsdTWkzWz3uSN66X56mxfrI/f/QJsW40vVjAFwTHZZRsdzS7OS6d
X4NFINoKt8IfPwnEZ49oNon8ZzKNpcYDBJk3HuZj5XVx2O4ZWQALaNabiJxh
3Hue6NIjzThKF6rtbpqG8TuFbtHQheChprDSp8BwmbscMB92iQaIOJDYq2LY
x7OSL11T3/FkG7B3YKQ7jQiZWBVhARdo38Jg3AxvUWbeOB/U5gOExb+g2Z4L
5lfgeVnD6y9YtToaRutbOfT2vqFlQ2YtacWeRL+YFfC7D2E/13jygsLgS8Dv
kuiAvogWi4nvosXsYpixiGESNjfCscLOhTdvLQ4YL/sxgsSSvWbWWMI7c5Qv
PsqqEpmempDH5bLswh9I/TRYkJQoVzinmjqtGn2+PI0riUcWfEJN/3qWmSCB
mSz9KBj3fsL5SNBGMiz6pT7w8BligrhNM0EVLn6W1WQeoSUTk/iNpCyAc4Cn
xmd7sjSXHXJJ7kD3HGgF3l4xZgHnx7j9bjquw8mcT5b9eJdyHcDRy7n3lXMR
gCEfF/W/5k1Oe+1GjhevgiHrtD2+zHqS8avhSdJdeG4q+ubmZOv467Iun6KS
piNqLV3TUzcrbtaHSw5dwoNnMIeP2dnt8UvyG4UG4m0FBAAkIr6G2yI0YJWS
U3fHt8gnLLfdb6YSy5GbZlDHpB3cvFwse0up1wXKGhS2kHQe24E6J3d3w4WN
MA2aPDcNxGrAHDPVfk2dAdvubycYUTMYBx0QR70il+C3q29e5249D5ndw+Aj
gs+kkn0SqNCSd/ZOXpe267lXxkM12ESapc+00+gw92FmZ4/hc9EP/o6mDeCe
CCU/XE3NlNLXq6UkIKXTr/NhB/FoJiXC3yUCCPo0ISMUK79L3rmFwFKR4+xw
A6tzr6OhzhvZOaUtXlTdAK0o66MXOYZHYtYXOyeR4jS5vaSSJVgtWaQx6mUr
ZeFsoInS8GsoXAebIikzty3N0Kvd4nf7hcPYxESorafZEZ938DjH3g7iUlDy
OQ/J+nBWsQ3msLVDbX2Fy8oBXs8ujY2SxEkX451xKztUxPx5gW9nVno/MBml
k4xKAR68Fe/DgdTKG1Z+wSNggS1WamOlaOcuzkhV8Y4Zn/pWsjMDIPZxkOey
hE+BIW1ZTvW5tEJrxUNoWZ+1X3thfg2mLsMMedi/BDEaN2GbQPa1BfHVyi0y
QpLM3CCj0RRW/VGyBNL79DJxQnnGXJ4lrL6LTbwxd3AFEPJgEi6cGSTLYBST
oTQqdGMCui9B7MmaF+F2hIbhBW5rYyqq82cx0Yir+OoB7IuZ0I34cTA1BFit
fgzVDXktBI/0aYHoytf4MUT8yVNnm+D25ec+wa2Tiszf6k+cFob9k++pbUro
yQlvPH6/cjxTu686IkH3JnK/Yu3jzc25gr/GVeeVk+R4cXngdSpsg/LOa1Vf
uqcVwhTyEHezm83IbTvAAy4YgGzVRBV19PS45VrBIuphSeAzMrhZ31qnNk6D
679DCqxXqySAufVDTQP13oM/SXMJiCgU+Fadjzfgyou6pSFDNN842fCNDME3
VzcS+plSNnHTQMv1uf79xccwWkBMl0DOWYSYXJliAY0AURKKXCOXWWLAUr48
WGr+sFNZSTiSt3q+bCKpBcO7d27WzKjdegBPN85UZRbOdyjMSGVQVC9QWZ3Z
IIC55FamgKcIhQqvgSAj0Kbnv42IjoPyDKQJoAOVf3kewCa6KWgIPpiLzqQM
wGi6/24LAB9XRqvWJuaDFozccYekW6xjH3Qzc8FWxQY8X/LqK9x2xs1n70E+
UiiOJEaB2yGR1v34zVzXfKEH3I2cWtMPJ9kxIjZxSEWkLTGHTJxWweqZHwh6
Qsl16HNIpZyUi/ZQBNpEdfoJHhVs0/t/gGtHJkvl7RLZAFvx1KVqig+2OnoS
GFsHUNEeovPa+x0DMbM1TyJgh7brcDRclddI3plBF4ay4okUQqc+j6etDhj0
8j+Y43+N2rKemWxLVSty5xuU1Q32nw9Q/Eds6+iaR6hJw+FpXFLVftJK7VnI
HKYWEU+fcl4xO7ecBN6WfzVCDWx8xsAsepVZtXRL29JNOXabuxB17s846A/Z
ycQIU2/udcxt1mnBm8z7WwdxUwohaHYKggfPQjR0rsaOhtue7jvUoKEN9Ap8
gIsJhmPrTcpg9FnYXtdpasVS5+WATfzI2kCpLuHkYeM08eH1W4N4oUlxgyEr
HHlwfkj1g0H5GuhPJmhxxggQRovCevH5cYJmX9/Y34f3HXhTJjZyKPjD8RT5
d8z5QEOBL/FRlomsxsBH0AbP/BHTkzhmpUGlOCPU0DhtmQwT1RvSAZv5Mnap
Fw7mRA5F6sZf9/eHWNlNjbIHDetKQpyK2e15asFO5eNzwLp07z+qvyyiohtA
/SvDmCz/ZBU8tVvG+ubjiZDJ6/L6yHWNPL5xQBnubN2zI6GZI/Pp5mM3PGEt
71j1bSVX017OLm+WKBgjqyJZm0v6SzEyo4YcCfXt8fhQvKF9jjY0Im3g1BKH
2LT24X+giHxyJf1F9tNmmF+u0c9ohGN4jW0xayMPUXQ4hqaS1rUYT3ediZZf
1sa/NDsG6w5N9Z3ChZ5lXZ2n3cSwRSC6B4YNhk/Dk6rHr8+/ZrEPZqx6vTPL
2XC6MSw8i0W8aodSLLy5oxZQltfLvOWy2mpAj+mW/48FmPzGRqYulfrEHSMc
8rugsYLICep1qfAOIyoUdSya433TklATen0Q/HQzYyXr/xM+EGzJa/KWuw8S
lxvIiPlOHPgtW9zMhN2OVjZYeu4SW5sgimQekJkArbUzKLW1yxFlosBHAmPz
1sMxnIdYvbvKOo210BEycbpEVXhaJe0dSsgVYxWVPqVlPIiEY3XNyW7CCXM2
cvL03Lk6TP6G59fwFrHLnv0myToTcaCeKpyd+LvS39IsEZhTBDNTHb/W6dP4
/0x6BJDh9q+Frt+Ectf4iDviiWTog0V+S5mxOwn7mkUEzenFYwn2LMD3OFyW
pSWZV+dvF/LFKMT4gGc0ciXSB8mz8i2Vf6TdhqBUiWW/JxjWM7R/twm7vuUd
hIakbcbwOFqW0dGcSGnKvRUyMnIwXu/g2BIYIgOuvZUT77DpD/eRF0L4Fs1K
ncfNL8SFOT0DMrO4z21bxreP2LG3Fl5WjF43eFjefuLLoGgylKFwsgj/dmSf
f/09D5XZc5Yt4xs+bfYL26Dpqwlw+ZUwKv/j5axOENRnDJ4M/P+T7nF6XL9u
BgoE9d+BXVyQ/R56oFkXUoM8MsMBtLIkHpZn/Eh5SaQJuTZeT+7Vb12WbEaS
LDxT8Q4NDGAz1Dxd3kkHs8KbfwDxGWL6FiV+zpWB4Af4lSl0J9ItsawSqKHW
A6w5YUXZLiKvc6FoRBVb9RHK1HB3en6ycE/abYTyrg7KtlzFW2qbiZFPdcE9
lbFX+kYcx+oxxr0NToBFwQt5ZF+q5CKIOC1Kn0eg2RkG5AsjmH8MF+23/MtM
eLRwhthNU2eJU9VNM3CtcEhNocjm6I1KcDLboPzxJXtlUYsGfBf1bGo4vICT
bw+HQEyGFLJLNrXYxpSOsIndaYCX/uVQO0ZT7mULsgGaMqwYuo4rCyrUy/gY
/Sh2FCcopy+kiDbVy8ibuKoJn3hOPvo9ELIVoGPPEL1xKdBho+TIyBZZuumX
MYCuUljd8hv+YKQMaQzDsDmgQ+OBVoCEqkw/fa0wBuBJ2NDTaxkmVaS3Awyr
nK0sPvKYmjOz7rmSTvmL8a4Zj9VhK7vkm11uaJA+scBq0iBfvTwjfLF8NmvA
kBNsJ7PaWvF9nBopaWvTgE5YzzupzUG8AuPYo94h1QGbXwtgJQztlwQcWzB7
w+zWjIn1Mo4VUR+j6qn1JkcVqkeAh5GgmHAz8lgYS9imtU6D76i1sVf113pv
99La2epFWm5opTeEicBWI+DzU1eqDakgh9tZg72DepmyMsyUN/90I6iaFrSp
DZUnuPp+1hFA3WiPMZVEbF8hl9l44Z6tcHNtDu8PD1yF3FNb5uDehPxbxScM
nfLIGHzwo44xynWgG1Z1D0Kk2jrDJ2bfwU1LfPYoxO6Es0i1dQ+utvxrUjBw
2qaot+XA/F4nAHpynaw2+gMo0QKJZwavNbK0W/0pDGkUNETugj9FrxxZ0d+8
7JDViN3Tk64B4mTi7UNl5g1SZHOUnTbRU9dXguT3Cr8npXB8kDDqD8k6yLtF
DYFBQDT17pbUj5TBvMUfHGHsdZf2WPRIYTPFCQVHT/SER3ly3jjM0qgFZ1xl
dWsGQJzGDWBtHdXWN2VusQbOcRd6tliOCAJn9mU7QjIJN8AIdBo9J/cG6Dak
YNSoV8vtWmfuV9nqlbBvmhZx0RsUDEwn6ezfc/MyL6F7sZbkwnkw2QoG7EyL
JGASRcldcGXtvXcZLpX3LVDLM4q68RDPhH6ZluTGmcky3cCgS6kNRMX68xJ9
FtGXS7DTjxQ4M+BzGNq6JzFJzmEzXcS79tRBzzvF1rfRaYLxsQ8LEhst+qAr
O9b9YOWi8qebx8FD356e2398sCK0YdlHfU9aHJs/+0NI4Ao6Ajn7UVCpJ+OR
SU0fwej+82n1NvpPBjcGCuWRyehWoimVfcwk/CqlQr3GWT6sCFsRjqttO9GV
i+Ij0Mfbwxq5Y4Uxdy47uQk4wxctU9nQ+VfnMJY/NaBKooONa4TI9KcYREZE
IwZb/VfdtNX/jBMsDoR9E4Mz/Nl7GmmDX7J68FseLjDOM08dReQ8+wPtkNck
jgdo3KeptYgudG7TEg9nGMu+Ot08eMQBry1fJyuBsksJPqEWA7U0xHhGWWff
iIp/l2M96ge68iW8LnKoR6FXvGNqvhkrnKViZje0mwUt4aeKqQQ3nAdRuJMl
6igaPKF5xIn2nuFmUEIdbC3ITK8//QQFkaureCQ+8RWABFzMIx/BCtdhAyMs
joxn8jFToplU2VRsd3KNTuexXXHm8YZiTrBALQzJRX0E3HNM5Qx9LViWTKRz
KvMQdniCsyGEEDIO5wmL1qQCATg5wMWww2TVvwnXVnq/pNoAjeiVebgvCovm
A/iOVrULC+4nMMh+ZxhNKIq5udp63i9QiYXygzJ7vqnWOc8rqRePwk9KxtTJ
f2SQznH0DLybXa27yunaxXNC+jDZ5JzRMYyTZ9uqSBIzn+HdVTxrDl8QZjGk
G2+X1sixVwAIVWt4RoarkZTWcDCM+L35xaH9J6A+k1F8fZCYh3z2m4vh2DtR
8xiTpdQQYFnzS8sUNCyX1B2Zckiths+9SjCJqQ1psomBqRBnNQNV8vQbSk+c
Le5VpcsayRYqsOjfSS8G/hcCf+WaR5tpFK4CXJ8AJPMD76zjv/zUAD0hr9f+
JiqPveA1lsLz1hPol2EmeFu/bB2/NRkT0zxQvIQEanPmJiEtcVKqLJMdiCjn
tvhhXpXo3z/6IVOIkzuTl6TA4GmgtMKnSmXe2ZBpuBPMArMxXq++WiJzoFkx
kEbELXwBr8xVIgvZycrVvKjE2D4jGHWayElYR58LnFFALlbDYK9GVys1L/mx
6bm3nlSM7JvDQ2Gma8fE9RfYyY7J3OvW+z/zcSim4TJMWhcXzSNY+nkCqMY3
Kbzi5ryxUdbvvTX1Wxj6LtFwHmBmyJTZds8VEWXbhD/y0X+61NA4GsmewX3s
9Mi2s5odXee3FkOKQBlaBXeeiEUVXRSS9JRiIPKlV3ElGgVVyvhtsuY0H3ue
3nnNVILUJXqPP4CpVf/9TtddwdNIW7ZzRkQ0MReHCcihizjkDz8FJOMXJuM5
WD/yZxo9d7aYeqo6OoKuoM8bdC6O6g7Dw9+yjcPDqSfPvfexEjervYkD/5d+
HN/k5h/SCIkjqNj+unWxWXX7TC9biXH6pQqj3bhWLroKN1jLEJDwCrgVI4Eo
o1pCXaPsPmbceilU97yP85XoC2p6jM61w4Fx2xGuf3gTDGddr8g7QGbSAAzB
mLLeW81LmVknbG7HxQ9clcQO0Mi7lZqZDVKmxk6jP5q5v262S0s0VTn6smvx
ocqhKuXherhj00EwLeii+fkYgRMgcTsgIN0tjwV1rr8gow0ZcAwgvrp8BzwW
Ux2knwi6L0PSp1qObH8+Hbrm3WSMORJeQx86xBB2N/hzI7+Vy5EsLsWntfd4
m7fLk39l1EyjLjEM//zzogOOBW1X2qxkbR7KpoL37M1pv/7e/GpwUG21GzP/
kHaoYw8c3Vm6QneHpj8axe3jqhe8bKeGZ3n3aplld8QysgXYsPXYmcNStSqO
5IA44vKWtovbe8YMaahcsrCi1j3pcWC7eRkXaqQFrmXfOyVufrjlMRm9bdJK
bKz1JYmAr5n4UgwGrSKphpJfHXeTGv9bqRXOuI0kI1ycyEXBUuYa6Jj4f6eT
xfsQzul4bByTZ6INX/BI9SSuD2GRQ+sCWDHv5dSYHAdlOqGirEi1Ck6dcjDV
hrHmhXeZcG6QRoIZoZq/Jfrh4wK43nRMyfN54pUbP9WQsdREfekZTSkmcfqC
EavOjQejjYQuxOoFzmyeGP1hNY1ScAW6GUQT5jIMvcWofzRt+ISA23h01Tc3
E2GRYCPbloE1kU/c0UnAk4ksq4+ZF78ZZHOCHpmaQ/JxtPurRCcM2JH8isH/
7iq+WZQDvOF3OBrnVY0mMaKFa1VhKEmwg5M95r1Rnv2M5t5YHrAYw7pHHnZn
sOpO3oEI1kcRSNGAP0CdQEGD2vZxNyBekwOzXHmMR5OjaukzJl73tqdq1RMd
pLL99RwiCj/ahU5uBv9KDm9+Im50fe1Fo6gO2hxXcG+d6EvUJWaVSciRfTIY
mCfe3XumBSMnJr6rLU/eo4/n+NuKyDLK2ZjQN/d8+arPfFXrdT3Yg0y4n/p2
Da1GMe/UcNsteAxJTyQ2brQeoMlPQCg+YhRfttsx9ya28e4MiJ+KWgeuQLSw
YLN+gEp2m8mATjsls9MbVCsVdUBc7f2JYTIuR9Nf1SLmmiafGP1zcnp2M9l+
peRUWxxlDN9DezldIlzOl+JeNbtVpwH3deeDgfYdmVEsscplKVvWtbeGZCfQ
wJoox9Q7AOpUIK3oUeC/9PROsk4CK8qokABjdtZenWXOubg0KjbAPcuXLNA3
0O1fSOtj65uIaLC8kmoZIijdafH1yzu1O5Mevi6kY6zTxq32tH77l3e7BhIK
47kiVJLiiWbRJXlRVGEZVgjr2sQLmrdPnWlJ258tv6UzjZNN83v+eW65fP+D
lIn5yESD2bDWqC6K2oSHPHcnPAr8pRVwlpAzP0nhXajjzRprMhRh2995a8jf
5fX0vcGOdYZHxfPSzQG9dVyx28OKLoLhtX4qhCAj/s2/s320Sw2Kro4Phz51
fR3xdksyQk4HFsGgeTdah4euAxw2GM39XDX9mwN7EuPpSsk2ZEth3ExVoPAo
PRjEo0GjYv1iF6me6eVztrNiZdZF8jBZgdtABSpKLIoWS7xe607jcW6hoKB8
mFCwSR8r7fKFQXgGoeEEBXL4Rn6BZzkdKYhKD1ky0xt7wY+7lWKz+iIzmcdI
2G/vvYvli4wXMY/Qhh4VIDJ4wCmJIZoRaToDWOTk3lHI/17welcC+ZoLtWXU
wHRrAgqM1WlKnLLecsc4On1aUHzCSK9+6drdKPXBEjQjc/laWSY3cheEyJFH
C8bIWHdK0KZnAqgQW3syOXamHd6UXyCUkN49NTGJL1Jjem5Raq6cCJm8LsTQ
0F2kFyA14NHSZ1t4lRhj1dYLjJZFIiq330G5MkQ7HHqy7Cx+w3CMt1dB+9/X
7I3EIYpCZCWESvBJHYpyBVlhqDSAcFDisCzGDC07Guo5RAhN4peNBh1VHGKS
dTaGpwH1/Rbpo27Mt4z45y3wJhx0hyddyk6VHlX8KZkTI5ojPkqykOZxsPzG
tWIU8zIfV+NcCxbj+zE8Xg2oOZiUd4Y2y/IRh3PYQDhlwbntD9roijgk2Hcc
VI+Z1l3hQ2Q50ThnjfonayC8YDV/9i12WmweYKsNGhpVDrLGkpZjm/FZNfdJ
O9EMz0Cyds63xMll4eGPTKsbWHbgmn9fzL95/eezMov1CCv65gCuAyd4Of3y
bbq2PjkUNICl+dU8Al8L2eAGaF1mzRBuQsZKpdqp10KKAWidJtZ1hqpd6/0S
U2dQdXbxPS9AcWGo7q1OFhazs/SobhyRAPNz/ku2lhaOUObPstsOBuuvFCoX
yHyJmDbn0VbxihVIemw10Mn9GjHgMNOn6tHPHxL7rG3mTIMyh/WHuiZDOlGr
M1g49S3oli0dj88UoVT2p2fgj62BPVAUBKQQ8wrYkZSzwWxV/VQvOIgy4LWj
9WgvM0y99A/8BzdD97bQOuV0t8woRC5ahJgK97ng3oHJgrNZgYRVmRavXoCq
5SSwzNZtc3DHYtenO8Phmo8JjnQBT0BJlGQpgk/7Zmt6s8NPWQqRI5EIndHs
8BtjsHMfJjbnlbvd/QqJ92nmCydQWiNLE1el+bY97I/1a6cgtSODjPgvOvgw
lxifheeq13OQNWKIu8VeyybYkJtK8oqYNbqfw0S1GecS9Y3bzdd7haJHoHtC
bcRJg5c0QEc7/wAEsJy6DJgde9JuZdAsBNKXQW578CEbrZFvBY1hV8X/64S7
Lvy4WnjyObif/aJ3vWleTS8iWMeln8AWwItVbK0Cqeq7CW2ADl5rdkdQuHQT
YdoKA+qYapK82NJCyZtH0EA3xLgqIvWokK2C1pbaJuiRDxFg20zELegbmTRz
MynnDAotvfryQa4vGi8aqEWyi3stUzTShq1X5rJX6tUinFURo07Klo2zfXKq
VKloI23X/zf549fcy1vuaj3cXskVZ5y131MrRloHQCMfOHc3dxNgKXCCkyzG
32jDm9IzQAkbP3Rqe4Dqfx57TwNKQbQQ4TZv03tAfE9uoKy6tq3hUcEALs/O
Q64E3toHq4a2gOYQruuOAVgyPzNxoI7AgEXldMo41EgL1FieOFpG53hPzteq
jNKiwLg4088BpvYpYfQL4mBJ3HwArwmUAAdcRkkiBUScvpY0YWGtkbvBa7lp
vDrnbsDDa9X9fj+yMfiGtkVF3PK0F50MSBjx194zZxhjEkbCmxkbtN35nwcv
zlq2A5QQfci2g1hn/Dmcr1rjQMP7LdgqmoneTlxXSN2AgGuxsDfMWuJINyL0
Nt0I4BAygu4p4CGQFFm1OV0bFD+ekps9q39YmTvaOFWCR43aqro4Jxjgtf0x
XzQVDszx+jhTTLaLx1EzhXtl/OGcBHDBkvey07KrewW2usPKlbVix+icYGDP
sBR1fXeZ3bhmWC/V5QPWsX9iwR0tuOzl9BU/IIFY/Xe7pmlCmLuJ1yG2sCoq
tmAGgK1kS85Mdqv1FWWWKU5fmIR3jqLW29gAYVkiaCL5su7Lp3rBJ2TO6dif
Y4GLY1dHt9r+ioAI4PaBvWpTUezWGHsiJ9ohXCiC43a5PDKLNWfECKeST7nB
MhPZxrEI3f6nR16gOVII08UZP8xPGXtZlX8NhvKjBt5DUEoGquj+G6/tNIam
MapXf90TjIrn3e1y3aIkEmw1VgdRXlL/XrMs3ZF+yU1dKDldICTk4qUmW7i+
ZJjK1XwPVyx1pjaW6liWOI8/haswYq4zVR/5x3X6+uIaYKFoY7SxGRAEDNQ8
8ff+m6Y8OqK/fFK9I8bDpIKpEzQ1eO58UC3mtygKpVFvJJTTLStosV2flgW5
hzLYTRb0uEQojSfovfR3AHXgHeva2lrrgI1O5hWMzOe7olRxzBqnwieTt1fQ
WDeU1pmeIUchIASf/OcESs+myFnw0dwPWiTqLpy1zPlBcHZua0B9paehU9mg
Z5GJQHJlu7w9Xog0JZEixW3rnbhFzH42xMiEzw2mPoQqTT5ubPGiFJ0TzaGg
q/zGKNT18Ok99p0ibLjld81IhBotF57eTbGAEHSa705gRZ3XGDvwmhf17uUk
z5LBpiPPcgttm8gVBVCrjydJOBxPceOhHvEg/ppUQZvugZXgxrbrkQ/8Exs2
PgUzVfIN8lxRrt7ajmYEglcC9U0nImu2l2LIIOXMv9iriDiaThzDKKtALFEu
sS1RXrh0JtuTbcNkQ2hwhjUGn6RtYpMzwYRIv6F0tJb+LcGNFhc+84SLAPwv
EDacBhT045InWiCcADzF+IrZSoQdOr71fCt1VuufF+bIfkT9HgNVULEDh3Vk
f0D3THCFwkF4vtND9Eypa64cHzgQikf6cUJTX7ptRQE5s6vy4dW8DerK1kQ1
XQFyMNDBWIyiDWAXUqfFKO2uNb2umOHNIGzquVJX1sOx/iHrxLZtS8jCrfso
ApBeX1uq3gHJraI7ya8fbgE6IC1Sa9u1YvgYraLd9Q/I4LxWDphge9oEt4UA
1mI7nYrT+dtOTUt7naHnf+geMy7pblJqskg0//By1bJc2ayKe1dWVYLh84Ii
otCcC8n4/US2CUMR9KgPlNqbkb4pvo0Obz/2PpP3qj7wnXDh3xP+VH5T7slr
uLEebwqlDTaS94UNyZo12FwNjONx1HrvuzqGLW2XxVuRCDkKmjA15x/ROsvr
IEaclesiycUX9mj9u/Sfhzm8x+lW8yy/8eJTaMRbP53wuubZHudnamJM7MLP
BizX3nZjvViPGyVYx4mIqp3hdVX1CfN3pkHNephnc0tL+8mh6H9QjvJ1ONLp
y1Bu536EGnw74lmWz7U7WWyypCjW/GtQh3lDnGXsUQ2qMe40Z8rMqiHIMQDg
FN4cQLk7n/+8Fn2dzQaqUrOU4EO4C6MzcalLPKsDl4flJMN9ou8eAkGhjzWq
O9RbtG2zhUEtQoqkgS97HOAW57nQZbgu+1hv0lv6duaA4TtMbXfKW8VZ60xK
LFll5XjZkeLctk8wxVhPsAB6kUVo0BZcsciECTTavtl8/6tYCtIujDbe/YN7
isJmwjVtEgJHuMnmhcSTvoZC+L5J2QQcDZ/AYjEIcpgP3PghUyUQDhmoBxcK
lswu7IvbmoReXPJI+C6PvVrZenoS/ZmohLdewNe64bOfyqteWeuIqYfZ+ta2
pVF7BTBqXHKh9F+TgEZpsC2WI7ycS5l/Jwz+N9vBh2lRCc17rRLgQLRCGZbW
Xl7rO02F5M26pHQdrgwVJWNHp4rB8xeZbj+60YFTl/rVOl8IaPupBnts1PdA
xxEwief7aByj922E0jJUSrpHlyNRA88CfVEzvSYk7YaTtsFquKaNDRsHWAHd
fBTg4C5VG3oZ8JkNVFIH3vaTa7143nZxh2Djx/lUTIoA21qTu9Ztr6waJRki
txQpcP9LxPTvnx5aib/i7j0IBcT/+AI7cDXFvXzuyAu1juyEir51c0H+sS6z
EdSexgXA6ai7C2PDfbzhXehtL5OJAKxLttcPtDbEQAqhT8OZ8RlYI9ySq4Z7
/gjYvVjwgNtYy6cJafVAffwyUy8jjJ6XT/rtmi7AQ8c0+KDl9hJEwE7h4Pdi
rc4Z331mhfgvLymrrza/YOvAyLxNGLv3beiT+glVYHAkOJa4OJCly2pVqxo1
EKylmK/j4UYesQjoXTWXAe55m7kTRJmoR38YdCVDhFzsRSNDtWBgP3CunTxH
KoxJ4hoPtBsKknO5uMgQNAIKM3NX/jd8bF0XCg2GfFt6TTJyK0lWsrb1Kr1W
1uUC/ydmm8T0vEO2oggVgzZRBaF8pjjB04ASsFPUuDHiMTFhdDPgsAyTZ+Vx
A5WDFt9XGLBbaEioosgJA8lEm/sgc22GAEYgXbieFP0nZJKFLQEGewBxyjyX
VZadxarrnLaYbxcZK+oHxkRe19T6TNSUZin1WpKMbYeJ7DcKWbQzalN+wOyQ
snGC6Y4zIC961PFl1AVY84GBqSEoIh/nignBfK3pyFah4u48hISrSkpEUClf
THy2BTv+tlASXt/85lLEGcNodqDDs07pOzDViM+2ApAxkB+L6YKWeg4CT0PB
HjZEOSh12HyJPZkChSDqy98ZNN18IoExRkRDnObiSSpL80oUbeMAH5rSnlAs
qFTYcHPcHugAqqDpQnGnJqVvdSmMJN38CgdlsVyY9nb67/16wN/OUsMQDQlC
5doDSw/yf8nfgnbH0y83tINdAxCpCz4aNeFs5JbVVAIRm4PY4Uxx2aXjVAZI
xhXRWUUoukG1AvfzUAU6mGUD5IwYi0+OabOF/ff7AZsUwYJU/JLbmJshRNUx
+Y6WeEYAzvLnqguejxpargZX0vrJJsLj50657Stv6avjuWl0kKxbpwxlRSw+
eRMuz7CXi655yMyhXY0yeo9r2tZ4CauCHjmJQFtOq8Xn/bt//blRJOi3rEcy
5KVuL2g1kHQSwMeI7pfdM57S5IxY84p6I1+a/LzhCTMxnGzuT1ZShwh0lqx6
riR6qKgT2d+gUOuteQqe6chLW8qF4xhO2ErfhvjkAJDRTyk3YNvHIqgc0DmE
i/I7L8VEoUU0TiOUpZtVWJYUhwItRTmmY+tYxqg93Xp87j3MGjeYR1PwkI7u
LMQCMj9hq7YntHdUDaYtAfPxkktsU9Un6rNZazuXt6sE4ujNUnnSZtYFOXTj
Nk+Nd30JDb10x2OH6JfpODmUpL7H7hf5pzTQPZEbYlk/13x3jzNZKA8ATHMo
jYhHkOEkJtOjQj6n4SDe2y+zSB6D51fkZwWF5K347afrEzupvkwzqVcERGiX
+TLLezzcN2c2enH9XTaUc0YKp2dRMHCEzBsBiN8o2hunyeZIkT4AObB0HcnS
H6/pX1Lge0PoYkEQ8Bel1ifiFv6yutNIG/I1nG0Bm/sGKqdYvB1op0Td5ItB
phZLzXkgkgyo7mjzqV4yMv2etYV5dErFtoHM4ce3HIPm4Mibu3OkXThlKFvk
EWnxgl0qYiSeed0QA8grLbeyJBCY0Jhzfx3NYdGT3lRoA1tqMJ1/hI7I+XsR
MsR5IaVlpEcRfqZ+Kg9D003DZ7Xrxw+J0VQtzwzW5jy7D4Jk7BdRLUP+mCkv
njiZp2O8Q+vIt+H/ZOXzs+icXHx6BHEWf+N8LKfA0FUjwVIjg8Z6R9mA24I9
AArlrea1n+iM1sFspeZTgusWHkYGbz8zvR4CibBfulZJMq5WNTGRsZnl1LGo
MPnNTh3NrJSA7krSYw1XyWu1aW7z9RdUNFkoss7FUDW3fhWlnDt1ud9t7VLb
eyCjsXQGs5W995f/PDF8UjKnmdEXd1Oq8jyQrlIbpueUDE01ycoa46EbyIuo
5fH3XP8ET95rLQtdNCQoaO3eZXWxQOLmmNofWn7Hrler+IStrachdPRQ8J25
uXSH7vnmoiwHxuq0dVJCoMtlQSmcRX26ajMczlWfCDX6F5b4493JmUwAw0In
4AqDpmh3kPMy9NKTLYRnbxL0xOvKe32s/MGbhz18UnU0Vn8mLsNH5Jk4T7Wp
TWZQbyGPuRunFBLbASXxtxu97AfALwfwSVAe8SeVUBFsjpA+HfwyQqetYQ9D
0E9vKNsN7JlSEBAi0J/LqSi9skr17vLJtnLKvxEsKTzdc0gXNhwnEWoTWKoO
7RHVcAF2ilvjBvhiiRa8UbHmpsHwVcfYSNPQF/yAIhVK4sWnQvlHwAffa0w/
Dta1mPGCCWBG3i10SmjrLG5FyZCg4tAeLow9GSFer61OIjjuyP1DeQ8lYek+
Io5wVAMvJkbiGzgrPc+N34Tf82yQERWluHcnTR0vr1T7rRCKU5dpDsKiaQBf
czTnpl2AA32NfDd5PW9NNObVFMNj602sJ7BVRz/aKv7ydTr8dvwnFK1oCBUO
3FD+vl3u2Ok85RtdP9qg2RlPlNnSk8l+Qq+J5Db0Yzunmqfx8POL4gD0H01H
PtJ1PsQY7EHE8sNvrdBqAYRwB0WqkpCJSFK+beS6e1EDxrtY6dEtDKmV3J/Y
z/9YNSTWGPv06hDxUUnImKPSAZIyur3JhXBb+LgYPMlNLDMc4v1FpG2SZwjw
p6wbJhu0LL+RJXA/kTS+eDCStMGfnrsyrDu5ZGzDeQhlJVBIa2JkZWAXZKdt
J0NTa05dQP5SiJeHhJENQgytis9oS6NMV9dqACG0ah3/ZW2gqCPVS17Y8muk
E/PYb3V/31fDtYZp5LaY6cxAVnnCLL0o1h+7BlQ5ESNpkjgLs2jdnUfnHimL
BTRAuP2wY4ezR2PxOFLLnyAj9rk4D9ILaxtSzmM8CrJl+aTmSp+bVi1arhE9
wHnwWXh3LwjcrQKSDosYxtf7M+iHeK8BR4FEjr4BGVXEQ0gdXeOWfqj9CWcU
46aed02XYitoByfRLNaeRwJW/3kWtXhEByLo1u9xkXjnWgFziXPOcKSOystP
kWCfkessXgTp3HHm4LSP9UqBpSVEczEp0FsahGitfdWlpVmaaRHFbVp8AHh7
HeXE77rmJwvlOU++ZO5N3C+6nC0z95mEEknbVuvYhtUivH2Fcx/EWftPpwk6
SuCjyLiblrcJalzm9As7YE/G85ha97uI0MHHMj0baySzqyVLocbWRLrDq4KD
t+hSpP7LrzfNdmP3xAqgY+/urB+1YWxJuGVKNQwyyyhHrk8msheExVRxB7xx
QNHezL9T2p+r+PCyvikZdMLPu1uz6X+5z1jkEgPu1lgToNKSlWpW22LLRxua
/kA4lENXgNIPmxSeA3fdhpknKLvHt97O5ZpJk3UA1EQiD6yivcv4RWlUXHAF
MV6V+5JXRebYku1/3rbt7SFk75r8CGJQGzsid9D88xVN573gn5KdKbonCsbk
kVBjfMsIZf9cboaWZvZn8AFAJmYP65cwbOuzIdvdZLlvvlOFFYmQz7i5xkrS
aTH8ZiJ9YeJL99aXumj9SMn8veOuFbKGvXG3bvZr1JQBs72pF/XMBmLJBNqV
N8Q8YtwJ9JoJ1f166qwT/ToQohgBwmnIgHmfoMFx5pWG8WHS0KeVIpFay5XK
WwKOIrnR6MehF3mvpwlnJVevhAEK7o1PsBcsx9amcKdCGD2T2DEyBUH43Nnk
pWRr5J50vMKeR7kgDOEwGPf8pW5wbz/Obb7VuqsQjzNdJTvXBSDvI9ut0Uwe
/kjBumFf7rszhDyeVHvA/suX97DJYruRwHVy3gtZ/9dB7VXFnHUyvYed2YYa
uVXywGFfMymGjD9DxbQJpByVCTrauwZW2l5jSuXcF2zZrJUvOkE2n3bMWbgI
nzZXHRXkrpnA2UmBzfI0/SGJJU5GfWHcwocWUDKEPf8fvdXb2BdNY/AqevL7
D8j+Rfhet9WJ/7p0xF87nmaBQvnXL7VfEBbV8QjmL41hKM9bW/GXlgMU6L5A
GDD4xneTJN4xd+9CgRJcSYxeBEMN1uLyAGOdoIU8/iTEYuk9S7fiH0nRTk0d
gTgmGo1DzB/RgDQm+s6grUGEtEvkRQqKXM4McKS1wBXYw31oi8fWLb+jrPPU
fnSDv/XhoMoervTWyWLb6iH3Tupj0sfloRkS+KwqvHAuESX02khXS3vHeQrN
l+DcCvAY1z5rzGcYOmqkkfoJVtLK2W8roVL7e0/a2kUSgWECpY5j13neiLIi
mperU87EGyRCmcCA9/mSRP0eYJy2xS3kvGSI6/uPAbNKlgfsP4PEmAlTiHYP
eHVXii1p9jkIxwHVXnUya/L/4asVPHGv7aDapO8k5i8okP3R35OlInLb1bXI
Zk8vFJI/lCgVKPILRdPfW/3j4S+nmmiPtdxfkbOHMzvan3+0L1CUYRFWY7uR
gJOfXAkqmMjrXsXfzBcYXKK1c1ADqebFoVPjLqQ1p/ZkAuIvprZL1s4l/lko
yztj3HJWW7Aphz+6O1kK+BHVYU+0VLX/J8h585ZX56XtKGo+E+WzMWs2GU6G
eWMJw6E2P7uPDncXTNB6vXNMLA54lXOvrP1CvNeqgsPjwQKQZkDHxRoUOhnJ
e05VYlGLwMwcqZClkSf1FVOnviG5yjkV1mWqI8o0VgVQNUgKiQ37hUmmOYCP
fq+6eDrm6ZQjxTqSlw484baus/izUSYxs8n7xQ9H+Ww3iSzZtPsWU5bR3eDj
bBHA4eHSG54zurtrl4qtahhaSQxACuzghOUEe+2473135XzxcjObteJU7Yz6
xhR26Xgof6HhCChRuAG1rsz11pr0SEdBTpgY3XIL71pz+boGLk4+29qBjBHI
6gIBcMnhcX6Y3Y6L2TMhGDUhvTQiOR9uh/Pmj551eCYqtUpwgcWaULDWlnVf
JoSTk4J3mvynbBzCUOvOcU2/HRweSqUidCGX9HreZzDq1ZdTVWZc5iM2lJWC
xmt3VfhcSXeGVMuc3EL9AQtq9LWth4Jy86IEegy0YT9eRN0VRx7g0nhZ9pxR
BiK9ri80k/8XG75W+WU3Wb2QSrSWq8PqmHg0wH3SehDkwyYncmV+5EnKYZNi
v6aVKG6vSzGv+c6284XHyFNz6nvQ6sp6tPzRZ7p38xHE+gCOO/gT5nBM6qxM
a+hOLUsTzQ/U6xuwtb15UP5JH63eKWlv061N6nqPKIvjzxPFITN+Cgj0rfkJ
uT+ky/l3p/VOJm6pQM7YXNjH8Pp4AjkNzQhnKFy0l73ETGrgSdeoYPWFQ8sl
hpuiO4RvlNvKLOWGGW0Obeml9POEgRoJDhZqavdhFgHzvAbZE0/vhihx7Xza
2jKRDPRKRXObsTt1nufs0JcfNBbX2pcJhcC/sOsN6bxo0++l8v+4GRdRRtP3
IxNN26Nm2wGxXFlawWGJqnN34e2quFfnJbFKqH4ApMNv3+cyGvwAhIlHmHPS
5K/J134zUpU6wlIIAjtfCXeQYPaf9RpXyikfGd98a+6YLt59Knm32sl+r1cA
4hf7zQ7XFrAMI0DcmqsMkuzsT4jPf5JWMhPuY5aJwpBU7PWhZVAD3zgU+4W3
chLFtMYG+xefPRw/nSdaEZGdEWOK9wkGeczQtIyx2+4l7uShNXvX0nv5v6Eq
mGJ4O8GhIXBqwOtkPBuiwi6OU7NqD6paNDtfWeUgsWHYN5ybPWNcRu0dfvJt
1endTaCtPOGLqNxXfWn9jiQYBDLaiICMp03YG5X5Z211yUTbUkqAbSnSA4Lp
zJzC+rQacYO5WhdY7rQvRVFp3r+lhERiubdkwbr7ayBTjBbYWW1gvC1r6tly
gmnJdoqk4phhXDrbu27uw0YMhisem6n4aAhiKDPnUhfeBoORVAHEw8wTa4s0
iZAMmq9xkcmxZGc7PG+zU6ON0D+PSHktQ3nRRMACRbLqmiY3XdUQQcxWmlBh
/GLg1RSFZdeDWOl+jLf/R/IS7yMfcr8GL/3wBb43LNC2Dwy104YsPnTmnpQX
TdwInHTho/jWMGnKwtLNvAoTHI6X2sMDrOuEOXtqFU2HMo7RV34obIdouE+m
3AVWS8/5Bdy92xyeRWEbND4r50sxZtNygyD9jkQ0EgN2j8mypwqhlHDdw8+1
uWBU8kBgUq26/XSR4LqH7tQzagx+XX+YWp9UbHIqssw6xTQGlZ+jwJc9baW1
8SjkHV0Oz8qzyFHKTr/1qkvlUGb5zludBseTeHVce/63luY21Jr+TW3zmuFf
+kpd1OO7c+XiWQgh73r2QetT7VaV3GxTY50clkTsmigIx9zwdVtjlrFRfxRM
yTT2/47/Z9vu5IljfsaQSj6AmHn25Encyn3w1NiLaJ4CxlBV53CsPnSOnpG/
tEiBtdkNqtYYk1RcBtb0i6Sh93MuAa42FuXxWBCyeG+fZyR4Ic8idQk3b53x
9r9Fc3S0IRQWtVIb4a0WJgd6XmQWUope9lWtZWKnZrwSOKAUmSiLpMvAedEk
enV2uLDbCcMP+9jzMzgqZLOK3RXS+VA2sq+58c4H4G73BBDof/sJtLsKY3Bj
hMW+phYSqwf74ZmEaBKvj/dDUgQdsYB7qxGJNB4rPFaWiU8ISQeiioH/oxa0
0GVexzieAu8WoOuPa1L1BABqz5aCjkevm6pjNXiWZ1CYHXTkHhyQ2GKQds29
X3XVX90DPVQOIGwBZskFmrVckTgttikKrPNNTDuV9ttKlMzd7hoOQcv8zFcB
xLiCYZV/A6LxU17Vm3lob/z6Dt8b5lqxW/wtZC/O0jGvrVR2npDjO0FpK+nM
P1URujngnwElTgTrQX4F/SMPzgwhUNahUyQfFw3mkbBDFvEUlDHXOSh704E7
LY2PRwT9rBFInp4nWTFH24omjVGMilDzhWqFvM1pLG6omlvbAKFcNiyXWkqm
WQTeb2nFfiHoS3onahwTajPyVRMZztjarW1LGNpMeE6lNhAYWs2ONkj7blBX
Y/BBAKBSUkI7aO7e1GZ5MOpOREoifjNt0CR08EAqWcw659/Yh2qgCP5bfWym
x7w55W1AA77gLyYC/pNGVxkko2mWvYaJzSlO+Ppj/oxrUQRP2O9EiKfaTcDL
95rGLH+3+vymPX/M/V0KaIzL6SxadfH671DAdDyq1IrelW7Xem/GVBNLwXeW
zNgLucbAECFVQ1Jskpv7/+H7PdfRduhCNX+536EaBzjz9gm1BI3L2HGep/3M
M9DcHHvigrNCMYp0ygE7zF3azIIRNPacpuQVFD5hgQWKMbO2JMC7ul2YHVgq
rSe7x2QPPRQ+lmeT9MTQFXvOaXIMb1NfD/HqA5U2xLq/Gz57JpSxTaHFRceA
VdyJfNhOSQu3QIp5o/H08ebKTDLEqXqQmFjNSWzkOlxc34zh0R53g8WBkBhY
mVUyDsYaEATrxPll2gSlaM13M9dH1XfUsYCmkPkVNmiICGV+T2a9ZHYq4eRg
OSadsm/x0sBBLhOZ5L/cAjxm8CP/wPu9pUT8b3Jc96KqCw751MixOpbTIR8U
9VDL7yj69G5vXUhrkmnT4JoOVH5KILL/NJLRIXdtfzSyXSoHrdTLduwZ1A8X
jgxz5gzr4kaEPV7cS8EwUcYLOhqDfT4nm7pctH2zmK6i2XdOIkGoI7jiTEnV
lvkLc/M8U/05OLCPqT78LVeV6/dG8wiikpJnE8jO3DAxEjD7+oP4bMrm2/b7
IT1NbJZqNjvjL5jMBvvd01hVvUtbahAsq90IJkEvP80dtt+vN42GZPbS/xao
Q9EFYd7u68X/BS0u6S4IOHnlzBTl5fvepfUCumtAaCny97aXBAiBU9IIr2Xq
Gzf/avgkBxg7nDloQ9s6bPg0MlqAGgb1Y1Dl6QlXn0E7OGo656MnUrRzUfk4
TQsXad/BzUwxK0/7+LQIxF5cbwBzUJTgVffz84VS+ijGoim/F8+rsIwvjfqh
l0uqyX2KJgCiiK92VFUmN3xJstNkIV02UnUZDB1ywMmo3RBUv/pU2/GeeuLh
Qxt4xgCCpJGgeqw4CIDNFRjTxGT69axLzgOKD3ckOMqX/paCSkDnAL3pFofq
KI1IQIRWik7YTiOd8mbwem7JGWrTGhp1xPcCF7Jzzj6OMwgSosGTCLf/8EtB
h76F112pdFql4x84lEsyRxED2V0ZyaIK9MRHClfBmatQAiuavv+tHNO/stj9
lH3UCiaM3Dp8nJap29lAs36mvXB4YMU+Jn6dgvPzimSQ6mQNWMT4I6GAG3Qt
+BEPu9hC+rmdcBMXdVyCFYdr9S7fVZQqnqVtx3zeDdooEsZ+eJBQJRwmPgD2
oBszgYWymeexaVke6pV64TiBke1pGF2Jf07v4BMaRtVz7xmVZz1lVoq8z5DP
LYttNU1SupH6vQozRl8tRVywnoi4dMMAHZB6IYf9hTlYjBh+uhIEnRRlen7t
jbM+WxISUzfJUnlSu16cKE7YL43QYaMiw2IaINgnL8c5ko+nq4NJKoF6827S
+rVhNRrFMZLTEKweBcuGZjyGwUvrQn32I84hPHSysTks9senHjr8fFUsMmS5
8W4dGv96hpwDJFR+g45Z2BcJuwDhRNDtQDpEqa1pPI7NnCEpGIIe+HZPn6zL
NnB7JEMWDdXyjhSDtCx6ZAfEVtrH4zUvP6BPCsztve17AYxXLu0botJ+B/JT
TkkmNihVFrqQ/03bgcth3qo4T+HYi/dX/8sLt3J3pUfamtz/d95qEzK9nH5y
K1pddI/j1lMQFOLzPzTlOFxaMIEO1ONTTAdqY07vbPOX2cgDBUPDIXUqJ0f9
DVZas8hos/9RQj67bCSF5lsxW2wmRemVMT8TwTUDg9j6G2HUydeMX1Xjxj0p
6TpEtQuld7Ia2mTISbtlAz37Nhj0Dn9a1r52/PLbbgHMokXpg7f4+4w9Rs0q
wGdX2MXZC14YpS0JO62GqMGoUI6ERnjXjUYSs9azCej3AR+H5bLpHAXjnQGY
tdEVgTQpM70Je6Pmwfc1RmMF2LASS1n3s3PWi6oCASjdUgO6VId/nKA+IJzJ
QUua0tPNJSDYlxk642FZEXgZCkNEgznkz7SkepwWeluaktd/fqpI4xUrLhwA
J9CIMWPyofW2mg0dWOXbb33e5P2bDGT5b7M6fr78wWCuJp3o1Br0plLJ2OqR
8x7+1Who0Z5SBM9sudf86wZ50timHssmMZ+BR20pHSPVSw84pOgj6dyKHEsF
2zmVlcMwHXKtHh2yPz/9BgrX481H+7a+O/K5fNYTZiYf3SQH33A2WXwjxOvK
0hLn7hGJa/teSpHy+7jNo85VhxVm1At5bzM5n854P+U+LbEc6Bv+MrZ6TDsW
dxmjKX3uatiohdJ7hg8JziLnbs2vLSPDQggDfdG/lgtgnCh7/FisKYuRNc9K
CMLS2kWbgNPU+intJULu8TVqcexNf5ND/4UWUwnFAh+aD3P6ZjlnPnn51tgv
km7pHRMpsYpou6K2Smyq41NOmt75JWaX0TrYCT/iAlAyxCr1JyXRDzRLzchZ
Z+OIW2QNng0BOTnTOwkKIEndFK0wbfK2vGhk0IXROsyDMeCHFmHe9hqHXvvV
yLJT2Y1oOa0+UWE57yAISIZTAklArjmQUO/TjjJWD9PjKDZxQRntEPdrLqCx
USZNq9UXmxZ3EAxk23H5L4awOsQ0s48iI/RWOnyDffrC5jjoscTMWW9cUKpp
EHeX8bMEtwcQdzuROZArxD4eu9b1mnZDpELasKFi7MKelIoq5PdsNMUgBd/e
dZw0wyog3WVeYUOy3oIJ4iSy77RJGuV9NEfxEfYKhBfILa7D6VtBobdyefgD
BT4SqBsoFdPb83eY0kBulcAMJYwcRGzSkB2gJ4yA+wfmqFANQGJbOfKgPz4G
MOX2T80qOMav7XotzGC5LTw4LyNEAq93j5mQFFsb3jKIyEhie+qJHqBhytIm
cT5faY6w20FBc0yWE9IrkxailLlUBZYv0b8T71Fv/PukyR61lr7tSVMKlofB
PQtJV0KQyNSEOcDBYI3+zJL9ZpWd8aupUPDQJhL/uUd906ZPoNmwSpS3Q/bU
zrE1XDVE4Gx9AF/nnSz4S0YTr3DRzrsz8ol7Bmz+bPKcZKTxQBrKSG9U+kcN
mvYW+klKgKtPtXuR39Y6YYCWyHaptDL5ZXIMNT+uQs8F7rwtOQ32VWs1/uRg
NjYN8y2KKTQnZwMO2EP56RB3lDoSP+vHyYyLxVJGZoe6S4I5oSnd9ucI/Jqi
/G9kbnd6NJbPsmqAPIFva4/Goryz4lAMP4487a4evYios6g1KHaE8/W0pHs5
hH3g2ukzfKDThu6K3xdeRW1F9aSACjbXMFPXvD12OzYZd4T9Q0mkp7gE/aNn
VXRsfNXs8k/65eq/MCq504vCvMxruFOO7wSVJUeh2V4uofk4KtAUWNHEJTIi
zrKwVNRZacZIreySv2KXY/ETC4LXpiIl+vHVr39PX28y7C6AJ2ndSZwPGQXq
7QNEGtplPo9WxjlI8s4nBTNK2TZDzi5eB0P1g6oGQ1FHK4zmaDEBll9ypkky
+X7ctNxavmfLh3+tl2+n4T874W4/V3wU4zoWzFbzJSXl1lXArJVVxGTWu41D
6bEaBqIzvK4l8W3wq4rFYb5zei+zhShbl9Ze9XFcXkBbdA63BS7iNu5jWU40
keA3Bd0UFB+9vO0ONz1iDIA10cSg4QN2u51w+anSqtqs5lcE57A96HZfHWeB
BF7ZIOkPCMsbf2c4sWF/yqnhj3M9FN5u6VDGRphK7NJ9quii/tCOli5rRbqF
DIRQu3vfwB/liAqSLrKzuiobGx7yskLb207vpBUeYBEcHEKdkxnK8VL4IduY
IiLYcy6r21AXPFKdFccKn62DwW7iW7iz1H0HDKXqPwwUSE8XkU6JhrJjm3NX
lsja5EMK2bkavd8x9ePJnkvSIHC+NirJmX1y7PAS3K8NR6/DYhEx1DW0YFwG
/RIUgr5ntXBdlBTFxOnwqa83iI239vuNVgm/b0FfzcacUK+lCSJnSq3M+02I
/u86Quw0RtxqkdVoWlymVHdajDj38gugW3XEJo5+82wjqdiyiVnwIXg51XT9
gI+TjuYIZ+nfJqzpXhkRYvJv6jMUkHIt9QotXGc1gskUkhh6QVEyPpJ0aG3B
Sr8qXNjgRNo60nQ2MBMqrQ7nAlkdyqqfZuYp+8Nb6G86oLGhUQM8ZUbAiW1Z
REPLIC5BTBo5sU+PuDe/7uUvZOia6I0OoM3CTJ42G8sCFG8mvtQ35TSudJIi
1NujqmAzaeWuK69HXq+MbqwDzGKplwCrJ92QHJzz35pd+r7IVoaptE+PkU1i
Yb/kUIfzt4CDE0iK7Oh0BqOB67K1S13/s84zNP4ATl4aYpNQS62qvqLXg67T
84W6vge9eDUPh666BNTKvznb2McVL71AJTJzZ7O8nJlDvW37t21CCIhRyrwH
8qZsQRf8S2xYn+51jT5zGYAzwRmNdYACNROg+75TdJ8llZ9V8s59GtFfyw97
1CosQR+0wp9j3LQnHfquHvhTBJRXwmVbi1fXJEixks7mRJC7TMJsuQ9v6jLV
I/jxIqhxEpPOphqioIIYI8g/Xl7vc+oKMG8REKtUHDp+seaHK1HainjhesxB
ZDqdmhoiGmkDLn1GDAOMbjVzwMAC6KYSslh6e4T6F6lLPOQZ7EkQm9PqCcAZ
kPuufu3buHCLOzEHGSgi3BRa5t019JglitmHP5qZI4nyYt6zyowBkRavD3nw
mUFHlUfaq+Iy3uu1iFtOw4920aVssqH3JOV6m3/bv+0tBEwbVduNh2h+/Cp1
nCqBHz+wE6s2KXANLC2+5AjGb7Eeq0gEk77Jlmrq2YTvEkMhmZbjyFgcNRyA
h/gbId4+GWkPU3Hzsh1DLDuxJBP/L5S9dn3IOAgXutXdD7ydAPOhLI0rbu4L
1NLURy5yLKgUj65yvjgzGEG92pwZ6S0Lu3LqWuAwIEUFbuwLXL/BuuaLFO0y
GG7ryQmvY5giHKOK/eUjfnjFCNIhf3rERzOqXe5YhwHIBQnDrD2vCPb+yKZb
23uBX4ZLE+fhUl7ErQlZu46pUvwpYgioXe/PKeTvF2EhNoNnMdihHqQzoOg6
mP4WLFnoYks2Xct0wStf7I/Qw32ytTbtNhaLAkbQQ5Eest9QCCiC0LBho+6s
/fNNiFzRxSmptNrlyceLhUsg7+/2zP5ETqu0nFWPveL/C+j4Kv9ZOTkO+i1p
82OeGPZlFR/GnUTEqsjlo/rwY1F388ivsIeoZtQhFS71ZhAy/+0EAlCRqWaW
Fy6dyLQOMzWzzW0JvxI/LaNNRMIehh0+ENvvsZ+CJ/yMC14ilPn0ByNCxD36
Dksyzq5Oblzvq/ITB7vjg9Rph3oRkmSHQJcbouUJdk0LXaMQ4m/KQ+O0QKeJ
CD/1Tx1Y7L2Fs1JDJqKrfwbKAPl6+o2rbs2t7v5RSyqvwI9A13MZIn2kGzOd
Kw/Ctm98aU+WZXy1fQH4SJD7DuCjhv3YyKXEAJKO3WPE+oLS9Hzosofr/6Y+
ptqINhPxakx8AogUKSmpOce4erm3FZqNS6g5UZX/K/SJCp60EsD42NYvPz7t
GkyeZT4slr34SuQTGlPbkTS4Cu3DJZzFG48QwZQXxvOwUHH93nsSAACfEKVM
tejUUyjDTIb18cOnojKp7MaMn84XTOKtMsZnPVwjXCNerSWSH0oocbLkhAQ9
6aaEMJe13PsuOd8yt50v7B34us+auIqVn1H2Q8zBD27tOfm5FVhTpt4Db80A
2eyrbRaDguqaehu1u2CulVZ1KVLYn3cBpG8wB2g5roJAe0thHpKa+OqICqe+
kulwx40tA6QsgCzlmltmAqLplKS/gyf3BlKlTTSRZSnHO/qboek3oUiDt2Ou
PXzjGVvBjCFNHJE2SNddZoZvR2WaYtZNHje1XRbeWoX7pz0r6fF83HELvd00
vx3rXRyshtgR+ibQD9ihPsiculoxFZ+wyiDBD1CzY73uznsDZx6ufoH3HozV
sKR7wM6InFU5BHB32rNdj+RPhFNeaNbtM+xLauPXH1nNTkD4y68akRykd+p4
V/ZccE4N4LBfOYRMACYWNxcpZDymFse24lblWoCLBZTgU0tCUkXF7FCLQQlj
BPNdyppnFSgk5It/pQogNmpfer5XS240aO3LoTftnhqXo8QbmgiyB4Ok8hNB
SwqZ7Hbkv08MHscENM6cIU/DybUHThw1y5U80VZenh5K7ig48gfMxP55nmOE
Uivomxb60JPNPYQTlbRb8kqu+HY+S1qIEgEbgQALEY7dpy7SjDhECBZ/hYom
SIVZYNG0qvVhA+eb+rg88JxER1R510DFMXjMNtwyzVL/oy1YjFD43XF3Y8++
vq6gT/PGi+yzaya5BfWnw++IopHgo+sT6OJPJBm3kn5VpXFpzoqFYrg0QYrn
gVowKQSiyFDZ7KlYFuL9EakOpCcRBYIX8aeNoeR2c+4n9YMG2B4bcWCn1Rvz
4A+F+yDuL6BUOjzWd5a3ImcLz81QNnPH61/xPGBlKW+m5r4uZONp5Jm+ZVGy
3VXFxl+N6JiXhKk04UnsFlTRsCtbkB5R1E4u6YcnMPZxzxvpVb9R0L5cWAJq
gavIOjrlhnAVfXFKVTDPZq8u8SwFjfcoQxaQK4TLoBFDd6a06eiGPZ59WIC2
jFjzLzTOCOvUg0utyi9Wn2nXRvyPek7eeQUowo5zGUJiLjxZa7WQcWTsJ/ns
C1f/u6KOeb/StLKACH3MCGO64BJgJqE2O4OtYN5JaXK1CN8UIMvP2mepUjUt
5dWK13jSFJEFfZtsLv9SHm20TqgChLmGHgIx7mz/m/b2lCe3cAY85yonaw5Q
QBdo6vs0+EBozwEEmN+NZsqqN12dJnEH54u9UyWcgPZ75Cc1N/sQlpsJPtrR
nfb5f8/YBIjG4vY83cy4z4d2v24OTFn/0u1eH202KtORx6vK/yOI4uo73k4z
0IY05Ia/fZ8s5rN5eqmAMrmSjc4Lf50qjrWjPK8BSsDfUUAEpfNHoetATXPH
ZL9sFKttv7VH3Nk7SxlD6qo7UouklcNWZdtxy/pjLfAcrd9D8EjLajvljAoa
j4J64Ivbe8mAI31vgr/Y0c6K1kYx5jV1nSmInJn1HMmLmqkVNiXOV3Xc5RyC
lkrhUMSKWhQBCy9cso8DerxvuqdMEJCCtDsT+MUDkZ+AI9U6Z1MsKRSvZCMu
R1BTAVdHVf5bp9yML7Jb7e/mk/LdieZ0k3V3TBRfvnjFV7PFlITT3fW5rk86
7q3P+51fm/VfrYvBGgySTUsbOlhCz5rccUxot8kYgA05h7yvCYVlG2TyBDGT
hG0rq8KdfBmWWK4Ht6AgVrOhwp/oS5fHmmR1IVwnzTLp/PSmlglzz5jZCEEA
d26YfxvOHt0khT3GWVzw2AMS0f7BJ979bDK3jJQJ9sjWGGE7VJATKUpQh8Zo
yyP3ffoEZSa2oiKng8S/obw3R0w8AGBrPrjyEuNn1tQDw5haPl6Hrp6JkBjy
uXxSBwDnRHBu20HcM9AiLgaU7HJzCQXbo2QYJ3VG+Dw0cyR2I5j56Hzkl0iC
OunwwD6qmnzQOrYOWGnUhxzfh00G3WMUaat8DDfYDZb6jF8oOtvEJC+cZhFp
BPWrHMNdMjvoi9qjCUsXViHjbf1jE8xC3qc3CGPD9tpDBjzCxR+QNg4O++CX
FY5w0LuVttxifT59rLQI2rym7tBEkc6yd/iYQKZ9vhNaniLQR+J6YxM4Uojw
juhWsu4q4xbOudHPdfLWukDIrcHnngQ0i+WZc0D7BkuJ208Y2NG4ztpLsYb8
JP4yX0e/k8d42kekWCC4fkp0TcwF910KAwu8e7tTtZwZP4OHorx7ZEei0AwI
koV9qInCynYr4XeD1vWlhfpKQf31yj+19B6V33lTk0vA2alesyZBYol8GlBJ
+2Btoo3xLvZnPEobSCdUpNJCZ4XoyTLzAPvqI5o0VaJsBhAoTKX3J160dFi+
5QGbq6BqkmHAVh4BZBnb9o2cRHmIupumMq91zJw4W38Fk+thIdpviCs1vLc4
CciMegbjOrJd0ruc8YmhEpYYntCGzD37ri8xiuuUDzZV+o7Wtt0eCTb3q21H
bTqjcArA9rKNYFt2m9/tB/APAOgwQTW0ldbBWP+1W1ofHWehQE9srpJ5T8Ct
GPJPVQOaDSFO2Un6yZ1Okbt7z+58uYVO6gybfoICKaHzs2PHJ95YJKFCk7xY
b7egj5RtPeK5YJEtU1B7T/LsA5cBBpiNpXynjmTuHEXJJgBbYVbutAF8o4nj
ihGnixpgQrWiL4hiB7jqX8QaLWg3PHMyF5WFd1e1fIaWmkE1wHngBdJgFo0s
viovbaQTOmgLqKl7+fGp5IEVeEel2J5WBleZQoPJSlV+nR1cbj92+p/xKwxI
RhM+nkLflkN0r7yBtsVBzKpNNF1jfByqi7496VIeb9csKudlFzZ2BqR4uWdw
6rwlDLJz6NDQuLJk5/DZsMjLHU7ToPwOdIVR1xBUAyXzIAszRIzsF7KT+iSs
XB++uDRz3tCNaktLtyyboWoJMReWF49Fv7/0QZGFLNqhVa+sXWS4XdN22qG8
oK3OMoCy190kJgBG2bFX688n7wUA2uZz/O7EfvV81tlu8yYHsFf6E/BFy5H4
k5tvZihC+G0DRyfIiuNlpgQ29xTmSItAgq2jO47UnVINqABM5PalfDqggOM5
oPO/IuwXlZiBopQ5GPkucLOdO5EXIm5cIqghKp7q/Dm2DN33C4xhkRsH5+jx
4R3ZO8/u+TUzI+N3BjYJyWltyBVAVkpcSoj2EcE2umRgwUF5X0RSPCypu35m
efWJg2v6ysX1Zjgh5LnW2/C9WlnOYLND9hgmt/ArpkINOXO7GnAa9Gqq9WWf
qpAOlGJao3/w3gd/yFl+shqv4gy+u99yOZBxO5VFAMXU6w/ihAG0pjbiuhbw
Q51DyI8O8vtugKoOYQrPz/nSc9Q+PN3uZXDUKP8Ji7cXyQQAWxp4A3lcA9AJ
40z6wbcQBicc4F/VpgjivkWhbKdMbgsZNRpxz6nSWuKSrOhFn/57lHiPToaM
5GdxQ8wd29tJAqM+mljhgtK+5+nhAx3gD+nxbWTZxU0GNvlR/ExrOWqvujLo
Xqud2Pr7gzj8Gilb7DogPydBvSZQbXzT/kqYuG8J9gxA787l5aj1nmBy9oc9
vOte+SThm3JmfPq0uyMpAz5tqUh75PeV8teISKsGukNUfhhWgSc/ZdmE4bv5
V8euPT18yqbfq27yblXNeJub0iHVQ4BTUQeICmWF1HPX+F9z6MTxsXHNGuNt
vn6VmF1NtiF8Vv+c+YlQozRmAZ8Y3QAnv3R82EnafWnBSoxIUAhAbJRvaWhA
Oca8mLYzFTlS6s76a2FPImBJe4wF9KJfsu2UPB7GRv0Qx6M+gavOd4UQLyuQ
xFP3sXarYS2MwPQKF1+SMYnkW4Ylod1HKJcZylXobB2VNW+O3UQqfBC/wOAl
nU1BjhgwfbIRWoUy5ki60qLrMiI2stOLxfUqb3kbZ24aL4sNAMwS+gPsN+A2
zu97gvAIwGomb8hDSKPnnMntk0wAiXlRM5b2b6ioUr7IKd9GQ6DqtokncCaj
X2aAgWtUtxIKIihqpvA3PFU1Q0I7wMboWy2iSUyFEMe0vxOz82snZvAHyXtS
NWfje2hgNt2MoPIDh6NU2VXl6vySC9AjzZx0TICTEuS8wFR4SgJDEwvTNby4
+R+pedWkDmyjHh7Uyh2SfAF87O8dnCLvFH7BPYWwFwNlIRSvlbb37fgnIdap
XItBclpsehYn5iEYKOFcfrSNtVkLBFsJ+ZF4+jXAtR6L3/kvRLIrphP/tx+I
mpp8HmZs4z0ZVtFXec8IYkqWi5twaWeagoopYjE/TzfoXqcb8c1JHAd/i7Vz
s7ACU8XmLHWBIBFogJ6axE5mmPANFkHo0gbFbRVoL5WrmbP1+ZkJ/+kvGTcZ
J/dhR0UN9yhoAYu/nlDxv0oYHB7JzK7mul16OtQerIG3RP7KaAEgdIQg8Qf4
LSMrZtO43YdEXZvX9pauXAxnkHXgss04UfSAE4BQJoH3d4hllmnENMfHVL3G
avhK2BF1Fnt6rcOlxewzIrug0B7+/XdLsGsHocaKkdFgZMEdCrJ2IsHS5mr+
z1dHX33Fez7htWZkwbH2iXRchy2fPI9TA/1LuBR0W36lKTd0OkXx6h11Ej/2
VUL6UAhegpf4xC+x1X7jmPagXHS15Jue1tJwosLyW4siERXETZmBN1VTWzbC
GPXAy8WAG0Cp0RJ+sdzm3HwIFlsFFxKT0FQ6JqYentVf12MZhueQY7tR0nt5
WymqAebhopsnYUWCR2nub0WNVJvpGq/TSJG7iky6ELkH6hVjBimiE4atnZMk
rm4ni6qux+HltsOtTMuZQ1YzM/1zwVyYwEaeoh8eOVq2ftEEXxtcds1lkBX1
2ZxpTE5hONL7ZJP6Gy2PxKcA/emaOnLQnc/V8DeZjwU6dfbmtYMB0QQ9r2Yc
PcK3TSMayOzsrfYez7H6p4ZPVqG/UO8jrPtLloesMNZdEa+tkDQuF3wGtYE3
vVyXSJYVsVjFzOcrrALYUbAij4nW7h2bBJtKebJ5xrfmnZ/WVMSEIlPCJKR8
YXrKAAMZxj4WxksdlIzpmmEdDAiy7/+Hg1C61Svl0GjGGFSxQAigXV4c70+q
/q0911u73y9kF8Zu0Lbp7dlGL4H0XgU6MiGR04kvIxSm3JBWuOLlCsDhmTpP
PnoeSkLOzM2rNtNBYjm+Pxez58uP32kGak5IwIzuUinNSP5kn4h8Ut08f1tt
08eOJBgE28sZFj4JAF1U2nfq53qESnseS/BDDtPu2mZlhkvWwkger4Oo93kj
+c52UH/A0RzxYg42ykS1neJrueB5Q1Nw1GcP8/deYa/9MncG/8qu5j5mutJX
0Qkhx3y9uQy6Qm+a8K13K0IkX8buZisdOjhB9Ey+/HMFa56J6dxmnqVEgZQy
sbuZNAV7T26BXOsWGg1EoCDe2JXyKfISgXpzDKDdRCHjp6E0IT94pg+VCfMa
RZg/bvSUDxL173tr7yvqDLLlgp0N9hNmkusUPTipMPWMrApXRwzZkWPkcw0j
0+P8wFjdB7PI2xQnYLjwnK1KQBPlHacR6oXoT/zvj/bGMtfcw7E6qQK9z0KQ
8uPQDI3HsP8gi8zIZrEOEqs4MzPjHKxy82n9ET50a8+HSUPhbehtF97oQVT6
j0W4cbr4uFK88P7OIN9iUpfmG3QxLEyiFTh7OL2bpMc/wZa1liCd3t2rDrto
P4pRlQVbAjdCLT3fxGVsVWIaLkWrB/6LX5XrHJ8eqLMG25wivdDqgOQm/lzg
D+fmB6cohnptLg/4qeUEFf1RodbUTLO4d+eAJsdjlFj/Wwr+oXTeMne/rkcr
OyZdBlRNSRKfmA9oyszaR0VQ1pwiDYHizlOYiQ0jiOd5h/UaAng9Ayr9RB+h
Ds+cQEXaxhqUBvZZdQXJrPklrYG/eOP0Jn0uUBi8Yud+tpKEZcctOkT29+CN
NqSloRf7rSbPt9RsOe+SY/aqWDz9ngZz2+A7c+GKTZiLLxA467yJwlvR0o0E
0KleAMZVH6B48l9mBpCq+HYqhqDaWDIUdBsK7U/3AzN+ye+7szFl4RLn86MR
reh50kaXD0SOt9lGL9u1h9ye0LAMmQKE3Fdqgb3bjysM5Zt1/oVG/iH0V9YL
aT2xnVVaa7SVymtOpblMSzfsRqZgdjP6vWbmB315vYHFbi2BY7/qXsvtf9zN
ChRAmUmSNvB+oBoYgv24SY0iDS8pyu8DvE/P0mOp9hZR8eSkS/9c6vUXj8jW
wrc5cwNa1GLu7OXSeuW74LVwWe3aBfu7+VzfkiX1RPvpPq03c+droUM4Divy
ltYDTP8O3BabYMpMZGw2BAJTWialpTpn1GgR77vHFqfJgf/Ei3hrADVAE10F
qhfp7ITN9pZxyV/jARCUQLQ5sTK5uZT3y05E7pIVQKrEmG8MIL92SnVbeia+
n3b9WPA3l/vrlYjgETWGFRdoQwx45ijyZ0tzys45obZ6gInJakzMsBBYH8uZ
HRW5/1pWQiNzckHcWzd1bvorPlIeuyDEEC1PZULyWx6AYnqKVCWANEkdeCLh
dgICZ+uRQwDnobK16L6PjNy6n0Bn/Mfp6Wf6ACVfurhj3dOmgo3xBPsungsc
F/kQpmAtxyKL2qkhFvN+pYezmE9qlkkTyKhtDORBG0B7s8I3kWnW25Cr1MyB
MemCCo5MbM0BbeqTrgEHD+DL4Hv0HawLcOnumwpCuZclGdlPuO9d950U9JcD
3tXTttJudBym6jqd8+xv59gmaIOWPwhwhe/DEBH1+zlxfQ8kQjiHtE1iEFw9
k9pgy0vr2img5mxQzBWMuEEBDJzmJ+Z5f6bsuQArGF5+vbCiwXkd4W3kKu9B
lFE8LwWFASzQVSSfbWkmWh1urVk+VqkzA5KUjXLNrNKUYlC+aFLYokqqimmh
2PP/Xf2tTU/ZXkUzjCPiufjfkbHO0dMKIdBt6BkFXm9J7eJZVZM/bhRdWvSF
UHGi8/e73h0lyElFSDW3+ByPcw/TpXU3yDH104zD+G32wlIXKfIa5n5hAOMs
l8SP3Ehk2Y69+hSOrVbT3PXgSeD1/VtvqhmiBNne4KDAQv0qeJgN5npc8Owe
5jZSIrAB58F5lnXu+QDAB2t2YFuEJAbmBKUwC7zz47reK2QlVdSNqfnB56uZ
3HjztLDWgDu+p0B91oAJmNySb4NG93cAcudK0kgSeUCJF/iZcJcCoSSYumVZ
jRr9jUuGyvCvbVFp8TQCArWGpKCpXOzwuIN+7toVyM4cvio6wo/EswqZ9X10
Um0Fs1/rwgrn+zOP4PrD+zmTo3PVbK73PKpL8aECLul6r93bB/4eI+nb+NOF
U0iulrpwO3bRm7MCIC93XFznacDH71ztYt57z2xw1uBwknrziBbTpt3P8W4O
ZItfJf08yDHGD2YNonQnoXGgYZYzD4h9gw4ZFMvNnidaz91xav/94fA3sNLF
JhmN5X3XGx+TTbG9PxZbpKl70To7wORliKs9oMOrH8Sju4EG3aXyGhJAYY3E
i1cUX/CZ6ArfgotbigRjVOIRJvGeslTPyjYJXMdBSqcUkIsSQBqyy5aag/FK
7E6j4qq+81jS9do218DAFnw2t2dWQZqm3BVVKlDXVGSDlvgfsjU50hJTFctB
4+3+UuL+y3r/RFSarEBQc/i2P5GwEDfWFQ+iJLb4l3VMxQdgdn6tF+AcbUUS
hmHcrm3LSiiktAgPqjjSxQJdNZQn8DDyAAC24QLKrMNNRsgA7EC7yisJbFE8
d00Zz1v4nIE0GizsGMQM6gCRCu1ICDX+lyCEXFEAnlsMcbhJYZKI5fMalRqF
GxAAjD6SBl3tUHeRsejv1osuDG8v4h3m2PMeP+2TA+EtuLwd9+wNWGmQ4Q6R
dxHTgyPOd8iXsG70CARU7DJxWvYbUQScEdMgs2gqjU05hmkQtUJIdTwbhZl4
R2Yktd12e6nYK+PbxZEuBEEWUDRoIkEp2nuU62OMvuOoM6/TxH6NbnsJXpZ0
FuP/HMlepvIUZheGsXl5JDp0+QE6B2R7LFNy5nt3ALaWOVDrN5jJBBvfePmt
MIhHinL1viVapeWc4g4Ky9++wYcIE5kmIvgVZzeiE4zCeuIvuVPZz98nKUSb
PshWYyBrduHfjNkD5d64kY+hR/n8v3p2KjrDXhgGQaN+ueDE7ijUQkk1//bB
NhIuTeSgrl0+MCtubZY/j0XgjWvrEfG26mXfSRY1fGSvfZcIETPkaqTD0/oo
Mdb23wTFXYIYyLzast61NLbpu6IdO/CAWzBKz12dRaMNNqlqNtELRKyVUMMh
PQBa+5C7aZias+cjE0ilAMq+LJg7PZU4g5cl9A6AiUdskquBr2YtaDco0Lg4
+62XvyKcvNg0ObI85y74rRsv2FKLTESsX2vX+MumonkwSCteCJg/p2CmJS9v
9lHh9ukM//G8S9jnKMhL/V3L7adqQD6N/Z0utExjpS8agAkTZAeyYalvpRw7
lX08O7j5pu40m64W5IIwvROyoXQqSVQvRz4ViGxG2Ak5WkeHTJON75X7bwt4
ENFPu2ni60slPZu2ZLHyWITo0/n/SBgngwg5I6A2puJ69kFeCB3qJKWhjNEF
x29ZgNe5lsmF3+fb8aEJdjt7Hz2J276vACMmWnt0lM3GN1u5HnNdEvrGTNiR
RnM1gSBm4NqQrNvCdoxrSS2+v1Kp9Uyib+y2MvB95CPjrrc7jfOOaiOYFEPY
X51eTVdDv0eNlmHZbDnYfZl3cKXPPFDI17IR/N+Uinow2LIOS12B1n23PLg/
S2x26SdCFTvXmMIDuswoUEJjYgoHA2k4e2xJPF114RaJ8GggC/sPuHhWdXdd
VDlHOTPwTPZoa6i6wxmfZHbp8u+ZoNPNp6p2+nEP+FcFsdKUAzCac0AH6Thz
ftEN1dgXTJUig5wCVAPaFReK/NkiM4OQ5fPnGvIO3416LDXlZHSWEwiR4pt/
yHnOJwCYQcAaudnbaySL2gm0wpw3a0BlmRsbefPsGRAyaiI8Cviej5s21IX5
L22k5oB3JSFqFag75W1iByLY1EqsQjgzrpkcZXbrns54nBLTONb/WGbUxE99
LqG7Pc7y6WohIj0kd8QaRVMmtj3Y8fxWKu4n4QK384o3H2oTY/Drn2CJfJEa
ZnWfPf0wnQRXJFxXQU1gygY8uJk/vU6Mqu0gV7472C1WXrcXzX+/vVrxMuHG
kDLp4Uk90cK4WntbHZ+TJ1KXI5GTmt60/WkdxJz6vJjDhWrptOLObXp4/AGr
IZbFybdHAW1mmSoPP4QdrB/VpC7SY5V0g7jHysPksnblI/1bgZOBkBZyhl3U
+7h2V3KUpVaQL8U+4X8BSTu6i4oBS+oBXJLHrW1S2QyGWgS9PvEhk/vJDPqE
SqTPxlRG31RBqChB+WlgdATXQ7/Zj+CQBkQexNX8pjlNkHA9uobuCp7eNc58
wj+YnWuWsxvywg5MJUKrD5DeFLtcdyFfeJR3BymwPiElTmHW4hKlhei+2es5
HWvx1/7y/lVdtUrO/iNCvEAGe8MFV4f9V+9IYuu9Qo8Qx4E7RNRvS5Bg1cKC
BYdQZP2wYsihDq7bh4IJ5vMLz+cZhlK8s3p7668pJDrF6wjhybAu8Sd4YdW8
ACdF4cUEJS3aM5r4gTxv2QN5pkcE/CsTV/YdWjV8lGwQwbT+2jplOOK5PJ8z
zoWhrs30fT1d2xlgDhk2mb0WLZ6PSGHbabyr+1fmqdfOyuvwioQdUMzpdjL4
s/3ryB/aZbxUkYXFu1pov3eHoVcjexrID6Q5kGyRY1rmMaGVRBKyvEgt4o25
d2g0siBU3wHfeIS0GyMeDzkBSy8Vl9FSo/GgOx0UG2KcBvjamGXInyFp0lFY
0zPvgWxbkR25itQX8qvniZeP7P3xUrq63UrD4s3gNNevO87JDTtNx4nDi2j+
NRdjVgGfaZ3OeEowF5ZQ/rzqZe31EKWVouabDryHZrXNhqjfDZkwEX37zcxZ
6Urgq8lYUVaYqA7t5lTsk+e+qR7q3Czad/BFSsnP++qU0zaF07QTPwrw4nRx
iGW3wgG2rufx8Ngye93h9dqiwmDU0LKcadGC6VLgDwC0VcjzA7pVNSwErwTH
+d61BzqeKQYzl+g0p+OdzdoQiy7zB2UGt9yf1uPt4+7SK8caZvOygxjnDtSy
qXMJxsiZzI+YJuiIG5u6qCh7nr0bhNfDt7BS5UK+tPeubVzN0K4gqEiOk6e4
iPqDazssaDKOXJM2d321wXaP2cyMdUex22Y/YKsMK7gOgL5eYAvbEDmBAbFD
4orS9/g8dUxptLD+IEIpFDcPGgnTPGWl2cAt7gDp4GO0ABxlOXCJ5USd6BU+
Sfx9CIslGX6coo+Qivk5qchek5vzv9ouSUS/EZNtAY/oDtL+F5YD5P0lK085
/nxUdLW4olIQwX0n2vKAYiCPk5XI9qsIQbTMBA1x/NxLVJ/jydhJN6AAL3D3
zVJEhRsrHsJDYuPkhP7cD3balN0HBakJdx7F97yKkY9wDFCqbGoKUxccwsb7
DwHFLQXMtUUz6lKGgsEvEyhHkKc/Zw9y/TMMVxe1yLgBkAmnzMzmjjBF4pcY
wrvX3mp0PX06B/ofvzKdNhBhilx/PrRbQ7ePI0Xe/BYUpBNsiUWGTQcXTFDl
FEDt8e8nUTwDWVHsuGgq+s5hEmhG8QOlG4y5AH4s5/5JeenC2xTlZZ9rnE1W
uyJXkFioTXF44L0FXWytqUIxKKuoBBndTLf9mMRbrj5VvG6HeI3HvObyL3V3
TbH/zNL9vncjfukC74n+Q5NQ/YcggsJvw0rtvp8epM3z2YhFUY8Ua/aERiNR
s3/X04Yzp6/+i0uwx3UgjB3krQM1MYYhX34fhgFZVximDvTJ4Mih3EfdoiN7
nPlHmObGuFL2mfg01s336cl7dUL4YfIZzpoPc3UB73e4UiQQEUArWiwOWw3d
WziksktAF1A8BH/fWMTyyZswEpwIZv/Y8GWKd8mLgY9AlVx4BRhWrgHAo9Of
ROxNted6+pjaSaD/fORpazoRWCRAbkRALGABQA8Bnu4QGVmcyfwqjp1gt5JN
rYYPD9Xc3p5yxirUeU6nl1NOx38zZj2aL/u3EdCS/+h+3vXiuovJcTr8TFvp
gv14YWt90RcUAnIf8Gv26FAJhJ4qJPgyoBH/+9B0zZbHABsY5GOi9r6WTCvg
7ZNJGE/NDLLKEqF07USEByVTWxaFqxYGa/99jQHKMHwIBKid88ofBit4vAtG
xjcD+YH09Im1MxCwUgHZVv2/f09iORdFEymEXc7QfONjsLo0LgDLj/k+SSnC
Y7LGCjuask8Vxf6VxHW8b6vRWwuIybE8/pxIe7DIoPXHraWWUmiZK84NZitG
kBNTfIBHfUGZprSsNeWKXt6yoL1Z1lke0A8y81v3SUCHftySybaphpHTx/vz
tPiNIwk5oYSgVEXJU6aqRGYooy1UqcJOibtdILSaM/PGw6SupBtE3sWcWhox
PSHgCGrBY+WrxrKJttx0w0nNOqYtDaJqL+MDYCJLmqr28sqh7/S5GgaxVSFG
Oqz3rBMLVuQRTAr0GWcHOT1MxuNS7HeURWX5jnlec6Wf5yDuMs35jARtQDoZ
H6c0yuU+SkWReo8uvAT9kFgfMwSlYXBjWTLVJdgIirkmx4OfYqboJDtnZp9N
h9zfsfuXmRLeIt9EhfPFxALmDBihg0mTWsSQxBEGjJdU9e+rjUg7fQyTE1Co
gXKneokZPX0ULFP0E+16am/doSxzDclZu0tBEoc/6gB6guRvf83BQKiu42NL
Lh/xuQERnbsFpx1tIHZOCFliFScXpnKjqlVIBOTH4XInz3bqUynYs6TjMXSV
F/vCLKcEtHxoMBNJ8y+EiHg8eqKoF8BdqXFmlmAikP4ndQom4kpEZGFNKo26
eYkpr5a5pg/4UOKuWwQuv+o2gYiC/+EF3ZOgHuQZ3Lmpt3VrZBCCgHDHGWO3
0mzTsQkDnIZ5/MadD1aoGqbq6ddyKVEhqib4ZUWReyTHbiCAuVuLph4OWWGn
E/0yo3uXrDPPyQg8UHSOkGVjJrOBPEsL/rS4G7WkueAl1UWN6hMssv1tgVnX
4FgFwUhcmGhTeaTryOwugDYd+g/YtaG1icwhlARvNaYJJ9spItMRfr5iygbj
SvjJgvlbwTGi/QNmSvlzev1Qj7HrEpZTrqNpCqfKTuLQZBYv6OjLU8F28CFN
KTMx7QmYJwvKHxNzLGwqARelZe8CcJrSv8P8rdBq9liKmzY5+x1UNAkfD/Rc
p759fGZTpleUvShkURQHiW2rwb1mi/UZDGb9G3XgG5bYyiO+f2Zl7+XAR2Yb
Cml3Z2psjKV31tQP4AnPE/FSL8vbAgkdHbYfU18RXEYxvb4F4m1BFpWcQFas
4Mp/CqlM8IYGPFXxcB/qDKhl3BDlS/WxK6VRSJ/fZrYITJfQVO0erbc/1yPx
mDDZwpzOFFQEuzfglTpQMwwV4FaIm2cLa8rXT5JcMKW3yRwYixVX52CB69er
ifdmFCbDK9XVmX6JWCtfaHJXh3IfjfazpIE7OKRWVEzCrMvZvbb6rk3D4iuj
D3IWUpzHaHNGeWlWZaNY+zSKBJ0elRSgjHyR3qP5hVyEgq/A+35FB1H9fanF
HYjdu95XS2owNddW2L9t5x5ZrJCx5S8H8CZE2D10ORiNvssyoUAJVrpm5Rfd
epE7ky8OKsqHGlHdtoC03iao0XxHthgl+w/DCw7yxoF1rAG42cCe0zuVPdyE
XCdErYnXj8WT68KUmX/j1M+vwIXJajxNJYvux7qVUdEGIYlHr35LIuI50lCk
yQ2HTxuTfeOu4gaQ41wG2ml4k0YGUwOyl2399wwV+JRKRSveGhbg0IYGXit9
xDHwVbqeVV1fUt7RSyyz4RYl5FeGj37JLoC5TXLiDjqhZj+C+XmHinPiqqZB
xcZfR1j9Cgz9ETAMJFaBom2cEoNPwmgEUSr79YKVP5s/p9sUhVlaH5uVDHXz
MYg9k4RVNGNUUGBd0FfQEzTbgzym27Q+QULxtR70ciwuJlfKU1sn+Hc6x5qr
0dJIWPgPr3vA6JmMTdPGQfU63WaLwlLegO5bG91h4o/6KInAHp6fIAM7Ub4W
DMcwJNcySi9yALeWBKjhOyPoFj+30HTu/Rai/NRtyGxyZb6g7kfIbBZnCsiG
qHwyXRJnnzY/LnqoUtNcq7YGyYthS2l1yEXQPdXwUZVXyNCcsOtKkm4Yoazj
VFT1EQTAcjyeNZMj3mCgH1S1Snb9JCZnQgx4LM/3TyauRA/YS6jYNghNzFeN
KbBRc7TQl9MoM2CrN3wBcgQmLzReXzm+ZfMvwZESBID5WY6wJV54TkLw/bFP
esiYeGga3S8VnyyqwCj6AqO23D1yGplBgwNOm8jtcM8b+lkDwbr2biPAjMqB
TWXSyxVA8de2B8xCWZYC4+O3EtJYYMX2QMmHtAWcfhu6vG8NCYr70PvC5z20
ZFBJgEquGW+nyUgsq2FV6ISIcBIaUYNqnTZmF49Mruby+0qTw0Kec6ftuqLT
wh/uLih+QREaO2wzV6BduDY15geu5jXrY/PHUCFnNoX2eIws/yFc02B0bvPG
L5pRFf2R/iyCXNJZEKQT9icrYoJmj72xVczfefywyaTbErGw8qT9jbv3RSZU
umN0Mry6+gzvNkbrnPYLdi5FC4zTUYcuHSCF+us5h0QSkgpwBS2ZQyBdCzy2
G5o7qhfwaR1S/BnZIXeFEwVBDxXAZKGfnJGnfgI/YuP3NPYVyRVs/AfBnxlF
fo6cD86B2swNeAHu61ij/znla2Y0leR8Pza5/kD5KdBuvFuRKfpOGVrnTkw/
7/phswjZEOQV9dihKoy163ez0qON8Vvmyi+fNXi6FC4/Jpbj2bJ1Hdyi59fU
IG5htcDDfzpSiziLKv7+i05IUxAMbf4pvLb/p6+kBZkCO37FsphQ7h1cOUhO
OVNCnpKZzeXe2OSK7H2K0WIocdFXlZeIhoEN97+MoS5kjwXO81gUxgb2YTd9
A5RUEeo4XYwOsBebFeXZFIW6J1Sv/Sl9fAGQnWpGqABdvv3157Uy6Dmpg7Aa
J0z2GHBEfHH9f/E0O13nAGkyR36gzf14/tussrE5SHRhdq0k36+ZFCHJUAvL
vpLDSYJYw2qBOt1BvSo4MYmogFgWT/HrVWpudKNnN/XJRCIqZ1lwR8tLNwnJ
W0xOQMg8fr7ENMwj45hl1P523UGtWyGfGbPCaDdcdAxu2ahBue4Yt/VCkxvM
TF79l66/fcihlVo6P8uvJ34KAezcvUbQxlyu+1591gt9pc/5nQ+UTLAQkiiX
PvRl2XYJH1fsj0FwXzErs3iZfQz6yocQ7NTZnp8RK5zhrKXv8JRmit64zyVP
ZKGHM2M/02ASwFaaLW0sqzDZ2It2/efTEKGx/eVdcMiGdsQWcQGvKeHz9UGO
ujd/m8jAsv5s7lY5pmyTg88XiRYUKEvK07Y73SdEJjx3deTJO+N1iVwnaeqr
n+BCGblBtdI5k5duxyAbYVy2zWneR9U7XsL3YFPzEoTiA0xJZqkbra+M5wzV
GOOIAEo5yoUxpzZgHxvhnvnOp4Zbx7OFXyZwsT6MRSqy6C3RfZ9vPFxoyuoG
4b8HMIu8PJM78cW2vFUgAifdKU6RgPsNyDu+DXdzl8qwZLD0MMoNXVHdvTYr
rVAJX+vHbZ0Y69I9Mrh0IOc/F3dY/qxj94l5xsq8yEmCVw9K5zbx3w9s9dX/
eziYf9yKFyx7fbq+aK42JjpDNwdqpIdMh2HtUbtiHP0jpuC13ipnJcNY4V0O
r1eHPWwZe7YW6uVSTM5gY9Gf78KLQmqzuHn36TOb9DE/hPZ1bpZfWiXjPYPq
YfMiyUCjEN4ZaIr88cJDb8ipYrQOFlLhiC8fYDw0MI2ReNUL+O5J9epm8eoE
OTk8R/5u533C4EreK9qVeXYzAfzFH83aAO9GY2AfRNQ3BnwFHMdko+EKIDLi
4NiQ/8qdaHdtBNfLXgNxfhPP1uuUZtjYCTXUnSJllh3bYI6arp3aXZ9RGnM0
s3W/nuqw7yaDnZBg3r3w1urI2yLdZfQyuGjN9bpos16Bp5CJjaQe/poZnpUQ
QkQBblHzeVA6XlBpQ9uEnbt2FNBqK7P5j5ISAmaCAi5jW2ds5+8KP5kmOCu3
zdilJWAQomH8tCB+xbCWpEpuu8TjHeWiFzeRNJhc412nLEhivX5fjMkttVtR
eOvXew+ICzKtV6r3c6UPzgCC9vhnxmC8KMZSXOO/0hileMAVLWhFQf2d4vFq
82rfuff6/bIittGq1UUsR9NN2lMdOlZcI1NF0dGXQwCjRZbpstBaeOUxyUCM
xpQSu4aseKjDMBwwL9n2IWvJazZnwlSCMKq427ttL4AoobZHJBy5WKdOmzvt
6WELD2mNt1B4fnPOrm6h6RLhpMA7Ia/HL8wuUWffj7jskYj55Q+ogbtH8lCR
D3Ea93bP09vajAknvcMmzS1cOaRj41nSumJ4NJr98zlMY5C9jNHyfSDPSdSn
jJBKAKiIN6a16wybo5EsbEFr6XzQB0Vl7QVbjXSHwxgqkFBMhIh9jP1kTB8J
3lpbAuVWMYBerEDYfUadwyZqS8cptEJL8iJ0Pfnk7SxpS/1kzdfRgnegp8yz
RdP5tLrlOC6Mc9dyWhzQ/LOOCYbBkyqtYZCK31h1Wnzz5RShUDlX3wq+5V+v
xoENWR4FSVZbHoiWyXLI7sIAFP6UqASsQbsUvxHhqaW4FRAyraogyzhSjuMT
y8Q9LO0xAxeSfmMpxAjrikaSXU3thHawZdmF4myZfeqtVfWWEfXKKNbRCYgA
dpxji0wOSmJhuJGfDdCS+TRVB8TsbcY1gVlXDHVA5L+ge8QfSo74X/W2EcCA
U0COeMBZklZs2wvZEDJ38Hy7sj+p1C/o1g1iJhj2DSjj1/ynRW5Pym5Ratpf
WMA4nnaAgunT1ktz5i5oEYR8ODjzqgWJzL8zANAh0BVUfN224lUMZTOsyexJ
4/iyW0Eq1yISqFSBuBriS92Dodv0pepUl8eqp2jQ4DzFIjlaRklnOoFmdbPg
tYFoj26Bdsbv36YUYadLBhzsRNSgaiMNw//AojTToZomGXZXxHH/7nf0mRTS
mOrO2bAkI7xSkwtjOutMS80xsskiBg48EUmpHBy40D9q5ROIosoRjZojgFUi
fYugVrlpxmwUuhKjwlXbzknSx6GJw51F7EAYSqzfXnzFoVXT2EhDrLweZxvH
FCqLgy4GROYhfXWHC2+b2kK/Wz2muXOGkptIArSc3Gs5rFi7fwQuETC4JisV
wHyEDxjxg4fgoXCcrK8LdA64bJwj/59wvLOT6mZPxy9GavNKhFeEjCD9yP7G
vBAl11RomZ9wWG5Au0r1+0pqAxeIFUwcsjEoNoEcNLalCZdQ8QHAR76qIBwW
DzFH5c4SmQvoADv83PuKFQWdjrQcDjGZqHw/00+mc1/WmhVEAoOj0Eds3D3a
bteqY6Is0b1WEVKwqdOAAB4yIfj9jlGg3ouOT3JGa7DpdqFWQhSoXzbibKhr
3dj//s4qhKoDf020Ul9LxkABy0SW4ikpBMxVjuxdZjVRURXogg5SUbco03q4
4XIibIzXEtyduQwoA2anKqXyvPGH74eywz8BTsAQRRpTmmOhnMSDlSDvt1xC
Zh63w7fz+fzOnShNwX4v/+uk+GQLj2bh+03r9e3BscKkV/tyJ+PMbyO/M4AG
qzwXjdfcLl8QyMJhrCFjUzbU46ES59CKFNqwOPtNoGfRYO1TpTZO0bcIGPVa
4lqQQ0TVlkkTYzszhBQmaTKbjUZlPEOW6lJWVRnk5cbg+tsz8xbHcb4UJ25J
LYtebf6to6ZeG4QJAKowbndFc1YJT4fkVtXC0O+w+MkDNs0bUZxpEdnSAFfR
9ILgUOdd3ywKG6PFlYA1PK7owyVOBbro/8XeDgzIKN9X8EY89W1iPfFUApCB
A3GgsR1FS3swbFLP8Ic7yROoWAaJO1ZD/WR4BvR31fep7J2JY0tuK9QQ4+JZ
TTuDme7L+IIiie0SZ+SMOeMryD7bsULXfJsAfOQsxuoyiyPm/O11yLykgnBj
gHGVXOM8iKB51VCC3Vg2Y3cu3XEfC7zrhelXcjYyWgJbMxdb0Gj09qVovjEy
mTdfpZkxIGk1yEtvo+fm1eE3xtrGsx3zjNqplyiXE98ozIKA42wmEAIO5T4W
4UPgeTdA8nNiUcsC7etslceLojsM852rpDQU5R/C56lBgHXDV8uWPBugSzWI
QM+AfkmE6mbBVHMpRjkLVRhv4PnnI6lDsPWUxcFAi7G0KIpUf5u1gvj6RrRX
QcjLb/ZRtA8V5pLmKL9H6WzstLrx/vK+EMMLH0O4eV97zwrxB6q0Qtt6ngx1
gaHqwq+Yi++dVKcbBK4EwolIWkR7W5V5PBB0zFCu+xhWIrv/matCXXTlRvR6
JRkqi05n11XbJlO/MOKTkpZj1vt2vwA65JfXiUZtFzW+FvIdQOwoh5thVYPR
VGaA3K253W0+oXZ2vwhvQef8uQ9n8RnyO/dMm7L8hBunKnhxwyReHXOdAFTq
bcXKyPyD7ySZoNM1tFE0dluhfgTYMOfb2n66kD2O/rDqMpIo40xwoQh5TrIz
PS987t2a4S7DbhLH42m2apbNxmVBUhdqZaMRaSjqaN/j3yCbslix8YtmBHFb
393cgEZgspkdJ9fT2flUGbekeY/gUHRfEAbnw1yXQsmlQuDoRJraZNSInp3E
IilqKwlJCStBaMD8N+pMvb27VhX2ht3oKcZeyYI+0wZFXEmwMGrxw1MGH6gs
aQf03PQE0fNf42LgB9EsoI9PhtPUsZ+ZcyAUZKmMTxiFxX2j7I1pn0Q9poyY
TjUOFF45JqbBA7fdpJEdyeTa+/KZkWoLCZhM2i0T9WRdAF40Sp6ATYCKTHt2
uxUwIVbnyRnr7LWjWEZhMgp/uJU7ce685RbMS2YAi/nvGtzAA7dJAyo+oYw2
yqPSQpXmxLWVTwU4NMGIN76NGhwMlNM6g5mhhwthrNr9Jy1E74CTL4DiAqkx
J4CxA7IzBoT0Rfbxu7BNmP96O/mhCwYvSh+0G4HgipQR9YSiZEG9dBOf1F6A
gqUtrKo9CQvE7svw9PFC+lsU+QIkYZBTHAD9fBmE767rzTG+S1ulpz1rf9/w
ips5t4gF+A7ki5eH6Wv0Qpa2l9M0GsNQ9XRDfsb+BRAG43eXrJecTrdSXh9y
vuVkRHf3DeBtVZg++WfVCNclSdwU1CCaPofHD4QbyVkLi63p/RXc4K/5G1OR
V6iHkAIgYQrGQa5nRXyaKpwfKhEjRuAqbp2htVJLgJaQACezDsyOzVZTuQn2
uCsKM2QCUGAwkDiq833o+boFsNoJRDn+JBhoC5o3LItxJkP1PxJ84SJL+V7g
oLODSq/Ou2+x17hi/6Pt19NamjGwYfqX6ArvEk7Tul/h+39dFnLaLs4D5u3g
RYI1UCBKKLtc2EKFS2iEemC5v5NW0SXgHjTRVRKLpaPwKWiAHgoLFJmHoMKW
MXu1WhEBEmSkVKQ/YISdwfCYnMO9vDQ5EWmkkhyJlj1OGNpwV1AtToFIeqRN
K03fJGPHE/JACYHWJGO3oHovxYlge7noLNsNnjKQKouLbwS5gktVrmT3n4QY
5gFQg7BlqPsj1P+y3zAJ75/WP/W/8wywJb3qvxlAec/5a0S662T+G7yNehxM
gMZo8fMwJDjqpDtkE0WGiNOjZqi6mmwrlvnp3tfGGLscgteWblnu4vff1hSW
3STF7JJ1JE0dX+S6joqrxQxb7pRk3a98knWSe5xug24m12hkTqeA2mmDanlj
6ghAJsrYrt2Uxp0LNkSSvtnlBVXhLzLNlphX1ZvxTit9hupvQBT8gh3O9kL/
a21F6he9GfQVcsVtArXYy2d3bJIK5PFj6kdpCRh0hHQhgoqAnmORBdRbLFBf
XWBPPzH2d28sQSWQLylQNIF8w3yM74J16hiic+3Smvmaqx74DN57lvXzG15d
vPQEwFq3ZJhEim2TS+VvSyzaYz7hH32gcM4ZiRhTkwL/nAZ/wHU1KPDwGR6s
dygouOMPVoQG+nOF+ightr6ZzKEQPvy7J+Y0npwtb2/ZM5KlwGLh1exbMW/l
Kcke2X7S+J/KvJa7ipnp1h5GEJnc67rsXv/5iPdT5M3SMjWX/BsC3T9f4yUS
RhemtoNADBGR7ZLn7WLXKnynJmL7pcOW6vdUuWbELdSM7sVYI8KSMU+G5di1
yyOpUjOeeMl/li9SzmrmTFJt41yFRxYgvpZ2pOxl5n1RfqlTYxuuFa2i4ldW
rOmWe4rvp7aXv8QNCxk69dUtPoVzT1biEUipZ1VULG9eBWWCP4Ga3tXcxmbL
OgY8OcaiPzm/+XuH+wmXSwrnrQukQXchVJhW823Q1MVjQNfYhjsmKL5Siz1n
9hpGoP8oIoTx7cWN+IYm1jXP4StsPfR80sOViFPWzHed/koniiU2hVIgRcc6
fGgzGiqEXjHLqvQDWy65TeNrdimD3+4hcjjCqoiRFSiyzy3XuNfrTG1VpJkc
8GruxmL7eb5RYR2ViwY4Q1oJxLd+ogsS5H+YP0XylZz+gKVKFu+cVvfoxdjm
GXeiYRu1CRDhYy75QXyBidqRFOpye1iCCdLcx3DirQ+EO08Cu/OBpWz9Sths
9CPsZtDmYsT0CjR5HAsZS3MMV2eL35DccRlaYiBpXaQpJPLWwxuJ60ol9Cwt
tBD6DPoQf5+7SXchAJdwvBi+lib8OrSE4NboKqpDjteQLFUQ7wV5pLA2xTVU
GBWnx/xBc87OPvxMd4TD2loBD13WvJTTOPlzRug6c7xd16HfLxz279CMoUN0
Eq+DttZRFWpemSaKDxc9VLbME6A/9rtUuHncUaY9xl9Cx0pd4J6gDR37iPNY
TjDs2R+MaE4MtFbEA+4ICBr837iugdj4FdxhfjarvP8m6F7vSh+zMO+R4vmk
sT8sG1tKNSqlN+vjKu3yMJqXm32xzyOSKzyzSNQy3OjXUGUHT/TAjZ3zq8gU
+Keek0XU/cJF0BNdrdSMinsqPpoSBvj8gogFttQwKmXiPgHKi9PF5SssNpYt
+NaNJYMzAN0ULeKCADWXBZpixQxtLcgMh5P1fIHbKDOhP+Oh/WJkv/gSoezk
/ExUFzcYMNrTM1JdIitXTwDdsKHoqLdkA/F7oRJJUBVEBUsfQRkKMC4IAp9H
GQtPTFfm8si9ND8sh8/x88YZlmLA40a70dzQlkhJtG5a5q4WueVp7assnOLf
POfwTOKSXMKBUvOwMMoAPOTdSiKiZWp+zboRGmkuGtr6OzOa/DR56hqn8MpW
3okzB87gbFeul0+IAAdSbrocvzszFbVN0lxVhmYAZi2y2ivOhJNZ0rfgVZpv
2U9lx+qb8NMLxwe3+ZJEP7Aee7RCHtHLjeK5jTRReIVGQACig9DxhIDig+bU
ENfBFJGgOPZMJAzGnJLXRPOPz93VI/XTzSXmNWZ4SM6eaDjZCCybMh1gbkSd
UOYMSSnBq8TwPFvUnaLPQPfM+gu7wZtxYqTRZs1qsJoUM13BXC09akifsnMi
OwJuwPnWegfZhfZAVSFP8vM3HEn6fvg0iw+EYM7vZiZuEWQd8Jf03FI+9R7l
cVcA4/BTfzwXRWz+Lo+GFkHKHXg9ggqu0rlfl0h8q1gL5o62kIE+iBMs6dUV
r9FBkpox/PQbDg3CrUtXSJefAI1YJTWoKbpXnobm6bdJXsP6FdSJeTGsqt86
QBPttm1i+ZoIZ4RMrZZbdFvtxiBrI7PMmcy3r+q8lvixZZFHcAPj7pfBvoh/
lwEkO3CWT5r+izfvy5lEDyoOsbUmNBQa1aVx6DVZwV1I5kD+nAqCzzFcUlYK
RidS2Mme0oL4xZSAmLYBeCQz9nzURo2eeiLUSxRpSOAn2W2x1BYKkzL7OpYR
rO/u0xnsObVLFbVM3gGvPsoktFlTFeA4Jsrizoch8azIDgJwnJJ5/nfePIub
681RZt+GNa0EqBNP/3mayjv3LqRTTLOM1OEO5hh800eKNFITF9hh/lf2fUA+
pR+lQwGS3Did1bHIdggzPr2vaeXZFGFoXk1ErBBS1GthszM5WC0aAuvUePbe
5kRMr3pHOjoSj2bkIf3jR7fMx+Y/s+2o7Eykq6HG8W3l7E1U203GkYJgQGia
sdyP4DDB3FlaFLiCbl4sAEbkuQweJgOsvDBetWX6hcqY+88rjFz9nOlu0xUC
yrp/6vrj0oFGlwIF5GW+4Rp6Lf8HAVrqk5bZ8q4Heq4ihuwypTo4P4ih+04O
cTS64NXzwngXnqG5sd7Q27ilqYi/Qo+Ezjw1f+ULSGn46Fn3VFPSL+mtElUC
xmlKlffSOsa8tbcbjynuKNoCr8OgDnAvCK8Sxct9ZFaZdNWlYvnxH7pOXcj2
QMpN2uhxdgAXL/Er36klnGq7fcuCp4vKjaN3zBtzyicTUYT9ji6fEBupzgL+
JYHHlplQxGT+QJHBL7nNiCn7N8WArvi9JLLuje/Jsw3ZIbnBxrvgIt1TCEWp
MPbodaaeRkNvwkHG6Yk9rk3u7MfpWS76ZeKYhpojp8X7Za7f0+peTwj/8xeE
HRhh7g3JF1NSfYIfymSD7RXNPsVlBocyLWLOWOAOkVm7MxG7tOnPVinraweo
W2V1/7UAbmubnkePSbhcKzNFCgcSSb8UlvziG6UP84JJTuo/MRKC33NE0OGl
KNlM4o6UGdRPqgXg/PKtlKM4c6O6MWXZMDO6+PrTcxDAuZCiUpGTztPNJOHA
HkzkUvZy8KXEVTAOv3vxOnNqCbSoS/McYVZm7912kDhn3LPEa4p1xkTFwDO9
f21lY2F3jfCY8DdT6gkXHHqVe0eWp63ONkkE+Ss0vqP0Q5zxd9ALbJlYTaMg
2t0KyrYWQ7oUKkQ5Hhvei+rxVvtqzBLLiJnZFhZd67+Gs5Mx5AE0ZgxIlvMI
c/WoI9beWh1y/6BP7QFr78ihv5AGkwBNg+pLq2g0TNsuZxJfjsnDiEXLahr1
G01q+dbpR+mUf/y+SuosEhIKlq+IlJDXGmNjuWhZdEoiNdqpaAJlm+MdEjnW
LC/QV+kSypShZDYLGj41o0gHWLOLQZ70Ad52eGLQv1P+Wnebx2tkXDE8FFZs
B05kjJg9CuJZleW74X/aXMwRmgxifuRwBeInL3eojAxw5v6RKM+ikQ5dIIXt
RKT7AFUca/Y7AFHTqk0YMkVmaER69tcKyo78Ei2HhRZhhxbRMXA70zFSsXEF
sySX3rFDNvTOKHq0E+CMwp4rYf1NvVZrWTJMMLyE2gIlJYrDKpPqDKaoUaNk
I6hrh99FJd9zefn4lNvoxJ1JuSyKmEu234Q7SnCkSvjBHFxc5mPLbgp4B4wI
I4pKJIaM/iovkT9s9K2TLVr++9W8Fz5du9GkFQHU4AQ/9E+kxaOHKxI4jDLZ
FcAF6P/pN4gVqXnWf1VD0NKfJhNRZbJMOz8FVsi+MsC66mRC4VIBh8K79YN1
PthBqJwa7ZI5JRpEbalB5iPChJQTLAHr7T29mvB6+LGzXpKLt4YiNTWWvYE+
iJ3ENOPR+GuZibKPxAUgGYJ5i2zy+cxrDrMALB+X+mjYhecGbK8Tvsoe/2r5
z3w+JJrftafvQj61HUp2mYb8UmSCHmHO81RBkAKmLVjV4ACVGG01W2IXCryL
AxupcChUk/700P0nxuxHxMmZJ/OkZzX0lKKNNXlaOe7cjVJm4cSWXZtLY/M+
E3MTK0QFFQA0+JKWdrr/F+rObi2VZo97LhQ15cxYgLNnlBUmXUAVvXlwfVdi
5F12OZSUbNmHXiQ4W5spNE3j35SHod+FIxWE2QuUCyvUFqXrf1F+dVgHSoPu
/aUlMaaZ3AUnjpnqMcnseP6sDGawZyxQ0uFJbcNrTVI49KidLT0Tb0b6IT7h
4sBhkYat2cUDbu8Iz3CfUyG2fgPyIbLE48U+P0tzJmDKGFJ4f4DGHuKhzy7W
Crdi6Sjl8ygh2eQKegz0v6Gf8vRZw4IvAExnWtnjagX1fdGPAIs08cb9/2xK
64Y2wE8HMnVBHFhQZiVnHKXBVzMBnZ5A2lyGsNudtsj7o8sC9BNWg3455yuB
F/IDq8RZdW46vr0IsB2ZC6DpLXLfaRPx0G+z+YvzbLiCJByXn5yOlsW320K2
fgBONVcZySCp/eTSRf7Y/WXZhoXHVZTtb8doLuufUJo1z+8n9v6A96PAohnd
ZciI0t4m9hllf5JLsLhsJ7/RStDWrdDSv7NYXh2bwtQrw8dKv6rICwuz/q6c
JrJefjI1qO5BLIgvk2Rm10O9uRvNjS1el9MW4EvYGgMEtgm09T7pTPjZgJdT
4FOYWq0hIEHrLv8kacwYUL4gTL/qoGUGd3qbQBgXwZCNeLE54AhH5bgrq1yA
tEAxXuvon1wbR7jU5FhbOHCSBOTXOqW8cXxyKYRtuAOFG3Is4DR9pWc2foVt
NeSXO89Ml+Wo/lQbzOD5ko4dmGdeIU/MicuqEuvuZ99+RHTi1G49DjPIRXFA
LgGCjGp7iTOLCEK+S5VqKh6evnS0M5ypVDye5BGmgXawtK4T1Pd8w35wIVFC
175w4Pkd0N6oxEn//7rIJ7bbE3wkiKrcUuk5+X/nHMddHmr5csWyrJ3ibvwf
qWHi8WRFh71ZNGZfB9Ml2ZHm79voXOuIOaUIZo5VPXiLGesmLX7FPcF/vd6z
4SoNFsMXFMkyo+/yRkDjJ/At4rxn0+Wx2ETx21YlCC/2S6tiFJaZpUDxWCt3
lyCun28LTj+l1xgOGVB5DlV8aTsg4nt5DRjCB5xTcZZR71PEGidUYYT1A+GJ
4EA+EkMpZa4f0ob9eYWLVFLTCMeDZvrDUiEZtVwSv8UVSJlHgKNm4RVEJMG7
utENTULPd8U0KN5Fi6jWE7VvdH5idIkxsGljjpEvMOSo1gU6hwCZFEgRk3yo
14ZAIxw8Oo8JN8pDkecYi/2ms30NRfYZi9Rm01Z+X7frtfhox1buT99gpIap
vqHRpEU3Dy2pTcARUh14HGDQ5wwJeIUz6BzTFcyZMpemnEvjNyJSK1oXsd8f
dJy+4IsJ7jjOKAkcNQ0HcfbNDTHWMA1o/HHq1lcywRXS7f7Dqn4lVvxUBCJW
0W/YOiiSiZVJO787VfUr7OhrYhiDo8nBibxFzWBD/qxMUkHlab4/05Y8lOZb
X3miQTgPvgTt/PXVM6bt/HhEaGF4iMuumcAwjZ5oU3BTYkc4DFWt1SxE2Gkq
zjvS7Tu/FAjrdp8yg1zqqoHaYmPrx7O5sm1mBMrxEB4SRjlXNpRbufx97yeB
RCG/gOskcsZQyRZoKHv2oWsfVUlkZ4NyIzX9uSsaM/MPPjk6taE7ZyamYsis
GxA9JPMccLMx0acPFStfHG5WDg2T6OXIOBVMziyMysaD0aPHqbzBo2JVIEit
Ke3EJty14/zXgTNyOzYWQNvJZUDMvXb4V8e6k/6OShjnWPIxLR5Fl8rd5aJ2
GghaosEu6GDAiS34z4RERYg3IDTRKgdyy+whp5UyRvlMyLBhGL8ZO1TqLqKw
NfwlQmFuzovEQ8a+ueLv1Kp3FuSc2A/bu8mXOGeIYAseHKGLbWzt9dr8O2P9
U6XhbFC9c44KtO+UsSzYacr6wgUY/k+eabENusNLOAkukBZVK2RSA1ZFrJnP
tecc+f7qTYdMNb5jlNh1TFjS4xHgsEr8x+E4EogYMvW/AZfQTJuWIVQ4sT2w
UNnhmexa09u8GSkdOeOnAB1LOaAe4Ze0SP6YOy2DpbTT/V+rcnuCZDgrY4gD
07YaoJ0g1vtmRAaHRBbsXd2K1cutXdS6AOGOrTa6E5ChF6xGqPn7DKM7k2Zk
Ug4cdYAOEUpd+6rrsnPygiwcnasTWGSlaEqUm7rah5r3Ml1hyNJ7rwgGYUmj
sZlziO0iPNgeQBPcCfjb0E1XXRscY/tjPxwj0dtMnvdqcohzzlo28TNIIEBu
82bacDHG3YEUMSeg/ckhBAYF1K39G/TfqG5ImXgflnD1sx1yHmlkjZelzqbs
HHOCTs42hyKVtBD2DiS+UBAPcMkt1N6zGjDc9fca7CUKtsL6wouK96vJVBwi
ARfonS7QsNMMJL3JmGmTTcgMPj5kwLgEwWQmXp9MP6M++bCC/Wx+05FzV1R9
fXh+eEMMDnD5LsqsgBJBNBdaMe468Xceod9FXSlee8nP4qw2pz4cav5DQMti
SRR5dVAGitzRN4lyQPCDd644BdSf80xSsTFxH0A07h9HR25zYz3vFYYu0dyU
GFsVu9su9r6QGbVbIo7wfHCbvlhEXJUdIEr3soJ7Grwg0mKycnKDFF81eUyi
JLDjbTZZhj64PuquTtR5yzPr5BcjTtbHFD0NRIyzgC6SQWVOa0Lu/6F63Tog
Y+kQNkpEqIU6xlcw+wmQFy/mJFZh9i2qJQfd5WiAiKDBjX4YsaTIUYggR2sa
Nrb917RM672ZemKhOuKLe98PFpHPJbQ+sfTNsQEQIqOe1T/JimeDwm91e8QL
3UVD2n1F0pD3AuKbHGR9NRKc98jnb3h5u5R2rj/GXkxySGEvkfV4qS24+G6q
/UkMuAP3H57kq5+uTYaVWqHHiy1GQpw6e6q2p7hydBs8FcpFVvVKT+hiTBb1
GN9fVS47sNkybWtpslROf5unJROAPn0GW3qfAZHeo64EtZtoxAyYsPhkR6E+
hlHtWSy6421lGmMoIMtSm5GJXnj6Q99LRSr96CCUWP7xKTKYvCB2gz0Ylnnz
4r2aHB/DQRybQPhIT96O8lGU36VwvD17TIv9LIKjEC/yedSSIRUaCnVE9Jir
sD+ZiH2/nSyLantHxog1gCwKoUSN3PB8nlZqBuj3XJ/x3FtjFXuqwlbbxN06
LCPuXOe65oMx/ie6b0TIYWsOxp6BvqYoYIGm5O25AM4rgtou1H0CT7d1YpQI
EQlSUuXaf7l4Ir+zcCw6XnQZlJsgyjYVMP8/oHajpXbnqzrx6l1x4XCg4glQ
qNXV84h2grznxU6zLv7iMa+0HhrnK4j8NxU2jULahy24Nnjeb7uTLAtzlp+L
NqxzUhcKc7um4pxblxQm6oeu6XV0y9SRzcpTsbbGE3Sa6Qjsr/PZww1bmgUI
GuSvX3BjP7aSAFRavP1hHwcTnTuwA10hZX2IFr83dcAGMlmZBXtz0afYbHYS
zEOcrbA1w1v1xwFOV7t0q7UhbzUnuTv2hLzG7DJU5qdDS/eD/QHntef7MLbj
7Lb8Ns6VYP2BRgvfu8MqxJryTB0wk64Pd4o8v93jD952bbnFhzqVa67W2jC2
rJc6RiXtv/fbemaRLkfxqQleWWo96h7mMTw7cLbaX7C5mLMywV2GjZicXFJU
r0KxA38R/UC80kYxTD8XGgk9XhRl7oqCNX0im5nkm3ebC5tvSWLZqpvqI6HT
85Xc439FHLTlKKJ+DC44GeBMYZC6zZ8xAxSWGF9d3lzK1kqkdSiqWFHbY3uD
qQwzIB/rcXME9hFOAyf+tHMfOUj2Tr5JEj7/QA2wpd9bT1ltUnFivbSX/XHW
ZVDi0YcRewU7mhH52J89kMppCvuJlASNP+u5sDE6rj62rRbLh87czFxix6IN
2RT7AGrHa8f0DRB1S3WsIrn+t2KPZvG1+8YEjRrehxv+9fTTx4J20pt787B6
uhfDpoNv96GdYc8oCY7vT1EXczeaztZ0kNxNI31MRn4vFtfqLWfFc5UrbthZ
/eNU5zgVYq6Mj0a9Jm6SWFuF+sG9RZKZMcUhWeSYQ/6T77Vb5esuWBnfoDkr
DoABNDvpH11sYfdiVHfHdbuRX03s+tGlD/0lWZQjHj63JCJbn8HsIbBHmKh/
kAaUZcxchCF0RoGgXXN1liFdcPGPkhKyKfQd8NzDtpXg2/h6+ZhDw4+OsT6n
aM5AYDxxoz2D/x1W0Lcyfp9KPKmDTEtkEIVjrnwdMfFUU4yjUGTuTcvotn3O
IXF704W17wEzRRPeH9LJszavlNdWn2dx5M+G7pYg/Y5BZiR9YG4b5l188Ql5
K1mAURRi8tKA0D061A0K8aFsNZZvICE7AE8/VBICOKNfHNt+PO4tOae/chbt
ZQpPTo9kqgvo15H1c9V9s6M2650SJiVAYtQ6YSeKj+smLzeXVGhlVcdl8lqY
KgD1OMGicnWWZfwuVF1rLmSPcKdx3sxqUzfyfSXley8VfVAUr3O/sCR9Dtcj
9e0E/qiK9R1vf3/vQX8zVXn8P4kXWMQ0nc4BfkMNirxJunt26af+JB7Xitm5
n7Qd/hppWXdw7NHbW8huJTJMv8nzoiqRegGsxpOdXACRni2HIiW7gDEkapQW
JsXOWzO2X2dTrxJ4STQ4NSr7TFVRNCyZLcBCXWZDMTH7dpavs/pY7t+111TW
s21XsDJ+W0ED7OSaKVkwvbE7DOfyWwx7aMGUDC7mz1ty9PxcsPZPscbpsnyX
3WEJQu5eyHTnEZlgyJUcxDM1f5x5XukzRaJ95rNlH/PmO9BfBU7OeTEzv/pm
hDrugr7G9mUANVxudcom4SgX+9ndDnKqDP9zu0gLdZjBfCzDXgH8P+PGdAkd
9Cr0iHIzTLOo4v7C5OAbw6xFRG3kf1lBIS2HZ5OECE1yuNV9H0psyRWhnS0W
KkrdVA2zR+V1OQvbKvf7RqgQGjfrbQUoEHHauPQnpTS2wqnCWZ641Cl7A8t+
+y/LQfjNmtUNbaajCjcfo13tFpvi30xW2XUAWtsnN18heeHCj60IW2ks8ssH
AIaMJmFbr8jdDOVCkLkruODj32XNG2cARZ1NgP1Sx4pw+EvDD7ztQvu4wGEE
QR2BaVDnc+SbIbNeCH8GamewkzwlzaArOSuQhJQgnnO0dvH44nbzfS5cDQwo
0WDs+HcBD36iH1xZqqyvfyi9TDqqUecqui1pl9kW3/H8IX8Z07Ht2KkqiHdR
nvhvQfnuZ7YM83feCC+KYxGUSfNGzXyy6T1hUQBRIsvuPYPAEYvYGvZCZinR
+D63Q9RRgcDAti3w2UKgxCQwdGJvbOEjBG9Bhe/GDna2nkdQzvabhEg/7dXS
zzMbpGSESPq62Wfq7Gu2XN67qkolsgEhaX4ONARuOzFbjh1NpofkJgJL1At4
gMGPcCaYP8Zk/uM8DDeIQaesKjA2zcpxunODGFEEOwebfHcka5N8X8FaZ73U
JwtJ/DLKDlH4Jne/IO+2EY3RftrphuqQ+0EKlUzISe2CozDJvckhkNE68k2z
07otoPkqiWa6EgFbjoycxUhhzrRr9X9kAd+qgFVD/MO4cgZCwDW/yAVARlF8
zrml0fsWtR0FCNBFro3OH5MADXGLG44utTJaqtNrYIjeOltbRW4m4u/0dPtN
8izCwXCytJyk5yyDGFL+jiNmvT++nKOnZTEDgXzmDuRJrGzJjct+oKOp6zd6
vI5b1jq45aJuJN+9xybahzcSCB8ehSohk4zTCoUmTFVl6nX+/k6kOkskxXp+
6vpukw8cBRXoor6laQmyfJSEEPJiKqI305W7Ucx8VVvsM1Wz65ubLMTJqeI6
UdVV6sEcMJddOEtZZlq65TaPN/QVIdMPa9h+tz2ZgaWTM6jS+r1DyT+Zg7qM
YrKWbbqhU0tTvBJYL+/iaOSFe/9IOItTVllUAlBfuWOjfIFs6XWTHelDrxhp
AiiRFmRzP6XIPD90yaA43yHGtdw3XxUx0b2C4PtIXzKADxgwLHJTYZDzpVMH
tsWUPX9qGlOOvNJtt2yP/QLSFp5/KHBzWDdPCYfSd5wZwh9q79zD/BiOEBNN
afaic51TUMMvAxBzGX7vtv3cAToJPLAkWqNuMYrDL/rI1lY3BgU8iaO1lX3N
X760YP3MTTGfKaCQqZktOTwYaSzbyFCWuqzSvXzjcbfgzitpY/7ShDdVwGOb
MAkkyEmnOKKzH+552dDoQVsyBmSVu58VHWyaJn4urW94WiCy++ybGotqtT0E
gTjBd5xPBZUD9QIQ3kSROkvn9R4he+TickNQQ/XNuF10/cghvaIeUISaoN/i
K71haCH2nmlAFf07zffAoi4XSEVjMZnEZEi/PdA8trOBwwyGSXIofyTX5hyD
u225krjdosD3/vPzqw69jrhH3m2OHmMjxnxDsnIRCpeiTody/13QnUJ3IH8j
t9QbAz4oUP8j1l3YYOBQ9+8hf3oOFWXSTeaAi+e+bc1KK21HmEgztm4niInL
f1F6sXzA1VY2jeUUObaIHT2qNMRGs8n/vgm0vjAPd+FMpp6rVp7QxBpAwyge
IZx4SYAERbAkRYOBQjY8giF2jjzzX7cPLieZr4rwZlTVYsYrADKJ60yACXov
+3STkC+7NwNHrm3aMKrrHF5eiKYZMmYRV2twerEyoIdFwDiGVVmVyKp6yggb
4L3OcbftvDCC4dJI+9ccVLxifHYnx1+VjJlmlwP6RzQV/KjmGUwLmrcmTtGk
znucowNJey3ewfjZZIv8FWBUqtcfx+K04/ce5Nq4vjMedVu1qGzn8v3bIau6
l6blryQGNDr/RSvo6rHzqpRM76o027gqQQG+HCH5dG0ep0sS2oA3B2MAc4L9
FSfeNMLgZ/BprQqBRL/f+ZUKeLVkqlfV5VYH40AI8fxNA12fEPAO4wNRYtk7
HPEpA+jqoZAdTKUQyTOGAgrbZ4DiIiOy3bYLiPe6stAtLSbGM6xquEXJ38Pp
8/9kCGnen7t1YJNAvTYVnfmGRERnp6c6yJVA8IxMLgAk6KFyqdR4ZbV53qyW
tTF5/DDntok5LHVvM9PBzgpgmZGIVXNBmy9TYdIHwsKfc6JAdakhvXURaoDw
ZTEKnMPSGvzIjxXJNP00DO2rwyu68CYgXjcy/RcZfXjN9VBBdXvN9DluzRwP
nr8RTQTadKEGvTCBQeVAOFzQjbsY6ipQwdkOnpuYJPirkffkAkvnc8gZgtKI
B1FkE+7Z3fBfEkGavIEF2sKBqeiwdbSBOUocKy+DRS3stSooI0+yE1yiEJC7
rsF9s0q9QLvQU4yPQMUa2iEZYyLOV0n1fTpFogVUj9ANz/+NkS7rwrNaZjtp
KuANueELqYxNkKq6XagriM2OAe/7ov1apVls/Yy8Zw7l/h4FRqbVRR9DvDoh
BQvqOojQTJcIwYMK2/nsLGIy7TMiy2Qg3CqFgWfve1OHWWeIHmXWnF45EzCr
RXgN7dfACwSmLk/VlIPyf5hUbdqnVBS56l8tZsVCan0/fDabMDrezjD/pSit
7I72p1yFx4Ll6OI2rZ6quNZShmvIRfk2+po21Ir9hJCPNz5TVWKe8XPqItoM
10CcDFXNJ9JS9kTp47/tXdV5YyAUMLSrQdMCsa3LSVSV6ytKEuMdPynoiGGq
A5FHiAau9ERBQ2FvNLtZtJhhUfTwDzAtMeRyyX6MPzJhgDdeCZdzMRet5Pfv
UYXyfOGNWAxL4p7lRJtDq78gii3lCAHQBEAaJ40Rpen6l3/xEKr/+a3bdFCk
K/g4XPT2fmyplfNj73R/goVnJelr88JcnbeyDJb0xQvwBx/5DfnIy5i9rhpP
STrMexbZCs5AeOQKOedaYHnVb39BbhvchHi5RjsHK8tzmHbLsVM4Z/cp+bxP
rNRU/hLjVm3bAH2EP0sRSr6ZB0CVuEqQ509WYY3ngEO7hBdz160XfNpbwRiq
kJpO1bYotQvgf2pSRXZONcG9yGfpV4eQJwl9JbeQ33vv9sVGVfPUkgzt46JQ
LOWuo6uTeezJbYe083GLZ3IvnLE9NkMcuRU3oO8VIKJXw0ormfO5Z/NYqofd
O6QJ49f5xPtb41rKI5G/WQ3rVVuL1R0Iyx3AVhB+N4MFnsf19CYSvGYIFUf5
fyQehaQHGGNgKLGvPLhbiUMbgauMk9927ycIRmbVf9uAkMvnR2YZZJTkzXQs
I2tKdgR59m/VFztxrBuRtilDo+VVvvgUJm1jHfNQum4a5mTrPRaOjlYS29nt
s+f9bIjo9ekOCGUnt9rCflDGLv/mpazGj15uBAHv2h1SAPY1MfffNZkjC6wf
2OFblq6ZQOrHOdUiLH0eRv55Q9hk8KdZq+rJ+uizht+hRVMgx/z8nFg2j9Vq
2izGZXDtaLStRvzKUrDfXus38hLH8fVKa74Xcj1vu/EL0xHi4mDzepA/w4dL
f1YkbLsi0KwfflwNFB/SREmh7slJdKrNICdDMeyysIMsniFnLzvvY7rcslZk
baDGjBHsOIpA3jXh9PM3WJuex1kLKDb5/pBZzhu/uhiH2NTGb7pdrBwaUmRK
4N1LZmSBulpYXTTpG2ldgz2E0BwUOZ0x2xUOIMffYjtTh65dAIDMf44vvnSb
snVZzrEuUMqsMBJaTeVrZ6euqb0yRCQNFi4OdXfTfOuMRGZnmG2nxv8lK9uJ
bE8RNCDR1ECTw3DfwTRS4u3tSdsqrCOjIs2uXrBWm2OPW5RRblsuJyiqmsh4
SJ1F/oC60hl6QiBL/gm3jCvd1z2WbNwCjXoLkHcUdsUPclzMWMqvSWvLumEY
oJNbqDIVDKwAIgF2wI6vq4NLlm4JPVK99HI0hL8pmOKfxXkBkTB6cEaOvJgK
jTaqEg0L1Td844nZaOfpEMCtxRttiyElMGstZtvTbLSPbAjWlfr/z5/fOwKf
edAgzkrUeSL5VyBdvxZLdoAd58tQk46C07RaganGHRgiu8yZ0F5xgMTG8Ppc
VDawUulPQac2BJlWpNbLhKuAuEsG/8a33m3trEl1W3DBMnDe6Gtmpvsnfhor
+WQF45JZxuvU+RYMiB7KLmNbGeNIJqs0TmMC+8dxYW469V7XqvT9mVKFSMzo
il4KSjPPFdwtQTfoGavOFicbMa+wExwUQnSn9UEleLECNB1UeZoBbQKzG/h3
rskePRcVrgr2n12LrqbEg2bkjG92pa1kZfVL0rZ8cS4lHH6RQVjxk1+GCnw3
7wx4wSkV54j6jV0HuU+k1RXf9kHgbxxh88krkFrbzeXcopQvJ/uygR3tSHPl
KqYrW+9phb/81mkTdjjR2D+fXvJgGfYXfqr65LLvOuC/FjrBq9A1LMSHPTPr
lUwNus8fSURnytOfmCU5bOdu+rzHxBl5G+XuH9tas3NrnVUzvqXXJrkZsq0y
DXkjE1yVBCFAjtageOElH3dkxgV5bBAvd5mVgFNqZsVNxXjNdS/k98XUMg0p
02Nnfh9T3NpJ1uXMXlNQayWdl3ceYf13DJcuis/fTFc7Q27vVmYAylPUxCnP
1E4NtwB4RdBQNGcK19OlEPvepnXPdWLNkY0SFfH40ZDpJVb0Yhm2f9+9wUZm
1KDeq1Dsf6i6pSeyM00U1mj3ge9LG3UfMY1j3B3QFF0p/fl1aNK28kht8+Cj
q++pYaZ0tRLKFo18Nl/Au8nYlN3vrpfCOvOHyl0VwZnfPV35KMD12sD3LzfL
b9en3X5BZ02jX9VVjGQyzTSmdrQSQ8EtiyGGwIzH+pRJNKeFbS2UHzwDcvdP
8QZNofd/up3EoK/dbYfiNQTVlwjlADYR/8ShmTpmvo03mXjqMnB7YxEL5mS/
4wNnFLVj5z00ZyTROOa4X4lAcDWsXMmYs7RdvfCHZhu70Klli4JzXvmJTyq8
RUpitio1+vOu83UsQmd/Svr2r4ERsXqxKWswnZMaE6CtJgdoiVoz2w1mBa1P
p6EouQrZGljHzDequAzPOuwTgSBx38L1sTJnoZWY/ZLidIiRY+HkX4CXb1NJ
qIwd0c3KFP+TcJmwjlaZI1gIV8B1vv43PbjzyG70fcoV4oyldHESvz5XplmA
hvRrDa6zn1NdebW3aRXL2ijUElAAn7YjJre9wSArfJuC+MhdtlJPzP3yfy8p
UdeNOyUg9LrZvLR/owSeZj+DuQd1N5vEip8LXrki0kGpu/6aH0iDxMTf+Qbz
PA4GQRgmfkgt6YyTGzt5J6e1hJF7HUuglDBjvcEkQSOebfNR/j3S3+coIqXQ
ZodhvDQUHs7g4NhQGErz073Bfs5D7GgEQPypmiMkv6DrRyyl5J7hhDLXmeBZ
6rGe2NCoJDBQ/I6UMQCHb2w6OgXXO9Ni/aAWoH5RHuxlJg+zLvilQqXakyWn
w3Y3OO9eVe5jBHEGaWRWEMtuxx8zUlYk3hCcSa6ATZWopOJ4/vM/XFezgxn3
l3TtkBHKU8KbZxOgSKnFyQn6Ssre9ZQIT62j7o0o2jl9dGUa93ZkU68vwKpz
N4MtiZosJ0D5oCAN1OxFTZtUnyLdCBWXJdg/N2KIsSKrJMM67xDFnXoN2Q4r
socUpooLsiogJWDo9PPu8g/oDLUqeW7RVu29qNPN7l4Q2oFyjGJkbqv90xTW
nkYKG14FMv1iu0ophQAS8Af1rW5qqHrIttit/WHu8GrPWUafH7cnnoVC49hn
hitb9e9E/39Fl96T9w0wwA/cGurv9B9PUrRjQxDmPfgPLpC/w48skxT22BQg
42Mzq+mSBBg2pZMibpgU/r8qqkTpsjJ68iF0zzc/fXgEKX5liR8fq8+zTOzt
cUOkG+EESRUU7zW8NtSYV115V4LcK7XYZ7lm4bP3lMBkHfh8hX5dcWnKFWPz
U1qS4A/F7dkKeLB/5fVomfqk1Ar6VW4X/mZF1LS9Oa+wi+GgcujJJrtO4EvU
AH+NqpelUS4A3X7jduYFBUvseH28GKBMRth43HcS6OLvj1T2AMOWyk6RxeZx
BPKb2DCkSZrXxoc/TCV/1RZ3EAIJIDfjxxvYHM5ek/Z4cCJrMr8YvGLU4cLX
LmQ9rInF/hZcl3Wkupc8S/xFdjhthFSqiARK28IihswYfVs5JHkRTCYDNLO/
1oUWdPu9Sf2riy/OD5oUVOonRcJlRJU3/4O/+yCGjzc3w+wHKXDs3TBM/oXK
NW85lPJsiJoxAymU4+0+XYT152ELSQTDTDy94xwz8anyzSlL/neeMXt0WlvM
2g5SlaUcOOakdn5H35SBtswBypsHWMPZ2wlvoYU780TBJ95DmaXrmPV8XEQn
q4xK87iNpY/Zx+pItHDMjKl52SYKOMaN8IUJQbdu0QXRGSqE04BGLZNWnkBC
38BJVU8HOCHlLMXGeEblCWSsx8PIKqg2uXAUi9PCd15WR0k0XjpmGeNogR5i
Uz96HakC38WkbXIO/nkLtXrZ4XGDn1j3UUfb35Z3IZoOoXrwfmiLlMNO1OkG
j825Lk08GLp0OwI6nL8nlOeMrBiopqYhC48uJtGQ588Np3+6OK5y/8ciyYFS
aagZOX5geFGWlQ5oZRIh56P5cwSFUwJENRKLb84lmrTsAlmh2LXyQNFS//7c
boWA/lCdjszN3/MyB0p8oXCkYnAqEPeSup/ZaBbwFp/EyrM4PduYnI5M1/k/
zQ2l1BhEJLuUv9R84nmQhBTjF5Jf7BOfKj/hU2AV2oYwyAltkVXb58xqVevB
RrFqAr/iBSK64bpB3Fw0tVdJ2dGd1xXWs3p8+Vhf/FlKLTbG8iAhHXfgx63L
FklkDEuLAzmC62oncZvL/qaLF6FMp9+QIX5rES5JQHBUBjCumfqHJghytXb5
WWFG98qF2X1jy0lfizyt//C42+q//xgcGKgjddPbNDCdq9bDY7fSj6ec8+HS
a872dYVxFcUQ6P9eyjb9jKF0opaDn1wTiFN0tDlMN1l5Upj44Qj64GilGha1
26k8uLxAEUgBU1ziqCfCnq4yN2n53TkrYDX7UiTtSLxO/MbD07falRCNEY75
3N5aQiqnuTjSYhVrdoxnCXl/Ko3M200mrUhAJ/G9u0dh/bwTE7nyxZWNuweD
a6ojfilu+xiFvzc8HkrJ9tuU9KoLh3jxCQOS0m7oW98Su8m3uWyDHazc53Xb
DyWfBeZAeNXUFzQNTxcT5OszrgTDXBCDE7Btp/GdyQyJFuHH3u9XjHSmoC1w
LZT0+qFvXeobPV9hFZ+LQm1QxZrBwjIq75LCHLQBRJmTiXP1IRCSO3As3Ju9
P9k94RvW6nggYnCS5hOV29Xdh2szd4wKY4ffe4OA8ESo/cAQn5ks5GdbkyKm
8w64ZgrXAixHrK6m9anfyRSxycvWw4q9KUwl3W0nOqnzbeMpBMqx1Ft9jyIS
fYd8cqwWyb6/Ha17x1GqpDVVb2Vd0taDiEYXckGd+o4rr34DJ/vh3PQBZc5r
3G54JW6TOQBYf77geVCC3txKD+UzBBrnm4qPWSFrkQN8zZsOP1dWN49Z64re
aqOx4Z8fK90Ojs/1xTZ07f4CjkBahwW+moao9MMHkFWzFc5nSuLxdP1HnPzw
bsZTQjelfi6xp6v5YUS4u+Fr+CmV536AbAeaAuCwgci3nJ4LoMPjgaYne1cf
Hfv1wvd3/NboWnr26TXW/jHcmW22AEYqPaZBc0y0W1Hydz1p5ssHl5n59IA6
OI/WZajVH62N9juTE2a/V72IDFQSI66XkXawAZ51dBBQs4xJIxJIeWX5imsR
3fKQO2LrQabPDVArKYJJQ3Se/UjoEHkgEUWKsigGBe6otG2PmI0p5oHedzTK
sduaXl5TCyKgS5nsnFVGqfALC+fCrQCCsQ/TXoYvhv1WDSHujjpKTHWaq2zU
KrrogvhQOtLF5xMis9vkvUYvZhJ5Q6jVCQ8Lbebg5oya18JIT+GCLAyr4oV5
2NOoe6l1++gH20A1L5Le/us2NTejZHq1w/yAd3+KTszx1iTiZlMFYagGdqJj
6IsQwKj8lbVu4cIVeSNbszCCcFIDQRMTVh3she1MD7+6oszOVy4ZKh+BSsLM
+rHjIRzY/STZCuyl4GfOXE/FEuLf4EYE4AE9P2yOCYWlaLMNFrDL9yADAQWA
0uk4IDfDf5ysZdgfLRgS76TQyUlFjfwfMRPDdK0zqokKHMo+cgJ82+Hs0/jW
opP5sryqIIlYfDtHbcQcA+rDcmHmpjBdDNh/OiBucNFsRcJTntfdbyFFNULv
ZNDDEFhRn4rvpe3n/1ciopImGm3hMCLAgPCbdU9fNzWq7I2fY77hgwEzxyyp
gKc7pUVVC2Luj73KsfM7LgNWt0hwDDvsx9KCa9m6NfkLfc0J0Uxrj2r6GO7H
j9bGd8tIpWpisSbhTqRdOk0uQeMBci8WWVIKYR7gZO0NIgMnvUuAuQpz3ZSN
R2nEg4Wk/wP+KvSmuukQm0PietQO0JKNEzuz79pIjpWXUMvSvDO1MG7QhbV+
4WoLw+nPgFmJQSZAclMkRIfOM//xuH5UvpmJpsqEyrtAbV1U8qFspPSy4Nhr
1N4lGVI1daKVcXC4xg3/3a1ycsotzoPDa0PDkCA0oJIFn4oGvoLeL/2FLyJC
ZmAfCGN/uLScFHk+StbCy+SwQkA2bXiiCD/zNk+gDC/mvrCH+J4BcXyXDltP
CH7KJ04+Mk3Ha7kXCF4C8za5eGSfx37zsez8Yjhe+hoaEoqU9rVa1OoBCL1w
rrQ7GPLbY8R2SiNsjjZTOEOG+dBOn/MulIF8SuvWLsb+pEORhHqOmP2LdmWM
B5TpzmS2Xt6aQrAUAE5kqlLdyo9hMOHP15c6FI17lgMa8u0ENfiZgyCkASdW
U/v1hGkYlz50+1fPYm2BTgi2Rkr3H9XLKM8PnzPyqfpHEPx7OW6IoiG+83WK
EyfMeqHZaiE+GiCW+qFax/eRa7Irw5mC3u9hVoK0PYAJ/0HQ88dikYj3F2jJ
WpgImsn36330Bf/HNKoKGP6pg3QXYiq6XHbLyB6g4TD3ZOBLIZ2Wj+gWPWeK
e+NAr2u3G6VAznb685cKdxXuXykFoIHEuDyF/CLRV17PXCutvoZM/mPR8FCy
2xoqfGClXItT6qZpjeqJke7YRm/xjAj95UMsHKLR6Hjl9kwLXQ3a7ykdUs7L
LVJt4RdN4KsiI7nCGuWFGt2szuyHNdE89ZHtecRX84mjdstVHcfc3y0kCg0T
14+eGfHBVXU5C4Onv30uK7VQV/anmNkLMeC2oSOaneHAKvWZNfcNpOhu++/t
a+uzM4q0Jz8WfAgtkvI5xZCCGzJZNdDDyRLVRbA/hyQXTo3LvUX/obXVFlPL
tVjw6vchZQG41dI90HLrbOh0dYOO6iJCzenpM3QnP7hRoS4HpjEmT6gYaX5E
OoEs28XybdfBA8C/IsQK5bR10eEBsHAZxNhp5BxV9ls37YUW/SiBK9Dh7KVI
wWIVagqK0OuVHpAKhHt7di6KP0fVT022s5DyoKmauYk6RP/3nK4Q1IlqW5qJ
avuYgRKTvx7gV+bWM9FVOSRTjZY9PIWQVjvBC+8zNfIIkZNMa9tUPqjJlQ2U
o5FXds8x51J5cOmaAJSgIgEmI5nBKIclnXEobQ3yjMyvT+CnFIsWVJpFGuO3
uq0t/VDNeqtwrp5Cd/KapcFA17aLrGLtJjdBr+G5Euz7fyL1E/CAqeM5JY9B
HiarfrOS8Jzk6/rmTJKKQGtXrLHR6BKkqV/jdHOTalkPa2ZWoFySyoissgi+
bEzT2/OwZpGSCqC8QQMxfHAxcPgwz4P3mjlq6pBB2xr6yAT+ayWwYiUBOod+
Z6j6q/XCkk4Xx+u/ESI9x7zza95Ml3aWyJkDCisw54eXmh6b1PX7sUx8kcXL
G6GRGIYLsBuyF85sOv1EO/bn2PG+8GJqyc+dUxZPyeU+UeKXLQ0CW5iMXAak
lQA6q6iuBRqmPmXXsbZtK7Hyst/iHpCAI1R9vzw43IOxGYuQwZLqVUzzFLYx
yTOAe3qRX35/HwguJZethS87jTM4qJkG7buzekK1sd0EF19HEvbr7LrJel3E
vVuq0+UXpfxXpPOHp0EoV29qGfFSkrUp/1HVOVzmv/UHrtWN8XO572I41MUl
rh/f5sJtjfJYQ2ja7sBTeIFOglcBUyy7Ig1rKrwKNTWs5rVnDWJO+2SY5YSf
xuRXQ3PB6y3eVnkMegQb354qaw51EQ6HWZAjfCPbtW11spI9VcO/cg3mAw6e
VbmrP+CmajAN7I6lwiHja1TaEltsjMcKAmeTnnJWD1wrnShNr9lym7o96An9
BTFgY1dgjvTtVSBk4s+wxmJHud71+sX31kFdherGgiHrccoilGhFyW/SeX03
yC76OBslaWDoIk6EDfy4Z8Wz8GeG/CkYoHeiPawGgOeUugZl1lpnCy0GnHaZ
hXj98h13rGhZuzdmxBRxMpJvHQtPK1Ssh/dUUCWu8SdR7TUFt9NyXRnNgG2Z
jQRCN99a/9L3XEriSm3cU0TGQdZKSqqTBBXpfB1dhe+BlQo+MbBDCsT+2Z/C
iSeRDzoQrc/3mKAjgswu3gxrt3eZYPTE2pKHOqrcnIuy34Z8zUnEAOHG1D+Y
Z5II34T3I7eyH+7vnDsNLRwOCly44P3dLJl9r1ZY6Qjahtm0cvAbDimH4C1i
+TUUIHJkOPugSw/g8c2Np3mkVd5/ooo7aCaYiH78C6Pa0P9GMgftXyfYQBa0
nPKFlpKegRrG7ZLop/JKCT5BL0u6iIA81dlWchMXQK3V/20at6AtMokQuKHR
GINAOF7aSd5CbVhz5tqoApCau+UPmUM1P+nDOLLkApjHqSzyIC0IopS/+HkG
ObnOSAOiU+gCUKAEJ5lWGrGvk0YxzOlRa2J+S9RdZ4r/0nLoS7yLLHDHAEsf
Qz0l653DnhBxKyN9k8dfCCqIgxE9VFSBuHnAj95JJ7pFoppnJ2ngfbhS/FfW
SCgf8/CuCyrjvbVA+x8Ej/vlNSNmyNSRLtCiazmbedOI7x1PCTSxBnqxRrQU
1xbsigE4iDPszZVc5qyAyyxrSdsnjYG8cm100Bv2PqHsYXXyd3uaz+wIXgzu
L5FX1Eft41NTPTmGoGK/fhgpjS8xFRmcJtGtjEyc5pJhsTXkQ23Q6dNdlJlk
nm+0Mqmy/CAtbnWnSgIONCXc01u9p4Ng8yvATLwSeyrihlAH+0O+y7j4Uoye
7LWZaZRWDQjEj/kX84VUhtM13iGOUF13pZn6eZDwlOa9E1IEWfCVn4aXlJg3
gF+NYzYESNOGwghfSmarMYdsBEG5diax7SkVYfzl9D7DD0J9PiDhTllMHIgr
sL4wa9QxIIXFrsEKZluWhoIY0GOdXMw3lmzvYaECP/ltGUu0kh3K+gAdPe0E
ep2Pr37Cv6mz8oWopYriWNbecCX8uItDfoSQLp9wmbSXjx0kVu8QAEpNt7wH
2yP2Z5kFgVw3rLpc5AhjLHb01Rk4VMnhmE7kUoJ6OND124Impun2g4/XO5/M
K9Qaa+qQGmbi0nlM0Q78z6NPgEN3387jtgoR9jTqqLd8M6dBkgVZsnz2Lk7y
TQd5vUKx5ta/9rdiw6s2zYp1GHMCklLcsLEYn/kTINrkuw/xM1xWraO22VXb
cfXeICeldgSpueizLsylst9C9KFoVPPHHrF/jlDj5eOaPMddn7eyHTzRsfxv
imR4QzuEJizi4ZiogiiocsvHklnp0DQI8HX1PHcqeBL6iznDHKkRkZjnrF9Q
h/QndV7Gxqg8CelzBJD7ewzPx/IicmDO/1j0zUKIlaUr5kEGBIRmnCXawntp
ipqM+qVw0FEqUJskMyxt0MhCtCg0iMXjGPbmt+AzXAMTT0ES+l9A1RGQ8Jkt
pInvJqUwffLlhJpCkDGjZ7e4d+IDUa/gsbmKWEobb8pNPSUUN3IBr1G0mpMx
i9P+JBPPbIbLxdYKrEH3hiVMRfMoFK5b/0zepBXMBdWDC7copBJCLURYjkUD
6NPDH+lh3AgG6xCIaenlz6hWyDbeRReZmVnnpMPNCKh+lU0/pLjcPo8/LDWN
TsMpxBoOxh1bx85QUvJleshrNnZiCx2DDfolpwrszcNxPwazQc8SDI10IRKn
O/0wxbt/rH1/BAb59nrzBu5lU+rpCdOduy0WPaVFV08wHRqZ35+/X1SZnfZX
q6OClPmGuaVRDE9CRbdn1/Noyi9qQ4N5/8HzpBEa14QN1vGsH2up8er6jcpG
TfUw4fOtF6rk0IZNGMBv8k9FtM/ltwiZV3lzrBlRkguL3aLBPWIB0/TLAM/S
1NvE6Y8w3+JBTMcNur2wAZKtjSQmto8qWYIxQhcElScdf4Sqn4Q0CZSfD3Y6
Xo9f3XDOUohgB82Dv1HikwsUIj2VgsuAbRSB+xUwUVxEs/JVG5KRny4XEyd8
S9amYUOUmRw0+VYzORVm4MG3RYZfEhScQrnFHc/B+NIvQ+hk5uCX2rqCWcf3
zCDA+vZVzege0Pwxxl6/ATsnV6gK3D4aYxE7uDT1cTxCLZNG392fZx3GYKn1
VkVfQm2cmyj0ksVUxIOti1QT01s0Y3hRhYCQAiUSmmbhsMC3yzgzusO7kvEz
D6pqkSlIVlm+9NODn/l9qVrSNpEWEXnc/DglHjkh2CPY7pNud6iqG09YzURe
mOgzK5uqvRf16NgOA84YKEshjtdGW7WXMo4rcz+Bob/34j6o8QSgwgE3wyQd
pAbeg5QI9KTj9yTgXqk2tCxScgjrgRJgYpJcBcsYZE2VWwSMtlxAuNKWEQKp
tTSNTeRDwpDXWss1XkbfN1cDfu8p7sJIKQltsB6sy2n2xBBFbfyct04h0Mv2
D3Vu5rCasrq/VJvAqEvNTL+eQbIgQI4ohuYHhlA7Y0iS45Ekug23i2JfUTU7
orlCuX1DgCu9i2yIcclkg60wErVB605WNHLVaLA3pGYjCdN4auQGQ0gpm9sZ
ZfU3o7ge78LELeuTwn1KeTFkSurpYOnQgLX2T7qpEv2+MBMOpkLph2RF7YKM
qn3aHSEbIKlvqWle6JkQCXW+rl0hXiIjDJRRhEhsutoXTmzs540nr53ujSG+
3GGAQ7P0iIEOH0xavu5sr2cnrG/q1CxsbO49S6sto860RB8aFhgh4lIY9c7A
+nGz8FmwOBjN9vy474Y8hWxfTPNcUcUmByf2bRkwAGxF61Ai+Q8JJkYo9xAN
hqWUOszhxP94DrpC/NJjyXabc4PnuLMBMf1NFagbEXQo23ffx0tnEFfTx4AY
tOzscEcO+qLtdIYPA9QDgWzNVJRSZFEIn7mNnp9WekM4ovOzlPtLPns6AGED
FGxi7fAScmWsRqDsWJA1YXkL4aVxEvvKa+yqd0co/LNYvMIoeMZOZ0f2ukvU
5wUJLXrsS9JLRSlvAIICMV8QHBdR8S4/SUtoqbRpeL+nhuCX45s8uut/Bchc
YBnYQ8Od2SolijNrlz9PrAwCnaB9feE9KR71ThzgDVjzIbAgRBXWNJKYffRt
DfuQbqtbR13Vt+FB/3mChAGWXWuuQwsEj+r/zbum3o3izbO2NGUgpPq1ocjq
Z9UjQ27IWF5kpmhjIKXxOnwZxdPHgp24CggtCoQgNv+nu5AZ7qg2CBsqqdEm
FjpNISmyJDR6k0zBuIjEo8X81I86dfKDeTu4D0v6c+liAbLF4qvpuiPc+59H
nASBiaIa1RD+RQLBkiCbeDhZDOXdcN0wPhvdQ++QCSEdis7a5qnLHwVEVpGy
rBGtnd4ISLch3VRgL2PIZdozMH/5itOhtKlyAJNndeyxCOQYf4B+CSthwW9W
gDEO3ONjujzdOJftZmbssAwVsU021eHkOxUtRvATZdZaCV5ojqtS072Dx6cp
9Vjtjts/VnRwgN0HnHXhUt9VS+UgznIukAhG+IFPlxe3h2c6k7/h/mphMybN
+QZTvS+raml3faS4XeKIujP8GPfmhP/kOknl/18kurhXpdAEUm+1cm19CpVZ
hFfqv4nqnPYyjD2ulLs+olTPkhymhNgxNpg1fOQRGV5GFww7G4hAnOW8InOb
mWBr1orUCUmIYyiD9OJGWViRGa7GgAtOFSGg7OWu+PFXkdJrUpf3cHkvomdE
P0jQVUmnXlF6vj3TERbDcOqea2puI0M6edhBjRs9GesFdpxh/TnkQnbwkCw5
IjMjMP78BQHyrfZ7N1eUebuhwpD7fv5z87022gma99TVfWz70P+zw7z9Koe7
8knDiOMIJH490UlAorFeJUhTRFZzy0WUCJTJYn0gWy5XlMFsfmVqmglg3/8o
8nEIjWfG06ZqFXxVfSWM7+tZp37pPmP2x5klIrPgU8kSdchIxyYnmoPC2LbI
IThGElo1HvSVGaujUx4Qva0xgyudGf/wzCjEk3eDAjDKMfomL9x8INYhAWm6
yOMAY70b4ToXsQVVd6Z0c5YCiOZ/YY6sSnP4BNHQgtCaaDy5I68me3+UsX8K
XvHzQM1WZFVMs+iDd0cOckHe+mBfIobXYEK9+0vxrJ0dIh4NKsPZC5kknLbS
YmvRdDo2l0uTLrXIrUWbmFDKEhkjwTfkm2qW1eQjHEYHB+9Eruhsi4je02su
RmPmLOjrUGHLOY8td5VQLPgyVEyfWaCTSTkeKFs/C2UJpk+t2vtO4Y6L3N6M
rbWip3vzX/Y3nu3GlcRD8/QEFK2CmB8WvAGjFIQWT7dVnj05KDf/TVgQoZBt
I7FH1H6JY2Iqh2oT+exZTEBlCoVLXSm+xl5xcJ48jfT5ych0vtDjsTwEs8zT
L3dQsblf2YQglvfwLKYlvflCd6K/jRSj+CGJ6z0BZ98Nyb4UUb0YG/d27OWh
ci0W11Zcd1uyQuoc/1/f+Y6GCHEp26I20fkQjUvHr8X7y1NpYM+MlnLcRd6A
35kXXCIYHw1DKclbAh5QEkX/GSvz4vZ9lzAxyyqN+s/Ft95OQm2tw6zD7b9G
z5Mj/F94gHzC3NeaCukm98mJBon7ce1PVR6pvW45cyhqPjCNx9C+lNoJ4+CQ
8SWrMNBgVAB7jdOW+/iWQLvZOfjLmEgaMVyRA0WlixtDmvq5UFL73v7IVFFu
xjS/DA9OKJtc1sDVNfhCD4LhGvuRIaFK6J4j6IB+wsOpPoaQSDWb18lXNHYr
Jrf5H37F4FMn++4VAngTmcUuMEnKDsi8CuBSyeUrm14frj0ZznOSoMLvY9Zx
C3NVMtW8mV5LKeJIbcfiJy8LFwS2yGmrfgtJ1MkDx9DrOV+COwtDNFQcBwGy
EgF3vwnrSN7kuI8SNg1zOp23JvcwsCxka7X5+Mdhgnmlv9rGtcBYEkGr3i6u
XHDsjFShCePrm1xteKaAcHfDH5iwGP0wZa1V0urGZgdnmPH1wu1gLOMZVZcx
YHXBWjjB5aVGeo8EQ9q6fsGFXL/q6UKaEx3i+dcMoZJL9nn7IuSmXDZ6AtgY
4Qi+3Iy5ifzvOAvmSGSI1F+BcyGSJCmkChTJcgg1ydEcdCImzYO98V7xPl3Y
KicPnqUwC+uDvxutDctD5AoWOG0xq/GORoaM7u5Kg35z4RXYzQxNvKDLvVWE
EgetjQsqkB75t2LUKyrlwHhLnYdIRIhKpdaosq53Q3uOdNm+hgo6PVUwKRHm
Ejm0vUCQ1NrHSiF94YLtzRyZ1KBs3idAd7rcf2IHUv8OJZFoTDvbqU2TZufm
k1WHsngaF6HUxR3BW/XdvAZ9T7UzSSeruAoekcZpNIfGjZOiglQzJQZW1iPW
JvrpGPBdMDaW0eqKgRMqcTg25t8TQG2BrP8fl9fbhoAhaIonolICcuWr6/HC
4lWOP13WlhjDzw+GXtdZO3yo7saeSLoyeVfXVO7r4YOGuJIh/hqrjV/x+TOf
M4mcVH4oUOqNQIxQVP3JfoSRESMMjP3zTwggNEaOqpd+GeqMzSYqOUOEUcVf
3gdv8Gmjx8r1+Hvl9V1rPzjZMI6A6elIbZ8ZHx6Lpj322fO+2NaDoX+fdlBw
srRtoRDHOH+KvlInCYkgOiG2/cTopTpdJ55TLkB0kIGmTbsnU4r8DrzACJ8n
o/FEK3WwQ3K8hBhxDIuy3fDlXjxYrUHH1vCS1mLv+n1bAK9DCnWqlAk7cCrQ
TVkTNcVFWGb+h7qI1HPFJPI+DZdzurdTVFkqvxu/f6QRXe/GcReSt5MSlTYC
BU+ppgjSeJinmA5Tle+pb7JKd2FLnom/+8YJb8QSjfsrcBoZKwlYmieRq4sF
+3hpFYzklbOqGg5vslHDvPutCl18CTJ/NW8Ms6mg59SUwr8MwMG5OPpY/7DH
OUgI1NOu7yXP2ODbS3zcHKpZxCRlO9FCN2Z4yWYheauV3BaWTVKWMyfOE5kq
fWz6siNKLuJbNAUBwR5g3JnwZESETC7l4L0e3Sk6ENQspNTuq8mJR59xmd/4
0GRdPkk9imX67dW4DpmTKDC1vUlfaoqesfR8Peik7VnYmLSEOXDnJQFyPdX8
tbP97m2QpI5OOnveNjnKgIuxF5jq2VkijqJmNGKNC93UnstEYMSq4LbzFz4t
EQqsKtvOYFjGuVt1sYFJJsiMIHY1OmJDg32GZbSFvVvZnaRlnE+Lwxumg7rw
JQiZsaSBbT2fFg1iqanGTawkyxGaFqVEDpE22OzQX89Eam3KCrCC88FuAvFp
OlxgARRaEDZcOQI7DuqSShhcQJYO260ZwCWTsQmVndXpC5bnzz6LiTqCdgeO
4daMT+FRxiZSLMJchaOjLGnqptZRt1XLG9lr2rK+QZS6tNQJHuoeCEPnRzYR
nV360/lO8Lwu8dxJYDAXPhXXhIZ7FTT+hyjJhOXRMR5laTdxYsZ3bNLFEDTO
JyttTYEKN/ZeJ3qHmk7pBIiKu9QDFT2qVB2gxHuDGv+GeaSUWSWt5n+pVJ+d
BkPrJ/291tR/5bDHntfMX9UnkypA7/rxPpx/qvrxp45KQ3ee5Db3aM3OrnCK
dd2pt0Vz2Ohi/jO9jf0TiWASgQfWuYuHidJHvPNoGdYsuBMHIuJi3y+ZVn7i
2siPqVjS3hZTdr4KMp+PilUxr1/GZ3o5OHEdUwUakK8j8a2JtPNjJEGpiIdn
qWjZYnTTApeCS2vvU2z0ICR0u6PgyTTb7CVekoSELXSQia87TThMdbXIW+Jo
aoxqF0Qcn4M0yVRh5ZWp+0Q1EJGjerwxzD3aHKHKjgO5VAS7REFGoUvOzHbG
ZlupNejaXOPa03MSFOHJlOc/8O53kiejxDHXy2kD/uKSe+UC7VxhPDlViIbF
xFFQyGjLHlq+PWLED8UKnsgkB7ccCa3qBnagjkxSQJo8kJ1LHw6j5kVNy0nu
GrrKoyFC7D1JV4pTT2fWnMV4vk+Zjp38cV6xCaQODSGyLcdBW2HRmLK/82y3
a3QiVfxs5w4Xo8y4s0jevmhf8p9DHihggczIoSj9zDOrgVpeB+0MNBA8Zz9F
zMy7YwVzB381bkPUSnoeOZVOF1cQ6B3zoffXq0OTFG05LY5ysHTVcZX2SJXx
y5RpZoSdk2eIpwtvGslCBSKsf91HmutqfL5Pw1CaEPIMHwG0r5LxWj/zA2FD
s1qruTdKfeT6YC5cgnQISnXfrY686KNe8H142DmQUQFHwYA2gPodCFVkNwAn
NQ6mBpi+sQQJ+M6lfs6ACtyk6wW/iFeD4ksROqgLeO35QpbXsb0Sxr2Dp5Cu
4vkMbX1v6ZfCBTf0i+XkgDbqIBsFOncs/bBNprb9hiV0TKdxVk1SSt/u01kK
62Jza04134jQkn05RCUscF3j+7unMTb6YLj6xVWGzhbh8ofiXODmXtwdYy7L
eEcSprLgsKTjOrx/7O3uQ6OwZJitugZ1ga5MGJUfA3cglyha3VckCv6PaknC
Hrxxxytm1pHr/zZe/Sx/v/S7YwUIokzhoQ/tDjbbJCcBvmUaDpKeSiZiCd2c
8v1ti4ZgP7wvsqG2YKbZW+lrnIsCvynbt5azhsfnwucGWCF5rDckHpO54EF+
Td/L+m1zxGyRb47FwOWXw4VqwMT01SYdQgYQrl5lvEDhLwr7jSbjUsgq8fSc
PYAODvTuYa1MJRr3tOe1ST7y8Ti20QrNwNaR9sFIxvt3t/xp7Z7mm5GUlcft
QdQk/jOJHEvH0exrznMfLaGAMmZw9SFaBSYJ2DXTkwLLhM2C2z2Jc1v7cX2W
pSUuHYKffBOG/fB2hqNPo/pQzXhTP2rMpaTvyjiBJllgKGAdUuChSB1Tzjcb
Li6amgwn2Bg+sJJmca2e5ZhWwTa3NgscPJW6LLplXvAHTY+HIt8htaD2GfGf
hfLR6YlBFlX8+gZQ4Y4cknKZ3fhdW30nNO2d3kDkiVuXONO5QjL2ScZrYOyk
8Yqmu45FqOwRAZgrqf+suiG2XqWZIwCxgPqosb7tfE0xr0ny5CL3yAgAD4hM
3pBvGXxPZHRyQh8OYx2bMffbkq/KkatmS6mPSi1wfMmCteTMPXaT3hCA2GUk
CnWBUdoMkQVav0pVcC1r/8Embb0ZDk1A6dDXAP9LZow4rmR1vuLZdsr06z2R
O/+Bki+EB123i0rucMMA9wU40A2MTxfR4Al/e944oT5XlHTaE1/5oNjgTT75
SavXBBAzZBowsrQr20tcpfFp1w9RTVV/o6bzUB6zxrOrzOVly1fWQgDVBYwT
1Y0zBeX8JJdNAGBGpot/uxMJsH6K1yrTRXMVDpPPDBBpNqe2pjQ6OBbScFsD
ppDO7negOBWS8KoxWeSCYhKVM+LOuhgY9nK57O403Ohh/NgYP2r/K3cZ0rI5
b7wa8rpYfCPKGYqjotu0BAUxDfCjQi3G2G5F1PYD8XlNTBr9Icq001dnJEOQ
idoV1N2eYD3Ap5sme4eMqsWLhdxuQMs+XA5cuGNuCJ6KE9EK18BAhnB/xn0z
nABd7ctK/PQXC54dzeL78xtKcBF2dxeJyo9MCpiyQE3DrD3Eru3eX8xRGtyh
FpDGM/ePK68bPVN2KYMPLsa6NHsw9u4KxEN56OrGAXBvL2lfAW8EtHJ7FfHe
yRc8pNDSfIsGZmlFIyr/76wX5pzsT2Y5R+dQf9t3M/ktxE1OqNnbvx9Tlpfl
mOPoBVEn0cEN+t6MSYEhlRPqtE+nQfYUSa0Aq0B2PdDfHmc6HzpSUzahK2df
d1fk5vYAOEUu0PuIuqOBNPsQ+mrbIDGAOuRJqb+uXP539QIBRcSnqm4no9T1
MnOLpO+z5xaAVrHmjwlRYWuj5afnGbapeD/QYoNAnW1R3xVdoIyo/+clrWGW
4mWnn+tA38sv5NeWngALnnyNPKcYtV8Ql7k9sy7TQchiBEDOzU2oQVbAIgME
NSJ+mVyqml2v4A7zxJOXLd3Y/ARY14Fj1+AY0gyrVDL0OUyPb5yCCXIDT2i+
KM5laPLvVgTAOChNiSdmKCDqsTWWauykcfOGdVjaxTkYx3T++ZwM70yw4cRS
7jQfY5iwTO2t/U+tfYv43X3tybEI+FdSKkv8x2doofLuw3oplblYSqLoqFoy
svz5lYy3jIlqRFUGeZjzSqQ0cbDjvdcap+KKvxnftYLoprQ3AhLuSwikh0Uv
Xeuk6fYkR0vrY5ScRq3dfmaE1sTJVhsXc+f55lgayiajZ2gr1fZY+Jk4bqBB
IIBq1IhwE5TSAGzswgBYcxUpyIXgqmIgol60VoEnajWuBcQYzc9DTeNb2Aoh
EPqIMdW6u12YxKzym1KVWPCFWqZhCQtijWYw6oXpH7JrGIY7a8crGFlu8Wpk
5nVpl1BVtVlDKlJOeqHT0O+24ZlsEpwMIRwYfhdxDRvePHOrhntOqaMrDQPz
uz/zCjeqqFfB2sBjK/YrU5CzGIcUM0nkP4aMdkHs9Q9lT96fPXyA6WUcdR6u
v0epw2LU6XaPs44jC4/nAgmrBlCFPEIoNI1V3Rer/gc5ho1Z9gu68oQJ0q0R
wanC9qWYn29wp/5B5aJF9yLSX7WvHHCABJFoR1srah2bHx4rFRQdPfXIUmv9
mUtZxGzPJ0R/XS/FNuzdGSn9lRB6uZkCYtr7CXlM1SUIoGPnLz1fM4dBRUBg
KZbEpa7uEYvltYEFIgODLOohobwExxE6XAd09CVV+9L5WnDK9abs/TNE/CjH
iCCTrZL/bHOzMc35SOeOJnf8PAojMKsiV/qY/xS/5/dsXEsmodu+e6xWgW6z
8gwFVI0SlpJSc6gnfqje6MO/lZFfdsCSu7oBqV9UgRBsOkJbtW8gc+CdXrsZ
PKH8lb8/myxxfYG0reQX2++rXd+4t8K3D39JtFRjC14vWcfgvePOu7Ugneb9
1ezrUt/TP6NMJ2tpPr0cS/EhptI2ne0u3HCq0DaXVh1FmCXNz6fpZw18j/k9
TmNMRi7wPfkmZEV0UmUI53BLhpR9EWUbwZeqFjegzsD7g6Ajs65For3PKzwt
6hSk/+8yuF97fMvXgrX0ATFSJ9YhNypY7OnHACtu6UqvKuyuM2rScx07+K+Y
3NWghVvlFdhdlYIFLwdmM7kY4NKYhHVHOuHwXi+SZ8vbV0SIBIWlPHrV3Ogj
hDdM/1too9uuZklHthmka+Z3c1ZquKeAyfWiP/iHQcb8DJ3A2vI5AdTJMeUw
uq+3YsQc01Xko15+WKYrfY0kI1XaGGC+BTcsorH5mH8r6cfJzpSy79fFPUzc
5cwMC16kZsH2T48p556yArhHdoIHJZ79AOHqyUhf4qURgCsfrV9RqQJ9nSTY
C+mDfvL+esUDKxeAtnyficagSPFvkZ1LPU5JohU7h4A9s+LagzfSGJmSHCen
zMUMIhdf1vm0EVwBWhWkiMZjZhzbvI44JER0PSHN2N/f9LX80siPaIYbPaSy
rZz1Ge8r9KKkOJGjyXnUfrTTF4Ac36WTufU/OJE1kh6y1/Ijw5Pkb3iPQiRX
Ew6OZP8+IzR+DIio8m4YG2oMVWhiBaN6BJK8Xtr+keOHfRzC7hYHaAfXLpIK
VW4bM+WxQVvkC7OS7S1J4x6EK+NrTKu36DgIe7OQtTizH+XtVzsXCIZPzKim
Y0VIeMiCVuQVe/sx4Zs8oSh0f5a4fvYNvt6xWTKC7nacGvdHZqqoqZm5Fqrl
+iJzDlJ7YEBe6B/uIXgUFimhsY1DQaHq/XUeQPzgfrjgcktmR2S28YzY4uMz
TR5x93GbL0SykBLD+RgeVE0t6g530IEVWDalXtppx7w5kdAjzg8EYH/Dc2lj
lJ36KCVsBEqiB2pTEQMDkyUjIUORCd7ldyEL0U+1t8UvSB1ZZotVjMkNUZCn
2LKBT2QFCSdk7xoYLRQ1Ub4dN70elVV/fili2OqXgcDkehFNPvWJ24iAq5Ds
VPEL71zNW0x8dL6h5zNC0OQRxBxOQQJJASFHqnJeYdNbzidcYlH9rDYtkH1S
FbcmwvBZD1VfDYkazWHW435LkaSflJpIY3cPEftHPH6Y0mU0bOrtXmXBkb0S
1cJQV/e3zAgkd1nTgS3FdKivCk9Mug+SCfh+oRK5egrLcb6TL/hf74N2HCLP
k6dGbF1+7o5cBAxVtG6/BzCiihSxo/NeVpYDSe470BmncrmVr9rqlW3t1E3Z
KoO6bOhxcojRdQXdp/mAC80X+iOWd9S1omHiKOQ6ccenJEnyTmv+YkI/AQMs
m+Hn9S6E6e+wy+Od7vBPOXkJKTfKHl+pAiGCD0pxY7kDD97MUTRVlBrxHEVk
mDAG6gknLUhGrCmobcTB2DdyX8oW+SNbRDm4GPD/pNFr0bv0FmTPBwqpRttE
yBSqcLkg91Zqx2EFIRtpNZinbwzbqB7XPy03369EAkUxkIF0f22eZ+FDLLnN
lGz5z2iUcyMDDbDTrnEBDgtimln50OXIWyu3gX1OKZCPV06BzcBALwc0mOVI
XhEm9nqCmRJgMv8pOFSC/h78+0+gUaA9wv4aB3nsGclIlCAeRmw02Qeba7Gc
3N66s64gMn3gbeCMih1Mz1ZxNa8Xxhvi/KFFNDhhx8TjFuNab+ODgrvPu2sV
SlxJZYjEN4lw44GPPpFgeX4MIckDLd879c8VlJUi/4kfRlebaPB63MfgOy7z
iiLOOt81Qz7hG9eICx4Ga2wMUWBQMKvT93xSBBoiEZDH9bQV26b5hADucHP0
taavlSd2fPcHD9KsqhMTvDGocyQPKGjNTNDdqdDXzTAO3TyvWl34IkviHfRL
BjxKW0ilsvHju8GrhnYK8ya9lK2Vk2OH3+QZyA7vPTtPb3VlvtM/LnQR+luc
QL/N/lv6AbCOj44ovOhS2uubXO3xHqiQvLLRMC9tWZVl2o56QZO5W0e+ootJ
S8SK9tAWCKq1AT09ZdjndWLZrEvOFIaD/0xYaphQMfyuV6Y0E4oq+927VWXF
8ad3eQ4Vi46ZgkdkWbENngxLIU1hJGW+48OKixwWqYCogAy2QhwjQLx8e6r+
5mOo5UarJ8CKro60ba0DZukFuykBa0t/5rjkAXZLtQiy0sOWz2dLg2jKd7mD
u6Eow2SRB95wkwRhKE7MzW9nJ9uIEdqJQQPYf8a2ajOssqu9v+jOH3gcUhT0
XsqFt6iFGfFLlkFgkB3qdPlmZO5mZS3PgkPm72/hGQxoB4WeKYt17QMojhDA
y70ih0R9BECmVFZLjk+v3QdhQizIY5FtCx3esDUVft+XX9yYPZR9nLKF3f4e
IOALA+AubY1dyQZxaJzZZ36B/lXkKmVdP3Zd7OTR5UGaR6sBJEVflyTMut8Z
xEnZ11nTePGbTW7ViDKUtqRJN+QpY49fIP4dDeyY7b8O24PfK/G3WfxHWFmy
5tkEWdPeBH8R1G839R9IHrmHzJwvLrVS7abyFxaBDKwo+vjrEFf0odbhu5os
lVOeYY3IG5P4O6omyxnKpOHy33J/sYTw6PF4jmcUc0YKVX69l8ahrSXkDN+B
l01qVBAheRRrGosRukwAcjZVGElT68+AXYSfxD5cIVGcqXWtTjax+kcGarBl
rtqWfVbBA9JtCJnYbfq0mSGTqesfnkBpfVTNdvGR/D2vjKY6J9aalzO26A4t
Od8ohoaOsT+EvNIV4r46R3XUrE8vWM1Z2fyxhK6ghkGscJ5mbvzvVrzC9V9e
BKrDiTvX1B09T/8U9z4r7SASy7OUDMfShVh3BD5JsfxASGit6fwxtQsQdcrM
15Q664Mh8a7OIoeRcgW9aUWSHz0sqhAjtCsMphsSpjBdKo2NBKL1VpNLlgBe
rycwMIu0UwVFE0KaxzvJ8GCU3pmNtz5PdPlF8yOnvy7weXh08LnZlEUQF3OD
voUlVJYXFkRODjm4e/D3IZv3pjT7dl09ulozzawe8IVMeHWaEx+Jc/03rv0s
B+SJDA8RSeTloqs2ISUOcvZGbv5Xuvryq3qSSQCU0/F4ssRcgEyv/HYmLDnk
9pr93S5TrtIo4LOJR8OW2rKsqWK3aUVGT+bIN26/TLsXdQy9dUFAPY7NYyDm
1I7S3eT6GbHHiEhQtSZWUOK6T70X5wJ7j8dkjHrqdRQU/6V4jOmffCd7vua+
a3vjoNZiToFYapNigztVVsPecubnWrMV2QZ381MCegt3RNxgyqvWSrtdJ1li
SbUuzvGZ5aq1YJSK4f6hwlf043cKwv8/r7Z3mhk0ElHDgPVo6BwLe8LV51jr
T5roR4EVs6RgdQHmHxvriCDv8WKynHIH86Mcn+/ifEvG9lp9ydYsI0UWlgD3
B4aZ+t/3YZ8QiQIm17A/OGNeNVb3EvV6izz1Jj9hiwcqdnKuyP6R5C+rbcq4
Knw5c9DT6QvBZlfanITqdnYn/sziPUQSod4nHfIyt2340a53Vz1wLFEa8GX1
XXfsAA4mWDCPX4gfpW/Z+rzWMHfE+0/UQ7q+UfOctK9G8NsaaiMDI8+Pn0ky
QKlJX98+5zD/mxj5lUkJARYG9T30q9MR8iX1IOqPWhHZHdCUZwQgeu29hmu9
9ZTseKItrEYW1qwB9QIWvhw+kTKtKchjJWxXV0Wm3bb2v11lVuDFcBH0XZ6H
o12ac9wsSFJePYEzPGRbHDtgc6rAXtAyYPNgGxfMaON1rR3VscuDPricx1Vy
0NVHgwr9Xp1I8l5rJefOe3ZyP1pDv+Vm40DwshQVDbXvcTgW4wHQalxLQhig
qPk9h5U/znNfWcZrMEF2Q4cqmmyZQfwv/NGUtOkN3aKXohjod0FuL9ElEu86
emr8MQFmrm/KTTCwfaXVa2kuVVwzu2WT5DPdyFwrI83CBOkZH+vfAS2RP4/w
xe78ehdiNQkzr5G2/qBUImymd69GeswIjeSYQ2+p6P+t+nJqdKMX+WAvK8xE
U6+0cO6D0XZUzfJyvFzTVaCaG0TCOsndJ4paE0+E00JSLriq5YsbZGgXVd/U
bzZ4KK2PBWAAQRcyUB1lXvjVWHSv/j+pkvM7OJqRwbal6RKwkDQqGtrfaE/g
eyzfwZ/KzPADtmFX9dpPecwY/5pELQTTCCrTOxs0usMDaeqdJ9frOwipET7J
vXLqq98KsG5zC70SDJZLHl/ggQ/EoxpN8xrkMXiaYFvUzkwCNl7dTaBdBxFs
degvB5yeaN6562nMrMkhhl5hQ5JyAQ6zTRH1Zoonf5NXg6QWuHKHkSS4hTKM
XyqQCiY+07EsOXAsJcUbTnTbAKBV9MdY0pfI7NHk4wkEKwCMuh2xXlZ9xpZy
xGFIB7NYCa/06Kt5JfG/STJzOjGxOp/w9v2odRVF1rwrlTLDo/BMEjJqLmEf
5sSl0G18EadtZHH2Xvn2zPO3i03TX5oEn2I6JdLxvl4wmLx00kyjjJ2f2FV0
Lr+Zi2AHlDPZP1XI39erHa6BSZIZ7fTUTrk8gKRMezSXV7mxT3ML/bfjVZjm
ltF2XGJCj/ByiHgXV1zjtHGDOPVjwkpnOuvKd7IzrlV+w2PoVwsfElkBdO8T
yKKJ4PpRtWXQ1wnCFi9MtCvAr/KDQSrt+wk1Ssi7AiqP9URUnIPQgbCBPB4z
EUwm7eMgGOwJJL5mPToqyusVK2RHGkR0q1zrsTuQAfbWdTY/j4k8jdogvNMt
WmVJCJBgq0F4FXVPiv3AbXfkdPvsl9XTUGt/O/Vtip+/bvcwkNBRIV4VMnW6
5X7YL4/rQRxCNrzcw+Htk/lQ+q1UStuqDa5JMNdHvZbci41IDS7g9cTr97dV
E7I90qdyZ1L9AXM4oKgGQvboqU3NC0VHDCB8vGCzL9yCOpOeNlP6hpmic4/y
JtiuMzjnJ30dksdaprESFU/7gHwwuMiUbbowVfH6D04m2KeLlsKHJCgD93nl
nOo8HgAURb4b1PUNBtwtQpT71+nPzl2vHsQgBDDraMQu/nxsNWX2UcPxDe4W
rzb1HjLcb67nJ8ujlMnwPYknD7L7DYcwJVmmks40V6n5OOk+OBEG/uFP7qrj
w1Ds/1S7uJpN+3QynsWdWAIBsv1KNllrovnjPDHBwoy2tbhckRl7FAJmIUce
3TjByWXG08ay+0ntKIKbTfxpiaIWKflYA6WFJWyYaQ+Ap4GvzuZte8LBxNKk
1m1KaF78E5bzfb0gzbpunNaWiXlGCSlagh7lSP9Ybd2qLk3nviPZRxL8RLjt
3KFJRBvQRZ4zLeqoyeQ8apohqHvao0h2ruLgSl6VYpIn968qVekdrbo/hSVs
xrO2BZEjzPVH/lx0dZJqcbkFH2Gd2L22ZTFB63tMCXZc6HyxVED934qxl2I8
C+5C9WFU/ENpodgELjYidBuypnJwb/6QLR1W2f9hxlgIoiFlkKBb1taNlH6X
R9C15GPgMh3Cz6GTGngXj/JieVhIsAnhJj0/j1VTElnuhQtOSoGE+CT/KVAH
wh6+pehyXs4oWFx7ZPOVwYuu18bagiu++JFKhNJE/UK+kUl5u0GXwPGZotgf
KdQAfUw7rU0KkgcBVzJPNcIoO+RdsMIxXHXsJNs//0Kr1sVayx3n/BwDa8mx
pRCmWij+OBvc3EfljxXEEEU2WDpQJqOfexpIgnX2FYK9mTTRYEAwsbAWXAvA
Ghgzlm2y7HcKUoClDbBnz4AOqJwucJOWztIe+3J+43kFD4AyUiLNr6Qhfxqg
KGNX48ADJs7DMrkYP/5EKjhctRTiaMvgUb7a4XiXN+WtMj0Ehi2XmntbZvMi
QmlJBPE/0oy3Scz7paA+DS0cyORE6ZkhcnQRpg32j2Y67+E9xFqRRCQyvqoF
u5NfRFtO4Qxp6NtjeOuRmwi+QuIT4J9UtT92jtatieFThB32f0NPxmckNdSE
ma+x5VBTxIgqAtzOzM97U/TulN+2Igd+K6hbJYRWCbQPikrMRJqU8WxpshyO
59i72ni2d34z7uq9lwvKwXGYmwTC08Po8ZuFn8da12PiRZ8u/Wkg7oaQsDDi
kQ1v5jK4t7Qy88xs0pSIbmYZGOeMb3EzYxeUr9vP/rldgGLgSp7zRAvPlgtQ
WWsee75OiivNJhgJc432PkA3BCB6gAJl3KiDy8sHeGhyLaarP077PmeDz/0J
JDbEhuOS1ZQ4Wlx2769pP7Tp1Cy/FbRgSmhnvrUwmflRBeMqNJm4nYAeeBMB
CFOoOGXI8MfR5Y+xxDFSPPFh5CNfXa4jmWZLwMHeFEGVt8USjFBR+u5plSUX
gK9DLi7bqVilyHad1h/xXMUSxT60707aO43uoChK/6Np3Gv4QKc/aPJkGnmZ
iX9jncU11hCXfic33Vd76ow5tuULzt+QjTjkqbh+FlZXar3pZ72a2pbREHdS
GSfPmHTjtxU4dH/1N8SZgEQKNf2MnBRz4Z6apCpbzIYS4dqxbrxv+zzhS9ct
dAcwuanoMRSk8dmYUeOkqh+ZnYDKZLq/6XOzBHCeqeQvIcOA7RYeOB7xz25Y
uN/KXUAHGB/eYeczGp3pn5qi0TO+v9E0foCmwD4IFshBjA6L6X0n85XK/qeq
dYT1C6DKQFhf7b2JFH/XUEWj4DHGO58jAzp4plKb/eizzQykWlqOMBqjlyO+
KkYrq428W/KjQubvf8hu7NLKKFiKL6KgvpdgHjTEkViTnTdzBBMD1isEwB6W
h5ZsoY2I2/G+gCjyU8H0c9J1WA3cQ6387HnrPGusy8dsPYMgj7YmiL087L86
MBtoe6zi1pzDqS5QuAqN+uQS9McDNPFpose7t/T2yQwwq1JddOx04xsxzEec
LCjbXbyi1Do4VPBcrOkrluZYF6or7i2iCr9xKslZ7FSkAXzSHMykLdiQNhEz
irneYgY/z6H9ZpastTdztQw2v6Fy4D7wpa/dAk2Q1ICACJAu6HVuY5ba4s7S
nCMlplkCKeIgRrBNca7xIy6LMrlt8Hnw6QQA55FmZNJk7xxL85gxSCO4RUJ9
TERd/hUZQk8zZM/897JXFo6NyjlWhrtKeQnMgW/Ep974AkWgj6Ugdx7lFxCP
jaPfBFkbxZ/SIr8zxirl6kjABk33zL/DSmYj5Qozkq0cAB+5kwotAKPGzHLN
QuArt/j/Aa73XwOvdC8iAuwpK6brnM8uoY6AuWWaZLfpb2utK8loZi2Vd4ED
b+vfM5S2WnilVvTSBxeWJRPfnwmEwvmzinCKOREhuofTbc2DJmLu8/DpIkdT
iRO8++veRyhknt4s3ITCG0CJNUyK8IRaNq2OK0d4cT9lQqcFLHA/jnykvPGf
1KPHC4Zz5C/nhHVu2Kfyk7Dtv3lNrC1P3z+3TGvmNmEovgF6vXWmCk81nlFL
JOdrfknHi/tEtgBaIm4ZqWhC2/Zk9h8JDxBjAjrqMzDznV5tI2hlqUJsbf5Z
/vkTtw6AbiCkYEoK2w/OD2ZBKchpAtOrqSyrHEowc2ilf8COfBDwveLNdHE+
I4SBj/OzjS7mYjguWG5XiOiPsGKWWj2bNhmCwfXlzcC6MfASc1mQ8G7EDhEN
YBRS9KZyI7tYtm8y6r6raWHasl9ozQ37jZX3z2VoOWeJJJqmr8ChzgBejf8C
1ELWq7+ImwC64/r5U1k+5GpbAuwkzgsIqTsBmO719O1Azmdnjpuqg0okYZ8n
R4pp7nIXayECQSZRVKBE6yk9ITlHItSXfoGRSDvegXfLTBqmKjHEicEIQ6UV
HfxJGeaipBSNuA+zU0q77yZa7eyleRbLZfjSb7T9RIEOpOTrlVe4y0GwajOb
Zl/WeXErsLoKx5tB6eRQv7Gr1jx2suNgTf5g6AiVL1f9tQFGEtXsB0ia3eet
d1hGrm1PCT855F7j0i/j9qt2PTwwvMrWsrsL6u+BKLsvB397T2lXuKTMFTtC
nSFCoMQb9qoJ8gONaSYSBkMmctfxXFICcLqTn1Hh7MXS9cjo/PhsXR2m2z9d
y5EH1rd/CTZzKThfodNXLP1yLzuC/EPGFBss6DhZoDV6SjPaSBVM32H4HmVa
gLSvVJkg+h/wFJxyzp53e+ouy5w2+hgAPjb3mxlHo5raeQYsErk7yYkP7H0z
TwwDjzLTpcoB9s1MCfiFJr3+0klFFFEqeaqezDTD1uIWgfxjle3+r/2ZdNmk
Q8JABEuX4z1ZdbPlB2r17XQ9KGMjScVONPa1P2jCOYkFz6xYewFt6tH2ne6Z
YMVYm+ch2Xrs5o/kokUpUGTjtveeXYyvIuD4HUtRhBVLHjtskE0LKpgmSEQg
ag1t4zpOIez0tByBlNfWKq9pTreDuuD35xa7+sufJZmHkPL9Ng8ROdBAJ7tl
o7PL1KYAcxMOhCQOyAnA2AiHsRAig0ypP/g+NaTlgBJc1170MZgrca4W4PiL
ac34AWXOBOdjEGctM32u78VSbAsTHymzz7DDskUO70tvuHqWrFnG0EVVFqwR
EOvDzOprPMZ4hNzjEC67dhrcf3bd1bU4SJrbTiCmAIaZnRApVnRIl4zvMp5B
E+NLBnmk2afIQEGBAi3xkmQU7eua39wH9it93mym5x1r5VN2sG50cTdMACcT
mGaCmhZflFpOds2m6VJK8EvmvU222EsFgHoPY68VhXQzjQYEpQzXcxolikyW
44mFnfNlXju18YWkdGmcEZaBkrl3ZFYt81JIFBiGh4tcVIzBkAnz3nsHG5VE
pnX/ElZvlM9HudlMWYjdkDZvzZ+3S/xgT73d2GEsGmtTV/HDdTwC6hsIx4kR
tb1+19X9zSy66ezmwiZ2pcyniSpNGkjOGR+8mo7wZhOlPHlS2wGCJIbKrjoW
kDPb/mGMRXcMeNpDJgMYUy08gT70XFgSP5I0wGxpar4uccTFAkPMejEgeaeK
YVQOxCgBvKcZO8oc6ACE3Lhc8HpSzk+VfAnm6JbnESl4jx5vwduyR+LGyRKR
7kRo/utfERxS2i16d+fw6ZRB4CjJD1W2lpqiZH0ghN195FPp3OLIzftEBkoB
rBQ7bM42QWPsQHwntCLd+THJ38VOx74gfcYMi7j7vGjQT0STB56RIdtDRL0v
vOPZJBRk6kZZSRC1SpkoswHUWDRXRh57oG2sgL8gPqTeCatVtmtS0fDy7aD6
NRreJ/NfJWPZKbmNlMq9ZhI7xxgZLyQhkhHpoFO7wy2/D8JWBuhHOvy6Sem8
VvXYHcytOcXmEfJyvGklt7prvufiUXtVGdagSIIsa8ZgY10lbsDqy+xsvBYX
5b1V1sZKgp0qdkdh6jOGz8KwjJ85Nk+C6aY+FbW8SJjcAo+UY8wcFDq/bVqd
oFpAeLnHOQsPN/xiR67Qw4iOrJ1OmLMoyn05/PcNc9HizX7Y5/Fo1iUSWgIw
RkLTyJ2SIUMe+XS4ez7Yam9dZMrI5VzCJpeMcleNA8LOlgX/aIeshSCJLLFd
FdmdLhvUobe7O6RcdGouJgXJWKm5OSA718bWFosLIw8pU1leMtkqYUB/uWGq
h5eM1S6kmcjFWLt0mMgf/5E4I8Ill46Fa3OcsBzVwuA1SFTjEl4Di8/Nexak
sOWgojra7Uz9RgJzFEk6ZVobR3ax82BwIuFXKGQ3XAFyyg1ivRLoVZubr3aT
u/YUwD105RXT2KZeg737FrG+zRXshgyQwe79QnK36j+QTpuqGw+s7KGpV51n
E3p/1eGZgO7kVu0OoQgj1Fu6rZnpIpH+GmLtDc3eKmf6fbnZey+j56KEGMH3
LcLelDNxkK1eiLs85+ED7iTJXJ988Qjc/kkpnLwXFeg395AtWr8dbfKCYDFm
BleZKAh0QHCKrHjMhDZLYzWBD9qnDMoPQMXg62k2+XknCDCw/Kdxn2oeWiOy
V36DlAt+gtjd8n7gE0dHsteUtT9k9XVevOj3pYlpmQciVmx/PyuRI0nHTEVJ
72BXteKHjg9aikx5j6qqaqK1SCQSlDEA8R65ZsDVwxdlnK5jDbgWafOx1yzD
jz8R+4hcayHyvSH7TYlqXHtY0iOQixB/2mYLXUmplHnJIwKCfr8HWKneymwz
eLJrSPjWOcDgMY3TZVO5DBSspE4zjVJj4KzFFV/ItC4AVvGmweNEKwyEKTvq
7hWFvuzMAlSh136hMltTGia370th6jfoVsX0MyMKLHBG0ehdE0oD6VOd1HKx
xbjP9Bs3vJP8HDo8ELjSDrkSOkpiX2ckysQrhGsAc+aYZQNxYva+uMkQTYRp
by9tkhJlQsfGqZtTj0u7yaFjexLAoyyPhH/EWLMKfeBcU/pg2lsIhZp2J1oL
IGBknCIBBd/pESKaS5Ih/6EtU9jXVJ09ndDWyOLKOH0Mzsv1vIpn83OGBEfN
x/pLJyUVkt3P+FimaLpF5e0fn8eAZS8JtcdZzXyxr9AUmpm0JhNw4AdBYCrC
ZqTMn6OGuvw2PyhdutxlbRLe5Gu0yoKdEkJZGwNq5taN50zVdFnhppfcnNwO
MFC0HcJx38+Blxf1bhaj4oV9w2rqoKFPWyRwCEhO2trz8MQDNYFP+5xHDo28
oo0uNXypZRFl796LRlDapdUprzMNfav5nJGgnl7WWNAvrF2aX7Ihx2E236Ji
ZEYmwgt/0D9zi8ar+sp/c4urYmDVGpUsF+EgCpSoHmiiQ1f3a+07zt2WZ3eB
ud9I1bArmrXv0IRs0iOP1iZda0BbD9PA0RQoSAlZRf1r8y9m2WGpWx/N8Y7c
WCR+dIRKTrF7HmyZm9Jnl7+2RrG9L6+Px0OquYcKG6BEehuZsoVr450ucoCw
op9La78nygPiADXmoXgdhpTYI0V+HrpGLOMyGcO5eY6wjCJfPH4PHAwRY4hy
orrV9AEzQFgMOY9RIBVEcE3Ne3g6MboJOBkWOxlaDwcY+eCb/Ti59MyqL/Pn
rJr9fkQ+24EDgTxfiKWgMwXZxDKk3ogqeUP9Dik/ZzDWclTLeCCdovhxWL7n
LxSzzhYGOiuRbWBJpTSfE1oPovuq3DLyt2ed7ZxeR+8z1YkUdpI/dV+rSZDm
ix83LYV7aPIvSljtku4SL7oj0xuvgUv7a4V3Vifn8aNddvgk+2wJeRE4MaT1
Ra7Z63IGsT30kTWq39PBFHIwXY5Dx4/Aj7k8xJIPUKY8IIw/zF1bju/487aV
MGk9NuYC2SE3fJTCcoHQLFw4/K5QrOuwRlVrCjlN1WNCsfbZaiQahZQsr9eP
WtmM/Jd8S6p/DhngED7kRXFwBOgbNP+HpVbzUXQNGnyglz4sP3Vhf6gUNy5o
d+vJZdjJZDM2dfrYdZayF8QaHBBiGZnEHAzbtTc+DiCsrK3Er5AV/cnt6Rp8
OiPaxouap5HReg6I+dsE1+4w54YQyUnRTOisiFYfiPUH3sYEPh9RTAQy6dyb
opEqLRl3Qa0nlVRiiTiCbsj9HcEJ2yv6FMigwRMgdmOSHLx/YLE3LcDJS2Ln
jt+kLsWWJF8sIkg1Due9Aw4q6vt8TKmvLrKTYKzXbgVv8liVHpYd6or9/YS3
9yZv5SKozjgmZmJlawm2Jn0VQ6KZwQedeqz9acGdig3KHnKEnl0c+65VZ0PN
WvG2+Z6pH6Swb+vmtFVZv+Rj2d8Wry/9ncvlf2X2QHwRB6+VMQUlCu15nh3K
ti0b3vFkeiw1lH94SeC6S8QYlfeyHGhqULH2G+lCkCprftyWvpKq0bes1kSM
F5y1bom8MHVDPnLvMgL7r5qmtoonk2zG7NMOwrahVfMKEaZ6zeljSTlbymUD
lOTGAexb8K2EFqWhCh90tmG5jndXbkMLVPq8TI1727A/w1gRCVVbEE2ZH4GH
aAmJNuMz0ug7EG3oDoCY3hzDJdxCTir8tkRys8LJMXxBZoWRbZLt/Lx++D+P
6Vo8OMkLZsMD4zCsFtXjjPZW1HdmJGRYzGrCOUf5tNS6BtOmSueyiD+kUFyR
0mZGbW7D/Yu1F1leAJ+twDlgpPi3kjt90LsEVWTjWqptaRtDllqib/lpQLYO
DGVVng3RIz5ijCO/RZE2EtaKCui89ya2BcKu8kmeU5lZDmGyNWYOgUt3HjRb
Qd1vM5sF6ay+pOP88p7zwT3xgIhgb9YyLTe14epZHh4oxsM0cJu50AFjqfL+
7el77JXC6ir4Znqatzjuik1X/VTl72UCsG/P1ju+7SSopeV5Hulv0ALJN+j3
6JT16FYu0voQbS4Hn3CKlL7VV2bS1go7hCYpZKh7f0v/KU2S7FAT3fdrL3G6
R+MZ8FodR9lG5HuquIgE0+xYeFpEHqcbCutRf/v2AqTlEAK28+SFcxQ0R/cU
GsADkMJCLU+ncuBlvac1/2ecIY693rApEv5q9X/pWt9ab9JJAReN1nHN2NZq
YxpnuqDOEgahCE3qBWdxRqjGm0EOrFLNJMjizWbqZLSjSA0uddS4XHGxPYjo
l9AsfnHOAhZgsSXU7sm1E/LMa6BJEuaAzxGlIHnkTT87alNR27WNnmnelJI8
UQdacp1atzoNT9ej0Cuwc+doQJcO8X9FxRJHGjNxADLu5vy48u742liiJczg
1uYjbI5r70a5iF2D9DdpC0sgl5q30VjFC8nwXFN0VoVipF7e3sxrMl17I/S+
5nbkQdZ1xDSCR+7Wuh2/4Jt97BUAmmbAvTNgxkzt4NfjhZk4nvVYxr9bFL0u
cE/xGb/tclxr8pqFL9Kn1otDN3CAlPghbl9mKsM9gnXWb3O+CHwbMqQ/Nvuf
VEZc3gHoRCR8B6KwStg6xaoHGe/08lkO3sOo1GqFGsxs5XQJe6j1iUTr0zqD
VDa4FKsaMa4sjneHFbZRsRz4jdpSeUTNu5zr5+T/n9LM2hE0e6EIwvAtFrxY
Ym7fwwztClq59MLo2CsnLPAYmFQrnLK9Ulq7j/DU3W3XIgTzHeB9hS/9T6zO
19XUJq00ejzM1AqOUEuUf2yXA0WNoMC5bc+OANPc5PQEuuFeM7xWE03GSsdC
t1rhaLPgMqLmWFnERqyj0MMuCmokce2ne7LorzEu/x3KqLHu9sYzgsG2pdx7
DaEs2QKsS7MRZ21YimB7Lhci+kA8C26EggnKkEZ3TAjVHt+bbAhU59GR5IZz
dmzq9JjnJJE7Ydyqg65x2FGX68Jh8gfOoGIz2ztjs/j1xV3zdvEsSc9fvChc
EGgPfBOyo/GEImiyvjFwK9LbW7SB58ntJHGmfOipGYaCFf3mt8lrTgcNegen
WH/rgUpnAAjAA/DYEmmsoQnZxz2Zyzd8U/QsCn2hancM4Hpj3YYC+BynMNxC
QeFg00mAOTsewb7H69a6tQwguTJm9jZejdj9W6901UPXQ/qU/JoLDmoRX07n
u2cVJcVfDDbRgwpzmGyRaRGNTpBmLIPZp9Rg4KmoxYGkAPogxGLQ/1Mgs/Lf
EtB8gCU7AVfl9QR9OiOQaYO7XCi7rfWK4wAzd+wiQfuyooqEyMdN8yqpUP9c
GnLFNWU+WEYI6oTbnL1+sfzjAT3PJw0bKqVGATT3vSFXMg9SLiPLT32cC6DI
QhIFpZNsHIs7edHW1jnWJT+VEPucyCvWlvOy1URZUlPHYfl9dWVm/yEo0R61
S7Ty5niIyekArg78XNMUKqD4CCIq+YDjqtsEGtVzA8ngpU+n5fKR9Z56rMzD
9xU+vAqU1e7f+olTr5ermoU81QnCC0i/wP1tthQ3HeB9QsnwUV1p2L641scw
qWE2EeWesFOrvZgF5IxOh9NDHRSZHC4WnBplQBDyDBHOERn5jE7r4qs5hauI
OX7IC1FpdAQoCBVF+bwHfASn+yd0mTiVr3wSM0NsLeZJVbvw42bh1MIn4aM4
SkqQdV4iupjdRs9IETv18w7M82pPRr6h0wT6F0abNQeyG3NNUhBf4xbHPA8o
kX3PyymQKYdR3atoKBt6pyzrxvXVYaITPaJwOBizEdcnRhymOQk5JKGNvPfx
dtwaa4ZF83hg7+i82D7urI0YzSYx/7+N6c4V+i6jfMXDPpMRzRfdop0UWBsA
A70rOS2Px1+BLtiDvrsCsSZNPe1E6rhoYbC1UkQyPHD/IOu5D2ZbD4ogHtzp
412myMoEhdF7yv1PLDIhbD7BMupXEF6flUxHhddneBbm50fhMi7LY5aWaVwl
vh1JUpraDqixqZmXG0b9IIpRklhcF6RX/LoEVMyzHIDeufH8TfMH59ScPpCh
zAY7AaQntrKPi0/T/47Gy8XNlvEuBGnsSDJPta5QYztfQhe/PxHGYm43LRaM
Laxh871y0vmPVrniSc5ADkiaYFtiWkN4GYG/vkUNFaSPCpNso1rVhdmOpVig
5l6DJgpo7UeAcCGUgrN+hyO9f3zouHDmjz43txa/x7mMBAQro4FajXrEmxdG
mNHFO0dB4bE4/W83WhiPN0EFcV283O0UUsjYeax1O3f7tRrahEFPhENfxhjv
fbWl+Cb6LkZPv0yctGtMkrJNGt7Ej9P7hJQULNfIMG+7k4ZEyVz7uPAj1NI/
XtKD+vDq07i1dIYMZcyyRGVZnjEKXLLMAy3ItTvgMHknby7Qlqi6pqaobbd/
3/G26Bk378M9+XpxbWz4shtY0EaSbVm3m5mmWHRDn39ZxL/ht+hRof068zCW
hwihharE8HtheU6Vo5JTe2mRf0s3i5VjuJzFUkLZQBi4NDxZIABdvyb7LjxR
BWnYI8YuWi4EL5HkbUvetFUEOapeBpPrTwG0i88OxOrJPHPz/bM+DjC1JuYE
Y4NWEW6oaWR3V9av15QPpApN7SncBxf08m0ckZE87Gf2VmBq7wK8S+Tn0R+a
BS7LEBY+H33gIlgwtHU+fFm5P7G6a8UVwUQh0godYZ/n/SV8EvO3l8swI+9/
a8TA1wqM4VUyZxA/i6Vh5DBUXH02VQmQKnI/UYa1wbXu6853adzgbVCpwiiU
yXopt5rDd0n09aynY37/c94lcs3iFgK8HVMwA2hAzzIC5sx+l585+dgz5+Pt
xZPxA0T16FB2y1HWF9S1iK726jvy1fIMQhOlECEqGQSIBKgjX/S7TV/I5MNT
dbWMd5m/WuE0Ua4xeOenR6QMQeK0ewPyIp1/6tXm6UU+zzsruH06iE+WLD+u
wSg2BBMSJn9CPApaEMtX2sIa+bnAclLlxZ67WUg/c1eyKOAhF0I/cT3F8WEE
VisIlm1TkXodkUhnkxu+zwmnfjiGWnk9JzwRDMbzOFAV8MsAY9C8YCRiNMxP
POYhNu0/InrMcxMF28O9BNY3k7O3jxzeuV3p9xaRcB3fJ2ZaE+u+kJT1+pgC
FVrfSARmVndvUOUX6aSBdQKnt6OJRIr4YWYV/Y2aZkUHLSD19RzMpN008Cqa
aUhrTcIpj1DVBmApQairP3Ados2GM8QneNxaFVrQyFGnsKPwvyrwUe0urHQC
jcVhWfHdSDg1Lvsvt3z2gfQQqhSXsAQhAOllvsLgRFaLh/hKvI7n01pTTOIh
K8JnyLInuBg6kKuitEkubrGKOQ2hjHIAgDE4rDnCcvlbmOFHgh32sFfgcti3
9Kysb+ne/RYSBEeCaZYygZet4j7eLkQq4vzKf+1BbuSoMcqio9wqZdtGjOds
hVFwqDmklrwUBT5ZAWWh+FAY3DKRFwRTFEMBh6i41KrHmYtuQiPFAEpbVhnn
RfJJqRtqGbsYt+fhlnZl0exv6/ZYMmlvBP8ONEwJycMXvlSbRZRureszGuXr
QtpDISSttBbv24ruWZb/ZTThYlX1TDUnCcOrvYH4V3vLr7Oj9h0jmghHdyOn
FitI3VquFHRtaVl2y2LZ4fAEj0m5xQMrpBniPPBscjwmtOGcmPBhxr/bq1NM
1sJHKk1+oaSq7pEtc+Grwoyx/ZybDmv9qUPyatPIJyA4u1vUoA97vnvPxfSA
Rh3GtZApyXkzgzbmYIGeQvfB9vPL4yNTTQIb3hPtrjAcB6YzO4X/kpjbHPpS
2OSN7czVfq/U6ndVWPJqB5U8D6BebFbnt0zGLwo8NfkBju0hh3PZub6DiIV9
FdzE+hSgBO9ajlvNdo+TOHFR1ZKV6L6oq3/Zg0jtlR/R7t/hgtRgPfVDJQUg
OpGrq7bpR57qRBpdOJa+YYl9VWsp2P9CX2GzsRJ5SBQ0XarXUmkwVGgTfOKl
yW1ForkQ5U81taBpm8iDln4m3Oe5vP8/6RT0zG+t4uEUhf7HOF/Cyg4czMyF
ZVgqiCnrmnL8J7xmuy5/4nJFn3ceKBylpmTQMgBrr3RXwMAn3SiWoXaQtXdm
txdem7akMwXiWzlm9aHzvo3IUxmD5+zm0TBI+kiNdSDgbwNaqHs7UQCFYY2V
EgsD80bAKu/H4a4WPs6XfFGRm1GSyv5GpSFQMXn9kTGzY8JjRXfb8JYMeTe/
7aBziVCDz5dFZd8frBoUZNnEhBdQheOz6Phx3hrGWrp/sxxkOa0RtPOLRUad
pHZ60Y9r2UAMfRSO4dFDV9rRZd6yXiv8Z+ZxOrEoixAVghWy5i4EU9IoQtU/
0Tu7sRth5q1hHvjppcPEKgiHtLPtG4Gd+HPrCgPAMO9uSTU223YfozclHVIR
Ekp+PLDAjg2cPCxdd7G7du1ro7GSIqxlgAmQBZYknSn1fkwn9wbTpAWUH7Au
yK0OKvcuqCA6GG1jZpjdVTTtSabdlZynn3ttcyO25vm/j3vMiWu6HT98657C
dy9KOajqErN6CILy5SEjEbwCkQ2mwxDPbA8bCCSh+Uv4BoCiqhwqMYQqpXfa
iMkI6HH4/+d5F/zHOYBj9Xtvyipph1o/4HC4WOHWIA6IvVTW+q0YjaI+Rrzx
HvyuQdu8JAxxyuYvZEa+t+bXRzq6QL+HPWFcn/JM6O1WY8i+b3soX5/7g3f1
Lv/bl6Clik0xIk0wQDDz+0zNsICnWH9ARahtXkGOEQcra34dWGRTzK4z9SeR
MHfRpkiLAild1UYQAxDAo7B6TLbepAKRsbnSgTdBZ4dwOjaSsXg1VuBLJawo
/QQwm7muS8JfayA6Q/6MjpcsX/ca6AFOs3wUoT68937t7aegCv6eLRFNr17U
CUcZzBrQgmTVypqBImNc5vo9Dd64q3atcfud9vIaA41/wCZhn0RsUd8jdozi
4WZ7X6327ZULO/JjL881DWaScSh4Ae1nA/sDOgRbJ60kyd32xsp4Hzj7qwX+
WuXjKKwkXlSZnVxT9OAGgU7cd2UUi+5zDa8G0FXis2sHuu02Vrm2WU44zfjK
KjMQzazF0k42cEoH70JJOOGdBsOP6KUoYY7oLo2P6Qgz5YxY0zJva/XqUrBI
uz5iYy+r5YQnvU4+YN5iaKi0HUjvg19fkhmY7UuOmVzBapUWOAJ9wPlI4dFk
TKHbSitoD+aHHE6OPSC+XGW3Xees2RlSK2hB4LHF3PnvN5wW6/UguFWeN2wM
MtUr6lLn9srrdujRnbQjxFJgjACi9pcdbhVs+Z5t9hk5GRp8sxXvHtOI+j+4
3RvIdf8yhjWukvybjxLgE3z97rCGTPppqltZ7lJcq5as1HnN3b4XIAvGdqKZ
RxFag4J8V9kBe8mXR4C+SGe9pgXI2CMYy45ubJoNXMplXd5doz/aAF9Rulif
6HgkRDAChJ4LxtB4yl8jX4dTZqStME4p2V97Q8Qfi/Cj6XqQ944Pv0Mnd086
UIZ06r4nPZTYN6kW+5nNK+Pe6a9pWA/xOGBa8nOxh7ZxABISSX27BsSDb9Lm
PrARy6WGdIwQMju/rOijKkxXKDY/7AALXFOiFLmpw9eTmI51nT7d4FhR6Mt8
RYWlOz4wN5JxBOMl/FoJw0yjHi30Zrc6N6V1z2P2B5nOgdHTTILSDR/mLbsX
AMs7VtvrKEOJcgvhTfefIWEFNpSzupWuVnxSelot5ek0ONVbBKigVDv2NkRy
yhW/sdBNNiJYMEOObPgdJ2erzHY25u6hc00DFKyPau1c1KL9Yb4thhNUpNyE
xR0n2YbV9ZfkBGunZhDWsvq5u8mXOgHxUmrS/6B1GLa2zHXf7+DCA1/cORYj
6mUEOkBx6+kdYLqW/vo0LMhGn0D3NG4WAlFgw2C1Crg4Y/zIwoko3yu237ux
Q5wDiK2yHIK17S+Z2yalfUud4vnregNmAkLZD2i23CIcxE3MVzL2n7U5bV0u
WA69iROvVhgDnNN/1vx85oyO+/Y+2uamEMWlaqAZ3+12kCN42iVC+JFyMrBc
PP5TjqX0ifrbzpJ9D9K1VWy5X7+1hHBPkBkTSKvktP5gJKy0RIMupkDeu7Yw
LZk11jIYw5QtU0bQBBXUQ4KhbSYjGEDfRtq/ouaZko6jXbUUBax4ELKEX+N2
zpX7n+JaevjAIyFz6g2VnVNgyjzcb+szODyPe7O5r1A+Ouza7KVSVvSMgX99
cayxU6W+69LsauTpAwVAcusntrgg4t6CzLCKowEfD6+WCF2eoKWgN9/KOXo6
+pjC3sDoNOIUwJifqQ1mmCuzcel9woAuljCGcxIjSyFTa8y52FK+b5HV9CxT
wKgSIpK4N+2/SQaT5GbRkFx0HLGeI8txL3h9tUIiEmWCdr0x1fO+BW5oSvPK
Hqb7djsY7NL1S4kb5yk4+U2mEsSUuLZM+hcoOMgdZHywJDKIPuenF77hXOVH
yoLAsfx6144tGAuLRk1PjWuZHSCg2dsx0xNd5Lm4mp9TqBYgbaCZm+wyDVti
aBFy8x8BrADcQPsx+409MePedmqefXLAx4wG0Af2gDm3fGA9Hc3v7B+MII+c
E1MtQVGCk9or2eUL2muI19d/ouD/BphgaS0CPMlAdYACt+Sc/yfrVtljDtM8
RzoGXO7hDKYIczBSVAsW8e+LI462NTN2m5tPEaYCyf9IPM9TT420/UcHxP5T
kd07VcYYnlxq1I14iVoIM7uoKbU06hGcaWn3HYJRgRfq53uzRIcNqEeMbBcn
1IpJGtAumQMmr3dm8IbaJxH+khUL+jTf1GqGoriOql/ZkHnWDoYVnUqRlDY5
C/Zxa75oeKaz6aSkR/N9clxeBtNhnPtCWSincTDeV0qGlqq//f9VSsHl49bd
KCzZTwpe0Va/HIkMT8QWPda9Lyp7sbYTdx10S4Zq2kEyVybrpHlXYOW5lN/Z
fZMUZkL+cCoZxGpFBxzV/YeqeubjsnCO913DrqmwTBjZp9gS8OOqOSQ4JQ7+
8zPih60tcUdN82u5b3ol6u9NIH36wGbhOX+9WzwrxZiyVJFIbngnU6WUWH78
Y1W3kN3C1QEwoSZHfLgQkvRmuX4LcEzDPKFM+OCkRbo8SAzl4Z1WkC7XAK1G
wES87eyVVTTyyL+GabOLtXveyj7Zyk/WLsiZZmme/Ind1ttizfS6APJvZ/ST
j0MjkqPk6uPSx5LodsUdVrBLy8WwJ1ybzS4ZfD2Umzo6AFMB/7eqnRKFA8GD
Pll1ccFigklKPlv/vJ8IytADx5lKMjQeOBXHQ7FgOrraFSLd/qBn+q1jx8Ku
K5kwvy+mBzEUMdZcamnkjwfY6HHrLqF11Y49VUj9bLBhECWy7vE8PdaJnoDo
qq3t2eXWfRoSWhSEbOctcSR9Yn+L0t0QfqURvDEZ/HpJVOfIbwrmpjZygYMG
9myJqFRD7wd2Lwf9M5UvmJ322BYeQeD6au6kAoCW/xXQcMXvqxCj58z45nM/
34jJ52AAqDylq521tOju63uJAee9k7FeZpHO+2gummM6o/CfWUnD2t2DCwv+
3tbv3vfpn1old11Sov2IfC3xysNdHs3fRNKpaZOcd8TPZqs9u9BL/qU6vBZh
3aEiSzYdfseIFdIEwb/WnoTYkgcJrx0bV2ukvHNS5H3jy2/TZbhLl1fWvAY7
ZRsBEUIyLsFJhfaEAPX6mNObrJ8QHBhjQzPxj760uYxElb5OC48MWBvCc87n
VKhVoVyhSNoJT1YvgJP2afDI5pZtO9OHDajR6ideJ+4CnSq/0gFYGLENqxbn
XtldGs20JncMI3UlQ62XCkYPJBkmQr1pEPGValuOkDDfpOUgkT1X0erjFuRr
3Dzq9aWvvG2nqR0EeK4FKxkbf7FV2DSMaGuch20gtiVU5r7wW3uvN9QTDeQT
jJ/JitpS84vc+rk6RxVIk9HVnsO/OUkqGfw8tlpSkGe2cLk836ByAftO+BoO
Gs75p7GMGjK/ibx4eWakBR0nXx8dXdNfInQ7BxNDVGpIohIC65LhqAwU5SAO
A35CxwaCKRu0mNXDCewzAvAOGEGv7WrcKYknTt4wg5lh242mo7KjvanqESGr
zhu/m8+JdWqHUsYnnQnXGi5WPaMDlz6ALJyfYVGGO8xuN8CP+KrJjz8wc4r/
B2UCvAi7mt12uU6WFqcV5C5fd+Gq/iiwddnA46DG7ddD27kSNOttIVDUCGLz
sW1WnQAwr15AQ7Jq+0R6WHZjo3z6OWsUHVM9bheD/sA6uOjYjLxzG6BkVfD5
6rKyhyoWvw9x///jCLinQLKd+ZCX9Ek95r16/mFvRDj0+ZYvCI0Xswnkq1Ls
NjzESTamkNQJQKZ+sAf0lxqZpgAySY58qDFOQD46CXt5p7QdnIfKgBGk7VOJ
8kMBNRT6moqS9K8s5lQEMXjC3izz3kBtmCg99cKxokr1rvtKpaJeSbaiJOFe
6Gk8DBMIQ0h2pkMS2Z1WLjk/ihzDZOlY93/EZmAe3Jfbhc1/ROJkdNe97cqm
bNVURZzNUUcx7YnKKcf9tYsS1rFsoV/PMuPnsvoySnaaUhuuGP5az17pyoXX
fhQsN/DppZ4kVUMsqIORKcbyQEUfa0QDpY1Iby0HA0AVaYmSlPGShF0mPdCA
RWUfYUIik5U9o4zEZmrjbiiAZoN1Zu/mNgd/P6olsw1BwthzOEQywx/SLaTT
kdpX08AUYYzd5q9rRV2NulZQniBKWQOrViLlH9/ME8OWKKB/HU5yjyngI+ou
QJI6W3AWJH87qUvalGxJU8wspTPl35OI+pjJs5W8nYtQ/m3HbPtGZhKWHfRk
8XlQcSi2rlCwSuFu770aSuhW7rwRKx0eX0RTfNGPWBo4/8vN74ol2nwSTH/B
xCCgcdOwFpmdz5gsIl1GQliXr8bRJiacDOqS4ebc3d8EUxpWKWVlTu6iF0b+
yK8kgBGvIScWZeFguv5PZsDrS3RgMgN1DYMUsLxzrICdsFjfzfMMdRKTZmFs
qwbmh4tIpQGfz68cI+44ZlAFNT552/cDdoQZmzV0yzyAWgdep9XTEHU/EW9Y
52zpQTpXQao6SYjLUXzURw71BDmB4acC6TsI3dnEn4cmxxtXpTW0o8uUlRZJ
6umDbqs2l2IBWjxpSmOKq9DgMeWTYAROztEnJWdiIQKyv01QbaN0ShWvqAvp
cBMI9KhHqFvKuMe8AfgVv9Ppv/pnGR2g69ev4hAor906bSdpjIAR0A5+Yr3m
psmmdC3kYtYzGlrVufzOWKPZ5eO/L9w47QQHTjKQQ00utiEkdqe6qPdwIANx
hYImXH6zRp1Ug/SPD8akygmhPqSCF3NpsTgiZMCw6x8lJJ0rsSM7+JIipXfv
PvmOe7iGqgLq2AvFLWXFKDTMOnAbT1oOGnA2N5tAWVsTqTZYZ1hcezfo02ox
vmCDZC93hF1YS2Ae4PCxawSofyHLt/ayMt6Gf6jwtguXXRl9y4TxIkWsZ3VX
tEzE7FMqdf4HXqH6fzrtFO6gCBFe3qjOgd7fv2H7JKaprHG4VzLEdNDCq/dw
/AvGAz5DFqJ4ZE6MXbPLWD9NjudQuG/CK4ti87L92ZVD8YneWcUY0b33xsI5
RWYrR9Rdkg/R8vLxKmztOkhgz32pA4dRmq0aWoDTk+A/Gk68g2Bia8Q73+19
9ct4pj6DOyOoy2FynvEK7AO75As5MZ266yq7jIBIwLzf/D4VUFp/BvowF3gL
2JoBf3CvGkwQwbFbSpeHQX/n8zeC2/6eW2DazoQs9pD3E60PKPidsCiTOvZM
QIooow/DUuZPspQ7qi4Ce0Vl0UPEzwGb6A+CEYzykXhIys4tw/b40+O2jSZe
Oc5KyM6kXnOxi/zIXRV/xFBer8ieT219RWeI1pfqru4Csrc2XigFZF/PyTky
USsszhyIK5xYVcWBMuSjT/nTHb294/AdQiwJ76jSjyWlHlu/7COV8FScoL1U
z+DHLSpg1wqIqwJOrdi5QwBsP9WNf9t5V3m+4l6rIZHPJwp2HHAVbptph4/x
09ZLHky7SbNZ6O6BVE4gKdXGFppePHbB+mrRkjI1zE048aKA4aaQeUl1hpJ7
UBjNt8+C+14mb2gbTkAW4wYCkFqXA10KSZNMhBhl0731ZUwgWkLY0x6YPTER
C6RPFfAMmNF3kOBjSbvrRGVRVK2VR2FbrRv0QvXZqFI8G+anbyDBuqU/9We1
USRaY2Gfg/7gwgpyuj6U1G5mUUnnngafZxfH4Bb2euRS2+5gFT7+Xnh40d/d
9ayjlRpdFWFDPV72ZRg6fhgWvcHDqMgBCIXrktf2N3pflhEnMVE57qJ7eYVS
lwdfDxj1qyBqMBk7vvl08X1I4ErELP7zfBt9nsZiUZp2TjZ65pfXD0v9AjCi
vlkO32GZIPVP/XmczNS4+9W7sFftmB4/1VOu6n7k5mrPTlaqA5rEYBsfFJX7
qvlmXnQ8eE5NamQm5/bjqOwoB+fqyIJzN1jUPnRO7FIHsFicOl8BYaFMf+Tu
nAis0TEx//AIxHZIXqEwvIreSyesP0hvPghYDKUX3QKvA50b7mCncTeOetAW
a6dPdAEAabirHt7M0OxzBDa3gWp2p2QUnkDEt8vmM2yBGDzaRbY+a0cBc7Ns
YH4GaclbBigleuM2WByrtBTRQ5Nu/rXIYVSBB2drr2Tp2YtdrjKDc+Xigxg3
uJMXwUrHonYfsj/yfbwpDkMjBheJn3IiqMoxFYJEwT6FsEjsRXWrzT3coC58
OFk31+S1JNzHyYWTsxbRHTOkiamnJ5AF7fDxJSOGKgn2089VPUBp5A5td9r2
jtW1gkTJ6sl6w2ILFp6EZli4+1WPvt/Mr4fqnsvz0rFBPJiy01fFAiDdhksO
0GdvSQGFcsENMrNeLKPeFWQu71SlH9cfFrzT+EIzmuIAlD5g9yuWoNKAX9Qc
5+hD5LKsOANn2D6qzFnUTm0OMIDGfTAa9WfpZ/hYjIa5o5A9BEzfzwa3YT1J
JuydOBiXOHBF+mgffyULGv2T1PpEsOBlANKQUYXUFmp0GFy4reKmbpKSK5TS
/Urqavyw+VrF0t4T4DoA9VKeymXpsJdq9hzTqY4diClFVSuNhwhSWLmdH2kk
yW1aCLx5hhw+TKSzwwYvJQUd4xSb7tyTRvfAfU76GI8dLYYZTSQlRvK7uuaO
nH3COgRGQuAoqN5FKyWZ9qF69aedi+x682ahn34tEGw1I7xU4dJLpNabLECL
WNdO0q2VU/ClxR2QfLEOnaPhTUkPrbIVxtymCWWvRNqnV3AFbJW8lwcrAkHZ
HjZQH56PTXedy27h2BFXbNDghk/X0j1MvbqSSWBFmgfKyyJ4r4AuoDM4UKLG
CYqX/peLaN9P/8xj0Ug7030MG9nvdNCtGAfPJ8y9LGVAH0zFKWmH1p2SauN5
D5sbJqpBgf6CwUszeADF8nT9T6oiaFOpMxBe1rrYKxva4nWjcv4F3cc8xV8z
7bWoRscMUqDGDw35nUg9G8zyC+QY00fTACNZifMzTgzKvI3RfKUILaJ/NirV
A8cM9x5/kGwVxYWsrBPbJjdQefFTHvQfbiRkd0bSZ/KyzFIlILJlfIyVmAwV
MVQfitB4v2UaYXgtm6SLLuEf7DS8E7Mc0BLw6yv96eVlz7Go0EUzji35ghU1
GGqKKFzq5uuYbrNlWE2s0mW12o7M8iwHi3RuhYqMuBXBjSeTcIOriOaEjBOB
TolrQZFdWZ3xcTZ+28XVC/kjKRInPoSk1iE4X0bHsYh0up/G6Z4oeqPZMlby
A6jtjbDw9Y6/Acxv3FPAWNjS7L50TybYw2ZYW99Z0hIQcU3xbagtwm64FKhq
aU0hMymFc5v1v3SECfZXzaCcNdMH+nQr7l6hQAYdbDWgHBEHOpoXgyc5JyWF
Y1Qj99q/YGEb+lwiCIvJ4osLPBlboLXkD6gbSMW0dHAzqNziyNtz300ZXC3G
UXkQJd8abG18v3IQW7Xpqv5WVc3o4UZTcxb7sIVaT9LMsLurTJirwkQGSEpe
QBIXEosrZ548CG846Kod2n73EUL6nZcPUPt7mpLm6g7XIRAEe9VDsUHW/iH3
9ML4LncBRiYHMx4Z8iJBgM9iOOWVPwmDI3h0E9ulKlNBcbQ6uUAB27FHWsjT
PwWRGymcce43XrF1WJeBhaNt4SujMe9E04CG/jSbW/sl+KHbSqsrkfMPMMN4
ai1afMdyxzYhDCc9kEV5PHujpeH3+p/4JsYQbHOH8WXOZfe+uKeP8f1DDzIo
sWdbjk2l0CmrVRqsG7iPLIe3CofN6cV1kTTpiLM7W60uN1c4aZN6fMTxY/U8
eE/2Bof5rYHhsKZrXovstTa93WNXcS5PI1t/pqTTx8XEhwaIbrr5tk5safao
JxvrbvYvLY2lt4L0aZpw6StZxwga0jNCuTeQolEwIXJRB5t2XUpSGoOk7T+M
S/MIYHvQqWhOnKBftB2eFGxfl5QHCF3CjWBgsz3cwD/HQcwW9Ef2KT7rrGCW
XQnlH8iLGbTs1wWapZL+ZMLJO5korYpAuTBmVt99c5JLIrGWP49tiKiPc6n+
QgZ8BbE/dKpja5JRGM6UM4g+lu0kZmXRRwWASpjl66Aeoxe2+ZMJopbJ4Jnt
h0p2MmLEY2BKTX+Ug6p2gbnDpNu6Aamb61E/izMaFxMPcSG6tkX7Hb+Thv9L
lcz3hcfU8AtwtRZn+UYeku+m3Qligcr11eyKs04e3Bn7kabqBMFodR6tf7IL
ypt/TaVicOsxUjprzQtBcg6w/O3VBgt29p1KENS5H3o0fhqcQ71M+T4HI0yn
wSmA7/36RHrgpORu5/7IC1U27HPpzVuE6pSfEAtME3bjhTpsBkoBRigB9iHd
CQ0MTzUIExhs0emjQdFPhmfn8iBjkijhP548Zd6HM27lghi+YNDWiH1Nqx4f
jBJ6j2GB+Jn6pf9RuTE5+kyGlZYl9oGwMQ38tNrFxlc3spy6zx37XPIwlhWi
us3ubrgEpIUGOpi/DQU0WylGmSaVnXil8UQcqxAPCjECxfzAjUwHIflsQDwD
pVliAr+iOUSt2DAB6I1oMvUbK65x78slmIMweIWwwaVAoNQvPqCH5mWtaF9p
jN95ZqDRsCGiW5cTCuYvhOtxoM/WDxVTOE2+uAtvxQFOOxNKlzZ/ZlXQBHFs
SieZgUUyKkzWYi7pmvDsXSdBg1a0lTk0gcGgMUJQgeqTJIGNRQC2KzwdnsDk
g69ixRNfyxuiQgNdom1YUE019huZImp91gaNQneYz4mFeuA70+YH3x2PGND0
H0wLzT/2kF3V9IAzXQFiOcxoYj6205Bupp6Raz6hgkZxhdkAWKWSZ8OInurl
ogf75dCQzmviI2sT+Z5RC2fZ6zkh6kICyQRPPTnETuzn4IqXDSLO4AX7DMzs
dbB+qRYGmE6KwHaUhI89Qzew+72w4gsLy861F1eL21OyCjm5zh7u3Wput6nZ
9TkMkGoECkwyUBdsuXVJ5+ApCE2EqKMfNfSRb+PSYhvr0Wizft8ydGmo43ni
B3w+9grb8aoXffEjg7Vdv2SkJ0Us8IOhB/F6/pl6cp7bvKO7Scp4D+4zaOxG
F06+oLf06zM7oyC0BHEdoF+cYf95LguQyU1ct/9CJrYgazDP7TAugCRgJ5v3
7KeFHvXR993WN3wcR7iK9O5kTaUyy5K0/JnBfH/PkQFufZa6Wnfbl7qUBp0P
qz5OM6FSsUrrM2DBKTdbOyOm7ZMUsGt9vm+EDlPL0PEL4dGBvaGMAQqaRFWv
dThEdUa9o3azf/pHtTXotj8S+YnIGKOEnp+gOGjnXjy5cIoCutF7sf8JvBEI
Tf43phCy9H39vlGyTZkxE5hLRwslNLT6svOB3gnZbUxLgOc0r6pP/UZAOZUN
WZhwXWLzg0SoNj8P6Vevoc2GiufkWbxswAmEz0ZVKBwRjizegjLC4hcJ/0Hj
KRSp3s6pWeI1Y4WW+BbwQHih9NhH066wtpM/XwfqAeHeWfHXEw5yWnTlNgKD
+fVdtBtu8VQIbOarcOFFWxxea8A/x2ttrYLbJFFteTFox0uHNi9JVybW6Hia
ZXTMW09aupSbtDa2gZ9qn6z3+IrVpSTSOzsWnYiIwjUljF4RzZ+cdEqnjPVd
ALalw8dK1eHdM6wIH34ulByJKBuGG3cE8R7Gf3MFqYZF2vN4ChtdkgTtXb1s
12Drmqkj8D+FTmxjbam1rzTkpV8oCIHkLDD8DQEDOm3RX5aoRTGVQyG8vkjq
KBG7PduVoAx9uHqf80sNHWkE2S4trhXXPPGe6pCow1SYrzsj/0A1s09EsHwF
m8BbpMeIPfcZIDJQjs7qHb70utw+3CA68TL5bWwE+DRXNrYpmw0OaCjpNwDF
tdekaTax92T11LO23cm9gBUQKhdKy782oWRprwJ8z1DD/dabbHL8RqCh9Yyx
UfxKhNYS9fb9E4urVG6eM3QO2JLgsZYG2EmIgFPO283+BFZXW2nEhREzjJi/
BJkS3VFypjR93hK8aFOruQFJ5DSr6e1/J17PSkCoXEC7c3IB5saBiXjoLs+v
N2yS/0KwJ7c7NsK8zt0wqgXpWUTtcuRdLf0oM46df6EXHex6Hn3/04XmCkJ8
VCtrk/DNDo5Fps/s/daXI2nEtsdTpuhEhVFCOf3PF5xpSWSB1pWW3tucKHnK
3+M9rC3UGCaZ/iH5KryJDeqb/6oyRk6xthEALE6A7q01rF38kVWPe5zIxLqF
byEAbPERQQ/TWLffnItwHY2XH8W6JC+97T2w4UsC5avsMxwSr0J9j2H5L/AG
2NYp9Tibvj+CI52F1OaRvmI2fJUcsJUKGIuQxriJ6VwxURtmkwlDLxbXgEeL
/SPNKG7q9dtBa56/oKSA32YaRXo5KEICXlbed53CqMzZ5J71Gcc324+RcY25
xIy5o/R23kbASx/sWJxfXMLtu/G1gm0g1wd/jpK7cTIQvpQRkgQFcGLvzelE
JR9Hbr/3dpFe8cE+2tpT37K0+iufjOLWRhvDZWAn4fbzhl3vX0nMLwKlwIX+
4WDJwEED81tZql5MmrW5wg13emsZhXUl4j8jwYAdkRS0d+hTwx8JG20KXffE
Gpsm+rWWu41pirMSLDEsKTNl6sYueMdbNWJARi2WFvDZ7WwVTep9CvEGYFEm
nBzQ/qnt3obLe6Z32cBcB5/xA6LjwULQXDCeYQOy1577TUrNHGTc+MEr8KCu
9KZc8uxgMx/ias7DImVkkXwpU2XzidpAJGzXJy0RQ6QdEUUYsSQ2tw++5dpJ
Pcxk2L1WyxEolbz3NRn0JyLed/z/2OPSxSeYlqaZLhycqem6Ph7NiX/xAdo2
LOIbb0+3A3leHUV2J89+HUkhTvx1+PhPoPDy9Fn8jePcwSBhKUeb+5CeeDuJ
6QAr1Uu6e1Jtd1Jyp/ojkvE/0bSMU8veyONB5Oc+qYa5K7daCzYvMksXBYKt
5tsuV4UMkWKkbIu/NPCqSgyz/t5eTyslx2EWpQ+ScfgFBXepU1Xj4O2qOLSm
LUMdD0tg8syh3qM2XZTIhCcA3QWfwyRyUFuv0l+NrfNxioDA+ac3mnDGSi+u
DXF1YMfsTxfNdZ6cdmdBud1nmarwBtaqm5xV2768RpNJ2uDz8lYRuYNR7HhS
P053arUgKrH8AddVVkV0dqM7KWDAaI2wKRepEfOfZH+0B/r9SrTN5OOXZF8F
48UYLIyBHXHFJJkqdx7gKLO3y6+C2hfBiPGhZbv9PVQQjlEe1ExEGtf9jCZY
NR2LYfV+4O9Fl7pyZbX1XKsByOC24qWngjxbyfWGxD1rNn6habi162LQuuJo
aU/HfAaCVpwZ2FWclz/3AjqpjO6jldgYxidW9jWP+9xig1FnKYWIjf+hLmAv
EI5F7d3gmgv7rrk+/uWs/D4noa+KqZeeyc4tIQdfYWN6ujj0ahfxVt9r63sc
iMZA72ZE0fhHaNu/zPKhwMdAWvnceZyNQn1Er7TJB2fkZngDNjXl5tSyqwxk
kpFcg1o9n7j1ppq1QjvfXNtYZY1VDDkGDhFUMOY3ugvDdDqd2rDmloKyJw0Q
dhgdvu4R10y1152r1UJiROoHHzW/dSnl0P9Y58OYobUt/YQrcLGtfEFC7NaE
4V84lmmHLbO9CFghxFKYdGILsCn94L2e4XSUD1j/Wvh65N3jc7sXpGPP5Dm8
E18pyOa71rILEpyGiWC2JFIT30jPwAInm/4V4MfgB8vhlLau6pOg10Mao/71
cLeR2K27N3Fl0+WRHofX2xHL8oBEFAULtrmUiibYhAoTOcnn1B+636kJcT1l
0oViHF/ks3Lz1Y2m5gxK4i4MfmlfUW97RJVdjX3cYG8/YqpjMQdemXVejrSA
kPrQuohawVUKxm3J5p9KPMD4Kjb0mkKpGcEmy/cXcwz1EDhNP75wMJKi7Xw1
uP8qtrU2NCcT1ImBrkqADph8sb6/6rKxu80RcnD8aLOqzkR/ntfCqlOXk4rH
5DnhB5G95XW4lVhhiqsAzf+JCowJYMKD0rBWjx/MWuo0doF0M8A+GLpvEPn1
6NueSJV2DhVe+ESPhTMqUV7eV9LYe3VUQwkZTabX8WWH1DqXR2nRVn4+9T5o
NUqWKNJxfauNmMBN6po3jZ6dly67Gyyf75mdlR+50F6Fg3mOJ4FGqSK/MU2I
JU7XJk44oTSbDVDjHbfERrome2N/qQBo9ItNJMWIDlQq6GUlzrAltRAy7U7i
z7KALhFujxsJ2uUnjad4bS4N6Sdlq+QOYV+GYl2FdcvkRq1cyGs+xX9d0SPR
FLWCp0rDdhyqgEvE15TUm0FsKO5mqCORwWHXYldk5lIm94TdSA27FERPPC5I
fuKPTw+coxLt2mOuE3bCGkwTRAATEWRtsHS08Qo/aVwghYLeJ+Fzk4pwbwqX
lTSi5/152xnZbTFjbu6bpRl+5GRWYW24HS+/9u6mJWPusXZioihDu/BLb5cG
bhPBKwv84Iav8Jg5yiuRx0LDqeTyygfuZ1HY64uZC3Fm3VeuxB7ey9kq+fyz
b+aEz5r1Lqc/rGAmgxTH3/jJrE0FY9uOiBSh3T7UmMHJHEU5Agjx1jHZLOnx
1shnIYyldTT6bUiwWhIczWgjAXsu9XjGwC0CPO3ExkOzqSQlmLvPmQGt50QP
MgzWb4Rc/s+hIR3zShkO7Btu7AUGZGMnVy5fQVpFz/9W4y/rOLoCVw2tgIPL
tfM8OUa1sVSiVLqbnDqB84vfmiG9CMu35rYUdU90KqXKSeLne08zGALj+8rA
ZvLk3Oz/K9qzMuwFVwgW9V/bQ/mBQQ4IkCkr/ytAtO5tIls/1/klFm2mrzzd
gu6fNC6bZ2TP3Qf3uNRAs9MkEVT6yyd5OH8SFj4rw+6QsRM486AGVgnXpT28
2GrNfA8CgUj1d5R4YPFbyA86TmWxcAaogE01JzxgLK/2f0nNM0nr8w/DLN8y
ns7+Fr58yg8vWpRo46DrXGRzOzsQL8DMZO3W+MdFhbW0Fi6BvknMwrgqZn2L
jkYFcr343DWkAphxT6NLqMjUDggORcILa2SgEicUfO2X0dTo0t5Q67+s7ava
yrrQt5JY4/H/IbHm5ZVYDC1eaMggk4IpGGGmv7IeYrl7kt9C7uRQW7q0R4tz
Q8URrLpMBGr85GIVr1ztdE0A7fTH4LxSyfO0/GlUaaUqYvxG1icjvvCvj0XK
NlV/XpD59f0t98QnyBywPQYTQgyrY8rULTI0ReeQzBhJKM8JVdOG7t4tnRPF
IqB1j9IOVcX8nlH/0QLKsNHZHvODpGBqkD4Cvm1Cue1iutvTsmtnYEQKuX6M
a1x34p3saURkNpsh9roqu24QHXS5e5Vxkt/QJOOvi3LBoecBZ8gJleyTkoGi
CZMamBsGGJQLyVfcvwcgUPeoQIYts0SQjTcT8cqxrsc5gAclnXSLbQOc1sGp
93vmbCPcMSx9hJpjAIwTYDA/E2YOgfbcB3XTZLroYdpJpjCZSDmRlhivJUcM
MGe5I8/54llRlDsEfx3yftXe78fZQSVlbR7dlbYxjsZ1tLmkcVqYNyf++eke
/PkMS+CXC4dyICL5xbQnRo/h3aONhpj/tevOO0+A+GPkbqfvbrLnjs15VqJJ
QxgvPya8Hg4+YYN7Fzl3W8rOxu8vbXlTjdApR9N6KHkPmBdRFThaU9+mTkL3
xCFxtzSmfbAf2gziCx6G9X8WMbZqN1bbvuoi/u3af67RqMofeUETP87exguy
op+4Jv9wJ6kaNMS9yGW3kvadCjtuPhFMBzR1y/qnofXXsVYCjqEOmf6WZMA3
oOcFccd/vLkpXe0mzPEzveuVGzyQJg2WEcq+c5DAO7yUhfazf4aCYS+jp5zr
+6dNix7a68lZbKhZAH3qf8/WYbuljveM6X7l+wGWleYK5H0uOkHbL/hIOAoD
e8x5TY7yUaV7kVRFqGwqpU775Njn+ya3fpEEEAjPlBvAp4FQqv9hqNjcAS7N
QBgzK1cfFuiA2BMUY68bEQyOKTYwiPg6lst3cx30XM0laHJuliVz61xDaFGx
yFheEkA7qhAwQ4Da+sTfh8JqBHUEmboxSHlU3WC0YoExAQVUUxvDWHEUSHnO
DFQXYekrh4RhWi2PXMHKfwaTdFaNBsn3ExPEV6jFSfyKcoj+e3MjhcC/zijc
LPcRONqoGG6Ag0FCxAJLmOPJwoNF2G6omPo0YwLilvoT+h3dela3YhVZ0Da6
JtZNpZWuumwz1pZtE0uXVzfeNH80BNpAX+59+sjI/06R8ku7xVGfqq+9EpkF
K5PvTF3kZjo127qYliK8PTTbDZrCXwL5XcLrblJF8b0pMtV9gfEmuqHZROGj
P55BUH1HPR+ExcWTc4zI8eEBpQBxGxwlkh1K85KGcmbC9WfRnnSHx2FQPFA8
7VhnM4945GZYe8YIqbNRMmZmUhEqai01nIktxUKrY6w/8dOiPzL6jhTfwM69
5EhFz8AjjzqkKMhgSM5rfP2fcO6pvVEug4LeIHLiRIO4TNh4dEGypzxsG5ee
nvNNWm4sha85BHYq8/1nFzDrNn8UIha3nxHR5PW9ONnTssC6AKucfjBYUALn
zle2U8FYdK2YpkNcWlF+Qvs825ZD7otlLh89C79U/ot5GBETDLxLX6eHlnvf
QE/iVcR2gvvIgnz4aKqKGW8Ew2kBDGlPRKhf1+/iQSnXPkLObh5+6gwhinCG
bZMTlUMj4kp3bz/rT72cTLB0N8iNktH/Aw3EDoPhGa8Flwh0tBzP8V+KpQyY
yKmTDjdD6M3WXnigs360NQcNw3psfEMDKESwafUgagGQ9Kn+SKIhOAGfJb/G
LkWzj47z189TTxKWGbdGqgeCsVNhEaZsViah5Vojo2Pe9R3sKLuESubCF+3b
1f9xDNByEBl+4WN10XW9hHmuA4ejG4RunQgfTkIuol7VJlDTzoSjjw2zAiX1
6ZQoW3kLf+7AP1ntI4fTYr4JheKxlFRR6WXnEqHHb0W9iD7yWBp7XbqRNTle
dJovDtRtCymXDFwT1dtNdOEucit+RSUWgVyYjbFARSY9N/JNquOJpcxM2Au7
Xm1JIsdmO9IYx98fWZydAs6l2ZYA7kWzFb1jNOcvMfkqcaJcdR4xT6XV/cyw
nNm2itXbKaTg5+qLTq7Mm2WQ3SncqUq7CWYbMctQztDBdbdxRzgTs3M0qalX
dqAOYDoGJRBvOEWqPCVTYVIno3abrV72SF0y1FSvB4zWWp7h5b47rUbebmDo
9gly6+IoHXJO9C8UUC8CGZcIbhUiRXynwr3Ay1NYeh+B6dyDwQL56v0NmV03
o55qY0P7gZTeoE/PwDYzpk0MOH5ojbzrc3Mtd1l+30DDyqNI25XWAu/WwZpl
Vw3Pw5EXRJvRwKjRVqXwM1EK1kWmncz7xKGEeOjLAn8wpDu2nyxYgcdt6D6j
HUmVbp7Wo2wRZtMNO4sou+sfjGSE9xlq1rGthotvX9WNjBJ58W9dqmymimYm
S6V+D4IhKhPOA7LvNy9MzipX8atfJ9Oi9073FGVWaLp0BXUa5KjgWik2n1/7
lUw6Re+Xzv/yM1IsjhFk9rTHMSCHE2MFXYcWGGQIMVFaTpFmpRYU+j9lfH2f
3tPrpjMkQqEGKa2uCa3FaGhQqOHEWcy0PpdpuGmh6w4Ysa2+HjhH4y+93s5d
DVfatSqkO2v8x46FPMU6rWcWjdJuqWCLNyi+NIeL+DpvrAa8rsyKvNXcKPrR
/BZsLpumhW5aLCvkwx0l+43DTcbYNdmBrLG120POkrtBruoprKwPCP/pRver
yR2I0twc3cuYOW3vGa4A30xRy5bM1JDfgcdicB5Uftwz1yMwhmNjSki4jeNC
fxVIRwAwX1Vv+uD78v3ZoWhuxKQiGfdTlwM/mlBdUQZCulSGCeUPa3hO/7og
Oi1AW0+xyrBseZvbomKOdcCp+PvEEy8yUXgbAKDdCe/K+g44eJnUb9eAO+sc
41wWwn4yzIwkL6iAYKX8TvmZNlOXVknUqersKS/rZM4kWs9SYPCshBiZA32i
oeJv1uJ+3WJTz+8kLX9HRWNZZluKmNJ8IcSVN/w7TtmJoWfl7z+LKyjfc3Kq
ZF+RxpuseI98duCSh+d/CW1t1rWKp9TagpPM32iagGith3ExpSS6JDfG5aRb
n/XrIGbX5TAvdf/wAEKy3MH7rGo3fJx9YffFtnRBBmpI5RzjjnjN7RrsaEAP
HxwS61kyzg/roevCn7q9w+sO8s6hfS53D3F9rBc/YlQLPQvQlrNZ9y+pZ4Gi
MrYKteUnxGk6jQpe70O8D3TTxojTIKcffPC0zJ6ZWncwDjbJ1DjdU6PnAz0Y
hSEQ8rve1mQpzr4OIDkTkRVBbDIlHkWvTyfEaIvIKKr7/1+LvAvHSma3qP2P
WfqYslv9GJHhMrQEnmWzFi+UJGPkZB21kWbq1UG59yAlkjV1l7JrNe6EUo9v
7OEsFMEa4Y6DlTRCTDeyCQ0DxGmDtxi+64arYAgBfSLNhSgApU/AgirItJhO
zieoOq2dGlJualH/AcTp9lTLuyJvYBEaPJ9sLE57PSY78b3ri8BSr9AtRj3P
0/y6kUt7wgwWawkunetJ0oW5wDTGCqf7rbUDkS2g8qQgxnQcJ7cIFyWwg1W+
XxqD4Z5kG3m4+ud120eAFMstmR9JPlkH3sIGF2jIb0CtekEhOzRo0eEq3adB
Q5uW6Tx3wzFhL2EDbIVLvag6ZmDKbqNKCHYzQid73hAeCm2y17/v8dBnTgUS
HeskkJQr26t0SXd4BgZVS+F6K0ESvWTzLKrls4+6i5lNfxLxiOgg34J0/pyO
sE0JZDr30RLbX03j+1xhs6zq2bihnigUOjVXeiZRkCC5CQGVjAUkY3ElEzym
AoF0n5HZfsSCjAtiiEY9mLkmArAvYO2NaREz68rU5tFsV/j6woQ4+JhzNs6i
NYW2538bE5/aNjYY7dAGqZLygXdd/AJYpVFB+/HnIjtoyaYXqbaunHlH9AZz
oPCoi/snV5EP0jJosmzUO6kk50QrcTXLmYc33VHG5XJfUPMumYV3cMgxqaUW
iAy0dxO42kCUSaU3S47aoWdzbtJ4w5xqpGj8jYFNDZHLI9zv0ixMbUAKlxDc
AjzzbURv47S99oSXumx22PuoG6kW22whwr7X1vPmGIpLONw7Ant30x+FmF4x
3EDiKk+fkqBoLVRUCBxMMG81rHMiaUfEUAA7NGpLra03h51kwVi/SCUAv0hE
y0MelBBL3Iy2YUym0ix3z9cRPEmXIfMcDPcntWey0kyXAngFQMg4kAKcvMyS
eIJCCYHZK5w3NwkIu1xIEWIs/nXxeIjSq+dd8SwEpyX76S1vaj/+rxYkfXFx
NcOCy0iE0ec2ryRI/uGXTE/jUYNA19/bSTsNcfeWYmuyt6HHk0MIrHA4Sapk
fEWFxOQ2FP8sOaRKfGCAao1D0cIeCRBgWd6EmhwZabTNno9zmpThTYOhNZZo
ZmhLUvYjUMf/QUiqjK3I7b2/Nphmhmgb0/wfFO+wW9OTlRKjCk+vLnQbl6uB
UcEtc0uy8xp8eNEFTqATvq1Uv8I+GJDPBjNPIpw0xQ886sfXJTS1w0+cfCli
4yO1nZMS3/CqMKNoKBeifTtFy/ePc9GWKSUryFO/uk+uvvRR4phiFANdI2AI
NYvZzcvoAID7q2h5j2F8hVT97uJXaqD8Ci4Lw4rL6bxMUjwNnZ12NJWkPvzT
EPp7Zx3YaMw1PgPCFLz4Ix3GJ4dEpBjCKobPMZQ9ivHC70HK9ch+Ii15xnG+
H7dE5fboUTA7rSrvHx/zzHr6v1GeezqykjLbbyahbhNW3TnUj0eiSlvqQqur
6cqWJE53O6TQ8VG1xI/D3DOzWDeGhxFH/XnX5WtVgBYHgLi4GEQwEf9v1Xzy
mmoG6xGknStDL0bYQ7qo/G/mwLhRkxfdrsy796hEHQbQR2PtLT9BVBV9AEZL
6ozFuoWa2tAiW4EQ7H51kXNSVLTmxephWYWMK7qKjx+fg+gOVG4/gNIszQJf
zOEBCwEYZj2Nz8EiSLmy0AHOeQmmSu9BgvgBLYkU28PCYtgWTeB02kGpqP/J
PqNgwWyqE8su0nCA5TFSUvwEf1IFaeNdoS4BR0kOzj8NSt3fMe44lG0NYi1W
40CPl8VMzfD9yWeQF6aj4RjZFUknaSs9KlY4ntXIXzn3p2khFptAi2cfjnxv
eNSfOEvZHAkst+c4mrwvw7RKUxXOJyA+22mi2XzKQk0HV4mtvlyPM4UiIbkk
omwOo+WE2n8dczCwajW6WlFvwKok2b1w5t6Mpig/hiRwd7Y3WQkuMYi95reL
LY+RreLSXzinRfwwsQALq1gSf+CtG81DjEyJsErY4HWIJH06xkLS316AeDNw
YRIJBSzd8NiTZSUwPpCn2LnOwuUJgZ+oQDlLJv9mlEQ6drM9OsxIt1WL70pI
o5xolNF9VWMmmC+T64pTTuKZKypdMNm90/Tjc6j48KS3xjod2Qo+ylCCMRxN
k4bRcbPMFy4zoJaFvHiIfC+gkAbtvSZEFqYXbJBwYtm4ugjH9Ro5goF+P+A/
ydeT4f8aLqO4t68is4Tfy/ksUQ5T8zhVjKHDQaFEOFeoq+R1yhUpu7lgm0mP
U9seSGAoTjdDbBVnAU1pyzmo5FokIKqigqV7v8AiLi1PwNS49ob9TbKzlPrM
IXWxvRdOWKU4EMaJRjBhXqk7SvcwpP+meW5fKwyEciR9VP5Xg+IIi2HHrCbZ
Wd3y8lJjz+xrvoyJpP8HCY2GLyderOoiuUKXkdhIvyIKcuNqNfJvrpOuucO3
uV4ysrub6gTtKztWeqnzuxPZppBIDbIH39bFW+s6ZP/bZNEqxeZZm1+x9Jnt
ItJ8IUu8zjNUtlShbVype7bpA9m6H78QFPdjYD5ISF2yqWDkg8eCb1y7gT1w
wdrJM8VV2B6+9MnaL8+A3BgcXSiVfqRewHyyGgBi+QgoAamCfL299Ohp+8Rt
iKud7SiJAK72qpJMB5x0Re48q4fLFxu2xFfa0zOfKV10HlN8JTGsG/yoXU6f
yHZz9rVcIgVUnuhhHT3CTxrqgXWfrAAtN5cL9AhBSXogd8+WhOI0mxaCUcv1
JK5X/Mk+PgTcYeBsLaOnRd4jQ48nwPYfo8vu7aN+G1+cb4jpWpozDraLpZzt
kKFHXIjLnRNZLD/9fEmoXXXB6iqyJ9JoLwQX9lkqEQXvQ/M2zUDc/LwErf9O
tut+xYAExvZHUs78OHjPVr7grdjjuvzGfxCMl97bxAZfUixw0IPs8L+dUa/t
Ja7XHpx6i1X2RFmYuFpkoPlSxn8YfRUvlyvy1ZY3cZDb9D++6TrvVxqZFzM6
tzYIJoI9M2GLdmO0J8wb7WsMuJGpiNJjzk56xCgch30e9mw2F7zWh6iJxBxT
pJyCZbFU+1taRpkKkDr5bIx86P1buoV9bnSDNNvDtn8cdN1ww3Xi7SOOq50V
v50Iq3bI64UBZdJUkjtHtHts9133bdUE8PlGuF04/8ozzyYebfNQ6NoKYVef
GWwhP6Q1ZL3VhRYtw42RbLo6npmY4cEDoWJN16EWocaJpmIbCZRHJVv7BQfw
bYrsqUUUAQFx6JiVHuyS3YnNoZkcxPJEgboFYz7NYJzTgakmY9rZClSkdjYZ
0+6lPAlbyeqkXBtpUBTkuO9nvvM2d8C38v/IB0g97uzi4mwNz7heG9+1XxH/
vXOrbrjy8znMiqbndYODy4usLwE4w3Nma3AdV7sLqVPwVrjMfcN8lbDTqGPa
avhvS2zJY1BO4f7AA30D+gfm3KHgYayYuNt5h1MmUaAeRQbzbrYYdK7RI4Vo
UQIrhsx/72CFFGK7FZ/NUHXYnNN59Gevl5n3YCBWcrKwAY8CvFrH0UFM6Zsn
hmMP/51BkHj53hvQrGEUZrnrK62U0gOFE9Gh3ewHfAzc8WD+e/0O9x3YYVQ5
iIauat5v4tPuFQGsiFos2NybWQkqLdlawYnOlzjgJF1aDoqrMoQAJWS8tMvd
GB4FHpHVM4OcFnpml+omufwhRatEJOQyqms3XT8uoDLfnUv3Ma28OIFhauXy
x8XTMB1+aV96aKtZ9fF5bQF/POPNcofEkUXDA3DGpSLplZPChNO3JFbXodTk
esDuj/Dr/GikOhrRFmqhblpF1hE/NiB6fOawVudVlrGC0UTS3KpC1kOX8F9O
VZCVsOByM0KWCbphlWtvzAs+nCEIhVVTfPeks+r4Xs6Kn/EnvQhvHnuQupRR
eM/2sS/TX+jH8WNcuMaHjHLgeHqTQJbG0Vb9RVNV8HtfUqr2EhPFkTNgAz3l
2P4oi1tiKlr508wXljAYb564oCoqJLKM+yhCUOj+aFF5B0sexhAbztO1Dvac
/IWWOZTQrYaQWqhE+3zLfDu6aJhVFAezHhVwxvHYgCBihcIuFnqf077wCTCS
YI4ew6CKE6sIGnmFcjMuz0sMYCf9Mls111FVgIJ11cyfCQad7fGQwJdUtOKY
ltl0BKn0UuDbtIzCsBWSQiWe4EXGrU3aJFlyivOjcJhJFO/b3RgWpRrx2ilj
Juhy1r2jb9cy5ahoXBub3pEFnP7M6P/qa59witys7C5YxsGQPhMPh+KwrA6E
FNXClnbjTpMPHakp2jqOyxaWFK5wiVEWQzIGGaaGb879G2hZ2lJa4xBJH1WS
MgEBHWIWVAk3M6YaAGks7XPMpfKOYMCinEfd/6Ki/42k+OfBtlYRdAgAs3r/
LuCbiYuUVhJEIWU2c6A/crrVa03yscSdyINwKSVRBT3RTzEL5YpNsgjetAwl
yA8fuuy4juheX/lihpejWDsfx9orBFINporxClZHUE/MNulwOxn8EUmQwWqX
j92VjKpuN0oqecGW9J8yzXmNX9puW8BxDa8DsFg1O6MZf6W6hUZ4p1wTvk7j
hU3D8vhZdc/PG6EaK5Q+84gGmtMl7oWB8b5dW1COu+9ZQZTkv2i74yPEMOw3
2SCF5niXWrmu+W1H5nGpTMo8JyUmc9FPt+Nxs+/vUBVzqnGMmhF2Ks1veQS7
7zgnoHFuiDStzxXg5buiwWAcX/xBMEaZHvQUNBsXZdElPWb6AgyB3GJvlJKw
neJ0CvQHLqRgZaLxeeegwkFOuj/UNGGvZXLMqCVyWUQ/KF2AF1C/UUKaU36E
gzXXLjXrt7pWyS33MJOCd0Zw/e+uC4nKKggbh2cbQdzN49OGWObILZrfhD50
dPbGvei+yn7rsagoYsFoo556UUxw6beaU3WkuuT856yo/aIAxRU6ORHQUB+2
Y3DJJ2kmJZ9fpSWZE4rbHssWt5I5uxZlEPN9JIZ/hwBZFz17Tkq8eQkgv8tQ
Xoaiqw9vADWqTY7e1+0jhERjI3Wd3Mc/VHTCtLLPMeI4nZTQcU6OMnnOAsXP
iWYm7MEDdIK9/b48mnD/Nku52PidVzx6WQh5pOxqOHoozyPBrqdekM45z3oV
QgaVYSM7SlofkW/Nyom9ZH/0FUQAovCGDe/pHGk2JCNMeGAAJK9Y0Eb5OGtp
FvqVCf1UDnDreY+ztHxtBcllmFeRQKgRZFuiHQ5L6miVMNTJ+ci6yNAJQ19R
2xE0OtNvDFD7N41Gom33azKKaBcwGUyy29SIhWnq4x47KSjXWiDMNSHUVc6v
dDhh4a3B03OQclCpa2i0AHVFuEiqZK+Wq4OoViASOB6rjtH//sApF9+W2YTD
0SK60WRxxFKnUF94HCUXrBsjyufD8/17CHP4jyoNZwXbwUonSoo1Q/17F/fU
5BjnhZVHeWnPxMMcAc3LaYZO+OhnqIx7t9KwOSvKnmWN+XvY87mikligD9tu
ohDu0Z6a8ItV5iuhkRppJCqNKmTMj/MHzTaT+jYcwBG/Jm3bAuW76rHwPEqj
KxP6Etf88dsCYDs4VezjMbSgPswzkeHX+VLVOF8/Vs001BlDkX8a3NGmn2WL
O+ide8b5bOdRI2NtgnwqrG1nWIv+g8a65sePrXCC+LOfRAUAaBZk+rRxcmKF
1x6YPQp4oH4kD4dCorGUDXfkz0AIywWvTAaRqbvMvbCBSfRfcIwPfqTjtdpj
SboWENiXYkHQfsKk+c2Y0vYHH3DMxeB/4SawveXt8I72w87N1iZirbmnCBVq
dW9lhmdZBiv0Rjj8QwnNFNe06et12svSzBhdQnIYbPj6hK22RfJuWXO22w2v
eBcuktJKauSj7WECj7hvpUr5jS2OKRpIQJ3v8Wbe0yGAXKA8Ruvl2R9IOA44
g2XbdXLGOLp50WWR1dyDAwmWAddUd1cH3Dr3Hg0DSeajPlxrCs+FHdy1Kn2k
64rGv8k+9Yc0yIYuH6Alcq+bXrjRDX6LHNLNeqWNUDvvnbpZUQ7c2lLJT01l
67SsaMHubO38ED6+uc8k50AM8u9/3Z6WzHGofLkNssC8rHP2hQQE0UCvKDEG
g/NiVEXeXdQtLjSUKe856U6n1mAPbrVaeRwl9yjfwr0rJrvWtbWOQNxoHJEI
5r1Vtls9sdFUior1okreI1kjMcS3BAHpThyRaidoppS8bgTeJ9fecdQo6Ioe
stRPxDNvd6qFJSdvY71Lb36QzmvqW8IJ/eOFTQw4hbSIu4Gu/yiqC2E0YU4+
MYGFQFY1LGvrtPlkcII1xJkB5qQ8KQbuwJmOwW+xQN14XBCHdDfzQPwqwUVV
Inc+CA6h4jzKyLFao0SJ7NT7k1LUpFjei7pz9thf/CuZXHLh7+I4guXbJ5PA
Ciucs4KXRirC7/r540F/m9uXOevnB+kGaFn29wjPnTAxYrWQncG0LvKz+b+D
U1fZZg/5TjkbAYNQIdISS1hTukWnvDFdgR3lKwnOUaV7m6qVYQ9RrIoK0K+g
ppvG/BTs7J+FtjdnBxFefKzaE8F0cmCrikN1FBkDVzEaJsEnQ2bAEuauJ2Le
gDBJ0OpBDQvDZJmz+YJVeeq00cFAPRI4QQOvb+G2ctZyp4J7mhO4rLWHDyJ0
1CIhCh+xknmiEqVKcK/4EeNX9C/lJnNUgzOm74rLhldaj3Yok9zoJjLrJ0ID
cfIFJvQMDvRNsNzZfk8nDK1wL2xA0/FsqBKIuyPZr14KHg8tc762VjrlEQ/q
0nwjs9Mdpeswcv/zhY1KL4Ht0g86Wzix5XqUML/0QlHLiWVM9bLXQUHlTokl
kdRmrpQsvoKUtaadKzyunohFCZbdagx5vJW5B6a5czOrtrIpsrh8Q1xvyhNe
jPPnENj4NYYnlQdjQlsnyMUvJdEFSWUooN5ltIrn3i8dpzgN6LD470uzShHo
SP8oDZ4h5SIgD7uwChBGSRmh3X0xFMERNXSEoiAqhLS1RC7RfhN16qmjY190
zrQpkzYPN/GX285/ejlr5Wvrgh/bOn/R4u+Vqwwu8zgz228pMv/75qJHmPI/
L9bL53bzWvH2ZS2PryLQbyFtINpyIvjggK1XRFhuO82QZ1bkwRqRcuwCcvnT
Dgh0vG2Bere0vd6+6kM2SpB3RdACME92voQF4R9mEo2BGVVBda9UGfZ5x7oF
1oK3I8dadP83yI8eB28rc96cdb5C7NNQqX9Ee7LqwLkcrxSvxGPmHaM5aHTj
jSDeBMysv5zreWYDQsOF3O4JASUAt4rG32ucW1ovZa6B7HFH4dYr1LaxW3qv
l0q8pE8K4TwdqeHzOoq3rcIQfUlo8Dc372DvjgaRBy7879Fkd86PrgpQBRQF
nOpUcmEa+PYXITcumS2LuEYn86KZLm0+NIIh4MmOYhDxgiVpCi1J0N0k2bXi
6g9NbYSKrhT5JZ/DRsnOJzngJfkRsEU6g0xpoyl/60/PAF/jekt11B7YGf7V
DYFKos2VZdRIYrxeqEyXv95C+g9EMjQIf3Do5LPq7FPwvuIUZmYwKdcsIiKk
hO/CbE33DIFj+kVYHXaKkf4AepkaXltYEFrnYSRVMhAhbebDYcOKEZcn1qbI
yEMuGbeI+8PrjuMzoTiZfJ6gJYlNITrI55jluMweTCdAh/mJUAyLouMrrbDr
pSYApRrwjiJBrzjwUezjEgMve5cpun7SmJzf3vCdlrdN0HQWGLYPwRVbX+Bm
oSs+AbbsU+ez9wc2dWOYvPrbRS9LQ6ZRKhpzD6O+G0mmkr1vjYwYKueoYfAn
gv+eJhN53E8U90BBltTDKKSz933Fgc+pbzj1bS3R9E1RAy7150y6zruqtdPj
y6hi2I2MRw0ZQw2g8i3N27xZAGPTsOOVcdcmuS08VdkIzeqqzdF62qlVV6D2
TcmIvYSy+so+UPQ5l2kTVIIbwZvZ70j599etdqoeIaKDXbVEcI+ElrEkbYzF
GLg1kvn38SuZg7SPENsSrvIt20zJAvJ/UDWI0i1jmtAr9fwv7V6AY80oHeDW
4npASqbHCfM5FQTfCk+bZcmuSSAfMpgFNHU1W6zNkMGSrVsR0nw+A2Fh31Fx
ZdQfVm7evaehpSkTCMRbwEBnVqAOmQ/xEuBpyp0mQuj7aRZ2zsDE80pyXnQa
uQ76aXINGF1pCT2EEUtvMDiTyJs1Yn6yDvNN2vPeLoaUQG28RPDIvMI6XEfJ
X0O5oAHS+94Yvj2rOcn4z7zm4a2J3nxdkh9CHOSN35YOA4hiSUbk+yabWk6M
wbyJ4/4J5kRhQD+cjy3OmbsU39GvUlS8Y0a2y0G97r3Hutq5q8r/dJvJt/6C
ahL2RiTIV+uyTb0IphPCXCB7REp0lT+IEciRHh0eddg6BfQzHi+PBcL9dPYA
SMZu7tdFQ2BG0cPBd21UWWfDmJGhEkIGVTMcH/u6loFOkOqVfAjfHt63I5H2
ONxpaJxWSdp5jFo195wsjRMBOLOzGOsUa4FQ39BHJP+BpZq+lr5wP0iFpJuY
kip3bFSfprQLh140PrZrZYL+NaMDJ2r5U8f/KMho/K5thsmn1IIVL4DkZRqS
ra3rehmnjm+RjF7UlX7+3np8CcTAkh+KaEZ5JCZZdCKeKrp8OjsWxKLWR/Qy
V8LA44kjPU8iOo8HKcOguh5E1ahXCg1H/DIL2/42pF2tfxJolaN6YSpUig78
VL9NqYKYdhvw3sclrR/N8hDiKQ2s0JKlQIDbLNHDvw23rci8kZDBhzVJRgQQ
h8q95R7TF/NHPkcdlKzHgqId8C4fO8IP6msKObwOAKGueLgoOoMj60VtCamq
TXKKyc0ocPOvriF99S96wBdaH636H2uTVMYJn/xgprrTQzMX5ooK9sPWSbiP
EkXw3D6WIyOkNKkuOmVCpboV1jQuiW/GnBwOKa5snyzl/+F15aaWmnd/qpoK
+OFW2hob/TwPqRBMTX5XpfEuv2C/a88Q1xLOPls5mGV/AsUSb93P+TSgWvku
Ousik6ACMoxxeMVH7mxNmYcqdGKmzpGTFbP7yr+YVjGwZrrSO100Rxg4SrWP
D16ZEIUP/Kstv0xQ47TaMOyaC9l/guDb5OJHFnxtyoCJt8txWF+TSD/bQGjy
GpEvO2/fErtV3pMo50lbc9lMYhiM/NjK+wUfucb7f2yzS0qeZpKcDY6ju0ap
79HA/1v4QIVeE8SOzft8bjN+dlcbjT05C8CzWFz+qGwbrmy3xUlo5+PW52ZB
eTOfr1YehlwIpIDGQWVqQFkCJbkFApuOcx2pnPu7a+tbifjBzOa8yHfs+i81
K3Fg/c4+kmUW2dd9TUrpXU1cVAgJAiLIt6Wxn5yC0CythJ341bUBbnDm2qHt
qIJ7eA2dqduk0IGyoRHu3WFAjf4aKV8PUn6emBug8P2kc7VJ6RSqWhP0omAP
NVed2yKb32F+XQHWkTwvCO22yh1d1gELmvKo7lfcXDI+h+XsLcLSR1JM7516
CtyQP7o4idpble5lU8AFpFfwbGMo6I0Er/bOe2WtlsXLlazzn//20LTCBM/B
yGyBdiRlKXZsedaBob/40hIXPYKd8EnuAkVuaE4HsKgkxlF2AMhrV9cg4zpi
JdzUj2gMRd5jR5gqz8QYRJhsd5OKd9wQlsR+i9gzoW0E0m//yjk+bpvqx92v
JpD8nhC/w8ADLs7HQQRCo/CxAhWa2H9ptsrlYJ4oAn0sUvGtKWw4/tyUn10C
oPVtHGwYEaNkA3pFtVTdoSR8By07jBAUuwp21Swzh6SnI/Y/2JdjFWH3h99V
pTzKTNgpq3xWXjHB7/V6/Mpdps+kObSUYM77e5q3z2ySeLgkDmHpXjRCny2X
N++82NvZ/xkDNEp13Lv1oASneG7DA72weqSleBvpEMlTQMEVxlUFQ5CxarH5
+h/v/57h/8l/pP5exL9SwbyQwaxCBvbrzLmNpFBWEcheo9diztj72owCdj8l
yDnGWvDhFEa84YKQHoUt4LxKAt3QhOV32KyQhBeRxLfM2A2SLphoerkh4puQ
Mh3gpUU8IByZrWLV4cfiwPQQn359h1lwc40h22cc0ZcEozW9smlhqSeLHRlP
XnzZ+O4T+txudEbGIef9UFv13yOmKqqXKxxJLgEfCYhVRLT7EuJEeWvo5bla
cS1gC1WoWwW6MWw+yWP3+lG4RnA0QRwMmVEshu+ZqKNcXZqkqO8vaJNdwuLo
smgsIFRc0e+glKxPV6OmKaGeRNdWU7ZNN2vBu0W+EczTg+WE4P8E3Ng6wgzc
rMFqpyom6WQWBNNP/PAdGu8DzI/WRtgvRUD8WPbw1my3C0m7FRyan9WXeQnH
sjdNLgp5gIHVcRfkyWlUrEJgAXpouvZUn0mKikK+y+aJuGSdlW7YCQE+AxLZ
7V7CJHOr2mOqmJKRAcwPERu9XV2V7IAjbET6TfgQJxUXuuO+asSnS2qWnvsl
hClfE8CQ2ZBSeQTM8+0bdJ+R8HGcn9mNLBtHnwFgnKTlNSHVlbBcapD+BolA
72TklUtpKytv92fzQctLLvwhcii5VL/ef77acfAfvDw37a7iqVJEoEQERcoc
jdh93Kc9iWY9jA5F9OK8qsFX3OnFCMJ7X5lVBDQBfPGxrvmCn7u0Jj32x6Td
aFhGvAiZeaO8bI7wnYgQeePveCTi3hEgW9H5Y9hb4/2o3S9icVTRVqzF1MNN
/8x8EX6Dukx2se1cFJKRFAb8lUpycHuo+GQNnF/1do35dJkVgFlB0fuT2Lqi
I8pDsBPiquGhROzriYVtE7ex4NDSvL6a5ZArR1eGs+wcRYX9tFOQy8LdK7Eu
vMZeNXFY9Go3Ks2diqxrpfNkAtyRZFNs2X5D9Eta9KQC+ub2cTTJlU+O4501
SfzWbZHg5USfv/hWe+JLf4nxd6OsHVJhzRJlO1OICKd5zoSe5VaTQGehaKuc
zYG90MRc/L+P0dbi+f5goIjlkeBEC6dM9kSb9JBBuJoXgkooy8xMQ4wAG6bZ
GGAZ2FVRYvRhRfj18JM8boH+3zp8GK37iimqwpzg29D+4wzU43B3VtgiShWo
1Bb0AMoTpFrL1d8RXn3LWFe2MUCGUieMZJErUUdkInXWMZCau4Agc8Yb59e+
aDZDhVj7WeWvM9wJVYs554UKRawpZck1OmQ9RBBYyQYvKkQtLB7S0OI82PmT
u5QiSqcB+wUTcxXE+JfoEIDkPNnDyHkb1czeH6PDdBr2fIUpf+/mRC6WMUp9
mXJvrRFnpvlW6eZ7XwbNoy+8/aQCwQI3X8A6ZtqxV8E8L3sYU8bCzXbl4bP6
7YZcLT6JrKknBcBN7dyBaIjeWrcM3ClZOMrLJHFa3PTOrmEzMR5OeJx6fJJZ
XaKiKjvFWJA9DiA07FELR1KpXiAhkHzaCu+McTxln3zoUCFnjy4mxggDAohy
38b2bkpwYjA8nKTl1qP+/2hHGf+Fc7xPYz9SK7w+93KIkymb3xOEPstH1c9c
eVRyr0bx0lgF2e41ecaxPiZPFEj3kPjTE6xE5iNL0BsBzwAbXbaTYpcvhDam
Lwtmjd1sVgkcP7VdmsucTncv8ZVWkM2Ol4RXdVPi8pCKBEWGpr/L2Sids7/A
3+ro4DUmZj25Zk1VpHEU+Bo4Vrx+ScetkyFCwWI+pUsuvfZTr+ZdEKStJV/9
hUW/9ITKSrD+9RSPgRcTvZDMOxrej218KNEEUDbOUFM42Fy7fCyI6DOVfKjq
6xXYLKfH5PwqKGRLrE2sePnFFAQyb9Zc6Cag9Z8+17a3dGgbvn6ie1tMNJIr
o+xgKBQmMAsYOXW0UrMohT94haXoXPRcvUj+pUo9DKPcGGw1NmOyfACxCLRe
udirYvdyFNjf8jx8+kMUOOHdIObU+8R4mEiEph2k49hpJX9rovU7lt8Zt3Uk
Lqww69DUlB+TSj0K5PJOGD6lO68Orp37qJlEbFSqJaQEF3aeY9T0ffSKelxQ
1K3EHCe+7WS+e+ryEoayNSoi8re0iaVkAPksg6fvE8FwhIRU7EbsPsnh3cST
tln8zZM5QdDtronI8zciOo5rUZ2Xgj1qOQvbftjPlsB2qyS5AUF4jbDHDODy
DVQ+r4Z19o2ZaI5Xtdo9h5ZcpfddhF1XS6yOxHAXiquyqxbE7io5VjD59jeH
sHUUpn3CNF/Gn3G0iPGGjKUXiRMlBlxlBcP+Vs+yE1UzGQG/xVRGrqDWfzu/
4agu+V0cY+3q+m1C1yOKWOWqKUQapU35bOBd5P5AJP4TMhmJKa/++hBuPxmw
QDvoD/6CtPBNQPXnAz8OFjAEE7osQIJN2uJFND/nwY5Do+OmDO6w6L5lsKst
AjrEpbmYPfcD+TF4Cc8m9OKGv/V9z2o5UH5JlhCEAMlOVlF7dq/3t8aDtRaN
aPrN/HaSBQFB/50cDMH0r01x5FgbyIwnbI3+k8A6JiJtF7IJhKbI4oHzIeiu
/sfl9BpAqJ3yqJme9VnVQohbuoe3dsfYYfnP3YAP+Qlfarieyc3k5nezIm2D
cfCSkDALW3quIEpaMdq+nWWOFzd7kP6Wp9sghu5GWdE8dOKxPSLhODQdoj5E
ova+dCbayaJkwrScDJtw2ypGy6zT/FA91pWbBnN5htMFNSeE3kijuelxd2zh
qGuRY6r8y6lrAze3k9bL/nyObm8z9n/esJi1N68tBZwFTaph2FjzPDoI0oTk
GJu6GPPb+sRmlrllQEKyr6UHcRo78UsRqM+VdTYEXOegnhDCMmBXIx9+ZpoE
cjQS9DFeP2Ff6NiXiTL5So/UhfJyNwY52CQk1/HLY/748OslVns0xHAmcP3C
Wy5GrSllmDxgQGwGkwiBqCuVpafN12yIUSW3qN2ZakV+qA9ofKGCbPqL1uDX
mQy1sVQ6v+WhJE2P2DuCScY5uMPfQz49bogYlFiGA02VRxsFiZNcIAzQZCCi
YqIi2i0zORkR8Mp9GePBicGAVYU4rcIzNwjVbRalVRgyphSq4Va3ILKeD0GQ
PuoIATXbA1yZjtB3NA2Opf4eyQSujlRzPfBPBNbOjm7zBUfz9MPb19QBAjNf
+Fylpt8R6Jqm9hgNz+ZwpZTdqGKICze9gxgYL1I1RBPllvpcWjh+fuQO6tNG
wbzBSqQFI6SOk1EILCmhJ8eVbfb3enBnq2U7+qweZdFTwABvPnej+e17Q6JM
yB6cK9UGi7CSHxwlfFkVAtXN5isd3aVwk8rHS+REj0D5lsjjf6GCisWJTJ6Q
h7a7Oe1fWn/w+NJ2aQm8Rmu6qj6EThcRvdXjUEDYwb9KFEXhihDjxII9Wf7m
O1FGwXq+G8mLCUZQ1dgXmPvHORGMeBB9yb8hi5IhtZGbMNK5WjKjby+VStJb
LxvMVLiNgIITgTlxEzPfIHehjJYR+LhO6hmCPxv6KYXHVgGbjwpYJOSWhaEW
nUo00mIa+F6eZkfX0Wb4vZrPecK34qxZHC3RNmOykAOVUNt+NCKqaVJE2fJO
XMIDPX+5ENoO95igQvgfPsRgPpw9RG1i3VD+6XpfjS4MgazHxsRY9OoYbKke
ztYg28JfdUC4MDf7TBbeV4llUvlOQ0gefK5+HawYP86OOhhNrNXdQDdEnXGR
5fNgf5b0uA+K9uS8YveIgFnzIpNnYg0KQBOG2A4x8PFWrQxRdpXcc931hWNv
CSsW+UDwEXbO+9CsxjmrzE2e2XyyvcFJOkNPmwsy3GbAH4amWAl3VlD0KF+c
WoKWwpo+A1NXTAA5W9rLxbXGOYFzeyKS6f8nolE2nWOW43e87rYLtDB7Olyi
slGkcoc+xkBXR8ibRGUBPnteZWfWsPt+7xfwRnf3YOxlmC4u33aLpIIKBbpQ
OsnMHAJP91bKMmZjXFJxd+11eGz/voae5a19p/ozAhPgawevKTlBI5JhFLBd
/TCR/bGJMAqG/NaL6fVXoV/Lsb33ePko/EbhagNpl3zKLF2+yhVMpGZsIkfY
RVhdvi9veMYn16jAzp9+jRgYI5vE/AXtb0UkxCLflZ7i5JDcBke9semdY4Ks
lPGmnPlx5V7PawErwI48IJUtcfL5X1jbaroF6WEBfvnrXbRDcIn6Ga5hTBO4
M0lCUZoMfrLCq6ffUNQ+zm97lrOrxrGHu4dPnW9/dA7T+JQbH1LE2sLfBhQE
fMQPb8uL19FW+Xo7ySxopGcQ4cvhWNrsD875gGE5Qf54g8+kNvFfYElyn62p
maYBmNoThdPpfAYSt822pG2cRODrHBCvZ2SM2ANVbsUxI28uV4P0oXc/Rd+p
myvwlLuKtadPn5Sq9qRvfv8JwZQ67x/NN2KUQJ+wVZ7JrPl7f2vYWMCQwVz+
Iy+9pVHWNMcyhpy4AFW2ffrsEtJNMfgt75FUPpFv+GH+ZbBhB2MTd+IsJxGP
xVM3G3+NPoACcpWTDLLMzbRQ183tALAjT1V6K3dWe1wzLzaCH2cYjpS5H7eV
DegCw9K3XFGNB1F2d4PPifa40YKGkPkVRkYB7HmI8/CCXmZB4ekOYNtJxV0P
x8/g6oOoKWMCfF1C4lKDYcrYp5OjVAMyHnlDi1/kFznTMatdHK+Pf6FHV/8H
ZL/oPGcKyiwpZPUuQp1FRMaIvGQc6M4EpKFE8S+EQS25aTtJpxXvYAdWO303
anVvar5BB1uYa39OpCzAYZdNoFq8YD9PL7ATjte2hta8Tumy6z+ednFCIL5A
yIgxFbpH7ZBz2NWzo8y6td78n54dUwiYOWoGjuZhS3j3DcdBQUuVnzpK8lCV
m+xjpoGQZg2vGENvvil7fpZocu4dPCsFX4ZPX9WrMdPH5LrPcyeUPtVN19LD
KO+ciLIztZ72/a3RTqopxLn4gEESWFpeDpJ6KBmVV15PHghcfC4P8JATSHkN
Dq7DFfwBKh6xGcIkRTc/8kQEA+Ej0Frmn0xORb7j4V3QW2KYtccB1TD/VTqe
I+K3rGCr8fBAFHiOaXJUsh6NZaTHmwqQ7Sik7QRO0gZMuo7DHEnTUBgIV2Wo
RH6bvW19v+O/+HbqKHFdh0r5LYAPwy25hjP8RBp+NxNkLtVaTlzfS9ChxVFf
KaK7v0+02vSefxvsXI74H8EgQaYePZyMOJ7bpXifXZN+zXwfQFtWSuu5zxly
ny003rR9nbGSl6K7ex02nDS3vFL0WwgHzsDac2JMWD+Xg5uKegyx5BC4ldRo
uXdUVJjij5jVQQGD9Ars2YP1cFzgxo7Cd7Pdug7mXBdSn6kOOi98Us+isu+h
Ikb+D7MrxTpgpZnF91w6PKlgaHCCH3EpECrJzef24GBfoH2lE/Ci3fxLjLoS
BgjpahUHd+dLsKagToU9A6SyMHgCcngIpk8f4WdoJXNKzzlHkOiVObDs9/F2
t5Re5UVh5BJEQ4mYLTAJTM6+tz99Zr5zu5497IaKuSsRkCxBhd3k9sVDQv13
AMzbKJatdZmEXpBQhos6gZk/jfr1WqpXlT+kVsw6nVa1C5Cyk6ww2fL3kinT
wZhjqIBfjdyRrzcbkSAtdjA8dKPV48P8hTtjmp7o8FplV3pYjV5khLH+j/uj
1O8SarsMwoCxURDnpbYVyAkYKKsrGTR8kv3cIuIuCDNXBi8sHwlNpoT6iH8H
ndgt9zgO09IyFxNGuctyukOa1BegV8QCTazHlGFhTwap+V/+onD0O2XduvFs
TrmGpM5oUVA69kBKY+el2tVECt7/G4JphtwoSXKKhC7o7zVOLjWvap6ihQ75
qPVyhgmm90XRwD9SRVDErBo8L0HKn1xMWcK7aMp49oXsMCztaSw86UWnlcK+
awB26kpDCwWgrj2wgHf3ApsLqvzqMxSVur5QdxXzQDoNXZ+/XL0C4A++y53H
1hlA/3dcW+DV0jduej0qxMyrHlo+d3XGPpDB03a8saS+p5aOU2m5QKHZO16S
+cDOQMpCZxHBTJdRi6D+ilzCzLDo+WFSQQRVF8gUP9TzPyFBpP27HVv8/E2G
j4l/zunYC57mt6XF7TAxpud8AdJW9RVjQBCChuKgTDB/Zo7vVqZ8Vx5MQFV1
owFZ9LVLOaJnRW6mfLssrmVZ6CPnGd4IPrIIDD0qMAFiWAtdv6OJ9C6R55+1
+4y5rx7gv1rjFmavqdovu7M1vN4v0E2RN1bYExSYDagjNW8K++FNgqExiUee
l/rl/6zox2kfJRwy245pNCD68a64eD+D9s1V+RKBg1ZsP6LzO5NhSxIgC3Wq
KSLT8G27llMr7TBy8XPYaQ/7Kkpg6N0pNHdVS8gcLkTtqe+1LtA5G4/nWyKV
hOyuUIqcpZAbAkij/yUdHt1cbYLV/p9MP9KQiYEQOTdVWoKOxXjkzKU88TMB
5WhgG7bNT5GKfnYMVQ/MvdUJbChqZi0+Mpred6EgXF3OoaBLRtwP7Qk+VSGm
ON65Tc9lgr3T4EiDaECMkyDOqH9UPcVNbLf+RNkDkCity8T4x6KCQOwNTgGY
FomY3kVl0zlQAUNmhMe0hSK9yF63+wbF6P0aD0lm1Wi+No4pH6AqbDOpq9lb
JokVUrZNi+XfhBbMmIVhcnZzlaVYafdSwOoH+yODe+zpOgpkzKvd4rkv8B4r
vpEOvhHZe9tUl00EebkXRXgCRwYBRXTsuSuEsbeTFckM1qv6wnnEbVF+VK6g
URZd4VDnXR46JJV+7uDAvAtgKTcXbcQ/bcMGHO+GOYA9ErbvEXgUwMKE6uBj
vCpY71FkpJthzSF/N+J6lxGvzihdxUC8leCG5haaLv0fdK7QreVSWw8PkctX
1Zu06qlkmOY3oUvlCnKMU0R0DQmdYZwvZHxeTS61DrRjsmCEs0RsUKZXKKYV
IsJIrpvd2TxUEzkMne+o5FV6FgnQD1aN57IPxLnl0JyE4TbJK+NGJkbTWPnY
fcKdCJVUkZrcNK+vkTae5ECQ05Mpx3UeumE7HfA++cLQKFCvpITJ2svCc1tO
A+eZURTzAvuLYCalZzUXdL+Jg3qKy1HB6tqkHWP0q00mdtrpRaqeKXuTv17Y
Y6YxaqtP2Q7Nq6eO7hEUm2mJKWJufPp2+jZiA/6dcqwgB5L1TLootMo26yGq
YhP9doGbnGqdnzAbLNRqwbdK4xpn0RpD+Y6uxAuHwPqBNE514ifqI9D3uisG
QSd4RCXREJQhp25mIKSlgNVGFKZtCEtsAwsLQkMRqVkqX6AP4SN7bCLLQbld
XrTwvEtsxbzFpz1HSttgKq8THgPcxs5New2o9ux181z0QhFO5DxORUsBTt8G
U7B2jvE5LM12fDQd/7Z0fFWW3lX4VMDOKao1brRRrrjW4kxuSaBLcFOKUFdA
F50mktleh8xfgGRM4E8YlHja3ePrYqrjNCvss/04UTvxdmNl5r4NKOhtuvgd
rB2eBvMCtxSuAZ4kmp4tEv1eHoEqGRzvrZB/NILiAjWzRgLxORHMe94RxlrP
L/ulJUZdYLKldnAhMACVb+4jLUfSAwLLqC+9Eu62DjDjQTj5csBoH2lo+DPr
zA3QhMx2RQEjooOy79iRjSvFAKsOIVKE7u1H4a8JVsnstoLo/Mo+fAaXtpv9
bwPB+22/caDcMymvAWT75o/G/f2FsxYSR73tDZ+ju+KuLcfZLsT+Y+fOiiHT
BKaUNOPKUuZtDvQK99Y51ekiUFC1U0tCRiUnrAqnxdpZYarGqScYe2+sv8MY
uOhhIeDmAQqM49xqQUdXWfmL6xZlrZ69mJNXPuByCAec1KDX5zUV2Jg9Z9o+
noi53LUoQvAGA6ye/Wjt/pM/mAtKqkg5eQ+J2CaL/5+q/oqlua5CBwVIg6b6
7F6Y4R4s8vSHaQ5WIxoffhwhzXPPKSHJfa6c9EvTgY77/rx8520Snz63jg5J
2NCbeecD7UoAohWx/2EvCMwjqAcJOfLvHzDXlXCMV4NoC/ynS55kX4tUArc4
xBuGt0z08IfKUjlbZaiDU5Q++/MzRX8sVCpavWU+5tRviAVAh+OhYyFUOrz1
uUmrJTEEh+qjBrbBQA8nf3s7+/B9BFPUElz88GXV9aC+/5kYNaOgKlsopetZ
mvBOufK0PYW/BiC8rB7OL473LWcdTc3Ec6aXHeJJtSoXo5fIDeuSB9+Pf2mn
61wzoc259TpWbh+CNpKGTv+bBXBeW/kATCBLAX5BNSheuV7HnF0GaRaO8ysy
LqStCKPj6ci3C0Q4bWgxu3eFb3nEC+wYKZfSVkm6pfmqEVeNmYBpQiHlatnB
Ft59GKKoT3xvqxeKJ0osDlcO7Q5AAYsU3lzrVBXWu82qapTnPw9dej3wfx8F
ftlK09Sy7sc853WVkEM6rS7DiHRuh53qO8kFZWwpdP2gfDt9AqaBkUcUELRq
SAy9pAsIVWS+mo8HNwJRzuOGMC+TUMUm75RlYnaQg+kygzPGzE848vlYGja7
6oKRWOqIFbHYpLidLDrTXB7fXwqW+e+jPDesLw+XmTjiUnZXyB6QkVO6DHGx
6bd1lO/A/7IODBjBeEfh0q/5nnIHAiUTBkJjPp+KRM2BoaxH5tiMkEVJxcYo
huOUMa2dL76CnVxzeds0QPE3yjCtgkoSZaWxMz6Qle0pzHg/6wJv4TPT5YCW
/7RFaHZXhRc0ija1zMt/1BAw78BeMzwtS3+AmNacE2OEAcZ7rrZkj287QMvq
8DdDT12BmNE55AvJpj+Ai0Xv6eLuz6XJoC7CIadrzUYJys3joE8anlINDRpW
8GlGggsWPcApLtCCLfQg10Aaypcz249LrGHK6y703I5VjRQv5XgaX9jWBheg
TTBF6TbT0QKWUeR+3Iw+0BRN5IIiuGT8RZ6RiJ+9PeBg2ZIGre1wM8+dDGjN
2kombLFK6wsNOaO1uWXsIKaDRkIeaEbWjGObOxxkaJDrOp1l//auej/dQnNK
4ZHAyT6kbpyAbxpSD0gdScbydNwCPpSDPBFPvKbiIxjOPgfwPZH9tsXvYK7t
C/0qRzgUkiPZ1CUnblQZP4/WVWqJE1kdVrQE/SKP79AdMsL7k2SY6GOAtpCC
Id25GuW0o578jTSsPNNUZ8uQQAxeprGd+dBnQkY+cRXFO7d52jhTWgSlyY4c
AAwGG2L/4uBMbjR4gn2E4tRcU0vrv9ovzzFqWFLmInjl2zoji/ZN9VmWZXYN
sXdqF9Eh281igqkf/P49uZCBKNW2Pcseg+YZSNGZ6DE43aWiGyry8WozsWOz
4dkkOa2hCQXnqd5svEcormBkyDv0KMIgGUQvUQESmmnvorRiXCl8AQotAGOL
L+2rSLqpgiG5dIQQdJiq7+chqtxTn0X9W8Q+r8BlOG6hXvowu0XOuIXGBYS3
E6snkuYEmRuFimVs/twVUlx2F7kXWXGNZQfVGP9t03JzHCHXLFfJ1YJPqmsj
HIrkcZmCQNre/9FV66ZMmZW3YpWR/mGSojrFdWLXYwjEcWagjWb0NjhPu8YZ
nl8/4RIV5bEJyY6qkisqbTJmv2UNsCmJfS7R2DATRWvu/Ie7VEhlpZA+jW7x
T+FnKy6PpyGmcJmQYPubM1ZAfdsEJW39JGsL0VD88hkV0XXKM0Kv0V32DP0g
z9yGX8IKdnXrUpJ99mCMObGf/CjX1d0gUfUjB24PyGE8Ysr83mKCK28h4swC
zwu5TSe2lJql0kFRh3zjgD0dM27rkP+CelLY1J505dDmDiwr8tqbsRD64ipF
HLZkseU8igHcoK6/OcFOZOWs1819b3+k00bF37+fJUVBhQxo3lQxP1olE+Q2
BVsiqbdySjmIbJ3rz+orcNgf3iZZqiBZPGAlwp4bukx9u+YG00VrzJpZtwXc
WVYQyMhMjDqqP6PXbY3AXBnCVOefxSrwoJ7hnfyP3QLIYDAf6meyHSCNDCSX
tlrHot/JiIyVxMyWK9FzsuJfhM5nRuZ/H94nYbu5gJrUAZONZOmKKNMtioA6
GWrBr5y+XI3bVbeINEtfGYrneFC88alFo0JP2MDDD2SGNy9eYcjApvhYKbsj
ClfATRnMHrUbUDvSLE6Ti8sWpSRW5UNNMC/ncUOqDlSWVwcaSndOCrP4oCWX
6tpQitVooPBCa1krV3vGQlVtf3U0YFzSKgUQ+qrIHR4jw/MiHyEw4fKyQeoQ
px18hfZvhyVD7CyvzUQJgRSFoIg3+QuFYF1DYu+0rZReSiPYG/5RPAOVU9Ze
eFCjBJFjA7opmku28vQMwA4vddva9iveplGvh1KrC4pf3GiMhD0upe63lFo7
3oUR6px9sXT60pm19Ud1CqQ4NFuvr4u3A+nYdQXNr8yTawk2O1tnfXMm/xQw
JcYWaKTh5h4UDHtc5SuUL/KwOKJAXw6CIobJ8pmTld015oficbwBeckh62fE
3vQ3cXkUOzPWqT80NZwmRx1kyydDcfsMrZC9m+T8IPqZPm9vzBO2qHGWsNZn
VayDk7FQ1p0gn+j97uGdW3KewjAwTEj7O/han4/7y/NAslS4t9W+TuVCSQpk
4Vl71wBSBpVokMmJbvSMAf9adGKBdFuppYm9MoAAVaoA0H1bbUjM6L+oaiWs
C546pDthLeWEBtx7JntG/todKSgYLfBuq4tk7Pt2J8/j1mbvyLnjx/rlrYoS
UkZRMA5OWHHguULxOYKmf1bXzh0OEQUxYpPQG3FYofNZacMna+CyJYZO+Y+N
LjjlghafykJjKmvmFVqWUUO0H+KhbWFU7j7vv0Xv9B8Tw/HcEHcDYTWqyBEE
kx+ZQKngl455cOBkvdvx5UKtzd1jTMPdOWlEQmuErskrK0U+3G8IHr3ePhQE
byhO6Mq/4lGdHO5Q15HAGu8/bFHjzOty6g3KubPtqnAkV2UAOqFFdRMw0XnX
XEQ97qRJEETcQJkmONY+9o/Bnl3GGQVif7BGI8etUcsrNR6mc+aVCSFUnHsK
cnPldBTL7eU/iK3kl1Zcy/jvs/6tR5zByMzAZDA1+6CU2xS8Qwothkve4fbo
i64cszetTdd37bfxBZx3GdmV7wetAHv+DXzBFsqRewnuJJurymIQWK8c+qty
TuiHKcJK4oKf/bPJv6IQtw1Ly+4nM7/MXQjEfbUuOdlsYtxXtHQXHpjxtEju
qYcWZJj5hRhy4mByV1RlPBUqpBaxCclfMYU8AL+pXbqNogL7ivh1e/o+OAR/
UL63Z9HlGgZN2C2u79vWbKFDBb69WKcWENs2YdmqZuXnxivu3yJcUYCBYjdt
rzBE2XClI5SY5YsrDcfbcLj56Yysi5lwIOgXPFj7lwjNKS0IXXy+gkJkQUFK
EG/tTBQIWDS+ir27hweZgXOV5tK6sMnC/8A3dvuCOJo4Z3uOZOBfXfvAn6hk
/jxjh07Ff51ZM/fjH4n/cxzXidLE5/50LQ9KiRe6D60CmpxpdhvwwxWDOyJN
Q4L5JbO3YhigBroDDdrD2rklVtQr5IhfBbTydvrC4pU9WIf4VBF3ij+S0O2m
MqV8y5QgDa/HV9tzFOgCFI5FUkH48un4Z3MfXEmgQ6fbU1OunJLMKUMusBn+
53tPIQwiBNb8EnnERsIyPtTauo3MPV13fsJg9ThTIm/XLgpDVtzrULoQWLT1
gRYucfUnC0P6kqn1N1B2TLtu4Jx/+yuJkqVV2P0jHIJmxs/ps0OxuRY4FIRy
oKCDLhylWNSNI94Z/ZqACD/W6Z7lI8YiJAxOiHeiSphMwS0vbIDdronsFBFU
c1c83Jtqhgd3dQXNsnFANYJcxACwwd93UgcGxEqde+B8ZwtHT69ncjd0vB9B
fc+MwOAqkegcG/vob9EHxlt15D2jXyHjc4iaIfe+GrNotLWRX5nPWn9mguJk
l1spQ/jEzhzArVI4CMeOFu+YZMfvyUifE+aKiozvnU68GmjXP8H22cT1T0vg
6pVnvDTuINhlXztO4VxNPFmgFxcIn0caqV4bP5DwK05tzk85NDaOimO0lJpR
08Danh+tayIb+bw7WSImZ3PaSh7m1mwvob6xH8KmzucSud3ofE95q19NVJmF
kCEYtlQ5SLzchDGS4DOmQaViUrizZMhOfdbiWja8e6xpMn7h8/gplJrUIW52
1Qn976QMlmHWvATvF/2kituKbmHrn1y6UjvaDNBBNbvZEdHfLY4P/JKYz5UP
skIIGRFxgiXdK+ygAdRGWKy8oCmPr7TpUuBLZzRkA8jQx58v/G3uWsw/ulb/
ft47OyMU4qxENtI737OOIlPLfXX2jKHVC3Rb9lfrfAeK6l07RlNmTFCZqlRU
lPskYqp7Q3w768RWdtC8/AkMyobQ5FgXWraUzGAKw/q6FVcgeemGt9W3OHph
0nF8sHNS8GCgPIFv130ESw/o6MSUMN6HXLmgGQ4XYWPTiIqmVNFs+5HFjddj
sBBwaFrxoPGS7AMSWv/MYEh8aCjPFxj0wr9iSxAwR3K2sJjaVFHDDGPdOkCb
ebNBAwtgYt2U9t9BZ3+pXVLnfxAZZi06ajiHdPiSeuAZWRNb3XsGGovsPGMM
O93TclNp7jpw9ln5AdfoWxPm3ID4mzivVrWV+E+xtoHAlBqRbnsGFTUK4h3V
sI5lw9agSMJ0qKbeQDoaN5lAlNGQZOJVkSxX/HKgOwXZP+T/ay6H0XGFk2/y
BZPq0bynVxfFWLQ367SNBtdb2HxNqbyv9LbLlAdfpzJBz6IVdeABgvU6Ec4o
Ix2YJ2O16eUD3mbFR33Tj0Tz1ukVH6EwLlsqaSCN0xIjbbob2hEb0YoaXSbS
kWK29SnN1W3caBL4aao9BThRjyD2TP7T+O76yF8c0JPB3+K24rs/VSvoCPhP
hwzxUGJCgMrO/eGSPa8yFGicIvH66HO5QqvhJxzJHX/BISNMCGGYmbBhhgpt
VrCaXYeARTWPKwBMuEKbnV5PV6Y9htITQqUAj8o0ffUHOu076pSQSpLBHp5m
ds/DxYc4ZYsIXF37mDvsMBP3FVOy+HSsqHWrJLI0aW/bRoL6rtwqjnX0zdrw
8gvIrkSwBZh6CqcScB3ojZqFEjf8DkDA5RDoxTdOmvF16LyGNjZTumDekdDP
jsSn6QJ7hnTCYwYrPoZtN2JYk/eYF4jX6ld91YxN3j3LKhL/uMRTVhqzTU/8
AuzEHK+0+TXUkLZhXGn6kAOpSUXIsoxCDhYoDUwrJQGtbOpkNgBGK9yfbwAl
kna9LMX0UeogpDBokV5ZC0zfsz+gJRgRLZR/q+10QpWgydCb7gekkshngUl4
9wZWTp9dHxiUMdG1NNRLmgx2Q3MMPxQRYTwynaX9XzdU9UUFdqd9BaivBLNB
eYVYcGJoacjdVFsi226EDYRFSPwnwEKzts6YNX4gX59tR6O/2F+x1znf3XJo
UU2p/cz6P8y4PG9yqllABouf304UWdwxL8e0qr+h7CRPVEj1MRoVvbKooJO+
LsKSKU8WMck5GvSYS4sbXonsXT/tN6RNSzFuL0Ruobv/hNV8sd7lu2QIhLf2
GEamyim/sNXDLogCM+U186ke/wS6uE+5B10TT+R2lLwINrq4jc/X+AF1ifOP
iEQ2uNi/NjFA2foWaOHVfQ/l0Ym/pWmJ9vcHisnjlxDgQdZqlSvFZWJjPfal
WJuI1gewwW+nnbOUDIQb0pE7M6bqLhvmFO7XBvmE0/mlLfC6I0/aSjqgKkhT
b61QDKI6eC1pCCf9DsgIdwzVp2ui74wuT0qdq2E8isSCUWoEx1Q+MbSQBxm6
FJvTnHP6Ie6cQbeCVc1I/5T8mza9UJuLPx+Sz1MUQUK3DDu37J9TJMbB00hT
ON0YxoxGaJppkm6ew7S5HzlHygA7GEMEqPxCMq2kP/OAsDbRkEKYpGjoJ8Ky
l52Tbhhmdqn/wakdQK05lNHpn8OV2bu3nOV0sbULuxrXAPgxXpX8DcwoGzdp
fxCI4Q4rcNFRfNNUbvx/4s6gUHjOedxbfg0SIzj26pGTw1EBJ6X8lBF9677q
+7V4k0Q7Sq6+36y+xx7VQ3kQz0Hms/YczrLOgt7ZLsWz29dYn4zQCJNkOAXS
g7hriI2jjNGP9D8zeJUcM8Xp9qQq2iN4Qff+688cezzEd5otsg/NJd+8iC1n
fxoUehJpB3q5VjzRR/94q1iBCI6/sdBwNYn6WTi3rtI32gqP93A2mtokGjT2
94hIU31zhVN105jdY+eb637630lhpTEwgoUSdjFMFZGcLTUVcwTo7rZGyE9/
lvS1nNK9F/1Iimvvq1dB6X+RL88Tma8jBIc0pAWbCwrx4Ne1c5pNksZIWuk5
cHFevop82Mjb6Nxgcd08pVjLIXEopjpmxcEe+h0x4qACTsSJP2rrzThfHLqD
Ojv7uRjKGw3rUcyqG0Ikc0oJqeF4gcm07Lv/GR7W7+F68TtjA072ApyksgRk
wKX/4Fg8qbNcc2l9S4Dl+wAFVuxI/Sk45LBH0GXxBOh7bjC3rdvGWVsC9iDs
HWKChDV1KAicLZ9cl8FKVs8GLPU/smoayQOsGGluZ87xanz6xBWW06hCrdUd
GSf4bRF7Oder/oOauFZ7vaK6AGr5VOyqLoXic0MY7zeqbuJZopl0cYzipMfk
cnkSysv3LBsSz0V30WGop3PM50baWxWwNksOqSwMGw/pJ+uFFdoo4/DeOX7q
dXDgXKMETBh84M/L7gzjhlR0El732VngzUgFm9OP72IYtCfhI7petpfN6nCe
dKpdhoE6JY31BTk7Ap8Rk5rAo0u82EtWcljobOwxBQyfgYF5G/25EqN6Voif
ppvwCA2YhuuU6qlMFvqYEmgIxX061Gyv0WkU6Us83fSRkgUNf4msaZuY79M0
FMdRK+aELJAHW6IZOqXGmsUy8VNlkP6cUkRwG7FsMSGAYbuIdlOHJEx+1WJJ
WFSPyaO/xMrgsl2Zpv6tbBru66qUxuae/77gNuncq7cykOgesX16gTAKzvTF
WwU09VofKHMdd3teADmvpQlA+g1lMBwtBXbXZnxcg1flR0SJy8s96Fb260wE
yqr2/mxBnikDvLxX5mPjhdxRaB0jW9n5XwEKQ7wceCdZ/JxvG4lWOtPryXW7
FTuN+pUM3mUcBZlxASDfbZB6ZmzrexQXngHeU9tg+YVSS92Xmw5MvUjOvYq0
4s7zN1FAWpOf1xjZ8Cdp3VYuDGBoCHCILlUPD2v+YP3+t68i275h+0+sBeW+
GIY5a/08AVNrl4b8Qeyrz/BQUIly1ZC3wGfMnqG1l1z82DPXxnsPbtZdoS2z
IKvmo0sJ5mNyz//9XxvkHC8GxsrZHLpZPdpvlsqWic5RYce8iFCQenSrJg0H
F+AbHLVbKzPsDmo+kgMKRy3BKa3qtDg8aeOvibjAcvrQnqJ/AXgKXtLifDED
jSIKZ90YFjRXb44dw/qcJTKat9/pAXEA4trcfg7X3JlNPWXGp+unI9NhlmLd
Uhhh8IY7rnnGUmuKfciigsp5xH1dbnw3rQEUs01+CsLny3Wkx59/D2ZLMZH+
IUHz4oRO1eoJB8DOKS3NKAlgacgFfegTcmkxqiSfBHhtm7QDkt6hqlSvmgkl
F8ZU8TirzkusVe5G5Q3xTW1bi+pxYHW4OHoxQZXjiY/XTDMUNJ3iyN2UFlrc
hneTJSU1SayRKPxH2KyaE7G/Sp1ttPXvpSNZCvDlrJJfE4t0CsuX11FPzAYN
DKtTahVAi9aSbhxMF0xwjLul3Ak9tUH3XYRDCJhdZz8bi/tQsLEKuoiC0MXT
qfRErgdILwjgu02vhFMClwfwc4ZXQMR50wAwHJ50NYYXpcUpPk5Te9zmVR5m
9/h72h4Gn0k7GN0eclbmxRisRdrdsLLfsRPxWKLEX9Iq6Gh24jHOL8gm21aH
TA7AA8yZwscWO+C9GT11FzKyVf9G1tB2IskIFAzyic68PIdC+QNkcyi4PXND
Px8uFy2Sz5eHfVPVlBMP43ghqjRdf5wvQMxqImG119TsTZYXXiv0NYXFZBo9
34VoCX0iVkrD08MHgoTDZK6wJJnl7Um2cdPhOb9beqEi4+W7+5lpme9KJ/91
ejpBx7vSdDGOX2cupPgorr7M83ZiPRBO3/aoFnHW8x/dHdmw1g0puzpletaX
Ljphx0gRms5z3Sz+JKmUD3bc0kgrfY2CXD4+772Ujlnoq8sp9hYhpsLjrnTT
gLCwbx0xEnNq1eS/JNvBLbX0o7oapIKYyYwySkWWAW4Xl1j4Xkikywlf0XQJ
239xjcWPy4mon+aMCkJlof+wMKEql6a/neCbWeZV7mwjaur1mmfh6HoOAj0F
LDi522jw254nYZQLX+E1PUo1X0ACeENfQi0f3AmN3tp28uoY42KVOQ9fPZ8q
9nfK3x8a+51oveNeJb94i9mdZfM9q8PNjBRf17801uAEO42Uvkbfa2veqmNQ
kIPXqbn1BZT67GI32agdkukZgZ0STm7aiAx2ipmMtTNiw254R/pLF6ZM92Gy
cWz58vljmpFtaTSzOPbL05vRzZvrvVSid1TpnsKd41Sak56u4IIMDL+372aK
jC+Ijn9JlRHJvhH2QytTxM+MWBzIMia+ozUUOMow9e7neXfaIJgbzEykpX/0
mT+L6OkhGNTJJqvqJxYDFlnDHb2d/cDX+CTeFJEG2INKJ8N1gShgcQQkvbeY
lxcX1j7ulfUaeTR8HKjavJU56itxGNBwOx8bzX58X9rPSwOMdf4s8Is0wBuj
ZJv+FhV37QSiVd+thR8i7VQQwdmvxS5hoOlQw7btsy6hNB3zPb0PA2zW9cXx
rvIqsJmTsAJa/eGnR+2ubq1vCXJ1AR/iGybXHoiuPm368gMLzwvJrcbi8Kw0
CqGms3+RxAQCMLPj4VG5/TEDqZnrP4r6+KANCg+JPRFYc9BJ5q+ARpqKPeKQ
eWR7eeU1u+ed5kxtDmjgpkJ0BoraTm+AuLFEbkyDA01hB9Otd3B+RGIhtoSn
9vh4m3sIrPXw0a1QUoAKAkd30Wkl92HJugboZXsUs/BrLBsHq172Fid0fEjk
ZDR0YqSCIi2SzWi+5zej1DKlL6gNMqVnnLErReXCLEyUAwG6uCkpYZ6kuuLe
Ha2U778TcgNZTryG84ZYPlNi6mtvbft9UIUGDI577bMBN2ws9g83EGwrSsFS
hR8vAjTiBrxj34s5AJ4VJE9qJkAEAFBY8aPEzkYclvg67CZv6iOFSwcE9aC6
vDp94P8Mb1Jwo9JyDbdN5zO3a8TEmb953VjiiMRpi0sTwQww5LHNK60jR4DQ
r66SE5qkAOlon4qQ8+60wPwvVBTNn8sv8T2GFA2t73mey9VTrA9k9r+47VOr
VZxlL/bDCCMi4w5gBlyTK43EuYO9PnUAsbM7P7DAFROWBw6syB02YIDbj1pq
1wHOVGglNTb5oDCns4Wj2dXGjULzcN8Un4SSZXPcH+F3UXQdyH52x2rkcBip
Qr/UKjHtywNrABrES0yx3VLD1M1ruYOz4CgITp/r/D3Avkftoef7SN5yPF5k
3/O2wxxZyuHlOpGHOQxogk4XNsD3f/0JFrTja+QWWdGYR0S01cNvK+nbWZ8q
hsvbWRXUZGM5S5e4rOW2szNknuJK4b4KKfkRt2Qj3K3hsdJDrCwG99Di8i6d
BDJvwkhNFmNM7Ywgpyf/CgpVUG50Ef6PQsS09IvWsig9hqq0jnOs4/DzHlkh
Jn6gfB7hm0og1jBmutm6pY0iYTCdPjXSxJjtyvlUiWi+uXiJhQ9yER3ccfNi
ldkprwCKn8hFckST9bc+Y+CesYI9hDQFv/3iuSVaR/oihOGxLLwbMK0C99DY
l1NDdDI9k1L50wssTqz2gvIYzsQ1hdWn1OtLxeb5LeGnfVLAM1ZmUMmsFxYQ
/IIQGzukKuBfttsmIm83efZnRSTH7RNV/VOiyvuGQ7Jx+4eZVkATMK567QhA
MAQLSYjnbPkE9jN43qZ1tmI5kz9VBPP5kI3cOSfP5pNPRqiOTr85k6YN74IF
7mbrolaGsIaRS8MYUEySMxWcF1+KSO9p5+B8LuI3+VdEpXLb+UHMCYExHi3u
zO5fNzAE1llRFmV2WSSlX3Dkt505eNgSZ7xhjUePNcFEevxTZcQOXHDZWBOS
MzqkGXV2SwCxYjVCDdDdfLJFaIZ8vrgP2g/2l5oV8exFelo9v/SgndAe8qZi
ZTeHnSi7sHt4WV+QUhmubVrAsKwSe/l8dNFr7EDm2Mu12+8PHvhpINg08KUg
efIETcCVuv+pfRjTCbg3YPaJ76D/6jSci3hdrkjr3o3/BvecSsySrA412QHd
1DYws7Ou3qZAPgekUWQAKvYhjRss3UcSyYg4A4o1LNwRojjNqe292jr+LXLh
NtAb+DZTw5hgBYcX/r+4SOf3xRlQQawY3vuQVDpIx0P1YsNkUlw8/OeeCugT
jxPoGHcQQHRTP4IxZCwHM/HWq739HQziTYLNCgb6WV6+EeFMH7VKk+k/YotJ
IpjB/WvOoRf4AQaRNapgWxi1w/gzKJshBOIiH7Jnk+pUPyr7iTdJOKneZ8Ry
fX1E5F9EaAUhvVvKv4xFNoyDqjq3Pm+JsRprSl+PJOLzXnZ/I8jqSbeXl0bG
8sLiOsB19xqLIKDx3RIHK5g/jRVeUr+u6rlzuhQNrasJ2c6GCXPKal4H1NiU
+1RGXXbaZ4t1WnZC72gVYuDtfCj62wKoHVZz2QcMU0kkq3ziGQQ8qNLAwxCl
POJVOT5gFClLbZJUx3oZhzJE7H0le2eRpsvl0JUciRYdWoHXOoflpxqmDOAD
fwxhEBcWcbqwtRx79SST4lDtqImpw/y9aPKms66BeRaNhvxZUmV/mOAbZ0Jt
4Wg1xM1LfN9vHoECZT+nv7PO79qYfO3Y6LXTjQrYSjjSC9Pge4BlhUppVpHj
Lw1gogiQPgpWnnCK60N5KcAnOD7UL1r4V4yfq1DqmS87WzJPdpTbNpLmfq52
vl1QOKAENCpRl6g+4chSfNWOdPyxVm1FjNSwX0IydtDaLDjKX5kyedpJCt1m
mUKPZa+Cwer9DWROlkXpySps8nUhSABj5ebl7jAGoNxGGg6riPIXjDLr6g/h
EaOdvDyHH70w/qXTnm6wN8fOLIBRRoN30KR735+ufpIyqjAcIbA+XbXTZQam
X9NNE1w5xDRzeKM6jIxJxd6hcAFvBpAJEYH+F8XA4bZPrR9T8y48G4p2SeCO
d/+6rdjQm/snPCEHsDuRpMOmpn4/+5NL+nbvcpBYNT4t0kmb14EzxOlUwguK
O8MRsykEViVGLabreoQCnNUklwH7jgbLVSrEk0XFcGi8Zk5R2ZmjWgiVc3PI
bGrrkn+U79IRAPalfZg0OQE5OwV4WeaeHp/ptkQDUV+tWr/x56LSfopotXzo
NmZPJVP8wYblOyRcFnuXcAhSDhY3lozgCGYpz+WGdOMiTgYiZtI5vu5S8pH3
Qa7B82zin+bfeWJJiA1bzKGV/1mEi61r5b9IkHpXadIMiIEZD9c/qmcT0iuD
GcaejINdgrI0p24H61v2HpCvH7COxIMgCIwOgyrevjQBJR6Od+7iQnus6bPa
dr9UB834eddREteXPYjOGClxZOuz7zloaHA96L+4tWpO6F7JTwnNA3/IIwIo
Q6l9V2RxHqlW3AWZJsrbHtQSzJfzZGt7sesBme5o2QPaY0iJZdyms7ItmM6G
IUNtpEf/oPMyRRJyO0MJKymCsvVScQ3OPxFsCokMKupb5wHQSrBnUfpun6ZK
M9cOBOtd78oMjqDkssx6Pwejtwacj8sXPNPg57r+nLgU/xDwyfOTkgSGKLId
9G3QGe+1ynBurcfPHNK8QuZ7tHWzwmDr7lSVVDtc0AKIBtTeYrn1Dh77hgaF
CIdeGCMO5PzphgNwNLVNIq7R31sYF74L/nNQQPZ7hgey+pd6Q6+FfV1mNQxP
JgWqXksfuS3haxOc52RzHjbihCyJ58ZXS1QeIwMA4p3m6SEEF+vkFRWmQdiG
vHmejmRMAnwWcCU0PNfUx6HTcERHg07plFDDtZIqnILzjrNVVi1GnOcPWwpv
VEz+sZpIFkIdtfTKG5lYJWzyCsou8fhkA5pHilZj9v1F9+eDfLMmla0FiOBC
HRVlryJ88G98ApA+deT+krG0iLfNacXjJDh44zlOVSTRKRAXCR+f4b390e6r
zCfypv05WLWcKAMAgvBzi5uWEsixwCXESEvlLHpH6Z3N73j5gZndFxnMjPmg
OisMwne+ZfntuxUWgUlNdG6t4m2azYs2vA8lC+GFNqV8GXPpr/ZnID2qQpm7
k720HlaItjZ2gKIwKXHb2w+nzadjEfoyF9gpPqwF0ZgbK7ZoEb1+MWToYw7S
21fZ6gPjS8GtAtNle92obZM/NH69cvJSuX7UWpxGFcJo3HZyaVWsLwAxwd7/
cioLZYoL+QE+Fn3w8d4zva4pVW++nuaRTM7Vo2auOl8Xl10R/hf6rvJIJB2x
OETCV6im6tVID6rjSUUVp7/NvHCR8wk8KH5bnMZBMDosN+28zTzcTfmcW8qJ
iQqCTNx+DbWfOJf/1FcfFhQvtLhCvj+3KPE9mxRpNvMzFeU78fcVisCe74+x
HWjrZVlb0Fr/9ECqVa0sODsUSUubP5N7xBLLwEXFY4b28zyldJVKyORtNIpn
lcSdWZogxVSDxNcJGCIO7BdnscHxBq0jYskUie357EPDmOPGmkWBvz4wMxhK
K0bO4jg+RJ67ycmYm7/VRv7qZ+riwDTdp3Twj04Os/aoAYFI+0OZgJsieuvm
YMnBhuF6663Or+iXr4t7sJuWSk2HFcmzAIhIjlbex1GQIIUxUvPErD5tKo1h
76vUx/Ygi3/iG5X94UClHeY1t62cvosUOV8V3O5tDeMzzJUzkkWc5dGWGDFT
KfXS3KSS8WtC95/F/+DEC1Pi0TawaUGdljYP8CRXCmVCyfOTNg/+f1Q/BuUi
wY5bWP1BfAdsz9rsS1UYHb+EqucNX4osLq8xt8fAehrnrGPWE0qzQ9yTGDHn
kamN1sT+TxA6V+TPc1/SmImMYgS6QAg1dbPbNXX5WJMqcfkijeVmcK9o5GC9
emvzbWfMWQBNzqicU7439sVK69IAUQPJTFfCPFULs13uz/AEdMMphQdhL+T5
kXXddi0g6TlyR4Ri3OkpQSif7IPxZuKd4WrruJVfGcnTbLfMUsN7d3KSQoz0
098jlYioAhg/pnS74FWuCfzh4nHQWYxQuz7y9/P7oD9YRE0Et+Yae6daSSkR
HRmhzsHXaMuHqws6HbFDlS6ezGRke3pU0ZlwhgdtyscuQW3HJ8uR90kqBgEE
Kso0Ckd0TVyxWsUc7zRnOiEIJt2yR5qZz7YiwE/2q6XUsUpsCQzt+4EyAqHJ
RaPSImb77yLubLaM4ywR9FFLsQg6Tw9cZ09ndrXilTWTNbL8rsKzgtu9V5Wh
E4c/KV07W7acmsY3X+1v3Kh4XqWIAdWmmDPppLbaVFx9Yk9q3LSJ7+RDQYGO
wGBFFTyBdaVEKx1WYtua6xcnY8da9eqsGpFIBkzs7QIZ5vh08s3LwsuOWCPc
EmGY3+3JDusRhCDep4OVJvBoxBw2i8Qy5pvfCIB/Qg71jyzXs9OuIRG6Rb/d
bBi7Bmjble6ihct6XJsaHv06XxsTqx8gHz4DlcNwgPKSUCwqL5/XqSUWVyW6
sPdfsaQx9Yj6jX9Wb1up6oAoO+PtKc1Sp5fh1YA2MdbkDyz8sBre1pnp0frY
kpOeaTs7Wfpb5SWZIJFuIXhetgbBp1wcVKjJ8W/u6cpgAcUIwPWPjQX+hSRa
lThu7zZZwylMGvL3Q4EJqzydywq5E0cPwF8sDw/IQUpgfttX2CuJiSRRQFkH
fhMTUiy+5nncZovz6DpL89pOl8R9nwpg0WMCBFmtq6C7z0OQrA8/jj1J/60w
W/kaqGXjdE7bcsJePZ+2S69NbYHXbh7x9NehPwcP4R4gaVBI5qcsMN6Id3m8
kgLwtJXy9gKdzo1HxVqGI4nlur/Ax+1HtcJ7LBa9p8Y1J2VwjvnvfT7f7LqN
e5YXD1Ld0PzGEG/7j/zaLc5gbZ6Nxusftw1J21r+p8bsNnr1069UevQlAmV5
r+3y2FutcFKL2mXWQgERiq7OlYi74JuzqEswP2KgTvQO/Q20jdC3nReM0TJL
Q9csTWbdlYPkV6G109wHbVWnStnVDnulirwPBrKjzBAmXl1ypANnBpoRtXGv
xPrC53jZbsvLmHqwDgXi90b6oHziHXKisPxP/Gm7UmmKC3TH1qa8kglYX+BB
U6w3AhzpMPBErlvqochHQn4696fMisCRSCZZKspc8OcrhRF3fFQQG5DjtfHW
88nqythqGtnpLU052vSHwkNmK5p/itTCuk49j3fir2x5QbYVPl8xzouW1Z2A
g1m8ifn1wyk0wkjfZsBuNhC7GCfWifQ7hmAgkQ6YhBoJPCGAadx3YXLjODzW
AGPM/TIlNvjalvBgnpX/u2M0lskzpGyWB8afrMTRj3TaX3YzMUF0CGgUAKvk
NVQsuSUjB5pDYUhZM923Iww9Zhx0vTK/MGYCyw3rojmgtOgJRcE0Pq+w7eMV
XUCHLJ0oPRu3GC9r6K9eBwMU2sW/bWssDwohytXtqSuk9giioX62Rn59ZJNS
SXsu1r6MoVg14jgqSoDZktLZV0Q2wYUOGV4nFDGIG2KJLImfLDvE3Cj6u8ve
FQ8Vdi/pzBMSekeO0zNx6BgP7Nn8ecYcg9Z4u8AAX5jPwD6jTvZVV7gqbL6X
55xYEF+2NYOSzNtspGt9ChwHoBV2j909VjyyHys80bY/sGCBkLf4eZLJxby3
/hFRlJrH38W1BbTkHviWoEKNDFyZfrkT2U5/Uggulf80ve/5g+MgpE7OR6Ow
wGHQY/7QtwgoTTyMBxzn86SAeWOw+unhTcfuwdJa/krjX6S3oJBn052i1Z9r
LowQulA/k7e+KnpFlZ8uv5t1l0JNSHf6vzFVJ2V2u25h0xiZOSLUTefkZibZ
oo40JFfUbvZ7+f+6m8XWD4PKLXqdjbSVK7W9UDB7tYpbYYE6+RqQ06G/o/9F
7P2mre5yf3w1tr8dSYMkd00EvaVa2qmA2MFdbJgLhoSGUeV+gB1bA5Un5sfP
osEh4yKTj9JqVxBzswuFCwrc+BoU6YHptIiINd6H294BHpOEHWPUIsgXc9nY
ts/bjbX92NjW0qp5vYv6dxy0SPvxWUNpQMVFbDwvIwLxTrj909CdWQWawRM3
6aZhxbK+YwL3L91CU078GCv2MxzfKSQ3fMc7mqmVd/lTJABlM75TNmjGjgba
TSnU8r+AiFul7DM0csegt50FdqqBWznHboTH8es507OFsSJ/QppUFekX3Tqp
U25sCyWXDO18ScuqrOE7nM8tmML4XPEaWcZxLSdrt2qZ3PmK/TF01/Ylel3A
NjoKi6BJMVGcRMPehSHfaSNzhaJ6Armc0P8pUDjjwo/WLPCCRPRBUltOFVTJ
es7FaMGcVTpcqbdPyZgSRjpkN9oLCqZXqsefcvpqyISSOJ5IlzOBGHyHysHk
r9n3OggvdYvrSDLvDWtO29FbtMK9K51l0pfREBsOqVEWkTBlqQDo84cdH7pR
BJZRE0ppnQ4U5+BMbsjynSjPZPRjC9/icnAu5BDWKBl7pBaZ1OQwq35z4mmy
hx/WwMWYKtna55e4YMHxtBR4+s7OuvIGjhf/d9szSvSTxHR9I5Kp402N1j1q
UvnMGNliJcos9/Oa+gdf5T0i6xpr5ALlGbAHQZKuNwWwOon8kSQatim7tyIr
AbAayQ0KuC7k7P9rusiANnvVK6r9Pqjgn5gfcUlKyZuTlHRl//X3SsplrMwU
sNpPsnIM4WOiNnShkZSd6U7pbz2IDUI3Bt7v8ryIPTVGOdL7UcAsN5whN1Qe
eGnauhd7y1qVXiFLQFCmb+4IHkDqcyG6CHcpQGGHxYSuyGyaS2rw4i0rGm0F
5PzYhayiNtkSqPPTIp1cIp0MbLfrPGCEoFoG+KoR/fv41W9UFbtQYvFvgF5q
as5+JvtKRbkrU+QQCkq9Pikd/c+/UTqnvRisVMosLqEXYqUISSxAah0xop2h
JVYVHKg6BWedYBQlpv7PYbMHCyl7HOPNo3R3ex0zyqE5Vq0HwkhsM/vq7s9r
0zXCKHrmOrTXlKMzJCqTOK/qfox+Js/nXIOpD+pp3HmGn0Mhu4esTL3rC/BD
KK5dvhlWwcdKBWA4h0cOypTN8FxwJPMsi4pMkPboednW5PsrYr9A4RsPW87D
VNPUisxF1UC7fSVwbU/5gbZzeMfJY9IVMexqYZ2iClSVH7OJbpTAf100i//S
W5/8LYfVIQtClw2CzTr/tSXPTVcR0w66Hh1lisLXkQ+wzwGw2dVUxv5Ff1qN
KP1s9n9PzHwvRMnBErJ2bmcE3iX6G0EtpGOCKieZ7dQYMxWkHvjXxKBYVkTV
lpst0eCfMSTgZrAnwwgeo4a7Z2di7C5zo8S2JKOr0/KQkcYm8xNnBBxk6453
+0tOvCejCZqj0uEwaKV/IT34qaod8VyyUIR1ERsC7aUKD6m+HPV1EYQt0Qsm
zqU3tgS+md6Cose51zovOpnHnaD2j5MOPLxkyYteFtUdP5RsyvG5z/sbec50
BP/CKSvBbe7EDCR1P8y3LSaoq4Yu6h86PW8JlHElGmps9bOxeTZqymidzueF
ZPogAo467pfcl2mhDsp5n9w0al8nQGjqJl1OKI1Z6y9MXojO4aXaASKntq3d
CPLTpE9dzWhtrgSeYW66LvzZEKDC+3fPetjZRPrHfYb40I/WrBhLLVKsEDLp
5uDXnGNYZSWCmKQf4lvzq9rUk/Ilv41t9vWhQGUmEOsMORFVv1WEubhg10T6
D44gi0jOLg2D9iPt8cWbJKBdPcb9dGJVDa/ZdA68RjOERukSz5hsEMt3nq+8
jGTN6AwTV+XvzjkqA2/vmk0WCPIQm3MbjSUVczyHE9I6+JzipuhINGqW7Gp5
EXl92ZuvA5LgmFu+a2IX7dvxEEPHzI+f2oDfFAn94D3m8QHwN5OrHISAc/4R
ug2pl6TlmTLvtBueGFnIFYb4RDn1RVykSStWJlbiDEENluwCfkMyz4NGBzg7
/oO5WUdm+Ioyt8/nkQUegtV9v8ToxKCYuYJYDeisbpHOiSf1uZSW5X39bu4e
G29L7/7kdFkPjHObkYj0RpruvQQZ7yGmHZJ+Gkn8p9H2C4e5FneMldmIx7Dc
KKAyTGCTujU2zOmgNW+uD5MJ19EgOaSFjR4yAE/5xYagsCm0nI6x8ja3Yyxx
1XNoVrRRYNQg9S67S4VSkec/6nGYAJlmUNSx1B0waCMjIQcxpAUVNVrG1OX5
B27/OXlONFYvJPtEKgpExmOYG+FuJGyXm/bt2CCnzEswnTjwaNrsYeEbRfqJ
n8RkGUPx6LUm0Cd7b0CVS2nYOYN4NxjjQ4yyIl8MaHpkeL1J+Pu4SC5ZGOUt
ayqCjCLnx+FWrSARHHkSBsrsD4oWwW1pd5I/0y0bd1kPw5loP0qZ78v5NqKJ
PRm77uSf/yCPbHVBOde5QU4JgMg6VloP0wI2rKamrp0zXtDSlkUnzO2rnRj0
Ku5cqVzawpC1zDChjNeVnPcXvreguhURHWTrHUSA+1VjN4cKKhwLL48aXUKx
CtDFOhL4i9zP7kkFffftkarcl0lRS5tUmUO1iyPljTcgjBtIirT8Q3NiYwoy
WJHlMOVtkh948p4ymKMdSRyvJq9mslkyIyaKuMJuv7NfnWaB92XffnRMamLV
9poYAMqL4VWrlW0Z9FQyThLQnEgNenAl9tpueVQKQQqYfVnLBkIjtCS8xUrg
sSNC8kfBTvF6C46iRxTT62ja9cEvPGm1ATnA3lV0ptKCnfYMxdoJgM7wOvOx
Qhc4SXPciEwI29JIXu9oDvdDcopu+IEL5ficHXp+Et4IQ1VdviNoP59MT9Yb
ow7flhE+x7AGCal9dwBwrsEM0CD6EpaO+7kUluH18zjjrWaC9Gwq05mWqMic
nOZvHYXpatHX7qO1IgFLCeUSnwqqPxmiayIBmsj4BsNc5ldeUIQ60be7fO6q
OXJr1vJQZd4DlGcMod4/K+ljLKW31aXs2ZGgjpuOc1DhBmK9YxxdJppuY570
qI60DEAMFbriD45IPrmsqoxamxJ+zRwqSMhRmT2rJvIMWYm3eOkiwVf4k/3C
7/2XvfCnohB4+tIbuD0sBbRNgjYhms5OvC5XFIGss8CkbFZHNdrtgda2bqiC
0Xesi23qQppDsJ81yT4hhKY2lQ+F73F4eO1/y0yFBerJHdtdqIsnID+2/qO0
kkVhJg0vFgdwfmIj1Ak8qJoqLNWOAD98QVa6jBS5u91ECEMgTcpI2rwNpBKI
EMQriWNn8OkWuOztRacW7Scra18w3u8h7To7zpPE9Q5rx1iLA89VY76B4iJ9
HX3887luK8lfwETHXXaIqKCJDILMNA2YpdxvdUO/XjJnH3EMtoSVcx+yQdY3
7oqWmUOvjc5os5FvcpHIiTRXnbZdEPSH/AF04krc9SvZ/sajxY1IfEOUA1aT
P/UYe/vkzdMYYWShpQDUQcUz0/FNhkxWa1BcXSBxkPOt+M9XGE/Q/9FBmDof
tBpOmXBQKxmyzGxWhTLmJRBZjFqujYc17C3v1TDx1rEbLeJMPxyAcixqmkJy
39G/kXNOvA6Mmb5gpT7FD2Ezi+orhy/wCfrPqB5OKVcCZqUCbr3/uCzHdr9v
uMNh9tCQwoaBabTcQd3bmhbVooYr3Eld2NTefxT9bcymTXhBXuxNl8UIMUr4
eNihn7a+zyxUrb7QqXq6yMBFPcD6JBVWXeoW7BPr8Ma9M4LwP+1+ogz3A6RQ
kVR4LwrvlIPM27tX+zte937abtR8kAxeX5jRZFDL9U3cTiAFM/XcyCN2tgFM
YjBaoqpTI3XshqWEajGcVsyju6VvvujVBqW6Xx+U49xbt8vmivtxybWM5bWN
rba3Ddj8RVMK6rJkRCBY1ExZq6sieHCglNVItAyLm9bSA7JSXt0qXbVCD2hc
rWttJd0LEmsMfaLBD2lijrBUA2fUhRgmxlzDwCJpZNR32BwQgqBVFVyj+VLI
7DVBJINwZ0PZo7b54ZvksQqdUPqyklrqntkFTvrSUg4UkSIMDsFJiJPm4CLL
EjF/7HxXjy1HbBOB1fTgTI+6E/g/hg8kx3cO4G+4ubCc3TzeG0Eiii5gNq1d
CCFGAjJKlfJHMuQ31SVl4KoGZ3m7RM3z/BRKQwc0/47Gi5kST+7or/nemgDm
1iF+RWhcz+9JzRsTPej2Br9HYbYrFJrAZvvXEEd37MG6dZITXLlPwzJx6jMq
nfpn2ng1eI2UvifscJ7z2hwQGp0DgslWPQu1SsUteIzf/nXMSyeVSDSDTjP7
E5TMXUNmllRBM2fNT0OzaFRmj3IqWysCuSXT/g/veOTlsLKNk34rugbfyPJn
43NLcaWUoYciZXgmB96Kn4WehaNNhyu918J3sFpb/xhsWJo7VtiP4j1XsWgz
CY8/JkZG+nGHBl8/VVm5OZLrzV7JydXrD5D0RSEaGVFUH144SyA6e8xXFakh
U5mEgaR4tK2FlSHZ2KumbIM5O+2q3jkvTeIC5AKHwBg2VgJ4kkm6V/MQ2YJa
J2NvgWEC2dpD1OKvbvSh5Tm3s4XjwpxxDi/EQCWnNLhJNHauEJA9dLFuFJd/
I/AOBolzledmfTz8xoaFAn/ZeVqm4queWsU3Jcu9mdey00/m0nDrQLY3iVA9
q5/KWpXcRMnxpxcJv7chPM0vtteI1b67Hl2NUCb9JSfNs0rjX0F+sHMBi42y
6AynIhvb9OBaKkK9Fm6ULNVZF/FbngZ6s3+YUqn61G57FQW53UzwuK5pJeZb
gcwg/dWHMlwHa3jsS8JMOlxFA75z18/5qkrXwYFdmbC2EzhzE6/GaDK3QmFW
epW3eBUHfCNGh6GOCnpK2Ke7rSiLLQInzPZ4iw0JZ/ZCA24fH5KhOzqAq176
ZufenQPj6vaHewwxEpUGtT1u1EV/JGWumpG9ojlwNVJ6Mwo1n3ohvl/LV5BP
mkwldhWLj+FHqo3klz5MYaeVZHBFTjTMxFKWTwxOnNx64+3YNM2DccXuaPIE
h3/sTZQDOhLSQNGAjbCkiIlUc9GzPi7q3KhMs9BNIOtL2IhT54Rn96TvfvVh
g0e/Jq6nqiZlziB0K59iZsugpy/81OfsS0IhEYdq3lqm9xR18IDW07uQDoqv
EiZ8InHFtebHhfiton4i5pYZQ+KktmbqL8us2o30m18Wbvw2IqACcb/R6Whz
P301WyDZP672KeQtuPbIJ8KgHgIUHB9wwr9b+fPpddt1arI2AAYSuAz7zv+Z
rbDXXN0Y9mwBrlERH1dzUY5cP80ma1QIk8Zp7tsi88v/qq1KKnWLDz4Bz26N
M+VHMnuwe2V5Nixnpywz/TFkchP/QLxpFjgiGShKmKZO7mHlR2EDwL3KBxux
9051YCu3EL7QnnuK/Ui7v1O8G4yaE4kfOc03nnZHz9Mq8d08ZLqjNoXOXWag
IIwQIBUtug/XXqU1a4MYd8oAsiS2xMcaC4H3O0pOoxnDCeE5ebBSxaHkLS6C
p+S1dXFuoRFUec6Zmgs0y/9W0ClSEtzSsYJ0kXfxw1mx8qGBR1uxytcGeeLh
8yqS95o6rONc/tUn5Xg2tIwKYkIL0o/Q4/LxA+mrHyyt5C/OhFJTaAFsPLh6
o0IIM/IdZyCWNZLPQPbvIzrqAHs+KWbYsuBvvWBIAREWYbkFSSjqqLK3yUi9
bUWZujUxyh4sb+OtsE8XKMA9MDF8s8YmJYYFIuA4UwdmRtGFSYWD4RXEilZG
EFjQZ80Fc7b14SIb8ClgZbQftN1kyY2knBUissAgO4s8Xs3337MjLbeOF3e7
701haNwLf7uWeKpJJiG5JP+lOQdE+adSeKXALxPZYfPGvgFJ+LMQzcDFw9Sl
SLzNJyvsWDfE8n9pTxUfRsTISxAWR3Y00jG3mrMCphqrfVxrgVXjgLbjxAmy
OF+Vy/H15g4KSD7JLkO1ZYRMZ8S8uAYnN6ES4gEDhj7sbREixk7R2OoHI/tz
Yw20Fgf1PPycc3I3Ut6/zWkQsdb7NYqgx0AWD8JAIoRAIEeFBaiFkXKj7/JZ
VOdKTAd2bcFCZPagMkikLrYDzctKdLlLWw87W4f/+wlNfwsuhpr1fsGq5xxh
qM8cbESTK6Vl/v+8dnu5rPsuBuGPJhVYi8XxkifdmOu8XduBcyGG239H4I/f
q4p19v3UEzbpQ0RmQo0ZzNk92CQi3WYjdYfXQSlYsVt3RaTBIZ+PpXqd7ncq
qqp+viYBMaOeZ92K6gL8I6y/52vaL4pT3H3qbx8M9WjlfdWkYmN0ukShVcdK
0pwRss5E1x82UB7KecsKENRB4R97GK5agwVg1wVZOLJ6ky1pEVgGFP2RhNiI
6QWgau3tfvdRfC6U8CwzyiL4QM+wZb1tLUy377RpxMDygYfdrVYN74kyKB7+
eMX/IlW8KHGaBQQ+00i44jpepLaOK+OUqYssR02OMPBTb7Ft7xloEUNVxmB0
C7Ryw4EaNdW0iUqbiSPSS3tgWvnXwfiuE5hROcBUO/tivixcP0x/Omna4/Tc
03l1LvVmPfly0AOxfYS/j4TgRsVoFckYWO8MGAWeWl/UfV/9C77Rr0T1kwPO
ITHj1Bxj7I7cFx+znrHo3eNHgn2phD9x7TX5ldRRfvn4yzBg7K3+Xwgoz6Xx
JjTpZdJs/YKtWfGtVSGBMomKjVeZoy5l/Cy2lUMmOC5IsZ6vqcuYcEqmtEXK
+TYv9U/h87RGmX68AaoqMzmI1r6DhbJc1SG98uwdxCc5++/7Z2EtlVN1JmVV
10nPDQrAwrzOJ9AJIqTY2H6L/Vdbf6V59jUH6rz6R/NHd9FTTmPrYx8s+7r1
H8HXuLqg8PBJNlHtRgHGD7j0zf2UN+Wo/ReKH/uISmy+bP/5FWqnmd4WFYRe
I6IHqKP2o49f8HMjWjdET2xEE24F5+FDkvzlUWpU8xYAlzzcFQ8I+InDAEDp
SHDeN1TvCFDxyNpfamm6Cg7CXAEyuwJ/HVz8BPuGHX+hOFtGW0tCVrP1YZIz
0FJ9CcmgJ2iTjaHpBVUN6wmG9o8C+T7NLhFjgmM1pPAMgOmsftBS9LENWvYf
wcgo0x7sgFw9fkMTTi5SLlVarvH5KWCJwemj5FJ2x4/28P6z2HCa6TZlsBb1
o/4Iiy/DCYAtLNfm/f3/X5IQFrNDm22+wN7IJ7qm7tChqWC2bNyAE46x8/Yd
illbPIx40++kWU85Ssp8z1GciYUr4/LooD4bRzI+C8F/hI35aBk6SV0vWtJr
0IpvF1BB9DI3WUS8eZmNiOLIHe+0VpjCHArj1X+tPCxK/STTdb3ag+IJxL4M
JjOJlIp6Nu5A0ivtfcQqkfO2r3yIwphUC25gYu9s+++J0mfo7Oe6RuKp31gu
Xw7zAFqlNYtWVgU8fQsoIqOp5JZ3tb3VsfdDMiS67UKAngTlg1SaApFuNhN6
j+7xi5yu7fKMth+9XKPESlfuVWmWLeuyBxvb0kyuF+5dNttHj2FLHbhYnGZq
SU8iOeuaq/++1jnst2CROppzdVZinXnGYFPSAQzARP7F5k53xbiiZqLeeLyM
m9+6GD+sZbucQwBba5lifQD5guxSL9/VIYjIGrRZZgyisR02fbs6MUvM+GGS
3nCsINjGuq65Uy6+ATjrOLclhJYGZUBtBd+giLL9sPhiSNAzXolFhKxQeJGv
Bs11imO8av/H868IPwpBWpvYfAqGdozN9rNWGKjWCf4jSS+XHKuSTtVuYAQl
+wYbr9xA0OVCvN7cs7ZiabBGCiyVWEJUF0D2nNm8dsGWGOjffYNOVEUAn+tj
8idhvpmehcJv7eqwCwYlTibyNjK/ODEh+xcoqyf3gxXTXdClt6Z9lTUWOQvD
X612brnsKTMlsZe6eOaUNPfvcdV7SZnW7A+0968ioam56Ot0G5svKAoLRaa8
cjr3GzOkcLO2VbYDNEIxSx/VQoFqVnOs19SMv0dVHgNm/UQ6uocgJ3OrjLdX
g7+wTWg+yEqJ/h08OOqJoDsTTuOhwfWogLZ2uH356DqEbhOyN5EArBzMuMdv
XkIIJuPpT1k+mD5vFIwMM9x2q/2CfqDTErtdO5DCPn1kuvpgi2OvB/zcp6TY
rSxMre9BHComxuiO/fdeHpOBjF9upd8MYGfI3njEQ2Y5q66Am9MSE78g5iRv
WmcXYrfgpocz2gvjPjzpiHsGVUA/FCW17fdPy4gbpq3C+MG0BQjvP3m26SIa
bRIUUubRYjTAcgcEuxLdt140gZrESaslUo9if8xVISr3Vga3eJdROVE/cgYh
Nwnqs/U34a4CDEgmDcxa1N4Ftx/dOOHuBa3pcFh9gPn3O0/A0WCx1qHzG9rf
R70pRur8sYbZOeMl2sjdHXDSG7xMPO1ua3gnJoPADNEql7lgFW1YTQjFy7yi
r7PL/ffCgCjaeTXrIa+v5VCbGTo9bFbRv4h0pl/kdt1b0Fwny+j1pKIipWBv
83LiREFR1KU+O5MBFL01IkbbTyo0lh3mRSuQvBDBe66ezayMFnab+jqDv/16
X+HN+DxFq/D96C0/XvWr5bpt0bAE+h/pNbN9neB345fq2TqDvNPSQ1IIwewd
L74v0pyLVmLNums5y6ytwpoGfI4rcnCbb872zs80d4/92DOTx5Xi+VxIMoeU
iB9yXynxEXOZQZXnVDJ7AlzVQor2A7JF2RQbyIPWq6IVUNI9tSCAbvH/2Xor
RsTqy4u1UfKEq1dpctnN3PCGDPJUaqaA/S6TH6lRY3m7zuKCg4aOuxPMatNC
oOg1apA1wCcBpPYbx5g5rJvrw4DYXNeSFEwe/zANSfTJl+cf6K6bJOF7UjKO
Dn2+m6LEQ/up/E4uq+S44k+PDebUBbKMWgThBSSmZTNrwJcwZLSfNpdGkc5o
zNPHlkKwKjj7r3CceRJqYUp5lEcTQlcLz1lVWI+JvC1p7gPgE5Ipq7hppx6C
xg9kFbJVwv8nwtiLTgKuNctLO3PFsgX4TX33fbj0mt62fWLAnhY5Vs250sl2
CkPFKAmhfDGyBmS+eqzO+DBde7HUMqg4RcBcb/pn6t50qMHCZl3va0XQ0ku9
7z5ZzKp0kcjQJLJOD9i38OWMsJ8uicuYjW+xwEGPj2viPhttk9Wj0eVteVCS
j/IWwtbSsLmAb1naMP9ylqhNQfRCNaTrAlCA/Zk6V5gWECegugJISddmhp5Q
hMhyKwfq9CP9QuyKjzUwoAkZSZvPIByXO0fJXBI2axYnY4u6wnqiKisLzUdp
RIQKmFYaaB1z74Apc94Zg5e8B2JCtRWGBu7G9M28q/pnv+h1oQa1nASqYKt9
5Fls3mi1xkvv3wQ0B3NIvHmc9hHhoFj8fbsghVbhTkAPN4nk3hP3zYjHjgXK
LtIGDbbzrLgStlA9pu14a4vseJ66p2EV/R/VFuERJZYO4imPYaclSZGuw7JI
EWNqIQ+FLaF45WAedw8QL65Tic5TA7kMeASUJ+MXxqYOex73qIGVfklizrfT
UzA6xZ0qzvlbW4XTPVIf5rTkOzI+NGIi8CrfAddiPWMoV5bXGnx15xSs/GfW
/vof/qVTlrhK/ywtpJ1M8mvDz6zH8DvKjYxnNGLBxDq2K4dzju39VVm0EEu0
2zTSwQ6G25IXae6PfXTPLAWLjVMuNXuBbMAKQH0KFOlPzpbQYzvMNRa5oreg
DT37HK5nEy93EMetnZN1CAtE5ZCGx45G/lfFiLrIek3DXj+mEKV3LvELBogV
DLPGw86F64XhF21yTC4dc4bHWOYyUbLJo5ldE50F/ufOboCdE/nq2efBqqCY
qRYOgoIbaLI+jvqLyODBTr/QGNrj+McLEJ0CNwsqlW0Yzs23I107XoyRq3pX
xGts0MHLkufOUeTY9ODXLV25h8m10A62ZqZCUSZgs/TGgKWRS2Z/5tsumJ3+
LdgNv3AAINd1Lku6RZ6athZ8fHXRLGKspSUuaQ7+pXbZ5HwzSOTK3BUN3nMr
yKFm+1GCceTmE62ygsWTTLpplpSZC3ZbfrYY6DS8cFnfftJnOFJ0q3+EYnvv
vLZjFtWA99sWP7b21VmPykuhjMLR5VuZDYXOP2W50WllSaEWrQirvlZvRtJY
szPLuz4vjs+tj+pJEThbT/Behd5Oly6nINhPFpMQJZJS6u2rTyGG6a/nb8pC
c2pvgYDb9GEEJrit89BGrDubY4UbvHW7wcNPKWSbC9miFBpRRha0IWkpDzj1
geJWefnVc4qyaRMq1zkAk0a1dUWmIoAFe911j8otHWjGUhBaDc9IhghAd3VR
rO1fHQ+hu86GV+vFmKBF9faZy4yM1JPbGF1bJw+92CYzOGSSE3vX5/MnjSRR
onKMlX+2Wsv3U3GI6oJhjUo2iXKOIko5uvKGbchqNPy500xHMEdINP6Yb4B+
V2IXe2BoDeKDUJ4j3w/xSMWjINhAgqK4MUOq+ZgHkiLUk3jYIYMA3ecys7ko
ONxgpNwKakd01NKXy/GQbfj2JaLAx5PL17iPiahUmvEhA0uMYeHf0RwKAhQZ
2vlW1PtzQMYwWZP5unk8xMVSVX4OD1UVnwNRNjqqdI5tpJZ2dAODo8eZlf8S
i2N8CXAslkYwYRSmRLpCGUZ1hG78rstn4+JeOBWJ6L7RZusUSI5QQTuXqmSJ
0jXXtAHjbXZlzXuyW+cmVA06yhaoYHGM7bWBsvZtpwXtxlIY9iPS1Fb/Sy21
IC367gFGx0YGYPAgxDXxXN37fMXJ2KZ3M/UQWTV8Z5HZPILySJjCzbspfFkQ
32EEotJsRmwRihE9Dda2ww2UnH+tUdjpV0YxoAWBJz57cxfVo4aRmlAQ+KnD
IgfN7u6jhFqdLaB5GReN+dVidcdM0n0OZuFDei3uyOcX3p0jonQuL3ONxSTs
itltW2L0zHr+LMZniZLIjJt8Y2btEkUBEX5MwzIbsWSZMDdSRUqGVDywWe1L
5dM5wsmkhZKhFsPTmEnRl4ymg9hbPnGkgp+fYRYOF3jlB4/r11gjV9vDM9Zv
3UkVue8ZYn31B9ior2/U3F/VyODS9sgfwpTryiQdian/OJ9WYezU0IKmFxSM
EDAUt+XOReWGGvx3ZtYhSsJ+8NZ081uVsUaJ1TdEEtZudUH2+dzLdyHNYTpD
fboQ70Q8T7gEwi0mmb7u2aXxrp/m5i/0NF03LipEoJ3W1/I0Ogr77N8dvGr4
DgJyi5+lsCuJb8pkNsq6cDLOXWYLUY0QApYv/MDlIqD9GAXYtkFTcPENJoe0
PpUIi9GgQWzifbJrp0ZRD6NIRRo+W6RLjTryP1Tz5GG5ajlMPsq8Z9WkTEYs
Yj8VA0N2mD3FUlGUBQRYW6sl0zrYpf+dhS5QK3tIOag5myRAKSm14weBOSCt
no4Tk8QFzSTzlzOcCd+oWwOt9ugNpaVf5zQUMIZgVtEJruy7uoVGxbTCIGAF
W2dlpCMYXr5pZOoOrAYn8Up+8aKirI4MIfpsNJHew+yuH+NuSORUodq2KfkD
RRlMEwBNCyDWvO8rWDLoikgSWfca5wEqHgcGESSRdzmfLvhMGSZhj+gZ5FiM
I/4v14muDDEQiS/yZFvBKLSOVg0fTvCJdJ+jZEkP8Nb2ekm209A3hi5AF3Jz
3LmqvJ4Pl5kZxh4+1O9GlUUPeZTPWZfRGjcLM+ZrEcb5dhmqc5kbs2sqUNpL
oqJHvzv+3AggKV9Ja1VnAdjrRS0OZ8NTM4GGGx0TrB0R2xk+So7bwHAIplJw
YLJ8J28bbm3D7p/+UM1Ka+4EG2JGAkDPpIWE+2CWrk6b06NuKUYA6Z11whbH
s6QepbktHvFOiRP9pcvM7gFSs4Uft18tGiJmY5Lgcu9f0hvagzaYb8J8Jqfb
u5ZpRcIIkZp9gRV7p5v+2TEiSSDCtAZqOYhadigT6Yp9EgWiUNgxwkr0eNGJ
nv+LP4rgm0dWXEBZef4HPEh+PPjhEyAiH8+/WEnOux3lM9LQ+eSMY6Om7rlA
Rg3cy4AX6rPGSfXUeeJA/Uqd8ovxH0SohNo4fRcKQtKawu/IV5p4eyHrHipQ
SizPe1nWNh4PFfc7351/g/bQCC3KUbLDcCPd9D3yd7Pqd26wme6KY0Ye3wVt
VCUBeI0b6ED5TXCoZ8AY3txCorh05y+50BVYIRpHqWYOWCjDacGejsCNq7FX
2r7S1iYfeu5kxzY1Er4q+Gc8V4PJFL7R7i4drknPfWEdkjHLetcdv2RyjJRH
NNQ2f/JrMgGqgQqBurnhM5Yh/jrqusk0FZYLsN/gdXxU+oXEcvfmXqqZbMzK
N5dIZ3cr7Zq34+602fmVfOn6Kf9Mcrv5qva0NveGHHdAkfjEhKC4G5jTevsc
RHz/Qmfb1iEkIFY6AYz3yqh5x2NRzuYZRvAm44wEhcj5dQBmiSA9UR90DmGB
RbNeEcgsMXAvmSfK5VU/YCDyDwriqEjFLJqz6xlT4iJCtM/IruZbE3QhmeCq
Q4rNyMe24MPhk2+hkJ8xVI6XGhgedgupk6wIACETZqegm7OSg6em/f31/rFX
icC2HBjEqopiopshQ81ficUaFakUm/dGWbagqJEGriQW7ifCPYuY5tmJ4xJx
ZTuIsnTNoqJbarCbynFTgxAaNrKhPzkzPeAGbVU1LrX38ka5QKj0InCHBW+R
FAc2GbJgeRKuWwwrSp4ANPy3H9fsg9YviViVQhX++SCA+TQQoKwcfoeF7hsS
sD6uflNHCXEAt5AO3SEs3PU+O4LNR+si3/Okpt/w1SiCJfrAl2YxAKwRCixO
gXdL96qE0c6qROQP35Tpoth4WQJkuoRzTUoe5nTUGbxvuaF9PUWvYMSjX/0V
sTcNvpM1uVgLxLlQE8dX6h+KkFzo083Dmp9cZ6L2UWc3jlonxgZQgXiVs5JS
cRNXBsjCtz1M4KD5mwY1BNWfQzV/2PqKOS8dn+hBl/O9RmgIAQoFZ9H+BLmF
rJ8RP1NuCHa0HdnxdrEvpK6/Bf86ait+KVL5z+cB2+1tkE1fYMAwSlVGU4+T
CoOmHMeB0STve/UVYfM7sJkHv8WZWF/rKCjDRJOKO3wogCZ0/4q0DB/KtJt0
zJb2er0neKRoxJuQZLep9LHBLVwdlPNLVvYf53IKEtg8Fb++U1ByPCehty4u
YQbmsY8hrtdWY8zQfeOLxsPQK1gpAilbxa38hT0kogNzlf6PeeOeNgy16AUL
1S94bTKAgHY59m/TaTXGewavVT1mTE5Xd5UXXmngUHMBw6jlCq2C75VHX/HC
dQgr0sEvDpxk3rhcVvTghg0vmA7dzh4Ifk73QS3SXvADV34R6tt2INkdvr/o
90nHSzoxjtRmg1SRJKTbmbyPzpzzIQhupQLAtEHRC5du3aE8TGYkmm2nd8pQ
pLFYe+XrVa0csXwKN+Hp4cArcaiNlEN6SmY03kJdpV6tG4qq4sSktr/zGxEt
7qVq9qLn5Sxculp1kUtrQd4xVDcZfB1j3NHgud2yxmVXXxCTA0R0tqT94TH+
s0hty4PYWoo7EAbNGOUWm5RTOFB25YpfZgIjICQEdmOE7n+hwrZdculPH+AU
GjoRKQXBe7F+zy9qy6N8TnUX/IGslLjBcEYKljvStP7/SO2UOnhpi72o2zlY
agTEeMXlfWtWnPYcmwUoqK4dGVDFD7FPRKobS+NFtIlOYL/6pcJD3/aoPfLa
Dw5+GflmpXmr4TBbTfUul1SLGh19QQJsV37VIxpw1rChgAUonlUzdlLkB2YO
iSJIy4q9xLlDWsyy+vq5srDwpiMPejHY8+0XBpD80nG70i9iPRZGFoBkVZgJ
kZveneBsnyIUPSQYugtyMZVCC1Kj+B2T0u0zROT+TF9/wFfwUcD23RS/7Qgx
+VYP8BhI731f7RwAEHJA6Sl9psGBCzz84zzLd9+exfrA/qDfI56RhruDidcT
vddeu7s1CWKI0CAOZ8i33k0arFKIeVGNlZ+/jQq4W6kDOYBXz+jIjze2zXaZ
B8IAZbggFz+fE8nlLvW0g1DojlOh53J4TFJnamzKsgh7DzNnS2uXtVDgIuTO
B1QhidmU0uWs5HUL2qQvvSdLDhSuFxvCaxc5VFPIBuoPjCO4R2TJNr9qTp8d
jf5FSexgK3RHWBWDNgxzYugiqEti6t7v6hMlKQAFg6+b3Uve3AbvLqDr3sY+
OSNF6UkiNLVA7s9AcRPsaslONQl5RuikeN8h20rh6i9/imjnmpplLDicLO46
CB46tAeqHiTnLqS4J8Va7dguXddrG86/mDkyR5VM7zb79ae5PqQRXwlBumeq
yayBAMaVxs5emz0D/UhmBODPNhaPOm+g1BzOZHCI3PEjXBG+WMmbZHvZc3xJ
CI1+ejp2XRVYQgQkLS+ZA6XDNeRBSxAh2Qtx9yZ7pVDXaFdfJXFqoop9fcNz
B792ZYx1eRwZ7LUy+hCLTFX8Y6C5kWV+mivw+Y9w3lFaXzmSNB2wis425B/u
NNczoIHgvuMEQTV22ArSHbTTt8NtIO0osFz1sXSyLc28kmak/uY6GQIQ50i4
cngWgJVh+ZUwOunqCu+ZAgeo8pwxcISw66ZvRgIYVhBMP35j8UWdiMVQlyu4
p6yRLrFcDqtiTLTGXQZyRY9Kg1un5Mup28eQJFC4IKMSuDTRu4btKRtpFC0H
lKhD/bixKubFYB3TBVbgavgqBkUPK21gI3zNv4Q7Jy//M84s0n8A2XBgta4K
dy49ltd8rHPudaPSw3FvmKpL2Ls94w4eA3D+Hu+oGZ3j1Y7njJ+XnYSyoBIe
NyXujvAJjTij6Ex2nDsKuJQSUdouiqKiNlLZjfGTOGu+79czbUW/0hY1d31v
2Sf1TR6+OjHjIhzR8n7oQxVsDIguDdgIUwsZ4+Mp2YyEmNKQgpuloI4ywWYL
BjFmugVI3VSEx/CJMkyHioRUiG43LyP22JLsDjXXomKTnIRt9ku6WfQafpoO
gdg7ZWdwoOt/Y8WIRpBIy+s13O08/LIJ20O52b115M3tnHdV7hwj0uC0BpmN
+1NYV/3rjIfzYlbYd/KNz86XkxX+QPQz8CqqtBR5xe/LEKSjJtUBglI8fTUa
eRnaIN6L/JGxESve66jfyxYeV3+wlUhe99ImQVVz1nF66mmONmK0bFuf+GPW
oWrD2oY+9VGYTA259ohnTQ5ri5/1gPL75PPEbcdrOa9ajf2O/UzPSX6L+43u
WDtjm1RynOiZ89s8yFNJhIymNgphtBX3O1xrMIiT01hFbg/Ueuv3O5phNcZo
9ZBdlJPCTzmqGxDVBOS6274LBfHiIKi2frCoWK0uZbCwaDeCgYYmKCqshm8f
c/vZfzOzDZKpIPjCJ0KWWJSk719Cyk0fI+8ra/e3QDaDR/us9uuZFh/kWX8V
N9fX7bWqUIvC4RXpEq+PTEzAAg6QK5b42dFePAEv8C22QXDpphxuPd3Jepsf
IXV4G2UzHxij6QVMIQv8iWhue9TcX3ULzGKOClLDjGy7jffHS5IgclHHKZzY
LwOcOIm6HSK2YbUwy7lCfX6tM8bE2UyYC8lVPap91xywl9gx5QwdSQovi2Vo
PzMjD2r5L3xANxEzJeWfelkc0+Nb1PM4LTLdptzFY3KLsNGQvKaMDRDsfoD6
Oxs9ArEwYkows44z+3mmPzJjiXamVAb04YIzdXx07qu/xe6OKCCAk5Ii7ufL
ViGn6GVQ9RkX+DpGkMuRyg6JWKLR+obkRBtQivXFcg/6YEHZ7U/zQxzzYx3j
KFwquaLNpI7PqtQuEsn2gPBEAWTF6+8SJOTFoPx0RCXO7bkfvgtS415iK4xz
zlH/i/jgabbytlrziGsBqaIKZE2EkKohvvSJjG+uwK9TISySM5axtP7AAnE2
u1YqRkC/wtbJncyg8/OJLiMfh2jFpQTtj1e8omOk5Er12T7i3v+7s34CR0NG
DnXomreTTnCjmC68C61wqe/K6PgmXHU1RkwtR6tbmorjum3dqLVe8WL+jlqN
NJKE5ysGmZ06+prlTvdKJ3987EWWcoskX/KgFqDevfyqxBQd1QgprETISwC9
DxvUzwns0HEU83dcV/fFBIyKGbSVymbnt1JCkOlaz1NWOtmrTIH+dOzroTN2
wwnQWnHk4SN2e3mnAR71CprylJCGA2MRjndSEpy+pkSsMcwJXvPuB1RksSls
XIeCAKP0kOwvL2IgbIfiCIIuv6g9itDuPUrGe+9h8yECeqX8FkVMOxLkZM2w
D/k6RIRXPH3WLpgek/+R0diKGL6N+O3d7cjor1wlrlc8gU2alMSm21zASIu8
8AITfcdaW4Bdsu2oCzs3PtONg9Po2q3kbJ1BOtTtWH5ytYiCEwt3ldgQsRbA
JAPXcRGkeukk91iV6jfAj1YL7YMyOSvUm9uiRYrWvIOpGKo3TxjdkIpCVNfK
4QPOHyhhGhu1v2jZLOKX+7aErnVbfQuI4C1DJRCWWo18NeXC+zQkcoQcjSiX
oz8pJaGdIsHQMECA1ya/WOE3tDnhPIogXtZTCL+780t4LHd64uX70TbCFB9s
S/CldyVCd9HWA54HJZdo0MVUxgDNtfSACE2BT/G5bF0/OtRcPtZ/iOoZUGXL
zQPssMq32JZY1d9H/BvlXyg/GF3FmzGbMw5o4WDcffnB3JnfmM6l1AaBWJG3
oQJFDN9Zx8FuY/gVLEapaky32J1XyjQHC/q7d3wCbk5BPXLdt/kZKCrw2mMH
U3Vp2fEDhFHFY+WBj0ICSVEfWvjHN6nliYTyya3nch9SYlbGceWoLFkhvZXm
lz1IC79YwpM3tsihkQEqTlkRA0RdQA0OtSKpnAPIVdCcs7CmvV+O4lu1oejO
7IDra8SezYWesR3AJXwHQudTSJCt4um4ke9CD0njS9YLgdTVRkRo37UTVhkl
l3EmoSE6/6pVApOxwERWkWqGMv4BqlKXf/Cp5gNvi1SkSpdEV1XSbetIsZr+
qNGJQWjT5qhFjaFBxGOhBfJNOAbG3k/ttgmiR57Thg72sqx40m46L6Yl5W9B
2EVYz6T0Tl0qL5/Xq5EU8HL0fKh/JNVVipq1gV1Ke+IS5OdsE6mcSfLEqqVX
cOR853p4laLOTe1wGINQa1eGUxTcWl11ainVmmnzT4ibH8sgHxkyoeUegEAU
9m8RXTig4gPcDQ5SF9y3P1D2msqSR8n7rqb7QW76sZ8k03JguvX7yC/mltZQ
rC6KbO9uuQx5vMwiPVVMK/sjAteDdfJiobgw0jt8e+hrj1Ii9SD2OEF3otXQ
PZiJVRsfKfVzU8n2SwBxWXi5ay2mBM2aFzDLjKE1taCxBNc9ADP0pMysEDNQ
YRsUbzKQa7frEq4cwuzXmTwXQY7Ta4aSH01W251Xbi1kkcDtT4IOjqd9zGl1
Lvo6bHOagLgW4KNlna/umyJivKFIkvf/BdI6UG6KyDB0eLrRW+Wqty0Rv425
mOXoTSTsH8letsltokejnRdNLHz+/4XUz7bsBgIbwvBwMigPTIv598qDJNoA
8FtmQDzgieONIGtWCkvUEx53oFdDD3DoaHgeV3dym5xMzyzI+XG0fDUKm+TT
mF0LPtAfqmH7B7f4OurqtMoRKGuMReaBdH78/F7kGiAJT4iBR6hagyjG/MTo
rMg+uOKrKJVe6B2ZyEdP2VL1fbPpH/cA73SjvuTBRUxXZVYGVl1QxHlTghsC
Sblv9yqy0rl5qr1AaGdEQQ6nlGtlF/7UpzrdzdFeuG+TaQhKrLEQGn09NmU2
XsTZzKtbkKcUrJW2Rlx4qi/RsCj5OiyDRGerYLFRFpWcTwyTtISeChp7qHjh
CiINl1fqjZ/GWftWpTEi3oCJnjBGffiTLIo+LklqjxUyhraj1SZ22qqaO3HF
B1rHno3Z0UYbBzyOkvqLnhiYbgVNOaN+0Uf6rkouNs0oBiTsGd3es1ZSCXoF
oXhZT0J/KOc+pok/aKpQDTWla9ypFBCeZOEERpfiWTG6l6mbd05SqicRsOQq
LoujGsP9OLk5rjfLgwEayRCOwJdCyb5rgHyEiSfpKjn0YlGA6y9L5iUk1f4S
o45fjCgVjGoXMNh61dyCCDnKYb7KqiN+U+5FMqDAxYDoQsaINqUcN9cYbc1L
N6NY6DdTR43WaORqGByhQv/t4Jh1X5Q2l9+lblh0goV1AqHtVnUkmoJIYg56
cCZ6QnMnnxTvwBDjPfB70oIUe2nu8QYvLKCdzTPzKQjfRnS+jmdQwmSzbkRU
CusQG+6r+sC/0Lg4Aj5HUojt8kTAJjnXzHyq6B5fDWJKBlZ8GcgKBH41/j+D
9Dkqa2YzIodSQuMoa7FFOtf0bpKJ5GsNWwtPD3rgnrKUKLswE+qugUWu3/m5
FQmtCE+72Aa2Zm7EFoGXxvKGuEsrk91X/+0S29dqwvNYtvN/U/xbqtZYvDwv
ZXrtMMLLHVDwsnv61CpxGZyi20215BZAHm6S0jQDZ+Zdtn+UWZAvmr7ZVNhB
F29LqpXpL34gjV9Ho481fzAY5a2/1WxXAig3KAdwjRlrTft4gaTf6ilzRgeH
vqDZrPlkWYdezb6BV7dnANyg5HeRcfbIN9oDCbvx7fMHqGHzLVrxjybx++8x
/ztDgHPdkBKCCYSxfLXj8NSPfO3GAsG/SZW80KuVcD3V6lkvyBoRa2dM46T/
rziCoyXSRcKP9hYW1hsqhY6R8P3pzJw+0v7cXuNsxZo4NjllZUCQsd2IGua+
XUHQ38Y65d6McAD5pWBIZRgAv5teUr0/kvtSl3Kt28QzaOXFFxn4t+bLI2zx
W2uDHOtex95L7Tzl7KrLtQ/jHu8T63KV0IsaDhlfFXrLFXI5+EK4wQnCZi+S
qhSFZVX18QMn1QXDOHBRcCfFcH6GgLawJG6HniqfGyi5mszZQjkPHc/o8ySm
KVh6QwH0VMhfBxAW+NM7fVZ5cTs2iSOCz9qomc6/WTlRv672yV27/DxOy5Wa
+zZKaoDTJEJ/L26gYb4bhEC+zzxZu/Iwk3ZOfhp3dHln1wVo7DMgb0eKQuB6
B+CxoopngiNNDo5B9Y5oAooMuKsN3h6uJgQlq2Qadfcb9iF3/h3YPY4erjKa
q/ocLRvnAef0gnuclbc3dU8UZq/O1uTnd17F7sTcuizSdedP+0BFBpBpgLZg
n1TySDGuLA8/0YHZ+NE1/gTS+JXxwVVHmFEakMjm1InX3xTqatccqYV2p8Fw
mGFhHiriMrCFx19MK/rE/pmEpmA8W/p6PEADlVWwJPe5JqyoFyvTzKyuNCJ9
BxZJ1NBSlWGyrYeORTgb1Of7UwxHb2nHzRVVcs1tc00O9RNE/aU9R22BiMWh
Yh9TixL1G0sKc2cGv6Rf0lhjhR1o9+S1SZO3VitW3p1fR6fvWowF0o3XLWhI
5owgoGnX1DU4qKteMjL6AOx3eUEJoUpoVpNNoGOs3b4VXab1c46b/Blo4gKx
aq+vTGN993/8wlsR/Lcl2yYTi18ZpevD/VP3pWvgsAYwTFMXuJ8L2A5n7G0H
JZ6/HDWjYy2IWZwpf+LIJP7qEXP0wX7GHjZRoqVVr7V7i07LcqapTmeeYyFq
x6Gs3kVtsbsnFyfogCauOEhzvycOBX+AGJKgB082vO+FP/3apF/UCUGeoIKA
pJAa3EMxD2ZKyvyxwA/6veB7unrR0ifyeuvVDInFh++OTuxcnmNBnGrqkVQz
/INqA0uUuc+7gUHleVQi/9YDp9qDUfK0ft3Nu7pl7+/8Ms8N6my0XFL4HNGJ
IKku8EBalJFe4+sU50eAIkGAeLlZaWH+hRAVR5+mJWl5JrGpDB3YBPlDO22i
tpFtuxMXrx2Moz8E+j8r62d2MXvbJ/b4dNUtWCw1ZvBEshcwRX1q9cAuzuTP
GpOHS4VgCBNPMrbORdYhFtAABioSXZ8IuU96MHhWgQQRBPBEwB7LLV9JdIuf
/cZyR4y91pE1rm/ETEdhkMYoPe94/12cGGX9KaUZOgglzFebqlUKZLZ4DHrF
5U3q3efd3CJkLwXaAJqzIotMAp+Ydj/0hsZRk8Aay5On9PbQfYG9xpLNVT1w
gFoyt6P2FlnUpgYU+dGa1IYUVsAvX5aa5K8CgGPtZoHSuEjj5Uv7bHBs1vkX
AKd7sqrAHinKPUVS4Avk2xzbKdcKTH1pLjHexeNdKRCv7ehlOohkTyAth+dn
dS61xM1+Mf2gfUpc+rqqF+wA+HV5B4rq6qPNQRIb5cOf5bMw6T+1izKq8Gvv
S2GCtdVBpT2I5WRPkcIRqVh2AVp14fvCiJoVShl9jqBnjT85qQiqiW2sCAmG
s9MMM/KLAUSVVwLfMpJJ3QH4J6bG/EFb9dbm30mLRBuZ4ZgTs5W03V/UiaiH
/LnJshYskyhXAkVILcXZSPk9pF+HLF8AMCGoodjchSXv2DPMs2yLfcaGkJ3W
C0WomxPAfeuQVPrO1wCy8C6q3niES3B57XKtNKbmO+MPgMT4X/JDEOCNobmb
zoTcIGqsd9NbGbkviXrg3UWHNWgQLWxY1X3e+Ih8I2XTeNDe6enuohNSnfLG
ZMffkVRvLYGNdt5AudcwM0TehIh9drFlxshVforJwxyJV+wTWC8CwIvka4CJ
dOEMMsTw84DofZwZLsYIyb7ZO4kMWxDPF41sAPHLXqOtld8ny9DmngU+M9wB
RiN04HvWR+k+Ki+hrtsEhxayQjDCrLpfTESLE8un54XmrgyFlvK9SRkzLiqc
WErzaQsT95z/Ike5A+88jRIbtnE1KDa1dw83ny1pOQqQtseIEesuRxHxE9SO
8RtsBiDrzD6aMaZtt9KsE+MPEDkAbaMASq9rPo+gBiZpMM7B/YoJ7CmstFzv
813/qsTpVqJc087pN51Zass1oz3+Uf2sQXKsjVH1F45yUU9TgnIkaHG0YlSO
iK2GvVW3x9MEE7+F0XxqtCkG+JJYNz9yMmiSLsBNcr8nFDwucvjOQRWWA9VF
7gVTkk2EhX3siNexM+YptfrGoEnlZDuAB/U7VVmKnZtVvcFOEWn5iaqnNgSZ
BBN0nZaBIg1nhxL27L6SXIAjrCBkhOMEpow1ntQtADqo2iMUWx+5QNx8F/jH
Rfw9xx3WbVo2BCsLwAXqibRc4k2nMAJ4j7e6w7fnI9pGSi3NFWGxRpY7pScN
xcXq1Pqml195tvmIoKQ2Gx8bBFgBxbl9Rzf0+H3hEOmYNcbp0hxzhPxVqDXf
iN2rrE/QNZ7V6I8kihrCcWdU1Az0UPOU8LJrjbCkY4YquvGEGlwot1GcJx1/
SOpdA4v8175pwOixmBhMfjvCgAn88qi0jZpw02i4hAaqB8tyWRb+sGljkntX
gAfRKtUt30WPReo05NWaGg80QcUFSS1X3I8reBcBQ5olF4qeboPeXgPNELov
JSWGyoxRZivaCos7V++FWmOg1S8M5sb7SDwxosWJnminmcd0sQwbL1kmz/kg
WeCD64YRJfU+9bvvuYBO9/DA038UlO+2vPJkV8KzSmDNWgNYa/XIdN7iqWoA
/u2/o2fm5b6Iybsbmx0CC1DZIOZPqlpSm5U8OWcBqMp23xXHXz0GyPr8P7Zl
0AJ4qIds5+GL7hC62vgUIwSJGIMJV5SyyjPKSUaD/voQc59zXwCu01gku8nS
jF60K+hdMrdy44p82HUD6cOfUOq8VsCi7zrG257TmYyZz4atawITqISfhJO8
bDrw9jdFaEKFjJwFEsSYsPq+Wa5UIhW2rBR4JqKH/NFqxil31WNBQauEDzdz
EZOcvWOLgpCdZ0p0m2ZDEtKziDmU1uiaPpA8/aerizDjkKTU3c5gwl4pgDhD
Ecq7HINXlYm6Ch8u2Ugzu41XRa/5h5Ef7F2r/9P+Yqm1G2LMLUpyMe6R4yvW
yJRMxbWpBr36OrfJbi4dujKV7s+ZXvRvOHzIA+WlDq1R8y2sWHt5gRDpFzy4
XGX6PNlUBLyIdMEr6gl49pyPdSuVtnVwAmd/CfeI6UdGFVruBKh9svsjvwQx
pEh5e4MmtCdVoprTN7qwIygut62FUsP/DWYdzSIJEQJqUF5WN+RvlweJbU+z
B3TXPMlgHRbLQdqdeS7vaiwuL+kkE7SPlYeJ0vWtcsEzJyo+g/qwkPGdAGHe
t+fXWidRbrg5Gi2C+YGdnRJ5WVjIIVQc45PNzEHYvB7fUp0iu9RRzqgx93FQ
jkFjTEGnWuopLtOqqqLvfAo5adkru+UO0KRiKYnnUz8XhqAmigZV6TU+JNso
aupJ8/fZF9FjGR4nM4PEotaSkV/TjCH41beG1Z3b8l482MgwpR5s8VxFoVI+
1UsB9ooXBna0qnUeEcGzQ7Pb5nk7aCEGwADuGUt5q4F7xFh015PnYdK4hzaz
Gltf2uQW2zZabJPWEGGX3uTszQNyrNaO5TIkmCVqOfeHPouF/5UeERDeOcC9
ueR2hWC7W0HuIKnukbtvj1r2xUvlCOJxcBt7mmvvIQIXm9FBLiMX3GsCaE9Q
OZN2UvnxC9qhvKAwUCVVvTlmdK6A/wRElEg+F+mPSfXAq8HgkMj25bTe+xYh
AEGYOx01/4mcAeUuFSNogGTkOlhKQN1rP3dmrwqX01ya+VI3XliUhqnOh85w
g4YNF8KhLMr+Bu4Sg9wXkzJhQqNh+9B7TXFKcvDbs/sRFQUUaP4kjtmrP06p
WIhAsbVS1IVSFISgpRnjNiwyIuQP+E2veXRe7zwU8vBG5ANPWv8YqB6DM0vI
JFzJKY/6ZEZOgBfFRKre9i7CLBDPS2wMaIgLf7f2r8sGfE9Hh4B5Q6g6A045
veRWOduSGsZPeF30FwBtcvSjLOVIE7rmVc9sj1UR6yPgJMUIuMPIMp7rgq7/
1TN0h0hUWlh/dIbVlS0cRaMvKZwlF7XMJxB8U6VijYQc4UEcMR8viDKYefEP
O02PEuRTv8hinYwdx1O6RJ4+mD0cGuJ/FAGPwvZHIkmDg0zwyPFP/3HIRHnf
aXYXXsUFij57H69RKJlLlLc8VithdRbpGXZo+T1hjAYCdmR7xkYb3j7QbRAC
QNY5mhq1uF4AOEK+tNszrsJCI/8NNnSQNNc7IHH+FCft9rsuXWXw3LWx1suL
5NGQpfb81AOwbOVkgQ3DSfJBEe0Gu8vHgT0LDlm9TABmUaDivqSy2Y0fwVed
EjzFcMms0wy7w5ArWGFtJOl+hHUSzgaEKYruFsVBaYhL5nN+T+NlKsMvXZjl
rkF1H/C3x8GQ83xSIv4KiWoNUOS32c8F7GtCtWN9TLjzmnWN+IqNFkhxL4uU
yodTfVxqGzCWbBxPVsDF40QN+Kge1VixSOOlTvNmY2I2cynmdc8VoK/FRCuB
2G7TrECuvQMa88wcASzwMit/ueBYkBeN582IuZ7YXFskVS+18yBY+xKhXyvX
QcSsisKkTkMpVMFWMSCzvBM7Z2QihzkLQ15GM9bVomut/h1IAXIzlEKilBNm
QPT856bd1df4Kb0bGgkndURmEL2so8ME6pkT5cBlNvdFFV7v6fAA2j3OKf3/
sTurqzUVGgpJW9s4/dsL5/FAeCeYJSOAPkhXgmLnarC/n1Ee8ZME/Fzu6QYK
XJsR328o/ppxMH47FCCzasmgR7peFViJ+OpSMVNFpPsc4SwH/Ab9BKpzHjE0
sdNFldHqyQFXxdBJbMppS0Ec3NXOuNVNRatxCboalJw+V7IO8J3Bl0fZGbCS
GZ6TlbzuGMjKSjVajInBUIe1qfo9r/fKkw3zEvYH87ZAZ8ErKqe6uEqW4TD6
8zWLKGjVGHloauM1WsSdERGLtc+3KicK4/o//Kgdci/YMJEvzIctjE+ssG+0
0oj5daej1pgwDc4NFlbWV/mGiff/WIKkjdtyz0dxc2Kd6dtYc9CvV+CQVhT8
0FdMjmUb0lde77pTiJ1BF+lo7UwxlEN8CwG6kDA32ELMr6iYN0JR4AlxQA+n
Rh5Oohos4rWS2jPP7vEhNGLbLz6ipSWpLRGoODYhVZ2HtDebgDMGJmNBYgdu
msb7XHk2Shd/R3j53Gfqzo9r2NZub9gq3Q6L0NTzDrDMHx6e9VjtNc1HpMRK
0o6QmdN9aMlboOACFt75LgXWTIjAZ+pCGOMJUo16scfh6mIV6Can51p0Slc5
rLNamcIl3sndIdk3OIh3zFENWnSzHmyRuvYu71siT/8VDabDdyMbF5C78RuA
JPI2C0DsHVsUWMXXHPwYco0Fo+MMs6eKfR3TzJR06t5VT2RWTr0BuMeI4xh2
w/jp0jDVtMRwCUo96exIh1fY4Uh4AR5bYerIl2L1BQFzZ2lgRD84+Q6KenXm
qqcEGxlDLyf7VLSs6U9JvctPvXrStmFnnKfShWkV0vdQWh3C8HbsNRamBw92
P9CB7CdKqXNUIT62mGhPY03MDq4G5AOyCRi6YsRfHO0tEvVB01K81LXxZJTd
lF6h5Ar6KBGx9IDy0K/nrXDCI1iznHn+ZXrSs9HjYW/j3TMESf/mcFjNF6ho
mC05IgjqW8kctb3XI4ACJr8ik14oI5RsB8JGg77K90jsPCqsWgZB4BXNtkBL
GlYdJCyq8QqH6fBbLQoKt0X6jzVWtJz7BaYZEy3mxAGvQe9ACt4mwDg0j+sF
lfHxEqfh3hcLQnCT+UwS/iQp8IRu4JX5Jo9yIsyx1Q9EeGwtbCGWDMisRAsq
gWC9QU8rs7Sl6ALV5i+w48kmU0fFp8XK/wpcMC3AmAkfyvBr0YZkeOn/t1bF
zM0X7o5CD5bm8g/fo0I899II/MFi61gK4lirNYk2w5jR/mI3dGZV3BQUy/Zz
ELWkgrVn/Lc5+q3u+zhRhwgZa+kD2Oi81Z9xbzYI7PthxAXcLlLvGL+G83jK
IFc3JQsEyuyngSKu3DyfEd9ii5PKXe5fJ1fh21FQ7hJoCtypgD7PFPwfuPb+
VhiSYJSMQ7HPM83AvmkHJhjGQOZ//F0wiV4oGKyRXxJ5kYoP/5TP/pWmJZXU
/tLzQJ+qW0xVF9DTUrXKpwlzxYTPo5ULqAlNXJSfhDO1xwaPAcoMR9yKw/ai
kXkUixj8iUTvu9lcaQM+ncbeg5O3y/s+VJ7xP8FVb3TgcBjG1WQXq2C5C4lt
ArHFrnlVJimgOPCav36mGyNlNL3qLBLUHuMPumqKYQbs/y7kFA5UM7v1Qvne
KuXUrtBHBS3XpFBpIMXdKmn+kXvY/7UsSCIVnQR3VksaCFL8EfBOTphK0eEq
PpL3E+cd7Jo6/jAktXO4II/+Zgr4obHLWaDCsNGZg09O5Woot6YxUGBSBJZq
wPxiPU+Jn4ibV6jbnFozZttNCGCrp2dYzUmHoJmvrOOogjF2SsW9430HXMq/
hE0vGFOJPw289VIXib+qcOiWml3519PbDieFeyDG+UTdo7PaXWaOLW+T1wRK
w7+Y6tNd/Yj1Tqexi0qipbUHNvX77bkIjE0iGrSJqMZFArO2T5ryV7zzmz9s
tmZk4FFV2Ulo4jBbj45F46s4AsclECSDkEL42qpYnkuCXzAf9Dc9KzZG4Q+d
27KlVXANF1NVzIf/ok2sTmpNoZ9WTiUo9RpnsQaa6K/93VJbg6i6OANuMZDx
uIBcJBkCXK84fNIwI+gqUTT4KtoI0C/L5C4W71xXFgZAcuq5sjMkDoOtUgY0
kNmAIHpLjA9dNLTZJpukjeXWQAZTYye0dVhtCIBWTnk4eR9gK4OABa+3xCMk
OfFjCIh5X4tdOKybUvzUL7USsk2/CKnAkyHhiPzV3McO5Rs9g9T9WYNLqahM
CRlGbkGPEnUEwKivp1r7wnrWPo3ashS/M7SWE+QYVoGwI9MTqeKY9LCtqeHX
f3l9oKKNwcd0aiLPk3H/9nTfuBYSufgimQpusLu6rj4hJ25suRfvn2kVhFxw
8R5Dqmy/RqyGXnQD3/IzNagAYg+2qXaEr/0AkKWi3f0+A7aezpgQPy3yDIoX
QeBpZ6qWyzFHjfIrOxwSOzoq00zg76vs1PkojJvlXb6eOQeq1ciLzlI2tWC5
+2jV/UxvmMFIofzwI4+exbHL3fCqvmWhneCwX3wmlIuGmKpzRjnMVwfxoX6A
hwXGAofVXPgVNuysm3MZY+N1ye90A9X2IrNDm4pnfzoCBfeR0ora6qWN0QVF
9Qh6AkkOEN/e97gu28HaHZ0UmsUAOemD15T5aa74YhSFRuNLlpGkuXiKnMa2
onzd7hQgS/484K64b8adjcrD8E1gpN4+6CfXtA2HD5/Fakg6sa9yBvmKyiSY
Mniv4qmF5ng6ur4GIi/T+DExkGmYjmN/j/9QZRktaoAhjIxhKWAbDhq6jky4
mpxif3Fko+H8J8DBjydwaMhGClG3hRev4l4J9krb61/cs76E3VqYwQHCPAwh
wAcPv4Q7Max7SlaBv41nTZODVb2dGX75OIQAJpYFZN1Y+03LVR72qgCHpx7L
Bxw9Eeu5L5cawj6wy4LxvEBzPfWSP4t1EacwJ0AeX+B3cy6cQ4EbFIOF6ZNF
5c2UMp6fd3e/s/Y9FT7x3EX/xNja+177oJ2ZQj0SIodKLoYxytqpXfmo5bpk
ppo0suV0R8exX/nfbhZ/Ik+DyQChrEDt5y3UVdeEwBuptIgOMxAxPn22WEN5
9QgCS/xWI6LBqKd+ByxCmfbUgkXr3N/mLrSGagXr5HRepsKW87s91Snabp82
YAXiAb0bGJyMNIc4noR/RbMnul3ofXYXwEuOCi5Kj6zpqlFxrbbdh7LUu1i2
gmJ1ncC+lQaLKjNjvsRWNTOpp4m09srHIA2waeE+jQh8jOeQhIyocD6enqS7
7i0cxFacSYbK6kqCxls2OO04Ru/qvtIZLWXciLiSmAZOSlFsrspQfy70X3Mf
KRR5WkiRP+a/mhpWkusSRss68GmnnqDRx/1oziArsDxhfizjzoHobJlaJsf0
qLicyjpMXEUkzWi9SfiRETZUzK0Bw2VtU57S2qMA3m6dDkE90Ct/VNsv5Ftw
K+1TqcKu+jq8QxPcFJVuR8CC8+vFcktXCnUqHRodidwRXFTrlxraO1Z8wpeM
areIRJw52dMtlJ+RzObU0QijbAN0FtNXZ+hu9tCtXdf3D3Him1/eOLUTEPXf
GUng718Etg05Py54ckJJbzhrA/vI8E6jjX3GQLtpCXz7ogPZ6HWTLZ03oqgW
byRrZQZ2OXUyImKZzcuC8QVkg9M9KC5MQE27P40+GyTTTm/jMtGAKJSkoIFy
QyhaR6ddsat2lkQeMeKWjkNbdr+jctD0Ou0wddeymOBQpFznXZnm3jZnPX9P
9ll8oFJbJLJLRKQY+NPl+dgp93lgn7V9uDG398ahsZfJeDFzgp8zM+176fY7
FzD347YC5adMA70B37CDZrJQlQgnXbHdNyC9fp19uworzCFw27RZlIksgXUq
1TK40Swb5fvcJ47WtAf8/hY2q2A0h7FVO/KbR/8iOykWBmBzGZZxsre+Qw2H
1JGEq9y5+Lom/KHQ3ZlCX/OntpNgfjlcizD07gbhL0NJmeYkB+L8t61934gs
zBK+MD8a806NwzyazuiN+IsNCDiiiTuiMeLZ/KjA6s2YyZVEDURSQnT2+GLM
delKm6sazNd2SwmNGG4pHLd8F9hZTT1qtDgr2POKKBx0H/77AhPCva2ZQvza
IEENzcY5Oo30IiOeIcjKdkz6uOrf45fet2hQ2QgMpIlz5IqUO+tizkYNJDId
tI1joc+g4STgrAht6Q4QZajl9CM/uOXwFU92wv1sf8DHiQvxckRmzSLrFKAu
JJfNe2Q2D1h82h56IH/u1J0twkjhNCub33vpd2HMOFXPl+MIeyfHcM6DZTH/
edDfpkgsfTG5W3H16YirPyFlhCyR3xDzJm6ay3PpIeBiYlD1VQFfSRzT0Yk2
UwoKQsRZ3LiqoxGydZ4Lupcgqhumx5Z+iegHbWH/BPD/VgTNUUZHoEsouTDf
cl1HLZ4ldjuCg24+6unRzo8TRIQpJZ5GARH7LLp8apnKIXrl7+e692ztfAJ7
cGCyb5JYbVF3QQBwggnzVbomaA9fQsJpOwTxDlrf/NpyHhRbLsUjy+uY9/69
xHlxxQp8dq/guCoPq9K1lSgTapQXYU+DJEhS4irevoE4e1k5E7hh0DvurU5i
yhKbJeLwepOHxgDgIK+q4ov6gJ6XRw9JndnUHFIPvPxpuqY6LeA0bnwDYZJ/
Kgp/YtF5fQaX+M6nuR6Hxc6PfwS06bUD/x2cL9nowrDlY4J00+YpDSPhz/gl
MAG4Yti70tu/lbCLVULWuXk/QrXn7zNWAVWRxkqczrOZwQEJBPz2BdFLUCfJ
vWoiexJyWHUtxxEaRYujFvdqBJ8+bUiiDMpIxtt9qfyS0nwRFuZTFnmy2e/E
Uctz2OBHF2INtduGt80Em84cojXvQGSjjOsP1PxSS3uKb/bTKlYcz5eTMUuQ
5+sZEUTNUupaDebQFv5hQTwEmPmCbmd8jKdFwFaa+AGhYWXZw5vMycE9ZD8k
YdaAyBvUDqzg1EOEYjkwrRO/sUvWfL0sNyE7rczNaT50e96wDAwB+QBrFY2/
wXvhJ7CdPX53uugPQ5enHt8pO9EHGh+J51SQc+/073E/+QGDyS/2i+kB4Iv2
mAP8BrwmMts0zMiJnj5Ql2lfFmm3/059637qZ74QSfVL+JRuKVtIo5WkXMFs
0l3m+2eDcliSksntQwc03OvwVUkAUjd/1aEK+dzJQC0BjjtlWz51S/nB3iui
CRzqvJaQ7tGMQZ9R4MVW2tyTKrKbznXT6A4vWryiVShzxrGNqxHBLzTCdOpa
wct/tYmhaXjLFtw7V4gDbQi+LEsBycImx2BCKOuQUCP4HiXZD5iZPQFa1k+Q
0zdMKAZarsBRGg3YI/J+nEudnt0KV+AP2e76oBjwcX2SZKDlZ6ag65/8wfTX
p75XFaoSKzvdIyUOOo8Z+d5+VK4I9IlfTAfEE695GxHgeNExlwWJxwoKR+eP
+YBK2LBcOGAY+BrvtifZJW1OoCIkGbFCS+gGv8pQLgguwqEhzE+xYxV04Heu
Of0hDYkEaH1SVbz6EMqZVGM+WQSN3s7b9o39ZhfloOq9MoVZ7bljrFGa+Os+
lqhMt0Ve7gfU5LKkONFhf6cqaqHe1sOBpj+CSlyFEVdvC0HegZNEP1E+22qA
Ltv42jgGmV1ponsDe90PSejLB58WVIkYx0LJMJeJlW6nub0t3rG3Jw1R25qT
Qj9ixIL//GdlprtaPy43/aQEo4HV9uSCObcZbMwnGqbEw3u4qY/J/LU6MrdS
xFoytwGmDrzraGi+nwmjsWTzx1Pz/y9zJxKM2XXiBckcjqXxwG0kTjWZh6GD
F1RgrLo3lEXqwMuMQZ6DeqfCRFihoyvB21T7tUQ7MA+EDjdGM8HvEN1kJNUD
hCorgFk0DG8aATZv5pKyJuRv6xJXCUH8V2FVjAlv9PQbDofxoxAAQ4dQXT+9
4Om+xdLmfyz3j8tdBGn5drWbLOacOphDA2neA96hb7QS6O5ZMF3F86rGXrwd
s/1AxRGtN0IPNg5XI5KWuIWyXRChtcWtK0ei98P8w8T6IlFJNjGImVgy60kD
Z5jGQYnqzE3CBpI1B9scQnYkCkcgpH6M2otJROAEH4Lruzux9j2bzvche+2Q
cvEtRb9ND8Atrg19KUSH5HNyp5Wo+7WIj3Jllj04D+s9nXQMk00cHsHccdDg
ew99BjrKlLMgYRQIqt552c5uDNK7JU/8AV6efwPGerWkZDRTz65co/XFxJ8N
JzLJTFCgwtblfVaBIUXo9JBtj0IO3pIVVOTLflo3NKFZR0t2R/8yl9WXr6dZ
2j1Scmk0AAc/dQmo3ndDgpouJreSYZ0c8CECwqSkm5nn2nD24ylDKlwwQTMW
u9OLhyjf+ijMWXSLzfQVfDQEmlYImT6lMWStfj+ZEdIXHlvVBCB1bwZvFznS
lZgzWZaO85oJyMxdb+qie62nkLolDRzQK4z51SBHrIXgzu4M88bnt8uLqL6Z
hfoSJBniVoQu0/3G14N9GFLt964j45t1yQqTOsv7bgiOIGBeGSTUtcgNzPbh
cxcfm8s0bUPG0dIAnIUEmog6d4BLWditODnFCsgNWiwpWvJ8d7tGsHHcItS4
HIlcV57KoE9RsQYVJmuvW3g5CT/Muip5hSakX+DPM9LAl7Qjvb3Ak/HBZ3Xd
QIDXUpVtYh2G5/JJf9ZsEfxV36tNoivHcc1bnxELDppkOtDqgOQDCJ3o4gn4
tg6VPGxlHLZKbwP6sO4CdgITw9M3ogkZWW/5YLdstCCQ4YiAHjL66IUkehBR
+e3od9Lxn2w5tIKi4hJyN4eL7Im9XyKVP2i6VrKg87zZ1KrDSwDgv1jw8/9K
oHPzjErwKE5m2DkpHhQFvwVRBICUjx9D+JyaSMZ9M2HAoGf+uBrJTTAiyrvG
HEL9BP5XNMwiakIAe+ShP/r4oBlr4IaFhl27+Fzlmb3XlrgitkX9dtyLVfqO
d8F08zKNYssiprvdv4gKtPMIHBMVxIkLPpP5b8g5f+0TUhF7cuTEhUAXp0NA
k0qrFjN013Ny9XQA23Y/kLVQrpWNHvsH5Mj+GWemx44gWA4dsF5SxWxHzuHM
PJPaG/J/gSHlVCJRytCDTYSkodLjg6tsdl7Y5cd8aUXvxzoRbqI6nAH7itmB
F1EB8mfA9aWnVi21cE2EhRph1mbrSCgocFcGSODq010/AdDKMSmB4wYrY9wD
JgWwsYhmSUCxA4p3sMZzmvfjYSzr1ERnK5Kw03MRZQHJFMgQBGcq6Decvhej
ZXv27zZClh0aRcSBU72pzZUBIl158CLu37IKbJGNRKOvfgkY9cXkpOPVXEr0
aBKibFQYa1544a7EKER9TXD64qCSdI8KXZTKn+9JUnvHZPF9oxo/nDztTCF0
RFEJEyKZ7kaJpN17hTBKr5qLE/+P7oW1zvGXKLfCkmyLPVstX1Cxm2F8XskD
QTOY5Ljjn3aLcBm3Y6V6HirkRMae3mM5LMllxc3kuhTPoEr6cyFbmA0Cr3+H
6frEyNtyT/9WTvPKFPe3d3GAlEtj6U+IfkNM1NX9IdYzWI/9y8o1Nr+up7QH
Iy3pe8R7Z4Ga51WpJM9hMFozYSYw1F+/wsbadVtkn+SiRgx5KbHcLrSjisz9
dWxaXGP9eeZwmJ5iWPPCYIhBu1RXBbSHUtLaajMfnGwLK7Zxx6oOtxVHAebE
6XqIZsxPzFOzosFe2YJ5azLd2wropcZ5T6kHVXcbCO9HCiicZ5DrZFf2gbCf
TqJav2ut4y29kuSINHX95z7PkVzAMjrd2z0rONDff1RxpG/zwhZUIkyG3N5f
Nu6GsMzaqHjr1rQlzOvRIaQG2YO5n2b5CDA7mVWtk+dUWaxDiyG11kz8uHxd
vgYNmIm1NsHoXx5HWoeyj9ZyMk8BqGrdw7R4F0zuRGl5KPxJmFuSRauJbwCX
keddC3Cb5ik9OtruqHZykfP0acZaAoNxFSt2r2JYqwD94d7Hs2q0uqu20Zhq
otzCmmcMyE1+0v7Xm3qzK6yjpAMIN3ww9SytU0jW/YD8YAikjMC9cAR+zrAD
AKhgWprMN2gwJ1vWn1mBkNcrV2/YZk61RKatStcEpNpacN9iUv8i78jjZ5dd
PLvW4NogSmKipeJytZJTr45g4VKeWMg07aCtAWumfOemr3RRqC+vbQNtKBat
YjSGYESvk+GG+0sS2LjaxmnLERV7d9aRUZ5Mi/Nu1WcfDL9LcgKgR5A46YYQ
yDWLWzVRObrrz2oK280dGEO/VW9GNwwAAknsxSn0RfEZww6kiyNzdqFrxnl0
Ms9Ok3LMEGdWfsHH7kocW7CkchC0kDGfCpN7dQfrGE2zo63u7Y6Oe8//TMSX
DMr1779vw9xPOvq56jgQmNWqIDJKH7F88VMNWp2P/1xgaSQWhja/Ge87o2/7
qnHZuABSlX7Y/U+JZLtXPqauHW7S6arQJFTXjqGdqviSJ+XAcR6lSwvaWe88
DPAWtUlF6Cq1yLyVN2IzjHMvAZcmr/h0baRhFacZPN99AcwZFE9kqH23T7RJ
2Dd8g1dEnA5VDq199Hl9dgURWZLev0TL5ifXY21msJw0EaNT/LB0s+FNVbzn
aUh6pADkfrB0MsvjNKnsz3RXrFiw0givHVY43XpH2QBdxEqW/VsUxp9aa+yt
+GYiy6RA15qT1ueWzeuH9JPa7xXc+Mx8dP6fi9n9uQ2TZCOAQROGw9HYotai
nl2i0NwSzRMHHOAisB1gl+YsV76nzNgFzVDP6ytY/SYH5xePT70mv4e4C5lP
lTytlOhnbsx2kghsnoogYod/KsyhAKJc0yfmFCnW5jQCjiwaYpTiB4dY9kr9
BnqnAFMMBu6orhObg7JQirqoj4kbjVuWvPhKetUyOFPniqG4JT0gQVRJTd/L
/c9KTDQR3g/wNwaP1dP2WnnI0jLorZ5bSd5gC3DLIzBuE8PEWcCpArmeGCpM
to7AtVSxVFvKNVeveyji9w3lUP+H7OrVeiGbIhGgBmsKf0VAzWUQ00d6Coh/
8TVX76ebK3JBVtJpFT4OdOVPlQDHXSpkCMeyy8r07MKC5EvUfn4kxBra4wfG
BOjIZzsqVnJ4n4GcCYf4rnWBkQjIUQHrqzOjVNM/+ZNRysncMAWfFF+wexxx
5h3ZcyzMVVUjJ9Ns828tFvlRrWG577sgOcgnaNdKiP7SqzlqFSLP9taMsfgx
lRopBzaQSfHKjyJmo0Qf+t89hxlNm9JgNEpomRKuvWStkSdcQZMuZfteTzOJ
ovdMJCkvoWXbOYhxsddAxRztHlca7P5YkFLL8PBzwJXa3z6hxfeDrVivf83R
FaJkh4nLX8hPbnmPRk7Ysp/JeCapY6HXC5Q9SpP8rnLA41nsqmEX94ZyU5g6
WPp0RCDY1vQp8Xu7w44rKwL1+OrT4e7ClbYQPGErd9108MKVC3Ekf1WibZcC
AJNxB1KaWbPt6zp6j7NdiupACUpfkVa4WnSs6A1ZtKe+D/fFOsuMwptK9dkl
tnkzzZWZUZ6wWyhoFWOSJBaWmT20DfaSmy17pM94oOWuuGMOHuXNOeZEnRdJ
Emm8DlezEVUsv0bQgBWIFNyYd/M5zhn2botHIKf1uQ8QzfR43tEXK5oyktyB
ZiQWLyd7bb5AHnCXzRB2xwerBWeb0NN0LZqWgwOrT4gYBXOTEOQPAAwsh9TC
sXymu22ufKHsutst/oG7ncZjo5YcbjZ5QWi0zetMHkO5OfXtC2Fg+a0zwlW7
jaLKNnfX+4fRRk/Qaibf2Cr+QcEUhy9qGTCS8jl6W2HIfNZu2BxFhVnr0m1x
VuVQAJGiFhpMqOiuVZWJicfnSWEfdTFVgLXDja6bDPWzfjwHWkEr9jHG37W0
j6n4bq089GZLfpWIK9Z+1BXFZkVAMhAoKfg8RsmGIZgr4OdSySn8D8mg0lEl
F6knFNZ6++Rfa+fcFDoZQy0gsglNqI7F4moK9JnagxzYzg+Xzodi65T4ZMDr
4ajIn7zO9vf0bEP2Qk7QJZtBJMgGsZT4LgvBUEb53TncXAdiYQ4roXdnL8Wt
wAqvRJx5R7dXx2v1ljpXBc05kvbdXeX/vdap20PuNPyCAX2W/rZukIsg6VJu
BzX//QaCnS11RSlF+4DqGtwMErznLITcimvVzENAxZmcbiz30gonIW7XbUai
JCcWrhKu5wdRT7IvZepUfOcao7MKXms7VcQTzZDL1SDsq+Vo8e5S7EbmFm8R
Te+WOIxe7twDQUK3tjU+TS8c3Ovl2tpt5WlnkztnhfjND2+n1wbs54LCyMXn
ttW5HGdYmmWJBilv12biZe9K2ii8JMtSMYhzlMtl/0NNzYLR+1OC7k2TJxjz
Kpqx6w2pxoxkJmPPLGMMDgZc5FvLhEuWuAeUAn9o+x1Ues58N6L24Sx4StpK
d64o1QCB30odZS7bOoPHp31SUPUwC76o5VTuawL/RBZzRy/dBpK4eDPsQ5Rl
kzZYYNhPZMaVFX1a4UhX6S6MhSXnOep1s70CQG2+QrE/rrhQ63UgNpgHhUYm
uzl/U8J371RtYOGXk2bx1tPOKNMJCaJn8hYqfMcgQ0icca+JcjJCtf09Y3Jk
BqgCusk3Iyg4iNxC0s1HYByzxTtQ3HMlchF91vYmmBECbqhU+PhAGO8XPq/P
8lSCS6FmC8xNijPsJBoTX52Tw51DMVyhv7+67N+vSYhEDs53JJmaQgS7tO+o
UiIkD6eJqdjP0icClW7JbCquz/K7fPInZgLSsrJrhkdxZNBT0AwGEtAYlJdj
dAbvYnWnbri0nrHBIekwkmOGJ7MU5lHiHskYn4UPzwQsMwXzrzuxhPOobEw6
sltE5iUksYgmvfoVnvFxVqGPCT/gEzSu/U4MxPbwNEicsEzFuwaJ+br1EMoZ
wCuXzb1Cxy6KD08CKPhs992VeFiExniOKFyQKRWdGwJofvT94FB8ptk3cJHU
FtmwVKQ7lJiPLSf9d74TYM4KDTx/pFM6SxN8ilnZF6kWKpx29rFa0NnaaL04
IuuUcgMLSJuXnQzOvPp1k0U4K1kMTQXcAzHbe31uEb2Odh4dI+6QjzsbkbpA
QXAgAuanwnusmkXvJaPCwyNBU6AudfZA6+nrI4DKu9HOg3Fn5FiBhuGzB+Po
qfysTYxxdf4S+whtGfzv20qAyZrZymo/ye6bejcIxgqgQhfiG3zGmlDlrsdp
7MHbRidWDGBev6hQ/1vznn89Z78ZlyU/VougvIvtGpdZBYJ6sZHX3h6BQ7px
Do6ihald4BU9ijg6pIZd1gBRGHti+uq2mcGrc/Q2wYtdhQ3kcE+FEm5iIgqA
ohgrYP7/swE+w2CDE48Ns4NdFKbalehJWlkJ/TKS6CXkyu6qfyg+UVZdl66p
U5U2zwdqHIUrVKYTDb6moyQgwdT8RoKQMJmunJQHZaroIRpwF4KkgGAiodAU
SBIEd726nBmcrL1kB8ufV67IUscSAbtBEiAWPL+KbtWU03ZoThZCeLMFfFTM
jf6Rkq7DZLqDoN4ScR1Pr0vMWzDw+UCgT9CDi820tnlE4sLL8AqJlw/5EiKC
yxGALVW32YgdI/XpKQmcmC7qXlLSH2zB6Jhwj9nN+hb993q/RcC6EW+DuQW9
ZHFaQ3ZgLx7le6y7e/ItFQQp6iJhEgpbhxXV0kByLtHvd7NIqmMSDHY9XTIO
vFxliquMNm+Y7YA9bXSsgY2AsCWJNzQiFh/H/faFCmA72U+Pe6wZ48rv13sE
7GPbPqrqck55ZxHkQgRL99Z4LWNSlWGh+yFt/txG29EmSpvwVrEH7yU/NBax
YbfjUzR07+9+/t2e/6rszSGG7t9p/GAjh7NOZ7rTbczViF6Slp3rtA/YGXHQ
v4EoBHDVaEEX5pBcgYwMXUGe5j7jK3RpYJoMxXpTZc9vPvAJvNJ/QHJQuHy3
x5+emA4kdyHwGnRSE8sEcstKgAjK805126vFBRkv7Fe2s3YxuS5qivHTD7iK
TPw4rCAjTScOkkd6mtqMtDXGIrIOvRgEw23kdiA33lUyrEOUkcKWyS6WjFXw
lCEmbK4v2OONzz+/faghSVIpDEViDOOJwAj1rPzeLFulndRF9QRuvcX7pBFt
yJ9XvA4S6X82mq3c1nNAiUafozNhobJRnisZeKQ1ePuG1U800yDCqVcCQ7d0
3L4Z0oPcxgA8WurC+XI4H6N3JJjfPKrbYABl2HPdh5S/xPZhTJndhMVECKhQ
9lsBcwAodKKC4xIbbDKyqY9l2DKs1BC+17bcWqyKpxXsNSgROn9eQuqj5uNE
EL7+ADxkGImtq6xRrXg+5SWbOzAT3OH7b2yTojOXaGOmPrE+87RQ1T3Mw6lj
1a+tpLOoEtF4f4v81P/Lh8cIZvc4SVSBPQ5lhZbat41q/oHzArJDzhCCh1EV
onfWpsulxzLBhHhQhhtn9vQfJXMbr8pa/8nqOYAI+xwQJHOCNfY5pOJOB0g+
zrN8irV0UlBVOmHmEhHKUg7X3TggDYs2g9g2tw8iIKPkouiCx+c78048dcZG
i3n5/y9LP8JGaQWti3qgi4b6lRBQxqL1f/cCfCzZCcsYKG/dXKDqJ/rJIyke
ejFZzjQr5iV8uy9d+wTwkUJxCpGlxFMZDOoT/xztt44+feoQhu0/5BlS9tfP
UnVZkN2D+ajxGy4VgGF5fgtfkcxI3XfgCbvtcPem0mEz6KvffP/qMXiqqavp
qdMRmKQMnfutKdS1R5u2hdHoCRVcOZN2k+PcsFa3VxA/VgkDcDswR3jEVywf
GO37U+ZjA8T7OJ0d279SD0fln8Fd+R5WjVTS6rnXUqtKyODHCnPo7N+5xCVB
rPUqpqPxCDAfpmj6XhF8jVnkPj08Rfp0LCylZbO4oFo22EyEucnfzNoGiid8
4mdV2IF+VubS+Vjwh6zIV88AwZ+MQZb9oaz/ZOt1CJQ4q9u3Gfb1U0EVnMXB
DWW7qa7WDb3aQEu2K2jjoxd1/HF8LoyGRPqgSuZ2zcapFQmLTPFImXim+tUT
OS7CSeJUoCzd6sgfjQcJO+TMaFq7ZD8sLNcDdBGtjaj3r+rw/Dk/Xm8asJik
j3BvrVg/PVRiogOAN10QtIQYNCPxxvX0L2IjuuBtJgKlKrKUWbXdjKFJmfU8
jrdY61x03sE7h3I196B0b2EKmtXw9JSTggRKUlYnpPAfFJ2bLZH26YtHxDOo
zdkpigjbZ/hYvAieAd/bTHo7JcjWMTVngN0UgBGohP541QDn0+sVIs3m9qaI
9n0Qvj43oWwuMbtcoDdOkdN3FXGVy9FanEIvmnzKd+xkQrolEsMSWCiwH7YE
mWidRHHkiW7/KsHOhvXvmz3qMojQnTxUox5nq/1qsbLMGgt9TpsPcGxuK/H5
l0Jfcj9mnJaOvqeuE/DASW0mQVrRf1RR9IAA0MDWhzUNpjgbPuQ6+W33arSf
z++XJ8Yphi77LGX+KjJ0KL9t7Hc+J0N1RFrrGOXoTcYjSSxfZtYOVE2Cr+pn
v0NMgux++hNb6J2MbvZk83ZL3jlKxsc9dWxWkbHJKR7s0qkq+usgm2IVIVi4
1vdixbKGDBNprpGbDZEyDwHMLbnLRdmh8CdbPUlS4OM/mR8zV0F8BOd4gHRh
76DcWxwnE7DZxFG3FgEE38QWhFsdyKNjPFwUGbJiIcvg17P81HV9RtNDErmT
e4UrLLeP4iBecxKC7VMQjgvdANK2fqAUZFuiKw4glHHU8K5oksAxvAUxGEq/
PUBcYIt75PLSc3xqbnGAPlvvkoDdinUZecSCFr1c/mqqnn8FPpMgR7zdflCH
4dMARurW7uLmdaljal6SJK99ABv22L5rZL4j+gJxf1v1S8kGj804ZAfZjCbm
cExYLM/5JhfzP1ivjbkCw2N51IGUjMobturronrmSb/Kd+ci3iYObYHV+R3s
pMsdxkB14PW/Z9aoQxNddsSBeZAH765AVUDEHUBAeiOesQD/escNVQz9++0I
D0sGjY3h82rg1iQH8aC5iLofwclhNB7y4zznpl0JN+oDIU5H5MscSg1Od+0p
+FukxaltHx7tg/JABzqqifp/pVDUgUy0PIBp0CG56XUVULuR/5XDKVFTNzDw
T72sS90gl2/EC59MC8DY9Kt3awrGfSXYY0VMejuo2tJF8/tbnX2S+OQIO8+z
DyrTifjfMhzlAqrRUNpHKdKBbN9W0vrPmj1J3+k/P+LzE4C1hyaEEcawYwmI
KUcSFoAkPxnG7j4yEiDcXQBOXfaAWiNRZ8YHP4Bz8d8dnKJzY5q0oTyXhVLP
yVgSLoOy8PG0uueRGjONC3X7SIfmx+CwxFRbitV7Q7NPSfdv2XDqwDbaygOe
1cHNE5+96EvkBwsJx9bPBDlPcX/WRAmkEMRzxmoBLtGy7zi+30Astq/NNm5p
FAnySLcRkVnoAiakDKKC/GkX0tcBbwsOsU7SH7UbEBhq6Cvmh2fHXb9TG5lf
oOxPbdEE4uTmY9zNP8zMvY3LcJZsYKQS0byYe/mh+ILq2NggxRfAhXbg6Kq2
gPp2b4CPjURbgCt1TehO6XkEGIiw4lFENiz2IjAWVQSmSQXxSLw7opWI/x1d
Tfxke0hMpWoC3YHGee4IlBX3m58ZLMSVfucHKvGQyOonZT8h6oYT+M/R/69N
AeF8gvuAzxo/GO0DwqHX4folSkmGp7UCyhAS5zoe9VNCKLE7K/vetsfnCPH1
Ke/My2kM2if8ehNvar8Q51GBFZNucSBbgCU9QTnqouyoYD3SfgOqTrCoQV2R
p9/YXJWfq64+UqDqTk6SodaW7uYp3m4hffdOU+JrssG5erfNYhvsqEs7zqdF
PxalXndqnEYXYjXMpQQNEOvemmWeg+uI2lHj9crTG4FZcdvGGT3SGUMhEt1c
bLouffSPIAoFIIm3f/x+FzIS8z5TCDj/NjakY4ye9xIgBOxz92rXmTLoqJpN
j8yF1PQOXITV9fy//BHVwGz3uscFfDBxTb0ingsrJ46Gc+Gybgy9OkzlpM2i
Hvbxfode7DADF+H6R1J+GEDl48rmiX647iVJmK4h1W228wp1rO+MhXljr0Wz
LbGY4c0Qwa986OTU9Ml8v6GcpiOs9txZYhv/SSxW6gAbTE3T4E+SodicssPx
lFmXI9PCzj2Nbo1kKshD4e1dnZV0xzyJNfdZ4t0OCSfEvTrNSRqM5x5djKeq
dhWrk/P5vQgwzTlSk3qk3aHK9sFyA+Had8a+U5z+H7PBurryOOy/IpN6enhO
eU8z450/LgQO4vJ2/LKLkcsk4hJimCbKscST9INjKSvg5YYtQQSBUU2L88aH
Mh5u8d0ZklYG/V6FtJs2O7XIo1rYCGP1rUxFmaqScEMaGkvo8kTx8Uoq8Vll
DCu9TZOjiC81cmnEaan2a7I520EscvrnBBdsC7KpxIQGYoQHusfqfZksnZ2D
peDwhTj7SsNmlswmqjOniiaLiRSA4xaW1w/fbaTWCbo0U8PcCrekYEp9w7/e
JGZ1pZoEr+U+dvfzNByAwTCSOPN5RfWGIqynD+PqBk00YprajplI4C/w5pW+
7PGYN5O5SfkSgY2pwqZNHk4zVV6oIhsU7I/pOXmbNHwtsF7Q/h303/Jku/jd
c5sDxdxOfUr60SDbYXu77lg4LMj7crrUOAd+ztoKx8eUGdT1dfD4G63KcbLO
e5SLNXX/vcB6icxJojCv+MTxTgmMLxrebnnoAeqBoOtIQeN/VWuJGUxpqPuo
8ufnRoWKOdyWUTpMFBq3/8QdiZxe9LfMiQ1+Pw6WHTlLbqn69Yux/SZTjOyF
SJtogYhCrm0cRMHzxi3N21CJHUkf5H2eQLG3Q5iF2xBngfev/Nr0b9lO55FY
JP73HXLKBZBbJCS/IcDAyTFFV3LAwr85c/LzAfgKSJRW3t/UxJ0DM4Vvv0gH
n6yidjJsi4GXPHVNbtl6z5Oz2iWuKfaVJEoEhm7xg8dCXRxCI7Ea5gXTehxY
c89piEJwrwN+kechkGUMcCftL3N1mh4Uc3y1Eh5RbPnMrGTQP3yva4+o7gEM
TMG2ITQvn+oH0Ph8VMIkBs2ZjO/sdvTo5xtjIr0OFQXQErdZ+GCQXfemlv88
cZcHlEf2l0I2VA96S8oskKR7iPsVczyVSRLeA8lpd1QII+A+N46cSuE+P8/O
ILtwM7jdr1dcpNMQuVqVTwmRrF11WDLgWR63L/hzIKJa9L8Pp4eT457jKGQR
+lU2o7sSZhaXjHOQFt5jYp5/QgFfJ01PL7ybM/SBwfX8ArzZF0zBcy4W7i8a
NlQQKHg/CgtyiGmeDpV7lGraiOou4bT8SH2OsbDLAIHG+rwYY7nKEIQQDq4y
Ac3XDWrlqoUXA3IWW79ttPmaVf9EFcCEVDWxBXNz+wkyeHKJ88wx42vvziyp
zsOd0NJEl7K8Z9fuGofWped2vAQ/KJSjcJSJbIZxiGWx5X/gPOFm8cJ4euM0
O1EtPwVqh5CTHnoi1ZOoke0X0e3+WCjnXeheiIed6yXJgXaN1pSRG6ASAY7+
/9+PehF2Zit/fZD40jLu66w/Pq2TNUcKmeIJXe5LUMgLap3z3xwi+CPL8qmO
yLVCFcJQvRAlZ6mKIfyKSyWRYZtFPkNetL1m5isRVZYYGrWZDroIpkPKx0+p
ssp9bDrhfMXKPlzBkYPUU7YB6HMR0iOIjwDLfAoa2QQOwTbZFKSMcB8YlNb9
Nsg2uEaeYdRZ3TbIWFsYWE7e64m2eP3AufWFve9iVxJqwaZP5DebCo/45OEH
LcwmR8OikwlTY9A3Si7Yb6ivIznKlFvaObWyXVjlg5uPlSsIZy9QhESt+vjp
3tzBJ4e6Xso6rQDQ5OeNqbYFviO6HDPxxl3KjUsqtm94x2JOjK6Hwo9v8OKA
ud6anTD4ZNfNNa7eTAbK6Rh4UY76jGm56Dij2beInNZtzxWLEQ1mFNRbCLdA
fTxe3KdNH0piEk84xz3Wn4/YneBwGm6/nmeGiBBdxXvtGOhBSUpgZuVhcSFv
KwshypCEwtDRPNM644TjVzbJtU2qIQeZ0PB5Q48S4BNERh16W5gjO9ZHLFeG
SlqdFRtjqXRj1vU6sTWp7hicHqgTuSV3eaIXI8k4q+dsfDyMWVwH2YaeM2M9
8wmbHhvs7OS6SCkMVlm+/+y0lHijXYSDdTgr40lYwdP1LyfnHKB+MbWbPGeI
NgpCVzPegJryuR9HZMPRIvvIuFOZ46gkeCMO7aLSUzdTt3cZS79rk2VSr/0p
yGS/hvBEFVFDTrkf6VF0lxp8xJptYnEQkvTm5AwGzhSRp8+nZybpMCsQhaZl
Ahmi205te7HPsMOP61lOXolHgQF6WMmvbSaeIDT2a+sqUqgq0WHhq0oExPwN
3dMdYwDyIOisrdRE5R7WqxtCn3BLcKO9neitGi0nv+uIgZRbcD/HgGiwN7/8
uhE7Ha+SgcvpeTo6KCcY7p8SbYuhityERqPGOIlhpRkIHjOzLd4vTScjX1XG
GvG/4r3EGlfKGCR3hndN6RrEhU8IZRkxtqhApoUfDdHGT5m3eq0qy4vAazJh
q9Gs/Of9YRAyGxPS7LSlmLdIMyPUhAIdMHy3HxXpaInZXfjIaLxMbRSTecdZ
lDC+X+BFK0a476W84nJggZkEcSjXoQ2H612Tp7M6jPJ8FKgggZ+5mVzFDX2X
imzBI41LNRD48Fg8MJ9I1tzI7udWMS7bdpHuWbmfZVI+5qnL+1Gn03qFIf5/
JCrL7baBjXzRCggGYiyIF7toN2h7EJRXdVbRk6vsNfzWfE8a+VMqqvcUSKAz
QRsfr0SjqMQCniK9my0UbJX1ca3P68oosG86seLHdrBi1wH6HXvZaDwURDDw
sgHZj1vqX9a8cGirHpjsYJbp1UW2kYZiZ6eI3Urhd+RvjmUhbmc8Wazi8Tjm
8fPk+DtfbyGiMaLSLijfP9mGznlm9Xfu0H13k2kas4ci6cQi1iVAUvEtcxQo
d5A5iNwZ7FDuC1cPfRxnOAPKbzmA55WT/S39zbvJ3eolU0P1GCefxzDwywwO
+YmUCtTzq978Sdlzw/338QrZdL0eM2hbYHtiDciQf9/3OfI5SVUrHN8Vjchi
4mUe133Gjuj5+xPbEqL97m2VJEo7ixgduiA9me7nTZtLUp72f9mQ/Wh858w/
SXaKZYe6bsdOBWt6XcUgfsQ9Jm1GKQNG7pvIFHeaPcEe+c9M8noAP16eO5uY
862O0QpVOcRlQQ4rvb9JFnPaa7hpocEW2PupgZQJ7URgFuoqKxkueVryZBOU
fpXYyysje6+2iCPbAlalJZEq8icAhYde0jnGIDGT1NgN9O9ft5pUIzNUa7wG
yMYzoTAFrB3T47DQEU7RJc6Mk+MlQ0/rlOKORQ+V69OUyr8bc1U0CvffDM7k
rM5CGE7HyKU8CrONtK/kKPm/AJWmNndLfYny7v8Wy3YHSAVzthiWeK/1ieC5
WZ8gVqNamvI+XiVqSNuT+0K7UsL3BQ6P7/zuBkjb5KZ7MTxznstE+ziaVnsH
SVGw9i+YMuUijn9L128gidB6aw1ypOOPzfzrwmhRcLfZDmIbLP5D/iTBCfBX
Np+JahrFTwmsJfJZCoRkE7JlT2htRvCEiCQ4Ljsh8yPexTADFXkkLDNq+7FY
YbVwDowiZNGfQLuOSuzwGVBhpouxvDuJvLnndGa+yvzTV3DiAJ6XUAUzqU+j
jWVWSemGYVB68T5rf+QRJ+kO6ZYYmJ/o32hy2959dZTHg7eXdUxGwj5+Gvnf
ZgdLgTzUq7iSLQn+dzPQ+zP4WBareze9LO9Nax5GLH6CfEJTv8LhPS64fpmt
dG/PpL4FGabtlXS8dpfVOCdX69NexnUXXQno44b+pP7MjNj+a0P69kgsDIbO
UzTn2d9D6YH2grKzJzZ1Y1CJNAqji1ykB8pV8L/VX9EUPh4ZmKkkY8E5evJW
ONnHAWykRThDknqVebdjDsiB5GgdqPK2RYlBrbrUcy9BNTMTIm6rCcd7FpJl
HD1WEmQyfDgxjHP/wy4mR07f6n0CfdgodqWBF8532c+r6bDzhpn+3ZZNcWRH
zYnTwGWI2QGbbItY2MX/4yz5EJhieqZC3r5tpLDnm7w+Ot//lox84UDP4tyc
eo/DUvhditerg71ealyo8/xXfJTaUtmflkUiUiRCpR0SIAWijZAe7l0P7el8
XrcbVLPmaa4voRXsEkEmWDa5yKZnkL5vZozYSgzcZSeSlZKqIacN92LWdOAy
s/xC0bSDu7kZ2OnovAVtoB17P7eJVuTfvoZpptHIBsZ7rwHVC/sjRK7U61iT
8ZW7vRtLwFw/UFwuaQQInAtqK8S1vxBNjVFsvJwKZL8v7PexfkpX8Td1H6q6
oEfyVPwHyfU2xV29e++fk6osG5tKRAi8JJNmZdZTJseKuE1aetJfz+4hotnO
FaMj1fpwEQnYKKRblkguWv/OnP6xbpn+nZJo0ilFr+FXpnMM86odGREwt6bj
3f4eaCsiMxILJ4AwXJDtrOdJj7w3gRA53tzUzmAOqAds0avbd+LggVMLRjdC
G+7aLQJVzqszWICAlZqupjy+dKj50e+jbPTB4cMDVq/DvHFBlGM7TUHRmWCr
o558UYuSMqVe07fRbCCAdG6IdVnbkh/61DFffAcoTf4GjZ6or7W7tqTw9DoB
BzzmRgsSjR+ZqeULjccm0ltaYpyheXE5g6U9nyvFwkcBFY4WQxn3UDd1FR/Q
pOvF23+C4lMEeOA2XN7Ml2Oxl0LNq+eukLkjTlvYV9i724sY/P2c3oTMB0gr
eCY/OvEFxg378S1Z4Ku9nmHqrtw+n0YT+vrOUfTOTQazUbyjGWAK57yeJlQa
txxYkkOiqFCiDG3MpU+iobQVZDUIIRCamhXqx9cEcq+I/KEOkCyJTNBtTWRY
LW0IRSdOotWrAYbpedg2FF//74pnZ67ZZ0zsCzN6Ymk5Ua7Cv5/k1uJEXbvG
DOoBfizRZLptOAecbSghgc5D+RlEg65niuN5aD6+/txky23UwrHGvCvFO6g/
/b9RWtGzU+2Owvbazh5AlVnBj1m5PtHlSW0PrnX6uOxJz+iqv9XXrx23FIZG
3tQ0Hg19rRNDrqTSkm8Ep47p7lTon/9UHOnF5FQPuKQlLqpocQa2kr/DRsSR
jSQaX0GyUBNdIwT9zQldRDy+cg6TalJ7d/KCucrIHb1e3Jyihc5nezpSnNL6
zPChuM9im+eVTxo8usmWACkj3Zuk5ysKRUnDGCjViCkgnHQ2yg95B+7ePOVX
lqCbLcEGi1Av4cSSx632rELMtCzVWkTH1UnEI9zN0qhGkKT4pndREe2M7S9a
B7mqKP1TmiAZT6cQXQb2/IdE6AGr4X6bQSCpK2rLAjTCm+pBWh/WzPXWCwXf
LoLR7ShLGgg6Fe5YmQW5zaOv54xr02/B/+yLtQ0ZNkasUQnfaRt0iWja7+FU
5jHtR9CwUMCVCT/R5sH/CkHl+eJIrCIBJe9DnysHnMmZo8sxy3l7Jsky2zDK
Kx+kJH+aw9aluqAFOEKJ7OwQyNso+X8IerUVyaj6BBK0kyeec3W5nKIQrTZW
0ykpnIzGCgK18EslyFkIMPHc2t9PP9b9ipz2vws2f25vipohS43naWiwKnib
REMmwuYDS7+gDUEIq/Ngty3FBsrXepPVrJyac+5N/EjIHRJV8mKXIO538wop
f2S2zMH5QomsGuXU4QgrSpXTda8UHV22eV5BWPBZBm5u2Q24HOWZ09OT1lG3
qt8nz/fA+nNY5YlHRXLkkJCdyRhBuYTRBMHWp5EzE1uoXpnfY5bRuyiUcRqh
uxsD4FDvX00P9aOGz6y1Shd/Cu2WBNGzkLoSpV88m22tbP6yH/tujMiON8lH
urQv+AGPtYC2KuKZwgM/1cnQrkVyFsARRzQTRcVxbtkEkMFd6gYM3qJPtkG8
azaY7peGqFr6jwPz44+yv/8zulgQ393Pk0rIJHu20DPWNvTPRfiR2195u98X
JqF+og0DP3iXwWi+srZGQu4Qi2Xs0pySHShhR9bvBWr37LjTze+CSYraZ20S
f8uc7TO8c+xqkoIbbE9H3LfsI8RYTZMw7sV//sw1FYmg0h6O8Xe7+/o6sCsm
XiX7Oj85kMqm7vaJqDO7yRGxGPntFj5Uc1IznDSoCbG1fNQG3m1Y+4WYLoTL
vd+Hhb51wj+SaBu7ZbyxlPXHyYuV8nPlyCzbP7DcBtYPzeE8JmlZWJYQBkh/
5Aoc5R70hqZjoctcqzcAcBmmgcfB+mZnt7hQbmf1zWXoMSt5YIPWHKFUfm55
GOp0C7kR2ksmkD5tG/ZaNcntm2zdDUKbLhpmSolQr44M1YCveavoTqaClEay
DugCWQgtDZ0Q2UlR3z+FWOL41fsCnofRanaL7u/97/IlRv+t/VE5c3buoSU1
zOc/CNlDNQCwQtJ1Kf9F8vs4H7QN+Yfba8LC1qc/jHrOkT/wJ668UTPun7kb
UdNbug5A5EPx/nDFL8n3EOGoOt5BT0Ydz+GQm98bG5/atQNUYBZkCYDEvAKu
WzXvHp+LY0AmrE6Jr/ylCIjB3jvRK/l55mksa4/KVF57ebzGihUGiU7Nhw+J
QIqNDjygFWla5DoYplOeqjwAOUKkWJBu1wtCJNHIrP7gTwH2dMcdO/Ik8vDC
U/AmotUAI05FpDHDbwq+VOROnw2oRQit3LmhE4TgS1k7eRjKgCDo0OIhvuiz
boKRID9nqQmSMAs0Drg8B+chpjsOiWmgTO2FLwRxwkUmJ0PQRrHXXimlOvqU
tYGdtmChnftmsPhiZ9d1NDtg9u6NH2TG1b8III02+tXefyh+MtJ5BlUy/VyS
osCJV8zTmvgQi9IaiMeXR34M5ePElqtodFQ7R61JMcp8XUa7PzYNA+XgezJF
KWyUd5v2DM0gY+XyLd1cLc4GBiZBwsoT9sBRbQu5xBPu1sMhmwTmkbgPZ2P/
b0qZV2wvZyQPsDyiqHN99Akmsf4/ccKuIBVQAKYVGybNJs7F/9IDApsvBmKQ
H5Q+0wfgi86jBhblsyA3zXXTW6NAxV2zdpXS2wL23jCs2vnKDPcqtWaiK4bS
zWQdB8W7zaV4HNKIzAw/vSmkM0wNQ8Av9dH5qNIkSzFuJELFJmOcQFrkN3vq
t7KEz2XwILVnPKGf3NPAF6UIxhaoEYwY+slxwc8ubyYNSvKnUC9+RPLjUtaI
faIY1iDk5va3Qh5Pd9mH3QqD77vGax9VrlGyLt6nQh1c6inyHVcYYoqqUqK/
Oxl0YR7Jy+yH1NJSid7p5S9uXfXUVs5RcXCiqsfUnyu4vBn+jWSrs2shGLIv
2hKn2WjBg5m0TW1O6PBxbBXcVe2VhMACPCBGduzpPRwzaLmp/ixTxod+TkWV
8bW5QCjt7rNh3D70Mq0TrnHRVF9I78WL67/RUw4h2nE29xCDrURqZROpYd42
uaYyGxbm9MExWMqlbpp4oqR6A1UWgu1kr2xZmMZ3ptWqzqeTm0RovdBnZnMl
H7FK3FD+Hk1CabtvSrHEABqueRvSdSpih95VKysdaa3u+2Dr0KWfDHVRXR6b
78cD5wK4D+Ax+4QD6i02XnhT+kBnijcNJRzr84WWCd80JrSc1y+z607NDmIO
CLl97wYvrvmc3FSxgxjROIL0hqxsDZfcMBOlJu44N7PJtu/FdE9o2DBVWv6W
Wbw5GBhewN/wlqTBTAFQHojbcUnqn4OLpNgiZW10EZmvhAKP/D3JxhoaKgHT
xhIgozw6Gkfs5tV3bt8DN6QPiVThTEBU0gu6yYoHi3kqMJ01dZiaeiQ/d4A6
/BTjhtHg3/SdkHhsoQZ9SXqINQF42qYQzautmc3k6js1lvU6die471Xa2XX3
cHWEFaGstg7rsDIu7cO4j+FhcQZIsGYQBWgP4jHGE6jgOf6GRROR3HnhsPIe
ICzd7RpB0ZG0CNwrgj3qrAU8XVoxqm+jXbrgefh9j339w9KWu31BBRtOUClc
/36nsotMwgXiaadURlChs4sCyDtX4alnCuo1HlBgJpSOqdliUbzz+8xCzTDI
zR3FcDul7K9sUae2wyEVbwUnhepGHdwj8jeoj8AjXWqy5g0yi20b1WEdNO8S
CD+ZyyowZUmrk/lKF95yEfIly7oJBT1G3Djwn0gzjpk7agFMrwA5OE6q84X/
L1+mQgxfcM4ror3mhvBtSGaqY/53p/D29mC0jWESn0e37//UbIuyhXXWXsIp
3r/fqr2OOQWRqehWE6wrVCnRbGgAiCG0P3DqMoMQTI7gV3zniy5FLhaqU3HU
33YJhrAsp4Fzn1a6nMarWX4h+pu4RvPoqh/pozo/BOAscTXuZOSX2DSheU6a
8BTn9/RfQPM+qKrh2mEvSSrP+qR/BFd1zSmEBX1hdStiuKoJI2I6Fjd/Z7mT
ZfbCCIXCvoTTj8I/CczclCj8088LCUc+MTlUAaDFM8p1KXUZFhReRaPRNVym
DGrsBU3hK7cdb3qgJWljK3MgxraDA+fJV2JM5r16OzU99NRHZRncBK1FVrVA
QxS0V2ERtdhF8Vtc+IIjrNUVdpMlVO0htFb4XfRwNoM+f7vEVYiayRoTLQOT
4gKcbugafJZgA1iC0CsatMVJqOHSvA7sLb9n1KrT4ayNYxZIxb6LkHSWEs20
tIpnkiM8O7s/PQZaAwPExCTtKavAJbpGMW8XqGVDOk7EpNoE7zgAdrj73CHU
H7o9g5/A3iLk4PeWSlqb0ytE64iYkPTC5npT0kz5KMjcQsqziIiFuvp3ud3A
Kbu1u/d3H0syHZkuSl+KYdAzYBCNDzOcnzrNjeb37M6SaMmaOydvnTG9Z7OX
3+0rLiO76QAFeW+x1qa+qMD03zfOkLPng6AJS71AKxR9hCi6Y+rAcCB4gzRN
Gh01ZBvGxjD51gvnMCIrzQOYY/VblcbSWraUs9JcSE03Oe62K4hlYTm1ORhv
RYB01dQCN1fj0/Uv9bMXSiHtKGo/OWdn/YAKKqaBq1KAL3jbL9nLbeCGBOho
d3h2dDLuVwOo0a3kwhf3GT60oSVmYxomxFbD9xZADC45ktDnPMLoA8P7W5FO
AuJGi/V8hwwvWX/6RmaUsehC2DbRcKEOZrsGS+vry7sRYI/YwuR6x3ggWQeM
KTezdqA2uoMhJ+J4HmIOUtyF05zki18oPJtOuhkOrz7UmVQn1qtL+/zlbDPz
87pyp7hm/bCsFY7qRarlw1ht5Hl4MUcMMCjgxdfOSrG6h+XLqCcqsMDeuGB9
L0Eo2tvigKYISnZCd8PI3Iz6U9F6Ct5BgAJbjHkzOE0IA8IQCNb5XldAnPcD
eBBk7a3C5MrJl3tHGUpBkhNqtwqwOkZc8CPcpV0GczoiyXLsB7Fbv2LLCbR3
14HhTHNDDuyYAUbIcBeeGF7CT4XpJMbK76vYxqXGFspqMjxjEayDbD4MkmDz
O7dALEdxooTIac/OUHxeOk5Rpow0vAGtZSNA57OkNZgW4fzpJYjh1yepatlK
60cgefv+yK6INZ/bOpmEOoQR8ne6HEROIzDDK1E+0i2thI3IeV7ySFeqEBP9
l+33vR+XbuxuomOqC5Orf5xczUI9/9TtGm9srT6AeHaxL3OG2nfTh+F5xexn
OEU2/dE4RHrhBQcihBvZNM1JqQ/oM4s2FTwIPihMUMZ0xRT+Ji2/96tkMjJK
dc4Ldvb0+mXgpi+VlKe7Klln527M774+Yky3L1c/m8MQrw4PqGodItLV2ibk
MUJGFvdWUWbwG9/S6hjO/+nDHjc4zO/9NHR5Gr+YJCiipxSWal22K3smUrKM
MHSftAMJmNQc2s/sS7MW0fxI2RRN6wxZ7aVj2xkklRLbcK8t110su2fDyNQd
PxsAu3fOhnkPCs1isqSwzUPyCERg/zszSvjt0VeIHkVqvNOvrEeQ02BOo2ob
6Urh+RUO1zmvb7b1bFXuXaVNspWjeUHMYFeM2jwrcOTADJEMZJwrPway6Oex
//CjoCFxDcgcu2p4O+Hxv+/uixaYb2Zuhf2vMleqRyn5UdYo3ehKPfafyAsi
oCDSkj67AizihfTsiProAuZOZW1gdroU25mwfskIev9picZ5jCNUD195bjGM
FjMwnmtkIFZy3ylkUwjM6IZmZrBUUox7boo8ivgKFZW6at1HR6FdSxdg8isC
2MT8notZfNQTobXFsnwmF/CMvjSzKdb529oyyCLvDW7T2gV9/ysdRIImdvxb
cJaqjO+Q7PkeGeCcInRMMdqDhqaGBf5b/3OXN07nxmj+ewcGP6syfW2MGsDj
6WLkw4+wkH/6JevNLSJOGMyAEPkY+X+t4y8IF6ahuIpryP6k/FQ1XDgcbmmz
7i587ULbT16k3JnD36PWb1I3F8k68pwwP5ASK2iX/QhQtLAooUAsC/h9prR+
p4f9ECFYZVk+kdmb86yiTbd+pg6rTipCC1MDoOe7HI2tSw9stTdDiBCbL4Fj
7Mg3DBBk6Nxx6KvArjIXB04vNIFwxRncX5BJ6mrsUWkwJnt2inp3R6KxMx2U
oHQHQ4afdfIYLUjVPkLneqFUX7mY4EIH300rRDpXNEqdcLcNfwYZqrBscKlR
70oMSsEa0qCGoz7v6nO42bg2LDhgjxhP2JhS+W1cvYFviHapzV5PiwfUdwQd
RZ8zTCHBsXdircp1ceHnpf8b3A3ifWxzEITV2gbKWgg6FbpksVcPk9/mJzYW
8UbwxG0hxZJg1X6JKUUZb2CoTrmS9QQrodIqnTJWhke3Q9T95NVfsSo9FNM3
wluDuRiU8gKxh4GbFiw0pr329D/NxDosHtBDB5RFJeojpp55HhY1VKWrUCJR
w25yHi2nqyPevKFrn2qcc4TifqrpzOuR+v0uf1vTb3jqzyRTjT/TsJYkid0Y
XyKJNQtNFo8U6GLCLCMJMgRyw3YxS1CzS1rykXboHB7erPhxff/YGHJS/Gx8
DXZX+75Km1qpXrNNLbeCTPDwu64v01/MOs1qnPDes91hgkw/Y4UjW8CPYWv9
fNCz5wOaigwUcH0h672ML5m7q1f3x9RjQFzQejuzCsR0MQiOWmFDDrxCDTK9
ngCSfd/KpvMXGCLxVChJAJBcbsBxUaNfVwaYUW4HHUrXvnHlSTEs0amDmiKo
1wIuCdO1Sfjc82Rhh42OdoHP/O4MIRwlzgZdP885RVHt3mHvThZHS1kEjE8/
tEhenZA461EtT67qmVVE9cG8RDMYUQ4VK6yI5iUf7eAvHCaWTiKJmwvmusdt
wIlAuMfQDgO4OJgX+L2p18yzm7csLqNd1MZFflZCGc/4xLvCzDNHcJovPsRx
LnCw9bbqzIE6/TAbcQv28aCL/wVKyVdZfOUPRZ71Frgg2VwubvjHq6/zgvGm
Lv2bKMragovgT0Im33jUJ29ClphQ+gGq/BE4+M2C23V+B5/u4iZh0CVMixFD
sF58Dicoa5w/6kFp2a3OVQtYV1kLAS7L4ZPuJLnbbx05TipRRMAWA5tbC2MZ
ioA+SfbWrhAvrL/Y56P/O30bJQRtBhe8dYkz9XKfgkgn8WEJFI7irkfMW57J
U/2zkMgBsBnY+wqK0ju2z8fG0xEIfgex75PFu1XXHKp2yupj6SM5eNc0AOCc
8gkWjN87EtEJz8z4q5EAydMMzeIwjrgoxp+O1IlNvZeLYcU4s06mqJorpwbb
yPnuk3Qz+e8rjtcrfz+RUtpMPJTyBKHvoWOmbDMTZH2dBLp6XNMrmgbW736t
dizow5x15YqjJpXsqwdIhlfzFU+fTjJQNf5p/ZodfZOUAFKFGEUX5aonS3wL
22yy7X4FXa+/q4CtRhs7THtskoJkFjxSiD3FI1BVgQKdi8lpv26+NU66l9Xa
5DdDmjMLG2KK2J++yj/JoIJlh5PHtDDErV25ZdVz1Y5g23se9nst87HxyJSS
SjFyEHrB//Wf0CKiV9PT3hj8jDBXjOji2H+56F61z34N9HJQJALsGSBnCryb
fvyAxCBdyc1DF/4lU2BbfVTfYMG0SjF8smMXWeRda3lNnUDuUGya3EIk3/v8
GdkSzcNVdYPlZos3r6BVdYrtvJf84Dy+1sxYuV3QQ5rsZq9Brc+pP53lLHZo
AZGUBqNK6gYqxmJuwv1e0rcfj2bgRs2VRMiQIoCbG2zbgClrB1KbalkaoDlY
/XfhAuZ85uZU43FZBeDAct71PLng3oCptbw1Wi9GZImq/wdeZ73xxqq9elce
kfJq06ViJAxC423evaxiGH0+j3a98A/+dtxqIfw8iz3aiI1vOLYyryMhWo3+
mPlIZtI2a5PPv5aoadI42/g6gfOdwG9w+AKWn7pLLffg+lnMuZu82F2eo8et
KEqbcavPbIpjawIwTqSyydquwoopuikehVwH2uX/Mz7fXeSWA6vCT9tUR9Z7
xP9bfi1awMqeBttqv0s4wxcu2vivjbcaokXqp5BXnLs+nVG4+UntSPrxtLNP
6cGzYGDvnMTPtP997TutimJ4BqwZe7mJxsU6veZwukAjR8UEylvra2+TKHx6
H2v+fnam9hl9lEkX7ABUt1Kvp+/VErfrFmPLFaTYNvHAxjMfdERguecYd2y9
obVTNkjX/SBSnbFmk2FgJuPAEU7M5vRdl653tE+dRR7nEbHzAS4q36s6FzX4
a2ryptdMDxyhgEDTXR4S58K7kXcteyuxF765yGeTAJT/SmxnkcvzhgYyyBDd
owWpAVaOXkwGZBxPQa9eHnTy/Phx4IYU0byTLrV5Ug4MP3FKwsHNkCJYy2qV
NQDlC6/9wHn1OkjsWx1ZzWM6cvNksz1Z02IU9FyHz5A7kGHHkfHLAxQ8KXsG
TuPzcAKqSOwQ1sEO/8I2mUqi+zPH7tJKg+09noVYZAsmrBQfbtWkOOd/yodR
AzthMwSEep92C3xxBJ/4ZS6ujA4n9oK6/x1RnlaFIjuCHDEJ6GxfFz9askR+
SnPWZTpffNryXsJCo6JrXIXeXJN0LNFjx0dCxSL5Q7ZzRhUWxbNiF9IKYbYv
o2dprN3L4MPmx/Zrgx8pc/i1LdSqntCVCtie8VQPgnhYXEk+f1b6rMIBgkOm
ZHafTHb6SV9fHkaNckcm5DoqpC8NgPpu7SYA/ov9FVFwmcr4pFl2qSmB7EWx
dEl5T41N9ED/+j/Itoh3xGBhLg89qDbNrVK6fmA+GJC+XAZ9JHLt0JoqBGDe
imrU4uIS7TA9fCbDfVcC0G9edboRiJu2gBUBB7jpCGmCcjEhscntFy2bveQp
TEUKxNIAPIYUBNZ0epDTfSBqJokdCt1mm+YDKbPCo+DjW1fW5RX/hLN0Gsi7
+gS12C/HYCg0C5yPhMWOPxQqrLmlt+XsPz+j4BG1NerywbsKLDX9otk1UWpH
qeQIBq25XXNfOISk+wh3x9clXkStr3rjBoVfPXWoOVENdWFoulYSdX9+Gnz3
aI+LdTj+osnfK0i8FnVyKLRA2iPmpHcFPrBR75peztnK4tdjfkRPvrmr69RD
o3w9IvAAzC+o1VJ/g54GEyy5I3U24aILtSu3Hch2gOA/pjXnnGqcSK/VzKYC
q7jdLhYZCzXT+jFy/vSUI/IN+Z9gudaXjcgVVFPe/wpkH1xL96pAPPifxtVZ
RVygxnPFV2ZlLXcuDZuDBxlhoAKjelqvVAYsEukzpi+K7gA4p5nEgA5In+Gg
2EHVMvXmaEmgswr3hOxjssJtbhS66BeSBRQjTHG5qNifbtNnN/B1wjwuobdf
z8zb+8bC3sN50UGwQEu3EfGLm+msz7CJaUbI7NQMe6jVMcIhD1N/RMJqTm83
KRs1Il5A6ERZbyYKeXNScWtyxveNVLgnxb8UI6ABxs4YynMybetXagAL4oDG
YWMwbCOV69nN0q/Wl7wPTEecsKz7sLhRr/N9E0+Smmn594Og1MCyH/tcwBm9
NZcSj5clPVJl+LBw3dKHJ0gDWvno+z2FyaPJBK8vskRNXkqgZZEJu3ECkMRX
sXChDJVDOqgy5d5g98fwN5bjHysFXXhJE0X9WmCpKKxMg1yMCwJ9071B8lPj
Hzeq3SSTOzFspXd897JP36rEH4WpWEFg9F4Z6RuciGgbjAKrwMWzGT3DwLyP
AGDQFpekLstz+olbD5CuusTTyWC5JeXsSAVT7VJByWED83AJ44UaGSpepbxe
6UKl4IeLWfGuy918gwcqobQZFMzIkk1wvA+lexf+6icWPaaeF+7U23PouYW8
9FnTXPX1ZIMI0TeIceupfmO3XTSj3ZDk1ByF8QEGqUfMoHIIzWEkmFxCvXtD
Rxrg3/Giln6sB/F0PqrlWThmtqWtiirki6LW6lwuEbD5rCm09GPhEslZ78Jy
cslMWJpX274U3zhKc2W3VXAgyPWb4KRPrypwBRwub9nRUhR4Zqn60xgnNaIC
NZX0Dx3+jo0OBqWaMnFhgLziVzxYfNcpzoWCQ1XNsVZN8Saji9S4AfDgqM3Z
+pCYhPDiPPlh3+yuY08Y1E3iKj8ZONk/x1NzSCwSYkQe1BeN1D9M+PXCJPMh
QI8q3u+nxo/vZTzy0DJl8fJ/zP7HsrpTH7rZjZ+TA7xQVGpeHHrhpHUKxBf3
CcIrHNsg2HcWKUjiSL2uv/eVhPWDkaJH08C5pIZgc8wwFEtpSzVD+xI5j01b
l7DVhQBeK5l4mmJN8joUS9R+brCG7G99ZpxAw7lEcJYuchFJDeEF91m8+mKW
kWg7oRpkhv9atipIeYL1oi3tHvahLw3lCzjQ3dlh/ZqcVUVZNSfi9xnTRfPB
jF3fK5lLKOfsq9GosG1qjEXFpShoMgD1U4+Bi0D3PkbCaokOJjORLTjdKzCl
aFFtSridCxLEPLEqXI293elNjC7Vse7vMzr2KcrAtCYpJHgsPAknEKQjjw9E
jUQuZ3l5tNmFuJ+CKld3uARQhkk1yeIsxkvWpt85EkuCEVLcN6garQopCvo7
pBPaGevOxYXoBUbjSqMQ10eTArzJs6e9MnJ9MCKRkEpFAT5cFzwWCyrPLr02
BwHRLxhyAYnBloth6TaV4J4Sx4iH2SLMP1sMbviIUTZQxqDguzaQgoBvnOTq
WWGLKVMfCMhWu3PtxMn5OXe+1PjwwjP2Di9l0JQryHgBTWAmBYOW4lp3sBRW
M1cahhi+YwHukFExhVbDFLLgDPDI9kNTX4otYLSVgy4DcWmQy4CoWzZXDJ4F
JXD55WY/gtZi8R6wWA8nlFcaMz6yaQWmpuqBab0+VOsUXoQAUR1sjK3PPijG
7KAckzvDW6IIFEVt4dAmOA4bJkZCMdilip8CPbjAOlRWXgnlxvaUFZm/G4JU
RH897/kTsOZjpGRjte5QpPXSF5S9g5u2xRNc4Ml9HjxOXlbOvj9W1TMf8djf
JZh9Lzlw04kPvvOFByFaLtmdjCdmC6anFoJ4wvYmoPk/X40c3rO+sxwcHuVx
JnQWr+yfatj3uuCH+Kzqm7K/60gfbCi0JhHPHrnhESn44eNNvQxgQxu+0Gwz
z8jYG9jgTmtAg9X43nIeybZYmnfM4O2P5z+hD2fNk2htBn2+9NRgaudwNgCh
fAA80bNQOFz9LiDAW6jphA0tFzzUtUBxZBW8z7pJLDHOBm4LV5Rq0KdtlgKe
tWaSAEn6Hh4juTXqJPplYpbg81CMU4xNFtj5wnyb6yJmdm7MA2jIsf5xSaIt
5xFMl7deEAZyaFMMTCQeaZZ+rRjmie4Dc2yq5SFyvVD+vGNT0AEmyP2SirU/
DWR98engsRn3eupsspuK2l6ozGsFvJzssNtlFFXIfEUY/IQ1e8x8OMOhgkoJ
VjaWBpWoNAgPnrYhMdKKzRJRL1i9IGoeo6FEzDgXAVtGI3q5/RTQQwyqFlJ7
/UiwO/KXYDphugvtlQybHBjBtjHKn9oVIrpz0rAvW96VOCOkc2aV33zdIS5o
ayZiBM8gCNG+RfDOFTQ8X1RFxXF6A6Qf8xxSKIxOzXZOa0UK6zgPQ6ME7Uck
3Q8NIR45YE7YYsq5LiMCewvtTx3QObnvPYRWL30ERzjnImCIHnKX4DVo57RQ
6nV6IU3/hcFAq9mSlf7hHqs4DJYSaD+T0XL4VdNAkpaElXKzDpYxwoNTPyvL
MeCbXeL2bXO1IhEG3qi65EIEWLBwOw4lGGpDJa9+zXWPia9wkfcNSXN7xVGS
APoRptGzyeiH82YgSEso6rDQCtrMeciaY5i3NMaLc1Z/PTPT7x42Jb++VY+L
PMjDCSUDmItOge5mJUIh7FVqlQJPmDGY8995PU1ZjXWR+wqDfcHM4rNGIHpX
adlwmrA/NP0jr1o0ldjBOFbeHQRTzRwhYGJxjjeqcsK3e1oJ6ExEqlKYB+7v
XkMMn/L1xaz94hxpAmLTUUDLE+vr5RGCjb4pc4q5A8xxFx3oMFiDDAmqBf8l
WO2XF3thK6UBukJ7a416IA3MPimXctpiNJFs+OZsde5KmVybHP8C0bU7WGHt
tW8/t/B+lDXbdw9T/jOk/QCTLXc+QMPuN4IG+/PqiCjs/irr9Vg/pwIZvxV5
Lv9EC3QopVHAZRA/AMdyXgzNhID7nqBQwuRQYAeus4DqUaDrsCwm04BpahEp
DuVtDja8IxQY7IYm7vtjBNVd/43VebcOYbrfwK/gceenXvgU8PA6TZtZsW0C
3MQWu2775aNLtkgyp2HcY/5XPq4xzCsi6WzXyyGdxRgihPKMaYIY6hSwsycp
PMmknkxdAI6WW4z1RlwW01AaeVgvoRLVll+XQkwx9lyJoLXJieoe81Cq58dr
oGMVmO3hA9x/fHopqEftWYZL0DXXGybh+aTNJqrHFd2fzXdgm2hEzNO6Ltg3
QPbYsgRbH+6642FcTTd5V5wIiF+ln1RPXKkUyCff6HVbHTW3925Fpp+U9L0I
HxynMYqTBt9r0itZ73oMeyIQcttQgqsHgBOR1W4+aHadnXKm6xN3n/n/Ikjk
WTL5fQWDQWXW/fRt0y55fP5vlYwev79I7Cxf6TeXfX7ywZKV3Nm+8SHZ04TG
d0IoNzHG0T/Itp3aFNylG9VhiPgsbzTL0kCaJ9BhqWGXaCq18YhIECwUDi7m
LdnbrU2fQqan3ZBCvS1WLl0ZUstE6kzBiRb121hPf8hERrdvAapapJdITP6x
XOKe2Su/FQaqDwSH59bu9B+z3+wsCX4pj8g8ZjYysBARtN/tdBpoz8ND2tnf
voLt8b1CDLfM8fbuTquu9cJ+0IhTvPYkFjHdRV8LdZYIu8Bl/+B12Pe/BiMB
IFKPQotbDiecAe8NYlh+JO3BUSdJmZN7H/O+eOkTsG6T8BQ/MFrc/cDBMegF
N480O2XpaIMSsRlYlfS6/6xJCIQoMYncUgidJEnpGrEsfWyBAb8z0edtPg66
3H0IqkRAYhoflP2bUMu1fWajo+S0Zz3MR3fz8NKH8fOp33iJvAriUrH4t9N9
9USgiB4aPpI/SPfDNMCEeoTV87ofxoNZZL463ekigKVAKqdp5PJuRoeqbpnH
Jztgmnl986hwkeQAWT5kO7BBpscqImdo394ZWFYRytTtoqsXfK59DBctAMCb
iPnNsTFrbYr9McT+lEMHiuuP6ygDXYccDyrfjwY4+0+vqYvHpaFCu1wd/lfn
KrcKacSLLTnq5YS8fgsQRCv/y8gEi14yfRSIoT2O/TlZNSJhfyGAA7mieEjg
Sgbnbbx4RKFeRMMTmzAu7PByq2Qm2XqkfaLepH1nw63suEw9Mcuxo8eKpqG7
B1emQYAy3CPupivGPDA3m0xzX1KHs9Ydjimrtf8Qbv9CjtCnfrIwkvbrlOOq
e5sRTpqM+5D6Br6t2TucacZvyhCSfITLHDeY9rR3iLSlPoCIIWzmgEpz/xzR
GS4uEvGRDf37xik65CI04CtlNjfQAGRxO2Skxy8Wb6qG2jASsaAhVb+ZEX2B
hks3ywiS3KvX9oMqE6jRHTHxuDDsx97Ux2/jJkHLnSbrNMbLjDy+DnIM2YRJ
V4bEGgghVBGjKYgN8aBcMYo1244l9FIougXJ5Hg5ESWdfLXZLQQjwiEkOaR5
NsdEexG1OWFsY1cz7qJwFumCRk+459cwwlO/xJ+QjuJRW8VhL3OObAl8FPkN
VAk6QNQ2j8ln42YoSeCv1GbalbKt/0OKkvaRLMMkqxNy+C/1gDknc60DqCHY
Dd5qGxqSU27wtAOQ7JzXet+wTE5csd5k8pG5R/5zJ/ZT3VhY1gsQf7o9k+o2
SEO2jTbv25CNPIxIvm13gmRrv8fMiz2xXUC2AenH46/z2p5NUp97f8Gyor/J
CDW1e7Ae/kHok/YApJ32Eo6vth1oXZU8pH/G3NR8f23X5IgibdtKhQiN8Lim
HCV4/TLjBzs8dpd8JtH0HJidjlXIF5YJ7hPgQpqYYwcsCdbdvCqin++P6SuT
xlOSrb9F/xm9f1wOp9ghHvuRIzw9o+ZM8vhMZMxpw74CdyRLBLrPGrMvSKPk
x0ISueZiG+Hac6wHI4YIGRVFI7YQypf5qVigXrOxe91kUyr77qxm466Rth6X
9zkUmhPw0coFAs126EEXYEaFC6u5tgR91ivamim8kp52fihM5ifg/n0kolIE
apqm86IH9CF/woTYNVzfChz+QsMOqazeVnVLD1bYtLiYFe5dqngXwf1uK4Uq
MOGtBvSc2XIc2ymHch3od9SxaDNugwN771WEuK+sav8pLv3OhSXeI0+NY6kw
34T5AyxE2vo5wJ+GWVsdlDkSYzPVtjvLdIUf2AyPnKsyYuYujK+aK4/w5DWV
TxaA27rbgmMhypOEOlayAcLS+nvJ2CSnSCULTd/1hX9HcXYJCu4dYe3Tnue3
S8iiPqxnWbAE6p2OWA4UuVmd2CfkhgcAzcs8yJT3ZSwe8skWceKyNinEdVLh
r+9DZzg0baDesZXK7f6aiPbLM+b6/4oYjdpDAVeMiEKCKOtGxBoqcihB9M+v
E/m54og627fsIsd6yq/HIOo+mFW/mDvQayGf4w+s8pU01MtaThQ0awom+pJJ
mnd7AypCN9qJ23XXvlU43lt8ZfIZGorO87KMm0XEXObx0syKHMeF541EtmdD
7YxBXthway49Vx/vgxHdFnNh4kkKLr9F9RqBlREh6KzBL+2wBUEbzG1MYBSv
DYHyyz9PgVNNOldY6d6PpVGLcp/9vTul5gpmWScPZpMLvrnL7C09riyRABAZ
Thl2wJvJTgVMeTKVo1wBm/ON9ty18v9u09WwhGySf8dy2kYr5VWxepIr7Xaf
EAVw5IUmPIwJHj9Al3Pe77qDeTid8Nt6NkCUWe0BTB0sASdiwre0LrAkM87t
U2VnCyXyjEBjQiHD0CQ0NVixUA/5/JSk4TBDJd+3o4XZa4dhweWdoUTpfPBQ
Q1LVMssFPzTynakjhesNMyp8aj29Tw7BsxBAd/KwtuWu41llUyHN8HL5jVV3
bkFczO4/oOIBp4fX0d+ebkt/PjNb0uwVDb7WTNV0LcXDxhT1Rfw8MzE3SVKe
NPE5B9DxWe6H9WnWD4N42nA94VESPmhNzlKE8RJX0/7PUuWohiPYAus4Aa7g
PH00w6n3zeIva0sg7QRQzBlWYTOMR28x/jowTuCWC2kDfv1q14bVjonkAshq
u8Va3WhySsrZsKXRBAKRwBB8QEa46sxPwRgZpIyQEaSFygy9B8vSAHV56b98
eCk/FWRAWevFBzN2756aSIlhfW0qi+3hCpoT/SYAHYOU5c8X7lN+mvHH8SoL
PQl0FZMShum52DTb2y7BmeXn9RKWeXb9JRmkopCeogLGfhpHkXKepiJpGizU
sJk+aaG4OL7ZFF2OgTnQhzNdYKsxJzsjxPwQVfPO/prYFFNitOEIzh6BCL45
5U0iebZZ9XmvSR7j4tbvxBS2MzjjEwUnhGSWwAotsdKySiwJ9GOUL7JrD+mj
oygDKBzyjaA0Aa5hDfeT+Y8pQiipmT0lF7QkTR9A0TP8wOmpmMBVE/Z9p9iE
/JqA8jwEHNbtFj+owNH7Omh28T1nHyaAXeEvU0q9ceTlTNci3LRP6mOBx/Bb
xW1LlOAl7za1JxIqwTiE7YXYLWvynVzPSZQUGh2EK2Imw658Q5x4b1xmhy4m
+kNrJAbFTKxq5IXXEja3NPIVM5kehKwbba2eDCB7pPlJO6W0b0pTpblIzOrj
qj0VdEGPqOjR6x1Qn0JMQmdLWQvD7qG2Nxkiq1rPb/X5ZI3C9dvhcVE4xl6q
IYEY11aJJnGG4VDWj3RkSLWEDAhYRwurR3dX3vswIvZ1lhkTghmvdTJqoUk3
C4Viuz0rShIQmGoG4JpVWyLi5gtUFWsmH6/ZbtPzPVtIfTAV4x5QnNbnEmLn
B+T4H96L/djmun+Nl2oKjy8IoRrQ4Vgfzahoyt6WCXzztbcdA1/W0LGnxiGT
GqkpKDLcySoaqruV9Z7hg8MuXZDqYwOjeFjIQS2yXkF2xoIY8fKwjfntxpM+
3LStwfp+62duxA/mSLCe+u9NjwIfw/kpJIHW0LuS6wF4OrgI0JcAqu1wTnI/
dSeZHdo+jLJjbM6xsye800BM8YxhH9+q6x/1VDyC+67EazFLbYJiMue6pfdA
pQ73rPnPvRoIGVfjJ5vfdXuzl7uByf8zQwGFieumcDxbltWHe0IsHZbOk6jg
xl9gJQb40tTu3EROrL93faJ5RXFzWZSg0P1Xe3H8aHSAr6kn7+66MbCGjEi8
DUjinJc7g4zsUl8emauCih7kF2cpzwuDelvgp92HeANJLPTg2mbIUSyUflPb
isVxa/q2ed+SHKaChj9DBW81f23B8icASXOZsh+988rRedI58bBG4qy2Tdg+
3HX5Im9BI1j0rP6RsRd3LK1zcJvjkWat+VZ4kRombbg+iIENu73fSpczAqY3
iEfcvmMqcLYR5csR4F5fD+8XkCz10P8oyEAYe5BkcHMYwhVtkjc5vzpS1ZcG
DnadXHojAnBom3c/fAGc+yhwpBQlijLZ8BVEQ2oBaRVrtze/g8YFj3xvMYry
EXhE0RsOZ0UXqxHaGtwVxY4SiMXvr6VdZP/jTKqpTFbnkqzp7J+TDVefnB+1
O6BgM2qRQIj8AdTOpfQ6YpGAGYgNGd2oiFhndZQxFxLflyQKdONgCqtriUOs
Dco42hCbkIUFp4sBW6InVctjYqVzdN2BAxCekdWpiu/RFmf3FtWTXaGx0WJT
1vZSiYY/Vc/1LFLSaXhLa+621tQ+klvaNnNOBua5g7q+YSUDi3COgWWnkVjI
ulgNu4aeLrmorjI54iLmzB8IzenQcz+xe2Tt/HCS0M1HzYngY5MqAQFfbiOk
rawG1klVZaH1Msdk/ojwgo6FoJ0VH56gYK2jxg/wk4UkEzyZil6Ly+TNAX3/
E8RurKtdEZjL0f5JG8l+MpGWWkMkrT0B9yRqNA21RCf5zuqmHHPdCujpmC6b
+AYChENr8LPLqDDRhQIAWaAh+4473Mg5sAFnnzznZGt9FO7km1F7z2xR8xWf
bJ1DRze/pmm4skbbGvwa3ycH3wnadvOSHMIexpSf1uipvqSWE/saMYscqbx6
sFwwdRPv3hhvvcbJ2k7E4AdLsbnAr2Fv4oPxxniMKAKQjCzqRNrdDwiAKtM6
rOszNkGvOogkTcS2e1pB3rukdovS+npmGfu/mmIMzxy4ZtHlSy5a1eK9pqGs
vRjgvr8YdLlcCL4KGOWHF3IHdLf85ySMt/XFzV1WNQdBJteZalvS0lAf5aLy
p6pEfz0HZf7LkbGEGQLi/AwaFs5/2jCjh8y4T/Sezm7njLrJgvvebm+ABHPD
TDmCRBfPOpfNzFNdYuWbozliPpSwfzFI7Y7nqnee0FEG1WuL16RlhzJOYPve
mbHHg4iIbSIeaKK/qJDt2lAjCndYp/vaMq2M1PcjG1ER65faJSBvPoqcQuu9
a1pS/cQL4Ji7CMhu8dxKTL21AjROS0sFw6jr+Zl19nD8GAkZT4uI+vNR5R87
0iy1NKzc3gxee6CqMWodj847vhE2RXmnveKgZS73Iti4LzCkOELL0KzTGWrH
/cvNSX179sTvkTTDAZy7l6TmWqKrNmlDvd7IBDuAGkYbAMY2FHKqAnPrQ7xa
59oYVq3SZM74F1XQeioA014e0c/QnrjI+aWL0SuO+w2/Dlm+wGyYQy2zPi0m
lBH85r0TDVJaX/esRtKvCxR36eJ34fV7M1rYCCngD+M5Z8PoDXypBilrIqjX
kxB4ftTkcuXZC9xpn2KuGZyBV7oOStjHsfQ6lhnU8LT3Dws0Ub5gZINHydRk
gslTg6ea2hp8jOMbefx9snMveYsMpJUvW+rbEIcTTaIermbch/5VL14wvjaR
zF7+ThDaAkAyp8ij4ZNDBEevsPxdE/jHMm3YXQly+T4vWz5LGTQttmpt0Kfp
15EkFlGoQuLJEMYnx85VDzWM+B9SoUiphnKQT5N08WB5vHddBVD7m+fPyDRd
I+OjurERnY4fkhuH2IR7bQ86VmIoJy1n3ZfY/v4a1Jsw3oCy1ytEvZ2pbBkT
j88+Pc38QWp6Y0BExLMmu+F0A+0UJy6WUMnq0U9dQBbewjez81Ino22YOKNE
dRDTdZohAmlp+5fmI37BonWGnpnKKD/a7/S6LA8+sZR71mlnqncDMVPOZawf
hTSmYbkVOGa//C3FndtoDFMN9QmW6sP28C4ppJuTEWsy3hMBuGdf4dcNa3PQ
57lVLqvjX5vNF0202XqEY3VnMWuvy/fa4m0WN/pvGtt6L67kbLFvn4moVt6L
J3m1gr6T5vwXEZb+xY+ljxW9plQOWV4dmxcQpnU3Ky8qmPS6mTd6mo2oCMlb
e7A6V9Xy6nPgPVUskdro9xDHCo6vHpFOaxmqQ7sZCqd6mGyGqxV7grbMyqKq
s4BrUwzuiqybwdkBexNOs1U/Wq+Bo29TTOwgE7t6uI8tLh2sXs+dJaaaNMxv
0AUgyGcogUzXfxytweGycpO1xzceylN1Cf3s9Z/AC1w7n8tbhzFobNoUC4SB
riCo4weUB1K+E4qjR0ghwniDqGtwKSoPF8bCohVws8gqoaNAR5RLp1WpElMV
rDCOh2gfi4uqga7AbrNQqsY0mztdU5uAQaY8ZQGXc8m4TnP844pyO86TOtNN
ZZcxBgSFnoosTVCp3BUn1++ufsAwQS66qFYHWwirZTiorXlSQSm2X+opqj+D
y5q/C/KWWKIPTxEfNOSZg8J2tCdpcx9wL9h9zpuIgX7QVBei2PRfPfUVYY4a
6OOiUYH4bJfz+IkboyTLgyB1JCk8aS++DspZLgLWzaXU6Gc3EgDm4jL9y1li
dHlvOx/g1E2mIrEptAR5W/gAGJOHxagEOoVi+TuN/1fRPYB9vcj1/RktkjRR
XrMncj2UiKNHNwMzg8NPJIQK+UFCZM6yeqKGMD6rCePVpuHG1XGrpY5ptBD8
GIWo9seihmTQkGcZDuC5dnt/A1wpm/vgbOEZFBjRkjNnvZfWYrnKktB+22Bg
uRNJdtF+zUge2a9qKgOHA8NtYeSi6H9GPXRivMA9w6Lu16QeH0FBs6cis+kn
3yUMn/R5ukIUsfQe9bitIu8wuhSx/j83pSVVrwX3VRtd6LkYeMXLAFczK/Sn
SS57P4Dd+fpA2r29w0szGEXeMKzKwvHTt0cFJa0tgaIFHQzrKB/LFGqi6ww4
q4+12/6sWvIt/INZRJ2dZ3cQdh6mdUVUo/tJMFvE81FkT5tOcl9q7fRTBq2b
isim2LtSQZluz/9gyonl012f6dHbO9xobb19bJeH+LVsdvIIEsT/2Bs6Uyl4
iuVcAvM8IIBYeqmjU71FkNVhsZXVRa/5pRQsTZNUe/exgdZDqe1sA+PNcXNa
g6r/fPYTIUpFv3R0qnP8PhP5L6cBkjaTHhGLMnRD1Ulj8qx6EFzelWps21PH
rxjUZ138NN35MFWnVgBCxIVQEq1xIt1/DoVdm2yJxH42f92AT1moO/nvfvJP
llaDVeDUPekS0qNJwejBfXOR5wP25NOzzK20gkslcmQv6YeGYG0b0tCSh7KU
3zENZI1HWoWU6G8BPHx+3nE1cei9OIa1NZpJnRF0G4RlDO3Ag0tYYuMQZ0u1
XvYB41GsZ/9eGfa4D+Do0Yj5SJzq26i+RuBge0yZ5DLWtDXG1zrDCKxl9SJL
DN7Mv535EO/nO9c7OpdGro4TVfbw4Wx8vJYetNsHRHvgxgYKKlTpF5zqMRac
oUlInNfM4er/GO3rVlPpRsb1NEDiVU0L+SSOEFIMaYbntiOhmeCv0jCGnQrv
UYtRgkjqEaJ2hKBREU0k4aD/OUZFMVcdta9kYg/MKrbU8E/BZx4RtnW2qbuK
Hnf++QMKF1RS0eEWdUKZ6Z5j7EBIm+rM1stp9KFWEOQamunzswMtnUHJ7bie
cIC/hToX9qZTnDlJWUTXhntm6y/SLteE9dPkxwY7CepS75hpx/hgYzOK8LmH
GlfLWJ+Cl5ih2swItZFAY0Rv7vhPfOJSbUaz4alNapDNfl4/mPrE4v0LkfgU
/TcbziXW/k0eQySbpGlsIbhqGGPJakKqWUkpJjjD2OAvP5TBfGhETPuGPF77
jWflgqF43TOAQXrnRQF2+RP3PQmCjo2vbe3/eT/s0ucAC4IvN4vZ+JiuvOye
1N5HJsqEElm23WtApyWB3wqDYh35vzSidDzyJDm9x08a1UkMxpaP8PnBVArn
Hs/D3ao/30dlQn94/VJglZdj07I9PFfN0vmLoAv7GOTGB1KWUikPCPswWbgF
1PjXFmF/uV5DzQEgHCsjrMVdV8zg8ejT2aSaXDPdOocmdo0dYHNTo0h9e+5F
b5srpebgLKNjGHrUknjVkk5Oxob+elQxIdhkBJXIV5MSY8VvKWAaVaRa+7CQ
+8fxksT3EEvMCecUCuYjyoOdE8G1tdtfAvZkh3YCTCaQ0W2ySzioPkObUp5L
V/S4xWWZUEvJxN2qaUJZNwpdlNPImP6u+nt4sXzb0j8tWWu5XnWgdMq/jizD
xMGqYooonMXgnclZH9BwY16beKlv7RUe3B+WomLpybCPSudCraTFYDdXZibs
iEBJur43ex4taqn8cEWQKbJygFHJ5uhe8V51CrvRdKTfwRUfcuW1S1rzdc+g
1KP3KepaIBROCNzHw1NOehpvduI0gR5mflMAZg3uvXGIq1RouANvauus2+XK
6UZAKFsy72MAbPv4RRWRg4YgZVgYPaI32ZwSm5gc+deXH+549iKK14UVQRFz
/ou34dsQNJz9a7OXWZ45ySodB6VfdwthWZ+r9YMRgwZeGlo5hODMqhrdNYj6
4nOW8XUK9DDrR6Y5oix2sLU1qo5tC28LXyP8Z6SqWudpvzXPUIluQuFYnjoH
zWmduGAUV0UOVJUiBHtYV8++zmZy9p6DsZdUJALD7gdy4p1EeBVIBdojDG5y
2U0dFrh575gaqKjv8szTaVOET3/qq6c92AU2Ns3wGkivP1xgITiC4al6IBvz
YyvLTrlwBfBwEC4xqHrSnKyv1F/TdGaMnxnrpzdNhQqJ3LUADsoMSOlaKqow
uszHNZesMvvxx3zyN2WT3nEEWntWSItJsynFB3j6kUXjQRhFTyCceOUvUCkv
dLiXiCHYGaddk6L84VwTIxvpl8saLordeZIenVQi/VqWq5WKhNn2ghcf1AYL
MM4l1ndWOZ9vWXVLpwZaIw5AYw+UIAQTfdAVftAwBSyuMqetJIkjMRRpnlq3
NcfkfS+DhNGgJxkMa884UEK9SnQO1mRHRi3SAxIX57x1UBmKnEEcIIvsx9xl
a7Q1FY4lrniVOwFTbCTk7hGagOkpwQ/j8piv1wVVTqt1xPiy7+v/j/Zh8CNl
wYXu2N5bIeU467hbaECEXgD5zRO1zznMGGp78ibh6+GS3A5E5wj5IL7qCAOj
k3LjjNcwp8vpEK53M58TKvGV2M1QIBB2XcaNbS/jOOZlUwbaz6tjFuYfsGtM
onIR4Deuju0pZXtmaETSh7xlDBoAfPjdaHNCUj1Zwd/xwvLdibUw0D1nKqDA
ykpYdHucsGoC8EdHj5ly2lFs34+wrRAYGMbVUaJbdD+m/QjPK0bkgt7ULXDv
5lJkEmjodQC6zRGRASG5NFL3jISgbnMsM4HjECTuMXq308CKHPsZtsW5iOZB
Dkjs/TmOZnONqD+ROmUOpo65bruYXc4XmEtHXOpTrzDKIFwQmvhHXwAN+P7U
t6F5L9QN3ZCTEJfSjbgWjUsF+h7nWJMLpZeoIKPDbFhS8rWvJIR+8VicFwJv
+xNMG1H5V09wGFKRMVVi/NMXUWuXTxAg41zcx3JO4bF6FADTZWZ0m2IKqpX4
Rwvqz3oxusM//72H/mVwE2IZlxto9XMzwhiPXwtnUIJF1rL7m/9aNopV2WRx
6UK9Gmn8mdxQdo7E/FKhQPVviA6MNOXa1ThprglISbXEduStBpWIVmi6tCbE
kdbpdDUt8Q+lZ122YVhzJ7G5fNzFE69LaqpgtHZHeUf1Q29ZSZb/ZLG6zR48
MbxG3HsICqD01s3BJxQ26lBGYJJM/DNmsiWIfx+WBtbqahRSOsTIt76/S6qJ
cmL4+Dn+HMDvMVsFg0ZEx15AfRWLJ+0hA6W6M7gU4Tokh7I/umLXQ7/EYNYJ
nXTzTsg6un3AztKPkOk0FYs+DlnBIPAhcJewZs7sAtCB4jFkNPeGxWG1b4jg
Z6ogJ5ibrQ6kt7MR0q8RkSMN/Y7eBN5Gevn12UgnPbL2F1FPC0XuioEwBaLg
GXlkPvxCeoJvrTdAoTRBnaC40G84b1dYef9CZP8Z5ESgur4cDxpKVuUrRKNU
Dv2vDqMtEDXX9kKksi9rdEflu/S1XldlCq25Gx974+y7Al56EcT/jtP57jcK
hESB8juBYVEAnpTZFeF0sVhM3rogcMr3q91YoRhviazP8cj0MOtVQGYsvmP5
wt4ssTBU6D4/iD88vr9DAp7zD/1DdEUojnaUK1uUp/gOcR2poGnp//ldvAPW
P7r5ZOHgbOdbG8fuo1nthhymV1060ZrjusmpadwhW911Kptq6hP0kK5xSREW
AL5NyIEMcIjKZNXRTD+wlhJOzC21znIsOmYG9d1LlModSJVjMDIfa9b/WBWH
uCUsMesOv1/ZK6lBUeKX8oXzXyKqntC7zkxCliKJfauUPKC58fqsY6SYN+1K
SPhFu3HMrXjdZWCEGuEBZz8gP2N4DARC9AedYv1ErmPg2xMrl6H2QttNAnKN
kcPIelQEsuc/KprmC+RhfOzks+1QDLB2FMuz9JDi6Nb2Ah5h7jFOi2tMJ54W
T0v7S8ApzZDaDhzzUdz/voHKtI3R+cWd2WzPXf3crnOnqql2D8aLuMknDsyT
MWpiBoybPQQv/oeLiht80hvC1wDsY/IixDUohNTQMv/KyR/I41DrgxTAdG1Z
+lP8invHEwoc0VWCLtF6AN8HyzqmR3EQ5663lBmPCbtr9qCjS6VvsGUxEi1i
7xbNyhN+EG71JXeaxX4jTOS5Sdr6ITyDtL8bT4WMi3UhI2oRbxFF3n5RrF+O
NmIJK2wQAngScszYmQfTYxHsCpJp/jzcZmtPX9rEqbjjGIzO0oGXTtuzEVbT
UpWjF0F9qTVAy/tcG65/HIJmOI6T6tqM3X8lDJHNxJ8ktCljG8wGFIgURfCP
PggiL8zUxa2ToS9U9bA5VpNr7SefjK6JZI4HELjlYFP2ytzlftN1Y6tfGIJZ
8B3xuriamViUrarfQ7UbD/VvBMFHOnOaYFZ2uQ4TWFSoJVFz0bIFrq87c2ky
hj8m5ofKBzus2lRtMC2G/G6wr0b82fFE2rUD9Lia/vj3WKavJ3XoHrPOBjiw
O1+8dIgiu5jVSVIv2RuDyGQEDIB/WKIY+R1SGQGmJjnMT+yG0ALFPb54J9Lz
0GHptQEm3eOdYRfn3PQK9c0Yfz6+6YB4OkxuktCi1KjTLR/w/UvpOHPrP0Iw
GD6Ok9XQZsI7JuAU30fvtyQRa8IFKlX2A8SeR8193cAH/IOIT+CoBvKClo4i
mZ54oewpgnI4gplqEFvhBTbTnPVhW+z35wig3FsjCHKHxsp5VjkvBDRJUh/h
+1Nc5Vm+cTPJIawCtdWK4W5JOBBqGOJDheCTyGLqXPumf3T9zrOyPtrc137H
zAXt3gpdM6JRd6RXw4dXzXBeDZZ5GkorxZRBwWERvi8EYnAqD32MdQXfQooU
rHeXWRAUbuzHwoBhvIZPspYaUGJ02LZX6BwD47CDvmW/w9c2+hICLiUEch24
H6jPS0qQ8GGRal24Gl0AEMys6PerNK9pmCBCKB4aPBU1fkvv41tVHF9xsKOL
gCMplna+C+3UeulK+RDPpTiTZZvpMUPqaJAeUVhmaO+2CCJHxSSShy1MuHoP
/E9IqWJcnOn3lyfn8PTr/dTzKxj7wiT96fNxu2oUKRXw8cMBx3tynC35yqje
8aqg0I8CJ/dKg3NQbXZBVe+pEGxncikNpO1qymbvdRcDNEgg1lK8vmY3gAjU
ntiZvXOvuBmo3zsiKrDoSm65naC2wBCUtVs/79iEeBfeaFdfdGNFI+M1K/na
Sb8kIOEP7zfmCwwi2Uwzbyt7VLH65ztdZfAr+2CR/n8+D32xJrK3wGlqaQeJ
wQQhUVThGaGg88fAcwQdheiB1U0NKEm1mDs4WBe6suKeEE+lgE5nRp6cD6bj
WDp2uChFHLbcSn94LqfBmS4KHKrDJETKZGzPeDXC8p9bL6FntV9DDPxmSvm/
ZWpvovlF4qP8dqLj1cUE2UCs84sRdT5r8Dv4nKMIU3kiXfuSsa/24imFu3QK
zRsv9U2VTayZK8iqnJOVpAIDxgoCoMn+Qi5YW9NQAVJ+b/dqKGlvfhcd5bwb
AvBoeze98PLoKHxM6rQlV1lvdLzGmTkNpzraY3FDakoW2yk1nT3EsKL1CW1T
cY0JjuhrbJ2vFzhdkUzPRnr9XvGMwpDHlTNW0aj1syRPJzYgiRknHVEYLiKa
XJLRLlFEIM78MJehsiF5FGx3/iK22DxmsNf/kyEbPutftH2rkVvJBcIBSty4
EQoWq2C2coIgxe5aMfNmK/p2DeFQEam0uXEOqFTAzsOxLgvqxyZQW/HGXqgS
/ga6nCcvQywQYIFn4zk9g24sR2JTIQRMERZmfsOQbZ/9y6nEzzA7RuzSDJpu
Jve7K/QEUh5NVx0lDj8ZQ1Q96aM08INk+zfG5MzZ52M8HnBkocawAet4Yjvt
IbsNNtw2HUEtZruhsJGnzcAo3DkHZnQo220jkqu8O219wfzQh3Vss1gbQL/B
wFXVCnV+EoRFO5kruCOG9aDcVWjiCYD3vxuj9U0TGyK804hGJBUinSsA3mFD
IMSL5QgR2eklEPYm6ua61fKBWccnovcpvOh7PWsp9cZkTHePZOs6MJaRBlRs
tKApB14OHwIKM8C4u30Mluv6e7AhZ0RDGMMDferFIfIqCDqfa/sRkm6kMvhX
bvF2zH5HTTBEarLxa8A/RrXa+5CqWFIrcm0BrWJovDBTcY2ThQ8D8kmFKsl3
wX5y0IqoIPwFQLW9QuhpczUAU0ezpX7/vf9Ufsw7v/Vooq7ICLW+Lbmd25GU
PCLYoSR/s4WPNpo2PWXbChoxQz66nqdmy1L34wNjKxG02sLu3QE7k3bK4B7x
+gzPIwcze5whpyFM5HD0CWvtgz0uG829d7XGozP85SF1tHbo+ZaPEAj0CyH+
et2USQB9wKGtRvaP8UB5e/hys3pEuuuRqql1fpPIQDyVZ7tZikNm5PC5JWdd
rgNdRR/QYtGVQLFms1GI30iNTAFdz3ecfR9ansRh7szqQULR38gs1lSbMgYw
tku8LbR2+D4dGvSNYx95PgPgIDJpRa4OQyP+4m666YMDtOMuNH84rPCFxRLs
3PCL8I9+5AvRqkV5geQFPi5tM/DiPFuBoTXzXeNmoZYCLUJWY7acpNavwgto
D9ulq49832DIYpiP5Y+uCIVmvwJgWpamNGhr9Ed/Gi9i5iij/vWE8XK5C2Vz
ugQdGOMqnEWWjWwJ/k/4j8mhoGjxKU5jx9yKcOkSCaDG43nYwg4lmI9yia+H
Y6dlUci/quLEQdXEE3VFdqKBnELqdy8dktJdRDGJ/f+Si76v6jpTCbZBkQdu
pXOwFfQ/Z9a6coB7crWCX2YhAEL3kf4UTDgakrCCrJREUkEsWr9LdVwuUIj6
2HhbhRdFaV2lV8LJ+DKkgiNYA1JOdgtfjtlPVwKehhWjoHJ3l9xvIshP2iaT
W/lKNMaocV2b2hYQFYccyQNL0LEZmmjtHIjMou32TyRhyZzcsXgi9fdJhaV6
mcuRTdyO32ccOknwSSd8YMxVsf4EtsKaGtaBzgXv0OwSrnX3CLm92RatbUXE
CrFlXyvKRpFey6+palIQhBSWEd4qSpSGbGkcxJhexAYaA7MhlRH9MxIoDqX6
7ZOG5lPXTpyE2B77raPyPm3bk98NAEVyMMWKUpzrm46cFZZuQyM0fUaqTTiJ
BdzArEly2xLYfEzXqyQoZBviugD+O6KenYdEFLP3iTzBTz311JgzOne9JZXB
Iv48CRZau/H6MomkDxIYyx0IxubCnG3GY1jJCChmsdTBndYpcaMN3b0y2N8v
MDhA5DOjU8WXzajb5bPT943ISv3T/upkixMp9CJdC9ENxZh2sYc7KSNILJ0Z
ETDUeGc/UrhpjWWNZugwfAq1PV0VPNOmGnHwhkrPq2kxW7QAR/vnMdOuBJs6
YW4e8bGWDBFayeAmNGgUwEDPSPjOj/M+b5XVuN+c1qtMfl4KbeeMyadEhlR7
tf+eWA6xRwTEufBoxLFL7hlWtBTGhgQJbj0qMS58e9OSFY5KAf4l/Jbwwnii
fk7ke0212MzokshNDmEF3C50nvXpRMnHlz/7uyPDeJQfgohSqubGUrvymdk9
Z7EnmQKtGssA3rtzfUv/rFa7gW/43GuTy5nQ5Zn5DYhepH4Q5B6Py+qEPrM4
WczJpA33x87QHDdC+ADp/L/6Yp+PIKBtF5CWFnTRdbnfkUlHtpSrEFL4MN7+
3wzNMq1MN1nzyEavcswD1CkDS+ZLYlHevKViZp8rWc8ogjYyKF9xu5p76m7m
P87S/rg4hjgQAETSK8LIF3n8C9xpKcrgUyVH31ysZ8us4hSTHA+CWDoaerRa
ad6qbWfIY51HB7m5j5jiYKCucTdZF6Xu0sua0L34ypL9owz76HZ3At//6ASD
DUVS3VqE1x+RIrWHBd7d6d/q5TquXkrN2jNxcw4C5b1NHfy1RIDmVnHxCuXR
4RkCbF64k041ZXG/OxxhI2tJYrFjJooEHU0Z014Rf6wYBhJIAZEw6Fs+secA
xfCdG40qt3hjBFI7SFVgauvl9Yir0iFBZPFeMoPf9SmiZQMUbfxVS6njQU72
/eI3WosWaOTQQIc1SUFUhx9T7kBfzej+sClhr8aOHWzcBHAEO8ooL9FURlI+
kRT7Vj+lbyFZApwyyaRCk+mEhLk7rsvZAjSn21FFHqZSAAa5N718332GLy09
QhZPDzcH9egZ1YkilHrLP4gGysWxrdL6vUCM0Tsl+8o00nNiHV8FJCDkpgPm
guuemRGVH7DqIgB+jcMROWlVdBbr8RN3ssveblnUT+UP3DK9a+DaSj2qIihl
kz45Bt3e8/qkAMo7GLi4S6EweZufZNXDMI94gHXXc+0dTJtbMgJSsO0Tlgtm
4cdHD0HqO7bPSj8eOVaxLOc4LzKJzfxtAbKU+HtpszpX5JHka+NLEgGMWBYi
uWC6Ll59GwyeSRr+fehayLBC4axAGZS5SdJKrIrc98BE5P9v5Hi/7Mwvktly
wy/0hB04rOMnJDTi7BnvP3GWUqsXTBMEcPJyyhR3zTMldzVOYE4IfZPZvx+c
KhIJi9Y4+JQetyPkj+Rdu8s0xgh3EH+JHrlpSOfrES33NoUDYVl2GpEk1Ew4
jV9meY3GlnLxAM3GtMfIqT8t2Ra4iQowCY6fFHViogkqIzzQgVOd9m5xV4/p
vXLJC7iYJ1nFRQKoc8lKccBQAI51b5i9vD7Z2uMmAjHRY54xAbGewslQdY2P
l0Jzu/jJ+Sc2gGTpJX+BREfg0AvdZu7PFgx+HDI114PZ3U0078EHqwS6OpRK
ZezmWz6yxCxgZ2zCMOJFCJvzoPLLEPFgiWJpRoHecytkNLdYqx200I0JpBXe
Xz7KJaeth3OU8qg+U++9EumNBAEazhWYoEvK9nDNcBKTuGDL7A9T+xrbon0z
sO8bIOGYwL/d1cB57k71+QrY0Y5iCfCMt25hocwiNc2lhJ2M+W0evtc69Uau
GH9gSIjRcfl70sekItL9TYwAfZUaKmxEc213AxlieEntQXCnKMuRiQAlaYYS
NSxHfCPv9Zp1rGr3u4kKsbu9Kn+wLZPbewW+ZfhDjXGB4QiLWiRv4O1dzrG8
UYOwQ6HfiwxdBKAfPPVAKNAu2jJtM8xm74rCDycge360Y6NLiyqzLExu0HuU
zGq07MQNsoL8bX4u9eFLJXNX39RkKDNhoo7VBTDgESs5gELv2/jEe44WuMDs
2tFQwzGE0rHX3y9S22ZDVJFJ7pxRU6peuKhhN3fA8cyExkCOUVNC9Z1LCxel
UsHUMlMlNyJpvdlNp+RJpwVRpneFDklUxu2lRHmEwhPnxKiz2Z3e2fjfjxhm
+GdSp0tTTBGz3k7eiyNASETQJjyYE4dgMO8cxXDrwt6qGVCNusL381ol4xxf
W73V1U5nqDH+dnzvNZbeCsa7ZSLuh1wU+S4H3cRyIPduTEQsfxcMpmTRpoG3
pR70zdZkSkz65AQgywWweVF+RAg2vRF3GUuwEnyMq/4Xn/aEFJcFyVLJWxVJ
4PZw+pKm4XF1wOtYQIFMDPBZqcaL6RXynvbt92y258AMGEBtFotpz5RTrHzG
cvyurpmF+uV0/mPG4t0Dq+q+wOq6l8gRVgRQO/NcbxXrjIe+10NSVtX/Fnr4
Y9MGlpbKbtww9vCy5IGAUhD8NJZhM8h3kzPsi9z1psg1EfzfHpvbaW2mDeOp
dMsHbuixTKhCssd1v6dfTrch+Ummv4FszvscCSPjqvEpcB1dNcAwqSp5etQe
rxXxcSvxWOobEq65Wmpvg3nJHmjHrEONdIDcRIQhRcSZ5Vi3J8lrjNGROMUr
spntyrc9XRz11c3aW3FYVyYuPuxJ7cAFnlEpN7fBF9/4EQ0YIBn8CpvVkZ8h
cBNhGF28Nx+ihd4gmAp3hrmFITLQruw0CFxaAgy/2/o9Daqvq249/8vuFGih
bJX2UA147igYVCZ9cx8obctCrr9mvQgVeniG36oET8W3DrgD1ih6ZG27TFMA
B3LKFPEgk395DvusITcveIjGAJxE3cfu2FM5AUttxeguwBrsHFsMr2fhZAPm
US/JLCh/pFy6oVyoF63UO3mC5dBe+kD8v81dAB/lghmwjnyonB/FHbYpvm8P
B+hXX0aZSmXjGNVQ1RVAAp8BTePDk5sbjSwFhkOJCNPnV1qqTIvgLgoIHzVJ
GvTbzznmAHAayIsNDHI+hjPJG+Z3IBs1JZRRt822zOuh5zNoSsf3QAuFDzi1
Va5e3N1DKEH5OuDwQAW8duQ5uVWbBU/JHOzyHSi6fWPNGmXGn23X1vvH+FGS
yBQZM1CEAZTtNlgJX4eeahyHdY8J1SSQaND9ANK50+HDDoldoAC3enJD87bC
S1PWUuviaqxeTJDKdXygF/2AscNe2pA8Q10EGI3J+vHZVQi537b4HyyZMcgH
ytFeH6tPWUtd04xyLUHn79CcnEqAEjAbhALONXw+ki1ZLm59dHx7NIEnZHCI
nozDq86Lj/wR++9q4B8cOlKdPxgU/EVPHgeYS5YtcbvRodz98tCADRd4V9Vq
snTItZKpbwNvCYwkhKBJpr34Tzsi/u/UW8ExDvncSZPs0dQxvBxqi0k3SvNr
hRVlyTCCJ1tuJpE5DU/RpSo8LN2ZqxFa8Fs5hR8LI+8J+ajYf6xf3sr5lkgA
MvzWkok4vjuwSQesPsYXBDwczFdAAIp2wMry1ZmN3lTMOeBh6ks7lO4lWJKp
WL+1XybbwQegvUARAiU3WA/RMYKfSlDx+GxBbbs8CQNn5jCyVkyTa37y+Ycz
/Akxhh3x1PaRMbIjCvUfppcre3H3r86SZnf2ByOWUxsUbgoJargnuz+sJ+py
LSSyrV2v84PWFLa1Ft1yyZtGw5eZlwf13UyoOCJt0yHxLVTZXeVY5vsEm7BD
ipLFxgTmYqgp4MBzOTMP1ImyQwuv7JSV7FyJYp4L/Tbh+fIbZy8gz5ROHVOu
gJzcHwG8FJzXPybd/iU2vVFzNpWjPdZU0mL6DNZRfb8RlB1s6ORdweqIrj95
HVXdsCwHiVggkhqyVmirTgshdaVLsleNrsM6B8YPa/sslbT0Q24oqDAZl5Mp
qsXQ4YuOW605ASCDoFMwuQNthkGtXOt27Bml8gzvekZ+iytvzWxSuCn9V5WH
5+ceRcp5Auk2BGpUx/AvwLNlmuLjkl3A/jYlhQ/KZUkH+KrhqRNri6Ri8oQL
tCgUswRiexHBmA/85crBSmsqLIyQEFJyxll04bOSfb16F372E6ZzePdmQ5MD
hQ2HcDGslEfaxWr6JiRtV3W2sDYtZx+YwyDSWTrKVBfuuotgJX6RnxbIwOil
AM0B76Wk1p3FPAJWAYZIObJv/JhFEjMRskvQgJdrzHkQSH2BX0mOPvym2gBZ
xLwOgQKavmjQgkNzXCjD8Zw9DVgwucexZWqZtVi2+ImQ+giBbX01tVTsu8yT
+Fd6Ra2ppDRNliLUhgEA/stp18drBHyf/e4wGcw+fo8XyVxLc5ACql2EH41h
jivoEppBzTvQbSH0g6Eqos9iz/IHIbcFrKbZDT6CaqyxiVdBJV2XL/7irsiA
JfJgqmqDHhISTtS9Fyfm4wK6xB40MwCmpKZfBUkCumdfKQ7LgGOtA6MfLIzc
sxvSxHxWz5NZWsOFBO5EOKn8bZsU1brXVHsPaDZwRZkXOfNkILh9J1dNAk0p
xD0+132PLlDbErGhtJmU2fGhBhheq15jl8Ekzz6ATqWaWs9WeTSN1Vl2lFVV
R9HjksG4GGrRnYK4SU7p1OTYxuWXqZTBdcYTJlU4cBw/Vk8YhoTCUt1nQBo4
7/L5N7y52rreiDrx1QaKQWoZQ/99ZTIFWKGTi2jdnEl+pnYukXySEBZA4K9o
tOgsbdfRofVirm4R8rOrJWWoFzH9ebVlqnuAC6nUVpHVTVks11ScfWmu2h3I
+i34p9TZiFiBwnEhK0/CpKZmDrwEwOv1uh22zg2iI3kyTbTDrlnhGpHYIPwY
GQYT6nP/iDLxfOiGjdcG9SkLeH1BtTv5LHiEXfhXUFgsrtnr0yrP+4sMVS4F
CfEaXtlOYOMl2v7x6u8fp8qcRDpGTGe8nkkE5euh49Ym9QISJm4Mn2DLHsi7
NlQX0Pt5NsLvQoG/b9sIasKlmhWZXYp5x5rIjEfhNkIfrXq8HhqM5jSzNHD+
NRwzl3XCRZ5QWjfFEMP1n5VWJ5/075rSRz0OsDdrbYoiDxvyAs7+WkZ6wCE+
PlJ9dO1Od1W0dUSkXbUaS7FlOv4YCq9VGr2zos9EtFGhUA62onvgQw1emTAT
lW6dGmPn81br3lSzJpI1QV81AuF0/EKFZbWhehTEMelZAHJmWDOg91pCDKd3
s/BZk1Xsb0ZUJMA9YftdKzABX7VF/8DHADvQngnv6IyzgKbEEUNIZRhwtjTA
lWzrdpY7/xZOikpw+M3tgZVF0WMjzgAjKf/9QG2MzYeaEDWmEd1nuE9FFHQf
OIqrgsj0tymsWyC6UMXhmDGMaQePTHgPJBA6cXx4D2XESLIYRDqjzCLztIA9
pzozvuKVMN0qp0U/KZUJUfv46vUqSg/hgfaVNdpp30eWujZGo0x4jJ0X8Xq+
ToV8d+gYEKY1OEzgvyAKBx7K567PbWpJ5yXalGgVN4+0lCAFp/bSjBzRCtRb
tqJLNzSNuOZLsNTkSE8rEPCNH6GEV412zYAe+luN48jdb8KfW3LPJr2k/8t7
TB6TwtyDJvdddLyeBFSwccOVZZQZH1E/h+QCf9tUIZm4fLnIyzMchp6gYSi3
484eRktoUKlNf2FILjWJLf5ostkhoNN7yZQzjNLIorAaJ+vpyeT6qKAb5Wya
v67PqXYDrOgHkjL+02djrMMz+31nLAjdjM60cy2CR4vwhtnxu3N5MYakCmYS
jWi9B4kQm1zRdr6owf6KzLc120v5Uuinrmw0rKTW7ncvoJD8WcHQC1IaAxoU
1ekZOf53wzF5XcH93vYKdjxegumvYy83uEfCO5hdwmtxVRJo8F/2JT4usOSd
csppsXughg4usLL5TXJdY6Wd8RqTl68fTX2lf3XGcBr3aBdL6vkL0iGMG5ix
mDaa5EbsDbsRTpoZvrPWo3UMa+8diuS0tDcVltYK+c7TPm1qg/CXt4qRYI1a
nIgxuSxm/4LLDVr0/ZxOyAJLnJvzPJ2HkvmnmFm5MqQ0rtqGDxcyNKLPj9My
7KmFA7qxspVDZIxnhGV4huuJXcCsK2dpbFN3/llKb/WOA1vSUQGpGyLG1eXM
kdEuGBUxe5psnGBdE0TUB9dWngnDEulC1Fk9kedlyrgeiLz5xjvoQSIVVjh4
Inm+4tM8IWLuGGzStyuGREv1k/dAN8L58JKUiPXjBWiiUxV6o4Shsu07atiI
ywTIzfni5byvOJDa4ylZASTo9xrhfFewWSdbMdGM6OUy2ZGmqfiosCt9N+k1
o2sC5Z/PlKBwQQMj55UYRdltOEDpbtqUZTUopxTFa+QGiak/UkjsxbdHmIPN
9o4lhqTB1eLwdyvS2QOWIvbrQonb1k5BtZsT+S6A63W/afiAXTt/77dNY+Hj
hTTBTFDb+kG1QUGHjtJkt/1hmEa2DY8rwifYFaCJBq0hshhtnQ0JVaKx3fkD
IzslvdghufzhENzWy2WB0bQvGfRnJ4BFCrek4IvgsAJe35q1B2L7BjxdJBWc
IzWuv05KTE8L8Bmxo/R48TZqy0b6+MDOpSO/bvg/Hy4Qm4nIa4WGE0kn/p8o
lhujjj0W8jIJPtMjVzonJ1jU3nJBC5Etuio67yMc5w0ATbS86QAXGa+qPxHc
ybI6C5eg+aY4RmgppCn8qYHaZu5xjrt385JVmHdBPUOHqB4eCEICHyk7BuVy
Ys9BmsfZsODjZf7KF0sTsuqf274npBoC/PrLpbdXvj4X808FyfsTpefxlJhB
gwBjmNK/xSKl70gBtf4/hiXYZ8NNs98CKWhB10NNs3+W+fRP0JMiNbd9IkdY
cLY66/FUnt6PizeH/gz6C3+/xgjwIPgxd/cMhhyEgws5EwHR+EKkmbTo3Ief
JVgDKmJAjDXOn59h1pRiAqEiGaECfcfOiTA8laS3ZDVcomPWZdJuhuaTH5HE
+EwoCJxIQAHBBOdgAYTUsdyI1Sj58GnbZakyFGTAxdTn7t9yZi5UmwfkrPVU
yZlv4rAFatrC2XurVT0ihCTt5BcA2drlP1i16lSaIdya3vWAl/YsaxxGE6Nz
Vvs/FbhTX7agELaeFjm6tpSsm96gxQ+W6yJeC5ytGDQAIOZMeugNFCU81CFv
tRz3Hx787CBPxsVTLON+HHIelPZxB2MbVebY5gxYON+nVp9AqRgQGF8e1sYv
kD+IxgkF5kMhrdhmTzvr69e87fMsQZlmrhLZLxdaWW5H97HWYLAjMvg4TVow
bwkpfOkxjAKb3ezSYwehfxYNVy5By3lOS1AGsmKnh4n/xgODkHvnfj8cV6qC
MIhSdX30ZgzVTJnMp2x2KPb92+J6DEmxs4A1LSYqxFmUTJRVUUsZmdXZYEzU
fKpJ39z9b5R9bfaKfthclSc72UK/iuhpZRQzoUGNY7g8o6ly9Rkl5kMWZMdF
J5FUlbZKsmwAgGhoGzbdEl/eutMg4Vy3N6gJE8j9Vzc1cBqFJkinj07zCjMv
IqtoLKTdrczDm58gKTOTS8Nqoa8Oeeg5d32TOokEMvIV9b5nsyiK9d9+VzYY
5NUNWu2ROI5PHoo6L5e/zsBnnJBGF10AGTNUohMNadYYu55DH4d0FxoIrKbm
/Qtj6Y/7CV6NtE312YmLj7Jze1kIdfdhqQp7oOCEpMbRcytpwyMUYoy5nzH1
pckwnEehJr/PeX42L0kmjOFaSynC/as6G7qoenZhM2rbqPNH+2VzExFjOs+p
vk8HBHGU7FJZWplUeqk1FIF4oTn3CuBt8oxcC+vBKmrNlZOXH6Rc8A21v1cB
q4lCsjO0g+ofQcj2jZO7wiuSELsLs4a2YpbZtt33z3hacIm/HMSp7nYdtdT6
XHG9ZvMJR099Ks2D2tocjTaWCptgCFSqw6xNl9ihZpIWE0QGE8mcUVi3kp/G
DqpGE+rx8LYAzWCEAqC//W4A8L8QFo5xS0/oeDV1Y3KBMIeRTOODPVBYDIqq
RDduUbNPOxQZqQe2mV3L6vHL1Wj0kr4KYRq7ZC/A65D5vK0YizkaWwy9c2O7
ORj6lg5lqQ5xXGe/Ja/v+24TQkcli03ucziqde1PDzbmC7AUEga7XvyM9XcY
P2GbJM7GIpQjV+K9X2mQgGeAkOETuxVrqxifqV/JxrD5qsIihkZ0fLzX4ssJ
bA1Iw/4eEmVrvJv7CX2uhflLnqFlih5w+rDCkzhs3wK141O8DvnToVoxinWv
qcA2FnVX+Go/LpSdHMqLG6TUk2aSrGFFs9j9GJflCOWgxo23XwNTTmJmnm+E
Qh3nqf73Ha851zBcf3PNYhdoAOPxYm38wbQm6gb38T6xITtxJW7pQQ9RYXKH
lmmfYByqJz/PF2holcToPUjjOHB+IsPNSnMJJpnbps7Y2jr1v2z0NyxxPRND
DDkikCBWF4UKPK+wWqSii7x+QYMTLfixbVtP5PhtjWeeh9e7yozCgNr4kL/A
o0R1hLqR5aBxv+YxzqXnGjs1fb5x1VvYG2gX4bvHnDCOAmcF1pRk5gmsM0ES
KR7DE54QoWxTr+Sl08XovT6mSvn+WQGxwLmjpIOUi9Vj1tpzZfaBwyC126ax
5CA+Djf58IePKXMsopb/6dra8/7T6Ef0l4Wx+qE9mlSYuwR3lQTfjvqlAuMq
17Q62Tqmw2G0g3KT4RHSH8jKllV7ZVoIU2RiimXiNBD7UM0SKiH1w9Wy62kD
39j1Hop4IPyyXPfs3rNQxj3+vhjvdUsE32jDWyU1VvbZIqOh+nyY85GOA39u
jutWIBOquvPg5/jGN578ygnz6Lcy0kLpcQ2KzM3uuSlf63kBZySxfCVxWdJh
LCNyA2D7N5e1+5kLajAbGhcxvkAf6YJ9NTrpRDC++mgGVbvbwhglNUuT2Fht
DNsYQxNwA/pgX5tdt4gI1aFH4FT8h6L42Luep1R+8dlOPuYhKXvWyb+fR1IY
VFMPwcSKYT+c8T1AYYZsSIQd8bNCjAAhAZwrOHgUQgNyihILNiKlkZbnC7ra
acsc4GnvhVTJkHp/k2XjhJUb8aN5XY6rgziRAWyY9uOf1qItrslegJrikeDR
vDvtcm7N7pzK8BvprGSC6YEmTnjcQCvlGjVHHxHm78oHnGXbQCXFs959FZt6
wfn6XmGGjhMftDGKL0XAaPWGietk5e7d7jZFmb+ePABYTlfaxfq8Ghsatpoq
bDNf9CDT+7Yig1rgH4kCHK5WN1gHDl7EDexV3JbQDCX5fW+kY7aqxpLQ1StM
A0r3BvSBtbNGQ0a3zp52uTlRkJQ1qsq6n+TMM1WgKa1f4aCZdRSGgabhS5QA
zQ5ioopuRVsBKhnH/xkjlDoa/lSlcYzq50U5sHQ1Hq1hI0HXDF4eD/Ps3sRR
jKUtcQr0fSaY85soeIXBsEnYMvm9M6t4NomXr4ZMm73VT9qi1hV/jkiT16Ov
GJ1t02FlJd9/Gblwf1BpVKYAvDCy50dpqCWpbF9ewHQA84OzMYwm+hg0lilu
M5YJyJ/b3zrwu7OLGmo9hqGdfiOGU5JTG9iAbOl8F20Tndetx0b89gORIdo1
Kclj8dz7Yya61sBpoGiKMfJvDXgASelIx2LCNvfFZb43Fhci2r0gQ2IBvjAG
0keUeTjGSNxY44KmRs4L3lr4kMf9cfbTOuERAuGCnKSq9HlPdEMaiA/hED9h
bL+Qbbl65DEmCxBqnbgaC3IBrmwkA7lqZNLeHcw2y+hC8T8DcYACZOdtrupI
NSu4vpk/odKh3Q6ZKSW1nEMMgXmt0Wq7gQayvJwg0o2TJEwiD9dXtPVNC2wj
EEi08R4bpHZUh6bsKCX9nz0w5Lxot5oy/0HK13RX5aaRJyeEjHGZq9U+J9Ia
r+eXTXexz8+Sr1fhGIeLniAkEZg2MSF5cxW436DClzjC/luisZs8EnRJljv4
uA4SOy0nInLGtgDQaCnSPgr6tEjXZuqRTdC9ccaWm/YNPXLMKY7MZE2+kHFe
4y7GHGdPTVpPL+8rwLpAZbUzh33chM5yzb/5CQSuMnJQkpXgTQfVf05SGi/r
TN7MrkJyw06dO6oScdin6LqzhU45GqYlN74KfxYbWX0z9MMKg/2ykUfeLmEK
DjW6pYV/KKI2sivn773FT4BFyFJHkLGDGpwpf8kt3XVo/h+9HJOfN1seZs8+
XUTT+OcJq5GBJMUXtlwYBrDbBYHUeBKeOzn8lUNdajI4bkKuG4Z04M45DebZ
xt+Bq8CU0ILytI81Ox76FhGaGQM39ratU8LNkY7FLEEPK9SFYXqTJYmjO7c+
9AFUVzmNWrGXjFTJ//90NrTz5p0JhTvLxr6PT3GQ2x8siFv2tlshhg6cHsUA
Ng7dHFystByejv02A7c1HTkUtoFWlE9VnzihA6C97I8kfrD7HfjdUoq7CYs9
T+jbQlXt8RDHJWwpJ7NU4kqi3w086Nq6JhsuTQvurN5esHcxSJQOhd0ZrzZu
N/yzjsAGvfQysv9rta40TO/VmzZy+M4LDzZ+/cSSkorGZPWOUY8mEgbw57G0
+T+3GjCwuOOOJfWaB4MNg3Lp8PKPTSJPpWH1qkLDp7I1zdIBXQ8sqwIuvSbY
AIuj1OsgvdHGSmUuuzIvdosP+7nzEghaaqk3nD+Wn+0l9cV5K7PnuA8S5dfK
tHfqqJd3/TAL/cTGlEeDiaYW9GkTiOuogLpC2cDISwhdd7PGz1+WjGr4Yy5X
KuGgjVoeK4TcEv7fgMTH8C5O0p9PEAE4h5H2y4OvKMRrZ6M6CxuN1IYDM63F
xw0rjul6deq3l4UbLqFr4yS3FdGqHGmf8EiN4TxbRNAXi72VffijXODzjvcM
9d1Xn1NFAUSLQlXpeE76xUq+flcwbBZn1G21/pqvQk37IMhwQ3ohYyi8/6y5
kb4EsrhGB5vWkbq7Kejy3PJZQO2erDokGSKnN5eh8fwY1DDZzp0FD5D3nR3Z
OtZpiN8GyvLS0F99fUOJWv3J6+ZfHl1+/TdDvSVKe5ue9NacykpwRqFtvZTg
zwGDIFuKmVXjn8r/ecSpK6FZ9XsjxUh43h4tMNrHwyTyBxK2Jv4XhbykmeEU
n/s9YLWWFwTuQfyq1hbsMbMY2NLOluwbP+Xrhcl3x3BHaGfGiECyNWHaloLW
HiY1FcUYsh48lgEXpHfpvgL/zoOcEIxxccSaNHhxj5xGP2MS64ceJtC6Qjb7
kLPx3oSXKOxpTfCHMTfC0mW6QrCMM9iGqhVROFMcZ6CdIg2grghGm2I6qvZJ
TWz9nvM3IVWECNg5wNTJOfV9DViAlPGc3mjYfxokfsbmax/jVZ8SML0rN0D6
dL0mPb+utL1ztYeh3nvdKyn4kFsZqt17XfXga/24HsauO3+qnNBZjx7+aMG3
gmB/Vxgy5ENVkO8PAXES4Kp5JLKxvjGBs7gY/K5h9faLHDG2oT9vFhItaOGK
wuorjKOtah/UdxNB5TIHzey+OeDFBph7rN41OnhfiAtu2xRZZ2wmYCKjGWJS
S03HwoPH9JYu+3zHXlq3a1u3WQ70MZOyAvWQpqYz8xhY4rQLyuLgeMqgp/38
zWvzgiiW9EpEG9nmoNSsHqjagPwLKMfuwSuJvRPU86J4OYKwOC2+hIcKGcBm
qrRl0SzfAqR95qnAr3Qmm1ukZorIu+Dl6ke0xCMlN9Tmaf0KHgX0WYVrj5Zt
5WBYm6xT9lPcqRZVwUh37GdiN14gg6dyWqca5rAaYfvLVZIIv6Zi4QLq1ybl
WLfQbZ0OepOe4bWNIbw9+CItDiJFmJkkii9+kxjmf/OdmAJWOKvTAGIQrMun
5GF5qCDycCqGI1Lq7WDcVRCLVCPinz+TFmRxZ3+VEQG35gbHGYlSO6xZAp8V
bFXKrYLwKyJqNtmePkCRElowQkGi/z83Uroys+UsY/C0DzzH0CeCbgNjYbBj
s0Kvc7GVFVLS2+v9mgxRbkh7yGz1FSx7xSn4TqRA0rq7IJGTxT2rL6yJScDi
dMCMH7biVohXigIcmSZThapOYvTOxEs3+jIUOdHZsIfniMV74AKEqNqk4swz
dssMYG9fpmT0SKraTny7xkAAuraPSTUB1AcqvIOKy1c9eaYFeZPtyf/ZiqeR
2tiR9RzUlISzH4dSselYq1nwERDWMG/DPRGh749efbf38W/KBFkRcW5S9/IM
oV3qidKjoSCeXgWTT0gdul9P7S3dyduMJhTEmVG65zb52pfXGgmXX/FNF/w9
17zkdY5L7sdtCQNZ1LOXuvH4FnkFHZ1auqrjepLjQ5ilUeXcCX3pVRdx8wwN
e2imlhX23RaR23AMMBWSDYurUKIOY6Sjajg9aRKtqJ61O4+KzaaBW00psee2
9xkRGdEn/3iTyr7D/itRigbddm4vziUNmjPHy5D8uXeu8U20l/xElOQrIeWv
lHMrTJ0YqL0xCiGgd+Q0xx6s1iQUTa/wm69I9euoxe2gT2iq1lO0nw7YFPYm
4EcZWzW9Di6JnE4K0zHpXuxeRZjab0DsYfAS+O5zc8MYv/hnT4w8OTLtqDUH
1EysK/T7tE0FCtDQIxzo0zKeuTz1yWIQlraX2XUVO/fmDvJTQ2mG0xrtMsWG
WRn1kDfxO4/R+WUGuqOMNErvIa4P70PAriN8v6Z+0B5+eaBlwmmbi89/+mW/
yA01BC1s61tFzt0joCa1OsTxZvXuAqekGoTD4fI1koiOBF5E/aDXp8k7z3BN
dMWHQJbYS8D2XVVhJW2sRwK4sWp74R9zUbZZr/pgq1meL3rarMufM+S7wIM0
K8yZmm+YyTm2Jnv/UlvjPVzZqTk2V/PahD2zmeuj5rGxwAhWjIOy612fRn81
FBWmTQy9sO2/SQ+yZz+hz529fqe77dd2OT/BA9Ps6R2l19QoKJcvHGPTshXi
v54yw7yA7TTC2RuZyAGNblNyYizRIX+FDb9uaTe86micpVn8x+T+M1tYg6E/
Londrp89cMRvocNeYz7TSr317RzeDh4JHd1QcluHfMdYbfutdMvTNPkjWNoL
9ik0RvCL1zL2mq/mP9iomjpwgmMXt1+bjePxoHIoO6sa+2mTv4LsgRW7/Vpw
kwtISkTWluvfCU70Cea9X6GE5co6YkpN58zyt9cXaBeK2qjKDn7bPch7Txa4
jhZb+QlXO0p+5iz6MRfIW9fy4D6DTPhsLms0cpndTP8BgErsRgVFDEqkVo/9
p5V9AQ/1E1g5U42IBYY3fmkJU89tfzV93t0NLk1mO86wtLswp+RTr8fr+P8A
OSL/Sq5nW9M1LJonX6CF0wIcvbTDcuM/DTgyNYj8KiqX9Qo0tPy9VBcV20Bq
fSqaBA0PH2/htvaKHfdHA99gkOVrFvdh8vbp3kyCWx81Fkhpnu0svhuB1bdL
8Yimse+tzZQ2UUR/NzmGlIk+YaFLRYgLaPu6GmPdvilYDG+6GrvrTkAItHXb
N9JpRy/YtZDuyJxv/caTamlP80laBZey8s/YLJ+Si5ye/nPrWxpFJgIDDdfE
02a2BV+ONRqnQ7CgWvF/SgCMFCw3H/p3QfSJ7MxJyK6JYkI29Hq09145s700
IeWoFURUAVCehlYPBlny8hYdFTJoyQ/w00jhh0J6A39UI9dpIHCccGhyYLvA
NjgWmqFbcV4/WuVWmY7/+v2TCQGFiVBLCHrdgzDq9xKDpQjkT2xyOfvC5JIG
G4ZozUj8suvf8v4hpHvY3Mfg06kOtj/uG8Pe1cTE93tBNdEjDT0UldrPTEZc
rA3QDM3OutEhWhvyKGO2oDS7JTRQJYNcthlPIEgJTDTrMOhdh3nHxvjvb1Jb
oeRhJbkFhMOK3snuwTo6VC8GsRYhJPT/uxWe2amPlvrKkoXtz33A52cHGJ5X
P4+dNC+83U5Z5AdPrM+eUCGd5Pv6EZqAlGx3TTcBD0OsQVU44OSbHD1ivxcR
/07xBJtn5tFnBvp8STamkQyxoSuKocVPodhIfKW8S2X+nikma+YEq2Z1DhGm
gFwIT3IIyEqol6WBcu5yKuYa1wqj1yRJcWsxIKbjfPgtpTp1zLyv08f84xqu
ZE8jEBT3yUSc7foYMykqWCsahNeaa884ITuvFo+NbPDZGJTlMP3rlJYcA27N
1lFc10N6xEETotWrOf2g44Q5YPz4nXmZIR4no0bl4u4K918wifds+bLvmK8D
qpX16CVFdidVttKqks22um/H0hJb7ybZggRi+wycCwC2rA5+/hpO6VkJviE0
5JnHrjP1mueexW/yBJf68CB5GtQNV3rI6dpdW+EFkfnBchrMrEhXoDBGfOXx
5Wd1VXaOSbYXRV7/A+RrXn+8kPOmuu/3CaovCSLV8DBY/49mnlbMMjMm8wop
pBs8hzhe9GbtwF2VGeNnCUAvQZW/6vg4GKQNxXKuE7eNjYV1HSMR1cpzRN3i
h1vYzYqsGGnbXzbWC1K7xbjndS5ajFbHE9IP7IwDQgtOhGsMFrQx9TYfh4h7
1V7+I3tBHReMTVxyCt+tz+y1RcZKlYa2h6EkgWonCA2LB9f5h0TjfrLF8Sk5
n5VXWEKGzDmT0NJkRaDdSwIw4D2lUlWQYiJ/N6EIIW+nm4jFXfivE6p8x4mo
mRDfB6uTuXDi88GpT6+LHRKYLb04WBx814n8wxwK3cLh52PwwxH0jjKSYqp1
LmWrUP8MFTGWzFXHmMTUfT/mBpjYVHEGD8dqbHG8H8uGZEKJVDGSqKk3qdtq
zxECm+T0wHLiQvBNGFNKDp4dUuT+Utut4Q3AfvuVuY0XAO7tpRYb0D9kaLBi
HSl2b7UJwr+tLNQodvyYvKP+t1as3Cos9cPvGqmLhdXyK+whHvWVDE3VRyEN
x1XBW5UVzqBF+0f/sOt0fSQ5uHRbAx876S6j3utvB6njPW2FScrjIKfsNOzY
DiQ3+Yfz36fvC/auNPBvA7fAJmiBfw0qA5ItxxPPM4uMD6LvCyaOGkC6vhVY
NGio/a+5Ui1m6v/AwG6S11geDu7TdY9GgG9SPIBZOR6+hSZpguPlz/vwoo6N
mPBppZ4D0Fl9fLJV/Ghw4YndvU0M8IZ6rTbXIp2CKbD/MPBAcxufC71i7Syr
sMqeA0PvuC/8A3a2Gzgv52jFeZYmrEj1XyQ4g6aS/O2FL+5TzELL8auj/8T4
kyjISYfd9huif9Ht96Sm/RVIeMeYRPv4MyfUasQQ/t23ott16fwahBwpGSYc
SnZN+ivvKrSCE480yeZvnDpk1X4rrk/sMlMkKr2MeRkHyogRruPsmfG4/JJt
0zUS3f3hsvz0S0D26Dr+cTydQnjfAVr99whcm0t+e0+KmActV0B51kBoT0Pw
U0/C4OKtcYG841jiTjOX966AYZsGm4sZ1zDD3TJ3oLWv02abMkejSlmyMb9H
vYkB6prNchoYECn3NTWJYb0qUr9HRF4LVCXPNbpI5kerZyPCwY0PSqcvmBGM
1btZD+sVsVNDor4PZqYryTl/0XqKHfTDECigQaQ6EBwLGjKMYnowhb4exOrK
shqmNvpaWCKCJoM4rGqAaNbXhai7D+W/SAexqso2r6oadENnBSE6TG9PCyC0
GnhRLcJHSGS33vM60b01U409MTYDS3giDcruhw36D0Z+0wheuXcq2kTp4tBP
xJApTtUr/CaFNHTJ7W07rdTeS+W3Iya1tExKqromOUc2bOUwezZ6g2V2p5CS
qvPK39N0EakQPsKW1C8jYwPFJg0a8b07xn1kG/LBvYp4DY2wp/RVW1vfEXy/
0noDXdygAw1L947dcsbB6FHbKleuE57z4HvCIXcLzu38olHWBDvIP/f+oDPb
90TVVML+O88/CoOPokwQmtzDfDkdBDce0+AyQ6kHESeI4DvbF/GLgGX0z+Pe
ZADirYkFBAt8uXVQOOUHtnzJuZmlZ/7UffmeNgxOgiGZCFkIw2+fn4ugvnnI
KeT9xJkwZNyqBns6cdm2wIA9toogjl2j2ibY68ttwNz9knkMV5DKlz1hKrNl
HTrVtYseL3ISkKgYZual3h8pSzdDUmP1/zTeIZXFzpC9bvwqfsAyMlQnSPg1
YclIxKBgdcDQ19tgEMp0olDi+Q7cSswdIiWKuTOnE3arUbp8Wbr81qQDYrBz
FKhuOfsjJHxy/8xp3mUKLfmV3JWMc2Grih9VsBfjGlZH99n+AtStBnzbTg1p
ImA6d0M8piTJDYvlUvlKuB0nJePGaSN1jwW76YPEOURszMn3q7zpy7+VWGsm
Ab9WWYB4j/ceY+niFoC4PCoKVp5jIYz2Fu9UgP2HV6U5QDHaww5MCG1a8iKI
b48KM8qLGkm1WfSrPXKQD70fNCemAIkoDN0xge9Iq56cCweXS/UVFkygkzRZ
wGP4J4I1A+iSqR74sPHIfOvaJm3NQBuz5AmPB/gQCkzlYZUoOjkznpy1vN91
eg4iThgfsDj+xT0lwzm/1I70PqPqL0S0kwDALyVet0PJqY3nLB1Hk/1muYA3
+T+r8TJUarPkehlK5szDtxlZlo/MDiYkqKV47kBKvnwXBANFZHHA+ybTwuIS
nR9l9CDFcl3CWajPtvLkhFLzF3zC2cPp+yCP+zlO6lOZVxbIym7TZOGtp2iY
ZO1UqqI4Q/chCvwRDKaYtbj/2kw3AAROgeeUS/MJ7mB//e28HfUlEF5odF5d
IFWzDxg2on9Pjqfl32YhlTz1jBbCqxd9nFA/UxaV8LDYswrvlQjyR88B6CdH
1XQ8NJj+6ScqA1DYF1fSI0nhSK85TwiSg/jPsgcqEsgMz0hRAW3MUK4TwJD6
Y/JNYpKK9ORueGRBd9bGAbAzzV/Wbj1CJJXorg/IbbxRRhmvprsImRGSsvnl
fbx6bVPPxgGyAjdX+GT/s2XU3+YHVLZ7ITClTWye93mBeeQIVxOuY/REgZG9
ogiT/NlXM4p15gTLVEeA4X43u2f9XX3vgWsUEMLhXX/GIbpIhLko04jIE5tz
EajOWroVY8QEePi2GRuL3e3ngsaqg2dqSHzKjD8sY9/DteX+1/koLqkKf2JS
kDm+A7W+Y0yZ9bIbRbqXGd6tTYsgWY0ABblzXgax7ppVOyf6RrXEb78xgj6y
1Tg2lWnVxCKEHTm+idQjB1QSaQytk5rJSoQ+4zHTk2j66eEqPqR8qxgWudyx
ffrKkIRYXEQ1sGlVM6k05FOcxPCCafUj4vgVPO4Ik5GHtlHYVS6zFZi4W/1L
xm/DS/RUXwSHksYQ7Np6dHf1QHf/yEjViJEp2gH0n3lm+waBHVVil5kceGvM
ncLzi2HDTAFN2E5z3jn9gePpPTOsJznUELA0kmhcdhrOnKtPBu7JZexmvjP2
TrMtTTCXOJh2ZUM3jAaaMrW++VLaFLBSwF/qtrtrkTo9iqagPDP0T4L3PzaE
rYJuqdK0NkuvavYyxiDaO+YcMfM4cvA3RYTMeITQrKPvILFx2GkG/7MYKhEb
8Rg6K+6EBS2vsmNSQnSeUdcVnbk69yfLqJQ/fdRHzIrdwMhzj+vS/ugHrzVp
LBirqDrNRfwzQMeXuqcN0jdjl6kUqxMKw0KcfkotwRq9as6qowspnivsu1rS
8kowOWPXj1mX5RbtzHwZdRY+2pfo5XO7we380Fb4e0xCKV3CsV2t+c2uhb4X
/gGwH6P37K7JJy6hvWHuDc+T/cMu8IxDL/mUo5APTCPFPsuOqC4UxGnehSI2
MXKmbl+fQbTELlrcb3E0Ta0jx4pwkZEQWxt77ZLuRZ5Aw0puDowdlqMmZ0ex
wu9lsfHgjT+47CDSZ+GDCSa8/TQayfGGezxe7rcVPLGcFsaaGSRzEw/+NeXO
40z613XBeWicx7ClSOEhtosF5yQB2/9EHajeJErJMiNzvWNa8izbm1E4cAKL
7ro1zO10iq+pMhOeG0xAc2M5bffPsNH8ccsEIY8XEyVKGOlbKh3CX53/x/52
qIBsFKH1G6h0nKBSBTfHT5zK/bfWwZEk0Rb4DMbr7/OOHrOh+qb1bOuaGlEX
IuZrVGw5Dx/LUB9FmPBXRc2HxjPEo1NNhrY9gB0xbko6RLPJBOo661xpOkZJ
vmAolLocCSAYsK9I3CpI1yIE7M/0/a/LCpXcXGoQAGsonEqtrOdYQCltd2TS
wX1CNkGvRG1dCikYq2WuO0NwU8KYPupQi6beQSc4bm1RpdH60U7C5f8zEsj4
rtLkqPu0LO3XWopu1oKBIvOXEJhp0CAMppYUb0B6QSuJzT4Yl85hAry3bCEt
D1bh1UpqNHvsT2UF6TmMUQcA8H9IAZiEQQdHekbMFtHDKJNK1JmZH1Pq4pYF
HnTW8HXrdYA2PEeSjUWkKFcYV6BaA5H8553Ex1YnSrZmWw6rKxlOAZc1Kdgy
ddceowSyEH1hN8KgsmIf5Pyv+yYuIjbcXJm/Po4s1lLAz7aPXKKTY6F4dQx6
+f488Za/zZb7a4LyJN+l0vDUL8IUt4PQGfuMstLxPKAeQNvEJt4A3j+qAOkS
F+OYO0iFkiODKavWJQRYkpW8SwlAt617jyqwGEKC7fUzkZwLNNPmlUuFxmMr
j+FUdZmtiFfqj6q+hlFlZDHIm1aarRfTgP12Dc5H6Fcl6sMn+OxfnpK8Yfwo
7XGKejiKFfhLDr0Hdj82V7dKAFaubrvz4AOyu/LldXG5K7wTYmrKzh5soFEX
k4Hhb1b3a9Xx+koQrAkNgeaRViuDQQatCouA5ACIfpZz8+blmqcB9wgBZyKC
4BOZHl2d0oG9QYhZeXSoXpu+W/zJKLyKtUbYwdsoLw3Q6lict8wt8FPrF2CY
q0+7Cn45ga4nOtAgRZnVyKkqYWYsRUWSdNOcI565w9inf/QE31JhPdq+06/+
E3ljwiyYt9Ip4U4JcmClXmh5dHFX/aNMhJ1nk0jOVi+/y082gr0nYTekZPHx
giL8eyweu+SAS8M+fmFwdqkRV4pzPCUnyHmAw80at9H5Flxb/7uF2Of6ISTd
vwJVwFz0F6UMo0yXnVpo4OGomDF2Q4GHQ/7HHQG3mRJ802S5qRC1hRlBoq/s
eWGgBtcDNsmwThG/Ow3HcxiKtlH+qtF/AyvAlLkdbHKI3xNCwPlUZWWtk4nk
RfD7636JUSXGI0vwaNBUdLL1dDa8qeEYeOHThZgEhgM9wdteCjLpWRBGyIvH
dxyYyM5pYrZnwwoBPM2E1W969OUcRxciHAAlsahcH9Wm9/7KzRkGpAp1SQ9/
FVo1cfdx2CiZoC1GtVf2rFuAAyS4QRnPQBvRp3+H8ybi942aBjC/SmVG0W8R
y+h+v3e7I2uFPxYUvfXPCB5xJhPwDP0ediHney6LcqDP9s921DR2r+zo2Ev9
dkva9VXELiXs/O8vZ0J9KcdpZOoT+lO/twEu9DsPCFy7raprjjbnTOMMeZuX
+MlzSQZZModkr5/wCRmMQav0cvz8kQdmXEpeE8NKQTLLNcRg1mAjzThS4nHb
NeGnHqnjRFpWRAj9woYv3Mo8YWbj+pYmm7GK5wJZg6jSlr86lyKi7zo0m4Ih
CSWIzrRCg/XVF1QtKkgYlExkQwxDX603sDCmK0w4s2hlGDr9dhOtTt9oaE9g
Zz3XOYyhRUHaHcMkw2eNBriz7rzBwMgiRFJHQFw4KFY0OjKEaE1URANpzGZs
X0+YB8V2QnruhDzAg46KPhODN4YZV1Hr3VSumhoNOKXJdHIq2er0dAkJGkXR
oxLiOcrbYxZMZ5YobdluFxRci9bXmGuOyyPhBowzwTiXp5+wV6SZktOatQiC
VB3XW1A6IdBrP4ww0ELu2xAG1ZDlLvlNZCls/itl8x+PZjfk3ob549n6je1T
QzSPEUGe7XGuNd66xXEzeSjNMW04XVxOT5L5Oz+9vFQN90VCd6VcpG8b3vSx
oQj//QugLkxXxJiOSmpGKMkMoTmlfotJ3cw+jL6sXIQoPUrlodO622uqTFsN
e5Zdua4tP/7nJcAjGfTzadDvaDo3+54pBC4BN4hVyPpPAHyZ/xO6GIzshviU
tHgCEae/R2HP1J2KfEEjbX93tunHxwpcTJbGr+CE0R2nfJTdx9mWE47aOLbb
drVOT+fqSZc1mFq9SPP+J82VTxD6WUqZT1KEHsfZY262wJEZnRpqYPHP4fcU
7EeKStTeIX05VMYKbjAhSBertDGqmglY74ETkXq7/wW+sw+R+Y4zadsgs/PF
rIN+kU7cdnIeVJlSNr6LGDw/+gekZSW0P4Tr0uRmIyfqWPHA6jlB/YxyeTXh
idTE9tsMIrN16XqJL8iGepgTXH7wqVN4PfLIymbo0to26vbzRMIra1/L67io
zI0hH4x1bYOy9yH/MIlV1h9usWDiR9z6i+BE7Np29P/yAqOGdJRYWETt0xlW
s1iHd5ZpxxUPrRai/+nwkwFh9chLFuPxEvKCN5+vnuRRid4c7jLSIN3uS5QU
UjuPpeZFMYaCAsvGc/jNzdVH7+q98cKdg78nOUdLCueES8l1+Ou6kKE6dsTS
SKLrshVkUmtx6S3zaD823vWGvo6kTBlirwDiXOz1wxComWWOPh4MiQOtJO67
tZe5ENWebMYc25PGe/eqGZCwK37NPrdpSn9tMV0otu3xxhvNKoasXBwN9nBn
Uec1n2Pl5D97fAE5VE0nf8OYWPJksu8W7wYJGyE3/oCwihmOEWHV6VWsz3Ic
lyOJzZuHgF3+9A608TgsQYUJHAn1pAzUlQM1qC1XpnuYerlzPiszGLekCGQs
A2D+zQg6XhuO2Q5nMKBHDBXTIjg80AMKQlp1ysbnyejjJNUvW3Ne6etcDQ75
XIvblzTwGcbD/D2lOVxiZrH3ZULnk4KZIgx63rKagnT881AGUPmXfQLEOEYe
HRNtzJtBXdhV0Ri8Jaib+nEKjjO9ccAS/SV+DEDZE0BXRnpeiVSlAwaeEoSA
LOOVIKw+Z1nqeg0ZocaK6UjnZuzHrZyfPKG87sTbb6/60excqGzeN+LHxSiM
L3D8ozpWBVGgaymhvUbWIqUj4UZ3wXGG6ZzpVDwxdEFZ7ew87/bZAkYr3S2K
8OsH4aDCOz8Ykwkp4dGgyRnIyizlQaF2yRt1kpE3KX4MaRxUIHNdsTfJ0OAL
D43nIADg6hDtOadgXLDvlDwYuO3fddLJKOJsJjrPnBv6lmsQiwQq8006kQ0G
AnQ3zoP9wpYNPpskOl+rg3lx3/BCw3ZKFQzgiPLA7JQ15i0QwtBQGGA1s/8R
tnw7NA0xhJlxr5cIb5++Xs/hPXJ/FabTAMMu4m3PD+b0GUiFs+73LLORVQx8
671739c3VO+4yXYJ1zaUqISttSWPSPhuzimyb3oXMkRdvT6D4w0H6dbHtl00
8qwfd7LyyiPmXaJ5U4lhg1og3c+tp47YcNkgZ2Uw+8jCrZE4xyjWMW6DW53e
/d7PmimQ6zqVvnoQOZoZLh26BtU30jIIPVvg7mBySH0nTlpefsLa4K3a5Rx2
txnD2V3mfOTqNIgVSuZE+w2kUkVSDu7ALo9xDaQZQqI9zAW8aU7/pDuRcJkT
tKh9mNM+fEilABy8oxZVrpl+JWUocPBuYvz0Bq3QbozqwXVEU8b55b50SEO3
2icLkjtg9oa5xpp23yHwiiqx3HpSPENTHUYotemGgvSyBz+JOsi1SqXSW7py
uckEvZEy1ubVyxTmg43e/AHR0CrSs50x7X+Gx2NQOhAbyZSHCC8Wy7b4mZOK
rq4VdUV4/rmXm/PsLEThqzTwpyfzPUNywHgNk71Z14xiGIYYwVm32YFrcqUq
P8LXipk5hSANZozDawtbQKgCzKVsvg9JIzBnUh1hLKjS8puBlRc4wyMZEk6X
ISaLuhP0Jdc0fjeERFXM2OaiZzu94Yf/AQzFATS2uv50EdZ12hvYLtv1ZtSb
vDqgxbc5bB0hTy+Bhfmj6NryM9oaT2e2HcMh1fIKvYbNDHH801Y8mZKSOsdE
OVGYKAqh28nJaDOe3eKwGFG55yfBeqQgHf+MR5dVIaoHpRmjt0LtN2bIfRZS
5+w2iw+SVRX8QgHx2ON7vRhJy/hQA3FoTx2iI1rCdvhImIYzXNSbKMXJvVmS
fGM/c4xpXSfV4PECuGGMfKmaKp12RFh4ilhOzBTMl9DNaG3CdOFMj8g13jJz
cJSHAN2UkfiBAuexaNKtG7xcxzGCugAUKiyjuianmY9+HA5gmYAC/wrwRB+/
IQ9X7rK5nZAo7sGXYD6/S0p3ISK7BO8YGr8+bAEFcn7J+UkMU2GGhRHWc+xA
HcsvfXBzuqBOEvHVgjNskad5MeUJDs3p2L0WTPUUmqQ6yMqqyVTVmBYTzGlL
DwaBWnXpceWbfxx1BYD5ZxNxb+080lmVUvKMz5AvzgT4mNHtbI8IYK8a6rdW
G/qQR7hR4hoNZxlL6tlVwbYJGeotlb1wGiUaJkfe3ldH/ghQ/Yt4YjrcO+FH
YbS3j9qvBjLfny/LWi9QLyDEVuNDWh4e6TXVlbLijdjX/fpF+Q/FC/ff/EUl
oF6jkojGhFG4Nqqx/j1db67B8uPhS/Fapm7Ry4ki2DVgI7xGQf78srrTlLen
LiUK6upGrF/PDa5ITAd4m2Cb44kjOg10NNIQfwBkbBHhxCNGJgkBOUlsJr8J
U5sNvXrF/jJ6NTu27+NKF4/j2AV+oIxFHuPQ0npmZvYHsbXHpn9WjuTztLqp
4zCoY5THlNPvCk6SckXfNwCesdlaXqDVZ5ofL/P33WDNXh3Gytc1IAU1BGOs
t+uBkgTLfdmEconXMLzE3CXCNyIg5JRPMFYOG41l9uqakIlOOg4GRXtYV+BG
4aCuh21WRtm43PCgsN3DxYyXUL86xwWnC86Q/lntYY5dxpIrvyE/KFDeploj
g8fLGXStt6rH4Cpb2l5DER9P1OQP+5dCZQM8zjAeEpddpD0NuLLoOr7BrTgH
8nM6QiW4XT5R2Pq+HbzeiPJqjWp3QJR3/FTQ83LgDOtRs3fpu/NoXmVE8xQs
1xD+bN0rSsutDMRVPV/qdxG3WAurVLrFr/q+7QesX8X2ILve22whpC/Jw2ws
WIMS7KYIYLr9BVzkOe03nV2p/H6hejw8asS2HgJfNuuVEbzVSmzCn+u62N/q
Xri9L+KoVn9Yr8O+vtKwJtEozEsHzUXquwjxTuh0ALrx6vQLI1f1O5TvessG
/A5IyBdR+716SthTf4VpClb5gB+oYookJcfncuZVf+kdfbHLgqZvlnbg3dSP
tJ45QKAPHqtHIQGGBRVAJJnJjsDwPEZfv97Pt1zVZh75U8ZiiMIxa0XT0rCo
U3G2oNQRSfb4kPboxN657Y19qE6GW4ce9MNvOJ0OXvTkyzuyFoT32c3Hitad
OkA9OdocQE6SE5iRdcvyGOYbNPvJ50tY2Z1bsu8GWHEYX/KRvSMGxQlptTMF
pjNRu+UkQ01Quwqu52Y0d7fJVaufYtvqG/667AyHncR/5Vf3mmbJxeKFpBMi
Ezv0xR8x2M78g5r+iv/9vL0ONSIpcySMMf5XmpCSRrnYAFHQfCb+kUtOkPAg
W2+a8ACQJw/a0/4sinpbnyruGoFsOzOKqV43Nz+7cxY5Y5Ek+Bav2Ysudiqt
vAu7B7OMRDizNHQ8swIiXXSLQDytgYtuCp9nOq61g6Zhm6cOdWUe/AT9oPpH
GWsQ168+eGj9opK6mKfdzjAHsZ0whCwgd86l2ScSzaDuKEGrrcFup8zWMWfG
tJ6GV/ctCCHs2QGp3IktmNfW1+Ie9NfHSuMyswkts/AZNVNv/OGE0deUVfD1
SnhQ5BxKwrMPempf2i/YPoTU4zFEsBrQOud9Jq6gRx/8QcW72lSQBzfkFWyd
P1JwQ7/KiDGUXH/6oHZOoKuhUEOPQlRdb79aVHYyqY/DfH8ryUHXhAVfRDdw
qB1+0WcgP0CEkRlHkZBAK9nGHXmqR9J7l2IVrxNHDOL6dZp7aAZNYD4m37S4
z6snAoDz09EKmh/LACTyGSGUVd4b5HXmsRL5DDgv/lFJSoCy34qp/9gcrb2t
W3JVtv/1L4dVmPD2xU2a2EM0Z0YxituSOE71tCauW8XRGSVJpS6nXcHwkoBq
mulCjBF7CcmkMMO+Ho3Q7ijdllkSDZI37Gjy5rrrpi8yLCX8RZbj5zNV7Y5P
8DdVSDLt+tCcm1pNpy3dF48d/O42x0EOpRocjb2Cim0zEHH8lAqW1gTPwM9p
4vpcsa0OdiCWkGEeo72/epOZ70NK0KFPSaU1pbegRNQCkbT3wyGqo8er8nQJ
zSBRuTlVinFuWjQAQHs3MYD3jd8TIz3zXiWYGTdmDdfNCvWdlxbYuAp5PXWF
ZSUWRk0TlTRq/2QEKdesr1i3zB2BdZ19ThjuuL2fiQ1RPxd8t63rqSUecIaB
qOLI6CxCEhCF0Mx/ZtyxjuQXzYnZ/CVFPrLrjboYEeRpaXCA9LJM7QPQpqH+
/95g5N51kMnIo01J+YI8p9e5LMhyg1QL333kljpx3bTrAUBZHjpRysoq+Mf6
NEmZsnIWjRc3Wqw+MnrZsTji+ZXtlzRn0Bt3d3ILV4V28uE9Ike0NfHpDV7p
q233CUxk0y26odHnwMNWDmE522u0h1QR73LHegKzpWAWso5is+xjFLSdtbR6
w5s1ihuey9M97Nu2heZVjKt4ZEREl1XbafWQi2Ee/WtJUUPnVvLcZix1AHEm
/wNduW8ikSBizFVqLNtfqyyezzBIiYZ7tZMgprks9jdvDFP9KdzuSOQJUA3Q
j5yGvekqvQVXkyG6vW+EmYyptU7gTjPf9GUHFB313vW/yUBExGPTj5WTmixk
PUCut3+G2ad6U85YrUSfwco5YmPRC6AA3rY7joXYXG0u4MOnpCTSJEx9HTNl
rvn4CN77QqfyWhu3bbA8NvkY1siFA7i06SEbrQ7ilxRf/olfAPgoWbU0tR6g
tc2DjGocDJyHc09qJkst7/U64pv3jhmyWKyfXi8/hokcdh/oY0A7x00DBmDr
M19q02orqgbeDp14rUa/zf6VJWlYgIMYfCWS9pLi8XsFW2I9uh7wcRIi6Wt1
P73J2vy6wrLOb2mnnMhaFEGUaoSz3jqewgg2M+3UiW9F8NS5P72p1ySEKMi/
WeDMnMdOj21hge2GihEK3puMw2Qf/yryOEIRoD+R5XgBjro9FLau9yerRFOK
Izeg3bbDn4cRCVbsfZKC4y6DOx0hvuiTSO4SflYz83IHKJJlaHsXfgqLIU1U
vslECQ4Jz9XZkvyr+mzvl+htK+gARSOxHI8mmOajHSGPDPx5hfnXKlZQmHFm
WE13Q/WqaZMl0Sm08LVG5JzlCQ3sn6qEIN5LGJs9NC3DzWjSpHpsWyA6QkuJ
Len75O/pOpcQUmIPxkOLhVy/PfsZnV95zTS3eYHhOy9WjKdQgTquzqvlcKOi
e7mz3JGGePnMaGQV9UA6qsMGG5Y4qCkxB4LvK1/ufo7gfwfQXPihO+rtcvoE
ceh9aY35220J/rSpNTFbCtxjntemJPDLIFP8yKGjna93db/o9AC/WDvHCw0f
qzdR0VhpeQwN/OTfiX2sGPpGC/1k8huTur6EVUFEGsxdbjRTTf0xlF2cznvp
+3XAIcYYN69HoDN694zB3HQ9Yw78XB3Zj1KhqTPkj0Wz4OzZ0jbgW2jBgIca
YX4IrcImyiVcx5Rxofjk+3sZHyD0vt6fu9Bo5nh5BeguNcer1WN+hDc6sF3F
2LuKCBBEOt0N8NoUrpDZxjeUPWWwEv7jxI71C2LHF7h1GeAvnT/pPycmhwpJ
fa89CtmHT6HcK8vNAbnTrGQYWd8M5yJhjSNla07Uh6ngGcpkYKiEi549+K20
Smjfcw0q+GnejWzmDAyaWhIYBfF0QuAAc2yzKayAQk56idf0edV0XhiQstoU
Ohp2yLERO48pa20+HgKiuLsLCCC0VopFAxhAgIVIG4sl/+95PAvr75wKtGrs
vd5VEwsSA6+0qExwxA46eM+Eynx2guT9OHmU5ZYIKIuqwC3OVp5/fA65Q8wc
OawYrz2bz76da2tcp+JmHc4Ijhv8zzCPyZ5oG5iU749acAi/1eoOJBMRSUfS
P10j/FhWJDDnSPdLKi+XddaxN5ziypOfc6kg3LC73jzEBiwqy90ytiJQydrU
K/Wkp2/ZkW1lwYbIIFAe8SS6VBnHi098GkV0aDrbmsftfBJZEmyW0v1Ul2gu
+HjMyH3Ia3HuAVtjeEfld4z6STmTfPmDhmhkzPCP8sMBm1yYg1bYfZObz2D3
N5JqRpV6w9lqcdIGqUkYC+X91OH9Qlm8lhIQJaCXwfZzlWIYe1FEBlzUw5so
50jZvQ1sxfd5swyY7RhQeegFtNh6pY6Cx5ZiSH/QBH6pR+nJULSsRwXcCedI
0S7JOEMGDeJG41mJNQXzX6MnKmQYSc59Q4lMfeFzXPajsufhYOt+FJZuw1Qd
D1U6QCw+b70pfFnNzu3QkAS+LUJyYmbGnlxpU9uJXqhGYu3znqjTLzg84PoU
VsWPxZ21eYYdnwKIgtgjCzH5To+MkMYkD5sLNBXj22Pbng1yP4e+wdVdjdWH
0mllE9qbIL9vyPtLz0HjNVlLxz5gaY9URnE2awIBmTA0m63YHt2R4ytPvZ6a
1FOlWzbrojKPqV8ZXDhi99h9G36vuIm2Crs27I+I3FGMBuQyKkeDBpQnvQBw
LmoBTUeV2GyLv5x7MunahbYW0GwyUQtLAiZeRVxm3mggR+WWPpx9PTZT+VA5
Ld0sMDz+dRwbtQ1SoRldFIOM2J9G7PSE6wUIGN3ZfkT+2TZARA+aHax5jDDC
quAVbSst8xnVohy0IzujGQnSRMM5vL420GoGubcdjw7Rln/BCxVKmG3l05Et
vaADGOgAYjc6XJuWNDD3ae42WYY98jerdYjILtcdCkMfY1UPm4Eg0yQqt/zs
zRcNSyNQy3cAatL1JsjK0c6r7qv4AQDDIbr4XiVz/7O7VKIEyrXGV14EWoAp
IBGD42y9SwGt570uuZO3YIXeeInWhevh0dhCFC+6LuxEEMTO4O1ip01CS2vx
BOPsdqcF+xuCviYpn+rwETQ8ix3blpPgRgc65QcbImwpvBMQ+CA5kCaQ/9k+
9i446hvc1ntRd8YqYf+xjrNqic8UVK4kHPYXyyngSJhhl6smz47nxTnu8HSi
XR0pvdQx982TLfIf/9XweGaPITmBbBryhgsnq+4QDJ1K+4XdYAOrlmjJHBg8
VPgn2vjYJ/XQ/M1GvzcaYofDKYvQPcENtm4u5rnb0yEGcgXiNy2IDt4oQNyK
HcZjcZFPQ0VqnpsBdZpGJ8FFgPS0e8hmHiOVkcu0UZQahASFvS6bv7Q7B7bV
ULN37ONk0NzozJrjiIVH9thmR0KCVRHTNtMtosEmDAJ8bO/VEcAGmojh7P+5
itItO4CHKGZ1+0dcli9IUzy8LA6iXdL512P9r2fG7pzvOk8FiLaqtXPvMwoG
0P668PGFh0Jr3YfVrbVwwVCumpjjYp4IXy2YSX+RVcRtf6iSUit24mdfYn4P
AA1nybhV0zgIDuNM+KaHOrrfqPCi2nMiS9LCcTKB3d1j23FYeEzK8HnxsbBl
5i3boozmU4S1yqYbj8BeYAVs8z2a21Yn2KiEvFUKQSo8bYbsiARy6QcjSj6j
xk8HfdV3dioZlFgqkOxXJYLlEJE6DdukDf/mZ/9J5eWH6WC18FtE16mY4Eop
LAKaU0dVNYrZYdDSEnULAYhBJJz56IPHbc8fp3NKZ24Gs8Y87WIS9S0NlLr+
A0Tz4pKtevmJJv1aqDzOZPq02XOqq4qNoht7aAWL2YTTbVXxEq69tAs0852b
D6uGt9QoBy4tG7tAN4UUvL6rmUel6A9CMMzhms1E0W3ISp2LU+sUZLEKO6tA
SrupCDunS3yFE8GDUDAnlEdhexCrD/zC1vkjHk3pdnuHvIxNjzIoHTxzLWXO
0CwzVz8+OkbqZHCnUNbLS+Wvy3BJcbxbNo4M/gRIOa4BH+kV76xIj4kE86ZO
XDT8wQPGcv6T5O1VFJO890ltlSxWcYl29MTNLp7AGKC5qcbwTGxbxKnPr/YA
lWamk50c/I43jKlOp0Vv3r+alju8/dQyB07l7HYWjxn1KQgCgwy4cTczffC1
VzHJTfBU3dimljYmeAUaPY19iEEpYVB2rWhcBjq1XC2C8XIeVucSGlY8xhQ1
c/2ojg4A/jhne5s4QedWpV7DMEjzoyaOV6d70IN19ceBfigUgHIRD8WbOEBz
cJdu190hosy1HwGXhB1giiiaOAfb9JxnJeXv3Pu1CzmKJOzvmpFfCi9KUlJF
M/fMTvRRXTLbUwX0NHx3B3DWKi0MVJI4qa768fp7WhGmETcV+s4sJtmoCi6E
XUx+KZRXFUsV/Q3mOU4ouFXC48zVQ1UHyJC2ROW4S/krc843yg/dI8Q8D6Yj
4M+3LtX/uIoi7ORJG/1hKi7w3NLm6VyUpSKBsXV9joY/h4K+B1jqLtgRHsHi
hmAfytnBztFGr9ERHcJdfQWboWNywK+aiLg/mFFhfPV3uozTdLb0B/5L0KtC
l2n4eCZEOGZL9xhS03ZHwgrQbjeWJZhRvt6N5kJPipCFhCUvJ1Kq8lCW+K0b
3hELALqcMnhSJITkB9a1cOJMmcYi6SvdLJc+wyYSh4eqmdKYyV1UkVsKxzan
70FB6oijOXzGo5a3olNbBvt/d7nz0tFvYwtOYY/MefjXqeZrmBPT1YFbjp/Q
p9uMUn0cYfRiQEtsoYPfPMKFn0xyh1iZzqSz/rGtPuiGVd93u86o/qW7kRT7
ga3e8RZ+amW4636jRBcP1cQahAqc1rwSukvzb7cHxUzwsLdLJ37Gv9c0iven
XQvN08C7vdw+NCzgyaKj/uAOg3JXrYRhF1mOl7vavOcov0FmzzEIyTJ8y3UR
SS2HbUCjats3yrrdbsXCEoyom95tAmcW8SxvkilDe4dRAzFncJDHSiKlp0uZ
xnJt5mQJwEhuDkFwww6ICv9c+s8DZ2TQDQSDcPYEmVrt/Xn6aqFcKXvKuV0u
casXT3eqgxx6Kn3DgHPoNUQEiKvJT5FnXqdBDFMSWRRstXKpAEse1mZy78vx
YHF60u7epwM24WRnXJCxMIxC4U702lNzbYpMyCuE0S2e3tQ2SsPesXrSHEOT
WZQ+jfWym0d3QGxw2b8oEATwmlbfBH2ofHJhtI/3u7tn9+GMsTsbFMu9GDDH
4UA52RFuhjxOhmrEtwJCAA6/js5hOSDabNdGkiwa0EyWjqyQUqv5FviED2Kw
RifVQu4f6umgv6VDcrSUqDgDWhfZ7tOG0uYfQYA2rTNhw2sCAl/gy+l8OxI2
IPnsLCRTu6pvOgnWFWUGpz6xmpY/j4cfDgoAV3k15AUaEcaDE7fwW3OXc9Z7
rQzZadt65fftvL9/fP8wAG9WxG+VLWO9j5aKFxoqOtsTtXvgEMoSYfUgKFz2
Y+HG8hXQLnHy6kXMBkzS+D9m4tN8J1ojSlDYDlxvArfOf23fIMqRqI35Eq/5
KSh21ErXntBZf2t3AkSjadO1briEf5uZ6T+NhuvSO/MFbpYXo1EFvU/uH2BT
oySA7W1Z65TyxedLSdQkO8OsUND4Z/uXItJHmO/TFjiVPlq0xkrEYbzmAaPZ
iG1YGU5YWd+zNlPlKfCPRtavy1kikgP1q+rhbKCb1Tr/eLYlfFAV4mZ2bv4b
Vp73lDZXV73Hj4DZ6ZGnrD6dSo/TtIxrVQ79/DXWSjTkSFYzo98OdhEtFotS
J1MzQDA0m1WNl0g2Wm5TDPDDgtSVAmF81Cbp78jSXNEowk1vSPeu7TqMOs81
4WvEmNtmInDVJpVehgEEGu8f9Ulk1LAWzM1YUubJifAZhA5XCiGsavxHYuGv
1fPYuuxTC5tNY4DeIvfG9A+BPTGRKe0KcZNSdew3PG7PZgbdxMIzcVWcTLSq
n9m8mvYMztPva6oJJQ7JDcM2OK0pNLcsDLxlMT2T5M8hG1wHqL6llsmN1gtE
i8HdzN0WOqnoukQSrkDV3s6cThFco05an++Ut89e3KrFPrXDAC6Iq1n8R3f8
iiAmiLX1HuuHRK/onar43YbUjdtAohgDGna+6uv0SC8igb0+feoOWa5hf2Du
7HQbzf7Gbw5WNkEU0zDwsbVKsnTL+IrqsZe+152P5qB6I/LOaco4+fZXSXYc
HGjLzIR8HzobY8AsHGtKkfchwn3HAv4NhlNBbHeB+YvjdTl80UUIZJrJPjj8
EAkQaCWmUauLuOk3xGv17rwWNszYREUR9WAu4RpgFBOJAIRcORsuzUqA+bJo
0Ews5H22rTP+ndQUn6RuVLHmMQM+EBiLMbgLHnI8DNaKwQKWcjS09+gCliQf
9m7p0kkp00QrIb2XogZnzSnzaZmrtOiVTWyjB3obxhRp9/jqkH8r6NCT9lql
uj9xlFS3/wNyVYlS8/xwKuWnmHhVlJKpawdcTG4X1HKuIcm1eLJX9eS4w6va
k/0vUUiRr9VeSfawawEbLqzH0TWuAW4Nx2hOrXRedilC+n1VuE1hGNg7e2mF
lXuBHPTVsyVUp3Bg4x1cw6Sxrh5wxE66zz1VRnZREXrzxvqVLzmr2rLOQ3Ik
Ep/n2qmApHWVMkshUMnb/SRl1PKjfH65vLSxTtP7BR/zEu4UhATgzGldbTYG
QDiprfiAgdOi/6LXqySAUq7R5gmBYjP3lgLJ37hTvwFefI2D8sZAL13B6GEO
yVKMGPNNl1Y53WKro9bWPq8T3i3R0Ik4oZSOaMxrSPvEdtFLEI8BbPvF87sE
jZAw9m6kMqvXKc3+J75sS7hUuRPQ1caSKGXuLUCfqtVkI4tXlKUfuRB0zeWD
QkJgMLOz35TSlSb06y/LJ/qieRvYWf4PVErx2bvqWXl4Md4le2oHcS8q2x+r
0H0ExWqUJXhFU5t4RQZ3zMk2nCqlsX0+PVRx4GfnQ/BRezjTcZvyBi5ZjTiT
VYXzIZ4gIhG3mhadAKDEIC9kNVIQvQoZs2e5xHwvEqKty6fAVuo5OW9FnTPB
9/KHNlY/BTdU3d/69+tOdP08HD5Bewb1Q9MCad3+/wqOExJsJa8yh96GadsC
NYuB+vaILKH5AhQtZEIJKV2ea4WAaV5fnCk4mUnTorBoamPm8GzQbiPc1LDH
Wa3AgaisbldoEcGznG90zVjYekqKjbjxxe9urSSnnWjrYw51ws01GcpSUCOc
OYypmyfEpmjLzGLI/cY0Mii8nLjKohp2XfsidH6G0K8iuo5K4F4V3N89mfOo
glxxl1460RPRYJF/VrbJi9wPQBNuMkuHZo60oNPp3pi/BleropWnuUuUcTgO
e6YJOkrLyYKtrspwd4fXYxRmgZMLc7yybnhBswvYXduekDOx0oz7PLS7QGjL
1FdgPtOwhHRjQ7k1q6nB1ehpoJ+UHMLT1WITdUsDq9BkcArzxMp73iWng5KG
AmdZcAsLVZx0rxviSahSXKOwgoEB7nkvrPmGUf6Ld0+q63EoBeGt3TJTaH5+
hDlBZWVUiCWdq1GApiWa/VtbaGzGvI6Rgud8YX3hGFKUFNYe27LrkJqJsAqj
A8m9sNfbPpL64l8HI7FegGEJdZA1gt1sYXnyKjoUES2pNsi8pWVIrK7wHedb
sub3wkKmU2FOTLcrr5FdtOSj3chPUunBVOQRUgpS1y0nOYCIq4fPAO0u13Jj
tUMOfWSQQ+qA+1Lwm9rOFwWbIIJAvhIdSgq7tHWmO1m8xg4+1diMstQ43e36
9fJW8E3i7G2RAhn9+/is/vR8tTf/9C2X3PuTUPy5X/xBYBuaxxENGl4RtNPH
DeXtJsTzpYr6Nff/zOHGpeuiyKeMgxP84BCtZ4IEI++T6M7nWI1KwJkkSst+
Otgn1vaXVee2DdkvU4U9pHMb5CP7/Gv2Ao5NtCqOBqiAV3BQThlLDl632L63
COGAEAVoWoM5LAiSYP02NveNTEPrCAhFUrloMUZUuy6LXFqWlqaOzXXdgXtZ
G28fbYcmOqFB5ynJIloViJntoGjGNJ2XM/BSxFFZxOXnf/3ktG5pEE3oxraN
C2iC/Z6tR8RucSENNkkYF8yC8qUjCPny1oG/19JWJQlydedXpHq4muXAaQQq
/2vtREAcLw7Qphjk13HVg+xwy08Bd5d4V3PNmlbPS44Sw3GeUvY+GB2nbfiW
GV23UWEIUtXdx/+i8Et5HWR4PnXRwSQFUmhV2g8XQpgaPtijuf5D7x0B51mi
C1lJNLmHxznc1LXaK7yfQ7Jlj+Bzv3fonKsi68ktpRIWDK6gzxkIO8CkTbiS
gYzd2aAsYwmiguNFUsTLaIbmEK25UGjyYbcZQ6heYfm81cw7Yd2FvBPloKwz
ArpmchHuytYBLQ7lNTFOcUIRqZjxqFawxHrH/A0VhXMMOW074kmFMgffMOYl
eMf9DqJMXHEI/osEuWkkgeyO/sPYcov5jmDdhbfsBaTxp56n6Tw58A7oMaI5
RnvYeBfy2DctDGZEdBIjaF+1joFvdSvfHvLh5MLUhTEUnA33wSADDkFf14Aa
56JkF5BJN7XIlsbRp7P2xP4d0EnxZYOgEM5pjtY3DXsmpG5CdTLPepR7X0/t
s/v/bpTSkpQ9iHqQS6Ux2zMLcUR9lZZQNkxy1vCoEju42tPB0RLbUoC1+ITp
h2BJFMSNzjQO5Icih4ZyYn7jXxU+8IEfsF1KnmsAyqTNwzWoUdex3QdYz0iU
3bPSF0MrYsa3Yt+KoeggVnv2sGPZkR7zR5he0iIaWAXr1bGSXFgpcnS5tPcT
KjGcFmFHD1FkesSVPYrWMlxfAIdTuyo/xoN93jeYhVyZnmjtiHJOZDIykniH
55vg9b86WXJtGd8CDKWFAgceJeE7iQVusoM/XdzOT0QQzUwPYZ0wd7nafHAx
tI96bdepBTB1cE8Owx0o53t88gTr8MI5hxrXXkF2bU33J4GbVseoz1Emhbcc
Nb4eRRGKMRMypQdepjUh7Rj+lJ/7kNY5HV9T5HClELs/FHm8F0Z0UhSzd0yI
jY9Vc2fIWdJlMnh1BwKN4tJ/mzsbG1CY653VXbm60xkUqCESN1fQGzFLgXNz
pNIAjraFbyZc2FBQznHJV5/HGStq5ZcuqeGCT0VUzBB1l5zk8aQVly2wsLhu
IxEYs9Y/SFqcIgA/fBBfnMPk0NU3dyMl7c33g5l5jCt95kV0XJUj5rZ90xKp
7OVEytVnfGVfZEyRKR6obGNTD0+wzW3jL3t/3K2YY9+l8bL3dSRn1V/cWKj2
9m+lJ+KCXbs6xDLFTsi+FHPUzMVT7qdyf7TToBf0OeZJDc6SH3wFqRVJ75uV
TtEjFYoqC3hCI5cMszsoamrOCmsI9Ma+Ju3xKjMMgJRvbGwNktDkJIv+Jaua
vJ50WfFPYaTbx8QA/LUNgfC4MZBmikZOJ+Dr+FBj//ZJxxt8KVpvQfAmXQYk
VygOOuWillAjL2TW/SXOT4Z8jF941r39BBoyunxdjFmatRvPkTu7+R9L3c5U
pNQF7EznZaoA+yPqohrbPs2Kw4pqA7E0gutZh3MuidnC3n0dnrN0zqlNdyPb
2wVOJkrXw1+nAjBGMDqlUSefPXtpN1DIoTYQ4C4tLt0+gt89tJhZhqmjBWVZ
7aplryaAvLOd7PsMt3VPkIbpJWY/jEKGTB9lOCytzHfbJNXA+Ov4RD2iU3s0
S4WAGjM2b21VUGP3t8f2GPb6B264NJc2P+me678fdYoO6OuEkoj20ATM4+z4
L7dQI9Mdeyd92t600nRHMnGeibwK3c9FpssHRurbyNl9gZGWbgZ1MNI22BH9
D1CxmD+aIhKuAeLibu2BiWq2j1jG7tEc+ghWVR+HmLAt+G0I7kYMow4p4M+O
broQA48xBbOmFWhSYTgEl8oGpy5xcSM3Ijr9fimWA/xxMIB60AEb1Ct/V9vH
SYGkpiV8oez4mPOCo1tmpNUHGIrPBrYmCvgQ3QgzKEF8uMlSZoqk+A06OcL7
MaJlcO4R81uWZ3XZnRl9wKPW4fkQU590S6vFCiT3WJaU0sHokL4VFlgdOxPS
vudTdqYGGP24VxiodJnx32bOrCxjk9aJdhVif10b2RrE/3xSYk/7CXa4gxm3
9ZI9r18CkFZ6uQU+5HEuIc8MeiCOAUqi2NazLj72ctBd8/X3VWPVMp339R7f
MKlnpeSlorz+gT4LfyGXFUeyCqK1SViyPeb9FoEEYG+SMyWT1p+54/Phj0TV
ijP3W2N90KmTvZClWP4xaf4rrGRrmysmz8cr7qgkvvnvvT3QCr+TR3aAxmWB
XGo0EuVArbvpWTmNndeN3km7XrWV47c7Sg5PIv87lgAoX7hdBGCU9Mmpioou
ovodwZInytX6nzP4Z/o4Ckg28qRaWLamfZWw7pFjftaJjOEmkVCJdKglZ+yV
ubkDORVlOqZMp61zPeUM8Dp6BzGPbNpRrFKfOMf9/8Ic81K4c6Qnjz0NdgfS
so+30+2OgAKCtwDq7fbhrBZ4AxhxLjZcst0nVTJrqhRnDMoTpTdh8sK8YWxY
xmgBqzxv/4bM8q7+oWSooLK2lud2qhUNScfieXZKAmG8MINP+rnHlvIBfstD
T/inzubd4pn3TiF+TMLNOF9mVlEsYE9EsakyRAWh03cR6p/1iT0y5PYKzyoH
5vhnPT26Z+hpMinEytZRMC5eOMM5zQ1bILlleTxwgDkq+8/FHmKXgZJSRYpd
NzUnaAYoG779ua2mmvULXF+osmxYimN/w84Pi8Q+Q+IVRTwSTipSKCPPmXfU
2iI2nfHolPH2tB1RVPu520QGN8CPM3B1hyXXrLdo8yrJsP+i5CPLI6rOIZvN
xYPO9uy7QOCR0glA8YgCbZViUGtBPZ4mZHtijTKT5k7uPOtrJY1t2aUk9saJ
6gS3do+Dvw2H444HHi7Ce/64d65+VZyjeitfWHLqC7ftbAPWCbxQSEWLRj8O
Rk1Qf/5jkrMY/fShkprWx7ase7XNxmEZfZToGy9qWxYDwmnEtoDnJ77K2Ulf
8E12vEfcCt8ijuaS716Znq74LVZo2P0B+L7Sf0vE/cYnPgkjN1UKmQELuSOy
0T+O/leqs8YsyPCM9IENAy3zYcqmODlumAtxZxiTfc+NvlgffQFWfFLQ3jti
ZGOl03aw44OJEh7/btjDeDLqdz9wQmDQ7tsSK3RbGQJFE8pzEjPD28yQTK76
ODM9m1Ksgz32LwMHEGT/iT+5YoFBVr/Q36ZXuNDbg5FE4CX3QWRCX8gqT2uf
O7t9nYjiyvBBBxjSTPzJbKaefKWhBAeRpsojGCZxKJkiPYrnn/JeXE2RrHrp
MATP3RR+ooTgGsOJOFAJpZM4DPUS6zM9+LpeZyHa+cy1rP0/RFdiuSfKVr4t
6QhzAm0XuPkSqu7U87Zn9icQmA1D7YtexAg3Ptc8I5B8cKRGtrZhHIQaza/U
AL/6PXiEzZuUhJZ9xEFemPmMLY0hCPgzSHOil5lEGmxqDJ+50OzqJbpi49hQ
7m7jRbK6c7BKo4TQUWxmzZw6wXdjq8PUmIKwa66xJtt6hgUB3e2u5zrkU3f1
v8QbfYZ+MPzJctVuZ5t0pN1vXgkW0URvEvKpZA9XB2Y2lkAD47O72gOwtXX9
bPQsdQ64fLu0N1mqwVTSTIaudvcIqtQ5FFpFMNZpk5CgKYETojjaqbXc3Fdx
fhN2h9erFLokZA6Zf6M9ER6mSTPGpukSVMxGPMjQX3SQpe5k7zuhD7xAtO9p
1epJxTLnjRlY1y43cJW9olDd0KPvH9HgE+9PWu88Ji3yo33OipYeTNaIU/fE
YR3gRWr6AMUMYFXMdjWd8F504Kioz3A7U7bAaIMFqLDQfZ/bteMC+HcBvAWY
/ob+sb4B1wz15IDctqLv2DgYt5nBRDVTeOqFrJl8SfnSb5phC2in1nMhF+b6
aNeD92D7jEli2DJt8BR+092S5DaMQin3M/d6jHbZSiWPQBj19HXe1grXnPlp
VSc8ZXbuRBCOodPqekByu1x+lPtNvbghkSst3SJleIP6BZpe0iZRTfPVgqT3
afiKGf+65SfoMLXdGREOfokfl2rbTKInZ5jc153ce4NrfodfcXldO2iSH1Mf
o+y/i7nr5xaETJO02Z/y8tg6mjRLMl/l2NLzyccbAucCH0LxxnybelfdaJZh
JuWNDGn0Regb2ed1+9MLyY3jOZCMe0Gvb6/A+Tt02YKh5wCmNL8B7d09ed7R
8E88MYdlqahdRn8CTTkzdLlOQO6mLb905lnVbwTQUWSXHriJgRVPxSvCsoGb
k+M5UHKhT6HFofcoGtsXL76GamLW8Gwe+R6tezT1z7s8SbOfI0nBRCR92i0U
Fs7fGvywLkFrDMxU2adFzgWCY8a5SIJIaZSfJA1EcEKJOXw13FgjXWAC73U0
B2zKjESjSvOiBTKDD2+g21W1MGGeqi6KeIfy7Ayeu5dYoKIpxpDu9JA9pMuH
qy56Gmmqm69p2j5WRJo2NcmNySvzhjYPDAgSHs4fM/g2ubYyCrkFWODQ74g/
DwarZiV1Z2pGV4Q7h51+EUOfs8rmDY/B73O1HS7PAr2fVdTHmB25rhXyy3Pf
g+YWZwLZKTTb+Vr1qvtP/TeVxF4wsWOPuWEpin6kyppILUXxUn8NS7mkzvcK
uO5PTXZZ650rBzgAXrBjTVnUS6Ji3DShChR8qxGfs8hNX6Zku7QZo4b8k1lY
DogvcLTb5YRQ3H1QmFjeIAq0K1aDv0a2C6qDFKl34Tegw4WtvS9v25R/x3OD
KajfwQbAdCRtxbg/UELBD6GdSwvPgj1xv/urjgOlC1Zh7+LDq37TY2KnWoIg
YnltPvbcahYzZA12Zkm9BYnGcbXS+O35bFq1+tIAgGQlTUCRE8iAsgULlrjs
kVZELjGAXgK2FxTRDKM5lLVPP3Sf6vAG4aSsXAPvaH+KuACwR7V2y31H52p6
q7tl80IaiYLyUDYOuC5jFUhJNbl215kQ8QyEh4JcwUf5HLn3llAJpVTQORXX
nrUZ43vpLZg11fjsCGSo+snYcKzwqhm1DT1XbOla3XRcH3AQD+X0q+QxXt2c
bNBcBky0JzqOfZ7Xkec9SHUudrbbMbaSIrNDZv1kuFcW2eezhLgNFfmd02LP
9n4J0DfNSbDs3j8IyEp4plDKAkiY/WIfOGtQyH8mqGn1h75I8AtklZltHqzJ
4HmAEnjhtZshWUrheZX/VGnwztbZ34WyRQMD9CyTQIErPnUL62qHqwHGgI3j
rO6qqSZh5vXNfxzqsSmBWK5kAtoiTVMVfHr5V7k6ip3sXpnERwu/25A6+qGb
xow75VESt/gL5tIAlRtqVyKb4XC5WDwCU+kXCNQ91kiVWEhd8+QNprqxIff1
XBb1rJDCz61Y0ibH1xccJn0u77E5LI+sK9kydbOnMHtmHct6ZS9jjPuXrksb
OMYqJtdv5BKCjBLAJDESSLuOhYumJP/EU6hIfQCFP3znXJkhD4i7ptV6FPmM
zAgc7Yf8kMthidupV2LaNg7aJVZ9OsxRiNBVrT84+3ToZL5m++mk/txTXlyi
l/w1pUD4YRj3nQUJ/7SG2qNlSvOdPREmAayao+14nW1PS7FzjdgaIY8w7n8r
wQ/Eo71sZuHw+iRx33kAOpgtT3cp0JgXFjGDtRkMv894v2pBV+wtVrYJDKiB
axAFoc2UqtYOc1hLo/7qAqkwO3mQrzRbghQYFgDmdOI9AxrzjegSj4rY3nTD
nYX5AakfEB4MmwVwR/sE/TcYWAFXe0M8c/IAm4Y6o+Tsv2WHuH8VZYGUQTpD
YAM2mKQXfKBj36S/gj8pkkgsRJulx2KDOVxBwf3YQu1b1xoFPZh9NsjG94mI
opb9w6l61SDJTSeoQiNdTHtxStnWUHUOdowU1tzwB29Re4hp3b2+4XUwueOW
g1F/G+30/trfhv/+WSk3CTvltMgv8hqTLuifZBbYuMtZKr9m+jvxuljVu9Vs
dasL8GsU45FMk2GZ6KUTFw4ZIG+lzrqVF3G+4NczqjZfEGOF8qLNUpKhk435
HZfEz+KkiV+FjZdfmcBMul0lKeNxmu/B84qrbwa6MBt+/bRThSwPqtzHJtr/
CmftQ1TORsyV6pXUc6Q9vkJtumZb2LMeAvdqzoxvYLjj8+L7QutXVQUb49Gr
CrIoLfg+YTrVwapHYnlRItSbtvvWMUHd3IGjm3KhgBx/BMNDTyBtM55gWGMq
nVfJbB+0nhN/yXfqT722dbc5e6QBNKj3vJUOnc62zmQt+GVmIKlK8FoECf1j
qeB9WRlkFFKb/sjCZ4RDxqPRw35BPUSQnKy1VVFhbeu+STJvoWHbf032HnNF
Avz293Ok3cyuNESZI1/aay2cdAPpVljES17PADm/DFcZ64EaAqF/aJMXNrUY
iCh/sGCA5xlZ5vIAa4oMoaqsVZanAe7KPQ/dXICaiLeWT3Xhk1ZM8V5WZTg6
FedZ+hT2S2GoPpURCqNt+Xi/7gvuksUSYGrBTzo0jXfzCE0Eq19CryN1CEzQ
zbaHEmuWII1v+HPmC9cxAG3I7KY1Ml3vPrCWnQcYzXk0r27eLHaKmiqHodd6
4XYzrBobY+9PfpaUvkH2LSuqxkgXHWkj20NI+iLXhgSrdFR66/OsL80ouMgR
Uo2QVUcUdwixA5vP1iaPs8ftcmXpGwUrf1m00rEy/9wvd+LSfFx/t/nyBruz
hOROa3R6gHHb7nG5IWBFFxDzkWXk6tiB4ll5UpZxhCL8ZB6n/GeXzR45MkQN
bg4fcyPFPv+4yQn0eumMBqIGq/Dt8YVK1BGQCnTlLRXSkb5pctXZ4T4mtgtM
NBK1B/q8KyInSt4IKLO0W/V6SweTeuXeMNzzQH3fB02zhSZj9ZGWyqPIIGYB
Jwe1T5IAGvC495PSRNCU3QaB/4f51EqDap5pZA/y5HOvZI6yrcOiDovoMhYE
55e3mxGC7f4D8mNKVPwxCQOSuAKBH/lG5Jl4aMzYyi7/rEWVHmnXn/3nxkPJ
hyjncMCdrUAmoTJ8H2B1Lc/TQD6VT1ohFs8v00NUsUwL/fJwly1CEbA4Lvmf
jEW5vT/Ol3IRId9tCvOxx5GaVto8EF5+U1yan7MjiYYoNmO+RtP+WArIIRoG
IQZGKQDFAnxEtSOqGSYET3jGhsWPG8DL4wu1QZAO4ZKmsyCWt5Ff1QTs9PhD
gcDRY4N9hZ7LCwBjuCg3m8XVkOwiczrFK+E4uOImYhL30POmDDGis3bUtFHx
F2rQQJvIxN1XgZhyb+4ayjkDxbdjIfgMhU8GL/4fwNNSdz2uWTQO1lxFqRbs
kU9Nh2/FOSswvTp/Ugx+u+HjfqYMxOZ9oOJNGajK33ptQdSGtgytmhrvpzWw
lpV0XVavxKSMOrfsOL9sQOhAvqRiQu9aX+pEL74AZM5bQntit3WX4TfdjiZd
65vdRgt3zTL2ov7DCT/Lq7kPDHnsUjhACOdTCOVgozJD0TmaejVngeHGB9v2
HUT4I1eLkcRtNAkRsWrXtJH0ezunbuokPYYqtlLVANipNDq0j4016Eljpi8H
b4gjaa1DeRl9BbJ33FV8RsiWYCfXq0ePujWMDwnAvLH+0A0Az+RrmCSShSuT
sMk5QmZnksYnlW/fcanxFRP5Q3kQndcSg5cIBmnGogHLnEiUZYdZocdsDrKj
8hnT8lB9KHITpMWGi1V6J9DSyyY8Lo6k++pWNQ6IRFDHMdq2/VUCVC92k/yT
ZlrbfgoEn1wlkLDuRaNGXx086xYVvT5O/RdxWwx+wZ2X8E4mkfEf6QTXxJ60
3aWw/EC4AJOm53hAQNmEsHV2wYB6nV1bS3JSXA6FP7NaRBxnM6sM2CaaMHua
6klGepKAH+lh1fB6RXE84I6dwTcFjnAkPtYawykqk6gNCCbT3VJg47sXjVdv
6Xf9FrNzuGLBvBaha0LvqVr/RkVvnjt5e19krj5SiLkoEztm2k1HzIAVh4nt
RnpHkdfJmft3Ob7IJtl/aLPYJ8eMtSZTceh8x5KD6JQAmN1YSHCkikLTgxMD
yZyhVidFZveZmMWw198tOhKRRXwd/ciQqxkq8c5EwJNHJwzxigbk2cyxBzj+
YkroKLqUxA/8M4TtoFpdcKx7KiGLDE2u8ffmC15OerBuLdzo/lfa5edh0p1h
CYujVbli1+zocjc860Uu6X7vhxDm9sm2hXS41juNiWItk6kE2yXtkJn/0ee6
m3GDdEoV34pxe8pdupveFyFqBbpmrQv60YpylOt/+N1nhxZlgG2PpaU5Vavd
LTc8QctGX7JCIeus4wnoju5YWQxBa1dxjxo/JHlzwyoOECaIUqhAjYDbGsDH
J26A3ZQS1560ZEEsVt0c/WVq5VfbjuvqwViQ7/w6f+7CGc+P4IPsQnLKTfIQ
rIgxjtlIGMxgyyw7Q3MakOmFK2vzTLfJYCbM1Nsnc6e92z+tcLAfWesQSSQu
8LmcDErlKQAtm0kQCfe2oQc4UsDhSvQ0EsSej3xalEut9hAjPFjJexUTBbRz
sxLqb1DLbDdUPdCalfpclJXEy/JjtZT6ssnSGmi3WuQrrwiyDCYZMYXqQud5
hOXTRXmSFPczOutvtcEvhJxVCzyLQefIM3OlAyognxcX+v26V4ijutGQpoAV
qehFXvLBMzqhxxk+QxJl1BQ6dgbpVJGRvZFOaiJerwo+El/W8YUtXFi7sQTv
tel31d4BqLa4M8fBkHb8bivTQeNWrw0/W39iyVejGmkPp+ON4bQsXP/sLSTL
ya0fXjx/EYevRE85wOpMTpJs0R6UEZtPa9Yi9SIPpWFrkrTTqvPd3l/WdKrg
2lCXaKuh4Bx0JndRWmztewjR17fpYCsvRHHZ3gPuJN3Nq+wyDCmKWQlZTEBr
XlWCaSGWgD1HT1Lz6lHZKT1W7W/0HD0jJ/2wsPGqw95MyuW1wQ+jb/Pf/LU0
Pwlw18vgYAln9HmATts8HZuMQpSfPAiI3A4NCgBTRJ0F3RokoT5vMayG0pDg
fAfaUXM1WjjIX+DZzF/2cFNPf4HBczurTT5zuJlU22ZduoLg1Sv0bj+vkUXP
e47bZ4hd0A3mrTmFzsfbEdiJp0V3twPAM8sD1kuRx38jbz/fGfdZ7Y2hfHSs
BbYhlNhvMMiqwHnle/MprmzS4YLPL1DYu0flhHRG39QMimzQPv0HwAFKD5vn
HbbuHjY8TjZQ0jYSxSUlm8g5GhFDrn0EwX/152S5uOsSWY6DdFw8JwezmENK
s4VzZ0DFXr/W4errfMAuUfMrajWvHM009wiL1akRcfHlCzSuuKoBAyCTWaf1
6GQr9qBcKgUH0+mRCromWaF/coraGUorrjWptq8Qr9dJkjCW7BGYohWGZ6O7
7WSuo/Mi5wTUtzo5GwaJ4+aGSvkpPH+KvTzAjtO/fj9IbsWjSLHWgLijP0GY
Azu4zwtBhywPxMDEUur+CrBjF9SJDFUDt+YHM4i91bHb/MwRNmv82l+thuRc
zPmGXQ2vPMCnZCGuV1ibY5kOdX4H6dELLpApJ92EnOCUjk0ez/pWvxFbawb1
pDpwBLJiBo2+U4ngBAhj2SuMD9eBodVWSOU/nQjcISHPauPS9O8ELCyPgViA
DxU6CLM9Fvg8qOYqPlC6FvW5unz+ZMcsS37m1pT+tYgP0M+H2qdyqgkTFmJR
QOUWPrF0i8GqRd0n88ipWF8RLbvObq3H2nFf2gZKckhhHPJQO8newCFRztgh
nYpvmgFMJ6hahfjMRr6FoneL6fEx9zPtp+0nxigU58WCL31xHHJx/j9h6DxC
C9exjx486fjtj2cFiOsH5tWv60ziHdfcD1LWbaeJ99v6o7zLWasiHPtRNNij
8H6JH0x3V0l19DlJlwV/3m4qQ8YF4G3I52U3cGgj6UmaoyCzATSHDvcBglrD
eDzQNzqRz9RjIzi0bly+y9bX7vktzC/l0sufvv+ik0VAyjSnQU5YVSFV6OXl
LtcVn7UffO5LQyox8dgsOb682IVNngGeb8fy7l053xd77RuSxQopGNbuxWbT
z5JoGPD+zr0SJ5pEMhIJaOGQEdFpfdlUOsE7YLZzFBBY3q4iCs3hUVc4jgR1
DzW76qJ622t5KiqBnx2Dh6YFxGvDJoiaF/rwc5aro79Sayl28WdDRCD2ZG3g
KpD4V/vS8wjdYV5gIhm+AmeXMTFgZBvA2KtHfhm9ftyXnhKtOA5vkXdAl5YX
UD1mupFN3quh88T57ERMXPdZFkEBC8LnEZbXbXlARJpMgvKSo2K1biaz/01b
yr2+p3av1Y8Dh8w0VgwGYnU5vfsw/TPf3JYgtIXnhOYe6iSDpXVOypCpZlju
qfrSYrstFCXFOOgRGm3p5RNnmbYu8T5kCpPJ9XrXph26CfkkadbPLOvxByrp
Yuhj5XY+ULg5qG7EbpQDBVf9ZhSilMlSrmVxi/63AijcurPo05bt/4Rdatcq
02Zp9bSXlMH5zenXo6H30aw51HIrIqYdUSXcRyfci/JNw9+RMRqMoPDIADxi
Qpq7msElX/rVVffo79DRckN60G6jNEeFZpzzkUnUSsPMggyTT1R+vzF4Sm4A
z202CfeQqYN+tmE/yTrt6nZjmXVBuZ3hl09JMJJL1QMg/DeWt9bXsIG5MRty
7r7EhNeQ6qOb0vIu5mO3UnbBASIDCs1hSLkif/wWx7xsz93CHGT7VDCGO/0g
Okc9YISklPxCE+VGUqw5txKyFrKBD+4ILFKQN9ACvzn3JXVIqF2Lwk2wQXv9
U2RRBIVMg5zh1gcx2UTPmvYmIVSpjH5W9Nup0ekW3+sqR7zsZkrRCE54ApqV
x9c4LmpACX/7e/Qd03nrmhp3Hbbt7gTOJNaR43m4tMMBgCbDJKHjf51j9Cvi
E0yPdJYeETDtxxtTNitYJqLN6+VNF7bzZj5i8xqw3hlY6twojGJA6IJhQVkz
71Z9KqdjzYMOsAxqNsX6qZvr5WvnTwRAZPhC+33qng5JTkZrFrEqSavYxYlw
YYI/2TFkyiAcIWdpOOFzglkIrndakiclpC8EBWwj6CbT5+xgvhLX2xCCIDp1
wJDu925JOgepnCifyyPlE/2s6fcLu9zBhIqxRBQnvJqpntin9FDF2eVI8jlB
YuHeMYOiQnRipDMglNX4FJob41vklXkmWlCBK8WbzyN/KUa7Dq7hh+lgGlru
gfAlFFVmGZL9jbBh1ulk8I+XHyjCFFN7rOJaefMgoChebOOWx5N8YJvLNTER
UDFBT9IVEyk4TderZzdzpLu4bfs85lZEyP9M2M0/5liTAb/m0juhM63QPrQ9
CBUB4i734t68xVsjhIh9uT6bBi8070b3o1TGXE4hmnT7IjU4GNRydXmM1Cfl
ozhz+JVx4iUeKwCrWsakJW6Em3GXqsTyQhJs0jU9nSApwPjwOQm2iz4Z/qXH
m7RG+1PSrzs2ChFVyi9lKnodwxOlfGKaGPecUAHUHd+XeWPURSABl/PtNAlp
qHCKDVaiWF8BTuFlYf+HCY/eUTp0rlfTJ/ZRSHmsOHSqSRojpb76sN6y/c2g
Ndfzsi20xdz4F9xDyHRkBONfmhW/QS3gulagfnDlBj3+zYwFotUvKUewE7f9
QEptUraAYlYB3HUhd6l6i4ut9XliNAFIwmOPa8yyW5pTguJhPpTmIKO+EWmU
B1Y1TcPUfn6d4r7UePndtcgGddQl+NDoIi0LJsXGjnHNVwuco0953DNsT6id
2h5RMxTTw1FWDoH0yESrFiY93zn9CMv/G59SiT0WT9dvbfEgJyXThPtSKkbW
G3JKx13Y29WJd9u1wn7udZk+eLTpU9yZFKdSKqHMfltlGNfsTEXgCI+IGKau
BWg97ukM+Dh/x4hrA1awh49vNe/RMHPJDHjdXAoHu6qFTiLB4gQAzgZ73TKw
0HtE5zvuXiRQQjcLAqB9AsMJ+uVhkOzNqmL09nYsekRVNWEVc6YyNZeeY0+z
0DZWCgJriAdx1lU5Fc1GZ8W5efvlF9VMoYJkLg62pBLkr6qz3L7aiGXiKYur
p4rQWWF6fCoKjXtySYjKhENjwfStOuYHnFaw7GAUl1e2kNbK90YRdHySGfxC
WOaGIwhL/k+cFAYQRHNPhC+I4+ejZliM4vLpuKwpWVIjaoGeuNsqlZTwZPJT
whQ+ac8RpLIOsibcna8ZQ1Dlg/aAW6iDgdG/6QWYXRZVKptPQ4GnDk+Y/frI
Wp+3SSlAd+MB0mrI0jDqlVC1+cmpvyvOToOiYxs35JfDgw5Tn4O0kREAPr+u
BKTbj3ZoZYgIAobeJe7ffsbF4wLessM6YlmduLynnCBr1j74SJoklhQmoz12
GIKqZDgqySxYGzxt1nbA9EbwJkmcQohnjeFJ5wYm+X7jjbCK+0C+r00tMehw
rJSzNnwzr1BNzj80vuCg5bLwR7y/Wli9ibYbSUl1JPcjyN5/JqpxzcHNaQAb
P6+mUpc5UCoIr7eXkzZhQedDJZ67LSVFwX1bOtfJF6wzCfqbCqvGNYeWpFgz
aEBtx7P3OZbY14+rog1xjplYDDiaVQakm+2ARM1qeEy2EoPLtbldTqd8Ikyc
9sShVwZddF8qkH39J5tSBzpd2IjuUnuUlEuhvyZn3e5+r+yBFUu/tvwhPxaN
CpTiWcP2sd7HrimGD1n8I64FwYHoHg4zZs9/0TpB8pJgV0qkvaNLaziW10wl
AfQx7Ys/xTUkas+Rk8pgki4WoIev75tIvqke+5n9buamiynzGtrWltn1yXUS
+QWgzwOF25cg4aOdHLIfTzRBvpctS5LTPoGt+c4k5p50462w+YhvSn3iOu57
9fI//8Z0Q4DJpy5KUu8Y0Nke+aWT8J1usvDhQwXRV3MOH0vzvjctlANAZoAl
q7pow+dAt7/7mlwdZwTsz6THQ/dXARdpGtF8xfkIOl4RXjffs/rYChStRtpg
cNZbNxJZziVPsZ3sO9twHPjW0W0bvHjcv4PMeww0+UrnIvMriSGLCBnWoTBx
umrPFNxZdgDWj+wiaQR2+e/oQmL5HNVkmIPjGKzXFVKaDVep3lQgabgYGrZn
G/VgYFJf/SlK7hrBehGwpmRKxfNiglIaH0gz6cU/ryiCurxpLiHVKwnK2XBy
fsV8mcqWNyQCp0AU06vBXGphjIJmEaJBZFMDq5vuC/VGx6NPLvSBRQVoNYgF
1tCgxoM/eQC2I2EMwl7OhMtph7cEpt/6I8usug6L8JIVMvrgOmBcJ1EsoCoO
CE2BCDmDSTvoKTNQDUsLZ3wP7Nqp0BT64w6AeUmDU8fqJhfygNPgaeXo3fSJ
VPilZYVue8bH97M8hSXEVC9H2gkIOtyuqn+3wTELnHY0YFiehUZXrSc7vc/c
ZxXUZXcqr2jJXDHetCKfKcRpPIxCu/ggbug9ECiC+m11I04Z3n2tQGXFIWoY
BYGvEHqsgdlfYr8shorNccggqaSVkKfxDPj/UW9wcYdALzuuSVZtJuO2gF/u
eaWOC6JKTymDoPY5k+KN3v+h1arQHfKTxEDgqdbgeuk+GLBOTke3N1kP1iCy
neI92VPJ9pPsKnxHcEe20DMmLOXc6GDmey5+0R5vvoxpT6RQ5XTttEQkKrXK
FXsRpXa6pmtkvGN38xQOf1vUPfHlWUL2ptAZ+NXwwFZtJIm695ZrS3VNUzE7
gq31Gx1v2UwFaRU5TG7FdwdNpRTdd8XcweCKH/VQ5MghDtT8L5ye5BjXDbgH
TWOVZzwEdhkiTVaYysRzZapaAotKSP6UtSv6Nf+S6QMGciZx0EUAuCEf+u+7
H3Ot7nG87q32H6TWVrHCO8w8HDFcHePsMA3f8L7C06lm1rkVDT38yEE+CS6X
cu2sVapxOJyuQ4Pu2kOsdIxIWR5VRQsi72WON7XAqpxEHmu5vXmHcuEz3b9/
4kR+fUiYCSSW+373w/CbTY0cyefBdwRHNymplXbVW2PQO/E8Qn9UnKQCFZQe
8M/9TYZoddAM1Pn4JWs2oxTFLfLbFNSy28ztHHoldvLH9T9w+s2d84kKXwua
ObDM3OJ1h0rWv2AEcn6miVw3CtvH0eZxgTo5m5PmWFcooJGVj+XdQjMF21XY
9I+9KXLy9k2hgT1c5V8W4BOA6fG1QKSutrDxA0/3xP3159HnnDT6gDgbKhvi
RqXB33R2kcScvfQY+V57Oa1bPFR1L5+XOxlUj38NTqNrbe3SlN2JI8ZfL6bQ
V8UbvjUsV6lUO8/Rc8UHU8yvLrHQElUg/ba292N+ltMTmRT7VuwX7S9ohA3j
J73tu8/tf/Ocj7mpOElaoapfbrpPNS5MlLm8GOvu7H/m70mvGSaoZ+qB156A
EaculcZuDB92H8/7yDl+IH9Jaqv2RtMzX9JeS3hxiJxysDqOBA1zafRihFcD
BU7MzgFi1CJmZsrD+D2CpDxTmf9chMaY+1RoMmC10N3fw7P/8t6VLLc0rnxj
5uBvaVz6dyTMXOB5RYLSOIHUgQvGajfyQegG/81dNILakySScywF76DTW12C
WsfUlTx1QtWx6UiOZEsSRd9XCXFt32hMiXMzLCsgka52cu6ILVSyT/EqNg/h
K1s35ymm6A4SnOvEpSwNkd0qhaAdm/58r9M5NcpEGH1tnqwiPl2AiW6vlOqQ
J/xlAoPc16f8keplPvdk5Sz8HdgDHWWDXAiTNhlYo8bHp6Nkvx6r7WN+yF9n
F8/TNweV+LvFe8letdWj/kX4N5oeljQpxc3kBw5RWUEV0wMfIBZkPxDBMFtR
5t2ac1VbC7C3LnsusYKHEE0Q3TVQvpAFV9bkSZcUxEBdhkUfTh7p0htp6L7B
yhwfIR4LfMNTxLz1S4zCa5bNbHPGK6iqP2ciDbn8B7ZZi9bGQpxX20d30dVO
BPLHjO4IbAj9AVhPyiy/B4wOTUCDxwNM6LUKCJlj9Y23K59MwL98hcH+yLP0
1X1jz3qolnqN1ISKAVEuD07c/NmrRxkqAd7e8pjH7uc7V1njPxYyjGZBFXA4
6GjSLyPT9/1zxEBIJ7Wmxk2auTYSP2Oq8abafPoBxbI4gUE4ea1HxrTzSYtt
HO1d5vVWkO86f/EDjpFi1+nJkXU3s0iOD6tWBp0QZPJMuglvecWzRHSyCYbE
MnamkHxUxUzWJPEP97Fc5x+fPyyzXLbULPLsrTbuGfYc9zEIKsJqXkNZLSZ1
sgiXVDjkSz/4K9niXdm4Wq8t8Z7sfgC5wCr5bZAbsdQAutcM22Feq6Ogsvdw
rr3r8lg3TRZ7cczXb0d8dniB19R6ZqB1rUD0v7by3QvA4pr1XZ2jk2L9Jjzh
4mst8if/G+dS9ezRDBsXqFA01gmXP1/xYiJqHQWIdVQVIZa3l7wK6Int9ScP
tqu/DoM/I5Zghv+IQOMrOd8kS1IMlvnIUCG3qMkz4IfH0voaklkQVjcEc2Ds
0YXS47T3GuOHiXG5iaVmmcbVAqmd3G1COu4JJ32rVS73+yc4kJVHynqysYrG
l2hij32qKoN22DsD4KCy2ChpG6RcP9c3AgiY9I484QH6j9Pc1plcCDivs/El
mM9q3zzARrky+1eo30AEY1PMDpFXzG7oqFYgEipPvmvgsf2OnbhT+eAS9yeU
xHTqBQHNVASXznMJNuGArOMF4ItMOK3VBKy7nY8EpGeIYeF7pYd0gx0rTyOS
6YVS4vOBYNdo0FdSSZlvnT1l48712h9Iuu1MFxtt5e8iij1FLjeb2uYTT7IT
vh1lyUUkz788Qnsl9wNCE+gSK9K2/cCKDLYgIbbK7ZNVpCt51JVU2CSSMVNR
Bg0pYfGcJI8MB98PNUe1+Pcxe386fI5qGt2Udr56Dqe9pG+dWXP87soqU5U2
LmEnUHS8sKm5grrdLm03/px0A8S7ybMoq+Lebo4cLFtLPStMyT6CG7aNBYBV
7XqqtkcfKJa3wyEHBaL56n+THcUlcERiWwBfJN0cJes+2e3hlvPRCnueCQK9
/SwtDExsRp6HzytVNJxjXTW/jGHIDWn7qwvXX54+8jonXgaAXTQiFSdjamAj
J/OBH2YwGNViQDPUuqLUHsUP9VOLVZtt2zrhfWNKh9JWr71pXRO1OD6nUnF7
51/o5HsBjUsYSoHbZzbYUdiseMuGGHsaCKppTN6itYC0F09Lf8SIUUipsWp+
4jPRwbnn27BDnpKvxmuGMd3aj0uRcXHhjjIK8FwUdLH8DhMtINy9mOwZN3j1
uukH6ddQZXXyjTdhQ0v6+Z17kSizy/uMRG8VF+4kESu+K7SvRmWvnDPYbKQn
hACY4RwHQ6BLcYiFPu9aBqmBzBI1SkUodOFKS7/wM6dBkNlf9ui8qug4ncbV
JDheQ4FW45QjTgPIiP3e1ZIR9YwswRkQWEwBfteSW+Tu6gms9WdWgbaYXQIN
xftEBeP6Tm2tKydJBcZiCBos7l/EpJD/1dWZbwjR8jeokEblV0GUmLJ/dA+l
D5pMfjMj4JhHjpqD7LZ8FfdgjbhpxYR1he04h/y5+GiY4y52UsYwV0ROOFh+
c5I3ZOk9LELB95v7u/SFUYJ2Cn6T+SSZLV4TPuYiDM9oIBnjVY6u8f7VAfip
5ywvSbqIjEk2IUU7xZbvva/TRzNpY9MnCHOaPgb50U4VjaQGLjZX8va3axxk
2typcUMrnyujZdU3LFQxY7t7tIrWpzZcHwMvd4BgaKaF8GhtYg+bUDXvfbJ9
t8nIPM8CPYDzbrKfETTm3RQFRpnK/at+k9V9otOg5GqsSgMQP0xPGGwIXNVQ
I2zAXUJ1c3C2LHP53RMJrgWtJJzVkGL/iYomIqTMTySUV6cNhwF6hnYMTZdz
WoiIHQs3hBvJ5PmIo5fga8Ck8ilZZlLImw4ecWsxEJBS10bQEXuWPQroCz2j
mYe4SlCcfjLGXjL8xHF9WrK+8kAkZDth/EsAOOoHt0nquy1FoxWc7R0rHQs5
NN7++7/c8aMULkw2kqWbCZ6gETtoe0LM1KprbPC8fDfB95O+02Y9q3+aOGAt
UekVrGL8wA6QX8n2WCYRWBwOjhL1COEveQIAtj+6mvMSa/BrFNi1mf5WhZ//
m5G4uuEIEI3YGI67Gt7yG+5iZwft1Ifhh1S+xaLdXAJ6ybRHb9lDLe3sGGhb
jIkveJQUPl7Hi/YOeDUTEr/+CBUF3MMmDhrBc7JmoCYx90dmpjg5isXdjMo4
kbnl5flOXG156pl2PjtrcbEZ0iPbaVql6290+NhTQfvQt9rXFligRzTxa9L/
UEYN0ZOn5ls3giaB1Ibs2McR9ZLJgso2NVayI388duZy0ZI2UeXNJW3bzyYL
mtauct71bqG+8MBU/TdXp2/Z6aO/HiWAjRNBS+X+3vKotQdFuLwBFW6o5ZYg
w3MZ+8npfMszqacfL2S9OesOUo8TffmBC3cHrC7e/mQOSdnw4yW58T7addi9
qHnDq6Ba0Y2Q9rIyqdmoB7sixlnvw2BI2yHsNEqqlwDxBNY0gwkEKjVtX7t0
WJy/P+E4qfgz6SIX1kGaDdze97R6Ce0xN4FfBow+4IPSLA/jpgk64PwW3K5Y
S19CU/AtXRwmB07cXFPX13TXY6TfZJgxgrBV5ctYFL6A0mEwuCQUtD4vjDID
C7rqMN2NwhJmg1mSzoVOSxjNgy7g944V9/Ul5MreZQUUbjILOPHZBa6jroeo
th0+pwqh9HasI04ai3700cUWUIqEDDwE46Sgh2tGJa46UqOsqjPmLBB1qXmG
tztaxoxB3VVVqHc5gPKzHJy29dRHYjHr5ZZ4dEuCoc6fH8HyRHZmdFn4GMy2
aG3LW09Zf9tuBjxkiZ0tnsfah04IU1jKQBGXO87bvxt0a+EB9GEedu0k2MbH
njmhRNpmklEWiYoGOOUWRzALOh5Y+CBDsRXQN0kJ5K0jtCel//pH6M2CTvt9
CBpNddSKc5BhUs44mFLevfQxc6NIC9WZ9Tuqg4xLqr7qCZL8K/D04bpGYfWK
mYpBwOO9lIbCpt/KVUYlxL2uC+z3wleP35VT1FVVrs1S9fMVb2huyH+0AVpQ
UtCMr/xTxW4IJT9gv2ugHBOXkiA+D8nypZ/JiRWCDnAsOPoQcYIjDuVqEdga
YyZSyzomzr1I7D2pZPQcQ1VuVxPYjuWBZ60PHaYw2QFPkmKu1AiyP0ngYeC/
lBX7LQorsJeU9MbcCUY265shXOmMK/LceSi1VoWSPTHXga9agtIDmttCwOxT
fu/KdtShU3MAGLwgkdylk8IAU7VFMiDdAz85UQz5KRYXIFt9qugksOtM3LhS
3uCp2Rn1p0kkPUlSZ7/kdjacymtup5X+FxpYdVIq3AgZOCyM7O4BbhQUAl7z
5YF9q0tZdWejmtKH8PyAeSbbSKlduZW3rjelVXkxbHg+fdLZcqWJCuWKpfQH
7ntisldxVKN+3QfAWwGd6srywPBeaxRnkI4/IKj9CMY+cSgUFIKaL4COEMfv
GDZ6138MvhBnBBwT047owSaAKFn0nl22RMsSZiCT7JdeqcBVs2QKUD1L2rbX
0ISK1wdZdFxJb+k5NK1b4Fazxo+5MCK1Y8FOZjO1RQu232iGTQuJmv0XWef8
Gs8KtnczxUzCWrjmZb6nv3smXInKPTnhA17BU3jgFxZAGgXHcReCfKJjYT0q
GjoZspeB1PULRqdv+JTZY8vYam3D9AEDCEnRuYFiqYU21zx9UUtIonf+EnFE
Napv6q6SNlirxZuYBedFrvRWPnm4h9QlVbx4EL+oyRDSI9c9q2YkoIVEEm3L
lxqwOcR9KjLuIFxHzIgPTGdPyVFhHuPNsisiBDamPPjD2MbbLVX3OPkk7HFd
g2ByBTwEqpJ3Cz0SVqI4/30DTNzciiF9SxwwSy7nXXjc0pmhKwL2EuQ99In1
po6npkWELF2Z2zNhhE94CTBQcznxhzqyFgClhMt2aRjR6GiE8hOFeiWoMSOH
6cwgSe0zJLp/M1etd+Q4Kou3q7i5EBCzInTdadbWIja/ROW9cKu6GblNv19D
S0GgN2EUbq6e1Rt1SJR4gAoXN7g39Fpiq9EYd5dkUmJHaQj9i6xIIZ4dVfRP
fPdj48U1lmZBdlizx4jpJ7i9u5EUZC5BImeus5tfc558PG0qKtKcrtTU35iw
8XoOUqlM8sLXMtAgd/ZT9HnrzslrBCaayjQAkwIxKfYwQlwTj3YaXJM5PdJo
z6067lIFZyzeac0D+aj5uRKnKndV64Wr6xNulVJA5M8OiUcrA2ubjrOeEm70
PimwOkgJEFdqx05z1MNC8C4Q9DLHPwFjGay5IHmcroRh3dzlWOKsbGSaiL8T
eSC/MkZ8LvXk8nKlbSgK33r789lmlJIlUL7tNPAphyyhSNU8TqdELLhGKgn+
kbzc5y4UPdESmiv5bxqlfKoU3TMku1c/9D1086f0H0Z7vsOPbndgbNrZF6CI
JaMGXVsBEB/jTZVMQY871yrek5iNUKyiupmeTHKDdAslH5Qw/4joK76gcKqF
rGZdt2RLP0uMahtejm8hg3zc4YgcZMued2jfMwpvruLXqb6oQoiUC9i/anCQ
xUh+sk2i5ProR2W4Awox4B6JR4H74sRMZIgO757o+m6NnEhVK48raWdyJXm7
/Xq3UjfwhNkngmE04DSEle4FHlFh2lh8yzMtgkMIJvhnZgGgsrUKrNB6+gar
wKuCGKwRGqN81ihA1LPejKkonljzOtOJu4lfRih2dShn55OLyMiVxx5AClJo
b7x3kSSRAT6Q0la0T7sjPD8LWunL0zPhDLZsrBlqueF6DZ5HECOlIvcVXzZX
TG0rKahsP2U9TSSoNQRr/xgVOOSR5fIiea67dNGo/mNmdUcPdbx8Bv4VPXek
jF9K1roEC23U7T+HVRVkzFJXcOVVS5uDoNkPW1N3Ib7knixlLfaeb2VIQ1aQ
/TXln/Gv9GE7TO32obrjaQf7T1lcjVpkPfEY0o2jD5mLNHrS6rk5VLHr5PPC
5523Zy7nQFAQJrnzuaty1jftFckcfWHSjGLwsYeUsk3mzgNegrZAF6F/Urm1
ZMItWTueW4t5fCWZxc1LTa6JWw8q1rG2vOexalCyDtSgsYtIQ0nVazkFk8sD
Vlg2MrB6bw7Fu88a3iXbwSXsFwKT5C0BnG7QO9umVSE4aQu0yAru3snq7ba4
HQ1hN52xb4iiUBRDXS1X6xEYzOuLTtrBfI9Lms9qFWQPJdPi5jH0EzC/E0nG
iaqVqS2cby8EV3E8fpqosnMKgKpRs8SRRdhgtBiK9yJXwUPcAvw1s4H0SSpz
a8P/h97vP4Hlj14o95O6HKBPpmYPIF7XeoxiVqUB4S4r2S3Io7same9lslWe
aCcMob/yMU+JJOWB/Ugm8ym8dcLAnn1sOw2en5lpuaNTUcL86cYr1AsGC3WX
fIfuCvR4rdcrXzhBgRQmXUxYi5mW84Mn0al4zcgx1G2JZqwwv1lGXAIpjuNj
qkSH8tkgkigtZyUuwHUFCQaEwSW6qvU+eqNsyEYrdcTdQgXG9uH1yZZZeEWY
6wXstuYu9+swPk2nb/eyu5nMCIU9E2M7JE35ByF9XwXr5bx+NceaTEPvtp6y
Nt4JCVDHgZvZevtE+Lfmib5YpTchk9gjMh7KD+iPK5XhpF/YH8/ZfBDt3lN4
d3LjzfkemkpUMnjINVOoPwHB4EEeQ7xrg4QGlftUjIJ7S4ABe1QMCnQ8/KJP
BKo7IJwkTtjUBL+VZYYjYmHPH19x8uvxkX+f/ltR6q6Wi8lvDc+BcshNUkg9
Qv/mq5TqN0vzk4C3KvnTEwMKsmc7L2Ay11conMSK+FmZnGdjtqHPhaf+mrUk
2DE9v21ghSuTJfjD4ckW/aZb1674abftcbbwT+PFDr+oMFQt/i+Qm3ZJ8JIf
2YJiDCH0S7owSwcW26L2RvvBnHGPYZusLWlTZm2x04kgysBO+AZU57Lks3MY
57HqEcPQ19EwUCsUNlWqYkd0LCq5P6GDe0x1oAGluv19LBGjdXZ71muw0pCS
Rk1X24MgPmaHA2sMHr1rMY2HYuarHIvvXzUFHDzvuD0XCevCaWPwdLMne50y
BwOt1g9xQQi0ogAaCGgdKEmvg9CjmbeKypjrwqPZmmjiaK1cWup4aERCFO6y
joPR0iwomLg4v7rRMcFvzhCp+9dqiQPnkXTleB4H5ol/s1KewdMXPulNBpC0
KPm21fK5ueLc7rnCRp5at9WOK4LYvIh33aDl1HFdHQKG8U50W6wN/KCmzgu7
MLb7p5faT+3zBLuw7dg1oqnPY+I2wh5O8Jec9SchNnlD/Dmu3E2NwZ8evwnx
Gl+10Ojmw8Y9yaB/YJSmdFtPWvGmMVgIzbNlSEwohdcma/g6EQVjhmkpBOlI
QW153TEcKoaVVLg6gwyV/ZcxsR78ZuHdE0Vd1SQPB+8LE8QJxaTiPr3s+mdQ
QhDYSBp4sC1h0LOYNV8Xi66NH9PIAOc0O/7R9KU1GpV1nhZZa85kdq9X5/Az
vK+ujCjToo/t6mhxLNat9I6N8ewIiKvNl/T3I8ex0MtFq1DiauwaqjC64T14
Z9o2DDrVZN8bA3hHaGxdpR5rxBuQX/O1jykK4UEzanHY9vCusJg4T0LMFkZR
wXE9/MMx0kmR+sm9hj1HnqgPLazZvp7aC+AV7Hi3qSVbZmUjaXgWfR3fwFIv
ZRBbbq99RmNAQU8EprX3/lxbLmYyTymVHSa5b72HYWM9D0ULwmj7pnJn2KFM
K+OXGlmdZoehhlAUE6P0oeq7vC93piVhnmlyrM7LGcsX0BzKxif7bq3GfzJp
k17h2fiS4rPMOfSMb+TtOBT2qIiLpK967veOtGShD+sg9vlwIrcVH3jOARov
kICbaY2gwZ1d2YY6GFMbnhE3vnKM7MATGjUUhwUSY7Ba4SJUc6wbSXzi9WJC
G3s7Bb/3TRy7wqnPJsu4QArAkXuMZm1Jv6RwVu8tvg6LKBK1BJJOOlHaGk2U
oPNmvgN9wmNdHkZTuD75ZIWJrddtSlGsxaKROyYW9GdAHUx/nZ+OAgYoc1WG
RNLYqoMXpLaX9jeFtkDlgG8eX6i2NKXNCJXDSW8kwPcU2535hIbeDEDklVqc
OdEEhDXbjZZ0NbPSNTQ3iutc6mKvJDlpFl2JylXfdS8I5/dve9DHm/cMRp8p
RD5BvJ3X8ltfLDijv3bJVLw+sSdb8PyRyoYIg0ZEGw7SIcl0pcwwkm55Pl2+
fMKm+SYMYQwj+RG8h8I/V+11TYNBcyFUnLdbFRg2wsthEfM26Di3C6hM93EF
UzqZ6FUPrDX0qAbKZwf/pt4N2F/T2jl56R1bMNcTETw7KuGkaQOcERaEF+Ri
KH8TUXkoXWqq3jQM0ijQlUub8KVwfGd8RjkeJv+XljQTyrTWJQLwa2vk0tI4
AmV/7VtOJsNKYTBjy0p12k8KfLLcjnVcd/q6gLqiedCjozkf6CN4ZFxZ7h4l
elO0SG9Ng91vYBTNhszxlQ3tV7auuDt1OuES8vShuRXWBmtjdPHqk89bP7HI
ntZm8okVmJ3+2vQpXUuL5SGl+kldwpuA3nOQYywoHcEi6osCJc3fE8sh4Jf1
LKDwQjI09AbLexOm1t5bKvaPyrJKLeX+VooWgtVB/bJ/cSjQ/akUFyWmtHAU
32Kkcx+3nEV6+Jjk4b150cguNveSOhciK1UfB7hNbdPis0nn+liZuWD9yVtx
bSoVBAOgCdgR1yQ5HRNeg+9gbAUGhNB9opp/N/nygg7zwQ/taaRYLv0fPxGY
izi2dUGjGQEjBjUFMQ11LmCQWVctO+0d9f3hYrLSXZX90ZErvRxjxYEYoBkJ
gO4Hgac+mImgJetJ2hmwAGeSp/ovEQWyVZot/94i9jSgOGRnUJXb/W+Ugmo0
AM1wQgqhWPBLIC76gC30/tWpOl08uGu6tcB672m74ejZ1JQNCP/bWgHain98
aGICwACCJGionbVuReL2hXr/24RjeRaIw9o3j4DNlRmKc45RoiKAdz9CeVlX
T07BZWO86nE9mx0Idso8mlS0XgLixKZV3vtCIlcevPwF7A4OIrS2tdcnMRNd
1Bq/kgsbWYZcR0U4/04lJVuCsUYGAJ9t41BSKtw09yu3iIOjt+C2reccAUzj
JPPHS0fTdspCbddVDHM2gLEwXQ//pTMx3SmqNGuwgdfR9f8F8naRmOoX8EMo
t6gUeMfC7bVUKwyEDFVnVB1XHpTosAUqqDj2PYIXDeTHe1S7UhlWeQKXe8GQ
yF8f0e1gL1/nCOZMBw/65V2NPAW2JJF46TWoOk3i9rPnJ/cwJ6e+e4v13ibJ
6wCm68cEnQ1fUS/1kq1CItQklJyQyo77iQud9qQbItbHo/eeiGwI4x2mXL7e
PYS/OG4swH5LFznFceYL/JbfL81Q8WzKNWmvGqHAx3Tk6qoUKwItmdFK60sm
ua88zFB8xesBHI4zZYZ9sJf+g98YRrl0vahEErPWWkdn486D7zx39XWoWEvs
XeNfwFQ+Eo2Z5XLq/cn+OA+IqJdaDS5wU7fQYto3rF8OhJPvjLigzd2Vs9xj
S/07YA2iknNgskNVo0oXSD6/9jsIAkxi6nhqtG+TwQLoskBkL9Jn88p+hdqm
Mmu/BdUt2R1Byc8jFyzDPU6RHYrsY8ze1ECC08+xselobkeFaqncGPf6VGRr
ST9ODW5cuG3oq4KqtJF5SCRPaD3QUH+N3WnVLp2Pnn/gRGFMFfjX8bNvXr7z
iwS0r9TCcqqJdfuQqS0RiQkCXNhVjSMTdqUOaAlcqcjoPw7vgzp+/2catpnw
sROjBeF7FxqhMmCC7BQxrBdkUrAv8pNQ93fQcilDY4n2c+9ECPe+y/kQwYfA
0aeTkp5xuiUad9XLiCRAXMfnt3IroOCcFttHKSVsniEym1yjyFpYutbvyXpM
wwAOrHQiI3X1XjOBZEB6jnu4FgrfAofBMEEaGhraR5PhGYN176z5QHQkwn6r
FhAohNh8tkzJbCJwYi5I6FPu2c4GdXogBjXxcbaM9pbaORtkEg4RArYtEu8Y
emr16k7qoqvDuq4leEbBoM+SthckzBrpMHw3ue+E4RhDtO8lY2VkJs+UVy+V
0mlNqJoFLYhykv6WaiWgNI+J+UydJ6y2rVoeSzUdhr/8rE72jHsEoREmDjxJ
twbs40OXQ+fXi+LBgHIwyOti24lt7vhkOOIEKuzMgEaWxf3rCY/8lwCLtnbG
DQn3x3iwClKZCuxcwqm1ZSoVI7uuxsf3asrdm74Ss9FzST7aY1x+6jhe94n/
ctPJprta0GMZV+CNmX2Ql18wq75ulkK4VvniZrlrAU2B15Jya2h2YVMI/cGM
vc+btbmIH31YrtiaHRX+N1BWSWn7WEG2yp0aE5K8Rqdurv+ljnqP28sxCE/g
rysfm7ydBVvL5qPZjWyNXgv84b5jL7DgaW4s09e4iJ8yQ7XWOLuZTlU7aUWZ
tN2VQMt3ka7/+C2hvUlgHLkpnJ9BZj4uZX3vI9h0Xn26UK78tVbjXhxiT2gN
L0M26E+ERPOwU6ekg6K2649w4OUw4gnbVFqk5NBkTatjLrC4ggv3Uvs6I380
IcgInHkphJbHAKaTISfH/J9h4f+6P/DjczpZKaHUrKCiTQrxl1j4FYmclS+9
UUZP/KCnplDYP5t6GnFm9nGxh8o+orwlNq57AKTMj43An6wQIsF2HpgCGdAz
T5YmV0XxZ8aiO4V+OHwGhEMFb3as+azQ5MjGNgqpmLYjj9VI87VGTGUphDPy
iRy6cbC92+f2vtwl2u3+iZSpjDTUoRH/hUcXjAKdSfNcIvOcB+Qr8KsKxU7X
InFP/PKaLH9eDa8B6MSh57qAiI+MzEdSmowxiSSp18EcIqvQeEXFXU0tbq7s
pqHATd/5opo6reTazhihph1MbPYsZ3HFbWwM36bQjN7LPI+3uTJ6V7CgDD7I
Svv5Zr5O74xjm2XmqpGvOeS0vPc2oQSGo0X0A5ILYCDIvckzOVSqRE+MZied
7oK8lh39Qya44WV8ywDMUb0q2W7ammN5OGyXf0FTfmMNb55vdGX9JztOZy0V
x2LWyIQcytrE1sGB/Ad2PW3ASAqrrokH1+30tIa0DRQE2AiEvmnrGD160KXx
Ex0fVBy8149fUN3/Pxi1b77TKBAh5NSlvEuQpXPf7TIBvnVDrplLjdXuGPnU
C9Vg1f7uBeaegP1YMzQ3yrWAthoiurqwrVFQF3J/UEWty3FRXqd7GfRy32fa
y08VMkuZUqqdUmS/YuC6/eVoNhwpMeXygrqLJpf1Ec0yxShBxxiKPXENbsjB
1WffJExr4dyiJ1lzMRTQIOcbBjtGEJid7oQ2jpZ5YROxmzw8w0WiWAaOhR1x
eGwLpxeVHu6yNK46Qs2AKWLAtyqaVLtjod4l5ZhAu2WsQ9ITqKzKFRI/hlYT
V2ucvkItadtcpCPDGhxsrLdQ0NfFL5ii9cVEZ4RaqxZpk4Qy+TLl/0AaUTGf
pHn2T/e9UcS0ylxDsi9YIU3IqfTQKTW0x5/ig5ETz7A9zTgeLYbdfanQv/fV
5d/DGfnoNeqw8llKfWXweEU9v7G4gYqdTCWuQt4yy7FfEgFGCKKO2UkyjUTt
4DdGMGNinZKQOPi2/C6MKpN7D7BrHummlW0IzO06WFPIWyg0eEmGC75V+uMu
AatmRAeGxm8aO2WTl8CCfC7pqjsrWYs6q4lOQa3gdikr0oPAxV8ic1Pu1Vu2
g0MsvbWTzJENYpYztn5BQYaQ9DXEpfTjLDVa4eyBG+jQKP9WQ6YtCM9lZzVm
0gNXUodtvwR6YUpyqct1ut3lP5pcLWTpht9bqlSkDzxdR46rz9WKRVfPajjO
naQD/xav6J7eDUFTiTJ/Lu7v463QGz40+W4+aQ2gRbAA59DDX/48Lw+vKs9T
qiEGkocBKa6ZEA8RgoReGh+ebN1QrclU1zg0dr6EI48gbh8NriTDwXWpRNJ3
lsltnHNwls4qj/P16APHmGuqVVAALWRRKLUiPZ5K6oo+fAQm8NUV7ybDMYI+
ereINcuOe1Em56XB/yaQul9Mt2MvsdEKUE6+JU2BGxhXdkdrwK3JHgLCt6z+
2UcNg/t71MaQgZmdheU5VTgZnRozSMDzhhuvVxoaAihLMxBb13JUyBS3RUw3
OmuAVHS76Toz9bqAtqK+Adn/4z2X2dcpoRWZD/hrtOAIPAYj4iZBRy6vwM1V
kZLWNiTFgb+Xea3z4l3rUpN9e2XcvP/eHV3DSXHLY1aIVJAkkfu75knVRp5r
8bIWmXqw1Wa7WTAsJ6w/Xbx7gxI8yXbWdYmo60Dm58J/CqoxHgBY/yfhwNJ7
Qtx4VRjW+zzrpJQnRH97YXz/AKJLgL5+HLawa24WbqDsvm8wOTsgPTzKEhPL
/FTZ8xLh7btYfjd8a2yiKd0fpyx9DhK6ezukc14SkMNZiEzhbxSM4MgjbBhV
hvadnJSk9nmXt/7Bs3eHvXE/kxTnNxWiiuIHmIMK6mDgLlqChH1oL8iu1rmC
qdrtO14+d1J7pCH0Dgiss0rik5blIrA/2g4NA9mIZ6ZFK+cUQOVIxog8wuHz
m4YEMD9tJAbhvXJJBPkhw2O1434qRtQHyZs9fEDR5Qi3jNLlnES49a5xijMN
mqMtziOpzuvf5bfwxhnn3Sic/bfenYFdmMnraOiuD/MPZgnstztrxQo7zsn9
a5+DxWNpz0v5eWoo2+p3wuJQ1K32NedLOInd3aRsyo59e8wAbl0EQjJa+D6v
jOPg7hJ/KtpsKgH5HkqjOkjrFNP2p1r+AJW+gAfgMenxX1Z3AoRGC04JHJYS
oWxg/nMpx1HLW6bHKO46XZzPTxOoylOIwB/AsXS4PWHaIWSN3KANnnU9Y5J3
lUDjgPMyRFGvem+nJi5Snv4exwWdNAl+fcGhPYKbcXJPESjqC+9O5aEXzzeI
Mts11e9AgDXIAnNAjlhsjsoyGB+TpP170cw/p2WwTlXbOAoKi8I5jDjtqlZ5
wuhTlqcXZjekyxrCnWO4G95TS3XOifyvrOUOS5uuv7h5PdqR25ABw+J1yFn7
+MRyaAwLwcNQ+tRrPea46Zs33z87XpKelnkFiFvy16aMh8i14+2+7LvVqQzc
YI6Z87NZKB3xYs+qbe6XWe8L5NWXIob/7P8Et2hMhPXu8USVXFbOeUld5HEI
JKHq1gWpWYrh4ttlNViEkdcIInyjfEQTLPkbACJzCaArDy4bD724OW+Oh3r0
yEWS3L2wp8061XZ83JIcUBcuCaFBjq3UQ0iuVC90CBJmu9diMydJCTDELvCp
x53z0iISdSIkO3gcWJWs5Jfdih154YbR4J1iwjRhb20JvTmOqcSpUrMmzZR3
lozSuwFBKC2jg+ayHY11+4VMhzy48hIx1/z8qgYxZuX2RRy/qyQ8ELtNrX/Y
tyiOdhfABHF7B79CpXmDUrp4dS4FtbzXlMRJQa1lrSbAJ+zJbQmSbsVAGn8f
QWC7Kydklsj2WJcaXX8yXZRojneaZ0Z8QPuRYhdoGtZ7khtMWh0Ew+EFxILX
lvlaAaTPq5dIiSt65mANfbVAzecAs6/BKPwZUsi2JbvPcqQxMa5uVa/G28/t
vqfYND17UOa5GeTm4V7SLKjJKoV1+gLKtUnidqynBr5w8LwSRNK3V/REOAb3
mlPQOw6HYU6qlbdYq6XWB+0raN4erJ/LMNZLgc/7ElTL53Ncl5+BB6Dt2ia7
eJgSyr+/xCWeT0nLh2aeIUcnF6wcJYb8iRqe8mjlo5VutglWTVZ/uDuzFAp6
yRpLrZtd+5Gfr+Gr/jYY5MQXAOiQ+dbLCNlA3f8bmnOsDWF6MuFqh4QNbbY6
E0qPOjqQhgSJySz9XQSyWBT65pNUBOT+nYZ9JpDhsCm1A/nTvWy+/GtoNJnx
nGu03jgJwS42j625EZkzij/P9Nw45oYYyxTxahOtHmifKCy6ZyS13G5E9WJe
YqNpaUeAmlHi0/zF+o6b8vmGP+/8FTsKhHe7iah6q8EMSp4CxU/T0npsPPp8
6OlAeZPJBZc2PQHYHF5HrWw5N7gLHFzWVk8OPjAMddmGd3Z7191D0fqRIXlG
DXZxMo34Kohk7vtZsvMQv1NfTSdaAMNKXoCx0DLBsIBDbu0oylvcxSoVIILe
5uygdemCaBdLY+YxQmxNjvHfYGXM2OqJheFAa0E60lDwEl1TvNVafo4DhFte
ea24qii9qZFavbTZL/RZEm9jlls8ZZlfB0KHATxoHcUc81jvDcclTd8LaGlL
igXNNO2re1WNQi/f7E9IbeaSwD9ivYqmMmTTlp2jA8YgWwf5gwao8Jes8N55
G7viZ8r/Dy0tWfxISM+gS0vP0dsdJ5hDhlO28MIlzlZKg7ArMb7GTjE/45c0
x6Ifxpjmh7ZeFa8jaaUqKYwHtwxSFnVwm8ifouo0/Pty4Nt9FK05dUG8mZ4J
kvfQapeXF91gvZ3MnJ9Ys3m/Zb0QGcko1Tx7MEPMslsiU+g8g19ljTS4dPvM
55RbFGdXCB2yCCAUomjIyqL12sNMiVy6NwWu+r+w6Z+TkVanUpk+waGXmyIm
w+h8unQvADoL0vvwUFOJl7b1bQNO2UIrvvfG9Jg5y/DG4dfVxSDePvy+aQPs
KKgNFg+n+149c1xCPz0m/CNPqy/PS/AsYYOM+yetjAgWIMAtfiibrkcNrCdY
uxDSqMAxof9eh6fgzKlXqWPQyue5PuzL4fceh84VtzA5aKjIXB20ExVP0JOD
KRTA/9//996Fn7g5zAFKMAIY/wSLe7FqE4IDWlKk+jzppkuT+D+Ypj7GEpye
77xlfQYYMT0c+reG5LkgrJfCRLGF9kGo3SEHzEm/OfzlhmDLmNE2TxQ2V7E5
kkSttCdI7jnkX+Cd3sxSuwXLR6YGx6qaKh0rdmtXQs1vK9CAlRKUsDkLhKuc
obe0/jtFQRE3Rv7sL91GsE4JSngFLq+UnVG0kH06bllRFgRVFN7h/lcucwMz
J7KLnRoXULW45/bhJHGL0x+qjOjQBFf5P/EnrWKHbrcnCxc9N1qd8X21kxV4
zHxKspMYK6Kh41LslIciUN9keiBmKCHuZp0ItOUNgE9heuzbmw824gztUJpP
hLewbPJ4BfQ+8rn8wZtcVK941aEWl1gZrD6KfZEVl8PkIYcQJ75W5ZoBDyHC
XEvOd5UZocWFXjZ4ucZYph9SH7r1qYKpqcrABveM94/E04mZIk4gbRBk89Zj
JYoUzxkMNZUVSpEf0WyYXefsFai4DriVECXtzRgD+c5+nCZXC7cyU10raQy8
bqq2BYMas0xuVYLdnAiSn022grEmjLkGJZJqaDNXwUiV8haj03u5a164lLPY
4JF/mMLQnq9PZLVmOCyGOrASu6VKDqCjtBu2v9PWBxiCrflaGa2ij1RvDlrz
KFrtDLKQ0qc+LkYac46OCf8VWk45xKCFVPt2Bdf426XWFUlp0JvPNSkU0u7f
uR8IG/cDHnq6BL3ba5RInOmt2eJ/RHEOCRiuSqdwyEssFAooGHhzz3KrVD44
k3+i76koOWGTcfkGAU9eR3K1/Tf4x2eI+l63VSSntyK1KWDufulJlClWt4ds
LEIX+GDISuSTcr8r+oY+v7P3FYLsx1UxnBmytkc2LZXf05Slb8iNdBmSmjep
fwxpY496sXtP+w8L7LnORxTXfy6vJDFXUgMwGO5fr6JY9o/NMpUampEG1/VJ
JQwryqwHDBSVMtEXaAEvA6vHBeeR0tnmY5T9sJ+nlAmKVR63k3IvwWQ6+Kap
0aHC5966GwP2BC6pe9bC7yaqMLgcXKex7WamSGzeOImL7bANbpuUjcINqljC
/Yw+28xwpK6bwydfsf6L3CbAKsH3DfkAFrrr2gM8eWM8ivhqLVXzzv3gIMoW
NIS4TzR9zwh0ZwbHz/jC9nliQll5tpfKgqeLVQu4nl+w2Blu7JJd2jAyFAmM
xeU8+a6uK0mGKHUDZPMzOW/znOwUdSdqrW5FIbTKFDn10+Nzed84bU9/cp3C
+90tPNtVyTAAQ4HINf4THHWgKumpQUwo6VVNXNv16MBf3x+tMWF7eTD5SECq
DtM4sg/hvmPBUl7tz7ZxTN3vbAv/KWhEKRpkryGRXc8xNCxdvZhop6294e9l
nnYMYr4e9R41V33lqZdnUiltNT/J+ZvfGop0sN4Nz28r713x+qbY6HcgP2Gr
D3Zt7N8CZMmTTDIwpw01FWezCiNeD63IyK8hBRyFfkvDkVoI2W0E3VsPJI0m
U2G82vzSFsuvej3lNaEuD4n0l5Cid3ET20oFRvmdUyHbHe3RDQBpydva4nxs
wRy4Bi5tHvX4Ux+Lr4/oH3JA62Vz8QFvZSi0vl7PjDMbjSqBw97CepJAHduR
d6GcT4Kdq9n/vJG7ITr8Q28YaujY1p767hdn0MJAMoVehCJi2hZYg53z7gFi
27tSFErZK5yUANwQR/GVYf83hnGdn+R3Qk7a6x1IZgImXJYn1t+De/BAF7W2
yNimlYnCVtMIRuCM2IbRpr7XWQBhwcSiuZ+5u1k9FK9R1TQquD5fhzzORd1v
l/puljUUJej4Uhm1M1d4/aAjvUdZoWtmm9IcfMGBjTdCMdpmWRy3AU47Y6Dc
sO4RDP7hGyXb+r72pHPmki47eoSsWYGdKVJ6qeTrM9dlSVGm7A73Gbv1UiB6
759UCKppwGSvxgiJioqtqTP9ajwJaCrhznjpsw0uI4N8JSG3tbT86TYoUkuX
24AhspB048KMEaq4zaA0pskWI/5NXqCVUZ0qcTrKvTaM5LYrGs1NLT23Qc3P
fL6Ls6SSz6BlxRn2x7gRZVyFHUdrPmNPa+1i18XZ4/pFBpTN7v9gloKiZBVx
lmJix7g4K6BU+q1B4vfLbV8GGwaFgBYpHK2i0MGVNM2fkISvwlSrX63iN2Td
iWq+v4Tyj9G+2JkbYB0SewBKBxaV4te+WpogpvbdiCif84p152BlMCQ+1Rp5
MF9vbpBJ3nkr4jB+EW9YR2wQ3cpAp8bCo0f7F7EDZR35ZxaNbXCS0Y9Jx5/N
OuNg3f+BzKQZ3XUXT0bWkdHN/zLUxtyyR35QckOlS4fraB3m/01SmsLfjCu7
qb9ZMylaRQEq20d+noa74HmYcm6FW+efj0WwT2uPzrJ/o826oUOm62sxyo1F
7XuWQCuNg9rEdxJmbgxjbIEVFgGEAFQbNgG1xdstyjkG4HQPC12SlHxVFhGj
nN/UcLRJMFzSTzRYmB/teqT2h04ZuHA+pyE7QkkBx6Y1gQJp3JfPIAQnMVHQ
DaCOAeLYc/ykUrtlpFlx3CbwHTQ14/JIBiLN8gNeBk6beAoeDow9DhIzIj0L
tD7MF7IMD/lvpFY9Jt3Bmjsc2KeOYGK67ufn7dShvEDnlIy2YjNARminc306
W/5E66WxMi1TZhb+HGO3vQ4BdroI57Zcljlpa4s41VetSPE3enlnZC7QCySf
12XFRlmPw2fWqoys+/XVYsHnnyXTKlZ4iX+I+HlxxT+GaIdFJ5jCuzY2uoMl
YJE1V7FVeiFWBVG++WF6A9nfBlsWZO1yFjSPvQ9ukuv5PygapPeMe9+5RV3i
9L21C+J5F3bM0rW8WT8BqZl90pN8ktrXmaxJxmJP2RHW9bkP9MLNBihDY8Z6
iwdiJ/MhOUdjHXz3AgLsBKGgcmigmBt+5yf8diLbVceFE+Lg+MIX7XJfzHgu
KKj66K7fvlgRHeiLGx5THjLsL+HEp0RCW9IjROBsnX8Gq4m/iSTNsAgDWhiO
RCgg3cM22XmgVDKpjdYmc1ZYeOiAhyXKzkdazgLfh1P0CgK+VOXUgbrQkv74
xYM8Bs4e/mNu8nHzipBHXyonmKXpUC30cxC7c8TznpwrXerFCMgyfeiXqqbP
Rr0oVjxfphSsUhKrIK7mWniFoN1PaZPT5Ezepe50nR0Jh7jAPtDMw1QeYdls
F/mgs9av1zqcxy37EXKfOs56/ljQKSskiFYmfLaAFSTgwpQD3viZ1oduY4pO
4aX3HrLELgmxxQHrg++mUEi7Yt4d/LNdEWG/ipT5utYpE9vMs//QSxnagQFg
BYh0eq1qIiuMH/19IirgjbeTDwOisCLK8Ifj2AcRyRVfg69q2eVX2/i7v8qO
segbc0zt6RLF1KGSEwtTXd4Y/6u6HNsM/iHElPuYENSyPItGcCRU8CGR3/FK
n0qC89jubs18TMa+x1o88rZ/L3xCIPNNmb2NpgByA3H5ayOOwWvmTLDK8tDv
REyNeXvWx0kfSGLwlWSdX4pvI0g/OIZYSrzQ8XI5AK+DAbBOHbMFKnBACVXM
SZ95ykcsB/+eu9aoIeQsaPTCjwbo2dhA2D23bSCn0XA9IIY13np0NZSzcxmp
LVutiXA9alFVNBXmVcV0nxyxYLNV2x1oIYfMLJSTXNQDQi0LGODQyLauJv3R
KBCPpZoeUAn4fd+fBzv7Aj1rHmo7xdOp+g1tPBBg1SQ5CGMpWX5nq66UXu7V
O6V+YJtFe/HTIo7jZ31FaCA6idRaQeaTC/P4yldQnPSCCsGEUddGw2ZB5na3
MokaXs2TK6+BHGJP/dJQ56NrCKojwJRZQxQNSx97/89q41zNcCEZvFHLiapy
aFWv1IjpQw5flF/Pp6giwr5++9lkh4M3ojupkn+8x6/Zyjdd/YMcXJaXmgK7
AmkOL91hQWom6JY2XSjdynUsu+tFAQMwwau0ubr1jDPCkt7psOOLpNCMtGHd
QGGCDl9JDavZkFeBQVm6Tn3Ljd8yxS0YA3FwR2Ay8cpcVB9tVdbIgBZ9B0ge
JpA9BALNWPFWdiBZmudWCOKhnvF4De1ZMJJoiAi0iNNCIhmB9VBvaFy2JvaE
5P0dQq0kEvLPh98NE/kBYl7Ixla2jSFmS+5tz6KyFNpIU1YWbhLUlJe7HANQ
Bs+QvckTmuouNPd9rnjc9AXex7MRlcgdgcdPfdz7tqd/fIvaH7BlZct3dK5p
WU0J9bOoSZtSrEfJ9zn+IePP3gnVl2XEZ6l44NKLKYVBxJ62vkYysBHLRTGk
lhhodmQG00ffyK3L0rVQrIt94fWXUBkynYUMtEa7lk61whn8xppp3HbCOMVl
FPir047qjYZISaxxz62Kke2olckAe4qgEVtIEV4v926l+oyd5CUp7P1YBJjh
/zNJ5Wg1UbjqEKIf3/q5dmBVk+6vAFVUlo4hP9pGWOCBBJRNbNbt7EsmlHAE
EFHuvGxEPEyhl8NijTMRp0qtNMhQEWmGg7DLYEYAKJRH0tO7UAsDSqPiqGw+
Fk0QI9bfEzh3bnl5iyixy5pQ6Ow+nXBV/z4+BsWhpqZpRj6vwLRRwnZmq+5r
HuVfPErh1Kk+ekOBe168RSZgPm/mYDdLG/loe4asZR6GkvhFf99/uzHga6VU
HMIv7BsXI8QcOBMTWpG4HPqPKWz/XCYY3bBhOcfzGDCxbmnGYY8Tx+0OZjQl
C95yNntW3ibhXw/ptnnyRkI3611NV2zb9SOsxv9UgeyCGov5R7xD2e2lRtp9
Y3YDzEbruJ9Geh4DRmw1ZbWxnrbVos2TheY7GIM4WsL7wAEvDXrqFgO9imnQ
E0JTSL8nuayT4iSCkAimqsKbHlXziPP7Xqv4IvxHrVLzuL3IUPyRXjCTMs7b
NVDA8xURdh0UwDY+Anqk8MrZWMO4Xk4Wo7CM9dQSjucKw8jMmsU9ZdJy5rac
uEObM48FUaVGmFsI9pCR47jKZ7vXgv9WKryJk/KuDc+qOHKZG0slPrK0gZqs
qQ9hs1uytj3+WUpgn+mm+VjXhKCuUQ3Xbs/z2iS+rQ1R4mWIUVMKlAusl66I
R+WSUrninhPiRIaDzENnv5Z422j4wHfQTcDuFwrXo4YkgdwB/tic2Yo9XBBt
vOHeGplnO46q0GqEXEDT75uvxPhtljFQuQbuz61pHeN9jiGWxJ6cMLTUwGgL
kU8yc3P99AbDvUgkQpa34pstLlWsX8N3Rtf9P4XfJLOUPp004vvovC/JHvDg
uH5LvHYt2vczxchQ/xd/3oaMZcurUncqUdarFrqnTj2LDUinBB0lv7Vphadt
JzXLOTp5+8br8BhGWe0Mg/pIFgTcasGT1A43XvS2iz+pvuepcrjf5VuSudMF
8eWqhwxF1Z6UVi+LLtIDKZ2kY29wSjB0ECAHf2weQRnWFE00m/ZIxTehEO/H
zRUw93lYVYiaORON/f5A+cYg90WCem5ShRPFvaxV/aGYQGTeedFQJ/K0TaNO
r/tbxcsQRlruoqRNsoWO4M7P+PK1lfohHtEJGfTu3zBJxRmB9XxQ+Dq94Fpb
Y37PXTISRcuu6vhrzs+3tt6THQiC/OwSKLxs2iA22WByAOBAj/0/WPxe+dcm
SZHuQth/7x9a80iVsiQtIORoEdSKI5rPP6285gQrv6vJ/dR162vMDC4DS2JS
kFhJVE4lLklESJwzwUo/fVxHlTWESltObz7y7y9DMDnJr2fwfR/CPikf6zuu
gsS0GpCMPObac0ja6iE6XaBQ1zAB+rdb61bGMtj80ZeGKa1VuxlLtu0fwClm
uqdj/PxD/KBO+Fjki7wptRxZizoHOEDuPjXEEXzfryyotilAS758WZRTESlF
ySy0dOjXz4Gb4CYcGo8Z/Cmg1C2wWwR0A3TeU9hIpZju1qhdnU3YVuIMBUfF
lcHbuTjn+xOy+ZN+F2TslEsQQAtEiP9CFQsb7JtW4KoRR8bBhLfMdE5h3lwF
NxnUC5NdS/sd0Xn7wkS+PEfesUYKY7PeVbUm1nmQfcAi1PLTfaezTXrW2OUq
4Cj4Kq0nY2H5cmAxBbIvWobNl3TnOX37D1sPqf34mD0tqvxf306rLJ3Sa5pg
FXSaKgjicUOUKxGCC5b3QRRk0lg5dBj6kZsQAHBO1Dw2SH3DrR3ruOn90Y/q
8Y4QjWQDzhLkAelN2jd2rGbTjIWTxwSObm40LF6hq3ooIIbM7G9aUOZr6cyM
3qwtfl52DpCOs4uAlNOHLY6hyqIc/goz6aa4C4HqdD1AnCTA5pgFnnK/cGS6
5rLpc/nu0WmR7eiAJzTJHlMK3+0x63uZmFE0kIVe1+Fz4iQ6SKF0myZULgpa
UBRlh0G3Bdqo1MmNnYyg0YeLkgDgLK6NjuM0osh6SwEl7+f91jwKFxrjDoSe
bTvKV8Lkuo1p+ztuvJLK9lHBXCQHe1ZQ4hujAeRkASLj2ITkOn1eGTAnEOy2
SUzc/95gsFavRB8Z+oAFFfdp59oR9axEAHc7mLqzP2DnFHbfFCMdhUMe8mX8
edtVppAwnMP4l9kY26sMqxOMRmFQqVeo4shSqlnozBTMv5SRK5qF+ggnGYhD
IWDt3oBzTY/KOudEXjuchL4WFDoEJg0VQtKMRHkG5HwTYb3yv2J+lVJ8gq0U
ILY7YAZqV2S8ONweh1u8YQB7RPmYEN2c6AdogjR48dNJMFskOinCuoF0mE7s
We4Hjh8UU81N8jINgWFQi8IjZ6MlcNY2GLrefTYiOQv1GfoxbaW5c+8iVKtv
ggSqWDT1iP8eEVmBz22I2qh+awmDsjX/eFx+GbJI6RM2Xwqq1QKh40jS3y/r
NaoXnJi99yS5srbunzGJvDlJPs1JitNBUNPftHm5T3gqDy2i73DqlRhQwDtR
FgLq++Qj4fau9/tXTbL6p7nf9zHjsb9QDeW9mWVXjB9W7hUvDs3eSbjum+ps
Yd4isownvbAuxZoKDzffPYpTrOk3B+gm51+aQNVsxBvXc8xHyMouyCxSGAon
3CJiT5JbN0MEfrCX0y5oz5eMjPSbviO/4KAysFb5QfjxiycC9Ohofm5zv3dU
gL5uPBs/s/knfibb26ILzQKc5Ah7ujS7aDWme9TzT40+4TNnhfFcQO0i7fRc
4L3yzW5+UpYRWzwImwEGR7xNY18k0ARACPPsmLxngHnjOMf/PCbPAb+d+UZE
Pqnvau8OFZqpXd3K9pnTjgwS9l/RpuRy1bYKqqjwR0kONaLf8Sh7rG5HlQIE
LkbVy552RtIAvFBSyhVNyR0J9eSFfLwKNQe0HwnE2a1F1j8+Lf3Ny2di7/LS
O+N4oIAjp1RKEHuTATj+hsmVZkLV2ntY4Dxs7qBd0IGcmKSQFNxUxf33Lsg2
URPLeftSGWKk9a7Pjs4Fw1hbVuO/WWnOT1BmenMA4B8pgoAza/VbfZM7/BT1
wYgGuxn0Ni8WZB9lijBwCBia/84Qvb9JOi0/z2GnJPWbPF3KndI6T0iSzF5z
6uhb8py2bzSmTgK8O0/Xe+tYFfp0fXv2djaVnb3c8l6PxFn071oIvlttey47
Vt4HJa63zrT0kAMCO3wnbasqfWs4vILtO1Vr7oZpI57VwYNXqODU+XuxPXZX
yLiQuxW3H4nSNgEQ85wANTjk+sDztTbxlv6t+pZ4otw1PrCXFsUqeWe/YfRC
9jq3hIi4Uzim+GEKCHB/DwPKvRmjPn9HecH4tNgit3EnnpeR6BYdAoSGl7kA
4v6uv9TDv70t4ID4gR5L8qlcg62aHRMmloTRhkIOYm0HLts5UFuYTOJDmyz1
ATB0ABmYRR6b/LSPl7dL470KsgG71QDrD08qZ+0YOFd4e5BQPQQdzlbzwtUj
8r+cAPOZ3JVkWyme/BN4k5mC8tnuFQU+Lo8B00O4x14djnxpYt9m/V6yd9LR
KUVN6bqUfj17LnqATZHJsjfKbvuA1iOWvf0ZPp126lK1vjXKL64uSLt7nsGn
BDvui6xSYnS3XNYhuI0cQPKtJNE1O4aGlwHp5fuKMzQiXhaKac14oGBB3Ayt
1u1urUznFKv5eQoslosxebWTWfs9OsownSHexm51bPFlGRapj3FfThDd9aBR
UMKifGoJxCb+Z+K/pFUA8MHC6uoL8boPnbqZL8RArO0eGUnRcV79oEKqV2RB
a8iGO4SBw5whgANV5pxMtD0YDoorbqeZ/+6PBfG8Th3knkLnSy+fUkWBYn/e
XsJ/L67CkT4BSwLs8Yqfl1l7Adn3mhuhRpSfWCLfGlQ4YFJvxfVhxsd/43ic
Aoh0ipyrVTgyUruTHKR3BBW+nMOh/p0I8n1maWK6FHaa9cEBCWctIM5ogjq/
xCRyU1P/Qn2Kx0XhsZSleNcP+G9ibRgOgKSgXsbfuKtfkyqsautXrP++5o/u
HU/6/VL6SR8qQz7wAmzDqmobwYN4hh1jWSDNIL3thY2hg4AGwdZBEAhkyvlK
DjdpeY7+YmnuMUpntjniL+Rrtp9a/prGybmVqFslimbLXbcmk3F5RcvaMdf0
9IWpPNg+7WjzEFni0jYlOuyYUGRSsasmyPvrM7SZxEL/3uBMXNA0Wi6hS5eB
RTaCJekoANoU7Lppv5E+m2Yt7792lypOOCmFBl56tuBahN63QIrWhcr1lcmG
SoQF3xKBHuDCBkbpKUAgq96DnKwnBmuBPmayHLALBeRyrpznQBM/QwCqipsT
b48ukJVL9YMRE9omU/AinuBf3fUtHYsKO478+WnOeIOnh5whRB12++k2s6Kt
12GAm2pYXwZjxNoxYMKZjMEMwB0lUp8iniW+rHf3jdqLM+EewUBXwx+ROtGr
9LLL1BVCtV887LVJ9kYqxH8iThGyneKFIPE4fE6b76qB7UivWjBzuhaAiOw9
6jE05KXMBC9UMa1tVgBGFPanGBjEyUrJtObobWQx0mZ6vxGlK6i02JUzqpPB
ab8nlbe1dm8gG6/pFjaWqwt/XI7FFV2S5ew3TH0voJ282tOwcXRuzF3w9arg
ODJfyKGpK7rfladczYcg1Grkkbz24zaLAbeX68aCsDJPsBb2NysHrkuPXcPe
DiuRbxUJU41Fz98s5pNGBb3Q8ygLsgQ/mgrWgdazoyn50lfY8sA/mwoHCJ6D
OI6cdPRvvXWEwt//9eDBB/waS9y8Ai1wwMiWFGqiKF7fPZMtWzHtDHECPG7j
q3sdZ2yFVMAr+u5GXvqbe6zDDli8JGunOoUtWCrS7eAthBcVgXGUohqU76HQ
0gcJ+k6LTI42wq/6HYosGZrSnKoEamTe9o6mop481Xo1CWETEUnrGJRx+UC6
tKWneT7ndCQhqXSj2MKiWaEt+jdFaeTtndPU7kzhugBP+L3YaLeuFr57bwFt
czrRNneV3RDv5zJtbPetEZi+5SY0mOdFz2gA9e9PIK3d/lLPljxa9WzrD60b
G8rFx5/ud4TAGVfwA76dOg7l0dPs04j21S0fRBQt+sB+n0ZRAi0SsZ2DHMVr
OiifWOWE9MfpZErKWbItGXpObTo021uUWyDWyl90Rg6E6ZOKQZtZZt4wBZ2D
b2hk/pShd0lf4RD+jNQWn3hvoSlK2P+MZmbqOlLRuMoHAIx7ESJM4ZJ1UxGe
ogr8N9xDzdwibt/XipX+xMFjcW2OxG1M+jxcZNTtJk0kjeWA2AL7cDG+mUia
v4jUvHkhJgHG10ejqwcX7oEVtT5LzExLIS7rfAKJfsv8T2jDinmclXWtKYb/
fZy3FEHDNdUYUdfEgLnUzg3kZwjXGtVCNW2E9rJbin6mKDNOyKD0FIH9jc8f
r9wQYsrWSD05S/frS+uJF0iujKcigAMB+t6fA9OnmOXn3fT4X2MQvVTWSPgg
CgVUW2boFxN3znpgJXehyqZig9z02jXwOQ4GOzrQQa4eOcUBcDO9pv0dGKMv
FT76VcCvt78GOtHfFMYuevyDdLXbdZe4MvIWIduGjFEjnvX59WHT9e1/99k6
1PkiyYnmOPO8k+5AXe+V7OnlMfAWzgwiqPK8JAb/leCxRveZGRklqXLW7Al4
Wt4nqVjorCUdgeGpSARNNtgLJoKg1AoE62oqCp/5b0C52b+za79Zl28FhoQ5
y+1JGyck79fzgE29WxAhWEE81TOXNV2JwEzFGG50XyV5OxbfHFwSQSzYXm2I
FEEbXdhOrIXg9ykv3MPFWHwPIQmhY4hQKukkCbR7a6mgDH2h6PVWlSS4EnKj
UI1CMIcUdjxn/doNy7qjnqEO1zxFsZK7MI280xB7Cx1dhP7GqoOkganCsHjS
HqTtMALySDhbUdyqadnAxevgDCcuwOTFzTZ6A8GE+XfMddyfyhqBNNpIg4gD
2adVNaLqe2wUhn7YRF7pxgoiU6rIG0yF5LtCHw6tlcpwxj50BUcwYi/RNZTq
1AeAiL58O8rVIFusmMnnRESap3QwDrKYbKurVffPLWY3qlCeumyeEehoUZwL
tTnMvDGtBPr7yX8XUEVZrOpbiniQDouoR1xD1EQWiSovHQROal05kqg1AV7f
ZbOfPtwT803aYXAm5Rs3FY6k9iVwLh+GaAnIgTCL38RDW2VRGprB5f43tlmG
0xXX9V4s4RSbDZVpP0Ra0MLiV1P6uxKe0nRFot30SZYKBi8inagfHFarGd7r
SlL+iniE+O0e8PY5XIxhOrflQ/3urIvocZTvF8X7zovLIuBIzzHwvgP1X3tB
utl/CFWISTW3ii5kXFUPQ6hY7EGadbYxXRdCVWtK7fKmg38vzGzKLCQWGr5p
+joM17kybOlbkOxoDCq4E2VhLRBDA3Xxr1op30rDUYBo8J4CTYkuGfM1jiYH
hMaNew2JzDgSr0gG241BMdZeOr/6ao2LLZ0/1kHDgfSzI2+LLZ11tdcYqZF+
I/ogVLgWpOOWFc8bLpFgK5ZvOcqrECzd972gljphMmdsxCSjlY4dZPGk5pVL
pgXcOmLmR27CtJ//CqIDu+fZXx2zI6QlsvKDblx6Nqg7EK3mFhktJftWuLPC
d1hvSb/f63FHX0IZqQ1g5rgjSmVHtrDeEo+8d8gwKeR++XolwDL5hGuCP7Fc
RqV6eD5gFdBUT9yamBsPJv40nD4aOtONyXC7l9th2aLwf6ENC0wLkD3XUQ/I
fQstmV65dWB1ziapKe/e9oH2/IA2XhJK62Qwnea6hQDD6nFWV6WgkSmCGTJN
Aji2os3Xzm11oZdcxruIlhwAbCovoST0gN6QeMbor9u058W2TUx7bDCbUjVU
RENDxnfRREuCyKdu/RaaKJFgdMkAZez14wo4++lZnvlGYKz/xflQ5cfPC8SJ
/cA6pMDncCSdZSgBfn1yENQO2D9Aci6ApnNUyKBbdBsvxzsVd0nYvDLdAOeC
jJecId+ak9VCMdLbimqNQ8t9kZUY8K0ZXbK+t6Wcb1CLfT6WONlEI9uqFeja
K0DDnYCns2s1MYUcIEjTrSKiUZ6WRh1kugoMTtpQaMIOmQZ/KN5fGy4A0ats
LgWG/jEfy7dFz0qXmnYzXhuWnVNqVbS3t4of5UGWAqNXvQ+Sjm7Lhjpkk2j5
tl+5gFCpwq3I+kCif9/RMsFcc39wYGw926LkZGwRK7Xpo/ggtw2nLN3UqIFg
Q0yNR+K0Ydy91o0qOY2fIlv8aP6Y9a8/e8sDKEj1OIFM6DZAZKj9V1NekW9s
J6ShxVRCr/7A20Kq5JmxP9n8UROtF9KRi+F5FyOwm35kPq05kKI07UJsyLeo
4MVGiVs93TCw1g0qZuIOlPU/Ucw8P1yW5t1IxGZdkSdNSVEPpo6Fk4lG6UHy
6UqQbybHkDw9I6wDSu6ijjIKeFcBWdb/neY/qLjXKE4IfU9GsiXVZ4e1S1MB
YvekhGBP+F5qwXFqxte54WX66CE1VyH/Ma/VnynhNsFYViZdsyyrLBDxCfmh
Ha7jNIrmwn8v/VETJcCiU9dw5Io+sajLTktrlXcMmjF9Sa9Tl+mdEUa1NyMG
JJCv33j3Lo6jZIbenJDO8i4mZS5bsAfGCLeX7UDeVisXldkdz14++J926K3R
62w+ainiWu1jzFquWoLQk02hLP+HpvwUn0VLQ1h7/vmUMkBCSHiLKnhNtSmN
hisLtxPykvWvVJPsJV1cGBh6SPpPXrbpN/3e49urjNONwMOMF/Wi9ilmb+1Z
IAEXzs2Q0KtZ9YmCbS/KN7MsMzj99X9GiFKv5Yflo0TO6BWqHrgTdDUg7oSt
r7WpvDkI2UodtgglnIHQWM8jzO1ct5aeuWjFJnWhn2xQ1iCjANV9uzMxyVOI
GNBSr5CAKWItuP2Vl9Ox/FbJx7etK+aJjcl9nVC68RakAT35/w7xoWJqeq2D
AjsnhldIX43jgp5rClzzVvuWDkTVZEa9Ozo0jtHpecn6YxSS+ipPSKlbkOnR
PjBLS0ypDULOxc9ksOjW/AcPCfRw6wBnOoFRjER41Da6bKNh2/qMPqvN6jTr
sW+euh8vfyiVRkjs62ikHrYyagVpDjj6RCm0ZW6TAUqqbjAPGH66XZ0BwjuK
5iwqb2eomOaouplaxrqUiiRMjVmeaAvUTqvhzv6KNcqRds8jDStn8JNdZunv
V0xvo5ZW6yqrja6fJkp5gajIhud3iaCS6pZ/6uOZCZqyDE6b0eTxV35a+xn6
dqugJCkie0Msv7Lx3Zgqj348X+NXAm1CkGrrMXjDYN7QS+Mcisij2uF5chR5
j7V8BckgPRErcxcljISOjpdV3EVqygyJ4zZyeNnCZpM/VwLtYJwl/G1SI8JV
cn/3ZZVox6mAOSqIK9UqIQPbD5oMQlzdRjJlYKkhjO6dnLWqzIfP1DvU/D86
xRxw0hf0D1EMikRyK6DyKCwPIF2o5lpeL/vAORBd3VahJdmQ4Vb9pEEnaNwS
sR2hqVWXr6ioAF4DVdl4ZZnDa5H5OSbFVs3pVc0sa3XIZS90l1lvR5+vP5RH
xiyxXZquhP9WN/J4BZnxdKCFd8WYUZisN4n96IOD6yQ7Je70cz2KBizoVFux
YFYVu2MocEpzH7BtyVuuSDYskde0VjfJpwGNmrk5/eeoiD/vc5UTKn1U92en
Qz2b7crOscH9OBH9FMJGrH7KQ6MfZRSVT0Q3qklqtYnc1ttliuVO0B1jlrLt
A6UI39RRxvl8JCO+C4nQGzuzSjAFvbDF5ZxIXGnxMthHKlKiIRdovb7ya9rU
c46b3lydRxaByetfl2JM58FcEnkHWLpBkD+LMUJaO0f0bf0A6mD3gS1OSHBv
XaKB7CFmYSEO4oNhObeAy7hJ1Zt8BKt+RQTzPQdozCt/KJUoF/N3aOUNSuFA
sGxri06ATpiQlyP0tahf85TWKuBnQ47mZug/hWq18gf1bNcGh6loA1o2tRPd
HbNijrDno0x49+gqZidQymN1GODtWTeuCArZq8x+dPnlv7nXHCMAepnnDcyh
lC7Be05GYtFvO6gf2MX48ACG2ZAK6gxyetLWuXkaaJdN4H5rpJW397zoxrpv
ECqqYl6ziLGeJw9rmCDXWpmU3JnObsaCCOk9DQfaY9i96oDwupODpGFdiYYO
M5jz7GZJhcfw4xUF/e1J7wMbTQaVGt7njAoxO2B2ipXK2y55plppTPBkqwPZ
KZmRukR0xhgupXdzUt/ksxZvaWZNmwhf0Zu+iyjMglu15nNOMQnvD526bj1M
zK6fNE2D13bmRFNyTkfwg3gsRF0o82bGRPFMkjpiMuema9UW8R6c0X17ANCr
2xRqk3ceE9F8LmpROxEi9FxD1KlaKoFmSDFPJaFP+C5Db730UUJ/L1trOchg
NLJfhITS4CuVfWdpxJ/tnLYUodr/69j1HuJ10TcgIwKlxhcLgHjSX1uCd1Bm
9rU4JPY8b9OKbP1A0AXBvLw/n/VjlHWB+ZyiDNWgpD/nQB8HCAEuCDEfU9Gm
4K8S7MJcmmASHJEYMxALB1izm0SzD3oTxmAThF3I/X567QjeCyt5S9IcAQbI
ox9UOxMoMOBATmAsROFha11yvjMyJ3wS2xuHRSpTC9lWLfu93LZfM8IB9KM5
RC79b35LAAnSUh4tytRsSUU0GvOsX1u84ERVzU+4bOhzBJGJsz22g7II6VSZ
4hlc0Oy6Oxi3PX0sK3D2+nMgHNsLQGdbQFAbcljvZ3Pr5QPUmuTdeXo4swZK
R9osMP56mQN1R/Mn9ZgRKkgYIweBEJYrSVzytL9so3G9k+QiGvLRJu0bw504
d4XBJ1PDRgB5tWWzFn8+VelcYprU15NmJ1Kl2kjeDwzXC0MceSqEzVZe+Sku
UZXPDGRrXdrbgpNMeW89slM4S3MyWBaTEMnRr1IA3FwT4onqdA0kwqF3oX9g
hjEGN9aF2le65DdVy/NlO5M9ZRT2TUBQOjcG0tPFXbNluHQGG0rAcmKTfbfQ
KSn37hkGTmATACY1Sjb7DoKWuz3jDDCut3qeTo5Zpjv4vtfGDMyRvA0uEBD0
hHtTqCZ/9ywnPL82Z7N/ZxTfiEP8sTw/AwpSEwOhPgghzA7RdBsXC1189IUy
qX9jQ3MbgmSxmCJ2k/DpYCvCMQUX6W85bx0BT7TYlRXULjxf6wrEUM+WLTK5
SjgfM+KNxuv0E1ZVmR+r+AWniJOppuIlKvXwjOkE0zDPx7zmNo7QwsYvhh3s
uflEzp5CahIzmARXGzF7MNnZoOnBIZfeGhLXsFtJ3qfc+jN3Yv+yyo/8CwgI
bemVvgzJwiYmFGb2S+An4EkoSAvwOsWTo8w9kNhm0vztdQT2ICWaxTZbzvFj
vw17ftjORYJaKWnu4YtmxakF+/px8AESHM8aVnUTH3/rzQXpqihzGzaOenN2
xJlSwXFyglLYG6gS8YQrI3lY+0+Tah/7pq8oVl6pZ4LUaZs1HUhDliwXByJm
hj/K3vut2XrqlxOJ27TyjhvwU4ZfY+PK78wHtzqOrfU1URCyQr/C6JWQ5t/w
kvLsZGpw5CGwgJL1QWXu9Ukbp4F/d+lzdhw5cEW2BAbY+so8pKF8fDFIQow7
yFQvvbCfigOgDs8Bskn3F5dT4cT5WQP54fbxS0x1VF2Apz/a028ndXfZzE/M
cBGaUm6Y6Uf5ebVSCpixAkvPCRLXr9esM9dAsYtP64iVhH460PDO9xBaYvgk
POHquNvCD/TGb/QKIe+Yv2GegJEt8LYUJ7jYZ84CWebAeOKygYVf99RMx6yg
sQzDEEuqMjsq43nGSXJT+5ojqeitLubfhTMlUM/R9mWz40Fzb3I78rnDDE31
cPS/rm6bdnSaBxszvWql+LSdfPU7sySCExR2pq1TNr2OOXvMoEe2F/pXwM7L
MtsTeoRr3rqR8+X6mLC+q1Jjx3YkRE05y70dBUHFGa6O8lcVHajhaQwy78d3
A3T9tqJYcRVhNpoEB4QY05fGwYPROjdOpHWHrcCaPRI7bPZgVoQEmTl1mD1C
LqoQq/tmJc6OYeU+D6dENV7Iz9MWIHsOyh30dZbVesCiZiQLEv4lUN/jyPmx
aO7OB8DZqhBNfvjs3tOq1UsLxHR3LlmuJg++vCWhYnaUipnUjQ9EoizgdF+9
lPbWlI3vJiP2D7vu0iOyLtJQSF2LNQo0XzMFVIyAT7rg9y9j3DeKOODv7w5B
ruHcIoxqqpluYqn/Q/BWdgJXDtj9lOZIlslIhyrTK/RcSJA/LWY5Wi78fLGT
tIsszBSamsTawpqP06vwTVM4fF+dslEcGd5XXk4wjvkRTaJRHUTmvR2kednT
jYDciaedhE1PE2glJJGuV6VfVBpLJ2uLzaCUtP2YPGQH8z5q2fa+GOqJQuAx
lxMlHxM+NAGvYFXdjv+91xzfjeXN5uRR2FZNVys6rhsb1r+FwNsXwsLnKG7B
XsjUw284t3zdsO3CaZX9VsPOoUM/9M3u+1WTJ2HJNlvSXW4+8fRedCo0bfuH
i8baMmhxDiGrePqRxQSob0YkBMuvIk+N8AIktQUmlMWH6sKEDBNX163KO7Jc
5wCFIU0VHtoptfpy58KKjhLLZDx7lXl2HIm2rG8Dk/4yVxg3V3vPRoCaybI6
0QfJ8mx/CkIFsB+TbFs1yzUH9rST8BpYsUczccSyhQ1lgE9TjqtPCA6Qg4Fc
Gbgtkxd8DCr0J98JBiA7y1ET6maoqkzboitprkJGaKfgZcC5KHfya7ii/Rzv
/HVKKpxUT7eUKjZQkaArXD0vtPtbXGO5YTnSXn0TUyTFItmwnFcEOTErbloG
dUh6HR8q68q7zzTEJrPri2/2Fn4135zNAxGINX453Un1dB1FW24T+pndSRLY
S6OYNhcL8x2KKm3NSvJ7UuJBauPtu4KyVcNanE38LgV3anwelND4c88BJes3
Cl5QcDiWYmKOLd6ZDyJ0d+T6OsfQlhOGhCcHdUjq5a9Bh+wzn5kT5JNzyNQm
FSC9udx30HNXunVGDctL8obSO4OzJsqBd58uVvFBX44BP9vQdupV+cKBWQj6
7euS1kPrVewA6yhG57wIS9Y4Gh0whyaWs/7OmCwME7kSmGaZVzHTQWANxPqI
6Hb/FGS+Lq6KJtJpOTWicDhPyRrjKRBp5j9UcRN42wmy75QVX6YlmuIDYr19
TJK9Fpao+MfKi7VVICRfCtlIlKm/Sobba66eA1EaGGaFjErI7+RoyfA96GTb
KAh+7TJn1mmGdhv8LAh/Og1waIOofNlOWKIXNmkEKkhQiwvl6dwmfm9jVJe5
wSOCphM2o/K/bcaS9QcTTOLI5UDgMTSV4XjTcAp6A8biNngUXkfX+jgRSsBn
UKh5VTfoKe2ULVK+9BdVL4RzLrabKIW7AxYVwyjVFxlVAglzSdpJfCEHYCsN
TUyFwUKR3w8+o1FFmPRe5jTZ3rKl3Mcf0PIzlqakgzDFFwtDB9OIeHN62+WC
m4DMYwsM8UQRtG/CBJA2aBsJcXpXRwJitkbhzIZpPCBevyOauncQ43qsnvK3
yIeBBB/i8pqB+cnwa/Dk2IJbcLfMwPNLRStsDzFGj+AX7aa7lGfcXokae/hd
1rC+7ZqiSIxDp29pMTNm/HA2KEADQo6Phc0eQA1PBMeciiUDBFgS9ZwdWytL
2DiHkyFRspxRxIlYZ77XrzlohXx6MjmgMlE0sDb2uHZCYD+se+PbGpuT6DDC
7VRRIn585BHJMFrhALSARrFATCtQuoewZVLpxiLWbarjZg78AHL2fcbzdGYc
jl7ab6T8O3IPh6lAnvxX8Rz/a864xtkFWKyRqMpZ/rIZDQKvRjNQU5+DDL8I
F5gnuPGFKQ+ZJRQILj1OoSoHNpDwjl5wWRwFEXzAkgQFXumHgY1S/8kOrGk7
+i1I1nO5qqHiOmvcaYoFN1ieml7LBx7y/XVD81x3gAq01OkQLTAifnhz4WnE
JlWBvXA9dWC5delh7bGXQBtzmV2FCY5fxGFUYW4Bd/AekR1DhI0ljV+FeJ8U
zCswJiH7ZZe2cbO4XGE6ypo2GZ+npwJkUKPRlds/xbs7FH6qZNKIoCtFFnic
uk5hjYRallFSjoBDSf68wEXasVKVq30wKVvm8OclptdlzZYbRlve/24E4+sk
HdofJf/Mi+h/rcnThQ/V+a/ALUvpn6KB39ptnyXUOfMxrXl0Qvj54SsRDNUs
iRZkBEVU82ZXN7tw8O/TnwV1R0+DR2eLrcG++OZZKdUb5ANWnD+QJfGafuuX
/qcvfLh7ri4WmLjtAe2h++zGLQTjDW8Au3cIKWbLhw9cxUc75WWNuwh7H0O9
/weitsII46dymzuV5qefXDhZJH7jrusMWiw4EcXtnuqSZ9oZDekyDuTp8lM1
2/HUx+y/J5LNn80KjgI39hSlruglf1YxhuXTg3zFx83wIW9Z55Bl6tdzKOz8
IFJdj84cwRu1QPNdIpqBMU/8HbpGE3W/FovXNKc6d4c8OHjoF6HQ2gmnnCJo
oTtyAHXpfDRKUgOZ700rCaeewZr12bfSBktPhogiFYMBc0FNIGfey8nUrbPR
JJEWJPKCt0Dma2HeUCnrEH5l90vry/qUYzD36NZc6UpOc1V45oLXYmnNonHq
yZbrKhLyUh3zw4H74tHnvYKlo4m9p4GF0zdX/448BcYcff7p8mzBE0dJAISW
jKsjz/Pd5yAbUb6yPJVyJYDPIERBXjfzB3H8jHKQH23feQej6khuY8L4sKjX
OwlzEndarBFfa4zXNHRspHuuSvmLUV3IPA78TBqD104E9EzopS2WpR4WRQzT
eluBk6ztX5e3GSHVC1QRcRkIrB7X55QpgLAQ2DzSKbrFQstTBqCaLU04W4jr
AH4Khqeb9cJg/CctnQ5yEpjPX0oWD/d4wuayiKk+m2bSHYCsa8zKc2IwhZm4
9OGZgNnM896h8G9GKq5iBlruLRlGkegNnhokPoIvdrWvqSf0nBR9EZ7rafVl
3+XFoQIQACrXtirn1UVQXnIi2m69P4cOuYM9E7hvdqkwmBnxTYs4PKdRt529
t4agwS5he7KzGLRvMMLTN533N7YYr0UeeJUQopfU6Inv+0LtlIipyMYiODcv
WpGGsxnujMpcbm+0MlpA0En5K5AgYZdkZGVaziBcMOIrwwhL4dfFWZjQ0K9r
1Y7U8FGSDEV98snkdOQsOpO5E9e+bDjRNt+W0j0quZkiJ4jXOJLBtRdG1b1E
HDW2jLBF7d2CQ30x5UiGOtgSk7rxc9cX//Hged9JSE0s9sccF/Tj4c0SlyoD
w89jOHo8uOEX7QI1MbJa9H6da/Ohw5KiLklWXKOWw/u64Zj0TOovtV4ppFgp
c5MXMAl0ImnZhrO7VrDWXJP5OSX+Gxr72+EFusEjCMXhj/80RnRLOWpqcMRj
ne6fDoJHxqmXvUuj3EyyVzfiSqcbc9Rj1FQebv29b/dNPoiBFd+kLhmpYQPS
yPPsqsBBxKFnQnd9tAfeIJwEfKHFhlW8zREscH/Cx84vBPw+txMag1gFNmFY
p4xH4/KJhY/btDCi0nMQwR+dnzcgGGZBIq1m/ggxDfFix/JKPzBz7kHxDQbv
XjabbI4ckl2KocYjLvvi1EyetxXFoKOHwrQyWMUSLTzqtxosCO7RBVxR/kga
GLDmytmUxeQMRD4rRfb0q07+YwdUF2GM2bz7LDscQuVDf4/iLYyQVfSN66zb
pqNt5aB6Sam/uGqSx6v7TVMmnY6cox97AlS/14t9qom9HnGfXO/wUYmv/kxW
7ENS422Z61QoWuThOWA+IwETv4U0++D08eaiNqBIirBQttrBC88USYl3IIjc
R7Ngl6aaV6U3eL9rIdPo2Da2CZH2JlTk7UIg2a9Vz3tVaWK0VSR05gBPoBKu
XnaCEWkeAWDpmeAsfoZmdeye9f54otTYmhjoceMrxOxRJsr247cSLtpzUebX
6p03cUcIqKg0y9bVcGiX8LgPfBa4M/Ll8U2z5uhXDaCmZXfZwlNcGGF8Rx8K
AMXKEcfw9xYALX0kHTisadECASHzuN3Ra6yh2TZ1IuunTodjS7AyTYxFjWcY
WBAt2oBPmZfK+GPs8ZKIdld3jtx/7aS3mLSdaUjOhb9L+QVxSwDOhHqIfGF3
z85mJY1vkftPnIz7Eb4yFXb/4KUqRE35lMtQwdWc/dNm1QniHQ65E4f9qzK7
w5bUMSX9aSWKrmimBEe1ywn7nL/EXi1TEtBw8mGlOSAmvLRbwGUbo6LyhRl8
moQI4rbqUMWSzR/yX9ge051xfXZgWpi8+Y5jPfJGWSScg5tkMzcSp8qucnCM
ObIElb38h+lq2OVMVl+X/Y9tprvTpZSnMOd7CHu9yyJfe/Qfik9rE5vjB7vT
r5ByO0c97ah3SWKf9HQcQTpes9JyRmWZyP/XWJNhgglAKhIEcDyn/0cO0iKs
JudVg1TwebOm9gnPTifjtFBObhnbGBDpkfaEzosdNsFpYnsWenWcjrtblJSf
3AxkTVd/+OuHkSqF7Ym4jEhlbh7HEQNnDtRCKo/W2CqUrrW7C+J9y2hsYqsi
eo0TvDNc1HvR8omb+IGrIrBe1F+aWKICAiE8GFsGMzrYmArEXtQueNfUlD/l
EQL50LD2dBgwz5RYDUJy+rRaWimr/tdjAV64aLv2dzCPlsU4XrMIjM0Bs/Wn
3BT0hhJDSAxipCOJ0I7b5GQgAwt0aPdVG3dm9070A1bVrm6c7OuQWzD+1EfY
dOKhlSMQ+GcrFO0+F0mNFxEHHS13sl4/A+ph90ok2OAttdMSSvLlk4c7/C93
YKEcNHKyYASPTVEcJu0MnPPdsgWVXeLwjO5JaYGVQ88LTWA3fw56ol98nxRa
AGocr77nr/aUrfwc7gBIAMMhbEeONsyrrdFsz2w42Nsd5ULjIoEWt6RR4XMS
grXp5HqMYgZPf/KJCcs2rZuaq8Dfs3S9NS+xZTJRy/tv8XV65r4k4AUWnjLH
fHU5x36xIa7M+xH5LF9yhhYrVF29UIpIhvh2uAbXgpmna8WzIH+v4E+TVnxH
5DWzG5uIx4y1Xw9PhWUd2tb3z0wSLtr367LvlvVFNyOzvVSqV0PRJR9wt2iQ
vAy2pEeh2iYTOrilOtSIRv21bXhBT0QG9X+1mnIfrqkQ8PXClQgwrpXOt4L9
nrnSpGgzbU2DNVOxPlGnLIU+VwjEOlL5esLb/OxJKOg9XukWfvHEXGy+I2yI
h76eC7KE9Z+DIVaIxdIYXfPRFBY9OiMdnu/V554ZSYLc/WqiTK/aG3mmGTMY
HyV8GU1M3bjBriX+iqXz42whNlSBQS97FUDV1w49VN4ZWYDswVbOQTqP5s/v
Wtdf7X8ZZq32eYmR3ZMJhpLzVWTRs7BBpmGaC7RmrJO/AzS2A5fpLO9Ik0X2
OWZamISLgEiVtgdmOMPLprX2caibYC5p9a0aVq8M0c2I89YqtuAGnFvVZs+M
xX0I/Ee94Dee0FKo9kyGRYoUlfn9WYJnA7FPhRSP9imHkTHKlrrfMeCHAkiH
Z2Nut01lib7fV2HqzcMFgWZpOCZWPbiafUNA92lX8w+izeRp5aqzHtnNhfi/
yklU3b+jqcPtwv0RkSVpzv1h/yzygfK0UvkrO8S3CNAwodEdPQinR/k4YWkR
wo5gddYLPhtTA/1I/Vqy7j+kLxYz7myXmSvQ/+P81aKQLK0rHD3MO41fRHc5
xSHYL3dfSVAaCpBoieWFhKdB/gx80ZcOS0uZCEOmjeVl4aXVfwV26Gsb6rQh
TOJY0F50vOzzVBiq3+djhk70EuqZnPaDYUBuC0Ezl/fLFtXLaJpWf6vrtTJS
1CNOMqdpG/gjzC6fsFNnnS2aQuHo/e3hC+ciUXgqQfZ1OZL4hcrtqWseLjJM
YVtsgeiilEH329RXd49KoEP4e66QnZP7nVz12ja9oqtN/CsutvnPyYn9xomx
Aczhz2JzCpWJqLoLJF2jr1W4JoCvLUQOOgrBDuQGYqjB9srhLJeOjxm6mRJM
OSbM1FQKfPoPgsiHDQuQdBV4yCXjVIJO+ceuXMfzJWzVW/7npKoPF+R7nD8O
7yGD5cda0b03CmfwI3szppx2lqmE6K1ZSKym9JMEBFS1tlnQqCk49wMY5JHN
jvXbl4mM51r3A/rkZpwOq6JwmHe/amRZRHELldPXzkw0qfSDWGUc9ovLtZe7
X8MsUDWMsLZYqV5EDEqZxAIUv9yZxvKKlSJc2qUCIdwn271YavQHfPCEhOfg
PDgQX+5UoXvK+s0jKqbFq88k5vuFVrouVSkI8WOoBK1d4HIm7X2sSCa1SGgy
l3adW2gkRcrV1wHJjmleWGRNglzhFHCd1ntQ75O6abVhYXfGW607/ERjIwI8
+tjnMa5ffjE00Rbsttbyq5tg+Agds5f/wz58rMmBJv5ej5OVImQoYMM3xUd2
qBTqBit4GWsQ3+rCPojlxR52AlErU/sIsIeSrL2kmSZUTHUoWQNtcu2WL6kz
uRh0VqtAFGrGdV4CsLSwkmcY41HxZ6udUeRvWjMlJEieuSac8VdxtRPOmwpL
/BcFZmMxuyrbarbhu95daxI0YBtk6nD5Nd2TVuNi5jSS3U8hQi7nDNXRW9P5
vhYB/O8SBKY/Xx07sIaTGS9P0D9NCzdf5SVo3gcHTiQ3Dm8adPfEgOaZTaan
N5W5dBZQWPGhP43dDjCi3imXnLy7rVRU0UuvuOG5T5U8OX+0XOxo9bS/s46X
hG4p9x+JJrdgHw5vbjUr+T9ovopmMJ/gfiSw8rJOwNn884yxfFcS77vFXZ2E
mBxxFojySGI1GhKOWjVr/cVmYqn5HhpC3WP2y8GKTBSqRLWNgiGJosiXg4SF
H3FMpEZPGICIy4yX+fHGhc292fBOZpBQrhUmtEOOhoZhXfYdoyLG+wNbcTFu
MSf7wxkiZ6JChOF8vi/lwq/aLoukAJSkRZA2R5uXRiuliBmSkOXqvtmxlsgh
biwvxkVXjwZn67JjybOwkdQ6ViC+OWAqvKwbBlxdKrIifm86fsBqaxBhn451
Z57vGOTnp7O1x6FJ4Ln0HOul0INMW1MjE3ycTYxU+Ey7cTkfyoRTFZndzvRw
7pKeazFEe2ASE87q9PL/edbIlAd7tnS7iNlDzeOYZkndIUUDej1pSEU3MHbh
ADVoe0IhfT4V0uq5gy2jxBfREC9XzLXv7QCr/tb3h+nUFdnV0anvZF3wkRMY
fv9J58ZuiP2G8fA/nHGaxsHGx67niCsrB9QI3BFBtyk4SoiBsXG1IvjKpHd4
/HbJjhJoLB6spkTQTpe40mTJY3wMD3MxiAUTCu0gccEUMbQ6RJEPb6a3D2jW
sn5Sb2U0FUeOW2oSXxx045+MQO8ZDtklfSeVYLE0GDlSz81lDOH9WpNnAEOU
Q+BbB5/AhZv/gyhlGfz3gMS+GV4eSQ1mmL5vl6s49eIsjxehKEKMTaqU+qo4
eA92VjxLVNgtDKKI8dGMTfy4DYKM2OlFtHcWuSSA33G5VDmsFWdkrncBfPcO
5a8XJ8rZuGx2feQa1aTodlA3kUqEQhktXY8+Rs6yFRfzob7xWJuaj4Rb7Eiz
YXvNQUV/mONXFaKjsCPnRuHFRskRBAH10Smkh0n639sWJi5adiC0YWkVO2y1
qfMI4w4jbPWE8Y6P4mtSHX2oHEM7lbG/tGn+NynCzR0F+tWWozVJ3odlCOOM
xUDsCmxorwc7XpPt4/v5ys83Sgn9ooHQq/Bc1sBdRtAonrdxfhcW2xOWkI3U
zuRtC4/W4+cBnAzApYVu8KFiuq35eE6w2l7WNIIPJ1mRQgeAfWh5MLcOfGEF
4veazWERzFqqjfdJW80zR21IqKbe4fRH7T3c4XXLVBRpybXSz/cWrjrY52SB
mAhNfilV87CcPQJInSQXIlCRXjOKvAXKebE9EdvboxPW9xkizSCMe//sbN15
fAd32BGQ7wggNZjtijmTWeAfg2m/XC3hd/KdktDfDf129yQFwmq2g8UBy0Qq
suvLUWPKNPoe494XWdhYxlAy1C5n2aUbmMu+BgPpuzooPqFfYPklS18rWooN
8+0EBtlurMh5GYCb+3EFU3SpyJUTm+R1mU1M9zIAMpBgeScntOuYStdz5zab
vMxnmO2YqR9q+ybnuDDCY4A0XgYF8FI4Hz8DeLGwtmKt7KUPKEgA+OFCLnWW
X2tg2XWnNDTVOfADfmw61gvDXBkv0WNyjec/8xX40CidFf5UP/9w/QIAUMHD
1GUyLhEbQVtiScXnYnuLG9yVIHJowRwHGlaK/7CU6C58vnVOBAiY1QtNE3nW
8s7ygnz1mlcLkQAzKGuwqLzBPsS3KPrx6sTZEwIaX45bC5lD2RgAR+hpZ92v
jRmG2x1ts/TumxPkcAt9yHxTNhrojko/J0J+E0OS8rBGEwsWIcpfkzDHummQ
pk1SoD7zZHZF0UXPwkVGrTBBeM6est9/+VPgW366Do0Xj/10KlnzYbag0ywV
UwuSBxQwPpKXPjgwM0afkNUCu6KexHXEAAfeGKXZ9wR7n3DBr/wUp0JTzi8J
maM81eP/TfLuarztaWzxwqCRts8Vs28H3zHWbBA56+d5FAl69c3v0jh2Eh19
dx53vgVxwbeXT7kvIqumGDC6goiKTGXguxsmrzvSC2pz7chSMnHAkhov3ytJ
x9YpPPmc0EpBSk+V++DKueuhHlpp4Vs0Zs5AkfkiYFFEoMyC+e8VW8B3SxNe
wwYE1VDa67V7FhlmqlS2MfliWH7IZqNMnTti24U1TY0Wc13oJFl1Te9qzXQ3
d0eweUTInkjbAUFYptuWaSReaJ/2H4zEycqR40QnL07IGUhV9UqhHpuiSwRN
RG77/kgvGct5GwffTOTyFC1X5WqzbTwlajWxJu7eKjQu4mkVOnOsHDGOBke+
fmFm3A5y37outvmS/cMw1UOae9MLdHuK4pcmxJZfJHUEfFwr6zjqtuYZwKEX
kG6WZztJ0iY5A7liFhwQMsl1Z9D5PQ8cSw45qPA7so0b062trDeEfKm8whNe
1dml8F8uQp4OyzGe79jlwSSmJHpi1EFK6NOhu/eJuaQGfTgU5xRDlxwcO4bv
GkxXbo1NoZ1DIspxrNCC5lUjTi0Z9xO/0t8Cl6+7vEAc+hv1mfAtIPYs5gjO
kkANB9uT8R0VNlLxp/KzqRVOAEL+Q+icMp4+oGCzyqh711ESXP1G2GGmIh3j
F8Ia3DH8vSmOAMrNIAKhoS6u6dShoAcCIYm0+1HKuavmLBRRa0/QMUEqWWab
Un/6fs05OEH9CL5XEXfHp2rKou9wts7Nfe2ob7CCk0yh7op3G8sngtOH3uU1
1ZfvQfMXrfFnfMlNlX487f//2o5ghnvRH9i7iNCv+dH+pQNgmcIId+pkIcHC
znYh3PFHChK4xsQowE02CYfyXeqo8OY+KTh7iwKlCsbAHRvgL1nhQ1FxJQj5
5n4hwytBrQudbT26twERQcYlT43HLkVXmW2pRVDQakRuihQ7YrcnSkEF92RQ
VzYPBj2kDPKmwtRlsqjoHCgN5oBrjpn8iJsQFM6nX0mc9gmkKcDsyRxZgUhB
LSn/XHGYvQyIwN8KaSiMro0tD4x1bwA9M5lJ3gOzqyFP2mRDwodYUa2kqSJ3
nSo1k98jzVooeLfBhWQSIq3qqXWJK2rirK9+qvUc211LxTlWjGBgoz94ci/u
HBGZ0NW3vzy0WYTjwsaW5ZaEIFWgBbQQzLMer90vSDisjZcHVZdNHdralXeW
0BdU84n/89+3nDah1vKaQrtgLwqxV9Zxv3ITCJZHomWdWk2wuHyYnXQm7Hep
rUpZM2zJ+9eQgaeKlyYruahe7gIXq6At/jRU2Dj6D2blvkIm07KkL31WJxkl
NL74sh6LhfiCRA0MfNZV5+9dUfOIwR35/f7f5vNBegOtLHRFvdt/ljyjyUye
KGSKSahaOpN2lM/TkBOH/xlOvxEMWRAoCchjOhLWhWTkNx+ypVkkCRADp25f
w6sAfhVHrWQnyO8Oz9gDaWe9aFKtv/pNaWU1GA4aiSUoAaLpstj2QOCLd1f5
XzpCzyd1EWC9m+Q/JBM4NHj5Mi36OvULoavjwcLRNPlb3rHwXFF/rXjQLewp
hmd9bXalchQC9OKPJZUg/hMkE+cVpyoNvpS/A9Acokjg+4u72ZgqPJk59pZ0
XwSSjHcu0WB0evNwBdyEgUbzzpA44PAoEBXRWvK/a5/MO2gnc6FUmwJE3r4j
gLdoxlaIdurIFgXmW8qo264d3MO7uaB4vo7lJqXGiB9A1znQPV/4Apcamehf
uehGMNe5JRq6w05+lCzlqKJS/glmMoIPa/rpj9g3bWqxwzhyKc32O4AU/lYZ
v6oORDvKaB9LDB33EaCge1mqDXoD06+a2VBwyYDighDbkZ8Fhn2V2ilkCSap
ggqSkuYpIxxHunZ/aJ5M5aLzkIPLBg5E44e1bsKsWKKHy255mCJR1L77ExUE
1yTYPEgpv43sGGx6aW71sAlASniKo3Y8EFspOKEMNdYrPLHdfWhhGcXlWot1
OwpaNxN5q6+fq9SHj7oMPIWC9T+iMHR9ij/2tvPWHuDOUoPad011a6sc0ewR
iuEx8IsPrD7KPk4CcsTw/xfqnGpo3EhlWEREEbOLFHVa21gknSqATa0w5dCl
v2rTxsSrgMJnpltNO3Lhb0y5wjjT3er8GzbBpSmHtHH1ifvrqkciKD+PLdJh
XzGtmYV7ESiy0hEo68dc97Fk2kk1rqR8gKFtXDqf1Qlyqn83DVCa1ReiI60e
Y6ax/0yejJyckQZ9sB/HGce1f8ENxvp6+1Ub2n3hQXEzdSIj/Bv3+fY1wwnA
+I4FJo2YGj3FKkVwQRc3fkyxD9ubvjAphbACeif16X4A4lk024DiVKxc8m2P
fnPQbUPeHOnzOs+H60c2i03Bcx3CnJgYakWY5QWvOEFgEb9dXQMH+4A1Uq24
MDgaEIHae/B4zd46nC1Pg3EcRYsxgi3EKEXailtMDiSql0nkYxrTtkZm6F8p
SAZodS2YR7M99Bu9VK3jYlCA6UDFZkXLoLp9QmFrECNHJe3t5IIjkBIQjmoN
Wh+3L9vY1V7rDC1/a0I3JRq/zIRu8fxkohuXq8LkJG8ff9UsGTSK4sYo1AEJ
PcPFJmXRiOatw7S4lTQ7cSeP/ihfSbWH2zdcRLgs7sl6v5CbPVRGaTSzminG
R+bSRhPWdpW9mcIdVXnKfTew/X2vtnvBOHH+sat7ufrB4w9/2ZGtShgj8GWo
jLgjPKiO3X5VGHcFfhcr6pM865gdf52n+2idqFQqyfC3uxbeMIV5+3jert8k
ZCEKFeM9XKd62NOiGIRwrnju364Dr4/YVlv3YBO8jbQDelIS1emb2dTf/95F
utNs30sIm78ECq73XBFNAUF9Ceew3g+i6SybRgr/FAl0UHW0eyuchJcVyAoM
NFcnte9tG/HLvbCfuPFGl0AAY0ZY7lCqJwAAhEqWRMpe2qA695yjlg4p+PWi
EMAsuqG1c5qevTXfG+4L9Z2ml2aVmFUocix5WX4LaAWHC8zXPuEuRMq4Fv3R
DX+5/WboZP0dcZACQMES1I0YZ6sHQF6fZywP/JxMA5DhcZ2opsQIU3YFrQj8
a04c3W839F4nVaFZ4hQKki+7EnjyWjNCHbEA5pYW1D/u00ti2/7Bpjj0IizB
Dzswdx0zswq6CYG2Tpay74ON5g9aItV47snrewXnSK29IpxgJpaPMGJTN9S1
hY63s6EcwsT4847kWfRZlEWaqqGoayC8OmCcBsU3h3mJ8DgF20ISTrDoWBMR
sAiTXTDKDfxM4PirOtE1K3NkVLPI2vEkiO94pZdAgPi7JtfnyPTJWJGS8GWL
+3IoDmPKPDQyN7jMGH4p9hMKKixOS+ebyFt3RfL37jip4bCDPAX4Qwn4GcM5
jrF5+pkdHC+aqpisq39B7Dmar2Fzl5OrhXudW/hhWN1oZ5jG/+crRFaJKwDW
D4inhtrEHb/+OHXWDAUBM0FXfHWP6QMYX1Yha4Qu0grL8OAB5XRrrSNsbbGE
YXqGPROVFy/bWHwMtfDrdzqXbwV3GhKdXnfVN3decqIhHZzQFt7UIUhdeaiM
OvRO5Hxw2x39WE+gYHbqmLm46bEkkSncK8vqYTiHLhMkaVlAUZ/tz/o2yG0G
iRgPBR06szjihTh6QOufmkPqDbWwquZpBli6ie8MPHeoSCbqG+/RH/XRcy4C
XxAypMqhenDqXV9kKTsnevrEZUZUxvgTJxkBxXgCZpDzN/23x1YG3oL7a5ze
zfNxBdHc0o0jgEpe6tFv/k8SJ+T9BdGLtg2AQLH8PDMQFSSaEgTaDT79uF1L
xDEU/BOWDeThJIgXe2kGUornmW7JAzYG54itw6JBEq9Kp9ZbT6JX4RBi4pjG
pIyd3dDDWrNeMJoETbGcKurRfl/GUEdVgYMXsdDugssemNv+c4sctjy2PbwW
aQ2AyrfJIHV+MBgBUDN0D3XBQY3wjF4hxNLJCrSDTlrOoQK8TkpnH60Y/bVa
sPq9Gne7BY+w1USKTGjqMTfTdjD19IQMjK11uqYQhUSYOJJPOPUakcgareUT
skaUNpb6S6m1luJ5U7jIWIYEZlCVlL2Ddvcd3GxM1CjSfp4ZUebucacdsUVB
yP+WHJIp32OUHy9kesElA38msZTSPlCDnI1COG09mBbszHkTT9y2cNqTjLkr
AwnVGEv1nkekZqlY23d4gmsVki9Fgv3BVWYRMWc/9hCkHt6ndLiIkeRAKQ7s
SjnrPK9XCQjucRGLD+2MrxiY2juVdhjXWWNjkj2zHAnnVJlwZAc1ckCOYmaU
TDEpqG21vd283RhxMBJWas8zkd+HP1fUjE1hPNenyhcjmte123Nf9NcGe1xE
ulur5N5hKn+Y0b7/9GroaOj0jwA+BJmeQ6U0q11qyZQ9QXEkorhAjJMAl2GZ
g78NBxl8cz+z5JzxfMsuil3qCMaR11PPvdp0GJEz4vohPFc/7iwsAjlUmfP6
tsiddCx/q8MY4WiBQyro0xsaGY3Rav4z6yf9Ejc6npD+L8bNzAUqmHCW6pvL
8Zw2yXuSEpTNof6G+OdTrYfBi9zpZ5Zvb9QTA4F2ILE8Kz0Vrt5yLXLn8LoT
Mlqf9+MHRmamMQwKRf632271bRolDiWV2PugbIEYwi36oj9n9derYLP7Z1A8
K0JiEWVPNst4uMsvrGhdf8YNjddA9QgZWV3sNYrdztec4MCN5lm2TkEolkjA
O8fL6xs3jZ/LNEC2YsHa/w++i75XEo7gG9/Su0OHkgQYd1xY7jt5utgpp16d
F5ozgMOUpArEl+Z3PeZlXoRsXVNfHO/iv9tnIFmxgIXChFRe08MNhQ7Fy1kb
aTRWoDZwAatxuh+o3CCC3D4pCgoo3OaXi6nlmqQYEWaUKNasb8llv0riFMS+
UPub4uC6WKoVPRvBoWxiShqq3L2+X8RxQtIYUB9Xfa6+NA6O/0aXSbhCq9R7
g9MCxSsNg5mzMZybniUJicC+ANZxxdY2EIPX9YFP8uDm1LnYI41IgHRXG6fl
aUD+8fxneqBp7byluCOjUEXetqp30rm5gq0In9RBOWrkxGgyP0nzznvcyh7X
7imguFeU7kt2Txm6npU+YSL3+kal7OKh1c1aNmaXfyJpItw4iM9F1bXta+YF
vhxiOXhbvhY55V3KcXFwTttmOn+1wuQFsqgJrBF4WiRyiiimPpB9cGrX+4WM
T6zQDkVyooU48KDD/HoUcA8JqnpVbplkyzsD1MtJPnoHl6IwHxvW7yDxQKLK
jFfBB2/Bx+74owaQGnE220b9BqjtPyjAK49sBIA8jtE8/rqkLIb4P2+p5ESu
iHOJItpfbSKF9ZeXjSbIygxyrXoWP2dh4/WLnfTtwMtCuVlmcvSsrZB3tQxE
scGkDBwqvzprs1p5EHsxu4WLCL2dV2EGmzea+O4kgSxDL6qDKStHPCvYQEeK
z5CYeNdU0BNeUG6y2gV3SxYSaPfVTI4rtBW50P/X0zMwGsrstZ1TmWHIIalY
/6OLUy4L5ZJKqxr2XFaao2U82AjdL1Z/lIFC0JK6mThaG1LesSf0APwAUWC/
GsrGMCC5vH7tk2O5A3dEXH4D86d6fvRnGswDgE1BlNw47MkPdCyNAEUWbW0/
LxIqKCLPcaGTUGISSwFMW6FkvE7tTd/fsMQnTNdmIHHV/5OiWPICWW0L9MfP
FVEMkRD6e9vlsI+GTbsCMa8MDAWkyu3i38u4Hl+Jz1zpPA/bgOBO2ld0P5lP
dbdlL3SqQOwZ/sau7bORaaq0IsTnrjQLWzZG9Uw723P3/eZwU3PRfrYCYcnH
/5WS6PtfwKxoeW3i9CtkSJSvHCqYefwYjhX3hthWSPveVUN5djrxn7qKh3KH
ygIJr9V7khLXsoWZKLZJe5f/7WjJRV+rUxD9kStyQ5ITNxPZbcq74aENmYTv
w1mfVH5tC7LjSyvJXzlVZ4HR7MCqP+KzyhB01sUufANhDAK2fusZjFEAtdXG
a7jjt1nqHyfznyAT4Fs7wv/M2DMpwtAn10g9QwJTP/mFF8OWw+0dWzfE6Rq5
/0tcvzCglOKXCoR/GowOalnELPXvn7qqfwUz4g4nWzw0uZPyTSWgsGs1L2w4
2J/mc85Gu3QtLCWp6UKbFTda66QWV1CIX3rWt5LzwoGEpUsvqzJMmNQk5ds1
51O+LUT7+8v9M+klvucn3DeqBBTVq0q5RMhUAI5nO1A4KwM4oWpdrMx1mYmo
3245AhxO613fpbht2jA78KQiO/bcKZ5uV76+ipkuFrpRwsQ/Jv3DMiMizX96
piZv6y2piQGZOV63PgCA9b0MnKwlouVMq5KpmDTkeNV/Q6GLLZtVRpA4saOm
2TUrX3SATNPNC10YH6/pMwCW0hXGXeXBhsYA6BpRD2GFbwlOtUZw8TCH9umt
JWk4MzohQkN3D/qzNNy7jzzpOD+i+Bi1ECn4IAitBDn+WLIytjkxxZoakvAb
qLDBojK+hVIqOzVY5T4k/XyGXTLQEN+cse3SqfypRIjgzGZxmvyNGqgnmHDO
oaG/6kQbtTUZyoyKab5IoEtfEagSG32+eVIpg+9uiINt2JHzOEIg/OUYYjAE
hmcFsZGHKWuCNv+VPMX37OLk1DxzLNiWnNGonYm/v6YO/QxuM3i/Lxk0xZIW
NIcPplYk+qOuXpoifl6uA5iOCRrk6qjIpes7OeJUopWVAc1wf9Dy9K9sJF6y
Orz5N32TFc6IFvdNVSLR4LNY3Gq5BZOhtff2GOXhV6GgUjmw4JPzQniwkkQg
X4I8yS5PEQ9vxfG0SAJzLdETa4UE32eqmEpbN9AuRGx1a4Zm7K4CeWqbJ+eC
TDe9OgzoEmBZUyAXGEQgqe98RNVPHGAOk186DwpRipdYoIjIDCG3Tu7K9xWB
4YcehglbiV3OwRq0bq/DSnUS0v3SPwbBhuO127GAVhGCgQSoAMg4Uc9mI1Gy
DMniL761OlmrfxNJ6C0ZAIMKym5bChwU35qUjekPAobxpjjvacgN6n1dWHfC
G+iLcle/j/TBuIkV7sGcvKoDo877FtDIkrKBMMLns521bpPGf2xH3muSer0/
U6eyJplwZ3tBqtheYCvmYQNecY7Rh8mkc+G0pLh+sUL4qSFfDec5npjQ7bWB
g/5sEI9PtjFj1SSUTT3Ygs7P45maJ2fWRk7lupUtMU9pDGjWzmVWm+I+oK6T
QHlacJVcgJ9ZrQhBKzyNIf96yeVWHKwsv4SuzBvMVS71FlLq1uyZtSor3uHe
mUweumcOMmqqUJocUykKdrXWA7tYbU/vRiJgGoADdzOP93/it+DH+taIbSu5
4fvtuE69u1LSfbmEvHH/BzMJ0KZo4wuTt5UQPDoRsrQ9rXC6mFTJDZ8JSyPC
PuC1CF7ygFzjNQHEOyp+IK3n5ho4WERSG2ylO1+tLSdk/AJNIaqIM5X2yMu6
VYWRTYjMYvP3tnlZDgH2nT5/GOA3GJ3EpLC5axbvTZ1YBXxCyItCW5S86JAd
S41gA3vLnqhUWSswuIeAPIaAv0avdGJZe+Gm3ggPKhLGIotq5486BN1kGnP/
LwqpNsXz/8KolwULRDKrhlqYABtqWGMmKthfWzanZOpIXQuRHDN8RH2gEHjG
6GH4NIYFXgoiGRYXxo+f/ESU8NKR+xC+gBqvimBtb0071k+UCOQHAp7j4B9s
o6m7l2e1PSV/SuRfP1+fibCZ81d2sCybDF56KcRAvTuTzuZpNlTyJPN/+l7j
Fjmwa3qr0aBv/SeG3zlpyJL1CggakUJ4LiJQ1HgR7T47dulUgsbdKluvR5Zz
NexKPLRyGJmd0z9gqQx7ka94lj8FAeCu/Fh21yUblR5Ma4LtuvRjm7YShZFo
DwMX64kF51reEFz0aBBbpAwpAQ+5SA9c1UywV7IxoP64Xq9p+U73OeJwPFES
LN4nq8A/X5EhjdgG8OB18/U0/DS1ruGEze9LnNBreBZAzgsu8mU0nXX1wE8t
FWda36Ld+tB0jhc5VzuM7lO8lvquH2JChsZlBAfEdEJ73rcGW/qkr7xZNSeG
gpQs0DWnAh1BuenBRccrK0NzzH6ZUYuBZOARFtJCukkf703h754Fk5kH6yAG
FT3WhTbBK4ZtrnLTZJprhPnbbnyGJCPPCZ2gKIcZLJMY8c2PVi7AJKdqcZO6
UHrhNFg+pcms29BRp9lRGL6FjnyBSVrYfXA5nO9X/FiTD5gVlej9HMMsleLa
L4tDHHW4ffBFvQzpsOYYQV53CNqGtR22XU3osQI+2fFsjIauw9THXqW/0Hld
UG3t9e95OpQ1fvkT9XCKrz59Y/VQN+C4rteSnR9/A85oQRoX7Tv7dmBtUrIm
j+5+Y7KYOMqtiC3r9sulFj3LvywmLtNZPHPF2B8+S/pGKnpC8D27E39Nsi4v
L4CAQ1VrK1KTqykn9F6mAS/7kaJBuVsJmed0TuplWQz0Y6nWzbfzrzqSCWaP
JVIkTl2MOYrswgyv7K7avKmUOKbpfUXL3TECmlWlzReL1JQknW8EHNRFgZgh
G8z8eZDu8Shw4sjB3ZoCb0kLD16yfi3fEbBqC++xjZZSsQkfrIvk4bh5BSd4
LArQ4mvHrMSj2sMH1EMiS6YkwcAwHcfHuLLo2uHsbb6Fh6YW18hRmKUFA1FW
j9SEQ7SEly4i7yXb5JyrkJlZ+hg44BP0N8jfjiNx1Mro4xUEQQgMybi4TFa7
GJLZ+oAY8Jd6LFxz1twVjYltOOvbezBTgt1zXXuisToDjodk0JfPa9E1Zplg
NQ2+6AIdil9aXJ3s0IbTTgzfEAt/eDTFv0adJeSDREyCCbBjlNdPUi7GSoSg
aItReosM2LCb4aeE5GkX/dKBcfEgZGAyOo/fauQ12sQZfrWKTMgo8Glf83dM
rDLIbD82tsTpxYnhZsnIZOGV97AIsaP+x1ck2fxdfRmbpL20fJtXWlt5LYz9
9odWol/Xdu4QTVAUexm13m4iliHEfx2RudJiDTgQ6ED34VhknjhKjZd1Fvu+
NJSBci9p9vT5cmU7rA5GDFFatn+KbAS0azcA/j9qdlqLVGWV2bnDHIc5F2Rl
fUmzGxIhhYCYtEMWI+99qGco6gkWuYAIXc/Yu0Fzz3T1UXnwmbVAnkgd80fY
ISd3YPpL7Ll8/9yV/rgmlNA7yBZDWJmdGSRrrKcRKEsLrempI4BwDtFURRdT
Fh4eU5O0u4MTliEqhMH9ih7J0aHbc5INo0G6nf2hWALYENd5RifApRWN4dZS
GNUC4QMOyL2+3R61ESQUP6uItfcNVMeqpbnLD+xu4psRLWUqGmnGaPrYeW3K
AOWpYJBg3PXg0yF2nF/Id8Q3rjMN73cjKVb1WlNkkXCoF5S7rAMD5gk6rR7r
uZrpERZb2JpxDm+tikQfsySu/1ijiN8Pw6uBvf1osLPJrN3wbKk4vuLamcKd
p6h+CdQjDgFaLz5y/A27PciEHh3ayTZGaMWesl0fUaFkr+dL2zh8qQJ2ym1z
F6n2KPuX6TWJBngeaLPdcbmyL+dYpYx8JwwcqEALw2ka3RBmYRlTGylosBR2
Ys7h8B4UDpR5MdYY0QPSvNShSWrwsZg9nmsrHS+wxBKLetuRANvaeesmLIBm
VV6f9IhWykK6WMj8ltz2TB7toswXU/APtrxs/mykOmVerDTwgq2gzw1L+UtB
E9ck9sfdT8sb+/28I+Gzp/lRISVIqHEM4rCacXcp3Kb4X8n7rLvzmrs/5lKP
JrahF2H/Kvg01Nx5xP2mXiErxZ18NAnpulg/Epf/IRkvSfhFjaPk4L6xAw5Z
pDLTcTWDt4ArtEUkv4DhQ7Kf69YQb7rK1TCKn8nUDG7257KnvKnPPn/dCVAb
P1+KftupHvs847Tu/z2A6E4i6wyRzeDHAq0DOvu3DGIPH++bSmSaHMVhOvsS
OvE6lNHCWMeLTz++NeTws4sqvTzTy4j+i4zjMV92sYsd7HkYk8iJPJktHRlV
e5914Z4wdBmMZyY3fcpb3C835Xr7GHCfWbQ01GTtjXkB/OlAIMnQEsdXo3Yk
g+j1mUv4DvjvWNhmezunRBv828/Crzeg6bHFkjMyHRo9iht4MkRJWC/Yddhy
e5Pr8jjDsx2vP05e5fCYAHK+emo6hH7P4EN/cAd3sylJqvil+Ks9WV4Ut1cG
Ae9OmMzpxXj5AlfqOuTIcrsEBN+BMVWoB5QSJcIQrBy9ILrtzCEryrNEIaTl
7d8p7VgtORx3nT6t7nm8+f2gjvq2YZ7ifvlFG1KaHkmszWU/tFpK+e5WSCnA
P5dXkQE7/XMv+b7EN4veFsyk+XztW0hR7Gu5RDLx4GAAH95HPSTRP0QORydk
ypKbkqD6P9TxCccKrnlZnBm8tOzSxHn0sw7vTfqvz86MK3znmQyTKMdU1kFK
WeDlmIFUJamq8p+3MRfJ4NyBdgJk8DRbArht2hpAboNndLnPNliuY30lMIVo
Qki7gq+OlHQPaAS79Ex7hB1O0qaQ56/BdywALkO/aP8Xhdmay7XOM2dd6k0E
sxlJMb5N9EHw7bLgGDfbJLuR7ZlSm+E2tvzny73k4yuqw+VjpANZThKymDmB
p7IRC0QZ43/wcvwjqgIxV92aG52z8lGIYRn3XiA17mtBylKeK+/uYFsb1Fuw
ECEJnPpjwJeymJ+Nb+hVB2fsACW5zoXDAMTSVGCnmS1UvK8GgQqTI3Re9G6A
H7EA/379nazeYKUR4Ji7voVr5cUb/Sxi8YpjRrWHK+N6jm0phk3072/OHixQ
fngAK0q3iG+5a2amcEhr3rbFXnFss/BL9E9hOzZt8Yrw4+Rm8qj7W/xNdabY
3XtlZ026qxVE27DXdNARsTEhbGI6h0WYupbgnLofZka+awvMV/CbLybNZrg5
b/H4lN7yJYeRd52DZFxv5xCvM8b0FyR4q+Zco7owpLTcAzWVPKOpZeXq7ovK
RcrPAlU1UmrZsBdXwGI4nanbm7X++VDdqxRTWH6DHI9Y1TqX5noKpT1UvvpU
ZHPpLFEnbgjzL8RlXRAf5ObC40zKRlgwXHH1wO1mDx7q3+9S4/4L/eET80ge
DKV+27mvu4UsYDeyEUXs5RzVCoZ9G0Krn8iGm6fj5Rov9ZBhm1KawcU7JggE
Rvpco/c/HUwQK4wDCstL0t2RlpC1TNEufqvefnHOfkZkRqoauxvQraBZYBJ7
gxl/7X7hWxoXEVt7YlbyKpv/53wV88/XN3WtuFbvcu8chtZN5svc0aKMXVNA
yBKOmebnB31GOjjA9qu25H87TdQRe2eZp7U8mQrZyeMGvX4RBPC0d+QdORGD
ZONu5MmWUYUUqD86EE+exLXHZssUQkLziv/gztlut5fOR+/SjfyNQbScBSup
l0WRWbhV/tm0bPeeSSVVxyXaSJb5/AsYYa3jjzg0KDSF1rP//j/9TTxmnqzO
IzUHSM+SK5WISJvgFOiel8/Dr2WvDEpfnD1VZR9TrejHsKdVKKpuQNV2TgFp
cSXHzgvfuFKV9Cfd66bw1+YO6oTkKSbDgBE92udru+SCZkT2zyEPApb12MGU
krwv6k15gQk2HrVxphBOQ1+MVzbQp63/4GOQ3oY/4R1+M60uYIApYSBpCmEK
yV87ru5vErT/B6wd7ACLb1tTebat238ubvFohdDfSumqt5HujfcTTEHqVwNd
Xy7zyA4N5gWWcAWR5hJnW9LaGCHX+Il0OYA6r+kxXiaWpvFsvPI5JDsivgr1
+uhnOA0+XYAy60usU5GOvGfflE7Yqkdx4RmX/bDtde56559IAxZetEiLKq6s
RNJh6+6UdeqZu0Ll1poigtmwDotYx/jeLwrL5cviNax4u42NC5eYlu6osz2U
vlYgi2hOUWg+YtoTI84KN0zIOubz0FKNseJ3V5nvQ8oa/p02VZCNIPWkkgXT
xfzEagZhnBla+DHIWPDUPFM08xk2bK0jgXO/YpyjOdmBxGntJ5FUyUqlJusF
mTWJFT7f1rm1S4X2/u1CMNU9fmXTMm3N6dHa5Z+r2zc1aWx9c3fIpyASj1TH
pcyGv3c25pAQJ+2Lf9C+sGAq4uL6Orxyt6zZfTiT+lRYgF5xO9LkgY2qCe+R
C21P0ZUsYzmy2vHqXouK5uybQKOPsI3ePLbi7tV8c6moGw1stFTDKnngWvBG
EWN3SDGF7YUFzEHtXAGBZdBBWVNXpmDS2ZyovFT1GigUPmrNBSRwKFUgR3cH
ErTjgItILog2GRTJLGB0rjEep5LnYbx/Dcld+GxKtv9sgy3f43w8hv3/JEoW
GqrgNW7GqUhFOLxp/EJpg9bU8qvZM8RnZh0ojGfymIsmTngV/mkwCqujkmf2
psRpvdtbjk4lCyKNkSR3VeuWm70k3VqoyE+rJ4MdfzuiSIaidZQahGHGLA0H
KDi9C50emFmJWDdIbd3xdru2Mr6NbKBez1aHVKs2LIu+nScciaKqfrLxhQlU
JgaDAsSVEvaILBjbhA1Kfdi2szRfk5k2FMtHGiaHumZtDZN4a08IL/zWrnI/
F3FJcmE7Y2gQGTLOnFsw78/eaySuZAQhp+8Tfg0FJ6DVFgTc3B2Lyq1f/lQS
U7gf37ssTTscTh3OB2ZFJiu53VE3cqEVDU3M55ffwm96bkt+StqlJrVAcaKf
h8Oe5geO5tzuESEWSU4q+Fz/yBU1RxEYmJ3LRDFpm095AFnEJFgHVM4FAXhN
j6CpOcW/ItY/pchdbNd1MzvDYZm9TDlyd60IgZkCISxOkRuil/YNH+1nhC7+
zu1AdQU7lAmweJjdFvZLT0zNWKTX5pfOjYXrk8/cdPyDVCDfzcR65SkYsZd7
mIYy9BwEYoS1ciPDNwDPLIrbCrbob6WgjTLKIByETnc5zGaK3dXYYJcivS60
6wetw9XJcp3cT+YSQAw9ytDd7FYG1wQSDyU+u6frsF1hEdnnW0CXH7drkLu6
FPbksDHCjou23Rssc5SKia5KVvCp+ilQQ8EHDwF2MdnxIQvfdJQqh6A8mvv0
wkiPw6m9AP/ngbUk4J7hQiTcezXzFQmhyhQzCFduU8oVMiEjsGOL8Ew3gyxF
fx1yByVXDWZwz7bBEhWQKEEMYhHYdHKP6w5L9YlssRhBurnzKWjy3+G7orS0
+QwbeurTQuoHGI2rxAu2BVG+wj30Az72hLu4lcbqCHd/h57P0VbJNZsnfxi/
0Bu9QKcG+RsFPmR3YvnjyNYC2L300K+YjWFno56W5qHxv4ag0X3hCFH89RkY
8iqF72oMsYFTDVInaep71ZD0Ac6Pjhv97ILIlZOhchSWj1XMWtx3SoO7NPc6
O4IgO8j+uPBsEOSMnRruAh847o6TEtVO0jfIKHUmQAHx5ONz5gIonm7ZAPqu
JZTeNNtAoW2xv2BgoXVy10uQFKJxNzCjeard/g5D8cPi8oyXqWhYEuPhOnOq
7h9MXGO3nt5omp6sRoVohJc9YpK1JyloN8tjjuKfCEk9wRfBpPyEaqD7eFnS
OyQGLMi+eL3pAqryICj6R1I+v16277v2qBhmtN00MIQeK9Fryn/PBrWX7RoW
qCXJq3VAdbayf8dG78eORSUrIoZ+bqVPjdmUxBeYsmX5iV/7JpCXHHXnkLQW
vdmtKdoD0mDDAX9ADHu+hRLnjV2fCaN9kv4NjGYYBctNPaNokKR/pNKVLDnH
G1zjDn2i/5Uu5teMBqN5wz41IJT3aCSEDjEia+rnKyYMsyKPX5Bx7RM9x3F2
pzU8pKuTc1ayU3xqtzHHpyVSDwZMp8hiGCGgC6RUGexyE9n3DP0RcLNECtM1
n7WB7mKJkLQEpOK/0hyYq0stu4roDCuAK1ss2SekFplvDNfMy1W2cpmnwtJB
YPKmQAzoyZPp6GEPJcHxUXgDUK4Vf4P2KWSsAooC8plMSUqJBwNHBxhdGyK3
SedWe1o1quwzyBJfl/KW534Ev2fjHOLNZDBlJuWR7J5Mp6Ahf6YGXAH5/fHv
jP9/5ziaMQMnVS62uWnf4ZpiUaCHXqJ5B5tLfYAb3xj+4TXuxRrLXPAjc1IX
yhbVEZUHOl5h9xebKqPo0IMdOeIQe7PYhC4GHx5ZLO0wjPEdr38rxNq85iRh
QzHFoPng51p9eXYWHsO4qkiT27+XuY9ruEbglsBsjyDAXBzVDWXiep3yd9v4
I7ommDf5JwehzS3xxmkfEk6aANR2Ocqje9yduokaYMWgUkW5zhlHulikgPa3
bAC6NAC/+WpgDhhtXE5c2kwgifsQY/4QIkSjYMoR7d9JZ5s59LSgCLYXoCse
l6Wdn9KnowC/Ct9ZUl4hrQ5bqWRmh8t8PFyu2aydGR5NuIxQdTHQbiZ5TIHO
TbcDnik2135A/Uu/6NkFzxWvhmJXA3x/xO351KNcEixDqapOGCLF7UyB7sU9
RNw/JHC8nYSG2AvQ4NdJxFBoPbP+AVdwcIQ9kUTUUqwv8IGJPSNRccaQjqFS
pkpDaiMREF87yzTaOR851ZT/e8imIZgJES0gi6N1MFgGzfdFrvX2kee4Ro+g
+//RfjWNiBhHpuhs69r/MDFnFkYPGms5uhheuaBZOA3TELj8eWbIUKIJVFfH
exDFZUMHR/QiAFtza3+2rO6nKK2BdEElwF2nIycNCuuCN8FRZcqPqZZuAxa2
nNgIo97uAq/sLNsrpN+4/O8YsSNh1YkH9GxoHpibhmMC3zYAAIP8v9YmunjS
Bw6VRzF1GDoO0SI2U6j5RP24kcfj7MTF/2TnEsrAgQBybZN7XzrRo7CwD6Vu
YmsY7cs7luDwCfe71zcgXjKvSX+7mFQ09Qck/B3rnsXcqeSXo2RuII8sHyjs
TMztigMmFhJOWLjr2k6PCwigmCwY29RWRZocwNLRkyik51AM8kn9DqHFe3rl
gwZvth5qFLNeG8zKD5ersK9BpDkBq2QgrdGn0qN9b4iAFnecLlpIvw/8/vS2
VOTHplJE9YDLRI5zfcM6XxHM2RER0F92dHSu97hIMAOcqig/f8TbzkSQVdtm
yUuZw967Xiyi04YFsw428xLK+4YUTl0Vil6MOYYk6nDNWpcpXEYNXLCicYpa
xDAIKJqdgOxHPGNgIqp1ZuaYtJywwr/4wWqbRDbwR6MfZP9DHp2/R0ODADvS
8/1OuSMhG8oPQWtTeK4jr80oygsp2vZH3fmih+R+hn6L188DvTXUV3HibfKO
yLlQo8UBo+UF7CMAKrHdrgEiePskON8DFjvmXnqCQB8s2vEcwv2v0y998be5
2zT5iVc2dYiDRDoCCBvSWh9uZfiAkGbcL6reNrd4ImDojfDuUf+2bqhXm+BJ
YEAvS2WX4FXQIt2qAseou7ZJYU7lOexgagUVStj4AF+TMOoXw58yVecp6TJf
O7dHTYeu4vwtHRscnCAW7Gkf4zj5Q+I7FQ8xXju/aeb8cHmLPwQu6brhSv42
QXm9ZmcDkEyXeeR7G/mCLAriwHHl4roTXLyDKaA9/KmbN0m5lbMquoJbmPBb
O8V0Q6tivRM4l0Y/J4g9adN+UCe7ENKOevOKOtFkoDwWRKjy/E9nkRJYmBME
ifPyWxYRz1M8kcQsGcuGPtbacYNZqIF7g+MfD4aeczoMTLQogsVJw2bQkXwX
MHgHJ4T4S8ReOGum5Jo1VPrmus40dsZHw1Cxb4NoTkXd44GO7w/Vyw1BE9VS
X2Q8BGBu7+aTgfgKVDsrNYq606KtKLtrGb8S+desXhWXeSc08RKbqL8lATXW
jnCDerhWACVOZC5U2w29gQxlL2QkO2mfVksz7w0fhwCrkjJLx/IZZmMbsAaS
2uGUJAAIi4IX/LJrkwhRbyFA4d1Qp1G4heiT3ejTFJmH9PlWiTLNtuD3TZHU
foVR47HTgC1FfYiqWAEdHsC0ecafsK1pIeHnB4q8BfTNRYew9OJ8B7g39zqW
wJmQvhG7hBlkzb9/iNzax5K+2pNEOae5EcYIM/BmSrrLvqJFqhLBdaJL13ym
0zluRs1amyygGmLsvbkTDFRSaFHv6LoIgloFz3mck6TLNJaKdNPl/1IXhDJx
Kpf2N1+/Z35zK5Sb/DSL5ZNjmHax3lPYhn+Ac//WVSclISOfVgabTkJRlsAW
8b82IXvj80R9oImlnol7j+Qm3j6byZaEGsLVIKlFkkH7ZVIJi0te4JwYTBxN
/jjyYY9SRRC5wbE1Aq8AgIFMBTVEWNZPmwwAfXKjIrWt+z8i8jPNQU4UqAy6
h2TnX8NR3Y1BUuYnleXvXl3qo0Qh6HXlO4P5JDb+n18MxcAjxu5Y/GQAaNto
eWVkmeQacloFEnjyF03CDfjbRfK1Nz2FrltqLnKa7BCk3p9I5UTUM0GweqIj
wnPn5gN2SEcOHvhqF4szC1gOue6xZaZWee9u9uO0LOywDdGW0zK5/4wNbTgv
py5ZT6+dA2UqEh8SoSiFerAw9jl6BF5Z9uoBEfm4GDFxfk0z4VEU1np5TrJN
nx4y+BedS5eaOToTmFMVBQkwXk3tlvNunpTl2qzcYldgEW3QhfwqerOW0uLa
iZPnJbq3nXvpVSY8tBcEwlUj3LSpnUyH32HCiwt7ZHrePFeseq5vq0XBw7wm
oULeI5Y7qm1MUKsnN7RKnLN7rk3aEhShqe2u53n9216C7alUlx4ZFtGgXNP5
b4KkjjJiT+lJUi/LrqHsNZVsnu9KJnf7W1CTDCRh2raupBRQlZ6g5VVxefL0
zwwIu4HzG2Bl0Msa7koCGuYpQUEwo18x9O7OfcC4qCp7B4fW4E8Vb721bhEZ
KZj9DyhphaRVZbNlH4oT9vLY4El7Q46xNCjRuAg2xniP0ihXPpyoyYd6rM/j
Pz3R6L+nDHFpTOeeVjX7iPjANu1JgfynjlsI/NFDs3nU9Bm0g1nJRKrshgPQ
2kxqRU8CEK+QzHMuCrSfQsb59ViNJROIYpFr8PgDaG4EfGLwdK6qrVVmWIMK
TAK/lrwQHBthv4D8j7uZYRNLLNZ45wdq1vzMXuGpF7EUQbOQfsswql20mBXf
0tL2JwXWuc1lst04Y391uDJpd25U02QbiKc0M/GClmrVE5+z4e1+IDzAeF+a
7pKKQzpQmLU55Ia1piQlq3DyMKFqOhROI2jGBxjBvXFRPEauK6HhVRYu1qgX
ROqQ0Dhsh2MOQZ0OcLBTGpsmZwD++sja6LkXInFzTVNYoUjgF6D5GICdewo+
gbL4vmM3xxUpbC8ixS/NNsReAcUxcbib599kOB1IY2axaVNybeaeOUs78Nfd
+BOZPfmJKQ0KUsqMK2ZtprN7SS9dmEvIEU6+73A1zDtVzQ0svUPVHKX7GM1R
PViyyaaHF/34I1xJ/RqvTSdqQJIxMcMwA6/FGXMlyzGQl518eGvDJ7mzE3yJ
utufdYJvklyBlj0rZFqRlEdhWXGjlGT22nA+Ny65Rmea63GPH/qLB9Y0nv2c
oPzJJ+dFGKWubxeEKxekM9NqN37CZAQGy3i6QRBZkzP1e/HqQDhwpYH/wvtQ
KDqppWulBu3iLlgM7aiIXgGR4JHmhEQ65tg7PP4LlNxzFBKLg6Oe9c6Nsreo
ddBZoHmp6kjcGSkRswpAZJAXmIFcUDvqD6OCQv05s1QtcfUDkFwN20Sjj62X
Gy9oiWnU9/tDgz0QpD/yTm8UDDBS8Z4KsCkShh8mtSl4wKAWQNsdWr/VXaR3
g6vp8OzFIoh/ao5x1EkqKhiWtHce4FcJmBQT/h3zzEwCYlZ3N3OaV+XsnVk2
l0oBiZ/dE1QJOEY3pD+dYzkFr7Z7Kdo+bO305lSj9vmCK7Lh1Lgj94/vye4h
oOAFYaNME09mTgAixCwOls+8noeWTfV4oJ91j29hsV5bOW6Pz+F/otxoRfR5
GTJCiXks1Fe3Z7CAx0bOM2yFD6GWpPN359RR46yxGOAtcjzE/ZMF13PtaNxI
wby0Akv8x6FOgS8d2bjLBXNjRo2hDMUllbsCmJAGiXtoMf2zQXXSBDxuu4Va
N2ukDgjprQyE2udfhtCoUDQqrLqaLZDwEKAbk5ukYTaNIu6BDaRegwyOo73C
olJjjChnQxUG6yG0C20SZxYu4wuHAVg/wZAagzQyh3DogxSYFgnAJhLyf/to
6xcUQ3P7QEYfiXn/Lru2ZjAF2KNcBplhBKP+sToYc0QI1l4PK6gYHqDHGKPS
nosqBXJOU7hZJKx7wTqjTs1i0PPRFEQObXUR/Bxlx0JTZPneyFpqIWSU4qAa
fHa63TDTHYrdw2Ha+H4o6RfNZTZEGazOJ8auWYbZteGiciMTWDzwUt1vmEcg
fMNeM73u9dlFzzOtTivdd7hiiZpEw++UQih1BIwcnhUou4hIbieQvsbCmeu1
hLkdxO2OLuHKuy3AHC2N+vONmprf6cm+G+Fp0m01uHdBJmRyF13rHxj20JhS
k22O1zchBcJI/rgNkAGO05b6AcqFrgitLqkT4yqDtBNAcSUBGIgWV+691njB
1CpH29CqbFtXdwmOCHxzk+sKOKmURtuN4jvF8oHu7VFjIrfAfI10vkD3bs2U
hKpALEzwSj0VHKp2dqchSu49Tt6qVLq//o0L7qBB11DAr4iDFaQe4pStuS7A
vLtGeJ07+1QO82/8Y/mUbqjzktZbTGbnEsLSX2sXDeXqGukyhiSg/SvqpgUc
xAiSa//XHenW45z+lAR65LZ7hxmb0Lq0SCLSbkrDvYj6Vy9MPyK/xB+fx2ED
MrYE2h0JxR8sgfVpXG/3EXewPo5F+0Gf2JAT08gZXUq1ZgU7NtL1P6AdOGRU
udjlmLLf3fWkTe6r1LkTIIiJWFHsXzRoYkk3YeojWEHGhIUp1ob0h/mqB0Ji
7WpDlMKBi57vlOp/lOCrwus+gUZ1BUC9ypWruiWiCA3tkX3ouO30F4pmqI1k
1ozAZkceXyrMX4LEsuVMy/UX4oEM3xVd9rtaXEDZNiwxNTgVbDZbFgrcxMqT
RnLel4VU9TfHSVsRrGekCIDFn9cLQfCHPtSJFJC2SBiTg4iBVXVjcICJeHJ0
8K/TNd4p0iZ+8lX/gb/f/t0GN/yw42JOwx9yuox2MHSWgzeqzQnCXMb3H34G
968vqu9CZPcQZeqvwh688K8TW92jaYUfhaElWHgp2NjTXLW7BamzkI5moFQT
Gc8B0WXNhSxzbDG3adDar5yqjZ+Qic5JG34BRiaxMpovxy0UfnFyZi6iXUu/
TzWBR/OqUYuFleKWgIqWqvEhI2WfhfXV32aywKk2vPyVvYUi18FKzd+XiI/7
olKtLRcuZr/iriF8kcDf7PtbZY4QtmZ2lOtUWZXBrlrxfOV7DntNlqMHZfPb
sj2GDXVZZXkfckMMgqhEn56y6+fn20UvPYmvPEGd7J/NFi7T8AB5EWer5RJ2
B3ZR6NWASjD/QjHUUZ5dac8fezC5cKOIAKsd7ETFrH1WxwyR6PRRKqBbAzkv
R5lGQ3IJd6av9nQEvaGxCz0v3r+R71/fI5JvY986II6Nl/2OKaot/fhL3XUd
bSzvu+gCL1YguBkCbX6mq+PtvPb7jYtlqikTE6/mPMKYE8X4PvUr5cgwh7o3
Vq28HIBRXBrJ/vD8znrZnJeBf/sxEbjimN0MnGF2GTeEbREdts1ZTE0VGP+u
3IPXsYso9s03EA8wrP4ZQt/NvuuQHrEZ72cjkbw46sknvShHGNQ0ps8OXacT
8nI3OAGz+LPC+eLlf3fH51CI2v56jBEabkkLS5mEqi5q4XpPfCW48rXYU5wv
j0svCc+Dj+oegK19niQC1raT71f8nkCGhxE2H/iTb3KUnJIEM6rvnfASNH7j
9BrNfz/gJ4WYJhvNsahCigfrQ0EEsn5MfpYElmr3W15nvNRrljHQvwlGGQ/q
iTK2B2SCBDa0XOyJ4FPQBEMY8roZdLSDU9MRyPXS6Kau5clQh+JgtBTHkMEc
NiWXqbskBQqmflimqj5ImI/kEdj/8+cTOH4qbWlzQb7GmCEmyYixG2As/NGS
iFUBmVQF6Mgxr/nxtQhp4eTBdtocE0YAbdzykPZaKNuhqVE9aO5j0wgZ/OmL
KPNWBSWQLy0yQbJFf8M1G7ceVT45Cyv/LP3Mh7lL7S7T5O8psKnqG+UJtlW3
VS+70M4XZFdwtyTCPxnFhsNAAQZvqC1J7D8qpmtwQwXF5nVZy2aSAu4jaWzv
oGl5ztaUG+cvj2Yy5MvUA6KPJuWz09mMrvWCO9otv/aNNhZ/V4Q85MZXq1PE
p+ncZx98HWj+7Tx3m/tduM1TOGmiso9Qwf9K0W6+tDLDvok8ZFNndrE1R6YB
40tIZ6JEuvFhV18ijATBIv5+67w5zvH3w1tMTSVDilqETJ+HgAkVo6Kvq03I
FkjyqcI5bjbiQLF83uoLFrsVO8xXXI5Ac6sBk7IyRNn253i8iGOmsSwu7zHh
0/RjT2sTZ6xV908WUBVMSie9zXgi0tt8xjXV/mONnzRcgzGIAXwocxDMB9LI
zpxwR38+T2XZEqerWalLIQrp5Cd5eLhNqnn7i9vG6Xo/byGvKJOLnDCErQZp
3oOlCPdCMv2tEHyeGZF28w0aQ9JytnSD5lwHgx3WwSAgFBG4NymgjfD1+A4w
EZTf1jJa5O0NO9WSfh5rLRk2deZgWu3ZTFKn5LMSv/FsxpwkTK70fei2dg4O
fmN8in1OvXl8Bn9ffYSVACuO+aMPmdQdRGTmFctSdp73o9l1EgiFhB16hwXx
Z9qNO1VVY/uXx8V8GTtXOsd9Re7bUuWlfwb+npfYDdjgTDYnaDaJOBr+v+/k
aBRkYrLB1T1HHnUoy8qfbPpyNCdO+nAFQJrlHfv7HbMcpp/ejStdkcegQ1nq
KOgtnMSj/BwJeK6vtZ/cCFuhLfVxrETUctZsIYGopft/V1ZH+63KfcyJ9cLb
c5DxcA9CLKLMZa7OqJFqS6dmPUgcaYAHKlRbCyZaWmthfU5m/MXYxMRnXJXP
T5YeD1fo/A+bVgtfQ/ePkPUar69HsN3t9EcYX9xVq6H9wcngbGS4GuLGG22K
RjjUtAOuSBJPX4qlVw8z3uqvS8IEaF5gKDwd/w8OwGb4q1ZqBVNDpu9tggMa
Yvx5VL7IA/G82BkEoFDMhar5+ZIELaJSC8wM05/wQ/gmpQ2ZodAT8IzbYzAF
btGYh67UB5cD/GnjS5uqHXYMBI2mwnp7E3A5IlzrlZTTUFhbSlY2ZYAO8s8k
I8ruav+rxAdYklsqdzglC0TKdSdQtpNh4ZcXuHM0i56MV3CUM6AuxM5oZlHi
CB3zvhXnIHDypIH0iqCd5DsorXxpXRtuGhkIP0j+5iF8tJa6eY17bbR1QNok
5enBVdDveSXA+CuPKOMz8OEQxuTca+K7djFw4rZS4gBam9i2wlw0WcVezIwU
Ik7MzhQSbq2R8Khvymr8wX90MsYNvD2aj5ppZfqkOAuHK94otyaGJDXDp1kg
KSt1TlXVM3Qqmpk29UDo/Ih0PDfGnSCg0EbDBgnTOSEJ1tdy7NubBQB1uIca
r453w3v7uZSmAyWcdavwJGSWLIgFGNNjZg0MFMw36Gd2WWbHRLos00mq27uY
94tyDjMP0aodNjZm/grQlvahH81kbEeaSG8CHh63+KOJwaN4Z+IXW0IX1soL
qRDl1p8XjA/n6w/cP8JLLECPxeeqOizqaSixGPLcqHvrhnbPzxmDPF6IPEhD
STpLfhDF+nQwvAcmGQRRor40ImH4Gaqth87B8fv2x4O9ppOtw/ZDyvhe8YdM
U6ZS1u+m4/hBXoJrfXsd6OQbgHZ1yOJ0KmqOkio3mUSRhE6l7pFz6aKcixHD
DzfndNJK++HgWddUfd7CnnzSKuczzvvBkNdO/BYTv4vxlGUL0sCVJgK6YED9
hSAQ1zPrHW9VdyV5XKiqkcilNyrRCOQGWvyAe8hWG5DoIrmTWQCBHQre7ffV
lUVlCOaJSP53VS3/nPvnMXpVLGd4Ub7qH7E3AynizjU1rd/LBwCg3f8EK3W6
IyIl4zOwJQx3OAe8/LI4XNFuQGE1PmgIffJNgiHSPpZItJTX5TlzZLd6nDEv
EplcwASbcL8WkGKjzyDDIV5e4UFGO6K34kXm9TCoHWUzXb0FSQ3Gzk6ixL+E
3GbofwXYebGGq/PiC1EiMMx7mA+EMfGB6azlp/G3yGPeN4bBevlPu7wN4tlF
/LADTufCjO9Kl8OrQ+wB1QEfXbyPCkJ9StBv/bDW668k5RM+s4APceTQI4Ph
ekncOSyN1b6nAdOGMAJphOzG/Y2VKg/i87OML5W2WlXQNqDYl1Whx6cbU0Dz
HTVWDS2/LDSwOla1dzbQElg8pTDHWyFJRL2y8pkhahQcSHJTaFf/PIethWqX
kyyh2eg/XaqQ5AOX/0R9BTRsfUrbIRd4HHgsL1sMoAk+JQuhJ/6k2INylwN5
YaZ+vvk+29ACL/WgQGKWv7OHS6zR6opMaIdvXRD1tsg0GSPlJtWjhyukPJfE
gJ46y8ON9vrXK9tFOLWgIXLVNV8PHsXSV8SEGsqKpVDYMfDno5dhh8jJPmFJ
n851t5gjMpv3wA4wtA2oo4fr8ArWAtWv6xg+50H1BRpw5MsjjKFOqGUEWPvj
fN9hRnJ2jDyM/IBd+2ZPWDmF0HKZEJN3aCUcH5zUtY5kjtBd/q9S2+76gUBv
zWOWHG9EOvytxVm9u0DVJ+pxoBte4OfSCy4JcPUvgKnQlO7GuTmf38/yeiGY
2vgEVr5s9cPTI7m7zU/cVlW8dLusp/nLZQg+2o5r/gZGFwCWaPlG4ObiEZqD
3NjL7rwcH6Ue4kosoUBZ0r9v2ZyHKwt9gcyG5EvAV2mZrOXVGiobu6Kk9qDO
WDvED+XF0phq0VPgvVnyMOKGNUGGOJGQQvYi+FUULWai3c2llzOMLUx39jDq
aNWT/yHBWfRGF3jchyxXYzr13/CDo/hV9pgh2Uq8+TD0BYo4ITsTFRxvOINC
9m3cK44ABoBSWnjok0+gMZYUPTh1gQTTV157mD9BsUcVG5nZ8KzctF+WJwq/
bExmeM1FbqAxfQl9xZvmdaIuGobL9LW+kWFmJUW9rLjA+lmpDtKL8EWslKSM
fUct9v6cj/Pz3WsHCeGLtUlE2k/fEXWSJncoAPu3VbmxAc/6PNpt4jwNca6q
jjIlJ87uoJDqpe9agK2KceeJkYjA3sSSZvkJX7kosiwMrMrPLcfM2i/L2tl2
5SUP+bg5F/MB53ZwA/Us30ebZ02Hz0O1CrWXj2W1+FvKcAZjfOKAFzCJAzES
l2EyOqFMn7R1FbOJQhu7gqe8lV9sAgbkx+6Q0LDpVv6uqgHHbL0DMJnOrOSx
Kl8DMDjrOLXcbmthVYAlQpo6d6KIo8MomOx4zyGm/DgVaPzbep2S6pkBdN/l
IABCU8ARHCN4RdcjYewoUGWUNkd3n6W4WtPC6ZYiUn2CiL4Jpr8r+e//VXkm
6YWVIb+CsERQbg5t639QSkP0dqDeUlB2srszfEyElPnSk8X6z1yyD8ICydSm
VsKFVWfqzOTVrRX6238mQSyAUN0NwNJ2HLAuUSmHe08f4eFrNpQRYl7+fJcK
99ortR/yV4yLpABD48Fqjs9h1HKRJF1wOyn1vZR8uVCk7JOCz8sk8TZ8perK
X4/30yDPI4/CqvO7muc4V6e8kzZbp0zh1yLAf8OCnCXfRaY5O9ibTfF6qohb
PlwaI04i2QyldF4ccwPAtyNH3EpI5WQmOtqu3fy8pdSLmvnJr1V6zSou0Q6l
Tc6T5LzHKwU9gxBE+V1ai/nEJsb6+NX4HTD/z9nxzOOyKKdyDKXNkU+S4YuT
8vJeJ/xAUcUwfse2d0MVasRkX4P71+f024dRNhZy78z6Qu+B+WTdTWIh70GK
2dTATHf9fZGUOaJnBV8b7QWD+SMpRig/1xoWqe/rvbeKXOCxV6BI7i58aTL4
PLIb3dTA61uUyeFB4cpqu/Ms+5ToAwouZ5yVG6mvtZH0E3wtXisoI63ToTIP
Be2dqRutBXEimueQZ/h703u2Qa2alk2OfohBxQqM6od7pVg8b6PLJSPuuWqd
XI1uSKq9ayrlSPw2S6DpTpkn3PuQrLYJORbQYNkBppx5F7AIBA/vBVLCKPUN
CxTvtAPZgy2+ugpL8EowOmfMBJJv3s/0X30fbK0tdYU5PjAMs5EP02uJz6ra
amxFSxxuc7pkTUkD1yqblHMjCsuKdKAXBP/1oLmkGAYQiVuZBjcB0/pAAhIA
GS3lFpCgDNCKCHgPZnPJEoq5/ikIIBmVBzCyVfS+jIff2dE3C1G5aixhB7Yi
9QKkFvX1fn41/HnYtkwexCYS/i/2MI7xRh9NRElxg67b5DZvUhMMzcijxQI/
4GIEbj973teSUvZzab4vxm/Iw/BzxHiJVbOyQfVnVawWhGGckVAvvStwAJL6
qIx03zec7qqZeqqa27GN9Q3Rd21UPiR30rryeNI52V3kc3ZrHOsQoWOAKQa6
3HIzLGUhYBYKCPhbERpTmEHJGLM2sAGAWV0ziZh7MWzUwdZnTPmD1mbVs0Bf
GJx9VA90T42U2twOgwOgPRgBYzd3F6rsaZ2m4ff+RHza+x0rgtdOGV7ZfGTE
ws/bf9YRHxe65nKPCIAWRHoN2HGxtUZkacGQVrkkHDmqHv+LIL33s9QXs2tJ
F0cZvVCjj4mG9qnoVLqpSSfGV/Tz4Nv9kar1XKuul5uD7jUuacCQ8eHRVF5Y
LoYeaGXTPHZJoh5LpoAligsUgr/4CyJuVIFG3M86JndDHXZQMTOMbIbVREdy
WkcxiZHOqH7OW2XhUu3ErCqkGc8eVMfEDHGUeL8NuShlpl0G5mOE2pVi4qPm
+LdtoIRegEyAUq0VCWk4vWDXPAPwcty4X7G2zCiLRB+UVaAdqmG6nTW0/C2/
TW9wv/06QO/d9M03M3kFjt1DxVKsCp+cZWd5GMfm6SJ2KT6KwJuPwUdmUYie
opkTkixrcd/Ne+FjLKRZxxvbxRzJXpOYeMghU9TOr0cD5IJZmL+hHdlhn3il
pGVRXK1zeiVex9vPH0Y0vCOFxPK/O7WFnjanuTWuFB3JlUcu2R8JaqwJtyZC
Z8totQLzn6gpku7Qic7qdJCDM25qSPNW/u4ePeUnc4hY9spvhaxsgeN9UPsV
S4mcHFG0JIQ12/mLNHKR/MpgSHAhcyzsM4zMSRHoKsIidOU++6MiS5jJfVXN
yyKmHaZxayNpaFVr9QLFDbctg4MYDzu0/eS2oQ2N7nsp/8IORn6peUOKy2F4
8izRP0Al1pq5UbGDf9hVE3FWyYS5qCsVCORVVm2fR4WcLbcobG8sYmtMk2dF
FcGu/OKDHIciT1KznYK3RLccLYQnz51uzMTynVpeQ4VHuBWMiUgRQ6rNVODp
KawDjMKo8/rH7dEU72Ld4m5jDAOKwtCUdv035ykxu3URSBnOCIfAafpdBkpn
c0Wm1YjA4AcoywG8XIR0sCJfLv0l6TwOEl21lIAH10ht0Uw67aUZqVQpb/YE
N5IiHTjB5B7RUxbPjdSoVS4b26YqbGevNYGls1cab7EUA9RxqmzHkf6yUxut
LxWPciFgflcyZ7GqS8BxgYlsskiuDJgPgo3p3mkMu2DIfQ9cFaNclL2LvGtv
Jp5Nn+EjDTg+OA/+HJD8vcGu+2ZT/mLr5W4Rugb0wyxc1Mtv+KF5WRRnDU6a
n8Qstmu1UfJaBQaorOT8/q+E6XrltwmaZk9mMh4H5+1ReNF7wmKqvDcoWyxF
0w4fnsh7J/6HA4OtmiZyP/lBEXVCEtZnnWcztoZ5NPC2B+cdhFDRs4Ky8UAv
vuUIKNkRqkVYpvV8ChMZn9y04Qv1TWUrbTiocQ3CxByqbbYD1lPzHLE2x45g
y2gJYI+A54Xm7w3A4OYkgEcDdrJAJl4ZDtTGWa255+6yilqNhcSyllSgzcfu
jfQhGyb8wJ8VHegGaTAYJYtV+Dx3M1beF17wDLhQZDm48rTJyZeIHyOwADrN
KNPjB/XOac4ug9Pywyj9U13NfFd6/r5nmZPP65vb9kbktGZhPphDWRTHwgg5
1W/drMByrn1kVEOLXupXLkBJjFclZzlocxEyR4CFACZp8iaIorqLbztlaAMr
alwUeAnB3Pcz2JyZDgckPldCAlT0MyJP1CXe0wX9XdflsLcHVI0tnLO8agKP
J2GIHoigiluoc8cfTsAMf2UCy1AwYvdytUhmKPD/FvPjRyoTAhx8efuH04qZ
gswoABlRvAhri73FUIZmw57DRoHcKMIped2OgU5uMIoc4j+afSWMphhgx7oT
Gk4jQ15RNzOGx/1AgRvXi4yQ2oMQg1QSJNFrfXjZN5DAhwH5iBgeLMdshqYd
CmUFprbf+3pC6HOOad9r9a9cKucFdxTtSc5DJbC/fLxHsGl2lwUiCbWngsNN
XI4kxGrwtaSuFGxXCZt3AQDmnWfTrYHzWJ1g12jHQgpXk+yAyr0wgdiIlgWa
oJDvWsS99qSs7ZdDRTvIK2y/bsus8OsHw2XUisPyA1+Xz0Lj2BNVtuVp44eG
IEE5F0MuOXC+jlHz6OtkVQevlPfEx5cfUGpnv6QfEQcO9e59sH3qBJFWbFy4
0TRO55r+4V5cP3WfWooVljvHWc8Q+mAGtUs8NYSEGe4xH3eGHLKx0Rb2obMz
eezPrSTs4qIBQH5pt8DqXqJuyyIqHenXhqSAtHLi4YIxY7q+L4x1yf/vghK2
0pzi8SZN3iQoROi6ZSBD0mgia9exMnVy5w4ghWrvftzH6m3XraTGMqX8QrDw
NkzLhouJENqGKCdmQABvfhQtBfE4RznWkJ4ifu7MFjbkp9Xn3M7Jlim29aHO
rNjtOrb6NCH+nzXtt8sWRgdg1LY9CMD7VUuftc+xC0r4CDqzWZkCvQNYedpQ
XlYCTypMRWYfIRyhfNN/3cPbYWvXt7kgv5MdaxKDOL+TtrYAFm5EKauTKinx
Emb4UDOCuUCc79UruYRkabN11+dK+HesTVBpj/tpW8jSAQ+y8pvUkuX9s1ls
MUhGgTXTaZ8aB74DqP3vE1FsRwrYafu1+4JwdEAgnr2jCDSdyV78uoUWb4XL
rwnGlj3aW9Yl9Z3xmLdAeJ54nVxUkfa4jVgGSbmPJTWUcuGUQR2kUnCmaGhW
ds1kfF+ZyVaQ4OEWJ1E66+JCXRZ4fzHPgb+KmhgCY6HYMQhbody1lLcXHajp
Z3MtHCQmu6UlqOmkVisDG6DRCapwE/+pApQSwyAxVt+Mrex/Wt6rdR2LUYzP
yF4+yWmJpddje3Z1Ir+x+fgrcI3QLZq/dBbdN5nwEldmdrTBLfgvu9ULxWR5
AwnxiZNJjujq1dSuaB9pXSb22WivaYAes7y009P5EfDi94G/SBBgF0ZAXAm6
1Slv9qfCGO7ykfGPr7V5kCtltjv6mENSbAHl/XzVi/AZ7w7i+FKUoNpQQUsh
lsW96ty05dISdE7ntfpobmHNhbcttqdkAf5Tv2T5xJmhaWAWgVBYLORMbEpK
QAeXjIqd5rf9LP/zSpZNP1nPVJHlA+IkSnGV0587WXEOh47ea0cWO1fMmNZ7
FSMlABOJECNmV2T08OmAc8VLMjMTgTONkRzP/jlQJmjdiaHbdCnjWcTCTVJ1
4jd+zbTl/rQGES7sVUpiQ3I1FbBbvH5cBro8AJBcYUTj3zQCkdnPhA1taolx
te1tQuBvFBBdokhJIdgjZxG91WFUEa07xMaQcBMJahzX4Gswabd+WsXbcDMI
wK8hDymZdOaXObnckNa0yknvAXxw7HXWmiilPXO8BfQE5MTafRlAJBA7nUWv
kQK95LPdA9v05SfBQqdYcRclI5C4G74AGM6Gcv5CNDC/S9wf4ai4IwsGW6tK
d0Y1dvh5aPB/dEnYPL0i4Z52HdQfP2grLyzDUQz+F3LaqcigmCHnog04wQti
2hhGZ7sH+Y7JQ+nTf3XLiFbZ4H3GH6wH9ui9x4Kc0WjWGI2c6ha+MlgTawVM
JXiTJzIDS3z4i0a6qyd3/qjVoVvlrO3Rtirxu8fJdFwihfEBB10l7odk83sC
Os4TSnB7McaBuDWKEw27fFZMJoUfiYnlnSnBf8wjQXLG88xvUc9eMQean97f
fu8RaBpjN5RFFE6X8P3K3hOxOxwW1mZU3mGgGNXCDPIvR/5g4ia7fPisaY5x
Opw8gGq+pQN7/6jryZ8YG4RxzDKj7yfMKOy6aDagbheT8miG+0qiv5Hyi/Jo
hmjNj1xRGGehxL5YnXVwvUF4VKRAjVOy8t6Cc50yMPiE77VqnGd2RWmpFygj
ESHk3pORUsbr/RcqXMUYoejvoxD+fz3veR/+XJPtA1BqJ8mapzbH5MK6Z/5b
IgmwUHRXrVKTjmeG0Pg/yuv0FUeuwrIQq+Asma1/VVCo6hJnDELhQI49rgGP
lYjgIbqnFZ0SdJDXDmVIPFjaBtUfJkXAxx0F6sZ3MuvfB32ZlRNTtDkDZBoY
zrXhwiT19JyC+YOh8xP2OOWmbyvXfOW7wr3X4fiScTyBCqf3UqKpjDrwB87M
Nm77bkrPBpzLIgpOgzOFbzbzn3nM5O8AGKaBUdBWN/GRSU/WN4QmX1xf261H
PdHUVafXbeTy7ViaeQB0tvEmzIIYVIdWb5u5Q3z9xHgJWd3WdNDSMKhkmpn5
2T5gX43sAFrabooe/b+nR0pzbWdBi4zA9VD6v8JPfLccL14cXgOxIIV7gp31
4zE304M0TXVufToUuO+7aOU+8dNPz93PtmJzUoPO7GSuHdl1zNjd97bTn9X6
3P96Q/G2SIwL2TUMXStTiFc4YtFF85MPr5LtVdtIdV5IULgmdWKK9+u1WMbQ
5DXZ95TSuLjRwU+M83LKS/AynFtexd8lc2817JHbhhM/Q55z3tn5fPGARfdX
wrzEZAizMYsCdHhYgmxltKrI1z7MUgJxTLj28jcX3EUNhK8a5zeQ3sIw7V3b
P7Fxk+rnWI3cFsgmFfOeDuXVCyEyibCZfMrurI2HFUjrRgQ+hLOEJGJoxgME
Bpseh6Eexrhk2nE7BkEjmpbE9En2KHPoX0CcSjCALDVAjvta7uO7MgjgdTV9
+KsoiLPSP4Eg9wZu36iPz8BohgCxQHifFb/D5I+X5YzlNNqNQhpf2mYieD8o
HCbkY3z2DiSNYQPJIQGWsSP1Pd7DH+pA3qesAa5pKOceYC7Q3l/OTGTz77RJ
XswYxAJMj7vBuOiS4UuaibubWujIS/Se9g5bejQVtLMo5LNpVPYIv8umu9Vq
k5ZI2aGLBKTW5TNzd3YJ8QCbXpm76FGn0P5Utt9HRbBIvNXI5TmAisQA+rU3
nbwrRcgeZVN9jTkn8T+dcK1iqjC2/D5O97Ar8B7f/b2tNPWHnZG3B/7tT9cJ
k98PVZ4SRSCHNNdf9ZvjJAuocRSaqsHe20I3gt7XRM3etx9xZFD1BaR/S1gE
Wh/uvVjveCwAOydBMCZozBC+VgTVuOyw1B0821llegnti0x+rTuu8NnmuxSX
nNIU/0mwcSnBDdlp2hM18x2UmYOQKekJ2I73ESbla/pY7PYiId9nOyVM7ojh
rYpGSUj6d7ZrhYR+oOqSOn5xcQneA2e6WdKIjK7w3yNHuq83zvRXE1ch8ofE
Sup4cCCEctpS88+TvKbD4T4eJ0Z4ef9YzdfyQd5n88LRthNXrU06PptWmLY8
114yUdCfR8T7FcQIChwRbPrcHNTSy7jWA/oQfOHBompy2P3WLzxz/OUn8HxO
alNnhk9AjA0LTPqxQHyIVCGz4xDpGOcJPPiDYxdmXuSoxDu/zlVmbr/ZkqZL
6nKwsWnIIJm4IowykF7QFGA6W2mgKwEO+O3tL21cVCjtCWMQHFGHXMJzZKId
LOnM2v995h68mkLOe5MmIXjrKS/+fDI3uE7MWse0dHW4tk6hOWW8bRIzRVVZ
aljB0dgJiYMTWxNiGT0Y29/mp+QOy1WOuU0zxT31OdIHGuyN6vTIGTX+krfE
OBBpTeSjhbaR6+2DrtiMB+mpNJNRE6TzOq+is6/16bQ4XejbIYRT//7wvvK5
ZG+oMWSqlO6PzHx3zEr867PwiQqTXjwkEtUVd8QZm5fqzRKTgHMKpjWuX/mt
iuaWq+eMW6h8powAFxsENOXtIqrJboU34UTqkJziptVrilSHYkrvLv+ZjHt4
l23D8mQHbQzMEdrW3pajA5aN+rcDBJv5oAnPPnOC5SoYEQzLI8Qbqo/IBOZJ
4Zt57tILQCKRj6kHrhl3WeS/fv+MBvcNp4WiowUtT08QApZBeaLyw147WAE+
pEHXsVzyHD9lJeGPMfYsmBjKIAbbJ7Um7b0Hp7pJHYtt5DSgSlMqFdSHkykn
93tHY3q8lzYW4cDEl0qfxuQmzzpA8RoxvIV1rXFdZs1Wo0vIDj3gTQ/4QPKL
/xhdmwXBAUkSxmrqPmoS4zNxGg5o2hA2drSoA9hyiUDK+OYZmRrMUbSph7VY
mo28f9FmgxRXh0MoWFwIyfCVFBdvO61kwocGopyQbxfQTJlvJBUwZ/qGrs//
01J9X2/ACuBWiWxrwHWAQb7gCS+55aPOMgmbmQ+yNXX1ZkZS9f9GxmUD6zZ+
bFtJKQ5/NcZSDY/8sTZDGyQSA2fbIDg55QXaq2wcWBcUI9iIl+vQ/7Sa1Icu
n+/IFWkpnOXl1pKR1F3RJf9efkCPqM77wQDaaPm4Y05wMedhVOhBKPV52zpS
ZNSX35MJu8mG1gR9NnFWQjY4rK5Nd34pgnUqrUFQOtiHkrL9euL1Ny58u/nf
h6y2mMy6qCCGKg0Qn+J1mpK3RapydhRBhYrrsJDQlOxo/OyUZkCulVAYvqGU
MbgewQ8aS4UnUu4tB1N8Hu5MfmZAjcEurqVjCHB13A36msuK2NtpgnLsn/oU
3h7+O9g+R+miDm5Nu+HT0P28QnHP6kjEQQxxaXFd6SXWprc1Og6rRKPQ6czJ
ZhgK3UNVEUuFy/tyY86rMnnCQa/zpitjisPweeRM5ReJmIl8N7q/iK/R4THM
JhHdvVgWSIH1Ij+2BgvI0caCppAoxyN8DAFetvw6MmYReCAOqTyrl+H5fhnt
5QuXSpJ003kOkdquSkSbldFoFtP9vYs6vJ308zL+DyV661LGz8jZRYMu+SZ8
XTPyy3wdrbZkOsV1bVa0wjTBLc6SAXa+qkx4v0W/g8yINqLCxdtQo1zR/4TN
8UF9odwpXKEi1Exzhg4oF5ToLdlr5t6N+SnbTVS9aZJDcXxxhWiDkQDsLCAI
gMnWOWyYpM+QDRKSETa5nq9djNxK5t7mn8X4LSjCk8ZZMM2vSX4ATr8MlWm2
IrO4XD7wHSCOr7m7z4O4Kbdrx90OE4sOHXgQmAESPAtsLYfGysfly2GgEIUA
TCXSCcYnYBiegH9YQjFc360NZbXV2On5UambPbwJvhqTAhwy6BJIRt9DA9er
44W15USyaagdR93VomhA/KTibqq/RPCRc2XjMJY4S5Q/c9wl7UCiO4QOm8C3
AfU4CcpN718rIqXFs+oDLbimsdcYDnET9IXbXDHd/OqJpaYRnLTSiVDNBgA/
KruQdXrGvWc0Ggc7OtMzkXenzWBuHSjxrCZN2hqOCneME08MfXmxAYeMevKI
XVwi+jus/Qeqlo14aKj04CWzgod3BOLwIFsWKfRrf2+NOey7lP3pAIoz0maO
dIGUToZn3oRA6UwarrBdwrOWwiAwWZXCXqxcUZ3DFjL+zvJtpoagKMjBhXXE
9qRnMgAR7gvbhBqVbbFsKMybZ88jJDYJTPDdN4XYNCyhq68ub8S63bBn6KYK
gE/8xT7+9foOE/HYS9Cllj9lU8qIYqzZpuK7TUCDyETvfFG2p0QeFXzdpp4p
mj0GaBRoiPV7eS0UIsrJhIdYZzEOchIQYMS82mE8DGg0Zw/qfl4FvWetvWF5
dWjSvi9InFrO+Pbsgizsavwcdtn8cbrGaqyHiPooebA+UKQPCZjTbY7A1b63
N+5CsEaQR0ILBCPo5FCdU68c0t/ZdkC6859hBuUJ7AuhZ7tISbtQYio52Gqb
SYuh4vkJV2D5nK4JfhAE2eyt09ZwQO3xSThQdcdVuwPcfyGUdEReAMy4eJ0C
ey+Zkz/cSMvytYwVF+mEkYw6z+3Xgejz0VWwQTIQOVuJx3GrmPzaDQIOhGm4
SRO8eGvJzcmn/TEA+/iDCrnQPhyjXDFrGDVA+KhDWs1kO/B7vOhnUZSWH7wO
KH7dIK40/+P15qwlft3BrN55MsMjhTqwNMM+fmdSaTHjKWn+O31D7hG06eE0
SlnbeToU9Gg0u0TktkpTdvQHNRP7gtMjtm8dck0eGiTMd/qrVpDLFamFwhHH
uSpZkP1MZzUmlg5RI8pHKM30RMyjTiRmRG8keDXJPir1GACKq5CvkmC2QnBx
Y5v9+AiPUDk5Xih1vBUgeccCy0mkCbW2ePAMT0ZI1Qmf/3Asc7IrwOTuX/Qc
dCcFHvuOLLMFYO0GeceE+MndKoNY09Sv/4C+nfZHQWUTBHV2o4TlXAnHrkwv
nzoMJr6yqv1lZIh9OSzqaldflj8x+TFnt8kTSyGVj90BHdBq5M7V7P6rijLG
Z/HJLCK9rVMmF4mC5RAgfM+VWRSagvmWLLM7ggPvuUXNd54uVwiZl8PbjzHd
0Z1tAdipkHrGpspWVm7efFPDQCU9otcakuI6KY4JPP08DVR3oowTkjecE/CE
JsMvLxu44dt2r7/h5950BBpSUDDNa2QzvnuXk3lvBt9nEhFfgRlOffkD5jqN
a7GyuZ46cj4m1UsTAWbkO4T2rFzlTRedr04RIB7trmeLbJZXO7fQoB3EVhJB
H0LiAs9p1V4/ErgPTAl9T7fZ5XGp1AFW6BwyVGOIKC183P+ax0LzvKLF2H8p
CE1dn/SywdzLQezR03LaEbbhj6N4O9yKH2yVSv2dXTIemN15CTIPNdbHAJGO
O55nGJfviqvCYuJUMKcCIt39NfmKyYVyEvhPS4NmeIPeOAH8MiiRAJJANCak
YexRryN/nufXDNnioE0372mhR3ApciFKD8gbfGt8MLgXSkVLFoKUB2d2vPCK
uJqnR344kMHoFPrpNNms1PjVryO9fepkFazznQ7zawc+3gW4cv1BIb93pKm9
V8V2QO3lNB58KWal2XHQz0BGXI2TuOYm+weNRr7FMr0JFTLCgPyzKFEGyAzP
MzP7Hdj9mZFUonOafLseWLfLr0jpTBep+SUxDx8AfGOUIjW55kmAqehC4ubE
rNv8Qhs5pXVGe/Qg2vCi5iGyL6KNIjcbNT1hvhI02q1xCAW8Jn8SpmCBm+/0
l36GJyntGjeiqmfDohaDP2yxadsrzKASUlTA/QMiJTdKNEdivC5pe5EW6Cqa
vLIRK8mLou9dgjEXEMLl8F4p+Ke/it5oHrVAJFf8BaL7qAlLhNR994FS6IRv
zY2dQSdJ3E8IKX7wpJJ0y4zGi8+v0RnhpH6lN2mUkO3IjBJarT4aHVuqJLox
BZ1WR6kHWkeBf1e7pCVB4+/bkP+b2ionynTcnsnvgF6Y8davLiPcnJOeqkYr
LnLsRZ+UXx6+LFTt9++WoDYyOUcugw4Yvg4FjBUvWRO5b/2buSPMeEnS4YmY
rPnXJpDmpmmiXDIAWTaRJKnyINViH7IrRyEdH2A6n0rPG1hwobJuO/mdH/JA
8VfFcDUDX82uDQ/gLhOK3P10UYMK+UmvV7LAncaZwqtGyo7dUrbkabmk4OXd
BJcUs2+l8RgOgsBKD+XBNwlmmkiicynHM6lxZyIS+omZB2UHDVXAGx9oXexv
glnV61ZEOrnsez8IocAoHYEnSmvuIczyCmZUMCp0Ari7/Mb64+a5TrRHlxNF
DTeAYqmg240PTwmZkPh3qp7srIcOEOZvGjisU0Tm0QAcDBLMaEGetySDj9eq
XFaxY/9cvxJ5c7kJ2YNvH7sM8KJI+P6eB63BN8ylFUEKXry9uPIX/BZ+yV21
9hhCH0bvWlcJqaOvOk4sA5++BbNsdwx9zS2rI4NvI32Eqn1vrM8PTU/pQoW+
YUkwvCTA7le8fCKs1No6vMOXSx7MKcE9o2nLX0YHU2/EhXnm7JrOqWXtB6TJ
Kd8M+ELGRCD67K/eltWduXKioHahAL50aKT6eK76f0tShnjhe8r0ACtlxuDL
VGofsbUvmqBUOYNIMdbCHRVaQ4mSs9UfPMvCnwcByYc1sEhDp8KgwAnlirag
WnkRa3QxOUm7sfvBiDsMdCKrJZVGaZU+aDF3YWOrJB8+wpYDrkku7TDusDPK
ijBeKkTA3m/0B69kzBvIxYCQ41wRQaYhQK+1a5dpMk5TDmbYx3cnetvUUjHk
sGk69+7CZNe8qETxpT0mqPFY7I4BA6YUhBnAhdIGWkAnGtDph2yFJ8Cz4p9o
z0eDUm34SQMSAneBX2KxZmXUfJ/i8PXK+yYY1mU7zyxXquPQNwAqawLVNfVW
udqJdQAy9YVovoP49NGP5Db6O8jE3XkOYh9WuUB4S8BxkHCb+aT1+s3Df8YK
pBNHGLhfWbwJlQG7HrZeYHFuwN5ELLLl5C6AtD9ZASCaU6QSYydVyQS9xjBK
9tV5RV57njJVojJVLfWP6inGV6UDooU7b1o7R0StKSgwH11UemUXhqjKB6NV
i7MONohe4omAlGF8Q3gbMOGXWjdVDSHluwFPQUt0+zz3V/1E0Cnw2gz8iA2A
I5ak1VBwZ/ER8xzkglW0yFiNABY14O9SP+Z2NUbkcs6RXEiFXMxTu6IY5O4m
FMR6cdOiU3iowTj/VskF4ks5VU1YjqOhh22YC1bKcp54uo6IItB8fslp1Tp4
CHqrC1FwVZICvbQA3bcMEG3xnbo9+P40ohFe1/SNnDDhrQ3jDY2qlEBxf6K7
quykw880AtJ5L3Xo++NGhLWnIJHPGcCFjys7VcJrMyLMSfHGlotr5AVy7tcD
S1MsDW7mhUeXwkBiRUkFFs+FBqO6N+yIbOs/SEI2L0x5UsxfN9mg2YPMAxMU
QsFbz1ccbkRUIj8ccyNnoIRoGsGsH9qRdOgiNf6+h7ZxNtfjvDK3UFF/13eN
WlMtCWbwfWkcaMpmDAibWcHWOvvXvbdAAoceVMDHOqrdlxlyV647L3c9uwhu
BLMYac8lvFp0Movhhd+8WtsUrojOr9nVZLz7ehNzmYeH2mxK1DNa+usaRuBC
SMQ/BSRAcz1eRM3cFAPePpZ4SFOotSPM7Xbg89lhHvawzVB9hoCpPS0heDlQ
QNn9O6NcwJYSvnhX9xOA/T+B0fYvsMNdv3EKehePuQCvZRhyJAFSnlnTgEZD
6pJGQ7reLgqdw83/0ZKoQPFCfSBpM9CV8wiquhik/+KnqXYFk2WfCwDR4nSM
1iykepKe54s4NQibP1trYvN6rcz12+WNjD7U4hEfdsfl4wUKcOZi9Sfx3iz8
Mo1Ru50CcctziNzZkSYImev5T5hwYrMZRo4XuOZ2foRjKDr1VbX+IQT3C4nJ
Qe32Vay9mYJe6my6IldpSR0SkHRa5AWaAqCB843Ayv4vux5Nr/b3FJaVs1qZ
BvwErUvXH4HHmV3qNUTlyRNX2zW+xT0i7ubA61TClAkEG2ck0sO1HsslhXMh
LEPOPcxekEvbQxwmE9BdxoLAOU8HNmgswT02cr7FHklIjPg/1bBLS9rVHNbC
S2SKzN2OHP3xfkqDNuIbMlppZ/FeAgaco2eSfaXcpQcgdlMBvCml1JPecMCs
IzHP6XsqpmEONn4eMGn31qX/fVOaozzbSLnXcBiv+eLedPWzZqPOw4eEdecH
xmZdudMe5y+ufmxuxKag4r6nv8n6+ppzGZyxuL8N9N4GoGF8FCAf9StnDal8
0JJyPTuQZSmYEf8NlU8xT8+qwDlXrsnNlQEhTi5sjNJDcLZ4DfdKxr8kv1E1
TYDTFTVOGU60PArp8eXt9mguzDaSMCNWfTd1YvZYTuHG12sw1r95vc1UqXcf
jtuTlfSGsdwSVFCUkKYKzjRPhilCQlWsXJODSpsC1zVz94P3AhiWgYdMarTV
6NhAeZdwp03qzdohvQcCyjq4HEKoctrdL0YmB0WpyI4OIddbB8mAdbtMB9cH
XoZ9rCTe0PNVgYc9WUy/QuvGDnJdnzGjogfGpvuolJVj/YjqcHlh4FFjDeju
B3HkPbqNxKrMIdQEQsEWwHba19uzpzyt1hPmeBsN3QSWGbBmGSUE+BZDzxj2
+c1sstffAc9KGRZSn/fy9K5Ljfpu+skAqfpph8OUyYdCP7Exs/tFs3BrXL6A
kXfZJSiw/vKYCUQLy50yUD9JsEnYOK+LdusUWcf3ro3Hdji590g5yCLJVmmi
e3tBtHAOoFX060LtnWCZMtY9Gb26YWprw5mJRMmLYEyj4Gu92aGuvKaFvkym
tCZo09pKDmgpHUmcKNybizZ/fx26l5wxWLhkiS0wsyxzHYTA0+SUNhKEvgBG
AhJg914yaSIObkmb+kgHAK00CqVcchzIB9gWYqbSLqFSBvP16QqRjfhvn7ub
ClZqdeKCLZDnn34ndN5F4IGxMijMLE8f0pnColu/eGDZfM7Clr8Z5G7cfpKc
YLT+oIxo0rZwkQERZ2ZiW47s7ZUol6/BKlJYbhIMjV/eWZ749OY0zEWE8Mnb
bmJFLarocmV6VLXJP/mYDC2BreN0XTuUczyfF+eKDmc2EpjtyKoetQUpawSZ
+wEFcFGBoJ+xsbljY23lqg+D+pEDmRgN3AfXkqAfxj33HyiqRp2ylDziJLmz
erwLaojkUk9lIOv507gnyvTmZ2FF8l97kKGFtQpavcI2S7DQZJ1KY8cYp2be
1mN0ICoj/l2D4CBZ3YelLrY1n37rMBF89DPLvCn75hCf92Pvgv55wYCkuUTw
hx80npIrG/iHOCICXhUcW77Xo44phQeiewRMdi1ydM5ZMxb8WC31M6q84C2F
rh0Q/BVo5yDIeTTyBVMFJwEbAVeFUyq1GDjXAxvXV11i6lruFuBxxzRo0eoB
Tl9RwOoB0ymR9X7CVtjze7gplIsNzV00L0KcObgEcbjTi0ki04xV8qZbLI52
XuUSYv7vKjnFZ36Coa5udlaFjJ/wdjqltL18IJ59GZFsuKnNs1S1/0vMit28
AKnAAelQ5LqHq39R6HWq49XaPFZfNAFp9YPIkM17IyAXCFEMkgYiNCf56J0m
ALiSTAuuYFyUpFyaa3uXDgN/qBOuQq+3WY/S5ILs+xDb+nlTLhktxUBWBV4G
aQtTdylWRZA6O93cWAYHy5iXmixZ6j36ZPGrlaTCIbl0gL2RtaHeBlmfGkEC
VI4U5gfqx2wJeiTiOMtjhTW2QsXgXZoWjL/ZPf5h0Il5J3lgnXAxwVXEWiRl
lrEEws5/vXPMMbS4i6KafJCcow4GgQFREAna0aNZxHBHkR+nqtJmdmzLtt9C
BAWEwas7pk3AgMOu93/iaw2wxP7GXKa+pKh3oY7NP4Q2xk/8+uaH1gd9b95S
6XVpdDICZ9P9qCLoomSOR1uamIuDXjbIRKx8orM4RHUFko2rM0zPAKm/yN7i
dgqckv/SGJDbM9M+rerzxCRB8KJppZ0Xw152ZwBNbmhhGHarfqfdh7dzS2gk
uGri0mhg9AWhRIQ0sOrKrNoluNw7cieLxgeEeiHrdPdW1b4JxwIB5/ERM00g
KIueyWtPhiYFCb2mtJfemiyaWjZE7VGlAOIeP6tWslZJ2sUo+lbvbMOw2pvw
abJoKGXUzT59LXlREmDV5dOdbVXsKL8Z/inCJl2I/kQlXcu41kGO4FezxaeL
1HteyXL4bUjscMLGymhjmydXwBabaQo0a0MH1hzmz0oL7Kj5ajqe4M3IH4n/
DUQtrAptO94czlIpy2cDHhMdduZgZaaHHzuj20A3oz/luPuKnjI8hPJ9WIEW
deJmeyGX5lPsChaTq2PvApNvHrGe3yDTqxjlWBYZxwL3g5GAmBH2wKmhvBuc
LDC7ayFdLJmh72r3zcWoJOWPu08r9s2si+kTmHZ76yd+3QvTxWCyMCV8eL31
sf516XUk9WnuMfCV1P6vtiE4fUBdYWTNfLaHUyX3/HFW69BFR+U9C12bHL0J
nx/zaCC2REbrmOBcJT1pc9yWRr8GzVzYqsuV9M1/CUJ6mCSUG2TjdqCfx68N
0NK74w1gltLqfBnRfTc88uUhxbW2+eeU0HUhnq87VwLhpesEebLo44Ltta6m
jdPg/u9kIWdOxBt15QPcI+8zOwLThoHaKPxqs2owGMC51/NAaZhkLp8Odz+t
WvAwSqeNHP09WeV9E6vM3Joxu3fi0hTXf2nctgdCKy31obig0BcL7T7g8wDv
tBCBEvdFLA2LQ7lmPcTsFju1DM8/0MletynFNWhLmWjZTTrmKE2Ep62MydaP
dGFzwQQgBgZ2QHmiQ//POdlPDoDSZOYAmFiE4aWkcrcjgtfwg4lG3hvnWpAn
k53BiMXETi44HzdCX8tV3bC91mPcNYqpdjUogwitS4GJSQ57IdCC4bHPIQ4e
6UzDPPgFhgKNBGaZxbQS0ccEeOMRlyax36UyLZss8SUrEAPFQUV6HjeafuOy
Tls6cvmM6DmPxryTryrc9GVTNqP6uErrwzFOH4PB+tH+uXsoi9KSf/afE3UK
HFN7CE9jw2q6N5QNpKmAPlbEwEaQfaoEjVnGYOTeIzZhNqWsSKQMKDXQnBC6
FB6vYSEthey+FjNvbKdKGX8aBT5rEWmds7FDoRxHO7qsZ26WyGbek4C/0CB6
adCejd6FigSt5rtNXfhIftdGr67c6+RvoU2550uXc1JERqmn3EiulQCcJPg7
rqLRI1qMZS/9+32ylpHvzGe6HRKS6besdNnDyQGENl++XqGzw95MMZwOBWbz
YMlgc1Z0vRJuiYzw1Pf8Huz0vLG8+JWmyJmG5vawbWnc/yBH43JQH2oo9q4n
iYxAfFJ3jvMx3HQFAtD3sFFHgnDHkJda+rxh/sPAYiFy/XW1yi6TWDYBfU+m
gv2ske589c8CcK4CbgXmCbyLxgM5dj1uy+FdRjw/vHPZa7e96/pAkJcTBzHv
HlURHH5JwpgQIMD4fHAVU+8ZjD04P/1QeNwBXygYfZUR9XZqcvOODPNTU6Y3
kEPONKoJ4kUySOpkDOxTaBRdGkWI1Aa7ZuxlNR2GSAwECmn/fIjZBtiqjMDy
F6M7npDXe4RW+FIa9616RiMNPrl11in3ruf6W5RQWzONZ6aluX7B5/6ni/jh
ciO9dvHWbnUA57y/MrMO6fHkK7Svt0Fd7bIHPiJ2883zza9JDF5+SNg49n4k
qO77AtIYWUscPbMwl+62W8STlarVfaRYCoI7MvtGML7MqgPYyzg7HGgWR2vR
VR13TKttpNtG5x8h75BkQsA+KJ7FFoGR71ICCrC9xLFcgTq5QsDJcowh4qTP
l68ZKyP65n33Ti68nwUCtw2vzEEQ3dsvTU/OIjgtAY82GhOE8Sdc3GKJA6ux
KLtjvQGrZpDassMqE80sO2KvojW6WEXAlds9+Yj17gYJgTxf9ASx4WowUk0i
e8SjE+i91ngPIFEdOwLH1ZcuXn0kyDgC1G2lN+Rw92FxncvRN4rrfWslVsZY
YBRekSRMpVLop0I5pQqgY6FDNPhzQFlNu80PLIF/lXt16amjoOh6Zq4yP5ZL
Qf5wTVfTDZlCgLVrSekwlz8fe8yCoJ0OCyG+zpmZwRokfIKiDwEP1GflJDrR
p6/ByI68HjjE1knr/oSjIexKa0ckhUrAGZ7pRlu0qbewh5a93KT1nbODoo3T
z5cZADw3kjuBpjjFtvLMFGVFK6acb081QW1RhfEm/dbJLi5mtcIKoI0qQnCH
yFpVa+unI17+uT9ZVLQs8m+/CxLSUi/0avAkObOdZGIWTCNcX1n1xU2ZNPgd
lS5JqeLNvncTou695WaYJ8xG7sW05PN32mtSv6BIQwjQPyaMuMFDHOLSbQ9Z
Y1KgchfVW1uzA96PgvlPQME+dcHX3GRNzSr9GPuvvMYSlBEE5Gboar+mvVxH
r1AD/ygPcPHZIBuPaXo5+B6ShD+fsOzDXVpgnzoxvpi2sosVXhziqV/8oxyj
xoFjk3qUyjuRjQ3+XPOP17J6L7FdWl/8KQrcXRem/hwWeA3QUK0QmdApXhYs
ISRrsTCmY6MEEk+c+f0c1A2nP0cNmEoPjEc9r4bj/1O+uilmeT8SKlVf/CA/
OaeYtUo0g7C8byIoHdb/hca18ftkpGfrcwq2ahSUr/hT+ulsvBbMA61L113f
UZRiRjFSgoO5z8/8oLZx/WZ/7D6/hjiYU6oIRsvY29H7o/Ye9XaTflSvOkOD
1ySexq7XdCZbJX/smtxTV8HKmpgtfJdWu1TwpOp0NbaXC2coDjoyjNAqYq+C
EYE+gupBlY4Yk5lJ1TDH1zqCPMAA3QGefORF+F7Q1tLWKXulPGSOKfw5ud1P
xHEVPpKcvDXoLUqvwn6IoOuixOoyAAn9ydJ2pGhJ9fR7llEsnsUihl9+6kH5
4Ctjy/K5oXuMJ3mdIJZX7dgkGQcm0fbp5roYjqBQp3qPgZhU35/3RgQ4AbTG
qdPsH07liZs2RhkqUbTKNvE0dZBVJA+tER6Hang9qU/GcUJ/dIRjBcvPiUWu
PRYpe5/5uYJMsqQij7jYg4uOTPOteNgpFpJ2Dj7KvqxUp0rfYP4uzqPXgAbL
XLCI1/YQmMUbGow4mHGQpy9LlWAxHl/CaQHQCZXwQe5+Jr+Jo30NishYiu0j
X74NvwM7VFHSlDL3JgMlZOAmB4kc26RqC35JRA4FmgY/fHDWIi6RF303qdRh
tVA1bzABWqcU3WrIQOK25dzTdfL86BVYbP7bZBilvPE5nCLuUktVqbMPyhii
1ja2UlWVea8GkdN3jpxxLm9mHU3xz3yVBbintmvpPlSLy6x4Bt+ulIo/bsD9
qMDOPdLrFZwq3JaKbx1rC627aaWq4BKry2hwMgYkNabHnXN5grH14jp9u9Xg
4K7RmOa3uOFRN/BdDmQSbLFsajjMfXTMk+2r2B1cPFzjRRtVz60JSaKJ7cLa
TooWXDfFSvvzXgVvGmaznnNGf++57ltHRHic3WQQYRxzST2Dyghur/eGLCU/
b1n7sK/8xHqKcLntphpSOprNNvV0SlVMrWu+HeUCwYSKCM/Y+udzEMaYcXlR
c9TevNbHHoO9Elxr86VqApwIt0w4CU4102XB/ydE5T/jmqdTe5FizdD39TQS
RT9p3ai7aCozrrQaB/E+2ZHU4qRey3CXV3qRv2f0UW/kKlS1K+oPwTXzRSHZ
y0FKtmt94B6Gd3al+0yLR1RK4z0CDVZEOxNKOqZrJTZPkC+HCeTz3txW0zAU
Wv3yIlhfDiJkhkfetwLodOXWRxG/ifX7mFSMiX9cr9G7w2QVjoNe8gNqWB8q
eJl7YsrpQZBZaq82FCsJ4IhYR4WOrsWtqca210cBLLgUFVFF06y5MZJWPAvQ
OjfxxhUUJgCMpterzrHK0aFnwqT13mYHnPBsgkEomOixghsC14Y8nFeRCyr2
bum6uAwcUIXxPbA8HuMbuV2ddcjGwoGycOoq40yA6BDjRTjsiy2zjqKDwzuA
RawgahwcNMp3L1RRAs2iSBLDevFemoitwtVA2ZP21uPkyFll6k7k97wzhyxN
/b75hLQrhMyQlSAejr2oERWEXloJRHp5LF+b8p8uaYJTTyL5vbITMW+5jDwY
PJZwrpsWJd92HV7eki+H6ChkF7t6qd+99N96qNQhJsZttwqCZmUDYhA66/Br
P76j7tDnb9sAwg/zdPQi1qjvuMJbBE5qhqHYEG3JmxP5GczB7F34IvMYXI9Y
V3iQnaxlvSsETYW+I9e/CpGJd42H5R12aCjXCVhbbyQ4X7e++Y00dph/SSSM
Bxa0RngfWIKoV713xfXWYFD0tE5z/cO8UUG77N48WFsYP5ZJ+c50kUYXjZjv
Qjq0/ZwXzPfTIBMlvuPGc65sI9fdQL7CCujvtYH24MFLyUMJZDLiT5wOFSQo
zdmH05xI3OM8lMgA8zfTJUNwvHCB7ly7jJ8rBexrD3Jz6UynECcqqPpjWDs/
5ZVMTATeCAq40zf/sZ1GphdFJMg7/hfW7XFXJUtMltyr307zstg8Ugv4qNQY
ZlFpz0i0FguaRpvcYAvVPVYz/RvyX007IhnSlhE2y0ZpH7TOqs7e+xyI4CXo
W3CT7uxQXPscru0pqIXr3P/hhU5fTT3BvhrkkWrx8bnN91weaUYXeINeSy/K
nHPTG0KZbXtBlsNxa/aLRVNU/3xIj/jsrJicQQtZZnuVTd0lK+wotiHuzdsP
hGD7Jqg+oQadJM/sNOMcxu0VeGbibOj8YwlYzElKkyCMf18WeqRQPvssRli8
hQ1lPluSktOXRRnMapvgvsikR+Dv/INIHe9FR3Ksj919rrl+Z2raXdvuhBVY
U7J1XbSXPIb3uO0JcqZ3IcsVAreLmZMpKDwevtnw2vUAXfoylEjppb7u2YsZ
pJyknrSrcSkQUo+vIKc3G0cQUdGniGr9lAgODW0dNeOHsE44HzNBiTzDx0SE
YtWCDs8UR8SdGDYE4CF4+kqOcnFaK68dEEeuVc/optyk8HnYMgrk89zqF8fX
VX9igpOi+oxlcujPzVoGeUCUWQ26eX/tZ4/2PtOZj+td6ceLI/bAID8nYBrB
XfLQYB3HNcYY5AwbN26ukJJVR+bWhXLzHyRcn/8xMesb1JHARn6pAk6ium4S
82Day5tQo3Kpv35kZYEVW2FQhY1GRhsQkpO5UyLUt3LDcTDqTmbbMcMhB8oR
wkErjBjxpHsZBn/ou490NpExQtKDgvJJwhbausKjwl7ONrrawSo9tZMTHP8V
sQ85tNWyk485Ocsg3Q+lsm/qujMMKBQI5oNtL2G5BHtVED22xx2t1w9lPNYy
PedSFzaU+PO7fSv4ylBMUtm5Gf7ShB3b9B+NSCrIsAlZZGMLbxmddfOKXZ0U
s0L2hiZPe7fnyGQh8JEu9IMDUuBWSBmR4HCWUlq9Yg9bdxpByuAxHQZrgwVu
XiEesu5FDZoSiJMISjzXDti0Od2MGhPM8cPiEzklJ4kXFMrwX/+wW7ZyJ5qb
j8PtHfCyWpqzpLfxpsvjSUdvfu1pR7Kgof7s6UFk4CO6vtC4M3Gq462ZIq2g
8xQDpS6RxAR98Hi6gbvMPE47jsVgus9YVZ0HLGkwwR/q8Z/ARr8ITSXx4S/y
pcWHlBGVH1A3T4hXH3eBgcxgyMScW3sHrNBuQm925AnUsn7wWKlzVTNwxUhb
BAj9KZTeFoJvvI9ebRPFCCcHeq/kF+d8IZW6EDKGHk/7zk6ZNlhROGT7f5/G
DZwfJYz0GVzUNq/yXyD42Xv2kviSp3oQQmzKCVXHsaSsbmzYPRJhyqxfMgDK
M+Bh49Tis5J3ggrjtLL44sYwUBHHsOj/MTTNqpNnLI2lT70rRRdRih2iz234
3ldLdKBfstD79qq/OUMEJ6M7vKxcjgsAeHr0EecegC+aw1g6yCLZ48g1wEd1
BySFysNcjsZPSNAUwPCGKsjmfkxttDjmpsv2aPq4kQwCqC+6wSdwk1JKuj18
Hu1ZH5Mk2S6kX0tvM4GiP+uWGuLyfgP4pebUihSPr43AuJX18zv5bCmdchJy
1e2eJ/dvb0neu0x4tihHjp1ZJa4Q5EtllRfkjHrjYtNM2tqXna4nv10R6EUL
Yv6V0xqQ9T1x63JrwsJeAtKdMrgR0XBOaMkz12dpcD1l2c+GCGg05Pvi0g39
kJy7oGKEc23pXJ86d3Lhnj6OaTBhxNySn9pcqww+Od0fD6bVecqNBbPcpwst
Mrs4dI8g4jpVaen9qwYepUVfltatOl3ia4FmgaEZoPpgkkZbNdKznGF79eTB
9LZh571jfbJeTgP5uTZcVlyG7DK0NwhkX5qYqGxfYjRPJtwOmL+GFBhNT3GO
DbOIVp9Uv0k0XUswi25OWe/jHIUr0gy1tNGdFAYGkVLRUoMH/uiltwiMrDoM
s5ovVgZLhjaEG7VvRrtCZSwIVrib7d6AW9Xsp3JJ0o2+0swISFpuey0uFcQp
GYIN0vGV9rjf+54F4idCMaYkqi4L7jE0wdnQ2huSFeObRneraiPnbDuXsKhW
tF+5YQeUn1DoaM4VDp9ZxqPEA2m0ZG4AelWBApj85i06HvAZ0CWA+SVmERy5
IrwKq37+7Z6kvaCUhPSVvBFvRoaIUcolySxoH5Ryzb4ayq2rTfecRksDjkUb
dZGlJDNW9hqsFd3yZ0yScA2ScTxPM08S/FFE5t2o22f1CVJbL8QU3RvbGZUK
ghF+99hQWHo5T9hI7sOD3s5QbJ+mK/jKDt2u2kMKyrOKfOmr+06KyNTrNHhy
fPCu1TeEsIk9WE9s8MMHmj9QrIcgq2TyE+qoQumY+D5RSsCxsHaaipYEVjPG
SGynEFHN/Hp6VOMYtjglN8GJyOLe/0y9NJOmZ62X6tbfW/iQB6nkcFD3Mphh
CkE70EykVJW8cHwtvZ1se4ia7zU9obap07VmLEMh5MUar7/Mprrcj6eQPesD
JlVlRudBD9ojPRY6xddDawADVn3qzOu094pzhKTcVjYxcGQNy2FYVAhPbYc4
amnPc/bBz3iBUpqxd+xBPdTRLToUib6WaCaQP1GslzQvcSJ8aJi2xONxQZuf
7AKYe1xYKfSOOEdqmlr3yBO1MV+X4j7/Gpzw21AzTeZqbbj6afXVoPvs6N7m
aAOKNBxbkQ/kAhkHbR143qikPBcg8yG4rR7RSRlK1waHacRn2ouj5w/SrrXs
vczrSbIrdNa9t9AHchMe/ZThRNU9bCwhx+nqkPHox9nJ1dKGW86uRs/vYZDY
pIJSUayO10dqwpJh/Gw01+J9VFAFD+lxgaN4XfGY40qVqsP4yXy96RuOFH8l
unFzWSUx2iKbfpQpkb8MDHmeAMfgPMPrNEIfR1Mx1YNRSi8w8WpDuAaN2gwm
Q3cCmCxn8Urj4pjUFL8Lv/H8li4F4TTrS9k4spbT+sJE/idc1lbDqJyc2lTD
xq7rxSNZ37U9wK4vLXBCD0Fre/9bVeIlPzxmWigxneOpVArb+lyEcvbZeoBf
e38QKp9xharLbA4fAbuNs79sga6iJovPzEyoR00E5NBd/vClxrYOoEUli+Hg
dIW1Le3Bs0qXIFsDtBgMeFbW3Vqm7EotuQtG5h4RFltfZhcxs8Ik12RUeHPv
74pKGeTkBqcnLlTJBF2M52sQoHs/Q5eocnJyo7/AFZcBjgjj6chPLR47Yyp/
srWm+IzYbRwi59tsyphx0ShNCrJBAjF6ePgCvm/metoX/kczjgGxV3TIQ5E3
u+McR3oSpi0Yc/q4DuOTJjKYf1Zs+nb2rsqFgxKnyMS/nrGRpqevnL5039p8
xlmL6AsQAc5s6b6duIO8+L6nS92K4RzIIkK7eLsfRevuWJkbx1w15gqK6+cO
aCkIRiavHMpBefsVz2UQZvszoau9Zc+cqjsb1zhUjwyvihcK2FSYo43iuR4P
i4/Fphum9dNPf7+04Xu0qQtxMWFo3vs0xgkTeNKL6SQ/MSw2jrHIVx0CeSWD
oW/CcVIeExlkaxn7vqWYew+rvansYy8PJeC9KGm77c8Un8b0+pvx+xFjnTIc
R9umiruo80RgUQJhW8HQx3GbhlKvPITbfXRdADKDQNvONdEJA11SCG3SspOU
Vx6dfChAfqtNEBnkSDeQFO4dRf443rCCBnhw+eGhriuRKQGVXLtx56MdlfKJ
+lu5iv/xpx6gQE+nELSTkWeiaLtlU4XOZMTgFGtkPN3jkMhrnaqcXBq1dmdS
YIRTiTL/JgbD7kQnCsj3/7kHdSoSWw4P5MJJB0vh0S9GxYJzy7uIWAO7oC+a
F8OFcryV/OXpWdisnwp+SxHcFIYxg4O7doSmNbXqhMlxYDL0Cenmr0c/YIa7
0W9OzIEdMmCR/NaWwWxIH/7DWco1JKzW8hpTz2+qIngVZtQg8xOYKz5XDxMk
kl9f7zf3LRQaRarU+A43MYr2aNAgd7f3lI9CYYepCbd6a0/B/0vHa+2k1yxw
483HeRsyeMlBXZAoGa67QYJOxNhQ3ZD8o+3ADv2/4VdpjzhwaZTG0dPjPrYw
nDjwQxzMht/TZ4x1qf3WmbaZ4BPUI3yGrZ/eajLgSQDfAJTEqgHuGRYoPY7M
Y4hlGh+G/kMNO34ubBrxCxQFNiRDcb20XNDXe35+3Yvx0B95Rn+38dM1n1Va
nT8yxlqggXGxMOsBv/aCtl3AgO3vqVbs7DUuRVbi+Fw3nsMYAYRrZcy4PvhA
RI9WqyuYzyCHj/Fn5VlvILhULNn8ocWYQ/hwmDHhiubOgTIFjWWpcb/oHt3W
fqrmEKgqEthz9sSCjy6NdmUwDifcQuKn/MpxDwOOt9rfrXPJKrzdMq2sYSVy
JIKk2rWy5GmjBfMCtiEX5FRMs9cZxgKAzse9pctfmSKugHJdopLabsBek3mZ
x+TIf5oe2yAqe90ev2aN4hCnn59MfFcXyfogH10tMFVNKmHS1U3mgVaxvl8p
lYKBtH1jGXiTPort8q34+0u6FNQ8ZJkXQnLwZyAEqQ4xiUEdFdlkuQi0mYuI
8p8fy7mvVoyt9RtJYISPnHL7qvAqTsLJdVcSwvwlaj7kXC4ytSVZ9qnj79wg
JrpNFRWs84+xthEGztTNbY+aE4CAjORMLdDl/Es3Y1YBPkoQ2zwVKW+YnMby
ZF1siKMnlNXwF5rcRxWb5odu4kc37WOq0BLYu/ayRmaG+KkMma5xLqR6e8le
ZOW/pyG+a793tXuY7gvEdr6QG/XmXvHLVbjKgK/yFqlkLvBlakFMzpEBjeVL
inCVFS0UbRgIUNwJSxOQfOis+nFtIkeVdAoxDb7pdWqMY8VoBYy/LxwBjizy
nHQlXAoQuoZrgjP15FvSkTMdlSnWXEjTnKYX5iOHwHlvGJA6ipC3kJY3EZpM
IwnJ7hhAZbKQkxMmZPQOkKj3JbuFGwjbwcui1ONNrHh9gwzdFGp+4aZh3WbY
r23sKPPukS6taEmDWLxiSjzhkq6oGCXkn9gDY1UQVNZcaAm84KK90cBAn33A
N+BNwXO1fTjnIZSk5HeO3fWs1gJyhmqoPksu2CbcRQl1VSazN4wgXbcelu6k
Af7K0WCQ54JIGM9uGOcwCZqZjpqu7Bi69gIX5XdjqeeIdrQhJ0Db9Lowh7hk
OlTpoktFihipHRI2lxQIXvfhj79joy/l6yGPU0rY+qtsMCDgx4BvDUtp6cN/
9OP4VbxfyT/MLApPQM5L+0T7Q0f6XhGt+UukBwPUYgx7AUqdfzhxDiw/Whah
lM3so4+/0pvtupkQR83hI0MC9CVYuQktosDtKwOsEHNs2vQhyhqyYlrpIK2t
u1DO1B1ZWUfjphBdD3nmwDivPtybIS3uCyq5rEdCTL4fpeovTV78woJGLt15
5d0tatwMtqgNmfcS6F38O2EFIi2VNxefoNyWlbEkNZe0w8p99ROT7iAA+DzB
86toNKFX7KAcSWHp5Ev/DGe65wZYJv8I+kuWYAZ9Kr19+8/E1efp1u5D1mVo
zidHmFxYkQMZSf5+shDrvVF1ltMe6V2M4wuHPQq7yzjGcLSuJwkOw0PJl4eN
gU9QoDzDtZbCemGtmwCdSGpJoYVj2xPT9sjL7oTEPU7ZboxQwln49Yy6pfYR
RScCDCipncRgnevlHz3RNIXBvaRQ1ZIV+O2RkX96WuCvQ+8pk2QRLCRN6sAj
d9HfIDpKDi70EDwC/gQpqwMrLBk8w/jw1rDCGYm3OGx/j58DUKKcf1gGdqnO
tMLG+QujJHvIaDcU4onFPqdhwBqHFNi6iNH/5/ucvbhJWkRe0DKY8xEOxBIM
3FPnhmpsnqLVJ98j8fo7egAH/PRdWEDn4/Q22zuzNA2LEr4d2BgErisO1GE3
JgFB8rkHWOrAVCEW1Hnpi7LzMqcNGAXWTnkHVVm2PbXc7jkvLu1YdLhGjwor
opowi2DVpKvdWPVnCpnZhMSf5vXjGd9V7WA8ByBLndsIa1bnvzOXk5+RoPpq
OqvIw+EiAAtvUXhBRFvZr2zIEHNYZQfin94+jY0gvAIqkOiEjwXAX+vRCAl1
A3y9+wZ2HnFrTXrO1lNzC8elIRx6xDveAkKheYilZf3HejC048hNdBmlUTcs
VCHArtPtksYMyFBHqS3Gyo+GY4z4+yIlQEeVMXTrFRiLDSlas3bu8dAiQCms
BfR/JPaUtlCg+9VV7y+jFDXw4w/sbJ//ZgvDWlfMpPMAviLNTOq4vxJVc+iH
KQBnUlSnfitk6anX8M+ykIkoD/bDy+albMvMjG6smxmTIL9QEJxYE95fT14L
Ly1R7OjhLcKklQX5/8Qnkq98Ut9dEV0b6sDHoUa82kwiaBsdD+7+jP+jn13Y
Yvf24F28IdfR/wwBPvmb9ghhnUAnIsZSpHbPU9IJsMGeHtuEQ84IGkEm9x2W
yreHSWHM8wLrmVZgmNOFZdl1xrSM07nod8BtvH4vMVpPiO0kbgDVir6H5RDV
VdZ+Gr7Hss2Twu01CM/zqtNmUnxWpTad523OZmI31PIIkiBhOcilT4g7Pimz
aQmfeDmESDPixlA7KPmcDMuyOeKnTcBeeaosp6u1pN54QoFcXryoivf0VtEL
EKP2xy6rsWOa1SUorNX/wKzKBUThF4eR8Ojp4z+1gBT2YE5poUFR6WTU+h/g
Auz2FCtc9Y5hGdZA9gN39A+ncMnXdb5dTav/gHt6nl1heX0Uw3ttWpiAVXyt
6nC6VPEtiMqmoSrg0cK7+LVZkjzlQZjFh9jq4lqmuXv3fqm8a4+pUfDiHX51
FbRZW2FSWRc8HhYhfdQPLmE8CQLzTSnW2RH3pMwi3AMf68wn08nzflB2mpn+
0uNQnx1ADzCt2Hy7uAojmAsjc6l2l+srqRUMxywGHgwSIoKq+ipwJKCO+a84
uYZMMNwugg6kylpoRvwAfKU3LdwZ5rHdagITqhg0qWiIz4m/C6j3xsuLLHym
iS2Ip8VzmKAyPiBOIaO8YswyG/bhKSUwRzZJZBUmepn776BeG0Z5c6eJDoMG
9vkI8WYvXQAvNUBKTEe09Jo19lrPyyrKFc3Y12hqk+D1OratU6JeIWxjpatu
/llzqiEsZvOy13qiGOXaMtKArUSr0zP6RE01nndrVkrsJnUXIPhMlvUESM7D
qcwmlocICQzd7joF6ms+/h52+UAvHjoV78lEdXSsmXNjNmUSIcgFi4S+Ou3P
0oY4YP3tyZJ7fiUKT0kLrlB9T8E5HIh2vAQ7doXbfh+CB5HQVMY3PrjztDdE
B2zePratlWAEXVzUcmRhb2QU6VXhCtyGfpcwTMkc6EHGXLsz+oLYorA2nXZq
L2k67qMLTVZdAld33AitIaF19sFNCt8B7QG5RYK8zGno5yPetL2SPRPrcXjT
GipBvB0SPvOIjGQNICd/FU/qgLdNinIdErnB+pEr2A6zkMJOGDre4jW9grPS
MTTMMVqodwNR724DE36tcTa1KFQ7dyGpryMuaPM8UmNM1io8AuGO6AvngICL
JA5YJ1jYXTZWZQAo7fY152MP0oYd7ZCVEMDfMwy3zOFb+ZXAuFQ/+H7X68eo
35e+B2rfjqHy1NcYaqcdufnL5rhViwLjsdd8jaFwPd3ig44V15JHmeTFch7Z
OyTdoZFVEA3PHIvtyrbWK8b9WDXm5eYJu3hI6KXx2kTzFGvnWoI0CUCAMwb/
RH1fujhMtQdI439EAS0jQMCVe23I52OpKL3OTNuoDPHa9PV+GKCqwYGrYnJD
LYrOt8neshcg+tyd03tBnDto2VqkipHqK81sjAfDc8olhZRo8RhEh0+4XObe
2vpL1Uw2NwlRHkwrFJPxxmK9d/SvGn4BF7TZv0ULsVZS1JfOFG9qZ9vran62
W1z7ebqdUwHwfBEOOtaImIMR27bon2N9VwWyj4mAxQ4qB+SCIEKTAKzBAVXF
iwWJUnKfOm5/ZrmRcNvW63tZOa8DZymr//qpYAbIx5+83fUgiD2bTqPn7Lec
vR9dYLBrhxqZCJZ1wBygv0cQ3QF+xPoEfpJi02CCXmDtVkG5aaPGXEczO+kq
skGOWQZZBHDWv4kpeNLSPsADyLV0rzPrK1tOdz22Rt7+MwRaDIUr9rEpdZ0g
9ZFTLp+cHX6m8ljS8to+clswWuPPq/9va4D5Wk+mcoeX8mxeoKobDqaAoRan
qZ6SWwqC0au2q4M9dmHOPK3yVoGpkRLjrvPxtOxEC86z+S7CCSLj81APB9bP
Og8BEjAN30h3CgBN7cz+9lt06+RXux6UA0dKFcvn3D5/bz4+VPSEni/U/uCf
iC3IQUZpAhkVxBJ9SBaWRbouV9HZOoaPVCaG25ZZertUyE2UbPkUOt1Zfpx1
2dg0x2LZky3kGJU0OjUfjAs9zRUSDaQ6tQU6Qzkf5o1wTg68joXH57EQK3aw
GTQfRE1QzVm6QTJTal0afnHZM9680vm4H69k/AzZPiKRSIDzOkCU9SBVYDPk
Rz+eeZav3g4yVK6OCfOTfQkBKVDAwAXefpP+QlggA/swAMThnQh2cuD5l6pV
ZcrsUv6pIm9wlcsCAPjUM03tGPUVKbQBkrXmAmJHVZ+ftqv7nK7FMOmHLcyk
hiPK+xVoft7dQsUNSD0NDjDgAadjYk2R9c2Tcg1/6SJJmYF9A4ErKp75D8DN
Nlgc/DkGzHXmNWj79A+tgYncY+92qpTFC/lAeqTDXd+0+gaiJmoNcAm1ovP3
wcwq3zMcAYkOkBmAYOMU0cqn9BGP4ZgEFa9AmPSQBQ4TP96+2f3biWBG4Acw
HDqiWKJiZB3Hf1FV7m8djEs48RcIwdU3W/VBt8GpOlNY45zrwbVd3v8RP9lp
e692nEZvtTPk49ZitkPK+86sseWC1GwZvHuvIdFGzQaJFBmjVheYSusLB+nl
ODoE8bAdfx5MjkQcai7Cd0twXgq+VoPcYpF7zcYmFx8GyL8oiIoEEGrM5nXp
TWji/kTlfQ6ub5AapL7ll02f8ODgo2HLmDsmjmTcWDwvuT6e0mzanq3uCQGn
R0QIMRUv1iH5JZmk1tft+2cQv+LQrKctvTvaHopzz5h25tcHJGlsz9tst7y4
6wQiFr7NcogGf9pifPAc/bhwbj1iYICKPEetpr8wRd692Nt78J1CCmL/mWyu
s0Lqv29KQuY6OfZd8zOnS3WfPL7ugKV9ZqEPLzC6XPBEBPVuaq+xtv555sFH
5NMcm3/iPvatbk13xZIOtXHpCkQXImU+Y5DzxxybTiPV8R+c3nsk+cSrYLwQ
NgZ0hTjunwdj6Z2u+hJN2hi61teev/HJD8uSuSl6A+H3ksxbquRBnzPefWVf
RRclzsMHj1WtvjCI2tdmL0BHU7a4hLqp60MceSAjbBEEo4ZFOMdZL4mgl6YQ
fTDGARTzAI7C6c4OFEp7qswUCXZhlDLHmr1Zn4KkteDRBH2i2kdFNIr0TZXp
nWMP3VB7R51GhWqwQjnp5NW/mQasIEBjOcWtiX7OOX2wBEBO0onIahCMfpZP
SrqcoZukz/8HBzPy+oGVrnUMuz80zM/lK6OXNcwNkWA8kTCCqAB7E03HH9iN
jDOZkhdlz1oP+F3YA8HaTBK0KqihPItyS7VB7cugbg/7L5tbz3mOgUY/BvKR
KYtANSe3E3NBHp6C3O9PM4JD/vCLf8DuJnEUuflP2TDBf03L62hf6ChMtN3A
Cxr/BNo8zGgavr7WZE/Tr/0Z2M4Tn58tf0fMqwyjzYerUu3Ttiju9jbjb40d
xfHhyjkhrw/lclolANZBnLwc0cpAX0oHXaT9PS1pbiEMLHoWDuWkYaYGpcwh
FDYVUJCRth1aa9gT7fmw1Yb8bfQWlfcejTh5r9dAVDLNsp5b/XpEofg8YjaY
EVcIpw3ksH7V7K9YOPII9xD1zMKhBSWtE8cjiun+j0fVq44aWUmHDVORMstu
nXwcXM0moGDRhAnY2hTkGGHtgzcQS3g8JU22RaRQNfQUCgbELpO0shu5NbL+
L88QQ02KAvOULWH57+u6RBAqdUjwiVR3q1mLrPU6tWSbjhOoyNZuv7pGIjOe
pA8ijQsU9hu1rNgHW4bd1ENlGKEESBH0t9rnrePpWBpOK7svwzVvZF9XpY8W
W/8NURoElz1Q5/p10XZb/tl/UXspbHGuZPa1TFSIpQzyRiXJtrucq2ce5VGJ
LuNXjMB4cl4qcKtCBPXaDrVG6HRF3E3oMANfb9e82+s2TkNGNOnb4ySrGKUE
LKlJ0nw1w9jhdJkC9X3mx82/yJvwN5XBEevPg70XGkxLAmZcZEklMF5cQxSY
7lOcsC0GnDE//pPsrBiDYDJmjYrRyKPWfFlzaz4khFOtYyf+nj+4AIgyfbao
4in09Y1ykeTCfaT317T4hWKnrc8WVWrMW62NfUvkPDiCsGRbM/fv1wNNQzvK
Rbxd0n2rcotMxgYI/rdiwiAqqqAtyWjgDQcFDDjUjHn4CHtRH0S0Ff5AcN2M
G7FHh/zzrBARRo817rj8FXDBP9s8hVs6EvDWeIbP0wA8E3rBTRPx0ps6tDE3
M2ZWGa2lQcqZyvUBRYtlDYrdDUC4TqU02oUnHAJMfnaO3oBPlqdAQeVd0fZ/
S8xvKig+kSp7tU/M6Zhth0jLel1rs0yHuhRSWV44NjI84WE7Fl8Ih6qBGU3V
uidScsdYExhi7TAXkuQ+g4G5RJ5BwQuq6/t/cKpncP3ms7Kut8/SEWyXPpks
g6Wn9f4/CUlCbjGmRRfoKqoWnI76iBE582zjW7fel0NRXbHOuVf2zF/7HhVV
YVTlBuAK/qhj1hWH+HTy/l+M0s/wd6WkzxuQRp8Y0fbfVuBwCkVwgE9/ycnQ
2EsgMJeB+yMqMbJSuzftzuSSex+4myaGnoF/PtmbW5TZ7K/gTbZsFau56SfV
W+1M1OTHdvisYllxHhR3YSUMpjyFdD1C4gfKBwsJgH/vpnjymjvpdxHXuPio
nvM/ztVM+dTZNcKrW1HWjS3In3PBKhUvjTzTuU4Ib2Zz63sJriGTYkr0iMKk
ofW+SU9dhJHze0J0UgghZQHe/RVyvgDvQJs5Wa20eAxPg0+lI/1Cfm8Ekr4p
8yMiHz0bvt1V9leDlfXMavwjpxjmQgEeU3tmJfUbDK/K+tuWtMywR98UKR42
b53amkQ9Hbrd8c1B+cWDvhO9ps70PUXKJoCfcZxchyidDN3zIFc7dg8TKvS0
CT9mS1gO4XHH1vEjAzhTBsYoWbZZsubF6UkxUo8387h20dMDi1udfRZxJb3V
/LjVLVpPb5ecbkaT7GkEtaf5z8PJ9BnNRt8uEoapBx+XnXLxhFLmSJdc1OnV
+5mMzkK26h42yA5vPBZqGPDEM/hGb5+naL8J2oN2mvrB6L9m/7QXQTaufpTg
Tn5WkJ2CvskjM4J324Y5fJ02daQ7dmh8ThgUayzXuTaG8Ip+3Bio2zkqEzSE
EiCHnBHhYOU1axYbctP/7AnTr2Zq9a70mQZbZkZlVonIXNzPq+mKcmlmqyDQ
x1sUNEpRVYS6qF5CDeMffd3le1jhZzX6bDMAG3Zqy1MfaHSht0q9/p01EU8O
9CiuYNzZQKkJ+AHX3xwgKUiUQe6u1539knfIdjNHLlF0PIfw+CjVwqhOTnmq
2gjLIJFZpB034weLmUSxNNG3rV5oHmQ/JLDb3erfAzY+shROFcKMO4oTYfTM
yu+J21QUINLw+yBNt3dNpLY7EHLp3mMkh5f3L4qC8ztSglwlRexyf2XeWwKj
mIZIE9BC0FmRCT2N/cMDdSjwhdZyzl3tJKE1bOx9CQ+1J/l1zhDNpM/IOvOD
gpgHw8pOcSUUpfXboT3jLtUh7CRWhFxYFdjjZaAbAink1betLTfHSUjUwSjL
bQmvKbthK5iEdzkZNCsTb9YdohK+ilOawHNVLnSGwpJtZJ9EZXuIfEgRMmb4
KtUuCbTKH7VfAu+sSrveA9e1pawGIyRF1gmVw/yszJJDJu9syH9gBRy5r4AG
Ny3Vznl2KGWujAYefERPIhroGk89wpudkMAH/HNfFBd+Dldme7yGAfv4az7e
SRMa1AgHEwV37h8S4zn71+WahXvZgZ2YOVrLTCDGJEna09HpuS+JtgrCw9tf
Qyx3X4t6h04dmVSDp6pyHJttA7o5aPlPqt4+SYb82QBZH73QiLse+giyoK7K
tpyLo+5rKboG10MxUu0jX1ST+bpCA4RtaPNsn8l4B4aohi05XKKaYo/KOUw4
mbp7Fch1iOyjmW6D8L/Vx8cTygioM0pMFODJS0h5owZFKcCfNvFEn9YBg/Xv
IokHwkJyQ4Q3qNulJPMNIVszybtjohXOzK5Zc5q0tr/X75NzxMe0/4ytrioi
H1oZTgKYqeIkKTuF8vaSwjcDNoofrSrIlDcqDV4mgo/HI9fy4PPF313NZAT5
nLBgw+NCd47G9z6tZStQEF01WEz+0L8TWI3j10bi9ivMSdOjuSthOPO9kCfO
T1qVd6ueA31FC0b4qjhmN6AGnV3IIQVgXua1wSUZ9RM2xFu0NrDhso331dMg
rzQIZ1xNTcJqbnely4Q3+Bi2BMKrildPR2OKeqs0/Cp5RtTamoT6OMbg/Esp
cxpOoHYBy56R4MEOUHGyn1ebgBA+FqdhYTAX7FatmnqdXbvhMx9XMMMZ0lJa
ClmKci3fwoVIb0gfBqFWasmT7UYQRVitDM9baUWscT/e5ylm5dpSRgrtwoFq
iPWc0Lh+hLKwfdB6WA4X7EheSnUimfcLmBVL5NzoeNaR/3OKTusXNhapRxbX
tbxd829bjmtS8fZRtq6IVrLYRyJjYsbzacS2vNPJV/8ZUqcUw8IjnpSCmxjU
basY8nF85LdTNKS0DXX9JsPsK6wiwWXc2VnNO9RaM1ggRKp5ePkpWKGxnNLH
Dn9lg72DVbYHehDqo37j1rWrhszfLNaAbVHwqf1EEuW6CK6SNHTgqH7sMOpR
w6VxlHe4Wc5IQ575sSc5jP8/C98AdbX8aFpErA6GrJHMltsmx53+0a++d/kc
FWzCWafuhpjztjEI0b8ayNd3E+cLAD/Lt4Z20qTVlyPzPR3T48cJwSd68pWx
LWTLUtnwkTzom4nLscXNGVPsifhAb5yXEPRltHVVBAYJ8yI/5kxCzqHG2Idb
aXSCzNRg5EUHcj3lxCMG2NO1RguuHcmK4rMvcddjNwsjoVZFOSSLWxMZV0Xa
eMGkzJPG6/d6L6AwdB6+reJ5qXg6SzeS3pDKSu9dxHIW68wcO0z22HS20+kd
t+kRmndR97aK8aX07mJK3BnfXLLyUU86P1FwDZiEIrBm0cHjtjI2dvawy/S2
3Xk0uBoLbEG95zLea6WSsBxkHOgQcEHa/HMSgBiNn2AHx/4W1nNxPNN9Kkn+
iZixwdDc9vzrqJLdS+u4jvnPoFx5rInDylsD0nIHdpHTWlPl4LatRGFL3yDD
3qbxIwCENXCqlNsj/tOY1fFmHEqgKgoCJRzwfZp96ClY2FYuWZsB/aYHMwmO
seBM9gBXWhRVIAOCbfI86ygt/bdUrEdnNNay9VUQ2iHAluwdFLomk238jv6k
87zWG85L13lo8bOathoOfCSNfapD0S86ou6HMjHilhb6Doj7GbNoasUPrxIJ
h1U3x2X0/VfN+wzQifG/ZCCTRvztM30UuiwAUkPxd0IwxwmJZEHlWRUqdPSg
x2inea0We5OMB/wXc1jurKti5Qz+2dAoyZvsHo7NWrXSWYxyhOmcIsxB34Ih
vwwC4l5vYKCIB5YHcDOqD8wfa641K3wZtN1qNuJBFXJ5XOGWsQyn8Nf8fIKz
v0p4h3hxTPBmngxmQoCoe9lf7vs3AOFSKbgTFFlAm0H7Mi2ofkd2pPPnLH3U
ZXR7Z5PbnOL+1wcjmQbrrA54TTCObmgzxYzUItUXKHvhXeQINP4HomybpjjZ
e8e0otZogCelPFm1en1MeJHyscatI+mdRqYCkBSI4pRDEK3ddFqDCx+cbH+M
N8JWJ0kOVf8lSQA4GElFmzU31dvsP/eldZ9ifhEU/zOLCNhPTMf5GehmQTt1
F290CQhYNvlXE6YxmdUzOaBld7/0BFa9fE+AdfFUl/d4KptPw4ci+QrdRiPK
kBfHRBfL57N922IJATzWZmntmYkWA8kHAE+M2XD/OWZaqCKuMI83Fy1G3arE
hHLrO/Rx+nS0iVMW98fO05EkSuQ6M0qMD1InATnDdR5dJUsi/YQWH7xOendu
1FdtArz3ypukMClXlqlAlfxP7tmgTuahIFyVXEF5slf30+XjWLvNBiWsakTw
ik+CfLx17bepgWjJIKSGaR9qTnO9KYugecjXWrfuJMSmbXG53dD5hUqIcU5r
HtFYQ/KnCwip79DDu/eE2GfWZ+MY5TqqHfwhTDE6nKLPODxT6z/dKAy7oukF
a4XDsiWZU/DMmqE/0sp/wet/yr8zbRvIAICG81InS8lG794MWuoBbUBXNAnf
9EsjlKjJRJAJGY3I+mZTK0RiYiToLX768PujmkZ5qSIHMFAawVhC5Xg19JbB
KS/bwnKJUvlJB7udGX45O2pHkOfMLACvRKyXXvXa/KmrBzuoi/4dDICMuZyH
FidV91GXRRFmWNQUHMTOr3E35f6SDRnJRzhyrMpqmnnUySgGHRSwVmj3Fcot
NozJSVw0x6UbRVvxifd86cpEAADhhfR+t5DSCJoGuTRmejqE3HOybziKahsy
Ag6/5TVDvZfoxuf+YFA1XBpnmBnhqRklXxu4GnNo6FoxqM3ODfOXOD1Yr7sa
M4sqVj4MYQPwaBd15Q+O98x2v2iwOn2IB8da7CLY+Sc+p5tCcWkJqk34jjC7
S5No2S6ljs25/N6944drKY6FTLNynJTwlF1CCxw1iA06lahXFb8FvTueXeUf
et6gEveWLI2Cq0jjLl0KkpDZ+OmkWlEJU0mI5vdD1VGyMtRID9kL0xY+GkKq
pyMTT9KuMFPyLqPKHArrHX7BzWMc7Qtew6hBFT6Pm/uuAZFREOn62xWUPHDg
cWFCszdfcrb1AO8kjVWb3sA8PdaVlAZGM6fMSMETVzSFTt8q0rRvbqhUznmt
95jlJrCDLYrF/8/5QIdgUa1ilgsdsRulNp5Tc+RA9ps47DEu73eKf8AgYPE+
dcRbJ7wr2FB8XEtdtMTC48QnXu5LVx5aWQJ75Vim8jdp2pDbof4YtV8a+u+g
BFLKr2ckN6r/tDdpAJ83KdvtyPdWCWNd5WpvC0/fZnxnPUWxfx1uIB0U5Mr3
iiNRay3JJhlkk2rVJ1KX+VBKFuQrkbBifkz+FlvACPiBhNPB2iOrI5U4zhaw
afGLzz1A0mNYNy6muEF8R50w0MeFlI7LYLocN0MbdpTNkwCqtm+9CV73X0H0
86JWOMPZLjLag0nF8K+JrI9GQ7YnfGcIkGq/oKOyVrrHIG9NmqBa6mqdsUBh
K4DVVESBGNM28Cvhp5ZfuLP6tj02T+h79/6WeBG8mctMfDx0jKcbHIh7cZCE
xUJD8PjuInD9KCCx2J47nZQBcUQNH99IHvWSSZZ1B7ByAnXmaWG96gJIXoaS
n/Y+gkCCDnfdTCKHsfByhkUxson4v+mWt9cpwfwWOmxZm3iIrary6WBIxPth
ND01XRGhICgpU+aonZiCzSD0drm88ZnDO0BcU8pC1lX66n4hO5sr+qHQhFCN
Qk8OnBsVcn2vZwwaAWGx2v+BdD02QzqzABtpRmc1D22lZp4A/OxdqJ8F7nhO
MpzyR2WdeF7HlKmL6LCK5pilVkzzuwuq9L5h0cmSkOZfBg9XiWxGFfP3N+17
KTL6CB2CtdQXt0voBmuGIYMCs/vb+XV5k9CISsK5D33SM15XrEjuPa5f0AqE
ZpObkUBpS1BshW6GwG0VGrpCUO+J1LdJF7P3z2Xa5yKhIPuIohBNTeOEiOG4
KI8G/8shZISaVoMFisGTKafJZix3+/WN1YvGFImzg2i8PAiZ1Jt9GU602ZOe
qSw16rhUC8+NAtkHSLBhTXeY9qpMYkJdMPbDlUu8yOvlSoc8uHjyRafPkgQG
mDCMEMkh+PnXuWn9oVlLCEBuB0CmIWONzf/xjCfTxQKRyWiqwAWYEdh1BRVM
61zUYbTJ37yYuiuyV6npcy0nKLLSYuJPA69tbV2lfOTg8xwo2mc6uNlVDYTi
Tbpog2C9DEQi4Sl7UMUwnNTCJEK0u1vjZS7/W4BgXZeLFrk53rDObZ6CXjpd
kSUrbo5+WWygdTLj8AViCU/wG4xnRvjl4tAOQOugjztE238iqQu9rmwWuasM
BrrVe18ITFMIEohd7IwEx0AjAWoOyTBSjF1sYtzUGulkRN+sj3ilgcaxWKLD
0xgH4F5ily1J46KToBpkVzSWBN0x48P8wZYMCwFSCj1AghtE6T/BU3bRqqL3
ppMtg5n2Uj6aH3rxxJew9le/0r6GJFNDSw+76n9+2h2rReBvSLbCq90Tz5xD
xT22CAWBeQ2SMsXwF/K0wzr1efh6SspftPp4YufNCI/NU4H2Idgsi28tENXS
qyfjeihNKW2fG84RLGxqcx8D/FGxM2mHm1hdgZv+POXGZQR73lQdY/IBg9ie
ax2Puwkr/MXDpLZqOwC4eajyFe0qE+U+2On9AGgtZq08L6oO52mItMKgtbGX
ok16kqZyOpNhHI5bpWX3/9uA+P88aqOrg2R7CHBk7PG1C1vBz18xeILX6Fia
zFdlNp0aFhhF5oncexpmFVQr+VYgWdO9aptbrvpqbN6eglxeukcydsIW8c+k
ejFgfIhqK8kIv0B4ejwY7akhihNZdyAKo9jBynKLajnwrX7fQC3hG6X8UZ6m
EfOTvrDTBp9Gix0E+1hs2AJj/SSZjeXXm7cOqmbK7ezfeQC9M+8OTkGxUhCl
aABqCsLk3OOFxAzXiXgkCMefVRRjb204buueDhHVzZp+n001mEuUCTAYjQCq
EaJ1vhkjE0VjLjlFbkjGxJE+dzD1ZT4BGevTDHuxN8Uzs8dVtVJOXNfru+ov
X0Z3rt7hovBDNvv5zrqblEbRaNCC8Mw2NYAU/HpXPlzmz4Se3f9NNtJQWN5m
hBydjiIWFSZNF4zF+o+CzecownDKvZRmTRl2uqR07x6G6QzMBilqyAGRr1FF
TS2MjI3RUY7oFlWIe1uezgvjd6ja61BAqAFAf4Qrc52yL3DHk3nmb8Map0DF
9ApjTmOSPcnTLbgCOAY1wN9O6k9NcAKatxylqJbR4/Tn9SEav2DwNc6FEP2S
KJvRONAjqx5S5yoihvoP6yC8ox+1LkYSB2Zb1i6t2MUzcpoOv1GRUB7vz2Am
hCR+raIoSX3u9v1zVQZuwhv4PxdFnoJ5EhJQcNxmOTy30uJLrlFVT3Dlypu6
NXxDjqCAWk+olSqIM0FrBvPmufvm86yjGkrDMsfGn+RwplRtE0/meNqYvWCe
LIuKvlEX4iHMu8mjV9M46OwP5pP4KsIM6+55NLXVW7QpcbYA+D/xDcYACCQ0
YrcZyUoCeARvZMeZV23WZdij9p7Y+FHDBC2PT5Jx6Rnm0iMJ4G/GoPfEc4QY
TJFEMiCoT4ffC+aMprpAhrJ8W/Jc1bCm2y0D0SGinvjxNbaFT/SC5x7l/Sbd
bV/NPpuVK/tSaS43oqS6DjqsZWX+WafxkommxY7Hvx4SQnWaDpcdDRzeZIT0
6SbPuZ0nNiOCz9q7YoOjXgUmz7HR5f7E4N+0+SBewZGCQsRcLGUpqHAY7nNn
EB2xt8Pu/CfVn0QFRxUdO39FqLjZlt3H+BYzRx64jrfV6tFrs/fOkjTIjLel
BemD4yBKDimJ+tm3WTwBkOXHol2aVrKNlCPbUvD+pSzbunj4/8SQ4AQiMC87
z6LxmnzO3pP/xaY6euD43zkmxPiJIAU8xHnhv94xjpTHDfLo+7WlnzOezBqr
LtR/DQdy8s6/5OV5LyE6E3JMBh2Jrx/v3W8QKothuqB2Pf1xwKk5B0qjHByf
0T7TrE5YdiU8xNU5VEE8Oa/Gfg+zgKL+5xpaQDoy91PgzLVBP8Jp3rXPdt44
b2d4wCYWgWoXyeM8Uj8AABUZS4AkzyQG0Bwj5DnzSBAVNMOqliWKFBYp6jy0
0HfrPJ3Ba/059d+OVgFHN+mKpVNf2/BWj8WIdt3ubMPjV9NONcab8E1SzPhc
Y+7w6bl9TcLzEcsaYcrrJ6LDZ3wrgDK8BKb3VIRG7laVFFvWBgod2t6oWZdz
KXnGsMb2Cmfl1h0NYkrSTYmLK7LGwbvdHQFQVA7DYwz6MZSNx/B9yq1zJLcw
C+Rew4R8C00RutJNS7FfObitOve88KhQ5CCvullj0qhcFDSxUILv06QFimsV
5tqAdMKajU21GB5ivmGVp4yUklG/YKIUAuDa/bhpjhQv93iQdCxszabHzXd5
oiDUmb31WBpNrwb30lod6tZvomLPWJVWFXUXJSFPPYhO2LiBIsk1Aw2DtvgH
ZQp8bikMHiMdafwRq6pdHnsw974AiLGq18C7aEpF74XsQEzoYv1+8is5F25S
eU0YijzdRawjnRyOVOn3fsYe8iJ6C+U+PYvjwyy7wfb/V+M63esgNxrqTBTD
7jnbcjcdwdNWOVa4tJGpja1W8k3z1GKJQpQOiizbQ1e8UHRCccsZ3XSrMBAh
Q0kDySsvoe7BX04eOd/N85BWZwth9saUwIuClEcPzrpAh3jD0/UrQR0MtEtK
I/VHOwGt1tSdb/6yUNMU9PWK+fDw8cNTHKvleCBYQhH//Q0vsfp3WT1Z86on
MCcpFJf/sJbSE+gisW7SIOB+UfH9sD8lA/IL5yzi+iO35xFaexV+ioiT5khj
7uFE2TQGCcwKhCPVLuWZahirhgGOw8nM2/0flc0qz3E0/3Vbhl2huwkBQQGT
2enOix+/4y83EvMU0K8RN3rlFvnbxDJZzgIBu/pM94jqcjKlDvmWnlUJBlyp
DUHfvTpG9+mlF7QWeaHWSY3vN7Dan0vDOCNQZLOeaQztcP8eQFeh1/E6meDq
EIoD1juN9xTveKjca01idXi9jiuIEEbUYi/QDf3hWuy1wIRFepOQjUloeMp/
MD/+LubbNDkEiAQ0HydirJW/a/Mip8eEF4eAEpUTKYuoOTTapJVIEL0FjCX1
6+IR23woxCKChDqCtQnUm+k5yvfVt280pXfKoV5mBiHaSEm3MJOCMhcq8S5N
DoPxSv/OB38fVdc0By6jUzcD6DWjC6CwWWTeHTyN0Ue/+bLNjgdjLJmt9QMl
J6V8jfvCY7Mg/L3aIjOWX51LztRq7wowzEdp50fwpeeQ939u/rAZW/kIKIsJ
kHWgxT1E0DUt9dRQ7vP+DmtENEBHIicjGOYaoMu9jEduGbV3wuJZ7yg949+T
KHv1MrkvsUNtNKwNEoy8Y0GWyRHD4RS2Pu3L8+qMej94Fl3iorZmNdqWhiaf
9+bXnAmNNgCUjSaMtXD6U5JJlF2VvC+sbSsQem7SjN4JHpTNFhjHS5b5ZTmW
PDKV56fufkIgYf1u2uajpQ1pawo0mHkskYu+DlP72Q8UgA6W32v3VP/A4jth
0e1+XEwLyD7AKFW9vKxV/h+ck7Dp0S/OApYJjIgwtfaUS+17Cyry64EgE6bj
HcHSjgTPH6HqbjbztwahBCfq1iyd3EJ+c1MZw8C/maZ3wAeTQ1akp7cVycAo
/53ws9JlxcE86MZUl/eoeEhlTM+QhpGEBCN3prfc/kAJrPmrBiuD92BdmnDv
dS4CUHGCv1nUqZ8ucoh1NwwuTGfQlXbab0+CQ5owyD7+nnT1z2fuQtWTb9+C
ZSTi47mdhSwbrrLPQQiLFR+rI+lOcCZ7ukDhnv2xoxJUo3M6OitTYwQ30e2c
qrvxfNPnmPVCZ6pL5GR006s+NMvZeoaRF/mKhssIhfVBrXozxpB4xfcz3pVX
qW1IfOULDk1EWzv12mFR5YZCs6Qr6ST0HhiCi2yWeFBv2Moov457KpDBBVcj
ES8Bf7ekHMLGQCKo4Pe3GGxIpnY+B5PeMXwOM1GSvzJEOr+oQcwVkW2W8vq5
0XQCbKZTgKRwXlmaUrXXN7T32Q5qDGwKwoAGa8IQolpEK1SSZx+3KhF5ap91
w54UeVYUysyPEVaZn216yLPZj2RJLQebBdC5+ORwto4bWGTkWBpEuHj+voeh
Q/vIXoiXHsap4Z62idxsK5SuTjTfOCPD3VYEEs3miNEPJ8zgJezla8hjG2E+
1JxkmBmHBcxbyEJYAloy8nzll9do78qGtCvYr4gLi4Ih/RVNKGYNxLukjBd+
l7rqpvPQIsTGSFUx1b8dMbBxpeOlI5/AFav/BnQ9UmH4P9bS+T352Hk5kbw1
WzRBZrheq8O7ttdDXX2d/NKO47yP6A0JexYLnTAq0zHbniGiqfR2RUlwykL1
FXH3FQYRav/PYewKaMoXTi2phxmbEMuv1igBSZsut2QNe/PUWPl6ARu6aZ0U
g+jW9PGTsqXjquKY55k3Cx1LjBFbDBeCMzPhvGlLPR3jeUrjyp1n/mGQ2dTP
KM2QybeFkoikTF4HuJesRWChd83y5KckRkrr41Hz+Dzw4EYceQBFVUGHD/cx
RYmIYFqK98AA9nUPDaYvky7tsp7o2xG9DkSEV0pP+X1Tkf0NHZbyVIC7SVes
Cl163ZkHg/itu8nbaSLsBCZwTniaVpMTorDLNZaCjCPGwl1ZfZTtJJpt4BJH
1TGO00D60GE11wC410uGu3m/lbmuCI0t6+dArWq4D5n4oeFPhhL2gtg69S3G
xQ7PW/nijYDU/Uk1EoEI8JAyEwSyAhexkDiKcbvDXS09Y09Vaf5PY4OZ7c3u
5cdTjCdaQwJN7ibaDGpRnlQZ5O++AsNNQAX2yGL464HfBRFMPjOCstoXInnt
+Ffp/TySGBtmeYdYR+/v8KPtNkbBFADapyfdIQ0T93FFb6jqFudARuf2yaNC
MAifL5/SP/VA42snHD9h2ZvDgt3gJs5xd7h2IOHgubi2xdJ4xDbLVdRVjxEY
Go7PtRptGwV3PJ7+xtQXesPsbiudrKReNx8Co/oo7U6RKUM5PZasnhucXDcw
tvQLcTjpbGPCGhrYDtLu3RyT7+7qPabzLS2uLMwjxEUTTVhPXcwvmTUQIy1D
nU4PTg/J3Yb3+urNrWCNYA08uiwXGqRt2eTUoHglWKMJjluJdA5CHiAEoHI5
jtdmqJiSv7cuqUmMx12VBCpzspC2xm9QYP9GeEgpUoXnUFA9Sx8VJ1oHFw5W
dJRvod3/pidDNt08/hPH1XoQBlduiFrfoyFtOvvxx3+PoMOine2bQ6tZkM67
a/FhrwRZGVxPfTY7fFKK8eb5yqEv32JM/1dyrGayFJaP+nM1wDy7yO2zQnzQ
yXtF/OCqQm/yPqn1xxriFiwE0TB79MRa0BiXYSrWkrJszs5+jnWG4mhmG0cl
lRFdq+u6+XymFNWdSrwFWphoI07FGIlkX7I1yhS0Xrw+zzEhtTV1VF5Rgo9S
LZez9ajgE4OzuScndKS3UO5AnGUN+SqnuRQFSEUCs2abAcXaa/Yfri3Zoq45
D2k5JlpY6NXUQzhRMaV8NFFQfCqYmz6ikghuR3wYTDuGMn9v280TrpPcRx3X
Mz5agj54TCmSOIFDGGidwb9VMj5kzT/mmZH0oim1s8hhQpEDhYeLvzUIXvfn
Mcp5BvfR5ZK/Oxy1x0AI4TU+Wh8VJxp7XcH2kSt9wLN9xLXnDcFG+BxApv7H
c8CTPLCgbdOMQBkBxF27TtkpSGvAkouZ46L0c4f7W/pwKcyOaPpv5tHPkZxg
2VKC4aue/0XCTwIiP8gtqNxwz39D+KEGXgX5+YNeV8OBnOMFLcCwkp1wsOiq
J1huYTkAEV3G18Mz8NuGbWu8mMAR5IMDyAR9ePex1Wp2wv2rlsP4HIpTZ3XP
e9lMRmS6vs5ymVhx4NuQd5fA993+w+maTyTSVCjOlmHIIIQQ6NQ5C1uQmjM0
iLX7j0VYpnJ45JFLXmTf+HRSgDt7WnXPIEtXHth3xbPt1xmIdfGcc5kO+FYs
AxbCnXu6dNCEw6Y0mrgn5eEt8suBeRcNssVF0MTtZvNR2rdiRAMHr/OOhaE9
jk2J4HvPU4lexBeba9rwqqxP7y057qZZnhVgdrJyCA0zN6qiBcydFZWXyjk+
3BpyOhLvSaGgACJPrlyEabJeQEaZpm8x3v1OyhL+2voIvMXT9cW3LJ+7REKa
Egf9XmH84GWVPaYZMyS2GwPpRogb9xXpzoXOZNzTOYq+Q6nx17k7sbbo2qfT
1UT6SyDT4rqF5CX5pWSdJiCh9rlPYJVMYelhK/NrWfzG8IH06S7xgsfxpoGF
dFWX4Z75jN5CXOiavo+4o1Fr08HBDAkc/M5eCMJeW1U2fLgiejR8U0m1utsg
dJN87OGgNJiu74NDGaVOBlGoPjM+QlOf9Gklv/EeydfNRiH398pfnLYWwxiR
nKSD3u3nqYN1mGjzP83dPWMXbEERpLWcUePrqIY1sUtUWNTMLw/bmNhZCHt/
eMkUS7PWsxjfNZI0ZZkItGnYQpzyBIK3V5X4DjDdQ9WHfWi7kVumCQdSaSZV
f87xhPCmgB9w/rfDOWAc8npSMyCJ6SxFhQ6a/qqIPq866OVcmSUEdGgJDP4Q
qoQ9b8iZt6Dp/t2AKDL9NyuWT8r82zpyq+2Rgz4sIVrq+G5r5tYOWrigs4uA
QbtuYXLo+alQoVLi2vG6tYkB09U85UXN0PNJLC+Dy7eB7guULnC9dqXXFNTo
e5D42kWz4yAyIDBpfLAjNuAvjmouS4MA9dVYGHIcWJ84DGq4vtmAkh6o2TKY
Hd9n1wtnudnOq+yJnxp950AYu7Dc5fakGK23oHWuQgLivbsHfM7kaOI7Vubn
vz4WHCdpG29nhGjgmZREMW5usIcX92307vVKLWk208mVTvDnsniiHFrGa2yo
GUNqrcgpZyk/DhiikJMrnGd5KMKM5vGeox/YDu41z+hvaSWXSrzNu5Y5h0fu
W6PZxxpCT/9pIVLFzWKkNjjRqhxxeX0UJLnwK0iyIxu8D+bJCAKFyuLEZO/2
su9K38wxjw2P21TkdLtRQiHB9HgoFw6fkj7FXN/caEvpITmMHk3rk04iRxae
bCjbotVVpoRVirVriNpzPaHAPBqaewjZ6ykUjivkmTz0vM37uSgDnUQiSkxd
xZGymZ6Nn3ElYr4zl6lgDkheo3KGXLJ9YyppLuImeP+IXp7rdm7FmmaQYtYL
HwiZ2zRW6khj+o2iHybeeZbDaIAfygJICbx3z65AY9OqeOD0uw+r+NPwSz4i
jI696s2Kd6FX+9P/rnN075DqUU2UVhrmAyfraPTCvYyFl38mOqspyVoJ4Q83
imsIXU73G7/pGaG/5mTMHHW37K6eNMDH82nFwFg1+weAL4X2AsFphmtCWyN7
34/UiupV2xLE4enWvq75JNwaCqBBQBfdKwzpls7PARXwwI7sAVMF3rcy8bQ1
4HLEdK20GqwiqGFIz3AaQvsHPL8epZn7XMwf7gOZrjxpeM1eMr+Kpb0967m/
D+kCN0N8MivTiir7J6XQ6VfXScMkxfSdQAOPS4kVxMt65105FeSAyX1V+DGJ
oqsk/Q4tTM0CMYnYWY4IxDQ9Rd4LGOfYfiAozBKzGVy7AK0RNG5wGVuFNOZ/
Dw/MwNE3mUL3wbJS1F6zPJSTlwywi9Kjer4vSaTsS510WGRo1qgTtp8Uz5ju
rfOCssm7OIF/sxTZjRcFMg2HZjDg7rdDJM9TVDyFlxGNzeTayyZhKQroyHuv
iEVUQEGKexDEonc1B6b95FQfIFA19iNHjlnTwlK8RuYyGvM4nED03JA76ux1
7kkKCGI8qs83HHBxLptNlxRLYIorDO7Lss2ROCnmCkFJNy6s6ebiQKODJoZo
h0M8H53025Q2DV7jar1bNbfmdHLZ+n0zzDTiSqRORVDdw2JYn9nCXQZaIhT5
an0CCmOkrLzbjg1t2AQiIxUk4Pq8scp29iG1PZvxnCjMThZUC/atGVaYzWuE
2146iP7pfjQZ3LWlup6z5aYuNiZoR6ZLllYTQ0Dce2v7pSiS/2LBxye9rSXn
2lUg8zbgk77hbl8LpN8aEDxCk8Yhe++ULvCsCvWTZd0fCg32ypO67wFxiaA0
d6tfMRGMcLUfNv7FCEKSERMVN6aWSS8P7VDSYNB9VcGVrPPsQ/wQGDOG7Zit
bL84zehN4jMRHdeo1c0xGE42RiWoT/qO9v2V5Gu3QpFVsCqOvGPom8VOPPeY
zUhelhoiSq5FVbIJxge/fHZTrUQjPllr4Sv+3flezd5I5QEki97cuPjmJFP7
vFzfr7+QzITGQpD+7PPoGFGz8q/Fv0pLwVJJAzu7c9JizZtviWrnSA5Yq+H3
uhlROeC9+CC5An97FJ7DjRRTsowiIghpvmOCsNuFm6vMVxEmrWWGjwHmkD95
KqJpNeM7KFYrmwwiowJcqLnzAyEuCIC39Zk8AfAHGqkgdS3jhuwm742KXL4M
p2uTnq7JwGTJWLQ6Rb/PmPvWYLAinILaCpgHZeMWljSx+11K2tkeItbfSoqC
t3SCk2+2HUPVgm9izhPznSAgs5xWJGFtELTitCGPix3L3R4lu39h92V1J4Ji
3lggjgNdw/LHwwEp6DG6PMImUo1EOghxY5VME0F6bKd5tVyOSAbKbm6SFB4h
kysY2M/WsDXVlUC/DYVA8iNI/Cw2Ne1h5sBW2e8mHcWmqgA0vHJ1PJTzHE71
A28iN089knI3gfyuZ3UlcEkX3oJypE2Ig8VUvRTGNcsE+vMkt2FiQoLobowD
t7mAJUKU0ZufIAmePT7uNnRQEIl9/RygHeguCOokCe+8JYB35EAgqpYGKHaE
/bOqexPR/wICF8zDJRp7bW2yTBbqMKWDXsmzokzt/T5i49WJrsvlevI2UTiV
l+iK6hA8bB9Nz3mdrecZ/k2A+Rur2utinKJFvA1OOH05twf7mYA9aP/sGCDd
foOJRWp/3pPZf7nlQv6OYf2dzGvUk2sThqXZ2XmMJa5ZibDmmQGE95AvyTPj
6Xlv7gaT6hEPSHBooocVEsUCKEuvx4D5oJ7ZXOh8bjQzhvwA0X6zdDWCRtMY
8F9T7tVCjhxglCdhR3kh8QstAVakJKC5Ch/6OR3G/mg65ApwRY/CxQECHIcN
0/WnXyOPYIbSnGOOEI52GP/eNWIs8uBkqIj2XBJIZDGyZG3FFCYKiNuM3d3o
FmgaaFt6aT5Ou019D9Vmxn4Kj5Ud3drCVKR9xFJsiuLpgG55v5bPNnLTmsuS
ToiviljRCOjdBZft/sNSbCrqJ3v3kcbaQA3J+kxnU3OUWZeQqMsopeRBcQhq
/bkkJ91tAZLE0qmEygS63EqcQvyFh9qqgzHyOza8brxOiMROH8uqx4l8ug30
rCCXu5C83SrDnvBspqaoECXeIbyp8E7RnM7q+EYo/m/Z/snFDbB4eevMtTfy
bLanN3F9yMKe3MMQT1Li79G2qp0tqnk2LKt+ZlOV3HoIzo9FbsfDyPEBTd+J
sl2zsS/beMzDHbGR/kWC2sX10AlGxOk5rHKN85lndPO/eY+HElvkFIPBxVkf
aHtysg21wZ8ymmKokwZk+dXLQWqcvrF+Vi+3HVtV8fuxtfC3hbsRyhzn9fPR
mlLSGJ7oko66gNqYM2rU6WbKZsb9ke9fyuZuxH4JHr5j9HxBlZ8XIJ88VPfN
yrciHnbtdJ04dyKgJf4yeMCbPhhlylGnLEiDafHfrthxZVB0I3Saz+h2MjlL
YtyEYNeCUg7tchQtxLu3hgdwSTwEGxigQdxOoed3hycrwvXu8itiU+0JtZ0a
JVn7pgt53/EAMMIm0pZdjTH0beybm1nwcIYLegwbEWol/+HQzx/e0Y/XGbBI
KjiuvBdIpIwbCkuTK5hGH3PpQ9loFq6mzmk/kLbl3Br3QBB2d7ni9mjlt9WN
b/VYclW77zGaeyJrg+21b/LnF5nlVlOumCEpFRRgY5h0X+MliUKWQv/LjYUp
Dmhd1ZkH52J9hJmpoqIywt2xrdEoVGKRxHEq/Cx1msgIa7rDl7v/tDxhsICl
EPuWHt7ewnz3LGDSKtlqKMdNYeNCPDbOBGbxqlz9eZDalbrJ7BaQhXbf0vKW
MdFXJCVu5/pW/pqTGoNo+R2oj9F2XycrxRnAjGfkxd4Fki1p+lHB8PubZa3Y
FPIueEpovNdQ9R/Dk9gxFJqjGwrjhwZs6mSmiqasSrSOpKnl/gkrI0lmXhpB
ablBH4AsVHTXW60sAc+nhEDCymbSqNEK+Mmcwcs5sG7cOvvrAKvdFiSVwmDI
nttuRjLmLu0htJXarq+0Op8/5r4dZTq/hymhDhSPFJdDoIMgdsfiZ2p71Q90
Zbpb4FDSlPEGqNCxVKr4DRjWNDufr4uhjNwYS9Kt14fJ/2q2YZf/u2l07Ogo
hwrx17lC4JsjZGoT0jDtEYIXboySGsl3nhYozc5wJHx+ZEa8ppW6Z86kdZFG
VAicXTNhXELGjCEhMjTQ5ym8cMKNnb20S5kX6tpN9A1I8KnoWDM4QW0TUQLR
FH6yFvhuclPniAkB4JiZwrz9FX+AfHH1oYKztb3rH+DuUy9R1/Zg8C4UxQgz
jO1UtrlHAA/Hg3/WdzataCaFHpm2fsy+GShqtDsEyWQ0l13tAaMp/4dpdfA1
R87YroNcI36fz+LMSa1LHDrPlZYHnOgWpKKqm/HzHSI/AdDndUWDMMi/ol0y
V3MsOJDAi3gop3Bkomyycy9y0fnsBKzxW6SslapeXPytOF5ow/qu8JXWZ3kM
1o6SSFN4IIxcDSY6M6mkSwSmAT5kdX1Wv5t4kTmKS2V8vWr2rAxSlOoWPAxa
hVLrNzntT67/jCT6awx+PGA5Rb4vYfK8V2W+zyo26f2btHvpfxcYHfnZT4yc
LmnP5Grc+WYyvdRnjZyPiu6k7cNcxDhJ2aZa394izEgOibmKfstwiGydvNrG
h1thyUgbX5xj0+nOAyYyMGTmr+oXmYr1CcPIZHcm2GKdgML2/h8Aovo2oJVV
NtSCDPQ44w82VLAJViF/qsut0ndR5+WRTvWBzWQv10/drkHAribKNVJgvNIe
pazWXysnULIJbPF/lIItDZocwSw4uGc5GMjTuKSh4It3dBonSA+uqU7APrNv
r086NE9uYe/rikYI82ZeoyaigVyECrB3V3QwA46GS5WA7lubQ7xhB3WJtZ5d
Ks8do+UlR7kpOGN/XmP0gkoBR+O33S6WkAN/VVKF1HqxeHradCXPjrLQyG59
ISH26AOIWRntc9YcvfjEx044b3AamawTxQZ4smSUkzD8wMNrIwBRgc9/C53J
pkdbWmS5YlxqQN1nASrW9iM2R32a5ZKW+GdWsTnj7SxegVumWdTNjU0UJrmI
/dFW8cNWg6z0hNYCEIEtWZxeGY9gWOrIz5DbLxiDEhDLdYm5YyPmtEHBL3Dn
B8TXVaX5SUBoLalvEIziQ0MYMeyRp00FXs/PfgWO2fJ1CkBwFsDTPUsoYWnA
09LyGRUJ4ZGT4uvlVGJZxt7cSwVDcYiITG4F5DAropxs5GPiO8EoVvhdysgb
7cZpt6DSVwCwvpP68FwPmsHMRMxGQh8KKcRVJyBiyztVpg1TALqQDcXNDW8d
t0xX3ON1IcYokIF2m2mgceoTewkFFnZMgEqNcR590Kj1Synkiuhk+SDINyLh
S7tA1bdEmAwfILzl9Ra6zD6nx8yAsE6gtVWljdxJkDviLrWgSrWDxObqMxVy
EZDvaLivcfimtWBsy3l83e6RxY4O1rE70XquktyKbHciLLcIafwcAlKJhZtM
vo+uhg/TAOlf8h+EZF0Cu3m5aEdlWzRGK56n1I0g910u+YvdDwOHM0f5Al+X
k7KySyI9OoFJlmQ6uVPXVrS552fRD8pY7UP0tpd6xm+yRu3IGArFoBIBpLyq
klf15HkEaU1zHGidtbXcwi6zNFzp7MGmtR/4kDAy6dkhbQeV63/AAGq0i6rK
PxjwrYFPqg0/ySWb6FdbDPA6559//JDz1C8WBoEAo/lmMPrywMc9d48RYwRC
NHS473zTQNr2ue2VGKTim+RGS9N8ontN9Usn4yzOHpuEpk5cp8eZvQsPTn+6
y3bltXxCDUgwsVmd2MwOEUSAsQV465hT+sFiiS8y4vblE7OyjJT6YxCekbqC
cP3A8Ugs0qvPixA+mPJH3UWmh7IY51e+iWkmjA4B9aXMKVer2vwAk+Qow/z+
6r6FsADMBGL5zCyR9NeQWYHU/OqhEpPWtuNx2k98YVRYzcO0BHA7KWg0rdNM
rPrQNux1K/HrsSCrfyAWYUUyA8VXUSRkSKi9datXAU9despLAilQ528q/ppx
AmSs0BadHS6v40aml/sNZO7w776Wf4EXB0pD2ZXpvBfuK5Gx2cvypgIedtv6
93GhXWfYZFKLmWi13igMZe6NTSwelGY8/5r6PhNuW9/sufLiVDcIlVnXD6Q+
Rygq3zetvONKad9y4buZflI2puwC3gIiMyHwYXdOY9zDE3moClMTKD/nGgMD
k4Rgqv1pe5AxobyS9xPGl/SuYC1oldNiBKpR2JjwlQoAYZACwFBqr1wQkI0P
12s14oODgZ12PX/RA9SvJm635wphYEUPARPiu6MFitM1eqCCkDDpWSyMIKOx
18tBE04LsLdZMZAC9uvrRmEFPHV7VoiRGja1rKbQ96xS6PpaKK6UUOU0EIpi
Fya1hYHEKtaUPPQPtkBKeIgNGs4agZL8uP3rQ1AX6bDDQfZo+HmmybAulTtd
/wvhJOrXSOwLuW78KVaKT+ErvbFWXhlGpybeOcbrqW9raW28ucsru0jHs3P9
JU28Y8E4b6+Gx4XQyGFBqGv7tqGmSMV20E6gVSABUGTh4ovC2C7I/+SqZ4bF
SKy5uBFyvLdA5qYbleGjVZVqtT7fYQ3aChF7yz07Ptxq1MI/xyguL/px2sag
s9VkqmZKjatFpLb/RPxFVIjhQnDL5/NF7hRDHyxHAGzU+PeficRz5nzG6esH
8e/5oZ3Qm/GmWfKFZDp4a8zGBYU4k2SNczoudtEg2waOk3J0u+XK8BkbhPGC
RmS4OpNpHjrNjDpmwU6LFsFcrGF/kotzk5V4YqE5Ga5XTOBvaXK1cYb7/2Ok
0RtzT+mgiHfQ2/d+lqiyNgiV38bszrv8/Y3m8W3gTxzKcLISk2aNDehzDVno
rtpWhhBu6WVnQS5pr3pHYrdH01YptvaLFswfZube1LN4iiBOzl0LLHFph6Yr
iVHi98c5lazlWEFHWylW4yXi5/34xIDFTiSKi78fRdszSqQV/s0ARcV/RASC
qMdpeQqUSe8QJrb931H9cHVFn9WJwRICYcSv9ZrW6Y5RCHhb+WZsVScRn4Xn
6w5bbsFTKlv0RlLbSBOTqmRODPoNuQxvuABemFJz3PrY9Vi2RVd66apgXiFb
zRf6wCkLVzrV1qoRyT89Fug3lfuXZlyv0LMQyF1nMXVlxIshicTXpsyT2ptv
WW/yfKCdWGR4g+2Urj68XY7lmyAI6z3eH/KD3ewCl4Yzn+8pmyeUoYrEpwan
fF6c6bSpFDW/pL383HqUkpumpJxrjK94V/wGqQMGVxe1DXopoX/Bt9shJtR1
crP20PxAheMLG5BFVlXjGU+BTmyAOX6I9yvYegtMGnT1FB4/nPQ4eaM8iL+g
JV1Er9G4B8dmmmoHnNjQva3fbWHOIHb9n6lw0AdjXmNk1SMTzCqlbtSbg2st
Inmh4aPvZsMt5QkOcMUEVCDVsvmmIYWm+JYkd6Nv8a5uzGRDEXHxMeCY+MZI
d1/V37E5rdsPMcGKkeV//2VcJvN4I8DNOumif4mmfe9qbo0IwJ+NKDUBjU0/
/O5kSAv0AswK7zvJCYb9zJBkeDQPILbtmR/rM/ztr8ouYUUNJmq3UGfG/Sbp
wLUWGGjSk2JXLB0uE6tzAU49DtruFA9OBXYQArXvBXPG+G2KSwFFta1LAz90
INs9XMlj5VgeyVmlroeHg/8oPg8FqHllfkNvpFK0g83i1PL8//+lFZ+OCMg9
G8+bqum3dJffzI87bY7DXJiL6aNAeuwOxzTK7FNgWQlh77rQIiD2uQ4MFF0U
iXTOWVGhJ/Df6lsN7m3rGnt/+JrSzUVusN9HDH7P7awb7TyGs5+HMq54D8L2
zsndgtjaX2CZ26efRCfIB1ImNN6LB7F7n9BEzQegriH+x34j1JKhfkOlfb/+
t5Zm/DbRHBIqfN5++ZACZJ9cQCMo0fYcwwsXTFk0x4Dyjjb4KmUsy5IHsS5f
O5hjjbZTWyc5XefoEL0jN0TCWjwgwjyvJApQrTuU7bB9UZHJw8URkqadRJ9a
pzM9AbPrpFT/BpXcq8SzCBpsNTjJMWT+C72+HTfKL4dXYMDE6YJNP1+MEprZ
oazPSOZy604xCxSdlvj3bOC9yjq5dwkQeACqvnXwZBa+ykRY7koMDzanEoR2
Pku+XjYKzWN1tgpp6pyk9EVnq9QvE40U238c5JTknecsUfQjkwUCZAj/Zqr9
0A9EcnUj9sm91f3Fys9XTYuM/nB0C3h4g1iIj1kyWRk8pYCqx1ebho8SV3JY
vBrr3UN50/7QgY67LyLE+jB97JOzvMv7NCPDuBxy3hOnaIYbV1W0nVYeAiOv
vNJPbh/W7Tk/r5PASVdePm8zwjPaesO+34oftBwApYMMNK6fxqy5F4PPPW5g
C1GZrnSULPYOb7Xq+gZF7rvhhA2pcfIH4tTFxsRLZigM+fpvylrO/rvLFTLg
aMxZXk3sIIRYvZKZqnSrCAPzlXsh6FqXK4rL12B/1j/qv0bWbey0IgnwEfCM
KIbDqa3kCE03Z3TSd+W2J/BBe0Z6g4TCwO8M+3rnZW2182xukzyJlIMW1SML
uWE0hC4mgca5zL0M6489zi3izm0FmDZFQWYUHGGGAvV/fWYge3tVaUnmfp6L
NKkZQAFKJTJJIvTsQ5ivIoIfNK8q/5bypPC+cAD49DPF1zffj5/qP9EXaNqO
UEn/BiAJMr8uhkROX5jXOiHosAUj5CWlQBnxwpcHTA/ws+b4CxGZD9mMDebx
m4SkoBfFeeTd+i79tq6hdFu9qZXc5FDX0U3yhJz7vqS3SNWWphBuAxMzSyAd
DKuU+5M8ICGvNZRUEU6Hxa6RkEdWT33sDGwhDhwF8q8GSZ70vdEPO66w6X0z
0ODLOpcX2MAilGcGujdDZdgaBusimyrAcit8ijY9fx2nA6r5/kNkCoj/pPwJ
Ei2VeeGMvFOFe79yp8PKrNIHKuUlxeySr98EUthI4L9ApPCOhAgW59ZNxicF
Th+Ro7bJdW7NbcLrQT/QBXv2yEyiNZzG5Wj73Q9fr5+gWuHby5TL3DSZix5T
X0DuVavPMIHniMGArcMe6Y7lPPh9EROfvRE1kkVDJec7Q9f5kPYgWgwf2ubH
83HkLcTczm6mvFxm5an2hjEyDhq5VWso3NEfpFciRvlH2GdjXFRBofDFLpA6
sr1oF0DcInMQrHjNO2JhuqQrC5HDtqu5gLUc0T1tasSNH9nUsA8q+6wZAxll
a+V7t0ewgVwgEtQsBfv4KPGXZp1Mse5jJLbnjmRgxt54ISKdKdnw9vprUB2J
pNp2TKDkiTDy/6YVd7KdReBKK+d2aI+iUo9hzVZggMnzba1jh0UMTYxmGVy9
co0O0OhmLjYw3idJfH9wGYTMw4DNSb3t2Fno3Tve1nXwmvDdemDF7mSF0tZK
uDBWq4EXYwa93X3RdJT26K1HBKBnVJ+4dNR0iXgSj+Gpy0/M+gKaj8a7+X+N
NCCXB1doecmg/TGzLQOrgP3BPAn4DZpG3puVG+1kEzsdPr6BC0M6DOQ8Umzo
t4oBk+lcjNOjiJzFmhzn5XRcL4teHgNFDF0AQQGX18huWU5F8rt530783/G9
ZFC4XicmgG/n88eHn7EmcNUTFc+Pkj9EIIMNMt3YEnR05A9c/HwNuZOXrQyQ
+Dg18xboMKdz/RDS0AiE8vpcrICu8S07PYaNHr7Z6fFvyLY38PJWpt5ZHtli
jzwK2X8doht0hRRw07d+9ymrg/6xsxaBWGFPISFeh0/TuwVNWoKoTQUULu+s
gy+xOz8unMxpyfQQntPMBNZO0h0YV9UQvWN9Nx07Uf9Ju4pTcjfTBI7ThG6b
ymBzosOPbDfi8bMawvVZZawwalOyUF8kMOw3ErhJxMlVsB5CK//0G5w2pdJa
exW9oOtNTL5zN6mAL+S3FGTNPzd9NAYAUGBDIN3sGTwvEOfxzDgcu94k1DyW
lFidIzen5adsncttQZDPK8wwztSfyUd3TUBlVstB9FN22L1RV5xE7BM4NoBb
wGdaxeystsLeo8SKgnpy1qP7m0o7fv3ANIhB0NO1HkmwMALpSRD5UxYTmJCG
XMU/VH8DIrcnv26FAIQ7yxhCE1gs3Dhyn2pcMsET+PNdpx5N3KZLwXj+YANQ
6AzMt3Yj5naGTFIo0HV90H6UyUjaj+xQn9K+n2/g4Y+tLvfsuWfgcxvJ784A
L5YTt2mckL+NU7d/X4QZ1rmbw93Zk8FOlgcEGsZ8eq6TI9gZEtAy+9w94Kx0
Z9LkQQw8MNSvh6t6bnEInpfQeevz7FBJWXyWlOnSXRKUy5srH6lwPfdhEbWS
OXn2sKFqghMCEpLeyJROUTlW4BAxvSzYh+LFZ3MwHSqNvUJUBmaZbdok4tKj
gAGPJ0J00cof7mT17PF23I/9VN70r35BgHwVVFm0bodiaPkvdzNYYjar9XvO
hbYcwU7QshKNKea1j1sx5KrwSQQ6qOWy/cm1LZoqvNdxo8MLWbTKEhmy1Lx/
bsRQaHyhefYu6jrtUcUlrvVzcqPx8Lms9SW7wnde5IZWaQnNy22tY0yrrAuy
wsdnQeLrz6+HXXoEZTi4tXFGDx2ykXG0KiadXAMEySlJt1td21D5bZFltamz
ScpHvusTdJrBiD76KlvMiKNJ/DLHYUiAHs4ezPUXRz24Z2SPVJKP6Al540XN
NCi16mOkPV+9M1n/m1fvut+qQAOM3jX7iPTs7cqFRYXe02I5SG22/uBGiiJ+
LHnxrU8bb8awzR8Dorww8/S9XYLTybeLlKPh76gfXxwIFB/rv1Lc1/Hnxi+7
t5bjr6HW0gHHM0DpIjSJeLZfKT0ibn8PkKw2GfYHypGlLM4NfJawDUzfaCPx
LbZt3/54WMZ4u3jUe2Bw925piHmU+nUrk7OrndkAOg+POZYWAjqYM8t/j4Pf
I8ArRt14aT4jhECMDl5JL6y7E5NjrROyxgT0CHhYlXdRjusnrU+rAsYBsO7f
Addzx1Po/vUsGzI4o2Br7DZLOsa22nXqpfMFx/oN6bEFHAx5niAnR9nKEre0
IwV7cObuAun3TE/qR5WqyhtYsDwYc6dEiv/2dcyNJqmJ6PDPOI7g6dug8e4v
iXmAmgZnWCIO/G1vfBeRImo07xBG2yYhOTUXgxmuERHmA2mpqIgVL6n7f1Iz
gkL3vLNtywFRmVP2K8cEnwPzQITph7/wO23/IQmpJjxXfGTxmehWR+o2ozoJ
jy64xmvC+Gr0Ma6dR4G86SUbbCg4aWrH2jcRwOx0mCs0Lfz3Q+Dq/x+5JXOE
eoTngV6V2lKUII0TbotZlPCAXZja5jsnGRaD0inyW6YIYk5GK8OF8hlFhZQ9
dUKNxFI4Bzw/uDudevQGdcN4eJCg5uM5KFKppUshoKGhPc5DQw/T36ey/cuh
yAWOyF2OU6qYoHDv40tHTj81YppXqFxi+x5BiDNan3yr1bzSjxR0AFVOPGpx
i4EO9BizuSoqK2CQHs0lMjuA0rK7MMUeEdl+mUnqFdqK2t1VdB+sh0fqEv6r
nbvji+IX9usP2UhB2NtBEVCvew3hU0a9ADouMsAXtjLPTm2zfzcl2Et4zG4E
8q0Z1P/+fsDMLgcACLNzVslG44USTX86IrqFX35/A+JgX4ehrvaObl7EWEcp
lqDGH5vo9IIz+To16Bt2PqqDHE66MzrlNL0I43uGpTPzIUKY2tI4MdUQmLjQ
tgPauWtKnT7GSMTX7v0kjgNoe7XZE8UJ5G15rMTd8YmchkfLdgJKg1eHyFLS
mMtG9VSqlxLwzkLUZo4adGah5YrseZnXD/vdDJdJSkDrjYhs/DHDfqVF9xB3
RMBokR0bUilMH4pyR3hv/+y8jrs6edC17024n14MFad0zhy/CIuBrfqqBsUv
L/RDo6XEa94uRac8t1YrCZuqY/buGE5etTNabvkPOOpS+Wn4lCNrVU4DIKxk
iqsaRiTXIcWqyP2mPOsV9oALMJSrP/e0ieD7K6ilEUogqpiy+DN2WUlfENbB
U/OnlqLNE8i/42RvKkOfpXneFHR3uIdl3wroWICZzsePIrOIs4jZsOCQC2pa
8JHR50vA3ouYRK9fRQ6eUFKK7P3dPaSyqnWjnUpGlz91KnDqOl6YNG2SwyGE
NuQn+Gujr/XJmzh4zhCMFVundSLg/5Gl49hddDG9ZKMALD/jS4OAtUgbyV51
6/fVUVpPLwmaofBL0aK0w/T7cqoBAkDsMRkNHbkEPC4DGMgML0UpEBhtEthM
hZdZX/hcZxeydl6h+110pFXFwa7Yw47menqocYQEkCyQRHEA18BfJWZLATJF
dXReXgxwQKzmw+QLR7MMs7qKNkFfLyvhZyUuNZvuNLyFPCQrjT8YcRx7axhb
O28FHaLK9SevnyLrxgkBC4d4P4MzNrji+DKJ/GXrKcuZ+nWVLW3dgwWMwnSE
ybNf5tTtblpNONY05jrunnNpC9N1Z3PsdeJ3uzin5eV9djQ+joFZBsj8t7eB
bgyCPJyoG2T0EJf7zSwhup1BnnfDYXxDBuigRf2GJ5/XUfCn7QjZTD8KQhcQ
/0ejI2E21VxBotfed20RzqX/eVMd28NU4oNKN/r8Fu0lXcDYL4pAS08Mp8NB
dsCRYBn0LlrLdVRSMAbG7cViMsIyP1xCQCHYOMx7P2uXqjU81giREBsM6MeV
QmYpsXTOBcL7IbnyNv88QABMLEJJpCObXu/HWRhwoHQckExgafG0W2Xi6C7h
R6xty/3rxDuHspS+mXx/vqX3oWri9sjVJQkbW1eSe27O9uRAWRJreb53iWNK
L1ThfaGii9ju83Km8XgmwgYHYsbQOV2fFWxiDcnfJh5LOoNnsYOPBRfqZ5Mc
XC+8ZJi9uIcipL0NvymdUnmvCmGGHHJ4yPYyu8vzLDK5DsDTMse0JQBmMq9E
o9KbhCBM/0UP1Ijfr84oaWvPogvcvHjKv0vXgC/JfVQh6j9hVH26FqHgLcP2
TotbF6tNxytoxOPCY+8rYi82LAh9lu73yf0z1Ur9eASGzWfLrztMFYM3vemm
dAa/MBny1YfI93zcHr7hkP9EFjPErSzMMiu8+Y4oyOFkgrrXoyJlkZkyFJMk
kajjxvdV4eji204xDrVRDHZauOAaqN8AMT48FbC0HocMS//uMD7ReySKXbPV
ukJnpsNI1jjeesNXo2v6XNmul2kpIsJoQWVPCGmdJ7fbYLxNHr2LHD2oEQLo
3UjlHRw5ETjQQAQJBA4hbWuOke4iOAw/zNjlFxb4VB9YSBIN9BhgLdJ/clp7
Vt4C4FbWyk9AvT4Ywddc+CkFNUHNpgNltMD/ke9kPc4YglG/qBxNgv4Qgfsk
4uHuGC9oX9PBnM78ZsXpIvtL/tSKYSlCrdOQArpDjdDOikHq5G2/n7jau70q
IdYOLAhXtNre6s8zCrXPQBGke5incg2uL+j4v5i5k8ZeaRZKHZTKVuMv8o0C
HNsEPyAPPB7yI+On4kbiPXE8uG5WZ+Qc/UFC8nHGhwak5sySXB6YGf5NxpXh
vCLY9FSpqc8M2eIQkzOsOlrZ9UiUGsOg0Zvq0++KmwERuwPSDGKesLqNTEQH
UiRUcoBOlyznksQ/IZOih2AQyGigEg2e8zmOVz0ZeVE0UfbBau+1scVuz2Np
taCoQmO5ZZTK+aP4s7r07UakfXqG+YqroFebG8DvHo2GlzpMstdBhrqZF2WW
MeJGlohtJT+QyG0YGCtyW5fKYgt2LIEtEZABuZsiL0BjyFxZl42bMmIDWjW4
sHt849RaNv3vDueq6XWNnSGZM5Ka+7GCAbs03/CvVCFT0YL11jocAXn1CarO
w6Xz3xQ6AUEBSVcNsq2cZndVSze1mFpDCPYkMu+t6ObhNede1ni8KVb8A6rm
A37CW7uK8cn+ufAsUVDpjQWDD+bGcfA2n4+J+qwHt0SEYlyexV8EQLRWTP15
E7cwsOTJ6I3NttjkR0HiZKhyzUH/Oi833+12zm/U43APsL0oW+MWNkm/mEVy
qSyK4XyDsPxWu1x+yQ/x2AQ+dDkEGlWCClYyIWp/dnhT1MmigJeoKrjsq4s8
xdF1u9uFZMjxV9WszfXCh0ft9oInmsFc876WxtwuWbT+5n/9XaX8KySu7As/
SoyyokysstJ/nJZ+xJgQiCCN1qbu+nGb0NwGmYqjZ+UvFclaiIwEJEYYbgYM
gWD/OdJuU15/jWLBQ8zog99Ku/5hWMPg140f3wtMspZHXUE+SRJ/uzT5hTE/
IBF8qRvMOvNq1GN5qx1JEau8EJn8LL0X4ufOqLAeFekp19pbn9dVgXRHCs1V
yduJXqg+uJQBm2FClY1+BlyT87OZALFbJQoO1NOhjQ/Fy/1orOIpcl0CNUtE
KvrBft3eDvE5F/I8Utd4VtQujXYrljqcqK4dxagb5B9JtD/nN+YIPglcFd33
3f0/mBPhxsuOMmI51x6hFTttUG0cSg0B+qHSTlBveuG6oN2PXZDLSYVu5Vaq
w8D8modadmrZgV3XE9mxzpV5hTY5BbpTu9r1+oelHi2OSs2ynSFWh8Ilqshv
eWS+uyZe29u0GqPPAA6jz/e/empS/y/L76bfBTPWXpMOwiETisMbVRMwalv0
soStvtopcrj3T0Pzw3rxx3N1AXNHVVTgLANumiCJGiDolSCHPKSBeV5G95Bp
L9GT3G9J95wqPu5vDq7vI3CG5kPFba/8eDPWwsm5WE9H365nMTnVHFitoatZ
dc9bPNrH361+US9kbAlA3nX286kZh9NNH+GZz2j6l3GynZNDHIrfGJllF6pA
al5xBrTowvaoAXXDbiLCCDF1/mRkpQRR478P7wd/RoSwoRGoBC07V09Z+DwL
YzciosMXp2EpFbgkdHtRhGo1u1dOzeLtAXPaQ1D89egmGG8RRZX2iDOgoTOV
XxWeDB4a+vQ9wJ5gd+a3YYdASVOCBLhI8wgpQ2jdcMcqKWTpV/RT60EVX4YW
EO0TjkfUKcEt7YPdazSb12h603Twc/lG8Hdwq2BQbrSoceqMOWR5Ho57ybbl
4BwTNWOT2hjIYZrQeNuddanQ+6c8cI1fR/Pik3QFCakIC4dVWI5wNHaSjT8V
ro371mQoeIPQZdk7zPIOFjoSFGUvhUI2BqTIooRudypziROMmpHORuTNFPPK
Oj6HRCZN0zxEwrZtUYET7ejNEmXkhK/tDFgvoB5kU15a6tD48C6f9evUb+Yf
z66hzLVCImAeLrXoVUEVT379Bfrm8vSTYJZqtCz20JI0c4nGlVQW/eIAp0YF
YirtcPBHgpAnD0JvCKq2cl/X3XJx32314wDHLuLXQ/5dSvmBgTv2QVTyUICY
IKifn4V8UWKjeh2rJHCzE55jvWwc2NOordQqJ5N0blk07g0VWIOskhiyCQG9
UJ4fMcV52B5lxthvQTOp55FVGrT5XjKdwRxfboNHQ0x4TuWJdLurWqTM8nxQ
V3QR1VA90+8ZRRAws016UwJmDHPuK8+QKAIPj37Ub9Kc3/pYmuF+OZ9PlT8G
d50ZUaDqHdxduHVzShXkzyOcAp2sOaWdTrNgCxlJzlV3QzgXnu8p0RdxYGPx
lnb9jhLYmPZuQjnCWW1z4cWKUvaa3CQ0jqolPJiXCJqGKVj6n9A7OS21Cm+W
ilBzvzaot6zXeYT7ko3KuBfufFJ1/ay2nKm/JSpdbyPIa7Nq5RW59xrOhcGB
CVlaoOi+y7Viru6GoU2TL8QNPF6+wdaz6zWeMDD/dxZ/dQoKBIqr0ISDl8Ma
BU2+BgngZVWWG5U3Enfxm0twqvomYrg+GoFL1Vt09hhy3lbmMNC5U5k1CEqJ
k032a7fUSyQVMmrQPFEoMV7f8sCM2HF2xtEPJLwDledhmK0wl/T4+SPiTJr9
WVmHf6Kzf+KsadBLdWlnlbgshMGjevr8BNwGHMhKasS+Z6FLOMDZpvM50iI/
HPvndFfjDBjWbNS+ZjjvyjwVyxstczi38F5SWkbc8QMklSygodVbSNa2kE8s
RrH/0OXimwR7Sha0zDrFUNJSGPw69r3ecXjb46mPqeM7Bdl79SG4/xw/Jb0D
hl1Su973NwWTx9GOK+zavz/aH/iv7hGPJ+GVVmC8zTewQ48YyvtmaQeCrIR8
qXMTXN4+aVbMC6pOcEnLUEyKt0LAhPmdDlt/WAaFNztMZ4e+wIOnx1pV5tea
UvxReNj6dav+NETuedCJ1opVqghgDyoK9K51Dlc7Ryg661WH+Cv4U7TYYrYf
/Kl9AvPdxkZQ3lBR6LaXAkLbIeKWySZNh8SPyA962blgTmHVQqY34gqqcnbq
+eQWqaCzKgvjffEsgIzoNjpu4L4e/kzLIEtPXO/H+8U1TZEJ/bHSrmq4uVz8
/+jDJTjCDpUprpgNZwOVQPCNGtfB3IDH/BDZmdkn2g+IKixbn32/VGP8FUz/
qRpTTveBfj92GXpbhizuBPvl0z/hMbNih0MguJ0C+cSqhB7YRorXuGzFPWBT
tmEqnvNHmFAZr1CqhkYGk9TW71aS6QRlbi4LwoBTFrRPXEnSTiFju05HU6gR
4zxgBw/j3t6u7JnVsAL6V7MowocypnAXo0x5fsR9hOA80f8s08TaglfZInj+
olzk46hqfULkZJhLxx7qCRUQL7TQWBE2lbMMlCRQ4w+/WPPrth0zeDB2n7gx
BGn27zo/wBfU46aK2dNzzsOsoRVRxBnkGoo/bVOcGLUFQG1inl0+dcxF+BSw
UP9pSRHwDfVmo3MBkT7ftC01YIlHu3zPErvRQterR81YvdM8w/2JdESpIUxs
1iJg+6YEG4S2hZ59Msegiydp0ar0SCZx6+Fn/+bcPUNGutQHAY+VnhAGKU6I
Oi9PTj29NTSEGY6otGnHhraJM1lN6Oelb7lxJ52sSbBit1h1j/3vvxFmoUsf
5Y2b4Odw19JVw6lyGDfoE4MweBuvuUvWYf6JpPHvupplsoqJAcq1oDZBVJKJ
JYwXDJ2WYhdj4srYR6vxhmYtlbVc8PeUMAiciBZbzL5lO/grfi8IQkRGnh1C
RMuCgDPEinFzutYHFL1CsCGNV/8M44Uo2Ehvzd8lsLLlatC+Q5LSjrWFDBOj
o7aUwfDVFdE2rq5tUmCo0WNPizLNKf+/eMG7Yyrpyt8gte4Y9yCPXvy4eZhk
vblblYLqyhpCOvyKrTsrKhk/ea4usTPHtOL26FHN3UpL+nd3q2phUII7QkPC
467E4aZdWKpZ6smlmoAK5c5cL1sBIdiEHpluBksu2UUGB3WnSMfc1veBhyP+
QV98DnP5wcqhpnpHpmBPHUTTkxUq9KpxP54+k8ZxV8nWWRfgRip68LsQjibO
hyxabZNlv5cmnaFGaiGRUj8XLRb3jfDjop0824z2DAja92gAdSVmgrCM/8my
/Xe15BTZFGQ6YI66OWGT8HNf8xeWOg+HxWC5UzaTcGqyXPYJiWPbo8lZL1Jz
rZVZf6nsJJSmGf/haneLs9bE+dHGWx6BjzecqS3t76lq0Ts8bdxgIE6HpnLP
S/5nN59GxZQ7FJKJ7ajVhLo7ftkC5zF+DY+byeo9AZrXKPyUL+iZAV7m43+V
xOq9XXs1WG97iljNDuQsb77wnZuP/b6N6Wp/y3J9orS+aj0JswQWaxGONzYz
djI8fJRQ2lpJ/nyd7p2jbfJyFwjunvldnmP+Yq/nHUbPzUpjjSNQ+/tN1OIE
ilUJmpMZOS7O5s3gmWXKyhU8CjOmTBxeafBVbJg8rRR2b6IEvOluodfgTefM
AENHkzlr2+gHM71IQTIZ3V0CMgzRIzSbvfVGB8iQPvxs5SnQHa15i2m3bZI2
HuTXT1/bwwrW4Rve6BaHkikJj8zDAzB8nQYJRTtha5pfJtbnKLboYRwN2bkd
rFNQthsdGmkEDbq36YATRtRJdLzOPRHlhHPghMm5BXefbcLwUHUHLYvQ18He
IXNrwFX7aFlt83xe7Dfzj8T3s+UPZenhihomPOsl8n3k86iJ+vlDMbpRT7bX
OYAVb77YMOJtSofpn5YGJKxSbyFwW8zDVzxD/X33P0NyUlNH4xOArYIVakcq
7eDeWzh4zYL7Xc0Ns2Bv/BvG7h9pTtcqdMA6ZJGf9ULj3nl1WCuBfwvJVyF/
kSN3ryp/edQRg606WbAhulwHQ7qL8a8wYT7w00t0VvBKc8nCqiGx9aqiy0WT
jj5bhQfefCqjB5LJyEMnNvxPecz5n+FoAClC/5KWjRa4KDpfQacoX4jIa7/F
IZI65ZRtF5A0w+VFiPjHNvI4TS9ccEDrGdfX8XnLiRWGkGiWHb/WAwwtFk+N
UD7jmtT1icVtw6m+67eW0DcEuyu76p+0tyi5QP8zHyw9U82JtlSB2ZWrvLuc
IKyLUTmDh/mt/rjX5VaFMLI6FTIP/J2BZEUg11+AFuhJqF/uWH5tugU4YfcL
oe7P32+E6cqXotoV6J+B0KN7zWsC/AxCI2Mptfma2iBd3MzDEfnS4Bp5y8Le
t34WleMqWV1qaoA+Ohek5iqqppgqOoR+xwehYDSZ0s/QbheYK2oXMcZKuY8J
iTOJFdYcx0f+WgNJtrCauo4JkifXb2A315okuJGGWgKbEFuh+NVxhD88qtaQ
9BVBBxV5AetN0DVpwG0qm1avFaxzLZj7LWDDcPdUmyvFCfc6OIjRQ62crXp0
xBxOB6YCuDZ1+p2t9Mc0mpALfPg5Ny72vZ1vefMYQPV/OURr553va2ifhAwK
wwGcdRDh0zi3Ick5uPspi4BVLINJaaZVqE78z16GBSWnskAux+2xuSGS2s4L
vt7b///5lUICaTiFNwdPA+N52iDLvD17SfTPwxLhIjWn6p1SZwbaYWtI7n/g
1MVjDjsrYtlaCXGTSa+XS3cu6fx3QLJeu0QZloUL01bnqoLMe6S1DJ81hYxh
JCAIvPO9OlDf6Aoy7YoMPoxv9W6ZlG0AjhevESee1p979IsRCJgdhWxFr8TQ
3yfivOajXouxg/zpFYwilo+fhLzmxKgaR7VpRv0UNK/xGsuvoIO2Fv4hi2MB
U4hn9TU22cAs1FbHsHkM4zouPyZrJ11j3Zycv2mH6oLEMbArcaKsPwqMs8IQ
yUOm/IhOwxuaTWvkp58g++VeodT8AYky6o3nvufXiphYq4znyt5eq2unoV7T
G1OTYPT9suUAlJv/LMCuR/TEurbXgfUr6MDVLcMRroDIDcfBn4qFaHzjFNeN
kO2oR2dGgP1ChjF85XV+av49UdXTVnkmXc9XGGBk9vpwRNPC51MqdGv15Afx
NREamIL+cpUePoii1k4e+RlxZQdhIJqWYuH12LWjS5bvnCEebz7FaMc09vsW
bLKASapIXRTL0vE+dJ+OUhdEPpn3ryMFtolGQvWR5aXt0Qx9lRac/bL9gU3W
VdQkxE2I2GQ5W40jkwTgmGbzK9y0d2Zx1ZreGDNiob8reH8olxIk1BxtCrLe
xNOtTCsfSMQgDplVo0Uqq4mUalx+JWi7vzPec33DcXWy8VxPvBZJuSZzD1Jr
XgMxTWcWQcy+cBug8Arqq9kvPvakf96Kkt8KirlfWHd4ipLmDoouItuc7yu4
oi8lXmnKtYwIC+OrhAqDpxrVdH+b0LxDpRtDM2xfzaebRK4RbEhL0Wps51Uo
9L6etD3MvlUycGiRdkvphDytbn99OL9T+b0G0inD4r42GMe+PGB/75smHwHe
ff0S5afephDq0EVNY2lxRPROqz3vMiT+KDcfNmEMpjG6uC4s2cApyGH4FKCV
qtbtTyhd/AiNZfAoDP8daag83GTnWvTIYKdsfSNLN/5jnPx+8cRrk2SZCHUa
B5CxA9eZUNwpIkkfYg9wyZu2xepjxHrbsJhs/hT4WglkOS7cEsQlZc1s/q4P
iWDpsXWD10HH5fVkUx6czkGd/lS+FKtI25u1EzSYtFCuPgaUsSXhhaRN5bvx
F9WThjv3rTHd/WIEIdl9UYkPmvFUzuYSCCc2u6i38dOKD8YFO68moFKIWx64
nI8itkkuNu+eUs5l182qDvMphBYT2o0BL9dF+ZHaTPg7l6DJuhBt5S64lXiE
JkXDgWzGLY/HVnI5BjY/Ff78AAEyN6Cq0nE7HozIi5Hk/RlHfGbn9KU96pI/
seT6xl7Kc9JyFYxOwtkoWQMcm8Q9tD7NSdLvHRYOT8+7S2sfCFPjIknNPu48
WJWCFX8lUgPHp9hDKQ/Msj4oo+F9ZKgazg7Fz6fD9wJ0ya94ZXiB1tP0g9lW
8GTX3HN+qoam6mMTWf3UytPiEEw1JEMyQC+h8tqNdfioL1DtC36L4oSGBy5o
1tpaJ82pVjDReHquHc9KI2wccSsahxk9GTBxwtAG5zMvuYMiv0n5/HFk2zKW
+iklCAykGDpCEk8XwfuKWDDxon7v/qOqb72xayEiL+v3nWnow5PFokbu2LMG
EZSnCdbnfC8wm9sxtDKPROl1xV8cofJGmKvJEfaCTaIL4gAbpbtLSfRd9MSC
PUBZZSB3OuEdCbKzpPdb2HGyaqXYwJRPGzHKo88tF6cAfFOojn7C7Hd2qcDD
P4UpZwb46X1/9LMilvzJM4MWM8muqJRqEHJPN5oUU88OdHUjdLFbFJJeDfm6
8tWodGgstv5GM9yzk3pWtyV+oiyKViXJ0Oltj0C04zrNyKqgdxBiWzMncf75
Qrb123C84uSpcGSxgZzlb1VaZKy2qRq74KiE/+xDQobgcQF6Mik6YBKmZTWC
AuXMxHmoKQCmIZ/vLDTWLeOIdRv2chpmLnQl042nWwfzI8aJBh8RF6Pj+YGI
/w1qDl9lNVsglFnN09JIdcdlaSIAjqquOmbhDChAKm4cyC2Id7/K4yoGXCOq
LNcKb70ykLUeZb9KoS4NUwcsQBIHKxNXTqOruSR86bRGAtcD5po8zLFxMDPa
tDrrbK8zmJOzeFW8Hf5CcRi2dFC4vthS3J+fkrel+hGJdXDSHMTfQDh/EWVM
ihIZ5GS8EIcoZTkeF+LPdU+5QUCaNCltmZ+P+iHfeffeAlc2FjSPr7zj/c4k
XXN0KsDCOB2E2WUo9pxzdcfxrUXmfqZX9bc8DMALPr93U7v0f2d6sve2o7Xd
gnAgG6jh4vagvNKKa9UTGVPu9TjZxtdDpcHuk5CtibLf0oE+j6BmbxlQu5YT
ymuMyNnsQYsVWaCVIvTHsz4UmFE8BrLFG8oaFGMCzGo4cTnLWcDMFUbTyKUF
kol7tlxWiRxAC+Kh8SpXcM2Hihm2tH+RF2fzVklK/P8KGw4S/EBfkesFjdqB
WGAPuFTFtGKZ9lBEats0EEdxdJ7Gnypl/P+Nf6I8fb6zykWensApRX8HWWMr
O+fp+NRcgBv+hsdMrArMOKnDKHZW31pnA/RomSJV4mRLVo643ZkjTo3F0nxj
CsqEp98PP3ti1MaaRHvcqxMStdoRCNpfqdf8P3oko5RVgJ9o0nH7QvQVXceW
CmsNyJoEjD64F9rtOru3T/6vQM8t3DyrIxxsUaWN5K1/cbykPTWqPbcnuRYt
Re6IpKa1n3Uei886BaF81MsiDZxIP8ocHoTkETK5zVnOzUIyuevYdfCi6wH1
shII7VY57vOtHa+01C+X/l9kza+LKls723Oa4aByrtFO+cth1u52NTbbP+7p
koH4gFdi8x0H5Y4b/ydrQCYW/0S9mOxi9NTWg3clP0a04VDXc3ODa1XnLEKp
S2xWlYBuoHjomxEidyi8kRFtkwLwKlLBlC5V2M18iaYsq+wlpAbicuTbRxlI
gMRQiB40q7v5CY4AQtjpCGNkHEhhceIOqU5BBGq0wCgwM43BXcvM/9ZCdxty
N3Tkj7kjNXHjR6mNAoup28agqoxA/GiHsg7f8Y8XdT+OthbUEMcC8P9SUSZu
kWvowdXCr2Xpm3FWS19jUlXb+Gxnve7oQwMPWfhl7veMAdODXARfBe4YBEfd
swB2r2CrX3HNQcB2FD365bHffySU6kP7wH6f5jYWmJo+4Cw+2vFYi+iTviUq
kha0L9/nwsp4KZVUzP0+Ssg/P+xu8pk+B4+VL91diZbYkzf+JFP8iZjezoer
VnnQF1OnEQ5rQ5DmtsIAdSwsko/BJ9X97q4dXRx/V4ZvlHG9RQRQe8xB1tWh
2Y5obVjX1fEFngFCmptwfPZKHHEQzRxkcq/gS68huKjtr7qM9oyDaFapF4RE
FESz1bbhKP/9UNFoI7fiChxFjLyFWTlx/ZS5p/hQIJdHMWJWiEygpJ4Nab5w
MRCd7xpdmjRRbhhCVxPHDpXaSa4If7HNvko31I+ay+K+cp9WmdShzKEDnags
O0CmVJw2V1c70D3XYPZsobXEo+d6EXFjVMD9VOTTdFZoc0QeDCXFVv8n6HmA
Whj1bpnnlvfExkl4A8Ey3bTsq6RalIoCVtJ0TE09puwq+M0w8WL7DztLc5PP
N+HECw0jWtZbPWTmePnvE2fc7zK94sqr75DQJ6D9/lf76Q/4oqkPASgtIMMW
wqFMeaj4flKCwZh2FSWsu65UVg1AQ3bcu8vdFwtHoUILKO9aVnNia4lHn7oA
W9KWT7x9morun34lMhIRn1V+UUHBZMnFp0NXLINgzmhilK7dDsGKhdFsV7Po
7FveNcsBjsiJcRVKAvOCu0s4u/KmDh+FWmJnSajTx0s2pN743YHiv4S/MOsK
UAcybrRrbMgiNsxAeEwK8W0d5wmCTbztCNNRAEhWieYcTD2XndletIXsug1X
10a1OyUDzzv11op2LGIsiP1zajIZOZuhlhtARloDbRp48dgr4JrFhp6yFZwA
V6yhwRB5vvByRyFN9OrN6pi5ZpC6LBpEWc+RK008SfIO3WEFCHuEGoHKRNq9
VoO8ooiLEo8LilnTY9+XPCZ+8sNh+KZx0zeWF4bqNVMiAmEoCpltXt5NLcPY
4OidL4pNsUN5rkfSrEsKwHzRo79xqrDtheVqc4uTAqq8kn0EbT57zUeQ33Xl
yLeKlicWflJ7dZreehhoYRMWbI1cemOFz0wG1dch9DCjK3Xz8CCp+BHQ0VIs
dzecuU83gi18UEAusBf5EnaMoJqaWG+hSFGIXC3pTqdYFpLoJ/AauSqTUKA7
wtpAkJUaPqP7GVuHrXnlyWWR34u1cyF/3Q428bydMABwsZDw/Hu5Kj+x6AQZ
fwtglUqqtq53ePxsQCtIKjM0tFuGguPgYE08K02AZMjT5gaQfxVA6ESmn6xM
hE+WcsVth3N/h8AnKh8Nz6J3xoDcCNwUC7hBjW6yVWyC3F10n0E3ZueN/Rlv
l3z5t3Nv4co9aywd2J3bdFVJXF+yAPDWG3xxcEg7CBNPM/q+EVTzbHIaNyNu
Fq32ifLUlw1KNjWYUxAAC2Z0VqG6VQO5/lmet1LbJkA1qHn6heiuu0UijPsX
twVSyBTnoh+FLHrxhTIH4OKYHkIVqXE0G470fAtexwAo1fxzs60YcpAjDe+t
TiS4NOOJMryFBPLJTyexu4lhq8dx9i301aNYLkAEMKRU3jHqjX7nys2actGA
X/em6caqjz4vvH+HVpVAemli/k9dyaP/Xc1I/x8s4cmTKIAZN2CRTTq5bXit
UVGbj+uFR/cVftd/Vg8jTZcnZRSt2f52gqy38Lcmsfzps6aJNWi0oJdljV8K
ZeY9+pIKYbG2hBqGMHpALsBbHEYn0ynj+moT63Neva5GU4LFQq2rTn0saF6M
/+V9/nFAk20it3IGpWU1rFzrhK9NI/jhfpO9OvQexJW+Q9StfBu8pAtqIQmW
zJ9Af9veUtU+Q2yJ4iYWxIJcsoemuAeK2jcvguBc1ljLIdGmVZKF1dZsAOCZ
X4WTUbCpmy8QMT75DKuhVdL97HMqJaFfA8MVLUhMSG4BtDauBEk7EU3x1tjL
6+Ghjs1EXp+lC5DuKbOSSFavicTkt5xb7afvi02VnKwTbc+w/PztyRLgzbVd
tKrSm5tcSUcH6NHGAgx9mbCnhxuzeR46rHHQJYrtHm9Er0WipCinoiOzleTa
Wt9TExgqE7/A8bRsVh1mBchZd/SEVQMSoZ5TXTAXs2oujTZWJUa4UwgH4U9r
oXgQTdmqPanzGbs/gSg52WEVCBzJ2fJpDB3/88PvONdkkRAzVFnDtFHM3T7x
YkUtzE+QV9Sp428XM0p2D1ciQe1tvQji32V4YFmLbd3NeXsymgv6Q9CvCxs0
X1gA5IqJ2QzKaLStIxnsTjPFSq5fL4ml5ekdH22VJHIHaLncUORB6HvQW+zB
OXXeHr3ESFdXj5fG6L0cRoFziRP5tHVsTlyGsKg8qUVJzZZYIlfYfMJTCaDg
1SltarF4djnExkPWZr+9lF99lfLqn016vvIzmyEJiRZdqlDm2oS1bPJSzbZz
eESpwgZKBjYMptq2ZxUAPVftZbTCjMEU/xV/pfQGUiTf9nvo3GeFirUJbx7L
UgF+uuxFJAYjH/NDeF7Sl4hw+oDL2mvRXEv3huGR5L1omQTrHsMYdWA4jwb6
RZgUNNLIkdAqyXqH+aIQoN2vq9ppJipmo4CxCVLEL4MJZYFG2BqUkDcuiiIp
ZH9KHKKIYd3MGlouhAgzi4X/kGMuFc6grTc5oJkxkWuPuy7LvvtSmzJ1Hm2A
ZfTWcTQuQcdGFICkyPlRvEP7rtpdiKlaBHkVSDHMOwo3qukSSRzdrqz4tTq6
RI9nT3hCcE1n2j8azX9Uco0Uq2TP+KdsCM3Kp3cWUMd1d7nwbp4d4qC6ucud
M3W8Uv/j15HISgTUmfUIgetB3khW5/aitIrhsLfh1tqrHN+PhwjzyaYuOvHr
QPIoaQXSx9B6Ieqf63xtqSeKZ1j17sbGxwrOpxn9lG5KplyIXQEspWUZyhSs
gTOhidHItl5mHAh46NpRvoJsAgRlyz1k5T0iwppCY3WUHrbyyFAJzBI9zrcT
i+Fof80zMPAGK1bavUVxcUDWmKLv4rNkkcA7oJDk9U/wTlVd/4VBSICpb8Zm
S6Bs9XheIV6wSVWUIFQyHupOGrIgMpjuTdtb0m0MvitCfaRa01YxKodfrrSz
xs6wZqzFvBW+Q3Nrl2rS0QWsoDm6wYuRS+EQLC/xR49HwwVOIlxuoao0P1az
Ov5u//ihxVBXlxdC0tgZP28UrMc/UfpQAngRj+pPMo6Su+d5S+THt0oFz2w4
uLggu1/4b9np9sIsXKjJ7dHN4+YujitjrAZdZTeQjXrCgPT5pemD7ZNCLbPV
qUgJhVq6owIthTkDgYPLxzjXKJp0n4kBSQHmgXnPR6L/b6lYqRsuUT77AlB0
tbGrINuQWJiEPWONm6Rrq9ninWyt4OeqE2eAADlH4/eLiC266hNyxzKOukT6
GRZzkvq62ecwRfgCOp+4seZFvGfBVcrDZHHzVc85LG8kyYrDGZlXTLmn610m
i6cfa9Zwj2SodyWBF3JJK92VYlSMZCHmMstEx1N2iE/ZGHise/9UyafOCKw5
yIlNJLzjmXH7uBeMDkZHHMMt7+s1E3vdeIyWQgke1pCziAXr22Sr0+BLeH3a
SQ/r4lnhlzDRGWAJlcJIZBXcbGf+YNRHnWFxoPnrGTrwD7R/QHE0J3SbZSh/
rARGZLKgl4YQ0imHUctMhUcZ7IxbbHEVI7r0DSnFL6E/twgRk6MIJGuU8dIm
r0WOOgQ8FQR9yDNHB7l5FAYfVNoqiucQuzTe5GfTiGLwqyZoCaaBWq0NoxvK
179i6c7Gbf5lIi1MSrg28i9X+I+gxwNRVHoFguSbjHc2AMdVrdezNTR/c1qy
hhycm2ptsRxAD3ZjHnXwkrU5D3JEOjpD5pg4jSnKVEMdkFxFcJ1dgjdr5ULT
p2+4bWynVyqPdckteytzRnGrCYUKe0H/a7A3Jt6ssapZGnsBMMlbLfNX5egs
lccas6dtN6RMdnfMmnRJT/DMJg5JBHShXQQfoko4PUKiSswHneXj/6hnDFjY
B/9b8rk/8h4Hgks7ORKjVSVOs2zVQpqfvedzuya7+pKOAU2TyscHzP+uwfDZ
2zVkCZAn4gaSTe5tzVy57w3SDmhmzd2SuUyKsBkiNsQXd0eD/dxk3a/cIkJg
BTGxIdTeCcfQB7sI9qdAzZtUWaYlFTz3FYYGrmWE5cLnr7YpRC6BA4U64Rl8
2NU72EuxCsuGMjul5x5Tt1PAXzta0V0fD2LRXhh2piddpVyTSxr7D2PveaZ0
CZ6HXZKrerzvDTmJ0k9+TypXlW6pbHuEbGK5SDHRSTREP172118tdXHi1GUq
x947nB8JIcCDBJfGWC6LGIZUB1ku+mgQ5VzT6YAU+ZezIKaZpqUz+rQVheqt
GctFdH4MDkRkYn0MXDAZsc5al2FmpH18GKQ02FhZVJtrGvURBICxTJIEoRPj
jOPWWeKkU/VFnij/UWGG1xOsMM/JHp+V7CQ7BQPnjwQgOpNpUP/xG691tcX1
BsVwG90brMwGmL7WZyEWLGplNWIOf+IUVryJ+wlLBcFbjcckXG0mTG1MRYNT
ok5KcYZouxUTwjz06VwmBLRX7Z7EQCbGeKzqHCr9oAElFBf3+6I1iRxU5QXO
6qvvr4vVCLkqqsYxvC2p6ANWguQuqGQ8hweFVjNCGwRgaiSfdwGcIyGIYNUE
W5OtX67EDPqh1GQn9Q8A6lZrdmJIpBKqn8Z6n0yAQpNm3RQS63doDrzeqj6q
4PfVlwYwBzLSN1H7nnR3K8z063oyQlrSfNzxQ0Y+XgXLq8LfcsnHNDFdIUfp
zIACtQslJRSF6J8wOcvMX/y9v/gJ2w36L9wAVsIuO+mLNd9l/8s9kgnEAWY8
IVN9+cwvNPyOPIIusOuRehMyg+/oY7XFKi20rEEJRqvo7Pj0PCiciqupv40F
8/oU7c39pRffNgAPZAzLEMgkFoKnZ5/7Dtwvpc4rrNTdRrXlQM+0NrrZn+EM
micckmU1r4QhwNjiOiFoWybTMe5nkUqDdlhB2T7NEtTeGRsA9O0Qk0qJm669
KPBmzSgwSQGeSDyJogDNwAxJIOuXIJVGRsQuqYc3kKvav95/P5zKCiKwhrO4
KK2Ipcte11qeyFFDDyieowZC1sklfkIFGIhVpI3/QwEKOiFkDFTjWPMKG/hf
GMxyEEDNxhmuvxx40hQP7mO2mASxbfvZ0Fl9Di+CyRuyvOSHhQ24Tpid89fB
lAD1XY/XarM6re6ii5oQJuWZT3lVWHADC7cbzlqD6vdKFLdzuER4/crrCGvK
/r1ZXiYg6f9G3aXb5VzAe0bgHjpGBCCnunLaC1Cw40GVAtcDirT/gaNUmRYE
ZIUg9J1uLgZ1Ke0OEw54pwLcbvrQ3un3Yyv/e84bzbJn32TJJjdZ006NpdeY
ri17MnXZnQkBASvC4vG8DfqhcX0i2PzOPydWABcg5iAOp7b7Y6V14yxZGVQF
pBdFVIFhVZawd0C+iDWnXxAP6QokuJwOsls1bwClDsly+W5VabfUAovrECEn
EB6FwzgiaQk4Ruf7rK+2jfSAZTt64+hnRuCLDQg5lDbeytlTSv9i+38JtZSV
jafa9PqL8WuP246nczJwipjjII+gdEZiSQhPiBobp2ev9qzykGSwm0JuAP+w
fdurss0o7OwUgXtA2SeYxm5Dc5/qSDFtAltdLp9IvHULqWJ3Si1j1IxfJEFm
3dGpuVu0IPcdqC5kSdAP8Eo3ZgtKGPRVZFmWQMCuuSq/pw0auuHMDkM/Xh4Z
eDIUKC7QRIk64xJ+kfp8oX6K2qe3mXEGLs1Kxp08+qWuVIaCkU4ZZJdnNVFR
jpAlm4D84fuL0YefILi/gHlTiCRdPVhw4pFg4TNnMnu/uXZt10ckFWCqxeJN
mbH4BH59E9VgE2gCrTfYPRzMI5J0bamQJn0HUEeG8MCuqN2Doz1AoM5oDEH4
LdVQAKh3SZxyEHJr+OwhxqzhaCrd1zuSss+xjnOKF7+G7imfgz8wJx6cOF0K
riDouf+7nBk8Nx0dEuQ+U9GglRPZSbsjKDxWZ7drYYbVkMG+Lm59eiptF0Dr
ReqjASQqx9K3iEqQeHxNCSa6w5qtM8Y8xBjGjztWdwBjcE6EvgGYS4m+9Qee
Y/HrDc66PVIRaF9LLW9uvJvzH98IajAU3gu7gGR9E/LP/WwyG8pn9p2haO+4
KkxCCpSddvM5842B5C4eyUpS37WUm029bde3df7+g6jJEbF8TyfpQCqSbUSZ
wWMZkeFTRaIa9LLKe4K8Xbk3Iw2yf3K4Z91l8/CFWXU7gn98cb4yb7V3tkey
HZ43ZKKgqMnNAaJAdw9PnKTrOiR3yzGptqMunmX+rwZcEKBoPH0M6KFkvoDy
pFUOm/ebPMWcAByLgsbXyGKbGFTvx4xH2mZobsstzlGCcL4+9mp8tCpCs7O3
DWscJD3vFePZOLQSLWpAOwYdAb7xn2LQXXUJ7+RwYL6vTj8sfMyXRNtYnTor
HFdvl+9hTGqhKfAEV1/tQ+sQ6udeWf+bEpuGcPwBCpa6iwNI6g3yeG+3GNnL
0Ddgu0WRs1K2GnfdgVUp+WIBolsVNqifenbm5vwOj/7v3s4lQTIxVpI+EfPz
JiKrRj7c0UhVfYog92kral02KlcRh5uZI6560m5yV0bOQvh4nXQjJdvf2+SF
n0LEWP9Jr+shHClYq00bwpWe/37oN5+4Fz7n2X8L9zM2KhdlMfaDl5PZfwEQ
KcomkJlG0CZGniv1kGSmYTSimNX+gHaVO7BrOB6NbEVr58ok0oYh8vTEyINL
PoMcUK2U9cCmCt8LpkQW1UjvRj/GI/nmznhtnNGRojt2eHFzc5l3AJGRaXf7
egDpASB0UCwVdcdg/yE0r/oGFdSqGSz4dlpY0G7EhvRss87facH2MFpPDvCO
OtJmjJH5JsqwUxubIGYv2qz1r3GqQijK8FkpyyriwBKdVwkWUudgPvhQCBb3
Xazk9L9OoGqBj/cZgsufSi7Xw5qOUJZIX/0IgnIYDbQEMC19ceEHQjJbhYZW
/Fmy5NtZy0yFPb5BBcfMjtj+MbwvjVTdAaFszd7hLmelv1v/Qg38PuYPjzp3
dJKsFtBs6clWTqlUEiikPvMSu+1I1dcn2V9WuddfaKurZ2cfUDmH9JhQgOjb
FvA/WKntai6Uc0CSaT8mSwNYsWQxTVDMgjcZxPsJ2O4887vNxw40qRT8ywsC
oH1Xqluq+L2PShHy/zcaUFyM3pWcK+VBcyyXtpGFoyYwyLMa2AHjj9uykLVe
+pFM5BrF7WDdmXq3pczwFIZcntLqyFCwXJzcWWsjKQFj5oEYPIQ7HnyIYf5K
NLCXd5cUjHvWGvqw+w8vEEBB81maZkEe7b/0DSTB3cGRhab4B2KduNMxWv9Q
kc6Mkf7SKvryTVs6UoTY7zvahc89tf6I5j7ZrKPiQaWoHmrI4EiyX/X+oWoG
PMajVrP8CicxDjy8S9X48Udld4KTuIVfjFYfqDm1F/QziYK+AUnziPbQtUbm
oZItm7x19M9U1qmH4mLLEhVAzedpi8bFz0VO7D1rXozcSlSH5IxvI/fgiD8+
hb6SluN84edcV16Jbqppyp8X4x9ByY0IqiTinoegEvmfjgE2ezZSFTbThU+x
4Ovkcr641lzo25jHbChF9AVQvnjBotsW7Zhhr1Wbudv/7Kv67wlu/6ksIkvp
JiBa49lHl+r2syzK7autVqpdVQJVAvkGPZo3/nI2lKvMgdei8pZniXuWKUgd
ozHEBqUgbbXEMHaFsXh1p82Z1ZQhlDt/q3+if4H0pld79OlEFlYPL2+X6HBn
ryzh1+KO38ZRM4VVJKM3sk3PwHoaJZ2HZIpG0i7tura5lq0Sj0XFrCmTyQ+u
u+ydeuY4qKcczX3jO+yLFv5oyfgXLjJbqgTEugmKxHmqLndpQBLrSxgWUbqS
YekYChsWQJWtCQwwXhLX3+r+9FbL7A/462rykdL58P0v4PBaZP+4xvUbHIOG
LK2KBwVi7/KNkkuY/VQ3pyP2GCLYR6D871rmVFf0gcqGXF6y2RirSKhKuyy2
qbciglZgTv/BNrdrGA3eS36/IJ8MEiWvyPGDU2mPsPHEewzcqcWXH/3+Gw6q
Q2SVVu46sug7ddh5fU+P6b4AnueCtL0ze3rQCpF2Q+4sjeiMNYEG8DXfLYfw
FRvqaim55N5a1sZHUsBl/OJrRNnKV1Pb33rKXgW9/AvKsWmwW+B43kNnREi9
gmz9tNC6+MviWuEhRv0W5KlzNbf1OWM50SRXxNAQN+iMhUcpXE4wlPOj0jOE
TCckgxyBiGCctjuT/iaamrLt/RQK7GieAzXABgmmJvSkByvEcJejGWoE+TjZ
3Zgsxk8pUyxAjyVBQrtTkvTI/xi6vmrznG7SSsX+NUqQNVQnzhudE3tUvt4P
7Dm38XV5El4zTIWn2IDf6WgJZwkaYESZOOSwD5Ia/cSPcOW1GwHws18SGeBj
S9/QJQuXEcecryaJsOtFRcXiNBDm9oTrjPrV8y2rhdHb54ahZoSL+BjQ2xDX
2OJforLKKG2uVxLRpkB2YOaMlSPuDDLxzy+fITr3WUs9zpunBczxFzhnvzVI
HxGFJ3u9iKKoJrBAQO5l8h6LUB8E34kgb8lOX/eVXybTmW2CwzLNw9pvq8oV
x2FivP+tx0QGL3I21Wi0kdRxE/vv2MkZGo5cJcN/w4T6WuFmDzxhfaH6ZfvF
rwU/iqq9LYEQUJwV7whwaLx3n2XpEEkwRzUjAwmwxNMTh3trS76959rUgKvi
+s7EOf/qItkYAGdrNyxbLglgOYUp0KZFskDp42OiYj3AAv2g2+kQW4dAg9Ua
4KPYyJwDJyewx+vhccGxakqiA3nKjmTyuGc914R2Ib6l6wXa8ogJAFNP85qW
mkZetTAaWoIwCLsW8sxSbBvTt+PCORgHjAMQwuFsreuT/X/JvOacgWo69j8q
nTPIyMrYad/GXJ0/CLiXN2598RQ4DjVaXQjhrORrG6HW1AKi/IaufZoa/EBY
llLaXp+vFQ9Nt8SrHbB4YQrJSc7meQh/znnPbfVea5WpbK+01vf/86GqkG6R
FEaIzsLpDbOe9o9PeNPS0xO2cyKra4OioU6wKgkdMEuY+3b1nKI7VPtWTlfY
OdDbnSWHtlWtqvonNQfjkHxwxengaPNXHLqkgZ7DdKGlV7P8/V9kXGnvW834
Ex0njHyOMhCpiRkLRmi1NMXWQqiUJu9n0/z2eQ0tGv3tg3F7HG74KX4Tx8+2
Y//GnomxhS0Anx6KeRX33L+UO17iaFXlWVk/nV3+FX+qijwm+bUnZo91M7jp
2fbPXtCZx9moD9RMna1+PNOiw1GqNgwwDp4YGMKiEXe1orifYOP+jD1vIPyp
5t8m3rZf8tg2095pwBoLttnIBpSN2kBkkfQZSvZfoObA64+OuquM8QctYdlK
+UO3coThAEQBaIixH7L0t/ddvijmXXbCrYrO9HyuqGmcYWXJMFOvvGX4g1gY
603lJzTBsMX6ywa3nL1+3CCHYcymly/KXmx+EjUn6X7b7eiEDorM73vMspm8
Jx759fjUJw/uOtpNXhacVykrKH/gsF5lYwLYTjrMtH42anSqwSVlVK/rg7NF
jW9Z1LIRMqSST0eWaGJQ49dxjwirymU9mjwz1Dw9kX2KlNp8N42yQnI+l5u3
xZQHcIloNtvJS23YxqeYymOWjmEoppZg408NQH8bXMNdhJu0fCgytMqi6ES7
hp82/A/m3mkvCIYU9UxkOcik8pV5N8NZ4A2VjLrE/u8VurPZQKYdIWq7itHE
dycYDCaXufJ/yxNrIx3ldN00rWr65Skx8GaGbR2xMeQxZutvH0YxrpBsfMjC
BTdLeLNFOv4ZbRnB1PKULKOxreXoVFivrXBU6c3YMXJcwvZCqN9NveScXgw+
pzhKrFD/Ajhpe3U2ngt3s32DEya7HY+cUTYPV6dLHnD2DG0re2yeUC3whwSj
eAIwbpRO8KEvJ7iRwEDFlR+E/+6IDKMaf2EMoNBdbk69jEJTeu0OXa42lwuU
ucS/O+I0sBsPkDDw4dX+JXkERGtvAj+1ksPwJi1VvjEW4nEJ4iH2Zu8DM7g2
ypnKOSGKUlt2WfKdJ8ih5Fb4+E8Vh8xE7nNXSMHxuU+pJK7Kdhec6pIRAAMl
T5jwENCASOcsh7pDVko1N0JCnp746eI5DRMLFK90LPr/3YDumURZwHw/2y1l
LcM4xXetxN5w6LM41JfdC2IbZmVhbzlLBss5X0O0aS7D5MLK70iWMh7hbyeb
0Hi+gOaCBJopyG8fNFMhVYAZ38i2cscz5k1hJTz4ybvcAzHRhPS7sS/fT1El
BQpogPC41ur7CbvJlhhnpdSwga0HrWeWglp50uScu1ubY028ln7SZppdWpSx
nnkwUXlhd1ihJjem5ijVp5Uv+gNAdO7kWKsoS99T339w4D5vcwmw/oi7lOjf
GubjW+FV8xrXY0hi66YnMo1w0uRcBuJvJ1oNqZz636GmWTyA8dGaIF8MoH+l
TeoC18dNRoT32TE6wm0r9zcIzW/WtQ4n4wtMxzlBOVMTEBrwlwyc4MfBAics
jJfSNkD+GKUQH6Keyn7w/VafoIRvuWNgk7NWzg3VeXcvEft+jPJhh7Ssutmt
A9oYHW9n74yRWHAhz8OdoXCNXKtIzeNBLaeOvZC8+Td4iu9Jaoqzxhx6lPL8
uUp7h6yazZqDEeFMZibYNvuUQWAFsPPhSMQq9/qGtVQy77hqNuuJOLI8ICsm
S6HYANGicdD+pA0+OjmpxCHPmCG8lII56WvXJlqFEJBPeqFBQ4lia7LGzedj
RhrExEtN1f9Dm9CuC+ndPQ6+Iqb4ylXX4m6nVjM6tiwettB3lvWJRVdim88C
GK14ADdJI1cmVkNc84aTWnqLpUhqN5cpYOz4ys1agYvw+q9guyTvGw5pzleK
JIUAc1XbyzJU8hthVsCWJASKeroAVKeozZTFcIgcyIPLme3fx1w5332RZ6rA
F2+iujumNg8ntpDFWO/mQF6+dPkwQaRhaymnGblLQ5JJUycJKxMKTWRpum2+
sqGiHRpuhhHOuu4aiPEEKMW6TJV6yidqRWunuX7l0R+zi7QOBLBiHVfnoJ70
TGIEy1OGaU4mWAdzD/Zg+R04u+HSaSJHaICGPYLCTBclT+2vWgcNJlih1VlI
UdEVXhoc9GwoJOkGeNtqLzTOp8WkBkqdPfiJCuH3uwCn2kPHDC3nsD6MYrXr
d4pe/TzpN7Mqdh5lN0fvQufNml9PfbeMzDqJkx3nEzz5ktORTx9vB6WlAhLt
MA4gbrai2unf64qOytIYKlnedQ2oXwS41ePZ/WfxA8d247NLLPUUPFjR7HuQ
xY1ZVYEvNx7EicmCUDE/0qHSaYY4n21AlnYxuwsEtLaRL1mGF2XR54Ce7CW2
sEHhg+UmVPx0vRrGtzJ4YcWDjuq1AKkFRe11RCj+0ASZFvsqZw/4wg/lcNIS
QoSkIYGtnAcVJMjLnvbugG8lZ6Xl5yQq/Cn2s1ZRAD32o+IoqEd1CF5I4pap
6GSCC7EgjD3SUNDJ7GuwOxqJgVtVXATGcQCYkSaDeMOEktFW1YU3De3Q8e59
qXzwTH6rn353qHHhmnxzfPROimP3VVTq9mznTsqB43EmFWnjoHHDM9jN7/aL
B3F/4+UrKJJoU19GCazfGQ+v3qSlMRLnOwQPBbpnD0PBB0PnrzsrJms+hkop
v4JpazoJBtnlaGszeJjfwvbFVMKgbsca95jWmrliX9fC7G1j5vqDsPXXzuxI
sBENLe/Y3sFOB7ogcQE8DuW9zbkcySJGa2i3MpiEoqir+8F7XRpkXiNljRv5
Z7N7rf9Fd3XZCP+iB3GgV3ESs2HOMtTuRKv2Cxl6/nb0F9GRce68tknASFDM
28l91Z5QjFpAPI6WYwou+7FwRWV7UUXKfKGlFODjkeOeJHT/j1BcIAkRZOmd
PN32FdepMpuZwPDrRw6yjZ7UZOFbzwzRHUV2JDXtjZFk5AFokaRztp5ktbOK
zvwEMxKfaJRt1Kvne7sRaQO5Nk78TpdpCxYOoaLyRlCzYKTUw6Cc/z7/NrKF
VUOIe1gRLzrFXFUPeuzXwCDGxWxZcUgFWr5MqjmzXOKMa8qxWjSekE9YPJJL
5W0Hcaaj07vITpgNyZjVVY52pdn90zSG2ZHi8A9BdBzhB+IV8wwSA2t1jyJE
sNhohB/f0ZsveztCIqQoMCNo+ree85xIkm992VgfN7NQs/aG8nbR8/SMLPm4
8fhxpYgGalONVluYnU0JCsrTp7U9qGcuOOdBaWM+ENvTKSJsY5KPzKtMyKTq
Ihm9s4nGz4RleuT1XLVA7hl/5b8NgNWG5j99I5ecANGH/jSgzkYSZ/idlSBJ
w3++q9GtAc3VXXtsGPGR7SIKvV9G1OZd5nIknpnlzC3HYKylCoVNyO5NvcUI
1iCdcUAyEUE2iX3MG2JFs6eYluI679x2wFvrQDzzcF7+UZATPChS/VWFX6qV
qFhf0MhweXzpN+mJjustG/+PfZdiyRq31oJhyBDOtZz2MJjLSD+YqLejSCsG
Cqk37RpXAPUnPLg1McuupwkoCJ6ZmrMlutND2DMGdNXaogLc+lC/mrXgtZ9W
7Gq3Is03RgL6Ug1u98chc8emYUIRcEGmtYL2Fgw/mWxz7B3iIPGO7n+Niph8
nfL2B2O8831eF1mOlIVcXyQxfDxcYkTbH+rsePaA2WFgJTUTS3kSBeVkK04p
3m3OPMCJiA3YTOGi8c9LoPfvnzsSr2ptw4vmFDX/e9u5sQOuA01U1VXCL5T4
k/OvJ3g8EL9UnY/ixI9wICdR0olXDyoLGc+LWDYvB6DYsldzz/L/UATXAYg0
gn+3pbOOWN6ccvL+0jgiay4PWDzVddWSSgjLwx0VvYKE+tLyepOioZp/q9Mc
KZgt9j7wqrAxtlMfsEwIcJJCmiWZkTZDKLAygHC9S9ucr8F475lOgqD7WNtb
8tM0t1W9qtW1w+VrfHYfN17WRdqzMs6EpD9WQcBUwy1d2QaCiZzf00H1cBtt
DE6nyOlyG60tjzXpY09KC0FIvNO+JigO+gIhugexril9QRSu8Cx+KywJKolP
sGCzczkXj0eqWh+4Eze5tF+0OASk1MksHxkoAx2TCniOzwa3GmXWkUb/O0dl
Cs4nJ1EUoIC/Ma95o8QoKO+0b+QoR0ntsHvWWpnDwsoyjWBcr1363lAS3Vty
vGkpGE6jY+DbaiuVeB/ppwKVjp77j+elzj9EiKFvpZx1A3xbgcW4G5BO2sT6
9kaPbe1vw7Wm6Chaoz1lpboABpuMlhidgxBP3ge74fkqRVtNszcI27TPGlmT
Fo3kTdneLMBCQFxRhIC/G7DPBHYOUfj4mPCIHXA45NlT95cf6cR13f4cwkUm
m+/fT4TxR0Q4ZxAy2RmEwCDSgQXJaCX1qBdIHIeUrCm4dyTvRr/xhB9fqCBu
TH5IR+9aowqUvot6Jav31QzyAGfwbcBu95HjxAdiPEjNWp49AxgCUgA6uRwt
SlSyERu/OLQKIaS5jcOITB6mpkVY8UQiq9HyelqZt8jFlcPyuTFGe14TpSvd
3afhJKEIOpWW2kBJTy5NFRqoejSmkXoANGo9JaM/uDDQR4Yl7xMkt/O55hUG
r4DwthEfWRAAmEuYXbb4kxWZ5iw52Fk/ckGDfiF9gIbC51V81177/NOn7o/L
grHHgz+4QnonMgUdIuQz/GUAl2YWDOZW/VSK8RTmNNy9rB8k8v4q2zd+P+Ao
Ml5dpCHZ1iYrBgVs0RSjBhs08AOLuj0EwDRQvA9xnMU2LFN8O7VyyKfj2S3N
FS96LkGM7ZAjgOvYRDk4B2jF9qhJuob2J5wvspTNGPuK0h+mFkuYikDbhvla
5fSylcJgtA8SnUUvLFZVCj/wYZJAENl4ky5HTk4t+LLDvdxUEnpxOojGVi4M
/eWCBPtCZKnA+Ijh87AfgFJbbOMUipca8aQbcmJdhv4L/1HSbWlkvu7aFzuR
oE1++OuzNFDxKoCOu0Bcrq/5PbROOukduuXqDL4wrjni31SdbE0riCee+RgU
aLf5EhYtC92R2Nht+evIHB1/mh1ESPtiPisdqyW81+PMMC8YP+YjiHmp3mM9
nqzWLED/LSwO6qWr+s1Fq36cRF164LVPy77v7f8iuKmB2gs5OptOeCxL7I0U
ljCk6/6ZO+EE4LOXiu1CUHPSJp72Ymaz/l6F4iAGUe0dqSZBsk4SMa79ydSt
5sIFirMokLN47BFYhv7txV8qwVfpUSSXwhj+JwVHk41PAiNEXdyVzuNJshlp
xzb9b1hgeMjHm7pEFAQdEhq8MPvPbUSNWja4tsxNKvwSpCSHIS4VE8XgfF3h
WR+esfJfiCEcXJybEAkWlgI0REv3l8ib21GH7Y9mwVy0Z5kp9K6hm1drQDv0
Adtvcp14R+dYcBrxksNx8zwqL81CPAz/HO5adJ8OodShHGXNgumWUC87inn8
6wUJqgS/nVLorom8cGfnsWSaD6MSW02yOf/jSZxAvrkqpCPsk2UnkffJV5AO
NsMbmwRInaKBw2fz+fvZqACrJVPzCYjbjsNRzDe1M0EixqnFxz8E85QLp7WN
dGV/qhjY+sKVPKnhC1iTO6UPs6mh7Rgtw7Lcm/QWyKsvBKIV0e7lwr7SxvYP
nce7bqmDCgDzHIVmWIdZIg4pkPFjxVGFQ4y5tQSTzixhoqAp0Sl2DbDTl4Ue
MiaCp9dfY2nTF7PW0MTvCp2XudXRPDlBIN8cQw7W2WJUSkFbu859KeQn9cG6
OiEpj6CH6oZR4eCEPkXpvIAeJwr8l5kibuapEk245/I4fVJoF8hOn8OXcAOm
l3o194vwj3shyjt6HrDEo29RtQwUaN0wv/HLuA+4w7GRsDIHSIKuAcjwaZS6
c7hEOz5coa7SAdIkg66cLYApkSuZQpRVRLvnDy/hdHS7ut2uiKMjkbzX5IDO
USK31UFsoOz28OS8Q6zj2EHHPjZ8iZxnpjn+Mx+9ZV4aygia44kg4c2Ys1gI
NlTRqdTJIhAF9DvX78QOscgH7Ke557PK9AAbamuTYxLbGkhycPDoeWRumFjl
Y3c3D8yL+zHBjJzO40ah3c8MoYOFYmpDYXf2+V1sFmEY2d42IPWDXISgJBee
mLsnVFzryx8wJkxAe5baZolUpuX5cOk5XyyKpuxHlRIyzZ/NYKBswQ5ilphY
mA+Q0QQnbgFd9/NZzs4dsTZ2zaU17j/Rtn8L6Ub7x0urAPKO081NlNIcsTc5
Xw5pcNX1hht+a//xSgM7Gnvmfl6Cz/GVXwWpKs1X0D6xNAsNwICkNVdkN1aU
dpvFGOKV8AsXm3oGwubeFNiyey1OKlH3lZTzF4Rvf3ypAGQ2ryxApfByNpyu
hCugQ36eNgYpbCr89uCK94gc9eIvTB7O9/d9XO02q94wJ2vKVyxythTBBxAp
VpeRKn8cHof/DiVWxPBVkrWZdyJ7/AFjrOh35k3LnG+pLG5gqeLO477xTYwi
CCdh5Ln/QITZ0+M3OcTeMAy0xV1c924M2ldAdQWzBD/yqTTPFZ2rjeYGClyv
bS81wDy4xt2Ru0LUDVapsGiKlfIQGwSPaGaHbIabvwQUBX2/+a7INy5Nu6nr
L1SPuWRS0Hpa5lPFcY6++clAG2BHsQfpR3OlAubO5soC7a79VKRddhPcNmn2
o+0Btc3B/FdgkF5qnO9mRiJe43fM4LNb6ZuDABZBTrgnf9tLgu9xWs0QIBzf
i5WOpbh2eC/YD/cEKvNnAq5Wv7HF1W416uHfC+Ws7rze4VM2hWEeZY2R0S40
VWz+NfD8j5Jz8yPFwhPyuknybmynoVjL8IqJ/yRE/XDMYfkHxUkHrbUVPmHQ
5W3NnwUg84c2yR24ChVpm5RLoLzwSL3H+BcQDNFhlwNOROxe5JH2gJIPIf6R
CaC8/iruNDne6YO5K1xqCbJPJVP7biNs1gdKkP7dzpAPE/9FMljCSdJ2FS8l
8iMNw9IZGpXpFdIJWnBgcWvpkqTVYBPwcp9E6gfL6NPMzCjNdNaUfDe9c3rC
RELUSoWKf3Mc6/0Wm5Zs1HJ3ByEU9kDogdxxmo/nVNk1XsaYKrCu0T5TzpU9
2xBdUihRO+6ba70tqqOLVHCxRbsHgYP5J5pcJ7vYco86C18/CpSvn1jh/nH2
+lP64qAG+Hd8v9CCTms6RRDOhPqGCtFHH8ZF4fNS+dzlvMdaU3NQW2wt8ZYm
f9Nfv+SZRKgPx+9g64ogGUZXY0Z0ILeETIfShrXTU75KuXutV/mb1zZreQMp
F6hFPzdUnvs/oOJD9R0wYILDgxuue11piMdiDhCxLSpIQFppGLLpO008yB7t
JS1lwXmkLF275vi+FDmnktx2inEKG0knTvi8OLpN2FV25qaJvB1TywxfK/j0
t72ScoS9Zr3d+l4L5izOwC/YK/f4OpWG+WpsjMTd/buEUAlQIRKdwGYLkdll
rqmd+UVhHGq5roHhmFtrCGTVxam1M37jMirRtuTn4rmEPh32htrI8e7slWe1
0WYbRYOST9iqhuPcW4h21FhR1nlf47xmYmv6baD9w2cB54IPdJYhpI2VYy8U
Rx61DL3IZvpXW/RkwfYdW670G8fRCMghvabBVa9M+w4ORo5J1Jn4ls3yA6ZV
TaYMbdlTKotti8tn/lYHbnaUbSURzJl7cus/JjColXAEGymeLjrxJzLU9pCx
OUkOSQrVf+CnEyAy417lMbfBc5v4JkIdnj7ZctB85K24ksn0QRGHp9+8ygKL
HPj6ceVy41dMlOa7PfT22PQvn+JqC568XM3/Ma/SbUf5iRIvm/o62jmNaZO5
aeYQIy6oSTa5GDJj+qCdAwXIjkBX17hgPjVF6UBc4EWxdjdfkWM9XVsLap7Q
SMskUXQ1ANhNn3JOTkTXw+KHjFRbkEhAG1FbOU3tyKNpzsF7NHeuDBGBBeNy
ciiA4C6meG/iXKHkX/7ZXnESypQpEv0jiG3YqQLLyhnXdZ87jWpq3go0gp3a
b5a6bjHQ0sGNwgkq29VHNqVPi8rNVRqY/1neGc31T2R/siguJIBZYnf6UJ7v
ubQtrTPXV5bB6a8r3TifCyGXKDILV6IJHbhVfcVVdcVuGdsQ+UH/MRCvXCrr
RIRihr0g/2O4JbYLgtpm6W2rwL0jIyBV7NoCRvu4nyXZG2IAI/0q2kqHZr2U
XiKEkP5ePHp5PsjgvClRkw03bIhb4UnFINXGn5v3f0fmmhqDesRbHBp0f2PO
1sVxrV+sIf7RdNKaajiGMZMYxTmwtnU7w4Nwiu+AbO5KfdxOe8ghtqxo1L73
3NUfo2qE79hZCoCWH4KA4pT4nbmiCAUmGMEigIw4zOcDvE4Ly8lttWgcL22b
rAhkGAqWKGcEYGQSBZuO29Ct1oCXf/IUBoDsotHjyNsN78K7fHP+ltgeBj16
mERGPcZorIPAK038lK8UAbzS1ooVH0A/AFtjHC7kFnEyF6bhJ8bLFis+iQ6D
P9XwMvNTJDTlF2DDPoSKpIBC34HkYYpJlw/xx4KPq72N9sf6yBgFarKLErxh
l4+Zqz15WJkb0e0inm1Uv9xrqM/2S38M4h/S+2atnX0dmjyaP10c0ZhdyWoG
7JVHlqcUdCrUdiJky8otKSi0DnCh6US/4Gce54Dr4nK42sJOAF2Nh9MwZG+7
29qvNuhihSTAXpU8OGlgGSnM3CvMyq97grbZeev4JBEQ1nAHQX1Q+VrFpJIN
/siEH1RdvIzGK+iPc+l/n10oquFwGUVc9Mf/X1b6kK4YBG8ZPtA7o/WWRSIN
lGYosDguaUlBQ1ivUdvr1VqcIaW9XWOx3wWlrCOoEgRO9R0mOTDBmtKMeMxI
Qe5atREo1b5kAzxdqg1iqVEPir1BYR/wtbOO/miObybKpvlutivKagg1VNYn
AsVl/jcrf2UDebo5/MPafdg2PT+Bu+rpxJBG9EHXGwCxD40j1nwY+0WBjFTD
5vlzz6+BU+MavzGzndTABsmCfAXJcx3+AxLeN8usIAyRhjXoT6xBuMdjVJb4
44RA/lLV19+8orzUbaFlLSU3BXQ/qAIQfrrUHyvT81gRUQ1mSed9vOSS2Uxl
r0jKC1U7orsIMLanDqLaNkjuM4IrXD0I0ZgMIxmYJnPN3zUqra1BsibzoCyH
2LHMjCgyjXbKDXf/u0IgRwDyPqKrsvIDXMWJo22gJ0kcJHXKkgdXdFbqKxDP
bxKrPLXccMPEdBZG7uATUCCA3Hc7AJX/kw/4D8PlAmYItNePBiWAgPxcLYqM
YPB4cb30pVmH0NzMSwup6V9DvD3tfVx6wadEzid5SP18Yiz9rABb5UE7Osv1
5e6iZeZOIb5Z/YWpF2aOlxhAZ3lougv3JyTdqd7MFrykZTIZJisPWEvLY0tG
fJFRVJ2lJEaqGxyDgAqN2A3IJAk2BkjRc2jjzFhEwPSH1npk3YQTxC8B2z7Q
SnRxrJrcyp/aMrBIJpP/PcktVVFJ0TfkRY5AHneoJ7Q7WayvZqvwNC/2vl+z
0gjgYivDSWQmGC3DLXUhiKVUUjJpeyUJKgwr7qJKxqisGCYpoZW/3kfyeGsG
WPF/Qqb6GnwhxWEpWtdWxVchO9zczG0DYCB9xG66oxDSBk2bVtY297Dfpyna
9rP/S9oDs01q0g26AEIIymcMjap7RuDFQL/9XaiQ6hgJbMLmeZ0VYgK78IZR
3FnckYeCP48i4JIAr+AmXTbIHV6UysvNOO5bCCF+V/jH1ZkQGVYFa3KKFGHC
pNKmctIrdma9RqEJMuOTMbbaMravtkhDw6J4YLV9cURwFwTOROD1muAQMPwE
F2FJszll2a7nFLOSB8j7f9DddI+6DoCUXJ7wBmnXko6Rb7KNnoHk/tb836+Z
NN+vIQfYOyQzzJqrtg5jFwP/B/lNSQd9yAFI78PMfePOxFB64E4X96NaQUw2
yvXGCdbgzFAy4QU3/WTmCMVeFzlISMqux3T9U/h92ssWibpnzMDFW1Yr2W+R
305d+yA/k3vqcJr4gPT9CqBui+HBT7uj8K+REA8cLtKwcOPT3P1dZ4x/NTNR
o4Fzf7m4JpEvciTmJtJo+8rfBtXz7fCT6Pn0ZGxfIiTvU50usi0IxIkZ+IDK
h4Gmvpah87YJgCTg2xIey1LWMdT6pgNx0dZGg9FIfGT/rXFBI3XYpLrjTQD9
qTHz+gt9vr2J+4H41oOqtBn45/GvuhjOJqVEzh2gnA0JeuEnt0nyLS9uKxKY
EtmekuFS/t6x0F6sCeH5vYJBGMUdy7h6U6M1OW5dUTBs3HZrQWQCMgOrrKlh
zMwL5w67TAeMEpQxoYXbQyY6+Ob0HwgITd1IGxc0oEPVJphQLSggGHzrhm/G
Nn+UX7egu8I07ECNTCOOn01DRLl0Z9zyeU9n3+U+bPBnya/+fx4mMzILeFnq
+sopbHWp2kcvwBqPzFZz/OaW07NMCh2vdScLIvD6Fj08QNoHBMXJ+D3jDaOs
D/I1f2saeqhNA4HefsocGc/vM9lvLbDtQb6yN1SizWxP0YCnP7wQ/O6/XI0E
We/cVZngMjjVDyQo0hqXj49lxqB/SNKwjcea2cjSUsE/hrZ5d4yEeJi+7Oud
iA0+wAMnw5Bi2V4pZcqRKkk16nrwM2mYCThtm/gylPGwF6GEIGXK5lG2Nx/0
KJFufJje0HHSmSSY0zGel/HAR3F+inJgVrViE+f1Mrp2BgXbx9mbU2VquI8P
Ch3XAN3OnfrCYCNaCrwQI9tH+qjMR55C7tD62wEfly1pOSdffBI9wVckdJVN
AwC7SEUimuM36saLXBI+S1sW6xUVkSU2YIOdTszl4Hk2HD73wKy20oCLJhtk
WP+O1EsKM2nDX8/VVmhKfNjOxXNwnJrSxJZBl55VXQWZ7wbjnv2/8UEQh4SN
h87AYe9EuDAj70Mjh2B0I0zWi6VfEQ/e21HmtnPMhWd8tLSKKiIUuQiF/B0c
eJkLnSb+V0gLtF5mmuMDrlpnyCLB1Z8fWUUaDRamq4hH36cam1Nvr4B57Msz
NGwS2ml2ShyKoB8I9CX9SjqSXB35raFYj61iKcOJ9LTIO20mo6MnsoVuE6f7
f9vmC9C3DOrVH8sE6Tp/Usvf2ek0ocXpqrbnu2DjEMFa6oi0BmRobxy+aCXP
JHVS0XLDlKeuSF4Y7cvuMFIMAqNMqoa+Q4/QvZTFay5ehju8BrFRDpKciN5C
mXPqBQare5HisITlY3NtXl5VGQ/HueYafG6yQFewyZxEotKw66r+yULylvOR
yIg4KdCFWlHZRMxrMBhlenhOWmYR3iX0u3wEZ5P75ea7cMG2Erg/Lr9Ir/UV
yVvMi2dknQuH+UOVi1l1UftWGWNeESYvGeMqfkRToYrpaSreAPmbtkjoOZ+p
mJSKG7NJtX7ZLuShOVNaHsb4TcftQjEO5KZSE7gib9sq5JzaQgpjOD/n/8BN
9Gg4Zn1I50bXIYW93sOH6pJWwslGzwAeMxYwfY1t2yv+h9YVXWMaUkdU8nlC
y7/eFJDw5GzaAmDCMxiNAtGnx77ybMHBolluL2fFrpxyRmfhzSuroeEf2ElK
h6oEJ48rKLDOsNcKTujzg68A9yKxVQy0cDg4ndzlr+DDq4zoF3bhTcUlS5dW
L/Nt3bQhoVX70V+qQd6yUMSphiptphtTR2mE4fE5BqKF3ZzCGfk+84gDc9Vr
LFOr8FIy03gd6aH7ZUOgiTYrvvqBBOuHko+C1atps8zqDjCB66s1qxYxrq/x
s9MyRO6+QQCTsTGWu2Pg4agFso22aDVNwnz7c1wPN6OMtvKKAYtBCnhoZoRM
3UF/caat/AF0oLRVgCUoBMKpF35nyEGtmJ0qguKldRhhUhDNJniHXFSMh0OT
EFAHvq0Kkb0iOY0ukMpvXhqHVXbPrT9+wwkCd+6PWYicvRbqcFFLxkYTeTkd
czo/pAIm6fzlz0q6G3wMiAVWNEwLfZKPb937fxhc/O1GLpjyh1fbKAqWw5+h
a9ixyc5lrpvt4rQyL6RSu5lioeY1oYS1sGOnk47AmFNm5OqY1/lOVV4zKvTd
5r9tZurvNO03lx66EQZxrN4PKYpH9osrpfNDbD1l5TqE0PModeAAliuqvtBr
E5HwWTztEVYgoMJ6Y7XOfzHdxW9fTvPZQK03GuZLttORyp99yn9ojuh6+Nhm
xWilDD6EHNHmRra99WupDf3rIIJci9mgwZBwIwMTDj/O+sKpEHFupxTgh4id
sNlan26NbKHEPUXuZebqlJ5LtGz9kQL9wtTtQcnk6EN1yKvVz3F6P5VWPx7v
CTS7ndKEpI47OZuMVreA2hqcGyrlUGJl2xHuVzjlzZkLFQR01OqIEbOkK2LU
WbMeWkwfJkTGXCojEW+NkZmghxFx7v4o8Ozh7H6RXkVd3L0XNV32l+2QwD1x
uvx/WFKhvEY7/NZANa9broo0pgWJank1zz0lYoViA2E82/ou0roWGqIBciCm
rOhRpfpVQphT5LfeyySNVpoRrpwXZBAbFfcG44EZ1rkCL2pJlNw8Y3Nvtbj3
f6p8TDN5ID7HgNeOoceS+5h+sBl3vOgr7aRjEA4hp2ZYIr+4lUbPvWjiZ/Y0
x5tnmtZQX+pIw8ghsHObn777VvkGiDWRjg89IhL46SMKYhyAHyPvTFvrl2Rh
LqPRKA2GvrxZ2XfKh1MRXjegB1pFWACCCfgDCVa4+1d9xmFnEMR2ExUq7zez
QPK3UO3iCbLVYhcv5kB4YCaxVkV0BfcC1PWZyy2D26q96cnUKDt6ei2VOxJL
988Ni0/SaXd6PdNvm4oOSDTn0wkPpFpj9hxGd59Dt0NiLPmCRLBIruaNe/TF
K5I/DDj1vobaDpeHqevBCjbZx2joPI8Fc4yPUH7TtigVa27HV7ZEyZZyWNVY
aRO8NFBQLhQLrurrELnSTb26RSMtll5WSfbpHbXPYqKq4AZLAnczUDyo9NZ+
+hajvgn9JdbgA4zekIEJy6mDjXgSpcO5PhqtS6CquNIRy4E+zRdij9ao0wya
Y487G+B1VTxGa98Ib3afejYgTsCuCY52IMmLu6exIN2UTUPt2J8S1f4BwAbU
D0AhkNnZ8e/+4X3Fmt5/F4DAa5h3lysWsY1Qo1JQdm/GgqGUI3NE6QFb6KQp
8HvQ1wx15ouch3ZyXRGZRbWWGhznLt0x8nqJNFhiraQiwQyUufiE+J2+GTN1
Cfsn0kX3vEbCsxKM0Mgnj6cicx4I72n88OJWyLGPT1QnTWmyzL8PJALC8dlh
HelxKRkwxOBHvHSxzTlBThE9TyERp3rpqsLCQj5GtH12+o6sEMrw9g+Fh1+0
HALbS7bh9njllao8Ga3Ss/VP2FSQjaJfQEikcHSlXau/kPam3ePmqzChTxfc
Liv8y3pZ0nx4tHWWQFaUabT2s26nPIrHgv8BsuvHQKxv2jth9IgQwdnajucP
bQBz1SsWb5uthEFgj9gkF0jxZDfZoB+ANxqbeTVvW6R/AuHn7Dhwan2aF0jj
7PQgPNhhiJT3VXhGlJhymIqoSqAZN/c2cPeiQpraN30+XibfWYE0CveV53By
duW1175gCtTzozUlxH3+A2Cp89K6OO8tMdql8VJaaFvHdE0RwhY930iijUEl
HiANOBcAfD/hQWrRvu/rbvm/QlFafp74CoPO4IWJ2CyBphY41Y9vDdSgJdj+
wnImr6b6a0rSRRSoGe3NtapUP9d4d9dh5LLlNB5OGK0B3kToE2QNU8d4Ijt+
J6Ts+nQkaoZ6UPv3re+xAcVUwKNYRJp75V1V3vDDodbZ5yVxtNbxt1lVli+Q
rVtISqreDB8vua6amBqcau+//sHKVjvTtAGeGdqlRnv1OQiTe5VUzd1wXENe
hBT0dLAO7/Bqstj9dQT4r1T9SKQIDXnlpi9cr/tKip1wtop3tw4B88LXJsCo
bldjzxa+UhzRfmYQwsmtOzsQnHBmzFCt7Vw4UyX6ztZG1/R47baEQNp8OqLd
Kqnt7d2Xi18A+eKMTkro2DHSuGR75070xZlphz1iHrzJPB9Ieal9KtDbMQEN
EpYm8zX/j5VYdr4pCurTAe7BlL/XdleIXmFdGfQuuW0fJAb+n0LV0yGzh8yx
aW2fzEw5ayjxYn1aPS4ZbRYg6IWVQJNE2q5P0Jz9M4VtZY+YcWh9c0pqtuze
yzGY5ac7/5ftqZHyu0PtP1mGUqCHfopvSXgPIWh7sW6+FhA0uPWhQFHEZyP6
llQT166T7GRPWCcLPOpYxzjyhGcxw8bBYOhBI3RIhl2rEMFvS4VzyxsB3uM6
Id45CRuVCrcK97i0kPZXTZ9lzN9bZDZx8EnXcf+MMjevyA4aEMntanpg5VpJ
c8sfahoVFnmaf5tLN5uapng6wYwjpA9JI3TZUfuy7VKf0KGzoPMdCLpEblQv
kcDr6Rhulmje13HNHkc3c619ENjYPIRYWTABuxdre9n5IY9Il26xoyBCqJVD
guCAY7zQd5iTmxvmoDiFg6fcBuUG3Nxzb947gIMHDNKK/sMx5eazOb7rM6j/
JpzUgK3en/SBL/hfQ51m2GNoSwtoJTOteXhPOP/PyMv82UrZ47eK++2TaAsZ
eVx7Pw+50pKHp9EBQZ+KwIEUwYBwHBYc6GbdwhvrQwGQSAJquD9xdDu/9qK7
jJIA5HxWK7OhmG5PFLf1mp3DG04nzdiSw8O8dVWcF3p+5dqPMz5M5IDPuOEi
bRJDD/ESJsPYHQqi5HUeccdv21Fyja3CQmlneot62AEbgD1+rN/kpUNQ17Ha
6e96qY21fa7PuNTa8QxMVzpO4eOkfk/ujMA3ORYoQiYqmzEJji59g+wDfia5
i/m9GinJDU3ZuDXNHbQ7lqyVs01M4Rh/mb81UgOIkm8ulV/lUMC3pXACk6U5
RoHc+GX4jYSnxqKgPGI4H839GEvmkBMywiy1c8QlKF1L+tGnYH0P8fXTgJZa
sIJvI/QuSCUdO9K7QMDUd+Ag6YtizmTQy+fLiH0f8Zhy21clE+SEEcb+rK0Y
kQNN17dLas3EQztWw31546on0JQt/RtZVldiM+h1edi7lN6+Zl97M5+rmRMx
NihIhUVw9I+kH2VJySKbjvtjNTZt7zHnvxbq7gHGuVP+0lsblIVGfk3INxhS
F+LZzazcTglsPPbDDnZN1rpdUWikl+QO+PfngGrWUtdxF4OgexN84gvcsWUN
gTmKpE8uYg21LLFXSluGInzO+xnbYQeCPve8cX7B61B4qPUujozSzpY7XMEn
J/dO9AleLKDrId8r8y0pKv1ar1/HD2Z+XgoxVCA3ubidD0+a1ZufoVcfBHBZ
kwTbiG/VsajhVhJpVOpd1kGuExqBDWPg1MoApkxSfQu29sH81xLK0TCLGf/C
jMY1ssUgDVqEU49z66lPX5hPmJbbHLZQgSTdh1vohCkNUhFsgJWiHyDfkdIP
RxQ4K+q8pbaMv2V5UTDrHByvhIYtPK01oCOtRawZwrTPrHzWa/cWgqjLwKgs
cPqYOprCUkQ6Qn7wGlkUzU3iqkNKPwxSKsj5VNZLcex/WumM2MgttJ/TKEAF
KoOZRV7x4NDXOrFV1vBNLTlztxEgTFHpHnX4yW7aFTzwPi8NPVsplhmLEl1D
VgGweoIbnA5AKc/o4KxFV2/x4N/R+zIouH5iF2jIUcU2UmsGK99fm0IuY8Ca
96XyECLDQH2rbDlRPa2+HcOuCrRRTQvibPR47T8xzfn9ubnknZMqkmnKN2rT
ZB5gxJqYsx0ANvHtuIfpXanyLFnnhigAo3aNBNSOba8H5OgkS1oW6DkRWqZ0
fcrwe/qFPoNjs3P/6aCAoMulHfmhrDjz6Wi9RLzRCcG8tq8qMP1bqYm6Ppil
6oG0CkDJ3lZ9mqyHjvaQLVhL9hAFtvxl40HtYOQb9F5eiKTVUOUNmPhameh4
blAGXFKFiddKDkNKddi6WF3y93xE6qTBhemAui6QW1A120gg5ezXOdo3+838
clXkDX96I89Xp4AwxK4gzfGLPbpqXgukaOSFWCVwPPymVuFnpVhmjxQkUjcd
ERLc+7NKpLS76JoPLKH0JTrSfReenbg70x5pFNijcs6qCzZbsCVerK1c4ztk
OyjyW9JPwaJ+qgmJxHGOjeSzn9jKl57OLc84CRstS6S5BUGAJYACNTe0tEMp
VDa6GljXDvtRmS9R1IfGuNHeTXN0FsvJFVpyNUvL4mSnFNgUG55sxhTpbr80
rb8DwPUib+nALJAzC+p9ET+tFicKsXDz2eFNl84AQCNrSK2ZE6NeDl3eDs/u
/LGQ8mMQglxpqQsggYjEvuF6uAMKGjMSoKvQ3GVPdqlXzuXuxmHcW56fatXo
XT7V26i1W+lHT/iFnL0aco7jgRApY/V3WUQLEOnDERGhby2yukiyv7lZItJi
tgM1wnRSgb0nCl750UCzY9EOactXeVkZzyfG8ZNXvX2R+KDCU5z8U4P6hePU
nDgTd1sEdb2LzFvEyy3yKGz0lXHWpLCy7GK9SXbHeRXqiEzZ/z1Ni9HELVvC
Xgnsh/o43gCmZOqvLKF7GWm0sFSbx3hJE1xLS27CXjQ3FAoEA4wzXIcmCfcc
YeTaw3f6VqxVhPXI2SJ+XIhv2zPc3NoEEw+FQziszqOlMWxgKdqeeWZ7Mnup
mH9EEOK0N9dTdo9zzHKNqROGZzTifaX1X9UCVl9DR4KAAWDnohcnT5GJ7iYR
vlxWBCQbaOZKsPuMJ6KyX70hhUQDZ1qoJWvaBwG+Vwi3jQuRVZK0/FZaphD/
A7nZrzv0KB1uR4T3dvBUrdv6xQgrW7g2ja+5gah9KCE4a82lvHZ3k88kRDoz
uR0ZRrZjj/ToaUPNEDTl01T7eaewh4crOl1HjHqmqN8zllCr0uMv4yw9qz8i
MReeif9GsaBzCGg+vPXH1gIVcGeqKw9xZlH91SAt1DEOet5F1VDCJAVDE15P
t1mYq7zx50fMvRiu8riMNF2escU9pcdmn+NY/D2EtWFiEEo4MK9B+EwLX05W
F9rNmC1Et29eY7Kw06bxGupqP/U78sP8ycO/8akN2K6wXbDbyLj2z0KPY0PG
yHMj1f79YDX9TLuWCQP8chGkeCjO6lqaxu+6cO1z7gyTdO7AZVyu7EQXTM0A
fQ61XwkxCYrOAJAhVGen3vvPqvDDXWFPgRfDycyOoKB+/BU8vdC4hfacjMml
QQMlqgPlP5kSQHAyu8EKdwwx5QtLzIrjDPaEb3Mzie46yEithitmiVi9r3dP
Pu0gGCBV3eLegpKk7A5TUCR2IQ8Im5DcN1mdYxrqmycGDKxUGb1AQK7lRxzJ
2D052UHcbKMYLeWEhzryDcKCxg7lasaiKx8EW4ZkXRGt5GbXGf3qZpZcjC+5
zx1kVxvMc/WY7LHxVxkjWWH7Y+6OmFH68y8B+2t1p3qRzLRauZTEfbVGw42C
s6WBiEzrsttbos9tPg4GuGGT/qc4S4RMJVMkudz3HSFS9IgfhzFAS37ISbgJ
BjjIRX5tVotlI1buGcdf9mskRwOxzKIpVt0u1rUm7Xj8vYP5ycLCFjkrjGRh
TNHzFFLTZXLByrVxxP9gOIZYPnmEB75kzMo+4xP0O99UKfXfGwl6snaeghIx
F7fsNuNxs/kh3eh3nG3QNFKWI7lovJGj7hA/U3+dHhNBotE1R6/yLw8b6KAV
AbBpufBmUu+QXFDq0g34KxAb0AHo1CwIHR2RZnVx4Kmj2YCXHwI9CCDRSZ6l
+yHI7SxJZZF53rAKIXieIC8WpsIHOUcmVW6fEuvs2vlaxVjszDfamZnmd+vL
9d/bfbwbOetx1XSWjhUeLoYACQmmseIyV0KA96/4gmw4BUu/LLwyQkWZETr7
Iy1FC7E6fFG1m5yWIMfVCaDZFgt/lqkRG5cjShqEV/tdP42EYCHsX7osZYSM
qqYDsq7HrfZobqVTbuAuokWgrCNh7d1vbuTrDVPJyRnq+dsnN9PSSmmSyxea
ERI36P6Agh+bgpUQkins5RvB/Z39/4PHjVgTmHzaIpNQBzd9e8J7zz03ZcdA
KbYIYK8tKKvzyXFdDNsAPUKDu5VWwvRJskzf4dzooAwZgegUZvcUJ34hrU3q
JKoO3h5Rzj4BsTB1EI7wj/fhz+JgDTWUxFcH0c+F3LWPr55bn8wOK1fZCeb1
cQVyMZ1mVQsBmtrQa8/D7fUwgjV8QJOHyG438330+SawHOkNXgtDzcL8YIhc
nYE1k5KU4PVyeI+hHBFUzzpm/TITxE4jvTi0W0bqtCNJ2VNlXNCm+UbUWb6v
C1YKTYnPcBwQUeTHgALniMLg0T2zQy5cmG/3dzmBj72kKh6XpJNbzttTxAE+
xxn5+iheToMnOK3e8GtMYE5hnGxhFIYiofdSJxnCE8RkDZIzMqK4EynCCz0N
JbMBhs3kEFgvNISJZXtiPfBfr1zQ0pdBBZm5uWiU1KMMH9M5jrG4Wn/QHI8L
wPYaDAfP7FN9w42sZloG9eTZJpMyC6EBRulFUhLLDzd61cPyZoZsfwiod4Jc
CIYGhbTHUtjHXgE831Cw0MYwMYFsqVTlJ3g7cnsPSmVKz+ZOKpqPjyKR8ofa
9R1LJv7ZYyfcpWtw1k2Pdfcpbg+86CA0yXRwJhCbvFl341E66vW+PBZeQ+vV
rSYcUm7Vf6y3TBzmkLHL9EcnIN6uhOVIOfIlRPjofpoKd0qF2OiUCXdmlquj
DyVKbJlONA0dYBjM+6wkzBIm4WJHWW9LgutdsiwkZWBbDQlC7t1Hr8K0IGp3
r1vwQ7H28TJR2xoKa50bH7Gn6nlKQNdeFhK/nWlBfR90lpy7tq67B/fgLCuM
WQNmbQDOnUAEehQDtvAd5hh+ft2998qxOliADl9CyGC3hYrN/zWD6qiQ34m1
M/TqxgwhumzOkec9VKvqHLZnEBxYkDzR4G9iUFovVAWVmce1ujVF0kYZwOzy
kS8eBww5XfLmxAKza07Dl1DgzZL0XqGe6w+hSLYIS7+2pwne4guI+G6VPpAq
STIo2OJZF7YxL3wiL2YOLPIrRxHM5GXUXioY3t1gvw1FFZscn0GlPEL0GfSB
MzGUqdtPauILnMWyOSP+ZkI2xxJMoNLG5GkQ8TwOyfzwW8OwkTYdDpdGE94c
GZt10l0d4Pv9HWkoHEI73XKk3TYdyo4UnayezcktSIw4d88zRo56oYVQzTcJ
UU4Cn7FK176GbpNP3gJEhoj24cB/tmg+H7qkRwXyZyQymOILfTcOg7E+iBpX
EFkkkLfbaOt4DaNj1NhDfxf27bAM6fN/SDn3MEhDNnoz9GtTWOq96tluFquO
sH/yLy/dJJw7VrpAThGg8uS9rd6r//wTokAclnHuEo9wubC1mWSckyAaiaWj
1DPef5lKGWYgep0x9ewK2xa90jV2RqM7j23zh1YzekkYOX0xB1BBm9xRGPib
J0yJ7pBJ+R7W8ceO2TjDI3Sua4T9BgTH0jHPyUv5keJm/E2OKTAa445aRgF3
XemJQQsjmHVzX5VgVWSwGi1sAL6KbD/SRZkZY+g0cz7Cg/sFRCXgUSu4K85A
fwENGIcQ1+kq9gOh7UtVT/pR6aWBYxbfkQ96y0H9OIDcVKsbQm0ovIspr97y
McixxA+t+su47+yMnp+KgO5yKFFhPzrEFbjwMEqfZCMQVHsOWb3zMNGH9oAz
qO0JQz3zMeQpEhecm5zONhxc9HQryqd6XXYNOMgGQlGfwl04bI9Y7vM8n+nq
ytgoz2N9OdKvk2QjrotTpYYSecoTR8sbyywoB21hTen2AKrFWiMlvqyOJ40o
qwDhohx/nPSTSa/xkcAG5OLBdNH5eYnHa9kRoyD1FjutPk/5Al6/YxFj/GtU
vUzHIlTqbH3Tl0kv8/k8ZFz8V5Pro+iF8dCyDmiCagBbL/X86+NJQIW1TjnF
i7kDubhsoN71ec1w/hpeMDlhG2rg+oP2QeaySL1VPxHNyP80eTfIMlAmE9Hw
ani/73PMCYwCz2aMPtQFkmz/4s4wDqiOeHLglihkgRrVkMdcqkz/ZObAVQfx
Y75oEGKxgbm/k0BrSBpks9mBMTv7m4DNEo+9Rbq3QbBdX5ZOxkw3DvhksV9U
Faa2x0MMFNFh09Qh2q0a1oyFbb7GPB4NmS0MIzros2xwH35K4sHhjRNQHqe4
dne58IkbLfVwUymklVuybilI2TBr0MPFjPZOOmZv8G7tiLD46kpjWOohdAhq
k2LU4B88ADxW94L7hV5Q+ZsHIKoHEmaPAlZF+mN9KF7vS+fc9qasjC4ZbeiK
8+zHz/9QPKsHYPosJypUIj/+bf9IoEqQD58+agZKg0FcSO7E/+eW7nDms5XU
bIWJdDdqPzVorWr1+O1gBDDfh/+dLYA+/Afo1UQ1pHvdN03lukntuQRqiBqx
eZsiSEt3vREOQoV67YYfek0cxd8LGpaHLt4jkW0okMq7+8BVmsyO+sP+UNGG
W+0Ul/9YaPjGKPh8t7uuYkFbx/DZQGt1cTL5w76npChhSamwEzrNupxCZX5M
ioNmnfptPwjIbXeokYs9JSXWJcxonhKgpVKpZQNAwoT7VYn/lWRbNJPdHo5z
4ua/w241DD/Kkm5HOUd3QZ2UrQR5bjPR8KKdGGGVuP84afSY11bxOCsgf7Tu
L/wCHnwCIvGP5LiOiNT5LN+yAKhDW+rFVPpR8c6nPoP3aCEyklKI6PEy1bp8
0c3KBG/FldBxDujzThNNEKR+ikIk9Ex0c0sanaYVqHjTM49gm7snqI37Iijm
cEXPy2TOEgXBqtIPp/cNH3slDKgLQRWwdXsA8UbqqgceJg/uG8HObD4kuqkP
jpyiAJD1xI/u0k4k58j1irY0aVlajFUdhNL45s9ezLNP9zvROmt9hEiTj9XB
y2FQ8EuUECLWi9NxXKGx/pci7EdU4UPSAR8L0jlVvnRnIWk3ZRMobqlD6de2
FUzAwcSpc45A61dTWhflBNF9WvWIY2wpleUP0EYVtfAsDEgo5Ou+lhWvtJlO
uGy05kLm8g8UhWXa+DvacYbBuKPjVQfDni+rSrSBuFwq+jWStdo2iyUNtmfY
JYAU4drjI+6kuW0En+h2VKnVF8UkoluLFTUUu8Ef9TFb18tYGnlRIB1YL2mW
6Ugp0QcLUuNX+OoZDulUfLRwhqwVEXkPVVxfoKCGljcSf/o6iz42gSEV6vEy
ouqbp4S5OSHflKm6XOogtlX2hBsi1F/4GyRxh4DmDmKS6XuznzVSVV74zng4
+HfNI4+O4/p5zLbhsynfJLpgKMDKntAZ1kzBWzEgYd7wt4IiDUW1Nfiz2oli
Y/Zi3BFYncgNia9H+KzbKt/PVTo6QiQslEPhzny+64FI/zsuFotO9bddjA2G
5j41Eh02uDENWtGFtx3dDPHg2Pz/AhOKT3xV1Il+bogA+f3iA3kZnGxQesGb
a+wDh0UEa+F9eU6O+P9G5+AqaeEMMC9DmNxBJ8rBxOKLxKW/TBKw/sqcuM2u
3Da+uk2YivtoU73lvYa26dFkL8NFf7M1tNX45xKqfOHl8CQek0n16l3I+gfB
QeoCsQDdrGino5t7dC8uPflGcldy5r59f1+4SSetGB3EtQjbTDkR2yhdYrPD
AbBJORyRx7yAou5cSx1+ftWh/aewkk+JUl7T3CTgZhYrQHAHNhST4nKEMPMM
szIZx+IKyVjfx2WGgpwtVoq1O3PM2XYXt54ZgB8jKUVLOp/klW01zpFHyfy9
lTBqhzSr48URnKK0qyN8oKN9oBg5JikOayCt7HV5Aj0o4prMuzcpubPgMKB3
pfCgiDOzxx7gfvydSCQynkABsPaoZ3nmykD+TrsdOmUEL7ynMI9O9dKD/Flv
EZW+oCQyAfLHrRjylJPgml8gcd7eqtiLUxz2dQmOonSmjksth8N96bIZZV+Q
bAhCjSfXbvccNxvKMlFpTWI2wo3L3KnQsxu/6iNAKPNhneexE6gWmjjz8dxv
tzQ90oLbhbpwGCaft33htP3cB/hsylKxECOIaheVcox4DvEiyADoNUiJ6Uah
2ZpflCi0lbJshgZqfOMUrnccDyO5e7zhjrmaKTCyj/rxbjQ/Y125d3kPrcDn
fiWZRko2v0AdxQUvZg4U/bJT1bBNtt9V/4kOg4hEgXRKLyEBJJhkyU/gi9gT
FaDH8MoEZpHoDy38IEXmqUXCUbNM6cMTLzpYO9RIn+4AGlQQibLketnGv18Y
AItLseTNgQpxzqUk3RCvVIXKwhbNqG2VmTZgWuYMPlwLH4oiNftMMjqGG+5L
sAieeCrG0fC+eiqnTcoxqoxUf+o8exs3n5j6kWJTXgvMXjjsozmrg9ML1h9h
Xd7pZfpFMDVIeVvYljHHMdlfTmMjwq02d45cp67vcuKTya2JfrieRP599Onm
pc+g5pgFoOWHQMEmxazgllpUMDWSOsRrdZth85nkutQePbrOTWCkzZldRcTF
qqfASGJEpoxHX0u8kdoSQNu/4k7ztT/XuKAdcElf4uGfHjcrjv8m/rvwgEp8
9oTjXUfyzPPtpXQxiCAlO4iKUuGpwKoiYMfEmkLe4uNSQhTiDNj8i8XR/yHr
4nJNmWEECOsOoLT8fF2T1MsE0zdg9sLH6zOeyuLCrggAWBKBMEXcnT7kZsYN
0DKQsWTH6Xe/W3v98CaA4lEbfan+Wfbzh810Pom32C2PoogXascRbLHhxPMQ
FQ21f2/7SkkfwBqyuuD24uGITx0/t1n36HQo89DPnBvSyd9+70p7zj77Nr5X
bjxMD+Du/49Clp8EmFJS/2uKBaZY1vMSTpgpl6qiNLqo9OCyrZRCFnkE1Smr
EpTSrGD//K7UTFZFDbCptwxcWAyHG6KmK0U1ZAyCxjQjvCVl64JJfWWDzjR2
cJhsxrjFK1+MxbrMhOGNvt/SqDpLPxBYa+iwKS5WTwygFDQMKT8d3idJ1y5l
+2gC8qR0KcGv1+ghfrQzwD2SljBaMYLSoTHDfOs50Z0hhnKafK5EaSdhr/m2
4GcFPf1W/7VWk1RsU0t0hyT1wT87I2Noi+l5AF2MAYxQen90IXI37urVoN/x
EeZKRAwTMfQjM49bKZ6jqxmEFGkoyJIg/FA6Mv5Iphrmf9bKytwZyqAkGydy
0vTes4F3FYAUilxdvPViiOirY4z9MRtJrbaXq9T27rrGc8FdGx5Ph8EFVusf
8zlKhMrZoBFnlRPCEUjz2mEO6UjcxXNl+suii2pxW4FKcomDt/9T3yAGPUTl
TeF2qyh0VhE1R+38xtx/nHGcu1qcVailaDApYYlQpLmZsKgM9MnC/l24P1Qi
TSeWDOazmFShYvQLpzx9lmBDa/yhQtHPjCvj5TXvHUQ3XA91hY59y44L+LQH
QLPSw+vP1GRf24usFBtpVvY1eqBEJOvaqOQSxe8tGgrjboxuLMxfHSWhUmDD
eXaQSP13huoB3sEXsj0jHZ4x6FXOhYZ5+iYKLGrDkVib6tD9+q2yd+fJJHCA
fs1iNKedIZPAGj3iT/wazAhinSOt/8ferSSLZ9TtT81mbxLPvMhb+TgqsOmG
nfifbaRIA5KrUdZLQGuM+DVKqZP9hqJTtvRTaL3WIdzXz6F0avQk3w8yujLZ
jkJK46DJK/s5+/HAYNJA4DOm9EeJ9RXn79UPOdmvXj9zmpIr6N6Vq/Xubbx+
IrXiXWVmhYz8A3P8HUDsCyIvEDzUO4JdQLfmefFM2itlXMVS3PjhKnGy0hv4
1e21E1dZEOQdQ6Rk6FuUPWCJKm7HZQYyUE2iU+2FjK4ze/yxa1DQBiCtqnuy
2kyjXr4lC44kgDQk6yxWEizSkZVleql7+PGb3JYseD1NP6QkPDKL/yzmG4hs
ZZtbALwiyzNC/3lcjJsibliJ8zJunICQKjF5RNV0NF0+lN27ZVtBtxHO+L61
ZOr+PItl+BH0hqr2Ysdm53oBTWwP8oW86KQrVmi3sbR0byA4XkhBqUuvsgZD
XwISvinptfsHE/4Mx1mbC9GIAAOS+JPIIeT+ySU/1nDppUuaMbDPKjwInLM+
XuKC6grnXPaq0QtuM4rgPiPJAak62IdcOpGeCp6mgkdA/PmGHB38rg9sJ5E/
pMRAU58djO0L2CfgMvUKfosBvZeA6YfFqGGjLjqJ+fhNKlIi7+BWOS2hR4uo
kZMGAC+NRDOcJpDfidDTuHr2YLcJaA8iLv/8Q/6jf+pGTRJSliJNR15blqcr
0kB8nh/cDZ2efqbsGB+cAVpOgVeBL0o4vWmPFJHa8NflJNS+bosKVML2Q55s
ehUkcjF6zGAZ3am1Sk0FdCwWyAxPM/VEBIN7WALx4fWlMc9fqO83uXfW9tFe
fOMlz3gB57TNwyKJtiuoAyy2KhjGXkql0TsBwm4C1azXMAGHdgDyRJJeUdjO
zz5XXu8IsENCqgSLz3PR7iDKdkWg/Wd0Bk22O3oYfWLYjN6G5wWnVCXbde9b
3JoHPB9UACENBKy5gZQaquAlMKUee5Xgp/UK/qrfOmwO1XXPCoAwdVqKA51z
drezpfRMZ8PjrRfjBhEdqJiqn+5cFbV8wWoU0Zi5VQRYksy0P7qFdY9yXNIm
YNDg+yUg0ibp2BN+UrFjJYJCEdFT6RIz8sUzJid6XW8E9EkmZ+GoVkmS84Or
/AJW1wBinyBBigTuReaKHZt9TnYe86cdlFeTUApAnuQQjYXM01GYHrJf7wkQ
EkCBlFx+CErz+kAgV7WJBGFTjujX5Jb0F2drtdBJX93Kx1yIrdaZsbpaZ6Oc
0hpU6/1uVTQnLDp3QlqSZzCDkQX7PChpdc0cm8t/jwxE2rrUkJoZEXNBkVne
ZB9OB7sKGMkc8IqyDW3M5/PazJ1ptlalXxjCdeeRm2yMHbCd7VgP/WUsRr1e
ehqK2cJTo6u48j/FRwtP4wKC+1oL+LxKskYXTW/yP86pf+INc49YcU/Sx9Oa
CC3BdjS8VjoeM5JDXt4iyruC/t/jCv1takFmHOzvs5GpQXxKFkaeN9ngF00j
Ql2B/w92fc3uzVhDb6VyUi81qp3nbeffDBZYnw55TSgt6DYEvTK63FKTwvpt
iBaviNqBOXZbkysf1sEEXbgwoz+3JUlofaZYvgUJ3ivDQiZ7d9PhYkwI86ym
89V5BlSk5hLovagS/x5L+x+1Fn7HOK7IKWSUJBEv2U6eIxePnS+Xoo5pwbi+
zmwFXjWeP4A8nFTjSSneLp54zKeTqKhc6Hq/oHNQL3s8PTTZCRr2vWU8aD1i
MrMUhdDFJ85P7/3LGRnBx5rMOGiYWiJwL3c8OIyK7ThkzTWI65a4RvalFXpV
GfD9j2ZPBTg5cgeg2Pr9k9Yez2+lx+GIjdE4mrnrFsazL9quvpfCX4RzQzat
0fZS8AljZOuUdFRiAs9E6Azl1wZ030R1BcVXHgFUDyjQknuVo492dGJMvxMH
L80y+CBOG29WvESgal5K9MPucpUfjgasb8VV0fgHy00zbul2bIQouFNpdv50
ZfKWjYhf9SpFrC8UlOvxlF18ssUlXCVOPsofRdMExgKacThxb30pWy3Hl2Pd
ComaFcOsd3JJEZf4XGFSbdUJ4fufMgpDv+bJv+bffD1e9tbG9ObFdSroYD9e
0wh+8V4usmiudnEgeIt/Q81VdSqNMV1bw0r8aVa6KEGd0lBLyQrtKR59jYs7
r3ZE9XTEXvFIpU0nV6CxBzjRiarNSlSRzpMV70OVnZSxSv7CPp29Qkf0QD4N
NunW2dwN9kOL/X3kB4M7tJBuHoTLgRHDhHFntJEb3IdLgni+3YyC5aqKXF1a
q+mrvNR1AWGQPrXvzSZtT8Z/Em8WelnxoohCLzpbHcAwmjBK7JawZcTv6zvW
gbtQ43PVawIVHdraY0H2H55Zo8sy0Ar5xEKRByrj4vjpmCMYNZdGAD9Fp2ex
XvKtc3DIxlOjLtaqQmvJvZncA3XH4Z3eJE5gKlY/z/nH7w3ZGXBv4DY1uyaL
or2noAh9XpvQnkhSJBYJOWzkxTHdF5xK/qIPqBWYGEnUtSJV8uPmeHDX/OU6
uVcBANIBJGjG5jUuHMK7KSxjD+zONd2ArR0ce6T6Qun3zpod3pKbWUrqxuAf
04kDw9nO6kQFLDLZ7PkXbzgzg3bh5x7BwBqK+vvp0XdY+ozTQCIjJe3eQpbg
qqrFV62UZSs8IDMgHVkT0xq/dpihHPaBjhu7Vuy0eKI6NlW7FhdUxMlDIQGs
H95zBl56MCXGnOmXFa46AWpHxZc2pq8bKJXmC3X4PSkkYuh+QIXWlBXh8HSz
WDEQEC08iJVZ4JwKdapZggbhEu8j0/TqWf7MN+4k1LWfkMnVtAsm3Gku/+KF
tfpROvvY0VEq6r6e3ndsbVqVFXTmShJXI9twS/GcQTJF75k2y/q2P8p1XqiZ
G9oAxIpBJ1wQSPRXdfw81UOaga/v8QBXjg6iBh5KwfJC6BeNHuji1qXkYRkT
gMx1IK7kLOs0AQiJzP1GTD3VhI5CWMzXJI5JUbqEJvMRUDK8lhpeIOWDk6Un
3EKBKy16QSu7V9BbQaHOOVRgDWVu8iwxGuEcbAUlcFElaN40LtG94ahBfwVg
3nW9+et2o2J5G1YJLt+2jtIVWIBt1ivH1EZHRIjQQGwwoB1asK8TB+M7GuzN
HlzNkAMx0jhzn744XeArXAWd3v6ZEfSMWMC+1jfH+sCFkgqm5hPLgDcZvOya
mFvMyTc+qpi8xIQ82VlqIC8KLknCzz+qkLJEk/SUjVQaoelKDP9UGRwF7I71
JRnfK0df/j42aGES6UgEaVWgy2f+29X/3Y2z8mIfdv+i3J9s6RdezAU5zvA7
oqSi2ctYRKh+Sz/E1ct2d9uyf3xgSebO7hSNgUuLRRv6EkPHUTLq4xrFkqfy
bvosjfrUb7DZl3IilPUUm//FGK1qUkqVi/E8mz4NyJkB6UQj20XhCgNSCxuK
S5HmC8a7vTqzKUOyf0ZScwrmBXfgxFNFiXBAXDzsyl32W3vR21VzL7LBLlx6
uN6q0FmO7YoA5bbo5buE0U0KXvgK4Q2NVcvOTwOejygy7ijHY3s/3Q4BXcZW
xECkvCFk74OE1+JhEZcrJG+mqQdAHTbqUB7GpdO3xH+mt0606Q8mRBqu1jem
Fcs6E3W80++PHAIWTUbGzZPZp3jJhiQCZq7aOv8TcO9Ca1BfCv74xeVHPyOa
hZY2hctOigCOz8+8UT/yfmbbTYQryvOhiIvOwG9LKiRJ9CAUoU2xup62ux2V
MTYHzzXlKJ1LiiSbV007zhQ0DWWOWN+wjMKjKjB7xT8kStRhzmY384IVfzlo
FoaCx+Jovuy3O9MN5jd/H6lg/rcpFZRzVMGoHIsjWMR0MnBxc64AmkZNLRVQ
csx0Tm1rza+sS19/f4X+TaTUE/htpOFINfwEnLkAGncJsHLCleLjkwX1HRLw
4tlmsvK09aO9ICvK9tGRf8mtvEXp25udP4r05vp+N/tnDBEH9IfdWEeGHLoy
N9Kh5DpYN7LNgrf0dGrQMYaymMqDJAb7mXcf9EmkfMF1coEYkYAwqwzbEsEI
NhmIqX1S3fm9MdUbzLSR/0QpfWr6WwnlL+4JzJ8LPVw5Nz4CNflkYfeA9nAr
0PcCKiBordFB/K8KHeFI/SxhnMO2fm7q1HJRDLBKybBHV+Afh9EQNV//r1b0
rbY3Ng/qVN0hFt4TP+2b4SK0ojx4qaUfu2bB5SxrH831ItxRyvVj34j3oodi
5gi7QXu2eCgGqC++cdNJZl91ZmIVaXsOmSdZfjat9OdD8dufdMDsuT9AKTbd
8/sD7R/vt9iT/wiAAizpvNjdwgd67Og6YZYz5mOwCvH69G4rsXlsrWzanXcn
kRspHQDy+73sVoCLjzhjLaq3J9h9a/wTk75FyGA7Vky/sgK33voyNKS5L/oY
CU/CaEoe/bdffP/7XwaHQVgIodS+e782lL/NNFakeTmj8ZseCuX+HaSViJlL
RgeOCJAvtIIicL9aKCkv/R7F7/sSDqX/yJi+l0MjBMbGrOdZyAwntesFXIkM
o6RCmz3PBotcsDDL3OFObrk0YZHmlQIOyH89/hZyQOhohdHdtnTUKXs3gpIb
rUD4QN9L3yNkz8Q6tPAif76j13ZT1IXJXLHzXlpp8Kb4hiuq/sKzbkUKQPf8
EXEBdOL2pLDjNvagiXQ5qsRpyuUP97mfMs0hRTcR/sr5L+d6IajfcmzzMhBa
shfQJgywqcp3SXDERNHHoy7mXzKZtccVw7BStKonsB9giesMI+N6u2t0JiU+
KqRdn2QXBMLc4tHS/ahBkhBeqU7stSgzOFo03ceaUUQaLXTuOyIqP4foe9Pd
KfhW1c6NO0BHzWvJ7xl0o2NIhhhocERd1XL8w/tqXV00klbgibGS+GLTySvh
VUvKaEY3sOORoyi3dP1URtbRuA655apZQRtP00I0Ot3wGiHKYI4pI+g3NFwf
qFr+PgTNXLtSb3OHoG/G1clbTbDrprRF3fC/nuVGPWm+OsZtUl2qad8eGVFX
cg+or4Kv+MfG0hIMFlyq+EC3Xo/Rmth0fOF2I5wcPQbddd6AsM8hqR9CUspi
85Bgde/k0CGDdhoNDd1d9nZkJ5F7B2ao6Be61MrJcf+IL2RlLkecWYIPL2r/
QSCXRYwN2XsQl1uoRjylSF7ukQh68wA4hXebC2FFieFLQBMlc70lUE0H2Qdu
LdtMIqCAp8oPLrL2rWB00DH5KSWSHBOHqEtVn6FRVzMEO9PaFE3YbAOUWM0F
Xm0gODcbsz2SNaK2qyg1RPYBpbjpjOwy3b42+hx8kQE+2x24oITW1+GHpcHN
xvA6IoWflhXBoQziS1Pwp37DzofV1gtdsjbzvpKCyEGa8v1DSUnK/OgPo+vR
6VaqowKeGyvhRv9qUci2ul1mP67JwAEk7rTfDfno2/I8HWxIYH1BOGg/TIlF
a0DzTmYcwec64hB1jqmb99woqtb+kyWzqWlx3wNh1nmnJFg+R7Zrr65Xux6G
8L+WvfZcHGs+jtVVpcblVwY1ntL34dRtpyMOmCreQEZ0EQ94MtwNWMP5siGE
Xz630eIdeusvcuwPVkYuexQkNsmuBPa0+ndfyFAFz8SYNn2pKRkxJGYYeDGk
zRSzjIzVMPK0lmuUOdvXR9TGF03hRpGS50D6T8RFIaf4oNGex7YKUMGK8v7v
LOWajUi1Y8U0xTVTGNiL4ETkSHSVkVlTK5CI/mpPq5eMOpPC20W88aXDmlxL
x0v3UcODAK5kV4V8fEJTKnJPPZSZVXKwgPTpdz50gD5BHUliU2UGVtHDhoyH
Rdk/2gKrd+qeQYt9jBGvPj8Tu6w1kdfQvwk1/TAeoYN84jgKM3LAEShq9Dmh
eC7L24QRkNK3+8OJrGrTsiVjsrLq2kvDBNijFHxFMy3pE/Ya91qG9Nv2pa4m
TXDzmdSpCGvW8VKJ/VTdYNs1sUHEVHBsEMMx1qQW4x3I0pzhXHP5O6JFkpdF
TsaxnweRmyVzPSyv2SGdFfTWda5SYMpELAGwmrVZwIQU1X/ZROp99BdtkE0q
bVzuIoAzErswMP+ItTZmXL6X2IQG8kWuNTm7Xn6rCrRA0RINwk6zfzhjSxXR
3oXZhXOYspTTSF4y8Lsx42zqXNAmPiIKDMmX7Cr8rMQChIDbgbzAN3SSkPIS
nisdMN2J1ua+CLE0iuW6tvhgsBfwAhW6ZMGU0dzlaL/04EW1YkVYPXIdxdAK
RdSwUqoeXFnyy6ROO+A1D8sEhnzivY4VpdaPAlCJvjZx+53PesfwLS+n4tku
4pRPAyEILwb7dSSlRVXOe3ReIGfadEqQbLOBb+EGdOW/IZ0W4DwLsbFNonkv
9tbC9AbRuueLmwQlcIXuPvNfSHOJJIVS5S/0Oib3KH8WTBZ73fCzYPro+H/l
h5I260vJVQox178LU6hqEVYThAffSbKIii1chhyWDBiXg1krdRnyB2/ydotF
BVeHezjY3Dpc/1NsI4LbgzOIP1Q3K3vcCYYjrjFuna5uBHo6Oc9OHIZa8XVr
Wx5y+MeTJ/oiG1dQrg9LYI42iW/cGPhi6z7SFuVtpyeMnV2J2agKAyohBBUv
v4KGHVY1LQEpyPY8sREDEoqPsdaePM2pY558Lr2YGAuOXnZcCVuF+YQ/jX9E
rtzyg9MnC38r4Z+eO8c0owLXo5LlvRYa8yCbIWSjvxXRQj1/9vLeSC37ZxBT
HqIeMAQF2OJYd7fBB+nvRoou8Y2MVjVACniXEXjygFWb7wlWiKuZhnDGt/Sg
AqDw4/mhg80PmIrXyBQT+0TsCM/VcaDzP8kLSpwn6wKrBeWYG+lvME2JEi2T
zuZaX7jIZeXGpuNv+hpKT/TiRCgOzg1L0nUzST3edkQpGnl8t5x6BTjYq1lp
QKI7HuiGVqbV7EfqvcZCoBjkgtku1bg9bZx0nb5edurVXeYEdZn+y6+A2fWV
agFgHE2j/T6aVBFuPgtDG9qoSAalnUumXQw1U0mMRvI4vuGFD2OUTVdW2JWw
4Gp5KNhY/oVRIhSdPgt5Xxb4rdTNZKq98oB8fjEAgnAd+tkRQfGv/o/D5sKM
IrjA3UaAd2WiHr8u8f0Nhs6/wKQG53KP35/W5KJoHcxFQNFMiD/6/0fbzbT/
7YYluuuzz+Nt97wC/p66oynFqLnrPLti/VcSoFzNs79QURx2xHPbICkAD0X5
KgMY9VIwZ2M9Whg9bAelFFTWJpCbEXaAJPRO+BDq369PYBxfgox9fVlWThEC
xZoT1K7hraa9P4mUvALyKFtEeWdlJYNL9GwpKLVadDXXaY7JpBPtgrcU3kG4
V0KuucekOt20cH1LaHVQuvC/b3Ur1eeWgR3jXOCGKlaTDx/RwxRt1OCY4TIS
gKyZngv3kd03B4losRCG8AIR6YcgJC1quaNTVgevrXLS8m8Yl5BP2leFHFCt
vvAHE5O0bxBmnTWc8cpBPfgJwhHvUrtYqN157o0CBy9iX2T803He7Oo82/TM
3huaUHHOHfxaRLW0PQLOZbZ5gVsVYD19Z18eIg22yJGyvJ24WwbJOKGL7PxD
oVDE6GaQfF0Fz904wTv0C4ziknb6H3R8WxrAh/81C4gp9LvmgQBYclkdT55Y
JcMEbzgsW4xxZnY5Qvmpadqx4m5dYV5QKiHcdIY8KuWYrSMklFO5m3d/b9Ng
epZJAwY9A173YPIY8S7+KExcSTmRj0VTjIiDeqOWiOieRjWnO98fiPcB4mce
LB7OSCZsvl9CUvE6WDOspIWBMCMnpuwc3yQ4au8dIePqlUliv1/+5Bod65LY
Zkyf7KUfDWhusfzwmyuFyOOe3xuwJGEE6dpoT1GnaMIziDL91TCt6cbSXN1v
jy/c5UpW2QHtHAk9+EQPpnCefAyF9Ao2402jZRMp8NkLop937af/pYgktYFR
QsDODDn29Fey1FyEcZJy+UJVR/juKQgFwKsRutxPRDhsUf+ZfjKOCzCQDLaz
9FNeWguI7gc8dcONXzBl6KpbwELTZc4r9VYVaAWJnmROATIlM+orIxD9+j+D
nBtBOz5J8AwCj+uwiLVpl5DH6y9Av8lyRojnmKeWgQBajdjCwjJIgnMjV49v
b8mlNVRr6s26KUYVa3ziXjRC1jhoD3HJlcTZZVdNjlrUxZmKYG/figqirIWB
BuNENPnputTjzO/4D53RKJUtkv9q//AaymART1Ro9qM+dIyHS3BfAfZ9VuIH
dsbsHXfkr0WBzcmUMy7XLZ0O3UEdubaLqAMq0HXqhHsg29dNSYsRcSPFFokC
2C9atjuK//Fi5WijceIpYo83eTM2DZBUonNEOPDayQF6u1LyJ+lnXYThiYX5
ZBU6b1dieT9Ny7YwQ1vBxmpC5mljqYxllq58bRXYW7v+4X+iazDS3mRCx9Ex
L3s6ae0IOBacp5zp8kWF4CeFBNdnnNW5iJoo+sSdEtXehdCrOKQWsq7MHYwX
45JJvbUgpYlT6nXbF3O8nvAwT5QiSarfDcUCE5VW0pV7XSjo2XlV38Iz9Bty
xOZCDPd8c+0X15q3HXXU6rDZVsRuKdANPIfUF8Sma4bQMbdmgGrYxvTMO+X+
GKo3PAMKZYzBTkx/2kTrbQnEfNhIvp2xdJiaiN4TY/BLJGjtN9fPN6dzbsYE
uRexPaJqDZ/c+mtJripk83GLCIjDLopGO08tdLgypabZYVoSvF5+lIIDL3vR
e2GkNRNGp0lQgkH6yazyLDz3oWr3uRGTD5xAjTh+gmA0QLUHW77tG/ShoKtQ
xP8xYBlc6u1wNyrfYtyEQlwzIBdxHWpXzGGbQtuMgepyTB2Lm+xDGP4ed/an
2EuiSw86QcaiAO6dy8N1t/zghnNjbkjq6jz9W8kpuTcinIIF4FBTBgpL8Jb/
WX3nKjvkGv1JBHJMZqlhx5gDfAX4c/Om7G5+qfG8AihPITmYQuPbwIj6xfS8
xlScajnACPhKgATdG5XjENvVMDx8ah2dPHdIfoKmLdqCyZIG1rqDaf9NfbOx
qWjF+XRGsb/j+tIeqJOQBEB8cQXD3fWE5zSkGgqdir2WbbOnJuVY0a6iysiK
7TDEPpG7nI2f2Ttxn+p+qa/BBSO8I4qwhd7mMMzDJth5MIvg0m4DycQCQqXm
EFd7L4ywGcse+esxhVOWw++oy0m5NDPCZgPS+dYhH5bl4cY3+DSq1ubpMMub
kAWZDRhJXIEhCsXAShjcHkRhXT31bTOYvN1g2rj7e3TJ41qEdoAOIUwRzDyB
RaEFOc+FGr4Bq9TfrY+7mreFBvQoyzP5YAxdG6CWRCF2qE2BSOjeunDAa3oJ
iFjvAKZ/M3jbHnNZbxnEpE3EN8lsIpgS3W2RHqQRnWEvoO+tP8uz5PluO9jb
qK+nTLAaceDSOH8ujlJpmz4ZOYroWSksaFdOCX/OlFbI70qmOIpSUt+4kbZs
Gbwqu24Yk8l7CgDrPEj1R9gdN+q8LTlGfYTip7xL+ClLw+/GPvYhZaKjQSeX
XIlo0pQ0Z1jSq1chhXpSFR8SyqPOyLI0M1Z4qDpfYs4ckoFWaM9Bi1zSR6/w
MvI1yMhd9SShE0v+MIczM9Hva15tS1FSPzkPL+OtUsi9vC6P37JCR1PidXcY
7czNBDrjT6ra1VwAk/T3lGvfJEE46yOXLfsbn6dlzygnDoxSR3q5LKOA1VRe
L3TSnRBB11ZMX5U8ILXKI9QXJFerTymW/4l/7PC8HMtKAddBeejNchxYwTZy
17Q5nU7M93shxXdpl5Ij+aLkvV0TLPGEF7bVKJmz8b856WtaowAj7MVkSwQt
Qo9RhcGr4PkNzEKUU6/5GlsZK+kEooU6w0tUpHdJF76KlTn7nRK7dc0nyeR5
DkU/qcm1EWNoetHmVx+09o998fz81CsXj6dmxMc9crpQlQFgpqk+wyQaYmgD
bhhDrtlD91ND5v4ZPkQd+x0kcGIyv4BivbdqC8rtUMqXrixWvy0Jy/bHB4wt
EDTfat52pPymD8yO07T1Oe23D6ZadD1sSunsyD22qvj8e/MpM/J+a5k1ewKI
v6xIUtzHefbiunDlvn/vx7qKr0UdH5rfVSC/cKAwSfSDdmIOEowde7L12mIz
HHa2BMPfgdTaiI8y2SiQ8FYav5/2SY2PBXQ4mbFurBBlO/IZzzURVtlo6qZa
85ht3RzgbdNwA2wWbBFJ+WTtLjj/GGn2rlKwOR6Yb+bKaj12DdFqadJEpDTH
VFB071F4lrPiH7vedq7Ozi3khwPSiXuPI/6ISE4ZNlTrSysdEXtsvJEokX94
QqST6oAJoWrV5zCoZxU0a6O0nZ6rhAIUZNltGxlLYB69PuulMVf93kTV0O6s
8jZjPMNmevy8aNf5F9MGgU/sKGO395IPZsqAGvXPybA3wRs8zrgkA0QuRmdS
sXhCKN+pNDgJ/3dOV6Xi+C7DAmfX6+eLsq41huo23lF+pkYmXUx/iAoRJVFk
3h1lejuTVzwL0cRlUZRaQ/MlAEic3gqkm6/UOvBZHSg+9lkv8lljh8A+MHNt
WY0Caw63q99tv+Bm1f6MtZ2LXGjliPGzuVaXvxSKCMZeuFAveJF+icvIPEyR
pRVsiIGw2y8mNVevHSyjRL2H3fgBCGZG3PUqZhkJdtduBe4FN27FHrAns0xG
G6xsIak2SriWVuDnB9mfnoghZrHcT0kwzZCaC2EAwCDcOSYLLbHItCN8lX6E
W9ekLCxwDY7N16kmAWfT1Qmy+dcopY9IPJI1zgVzC2/tk4jETx5xa5Hk3ZNY
SjoIVGwpIMYbQlz1sDMPbOImvy+SsJs8fwybko5AqfVfe0AWxmUz+LZCkuPC
UWnZ6xRIwaUiknzi1JHcCcwjmDG/tXWhpOldHfjVDZOEnfoOjfyeZejVQKnw
t4rsySdYVg2cYCQg8dEeFZ11gN0/3JLUmmyzxjBXaIM0qjn+zjyog04qiTSc
VCIwc1wtTgyQZy4kVYqnyo0x/qUYK0T8UHjrqqLEvOBTB3H8Y0BrCunUelHf
XIIPFF+xjqSFys/h1r0MYOdI5O1voCzJfMhGb6hs3nGG97yF8iafFZzB9qgN
Wg4JIJYdx/LaYra3pvmcBSWa7do/WsqBiHrZ6GX51Fjuy+N7TZhH8JKT7GbI
LXo6wkN59CTwKW1SORawnQjDv1LagkTScj0rgKSzWHyktF9ZkZLZ0mriLTHI
yuR+SbGjpjS/mXbGjh2HkiVDtssI0JyB9onmVhO5fBHXGZ2T0TyDTYWJlWWx
OwGxptCOYuR6LPziA5WBSdu0axQcdeKWasNtvGy4+AgNuO6t8ymc6aq57RD/
hBwkaFAbbbNRViVjH5lxYlDsVtpAEVXKUYXXwtvQcAAR6utm+EUXmwtG0lal
a+ORQx2n55eJG3YHaVeF7WNqC5PO41Ww00pZiPlkAsTAEXj6hGGvbJyPbsC8
gb5SxMwoyDpfukrWMZ5w8BN2OBxAku0aS2U23BhZLFOsHPnY5UCiirQ6hW3S
6ivm5+Yx0LJrli2pV0fR7SvvArCB6d1qPgOzTbSBBxr5InGmwLOjvDT4Em57
Ylb6fvhxHSEaEYNmsvx2a5goBTr/+uOLlmG95NTg3oaP2IqiyjhFxAsW0NRb
p+gVp0b1IZDwB/zSh7mylG2spw7NKVqrP/iWIwMZzSxDzsf/AbDaPZMRhb6p
GO0a2p4eVbfpsyy2bHqkZdAl+fYotL2e/7NaSriI+YFHoozCcxYyJoNAlsbs
F+xmQhAhvdMIPzzMOuflqs40BnjNezAVERHspIY/3csESDMSy7GSAwQdVvdS
bil8PNizh3cUjiyExVcSX7W8VlMdLB/wwoRm/Xi3ONfQa8YxlmWI71orKT0v
hzfozOhlcU0jSua7fFa87bijK0nKbmzKI/I6s1y5Uj1rl/yHbPX+JHZigbov
+pVG25J90HIkGM/0CfvUBpqBNdKRDpSSJuRdrHMWBWOnkgENYKSvz6oiZrcA
DrwVsp3e71vUgZe3TbQuAUyAAEj79p0QNjWS9wY6D3RWtBWClTJbGKjumiOL
OMtw2o5KxWXEtngvqoOkBpi0E1It5JTRQlYYzeaQ5pd7WUUbBsOOKVp3EyPi
6RIk1Qv8zjHW7uhDg/dXusJeG5u4tzIm+YCZYTc+ZTP7sC9Bw1HUY4+1vZUs
Iv7raX2nLkvb+IU5r1uoyJmjKBIhbPV1sfNQyGIKY+aeLooQR6w4aBwFbvJo
8Ywf919cPCDfGZ9Zx5C+2NvbqxRMY8s6JQKoRz6uIFsQbcFL8/NNIgw48/U0
/36F7v4H99iqLuVwntw2j/AE+7PfymfNkiIjjDniDiwNaRsf4KyIqWPVRM0M
nPjtReRB9TO+GqX9xdqFTCtUYK60us9sIbjUZpGYMeVQmBrA+XYQut0zMCQ9
sGzppLF83ki+5oVWsmxt4uCi1GfzfmvnocV0Ehpwrb6uwOiBAd+anMvko9O4
0FzX1ynpoSSG42T8dpt+2D3hmxHu9kcrP/IUuGAoZxuK3RRSRxTeKIyWNCf7
QVjbdgOEhzEQhX2CLAl5QGhrJoXVDUCZmUv91Mr3oogsqPN76x8jizZKiAeC
0Rktrl8rHU+ZQ8Ho9Qgvd9QJaGSZFnvZ8SvGz3sAAKtWZugUE0VJSTZKlaGV
xSkgpGNyCXjXL8oL0MRzCVeffKkWf/wEtGm2eIYpbx5SsNHsDrxYsjxYRuhY
6rupJH9xR8VHp04TxleElABw9zKWn35jun0o2Jh6EdVeusCUyRqogF5Q7789
RcOPNkAQrY+zK2VSajlptylBsWkBeUwwfycCFs9/IjzCZQklCeRGJ31cwnQl
JD50yc3syFitALNc5uOfCksmCR2BzaP7LYk1E5F2OKBUBOQxl/1kX4F17epS
K6y8DIWd5iUx2fv1C8nNuWB1Rooq+Ba0TdrROhSnUBtna32VWxXyEonE2VH5
ct9OA1u/xzaM+iQ1SVM44EEnlFU+MWVPifnhsQbd8Ojnblmy2ioFTdaXE+fF
SiVpNAbNb10fSZfaS4C8I08lyg2HXS+U7tz20AFgI6o0ykACQ5ZxTBMXnmcz
tC0cI4Kezvhqe8TXYb6U7loXNoBrCokAtA6TOia55Nwe/y7jZNuZmn+3XTe8
ZFcWRrCJEPicU92muWURZji67K4TXCJa1PvpAv/MRZJxvkaA3OKTuY0GlVYb
TOBvvs1EjImIkMRkT1VkM2ksKxny9Gz76yXhjxrvGirpK1zJzSN2FK5xs9cD
K3CFi8NkidwBmbZceIusFA9Qx77L3E8Muuy4MRaIdY6U/hYhuf6wfCSsac8b
0Iazif8ObE+kxqZCxjArIBFiPhDv7Locba9H0DAqX3TsqLK31NFX19LkCCMQ
JaajP+G8819lqz7LsA5ZNc40bZitc8Iyn6mSjKmR1eGriBVaW3pWkn1Q5k3V
apHISx/F6Mzv5RX3eJKFupNd+aXH9l0wK2GoI4XAUjaZpPH9idf6zZQyon/i
RTtIiXcm8mL+IIWIrpl950tbxZTwd5jG/RVBH5dj6Avdv68wfFN+AwVoaeE1
WQ5/w0TGYGKBhlxuOWVTufFjYTho02gC2KI0x/gphXswfNLzeTB6Wod6kEXw
Sk0XUQhuR66XNEIXaAyxYGwYZgylauinTgg6ww9+uKoJRtK6ZMfmUYLWco9w
25AzPj3CEQuxuFknc1tGz/nOjJNZAWbLyM6GS9boFUFKtXQn+tjQxME3jHI8
gn2MCfvzm/tVkYhqAHpfV+5B47YmX05cPGfEeVNYrn0zFj7GWzzz6AIFd/TM
IrbXgvL7UQIdVTu+kNq/V2r0rZh0OMoRoqvipVXVqZXumNFpSJndu2aFgvID
eU7o9THc25p1j1k9T6XceZhlbOq7sXINw3RBjI7szqwoUiF3ot8S+dyzax+y
Ltw/eM9pU9aOzdqhCGs25/0k2YriwV/jntEwSL5A6fSzsOLCg+A7c+fyVAo8
wRUWM4RsOGXyfSsndVtx8h7TYHkq2+1E+jBkEmOpRzRgNMAKAH+qZUPCtWCN
tgAJxUZtQxmV4tLigRLD/XNpc732C6THfUh3UYsccVpbasKCqmx81Ol0TcB5
m86CBE2oSaTJua7GZwqDwTcaJDMLF4/DP7noBIed5k8LWO/aoZbUn7GHq8Hn
HSkEn4kjuDQt9pKzVOoMoHuPJWekculcEdirZbbnuSXtjKnHLDKpnVJDlYVv
w2812PmkY+yTbkCePTIgdAWtYVveC8BYscnHNe2rU4ZcQQuy+6IVdg8q6ICu
JD5dfOzehYYfcsQBtQ+snph1mJ3oisWsfKi1X2boKiWhawk8h8gTA2jOB8Qa
Zu9HJ0L8Apgh0jsuImfli3n+Vsof4qndqE4oUrwPrBFG76xRRngcpRXEl8Ju
H+S2CYTizPT/rabMgv0wCYAjSLqhXthpUW+AvHiGBPUPuhIeq1zaQZrp9Mtn
xX7ePcYjtUPnFiCngck9NH3UUILpQ9EAVOAlyUuvY0padOQvTcXH5/cHx0ol
+u13PcgpaSy3XAMTr/88EkcuYcYTtTFmFvaYuOV20QzJEmybXW6FkuV7xlQk
CT6YhKG32UFbFFqdpo0S7wAxwYcdoPW9X3IFhlyRjJShvJM26r6u0788wNHs
9GjoC/DqFQDA/tWMYLmcxyqBhdF1Tu1VqofXWpuv3rg8cW6qhrG86RimD07p
NpDLKYmwH7x604SSs+HQZ3TtLR7KrioGAZ2ztL4J3UrRVu6TflpNZu9RUHwY
HwCwz9TU1oAQI0khaxBsxn50fh2LZGppJ2mxHRDCQJ7oSdoUeCBVpcIetXoS
PV8thViOS9u0PX6EogE8QYDoZ5sP17p0YfX+Ii16sWArX26g4GsbPJn8PNgS
CO6JpN55du71gDLUarr0ODZW+BUtWdAf2BPG34LxKMYCttuXnFCYhIhciMNZ
tQH8s6ClAmTlCXP053ujyTQ8pe/Oo0yrGYaxeBYLVR6Ur/LbJY9WcWSJGd5x
qssnvWIFdh23CK45Wrqy/yNl4GwYA+3CLiVEgYR5EKp+IeHwuiwmTaz64DKk
nDG4Z1AvI5MulqyCrRLaxIv5Ysl8l5loSAnhtVoIMB9oH8TkdZEw5UsWjGxx
1fM2mIvcNCNRnoKgE8Seb9lBvbsgl87MRjsx2bMr5tNMPw2/LMN80yvA63r2
+VBsHyDtK3jJwhVVA2Rz0JizojDS4hF9Lg52/sKMfaeNrRViSmzHyTJAMQlr
OAkfA79dcv6yyeA+1bhyxFxBTEzDLd8RYH3MgBE2aWXRSXVlUuY4WtTvoLXk
iLX3+UrDx7Ou+93em2l92nwAhKLsiv+R/uVoG9rm1GBCggwZ5+miA+YjVuCF
zoFhmeGk/oqg8pyi1gkAIQ9vW4zPK3BYEnQg+BVYTmwUvjCEsflEo3cRHmN2
UG3pdSzBNtbE5P1iAEC1M1z6ofR66SwD6E7J58kZp9Id7ugeWgQ/NLwgq4FW
+3uSIphcEru5/E+KKkqu+/CprlsQd/0cJkudxC0OCWf582YkhL8uMkvp1Fy/
hN642FjsB9sZfpMJoaxoTjkJoVYvnRTzBO8c6I6hdSSA7YjxH0h2ByOuPy1J
TAdPurU6fHnb+F7q40+jLrznWS9W25HYBndvSh/YSvxy6xNCU6ROjo5p3V20
lcP5HZ3epbF0XPRtKNfen1tK4QcHP1UvVNBhabyHNV3OSc9zydiaQsafTJLG
B7mzH8TnmN9OX60xkMGQMxL5dZJL5ji5gL1iU/7BGwye6m471ZwG9aF8GlcW
2oxP2Mo1WUJvvS0Y23FCvXG256+sVppoe3sNt+UuwGHJ6p0yaOcRTzlk5ocS
ws3UpQHJ3EbpeJcsf6WL2/qJHt0IbF7o0XDbJ2IMLARkTXJ1DyV0MEFeiV7F
imCuihyuuIHExfe7ITFeswqzcXhgflt9NLPs0x6kYucBLHbZW2ksQPO/1zCo
5/f/szCxpgoj4FleAJmOIgmMi8+65KsfRxs/WyS9en9CM+pFL6lYlHIQuhHn
lKmWE9yAO+xdMOqpIcAK6X8JgWlRorsFOJVZ3Wzd30VfWXs2Uh0/ujiLIQQ0
IDi8YGq05UzO647hhuq0OX4JNfOO30auODI/n8GKeH2nZWI9NP3Zlri+oU6i
PCd8IZOL0v1uI4g6zwCcWH9e7j1YOfdC/1vtL3p2ZlbNf5q47PQpaw7ZdWgA
t8H63Jk3hZlBoD0w/QWslNZzonAK4RszpDlR0Zt6ninM7IWroEpBhNA+TiC8
VhF7kqwThVWeONB14jqjXe1/hOy2uBHKJ6NXZHzhQ8dBKxOrPVOwoshGDHcc
OLOZedLTx6w5Qr5teWnFd7gPl3JQV/6rDFJjB/aquVICz9susp8/EtTZvEog
qPZCsi8qjJ7tRmQlGGQLGVVvPL/yP866lth8vQIUIWo9DOfkGDac/IeClAFD
xcmwbKfPFFsv7JMDlnj9u+kCRMli4axdkrpfgm/APnA+f+j3f7WofJn9zfpm
MyU85y5Y+lwz7/Ozia7i2yurd62R1W3KQ2JZn5quOBy4UuVvzoC4yMnxqRAr
CkONsObRhSWPf/eYgiuoBemQ3un/Xr5XFm3pY1MdxEiDnXIb/wRQF0SHaf4b
Kl4gfsi7RpTBJhau1vNuO7/tg/QSXEG6kCaUpWg/Jzj3RD6PFwiKObmHZlCG
B48jBKPNBkPFbbt6+93xds0Tv/0kJBjoKOpI7If9mhL+wMrK2vwuXdo/KwuD
A8jCxjpWcJumSh5uHHNEh6lpRrmjEDmhdvQQqVjY8fVHe48IJlPoizOiLRcS
GbgbJMm5M4TTdr3+q7A7hbqUMmLVXSjbPYxQ6cI5P/l3UFzgD5TW7V2Bw6nv
CNFclfkYlZAQxXWqqQps4x+hen//2y/DZGolnbQFEVIYTO65EwCzYXTKCmbz
izIxMK61JBEPrFEz4iiv/ewgUefqKDGHyGoRNY4LqAEMxC2Wv42NeJqB42ia
Vpvgafxkkpzs+hQhD6juzCGCeHBdQ26AdSMPdBCdhUBHvaW8MjuwQblGARQn
Q/yf3S9KxGlq5WNYl3L0VCC0Tifq3fYboe17MzRNgBMFqA4tzHs/q6IGIgqp
cssp7okk9oCqQkCc8lIHeHlYjgUQtc+R9+i6KqZV2+NcRW5UGI9NveGSXZmA
fOYYPiI7vO+Gr2Sr8dntvqzVCDwh7+hmg7ljw8tikihSs+5z/OnQ9Q0FQhJ7
q/JN6v4jpU9s3AuzFYHe4YWZjQQ+j8RWILhZdC98qYEID9c1qp0PBApntILO
6t+67vnR5rFFrJfj90isudt/OkYEzC7oHg4EqSls9/77Unt94wWA7dCii17x
sF+HgFo6taacUIPeNtIR/vGuv2OVO+alHML9bbH8ZLZPaGKiBacwsp2Awyt8
asBWZj1VLLe5L3Bp79UQOPdoDh+4yHIl1BFVt4gJ8FVP4W5rhVBjVl/eO14q
LdZKTtBPJK+V8vqulitByxAFtwdbshgP5wVw9GiV/3E2Bc1rjTDOT/0nu1CU
ZYcsomUbKvZyZriBbnZvmDV9B/9+1JT/3Ygw1WrFl77AWBjbdZ1oZzGHDEKA
UybhL9nYlHOesUZE2DcE8/aE+wunBmLNl3VqJCB4Nv+T/AmGXiXPnbO6+dyz
797ZBXx5G/rSTnZmsXvZ7722CYXknYB8ZNR8/9jXvOfDY4TigZhap8zphBy8
QgvTJxZe+q7hfGkfW1srCCyGmitmv8j8VkH8/DL8PgjAjDCBJrXRFZvdGA61
Q+6E5kCqvLcwUFGc6gWb/bmPpSV6bRp25BSg6mMt6e3a55C0W4XeItTD2B/G
loPNjYi9iUfBpuJkeGm9g7+/WZ2fNvsp5alr/JHNTJZwCZ+B/6VEjoZ0gO8Q
tmhT/wHiRnnhJJpXgvrnyTMwZTy/uDdzmTebWtPUGK9tUTmHaOX4oZA/nVZv
F9bHlodBhS28M/hS12yLnBHM3/NWcOf3DeEGI1xxgaPH17ykH8I8yW2Kvr/d
FAqu+f8kQL+sAxcT65wh3KcG4SUcV3EkKz++iM/DsZBsJxVjPxmW5xgLjQ1K
z/1fRIOiFKiqfIjLsA9OobTa3jJ+oKBxwbJAkVX/ry2c4v3Le6ex5xbXDjcR
oaw7HUkxinGPYGEtf2n1Cxu4JmrLt7uQbT5QtDaquHboAUUD5LmT9FBQPdkm
iMaC8F3ykAQoLp/CbrlM3ADrB+PLRpN9puf9mfSFDGVk/s+GJi3sebzTyjr8
3i9Z+0+q/nWD7ZIXp7q9wG5bSHfsfRHpA+7RF73Za1FmAoUwiaua0+Uam6Xt
fCwe52dYTustTIBIhPzeN0+sWx9WwV6nCmPkFAwGU75RIj0qIdFyw8gxs0Mt
gKhA2bTdNhHFCJtX11vSJH3yAjkTtwzNsCYTW5KdWO5MMmIFqwMszXzz4Yvp
UFDzF2OIwAYI/fWvDa6VUC9rTWMDkY1nAameyeptTSTtq1a1VqiHrkIUEb/9
I3pNaIer2H6iBL3QsVidDL9/5v4cpyQokA6gk878SsNN0/v7nGIPagy3tDGH
S5wQK+ZgNpb5Mamw1HB4MB7FcjH2inrCHPsNbaWIicJ+qECJO/qj6TNR2m9E
wzlJGhpe5FhoEmS6PvOC3NKYs1Tf4cLb+1Na3+5bMYReK0OVGW4pmdZ/Isjr
82cQa1SBZr1MomaTY1tKihi4XhNzmx2PnIyFLWGc4XFtPFvKpdbvrZJHYPC8
yQYoZ3dOjGv9vSyXWFzCl9QjC6LNqTTXdBX3loV4OR6vJDSyKfZVtExTIJwB
fO0CZat4hqhfaW4DbtJVcCue97BlniNTaxqIkULteAcNfrAP9PZf2mPtZCLq
C7ujWvBFQ++0/GEpd+z3mZY7coCLBREq1uIjLMjcebr5+W1wDFLMUR+quRj+
m4CvXa2B0b/P9CR4hCtO2AX/5swVwLLatPSbfzCRgs8TPebuI4gepIYYzQWo
iDTR311SZcbsNDVQiPohN/KCpHBxmLRUcLc3+EzJxvtb7g2xDtuxHOwnez4N
fGJD9YAp3Gp9Ls2kFABTQkJ9hmYwlqEX1DomCCZGp8xMSnVTTJ/nqI6B5qO5
Gyur1iafGPzr7jcNz0JGWZA8AxcxbMRD6huiWKxYEwfvSLEHC9UTP7FfpoR4
5ca5bec2wgQHfXlfCZsfAJHDZLWkW2sud5bDCgMpKSqhR0pltPbstd22T4nu
OQXpPNeU8FUtDxpwE8qIUehTu2zaY6vWGCYa4SHOF/3GhWconodzMd4wVLef
y57o5bBzTsPiiuqCBpND6XtC914BT02dQJn9ffrRxWp3t4YfqvFhV6o+iRJV
z/GNlubFGhmaTHA5LvrOlHd4vMjgP2/Cz65FuasVrr+kNzep+uLjQV93Ue/s
3FmHcWuZ8KHoes35vdpZytO61nElc7brObXbshIO6Ml9sCbjV9jRrI5i2tc3
y+g1gofHl5tEzn6zo/m3CbVgBgmKClKRGTvuD226XdHvJclxlqi1aEIxyyAH
zC2xtEd7WbDEUFvHkntsn+jekxlE/17e4Unspt/foqhbJ1eAQpkQ76DfV75f
PgKG3VK2aYZlIFIb66LXmo0hE17Fcdf2oQog89T3yCQKLm6nX484rlbxo2t1
d7HBtMr5zxKbrHkG89tUxow8HnVq9mrl7Ixq3dpEe5OUzOdK16gWPGtj2kIf
LlcE+qoaICEeoQRYpFa5bwiIaSCqFGXd4M1XPVLAfRLWz1iVkjkVBC6PZs7C
NfnGyWn/eYgFIHv5Dqb0BMvSSnnTvf6NWTdTsd1VxvnRoI/R9fN6t2QXA97H
dgKQWDQlnX369ePHLZaV4i3Wg1rK4Pxjdh8u1PHb4MRwNQKWKUy+r9cQ6WPj
ETsA+Nh0izHPtBDE6lX3r6PCmbP5nGb9AV8Z4WoJzI0gzoK1uuaeQcx8nTtm
8hapdeHrXcpmWq/1UrfSUHWs2r6wqbmlXsVmU4zzxgLUR1/UPpGeSEw5SDZz
s89i5W+Cg8pAMBhfclhrKUfaBoeIzGYrL+y4Q0P1YgJWCnDoqpkkDuqsHFhR
BqQe/3hLFoq/gV442pqU/fCaqfEHWSQ3BEnR7i9ksin32kYpmRJb69MFohNn
O+ExJrPu0ZZ4+mKRo8yuVNNwroxioddFFauE9F4LUSwx4tRHGyjoT3NImMFR
k9/kKCjhIjJ74HW4VEVLRvTkkfXYej+T4XBiWPusiRPoORZxgjWzu5Fc085N
8GWqNcBOva8o/iowvmSM2Ah+qYFR17N7WEp5zb5N5khyHagdiaYgXUZsB2cv
d6mxLC3VmjpjsVrbzu9JiF2CEdkJ0jQfOkcKEQ13tMcDR35cFLOCOLF/tEQR
k8+CO18GVPgflCEf3pA5FbUEPCmnMy46lG+iUo0xG2toFtQuEMMLrCL1jQmO
nqBBR3LdxReiV+FYT623BckPnvcEGypI0BwOtTdff4vDMhmrbGFZ2BHfSHwb
ss0csPVzX42x6XFFAX351/MLduNvNcW/wjeO9U+PPCN7XR5GsQr1UsSzsLEI
rttQMZByAO+PVREAARDBbWn+Ocy7dH3QcbbjwFa0afGdXE7KXaQsiSm9Jayw
leBw1XePge0k2HKLir1hlT8c8WdxtLD9G8I04jzYZepY4Wf2uClnQygyLtyP
XdiESyOiRcPwZqLAMYKtJp5F6VUvvXiLN1KJ4g72P5R3xOlJe0fDbNRzagov
EYLF9nFsyJhht4zy50PSSya5PM0cg4XRVL5MMslCOwMzLVNg2SrVH7pGsevd
u7eihJ9SVL76J/FjT51JBw+6yYg99eLopZP354rH8Q/LcAYslQMFDeR16wPX
IvQOV0tx+QnZqgEhUOdW8AOYB51fzLbqvS/w8kdRwGvomZQPbb+LBi58AiTg
MAgs6utSLf6fMetuOX9dA/scBKMK6dya3B4AJw0uPL361+THkugsjhD8QOn0
VwgK8cMsCcDHfJ9QqqKdM+SZzayOcah2kqJrTvlerZIxFlzasxu+ikt9fuXD
JLfy1qp/KHqda7wX+uPT2fKPBFEFU2oBXIOlg2Zf9QZ+s6X4dpjmcS68kgpy
AmNtOgKCpIlf2Ko1xqUAFWZqSHYQD14+N3PoqeKijjZGLG+6umECA021COlc
Awt4h/3oFeoqY/BUDNJPOxVQsaDT681ogl3X4qP+kBuLx1AF669Gck1s10mD
fsZr4SNDhMICkv/7AC1nLP8uW7FNyb2poRRsC48EzR7qYQaBQLt7xKeW2DVe
CLQ8TyxpOQvpBXKm3Yv4Cs1fDr3TQK5WBCQakwNbfUm4VFcsb8jMpSoJBbt7
3DVxW9hLStLVNlzBRG9DfCMVaCZNXUJJWkMxaH6JV58QUHSBYJMHdWOnOKNc
ZxmxjM8+NgoQrpF5yjnPtG5aKahKOCDDpQeQ7YpRUPJteBxDUx7rl45EHGlu
0Usahls/8EGD2QBKDkWBf1Jf3Ly/rs1mY+3yWLKF+BFm7FWGAAOTyp8BDrf+
fcnsFu0iiFzPxGbWBwoOiLucxdODFkE1sJx7Rp9C2q9ERGsX5OemajIvtCqf
sdkzOY3UYSnIKTnKJZbLHR3Cg67XOQOev6H0bBohA8oj9HehdQWfT/VuluN5
7/p6gA4mBLDuPyuZJdiogRidfocG37sU33qiFc2ncfRdjR1T2TWCYF3d74b0
Mw3jhfFqzPJcHsJSEuJrohlLs5TQjQXEw+mqmBvycREAA2RLna17488+Sv3V
F57k8S5pd78kncm2rq9k0ksauwt5ULrzenYpV2QmbImSg14S3wqduy0cHaCk
rPbU3mS7nhKCxPQBSMBKXcWckgm2dBIiYTp6GNFjfZv4g6MktNdUCQlpEJ0w
atop5jkLCfEA2QaBvFOkCwh6Emb2kVQnN1Cfuhbx8QhkuZmb8zYSlSXkrkkU
ZryGhaiTsSi26wFbr9LdLhFP7ohAdOqYuW+ZBpVS+eDXg158XUOb8MwJOro0
jN3a6sagZNdGD/U/DfVfCtGKf33h/t7GloIjKwOU+N5SLGFvum3n0DdwbYD7
jsIo8Pa1efi5ZsWEkPI5UF/L+8JnbWW1xIkixMlNLwjL97SAy3fpsjI/A6tN
Sesa/T25W1YCYm5akqTn2i5bNC074MpZ81FZZlVoU7hzaaq6p3Gxv4L5Mt93
upYMc/Ylh3n8DMkDMDoiXILrI5sC6hfuyME+13vP/+gdQd16Y5ohmlbDRPC1
RGejzSpSMRvjlhojgpVufdRPbacsc/jT0EnPTrzNeM39kJFRkxlMP5lK1fhq
QOeuiJ12v0L5Zibf1t/oGN3K34A0eEGKwh0NtfnGnI8g8kLDiMvvGUEEpwi8
fNBLDLcQ9QkjzrfBQQSaX9R3AzO2BZALgRy5RZnMIBZjdy29vBMRHc8bNJ2O
Isk/auF3YAWnzQDR7L8y0rWkPQKDIaeGAIGfQTbiKCy7HuPrIxvecJK8x/c6
Oio+dY7wpsdcqXg80ix/pRwUeawMH2UoTKY/qjUuswyk134so5hNpJcQdqis
CTBkhTcvl73GGopsQAxPfsE9+80s0pusKt/FXMgHpFsiKABX0GQbB4PXfIkh
P6+SfeiQXNgxEOBS7P924NjH1FEDC0cnghnHFDAx1koqAjb7mSxgNwvW1IE1
mUtVNcO1nVr1OTW+aSQSbMJyKloeLCngDIMwG0f5rMfIHXY8RdQV6+NAaIFi
V1b/uCOhjx6hfDNEnQ5CPY60xF8opHlNIEQnXQO5hDXdDypYXN1IUsOJP/oh
RZ5wPuKnSc1Wyrx+L2KWAdntH5TR5f1yiz476c37x2yvZwRdLpi69gbNFY5L
D3KHlXNyMjCsTNLNNMS17biBK5JhtfHeJatqHH+R5F/WhTGq0hn3I1i8ZIf5
W+mqTI6k9S3faNZHVqcc/Q+Xa4uNIewrSubzo4qZEyRHtAbjNXVWA3gYFN0w
awogFgclD9IorrXP+tIZOiGmki1oBcLwA2ZqLx59Rl2CSm2Rpu2M0gXpJH1Z
N4RjstEwDz/zxbt/+ICkOsUOJwvnP3C2wlWrTa9qDCEm+vWu7zv8nA7w9LYQ
8p4KFEJtWImgyKcmFxF1GjUKLhG1G/8w6VnwFJAsytxqflJC1m1/IIlVRiNT
0JVhLz9QjG4SUbKw0SBggh/+8UxbIViSwFYawlyl/LSH/yA6kaiND5KUG1uf
1jFQXJULWkfTJ6oNDa1fIfl1/IqsFOsATFKRBPforolFAAl1afPyUAM81Qvn
lexhSy0XDisQLOSkX6PpDYca3bsc9ESqMAfmyJnVX5pmnY+Vl89wa7iOwIlo
HCvKD8h7r0GRQpOL1emT0JiUyKnygiBtnZ7aaNsK7wl1DO18MqSzoOK7J9Vu
njY02nFny/8+i/DPZZoVK1phktFJPyyspEy9QaDhl9JDXK5AEf7T2psfBtAQ
7Ny1M9IxS+8WS6gZtCFDCQKTxTg7TtwJ8SzSyUVexoJNpFpeDVjc8iQSePLd
vGorr0Iqrgdce5vkwyrCvjmg+jWsenePNVyYQ+iGkhsZWAacHLTnz9ATEYlW
pyLKNBbq+UXNj158yVmjYy9pT6Ri9YYsp8VMa8sWB7ogvGduxV957d85fl6g
UKA1954JlW/Fi5wCXgGdapE6lJkBNUOm6U6LVk6tcpHlLrhAKgs06CN6c/5y
ha7YYx9wjDaTXUjvdVsdbwOVKW0YoKLqssdfWC8WOsOHF4WTo9sSoYkOtbB6
zuKyzpw4AzYdYYTBEIcDDA9R4yBTiEy0wBHb5taV1gleqs+RJha0zfc25Pzg
rOxIxZwWmhj0Z0Ishh9rwK8y4rd1HBPSvwvsuEPBbEea5HQaH6fO8zbTIdiI
Xp21AbZW35KFJLdwQr8V4kANuwM3HrDDIA39brcezF52THkrFQmTljpuLQPW
70WtGaZD8kPYaEVDvMfx3A9miNxynzPnc4agB+JESk+sVE94Jj2B9ky73IKC
LNg4za/j2f8A9yLK4QUq/w3FJFegareK24/MalY1Mc+79OGMZNX81mk/qCZI
pzGBMD8UEGwrsSQK7SE1Ml4HpD8GowxYkvxEy0qmlp1nMWQ+H0Jg0z5NsYZm
BysH2kNxCIs1a8VZuksboFLQZu4DQK5r6BsTR4XAHX8HU0coc8DOhEN5l7M5
ffbZMiaAbMWIE8wGopAipjn0IU8V/vRo+/AHTIjEoYmU2wtQ04DepxcnVLpO
yx3XtTai9F1MYdkAlpAXO3jwlqreLUViRdLrVHd/XMXZq4dOAIeYLv3Cdua/
mIy//yzBYtGNQZtVhfM9tXhsaBhyuHNdHuzQAE5oulJeTT3DdkJifROoccnY
xj2WaEEexayT1hQ5XjCC4xJcZ2RI3iCFqHbOQKRRN43BxVMQWEYzvgu7lcVi
mrm0axVYC48JHQRk0x6r8IFCctPGV1RZkPHOIA+i6Pcw05ezqplRBSvIl2nZ
rlUBdIFk32ENmchpPn98MiBkJm2TSS7AF/l3mJxVf2qUc4j0dsU1BLmB1r4F
aCRh5j6mVgWHp9L4UyvdlHLuolpaI3g9v7b2pTO5vhBu3gNG+XyuSxLPjQv3
4Y0hF3oCdOqbPsvAsYLwb+LPcvj9NdtlERK5HpPodV68+7FgLhVl65YFL2zN
c2tr1D1yzKjaQmsjeTX5P34GyeTJIB+xsTVpO9JDyD8l33hwLmGgsl17Vrv3
URzNnKGOopBVJJk8Ny2FWT9WoGvQGXmrHsdoQqhhEhEHmEDkkcEXjttZq4F7
maQ1faKYkE7wQyY3g36nd0sMrGzCxoaxc5I5kZagyqaghkPfRSU3M1SjkIsK
J2hrhHei1cRJYr67/IVpm7WwOwpRNEW4BrC6c+XNww01Yk3jNNBSh5JkMBL/
lbQge6covCvHRzjoiuSaK2F53bzG+7VfWYsoyp+7UJIMGb2NXER4Sdo4ObY1
yJR062dw2P9Kxi+Rjh3qq7hucLkjQESLIti+uq3KOJmWJG21q9kjOKzcAMp2
zeHXJMpP2tTtnD2PlA4n+7np32SjRPKHNaVold8Uytu7NNWYAJobJUgToSz1
WsAGT5gYGaWGetaiDR4JD9j9AfXVJ6ywV3xntm74CG7//nCKOUzxE0VdDcaM
yAJSqC96eYserKty2qGLumKVsrTa+K1BcvNT4cJAMSJqwXRNUshdgLPZzV+g
0mNoEAa/NTAqHvQdyPacvrV4UtmnE5x10kslLLd03do+5CRN27GqLIwlTMkY
kEyjrAGhQdfB3/jpjIaX//M5YbpCkQI5muznBYHR0wdQR7gPBupz/NQjnzuO
g2Ny4glJmW5q5OZFR16O4xAAO1fHIvSaMUxrpeqY+NLW7NbJzEuLt/hORGsN
gAHDlods8i7cw3/0GoKtjFeb+TXl77M6EbCk8RPkbz0t7gtUfx6beMN1wBsB
4a5nGHUROwRIqEsIYU/ykIIssmV1ZODMfLrlyV79i8ZI4LZ42NUOii0HzfHx
dOMSeVRFn6kebUO3DzAnGp5TqLrAqdqQaM/fwEaMQ5N7rV3AWXOJBXDw/cFu
mi4J3Sf9w2Gq8h3jnhDbUwav18+zXVzFFT0WwD2DLtDCAfUrNtSBnWUVuwzl
leJL7p5/R6vO2iRj9kNhTfMdtexuMuxAubJlt2PXgn7dNf8ypjN//UN5pFRB
C00qTTZulOHhzDWlSAhS4MUZZOI32my8ln6kZr5e8CSQBw6ILdtKo/unOoVf
GmmPOTc0zUx/UPl3v3nQVnms01vFbozoVF4f4UTs5RO2UxjuBv9nc7DJ34IH
avcZCxSWpHUnLh/0E021E7aCtnIcO+mNg9szhpOXHVyAc9pjr+LRkArSWLu5
n+uE5bfoKljZ56QKQm7IXeAKXD2QuoaRFrjvyHuYB8P0sUbQ28Soh+SGm1Zl
RP5NqZlvrmikqnUko25LkjXQAMbTxYl4OsVhN45bbNxFjnyUDmkG+oWJzYge
rABDMmurP2ybuN+FzGI3YMWghm3MtXhVFtLCEtQnYo5A5gh2h4bk8//GP6fD
escUWKx9Tlp1UkhqL447W/O0KpUFEaXmqHsi5/V6+77V36rq+cyYDWSYda/l
s5g4MED6k/MrDzpTqpwADcePefktB0F6qvV5YjB8dT66302yZHDTgHQ7dqVI
XCpdApO69MXVN8Zffde5s0Utt79oaTsyTDySGyFkfkQxS0APMj4sS3tJmDF6
+6NzAuYHyApgLEvKBQHj/v2A2LRAL96aKg21fP1rIOi6hQ6ujsC7L+KqiJ1A
RdYpf3WYpqn769XOut6dSB0YaQ9WvOtgdOwIUJRhb+TTWFVm74LgfPT1UF+y
eA0cbHwMUBw3MYlqrQmT7GRl4lXBNgD/lHDcmyZ8uWUtqjp4aaT+/ZMBePVJ
vpKXiPmNE2yx67gL1ZegrX0ZNJitRDKxuTRdphfp++aZVaEvWNL79j3sP51X
Tt/OVa6r+kyIYRw1CLtYPyQaZzZVdoE9JAFSRJDcPmLAvrgNJcSo+kPqULTg
zv7sJyVKx/34pH6658DbN8431tTWbxeAvlWXk3WCEEv4RYvgyHlUmkF/7Jo7
krrzPEdFnNNHmY8OCMjNVvig2Ac6ixPnyGQZYEH/U501Dxo7zjjwdHb2n4Z1
OVdoM2tpiM8lT3QRbnKLTsvBuljdDfeXmKpp/w0FZsOPGyjQ69569MVBL7ZL
W7bSrTdsO0i4Vy2mdRkDJR6ekwuw5RuHxS5gto4T+/DIH6KfSP+i4eRmr3At
T027quu7rhWp1wvgswl5tncrz7VTWq75cKIZbunZb5WLYT49F/74uQCWTqPT
9K0/fbcCJDSVeqkxLGauzWSxKYH+qxkgvQpT8WB5dU7MUWhJy5XJTDvxeF77
g3x3SX7XXbi7qJNREQWwJElxerrzCHzL2S1RsHfZWuXHT2UoNRyZ/pU3i34u
QgdIn0HKHMqoXGgkco3TPDomrnvqjftjptWvxyyH5Oyj6iK+psqGexHXO2wy
rJTrUqqi28mvoaCRlfFBAJ1yjxIQfW2nMwqmQtKPLof3aiUJJW6YqT0tVi7l
oiTLIIHS1YOJnfFvYxf4dqRJJdUj5h7uE11rfRwJM6uvxsSUW7qQ9EQWvkcp
IZmZ3Bx3MJERdWaTVEfRa/hI2l+q/nfj3mOxcOclo44kSCjqrAikzo9sFA85
VASwp5MBG6P70Jbb8pMOdD4M6hB5WAeLaRMVGVSG0qCcrY1QNG9ELY/cpSrS
u1JHqwWV8pMEtiih0ozNFogAPophj76uf4lh1dfySddjfKZ4vOhoOen+90EJ
jfuC2StBB+ozGLsInbUXr8l5gucLPGu1K216Ti+oXBtxjoNxfWB5vbXJEubO
jvlhOorkXPKHi4euqQW42RHTQU3Kcg0l1U3v4NkXAEMItoFDcLwaegnIfI0z
/JI4SFC7Iu+Xund+kpuFrlETldefJi3v4fDwVs9/ioowrOp4IEJgS3gRDoml
XRfCOftUb9cHWAtDAB62jwjDNLrKy2BMxXeUXS8ehdrOhpZH6wn9Fw272k1k
iyUL7aDFBywlvZpd9XrDA4J4Fk3f+oUY2u2nN1458LZtWwPfEtpbrBvwYGx/
b0VN3KG5EneJECh3JIG7HdjScZKS9O6Th0Cj0BZEpzPszU4DcG6bZgUPdaFS
0XSYWjdcJ5ABA7Y/Crb2CafRYjBvzoJPzOsR/YpF0/qMfhkTGxsFDjdCsCaE
06rgzFnnrdm/S6gothuTAyqadCrXQD6iddartQAkkf853DoH03H8WV0Ucdbj
Fgp3qZ6axHeG4pK/frYUBLkVQffi+KNm0nBW2JTOKHDxQBtSPiOA0zf4jwOw
4yu858MWByVHnWJvcDyB91prpTWGAH77jAgDhr+PInvZFXphGmJKgE4sMoXu
MpDx7ZfuYxkiKjCiPhpghQCf9DfEzUeogA3LPtKSfo+8VmSWW1EOSZg96x3t
ubpCragFeguHr1myHzytBX2eRz9QNWjcxgzM5gXWmRPdeAlwkJwpkSHL9iYp
G92g8A/aAfY4nmIoNj/Vjt+tjA2h8x52K6sAfrd8DRrC4+J89P9MVDsat6GC
PvDayEg5wWTA8L1v9DLQq0FUPHcPLK6fyCLSz8vFU7U/CHojN5CtUZI9fjZ5
Dlu+aJnarn08cMYmlrYbFp7BAamJnFU2JVT/5e+oPoCmyU/9JMWxa/09VQcO
yqWZV/PbBveNox0VZ2ITMqYmjIHbKWGNFm94W1ShsMEdl1TubHlAfEVFP20G
IX/8ICYJAZ6pX4knf5O9TSLli5IQ4GOjV0CNQ7d47yl2wB5tKBZ3+0iIAJLS
h+pqFS++DlbBBhAxJQpZ8Km+RppiO8KQ2rdf8eHjRv1LE0SN4mViuBu4AXbW
X5hBX6xIjj93HMEUJ6ooC1+pqJJbLgXG0HG4+ocI+NfcHersqcQ7UEN8axc2
tQowPjALxl6Z+aO8oBSIj7tNl5oBulKNllQ3uSNIHCNT1aFetlVzmonDix/a
NyxjcE9GG1gjPv4P6cOlwjG+DyUvNumQh9bl6qsKCTRzmKOxq33sO2lv1E7t
53qIb+BJAWi6d3g2Zhy8389swXgU4kK2wSXaeocjWnLU6bwlFWi0vj74CXhR
NinTUJI6lrZvx+2BAu1sMLjQH6/9XtqXf1/g2XXY48X8npZvlV/nkEseYAUP
TAu07XbGNQXIzX6fKcxC4wZiRyxuE7ASwNv78yRYoNTvQ3ayHE6DqTY8vJ7H
boBIa4aht6WRcfNGDktBfUPeeAipQcb6IBK1V43+8li9YQPw06l/GVN+nxzl
dmjLhAGrLoqi2WFX8Qyxp+cf32HVOSiYRcRpdrlmng6js1lZ1kDa7cZPUZNK
qufLu+T6chRaMEof+UyJ1KVUK6lMFqVfRaB6kPEHQI7Y4ot/qbH6qo1dXZv8
3SBnbeT23uuRrrCqQ58yeHM1AER20Rp6rjL/XanmS8Jb6u70sREHKBg7PtsU
LbrjLzhHamshXkNKra8/abCnWe5LcT/VQZZz5gHEDmaMrHc4vqul8PZIoDmB
YQNeUlK0Ou6qFmLqHXjx1EUkcJ4ClxK6LmRAtB3/FR66xDFW50URz446qBin
lK211pO47MA8s1Cks4NlVyqWNWZLa2vf1PzweQA5XXGvuewpaPwKndl7bqHK
w8slCxQotzhyMSzPtMFRg8jGtrlsHwAXS7B+ANWledYvUzR2P4NKnsPNP6NQ
DjdsoI47VGEMjuu41B2QL9INS4zhe/QrmXKkP/idZx+ewCgWbYbXUX8xXORJ
bDymETFRRVUUKltIaPzCsuEb0cActFJGMA8SXuTvWmWBQb6/bLyqXQjheEWi
IbG4c/mSkE6sL6MBiy/QjIsJWcbxY0zR28etVe341C/W4d8Z7RkSD0EU03Xs
7y1a4XI7lv6ukklETjx85aHQEuTHdnX1QtVsSuu7DI2/CHbTkcU6uzRQ7Jg0
1zSflWIlNcPCmk/2bOYOybLWbnBy1uMcwvsMNHR6YQ3sk0jYBRqKh8z8Ih9r
wNfCrx1s2h7fh5M5Iu3WNOe1ujfgqPUlRK/R82WyhQcYjKw6JXNJMoTDVA/c
ddZ3FCg2qeOri8BkVDxvi4di7HTjsl8GKI9W3ieYCo/KLTZY0bR9FEBSV/CQ
NH09v1mtsrguj2PavXH64sktgDRX98p9Nx7qtzCBgjroIpU+7X/nt0T8YSDA
3dVSocr6j6Jxt9sJSedrLRhNzdrYeGkjFjs61M21Ow/9odYPx5pjNYF8/sTS
t5wYuvHWb8UA2qWZ4j92DIiHENka+iiug/KuOuEkW6twdetR1K8qIb0qKMZJ
7YpfTwZC9HHvwh6UJt0F00zB3CRRxE1E95ii+rr2FQzd8J1DBtlqXxdxYqL9
Z1VTHw9cLvefwF945Z1zgRmh7Cq9Uekg7iVm1RFN7fkjHh18cCqadodLcFv0
4qDSPvwVMo8cZ0CuX0StZBXJ4onmNR8lLHG1UQPnla9Fw5sgSBIP7QCdt5+W
Gju/JoGV5PuCSrKaayR0XLtupP27BFbMKbYUoViy59aXQwspCKdkSSaV0EKN
npy7nJ842VvoGdRCQ7fiXpybpCbe8aCecs/4a7ov53y8R9tvEBFwRZQ87dAC
vlEJTva2NRtYK/1OoN5PWS3kVtc/SSIoCShK+T8Rsdjra7Z61H3lvqNsfv4d
bBMZeRPF3ucaQjmtcYgKLYxlDwXuGmz82QtSZgpq/2wHzaTeianOD4CY/454
TnWJS2CTcyyxq7DKJCfTaGal0MzUnylra/GLAvuGlM7C57noc7s0qmGIh2pV
0kvTFb7aynXKshP1mYcyj1T5b0S3y2qsaAQTUkmtscx2SZTJJnGR/NYdsHL2
qrCqdDXjMGpYFHHO6f0gjdJ2s5VHd8wscL2nQHFr2UMCTba3MbRDZqMgeaHc
lWRAPg6fl2sLiJ24r1JicKaDDDFf+WmLHnIy8Z3Epvv+MipYUMrLaW6ofEP9
TECriNsh5bq1gUEPOqvheDc6GGb3j+vuOtyuiZ/knxiUZhkMPFW/DpJGur/b
tW+W+wOYckZYpwUTpYqJ8hMVhTUmIAIT+MEYfBS7zqbN8/sd59jaF1/AWNIi
NueaVlYa/2wTgR+IFSd8STRf4ZH7ryecqLMctc/mxv3nGwc7DsZxtZDbKTCJ
FykwwYXDggJaH2IFcm6/zmmtQSOgWykwLpYjobDTmB4yCcgjMCzexbBM+Oek
qvH+hd6lwvbtEyz5U6RyGWfXkkPNcF6RQq2ewBnvXXrrZ0FLchIkLS3bGShG
VJgHERscMCCTsUbcD9Fa5Vfx4NMFzf1TkDCHep7gfql1992q+t/v2OJLhqiN
oM9driPJogAFFnMkrPMxzdz0NTlgoePaQZw0CXzpXtrLBazQv0MOF8mK/WT5
xuJYG0jv3Kd+feEZEs005r6Ql7OqXGjFa3y8Rp/XLTAaNYtxYS40dAVGcXIt
C9vhbwiLxqNHd+AkNDnud2kqW1ddk+9uYP1i5uIoDuuOO+/kNZXNHfVXCOLn
+7hPEww89t9829eUFXLhfaBnPRekNKB7facA/CtgjUMhhOHBfHgvoe9bRDom
+8eYJ4y6vD5GAohl2TNerZL92eLdlZlIOVQWtgVrAWSQ8vxpodozZ2REoLln
Ki8ycWMljqsFAUeIhK+2ZmRLnVcnKkMygLz+SmWftcdV/RD+rR3g/Z4Xjzvv
LmgemsNEZDNG/5AwEKkLgDtDtbnm78L0DbMAOmJyuUWFBMHQetQ+TvxX9IuC
onm5+1tzNzuAO8MHI/PwB72boluyj/EeeGgm8FVP/RV8WNZTiQOZurwQnQVV
U/MP8bRRPPnGscflADUL1OSUZfi7tUXr+YHDu8vt42VuwhSPXTjrg/+Zbv7P
46LN6D7iC5i+iDKCLCZg96d+ibcwfaypcx8vkevt9Cdc8iTQiwCKjTY98yUa
RvlscJB8zVdxz5yBysJPtk111NypjJE93+a5fFKuvZFdCLCy+w84AMLuNN0f
61sXZEk+GNX0+LEHrJvmL3kayuuC0iYha611upe/BzEtevwlrLKzwMAgwMzY
6CG2Pb9eskqc+pslWHcQchbS7Y7GJM0IVnJO6UsL8knuK81LArrcLYRSbCGe
tKe2uvB2RNYYfDh+WGYBzpaB0oog3S7668GC4MAFB2mgMkwchNULuHRHXI52
1W0mCBhbR91spDGvTj/RorUOHPXAnqzdYf1ilb0pRVDOqM8TFKH/JjQwCQsq
86KbqZCcj5hT1A7u1v50/eJj9gwfE53dl5kFU2PJ2By2uarrh9RgHzHZo8Yr
Mpis2aslFPg1QFtLnfwVwJB7FLcskf59CcE5aL0MfGncjRXbpsBkSg3Xau1N
TrlpbCvjNu4cmoJ/5fc8NUbKi911M9y09o3BkFhMZCOlRw9trz3mSaWSAOau
8P3553tsYHVrR5SRUJ+dr+83P0SxN0M/Ma0qg7+8bV2nRKU3QevXFsKhTrJc
0YlO8avlrdkxP2EVrNeHVzKSovfKaZ5y1d38xAUXfEvCLM82tdULMBoOBRKJ
WsMxT9X2fc3K3Ao+ObzH9UIrKiT8a9aOyS2bvIxVPZ7IdHyHp3xAswZrdRfg
sPLqfc330mtnDnix3FOPGg7PMDaaPBkoxENr8qT7KkdJiD99ohmxbnkgyAu6
nbs33kUDdTD7IISu1W/FA1tjUqhwWWvtAU9QtFoci50Nce2hWRuzySpqLWTD
IaaEzTojFx4PHUaf5wIxAh4RsaRei9q4bcNJvShBHyT3YOtyz/L+mlI4QA7q
pM1VoJJHfIciA4HKjVkK/+K6E9ePh7AKtDJmMWU4WZkBbMpKIf0uJACbw1gm
3hUOiMFNJWe5a2/vVZptydNvxiIPEly4XhbYF12oOjTwyeUUk3jfRowh4viz
reARaCwdP57ke9a0iqTfjSh8t5M9ay5OPK/8YAc+CMbsI1ECUHHYQTMSyZiC
+y6k6GOGfn+pcyAbJuka6r5mnf72At8rg8SVPOupd3Gh8978tCF7/0TWGFk9
0Pmzs59pI2xl8MFNy3vtYrhFsHQ0YwYHEZihrRsrfJTr1d5JtfYqPgnTEsIk
ojb5/j+qVkFy3+850o2a77MA9PGw8mCMeZh/Ex64mef9+HeSIGjQlBtbsQs/
UPmdELiYZAs334DQgUz/MkZLH+m246csr54UqXjPqia80ro8q17Ru2mYQ12k
vZFRPqSURHqute0vYpVMX320tMiKuNfsCUtlA6ftscpUSuvpAyz7JhBN8M2y
Lw/cwWDI3nc6HnpF0DPmit6P6B4yVL+zzx//CQWeaasoQ1IxVaUqDy2vbdMM
qlmnEe+Tp9sXFD5S+/AXJP8fzis1Q+uHxCv2gYr/YaoTj4aWMtyWoVhBPsm/
FW/lWECA/kFEDIvSYYWqxj40EtUWkEAtupuAvW/BunXGhZmP/xtyIkpPwEIf
eC8QUFMgdzm3y3/b/20Nxr4Fk93IKK8Y3oGXYpLOdWqjhi9MWLZSHXqu6Vsp
1r/X1xB6WGr3RafLDJ0tRSoe0anP73hp4fKCxkFeV27aUeTq2td9j/0ujwqe
7OGmilqiVXMR7gO707LZUP+J2aJ1bKD2lmSjtwQ0kESEwesSOLzroMSdkSVR
bVaT4X4M+TY4hL1/6I44r1pxRefH5IkFaP71nLyLC+m6hZmKsEUpPcqa4ey5
6R09HwHnToLEOMjEryTYoI+f1qi4qmiQZyZ+sGkMxCw4Q553LIgC145ZlnlK
k7mpsXv6+OJclsJK6A48pOyMnsZUDbMi39+WLiPzbQ+DND5Cmxo37Z6Gvat/
KY//ToGkOEbo+DowJ6jt+V0WrQuAZCcIZs+7gI/gQhutfNB9jc9B0yzBJFCO
HTBfoihKc2D4F6hXMGpDdANwFYEOwGLoirezSppWMB92gesqa0JfaXAzV3wB
7wSvqVzU9iOvHtF2yfQaQvomSNCCh0qG2K8mqcukhoRT3506YJBa8A+vLJ65
Ow4rRqxB6KsqKGSwcCYT2wEq0Hmui90SbZKuk40daDFqWd1bkJKfavzx+CbN
EnbjQwZYJcpEM2fCu8kgvLTQIeFAzQC28wYExOrWFICh/+HZZ8EIA/6Y4rFb
RDBRYaeMiNHpkxQB1vG7Anq8qX+o0bmldV1lki/Kct9j2rwPucP/7WzhQaQL
Gj/gZ0wGJtXNAqpT2bbPGRYNRM0jj2rCkUbLNZrN6mgXGol2w6iPhv6OtfZ0
EYHBg5UcG0G97RBgWHaDD7hqkmDj2kq1+QcoIYueOOulsN/gKKaVI1VCUWHy
WFrXPwo34o7v/TaLrgFEtczfE6K6T3jE7rr7AEu8lXCZZZGormM0xpjyrBJ5
ClraRqyw3JTsRNcwl9vgA1wIJ+IoituTGc+FkjaL31oxwupC2qiI0ACaPh7m
ms19/SjgfewON/IBamAB6pn+jbL76MBAQf4eg7i0q0hHT12X6MWie4yokmba
i6A+Ylj5Ur7qKEa/9lQJ+6qE7bnD7BG4rgY2PHiw6ABqO9aedhlX6XZ7CH9X
4GDrc5nmd2JMkro64i8ExUaAkDqICtZDSy9nzWAW2MBi/19g2XU081qEYVnv
sr2khz3N2ACWTeMc5x28WzgTZWVCsQE6I5+cOuT3c2V8EtDlShmjuLAmpLtw
218LirvX8cn3lURY2SemYQ4RgPplJ8Rb4axy7Qii7BD/SceBVlUs5yYOVgzI
APKvZNNBvZrBQLO96AMEe4xz5r7Z6tdZiSx3J/1qYOKoDm7pAeteh6WDyDFi
ousCDYCsEKi+Rv2keFQXvkR8dHqfLJzy1sFBwVuSlb+ZmpIiIze4K/F1Bk8M
3Oh1C+HD84ScAtc7m4vBscGQ2gm1Cnkut+evKD+0GrdnxUL5iuIoXTvrkyYG
Ud0hJR6ms5NCRf35BTo0CdZD5udj++QvUkf1KINYLjrzT8F4dPqHM60IPjoS
F9rx3W6h+2IRuXM+NsMkhiAdz9H1C7PMfVIctUeObFosynHBqznmG9DjfUay
lBvXqW9U/+VdTxEeXbzIEBm+XUBgpfgutJP8iUMdp4B8bgKEiKXd4ZSAOkEQ
L/Vg054ExjPLzWzInR9fneCxqIzMAI+uyZ2gR6w4sl9lFuq/946xZ0dv4H7i
R4xtHRABvKPrg7zdY9TL+Z3MXkAvq+7sSmSOgcBCqeCjf1yFQcBEayvigb6N
3hVblayByZ26GRHAr54tY8GjKS5+S0xFwKetjqsP+3+ghuDScUuQIBdUZw02
HTF7fOVOwupObW/zwPWJiHJMLysR5Z7t2qFixh8g2wggJJXedBZUPAEbZ92N
XzWYDFpgoqcFhrAij2CZhY83LNra5KWohY3RbeypJItz5D7DN5DmwbY8VQPl
ZpXHC76juMUm/MQif//eG3EhhC7Kzj3J6m08fygqBl8bwKUOfJYAZHc5bfB2
osZzjOgcC6m/slbDYrxLCvJqQ3WQI//SX+guE6fcBDR6NQvQaEAhsZnt1v2v
Y9jeTobSzJ8b3k0nfVw/IeboOsqD7QglI9RsDEQ54Uf9HfEsvI+Hm/L79FAy
VwMgyCdzJu0eb3+V7kbjQrA1n52CpopIhtOUgEnneZUs0DWU0LCicX/Y5R4I
d5Fo/zuoFyIaeP+e/NJYp0f/BzPE+aWr3eYyjUFZURjcIXUZ9UffQWhsNqaQ
p38OG06+qahoYngvUWo8fPnVRq6mt99WY9ZPtShpQJCtwobCcuE8lrfhgzb+
pcwotHlsJDXBiMAGbiw9TAHjqoKxqfCibCmy6akQgxEvEi9gOzCuWBrG4UNL
Sjj6sjqxkjBrR5uAM5S50YAPs7eFyVcnVWkuLRCosXALy8mMVMOGnKEXLNuG
C9jw9/UAQv76jrMLk1cFXvLEavjKLrE4lOIM+XrW6bsqPF6+r/jk5o+jA9GJ
6T9Yqv90RTRgJLNyjpAcePMH6Y9SagN+F2GLji9H7mWQPcylARfyoguG7Mo0
Ij3QBaQhTJ8W0enbYfyebHPIZw0iGnVFzS07x/fa0FsLKjwXSeEl/yTUikzq
uLe/64vbD1rjtmQJ/0K8UvsgNHOOYAJY1uAq8XCBlmvOR5MET3MhayrLbOrB
E1+MyBXfqlBtqQ2bL4HNLvzZqoNQlWdg731u1j5HiVpUnT3ooMAuZlwCgOii
A3tYkppUzRXAB/1nbOYNHCLDcAqlc2GzBwKRMMqL/LxhmkvcUv7cbHp3EMbl
WaLUEaZTcPlLpS8syv9Ha+YTDXF26ou90ZNgylGbJUYrNyyQ11MJ/hCZZUXK
ZJPWU0jkqGfA/7IrdjkuAjMDcIJgW8pZ5vIDfSNxcQzVSWitLC3hdHTq+TWS
9QC1sFGFKRHa4G3rFSmSgqoeBVwDzod0usT2cj9HONYwPal3itIZr1dYgM+V
AN/JXT8kD6D05oUcAQxDQq1VzjX3V6nDO05GqxAncwhvaF9zIPzb77keycXJ
gut8ZtkKOPQXiaopyBbBupefXAQ0mCTa/NqPKEEVD318TuI9rx3QG1AWQ/4Z
mLIoAFmCurFWCsdgrV3bF1NrAeoo2evQlC1N18jFZHLL85cB8cxcEQ2p8hVR
4LY0gbA/UUEdgUfQa9i3atnnHZZ9b+4fSJov87k/lVnCO4q5YvqedYTliQB/
rYCbBVane8SoAMbkvbQGsAQE6Yqeds8PFOe9xscMMl0PmZod4vEGTE8f+Y3i
5uYPTHPMWkt2fbXHRtRFdmKBHQ0Dx1Wd8MRSctd2H+F+q7STCyqfB3YSGX4U
bEcz1IdiwxgDOSt3U8Ks1fKRHASE04dpaLzG5+wbiC2clgfG3/3gmlwY0kFI
FRfDSg/xTwnkTiJwOUp6Cirl8juW2+7T/lvkiImIf7ToEreWZP3yn1vmdELy
buyfCMtJALJJ3m09A850EwcQ2Gpk8LHZLt30jWaSKcHQhPZyn+kZ9HKJ5Nzv
zx+9BN4AWwq4VYoHN+QPAbcVIaoLhuz2BEmNTKZszhP5J1wMiMkdTS/jTfCq
QhKnkgekkxKYDs24O3OMHyBuKjkBtQk6aDfMsFwerBS3T3B+ZnYjzy29agbz
LFnzz74jVnDSOdnQjzrOnFjBA8tf/1BTGvxvmfAbS1plXQgfoxvQTq3X1LvF
vXC1ql1RVz5tU9+41A8+d8DNXh+RUSXQ+hDUxyINuxgrcM2CYnMxn7+QsL34
AwdNVEdPIdrXs9PkNQcOIbtcxyRgbzj/3j5Trktt57mlPZ8VRvsL/Nx5viKL
+cdQ6d32HMnH26b1WAd4vdOg7O0bBGj04y107yfchb4Ca5OzhWJjIA5BQzvt
+qVgN7bl2kbcxGgR+ajZMalhFLRVnEXERvcKX/9OfuC88gdb5bNbC25NHEZw
nKPo4E6WOr3HzGqM7/e3YufNbBKjHBrSM3xys6GA/uD5eMr+VuBeA2xN9kUA
IjYFdwWUQFHd7kjpbkMOU0Gq7Xx08fVFKv9epKipSkgoTLKe8ko/WwPpb08m
Z2Ql1VG8lGCJ/BFyIm5GNKnRzbFEz9eoisWYfdvumOZgySZ1kCQN/Bxjgc9Y
KOl7qbhMAdN2shPB/y/ViazJQ2tSBEWIFr+tjMV//fQagCZmXKWp82sweCzC
wGpwyNHY9ESA62Lpg5qXy9pmY9ZuImRSCQrtjM+5PGkU4L7vFQ7GORsPExiE
3DmzANQo6SSdC+7QBnvusdSj65JOb3R6bIi2NRJElalfv4cjLZlHfEmzmW6Q
o1YzO3onF0sFaUdL4Cpjv6J6Q47Y2lwcsvb7KCcd5kqy8eKjKczcPgJfL6tb
gB2vfHMqR66i+hmV4Y5lggUVj1hrUm00A0UkrQT0osk7X1DKiWJbUjGk6F86
4HimUotNhLa1dLYbHg4oo85xMvm2uOwezLFf4t3T6E9h41wPPlzCRa+ouiSD
KpJuzzmw7pD87AAXsWFxF3iq3pa2sPH0VCv4+NWQ3qNT1aeVfC2KRa8j+Lpo
F0lY9JVLC7AjTWoBHo8MpXT4xOIIbMnbqbjpERcata1rIhtIkIXBxGSjeiU3
voaEo8tF5bRcngdv32k/9cfibug7Sqk9gsA/gcRRRUw8x4Z0pz/9+VuVIQ5D
PdOZdydxbfpOf5941nktcHtxOylor3EoWMMgo/VcUfnrQ9BloVykfbPvbMDr
LcBXKZQwTw9f5upvXfDQwujXbQ5ER312PcB/puiOONnrFnEVtGPEUxf5NM7W
ax1941WAvWsyRnYqyPUMx5GrqkbhSiYvEu7RXXcuv7A5Fu2cfe1Ww5UVUV0R
cF28nrNtCHshPQlP/rdumBJyzmO7FNVidNWRs+i+UbbzGCNqkg1S9Kjd0oyO
rpPgdBvWnOOOpZtMI1RVaS8uwqLPN1N1KK05dWWmMyt0jMv8Cxhf7KkOmCPm
Hbzk2Lz7Yk+Mw+HyZnRU0/YRx9nb1xtdjvf6FHGg66YIAix85HOJB9YrW+Zx
fYmW6/nkSOzh8/D/T7xMI+QZ8R5Chtnx10RJxkie/kT8tU5xT2e1LZDqx8eW
oO+qPI1KCIHiBlhN52Kq84FphVz/7r9/0xyxL2NREEqst/HX0Ah0z4rw4Zv+
291bW4X8Aryx6P03T8xza2h5E1789gegM/2Tg4T7OuiKkwxEeCjXq4wP1xsw
yvfGaKI4ZjtGP46oIjxqI9OMmFmNmEh8dF89509MBTPTvdtGKcWSU1Z5Y7zx
q0LiLn+J4EMEV5HsoKy5v5pjTpaPo5AZsSi7Ja5OF0wr+brTMpO9bVcFVX26
xlgYgHmjCPpaITalkHzOF8u6GRMtqxUtGGBwlrNMxaHJZV06+36FgNW5daLJ
wlhDzYcsdYRiB3oRfC2dSOKQmOTUeiCPIAekgRwmvAYyknQCajL3jepqDDnR
fhGt/+MzTaIAYj3ydSQHWlso/7iseY/rbu065XnEk6JS2RYLL1k2mqfc82Sz
hmN3KaiS19xyU1kBCVcKqQTYM4N8yv7I+BtV7UCKKVmnpW+bYUVv8kIzsZJ2
BB/k6IdzyEfAEHoFIBcN+II10L/QJKQqeplRvIWkLpUdjLh0v4p+b0ZbNXd1
Eu4YZT6ZdFr5NFweJdbrxyYuub3AAjHfHDlASItunpSLqI3ogbN1uV9PXKHd
0bqSZ5UiomLu1i0gmzWfuHkrt8DL8hvUJh2owSx5muddX/RvDq9EzUV2g4Yo
BeW+yzMutcoUTwpais2pt/VoXT6oPmlxkqva9dPzUXroObymCAoJkc1itJIU
+kAZjcXpE8xGqK1nhP+H9V9ZZPzzrHHit7SERPVBZFvqMm2m5J/NMjfmvsQb
+SvbZlZb8bGTLeuA+kZ3pFmSkK5fO85NWtqD/Zl4UJKIsnUzvYxj/XW7d2nj
4s9Z0G1ojyFMAhKIWPP25WT9j5ViTI39kRxu4+DP9JI55Ju0qs8wWkYv4eOi
tbF8mJev1BP//WRcG4o/8MeuWCzcljl9Uy0E+7pjMwSYqARRQNY95/iQi6uY
mQK+laTxo7/isH4IMLQrbU9ASBcg0/IVYUjQATpoGLez6xIDcBBHYmc25uBf
IwHbOso5Tm/42IDhzGWru/I6zk7YA0gcyQCCCT1DQFTBujoL4Qyv4bhPEBn9
AYGXshHalGW91C9PFDsUkPK5OMiQDTYEUQDAITis5k6F0GsO31EgXhuT3Thb
OMBifPIVLI3dmdXM8IVXlGGDApIM7cHXtNh58pRbk9cfuNIdt7dw3SCklpBC
AAKPaMzvxo2CkzxM7yWUYQrNE0lYdDH1MjFced6eptjsjiTspRiPmKbgI1nB
ngz+geHfYE51bjIbqNNg754mrH4P4jS2yvXVEG1G8U/GyfBSXsQkX3VZBL03
bAmSpIy1T0Y8Qkv6MgFXSnFfr+Ig5qvqbaXSjNJpD/i89pejJG7kyxSnX+Bp
XljHT+Ho6kCfkOTYyyRv03TdzBryK597MsAy6Y/FvXU8C9BFcptpMwNRKJrH
diTuK83CxE8ZdzMJLzU+KmLAdjqLJjsJ6xDiBJBbTdEE0YsM0Pmb/0TgeD9U
uD23VI35h1gXE7kkf/mz1u1txeAjPUmcqjwRMa3BtHeljrZ+6tj+nDtkD0Vu
mu3sH/GrQF7VmfnqDotIyTZ9HYXX1USvO00yLZCTn0674Zo69Bbw99v3I0Os
ZaEbv5OKY348QW2fnUKxllbkNTQSMDtPDXAf2HSzvN+JIqfGGq84yW7Ad4V4
m9QcaxKWQPr8uq4mBHZiDAMVfQYYHCT+zDy6Njam5UqsLJVv21bdnil2n4lp
vj59U2Qok01JhQdE5M/ky2e33DA92thxghVqya8JUmJbDgX2ZUTpncrq5qKU
FgXxo8tXBgv5GswAgD9KmXmXs0zD370sl0K4T9XAMAkTAZV849YSuCNaBL1Z
YcdCFB+j6fNIqQ+EqtzXeCnSeWrcn3l2qwspuuPUKUHTMyRVeAutLYYHetqt
hc+X49+EB3CryiYr+xQItETPmbLoQInvNkkQTapZ0dK4M1fsf3Vs+QSPboZN
WYDs2jjUfpmJjBEq0inj9XtVbPW8SiQUnxk8wMVwGI99hSd/oragRZh+S2rR
r6NHziwg8an54FmeBexuiBfgMzkE+UvMuDQbE2bNqujzS5W2m97ZvayacBR/
mLjPJmX0N6s4wUN0DGVOl/T7qYUvhhZX+7TYRSwYUKEBqSJrIoq4txQxqo1P
H5WJGJxACJlUBfOMKkvD+AZD5ZhJExcPtvEXq5NRYzB6ytxC/SuJISehUvsG
ljkr3XRlDCAG/g+ylmiuHEa/Y5I+anR4huBSmne95EV4Dz+MWOkE7g5U+Hhr
GNOKfrRgAWva7X3izMSoe/nTZaafQw4WpyyPk4Pfp7kTSiV9pBpaMx2Zu/Jk
lP7V6k5J4LDesHwFRZ7fFiWdIQ5Yuwm4+pkmt/eT1L0zX/KIvFaxLPLrSwcX
TOBTjxH8SrC6z4Esw0SHceBYmeDyNrit5p6S0l9sXNWMekv04Er7RcVLPLYQ
4TDcokoHDeaFSQa9gCADzTUGdUG4S9A1POWp27i3W+RKcX+F0QaYgAJs6B9H
aiF0YX1JIbPngErXjJhp5eJo9ZXFd00gpfqvJkBLP30SzS+l245QyziZOxgZ
6uOFbrhib4Rt9Q3OeL92Wp+kcxaLtP4XTNd76x/PyrvI6jLtX+oJJtwmuQvU
CbaIlv1pgAXYoLejTQwOFz14jTSibI1PJGHiVIi/fkO+5XNk5P6xX8MVMXTf
opLtZ4GbeLCxP2QLiQXLMPAZiwCKrmq2EI4sEwLYGrCxCTNAFygpYcQDB6pg
goUOP1QarI2u6zLptk2pZDIvFhbUfuNgBGVSncJCuYDZSdetSTfa7Xjx/mYy
LsfdFSO5E9KG5K8FxitCU24cowgyC62/2cBRfY7MSv4EHQKek8aETrHKCYsq
rU0PWQcCr/IbxtCIsKysxlqnQ4lxw2Z4w4Wgcd+4mcH+EJuBUiwdSnsExVe1
OzC/KN3yUBD28d5Iwsog7P4GH754fZOvZUGe1YCH1GFYcZRsXzaAXd/YJgI0
quwL75QVw1mra7gB4kmt+hSeDGKG98ch7Xz92gjWydaxEComc4O9aaTcYXS4
0SHQtggqzzptDzsrWc4zyuNeOcAXJV2yR4naQ00FSU+h++L/hoXDj8ISsi/S
6yqLyZMgAVbXPcqJf+O08rmJTC2tMoam4DjKMH8Gaw4Pipy6Va3YVE8SkWk0
OjBIlb7YaggjeANaLzScjvatUunEWbe1QW9Sn1E0MfO/U9rOc8jYdhXdai1j
JBXYJhk9PwkM3ilhVWWbUqkzoANMwiovh9a/8ttLWcuNwHc7Sjj4qKMz/Xtv
x4JPwROPJPqMtHqq14wK9PRcyNx9+Jn5lGJsR/SkniZeEepASQApvxIlJvXe
TxWbOumjA/ltu2mipRmoO+3u6LPieh/ThIEGk0+6m4cIYPjm8rIiWrmTMvfi
IxxVWSkgEIt+VdUJjAs+ijgk+yVaWzLwaCOmVnBrxPWwDto6erjR0wyjcIzZ
7P7djM38vVaAmQ2061aqoLKXgWQP2BPkdnm6N3IkHSDj/PwFZPlVTeUfnhX6
Lm+Ph3APyIUARYPGXDHSB1nnJGS+VYtcJjsLoY6sfSHmKmbo9dbCwCPkV/yb
Q3kDMeKwgECJJUXNVheg0XzRQoj60NuMjm1shXJzeR1KK+4MAvzmTeDHZL4H
eN4mmG3ET9QjqJMc2LguE1gevFhHqG6KOBrAhb3hEdfQBWhsIGL8cwEV2H4G
eluUlAGCw+u7Nx8tfnEV91zcRm0Txd26Un38kYkiclXm+kFmLoegj2JzHr6I
sjgMcKcsLPOl7gqWSVDMyQ9yDvBBb8S0FIbn3toFi7sawTjxgj8LEndhWbPe
Nb/8iSETQ87w2YW43fhM3Oao1EX/y+5XyCUkwrt1Rm1R/6QyweSf/A4qrLSm
B9vgLb7OimPHU0PreBTUCxj/LX6AlisyXW3yElIM6FdJjeVbc25Mc11TqUNe
557a8UXdB/W64aaOXeiouDWqiDEcWrEw2P1ISXbJzgeAs8b3jRvtPkQuFjwd
RYaWEgPg51DYe7gEa65MZFA2vPYJcj3VLkOXxas75K4R8Gy5tAw7ogytNzKl
JwRjVCGX118ukuXwc6JUaitKGdn3yMQzXQIk1MzdZDj2jRehYzNlXdri0hFK
zkh5UcW+MKhI6lj5tXUVX1mKoH8/x7rsX+W4XOqJ7wfIO9szsxwZeoN2HyyC
jSLZf3gyz5R/6bzeYPVFrgidyTmZy7I5HJ1/xGHGRI4mD0GPJiyWSsqv7J9x
V6ZcNxcaEsNccEjXCmp+fy4MTbpiohLsBFN8Ok0jDFKrUGZt5b3Hg2RrnLKC
EWRARh9pn8+Uuo5U7ipIA6i6/QOcnZJzilAM18fzCM2gXhpTSh+FA8aB8tVu
faoWCO1m55zW8HUN2LbHnULvighSku50K34r2PfxINcVr3N5iTNj92hCTTyO
vNDElOgqQIptJMI/9Guc3Birbzo7c+Z0ytWtGOlF4f4jcinjw78RxgCz91/p
Y2LQvpV/iYL8Bn0qWipcHPTQ81DKZmnEqMtVb2gEfWLmLXo3EWqpJblNj3x/
PB+bGsXYXgP3+4BGwo8YmbInkHJoxNuv8bg/VVrD5QkxU9LUVogp9wbFqkRE
Ptb1xZKufPRBR49Mf4RasRO5gDS5obAXaZ1UnV6p7dNvEYGPGPAhYax42ajc
qPixu0wS5UOUqIdr2kacS+MVinQhiJWYHy+fLOIBKuuRYrAcxdxivgcRT473
wyU3pcuvuFsnV9w7+K9PzFsJsLlPjiJD6XfngEvbYAvFF2Mk4Az9Nx4DKrmx
gd0SjczlwzWCFV6HeWr9MHRXVn4CCKT8SacTOz9oCWKnfgOrJWhoY3QnE3YW
+cqdWOgxrMbmHWk1i8gopWQqVdGbnc3LuGrKZDjdyxvHpM3nMEfLjSHPthG8
09+jD2v4Vu3HVGgWp8B1JmJOMAmEc8CXYb6pj22bJjBT5Kx2kGDT9Ji1o4u3
ah5mPfi7AxCN2NStX7g23F+kCAgYUCbkuOAZ709f91i/joLZAd48DaJCPEj9
TkxyXfY+a3q1eIKA/3dL+Z1T/WXXhPU4D5dyi2C19bTB0g4QNTNd9TWzm3SZ
9gr8QOP+HSTdZRVpoNiRQZXsHn22lvr358+FccOfUn/6OWkM6sdT+3Vw/GUZ
Txfhw0HHWo7MRgeX1AH9mYM1Cvzij9eajP8yJPt7DeHa9N9la42ea9iy/zi4
kwQl4zwbPtz6wm82BS7P18EqluaKnmAzWskvcvIeBKOA0C5/BvopVcC0vgO0
vZ02tzNe2zd4xIu6TGl+sEuJvQRw5IcD9OmHB6S3pQwTL18wENzK9RyoS8C/
JRRkKCMxHlNmxl9rtjD5Mvma0kmPEzTxBefQhtw64la6MoNb/CAJo59MNWy8
zX/FGcXICbiICSQAmhsdmMKoeItPMzjN3yTxl2atsGxTXwXaSDkzFyA8YhZf
6CC4uzVtGApyn3uiV2QOn9uvPUlFJ9BHItY2RKqHuO2GMw6UtSBtoiLpKvkL
9fODlKvwE6B0sT+JvbJYOT/ucU1UgIwqlHDkNDbLtShdaT5jsDGsPJoxMn8v
oNvjTsHoZEua+DD7u66YR8Q/5OCuNE4lvvwspIVZ8Ta8Tf3qWYH5HncnoSnS
N9vjpt9S6wyfjK56NlbqtB4Zszeak1TvWdHSZLnlLw+JDsZMwQI6bkFmq7YS
6X1YfLjyTRZk+Rtb7JJE9CPtU9k7mYHIwgcMj09UN9wHkKQ1/iJpviZJ6Opr
32I52mVhzlgv7mT/8/fIKzL24uAm7DwWz+topR+juetUQh9BOY4dzx6Qy+YU
y0fLeG5nIdXKlbuxKL6ecPVMb152i5bLuyIzkW5nbRjhVg8se3mYbrqraSTm
PwHU21kW7eJBEvIJIIFDDRU0KZzyWU8FMhiEF+gi1y+BVL/1UCRrk5crbduM
+jsrqaSCAL8JCXUBeltERPELYwrRpwdxY95LDITJkS4OZ8gxmaC9gORK6TlJ
Ff1tey2geMfWpvB8iccwySpyA8PZijG1DBQwb7A/pfNfUB5/sqQVwgfXJTgi
K9l8QD6DM0zBbJWWeeGKuay1PW5mNkw1KnELPjWtlOFnRqK+gdn9sC9Ih00g
e6cooPhpf7urfGVSOnKPgyw6QO3jv4MwzQmCWyw5uURLHtfEMXeQybuh8ggK
9gMKpZJC7S09BITS8ycKl3ElHE7fJhnwNhvQabPJLVfPSST7N7QKjFCqXeZr
bSBJ82glHaKMnen7Ki5G9JLFDmF+Bhq0KJ86J0RTUP0b9QrQ+PYUggWNXYEr
njaU3/VYTnRopGerN0jdSo0swAuPtCUqcNnZSsFqZPdL94ZotlDFnr+yTJJ0
sjfSxnqM8XLsMy78ghXJeIi7LIGEccIf3LyNwjq0kz+Gc1IyW7INzAoXhV7Y
c/PWkngkxXmLhZuSgYdU1pCBYKD8U3REPneis51MrJbqt3O6jEOeeib9p6cp
MSoMhDatoQqxWZegt4v+iqqMhV9jX2pmGw859I/ajnFXiHzAJGpz22UY+pmK
XUjwtWQj0px2GDVc8tvj520KHEBSG9j67K4CNdhb8ZFW8wKwjou4Y4ZRNZ4D
XVjJO26ISyJ5KioKQFUQFdqnSI6ioel7KyprKRfoH/3wtUFRj1iFEyipL7Zd
c1ny0C+rW7vanSF81ZyuOfiAyf2FW8ypucpaGoMDhOVNYWL+IkJDpGMyZuK7
v4lZNLEeLmceHmtLYOWnbO9M3a+mOKDTtCC9kW+/juGVeUs3CD3CvIooRuIL
5lzb7YOikMYkIO3YICKsfSkM90dCIxLaxnnrfhAME93l+Wa8zgzpe81hUXpf
mnRt0QRDA6QdG2XGgujvT8koXFiTkLGOyO4nyVATDx6R210oWw3Hsny+GUP1
F8ZaJb6+TROIUwxwfFNJRIVt2UnyY+hx4BZZiNJfUNawDqse9XvyKqN3ATpo
3A9t7EITRGuTeJ9yvRc06FxiQxeic+kRUOhQrII72j0u1xgOko9PCFBO+ol1
+bNeJ5TVJbgVV7XAFagOtGcKrzNx80TuwhUIAu4TSDfqFCZ2Ecn7Kexwi2wP
0rS5wVuIu9A8C1s6XMcytPGsU4PeFI2CddDtiriVjJYEfeoe09h6thximFU1
K8P4ifDUkLlmK8dBi7GgIb/5tXs0yPcaJCTD/thMHz1syczlgm0P1IpAwqVX
JiGDFQH8Q7qecmxxoH6JzXOp1sFUaw2SklhOTm8MowiWX4vIlPcIZJC6LweF
grr1Kk9G/iYnBtWmrjCPwzfZ9niuCr6RzxxtxRPLsXR1+3zOc8rkAYQX/Xrl
LhHaNwwCDRxTHEWeIK3MBvQPU3jCDhRksw/J/PFiTX+KK6mnTEul4aRoSQi+
b/xKgAAzwAfmYvvkoizfyePiDK5blR5vF8LzmQkiIhx1Io4HI0GEvxkinubU
AQTBBMFxk5uL0l1kg2xxGH0qkSCXSoeSFnN/1gIDDJKQEmtrwb/5+K5F2mQr
EOOlrYTcK7GrDn0uNNvAOAddkelqVskHztCbqD7MrtV2F97UAuUaRmwHiXQ9
PrWhmMVABxmajAQhH7+4Y25iECq8v+OtjFInKya6gcNSq9Hqf7EHJg+R4rWv
hSXjDQdX8xCg0VLNZhbYGO0StZ8v/PAWs4z3c8onGbHd2OJQyib7C0pdMdGa
t4VnC8tnTJ4twmZ/nRxxAlvJ1aU2s1+kHcOsshSbhM6k2SXlCSmgOonoEzgL
e1NFZBzULVipoLyx6oMxbrnS/u/xg0qxdwE8tT/LT5TZjqsL9xEn6iHyNRji
y5jL2YWjRE2hOgLRtcYofY9Nf9TIPX35Izi6ZyrHfBK2jm5t/jiEG6bX3H94
PVJewJzplnPAqgfFMSmSdXOz5V3umFQCDvrsvrpUZOvMsZuTSEW9QZ2Pbb/m
0Wx940o7TctdQSGUIB/XpXfBGkxVNYXjXOu4jFT6GzZFaXHtc29c4a4ET+Rg
C10FADUDWIaaiVxHle4I+be75Ha7iBJGKIOKbMofvyLXwkwJxUdaFmtmouG/
bKrsXRdoIXQJsUJIc0surEGHj4PeuhksxGSQyn9cWhXHKvoDSuRcGw7ASMFo
8u+bJRt1CMHogokbkeJCMibw3tBoWbVEb3qsaPoFLu8Ldp5VlbGkw+CAwlWa
v3Qa/m8oVtp1Eehm1mQ3ttZOYtspTQbXuxhiXdX0MJp5i7oeACaDa3N2emfq
CZRd8IvTak2kge5dkjevcCju/GX7HSt3RLvyt7BWNWxcXcrkahEGCWpE2gGg
lD4RBOgzlCsTS0IZCPo9we02ukK2FItocwKQkBS0UaX2NcuSM3WS+qx98F7V
PwxvO3v06kj34rx9F+7diYjljbtQk9A3hlPGlukL0HNYq8Jz2cpsuAd1grrl
VM81BIRIFAIOATWaWrhzfxpqwalwTZmRylCVP4do7j0tqj4GeiYETcWofZnl
5DDnI3nZlp3mMnjXslDF7OJyu9SYkNme8cB6YYnAbPIpXh+4Bx5+NuG4Wrac
rUtlFMTz+YZLI1WC6ovs7ck5Rd6PiKRHcPhLZLHgmwFDZG9vRRk51hIKG4F4
STgGlGgonHFqRRt5CviVbG7LM/DFGq/gNkv9fpgoij4rXPZFm7Jjuy1T/R83
e5+9xnxv10zSHxDxTaDZ0YjHk8JhrKiwSWp772F13FdzybFK7cxCWHVJm3bL
RlCIYHPX9SBMFPs9b8Gout/IxdOSBkVCElW+uEBQKY7XS8ss/RgbP7xgPjqe
LcDNDBK3OOPm8WLH0kxjum8YxRQl1ntGbCkog5wOBeEsdj2wNFfHaUn1thC1
te4GVXEgryLOnDKUIm4dTPp2NF02DI/eVRAAOnEcrIEIulB3gSgwf1F2LAJ7
mkrO3kWWlOrrH+pQa3TWA6aHW0zBo8rdvZ7ePRAVQT0Wk/OP1evKwseB64QZ
ib2fsI0t9ARxudyquQW+PlmrjGHYAbzdmNO3C2uT39Ueghtoe5nKoWDsNgJX
OOvTSV9NFMd7PZSuLuFtpNqr7QgFGRVMnojlbOZ6a2AqBvkzMOR/up7fwaCb
NAYCkT433Bgb3X1kpc22KfK97mq4TVEsPqdtr2lr6E7TJFaMRjVCp2sA/VGy
3dqPF6fenPQQmh3t7gkeoLIL6g+SfuKfx2Va6dT2HtEsNhS6w3JbrE0HM/Bl
f49p5FZqzfqQSrDXdTvfNeJ7Hd0xE7KGq8cXIHl7JYhYgl9gyJ3VURX+DbAA
/lzN6KwwKsKL4BItKqJkW08DOKRm6qAiK8rLfUkl0EuHxbDYA4rz6CM98nwT
LfOisjc5P7fuNce8rGOlFEz4Cs8pWBIdpK6WsK8C65lZ9TSvFij6n2nv12Em
Pi0W1gyo7nxWL9a73nalttbsE1fp7jRjh8Sgnh7A1PL0IjGn6T3FaLHfdhDv
I9KQwUjgLOVDInhO0mCyMXkqVH/KbtyCBsHUnI58EaLTA3erbglhlEVTTSdU
jlT6cNN/eieK9U3kUo968Vj/pfdFoXGYO4wW+plKwB4HWzOTT6c/5aqEVlwJ
MrfodpPmrKjCRWZvXIrt65610UviF4OrUbH5XD4Ka743e875EXyGsXjrp39y
4fPZmmFxTRV2ksle+muQj/IaUAz5NPCLrZgD2LT6cBriK+tpYQDj/bhII/+U
keVln1jbPLAI0XgIFS53twWHOQrW66YIpBAKlmQTH7M1kaHmPb7+Ut+uwXfI
03YAVkktXOpU7aY4r4RKYu7KGjyCoSNEYeCgd7KxLZEUb8vvTxJCiMLXcoYb
FTnYtFQyhlSy8KYxNKbMl0RHW0lSBWpDYn7sV4gYUftxukn83tl1aS6Pd8LJ
cI+83sGa2XEPBwfzfGh/hOtwIxCK0khqYSy1ARJHDsKAJlQ7u9JXZLvtFlom
qCpEjbOhQAHWlfJA9Sojs9AX9zIPPw5cx9VFkwo3f+BwCKCWC1hNDTSvhN6e
rik3cZ17F1XmJNFtTJwOsFi5KgdCZFxdNShivVk4knqTeGWgImyDm3mNwWuM
uOc0R1hyJW/3UQun0cT/+E4e1eptZ615DUuKzDDAi3vYnNKUogpfhf/jd7ug
dNvsO32NnbH0VNRTYFMk9drVQfp9ITa2IYKc7kpo2T7DB/kN7b4yBW1B4psQ
djd09jW+DtKdy2EpYX8SR11OpxvQt8D+Pw4E69eKW5dUvsxABtqSlv05CpGA
1EHhZXKQfbqhdxlU9dlXHxCtvH8VLN9ofXM423O26iwiHcRJphNM+sT9I3ZK
LSIVdu62ZINiLSc6KT6d2REB+l2AN8PYxApa4vEhQZ9KvLV6sQ7+v/B4t7WB
CeJPhY94vHA5Du32tqsO/E/QTt3/dqXDwQMo88EFLVOgaTVgtGC74xIwhlnS
p3Fz9j15X6hBOZn/M2h0sonGSxyHl0KyaPWoUVectfFUkQOgOppvvngprPr4
I6796pajiJQDkHRKJx1gLauoGA4HpdXNMZPSJdAyk3H/fExRazEosSvvW67N
KW4u9O/LXMp4nvgXJfV4QCeT7Qg5+6IpwJxBucaU5N2ngxEHstSndOixj+rj
d0Zs1MKsu6scHwcgU+QXiIsow0lG9yCvzX/2Xgg/83xcsLNyZG203VlCr4kL
Q5pRb6rlg5W/B/bvaOgr6znzGBm5/ScJdE4dKyHLrCY19JQ79sdODu7Jy34A
N0Vdz2cu1y0GncsEccvJwCWJBUxpQ9lEj5PgkIs8HRooKVvER0/jfVGAVuIA
ru+KvRoxiB+ZrjaZ91DfRq/ehO9/LdyEqvR1Pu6ECMO9P2NhqfzV2BTCenQY
IbjXI6VUSntzLANGfMUQvGiXH8XhgmEbpZQDGuP6JNQG9htsH0b1UBb7EWyC
xFUlqcpe63GP9ZwOMCC4gis6NEG4pru0korMqMAjx0P7pWiwET+qCs+tt9oN
IldlYbRqFkJwO+m44HTyiWeNWwoSJrmByB+xWaIzIJ69oTS7WtCs4aEuCbDa
1Qpfj56ki03S15kCTW3aoB5kQ9Y681k413OF96xIwnScNrJsZPQuBqs3tjLY
UCWtjOdj+WMQggAJckhwB0SL29DtrslrSSqvFy2l3YYDsIpcrE5W56LgFZVN
TvQYjTHk5W0O7z+mCsrVhNubsZIcq78+3C1a2e5mLTtLraprcfUCtOjesCgK
ZL4vQcQa9mGJEUkijJoSdpm6MYzm0yGcrS/9vPLeIeu74KKJrXEcvKux1U0y
drc5Y98QF5b2vFPrg3QbK5dhCJ3cAgcPS0Wf82R8GwvU8QBgBKKz3sYUMCoz
VIMv5iiGN+jdBZvJOXC5L54b2VXioDHx0ItvpQBRhFfB4E/i8FV/jMeaNn0r
O0goZaRlAz+Edv4UA+JiX83FhX0pUkvuGL2nhPlezapp5P78Njn2gG5zXZvM
dYrQZyYzWjLoBW4KzfXLGGOHjRvm7rIWlKHngG2Ftzqc836y4o0MzdG5wtbm
ZCCdxlkY0S9Jl+BYzFone/0U0bqbQ/JKtu5163R/ed9UILRbdEit6M+pQem4
cXCpTvU2wbL4t13gz9SkGtv8tN8wF8B0/3949uFpB1yWt/QtCcDsHqgoM5rM
cTQMjlyLL0KX+EfCz3THZSd0bp0fbLCwJnd2ST2Z2X2kEt2wodyulCMeWfPU
qpPll02pPK8VHLXWsf26zsLZx9cfoNeE1THux0HycLXO1R+en2p9vMYU/e9t
p+yq+c46rWzGMuVeSu44D+CEcdtbGX3EQNKAM0zYZ/W+97WI6BwZnbhOFJdm
+0+4sLLziilMKby2FZEl+SVV6BfugdVnCdalvmDLXaw8H4IDnH18rPfLWX+F
n0WoCrgCMmRrl5tvk1DMIq3yA6t8zSdkauPtnP/wrnLTQso/RODybVXEJJfw
Ua07kNtRa97lUdQB/saBm1Os/Y08VN3yA4VRq9kUArxKyngzxK4DTM+0GTjY
UU1BYo8JVKP+UNK9JupJ7LAIqmuGm4wAVsE9tB5XfY6Mz/PzNwUe9FGiy7/q
/GG59i82PUhgSPXOCZsxgPzGTkAb/hFj188PdLQdAAp3wis1XGzOQXn3hOZy
DzvOwpd/DaYzbZHxJqGo1Vwaoh1yw+YLxnhqw+UtheXtcmYlnbGNsJTkF8u3
VabI6g9PLSClJnDJk7iUB9jQCG7TzbNC2QllhGq6a+UI94NRVtTsumgRrhP0
XaegmHWGnCKpmM3uWuL769B6vhjKhj+ObyrG2rrPK9RIGVDJ8RByrorC29Nb
dpGFOHQx8rOOjPjGd18D0I+i/avGt7hHIOGzSgfjpkPLFttKnB2qYwhcc2JP
kI4c+hd5M40e1iGvh5o3eiU7vXlyz5cSB8TLNpZBeohtZMk3ph1a5AwJ8xv1
veTlg9scj5wJhVC3s75mBhysWWKM0CsD3WqT4BBZb7TSVVz8KNcv9pmdV42f
KFCezzenRBk/wiTgIw3sxzDAN9nyuFFYx2rP9D/9UaNZ/dn0XPrk8jx1dLKh
fnyEJY9Hma2jY7PRl05G7xk/xJVys/t/rwFOuNVK0Y09A5xkyRfQQ+8+9Q8w
xeUKZNcU+bXfwjl0d8GSMDAqruzTjjI3nmNuXz5tnoiEUpjuY/cgUzchIZGZ
a49d7V6RAJxFm6CQvrVmJxGHdvDjZSazPsstH5Y4IB+lSGdK0/iaVJl+1KgW
zp5IBGWz3D1wtPGnYyPM6GY7hDU6qXrqpFXcaSpUy9/NTC5+Gi/x4N1oMyNT
HMzyysGwje1YXyK0G/QFWPhmWFBJVtNBh/NDMkzT2qiMNVBm+WJOTyko6jik
t9PM80OvSslYGNulm7fzzeGrM8Ugp9Pcns8vz8ch+3tKWY18jTIGXPpVL7jS
vsNumOGbrM8NPA2E9LCQ0ba5Lq1OCAK/Ihy3xyiiqkQITzT+sVmpxeSIg+d7
8KE+6aJLFfTRKmQCfk8jWJvJHfeyiUXhR70e8TzT8tyPBfK1McWsquI2UFXe
gBVINxmbq97NcEwqAIXz/OWyrzw3Gqb94nV81bZKCVzZeMvCAZel+nyhqfp6
SoU8l/wJasV+qSAAyYRkl8v5H9eCVnSrORst4xPB9hjik3BPPQwfgEV6lw9g
m3tU/TRsoh/Ws4XlMVy/9PpRAL3sZ+UU9MajvbqpOJSJvmGVrajCTlsTDp4R
Zx4fsuLgaas9mbQsZs/HRlgKa5yh24IM25AIQ75TOu8BDzIP9k9OZlL9nGLy
GVAyypVeedx5bPZDNcm6IxCUaql4Z5MvvAUOidIevAQ6nPnlnFwo4PjXCnDV
FsD/qCH+crSzypNdN+SPgUCOZN1J/oWAY1DmEgOU+PEOOrpSyNc4tNl4ogGu
b8tKjTCVPqOjo2F+fPd4vUQtHv3c+DGYYu5PcXDMb6ExplxWD0tYt51dNB4A
kkAKiZ9v9GG0y9xKjFqt+ACc0vCQF1goJIw77uEySOPrPLamR6KsDaawQ6z4
95I2hX1nhXvk64YI9/EZGavQz8e8QArfeqsAChxPvoB8CLHH42d2t1No9PAd
uJs2w9Y5Kr5QdGo6uwhHkYpOZIKeAy6gVG5Nk25kpxBUqEw/73faHNt8RdVZ
rwgIGJJlp9jQ5S0V/8YAZV5VQuYhUeZIYXMLN3OBNKMW/Dx9vr+Xkjr9YfyN
d5KZB0sbIzPqFCCiSjrshd/zvZoiShrXzySRsGfY4VTn+wy/pOeL5FEg0IVE
63qwknd0DIVQfrA23e11+7qkX5HmvWx0MgxCyCfTvyViC7DUnGHc6+oVyJif
B3D28KUawQ58orKgQR4JzapFaw8qaHqQZpqsBMMwmhViLRVMKOJkbCMgg5RD
jD/rTbjC1pLEg1D2l22hcWoFor3ubPPpBVXUWW9Xx3qSFuFd9CE4paq8bWnf
52XNQjQpbMPwRxAleXu2GDHjDcNjxJ6LwOnFl+fvLWVCCzgq5jzS0jgTXWWh
moM26XqyA2V70umQl8HLK484fsNT3rD6xqKdPgwyyFkYMhlffis+/+29dfaZ
bn0cVdtc7tcNz96ZDWNq8cczHWdS3EKCdWHPXwLY66tO3ZLFS6ZtUtn7wSAR
pI+S2XrjgRliMnE93NkVgdmnknLUcb5k0LYOp37Rs2hoXLiww+DEtnI+Q7rR
VEK+ENyRt7oH29KrUoFCLG6GghozGALg2Ge7bTvj/IQeNAdT/KaEIiW8Y1lC
P2kn3F8t8pK6zAIb2XuTtz4ivKNOCSpceKENDDzqIN1tKUE6JDh4aG3bEguR
OI/kZOtmsitXviJNAsj/BCypYUk0tUARh2tzhEJHeErcTL86QkljCSFIChYY
8mDnr+DePqWg585B+iErvMQ9IL7LUBDN30quzOxFKrpQmR57uQcUeThn5VR1
YKKApo+8dLpPQvwxdzPIxWnzihZmxuqGLM3IFMwyVV6moHzbUr4jtPxFXZ6Q
eu2+YWVgpQ1ZzfI0a49mxR0uw37IUDfOv1Jjau9sEzsORVrNxh6u7Ye+XqCg
r4V0pyxe8I7SYSmJcsz4ubb6Ms4sxDTdVU+EO+DcZ1DYv2qtuRM++2qSlkIS
Lc4GbivLeF1+ziHbnahbADhACPAxT5eu88T7sTK5DHdMjoAnN1pjvnfOD2+w
jGtyIJpyjCh7jPqxHl3HxUWGsEx0OjAbmrPBUTyp/PRedJo7sHcMcahz4Qby
rG5L1Y4h3FRZnKLceGSs0heeF+l+Ph5N5Vntd9udA+t49NC2a0xQ/05bjmOp
kGxWOuKOkazDw8b6yuFiADKgflYzzMl/YVQcwUBsZHqmNAE+lqAkolpDIolI
/c7NqR2eoIPIUdSFITi01oIcLSfq1FRmqB2TvTWJpGENfc3F2c9oHEsmJjVi
WRrAAA7z/bD2WisfwueZ5n2ftko/cLvapxKkhCVu1dWR5YGbVRAv1jD1s2lK
fMlDLwSJax+REjH/pNAIyiRV1kHlcE3ow3+qN7PskQtJdgb440loB1qI5/k3
zdXTBWu+OfUsSn/n4ANr8nPi3qDZo6raYP2T+vikVfD2K6rHjF1IHn4bxEy1
xM08ES4IsNzPXoIjka/7SQHNHgwbsP6CVRl5tg+wNgttfEUKFtEAGl17V7t1
1NOnfQLJ4EiisbiKluCNLI98XccWuv4kmNOk81XwRbXo8ZuJ7uNmq0MbVzEP
yKW/zc+Z1xM1SN7yCKtNC6GPGgAsWRhBlW5AuhcOX+feY4VF36UTZ+BI7MSz
xZCfaGlHz2uotBoFH5S3dsA5poAYkj72FCeVAI5CKT1GAChhN/Eh0he+QT4S
OCcilqVDmZTYuPwLS3iMA4+5eI3deJtLN4aUMDRg0KMJDSds2/apKMF3WG5H
Ag9tLmKB3flzA4/9BcoHg2+hCA433Cc81xGAZ79GPmpzteDCR2e9VVcFADpQ
Rqr+VCpUW5nAPQzDRdCuT454x7UJUpIkdSRrAw3bxB5a/b6ppr2HegxGG1Jy
WUWZUYSBGB7EWugr0MsSmklNKN2zTN0eiZ8y7w+BeaJBA1chQac9nRqwtdGK
F7YkP6k3Ipokqda70ObgkeDJeg13bVVGiFgNEezlGO2NzgonimbhCR4LkUae
OuSttoJ+ytvNu0mUs6RkfOfi82gV3SQDLsjbHWXw7BFogxYlwrn5q2wuAtNN
Z2BJbMs7ugDzHQpSYZF5a3Jl5MVT6l3O4TNwO8wEKiYd7ophY8LOt+g0GHY6
bihlKgkRVNAdITlm6AXjYIqu5nJru82eSDe73dTwb+1qKi3fw11TNlJTA7TC
qTYo0F8F4wzwGCxWxXYhNEWxoI7oXsWMDFst/r5fLiS6coOScAMW0slZTTO2
Id52cd+QwvhjVaDJy7NkjEQmtpEJ0Qn06T2Ey3im9XeIF8P/aHhiyujWDQoW
3cdI2UbNmqA813SMeqrSI93QpRVhv32N/oNE4PJnKD5yDTyoKLLfhWd/cUZB
oJdApradUEDrydPCShlpQc5xUijHjydm0wt00uAD+uwCP20/y8+a4CyRXytV
byBDSehD3QxU/bGgUvA9s7KHkEuv4kGr5KxLCxYsU8EpHG1FKQrlSEdzSVLi
c1mXfKB0rizOpD4JL5J5mwGSCfTDyVhBpa8o783fYIbhpeBTiId6OEY9yJZD
pXxCC6Y46+NbhZns46FlFd1wxG9cGfbrNBUd2vr/hvDoRH9di8pdSqpHlxp3
EArJ3qUJmt8hZYOq7QFA3cItJv+8leLQtrtL+jCu/0VfEV8P67/OQ7sdhk9c
GcKJM5He4Tim+Sd4q7AyLjkygOrpVE45QgRzVUjtN2eRmXiSsx/y3wTJWqUB
PNCXStjFxt8RBWDOiwt1xToDuIzJzDxiOa0hELUbIm2tmZcoKESTUtKSMBJ2
SKsKqUEzPFWPi+V982gh2O05xestfA+YXEdXAuYkYisO5AOiyox9gcuRrHg8
NJME20BluRJ7JpVwQcQPDNsrzcwR8rHrxPiB9pzZp5geekjmyWaMr7JxrJX8
RjStG8M+4Lpga+eLBdeOtQodASFR4VdWUCxOW23fy0IIQPXDhfOxuzaZoYY4
GYEF+o6XFSzKkq6ULKtXnwVqO+66qKXZXAupaNwsBISlBj2tVeHGAbBxeHny
/5wSXlHopmkop6XWqnrcsg6lec6UWaZTL0vqAt0+q3L44UMGZEaJ0NckAYci
2L8R8F9azfZss9u2MN2xyvqkhJUM37sdHt5q3manslIM94ysq5Z+hBhB+QoT
k0CV70FEme7QnMtqAkcrsuBCFROqgP29o+TBr6yyQhVy6RRFKujV5W4Nykvn
FqneZ2Z7z7cZeJwiZkqs61E0SV7qpahllOx24cMJNZg0UgzwryDSvqGFh/rq
/Ub3VVmK4olC/kz626nQ8g1ugDbE3H1t4fnNjAtjLtuZDFO4SGUWFsN3V+37
wO9yx00DwzOLTKBMYQdu3UMajFwXg87cucA/iva+dy8O7dhjjHmTQJ5RDPwM
T5BsNwLrTNT7Jg4aB14WwyijSTxUq0adxM0YvNRdVlR45xgnnOcc/hviOM0p
18pbnQr/aUrB0z5Oggm0vVKjbeZG9h49TVkkf82F7BSYPGMcP3k3TEOVnFLs
ryrXrp+QRAPN7Pn2Ld6BYCMsRvLOP9kB0gso2KBk/YjCgkHiUgIVV3VQuTMS
2i6UTp1BjlzkcLwxdxSGZxkUm8Mw7FWDUpy44nxIE+N3kdVfC+Hu2UDMKLON
4lt7StB5rwGk/GO3qRpaaTt5h4lTINuuRlNNmnEoejN8WTuSyf2IXDtKfByF
4ucR3CIuba6pRNYFDWSDpKIxItLSyYBXndSHCLRFIg+MFwLF5iqoVrsqL6K1
JH+n63aNnWmNTCt62qLx6IL51CleXNG7R3Wyocm+ObEWfQ+HuA39xcDbdmOk
VYv0oKkfx0h2Y3zwBoJ6VarJy4kUIYAqd7AnP+tEPDO7LGbA5tY7UtP4GAXi
QzHSKAMX5loYbckaSCMHw76rr5vcsoYL1a0/hrOKTJc/VDQZ84GZnNrH9i1q
BzAYZmvIPFI//7gcz34Y3coZe7hFT00oIfSXADYJKMahh0SyN4oPYO/Q6Rib
8MLJ2xweaTYy9g1z2KZcheouPCALKzXZ4B4RK0I8i+Eo31jvUinsuByY7b6w
mj4Xe8SbadLxPgOH9WhGMAGYzuinUD2T+nr10m7FEHcvIz4Uti4e2ctv1pT0
sio7jlbBlOg+ZTLCdIugjIKotgcyOG4WGi3O0ZMEM5or7AyI7rBiYd80lFLj
+tUGEp9NS3l6NyW810YvKBu/qE0M5pVF2iY8p6OvNVMBuf2xrgfJX9ad3lPt
WL1JnNgVr93I8tIMI6QYAz/aFALuZQGtdeLnPBDqZ3nBRP+3KxqHvHItwwir
SZGVHwb2MKYANRrEZefSUJvicRQJE4K0buNFH2gVGzphEldqIcz+B5oMHPWE
RedpXoB5h19T7nxAmjtVTx9GQtei28mtWJKZB1Isr0NY+FzOSYJX0JeMlRob
jhOY9494/maZy/DRjEC1BLuzqlQybH69xjxNVbV3yX3fW3Q8ArqG9TZdUZj3
gDeQpytX2R3llRy4t65Hr+LV7nXvFkuclhEA4fw9sHl6Wfot1/78s0pw1/V3
f3xv/ok4WMoN19t0O3ztz9cn1vcocTLeLyt84asiRXlxC1W6DE+JuIgVp+JG
Q61AC/WOz6qMqGkbpc0/fuwA9hOrufd7nrsJfYfdQPIDaMWdPG2kxFVoQals
0aAns5BwIJOXRPZCVxcPmk5aj95b1Oqe8LOEBiJyvmY7SDcrKR5gCZCHTdsV
agWamDe4U9qItwCjJ0Dd9jZpXlU9960qv0MuuSVkDZ0SRLy80X4kVsUEn8Qc
f67aPeUlMO4TNlevauM9HX689V7Sove1SVCVspvMOAy3zWZJDZ3fxcWoGJUf
OWbgoJkJTmNuC9omXYZdGyXNM3XbddvM1oCYPcSU9WdrS6kSdh0RX/fKpM+c
9tz6kAOVa+9hVAnSBkJrRonAfEpV4qO8oiJpG6MPHDjI6lep8jYQxwmx441u
VoKHgFy82+AVXV+bCh7UvKvCdz2NgkL+SGwkuHbWw1jox/V4COVtDR4JWjlz
A91lIxmQ0xO/vYhAvJ6u3rgHYgraT1xB8aooI5n2Tncc7Z9a+JQLO1hhKEDk
MgtP1xZGbq/qS9R9gphYewczqtsDKu5ajd8tD/4akLR6uoOe9jv/QC9CPqLj
A+XJ4YlQoxugFJalKKCMJW+ybk/TN80ZYzfdrqzOWw8Ece2Uegs8kMuRcuBZ
WORT5R2ZWJVaWJBtpvKf8kR/pYot83hkylbjaTG03bmXG9jNQJAx5VYxUoWt
A2z8MrI1hEXUglIrYimTbGIf8h9PzmMvUZuTgQWp6PCwaYbOau/u1/epwFt1
n8qTkczVcwEyieHyyFGrJ8VgUxlDWemlIBnUyf/pTFLt4B35Z5WtTZzvauYI
sCGLgWteIikKgWH2i3VMNt6dmoWffkHbaIZqzBqCnF9X3eooiq7ptKWRwx4H
rRhqOZbOOWVakHHq/eUyUJs6qG6sq+jYdUiwX9PWWyGj3/sfWD0I+h4GRwfW
i1hroBoREQlCX1CWo6Q6Rr9azEi+b2CuCHZZ/paRbuPs4NEHYL9v198FNlZU
dMxvLf/x09ycgv+fnBU8MlXgBe/ms2x1CauxQT6mK5WRHUFIzASxvwsNpl3D
kibHU85kn1+UnABN/ZpfIoZNdsuZNCKpDsn/PKKm4M3LkVaWx7aZiheI3xtl
lbNCR+cJ4zWgrdY6OQlUpi1TfIsEI/CiDQFlMoDQtNuoYEQFGX6tj6IwkSE8
OuiDI5MgSFwLnNdX3RHg7e1qHqTOIMONtQTbYTQv+/vVIBhVURDoVdnyfEW4
c3iwNqGKdUxIDEJJAj9VDXip/cnONDACgpfB4CMGsBYQ2hn7/lyIoWcBOwcX
IhjAqoUu380ofxNWVIr6I/yvvCUSaasyLWdNvdIF1sO17ECM/5vWnQjZrU49
mVGutLIPoeO53f/tqh61alhZB9dicvcvqst+37a/2ayOOM0GbVaUwbygNJK0
1ivy5ns6J3D9yIKLRqPWsuNtXuED42RdmkNZzGLxwg4kAqonNWo/VEMYtKo0
2xpG+BeTmHmzx8K45ltoVvzA8L7E0uQ9E0MEIvJpXhlfJUr9ghYad6DEJfWx
6+XUqEYovTwyfIWyle4ytb688aC2XXRfQL7sZbE2+pTZ815ub5muqe02nGLR
Wk4TZoQNfHcvKoNuTg9AnYLstGq95ibi6UKc7himnXBYF/TGE8hDfWkrTQmP
oeP9QaMR7XHSs1988SZVEv98id+2jhDz1Lx++gX8U0RSDazZCb4KfgCvRdCu
LgeZt05pDXqqUyDpD0O29m0E+ISyg+4ECP+uS2ruhybLC9IFUk88nK+GaYuy
YgR9VfSJ93OJykfIfeodOPe+BeGBUaPgfEI5v7ssJtaMUIOblMMGvT5MI7j/
hilGABZlc7HfxOOax2WNu+0GGD5NeLmvS2pUJobczhht6JU9G4zzu3yn46w7
CFfnBLMh856CzxMboCo6fvtejt8Ap6Cn/vjmjKHseEIgsIifLK1UXxaGoUYn
rBZGLdK2uw6AAzwQFjE76zhy/uHaPDSdTG7utG2nNtVB3R6CQPce4OXKWyeU
WScPbrAJhV3tF2GMpZTMqvLXmtwSmv3bH8m5Q0elckJcp4w1GWWwfhCRbt9L
QJshVNRFMwhw+CCg8bEGHkBJ+Los9KgxndZWC6saK+oJeEazWnb2sCuig2gT
IO0Pfnm/nz+0soIS12DuzW4/X55Pdg6kCptyXhaHpnyfdU16ckHlYdiE0u2N
Cy3cHd+dcgYfHH+ehmaGq/RXZxcXADyjG2hrhhyBg7OtpkqRr3ZsRa4VQmJ1
cUbRZN3KmU6mtt0JSzoliD7CeD2r6RQVRquNO7BNTx/9pMFGNDSNOoapffCj
4CkLzM3MHlJG9baEAM+u5/Zm8yQ3d/ohPpmIm1IklFd/NvpTe2wS9hPtMu2/
UDldlx9UHmpWfIfpLkC3NzuxxGNRuwSz4WbErHh1sxz7BGgsJW/Rk4id2EuA
nyjm/drrnwflW14Odi/YB47AQTSICtCUgW+ychi4ytFlV/7wPzBugezi1gg5
qTej1G4CvYvz1PnfjPyUB206dQoaRvGFTDMRTWumbklmHq9ioSR9+URUEZ/K
xv3oEbIc2/1JbSnWfEzLFp+xMpzx7NlmkkknTyWMi4TLEa2MjUYga3rDTEZw
DwVrxudvse6224cG7vmaVTNjjP51JrshirdTA1TNoSwt78vNZKB1dNrJAUMn
8ioaaqgAXBkA9dBe0qzBzTy6PvV6TpIqqd1VNAykFQNtBmqRJtQtxjhKuDPo
7Bykwpw8tZ1Ll0MpA/rQbgXYOsqZhSqppccfbKGJ7RDi4RiCVWZ+qz6UXUF9
NDP1wbHXRIyCxDog5V0NZ+/yFSi36oTdjIrN6gDf9GcLIRPJkS4PoaqwkWYt
AUmdP07ERy9X1J6HOCeSOxERxus6C7tBhQk9Udg8aU1X7rWh3xDXrlNW72cR
x7Yq4VKz2B2Pi3ZoBQqeTV25RhLG22iFGOkYqX9uw9hZ7s+dtVxH9TAyCciL
ALTcFPOL87PkWSnrCcr+6ZQdgRqBpJF07aHC4ep+eFZVzmFIKR4LznJyOZDz
yPyKmTVuX5PEhqdDcpM/YV+KztN7o6un8XMDk5jC+qa8pFjX7enK9B2Mvo5N
+UN/U5p0rhsb9i32VkUuNUXfvmcV2+Py84yjwA5XGlVkZCMzxT+hSyYfIdOf
/vWvnhMBMCeIv7auDPeXhZYySyjZBdySvqwsEOQrncZjMOZuaOLLW1f1wWpc
BFG9l+DxlSGyALKbAeA/zhPQS8To+UrI+Jg/spRZ1N6f5VWWo7qVZpTES7bd
4YOgSJdmY2neyaU7Ukb4bJfHogoFo4pDm/HtZLbHRKwmUg/Xyzdp9Q5A851m
qZKBBHsRmmvF7itvICchTwnOA9AADqsiL1co2j5BFC2uR7xghGyRskfnDFdo
S1IH+e8gphc5/bdtXQWKJ1Da/Q7hM3Z803rsRErzTvk/3+zgxoOZeENDGIs0
5YVir3+6vR5gYf5DF0OMAhZaWtLOrd0Hpl3dkD5yyqiIqoZ6O29GS2KRLqtQ
PACF5tp5HrSsB4R2sufqgyp2JS/2iCm2rbAbkVO7pxJoxEK0A+nkUaD5gBH0
Bn4m2gjACEN/JFdEb2xDwDZdP4Ctxfv8U6Mq5PvdOpKIU9nlzBqugqHeLlov
9jPdiMM9jVoBUpqyhwTuHH58TwDWUTlii7Vm6NV9+T3CLH1+uWWxJjmTmPuT
ufL5piyqe9QfKVe5ey/itw122OxJmYokUif60w3QBeCL24I2c8uFY9BAzPns
ODnpJDyXNgtxvpPm3Ns7HcNaCewLqLKbq9PmBhJgon+TSOmbP5Q+coBgb9Jn
QpLhEVXL/7j6N9P0tlWtwbbGhBvh7g1pSUaM05mGJ2WjJUVraIhQxzzupAPc
yvqDPSLR8M2QwDIh4BQPpCwpMm7SQWItqhFl8wvdc6KElJPtwbuZUnyM3w4L
T5h5WEdmGlidUVbEbpd23DyVxCuShDfz+7doKSFfM/zwH/HT6zIp3hSwCfvR
uX3Ev6BZzC9A7JFwa6+eTggs2JVcpA8eExj6zO5un0DknJaGtcrN289ipabi
fcxZLMxx2tSXl8oRhejTNnme0bXor3xgDeq4wN69HZ8e6LsMbQolP4uRJuLN
QbvKPHG0XVJIO4zl/0Fwnqr+8/bXCoH8/vVCRdSiMgR1cxKO5l4iuBbmYQhJ
18jesjrCACZ22nOmUhm1osfqAMXL1gaoMyLB4smzpGwu4QUv8jl+FHjjwNgo
T3h2KOJeLYar5Se8gwpolq5ASBbskqyX63hOqser0PlbIIvPVuP73ENMjwf0
+TwYfFVusowpdryIQmV7kF8OWIOHpeP8y9D+48mUQD8JjhnysUQK48A+kw06
HfMjwqavnMi/NcHQlGN/x8Ji47k984Fgl9UiMKhhpe/UvxG2kgKmWGSdvxc9
hvqBKhkc3VaXNxnBvB+p0K3l7O1d6PbvAwk4hHSEP1xqeam/W3o/7ILN/HwF
NADzBsyb+uL8bYm7LBWiG8ePIfPwEcRMDvNyhwaIjwU1y0Dj+X1TlvS4cH69
yku9Z9B78AnLj/rmU8e692tvv+1OXg4tXqEsqBRDEHyyB7F9Sfwr4j8CSboW
X2qn/FWqkL/pfqVohD/ZdGAHB3sBOytXEjHsCf6tCEmrHJU6UkdpCs0XdJbh
N19FBQAFhUpMM3kDoDIDA1pIqHOKQmqgt4h2aon+oTq95Bbr3I4rB0MNjCw7
Y4zmWT9YDptTEPsvQkC8rEJGfe1sNz4f/Qb/+XOn3ZKU1qPgtx2cLyAKsZXr
Mo6h6kNcUmUy4knerOVKZsuk+x4kVzgmQDZ2D3j3vXJOYPGYPsxrgQ1qmR+1
UFrSy2A56HboqgNxXjBpTWWa0MeuKTaj9lu4dHEg2OhvZdK1ghgam2bUUybY
RGOSc00Gr8ckW8T+JH1F2RTKw6unGDnpDUjyUD3NCZQ9sZhNV/nen3sXkVGB
rHHLHCMhsjUW5IGwIbj5hGlFvkSU8FV6zH4sJF8Q4zp3znJspJlvAuaZGumG
wqgODzz8zl0EBUczTZFMY4EY9SD4AbXE7EqpgcXprQPhHrWkoOoB7Idaeai4
+1BWlOQlkAjE0o8TQ9rhSGgbb8ojg01GvClcmWhu9GKsc40qaMYXo4g0ePgc
u49OGZ+VxFzig2tgAON3uZo02JWVWQq/OjSUAcAymrlPlmOs0j3kKvU4ejTv
lT7EKEy+Y4AfjoQIW7u2DPmcboMtOVGdAs5+Ibbz7hX9iZDB24j5vLW0Ltbr
5CRyoKizgUdcxGy6plGaWlVnDszxn9/u7CO40QifYfoIcRXHcGpwH54CPUNJ
CWR6nNpkep/D3KauaJr0bCAwSwaBHndL4LP0jQdyCP1/i2As/fphNGzjdqfL
Df+MVot+7mFxZItdhAlvqHoDTum4BtBzkx4P1iVt7Hc3bLKSa2LNgAGbVooM
iyn45U0IQpUbKAc5Aj18006NPovprwkfzGJ0mgGrKcicZj7QhCK3U1n18KW/
N4y5zKTWWJuoR8KODrMEjU5UG4xiguWrpI/TTyVtxH68AXCGAFyr2EIDnAIE
uKobBN3+SE3lPkZ7DSKlyoUiW/aoyNvw74BF9nHXCtDD+mWdxMpzTp2/5vx0
IuWUynAczNZiqLg4fO+I1IFwCfKwMz17jgykveeEzaY1ghKqssTsUuOdNrRV
uFTj90L615T5rg3+H5k/lvLSSVhKq3ShZc5uUoDuwjJ7KS/LK9lkrCHZO2m+
n0w7w6cv9oFVcmNovaEmS0gKYanGYEdj3n20a3SjE1Bu2LVN8j5JYMAddhfC
Lfr/y4liVJ/vCZ5zgQW5qh59jeCkETS1GRWCLYTobqhN+YwzNQPHNpht1CPq
4DbnsEJy0PE5y68cZG/dh834izMq+6id6knqC/NH8SDrpF+RJHd0SyfeU3ZP
b6iTKxKUwAjFyHYMYZ2e26lnj7Zol6eGeiYKj6FJg7zPzeUTN4e5Ur5S9qsT
tOz7H04lOKMOXvUqvvEODyupfAuh88hU5l/8YyCFbTYe8Mngg4yTVcY9LI+V
CRUThk3+i7HScbrlO0MYne7CFtO6s3TO4lqvdmohbiPd6t4ysyXwb9b4tPfC
avp8kcUsQfai7JUkSZYN5lV2PRQBK8aA8Xkdz3LAUpGOaWdx5wCklOkuo1js
T2z+HdhrJBYriG84+m0nbbXTOwiRkmBR7qcxonfk1gfluNgpyDYMbXMQa7V8
jtcXDc/F8T7bT82vA4w+ut1aD/RbWxS0V3Wf/zFykU8C7uQsGyD3iHYxLdiH
gIbIWpDKqQZiNcW3ugyEOfxb/PcuTcone0AXQb1/sExM4tDefmJZ1imMqzOK
9LcIlbdyM9vCx65uhERqzgPTxOxgooQQv87D7gT9GPShppjftpVlrSWj1ca0
/RP+Cnj7D20HBr9Zdz+z5QGhWsvBW/JBYWmKDTwEywYHz1RpsFBGO/LiF8k0
6srFp6JQBmFaViCGvzTzH1BC2eYnc+nn2/hfNXgKYip00bXCSMZqY7Ib9muk
G+0jVCdjw5a8lNWfM+sXiGcRGFva1chbSZyta18IdDZyln3PadYTJHgPIRdi
Za+oj1P1sxc19IMchmkXaEeOidmh6zetIdRhA2unpF1j4jm+5PGZ3P++rwy3
0klPwcAdV8/JB/MSEbys3MgJ7l6PSc1ktI1XOrg3id28jYYCAKuDg5JlHg+U
Cxj0x752VzcuH79aXnmjpdhZUNIBs7fVmXZgQo0TO0WjrAtSxrmZ/7g/0/hc
UBEqljqydA6EqYfsHtO6acg/66Isp1pfx+cyE0pzPeYYgW1gsrp4vkbSBbJC
H/r+09j/PfOBQMGzheEkHapFH8zvfGZNYwuGn2iF/zXZ2ANyvLHeSw4fUMss
QM/v1DRTmQheaQtGFVhO768Kkt3bMENlUzL+UE5rgvdBpXGmy6GRjL2rxRki
TIDGKOj+99uGK91rUFvQJRYrqM5BhnO/KGQ1Pi9WW5ISWkCdBssA1w0B1ydd
c+XnaBBqDVsDHqyhGSQUWyJE+MoqOpJZQN1qdZUFRH6a3vBrCaIj4sFNFfu6
x/7Ny4sMdH+E7IzYJIX2d01X/EM+Z9hjohE9FshZPQ/rEDutFmmy0OzpvP7U
w3+NdPzjNHZ7XmV9a4UAOm69y6iJhTqEW9bmS8Ejen7SCg/fkD9rGu9sExoc
r3+Th5OTP4GLJgc6Up6MlDICkvUM67RXsmbjlrzsuAZryAlPNZhYsz2/cBmB
/A8aRl3L0AYqVZfATQBgdtedPv/0sNohRF2fN6tw/gO+IH03D1jW028QotQm
UmuMhGEXAS5hlhbWulBoX0UEn1GEaNv9zn2j1pFvFtSlpEA4+H7QLNdVskLl
+zvpZ2+Tk0oEtKb+ljoXiuJ29jeHDZHihQe+XS/oNcynMzQwTz1sLPzflMup
EeSMf3cIt/OOONi7ZaOo0DJH+hScuNcQgH8G0f9mBjVuDawu13dAkI+6rm0z
RfYnEfdW2EVk2UeG0xt8o88/ff8Zo+VAqmLpbgsGYzsB5bsBurdPXIa65zJ6
JLTdGb9zGoCDTzY8hGHIYmEg5RqaSd2mZ10w+EeKXgRPJwDRmEvjd8tHdmI8
U7iOkF0DLA/jeBGGLKiZJBsbNyQYK8i0GjTeRFGcMrc6SvfBqDg9WInvab2V
86JXtyBIMqG6xHNF7whf+HDfGmWfJWJROUXoYhcYWvmM64au+gfjx2ul7FQN
Xfgwas1X5728EVM9Di5vQyoV8DbG1PDGkaboJCvosyn7AApSKa0xDD8EepXI
/2gQESyzZ56YfCPoC9So2q2lvafKGXgr5rgPtHAARLfPAupO5STk9m+y4NrA
sSankYO8sI+unzZCmn2TSTF3ZfW6dXo+6PyhpCO34ncwAWvfmYH56Jqk69ID
qZNxIaFn6z+0z0A2HTyp8vsvnv4pskMBsPbVkNHgerAw86ClY6Zt2xf2C1sk
15xRHxYK44NuHcZaMP9zZOUZTNaV7/PfjTq3MpxLsFvEIUlk2/dBMCUGq4L9
dl+3xDCTPc8OJ2fThTPrhNPWsJhB7NdExcehV1QNcC/W1uB6+pR0j1blT/wl
IXvu/yFcSDGx9UE+3szXe/RDn8Gz3E9HeRsNEjr4mmzbCqAbQCQP8eWBp4fJ
WXgLKEG6D9lzdEkvFxIsaAUQsDHFpvv6RCPwewr4qc7mcNlW0MSGjMuVv/aT
oilE74dkJztCLAklySzjMH2nSl1M5W7KvzOzT0z/82DOaONwNtzVxjOYcJSL
dNYWnrpXjZqZKYBIgB4tnu41VkOe63+QA7/GGKX8zPkyUrGP4PolTG1L36EV
94K41uoXZlx1PG2Stae5sdoNN+t8sfcd2QV+f3tlcG1zQ1xmYT0FabWOdkIv
yXY1QKGIcXc5sMwRohjKRhZTkSnwZ95kQtKveqiLmBM6xltpm/t/dek7VZPa
mGy2OhPrF2Rgx6VC8F+4p8YnaYZJAJp3AVmoEjUP9COL19Z+ilJDW6HDJmH9
KDhtxh1w4CydIMuSdQ9sksgWQz16PPaTNYN2IUGUQBoulS3ekXsDdjagBxTy
XNX3KfgOTDVHSQuRFZT2xozaRvle1SGgxq5DapfHFCKjm0lPqN16b8w1QJCe
J312isoPKnvIiOFHvk2H1Q25OwDmcwrq2L1mAHUScHW+5mdDBcLZqkhsjXW0
ajPakgiz/pI2YIZ75kFgzMMtkx/03vXjxSVo1AsLbiSpAeXBO1ssc55RegwO
8ytqs9zyNfaU6RIrsY2ALCLkSp9DcxDYnGYbDAYLjsl3gaK5VrfKylJ+Voi0
LcJKVRM3MqP2JoFB7C8U65RGVjHadiN7wsSkGTAUBIktGiCB0OxHAJDzbCMY
/Q360Xws+6g+WrNf66eNzYal2T1LVxCuX1526ATDYxOWcFLBe+CJo20/3RtE
2/TtZHu4liwVNFsAtQ7gbKyEiIlcOhBLIJPP/7a/53xl7P3pUMbfllOZb/Nd
GZlqn3hZlkoJiKow9E4ypGBF+I3LAHUY2OYXer6K+urP2kBU62yRClwIa8qG
J0dXVEdawEkBTd8UwM/b9JfnpWmn9rN5A2gyW5IWM/2+LveoRTOwZ1x5rEWF
rxwJz+pdV3uupJW1EILjVW9DX82laam+ObKjpGRj60Hn/+s/EvuVsfaAuSVM
KDZA1r0vqBeSzj8BImsGSwB7ZgkJ2hc6swlvMxWw6rz4XZpIHJcC5L6w6Gv8
QJz/YlAgc5ro8szzatUp7Y8oCHU8OOkBxg+boFuKRUEze8db+NENigYdzMtD
Qa/2t8olJrVXJfwkOr2Xj9+S7YI2+RdC1869uTa03Gy2AL9k9hZZCNcUTySw
z4ytto0kWgkUdTHZfwCg5s3IL6gGeKeOibjAL7UWlSD0XSTnpqJzoaPmboih
EVRgyXocxf+feYVW83jOsnH/RFzKFliIrFZP51XoqLYgCaquHzc/nNuYQZj1
QrfqIfGYtWV5s8AtcS0WeCo/TCv0zWlejYkwqiJ+n7m2DYmawG3gbNQLkyKB
U0wjugmePZ8EB9rrd/jrF4IlMR6cAUKmut0Mlfq+x+zrYxGWUl2g5A7jpZCM
0kKXA4ucRxUSuyxniqzXcNTNKO1iuM2vGg8e2zAYNZw3Ohonu7zVMWH37bf3
AovtseOUeG43WTksmjlakg9aZaYUkyJI/e2DZy6dWOLTQ2023+nKlTdhNrLg
luTC5Y9PyR1aoPpHsk716/T6NgiM3od1dz2wv2ocVpvkA2x047N1yOGcHlEX
GPIJ063fh9LMVMF93QSSu2LL0p5PGRjJMKWZy+5ROrMYoH+6uRtwrWcVPGET
RrzOlYvo/m98dS4dRKO2zi2MN7HmSD4rkGHU15rYLJ6fR3FOGSMu74F+H5D/
OkI8ntlPEKV5DQp+0GPDnM61q+5AHavDP75Un4pOqW/H8I35ZS9bWskP/OCD
gLKAyEU9F59hH8bHz6Tj7OtDvPfjJ0tJfSnzcMw60+BceXNzVxKERFTlTc0Z
AXSmlliU5pB1NfDfN140vH4ylyLCm61db+dqPbI4glGSWeTvRvU1aC7UrvJ8
wFnlS388FQ/9eHowcGCOCcPXZdFRH4IPa1PDKd1Vy57UtGWZ4u7q0uzsAd0H
TlKr8smN7mCDKm3J53pKgsErKgWK7dE4y6eEp6N22OGkhngUcRnJjPgsrrFM
3pXrpyAeElC4u7yK4ezu8tS/NHQnR4JpkJKKkHdXOktbkntpSek5AxvGdXqn
NqG/WTqPmoe120ZaEu7Es24O3wGxfIgJlUbuKS8dQNcdf/wVlzktWx7gVq7L
kreWcUcwtOru79AdoXoPdK3pTG+Fo17QEs1x15duhcog7ocErHsF8X+t69+N
Nyd9RwATdmW3zxUiS75zHWc0qEdRF2Msx2UF6IycHcc1Be4Kdl3NJKz3JM3j
WjQ4iQhQJyU9x+y12fM2Sr70YcQWim2SE+qZSU0mOTYfHUI2z6v5a5MiGsBX
RsfGez7KruVV4tQkKArhZ9vUj8ncTwQXZP289cH/VT2m4bGfoHC9BMDtiMiz
u1LSjmndICyd49mZowZLQOJWxm29UM+ZIbplXF9pCn21saQlZD+BJiDelzhz
yMzAhLy0oydlnXvsfYFeDz2BlCw/4xTn8KRgOJkk+8sImuEj3FhkuU9nrf7Q
B7BbMqx0xyBP2VMOknbRr8RMLqBVOjiO/cdfCS5LiES2msKPQ20XEG2d/Wnl
l1OZpr7Vrw75By171coZDhUdsG93d9dkuvNBJLqh75wOPppEz3kTh1XmWPsb
rJAyB8KGy6P3yb2zyDjsFZyI+6WLXqh4lQoINlcADUIrGsVycxRA1RHxzkrL
piUhvtw88XK7AXSQQq18LNTRqLfDeLoPrO+08h5dJHfdddKrReVTbwtFpEUx
nJo8tQyGK+npyKv2vmtYq2U+8flsVqmgJDLzqshXeN82/YAjc1HNbXsqPkre
OMdWzLyitaFgJidTcL9DngJxlUiIyFqyBLinV5mynmUBeV5NlcmnCMenj6yJ
fihdwmN/ji8JPDEjzq/axOwmL2PXH8q0d9/x8lzB+Dg+eyhDJ9ja89rrFpFw
VA1D+q3JbyL3EnFN3YrAyjkqQVpv950o220EaRVc+X4nTQXnfyZkE4WwiHNA
QazLZuq+tModqZ6tv1lB/7PVL9xooU0BP9uNVfEzwufWlO9JFKH2vGv1sqkg
szG29Tm2WZ1+7Fu9Pnts6PTkg5BUKr4onT4k3b923TOBt0TZnKrxfaDsBAeX
lofmLUWF4RwlwUVMKkiSD4tfobbK/W91cnwBgdKEnNtDNI1kcngmpiy3x6ET
KVgnoKyeqH/wC5z+h5ize6rbhXMZhsbDHQBoZaCI3hYJwM1Mr0keIdnt0UaJ
Os5DniQ3tUEmWeT6lOo+CCImAQfkdy7KNiZAHLUGK8Vo4OKsuiaui1GLHqYL
M5jWqH4fzBPGXO/8xqG3owKSSpu8TkPTJ9Ix3nK3LXArtl91vXjW8O+KcLtK
OLuCQtjY+UGKRk+b9SjYfzzeZ/lR9h5MitfQ2IKEuI91RrwXZn2nvwdMmQZw
xQQJ7ZFJH7ep21izobPo54SxiGrBgzfp/r79mFWeNxvYlkO/91/1YHWh2Snr
jDdl21N3wiEvWNSyha1uJ15TqUyPZGPYBp1sQYoK6B8ZgekLYF8hq9VS8dbM
GcargyOYs+/BB00Hqav2ErmePkx6+au7mqNBkch5Dy4i33w0tyCbcpMwMsec
k3PEoByea42/CsA/zbB3dEomfF3+BTgKv7UFEEQWUap6zoSr8rjKJK4SRFyD
ZTvES51lb69D2YzYV0HiVDFmMpm/SIfEZ0baTW9MS78bl47wwYqdszHGC+dZ
d5lE8MZ89vy5BsuuLnB0jAZk23up3FrTxasHMyaDCoqpZR6AuZpbsZ20LZQ7
KriDXdnjwoK7RHG4MAY/NhHJgEBXxsu7YO/JdmMFE2vymlPYpju5clDzl6dd
lUp2kZCiiagfLao9z3b3pS+5HgnEI+Sx7MPmdvkeimtan281VwbmhsYhh3w4
DDaCxmR3aTYB26gTRhAJ2FqSrYqjoGaKVXymbgAE6nB137BUM9zOQ99oSHbv
hVi/k524aQiF3Dr3azSEbV5R7KUwqix1VrEccNsxyJBe2Yhx8lL9+ADVO9XT
VZV2MIp/mZOZdXM/dR8u5F2J6hgJnMHfc1atwww3PwfJnZyQ0zbWhEoXJ8jd
rqd7WbU0cXkxr/x3F/w8jZ43yulvW12cy6EjlPcabt0nerSV4WWuRwZnPqBr
qDMg7OaH6kRgAxG73iJIwDx137b+0v1dIjo0xcDiiG+MHDFl17IvuJTzI1Zj
dh4g37KdPdENblYpOgUzYfzkN+w0hPj9iHyAPeoWYSG6I0FPbCdIsmCcgKxX
w2PgQ1NsgTb6JlJvWeo9W2UlbquZgCDWxblF6Im467+pWBfIKM0wzqMNTk9X
8erqtLg1xQ9rrTLJ0Y6MMcf6Y8HpnTMXOT1vwtHh8pl4XAJeeeI/Nhhqo9Ia
qggU+UFy/FNmcHEQtx73kg+JLeFWzvoYmmOZfrSVrQJg7ziJFfFVdanJbA5C
ih7Il7/zSJKn6+ybPXQdWgbeCn3qMQgTZGaSZ9+JqKsQBWihRN8NKsflZP+H
jG0bPC3zjGtco0+SLQFYKITj+VMy5tNRtQeUo9Y27EvaLfZM5nLGebcfzIgy
Txdlv/+AOBfUomXi5Zzy5MtOWKYFNhHWqarofWdm/WTQPPHC8dM/l0rIYz4z
mpPyDzqMW7PX4tsymHplM1Hy4xhhius2euiPgpbknR++O9WmfP7fLehepz2E
tVcwgZUUCtA366iWFssENHbPkcbLmkeFNMO+uz8lucSVrUi2KdvXSsrqp1BV
UxxeyBDg3hDSY3tXQFKZZNBgJOpLdDqGgDJ+a0SgGrRTWiF18tnDQShDEtkT
HGxjgJRMcwY5rI7SMETC94jhyZSmDzM5j5N73t1T8Um/yZPyVe7HuOXy55Uo
efDQyoFT9y9kk00fa31pKkBmdBPl+vLy5OkP9zeDKqao5D0RRU6wKFKD2lmS
VRvNbStzIIQeEvqxxLchizxjWlLD0BlRVYtG9S7ybBqgU/JdmpYAM/oYKTE8
54wBgvi7zsRawM0nKUI2nYKj0ooFJRX+OTr3uu8argNBiZpqgBGRBFkqw6a6
MnW2FV8439JPoMH4VJ/jGQeeq+Y2B9uzU0p6NNSpkIujdFRQ8sotzvxVkG0T
jDjeYqUfPgADMbe+kNdbRDpbcmR8c49bwvoVPORUzLmC8InkvtxYZXJnF00o
zGhuQ7eMPldlvU/UIAO1aUcrom58aC883u6FCxCz+TxaPTQTMtPEKQcmysLv
lL58CsgCsmV0zB3xidwhBZfAN3a0bNmPm9pXI6XEp4IjuylX4jn1cMWDItcc
F8R+1znhfV8Zfyz1OX773TnZsAhYe3WfpXv/cu5x4l5gx2SfDHkEXFNBwNoy
KbiafKDM4nMnA/52/PayXLle+IvzNv8XOKUhj/0uCgGrD6g+eNKDF8iZrHIp
Yiq6ZyHo6mYBxZkt20JWdD4KL833+dpeP63eSRhD+OG73rzv79OzeErlNvL0
y6EYe1reLg7XrZ4hfynSTIPm2g41sEQl97LV/N3a+xBr6EZW5BKguAX0FTLK
KtuDio2bw0qtRvGT9Ofc0IrlJxW9x5z15aHOIx0UMYeGK30oA6hWkJevo7zJ
A4kDro0c7CLwOGpFL9uHav6yTQW0JQKXj+4/r3VfgGD3paPS7Povr4ImjhTO
d9b+3OBQ9HiCF63QdouoTMRe35Vb3l2NnTMmmH5j3G+XCrPOkOwu9jioJYNL
a3GXouhkixlV0p2u62YkLxGybPY6YduQwP9aGKWZJibF00cp/gF0UOMOuyyh
1eqlq+tKc9M2M+dU8gBbypoosBY/fBx+B7/g0zbHL0RDizYz6wjtjOXSfVsN
rVgCMc7ZcgXqVpDvDSoVgCWHIrw3cEd0sMOejAqOURac8b+5Y/Krk+z0Zcsh
yPAzOKwn6raUx+TOy/2g0mMsIXOs5DOE8jL6wsXD2cJp56H34o2GnrAdecq/
1nW2xoQsHLyiorP7oqebjKIhRzCyDg3om5l60KtChyaOD3Uo8R4TfLPw8el7
PCxsh/Eq1uLATq8/OeQArQN57VYpnt0EBu2ncrn61k3UhDe3Hx2OfZhrSyIj
q9e2vvBKiD2x5qNo6WNpgLFSqEelnLpfp7mRBTRVP6xxGi99pPyfnuvlOVs5
iPhXrkIddrrqGhhuyooLNUxh/mwdzMv6AXBkQdElWJRDRennB5kuRIDZsFzk
oqpvA3h+JOV6wLxIxIqnHJiK7BXr12k0SL5EitEAhBJI7zWZ3pz83zcm3U9D
6ugFUsIDu3yWII0qHwJUImk5rkvMxpE/SW0ZorBjBLTMXOQo1RcyZi0DHx6G
j2K5YcRcrw3LDIv9ZfxXDPnYce6xOUJ0PfrRZFYh3KnDEA9KNmqkqe2kiRy1
uZODpY16/+0/+Mih+C5sY9q3hTPGug4WdfLCsQANdIK+PZy6CBniczKttB73
PQLQax1Co46IfIAnt7GeXSL+lyyj3A/+1nXq05FIrPMzyv+76739CuOF97yw
6inRJ2XcaIrVFgOFhHF+1bJkIawtM6ePERyuzK9WuprBLOGbbHkJMxSISQgA
Ik/CL9nKBmmaMJFTn+iEjsWaIQ3UldiJLC6xe7+Bok2CV0bz3GzRZtgKrcHe
ysF6WUFob3tI3gfIIaDC4SAQJ2m6IZ1bffCsJbgOazjBk+Hfs1Bgy/jINXdJ
/yIl1PeSY/dD9amRigMw/N1XIyn/crteMhykN3IDNJJbNjFicn8cZhOJ1ZjW
CqKW2KI1n1osfhue87R9O5zJvAmac2MOg+/4q2BAPfySjDIntDlEeoog9X4W
kgrwePqrfW4ueu0w8X6qq3NTOpELb3CXZ5tawZdKooHD2DbNLPU734B3m2lK
RX+dIuQ0RhYyq/f4SYSGyPzLUDvUNGQazlasMVU7puAeJ9gafKBbfpVGKQAL
1hwdmXYwU+nPzxSjp3pI4Y3oHJ3S0d/Cp4KJq7IqJSUrFTPKW9rH6dIvVnbF
N4i7Lb2Xv0/y0nJFy9CVKL6HuIiXQpclJZ9akSU8rmlmUftLW7u9otSNE8mt
hkuuJrbylvPpSlU96uU7xHF/ueBXmEgJQ6vx/XBJ5uKZQ6+CRSsL6NNm2GFe
ONb5OHRxXLA6TJNc3caL+aVazyLFQyoXkr77li+ovcUPGt+0L5iuAZvX4w+9
GQsxpL7DK1bBtIx3BpUuNKXt18qceogRuEDbQ2W8/iHIPvDeYvsCf2FK9bNZ
1gOK2pzxmX/Kvo2fvJd+Vt+9WL/YQBf05k9yle4ZaFN/TIIZ+5jMWIprEt4Q
bpGpeJliWrCEcQDjMWPtT0ByTdnuAH4bQ2r8DG1I+GWfwJ6/zXF/4OZMpbox
TeFKFIG/XUx791cO8QHCg6gpIfk44F1MtSI2A4hzObrG+/V0SIXe0o9fD7oS
kyafoVEO9dzFdlb5bmv1ow67OMAFdISkVWLUpq7cALncj9WlOiZlQl5qGzTQ
tG2tYWBK1MFlDhYuoBeSHSQLtweMhSeHIivYf/l4gvNdr4YMgkqfiUaW4piZ
oVy58syYObV96L9KGeqEkwvUCC0AK7dgCRwJCjk8d+C3pKTK7+lsrhEkbP/T
SUact8zaV0JAPKEinGHYGTKtKSoKIpAaA/4lMaqPfEGUX67mjhnAyhHLbIPG
OuziU+a9Op1LhrlP7RiSqq3i/C9pbH0kw+NaU9uSRCdPbX8x7pBCkx+aIe63
2WdADKxA9XPDORCKzrSUwCdr40CnK0xx5tc0s+uI+7p6KYe3s8cV3iDadXS1
AiIkbf33/RG/R/5GBYqs4Gh+JwmWNISEDdmv9dwRh6rin6RIaJlyjxTfA+B4
+blOBc5wpaxtVvGGlfv4Pjm80RpoDfHGrpcDC7NhlEWlaaMOaMVQWrvE1O4g
ykx5iQ7VrR+H5tbFV3t/F40CBzd1qZf9eBeyLv5z474kAKAB9mepQMfgMW56
PFr0DJ4FNp7StdWhGqnO40PWS0o/qkCGKA34ZvA2cIQuguV0IU29gGjpkcAI
AakQlJo6Q3Hz7LyyOtQN/14+76R2/zQZ+BV7a1gPi6qmuS4Gm17sgFiKRomT
STKwSsk/UizGAv9OWt5Fv3y/4zB6p8Ig9x23ko/T45KeAx2Adw5cHCMqCVkd
OBTnaBOQxSAvxFkHeIxr4M3JJzGyeBD03+W3lCJlA3YA+/a+nW6cMNPRK5CE
W0Tw2voWpVeLGyuyYQcsnqPpxQnOzlov359df30aPm9exxBYYqFFRmGZqJ9n
ErGSUXJu3i8yd/bDq4XHtk2dxb49prGXlRWWsKqgb78XrO9d6su5O5MenoTs
woh5j7ptLMIQzaNAa8iTUqG7kjXf3+wPoSID/hQmelbGky/BGNTch3XQY1WQ
cyLjz2r6kOSdCzRwN7xQXlDGerzibSUinUiNl/MjYHQKhqfyaeLpgBqOIwdX
1+v4is5Q7HCe56z9g/5hytkdvJZilu6zfxvICm+Ucm++sBdeDW0VdgpRQq35
dtGQWS1S3YF42BPV3DdqN6/gBhtaI/rGMir4chxL8kuG8uHtk6LfXoi1icbh
SXfD7q6BrfgR7d7IG8a7pX2fiNIu31DJa2FZ4ZfWSy/kEtGzSi3i1iojRsQ6
mhU8g6WuxySCf5eA4JKafIPtOSCoX+4E2UjTJ72fLWOjIVMO9ZUy1zUlGl3y
Xu9A6l+yh5nkxVs/EeJQD/dEoD1sYCeTYghVZe9dh+MbWEKGoQDb57Qe48eZ
pt9G9wDYkrt6nF3u+ZrT2n6H7f9gQyU3IbYImA3FmCknoaDNiqKLLYYMtjq8
wRzKFX7Ycw7GV50sVws6bQI1FIO4x0IBX7LUUWmJkyY5wAWXrD6nZzLWjzan
i6tr2rNFg5tktsCYZSEtADsd9/OwgHAB09nxJ1z0q+l2/G4EakW86RP0VL5/
kFLIbPmwNisWvVYoH5bjqE7osS5Wf4R61AKCZk2hTIyH7HRh45pkKNzLcjbm
Jch2JoQ3TzsoZHZDelmP+HIxViL3KmXHWUG9wVxlX6AFCCaCbo9B4fx0aXER
4J5D2iwXJHiK9g08LKtH6Ftzy0+675Y210zUnXABf9GVBWdYohSQqV9I0kTy
cPsfbG/6Z/DDJwwyUUnMZykjkssDXJA7bW4168CvZLwZFV/l/NLLFk3SGQ2t
2W7ESWs714ZY55x0tZuKUEKcsfbz2UbLRHZUn0gYNG3q4A++2BmDR7nmXSnS
rqdPJxVtxy5G4Uw2CxB4kJuAzUzLu62TUuecXCQ6b17mHpy7l6jj6qAKoHZQ
4KNKFI6QydedOJcXU4BCxdQo/XvVVKLaPWo87JTWl2UyoYtnovMgCvUi8fhN
dfEHdX74OvIl/+ZNJC97yvJCiGbAXZKY83KjMirFUROyRgYcCUurgOMg0DUY
dnrIxAcpcMrMRHbpyr3Tdm+3BHqbx9qgdGAFHCAsuM3KveTROhs/uwARZw81
X20G7yaxFr+cFy2O4lF0kal3ak4hWeGES6rskeFn755XeluvmSKJXYOJYTK4
5GVFpjWxM4/iN2hpsXlwEWxXgCAq+WuVmL45LdqepIhWctc4mRveXHvWbMKU
pIqTwl8aN8R21JpCcKnX6CDl54i8LbIsKIRyyK72xlMe7rW1IsMnYTnqkUYM
D09Vco3EpyMmXzTsJ2ejmUzuRSgJyOhP8daLIxti+d+GAqc9A63KubH5y7nR
U9B7rH5OBjYHR6o1SUVj3vZmpzkN9Ks7ZFdNQQieXQsuMF78rapH72IaLjtO
o7wKnpuQlyYbfWZGELsQ37pY9qnTUZtxsLQR5qwPXvZapOWs1IbqovSDoh1E
7gcb1wnJEuEIuUmug3956Ragw5+qBScL0BCsdYgcrRHwSzrleP8G1NV0c44j
QyNrO8VqYUZsATq2XnYGswTU+ZE8rJpRlwNKVehJbLsqOh7ChHglUuOU0mOo
Tuyvc2BcTJM5Bu3eVN8qCuvjIQiORzULYihzklczsHdMA/GEnJcma8JuU4LV
uYUgR8K8J6FMgmS/cwDmWY4ouZUqe+RDISUPQS2PyVvJDqZdcAo+c5pzYbOs
mw9E4GwHCHkD8Y79TkCShV1dO8vq8YaCcn/hZiwWURpUmnR+m5XE1y02+1zT
4VGn/iy01GZ98qucvGYiYWTsokkSbNg81T9jZs2gz+rr4wkXsQ1rmNgriRfE
bS1XSG1eZdOC/wS5TSbjiZrkyojs5bJuCoHbP5MkpeHmTTNCEW96KyrxBAvl
WtiVTvSAJNZb5bEvYBTSmcWsWbgiLVvMdPCDI6DqRhVcKnAXOS1OvNKHwm0K
pq9knRDTeAQucCPssXZ3taupF7RpIgbDthCWxilYBYtIymE8uQxRUqvwbwTI
xNYx42vKYqoiBD6lwBaFdiWy3ND4pz5VNOL3QCtOQ+ICqpVasK4rh/9hiz2s
l+s7IlDFj58DILX543GtfBWcOYd3l4F9qzeE7Cj4LVn+8C3n/WcggAhKMMyq
YalzujdWJDO2ZuNBGYJ2eFmHECnHfn2osrvtDPYkQGok6mAsAbRHou/1AANI
AQisEW87BLWcSIrkyneb51JBJ8R8wahRwet3kkEn6XbP22bMo8Rk/mfLG7cx
ZBs/C47sTgAu2CReUwKnpcmwAXqogjfqTTyQEKzof0pUdU2IzzW9y/QG+Iq/
T00xSjHzonF9yJOzTZOkNb1YpD3J2GJt+1U4nI3ck6ZXLH0QAQSLPFFZt/DG
lR0LKK8Udy48XMf8QjPZSclclfEPMrIaaczAZEal6ZC4MQMvxRh/HdbMssGU
3OMHrlpFKYTHLjT/nYAoqvAHLB5vJcIR9+5psizINb9Uv8pr4d5IMnW/WCeR
wTa6N1tk03cfn3WEtdAnt1dtmMuX3X6OWv69lzHOPw1y5K/VWCWShbpDk2K/
WFRPvKkexAlaYcVEFEW/ehDdYFz/pcRO968DmuSgTpkFzmLXVvVot1cg5Emp
Lf830NCkxKVCpBbOM8Ihs7oOtqx3PkFIh/bqiSBnXvC7s9IuWxLriuIzABnO
9Gdxp+w71zGOkTKvvWev2i4NkXvyom+UQLq5qtUpwYNX0N/r6ja/dU5o2XLt
SWHHjSIsExuXsZrbvDzcYBfu0J+UrbPh+GN1fn6Rrk5MCgy8Pu+oGCHyvMr6
JuQlj1Qh8XZDHXwkvv6Zb1Q34ub3614t0izzbiFmMkhsjSaLyeB4JUPSWGYt
TvwzazmuPLy5VEgtQK4oA/C9+oOUNlhJrakUPCmRVq9Ost3dOv3H58u7+Qpu
nJJAOylIJeG+nO4TRRmLiDr+Klz/5RVfd1Tbpw9DMdjMPdJlv4oR7AWSGrCe
yCoynHO9o8tvlQNV8S+Fn2KAH9JCrfRFf2tKNQpz22yT3RwKdMFeRb+uonfr
w3beeLZBLCAeRnYN2Gs6fWUci5rj1McCWXOMJfdxwb2kb94+DzoLbwLjQ61j
qP6WLHw6T8F5I5Sb88YWXOalQ3P62AZttDNdcKhWtr3UzBjTiqt9YANoiR8a
z6k+npYq/xRalhC/CGVOH7fAUYlKh8Lvbcbm4/Vs86an7jePGOS6C2D6c5+y
bjXrFyc97c8as2Q+93ZJbbzYvp2ZuYOh0qwOMMIG2dPodsqHLDazuD8Z3egb
S6mruFwEQD5yrxe2/d9KNXZuQhs8nUpbUKOZ3gngZxR0HC6UOSUTvezcotRL
c2xP3JbTAAHkCB5xglBUdKMPGDm4Orh844AW6NpcdscjwuGxCQ0VMkzmLxKG
5925RLQAQwdWMLiD1AzF9yEKKpCZ+zA6zRRHWFxwC3TXBSCZraaMiNJ2ZknA
zGI1G4CvW/Q/Os/egGjmbhm889gBAfmy59jXmZZd4GZMQ5jJoxu918LLosKw
vXqOz64riWhaElRoqDHgGeMZB10ed+KKRhiljGgRRd84tFTLW+Fo4ru7616Z
Qaq0Osh0DKMy0L9LnVhKBUfUnfnI8Nk7gewq2rRS5oJ+1+H1WJDI0MjKYJvC
iCJhe355uhkjU1YoFrNGEz4JPjzAm4QBaoXNU4nJDUJZjl52AwQDRC5X/GIP
ts1drBqSmhUWCnLBgWuhiAGB/uy0GQa5u72E/8JyLnKS4db+Efdkl/aaTVhE
kRAJmuD/BMzcKDhAuecI52MjfIanY9GAqxiRDlxG+oENsp9H+ub2Gs016aTz
tjZoVfDHHdnU+2LEnuk5mzicx6UkV2ymW1FUmzyzu3zXYAKWjC5aSpXAp8ZM
7AuVL7Z1tYMd1P2hbX3aKQSjBCETiAowMXbFE00hdeZq8kdMAAw4dVFG8LhE
YcCAthguHBXsHO8hh0wAygSEhgMO8AjePHDveMfeTJXqx3z9sARe9a7ZgD8C
/d0FFn2Bb2WJ+dnwB1cT+S9Kf+N/GwC0+pFxJYkBJQX+NNM0twLy1uhZoavH
skaEjrfRW/hmYAuFwsapSj8zH36XJZU6WbzspNEBn/WZbd6n5ZKPedFdqAQf
pXQQOVbuCH5xAfwkocFb2OOZdJUI10laI/tyCZUWTje8PUmLMJOAe1KTyCHi
wk7n08vYc94iGZ/5O4+LsK0+PEc39zBNghvFkH0ttoztR2UDkAww5Xr5ei1b
csUOr3luNMNVKo9w/3Lor0jiOIAdlN+lLP4aJ1+ATkow6nM0hLtjqY8eF1W+
hRZSeNEWA3agUOEffTviuTcTwZ27E73IlSU6qWMzJWepsScz6NNqUJtIB5wC
lHdzhl8Z7vF77bx9G+d+EJyrozeUuADnNf+fwRzWzzUqi5HFfWdxS1Rxycnk
abXJkJhQi+9alvez1Hjb+ziw9hdbFnhu1g3gPO6qJ6/zuFON1wCxNej85GXt
G2k+6b6icFA6Lp2GA17aKRL+6G2ZsPiJXNxsR5e/Y2fe89/LMWWtzazoaDU9
nIjGf52c049hSnkLfq7/lSFicMtkAr80n+ez1XETKJESvCXpa7K+30k5l+MM
BJaogx/QtpBUsxP4gT/+CpFu3RB9n/V4OXP4YOQU9Ki/Fz2N6cXuxg5uHY8s
SYGOWFtaIlgTYG/dX/YvkRwRMK7KrCWzRas1NGi6BHlfE/8RXsbOqX8L2hxM
jFI3qkF1ZUT3JGIY8e0y1EU44AtfbOlN0wiZJiBUU9FN8qqkz+TuamiNQmj6
4guExWUyXaJXZpqtCikaxGNMKmZLVUNa9+ag2VLLsVCURC8008WtTyxhtsbq
rZKo0w8Pop/YuicbPCPJPEX84nbTpJ0mmnDVe2u9ZM5/+j7EBOZJufxjC7nE
3Cqm9PrUBQUzHw3PG8dvXDiNeLE8+eQpcipa+E+GRVk/WtsB7Za32tO5WcQl
RLeD+ebWaPmNTPc+GhlR4ELZp/rSIL/wZOlzvwjZOmyP7NGqE9VVzb6BtXmu
qs1x+HgOzmkKNqq8iKxxO0Ah3XGpOOnid+VNnoezkEI6p/aPy57ZW0o7Tnat
sBQ++GvtVgT5+KsEkApnFFzcQ+9V30toK4vmD004JYRrwPCwedydngdnRAtH
alsx/2ssVjDAtuCmr5yXMzzB2t8e2cd8eAcu4K4rh4YJQULsuOXnmrqv5IRv
6B9QDZE2a+XZzMn9XE7X2nsbDIc3I+epNxFKpiUZ5/wZoEjzLXh4NuK5ayng
l6r3nxXviWbViykqldRsc1D+J2Zttx3jUfTKZuEEze+prAFctuYDpEBFk5uM
ooAUDdUD6u/Rg/27G5WxGgG0pCsSQoTh1ChurkiW6I15QT49hyvqfdRddyBb
y2IRMKIRmcLeJ0CBA182RvetMBKfCi/xabU/euGmUMxGwJ61lP7hYqxEakCu
ly7Z6qb6oRz66jzz4ynkTLl2OoLZF/SNmSO0XAY5w2+kfpR9jAZi17skKOkj
gwol4WoA/4Wj54HQI+W5HGoZ09CSdGTJWlFvU+xesfQm4kiZbaoMQczWWT+L
ko1SP3J8LV56d2EU4TPDXSi8lpIwFNyXuPgi3vfxWAxCb/KlVcAuftTK1HLw
yASgX+K49Pu7hmn3PTv0KlcpdMWFodRlwI/0JBMdUWkO4YvNDF2gsCtPX1Ma
cG4O+GX6VzpScpj4ANl2d68D31MmcdZWko2LzW6/CqtIM4O9lZivVtKQXG13
GeOKNoerx0oANRAHrQz8deZRVjIBgT1A2V9thH6vcWFF93GlRrQOZH1bP8DS
Xdi3Bx3Gt5KxKKTM8FcL6n4+vwUc4wkT5KiVg01ITWmikcwexf+ea8Vw9spv
6zVOvMK7pqTrjpT3hNrJWgC8MZgRXwARgV/Vx+WhwG5l2jyi1nqkUgshM+gd
fB2dtIUtI5K8Qi6UwG8ZtAEqAPAiDKLTKaSjulFgXOL21+/oBR/EWAUaF4qB
O++serQoOZg7ENzWkAsGW9DdadC++5e8MliflCgnis9aJpjBbGBYTFEHrW2s
L0nm7jv2NVrDjukBGS+EJ6znJ3QgOcsgbXOHT33Pu8AQbFEsl1b7NScWyvWO
QS0HH+NMfzSax0tIs9rH+0ZS8IkUZW7uSDz0nIHzytUajhBS/w3CNGFVCMdF
ZkWKAx2laSKv/zNi14g8LZe2urOC2vJ/AtN/YK/J8yWspkdvKbsv7cwZ+BPS
7TYgESeIgq+2dE2QgWpI+Q2zJfzfFkNsFo4Ovpp+lIvWVWBYSEm5/TeiQ/Z0
a8W9CtEWy+odS21fUf1+T6vhPqJeUIa+jqkbyFQSotw4VY4mHSW/OIawKSWl
Q1qZszTdhyt7/M00M1AR2DXlFPADL/zTi4fuG6T5IYXhX81gCOHLd9woGuBr
sAgf3nHSlWMGOQWf2ZJ2Xa2kT+4sa0px5juCjHe/3aGJre84b0cKXaLJwvx5
uN6W5nGv+6/xkaTzJA2SN2jmPpb2mUsb1prsWJAhZIOPzKL08zwcFGcUi+t0
bnxKMu8ku3NfXuht6TLTWm7uEFlt6vgNsTh+NjLSd8+ghsCjaT/6AXpoT1rK
13gtuqOmCUT4ftbXFkhJnIn18d8rlgxWvEZv9cAClop9jnT6hPeOea2NNRUe
aFLK4Iy9y01WhFBRLaeiAAeePYEJbfDDQWh60iJmJTrCb6bnlZdrzNNbqdD0
nDOf3ro1fbXfvMlkJHBOJj49xVz1fx/FirPghdZGytblWK+myVDEf3fuKWSU
kqLXKDgMt/dIAMeMSGzFEvSkdKNZ0DzCc6X+GpCfy7CiV8Jh2IP7W2CytXxu
i0e80FVtL3reIgW0nPJ7THVP/gWEiKL6LgrJQEJUjV3mFZvzTgXKoaMcyjy5
u+h6elAeisPSgsnjPpi3grB/7Tc6u78spoapepPrvKgcQC4JIbUtbW+ZXcS5
QgwV3CdJfthjHCUfuZSwSwstBSOOKoIgHcPZbGb+2vHT8yyebLsxI3vuB85F
j97wYLsmNS8hyhRusuhFjgKCbGmdLvuVVupxFIcFkQgEWokEU3gCFfigX3tG
fJBk8r8k5QCi5BSsr/o80OKD7VG4OTw5ep4N0/uwb5mR3m6bKEYoRataTs1C
qe1Vzttz4wUPohMLMNMIj97hPuMDDLZTxfHxmndTH4rcejOXQdJmiuAd4Hmx
KU5NSkvyE8Fqh8d/435gJifGTuwa12bxXiddafKY/2fLLVDatg7O6nGnsVSO
1KIVr74pGWZN1KdqYAfmKXddA9lT1/IuVTqaOdn51GKNzO/P8lDyfO5DWyHG
knNbxT7S+sh+AzkyhWq7Qzxr4zk6We2HdevVT2paO0IpFWEy341LU8wOPQNG
dm2RnUqpREeTxyDJ1/pli6iAjcnKxpfxR0ok3ZP9Zauj725WECFLkNnuwBPG
BYgwScIjpLKG1Pd8JnH5MY4tPQvER9DP7jUz4CzhdvXhK3TBILeb5BcbcJnG
4YRFG2+5C49g/sctbWOft3J1V+XfHgKMzFbivOYfFBHj/UfGdc+97M2To++i
lDqOZKnNX2mR7zOm1I7py5cd0MJcTZFrmZVA+QNrVc/s5iwXjUVE/ZVddoVM
XtJ/14T4ybM9L8r8BXUyl6597XQPsjUvFREQGYW7gnr5KGs7I/TY/a/UBdOY
xZo9omefyaaNCuk/UnW/9b5KDoMM49MJ0pBjJFhE6EfJSLCQsk0H6gQNJSj7
OXI76qeLaulf/tLTd2xBfckydU7uxLd06SvFmiDvopksaOCR08eDY/e4Rh89
cYPbVSSL4XSyb9UsbM3BONDpKndK7bsjW7PRIg3wvJu6/Fi2sO38Z8Qa4Ydl
mOIkFXRTEqC+vNHnzbN6WDVOyR7YeKPOSC+ZvRD8X52jRxv++MVZCmkBdZO4
0AqXhUnPDxggcXJ20EceicmYUjWmnHHNoQOlCsUiad6c2cxeSQ1nXEyPD/El
u/547Jr7RpiBqdfTX5msU9WhH5STT3KJqai6qYgyJixJFvBYpk0eum0ovVWR
Mi17IiGU2VqMvn/oQDx92awaiMWQJXPU4wTou3YtHMHXVaGkNgtLT978XrXh
8vceKv2iRL3z7B3/zisZGlwt554mj4EzHPb/R02NZu9hfLJ50wxBMoEnqUIQ
4qaaE6frZ9M9E4fLXVaAaftv6x7kLjHvAptQ6QssfxgZiNw1YNoZ4qHjXE5z
RjCliWpsTxjSdVpR2VMWiXfSVC7higiScZkSVJQWK8e5dLfTkVohs3lXhfau
bpEkRNll3ChNGG5TywhCYfgPKVjUO2mdCLJZU3G2ij6YIKU6OTYZzPVeUho3
AoRrAQJcx8y29GPhaPS6x6AuQKwLWwX1QBTLV/RKhBKzcmg7DZ/4G3X4lYm0
gE/uzrK0AFVax5HwwaP5jd86gf0rC1qnYkbMgqJBI/45WmYaV7Ha8637kHZF
Thqr+ibfYv4zmH9eAPtqZU6d8MQisy5D1dh46bTqIZBaHZQbXLsBYtuOFiNM
bVQJWd/Hliw5kKV4HRgbsX5cEoK0vCszoNd9Ean3l7/mlhj6P+pbkmQm5rEx
Y2EnOeRDzU5o/CYHIfN2b+bW3BebpiPw2L40z2JMzA0HKJ9skh7ZKGMwoAgo
25NRfnz4fDBZ+FjQ0bvfvhaTaBXrHWNjxbqbzqDTvvvHfYZSJs7bNQXsr/5n
4xyUii3m33JnfRLlCpFslvhHPsEI5G7nh49FLIdEWlrVpK2o9N2gIWD6qN4P
OrTT9SxJ51ibv5tLWgaAqcDPvn5HxBinWZsIWfmljmvuWw8ttJmp1npZSwKJ
Not1Jivbr33SB6cayo3DzWX1Bfdzr2jGomn5NAqUbXyrotHETzPmFkKA8GPQ
M22X9s/vlo6Y0U8sLJpa90/WqEIxTe+NyIsR3NDQANl8NJiXYMwThSg7T7Nx
KypCwUb9E9jxtGthlu+N5M9hiD3tDOVzwtwyjPUiEopTM5zGTLHUZbTLDQUD
VqK80iJ4hX6+JN51OC6A6dzu+mDsLs4dUqQOa72i1NEU7cK+3lUV8jm7VVt1
nYdm4s96HCMcLzwF0uYSbLTiMb0wG+DRBZO56DNIeou5l3+AX52j3eKeUlNM
5NEZWFwZ4gSgZbNGW8oS5hDvy65jVsUTLdP0wlZNO5twn2vthY44YSSj6muH
mptoM2bIUmJ4jYpo56U7t3yrz7IlUhTgUFKaUdqBFaQ+uiYFyl3Inv6S6UM7
teZMBw5Eu2p/8Yz+GYAefiuRFCDRSyf/H4a50KEJH44FsFh/j24MTf5/rQjB
Don8knKQyJXQf1HBJXEkMoUUSx5YAGUnt3dE0+1bfuUgbJot8Vv9OozN0NUQ
uz40aOQuWV5XToGIbZ3xnR4g/EtOANEQl/YOLCdw7+UySoZxYfqiyDd8UlOf
AtOiFjSyryhIuFjShBTVg1GdeEI2IvwAV5fWVCx3nyiFoE0vHLNQ52ITprTJ
htH/Yux11wMDm1DsivVO786OVyMwC4MkV0exq4DYJXNE+J1lhmEjNRCIZjRI
zRbB8AJ/4KWhLAAQAfs94nOu4O/UoSJ3HVo3VThvUJraP45GHZe4W9eB2Hnh
z9rS1Okcuiv/Q/GQb+yW79mBFddRmAOXSH+DM37WEHIKFz+vTrRtDEq3jRoZ
1FuxFUqUOA9WaNFLaugD8GD//Gb69IFTf3jgnAQjCUInB3QQ0P3/X5qYX94t
vItS1GtKPZA/pOU9Cs3nStQvYuQDrEcX+F786bsIdSv+oXn0MuGpnl5DBAgk
zEI/ckWz+odnh6ul65jzvdjOjQ/AHg8XCbg0VI5KzNAq8jvzfl3VSHcd9PkZ
YVJr44zkdg5rTb+C+2oSjndt6tRUZ3qth0z+JWv28fLDsc8i7VpwWuDteB91
ROYBsTyb+ZRu0pk6emPq7WQO/VE46CPaUTWjIUg5EIwZl03vC/moW6/Ryjo4
aMcdjnpAbbhpZkLdu8h3n/4aG8dJmG+5EBCSAZM591GcgmhtDPI0kFbTlTmL
k8Nfgw7uRroNB3gr+2sdSuZY2maAtyukqig54vqBjI7l+HyZB/ZEekXI1QBn
YR61iYClsblCWDKpqvUJtzLE7WXp4zfEtB692yZjgUwcYKxgVxTAkXbQi2Be
rp3bbL7J3EaHdD51w3La6ZPprV+C5ipGY3R1mLwTAw7nsJAdbGZn+ANCsFrV
cdP0s7rAXqj/7eJCtWLcLmndS3YW+zBVkJUWbu9liEcJ2wXyEgKGmlXfbrca
qjJ9Due+o/bH9+9DZu9wQ1RJCqeMuyZEeVbS5UNOvov1+C2coOBuO4s67wq7
nbcBfdjkq2yDreC/LcNAA39zHXE9+eVkl98HvlZ8qy7iYKahKv2fO9Gm4RMm
uNFrSG137lNtvenzNKRJr3KYXapUvgkI9qFxCniXHpYHJ6xgtKlROS0AAHyJ
3JBAOLA0xiVqG0fyU4mSFQzRVCA+BhEszvAECdueti/qGy0CiPB+k5888hbt
M8JBN+g008EJpORnwz+tZmAHo7lRs00ZGvTg61RJDy1H3J4uuU6GchX8Y4UC
csOqyJJIsKezICVOHjVY1xnHbJzTkHdhgXcV5E5J6mcPumUp42Pa5XuY7lEZ
KnbZDLfNzPLLYPUuRdpItJXQ7DgSAlVPjXGysW5kEMGmQH5f83iGmD9tjJUe
LmyV7rvJ26RAmaH8x0QsoCgjCil6Xtt/QnMsCNPTjPOzx+miYF7Z15HhM4aB
fJShnZBWyx+7EyornWF0iqKbIJq+WHotGqRlPt5SNo/Bx3tpkqH/A7o/PCez
wrzA6Wc0d2Tq9Mz40fEY+ciofYhXz05eWCYZQETR90C+U6c0KC8lv1Det1vd
U6d4QYDdI7t0Kn7evKZrVaJONHu+C7NKffOmImEhjMZcFrxDQL+RUw6YBYhL
uK6W8GeDp6TWbPVVJjr2FIShXOtz90ztXEOE0hqzoV1dzaQB6gn0bkDyvLSr
4kzIcrtbcQFu8u4FzDvaj/GYBThqr5CKvrhJjydBfVpFwIv6bS6zTWNpA3Mw
bjl6irKDa+UZ6B15s2Gf4IPPNzaHiTHL/DhdIWxYoa71AhDBtgmIl72dxLHE
p13GVTTv6kT1knA/yAtSGwA1nUbmuHi4FLPlUg+ZEk3NOqZHpHvYgWdEGvam
Gtah2MlxjfUvYXVYpzbN30BmpRti9HLvdQuVnmSb7RMXg+/dlFBpGal90q/B
AtBN19RgfVXAZhWhmcQQSrU2WWNMhFsSB2QPBti6glOunddCENTF194Ar7gD
1AgqV4A+yhshHlKmbFibsH2RmegB87A+5XzFSRD4Xmy72/Bu4yNEVMEBqYGW
31WFyFdWy6pUIkzcOTZ7SbwtKzmfBHa7TH3AAQo3vgfbI5BrF6f0ABle2Lsh
HHk/ui6xzCXHEhg8sMtXXCucwRwFfvoZfkEMxLAhkc7ZaoTMZccKL5UCK+of
Q/ehdS2pQw+X/I/cq3co5NHgHnLq7LclNJbKE3YEgCUHYlEV7IEss4ZnMVpq
EQc7m9fU+6TzeZOSBVPNltfcdnoD/wYyAMXWle2djycq7mfde4wHI2Pj54O4
+DPJwj5jTaJO7xDUkEkhc2Z2U47616O3+9YmQdI9r/fXb1QZA3SPZ3+sh2q3
IfGIY0CufuvCvjgeKEResjT6+1x+bSQdKQrTFwRAIXjcllHRpurHANZEwWDa
d+o43gn1uRWXxD7WASv7sNX1vcACFybhMnHxa9IntJReM5wPp226K/WKi6Cq
0epQjAGW2RjB0Dw29ysv9dpmau8p5kmpaowgERL9AeO/O/sO6nFpyJFuiZ9H
xsp5UTCvJGHWeQMutbLuB8Bu6zewzyaTHaeXbgPuXjIldmmlG+E4z/aRp/QB
40YvGVHqeD4EzkZF4iQ/7HQ9XO3D5WMZrDgiRDKIh071z709XHa2nWt55kqL
H7SfYjauwb2H+qBiC7EYiNoii9dkyYmghuMYaBjWpGBGexGPrldejpugtnLX
P5I4naBXkriYJisD+5inZMFzvYc+4tCff1BVRaxfu7WP3sZ/efz5I+gFhvzZ
eQMiIYK10obb2cehaqPxnmNOwGCiz6bpUEJpvPxoIfbIByN7NVUJPHQ7LmLQ
umneW8Z8jgiHLzBFm4YfRe0R/Un7+zOpNxdUkPxLzyUrWIn377qYSjWkMK75
w8syCoP5DKvaJ7Jzxl0dOnSXC0V7+KOXCwHCRBCbr0AMXBI7VqSfacGgAL82
DP+WegufbT7wqKXhDPK8B+zMLg3A/j44/Qv3Cxm8HBC0qRSzEn4W1v2amPr/
+Bat5kXBpQ0ypur8JMTAAJ/IAXRJlX00/KWbou1uocW8P33Vp+P69brloq9t
bo8iMKy5Lv9jW4u/qkLpg9J03M4bQ6EszOake34X5CNN0X+LJVpypKp/1I12
Kb5yOCIMnLAfy6nBgx0YctTOT0vVX/Z9HTVz8d0SdAKqTz+8Oaa1/OESi4Ga
loS54Zl7VAynTj3kXexbcSeAWgFogXyogIkdeNaLsUN6whEs/IbbwwnRe67+
+fvlRCDngwnR93Uumpfa4S4+uGdd3WTqul0EYHPw6WJR8M0r7mIIFA33pqt6
M/sObEKsLfu24dAHGdI8mmUsjHJFgMQASpB0EcaV0wbLoKpFlgSNUA3YMIcA
NHcataSRxhS2gFLrsvbaWo592BxO1RWkN7gI5jcb1jU6zgTH9XD6oFAI5YMa
LdcRBEOIkTv7241wteWEQmAqGfdjjgFrHlOYPeslZ4v0/HPSqRfmgpty10ut
tS2rSJbz5mbPNXunbvVbTFPvPnZEy0s49l9Jv8qrBWfjWqC7AAbh8XJiDbJZ
EsTHo4Am1/yNicQlgwQ8rR8uMdCg78NoqVrhpmc1nvM75Boz3kXoxEkQX2X1
7/+K3ajTnvqrQKBHoMav6DzWSv6qVQJ2Wr4pBlaBxmMxQarssRmk7pur8wTV
S52DOd2aQX8KBHyoFh//354WtHqimuATYUCuolfzIJtf1QK20lzFEmtNa0kZ
RI8GkMbrO+sf71JCh2Bfh4blIGvi45ETmw7VrDeOyJQPjHjW4OX+zJYGLQmm
mbr15/YPe+WhbvVEL1KD5auvJx3hHdDbVg7sWD3VroCJpufsc4LDXDb7a78V
Orj+amATPQrgpFqACieQZgmCU1l6NlvyWIGOFFKjDVw5pp2bo1N/zYXkbL1z
iOU051lHGlHrN+UtVh3LqRnkzk9gS+6eVdDosWml1xZ9kg6X8r4FtBezkfr0
SFWypKrTRv+zrPMBLTttGBt47n1B2wlg30QILZVyzKk2Ype07Mik73CZaGHY
z/UeXvY97BUXGSd7L1w25sxN/3Ny+6nR71TF5n0K7Yf1NV49tOpoqb57cgJS
nHvvhzWP6VCoRNOyAPMJGwdRNS4/JexLzjStwCHxqAiMiHm1gmKX5yEek8H8
wP5DAhyW11h2whzadWTH1rOgUNPNyHAKJnEw7rKc6lt6hmgjS6j4C/CS6A4F
XlkF7+BLraoB/QFMT5lDuH3SHgdzYK9Jc5PD2/d8h/AUT5PVVGCvAeO7SUac
/CvvEr48/P13rVkEAiEeJfBMckZQRFKZumLoSOJZcwYL29LHbKNqSU8+osK6
7miRq4p7mdjsSiHKDmojBFDjHS+3pVJP0LOfdYj+vB8p05Nt7LZcu3cAJMOr
CRmtLBHHmGODP7EqQgLAq6nCkhoWazuzzpVtofDAeN6auqjlV92A1J9k6ACH
jK2Ufd4IvEFtoHWsfgdOuxE9GRcaCLdK2myrFiXuNek7R3L4iuFe7OQTbN77
rm5b/d4WQ/hK0IIzj1D12yvBDqSv9xsIUjxmSn+5GtGiwLm4vhSAAadsG5TH
B/bT76uawnmxR23gM55a90r4r4RhzJ4Uox5M4hq5o+b17TblWvFpE1ERP7fD
AQB6NPxIIkmco+HdwC6OlPIAeQAL2P3kEp1WKT+YBrLfhEoNVVVMVgf6EXX+
IZoJJIOaO2ZHhDPVIlw7Y3XATTeDrwKMHMH8YiM0dMDsHKi1Q5PN/gHHYM5Y
hcFQVF+8iPLYvJb2MwzX1yl5pV/XZRNWhO+lpNKDr70ciTa3Bw829IFkPBez
dfXLp6Vs+vi2ohm/ydG6Ar+Oe8FId3OrTkQGW8bJg3j/aWsh6tFDJas02v4u
QXCpq0hELGTzJsvqRMo2/qeNxLg2To39eL3mHBjeXS+uIbj9gd3/Ab19wNq4
TTJpvSRGk1EayibrMjq49uglGNvtF+N80C7UNVwVlSGbjU75xlzHhpGR7Mip
BEMd4dp/fZHW4l/+fcrdp9pPqOZfEEQ/bysVirw5j0AV7HzSMURRarSqAtPe
mlMexkQT+0xISwr9P35f5lFVshehTqcoMdWWXlpotqAngUef9W17W9k8QzYN
ufWssgb07jfnTzX8Qs3aSXbDhogd/8EICpW6TDCwotuxq5ByFPs1Ph7IsIvJ
Tevg/moxx/oa3Rrkd7EVc8Wzd5bcI0eOXZVGdJOQMOgyeSX2FN18LHXdbCo7
/U/+/HnJHjJfsi/RAce6YxgY+SSSQq3pX3XxMm0lrnK51/Nx8+BMjEve3EU/
/l2hr8RY6MmbYg/lIFnJUcwiM1n62RbyFs81R+tvIruuH/b80jHr5Z9Xl8r5
PQMwNjsnzzkgfkt0t2/2QbzyZEleUQbBxJZPDf2GRmHL0svJG2F6QAWRmRWy
h7gGMPilM3ZLNMZpyjtPufc6XzOjm9jyJ4fY+wR0rPIfianmMdCO4Fz/l/dy
o9RMndeqJ48xAD12Maa5u3NG7nTHsA3WMK1HSqL8EFuceGZPDNgzJRaWSC9b
QRgfHRCsZxhtYGqdQ4Dak5AIkAjyoHZUpay4lgYocdKdFzGVebvyTKPpHb1B
2V20EvP6RbrkJ0Dk/TC5FzO7Z3vW5DE2cglheXdVLLwnjamAijt0KM+5DT1m
gMELNk3tREnejdMlIYbKX83qQksN9eF6cxXxnZMmFlEGgWsd4JzHgmAC0cQx
/KqKOTqRRrvm1MNVc9N2GLxxL38n2j8Iqg73KqBXWxzDddRl3WReQn23dzU2
4TpMm9a2quBUDuBBiy9eTmLcfYQNZLgGArL9HtRkk/9chOE85Z3T136QCu0e
NwfzHiCCFlKaDKYleTO3j7OMWilHGBN6zsyhPl+KQyXpC8NTRXNGobuUh2W2
IM8U1ZtrUW7gChYsb3KSP2uAy/VgRi/SDOkYeUJLkwLhCOA2Ki5I2uzPh/F6
GLMPXhWQ+6ovAusg8NU0xrV95xcNsVkdmPuV13mV6SACvhGrAG5re6dtdlpY
ehNVHGrjfE9WqOTrbHqCsThuiRLtmvuYXfXqH/gkln29j1pF6Nj94VS0KwG/
/2IcCzNYKEcCL938Z6cNGoKl/RWOs9aVG1qjUIgF+usYtPkKCPrLaNxePXb+
RgzRIE7JOeV+Qyh4pmkcVKbmePI6uo+BEWYTR35nLiQkBUsV28PqB2NFXcey
+fIuumgyxqzOClAI6ADzWqRloCVZ+6l6jluh0s5dI83py9qkhw9aZMLeZAd2
6e2m3sIgIC5rAeCXXccm3hSu0M2ITXuJwxd0Zw9szh2y9rJ0uEFBMBQ/SZmW
qHPWDjtWE8MJZVcZgdEqx5HLt6F6CWKfMBlM93wxRnSkT3YLNtjqlYOLJrGy
tYITI1gAGy7EiLT1TN7pvtBep0abVeljlcuzr5MCcCVCp3eSpERsbVbyI8vu
PzN+nAoIitlxhqo5xkitpDxSx0cNUxB9D52fXlVHr3HmeNY/pRGiRiqMepFL
6X8rYeDeRFv+U4LiD7yUZbUWlnfJN+5YorZ6zrvkn+haIyO8OxQQl3LmBBff
hNcTEbJtabDS+JDI6bJiMikT1oClTdVCspDxaVOBHvJD7nfuLrVl0rRad7/L
Koyh7Df42w24kzGAk6GgpZlf8qrh6qnhyVtPF/fll+CWw7RzH1j6Qv5UT4yr
zwjDjjcqI4SCTliOhUn9OkDisIHPiJqUVSFiC7RPusb7TewYAqM3VvsAPBoS
zSCGzqxzZJoBgBT6ioofP+56W/XrPggvu7u6vyOC5Irgl7npSa3sbIh9UpwS
JTSjbyw6POfXyWSP20n/aCEwqoAfSaLP4/pxxaiztZMrrVZJ0U6qFAib8V4F
AIFQeC9ef859zt5trAomt6bGuNxpLXSmHwfQxGumTxcx3VAxGE1isZ6TN70X
b7LJmREd7S+QN4qc1Q5PSHLfV4n9qSaRTPIHHcv2J4FglqiDCL4dl1Z7rRIf
HjkYSbYc7o8Ypj+N1Fafq2dkJqmvnnsqdY83x0F63ZQJEQTjtMB7ZQWGoMT1
zBJTPVUtjcmHpwMarjRGQjx71CGqrhl5LdnKDQ40ndKGst3stJ92FSolUpV6
tIfxSq7cJjMmwvb6AJLpXScoQqnqNtk9s4df7ZiFv2HAzCw2v9n6AnmOXe7z
LLmKQ3mJS2AALICoxrn59RF6FA6n3tAYHVhx/NeeAVQ5Qay5vcAjjMgW79ua
A4q5bNlF4gyIdiJQDvupiE80UhpY3K99G8pHjsr4SnvBcOGPAfhifjDIaSye
IjBzof2QnP0qLqfsIC7ZNdSVIR0zErfBXZk+wA3T30SL2rJa3l90bHbVgKNm
EjQDmbDGiMjwYNgphq7ZgoOQVTgZ7S7YUSi0s5ZhyCu2heNTU5M4MromZ48f
uzEsZRTDGs1vyfY2wcoU3cHALPt7s1NyQsGu0QOyp+M7BqVVDcvnEM0p2x4y
39/xMJpRrV98kRZ9i/l9QdfL8ZbWJESV3t4CVczVQNOnDvMallOWzmsK9lZx
LV9AAYCwmFCjrk4NbYSnTfNNeHQyv3qKhFG3U43eBJ7Vp1vw+bLp3wAFnFgR
nKceJ92Ps6HHR/l5sOmk/QwsbdGYZPj635wmNFO32SPPRmumjfGwq5V2Emtc
RGB/ED3eaYQDPtlxmXxI7HorRd0A41xAlBR6M37jKv3Oz4wPYDH0lQa/0RGN
gbk0+G8sZvsSwOCgVHluQvhWESwuLUqPL0+DT8gcFRn4rY+39rh6Bk39a1uK
eaymraDUtulwV4zklQ8CGce0jo1bdXy3CM+NeT8kenuJ7ENgqRJ7JCDbp106
cU+fGcyq+KdiieR4yiw+LVDrxmynmEy8u022UbVAka4skXeDUXy3wNdF5Oqw
oR5zaS/obrrQxs8nwZawxGEE16SXX1ftzqTq8w1ygCdjtObG9cZSCAFwLJFp
f34vs55RgWoc/qOvLUfCrLUOTJwQWrfNsLNSNX/+UlAc1rfcHglQ4x9egPoT
kP9in40iKu0kA+Xj6h6c7fbyswVHCVBcwYgOqcvBlWs3s8ojtlQk2OOj0AJ7
QMKogMfGaIYmsgOuQ+p1vTMFBu41eIuNDUCs8c3tYT3k6jqURX9zcw6MlMML
ndybrEl2N1jza37pYV+NVHhxXVeWDtthGV942PalXY1opAE5zLwBSmvF8vBg
b7PpVB8OKXy/L5ISIr5ilWcM6jEeZAAVmGsvFpRO03U6kP9fA5OqS3WQquAh
wGT0Kn12wAV4u4hTptc/BFLKAkKQruNADa8MvSg2SX94eGaykBX3OIKHqqXQ
jdvNszS5P1Qz+SyItdMG/FyQjl8dHifaK99h4zNn4qCwQT9heGuL4/tDo2Py
EpgjZVxQLxxx4pNoOQN5fP+CjJQ7SLDF9cDRYH5fw8ZirKHBWkDIEriKiRJm
My/ffOgpvx2X+dF5sRtO1+EcFoFVXrbxwTY4D7d0KgaSDAHGEoDgwDBUIqow
Bg1u02Sx4qu5/u9WCwcrQRdeZuXmua2m2e3rgpr/Ec5nbYppeYQByV068GBN
9kkCftQxsZJi0sW0/U+JdZSvX1jFf5cjz+np/QF2QqigEZvrgiMCNxdkGpG6
EgbxQKYtz93coorJg2uuCoAVokhBek0dDNiCQd+aqL8O/MCuxqkPxKo/BcJ+
lSXDnS2tL1ai8KL6lllNy4uF2WLqaTNXnzs9F8CsjRhXwROphYygKmqKVCCz
HcuAiQ6OQh4m/zMsqeC1Tg3hxTb75QfL/EVXh/gTf6JQ51rWTrBeJkuAE8Va
Gj/PfuAIYlhAGnjEXP53EH81WTN+EfN06HxkkypT86DUbhiFfdu/EPeQ4iUo
PqfBHRWdAsb6a3/13DCq5UVwoUtKGOrQnEbI9xDckWguu32Q0ePhf2LMcHSg
QZbg+x2WKoZCqmyR2pcyL9xMa1h+kLZjSrPYX6mamytv7KSAVZVil54YYzvp
nOTB1qj77FuxnFP9gqsB/7NCEorrE3/tcoe2p30rHV1V65wGlmqJAyAGbrRO
2AMX9WBSnJkxhCoQXU43T6w++u8xAUzQ/6nCkggDTyFqMMUTBVtqU35s8quQ
G+oEcHnXrtT4e5ubn+SL7bZSH6gGwyrFjYOskSK3oQs4rK7pBGRFIJ+P0ns8
LV/W2zLkZksvWAzzLvIGsUzoImGU35GvaB9tERLQpj3uKANkxlSnGxug286j
BpiPMUmj4EaqzpH95LjXkpQbsTjWl0jkWcK2oy0AHnGkTbsOYWY4ln997hc6
c19cU13jiDwxFIxrVIsDk8kWt5qMvWu5pyeZPAdjd8KDKV1i6c6xCMAZs2F0
3PLfBvDeQE6MwLWy9xBLJSPazrfSY82ev6CbZcafIPppVtblpabiQWPs6Sqq
5jaJ3xoyxiPlRCR/LhFO4vRi7pRgr5qR0X52M9r95VOcoQ+RtNJV1RUYrzhY
XfEknEEiR1v352ESYhJMjblRbBDM71eRqcnLvK9RoDBEUG2YiX5iiNsX4ZTj
W72srg8ywRLuAT85bbxBJw/VnT2fypC/Msp6+YOTWG0KLU+wA8OdlECzlI5b
GgbEooGQjewnmCrAehRP7xhSuS3CErj+qOLbRzK+Shd4lXKiIRKrZsG/yCWq
J5I+TtkrV3Tg6XlWOgkfwaSokHUW+xXemgICaexRRYLZc+RH+LjfRKNL4fRJ
VCjoB9gHryPfdpeF4z8q06yko5Oxu7hDoWRIuvEBbLFg2zU4sOerDcz1lEKw
m/JLm2T+bWQH9q9a8dSi35mRccDHgV9BkAde/Y2Xx71/71q6LhYgeDqMom4d
2drSIHqA+8pwKkpBt0CT5OXwgOIwrkZZD3bHmJpDMCWK07BAiMjKKBsdiaoO
bp05nDRp39f+6yrtabJsSElk9vL5vxKGuHBZNDmtqDYr+xPscUEkJbnKynnw
AjX8pVjtkJJbNlp9ZjCtRK3as5IQF8G6eqoFRW14k39hQ1479L9eW6p/xTnJ
LuIZsO8HDUfqZm7QYIse/09SQplurst0Cr2qVa14dAU8fTJTbw/vfG4/vBrD
RHm+9Cqbc76ytiag2AnY4YRcV5uqIL7x6a3YEvdTbya5cOQ0MpUjxBBJhEt6
T+kKD78b83HPheI3SqrNAovnvg1Qw5D+H2ywmHyovFu1XJS8ywE4EnOQ2Xi3
nq9jf+tQzuAwQJCaD0ApdxJbXaINwzianMs7cuH7edz4KGXXsIKsCc46lXSd
Jr/engV8SAtkVA0coICkacaMGjDB0ZOexzyXp+DwF0TlXFAbtIxOyQnjAzie
XOhGm5ssJSHm2yGVkoMFgRR9xqiFeqLN+8Q7nlObkQFYiF87lBaWTvHMis9T
rmL75ILb2oyKI/ivcyHrc/sZ+l1ZIHyKNhYrSdj9EnMblxBYiQCgZ/MfiXHT
qpaV7ookiclMgi3SJTssQQDV0vHuQ1pzAB2n+tp3i0C/E6/eMiu6dvvG0pCJ
mkUvu0lqTlx4Vh+tIdfq85TxYWyxR6CrpmI3GcbYiDhof2LhVZO9G3U2kdm8
VdKDsRXFyHPoxNO/QC3Cy6iBGkVglD9e9rvSoT4F0ID8POLe5yPNLMhrOcH4
YMJQG8sETHcvkU2pu5D5XzmPAKr7V4xlUqmOWlhjaZfmQNWBix0qD4CjXwaL
9scqOxtYuK3xa/+pjhlVjDH/37ir4/KnpQGg6YE2SnwppgpIIeDVyPBk7/xc
CfYhg1yavZIdlMieQJEU26UXHouRxednOqrgtysKQqtZpxATh053nxNGvDbs
5CdUxJkQsTFrWUX5HO3F+WlGNuwuDL5AnDNKIi494kFG3/Rgth8xKcAQtBHQ
YK6WC3Fkk9V3+FQGgki1ko6yiH04BDB1Bw7JV2hAHQyXbLIGLUkBtJ507Bcn
sY+WPD8Zhh1GNZCI0MW3KSKg4vjp4UwbJlkvfJcNF+AMgq3xy3baE785nYlo
ALCuFJ4LAJv77smR0I2pDjuvemgPRiot3A+hoY4EFU/UESlHUFoTz+Rd7Nmg
ceh4gGgdSp27hikgqIluhIGC4lcX4M2f4jULDA1PD1cb8YVHXj3cSAu9zmjZ
aOpGAY2IzEA5NvbYK8RoAazwLAL0v+q7mFb8GE9mOSJLuwXezcfz8Q2O2OnL
qpLzVlVhCVwB6X+g7qD0hjvqyl3m2BjJyV0fAPn8UyFtOF2vRK2Xq7CImANw
9RAN+2QJV+S1eOXFc1dL7yGBC8f8IOnm+3+FszF3/0lwtJA8Ve3eOUxYnwm3
yVYSdQQrtQ+rDOhVRaELXK0gkRQ7om6e7nVFjZaWyOJz7afdwrhPSBNDHgj6
Hr4Lj4qsI3wQkr4ZUprGVOTz82JMnTSVFdh4lCAyS7iujoL8svGdImqyUW/h
4aoRTgB6MOOOzieINhAHxWDCHmlUtI5cWx8ulWX+8WY/Hz2BEx/VydlnDYys
HEzrNlClxApwrIA7RFK66lv5t8iuHHLEQE4DpC8PmWDFC8czwU8Hi4ufwhYJ
aXbZrdxibHsvF79zzzmYuCqzAZ5JLY7E61/VaeoWIrKrRQIk9tOqX4I/xkP7
mAUXTC+LOpzlM4O2ogw6ep/rc90Oi0V4WR6n0z0nYir+MLNqecQtB5vEr1dL
xyN+J9IrkZjdenx61wxDAceozaZom3Im2Sx5uAMFGypuGf27mqam/Al704IH
a6v84H5ALACzm83aouQ+RS4XRHkB3xBUWhYitoLvhDJGYPhD+SpVdaaeMJJ1
teCbHd2VgO+pJgDpCxMk8MLnuIA4I06BIBdy+FpgNOAAel4OwjNOdC+H4akg
uqcTtE3H0+BQ9KTBWmpT1Mu0VGB60Lj/sFfQqBQj0AOCS23M+PVqImfdD4Kk
ijRTY5mCGSmsForeumQ3wlTyCtufWzwmxfkFGclZHghMoidW7rJyN3i0WuHs
vPfuO5qINve6poF4Ii9kfDBbp+6TY9Z1uTyeb2PCNVG/r/VI9AYN1gnPNvqR
k1cwcBnGUXO0jpjVy9MPWT3cRV2vEFHSbXG41dXdC5hzNmjlse9HpUUlVOFh
VrCm7tLDJ6H/+UFTHa2IsrIB+9xSAWc1zaPdqj93527p4kx6I07RL1HlFm/4
UlkfI44fMZWuR2XQT5B+96DnsTPj3Tkd2V84JfUb8+KOpqeKfTH8eoDe82d+
SLs3cikRpOvKKkBonTq9MQp6GIueH7yAsmk28YNdsTtKLD9KPX6+BfTj31zE
I45DhjzcQmWp9rB+8ZpY/cfZMk7tNG5oK9z9gy0a49LB3HxmVSkIcmaIME9s
BNsZyNJvrqJfAQvbVseqwzq8iKNgkOwIhA3ySAEwiFhDVTnRqj6SKDgwcVN+
aZ1jc2Kz6EVNeQwXGUmqakDHlHOSDNxd6wIRyvIyG186vy1ipFSRGkvB/5q0
Q5TnMeH+l+cHpbK+B6jFLUHGI0eqRihdgi2sR/CADCm7UtRYHM3I43xxzo1A
3uBVqO2KtSBaOOptGxswE1gO1NSZsVemLv3mNC+11FkwNAtsK5003krwUfdM
yq6FLa7/kD5Sq8FP4VTMyyr3VSROSZqar2nZSeyVim/uQyESE+denIXXFMTm
y27HSnX+7seMI8eWrIpznIO99R9ShyQV6m4V+qDXl4GZXFHGXLoSjpoTGDZm
p5OrxobjXZIPtl+7BMoTwnGij1XhGk/YeL/NMSNY/tjhDBsrmGdkjCtC3Efj
7FULtk7wMwxuet6R+nXJSKrJ8TY8iBiQZ5EpOgIBGwduQuxRnXZ0S+7zRNw8
nl+ir6hrTANzKTUKICcO2FbCP9+mrZOmn2SIcO7jejJtc9FY3yr3FIT09vHl
TCPmw5ZHYwcDaPX+LtWC3se7HMxi0d3ADHfNdaxCZh3LK5+xC1hVXzsQx5/F
8qd44VxSfA2OwYmDgRgp7bGEvMyb4JJORxp1m8wx0OGwJqTTe6xQYAkyM7wl
GY1UBOHCg0LUryTCZ7I2OSnb7+EbppjQVZGprwCNx290plBtXr2Ox3o3kQTd
cMz5drtewiXByU3xp5qM2qSU+V7lUuM9s0Fy8ylkBX3ncOMkhkQ4ai9hwrq9
dx++q/hq9ifsWDNASlZfkMnOS9shDTc05fxw4fn8/dgOpWI6uFHdHnTK6BxA
GTyxE++xZNhCsjwojqWo7hxqyvKKgUBL2QtIHkPuNWd1+XDFxySdgyKABO82
tcdwMUpzhLSoWqLEWFYWfaqlvIghOkfw0VPM5ffUoD1p3HvOFjEQxkhqR6RL
wsoYDmq8GG0pMctbKMreIYidEPkiTp7GqwxQQqDl1yuiPCWqadpdFdrUA3SK
+mEYquPGskNm+2PgfTvccgM33vh4fc5YF7URUdmOtLB7ZljAKDakOLE+qrvD
/STcbkozysIhyXLs5lQMNV1gf5F+3N3aXVHhm+ZzmKg6Rh49AojNCnP7kfSx
rjU/yq+WjJWiNKcbktUfNFOcVs8PUvW9tm0u9tbercNuFxVZ+HXLCSOL9+fn
vwE9JszpZDcmzMvC7Sj89eerKFu6IOtQwIaSddN3EV+0xGUhYGk6NARExL8l
vJtt5zc4uTuyB01maF76ZsNjwtVz/+b6SPc4gcdZ4ey16jx/z+2rH57N2QCY
lrjSM3z6W0tGN1vtW7LBc3rUzarD9yzQloeSRtWlotIP2zqv2tFmx5eLPWKh
6Cw+rlYWPFCXh2ztOK4EjEuGWagyWuG1e0w4zsQR5fBWwbiX1iV5rvPeEzVa
ANH7Ac8hWn/eNNRVxWyE7tdcUe97PUAg/3au1RQp2FMHC0VtzGTQEglejrXW
2dT+GskLe8bIwn78gRI+hw2Th6Kkb/BeSEI2z1uG8Wm74bYSc6U9eH67qJtX
wY6nV5SodlWglFxtB89sT/ziL1Bb6tG0m0JwpLNXFul1rXdo3/WP72/h/Bo6
NzHQymdHY1cNSE4LBsuQlGF716AOVmpibAEbji9FzfuY/139emkZU+ZmY2kr
SdCSif08uBYVoVKO3he7o/Js2aGf5/0Uvr3eUI1LM6FmeT6AqdwNLZrLKxhj
thSYvfmS/Ie28OiqNvYwdp23h27euu+791lXMQHqEe6+3l8UlN/Ua7aPkgfv
qgD4OlXPn15usW/J0qQIdwWWkJA5NKmMTrdXe3/QGtUCCrkHurjk2fP9if8B
DhKz/2Y5AQK73ijR317dDo/CYTob4TVnvMINPiyp2mwcQ7NmZuRief9aVo6t
f2BRgNPDHbIwm61JSBRSyX7dNH1mW1uoL1Jxi6MJsJ0SU1NMKJ0RAFpzekL3
rE/DVd5Rl7xzqgkyJhr12Ufg5zwBuvhNqI/p/hZgulQZWtJc31nR6Mns0/8l
0zZNkhRKQLNMyWUKYARxfXuJ5foINv820f0wpuXl10r9ro3lDUt7Wv6G0AU9
wR6wgrzV9XDTv6Wf9ssUNB3lk55iutxhLlIM8bBHT/hQnxXlp/Pdig2lh6NA
+wiuIn8hihJ2kxk45z8Zec91vOGizDqPFFDhQ7x46kobV2h8rLhQj6VIz3Kh
b66Sb4Taxsuvw1vAALT9kZPktcAaCJF41cJFbW0FnRBRZ0/IpmhcgLYdhxw5
EUFc606z5UU18wru4eSP2llAVy5A7KOeZ0g0eZmUu++xp+T7lZ+wEdvbDT8S
fiGIpxqQVbYR/I2OgL4dtlCZ5htqjycB1OS+fXK27Kk1CsmIyKZgX6mZ9y9z
9RXTaXYJwOx3AvuvoCjlsMkrzPeB6Kr1zsTiAGopCAcYzTnmRtuoEa0HOJmD
Dt6NUPNP6twR2i9CbDUfYvrAA5KOf2l741QCkuGmZpQHR5UzvRy9Ymai+y/Q
elQtOWDXVBulFbFidvE0PrUjGzKw7g++1kaGpfmNjSJG/mK59c/XlcXTv6lt
XO5cRDTV9lfKQihT7rCEgfkaJ8RU9BBO8dCfnAFsJ0VkvRNuwiPfGcCTw1Oc
ohoG5UexTu7ayU+xaZ5bYlXNMh8OFwL+38PvF2bmPIHIAo/2QNgGUtORCbYA
rm5sq8yB2AgNKSslZLOgbH71RPTrRexXpNwvm52pSxlUijpBCYtfYyck00GD
PBu+GwVmtjpM7GhzHNEBeXhN6Zpgd444PIkZJeVhiq2JiHca7/hZqfY51upi
IoQbDv9701UU/3MtRgWDaGpsIxe2cDsYI7C8P6jap/uV6dm2sZ8wjQ2BOTb1
7ct+3VgGzWDfPsvGrtzx93zwLZJZUHfwkbsEiUDJMcWzaERIbwxi2qvLxY/3
L81Nzh4W5jY4cythdrWSgjZqbzBKJeJJv8ir1Oax9f0o4XWdbyoKdT6quu8L
zMvZ4leMoW8q50OZeH6eoVDm5EiOBWqqt7ACkLYQ9LIIO95TKdvV6+oaTQub
rdjvjRq9pse+gZFZUWPZ+jq2I1DXtFZFCTgK87ZJN1AO4/OYHV/KDICOcpkZ
Hq//IsMcnYiT9Js2LaxfCFOYbpNNqrs6HIYwCfKl1sI90O0YhT9XWDsIiVVx
0keIXIyhFxz+YnkL4wB5goWt3oxDHxuIbHoJqTSBUgoaaKsEHF4ggyW96wDv
KRvMhjZHjvIjE+y71kR7h3sjr9Z9OBzbJzBG4YESm2YRUgdmwhHhTb1LIXuJ
FE9hDby0WnPavaATGA0yh0D4iOReSxmQtMrLcC6M/q/ahd45eeOsVnKQ0Z7x
N5Bmpj4lf/igH0c4MIOsYVZvT8DwG7xaebz+foz/ZQNSVykFV/o5t6sC02qC
JxGN4dulrw9y57SgV2q5jTLgeMNNvCzAMn1Q3R1fJQAl8pDE+wDpcH4APETu
p3CzNhMP5F0bqy+70EJEeAuw+uztyVgJCOYuTEIOo/OM9ascY3vRKLRMMgKg
ibSKqimzp7oblWqxd1fG/TP11TOkEiLGNsO2v5HIH9LGusu/c8Li2sh4rxEf
34Zl1nKCqd7fNchvEYZ2+alYsuXgZ5i3hrjh9Bxcju2AtPF1e4+aebtPPCd9
obvclnGJGIw6QtQbCsIE7oeltzUhpHxTwQKaum7jKdE+cDHuiqecUlF6SC37
CbS0XZbZ3FndzwREm+AQCnEgcSbRWx/zM1eKG2t1XN+3QeIk4O+fTxSo06tT
BjOIe7mWt3jhqsqiXuDuoPvC/I10AKaBo2OzrHHD0lBosPwFxTWinOHSN5gU
ZAvQCS53ffqq0INcxk8CoxMcS8BDufqyRymsskpdRDAdgUmZ4YRgstG2h4oL
gqAi7fbaGWghCokhAXmPocO/N0AQ0q6HRDUSieZfPq2vnK9Lw9J+FdPjWOZq
0R5T5sgvu4Me4IwojDLJKmR+RuGQi+6xQbko7qiMWgTcOG2DrjwNwwOudsij
GIF4dQ6hn/tBAhkcm5BQHMO9Csjx7W6GsHBpRZMCgVjYYaJyR9pr9WL7w2Vs
urF0yx5LfJYWxKzo2gMu0Nah0xMN2/tZwrkpipB1RlPsrqKB2eTuywokMEFW
AXSpNQPrgxPR496DD42k3EYAGit96upw+yIG2yyO/mJQtZ8RLozK1I7B6b28
KZUuGFA1dWG46cD10oZ+tQh1jygx1eXtG1ASWzNE4Nl6n0ZmnCbiQDvHqvKq
d5VqhLUmj90hngpptzW6kQEjDKEKveQinIP77Ga3MrVAETPo076NrNWrB8S2
znkedcMVRzZNYDNliK/tIsF0fX7l+kvEn+FL7rhBuMqqqxdhelbTzcsT55z2
sXcZ37FzLKWFqivcD3MHueeYxW1aMVhCWPAMI+ktzxGrQvaCbOk2sRmm6kxI
2Jhqj56g9LUBsYMurkEwkpfZZeVmGQGUmj7MukR6U1wN8/3Qi4g0w73nSBBL
BMxC4wIDtsSxF+RjwdAo77dA1zZz6eQ7l1CGn6urbVlrnqMT+pcIJe1NYS2R
cNSkVieASnsxbzLbdqX0UBfb43WH9UFWQ8/TUvTut+zYK3CAqmlnFJBFiZ0b
wgZkdnFNJMwh3bsb3BhNg7HY/Ka3cVQyOlVH6gA1SEogXuqn4ypsWnZ1YzRd
s0TB2WyTBbE0kH3rd/SqfOmBpj8WEuo67tUXZyg/UyCJCpSKJNeLRtioATzx
QnX/9jchc67EuECPNaGwWEn44Vt2nbQ8siwOUK70K8kL19+KzOIIxcdruRtM
1iE/uFEmxPBAbzE5H3m24PYgUOzn7qhpa//UkE8hcu9TWE6z14U8J6To0Qo0
VKxkUxu+xbWWjj5Wnc65ZNCHTrVzt8sFMxC5eV2e4eAk0Cv9Kmoo6kt3XXZC
cOR2x2KJiV2Eejwr/UC2/66+L0obYbr0fJTWGi/jGxH6D54vcwiLlDRINflr
wAFjIxvxiPOKUpvbc9yP+NXDpzF3Jx+jxMe6WFqTGWsKTAlLDZMMyBy+OX16
6XdUGW5kcxHDq4UESmhFwyZ3fy0R5W6MiTqLUUyQ+0e91HeoevgmidtStO06
y1LvRe1QwXFKTYrcOw+X909PTIMUemPMYt7zVBuWblkH1MKvFHxpR7iiRuYX
7vgvsAiXwrw5bT+8yXkUEQErD7Ymt35dyjlp/9Y+rVk/ZsbOsC5VlROnO8BH
+LJOJbdpvzXbB9AtPuDEIMFW1OhSaBUT+qzYj3AJVTHQW7p3/nleMsIFTlE7
gbswkTDefhBhKKvM/NM6Ac5iq6B/yQzLWNTl5eLz5t/+aqUKZA4dZ8Zmip+c
YigFFTPlqHrBZwKtiyWbGygRWjf4f2OXtL+cy3hEGtBPAGBS0w9VADLxGsl6
rm04TPLvor7/V9oc2K47UZ1jbH+kd3DMGCUdLImtUAFyF2CK+dFJOcXev4sf
Rv5OxtVaHtgUvfjtrYgpEnYcWYumHuXHydCvTIHOB7VtuV03q4U9R4vqBhn5
s7VY52rYiooOpCIi43Tc7mlW8HE06D1bvJ0Zeo1MyQ/I++jfcnX0yu1hvKyR
PyJ/7Zfdy+gkfqF3guk+mw0y0ramQBbKfOKKhCmDRQw1422s37Zu91Gstvt/
kcpU3zsD7VqC7jzZp7iNnywOk0tQ/ZMbPKrtWFoEdWQZS2SvjFoOWCpRUUxM
sA82oi88cI3kxruHSS6GXexBYhuwFclyOJAzTuu7teUDWuVael6or/KUFngG
emlvKg0S7TxG4rORx/tKLPeTznTP7SHBUcAMbS9zy3dm0ru5Jin+Z5iavK2F
taLNB0GGoEY8sutqipqNq80I0wBh8IJUaC1hnDcRClEqfoo325xDb09R88Uq
cwQB+JyWdtr8RKLqzEg9yNJrcJwr4rhwarHKDTUlQM4EK7Fbsf+m/BsI2Wcd
gWQ8VmIpoq2tf4ZgAVwl5ekh6wmkjVk9UZxZyDv4zf8qj2s1bBFXxnPNneor
Ij6ikOh8YT8dUZmOhlFubpV96m0fQTNP7p/p5vaQcXdpcn99KD6Qk4+JTlPs
OAclfv3x6FyyJG/vr6RNEIIYpmlkDaPSUtnTnISkFQiZTy6XQfg8qlBBNW/Y
cavZzQChHGHxSSEreNKCNOaGrd1edLr/jFQqgPpeTq8FxXYZMSUcEUtmHHdt
zKAe2YbFqDxQhVYCsNunWUSBAql2J0nEByde/KDUXk9SwiYdoNQgit8+9jN7
r5JlZ7QGRok45AkUsh5halTSAFfoTYbifpsVLfnO5EzR3hkqRlUAvH3/FRTb
doU0DD1sH/gImnibkPepkrSNspVrhNS7SEkpQHVWuEv2qHZlm24me5+SwgJ5
Lgnd+ZNvrTnCVz27JQJ4uwM9mkzWuR5L2bwmMgVhvBeBYfpVmIqx6GLl//5z
QGsS1IEbiDZgE+3vDHzMnEO0WTt+rfQCRNJzxRPLMDrZpwOw306IC5xjA4cQ
pQeQj+BCKylM+HrrX2e9Kns6IeUQwEWkhUVLctYy7IECDIL8Ynj+hpLPNzGU
wC30rupJwKkJ3NqmhGKiIvD2+4zmd3zYyaqOqOsbE73nVsCjacP9f4xbBHP5
i84syfFLxkS1YTFW5pa2YGo0aFSxFCl7l0kAs3SxfhFuUDipAWviLBG5dYzn
sLXR8Hqu/nQ9ClVhrHsw8HJr9ZrIK8z67nnCzS4Js112NJvUeVdUliZWhafW
wtyb+dVNfilGLHgaL3MGbbLR6DSmOznDRxax3Eeb4WnvGNwYRpn7CAnRZ9+k
dc7h6T2LJlKKvjOE9jBeuH/yCtqqtEsMmJudpI+XPV5/98qBscGwXycxYCVp
KoAlVTblFEsBmMKiEnlJF7QNm1kpzI7s1R4XUMkhkEfLL8kDIayojrfLcgLa
1lcOtigbIvhGfB6H9VJ6vD0BGWNCoDxsWiToGWO8DlDYKSHxsCHmf88gDshp
p01hs3P55BnrUTgTo0jFrlsTa7bTQWirOkBWuJZ5+U2IYLt65M88YZUArtIC
aGvFUREMAFgabfokAAY52uHOdGDL06PW1tyadUCd46QztpAIlrzOblxnNMKF
XeZzEblcFR7sBNQn1Crp6AX6f7DPMeRlTdg/p0uH2Fjr4OfyIzwSi7slaWdj
LoNUBzb42EJ7zLTGnxFEHGz41j5Te5vY/0C6cewmQeWWK8RfqFcFINk7d99H
SPTDflE1uzO79wU5UlxzmMeiPXM3PauFErj1f8pVEti1o4ozOorLcTjuQzBA
DSvWCqk23fPvnGzMcXD5snblH3RyCGxwu3pSZRxrYyO3qK0IHbJCtnT8yLZ5
98nx6OHr4nFNHwVdVbsCp5dgju70NSZET760X/k2kHE6S6cj1UUY9g3Kv5Xr
m0Qp/guW59leookrJxB1zMA8+LJXA8o7xyt/XDSoLgkyO0wZOu8QXqbt1mL2
m/YjrW5H+Eydf1RbgTlXya8MQwBI8Gb5Ew+UH2eXhJSRVIWChy2tz1Ijl8+y
j+qVuC+3nmBvS7rAX8LIvdGqmu5XDdiitzUQddkX15w7bjHL3Hy4ciaLabPu
+H2FXrm7wVluwNvHQQtKcte0OYZ3lmCjuEX696fYNHoMqScU/74bEt6fahfs
VlEGpb9ApMZ/H5Szjach+g6XKq64kkwsbZTPkxzmsxAFHNmR1g4tpTR8PkDg
ECljNqhQWCLyovfw0HdY6JK7wU2vdjTEERRapFHMJ8TeZrO6MPevV3Y+NlOI
VS3wU3SGr1Vrep2bymBFfz4d5DsIBv9Fwrr+fVvJyprpfmOmho/Tmltki5a7
Qrfka5tunPqEJtQhQXkcohSSc+TIYBfgsK+7Z5LK2SzoVBN2C/FU62uLudQS
diDM917h/pRWhb0Z/CwsvO4Bw+N7n658TwsoX5oSWnIhi0hbmXQok2Jk4Ut/
xOpBfN5ioeA7ZNGj2w/kLmPhrlCozCc2qExqS3H4Yq7OrtGnaYoQhBTD4wQH
FI5U9MXrnIuQkQWimXUrf3A7ZUDmgYMujzKgCib4AttRy0H0MzAoJzUS12Vo
dyVtb7ozz148YcfzxWNCaOMYBIDdozpBifwC1M7CiYKkWwzOy2WUNFt5tGjS
tbqjVMivf0f+i13jtcXLNtZNF7bnL7nhpJzhMmqYdfDRzPdWibrDHHQbi7gW
vkluIDqf6wjQr5+axHfA30WEtIZ8r7fYeiQz435QVReXMEf67cfzJXxAb/8L
rlyLOrrmxRRyn+RPJJFuc69oo+X2oodyDBlIuOilJnoF9CLivpZX5SCUtnjg
1qHQJUD8iFViQc2jX75lktZ8RXZG6E9tsQqoXhoD7T7cU12Uo7nAyit2E92U
3FgoPoRIFSZmbPPPMsSicYcWqx60XXwpNRbMkKBikTe0Oga9JvkuhKMFfIq0
szU6PdyU2gwwEatWvX6JT+KIMqkvSxNgJ9DUOg9AQZHzzVGAjS2BvbsxfUkx
SGO7g9G/ixgiwp3fIrMK+AfjEweV2NYDsVf1ySRURFv27LS58+DJMglRSr6s
kaE2QiRU2IHwYZQrL6b8r83DOm1vq2e8/ePntiT5iHltPGFLRRElmGmtN7Hq
Lh0UREz9pHInixviSUB3mu/MWp5DnruMf67fkRRRN60wOkITGn9hpSCzrE52
gR+dvCOZcphuzmxChg8GYLNvxOp8GbQhU7jghlAAKcQ3HewOQklKsxm4wEDa
zMePnmWFzmwHhkqKi55iaG3QYyfrUKPW9hXKgvef+yi+Ngvl9JbsdjTcqVXR
iqv4AvjgLzIQUO1ra14iiymL5++iG9AHlnKZx2qOJq96UVWqG5WACvje6Ady
CxcojmZXR62A/W8I/JC/JXBuWF18UgrrTmKkBcC7JlUDVNBEVdsz8yY9sTKx
6Xk23J3Lwg1r4GfORpoo5+dJ+27vPS7vOcgmVQUaX8WdJkmqVUrgSABqANb6
8HMWvRY8xamyJFatc+Sy+D1NXtVWWhvPNNdBzeOjDejRNMn4RUjvhAS0LevD
nUtwbFj2YNzei3D5Gmt7M0Hivx+tsvasWDMwmBZ0twCRZrPCIVgXhX4U1F/x
OUbZ9qJ+ZbK0yenVtD2EYhbH66ZzqasBcwZawlugAl0cy0BPian9uL1u1KJQ
YvKH5iaUo1ZUlhnVvz/jG5HJLHo30AARKZnN9wAZtBRgYrGJhwbOsZy5lRPE
B3+t3uazVW4H6m0LUPOLh3yHKJz3ccqyciS0pPqatpGSO2lErkOi1x53F7DR
oiLpU6sU2wxK+0Sq1c9QkYQlIvUfMHVqJJB2O4agqcI3ZtmAaSGte6Mh6vG1
AAR3m3KLmwzSLW62k5tw+35/UXCNxiaHBHmZuPIJ+fLN6cruPJ4oJaIXNACB
FnJe3st8yOpVgvwIAV+TI832Su3aTZfYPZzMurs0vrSEvRi2yXwlKLgJcfh/
cTAG6GQYyGWDopj38OXU2HAPjor8E5P9S4rPSuv/VKwtN2y2Bjabqn3nkZlh
LjbgGvnUlyZTSmnTYnKqZryKW+xw5OPYA5eN0BE5fOjulyJf5Ad4sxXWsXpP
fVKtuBuh/8qdNJ491/8XTEVY9LoWs0kHLK2OjYiqreTS7+0LLr8v/PZDwNH9
8eOEouddZjowqe5GhenJFk3+UMr7zhEpkI0wrZV/7EVodouL8tVLrSYVpKzd
xy4KoAM5gv+11w4nCgLyNIMCL8AlO9ELucFhCxHky38MBan2YziPZeiRTZ2I
0Ffhi9g8pkg4Z8HC0vUfdAeXfky0fXTCyo86kvoVS2mry/jIbI3h188hS0vf
MzbHz1FdZJc9GDaJITQmBzgE+UtW4rwLWZ1drZiztqwddTbMEpEIZ+tEiC1q
Ile6m+wXOSBhTTRgY8jt+bwoQghFSrq6vKYDXJeCYsIr2sxsR5PpcgsmytXQ
d2//JsJqbJlV5Ao1VVj3sfkNNV7cPrFEH1C6GbX2tiau8UwnHp/b9RpWi4+I
6NYawOQAgTswdLaTB7d2ygm/dj9dG0C+PqTpLxIPN9zT76/+ddFNZ7aIjFcl
/X38EdJ13ZYIcA2XRReJipv5iTwwypZmUzQtf6LfEMowlr54NPSjxXmLOb3y
3NmVTmkAlaA5067SpEHDwsqOoTzX56ELX39cI6euFvCOdCdUFCPywlHCIPZ+
QA5NkWnlJndhgmBvQ9Qic2ON1j7paZuj4o6IBjp8tvf9eB5cKW0dPvxiJ1Qk
EX9jRsh/7MASiyltKSI4nNpRbTqidnRusR6M7/j9ue9mLSuojW0Kjd8TZ5Dp
fr0B5DZu908mrn4N3W2MpqJFK/6/7fkoUog6XjhLNhQ7s5jLqxSis6Mp8PP6
K6BQXRnEjolFNQwDJSZEbdzb8tR+eYRQKp39XuLRetD/E5gFphyJYtfVqRtZ
ueAUgRbXxQB0dsv+Vm1PSta8yXT3ic8IcP/d6g7FxYy0at1bG/nDWVdArlmc
0bqi0UJvk44eU3M/uc/1C5ih/dBFAq5VOyZo+Ov4jz0nmHWJiNawOrNj1Jxl
S8HLsoLyNrlxSYF0Bgy3kyG6u4PMNiyWyb5YuwgFHTtckL0RKgp+WSbAD9V0
s0Cce86P1hPvUY7bD/uWV0wpQmsfdc91bxZ/6P6OfOgKd8qWeNHY+st34+iN
wRjPH1i/v1yj8kzkBpl9AQc+47+8Eq8TBMedhct5sVYvcEbeq3V2cDbwbINZ
nNsDZf3e5A7exPatmPheo3ueTTEDt6VJtYtqMzV1f7UlW07B30W5diHxCeN0
YjLa2P7HeL88jgqKit1hDCXaSmfvi2+kLSVzBAoI5riV8A9nfhQBi++bms51
FTlWv86IRxEc7oF+sdzVx4PkbOJdP/k2DZBAAFndUg6XLaGYNwJo+i86Qhw1
BJ0h/wbzu+TDNj7/2FPG0bjtDazFnsrl3hUV65wNHmHzG6iBSgiEKS+h2wU8
TAQ542EHFs8JNcrW2e8ZUvnt/j2td3/F14lXU0o5Zv2idA18yfF1b2sZ4KCr
1TE3CEq42Ul99RbazHq2mXYyd7qlSbLYUfjxGWTVYhb5KBaPFD6LjEljKA1l
ECJB9zhDD6XWP648Dl66+W6gcpEJ/UL5mPUy2PFphT+GxSqfGLcYgpHs6cd3
ZUoFadavVwcLXK+365yMwsBI+W/YAclXtbAQZKUB6MbM45DTP1u+F9VWbPNP
oYXTO452y//xzoC9RDiP19Lp8p0Aq1zZzC+jTeMR7ROW9IUWE5XdiaG0ysF+
OZAJekOEfbrWoIOIBafW8z3M5fU56MhCNkHlp8Tq30si6FfIl9qcGclMSKjk
uyRvIch5lHubBQMY9YalOgBGStAmmv/GrfTGEfDVQjiO4Dy+bOiCVf10pMHG
wqxTEx3iUFUA83RfXgi3MOSc+L9HSoFGM6xEAFuvw6QgGWtidzZUch+lBr76
8afnD+CRWi4l4YhEkHiVV0VxXf0a7S0+or9G/h/Nb3sLqDIYEY9RUsrqiIeg
slMuWKEhmxkzTPUChxZiqnjdBhP5tYgledTtuIPDILSSZpqThZuJ3Wujg3t8
ckwWic9YTt+9YnDiXHkvZLWazMlD45kovNH6imER1soHIFIpSAhPb80KItb6
EJXkKwXWQk74wi9fMFhsi1qq9TjmnZ2kdspHpFRWymg8aEbQoirbTyaM4l37
RZR2ULAWWi3sx9jCeHGolaiwWYqMgS8UPpxfaTxoeop5Wu/6/Wd1osC1FMh7
fJ5EkDWB0egpMvx+7miQY38nDx3CmiiC/vP6uyR3CZ5lukeBEH0v908QcWEG
0HV2q1UHrSgRoCDs2q7JqDZ38cTJmBkljI7+xiYUFMJi+wLA9pHgm4qGGTSB
9U/On/h3iX0qgCMZCXp4+WYADA43ecg7X/Kj+P2B/h3cJfXoDC+wybEoUkkj
QcfHZONmvVnnL/a64kgK/HzZMFzkgK488kMguubPpm0iOJXrCffOr/kesNpD
Dp4G+BWB4eCvh4ZL6161xuDKKkgb15DpcIF7w+54RBmGmm16th12fyj73d6b
wg7M/t1OI8Zp7hQf/ht+6UbeWjJtGIfFb5cDsx8M3pM77OwTu+IuCnjH+uZ8
8m41YJfG0R3/UgY3LlNWUtWT3eL/cMPjkamYop3zgn/NC6vTR6u3ZxY83vEG
wGHW5ptWWbdyp4TiU/SrJn2pmKfndYn3aGDVm2hKNsc4ooq6CpIu9mYI8THk
zzSm833402oqL0xxSKld9XQ7NvRilVLv6cKx7A54oZrlFkLEGt+KGYOlx/2u
MnFGc6kDMnTwM/I7TZJlmI6jtoLcithn0zHXsHpKLYnCConG0GHwCMVpRsja
B0RGH9518ipSPJmQdlNyga+J2aQpbUFwCpYZwRRy/dnMpX3X2KoS2ApBU5f4
bXIonAisiV6QO4xzedQFQudFaG2csXl3uW/7s+BIx4y+QG1M/y5hcQMHU7cj
z+lLKNdJCb/niaVYB5z+VbTN+RS7sYoNzhWmqQnwBuYhH4RgvFAQA/WJoJ2y
HbEAs+lcEbkj85VtFm27D5vJIDUrCxoswgjPNqBP0mf8AIBVYcGG+I6thHcg
/zXGWOm2uE8WwU5EnrYilBTOGrjpp1R+zf34qqLELgNAxKUgqMkkY/dT+paA
wML5EA502H3an1A0Au4RcxyQ/enhN9Hm3eg3JgfiuWKkMNnDywchVznJ5qUA
hJgnTlB4wh1Y6heDFZoJ7EOuFTK7/8OKx5IkbXL3gbdDHQF4Url5rSHDG4oq
/OSEKSjhgBkYV3PtLSb+SMcNtGSNcUEr3Po8+55jMseJiu8EAkQIaSA2E251
oijair5yqdFfYAGFCbK80u6t/ubOBtX/lhReRLJDwZ+gFg5asD/GrenpoyKT
eK8m8VWu/tMGAlxVgQCzXClVgCN29znKO74Kuj6CExEiwmRfsEzhQSwEV3k5
8YTfXFNEy1DYD6HUlspLnxq3iEY9sX8E+Gb9dE32aBMBSEhh21CZxVw7Wm1O
7sscvdO84qoJQMG2VTC58moSS3HxJk/wmLlSsR3hH1wdWBvCijR2chLrbkB5
2LlONG+92jN+mH+3HVfYPCDJesHKV51SvGcf7yVwdRu1SOgAdaI5RM0YXOtQ
mps/hsscRXwaSkvpKYdurD0Xq7iAjaopBeB1CUwnr10EvaNqhu+v5gueAdck
ydJmbE0ozM6H60NZ5UUy8w6t+nHXMGjEEFZK+Vi/lxProlXKS3266zPxTnmQ
aAQBSY9Dh2634sjKvRPhK5UML7obaol3ygjvsO5EUB0fRwn54tuq2a94JQ4L
R4SKc8F//mTa3hDXCHiYMdoGrZ77nlZUIFUEMA0mdVnLmiiJLz5yopczR0W9
jEsIKYq/dD3x56KDVxn/LWwuB+uuVo0EF9S576Q/SuQg+PsQdNvVSYzXcIT1
c+XPElj89fQ3EUEKClq7TKIMeqVaXee+2kl0QusR6PWEMqF07gkFbc1jaHDO
dw3cuGrCglE5mY0LaHN0bjRrCGoJvOokhEIm95WlnNqA8kkCA8T2dAGXRS6u
UTtN51dbTJUQyPN14sBI12rfI5xwrZlvfAabVctR4P0E5MpmHkKvm3pEOSDJ
jfPtd6/TwODZBnXo3uCHCdAafTndXv68xN8t+aNJ8xHsYtCMTVJV4u00h426
EmGAy8BzhGYDwshv3U8YBIteKgC6u4fUGCxJFbiz5ssDQkknPIH+2iRg2lEA
c46oqNk+mrVh8nW9czhCOHDaAGJtETu/ne6uunU7OlZyXAw0Vnn4yORL+/WD
AG4C263JBglPEpK5Q8/VO9Hvl0UfZDkIEniE/r3qhT/cYeAVC7fLUAq+Ir69
PLl1pqQUUwXtI7k6mp41EhPLfOrpV+RMg1o0U7prf/tXdUwI6j3k2hM6iWa/
DIqcP78o1w1PbV3u7deCx8rVHHdqlT2bwWyaHmALgolKrJ0Ra+szQTa/9pHb
CPxSqQKVwQhQ9J3Nvxtsdx3YyQEbYtaJjJHGYClwSUdmA9t5Y53w4lOkV8pT
IuFHXwgVcwSa7hdQwEnHEJwjHelubrl+Q+AYx8Lxwrhw/AxwRYVTxIUEeL/u
BzCXwiKfmmbV3AtcuMGMHf1RVN0vtC6lzhKK9rjGjrxBxsQiojcdjLdrZ9LD
gLWhb9N+5Kte6SsGLdCQA4/v0H7ZEObl0c1g8HhT/xBJ1mIXYaIOxSUzIJW1
ELHs4UfNYRbvd+46hJXTUzcSzkEo+K5ZEE73aAvottHPJbqUX5yNVmTzl8Kw
PY5tWUP4N6o4e85/5F7j/0Pqvz9BMafeD4Fzf1dFz2dMfzjWe6vUspM+ft/6
Y4S5+tIgAQ+8sgrEE8t6lRz/VQsMU+ietJ+uboddGOBBd8rjwd3/LGez/fz+
UhNpv1HL6RxxxvK1zfWPqr+LPH4PyXBUFu58rnVdAPCp4U8Gf0fX8euWw5Lc
8Q5cFzK1Oe2G4pJY1uZCsD68UnD6OTyvnbntYjm1DOaIrAmILtozKCpdkJPC
dhUjH6hG/NLItKT74F++lSSOE24KMBqmQO/gyXtLZTbFyaeKgKh6bm++aoXG
ntCIzE5lP21VlYqND7BgoktpJrJdjI3c0qdTaY+z86MDv8xYibMrKdtXpbnP
aZZrmGleXRdvRBcihxLj97Av+nQaGxjgwULrKeGoGdivrEjX6xh/8Njuwpdn
xjhf8oLTFR9jdmHSP8BeyMeWtGj/uNGQNS508SLsWKSpNgYzagz238SqMeRo
8RnfsC0bJVCKtrdk3d1hKbmDDMppKCIQ7uGT/EPBdpOuSYVe3GdsgSQuFbfu
PhouexlpbzrZofw93f7OLBv1BMDybcOTavZaJ0Pl94CO8/Fv9op6VqLf7gcK
omHI/j/Mzh+6QzHLY5tgev2TMXDOmzvaeySZrhiPr1i2PFUFpSRa5q+vj5wA
7xrrcmnWKhVv1/gRP12HvYY5JgOsTHusLKiT6Gsj7tThVCshqlHUBF7v33SM
pDJCO+t/nqP7CzviWt7ZVNqwf7VrmRTigAxcwTHour4ldP1y2rSYPF8elGvS
FjvTv0E48MnNWEJIilwdfVaTuc6MIVGGx60bUqq6db9Db9CCKPFGrRJaqWO7
Pye8+3PgwumzosNUzrUutu3ECJ4Ou44a7Xa/iNQi4BmkTs2ZOEF4mqoVsmBQ
H8x29dP5YtOe48fVDvVo65EEb+UAt4mvRZl+Dty1c6LNguTdXYkUiyZcyPX/
C/aBrxbhG1WjFArp7UigW4K+wZnCxql7QqmHAHmY0xh6bEIiJLao6rSNcpbA
GqlA/GIS1gwdTKA4UzUJBvO6Ah6XDL0mDZ1ImCzyvNec/J2Ufvlf9KLr8HaZ
Qo/8uJDN5zOBx8V22XbWqxdfiVzpN6R65px1CpOJcstj5pdgrZ1rakRPO7Un
qnlz3QETjEE8k06Xt5XIJlneaFopme49Ke+F6R5Ey3TTfmbzoXrFe/mgT7ht
S4IiROrE2d2dxrWsfz13FlCI7pVFs6J7INaJcqS5LXPQ+ns/leIF0eq+SGJf
Ua9mf5Zc4KSW6Ec5UN+tbmrI1VRXbOy4rwiga9SPsLWsisF+hkNIMkLZFxVB
y2SRekWfdKe9Dra9DxMw+WFuvp7XFVPilU0s+IpXz7xDVZNEndsPLQMRHVrj
iuE60wPyKQ1sZkF3qGi3kjYU5ySp01muC/kHwjma51jfOAK6Q971Xw73SYFD
paqmtch5YeQVL6dH6HB+rvkeIrhgTIWe0j5mIMv54bQl2jWV+Fab9y3eaahf
RKNk9ScIAfAMquoDveFjpr9e+FPGJn5WgHW2jJHPP24NhNFlyiguVr5+0ABr
2UW5oPqnaJYdnul/vx7x2XUN4naGrV7REmS9KnMmudHkIYIekjR51zZ9+cv2
N75Wd/Ks/fTg2+oABia4ZHOGzLK9t9XhX+/zcATdrzr1PqEVe1VcOJMFToI0
yX9gSVRiBE5gE9S4YxRpAFzij5/+Ck13CY0/O4UkJe8RuN+yYE6VFxG9XF2u
1qTFAk/L/8fQODhvlFrO91wGWJ5oSZ8Y4Y3vJCeDsfIac9AYfZ2YwuMotCyi
hejBlv9o1p7RFxWdWOwkI+o0BYH9VUGRX3A9XjxQkp7BCOALZXmTic/5emtH
FbyqEY8j3RyDf0TZh7RdlLsDJFPBPhMLZN5bRAhayA7/40ELRao9HUMQL8jx
HDqycpnxRfjO+EEaEnfbUpTltqV3uUhsreHQIU7o897jMWOlQQBQ69/ydu7w
yaxK9IO8jAeT1zAIrGb7i/C5XXrzNjnbk/Ot2ZAO34t+Lev+oJjn8Ik4NNtR
kXPAWyXA0nsc+sIF3i3YBD43FTtzoiI50UCr8B+R2UW6ZED6kzskQSt2hTMn
lslk/oCmX9JmjgSfxPiWv/Zt4IHmOkb+34jud3sWk1O5AFCHt7ZvfcKhrJlJ
Knl3IWAcvYaYHw2KXiwYIQivJwHodlsrJ5c0+q1a3rmPeci6MjEUzhPbtD5v
D8yEUr/3HH3leKTyE/O9h2DeKQgUJts3ip1TpY4F0J9zFQBVmxwO+XvIio9s
bc/hqgb1jPo+efVWPsJOlXfTrNdj/InpQUax/z9fx4HKOLSvwwdwtCPfsZXB
yZwNsdnmqMhzd+7KyaE2K2+hHGidZn3ReL6jKBOcUXYHl2JPTYzc6y2jC0NE
+DNmIMiWOk4EHcy03fCZsTAUF7/HycaAPOirmcyIj0o8hoYlt6EXjtG6Jn1h
+4MTIbOgGWH99N/gxjiuxQzalQHDiXQruupD8h+SM+HDCf0sX4o6v5QUlLOH
4tqUxdsLusSreOA1JSAhK5hJQm4xDLx/00ycjxo30lanXKOX25w+uvLE59qg
xT4Sarix1MV17fkkMoiFA1/fNeHs9gGBRCx19csZe0vNMFTmzcZhTn7SBw90
sqQ2N1b/HhqugbDJa5/CRfWwkBs1V66VkW+aijR54IZ4h3vn4sHBYmVz12eW
/jLSHXxjkq406BQ/wY4yh3siS+iyzH2JflSN67cMBnZQ9kwidgCqUKVQCOc/
APQsmJsid1Iq/T0Axn7xv6rKEdQ14wz4637sc7umr6n4+4xKJssJQ7zX+1IY
xRnWRVpWlRTsUOOE3DlZA3OYGXeQTKASBVFSQ5iz2KcYQJUfKQ1TorC49w5f
mxReViODOwXSM7gc82PSacKKpTDW0pv0Ers9Xr3JbhGyWUlAezg1k8nuRxz/
F2ZHsPyPRDrRMVp33sOywMIJcQtEvt9I/8uI6djGi/Cd6WfAU0iuvc0zgwps
+tFofT0RPst9AHVYjtjFc1846KEjQ4+MfFvd2C2xd553CMKP4+NTakrze4Ly
m30voWkGl5Ky9KeMOL8DjOxYL6niPI8BmHiFpp1jGWjj395igBqPd9KKBRvj
D1R+sET1fX2VbksKGmkQIpwuEPHR5Fbiz7Hp1JxixGhg+u0N036GPjOaXgay
s+WGlWnPfDoJXQUUHTOSOT/+XGz3PXp/HoKGzgRdosczEw296BTE/9JLk+oY
fnuQ6gunMIZYhRg9xLcstod30tae+TFvSF6+c6IOt3ISrH/pWKTqXi9DbwyK
5W+f1J7z57gsMWtYRY8Pjh2buO2KdB1nqCNg98gcjEHnRuvVfAnKcM3OaOTT
p/cnUixO+vnDOYGZ64j0CR1ao3bWQ3HSVb/80nxAvawozl+V0VjwgZD38rPg
Tj/bTsqMwNf3XApoKQhm0jEA7E4Pq/GRCn/P5/99bAV7sCYORS/5Ox06lwg4
cUIdQLeFQhhoBwDCLtw2l4N498LO3aOUDMX96U+lCHzpeA/9ytUmbsf90DNS
Bs5SoswF5EPUOlLQ+V4EjGkNF5osKySLIOUlxnnplK1iG6lgkYe8/UQujW4f
JQCu59L5qwBGwjFhucrsPLUOUo5EZ6vfCMBqGbftia1sF9eNrM3HiOpd1Tk2
1Ehu8RIlAQNojARXvi7+tz2nQ2Ury+2Om0h7jzcI2aowGO59sW2o5duBos3+
ZJ7TYQe3CC+qE8pCV7RGNYfxgjVNCJ+p/MLOHFE435nW1tCClZMsxZyIZgEt
tZOZe9jmSj4w0zCWHox5+xGrH5FGs5/ZsHQJs+Xrl9d7ipIVHyz1nf/fMdj4
moOjxCtreuuDxwXuEKnCkAjFoF81CsdoTIH0sZ0JY2qPpq9FxCUfhhaGLKJ0
rEqqAZdaotve4955b3BZXYvl1w6pH/rS/8vjDJSG8zh0rQHppKIMEBIcvPUQ
fBe4/ogxeCbM0DFIVvjDz4PQqL7R3z/Sky3ctlRzxgeCGyqu4I7qjWUIRv/f
IF1/HiteajOLxQO4rvgtGYTHz0yOCXoiVrVFdEXrQ3vj0GO9iwxUvfW8519B
eBOVy5IwkJX81v9b/WaSleldhXQiTL+AVL5s108cqwLQNGFSJJi+dMuocn5Y
QxhLDLogGIdc6C/kUzFoVSYL//u1AStO+hhlZKI0ODzxv6lCAGyIQcTFFa7P
PTTLPr47Vw0a1JVQE3O+R2/OYkA/WTKmLNNr9OWsEbUXR3sJxOXPe+b9mw8y
Xz7sctsfmXwS770YBX07ayfmbxcqeENG7KT/IO8qt6XiAA2v3+JZto8OYJOu
iStzP0Rr9lkBmZhh6pAlIJO/Z3WN7R0qpxYMRi9MuiBLC30rjlkP9AzRayYh
Ub3Iq00mx0qz4Fql8qGBhDeOJluVuEUv88SJMWqMfESQKNEghxe89gNolVw6
GLEjFhwqc/aHTduOaWla7KKB7lJG4Z2BggEF3EeLZ8AbOgrfsgv98n48az3c
x/7SBbNqPLqIms6iXUEda/S+IxvEKcLRIzXsQ8Y7Qs1VJKCpru9tZitWWdEY
JWQLf3+bM7TfBbIqeNhQJj6iDjj4hnPWRECnngxrJqManWg7c7JslWzzuuSP
wYJvpUdmTutGpdZuwDoNrdJwjKTttGcALDTFFd/Ne+Q2bPdwEKJzkUDXBLZc
cbTLENNeqLhWwOZHLUDM9N9EJRQJ1HTalMbE7eE3oXNJvW+vJIhj/+VJg+JO
Nm1H4Mv1GOD7NT92Rz2hxFcJwJJMbHB5gWNcZapRDDctYOsYEkJg5VuO6J6K
FzDFRvPI/m7LyRqj7jPXo2KAA+7e8sMGJuC8mRdSwu2ISaQYTlVGmuRFBYmn
mDmJCH8b+kBwFtxiki6LnsJpfHc93EJhhQCHgFS7N9JmCzkKWSYjkN0wtNLW
m3ofrsL0wVoeItNjmseoD9B96bBkSTmT6uvx3IGDunSR1ex+jpCcdJ8PIGPh
kM0ImNYz84taZ89kDeY2MrSGIdlnUZVIx35fUK68fTNQitG7PJprN/+MbyML
m7Pz91Se/4JVex8lyaSq4o8oYt/EDKt8GiX9sKCMtgAFb3iAVtkR9ejYH+ef
YNRzWWnEoTjxPgAn4gpwY8t2pJDfDWw2EwyzXEons2CAOqAjCz5QN63NrBQS
v5PYMVC8ZaeCOtfLzFlFUln+fki8b91Hp5UtZYuoGs6KvJg0tCgRMqJPK6bx
0cIC9KR78zqwk/VXJ1CibB/p4AhYYTQqMefZ0P1u9oeLAdyP8q3aP/9iL16/
YnM+OV3xiQtV/VwO4sqgwOUOouHlpJX4+7zLoMeUV1gUiHqdclpqr/8UqqEm
ZwvOJk6F169/63NVFHth+gOL/mB6PscdvY/ySFd34HztMGHBr4ZLCDLBaVN9
l9EK/JJ5WT90o0C0qpelJ7jg+EF8lVTwWvkaCu9ecyaY1nm/KCmk+Vi2vbVW
LzA2OaNF9ka/qrcmUsLACJ2q4dS2roDQyOnQn/4niJKKa1yGYsxjaL46q38s
M8NJy1/GvsZkM4NygumOkCfijZmnvUBJTkVWoe578hSH2K/tDhD5sTXJ9Lcz
uk503WVG2pMSELZfQnUP7Vb2aQLCh9KUijwCqP9oS1QUrcUFJagx+HeR6kbY
208Cnm+mDgrRALB4l20A2P31QOkMFwq3kG/0x04aNGD6LlrRF40I5DQDOKhh
aUdIz7cg6t4LuHqFzjlPNzyBPa0flSxGkRimhqiC7pxt3/ffcaZ7WqvTXLO9
jhZ3sU1Rb+tUQbc9aWKwFyMz3s4ECIbGyc0KYCDSSesqU0O+hyoVyC9Z9Plc
pC5bnVI/6Uef+A6dE03bGhnDRMLM2Fsw2Zsw6mo0zpj1feV8X3xhaamLlsvI
CplcuhGNmD5a3+pGEByh0AVadikx+pUf75x3Rw7OCExgw0v1Nhc1yAl5kdej
jTxO25eZoF+05j3tjIJ2tUXUGl838BCS/0wGH6Z+uU5STjSeDfNMnCF8dsEO
o+1tVXFAQVkNyzOhVrDuZ4vJRWh0/PfRb+iSkIjwr1yASvPpPISoKDuo4XeY
kDci9vvWGZfd6npHs+xyPyCdhh0M3KlpaccRIf7jCXnGLpCKdLePdTBcTQcI
LhWAEtBVozjuRsfi2FMUIcA8j7NC4JtNZ4OjClHdxRUiHUzSS9+OJBXBaW2Z
WlxPefgTJg62yri6IaXsCilTbkpwaE+tehM2OMHLG+NYZqRBb/Q5KPjxpTnF
sYPDFc4TbFx140BmNF0wgjRhmm3dG2dmlqq1RarBf8n1YkxwEA2Uj4cqQoD+
vB+QzNYLG9u/4rWm8zY5OT1BPvnnOXTJh/O0JcGf+ajwaguAMMH+CDGR6c8i
GBw7rAl7/SbLU5eDvD0IKnT7ZmNW37POfYHk4lGarrb8BX8y1CpFLc9wYhEc
V7RyGgsXgva7/m3gK2RKjq5y1Zdb3gNtvno4ANJxAAhtr3lDjePZCxxV1dkH
j+4cay2ZP6XJgt1DWiHjVwKPno62G/WlKe3l4Cki6BUwoCFdcZvU/oH7j3TG
vMCzEWMo3+eSxshJSlDBPMrlpsU8b6yFiQnuh0K1I//6q7BMHpXRm1t72vCY
2bTJoLQfSBoCrKoco99xyrXyR0msFUGk/kbVom5lHk3CgxO/FzizR6beZPsR
BDO59gaI3zP0wdsr8psq0SJqJ1rFb9PhH9H8350880S+zmjLt8BhLozdukQS
VHFJwTTWHAeC3UjD0bfFzEWrvjULakha7oPXCDZyuvNBEtE+jxLYfg/cDxxJ
e7LjoI0kkzyg6oukCvvAoSxEb40qvHu/u4kjqeKJXE1zqtLSXoPh0vz83tiF
e5H4B6kQaH6fXTWmusDHrJfpFOvwqsNVdWIsmNEPUCpzgqaVHtv99XNSXO9E
IUWqwGl/hWsiJzObl4m+1r+8tA1sMbBELdyGG2H5Dq1gDTyOj7YDOiggJiJE
52KQAcm7zW2i1LlCITypz0cJByXpUbCVnPINzBOGdyyYYGOgcMI3r52nbbe/
vdYZzfDh4oRellO53VlblP2VUwIiHw60WJ1Fx7psMeoi8pngSWskVYHskD7O
t1AP4kWomxgvxlD+IOzkIO5RUTOpcvJvOfQPKCJuL8o2da8YVbaozzx+GILV
/vH0YHg5/0vlSC1ivtWD3TdoKjPkBTQNecM5ezW62v/tkaYYbwtRMUu8WNoP
ylY1KkJAPpeAND/gcYel88QvXs+ojojk8CpDdi2hCvmP25j2LPO/vJbc6TxO
KDt3SwKJnOS8JJ0axKUfVi8ZMgQcHFPStoRc37TC9fup8YA8rSGVZQLWnpEL
mwmYvzJYrRrfmn6Vlq5aaS9gEwW9xKNxsdZOVd26QU8AuweJLiaBlCBrbryU
nX5ZnIjqF1iKhdS9Fmx3gO9jRmIxZMW4J/xtinDmB/3j841OsjUPR84PAfUl
ry+h1gil19hdy4MKvpM0xbpPhHOGzigCpYlowZ1/HIArHAnFGffqmBNbaKQx
QpL24YXFEZWVzuzPgvnrp85pYf0qrxLQPog95hjNXYzpSz0QFwW9Qd+VGIc2
j1OutcjZ98T3BtAtFab70NyS8MlOhsK2AjzpRUKupnuPl+d7WbpZoivtNe0d
JcCSb/FvsYgHzjNAsyG+cWeyX5kOYygybX/RZo56EfAMV0wbBgCQt1NZTqHD
iOrHAsMGny0rd4otnsNXQPPkrLBqhPBL8QhOqqeSl9gxhZk9hYlZIMFwavsh
V2o0T/ZFm+6YqCy6RGLujhFFNKhcL3bO8z9a7yP09Wp2hXgRXn6mKj09pzLf
VQKMjEnZpc3jrBiOLZuCYp8SEQjaKCwzjFIfnbXwVLPJolW1tb3N1tLvA6dI
hkQMEBM8cyUTH56tV0lVIz7FUpJ092aULzFNNK3fanJLDGOTIKshIt0VMSAK
/otZlVxZu4a+zTzLuH8quDykZWvWyQjuQHEu7dqIlzzZO76F4Cd8lRnKIC5d
hZpe+9TZSIONVimgPvYs2BIdOk/Nzl5IfUH1NLryv3IF/GMQ1NJ7l7JsOHCs
nP1otX/J6zahVrxW7RlEMbXGIUdnfysH3JdXJesZ9rlKaqqBa3yGjVCrgy0s
U5OMKJ6RbfkQOqeI4wYHPWoN+LN8SCsiIVd3+FtOGU2DrlxMwJddJO4XUQ19
D1DgpGtsSiH6aHsqBuU64msXBNqfdFZiRJAGg2dkC2u6OgmUY40mMJN+h8GJ
HlFZo+fbSJPowSUsxLWrqoN/p28OfLs/P2NdaD0MfPupC/mW4cxwiIJBkxrI
qvudxRYiA2iTmNSCZzAVZ0L99YnWG2Rav/NH2dqfQyrXr1cU5Ed5J/GohH1g
nKcZ/KYh5tH74XbIgULl5/qCk4kiAv+Ah42QvQ8vnV9f4GWHlFWblIG4ZKsf
B7fEzuSbDiWRW2EPkaK3HhOmOMYJ10K2Ysea9VLVbZKUGc0DY9QQte0ylPEX
99yprfJEWk4bLvBWPspKc6kmVYZ2GP0RWWiniiHWH1Nad9z4uVcE2M515/27
FKt+IZo1d7ycNXofN5rZ0sc7I1dmh9LTxDvUgHcPfhPHf3cTPERa/n0dg96x
IAHtCrquJaI+yuFSDgdjoqXaRThBtZ1OpMHRO5k4rOGjntpHujQJvnuVw3/s
XVccQbliLxzvRFIXRiadRkm9iHDIpd0cKE/iFsnJBEr/kzfENR5AXzTpiFgp
oJXdzO4/IAliAZuT0BJN8sJGAQCbHH890t/FiQH+jQHBrZfOzx+WJc73GC7g
XTLtN/v7cFMe3+UcxeYmnGx3JVGoYHNmrGQ4/ZK13U7s20KP2OUOR53WzIN1
5nIc9yUozr0WdeZ+OnkCEXr562PzOZGkS+IiKOC62CSzuUHV6JgZHeLfSCRm
pFcTmj5xiDXChGaExzUhdpDU7UwFm1fe3GvVqFtEOVaPLQTArVXskRc98pvr
lcQ7oi5cl+syP1hsajpPsVBLWFub8FFb8i7GfuFH6PQl1DI59lBI+bks0gh/
mlmXnH3NGjAQ4F9bWedsdZH4rq3hZItiIKBf6GSUYGSamBFBTyYRcV945o7l
zqmTYiEqFUhcrs1hfE8CLhBJgHVjtVVRKTaO0yW4TTvvTkbP5An/u9ps5jZO
YJ3r8M4Uekx5SQ1vu3S7Laec0uo0WHDrqyzvIOsctocMmDd7+VtsQeoYKsjV
HG0o/EXp8rABFjeavEuuBF4mD6lKka+jUbtGIBsvdkzWARjTFCR4U1kMNgey
KZ2yrRzlpvmFRSV0loN4/w5fVfbDMXJKGWYY2gEBwTrDLDiG5vCLW8uJv/sd
A7sm7S523Gq4Qcfg8RaErHYnodQkOsB15iUFQGUhGIRkMbYStD8+l6b93URV
Z2um1P0W1G2QDikKhpu6fiUdyesAa421DcrWof5xrRXE/Ojm8syylpjIL3eq
7vvZphN2f0Vs83ouES+PKK9pZRpCIRUAff6TfgQZxf4LVpUIZVGY3uhh/2lJ
7D3smFrqUF09V57WbbKx7ennBbdBtpjgLPhcO5VCOw9HPQFteLjlEbRX6KBS
R0o1RaxUnoHL5VXgxE1lDBHOL/af8CL831q2gV2/t1C17ZcfTEfrgRmXs34u
PdGUi45pc5xM5wuYGOp6YIHJDJ1Vue5Da+8YIDj+L5Jn4nVpP8Nxi0w2OIBI
RWMLTqT25pDpKvFA51hOn5U9jX7WcUw0NiCraWCSw5JHeJ9n5ft+ch+02Id7
u6NBBgQj3Om8Pl0WiPEkfh2CtcRjtCO6pfocgRzb8Q/m9sKsYBh4CggoJuaT
pVvaRmkd8flfYDH8RLqf7iy5022mf6Bv12NnA2/5xWbZGQLLmxqFKRJkqnIl
yZ2Dp9m9BAJ7BjbQ4mBdeeeO0eDF6ftIUs+SWPuIEeBLZ9DRqFArlgte1+m/
aAekeZZjtI0qfCa6Iq+cR3eTM9HGYp7rVKgJ4+Ay3p8pSn7mzeZFx2lnMq+9
MNTmznFMVOFAI/FxrTtXnyiTWfSazT4kwG0o96ebpQ3OL6jLK1sqZg4gOaPf
2jGH4Rbv3IUL2wzAtX6GO4KWLmUv5/sOI58pYgdfew6cqVVfedC8MhtfWrjH
8B5FAj6VbcBX+z1a1k+W6D2VmdmsWk+CibnLv6DuXJ7YB6tPBv4Aqts+bs0h
qzx7T+SQTXW5QbDd79Dr85v47v1/U+Dtlk9PiZABY0WXu3jYEdAiUDyoPZbt
yB/JZGFYpulSUo87da5rxXyHTA3tlLu+GlIFWW2ADnqVbxAS3jvAFiYpVSqB
4fEQmfKkPzg2PBtP8qjzMBcMY4YVzCMpQyR5b9HcDZfFZOoBJYuk5bvI/Sgy
UQ/JDw/AvjF433ruXcjZuVm0tBi8JIt1JD9VzvZeUYu2mMJgEG7Ag8cttAdl
g36OhomlFjSeFPqa1pNZ+TDmqxR7qI7k+yF/4GwBOFiDNzW48XKvcg+xxP0a
KMW+VXtjIGkjjNjLKWNKgM2zlG2S4MDPD8/9h/j8BK3U4Q+LguMTRoHPO1b2
fZ75BCbmis1DdKsn9A9iZStl+HO2g3wmMVeR80XKyEBlnyhJovffEclTnnS7
Kh9P2HXP7ixHxYdn7oElPtazJKQu5ti02nVseCpFRQ7JHtLbtftDB+8JKydx
QW6Jt6rNRv4Vil0bX62LiI9N+xiO3d0I2uIJIZu9yoG5j4oxafjcoSaRK4hG
06TyZNrLHBYzY9RBLWkSNN0a3Q5CxKIRmYnsyBSefcV00aOd6YCSRsc/E4xE
mVgZBq2X8cJ2hUPMAdvNz9Mlw2fYoA3oxixRKek/CTLH9F5vmPkbJmpiE/4a
+Wiq2j3HLEdmpzcPxNG9YFtwM3IueR+TGZNe78uUw3Mu2oKCpmJL/1Z/EJ35
3hXniBK71Ipvn6WNn61Y3xJMV7ZTQqUQa2ggHyzBN2XUwC1GWtM7MNVhPOlS
NkOpR1gluvWQhN+nKgMFbaOURagpKXFEWu8BxwlVEhyTNUCTIoAEU7FpuNTR
NVq++TdGiPnWRVOak2qMKytITQJAsZsdGdpC2f4r1n8niPdPYvwyjZnwnpUX
/pr9iWpZW3zjo5w0xEplGRIG3TiPPUC3RlkYcrNzWwSi8/DmUSAGBBEKv71c
TUvhId66DHHm4gkSNCuQy++hW+Xlj7mEUoN7t5JludJLIlgGBi2bCF3E85hK
nBd5mU7IZKON63PtWIUCtmnwaMr9KDAzpo2vNCiOQ149aa3ZC8j4dM1O66u0
b0wF1P9/JZUpZzS52LkFkUcBA86g4JXb2P65HnQd0o+v2xrjnpQjE8rc/kmF
ygmlCsp7l563IO7XRW+FRx8yYPhb+wJ8T3FnBROksA53/mXRHLopq67JWip8
JZcF4mqduhKdwKzAWZ1jWAd8V6EiIWbWQnQ6n9vLt1lrcB7En+Ida1O2H2k3
OVwN6eSQUkjofKTmKqBwYIk+bnqYB3wTcrEUqxmKtrtPhS22AfyJNDOY5XD6
zKdeZTfjGB25yKtStKo04m3RWcv1gllshBCJ52EQTR1TFvtdYxnz4W+S6ht8
eqzkiRBZwcmtyHt/vxD8n0eW3dzq87DYAAVdBTqfMmS5UFXNJIivCJSiXqC7
uEuB2i9znHG0fcmC+XwSE7mCea1Qvqc6KgBU5rrgNoshGPo2X5c17AHAWz5k
LdGV6cCgOHNfW/zRXmTF0FHvKiP/hBtwUsPpVAf4MaCSwwi5Xhfajim9Wey/
5ZYw0wmf+4++6heo0nJZ87g+JHGxyL3QmdmLkEYNnyxbxAsz2IJ0ZU/L0i3b
CwFGxMxM4E8PmFXWyuHGxJeC/RvYQOjhVa7S8LKalto8XWOevQTdE5ITpztq
1BSm81hmLbTNap19RunsZHnllW+cnSIwjto2PGTbhMTwAMPdo6ICwQX/WA3D
ZP08ar6uPcBRK0jm8E7lyHvnhjKiLelCOJpy2MgWqXkQ5kZKC5y+WiHH9pV8
NtpyBnBvUgRHIv2ukZ5eATt8gHmuBXEJF8FrbEqm9ptDs3zQW9iT+kO3Zi5S
arPQYlZmdFI1k/URn5YSrWo2VZBq2muTqcNW2qBR18RTXenjs3reTNQ8Haiw
e6JjRWTESo1QfZR4ptA9WWaYaRa8ZLe00jQna/ldOPOmHr1fo9wO45DSRkpJ
OrSMmjsQWRUsaa3j/06Nk4ciGDVzZ9w5vNWU3UE52igvsCyWlLoxepXRzL/3
7pQ7xTCGDByt036ECUHaOiJiFQyyXjUQeTfz0+7pho7uSLdzw4DiqTPzLO4C
6RBfUD3pAn90O4KCF5zUOf5DgwLr863zVTLZNn4mzqQtF38e9fE2V81+6HnC
QvssnPloymJXxj0JWPPXhQ6igcX2+ZNvmufCpoV/miHoavmUv8c+0GAJczMK
suOJyM67FNwx84SR4EYuDM0cis9X6Iu95dYp1lqpfDkFjm73sUu2vfkrGddT
RmZnpSu8TwGCHweBhO6U8zUPTcbrYvkrTdUJvIYwpmmjjY6a7RSLNt7nfKie
QlqrIRdPKm8nu2VBp87G9CSsOZKWSUvfyI8Be+cCBlX+4g+XZR1FSBAvgfiJ
9DTzmZU2aRywQ00fUMolDP+P2ZAr5XAXmhJc2dnz6TJ0Tc9kIlr+/jLzFLH8
1Yx0K7fhOuP0OBoRkLpObfkL+Hs+dFRJmxsvshxLULOANDxUSQa8akZHyPOL
oQWJTfo4PmjSALtd3BZBLQRbAbie88brBkereUi0I7IGK0onL+PHq8w3d3VP
PSam+dbN5qtaQvkTpZiiVyiwvrWGB5iYidUs5RgH5f2BRL4O3xruywZSZ+9a
RQN3hGRg7ChAVDUQgX+sikKfE0x1+V34tUSmP9YN7IDcbF+Am8vxYyw0ZHuS
cd8hHhOUOu037RVtL8OpJ+zD0OD4+LGkBrsPZJziiKPBtxmcRDhJ4fztFc2d
HgvnBhDFvEXx3NVF7B75gVOVZVkibnQsEkoW/X7UtuQj5+tLLi5yKFlwSh2o
+G+nPa68HI9R3qYZ5RXwozlwNm4Xuvu6JhHmYhIZokyaLa1mtvZxRoRukgaa
sLrJPXrYr2Zst2Y/VNxCOevZ1WHBv7eD9gNjOp82eDHAmddCr9M/ChYAR+pd
UsyLtE2QbXjOVGZ9FSyfV5omxDhfnizjhgwIxqnCBFVIcwdbspnHzLCQ47cg
ck1qXG3Ws2eJd86V6hWzhtMZpqKezMcYKi4DWpTLmZ7PPYcWTKIhXpfy5TCy
2gQ4+DPsrJ6uXFQbhXxEIlAiDwR/c6BDJtg9r6+FwTwUbfKvv4HZVXkHwdnZ
vEkexYlxvky+noeVLMFFCjMK1TBRv58EkNcSnSsETcFJ09H0wgh7Y4ToQLCG
R0zXKAftgDX9PAtlGSS1lhLS98hBa+PusvsEOex1puw3m92+n+n2jEQp4cuc
GM9wFbqeiVgCuKmZCkNNuZwgCbh/ARTOpxrfumxjAOuVRWW5g7XyiPMLplt1
zT/9+EmSxJqnCKKgqouk2wUZWSAepA5F10rdJ8CsuROOcXmMU2rmZlRvp72U
ixGLwmcVEnOzoInTnWV+wP5gdiMZJanDcIx6L9I/mysXtEXzZvw8sBX+S7q7
z01c+gc3N48dawFxf071Do1NAg2IO98QIK0HiKIC2iGfHV9iLGDz62L6pbhB
gkZDzzzEBfFi/v+2KIuDhq04KdEuyGO+Fm5Cch5AVQf+lGTGRgeqyyLmwZcd
KdRT7kqxAmQu6V0piTgxNeRibYKZ6q4vvtRCQYooxrYgMiAkWy4gs+0NPvlV
sJfCADw+M+KvDcKzcn8SINjQM6zR9MkbJO3NXlcV8qSXv5+Z2CHErywRcD7U
pApQACy7oVtVFLBDcLoEclwI5VIX6RMhjS3xUHehHIWneKfmMmalBi702VXZ
AqYejiKMF6p87jT+YwFpKsDzObOxhen9G0/GM9v5v3P7OMYrDriF4v/woqEb
AsTeKOzQqGvnas7kc2SqDDgdz0iq/JVmhL7ARSpTzmV2M8muoEiENjLoTfOS
7Kvid9Cxeuip0gKIYGuidlPhPRjAXrDrjnGfRN4hX0im1Q3bauJTjjxKbSMM
CNItYv5/keZrzvDaqbTQEwkQcsl/5Mz6NlkSd7g60UQ8qhduBdEHCB4KDyYX
S05i396jLli8i84YE4TRdn20+aT7lkRt3i7jNuYZJWXQaZwC8VJ/FHQUCkbS
1a0kAryhXjJx95rX6FOxvXAAVCDH4Rlbkc7hl7AGPuYjKx5t8krKWd3zbTik
WX78ybDkS6bprin7qeH06f3+A7uDZRkn5fza1dJcwTzHoA/1Lkfk34+FtMIg
8DhiGHCxwFWvg1ERAX2NZTNPh3tz7gIz7gZMLmzlAtagIfj5BJlt5KYtw7fo
jj89NTi95R29GyYuB8AhESpzywJXwgYJjlIv3paerzK3HXaA2gzjB5Lg57NG
2NsY/BWR0I49LLqJfbxxXziFE/kwpbgXcY0s+YZDyGjTLuBSHWzDb5G3oj/W
XVXJBFDhwk2uExlc5eJRVZ7lxclsxO6bgBqpUyRVlylO8ZLwoDsoTzu97AHB
mjdnOnUnNA7bejLqOY0WHuCkMKADi16HLr1ahL+vK1ZsGvXn8hXoQDLREf1D
XiaJMaEKe63NzgwAQv/c4EWQM/p1tIYzpwOSWciSQtytsoOTvwp9L2Sd9VOk
vHoia7LWT1BMUD99dMQVZ6wxfLj7tq11Ofvn7EQ568g+MsQK2/Xv+z5XFMuC
3TBxD9lnas/2eTVf+oVZaUeFj0Pm2bz3JmmnWNI6vHld+rainVhicFY6FVKp
it2GmsdvUL2Kh/WCwRCppwho961yYO2CzdNY+1J8Xg1fohUd0cLqE8wYmqcv
+qGaUs9m55gEz29/IcvM09zYtcnZzDiGnBg8+nfP96MX/2pOuwQD2H2y/W90
Ezels0or/wSamgSloycykmkNzrYLmrUVxoZ9EsXlNutxIVmzW2o5sKHEAcxH
D1lSWgBRP+WmWXL3LmWMPpGTsW1cfSAOhHklCjspbNfz5LZcFFShrTSbEnT5
3LGQX+In+h0YbesVGVQDoNa+82yeCipu7/7SHTEyRp00DoAf/O2ahj9REyrl
bJvVvLPHCdS3lENmfE13kjwT/Jur1IaDlLFeWQEWiebfTBVHc7UVfoLMj7IW
ScApYBbftDqW4xbmll5YreEcgYWAJYRN5dJzlrDeDevT4+aac0r9XVVLeQxx
faJJREMIWQUY4nFZGwp0SKKelwVi7yYSPvQsF9eijHfa8KsDrjXw1evF3qi+
OGBXqGhRKycIAL5I8aFN4zsaa5wJ7vTgENd8Mrdh7INjQIRC+8c2HEsT53MR
Mpa3YtM1g7Q6FBUmaTfrhwWBE5RyDTTTLnB19od4ytNSaY29+VnzRKLvUypS
qbS1sCT0hAK0bwV88DVUWklOSfiUwrr707kn1ps3u74PN7nDyDhebNMWu2LS
0nDUWd2uLYgW1R3yoraP21iu9e5bB6kFK08nExBxjJ6vH3Iewkc4m12W0jRQ
VNLeSqEjib8HXfbYgLTR6Yeg53gfRDt96SjNAHwXvQx4QRU0/9vTguQzL8zW
HGCpgDe6FXIdpeVXYxBW9OZnh60aZsBmQbePSWggjevO4KK36j8ElAeSD5uz
EwlJlMpyVvpdX4d8N4wDRNfDva38CVSUDhy0gaYsk79+EnqT3VinfeSuQ16U
dimUKLlPS4bms/kwmw5I0UmlGAQGFoeROgm5tnTAEaEJkCfyL7CnNlZeP27O
kE5lim4zzcz0y7ydmBL6qyRq/u2FQ8vkUKoDVDpvBwOxlOopQkpjmu2G+H0v
/Afafbp4oHSzU2Z8z8OGjaPr7z2vIfKuaJyg2g4UyISHjaHZ7qxCksvVDi+3
prjcIkmKNt0fXZ82eyWHZkj52KJNylumR2Dts9CElNbUwkUA9m7/klWmgJ3X
1FqRsOIjml5uobV6A3OpOxdqF1r7GzXJ6izfq7zOoCryBbpYf6FcMm8WN9Zb
t2pnmcyu4GaZ6ACjkn7Aiq5N/90hCrKpkEplB2w9/yc/jprwnjkpKsNuMftn
PKUSsDxUjLd0t2cQTy+5YIWmPdxR/bz5zuPk3nIz6pJ3exTcDwZS6jwopUKi
U+SROx+Ro8x+EnivfSgJMhFzx/FRyFHwxlscUDbOuslxsGSCOvnaiVaA5Q9U
tDnE6BU3/pxancb+wqC/DPv9c4dd7eBsi73jgb4QbczozCvO8taByOHRvpEi
FLWqoH/u2grPya72RH1e+A+8Hwk5Syc/o2970A7x7uOvABPNrMQl33469evH
/8kge8X4wQODIV9XHBVq6dRi+/tF005pcb1HCguHtlpHNj76DNbP7wHB4g3F
GP6mS163j8qsgSKQjZ/BAKdAbuPBQvw1xOSH3fT9sv2nRVVn5COVHzy6LHUt
BFRDJkcgrel9LozdiSu2TmIvau2iXUY6jzdFrDwHGeYcpQcp2pX4JVsrtYoV
waTogbUAsnWygHBhMvcR7y+K4px6lK14Y2izKWPNXPLhae8UUWc18Uo5AMax
GPV0d9c7QJiQNDUgPUCj2HZw6nONY/sEfx0WcAdR3iWxquPlKNuitqQRoX8z
ZVKE2Sd/RZAd9IlaLVwSMq/ug5Dd7QFHMXJS2paBoPhvpMd7P67Tk0oqhNyA
LW7pRnW29Hb87YO87vFoJs22HylN8i8Z9ir5z0uRjUNQLf3GPL8h6e6fp567
mwRI0daP665lJTky8tAR+oiLFNtmpO3Ciru6qvXTE5Ejk4/K+HfpQv8i5Bgp
k/Yx0l8ZIj1+0raTe2ULOmh1MsLTLOAuRARUWUCL3mUdbcS9bqur7eWYko6V
DxIdFpa9V6HYoAHKyAD978pXU3hnj7MfmyPtzEEEHK0VdMPAxSrOo/w/seZh
fPeIp8+kw1sjNt7JUzElIiB5JuO/gBTwlUenAPlle7dztKSqXWf8uDo8K3qV
f6MRUetszmFks7nl2QTry4+kaO1cEBnVGhPcRTDkLrKggjWV9R2MiIrQFcPM
OLp686DQZwO756qWb3ehcixIoQlKIUdWawX7kpyDVXElYjDetgCspdWXER/i
tWF6pn1lXsFb3exAbHF61FzZdVA1LBLol00ksqSmxl8arqAYuXWkRYsVpTTf
URFh5ELYhQ3fdmdxuFMGno5bd4Qik1a8QW9/6hfG60PObbCxlzAV5iRNXEgm
gQAGeTrbU4zONe5+1O5yb481geeyv5jR8qqrlKoTin5HvpPq51ZIpXrQKL7H
y1vb5IrnYi1C2+MMtL+Hz61sOIU32vc+UUItBSYU2ZwiyQCzTZ+xZW8BCObS
tHdMKYgs0GQwq4XJJAU9qO/NjQ2SEPPNgeKWY04zaUa7Qtft0jWqfQuGmpZ7
Z/C23SaZjZMSaoCF4lwxmQ9iKIZ4+6viHUrU1n931qzqucMoliA6+IdHjpcq
r1kqEXd/dtsJ8FZ+uaoAYR8Mcl4RbXjrIjvwHeeb2AdyJRUZm7S4EQp7Prlu
G8JgAbSf83Wp7BH8LPOOdFZDFeQI1aWLiSevp/PjZv0VjbDpbls3zcVUTR1d
sSha1N22euLqQrSstdnpy6qbCKY1TE3faopjTWG8EtntM33nh18Y0BOOAXHz
mq7o3fM8jISAd1y/j0rInJtf2ruP48ZSLZqbmpoojQ5Y3Y/SEZpHI40GrRNO
oS2LhuvyD1zq/U7xOa2xmstXKcAFcLhfBrZxnGxd7gHPA6wVIhXdkJ/Z1k/8
a36idQHB1qRTyI0f7RNC1rqUYi3d6Kmv+UxdwoHN/P7UWnm19E+QZsibg1Q6
z4fZCKnvQOIKmBUFu/9hYHD25s4RDSoO6LWyDy8SNDHJkjfpFhjZIG/jJy8+
Llhcbtya/cn8snuogelTHifiuxCO7nzV8WaNgjQPzlMstw/CLP4UbZCXZW8/
eRX1akqi5X0wxkcSZDP5VZGCcHtSqUFgPwZVVfedfg66ebqMfRJMmroZqw2V
KGcCEyGu1sPZiu59HSd6c/hCgvnMMhYrM5VjSsFxNI8rHe10q01z9Ni8M3zr
FGTYzPqD+EzdgqmsZ8cbEGL4kX276Gkiei7/jSGHyADtkyV3P1wZ37Q825e+
elPrFhxSeNKUEp5eOW8gyHlE7HAStgKuBQWMQEIo1Uc1Zt3doeOGGl4ium22
7Exwk4XW94EppfTF+aMZfshDvay+gOjcAWt0RtGIPMk0N/f2z0FTY0b4wjFf
e57lPMS4pzwI7ZbtCg3RYiS1oYzHZLFkfPhJyiabFWetVXKkdl/LwyEcjsZu
J/VbdfZTeincLdpuXJQe6gjTSmz83BKRyO3JmvWW1QI/l5PNdzWaTrEuSRPE
ZyrqBdTs3mc7qunlambMlch/MM/g5KPhDY/629KwW58oaj8UqY1zVvD9E5Nw
sr7FdbvQ4BQQaDcFy7dmpH5L6qJU0ulIn/AduhxyMAYEKzat+3buzKaRnuRY
IcCWWs/yfSWszfpofOtRKLH2tdQURwJpMCnZDjEliK9OQXipFAyT4Np6Lpvr
xH+aC7MhVYZvuveYla6Br63y0dlZzqM0h8I3Z68O+xwGJmxtbPKxLA4iL7Ls
i5DjRYx1PbyFnqIvmfWdasb+PRVnTogGlLyYR0KSiG6ph5+KWEU6GtwJEaIl
74vZvHGi5+dIVckDs0++S6Qk80EuTETZMjMorAFH/JhmnFwh6NLwOJvOc/Gb
7uhcsixgzUv45qjmLQur88LDnZwTdAuXKMMivsIGMuimi8J/R+G1U/KkkQtP
EgIDpvp5StAwMoUfXrnFMX1LKpnlGKGOzh/7wGMn5kJSbc2t5L/i9S94Fum2
01FW24/ZbvUT+rDx+nZFj2fS1gADDSJ3Yc/RIRKiNRfYeHIxk5lYCovOYzKb
X2fv8e+wU5x9f0gHXcbZPtgPSkG1uyumYH2ReRN/a9lfcrO8eAlIBtecbNhg
JMmOrPVJtL+oGm35RPodDycWgnTnYGcS8L3eNTarKGvH6Jv4vR1Du+mYzWG8
9lTvvuYfIDouXf/q+H7j4DEqoT7VctMVAGV4cA8xr4QBBhDxJJ9pr7LrpJo4
oCxs7Wd1I6fXheeJ00wSCI9/ED5djKYdj1BoYrYeDg4ElNyF8iecooe7kB4l
AyXF0fE639LMmQnBZAbUC7I/GAtrrXpVoAcESV9az404TiNecGjRau46L5SA
bClxzruD/Z2MZ3rI1B0C7Dxts+0ppUv+dvzsDYrxEKsIsvAyvpnK+44tYMKo
I0S0uSpJQoVBjcw4vqCBoNjNhzlEC1mipxwDcmn9ZIHYfXIwpm2riaGdxIQJ
GKsnpPJQ/6XZ6ZsYloqP5Sc0EwDFFdK6WlY2bOeg/UUaHPgNHlqtwV3ORhLu
YnOO0IymXWzrdWtSd0EwhYzEx73s2cRWEXAWsAO76XhpSNx4LmldeYbmGL0u
4PjYArvrLaSDwImQc46b0UAx+fbC1OudVi8kk4/lnqUCRFc649PwwhfZ7lyH
ls7gzgHOpqtq3j8Lw0/xSQnODsU1fFQDIMg24KcMeUNcnOzVmeDg0BmtFmF2
VXNJHr6WbuvCsuIdM1d3IIJpeghBm7K3I08/gVLp3SioMi4XqUmhupiPXnQ1
9JwA1EqjxyC98+HGRu5FY8ycWabitOAwVdnIR8XFzRZADD/Nti8Xs7QNOU3O
GG4i2IdXExQMzs6XRi9gTXibPy6AxdMQYMsQ6ea2aSjEC8vyl3f8R4g+raJ4
iPW0dXWC2ikRj+lZlHuKWkxWMiTE0RZCSm11hoVGYRNBvX0KrTNG5NbHtGQm
VMs4XIq4pL/rWGJaZaGBtOXwEKkdTWwCfCdROIHPPLkMiDSYWrLgocSbTs84
Kf2/kyKmoccKa+EtyCMQd3dGhdBXTfBXsMc/GuoDK7JNORUeKDZNl6ZO6LBD
tGzrGbK6fILqgcUkTM2eV6gDU/HSsbBsm84raS4MfqLUHg2VSdvz15T7xnsz
l/gIQJSHzY2HANhpUDjQ43aTlFIYHR/xiABc3+BMUeaXchVFXqyavKUV0G+0
5js8uurl5TWHjB4iaqZzyZb7+MSE0891Q+O4YOiob/gVyuR+H4YATSiMaqpV
6F3lwUl8PgLxgp5WKZNeT6Fl8l9jLydkCtM9jcsYfBkQSBEq16iaBK7DUZQu
09L+B5aU53gZjoxzDloAL2t570beC5K+tElv988Ks+NvQ3B6lwrpaQeZg+XJ
kv6GzNBDbb+n1yHr322tCOO5zhF26v7ujjFMmbPcOzFarv1silXL1uBYqIty
uw+Z1KmBVSsyZH7nJpgtLJZGPDDVF8mAYAdyvLImpsRSJ4mxklXKQlDOuHlD
/mhnrYf4cwLoDK56SLgzBjbfD+Y4AjHQcy6hodHSnLRsE1l68THhBmvENGR/
f/fG1fIPcDJ4zvVk9vvXUSgq1noHIIp+TTKHbgJ30+WcCFsaIL6bHYqwnkDB
PMhFNRd63Urq3DyFrwhUqvG8fgQlpOcBUtUrhQ3HAZIV89UptNdGy0l8ipD8
GdP3/REtoq7uo46PcZm8lyg9l63Gt7RJh4VhgzdQ/caDjAOgnJe2BEsgWb2a
EfKCiukBdfklCQB6HozVww3h8Vt5nEPhue/910WhGY1a7OOyw7Pj2Kh+FEek
G0tub3MAsJ/7SKErRFH/efTPlc5yln3hlmHoV8+yf/3P48beiZ1eGg+G7YTC
cY/O5bSE4viMV5kZo1rcE5poxZ2/KwqwCiMUYhCkV6TTWoRuMMXg/QAI7Yk6
lYczfYKNL4NjkamLxpMZLWHHqJ1sxY4n8Sv+JZeq9iYnrcrjxw3IH8eFgGU5
EF1hXKi7T509Tgc3sEryWG1RYQnPmpd/CE7Y7w+bL2GBzGacI2N7jrIbhODE
+ar/2xTJjDVfO1OdaYIZtmUyewOnCmeqwlStd3rbS+AtkgnESX3wPUUhS8/J
vjE+ocP91LohSbQTxWqhWLlwpuTAdHgcxTlGcNGlOJfHhkFDudYY9u5mQguQ
d+TbDf1M4PUPYavdHsnNiOl3HFFV9jqssYgyH3eSKdXIeZVYh/BTKhhTxHwp
nPz6Uy+rQ/ywqSn/jKT1ICcXUM71t9C6fxItY8Rvj1aP7Ie19uwkoswqKn6j
owjBwmODW6TV6JEkSlONTAMLCBt59T6ARG3X7hnCiUO/AK7Q1HJefTie2kOO
DCziEd4BllgbmxgR9C5yaaOR7Gmz+9a5z4PIP68g0SUidYOVe8DBzZNCa1dg
s1TJiaRPBecFVe2qyaeZDvf/j0kUR878GZ0XXPCTs7/Jf3U9JxrL/iakegIv
0klKvmI3KYHF+8JtEABoob0YC1vhvK29AEXvDYCMyA/YaLJ7B2WSAM+R3TSW
zFDc+GD3SPno+JU3cIkFXlVEEGKI316y+Rx1Igl3c9fbFIF/zdt+uSywu91Y
T/3bLpO9OQeePAgxdaxaoiUNfxIsKRVyEMVvB48biDHW8JwqdsD0jeIsrRs5
uoWU3yFrM7+icHr023n4SmNYTtMg3m5JJb55fGLMZmROLd5uXKN/TjqtW5Pi
2suhyuB+0V7SUNqpzJMxNmf8o7/2yL2EAofC4gV7uXeip/4JnM5QXcdbB4N4
FYJR01NxUtqw+5NKUXzUJ/V4KIe1ea2CGlNMzn9dYo+YAyFxTFGQ//Fpofrx
LTtknHeIt6dws23CA76stb6rt3ZnPdgIcrTpcY6LArmq6luBFPyVMzI/7ddh
otwEHF/gEfgqZ14tt4tHjpXj7Ay+453jvCqYiEBOPzfWklxNfhTm75+1Leh+
sK/z7rvd0z89+AUzJQ0kqJKWa9hNEi06kkyrI+ehV+rh5fA5sxnkST9QmZuW
gHPH9Bpd3AVBd1fcE91Y1ePL0jH5GR0TUmzjjNiTQEGa1bnDPgK125eYDyRx
jL5BkGXSDG9g4LTSMW+q1F4eRSytbeVrEptbsDBN/AhLoCqc0G7aqMyESlKv
DY5CWBBEM68aX5tsyHBQuqROT40m+YKGtcyHyngyzcSeSOAvh+M3OyWFUYUp
PqEstLVJETHV6EDl8tFQ3RH/3axJqKz36RtchzThFd9VPavR0uRp1kk9LfRu
yxQ+kMzCGkKQsebvxVW9k2GBS1ETkbvyMg6ou4BbnClwPRUeOC51HQirB81/
ti52fT5RPovsewpclaW8Fz+j4vHh/EQVelgUPzsOrLtY9yLuob0ibPlqEu21
rmi8Wu9+3vDwCO4+4atc8TeEE7MBdWq2Jeg5Z8k8vPhqRLhokZRZEzXqUi+G
KYIybpIHPTJZdZmTUeqyccheKC5Bna5oYbLYSHX7JViRTR056lA5FgFq001Q
KTbzbnMHs6qttTPKvLJSTBwhjJQqhHreV6nLfC08oThQg3qsrjMAQ83krXk2
zWrpWuT/Ua1iKHFmumo1/pbUgEgt8TqwnVPvD7ImkKwkrxk3eq6lIgkKWHfj
EP6H0+mYFWt5l+bCUJMir/TpSBU2NZGarMZSD5NtYSuQ7d6Z/H970zuyYmLA
xV3su0Ikt2QBCj2kq5DOe70xx8zOvKV7BpuMuhtg8JS0q/vh54pY0ZwJnXKD
0Azs+emVHe/8Y/iVaqryf2xv69A8bmoJBOFQdztCk396QGX0KEVz6XIpnPOV
WRJPo4Z/jvr6n+PddbHgjW/ud3bmv4eNPY+CviK2zZNECT8QHMax/+8ELwxG
DQ78XT8ZRnns9nuQrJA4fy6zlSUAYSilGeFyxRMsf27MUqZcp14EBYJlLaSR
KCXrH5ancb+Fbn3+JfFVtEctQNTyeG01I/CL0iu5EXjeUHthxax/a/N7g/3u
1PjZ+32Or9xnw53uK89UZcghaSrUZ3SBfS/IcxV+Z17E905oB9gAwUIFXb8E
bWOICndVOkhKQdPhp2CtEPsD9WTyK+xNK2egPTXcClT8+mkXsj/MLFTz8y78
6Yp0frmv95K3wRr0wuY6IPrdKlRXOPiuYeZ46zYk5FsoY77LCWfU9ceGzguI
RnEBl7v2Z6CuQFAHALjr7kNUfrv1frXmgRYoqcFi0E01LPEa+WDmYC3O9/Th
gcB3QwRj6EPJIVTrvlrb6DyEMY1XVte3ZZjehewhLQIvbxY5gAyu6O6D59bj
XCUiVo5HCp9EKh3lzUri4iE/6OntguWTNOsHBWBNQFMvy6kFkSOkgJ0wE6NG
zTHESNjA9vY9D964ZYwTPW6fyV5IaohPqCbShgjK6LpJpb0SzDGWleuxcxWr
giCsQWpJTQhdTAW2q5C5nGO8ZR+Zj22dXuqztTqmIRIH7N5qocZPbTcWnNwe
M0b8dY+6BCm88XLcqQ+loQ9E3WrkV8YADtmn+S43O/MMuWqjDrN6926xUVZw
5M8FGGWnJI9xMBES1oEwQU1xZiTd5iUlDM8vrj/Zx/cgrGbMizV1akmRXdR/
kEJwkRUANVZ981GCxQBOiftZ7lrxDarSflIF0zKa1kczWSkICbNeKuObbHiB
5lyHlldg1n8mMpzsazN5Q8fJ4sV2kRy7ZHItMnosAdTR51Jp6RLZA5EK3WDs
rd/a9SZYiwFjnHQjWnSV0c0wwpwSNCU5+uyzsmJCdU5iXFDp8Qinoe0WNaBn
qQMzF+btKAUpc6GkMZAloY++d4rX0GLarCYWIFHAVoITSae0jep1NF6w5VQb
AdBxdJZhImqa6poVUDDJ8F7RKWIVBvWPsXUuqEx+4nt2KNvLAT3DDrWOptIq
rQV2gV8c5mMMSP4pFjyWzwKvsJoNlp2RvxTgTbTS2kFL3heSqocQw6uDkWvg
HieJLSmXUkc+3Mp66vgcrC6GxJVP+yyNqR1yMY8c9wlGy7z7wAFCJrf993/k
sWk54/N3OlinVyt841xQIxa+Duzg5TH2OWT4W7PzOKvjDEoUBSotl0u7K7e8
BcSGhnwJE7xGm57DGjyNsOgG/l0h+kB+jL/4zX5KJIQ9krPAHg8fyd/AjSFc
oH6ih6ikFmlOezQofNuuqNiu5vPz8u8y4+dnefm0htsQDSF51winkRjyS3L0
Q1r5h04oJW46uQqpN+koOyUrr+mAlUaeGhATcI3XXY54S7EdeRroH4LFDJzw
StIJsh1YYl0b/7iXtu7yRAZL8u5Vffrl04W26+jydayAY5ScOw2OTh3yGIac
3lRiD8uUEAMbh8P0QEIB/OsYeLMjcRxlWuRTucDq3iLbmZC3zCYMmE37BXzP
rIIPJ7zehoDN+MCYCWO7MeFksW8lW8bF6t8rIfjxY0L48YASBtzshBdokI68
fxJ23uwFKG+7PcoAoJsUchPqO/3MGSh3Cnw0B7fzQJ4ouepTlCSLYFmjurQL
h7H5DWW3eB5q4dMTXLnolfMvomCQ65ZW6F8qC34w0iuwHsW07m8aaa4vEK/Z
jBUihH2IXP7eZ/VBoT0FpPhitWymwKIIpPinWjFUbTyt3jg2MlfGk9DIlcr4
EitEirnEJQmvMkvK7UL3Gjk29XZeiBRaduO/1z4EhAzyyBdpmZKwQT718FIU
JxNm5iLo42KSUsnhhwMui5t6sEpDITEhOxlRXXIvwMHw3Nzk/pOlk6EJL7vI
LnndAHSOI6UQTw39LbXP0pzhN2lDUr3Q77FruwGGRatbjgwdnnB4+UkJ51Am
VvyyueJENKj+QY4FFdy7E5GiO8+hyoAgarwcPuo+uL81CKXOiVF+8wonb+CP
3/1PaY/Xv2bne4slkm33PShXrPt5pn4Dv7vUN1Ds/AJ27TA0Q0jgQm6rpWc6
q+ly6VixU0h7H0ojsm0GaA1GIkKenbPnBYG3FC6Na7EHEooJKf+HIWLVNmbl
J4m2Hvbwy60mOhvULD2j+qHOrMWzj7NljP0/fhk94k0Ux5B9UR//joXQFYmM
xXbCLK5OkMumkFH58KmQpkxeQYyAGOl39CElcRTY84N4bdUwibOinYArXxdi
dkAV8Z5j608c4sUyoUbiFb8++Aa0yP8Z9zTfjuKVY1Nz7oyNG7nyoGWq0rke
/Z8ud4elDq9VzlPB6hDHoZkYLtNjZuGO7pVCp/jIhfN7W3eYs40QP0EZlu9d
d2zN0P69Kz3EzGsA/ilNzTG5Y4oW2L+IGxzhKSwnc/DCQQTXHE8m6Rb0d0ep
e/3k3Oh9frjw3LENQCBQ5AiOrW6vO96NTIW5J40FQmX/iDZ4ekRQL2gbXu6b
0xwjOh+y5+fA0pG0aHUpNnd9BJ4bCImcT0e8+RMH7VZUcPdSOsrNMm7nht1v
lydod4egvLHHcHm3EsM3mdJwNizK/T/ObESe0dzQhgo2+WEIaHMUQyCDt6Wd
TJJE3lt5QUBMqWta1GxntrXQYRDKjkdeSOAaLH8+K8CqHp1l3Lt7QxAAFmaT
29J06Z8GWG1CNlH80CcG0XzRzGYOQi1vvo2Rn8VdaGWspskfppmsPF6cfOpS
F1ZxupcXOlPi4hHsYNV7487q9E5sXC119v0VlgoeOY9RxvOg40aEo6hD2kgc
6HiL8cG/9dS7rLpZQOIoVNXFAqJA8GrKs07YguTQKQHKO0o45wjfHAivvA5c
Ah94uYHongMNLXLEis35rcQcsEoz1sLTK9DlNOqPJZE3qcp2aUk/lbmdDLKj
pibQ+6/JMfElwiaaPtU3S83+cRWw0u5TN0J461JQQoQBGi+L8n67d4HQwqhd
M8n8wbFN0N1X+O2BxPxJqIrzrum7s/iCxzK2oAhVaNmG9zvjqfGsg7vDiTmD
VdhQMyetocaUGpvr85t2/Wd7CV8ICc06N7U4PbR7+RXA45ATzIrA1iuoX/xR
Nw0xfGd66w1hUYKNWcVMU2KzeXeiogAbfwNu59BoG14mcQ1RDphmtyksZMSE
N8/2eUaXyAyCMi+sYM+h8FjrgA+4zyz6NZwvbV5VKihX1XqkQpReXkEVJEPp
zJE2K03Wv3jPwkElcCszYkIKguvph+d/hRjTkMNWsXKYG1rWrJgwsXob1mK7
m3/u0++RSk3vS8rZg7mhmfjxdR+tua+WNjktvwY3Up2xMESEgKqhvjcXlOhD
bbxaZASINe19EII+RxGjoFX05CjvjJwhihJ7Rbj+bc1YVljI22jxYrTJxf+M
KR0xztiR3T0uM3llGYgxmip0MiMMaLtKp13GMUhoRs2HZnyNdeA+K/2IXumz
kjNmDlfz/MS+WMaDsIxM1uNEK+qwcBMk4ysZpRMa+xXKsryf45A2S4bvZtR4
leQaFVGDUps/8H9nj70U2DMBMrMm0iL/rGqFLefnZKoJFNd2mcHQKnkeUaEB
tPbb/ExTTotS+WYOU4hiCtRrtVIyGF2sdTPehsgJHqjS6GXNQHhvZmJPH6ff
IqbpUf8f9JLlBWD3kVei4O6oi5jPieBjGcTKZJ7Gij0HsWsCLY1Ph+sdCop8
DCPJfMcuL1BgviRDbQEbnY6ll53Puw82OlFKUenAk1VREUtoNv/blFsfit8A
WSO8qXtLLLxdVKrfAZbTiQbYIr1NPagTYiWHWeAi/8a3KQYK0PHuVVxtXDQh
Xa3x0oMlvrsx1IIkh/C6wANtu6gydfp33IEH+ojeAgRbJlc67KjsrD68KMbt
tGGTHyEvxzO1O4zE5MlIiMg/dFFQzaQmLzuYH2H5RX68dJU5WsQvDIfGgc4v
BJ3dqQfzssXOLCm5FghY4gLnTxQyWvghnq/a81uRMln+fQ46Z/tmOBY9dEiF
qpEzN08aJI/rR0K24uoDQLsQYUUsky28wKLTUrP/Aax7X9Q1UNHS57AZQ7jO
LhndSXkMimCDSdyQH4zEBVnl5mqqY4rSDJfpq0MWxFJBd211Iy9R3Hjofj9b
rZNcfHJCJgBSoPNbFhfqLyzuNyxjvOyuL84J6BcEtaS6ee36Xf7a/UFIYAuI
zSR5qY1CVCuwAWP0ilaAhmJS/jucivM084NgA7QxRWBXAR2S4NeKtyG4oEeW
TRrhmCTweWkHB6GgEmnb4UeA7Y5Hojki2SY/Mrh3EdvP6RrZx/XFkGyZ75ev
IBPmrl/AWA/hsbFBj83ooVzcGovVXBMC51FRueSaBP7iJcYUkBjCKyj5t7hm
6eaShpJDHXNOzCt4qtE31qaIsn3lNBzBWSAzgl/397Fx1D5bC040zOJNMuXU
daSpcXGeQvwjYq0y+nMp8kn7tIePRRpRAb3fZWxfaKAK0PmEuxeocWTRx5QS
eyrggFpIEuDmqr4ypmNGaYqkdbJlV+Xv6Hw0NqzVzjuTqOoQ3kBBOG8Bp27W
0ouG3rUb1pGP2qp415YQNYd4T1B8UPuvYjDxVUpeP93WBWHuq3jcVBPRqI4+
ocFOBJKAQOmMLwBBNPb0i0A1SjmvYfQXfU9ZPyxn/Ha5Iui0r+Ij82+qAgVk
KZR7/+9ymfln+uzeYtacn4rIulgq+jC7LLHwxPmlTTbny+jZHOx3O31dIXoL
D1Auae1qPmZywlPgs5UaR97W5qMaBr5uRTJq1CtvT2u0+g1Kfjs6+4+zwlG7
2cbrPLgeqvP1Dy+EYz/lnTqVX3S7HWWNjcF4sGQWWirxOIYZTAp+hZ9iTs7I
/UAbuzIkeY0C9pIHxX22OJ44i0R2naGhxwZtqF0Zv1VqKnql079EG/pQxRpZ
OkR7985GJ8nXHJ/ZLyWHKtJwgwAVF2Yjop4RoeWUrb72QZ9PkViJsM7pmgLF
uayuoXYeZ3V+THa0KKeYhYWeuTceYrP2tlyX4AakSDmcL4zHbgXO7bQfcvUA
LHvAXdWxR0ajQwzfNSbMzuSdykr/0tgSHi97nUuEv7XT4DZfC/5rGT+xmfNF
O3zCcFNd14Lt9e1fzVfCtEhG/cUJ5LeC4xwSxFcr6jg5bg3f7qQ0DeTPK9Bn
0kK05iT8vCYHBY3cpqBArRWZLFj8ZFrGQ9F4zbz5fMvV7vm27TFqVAyHTedC
XTqIq4a/fqmkqkFg4L8pGkqj+aO5F2olxzr5yicaPqxd1d+WqLwaS2hDAZJE
jp6gTJkoWOqJ4uwHanlMkeQNTGx4y4pqHnr7Z9lExH/IefI5MRLn7XJrYshU
boHn3ZiyU1/z6VnamD76FZVza2+noPrWizNZNOlomrtwLyYxeGj9NBIFoNO7
Do7yPokCPLDMdDOrO762XkB16C2vONfzwFISGKXc4SFSryyQDsTuomBNCQyX
qXIbap4p2YkgZZ4z5Lyx3HLrB5JxUsP62kxmGLnYkDlZZDYj8O3spDn/o4ey
xWqc3TPtv8jkPCKxcKs2ss0mnqVOGmhGAaB/JW2mNIMIqoW7QCcFx4XGwcx2
viktxESnhah5FtCLFR89MIL7rmLiN9qeaNZxLjzE4cqsaLLJ15adFBaC8ZPU
fv6IZnuow3+jxGUgYSQKTO5h8eiII+PtoWQ07vGVZRHk8y4OrGBF1fPhWw8c
ZEODG2r5sXuCmyyV2YjY4JlrWmDOVVZCjDQzPh+W8eQTLit7H+Hlz5S7DmPH
Po6E8zYkfNDkS8h8kabFVYM/EobUOG/uKCUkLDOR/siNOQ9FFYD+8PuIRQgK
9K4FOkn0aAwflQOte6ZiVciV6B3puR6Wp1FUKYs/5hbnDWRWrNbQp31suNBM
kDDOWgN+P/XlsJc4IknWtBAyEQu6+4Er1kuwPSE1UkKuK2H9lH4BfOv0e7Sh
dymdu6Ekg5yQVJy6wNVG97HYPnK1qYV0SesAcBiHczg57xbZm2AY3+EShG8z
czcAr6JqqKUUyJzurpCbYLqwDPccZtIbSUmOdhxs+PVhHu+hT4rwOxKQoNlA
0XZSvJtW6bM50LrMAZYxg5+ZiILC6nUrGR5lhI48zs3z3mGBa5wNOlBvwwcI
ADdzhTKuRsSpOlMTk26gkb6VAY8ssJPS1H1c1UyK08tx84nRZSz2MN7wT0ZP
mdMTmjDgnrm9ywZF7SVjLQt8SY3j9DnpqVwsBKysMfAA4iK9LTCCL5L+mYls
COeRbQB+GaLWSiuy+ibGwU3Dol/5WOOeUk6zXZ7ptD9rem6Ey5nDzki5dWMR
FPdtFAdwCWhE5hKBg8CXLHWyaGlmCra93CcuZ7Pzh5mJxbEm5eGkyOz+X+Zo
EVb1WicYcVe8FBeX60A7h4GzzjkrhrFCbTcEj1U8pylThRqql3WdnN05RR9B
0Ftcpq6bFRr4P0QsvNYqoTPY7zODy8EgCm/rkzhJLZngFPBAVAPQDeoWoKAN
MplT+DPFLNdjhB4BCk91dMuiHeJ7WUZgaMPri+MmAVpWv9XLxvLpaujLam65
cv7DQuEHIPurYgCfdxDnWALuFwBVUFYMfe9OqdQa2k0/mCz6j9ZztTnd8BA4
PFprsJmkMq0Zt+dOtzK/i6H4t2Idkz+nvBVHWjMrk3VEzs8NWg6cbVRmFGkU
hsBwWWzFlguIU2CTKaMxGXCY9AVIuJ1adBeQWz/budUucjblK+M9tOzGwm1q
unyhUqpC7mlhcwGIpVtBDup4ppJsjV2X3xIjQwi5MV+ETHtG8Diia4N6phZj
EwnQmpsJW09666NrHrDFLV5d23imSzdLZlemBjZ2FhMx5SSRDQitdTwkV7iY
s2rF/F66gAmVBsknV5K8F0j5lYTnVt/nntkwh8F1lK6sp0Yia4l2hx8UOvlU
z3LAsQin59qa8SPjdesXqYZ8cTNYY8isMKzCEM0vE59/bGpMN1+ka9wbmKFV
b3gLKe0OEe5JP8UrCYYv5CpbNpKxSV3BUysiarF2DgN7akhdwjGMaj/tiQlx
S97+JWn4Ht8cH1vouUsGfbax55rdmAOtikCQZhMlkM+yRl+jwOni71YYFyb0
R990dO5FXCZ0Vzq5Yh3BwicAZ/hfdQwG6AlPzS7gldn71dZR2ya+znHE5KaV
iwvknlffWS1DGVTpQhmvdkTGcRVFSlx9cy7E4nfaw39y1npsVH5CPwYkHYr1
HfZIcQ1MhACbvE84DSXKjjKBc6sprPdJqF+DWe3hNkve2T+LI7VLC54YDDjN
i/Fwc7hPtj9rdhtxlszpEbM/240jOrYY6AQadymH7zvkvnhIqnHzF/HkX0uc
MPaPQi6oGla9IOD90/k7SIUe3XTQbuzQx9HEwtVUSRMZ4Fq/w8mr+VWXsXsH
sHgwgkHf47fioL59kAGEdZEF5/nxllJ5zAhVsdCmazhEJT04pJH5wklop/K8
axF8yJDo3tUaRsXkRYGZY1YQoL238X/28c4VobZyURFCL/5KdkSwBO6kzEQb
XRWfHHnh10yeM0xsY9CUdZBJvT5Rl1zOhQSW6mAWiHE6nn7I6kNxao2VW2yu
WA3wiGXd7T0156a5dI+aGMjO1QAzIpJaAVEvWM2c+uIvogjaXHftsX3xXG8G
PQ8D4NZh3iaD00b+C0rVPbyEon2eHYeHqjnv0gZcDGtUc2uyO2MHUw13GZbx
nNBmwwHiGUhA/M8T0ZUfK8JEP3JPibpHY4RB7bTlnEruDoB+aIRTBePz3Eb+
tfxJJX6eJJr2g2ZNaQRzDS6q6y0mMaNkD/7cix3YZiIaIdEb/nsSwUCBDmxR
N0wD93AOcknmMj4nK4pBZ6ZQqcJtLby10fer7k6tcXSw5DcPKZbJp0NRYPvY
ZNmMSJuSvvH+JM3m8rUDPjqWuYcjgCFVlHFveI7zil0RhmMQviXruBKp0h8V
GJVvxwme1p0lbFRJ63oYsm9pegpKeZqTVV3voV+tj2ll7SP1WW6OHmEb5ChC
kgv89iIozmGUezdJviNBMpzuxt1umgupt+JQnJZYBEdxoO7A0/XZvNJZjNoH
dThUBVeDd01UmvAh7Zc0ek8iVrf7PgFRoxs3GV+Tl+QnQhAKDWV3C+jG41wo
lCgSeoObg5lrLFUjq6Ux0QF377n2l6XbjEYMx1Rq0RL6rzGKJ8GR+hXWW0UX
quBcTK7ZTNxjbGm2lpy5RNtAVYbm9TmJyg7M5tIac5l+8Uw8BPER7KjRmNYw
/A9WXHidglAIXOPyhuvqiKDSVqYlu4628L/p6jh1YqSuDYMKJAufgoGJyjIB
LXYUcBkc9JzNsRxmV6fFQ5Eaic7giiDkw8Ei1wzfx/hHabo3LlRhMtgGX2GK
rKvpZa8+AvUmWIVo3PN1jrGpwPl9FG/AzlfKW32S/a55olSf/r6gNDGLPsRS
wCS65K+P0Q0sTsuhoZ/zIM+Qs8ZaU/7QuetFC13C/47V0aC6oqx8EuyVX7p4
lbxmocQhnfp7BowQWJQ8uDIIUl1eDcPeQQQjHaCFoGk0FqP5756F218RC+u5
YGb8EEtDQeGtlf9L0HdttGVsCl9C95drK423ru1j6cSla/QLBorV9GwBxF9J
DzKtods6+xt82NpxQSiSDdxBWKYpGopfVX+xcOIJ/4vy55O2YgOuenux28q1
5/nBfnD05I7eq03YetBboi8ORuvkqOe+rHgt5si7/HMWAMGl8/LW/sj/Zkvo
ji1kATAG/46j/pdhd8EmU6kWxVByZgCw2Dfqtb0242y7N5ukE4lDBVKoDfUY
ViNg6KqsysE7QuLOqZreelXhXl7yE4QG3eNL/t4dBE7tdvV13JSfkbkoBVO+
CyMEGi6+5PYitUnKzC820EIeJ5oCNDy6MnxTOCYQRKk//QIcpVH5PxW0AcSn
x4AkEEfw5r7yRT5TvAK6uCXCeiZi8+bQ6tU8REC/rtJ5clcm+ZSSaYRr6I3X
XS84eNA10ko+/FjJ9FC4dv2OCOlvcUy07hn4K/B0TTLkCz+AERUczC7PjTdo
3FmFSEJ5dEu/NWMb3LPzsH+UUPIC50viOrdYgZT6oC+rdzRobbk5TOru0iFq
ZBgloZtt9gQqZQeqCTV28xWfZ2ilmP9vhQQYrBKjzHTHBUt3TuDdFVAAmMqE
7oWfOMjjkyRRDtsPgqT5RShqauVx0KImjZwLiOV2dZ2KOTb7oGmXVHv71J7w
1I5TRoG7PBZgtWICZmCa1hQGcJpoWgW/2TnCRfIvC/suk2uvS3yKDVmFtDXG
NJo4RnkZ2D/J9KVNY3mRyLyzuzoBBa3oe2a+7vnZiFNxRx2F7v4BoJE9VipN
T51Yy+xC0dXYKgvFos+QgUVZ0+jlQ2HD7Lgc3cjLJCEG+7o+Won+EIz6XjTH
xuIRplLo5omCqMfDnaNgKloc6ccw3qFJXCytJ/d8dJDFATPRG2Nbyro8uhjy
/nT7hoAVF7M0WQqbyW3H3rfbx/b71UvS3iF75uVzgh2SF2lkefMFHrxwaAlC
fM5uUawphvLRMJzBYlvzPKrPh38T39cnf+av+iNO2aMdM1d3/DYIU4sFp3sj
uCAMSqbb0NMR4U7v83YDdFrFShNqPNiJ4RutvEgaNaxYg2teg9aTM0MMSe8V
k1JckoSwgvwV18tYmPT8Kaw6lxNPAOoyZbGAspO5QKBatXyG4sjW3rk96XCI
k6pODaadO9TCbcYGUBtTOT7615/ZianNg5zNh1pEf6Bdt1ljzYpjF7xZMQ8Q
TAI7vKJO4Sgj7lX+gQFf/Zp9foHGUVpXl9scQm1TTkVsinKatuNndSjgDjqF
oln3eL5GBv1vY3ALY1A4aZ4Wc5/+5Z1gK6WpMeZiWo9YkEpy0IrtxeNHeKIU
VNNBd4SwfjtK3JPiirLhXBR8FAaeoAACW15qXar1bN1K64e7rnpFTeFuwXtw
uS76oNMSuh7D6KSCpmtyIy/CdVN1kJk3cLu4XAAZGHcK+6PHsB2NR6OdNW0V
eBk/rL5R8uuNDnllJo4keMVOC4rwT9Z8dwWe0pqvMggzDJmOOidDvAliNnti
nLDWS/NjF8s4QBHgUWWHZ2H9sM09ZcYuDrJvb6UpajSW7M0r89XrVWp7Pv1g
2RHIv+BSvKqa+M8c2ULDdXoHcYl99OVH3LxB0qnbb/a03w8u5tHa1INCGPjw
2LfKPgVWjjtUZ5ZuP/Y7IGx2K7SbcXTAo/kqyTmccztpC4aoROHzxf5Afu5G
IzgE7GFfbivOsYenJ0ls8u2IQ0ihOZhZCMW4sHZ/PFI2ika6fp0IwKebahlg
N4bFGqaeZ7ysNmDPAst+Kt63peW5hhel9Qiz5xsc2/Isn4FvMUY8P3I0G4Zl
B8WLcdx0RCyXdMzqpbETyzGxIm7G/S4fuQE3k3wQNEy7OlTPuMJd0HXxm0Jw
uoX8hc87dNjb4ooAubRWj2O+p6V+DfOn5U6kFcLPID6/X85iaFjITA0ntHzN
T67it/QXDAsDW6JZBWBruF+aILW01qJ7d70E/LiHYGghnSgAMx96qkOCl+aT
ehbSMOekUgvl6eHjl+1P6CWtfUOZuT9hjagJni2z/C0sdi5NIVIMdtbaAalG
uctTvUd7tinzUvKcqql10+uzUC+qWDQWplM+N2ovtOtP+Qt5EQuEIO1mAiQA
Xs04LuHK8jH9TAFfAV6Knbq6rR5yk2HF5oTe62l6zb8GimzRjZazWBNuXA3r
ughwYdcmxOUzDZI3IWGdfqvsd6ANw0w8VfiaxYGvonGfhrcFU/wVKrqkkC7v
35UIQrA98JWqceHF+HJ++CcCoLp3bp+uIUJDp+CpkLLXJTZv7OFy3QXlUsmQ
wx4bUGma2qkVOYNfPsCfZZ68Yfx/HcBTdTmE9NaoNoCEBDkT5DnFhnhtksgU
D+1i/TNdms/sb4Lul4GJzxIZqkT0GzpKlxG97f5k4eb5/qkOskYvy/Z+llft
ToSfeNvAUuM3YyY0LobbPlJUoS+Szj+om/NkoXbri5P7wqqZ4e9wgJfrYmNf
T2/A9UbPbABafx5o4fs+w8Ku+9iurv42zHczVTs2zw5BGdUV1fYgmBToHCZo
uUPzADjsJu3dLetU3T84cO08fBUDtbtdcni1pbuB58LK+xBrAR3Mbuwy+peO
oafzaJEdKWb3A4fU/2soIlszHNPIONtQcuHse9HDe5ZDgVCLbgmW0CfBSgsJ
Y+rKEVgePaJ4dD9OOvhInz/t4f1SzrSvp7Y3SQO2K5v8Fo6pwnjAS3wZyaca
d5erb7qoeCA8uLxuw/VOkm45GnDblrl+YGrS9wRGJJu0tBh/xScKUZjiNJt3
3ai8yJKLw6sapRLyXAJxb9NH84sD0nJag+T6cp0CvNhzchsEzFuJYJD7ELVm
QgxGBlFa3i56bVQVdZSTuwqHvmWlWywTIyw5q99IllsMgVH6o7UNYrTSGG1r
j4D9+ervyGHuXHayqbXpbEZjqSR0Jn7tmNI74fAoovNb2ZQNWnHj//huBKxE
5Ih6N5wc2Txj8SW8ykZaIlOXOzMDueFXLj+lkQSjJAnHwSRvUrb/gL6EhJyv
FIXGXrkM/OSQW9n3hoVXeZ1qorRWx8C/0d+BabnDkwGHu/TFs9DbiyEUdh76
0Tu9wTgS41u+GXnbCmP8zwOWemamARWljS+KrYzn5MiKT3Ltx32LScnAYVF8
IigB/BOH3sC7vjx0KSu0SRbQW5rU6kG4JdCSTkIghmM9czzKPAk7WtxWnvpk
1SZHujqWuJHDIBOSwDdO1uRvYTRgeu/ZA6ZGC2kfGqLgfP3XiUsFD1j1Abj/
XZ7yzORc2b3YGixWiN7pBgKXmQT82GFyBIOJ1Oq8fnZxaxtODczAFX/SzSfb
XckOJ7XRge9Ffth4WKeBIP0nnACPcntdyw/vU6S8PHGSxapBqbdVQgr62XV1
q9DHv5YlSJhyit7Gqz43Nwkl8jXtixO/WAnJpp9O9rvFhvaoSDktNxnmfrKk
qJPO1Mfu5qcbaqXkSIeVwBSm8VCzGVYkoTQLVqNTW/gSFJ8Ng+F5ZbLDNZNG
be7JzJIOr4EZGG+HzZaxN9sqHW2Q3XmMH5TdiJ/xUi/EwfGl4HetLtNvKcWF
IzJq+SXoII4LxJFeROC066A/49sEVD3spshfsAjTF9CyrKTQBwtF3JpHZJu8
RIpHl7ccsFLmBpU/xeSxbejcfhzqMIDAKNiMOV8U5seYe4uFD6rGEokH9P4O
fZ/RJ8icqYa5bW0MY0KbzsPySs+sKUbSDqdJAAtIaxQ8k8p3SWpO0nNt/GXa
H7k7nURed6P0jSkHxwC2oM7dyWBD5582iyea7N68iud81QUJ3eaSqUDbBcHn
rFxGZONLacjQt/+EWHIbtvFFKb8Fk/BgDrG3vtdIb1pOnL7Y/3gtTTbJShhi
JEr3NqXOeMoUxmXiNdKrOYjnmj2PPByQYVWJVuprTZpYFGDxz4XBAxKSheaZ
Hq6VVHXpGa7CpYrOkZWSbU19zSKJeu127hLoXttiOj8XnttxtcsRf45GarNo
laT7SHqKUxtgZ53Z5rLEkD+MulGlrV3HQPQzG2kjk4sC28kHp6XFP9fquuiR
Fke2c8EKvuuyK004oH5PfTlgrLNU2PPIwALFiyPk5hpVVKlUAF4bb6xmM6tT
54ys97p8BFan5ZkkvbTeTOYP4v7oCwqYsYTEknFLkJPS7artfNr8ECV4Oe0I
y+26IyBa8LLjE6wFtmD0Q45cNBS6eBZ6X0IOwZEAz/xbXkRIGcyGuvJJVe10
bTFkfy49LBcsgj1f1CspWd64O//YcvI72ttGSWf18bpPgINE5i/8sUtKxiAh
ZLd7cs4wFshcTw3PR+owgD0TahYGzuK1hKi25FqGSPjXdN02MEBZ/hNK9QoF
kRuDYJlpsnRm0F0m+wl9IsX1Cx5XI/QLI8iqUqCrnqlyDx5DiSCfSrNlD4De
YfVa1DeCIuU8K1N/9zc9x/M2mmiA7uzafZa1I0PF90xpaagO0FDQNYfpaCTQ
k/JaeKH8v9dGS3sPjaWK8mPyBVgHbLsw4WhAqgPOB80gzB/6mf9c4+mct1fb
DZIOKc51C8SdJyaCNyT3YjZPk1P+p9uF9tEMurQFZYgdzwvU8aXYUCLmsPXn
b8rfaOnbbvWoGNTjD80UNqoT1FiHVUBYUBZvj7222YoI0AOwvwiT+RCEEF3M
R6sY22M70tIcyZsiomE53MRcHQdA7SWMSY0Yc2kwgDl3EZlfkjOXYyC6KWaX
pLk5MwowHzi4bkxjQvB2/o0F6QQWmbSel5ZEIJ3oGDWuF+IerT6ETIieLBE6
+qPu6i1O7tp0f5cWP0kulf+zeLbnb0i9H2qH9Asu1ww1Fnap8mJ4q+j0wu/1
t+XNRkun9mKfS6Y/cI6P2jN8X1c55G9lhvrTxs3iHgROMWuO7emcEZO7WMXO
V6ylNgyNiIXxgMUxxe7phD+Zv9IlP4Ki0zcgqX3r7UyXeINkLaMysRwA+A2V
RjEjR0YuP/yBksYwqBBzQ0arlIyT738Nvn/wBNg/SbxxccSn72IfIGYaowEF
fJ9UwOLYBrokZCm4Vhn4PeDg71lQTJd20au/tVI2Hy/E1CqqHydTDsAbiO9U
pwie9NlC2rGmjAw5Xni5475zUvmp+7Vu6aGCiFWTHvoiHORKArWkKhVTXgPU
Ml2LtNu3zdlyKxnz7ig2IbA8bVQQQKP/Qn26nYXUaFdC56OcmADdTZywLs6J
PnWkoyiLWgvZYeiTF14zWoShJP83tJasHLnN/nWDp02H45mQPgum6SDaHexN
okQj3YjXzNzCFvCbd+WjK4axE1qEZBYRXZ5+Dz8p76jE0jWlmu2M0jmmRoh0
OAeo4OLMIkGy2RLOou1nc0qYLE0Ipe8pFep8DCqgp4GGJU9h3vjgjdDZRjwU
y6OHJmCDJPPpv5GBMzj4QJ/XrfGs45FIdYFbELS2wros4D02VJBvIUkCGmn3
hPQlR8QkE63OjFR0BWZhkbgcoW8IX9dqbtA7Zx1N199r2GrSVvWpKDYbCNfW
njviYOt4EMJ7wvQKvDI4YzB81fAQ0vESbENCzxSQwJjBN77DIVFpxAz2unTR
cJoGSFJiWr+gazAfSZ8JUa5nZ/C1qy8UY2OB2h4X9T1MwUWy2h4hkAarcc6z
TMfWlPwfSVlu338v07U/zTVD/3th9umJ3Lpb3RUW+k5bH3O+U+g5D4V+iZeM
OFB86uBqw8sSul57sdf6yYcvhR5/V6joUO4WBZiRqzaLCqDkvSVzaIucB4a8
H4C+PKqQJjTZ8+fscjIAo/41AWGl7qnsL+8uUeY3qGCpy8etOuSReib+pOv1
HAclFclcz/Gcr+36E8E+T9FOQB2tKzhhC0cUUCWVSVrU9eQnVerLuHOycXlc
FmjgHvJ6osrWLfxjRdENCg5cu8E0KvcbBiHjacpMuwTU8VEv4kzfPmuFNyQ4
1Pfm3AhsXVC14uJXraHl+g1l7hnNkOm1Z4Irf80pAdd/09g3g2TXeGDu1oPz
mR1EQiGDZgEWKv/z5aui1re4d0kLvseCHEvjOmh2gJxlbMKck01kqw1ov4KW
nc53UuiKWPGWyiG9whOdBdik6X1StSDXqNIOtEWhMKVZ6WbHsFSS5h/Z0tfE
maQDrVOP12NruW4vUaC19V4KTNTECqYS9wvPSb8EjqrhzOBL7uHMuAsSH4XA
zhgVnopn6h7RwkcaAtmVHIH1qts2YSWCsBuh8RjpKTUlbwNJ+QVeojqEXb5P
qWEqXW65YicfKiHyudUUiqDh8oA/pNFtd52iQJZPaiOjYhvZEIMqOnanKMgg
/j/XjnHcf8Bw6CUJSy9rp4p+w8/bD+zdye2u7cbFIpoztAbRtW5/WUUDUT47
bj4OJB6DwT/PYGFvvtG/vhodOpweKBL3tQftEpQaZbMykBcGpES7de1VZbsg
/C/SQWYZdLkfyOwwX06e7Kjlv6vOJc07bELykfMtTBRy+n8xKyhu0NCTX0CZ
0qAts8ZfCU/90RCfmFHEh+lutrpYv+uHUzzlbCFGt94MOppzIVsChdLrvH/q
k1PvTYFiwIdWNMuFmeNatgFodCr4/S4KgA6MhSMpe/uAh9oFI9IFha5baVXy
6yNMcsPJVcMm2l/SAJB3prw1pBvIL21pkpWs0UyvQyapvk9wVETzrVVSuGem
l0NhBi2M5D7LvU9mvNG8OjG5ZeSOq00U8tnp0CdDrUAd2j5py2LZfEsO5NkZ
W2s1RLl1aqZC1hMSJ5f6OG2ylOEjuccCvuTU6GImbx2iAhZXqEwJGI4aLkeH
tkmkGOPVJAwPRxLxgE20tEQyGER+ajo+X/YSVvQmt1p4G6H9uSYph/vk/zE5
Hq7X1wIfUfKb5Wqd4ZOGTasvzMu+ih02zWgBpqJO/i0C0jRqB+ca0I9JJEEO
e5f2YbTEMk9oF/eV3K0MdM20busGAr/3CNDdLFdrgx+vrkjtpD+qNR77znwb
UVYLFPnN10u06sGnVxImkfTycZO58nYl+Os/QP43xT48UxfcuD9ws8WNCZSx
B7F28ZGfJeIbRsjwx4dxJEsUgf8gklXP/rb7cafjl3+AdX8U1BcYXQymQ3LL
21A434TfZVE5wYzvWn5D9l3BzAo7XQIkUct1tfpAq1Sr4wEgEnVj6LQpXeK3
Q5EPN2ynpmTvGhFeO3opzB2ocsJ1j2sLing0iQ6KD3Uga2GfUiXUr8shvauB
hKYkfjPKAzWTgI/k+D9ARyR9+SknCqmwTaaFcDLcou2caDOehRV3T9nrMw0w
FqynghFioXuUGURZnZmqSgzDydzLjJ3BiQ5SHTvU2GwWEC5h+4qxqLvqotaj
S/SrMI85X9eRmIpxU3zxu0fREdKeKEdfXYfSFJ63gk9k36/vxTO3Mpu5z3cL
DYqi/xPfOvEyOUiI3aLdye2Ge2dlP4AlQpieUwSZQev8A/kja259NarpCh3t
xNLEvs7whNqdgjmBuzIKHm33vuDuFtSN3geko4cbO9GrNsqj2jTaQVIngrjZ
fXQjza6PrmuSIQpAGpCReVF0VntCuuJPL8pBuu5hFfNevuOuMLWwiP2Bjbr5
tJp/agV8xvC+U2f0wryMNQwxGbPkXyD/rg4PWTvQ4EVXze4oNU1uNPBvT26l
Lv8LzKT3uyUt72RYphJ+2y5u/hd4BIpsGfeUAjFGMM51eiIsCmu+J4U0hhSq
rrZoSI25J+JZ3VgFXNjSYY1DnyXBctBIPbtjJIaiCT1ZWQOAdqEVEEPaTs9T
lmPGQb2p2DnrkinXhEsk+2sJTNPqx+yH/UQZQc+Wfafmo0WkeFoDQ1GwnKmA
YD4vTrIRyFG8pz1eUZCDYGGrLIfMPUX7iBRQGto2C5Dkxgxw9zM0ZnFqG/gw
+buzOE8qgOLZbfSkXEb2NfoleFAUL8RPugDYKPXDKjTG7Cmxm4ZNfdlQCZYx
wilUy2yjVK9uhx70ng+JD2dQiQvLcXP3BCVefQpqGqg06TwQmqsC5ena/jsJ
uqDUsTCC2GZB/DeynrAy/DRJYci8ppV3YVlDb9AFu8rZ16RI15Ew2ino1ruh
mu+1P1NX1efDea3AX/kPr8Hpa5Fw1foAY9BBtTHIjhVSUt8H6eMXmXhDbXDY
ZWYbFGFQ/eNXnByjdgDJ0yzJMP1VLlmcrIAnB9e2FdB6RlL/brXYsFT3Q/Pc
/GzxrxDXkuE8eF3OQjkElfpjjyE08XfFvzsf7nR0HfWJzvlAnvO6/3g6RJO7
IKVzVQhJ3rkxbyGTu3E1kuiOKfZBCzfViCgTxd+mY1fMo1AJeTKZBkvrXjg+
8Z8dxfLIfkSdpmFMAChrOcxi9c2WsGMVs1NGP4cxP7Wt+SAo51hoTmO+itE3
OpR/n6hePyPRtRidRSGTqBJ2E1VRTr1ZM/vIHFbypExGfnerO8yFEgZuSGSZ
h1LcRiVYgYi2Z/A14G5x1a/AF1Q+yLhRDL+IMqINMlxmLZHq3Mgi8d0PrpIr
zbsFwbHGPk0WBHXpEaZEVbotPfewwwZ6e1+7YjFdd+GRIh7op2mj2TgTmvJA
TF/6ZMIWCg+TIHul26iBtUr98MRbLAKLZR3pIpnDAtcCdm6yhZCOHdWf0P37
ulJa0mRswjItokITSEf/fZRxzejck4RGHBbl+Pi63o+O5tuH79Qa/luAqeAN
4FYuGeh0UdgERjvJgyBvBddOjUQ9eYv3EBJQNb/J5PBEkNx4SKC2fFVospxL
f6CGidoTWmdU5jEYDOtFK6XTxqs764A3tA2l4EG+B0bJFxSLFWWcUPLT253N
KwLCparr2iWkdEAuht9utIJpooeMq8Jn6CFLDSNeqI4rKe/gAkyoMZTVYyu2
VioSEoT9sr7THJsVhb6JNKRtUEsqf7Dg0C4lJW3iDvhX3dY9EgBZDJ+eRkjh
u24OEbrgDzdIb9Eq+vwyP2devkatbLmSflEHuqMk0+CqS013iWb9pFjxb/Fg
igVV0IrNFQ7zsaxMV5YdeYS4RaYhdwMxsG8drCfkrRBZXaYIEdTf4/THa+dG
PdCsmcUT3P6kexr+BGsNPpmEo7pQIPaBY7XZcjwp613jGF2puQjhk1IOiFFt
lIXaF1E+cPQHH4d9XoIrdWxWSl1qLwu3WRrBWoEKxeEctIz1V0uUa6r8TlgJ
zRo1XVE3g/8jedXrRUkSedK/GqsIbZbpCoU/ks8G945jaMUziW/EnlInxHUo
fC76c0933Y381IX1HOQiAX4aaOvlmVOpR24th6EZHhPGZoIZJqQc2Dp+sxcs
oovviD4GA03cO8TjnqN9qTrEDopXA+V6I2RXl2z9Gy0nxhj/HYV/FCK+u14f
o1QJEHuth8r26/C2hDTHmMY64iS3705T5XC0qIPAGZRwqxg7ANgw9KREftqH
Z8r240mjIts1Jp975ChDaTOZfpxhJAZjonL1g0zZQOr605CY3cYw2NPgQm5H
FQcD0litglPHQ4kFd5tw1YT7aHnBt65DutDNH11ZNcS3OAXgGDvau+Zf/mMk
SBjyzJMihm7ygMZ0tuGVAhuRtMpXkK0XtmpXh8h8FLtxpCAP6w6aOd5oKTG9
/TPgkFM+iw6UydZCE/wpvMtpn2TqwBs230nW+oEFWFvZy5aJdyOPToBzHm0y
3O/hLHgrqjmZg7UIsFQDSgEIr0jPGVkNQl9BZSFRp6ldfYT5H0OstniUrlrm
bXriXRqc8B0rRzfVRdBW/WTamTrcH0rKOxpCt9yyj0UBISbn2o8JxP+1r+xN
791K1VRFHgvsiEQ2ay4aILrPIhsiNC3ZRe+1DlumpFXRuI9noWJ/odORf8rH
bJab/YvwAaGPwLgnUEGfHLnqHmytBZVVQGDyL50u4m+drCDbfDGrJ+5/gAn2
5pNyY1TEvL+o1mToQDZPF36wTq+ER7kF1ilSieUQ1kreefwvuqCh1vEkWr5n
xQWNHfvq4V3KhoTUV2jqCXIcLTDJM/KdjuQZRyYs5d7ohpKRXBr7a7/A2+5I
x7BJhDh0PuFHxyQZzCUnnrNiuVkHGwN3uf44qNqwPAeRgTcEsv3hU/BW+HMB
La2KviEScqR7tPx0DuBJxnf3TMjIixpDOWhOEV9/kM2fgDq0JWSXHb8CwdXc
S1Vs+/zZzpbizoOxI0lvQD2DKnW/BM4PxdBcyz6i5fmpMgiFTmaWzwG/c3YP
ODJe8tOJcE90CMt4LlUhuI1lt9SnzTmd9AjYjg/esStyIf0dz53C7CL6DEBl
lu4EVbBfaTkQQ19M7Ur+BvUTvPX7GmBUsIhaCtapkbEGZfbAJzjYqwz3GirG
SWDQNS/Odo0xr/vJgN5eAfc1vznN6LlCuZGpUA/XZYJuQcZRkZPG2pzZ8VdK
iDB8SKSt6kF1VSBRjTx+iu/b5rw44oSIsHrbsKEuE0QzrQRwkXXS9wuqvkP6
6R+ymEWsFRiISzXoq8gk3q1SEasRxVJlCjlKWGiPNW0EOs/g11Zca7SjoRsb
qMDRmG/t1SC2mJXRHxpEowPxjB2Lqf+TeZWzPxJYCqE5xGJUtxFMY0DzsTcq
+7wqJUsJowe9JMfaRlN5V+1m69WnbDAEsVl/xZjbAvg9FCT/ZUhtUb98QfPo
kPrHIeTy8bbU9IfVSNgB44p33gQxcZqzcqMpm5d19QM7aex8fiEO873UVuhl
CTSDZIEFHmQIcXIMtfgPPGqN6pzKLM0dmu9Z/Xh9tN3qMXICGBTkM9ySAOJ2
XW4Kh7nWn5sG0ch2y6duR4gobUniGbp9U6z3lvnbSznPp31aUn462mrGlTkq
lCTjI3ZT2iIktx+Nh1QI9F4kjV5qxsGLog0r/qxKyrjIFriYXu7ZyzCiBUQC
de2eCpVZ9axxddXhf9QnEC0xZIPUg8qw2AHB1+10FgvGGbteep62ptdIO7x9
luFAFaEyB4gLs66DpwH78VpthCKv6GhsODhzADAyvYFtWQqdUWqjTGGghmh1
KvXzfTsmi4/RPwsi+L3GNHxOFnZlcvfdPcwLRqfeY0QFF+UHxdP5EpoECeP0
9LTDpeDMUQolc6vo0Wirby4SXA0AQVIts1lL93FhxtSz48G3VKVmc4SBTgxB
edKzu1/patr6IM9CvhqOmf5esp+XF6ryC6AgafK/4Eu6AZBkD7HSuYgz0DAl
PdNKFuEdEJBYGz8IlzPb/JyYAiWeiqMgSx4APqYdUaIp1JvMT4b4m5RNZDjQ
M08NYBdFfi9LDetVjBOrLUmTg8JTtTFsb4Pe+nG3UMS6hTyToSeWCECXo1+q
KrxC1kPFx9Sfud27NW3cCoCkMR2RPJ7oWX7kXk36xR01yRT1nQ6GIaYTlBtw
IOiVaXehiscPKXNfcPiPBHIEWEOeSp5tWlMoxdkp3+Hx1gvKf2qvVHJiXaO3
xxpS5406CIinijE86VyZk6dAYnEcGXoxaS42OllvuZ17SnLeIU2KZ3YV/jJn
efvrfmS8FSzNXyO24AkW16rRIAbyqPrZbAULHgD5XQbh1Lu6wwlxaH0eIqEG
4FjQdqOZ+3BEmccp6ICmx66NLxObNCWfSoIPU7YCJN4f+yP/stPNTiqNTfCe
3aQ10svQaz8J6elHLrUWDAlY6cdZdzKaOexVYgDqsEeGdYlKY88vh1hY7sn3
ssW7E1vhY/JABCW4EYUkJTJz/l3tAOZgy+pP51ItFvZw5y6LgTUIK4A/AjJQ
/q6Bk9dzpT959EYSo8UcfqQafvwfFTnrk0SQYtBaaq4/NZStZKgGDiIVDIdm
6awNV+EpctqeW+S/cBujHi9J6XVB0rdJ9EKU+CPEjKLgzGcQYiGutWq0UzbN
eJYJCXpC7FS6MjDNBLNBodCVLVfFv9s0cAkwh8oSuXLFCPesa1P06/+yqYk/
qaORe6Ab5WOUADUXX2gFWHAqpGLwUPSx1P3cFTBzBmUg2SHRMhcTRx6vVxVU
8OHER3dZLGNcZmcnVZGiLsqrpzZ8iRMYcG47OXJRV/nONkFZ5Rdg5hGCQXPO
YKnKcuSMk2CVsavwY6xpZTSGQsBtKeqABuHAoxx+Q+FVab++S8qQ88Aea5LP
eUUDBtvgfzxFsKyTpn0of+/l/JYiWss2PKdRuFdhlHq7gIP4SJ6kIQ7PeJpt
PwpKq4hEACRwj6WQV2eaBIEfZ63qCHaiTqWo/ZyqoBEX92uAott/nDJ7jY/p
SGCj0c0l73CEe8MAgAEaHgeTW1DlNETBNseoqH5+wLj3xtSDLkngTaxFkUzp
GCrnQ1cKtn2NcfSybHAyXm0jvNqcjJtDz6FqI5AJmZjgo5XvGiLtLzLfiGvm
RLMgkcDIVAboJNv83Y90qfRgnDG/FZDVuLlg9NwYXY8p2BasJvy8PS2M5Lct
QPP9wofIUBUgoYMcsneSZCZCzlztZvtUNYLj/KJ+A7XxYHxcUiIyTvyyopsH
XpdPEVxvE9HozM3tHWj5QHDudSX4wP2Q1S9TTDAG7hxmJJzWThHrQMBd8Be1
IxGhd/pjpXFNZ/M1HS0sm/Y66h4UQqko4XVlEovpPD7H7m6xmi6p1HLHQrlQ
Gi6UAxL0JkJq8Me6v3jEodZoGfs1NzfTVtDz+EcvjtZiFzru/48e/Xt8kdlU
2s/ccomyV/Zj+ogw97eUDRDgPxlskLlL1CO9KQPunhuM00I+QPS8+Z2mbapg
CPhwCWvD6XAvVQHxW0JVfpR1BI3hbGXHnDDBGqz+jJvbygVXlefpc8PGhu5R
9q8M9nPE5inbcEjadRQELlk7HoDytUX1+BC+cYpdJ2KTB0gCIvvmHD13wTSF
OzXZPZ31GOjB+vJiw10+1Q65Bt6QqyJKOnM3rIxIAw7ldMhuDYHdfFKkv2rT
sWXYxv52MMOhfVF/DdWipl5SklTMGUYNIp391aI4wBZ3us9QA4YiaEzFfjIu
7szE4vD6glsGnNX3+Q3y78LiLMVHJvSTr7FifSSsixaQQ8SoibDWZvg2sKl9
Oe94tKWcHxm1X2jbSOIPm+VjqWblUjTaXd8/yE7hzldZtFkgDGGLRRUqksmt
r+sYc7vt6QAYYIcNtejHBquWujTOh1yJ/nntHOQ7somtFjrdiVPHZMYnqWJM
TJ0DxUwG76oqkYZWCwrIPQrBLgrldSffS0ZTWXsDISqJ96DzbkwCrdKBwCou
quJfk0n1Gh6G4Y7ja3DweVWOc4tkaW49YkRT19KLJOj/ig1lMJJdX3c8qpPg
lwpXtnRTG4bPPtoszO2f7mFTkOUlxmGsq27lMoM9z0hSYNzGneZ1Ev+syvCc
kCipHNxMXyRqPwJdAglVsjYnKy9kgmPaQ429U4svOP4BDGpeIwPBIYNzYwRk
DnN9n2+t1z82zLs0cf0PXthayYZemkprBUoAeSctN0MQdG6GUjux1bG7V+iU
YZP2QkxF2MAnkqh5l652BT3AmhvR+bUpa+B4ykqOQgvVj4QvbxooeI0uFvXn
ULJEQA0r/3rVTxvlM5cs8SCZwFFzlTmYHeKKY2z4M/2TPVj4FjWK8KZGp80p
MBl/yNQhReZg7hYhtzisxrNGGv7ircsvwQFe50N7ZBZMYw60+X4HMkf4Un+z
MUM2xFytNSM0MPqrQl7GeJsjgi12g6c6qb8JEr5OzKxcGr27XaZNYoUADTtO
E0MptdBTjodMjH2Ckqda10fZnON/vLBmm5tD0OzogMgCdd5GMc4KyMlsWGy8
Tzt6osWPnI+OFYADHox/kVcUCKLuyL5mhNNVDU6Fu646VTnOBbdgTIwmOI6P
yKxfzPPGH7PbrXaCVBj6Cx5EYRl7rPOQQHxRXlDmaEstx4U4vnNZg+FK+v7G
0wy4FZeWBza8tvXCYBJCnHytro1fjth7N5aZ9gWi2/aI7rrWQLaQZMXAgEZH
Cp3gCAeipuHifSgZ2iPUAxI/nVhFksrQ/QDV5TEEcRAQ/uHAsB/SM8bkSswC
1cRmsqnUs5aiA2283nS83lTVAAcmT5+Ei5bVEYtKzkErtTYT0GOfiw+mZIal
Ho4YF1PzZAXVQba7Oq9dkS/MKzPBw3bHR61g/j51BXoGd58i+zalXgNjl0vp
i5xh7xwrHhUIa0s9/QvKZh/PATRb6ZYiq3bi22Z+nhtcuntWZmvj22a23fKF
t9I+epfKEDESDAGv/tHx8IivbRM5vEQuU3uzxbZBz0AD+eLFclwH5GCaVsa0
H3GnJbw/G2BGwNXlsSpLrmafIR6QJ+4J+R+JzvfzwQ0XdzENesYx/Bw47+i+
Qz49R8Wj7rGVO2zU+HM2o99zTGP5pzjulS79Wqy96EwQ0pOtIBSy3NsfEv28
aPwW6jxfFr/L2G0d7e6js1IXiE5Gnd7dwoR/Tq30f7EtG599ocDAKIbADJMZ
wvkbHy7nEKedUEnsXcQ0c1ZYSs9mr84LtP3brOZK7jldYNgJ90DgUuld75i0
8G6IzVpRrL3ld8o4I/xwKzlTNvekEHL0FaaVPsLTcwm2HE4bXn1JolrvoA/N
QtflI7onbeTbVrPzLoWTFX/IDxRBJco+NGLU3eeYws7pLWCZvGLv3X165Fp8
e6CkszCKYyxr0IHXYTOEmWO13l3QGCcds2JG1ixWTPX+pc+vGX8zOlFUoUi9
/RyQ1HHvDQomBdvQMoh6Fi6KNOc6zoDC4WbfC6I+wVatzdjtUE2IynAIBRGv
tmtSN+DW6JbiJTsDu4ADOTZftOjnXfMdhMjesGF+npSFueJMAfJj75HJf5Dc
pd0xHrJOqgFpG0fOiCg3y0jXP7jALv2gRRChBZk8G5062cvJl0UVRD7KjAMX
iZ6GpgiXiiEVxM6VI4gV6jbXHZq0BrUCjXlzmJCi4IklXgqCQFN3TjxiIzae
gpEsScX4nV3yF3fgEM1c+U5RHm4uwyberJxQLpksW28vVzx5Qbzg6Noo0VIO
dnW0UdZ4HuGC0UP+cimBM/lq+Qf8hzXef4yzbKuAwmBcwbZidosM3ECIGbwZ
1UNRiqTi+SDshg9mmTGKzHfG91+o0vmdyVMIrAkeiRpdzUcq/93P574HakKg
/7eoqlHFTtRcP6mNZeCiD16NupB9b2R3MxMopNbNbbqQ+mB8mOFExK8+drg2
XtiI0Tf21NInaeSUSnxtpvO+gxDuKO3oNVyQPedHCvOXDVXJoqDIJ7Bgt9mK
mUXpu9EPW7+wr4KlWxqERxVNPAFChgz60BDWKYFebtWCtyUmakabsNcxcenD
WbiPyI0bW+tvLT0b7jRrfBjfcSmYgEY/M0GvOFcqoDBtO8MZ7HhOdPIiDkn0
YJEM/pk6lwkxPkexQPqOoooTpxXXc6x6bBxIvqa03vGUwozQK1p/vc7q+69W
jk3IN5bzVuUw/OxDnOzMcFXbEIaXTnmPyPDl3RnIqixCmjV65exnVFOSHhHS
F+BImBiL7pkqQJUZPuq4BHSddyXSXzXifB16BaGiyMCRs+iChJZ8fwanoTs3
igmm8Jv4+AgKcdC13Bg+rcyUSFNhBLE63MtakMDThtRCxVvE8R+44qlv672c
esUidM1YYoGmwaZ+vIHldnAW3v/bJZELfe1IE54dj/rnxZcIdfEyqVkfSlX0
G3iWnuD50yXHq0dMwD1wlWr86gICmU8QCfiqrh6vgWYhcJIK6bGkWJrIGm5+
mjTzGJgoBfHGd33Jh5P/ULGKYFukGLFT4VSvi9G9tUZK2MmG8k59n8BM8FAk
W0iKpamESdxUbgoWz0f3eRDzjQVObO16adruo5KyxF22RSzjwOcu+NoV591h
VwB1+ZQUU/U+PC4nko26N0zI21FIUxPjMNG6ZXLZjGSosQdbAS25KylHyAoc
eWwU2x97kDVjyUbYnGU+3DliG7P5dVK+hTjAu6AvK56lhriKNehTizhV39n1
iGUu1BPbMqwKbg0qbwGMlJB8QeP+AzXl7Mk6jbuztveP9Y+jZ1VLCPLlvDP5
KyMEXTwXM7Rs1OrNf1s6E7bP4rLZqzUrkZnO0e5Fkj3/w4J1wBc6J0m+dP+d
LJgKH4A0i+hSJKSp1iw7UbqOsueEOmM4nm68cXNGwdjS68e/LHpeygXNXO1v
ECQzII3C+XNcTBd9Plk1U3YfQH3r3tRjUbA6tkzJyFmSmNB6jxK7HJQ+z0ab
9D0kQABjXOAcmVpsJ/zkS1yAG7oHSizayxJBpYK5QWd/VebGFpVn4AsE/737
x52muKSIBv7Fiujftmw4egtoy1r7ahK94rq33a0iZ3/0QX2izNrLCi6uOAgq
4Zb7WN1OmiQfj7rH7xzFlF7edZJk5M9Cz/ILhH5ThBERu/vzk6Fp9iwqZdOK
Ks26Qox24TFSU1FLaLA5BQueKUE7EAfmDnet93Gg9BnrLmhTOsCRvWkXNetC
A85R8Uw9+SoPWyY/7SMEaW4pxpqQ6zj02fjAMhI4m2+VcKW/kgO34mURi11n
gd+/iN1hMUkiCJIBCieb0pSCQGjNTV4nrnZsvYNa3S5Ql1Ek8ZYuLeTEsph4
X/ZT2GWgENwKwb2mKbg3iWgxuQLExa21uGC21vqoOKYRqNKWuXFadUhN6scJ
YDQ5cRMIuXR+HulLisogtjbwTh5YgNi4pSI56vk9W71gFJo78TQ1zF78JzR5
fAN2l4e4IGHOaz25zQI+GU5NFn4P07ecpZAqK6syNzOghw6ZmU7gKjnT4exT
49saWWgmnvYd4tgCSyT0+zYatCZ0C4NsRl7RS2WNZKhuvh1qxYjuVXUKhLzg
srg6pmuv5nqBcBjG/RQKplpLGp0Cd0la4Rz5b50P5FMDCalFFA/ceHTby5SK
you+b5qzzjro4Yo/4ic6lXiu21bJa7i8ymw1e7+0KkztFF5E+5fx4fjbQWmd
I1fylIvjh0ZBybkkgnJNs8BTTzsJldLUauG+AAIW1GcxWxJ0LuFG+TlhrbG8
MTD7tgo9KTHrVK5QNb2X80TAE+LMoR1dZd4QvavJOAAPV96XgJU67bnWSIdr
rLOg8sbhlzlRQ0TqjOjabRgh/Bixd/smbwwIcg/dhrwlGfSs0AqhU8qA/smN
4om5W+ORCo2LBCol5dap4aMv+NP37ygOmg++mw9BrI2Jvk5Ersh5LD2a1tk8
RvNWfq1qXtkF17H+3vjCjY5KB7ZEgY96UZjDGC7onZJiUrGLrl839EfJPCEx
aGbVyzp+hxiRILqlNqY82j4RbrY+hid2Q97Cj6KNczmXX1AdPQjC/jnXC4Gw
w+HfDGIyevZVqFYk6MX8otRXw29n7FHGVSQfuYOw29z6ilkfnIEOob0FsuDr
UlvJ2U0XCmgk2p7l3xjHGeLUHJ4AnUTlIQ0L8c+MYlVS9CGp8Cy824AoJHp/
qXdFbTu0QI82gSD7XcAT2vxwJ0CaeHbx6wt27VazVL9S9jov2d4EsWRmQmfI
SLMQ//GKCI4/M+XP0i5pB8oX6kddNL6Ikgma8ci0KeGkz4kUXV9GnQDYHpkc
v9b88+TaSxirZ5eY/yGcniW75VmiQwAi4rR+6OOZX/lLzL05/mOQ744tFqAe
UYJryJAaRgKTRawxJTRd31TWAWCAlS2CO2bAZKFOJIqZrFM7p2fEbnLY4YDl
UHef0Pbr0/RIAHDeQ+weDUoKtC9T0AZQPDqQsfYTpSu/GFyiWAnFOIZDIXJe
sxEBSY4i/lzsdlrnW+VUSObdoelgIR/dYNHpGm9RhYb2cxPT9Uqiu7g3vCPR
zmSXB3iHm01wN9el0/lKI4CPnwHcib3mXiz0LsIT6R7ME3l847Tc1bN2GSrW
4wF5HREgajBQUZHKCXR5uUk5ivMkZfHMvJzCWIyHqLIm/JPmy5CJ7NHeB39C
sVjFAGNmZhQuvyAZ9//AVbM6dMvigQIfceowFc2wYE8xLbNui5iWUCsO9lnh
YtxQj2qLMpXvrYt9EiC7kIuQxGbpLWqGZUgYM7bhzINrQyPvHGdPrc7bHy6M
3noNCRY1dZI+IhmBr1edvoWiqf5oaXsGewJsed5v5B2/vqEGENipmvzDupVi
7oKGRlpUIeI1RaTvUZx0IPu92wGfkOYkvE2kRQeP7s1gnyLctKcK5C+uJnrP
0mO6bWNi+MvSEzt7qsiT8X1HJBISolpk935Eqxx+MB+Tk+82LMYKRQO9Xmjp
PQt3NQlDkS+AwVxyJRdBN8R1J+xH/mzlY4kbGW7Y3R/gBK1z1xFI3qitfJ1J
NV7PzSouXs/AqKdDtnYRR8caUW2TppvQa0kT5kYtQptCCbkAtxayOw7aZOgO
RiuV6Kkv0dEXuYdtlbUBwbkfY1F49Aj81jAys5EpgIg5XPokYoi5ZPKS3tws
HNY2rskLF5dhicWShwShkyMuTYECAHniTz6gEFyg0fZlS1ESchTLdlAAGNNu
YiGOuSnz6I/xS+vPbvgDZ/WxPi0pUFzOHXOWdzzBJggZLjcxWyTI9ePGS2YW
0PteuvwGgNg3TvpkKwPrOAOPJ5l3oyPph0EZekbrxlWCG/+fYCB5i5dI6KAR
hFXvG2mruwWPYvldRq4k6i13GJamfP67TK5zTz3IBKRzu4PEJ94TLglgsIM/
xwWijoCwQoDQBSRDwauUcY9FxgbGi0XG+diOmIsWTR8Mi7QCCrukH3q0Grb0
1RwkvFp3J5QTn7wMKqrC9gRg6CEh14ILTNw4WPrd+d7e7BvqVsxDClflrvn6
DWmWM3mSz+90XH1QPGdaYcLcIdtUCxFiOuPEHfWdIB02xysf/rK60Tv2WDxj
CPm55ha1exb3W9q1rrQM2NCmgOry0c9dkI79p4H55dghiPX+k0XFwIMWJUZP
Ia4+dJ1kzFc40OUsTxilqRkcqys7AH/I0tr3A9bBUJdAWi6Hay2mWMtceSni
B+VUeg5CfovHyz+YrD4SNplvvJ5BMqFF5T7LHoQKrscUIH3xd7RcqfqPzuoY
RGyhPDWQzyAWq+/stPpyACTs1gpPjraUtKeLKHtktdx+lbL/DLpuiVUtQ/Mm
6cc3PoJLQHsu2YNfnB4gpr5B0AhO+UXSxfyPieSQ9E+FoXzX/F7HD1Ql8arL
8XEcbOuFWg5pTx8AwI79SSWo86SdIQJg8erdU/k3Wo7nyIn3y1YPyfSZGjRp
LJg3KwbR3AtVYmdiqPR/thoKDbHzNOEu7oMJWmDIpUrSZQKF0+H8XMqGpfkq
bQJVJEkCqQF/S5Efa44aRkRNf2ojKNKTbxboFETVNXyCycoq1bJ6jM/H8+MO
j/nJDtUgKg6JI9viaeR8NXeCcRDbimt+T7Wi5zf/4js+Hnty3frl5dfWhRH5
n79j3zebRlAG9Sgj3bBf5VwHizvoZlmqNcIMvUQSVYD1tuKt4S4VV6dw+19F
q48WzR/CvpqOrdV9n3T0vXJjKW1pColWj2AN/qHJVh4XgZLRntu8h76yXfKt
OX0/mKMckOJx+VDkOfZd9SKeOGl/A21wBHexmc8lfJw73EpXMY87mztv/Sb+
LFPmyWBJI5FY2r9iNTjeQbpRjzT9ZrfPCmRTrqtajcsUkB7DjPke9GK6PQ7Y
prm6Mwc8YmpwhdX1WYPi4qRFzrDzFIG778sCnnJ03J1hraC5gcm9UaSSmSS1
gqjr4F6FcvQai5QqpXlzRoK7896XKbk2G7ekFJR8oREYub0vovPKvtOcY4EP
ooPQDPIcc31miOtjV9gRogG6w+KfsViWjR3IOiDlFZa1LQjchymauWxhtkbs
44ml7rT1UFPG6SimY3zk+UDbE6/Spu95dtoRn0bYalOEvqyuSKYTgJlonroe
UJlx/vbKWTM+/jxS/ITsbr7ZLYCbyfGnGpYZ40Tdg31Twnt+/zx5pXJjTj05
zKTlWOqtLMBFiz0yoUYs9Em2eJj+6Kaub+8f2RA+Pr5CwKdcrO6HUuCmD7JU
LS8goU+GkoLZCTroHtRV0cgnn3USW0u6PuJgkL2tDjmYljM4Jfe76lJmEXLh
NmJJjIbZAWHQO2bejLm+mUsj05cMvc2AL47blbXsNn7qM5VOq8HdaR1W1w7V
5PBQfeKWNzYs7s7fdH99cQIDMmyeh3p8jOZUVEaqJ4t1IbbAXS+35Od+CAd6
jX18V+OQUyNnb/rPinwps8wbler/OMRllVYuiwRltQ+2dJ78GRK/GWvz3v+y
/KheZH0h7+Xkr4Wvox9obqPw4afbCkrr6MHdACDX2RbSJ+gksKvEjwqcpiHO
l4U41Zcfu/EV2Vtt1QifesPxNgXaddFjnVj9zxYiDJIGaphb16oGvmAOrtuo
9Wu7iH6KAnkMLHyFANgDFLlfLF924kQvyi54lTgUtImRKe6ZMD640ZdMmxyT
UAP5ZEK66w2ZOmuhLa8Uo9C5lfyNv8sZf4g4CpdThmg518VByJSNyX+r1GvW
2jhulJvxNewq94LqDQvLPzXBGj9Eh3bvftrM0Ln9XjY+ocRMeh/nT5m2NTlZ
LO+zjZB+PpiMo7vjofRIymi0Pp2V0Ympn8CiNQvmJmSG/pXN3t2c/O8yvkEs
s3gp/x/b4CJ/bnxMgw5RwDJaozlQNsi3KKpgsu20FylnDE0753PDnzh2N5kx
bGtYQ9xfE+RJOJ3DjG7bZudVkHjU7Ire+Obsh49J0Ko1NkaK5sSdDarW+9yG
5bMz8e0rV/ydNsRYFLAUjul6MqrlbByE5DhWpf7BZHWDkDdUAY2i7w3FkOD8
89p28OH/ElvptjkQwMTk3fAVAC11gl0vtLD97t8Bf/TZEe/eF5oiheoBohw6
4xQ/vYPkNSuz1SBgXkIeeZrjlngORtgZe3EhstatOkjb1uGx54ipAhGnSiVp
adS3S1LMgC4fQW8pKAwGeYdKQrRMQE8lUtjKu0TO/COeLhvgo4oS7GM5A5EG
JYDZMNW+3LKpDZWRJVtCw+/ctZkCOu+IVgB4RF0XIze9qrS1z0GbmWqHsMbJ
tlUEmIoxU+BpkUaRbtVc2YfaTqpslQBnqKRxVV3uQVASSE+o8bulwPmh0qat
zvxBJWAO6mE5122Aggcc5mL9O7UHl1FM6fgj3j7Z9VULF0lR/E2x5+RIp2gH
RS06OnP2nVxKFVS9osQ4sOVL+oNRynhNNzrtnupQv6vlzoWeW/wApnh4vEFP
jhVUgDawfoR9qWyv/85LTf7f5XhLxKkAdVdYKvNpjdVBqPZ+Bv2oFJxenNZ6
8sME9DfUVaQ+xOBYdMTNPd5PVSASWn8P+daCwXZ2N7VJXrUTmGNZv6e6FMmD
Rt3TV9upOuIdrGjIjSkbpuZamq6Zi9aHH6SMxTPmJhAIiYIUUrApqWmPCnYY
4tZ3GAdB4H8OayeMy1+Js/Us0CaGNDlipzpJ2WxLGypP94YKxfIyIlATPiab
IH62rKp55EYPvIUXO+5IgdpFqeT7UfwHxm5sThdUL1SfAs2faqaxs669argt
1SEaXwAi8FJwBd1wFlmbE1sezDc44oACZbqjEQe8GZZ79QZcycAQkoTnKUy1
JvG2Cjje/rIBqfwv4WfOZozR9lUGFoFVzfOhk5rEqwuoeWKmAy4kNTjXTGSH
Fu2BmZjobWXG2G6oNsY7aiJWnSCSdXFa7w8A7j0XYIQ+9TywzPkOEnouju5z
0jhsv5PS39C6cp2bBoDCW+TgRzh4MPISKcgn+/RwqmFaEXvTROz8ZNhNXJH0
wyPF//sltQmG58JatFUUudit1MH8JBG/+suToOwKl1feKHIbu/OvTnl//+1H
dhQRXvyxIr6V7FLMCSUBKfhIFCCM3YDW8yUS2KLI725GPEGuxMqMAEj5vq2L
qM3WX+gCNo1xWoPPXx4qchSo+xkVBq7i3BCBD+Lz9mmSAhAKpw51kQmbDfVD
tz82driJuJwY4GUe2mImtyNJ3P2DCKUBqXHjVsAT26rlisJ1WGHYR4pmOpPI
vubPHOUPwookCQ1uf0Ho433/Zp16XivlV53XJdC17YpFLDGrIJcQg6l0xJZ+
t8qQAAEF1fypxz1ACarKS+14upaU0XsZZvvUOzNGq8iIO7zW5cSZQIbr2vtP
LU5EMTisfTpBe1VovE18f5VFtpOppGCxu3Q5vC6CPuFZP0nRzo+wBRb/nTKz
x7aEpKZKiAJBZThce7A2GUfQo7XYKgvA6q3HSidFpwxtBv4bQ7fVFki6vbll
Pg+S/d1sK7vxFBSJYJkvSuKbflx5CYy8y7yhOQhfp9ck8Cy4z1Mc8yM5RxVU
YJI8iPrUbgtecLZVRb11S3eiVmrOlCzuCh/r3l/aiipl1blWxSXdIfA4FkW9
Mqh6NvbsXVniSJ5GFu5sHgyt9RMhjG6I1L+ch0XyifDZB8H/N9fKYpXbX+ZI
TZbpu8/r4PDud3sCiYtT93lvpQi50Ik6wCcp3E89KBy6zk35s18EgJ7rZxOf
tKrT48AFtJiHZalU4n2wadACzyWPPB+7pl0wn9gfWAtMtjLfV8kHT1UiTRgu
JfYTjAxC5j7T4e5dQoZQnp3UywUjpITvmTsuSzMGed6k54NIZaYMzQ4sUAl7
e8zuC5wceU7OrhENnMf+/n2JTbKs3Fod40j+zM7HlRoTXnuj91hx1ZMGq7ep
dlNcapt2DzaYHs2USk7FGJHUm0pxZoWngAWDE9cQ7neqV3tVnfDrZCeZe0Pe
PWiYavLVH1ZdCLbGy3D50UGjm2eWG7zGMv0bXiviZlkYcJRunQsf1F1VQYmt
CYd7xeKDS3NN+1fjIoCWFcYztsA6x+1QMjIVHEBuNP4ssoHB3L4jQ4YyJeCg
rheN9VoGjrpNTl5U7+0sA7E3nW5pQtKT6xZT6iJ0fluktZJCtJ4q9a87riBh
OByb7pngtKiBbhcAxbZeNLqXsUACxmYjNKGynGkXdRYwlfM6kjynmCmUb5jt
gcZTqx+dDl6lrWnszkUATnO/diIXHOFWE5suxfn/Mpqyg8/qHXuwO2HLPPgB
ZzrKdaaMI2WzbOjKEBJfDqhs61MzKmUsfuAYbSs3pzhwe4nZ7bgk35XVfA4N
Dpm4fRIVSbv648yxDhl6Ni9hsmNCPblYl6a6jgnIcufUOJJfrRo4SBv6rfSe
gOX1+EoCrL7qHpd+WUJhlh/VL1PEccL8YfP70h8lyXnpkF7Nv0IQVZMk0O/v
uacqj85rnX7j/PqA3x9rLLa/kTii8sZhFYIdglUERrfIAJX5KRqZEZiBtsDC
w9N2uIETVxAAe0e1UtTBI0DuAWDffyl/uf+sECohrT2/m377BDGJK3sL1eYV
jJzqu6LQMTOjTIqM6mNvkLxNuh/Az+32UYDSrt9PNkSL8kTJSa4hmLcGFWtn
pj6YHjuYaIJpeKkaE2j9laMge9OSaWWOm0++N++SuccHD2/RoQdESnkErCxR
MslWHcph99SRCzStb4b+9Qb8QbzDc+gvQ65PcMMY+jreJ7RkT/OqX1gUevZ9
INSl1XoyFQXgai/g6pNvgJwB/SMHaWUGjc36yTxtVbQ7LshlJThHLi+6yAWg
dor8aeJk2g1NzMHWbVFZXVPo9HJ4ByWeSy/DzW31KHtfV3LPrZTVmSbM3j7i
8x00RH29lf/VCwr+dhUFnPG0gNOpEHQkE2Er2EeEpaRFpnVTallI5VewCjvy
OgHbteGInooEiHXKY0McJHbH2XwgwqewDdSlVfc2PKuormtgvx8tNDAlZhAh
9fHZUFmpjwtWrYb4iCyP7aHaHlQSLBBQi8diLkXthwBbrYmm1g8feGpEtOIH
d0pIRYI0LlIaSbPhAyhhVEMD2viYQtHOJg/XnKZFrLZ6hbkXTjy/9yyrF0nx
NGzMswONkQtANyTpGB6HqXVCTq2c6pfmrIhtcEl+4iZEhDnCqGlbA7zR+qa0
7qGLu15DZS43mLJTVfFsvWFkj7N7zKz9YXNvCQuAh0W7DmXNUTmao3a3NF5V
1HSIthOG73IU0yo7KWzYZXYzWalpF5mV0xM+ZyyAGe4GLBrXKVpGeSVnZ8r5
YJuyGfgOVOllTx/P5K2CPhM2oG0d5eE3FWivhBAaRhwNZR6uHrVipPST63O5
nm5TN8r2m+WdIlaQBMeyAbU6AfikJxFUje52E6qW+8M8L5YxqNCfUA3EfzgP
2xEXjMhyEkRdQ8/YvNvJ+8wVuMsq6UEmyuaeDwNBHW0dc2nHaTno7QXCZKmG
cP6c6RoInAvraXtQBn7RVMeyrTjHILG4ylFnnZkrPSMMttN4B5knWWS5WU6m
9LnZJFqtOLAmqTLYCX9fPaPM9eXyiCC+1EA1cWCfaY3JJsusxzAhjxxdEqxx
2jCCznJDr2C/UApFwgq4kF+OWEQqlqySOisvBjXGrtQFV9hnCtxt2IsAhwAT
JQbOASZ9eAaQeKzdD9KzZI/ikRVOrb88b24XMfb4xkRJTYz6axkBVXTwT/kk
fcM3wtU6O3DF9MTrNafiSwagT4Z24dVuqxOh1tcXLyQawxj+nEy/L3bAxubx
gFN3rCbtkQ/NMIhsxdYwuEYNWgkU3sqNLPE8hm4b43+UATVV6w2hN0o6cZWK
BVfytX2hgpJ4uLGlrAc06lTshjnJEOiA8fUobkBRIL4Sn4fJ4YTkipPqeEcK
UDrWWrJGyBGinGWYGu8KRhyu6W0LTKHhJY6JEPLs15oClGfTWHKW1zjICUvl
y0cxxdLzEwuGPCjTrLAZTKF/XN4Mxmjkw5CE9DM65WEwioAsFDvVml1LIMli
FlbbE4WwFqKmceAC1Or+YaKL8gq2N8lAKotOe12t1Ku6NXDl05OBhvMPgrDD
vAun1rT8XsbUvpo633fx2vErX7l5qbs2IKoMj5DErPKri/B/GSPoASLndcEY
BRqSdAd0Lw+Q02Xj/wQcqUI3F0/8Kg0jhY3Gn4xvXSBZTmGB0Ur1KM0cpABU
9CLnAUXNQYJjE5LixPMxIUcqxflBw7wXvrTEdKapagh4xOiSOlb7rPLaUvdI
l5v9f/BSh8MXOGiyA8swibPA2LyDB34N781tkEOEF++7uW4o7QH7Z4ysQkTQ
qO38cH3lQvpXl4aIn3gzWkiCz1v3aeZc6r9csaK0ycSJuiXlgtP0yna6O+Ns
0OJIBAzh8SochfeIA6RoKkAZibdli4jzjrUSb1XQe7JfI/fa5qNJyUSgBN9U
0YwVVHTNLt8rliAzvCHYeqcMoA3TMs12Pe3xQG3/DFqFMesFhnu9mmNubBU2
h5r8k9WBz9ypjlq50+FHGWWO5vKUI4/39wUj2uQgni9amCA1JmHJ5oWlOXyw
VsJL8Vmvrg3GCf/338sPekGJ0rNKZm0GqIoGtg/0LM1hnA5dJyrajA8gtQ9H
xQEH5ISNv/YW14CJLMDJooa9nHlA/8kqDmBtG3mrNZT5Y6QvpucxNXjSFFeT
IqsuqV3I6lq9slyEk+JFdMPlgEnm9RixQKHSfWT5c9OtSSJLmiBBbwBLWFZm
EHlXPMFcqbbEMVtaw0at4iojVmhBsfaSvIeGWEErpoN2dngaSBf/gqqnLP7+
+DaI2yw1A/8SSI+ucXUlIz0I6gB3FcHfRC9V4o0+SeXuYRMsLg+jce6W2lnx
xP/qNt3cLuAKj0P7fOovVxlDFYWrd6rHCnXEy9Telb761w77P4KRAFGdCo7x
1MlVOlZtIcRbZRSe41VTIDL/bQWCivm6LFScV1zc68+rbVVYhlAZe1SdOdrg
Ixm2DPhAB4FRYXd4LIPowiyIWzvP/+gBMiSy9KmlgtvVLs55t021wTlOns/V
5qditoN5PKK4+YFytWVSAHeQp2wqqpTnSLLdl7oVhIhywbLS6i9mkPyon6kd
qf3KFgmqehAFvDEwdxCmDq2+CiDpubr6VtDtH3vsrD7BciRR1uLa5gZVAfwj
wlqdDYaJG+tNS7gABCH9CIZoJ58caRFnnDLaUtPH0Fw62qZVXqBDMBhOfrBY
L3fg4E1p9o+4WBOZpcpid/FM7rOD+ihCVJwDUtb2ObZCx0XQAAf72o5TVfGs
WohWidYz44HzAjKfFXPo8UnygSW8UlaHMjvwn2fxdA2jRWEYxfhSYQ4o3VxV
SzRNb8VykQD4ohanlmfONQXGzuNNvXBZzIni23ggI7GapWiXV2ROT4+2EONa
yrexxPxgI7O+f4690VHqBGr6sPdrNBn3Ky35owHngK70eCX1a/7JROlUxkCn
+dJh0kLxBTweDHy9m0Hj35+3dUk9uG6jqMGcFJqXWpU2P9MmnlBehSyu4xFv
ZKbx6u821Z8TP0h5xkeMsnhP1y5WmCLCBz019eiVTqLefXcI3bawdVGdZReu
Q5HxHpeEmHLcY4mQnSZB7t7Uuy5oiZN/OeKV3uPvH0Mt39I6ml0M9NZF6oCf
wp+ScQa0bVW4ZvIK7lr8AwdECA/IBlNzcNvb7hZVMGywjZ7rdq/kmxkM53og
wk4pwdz3c/UjIBDCvc9+cxvaNW84Hk/J0pdsvnymmF6kzxJAmnV16HPOHdJF
yM6aTm+UMO+BNuOtm/I4Cv5pZEH/F9/RNoeIs42ExthEPns20FCgIXPk5qDA
NYvCHQIlBoVxJGm6EurBvpn8VJgpHgs9o8tXms95gCep4nsqjcYfOuo2sCSs
Tnxrat8g7tRIad/l5OWcU/wTgJNmIrzqqK+CpXm693rKUkaekrCwyYgQDUUM
wnvqXT4/73rb1+Q0tgGpd01EMlM1FJlQ8JPQ6nOZzLb+DW7w3uhHeiwNgYb4
E5PyHkiuDEvFwme377Sw9qAuBZ5Q6g8L3xbWD07CyI5KqXZHRKA2Y4I+9JL9
cVQDk9vjikhcPZdOf5xVVXxaQQhhllxc4HSCRXZl3Gauj7h9Mx4ec+5gbeFF
XdX1HdtOI5C9FOkzelrT4evHW52kVbHu4oN9w5HfEN9VTYkomV4awKba5eb/
tvj5SumutXkb0o2ZJz/PeHaT4HtDrP+zEsRKNi1+Y1qnx+7caRmKdLPrdA8z
7fRNDbwmeyld9yKepoeh6h9NERyoQtAW9iarzUo94/kxmlNFprg2iHJsIViS
5Ts/ae6b0EGfOMxvpcFgtAtOzjIG/NogtCCHae3kepfIPfT+uHt9AUcnUqQA
p5WMR21ts06n2rTf0n5V2libOyTNHuATi/ZQhbGXRsIT8sZuGCLjd0Vg8zpY
PN7N3xKfW4GR3togjir75gmqHnxCCN0MmkkMDfeGBf+HCWmpRwIeOQ6sWmR9
tFSH8/np42R78E6B4An2/WbWQxsSF9YPj/nUDmK01c0cA4/6ClOJzXTb6rtB
y/Q1GnfbgFL9dNUMrEPDR0DZN9CnnJ4fxKNINm9Hgys3dw7d5dP6zLIimAz0
FoXYsuF7jwbpL/KgznC6RRcB8jMFLg/F33olFJf0VitFEnQ63akYR6D8xOke
54NsLq8fPhdS+4xXqqH/0olFJp6yKws0EN1Hh+++Nra7SEHYHjWeMD9BkaUC
0kSsXoNoBRbim2lYB2TROHh1HR69/Iy+kIuOcR5E2VmE2jOy1ubmTGQn0C3Z
neBYLSeqrw958jqIgRVultNEc+C6eWDQPavwqyLPgPmBxceWritQz/vsJXwS
qbqfx0eV4GpJlgVzymX7BfEh81y1iBKd+rsijHvafMmD+AMGgQjxtEH8eu8S
sQnEedcVboMQ4kfTNvKmsGgLD/eoT6Mr5cRTAcSbN2ObcMTEC1RtCVje2CzV
cs9YdwLnjCgxvO1CGywmKFXTwBpO30B96ipknoNoyi1yRjJAB3JQgKSk1S7s
Mu407tLKDGsHRQMY40Z0ePATX9Lk51zPCOMKFyNXFTPPVfEHKNKV/IbANyu0
4y1RSJYg45/onSxZ5R2FjzexDi6x/lqQSeL/SKOC1N7rc+x+KaYScpHrsaSc
IRSolDRpJjJwO918zTXd5axCdnhNN9hNkjX4JXq/DnLmcdkC4gTK0EthIJJC
LwvY+yap4i9ujb+Udznsu8GRWb6qXiGXakWcZiNVoLGiNuboBIfFOpXdPuB8
psgCqImFhhHsIGvKTqzqAvFndDWiWpQ+ipbdFlvflVhnj95X2Tq4p/ItZUw6
KnrViT/0jLI9uKIYi2IMmCbNG3qYD85z4SKN2tAPDpuBH3B9+VRCSCzm+8KV
zzVUcsll3zbzMUxf0W2dqIy7lGXXOQ4HkGm8V84xfpCvQ6RmmjXYnLK6xSr/
lXshMWtJML9OWxiPsLL0H/lJz4co89AIs3KV4UNJFWgLOryIi59KzG/7UgYx
Nhm4q9dsac/HL+fmqBdw8oNgqFK4bodkJY1D7+EPNtzyKXwS1Qdd1NeHXDnJ
i5tdBPBA6W6rSLbVGWtGaCFHjZ5Z4LByONpvztk9VH11sOMrovAcPsa+rc0S
b/vIAO9N43jYar2HElPWKR5xnW8jegaC+Tvo92+CxOv0fD1UpWsWctkwaihZ
wcGCbr6sDLYKwoPtVYlF/+Eb7EQkYT+8H95yiGDBNoRHitUOx4xVG3c8K4iJ
zt6Ou/gtvgWjAPprZHQzGwva+d0MngoHl26sIkUzQksbget3ElltzPKrGL/C
oRGoIbvP4oheORa+BsxF2pQy5L4gcJqjvFmSs2yOrcI8IVsbtI3WHgicbKQL
I9kqdiU1//SMpKqzZPd7ydf8gy9F30o1/9SrLJiwKDxOmAllHL5KFwgGIZLW
nI5FjLXnZoGsosvH67qTJLxVTyqFtMIkM+x3TLW5ChOpgwJzUAoaMZNr4+GK
9awtikhMn3huYjFR4gY2Nhm9CPmgYo+hx6zPu83WCOOC+1YNPU0Ppknm7LfE
s42YMFzP9KZbaX4rrzI2GROuEK6C6KiktbKuB94BsOLX3oLIXEZtfuWL1cl7
mDT/Et5ORlYWvkMDsOD2EFksX+uuHFeqRWslRIxew9OOBfSfirA+TM9lwtEk
8ukl6H7jMQIS2c5iMww0OgfbUi8BSO6VdvSVxQARB/4LBmcHWj7IGgwNzv8n
oRvni6PUHIi7shtQ9klHbiFd671yJ8542SwPuVJwwuZn2zHzGWDzAJ0rEJin
7kJm/RZZb/yNNu4YvE5o5neFP7Q/pA6/unRGbKNDVYN7K6b3bGmA9UDOCkVo
zEk3jOzRsrdSlsakARoFFRY5fc8OMeGqOUYK8TLXezYv1+b631lybF1o0em4
FRT9MiBxZKGjufTfmhB+KBFBYdZRC19BfItYlzxv7jcle6gBdKUSjLvFLFR3
ZQZX3omuDcgjztKhJIUFxuhoP66V9aD7Wttm+LL83Nxtp8QQo6HoZqqZAru1
+TpoRTpzcdtelFxX/ycuH/3UqkdmUF7Ikq9nc/cV1Fefl0RzY0pn0E4pukqh
v8aRx3OIC/GSYpVZ+z+c/qzym7JPNQ7PiPcrbyMUpUXeg1s39I6u4UdJUor/
grfmkHQtxZtbY3EcGQ86f1N46kbxENs+j5h25AFeVKZr0D7jxbCQqrTNMfuQ
BN8Zuabb9f+ffAsnKxXbAM8gbEpW2q+ThvqnC9qZ3wbziuHsbu4X3sevmRAP
hLHb64dKtYPGBdTTQXQ1GI/Vvo2RzVjZWIBFQmlHsDQmbbaH1mMdmOoAPtYm
nDoS0aWPFY7vmZXCNrtlfm4qX4u0+6Uza9wY24JAedjnWETVE0dwTANofOYh
ag2lEsXybCu/KlSKaPNECm/D+114E1UPFJRowoZjKmC6Fzt/L5M2SEn808n+
vU+C04rhCob7ru1oqs4Bv1auPcwlTC7c04EukU2BQMkm8UToSbC//oqZi79I
rBBN7HgqcMbkDOnMkbW5ZvjNCSgRiIllz7nyyCugdSyB0vKic/gJF3eWwEhb
D3HL8l5u0Zo8/qiBR/+7A72fRqGO7OuaunL3xEH/gy07IFfPHvilo1Hvnp9y
8GZp61C4pCSIN2nS91YzbJDPONIWVFKGPgpRaOf+q9k6XmBNfiMWc8hEmMyX
GaZhKuUoiyj4wkvdoNQUdk+4369SKUtV+ewG6U/MnVm+R6GFw86QS3fnO1VG
/Kf1SpZS6XC7/chXWm4hqwokEJtjDuaFU7/8swLkXWU/NP7v75qCIyFyBKc8
Gd8XQxflMTeng9gagD2VZdly9fuFJ/7V/48m1J+9881Bp15Nz6OhjIUiKUoy
2izatpYvJEGbMXimhzHzHFSzuTklZI2XtX3KgfI134qCIjcKs/9mYkOpLYAY
g1J2H8JV2EcF1LrlDlykx705eeS2HLn22KEluA4rdrne3f357LCVSguRn8qv
Y11LZzN0R4dxmCqP7tvbHtpQAPu6jEieTGYHf/CzNxOs1+GyteDkkvdSJbtP
HF0tluh8zd4drnNWUfkZsr5KEAHVOs2JL0u6HE3a7c0c9RWCUuffeqOMV8dA
SadcBRV74k8Qhgq8gJCrCCTkjtgodTZHFDBHf9+sv7wtGSzatIOxBtWkBl7H
d9x90tH/0bf+6pWnU1sWKjCeGRKpPPcyzaKMNCKb3636JCXizZtkbcPFYVJO
ePz4d3LelEplXLbsskFSSNwbMjqwQ44MKQGXYsVNUjFPjeanY4sLx7liT1yC
Qydmkqfs1kDweHSD9pPkGWc65i9k5Pgw9ty3St9kLKPqBuAs/3LmBIcS3huk
hl06zk/eUxV/wwf7GgTp9esUMPbzjwdASZdzmjQ0fcyI98IlT/tJaEeOOk81
86hyBCTElJsrU+1Eyu+mcMf2XuhhVcaobBNaMbuRH7V4gizaqOu7ERkZioUD
qewGa7g3qjeXFDfm9giUtdQ5Dh++hbOytZhV2ntKyqFbipfN9/Z1h3dkYgvi
QockdmYXKveGJWh6jmxf6FsZKoEVMmZhppXgs1rwJtf0w9yrQ0KG5NsNdAw5
nfQvduqmWpnCshszCQsq4pzXjGSOQPhw0pnm8X3Bdd6kfE9vDoPGOyzvXBdM
tGRY/HFM1nhb9QnG/ExA3otJQ+gzq0Hhs41Q8NY95/YuwjV23icHjfDdBw/D
4sNSBTpeS1gqbItORn+wV3jVj81RlGoFmaU6UqIA62xoQFyKfNHD/yfTSZ1z
db0yE/VFEICzfkGuD9+4CSjLJDCkuzNbb4McX8kBhelSycfr5q24QpQpHoJa
fSSEY5OTA34mBXSqHUDYNNcWBu18Xkrykrvb/tKUSj7eXgOZgWqg5lIMH4en
Ej7FhuioIsc6mBPIU5ZnaRUVZwKKVmebiUXpLLjnFE4AlsT1Tp6eichgA4YF
XVklFM1Fagt7GpGcoZvbiN9G7iGwQyGPAqQDUTCiBSo7/tsAS5yvolF1aQGI
MS2QCgSTKui3MBf1bzKtaV1ePiJnUmmAQl7ISSkf3yVhgD9XHyzDyKPMVu8J
+13yWr/jGPT+TN9NHr8ONGSOvfrzU6oVd4EAAqFtnxeTEyiOfxBs5/HnzXFK
1VlH4veHyW4bm1cm45YgbaziigyMduihBKzaHZdXj8v3jLzVDbkimxMVuxMq
OXC3+wQIWDKwzQ+pYXKzOCbnh7Il2RMVU8IU108jqwt+XGeXkvyFyVRAROxl
6U5blX3CSsiZ0JpniWh70HuRuiotXxpM6B7SNq39SlEEH9YVRSjWw9t+jVxm
UCEgudiJ0uWbL5ygkHZN7erk9MvvSfGs9l9JhoeaRQGYhxxXtDjlJ/8mYtt0
KT3E+5ZFqqyUsh54Hld79s6uvkH2V+W/t/5+3NjK3i3suOkdpnB0odJxjArq
c+DljiL5bGUe9Ld3L8nmYkCLuma7M5zPZLkYkAKQQgeEyu0+i4GP5KFbvbsS
8vWd0H/Ie0aDDFDM3G58jwYXlarhfxHA4JND8OWpEJThORR9LfSzbNUGWH6/
OPqpCvJ+TU6fnwvU2mXbwYMY0VNin2JNgRIyY3NscHHLqSkxUXAEQWh0VrLk
f7+v546vHUOLafMtW7LTUI/jcKaAPhlXu6gjGIoeSL57dxRycx1NBSQX/Ws9
aF1isOsjS5s2m464+RX8uRtsaK1oqA7bs4E0mkBd+F4s8ZUY//2Uwu2N6bK8
JQOslsDZvb3SdjhKNKSy1iLNmSZiR/65D2jd5KK7wYAmFJaH1kU96A76dNro
IFw2zHA+qdwoxRXNRmm916qhwf+O6VK24Peh+F4NKiWkRUZ6Zdl2X5DSLa1Q
wZGULelTm2KqkcSqYaP5e5jaj1AtNh9cedwBYSvERqDp0tiM9vuBQlAbkx4G
E0jI+TuMmNsCJXAdQDJaGab3yWE278qJEcVXfTaTgxM8PB0c92SiE08pHyYU
9d9fk05A6nzryeml087IjB9yAY8AUrL6qscPoLZ+EeECIzMG1jvBznfxQsoN
wpcJ1nHFDUri4+fUelO8WYyWIBMXubt09PpEEkAYZxWT5tbGxedeZ6uXwoPt
BCn4U8I22y40uAHs9Kl/k62+egdBa/6Xf5tCBD2mBGR32qPKmh5EbS+Mawbe
HkWzkDuooqYQGQKr/IAcUlugejXAcZJNrdtTFkJ9S7UcNiz7w3wiQwMhJx2u
jww53vIeUSt/OBb1v7nTrCdaLWkUW8oh966EPxgNdSwhQ6mmhTtea1G47EAL
/sO6kzQiuxqtJ4FI7oqqfVw8xnnXA1lV16ogthSy2FmDO7UhVoHaNidhIGkM
sHHvhxDYyS89+ZPaKOwqMdymkNk20P+T6MgRVkFjZEVx6KUJop/ecP11JxpO
Y+eWDYgCFckRew/iTgrQDBpSp4OAFYq5e79Zl63ciyPfK0AgY9ywt+9LYQeN
afSU6+AbfU7OM/EjzcX90Sb4AgOZDj47QaWcCgaPPOflFABOz8R64O5aFm/w
W79XBVC0h4XQF6+5BX6K3wfCrVUyFSiB9ndeUYjGrPE3CFRqcSaAE89KRqQP
jEQHqSEt4mYPtw0KF4Sir0PvT4HsKZUV+bbflmYIK2djYumE8PQa9QzKyVgE
fxVkwxLVfsBL+12JU4oqaDUa99chhbNZRjAUNhGdCOOCnQ5+eKC1k87dw/pv
73n+jNUVX7uyAPpZjLMZXmlwBtEMEwwcQGENMzPZ1mcMSFHip6sZHvpncsmG
58dGrChxQqwu32jYwMSS7dhhvL8fGRJeRZar4KxdKE35tcohxHsPTeiPWaG6
uJ1r0GRQuErsgOOrDtm5pNsVe9zCx10x0EL6MgaNa83e4ARBBNlS+qbH5fA5
yXW2OtWfNdCvKFbdtPZR8O5Ht31i8NEW5ygZVIuN4NfeLOs9hLXEN5oLcr7W
7TlXFLgqwfejlEJIW2G6PXeKLB4iAitqeFMdbctiafxCbfd76oLR26IoHUpH
wkURZTncjyqr1pf29tv5SKKtZ2hYgFthahKmsxZ7KRt/vkQEmlKHDG4tz1U+
IoSshawtXDa8rCMx3j+cXwsNYSHXhFB/IO5HDxeYBGbzqfp6SYF8CJsm0rDh
8FydgkHhk+BN5mSJ/vBrfqMjJERr5F8JhqBKzayFyV7xaoMYrgsMtdmu7rrX
s0LnDTNLkkGPU/ag/eMAQfW31Guvya/76csDBxq4fku7ACC7NhMFvAGM4urC
/Be1/HctyPnIeggcx8pMS3Gozbh8KAbCcAZhKYoOC+OW8/B9XnixVk1Rf4az
/pYG9W5tW+jayEKbNhqbWf3lV0K89E/GAaLFa3+hWpCpu5KXhwQPHWl/rwtM
S+090IpMqOMsfHur2sZHzkRyawLJbUpHDq89IWS/xq4ySjEzCFGoqqhSRNfH
xmZC06vhwMlopHLeJorwG3AW05aRS2xnJe3SjTvos1WFUwLZyM8KtOkWxWk1
SZxW3ZskDxtoQLc291AqKvRHVl/LOrPgPCWGNVXGkUVctubF8D7a6h/O/DbS
3yVtBtITIbbVloq7r9+5nEi0E5QEGjDkvLA+ES4mPINPzdH7V0n13rXCGyZH
wmZ66cP/FaLzmeG0jaiZwSnBmukhnl7c4L79Z6U5KLkB/2miTwCWJoTqoTKX
b9xuZrEjUC+IBHZgu7EeVk70wNroQa9YP9okDn876TKP0rWOJZem/I1Osr+C
KICzqfHiIo3NPw5owHzXwQz3q2aP4BpecYjhXaxZ73BcoepKUqvKrBDg/h1p
79yzwD+6rmO23D8PYm+JLCYYUr/4I94Wt61cNRCgsqFWQqiOUMd0bQ8b10o5
XfJad8KfjCOs3FVrsmT8q6VSIFSDqTSma6Y9AAINQjHiS+Q8wGY0d2rkirhs
HYPPE/58eQLiShMsVruOaan3nwDBX+Mtv1RQyLvRpU1AzOS4/e5iIOU3rj6x
BS3CNHmC71qmqPIEjtUIYtPe51UIl6ptyNDR3Cvkv9872IUdaNFxrdZVlyCs
CvoKXH1nmB3dFcgD/M4bXKkiWtHRlDElwNEOrVrWO+S1TqFS+Z8lYCviQYRv
HvdEc5nPCsOm1Pj+zeOgkcaNqdfks9ErTuA64Khgi7QR7VwTvSqhfzvUg+HP
Iu0o+w1mn5qNHYBFZ0Fk52U6sUeQLBs0LMbGQ82LjnxTbhPX3R5cYLpOJof2
rTI8YAOXVjphdzKbaXKrPlfnP+4+Bf/EqYSjQ1Nbcc0RaM2t/mWMD1Nyi4pY
Ju5o2g+pADGRKT+wJmUoeWa+dtrsjYsjPNiIKh6QUXGSf197LDOsQ1CQLf9U
MD+vD1EWv7xdvEy0+q4X+iTnI71cVn62mo3R8XJWXfgEVkqCYOxCjmm+jzmD
15Fvb6WSpzhpMmNYal8B77xfgU/vbQhF76AcPBro+lwd0+moRHMJCUbSsEGO
DL7jSaisnD/IHNZ5FL8aA8VtD+uUEvLlcW/muokzjItKDPf6Z+Py+KYrImkP
xNqG+9IDy5C4V4tTxJllX5ztseTUAJs4qyAjiAY/lshuTB1IqyXsD9fdsIBF
1xvyeuezuPf+NzUrKCVJKdoMS+UKLQNkK8TTyvCRzfk5t9WReBCTgAiS6SKJ
j0vVbdfc5V9w3VOEHdu0XzeywKwMWeabAhJErFCWltgyGNujWcILNeUuFWcT
vfCPERwe5YpSBEoDs277+1CYjGlicozNTdbM3uLi3gFGMtlOQhoXA5g/+Enj
/xVw+rgtO/1mCr4h1A/Jp1zmY1E0W5pB4yOQuaChblXWzriUUM5XQwq479iM
uOYGsgxcGUoiyDGSk2u2meYnyjgAF1ppmzaDwZUl+hWq14CrrAFaQN7mUfP9
S52gGfsYvrp2UHTicwdCoddwwI3VeTzKLMVRjeMYox8vutRYT35ZbOI+ptNj
I/x5qdVu/04j108Swvq4OhIvo1/MTkua837k2boXs531XKTZ41Z51+hHY74V
yu+MbTM87+QNqPb7O2U7bszuvnXxjWNM8wqQwQA+uWjYANOQc3oLTsEYIoYb
rKrC9Sch2CjGTW5DqtoaIR5HflyiUksYjHILBQ70wzl4DPNkMwFhT5/lyOOJ
faBbQMFCyC/x8N14kuFRy0PP3V2gD7S2GxFt+6IpyxtRJb1tOXWswghQwM/C
D01LiTw2KqKa8B9g3MJqTO6slJ9M7AXQjlmTVYsp+cxn04zoibNSa3zieTkq
60y23QFVgsEmS7Y2Kl/KMwEoHLqvvZPICuqhNDpWrObU7VV6cDt6XEs0BL5Q
4KsJdRaPoVTXefMRCI8ENP0xIW0jSqZ8CqdUED9YfqyIW+BKyvtfYnX8bpqN
cl8cYHMxGeVEwysGUjwOaqOtTjgjDI7bXWuuIBps2OnHjwmBYkpy6rY0FwlJ
ECt4hQnc6yjQcKAG+QZb5brCN7BR8kCk8SnMuDCdKpvN6QsqX3oZVOVVes3L
VhhlPcc2VAcXJvQH5Pnme/vechU/SUPZTeKOSqTFt0L3vJFpD4iRUjqP5yU6
FI/ATBC/gjXAlQnVKsCH9BgE+itNqaw9rYPTRVWwK5XRDyFYsoLGRVUUAWb0
zyczWeCxgxHeVFrB+unEhZomXPhTE8KtB3r3DVPz4aqD8ytJcsrV+kqwOBne
I1JZiS+i9RtwdqeXie9/8CxRoaGKlhjyttgsFavDwFu5qOMi/gl26HEPh0/i
mLZgwkbjQ3k2zTumi8aXDDXQ5Z1LoWoz7edx+eet82KS3wXbs82zxg0+7a09
ucY271RWf7MrF/ns/WXErTi+y2QCuqpIdT85G+untNIQozTUfWnvdbG1nvjH
bj1Z5Xd3kzrqX0nq0T5WGX7hzbIFv5LE0DsNopyFLXanOIDhNiSe5C3DfJ/W
qwUrhSD84cAbL5BfD1Nqube7ztGBpB8QIDZfC8JAHiFSOoztuueA4XbtI7NH
5YetAdzSRxZvpegFgBl4yVwvOeJBj+goH4QglK6UG0aToHM460Q6EvFGRkib
YOHw6YkwkFTyyfeUdfGsytBQ1VXuALlQbjBBIjWh/fmVHvAJBokj6hfPb8Qj
d/4q+qAJzjoQmCwV+b9BhhpL3V/lmftLrJg51AbNQTIp4bD4D1imnShTfwhg
zJDCk+EwwjkM198kzOiShbJZ81metreF5WGyKPA614g0EF4go0b3j3EJxSwR
byPTQYEdTqOWVq1GHmw2pGY9oDRcrrZz/Gh6eD15N3x5ViwhG6NyrQj4oBIX
8xIgK4vjhskleQf2SBxhY32KXrQfaMCxmQ3IZfAEqvshhpcq1o//SrM0zUxa
aLiMBMj/Vkj7iKWaupCdMkbmrmRF80N0OtNGD8Llt304Srh3g140A1OtrWGd
ilzVkNjBnSFJ+vn1NsUGss57at8+KSFC+vNIZyMTBv27aqRHAPb8d7YpHSlC
qPEOAfp1z1RAsFc2dzpULbE4GRkqt7mxuUTHwK91d7SjAluXJcBuZTkea1Ry
a6IzJzEwy3MOkFdyTfDE2YfQOzCBa/pWHsgRFPPQz25MwpjzuAvcp3YKPNrM
2pRT26GHA9mY5oDFpql+yNxaypnJrJbaieWQV8y9euvcoy0/Kz458XSkK98b
j592FVhMMSjSMJ7ZHf5Sc+xvm83WDFfKlKRY9FJImcb31V7x1HU9nMuOIqV/
4LpF+I7HP8t9M1NdqnX2hgi8Ws4AKBBo0DHWaZ20xeK1q3wO+09nz5HMCKm4
JPDGItbQbjft0yh8lvz0zcYdq29W8LR/FwZm9Dp4POUaNtnyfhW9ceOmWb0c
mEjRVx21jbaZgrwx5oBZbPoZF+PPk0ZOPKfz6YL/40rkW2JGGFTw1Pazp8ta
tbjSZOUOUsM/VyYV3qAwiYiCwKM7OKa6ePC+b/ltLpGZwD7wnSoPem6/FaF8
LihxnTTA7BppJLWyjBk6oxDOsWMK8DUPIb/ij/hYI8hfrNtDEnXqJ0I2Q6CP
CezIr5IEkoNZ6XotW0RIDkqnL6O3wTHBYRUHotATmrzQ//qquunMuu8KEedC
z7zocIK0Pt8ikybo4o1n2mkpp6TVbm8Cdi+eqhb9odGqhjeyCtWjeXiqRd/1
AFHmzJqSb18/Xmej7IKdCH4l5VqlItIy6IekjXOvivLSOMN4AzQR9cXfpaeK
PgS/IPyVCMnrRdCdYL9YwEEv26wBm5Ey3EGoZutvmU4IpudZyEQsKFX/17px
OLAJbKVD+Jtuc6CIDrVw13BE5q5LD4qvOLCKT8E1L8TxSJxfCsa9GC5cwdZv
439vewA6E8VB/oX/S44/8zJiI7w7jhiqqIbOjIAMEkSJ9zCONXrzAfndPdPK
2WGL3yFzz2xVRcq6FHiGv4KSnpeyEg6sWgfcKonOdn07P2TL0igomh2/aIiI
OXtWo78PLxzaIHhP5JGMZ7p18tnUYO/RO/k/U/0iZnbsCYO2Do4L9ejglCVl
U3bgkXLijNBqtTedpQ1FX997AS24kI3XLd8Qhgclwmj5IKZPjx3Bv4MTdSFe
W+/syVX7ITpmmz56cC+/wBr+HZwVnXxXWSK/Wiv0/Phv2V5Zr6s5gd+BDOs0
e9UEL2wH4hQtR5Z8iK9Revq+eaqAmMFfo0u2XQcDbZVSzJffifuMWW2Rb5fL
CmRU46b6p0zAxf+rlDhauQ4v5FXp/qJLowzT6ePejcj5IHtHx8TZhH98EcO/
eo/bNntxCA4VukvI9Ykr9Nw94uE5lXdmWrq0seZXPv7lPI0xp19D02egXJ3r
M2g9PjXXcMttJwdWjOYzlcNFYSfsoEg8qA0dzYdskMd7npLh/b5aoFhu/8fp
xz7P3XUALUTzQkUK43ieBbsHJGMFu6JjYOWPOjo9zmvWJit4iWSJTFjBDufc
C181Lyr6pOoQ+qgND38SMpjGXlRPULDrfhsKy8/HXtXvzhOLS+x0pFUqw/GN
e1ZKwj4DpvLKL32rVS7Rfs4YpxO6YimUUfwRq07ySBjzYAXo3+P5SyPfyBMO
UUY8WV1eI6qtGjIs7uyflKRUL3Pvw5Sz2W2s4slPkxt9N2K8U85m2Wwvb8Be
nAXpV8xf94Nhde3ksXCpRUHtEhST6gVIwhjtMhX7LHtAsIjud08IBQUAjE7G
XMZIeo6O1h66fCOLiX6unRJfoQI7OO7dKAGJnAdVff9lVz0EsrJtB/v0oieT
tbrzqqfH2gta3/+pV+T6GMegj8zBw0G4PqakyFsoslYgZFNEVJU8Z42al1tS
Nyu8l9a/aUDfqfA10elNGFrRUQOhhDvC/egR9MlJhhGd6sNtQOGEAH9vDcaZ
Zyh/vaU/HoBIRp5Vmk+51+ZfHMt2DsuRADmO1J6V52j7aQeoYOmoFMble8Z2
+qNXE5m54wYOlzuVHzGmohdqzgII7aRmNRZeCQSJMbCmZvMthfcoz9SvZ2bT
v364J5a2LwVk3SJxDLZiQ3wMmwKvKh3bCUvNn5gG57mtnJv19kf8TsyREmzk
6G3yAaetBLFeM93iwJ5HAvpLfrHoJntUMnRR13kaov9bPh7CoovkTGjP3XAZ
Y3Do8Q+w91BGzhp2tsBdQXf2IXrxZs3haI3N9kT3Y8pq9tQ9hr7KbL0o2VgZ
h3RAn65Q9ZlLKUoFLjOucUUhW8OHXCo5Yfanq19rbX3vFDtTMMzXYJT14EQZ
xb34tWNrV/mfc6aMcIZ4GzUQHSca2bxKedepjiDvzE848oi4ZPrYDwHnMve1
DuyGGFcZw8Le0bekUFlyuz4PXoAkt54FcqM6d6L5oKQvV6ztWYTPwdC0QaWm
R2HmJWIHQfh17Frw8++J9fIZ45bXLN+f3gixo/nd841o94lGugShvJiv3QNc
oH8SXVu4Wh0Kb9rMq2BEtt18fSPj/ZOXY5vAlRqKjgRNIfhbJQ/AXNZ9HZ90
X5RmN+WfdmERWF3FprBTatfHxGxrqbx3QujQWTpyuMQK6zEOKBIcWYQ8dGwC
NHn6BW/wjR6e60pyVkGjQXsTODuzOqERiDDkdv8RoDUv7xyCrs1CjNueuNey
RN00T2Zhg10qiFNraBI/T0OJc5pSNygVoc0/85+KGuhsS1C8MgzPesg23Gp0
SxPU0msIFN0tuhNKv/+13RPP3+Semlqh+V78k4b4HIO36omFuS7sHN+XCxx0
kamLK1cgM840wqeJzlnWJMzrrkAVGKzQzaMpYiH0pmOSe4JYkddNQLm4CNtE
vXV+FY9h4BuFryVrfxwEDoHq4tGmSo3Jdu1eaVfgM1SCe+3OLwrYAX0SgDJF
rLagaq6vHjHlQQXL5kuKND+A8xaROUiN1pr0qoPYzD7oUsPyhl8aJTEPCpdg
0RaJYOfynTp4YDI7Jamna/pKv131mE3x0ztXtnVtuumR+ZeAYHL8Pzx8O6K0
0IZquFVLEZHjfZIsDOIUQYGR2leZwEJXDZGru0Uofj3bgjlg1fi6gn0880h0
Wu0zI8kmi2hsHUGJSxG6tVyavB+HW9Kv5nzd6RHqjYAnThjxkwK5rxvo/5q4
dn3oUk1NwyTQFShbMbgl9U3QrzScofCi/l8qkVWHz3zprg8e9sUm7917HUyM
Im+WC1CY4M+syMe6YSLM4y+HFw1jyPL1U0CpaEChhEbQCrPGc813sYK8ERvT
49r0NKWWBs0nk4dZo1pTr+DZX9ZmO2+tQWBMRexJjE95c6BpspT50KTT7Hu7
h/NYWOthJOMj/LKPw5jjEvOgORLmJiBvkON31fmtEhTVfXOSZGEuMf8CswFu
NwIHb6jOTF/qx9EBw7ZauU9FO1jWyrIxBUA/syitDAlMdyWsdKxhu4P3RaqG
zcs8hBKkSrqqh5vNj2q6ZFxblGAisdY7K6Omxeu9ObkYYZZ7EPX3+2ROZqWd
O9ehpCVAVFgYCS4HoUkrH3Tw+WhPuHwVIQrTiHJfp0nVjRR+FQfQj97daHsu
TAWyQh1koMmw2oBT1Y58Ca56NZdlqeijO+slctkP3QAh8GyYA3cMp+Aa0M5D
NVP/fewRnneeyzi2s+GkC4e+/Z20pxE+WndEtYTaCKEr5ssX84cuYzj1071Z
OVnczevC2kBRRVWh6TpkGLj4HzMFNUJkc2NcH7j+7fJczwkUg+GEkGeBNp5u
GESOb1Jk8MT78yMW32UBguVKaoVsZBUTLfOUvCptlYomxbfxSgwFwnkCJMTz
Xus/NoW+cYbbhgKOkDXVZ62axQbgH1mi7KHefQVaPSnD2Tk14+nkItFZhO8a
IFcGJcZiJG/qlT7ViuwuDwvZfeUOBDXlRakNXLUpotfbZF1I6tFRGeoQahvy
P8pnjh7f5ZQex80tuHDJdeL3nX6oBwOo/vnSa3XZu9XMVBHc20eKt52QQYtE
TJp8Ku2jscbbXsaluuN3QNsICfO8w+m849A17XF8COwhHJRmzrE5glNCWOGI
Ms3gCG+X0zqVk6dvNspUpkacu0HraO6ZVKB5akpLfc1EWCd0eOapjVhbUIgY
/qiK8AdtHylhNdLGf+vUCdiFqPTTDGpsLoX5LU0rUY7cN9tvvyUl07NKnzHq
PTbyVOUuuiT5PdWCxtXnkpUKolcfFV65Iu2zwQvvM/TPMAU28jov7fhXxn4X
maMLrwyEw0vvJtSw/ogEu3UmYiR0up7YzUIpEwVUrny5kyYtCqZn92xc+hAt
GSy0ehVVRMBwUrLzyAZb4dXgnR0cXUBR/TJEVjnnGfHlujozc1EiIU13muqe
pac2wJbv+IZBt1x5PBPTBzLvlhbf+YNAtqwa0+ZrFo7kdrTcP3x0gMdCk7U0
zjOvIbIOim7lmh8BPf1HwisocjQGON814ka8jk61sfkHoVtJStwSwrLU885g
8/40lplU/eTbmQ6WGbW+SRTkRa6DARXBCB28oidt6kHPvoZbWe+p0nD4jAke
uQVL/1kwkCN0V+6OF477rYCg69S0N1P6liM0aK4D0MXes84mi/HM1zeejwtM
fIi2U4CCLBaXknw+HnWRKT/gbK6ukt8kRVCnmbyIXXWmZPidmFYdRct1wkLG
cggf8YxjjYxYOtizayGwjiFH/s+1T0AWXE+pongWWChuNHp+8uyClp1c/WEM
X8HuIhs7DmINp7chtn4NYaw77A84CZAB8g2lyvUqWwttuCr6i/JOID96ivsh
dWRdCVda1wO8VWvEF+NOeAbR/UfXmT1OlcjZX65Un4CQIY/ICJn4qjgPfjch
qdXNE4G35boEvLPn6QYcgET0cZbpKFa8269L9oKuzXErb+7nHawjYKVe+hey
TLtP8Ovsml9z8paCQU/4krLLBt4K1Noi5USMJyXP9Fio7JkML2oYG8svDInn
UseXeuVzw0JxyycgQDFpOsMMnNfJMhV1Fwr2tiztJg3T3jckfxzMth7KQdY2
PDpIBVytCdC1R/Ozkj7el0EYc9fksjo8xKRpDEbnEL82XaxmsE3BzMwBX9EJ
EEnUc/H4r1vDzxEOiExmtMyGsuGI/+ehQyjXMo7+/QAD94w2AMcBRKjL87rj
y+9XiQqlHX9mydLHwTLBW7Cu4PzsGWczaghycIFcRLGfo7xOODtiusF6EmtW
RVS3uoHjOPkxRuLJikR2MKhfDx6vlgxIni09HU0BDoWS3tz64t4W1RLsE31k
Nc7iu/OGIzJ9T32hYLPWSiY4D+EfBW1TKv3SiW8wFySBIBy77b16qEDTy3aU
1iHudYrBMM63DZ1SfxyPnLZt7p+okSrhSSsc1sOjRBMQnDeL/7nHdqHnt+79
kpn6EtZ+xjmqUnr09Huu9nIALu0an9Y9t2Ve6gLe28QvyNs3/A/2oPiqDBYm
TI1GyI3nE0lO5aImdYSselW+ump61TLhwS7cDleozpUNPpaeAupUodGYFLm0
t35tit2KBn7wP2d5inIW0ihj1H4Pen4rzaC3djhdl3aoIcINklh2vVK4orCk
sN1aUxMworuVW7ztppooQ7a/HLUXc1x/jqfc7wfT8pOClCCHvcYzGU6phiU6
o17IK9FGE4lQuCieBbZozREzfr0qDK5QzePjIKJgCyR0Yp+UaJ5UMPB1x6Pj
m/PI2Pnkh/nk0GiIWYVegxys7spVve4akZAeOBoJOY2rYN2jPFobT1wr/MT9
/aVQ9IABfZF2efRMpWA0sZGt2e7szYracjH+OySXzRKNO2VGUPP1UG2WP319
yQ4yB+I6FhpLA5yNbRmieEv4kZN8Glyn2w815/9FK0L4B9xVNemYO6ZCOLX/
eyffRp8x6B8FeKn1l/qBpeCcaVwakEiFeIXBWb7A4Owl6vebqdzhz+2UU60D
LOANLvHeE5R6PaDunSWBkrmEVffhk5hS2Hg9I4uPYqY6G2zklh//NTOlFfGC
LGrVlwbAyKPRaoLNVM1seVtc1/mjip0riN65lqJJc+LtvaElw2lVTxqjGzQZ
xFd05cIvgbVBkSTS6lrqUFHLB68k10N3tdjBvUYkpSUUBj1CJgAFMr9SxF3E
WA4CiigysQRbznn5fX9AA3CkNVUmQZHmQpX6OaiUxq+XbmtAsLG55mNs9bg5
s9X3VaZ+45fU4h8ktBGd/+2SVzg4nDSLoY59Rm+UGRKkoahIvpZkx2htipkw
8MIHDPtwk/SCdHMMcAxibQy59lRGU5ToKaeLUsNQb0X1dLxskKR6WN2oU4AT
zE64k9rFitShkh4sTeHZnpBGjWKj47FN4pq5xXTXJhgOL8Sh4mJfxZU6CJSF
xKffTsrme0NVSBE6TLvA3N+i+9H+O5OBcZn4K2i21s5sZHHHd1sff1qEV563
VrNcYDdu7wgN0iNno0AXs4hcIJo+fCpNNSeA6Pe8EGKoQ/7GISzzKYF7sfcb
6L8vxTmhJDKLqH50ypoQP7/zGDOvkHQVL916n2EXuRKkQptBvvrGKtxDxlGN
irNEDKEtpn8Oa4TS5cxhuWzkwx/OPgQZ9TtT5iyyMSJCQ8bbhcKvFSmtsvzt
vXYbJmJTQ1lxhV3xZSbR8A5QJdvlx6C02zSyRXV0aVv/qfI1F4N1MgbNsZzX
pQKvbQZi2egtpWCgXQECOkaLriYZ3qo/aJoUwj2+D6MiZmGXkASPSUACrUta
jXZa+dlczxNxh3SlYQqq2OnQGlwTu0Xy/RR1pMZv0eSGi81UQn0mY3meZ3no
4IUV+idf1x7RTkI1cPc4MWSvcK/fpFFI9AYmG5OAgXosodUC4tYvzyiPmdEC
mnpuB0mDCyAS7BkMEjd7r2eY6/TYN577lZ3h7YBePv4EtwJ60gQdkcB/ERYI
OsOpjTulLntAqPxsi6f0DCagKDle9yXmLOcY4d9VzSuvavgfF9tN9MRO9auD
ZRebAmNZBj2noOjS62EbgjVjrkaA/Wtr/aXmY3itnNtSeKpEv89FeeCo8Ue0
37NCKEpey3tPb4bT06F3rNZl/JWMZzMN9zm3EzmHHmRmmQ/MzbkckbKr3VCK
4UK/SgYYOy/frsvpzt2yy6n59+VYZGhx5ZI/mV1KsSlksaAwTDTGTRWQIFCk
8vt0TMmnJjAamVo6HfUo0X+sui80sFLfx1R0IgA/ya8QfDAbXsE0BJKCHyAl
lutw/aCY2A2GYsoBbzaFO2jdJtnlIzrdPnIkEgIk83o7WDbJzIEU279F/zZG
HEDSmIvEY8ua1aKTnqh8c9NTgFdKBQdPFu0WvZQBh2LrZOxvCdu70mjasyTg
M41VVpvMu9qk8LanqFY85bvLjINCnypWCDiLAhXEVqQ2HDJy1w5Si9p9jzbQ
0i0Ax7E1eBQHfG5MWM7Qy4Vhu2II66gRJ9bBAZYzdR29gMS20sxwlu0av5ZO
NmXOgLbIQt4VnAK2WNXk7ImVpv+UjVNfAC7kprMBFmyP56x3ymbXIAMveZHs
v8JDrT1aECo6ZB3mIHdcJj39kTjAbjP3golC5kjQv8/yJ6EO5CRDRSccFZQW
3l43dMD2wEFY8sEGQcExj4kJzdQxw+G7NGo+5j/vLAh+ucDpqCgTDdtwK4Jr
Ec5jLTmaWvCXnL3nkjoKpinQKv9/tXBdMBeJk8hGRJqYfYvJa0dtu2Q0uX+P
E4bPEiqtndu21NO1ocVCqWJUgFLJ4ZVU5t/hGC0cuPZb5fiuf9uviW3Z+43q
+5wGnC4k+Y8HGGBI5ywaRHtFJD3Zh7Mq1ilQDm7YvGsuCdZIEExsikJnq/N5
OCRJY5cF54LwiH921mpeiqRWGbmDN65yFfHExUl8kFVegB0+V764SUAZpTGO
NBkFGdR1ryCWZiEb/LdSY98ROkTXmhp0bEZNd17BBmbvr8r+Z8rOwRIG8LQ/
jCHwSMEgvTeI0gNzSmnhjFM8A9rajMXvbeqMUlzBBgoeMkFudaxIloUBxdgo
P1iYv0IaJXMGCYH5QG+xKYHQKXF8Je7FHZk6tOXi7rx4iJGZNwHHyKctwTYN
G6maXDBctNQM6sEF8S+3/GC1B7iTA+RYju/iKxZUksucNyRmJVMz4UQaM+qf
dn5jfktkaYEZjpYedbK8JTc37SzJl5KpR0P82tu4Ixxiv/MVPA6Uy60JClC9
O8CsMOzKjOdsEZewjcASS0ONyIq2GZYxTUggpYjENqd1buq4WhY6reAeRyHs
6TSGv8MrTI6cp7cPA37M3bo2dOxxaZ8GW0cFXa0EhS8npOTCoCyDPgb+1GJO
BfdiOI/n+nwYZbfip7xrfedREFUux7M/L3j6u5By8ObNLgng7F8TYt1S+v1P
ewSgCFKy6X8U9qTiG5PegPP5DzKWSEGrB6DpESv2eHUt1Vailu2t8eKzYOyt
a32STDudnA5w+eE0vv7Xs4+wCit2GmZmHiJzyAucvYQSL20CaeG8/tPaSFuz
6YjUKE7ZcfIsU04iM+2YsXDgSPJXHZntVejfiFDlewRrFaHeicGFJBocH57c
JmbOqIpgnoeEl8EC2cEyga2zoXaDYgTL9I4pe49iyHdhQuYnTgoUhQb43+QN
yFc8FHEdJhhFgtOQgV/ak90Qpf6BivQGK5tMOHTlxOdEfPxQjtx7I5KRCPQb
HnYKkVsu+usd4m9b8Cp++1sEtkW/aVn1vZx4OyE1sSgWTWXNWeIv1ZSz73LN
qWhfTIYXgE/oRWRHpJXkX9+hDC9PlleYHtKZwfeLNc0+5RWWL7Pi2oEvour5
4j62/Rf0FKwp6rOFv8BC5V5wMpKFLGSqcrAFEc3WnkvEli0bRXBmRXUaP4cU
3KfIwmT4X0kYonyAzooR11hLpfQbuYaQkSxaX5IMNz1J3lDTZ+7Jq97SlhoK
ge0LH8MhSOfz2YhnLF1PX5jYIkaIIboYrtXHNvELJTvFyOUKymeZcrud8+XB
h9k7VMToTLSl06Da0RiKRsslZSifqh5UIrd7Hmu3peA/8B3ulheKqOp4TaQe
xeL6lg41+ywCL2DjhXHSCkh6z5KfzJYoI08akbiiCrUglweTHffNeO2DZAE9
/V1QQW6J3ZCCqBf8d2ViBiDYQEyh8G6P1MZE+XhmrpjnGUlE/qBk/iuzYlZ7
SU1i33n0/Sq24El/aUlcX4oZvgjYCfOB/h+wnAFMqmYBqHhliLV/1TTo9Ofj
3FtpA1y30FS8PQDJ/+NuUsUrrvFSlctey+LAmwOjCRRJkzy/93O/cqfs0OG3
gMa51FkblhfQQ55+but+0yDGmGipVjvMO/oX7E0+i49OmSCYLbgJqcIZSMrm
HJlB6B7Eb8fjTlefGYmJKcFn6I8U0YnCo5/3tarRkMXS+bIWi67C/Tz1rC0P
haA47wHuljF4+zBUSJkMsN3QMuot0MF0frEsQ3Qv3pwbsjec8Orj/eSTxYyY
PB0pevNOA1Ui1t5LEhnNvkhaE/GebjkX0UjmTX0vdYBEzGpvH+cC93Q0hTjY
THuMNQU2Ja4U7EpMVcPYFbA07xlUiAlPoKFT8mQcJFoKNR4Ai7b0OJ982ZcA
2dn4VKsMuTUlHhmmt85NlJO2aLx8QHrKTmyIZgY6PaMpG3mXy75CEXX1iGQx
iKQTVvMidgymi5qcatEfnG7wWc2ex/b4Zp8AQnRIlesBsPU1annxKIrQfaCB
hCNVdvBBm0t3e2h1Q8Aw6Zjceg8X2cFLmhQ0Jo3XOjVd7G3K7UwdCJp6de+G
4F2af0068G9GumIvEYaZ+xdN56IwRYnmPaAzih44T4lVj4bk8f1Ea3j9thJY
JCi0G5ZbdMcqVKHYNXPYgYivDOl6FOVtk3wvHpQlIvGRRDO0qiOhGU4a0fCv
gUQzATG+IvBTF3QGbCUFV4KfA4fTSorbsksNWoFuAhzCx+USNnv/LloANawF
CBWv5jO3zhgRytgnDigAE/YBotAF5MY9ZXszj2/IKYAYY0/8IJqTwGS5njNa
6kjcNGWCmMtx4YLuIoihDaxQ7ipojmtzoSOCrrwrEjrdThd75W9rCkC4hngF
rzJtTU6oK4mdDigAu/kZmyfr7FM5eTNvJXBvwa/WFOFRyL0jolXwD/Cjft5K
yQiqyTA5ObbvHjM+FBFS1fFI7WRzvDbxItpCnJfWL+o9Vs8zQS0q4j16h1O3
lkSlkG7vK+8IVTDV/KbGTaubVy8r39Q526h69wnZuE1h1kDSVq0fMb8Dx3fR
BZgUcy1+Z+jtED8Lu/M4sKOkF3aVeWcfwzQljn978TgYiTET59VXoHnoc2cR
MWrv/bMTe8EqHPzY/JS5jTtutzfl02PUnbAGD/QLMDq7P9lAGUHrrUKqh7rN
vRlXqDn42I69yrEgWYy3E4WHwRzyzb+uYOd5nwDo0wrMcBmeaKCLoZgO4HCo
GnjLk19hE5e2vWiiPLJmDz9+NG1limv23SkHCO0eMNFgdNW0SmOd7hZwxRby
mmpTTCTGgX8dOpC2yTkbDvN0ThMLyKlCnDJvZFQ2uLEgHaZ/OUhhRwsQmZTU
cGwPqECMP1ORTFD4QKLl8p4gjWGllaedEteLVDSYlRJCUy7xg1vv2sD2B/Y4
dTqVZ/9WvxsApr62smv5PwQ8FH9bDjNjyaZqbBFwodKiqc9bOjd1d58vl+Sx
La/rfXN5peGCa0nHrgAvKq4Bs6UID89iVfgpG3o3mATNZrIr/Qr8bl4KdB1P
YwaZyzKFvVL+viEqt1/OZd18fmwobivZu9YBSpWg4GVT65g7sUmRY6H1sVPC
mSkEy7UTbJy0uL4AY7XYg4YFhxaSzc+P5S59b0yDQDuHL8CWHySEYmdRNDmf
fFSw+1afFbR1aR8Km8xJmMFEN7+G/RY5jIDkXBuCkb+DbtS6WR9kD5K1F1UT
KeifLaZkNKLD/GhUoDEcILEEeiNRz8xkRd1Xw4gS/t+e6+4NYPTC8eC+w2Cy
pdpQA+rnOdgurNISBV/HMnIY4NTQoy3nLGd2JyMeqbU5N2STbbo4aMN7VNPV
Aq62RGc/hMUb8jcXDKWg3PyJzStFSiWRNtvgnUle6lUEskT7gvwpW/WyP089
gR7JVN9PYY148OD4VcxzU2Gva6wX4ul/257jF48dDcasJ4Dh3bOo/nU99ihd
ZALv7odI3Hwj+cPnhSbiNyCvjM1FmfhcrN97TycJalJFccnYJQCnuqZXFFO2
BliEejbCUlzVIyxM/01UFE2Jvh8wft8gXCNCW+gmmBfPTdLqLmOSDFoYFAVX
Ce+P6I5s4dZZSRTDAiV9zpVTCHtBHQGbcQPr36dcwbih5m0eTEaa3PioSe0r
xN6eWGe0VFJSHzVHxfbjgdyS6q2Ez0dhz2vfA7ZeGospDB0dCV7B07qQyrbi
jrZwIxs9oc0pMBsAbaWuOQQkt3J1wr6OBN9CUOfUtJWH3J2x1Dv9r2VNNaQx
+TaZUstn1hTfBXD/30ZaHiBHkqiO4PGXWAG1bELVoUj9FpZJ7YsxkFp5v92T
VNRQppTqeq+eWotSR/52ia3nm6xYVAWlXGYqk2dmDEgGRxyePhyXxL+C+QlS
gryP8eQibM/LwiU8Vd2J5+aWOeKAKqfsmBSxj4r5FO6VD4wZgg1rWnb8skWk
bb97uYPImzVSKpu0uiOAIi6qFlD6dxe+puJQILdByqhHauB1DY+I3LoCEsKE
tV1dULw/YNzrHbyCiMavcu+kV6L3TAL2GKHoVItiASWpUHDm8aztLHgpaFxE
P02HoZ1HohuU8Jd1xYmqTTxhbiFQcknOD2URJMOBmsGVN39pnp/UMY2vYNzn
B8o2MUVQiQeKFw4WsYW9mVpWTF6BkIrZE2VXVJqBZM2ym9GqOoOaBwjFLSf8
3z8d+JY45DsJDSuZPz/yzTSufW5CzVj1IsKB/GrLtegAzsv3rx+2gwRvEqiZ
BWDr3KSUgTkG5K3l2Ls7rwRoEH/rzdTbCbLJe63AhnaQ25H+FnSrsnGl1FqD
BlVHIuCSrG5miSL4Ak2m+HS6GCpFzTzg2CWS97c0p29KdRTFQrfTTzwGcEY8
kyiWwWSP5a6P+5dwZ6UmopXeDbBoOouaAmU08cPxKTcOK4lygZNgk8G5ZPJi
DQEwPCNsr5ixv8sX+vcW/AuE0rbkBYu6EsaPFuQgJKfqEb7u+exTTXIS+C9a
rrpbNQ1Wf1PRKMFktsEc8hJ8RA96v/BPbehUUaN2n5pClAkBITPVB4p3SqJ7
gnx+eMl1FgSYEVl8oGFm3XC+D6rkhA3O6LYjBdqfcz6YAikCNSUKhKhmQfdH
4rO9hm0sBO/oKAOny5po7yQwnynClcfINvRtJcM5F1r4+wN/gRdfBF2KjXJX
AprWe6AvSgCj8vGOaAfzD6LJJnlGpNY6Va5iPPy4DTa0ZPKkfFf6xoxInbQV
5AyCIsJ6j+Nf/aUlEht6CrknZs4LsYQ7Q4DvYmxhBbaCbbBHu+lSHYsWwRNg
HKHx6PO33H2om8mNEFwFbOHzjkLmlyb4cimYk2DOqsFZZULD8n6imfC6tnln
lFfwnnXZlYgBQe3+G4txw8L6OJADqmU8M77LbizeZJS+3G8Akk95olz8o7HR
I53cT6h8NAJu5F4CS8jIPPB8TnlBEzAP46J/K1kbW+3BIRCe4CRuJy4Q/lYn
wsAVRAW+EhvUzf0G7H6UFe6yFpw2xaBC7HWIX8bSCwKnu0yzSpzvXm74pc2L
Em20HxDPbo0X+CEZuQCGAGJUNWiQ40/brB6B+0OzRK+zGOpW+tLXwTk6w18w
W7D7gN43T8NHh4HSOnt52uOjSwZ3v5zSPquy5xFrEsVpCDqY28FR6Sj9Nd+a
cbSdI54DQuiWjYTnPGSsUsG3TZsUsW2xY7Vfx55ke4qySCFmBJk7HiWolxAT
lx5jgePST/PeGk46IdIGOBe03fjndOSIIpBzK/wrPGlNzrl77e82Q3qGyLG8
gS4e/l6v9HhT7qH3Lr347E0G9+iqQ8kKNmkfrKbQgR9xCZtDMt1yVtnXme2O
McnXPw8xqdkGMpJSfZUzOtH0T85cipi3jdU0gxuDH7yYLzv2reQSDC2v/HxL
M8LpmPXw31wtOdgkFRgfF817dXVSx+Y3NXCr8r8M5t6rw3ocrRxZmLrDQI8p
k19WUh79iSGGzSNlghTYiowDJ2sZ4MXA4Y8Foof5nuXzr9+UKK9cKgkMRJ/O
eq/LRNh59j5gVsik5ogmyqYBtC3zBf/xkMwFilAU3om6/tPXolxWmNuBYCAP
u3W9zolpbFRYM6qNLDFXmMY/sJbTRa7f/CXdXNkZX0LMthYrb+1lSP8ywq5Q
elkC4HWuSEZzxgPLjAp/sO+ExNfPJo3/F7v7ao3mmKZMtioeb7Zd6W2IRzF8
YmhiDL9TpL8ikd9FPprqVqgm8wINg2siuwyxuKBoApcXnQhT64nd5gBM7VG4
ffuKj429Fgdnn/rdwIDbSHsw2jRax41fUvnsxo51UHro/z9vMelVPzfowEhT
IfoZPg/+1yQ30N6Eyu8vZjyXHU0j15NxmsWvtwQYMXO7e9vfMfB0+YiwfrjD
zFGeBiSPnGszASVBxusyNwCuz8dyCSaCQ3Su3ZFoxoFZ1/nxZScxDo2idbwe
GEJ9Tjgf0dRQSqprU1OmjjklNsEgalXvjgizr2VBGJVcx0/Yhgr3IA7oVva4
k+nR78vPQXDDKHdu49svQl46clfP3ItH0zA0OPocXa15YYyRTJ0Cgk86f59H
CRK8MC9tU2yIylwN7/lXEXp0MUPdeRktl0Sa2ube4QA0KeomgJpoRy92CIiL
TwNy6IBGnep/9eJMRLp8wCA+Tia18uYHNMMzIp5ZtU7+w6ucTovX29pxHIk4
PBBqiJ9Vf7AAQqTrfqqyWZY+kcWD9Q+zxntaOAQKT3RgmxHSGL/Ky/1vyvL1
pN2Yx4tpx6joLpmQj/03MIXbYgdaT2Ue2DLXcZ93XQXXgRFGvTLomKUmE5/K
oTdiQJQeD0VEj/uqLOBijdJPcB1gY0ZltvbFnrQRKXSaYSxoCDndGBZzEomp
9lNMptFHopcuyKyke7VdZjBxuZ7FY3alIceKoEcvant67t9ZdSapMzfzIs42
62jMTQMGbwo4B5CeP3kilqBBgD/MjiZJHh37ZvxWVyQNw85PFF20Ui/SoC9b
GrVKyemwUKuN2U2DcDFvzZox+krc6A2pGX1o/tz4YK95DjxX8fyRjnLNHBxd
IMFH8siIWvLTneh5OxPjiMZ/f4DE69H+3edOItV1wya+5me+7/hvv3pK2apr
ducWc+Y1/tHEH3TFhvENbaMh32sfRXRx8s1V6TunIrmnRW0QU5zQV6PBZDkp
kWhOg8GVXSkbkPV0FWpDgamJx69WrdGCNbhKoJGXaw2WpXR3MyhqYrZFLR2w
8e35kUSrmF91eud8PaX4rGlI0dmlSNr4027HIDQX/e6xr/RZqfzXN6g5a5AR
QupNmy2w/iD0hQ5sN/WFI/hIzY25VmKjfpyiD5/U9anZ3vSMGQw6F/0xVxyN
y7RmxldaSuqp8+NYR9HeoVXAtZt4P6DlaFgAs5wGEv6ROQflJAHgjb4zTX4W
Qn/mdm955Mh8Fy8tHFrxPGlwuGPiWmdenn5fIdwvtZoUQzMbu/Ao/bqJ4HWl
sA9mWkWa62DAsO1K2xUpg7gI7gS80uTuqT8riIgVt3qFKMmZrejMRKA5i16k
qzbU9SKW6MYImAQqYSdgH90TRQy4YKfA1DHTe4efOuLyV49Q0aifUZtqyrrs
wmMoFerkJkxN5AdfpJTosKMEWEbLPZuTlieaVms8CKA8Lp7uHRRgdXHe7N4L
Bf8Hm/56wyAwsdYQP+o+DQg3JBhfiubnALx+kK2vkoX5zGdMiVcihyszvhHt
kHQFro3mB0a5VsYwZu8OwaYndPLydOWeKG+iVFURudUN4xX1SXM2p6ruBF64
VPyJb3nTTb2fQ0b/5iQHjI35NtD0OFi+1S/cELv1FmvU2NJt4W7fxfBDLKRv
Nmp0xNY6IeDAnV/IaAHk14AjVwQ+i7lAJho7ZIScSa2wYQOkTGSNiRxwzMGL
lXOLV5rYWwcAcCBvCppZ5fAbKIZtMauUWFDxVysQAP2qykT0sZALwYGsCEkZ
2sPm8ckVp6xgAsH472awBIChIbZbv0VKSLXwuJeirexbjQSPCt/GpEnosYOx
xbbNRzigjE5u3lm6GgQeRY67wGqTw+0DeFMhyP9pXRTzPJ5VmWMBCOdtPVqy
YL7bNvfkzdGYbI4xMbdg92hNM0foQfOkR7p5VajqKVtBkMCKSdLMI2T/uJ1U
cwnkT7XQgWmU2vQfUhYFEYNaZPAnn+Out3nSbr3qvuRENTTG7CcOLcKzibgO
lvFAmgftK7FzQmoDOlBAaNXQ/gmv6W/hfKCZ1Rfcqj+H8pdSJvADYzESveST
5Z440hGVfh2nAC/RxaVabE2AkgQ46g0QK98Rd9Tby3AND75BVvoexQL+ssH+
IFEs6VowHrUJMfkMgcUIcf7ZxvT29AfyAxWKo/LTbuJKRl0qcUNqJf+j69pq
xfT0xYXS8Q/Di/EpeWH1vY5fObrIGY8q3fCDpVpbRJV99ijzQdxCxHvob7a6
ZIQAd2r+u0EaGcVQdLRzh1sWlUAsA38iwdjw16xdZZOiEywYs1K01mQBQqMX
nQLDZnHsua5hpAEOgqL3816YE/lmp/b/zj1rHoveRiyOyHgNgy6bI2VZwIhJ
DwzF8p9n7n4YYG1CEK1f41SFGSUCdP3TntK25a41ltz/Z+iccLm67HZiTRSH
bl8SpU1Gk+8h81SE9/q0wm/cGQIbtc1gS7j04wQkeNsDNsW1FB622fS7k6Gz
A3noCmJT60slxkfrAssvNxQxJDKGzvnSUVppz9ABwAyCWu0J6ktFByjf2ZGp
LZUOyQjROvzEflcYif2R4X9qPbb18bMxdqdRGXaC5BgpSCMHhlY5ch4c9djM
OQX4QreUAcEXsyakLtEiuM88jedhoIDK3GgmKsx7OfBNqQCsHgig9BPAL5T5
fZ93DZZb0MMoEjx+xvWrCSgefq4sonUV2Ir0pXGWZpvBc/1EI5vhbgIyVRpc
ySEewJTR6NnEp2ghwysTs21m4YlgS34w1ZjWl4yw2LeOK4ArlbPsGNqEYG4f
b3sT0TYNDyK7ixjuOcqWVFTNMTAze4OAifF/WFwa2z5XvsIkQ8QOO1W9RvvO
VT0+5EFUrJb/aRKeM1+rCPLKmxJWXm9Y2bFzGbfe/N+wfoWlHb5S4rKMyXkr
exwsyPybweYMummiekmaiUGvwKCL2mbwUmaSR04+K2rp10nxDIChfoxNrcv/
VQzpYhp58iCokSk/OIVuYFWxLpVyiqKbnQvTjMwHS4flXp3v0xODmCAGfiep
pY4uvm5l9Zazfye1AotMxPCfB3E3PIYw1yUbUODbGYTV/uXHjqmmQ248uf72
6DfQqeBg7H0Wj4da0QRY3jvNEnMBKdYqMee/KQs4adBxXDjKHYN8QN5I/NJY
2O/1JWmi8iPbUtZKCQtENcvrbPGcQKRpCs/tT3ryhyYYv8W+vYcBqUQPKuk/
yWrTW6FUKLCw6Fik+nzKIVbFJ+1mqc39JvSZ7KzUizDFr3Zy/QwhUTcdH8y9
al4Yrel4YYlVYRll8tZ5v95E9vBPMdvsw0nwtUJKx758aFAYVD/uC4q29vZh
vS+MMOosrZESIGMly/86qrJe0fzAr6QN2PTEpXu3AsQEt02m9TmIG84WASMZ
dvSqfCPoOyVAD1s4luFdp77ZG2IT12FAR8McGGcIiM4WlpJkJya0squaaNfM
XJcQN0RjxhSf0hPtfQl2XFeC53F4WS6XTxlTGpv4SbCYigUDk89v9YgFVPWe
sp8Iphx1f36EZTNrJ1mEFOxZRWoMc0Zg+Q4W+Eo7LV8Mx7cI6fC8UxHCGX50
mEQHnXeQjej0gmqcajkLPjAtc3IhHFus+Arq4e2lwKC3Eu4TZ+NyqvEOymGm
O/iF0oCUL7tX1FqV8NJs6K2+N784djDDWjY3tY9z5fnI6Ne+k55ahE/djUOI
naqMq/Ko9/a+olVz22LHr/nwWFQ+1xYGASCVzy4gSJn9SJuq9R0GzsFmq1/S
4/PHcM77qKWbS6ZWwYfKmneNAs4l2kGyYEd1YDIOFeIhRmoVTdonhfj9K3eT
pLHLQItnjLXFdHU6YdbKDjFJ7jHpDH/baoKZTgDwds/3gwgmXHMBQuzjSWlU
LVxGqqQzx2ba9IGSCk4zxGD1vMff7U1QQxWYpKWxOvglao1GTkdtG786jls3
NCsg2zuifr8bnl/zpM3fIEPbMarVDk9biYKT0cxv/oUAp04ICUeemBNqJxXl
tPpZsR683JXhBLOKINNQu7nu9b3OKUCW9HX4jJacxUY/SEJVx6kB+3waVyGZ
Xz/DwQYb5k42k8dtq46S5KlQMQdmU5Q5q90h3et1twoxY+fuxdF7ZyKCLCro
QAsZtkpXZQco2EeG7E4ugJBVpaWvqBIIt8RBfAt0o3UFrKq9YL1F5cDc/Zvt
r+DwA0pXo/63V3/2oHc2LJnd+v9BuoXqyRcCkZtDSjz9B0jEVf5RsHrILCAm
aTIs1OKsM5t8dPyYRLoow7Fbc03fHC7Q8kdenr/JSQRBnL+wDGZqgBeax+TM
twkqDwCnPE8X26atnXCpQ/CVP3AoZXNszzd2a/D5FpjHngh0A2jYg1/AyXuz
xXc+mETsjc7FPZZYObXUIcpOKU054/2rk3g790krSv2Ed9U3jSDuRQTFoqGu
GYzzRGtPVYp0DhJsrOcaxIlPUO5uijx/5ccuF/Xque3mzpPEABlV6w5J3oUH
mZ6Kwo+Y5zEHe1tIjjXjG1GVz3GndXGVNvX79QIIE4RGE6yc7eUS193kiJdg
8dLp4d9Ybb4o/aKuYtls/ONCFG9Nh5cSu1reVO8TZbTqHVr+sTo7wQDOra04
Wk45YUGPg+2NIaG8UjSmO/DaYpLiVsX56BKim8B5/aMDN4E0rbakBhxz0MAb
t9paKIUV0w2VnWrVe7+kg7hNJyR3SzvPbuu7zm2ZzotXm+rkB4bB7EOI+VYp
c7J3jmh3AttjL+IlkRJ/D6sRuwpSuB4ce2CTkVtFx6KS2M+oTzgzkmU4RNhH
esxDKK28uMO32MNecd4H7I5X71HurMD8pkd5d/mw4SfNT//YBZseBAHBCl/O
CvfNdUsS2epiRQ4chr0dAsKzCKqyGZ4Q4TBloSSCT8X9wnkFGzMc6jWtrICb
enEGq3K8XGRA94Mx88kzNRcfeKUV1k1j6DxnYaLCZHR9mmHqwWr0HbmpM4/4
OEAlPV5doINt7enG66+Y53ooNvfgSwPXrCGydkQ1cOE4Y7e4bZg2EYnJb/1p
/wTM2hjmN6AL+b8bDgihVbtMzu55eBCtViNuEuFmYjdMThpSpPbGt+qVBbB6
rnO1z8usvBRvb1l+NXTl0VvTn51cxwA6tpNoa3QolJBkoO7solqLNVSqBvFy
HxMI8rS8Qe2IRMoxzmFYSrgmx+PxAPOnZwB/jXLRnjVq0taJJEOt0xxRdt8e
+vJLFRXmCgTO+kZjvZqXkY1Cz71e1YoBY7LMcNB3+dPDNDu6zoq4Pem2On9K
Eskebl5ZzRcdlguBwRyRstCyoAstfsP959hzsQNyCCfRceYEntCyMzyA7goR
moy7JLHU3i9GUx5NvKfpy1y19HZ7n8rHI9sqbkeMI5LD3+0fUO4HvqI3OWel
vsfSOpQ4Je73I2lyL/ZVVG2G9Yw/dNqXGHwNdqKR1VIuXyrktywIS0JAjRmw
+F/SWyqbA+6Lt20kBTeEYPJ6BdnHYKK+GUz/aqMnUKpE2oaT/0RqHtxcdKZh
ttXBL/+N8Jn9IZsi+ipz8H9cbi0aS9WLasxrpao+CePerA6sA8BodIDNrWEx
EGGA0Cg8tZpGVGTeTezgpiijhF/pBqXkMu46E+KPUVK52M9XQo6Q4xMHuTNK
RwPBgzQ4eSf2o5+5rIo+cDlTLwY61uCBRAgMt9Ui+AiuPSpfI6whythj930O
YTcAdrWY+MzIpLyWJpZf0nx6s2RSUbGE3hVanSv/kUiGpGSbLp9DIMi0JmLa
wn32vge52Tz9fX8qngQ/ukGH97kkyyQuvMpL7mCBYMXI/cO9ZhLTHO4RlltB
/LdPImz3mVpTR5oPBLhG4bqF9GCm5Ccio7Xd7V3dphA00n2PnCUhH6SerJzF
NFn/U3d6m7ihwEKfVpWzNSoRQQFKKQx8Vd0n4un9GTovMB2F5m0LRwnEfVAP
wlzoL8DZfryMw1OH50QD+NAaM/9G/rc/iVRdfZvi7kflBSsBMEbk6k4HvotQ
jwMU3K0b+MWhbC9DCm2M8Baynu5gVpuP93C6dMtPJRpIWH5hlH/zds/K9H79
S2qiY6Z3CdxVtg9M1ACVnMH3VbWzOCWGWazHWrn+iShTfNAGhxHIt7gCmYLC
X7DAt+znxKjoYFJAZf+YPQdc/eufDynAg8w6pNyRgp5gZNS24gtay+ayz1Wd
AXVW7Uoh33dUAfEpEZFvA7j0aVvHxU+wdlun1XURQp7WRZ8ZrYyTmLxAfLdC
7iUkhAQ0D80m3vmJ3cQdY4JqkcZH0f9VXlJPhsdNXryQqa5wO+eEvDXonp+v
qdBQADFta4hmxiMxHBZpFBTPiczUJe1qHW0ishUe2mqu7RH/rtpf+wmUIfU1
Cd/PqVm5LI0U2sRzwe+Ko4XCgK4vOE2Meet+XEx3ivzmoGHdvuMoToy4N2L5
6KT97WKMSZJop+obmBH/LtMHjH/G+SvUHJeTXcXhNIPFipr7JTSd8rhMH+2H
v3J1Vevs/iW48lQQP5O8uW8/zdHcQ9DZQfYslKj/z4h3GIaKjhDl7C4V2uyn
cilHsM1yNxJ+sGNubjQWtQua5XwC7To4ooxZVZThmVCDi1GVx28drOjMOtZM
IMxvDSFckf0SWlraN4VYhZ8ZxowoeBUguvI/HzNHOJ5/5v1t2si7WymrcPH5
KcfvG3CUznY/Xo23SrGBN57ykB+q/kuVBs+7lTRuK8OZS+BYdwol78OtflTx
xTXq6x0gZEwDp15/LMHp60ilj5P6P+QYl7tQu97eLhFo1j5GFzf8oFqwmiYY
7c5G5GsSFwwxjrvbxg8y78QYWz/lP2vdUFSjrUXuYYjOjD1zggSI1wY0TjzW
BaDbJbxzcXN5qQpW59ZOCwcs5pw5Sf/NVsszIo76tRNlUMyEYoX/yNlzswLH
436q91ZDjagqs5MTrm+EBon0Na8MFvHaRfiWSY4DUV8cU+va0fleiFtdWJXC
dFteJMc3BL3l0FSn3xU+Mwt68dGhW71+LuKf5lf8a/Trdq7tN2trYB4rJb0j
jIe+3scycpL0xgNhHcTklq/3Goh5Ovu0vTgpbzoUkJfB65vPhPIlaE9+w0NW
1jRFc87V5SUf2VHdnK669UUvxbmXNKvDe2ag9WkyVf/97TL9acMUSntBdQ35
veWqjKjgEejaOOw8rpko9Ex3+4UxYtrePFMwItbD3Fgp+86dk2rO2J7S9dJz
Ql4HgIuxYJ5Fn6TsU3iYsrM8lfNl5dH3M3SamFRwPtSWBevqyNQ0/62XKGH3
8a5Noonq/jKpvYBJyjJhtCboJdxh98peURuC6HL8cUfBd9KbDcKj1LG71lM2
+w2DjFIQkMQvWOBQgBT8oIrQDerplmXuMBizOntyu/kbt/sp8Ax2Qk38NViC
7ukqLn9Z95jfRXmYL7iBORaJ3RB3wVPc2SiHeHUWda2oBgr45+RIga0iUyUU
WaAJrh+ppW9WrrEIJz9yfljw+0C6/okZnTsP1YHtg4P1q8NikH1cem3/v08+
hmEGUf3Lf4sdA+NHrT+SMjNeyIBn3YFWUOMJ3h2at6Lm7dF7F8iMEEoabRxn
YtjeLU4rGRrClXipIlXT9xqNk/ncctyi4UFk+doOzvv/vyNTlOYbXqfYn9oO
ps2COVro6nNrjwMz83ZR/X0uJ1ywQnH8Y4RRGFFJFGgqOZ/u2q9silx+peG6
SF41wGgFZvpv36KF1Eg7YA60lLZ4rQWjjLeovGLDp+yrGGi1UD7HSZN1Kw2q
Enjph1wkKpGqxgmmlzqXNWohmZiD2k9pLWpWpQgKvOEs9frq5l+S2TkZnw7T
dll6SmsfSHBKsdgOrf3OivgkXvgfC5QfYIgL2fEChCQ7br/CVLFcaKG7e8Ko
hKDvk+oQ5iyFeMBuTha7IeCnuEzMp4gyBWEj4et+isIR6J3Z3NUYAA5SvJSL
RO4uYl+n4eL05o8oc+ciP+QEgdxsEBVpgAuz43Lk5eIIHjsHZEr9uAePTz6r
AawKFF5czkyspgN83+p9LJHq8Pw7JI+Zp0wk4jQO6wNp6ZVHeD9olYYLabu5
vQdI/u2i0XhoycK3eib4wlpsK7FZjrjn1wXso6gaN6kYYyodGYSeUlpml+l2
yXgq9hmFnQbfmBTjj+yisZTOvDM11NvG48emz9CUoZissttigo2UYZ9mJHLK
RLLHf6hjmUUyKsgYYGZvB9bLuEj9iYIpWqJ1Pf98V2PZM6J7WPspDNfxNkYz
VEPa4TPoXn3rBbgK1MVgidYZ/v1WRl+u40yaNNyHHl4lAak0yN8sWXmIMczc
gS3/p6sMN+SbWWUJsLz4OjClxn4MdkCjSCAEymuLQk971m8VR9Zu0rv1CbvX
YBLMRen3MRqlO1w5RHYOaBsqXLBbgVUj5UruVHzY8FSE+ddV4dhFcBEnmLPy
Av3cQKjeMFZncEbLQCLr+5IemeZkZ0/HfiHtBJgJ02umec9L3anNg07C8PCS
wMfvqpwZns/e/NpsKNJqd07pHfPoRBA8JUXosNcGDFuRuaBK9vpUyEIg8B6j
mEmeYXMLZXhTBjCzruTrg4mGpZ9bpSr3729N6imNC3xTysYgDvmwuVP5wP9R
VrrsvSzu/eh0jX5TOMQHBeDePP04V3TonYT+ffSfTEFmxq0uQqHd/dZkm0Jx
vBwA4TYQ8xEpPj0B1ObWpqdWi7k9v680pOBgZdOIhEzwqM/eHCjsOhlHZre3
mtZ+HlEkT3mK0hqZYrS0DTtCnU/kdfDE55b7GEmW3EkGRE0ASJLsDRxZCjwx
LInEGelJqdqC0b8uIGD5r6BiX7z2NTnj8TvO1PrQdKx7H/l1QGpsBUReU1Zu
HkfKJcwklYfgGTxpImtRr3t99LS1r0Aw2mmilYzzgPJ6/RqsvLt6e/1cneM3
rV4EoNuqvY4w1LdYtG7FAc9Y/drXtav/kczA7mHIWAd9AsCaXsEYxsBVRy64
Jy+uqn7B2N48wbGWIEBNIaLCdZrbCblqn56PiEuwnJCgPoS0nF1vdss4HVtI
ZDsz8PNGBwenDhv3aW6Xj4JgYT/m0yyfB+SaDacilR5Pko6zii9hYA/5MG+X
Q3x7dsx5xWgRKROSA71q/8k4yDVFoa104XShBwNEccNqUoaqRuq8+JwV7WXf
T2Gwirq00K2kZA7hVQT8XjYEwnhlWYFkLlKCOMyyQhCXEsCodcy2MeIGUW5F
/nhMweuxVp6e14C2Xqb5ngH6/DogXYABj+wfL94V4ZDZyuTmzIU2D3Jo/WH4
PMbbHMXQ5FjeuHAONf2Y5XP4qJJisg4a9VQ5176m3VqYf3uh7iEdXEJbZYD8
/ObK1DwdGfi6nbQWQdeb40mLace3wymI0kXSfRb0ifJVXZAqAhpa1cDnqWm0
VOCJ5T6/6KCcKF4b85K2lV7otH0Ob6B+Jld+0hPf+gJGtibh8FKmh7cnM0K1
zXdqZFyO8pdS6VRxX6P4Isa8OwxF6RiunZX3tdV9vKUYHYHrcsa6t3SZn3JU
D+FMJWN17bzN73hcyaB4Ze7qPWrcqSS7IDoKaTRgHF3B4dPw03sqZzyhNglL
ZgWiVGlceEiywM1Q46WvcGG5reWMXBSQMXOuUHNE1mvRymqxL0F6Y8dzjHvl
PQLzeP+7bo73jW2WOFaZpkKK2BALBGAs9rWHBbe8DvkbG/ykMsSzUSN4VFAB
6mlCvx1OO8ohKwU3l6HqSYTn7Or7zWITyowvy57LWFsaWMQDcg5+lfbAY5Q9
s6szh5rdmLxRq6UI8OMOUtAeKMmGimHoALRayk344UFpybaK/HmvLdf3prY9
nfQIC3KfB7KB1eyEa15HDYYLN0hOsOFQTHJ4lSOxV9BSQOATS8oRPgDXBwUQ
5vFN7z4J1OvfQJX7MThv2hN4/laGgna33Q1Ne9aybnrN4tAZ9PFTB96ShBNS
YSh3RYppcnQGR4plYtVZ/p6C+TkrmuNlTPVdSKRNFOYTQmorbdVmCOGCBxuD
07i1aE/KEtlIcl4fJ+1pfVumttGD6WMdgtGzBDt3cHQm+DVy0+i/2meIuhZ2
/L0b7cUCnfzpXulag0yRFTLDadMSqbPeqWnjqLFbX0ZI3F7Cr7GSyg9Nu8BQ
wAj/CNteD4gYzi+YzL+c/CWoSB4WWnaK/027ShVkvfe1isXb/mTtPlDdx/i9
2uVuiaeWhFK8UK9yFK3i4lLaYbg70Bf7TN1e7Wzc8Eb6p8gCj/kDeQpKcsEv
p3FUiDQpvLdShGN1JrZB58aspf9NGkIc+frgTTzNHzThcMem+ynNe/rBDFzO
yF0iPpJ1hZBGNEDicM1SURMKX3LExTN90O0TWm4K230YmpkCGGRsS4/eESCh
fIkfbNYM++q3nFtGm4FJb6OhFi3UoMALVW29LTcJb/ozAZyK6HZx5DQ10Si9
U3tX5eE/e7NuawHt/OyL6oqE3nTzd0OLdgAGzDAS0sreyVSMGz2EZEI7lg/u
LNLZWD3UCLGoIzEVN2RByDIXjjUsDj1aPKNguqBO6WflLo0PFRfPtZAt7JDj
TDQCMzqNMGp1YeBo11aytri580qsjYWQLqJ+/+lUVNcTFXIrfV0taM8CMIbC
WoxWLdWc/P8vrzGgGd7G8u7x9SGrHkLLXi5crunBnZDtS0JClpsb4ihEX6/c
a1K9DpJAQsT8Qx1DRrE9G/AqqaxRLjTTZ1Niiq52C3Be7DCA2bkPHSFiOq9K
qy2fhEYUbQleR+HfqVxwS2MyFaCCH6w6MONAkAhO4P9gF6aIqrpDDXGMseM7
sNgxkpp9qNe5e39exOlouTmnndoWAVJJCkLN2FdjxkZL/B7/qvSu87xvxUFq
g6BhUVyp2+OBKJzefrNopajWVTd3gQzNBsaatYAHnNMGLdKDnoJpL+j6OCXV
mgp+LQMH2lLE59MPy9llJDq4/IyqXokJ27DsCPu+pc3+rwS8KACivTr8iwGS
4aYSWzqTCa4cQ+2m6yfnZYVfYdecwyfCrId0uH10S+/8cPjWwaI/5SulVJQG
y6v4khfvR2pxcIZSIq32YIN9Tp57IMVz6njVfqLg1mcQiGll0Wb9U+sl9512
fjZZG1XTldV+v/ObxRB5lDuBwlwWs17mn/uFPQ16+PiCm8af1Lj7eMpVlWSI
wkvTot7o3Q99yrQaPA401eTx1WlSTlv1nJYuj1iuO/7lIgsh0UBgZLZJzqlx
N0I/GLVVUu3cRVKrHqj/sIB6uW+2dwoJ4OgRGhhV3QSiCn56hC6RwFy3BcPt
I5IiCdhhqnlDqHnL569E2RxXsf53A0bv00c+jCSYn9jMnKnhdzz738CXmdto
Or3f4QUgOk2DOAtRC+ePPfVTVfLPm6erYdXC6XfLYeQuRNjDttB0k+lJiZgz
c83jAYS6Y2ZLeXGAVnDLhrgEQWpfsscY338r47g+/BOWDrRJp4WuWppilu1l
ULYXdIfHhXcK3PtZlUNdhmnuN2nUP6DUkSLKmICy32nPts1xUz2axkGs0gMx
5G4TjRBHZaYWa0diE1x6sLRL9hGrZQEPI5wBXp7rJCLLdbkWTxwu1eR9e9IJ
w/jOhfKa0EKVmE4tD3+0vAtT/5QOl1a5FNPwkIs3lCgbQ3HqoqkIZvsRB1vD
ucYGI+4stZ5kSbc6kOw05aCsVy5XcagDtcsNvebeWsSsO2K8PoXSDDHhgzod
k/DTO5iVZ3yk8U07yWzCnGUdvJgxXXSGTRLqdsSNIBU9zcbSAeWREptvXPsE
Ivj3lxt3rJSGJG982UD0g2rY8I7OLUxofT+3qtVM4OJjwCs8w/Dxgo3Dbx5z
lgUR0lUXHScoAxklGzUHqiqr/ZqjqMeg+WPTg0mWRcWpHfrT2YVAlEQiHzah
R2VjsRU0Xr6vA+z5nYDbBQ2j6OVhwACuRCuyVbUW4dOx7H423NHfqj1Itgxi
M37GUWFQx7YcLG0KCr4W6MrpU959dlUpwqEq2Jv6Jq+PrT+bFrn7VOTVS/uu
5taFqOl2izGY1LRhaJgmowURbSbgBCHylslhYsf0AepwCbScVtuNevSbnh5T
omgNKfEQJ6jrLvFfnOJ+9/XJoFLov7VFfTN+uQXnIoMHBGVHbl2Eh/aIFYuZ
LmFVPKMkgygcM56p7be+slnrUjNIgWKuxZy95I8+N/+q+xJ9m802iytz3TqN
qwyz6JKu4eHdRvS0bCoSul15GqeK1l4TLEBq7Lsoo9XCzLuFFfCv3CGUmvpB
TMWQslipmOjUasuqgRVQdLa/F6SzJVxflmkszINs+2QwzGuMVTGXkISVQagW
lra94mhDXJncUOXs1/6wPP5nf5dts9t2vnRZU7PcE/HxB52r26O6vev5bzAo
E0AtpMzkZZ2WPR6cU0bFeWohmzH6kW24ljYczuH0tuFbrxxy04mzgGND3vCa
uWrod0v9Np0ChFUo3XirlbDEBmuH+20E/J9Cpk+UP7RcsIa//HjLEUJ7lwFJ
mXCjKSo++xIN2oJW4nRXUCMNRugZgJ0Oj4oIJKEY/Zc/svJfrA4FfQWl9qW/
tNd7LtiyKi9/KmjR6gq6VUKvOSSca9kcVmPmyNgjKZvPEW/XY2mXu2byLKXE
Uz+3AHT2sHzyXtWMfxidN1hGfI6e2/DF/rTKs+wvI7hA2BV3EpnMMAtE0b7y
IclV3RV+A/vVItrudwDI4YtpkcvP7Q3v3br6a6KrATUtie9L6i3kPSrtsa+q
ppveu25MXMMJpad2gpukE2otmDv0R+JInDQAxH0rvpgEBur3IeoFyp7q6QCn
Ga+YAKhzK85wmCTwjWpx3ilkEFmYE8FHpL1R+MhlOBH0dYYHCZ17G/Lgj6nj
6qgaU54Cy2SfRSaSh3MbCJOswIbCOTuBQOCUjL4Hkf2HBBkT1LDYUah5Rv+Z
x+P3w+2cOp+5wvHR9/I1sI23DQljMg3bgTpCf953zGXhkJHtas3Quhbu+V8v
DrSr6KGF5mP15/x42kyLqfnsH6Kiw/0hSKPp9/nwJshsVG8rDdsr6yapk7/s
zzr8CbJazBnCuNZIavWLxhx9aXBJrUH2uiN9VrZ0SWUOK+h6cUK19RwKNGrH
BAecPzDaRvfrGzRLgOetbB5uiMQH5A3YL0hkP3AsbeorAm9F7tvg9phwP1g0
fTGuHUJzzM2gtJYsFfQ5f0KJT3to2l3NKpy/aO8m5KfINt3UQQ38PY5rlCML
Y/gMV/zX/lRPI9YXN79w3BCUfN/z+cQ3N4rrPn3JcRfSWN8g2J4uUCNIpfUd
Ub09QAYm9GZ/jgVX5weCqoWabLcv6PXY6cL6RXmUNDMKcgudILEW3myzJiyK
Pf6PVbAMY3jI57m2Ybt7aPBV5qn6G4QgaaKlKkP4FzwowVB5EhDnq8BGmqoG
bj95orFaclUrX3avQFkfvrn9EEW5SBDmcnGgA/sh/y/ru5FMx0R7Xavy4qXD
/nd56VhgLa1i3Loxx9YfJ6etctf7u3EGRmpztzMPrboP2LEQz3pbwrUmMeBU
kvFcLRh89Ih11TsZvwTrei5XAmdE+ybsJn6m07+0TgNFOY19YRKksB6VB5F9
yd+2wvOhOZtnW4JgKybiKtJXbDyUj5Zd7Uya/xr77LXvML0quaFi6632fkKB
IAWtsAXO8SU6ktyz6wjDM3BBgsCG17y3l7vL4LLHlHi8GNu9A8igoMDszR4V
+sGmB5y3EwhRFOrbOWLo5CPJxRzd25zz7Mqjq7X2UYDrz8qdGlhkzXkAg3uZ
UJBs8bnxqus4efsot+x7bBEg4QFanrTvCxhwTwC/Mj9pPabRJ0ZGasIPlCPa
vIlOg+RG481VHSov8mxyP4u3GRnAz4a8toZzQLu8lqD/cVYJVKZMv8xK5FJ5
5LlpRLBzp/gk4OFx61hCONc+d0NBIYqUUrbcnWFwQwkf57fALgQuG+iZC2HK
SN8iIvgD4FAZCAVP7KPyzqyy6Ik7UllFmnk99ejB7pwRVsmZ3MDOzRdbS4qp
hIXMUMfl77bWzDvpOmudAtNSPQzJ3Sz7nRdS3GSJqgqdfHpnVUsLlw0NfDmG
yGI++4F585adzT4AOLCs9IeYj/tfQzURFgG8NhoIu7B3JPAq3mh0h5YeOUZm
JLfU+lIEsYLsuH8ApSOaoptGDohsAKIzgtH/wiJXGfua4m29mWMambKTu8tK
zKZKv/hEC3ORW62qxom4Ubw8FKO/1l/JDjds+DHv9DM8Fj5ndyq71uqEAKCQ
Y+vujNKhntVUYk/KPE6+xupDVhkL1EOL/xd2XPtdYukOJXovEdttJR8y8g+F
TJd4jgvDgZig7r1ORXXu+Le5QgpaFR2N6s8e+bnzL5kCxL3KpV/BzQ8rHELV
B6D8qo1TZ4nhqNwt9dJSGHkT88T+mx0lZEaHtGO+zmzY1qXt3BWRXfMiYGsy
AZ0jASJZWeQqE/2LYYHNHwrCqFPwlJAJFFCaP1at2FiqM5rTi9WTs1zv+jFk
zGrrLopMSJunfdRallB3Ao6Wq9eROkG1n4sJwtdt8+Y9Lrwqh9SRqwP+kAD/
GhLdJaIri4GlWAEcxKqclBm+MC3NIOU40aNKTr/P0+gYwTFLlpDnVCfsOsjr
jQvj0I9Lfa+pXVxgo0k2eQNHkfXkSbIa0wP1XTAe95MyRubEPcHQgGwRMTqv
OS/ihkPnP01uFvVQhM4o7FF1CkNy3RIH2MHcNfhAHTuvjB2qUqotCwP6Td8+
2vyXUjC5wXg4xbIG9GSWTf2Or3n6rLlIlaaLJw0nANyR5md3FTGsU0I8NHzf
+JAOPh6ZJMuPBCgC4wr1A3FH/yyFxDnnPOb/l5Ebywboms/v8HrxVK9hquzL
vhU0GA3/BHHDweYnA9vx5LU11Hm9DaRVzLfDp4F1/W0Mlz8k/mTax0MBQK0Z
ftbP5A5yE5Zi4zSgS/Isu8Axn/M3PSB0TfRkWbQoKsMVFc2uy+70YylEpOR8
WmkM95AujDM4adtA/AwnqM+pNzqXUJ7Mvlqdi4yMSQhtRxeVYSAoN+Hnvx2v
HU24eQf0WczJN7MZ4T+rJ0T1zNrqth1CXy8akxR5wW0j5pmR1H1ZsiVeXibC
q62i8KF3VqGIr2BwnfRPTWgBlYviYsnhCF4nLypgiBU8aPiczfbRm+aCbI7x
osVtKvR/X1ZvFlepCBotyERXTcTpBsGCgqUcqoCPqQdhyPgDm/R/99d09pMl
N6WClF7pFag0AhXN8jiB4N4t4eePdD6ljFFJ90HAaXnpXMirQSn0zVQTTJfH
POyY/tdnumSRRkHPb66MkpDhxy2/U3Vaj+fektLzH5ek9QgluTFX6CsHxYMF
r9xehj9uFKtQq99LsTzU+B7inT7r+fr6E2SCbZ1UYaM7FcRLK8NJculzSoZR
DtvWV6ixqHMaNxDtv9Tv0wSarAqtw+862gUuYQzKwOL7lnxCYis1ZeJP3Nfc
fCgUva9pxhTzy8NupbnuhtOyPRsY5SkP22Qhyek79OBiuEUNdo1ekHJZ2uE1
wmu2vyx2g3Jxim6qAwLI1Da4Q8DGkoNK4LTR7fDpyOBdlNMCHFUkxKpTzdEZ
/7f1ed1AbfHpekth30mZX1Aebi9oNzoFlHISdwErdZUEh9drAg5/LtoPuEW1
u2m15Jqua8bIF+r7J/wc5292YT5xFGGqmYt1ih6VsCjnpVM+2U2Y4Zihqhmn
d4uWeUE/1hV3K07JOtHYhMj28S0xVKkvbZftO7UTcatDLR3VXi62dtybx7I5
vaQGYJLVUt+gEHK6J+g5KE97U1ng3wTeIumGmj4XEsdlsSwn1kAuo60jxgYb
91nffOhj4TnJ2GXBh39IXUvfP7KEAU5yMpetNSqcg8ZA2yCuBojqX2ONJtyX
MhXkvBZDZDoBoGgLJjRD8whbAXih9lfL06tcdpe0sPRPNiGxVtrhOcszoLe2
CPWthDszkZoartP18Mz16WVaC5v95SfNH68s9ZbHSk+R/ao2KmoAyq1A7eIG
FrPBVbQB5G7sGXu+VRb9xJoskv25tQb17VDpAs+0fHSwaT9MmmXcJ4ueXqKM
qXwf3YvDZUx0zlB8GXWXqt1DbfwR5qXF6ZDabIklwLS7VRb/MVKCwDbtDFsj
IZWg8P+1LZcjPcqcxUPNP5avTU7xVKnQfwnRvTweFosi010k8eJEWYxshZDy
RnYXfxcINJj3cxhs2NjpSlo/jmCb32FMqzmVAgxVFr+M9P4/JeLSuaa2Ztzb
xo3mvL4QvNKeIYIkBolZigJr+GyL3zajfWCw2Dku17PZVclXpkA7wA9+m0D9
ZiJFadD4hlER2kYb0+Eqc1+u1yj+3xowh7BW/QjEfEVRhqDNxFk3Lu5uNoia
YEayuXcpHk+HkhZkBenaF0JclpvJTfyIgRGOOxIsLQO5kwYhjGyt2FkLbocf
2WhEZlJQWTLmxaFm4+yaJPD2R56axPZxyDvZcl+JblF/CPPmr5EloPScZheJ
b19Lb+jws6JisXLTLT0wTp7zI2pS5MCn4qSeG8k3ECN2HuTTzjxpLgvtgTry
gwDKbafgA9Dcr50m/NfcOYEI1NbetejpvutGo+ctRay7R8yXQgenF9+i7wOk
CaXhbs1dGqEUJz3T9QxD45AUEfw6ogQtJHPIw67+qMcwxS23jI4U/E6b5+Wp
BwlNNAaCt/zQ1Zfa9WQzcukwXSjzCszh2wUglR8i/C1nDbPKkBa8mH1kspoa
fkLYbqZoEvPyizYUriitZOVpYMkxg+xIc8/qsAXcYsMFGZiJpNUcrO2f0lZD
lmFO0trfJbo/cjzaBX1Kbo7VQu6JQiEHtyePPSoWWDYeQK8BlMofRE1hnbsb
Vo7ViAQ6THskN45zq+1QSFFH65INowAFQcqGRmCgOBKL34TZP+K1SExJm0f+
g8/SWpstI06Pth9dwAauuJ5Pk4PJnkcM1uL4ZfQmP1BMarRKVtvcfSJvWJTl
+OCY+hfYsHX5OSmvRYHgkjgfnFQ9U+ttTfRXtmqparQG0iERPDU09qyhxT5g
UssnZqjY6F35EouYSEuLiX3e/RxtyAMjI8Q78hn+zZVnTYfRvfzuM2iJDgVh
Ok7uJ+iFEZkLSHTCGKOZJx4Up3g/ptZfEjmXymGf4aQFiKCl+3JBwlQrKx6z
Nhy7A3DmYZMQe+HuQ4NxXw8GdQ4L9CVqy7ql84dm5s3ndhOfKi7+z2PkWtrx
RN9Q8KuzIY5RohJGG/Q0Evq8qRzE6s5mh6QgAT3QPRxz4vWR8Po07IVnAJlI
AhsmMmzsbcLj4AzM9zBEhU2NUrkx3li4QfrKw2McAWv4HnpCFV4gCD3zjzUX
S7mdTWrxQ5gKxGBdPXmi/oF0rP3Hl+UZ0uO9MpC06j8+EzySfrT8FxbA/8wZ
xdbrIDkzGjKQRdGac9Z+DbNvANNU5ER67/lrbHU/sORdpOA9CLVlK9otRkn8
QsI8SGO8DbAKJzxtfpiPI1kk4C97c/gEFUgc5seKCHo9ZiVPW4Jix2h1QWjI
/wJ715pAMQRDP0um+N1xujUB25yvrMj+E0PjR1r2PsvoU1b3U172cSwY9EE8
8B4TsW+ULmpnGAMWZILqBV7IF+ZMuRWgnmYcyurV8v6fSHEFBB7MunsV8AsJ
pgJ2oMUUKXLQVM+wrnal5z/ChY5sG7Zo8/HvOv14Qj5fLdgNNPmmC0u4FVls
R7BwgE5QBffTEzbx6aOWld19YHa8p16NHNscCMu39rgAeQNPEOMeBjagdGaK
tr0mnvIUfzT8hEpV8Cses+iHNVNw0rt5D3ak3rh49RhGFX1kGoS6iweuBIrt
LCxVm5zsaAgZz0r3DMhY1pq5ma9TWDDnxHiLYejePYhGhbAv4+9tj/ydkxb7
8bwwf99MEcxpMSNqrnE57ZWcJ5GWL6RxVRda+bu4gYx1rzJMaC2i7LyG3tft
3NaWbSbDpI1pVlJgu8Ng4EhUXAWFVfpxTFkul4hyIDIk54mGVd12D3N9UEEy
7g0IGe9wBSnXwjs6RDaONSm9WfDnq+0yODF0YIIx8/gOhhyiyoaRX7WzI2CG
DJ8cnlhqRHMiP5TFO/qZKPLQb9Bj2jeNYB8mfKR9pK6Mlk3+9BGYBVe+e6Mp
m15TFPrTrRwZBRB9AMhxPP8278Px2pdmvKnIX28osJpGOBvjJ8gvPokDfdg4
abfSWNyQnH10JSyEAmKECXDyYi2jSeJk2nCuzZUKQBd/Ju2lmZI74hJ1byX8
h8fu+gwUSKYgPtJ9L6UAFPCTxZdmdQGmW17U4LEHAgfT8rxphXOevZqNeEaL
YWpK95Us1q+G3lsNwI4uHsKrNhLq8RyDNdA98+lZZ6Zn7HCfoKJajmot3sMU
IRpyBp2S1FsBtrq2QJEqLr5g42c7MQu+dk/gcvGxmkt94zkrJO9JmjaBXWVV
SrlTXlHipxxnngGUFLchNAHZr01cePMVZU2CjGyTc+3JRSJvzLXxDMbQ2YtW
pFa1nvVwqTYZticvKDn30ZJ955ETIfYsjBc3jvtr37TFFvp1l8rzH/5iHkrW
Hi/tGE+W1z5IIc8oiyPqzqQXyQZ7bvTXUhlnzzrVKRsfeRiihmFGegU8yMgI
rOGVjajEl4TJjBnA09OHcvPdlnXLMNnwSC8UpfjSYDkl556BSg5PUulRb32L
U4zOKkD0lskxO4CwLAUrS+ti+3db4GW5mPzZa534zzf5HWoLjaQUMBeGCxZQ
PZwyDApc1sYPGOyK4/epyXuFMWs+Vqtn0ZZnOpZElwN+TwUP++nqUBSnWguR
MECamWdy1Xg1syiaBUwIrurdyHjjlw4mHRzi1ic7rfLXfjcFlPAeD7kr7RLA
2WrepyiSAEIeHoSffK3xzrXTJrL97llEsqlcpEt5Rv6VL92dOWjTo1RXzbA5
YCGx4FV0dQKlOGstldifrdWfaVlqjDIldZgwio4iyPfaVpd8Hy/DpzyS91if
+oT3H57fErUx16vSBhoTG/wls1AVzks5Be0QJzNI2ScjhFla95lMNL/h3ejA
jyPz69UVrcKdDIhM+LTTtvaCnpHfzTt9zBzP0H+AF1AzeAxxs/XBknPv0luX
9zVrsuZHovw+HatVlVl118wDrzsa2Y+WAIjTmlqH6N9PoyqYDa2kcKahhped
c6hJckGEtNG+WgjESFRcWjD6IOfPBM0wXapxqdRgi24hD0r1Z0z3nWA8KxjH
CufG621Wb25UPuPSicuNUHmgCFJdT95xMZw5WPspEzLd8u7oHoWQmfKzgZjf
gmPTl051sEjmD2WuNpwlYZaTeZ8PAHM4pOwipGt5st3UcCutTjt136qeQ2BW
aMnzbKry5PLRG9UKdnCKQ2CsRZfN8wG4j1AnXMpfZUadu4AyaTevaOPlrhxT
iMBpTYhRthq8w0mdNdnfOTc6ZZVqnmpET2YWtBWmVe00FgqZxpu650jwjLur
rzA5lh4B+3Wnj7JNK9gQvV7Hdr/tAcfw7G6v917IGH2CY7NIbyRCRhknRpCJ
hQ0p2cIngqow0dxZBhI0oCV3FeBbybWeORBfFU5T8SbIc1xvntyX29puh/ZZ
3kp1V3GoweYxhhGr5x8dJbFWxuPynkWmKpHtNqd9OVz1ehF9X6opZzQ3y81b
x6bU0Qs72rgGNieQH6U6ZajvOKQIvLHCBjBlLx4JZQVhjYEq7fw+9xFS3UTr
wSEJzCCucCDVzEGwrgoWBxcrdLoD8wJEHeMBUaamyzP7AGgCq3hwxpgL/Ka3
7/ui/m8IbPUTjL4BjZrsyRRZjsN2pYjyqsN4m7tYlimIbWibH9cDmlCC0JhA
lvys1rlJx4F7dapYSds5YGEd/SOh2WhUTTIGfhtJRA8OpAsaGJSNxYJ6HnbM
HwX7ZDmjDCZKvty/alaVGYvLx6m/KWmlFwg2RjslZpxvIYqWs2i9sY5R0BZ1
Ff+szzH8BqoknENBwNy6SdDyk2d5laGnn6yDU23KhGr+361W5sR7rcgu0OqF
fi/S3WsXL7rGJetOeQjfYQnSr5iVBW7A9xYtwFQpEyHTTAY7OqOTEbUmG1ti
T2FIGjK78C1TzQZn6Aa15z0qjWWYmTaFGAU6A5wk/QUPnr0w1ykPJOvpS4J2
PqL35BOReIHvrKYNkSmcGDwfCsHdGsxhhjQn3cMVk7tbzaqNqOJeiA+pifzf
FgHaEXT4zBxqEVBDuASsLPh5FFnbIVCiVCf2qrAIitQxJ3VC+jf7PSZHixap
Kq2ovbG0n+3uZo7fJ9jnjvDFLSm0wxqOmGD26nGXxce5vbJCD9sc34FPKnHn
2CK4/AKpWUaj20GOnPlJsNd1+Knqkgj6ScaArqvVLEHFGazW2HdG39LEu0m2
CqtC2KPWuCcuJk/dEpT7ehN75Tja4711vUCdMjNDHDx1vpC8nN00MtlcQsoY
r2hYC17QPAJVxzRi8lzOiXsXO68NyxQr7qh4Y0SYo5PV5xCgm21T/+ZABuF/
xl1Oc1pr3yTNe69IAtGTHbbWyjUkVS79Zl6OSbi/K0evGB1rEWFN8o0Sfni/
cd5G+1mbERSrFIwH/JFt8PaWlxwBymepRniHyf0yBInrz9qDLIp8W5iOb1Rn
qYJHfE15Gx1Ph813johiaCPeWerIlPrLHXnSppD/uAUenHMz41y5Zup4sQ1W
krReC+Ax/VWOyzmfeOJ8fme+o+BwFq/RDU5GveWzG3CyFdP3bJPgmxtkauTb
Jo8jN1UBHsrRbe69uDYmyPBsqEg5vvf6CKvP6skucal0z4fRrLHqXOB21q8i
qZs0ej1zu839LAuODpauEaKUhOKFPuces1wr9vcnnAo1QyxV66IjRufK0prX
ortpB1iIHcA8WRXM51OTM1NW9lz07knN/m4TnSIVCWuajFyMM+THAJVT0jnw
+WTW6XdBa4L8Fk3iLRi8rB6b6NIu0fHmEs/D/hB/xoaLAFlX7q/kVU6FVwMl
Z9vMaWV4P7QMj5bXLQxIej4yW4+1KRjmRt+383quyk8iz8uhrzYRyGWooxLJ
7WTNP7jJTQnf7mBGzfYFbmvZzzPqxSs+sTv5in52/QLNFnuTL+O/ZghIcvEu
mnX9YP/ktk3fwdtOURIQTo3ZAxivM3GDcFn3yTt4Vxlp/1W5DCAf8rSYehg3
iuHtVMjApz0zUNAumFv460/tTcD4HQjQd9A5DjjjfxMK/g6pDtr8jrvz4sx/
GWY9Ksmw822dLc5B9RZwTWcqwUj3AR5kaDlW8Q1PBi0buhTnv4kemlAiaOzr
O6smohLsDJPCAeQCEzE0/hC2F+IdaltveDvBn3VQZRRv1rnLHQiN+9iKGqDx
tzmEsE6qmIeDu4GE2k/5GDHjP67N+cR9Nd7fzR+/4m/EvoxWJYwR37oiA6ik
iScx/55enXRlPw4pyIMWqt12mIuldiyQzMkv0jeV0di5yYxEocJxFZhhDQ3n
6WLrpcZ66R65SjEUJOxkqBfotH6wqSkenyDN6ArVRD6AacSimg/ujNfOlDop
Sj4mqlwt+5AzLlt/VvpMVrDD2KpRhKGobr8ESpzezNNuckE4M5PuRcgT1AsV
P0f+G0hzsjstafl8MTpWjQT6eUHdn8gToApTvUOQV2/niIshfEMtPRjCKnkZ
0fvvkUVulOaE1S9QAjFeUzPz9pLSJ2Oz4vpA+nROPJObKijXX5N5GnDdy2T+
no6/l5skeaZ48bHhDx8Q5SI2pJ+QYb7Hms+5DdC++VshkaGIR8T30P5UoVUL
CQm3EaMowaayLpIYRoWSPqWWf2F6jC/eSqrgljOroQq48vuY3/t0L/Q1GTG6
cvM66nC5YCJHP3SrbiPSHDi2fnAhD587k9tfoRQhlc+F8s8FSZU/EArUafoW
PGobMNiHwa6lvuSW3k07kw2Rlm+wEqMFxGhVzb3uiH1ocyI20kGNqs3Shf3T
zXFm++Cw3EvKsYr5WudCJlNa+reCsu1Q1ovFFaHTk0TWDc5AuaHLbKalHh4F
jqAkWcjPFwWyq4+IIWuKdV8mKA9uEIBzdiOo2oUQvBGnX7nKoGPP+xRShPMr
2e9y48J09YpZMpf1r7DK/wZ11FVB0TWrUqAKneYD887dPLvhfSvwLERRQ5Br
sr37p02LiQfrxtQbaLFUzTNOFIagpStFhgRekzSKrXja46d6muZYtGWVwatE
0fngIXz6YOuLDbxUE1S5V/04s95zEkmQgrL+av1lXkMestUyPzDJfRlw22/R
rAmiwpPVHtXrNiA33f2qCgB1lYo9iGEvVMaZs1Doym5zrY5K6j01PY48useQ
M2SDU8LmKKf0/62eWy6BGSQqEFSR68HL080X5sgPEobN/wIF2dFgHpsFiJrk
IA+TxLjeYXO/nlXDNJpySEJHn1c0BXm2Jo2yOpcVY1wny6+dx9NchEayH+jS
DsldNyU0bFvfTQ10MRDL6s8eCZv+v74e70UoRAqBIVmB80mvZDwgQtzYtBW0
11CeqIjiCdYqDxayajSYubgyMqcKEhcbV9tNVd4mBnJZaobg+V5TC/cKMSGp
UnYl8gfv+GHNCZ27lhIBQI1NW5rhTfKiqOWeMbVoRtTwECet7HMbtMSiSMm0
fB9iqSTTv+yFumsLxwoUaAu/qSyS0/r4+ZOmrAtBanLInUP42EXC/hoHqcZo
R7Gb9EyjFBnPyvr2B2l+GQNpibml1MYUplEBAvyCjm0fZ6ixOOTIApmFqmnT
Atiubh57M6q8rEprWtHo1i5wtZSg5oWiJxIuYU5noT09D/SAl0ioFIqVNlM2
2LduIWEKCyvjqvQfD+ikHA4w5lR5kzqTiP/mvjXzhvcoQIeyb9oXAZnnnH85
ZE5xVjv2bSy1e2y4c5YdK2ti1sS7/1+AtSCZg6fce3m/Isv/QbKmgcgm6UF6
865wyJugCEb9Z0NNHhHsCuP0gsvKOWfit6CxvMGUT4Z+KvbOmbUXZksuLr6h
GQ18wlev+H2JonPFlV56vX5gKBZZ03YFMamRq7q9jRlJD/1UCRtCtHbiG6fT
33F0u4cz+6mmjZLQS7gKwRSmbwevyV+CSSLu9KQSgRVYWxAAZGS4Uauf5foL
Dq91qMtejiUrZPsg+JoiiyqETNBPc7OGIdoq2kH7eervq2+YLYhXX1SbqLvc
DRzbi4c4Gymsmlia26sG8RbEzNkkgWXg6M9WHcOizBE4pU5viwFf4srYc+pp
s2li3xSQC+YnTuZeuKAvNNNYiZJ4uxuLrSqhH55yDlKHL/wGLHwM7BeuvIgk
a7yTA3hkgDX2m2W2ZV5iXJkdXtpRjb8fGldv6uiSK+xiTVBBHly9VNM8y94q
e9PX4XLY0vVvVR05zzOePmeXaScvf2vgngG7iAU7RbGXHDNv5ocmQHirryY9
g9sQ8PwhzWjuE7oLXSMDCKx8hgfLbZZqnrBp7hVMyg0dLVxOLjJT8oXp78GF
ClD/IGn6OGLYuSV06tKB+iq7Jl7Pk2wbm72b7qEYqmgNQ51PZTQZA19Qghru
sPTUmw5Jl0/OcAtk2BUgYE5bge6UP2kfF75avrVW+Ok5ht9EkgykPhcA3Mbe
265UttfLEsovqlY/Lw3jkjnb8w+hsYQSZOscG0KjacEQCJEF6osLGTSyrSme
U8u0D53yTT1bmQVCjPy9nB5ph7TMfXOatsB5UZHKV3glw9e+toYaU6PyjMe5
kTFr9OiWj0ClgOtBvqXirCvailgfpGXRBDJEolTvrlC+3NxqvzRTeXjguhQy
VTMHrs2hV5P7KrcvvDR265yOx4uKfEEtWq87Gy7iiFqkp5YL81uKPRE/+Czl
2gfPK3Px2ejjf2iHerxMX2UWvVFD3pb1RkVI+Td3oXCMY+G+gzJLZFOlXzEb
g+bfG1EWjwZ5e0tygiU6qgBJ/tVQ9cg/7X9z3iIPcZUDayPsCHSmhaE0BbCy
D/M7y0PoIreKQ976OrxHrvZSaWLkFOj6omL0266UIwl23+xZIY7YeKJTpF2D
vJE3pYruaA1+o1lCL36xJqYa0/IB2huxb4AEewmS7X82JV91xlrSSAur9JI+
GVp8Ee+8aP356S0PMazWOP7dCtDWRMtnqsE1V8HNvWdwH3L01e1LzJ7dHy4Q
cCL2TbjxClykd451u+3pkYBGVZ0llV1zMeJGPGaLrhbuhYJejLY5tI+I9VO3
/y2R16m6CbqodDoqTSsw5hz4fusdrZOstLPFs3yVgNEwb3ABy3LgM8iF5PA0
XGzNuMLIFrmJGpFfprJIs6mEUrOQcizpk+kwub56bW10+dhZQZu/G9v62L/U
LrW/nogiJjowxG+9XBl7hvoK1TnTnKzcyO4c8SvzPZtCVjQiXv0D8uXpT1C5
6e/ZHfGQPucU6QJFGOqdzK74qGgGn+d1lMnb5UlajZK0E/Fimu06lMLGl8f5
D1eaT2h3hvBAhzacNB4zC2ZCjxUi+1cz+J+oZAbNJu8825SCkJtVWPJzVGUm
m5HPTc6bpOKwo90cfPBnfBcV2+TU87oCJ9GvKpgO4SsSZv4y68d63aUi5XTG
qCeb3KRGlmUu8thA8pWbVYU5QpWQ0wU31FCgpBBIC0zWROU+TR1eaKVr3o1g
szmlfgBD428kKax0bunKEmLww1Yge4a7CbXSuAUNpDuQqhg8Ma52cAflsPHA
aIdQ5rT50EOmeuC/8hQqa5OL8bzkp5pHrgKj2Kt7FtvgPaGceSZhYa0thXAC
7I3YdrdsJ/UH1G9icxjVdybxnrYuaJpGh9J2G/Xx08nLlW/JSNNQ+kr/ND9K
FImTCf27h+hSRNqGPdMZ28KJDSRBMkxl/qqteg7zyUCbNPVvGaiXC/SJV6k+
4XPPa/xAYGr1qAif26v2Mvxz/9YT0p7qAauNm0iz7CsIlcaL//KJeKDBU0ip
jnoeSGnqEmluxAuVhTJEzgbhRg82peGljEW66IWVqV6nRdYwrdQC2LstnrNZ
0eIY5OssCZx1w0vvI5tgPgd0kETfTnyAGZL9f/a4ZbRK2JVk46/ogJqpytab
2Sb7gF/URvgAX5WR7hYH8cVeQSEkfXc/YTMBjuyaEtfk/W2xgkTQhedUXOYd
I+5HpyJfgvRAxTUbtTm0pWZuJ8BCCt1bOPmTMcmgwZ1qrDngGjwGu5AZNvXz
BOnfyo112Pz26ppb6NMoc2NjlEjRdFrws/wrRdOTjSRIuo3ctJalRUhyiJYA
1jDK5bvTdNs3pjDtJeyQi+3m+H4DlxupaoyJOXJjiWEUVFpzdQkfFkKBlqJ3
59gmqusXj7Rxn+PbkBlzPWE8+wy1euWn091ukjgZ2glq2d3i6Rk0dbV3fpFu
0j1zrofMT6ulmW1Zw0yV/cR27BaMMDgn1mesd+Wc5WQ8t1tsUBlS/hQTzcBu
ridwJGY1WSH/ChP02nfWS9gLEh/uLj07Gt4BH9qyqatQ8HijA0pgJyTRKIuS
KVd/27AJ7TGMU1FzXMRIL6l8MgFtGMPLPTZIdd5xsl1fTmFd9y4Tz5nDrVd+
l//Zaz1Nf+jtYVA1tjrTExJdp3pdqHRrdbvZFp5HAWPqarXDVUmCqsMwSluE
7o+52rlYjrv0IAQYxvkTq3jH1QMXyBlIUV7EQuAf3WFVEpyWPenL4hlI1WBV
QL+gV3t0+QhrbeHUa62OUCGgdsgpdhIlVyN09snHKrjeS8UAgEB63tc0uvI5
Vv4t3cX7GokvibUhQTUuOW7qUIJN0SmBV79q70oJXvteawIHnpXT4Xcm+Kfe
h14GwLwLjDSyHlQeqvSWsnYi3AEMnD0Qy3sNU6W6YLaoJDPlWqyvo4d+Olp9
E41oONYF/d4mGHNCW7zToA/oHVIEICggGIvOk5CmsCC4Qo0IVNLegKx6O+aI
lPrbt5wK+BfOGiTyHbQ264Vrv/cT5GUIjGEdBiu4h5ULd6EBUfwYwmcmFj6f
qwz6xL6tvHHryCRZ8MtE1xoBiMrioiFaJr1CnNrJUVEwJ57RkF3YczXcfnYd
8riggLeOrZWDUBqB/xndCs0Zfl2Yi7FLR0anMMVYrBk6fDZCAqsHBVAROmDj
dYWnsihBdyGm7+nfGmdE8xxdfNXVyOo+//Tud+XUMKdwKtvLYs6Cv+71i5GQ
ZXLxZbVNhEJ86M+gEEXMaMuc3lL8zRWuEt/WTN1rn+Q+pqzTu+Ul3AGSEB3m
+wvmsB976Bz1JurqOWVLEZzVZ+tMGgkJc0RxT971b3bop5xGk/cKvgmHpAFN
RmuDdp/3DGWSFfbdsp1N5D8N92BJV3yXD/9ZW0iAjowzjwMsHLYSL6mM3orI
+sp0A08twmOGxu3n0SnizjU9hZchowDz155WD9S31e14ogCCDnIHbDFX7PnW
wtvea2Kgl7kDZnMxmKTipYFq/x1Fj7VOij4SJjt/2iwfmb9cbm6+rJT6iqrw
XV97TsXaRYfviy772Quc7DlvL0Dw4lIYV+PGVRCoRG0ZmtYlxeaB9Oa9tbIl
2IZicg1sWdV+Eh5afn7e+gt6Q6edaUAlmVjzQVUjBZb3jwpVaSIxC1IxwVhb
0gNm3A5LGyVj9cVEDgRqIulvbXRP9noH/02KlIho2ngmYtDqaA4xgsCKrWfG
5y/8ZQUZpXrJ/+/HAO5N2reZtdVh+SvQESLpRmBT9M4yNee/KQmW1qrDaLpm
jqWXQkJ9uCJifCbHkYQTO5D3bKnWijviVt1OLjWdN92/oADgJIBsP4Bisp4j
lyf+XjY8ILr1++lJtV95hU0TN76ENUj+xMEP+FfiJ/652pg6IjwPXK2XK6n+
F43Om+Qs8ypyHr01lvw5AAZ2HyI3A8+/cYSud69YRGwwKPXpY5AzH/NIZxtb
UewOpx3lURqy+koffl/Si/FJbgfc6HysEI2ZG7EMz8Ux8g/nXf3w8Qau2oow
4iz3+d/MCZBd0DUUujUkksjA538FzZqDg/NeFMpR53zD0kngadOwuWlxtBnW
OS64wOQWlyE7Xcgy2V1PLDHyaxOQuSpx0VdZ0yiA/OdTSjAB2Fy91em59oBW
5IKYekYOmY7cvrI8X64AN7f2P+h+x7kf0hWnxwNoz33Pr9ZW739FO93tt04d
SOB6a/sITV4hpO95o4dSOqi2MGWCk+Qsj5dCPxJZL6d3AT8hsMmu7WmmYcLB
5AuaNIeCqKuOxYyhr/zibFVnq948C98LCdnh8nhPK+eCjaV/3opsMIrBnaAv
rpkqbMkzYqxDzFYL6D7uYBA/K1H4CnuZYNMzqGecHXecrXSOW+G6InqIL7Lm
F9GPYwFIcTGKpAFMeQo/hBrXno1JsfgRheQN/aXXPbEX2DXiulSqke3LY8f4
Z/2TuDE1hMEwKNQE13wzuRYFpn6VltRnor9wvMdbP2+9DO1u/w9y2xjbA4Xa
F1GXDWCbAVt3S7D/h8zySLdzIyI7OLFJ3NitI45QyWWCHnsvUYvMSaU/o9wB
R5pv4XnCHd8fCeF2ekLV/3yvaS80sgow+OO0ugkvZCrTwZkm3jTW2t6o9bdC
OCndVEQk3dnQH4pInZORd5Wlmy4AnbINMVV/qbBS4JaXS+7B72zECP3unsZs
l0PlBGs0XMZ8LN+YyVXYYaz9AMnoFIOKcOs2AoQ+KISlkwIXJnsSUHv1iSPJ
nas3cOcqyN2uktXza1NDTcJF91hBUDfQV06kuScPsgNQnH5pBdVDncdExDDo
i4Z1YVKttL+QWOmXRiv1mBhE93LwJZB5IuKcUparon2t2RPq+mTaZZ8hvSUg
kPq2R076oViHXh2qpza0PnwecAoW0b7z11S2qsBEmD7/1eszlNCg7lmr1+ff
1RmUDZOV9MdSBfu9PIOGkKHlrftboXobXjmMjMjGGd0m/AEOTCZHEsueGV6c
cxpjI+aBxcexRYvGF+UikBGG2NOm+mS/ooFjuU/2hbemrXUgpZ0+sHbIP8yK
cQkZnd6mrdzDoqgr75X/W8Hv1jSbfP4M4XqvrHdcMUuJZ8z47H8rcKfSe5dq
gqYd+L2rXm5CSFoYEnBq4Id3j7k8ujJTHWJcPxvTCxRuVxOnWDfEA8d514eV
sUBDdJTImzEpN06BA0BshwZsgEXd9vcGzPkWofEJCQ0UTTdLoN7OkuQBjdTP
8Y9k9rZcS3Q0VyQKKDR8VgAfxA87v7L6Wvby/n72RnlFDULvwpifbEcIGW5a
0+xdLme9GI3PJ/UUxtcU4Z/dLufoNBZ0Q9IgruDcDpsC1dytXICnHCh24iuF
hp0fyH9tkKBWNbiURrtWgqEn0OUlXNuZhbkeXBLoD4gy306GkfyJgeLgI3WY
FQ2AOXHZxZbgFZ4PCDQGhpH2855kbfYaBp/vLbrRxlVRPt6n+aeILCQSKozT
YIcyeEBGIkqG2pA3ks4gfUPSIe4f0kItaRZfzR/10FofA0SM7Qd9sPjTOw+2
As1f+9/SFLkjvTF7zBK6zAZfefJpFDch7tRBzfDQbUUqtjDNOAxV4ZIX81qP
M5V1wAmRQ+qej/ub4//s6FMDXDVJcIPrXfwHbLsfuZWh5L1N9cmEKIjh8Ytv
Mdc7cU3gIyRv8z1vU7TGr5J9Ty9Wc/k7i59Mf0m5Ceh0KvWYF764vdrqI9Qo
PiBV0PjZ909qpqkiBY18tQxEr0e4NPWQmuQbpJgZhA+X7qL3eshfWOxWO4cq
9+qEY3Ahr+glbCq2uo3xUrwISqw8ouzbRT9PQosMGB774SZQ1mlxy7HcoXFh
3JK9JA5QTcu7PGAOc4vq4cdpVKdIIf/Ze4gyJlgaQNvhafWDPjUTmH0eZ+FK
UlpkfNRU1gLXmJ5ffaO0JFpvKyEM8JlcyEuAVnM5J0J+9OdHvQS5fjUd66GL
Yshj2Ogrk2E6njXsuSFdkJoWUaiJ6LlcMWxaGLAP7pNvSXjs0X+lS1th58bG
Dee8JMKSw+wd4AAMe2QXOraOJFGy4WdrcpAbdZo2cIBBplU57gEZWntAw/OQ
ozrr874k3tjSX38618cZKMIZk8wdVsJwYtu/rtAvaQR9nuaCMFp61pHHizz0
d1mYle6EJyKybtY96P6ythZZHSXAFoIUxao3OiVHo/DVPkolXStjcv6rxmM2
ofgUxotTvJPnBB79lSLrm4fIObtcMa6+lABPnI73anMxAoPldouHgeGie6Zh
H20a5Ew6W1poZ//H4vRAUPxll6tl1idu99QWIyZdbqx6WjvrKRWru3JHlQr6
Qw3P5XCwbknnjPkFHq4qrBMf1xs4IS08Q4p5pQ/QIlv9JKWNYhsNen0dNNEr
zKSYfApvyYiKWrVlMneYxROeBYQ0wsHMvlqkQi/Hc7gWTV01PblG5okrtQzt
WshyhOlfZVIS3krv05bTzOX4qsit99VL7fk0si+t7KRbhJO8VgmoRC3Pyw2p
MpLq/zDI2xBnBVQbIjHjqxqNFWisIFNrgJxHRu9rrS9XTAvgr/jzhD1MwX/f
eRKTeqh9EQKrr3TNmV4Ry0Lld+rZqP66v2BuuSU+wL1oG/OVyaN3676Zid7e
YCkryAsjvp/lc6iilZUfqRhdcig9NyuoFB7aepCohzcE2lL7GP/HxwDSy7G8
neJ7SrC/qcG7KVpN7wM1amoajJ+cWEVmlhoAvpkCsVFkfE5+akoS92jjunmO
RY3zlrk9myBd5nI8Z8ERVyw/27K2CV8r6jPK9fNxK8AVImwxFUQQcXqBQ6e3
9OcjsXH38UECER5YbXSVWtTmYBJN7q7OI/FpUPTy+gB7RPexA/f8rxuEEiEn
P7EMAuCp1syfpXSICysPUJ9JuCc/fE0/8TdMDrNJuBIhZLDcW8we3VYR8rLi
nZz2XzIDRuBB0vOAtnl5nT+tHPkt1LrnqsR0JqUD3l74ai/7+wklC8TCU7Pe
GNPrmV3sbB7fF3D00hmsJzhBcCWMbWJM04uLC6+GSWSl9iTkg9SXNMOJcpeV
vlo3fjW3XDOshgX04hoZ1q+l39Ws7E1gMKpG5h2IQjP6MJkWXb6V9BhgkenF
/EJ6Zouf2Vz0b25fTy00ldyNZCY8P9LtuRI6ypGmTdkSpDzyxRaRy2hWW3xR
mvN6u725Ld3ZNHzOm7cnYJ7KAGfReRTeV5nWqvTsnjtr4C3LrorMzGAaFM15
vmwR0++VTShp5W15duPx07liIUvGryMhBxiVxNHygtwohlxK1YonTtJmbTzw
lr2qYQNJW3dEM9EMGShmgvPgiPGEoaPhY1tSeZUbQG81uxZgdQrOqtxJN4qp
u44mdKARlFMVYV8yXz7sqAJrLQmpFVToM32g/mJFjq8TsTVGwi1/e1EyTIJW
qspSqw6XPWrKYJQwxxtHj30xxFWkEp1ilrrpceO0a5aquQ0bkGGLFTZgyW8z
Xf9622WrcSEycFVCPDj8fK0ty/ZU0BMbv7XFhc0eol3XmFutGD/i2ouDlFOy
E3NQYeKk9A4Ml7qAGeWF4TlET1KRkRsLHlnl6XUlYb5w/wj+3GRp/jR/B8U6
cNNGvdRAg6wCykqe9HGhxyrRNvY9/N9c1bzE4CbacpprvG8ZI2O/aFL4TdcT
7hSKR6PE1U/5xnr5UW85uz+/HC15r5EcDOJ09o1IdVJn9QsagllAaQ64HS4C
2JNzEQQucCCBC2fp4MLg9tjhp8sWB8y0MC/DsTWH7AdPBGJJ32ZZhV4ZN61d
oYHTu4xV2ayh8goYA+C3ub+eKmqjXC6O1a5W2VmEosTerp/MaRGx8Yp+pVHH
24dJVaBiutYsKXTGaopFt7mBXV7td5581CQL0XuEDBxzntEQRPIzZd4q0trs
/3uzSkWnBjPCzpKB6Ws4x5VPyEdilArW/tYhCzUDhuOXGBliH/558kCxNfm5
o59tz3ctSbaAvCzAFBh/cUhp3NFHQdNCT3e8NiZlWP8Y8NcaYEeTdXKNV08J
vyONxgEVgVMzoh3N6067ZhZ6fN5QRW/6BLUvrc8v6L1xdWGs5domcpj7OWQy
vAUUjr6BACGMWp60C7SrxpvXjUBlyj4FhYqZ9JaPfUB9Mxhej7DFOWH4r8QT
/46IlCSfUOvumTBz5qp4/nog9Zix9lQzXmwGU7pvC4fjKpi3QI6z1p8VvpPE
oSqLsDMICE9/VLJ7pjyXZUjgm10AtxnEZ9L320ZS3Bca5cMazHwKnFjR1zeL
Mnw8ft6Rb/JTkkSzmJlFTF1SDk17Hy392NLtPbALD1ogplVI/MYIzkYF5qXb
ywY7F02xWYFBNePQ/7IDUlSDnBcJclGNmGIu4Owc1bg8lkprZ5u5mWxsXIbI
30OMBLKqxklaPgglu+BobSE8BLy4RBehv7NoEvyCRA0HQhihLifQItr24/z5
CNP+TM9C8T9rn/HG05hRFF2vJ+O1LnU5Vvanoxq45D+wPoMOQ59WbqTEEwXo
hRqkD8w+zI/F7iOs2pAG2M90pBIoWGuASURGv/p0m0vx0k7+6UsFX0N7ErxT
HWi/G43PJUyOxOHVdpNKVpejomudro2fezFGFztR2XokGIho0Jxg9h/SOCtQ
MoU5vQK+r4yS4j/WSzWikeDvHYhwxCtdzeanbo3tWES4jAeVzgasoFtt+KoL
sm86PDOGuKjn7jjO+jW4tJPmP/dG3YeU85ma9Qas/3IpmUmQC8CcLf6hPI7H
4AKygFfahCPxbjGuwNbXaWtenBV/MjEN/P1M/YGme4b0IGbIPexh4m3GnPBZ
TNSeXAK19ZzuUPHU2rODDPzaB6Ej9VyTCuj2N8yXFruKYeVydd80Chmxbh9i
ZNuZopOhfFKkTuLGc6ml8hh9B9kR6hDi7oS7BkY9zuv8FpMXYGlt7V+7p5Uf
ybRBqdVzdAKoIkb1MaRnntWstc6n+yZyDVFWmuLLdizRxKrIUY6M6LdvWFdY
zbY0e53jNIgzM3b5yxNJckJPAJkEYRlhdFTkw9As1jr2N+Mc7ZQ8HjZK51YK
EbJiBHleRT/TkdvM/LhKHvyXaDYe+vtZwTpjVHU7POvMkYLyWEwXQyNT+MKU
kF5BXmIlm4c9ygeR7TAe9XDaWMWDJFNlcMdjERcpwjlvXng40rBN87tEX60Y
ykkTB/kN8zUC2cvEwBOZWs6e+oqMpeUuU39CLIMYO4dLU//8EpG/tgCQhsmi
3EGkLUsjY4xF0+6dqF4bHFPhRLYcPhCQGehL4xuWo33dhRiuGq6gGg0egff/
n3zZs9Q/4U57aCWbqa6Ejh299nJ4J5oA6GDmEgoh6pr/u+aXRMfiCXi/7+MV
ufRP8kfWbHi94/5JYcI3jwwont8MYj+yZQ8wJ5PExhgeQ2CiZqecLamzqVRl
UE+yohPkl0NeyuzalNNPpni5fLdLeeONHwpA5V5bi0+GGIxmMYADXVPeltuM
rbLmkE2WRhDqLN4ILtL/jg2DPYi3m40fqGVJSzNBZvPlr2KaKaDYIa3m6FfK
fWexbrSxlIHQcMs6j0LkQwerNpMOBh+i4C08TLij+oHMJItV7tyVQeFCDpST
E6btI6lsEA+o60KhB3uUHS79Mr+TG+CFDY+ZnEc2iXH9ER5HCgyigRtCkX2W
+WIcIDHyIn7x7I5bSQC3jUB9yyHZcxP+tYOtrRYl0AIkEATp94dSS6utr3rr
fAiZjr8XLqoq1e7xn1HPaUV11NO3WTWfoBawRlVI3sPeY06hDmpFQ4vKZP5M
CdfDnNAOrdTCnp6qUTxoRQ6A/so/QG57QnGgYbiKJ1HYReVrMqozHt/Rgaat
e6J6w6Z3hExyUJbXN2hwxsQoQ9hg2J1v/rJxDmgj3x7lLI58GTDdjnJq9u7k
eznFU0TSvblmQOqEfjA9nTG5NrzWfsTWVFtN4J/sNuLnZ/vWK3sJknY3bR+6
cJ/1Qt2v1fyO3Eh5wEw+1rXOiZw0vlQCSjeu77i1/Cf8p9y7zGubJpm7VzrP
Hnv2YVdtBg51OTQwXnE/T58zC3tx/zifxHpYoAd2k5GNLtFGLhBw2EZqhWkE
6R7sCqOtHQyHqT/N4sAB7doqkcNmICzqkqPmycTEnZbpqU/Tj/Y/r9ZvA1Nx
0FAsyc4cDAkkfq0nBa/Lq67N4qyRi9w3G1w5meCEuPWXsmoxCI0bcmU8JKeP
ikPFF1zuFo/Mzo6xObFxDJTlZZqT1R6bN/d6OFX5CAQ09JzHTMD28hx+usQw
svXTEILqhC/8K/yf40u6S8hfOMuy+EzokB3GpDrR55JmiNp5RQHVX5lwEawp
U/mrrWlHpNA2lHYTgURySic001NhCbaVdYaPM/lbMDAwAWxR2eFY+fcYB/vP
2rakGKXQbQRrFDFNyL3Sq8NRXUspoBqOAREBoZao8wK1Ug+uyNdE0sed5s+S
BwWgge1yQGbgejlwrk78PnRSSALxAYq0IOKMCcfvWAAM7T2AvZM9E57Qi8Fw
1yx5I0qkodz92erwplT8uDXtEj27Zr7MYjBYwGuKqXb0XQRM9fLxY+BDDyMK
tgClec/DXom7XP2QyztXtCNLVhiIK0/5lRKWMLmOQmPwEAoE4ovgdkhaXFZk
NjWHnE4ObXC0Sp5oRbbfSZAF6VSK1oYelsbyJwMSrI4gl/a8VQ3YC+TPVa5z
AkwF0IgtFno55cuycFBIKM4QeYH661t/KBF6wrsc3GYC85/qY5R0A6HuNylV
U8uuIm4W8IFD2EWw2S0Bw2n+1Xm5rcRviCQaink6uuEbWi2ONlpN+Yv20P3b
fbYZfaKoYegrGvZXpiPK729R0QVo2PuRfXoyeLiJi5J/W4wNgZmgmCOiQHKF
Hw8VSPoOr6+NSgMbQyhgVOXqgvG/ArbK4lkpZ7PVFMu3TDJ/8EzKIX/xipFL
rubWOPfx+N6R3L6Wsi9Ps5umgs+PmnQnFcqzSmgzY0F+ZDaplUvX0mMUxkNY
1j5bFOsAaSA0e+TnLwguKntlJLhEnV4LeygaYOqq2K0unRLjU7YHu/6ajr5H
S7W5nTzmXY7PpbK6x8k1FjwArr1PJCo/HFivG77lQi1Kry2EKH1cFSkGCQuZ
fi0MB8VtGmoWqqd74cBSE0mGEj7PlDagAg3yMJBXAVhWisixexwsWHq1KOYe
jqciQjwy7JMGY0QZkYJcIq7JqezlcKm6c3H7Q4gFJYDYsAXNp8DE/ptM9iFw
2S85Q69qFFmDTUyQSHhSN1SUPIb0lx8Uw72InhDi8PCqFF0qJ6tWMLrsJ7TI
KNuIxD4zQKXcJl2vSuqHG0swUTIntWLxGeiNk+kEhva4ClUqON2zAN8bq4Ta
ZqqOtLX1jGvjpT606WQOntAD5UoTu/w56ydDawZcxvRLykK4ahLNRmzhK28X
/safxMCu0iltriGnNz3VfSQQTJYrJFW45NRNp0sTF9RgR1ESd/jgr9QQVrQr
wYenRCnVCHABSLZYZ2+f9NwTFB/aJIOTEPHK6CXP+ztcdV0cQ+/Pg8Egwfj6
6EWhRiMWLzed6u45k4kSzCiEF8007C7ZDtNsAXtxrHq+3RdA0k90qfkhcV1n
Mx/5ugX/Tfd1mBEEKEv+X8U4Uu3jjqvUbJq1wWIEHPZQQAWq1vAaiG/Rk9QF
qd8CnnKa1d0TDIIbC/eu0HgwzU0YW9pJs918kULnkyqpUD6NkrZdCBHCNKH0
nIKt+X5aBfbjCm8XQ4zVcapiZdDUyhPRBrFzG+ReBU5G94Y6DraAKURIegE7
0gOrlf5xoJ5Zqr7WYeTVi4o95aphV8BlWZhrphB9EX8ks2ROBIasCC6Vv+rK
RshR7MLLQXQjuqX1ej4pbUyWmnMLLPlr+PfbTReOnMRXHqnEwf3kNjyBYK+T
KSbPTPsURV2l6Zn0WcwYPKbOFMkX5oujfdJmAl7VG36cgq8mSqDvRkN89mFE
248LXOXblh1R8N9SJlgb9ujlT81Ejna+2T/Wk2NZdNk3Ckei9/J7dVll+tOP
UzrUbT2AfJOWQvftFeqTwOuABdKCK/LQ9nXMOfAlIu3c3S4U/Iz+DrZPJu0L
ertkPKyz3ufWwM1fcJgcmql8eumRNP7/p3Xf0zqaMs30yAnF0SRmgR2Q6OnB
G9pUGBXYYueGpmEKU3myyndcZa8cFwfAxgiK1KdV0sB4jp3dKtyTVj1hJPDr
h7fJCeJdNqhuLN4X+QzRDOESZyYyrg7wIjgAIK5iOnmnXJF5yFC7gi4cswPq
/TZ59TR/T+FTbuKXo8UwyhQizLAv2eXvaKQnXguxBOd58uRVnobNJUQBVosj
vg1myoCBSrFs14OKzRa17ESf6Ws6HS3iJSN5p/H4lUUn4nQEivvmZwPrMuXj
8lNB4ZOULSAqjYZRD7YMDRbldmIk9RTkMpFZ3ntNuqbsywiQYlv8m/yjSOgG
jtKeTwuejmbDUp7Gmf+V156+ca+P02OG1G9UwkwxWAoiTHsBdSlZB8uohOIs
ogBCRyqwGy34Gb98EOOe3mH0SxaBRU9ckJlNQOwA2Iv7S25mSJ1/oVMjx5XD
YUbie5JPesDBpWyHpcH878eDsDllSUkQVySmGCdtATlw9JJlAxYRqN+7Lzoo
1pEG6eSAQ7xYV9kkQSyQAq2GkYtaWbVB3pC73PwrkpWwx+qk1HH0VGjD29ZN
f3ju8vXpBk0If0yj50IxKXF6u3OCWvkGB0IaTVTEkLwOZWsXzeHP4DEdlFyM
/dr1pPH+IFPAUCdNWJ0Mdo82d5ip3wKH32n33u8QxNXP2P3JluZuQMKAI/EY
MWmM9pRcIzS+QHZZUGEP1qXelDAVpK+ac9v7+cxCM4KFHcOd9h13t1Z1pklm
JX2uGi7kYvYARFgJhBUKeZ8V9FZXu+iE7f4o/5JrTJwsFZ/qkWke204Tzb71
p/MJQyAawvavI72Nd/d2Lp0Al/2VAJF2IAh7ogHZNi9zHC3u0oGf1p8nlQl3
5/6cqIEEuVrYRhgBLD+2X0hI665EfVziZ9lqi/ocg8I0fW/ZcHXcUZEUeL3c
LQLFWPVOcaaI99KGtkzkpmqc/EThMxSMHx7hWdReGQkHUtwyTeyXrOMc32iw
HLvOukVhWSQ2nY8b8iQCBIzBr5RDxKvxzS9BgM3lTJEG1+W9DGXtLjysPMpX
uFsmnW9XQXvTLpMOq5dvQ37Za9cMiL6GfcBnxUk6fvYpImcITl3pDKqOveVm
ZIgQx14Wo+LVl05pUHGlkui2HRERF6ZV3ZGNtIZkTYHld7ws/oCVmNUyRzM5
NBzd8qcm8twuaANRvDbDIYCy0vIH+Pclfy8yTY8cnpZ8rz+dFAL7ZqLqTRd5
anAvLEE1KYo3zaa8EdZQMGA1ESkiKR3HiMMUSwrf/h8n1Swq0HZpqYcSoILu
6ZDpXwO8zucXnt+jPxHWqbQBdVLbMGsY6j5q4c0+V7VWTgNZYT9xR7vxfDrm
7Umd2luGL4ShCsMbHZA9XlhID2QfcDbOZpVTaKHVPrGNOy5dtGviA6TSG4vs
dhMM+9zfcLpjfHqCYFcWJBml3lDirTrr6CCnbOJXoJX5KgYQ8n3Uy6qmsTAE
/J8CKfQcXjs8JRqwtVALYsdEImIgLQkNMSZ2vVlSZPoO9q1T28fy51LMIWKF
jDSw9kbSS+GP+ytewb02yssFfqRlJ5JWGiNlkKZM6e5c0L1n5mpp2i7lKQ2T
leEvTiMM+SXtPdBNEf7uZYuAaBt7aiU/pD96ZGFrQzEbTMLWTZ9AjFMsxGQL
Lfv0x9O/0dy8aPIX9D67XSRXXa6gKBs0voUHR1QNezr5AiY3qt6VBfpl9JvT
vVQQgzWsYlDVNhAgENWkrK17MnviZ2TjMWkYHymJ+6TkkTJYnoZ3WWQeutGn
oqG61OIqIdsi39ZxhOLJgiXqpL6S2FXcPNVMYZGLWdpWByFNrx60qj8L8+p4
kkndx0PC9qr8QYIURFsDE/paH5K3jSJwZlGCFINOQ/SCZMN3UkeAmfNngUcd
620AVE+ifR7uRRdJ03oPK0QRpigaAKw+efCyCjgsFQyz0coDn7xAHKA1V5nw
7jzbqPPlHpoAGIAzpM+gk0f1q0GGwxegfVHC9AFSn6oYHaaH3X9VWi641dbU
Qrpia5sFFMOSetdDoCEVjNauYxVOnDVUquOZfmIGclOqz78Mu1MUGJcwsv0P
xszWzH/N6k+FCAsZ8NlO/aH2vnnYZY+1Q5ufan2B7pOCZedq/5/Tf9GswAfo
kU7uTMvcxI8FOAgyMC15UHU+OEo4VMESZZzt/KmshYTx31QTYeXKmrdPJ8Mi
aVW5T2jRVtV/zl7UVW8dwLkDCgeeipt2eYbU96WGnLrXviO+fgWCqth/7o04
FMlHWQQGCHpNr9aP20FKaQ0AB/qMixAQ5QIhHN+hwWT+j+rVsI+qhq7mIjIH
sbeoS5gXMW1p06V/+orybSUva3qrGuCb74bVBydBvFKNFgXn2VJrj4B+NppC
klU0p9ls+ANwB3uNZ9m4EFaXWClNwEjvmfJ5ZktgQTsGFLs2jzlDGCpoLxAK
fWxyB1uwPIYNya+e0tm4FcBYsNKKaGolEG1Rx70HrPoclhBHSzdgxDVdjR1K
/NEW6/3laNrH4sW8a8lqYwAopcNRjS0ejqeFjYxWfqxAJaa9SxpFHvmNI/um
m9MwtNN91VAsI5hBxNmlCHCs3ZhFulYpRbH/3+6HxjyD6e4Yew5i/zc0DZgO
3xr4aqR3NEwIF5cba0mb9gFO0aUGZnmYj+mwlyf2njepjeRgWXLn1XzzraiV
wVBDMJtOTOWUQyzRitUyLQcuMHr6eMqspHWGUeSm4KpRFQjDqhv5NJFV6mWs
U2EC88EUXbRjNcepR9BwNp3MfElMTHd53WcmWqiRiH8bv2WBwJisfaFHAxlz
l1sMySzjFl6ScIbFjgcTSFkCoOUm4zZXEGI0HvJB+ALJfleE1GJK+ImRh0pV
eNKM+hW++0MyvAN5F1O5qDf+eNMNiYGu1uVA+Ti4AFUi5817Xz/303KJtZbF
3UFeZOUsAQvWzVwozhgTJRuG54A7GBWTWQ+MwVHtERoLIvHUT0b7C6lpI5Fz
w8tCEwrDbpF9Lim3OAbQQ5yAqQjOf5u/zKIx3+mx989I2t30fthcCjg064Zq
/ZDfZQ6vw/4vMSmWM8MdKBRiJEFA9xdWbcgEXEv41sk7F4U/edVdQyLMh6R3
CfbVzd33ToUt7nGx0NySANCBHf+yjo9vXDlXCIJ0wQRLmd2pydT2JlJ4gjTy
jHQVz6/OeLVacw2E0+BjtWSW0dBidpTS6L/Di3OucfFTOTsunddy1Ie/Qoj8
FVqlCSD4MmkV7FYhI3aNx3gWLDeFghzZ/XCxtp3HdGx8+abtHJ+ZAu1nFYIV
e1a7CzaKlvDqWNw2EjPmKlExNBm/R+tS8oAYWn9VFb7UzHXIXSemGK8iVAnB
mM6x0yXQ85/TkDBkpdmkCz2CZVf6yiOJ9gHCepT8vyDTTfgjLgvSaYTKx0cC
3F4/X2UdQN+rTWuyt2CnAcmIblKGbaGnJ/ZSikdahNyBemhXOaWgXPJUuxk2
ngKigK0q1Sib2jiDQbW4r7hpMl2g1myGqOIeqCA1QEBO26dP8fZ9VKSbtLQ8
sLBJO5HO6+fJSQd4BQPMlkUt0GDDpK2zb5n8ymsYMFdiABZZ/++ClI3Q63Q7
e1zwsXz50ixnEk35oa0Mjdqw3KkPJGvpep3O07AD3r9VuU8qMH30IcmKlvj9
PduPHPqLEBom4s4Qsw0s4nW29ZdJaKRqV+Hp+d8RZLo7/LtZxuemyzUDU7Rj
zoz4VwYUsggLLRnRRdY7kQe90B35BRlAG5v3YN3GN1ko36gE2RqB49IC1g/j
DH+fezgy0k92i9NsmuHs7xb9yfhvyzYijYXN+gZngkWz0nIf3a44jW1RyJ2G
OMi5q5LNbKUMTmOmflIYEQvLmO3PbPigWn/cm6ld1l52RQlTqZ3wY2HA1Tcf
D9kjYwTdYHR4HZpmTmaHUxV66ixyC7oFdSjXxL5qCvGPyxInBQj8ZDJGRZk/
7bJmNzIxAcKrzJEFT3wlQ4UNyia7tNzNoOrljH6Q6z8RNncfsi0OlF3WF+Hl
BkyCMCgGAKnQiJXgqEJubtFrjb6DMRNLbjvfvZQFS86WUzwbhglDn0I9vti0
ZqZdm6EQjYfVPuvcxu/6AMpOlE38NvagpCjFhyeMUsmwRaPPTlSuMh1V9UyK
ZFxS+3BOM3GhH3ul1XyGEeAZ3x+lnIqDbI+Uu5Xk7peAgWTPlV/LoNNrj9M4
IswOpALlBH/Mc2a7EcrfcZxonmv/PAT3s09s0Lh6NFRugibdlX435OkEXKUh
pYi7BBNIfYY4LE1/e+FWywTaMZvs5KoILtTX/39OhOB8sFhUuMm7yNZUQOSh
lQmY7yZcfLQvKhSb1m+bt2DyuJifdUjd/reMBnXequunWZ6U2+6WJilCjeoQ
wpG5+f18+Mt8P9JrOYU6nrQyy4lH1kgLKENAuP90CqRgl9iR3ssUYHSwLf9U
Bi2N+9FqbM7IPvjQfCpRI+qvqqsByBkXky99KW8z70m26VBJOhle4G1zfhlU
JHsShiy6Y12Nzwj+94KVsNi+uLG0ePCQ4i4fLYzWuh3COyxMDfARRxNlX5A3
3J/f4IildD9GCAB9UOKEXMvusqMphPla5lCMikxoFFPi04/R+5QbaQQHEKQI
V6Y2DxrZ6lDX2MjwUTDxYxjrCO95LlCcTaAfMyS1mmp3RKZC8NeQxH8bSQCL
jkk3kvu0fn5T1UGOqVzKpMnbRcHBzpcT7Tk3RlnEpBxHUX07r5KbGJS71/fv
G+Xa4GhKUkaBl+KaAs+Iw1NV+HSks4IN8GaSha12cSXCOmA9Qa19dWLCLR0f
DaJj6ZLpiyAGkhjJ6CCmeAosgftW0OmHUTH2r9CbUjX3DgjvPgw/Tcr/o4HS
S5YWFRjykDvx4nP36NoXP91iBqio5SmBZOu7NuFeKojqZgm85aUu/f4wDahn
6dWXtoheQaMk2r5E3FZBz6HAunoN2lCbX87ivS9wZIuHKbnizY1prSGRnF79
Qp1Xz0STrvQ/qSJRLTw+WupzL+rhuTyy+ORL/NuXULiemoQz6rCe8TeUZbY9
3ApS4bOez1Mw2Bo+IHTcn79v7nsaNRpRZbx9FQiT3S3lQBMhK47kSCNrrw9l
b4MO+06RVemsBHSuGb+2AtJ7Ng5mwtWcb3T/xpwie/ZcnYaAiDXpMtx+QyI7
YETQXKH/eCmbGCiArhL5bD5JqJQCfgVlw+olYm5JkYDjIjH8zSZw0O6K8TTv
rHNsEnwTqgTS7bbUBcMqLdftTwEYQaW9GzltvDFThqDL4wSSmj4n8Bfwjf/7
g88xJ64bjAefRx0zl77hsPvyCi9UuapYDsXl2WUHz3bmp7Oadu6nyDa0cr2m
+wFh2uKEmvLLu2Fg2/w2W5Pf438NSjoo6MQTEG1HpNiKHnC5RUuymKzGx7tF
IfvQ6yAeejmBbymEoU2k4UfTTVzScLUGe/n4507FonXmPpB3S47YyHpr0m7R
o8HkvpELJ0XKgQXvUWdsgi5RdM9l4WRVRIi6WnWwyg6PDVxt2Zsvy1p0G464
9T5rHIFwCWRBDDZaxMPDZvnA30ixX5DdurS9EGv1KwFl8Bc4HiK3ZiESvIV7
u7k3jfLZNtu9TiuKUuyp6ZYzHyFFe8qeGeDs8YFQ5lpQsVgoFLCH0ObZwTUS
ZdFFvvXqOdxVTu33S+xuy5qeFKWQW61BvG9T8y0DPhVZfK1PAxCYw9RQFlH5
w9m5ogtTA46r1SOTwTFx0CrJopD1YMqF6ZyghqbaMZaRdHCj8YcyBmFi2ORr
a9blB6ZnalJJ37PC/f+0V13BEO8jNUO3iUYP9Crc1KtUp2XxTKpDDD1sMhRU
wp37QMqc+m+I1QjhhggeeqN3Yul/6LhlnOUSd2dk35KJIYQRp5D2UhGxYefL
lxOdYZ6j3ZynU78MBGx8Q0qNLrhQIaWE6XzRnJIBOWtLmKSLvo6ApqIDQOxk
WP6fupHN6gdMl184ZWl0aXmjxETbHQ5wHMaDzd0TC71Dpg3sDLOGx2l7Invd
zy4Lmy5nzwt1J0Y9oICs00C/bLoJX9bm1rOdIEpVBIhl1D8EaHWgkrc5A5vG
0JoHZI0scgyrd7kBdy6aGBqYjqSo/CGl9lRIexQQ4yQWary5lG9E2OZID1u3
tbL//ah2KkO186Wx3c1JizPxbsJ8TJqJpZhfluGPv6H6zoCkrl2ZPWCnrqsc
jwdVI2vFYxlZVy8a+yD43IHS0rApji52Y71WqgEuOdIivZ4D4I1ykBYNiuDV
MmDMl3p7Ydw+EQm+qXVecofvtkpBf6bpxvis55LacRfVrYBQ9KBa6BW1fXQq
gQwibu2qo4wWdfa9eTTEA1M50vT9c2Y3ujzr0CZleRW/drWn0uexSxS7Ha3R
DBl2+vENUnbc6v5G6xovog4+1dVPRwZSsxklbWzE05sIA1OHAc+F+w8b4qlA
MHa5Oz9ntSjR6jI/PT0QqPFvecTbu8rvm+5HiqY4SzSBL0p8xpTweQu7OYL9
VBj6sLdalkl344DpNqiaB5BIyUzJUuk3A1azEyOUc8rLOp5VVK9kXUTmZWmQ
e0HUKrANwTHM/LRbTuy7OKyBO1IAHWTdHney0S8zHPPdUNmEPYVo49ZNyTLU
Mlpnl0fE+3CppuxJd16lFzeCJgPfKZ/EPobmuA6CXwaczET/qjCISrdn+Qrn
9Oa00ocwzoEvdkJV9ohVzSgY2su0KxGAFUeKe/CzCMkY5vZ49dl9i21ixMH5
e3bQgKrHOXYMnIrhEewzz5kLQf3oceUcby2am0uh1FYxQ1DbQAd4f+rnmovY
N9iUptG1/va+22da7/U82uA+QQsdTigE0PQLFfZzzbnEIZp7PnyEEDe/1i/e
IWcaOCScf3aBhrfBFlbuYAgcreXWTdWE5ytVYXhT/CqJRpH/HSndaJnteVl+
Mahg2L+S3kerxeGcnOzhRDd7e/0PCdRYZzwpp0XBTQp/QSJ9edKdOSJN67aS
daCoJYFNbsfPRJIzQyx9QlCQuax4tj1VTSvFDBTwbGCLm3hFp2GeAiag3JCE
xlcGzUvOiCYtWV3hF86ZZ8sOFORsvc/pHvzSOzx/MRCCmm6Z2yiTO+qEqwjT
IQp62J/dWj7F3omo3Z77VpipdpW+VTblkswzuPeTgn02MvCp8vwfgJVmjeoc
8aN2owaMtZJ/B1VuKscQw1H4mZKNJ8dfVZpF/vxuBUAVPpaQTpBIWVIjQJa9
G8F558f4zDCM4mYStZecxjhtlB6tGEcXBFh0BEgIUzQmixxTMLZyYXc6fUQe
LMUYIORSUqRcsY9C0giPnZZgsNRVXFmNJXAlspuPTyY4axrDueUMMIc5QkX0
iXvZzuJoEJ9aai6RrzUMFbzBSAQjTGWvW7Bxpa0kjMi/5ZkeAouw58y9kAIN
/uy97hS9FrPLQV4JgOxmPoWfuSPytzy7qXpF0tLVrsRSzhrykf2nuFGXOQOe
6ijWvMwaKZsSZWV5hh4gU7eHXvuKgPiDAnLPdXdwTJqCDtXbrjpz7sFHLZfj
Oe16JnjS3rUdorw6HYw8XMEWTcq1MX8Jf8ncMp2iFsq/W05ry/SpGk6NCgaS
1bE79SYfuDZbQAgkctCgbhpTBkrZNooY9Q+6d6UJEFtjYyO8R7bL2CUfP9eK
WGObjz6OQoC3iWiIORdOgG2+Vky8pTDKE8Ddqef+tVpu0HWABukZQdFrIdL7
4eEmOUbCdjaVj1lHk++1bk4o1Y8DPaiNiwUv/yaTNa/epDRx9nf7gNLGL6Ty
4b48f3fcKK5C9Mar83BGXU9gcTZ6iZqjTO/ga4GuhZwfPU1erZdopr1khObf
d8irRZ2K4nG5Y0Ryx3zkglgmuCsIPC6YIw1Ut9FHEGheotLWigAAwMSHwmHp
FyDiBqw5Mbly6pQlBHMxbErqsFUiO+ouUCIklDGpd3XOaAWiot2zYxHG9ep2
R0aRplnn0LjoQVaxZ5Au4ihpEqSKWgaccQpafVTKHtfHYr6zmJrOTVoZUDcE
CdeuFXxf12ZCoNjjIx10jhs9o+aI/WJG56mQUNoOU3fMprOC+mezZEOL/eqp
7olxqmKJXx67TDf/BH0QBGXhzH+VvKm405jv2Fr14q9MCNYKuwgq0WGy0rit
eAiVfgn/YXMimSzEDZ5oNpAFXgR3sJbRblKYZd3q3KlQ9TuqL8JQrQPckqFM
0ry2wKOf7WtzoaO7Z13atQdcMl+2fbgIqEf8dQKBh+TOHbfR0U8hNhio76zD
rVMtMHVpoI0tp94wMZDdaDMwAW4bYj534gNv/UtOJKcEuO2KLmDbxcitj7tw
xH34DCq1gnw2PGAzQpE3mX0v3a+1o/NdUWhUObHePhH9knUwCwcNlB3b1pJ3
vpHmY+hitdVZdvmlejnPGOYxPacSQdPzx/NiFTaKptM+bR2b3Tk/UAo/pWLC
jh072EwtiZxRfpXHcpPn07EuafgbmIEDoXWlFAzDHSIqZsOz3gylDzAlpXhc
LmwMAaX4NX53pIk/qOD2PsxD/2HvHrvB6r0zPpKvkkytnqypQqguVV+S1tlR
z3zYL05mPTaZmXqPCDmdQDFawTAMtsp58yB3iSSjtYqg69+aMXbZBi/n3Cb8
EJNrZPUpbPb8fWeCEDCGnj3gUU/WTKaPcCgg6mkVHji7EDqhGlwWl4/JjLBz
k6UgS+3cV6HTJpNz8CEcvDlJ4VHeKzwRXJVUnyzW9Z2VrqDBD12Hw+t2rm5y
mO3D7a3tKTqk97tZDkE6NBOI171AK0QkT4IHsLXSBMDMSiZtSqQsaWCogRb9
Zo53FvnWIA1HUi9hoN3qry03K20NyCLB9rTEG5id53jkkmghIrp31xUjXDXq
PB1jElsewU8tlPfxIQQQmkDohkhVcozqMNmJPJysJoCP5yeCkKnzvAZtGSsx
3ysQnYdR2Rl0PZcSpAxGkQXE7+SZpsuXF3/vJWnButZb7O5mdKr/f3lZcFGm
AZBvqi4LAHRvcwCoMXW2zdC7+acHScCHi0oMCDlVjQ+1qR144p3PnByMbQKX
zZrNbMk73jQxfsVdK2MHcsYAvGyfQVmLgAO7UcK0bPVA5vWTzmk3ZQ21JXbv
PsewUypARc0tc8ZvaaMfwwDfHW0XXijg2yTwsMDvg8kSB4gDk84iUxvQNwbG
WytKxPhpxXAZKo9wYif/76De+XcafxgEdpN829poE/UzreevwIzkSy+LiCN1
E/+IfvbgDdjg9xxOFLRRg2BEPuAW7WMXpJIMp9AOOHfjHIGoc68qF5oCRRVC
DZa9YCz3TFe+q7HACXH/k6nPW7C3dltNy7Dq+FwXD32mLhN4hY3uRhi2YHsr
CaqLz+FPXJQJeZaM0LI9xhblUvts0eJVVc3t7/4K15v/eILgJYGPQobk48zl
PSSrUyjvnTcUpDLYt9T4W78WoDuow2IwCJvSNGXtOdKVM46Ey1NDh/D3oNKO
QmLWwyPzRIhdd7bTAQxOnQbLwpFTQg5xfwrdEtSsEeA1bIjetS5Ncc5W2D+n
z2OZ3gfngub0UDUBasg96QIbQPUymnLgaHJnv3H37qhfdx0ALAus9v04SJ68
1xrWG2Jls8U/vqWyHkwK7c9Q3ZcesPLGLZzWDcYFOr23SUttb5cdjTxB2UrM
xbqw97JCIEvXSsEsATaUmuOMteJWnogBqj/GJI6f1VXIuBBbuJY+4w98fRp5
NSarGmqpCVVlmo4d+7WsH4FqslJrr1RiWuaZsFa+y2zC5HRhuLPnx2CLGSVL
iidinvSXB0H5j8R7iZdt7aKSvFVZ94TLF9EhcNTnZUHpYC3m3xfkS2hfiWCS
A2np9BqP2NzG+M3NXsbabp6WNpofqXLE6VP68QEJrsjXgA/Ssc2U5JJFuvfV
9Ed5a3RPVvSkzHkq4aTZvsa/GuJGaZnwNsCenZqSMaOl8L9oXYvCIIlIxoDk
PhvASHagOc++8CAzzveaIxC/GWbm+JB9S4M1d2pP+zJgVGIM81RfSygQggw3
mNo5Je7zKk0arTNPm4tiaPn9Ywo1/0iXOgh5hDOS6Ba3jqgfF/CG4OrQ9XVq
stRPLnxgYcWshDgLbvhcujMKJG2AiUOE/atIVAkVLEIEW/vXnLY/MDMmyuA1
MFZTi+lCYc6+e+G+iQ5bl50EqF8OrnkG9v2lvxpmI0e9HG4zN7FTInn5pAgw
B9o6tjmOkC42tZjZHKQMpZnvYOVbCBZYomhRzjApOst9xEre0P/kvuqzQBpC
1Le/fR6ugYEx7yeLQqGT8R0UANY7vvTNv1ARssCw8BSQ7vElIyQGbRn2RX6L
Trl0Sm9KAZrKL3ECKDJs3IhRe/CM53BeZ7oV2kaiBZqFlj7O0NKEWuA+7xR6
AvV0XSoVg7u92Oxh3+9nsWlzwSrFanLosq1QSjnsXkk8OkA+V0YRqn4R7/7O
Y2JJtls+zfzmP7Wh8Hvdy4IySM9tshYSgOokU6SFGUybkRTedpFiDA5MlQ4v
1PWJ5DwAM/Zey4TVtZcIUKFm0dNvcdHZuS/eGjrk9yPzaVCYhp16Zfg6FAJS
lWc2F6GATQONb/fgyUGhjOrxyfvqTo1d9P1vgmdlfmWWUBbB7p9CyKrwkbOi
cqE++c0dRRbqvtBxRk3Qt+sJ1Bz/213uIavbTizlyDBX0nQixHZth6YnkuTH
IFOdsshNodwVMvsNEd73uCUk01EHfCc/n4yG6Pi6KxS6EplHavk9+wq2mIeM
jT2ZwNms2if3011dP6VsOhmn8i/eWlAsXKCCA6ywZSn9dPJrZ13Wxqeb1VYB
bfYghz2q8PcpderCPIEZW3LpDp7Z2mQ8pAQUdN0PKvqpIvynX6VABdkkySVX
UPV+2JnyoJibT79EvJZNjLCpd5d4bS8kVsq1fWp8eN7LH6VhatZ3tbzb9fPn
hMlwkMfGXnf6AmgYfx5D5/6QPGUB6Dcy9hjHu2WCv2NTTZXXrWLYPct2Yp2R
1oGuW2S2nM2WAcI5jyapq4vE25GkeufVpezPIGywfd3tR68+ltpDqhUkhNUC
zTPQh5Ov/NnU6T/ThJ8NH/1MRfND4u7w25FWjhFWmqbqueQZHdgCMdhuqWgQ
/M62U33bcEBeHXu0W1vlE6GKQ+w4vT2cfSLTimhij0rVq2R9LAYR9tD7EKWN
NvgLUaqwb2wm/19pLPKvcBqXBJ4MOhzlHN5UF2nJHCuwkhcIjEBiI4wI/aGo
f7UDAcDfIAl92Mc0z4nTP2CHXSSM9XP6nZTgnVaKMkTFeVoiArnG5+DOGiBN
hsxiMNEiL/sRVoN+KSYL1AqBA0HbOG9krYpgZMKjbQ+oMmATeiaq2ZxsQODu
DMD+g54irtKRCiw9KZAc23h1MZXv850owy3b7E7hVmiFFI86IR/Z1BQRtNM0
8gt2LH+iq0AoH5bDLqE2/Cq6OrUCG34/0n/InKhV+aWN0QTVjr9IeKygEVFs
bhHb//Q0sjX5T1sG87dvILize2xe7vauzbHoU5Cj8cb8506X8pF8nrSqA45G
/F4e2IqTkDm4M4ZjA6FMlpiwSRc8YluJ2n3Ed2djNwEo4NFpbaoXe/KFeO1d
90/4OjftwaRrPHOBBJlfGs7GWjRGymC6dOpgOkNhn8fDjIBBspCR5iizDE9K
9Ku6Gkcg6EGq2wyqE5sf/F7hK22tO1W7lxq5CHMqFIbV97U3x8lSt2DoL524
bF7+EM61qcyRBJUvxDVvPdmsPZE574hrxeXbMp27ktfr37+YcLkf2C2zccqZ
kgiPpJpGdTpAmrULDfh4TJvWG1eSTcFB8lPlGHBY/jsRZ9eftpxa8NmJh2fN
n58isessbs2F+j0DU/pV7s5+u1xyyC2OnWSodKpuMJe6MSYpmvWQ/OUGV7PW
43DMds32SDU6mtB4D4QwyoBNQs1Os+jfIMCedCBt4L8VhEtDGglDdJkS+B4W
2W0XEePTwU900UQlDKyw6qtnT7SkmOYdK1mpukhEzwAU4d4ACIi+AtF1cnow
8cMxlti4A8Mfv4NgKa3ADVhQLTzBb1VRL0mnw/P54A5Ci/mIKNQ/92UvEcB4
5RTzXlhyuhg7b4IU+4BtefXuc+oRRRskkreHWZhHdfvpNWpgAP6+lnWRWpEQ
+EYszsvepQvpc6M9cQoA68F01nWgVA3URWV8r24Oze95G87Zxnf67LY3DRZO
LIXai4HQr0o/LrpQ7D3y7XNNJAJKq3KEnETZ+phlVIGiUX00yexpz6kFj6g0
uIE44a5Uju/k6sJyG5PRlefwA6uD2wIhylMLK2GLSBfTWTRaKLz3ZbxKK5X1
fTDF2xRUoioIMtJIKjLLClSyZ7KywFHtgD8ggi6INSgRISFkuuBtJxsxvcsX
NkLE1Q9Jf2H13qTt/4h+Vf+tjLPMnDLqfXeCMZHhywxCU9bEssmbumcgUErD
qMeGqI4Ejl4dh77x5LEVCmggLtl2HSmXQxLSwjtAlqqDnL2lafzmfdmjRvVT
1ymVDNvAX15Ze7Kf/IKyHh0ZlpX/C8FqL2asVTxEBRQKF1eJS9MLzgbib8JO
jNZRcRDpFgL3KmVzFnHjM3Zra1+NcDqY0aj1YKFE9+OsWCUcRkzQNHo2qArj
+6up5uWiAEsYaHMYG3HFAWJ8lhwBcRZQF3AdK65ms3T30dBbVmQiS+rMSd+1
Mb2+G/dNczQEKrJ7UF33r2F2Elnj48GBym3Kzv7f4o/vJsyyTU+ZENlUSj0x
T78Ed1uY3JimCJiMPdf1/IUOlZzDE6EUzaLNVEKOxSJTM/wLSWJ7XuBLglbZ
CQRPOLqVWr0eFbM1fIfcLF0PKC64vDwNX1JzSCzmNR5gmCT/kpKzJzp7HrOj
4CwY4EPfJpkC7BvHP6DxJdKHNbzksQfa2HrpjU7Pu4VnMdglNxmj2vgTpm+q
7vxEXOSKAyP+aga0Kx/mGTgWGEhVYb7baWEIruCBxaiR1+QLihzRSRLOVXIw
RxsS6AKIu4mUhmMzsOeJiNYdbN0ikOX9+wGlggmsk6d4Rsp4nkbnPcx5F/2b
yhpGEsohMzAHK1X+m573unGj70yZDOhiRkoDUs8dAdzRlTDgiavZxAzm8u79
lBxef7Dt/mU/Vu/4RAsvmiAkKAmJ50ZFGaTNOSk9UncW9fKjBZbVFlvJhDZZ
sOEyj2BvF7F3a4UAwGTYVweob2uRCEs6Go1bYZlE/JS96/9a8DECZ2j8agTe
HuFeuW+H9Pa9BmMcRmbD7c7nGtwSXz0TC2tRbGkjsPQTQ7mLnZyVdodjp39F
aqH7CTwuneRwLq198g8K1ijb8RxLPEHgVjv3h9z+EVSbHYz4xiKyBIhCGKlA
c/4ZZ9iECS/4NwNX07SnGumkFJJa5mIlH1FOvKxYQwUADVQpX8imDOiFWwYu
J8oyksPXqeoSE2xm1v8iVKmlndVsUS0sf8MCsNonZoUmPVvmHpucniljb5VI
A3uoUkp7SzX8tmJbX8EF8DU/Jw0hpe3fwzvsakVT81D3NVeuN0byDpqi/L0u
Oz9aOWs+6w/QRFOU+yRhVqNxgZO4eCmWR3t6VC5eRc/gVoGHzDZps9YCfRrw
OQEIpCF+MnTfpRyMPy8LglB0fTbcAfRKoWva4c906Z5FqfqmYG5eS3bzV5Po
aB3nF0750GJvog5YOfZJt3AvjHn+cSZ3AT5iPlrjbW9UISzuwerxJnlyUwa2
b+78Z92vnoAH5mL0NUbDpuIDucuKuMM3UJIZU9QYxMt0GXNSw1rY5wjdn9mP
CNPefbwDrxtxQ1WSRyvqNZRLQWeb+R1ElSm8hIHZSnu//6EuxtYGLolf48Cb
vPf8Q1ukpJxPlS4DC5VMu3joSCF1UdBzYO2dXn9rUcd+MOA8xzbbDKH1l6Nz
kfIKpw237TZYv7bie5agCDCUs7EKqTOOB+ecAqBS/aUh/aXoTwzRrccVjQVs
ecwnq9NkfxaOGrnuSZ+81H18YxNa6AWVAEkbUVaHqSUsW12lDQw0S4nq/OJD
4EursKkJ6pTqKYWSImhl1dSfnWrMfEUGscnY+9NrcZHC6S26XJZyfSkmZgU+
O0h+DcEdmQ88lRr+kvFlzxiRpNmlbQPOQYlQLirIhnSkQBoF5ARf1dbufn+O
TDZkggngeATVih+iiMJbMoi6sPCmplQ7S620449l3CvKsHozeIQU/aJb4HIP
J/FK6CTFjhtehvLSJQvE39Hfw/bVXZRlvt2Ks8oc7ogW4mGRDobeYgnS+f7U
BjykpyLurxM+w4TVrFDo/rbRHe9AU220zhclBE7sfFMXy8te12/Z+IHRlFlB
MczvEPux9ukxi2xpakkoXSsO7/LEuAv4cjYW9L25/32Y8qryjAnMaAH/ZUzS
G0bNf/LMx+Ab+OAM1MThJXo7yeyczF5NdO+HRAE7/VsPOGgEckGpIY2RvO79
vm698tGcO1k8yVxpFR/RcqH5LVkpbM2/jaeccJDGA8EgiJ97kl7QNxkHThlr
2beS//bwP2IiIAZLHMzSouvWojiNF3R3CioP29KOghq1MeQ+Yd3xVevLMHkg
UbuUF8ygD6htsVeT5G47Z46GaTFBd5BHF2Xf8QHnU/akZrNX09NtudgpEvEh
yTk1F89n5nTXYeoDfy6oAHiiac8iVDkWa+tmS6lX2yiMQutpmBgeM8g5OrnL
u8DpdfGGqRaOfz5M6MK+fyK9TDf0BFcGIiDJLuH7DMdI69+0e1YreTGjBs22
9sfhnyw7ykKCehrtHUiBtNj89MQuEQ2NB04w1t0un9WuBZretIO1/+JSbOsD
ROQpcpmEpr++lkd86EDMCyj1iUVV0ZeqoLYEyKXsFiF0NBqHfhvwCtf6xMXI
xcfjZWG7eSGeqU6Gwz6DnFOi38ZKXDfQHt5wnFfe97/x9MvJxdXQ9f7FNeAD
iqfg3Bv4sVq/8gEjm9zFpn90hzPmvgPS4ahw2E2L/I060xxqTH1YU083eo/k
uFAbqQzp+Qqrp48H4fgmySGzTw+U/GaDPw2garZPwbtXagUUXIOQRqocEV3A
RDAVpH+gwZl3Ie/VCxCozA+G6uKulUmAU6RWtYvKUWrUX2j42ABdGDOMVOm0
VX2kgu9V4g9zBxCfC0o2hUW68467Ho3GY0mohqM9ZXJqiRmQun0cNhDPKtC3
M1kYFa9VGIEN9CbcwpiJjwdAen/9S3qcuV5x6e9u9F876nkB9isCDr0jIC6A
diYnA+Nlg8dtSK02ubDrS80vFRbXYqWiT8eG+qTb1KZPLva0tFmm0N0jFdkF
hB/z1lwzhrhmi56+SGDinPYOOEJUpOkHYRfNq7amr/KzFo5PZQnOcP7Tesy7
yoJFRDiDvF2KZct7H9IHBiFNnGZ3Sjz+MBeq021vGLJ6MLZeRo2PjlrRtczq
wceUAQinaKXmPC3/Hio8+YFQceul5vRugEGT0C8CPWOTQeodke9kGaqWEy0Q
7JftMJ9pkZjukMxy7PZ97yYuVfepblJfJbEsjR8GKdcXMNyq3GBZ1pFmId5w
GHNal3sOIqu4asmfCNjjK+02yAicblgLvPk3nzCAB+BghTkdfS4mDegrQ7hX
d/7B73OlD26Qr5uTHOHuH7H+TD5xmJKRKsKVe+2vCzctIIkRh/LUWM72rEGs
1+Qoq/a4dcIsui+MknTDGw795mJxoErZZcbrcRDOErQBk9mhJ/hdCLe62+Nr
Ts6Hsv3aTok8BD50l0X3xPQSfonlFvSHDxBWgp6QuQkXr5U51VMY84+7o4Kb
BwNzmA5S38Oy1lfDQryNrnsZENUtTQXldNkaatGnAhnhEfCBE2gwkjbd//yr
sWiPUqy98sUp+F2pq3Bf3Qf2ll91ek/1OCCIJSDr6fb9fZAhHO6QLKBBrFly
auKTxNMYz0z6XfY/bmB06nLYIHsr0w7/1RaUd1aWleSUkXgxStFYLNCUy+NJ
rS+8O77kMaekZurUtNj/1dUo/SVnRQXP5ejUZ925kW/pFfRpZrQs/BTbc5q3
xtNrd+4anfUtfyagXITDsdV9pVb7SXSB5NLrGdbGDJUiclEnEmdCOCaivbWA
DpFJHi4/gLCTykEtGbrt4SRJqCRyTfySOkIuKMLg79vyDjvxQ9sLk4Z0lOm9
UldzRAiLaz/va6X8bV6pIWRUJ3F/kJFrNgF4/w0ka8OPLt+q4UBjvd2ILaCK
TLVxBIzk9122iq9JmHKGrVPbb0PZfRaBkSjKwcw2idsLQyF2SeKSs69hmHs+
5i+iX/qKU8/TnWgWznKCU+jchXssrSCXT9mU9PQnlktIWZrhZvNe7AgqJsif
M5V7BZ2Md/DZ8CrnkA2tmUAkyylePC2Kykz/7zK4J+YPMDh5hDNwUD1urxSV
vRqzU+LaiLyfOkuZG2wmtHxge0Z456b14gKPcaz4NEBBlUw5tEfw0MxOJjRn
SI2rNDYurDKQd0hWH4KriS9Q3sIcO+alqnqu7xdHWAGQnkYYrkiU3tmwqIqF
LLhdfQ7IaKj5Nx9TwWMgA4iKBy4lDInbwChcA5f1vIGjR4paG6LJO5AXseRs
lvaTyl/klXK9csp87QRdvvTDBDSS35v1jyJKnaadNKVY8btGiZ2M1AUoMssi
Cby1GSimYe0p7dM7bBhmkEsDRDYM/Y49YDPQJcLbPbhpzBeqLoCgQAh7LKVE
9VaVZaeLcKCgkouVuuEvvJLCCukSu0tsV7+BrVIyaGGQrA+mD3dk/OEVG10w
hm//nag54ooUFLzXEoz4GpY2/LJ/JrroB61d5or/7Sx5bPgHEvp6faEU42D8
0SEl5V4PZwd5Jn+wqiPnDQDDsVL8wXt/DlscotRntv3MaS6e4UzqK7qA2wT/
IB0I4BmPwoPOVS5C5siFIR7CNMRpIgPzazf6ggbEgVM1/YlfvgxrsKCSnha+
tlsAjG94zfp2fyiV4IP73F34EBrqjIrL6ix4sEBfY0cnkGwdZtEEFTHS5O9D
lxgl9e4rJsTRwIjhdl081kLmDCrs+NB6sPiXl3azCENWQ+OOb9/aBTHFG6kZ
HSihVuEuQbznQ1Cr9GcHiZfBi96Cbxttc1r7ssqdnA2kxwn+BARuDTFiBmQz
noZOS3xqBxHNzrwedW4NsHNvdAm4IXDZqMHS7SgVQbVJzJS5nIlrGgzTpzqg
Hj379fmmH5zrKBugsFih3WLqzEvd18fjcygWK5nTCLQDg4mNsyA5e5qDkdXL
kx8OQvYofUodFF1LDyuijbNA1saKMNgM9Uk7HE4Zs0YUGZ7UldJYZQVF2R0Y
HNPcSTXdwweA2DR8GgwEPZlbLNfNe2Z4uVMdw6ZJn5JRUjo3SsYACtKdM383
p+jywaoPm4+JNQ8Bk5V6QNs+p1bnd3331q2j08Q9RrqVlm2oHJpy/2FovW9u
FEBkzaw94RSLfgALzM1g29s6zVUZR+9iuksmKF99aTahNs4VejJVoQOeFPdF
2sc3b4aC/E9/crUjeXRZwMmV/baDTLlOYm2YIj8rggMWHjl1dYmNeLn/iwOt
9GIs/y5hZ6MHCtGyaCnxL+Hvh27g2A4zd5FdBJT5kn63QZMyX/IuX8YmKiNH
nGZ0wPnINaxKFxKXIW2pX4d65XyAMw/oaM7ht/rLoJyZtN4XB1kd4BATB9Ac
2skB0PDesWu7U1JQhdliBJvjuGdIG+C2rKc14fltC7hsUA1vLFLGFFZ1rZV6
oXZkD3eZFu+/5tWG6Yyr3NxhGwZFoCVvQ+LgvQS+eChEsKFbjRCv5JjhO70x
cL2TJlerKwEqLSuW+XqzBuyq6LJJtGzjhSYzOpzzFnlCOUdOzfh/KUV4U1KC
n9j0SGFZijZqioyHKJi7sj+ewuXZIiuOtuBKnp5Q9fB+KWP1WYuNwQa4bGcM
/IZFrzV1wCTicNc7elR/yVEZrFxix79gzWJHpn0MjJ4RZhadbChmzFE5fb/v
yA3J8e0+aLEwv1iCS8zktQqseWtn91oGnVC51nRVhVxChemWmOHLa6QDtwDL
BamYkmVKgCr+ArS0UgmQeXZfcpbBH17tr5G+esXunN5oPadOSzMx0MQ5N9mW
xWH4oDZcp45QfpSqwfKQHT3YU9QTF15XJZr8QsEzXrdRge8C3iMcv3LVE9OB
HuPzwzz8Ue6TL8e1Jvp12wgoEYIuOY/W365JO16I06MmtlV8ZfzJ/VVQdhGZ
VRRP0US2vzHf3eN0NrjgJr9md9gwtue61EdOv/b0ZX5JhclUlYNWuOKxeovC
EucT04y561L1LnlwgeZcYt8jGqXjbOvJZrT9xY9GKQoJXKYFUSoZQlyd2/LL
qA3mHF3gsuE6tWJoj/B0ABeptT3tibxteAI/ZydwNc7wmH8X3w21wMflBfOj
v/HWTnjH1Q7SHTtO/vlzRwqWRwxbP0rGVdvqzfldURiwfmP0X8hjoA7hSrjS
LE9Bc53Rj9WOq6+wj0O1Vtd7EGH5eGa37Gvm5Ypv3bYGVLbMyz11GZkVW+8G
oqm3bJ3vy0cIHMyKQ9MoZE/RcXqBIKyyF10n4LVtRfQ9Ygyt9HrSrJ3xiM3f
NApzF17PcA+vMNhD33JCEgZnAgF+FBHgLdggX+itjsdee4t7lRUihgjdmU+R
DM4ker3mAyyde2P52NtQJrZRj9sE1OeOd5DWey6ZAunqrVKdZgOHbmEvH5Gc
8WOMn8pQDudq6aS9oBUs3999ykT510H/kUeXa/6zgahJuMeJOj3QiQGARH6f
UpAhUuwTJFkWAy4dLRqB3DWigwA9l0f7iyD22XtE3Tb2uvFrkmWtqoFh4B4G
QoUNKAdWJU1zqKEIXpyugOIi6CbTe0NOwHDJbTQLzgzOhMKnfgU8+HIQFGCt
SBDbJroCaqyfLtabd3yZxYcVwLLpeVu1f6zOTvKyoRkeKR8yHfmrTAAcjzXB
2zAkRtRGpuBvFJuSe5DztV9bnIUyFDww9e4G9lUJZB9RtgPPUFvGkhmQWAYT
M+w1LPhzYjLJVXa0YT9y+sCT8UhnAp7NdIiISVM9J4dEnwiq5Sp+QIdcdyeH
KV7Qyvj6dFvcoaTCqD3/ru3TbwriyLH9U22Lg+e/Cw0Yxhfztb1RTMs3IKvm
B5rirrM1XxNGsJz7beeMoKU4OF+YDNvSneYcgg+DOJ44rKLT0q3rjiYpBUXv
39jjBiT4mpx+6t8FIIfZS0x5Z4GIrXHYjvkaLeM0cLBdQNuC2wX2r/7wD4G6
WAbBSFItiqC2H17kAX9HnfKGqKQqC8NXX6R6FnefkTPSMDlsxwaqd0zZPHM9
StwXUiiPIBe+sFmCvMKuvPMp50ghL9Ap3juO1jEqNthWjHMaR8tzrNJrD75L
9CPLSn1Z2YVicsON0tGsNIFuFfVRO3MKLJzjx0Fbe/XkhpxqKEMKemMoDAec
8RiZA4oq0y5uNyLr6AiA9BAewWGjIy6ln5vmCMzgE/oR/z2DM4cM5ygo176R
ozQFcxvH4Yc43/r5oYDpB61cOtPEk6fCGmOn2qYV8Mo+cmoJn6JSC4sVAumG
tmA2uklJwzsQCaq56mXgJGg9czyAYnX2b2sLvi2ovr47cYnR0qIcNBr52ui3
+gCB4oVymMjiPCshtAP6wNsvmkYuhVuzj+8IzO+wo/UytXcQSdQcIhTWVRVg
FOIjJUygsZnZoQZMSn2KX3u/EWV8hcAgzEhnDUnj4b83pKteaLTs0nOPKLjN
BNXCVa0RjKxdSaRHtmT9RecYx4OcePDhmccMHb3MumRuUV3Y3C4OC3ZR1wr0
QtKwIGA8XE2DdHUhIvNqga+fnDkkDMQhTI/LqTP50EVKHngkWdOdX/sWTTuW
/A7k9wBAL7ZBh5cOdE8+8Py8hjvu9GHLb7ThhliFQhN38quAENyoKs7P4x8A
9WFclrKe80FTrDv3p+tuR+6c/BPw41TLDf6k5bMcJiw9VIl3Cnr4s/luHZUx
g/CZ9RcrRX+eq/DkuDxM4Kd/TR5cfnnKsK4Xo7mMSRvl1Pyx2iWrtPwepkry
ShSz4FD+i85kEa+WDPz+AdynNaQHqdUwOLxaZ2g6dYL3XOXR2LC55YnVxJjY
IwoBuNjVvkeC/AD+XuC6MZGLpYrpHp9bJ0153o2VNGTnh+p0msplUYcIxzwk
EDNH+e9Wai5Z1GoyUrur1ANrwhk3hQZYtFy5LzGllsBinmKG6N1Y4/k2WrS1
WJddtS+swN/SsyaTTld54C5aPsNeFi8pbJ9uEJVoYK7z1+B3K4Cd/MytZKGV
tzTMV79ain0/qEUQayyt1Xtl9kvvSj3qVf63J1abf2U5MHwuWdQksj3bC6O+
IUPwnY6ip4BYbtSyCi9fWVMFs8FdsrnPuGZQBdi+GgDu2vXo3W+PwXFdeEdk
+wfBxEAr3Xck8b2aSALtUUS6j+HfM8nCaG+lgGBMlGcQtDUJ18B78+d3jxPS
v79X0QmHgThZbTPH4KTGiW0Ju172luzUjbB7J+iLV7e+ko37q+r8tCVOimZE
DPMurzY0ypURr+oSgxv4z8jRFkQofn2SxBrMuNANUVe6cagzbcNnJpANZmtr
gp+yEWb5Uo6SbFpuRXmBKOVH9R0JX13RDdnKpvEeR899Jq+v6zyhZFAq4gI0
ZFu7OmCr5RHowrCTL7fp1VGjTeLyzNL/4gjYLX2q2f+O7QeHk10lVMoqoZVs
4yh/aqrsGf3Zboo6wdGNu3OE2Wtz41Q4RmNAFKVOhAum/TtTX6qcJ86nbpjr
fdjPA0KUffEZdl/bzwllp4Q4TWALu0Jb7kLoFYfya1kSgHJGi5QbWtqoSnYu
b59OoEnfyyVy8fOB2bFsFkbDugr9x6raZ33qXzUhh2UfWJ+JbIa/CdDcgCyT
QQBiLSrTcN6imPRm/vcc9KiJeXOiP5uRgC7Xp9wK5B547Tn0hNmLn5dMJ0ka
s3Rtm85Aspk9fI36tVsRqX3uczIqEs3KgS55UxASXJvrI8Yo1QIjBZeS7RE6
3XB3Ie99QUtzWFHVkHjwRyD7abMDJYaO0NqMCnRnB4jYPEEMi92dZ21lGOz7
SvtOcIolnYEJtKaWSEscoWw6xpcL+bjPTxImQ8+iQsJeLYx0i3gTTFkoUaqp
bClK72RCSmhfqjF+nw1J8yy++Pq2ZfwnHxQocDZ4wyDyjG6bGiq3LdHZgFvs
FLRigSu9MYc7jDNys5WmJcX073nsNC/fyyQGtowrbwTQ8dHgUA0fA/NNY/as
JQFelD4pSI7ell9EUPTKaAAn6vV8S1pnid5br8Xvtjjm1mqWjPLY8uWYCY8z
9BC1HdRkPGfe7g7tc0t3o3qnwnV4UxSF4jsycMW/psv8IJRZi37Eve1T0Tf8
KR4MruuQyfZmTtzy/DjxlAi1+7QQXdBRKPWAcpc+Y/QuSluRsHxOZazqoj0P
plvcVSF8G/RdQOjpFXVZcfOlXS1FKa/0Og7uTPJ0KYOf9QBhubN9tbXc5O7C
Ni1MULgKa6nImjYUa6LhnwUxO/WHOLMjnoNuQ+DHK/72u7Q16H7k65YDFDFs
51/5ueXvFFmf+aiNW24kKZwyb4yLMjeNYeiNoDIg1BEEUPFl4M0H7aOr/jcU
pvMpxPyiL2h9y4ioBfL83FEl6uIWJM3gsKkYhziAnasA2LnVY6lVb89P8qfX
aA2FCSzL3ilnedu1Ur8uJOkAqTsKNRdJdcrcVNUag9X8aj2VsfdsqXMqWBC/
xh6s297Er+SBBzwGLKox/DXN6OL4PJhLw2RNQKZbI7cQ0EPzMGR6uBD4MH2V
rzcym4IyGV5HUqbMO+vWWYJrd+KHEsIMXz8vVK2LSi/uW4/1dOZrpr6cg6dF
eGejggyN9DuX7ARDgTTp/MjtQ8bFvoDVsQNK2FTwZkPWpOcN1OURfv3bSY/e
RnaiGhDROIfdWQ/VH/O3n/wVRFlSTHUbk0/6be+f+GDjgsIChgHy0HNhZKUK
Kka8B2zj9maM1DxqmuC9J7sTWWdVdXIlD38VRNZOYbdBFHqAmSmo3/2PwL7g
ZOk3iMTxjP0w+S5cB2C46weulkhbGkIkxlii0aY0tB+FRaNLI80JOJfAwaos
q50f4me2cgUhRO9mR/mvPNwNBv+Et6i4xk/X45Y5ZafI3p9t+LHjcLHx/Ejp
RxqoFUt3ehaASLRkuDjS12e2swt4DBJDJeC2Hvto/324JG37L5wFW7mArjoe
WRFuz27YxfJxlEL4jCGIm+KpVXVFQPTkeUOdCa8tW/3xBuWTixloFdN2PSBa
9YplifMF6J4YAY13K9dH3FG2eBguq9XG1U+U2t6li/LrhB4k8FNG12JCOvz5
akjSXlmFTzfTsEulheIVQNiRz8hymknMpqKjiPZbuZX958upc27QN+2vnlyA
Mq7lZ7SiE3q2Gv/VEDr8sDqbQ3UHAHdyI5lKmWpoSOtfmMassY1/k2ocYKua
w+hLeg4zAL5cB9B/MIfFjJSZGQ22n7L0SlIXDsn0qZaXD50mTYhd25Im2C71
1csSruSdb6w86LXr+FBI6Dq9MWpOpsNKf8thLcwoIV3sycTJ3Iw23QGBJPSh
WU2RhqqzvdTJ8r8dy/uRD1j4xAzTts9vCpGL4zHKqviMx/itlLgME8/D8BdY
4IuykSymSx0GEwb2Fu6O57OhfXyJ0Rj8QyisFok+QDAuL/RolgvF7Jv/eBoN
pNZUshYPdYxkc29851DhOBBfJGxs65Ya8hquT9W4tOvpN1P+H4u3H9KXlU89
H9dEFZ1YBan0fsX0fHL6LAK+WZHFz+7d2bWlwRaeqA4G97xfsgr+7c/RRm52
6/4m4vEqMGGwO7vot1PFzxG+WCM62YAJuZWubi3mOxW+gVdMzcvb9BfvclgR
K9VgoBUCxNriwv1ewfeQgkkuHq/53nfa+Leb+Wm59DF7siV0Jo3Da4f0UyrO
WLBHcsBtxRvO/xmQ60yUfdA8kNqJxboCVJ4n8OH5+BgWerL6bt84gXD3CGxV
zyuGoszb7HJZ0SuFwgJhWYuQt+FzJRKFkp2By83IkKt/BwepTbriPFDEwQx8
x6NFIi/CM+KOtlFvdA1dyelMCMMMGf9TFfmpd4XtraC4+M20tpW8IzHDpcni
Zxre9iouFp5RlEcIK9mvYEWDNwod2N0+n4RYgRWc8YtfLqqrgKznRIIOfZCf
E+sEBYggcJAioyXvvEgxUGvg3+UktIHDsGd6hBU4oygvs4qFuYraHpPMV9JM
A5EEJ70I7LC3cPM/CM/uvZI9SE8BFrmC/bB2JGRW6wxkjxhp6epBizVKGWmO
IQPO04WraVD4a8CsESKZOIHwzLopPjyWYj7gqgwjXs+GwwHOFCVW9KQA4axZ
uEHh4gA6woDJVNzh1Z16A4OGdDas2o4ERKdw+YJ9BRPSWlpehEio0twARrCd
78tfkTjF26Gb61s/txmZBxajrbA63s2Tsl4ekXyh2I0z68weoR0H7dnSla9Y
IzN+rFmqZf2WVlriN+did4Dp4BjbZoIPrhyA/IGWiYuyx9AmASY75B8kzoVQ
rAqPbb9OSo4ACBW3V/VM57OoojMGa8eJS/lc3/kSgjVmgGB/B2kz0xIHpAo7
LzpYA4tN12AanD5RreddpaMz/KBh9iMfx/ZWFd9KapRrAru/1A0BJ6CgFI2A
tuh4LnRnRdWkCg7AUkS1dMUBaZDsw1hcYHHIWfZdxKTGXNbr0mpSDSsuxPTc
cTd968TTA/13hIr9F8fZ1mkAarzmKXD83nke7p4cnw3ugc9VSZs980kYI2jc
aG2ZZ18TAUsyaTbKFjG0hip+mHnl1vZafYkTWMM9zg3mwF6kqmfxfLZ0HnBs
pvqFGajCaGqG5S37fuKtKpGR6zCi4oou/u/vj2+6D2+wfnymDmLSyepd0cmT
juwPzXaL79fSPqo3G5RaMu3PNmc561a9+kdq98e428tfuDVBdfE60hYHohnw
QPR+pmVMOn3A4lgPjoL/GZHuALHMh+QEo521Do2FOph3Dh7rTbZJA6BC2DdX
WvFDiS06w0DhUy9EQ63FVL5fskbPrWnDJ6aNQMPMygX2pmSpJLOndYu2uQHr
OaXt86PjdmHlOmWQvwZD6RSrs7LZ77EbacIIxUhU3uDjbbceyRfn9+slrSoy
F6Kc3FGNiZQL/2qTuyO6yvoWvnzlOWR5+MGOjUY4j3kyMJ6U15IHlzKDXkPB
438+DF9qzXkYnrVq4CJIfNHk/Q1EjDl7S2UzGlKWuAgjiD9IrLUPy7lJblJI
32+G6e3vT2lmEjb67oubrwib9fontFYLXEoVkdvx1Fx29qac9L/SwZnZTSop
GR7Gt6Yk23kCWWxQBFCai06sV4m/mhyMmWAiSaFWl2AVES+26TCWRKjOUZwu
Fu1I9Vl0TtECB/JyJRwi9GFT+yqQaOKObvFwzLan4NUgmxXM2x/+EQcJSuY5
D9XgoR5+xfXDwqczKo3hnBAYH+bnjnUkA2xtn3RJCteyLPWHjN/PXqhL3A5D
/gGTjc3AntkPSo4xyuaownCc7ZMHAPi9n1TyXQqX8j2K3yY2yBWGjA2JCBKK
AyJANGS41/FTjQJ2dXtIRhYdRDoIQCaFSEFm+/Q228uemCM44TdwpPuCnCzN
19bXrHQkp0MWMvgC4n/Dv5aiDfi/WT2v9aqhVYFORG35jkyPq6gHEs7Dh8Uu
KlzEFUCp1hBsnDR7aXjxJ4Gs0ILjWBcBiWVgG1zs/YHlR7oSHGHWtyhFFjUi
OAH6r3Yri/gpDMd+Y7BZEWcgeWIopS3YxDBQsbjq53UGRrC0RGBvpoQKglVI
+D9A30JbttXZQ+nuteMPdEmITzRVaZ6xQ5qPtKttBb1YzDNygXAzyocjKT/X
R/W5kJLtt0ToG2zqDxOuAMKDhZ7TztdzseKF8T7kObE1Xc6OZ4SlBZd5n64h
B6wX15QURfZgxTbL9QFRdtwaExdq4PyGLE/7TRUiAXU11sO06W+Xt67Fs3Jz
zRd+ceCxYw6Pxn/vpR7JDpgqHj45sv1PPeiA77oiE4q5Kc4fIdNHSGHnHHrW
i1/G7U8P4ttlYkd9rW8242lGYRft2AbH/ulHosxWp+I3Fu63afr35j33ylce
WuYXbzxFWuIgVoVfnNYa62tcfaznMQVnWnb04QO3i9zkKzzEhM7NGcyyj20L
GSnq98r63+vcRhlyKqi7RrdmlwvhmlgWxDBU4YfiZnOMcVHRbSv4Qj4uElHi
BRe6BMBwogq0ZtPFSaSoyy/1atSbdKvaJ6xFcLnL97+Q2Efv9sWFe6O+XZG7
QH9FII46TmHq7eGGH2ShnGaZe/ibaazXEGnNaaVG4VCmwlRU6N6OhoHueFv/
GVvLGULZs35rIky2VD6vgz30QxOVCjW0oAMNDnirIFYIAjOPdRJPlZkEhWGV
wvtpuIxUgrywSr0l+m3U1tjHKPei7mdcFA7c1TxhwMVTIScUabfZLXPjoYtQ
xOZUOXegoWaxOfR2rjH1CTdDV7ahy4qoPGFD1dQDoBAC4Yolb0vE79J7K39Z
Ti9Ifa9qOW4HMKsuAqNZvyjPtjatLgu1hYvbUBjMoa/yBk2Pm2s6wolC+LYZ
KQMYF7w6I8DQKOcpS8LcjpIp/mXL+grKyNF/PvE43xmdaiDY1NBKm+N9bR+f
ftfTdy3+c1PptuYfuulnN4t+bqVKyhPneR/mTxY4aYSQWXvgNw5jGIOUPxVS
VWwrt+EgxothjsfQjrzZCSBCbr8f07BSzSHAplxSGEM8Oe7w4ca/9iH/MDZx
TXNCPYQO9cT88uF242biwVoN3g7aUVqokPr2KJIO/M1JT5vfNi34geiApNl1
GIzyFRYYPiUVdvbefsBaSWJbPOXAawkAQYpbFz6kMozK14wKpvZiq4dbD0iD
/sw3W7ydqv4gLtYu6rdI/o5UfdU1KGWPUA9pweSVrMIpja5cGYZALwfWbLTm
vHG+xLKfQjjHpbOTp1nqC9W7iKpcbyjPlnddpLHWLeFwcx5QEwZ6ZDh/MF1q
0/smPXtFvwHeCEtpvayoqDKMbePJag3uYX7XzK+ac+ZDAN8dxg+GhkF38JF+
VOKIUT6WreSKW+800nrapBcQMcEHs44AQsU9nj/XZdKm0cO5Njs+LGbm91wT
4n96Jr2UqFKTda0f+NtL9JjnLUnxjcf9+fmyYEB35m3z2jtWEP4jIcAVa5t2
PlWlge1MjrVmsCgoCrb9Zj4e4l4inh7z5pYRbvx9KHi2kyxlmKY8D+MbPtur
Z4dGjF0z1hBp865jP+W8r7Dc2R3erjaM0q8M12FEXdpmW886YBMMHxz3FoNA
DMnFaU94kw2FDUXySCEzVL2TW7C9B34/2B/361/5zGG6qiwTP1uD7V+Q9trY
BmQPS4BNdimrPA9kjyHDhMMYIi0YUmNGuSnEUNoxR1K7qK9fuSWk8GQq9etc
ExG8icPSKf6+B8sTytpwgImR4NlSTcPmfS5f2jhtv+rESMrx6NPtXKjOE+1v
kvqfom7CG6l7IVOCWulVp90jxKUIGAx9PW+lk2CI1y2Bs/E45mxHbKb4cuUd
ALZ3wQeJ6AtULTFkhbtMUz1MVxRZr1dphSaR6uD8dyBbDmHvT5QlsmDjc+LA
BkpJ2cMpleRMM4acxWOuw1w8Yxb+UjB1RLHWcXZonE8xBQ7JljmjBQg6zsQg
69/mKmO2lVTzN4kxQjHwmSL0bxCQruFHg7FHK/fVD7PY+qwU8//3ldElPaui
dUj5xjnRyYaFFJwRUXpYWTxeB+M8azhBjYAzKVb9N6ZymvBbARaso15VHmZa
9g25bBrm/TNmBETFLJms3o1nz/g6cM2LuAJssdyX16myj3O3BqGJ1SizwVfb
RC2q3px6s1gtM2hZurIKEdyS4WsxyefUzQIK6RXuFfJD7pz4B1Yyu74gd/YO
XopEWp1/Q4ZvRhwdC446udWM2x9Hq9/vExu8UBwlb9QW0rxMRCbASRczWo1C
DGmHBqYSMMZERfbSyVj5IhV35kGn02C+6WaZENpXGe32llRvCtqzrdodDi3d
CQwFzEcmfASuh+b5G6gqztYWKTFBZvPZ+j3FZ65EoVni+TDYnf/JEBdrc92i
P/KfuwiE0ZAEhi+/uMqdZxz1Je+GCOicWw1iqywHouy7PocpclQIaomTsxL+
zut4qoPQzqm0MIkqD1N3xTOQ96aqkgkAz1iUx8E5ChaXAtKiTWloMBtpe/it
uG5g+RIvRKLxB4n+ylfWI5a0k/rFxDdTV95faaAAUa7dWOvyYUQzt9iaYBqz
x45WJ+T4QYD+VHlZBa/0GZjc+Wv1if/p6Opvot0wAD3VYwmxGzIIFQ9gr9iL
Qu5b9DHWp+CoT8i/DCFLsC107mjkhHSMT12cXHXL8i4SKQU9u7tViGAWn9RY
LP9+nEaBz7Z1craofjUVHzYSYm7PbG5KvNIqiK19/XPjX0KC1Y0bDPbeN1Qg
JVtFN2DKV/IfWDt8jFiukir/BkoX+MTtOHsN2j77g2txwlKC7HcOGw4sNczV
WCfbcQ5/cdZhxnz9soAISGPaSobng3V81dUM5XZQRrQz+7++dDM9zpcqvtNB
KI1Aokp4JrKBY8euyYM64XJYr4WEOid4Cs8BN0YfkVpXgkB2MxIVMf+b45f9
5qlXPBf+cAHz3ytiH/glkybifvitkmXg3Qpl8POLPYMIu0B5zoo15WlCMxBi
aD28iFMMzL1LD1eDXtS2dPQeMEHjrb8xFukqkvUtubDvNIMcFSrpgutaKLdR
pcCkhpIltykcnaFhi5ZhpAcSg9s3F+ISfGnOuEd2vJpWvJZ70CpNCtZgDVQ3
vkQNOfGmsmSNKE23Q6se/4lxeqP0rUIcqF52PHJWuyzLyk9sSZOeouXhSTR+
GVbanitYiEuOIFruOcyTP0Sa4EpcKb6mr+2RSJQn3cWzU/8M3A8BskhwXHVj
L+rySFPlwQRr3APtlBxCJsdWcpUtDuCghiBXp4jbNifEuCBwxROsmIJM7F2r
rGgzPc3DApQpPW1tGYSP9Z2X5SA+CjXn4W1yEjpHuLvSZ6wQDYbTZCMi5J3P
Zkb5VZkMEtFGHKcblTSxyYPgNSpZ7+LWf9irPs6mbn75D0sKoYe9hBAntMzs
fIds5Lo8hWZ5eDPcWg1ft426+fSACmhHCybvm2AzuaXI/W66TpBYZY+pLM5H
3W8UQjVWqqMRjz6pwBPPzlKNteynczRT1+m71u/R/OMQKUkVLs7un2xz2pdn
YqqxynXUlCwg+L3woTWev+FPDsRAUggVf9c0oFsEND0rqqAAWaXFrTw3j4vt
sok1QgTmf2JsX4lzLx3kMpAhqUrbCF8VkSus161CBbNX3OQxU8NmTStkFmE2
ed3AyjMADHNDRQZWsbWGN2gCBT/gyVz8Qnbfgz32i9nrVbRkL/iqhDVauZzV
TlcD5DIhbbnIfmVNxxkPhqOJC6OPsRAsVp4BOLwKKnmreBgCMKgEsdWmuG8G
7lH+A/tvaH4yXN5xlEtCppzlYTEYJjTNK21BZ+UnWuBpUVF3skDYw0KzepVj
AIcy94yhBqnV7i+NDmm8UTPaGiEBWKmm+K6ZeCAtGyBBOPt/tSQyqheTj9ER
Q1c+J7dlhcJePxA9wy4m+nYhgjoNJJdC3Zqz3cCxY567GidUg0fj/yuQQyzO
/RVEN1YX8kys6Flw/2CiucdTk5lXgpAUi3rxcLpXGHDZY/37QiuAVCASeLlA
OsvJZxG8OQ3dJK8VKM7TuIzawKheeCLWP9LS6H92P42dAhVImQJXbWN5vTNR
cwd/CO/tp24+Zzoqw0TV4UgJ68Cqf4yhAhXyN7LtfWJRQ49hVUo9ivMleP1g
c8Xvol7JYkNbU2lJ36lf+quF/h0vNv/FqL9lx91Hc7pIGWYORgBGpmTwBOmG
1HUbZ7M3oBZqDCxFvRRvU5K8HZSqMXLyUhJ7Qo778sqsOVEaJ1eA9IcY7J2W
VKMk9nPZoT8FdD0Q18RWPT6ryS/+JWaBTc8yxEW4PSSGhy34ATh93thhp2CC
+mvcbaL12Lb9sVBWMwUVlEPhGLpZy5ucFG1tCU+cGa0e7C1s6MXLAwMz6qkF
pnyfViDe22FaLaagYLshd3oxx13kj2lRwiSoUUEgR7XFHKqMJa9axoD7Qf//
nOL7YgEMQF+aRQFAbat8F15y4PfttwF6f4wNBNzpzJg8Bo1zVpl0PsPDkF7W
CAJMvAyXZ7Ire/UAgj9GpUWrIC5aCrCogh/DzFEPYGvl/ysSfWKkfGSpd1hW
+bkClWxaWGqlH1EbWWHAG3l4qT9ErJCU2iNJCj8BshDc8Yf0yXLNx60fJuBh
saK72ZlFB+wQ5AWUWuD1+4et6ZdeXm+cn1R7mPMPyNODOywHIFFLcT4c3AKD
MizliJm8HiBVes1IAK8CnyK+EWU9rk3eUp55Ao1IqbO1euP0NfezoNBjFsd+
z2S1ahiUp5tlv7WKKvK93FD7UO+ATjWp/mhK0+bQTboFOLrvN7uLBC/5fChV
O3FGx2sD+lAUlzjPTSdsekT+uHGchwYq4Vwvduqf0QHL6tJP9754s+Yj1Si9
ICK+dzcBHc1uHMn5Cj3FD0mFgeLzA0ux56yqsnxA/edbCf72ZEWYXOACxuXS
AaBB6hC05DRApde8Yw50bM44OH+uluiALSw1oo6bMKNA8Q4ZnOzLy98ZnSho
I4yIpZvq2BA1ivz9/CwNthlMgmWNdMAOJUpbuj2Kn5cJaRDiDX/ScteWwtM1
tNWbh/YbgRUXinBkkwzzSKN4INIlnv6aYTUOFWXzOkSelUfIpCnzYx7H0jfU
2+vLcXw4IqGSjn6RbiC4KQS+FAfrBHbuGy2wW+Yzd2wgIXjbKYUPrBOG5hcv
eHkxc40POEJib6VO1ufEV1HlGxL4hHSj/mbdUs/oFY1EPwZkoz+WsALNnFQI
4wwDNesWcE4TacFSBqMSGoy92bFI/SqMB7MTy9LFVh8Rq2932iYfJRNNT6G5
5xCBUbeHV9w10WXt04iGn3iXM77E4ZH+kwHwhKBMd+vYR4WNla7bWRlSRcR9
0L4pZCm8N0ic/TJQIHD8QDTn+2VhtDJhg75Nw4qvVUOSFIgPHa2T5Sd++df+
SLLLzIq0nU4ESgFY8Yl1lGuTL3NNBI6i5w/AaFXa+LSUar07+A7sBv74AjeS
lA/qfFkSd1kVnFtlOPkW9LJ5zeTxIkpL6RTPguzKhr2T+wJLofUfxBIg9muh
n90MNSbyFiPJgoVE/uiNSuZKKSX0vgtGFAz9/y+Pn6EXV/dw5xKv2utE5HtX
ZpmKei8Sr1iGRwbywZqfV2Rb/prcWtKUelYnVsK89NlPLglbpllE0XEoKERe
P344w03g8S2A3fNa0abGYnFaihxKz9Ucgc7/PhIQ3pk3O2gBgiS2NilVE60G
+D+y6C3IwE86nj4o0UUb+3sBqMO1QvvCz8Qr08TeIqygyvyAJoixRDEPQQNc
3AA4Xo/gfbX54H7riEJgRxaNcenQeAt4AXr2pW5QJF9EsOqPk/ZmQUzfViBS
Mu6IbEN/JobDMfv9jgDbRc4eqUfDG5FAHKhHf0e8maLQpXHFfS3Z+XqEn/aH
AaPyGMme8D14mq7vkpO4huY5B7jBog5OLgVuFQ4OhejHCNDTd58McgtCU5Iw
UhJDKt/qH8Mv4V9e+nyHzX1Nu+I4HwWQpkwzq3oGDZA8twWV51091NMFXdYH
R+BkUFKkkJ5cl5AzrS6iHp417Cv9ubQjh7K+Pri4e5tzEs176/Yo6WuZc4v6
qjjGb0XAYhT472PbtYaqmkL5U1smekx4CrKmQyGQW6qw60irYdPBaGH9yaT/
r36VzV3TjDGIpU190ti65FB3QseFROn7Po9R1EOaIN9TWRplvE4FVVt/MvSv
YdHZ13S8SPBLGmgEbV4NTffnbYOYDfQWLxceINO7gpn08Mdo6o0zhiHB1a9I
MnfWt3EnApZ6PSkk8TgZq97v/nd61xuDMZH2z828iHd7hmHCw1LA70wAdhdu
ksMGd7v4OsaH2qcK4M6iLrspFJ0S3ZQo86JL0uYJ0l7TcV/EIGPgvmQnNGP5
QVK39geGKqors+f+kTOjT2QKFDfNV3K+J3TvbDkf5HEH1xxcEXnr1eiszDY7
QEKRkJgZBO9L0cWnM9Bii66hXad9b7UeIcuAh1Q1RBeUnIpyDASdFR3XbxLN
8uaOrUEj5+AGnRflCfuy4snWqjT8GstE/0zPfX30CXZ1gFc1vJRCcyXEszHs
R541myROLrGhHk0U8QOkMcA9AIUCSCEwazfND8HiHp/QwnZ3C/WduJHV0LQ7
BBvHPkd9orKeFjoFtv7CUAtE0MdeV90aTG04FuGCT+dlEIez8gnEITvTtRd+
ETq8xGTcJIjJadMxsUxm1glAqGDfCoHh0j2BtOgWwaYbhWm5boJcTH++qfk5
sEzGgB1JfCkpOC8BKSGwyTbkV5phj0lpRycrhzHKJ7AI26osIulpq0rfERfW
+zxkainjTf9z8EZvguOF0cnlP2/cXQYwl3DS9UjMsaa+jI0tnuQ4oYY9DWyP
dHL788zuQeF2tM0YiHmQKKKp92jf8pbykbBYl1NdxyE6FFkRNugqJW+X3s/W
LdcMb7H00FMmVBIab3Jbkgb9xhODQOXgzIscIrJGQF6j4vwcqaoIXC5AFHAW
qndKfRim49Ymtr2ZrW9NwuOZUfXiMQhiL/YftCMTGObyQ6znubvvDomQP7r1
E29AWouM2kmH1tvz0zOlK2KavojagoNP0p40VeBxJExqM3XW64nYVE+oMHOC
aS8WwigOanppIuVt3yr4Lw6FHrHRT190NaDQBa3wHDDfYRjkBMHwXa4rLPW3
93fYCLHRPNQ29V48aZ15FUL4W2T+buTMW1qp5FnnNeoomjCqhJjcRoDgg/Nf
8zjKuWpC0PKH0jFb2ScW5BzuQnc+cBKyy388QTcgRiBLCwa/McccXrbPq69y
7ZyVL1K8aGFnp1A7Blt8miS/UDqD2pcjrNVDRgRvLDIpXFrRk3uCnqbKxT6T
8ridzuHibepfCJ1i2MzCC2AzfBIopPV0xJPCp6IEZezHeRkM2PFuH6OjaeGY
ZGUZEEe2Df2PHF8Vrrvk5CSs25J6RnMaPMnEnhowYgtlJ4tOAk8Mmx2u+vFB
3R4rzvZClhVmybGm73jcTkLNNculzv0xGChe+C9Fo2jAOxYsR2RkmU68v5v4
061tg7SKV6IUulFvkQ1Xv3tg836tRpic8TqEMpKKhh/uljVdWiRmwbf0A8sz
H3jt0iW2ZylFCDfi+AyW/kn+7p6qzlpcZCeFeosbh5mAU3TG7mxIq6avduAa
VVNzIgZUO/sE1/V2tZN2HVVXr0CJagUKGjwFwBkG+UDTbTrRBEPTnzuMzsHm
EVy26pHP8l3l98Ty0fRiYDfdI5Wq9duKbmafJ/8ebTjvVq1SEcL2DQy2CAS+
Mi+Iw2LY7VA61Fse67eoKNUfaRS8Oo9Al9/OLsZ3jUoJMCioF70HcREy0cVv
ADZqV4gfZTVEhUG4PN1sgHtqPd/rXTBdOls3BMNI74Jo1Qev2Cr18YedVEUQ
BPw3MeHlhAFtZwOnBb+QJUkTiqMx4z5pDEDTMzkCUawdrHenFdosxp3olhDt
G3n0iEV6oWl18ui7C8gxApSwRimlE2r1P66wDNCxMcjdFir9oKRkB8zFA48J
11bBUCbAIbnP5WLjRrTzgCJgv8zjdgq7ENbAmz8f6aFu2SE6VwvVq9L2FSKM
UI/1Xx0pWE/wEbbNDOp4oOcEYWUB5umKXU/04ttD28J9q6vbzps36mabblz1
Ck7H2Hj1fNDj1cTtLTSR7f4k92xtqPP/UsISbeUzt9u0qCxwHMvIm8uHYUR+
ztIGWeQeoJ6j9PmmqOfFf03L9chU6q7mSJeXtqcpiBQkosBBwp/mxHBu6A6/
HQaiv7mSstEXHcsyq7BfrgeMJzdzCDlfovuz/XbSfj8RswN7ynI133TY+yr0
DQKMsorS+ItfsmxV6jYTqNfzs2BwmD+uwVaxowZrlY84mP/n9v1CHra3gHc4
ujdoukRzfQUbrACFJ9X2KcVQD46zFQYcVMxEd66w3vaTA8O0kQN3QBeiVBMt
J7/z4njzR44T/7/ZA/Y5RzOLvdtC1jMz2DgCBYqLct7jhMkC7V4BrKkRDG+E
JsV4QaUL9Xp3O+vAprBP5m6QwklLvCd59lwhqWfv/m0h7M820vtSuhnbX7Tp
6wwAtGc2w4RhzdODtcPWFy8dSP05V+r31ZbAXFqkReczaIwCrX5kGynJ54i/
NZcEXrGBSXwqg9JBf0mXZLDZY87cT8rNMwS4+Dx1WildnPOZTxal3W0Tri0e
7OLq3HFeAQYWEwGGEMP7xAvfn7eb5a9op/RFsjrGFllcAGe0ibfGm6hixwu1
vRlxsyn+j9WkFiOapamt3YjHcgSpoT5Nsbtwbw0aC6X++ORC/6VIYuDu7xhA
kmYjlpHieZHEdel9HKUgkKDbWedNnUIJPLo1S/pa7/74Cp+r/mgG0lhtcLRi
QcUhnRP9Ro4lPr305439l1IO6hiqRVmmLGE9Q8Q4giMngzEIILSy32YYvOrC
TMjnPpvVdLHK2MoGxEkBstFOUhnWCFCEUMAX9uSuobuk7vJ3GWnrSb7VfkDD
SNXlTN9DRJjg+SI+nryojFLxEQBirwr+HThRlD7D+gdBLlQl+zXwF+zhkEtn
kbkFEkvs4T6vgE8dcapFXYR19b5h14WKLjIWpTstEgN+nt9hZhvbT/Ni9oZB
i4SY5ByOM8+K5qBe3gTKMkz4lYpkx/3KRhg2N9Jv4fsG996Z2hhFElG9bj9O
XaE+gIioljyGK6TxpWDjh5Atv0gpfetFmpO7KZ4N8zYCG+NFuacG0N6ZL6IE
TEMgXvdoiBP/VWRPOpMv5ySu2nzwyYWhmwyJFiqfv03iFJG/qdlToGQavJPB
VO7q5biKsHbo0KkWiiWv89zwuOTZqzNOYPuzQWkblDf2XMrjyAcGs7r8OnNQ
c6D3gSl2arUAJX7gnppHWyblZxB7LZFlQrAaOojtJLLTGOwua5KGSltFrjjq
tZMbgLYpBb0kgQ4BDNPzp67wtXpm/0t6Pe93gwAycPqt0Rx8Wri1PRFHOiMR
6hyzX6e07SoTgSEIam7tpJFbtiA3nLCUIhVGYpWbK3K2YOpgPayFw4CfjZaH
WEAINMrDYM6nm9Jolpii97z6GHyf/flWK2DpgnQ8giXwnRHryCuHrFEoD2GP
BRmtMg3RvHciWyLmYfQqHZqpa4wtoJ2SX2pvYliAxADMzb3GHX2MdURflOUT
eqmfodlPowww99hutw67zcVXvyH+5JZocZnV+s//o4CRNSCr8d07WWnMDBzE
0x9AebJktgl2gE55T/XW/od7br4JchNrR4OpQ3MpYHU25YG6nXblC5GHaGIM
F0E0b0M0sQkJx6MGXdIfIl87SFUuhUglYyovcuEbA3f7dgNgLMe4nqfmqWrc
YBScPTHvRlUYi4G0TqY5aXhFLPDAuP2xBO8NepK79iSL356ybj8l4M4mVzzu
Y1d9Iu2rhTicmZ3Y43vt8VRyNPVyH5DtRcDLZPhLREPzTyIPzIblbqNmqBSA
BgbhLzQKkhgOxLouxTbxZiC2HA1t9yFYaNqmCLZNPAA4Jems5BE+Cw1xSuIh
WjYD+g7TQ8VPxp8vxHaHRc1I7UHfos7YxDOF4Gl1EgOuC0tVMH0q/SMAMhbc
yCV8b3mLVWFGn9WM0BClTOedM0GALVhODM66RCEDoEhJ2bMcFs1z2z7gNkTB
JQeWpI6kI2fLVKuWzoWMX3ax7SVfqUJAgRudYnrmTkhVLsnT+H/6ebgEXgBw
NVb2C9jwqH4JAloKaG1BoQRNyOSLPuRqEB2xeDUDrT3qIXSI6HHl/pfi1hH4
SEZQhfNMeV+qSXnS+niXYK+2ArMvSQVlaOUAhNEDZh2x/tci3ZJx83XrGWE1
MA8TiEAs3V3rB9pzb+mSXZF/OJOa24RKBIEw+q3kPn/82lewa5pEIFOJl0Qc
mFPq8GoNWKdFRwmsSXp5VB4P+9caah2OIwhAiJbhWcA2kKwg2jxNqs8c96Dc
32hSva2HXz4/YQzjG2bgtV1w3v5hFNl84wkvMw4pDE/tBXteQO1C4vTQg5An
hLwUZ43mpmi0O8lXmczGv+zo+TrtTGavir+e723uY3jW24yoJv6+uAOFHN0k
8rVaerRD0Adj8GKskXxH3pvC6OPkXGTVhyEsgzQzzMaaeX0eaKuugAKd2wCM
RAdmATAT85z9i4RGzWUjBeA9dKnHz9ZkVqt5DGhCyBJ32fWgMkss2Y4Cvzjn
jnv0w+qCD2tYWRYd2QIM91ivdUFmSaNoWWUqsWki5YTqGwAp72xCRXn/U+H1
3eVQat8Cfgj4j33ZCLXJV1z99GMjRHsctRPZ7ciU++Zo59fSZERDf1MKZRA7
XEJFUUUlDUh7FGDAaA+fzX/jIKMsPVGjmG2Onq24iAd85EMaQiDBN+/yjXux
udJh+QqRHWs3hmBv43gFTC/eRa68f/HnznDNiuAFeknme6/qxC5aZlJY6qwF
N0A7mpS05Im6YTkqB4vjeRKFCaItu+ux/CVRIiRHg7h/97XH5MhgBBzW16O/
vD/jZklKFAZP9Nh1th2ga7vhdAtN7OOyVcqYYkf95ih1GPh6/0k+CDZLnj1/
2+VWlUiDwZMy5nxUDXFWId2XA7z1e0tVLAouJ9TG4zUaJqYbZTpktqODqwfW
uN3irOjkFdjcfEbBtieZd6XxOdDihMCKoaeJz7jApMH4T6t6ASgT4T8JV6O0
5Qy7U8YcLOuUwDYGGjxQKrJE6NMWLSzhD8Hr5srjObDXH9uisG1QWELTwf5d
PpAnjIlPEyPNw1I3ReqrQJZ3fjjfpQidg1Geb4lPIUI8G5yw7o77UCLKN931
vTm2tmCGLh7GZvKmEVp9ZF5qCX0XRM768Qc016XIfAf8ZbrE39J05vO7NtEy
udH/DuO/og6nlnan3tfvZFt4iGJqkl9g0YN3pOKRYpZe7VApSqcBvaTI2A5C
nC+qQr6HshF6SQ3uXGjqu1RqbXU2/pVUaBaJa4IC/Kib92k7UXB8k7i0Ks/v
amiAjbpvg17mhQQrfDQ76KXq99uaJFZSRclosYkWxW0hjNDZb/PVTUbdxQ4Z
H5oZ+0yNGBlJlcHUcP1+vVa2arrodDdSLMI4optAZwMCatYDQZW8AHr/QmMN
ySlc3uxnSeFjpKHZbGYY1Ibuz44JPu9zbQPOpBPdQQQ8FfggtVpYKIHJgcRb
0TbSlrvguifTMZOFiEGXxM1iufRIQudfahF+XYGxa+E0CuU/0hwBCKdkS+VK
oqtROOA7Dq3301mW/2s/gTqtH10LQl0NMSLs/jOdHI2puBhcc9t9Urrs5ydN
SThzwp0AfFyAhfd5YWVcV6oMREfqg3XWXB/klyzwud7PWGQJ2yUt6FW7BDTc
KaORcoaFydI8tRDVS4OfHL+/UheWBBMMsh6aK5k7xAXZ/LKDRw8Isal2zKio
i116ZnXEPa4gVcWXtELFzQmATUELG4XGCWbXmUg8GDe7wM6OblOOm8pB8gh8
qG4tNBHl8HD98z2Tb532plEO7Qc/ZlyXthmDzTXP/ORakumLztY4p8Cr0chM
twGuWXLyFqxioUMgqZh7aQkQbO27ojI6iOupebhY1NZfOWYLt0pEzoJwHV5k
JbDbdibEnu6T5e6fWy3uOx6Vtf72SuvRH5WCABGB0ZuYOHX1PtuRSNAiUfPQ
nG7bKJhGv8ahPp8FQlT/NNwqjNdcXevq67/UouLHoHgpicnnTdHjo1j7jRuf
t2Z7p9ePurLm7gpea1HgOcMxfL5mbYPq5jxbuYYjwTd8XVYbjR+k4d+sE9yQ
vUhf+LODI+wI/+i+Ci2d0XsprF+O/4Pbo4eEgB1NUfLpgFEWcZaz+gYv5Lwb
cJ/WOjyvMc1604fwJrjpayiv1u6nQf2im6EaSTfEAIN7QzvHkpxX4dB+/Ke8
JgCOk0VPKKoK9EQui/qCmRgTrkuQ9KcZY26e/n3Y32l3lVFzOVMd7qKKwmk1
bJE2ggbJZNlxb67aI8+ZFWQxRI4EmRQnD8aFBsBSQfS2CFkAghmcqb/7wetn
mzEh5tEhmnLIFy1Xi5TDEVHzRPnEZbHC9G6WdAe9wKRR+DWS21VH3YI4UO40
bkiaeJwWd99gRnfSMw0tIeINF5slVAkW5K7/Av9e+GVdvM0mVbQ9wyYhsSzz
+5knWyNpH3INtJM477VR+mjwrDYx+82/rEQv14wBslp5Q1q0A9W3nM0X2vCK
jNKWITSGJr7ASqEmPQgUDpxWYSbywQSUkeMnVuWbk7n7WFv/7xFTjrRj6keM
ESLJlvwhkMLhMtEZzy7JdXLS2OdDJRpfuLstFDIBMGeopWYqoIYDHP6aJLkn
GRpoNI1we3SzC8b2OgcvVFysNAW/id7yASaIYsZA6OcAkxrjoTwTA2XV3gUB
JW04wvcUAXiLIsaAvxEOrb0/LubZYP54ALc6cvJ1OXGuw55qbErZQmfzgiPM
0poI78+cZAVNhpFUdr391eSihRcAbBqqoYEUYfs9aLMh3S4nDzYOpGi+sjW2
2qhMFZ2cNsMWM2PsZ1bl/zrUSnwz/BEsEAslkKveXjiMraYsu2il72bbGad/
XSodMJl/gKmTGlbiIh2w8KVmPkyXAavg90zYtuintyyE8b3cq3QyU4gq9jB3
yisBFs0gjAqBdjVRm0yAynMQHpIg6AXHwU3FPyp6g3F060eosWe9VHyPej98
osSpRkBYgdU3R2gEpWVwC+R3idR6eqPujJTN7rIXAjVuatFJM6YKablszPHV
kmTWFnGpBLc6HFVbeGFOpjnbLyd/8eiV6ogGANOVPeIMPHOZoJJA7qMkurck
BYO5r8v1+pNqhvo3BNgFkOKioyJ3ioL4xCUf1aKk9MveyvNLBXwXAZDUCSZO
htgVrVg9L8rKAVD0EEQI9h5fY9Qse1JMpVAakpL8kUJUWd/xmP0H/S8dHswv
b5wLijlBjVPJ5746LKQa0roI3Hx2eHv2oWqZL8s+gGIf+JRr4jyM1/xIxLYc
45nMGdK5ACXVJo9CUUiJSNJx914kqmBmegrqp8RaRvVLtbK8sHjsxrWMWKwW
TWuu2Y1hHrWH691iMbCj9Z0LJuyV8J7dnjk5YjY+DS4UawNrIBA0V0c0RRVz
Hphn1wuiN1UqH8ZHtpd3dBBR6TnyioKYBQsvrzPYNJGFClbJNsB7z2sZDBfo
REkYIrbzv3XQf+RZBocsZA/b+tjrotYe8WRxv7ox7h2U4qMDw2sqAoVrDmNg
dWkAIQoJSMNBJmCbZctlP70P3BffFbo295VAgYb+XJ6Zn9er5ykAWGVZKaPn
uSBwdgt1fYgqo1vyA00law3Agu1+4CUa8ZWS2oBQButrzmyWyQL/VRNgrkxJ
EqBTZcVsldyqlXFC+/bVVDbfgoUXuCkizcXZMH/2ED6mJsKHix8Lk1K73Rn2
uKX53AjfVPb+O9rW/dESabmInc4DRgSduzl8ahVCDblE4lE29af7u3a3Qnjm
URaq3CjP79+oIPeAqkfvusRIQrWe5jdht4NxHFfgWuXwJ03Bb/o6t6LGGcKv
lrwjc5/HrM6SYXoo0UvzpOj/pbSSP9nZ6VDEYk5XxWYXU0wFbAIgCUAtQfwp
QIhR5sC2QdNrkm9nnNI4hK97VznJ3113KsGYGyEbeyMij9tjNPsLp/GeQXx9
nqHSLvpp6uKihaqiqWdtpmfRc4fMM0GKAt03WFC98WZbvnFxLBa5o9J/7dPF
yQZPJBpcD3Eto4VUv0SGzw9aBr58kfmQBiS7UGQrmvjujQHfKAQlGJ39vmEy
hy7XEpmiwdXPUWZGawVzJbXfSTfGiN7j2QFx4BWKqnDIFW0LNlD3/f9icQYp
r9ra+LWUhTmuYZZ6iZIlTVT6PMMWYG4hRTn36RWgXqO9gf4TG0tgRNUYyHWS
fzR4BFlH4eqhcazu+KTZ1MIFTrqBuJ8C0Nh8Cwin+wl8us1tZAo6luIneYYD
vQphDxB01BmVI6wW7Te3c6nBYXfvQx1S/0vVuZzWKQOAhN5HBIu5zk3OwuQI
Fn8itulf0q7hBCDgiIupFh5UPyhZbXAjS8WAlt1ri4sFgbfO+s54eEBP3ER3
lewWj4kdcG/tkGNYp+3gs+UPhsTsAh4A6gnKsWxLXhCzNbwbRGRuBBTCsq2p
9sBwPQaF7QeEzOJ1mbh714ABTTMMRCNH3pFf2mhHdYM23sx7xUfzF0oQGSa0
thLMWVfpk9V/XhWQ2hAFFdT/P0owk0pdk3tQdylF8TlombFId7Bapk1nwQuQ
0tVZGOBVoKGZ17Fz+t3+3skBVxPRES2dZkoQOC0XVuL2640q8S5EMTBQNTXG
7maQpaZGAYFD+FRPFwmYzZg3S7Q5gpqt0kkox6zN+Uko+DrxWrTC8omyOqQW
brOoQ86ny0eXuNgn3zvbD5e8LrddOZnRoJ6a2VCgFBd16lFC2BV6+h5UApuK
MNAzWXlV/XoLU4915QakhwQA1+g6ADwbaevEzv4j8Wby0r7P57zECfCZUi3v
neU1rJy8nDuzBRiDkK5gGTd9Bl+iNpSJhYcPB2A8GkeTspXzM1oE0IajX4BD
GW0feawxNHWR31Mq/ifkiilILR6PlTQdTY3M8v3nX1M2aoiG52CXtQDi4DFb
liQmO1bjLXX+R+sG4DOEThYwqYIa0VknLbsftlvesEvJdeT1bfVSA1gY1DYy
68Qt3R1e6iY64wV1CsEG0vbzhlzTVpRDd0XXiYitp+yu/SHk/fxOhETuppZK
DAVAh45oVfKy+LVx8Cwwf2UcvrVvZZcLlylkMrc3PITg5KJ1e6Bj71aTs3+i
npZpQNJWCsXPjDLAH8h0Q91nRkzrB7thezJq2+EDeryj1yfN72l5Cl7YWA+t
octZktF8T77lNO3wdvGo6NfNF/eLs/OPRtS+QyAbGUg65ObEzrmRy0Z1UW4F
mapP3O3OemEwgIw03YPtdMUpWmLZYkaZuxQJwMa6S+ClPt19mVbZM4sNlpVK
mbx+8Y63IfkOX7dO3+lhVJ0gPwGL7eWdvl0XZCl0l9pX3a1E6Q+2oFMN1f2x
Xw94VODYdHZOzG9VE/YpKR+smrvzLXO3I5LjCAVc6D7vK94S6Wkz5K4buymm
E2DRC41B813BDvvT53q64ll7NMq9q5/2yQsTgi3bxMaLIoJ/Pz+hMAaHNu0s
c6qsmDFBy3/sYX2P7UTAMEqIZBmFUp54TQHeIigILmk6xh4WSFTkfLqCMYUb
bgJZNQ56RUBNADADpVG9Jvf5UBXo2YayRNdM7NzGsvkWSmKX8tQxGPk9l//K
r6NnRHg1e+MDwLcjSEHY8vWHaDJZ734/3cO7oDNCdtz6VCfk9qizfAL714Xx
be80nCOya1Pe6T8NGwlrBrrl3Zxe1+XtIupkbajd4lRFXZS8ahxZaIu4xkUh
B0C3jvgraPlaSt6Ab/V0U1ZIlMcUk87ZtqhlQA1jMpbjCEA/MnaT4wIFIfqD
1Jzd0ZKsqr567LnlrMB59DQhaStM2AWj35O2hCFL7V1EGSgPqyPYMOIyGcVM
gmVCLRGjVeeNp437LVMR4LsTFSP+Rj2G4ZiDgmPCuYWejHblfg082XObsc6A
qHe5v+zqt16DRrL7HXtQD8j4byNLlzp3m8OzEoUC1Rhn9YYe+OsrsZyidcZn
pCtHU00wDxap5dBW6YB0JzbdHzOj1lFduysg4awyzBifBBjAOIJOeY4oqzm+
Zs5eFK0X7R6Mw14sioOJubEasLGjpT6ERDsPqFVXMOjFrLpi8MbY1SPNHQ/q
WGnTXSv22k7y6QC3jGB7oVe1Foyz8QhHkA5x33oDlRhx4Nazx7hDC7EnjHED
hXASPZ8ylQ5hQyOOjySb7v69eWNbEPGgxaWec1HSLNnJvITEUCcy0W7/gV6e
9jxY7H8428Uu4d4T2+AiWh58g297E3pouP/0Ynzoo1OWUwlf2DOXazvaLHSC
ziFmuGYcXZKLbXgnZDgL4N7D3DEeGS4XhLgX5vE/kY7b861dJ7s2uMr8UMMR
07rk6bS1LyxhQjmQMeZdaIyIAJDoFQFWAPvNEVM0mPOOLEjicL6t+6er30L0
FSFHD4jDqjIQkThey7LWi8459drxyvz5Mb7N4jtS1JZ2ZC+GpP6Y+bPUnSTN
tuj4K//TZqx/ihN1gBppoOBKmm4uMhVpVyUA0b3wJrpwPFROwYjmRHb4AdRy
K2bkNaL8MzNdpirL+BSdYBICpiIuqg/u7jwrOUc0ALry4IpdXqEYTJSWVFss
cdqTf6fyT8FUeiGwbnj2pwmTMFhVHS94PBbIobjknNVyFcMAo0PJpBLQ1rBi
+sONVTh3+Lvm5fk055v3luknXHvCfsImU22/ivnVCP/TBHDdZhNSvkPddZn4
c1kKvukgwED/4rM3e7wEaZ7TTORsTT0A+WNLA/XkNFpSeh4ljAkv5VtPyy9q
kd5vHYel5nyKmgSWH3EjHihaZG6r9VDeMs/odwH1Ykw++BgvP1q7vlG73Q/h
/u6dqWO5PRwuxkD7+fBvgRmtJKNuIYgayb76D0bQMY27Mnu6d2wjjGOAZpFr
S/1R/ErTVZxMfbUtvTdhtp5+ATmRSwpFdJNh8KcIrLyY6Bvbg5VvFBF8pm54
QY2Zlga8QSbIrMAoWG5908IcEXuN9bkY642RJd5wMVEy/am0d05v7/sGtSjj
GmsjuF5e8Yqu6mMSqF6DcR0BQnXX0gI+ccsHzlGmNQ6Tws2LB9t+szLkHPyC
TT5IxFcorw9Py3jGwV6NBM+FTy04D1TA+BAYJRq0QUTjqHAMqxa6NdCXspok
Q/rWObYeM7ti/Vq5rgtT+E14CGbol0qJxHdb7QlpTtwQPoHlA2ak/EQF/wVj
R7MbbLWagZ0bJFSE38FmXSk5Qwww6IHrIVeQfcjq/9a8lkTAdSKMbuLcpsjv
v47s9/mkoL8YnY2wyvx2Xn3f4Fqht2Uti6bIKxNIxYIY8U/NF7J3Ur2DgzHB
2oBW1tqB939sGcJLGyV6Zjjykz6M23UI3/Lf3ym9oDNZHia2uK5cKTFPR9Kp
+mAhXNNbsAyeHlCjUElGc2M02gHPVJRUhVseoKzkkkCMEWyuV25NXYhwvJzZ
9fLxOcgw317A/2Z9lgtwBfHXQzox9CkV7zeFVRK1QJ2R9Ai5vyMjJ2DNKZX6
iAVerJZx9cnxWx4FbEXr8wU3h9n85VRPSkfdiWo11h6vHgkeYKnS7N0HQ5JN
Ttzd8bopkamijfFa4mETf4mrIKfRzeg6JOJ08Qfp/2lNFodWNDVKt0CBStUM
nzNuVEJwt6WGQzPcp6dnX0uigEXxmp56CG7EL+XXXQSNKKzm33QSiM0eEJUA
2+hZrPwOeSFgqoasbu50crSOujbeVQ3Otx/nMkdi3nDE1jxQTTsi8brwsN1H
jlAqsyFdo6L8PG8eSBmsspwiIiaAUOQA1ycfl634FZ4I7hW43UuFjDwynEro
MzK4IQAsTdUkc3N3K6904lCyEYSLNJ2bbF+wW8QoaAd9o/peqYo2Nl8GrMp3
I5Sq77LLP+sLATlhCHEtBTcYhYmFV8kHWgKoa4uB2zpvi54naKcnXrabrLZM
NBrfyTKR2ZbpsCaeyPL1rT98C4IhL7I9pB2utYNVqRUTLx7kzJRY0SA9Ozxr
xLqImlAR1MlEed18oOhjkuhJtErLjWJmaNylcLIoGrsmAWL6zKnN9TzhTnHk
2ZaRgWwJL2thwpNIi2OTkx1pDjOdr+smvKDgGFI05x+jj1MV3eAdluj6jGYv
99zOBNATPbEVh/ST5mohaT/RNXe2w9+eSlSlBptraZqDVWGl83yvw/0Vw4l7
8wxDdNmMej88Fp5t0xs8krIiaNoIFEhjOH0HTgNSg3vmbj4Zm03QtQryA3V5
6QGWVv6wwGKZHvMp09ApVj93pDEEksCXOufVDWuyibWPFPYmahklQLn6PGTG
AIwYG7rZ5ETnQ5ZiVonbpfLfFuWCgc6jVaVOyp1jHeya3knS72u5XbUYVeJs
OSSPUAVj8Xwj5W+ixEG5E9yROByDcYiyZw93SwWVYzfADKoUTpoD/mBcMEwI
Dn6YDlPEhslzFEwQp3kLc8wwOldgC190J+7y49Rtr07rPertEfXwZRI/NBZI
nTH5o/4jSjkN2ZVCAbGGjo5QtGAgPTd5TFOREk2t33M6dJ0lV4TyqIyiJFND
zJfllAWR8xkfgmCrkHzsihhf2y89v93/WPKKaDzzRDL/hxCSMUEObFSpEZEA
K6+os/cKR38PX2sRbl6gZOfar1gNR104ehsac1f4vmKmMv1rmlu57c+xlkNl
BhrAQzLyN+mela555C/MZihAOXM9+yCMjux42hHw434OPZEXGZvn9ffn1m42
OAPiW75QbLoQYkTSLleLxbzneJyThVm9BgJA1ZZXgzKoVcvqsR3sASDj/PZ8
Ud0zqP8g5RHUqe7jpDSFGN7aP+DJisp7m3azj/hUYJPyjkdOXrdXSU7sF6yb
M0MBezxEvKgW4ruzArm5iXF+Q6kLQLDL4edcMnH920Xly0ouuS8yzkIrMItM
MaPJBPvx8g9+F4S/j9+waX/PilvV6DjxIIIpwFJ3rJyamFuyp02m6AuNm53I
My1yOd8VZZuuubYF8td4GmCeQjFWBoYvRGxYlqCKs7xvwyMnjbjurcHuBA7W
hCwsFoazbQt5cmYMEvJQYpHgMRWiwJDrApXk2q0wzv0kpLZnMZi8AYmDkRbp
m6NuN/TXrK1GztsUPDdsZ26rL4gKz0277leEnkY4VN380d21mybSYZUFBcrJ
qCCgYSWIgLtjKBUBqoT0F2EjmeHJYDjq2nejxmJgIafiOL5Et4qHcGCaELc3
IqVERSWlsyiF3s1vhvplncgz+YmGg/UU/tMI0YTmQ2sJl32syUExZYxmHsB8
hIty8gb9JBX0/2MLk3mFXs+jqvYYjSE+QE1qnAmImt2KshNS2N6n1FA1kKXV
N1A0vVYueg/XaSUrcPb4fyzeRF0Vw+sMGutb3os2trqUsD6xAflC946C/hSQ
e1STVBvxzCnrZhJ2vxeygEu9zZDCe5jrZtILcQkX788TupFyuVlTxAaKGXKk
u4rQjKGqp7ZaiHXGuZRooCBh3NHRe0Y9MsDlWZo+L7UmPlMPY/JQNm1lhKHq
qrdgeV8XR8/QJvfqlTP0PX+5DirNjgkWk2C1qev2KCgveAXBjfYjUxVaheMU
hBkfh3ZYWDZzLiWZlA/P5TVWlM6eZmyPPXa/jWYE6izr7KKiFLkbOgTt44OQ
kxsv+y5I/a63sTny92SuvUeOS+WE7dbz3DxuvL9y21uxHws8PLvdkf7kt7Em
pN3zYLMgRoaleCzRRiV/AJzaaBdXHIvXewJFf7z6tRu/ekE/Cu5PDo5JA2Hh
B86mYD0W/dhyexacmMK2sAOyZi94+wyAAcCB3SFGEtjZqcya5o3ifZiNmmoA
4EB8tiqXmdaBIb8FZ2CEVd41D7XGNKA1W67YsZskutmZmkmyLKajTtJu2VPM
y/PcgLhC3uJpUuXoIBKlsaAdxy3ibHyHBiwCKKmil3J0sZCdmZ0iDcKPSYKx
41nJ+7cDDYz8GGh+EljSdVe/IIb8ZWATY1UAHFROxDNyNyz/jei2gBWAsotM
Ad1cHskFBDRA8nWXsbn2dcfWai0vbGBh7Gtc5DtMHnTlNZam33LXVS8VbiDI
NSpMYqmqgwDcLWK2WFIulouimkZyFmdIVjUBeI6oTJDQ4szokNIPAeWFxFb9
2TkeNvoD1QNOPxKhigDjmSXtT38478N5DeMYJqZ+al40KHL89+qUgxSKt+or
ToroW+5Gxj7VQQlAkTh5+u8AkVZzV4rsoBfcX2n9+uYx/5kAHL3LfeErtEBX
C0/CuhRDtTdSyVegXiZitjITEG6jA8D4I6pGiSUHQpGeOFaimrJEIAIRFsJZ
WqHQUUpl9Xe1vkyVsGORuGSYO+8L8lZlrCAdq8Cav/aWK6m62Kq8zQkX7qHg
5wB3IfQQKzDdJ8TOFPQinrNClWzs/igW8j1Nn109/zVetLB4/ReIxOwvUJvc
L7rSVsfXWbR4ntmj0avmakeauQEa8pZS3/kDI14jHqsNjQagm3X98+6gAGE8
uHi6/5ufW5rP9dJWxnEFaJGdc9X/7AnP76AwxbJr7QHEFlZo7aFnpOILrc65
r1kigaEmMK3i+/d3arCGLWnUCCLFAcvi1qPYqrO4PtqJWSbyZn15/kiZ67gU
+7OFSDsdmj4GY7cyI2QndBUFEKzfY87mbFJaVnZCu7OS4tAT0Z8AVq0+TfiD
kS0/WTQ8l0rwkfi06aKtUOXDecKy0lAiYo2U5o29rh0BdKpbKGpljcWkZesm
QwaWepyF7mdspe/K7OxYrIdy6MtuFb7ZvS9b+XBjb8ewwMcXzjkoYjLWkrrn
9luRORJLKJQUnOspUcXw/I3/KBMVn+ns64XrJSEO87qxDIRW5a6wZljzeyNZ
Ym0joELCi0j4QpXXyTp3v4IQkjqc3vrO1Z4+Pa4Qb3X5NVizuzE5UBU+2Zdc
nzJySjiEXRN8I8lFSGOdMrQhR7ngor6it4FLjOSLkrYMIfHlPYr0HbQrmpLu
/akAS2aM5AprUhWsvmqeznuPEJgsEB/GCuUXz92Y61JsZ4WCgHDlcv5mXXi+
a29eVYf+3gwtyfo6oGCWwrAwRHc15CmWig+y40TuTbP+dBKj8dVqoViyNYf/
n84Ax8uzLkjXF6niYrrfsh3kZzBZQ67nspoaiVN389oqVTyeOvkavFz+GNb8
vbaoIVyMOcaYfepRxPEgBelOBzuNNWnrUhSiIeZ0GGRQNLSrXAaGk8RiBIrQ
8hLqPKBN3ub914mESMZzKT+Y0Ig4r4i3UJWMdumrwNNH9AcusoWyMJmqMDZ6
SDgVr7nBcaOhciKVh/Xiu9ZV4cFl4Qk7s72J8z5gYXuPLUgH8zaQ3I+36c0h
SyoSd0NVI2ZJcQwhIJjtXwQV7US+kKWirSfufOSWye5SqbFGhGr2xeJIkhhS
OwwkssmnSdVqv1iego/nmiW+nNaOBvwSTPA3MuwBt59jxEPK2Ns/s+NRIDD3
RZtIFE1SQKUpw8JEMtQlpXpR7gNNsRlF174SClvAhDsyqvUk+FvJU2Lzs8ze
JPEhthTvqAhwofBtPHDCQEFeLthgHuX/EUGPPWUoTAN8emtZHPqHzOH7HlsT
63BP+frTmHD4ynA0YutykdswBzkpLFxRhn75lZa+YxNUZOg1C04dTr/sNKTc
P/tmILHvFK9rtZr72MWBp74MWvJ3Ibxuk+hnAZjEnv0fraESUYNz1mzAbX7a
goQebkPtCQVjUkamPdBgb/ZHmAwZOEdXCsaDcuTTGyP/WjPr1tW3Pxx8CANg
sb77XNXiWp9OsSxDfYnB+rxT4/qtBVTyWl3IIt1VUkXMcF5JecEZIu4mm1Ol
hG+lIXkr8LBJhcsY1NqE1xnZV04eOGLOfuzXJASIF7HNA4DxfFzmJMcXuJGR
o+2SIdO2iFZq7Lxg91TuK52ehqnyI0EYbiCkAor/BO2MrkkQffHFoov7tHJP
14ZZIcoo68QN7yVrQ9zl0IkNd1Dn/FP2MIiIdv/C/QMeWXw2RaTi73lR8Idk
lbBhITSVyYqpg8E0LN+h06HGDcXey5wKl4fl6aZEzrlkP86Fs73lV9I37fqb
uD9Ggdi2H3qLtnRY60ja814vDndeKbg2QaXrEIAfXPifdwEgGP1g6Fr8FOa2
537LI+KlIbxF3t/YzJIADOqeoLiFS5SOoxAcL4r8jszY2fYTjyBvWH0XBYFL
wU0jRZUkWsbxl/92pYqf9ZWDFSrK/uap1BxCMtdN2pQVfKENRFAY4MEo+lE1
BgM9Sw4bgwL5WZBLEuS/P0hupGq5QK1Ku0DwGPqZ1RB1c/TpDzi+jVx0LlOw
Qo+Yx2yznHv1tTVAmNpQ4VlT3INzqrbAP+MPQ/cJUUHYbfeZDefZR8O6fxPJ
VTE1MkfMO5ilrJ4akbyQpU9J5tYQlOU52/JqhWnGse/RFVYk8/Xa6MWwjqUz
dBZXEeM+TSuejzj72s1yVF1fIxSGvraQjukVCYu09XwOP2k+EOjMhoeB15nI
SBvLyw2pBCzl8OE7cVTkZGTiy7eMhquL+OdUiFb+vLiRo42QknkjItZvpNDS
SJQ1qil8rwPPKKCGbKyvaB7gEcDbadBYImSi5tvoHIV8E0GXOwJh+SmVsFY7
CpKbci0L6D862FxaP8RtKg5V7VwZ+NkKNW0veSygMEw2EMBocZO7REJurZI2
rDyY9WTsji0FQqkbFxmZ5LBBnVPtZRzpO+UL5mru1iV6IPoCRI1gJpsnfHxo
Hg8XEd0txI8bwcF9Zw+VF6LM/Mdf0aHdIEzlKGCvogxDwcVATk5YBnISvCjS
S2j3QhE/UhdhaTcRfncLfTI7fsXCAkFHTuWRrtvHEvYgFTd6kWJb71gVmM3B
Synr4OyHJvCfYa1Y8BWWnDBqhHzbHU4crWjjz8mFrP6F+DdVkfftMQE/Msm5
IY9+LMplnkOaOrgNKa7mtpP60nyJyTDQXDCezXkldWmC71tPmlm+O63weF+2
Tw4ooks3tovEIuAgmQsdZ1RUOO8UM967TYRpULB+TsHGq1h3SwGTgqnJn1HH
J8ceUtuhqdSvYVEu+DyHlhFJxjiJ3pPkdLo9Jpw96hPjCS07sy14Z6b13POg
bB8iiDA545xrL6/lEnCMHxkfv5pMsszEN9hAeGK30TVkSbZeRh1p5qlmycof
HsUcAihPEf2oWpUdC5HMaBz+ysLmhZUnp31UGKw4L/ZUsMkvcuD5fwcvaIO6
yDG3hLFglCLB19V4d9FtzOdcWKml29xbVB9GcBaGBi5g70WFFNWSbSjJSw+l
ZhFXphwEec2ItGtWqVFQwLAonEex6pxg9AjcbO5T5KI+QDcnh/ecuuJn7xtU
zc4V0R5+rJnbWZjXFXTI6Sda6311cnb42vLqIDdtKfv4ZZ96r4k+L2iHTsfG
Voir2JMCur7ZVBC6ygvoClVmRVJidv7B36p7gSjN0U3Es88JEXWd2wQdSV6K
R6jNWq5wWaAVl0WxILPDvh/uy2PcptEV+anxI6bucgAWl7butobl51wb4SgV
RVzdw1+idsApBbDghCkumbdkpesEpOFCKuKNu9bspTGWdHM5j6wTzYCC6Twj
837VdFyN6li8x8PJmMnK+VHPyPz4dR8kb9LFARXQ46bORriQtxhMQcE95xVH
f253hJx6E0xkEKGHPPrhmK/vKAfDPSVF+iqA1wy/WQV/ELinuvq5+d6h4+xU
y36LH18g+WpEOEy/Qd8IrZ+bJFYzmfhxLjAMqnyCNPzlWBm0DKhqns/Bsqov
Vcw8rHlq+rSt3uOuX/71d4ycisGiL896W4piv1jVc+PsyswtE9L9JP8EjITS
Dzxk2nskhgGCCUrosiD5v0uKXQzv1UAQeOVG1qTSnjX/O0Tc/7Jja/VegV8k
aFspqtuiySVRtGgRZHxjDVBDqhrxDgxVjzzXoI5VSbQ2z2rZgTZJvh0ZOIH1
Xdze3GCkcx3dgRN7Xo4LPLPumG5FwS+upMlC0z1xYJDjcUvwKma5icRSetOz
DjjCqNBnLbyzQaVFL5MyugqZhkuk5zf894oEocPVUsT8KJDx8kNjWUK/Md8I
bJDh8qIN5Q/McbIXDRNIZU+T7ZI2mVqmppYGAgiFSEacNNJHSVf4mw+2syo+
QBc6vw3jymvE+1FdTrBorEgTP4xnID/TFxZtU2nZ+DjKwHKGA3HxJpkQUuka
bxwdZGSaxNehiiq/bU1EBkhftdkxG2F354p9KMPjO5Dn4ojWdefG0prT5BbA
a3v5dTXWUkJfZpXZzHEdCnHZgxCtj9eZdJ/5gfbD+fxNYTk1KPLmK12uDV6u
ZEpU1MWT5NPWiW4SXyVZNOci6jKruiv/mPGaRYusDUBssNdeaEcPDFzL3hvf
Swpole7jHoQBckBYFRqv+ap/exleWBij5UU1kWXUWRVaFi9umIhMCUT2Tx3M
nLClN++q1kaqkmu3ofmGSZxLPBhJywr+YmGTzyw5geNyfIzEERp8oZGOSmm6
7hGOcjn/cqwnku8lYWylv4u519V/yrJvVkwb2H3ZeJs424koFrDTiiF2Rpxv
GDeAhnvTxH2A3Ii+9SRTrkKtSUb+k6Z3lEb1Txk4YNJ2uDL+6gkNe+EyWa4a
KxexdPxnJuHFIUczHVMUgjNJzUjX1kRdWG3rCdKd11jdpo9c0xuGpmoSxPHk
s6m4C8JPaomHXL9MUfRPLb3xTwnnZDEqA+0NlT8q/67Pt0+ea39gZAQtNuJ3
DekXySrufkGk55dQFQrTMHDqktAh/v0XGy4YPxdA0q2+wPmUV52Zu4+pNmcv
DeeHxbTqltyvpAz1+XXpir6P4UnjehFQEqb+dhIVvQ3YiIiND6f8lMkU1niU
BPfM82CEJoOtcEhgWs9S9Z0VXNANkDvjjsch14NakrfUnxUWZ5QLbvV0hSmp
Rw3qlD4WyMd3/icZJGnmBs6Br2727NWz7rnWu8jEttUzA7shXLwBeQwF1wJU
ZbmjOuBuFEPLHI7/vPjiziTjSVe87hmCwi33ail1eC72UMPEc4j/Rt13ROfH
bWDzuDvRIYGLOWFYPpCllA6eSZsItyr5hFh+QRCB142azBzdRjQalTsTJbzC
3GVR7u7Lkv7zUS3XGPZuQbM0fIjjad0sZun4kzHKBQM/ad3fKE/UML9XnJuD
ElrKUKrwcJ03fodXSmthkQa90XwN5pE24rdwztSJ1zzRhgyyknMJsRfDX7A+
UlgcHn0bHidPzOzAGNeizj4xYfkX/M5qroYPJ2X9ixFoAzU46VdIyNPVlj9Q
o17QnPtwA+2+qMVgKAZGqZ9AQvWw9dayvU5VyG/M3fIp0aBbDD5zkh2JLHAQ
XAYMTB+jbcJyu9e0j/5gcfBuL0KsZhPv6ARNKz+xPlWzgsqXvtoCIS4AbxQd
6gLUA9fjVG7fA0OYfadSAmAdb+tGUqm/2a0Ovf1yI98i3enMk4NBW8NHa9H7
cLy+Gf/5Ik5OM8RKZjK1+Uo5RRg3GvMQc9XIcBqGkOwiEDrs4n0VFDISOXSj
kQ8cmuGZOOVXr/2Ae+dxXDidh2w0psfxL8lyQyECBblMbvJ337V1kAc4uXh3
+uTMC1s4Iim98KgUTuR9GkfSWVlhcL/3dYhow0vFZ9OtYWueasBBtTOfuLlt
oR1oR3kWT8l3KqVf4P9sK+wP5qOCaGFWKM9O/7+MTSZSJ7FpmY08mknS8JB6
+u9uk6oVIkVBcmw8o4lXHY+qdSgQeWj2+P9j1xFsv5r15Ih69JilqF8DyfvO
aFGhjfok3+7MWNT49y9WIKQvREPasjSgpZ+6dOjhbAUs9DZV2zMD4J9O14/g
iOYGpQCL3squMMbxnXqa+HiB5kYoMfPlgzbbiDee1dnsfumXlvtiwnY3jhKq
D3UQY9CV/v0yJKqrfmytpTPlYpgOg2OZpmDMSZr0G1dDycRL6elhZlxsXgES
+H6WLWI7FfK+So/bVNal0n1w3gKMddhb0++e8zsJkU7n16CUQAzxGc6hJu/H
HS2yoqz5PWINwP1nkURKpXGma+Q4jbAvfvIn5nraTHuX/+PcLxTTTdZyx+C9
y+cezlLfP44lXWmCoIDCorBJrNUI2F7ohhVFcQMKDkzvUvVgkwTPxh0SEOtL
O8xI2NQ3QGTP47ENSu+tht3syuZJK+bwNanNq1kSI1EqSrtyZtwlgQApf9QM
tMKqjmdu9oTI+IZeZmn2ihnxSZeJAFBj41gsCp4XJn4lYwuLZD57LAfUXUIL
twk9+IplNCgFQB3xeFPKJmIQWsuLTCsOZU7J+BV3RXDkHspzf2JQa4OLWlG7
c59JaVvQTF4wpAypKfMzrhhOqB57AeLTiyGwf973ZzgjcFWJ7F2MQenjoJIc
uJz0+Ddb212h3m3hyFgGKgbTPAPSUqmVY2k5XZAfPzDbDgyweWvvAOHBwDZA
iq/aktKRL6CEHcHpJpeY2xhNWcMbkQJocVa5ZLsx7Wk3c4X5qeXE8ESeBK77
xP770y9Y2fWqv81Gr0cVxZOe9nUdfTl8/OyoKpPko4NkNsctOzdq4mnK5bUQ
2F+A2n3LcCkrLE5xFF0dnc8/RqO8/p3QAuVlSgRq01rsWY+tq/nv8QO1PUkV
jMAQ+162aY1X5aMSzyRv9/eIh6LWsC0PM5OY3nDCdBLj1EpOSBW2yv+A3515
S2nUbAF5L4R/b2J41uIZgcHSF08ch6qHT9oEBzQ98S1p0CPJsS+0aHHVs4Rp
tSmRRpW5yGh9P7VfPQkcBFiFz3u2CD91xC14fw4JYTgQIi3AkqzzWCve5dn7
B6Uk2ajzWeSPp2RxQLkiWWN2nXbAVoRUY0uwK60NFVc++eu5BnuZkLXz9Cwd
proOr/7pBlUBARBPaioyFCIan6Dpv1JvjV3H+0yrNIQ5XaySjImVkNOlBgDF
SZCVEXLqYsqmza0fb2u5bRfcqvpLGUNcOCviHqRE8502eWS3dDRM1G46fXCL
JUkhBTdtGAqhwlkcD4QVTuFtxfVUtqdX1FBahJvloiGoKwDAGP+7VjLIgnXz
hBFlfx8yTDRbDCwtY9DFhcfDvL5p/8peMML42ZBjhtlm3a1IK8rD2bpcMC/b
O0TJ6qyHwVLZ+kuvgXoCjfXiRC6sGFtFwRIlKvJVPy9rnc0bRT20h3Osiznq
8SjLpaEkVOMVonJ7mXt2Vj1e1Udbx06B/XySmNRcJDK2WbaDzQiI9pERY+rb
jASOBkXmwCiW7yrDW1E18uSiU3unGbmP+T4qUKm6lwYz76Ww+EZUkPwVtXNl
3YOmSq0lIryX+uvDXvO/PYmUmS2uLfNCl4ZsmmbHrIK+G16HYd12mT50nw/j
lbTGFakqxpgCIFbEWQU/0Eic18BE52hpZBLW1CrJlWZwndP+ABek9lF8rmdb
1Qi7UHhr3u6hWhG4svbN56AtZJ4xwXV9smN/tEt9tDN+8lgRYaHVtK0HHkMb
w3FGdh/iRzAK5z5yK5cJkScv4SRGJsQF5YNzhIe2TWpopKjl0bA0KpW3hJ6f
rE8QNbMYS5VmFAc0smDPbwOVbJzX1f2HF2TmNzdd5KUzr5QwBjM7RKnRCTQu
ZAz3QWxcxWOuqs4xVpAMKc3JkZgRkFIjZZ9XfeeKYdl4SClQxGUiQwV/JYs4
0ftAVfkMunrISDSSl0uXuZwJTOchrR/oDFB1czBz9Yn35r9TSt1ngkYE/H/P
GR+8yC4SEPnUXWRFwVyo2C4GuSfauQnEWEGXCp9WNs0cXaOik2XHoRJJOFA/
wvVncdRnL5P6iDAMbrGdb2OkGVAJZwv1kTh1fJCnguAS998qePLGmyBPbQgG
i/+ymhOKydzmw8UmHmsWF9TTBlwoGkMSkifT3HyRawWrFghUA+pl2WVTs3fG
qd+MlGFFt6O3nDCNF6ydCmRpxhCFDjVMRWHI/9jypzUdrc4aVXxz91ktNoq+
5H/518WPmHbgqB9gkHkLkfOAbKjNt8bxxjA8OeuaD6m96CE4SAg+H5VA9i+8
Zah/csK0uEDv9u72fGRkM/034ItvdbYaJH+dTEZOQaf82plpPEN12KuyhhRq
6d2XSThp5QBgD3Xaiyb9vQZi8dYXIjdOUfhVR8Bmz4yc5DuS78yJHVJw//Zw
O+O1yDaMkh3aRKoQUkTq388Xn7H0LuAM6ejsmKr7lUYkI2ir22m3gKRcv4+b
+/h2gEBXq3peE/MYxty9xauPB4Ui0eCuk22DT8p2tD4prk8ib77Fun08uKpe
yAQaLE1ptkKFX9fIlLZdJK/pE9lZT+9nOV8gHpyB2wtBPeTnO6xbL3OqcOFT
NWEdsQEthIKQA4EV/iv+84p1ewa+faWp0kKSgDjbcJ/V7HaWIjwjITz2xi5b
CMZ3RALH1LG6ERNNMSQAF/EUIvKgVQDTDBgtDiokehK9DBmkrHlcijSIlya1
DwWhpqFCbF21UAGym1EQblE34TMIkZjax3Hl2K6W7qh6/RMet+puWyMaV6e/
SNle+lntFd+EPlL/CVja1PbYaUO8GvRAWtC0leRZxemmMzdxq39saM/Yozw/
nXLDew0jYgDg2sbtcgbz9cIdznDwig823mOuk8ptZEuDT5bxJDWsQ8lRGR8r
YyBIbiYgcEyaVZQxPCSmCUr3Al+JtiXb4i6xccfGmxH6K1F0J2SOIiepM+IB
hOyiP6Vp6WluXq6HIBU0VZ2tqJnNVTdYTjDnHmo8R5aYrULAE2n9W7HdCwgq
+WM+ucJ8y7F97prztLVaRE/5cdoy+smQBSx2PsgsOFsiPsgVKOMlkv5wZKGe
IsyRbG+a9Gga/Z41PdtOKQWT9NBeBehLUEtvoiJYN3EfmKoj10P7ZYtWj9es
Uz7Bi0nkP3K2qMcR46pPO2dez043ldE7wnfwwYkS89mgTm5xDgtozgpi7nMM
RmY2BCAt/xmldQVE91uvzRz3e64ZeNtKPSq9VIeA3ux0V6bUak/0b0HWQug6
WCmY3IqG1q8HXsJRB9v104kL6yWgFPLqb1qBsI0fp9ohz7/LnXid0UqfHFrk
m4DrfSGSOPenmiG8JUPVP1ArxDLSF0NgMiHJbPnabNSZsc+g/iYaIn4DiJLY
jglzfvC1zyMzMKIpc7Xo9pw1EXtaft2bmqhRheEDd7/3jQ/PbYOupUOyBX1Q
Gh17Q5UjJvRdN1rEFyl230m9Lf66vXGCVD73ngdQZlrGdK9WEF48tXsxWaNu
yy4slNlcMGOq5n8uIwX3ax2j4m6sFqihAj0e5rMVqfa079PSk5xqnCBDmOAB
YL6IgZVDBpe8oUCbtB6tIgDiLXuJBHC7fyYpyM9mghwEz/7+AIOm+s0B2IyX
ayi61zg4rH9nBgz8Ro7mPVegPi/PEQZId/pCoCuBsize8TbRPUI+xODL7PrA
qlZC51+EpaRTk5drloElOjudq3+y4nNSklqQ48gzaKHUxUh8F7m7VqMCnZuC
SdH2QHJKpdZO7bWH38jvmjxp9nIZC+jpIIL/Sn9ltCDKpd5uK5ndVzbCtDHP
3w5GiX80M56fAMJhvoeI+zSfzRV2hghBOEBC7/knlJIR0QTErwF5mwgPu82g
d8FrOd30BTdf5pv2VPr0AkG5KFn+xoy/fGJfP3coWRoYaMDZuRAYc3NEld5U
p4ANDkZRY9skewLX1drBJWTfRVKbuJBshmYuzUiYsvbyGOZVmTc3tx0SIdR+
ZP1p26671XlZZmsu4hCHr/fOnbVOVj2H9/WOna36Hfg3ALHqpxEzAogzrwG3
G7gXAAQwG4u7fJW8tgs89ykTYzTm0glw9/VCZZjrVAYj1IkcQUsii88lCwoe
Sb0fcSw2M6th+47wj7MfK0C9zebC2SOAQ8U6tTrqy2xjgIg23VOP8VzT/TNh
wQJpNo4yow1rlWfLjdnV1v4js1Pwqoo5wYrKhv7HDFDzzMrc7564AfLjoz/1
mWtCd9El54YsF9b02T0dxwR5FA+xctbyYJ2AiwAh7KJrlRbjcGhfb0kUCt5z
AFFWnyZV45O66spQkjjXIsvqzak5AAcPV/Bd1Vz0ZtHVOnHVOfqLXrKGQpbB
OtUKXdaP1y2VGcqnGHKF/yyYDNEx6r2fQlnBBN9Z5yEj3vEcwz2YvvLTilMu
FPq599f1F5rY2xbJrXrGw/B/FxR2tGNyKlX9jyUctqHnlAer/5WzUQMEknts
43iqKnd7QEcwZzTxKdAWhR6UsJ+HGlySoObYr0QD7GCOBcuCO5tQ1XRNwju6
JWNkx2v7KY1DyyFdnxklyaR2GFsvIZToN9xZT1K39u9HaBWXBraRVgqSF5px
k7Pj2VWb+gxO4ov8uYjcshpi9M5NVn9oJkJaG/o3gJx83GtILJpBn+cPYxMJ
FQgZ8Ct16ltMnVZzKtsnhy4fxRxx/l/0ylVn9ewK8FaxTZqWkHoVonjPKInJ
U64dcT9PINjN9VVto+YaAkG6h5HOkWNa5bKkTz36sjjT1A7tmV5IQAyvlwhq
3SeQSTilI07N/iF58BV6zJMfxHR0i+djX6trt5FXVMXvGMlWCdmaQH3hI4KO
YRa95A2HjbVVMSixse0RU4KoAGCfo3feIShsMzEiuaNqrhtwBtBNfavtAefo
GUSGxOnU0WRzWjigZ0pkRu/nzWyCWhww9R8mY1R8LyIOd0F5GZmUN7HvON5E
Z8RjC7U2MnYwxPRIL08fEl7qLOCJl7MRAdaZFC816gEu2dpzdXbZ47l4v6cZ
eQ8TnIeHM/CyI1SFfrRwoge7RXqljeXW64FL3fVqVozv54O+CsEM5D0j5FpS
KBUPxVwyhnTI+Y1xpuWAu9O+EDPUg7w5scragI6/uU7nvRMtoaUQtoXkRgW8
jY3W7z40QZ6tcGCI/s5PguKpeBtez4sBmHWF14uF9UyfZzjObg8aoahdLNZj
ymE8htmWpWvBpbCjq6mJPce9qYHPh8wSLS7enrYQAZ+tukkhsF8lHPV6u+YT
AMRogmoINon6bwIjIxH17uznOUlz/Kh38LEun26UGiBi1MVJa6dUzd7CET16
PJ7yx1Gx+YCUAgxN+zXaWuanIDXwwKLBItZvwbgFYerTTxGW6KAtJaR6Vywa
GNwwKgNko/9CfqO8WfGBE6yqx0LE8TvUpEHyFf/ZsRwc6ePyLeTyqqQq9KD9
P9NoWn4Fxaw/yjwOQw3onNrgClX/DrNYUVBl+Tgv/YwGjvDA/3tNjXLhs9Uy
Qj+8kwVY3fc98sHK9IVni1QTPY4u7nLckCgBMC6OrCxofy5KtBRmiots5cCk
q2Mnug9mm9Umm9unLs0zhlrDTQr6UWMmS6wTQIV8IK94xZFdq0xMU7ZMDASZ
eWwo0NPvVREhVjg4A1yBbiI7esbhUnxUJW15ZzyX5PXz9PvCnKyukvhhkn5Z
IuAIIcperrHRk1p+gcthDXuLly5mx5AVpaFds/rBPPBz/fJ2FBEh1U//DaTi
7oGuK1G7aJ6Efew8KPNzITkIBOPBv+eJze0vlLF3F3l3w3PJGhtOY1Aqzmvk
21yQ5bWmUbp/wORm1Ilm/P9waD2N9CSaQPmqeIol0tIKOkCkxOMGjsBY9rp0
jeKXHQaWEbcpzwVYHJAcwgUDQZYxN+X9m4+EqbPbyHqnWG7xzC9+o+7wfWbn
bsiq7n/nB/xqoUSo6Z6fXfOdXSoGItNdluWjM6mwYTsQmT1BtWQwtHJfP1tq
cVax1XrxyPR02C92+AFKabZ4fqXHywuhm6TOQ25Xhv75ZPjS/DexDRJhSKUP
Z+S+hK4zhj17igTlybFeb9Sld/2v2596pYqKS0FvnkWtInae/CtbD4Zn3ITS
nkJdtbjPpy3apqmmiTv8F09UjlrLt5wlepC1O6cdWHTmx85bYaU+bYY/SNnj
vJ6kwLZ4Do+he+vMbXUBIbwcPwF9ABaQFM5mbLfV3WZ+bebDctk0DeUvm9G6
OpAdRG63Y99yl0RbQ1YM/sGia6wgpMrazpUCM6/4hEx9K6pk399j30yOQyEJ
Ze8wDVEbA95GKBmpoanA3xRYWcyidWKL+koAzGEF5Ox4MMvpyrBXbKLqMcP8
Z9McIjnqOTRc6mkHS4OxmP9FXsEpOI6W5J8g8121tgLnOtO24R9wllv465Xc
EsbcJaq065Em55A8b1SuQh5GozmSgMboAeMe+blx5t+Ul3XsTPb+eXFWeINE
3jeueoEYPfTcnwGA0Ra7tiZbWcxq0iO5dFUwqGqKEjcFZBFdbYbuk+SA6wLQ
j0vE6R2JaxuZKqQbAj9RGJl9GdPXesvqP8bXZ4oPlgqFLOrzR/ePDRPJz0S3
8iPFUxFLi7JtyNda1PoZfPKpVVtJbyfFyAK2m5G0KI1AST/Ki935ID/Y7+64
CX7Ado3x1KIqOru7VlsauK0tEVf41JIvHea04i/WiJyfbJARZLclqHhBBvZy
OVv3o9nk1EQH27bkSxWD9QfORCNo5V5N0S56jqxHs9VWIQmxXMj2dPwxNeyx
1cKb/ffB3wzTbbRLRDkwoObPofUDjJcgrcU/wpiuD45k3ZEDlR4U8FwCLLHa
3NaqiUoiGO4UDQVTk/kBXIBxTKeh1vjQtLt1H701UT6zRWdaq8vGIg8uOgRi
tzNHwuyEZad53i8njkhiSgE/Sg9PDl10TDz/WqfAAMoDg/+f2gxtbJP+8zke
Em805aqkj05RBh7QdlBtpdKbMWn6i72JELqXNLSDLLtaePfESR2aPPoPQARX
CeaHdOn+nSj6heA3M5oIOw0U1BS3WFegrVo/LJ/whLxPm9riCAapJOxqhX51
2Z0VcTMJhsetdJZw2EedSWJfT33GzZ2zOvUyuK/NJMN1QejV+tjoaX9IxxIT
qgg4L/QmQ/7+GM/mCFkVMZkvhhGHUDktd0yKTGR1jYxSJRRMo8iJQcGJaP4e
HU7ABJl7/Cg4zTCXx7vR/09Gf2dGQX/o5VKP8HXfVK7mi7VRuQIkxfJ2Y8tj
QaNyeDPrY/RYebo9H7dttyOWc2P/OnEdBIWAytfxXzCO2nfOdsu09JJfx333
LR+6C9GjAh/aE2cHhyzVmFjhOUnQak8mmGiJEF1JftWFpIngD7Iak9HDlart
oRmVXVyD2Vt447rZLkNM0KfaYWmUclD2BIJQs1bzGKqZbkM9tgk5HLXdcsLc
VTARHXUMDwpwNv/tUWHe1sWQCCtbceFbKnbqdPfe32BVqTx2VfMPklnJfLvW
vuAY7krfW/4cQCij4cxINAkZuWze3unwKHNr8Fo60bBVzWhQ4n9edZO1JL+J
GPFBW0CIpyAH3oX44ergfhEhy3bl52S2+9oP7yZo8vjAWB2ZpRiLtgIyT59Y
CY6PHAc7ALYnQeEE83SZLpdxiAApXJtAO5Hcqm7oEJO1cN2sBkOcnjjRTnSv
TUod4paFqkS698vpR7r0zZ3IHopPVJyw7C+/h1QproHybsNw5VtU1N7Lv1N8
IUmiYWNKaQL2GVmbhn3skdrteyW8xE2dKcHxpBFXcF2puCcoYXg6T+whEtvb
FBcpxTa0cA6N2c4/dUtvsNi1mgJT3P7QKg7aG4L1l7lK6WarxFNQFUeCnymk
GbmQeGs9ERfg+q0osHli9RY7v1UhfnZKswNpHEjlPDx4VeS/t9I9Ft7KzIt8
ob3LG1DopeSG+/BUr1O6kq6Zdvn8AkSi+M8hGCoeGVevDNDoYqYb+cFqEL8I
SOFKKmKF6zcyqtPDdsPTjeXFtOMXb2I5IdbKQeh1pat3sK4W76ccaSFg4/7r
yoYjuDUL+03Iu2GFkF7FCp7aci9BCFZTtKc72QfmIYFUaIvEaH753tY2vl2K
0FtMfBfMkOMS5YsQXnHSXZ4HOiF0wFAniCoof8FxuMF1EOQSQphNTTuDFJxR
H/CRC2imBvIEWfKwXJBpdK1YQeP/933IvealkDned7n7NwscBSeCzwEQcjJc
J0oLAuT8MMXEA/8zXrrRjRBXr9fFZntYhjG/mZwOhAlFlbljvzxgkyA1b2R4
rH65S8++0+9irMTRVHnFzSzDsdfx4ns2tE5lIsrirlDr9qjBZJOGbgBoLOhX
w9mM0to04J3naLpBSYNYdWRIn0bpRjTR5768E2GfyXGlj5uNiLbOmat0E5mD
TNkigfeqjfXwAD3Fsqfl7AkXOwExOmtftL3yxRftHELGXQfa9uB/eP2jsK09
zcolkkq4qIJ5+GdSrl+5p6cA9pkeAMLMlssfODBuVFQyrtfLeE3lhrA+aYLn
DeNws9hIQlhtSwkf9uAvzFcWP79xldqrZV21892O7ohSDlMde93WYSfaGFe5
CZP9OH3JkPIr8fVCgIuEMPs2S1am0EXjlY5hK5J8WeVpy4qM3cZ25miToWeV
OIQh4WxpIYZc6nwbsOtVxaonYyOw48IztYnJaBom5Swki3tlpCR2GPZ9qLS5
P4x4vjt/MfOEIoHrWKj+0vAqqSf2oTS4kTTaKemM4ll4n15J+11JXoRUZnEI
DI8A9H36NVoGLwRuj6pFZePexJFXBHSBi4FBL1t9e3ccP7+AhN6I7sYgmDIX
pZAZmirIQztNYTDn8Y6QqBBGr16isysOi25cbR5KKRZTrJj/9KKHvu8X/StJ
wXwtu+oS3xLEt7+3b+x7ugzexpLaYUXpffHOrQQIBYN4RtpEWaWTPWhaw7mh
79fLWt49kGBbB8K5n2Q8vt6TTJkbNBIIlJzKx42hPFMoGB6xX5APszpYL0QV
E0YD8gPRdR10+Frh8wJixkCjR0uPmfsTM8Qr4fq/JrvtQSmDlSDbzCPBQ9zv
ohDWnzZdw0bgOhNPqaUgcEAjbErlfNLQquOOQF8PEEKrx4Expj2M738Ghm0S
jQkaojuwaK8OeObHH1YJhenWpMP2l8vjus43IErK3wBRPxUeqqed7+JI9jKV
466PwGl62eX3En1C1YeoqspLiH69aLW7YWozvbeo/CEBOSfnJHY8akiZBmrs
gFqnXyaurU18Zs4YZAa+u15dH0Wd/xWq1YIwfw5k7WQ+iZMFnY1GZqOiDgXn
1QU4oTvELTwlIaA+RMzLgl7vDx9xJSSMzsWgbg1a5tS5cywoxSOnBSKxtBn2
DWtTneKCLVSOtwlRxljpop5WhIFtYPZ2qyaD1kfre5t18s9JnH1/gs7db5I4
UZSksfT9rgBHZYx1rHquAA8HdnpxQVa2IovCrBcsucFM/N6DnIj9sL2wjG4R
wGZh1U9mzUYziQSs36lZXlJEKYXIk42wl5h8G/a53pXAVeScGzpZofqG8iDN
EMnR1KJ273q+1QeCO2bTzhozxBs4/4OjvsyXhTtCpcL1zPDB4bLw6wNrZ2Xf
tGBZBddlO9awdJDJm0ytAExP369Zaaft7KMoVpUc28/IigcD1lf96hq8+nxx
iiWP0ofNb0KnsXZ3tNVc5aq5iYLwzGRYWul+MXc5a4IlpUsRG4lvsRJb0ALr
KLUYQHB1pxT1rWEyhHYdTSX4Y20VLj7edZzNTfKxCmaZZ0qWopNd8E1dcI+t
QeQL//MEvQKD4U/b0auU71Qpiqn92ZLcM1dJx8BzzXgoNsxZtXa8fuHX32QF
3HuCbYUqSfzOwHRjZHMLD+SvmVDwnkJv9gInn8UYBKOF3bYS8mB86ac8VyGP
9OEzOtk3pvxDhr+L3qucFdVWQvH2iuEy7rSfyVOFyUZDdTL5itITzmY/2mB1
+sEuyJj3O6cOOew3fkvsOdrPsT2lmLQoRpsuu0GAUCgdEpm3Ngm4GUtK4m2K
vM+zI8kwpg4pYceyAjXcEqomC9dgF+G7dAahnel0ue1edi3i/y5J0+Ebui4O
nou1S40BWpemr+kDnuhoZVx8qvR8w9uZ7kxjHgSXGtkACZ3iATDuuewaYZwp
eTNrh1pZ1a0qixVTw1sW63iv0TTtw1pEcYpFZbsC1rly759cjKyaLMott2GN
CxRX0NSRE1iMs+WZ+AXEbaDix9gEdva2qGAsu3Xvuuaoc0bsk7fySiJe5TFY
+uxtD9PqEFbR70zMp/Z6pPLynEyPlOEtyJUVWbCfUqxt32TgEQovKrGpxVj9
+MOAK4YagpaYEab4nDtA39np71kuQsy5b7Bue6+iebbkcMf3BcXWFxSrZf4m
q5C40d1dS5qPPTSV4JO8k/aJWJXtlwf8RaEvnc2SSLzoDtqjqOiuFD7o3dzf
Azigy6Ke1n55jL0fTiax0B4wHF+7KCt9m7owiqt0y0ZJAFsDuCrk6nPBe3wt
bN8p7tWqcv2bBVU74LL5swxwYe+wEHGFfUPtvxKwzrnc6yk57AD2xW3+iAO8
DkA4PUIfBl2DrrHuh50MxT54ssetaDDopvNlvz+Ubx0Ae5oCTdDs1WDQII1C
WMItSRKe+hNrcbALjHNnZIIMlF/jqQsty8jpNYvzdJsUIZ63xdmQqV4lXObC
HNBC7xAVS7EhyMLSkXdfeSg1+g7SZngYYU1mjNVvS9nI3V7TNo0gImszx/Gc
CpvWo4zZVNMPKOQrqgRf0Y4apxNlQ+/rdb1vn3A9JfwTV9lihWN03cICub/G
J8+4MjJWr1sSx4aCSD4OE9Zwbs0mVTqRju+zmvXItPmKg6mmQwg+2XnhBxL0
gfJurEC7b7UaIFR/dX6u8GdsYmXg58wntY6ZYkZv0Y7/kCl/WWRf6Q7Chd1D
9UUa73sNlEqmrPDxKbFXfgA9VjOc1DP+f3ktus8xYNr5QQ6lp53ZOaz7X/+z
Tfuvy7fMgiv++MCZLtVKJbItvx9ng8OVRFjJ+UZZ7SAzurFt/FQDYnis9Ism
qRqpglKxSXFKwFoTjMMLY+6hw3hytGIX7cUdtaYgSdegUJGriUAY1b35MXOb
4N9DSpYDiNHPJrLYCVj+5EvFg6z5dJOiuxUqTDqziKNrcHaKY0/Nn5IPvTWK
jTfBzzeUUCQrpsow1zEfeXBdT5aFKHSC0B6Y7TbPq35nTFa6VSD8D2dcxn27
5spt18gJt8t5FoqNeDGTYdqAU7/ydC435gPBstIAc7R8EICaOzbWwYTs/tWG
H37ePUDSokrZ1+3KZfu0Kk+orieyIihxBCk1y4Ptqc6mBoemfDsFSBCFrbJW
rTzay48PUJTaGUXcFukljpIrEg+OVFzMqJaNbhrPm4AgT0Y5tn5EDm5SzXym
9Ge8ERwcaQ3okOmByoxf62plZxTW0lXAxXlNxm9YXG4ZeQbjVygcop3OEQ9o
dRqTFW5qF7zq6PVichtQa5PhTphit25VgfBmeMe9TeIUWuCOMGSVK2mNJue5
4yp0pC2aePdGw3qhV+j24cIxEjWYVQ4iubP8BePxYsIZ51gQnAOKgkLgaTMh
txbpcxKpgivW0GMZ3sWUeJDiVEdC3uJkyFxcfIXmUBdVC47axbD4+aiPODcm
t/KtOaHbY/qt9dHWVWntTxz43lah3darikE5NeOvkamp4BRX0raB/37EIwzM
XF2eOnsN4Dlb8Q1K6B+Q9BtWsaSwaPiwhmQZKaixQeekkX2enZ2HnqPFHy8r
9rfI8ZtLvTL7SPVk6rJbCtWI5dmLtTC0V1namtcuyeNoHniivsYjOwgkgQEa
wbHSOHvL4yzyvL1KvXeyrD6Sk6R7sVhXoZMytPFzUL/fUi7rVLnSXdirDFPY
W+lsyBbFraSthTmFM2VpIqEo4spM1QJK0plRNWPyxBMdBbdrkGB4yemxseLL
mA/YmANi33NOXwZ1tvriSYZNCcVhemyQiyGD9uGHHD/8ntcO2dVwgWmvcGWk
oY0yvsI8UFty+e3c9XjhFqNT2MkwEbPz81Z1tfc3LdqyL056RnBo51atRTyJ
rXlmaXE83HxdAFbOi+UIKMegdEhs1c3QrvWG8F8nPW7xlGMlE7WsuRLxImEO
I+C1gHn3awKlYLIuVBImD/hgbO/YLc2sZpcNrGalKhXXLeJPUr8Yn8c3S6X9
Qt0v2SShRcvvRfHYQfadT30t52fcVoolz8W3iyrmgzhiXAH7pYjqGo53v963
qO7r2+MSKECIEhcEATxqy+nahfh8v4oAJMexdCmAR1+eh5IJ76vyWZOj7ZjW
6h/4ZGL9zzTrIqVP2dQ6WB0MdcelNiLgBnwysDHbyC7NhXIMn7NVa6oulWcP
aCEWANlEE2yfUuzSQj7cL+Cwy/QQPTqQuSt3MkWMWE1u18rDrDriGKHTqxRd
IvQp9xkIHaiEvnqZTPvc1Qdt0pPlRzDqGSHkyz04Btu29gUtOs78M1lH4fF3
uXST6AwrRHRTC590iyKZ6NeisiiHnwMWD6fV5i6ouDotRLHm9UwhO43vL3ng
DW03T+s8XJ3ni4vhvzFKMNBBPCYeL8uIcqusqhq2YW3ql/KFsX0/kr572X2U
ABKoQqh85gTSN1GnynTpHNHvBMvKHKg6zhmTzeG5F6TwDZx6KDph1mmLW2RS
+rV3zxtInWj7Yv9uJL0Z1pMi19zU1DyH+C2PAxKmu5VSklp+He1LkLn0KQQn
1tkcpvirg79Hzy9zTsOpUPZGKFfWQFJ66bRtkZ7vUaZuHQJyYqdjOR96Tcwc
mlrzImG/P8A2W6g0CcCdUe5YaE0HmfQQGBn1p7r8qR+gWB3UKndvu2kG6qMr
Pl/HzNQRMgfusDipEONykOlYyQfClMqU9J/5z177TMdKOjgEOp0BtYP6Famf
DGOPVX2QCpUGoidJkjcThFnmWJl812MFu5CLJAXFs0HKn0sGLbUqTlpaL3e7
LGBXlezU1iXT4BuW3B+022Lcb6qfKkzK/IP+bdz/ajn/lDb7SxZwqMMPSenP
kGKGG0y9tl2twe+5yzSFZsIvRkDgav2TEygJ3VatJbCMLAWOXNZSb25WgOoS
eCREpiPWKnMgA6Vjcc0o5vB5jPFJxSDMLPnC9NRNWVyLwXADT+S/v5t7vLfv
+Bz+jtBwNDnrmB5UoVyi3k+FfqP/1jh5C/M84UoKx5uxqLu03l0YNMrI4BP5
M3GB4hYFtmxP8FGYQTugAcwTtWoG57Rh1O6dA03uXVKe3sLSunQ5hlHGTYJ7
2s65JVtHzloEpvIseUbQhBi1+Xuzl4z8VQ18Yxd30wtxg5IDe6EO2f2DALux
l52U0IP2MCIOKxQSQPBtTj+w3/f3cmC3XxrhXj3MkGTQfaDuTi5V5ILxtz78
YCmrHXRESKVVZ+colWmzj0BbTSq6tB1+E0NAYHOhPIo3iV1pTIukJ9uMfXtL
Doq13Em2a7FOk6PjlkM9v8pcojN4V4rvGVNHk2HAIMCMXS0ngFS2JuBJ+Dho
t3aePAQ1NHwpLSTcKTo9r1JMqwrlYBm8rVxuh4zssIE07NUlmc4Jn+pix7lW
lTe2osgj2G9/+WqWFwcVEJFBdEu1qBomzBqgbdrN0gOmlBH1BKocxC03pYQl
PxhClW4YHMIuAuRl+NA9KLTF6aRgeRNw0VRC807I6mR5c3oQnxI5edLl4WGo
pDjjb+pshV7y9RExFceI2mSJWdLi42UgrBQ4sQgtHcVKs08QN65LSM/jrG6w
7fKVxU/MxZps4ry2rrAleMiP/5KjDzWTmTeRx8H0bcnoo94fFqS8dBq+/iEx
qoAIaQnAqXYjsL9SiH8KK8weyf3h2BhBVR/+EDy5ANHlTDcAGrUZEFWryaTB
qtZFTYZrF73eAHaNvH+cQptnLhpdUUsjlwt7pdEyEBI+fvTDWI/eh+z75ppe
nDULAMlhvHYOtkTBixjOyPPOE0yt/0sDjEJjtwYAna9m6s1L9qWSK6RUVfp6
rpWFOSRAlxKwHf6fupt6x90qUlEn8qpT/t4qv8SOM5hw2cZtqOvvVIK0PSIx
YvhDfuHw1K0QygUKD6pqHZjEEVUxrg8mvK7PWfxvU7XyqGOnB6bzHuhe8ltY
4tkwWk8OXIkv9Gxd9wsFWryM2enwhOmKxsn4RAdqKT5h2Ctl7wCObSxEX8SG
tX9i5GvXFdQmELimTGk4MLKUb7ENnhowPR1UEXadOlnBQDyw0/p5Tp1tpX/G
YKlrmSiczoPograuxwSbNdzxaRGEAVBACqWYudHVvmsIaIQGuYgTFqyivuz1
oYqHVYareCg5NEv3wTVGnPWNJZlRND4GOvpH6r+YWdNC7R3vsr6uv6S/3/nN
QLWTTue1jJ6FkjiAvh0OFoBi3Y873SWpexUYEx9+PYhsgegRKAapeSu+zuf+
7KWhVR8l95vUt3DoGZAfbUk2IzeIfrSpRFhkUzAXy8ohv1A5m7Milk3NcLp9
palECvtMuAodPK0O+N2lN4huymxsbm1xmfhClL+HjkDn74fAP7pltPtNPv47
YDN7Y6U6qdJcCW/aS9iOUWYRAOn1b0OzbWKXIR+bUVVavmEONsZth1MUkHOX
ZiS7lCczOyMnU16zdqTqGFiwdMeDZ+LRUEu2Qk0i2Q+ozsWhu9/yTNyevaPd
Gv/kX/YNYXj/yoHnbrD4EvlR3veEV1J+/ogbiXQhmgfbyxCwvj4pj9G4t+30
vgbru8YVU0Yis+dOAYZrpOhZX03BexsLcAeOxtlN8teUeEIfwfGZpjPIxJlx
81XiNvW/GDdG8kswvY/WOTKQwjRE01ei2KmHZzuCZeqVxcai9yJuIUI6lZEs
G1dMG7v7lIfxkUa9FQGHUV1n9O5MoSaqwPsJY1ACrQzPUUZsapMmD9T7IrWa
laBzSWznIQtfesFqS91VpLy2JpKmcIpZz3p5WWm6S48AclLHpJ+AYayoIdU8
bzwA51M2rg5+gANlpt3tHkIZ2Is3ozbnnM7bcNUGx4J31AVyUwBqPwwL/Yph
mIyv9CG4Ql6wdNyX7ZdN8kCiQEh44Ud3cgYjhYHmP5fMEMxOTOIWUWcAnM+c
YNc7shDIcQDD/vq4rqDBqCRz2dIQsRFcLbIBbb7YCYMvLzd62B3T3Dj5ntXX
ymyQIwx7dqTQFr4MD+af0eLZy7uGH3X2j32ZtqlcLwLXNTvUnHIXU22LlFLR
rSeoRo02RwFvlbExQlJ+eGyZVsme/8AWf7U2URa5D++J2mKnmB98jwLpEbSr
ElYkyHVnmUtcRtgrC1CQLVUrrwBvHOeNH+6K9wq3bjBOGMA3ZOgWnn/D33Ek
+uyYxjs4W61nUaiyKd15Cde7JATssGEeYSlsmAiV41K31TKEj5xwDRZtZ6hi
0x2pmBVbprOkTz84xlIX4Z22mx0GofvhMjoAV4LqbtuzGyw4ExiYVekuvGcJ
Tddbf9qMiBQ3gpokEilCa/M7Kt22DtXuPPvZAGP/YEsi5K36LO+nK3//VkzS
e0XAERsCDKHxiyRyn/IIIGvXxNbvLiUejXI28MzByj3CA239m7r0eWwQgBTo
UBZIi+G0SX6qhTIgb+j/BSJcJuioslJ3IO8bdgf56gxCwP8NPqc+u4jEQkN5
yHnM8ske3Ny7IE2IHdyQDY10Qnh3FWtHzIdA0d6F7sf1UX+OIPD8RlAP+WeN
QrCIVedUQcjz7hHtc49HNv9cUIJdAGxSvvHlaV9UE9eYdpQfCJfkL5no1VTp
Z5qLEGys4rjteK1pbgSmMc4+OKIUeQxvFRQO9CABNKkIoYUStdoKtKaLryL/
cnb3aDYxFaLOj1C1ul8r96FLa0OWOCwuJZi/17XmaE6tVAAzZ8+D6OEsE9mi
MghntcqlDiPbQj+DqiLMoDETez9g8MoNKmbVK1jAlB0cGhCrumb9cFfuPCMO
VPoZ2Yb21Ms2xh5G+Zp4qfOdJFn60HmjOqiebiDq4kqUwwuziNB7L6nQfj1W
Zfq+NLiYutMHUr0A0TOk2bHjxsYds5acn4TKIAei5FaAduD5I0u6kIdQaHL8
IyFkZnxhsGLgCZcIg/7JNwpyOaH5v2ZXCnvYw79zSEs2B2yxXDpxIzcnft45
Iv38uck4PcgoKO+2X9jDbIVG3AfKFrMkcLUzZZqc1YdLEo3dopbNq3GHFvmn
VSJm1BwByPBUKFc3EmEa5AxfW433IbxqJrMr2iukPMorQwrkZoKJs65IosbU
LSz743kKvUNzutQRHAfOHfh8N0T2WtEyNMT081SWa6Z9+qzJQgthHlqpv8aF
eHaxe5I3QcbHWf5Y2nfBcyj9X+lKJLOFCB3PRqwb9ryivOCrIkfRHZqh+v0c
9MGpfRVLUk91Tqx9Ciyi4B5sMGLOft8mFUoqOi7oBdc78z8W6gZq/5YQWNpc
ordYldks8+Stxlzn6PTMDhtr4hbPyufH2VbYvoqUhQrr/cWT2HpayqP7YbfZ
TsUtTPmUUCJhxQlYhwa2oEcKYokWmMhtjGYJ3h3E/Gx9MwXNmk68ChDb208o
wOANOUXRyGLMq+eSBCEDceKwU5tqfdZ9N5XgbGDc5wHO7ipSjGbB9Vu89Myt
hOAjoor73aZgyKpqbLfr5BOSQRGpvERtOCuVjeCf2f4jwMEPzhl2voCfMbKR
XRCx8bepfPvDIUStF8YglKv4v2Wl/CESRyDVzKgFx+DKDj39N32ZMo6YPFzu
Rd5UvR9nHnrq59uAc0JmILgWLhltWVl/2d+5FYvtE7v8rwCJT3DfsA5boVLX
EtNSh+1RQMdHhS1hWWNnGbj6YC6hhXhUYAF7ZYOX9Fw3hnCR7/ATcvar4yNH
BntqRpa9qPkx7zwwXI1XI9Y65blj1UigU0H21jrANdxFMCbtK+0Iia/enspG
61ScA91xf7EnFj6seYbEuBX8vT0ekDkr5n83FIvn6Pldp0r3PjIf8OZv7ZLo
uuA027zCfa/3hkUVK5KY4N2KDwiKTv6NHjLieHafl2W+pQocY+EcgBuhLZRy
P/4F8yLLsNyh4T6CIQtR7TtlLhqrOWJf4ykgNDVur1IXk84562JGxYvNY3+H
ne+GCq6ShBpdGLnseN7coynANG77yPFgZeswKRRqK6Mj/0yJaOQaw1FfHEEE
lWxAQc8t9SGUme9pNeHoINSY+18QDycBt7in1pi1TzHXUnIwHnq5vVNMKTUv
Aos0FDTHR6BTfOLkcHlz5uayglHG8BQC2Smbbt/sNhTKaYDi0KehULETEpag
osHPkPu+usY30mPh8A9tIVMn8thWgW9gwFDgSZONH011d4+Bfm6x0faLpfAM
bNqdph0jqa8QMXD1C3CylGIJLdLKDERJ6grqHz2ow9USB3ehOmWJK6fzQLX8
svC8Agf2wD3NuCR4k+6vuQHfibgzpVrGUYKgmSvImk+D91Klmur9L1o2rVL0
/83bCIO/EHkI0pjPoSV8EyEngSLpWdAUrXGY5DZGTwlxpgKoRRf0AnitAoZ2
rw/eNiketDcttWExS58va1OPmNYyLfR/mdJbfnVgVUYT5znxAyGbhePF0um7
g395jRVLOUUa84TBYVIkcWRy+4Bhp6igLZpPpLXSufdUhV+eBapWRQMvGr2e
SPaVXWul/zEBKHJifGsPRk94gdJ7GVKG4Jqp4XWKB3vX5dOntIma+4C8g82P
TZf1o/67qB9h4nLJiZnR6/dQJhs/niLjZJFII46KcNiwA1FwGtXsS9qyf1ny
5zPYDaKUNV3kfsyxK6TnBZVxMfm0g/Mykp0mYbyJQn2i75N9XSwlAR9PA2uk
lZ3gck2mpx0xnrVA2I7/YRLJrao35QdXnbNCW6HT9+KQrAvY+1p5eG7347eI
cBF1/F3zfLkCdSLeQePP2CHDxIm6YvMHSbjJn9vQEkJfwp2mvZcHfsovedDa
gkm02LAmz01RpkGWGyucIVH2aF07l05cstUhFxQCoF5SyKmzqNVpIB4JUzFk
IMJqS38Tb34eq6XD8KSRkqTxgrcYJ9gmTelclNW+pwCN8QJF+yxlwZdNJ+5r
tqXuTb2+wcM0hKXwKoDj+WE70zn5jcHc8tPG/oOb9/zrVXUqHX6kBVb0YjfY
AHkQlTsN2jiTzuNzrwrmFdG4bIvwTP48L3yop5cuis3NfgJsoLckZH97PI78
DywAasZbzTzJfuEn7BOq4It7PqY3pWJKvL+JAu9B/1pF7m7KL6/LGaYJ74hn
Hcrb/q96K6zaRSpV+MvsbExvpnAIzKVIUfmB1kzKUMYZVOq0OT7YwFwlXJHj
9DWNa2JhduxCT1hv83rIbfSYAZ5EQ8n1hAGnnUcSktDfPS7XR5e3lWvEJ1Wn
LTVPDR2Mwioj8OQJ+XD8UnSUsGMt0PyG7RUCg4XJ+XWOq1UmD6xmHQfvJBuy
prQ/+paNVu0aJ8Siysj7jmgJKImefKLjwroc3yjVM5aPSDKC5Pt9XUp7shUr
twZvu37+d5FExkyAh/cuq+b8y09tPvkGlwrDyDhFjsytt52fvX5pSngzkBp3
Lx0oArEpLSL+yY+x3zLP485IZstA4K0YBvgjGbt9W8QWQ8xFRMIAiD/LLY1H
nHjuPQfa/WtDz4Z7x/GhNjPV0KjOH0t4AFbc772Os/HJYmxmZDrcwTolqLHU
+MyIvqDzRnyRf6GXk7PReM6Ge7MYIFywHmc88jLrtkJlqnu4GsY/V/98n59d
5LoYRzYqr9xpXp/rvsz+eCW5SeRUGQkwlynHR3QJXSXkzkTV47uUhhvjmgyV
EGVdaCDtOkQ8IztGS+7AKE7NG2b4v/wWZAF8RSL83Jz+V5ieEmKxDALBeMA+
ulowfYR5L4lo0fnjUBkHWSMlSpC93+o8fMK6wf9a50myXTsUCG8K24aU6IGL
ACL0y7zsRySACalfeLB8xRcX3/3buY3K9ipPp7bU7cJgbtV1o81PkTdkl2LH
L8Q7r4nh7EiBrXBVEvpux3KdhD3gBqH6RgA1B0Yzq9Ow+2p1GgwJfq+GlSOB
8Yu3kej5/5ZpP3NEpmBtrowOd/QM6YsBlz/nAHgE4SXPVCVzFtCWkgku6OZU
/9+6geCdY7uHlhz4QTR1RpW3tdVCiNlHdTQbgaThGTOk6IqkMNc+WQA7pez1
WQOmLc67xKLrMlVAvtYFn2F2Lx+9vLMSazLPlfETRwrCJZvJz53jRMfXMx3H
9zz32i3KZnfXA7f1ou2WfOgQm8xmGpJaIRtiB9Vp5j4aRz5W2LTHgg24nNuO
sha8NCj+mAf/A37qlHsBQenxcSajYGFOZdCdRjkEkmLACi35tZY4k3JWy7Yk
JQi7h/dOrehzVWFUkOrFdjwWd/gbOmuGtakrUMCS/rH6TQkUFxDr7S0Vom6K
rgenR01i9V9LSaibMyPaYkzPrYsDFvMZ8AFZWFwRlS/zhVLTO5yJ2TDXi8Z2
69ezT/7nD15ChzbkWLqj4TWYRr6BfbKYtskBoePYFEk+qscozPpJNHbun4uv
a9UnOrYL9/40WX/Mul1KjN6EeaLkgaWgWwKI89O9AWZNA5IBfdkcdzrXvy/p
VlcUPLgbfyBC1RD9ZMfP5YRANG8Z7Aqq8gG8nk12mPcNyUhLwVN3NRFmzm7+
B9+lE6hUG/CJ4cCZYE5EgczzjPCtEhVkda3+Tq7lX1IV6nB3WsjXO8mU3vii
TRGzenQO2AKELwlgpJ5umLWD05qVseROBsr+7gxdofDqtrHNG6XV5DW7hU6A
6ifYCZxy5th2b+p/B1A/iBMoIAXepeQ1PU9kdy+dwBC1ku3yLSwFIaX7Zy97
fH/52jVPxIJ62MTGe83PWXwzzSpdc8nu5vAodY2jE9su5kiPt+NRlA/ibzB2
aFHFiq5JJ0Kz+Tp05QOQOt/DwVnNvVVY7lbWiESCYQMVO0lsXwoXg3d1pxb8
3p2JnUAfbw5sTx3m+hviseQugK9oXQIn2mz5qbHVjLLb5qZa6ufNLdScerq2
O8YvLum/HChYS8UBqPBxZfIlCqFbKnEv9AZKG99CkrxjWcOzHfyAtKAm/A1X
gmxsldDT0xWG8PIzYxZpn1xafBHRkZCWESO6zg0rqPMvLkeHjWBvxeKYo3k5
Wes0De9sTfa7PCfCFMy2fTTyoOwIJIWW1Boe569fPrqg83ibatD2sqbZ8Swf
mkmppr2hzUIUIc1yopQGqGclfL+0kPy/NV8/B3qDxpbnykzfB3F1kzWHfiC3
6TzruqgSe5a1EoWdh/Ni8U4j8nnBb4msQX14WR7JLQh1XN7z3+/Ckbf5gMDo
UyxbGHn8XIB3qMWo/m27d0es0MYtPpaq7mYhg7p8iuwGqevklHw9X5zOFLKK
a4eM+13+YA25JEc8wDuwp8BQgKo7XOBeNAUxciXS1wFfkACp0a/UpJPXrRS+
I96RrfmeTovyXPOjdMjD0Vlvdh2gPN15l3CXK/CUmUHurE/QiytKmG3qjoqx
K8bBBuQUXhuYQ99DELw3e8oXjKfNNb0DL+ukBQVjfifyRhVg9NRvOhlGrSMT
FgNnhN/4t6OOm4H/Snd4SBCEniLmMixO43nmb583V4W9YlwEyeIMlLRtgY/d
0JX9P/KiiASOJIFDl1BV2DfpE9yDj8k/zaujsyBpbrwQd3THUSTIi6U3iBVJ
ktesw5KtoImq/Ap+l00yWOIvJcEhpcFyzEVy7sO+Ox4kANqxcdr1j1tITbFG
4mEoi4oXMnA353+xuwTviKMvUpod18WFYDRqOGhs2ap0Gy4r69DNUVqPN6T9
pB/BpumhLZeCLZVgx2xHnGBo7FmKXM0iTq0zb5i915TSUCykmxxLSgb9oPAZ
JE+N9i3z7LPIxiyHqB/f1cjmAKEj+5ZQ6+2GyGvOczisJZK3MXaTSCpHh7Qh
sFuiiP1YiuVsSsdE9xLHSajXhxdHUXp19ND/UAjli3PCM21UmBOW0kfX55rK
uJ+Bre7RpBZBdWsjGAp/chyktds9AzFNwoJp9DKVaq4Y8mOKm+TqqymvzSJy
L8QwwAIs4Jn8fit9QqPzRTRSWYbs7M8oNOljrviMxsbtCMGIp810uuGEDZPo
MJFv8l7DOZ6rAcF6KVndbcpCLDqzJFK3/varuEan7SZ6TXUGW+gGre8TpPAw
ty1/6/12OasDUFWzONwI7oG2+2WPe3OPzBK5sO+XKwrr4XclKSRzfwBIXIAy
/phOkE7v24Rd1xwaNA445U3EHxK4UU1iCctrN9jTtJX70VAhEVGhirYRlG0o
68fnxF9IpZjkHKCx2dmZTuRZTLB7p7RtqE6klddPGNi3M5hmalruu9XaIHrR
uoVvQNLjG9oyXU2GY2nQpSdSEmBnzqX21B4rfHi2w8Vt362TNQj/iJ4sxMru
n8W0oLjxBsLFYW+hg74Co4b3FNab0ZnPzAS5HWr90+iDMHix7A/ifO/xP/r4
ylBgS5GOU64SmGcr7Ww/eVURMUb9KG6KxPXY///ITqYDzAtBx+KUhFNVi30F
KI72FmhaJOV/cyUIvw4ETqXRSFsCCwbCUzbGMXQRTOIzfbUVhJcHQyUulx7m
FgXs1gkjjTvq4LPLDb5cS36ZL3Xm+eRhzz0DUtrwXsjXNE5N+FLp/ZMu9UHJ
zUQ+/yx/PQGMn7ddXQeua4/CMg0f7vYXBr3raXQAuV00PTYXW2wSDf4Kqpqt
he/3oPKrqpc/5kyksHbBK1ArE4zV4BBfQ2P0rj0LB+9UUVPgQHrJloUwtrtS
3ESSSSa/oTeqjSJIOQ5SFhI928e671E0yqrfmQAGE3Wwy3pY/TuScJ4IYshm
gXPqz5P97rif2EdSIWU+gXaOamKwPT5iGzvxyGfKU5Pc/7HDtnYlF4Ods1X+
wh3V/UQeX7AXftoxA4EJzdLb6FtXvqTWidC0ttsVmv6wDxjoUaMBL/eC0lmb
Ebb/iSvsTzwKz0a9OE/QEy8/rssS/DsHLDmxoh2dn3jqbsajKggMIvHOO0lW
o+t5oSvGvRSw169f55duhKcQce5oDT/HHUmfwCXakdh7tCOAzJ30pCy+Su1A
Dq7bLJEgoQSDXFcTlRl8zJXRQDPpDrhhskjQj0TYdg/jm+hsP8sithCvtUDa
vNyJjnv7Pgni9RyEdVkBQb0JoWZs3FDhnI+wxQKQ4HZz1gTyaNKFDryFe36+
7yW3J/k80ic13kNkyrBIYtQnvNK8V+RdK1vnpoZkA+zSkRNIl715N0c+cIuo
r7YhGyxXCpZENcfnmU+LuHqITf8VRwpWRB8kPwedZfNIptvTrcRW7bMw507w
Z5kezDqzj6o2L/ahUgOS1CMyPXPoosMGHvnWHdxLjtsM8FcFFbJC1+As97i2
JoESgFKJKHhC/MIYn/A/z6oJOCfyCkXVq4Yni0jRyboKazfUE0Lme1WNhtkO
G4Mk6ul+KQoFn3GTR/YofWnxw0B2dPOErLkkX4Lb4NPyOWdMhHdz9HG2TCOZ
dFPeW+fk9CSWgmWs1ukVtAkwgNH8vvcfBaA6C2/NTiv7dOZYgAFqE7pNQgCz
QPvD+83xC1t2p0xT8quL2tYN3dNYs44QQ+z+rZAXZ8OaXSgeUR2CM/YRNqcm
AE8fx4x3vp6JxgwbXK7Rp1bn4bmE199T8HOz9h1sUVmif/xYjwRe8AWlqJ4g
4ZWLcI7Q8itt+vUh95h2vOCDRkRlXU7QlOGhPOw60sQuKniqr7VRDBiNIT8C
d3Rqk7tG5ULuTgVpqbkZAo+S9VjgjZCbdXx8je74hlwoHNGBqFV+OoDBzuEH
x7aiEH1J+adnkQMGaMrS3gsASHF8fTepC9wtxPlYxavWWLY9aVUfVwtWYEjl
DIiSMj/Bo/TiobLIIbHkKbq14+iodOZIZEawnXezl2JaXhLXqYAYNUg/FQGc
KA/ywwWQHSKg4p/LU47aDKaZfzXBDFPxZZFRAp7Va7/YWpYOAoMcjy2GGG9X
E5boK5+dAzNklS6aUh3OmxGaTxgcfhAn7dZ3DfXpFzLB5+g8cNBm8fy3pcyr
okKOXUa502iaQibCPCkY7Nk2MaPT1xsqcyyfHYHatdfc8h2eNipv/tE6nrkt
lLGdYGhN/tKzs31hW8AmzhzQuYSr0Hqzmo1/JoWimvB2ahfppxhrFfK0UXV6
zlIgauh52hy19FqZkZcVEOy8936EVKtMCIL8XwyU8INCuWGY7uquh1VLgiVX
2bLSUuIUUeM+Kg6TOfxOn19lJK/B+MhEmxX2Kt/xoQD0PBV9FUWpi9G9mkHg
3l+uyiXx8PGbRTe71NHQE9XvA+oMEQlQPLCPJrqxslEwkHiloG/vQOpe99ZO
1x1xFLvDxMnW8NRAJy8PfQq79cxqMCKrlGHkvAwcD4lTEAOY0UPz3MVoYRoM
KBq7H4ZYD5jRUuWHb6wKpCKwkpwhn38Mff8xViz4nlLohTMYA9cF7klpae4M
wwPDjSCch7ayOCSCEHZdBIYl5g7xdxzId2u5oxHHBeJBW6HJ/QHSi7fx6ibQ
ecbJ8x69G3heXvp2hqvo8fmQ5zYyPRbaeO5aSIP33yEPSu7ZmWAYtHUDY+Qj
lUYhh2raj7A5TG+vv6jJf/VWerfrmwuORpokvavstCGYsO7yId+I/m1AJMfE
42kKdLJd6wF7TEjRqY5honWRGt2aFZbmRKWKuhXP1xmrGtvzBQG+a2nhPhqv
IcryzqnAFrff+tPE0s9SpPEU0ZditO1KPj6NmFMfAVx+wb5gxRuNu8lcBnQX
OcH+zDn9BCLVnmI1D61EgWEj1fYY+8SxVw9V9vSp2V2a21L8KZUzFGu1zC4F
DH0OQbXnv2VpTbmmG3TGklP4JHCsLPFsKUhQR3dzOc4rh7hpEon9iWgRy/oR
fy3giipNQx0sO3nAGRwG50ML2znFuqeG501dFZD7Bm7YyxNWN2nkuLonEcMT
X9Ik4k7OOxMvilAuREO9HrjpT0/SLIzKyxrJwggp14fyxTjBv5OKHfDVzpy5
r+AeRpE1wyUdH2w4m4Y8+USWk1Wl71EKWZSXI5LFFPqbJviZchyoripOxqnN
IxvOG8kv2WH3HRoqmoaiKk65s1Lv/lJnD4GtCXON+IzV3SvgxakurkmImmb8
e24YxrKX12LO1SBUCwS9TC0nMTZ5fK9/uwm7V10TwiRWjDIVA6FKivUR9gPq
tLeJP9ay0Ent4Up4ZaDvzcv0N8VdvwClCwKBLbJypwpg19IQnt3bVlt6Aa0s
zV987eJkClwIgkqz/em/ru3GWhjoHQIP0ZM2/PKr+MdFhDn6hkWDaINS0IEb
uYWEpL5FcVVIotRSkVHJNDAaBH8JSRH0E+N5jHVvRpMxrLF4YpR9Kt9XRBk2
00d2LCFSlckqK3lDBPs5fOB/9OKL806xcW4AUmK47d0ObRUaozQFMVPX58AG
GAxQwShlxULLhk4xIcxwbbSC9KmS2hJT174LaRhC37DIGmTx3OrSo49mUlGY
4rSeZbGqbmlXwMufrhVGfZJkNkEot/edf7JAgcqmU0ButmGukfdPlKCJw2Z/
DvIu13uTo53+LlbT/ACQ03yAWCfmQiuzGsyf5bi5roG+HTTJZdl6iMRJxWzu
8UayX8jg7GG9EHS6GI3+D0ngdg4e6JYcMF3WZcBLq41xxlVfsNH/y3lzUL58
j/I8Z1SV7SVK0BCQVdoJ4+KNPvwHRHJo5fI8mM5yO34v2g2nYog1KU+vOiBB
K7TDq+Dxkof9fWmdTK03LbxwCnp1Zj04G8s/MUgDZRlbeg1op/Kcmp9O7NYB
a6Ye/74CgVMj/E8SyMpxiGknrZjqjVUBHwX/zOvlr1tKQ7tdgQPPVGfCfAJb
bgKGBh10K3wFCS1DG16wafbw1bZfiXKujzgsNz4/hoTgFZJfEgVoG8QsKhZz
nWx3M8Jwljv1OIlD2nAHscuA1QxCXYtAcKHcBQCQPknRvw3En9snbSfb3GCM
RXf3Q33jap4phn4mnNBiHkFDPv877rWfNWYUEgIxbzagYsCs/eAf3dwAgRYg
tcIC/Sx/wiJQ6gYQU0zV6xmSN1aDEEUjdV8wy5USt3Q3hNrf4XDSVRchRyVb
EG9VYJZaIYrbPupcAUQINbTLtewtEPPnXJoCR2wQh69TLg2MGWp5IdwvwDI0
IX6ZKnmfnsO09JasbuSYyEWlZiK6IEaUYKSeGNCUxMPP+vAOJ2pzmp30Ie0H
0C897VIBHgQRZMBfFghlOouCrGNdvJTktoS3EOe4XbHY4R5grEn0HiiCddJj
0K56Prn9lbiF0Jt7LZIH13KV0KLlBP7j8+it3DdoJqHeUzUmrSZpvkrj9inC
bhPKyEK1YuTPjlC/p5czyBF5FVNE4QJJoqEAZyLc+T6tkTI2tebYx9jTkHSD
SoRZjPUSWUTLLaS+YwHwrkX03Jqn76cxelSw+Hiv20Ws8WYaoLM8w+2xkD9F
yE6n8bnIVezj761XStl5u6RZc/ZvkTJZ+W03H+84bLAy5lMGc7/zo2Nj9lJz
RznYl0LqOWT0W2QtFKn8MxCrZKg4HzGUJAff3i6g3Hj+86jUx+4orHi9Mb3Z
EdkE08o2U5/EgqWWo3o8xIkrvlm5gGSuBxg6DW3LKqkCJO8Ib4y/oBmSpLTo
FhbpZLzoTOo0wdACAAl+de6dxCGSrO5DHau27PtRhq58dgp9t+D3T7l9+poT
pcaHUwVFeOTrI9LTsp375RtyufnukcKoeNUGWpuf4vUFix9Lh29SEujF4hWh
f5CvpNjkTkvrAyn5UNfPSDqhD8+eVQDr6joG8a71b3On5LwytYM2YrHe6h1p
f34LasYTJFjTz9j1uxg7g2gbQa6swDe/TbxDmQe6VbQbXvzNY0rKrX9id2zo
1Uw2LPz6BqYs/rZhoJHyXOpESelTM91lMh+zdbFlK740XS+WT4wHl2p6Tu6z
N7V7UhW/n/q3QXpBQ8OJMrTRUcikRzOLElVuvsPyyGpf0bnOWQ9v/rKSAeex
4s8yFYr+22ltG50dQOwByR83+9JPxq1EmK2tQlXOMHcUfGdx3Vuq9XbkhHL1
WlWOcTF9VUeKlObDASDbBFkxb4Z1Lf32lkoBOtcLraY+zP4yCCxV8DSl9CuB
FGWPLx58WRizaVqmgaH6t8DeQwy0uRjlOS8hpr53s0gl7LwKEju8s1gA2iiw
W3qG39sVHdnl4U+l+xVGUmPcqIYTj2sqbqmXSRPWY5X5oxOALi/93W/LRmZG
nmJAMAeKIsYMyoblOR/bldz/WsO1/olXWP/e86yzHDtsWPwRPDXSWcqR1stZ
9NTKy7DH8FKPMs0azRpiyQQaDvZkf+O5QP4caCFpFrJNI69p/bUPmTH8AohI
CmRcBxQJovIeZnY6eenqGgGZ67qmDWwIN90+fpBDHJwqS9KJCvkygDbEWL7L
tE9Y+h2/yMaVm/2i5TDo+SQKVU+D9U1wKdLtT7s1i60ZhDoRzVKQLfGyf8ZY
Woqup4K/D8QgRywVgTLnI+GxWrh9cBgfJna1Gusu+rkElKTKxluZ3lMY9N7O
GBFeIrwq5+PAdH9NLafS4CEzbN6HXrWv7qlWoQgtC2l0nIW/aL5hEZGAT6K4
MD9z+F0AYOoHhHNHwFvyF4alSrwCUYgJYXvVyjdUW0/LB9Bq6Hah9IxRXx7R
/QCqp5O2aimEiuJLILxEipzMO0lzuozMismKJBAwBYI8SbwpoPksKQ4OWk7k
2tW/0n4SQ8gqRy8a3TPKflms2FUu/f7jb4ZmWEVUDira6crzBHU8i/ss+Ky6
khfLo6CdiFfL78Bj7mqGnxbft5aNXMLHMQdG+XzkeVHDOdIS3zqA4jzItFGp
8NyEEnTpXRaYvxWnoF3NWby649ScWEMb8JV9sd4E/jXMmkBVx9HXjYDi3ZTn
8iy/UKzloYX9D9UfF7/z3kUUaiiZP2lq6ryGxWPtC3b+OOtxCPwwtXorux6r
6tK3zxIsWnG/tlwrL61z10dUDUQyQALKw7gIqVhPX2Ry0IbwAmziG6UHr4Q/
w0e8TXet+nJCTBCgfevzqwn+R+uQtfl/R6YW++G7I5CVxRtf9ncHThfw08rz
4s5uqOjXRVDv4e5Dr9v/PCvaGHqFifeSKUxB39Dpdjr7VHPS7c+TKZlitRHp
jh7+lw3Z6vuwG4OgNvgEU+9z0dSED1BzACoZRAYlj6KJASS0jZWkhLBjPVEb
kq24CNVRwPbBYHJC+qHXxIjormx1eb72kBdmNNooOvRUkn99MM22tfUorvVb
N3/tjqqbGnz+a6rF/W9r+VdmlKJeT6xzwJ90fO/ObyNK60Grw3+5+RZXIWU3
D84Yx1aV76dHvHUte3zxdo3q3huLuE52IVOcSxJT49yFIMDfLjsu7Mu/43Q4
r5yu2+ho2huTQhAIg4rWJkj4zvtFKioNGRHUfbC7eAw4zrUhF6PCF1frgvMs
c+L6ZJ1r4X47M7t1srHGQC/CwU4zlAzEJ9ltpzoGWWau+bg4C2tk5gpY3V1Z
hEwPlTW8UrVObjK1O85p1EZ8O5xIb5KEoFfcWnRzbbKmIG95QXO97+BGHwIT
odlkeTXmDbf0U2HOMgBb4+mtNktshPARIKaKBNrPotFfIIBasoQwmZCnI/Q3
a/KTvzm43wjCe6J6CnlwPfIdbTcZAJFOaG+3HY9/5QuKAmEUIuxF9nSFLkDc
YNjNJ6F6zkK3gVOpu9D5QayzgiSecBZI77waNn4QfVM8A4EWXsU7uHbEQAHX
DFNpb+K2+Rdi22s9kbihRiqSf30Wrd7l+IDyNFrVlXhtljRH7dRLbCrjZBWS
MjFw+wE1EdKNXBvIA/wJ5+moDZ3rWYrjIR3LeCmKv9AsFgYTvIFjfQmBh7fC
tVhimQg/z+394biOi1Q5KQXqfUruUjSOdsNCHzYQaKTYxI10okl96xLaVI5D
HBlhvsyQCfQi6KTi/WbKOvuWQPmD1Nm50AA1oki+vYkpLvQDXM6ZpBSc8m6G
6V8TqVHaLxm3ZhOY2Yb0x1nKYDEwHg1CIjyKRgJbjtcwNErAlYW1E0Og5z2/
TNK7T6ek4piywFZA2qEgD9XpsFe6I/xy3HsHMK70rZGTk83TUxTXxewKtoJJ
AazNsupf3BL092ZcH8sKd4cG39aF2lW2IXVGOZnZBZIGTXQC9TxBUGTgaTxa
Fo/eG1B2OPkuB3tYWa/dKXvbzCFinlKbAIRjU+ffX+Q2/nwBkwWbwIqI1lXB
ADyTdy/S3UII4sDvvoDmzJRSe8KKiy0H8NrauMZUupZTOPzA3i4WFNmgvrSG
pbTAA4NVwP8TYTBkvVhELT3EMbRHvh/KF6PWuCK7yej0c73SYUu6sA48GOZ+
4RLKeBRCDAZ6mvtQSha/a8XZVZoSNKUMMsK8efmMwtJt2DeinujmDBROeFvu
ldZX4zWkaviw26ZCr2/YEkRp88zG/FQBtsYncu83yOdsmBzqBrw4f45uOJ0l
4Aj1wiG9zpAAIgaSqCo4fF5b+YwrLLn7abCMR/hXaz3AwKVPx0bFzIxfDDvb
1nr9tqxIh5y7NPlFwFH9KQFLpfqRPR9ts+mHUtGEi6PwTBDfjwH45xri1JbX
IIUNp+cEC4E+PRsWVPiboBXRU4nw8ywkjdvl+cz71FScOOhgJLSXgLkd3Dxx
p3kGSy47kQj867BJKbOi2sV+3df6nQ/91lF2/yKrIXAqhOH+x3/fhFYMZwyx
SSVpN3WmkRn0oMQ1fEL53j2thCFZ+w4sjNF8h5Q5B/ZRZ2iwR9RHl0D8Gdrs
SNI8bBMcIjBcRMRtr4161B/7B3Mw8zPhodB8aiEfCwIUjfnPsYQ96E+UX+2A
uKMavxZi5EEyx3Pmyn7tgFL525Ur8hxjwbt6GoiGB/an2UzTWVrA7u1yYwZ/
BKXqgYiqqcOmZ1MQHMIbK6/YRL95JzAv7/IhESYsLq6A2/Do2RAsMZCmErDm
zOWVgNTTAJC4XsoqWt2X9RoPA0V5Vk61lwEtzSjokE1Xv1tNw8rsXpvRYosB
98U0NUR2029BQP4+gmlEhflDSv8jLopSzA9bBQIHhTOGFw9mBfJCCV+f6EQZ
/Zw7MivUM0kFqd/Q+1tASurEP+gn1XFip541kg7BpBD+rJcfD2m0bJXy/WGy
IQnAba2p4qOSyRKreoR3Xwu3eKKo2Z4ExQPvuISShudk0F+F+5Ph1nWeXhqQ
Ita37KQxKH0TQ3WYs5I/bVE4N6rLDySPpWlLcexk5Vv1SFZly45Lqsd7ExZQ
/876j+WLld4T5j02W/BsRr53F8rqHIFIQWaQ9/bLAXP00ftMsFcOPd2KAVMo
+99n1O04VRCNCdUeWTFOxDHT+FLK3TJZMYKWfcJPgldc6LNtU9C4grg6FhOy
TY5xvDjmI81PJhKXazTcamn1ShxUUBIMeBh0EM2Ci5W+5JieUxF38n14Dtuf
VO/ln49r3Cs/PF7gYljMtjakNDGAQTdXCwpIShfCkByosklDeh85dEnxMJ3W
GCmmJFQFsOls5I4rnV3x0yKri4C8kzFwnPoKFA6NySdLJmE5bG77QyjfVMX7
/JrLJ+xfxikbDK5keiJlLdgCodksQyPeLcDdSrgR/Mq2EA7pFQzJgav+SPeR
LfqkVcWAispzWMWmJXNshMFw8HIeKp3vkuqTxgmJ9QS0ruoppgr2TppqUGSn
ffK/av6XbTl97g8Vk/5Xf7efqvYBozhh657t0GKAjQ4E7PNEa828eclAo9jU
qGm2ie8miHCfhS8LCxl4F3pUl7MBntZWW1XT9yHn46cVETs+rchFX+O5Z4AR
lbGVuEmGaQapXrSuVgDBrChVXtjiy2PorvFP/j0WblDxX58AxDh1yrfQS2j7
o1T1IFNXmgsmSgJb2vSEK/Cd8gLwcnJavLMgChgVB/zazJ4LPPp8RLFKchBp
XlkUbWynlf2uTS19suhU8hASS0596IG6h9UvnPCk4CqCJpQ5AujQR13glvlz
vuj/vaFPqOQaeQ75EjtR/9hinusMSxAnqQ3x8eSsWA4LsWtntCPN6TNEhiqT
Jn6RBH7KgKVS75LBzQnpkPDEOKpx9/PEftNLSY1tXrJKsIyxdF5YC4PZu7mO
ZPOr+sjahl261fiYPgy+QCBrmn2wlwlFcjC3wjJzji0LOh9U2UUUE3NgyG3L
ID/sF37kXDXA5Z389mRnKfKzUYni+YzJ+NfpygMQldfBuSGCLL98OMseBfOb
O4Ei+k06HkAZw5nZ2iL5YZKSWJmzNtYk3TfKfvng34krhde3zcacusHlsgv8
nZ1VcvtvwRgCtSkLf1M+Lx7EUPs65d7uGiBnozIyhowK3bNj9ESaPz2YSJgp
dcWVJI7fGBuTr8ltXxKZYzfJBqYC+0Km2tx1itcmkzSAGiO0B9oiGko3LZWZ
PHTjstTsLldHnfthEjgQzKMbhTAYsJXogFTOUM+oD0qKM/KCrmGnW9F1HZOe
pB1mF8zNXAVjfA9XGhqjvinWt7mEeX48Tu4axPGPeGcXyqwa7S4cu75Fn1l5
0AL2LOrrIaykEbuSPR3Dl/5TGZ21mc9xbJNnRei7GSZFPpMAkmhPt4NcbjSE
cTxcfvinxpeYJskvZ5V0N8dqdB2KbwnI6CoAB9m0Hc1tfDdndey2DpcOVbdX
GdIVPXurKHJJlc2JvDzPAV7jTwJ5r3lsvovyI6qVefjo0NmQG+yys3OVRdGT
gckBHE7fXr3Y6uFKu6yEgHIzJPEqEFLjhn7AMzAnH7UlX+TaRhODnCcHaw7c
v4xPvPQYW7Z+xyjUPFr74HFKD15VVZLOZ4xRZeCCRNPmoNHdAeb2GSLQ0x0I
VfPFCeBSNzEUPtWtfzpdW80WgF7/NDE/XFzfTZr5fgavepYSxa6c3cx8mcvn
PS2hMgvspBW8xxWE7I3S1BLvjbwDtsxC1jwVeQHRhP6tNgiUsmXENaP3nmjZ
dx0BVLgstsLVlC+4xY/6dN3QM6bkQVOkSgvDwyGXrzd5Bz/ooatr5ZzrMoo7
TW0m3JAv/vM9jL6znCuCAMKUeMfmmDuVS8DE21zaYV+wnfua2wxNawD95qOc
3kH27y/gl1wNA+4PnE/LLTpird1GyvnknCsYFnlF4vLKG6uoRTF95TkZBgXB
UQ5sILiBFSd2qVOXycxTToaDEyeduGe9QUEgfz7gqZeU6+Roqay2hf9nXDUc
G1I0bW4++pYpMj16F3ETbk7aOmNO2MRBEjZGeUVaknY49EfFwSKFGkWdHlYR
R/bxZzvo+/Jg7fg+hPitpF6en657fFUKaGt8eJm2WJRxTXTQFDAcqQCS/Bmm
sOLVZss1qIo19BEpd5xHDG+M56x1hhTLQjFlKMn3eumuQMpHJ5vAqwFI91gf
caFzlQuEjq3HDmXqA7fnFEw46+IJPQmIPEFU8MTFuRcwGBw2irB/WT2lFjx7
aC1F5loYua3fpqGgY/DEBKWx02IeB155sqIZSZ70jf3gwCY0bk3dcU+Npaf3
DvZ+zdbdBT6QKfAWEaMZjMAYKW8RFdGS5Ky82gkF5LDABzaf8fV5A5X2DbfQ
NcwC0sdhb9BMkxZ7aHh6k5xF/KRCdqLTj+rZyI04+FdSsUUPz+MAdyV2a5tg
sMykOGfYg45QTBwNUzlRUUqbt2p/NlRlIBZ6TAJXfR4tw+7Bo6KNofibUP9x
9h38U2XXyFpoPJ6ZEQtTButp+k9WcKGb0eHY0WGVFkvk2oux0EFyfU3BrBJk
zE+q/RZ9AOTM7nwblY0ayWFvfzZ5oAchEZE1qVGR3uui4Qib4Htsv6qiQd0H
9meXRP+pG2ctfL1oO4P/YVsJ/NeQ+Ay7tsBWDQ7d9Zm6bxs9FoqkwIYGSCCE
ifStdSpuZ33KAQX3QFPLVbRYdwZtmx/7QvHCRyrUH6ol7JtYmnbMZuRPhonM
cU5xZUTzOLGmmQurYRlqcJ1f2X9Ace23qZV5FzZ4+QpTh5M7JEPoz3oe5RTg
sJn+t4MkGZn8Ok0e0ddNQNGBDyICaYpqJwepQEqKPoofg8IQlozK5L4TIHEZ
RNJlHAjDzlbPhgHRUJUS/TmhIcaPmCEK/9fqIck0sCIMzHjO3qPUqcLm7cnm
Ha62V0zhvTZ7gwtI0GkVY+ra8mvT4m8Oac6vzFVelB67uDem+ishiiERFn6t
eFjS0JqwQbeI/7bwXUqtCpxtGvU6as87oZKdjgDD0R532PZJWisY66cKK4U7
jLYfPhZErjHZuF7ASyxWxvFKASb9/XCF3WgP9XLf1U5Kd78XZ9a70hSNTYEs
biXTAaMdQjQdD/nPcWqLfwx1N48zfWjVLWJaG+nNT6QIbjJFjOIcYgt0i0G9
pInC4QvDlPUjQYb8Va/WIJdHUOjmBTzjsedZl4Qo/Iz1uC2VDWa253dd6YT2
pcC3yB3uaH1bAFQpXmmWqkvBo1/NtYvMrzDVPGqIfJu14YefF/h79t5YhVoO
sn8T/3bbNM5ksjwp6BdbLP3GwQFDvt/vxsO1DHRtHCiQ4mitX7rOtMlt+Y5w
IewUXMW8LN1nBacvYxvilhuvtm6/4o9w0vxKLxi4Sj822MeZxtFmkmZtz8qN
0zSeGjFgDmWnFWbD2qhi+utveMoNFiCmimySYTQMBGhIRkG4fujQUwp82mfS
KEZoSMAKihkKR3VdPmCdQMFINrCuAgD07cUX7+36pVTnwoISLXp5lPPsasqV
b3uiWiTWquLq3ZVmIeqnlwhPsmBT1hgi6YfYoT4xgxitZxhlp4+cFWjDI1at
Jau9YLXHLUgfot4Wx1iBB4+c7d/jrh9BPlv/aG2ACPrazWK2GmJv7aPk+wQ3
5RCNLrbCoRyonwf04Kttg4JHFHUB/lL9Buuu1tRLd8f2unW+cleCWOaYdNXl
p6H2D1v4acsCFANclIai93/8PVv4dX7UJh2Lv/07kY80l78Bin8C8NDPTTyI
aROhnYqJW8TqUAMQKad8mNabj+5NfU2mTWgIj8kCbY79BtPDA7PuK+Z4IBQF
9DvOLsVRyR1Wxx6Lz6QkKNMVOrWjL99HnrCIx988mrLIlEf0SefgyB+3i74L
CkFFMn6pf3+Jlwuc1UU9nTCNgm6+ShREpxiwGmIkdzotf0k6r4DTCwbO0CyY
tLB2RH/tMeDL/C+E0NshPoNbIviRIv6qfJPfjBFEjSNl5rIB0OPfq8jgWVsX
UsmfoXFntrZhhRTEicznaj8PnmVNtKcM4XhjLoIOhmgH/Y/UtLDX68bstq0m
2UADrj1Fijnu836KjumpvhOiSZpQoxGNoavb1AjucE3jMPuFSvVm/yH4uNbz
iF3r8AZ0Ys5BVN3TMdiPXzTmB0iKqUVkRpf29DK7B+hcP8cAQFnYeDaYuDkl
5wHePmK0CwbA1sKQLTEyhkUdExG2t1atyBFlvX6anMOb7J1uUwim0sJvC7w/
bGigOv1PhCP++eahCKfn7SfV2eyPS/oIJJeE/pUanqy8Ut6k4C/aNOYs+w3p
3BuVMt3BxZVS8clicHUSc1bqttj0Ul5ITfRW+coMOiLHc2b0KV4Ln8Derq8U
cCU8W3Onv7amc2Pq6gNIyIONsZw+0iXBhLA3Ua6UppMHPvbyshD/HpCafOGP
k8gm9VLREcyORD+Is7Gc7mfOWRoRrgzwl6xMgRyB3E20mlZw15otuKoVHdE3
fznwoWyzbCvMC8ACAkmoNqS4GNv06AiS1fyM59ONDylVIQ8PcB8C5/dA4OrS
6JSi8Q8kNI4w0pebj2dmK/HMJN0QyZ6XNduXnvPS9uA90sgOS0458DbUIIEC
3mX0CcrJQ/XnLL3MDJbB2sAUev7zYsMPdpBzfZoib+vRZKYSdnQLQDDXHX3F
4VmtlY4562nUy54m+U4vjdGoKcXLHCsFAZx40WIUYY3V8L7HRyW7paTXfvqf
Pe0luUalA4mFDxRZzJGwYz6RPc2yQrRp/PaKXUVM7hCOvmR3F67gAFT9KfBq
7oMKgF7ElEu3AjksAjq2SxF0YlRNtNG+BboshT0UvY5EscgQbGxR3qORQqar
/wxSC6I0nePXfJtwQMWV6s6GgiNb1pN1dmLrZFmyzO7E4Bh4EKBiplPfxu1v
7u9+q5XKLUDzg55HNx6Sjs/U+NtOtFk+rhCZtpt+hMXEHsbo6VRYmbuaSCvH
4JkguELv6SWQOPAF0JtxzixvUc46OIOG4jyTDHayxcSeJFu9W39oPY1WY5Ig
O8PPeTrRI9uQlTHpEvUmZeBK1yqqGWuCPiAfarNLaJf+9T6OMM2rqU7Rtsez
DMjJzfL2eRBgXAe29hJA5bgQ9OgdyEnMhifsmofKzQ9b/JVwF3Vlyspjx7UD
H1WsyKuU9eYfSgKjm7QeZHK0BGeIPyb+HvAUiQaC/cRYVuZdoa/1t7LGNFA7
SHRW5zd+e+nAyAuAyVsxDW+qHoetMwsy6ctJ8X8fowD1zOKWOFkOYJsnRMam
upflxfkiBmcDbP1gDwqreuHeFG6ciKLLmrIUrUqsprj6PUdFbYOSW6ttqGqS
M1wIfXj3iLxt3u/rLUbBK/fOY8gfz76+7H4UhmHlFdksRP4nJPK6quCGXn6/
xkberrGqPTSqOTuS3DRj7Ekv9R3C9NXwHdS+5iRX77kIoM42WVhFwUyOLJEC
UEWSogjDFAaMhw00kx61hLju5A8ejRDsjASxZpbZ0FYstrgM69wkr/shOwab
ymfL1JoGSntxAbSrwhfhcQP6rs+L1AwTKnwCQcS6+5pbkilB7Iv3BAwcTti+
nokEEo6FfKuC3ErscldgacYPJPBsYXbFZb70Ah4Db1L4f0nOCfjnTGrBd//t
uBiGv5SgCb0AoXE6Ee1Zd9R5xJ6IbWxosIBeX8a56caM3bJGU7C43W8R9s/j
cEsgkrw1szbbC21Fc81bOd3QCC/QExv2i6oPECvmx2UpWXtWUkwdOxPUHmsH
s3Q8S6e4zjTOswpcqbe1jj/56/IUZhr+cInDMn+TwL2wVEUjLRmPkYXWrfc1
tjrjK4Jf1XFtdqF3/MWjAx4rTMyjTnEQDePwSYw+PDG5znyh25Hge0obqRjS
Y2xtopRHa8LmtZUxfa/I75Zcd8v7rKi1sdhbH1DQeDdw5LczVB9A/nCwX98m
7FYBQl1RG1D9Kdn++mNWwfwMAkYukIiEQT9Lql5xQp1359ZAbzQhXOp1SJvn
MjEu3K12iwkJWiw7oRPLKGsAi2GIiVEzSYQgmy9mutEiSOCJiiWXGa+wouMp
fLkgXxuOKPcVtPJyoGSrXWzD5r7OtOZ87TwDqjLKkjoCHy3XCRsZ97G9Rd81
s8e+TraQ4rotY4nnTUHmn2966K1h3Hnx2dM/SnWs6Bcde6sao9vWQe+cVN/R
jdrnCr5WIBUQgO4OHdnVtjtWBO3LUbizom5/fKi8SnO5NZ2633MVuoBnTKhZ
bFPEaAsbahaaodwhjc/HZN9NrU5czbTbRp5pEgZpntMsoh9L31+yNoZqVqcy
gZYQ8ct83LvcGS8LZLOiyFYKfESVtJ1dMuJLjAy5fQOKnxxkNZwATadBeLFQ
IK4AbICNSnKe2LEByPR+ontASSeGem9zE5VOe3tCJ2YBdFUhIMCDdoGr4WR5
NisEEuvONVdVMol5NAeK1g7rnTlcJMrslZE3Av3Wag5tdgOE7b1gs/VnIsZq
KAPRtx9KwB6Y2CDi0yZcP1xOJbydKQCArEh5ttkQPILtOgY8Ld/qaaPrgf3n
MvGJYqsyZzaLt1jxOjmXrzdgeYPG5lEYcuoLpSz7M4zu3I01xa1shPYmVe4s
Y55Q0zj1b0BBA0QTffTvDdfMqCjrKOZuG7KWazyRdGgucD6sydQhifCAaJtN
Jkc3wOPeT+VMih8HghxTk8Ypg7SJxKqwzDRIG6hqInO72ffa97ZOJNTfQ25j
JncbWO9Xa/oGc8TDAbehZsdFpkQEev/7EdFEqDoNJSzUEcVgEfAsdWL1MG+7
pP+R0kSIr3jhGacMSqwfsJlFbig7OoEA8wUKEmE6fhXtq0S6isKH+EojlPPn
zYM5HSb4wZszMYu8VsGpjdNGhtKIw9SpZNvu+3ceTQfUIwXFjDq4FXU1RaT7
U9M/lQ+rrm36rAcJoUHNu4Pyl9C5//67yIIMLA2s83R7J/Q1P/PunMwOIqxE
8FMe/BsH/KQrjOweEKWk3KKtIU3D3Zemm8D1cCtZ825wf1S2vhz0nfQXfIVp
reLaWOjQqEcMIy69O8Xg2m0JCUFHb8gQYVeZKv2pQ7b2VT/VC1dRRHDkvPfX
M75PjPXKsyp/EB2m0AkgNtAWBjVGmxyhCM7xAxAMGuUwKA4Oket5uQuybfFG
MRsXJQxnKGjy4E4CXnjvVwHinK2/756/HT+FPBBYAkLIqL3Qb2p6UGSQiQdL
SGv/WP4sMo2pMc6blH62yicEtbsu56tB7qfshT8WlD+aNsOABj405G7jIaEO
468MEA07M7HncQBXXKiUyuiYdoRswG/SqXuZunZkhdndnUqxfqajg1G37GUF
AjlvN7zBynb2AKuuKxFj+UqtOhnKgvPLNbvXtPMlf2y1J/XlCmbRt+jUh5ep
dLwQWt6Aa88F+SEY/mjjhxUuWPzi83+dmrsuAZVA9WtdbzYz+ZSCC2TzY0pI
ghMawK5Xxs/di8DZ9Fsg5wid1xsFRYLKIbQ13wgzT0dLB7oJhQGchJvQZGlv
wZwcfPo4oS8+AE1HBIRbVRI3+VJPCTBRdENKh3pMKxgeG7yIO7OrL7EmLGqt
8qWS9Hxo6sYbL2F7AHGcsztlU6BcWPrQRCmvj0zZqBMBl9z6RLopCu64rZ8Q
hfa3wRBsXdT/hQACwFvY4DpPNwacV3Jde9Fo4MmNqDPy+dQXcu1Iqaica0U9
ZI5ERqCU5zVaZdixzwfrkHWo1ZY4bi+eU7dW8fTheuoFvLK+tk2i1pBI1ENs
xCKRsin1wJ6mIYfoHW7wBN2NG9BsOLgHfHYzhR3V/VFaV/eHQ/jgcFymGhvO
FWPZCR33NmZaP65KsXXKwpsN2Y4kVv6SI+JoAqCChOtmlW3XSs8sLfDAkm7m
ojvTdQnUlOQQ1ScZV+7ibkhGQG0nu+r5VOgFPkpZPWBFKQVJzY92Aoft8m7g
fAcYYffBffB2jJlHCAyd+hS+dV4X2/mQd8TDdWD05Se7TZd3D/BOyr9ewRsd
ZquRny6IucMx2A7rFDDWGE+O08k7PN4mpvWrrpKCT+eY06sjraTIwrazudZQ
uTt3vTqPTxloYldm4yzgonWoCb6fxXp403MrAIXeX8pDRwGv/dXwkXcYoX6U
ikH/Z0BhUQt8aLX+ZEh80ZLLa0rYtbZfsNWW59SceDsu7jtU3fM6enXp2Q4m
+cErCQoKPI0VvRICK0d9R5Mqd1q7TImkzhW6GHMvEbDplDZqGF3M2BkoMrgI
vgEJgebEx7Y/ZQDJQFDltIZJyfNiBvPc4YZ6tWXeS1/KyTNuwz0AZpKpPrvG
c9S7LhzQZ7t3popZ8uA1ODY3Ti+10kZ1ElLc+TzyYzsfbmsebfjB25NdDITk
BqK7pxSyfM48usy2738lGgLrG9VTQhubFlhEJ/AgHXcMKlLVp7ISK4d4OOMA
FOv+DeVHrnpoFfoj25bsLnixNzbPt7b+KGqHTJS7YOlXE/GMfsPCJlg3WDah
/ByIy+ozSTJ2rlem4mhj9InYmN29bdNXX9cJ7aU2TiDhrSljnhLAjG3nfYbY
mItMymrK+xuHAHV1I0D4QMXA0BFR844KE/AnocS/FRvhECPLDm4Fyiiw38At
aOUNENGlq107uv2b7bgGAm767uAV7U+JKDX64B8Ee1LQNQ4cIhT5AlXj1Hia
2r7XWm/UivYBiNjuQZmFqBcjtLwi+UUmcXuD2urG9qAB1GK06A7+keQTtcP5
UJURGZDr7d/SWVgS/Ysf+Q7vmx815aXfKOiKpP9rAJ11Nnc3+fI+bHvQ7QBq
K/tm4cV4MS2TkgYipD/tdCOacznVWBClsDqmfD4YI6Ivzz6oFXGFXecZdENt
SRMk4Z3leVg14V9pqo0snfzX3V46xZjsVIfaYPKaDD4Kjwn6VyR86BBD5MTS
OZy1KMllpIWp/XyumS08FsHr3uKuwW+GiAJNiBRbtVrTQbyVp6FtLMNWJdoj
2Giv76ZxlIddcj91pl2B7M9cF26LF6Yse8aRIOD47u/s6WM2rVnmuoPOauYE
E4mj01k+j53BpLlntvWOD0bF7TP+5RD9aCFZoaj/CysqJvG8IkggvFEO6fEO
TGjmgSfq6boFK6upoqKSEniZWK//9Bpq530Vvxill6zyxw/QkMaaTD6KdTDL
qQHjAA8sCMn/6b8C2eQSAB/XrmCbWPz65u/gxW3DrFl+vWNhhrO5tK7FyKbb
fHbYZZdK9IvfMa5r1DVmhUvJHP0iBF9+VJkE1Au7wAz1G9PGuDmx1/osxitG
RKzgKZSZknnd5zg2Sf6431zSjzajz6gcKjhv5E3P429uAfaIu74TlEGmToeL
+S25tAJhVmfrghfBHKa1JHtpYS5qfLvUvMALScVAcxtrBve9TrRkeOkBqW8t
kiOQHPWfHs3d0OzR25EG24KLJGQlyqlUUhQP9IXmUAl3HRiIjGHrMJcQtxg2
kZ5IGyKQj7N6erGAut8ykoUJXxkKz2OPqigHGvtV2jFC2kr+Y2CaqHqUwfIk
HwC45x+qpZT+pBcTLRxoYTUaEORRcLiQgaVLBu/Eub/711mpVJxBp1VVLwLg
Du+/W9yxEoTrQvKnlMWVHk7q1pYixuA0mZl18EjSmck6+v2d0zAC+Q+5nuyH
dzRK7g4BCMxLmrq0cziAIC52+vxnWYyAXScIJetsESkDueEwJhNrC65YS68G
hAWRYNdFRATT7eDKK/W40WIk2ECYMNxqIcq4GMJDHrxzkDEnT0Ay8bgZd81/
k0WIYYGEB2ux6tgwQSnlwXV1qkWXX63vXvED4r3eHSfsasQx67ay4IdMuwUa
U3jmBiLTOf9T4kcmwmlHQl8EciVnktKpKRRkfm+rnm7YZCS+E89ghPehPy+m
zOxImf32Xj88LoJsXVCnXxPsQmqRAnX4o8KlfV6u9BCcaywvTJyrl6mfFREe
CB077rKdRXxrCYyVuD/vD3yo8TY20PGY0MqyvXFyAEoWOMbel+iHlHphFjo/
jCebBmcOK0bE+htvqbacj5Z8b1yb2icaOgubrJCrNLN21xNtawS9YrfKAGJN
bgzzuYsrw+bDAjYfbUUyVVDyISjtmTtzQwUE719GC+o0SZ/YUlUn6I41rh3K
oOjfWO1XJ35RyPe0Y3O6sF0efZkdH35uxLOz/kHeXV6GtA1OxoKKjUZDfSe5
SlxkDoHL0DB0zxXyw2aQJKg+WlCRNc8KoLupk8ITTvif1bICWusgBPYu64EI
AF+WprBXYdCUKmu+eDjFcUI7hI2fpBjg+jrUXcfEP52Z3+kWmmvVE5ErOr4w
Gu0J/lkg1V/0txVcjHjdNdXcj7tjur+NMgRYUn7vmm6jIgws6KaYeAa+sa1u
sCxFfNiWYCmWMUzeUM6hd1sHOLJHMDVwHIB9t32xSRNqkm6IxxqmI0hLIuUz
s31OmR5bVaBzzXj3L6cAzSIW7iSe3I7qi/IvJqWO6QM85loVecK/5L333C9d
QmKEHcHLkk1M1bNeN0Set2vw0D5U/L6E35V/BBazl3+BEB3vvzV5BNciBvLs
Wkjx7wirc1VKNvpUkAbFpmxOltF2PMn8I9xiEZUbyQ8dNFFnHuR773oIhMEa
PwedbW9JfhbnSO8+Ef0nwmFMHBoCnmxO7oTkSu10EESKZ+Rw+EuwZLzdoTuJ
M8TpI5OopeP6ozFbNUPgHCQ5OORVo+z6Avx3dgLKX0tp59M50vxWlYhNTNC0
89fjrLzVhVpHjWh0uCwu/IdHpodvopif3//HbFAUcxgeGca54GLtmtpN8LW4
6/9HGAusrrxd3QIlZRlDekNjNwwxMxxE1x3F0DckO4RGMn7UsSmmnT4lnKzO
WRtuxNhxsGm5ZU+clWxsvIjTVo1aBCRJVH4B1dszFny9VyAAc7JYsZNPMqu1
8571A0kl48xe4HJBtKVUCEMaNxm3fYeCdQUFULkOSe8wUId1qxdoLeJ28kyN
AxYUGi1LdFKvgfdHKm6bLlbNqMzCLe/bpRjaKAkeNfDK3AHW9X2JW3+HGVLZ
V2iECcRtxDCMW2sDdZzq2zOIMfcMoT8YNwAKlNYUUY39+GrUASUW7X7jlgCH
rKP3X6PKUAelFrXnzQbyKXR/ckc0nQ+Fdu4G5yYveHOmAJxbWT48kFfJxOQD
FJOvFPDPeGDSMG5kAhRMRxawtB+FSU/d2cyQwZTKuKZBT1kXU1FLN8ePZPaE
I9HYRsqLAUxDvoPMCc/WWBAIFaY+/Phaby1/AutsWdZPhHJjzEWtLHOmwpP4
699Qi+Rre70Jti4uwHZiozWhj8svEaoamiNcDLz3Oft8IjGV27p7Ec59Z7cp
oTYlBGgnugZdOkUafX5WHtW0057bexwq2VL/9vxW9hcvFv7JC3mgyIOYESfr
bls8JrigtHQDzgs3aRBsPk1RKNxSnyzFuLcGqV2shZdlOZOYeXi7SkFA9v8V
Kd/ZBFHyudRlHYU9Uu8XLdlB+SGdWY1nVFUlj7SdVKtI6WsbYAoSlL/hZJfa
xzglULW7D2gB2NhuUVA2e3Qam7H7OH5XwuSXiEgotgDouc2605l7r60y4evf
Gp+jRyeMpLTCFICYQeX5jNGM4eWxBaaweq+KG4QqgSAAMgGJMvVCOzNPfTXh
wKFnp56lWO5S597BgN3DzQmv7Ym6ClGmUJNfzZJAjmBuUvq71ejMJEyhn0xx
XyHQksRNCZ3BeTq8BXfIUt7ivJkWp3hPf2F5wS6VmVI88nSMQkXviesSRhhb
YeQJsqBQGQmnepEVmrPgvejmB4H4k7u1N6ql9Edr20x0g0eWRt/yBgIhEloR
A4MFI0OCRXYQ0NjJw9YKzHWqJrE1DnZMXTaRS0KXDJRdLcWW75c0FaAFpnFr
J9TFSjr9V+WrrsvD9RKor5ryeMaaZNr5c/rVikf2287Po4Poxzp3YpSBOsk3
aRnm4x5XELx3OSX6pmtqcYYeE1zJDQWIEC2qO/XvAMhgNJwjo5zHzamJzm/n
h0CuoiAHYxxvMTyskQ+4AqN76dWhf2/vCG172ZjDAS8bYY8Iy/b+T9Qm6Kys
57QRAOudaN2FLwNSfbg3pTYJ7ufi8T1f5F8yxMeW+jlanBumvRdnzSt20g/B
V7e+3A76mNOhgVlC7r6NRVgdvN9QNJTKJtaIboY2wbAKDyuN+qCR+PA3m5XB
YGX9q/BWbXMNBdUn6Osj9ttGFBQon+SeDOsEWnJ5IUH/I6NMgVhk2SassJQI
Tin/lqP63HrUV8yFAc9Xl/Etsh3+u16RLxbzRnJJx3qJAeiljnCN7Tc0kmnE
8+vR5+vI3gMoen2f1ZsHOfKPaS/cp2dTArGlT1+j/8VZS64JPMgybr+4z7gh
pqRHgJBzJkaEE1pueRL4ZOgjAGO1xTAPJhFazpPElmYOvU5MyQsGxhhImjyY
+siHfnPQEI8cw2IQEe20x1jmhHwOJShurp+AcV1qHSCQfZhhX+6cgggOxeVG
OZqakr83BMlsb31PP09FmWWcCbSMvr6DEcjF08X8PVrreaVLUBcEAU0oQASp
GtbIHmHPB7EwzVT8yseNGxh1bF/aqiHpdppzjiDhEvepxtt1psyDcxHvV6Wz
VkeP08TbeFaN5CTsdnpXCoKhZO+vywyQ0f6i8W9K8ZGvsYt6++aVRRpXmTzx
U+4Cj8txI5lG1YrR58fSJjz+3MIDPVmA4rmRKpyBkTawd4ZfzxeY6625bhP4
l7nLRpF8Q84+CIhDBMP3sB9HAxjiaaHqhnN0L5v9nXOjv7Q5nf88+V3JY5Yv
LqTe29Aa2K4Vvlzg0WUItD7AUZtbkAOHZAgQ+CME+bEqLdLGmPWUAkpcIQ2K
TGPBNZL4NteY4ozeOjVonk86fqLCSBl0F8QfZABcwQIBpZR5rgCPz6ID2IJk
q0XzjF8P/iVbUMsgAb/Ujm4SICZlCoi0YHuocfv+6o1bbxPCmxvbQ+GyxspQ
ksct2JWhdENDnSN9MCC2QDeXIHxVOksxVy0cj8cY0WXaZjxMma2vUI2niBWC
yk+oriGVOg4zo8I2qOAjLdqRP1cJyKVMlliHsg+FIvaR7hVCt3GG7OJV666l
AKL1cK2y9VrQjlss0pXdMwh2IEygd7qlcytRMGapSZTk64mCY6cOCyw0mP7N
NkM9GbyIk2FajOtY/rruDHwDNb0Sls/jFpKRV56YYMXFFxmKJV+HUqrXyLtD
UrQAtY0G1R5D0iij8ZKxhXtLTYnJs1Nzz2bz+K3Be1DQvWuY24u16ewvW3dX
M1tGuJ2zwkyk+xxne0Vf2UGFQk1RiF+gmaSMqNZl6BOSL/88lZWyNAU0pwO2
n04XiNHfcMuQFyOIz7vDw8XQfWJ4FTr/JoBJwSG9N1p+R0ys8DyrMcLaKk5I
3HOPnOEbXEQOM3fPdMcImlsUHbUMv5j2x7lpzVrW6zQAM6Ge2T3G7lalpg3t
mPdQ6+i8OfKpe9ls2Wgd2UVEcYQIzwPNNzB8Kf5QV5Y58yxBDCcM4db9VpFN
56nVrkQEoYpfQwj+jfO/oYARhItexGbQyUm4pGsahytGimgvWZYD5UaALell
JPhFeSvmfZiRpJnauU/K8mAjldy+Mx2I7eTY61pQ9AzNbOIXaPdaE/I7XCT/
XkfySSsBxmtg40Q6nGHjDscEyP3RR097nWiUyXoitYhxQnPtCLQOrNN1F7sg
CuW4PAIVa5lMb2j4W2fkDPhOw8urHBUoojG2gaClWYEQQ0v+eDuyfAA+xELR
rx29zzfVKoOJLlTzayMIWzu4bFH6VrgN9bp12NfCjfU8BGKYNTGisx8L95q3
vYk8t7UBOHsSUujLajL9WaIJHI49GtLk/8pv1Rno41KmepbKZsq2WW74/4uk
AkmZ3vmaziCCuypVe9JxhN6Lu5geclaCLmIsyiaVqVwH8mvu6HeSwYydTOjs
RuikwsHZR4A6qmj8JdNmW0C8wUkwQszZyRH3rhp8n8+gzySVY/3hetlzbBCc
xUzeENvX9XMDYf+MybXlsoA7/PrIh8ilowytyvwxTUgfIl5nMmYIaqoLVq2f
NTrNBvi/8bKM+EXXEhnYKGTaPpgIXe9cMOipButUHjDXZwB1kEC+72u8LmHx
d5JfeBVnxq00ACUc7qThkp8xp2tmYD6yZ18E3KPN8/fZotw/E5VvQywaGEQI
vtomodccuvn0BtFK/3FXrUZMp+zXA8b39OJQikoE58eLWff2XrRDBTfxU46V
UqVqNwSUf8DUgE2uQo8cM5BXlaXnYRuy+KAS9AqAjhZ9aW1hjNmmxKRDMePU
x7XtYuKsxbXzXOci2qRBwKuzuzvZ5KAd7qso+Z1JJ6DjW+HeKB6a33wIFR80
M8NQScdbKMuMf549LhRK5gG5mWsgt1DOM7RQY1VIk+KI1+ieA8MXWPPIeUbj
s9D4IKsLPr6TaYrCKnTodlZfMnp0iiOaUNmAbr/Acuea/waGX7Gi9jAgW7+O
T9EYZoa3pBpvzAh2+QGkduVEd2AsTroGCjHkaBl9c21NJxS6v92L5OGDI25G
QPYAH+G9TVAc1UXDsSrUI1dJBx+iA2wler7tjMyU5avTFAOlslGMiPdQXYcK
x6IY9C5DrYboPOHNU/TqEruBB5+cc+uq+LQmF9GR3obp25TA20jah2itd2xR
VKpboxmKc3ZRXDl++UbqqxOLeTeDm0NsFkm9pls5KrbKUBQkLn3ZS0f0oFWB
Iz3FueaicgW+3pR5WE5wiTzSzOFxYAkS2JyFdcM86Uv11k6sGloycZIfJGRL
eE1yiw+a1mbS4jXScWbMiba3pwJaNQ9PTwl6GGdVKAuGwglvSUlytqGLBti1
47Qo4ycdM7gMRB99hiuTTiCA5g/z4Y7SVhQyGumM3jqDhMwaGQurvKmdxiWW
7D6FyRjAtFphr8Nby3xLqnzHK9k/sliMHhWiaaT46IlOB2I75whW58Pw36nA
2NSt7TPoamWKBbkM8JqCFDZZ157zM4DgBebGvX8lkggJxaDviDXWDfDoaeb7
zPdfIWoyJ5mYh+wyjSQGSI78m4u2s4ZDxFmXzH3U/vnNy2x/BooSi11+8XEg
9dC/ZaD97QvI5YnQ7CPqVICFhYr4/z9+6ugJok8WjpOCs7bLbLSEqqEXFWuQ
2X/s8CAfwKPrOwbrue6YZafmK1YDE/wyFOlUKu2TGYl1GFt9tTmt1ypiCVUq
GNDs6Vvsj+c6ETU0MwCN1/UHb2NtiSm1cXHJ+UbAiU4USjnrky7DgLW9ji5X
kHw8+/pHsLWs6qqKPcfmY++B8KMoBs0MPkfAwxzQoJdklTamkMSbUz8kgfa3
usqfBB1qhiUaSKZvhpwkAJTWYqt+iXyl4FemITLwbf+ssL5VhnHlu0FvY3XX
ZF1CqN5Hojn/dSXvIRE2eCV6MfrRMrIiw2+MdTd6ChUtU1zPumCk93lPlG62
E/fboXauZs8rEDwjoa+/F48JAHV4G8+S4tEx6ABo71EpDHCAMnzm02WPxXu7
tYiCV8EVuj6lj+/kY7sBiTpi3mpfFAvI+Nm3D/j1cEpNmIq81wBTyOvuEZPr
QJS5REQ7ZUCQOA8MqD6jrzGvHLD6HdhcF5OnIODXhhxt9OelKrE7GnPKT4qU
QV3ysFILmhCemOKL7pzRhsb75jyHKDVGaIF38+w+kR3QFz1tAtCABR10evg1
sU3vAC9n/bXWPf8MVs3WMZyf4k/bFpLDNYS5GK77/0fB0bI0CPAuKLxjXt+o
jIrya1LUvKbR07mitNZzmiYi/0DZAvMg3ehBfNm0xSDDm/ye16vRTzq2IzhU
FJDnf9cqKo7uT07NGhif3YsXXlEbdVbPXdrjqnKBZmqfFcYudp3MrWdE9icw
pFRX63uFxYYU+Jsl+0+mvo5RhjuUYJHtXy9wshB1SrzDYGmcKGnZFZjH4DAl
EyxdePZjPIBdDLnrylC34kr1WFnyF7d4NpcuPB7LzS5TMVbc1hPaPZ2HYKXh
BW9AtM3INXvNpt9s+Tj0IEe4zAywTAik/cVODk89tCGcNKs7Nl83FVqiWUfW
CicTqk7kAqBLjRG2CEfLtNGhuJSqoVGOoARo1eV2qAXgqHha3xWEO9Sr/IZP
gMXKc6uPwRPxapMGk1k1JxwkNZxQYSDAvI/d59gjFRBmrUC7cSbW7jCvPB/O
+Kv11pYJe9kYj3fk6+9dY1oa9Bsb0ULwsFEJmv9mkA8uZovb6OwrKHOx9q6v
ugk+xoevvEOL2cb7oMZ7dqFDf/pOOl4w4PUhit5Lptml42WqHZYlqaiOAqfo
Tm4hKtLJfkbn1A66HcymAqIPHe7qx57hefQX54q1Pp4TGJxnthExxylY/W9I
dptmeUUPlr7WIb8MRHcVL0GaE+ixlcOIMALztxQO4DM/TIfQTSy0TmPGa0Ol
LH7jHGzjJyBU21ONToQVWZJOzUMe0SxlbXUXRREW2gGke3uLDNMGfB+8OE6s
QSTnkR7m/EOUDHsbJ8TTR0LY14tjED6h/Gdo5O0dOO5GHdBkoa7jCr637Wmv
CBeNOKjaeX+RxxMOZkfm55u/blz6xKVJsIdlwouSbl/bG3DRduGc9iXr/1+A
qjBUXNNBUl1LPVGTxPBjVtJPJ6iZp2B41rGDycmn6sNhQ8B5i14JFHRzglb1
lLmM702ibEgY8FS1cqrl9m+sauuaRcIqwktMZrZ17REtEN5Qrv5rlr4fSRaH
VrngMElNA15tQhdjxGF6WxhLU930kzTbL0PzwzkW2bv2DKS+ckKlCP/SyOCy
b1UL2sV9AP880b9d/g0yDdmE6JBg7ZJsX5KTC1/vO5sDMCrRt1KEtqFUIJPk
h05QADJ96wS47kob8rkrTK0qnzbktrt3kluKA10RcS48xTNb+9PkIA2ffb1d
D9ey7D4rY6aZnPXVHNI4fLCx1EXjFs+ovsLzwpslj+mjmtgxP0iww/gFzFzd
Ghg0XqmpK4Rb1wvdeVgwVMlN/ACCOIeACJ76fu1mOcuevdQu4i95CB71F7eT
YwqpkROuyUpevALLPg8AOTOwib/uIbz4mj93KY7lwXdrQKXVMwXi1CV5bgOV
/sHIDJB6Z6nNHhDv2XMI/HCgCQwmA6fq13xaKrT5CGhDkMDDsm21hKUIsnok
LYiKEVrBYirS7JcjqwGED+ynLQ1SEcr9eYO/PqbikKipWR0kxbif6S6ihLDi
jv0zpuId3NO/MzyVtEMqGHHswbdf+ZDDFKwwX3HK+EQNNaj7sbbNOcXA2Xor
67PoF40bC9/n4eUk2jWqWsel5QB2W81RIxJb4jm6aOOVRGQyB6hEk2/l13PU
Xef3fSAC7SNN02EjD9Hf8gS7fa64r8rsZLTHiKCJSwqrXdyw4ayOuFfT23iq
8r268gpycB9TeXWltLiMioZV0ZEu836cKUstjK9ZNC3NuECgrQuj3yESfw4U
A8afXM1HJ0gBv8M6uxHy9rdfGlOYio5T7WZCTevOqQrHocVcgPnhLX6q/J9A
NtJf5VIe+F645wTrY7WNXJzs8K4VET6/eJDGT2yFb21rgo+D7mE6NMSdGWpV
1Jtsn/rFMuPdG/JJoBjZ8/Lj/vh0Vgiok6/wY+X1l22o4NWF8MQl5+6HY5wg
B7NlbT2ICdWTT5ZIsQQXyuk+sM70eVbxw4QVWv/p2IcpBKOZSIFbcQfTdWP9
HXFhjYLDpnUenJR3baNBT3O/at1YDl9+vFThlzPMdWAR+EbdlOqTd3PuQkW5
BB3dAcfzy+XQD5FkhZfH+3spCvFFNkRwAjZdr7Q3c4YDexXCxun//oKMMdv2
IDYSrp7FFR6D5zTPp722NJ3gzlnazos64hXsfuhcL97F2jITot5b05n62jDY
l2xeob/3dU/nKC79Bs0ZjfQ+G8G84njcs40KbeaKBWhN0yCPjAd1vq0XQFDo
q9nEjNIaMduehmbs/1CVKgM4M+O9snuynyAaYWfn7VsQsiLOvScJR4yCZH7y
TtdnwY+ez5LoqtAk+uDyFFEtHlL5p/cf+AmmtE5utU7/s0kPUYZSUTBqHFFu
GSl+JgIFNnFsQp6tBmkzNrw4qT2mHZRe9vuvcw4KWy2N2vMxoIXff6dPXNTO
TaiNf3+aT0zzFZH0Rf3VF68a8mAs2WLQhl5TGIIe0TcBgv2tBxwX5piIw0gk
UIAtd+t6hfeTmA4GmfbA5+PqMZNNBO4LC4MFvY/cW41E2ClJp124Q8TWUXVA
YF4KoATmKOvjl0T4La7z4BXWqVI9WjF/NcZ2dhsaGbbbUs+c6Qp+Z7ZR7y6P
wcsfEqYM9RpkT6IYsBoEI8HdPi7sOgRF8b7YeuwtoXHzuTNHdARiuB23bxf+
q3sSsvDCR3ojWMjA66lJ3bTojP79gzfB+l8G9eH3oaS7/rXvBicjXDqmcrh+
7xYPBhsqX+cQdaAILzQtdlu0nzTREwY1SD+l7ZsVd6m4e70B8oLUdc/1T7H0
CDgDfcsGgtUIu102uvpPyRWPTX6l7YcOs39BfarKR6/R4jBnzmetjXRdKZNm
DdNOobpWGEhjFVfGJPQLMWq4UK7pg9oNqv3NuSUwvSAAqJGixUhG5A90IRW2
pQHAxkRblraIQQW+pgRXw4L8YeuBjGHLjE2Xq3Bel8TaP+BquEanEjfEcTAS
f5uxd4Poh/anAaUbqtWN/sC9qrzZFHzMOJBBg1H4VcchahGDcPWsQQpivtXJ
352qqUd6yfyeZDZgD6rrYe81i2xwoBQ2Eu0b54Gs+ACz8/cu7mZ7oy5Ux4jt
0b5yOLO0U7nN2WmBd2m7xRInKYxhXGFcSbCqpYJjTV2d0froMKyYwda3EEFr
cJcgx0jaljYRChvb6phK80S6bCV5XVciTM1V2UGwZHwtoHeNIR/JAQuMixdr
Apmud0uZGHU6iQZzZTwIY1N6xpb1vyxyuwsIo2Uh7z78vXJ7XRqbiytnBxVX
ybn2bI6TSdDsSpW2+C2UOW9BBzRm9bKqvzg1HxR3rQt+i9nP4T907QNfhSaN
BONBEL9BN8o/aiU6HVsofzTO08Bg6k42dPtcuAs+58ZOoXyvWky7kwd8yjNY
HvwldkzYl+xUPOIdIpX2Ijj3dalistyThtOyWC7HubXpUcJnjV3ry2hqb1aM
NVtVla1NWh6u4EFFYP71ZEEO3d1odimPi/9MAtshrp5XobhWCv40l/PeSo8o
EQEiI9NMw3pcgouEPaRtuoW5JC/LvHLNTmIiB6v4Ha34qz+ZioHjJZ8vhbqE
J6xdUl4H46L9qyCKdNiWk81vg2LbrodqKj4F0qTIMz3PGZYWx0m7mjHjUjwE
rSIyxT97mJzUFdGwSYZuewJfVVhs7mH47Qa/zlIC9C6IFRe0vJ/5bNWlw+m0
qfZEic8y6PWZIrYL/uJKroriKJqm4ejGil6yEAm4C+S6R0lQPbmOoI0bPLcB
jPKCFvRBx/wkgcaQ9wOPe7MtLO5OpqI4kCbyEpplIoSC9ZV5kT1SCDp0FmMt
NGAIM1iXBE1EQAizxpS/jsUKS+IucWpHgcT5MRUq5Skv+aEXdZ7JagsDvlSU
RhsPDA0w2G5rpXJABH9KTtLFB4KcUZRNgUJW3365+OKHouAx3ojXZB+rpKeu
hAWCUI5gW/xmo6roC4quBmV1FOWjq8zyUfOYOr7XbxvqKuKxHTs3gXJxTu7D
lEDCZVgO5NKlyZwj1dpPvqY+TFT70CNiskejCfNxXW0Whnwd6PyFstnLBT1T
7/YngOH43jZKsDHYoc6fbABfb8guLsb1kLS9D3ze2kdCpx6jApz0S98oe/ok
XPcgSybZ8KTS6RNE/61SPdN6qGlpTZfrr+Qn+3S7SatdjWna7pyDxW4ONhUz
dB6krTdY5GPtwFJlt/WeWLK3qKVEJtRRbNdAnLUjziOeZ5OcO7GXE/zs0Bgy
lGtqI63h/0eYnMnSxnKhX1SSIP/5WJ25ZluvROTMwlbbs4SRvXoUIKj2QgwV
E/iv1UAIaw+hfkXsX2v6f4qbYTFdMpros+O2m1/yC2qjacYaL8M/walkF4JV
x7VZ/XCUtH4QG/FoaPnNi0W8lVKEcy+WrzToDmeNhpXIzxnUE7xT906RpckI
kzYSgBuEytl2naivTEgIbHd5BIwqFu14uGB4gg19+daZ/bV2Abdb/ZgLdgQv
/4uvVAN6BLpSmdHMDTKluhhhZpRBenui0IlcXkOT+c+Rc7O594/wHCRS/Lqe
X7Y1oaSFauahUXXUKP75/gPfFEuniUDoCzC/b2ESEWOJZpqHJti8+XGLDn5H
8MjFVLA8TZKCLXLIBdrwXAqIm3vz/7oAfTF7EZrNqvylCKSz/EhI3ZoTPonD
avl/BvbKEZ516iBl3V/km4ObLe/0iN9WpggpdSoiQp2ly0yDZ6ltnn/cy/sg
kBSj1pTjVuNe1JzTMr9DpoZdIJYlP0qYbxaM+1bkUN7Wub6NX9+DB+hRkjuf
BgrR9caxEr3uT4+DelCK7S9KZQz/WUP57IGbk50Y5kbMd1LFJkU1vRh8w1ug
CRre11uBruhtBeAc8jfW/aFqaqzV+uJaqPBoV0+Sn/TH4uA+TNgT9Q7WEy1O
yT6ldLDnYgBMAeEil4ib4HaOlgcCe1Ns7PPHprAyEvIQi4zS3QvSs1wwHfHN
nV+vmPI4tEnLeD6EbFvvawlTaZ05VvvUvL5Zxq7NoiN6m668HDpFBPMOBmNw
8/sNmk83+Lck2LfvbfwnnHHYf+jQSvqkC8Hi7JAWdJsrJoljybni3DoHpios
kuwHO1zGoZ58B4vspzJheO82gV8riu9wjvjpLMJ+A2LcVXR9BG81U7xAKqKj
5XmyoJSMuuDUjLMYZInrrSlsT4dwnj51TPuClVLt57OT6+dsYYj1WEVhmBaj
hqFWe7fQGCui4rPv73CCLX5IYplUYUsUdHmfkaSDTQf/KYvX0yeoONCLWrv2
2saADoYxN5/LT9D+mSe805AYsKqAZ7k7k+Rwy0+rJxEBZQy2tMbZzI2MmLzX
IEVe/sX/C5blXL9iTEYoTN3Ed+4IU2Q088WIH891fN/UGBdVtj2DHzmjko82
desy+2Y4FycXD8TqihpWi2xF3sPH70Ni/7Y04vqV2O/c1ekHOjg3TJQ7TCoI
4KDZIMyCk5wdpAjvwQBohoRGDrFhOjW4MWNSoQ8kh5qqa7Vgg1VfMVVkVnSC
EnZVeEGjDeQWZLb5jdM0LC4Z3h5ZG/lau15xfhQx1vauatDb7vvHwHJCWgwb
Rnbp/GqzYe4lYIb+Xm9iUJDooUQQQTOo4k6REDJ7paGV1zHqp1gcd9By5B76
x76YYOytodW/wTW/YLKaMSC6WXxI9jRoZTcptGnEOUGjzDM8T3U43HcoIJBg
aW7t6EW7eRm1J1kcumZuxg7sLHWxSkSMkEwqUqeDwP2YQP/NDjRP0V29a6cV
jCsaHZ5/1d1+Zc4fbDzkQMydnZrT1haTOvLgeMhe69uH4QCvkA9x8tBSycGe
0BsAasZC+MPaaI0nHi++pW5k0jOppZa/Ch6cdSbkU7tt9Jxf/xpPVvsoYePq
oFapIKScfVfoa5drmpQlmyXd/K8GtzkELDWoLDq6whNz3PzZAG1w5TaM3LmJ
72gtPWkhYHCtv6P83FYuMv2jaggM3TSHGxYS58/OsUWlZFOxeThCCivoub+/
3uhx9uLveTeDRcTG3oK7wGpJt11Z2L7LxWuftLFIUzPWaqH+2sVAmdAH+ZpP
3b/eziIuNHH8u4SyNAZ7gBOHEOaNqlJA6WKltuISORYmGVmac0YmbXBGx5DQ
ImQouq82VSRUjlZyPIutnMq6IsRm2oNEUfNWIEmJ6mTuPMvxO3unzt/YcTDg
uFktF60AhirOQSAbzatuXChW/iO0Qbo3ekvvdH28Oy323OhOYCQZ6vF7LrXO
a/6nmRCEZUZF+AWg4utEH/8RpgRpG1IwYFU527ky/IwDf1ZRIyq+2YN28TlH
bmhlqjkVD6Xj+lyW35Ah2SIVaVJJcBv2v/YxVVeF7Lg0ESPvRWhxCOwXM2pV
EUIaQZr7ywMd3RItwkSOVuHDp8O/rPAh1Jd3AdAurJjbZ4LSm8LNUwR0UoXM
f/dob+rkjsnmHpWlxoRUvbc/APQoDuQAw/a6pMAafhiWhCVZnEVcKGkEeOGl
sV641V00tN9CHrubIyzifMeswnePqyO+yWjc8SGi/4fGHnoCpPKHZmpG9jK5
Q9B4R8pWaqAm5NvS/rCVQFxntNC5E/Hoj3kqlzkZ8HAfmdHaWBEVcdtjHz4I
QV0w83B2siMJjAwefU6vYxM22ui1kUHZHkiiB4/SRhYxY8B719RtfJmx7DSa
hKUt4KC1yh6KOzF+seU/Ov/6CLjItnJq4ChKcVgiT3eiP5QmnEZFpoOUqUpb
QisVjgA8jhk+3gsAOoUVSuyeDXRgoRmv6tqCM1BVIq1sMs5ynroOut3Q7B+P
aUgeqE0G/PWWMi423nQAsx+4SrINo/lDyT5RoYN8g/irZN1tiaOOlRw2cEKa
uAXmcYnsW5+j/GGcHTJwjx6bVljMle57xYk7K/lvsBDlzPUM5ZWLhBquGXc8
mdZmfuQmsFagwpJXynBGlAshkhvQ7dC2Qq0iJ+NbYTUBek2iBaG3+NEjqtnl
Y5poi/fZeviblKQtEXuQ1uu6SItud1NDEsjR6x8WpGjivbU5fKdM/FXEsb7m
NswvM/KM/10HMom2QNuAN2k7/RzS841KOFyMmfMpA0W9WPgtMQl0Eyj18SPN
1IYGqLKDPiRgrld1k2KVU8thGTqFfHgmYiw59zngndOTUA1EYwLiLKNamajs
96obujwx2LEbBgv7Xv+yHllF5keZdIgDhYVU9atfYbqYhza2qyaQO9WKTIph
832DWwqcYkOLe2fn1zvEa29g0FEf+qEsqI/2kslW0Jlz7KiM+82CldQAx15C
kZTVFNZ/uo54LYbyfE18yK4ETGtfn1v2KNWes6bRz18Piv5towX1C7NXXajB
KCUIPYiWDSQ70l2dAHJ/JzND5iCKAcYLaVbSrSlWTugM7SpJlICEKWrsTl4k
+UEnHudCIwMyF7OUCQMrdYPVg5mHYFgqVJZ27HJBtVl6cmmD9054s88tRqlk
gI2ww9mS/OFSYJ7gmtmoGjoqiD/WDrKwxXvRcKBS+OJY03bqps7ox+Noi78v
BAjfWbkaQnBdGUOwLUpgwlSIzae19Mdf+iV/hRv3shi8D977aifjEROmfXYJ
I9Js58m6LHjFOgv9qq0oh+U8bLafs0A7RJWF4DUPaUp4xfWy62vGqefvWY//
K8+jTzKeFbRwqCh6Ok4KFbdYVFETmK+xx7GTtqYTtdvPbaRxhHTcq27UZ4lq
0/BSitFnNQnRUYq5+Pl5v/h4OSI4x74bx92GOBDmBXu5hmT3r7aHxm2+ZvLk
vhUIgs2BM1mtR5GnMDoPw3i7vR7fHbJmBv+LbngMj2JBjbqGbdDSM0AzSUta
9hQC2+yOEN6/DNmrZEJ8i8IAyAbsps2cvwHluf+Dusk9q2cqmd8cIEhDz7PC
+quN9wWPKRMQR5LQD0ZAgNbRsHuSM9ijKSMVUHym3rtGCkDhUExgxVbA7acr
Ndfd/AS7SRUyHszSlrN0WgNcVTLNFtAkcPLpt6/DKFGd7vWq+IcQU94LIeAc
/qzhEhlO5nK/JBn+0vnqXky8PCLbxEjwa9sNO0i/PZwkSjcSBmL5R6lvBGt9
mWlGfP7pOgGRVgLLBrFrxrp6JusJm+UsfArz9D0vE5zgT6XpU/5SaMyDZEH1
Ov/4yf/W3dqOiofE8CXmy8gd7LI6kf/jCk1SDC/Pjgk5XxZn3ygXmeLZM86V
83cpSHJKPe+eNpoDu28pvPhQn9dNMiUhYtwhEmW4Oc4/POWNbWRRnJY6oSTO
LPodXvXUuLDZZx/fqUp5apL6cEVTASNaVs902vbyGTl9mDhdg2OkBKHgbZxU
egykTPFNN2rikZQ090Ofy7ssrIwuU9oPImjDcAIs33Aa70yTAOaQkiFmWf4V
8opMPqobZqeMStHdSoQwK4EAsQACVOp6nNv9DY+JmMbOV20txNH0lx65nVnj
90MTyL6eRp2c+i5k8X4vORGljy+sZtJuRHJNQLSk3CjpNAnyKagAHPpmhKVM
uH8l97IQ0rROb1j4zV77PhzLQVQJJ2LNLok+cPyK7O1iD6s0J+CZl0v+FU0/
FpcwmmNfOwpp9BRNJpaijgvGRMgxae9WiAiOcxuPY16Pi/g++ACw11eLidCi
2ltGatjViTYsGyQp8gEWUFiAvy6DFAfv6wSylc0kuZ8E7HSoLWPt9k7fFxth
ceKi3yMZufCHWUpUCgpv4m4yf3LrknjNX/oEkvm1f+MMcf269l2Kk6Js4jSh
+MxVeM/yLGizjMLvssPG8D7cA4GN//3gZ5hEvVErxc2nXHUVuFfdXWa6XA/c
mf0+dWlh/YqSjmhFigGf2pRoPM7vgMPag9bPwX29gfcGTLabzNs2jK2NPmny
x/tDfrN79DKPcotkEPYRGRlkenLYvhdGu519Lc1zd5NkrcHB3Xixdy4OsU7p
3vjqzQgvTXcPRuxQEgLwbmCDVXX8f+5I6hwS7gm/2vfBfl0i7umt5QXTNvvy
HvLclGwrZmYhUarCeSXKvbduGOapN5DIMw4cNczA5sxGj3K02Ksop75o2Gj3
OSH8Fx9hKSFVm73uU1wHrQggHscJ/09VBp0ia2DdhRR//iLvVnzlkcKR3o6P
aKcXG7gS9MbxVV1eJ7Vdu0c/w+exwuB9SmMkvJAyUYii/6G7RXB2viTAoXsr
q3xKvk9f3Y4KODdRriWrdiO7+/Wk6FE92EhOpial6d+3jXNRtm2ki4EOX9CE
MgOR5kh+jIOq1G5ZjSB948g+FruHTLEu5tHRrp0RUQzTs5Vei2q5MlH2laG6
3xLGVDR4Q/Fn5Q6SyBKKauE94YeNbE5izBd0YnMTR/q4x0incZGtVHhM6nmq
LWK7U0bfh6JnH1kOBiwsXThgTODw0UJKJuqsAkyxxXM2Cd/rtAoOZXv+xrW9
akz4sT6lgqQs0+2JLJ2VbJ/CMOFGOOsXAOBBy0kkxba87hs6vQJQ6Y2ieeEO
yqe+KyZf3S7trpzbxKEygeA8f6ZIUEiEtgYz4f2eeWsjxXjmFzKAm1OkCBCV
/+mZ5RtMfQCdq3mmZWEdFpVkGECRhSiQ+I1Fv4JRcm9OQPaGp+96eBaZsNAf
mOeF/PYyMIWjlUS9zcMmwZStPdYWdADhzDbG12fSzXgwDKfR3OhXs7Rf03uf
lzH1QuJ7+tt43lKk1kJ6lfX5fHDAuHCyv3gELPtwOU8Xi0zq5ZwveIaAfTle
4mSVhLrz08ig8QNSlMLGJD+vHM+gtu3d1mC+zmpzyw/Fhjx+jsJRHsBEOET5
R/IzP+Hp0DlzU3z38dpKd7983pR39GCA8tJ/7UCeL//5pPRrLnVKorKp9moj
zaO3vjaOMe15FggfscmufqHUfUNzkdzrW/Nea9DafJfFPW3wtC1K5Fv+kXLu
CoWFGhTjoF5zoBSwGpQdlEi8b9vzhG3E14GmjvNmJiWg5zIwA6SJNXvaHORN
a8tv6hIesywAv1+h1xgrJ/+uo5zTERZlQGO9kOKBiqQYAH5EgZyXMqlo2ZiB
YPVAHD4txSKsKFBAQ1gqpNBiXxjRGMV4jzrvBTqTYnoF1qi8FVfaMtcl/w72
/qPDTWnLwxJ0fUyaXz+KZdglojJj4sl1bTHjTHEmkF7L8JFww5KD5P30yrHu
4KP8Q92viSrzcd/HeuglIOni7LAaYH80MNraKX8qh2oCtptw4OMTsHEKhnDO
G4nu6nSnjfj6Pbd0CmkNVxRGouVI14RMei1Te1l0PaAGoX+C2J1l6Of133At
R1rnUrbbQ7BiyMTRj3AJ2gmrEaQPcJDre5WbmDyrUGMBcpvG1qXdYHefP6aF
OYqID0bbF3SuccqfeQWOGVuu0KTMAT+hIrHxyYwwb7z9drfE/twkZ/2XEBH1
AuYz0fj9iPW+FSY5eg2ri/iCvYQugurvvWBHe4UaLTdXAmF9mMFTfnFoRfAf
HtbrPhQEj+oryOk1T5OD7OKEBeR+/xkIHpxAKr5D+AXC0EIqy956EeHz8683
e2rHem77FNoS77eqV23ERtaTfGfIdqscwEbS8hxBLDdPnsmMZB7UH6zF6IKE
/eVD3o/F1HUre/iKW+xCiIy3baP1X8OjAlng1r3E3wB0hes2pyShPpkSScdK
3w/cB4ex7L3Xu/RziEcMWa83dFDVhj4tUK05US86TSMA2kiWyI7dTjSpAgbu
wXwDOwMsVQCJvJZlDsaburQ9HZ2nnBFUES8/952iuPoGT1UPRtzEm0MwkLqO
6UOFv+XhKrUHPKhzXZcrSnYotEv/pefGS1O4ZsZc9RzolH+GDdgoi05O8ZKE
I+fEYPUPDVwIwdy3AIekRRUSDG3wxnPsPfz2J5/vj9JCWyM6RuB9lNmEH+nq
gduXUJR5boRxuNh0rbBmycVdynIZ/crHrWXVM2Lqv226BL6/xCo7ZbwutqV3
xRymOWtWD2BcD1mN3nAYcxAATJDDDnDuOkoAyCri5y49G0dTc0E9SV32KxyO
qbOqsOwh5UVvKd5uaKJKqtdFdYPh87iRZ+6mITsdF6JvVluhPlfRyqyz+mRa
VwmFLsJb+9oOTbJXMPvXqnbetSOs65Co7eGYjPdSqYs8mBow9KGDYzXYGBfj
42qX0R2BGI25GqzC8ZRXxCaGHCIIlxYR8Tzx/FbkcnQuvKIYkuMCiICT75lx
IsuZxFCQnjZsiHVO6DRjtjsX79f9GmRKEfvQysnM956W2JTHkMYK5HLgd3Yq
zylR5/GFU2OGPfQ/RVTdQT95OzTjD5vQ/LET/ZnCn599Z9MKIlLOF68k+i9B
x5Z1Q1enTDKEaa/3jlCERWNj2Iotwf2FVblneB0uO6gGjoRGkDaIDDVs5700
2zL2sEExpjKa9T6XoBja2zSNvD6MGJLEEcctWpC4/bzUConD3WTEa5hXpEt+
yQ/I06233ULlmPE1Z8pk97U5F4eo2RohPz5Jkl3eBxnB5N1gpb/VILGL0LFs
cJJEz+IIPan+mFBzKsHsVVZZXaLXUzjx+s49lTVDuA/mQUWkYj5dygID55fN
rn6t8g12qLSNuM/TlpLE7qcitKgWKDYjauvzkrvY6R0TpOJ4qxK+dTFxT1yi
ctUH3vl6PXhey0jB3c4Gj/D0HR9rdDFzQpY28oB8LQvEEeuyGd+S5xKopwzW
uxSFDBQKNC9x+C1il7beDNRMA/KLoqwUzX+6bEmXoVoMzlAUpm64lVDHAj8o
sX0+up5CKbNQlF1D5uda29e1au9gCITrAsr8vJtIINIF54c7Bk/P70tjkBWh
P9W9YQfanELarrPJTaBs0JuxcMKyWiOYWjfd5WknLoLAWV7k6Un9VZ8sUst5
QRcM79PoNngu+Gf68V9QuZxHeCOdBpjIKn1B1YjLAheyjx0rs4JTZt404yYt
ecom/WJwToAU6gQCc7MUsDZu0A9QSJ6J9kWuPZwR4Oivxj5+4u7UWoUGmdlU
9CSM4KjA48j7I338oYQgN6ZQC8f90LDmNGuvjnueTrv7mbTSftYyWybCOP54
LGeWu0cufDWP3HGRM63FvSqztlqEI1aULzDz7UnET/cNCjoKwIePImsEoeMQ
YetmYSAylDumVZdz9kjM69uphcEQ9/oSL793ev2+i7UprdvrnN6Y1Z30srbL
UXpqZnR+XVrBfORhF7cK8L7DYxWzj2WpZ/d0BXAZS3Yvm3GtUGBqcc1/H3Ru
6acQJcdNDp8Ns9/8lXq8uW/ED6wIkGGuYiXTFBmA+2R5yvyfb1nFmfdbEhmz
J1CO34iKUxv4Vrc1/qUY77oFcR0LJScuEcdRxa/TEaBUWoAMOLOCKB7MJ4nk
ka31Upn6HYPPrjOEvgHYCncZG8h48G8TlncQEYM1CNQrTsyyqrI7BSgWSilL
MBYwskIuhalHKkP95hLxHx3K3HW4C6VJqc7mGLmK2rjA2o+bV/yeHiP3f0uS
xRHj0TgS3rEvZQs6MrUsr3/efffcTNwuvFDEgxoA172Bt0r4aFJ5U9Wk+jsg
qYe2kASe+5QWqtoaY0wo77auAf75lFB13bB2sfNMJ9PwlLPJ+f5ivirPDK2o
rrsSsBMqK8VM3c1aOmyzTBPqg/dWrpkWpEUMsM4NdTRt6AZRGekzRtg4Wgck
YUtW0D2kWI1d0tgxLU5fOSdWPKSGZfwVo8ZA5cnjSlRInisTGJ7xKTe4rAKX
traDM/pQCCSIaqbpdtA30qil9fce9cqBEZJnadECmiY0fCdxV8HasOEIljd4
p9i3v2vmzKp0kOs2Gjaq+WtczeNduqx0hN+oEBQYYPne0SqCt/PfP4XGYa7/
aGG1JFSXoXxonQ4u9MJz1IVoHT5K8oKJUT6TL6V83Ny1rX3UOBasZyHcdVlA
E8KfW+u10W2nOKizb8niIHcxrhzr3FHH2UsxhkB45BMJfRIYehYr/DsrIGlh
6LWDsRmzHe7cwRLDIuW+kgiEP6obvdMgqX4Ymvwe4XqoHxPvjTJjF+LwmA1i
+Yfnuz7OFVLld1VIf5mM0pKNT/PKvsCuvc3WkD+ltUqpoUfNxphllfASJikb
fe92qhINxCxZ1HNZMYfx/+HcviNcC/pwkVmdmgHCNUPhvJO2oxCeNNRgygHl
TwLQ7VoVQROlGVDR+1/DcBLZFgPKMeHkXAleoPwhWAYFKvW5Up4M5DC+SUIH
s/pG4zShdLugt/7CMIj6utTI/ppZHqgdcwWsfmuTOdnuTVMAob4n/gUU5Xjd
Eo8bmqzepsIfr8FU6yPTITrDDEAR0jnArRwtILRCTbPA99QrfRmy4wFGxyOb
gFYdqRiLuC5RsvIZEvLHO2fYQYxciRDQoTddu5prQE5lgrVivyzuss6IZ5ku
CEab8gstf4qBIg5NVcKnQ/OIwlPFM3mWw1Z33abF6SZOqoY2UpKyCNHdgDF8
8tOHitekUjYYal1yMMujAKH8aOdh/yMw7ceefcuPYXNt2ZQ5IICoaP5QQjCD
MbBFzgVQEeWQEDA1jJWWaMDfFxRB7OCc8BZBlTsd3gEWjmCGUqR3akKpcv/p
VaYUPyCuHRpJwGhL8+auAa2iz8lRPwGaG8rJJzYFCV8W+DNMbpz8MPoZeC5F
VO+LyTXZKtxLDd86kfQVi1qdCNJEACUGAdX927zm6uo4uwaRaepe0AokVyKz
iE+0oU7vE5fkhlGYNyJ+2s3Ybs1YzMzUVbjC2DhjgBD7BQ21X+fHDl3RGegA
LV7Ldha+IsSoAP9w0uNkh7Xc5g2nNUKRuTxRO/vb0E57KvksMvxPHZIl775i
ycy8RUd+enSyLBNYWb3pWeStnP9e5dT1Iayu6qjiPduALa2BPSW1DIg+Nt32
vaAeRUaBDv1KCyDeL/M79iyLDWIT/37rQ7FrQ1OEtLIHmQRSsw7Eq18TW8d5
KzYcBsCMAF6+gbURS8P75aF6x5N9GShqeXM5IeUPJCDFIXttzb7r9hKR696d
aCRHuGA34HduIwpEUOxTPMmAp3U1pjcQhJjT0VVhoY2AvMtxl0zWqvv16Yg2
LSMys76O/ABBqTklJzVXgjARqh3/ojx0J0pwkL2z3beINhq4zfIZW//5Oy03
3AV3aJsoMz9Ve04/I75eiB5SKBO/Z48XbWHy5F43a7K7an3LnaDWvLRxv6rK
lBDTNYF3hPAvR7R4Adp9GeMaXqmGxtqX30Jh7TfSqxn8+59gm7takd6Y2PrX
02Id9YbN+HNhuFcx162V8yE743ZIek8Rtda2VwcJzDvVTK6vtnVUj5Br6Q7s
ENC1JDku+glNITtGbc5sKUFO0utUIQk0dEOzPR+NqV46daaSKucnb4fw2guE
Pd401GwO1zZhClbGqJQhQNFm3ZVGHyvwxgKTb0w0c9FNP3ZSgryjOkUb2cp4
jfuvSmaHxrGiOzk+T/f3O1hFaqCFyXMbFjIwJkeAcQos4eHoyKqUuDQGRGFJ
oWr/7k1O+1lOVxJd4KMcikxxR8Y3VFIdeCSdmCKkb4TitJBPbu0Ll6h/fSUx
tqG9dAGTMXbxHjqUcB48/etDrySC3hIwCg1YpraTUiQIlJcfUZSJM+liOPek
hVfA6NWRAqmQcWYA2go7OvZ/2T9CitNJ3pZxre/LsF0OHfGZ+He6stRSVFJJ
gUSnbHcoxfP2HpdxGpRLByD/y6zaiwIl7osKzzFP6MFcEswbqSq1Ebc+1J4Q
LFDz9c+VUe+UGrH5qAPvRi2JF+0SNO9drKVWB+WCrDfCYlV4BWdT/D7RODXP
ASV97xJCLjtjg6nA1gLgd0gOdGiFllSHxEfvO5v7q16jWfN4zibyzGqyfO3D
G79+u7rLAtXF+O/XOn82WkjpOXwjFFpnuEBzdI74mxorsb05/cxGu6i1WHqn
vrE87ceP3Ws5Db+eYUos9DJwoQg6KQYhEzEO9DJZ+SGFuLyYDr4lYZvBwbzQ
IBWkSHKhrq9Er3rVqs5/jWDKdd7ZTSds2A1RJDrxsA2ndTUpKG2ScX1TXCse
plQ3GzpufwcIqB/UncBWRirXnQGIQ9Of0qZpJhifM4RPdVOR9bEXK6SbfU35
tLN3ZrSqaAInBntaxF3gu9FeOW5dmV4iGZzXXTm+rR/nghxP9YAVFLGSsCDA
8qwgLs2+n7KpBNSFffed8xfCOSoKYsU4MbjwkIt7r3fmOTYle0IU0VvrfE0I
ddXCQ7uY9KiVbwannmuNTtsH/s1vd5rBUiqJ1Qo3hDKIqt6xemcxTPT57aD0
MY89Fh3M55EScGvDfkfB6NGvcsopHuBB57Gdrgd9D+S1g0uh/5creewt8Lue
gosKAYrnTutuuMKvJwNzTkFTY+RN1S65NOnyw5lWRH8ROnfSKuj47YGN1Gl0
f4yb/7/jHdteheyrJxysdh9a3DQp6GuGG6bh6tFvVIB+ijJE3eemSjBYXLj3
UXK0/B56DrUBJ4Ey1WCBR45xRDMcdzsIDJfao40XLlcHb+7/MfNlt9aSdu+r
iZr2CRdRNP+NPC83OYy8xeDRMeg+wbgrFygq25PXzHrgQiBoFJVhtp/qOCrE
w/vO/xUIBJzkRp+nRtCMTIKWmcdkzGnU2BhXGVUB8G/BNR6XuEXP1pNOEpAc
pZDm9rq3aPqgrwen1zbCNMhSQBIemwO7Yhn6eHk/tgZF12H3Bq/IZ1vJx5Zy
Lb4tOeCNGSio5o6jXHl44IqF22odH3QJ6w6H3/sFyTrUtOMG5e9OqlkbWOYm
iHZFgEa9fwFk+2VHx8RlMkGTpOI7qhDQ1qhzNiuh3noy1l00AsWvCOxpvGGs
V0JX5BF3W9fgZA4/Q7kY/uDWHvmjI3pM+gnU3E1lmIc8Mb5mD+/w0oXWuYUr
ogi9nRbq92EAH8i+GWWCc6Mifkjar6CSulHmN9DxpFTgBNWGx4QbznR7wcog
uZPC/QbpQCZLK3nZmK9REMC62se923mh2kPzEX2bP27vy3uzgpLFsbTT3zD9
5o/Pm1ZjVGSHmIHn0Cn1YhyRvt2Q2hrggrSCpDwZGroHy4eppuX9fs/BwSGp
gMbXS95HaT2WYoVTlOvQKQwBXW5jmY98F5Kr3ntQa8vbDrPSt/4nAwJhqjKr
1YGeEENg7TE4UQK1g8NOqHnbT5uc+yGyXqkYY3pnLH1LrCcXPGyJ0ZYUZo4V
Q5t0cCXD/OAgPoP14CIeeJcyCt7eDe9vqFuGZjmOrl6gNWAXWElyTNyBL4kJ
qOfi1PhH/eXAd+0OynIS3SnzAlZFotEJ+DUKueGVrp9yG2/iI5QXuf4418QT
DPxda7ryEhTRHaTgmUnqObJ/ma5HD6E0+DO+HOIoxESfma/9SJ+SIG5ThEM8
Bmurr0G741s7BK7+XRGEXq0PkOLVq5LmFPxX5NXrb3mQxvpnvKygsfMxkzV3
XtkARwrDEfQkcgWTVl65z+rwvmuHsZC8ug4b0lsOWcLWXRt+hGIlodIcg0pI
qpLx4pggT59tkUiWo7i8CGyakWkCFsV2Dbzm5tgps7yKDLfw0VbsSeEaLpnU
WI9r/ixoA9aujnpxHHKqTHPtx1xkan40NQkOm7NnTBghmgSuD0rr9Gds+HES
/OIoHHWxvd9IYZO0E7MkLdOl8TtPwqRTtGVHwthtkmNVQBT78CKOmG5pgFD3
beWhCd1i3lzEaLx83FkWAgFfu0IZwK+qI2WQrDTVoQhG9czIL9KfBWC4mUTq
xsNtLay9m8L3dTR+GZ4XcayTNv3UAGC1N/VUCm01OskPtmrqGwysRytcicrD
rLsXK0ofXh+YSmX0ljj3gKCDbRCWJvZ/OO8k4/8/0Pma975MRdl+lVS5Fy6y
KgOA85gpZbNdTXoUfC0A7YrSgV1eah3Gg1fUsjkXfr1TtUNebKtE3Jopz33V
pOmHbKdCClLQQfLELMcZ2swY57oTVBui0IH99Q1Z8z+Ch/oUR5E8g0ypHZw2
w6M8FQLlPUpPa763LAbF5SepYHbSU+3ZbuZ165VL2LKroU7cwh95w7iqjmD7
YJ89L/oA3Bd0P/GQYdu4caK2OF8+QNLJ5kvgXnb4iS0Cyz8udUkF9Iq/DNlB
OnuOXUhorjPZwHj8LYrLp3S1/+PjIMIPmIt3SKXFmBbM0TbYddro8GNXsE1T
zdueU2AYI8TNm0y4SKbkxcwFoWQ+noXvhjdhYRM5CaUXZHqJlsawns+IIrch
OBAnwbsPtnTITae1rt3xk2rnOB9eooHZ7BY3g3WsENVGN7ja+g2rTWH+s9CZ
zXwx89pM4THcymbca944Rskz+Vb8mnmAzmRpH77QaXKCE4zsKGg/JVjeBjY+
bbZaNmDM1dJgMX4iib7hRwS6qqDQgrkugzrHzjUkD0CWPyKrBD9k/7p8kpSx
+5s9yqUExPuCynz2diG60zJ8p5oD2pZpypFmQaWRkb5RVx1Q99t3CaOE8yvd
7JVugSRbZFU6top5noNUNf7a3EkYhx5V9N/fuUXycSH392QeFqiqGfK5kMzT
YCB8PPiD2ONblcQWwcqxGZO7N+fn1/5EVriG/HMOeUJrhEu55rXgK330S3DM
N81diPLFhGcLTINwe0OTfkQ5u7BhAd+xJUayaNT3w/tiE9tTi6rT1lyjL4t7
aMOv2HCi6O65hzonDofWWDaEht4NQ8zfavkVNF2YQNavkE3X7mUCdrR0pkUC
71ERbxQFn56eJCFdrhQmATNGn+DpmWnVVXAbZAGi6UC+pWn1BU2MOtn4B4Bw
StGkxc4BsD5661ahb5Wuevp8pobLGOI+ZcL33Gs3a7M4eDj3u2ZIHgS0H08h
xW8syHM3u3AmuCFQjcKd0V+5A6IF9v7GXbVgZ6ejc9BRkqWvwu8KiAqOsP/6
6tvhs2aT8tCEcpxsz8bumskq1sVJPTomSxerGddOpAyHinsiT6IhDgVZPHV7
5LERMLUPpLm/GiuUP+nelcp7TMnhh/kD0irsY3//xx93mRxpFjKD8BUvLg2M
bjuCKAJZWqhu237kPrvIf992Q/ak7UHi3jSiGFWHNKNtqtE6GqzhQI+UObhx
DnlF21RUW8fkjx5NGKONRK6wZCu9rF/WWSghvcpcXQyzr9o4yZwm6pEwLWqI
V/HIYFaC9Bo7n0G/vhqV3WmhLpqd6VJJOAFBPF44/pqAS4rEv+1U8OvZ3SAq
BQ/e3V0Bjkstdyck65MN6+hm5IAVjgrBrmi8St4vQuwaI1ez9DQnci/zvZd/
6Ny9H7QkneCYHAW4RTXj0v6G+l72AgJc0YiShiiVz/cvCLUbu3KrqruLxtED
WB7jet18tE6ZIVsedgxeyI5FsQu2B3BiBbk9G2EcnrFAIAo9LgjcL7uZaAXt
Cb9TrH87W5ajSgXzMhVdFKLJdFJEq1pNHsdhdJ90aGMwN+/ulgFY8h8HFGqu
sN67foa0ZT27+Sh0ExpZmtoG8atXQYfuGPjK0rO766+DqazgOMsv4xqv+UNf
RHTcvKQ+he2U9sV35m/hKJpCVBn5BU3uN3IumQm5p5/WKvV0Cg6NrYDEB7Ym
BeOi63irEnCoSEIrkqmftI9iGwuuaVN3HZMFyLTKa4TvM6hWnN2Had1uqqv5
6rqW0biU2uJwZdq7AD/QP6yJdOpdxGyrtBZhIJi02lsY900htAreoDcjxUB+
t7Rf/RXVnxSzMMQGtGUwmnr885wlHirFvIDeBsyGG+08tRpZvppC/mqEQIv2
nm4aOLjR4lXiTx8kwTSP72HzcDrNhXuFxctXZImUBfldGTD7AsvHvxl61Tpy
lEmYQeIypTLCQaA2kiSQcQZxgxS9aZsJv8RlyfhROVN4wQbcMcvHyat0K8Gx
AIqfibpSp2qNnnhpbUsz/oCbza09Qe17opChAXO7vqcv16Ja/MyzEYks8mTI
rG9InavWHf/4ghibCJh4MDPWOsVvP2aVO8c2Z5q4SNqNQB/4t9zsXyd8MQpL
ETMeYjMBWdqzTZ7Rej05+xEC0zEVvn6qF2kvTxSDX3Gcomr3D7jZeqdDulxb
8cGd5yYZ7FhEkMx3H54GB9H1ap+RfiSxuPymKRWtV3peC6ys7ZGQQU3TtFVn
D3rLP5JHBQ31xkXaxMSknbXmr3Q+1aVXbs4TwAP6Yjky3jWoBB0JFT07FCDr
9ONYcu5Sfz0fGvTQBtgJ8ikRlsPFQ7mz1W9Oas9Q5X9acUXfUCT3eWGwVzVu
vTdm9//Eyd4cVJ8Fq3RM4er4UCP/iVg0ylYg3HQXBO8j5InPsKSKFaYil4Ai
kFj0yzq7VSopo31nB1AufgV+r586ax1mt+dzIhWQLRTv/09agmKQhMjmFhAM
E7KUORXdDP/AE9OgNlw5hm6LfdXlTt12OP6SMTLTERP0VN3d4GnLqLBam0c8
zMD30wzFJNE8d7/ob/Awk0jvWDxJl4kerDvTFq0gqrUHDTgN8djb5d6Dhxxm
DEfHtGg1Im4g46Okz7qLOX7diD6Z1F1T8e6PfOEU0inrzA1TIvIbzgapQvRs
TWN4imhekARUZkpa+JPYrd9q4yUMiESGjOvjZHk3MLsufie69eReOXdNP0JB
pLiHnWq23TF5l6CtnkPOL1G5uDVsAUHEmKA9xcu9PKqxzYN/Uayi/mKOZuvB
Nzc1FhXCjWS522pqxRJX43LpgKiooYLFyeYvSUbAFpoQTPCLMZ3R4aWk9HW7
HBWBrMF/YgLyTITo1dJPSgacfQyFvP3KCGCd6QYWXxolbD3hAy3qVcir+9Uo
p89PX3/NgUE5c6t1Sp9bZPeUI1Xw3sGodcKy3itTny27gO6lCYaTEM9czcCX
50xAvmsdQTeQkOK8G/ni/DIhxF/sPUbomj7YODWockj0GhaulQcsm9dVNgq/
dqQi9WLQB10q5inJ4EWl5KVB06J2X7yBk8rwz2X/VGn6yQQdvZd6fqWBZrfS
7RRKknkYpKFXwActXdaA2mfLpmVu9UJi+//HjQSqgdoVdyXSHGQBIugDgXf0
pkqSn6Apb7qBKz1PEEg4uHa7hHaqMkCp3s8+/Ndn2PJsOvsxTq27rH+eDHv2
GpoBcISfrUxR6P77bzC7XRIH9k44vYtqkR37EvGHY2gAAsMS5znzcnPeXRWk
ibX3Ey8II+5ogbHaSQBQlw1tZ5/ep93I/pbZB82cdXUDunEV/Q9EZIAwCsau
5khQNGI7ltoiDelxqZ5I87XO4eyhgzNya2m9u+ldlpZt0CI9cVNEGaHkhzBp
H9oKq6D8l3Fb9cLIe0EtkspDdFjoJrkCC5mJrzmFCPzGTpAKMiewcrehh/3/
NNfwbRsUzppk5zOO3MMlNf5pj17/6aWpFRw82mRqCcNcEdMMeURoOwQfM28N
OPRVVSGMpbEF8MbnHakr4hkGcPsN+T8j/9SCcx45zeqXo7wI8kDrjumYn7bJ
+sFtWIN0H5dKW5EvHRWuhZS/+8kjoFLK6RIIZPYdEVU2VItbaHPIvCdayPZZ
B46Ille6KQuU1lZODdIws/XI0rgdWtDOiKtEkRjcIQyDgtN3iBx14N44ppZq
IBzIi4P8IRcZZA9C2HOGpzLSJ/m1Z3fMp4BW6DM8DvfYeHbMXEtvO/gWCoTD
XNOWMJOJgysY4vaJNVGyMape3rH4XZpKk/jzZSPz1bqJ868wvV36Fr1fh7tW
KYG9XYWfsjenIb/tSVGXM8jlpFMZ+Mbfw0RHt8T2fiATyXn50o86TdAlxyFw
hOJ0VxPeVkmzbc3ZRWArBXXoFDdRkXfdv5/ezufdALBiVdJoNY5f4XAw9m6B
bZ206V01P4nCOH2LiKkJVw1Qte+DEi46AXo5F4PWPRBGVSNwaObM+KEEcJxC
hDl03b9cDEWKhvIxRwJkplthLXSk4+UhMh2zDTflKC5EBwqJY7INsi0nWxyo
Gmdxtq7fCWH0BBs8Ht+5tjLS5lRUxwD/HaYfZpel9gN1lyb4HWr2EFlw+2zb
BJleft0cNAVElypXTQahpJJT5Hih8WAp97v/Lnb1DHKDCNhp45PrO03vs8fy
sR7DWc14R5eGq6y6AQWX1ToI3PoZkRN58HkOV+H4+0SGN/4b2Jdj065AqdCi
zehQYOnYH0u/3y9SLnMOi2DQBGhXJ+lM7KijzXbaisyZC3O3l4cvRPbsI6WS
SRVRQzuv3v3M+JMTkpEjYH5lK4kJ/oPApsFbM8XLwNt0wTd2wTBjvOWetAEn
uhdWCgA+IqHT5oGQfLqqDNOHsM6/Vnc7/FFRzmBdfzL3roA2yQx4uaraY6kD
gTyUxfBb3UpQCIREQ3op6jsHVxAF/OcGERyN+Kvr46/x4YjQyJ3p2OiVEuhw
qVWgqKGaadchsgcjWwBTZNQIcroS0rEjjtIa4WPz7W+Wr2Xsq9R7wfYifh5L
Yu9syH5+sp62L1AIDsTRXb9X5ecfHWYTZeJocMmEZZcbH8aVDhWGVIHlroN+
uWT9GLmFk5Qk0pyiBr64OLejwLDy5CYLWGYs/7SAZKyXNtGv3iZDbpguLD0H
CWbp/cbdBx0/s9F1UWR8ttMMRTgMzmoM5WRAl76h7uc73Gl5de35IZwdrsS5
elFuIJ6tcjnfF2jL/7y6q+6QSfd6ksmmZD3lp7lBpo7OxlrtfVjEvCTakMUI
vf2/sxe1zJ2tS5w/Tb10KPvX2xyNPYFnMYMvuNigOvs4kECciVP1ujWk8qmX
VfOOHkxDoHu9VDr7A6nF3II+Ht+alTyFjEZAwMrjwkpM7G+2hP8rF17/gZiZ
gHiOginHx+0lDkw7nUAw1s4+BCXWSUtxIZCAq+9O2Mfa85PG0q9lZTKN9fdS
ol1EldW8oAfhqVZS77lpvFc4gG46J9YS657xMoXgy61uXvAm5IK7V084739N
Ih1pYu2ZVe60juUUlLPhBMiYu3q7jqm9RMPdIiBn7hYCA1MhoLL5tpVzT9wU
BvoRfIzlfhMqgO7kAbYsFqb3RUelXaD8nDTKHZbazbR6hqnanbFAgCQJq3ff
vgvW/a1TpckDBc46aTHHHgyfMqYOQPkef856qbuNbXhkrpheesFttTLIgLig
7qmHmSjS8miFQumge9nqaS4JlyPLbI00a/rTASFXOWvJ3vzqxt8mw/2edToL
UMd4n1U66swo3kCHbu7/MmcdTByrl7H7VAk25RdFbS1mAxlMf2KpXpKDO7XE
W8VcbYNSGhiGA9MCHCDPc3LL+xZiaWQ2lqHNjYlLJ5XT+uHjZuqimYoXXuzY
reO7eMtfbmU9X+PnPtXf6YCwg0AsupEJcmGd2kgQ0JVneVcVvS24OUi0jWd6
3vbnXCiAJAfc49A2NzCARDBKanxckkh0nEK80pMHnls/cIqmeXp/EVXWt/4z
7L+IE8mjy7v7ahEAX4lTPuYaye6eeV5xGYYD6/KkaoYAeUnqwCh6frEF0/pi
jdYTbL5eeQKP0bz9L/bCbs2P7+4P82VDwPMs2Nuiujpro3NNOlbFRQf6b5pF
c5ykTNEbhYSVUGxNybZbOjG6d4L4xWa9QEY222qlrslQPGrIWNEIj0pUB7RQ
jMYEU7CM304J8j7bc3yPUG+vRtRhf/bfbMS424X7lGNrgKwD5+Nj8f3BJhuO
YJz+k31HFCMaQ6A3q+lhJzpzEgX/KcAOpjNImvkI7ik0KWcGVruNow8e3N5R
l9nv+9k7PujXCos418LOlIotBceKD/t2zwrZfbXaGPxAQtjdjwocqL5O/rHG
JfaPkEq7f+MMm9YlTN4oO7ET/Z/PcX2XxPtfmhFNFHM4cURKAk3qQDMaOfHM
f+vIC0mk5+DJEon0mNs8+chUO4SJlWHbwsoiXI6rXQ/oaEkKjiGEq57vG6Tk
i01VB7aY543O1Ie/OSN7k7YFCsx8odPP4R0rr4xzFCe0rR51D4lig44PhJRJ
Y2OPWoH1uqrA0nfR+MlCHxLxd7b2aFN39mKpGbbi4H24MI5ojBSmHkY8+ZCS
hYjnOaD4Dim+SQSBiYD7Z8lYw2qbjHHuSDz6KICVfz1HdEofObm7XVrDNxc/
/JLzor3ilCy4cKb1tvjoMdXEmbQUtCagVZQw9TGv37m/weUcwxg2+cUrc35w
94PnwZ/UoByHRwMt/5IhCdDNqH4eNCahIBf9OjxoLzsEhSPNHK1Q01/YVBgU
DyH8m4lQ0FvZMyRAog79XvGMsi/ROIrZwMaLJRVzdAO7RNbD1z6t3I4hpFgZ
9GLSvUhuO8tfKkEAfw90cRx+xuJvoumGAPSxArfN4vipDUT4UdT5US/Nb5If
InuweWuOUYuTQ8BjyU1nAIKHbg/FinQgd+QS6hXbbOUBdkRosuiTzFRTudmS
BsJ8ji/euPujHiuZ+oKmvuwqdQXvoCLWxVrxbSLbkR9PwFlS0DexqiqwaIpG
if7AnidFkEGmVOANm9z4HVlxK0UokAS+vkfwty/tVdtBmSbBQgJYo01+IoUD
R/Rz69ej9LVYN5i/pvIRDvvgZ2RHwW/YIZd9BlIUrJ/Lh4nzd/KqMwtCAozK
46DFDmsL7eHFUuZVT+pcMCQTvfNtyqw/hQ+e70QkK48vJz4sZF/9O1SdVB15
LWoE67V/Ufb9bLsIEv9rHz71EZ1CDqopGs23SzNmXJ5K7C9WehICZBaloKFy
zQAcuDQN1MWYjFzGTLzmwCuQbBJivqNKf7TubyCO8fZijfhl0/W9Zbw/t+Ne
EZddmThfDscYAQQ4PPh7aHvyVC7SUrMTxyTAkx7YsSmhsuV2iJFJPaYrzov5
gBmWUPuUEBf6eyUF1coPpQYJuvrQklu0KIVb7kuGH/QVHsworVZl+G8R5qk6
Katffdwn3anGhIMKsQ7sOHLlpgmQeg43Rhm93opN7kgZj0Bd+lEjccvl/77b
R0NY2UUmRVrkORx4HgTFiAxZeC+Nhv5VlZawhFMb9QbSc2ta9uswVB1xa+HU
RK2WiW23ducnYU1hWw9p7xejn+rVS8xHTovIvVPJxMHNXb8rSEfAAaYQDY/b
mUrZU3gZm0hMxvaH65il3RTmYsesGwUOF8n/D+K5WzQM+IQs49nk3RsnSxV1
wcUE7CwrZfV6LFWGQzYdk4oeE0+tc61CEMstSBJhIsGbjVefbzNozUOf9P+2
dr2rK5CUUQJ2Pi8uOTejejUL0INUf7JXWcPZhoSJWRByrRybhe4qyVVMgcaH
vzALTqrBP+o5AYk+Vl8xhcCW9fI6dHaGW8bh4JD+YR4hAPMmDMhfa0bLlc8o
S9WRfJ/e6WEX7AuGLLd8QgLvoji8uWvoGl5xX1zjO2MlS14G6cjC/PiUK/mb
+8s2/Pv/O4l/ZaaiBHv8eRQ30q2xunnznAng7pgeYiJ4tz82jnTW9DDRRWjn
BfMilbBsSg7/DsZSOR34A4Ts/JKdjoVUB5P0ncqA9fyy1abbRsDGwYni2duc
6yBxqgpF6bQAdDSeUO238JltunC4ne//caYaIwRr0RYxUp2hFplFXxKVVEYJ
6Jgg/o+mq7BJNPtw1Q/R5nKI97jK6CZnBMexJRJK55WfxnLtABlZLNvqww/B
IdwLjAy9hEz9cZ/92nwlQ7XOeFg8tdzriEBFa2s3Z9S8Cpsj9rfjYca11Cuy
mhiTl4p0XNrDB+bUTuDaaB6KRDbuwziH2kDSbl2rA4QsJ+QXnbR/WdCGfr/T
kp6YtG4Wpf93eESlfGyeRxiHDQZE9gVqlwUz2LqWs/w/FX/8G0JvS3i7BQu7
/NG0+Rfj3vCLrnHAuDXbY5skzQqmHobE3NUcaydoFNg0IdQka7WFXJUokSrg
f5z2yQUwR0dMM7Og/47FFTK2ALqlzCqLTsd+Vg7MzILHjgMp+0Xk67F3ZKJw
r/ezWfC1NI6vgwvjNzUL8cDS44hSZiqIquhnHW8taxoMNpICbiFsWwbSmw9v
4Wbz+bwpXOYLalOc3Zy15ZPn8fOCUpRclUpH8I7z/xAkwTPHbecEzCfuFXP1
QAu4RNRp3u3siC3GROki745xHZ6x/JG63dxoLoQiEWfeairN+WhpRFg0lNqP
QlPhViwzUUvTtCZeXLx7sLvu1RXKNg1xGSW2R1/AfGxj2Y0KORn1qWk+GM+m
oDCMOvgBal0CJHMUJYxW6DKoLseRxnql3vk7W5pMBx/lNAfpfHakGVVNk2JC
9hFN7wuONAkS4ZNMBuuX3rXhQs23qOaXu4GQOq7na065SpeanQDJ0eJoyZWW
d5850ACJlhbcF5u0GkPY++F83d6Na1mMb2XhpTuYXNROoJdBqdUWEgVb4cSY
ahXUsXVPY7z5vHCzL2nu2EgdLBnHiyqBh5L5gPOdjp7CZSYhVKJVDi3pvMv/
ErcCkldxG4OWn7QXmHzHZJD03AV9Og+rzLcReQ7P5C2x2nM+4JlLpZZWq6aH
aORV+jKXmxwsGh6y02/etjIZ7tEovhwtDE1cUQEQ5W18tc+P0N1XTtp1iX2G
/O/QFciWfo6iwRzoeU5EtayFiC8gd/KsSQTCH9mG2asee8WMMnjr6ylv5rDp
JrOnCXFNRAHJjRF5QwmtDhaeP54pbYS4JDkpPmQhFL3I5zLQ5SJKIgYwH6uY
51eTiuxrhv6Kc18WZdjSy6L/53b0I/VXuvgJk65MIrSt48xwi7bTAI7UlcYl
Vn6dgrn/JW1vsbxQA+h68HjipZhjm3p7Te5eMnbiODc6GYuMhzmz7uL5GpS5
doA7DnpyVnGuQc0FN8KdjpNkN/UCbXxj6J4/0f0D1MZSzkxx87KejU51Abw9
0PjTK7zsZKxzP2sYCzLkZBMi5/jeqmEWlJoYlBc17k7ApXpxO7NiHx+G17GI
ShtftBoTzzMfJX6vAyuR1rHA2m1aOx9i9mTry5QiW++owNT4lDkhYyU1aJdY
8+mUFIzTYQHq2CXucav2NvsB4ZqVxoss1oVL8jE/QDXG9Zr9wHrbKhlKx5rG
8vGna0rbcur8//lOjC762p+y3kcSU87GgIxfi7ndOMNxisrlfezHe/Z78JcH
gxSQJw1K4j61se2ofVwJOvXweZEsm8yb41J0Ek62JPYKdb37XWwomQ5jtY+5
NjF2QjuonmQ06xNbIsCkO6qf/6HBmm/rYc3W+1ijzKMCy2J8+t7ebFJOa3Af
LY0NdPSXkJOcP4d5PegIGEPhObXksHFVnf5WXrFuf/yZ/STp4qwEsIFMpw4B
iYOJuYT+RwCQq0GuphwKuncHQ+DUqgFtr2eezvS4pRqUQQtmUiU2KskWAGJ4
y9+ofUNuoKlAIX795wk7+9bdcPutQIyI765J//lg7tgE7Ef5/Qrf6zmidNLA
xjuxB4Y0JqEWL68HDevRIonG3ndvkeuV6larBRh4NolTTp8F2vTo+zGEmx/G
M2doa06+EEHqQguwHlRJEf0g0ANQ9gWRMUd6fTkluikRy5Ep5sSVd+2R//Dh
8ZCA47YlX47FGDOGKc13mqXxo8LYOvme67Ai9lzRHCDBFWtclXB2srDS5fZ1
kyFaQGL0hon8G106Nlnt9XsNvv9yHfs2YW+Tiudmy/rV1wTDyRnEJ+BSjpO+
P3LuspeC80b46xU8ufTDcWwfgmqwtxBEYXV65xb5NNZ9FDURt2IOoYrJRXYK
NxODFxgzfGhZCn4en9RyRYUo+riBamdruttS1SM/fPk0u4AFLkyEQJjqk5rD
l+Qo19q98zRrHn+GqtCnQinhpGKi1kz9kiU5X6pt49Dv98DxXJTEauobouJf
3RkkPY1eYGikGb9Jg1Bo36vsPE/+aYjWpUxuWq+WOAkdBZSIiXBUc2ybBs6o
NamYik4+OUrYM60QjJd01/9IhDLzlPthBXnfM/sytgY1t39cVrmdbQeDUcdG
vhnMxATbtq5EFG8I/9oD/Syw7zp2Tztmjz+FWhWoIDQOLWeKA+iPsuwqOssF
aCQEq3LcN0vEMCYObc3sMX0NweeHEEXvfIihDAWRCtRMIxifnsSU/yJRP+NW
bpwY7xrz7pkBloqoFH8iSoPwvjSwT5JQvGGn4d+norSUrhyOTL5z6Hfsa5IS
99Gs4AWrpkjkLG+Tl9R3Vdo5LmjFZP9AOlJMEhXyO92zS/b1IVduNojVfoTz
BUSisARoxlBAImYVq/CzrP6zfIDv3zHsZ8kg4bzvU+NOuu+ORwRBLOPGXnXm
IIvc69N8HyiH6hiCCraugRO6eo1vHeEsBlrErmyewglu4jS48UIqdYo9MKtG
hXvQl3SA8n9v35+j/tcXMpqNLi1Olm4leYACRgsAfw5PN9saWegO1/cL1jDh
teFtqxF0YW+QWXIP0nlisqOERLTYDrJBagYISiWfX8RSF8dtiKy0XCEOdklS
dadX4+9WQ7PWgvLquJH6k+Nx3g3vjhJW0vEQNkeSHSEErgL2zrxGB8pngFgQ
6IGTI6k/rJvPLytRfvw6VkdTmm6kvLtD+84zScHHzQhXl8KgFvbY4iSt+QHQ
Jk88eccJ1A+mW/74m10OrBqj0SQ7hWDZ3vCBFhLBvt6WRKCh6BvcIAQTB69n
ne4zkHW5n5lvCYzBoetxCmKP6u9Y/fWpvjrlrWnL5YhSxXysgRxDLjzUFAyj
z2R/tXslo7ES1aOe+7K6grTyfBYPMzlu/G7mnGZ3IjGm6WwpaFtzYE2K2g7m
YpkLqhk6DaMIVZwKf2nfwBTGxFp23IxRFpxGuBJKAMtz1fwOgOpY40Yq9Wz8
vzxEiR44sKIB4y5v1HjVOpmv9AsziMLthS4TyuO/54tOgskS+okbmbcjdyXT
rmniBNXZflH/HMaYhE88MX0EwQTiwdOJ4mQF5FmsSac6q07UKUqFi03NMhvU
JINSdKQz4Vh22/Xav35xTqIwzP4IEAKQl9UPzJtsumAx6SH29GC80D+GkHnq
RZWZ8eslzK4a9cfhHqkleWj6qZfomdLRPEoIXqMp8P7qAP2TSSzvzwPnrHWX
3SyMAfHH68K/R3wSkAMHvxCjBzzczDJNdCHxoeLPk284chHUlER1GNeUHLPs
7ac+vVc51heljDb5awzCVPtXNtwdYOQoRaXC4CbpJaR9cNOhovFr4GSdf6Ix
90IZAl1vzFmJyTLdGDu7/DdZ3P80tRfVH11h3VYDvajvUJFYdp3nXQ/ZowX7
JWvPblE+bPEC2hG6zdCZoR6VL67a/U5a5UE0m7+mEDZeoH4SNXX3irNr8sHs
Bokf+G2x8fJ0/AK7VAlJGga8oolWCZIqvENhNFKcteEV2fvHIFFAeRXB5ywt
m1ZvC11yu/gdwMdT5SultiKtR1blZYuu36GpKC3ggWSCUibgZWA4WDMoSG7W
ho86AgmgW0ZD02+2E0LV5Vv3sB6d4Jj3qBYU8oVUokQ0BzA1bZU1ofSEm+5Z
dcA2FRubAGs2haY6rtWrsLAkpluLUtu/p/RGUGnE63P76DIM3QGUf8TxiCqO
5DLXcV54AB8sWMpAqzW1fVaiQTfxn94rT7JkVW8gcoKWff0qllNOc1cAn6Ky
/Pn6aqbxV294ewdMFq41tb0lEbPRsh35ZNH2PJkNnfv/u7fbRow1jFPHfA/h
SY2NxFOgzd8jPU99vaF6TEuVN/a3hqnQPBvpPGg5D0V+bVmNgDNXzgRqFaJ8
yB1/xued6sOWhLBeihaaq0X6kCkluxO9BEFEb6aUTlIENUhky0STe6uAUEM8
lA2zLSXtOaFwe7rO4RMX2xJ/2nNeFyednyn6N5ZRrK4WNCUUECrmYbAdItbj
hVXUuTLwSNbh1j50onGhub1n7KuGHptb5pD/FVQhPfxgRUuXL91fMIUVrKOi
lK8CIMGqEu+eLm0zfROVh9Jrr4x620En5FXDjDvyElIzPYYOCijSYWuQ03GO
iPAdQ5eYzwSeWQmejJZ5nPYunYgt4+fM4SKqY67Qpdon7Iy3Xqb0KbaajGsO
XsB7+Ff6PsyyUXFC4Dn7ZEt7FJ1cNz6oJgcaC3gSMtq0a1u6JTqm8vogusYb
GhJT20wEmI7Eq3Rnocrj1yyPk2JYwPSWd9EmpEKUVYdOMRkWEMWTidN40wwO
g6vPoHhTuMUPwekuh9Yp9qEkjzMsV2TeXeTDptrTTOrfF7SWHb47KcU8ryQn
js0RN9Bf0R3pgIdiRZ2fUm4/RZFFUEO4MlICLbZU0/MiQMUL4By1mN70QScI
3Bjm4zIB5zzq3SCyK5TMHasNsiPPJicFBZdb3cdZXd8h433+95Ee6f1smPI7
dx1VW/oi5YAaWnt+KCcOA4M7pw9pPzrUoAQ/V1BAXLnfj0kIbcooD7WEeGNM
2RgP0APMwcKVxA2tTHCN4+L4blXpwKWt0hESB22uK8nk/G1DaQmG+phNBNnq
zHDBaiw/QRW0r/1qAhhzV8tR8adll0NDVeJbIh5hqJnE/LDmmIdxS9fEei8W
tSy2FAyL8y5kh3rkxmz5qn88UhvKo0cK2j9fijzamvUsvot1t71VeUu6qZfp
fczMTRKEbv/itpsJmZ8/EMjL/QqlwkmR3ERKf1F6zm1MFqsyTeVoEwc19NGM
5zuE4Y4Erca+rC3mRecCmEXUKizduPRrF/zGLsYAmcy65VlYXXQclWoS3vig
+NpksffwH/+xumjKjepUi21R4xvHfax1htpk7lEAbyzFq0zDGJZrFXusqHpx
cJ6tot32KWSYavfnKA1SPnrVG70PoreAC5cunEIWfPtC1LlxzcXyfM/fFTGd
K+fGnyCRvHBTvBidYqpOE2STYG6T5HaBokwkS49Xm3iIqKWUiuo7XYO0dIJc
lXdoFsJ0RFbmhF/48+7cgMMvNh0UkE1PmQ3mNQFaIYoeF4948ERJ27rkqS2w
zaZW55+fOsf7Vn9mlljiF8440ba7MKXWKjL5QiGfWax0b/p/s1M7uy43W96T
cYzJHK7zgmSO1SzOuELAGraR2Bx0TmcioYlE92WHYUMXVrTRoXx5/iXa5OqG
Lau5RLc3azJwxp3DTnRaziWwmH4mtKYcFnFCWWkjv+RUOWe1PFnLoDIAEl/J
GwoQVfWFgLVKFCHEs1HZlnJ/2E52mYP0zTO0FNgzVN10G8T5ILhMl+ebFL1q
OFdpnPKhoQuXlzCnLCZcUOLsh5AYXArTWamVHrtzs/Z8zGSNl5WjPY4TZVRC
Y85FYUwoBztoDXXRCEbLaMXoyTSjUggOI9m9KQUt+dbn9UoFmIwdK7AASHst
/fhmUfS0RM4nu00H1pP4skdCTaD//1Q+0+wg2Rb0LvmRJD8zgpiCZu/2J1ER
ZlRZTh6IRbdsULQjetPX+8x6CPiXdr/TL8NZl/IM1DR6tnqPAvPEfq9CXeoD
3xfzgUc0UWfYt4Nhx05bMKcCyeRbJSqnbrj2eDQJA5RFLR1vWvFMhPqMYzp7
d1mbfRy+XFYnolqNuO75GyHCR+4lJvAjEZZuadHhHdfkomI8/oqt+N8C+LF9
oh3CSYYjWzBUpL39yj40fpHmcWBO0egFA3dPwYPx0w9WFKZtn6HbgeOXjhRr
J8djvWVzVXb7qzOsy4k7nQo+mf/Aa5qsCnFL59UOquh9Z0SnpGFhiB11Gf6q
dfgMz99bQxx8hVX7FAVQxQIA6I/YRNPOJOWFh7Tu3KLQIc2Rzc9swD6u99gj
GjzuRGODA23zdyct2+shXnF5DeIpC7dk5MH3ZbL79Ecp0WbHcgmL1kOe5fyj
zFfZtnA+J4SEtsrqGxIRrVA5+KzjJJ6rSv22Bw0QMxSnvGuYALjE3g8WUsu9
WB2YmNeSE1XOsqJYPbKSr5KpOxV3DWKbCNK6V2RtUxU5VBk3Kc/QskyBbjD5
DaHTy9bgWFQi59xqMr9/F4AJ4baE6Xkq20WNrwC5uZ//0SeKgsSCdYaWvzFG
Peq61HIvZUNPQxJe7FP6y+Or3LKjOh7fwvln6hI21xmdOMxqbPY3285/Igw/
xRSWBzcbIV3Tygd6rz3Vh8RNj/yBuI0L+beDBg/XWJWCXs2TzXHQqMQeFPrZ
Yzt+ywXjMp1X5mCHxydDDeEDJO6S1OijZL2PVXMYJU8tVSi80dUo6KVkyhw/
On/+k0BiNqCtP2qlT4AdvdHDRxPu45X2U5cDhPAY1rMpwU1X9zYySBasXYIC
m3RrQBb8RgXtYtGKsuSfZPJGUmi9mS+9P96WQ6Lwgp41S2tKrEXpdT9uA4KB
cDIXLn9MFJqjFehN2yHXM3vgE9uSny3bShAlTBDpfk9poHcFG+WNZDPYCNFy
kehb4r7vn3IQwv8sjOdRjbvcSOyVnZHlyqQiWTmAKLa6qYPJ/gUugeDYJL5S
PcyOD6G/BL6gVFEbQr0mTL2vWY2HeGqcS+ZFfR9iUW/1f6qbOo1Ng+pRXt7j
rjnruWFVi6OZWLRCUI8b4Svr6+2YLuecgT439BlBETyZ5nby4vsHCvotHU4v
SJ/x9q1gPJru3ii+iRFpxl55PCcFsL6y6IF3Jywf7wN5CS3k+y+H+TKY4rdD
PYBqWRtnlecx17Ocy2qzo0QOVYvJXH15Mi6aIZjbgDLfTQ1xUL1LU8D4iCSU
9EAtJqj4fszhUf74qQOTDwuWF5GQETXwaTyAgkN7Gy+XcQw50jRGyubnSZB/
93UZP5LXocz9qCWb81+ezQoKV4/IBOE/e700Rpy6L2cNIXIdeMD/EaB0I6ga
sFnm9RhMvM4YBV/eGDdEKOqaMqxzGq2bwHVXH5uu8kgMfqLJ7fYimVP4Rdhd
ZcnzgmBfGAkndMdDZEMMCw0wbmCUMPbUhVe+cxDqxBEcXV/bhePzfJQuDY5u
ICIGGbSHT1wMR8ZshcYkT2LKV6EYbNJnimket+/6DcVC/msgmxoCKtjCw29c
v6h/36CPLDqy+sxYViZLH96l+sT8sHShIIqJ2zRQN36pdtNvu5mIohlvavfu
Z61rOVfljhPYa+MU+5CO542E37rSzeoyHssiF2owMQQ63G6u2Ws6uTVWGGaf
yNHN5gpFH5+SWUl9ycW06rmll6IZmzbke2yyuqFEdiEWu6t3jFO5JPBRf35M
X4phGzrH6DC/HbgBeHXmdCKjf8OmT3SnMcoOen133HpXUVVIbF8uet21XqvH
DwwBHlOLz7ivymZlPsRn1zD7smssWUoI7PUQetdGHOU+3ndqRTSo1rKGsk41
IKVJrv8vDGic12/kgcBgvFmZcnIOEfsM2AUNuicQrERx+OxYPNp5K/etbAwH
QCvW5H+oL3VgFBc8ReCd1M2Ng3ifan43Pk0OmhU8Qa7FVcgPJbgbMAKHakie
tDhZYhAdjl5mNMBix8iXXSnnayJ7E4+jImGk8dgq2pixTL3adUhtm6zgLgjW
2Vu1LGgS4ed/gFLHxZYlsUCHFJb5z+iCJCcxkjEqcSiL2j3PYJXNAWeu7hWp
kiH5z9gTG0fNOTI15wwlAEujrNoIm6eqUg/g39UbXV9CWx5LftnwtNbgua0H
QnN091wQlNt33kDS+XJPm3xJJl8euigzv4bI2xrveFHfFFk4kbAhWfYaC18i
iXTJoUTIBkQJ2h3fDzyyaq6LxOez+fLfvcLJS3/M0uuWh6dCn9YS5Ey16ds3
YH7LCEjZGZhNq0AOoiWN5VrGkPYM2R1XTORyoh/odvc/Il+5wqH72geo0/l8
AU7NIIcvGBm9BMXQMzTN14hVzqOGY366mRSwF7DYs3b7LhUKVny+BQxyhrm7
zJkQrrWv+86b1uSROiVDaZbDQf7uYwI/5KN8alqaUOSdyWoAiXTy0NBom4rh
jivamW8xyvi2cnZeJDP0t3RVs5vlem4RrFJv7CkUlCO/klBMjHe3k9l05/bJ
oE6fqXMkdFQg/i+fc3fn4JwMDGgMEGhJcOmkdv8XgIfQx8lPTH9LTQzrWWZv
9k/i1s9M8fM7bGIxGQGQJbISQYNlfAmI5kDl1YObUM+MR18DoTu0Qnibf6Dp
ODyGdA1YZm1wPQtw2UD/aWRQBWK7ffpY7NvywR4Zp5kXz/iTHknmSCvCfVCi
1IjE+K0G8D2LmhyxL3kuDeCKlUOVWSOygYoeRY/3QVl4qI3NB5DiWTx5y9xA
iPiYX9mol/VmHHslJG6kBrQZATlClcw8t6XcUMlihEexqGN5C+awUW4OKyMp
YP0Hp8pNRixlMPnuwjgCkTLeKHZofocnZCadK+qivarm9183hLT0ubSKVkhr
fe8wgV/Vn24TQfHoJqMjav5igblEgoYh7igHK18cQvl+JH5kqhv99AhOIQNT
Jp8F4J8aAo4d3YWXsJg42mXp2mQMODQjDF7htsMFLyvxoPCyA1XkD7ppDn10
LTzcrZxuROoKSFIT4yymAywcb7gTPNsQ8ESemqGwEzakWF4vrYRjiRXc19tp
JTToMqIYKyNiz+qNNaOHdtyCcPkFmG93k/jnUCl5OsuZwrL21I6vjwc9xYKT
0cv+VCEUCs3mUxH65thM2MvUqRxPI0n70QEfzkUI6SSzeClaDjrXZSVUgACv
QR6XzzADwm7nqOcoAC0F/WmYTpnpID7tYRnvC0IkNylaudv1PkuZo1GkmFdW
BbAlgvemEuFBt0Ul9jt/foa97Ojeg4P9onZWXjYT8ZzGd4/UbJ7H/JEd6VHy
RzF3RB5qcNpPR+cWSXFahGSAGkzv9vRUyIhnQ508xy15Q6m6sOsh90rjLqqk
7Aw9az/L3XmDYZMC/wFR8osiNhvTGB6yXbYzH2iFiB9uuznZq8qXshjAZTDi
s6j5FFVl1+D3mJU2e9T3Bc7lDsHgK8VReQ0URy1izxxR81/CXoOGq0aBCSYz
+SOa0i3w83upp3YfISF3pdg2dwuNp7ZAZiMLaSrKDDfl1gpVZGr0boc62IXC
zS9g2/GVmlDuOJa9PUg5fjEDMUee4yIkn4ISx15HLqBxPW/r7mp7roerEaaG
dc1GWmoFChL82VRp7Dnnu8gP6trNV7r57Iw5iWpsxej//9bCPNj5IUm8ibdF
eiA94BWuBDkgyGo0wF7EVWIFRElJM235RqAomLlbyLk2Z4lEw7UfszqAQkQq
wLwr3W58+ERApVDXCg1uSsl9xaR60RU43EHEJ9xaWbNOOqK6/rQ9TN7DvrYI
ogCrBhtuEop17R25JCgZZtHSXR57S+8yOASvYWI8+RQHn6R8rfxb+y4pO3vY
0IfMawq7qbiz5HVWZnFMHA+FVcmPt0Pm4PB8FVsNUI9FBuPJL9sf6UAsRZbu
qYubb6QxxNaUpMAly31cchp+0cziAyA7qIWGTdrL+v+XVAUn/0syAqKbSJva
E6UMB6GBN52R5upTpjnIKPP6fZzRW5LTFZkN/BYnRAjZ35okmNJ080m2zYYO
ZQ2fUsRtRWPHtABZaVaPOqMud1O8pAD92wYBmFCbm30DnLryKfockQTOuqeL
0yj4O0OYI0MAYflO9pJWbZCPPqV5xk3p+wHi3biDF75HtKZULK96PPIdPuSl
6/YJlDT6cJt24r472gUWMLAaKc7pRPKY461P6SM8onP/dsnqXMt7XZea5sTQ
RqELQfONmZNsrLp2C1BZKHPP3xdvnDl86xTbXKZLsHrnq0Yo2pegMYg6+t0t
G68boyTaUt6vcJ0DYFjxd1cfVepQALZKw+I1ZrDXwux8+P+t5I61GQTZ3hLC
Fc2l1zZLrrNEeelD8CEBjnRRBpWzZidcWbSU8LUqA7tZftVG3Zx7cEW3QN7L
80+IUfIIFcQUdYsfHfZ6x3OK0hPjw+CaAIdqupktDZDdIvn9qxL4NVG8D5ZV
OiYwYfCAkmJe2MHM97zAeOhidRSJmwWwvJmG1n8IWUwlBC9RTNxonX8Wv0cY
e+pvu9TWCF/dn52BS5clmpdzSycID05qq8fwY0QRQmzb35V+L8ZNHBIS7O/8
KMb+1rr0LFyvc60qnuzeR2Tu1amlBc9UGo8OuyjEv1f/hgEHfKAlWp/9VgO1
1QeWdSo6UFwPxqA1G94Pv+v4u1DJn5wz6WICX4YIHvNv31XD4v6SxgLN/oex
BcPpKlK7+Uj30dEFyQT1pGB+N5C0ueD9ZCKmK7J/fTTFPI+lpCdtwQ96avBC
jnUacPJcoULFEZ70F6d4xdnOWudMKOiXwiuo81O2QgqnWuOVvt/WXjU8bPD8
ty954U+FYgoboqMnLUNCRQ5Fc5rl7lFRfUsXsKb9RJPFj2G2iRXNr0lWCm+c
eB1LE8OlcD0E/kYiCXhS4oY3WUFnlCGT9ravy90PAfQ4vKv9JnYg/Gx2ZD2g
nJwglkFjbTBhOqM7rHfdhSf74LG4kBsEjSpWuPpoC+syN2QQek3XMLHHmiM4
6r3PQFy5ggq2O/xFWxeh23MddNEHn6Z1UmG2kkJKPpF71ZpFVdKjYd2qHZqk
D01ijJ0kq3s40C6PoTIZ1nTqEpdQThIWoqqNeGMinHoQsTydxZR2XQQks7lW
FMB5psCAG8I8cs+2MVECaDQ6AJN0GIePvgSQ/+HaZXGjePLEzNGqHshbYnd4
8Rm20YjNJ9s1MZ0voNUh40BoGUNcvDj0HozNq3zdT3ub1eIh7gmrLZ0IOciA
7PrHJJ4BRkIN6KBr6mR+QlocDhJlH37adJh8szA65ZcoFUBAwcHszLqtGvBi
8Vl3yj1I2KYTHfPN4KgzWBEUVy4nE8+/NcZjAN7lWlvCf/j3cw7Q7G90BOAS
IG/h8hAmm8wUG+3Kj/Nqde59MUPRNvcXMzSdo9/C36u7Li6WLT4OsliCjokW
JySTdjpVK0F1Du/eupKn89KRWM8SNhRbtAg3bv38C087fPNG1vHXQ7CTRH5S
TkJK7jn4u4BetQ3heYIwBlPXgshgXzxRq7CRmyr60RgnPZFIRDb5friPS7j9
M+1qPg3K6cRRNQ39pmjbbiN555be/NqiYPWevOUlZ2zljQrmy74NPDnl/Zn/
tDD/6Op+OL9eO1vC3acbY+NR6GY1XHs/Q/A1yUSGPX9GWrg4wt52vxUHK61e
hhE+Cy6r0+xI90czaRlvZAGeaELmRz5i9RS7vkYsNonQhGQFKoam8DQPDqeL
FvJ/N3RIn1CPuWdfnmhnd6P/7WKBeugpWbMGco9F4gXd7OuX+ZCRITeKqUBb
MjRA/3xNn2Ry8tqK+UojtSRo3/E+XUu1NpK+dmjgCTF7SI297rpD19Ggc5dS
PqKkLUNNkg53bA3lJWawWmIvQfFRIjWkqFEf78BnJJKkQ58/kIUMwJqszXoR
gNBM2hduofk9G/2+Gkl6solBt3InkxGRhgPDw80L/h8Cw83AHaPBzHM++d/r
cgTNSd+q56TY2znJOSPXgEEXYM1cwhXRv8bA2PxhG34eX2j78FjgGGP9SDHU
l6p5i0uYnXcOXJqoSvyvLM4lpAFI+eRMi3WdYfkLuxmhI6RvgH4DWnfpAC/n
PAnYiONSm/YCxj9d5VKfTajv0qPRI35AZZz14M0f7ZkFBtKXu9+GI1uqQdxM
xgNqPOIMZdv/rFcIqIo5aeXflgDE8pE7MQVQqx6jIC5oc0QLx+vjZ0yqXwly
EJhgKCB/vDseVsF7IZ5YEJupakgwHcBiSlJ5vl5z3dKbgMlq3GouDid2WcNl
k+MKLAxzFttYKdnWcNiTY8+DWGd7Kz7oM4POzyleAwKYBXRvS4aGp8/DHwhR
viRnW33m3VY7PYbbIecTV7PtVDRo680XQw6MBgx0b4k9Ozq9612bw1DasDLT
VLJnhdVwgUUMiQqR2JF3/r/aGFHrj7qwn18egeoFat7yITxJqAXI3tg+TEeP
qm5D5yi2mfJo1W/38zvKNylT9vR9qWNdO3BRHr3dlwqgWuamSJuKdDR0OtKa
h2hcxpl0j3WJcK/Y9jYWHxKbyfAzTfMqUTCmTXc5i2Bzfp2XJVctQAW+FMMW
LbB8/X2G83x0dTjts6BWjDdKLcuwFL4ABDppw+0JoklgJ8c8w1kdxRhD7F9a
QsljT9g718viNe/0eWhFlNSVR468WL9ps6Kjj5IJDDDtfINveLRAysdzb3TQ
6zG2rmeNsp2F0JdiWqvRMU5bzEN4t+NNkIcWxHocWOyEU3hdDfWjq9ofE98Q
0oI4T6JQx/gosifMtdjs6pfVIYbWDAUDoeAYINuAMCnYd3bKdKSFS/pOZaOZ
81rNrbCVLmrcHcqwNilRbIG9iFioVp6s/4mzZ8OH9pcTfr8BhlpXHXYdwuCi
XlaUosVXq9hAyIA4UxVhuJBNGtiusPykqFyIj36qLP1iM5+RqXAMSI/PKECf
lPzKzdcy58G4OY/FlVo6MlfPqJPCYzR8HjaEvtGzCMgSNvc82Yw5Z7Fo8Bpp
riDk9Kw4ry67Xe0Q9E3EPMfTygklqUIDUZU7fjHyriGghKVGPdcVt61orncO
GVUUJsFMhTrwoY/o/wcrhsUdNZvz4vWrZl2ReZ0iaCWFQCTE/Df3YPsQ+Lgs
jFdKnUFD9iavXPvZVLKLkmd6lCb6DUAoT8uq7PUCQCADzsp6435j2hGURkgY
yBoaiev9I3Mw/0PieqowI5OCLH2rgDU25/Wg8nJ9AU4gpbG2XJsLV6WEju5U
xv+T8jrGgukZoF9U9puOwxLsWFJE9jVq6Jfn7+O4tlc3umIpcOYVhmFZ2X13
Ot2rQxM0itaK8fGaEyaavyOg/WhYgzIXrIDNw54F+Zu2IDYJ6d+w9g+iAolf
HJFK/Hdl7MEhae16ImY5NqzaQqSfNthb3I0zPFBV2MLKXD410jNTMHkKL5Uq
rLiwC/NYsdZl7afWs7/7xaRh/4jw04J+ZTai/s9pc5L1zx2laVWnf0MnSBLX
3zRrjE4f8j4yGLJ2Bvn3KcIAlpAf4kkcR+UjpVAZVmKy8UdFJ7gnLZGK4OYl
FMbsh3YabIR3cW3TEbLl5kZTFBvy/Md6eba7LcmQ80wm9RpCW8r4dGfpWFfB
pfwTM5poNGk//xUztEXQs20RCB9cit1lCdVOTlLXw/UguA6VwX2myB3vZQFZ
B01JLYmqUAdtxhX0tGdK/L8eaEwVdfP9QWHMiQ52ht6K4MSARnz4mX4j53HG
GQlECCMdF9T/brEe25s+Nok7PA1OcbthoBVKLIAENYpKBFcF8h3gD0hXrdoX
ajlk9rbRkCOFsJ/BPzAFaIGPpBwgrnYOX4Sq0RBGVRX+d7p4CObUtF38Page
N9RlFx++xGrudfcaVRXLmiUqG2rnN1cOmoCgq/fd6FM0Qt3JMjcV0d33LtJo
DBtkIJJkevVOwTlxJPKPZ/Ta5zb2m97ZBJXCjCdTbCxk/jdCzdqcvOHfMTrd
v5nBkbLA1vO8ob+Lz5XfsaMYt1uzt0yMJJJbmBSv1MgtXgBN8emFkarO8xxm
mNWpchAiwf2Bf+yEV98oVkxOjhAc4iUhLt3QTMkb45wCyMSfV7znzNnPimCh
ZSHQ+nsdTOOID9Adm0Xq15N7ge4wYZov9mpQZQDGGbjd2+hUf3uhDEi+j25K
GDGisff4aF4L95CKoI7g2cf2cUfcQuKpEJUTc9daUNnDYKCTlq03rgmHQj9q
R3xV0Ib5EzuLiR6lS7lriCm1ftCfWRUeW6OxHBslmdFKPYCV7o9z1Wq+sUdj
H/8GL3pRDxNpZpCvuu8XDbpO5MzpLWHJw4Q3pj1I6+pVwQk8i4Hvpipk+MO/
LDbe1a9CcNBLxOJprrTfznRd3OPUPyX7KLcukx8w3eBIIUBSroJvdhpUV+tk
iGeKX/b8eRW2sh/gjXpfElH8GqZjjgt2ZJMF6XA+WzmQJjuu+O5F2oAxdGi6
AqunI2ENGVV/T+9uMmGsWdUCbDFDAo6nmGESaFVQuuqU2Zjoy+Slcz5rpn7Z
DGAptlM24EKA96/A7T0wKtNG2SzSY2LafV5o33Py2aYq9YQjgx86CGT1sa+2
Ii0lIJBhE+7L13HUkqw7DBHVLS6pnvahWqppWR1ws8w8SNIXOeN6wiWVF7uy
7FRBfLH80wKuIaz1tswehQl8cOV6mihhrB6Bw0Gt0SeLcoPwKWrJqDPBid7W
RRiPPdj3jv35NOKGUECNp0BLhNDHOsTpZ7IQcj6p1ZUL77rtddBz8J2euHrw
saOBROB+6+3aPWmpdpgCPsEY//wqPi2Whu0kfTR4pGd4PBfcvL9PdcKTnJoC
cZQNlpEWJlPJ1tpFKnxZm1hJ8CfZZ9lMjuhKEgYcFxFrHwnt2uVzVWfRtH53
yinAnqSTOg84aXzlwxY2goC9HULRB6tESE60rrRUL/s5qRPYMg/fBTOwbBPr
vRrizasxIWy13EI40pA0nhRAcWn2EA67czVhpBcsXd0gXNFR8Jebxf2gfS53
wIhVRFy0IHZSTZQhqKEFUDMRIOs6AHUZrgC0INGXaeX9xf5n7T4BJurOwfdH
W7+cUAS2MOHy7Y9hsoxs1CQfxtxYp9MhW0N2hXjavOqWZgDDrDVul2Qx8TWF
DKukRWaCa/8RPVr6l6VNVTHPMhItOqyeK26DSQxBtgUqWtrTfuGvQzUHj1/C
g3tZ8FSGHW3010dX1+fvGS4W3GHNll+g85q4IZLYi+RRQ1U43OHOlTYd+UTg
mZSax3orAPo2BjxuU7hjPPXvXZ1A2bpVIrzZF3pOHroXhWVsTPyzgH7ERbJM
FTSAuxJ9O668TmOwddGaqxlopNcdAmVn8W2NeEIMGd2a//2Hi/M67cr0TV5G
fVzyadNGJr23QIaGxRXiQnTAy2k9i1RAA4I9p0rW/MeqR4RTUnLbjCsP4B94
mjRiWXACXYAAtA0OHRRvkPjjENBc1MeCfXOCkRpXedzpjRbDmG4Z4KPKsVic
4FEtTtTzZKccI30bFMAoenPRKbIek9Ol5RErOfeR8LgH6GZV4Bjzqj7F0Wls
s+3+ypeKA+IOvqUjyQVUp7ki/9LSxl90Dm8rzQq8FkR+1KqsT9tWMURp/RUy
TA0IpBEOGtc/0XYUmKaosk81Otwv5Xj+meik9AexGKF3N5hRdKuWBHwDnH1/
aIsNdrZCGHZp/zrS1lJAsnKOnkvjAN7YPJ8hP2K0JBYECWs8ahy2Ib0Bx7Rg
ohZu0wDe1NSKQ0ZFUO/ZjiSsqoTDmfwU6DuDm/9omUZNCdb62yhq/cZ37bIE
11ZhvuqVmskpxP/M/E2ggar7KFDX7Itk6umZXPL0qFbFeMpMvT0V+lgESXm/
o7fvFiWX4XMVgiz6JKmCackrClw1R+5nYlK/dsCRa9cEYm30aR7EO+6Yilom
Ao7zjiCb+86DClLGlJ5NY6F+rwDBeJvTJ65LocXuKCvP97WVjONFdFsLpeWF
TK64Xnq6d/Hcmt9bKg/ajfti4NyJXw3/qClx4qdVFfaQmJowA+dlrsUL6OvS
iHCQX4EAdhS8tnoNd1e8fVE1XA6lpfRIdYl3tjOifHADUS1eea4BQMvwNrBh
zVmXc4YY8rDJ72kTdWNk5xQ3y9c6bKpa9cuod55h5L76oB0bNMwsTWsoEuRv
EUKjW3/Y81tqjyX41w704lqze8hKQ15fr/qVWsd7VE5JzPUlPjUI1tK2xR2v
eXtTlh4hxxmMXxFxb5OJMmI5FY79dD+YWDKBn0Q8E9iej8z/rsUHm+oKnLev
zAn+YUBzYlZTIsE+ie6ALQWvvqIQEOdG3yUpx/Ad6V9exE2akI2DY4+FKPNP
9CSx+2AAhIxKQjD9+fXHctDX+v+LSMrgwkmUh3kZfMgSqcOpG+puOGSNfv35
dmLwjL1eyERFZFyiZO2SkxgcIlebmD79kU1SfxyMaZ9RXVkLwBezpXhZcesh
cKPwZlupzm1i6eLtiblaAmCTOi+5IV83L2giQ7k/tWWxJwgmNmbnM2dba/9f
P3bxMcHACcUOLqqogZlOWdeM91ire7aczCFCoQgj9GPpXiYGSJb5B+ux7Kud
LsPyEaZBpX/KRsfqAT1Bnq16BpkBg7ziTYzNx/K3SLOk5ENjclYVAnP1COq5
SPQUQJ+EaI45pyo9VJoUUYguo5FhMHaP7oammqlt6CRlhBaSOP1zUtBYR5kC
+OBVzsuLJAoQGWK5lPMQurY2qvFouGOK/wl6sFajt2jqVfdokLus8HTX2U51
1qvPs2+99b1Z+TLpLvyC/LyTd19cGu3ImW5hZaKWqvkBYe1rU9rMduEQjrwE
viEl0HvEv23hRy0Sn7bAtXcBcUkksILn5AjszJhQB+Oq1LumJMTC+4AYUBw5
oYzPa71SsGXhW+UljjHWxUMZRlktE0CiaP8XI0ItTf1QfFa6lWNCucHfJPUM
TyQp/OZlXwx7TAW8ojasgBE6RnTk2ppoC+WkW3nJOKT3u1hSDgfvpzlNdurB
EP+p1fo9yyre8V8Qq+K3TvMI4k7HKXwaLks+P5GBRmRMZEmA5JlSOvG8tggr
tvA+yU6FMUPczSdjenPdnnJgM4uZBe7uEcgBqZcDt7UbqkY7t0snZVRcIDdo
huUS3dUwBYiRZKYTIeLs4CHG36J6OgHcF8gKjsNfblbMZAru8S9d7rv233yI
0WG+6YWtrpSWnGE2agvFmorxkYQYMprPIbTMjm/cIaBYwiObCM4xnoplXlur
PIfuWtyWsOY6HbjIJWkERJmsqQZWTCxvG9GcJPuJLpysz7f80yFjivXBzCPq
obIZtufWZWsV1KsELdMLygIIzT2bR+IQuG0uD0vPahyRedA8F8J9jiYI/XLf
Xk2ED8R0rrN7dQ3JMAB3rRnoM4M7M8St3c3u3++DZhc9G4XkNEgQTmLj2acn
XYA7d+PcFHYrcnqvjFMNfIok+u5b+X0F+Elyv0zHFAUJD9rVBYeNIxNYYbxa
KHRFel5wTbQNHJF3PJDF/2E/rNGfc2I5dWmm2xWHYmX22fGo4t+jUPO35bpO
T5ZWc10bH0/OjkoPvhX5ouX2Gy/opiAhFEUe5PjpDWn2bcfZYLWokwrKIh6L
1PtPi5lmGuES4HhX3epT2rwyUj/MC+SUZEr/NKcPxs1Wp/kG+UUyVVtAlta0
nCPfMrYNMU2R3h7dEHEKl6ebfjgKhm6/vrpN8DBr40G8+mxevCUQYLENb9M1
gdPd+5zCsD/N01GtjCfadgCDiMrJVs7JXQOL747noPYqi4MVPGJNVbq8xtqf
2OxSlIlFTtQGxvQpMvleurHlkZdDBkydtRfH0ylyfrBfrPsMv1AJZ98cg3KC
lLVDvaHK8Y6ju/jb7d1SvZVfuRIqYEHJPtYdEHEhQe7BGRYqet9gPfF3N9LO
LxriJT/eQmBm9A445XY5NfXzufvMKJTBpkm+DJ39lF08FXxhKKWP9jwM1zjm
rL5E7anUPYJnrpqdWpwgqk/+gNHt6DKZ32s5ZQabxq9S4st8wDpHAaosXZdp
Kkm5ltVyxmFTkoDtmYkwCC59gpwlRn0eDr2lO+FSrpfNGpMqPnlwJPP3pm5b
iTvWMdYifP/8iDRXvZWlhBodrGb6AlekVjqNSfVhwwNXHaboa8Y4TAy01pVQ
nVpV2XkPK5qYzEaqdLjv/Z124sZ+jpnNzIYekjkM7Rr1r/RFzccXKmvX073Y
TUZEKUPiFdhzr6KDMVNlK/INlaFPfDPvlnQnhm0VrAHIIIlQSg1JKKytHbHD
U+7sKUixagRba1pHAUBtJAaoGy285ehBF93fazu6chlyvMlGFM8Mrx1RWPY+
idTlL88nFJ/0b7ptV28K2+a5kqD0Bfp76HLiLoyLrX294IlUBgxhPVe5qSyp
ObJ5hpNHBDq16H2szRQtpZFnVC/YXqAbXWVH1RVFJvfL+vmbnpzlLxybGddm
RK4+xL5c8fFiN65IiHtIwULxwh3Xjr8mNROILJhUTA0PQgSmpAgvYN9C6UmU
8cdoJ5ium+F1aFAKh0YukGqYmFxgassUgOjD8k4pB74S3N5N6XOknpPZ6d5+
xs6TDXlzamZo/zyH7INjVomlwxlbwaiLEWe/ZoAvvq1ehRG12lZuQXe8DiKQ
beTrID8gaW0e8zI20mVxg2R8qAEcvWS8TC1+7MXd5hbHATNUM2hCJRGTV2yE
wFAVvtVDqx2pkG9AcrjL2OpL0tItbX2m87kkDc6LUwOKlAcL0lVxKp3ORlvS
ITzz9rV+iqtWlaetlL2+uXXhfHrJqHqURJL4kwFS0AQmvKRI/TABVwxBCxjT
sSqpymUu95WYbdcDnbs/7U+oIOkErzbXAtlfDKSB2poNUofVfAtvGrzBvhUE
fR9HgnTDpfFJ4Ci6muhxDB0WnXQB6vB+DDqfzmWcuo0UAR1hfYVBnRuPMLez
Qje3QTlLpvYRKFJQB8zAGfbfkSATY5uYNgllc6UX5ZwGIZ2DQ2pQDnWlZcvi
CZYYX0Nx5hW1mKtmP3Ii5YKIfWUrcMznVW7/msb6UE5lGl/d7VP7KpApyV2P
/uoTtbiThUC9fk9AVuFO8/Mb4mpmlSQk0L+jjyXUdrEztfCkbbqrw9HB3VTQ
th4XA8Fmogrhm+dpmV5m6BfjV4btFWIwJvtFglUEqLxdxAoWwrewAJbqaGK8
Br++ZJ++DvXfEuvIUdL2BriiTN44hMFQ/tgTMFPCXgzR+N9anAFDNDU8sLie
2UQIia9jMz4H5Z09aPs7RRldqW3CSkxnScucrP2veF87LRvxqzQ8lG8dB6XO
7XQRffetlueq1k7+x18hb8pB9sjSVQLL9rSsbRMjI6b6yifuZCF4+j6MhW2/
dJ57ErRSlG2D4nFVkpTLjg5PKQY15ydIymbmcmYFD+tHvzhz3R9salvj52NO
rpmf0xZbwUL6Any45EuMLti9mploQQSCholbjkaVdSPnQczVr6mPNTBd7LGE
MsrTozKk3kjRTy6+sqgMPSZS5S7WPmh8iyc85GA5sJM7of5dlLlLP5m2lXNO
xqAxr/MCrRWcOtlztAXaWtz2qP78GQ7+UjeQgQUZ/ZQKHW3e1b0HG9qnoRCu
8nB692CMmAp6CvxG/o2W9p6nm/vQxczFgprrJaxrrcW/5Aj7AWii+eSkK9uU
/Rj8rLAdiYs39ROcSoHhy2o/hLDS87Isl3T56MaxpQB1BnIeAeWWgkLK5CtX
chGBL+0fqscGiypULDGNgQFA4pJshRGucvR1yklOdPl+ZYyRG01nRUR8oQif
I44GX2eFAYph9KH5rajt9z9MzGla9vXNyL0t2qJrEvbJZFiijcI4SU4Zcvl5
+im5YxZfKX8ASP+Vjw0JSJdtriakhYWQMX+sSMumJ4ItRcjP44EZnpwiQfO1
Jx4wLG2mNS3g1JJFoMAls7rfeSMYxdJ6osdXPtFd5OyGtYKcv23VTgzA2vLk
/zHncgg3dMzixwss/fRGRnDNf02SbPnkeEG/bFo+YSt2D/239hBB4We8ARDd
XCewfqd/t7Rvn+hEq8B4yr6UckLFg8qwiGPlYASMT/bCxEyXVidbloCpcUVJ
DisB623kN4fcJZUzB4+ChtGbtizNWGHpk9Wb9RQUcl6dVZ2Kf0KiQdcAuKCs
taPDTvRVlxqCdZ0DEHDd6uCbmouLnpG623Ao5glA/O1LlyfU9PFzPEdRWgru
HWWPLGlaoOkG3OIJo9jm7quUhqGP29Hp7UALwyQexT0jrR/DRPt0KzIVEF/L
0nZ6GoqDfRUZUueaVaQx2iCcbfxcd6usuGrWTah9XpwTCBKL8ygbxhD5QFrK
/L6JEWdss3GkhIS/iAiCOCS8BfRrywwNT1xT9jMnEF7VmiNgbAu7KppRVE6l
97bpmcKbN3dhBYQv1GAItTWgM7tDGE3gUyKT5oHKJTnA4fv4J06TpewyCoSd
fkRzvVniWD857csHpUReOB7ZYvbXGLVDRzMHOrMl4l4DnXtfea+b2ACYCrKj
H4r69e6eNZMNl88ZuDa6zQVTaTvkQ7+3G7UYivBeNvQk6s6pqcUfqwX8dwaU
dKBugDBH+MIL2d5VgJyJk3AbWoeytox7EIaAQZyWwrbmvwoFkK1NcLPSOZNu
0t6iB9P+hHq5d5ruXlIkEZ0Sc4PdMJrGb7mqqRYw1tF6tFGlXNmKabWFtZ0i
yniVqSWytIGLdCFjb5E1qdwqxWlP7Hm48ZGJ6lKAtO/xuVQFq0WcNYAe57yy
/3saKfmQa3uXQswu46CX4ZLGPS1NeAlrLcxFGUiUn1TMLu6HWlsmI1FhJawi
KpAyIM5f/5bd10CHEMb73lWbwD+Aqnm0+ah+QNvoDrdbRwlmO7/OOUjbCLTk
m/uDUtG5onbYbVb71U+kuL58Xdrb/baIDZY95dP9WcbozATCOz4IhrphRWAG
C6LjUVzdtEACNxM7IyWKi3mngrYsJLh/dEo+a92+XifVVJvlV+5XClPo3CMx
k04vhs6COgAgIi52gmfaqW/WDZ3VXda+W51h3KAwcyASfsCgHbuKquh6Sk7w
s0Pd/xSFP8ieFfM1hHVDHvmxfOhxBn531+RaWsV9e1FsHoxAOQGE34s5z0FD
4cTQ/g+nD5o9Iq5Pbkaxn/HEuPiAF1XuMiNtor3rGCGmf/Wn1YXAmNUeg+QU
kk09Kc5mIBCaLN33kkpfxykPhkoQL4VodeUr7erjGeGy/Sb++pz2PjkaIhv6
k26S+u8se8gHAnFP1rkSjEOdxjakSM712lDvFuxAq7OUtAWZwXpXxrqJMuG3
elsOfNWrOsdKJgG8sKdB8WXOgoOLBnmZhaS7xNaDZyVGQZtZxMOH78NXGEkA
letx+R8zj4co6gPFw3fuq/o/P/bLM0J3uZSKabTx3A2xFPtCSbAbn3afOcbL
oawf/HBTP9NFdjmSi8s3cEOtmB4zQPKjp1KfpzVZhwHj/++amRRMcaPOEmS9
SRbMrrPAT+gfeenmw7iyxBbk+jufIt+apo/lTvQMakRh+nxQoKyfTAXlM6U4
NeQL7WlFIRbmAAzGGHkPuaAXjxo8UYRby6lYRhP9o+5uu9oREzmjyf8dmIBq
0t7/r/OmAu9ztmA65fEmRw37j8rNlRtEHvDNYdyrp4diSxCvF5qtlDlIsAfr
3lpghC2NODWfraqBwtoyZW+TCFe6nDSBHPV87Y7xD+QMv6t6zCn4cIL8gpp4
sNb3zqnosjFlcJWnPwdxA7DlQ6WR0WnsfO7Sm/FO1f7+QW3B8PtSB5Hb9vo0
DhGXXVbKByi0vYLLfKzMmKgggMZU9sWeE6edmLP8tnfCJaP/i39d5ym8y7mj
9cBqtnRmmyRJ/hDFaxHC2u8QwqX9M5sHxBusmSEBFp/ByT+38578sjrGupNU
xqHjUWR9WaodPkjU0dyyVCZ71dkvhDjntSTOVzTnvAt8J5H7Q0sC5E9WS0Sj
92GYhNS4QsOLMLpQM9pTBPUnzigs5uqSi+YEkGdSmYipbILu8Apcm8/dR/0r
+YJ1k4UpT+iW5KWz30+2TbZksP2mbdUyNjjBcsynEcfG7Qa+d03uAvtiyoZm
HKweZR47crquLX0jqG7SbD5q3H1tuWXE1Qfk6u1v9LgjEsINXNt9XnFD1kmD
JfNUt5THtgOLrk8BAouOWeKANU1Qe/NBSWrjeC8CTN1oiZTUXc3JNYiE0Mz6
pVnecPkvUVhw4sU9aaWIZuwRuToavlqscRI4FPFPnCQllXypnNrpWdVnJsm8
P8YdIkxfXnVMt9rhBO+niTZ9/3LzspcMIrskXT1wyDXyrlGSymAeThvZt8gN
hchNKk6M6pUuvib8ZD3b40kTDVx/AwgB3V0ag3AeCXxszuH65W+a9OoKFnZD
l8B0qB8YLJUGRrCCm3HrVCLnhmzeBG/FlJRp7jj5I28wfYWhSDnW3yX2SF0N
t/UliRhUaAtNQvyAP+kIaZvG+CGE4RwaEpSioqNXCfuIrSpbLfCmamqjbzh0
OjTrB2Y9L2PTzZ0+DnmWjMehVlwF+Y1GXII73ucJ9hJOgKxNa3lkti+3Kip4
9kk5d8BkSeWpmzj5JD/I05p/hk8iMp0rxKvLdTWhe2A4w5pIoPKgd42fserU
5ddwNGHfbYe02cLAKvDzs4G0JlxwpKtmKqftKjth238uEkgAAS0kEb5pP4Q8
7DlBkoe6RHT5WGgG48J4TTVk51prs4Dy8SJgoklvikG7ZWo41sM38GAKBGzQ
0icQoju4ziHvUhC5MKXnyHgPUmxXNZg3wihCq4j2b6stizdJQbxJ7DRZC2Rv
wythid0xA3Iy3FxpKkWzW3KMOnirm12YrPpwIegqULV3M4eVvf3VMwlfma7r
tUdwlsFiCbIJTHndNq5ZiQm+WRgj6hrxOtK/hE/Vk/hOX0X0GeDndONHXREY
oqlKXrQ8J8Ngb4jFPX3FLKnAVEtacMfzzxGiZo5zTvleiF9XlNnYduTkboWP
oocbYduaDUcbEr/UXB8s8vmIirliWTvlPBRCULu15x7OM0NTDPU/Uug09a5A
ME4py3vgpD09s0P89ndpV9bhvPCKzyImap375jJ0BinD8AXFRghlmqaOCp+9
E941ivEYVEp3b0hFgNezEm42A8O5WuvQ5b+BjT8UevIS5RrwR1mtwpKZFABZ
SxfeHR+VD2DBAkWAwqEowPg1oxilwbG86NoSmoNGGd1YO5WU/M4oYPt0HA7H
GuX8M4TbQMtAFi4O1bqsks3rm4fHSnxtlXrZKG7zHEOxxjv9H+5b3PPAT2J6
clmuuKfWy6oFppUiIWMPxhS22EoIA+/p77fofoLONF+ychaqcUIoe6Agf/AO
FCbqZUm0XpU3/JJv5CVrVpo5KV3khysAHFAp2fmHSqzFxV5Xebf7SoJnvlLJ
+3IbcjcOvRdaPDf8/+Wc641A903QoNSIGzf0vQReeQQbK7V4/+hmGm8KH8Yl
W48DRsQc0GjjMtkOQIrqtA3FHDw6dJdgHYWYdbpI0WJp5Sbx6CkGM+nwxCdE
LaVJR3XPF/ouUBNpLW3U+SjErWPRjVyvhqwkQc3YyMOvfpsS8MPZnw095j1/
viL1+ej+4zUcSLrz9DS0Bm0zLEXZH9G1Qi31eabJ8fy17K0RU1p0NxU1JLmy
R/zUIQZNzCuuax95jOni04McXGTeKdIuyPfoyPh2uIDHpsA234d4PU2xWEd+
OQpr7gwPIKurX8Zdsn5+ODLfBs9SDCpGw13Fl9TmUX760ciZ1pgTclu5qTDn
THShuJsIKNudzMyOKw8qSiOKtbKpYlo+4Dxwk+bN5ycIkoDahI7CYaF2jp/y
16yN8kd/q7GvT3Eo6WqtiHz/W1yCK/NQt3VTC5vPxEc0RJzGuXQfAqFq5AHe
+oPBndsf42LpmeockTB0md6oREfBHUEWRu63Eto9ipq+eTj0iRhUQMTg7BS2
4zgwd5RkODGz/YhM35+IYqzwWh03wQMytsMsdGzOUdkMZDvJEbCajz9NPMpf
EuVthDJjJZVX4gpXOzXkoMqJuWjnQE+XaMAwVFFXYwydNfDBgRMiCcVdS5dZ
RcO85xtskO1+AGsy/w4BbuCcpN2E6GAT2zmOyzC9Lc/AhTBLWSj+5/r9XP72
Z13WkTO1lRg98m9Hiipy67rzT3VM0HIUpgxl2K7iFirSRYbQOvEFmHRVxmI+
KnY473ZgQLFRK3/Z0uY6YtaGCrfj5FyYVsuzFJqA2cgXKsVgi+tSj5VXFtMq
qUfWfTqgr2r4f9B4AWtdcge2nvXZmg36uR1Nuy6+R96/+H1SGrnpqZM1nH4V
YoZKOxbsmIUpzIilFQI4MEj9uBsl4+dxtdvUhVxvz2ryD+vYM6rA2iDL2ZlS
PbsQjh+otrnBd6igSdRn1MZ3kMFYRirIpVNlL072iRMjhr3tDMGY3s8UiH8A
FwiUgJwuaGNm8V0pHldI5H321xdEDXXDYfpoZzmLXButcpLpibZ3vs0689rO
Z860UN2kp4ZzmdmiTbnoZy0AWACwuSl52RhZEGoElaIJRFYswFKYNPwLvZTI
/43BTbDqXEenKK4swFIrRS56g7lwVP7+9AwSl6kXZ5lEVVBExlLie5OU76yq
aWR/tJkjTUFxyTS9HPqHPyPOmR+zIKimK7WJ+7sJym1yNY5GrlQJ1MfHjjy6
LaG4TsrJmEIzV6MadmBnLlWOl7GSZKs3/XEO8OKvmHEk7uniL93d+tmo72yk
T2JQsdn+VB+Gw4PQu38QHwa8kUqCzbvCwE6DNYs7S9g4DfE8/+bjT/feMRdQ
vnhID5aAxPlaMPtTZJMyYZp2WBGpRtJ7y+kMTofWGB85Pl7sGYmb4eZqCWxw
kxyGNcN/PC5SiIJ+3ltP7APL7PV/fN23wEegaNx22TVm8mN+gVDVFjGiQQAD
5jYD1uQPNFK2pb7rcazKMC+wbl6ARZN6w5Sjo0tiS8GuBYeKxKsH/+pwLLrS
kFUkXHH7opFGxsy9G8sD3kjLVuU92JxNwb6VxmZlxGqOSuPRzUpGIc2WZ0T8
aiaW0Ye0NC/kxolU7p0R+R1z9wN8SkIP9TUS0LLhDLCqyIQKPYclIRS/fe27
RLYE7grX20xKbJwPuwszqoEVb6S8lf2g4IynhHy/LSAz33sECJrod4pGYVcn
g5Q8f1KeqnNZ2rQQmlRnufX50QR+IpFRUm3/2wIEoHrafwPf94Crdm7P+5om
XYUlf9C9Ets4Ddyf68j5Ni+mI8EVyolVAG/RAh3sE8h4Et8ybyQnz062OxCO
eXjIsf0845oacoNEAOmr2uZ+UcftOwk/hThvcJWFLBnMWdo/nTW4bFj0YjYZ
u95D64K94ctHstZ/f3+YfR+kQ3McDEC8ue6KswySGCEbKLF/4Ri30pQCVTG/
Vl7d8o3pJ6YSQTIDMcOGyK3hJZErhr4iO/iq0CdlyNHagWZRFy83y9ONil5u
9lzxhd8m67byYk0WgJmAPqFweO2KUT3G+kXJYJqdGW6n5N6DZcf2mJUfxVh3
wLN2Cy+LBzpeclS1kae0dNiAQN+Ynu4TtgWNeEMsQ3vo6ThrYcxEx5IbX9FC
JwgNBksiOZFsOuxwNcG/UmBVNH8PLb+VONVjtThKojTHhOaiwHEZbmHi4rY9
v4JX4NgEXzFZc3v6QsX28CGgTnnbitS6NbcE8IMDTEk+v6ZCHbUpqJIsqthb
U2M11IMrCwA1Gvn0GZrZ9K/8Xg9xQZjJEwerq2yHXxcCkzWz4YVK33/iGXgq
GxUbZYM38+MOroFj8Km4GyLbeoqkShaWXWW1VnqCYyDPLPAphKxf3KFwYl7H
7Guei8uvY0D7UNeEtS1kIlVsINU/znBdFJcdc3raVcJUN8jVgkXhsNrrNVS9
oFWwu+nOESq2zwLBDvZ8N4SKWYntI3kOh+PZKyX+2u46EgnKN8Bm0b6hbzrp
kLHsdtHuLFc7O7AHY0xCRgTgwoIm8KRJqpD19e7sIhA1FSCgmP0EnPgcpeVv
EIzN3LyLFQh1YhZfkFGl5mguczmmwqIFpj1vWzbpTssyh0Kkrs3rqM+bvknt
P48ihyCj1ESJsaYWqIRQjeNo/KWUeYbfTh9b7dOJCUFY3fnlGv9tvLvLPrBy
e53L04ldkL8IJSJ1uH4rpEvWEIB4O9UdLAdWdougTSnXIHCqKXcGWqAh0H4d
Q0qsc2mILb4BEr6jdnPR2gA6XdDj3AjfxatwJYwXUDyBqGxTiXeDli4yxg+/
E19W+zdh/hXyfGqs7/FuXXd8eCra03diq2GOjUnRKrEBigo8TcwKdI4o84Ts
MCAxpkg/Fcz41ODb2PZw4bVDqEg51LTh2ETUmNwSTRrAcTr8f+iUpLba/K3b
piFwsU0U3d61IVAjtOd/KaeFuD5W+0jCpgUlbZjDlJMqmlJvS2AJRtCMEQau
5QopC6PV8qWSAC3N1Pn05NM6NAfZF1gZCA+utoLj6zbjwTM40SVGe7bCJtjY
7/gD2tz7gmG3zxN1dYKKPoaeTfG7ajZyDJau3mUyw3KREJrCfkFyHIboZTs2
Hm3KIfA4vitLRiAXGN9x2MDDzht2/3Lg71H8tRw9Mltn/uWvSXwkzAWvVBXj
pbfRwrQJzzsSpjHUyHlVlpzZJ2XHx5PJrYZf2dVT0m5gWEYAGb1dGumXc7Vj
HD8Izlxn3VuMM0x3u7lNH0xuRXJ56z6fXIDawzAcPzewHFDQTZSRhgKvPcDr
BDB4rwzsdc2noqy1cCvX0TfxhChH0FAq5nGMgRIz9wiWarH5Zp1RWm0v/xDK
E0Tthll/Y3lnbQCThyGWcvc9AZqYqOmt7aD2J2ERjfpyJMk/iELnMuS7BV9t
G5y8SapShTjit60E2X4F8f5NEuh5+rejt0N6GsY4AErxOkplQfaNly69rrM7
jB0XqW4JPPqN0PM2lHplVH+AkopXPetuIZjfwriWQgZsvkz5a1T8DYHxdeuo
svGwWjwj1Q7OZD5HMHj9rnsOhY5cW6LNED0DT1tWIiZAha2HmYSUimEJQPK0
3i0yXlX5Q3DPbDoLxRx4fOECrB1GcrLWXErTaOjbsJNi8vYPdwWtcUdLQIpG
yS0XkT9qsWmOYeJL6S8/Kpxvcwpmhp9xRLY3ag5Xrl+yBKMdgnbd2h0Ibkoj
NOb/Cf4eOC1Ho8WAWwO+e2vD25CjQhzZZ67KrxkE7wk1HKPuF2R4F2Xw+4yX
vZsKLBck/aMScmbkXDNReNYco41oM/t53B0pQ1CXlIoAltiL43l4bnzR/WZQ
1NQ96svHUo6Vs1efNXK7mq+MylO9/jZOZTcNmjPJMs8iZJaWqaZ2uu/qBVY2
eV0SQwnH3o4CeEmmVEPpkKxK6NY99RTSq4ZcWAxyTh7X4vOkUURxKwJMrjEK
dcIo6wAh4ZfhQwDexXqhD9BnBY9gb/Rpm6dFuqs6EHiDp7ur57WT2hjF9HCY
ENN/GMYkuuSb5P6e9coV5dPC8wnlZe2kYm5SMD64Lbz3nk5msqEI7YP8VVe7
+byMaHSrBI0l7pzyBv34F2GzaWuSnqSIF+Kw4bgyj4t2g/TQJJ2aFSyMYZsG
SVh7kCgTerJN3GvgaWCwejJaVuLryHRSw6k6JEMZX7Ix9dXxU3IFDV8hH/Fp
1+eIn3OmFoxQ71nWREvln2lsqb9Ri8vgTHe2SxwYC0cKx51nRl0rc1k7IVTB
OH0/pPhCZRZGnX3xkvGPg9TGskk1YVxQ2XFeZ1grtXBKj760S6IdmQjPJEgm
diIKAdti1vnG8LiFmdah0h+zzEuzqx7b+TLqo9PYP4eDnITdN0nO970+yF/b
Yu7W3XKLYumwOrmmfugzMQHMgND1XExuSA6Enq6eqyS6MO6O76VFNV6qKWCd
eWVV1sM7vg68+cm3Q0N50kzxg/yBocsYa7kAQa0G5kxIdxs09PUsTPR/+DKe
LyKCjY6aN8EQCmErht0MiLHQgA7Ldps1JcR2ehhJxk/SOd6ts1JLliBJpsZa
O9FfxG8uVZaUkNY8p0Kw6XxTe302DsoxsEGZs5/Ful9msORO9qCllnB78H4l
pXhNuFmIa6jlyF8J3QtYFBOwJmA4q4oKMK/aFjtQOCtj04yafUvaq1oRaOfW
2dKyyJ+8RJ8WsTkLTdtnHRVgdvKIGmuY/XiW1UH5JH7yxMrl2ALd/st5mWJD
4Cn6PMgsf6RfmSM1ZZmi7IO3RFiRKIhWjl4Hjl1EZ864wIw3vHo/4DxGoQ7e
rknQ0uRFJVQconpGRLkbXyseXRxOm+zYZb5HAYLy0PYAj7J1abDE91koQUkS
MkA0Pv5+0aji3i912+QUbl2tV7p4sYvaV4CxaPMJq1vynHLThr4zmW5E9DNe
rjJCm/hs0sgAnBt9bVxas6U9D94Vw4WvB7Uqoxa+AabEGBQd76yJfbKz4/70
+lbXJ3tCoYabcM24hqMb+vze/MSyrULgc8CaJfdsNR+qBQCwPyVzCWkdhmcq
sZfp5K0sjSFPvYjAhazaDdqHThkRZ/zyEtVZsJRY1Qr8B2O1zj0pZxRE8/i/
A2HHeb9xc9h9n4OczNoziaIDOiQUG4/WlhPPoxd5hw6f3fpUYvVVg8uhpsjG
jP0CiJOzN7u9EV9Vzj8y+++R6r3SaqulDZul1GlRNA0syQ1IQmhPlwk+vr0h
rlkDgrPEC8JpuxH7XuUrFtytn1eekJ76S40wY6ANUjZh31kmLoVjoTOsYbp7
+dSc/9kUMlKoJkW9K+dJngR6fSXVRzChOR/Jc40a8HCPoeEUIOwWbzYnVPi6
kDWpl4fLkq3hUqS8+kaszYTY4BUOZ8SvVjQgpVq5LrvOCEE+16AW7zEPfe7k
AYsxkWwEMAAWhF4V3ubYhXKliDduag+wijFIBdFt5PRovdBeXZaS3eEY1+nw
Bcqx+8jZU2aYrdjzoQ+FY+zhGqzyBodUuU9MEwnPluiKEHarpdo3wUDOwIjz
GqtloKBK5mqiXJwvXpRq92TZs+maYg5Nb1MWnH3vtp1suwudJuvV3MyN8A2n
HNpEPmAeEVOW0jhIW2dJtfa4jnq7076kMvQBpVOmd1LD23qByOAUeg2FaJFc
zvQb+W1p3WLJfJmlGb3h44t+u/m0cP+gjbe8+Ks2tYoOj966Yr0cmYxum1fv
14d2cf30Y7rxBsMVjqgkXg+Mc2mryQQhuGl7f0BTXbinQqHENGrbOUYoyKmt
n7MSGLHlaX84O/MgnTD/22qxbvjRPSRJ8Aol4ycsG09DoHuL77NXrM08Qs8G
X8iO4MbWHHOyhtAERtrm7kLdndzPa8NwnHz7KnFjDXEvi7w/4tkmfbq40KBE
ZOBD+SwvX8m84L12/ybwaWKKbNU4bXHo7Kd7gYLa84+aH6gxZfyRD83UjS1i
ckZv0Y/02Din5DqYd9C+ScFonAog3h91tc/o7PNkf3BT/RoAHlUzVj7/J8yZ
YPLEX5iGHrJxIxcgn9LMR2xPjJJ0eBKIbjE7EqxxYD1eMORGxjQC4mS0uxHT
ZegmmG2biXzs3dPYgttyXRSLBjGw0RCaDWKJpyHY0OEaWAVK/TMvzz5Nu3Nk
6ZijXvCDAQdXTI1kD2oQ0m/+AZxBMOVprmsvI43HfvyMqYA7DG5HE07P+vol
p0xbkLAIw4p1Sm/ylOUpwv1SoBHFB1ORMB3yLuPQdTKGBIm11So9QIzYKhC9
BVqcMK4ua1KyNYEvUhPqnZcKIo1H6hX5k7EcJc2XZBPX6Fjdgg1qxI348zjt
lMuz6MzD7l56xkdbosK4qW6vSxK0nkENCx1TnWHlOESWOIoag7lMcOi+/rPM
i7AUImlYJVXKnSJg2UVlToi5V5rO0oEYQrqR5QReUrrbsnEF1gJiUEm+MVzE
Ek+eldDwgGeV0c1Jaa1/NdCeLffMy1ZUDRv0+06/6g6Q5g2yRriUTlXKyC8g
hdfStnKao9MG330icohpQPJc5StxspvnIuVE0dxMJd4m84OPAHY9Wnogh8sV
7Nk6xMPm9NVyJef1Web5oBsfDce2aPtyf4HKAx6TluBgqgbHFKuI37u4QHNZ
cb42rM1+i7b+nGAMOs9cZCL7WECqyvutDGqYv0iO5CyguMdRp61dbQQ94ERy
ooaCDxDFiIz1pm3biar+1y5n2ZV27nOVzUfZVOotWoQpWqEii598MW99lHVA
lPMa1tawSl5qLp744k5s0EMT0lE0KKpI+N69Jvj0jOvb1NnDgZQL9mP4piuM
jUEENk/V0KBo6akqT9+fqBXsPqd6rT3IBXUka10pj4vNgZJ8JrowFReyZdjl
aJ0MeOj936skF9COLQoujPJV91nBdoh2bFfr5kG6j6BP5g80/fIaXaLByM3G
MbYfrr3dRGYj5njptI9VEN+x3cjRTsIvx8lI+L4jOsfq//WNvwULNKf67ncG
0j1HOArKT7wRvEDA+BDqGvarVjUqPuITChnNjBn7nIL3rXzbBcPaq5k0Zm/N
0CCaN4zQ+KJ4GujdLJBKebSr7CcvRSqV9a0N564YV0jaBzpytEqpO7HDWIQJ
wXCfPHQ3nUrbV0UPmi2DMU9ejAKlMobFchetY3VOjFS01udJyfjrMjtKTyfI
h7D6tefp2xHrP9dKHFVmqD4l8ZqTWmRf8qGQsG2ugGRiT3I3IYeQ1yqA/Br/
+m5SsFSk5PXgQwJqyNSdFc8hq6+hCY1188cgUw3t04megQAv5ezNTjFBQBu/
KDySOIDuf+ocge+vkXDHJwY24E/6dFEI1mX/V3tk+lvjKmhcCTIKhPeonMNK
P3bQ975vEyUoFw7mQgmbcJoIUtpjrUo1L3M0z2OHwk3n/2gUb1gaEg6GWYmi
juFI7tkX+zlJDeDD3NWHy9LlAASaXH/iYmTw0D1E4cSxKBpgQ2xrObN6w5nc
JMzNZH7Ymzjrc7qHfk8JT79Fh8Qp8b7qg3G0MfTVFtlCfMW38GStx1RVLlnb
lDR3qeP7vzk7x5krYv7EwVbrArq5KK7A8LwoIi4arEcZ067z9Hbw9tqIXSic
Z19dxAMJ3iG3iX4lvJtTle0Lf+eYjuDdKITiFSEHeHF+TbEqA7fLqeQq0HoS
AgEHGZNMVFfg4C+/7FnttHx7A0CKQz5ph9MbE982N85T5d+rK7+0XwfxiNqV
z7LU/cUNxaj/dfKy1B37AC6b7s0D/LCVXt0smjrUz8ZrMmH2ux+LgTxceqv/
lB2KGyZvJCksjueAsLWatzlPBcaXyftHEv7ON8gTkEAS6coqIbymK9xZZ5jT
j4XxiWAZiun8Z+OzNusig7QwU+efByjqAjzhNpE/KF0VgQ7kw0+vwDETRQk/
29a6kbKt/H39wjqMbn3Syoo9Dn/CCOftj/Eo7up+FtRyLkkz6Rsr2RXR0aZB
4b28uP1Rv/Kw+0hmbzjvoJ7U0xm54L08o4llr3by9FPfuG1s7T4cTVztss4R
x2lgZ37NZovDmExBAzZtRd9KVDBAGtmKYzlUZ2GBdv9ZY+Tgfn1apq9xbZk1
QI/QZt/ePMyvzZ2F3+FBXwFTLO+mebwsW9dlKm1MkjST3kJ9946CiXkZRm4c
snU7jJq3MCk6eEOiYWt3OMxSx+Mn91nQz5Vb4YMVMefctI+5299HkuRavwf8
eldTNOZWlTziTx2AQ+hvVxxuwPhte6ceRJ3VMDF2fR4vbk+X/7UTkt1T4orS
6Z1i2GxQXeA/pZDFkxhDXvL9aT9omf2W+Ni5p3fMN6a6bctIor0eIQK5cyTB
nOxgOI9R6B6mr3TlSa/IlR5X9sM4r1ZmUUVewU69sdzRxzMOZBtfNafOdk2f
2GcQX31miF8TFjq1DV0YsqUrXzUHjFvcUHHeTIIIMnOusTDJk25XYJe5KqW9
IawQGx1zDuwr7hHo6sjYPD+V/oAV08w0m5KgPjdDvxXEM0FqvVDxUe7+iTfA
gEURAYUlOSbI5NzXonAXQakN+cbKhS7/WG5Z4D5dYK/qw+8Ken52Eeve4pY9
gpBNFmNTaXfcrKaU3YTDiGNKU4+RXFj+zFspBjP2lzzwvOzZVZDzKI1rISU0
w0vB6k5Dd34DfdA9O3IUt+F98FCL2KuxfqpZr6OYoJeD1HMcadkv8bOY16xK
IC02aZYlTsfS5qqiBEphLmrhOwTDUZp5XkHl3mZqjWqLkWLLe9sET0DDfwiH
tKP3spqIgaRIE36/PzLHzKexXpXnG2YOqNiIQN7NBwMI2BrUDH9iScMn8tYX
UJNHpUcfNklW76l2p1WCjjyFrdznWkz8Nnzp0pp4spP5ybuNpnHEtvmx31mz
oktc9xLci63kYp6gGlD7KnaW3o2AwUn15RYalkMFkP/NxiUB39ZA/iTfPWO3
qRmHY0jdqI7svHlEidp9X1zg9ABGPxd11Qwy4Jk8N4MUeS7ojqMb/IrkDGxH
tcHNSlHncCt4hBcnp0EMXZHjMcJZgTEOROaiH2cqfoHvTM4XBKkaz98DoUUX
DpAcjzJk79eB35pGQO1aG+jW9UD9lQHOxCwM5Zliktv5qJOgye6xntrgY6F6
oWnLVJHxot0dXkqMK/5jgW2NyS+kC9BToVKUnR7iREmaCC0B5ile1Eiklo/K
tcYDeAlKOYXHe2EeYv9hHCuuEKHoqMyguklFxV5mftkY+Y/MLhMx39SHl+j6
8phEk0CufY6vhmSWTEqs0iU6WRjiyn1MepBAsODYyvk1jjZ+zjoKeHp8bTKV
eO/cbo2zaH++OJujBz7ah8FANdu6/khP1yG6GbNFkYtjyYIlf7fwfzbna8Kj
nW1ybTzXD5dvGGv2LhM3ldTnVBdOof8g2ftLj5LIl3FCW2hyw8KGi/XiRWQR
RVtYfOnO2Mc0fSlUmkWgyg4hB2PpSbAE3LrVjin+L/fFn8TxIM4rjGYD9Zh4
V0WDJgtCo95NMzcVjB1GVVCEh+UxR9cw2t+6fQtTJXrn3zMTJtHAUFmRMpJA
3aSO2pb0gBE2dWYB5HlG27txoWvy1wR4rMrnCNuhTRk1D2LR74OrAw5c3XEw
3FZWrnxfFIa76Qvxb6UwkCSXSjdeflEElufhH/nP4I9nP7SwTnptDH2gqAS5
jX1TtdzdXljyDL27EqKyVHXvfB4xJOL12a1O7yXUKkRfAkOTNehs+RFTyer5
AZMkBXgErozI/74kWK04Zp5PnNVcEH6m/kqPYE44dbdOh0ufWpi7PYKxjKjU
FHPi5M6ztM1dRm59VLzAFSeUzEq8BSmto8lNTKBa2K3rGMX4iw5O4HV4Wz/A
g1apPEbLTFMu6Wo/3A9wq+NeE97LxoYsbJnmuMZT9V9VmgDAxZZPHukZgQnx
gKycGcVixnZP/SzfhzZGhSdZrjFMpLcuvxU2uoU2FI0e+XvxckVBN801iDnF
iKtUN82ZGmDhxtBC1CK2/71VWS+FHTtRY51G+l96NGvUSsalmzgPSdNml8dz
bmpqzldjaeSLX/RKGNs0a896sKvwPZ9jFhzxWcNdxBXvsdG1+0EUJDo8HbhP
n4b9EvhKHPKYmaEuext+EzTwHteBO7Y5CXpotE115pagGqAI9LW8H+wsEJnR
A5EE2mdDRrEdkGlob1M8f+oDhnktD1bgPsjHRL6gPYKK2qUK9ZVO6fwioC0v
+DKttFKbaeKZskY02O7kwc3o9R/DUfidQ+TFE8LXzXyW6nFQCglOK0BRNfCU
znw292N0AiGHEKhw2k/eQyaWnNYTkrsHBmw6s+2ffwc2f2imTlAHJXdjn7SX
sVdLDoDD/T6Lxl2xp+ByBjEvj/e5VJOTFYLk22KlKdtnK9biiQoalAmkf0NT
bNTEypBVeeHQgf3JqW9Te09yXw713ZBF6BlA5qDjbN6dm9uCD6yC2vZoGR5h
JROuGTb5oHAFnYmkp6YZX0YkHT2D7+tA1GyJhPXP52xr4g0Bfb6Y2EqH6Ri3
/90Xbq/B0k/C3FWgL2Oz57vMRBmQhhrX8zSUaxkUoxKyZYm+s+f890QfStVe
oSRqO5UqQUrFI1Zc4mi/zLPBkdI2ev8rcOhd1VXWcNnP5VhvaCN2U+A15HOV
R8wa/dcvy2whJgyX0+WPFV3K3lbPC70jHYe7AkkEi3uat3hKDzjc2uBWWDyc
VjfcUEDc777aS3KYwChbGjBiOBqu5mfab4O83GFXIIwJPuVmVXk/670/PpyG
sVLsQlrd0JpKaloP2JxbWUaS3nimOU7pH2002tEQ4cIjabml4c7rNSJ4gvU3
FyMFNgx/9Sbl+EeUTFpQgXVfb18c+jJXjD7UODrxXof4Rw4mDTuXzB+zdXsf
/fg9OQLAeimU4TlBtDqbYWRDbv5u6tTJB5XOXumomYn1gW5nFYQb5PAtnXUv
d1OPfpjg41LKy0EYSEu1jrtUnRJAGqRHUQtGK1BhpmWX5qjzCU/CIIdnaVzN
zCEIHK9n44PLB0G46Rp5icrRA5ZpFwZ/ZWrmnfoP7yhrwcGOci2XQVky75i5
N9ShdX6WBxrkb3tscCyDCaVxACJFTElY0MPYQAWD5a+llkfir+l+5QdyZULS
qKsqsDM3uo76N51QycdX+VoHp5cXYhSLyWiLI3d+Ij6Df84ptXbuwiG3IN3b
VDP2VH9dupBP+agdBFZkiyxcc3ask1XuAl5B9z3NNUEK73UMO1x0jQ/JqpKl
4c8li6mZ/iI7BTI4jbGynA8/h9dHhE2Hr5rbtRNMxyYdT2Wna9eOdfWNrfMT
xIGxWgHi8mJl+Q29NPUhKOexQ5X3jVRyMVZp8ku7CnKRvReymbkH51d/w+yY
gImBJ1EovaQgghRPOepX8UAmLimMroTpZ6qdIMFepMI4sqkETJ4GSGAiwNjM
fZl2Wg9xpxlkTws7El/eHILiRKPBk3WrVR1WyycvFwW+vVBxfCY2Q8/n+2Np
eg0Jjg3Ot6mf3Oi3czXY4wgBW3UHYRp5catMtALt2cIHz4yxEgsf2drPgn5O
GhyffYFwlLoPJK5wY0TSQ0Al8jZvTbd08wxbgUx1hhF24RMV8w2yPF/JzmnH
po1eEz0dgvedWWRMPDCiqV7QxRmmzw/frUh/cqGnCBX5P6lRGPeowbPCTf3W
XXsWc7hMuBdSV3ljszed9tbbg1Gkadb2SUGC8ZZG0jiEEQVkQcudyyQ4Nz6j
cscQqTzoVORYS1Sx48LN4Ko8Bpj6E94ulpaJKBEHzeE+KNuXuGmJE2KPBYcJ
yiFyBL1n+n85MmLyMMMe/yr/YAI37xib1BnBwaoodUis3BBCjd9XTa2mbHyW
MnGhCxO3+pArvUpNgy1JIf2nwMBhbH/qVdfFFZYTTNuUACdnFfw6H12N/7Ns
xOIE9EO1N/hLtWnLpoSidY+YAXaDmePnya7QSJ+xoW42HHo6KSXMPJCQedMO
tZkdYdYNp3xXmtAmpQlyfmVW66vcq9LB83SmLmUqsTEiXCH93tVup2kTJPHp
5tVmgDXJoUQ37x7I6Wd8vBjQbeeNoS9eevuT4Tople4a0imxziTaiHTI2021
/YwOYtn4G7GntFewAxvJVvLv8bqUJMUsQMJOVMPcnIuP7hLOenOe/RukWsxH
yRzaoWj87dVCPghO7kqvcKbC4OsHWH5ue9gMWMbvR2Bq57Z/olAnrmpgbJfy
g9O+zCqYWVzg4T8IVaGUxbW3DuTy1URqMAN7sGyhlB9O0CEeVFgZxHCZBxIg
Vuu2y9+XnVjGxNVDMJQVjTJDJn4SlXyOjNovGwDI3HS0lprrew4SMLsj3cdg
KRIWlWuZxgAwQPUtKUtlKm06H0EL7GX1TFeAt0WSO1nSaakq371hTHNkrl/z
OV+3hxB/HLz2ghZwFbMBbMam31zn9ttehJj/4v2wNrqENoaN2zXRskQ3w47h
pvycEf5BE6NBaVho+YCf7GmtKTr7dmJRJ+SzqJ6T5ACq8ibGMKftw3VV7bFF
WWcsG+KwWfITlDyc0/q0VTKQtPHISLU7AUcte0lXNDFTroMWFGwA1LGePs/f
Pbgor7H1X7ghw4rdiCCUBNo9PXzku3AoC+kU9+xy/wVtjhClXbecf1AD0Ozn
rgk2+f4QWtG4UXAMv3dARZNvY/+xREkDotTnVaEKDu5EZ+wSGS9+VWs57Dj0
3gUUr67EHoizn7MKWLx8AZJT7HktBiA5QkhtWH7JhSr3A8Gipps3lb74Vm7Z
p7+PudguQ6QzDoeMA3alAJb3P74rFpWU8rBj2fLacP3WekeH0RPM1RQyh2dD
UIUIbMmlhHng3pnzTmDLzI4C5+z/JUlcbHTE7i/o3xEKAPNXoLPfhDOhSJ5O
cs2eBMwNeW/tDKeMOHprxJjx5/8ZeuxU3ktX12AyU2r73nxdfXem7riS3AwM
gfCa3PzQnD6sLQjdlLuoWQKZFlSm1sxSXBwxs9k/b2LS8gDoajjwujEVmj4H
98pbX6PK9wpjHNwlTxb6J5+Jbkgq+nay9SZo2Sk5rRnMu0O5saQGZJ20Umlw
7iV5hiPHPWEfwfV3cswAuOs7wgYr7wUoowYTyrL2oUX36iEZ7fr6L/PIgk3J
twX9oXC1eHffyN2sxSJfsu0nKp6NQvvNH1n6msy2grbTIyfv8W4ZyP1oVy7o
xrJhvF+3hfaBUXdVejmzpD5Mz91l9O+3hKRVgC1JqYbrJIxKBoD3hlqe69rO
y7dObGQd7UoKpUM4v5/T+N0igrNR7MivTAp6gvYCC5OHngQ7qO74JcpCk9zf
vDaMTyY9Oy8fG2c5pgoApAd8c96ug+BUIWvBmYyx7bhmaXKRxMRdcoqxUsnl
3AIILoNvMbDwbhtRBoOk0K/iarziF0KzEUrZMFyTDFhSZ9HUM8D/n4MtTGfj
0nZvafqtR2zIOO9CKw1hAFC0c1aMDt30KRdKzY2KlpIpfUkueFk22v8Y3GVQ
Xp/KZg6mgL/B/e7mzfLG+SeHKkqEZr97eJkibjsnx4qZwGJk9dxOH1U6l0E0
JzpLSbZL5RDBVIK+iERgv5ZkoRUF+vvXsvbWpu8oUCg9YwwixRrDkTq+7gsW
QGcnbC0oaYcDIY7aMk1myM1KYu445sm0+XS8dJdEQxRY4jWEXtvRKczwgz3K
XKWjVzS10qsHdeI4vtDPSCypbOArjKO+4OiQqttcEEhw06cXpPYkAEupYvnD
t6Hh0h+KpfkvpfiOHj2wxmRSrm0a9JiViSSm7Z5KDG1O6txRLLIpP57NYSVz
PFodzgS7x9HmrRe00KIepHpHjkgMbq0OR5R4hZjKEVlOcF82E+FngbiqWfXs
RPnG5DpRWRw2qYwH0La7+d1hM6yDxAVWrXFCI6R17QfPGZ/o6WGS3V9euj7c
zCsSLleykOsLvNo/N4P7sQsNl336CpORsh4PcuJSHlT/CgNTh9ptZkh9864E
zYLNUmoSDIfO5m+puccdxp5DEmS+GN8Tp9kgbunIrsHPoqN/hb7nHiidCFKF
YDjeNg6wcxUpkM03p3umOkXqkINHkVVhpFEPhEHY8beL/UoxWr4Z53T8U+wP
eO9QLGkLZA7l8rljgyMUCS6o/uQKSJGAXt1IyxpAazmnwsU21XRsNFOqW7V8
gfxHeFHcQJ81RXG+P/QHZp+wgOSoBSUwaK19o/cuP/h9KJ4pjZLK+0MFA7dU
bjvKHPJ0zX96VPleKqmDCDA86CsBYyiCdaUTOsSZQQUKmZ9ugbWUf3V0WEzm
OsuDN6N6lk1Qnfb1YohsRXdDMpjWci7DPu4kolLnZgJr7ZbZfIlq8rpZvfhz
3sytbPOOD8KIuD8fY0w3iLm85dQ4xQbOgriAETs0mOChcfhSWuyciQJ56QTk
UWmW8ZzV4650lt8BrXPKZy6mjSh6YWqVYq+bVa+kiS64rdh7IwTsQ8Mx0vj+
Bl/sTBQghr+Kv+Zjo2YXRrQ5Dr6lri04IhPvEt4rwqXxJYhalmK+DMh0CDi5
swg/kxk8ic1/UK9EZnjuEp+G5zjrxCcgnUIKlwyuQY8w2X3o66kFob5pYi3J
iLfSkgYuvYnoFAiS6hJ2EiPn969VsGSgzgw2JCenEVuIBGwQjj4YUU2KvZqK
H+MigMukdRchOaY7tJTqVzfuAITfP2NvquX1gJ0r63LbeUUK2gg3SADO4Ft/
dRlQH1qwwNMK4Zxsl8f+xo8SLKcfZKPXqdkW96OOjlJS+9IySAfBDACfT6YE
zUYwJkxBToWTV+H3cpyz3//sO5Ch7cCiJTk5GFaPjsgmx2CTHgm9V66Ga9My
J2CbQgxMJ5J9CIa8cqHc55kaxtGjlKWs5d0IEtgAuZII6rbGxDof/Gqr2SOb
bEysLkj7sRWNQ6RF/owq6q9xJH3QdKWgvVuCNgFIZq+EF/2YZPl0kvArSSep
Y5eH6YVawqejmw8L7oSaYkF3DqGatafmDaKtlb62JLpuQ2D3WgRd3DUN5wmR
ri1f1JxmkTZXZj3nhrRO0u/VS6OkIA/nC9L8bH199rk7gDHgde159Iq7h3JW
YD8QzndT+SwWJIcMIRg+ueJuXBChnU29yJix6m8cuoLEO44r9HYQEjtDo4T6
gRQqk+4HyZzmOdV5yivTkaAZFCn9JfDrVxIqYdCWldJK9l3Kq08+akLqrdbT
L5OrHabOJugEf1ltCU/arU/T7858HxmXnyyQD7wM241m5MRSbQnoS6XQaIKJ
dmV7fq0Ec0NwdsBt6E5coS44lr4RUKNPSWh1UTcKBFEBmLqwk28r3sbqL1p3
/0MfDyvANMia/HIfCGaqTgpBq8+3BqBc3XgK6HAYxBosfu1BThn9+dAJ1RBG
U0kloufIRiQnfD1h5Fcb1J0eyoMl2NzkribU82grEJcEYGe/JyXIw10MeQfV
xxbcedbXpLs1C96VQXSrfzqrwo3LZ14KlDVHl7xtaHGxQ78kFWDj1/VLUa/Y
z5LifEVRJyhP8bml9CdBz0u0lNBFJVHRMpnSXfssVrsmMnkjUsxx+Ne2aqsB
1LDB+oazjfrAmm819OFNJbY96b8ohZLn6dJy3eVVJsXGJn7ZMPZ81csF5/hM
jgdFQmD3hOHJ7NR8N5tJFyh5wQB+X5V91lfMae1ZnJqkKt6Y3CRIBToettnh
WQmRG40LKcx1fwA9pwhbMap3aHL9T64Hb/c8GDDPPy65WXaE0jAC2WqElY6x
xVOUbzMrQjjQo8sYS1FahKOltCyJLXyphFCX3pzVyfsHp7ARfkSuwtN/JOZ4
bx2MMEYu+YHm5BkzFfp8thu1miEMoFMXK6p0xS8u9o1hvlm4si9E214CTpsO
D+SLlcoQBnPfjurz9FgJivgF/8oim6CPvgG9JeWfLTAcYyX9K3mwaJz2k43T
seboGxdzfZj0zoqL5e9mpVP5v+lbevajk06aVhjLut1McKCbaXZ4Nz4ItooA
YFn3HEYZOZRvhBBVAJ4p1kE3l209mam5Po1rjdn37pgzSY+44cVcpCElLGfG
wPe0+sZJ5l3seNLRqj/6XK0vd4AUi1DL7Jw17u3Pi3zGeApGkme1VGrMu4fB
ExxbuPMb1cghU6H+2BTMKoDIOeda/ys7rNV+XDVoSJelOVeEKU9TLuSY6HwZ
L1g1AFzESHibzFVQzUe7idcOs20HxiRgqWs41pGj/phEMXYF06CxH2YMOLKy
/OCcWWjm5j5qvomLadUKA02BSEuJsqCh0i3n3dpcyk03w1nFcXDcuMn2pUO2
OESl4z5U/7/rlVSB3FDTSplJq3VE2+6fZWfoloQd83s9TrEEuuc6hOAHpmWu
t0mo/ozBZXhEuVVa3ql7SkzTEzanyvD5l1gmEyu89hGl2fz0PpyqQCVukxF8
NwFQfeMtv0G9XNR5+gFRFLo6ter5AWnfPt6vYu+xnCuWqYcGMu/IFdYtcFqR
Qv5LEG/v2U3PVibscDXitd/vvvec2bhprpeUo5qZSpDKVPLl/gWcnhBvr2Wl
jXedLximhtfk2J+FiSjDgFQflZdLt+OtsQHFDr0JQ6JESDmO9UTfRhVhU9sL
JlnkrDdgspteyurcimyQyrYvMQ27wVjd7isl3i6HXcMR7gbkcvPw5zeAsUHP
mbaLlbDNRxvNOrliRzKPZvnTK5pNnTDeyb6d1//UzHV8XObkh1CkTQm32tIg
GGtDoUmqpfh1jWSHSir2CwpfrR4vwJlxaMBhv9IYpv1MEHzcmTgI35c19HGm
a9eF0xh6qkwEMUS6UloL1rMdq03HF2CEYVamfyHZ7k0Dawvk/17ZvecnkrM1
0xxMHRHVd+eK67Wvshkx6aYcF6zUY9unFfNBIJlHp8kvV3FBee0UxKqbmQeQ
cH/zePcTbGGaiKjBlp9RNEzMr7m7j4m54WHMc30fL3M3N3vMD4bo8RIs0CtZ
OQS0ZdqEWkTzi0MG3W80dK8/R87o+JKbrMlFBXkWaq+GFPAnFv4R/2yqwETl
tdvqr/co6j7EygW4DgiYd26pLi5ki0L+Z0an5UfcGu64aLs5h+SHwG4Wv3oW
k5D0VZhhFtBVBneCMhTqSM6lBR8tuVo3X/yH/90+9fmqMH68YEhRm7UPCiUF
MnnFjR83l6CyF6q9eFN5rGQXubK/ktoTsFBMv23CNkml1BFieA4wtmZ00c0X
e/l1eMMXuBsdrw4zCWw14ydJRAHRCu0Tm9bJmC5OINNn/ob90F/MAV/HeRq3
0IWpDLmPE/4gxxvmNxBnTOsb9xUY0JljAOrHXMqtGj7buEc0E0FHJAto1z2d
K3NZZ0ZTJ1pduOfVhBmpJ2ujgzPYUhVyT8rNftU8f6iQKRvM7tHWTeQeqKQE
p0UP2epZUItSIzAX/u6HzNj+YHJeg3/YowefA5kdOePMtS/hKMMDBqf+SIAe
WT9pjBvP8MF+tgj/fthDWRnKGwyTOztDcJ66QsAgMj7UM//2kkkOXyVapTMZ
uoc2PCnXPfLEVTRygJNTWGLNZ6YasqcpdF6JRe1kT1A/pTESJFN0vaB/XFAg
uAH7/Hk5pF4ZZDA/HpITjbiBo5NjwSWVnw3TDOSVz6uFrj38JLtvxMMxnHrA
PjL0Izly05ABq9fmMFwP+u3s8MhfA+eNUk6lOThqlBlY1tztzjTGZu5AfZp+
ydVQJkRq6VeJsdblPOf/sajggg1a/8vU9C2sEiHILejic3Wy7iYAs0mtWySz
VXjS2qDTDgFnq11s2tsummV+Tup6Q4/gMeNw27RanxVsGnkVgo1fvk5EaMg5
H6Jfv8VLCIcpGIUb86jlovMIX+Qjnp64yKlU44mH2kst/SrPDsvZBrtDNUbw
r6DPt6Mq+5viVQpc4eFnv0qKrNZAjcteu+g3918gArACWzun3pKmKixt+ioB
kFEc2cH+qvOJoSpcAQ9f0jkIbdnduYkmQgzAjBgFlV6mo1LixNEIJTYeb1Bh
AKNIPINd2oD8UtN/OE+PBk7wxNyYmOeQFSKnRGvc5ds1jikGNndAX6YSrZp0
MabUfBWjuP8iyWqTIG8bskiGCYTYsqw9ecHWNFxFImVb6SofYHJk6vd/Xbal
2cc8cfE9mxWyDn9rBTj//wV6svKIFoujy0JzVY2gtSYnnMKa7k7ud71zl3xd
XnMcEKBIoN9Ez15hguzZNHZLWgJ+wA4XFjey2XACEXuD8XOBIcGXnAQ+xwro
j8WtfvauFCxDvXTSm/J9TO/+lBIKfIlBYxp4pLRup3eDqOajD/UUfs1338uU
OAqg4whsaLJxxjpx5eYQ6Tf2IBfQrdajf4mVfhLo99RAclI11xxJiC9N/Wo+
9hENxVswjxzpIKsDp4qdAFYFf/GUM+hTKkZqbie/OKIybtlsUPnDphcFgzhR
AI8m2Oh16/JCwkI08lhVedbjKsKOhoCp/TFmlIK3cCEJEW+y4gD6z+bGOfhD
7bIWE9uJ4IjcfZ/BgJ1bR4XzrPOtmn0yHZs0EImGJGSQp3RIC3fLOErXbXsU
AjuH6ZABv6abF9oHhvJ5ws9YDH4DpZGt5zhDB1SAdQ8BfsEBFoh9U6Bv1MiW
/249pTyILxlUMVDyk0OGU1y7FmF3LvldfSuuN1H71QYrcMblygs0XTehAW+c
2RjrOGT5KMD2I0gwVSFnP7mmFqkWi5IhYPzgNhlMs/H9GSI5z2MJ1zOTZLg+
g5pKA9/edGPEd74Q2/pPYdz4Am9wcp+uQ6n5A/L2R2ePTUKkjwSx7fLHnrJm
MH3TKCc8LvEnxZkV8hXTden7WHql/lFaWf/5VNcpvgjy9CtvKc3feXP1kLGo
aha3Qon0cVcQq3lommBu33y4gg9KBukyy+AZDJrcp93skRy2LGXDBqCONL6X
h5W0hrnH1fkxB77fm23p4C/ALhUNnlVu53j7r6EMEYCD5xRwy157PouBSjLw
fbdGvpjNrERET/mIeInJB8GgqB8ZxeWsOBZfatBHA/O8WKdbeVNOSkN+QD6w
9jPENGC7x7ltNErPgFtltbjAjsRMDZ7UP41iS1kiMkwlqAkVOzeSSAAQ/5XB
vddkTn3aws3WAJJTjGVfiPoLADyKmaUieavTNcB0KuESHS6rPKPXG89gNb/O
gbX3rH5+v6kX/Gjy2l6PBhWodVKSPxA71lcvi115TGBQQqoBcjrLjnweJwjf
smdeFd7G8lFo+B1SeQEiZFHQidA0hcbN55WKroZ9Z9V8l/cIuBZfTrkveqId
wWWDDJdDpGzQSsENl/7eT1ZB3PFPU2vOtNFVIT1YNVZ7NRKPR9tn9gQF+rWu
jtpopCSVZSFcmtRwButQIHfMc37xVefkME3hjPdj22Lc8Ljr4/OuEDoABKhC
K82Bxgw+0uEOAdiPQpfNMN4jS78zH6TbsLaKTHET8yvnvaYIrq7aV3nHDKSZ
VnQ5+WbzOwyANH2cxjrW4ZZWEUJxhLQRT5+2Pr8KP7Zv5V1UdWLQHaxmTFDV
qNHIYfcXcmb+ZgePA+Nk40BJyyLNxIBWXjo5sYzQ3pI75NvN3I8+RSGslOzp
NLhheWLQ11wGo6Fw8hfbFvhIdev3A2OlcsKgVg3c/q0sf9qSyBhay8V1kqB5
5P9yzsTAieDA/rMtKjp+3aEt+/5Vr3y9i+eAmU7napLHle8Wh/b8hsVnaFVq
Jso1riiNGzT0Un1PTantPmGxPAGEwY22lqfakDHS+99e7YFab8i9uCEfQlbj
8nguJzdqndS/Aq2lBzlzlGms0UClkK6rvi6BWl6xZrKtDQK+tpTgRQPlioAH
WM6RqR45yjnwkdSXAfQTUv+b2xYBCP54sAZcGKde55eyxsypDEKEA+FveMJm
lWWSn9nFJhCAngsVrt8zUntLoDyPwevBadTcQGiKpO6tv/YlMfbjJJK3t8m4
WwgM+EdR5HkooLtcbM26vkrvrO00UZS2+IOSaAN9beBimePeXQbrO6gLzAVK
+QbEhOOHpMareMFEF33FMNQNDZmcbFgoeQ5gGZG1Q0Whbay/Y7W/PHhRWyqC
q4d2AdWz42EWVFu4mZ74FU/u2CBD5w8oWidUNo+D/YrwMgzH7q/r5vPwxMQb
Dv2q6ugVRkjTi300JhzXlvuv7bi1D89/p9V7xOhRD+00eJ/xcOm9hsKtQiFB
Y2JJ+DoKogRN/Mxwv6GKyCzZ4AOVX8d33iMldF85418IWN9jBgStBGV3sPPQ
NJ7If/tNKj4Dvo38aWSflLVFjB3lZ3tgHrKgwgOJHwBrSfqCjGK6sCHB0Xdm
MzzAMT6V4IyGfUATtM1A8m76UMyvPWI9F9NI8Ex6qmwZ96HVaroDBUx0hjUl
WrThBdkoGf2Jh9812CBRNbTZ/7XZlx8FeOo5bkwvh2bXj6DFk14zivooGzES
5hSdHqhazLTu436++fn2xMAw52YIHpBvKNjD0ARib7ED857E3L+JeAQKdukh
BlisatjQVbcqzxwWS6MUurquN3TsHnfdWoHbAiRZwlm9V7f9EDIp3IPp4xWE
Ioqq3tciNiHulCGmX8KNg51xDDHVYOYSp1h9s6UacO68fvQR8MjjbWaholdi
GOvVS1Y3oxQkN8/hhXvMzHY9QLCCdoTA1Ouu/FGcmbroRWVYBuu4mP3AUFVV
ORM09kBHrJYJDZzogXWwd74bTzfIp7ssFph/KJCYmowKRPRXJYY/ZvcB5cMN
tibMkJ6qofbjG95yZJEDTWO/2MzFrUgmxqlA/tEHwxHnz4Ztfo7XPi2t7nlQ
Sa1lEUGkRRYm9eKX7D1tdZd0Xsvt/7y3yASSMQ/lCbD5YfPfUVr84cm2kyd9
UquALM4TC9B3ZIcEpf/bXfueB7OAwiTdKM/q704Y74TK6LGKnLhxzYIldiJu
4L+9poyU0bPISB9HiDom7w7s8gCS87iMs72wH4QR+iEqBwxzqnCxmmOtjHvI
9Ge8395ujHy8txD2ktu8tfz03CPZuun0xS66Z8NSXXncsrZBNRsUHvb7qJM0
nlfTXFwOed/FzAqBTyGG7lWMY6/DZX2XqZwDz0juM1rxS9KpoJZOK6+3qjVH
/+ELuXSGHW8u3YXvW7r5iEKKCDxyLL8Mv/vwvml7wkItNDDXMISW0FNHWV1p
plJ/vw4ykb019u0oUFzXpv0P7PeiYw8h4oUhVmF5bdEXVaxPaVNEg22p8Hju
TIrgRAoiB9zyWskL9wNw2LVRM4BdB/mwGgLvsaqs4PxY9ra5HD3lYoRKiIvj
J3GCoZXDHRCNJz1iUxCW/pOQ2IFT2LaTL8ufzpEQy+VPSbF+roYBugYU9rT1
rtIhYdx0+CS5yXz0TA0oFHvAZEogquIT9DlwIu+XQjC8LX9a1JipUu5Werf+
KRIabdIZ14AmvgJanmKlzZd9gvK83UZrpxA4Ye69PkEf++l0EChjxPOYY/96
+WAesmQbAHrlCJCKQ7EU92mhMm6iFu1ZLzNfVrYYbReN4hl8QTwq5qKvoLwW
L7gTtFwyksOUgsMY8jh58Bub8DjggNf2RCM8SkWfeNlCXGNE0Apjm9kjr8Rk
1dZe8WW/lkQnYmVYxbQvucY9ak7k5Uz0oe/f/xi72azOlArosqZHmZ9Pwu0V
/X+mOh2Q6IasPrXgOBOvNHffGkiJd8kHpUsCzyMZa9Uv24CehzqCXwZo+gnE
rv+PdeDq0UX284pRgRz9i+APebNkgyHb1CTOMD45dm/lhbPDWiXtfyOKbYad
k7xpY7BJ54Z52WDO1UK72fAcwZvd34lVZX+XfIS4SP7bM7S+oG9w+QnHmCNJ
IMFVGAYBQlmaa0svJ2FmpugPg+lK8wmCDVRaah92vRDFvoSWJsQa0XK3pJF5
e1gxkqsSIOgvDOMs/xwrzI3ux8kZ+u7mCB9R7WCGJsdYCWi/zH6LPQQI+yCO
GFZpqctmDhOw+IO0t6BMDgzKt++jZmOcW7a2P+r+kckckRQff52yGievJdKt
87ZhZ/sur5WYypDP7+0S71TXvVubBlpFtBvwkYe5bFuy6QJRUWIL+WaDpWho
VdQLIDSBbJpwgEWsUcxGkykaU9XCj8RNMZ14qc52m5FA3HdTYL+Xo0V3hhSo
WWHxsgRvv5bYs1hD1sbHEAh8Oskxo9KrXO7gB+rl16Ms/37XAnHkjpIrsm4N
opM7+zn1nIXaJICXRfOaPs/jOQkfIMKTMtr9rd333mL3antw9x0PSLjre9/x
KuaaUTp1tmGyUCQ+yKMN5b+GJghv1Mtilg7ulwrfRrqYoel/hNajsly+j2Dv
jO75RJFJ1Vt2k9yqNlBGy54q6y0KN7QqE3IAYbEYmfB8rQ1E2LWlo3TZi4fn
qgRp0dj30Oa6E5IO1w8T4rWWBF1WDemjqaQd41/lpztzUR4Iix4d0G5WWya5
6KCqYqs0UO5mfmD9GUBGjYvQw1acZWI2Hk6qBV1tIh8NY9rAri2ZICtFZZGS
MQKPuWsm+UdX7jme+IpH+gAznA/7Yo+uG8L/uhftb011x1B5o2kyY17jHxcy
/UEqveRQiWyXjTkRokyvk/4ELhmRHJCuX/0G+7Dau52+VzdJVoNK7j8k21pM
BLEiEZM9J8wGZ2EKRn/BHlRctTlrRXOTnAbQokLwYteV2oEb5PTldE19oHcs
hIq53R2KKzBjK7TQYtB7yvDI4gEXa/puLv4mdgkYcr7qjNQepo3iiacmKYwc
jdRYXJ76SZhX6rUaX5j4qPLDnBYq/eZ4m9nsKHOt5/hyzAZCwam02zmLjI7z
PCfn1FWWmiXny/jaNioOrNxW/gsGhehGsMuBuq43485nD3jeyuIYte4Z5G4E
cnuwUy1mXb08V4Y0sLLsbkvG3LcLwQIgZy3qPHAfok/Kw8/cPwP5aTXb1FjD
INV77YLBjCJqtTF//jil3CcjoMs0TJ6gdQYvSfCp3NZ7Ti66BMD9dmTQ40Ip
c1JGRO0ZvT+Q3v13ihme16n+rCDyANPEt7rD1XiAnBb5IfV4hNjL4od7OaPL
BTsSxnOdpIUy+y2Hq5w65AT9ADgeM4IgxQWo3g6qqWIiC28ssWvaQVzznY9y
Agli9eC+JR5iCr1VKZ1FFQ1izNmfQCtT3AoBjp/woJ7Ay7MofJWPYYpJnkhc
vMLNiAmz1+wV1+gcTCwUVauErVoyRH4JBp6kKr9LIFkku3MFAXnZNYhZb5tm
CChF4em61zc+/imLP/caKh4IJIc8aZWOiKmOc2HFQw4/34Jjv7CjDuhjNJTu
rivnj5HQaQcKQIzK7QPakLj9BzEJuF1MW9gkpcvbaYE0z0QOddkrNLp8Vj/m
5XuhUtPSehfP3buc0WQ/A83lqc//CsiB4VcJhHDIuqQd/5mSlXuk36Kq1ziu
edwtuoe5e6XgTZ6SKE8kj0agfUS+Ip1XrfN2iL7b3Dw0t5pF8uJqs1+ycZFA
mfyQMoIYgLEW496Ime6ggQLe8yTZcKGRlYAbwrawJcxBf7BiRhLUC6yfN9li
i3vUXUsDJVLFmGXnqU+6QcSQgt2n01MqrACrqgj0lRpET4dglXa+T+ga9RGj
9TxILEYcEu7/PpxDWTOFRqw74yIATB12EG8DgBxQQPJNWyKCl39Vf9fsEP6B
4q9nQBONZzWgsaQuHvv9DRYR8+mQP/ixpv0YGdXJLbHq3Ytahdld0oXH7rRQ
S17PfVHfqHWOMrU2OA2yXdLbeZze+Uj0O1kwQNNgNaBq3YYLOAU6Rhr8SZiQ
qYohbTBiv/FanVYj1pbUhFUEv0f5rASVCPPxGa+jzTliY7Q7669msBCSxEtq
s46K0IgedJc1mEVRWaWuTI1TQWw2OqfZLJWt7cWzuTtvjO+jLZSoahwp0OwP
+HSBuuFif69Q8PrtHWD/E9rRxcZZS9iJslV3VsEhQ1x9W5Nk6rAUhz7JKbDj
YHCxW5XUce50tvshnp0M6rnmhk5vq4ictOr6rH58XE+cqYfvkD1SSO/nLJ0D
3hLYdAisuWCysBsShZ14oW3M0N+xTnnlBnSlov1y5uBSnvsmg/BYzei1aXT5
IqKcyFV+E9QF/GY6qFjmuil3xLKfqlaW6tLwSWCKy/xw+yTyAIyqBtmyK634
/nNew3Z/Z1nDZ7EfjZ0HMBBXEHtnMUGEBc5jUhdAmKzfJheJ5SuhZ4RpVohK
rIFxVBK334G1lrfDvWxqiTrCU5Wc9uE2O6F6IBmLx79LkeJ4xKwy4Esw/l+7
Ncojf62Qh6yKLG0QGGSaCYNbSWMdZFCi69bTkBEDtWkBQowblM4jdes6DF1y
rY8mLYJsY8DzFXpYXK3cbf8kxUtyiZ5W4HW6eVr5R116+mp+HTg4xFsPk7cE
eHPWcotNdz0kPBxQxgODo91OfWbAQh8vkP8lY1nb94HADEgeiGFQ1k2rfGDS
1e+o1K6YCV9vbMi/knie9DRGgAXynRH++vNuXq8Num7ZRffkRDw7GRpZ0SU8
/rJ15g9+lwxN+fiioCH1CCIUK7PIwZsNGw1j5f1Os9rC0wvd0Mex3b52Logd
IdOKDuSA3uIuj8SXKD13X6N+rU7sryJoz+iybLxGX0SOFe7pSVKYEWrOhNoH
QWJw6oDVkY0H7VU+VUTs7NQPPksJ3BZLiX5vuDT/Ro42nCq/Y/UUW05My9fC
n16Nt5uzN2zd7rWV32voWma7Eq4x0+m+c9ZBi64sZjHATV6zy28AhjVZSNci
WHuX8+u2CfK18bIxGrw4XuMTmrlurWzU3H8ZlQGTis1oNo4BhfdRZ8iHJspz
0bCV88z/5kjo0txMIQEGgdFOqrJWp/2IpYQxhHX2Q2/gx0TcAeIiga8YevkZ
5BvqOfzwCy9FELTB6Nduk/IOP+6Bld67vhaHdhPFZUm0LP03Z2LrTjf1HOGx
VD0W/DqccskR8HNlPJoQOR5KNz3VjnmOmB8DOI8TXeITBVvdGXII1Tr1AO+x
ZceYDsjmas4CtPlhgpe4t7+/9GbeXz8C1cVbJgsi6LhCniay5Ch22J1a4tIb
Uy/EJVbsFVIO0kwIYaVrd3oFfRQ3eBq+WgSSJHBxEoUW3twNmYuXXpBsKWTm
ayBqBiwLQSg7HJWhHnAioFjX1ZqKJPKU7J5XMeJMAxGT2kTyqL08ni2Dn89V
0qJtwixqcNYgFITNZV5LtrCI/Fh1UHuQIotzRq6qWS04I9lnUnE5iK54Bx4Q
Be3uWthMd+4aO8FqwbLkIixlmJp6RaFeiHcwBJ4ZeVmTRZA9Qkn+J+ndYdxY
AHYIo/LRPTnmmjyL+40u7STVzzm6LybqGND7R20jG/spUKblMGMr2FE7Lr2C
ZN9JHkbYOayiCUOoc3mBOsd9EW0U2vAjoHCW0P2bEBON3T3SDx6+5S+rg7Yr
NrrM79Bs5sLFqtUDTJiAs9IUYwmWy3bWVoEs7sASa3wvsbwt8IddMReZ+S/0
FUAJ0yheINKjOsTeQ6bm2M9GoAd/AjIE17ZHIEQUEdU2lAQOShT6gTmBpsdO
ivIoJIQcDPUafCl3/OV+zzzEa3BdlmTqnlgus7ds+bAFqCr6wYabjDswB4Qw
fJ2ZflWf3lXT9zPlgHr7cwTy03ljroZT1xRbJ1BHVhJYlHhNcOIMiweWfkIc
KLfWMDNIHzRRmVarRKGLEmcVWV+cxbxM/LLteHTjK+3ZrzFIv//PhpJgCZD1
7IjUpQUCi9kIH8xOVHF1SqG1DMZBC6LT0K7MDqmD7j1h4pc+2Emqp5lGt/gM
KSw0yFdxxOieS81M+sf3uFJ0yDSqkkBBeMWnMq2wBQgd9+NNrkoATQTPNUfx
ZSrYk14gGH/4l7XXq2MAzfDfKwH6iI40l0DqY4ifiwmhXUc1yyUMta/wLzmH
/OIdt3/8+N+xI56j1wnUxo05G3NUKyIlOXtGDtsdFzKmqFJLaGwJtO2RzCrd
vi4MSU6A5LhrklCu2hYLKd0GFr52rkO0potQ8B+/xbJ/GJPioz3YCHPAZ8jk
LC026/uGga+MeuAJ9Avyq1Dv68344lgn2qFEVZpjR9BfGK2g4dorJUhHdT11
81Z++2oefQDaYa8eSfJVqxmyYi2SQMdGw4dGdOtAEVxvGO137gFHOKnkl/Ge
9kORGQGFyVYrVug8swTK844rZXuT8WWjqlyCR7FgoolTOInfzxb36ZcUuwra
GQaRLo3+tUlz5R7Adunf+sqNbcnSYPtcPAT94321RnCd24IJvz5ij4fy1J5J
euJUFdMCsAJXB6QI3bByVtSB29dMzDx9pd0MxG2hHJSZIU/LbOydarrJkk6/
H8tH2oxBDZKB5p8adoN5KpFiqq/kltkJW1svNZnlONH077ju84W1KmDlFbCr
PSp8uYU68Rgmv8jHh/SYBEXiO+HIwCXI4Miy+zEDFoxlsYvlgyFuCmxct0Hq
y7sB3YoYLSR6AWWYpDiS7oyn6522j8RbybGXLSEFa4taCnRZb9Q/0n08dK+2
cTakHGhxLH1Ri/3pY0du7WR6HfETRR/Kwpi8lSZ9jso8P4oXKHCbjTAMIzmn
aOo9n8mdF/ATUJwtamKW6v9MnFqcdfP+mYkXYUw+9bQYzglrAdfaC3QzVtcy
SSZPqoFa27agUSSlW9lGTa8piz0azVSEJkNsDKo5MRkqkW1VUS6MS3KUVo1l
8v5OB4svmqC94yo9sBoY2l4MhV3Y/GFCxJkddEeYJVes3M07TNahBt7Cpt/O
OPcxCC9LHWkgjJSMvXU768234VgAFNCnkilH4sljLhp1GaUetZQYDvJ6qbYJ
NUwT0e8XvdpE9s6et2bVIpushoINlBrJgY2RT0b1SHkA5UO9OGGgRf6j3x00
QcWp+8ArCUdKBIE05Msp8URLRhWVhmTgkA73LABuiu+68ZT5lcvMsi68tI4y
jVg/5phLlBMWaD2yQXSjNu8+yZX0nrQKSfFCKTNRk/KP12VoI53gsGZD7Ye1
pK9FzGcLMNYxGzd0yS8IX5Df+EZWEbAWUzTne7z/U3aAhxks/Vr2qx8RQonD
GVV6+igKvMZxVh/W1mefdQvzebHj0hCiYnoqkQszYibS/Zmb/A8XyJUJqcVq
zAdfuBq87+dqMaQ5GbTf9ecEYasMwcfLzxSvOxC2wIJQA8f3MhSjuUoVmZA5
vgDg4gwkOEf+gMOJTyR8o3Jgv+XkiS+jFHEOPoO8vr8XxXoR65oCCTprWaI2
KCkKFQXMsfujQezeBdEkMmyVPIcETtJAr4qpLAFLyXitcvVckJr656nZk4Zg
Lb6X+pUrgskKBaRPuuMwZhtJXJPX1TXQF/JH5ZuVWK5uudpMBuNKWtaryzhx
/9QAs9D/oTUUvv4E+uFQX3fmftJic+Cs6puu2t6+dvB66TAQ9tRjBPJ/6vAT
/kjYpJ7x/NrXEcUofvgJieUNLim7sFiBR+zKqHQyxfzQPoay9RNn4g+7ce3Q
1CZLTdHlesQcTmOtJh4c7SeUq9W4+1G1VzFqDBCFtRA47dcF0dwA1LYFgEAh
+w/wu5zaVJiYMY6sy90kNIpKYumnR45uITvzRb5w0rZDMuzizohSn20/Vp7V
vs0wnRY0a3TDMa+v1qJjEjA7tVRjptP0htfSTKkzV70PHWNno215nAO1GmSX
eAvMJE9cBw+q3oFYMc7gyFEoGv/po8jedEjdHj9dRv2CMAa5IY9xMG/r8tFF
RXjHn3vv7C7Y/+gdq7zq0sKH1mHb0g0+O7BthuCThXu8MyK+CXCk4aZpiMoc
vXqGhc/sDLJJx6WfKkrxtMwpTzKoktcH3ma1sbtL4k4W0LA+rIX9w8cXnjFs
zrwdEL0gsxbPIU2lLu+ki0Xwv3IfT138624AZOplh2zRYpEyVQl1Cx1PRM7M
yZhtcjmbpWKY3LKLW+u9F8Fq7/1IsccSLyOKwSOgA2bMkbFWnxhOGQjq5DxG
MAe/RqqiM8f/gY2BafnHyGaZrtXQMovIoS45FNxXZrXrdi+1gsNH+veslAEa
9lspu82USODZTURJSW2g7JA0DZOj9nVPE7jQ+Jus7dvRU1WbGvWBgBBs3DLi
T1b/fY47G/si0t2XpdfgHCJxAXDDeSLZQTddr3G4YoUFgzMeN8+Wg2QT/8SD
E4ETx8T3MYvkEGu1mpe56s1m8F5X5eMbCeUjxcHQS8hAnhn/TRP28tfNfUDe
c6hE//c3S+1HkujbtA63GDsGgZrSHYQinr0UjZh4oYpICCmZcxTcWgOXdTA7
SnPaSDPq16nzZOwlPy+/u03O3FOeclaAl47Ovz6Q2ZhmpvamURZMAJ72yOio
kaY4hFoD/bN7FM5FgpdpotDhVSQhtpx1MupHB0fvYj4k2TBd6bR70Ip5Pp/C
XItNMDGp1p5LQqbzlknwE3cuGXPTshhJJpuhsKtVbUpPYrZCdd7eUUem202V
gyFyZCOmwJPiedMh4VXZbg9ujpVDYUKxcjNof++2t7HSvM5JPuucWIKbno2D
aSajTEjdJMwr+wLH8nK0HV1rhQjIpzy6sEyHKJ4ShzBkcmicR63gMudP+f8m
OL011QoUzQDyUdceD2OVg06djaEJPYZnMPRL04zbSENNeVi/43Kp8szfZdW2
HHDpyFN/d1s/LmBS63SCSjFTDMnr2dsD28FxYMeSJ9lyIEXKnaH1E+NHw0HB
1TrOsYA2sjiHqULglAhtgE/K3kaQnTmukKt1tgJfhXXFKhwYMMDeZltWAA2i
IGpl0vq5CDPVzOZui2lx24a0xVHYzmsggFT5FaGR+IayfPLdVVJVkbeJ4aT+
/6S+VWevjhRn6DFUesI7Gfb0kAMkXdYeeP73n1d+ccyVOBpD+khVl8EeLODL
D/P3Ppdzz/4jl/Oca/rHddwIbVgBFJ0QyguVHlUeUWeGMRNu/McF36mqAizb
bVyRcKO27JD0SkcGLmcP2zRJBYPQvqXAh/lRUfssScmQbEoKyFcn21hgqDaX
vSteyQgvlzES3W1Pq+CL7snnFrXFuRaLFO5w2Gtm7NqL4fT8AjHU2PcKeW3c
5VWmjLSq/4gvbruZbeSHXd1PpljAPY8uVsBv5DYlnbqeRQhr7SmSeNEsitcG
q3GcOSWdEL2knau/sWgenMz30Ab5RJWyyLvUU2lv4iZiw1P/z5Vjr79ikRIy
CYunDicg29ucCRowEb/dDN4zg4JlURAqUAcKAdo1jYBrPStLxc+c2V0lBt4g
Xhl+nC5wRAuv5HkKOXIkkkQBqz6BhGRr2/hTR3y9d72h+eFEUQnHPa820X0S
2xrJtkp8VZZiLsaALgno7K73YLg7g35sxW28iroanI0+aSf89jXEOodTiYg9
aTpFF2BykcALCwXeF+tJVQo5n4JtIgxA/wUibq1s84yHfR4QCuW2TSGvExvg
BkQdtkPVVtAZv1efE+4M00Owqz7MOiDxOZgNuTuKDypRdoFuSiiQsRZdYK26
1sf8mfSAJQED6TdzeRuSuDnQ1l22I+yX1rA9XsOt5ejUymCAk0dtSSjxsCrx
y2ltLRuaqMLWw60GVXULzorP7VEyX9YDRnPO7vKJ0oy/OBehvfknaQkEmhek
tezZwdhSv7mN4eCxDCv48IwZSTqYmBFoF4f9qdGeTCgkfPA09zd7xTJFHZyT
E1APVKug/k9LmOX428d5bMqi9daZUSUa+c7Zd7K2M1Oux1sBsW9jxQXa8Cp5
as3XY+uF+KIooAWQvCRzGdz9qxqOdYJoNlUPVsOypAv8gBcIHYdCw2GZPkwR
7kc0yfGHHv2dU0EY1TAnn1UW3EqBKVVGzAtGXl9HyA9AlUNNIk4lWEbFOlcO
oVP7yVqY/GK0vPWZ9STZYW5cQY3qtqh8fJtl0qkFPcb2cNROlYgHjwmO1SDy
Gs6DX0ZK9AziAAXpZSvp78gTx9ZWPZHrBSsy5OEQU8GWU9KfFT75P8gQ6A9K
T/R3zK3+l7l3tZ07XP6xVv4D0+v+ZZmURYgchIlC35f8bkLlxlzzPZK+msic
MyeYl4D8YDR3ltpOvqpyN1LvKjAYYZuP+ThDC9j9z4z/xFVj45mR3un5+2+H
jZG4OjVVqnO8lQGFpkF8a51su5MhF/sAULxh7C1g+T+0jTMOzNIjitaHbspO
JEYQxAbQKPA5UmAN2qQV40FOjCh27UBSSYhx+KhaRMzpIw82qYBBQIPTwRLr
P457qkZac68Mb3nvOACI12Am93qsR7iQdhQA3S/LKG/NyY1Y8OA1juNIVZet
Aww9zc7WKOU0dkL6pqzr38mF8ym+H5PjFJfKljdw4glPblc10GqAMaGF6FpB
etLwRRdyV50jTbi070VmDMPdYSzqkZPRDJzkTScm1dFXoS3eCS/HQ0CcV4Kx
DB9RyrsSTTt81r3Fib8NF4Va4+vXn5tCcb5P7wH4ngmVLaZlYeBVMkquHYs9
nYDSSpTOcpKN0XcK9SGqrBobszBVGg+FhSPMTD9swMabXKwOTVEFAnVS9/RD
W7uoNETY2OKGN2gS3f/nNJq7XXlR5VkmxJbEDsK8WEUrbptqh+HlogzpIThg
dY8OgbQ891K3AKw/zm4YU/S3G+5JnAOxu63pOvqIiFfW62L23YoLZNTnLnH7
p0B4qcgULUL0fs96+TuPRX6px4l0HVwf2shz2xH+PZf+F5SUzYRNsXQdCvv9
whi16uOUa/ZLAM6qw3R+CC9Ng/suOQ6DwGo6rl1Rjaq5rtzmOUSKqrGsUQhW
gI3cJWQpnAdAgkjR0KLh/LO7K1IKLQjUp036TBheOy2Kc7f7V5VdzHOiEkFt
TSxFCU+pnF0c+nUhHYVsNfqk5ph6EgaTGmjYZmbiBH+o+pVzS/ctkq7gVptz
X8UWjacHN1N14fn2YqdZ8RdV2EXLh6g3fAk6uswHUnvdoLu6ROiR/E30/a0g
F0dBMYDNz0uBpQnXBBQATq//vHw7RD6sSQmKTK9Ybf2j1yOBzVCui0Pg096N
BLZG1ge71lvgyjjpQKEwjhNK1g5z2Yy3MDp6KccO8EZljkK6jj7pgv4Sw2J5
6N4I0P2RzItJzIKRQ4QZNm3royqMXnhTy1nDT9TK0rTLPaF82PYMCXkBajlj
B8+6h8MTg4lX2gQo2LTzi3LmNa+ahl8OTCE0fxJa3F/y6K98C/7MgkorvB+u
MoG+AVTPgeI9c6EeUXI8UkpaEo9Fvw4062s47s44Dfj6FsmbCUs5v25pDocS
b3QC6jJDcCxgRmFJdTSfjKRTwyrH/U0xShQNvRUpxTz7K60Y3Uhd/YS0WZqL
YbVQdxvibUuk1tSdOdlx4osA7eJgBVKJOS4RXF022+B1KW3D/2cFFnSevaQS
Q5GPMmT3aN2APTXx9vgYTMSvNQ1TFZYB8cPQem5/8mbSzHNGBOODOlVe///F
Vbpi7jRcBSxj4OhRNCS369wqEcagHGGKCtZKdG+IRUvvuKrZL/J3wVnWW6fW
07fV9aInICui68Oo92gSubq7s5fCICX62nm6G1HZmVxyKDzZi+46cWznzAbh
BLqLMydAu/eJ6KcSn3PQkUMt0mDDuB7sM6r2eTClAVN0DOTRPKTXl3qI7QV1
TRxO4KzxAom4BjLNVlQ1azva3YVojnZRKBu2GuDiP2HV9cH7X+TdM1OrznNY
x2huey+Hg4lK8maOf33HpJqo8GfOhCSsEpaZWvlRPK4T6EhCHsMrbnUUbp0B
kRdPJDxoDU0tuNU8aSznkkMkLewtZSfCS/8U4n3MbV+z5PIbEfN6gWLsx2v1
nOiKTnMot4PtYKaNHKjY+lAqK4ZfIISDM0nmJbP+oESyoQgnJ+ul02by03WU
w/mTPhl+bLhcbfB1gCBjMV8XPKkbO5HX0KGZIzwABMoaNCV3FRtD3GF5KQtZ
Z57OhmoNXm6H8Xd6NNasaDol+L+Uta4KvPo9m6tFT3OkTb4cPRUu6DoS4a+b
vlc2OFVmB+EFdEuozId85cFh8/p9f9oK96GP22l8Y4pQLzvM6mhLLp0mp9Qs
p/lgritDQ1UqaackCUqgqhXUwNhjvwSNWBGrjhQIIBiigTS/6wez7jO4CNu0
lPi9662v/Fdyon6UYdw4CvG6paCdongzjNYk1xk4W1m7pk4PRas3rBFOrCv4
iI7BrUHalJRtfSQEPY6SmX7N9N3fW/Rbt5RlGgejUtfYsjowDil3SKCHIQFn
ZM0CAc6jZUx0O1XbSagmOFRw30cqYGYi7gYy7FkM7A6ge4g95cy5LCJy3xnO
WmE8Wr/qbazJ0SgKIuO71l14/7absZxbgCw9a7qdb0N79w8K4X8oFhtn8rIs
uxFxGpPt7cTiNoYuHXQnBNvyCu14iLsvHSAirrrIt0v93U445nc0+/7fzrAY
BLC3XNNerLm7+zjoK5aTORSyE19UESjCCz3vDpG+mavmBV5fi0bjwp27EKv6
OJPeQTECI4jk1P32MXmAhl46sfu5DYP9wPyvRG3MNwRZGWUASb20ibhqUUFc
qZQypTdXzpyldq8ojqPrnmHwwzEY+l4MU6OchMQrlo2MbA0BglnJ0giYj8Vc
umMkMcN3V4OMxeCwM8p6FPK8NmizXR6+xBbCXlXqCtVQ7sD98hed4aNFGSyv
ofkJ0mIqLAeFRGFWg3WrawNW1jjCThTbMgKcOhBIuOm3fq722k2knIeXSH8v
vaxRQYYSimAxXWGR1EQItCzB4mJEm2f99+B94ieTDWqJ2ZsOKeXc/lIABh5a
wtDFM6qsBd+O3Qjj2BHOxdB2xM8JLScIWqK64sa7/QdBwXkT1jc7LvKLveNJ
ZUSMIx8s+RRLuoTg+ETMOPCRcaznVXnF0wk1IwXs4mqHBCmVA5zB67h5NjP8
vXAEfeq3ssl4GLm0dm2UMAfHniUpN3Ruvz7+8NpOQ+hnx28sYWY94hectjkv
shd2cXlXH+KOr9E1mSfIGR+xbToxhPcy2RUDdlThySMtXT4lbuMqIeCxoC24
/fFvPO6dmmWb3/PLN/ZuOlm1OCeZu1+/gv0v/TvLus8Qfe2EGzo308Q7bTJ8
5fvuuV1FQDr0xQ775gwVAJrA3QwDqdLWkP2H930/2gij+lo+FkJ9uP4lL0+G
AP+BgpTwhKDCeTXoB85eyNzLM4fRSf9phE2To2SlrJYsNRm1GFuMKW60lF7Y
e15yJMTNmn5Cd/82UHtk0ssvXoxkcPBA1thCk2wIOJ7n8GRH01foCL1Csp68
Az2+ol9bIi32261bYs+NQpJYQjEnSMhheEaffR/XEHkYxKgCUmKE1xY2Mp4q
FgKcbzJ0j+9i5dT1orCM26SWalffsyb4iuvGZvCwHtTu3uc3Zp2vfJ2ZXBie
choFUrV8ZIxySrt+RcOYpRXFofMOrCPsIIao0OKLcW0EwvcMRCWoZBLAkR4z
5YOuGscUmneC18XHx4zj0fRghcKSQZ4PRy3b67q4V5z671SJzteAtMauFNSD
umQRj6nz9oGGM/IfPJGxuZ8Tbyp7orw3kWNm1BGFoWmz7gYK6mtc3+nnhaxc
JolBGq3a3NCXoE9R1wnAcM49P3fRU5/WSgEuEs8t3PzstV+XHkvI1mRWpDmr
UNLK53P9a/2jgZsoD5rcQA2Zxb2VjVqTbLYPcHtcc7cnxcSeIaiiwPSD9D1X
/Kae2V97tzBNePw8bVZ55kIkZZjhvWEExV6LqDdSjbb49wn4obrpB3N+LaTt
z2I3jbWhoe+1k7bo2iKJMlU4gnoZ8AUzXIjSnWixdZSnzVrxl6yl1Rh3OQ83
zRKdoZzjiAGHB6A4WtADHEHzNawf/HOn3nlen3aH+DPnz9Q51mdnrd5d6s9L
j+tIMsF8JwG+4TfyYKHtKXz91Jtf0SVvjWP9afWhLyfNlavu+hq+4g8CAMd5
+/OvT+++NPLBMPlUrL4TBqToBUVNMhYOOGMFRoR0h48XXWxKY3gvf1g7HJMt
PzsAsBsQ1lNITEmxJeU4BRzPzuC8Yo9SdHhuuH5lWKWtzhHBxKDdAxm1KYo0
x3Jkw8XRNHF+FhSMKmaTKqAuPhXY+8uCvcpIKfq9S+vT/lEWVcMlqK3aZDps
Sa94i8yCLHXL+8EU50GExu3gYSokVxe18gcugvEZKTpELs5KQToWS84PhHA2
BePfVZ1E11gg1jyZe/LE1urij1FsymNCpeAJFb9QXidi7pBL9Ni3uUuVAzyX
FYtG6PhXxZqg5nNisysFiZ+GJEjfSNsJ7GyEc1Z1PPKciWyjWoKB2oemyjwP
09JWyPl6d5IF7imcwwvyjGp7KaqfSTQ//zfkPwyARPg0d39kkw5HIiwzif4F
/LnneKsJqBBK7kS4eUeer3aSAeZck91njZIRtHrhnKS4Y7pHm10wfIyVClB5
ueeb3PHhX8JWgGO4yK77lm8roZMizqh1DQAD6A6PS1a++zN3dA9yO9p+Hfe0
60GKlw8tlmJi//7uiusyCChCLXELn9xoewKG0v3ZATKrkl1w4g63A3mDaoYD
4jimPy1jgT16vE0a50Ee8S63TS9Uk8fvg13LFQWNM/elzipEvCLBpXB5/Z/u
LL8VPyJDjLHg6VL1x6swFTOPsZRML2wNghuRvUKvN5yxv6htpW9SeakuFWIk
VaLKIEBUKAhRlQUNnOsby3C2Nq5fVJUC4n9OIhrO3ZO4iI4gb9FLMm1swXom
rGqfvMfm+1lViRqFj1NJWJWE0EwjOmHPemKUV37xywZnKVoPqktSibJLlVqR
tf7gkQLuJJAhL3979TqyBIuKS17+xLdceDwX/jF21VUgxIGuq23vTAftuOa6
teGQiEjrxLiVtU7A1OLayFbFYKaBdwpulhvJuasD4fwCU6jWB/Nz3vTm52Br
PJ8bju7yOZHnm6umzqeeZho8weex+kxhqxSvd0+SWL3BVqNGUjGpUnvQaq1f
5/pA/2IXniGAlqF6IHJnpLs/EjU1h/XVEI9AQdDtmVPw4FZTKB7+bBh6McAv
xHPWFSh0VFQmsM9WAsxsxLtlHW6jPokwaThftKcdBKgXKr2XHBbjF0+5e9J1
ko5x4YjPZ6h6QYuMR9WsWk5bwSp5cEXWu4OPAPosLE8b1GZ4Cq/J+K8pTeVr
Xl7ZL+YNOXdaqY9F2Q6yCc0XZKKepdtOoyxBOZH+BrhQyDY7QNqU2TMikS+r
M0V9a1tMTN0s9yqlfp5l83OR6NIrc9Y+qMVd41dCe6mdOXYxxNhmh3Grm4wH
Q66lnYpJyzJ649ZUxx3bHNbXN7UoGSjKxubJ7eZp17vxCZ3l5/592itwVoZU
RK6/pdnjGNmeb1KXJDo76VwPbMeSeKit7oxUGKjGDV2lVYIS9RRM7g0bduA2
j4IJ38PFuCuC0pEtHGjWMK2XggbIuALoQUxeVt3sDRctFZho5trhcDvlk+Ba
v5GhjU1AH8lYb9tuuQGLx09pT+F45+cRpybMwVOdnWRuIjyDk5FyNZZ7mwYD
txwKHjouRpVYfc3+25hx2/1GQb6zagCK2LTBnzoK8i4cEOHqnp1ggHg2plRb
0cjERGN8B+2v1OTTuDo5ZO+ntBDhk298dDAudihTR7GJLnKkMiogMDELq3vz
6M1T2PhXWbscJD3idK94iW723wGWag0kDVLTFs3bONsTUdRlgunwkxnww8Ek
tedvxDVLt4UihY5aFVJf1BS4RLODB2wfHifssmbKB0uWS6usIr7MX10JVPul
1KQWXVx973fF40dcIMQuGzFx1JEmqknct08oICYvavc2sA+oUHtdFQDVrvAo
olSE2Eri7qGXUFeIT96cZBmd4wMEaAPSCnf1roOyKfh02ZOFJAuw00Gu+UUB
CIaJWjcpexEqb90FZYt6htdftUFgXxjHLRRVFsIGSJfNMzBLYu2bfMOPaf3+
FgwcGVttRfZ0TpGO8RAlNjF76S4EdEHuGygK2No8BM2J46/LM6TAxa6V9FPx
dJ/Xp3rYyL7MXRkvVx31sZi31sYKLTlP2tIpYqaJhoYLd4qAx5/Bg1C9m1Zt
D9g0WE0Cf2tRxlFANPGaIVU1TVVxv4ULtobXvKCdrYt7RMisKnfu7xnaJ1Zm
/HYYE5gTA0dLGoBnGXcLN63nf37Ctb6HExGxmnLL1yOjxEPANw7XuVWlwIRj
NPfLR+g9GBGrCoS05SqhZ4zjA0ZSaL8MExWpjmNz4Mj78wodysrgEvsQ+Kia
98qxBwNuuvKxt+hV4HEFYSrpd9Kjp9eFgetiNMfcHS/o4ZnRUlAzei0pd+LI
zlcMxk9uvBEPoR873gX8/eON6zi1bhdLI2awsKuabjGNGRhFKz8Iu+44gNxO
bb60FZZe75sPcJjnu6CSed0h3bbHRoZULRDu3RhNlFkC57KJ0WZG0c5yx246
/dscskSX15j9ZlXl7pPkkIKH6F3Cc4ja4Tu+SGv5fyKH+zrYT32eVoSRrHcL
i0cM61IHeTZyDZLNjpFYG7CKYxS0EyK2MgAY4Tvb3bDtIfItlbVl+NghlPRQ
La4+pkPE4c6SdUlB+LExVfnVl/AjP7ODhunoVlffXxad3UvlsvkrVwh7uxr6
l6ZUJGD0Mi2XxHfsc0FejA9daFtY+vtk/dHG52H2m4U3H9GeQ/7K+40O3okM
4umcMWDTV19evNPYGQ+0sx6tay5Ue8yYbp8Y4Qq+s1I1fDwGjW+h4jRnCfnh
k5tU+T0Ey8MascGeqnihs+6nBgrCJmA6IqV7WgO4j6HovZXslQGqcj276Ca9
WhP4HAVq7gWx5mi45MuiDYFFllkRy5gAtil0AmxW5+uTiTSJ7zb5rSQ5VkkS
l8441AY2ePVoVlxiEB7MQ3lYcl705EKt+7PejzVD3lDz0M6CvCovUJryXBv4
aTrJIUJYPdyQTojlUFWLP8agASzfwgo9dP9xdsBogDzqAlXKt/2NL0MFUHWk
OWNkN8rZleo9OY5k1/NceahA6D6Wu6nPVl0IsHzxCVIC0gRlUV+0dusHJvAO
RQ8fNN0CvFc23qBd+jyM6E1f9wHu/GPUGlshYT1JXHasKKVeSVw4cjdwdXFr
+hBrMWS5+XVqJ33Guzb8gkc1NdqR4/Am5xdcAY0hShTHS/RsE+ZlcohKcDQ3
fm+zEW0u26M4tqfo9Vc264Qh/1b4DkvXYEbFPMGzCEteWoGA3K2d1ofWNxCR
YSRYTCTU2eqXKyT02Pvkm9J+jVUWzFqjiFubZ1hfXgOrcjwbQ4G5i+wB01rV
BAm2Al+CyoxAjRSCm3bEtHi+OIsJjYo0aRQZm7UmCI4+SckN6nepGCH1oios
ZYxVm4HzJmrpp6Rvj4NbrlgCdZ+rvzGcbyNW8opPDfI8bufVHWoYo7Q0hsJ8
i9euB8NhqdDlRK+HWNCOW0Pm2FTtxD6dJ39Cimj+QLChm7BfsvfvjZC/KL6a
nHOLoYZZ69ZJqxgYuubZY5ZXfep95LwMWXsz6JWiwnFecF6kGS/X0x3m+Lpr
w1enXluTVM8c9OsGFHVA6+fMz8KU0dw3+qWhWtbFbNx7G7oKZLtWOFyIsGiX
Qn0Bw2VLHeDwXb8i46B9gEOW58QHFQfN/sJ95meuuUfr2ms1Z55jRuEQWK/o
ndKMAvk8CfDsCkf5Di11MvP1WAxP+V6LjcbLPkxhQUbyh9nOdM5tGysuy+Pd
UnRaAuQFU9+Uwz3PNAC517aO1rtVZ1kCGrHLTcVaDwfxfErNNozPWQF4omJj
f9MyiZKFKz+Blc1Z//tuR9yZHjuqqYMcwY+LhHDZT5LEIXOpHY6g1Z7IrvEg
O/q02966DsXKItoupW6ZlFNlzNQ0k1VKUqJf9qi9x+keMdcwTnvAv2rf1zAZ
fxLeVoV6PGF56cGMdxz1h+KxAO/TRLoa5v2GeejR9TgJ6r2/yCtZbUU86/Cw
ZUP2pDh5Tm7gPPk7wBeyb4Wjb6rfRFO6MG2DIddniNOOCItCK92wtX2WLdhD
p9z+9E/4MXd44vhAz+ItQvOi7YNagXCE6faJsrpAfRX95bc2TQ99yHKOTjqH
mQTcmSWzbON5RrTx3XoCj59l3JFY79qVc/JKvgCT+0d3dScClyo85EfL4C4J
5x3owRM90gM1K3iDD0MOaD0IQ4E71ZewBc2Qmh74MI3byR+/wZR0XDBHOKGb
nypTU+WQiuy4t7SpCr60Wsfl9XgGg97BWKQbmCkYtduqyT4ST+JBXKFksK1s
HpF8GHuHdQjxiI0JcrfsEP2JWFrvyXtU04VO4sP8OpvFSbs/w8vaRfNDAqZ6
AB1zUcSJ0vh6AsyZykj1wm51vZRt3lVkfs1FuREqGi7sHdCA50CVDnQA5CUt
XfuA84A8VOSLnjfP9LOKW9GJ916KhzU7gyybj0l6ux0rNVAryqJINgeQ27rW
BFeiowXNvABnwdvPD0Nwg7EARgmV24b9CSIVjgDmoF9DNTgpxOKuaJ6Is8xa
Uh1qt5Oj1Y0O/C8fXJJohPtDLfy7u9RkgAUGF/+VI9ECKJDJs0WXP5wXyQe+
XiwcvbmGCQIc94FB0+jHvlwPrFDXOyujyqrKDzfSzrAc8JC8jgA9VZuH5Gu8
WErOHYEA7us3kbTclYI215RWZcb/mRJicHbmyPLzrtRvksUiV+8SOP/b4nEm
FnhyhwWmyywPUR2xhh823cPsLgscwVpuvKRI6vPcsB4zMhOqIi6IL8uKUf0+
/W0FOdoTeGXojWTrX1QMCFPgd0CiXkH8yB5/a/OilJ2ZOGIM/jH+WHIhDhzl
SX759pRWiwMV77hRIhuHiTGTp5us+U5hY3ccmtmiLWpuQfGWd53YITo2a3G1
XfxHSXH+quj8jnJgpNHDReIzamMIdUcMThpWR2vfAlDqFuKNkZO5kVZFIC7t
3VRAmq1+Y9v2g+hw+1EwKXcUGQZU4m6xIzIMFWyNcdEinBhEO9g6wyP3NP3q
ZdFJ6sD2LUmsG+AYYp7VMHYcmESnmHCeTMhCrBs7gFQIvEA2bMtj7frANlZG
6fOv2BreOjXhlZhjaVOMvIQHVPGXdwFMIZZGTb2EL0ZiVt0YZ7NDB/iDyZ1e
+EvtTPWkM+Z7Y6d9DW4U7F2SxDud6tYZIhpERcJtRwKkFahZ3aUfVXl8KCBF
pmHWgFqC+o36792SL2wLOII6ZJr0QeSa7Pq+XjQXOniZVUvpVsGuP/NghT03
7kApV40V5YpFcXto+3n0CuamvAwBYeELRHmeYHF0u7frzqpXMkZnQY093IHv
Ei74EWmX7aUduHs/H1QOF1/9pOCZl5KIUFEtgBxfMn4UbOF/UCPfYBaBlx9w
MT2MGTMnDq9u+OmWf6ilcuXbPFfv9J7SMVY5FImraPcgCH531k+HIuMpqk6b
2vH4mgwTF6BPmkXveP7W2tfbLEuOf0G7clNSXovvglM+nTFQzt1vMO2maDG1
Xmxx4anYUdqY9SqgAbTGFfVsumTEJuvyZtZ/UgXHWOD5sSRlZ4ExJ1NiMDbg
D0vK65pjhD49rmwevfxxND9+JtmSbZhYs71YHX0T5r3EddOntWc6Mt4DZV+J
7rCMZTsHXkjT7oi8sMJfwlBw5dStjYguNuYQt/7T5CfTIq4w88XP9sPdlJxS
o0hGigdkupUgTEar2iKbTe0fuBoDsb5qapGmruhb5WF3k4lFrIdawJHrOigD
g+5j5Q5hebwfH/u8Pm0L4rEOVPH8sCnheK9q6BBoKIie2L01cK1pI7sdV/Ur
DsSKt1aSK6JdG7hBMbBLXnzZbyAXliqDJQKjDpGQzTaMjTuY5hhtit00fWEc
KtyYJ+UD0qBjPj+BGxB3mSUbqUaFbywgFhKyHaHQcox2ySEswftGUVy/pjLh
BL56+wCQmvAAJSoHDhMfbX1VEwlUHJDqfwRsjHObn/PgSEizDleW3+Ft0F8d
ldhtG2gIU2daqKr9+Bb+BszOedwz93H9WTeQBnrzK9b/ubrt041iB0asl77A
Cnoxa3r+Gu9BWp/QKRa7w17C/SvBVxX2+d9CD5S6AP3N0v1XsdTfRViQI/qN
vCY+1YO0utUMSggYhkbxwNZqLbwVpQB48MWSoKHbolopDAwKtojgvRwbyzsf
FwEXvMCTsZdmgtO1bY9fxUR2//VddtN2fPFsW8exg3g1at9HIKiGEhHfywKI
t1fuYJf+z05P+st6KbruE9gzuFWJWtugZgazGiqexkpFBFtJQJsmaY3ust6r
GfqZUF00MXK0UekG9763jxJcQ9BsKtSguNJY8J8gopbz+358KIld97pUx3+n
Fn6fJzRrT7hm9693bJ3UV4tKjN//nVaSn4TrhwFS2PUk7poTXkBH0spFY1+h
6sraXKhWGppxtNjjtQhg0P9/p4UeMc+b5uDpLd1ZD0UjAA8ZHYGMgPUhEEmV
2Sthc+C73Kd/i7sPzfEbUFM6ikjRBXGcoA0bPUX/xDn74HVWPY4LI/ZahJis
hdCJk+HoBdBZ6+I9n+609F0vHcY3cGLKyFu0tY+Vbngf6u3XLRIRKrqUuc3G
/xBMV6XG+0RzaDX0PWFsMiMdlUG/mp/9k5f7SR7hvzd0cInevVi5LQsk2j0o
TN+9oQNgWhB5I/WzAuIj5hjwnlwWH+k+YLsPhLNbfEH4gTvBNnm9x7nzgeBF
dG3uKaM+bxPc4adt+Lk9kjeUHfs+vkXEx2SD/G+N8aEuWtUrgIAb8fFPrkUJ
GUBRYJilOuQWRvaQtyJ2GIOU4K7wCg+oq992DWE/cT21POz7jRlNSLZgN3Td
sgBaH9+d2bnMAIbFQVCGVo9LzXfa9jUHuErJqvsR2PTEadcxCwG1SjD024YW
Puyld6SVYGFZS5rWaQMzOovNRlo8fSwXi4yETok6iDKknUACKkgvP4j+orFb
lI0jKLF1VBYmzM8FHjGxLHlftLlFeyC8PpDkI7ZuLzinhSp9gfcfMbZeudZ/
oq5uAd6StKgMk0zMjEJmdJiRmToJ60WCZbH8nTFcQnC9IPj/6vx/UfP8zXHX
WQWO7K+HgAr1api9hQCt3YtU28ExCvlSHrdSHzp+DvaRdJsX8ahBJb1q9GkA
YYBoRyj/5zJIMnWw6mYl557AApQ3oNpGMQO8gsLwOCeS6SQj9/ZIXsWMkpu/
6+BxFIGOten5KJg9VxTpRm0etOm+LW6gpUOoGi+HZ2OHl9Tb7ZguAZvALMrm
sJ+3fkxWHhn2Kp4oyCsFPsERl6lUdq+C5XvMJcDwBy+SHf2L/FNyr+3Ll7Ng
ac1jBL8oMQDikY5cHOzaLfiDGocu1J7LA2lwfiwfhpZkFnrok1DE9rmC5saP
yk+dzl159MxRF3Z9p3KgHve0fHYTUK6+J4G5v4ke3X8ZvxaPyJiYHGJbbwPh
uY/rkB0fXlNjbomEVLb0lLLs+fLv6XgbAyIu+VmDzY/7s9hmgRRPBTcOtlun
SUH/DVnNhpgDnbtMicnWIdT69AH5eJM6tpzvjA57Zs3goj3o3bNzpajAHNHG
f7KbSjaROCxbsejcobQBQUxVWhdfatq+gzdNDfO0vcubWGQr3SkrAKAkSzVM
Ix5n24CqNEsjiUio9ik7aEPm3xv0PVjCiZ9J6dbRqqUW2swB3BE8VQHoHWSt
MJuOQbd7NPE0JLnmM1q8IFs21s9pucercEEDl9aNYFzKs45NhSKI1df8mnM1
4+xr669FGdH/VTiOe0gPjiPp8IKXniugjW/kJUdI6jU5bQFX4m3Joi7BaeNi
G3Pac3JbyOn0s2KWJnHuhIL6rN25cl4Ag5Lv41gnBUa0LrFKyW7FYIjriQ9s
SFShvg6TpkNyLT2pKA5fDKZ3C1QeA+r6dM8GnsVBm4AdZZGFYb3YYYfX1Nh+
JaAhshxQpK9Dc++lXd5JNNqvaUmhC+txbxNVy/Wixu/wiONRCC+HIJxjK5Zl
zFPzmQp3AnO25Anh050QMa/y3nm5O+AhTmh+kAD/FONBALK49zzJrRsFDrbW
bgT9XjvDY2kMyCTHstzU+lHYmGuPWPdGsaSK3GTIi3PUZDGfAtpSyPx83BgX
bwT3t/dIJFJ5aSo41IWpahsvnURnuccTbYi6dhTxFoUWUaFGw9ETACZ0ygTW
jw2bN+k1eHxSmVtY2MoRF1Qh/cFqlhff0febkvrTQKMHgLXm1en+J5H8aKt4
aArYMtA5Zp+gHrTAkyFgPEgkL25kUxYEHKvn0AjJAJi442oHlBz0N2n842oG
Ez8e76Gu33V+tgA3rJA7Ww1oKzMen7vEt41Jwpimv33EeM40WCPKPFecu3y0
4jpODmdx153i1R3sndtaT6XF2ERTYaeMCOiO9cdKRwzTl6mEtkjiYbNSgHAp
GMesU/4TcFqOFAoOAq1C4AEsU37DB9JwlANfgdGpCNpUq7rosIon9XwyY9QR
je9FUZqpU8gqeYs9/dEs2DlhjygX4ctGh2GRP7fL4WDxR22qBdWvHlvNI8s5
ymFrmgf6qaCypW+mUbBs2AXn/SO36heThiZUaE9biE3HWa06T7a9xb0cRlFb
y65m/JcRSvtJ2Ninel/J/rF2W/P9nQWNd/VBJS0wg+r6a0TAYtzjHXrhY3xm
Lsavo0/hlxkH32bPogadS0PRP7OfNOilA4uvEogFRD3ZXaPKLpk9mxfbEh6k
B5E2ON76Vn6XG6/JOPE0bCrb0zR8f1932KX7jMVt5L9sWzvUiDNRxn0fXl/y
lTPcGE8ffw0cJTbJqLjmuWBOzQ1qQyPEmwr6dwAhrDSlMNfqb727G2aOPtgz
66CbkNsVFKL91KPvhseASlMvBrkLdiEiYIqRtnYvdLpJLQkavBB6Yws9yQMn
fmeiKpVhmrYxFlGdjm/3pXDV9uVRnVNsz2+DZr3eRP39Zri+kLZmxN7wltUf
Eo5HdZPuojiVuaYhRoMCbRNaDc3xdxMhkHnlUwQT92KX0HHrLIfnugdDgALd
9rZ1c6fs6ww50MZ+iQaPcXLaAE3COn7SR3NEz/iCAgQ7Q8/ItndsKvBhXhQF
uVJ6CSdAt8s6U8HIj7QtebCZwv6kM/AKYnCmfDwxncRSRfTw79QpGsmqBade
zNF7CBFB5xsTe7IMcuD+lIYRAb1eCz89TRlsSmqncv4s5yzmLMM+zacmgb8g
PLBdzBoSTqoMp8EsiE07yFbwPfENmw6Z3JTfrKwWwzYFHbF9WugW3gY18pql
mbcVF8yirCNO8FshQS8Qw8gifAdX6IgtwQ1dA6E/PWcC9fgrWXZShxPromtV
K+6aqugCnS8dk9aPPHUBrl+K74UuAL5ph+V5xKPJCuNuAWWbEGtp+DYWN3r5
hBWYyktlvAEV8GVfUBW7s+60V96PK64IK9m9yF9ANzauRqEwKrKgXlZqVmJF
PSLJcfifsxLm+WeGtuyXwHeopSkPRuWn2kyOyQWNQqFOxmixFA3U12zOdsth
7RDSseF2jDargYYYs0/1o+8Pzpa8+NSPFLXRcqMSWf0FZZ08ohI8X8WRwACj
GTs4y8nJ5EbMpaXUhsqyHcZxG4u6QmFsz++kkBqu47S7vwJnnhGXxdABgQ0l
3/XXgAWFpdqrpYuYoYmnGAed7Y9pcvBKgJRrRNKK/ZA0+BIZII253KfymPjp
FDkEFv2mqpO/u5WMbWnJv3vgdCtC4W0q2I6mCwMzVOjoXerP2jfuyi7Q4DaF
PK9mfXgTtxzaimX6aTPXqZd+nPApUEb4579Y8ifETKls52KbBnbAIQTBrVhn
P8vmy90c5/ZEaf1zjEg0p8XHZc6md+qv9IUin28vBJ8sEyzWDsIO/8eKnIEM
k1UN8EBd+4k69b3UmTF4jb1BMiQpaVCeRazOQ8BKDbZtAQ+mncmpzBQw3pvV
YE/ur9PxASXQePQIiQLnpkshewktly8w4lpbelbh2AVJ0ifs655L8LEru53s
Qc1DFWbzz4mZx3QQD11EY4G0REbnBeP9JUQ53iOQUVkDwjLepI62nYOHwpiN
mOkSziN3XiBj/aZWnMRcbNNUf8Zojg7xp1Bb8IzolfuDS8TLZWFj91cGu3+q
i/WUWAhbAeKgNASUcrYmQt7Xxor4T8Yh82lUJPU6VkVzWsFabZKq66+89S7X
gJ7hsA1C8WCssi8itMc+QyPJ6ecxIwymim8KvkY/1LG2Ynfsc0H0/7VINZzD
sAnBI0928VoB0Pq/zX4VF+Aw+iF6afiSFBFyL5F1sFAVUQpvrPepwVOhG5fn
YpX2qAxpQPzwjoEZ/bHwXMF9WxKTJFSG0MHKh1MIAZdm41lBBm59g6L9u0tP
13HZAriHndFhPV1kxPvGXZgIWmerSAe04In5/SaTw3deWJSL7QFhV8gulPjp
k9WHJaFdbuDww5uw4LjUAB6GeX3r+uctcmNGGlL/frW1SUfxalvSuF414eN7
8OkmJByGYgVkWxibFbgvP1Zj2HSdcOWMWYQZ6vW2Fd7tr/0epjStoPGAYwck
0xbie7tPF7p+09Xr0R/EMfQE9Cu4OQKMOtf+kRLWVQHhQ5ZBebI3VEclKVus
8IfT9Qk2gaFC1+HLeBY4WuGBGxLssImiBdeLVqwrfA3Yo8/rop97YzMZ+VIA
pfEV8dy/BuHl8IyfTb5ilnidd31/2piNUCgZFz2UYOMh5mPt4TT9APduXZtN
Mx3DDsTXUJNJ4o7b5j6QoEVNuUOsgRbLb6PjbcZSCQ8eug+jVLSwi/xv7Zms
UL9eWDYMJO21ISbIzGSPUsUtJnKw4ZYPI3SCcZ6qISM3f7Q+V8MiUoCEp5/U
BWvwsPRcTt2uOMczXDEMuvBd5KROzX/EI7vSyGX+OgkQttGjHhHi8xNAu1E/
wPwwzpDdpFgFut3irh/jmMLzyRvMt7rUb7LUCod92hdrernCwJtY81t40lTf
pqpLCEuju5WZOvNXknYmhpMqbwxXLE7+iBnCvOXXg4F0kXU7yjWMEhP4W7Y1
5fk6Xh4Ngkh3KqE47EZ99MizbVmVnoZclHSoWE70ltcG0TgHvAFHUak5dSbI
SsoJGh2Bze74lWAoKOMM4A29vBAhx8HD/clAvqca6NQVNknBrNgqZRLGzRuh
6BI6xbixkLSenB3ah7W2gYagWK7UWZIecx5L6rdPubOIowUR0a//aPY/nQJk
JxW55QXzunwxAI+WIOLmNa6TRM4KJ4GQX2CvAd4HG/c8TlRrlSGowIlreaLR
u7tH86WzZY4Mmh+VbJ3Qd/SHg/xMNTIeEJd6Y+XbKaONXgfgbDJUtBXQyWU2
GZLi4KvZgS1dFDW1uLFGyZu3pR/hM7QRmswYsHTkWULfUqR9GKHMn5yka4Tq
TuYnspSvFPiwYd4w9xDS6susT0B58URVREmiFya4t242Wdyz7tj4w9sYedVC
KMn+UG71i+n2k4qEr5l7PO12NLItvRpaXOEHKgV04OtiGIKTL4rtCegPSMe3
iPpjHlWBwdAHa+8ap+YbpG4pUC1MJ6BEO/6jqZoVzW5KSqcoWkGh2ccS8Hrt
Yy07mrsbhmwt1GyJ9SjAsAQ+rOILTk4DlVKHjX80zYYQg5kGwN/NNZBC/VZG
vDuCOGWTy+giTeWI/QjQQxeeCDpdsYVVgZLdHMdRxUF9AVMY1QagBS3g4X7g
QIqaGEj8wi/4bdB2WT3U7wP5HH24mFWKeVnfTgxzuAelPO3s/uVyT1L/I4UO
TzJDbbAwxkGXD5OIz135jiTujMsdOHU/ANQHUrcaZnTy/ERLM2viwS621ksF
pD3IennphNxOPfCczmUnAjCbHz1s1zjrDPWTCP0MKjvtJguyXLkKtrBNxZyP
0HBwo4SSyxuc8kT4Ur+s6S3YdTWkpss4x0Ca31DUzqVgjnChtx+K33sP6Yiy
UGq99OmB9x5i7H5EhjLWave167x4OnHgI2PdNPZ3LutCoQBEY/XLN/ToQUmN
T99C204E+KWo9Hu6vQsJx8Mm3JOWv8QAJba2LvD8lJ12Gl3m/C/CAO5BrKVZ
7UnYwnaB4+/kZyRj7YIFnU1cZrnUYtvvTIROsHHn3wmbq/Aq902YEUBIJAwE
NuUM5Itp5wq74LX6ddBpb8YHBM19jIz/AGTwvK+12GmZ6T7sPw7StS+4upon
Nt12o615C2EPfJkbzZUvUYh/qZPUtQ1pnHac7binqdd6GX654MrFE0+VS3u5
u/CcsqE+OXT8P77XPcgKGbz8WMGk2zD0b0pVhh5F2eLd+xgodqhCtm74XG52
586iOJEGqoQoWB4tJnX6CaHAhi6+jd85N4avE64HFDove1S7wuukV9kb9jUw
FEHoy7orE3FW06Ee5Ld9SAaXMAxi60BQ03OlERYUBKyXz5+Qg7BwPcLtLlfj
OEu8wOXbweDXbnhs1Ow1m2ADCPovJHKBx8pJAlfGoMI9UobFFwRkCCK3CnpJ
mM5V+un1uTBO2bKSzq60Flx0BKMumPvnTyikbYOjqepTzpROPO/AlNrwcCeK
jHZtK55mLE2+LheEJjbGcCsfhqkLzivaBn9/lsxBkm8uJiKddNYtis2c9oKj
yKOraOAEuJO9yz4SxfLPxNMNNFNly7Fj5pyfyKiQm5KphCIJvRUY1ud+jitA
eLaMug56YV69sY9f7cGfXvrBe4zwc1tnkMY3/ExOuO9qrFF/2J3Vms1axrg7
TkgyQ4Fv/FLjW3EIq6z5sitmQZ683ljy+eJ5wwYN3ZHekegD4ipZeYhCwSuR
sLPhjApyF6ErOc2umklbuK3ek6wTPePU6NUuk9sxWgCPioqKLACFQSTKt3ER
ThlHnERdDti3SrDl9NRcvGwmDBSiD/1C9Ooj+Aa3BHv9KIIlxwNrvv2icZKB
4aU9hd90hiT/ZBHxYuTUkNVEvYyvTao1fSTCrE7D83i9VNkixpQVLzDRbjRm
Wwhy0Y2InF+bw4iVQVTmQTEzkWSPI62KfPGkqUZHGFZFGociRFQygWYmG3If
FmYwhCiKXJ63EzCeN1BCmGvlwtLA2Vf+MR3DgSrUIyaOEK8FboTvB5xIQilb
vmnvvsSHUS7l4oH3QSKD4x8NjKePo3eynZp7c4ybij8Z3Z4bzLPbEOkj8swm
WOJ/g0uJ/pqOo5NiCU4Z4iEm1xgZjHDEZhamuGhiES+dGy9Nx+bQMIIRqjzz
dyeBupkTVZkaG21R9k5nT2BkOzw6fZRBHB2br/uv80fRUvtY1xBepLjwrD3R
e2YmxaIy1XESoNIsLSB13FiyvCKV6axoB2llL+pYEmbKlv2Mc4s3OciHsj1z
m2wv8UiMnItJD6uGFeHJR2eMHNwB3V0k053aaYB7i9cOPplrEh9qDg87GP5k
BCJqyJHicXuq9n3zqDHp9lHJTh5vFA6UYiroMu/nwQAhp7tLhvwSQVhBjStN
tUKDSonC3zLvp+WLxkK2xLISvBosPltTn57hVpVHJKzZKb3AhHbMviZnf3It
1hoJzhNKseXuv45nyehvWPnPDNzJIRHutFZ9+LwxSoybA78hF+3dfP0fX7Hy
YK1fCpAokSwOukEjM8Fa/7ss+t9sHKCbZxY00j67ttqnUJUp2GNVLEhv8ZCm
PvibXcDY3mx1lfpcuyP7Rjv8pGZfzU7lctl8qDy4LNGHVPdXn4gzZRqSw4Mm
/pm2dTzqzV2Cz8CNxFObMD2/EdLpOXbIhIWrsC/VsvZxjDbCmQ0bNgPldHWC
m1J6tx+U0HAhmmRoej1AUY+A3aaqBgMbaaX74SMgbgOFmFaofXxmGNWK37pB
KxPpyR9Ym7n5WvMnR9dNydUCbrD/RO06PmhzMAWIzt+hqTZfy0gGJHWrflm5
o27ZnJg4FFcDT8zJq6zWPZaUXfPg8sbzcB5ltgz+F68/c8rN+KFsHeUwugvA
oOtjn0R3+CpqBQ4OHsRI2rfv5pvybGynwCixGH4v52XkbE9IXckw7KYZx+nh
XhYhHNhHC/wCj7sBOaMXa8DzIAbUnR1was7lfaN6s7ni+gqbXQTDTJ+e0aqP
jCda9nMOSgZoSvnBPNbrzY4imSQdU1XibvLfoyiuCIFqcjoydypVdvVJ+fD0
K5GDviKzClQPVWTTcYOJG0aQeGUF0RUxtJhmjb6UNbkf0C9IgQ+GDt54hNfm
sEaWygOPRiHm5ZRN+3h4cKLQ3fVsQdt+h6z5FxHoakiChHLVg/IVyPoGS5py
iXF3O6ZGUKQkFGdituCBTAM0eQsM/qEom4wcmjOd/ymn2jVOETg9KAPvE7cm
a8s+2y99Xrvp4efj2W419rvRe/c3bNx9Ht5xsFA2rzp9XXTLb6V2P93BMVq1
I0SzhQwLQPAXRjuQ7kElOFASOdkRIJy3NaFIzsPtjUQNMq1upZtU7uXNG7NH
ZDf5TIEnJrVOjAzYBmFQRPWOTldWvtY1l5Ybfzog1dNIoYduH7Zm6dcxbYZ8
bf0KLiyINVkpto+T1s//HqpK3hcWoLyGQv4drr1DeOR7Z1FDQSV1aMz9SPDQ
fXEDvUyZgQybrOBxvPE+QQvaBF3trXxEsoXO7BgvzaWsT4gyY9iCWqwoOPBR
GKotIcHa+lj8H8bN/PuuxyiHB6Y2F1Kqyt44xaeiZ2/QEAPn/wVoMvUzAQht
G7ebRfPLi/E5suwKNUXxPKZ9gEjvvvxTjfwFzsKDnvojYvca+MLJDcwaeRJ0
wM19E/F8qTtaa8WvSGfaWjW5tE7x+7+vJeBcCk06RXKa8pJESl0yBJ0eCv2c
sLW6pNjrSo5I8vD2Pu4VHHXrLvmrvom66L3CyM4nF1yNKHjDUTrLPU5TyeL1
GT1nmuUigg1qwHzLVYpC4wSuxL4IwBuogwS3fSeJF4RLPG4ldjf8X+eXIBIq
Fjkgsf56UX7cZJolpRQ8ue/mG4KxTEiCmctr9briQeqPxkDkGgi7McGvo/gX
+M5osTYxXNrWvuUn/uJ4/10vEAMyY4LMeBiheh2kqxCGDupMUeyjdUeFuKk8
4zCs7DWBbC3vn5vh+gY6yjLeYqP4U5OnQLnREG+uX3vK7Ezw6Ocrkt+8zZFg
HWxpsuwYk9+8CXbSOYSULzx6aVhmgKfA7yCXC9VdwbqT+X37nWnITEhySyZd
qRXmk83IeM6mZpCdZ4GzRtg3jEYXvmiDwO+wffNPYlXm7gSlwlc53YJ6h2tb
p8sXtFBimL3KGkb/lCSo4wBQhGWnCPTyCoTW8TtOyHQYbq8KxzIf6riytlzS
oAcY7KolwlxVaDV3unYpU5dcY6BF8TZH1jR3cSH8r5+vj4cBL41zJ3MPhunb
6CMDSNOFjzWiFtGyBXCjBnggbatZoX+lVhRGxEiDU1G3lPs8pRzHOUAtLIph
mj85XZSgijJOFX2qYQ7t0XBPG82B6sDSSgpNlXSzC3Rg/fKlmtj8wJbmWu4G
16cO7lsu4XMjmGCRLAAY6Yj8sVk0oJjrcoEPHFO1S7f3Lj8f8+7sNiRie2KC
Vd2H2g9cp4mji6gwMDQkPGWqUbxGhM61alEzkakDBe3uYRmQcwH8PaI1l0QV
QnAFllixBu5DIvePmlAY5UCv333InCWpYoD9YkTko820Qi2DxnTHdzd8MWMD
AHbYn4MIEs8DMTGz2JXtQjSy7J52S6nrctWzyvh9sV3xTMRf+nWOjzTpKdkZ
zpej52zAy7XuzyYvXnZRoCxIzPHFl2BF+4qGKYwKAm2Gy6F99BLNV5sb8U5W
x6PhHDUAW71PIEF88ZvgQUt7zrOr97KaazaHO04FUwCsEUbXNgTzsoS9OdOG
GLwm0IBm0XDZ2CHHjm7c22RaMAqqq2KGaP1jCIED30riDzCqRnGi8Kqspxrx
ZEBRM8kZZBW+YEkjE746QSThVTthQYjvNtrolWUP9/WKXnCfjZ8zRreab/bn
1yT5PzTTNZZV2NZKrEnALdsyJckqFhujTkEjZRIUCGL3tRSLMcJw1JEwD6/W
izv/uCmXTzMUdcUNWc7my2HhLO+gdisXuXTWDxy09l9dkyyU6ZP6TuRAkkLu
Vo9+FvZn+c5sYJLVSKTlvlVdsqebWf5OuShip9XYK+KQASeNLO1JCMygIBpD
+awLCzEsNGGq6HpohGOTKN+dyOclWRbEr5+khj5zoRXg8B59x5qvr6NXyJ1h
zZ+i6HSujSrl7sWwlfFyiCQloaRKM+ujqSZ3035UJx54H0gSPC7Jvt1WNGnM
dr9Yq1UbxNfxtBpxgWek0+fB+db1ttRs0d2UBN19TkoGE+05CsCUgCXt3/TE
py+midGGVQ3udOTrQCV/CmKWh6u7uL8XqfWz6OMsszqQ7/MTgz5k1HN/bf6V
mDK1tHFu09VqIMoO1J6U5gZWwAWYwRR0RwW3j1vEHtEKwly8Q8D3MdxcBobD
SP5C938JlZyP/CK9SUBXhZGmYD+13RKJtNwP58TlSVcA6Kj7FRBZ4xzMHtup
1bV8eyquX1Uwqm7X84hsRG3wOQj/xvuI7fn66m3rRJit7ESIKHgGwz72S8/E
yS4w9zONL7SSuXapGudkX4N0OgY5QzBwe2EaLVVFP/YT6xFpf/hBlPfYQoXU
obRn+gfn0S8e3B780cuEh1OvO+wLCtEPEYDhrmt2QQboqm4wNZgMQrHqmaW5
+u+YEFAVG48Y/NfMY3NK3M2tsBFQ6rPw25M9FjRVzguE9PwvK/JQGupayY+3
G/ToP4BGvLDS9A/BNPbjtuVC1Ui1+Jyg9otyKLRFPs1qKrkXbUmSm2ZHXVRe
7qYgLW71rGOqkCZIlusQUg9/9iQ8O03CCpahSioeweep9T0bxp6WYREHVHdK
DxcmRr9fePLMW26tRTxEvhkgEfytIl5o/HK+5XfMsiUDipqgEloX09syuvBq
FmyJZJ6yyB/FoAwNb4MElRWwAojsB/NkVzC1+szPnHSjZuWyWY+AeDzGvgVG
j2ieJ0jaW8C0vycTKuhNp7Y8qVgaMaQ0FTkzDBiqslLMP2qawCEJb72y24Os
g383BLNtabBum3VuBIs8INWWPw1/VQF7ok1hKsIbNbCt2M+nJ84du/BNtp8d
kVs7oHRYEvedn/uFPriVoUMhipJi42J5CQ21pq8AhZkAAivpWhZhhyyWf2Ea
lZdgzBgHiDMwVdikZoEd8MpovshIh1R1nU2QQroylJGEvH76cK7aNohiySQK
bv+Maae+iVULGhKwHiF8zWK1SCpSvAb+bCrErFqrsHEu5/ByMZghlqHh8F1x
0bn9m9L7Iuhj44s8efdtscRSfpiDG51chfRc59TUa2Q4Tv7lfCAGKnzayDZ+
xqQ2J/7uRceeG0NVgxJPNTtG6yhm8HmETjceMco7x1r6wUHpjapwLrXeBRSA
GmAtrTDC9cUhDKZ0VjMAQ8m2FnR02cMScFfGeovLKCAiHZk0UlFwqyRkRjP7
IvNy999eBYCBBLuvtJCqbTDx5MVrMKnxI928OVTS9M2h/6HjHDRImUqE6RXp
/7oD3PQ0Z5eWtunf2kjFSwUiGjukxZaVgyKhkJbYOgSsAYw1lGAru7qKvFug
iZ9D6ARLLxi/+jHEh/fQkc+4FDtfTeTENeQKHhYC4Sv2Bcpuoji0eT9uJXAG
PBuaO29MH0YSiGeGCi76sDOC7srhyKo5LaRk+FIpxYSvScUUXRnrTKwsIP28
Gf2Eioxqov6EeE8qDm0XH8rzZTFqqy6zzL7Qoq5pUw8K1Cy7TCvpVeYS8OHo
EWsre0VD6dVKVeSnwlwTy1XFtITlnBAWpGKWUq0NFWg0ggQpLvBW1KEA+2Vg
giNnU9qGROAlwkNw0HrtSy0m72c1GcYesPjkNX+N1YJPpDAmXnMIqc3Qh2lY
gSytInQr8YV/RRqkOx35ntACoyqEN1WjVcKC/olQlh0olx6685lQkZO7z9VD
jvVD/isHWovJ3RaQWUdYJS699SEiUXyaLPxVk6IrCIrE+c2+pLU759ZZuVpC
B+2H++B1mGKEzHZrYALSR6EQYO/BB6u4ljjRI2kPmkR0P6X129YU6J6rPPi8
lk2QeTRXqJV3045OVMhqUs21MU0A4t164rnS4Yt6PMgs9bU5FRS3S06cxFfa
KkKMCQLKeevRAN7RFcM2+xANnGtg41aiIJs2M91QdNYo1Ou2GaBV0RYDUx1m
buTnUfwJErAtA635RyHRaWOCxV6TLe4FEtq5VwD9h5QYOrG9INTQI/YV6TVt
5VrZpNdOwJq1ansUjCxJ7vYoDMDM8r+Q79u3W7IFJGjLDpWXFO0YdlWEGRv7
FR7uc8N0kLmTLHWgpIcmLUwrgYSX6PghVqVzwG5t/xD0pc2mlPcLDN43yH0T
8BS+RgdDm0SgrWO7c0hDcNMb4nOqieIqhCrh5Vwf1/rI3O4fSv7HOUpnQLb0
/wO9KGHGlJ9a5XyFgam/ONWAy9xHwCl82ei182lLOHxpbR14h2c3K2DQIDDe
XsZzQKmwZ5/2E3MD51uf4AgfAPFuK4n6rSyOQRrsTZRTCQRqlHdWqT28M2D6
CtwCWz9QYnFUdPjTfRzwNR88paxK0ItGwJjCNJUC9csFElMm5PTWptGfPRF9
OhNjOY1INH810Jxc9ZMdo3q7AnhdaEbM6w5KN7ryrVXAmFgkWFBVQBirDzrf
/vczelA/AgBlNy1DrWIhGR2y6RciObiljBrTyP1X7CGH6Ts2fJbyAYDK0sk3
xPVrWWxLNfTnvqbO9uJUz6yiFDTCXVLGN3NAjmQAUHXUOigOaxqlPHWvohB/
y01gs6GQi8BX6lHp4ouXErLE+SmWMN+W9qrhWnCovzoEKZABdc5aw4dEokjC
LXA05ADupGpxdswmTCkp5ANiVY6se2ac++TrFR92fy7oze8JRobvMVG5r6w6
avWb3eosIxEi2GFmIpQt5wlrbjAMT6dmI0uXqoXvmtDHH5AqDbYGbBV5j3nV
IFAg6cT16dCcwYXsu3QthBcnsA33wZhPLKg0W/JSEXwo8nD3FPxncSaI9oAg
nuFt4iRleFECXVk53X9Rc9K3OrWm8bNeYAg6GG91yCdNSHzp12VeYcqO9zLs
RnK3o0Z3U6R8D8VyS0fChF+oDKZ63JArgt8bED0TUtJeOV3kZBgtirZgmHtY
7VARE0Im44qD0yt3hBnY499DbVVZBKWkHFU2fuIJauQXudJV9JzMYyB4Zg+Q
W4GSKQVvU1LD9LWM7TY4FNg6hbDHqD2W60ZNUbQhqNxXZJzhtbKAmI1fUCqr
GrnSL9DZNRfkBfzraSEbfZQCNRjq5ZHZIm32FDks/qWLpL6KDGhIW1YgfiYG
HWe/86HMAPBcB/POmAovXfdxk9LJXwcmFK3ZT2vtJ7nLLrBPJm7Ur1Nl/AcL
esK4DlWNe5ItYo+PEZ8lpU+Ntkr5JPwfPhzyxxB81f3Q5xjvjU5vYSn7K0zu
8iiRxS4wiLY159B+eWKVhzn7DuWHw83APFn6E7XTvYkP+J2UK/qWt4r6BA+y
UhsAfOlS7xWEzUrLLTTtboROSC/Bu1v4rJGXCogyka59KT+c+NjTnWlPAGio
F2fgU1pXEPNbdfawyfe8iP84vvMV+/53E8PJm+SuFGxdMf2gJJbouIgUUS0g
RBIsqUJrXf0qOnBfSkO0MXnGLucWSiT0ispfQy0SOJZXzHyG/5DaMYrneqtX
shM9WaZQUkrbfu1vqKMsZ0V5xYoCZjv2JJJH+RwA4xnUZzqRJp9a2UWIi7sG
4qSF4vKCSTKdxTmxWyvCFPV30Mfeplztz2MD4JB+XyfblsQzjBe59kwRmp4p
C5mekx2veoyb2dCoQgGW2o4A79zmvrrevy63ngNIJiy/8HOzdes8wV4tUc0l
jDjMjAqV/nJ7Qa9+jO+2a8c/nwaeBkOdQticWO5k3rpbI9aZv+GSIsio/3XM
jhE7j81Z7ieCNL3oHHHD+kRm4giD/0x/3hZYnf0iEv46U656xv5zGFiJgpX7
Gw/qgaTZUv0h+L2Qvo/ofPupfpgv7u/rze7JPCCgA4PXz++DgQE8Kvdk2GWF
ty4uakuZvaKF2ZUs5xyX7WD4a+05+J3kFiEvv6r9Ru6aHfTPIRKwOG2zJMPi
SevJA3xXHsd8DkSUOW9DQJTYX9r6pxOXkvEBxCchvIfbQMFecmPf6L1TFz0y
gAqYkMt8iVPfd2tJOXSNThJEGzBoty533KTygG5mhk+Ln1Q3rLYsFzl1cJ95
mQBi+VWzMsg4KUGt1DeEdqBrmWNpvqH4+bLPYOyYZ15ngoLjv6qu5gIVO/TX
kSgQdC0VuSn1e6ljAvVNklq5uTfJc3qV4wDOzGaHAhDlmJ2mU6Be3IcCfcrz
Md/R7+QZ9958VCe2ZbYAFu1DLXOfsOyzHxjWxsifwG69gFuLOPQpdVpe+qR9
Z/9e/73yXfLqFrkqEUHFmEMpU7aeR5hEDux9zZGeFGfS7ScCaN7KBXOmPTXc
kS29e666sJt9pRLkkQrXaJ44a2HaEu9Ig9ka1gCRxZKUvj/oDFkKqFFNBj1e
OUf+nqQoAo0j7UFRdgXXZSj1J0oS6la2g4Ndvcj3OQ0bkM1Dmjp7f1xbEtja
WQOqhG/dV9gs45O4s9bIV8cSmUd4K0BXJr5ytJIzKbgpq/BXz340Jl1sEeDf
JUTUh3VJJsRVvDs7mOdLUIWgffliVuhGGRGMoTok6acPWJNYCj/aCbAD6XNN
yD5bQ0r69TRQUTVWmihcFgbIVZq6HeQphFWx/Caubf9xgeHeu1sVP1WlfnlJ
7KCgtBxM5sK+vj2xyRA9TtHWjpr83A8cAV88EpBW1OKMPi6hzYqy2Q1FR4it
phtfbl3WAeipxXEb7MH4p7BhLrZUYhMHeW0DbIMOsgPxa5IkEMnJKbTjPSxR
ZppEaH87dvfCwnjCnRRBmikYbciFe/uBqxHbWupS8zjdp9hsVyndxhziJWjn
GDxrbkB51+/YngEP8UuIRSzxBj2cpjWgGHp5w07g1NRCUM3yZuKsMaVEkbUb
kfM6EQy20Gk8bNCJcjKnsxEvEtHHH/vApZ6u7JuZxnUXsR9W8EE5DLG3aLTr
CDvFDLHLYBHy75Ugy0xWQkyrZboY+SOSwSlA8eMgWeEB4jZAAE82PXUA69lI
0Hj28z+k05znmq6l+JDFCs0bB4Xz9neVxI6ikK+m6hu0OIKHAbEZjZeIm3zq
wbZFCwMQd+qY2qVSbY5/KRxo+Zun8vWjRX3pBXB7TZFhW7ttLNTDaVFpUuMM
nZgDsZMoTgzOOO/cfwnGE+mlFVIs7PCFIExRqLYByggXzVpvRjnQmElG0GOf
7GyLe1WhHgQ0gK9pzMmEkqMgHXkqCspKLu34SKYTe2fpom1TjRamU66rgMG5
OuG3YO6SWTMEpa52qNF4Mox1PmaqVPjIV0Ng/qTjPcvuc8oRqupsOi17caMD
/zkSkdNh6xWpJem6FD/krM55QBXjpparq4hwkG+1PJYNJK/fh4z5bWfyIQw0
Sp/HzarVesJFPRzPBXuXoQSVmp7C1Zzt9Kaa7gRrZVV27P1VcCHzDeadwZf0
xbEREdO7TkzEgQXArhk/1BXBEg+wq9q1Xz28FbCppNXJMmdbNyDAoIOVgIL/
q9wuveOr9pMqgGw4I8YBWr2Qo4uIbSt7V/zrdEv6dbGH/WbRh9piMPPJ53/R
4pk2ld7HfP0qI+WiM1x/hTn5nu3tj93DGO1LDgM7hLQZz3v/KqISg2dT1mZB
4dfJIuS3RpC+blpjiuHclhE7psOLfI/QOSJ0MMu7f9vmau4d3e7/SdsdgPWb
BgNsrmFQK/a7TKFSLA1HNWCxBAgQaUL5ryIWD7Cie240VfxsHsOZRYVAS4g4
esQmvYmQtPT7mkGgYuR7kFSompBl9O5GaqQd1oLqSI6XJBiDrfS6HrMykV5J
B71sHTiJowkojuOqz++yAbf6isfGLlUcQ7Q08jjdWRe/fVXeldU+kDMAyPQF
75hNjvXm/4ycCfS1iIouZ/7o4J3F+HtzFvfZHVqZ5xJjYKKuGBJ1uOFcu8XT
r0sNL+kMcSc9Lkg/ifFjLpTD2TtcCbVyRzT6g2MBK50ot+lxJYZxHh+A/EKI
sR8WXkrE2vRpa0Vcf90JEwqtU50I507q6tl6xmXjwfYGdi0tEnpDeXJynTiS
24LiJ4i0R2spHuyMhxnMag6xUcB9tjGpDzfEHocnx/wKFBbiab89mWXaV6Bb
k/er+jteUTESuIeL3ZskRADZ0oQN9sazh6MltOmHq4MJVmdvRtEXxXMACsRW
LIu1jOK/Cgu/r4F1AdRnWxEe78XlE2JbYtb/hcJ76qORXmjmxyDuMGeCimx/
abplVDUVCf3WmaiitKtyTSDTc2CvvBgsPFjDASXluyx85ddaMNlWryNde4HK
y8F4YSWJNDf8x4KJ4NQcFAr9KR7eGBfIeCGQrq+HbFJA5zJiqJDPREIj0krv
xVDVW7K0kX6astLeNazGgkZFmwtofUxi2yneyjvZp94ImoAJckxZvp3SZNx4
f2+JngzQGgoVjCoeu9JimgFSC/rNp2pqBsi8JLERTHeC722hkdIK+EjkWnlM
NOMejbD1JQZB+xoyxgjshEJeSIocOo7/IT/el7Vokekya/DwQtyQrxWPfKV2
4BeEA7q4fHYu/2fzuPFw5ayYTyb8swKvWIhNMx+TA0VyNIqEXzxYspvZNJOP
Fr6fBmiVb66juq/UF3O8/EG1ylMaSkQ/Zon+RLkVjZxpkM0c4H+5Jgo1gBE9
U/pY8u8J40uVu14UpsEJqOXdip7Fp/K6QxGW8FjOpXJQ1c9HTsjOMiA3FWaB
AFPqQrYaiVzOKmLc0WXA089d0AK73hSWUqYhAh63Bls6TUuLbpnVFnOFER66
kZV+QZqBsRixttEZseRBAZbwIG/JU1s7Lf/CkJ8czjRW/7PROObDLsKvARlJ
XaiLVy1oN7sD98a5ubSiwKCYuVUGwpNlPT8soM5VNK+QGqQc5pPO2Dg+OZQa
EMPWNz1GRPjR2WYczBEBI84ZMWYn8IKUvjkrKQQh7W9LdtC+0/3KJM9q+Vag
Dgk/PQQeXFjr5RIKhyi/Tr3rbV2e3d3Dzc0Md2MM9QhBHMnN0bj+fIqJHN/X
sPq/hP89kQKxTSgAY48VJWRd4UItz5kMfQkdhQnMhRPUrejabwW7/vvjZ8Kz
y6ZEPysuyHvIs0B5YH4a0da5cCA4yKoZV+Nl5GsvYrehSKAN4G0PjJtiu9Ld
PNIGeLa7elpnTXZ7pqGk89t8l6CokBwlW/2DNRlqKuNJdUdG9D1e6lkky5kt
7XowRzlNPAQG062z/E0hYZSSbAtPM2iPU5mhx8e206vd/SPyFbZ2Ayehn5Hr
cC0I0M3gqRxyL6KvXcz5Dfzd45J5/fqeEackOiLrFu2BgKUQX0DaivrdDyWq
Vj99v9kZYg+vmoztJfecZf9XPwvwXiYeRg9Ltht3WlfHeIYRXKTsGRWGU4wy
VDo6wa13nWrTqGe/wy0ggnj+AxEaLvNah6McK+QlfDEn66B8qXav9E4Z5TxL
7sNSSVZMXag+UjEdN6QqCs6Ok75gLUl3wS87dnwPTxjtV4QHaTMSSZFvaCiD
SFiCq/tpKLMLtalwV9NE4j5CPkppYNCloRbJgl6PrKH0GcuAPwDsy5DYKpcy
Nn4GJA7fFrMiSiT4FYknpTSKh0qXPncJvTGh+pxzd9saaZufCGyrYE4P/Ukx
36eRhGHahVwOubf8Beh3kk81n9YRIaSHcRU/sHC75sPeWw9K91FEvZN4bzRW
P5NfKxgbagd/ff3NMz+whmU0BidVbnSuljKgBisRcqALHy/GFsXvLeqi/zzx
yVB9zZMHh4cPZwacOGFCszP6sBVzg2uhR7bfNxWoHOLHlmCR0agbNYs1BC5f
FyPYXzYnqTiUBXlGUmYn2dXUr14WwzdXZ3zY6cjsmU+dEqhyXNLLtZQsg0Bc
XC+Q5nThTzmBoPD4ZrT2i8LEEHqQD5/rf4+o6IwTNR6hvG1Infg/NhNfE3iv
VXwNc5MSGkSQB899LcT8zMpOtJk0mzp9jIz/tlZgh9LOUzMOHMhy2F9+Copx
C6T5dCptl0l0sa+H+aRiMP8IzcFRfxHauLwcgbLMt2L0TmaOAnfVvp3usPTA
W6hE1f8V3T19mO70BYwvPIBLjITYBSdSlA5JMLYd8Y73c3/9gcwFr8YAkgTY
Wt1TYFPptaOdBTEcf25XeGeWkIQ/lQUJf69Sb4SYGgs2F6ZEbHHk+7L4CWs4
SM6Ap14O9dt/p5dpKYJTTv8XD+1uFCJnzqVHXdyIokVVhxWS3L79x7zQECKl
Jon4qON9rtCgwT8JTaIC4lCCAeKQQXM6A/YqqlKHneE06yXsVT4ChxNf4DCx
Z6EZ1ooIkmE1ht55mNev2Su/3o12rXjdTBIpDB7VcotSmDWJHkNVb07/0CIz
Da4BNZIF2C+1l4gHfNOR1540BMQSf59cDdoyv5cx6djuyu2xw17kM7a/00si
9cKk10bjfIZac5gR0DEZEnXmoVrDgtr4HsmO5jPVFKPgyknjt0Tq+Fe52Qhr
r6ww7hpEOmuwah5tQUO0/55boMzq2GBIZHZB59/z+a6vQZ5WbMiVJJik+Mls
s+yFZiXlZC5+WwTcW3698H/0n5dwkVRRjLtfi6ks+uDJ1PtdRIKpPgGBBNJq
yJOUDpFPwrkU+i//JPN+sRkEm9dX4Py6y7fS3S834rE/5/+ge2T5q7JozuAf
Hy9eHcKFi1UlTW/X2I+0QZZpPZwuxClirvCFIITnHysr6efvict07tD10Ld2
WEjc9M7p074yNCjn7cZcci23SRHq4EiC4d2ebPnHy751yEIQvclFIPMLDax0
7VzDhzm1O9h+JEGHmcY08BundWHhaljl6XcQHQzghRBDyIpk8HqguhOXSLzW
SHVcI1T8fABxAOeAAX0aCsEPSQPRdM1Q+MhbyVzBTcz3vi+y1YEEr+JPv/NF
f9bfudNXXbjCNyVTrKtCyfJqDT2La0229uiWnJuoc4Sa1WNnrJIz5Cui9tgP
dF+U8mIWIIFHcHcF/obqbo7ttFaf+zRcy3D28Zsz65kil+WK0JiQNJDyz28A
D3K1txJYgMwu5206MqYTp8lwYjd3osDcyb4du5FM+MoHxGogSFd3hHKfSnIl
1mVWp9JOvFZvd5KidzvNSFsOLvjJzmtQEN7z4Y/9bUT5Ys78VLGV0oKrANib
VcML6yXu9MKYvjnfkuB0cBMH6fsaE2jOZOMaksKESNySmvC2zVFVGmsDiOvo
gIIV7Tb+LpbkGvP4+pHZF2a5HrTntTUP4goy8vEOsWZ4u47V2ncR+l3ntDx3
75ESeQ0zAZ21NBWrlMohJqAbeg6E0zY8wmxNK6ojx1m8f/mxrX/IQREqNepz
F7NvW6Ra9Gq9+3pSuAFW3KrGXMO9Nhr5TEoOenbtTAlxB6BeGn7L8fFks/bJ
WRGB0lo5yYR+SjcQZ24rLlSWkzA//AKRf8v04sFpmYnygEnMlytK5dEd8NLR
cy8v3N6AU4HCilw3XL7iAHT/K54FdVrdrwSSQyikcle/YYvnzq/dz04wwDTZ
0OG/RTzeTAHzJ692B15d5/nfNg821oQj1h0t1CyBZqARrArGvdFOdoVIw1Oq
3AANuS5yQ0Ntcq//iUp5zDHRBp968axMqyyEHa2JoXX/zNa4snS5SmsQctVc
y0dFoS9yiRO6fER43RZ1uQzhWOlR3uJRsUgEqm6Cf2xR1XWW7xCnacCpn59k
9SEFnfAyHqKo72LpiaGJscem0kAvOQoFgRMkUCnKWgVx2NzEGgNssuLrbRQP
xqN5InrAAWA23kGmy3RijZ6t0tt+SuWh7riO2PWir6jIQa2nhqM2DbqSGyRZ
K69QIL85SI655uh3VfnkjxNZ1OwgN09ltdEYXPvxGpeLk0v3oGn17G+/TSeH
OdLvZPJfdz2RQvQIxo+WBor9rKkqAVeKV8q5fU0veOziyisNbmGdj+eBa46x
ZSSDonhRFBT/CxrWMQ7Wr3kIaTy6zSLxKTsS9QhTzx3FVewSJ6dCjKSvpqPN
KlWyqKA75/r2CBDmtKGALqGuG60+myNKNDvTqIaM4PDWpfen40nnDBwg2qBK
u8xmZwZAGE4fRsDhvYQexC8c5sQfiAIaTB+PIAgPUlWDZEjt0mAFE3azGEEQ
Vu7DMHdjy5uYLSB1Elj8Q3eIdYM/yRT7XWRGTrFMDGuxofueMNms79jneSoE
sBQU12Uyu6y0mf6zrx/Kory/QYBb9asO1JbGqdpStK95nZiltBfMSo4apFua
P3+jb5WxOQ9D76anhf0gmDVdSH+eBIFV3SZsT9n6CCsRt/uy49sYtbkB6dCZ
H5TJUO4W7hQ2/dB/HV+P71ZR5WWNJP8fm0tqewUO6srjM0MzbbcczJ6OLLSz
rXu0rE3NHMZtxFBtp4Zrmvv9Pvi4stuvXZZkBKPH/00TgsLYZRZzydxRQ2Vk
rIcEeSO+vyG6Z09R5HuUVZwcGD95i9lOKjuTY0f5TLY2bTAF+Vy/zT1PcydZ
rAX/99gTBkeTUJ26rMbDafL4uuEnJctCkWBmEGEbAN/yjxDQ4YVN5tO00ihH
xALnse1mTRvc4pyEswXQGe7RdwbZeq4PHom50AgxnFrCbzsgftvPjGBBVq7j
OjP7pBCBrYWw8kHExOUpkWdU45VV8IxkPq6JTfTaQb6nmZGrz8F32c7G5tT/
6+MKRij8251z7qHqJyLyEjYN4JxIayLlh9elLWwdYo2xZ4Z5godSU1ODqsis
5T+Np1Qhas5lD7qozln8GSqTpfuc5rm/nxtyXFIpjO95irFNa6SxTvkB6Zjh
vahx3cgW4y/D+3m19KoPvWRwj6zgjfRLGTCKJUnplCjKxlPeuDSBEsnzfxC6
78E+16BeF7HQscuAgUGwPVEwOB1UIYhmivTNgeVb+EiyQROsWG/BaGbkjmDX
Rm0PGqyFg9JydpOBM2iDeqArhQx0Nd8yEld4Qq8p1xSObKy54D2YajlPet+9
R/RbRASvKPyaG/PGXzsrX4DfgbhdPWhdEG18wbm5dNgvDUUnupAazGgRqyr8
hd498egOjT12HCnOlZbNgCx/sucXOrY/m2LohLMcwJGvow92qYF11IpN08/a
pGfyhpX/JyI68e2JrZwDvjpcfm3ZAm3/Ka8k2+gTGI0x96JsjhEp9g29Hrvd
Wcv+28saMlvyeFrq1sScXOxQK7JKFIOzGtbVvpmiZ8BIG/4VjSi3d8kEgF8j
Ly0vWamxjYAxLoz+FqD9eHGHq8021eBUdN8JHap5uXmEXWi3Sv3gqdtPIVtx
gCA+4lDVo9ell81+fOtBGihMtkPfiTaIpG1kshFq3S7UYmoUJGnNpaC1AJ+r
COaFNMzAhhG/h4B0B1ewAW660KDGZzk/D5/ykWLUT9QmIq6MlzD1wYLX5wQ7
1jX8/edme5ayeCDYkSBv6kmGsAvCyBh/OSAD1rDGyntDyQcx0ecfjLgWgW8c
bWHEI2rGl8XsiSFdQ2gbD7nEFn+FkVhsziVqL2C7ot2VpkGJaE5ejK+8vIOZ
c8SmXCcBaTwG0iuaVYbCB2V6KORwnerz94pi4FmDcfHkcm7NySJfZiYfYReB
aDQkl4Pq3NUMIutUN98NLH8q/jQr1erwtH+EpACQecst8umLh2dixBRr1+j5
3F9P1uuScgATiXGmtwMTtRPBYlZ09f42lNcU3Sh3A3tVEYofq0HjFoVf2Vio
aBNqysrM3DUtU4pXjGd4P260BmtJbQn2fufrGCGiXu86hBm5o4K5eWIYeoU4
YF4AV5mlZi5q+mtmpdS9QjazTk1KtJLGfd7E7rByn5h74nx0gTX/LXu/VDoG
NuX3c/+TRTpGLtHOVVojdcQBIRbhbXPeGJTOl2tKFALcgi8C+difwrunGT6F
REQldZ+wfpBsU2EVhAjoSOInyBWHzJ7h2fwTXhhu/mbtcZcFOS/dU0tEXeuY
xvXsydq5pdgVDmermBm1LCOJ0R0OpsUJgTMVeCCxgXrNSMnnPjIEmBzAYsQB
oEItrFCXPtDw6bDdkfn4Fx+i1LftPIodjQi22dRxUvCtXksnvvogWSJ7I3Uk
O/IH/Y4aHgTgNZDx9RO8K3BdXhbyLl0zq/DmOgdMf7s9hZONLYhvM2UQaBYh
IwCGdzlctaXe63292HVtlCQjxed/idhK21yUKyu+DoEYp4LfRzJxA9w9tnk+
lAOXUZ9OcOxWbHc72UhWwAfAccjd0JiTwCuUxaRPi7yeQJGw5FJy6Vgt+jZU
CDGOwf4ww97gywdODOdjg1ERcN4VqOopBWFXeA+0Up9LaevZzxtPATQneadW
fFEmnmIK3Ix3pvdWpadJESCCi8nSITjQyLToKA3h9qvLizmfijACs0bmeJS5
1AlWsF1WT8mTxfUs+VGn0Fu6NVEqLchLfKxSmkDzN9IUpzgxIx1CQtQIjVUX
yo/+9v6pCKPvxOMiJtDS3bMJoSwTNZylWMMpxq0KkUqpyrxlu9s9oCKBDoAR
1pBsLWYIp+l1vCx7OkWk5LgIFy4gPopT4tTEUVjfilcdK8rZ30Z9cwOS+29U
BVgBiNTWVS1hwj1lkyzsfXW5iOe95IWJWwWsRvoThYXUNab4mVElgO9gw6js
Yc3Ebx53JLP5LBoYWOZfs4MWWpZvVNaD1Eg6hJELrOjMCKGbDoXOLbGBVjqF
7xHZIZ78Qis5TUEgovWhtMtaFe5N7cCNp5GyyvWI5tRbhV5VYhrZOWUJ53hk
Fj0dnZFC/9kYYCRVWiJe95dqgTz2y4jNOjeAvvHhoPjU4lhzRdQ/IHYIHGqq
wwYKUiStUKgJyOLEJy0VhLPCO2sj5ewxPnlTC4EiMYUokTCH8vqh0y/4TGpj
uE81clEdIp2mqXnjj+7jIQmd8aAz5WTLGKSXwgRUqWcm8ntr3lSm3OqrKuUV
WXHuELW4z4s1DBZy0UuOLFqLlDjMciA3C61NdWYqE78xODBI4gj43pkMrsA9
YDmDp55WHyAQbJDG7SMdayDshBNysBhox33M2KfyK2Q3K/8L/MKLT5fxChXb
dIC4GTP62azrfm0Gt0K/o45uP3ad+6a1bOGVMgsTUFUFTbNXmUs2VpQtFLgp
XPLIAq5Ev87Zm4rVaKflrwDxb+4vjdInD5JVGO24UX5x/PZDFAs+p22L7gZ4
UAnpHKlQtj89WT5pYneTkEbz/t413b4Lnqf97cXyf7xo9vcDZz6JGON3SMHi
lz/JWj8tXtu1RIhcqe75U1cq0nGbfo0/mL8iD8DYg8aXiQSlLLbC3CvXunaP
M+fFDRlORHgXO3vpsdlkiVvQUPvvJ9mVQ6V5VFgb9AVQza6uL4nCWseSZGFH
xOnaBuKhaGoW6ibIoWJfqcb5CREXQi2qk7TO0pewPPG+RzVQtQ4oMvpoyyqO
zzBjYRr7+6pLq7TWwP+zZweibcle9D/rktfeaO0BCqx9ufngcNGOQCAvENDw
1fFS1vFBKbk00wrxsCTegJJOyBMuReV4aiWMBaChDSZsWPP/GeaCb+nc6Vn3
GLKUah1mx+3t25egFigY4pPhD31Wut/CTewmf9w6wepyVG922rhwkUAa6dYP
5nRknohjh62tjnJU7bvGVnlfsoA2htLIQzxL+PwvtSEGleMO/MTHx4E0b+fv
jXtOETkv0oeejF5OKueMZEJnFsxxrlMZnTyLg+waFwMFeCY4mB/pk98M8wMu
6Qq5Jlx4kVMrl8Mjxa6zF+xbMU0Cb7hkOW/OPFwA2GsCqN6xL+PNZj31PBhv
DUYcFhRh70PbedRa5JuXo13QjpQDDrZSc8ZcGnkcnqcr5jHbKQJDMi6DqLn+
eG1sZYJe/OO/A1ptrI5DwS1c5EYgfs8RjOU4iaeu19Va1zLNdmrJAwCTBEU/
BPjXlxBQhyGJvUoa6PVC+AzR1Ir2Loktzt/E7VSWz9V2vwBPjsKMNL2Les3D
hoBOk0u0rdaXEr4gf1UQ+SrHGHR1nYn7SkoL7Im6BQNIHwlZxeeaBIFEhuMq
IIbuMrMed/TK/r8Ihg6SqEcZdlPn9a3vmPh2FHDF53F5TmIbOEpGq52K0u2i
wA28+t8tZdRiy3AeQfsdp3iJkVVRU56YrmFwMrCJAexXpfzzXV95p/fQuikb
2VKu0WBsaV15jp5BgKN7xD7lB92tFKQ01Dh4zY3gzDUPnXcPLSOGr+q4onHd
wrLpdqK7UlIUMsgK0tmmBQs9Mc2cvgGAelYn1SFR58oCtqS/T1ZSqDKVFc1C
L5mb2fCRoLmT8KZPrdBTF70Uq7tAjX0VpGfbIkwJH80whucx6bBGPTM55EIV
QZ543ItUHTICKjWmCEPlWgku4Xscd8Jogf5CSwah0y+OK0//wYnyYMJbAAdd
lZYSsVJxn+2yXNWhU8rWFMveKatXU+6vH/9dIioe/TH6VRyWWCutzpBSioe+
vFi20xZWXoEDw5indxo4BwwfFgqkLZpBmLeH33BStbQDkb+/yA3vLWLbanSm
eWUHbT1iArvijPivqrmAQc0mq4zvhhXRcSczCDun0PoklIMNG5srCJlkf4m6
mtP1uJrhNMl517y49lBi0vJTiiJQTIIu9mHmfX22Lrbq7FU2tQXgWv/4XORH
lZNYEUzC90HHzTNz6pWsvQdl0eVVX6fk7hBhCCjsyn4Fg8MYHmBdbsxom0mJ
763BRDZ3H9Tv6xYZPJevAQdF271/z5v7fKAhnxEavldqZ/8Akz68dYi1W9ju
YhwWEXZzedqYareE15wnXow6Mbk00ty88N8oYEUxlKbzai3BQTm01ai2i2F3
DmghH0a28cfmeQwFwywJ46UOyRZOTrkFG7TT6RX732pYigjBLOkMS3B1gQqa
f2USM3rdRJMRoQkwS26umjB3j+qwal3/GvNbNkfpWXtGhy5REg6ry/xju/wS
qg9iS5TevEFUCueXD4Hg3aPsf/RODruPGHiq5fY97uz8IUrUWLzxUPSBWN+W
e+iKyIlseI/nd/shIR97YXNVANpJ4hg6uNOELFjZ0HMxcUk7R9U7IQsyTyjk
f4TmUbpftuJUdT7QvdD4pU+S3ov/gXloGOatUngNepBukgwQCNnE4z3Pmpq7
GgmT1v8lUAfFMrkcFG75VgnfQMDtjdwjBYZLPo0lwP8S/jyQxiedTPuHgcEg
cC4/bMk5TCwRqS8TPa3kxpqqoMWWscpD3RQAO9kEZoRGy6g9F6bDuP9mZFyD
kI6AhDDLkRCbZUSzoevG64rOGeVN2g7Y8Xh8LujUVsoZt70H/b8KOhm/gXjb
e+6vaxHQBvpWUAq3kxXTyL+oeqtbB8M3a4tZr/zJ7hcADdKqp+fvLGPyDAdl
1mVfzWtWRxRo6jjjihOQz1B1Ktt3Pe5SrlJ1bPm09y80dhDbzvKmq7OXl49S
aG7VSsZdZ28WgLwXOEK6kq1YFxXU0uL2RzN1xCv2LYRpKTc6ot2PuKVqBZAj
7fZsZXaXIK5r63YmdK7Xhn2DgIxe0/fuh8h1N+d1UHtVnYOAYmky+OoG/nye
7IoFqJe1hUMJM3UCe4mjN5vVkCw7py27kBc6rabHfdzQMwvWiTmruKPAVAkm
fUUipn5Pp0p17W8YlNMmwUILVaSJ9vysHl8U4VdAGRUSdvXbPtpGdL+Wmm4R
BBoIYxCM9Cif0s3DoRnSfXDFU2ZmEoXlAK/K0SbfD2cR2EWT0efk7rwZKf+6
uTJ01DlxsJlpfcLWiZyU34lZOutTznNwVywZO7r1qurSw5LQMVyvnfMbQW8f
Z7quPW4eGL949B3cx5AdCs56r2SOcBsSH8Q9SEFxkBisBe57tx+6Y8eczI35
C6AGeXgoVV8rVTaRU5crm5JOgMkgGiDw5UlZVSub/exBZGAm/so2ncUuLiHd
WobUF1dDrMJpstK9xPa5IDoWLsQ3JWpsX44Jw9wVs78Y6FBUdFm2oAC7l7z6
8UNgGf7vHYrGIRm9AzextHmM3w11Mzj3ymoQhg50KtTIkdOJ3crprUTVRKfb
FDeUVG4zPLgcE6gVERI26TGP/vphaTFgAjBqkb62zF3lJDU/z2Y+/N44SHEN
UW3DQFwSnpm+kX9kuu8BYBOf89h3m6JZ2qewIJIPo0WTzzH3fcuoYAclnweG
2EJJ6Y57GzMsIisotOLmVOg3IyHIXNic7uiI7eE//8o/VkwbmJze41TGITva
HvibxozTBsQI98z344thFateS3zljDGae3Ue3EG8ahL58mioqdHkpK/0h1MJ
3/rLPttFSknFn+ZgY2rni6RLsNqlhg06DUM7IxHEA2ZfrEybe2U59cr64Xel
hNJaVxWu+JEotXMOKNN+EVePiMeiI+zEwR/xiXxJPZLYB+NBYeuuXtCY5UdY
VLqnMw+96MIoiqFB79R9RcSDsk6JHK5Sta8urHv5iTSDP1sAdq+oNu8LYXbu
deFXOGQE+ERrspKanYpaXEDCu955BUQH2JwGdR1pAPlsd3kVACO+BSVULZOn
V3dB/85mGemZ9xmDiBqAwUYXMnQb8C48YvRGTh95YYVVovP+OL5rbKOqtNUu
2d6BTlnqdzrcDOwNppdzZxn1Rvpv08fzGwpgQj5nADYyHxE8zaVNMqm8bb20
eiqpFxYcY3eoYs0SskM2obdTWFoRpVY+Pad7ezg54cXS8PdJiWR3wop4YiEy
ElWo9ckVZLsfixOIlujUkYLn+45GopHxP4QZKdvqlME9ISabAvz3UStGg/BP
+BcAK7Z4wjZLEbRYasZdj1R45r80wck2N2g3gF4/874zv47MicaY5lo22OBv
qEd5I+km6FZIUOGL+R73NwpNRJHocIsjgEzG4iwNdlJw3J8uoJbe39GzUC09
KnBKUbijFxAjai7k0B7YREOuKP0aglRC+TYKNInSRajsP9g7GmHT3/78r3v3
BaS7Oumb3PRC1h32GgAbsi0MVRxPjAYj47JfQg56D9qvLxW1EXXMcMOBo/Li
AKMbrEhO+o2CsxjjgmpWJbS+NooRElnogMvGl6LS0Z+QtpXl5pnmnUJ0iGUD
zp6RyX7BmAff2Jx/J8DkYkiZ96AJvMwA1/zbUo2HZhoMLBRDfTJ+LXc/6xGu
yvo45MxCLILaf+VZc5HHbrEIZHIXwxK0VW9vXlfHwlPzt5bbDSMc4ccaHBWD
GaO3oZpRrclZFVLbSwS0bqJ8D/AQI/tjj9Yi83VYfY5g53v6cnKah+WqIWRI
GnL3NxUxFdMKNr0RqdYkUhDu3IX1jLqVQ9PqcmKw0EI0DI5giIZmGkgvMUVJ
GH9/2IgbxFM7MmWzLwb6wv0prrp/H8AokUu+RJbYuGG/o6K+Mh1ITD2/DsYR
BpEskY9rohzs7Aw+kVdguksgwbz/KZQ/nGf3u2CE8rWNJkhcm0713ZE/T7Ml
FVLYrH/jTz589MYIb4M4ficsXW2iD2zxkzZBT9CUW6vzZHXFY0zMUJQayNvX
+Y98QrTh0M7eUK6WJd4NxMCMtQN/2LSLmD8ngQ+im/o8b5F47e0fh2hgAvF/
4x11lNNgNOD0obF1oNWf0WVcz1GMKXLDuq+M1Gmvf6iZsG2c3XjGD14LUQzG
T63ekKOqK8tSXxpqGX+AGW0qfvPZ2MAQfuzaIy683G7d5X/HJ/yuqApUoHVj
MobIVX9IqNBJvUgqzkjhAqaAkxlfa213lhqlvWHp1W86Ecd3uO4T9HSShyrW
2Hi0NXHLqm75RDYQiT0ED4rPN00LyTveYctdlNSbuwl64MMr+3E7CdpFLqMk
N81+xT7fazo85dWP8ltbCqn2oUzyWuu+5yckdg1vO3kAxlH9K5rvqlSsYKu0
O4yD6I3wRV3H9iMR8fvrrOkpwUdCX5t+3hobIrbmlL7FGaXe2jbxDIoXJDwa
V9gTYw7+8L8CpUi41xYjHo4Qv6eOWFNPpNxxgGxYDn+BvR1sFASMXaKcDayI
GXUN2tSOvaZ3Isq+xaIMqloAjrJiX8Pei2fH4fzsdwUw+hIjK+R3rW7jIQ+p
3zoR+HenmZGdaCie2rtYjVVYRWWH5ZQHuc8qEqRv9n55ePlDI31Na3Vm2tkk
ZOp8VLb2jsZMoHbo/j+Gduv/NGIFyuEwUcXDxkHVNffAiYDqVt7PCTIll5B0
dQSVg8l1G158e1Mgysme4eI/+qr0SD+fOnMza6yy0VxPQeBlYNKTe8Q2vtXB
Z4lllHOQM0CRI57qi+c5K1az5eOMdpEW0+qgrpX45tJ6CXXfK7tkkovMbnpG
WkFLAldhbq8suIjizPkNBmLxYLpqClQ/N6OWqXGI+e6xyr03tuhSCSZZiAoK
FjU1J8FTh4JEU+6GrLeBlZH8uQ0gdN36d65lM8lvOFZhEKcdIp9SJepLMKrK
ZsufKicWTTXlcKd1igX8lIHaHG0k2j0L6r3LsEXCaHeXbp0A+x58Z0zVUXG9
iEdeippIUZhJCmYv3SQSz+78QlgVj58XFs+rTKh1CXx3KpsSnaGrAEFr+72h
sXl1WzRR7hzX6fHXc1885znAZ2ONAAiYiqh/0gvo/H+OM9oXQ+ceXErsce4N
kEf/UoK0hsJYO2sqNfkKEDBQr683TQp8bSb0mPyTXTpsB8gMa3khp1Au30xa
HLltXau2g3p3UsEioi2G/S5ycLRdv0IeiF4k5fLHWGwelWwtP5SYBvNC9MSa
f7TnTpk+JcqFtk0mQqxAfV1O+0nphxMg7lvARWTkmCNPioFfcqZMZ0v7Mn+M
/cZKMjqTzbnAW0Du916FGPoELV6FGmsv1KPRC66QtZiGCWlSDbeAv+GQ3vqt
xHM0g0yvt6JlQDWEz5KRCYKZv57Th1rq35djleCGZllYZ1zZZwY7NdPsEhPZ
RejtmUt66byK/FU7DkfuNXQbmDhu8zBEy5dhzX5SF02zDhhd3gpJHEgtWZs/
SzH4L9BfmXdF+qje4V/3TMGhYBXwQ3huGlsTEzhnMbr8lv7nzOGn27/94Ldh
epc1XtYHiTKjc2J9xDW4HWdiJE4zx3Uy8PCMcjPli5WPjuzqIyRFVSdevxXU
7mB03Zuf9deZGd9/wF2rNk+Y1whDO1bA0yWPxnPOH+iLpQo09HCLHkp7Q/AB
fKaLSxwGuX+DgqnXONkpKtSekzvzkanaOfoLlZohUZIBpHX+Vax6DbK+AkeA
wwD3lrhLzB9hKSeL/Z4IqcM/KZAjaX+E6RZZQwiql64hAApabqZbZ302H+UP
SGBBZyCkApL7vX7ogfcRcMokceWBxNOXDwo1BH2avRLLzj2j3LM0E3BsNuNL
y3XUIZCTTHje8VxkLp7EU2P36oUKgOYluofvCVqY3Tx35A0K19dIzdLyUX47
scv8mZ/4MNTrzvCSQfr04k0mfiXdloQnwAGrgihlLB+WIys/sTwwVK2NpE4j
nX/zkvzcNUWa6TRK/7mJLYbO9v6fONuwa1vM2MMs+vBnLx92Wb9uiHYy0wMp
JskBVjN+HJ/J/4Pl3rlcrP2RchK/yovUU+Lum6MoaDHKrqH+uXzSPnYnEW1Z
bGhW4xpeJZkInzt27+CDQispqSteJ/ntUzQXnGMCuPhgM9i5EaA4DFowSog1
5n7KYYgDLSQauYo0LLpmwyQOFw3d35Gcs0Dr9nGW3n7ZkdV2ivp4ZxUoxc8I
5xhCtVBiVajxOGumNsGBrL0i4r0dSzoYQNjoJIxKAJAWjVX6PslV2YgbSUBo
MYYDycew+7GGFEGzVVoLYswrslA6UHBu8OdAyMRdqUslQS86aCBUjEP7UzKe
3GDWESINrZcFZQuKdVoWt7JnnluBOWYICEHNBkGugik166qjO9QNJKOH0AcD
YMbj83B6clc0fmvjOwL2+eDY7NhsrncTh0C2Sqiwt43G5Z4CvMpiCZuonR3u
jKOT3visVg0Oq6fBNInL0X09F5GxZ/nqkkmX8QqAW+YnT887yXrVaFGedtSa
87cim0f/Bq5J5bW4tyRPQm9gLZsVt5+63cBa7ZePWnq3CxT103mRrJE06zx3
jIf5bFvDUKr4fUif9pg4bqQq/D0pnwfbqH0ibKSi+g+kqTsWCG3qCSwYhP/V
fXC9JMsYDy3qW8VN9ZlFWfAZjzWNMiQObGRpGDmpFCPzJaGXB6CJUEchDj4K
T5SXRo8GWbQIdFmLV7vifNmu+6SK7OUEwD6IJ7Wtp0htUNQKQHUvHtbOfwap
OBIzwR58nHM3VL3N13kcFHr3wiOyKjtg/Tegmwos09u2jVicB7lVP+Llpjeu
g+EhiTQKtA7dLkFzzNcm2qkmjDMVJDAPSkYNqYQeuETKqnkcO7WT5zzd0aFl
PZ0PshWMas/V4Ft3p67hCaZ6jjxrV4PPu+N5dISUrNvNsTkEXijeGg9vI3hO
FtOYZQK/yv/PET0iAY+GwWYCO4RxereKTgTp7xuXpCcJ3MyxZ6ydHhzy5+0P
NBfXrQllOO9nBGe6mPxQhAMbx3D/X5GV3QmSj6MmNXUEOopz37JypEUHvyC3
xVYettJOrcmJv0u8pSin0Y3sdAy9L3RXGDbkTwUfgzfPLmja4gbvuvshdW/R
RR6LdQefJNLx9ttRiv4uOi45bHdSeUK98DMcOV43qKQzK7lwU7kjQZZpgRUs
rrmlRH8lO6pbx0MjApQAhnNq6/2sbqn7WYIRXkrf3h8HdEhjhW1X7EBmf+wS
PYjE1vAC+nVKQ27ZHeQNZ4GJm6DlnzI8HZEIYUhzMSm7mCwE2a5DhyF6uIkW
sTHcHaf05q6UT+elX5N3VFs4ZH+UOhjKza1weeZjaVmVOczRIbzokjIvYxCZ
gywhjUxw5jtZIw063R/VB7Gxi8e3vEgigr/DoW8A1ENomAhWQQHjxPPUW/fz
8azi0RwZbn+F1Iu6qg3wiHks4mmL9JJiiy62aSYHa8/HoiGHdROySbsLX6xC
aE+03bdY51U2rMHDv8w1CGnOQRtS449fyd2kCdgwLjPhX0c2dkIC5VQBh4fG
eCQIvY8tf5RTkjk1uv/OL9OBmKRfHFevBEXcT9pkg/Q7PvO7baY5IZWWZIjc
8/pnxctUQKgDaRvoljGwDQth263Y6EezwpUWiHgNiv3TJ353KmahC/wdawNK
7fcS9Aehozs1X/1i3b+oXCMvj7WqgikQO/4kisVA/SwyNWxtuHTt3AAaYGbe
f3rfUuAdAG7siYQRv0EfFWA3D6eagHHCycfubiwXhqh89pf4rKdZT38haO4p
yJLJu1UH+5DGyDLnqndj45wGSvbOAdp4G7FIw14M7MvGM1BdzRn9UkgDM4zk
mHo7cUKxj/9ATNeklc+EoBTbOXVKu1QWYwG8nNSsnaI1cvQX2CuJTQvgyokX
EHQ49eYTdFeT1gvqgetU5HA57zHcHLnI35JB4R2u/s8ZHSEhkdWfwzvxSpEr
4oFpv7UiQ20xlpMI5GabAeGvs9K9eQHYWqW1e4XDMeF6IAVOcwscqmmCQkP6
niaHNudj247QoNJovtnd23ksO17qkihAya66PX8B0D8iIzGHVqVD0VUuSObq
/L2mzUpiA2VZevnZs9iAl2LWcHtNj9qbQTfHLbHfaOKaduer/tBKQJjkFVnY
aJkC+s8g6We0cqvvDuiEUEbM0y0p7gL/rYBCs7J/unH87TEEzVGRoX0JOMNZ
GlilKnwoMBby5/AD8u+W4IOWTclxkP6bcXdUxGt30RnL9KQ9wgGqrop7QMBS
JpfO2HHo4yBoHEa42ZXp+Wy0hiBWW82IV64rWeada4SQIG3ot77Q88XRDW3z
TriFBuShLzzAWnsPGcnF+pHp0hDcXj4IzSnU5L10egc/BJRUb5DbBPrDuY6I
7Na81j3YKSTM1ICEk+jzzxP4MyJK6AfeRvev2ufudi7wej3lG70UBWgEZhAe
1jd8YE5FD/75U73NZnmC2IZA+ct+TuUwGjY1Dr9gLPKJkVKoXrE3pE77dNu8
rCggZhIH6Ztwd9tveKSmdIWKmbVA0nnTOFUKfVe0+oq873gYiFBd3WtWB5mA
//Ug8agWVG4oPhe0oRpMCcBV1D3ayd7QLrDvCP8RbdGMWhL6KRUIJptS8jtc
1ISjFaqzYhomxsnQsCwmfDAlVwQ/aczXAilX0eKBw0RIIT1dcWlACY0ZhHEZ
qHhbITbEY7ZOJa934kahJLy/XoTeoPgv63M9cgCBiIxT2XQomvfgTvJ1YVbM
m6RQ0+n6p+wkIXUhqXIWXd+eLxHfXAFP2xeGYU50uPN8SXzB0E6ZU94K6riU
VI2eGLjaIGYOTMdlKM7FRh7njJphwhuq/RiKmWc7XjKghoPCwISOnLIDNVzd
gkMlmtoIOdFj4KuVECJ2einvqhYwWk0GxXLpUlV6l2fBbxSuntRExxImjz99
YcIWebt7Nftm1Txwe4lBVhBdyuJzIx7z9hqSo5fl9q3oz+dZMcZQIC3DrIvH
0bdOL6gY83cO61lMc9pmMCTGvSqTOY+jdlB9N5JbUMNqO5GhKCPhDCeXI7pN
TWrWcAbRRnBaTvV1pKf6Ikj6BVHSjuOa42ia9+JMLNCuHLD22Nd5xY0erkpW
N8ajPx4t0FtQLtSAjcZqarqDrED2uPXV+uYzf4xdtcdzV2ceuGv8xhyoOtM0
LHm4xQbPG3GU/Gz8U8KgImD5Dp5HQ5WXCCT8gtRj9m3QbH4HnO6fNNgA67af
D3ZIENG0uZgSnySC8/TFPxC/kupxANV004mw0KibohEDVOJ2t0ym9sVJxCbt
E+NCiBUuNRpV1yEgFLr1l95TyiNgJTGU8847zrVhwEEv3lgTpKh5mkE0rFGt
WrvhYtnQ1dNnpRIX/U4FXWFCwpe5tWoBtmLPovhUfdkKqsn6hN73E0MZjezt
gXc6dH1niotDHXDB73U046fgHdnooLf4qNeQqtGhCXO5MXxPwgw4WyMIReAd
5Xj+L/PLsw0GMhe+ElSmFdWNr2eAWbkDN+A0Zwz5jnsabLR+ZJwqxfXaYeF8
Luc2MP6/6E4DwLL98vU0+PYpI3MdEGJVi2JUMV/r6rtxrzQPxDZDtYN3PFTw
DVK/MMIsaUFfOY4VZElW3Rpqwy7Nm7rL9UepIyI8l5J3KCVGPH3rMFD8yk6b
zvDmYwAT9PKWodio5ubQnKrlsRrZwdH5Bn+CTUt7ho8evIgyb1gWjLCsKnPC
zvxhZZzohHiWR+F9s+Y3JbBQ6IRlrFfm2Lea8QLNDCA9W9H8c35dvLGAyBcc
pp0hnUVZDbC3ZvSWQ31KeqxPDNah0HuBvspl+YN+/kgscv/ihORIgAjhjE+l
fxQ8AlyKLp1R0n7DfYT5ZPwSaE75CKoU74CGvYL0qt1ltwFwpLgS3KFeZNEy
Gxk+IgD56FMHyRlkzJ/1XXGoJHoXXeqrgVy4ETwqKtiblSsBWP8O3sDs3a4m
Cngw7PIxt6Whsp9zq70OukUTKpMSekhJlOoKYpoVgD27iIsg9VnmvT5iuMDI
jcFz38gFwv0nONObp9ycXMY6bAQfe+IxvoJvy8x/xE1swr3lCyH89/EhKhIq
r0vG+G48q7nsAk5Z1ITs/oFkjoAbwUeKsNK+qaRofr2r5TbB7f4SmLsr/MPf
rBHP6HgGxkGh+cJF/c4BAUzdY8mL7qOM3+x1qGuFnF2BqtqXo7+mb6AFyy0D
OZOCGM/kCdIkXSwGxOryz6g1q72Mv4Y6Uc7Dj2lbill+ECz1S9qDGL/Z4PRf
Yl5jPoSq9maGR/IGvUME2rXyepF2JyOkuRDvRWebnmC+mLZ1Z8c2lDniWlCb
OTDT2HzqyOE4Yo7O2VbVrbgYmZwQ7x5RJHWA60BV6zAXmONH/z7g/gYBKUPi
JfTaAVtydAil5+KRdwqP0ZwnJRM90a4FyjXAOHf/CqBIKDn5T9GOisyac/h5
um3ethN2CURKxu7LHP21R8z/EllLaVv8R5J0l8kMLEGcCJzU7cS8nCT1mC60
XJSEmRs8rmidvBKNdsuhHy3ukegnNBeVmkfEDnJfrMqzkPmtax/W3inj3oxf
SWEjESHrTaKB8EhkewvInoZIze/Q73Yekz0phhAqVa+P7RWWYFGclDDp9THT
qvrhoOZG6Dfy0avEnS/KlUANd6S9qtcC1FqF8Gs8GCxvlWa6sZJjCt7rEJkg
zBVjowqcFAUHcG2t3N7DtotZYEM+3cOMhXObSKAv8fnRwRyqeyyoTZq3//m1
s37g0m7ArDqxRFre2/P0clrHE3Up9YhcLlNRiWASaVb+noE8RBQQKXjHdGSF
ADAAUGpyr24vpp3HyXqys1/oiQCcGQ/wHhAADbo2CNA9dnX+Bfh4D9mEkMwV
bDruJwwHAZb2MWPCzvqBw4I/coNicdyzPIPgkskn5YzInkdWrMnCoyOCDgK0
uQ4fdq2M7iHAQnCJX0JTZgnQiwdTN+E+6mVQ93pJzPUilLl370ufWuckkYce
YkzMOmPB08DOiZ2XMrLsZqI+cweivSTPyV9sq94bJ0N2Jk37YX94hHzWsS2s
eOenmr6V5/GsXbwTwPL4r5Zn+ZM4rXE2+m78CGDrAQ3KAO8q13qTXGOzNCnv
+aAFPDm3vowl9MsS9Fljq4k6/9wsT/bsVW/cRKTsLjDjRkbpPmzV1SNNcXWT
oW/hsQGtFa7uUWYUg3v0zuaT2S16DRokwLI8no0UwqdsKPu/i8+GJ5f1maix
r3JqJChDj9yULZh1qywN4SilO54c8FiAB2WQsHaBOcGnhEjfegOvuGT8cM/W
Al3WkW+k6u0nmRuC0RjXivndNqSRXHXiflegeZdxXJR4qe1RCrSfEjNdP08a
bvHT8mxDIpTAUA2DVtCACl7NhKlNKkyLpYPdEBNxuPBeeCkcYkqfsY59IM0A
tbMV7C9o49/j7cRlQdB7UvwKJfInbk+PTSE0dtL0LW5bLQnkyxWV6ka6vLty
sCe4laJPRbYR6DAf/GsVjQitrFwlOLLrnHM+0oFpnEYpUJCQvv7C9deJdmDZ
s1iAFOf/3wS2hcsV6Iq2wWo5cXj4dVX8918BLIcHBnEZKQ7H+Cj4/F7mr18O
dN1ECR662Rs/GiMgdbMNKAkl8YDLLMtBG2vK5U9Ma7FDufXFcDWsjJSt4kru
AOHXqv6DU6j0b495xv6m+FrVTY7WNR8dO+KZHDtjuRq8QGGNXAH4njiQ94SQ
ATDqCrZWycBLmXgiaxNLkTNSOv/uSmaUeI7ROKZW8sRQ+3LNnW4x5MbjL/gH
9tUgljhao1vkoXwxDE8vu175iKZDggXDUE6f5RmwADp1cOF/OR7ZFz/x3IsL
Xkm2N2AkraUAh9iqq7LPgiCJEEVVOFT8MHcVz8bh07lfLtbQ9E1HtcHiAHMV
0QtZkgsyM0F7c/Bs5jCdMX0+oFH5l2kbFGuTHjjd+gksln95n5e5WuZBpJjv
LqF+XosvIVUFV3Q+vKRtdT4PKpEmicnWA2+4KkNdsqUno5+M8QZs1t407tsE
L83ZvXBU/9uYV7z2IZT+4ZcuK5SnkEsudJ/5mVziEkmELWpDRdEWOxAOwC3p
k//y5NwJd9dMP1jmH9OcPUSHHI+ZUTWDuCH/0X3RuOo/agLDjgnj9mUShcPH
JQIBy3y+IoYWXsTqe5TXlpVAXXLy/HwlDzLYR2PgwMnmn9QkEfrfscRAUa4/
vVOrLr2WxTjsOUjocj7xb7YWBdIyCeQBZLYAIzsVQlxyynqfW7/rcfFe2MQ/
+vlrE00BGqDWtVUM+KE7qozPkVajT02VL7ZrIjb++Lg895vF00b5jwmJaUU2
08GNsCyQQm3LBNsImJh618p8bpFJpJUZceI9BF5vuUrkYQ+zcS0Dt3ynX2wy
H9FRSeDKAghabbsSoe9XNVrmPKkMRgFr6qVurQa4BO9jdz+i1ISJpxGzGyIc
9zDaMd+z/n+Ct1zlJFeCEPo59mumNm1pW9mGgVC49uqBcx6PIVWspZ3tN3G5
0umEWcctOoHMJI8M0T6rOc8s4qVwxa1yCNXPYqFW5aYYKyRCz3Xh4yvQrqet
iiNyZMaYBQvJUus9L/sttGXoyT04jNNVbm9zLo72J1v2gS3G2JCUgBuM+dUl
FEJaO+ctaC0EhTnoAPpueEW2I260wxhwU1yqHFxsBDlc+juc14cmPVEsrBWD
QOIWePv6gCfMB/puQGJYlEgXbYrJkaNTSHhMVdA4pFzIRq8qglDDkoCgF0dH
MRZL3dRZJvqgYIRlsEO5QF9WWkG0TH5Ucx7iEsr9dshccLzrttfSw0q4RfPd
fgMI/YCzCFO1nP+JNznkb1Ov2NIKCADBu7iCKS1NNVf/8KNB0HcqWhVmPVK8
8qs0Z4cDgCQKUG1GwO1jkpGrWbwGLOvmDPzzjAxOv7v/dNAPKfyyqP3ZBwgP
OppIljnuW1rL482a2425OcTIdfu9zJKgiJ0jJ3A5zm88GljPZxG5SjFCGgt4
m889S7k0B082zhzL7dh/XYyiTaOakwZGHm+rFrW3q7lXVOjOq6c89lWMj4bj
qR5brWVjqp0AQTXAGsz7RxjFhup5RTvI7VUJrHrlb56j5X48UBT9SqKqK0SS
fZTiEezQyKYmw+1BZqdmCMobsJVqezD830eRy5sc4uGYRTkjLAzxbX5ajR5l
OPg+5Xz3l34hzqVVfEX5cyoqddTf0wrF57GPdLHsS7+v4c6dPL/zJANNiOXB
t6ZbIN3WxTthamZ8X+3F3PYqolkZ8aQaJaXKHzb8R0gOOR0kJV2wtWAh28/7
ueynt0U5H0tk+l+BU00YpRT4u7quKj2hIhrgs1I0uRC0DWH+qtSW5QD93xMb
0ErNg9L/oiW15KBRb1wJbJqHsacHVpEUT+dffOanr2EELKK4hiGBdXyzbfRR
AiESUaY7iHKPOxii2B1EG8GyGksCTJJ1oZeOMbxWpKhGBUCWJtZZlXTUT2dv
4rRktPeZpTMZnrOyHw029u7bfFzs6eMCC62gblAn0hrheekDkbdx/gpY5KMi
YO6ex27oMh76wO/uvbBUjJ0NPPM+nFlLz0VQfBBP311a2LdPbgc/HQqPeXG8
EX9sAJYoK2x0rxPFKuJJTU84j4/3zWneb5uFBy+CYj0OwEUQz9Ded7JGzpH8
yzL6wYyGE95aJYemQUPel2y8HL5i+q/gYwqTm3iQfsAT0YFChThjTB3FXxzS
c1YVSnAbrwbG762C50DZnE3hwmSQ/V79KGBGw3Vmpc35GvgwH/d96zqx5qr9
usQMe+SW41HfcvM3QxdHoaSYmOQIFbvyi3g12kHRbWwnXtgDrw2jXfWb5bAI
S9SurUdGJIj6ZSpJuHj66KDtaHDTkx5Z7BDkWapjXsxcs7bsQG2MOq4s+jdq
8NJaFzObDJ2bwIuRBLwqAbN9BHjN6GtQlkKiq2rjzzHOYX4tKhqSt5TQcrcr
h/YxNNIg+49t8Qrb1wM8cNZGX+lRqbYUpmpA9FvKb8tp7ArD0jeJv3jgkuCd
3b1nXj32ZnGxNkYC7r8hmkXoS/X5YwYydalG9FKrLNedjc2Jvr3dSGdniZU6
iodfVDv49HBCe8qYWHLm88g7Rv6v+LnfHmT86j/OePtvO+DCd8GkqwKoU8QF
sYMCzTEYcAxBwGok6OD7vVWSJev07xqlOQSdKEaZFyoQF+kyptRgL4iAYxH2
atcjzF08/YOeKDksWX8nXh7wI1Go3s6VXmYtDKmlURdkBJtyHY+I07+VjN0o
G0P1XSY9dbsTavzwzlC2UBkw7x+BHrh3b3PY1irA/GSP1DErHlHkr1fYrcyt
BO1o+l/X2xv9dzMW7Oe28LC8PBNMtGdrbTzFUDUeu+mCgBbQAcTnM0QoNL+u
cR6f4d3CUhN+W3ZLatkRhupOaPbqxmdMgV+Kp98rev+ODiV+8bAzssv+qrdp
tMzOLgmA/1v46Zr030k1qQRU4a6OwcK/5RIwGbAOhmVqnml6Th9/RwI3KE5w
vDfE67gKNXl/7tSeVFBTJfjCMjOV0X6425tWRhX6x7LLVMuQRLCRUd0ksc9Z
hBfYDayWAJq0WgcyIgVrbknn9XvMv5D3SCa1DOT1Pw9kW9mTPvV1L+3dW/Lq
vVa+peGhC0Qw7oXQT/AKfGxltHFVYE5tfCpyNPXWzNPFgcdHX+8kR69O707L
RVRY9iUqucTD4z2zHJxRpqz7z+cxU9qeDqR8nzwQRT6QTcCqxYMX8S/x224D
GYOoisCrkZuWcxFNURHhg3PMxD9uipqUAuq9PReE7K4dert8YSjndVGWHFG7
ecyM62mUAKwhSen2ut61Gai8OPMF4xUPkqZl4d/yBMB6TqTer0hftC9DCsCD
eIPoOBJ06X2MN+wi+Qc0Rq58LgaTqoTBdOyx0knUMqfhKgfbOst22StbIb+U
fO7qVeESyAIzbqRFkqouy5c0mgLK5faCFfnz3++zgvTXZv+ofEsQlSg3XQ6s
WJJThGy0ohlk89i5dQTjDFg/5R/VAYcY938yl/VDBSosk+ey2opq5OzcQ96U
Tl35NpHXoMcJphlrk6veIAPihoWoDjngTQc668lVFpp2OklAf2xUNpbeV0w0
Zn7r6b2GZEbXN/5DBRY+ac47y82iT5JslKuqw47MjCtjZsSak7yADMYL0Qyx
NwT0sMgryUfUSvKwaP6rS4HYH2nG4wPqkTjPzHSSmdIUpY2DfmYZLpMnQmr/
tepV5vkBxmAR9B5RsD6Q3Z5hidUIceGJd0pQ2FcdCLEvhVhMXJZJW12KstQ+
1PMXNMpms1K462J6XYju5b3pzc9SHAv3spgSN3GG8hu9yTmSCxujGnlcayxL
dURzJ2OdKxTa13oDs0QFJLwD0G0Ri+3rTlYVNfIajB6RV2707ySOMlBuFMVX
FJv+ItftD9m+RdDPpB7S6CLn6gHuPphhue+nSaIbVrM+n2RWUUCREyLYRb5G
XykRO7nm4R+0Bo/Rs01qN3bBjGsu4cpjGUenEq0G+OIE/pQ9hxPknrnPX3gT
1DqKA8oCvS5XL5Oyw3SqkgBIQIqrqDE5rQj64VJ53W2Q79fyTLc/mx58LqFX
+75+Yn0Xfcw2/a2i7l6tGcN2buGxt56cYDdGrd87rmHDaN69ZK4hAPfNFuuh
v+tqwWPPCMkV/205ZcQdoMh9tNYdfkUCjW3NSIcHgRv5BH8TgExZX4TewDz2
pPjO2kzysRvaGbgXFSdBx3vqh8ff4jGs/ofZwZDoep42x9vU0p+KX/kQWaLO
Y+/OuLLYIhEkEZ2MXexSUndHPMFNLw4rCFRnTurN4rCAYnOD3ffDKX0tmZQF
+Jai9NGQ/8Gi6Z6i2N92V/n0KCYeiXPcSrea9YyxEOsH0sxq7I1/mTJyiPUR
T/CW2FvPx5KMKkuUfEbG2SKvdrmGKEB0I9tvvVMItsVXOHuARsUIEacZOxpd
O+IU3/BkupsHzQb0e7gNIIJhXbpo+p+/J0EfFs/Q0Q1okqawqMcpjMOG3T34
AiFtbEjQOg/UfQenmCRAKQ5/5LZSYtPWwcng/DkFkTGm9wO1SL6SsPtbVJ83
HqG3IRtDiH4ouGR/X2WwoDF9UzoXqAyDJ6r8Q59HLQ77dIaD5lcx9AFDvzp9
r623E4NqC7ziFcZJkTyJoP84OAqQ0/nSOOdwMEQF6j/c6dp8iqTI3EZuHKmn
I9JMwZLCaF269jhAHvBp1l9yL6QS9nVVdUvgJPlbu2AGMj2bvOIKfWEpc41G
SM5UyZ8beGlJ2RvnTgLGkAi2UU3kUUWxpvKyUdhj+WbKUqBtiFx0b3r2maMR
jl56h7HQHqdPfKYxMZbYN4XLnUDGZK1Uud9NqiSWb1SGigW0L05+a1xEm7Br
sGWCcs5KejFsC24HmALM5j/IIQ3SrTRJvz1xs8DEd2Ubpoj2VQ8dvMczSj5A
MJgbY3z/O9Z+2zLcFl0uTkjx1iki0KVWgtDGT6Pm5VG3dAw4Q8hkT8OHReQB
hUOctUHRqmaMnBPR7j0ROB9hDDh7DXSVhifEu68JomQ1b3/f90PjETy1iW6J
eps5LK7Kth21Xy042d61bziyEqz9cKTPvAWn9Si3EoSBLNeZQZ8BKpq8QiSB
yqcns8Rs5I/HntI0uEH35SFbuEuoorrcieeyVnnKWFlZnbvaYQE6jPZaqKK8
X2hbBTHZS6Dsyx6aCmD2It56G/+lyjxswIjVW5chwGfals59TUga/yH1TxYD
sqjD5RncxJKQ1xYyMesAtiSpK1Vsm5y1VlIqlAaplEQArqRqsdKM9PygqcR4
Y7ZxHmQBvqhT56Y7ifRG6+Qix/GVVKvXGBTb1bD88HMuZlwAn4+n0rJhmCuA
4vGdxyPgjOmKVwZmnCqv6GgPQWnU9pGNZbrIxKmtlXRL0FyNZUC2vbBPdZdA
WqzYEWjnc0o7oJlsJpgWhYoBvcoGqY1D7GXtRVlcnpO3vzV6F0WDxr6unGlx
ImSLtsmlT2eRF6y5ArxBBniICRSuOTEs9ocfFm7SAul5Ftx2C+tDmJBJa8gi
xTLWr/GlXP8OXoEECcSIk+e0J98yp4oFKy4OTUJdz2u0VTKlFuhJj3mPZT05
SfWlSVCGvxXpgLgH+nelHagxz2EgD2cuFIFeYcKXEZ+BS36wNjWUkRKFcZy5
S0nFtzHU5R/3YeGz5JE1rXa6OYk/qGaDF8W8orr+dJvozXPNDSHCPDbAaCwm
tTObVuuniOL/na/jWtB6T2fZO0kDkFFxqmy/Rs+hjoW8V9e3CNq3DFoBW34f
Dhkf72W4+7RXyFL259tq++arYtj+ElEBif0TyokjqQ7M0VT1porJWC51oqEp
a08wHQKYE2wqGqYeFqnd4nggfvLJIhi6R0Mlwz5ueyNtb2B6xv5mD0iM5JqY
VxKqN0SN97Q8bzMJcsASYCz09+dvc+LkXg6MPt0ABsLFVX/a7EDRZk04WNXm
IJv0nefG9JNJ0aBvaCzI8masfsFpCmaKPLXNyX2RBuW6xOe3abtuPQv28F+z
yarzneQFjG5EuD5KvzWJWC705ODQ/E+A1ggrbInJehXWPaJahtuWjfks5GDq
eQtvY/g0EFbmECvpLRCffPPN8kEcBug3+YxqX3a8kJab2tvLLFpLCfQ0YGwU
+Xxvq53/Bm6lBwKczCTDsbBoF1FvHvVvO0ofQlhpUC1PznYvvdaKUEDiJmwB
V6fGfqJ/ruAJ2CGnm2WADm33rQoPCWEDDHN98DPQbvIyU4qFav+ypbDa4I1W
qn3ey2FjXXcrle6wRjb6PBDo6vCtIspTe/aP3cPoJxxrsk7VFfburt9EzSO/
ChqTma4jpxZc7k5kAWDLb/9GvCpxDabLKB4h3NjiQvAyu0tUl+BB72G6JabG
fpkYwNzz3EMqtq79fYS0ve9HbSZTY/0sLkvxzhqg0vwX/wb/O98iNAPojsr/
YwBblxEJ89VeU9rhh/MKvCdk5L8A5qOpKpAoEl5pwLCQASett+nbElpLcadC
Dyg3SmD60qZHKN9LHNjq9DpxgpOLxAequKW/ldAuDV86Z507sqGlJN3sQxzW
rrvt6iKeOLAtyEefjyHNZRzJyMRmgyi7Nid1ZK+VU3Z+8a5t7Q3JDynz87uy
/IThejoCbaARLwvr42jb46xhapod5+CjzvE0DkKEd9dbz9of3yFFE3SuRJ2h
UJnuIwZl/1UO+jwQuc1YViSG0D/BzFEO3Kqw4KkkO0NGftc5My7QypAV8QM4
wpVO8JeisSecgEveeQza32LskjbxKv7N29FOU9VQQWvSg6URnloaenxIFGBF
pvuHudGb41ioZRGsGptV5BnRnULjBm6lRt3n7wAcaoyajzO5mxdquWy5IQlf
MFMmJ36S+CwSlYidVYQsN0uraeTf9+mYUw+i2zv2PMnuFIfEUmJKRHyLlcME
1+bqQBdsc+vXiGBi5ytUb3gyQCLXBthJUjct2/KEJ2mAbaEjpu3mdJSLCSM/
aK2R/NH2TtNHMHWkHpHC/80fz5UbBulOSaXX5gBce1GREdLy0ZFElFcVscH0
+F1N/5st3TU/KwYXPcmA53ArP/riLa8R14t1n23iD0+untdz+u+e1QmvCwg3
5HtijJ23X57iujF4Ro6GZnnV8ZlCPuKIhcEaq2zJxmJ8iLDL4L/pedcbDJZm
KhOSEDJ4uBnX75ka/sa+u9OpprPqsdSDSA7kJXsaQR2TkkWlT/6atw/jcvYA
FB6ApRnFxvOvQq4NQ2vzM6uYe4mdjlVx6Vqi8izV5RfxTnkLWV04ZRpI2DAE
UmvLflNlgaCQIbzmYw0O5sDM7aScpAtpwyEb3S1Ge3yLSWA7WDKz0bAlvnWI
aQWAzVROoYOjYXd3SC1bzedlzfdqZE8Q688VD0mQ4Dua1ox9Q63mrrXddWza
YWAa1n2+GQ/nYyxRioPkfjd+6A210zfpHMujqzK44wBQrQ4gCWjaMPpJwSV1
wxwbJcsN5V0P91f6+EApKu/4yyigYQBo8QXvLUJNuZtiFLqI4qRhZBqsICfy
VKp/m+7oBHznxQ7VGnNWP81tKM+LCpff6kkEVeqDWBjw1MNxYHean5S1xdem
x3fZa05jJyBim/4RiETgmbzHy4T5KjBlHtc38ruAfnCv9yo7ME9s2niq7cz0
btSmPrK+s9j4RFz5LoHz5cooyOciM2tMkiisaE7VjZCoX+aNC3nDKDX/hYLT
eLZJGGNqsjXyPLEUBpUI7E/q72TsAhPNGfJr5xNdnbVWRpJr0GC97utNZyxk
2pe1elmCv2dq+AyLxLhiRd+idVgFzO4ypFljMMyfoCLzfvz2AgzMCHctzbvV
3g/kot7Z9l6ogX2cL46JcVKHZ8t/YiEi0zUJtGWr+KZ0spTDQy2JA9/IBBNa
QtUj8gKUM/HLARgEzHjNAIz6g3QQVMm3jMm0Tr05RNyXi1OL5XjCYznvVJSo
q9G6gPKXz3xotrtge6WL9Mm+lkSlVjvrQIhca2qUXPGl488UY1RP6Y/1v7KY
+3DXLhJcm9nd2CXBwMqLFR9rYcsgzkBE3rtdtE7nt+aofNzB6gZrJWJFxFSH
g846ua3erNWb/xnYc3nUceoxTp7QK0di43njsJyS12CKCYGBudsdJIYhxJ8e
/1e7U6szKOLKFa1BNo/p+2vpe1OydZNe+3YYKsz1Otnht79iFcz71sdNUZgl
FNBgP9/sro33r/Re6VFjyNc3wrBnrWeSBF94PGM7FQfmt7x5dUpmAKeecCsK
mHzCiuz4CwYi/cWZbTXwsGhk3LTO9QgnM24dyJEjXdiu/b3wjhyrL65BazAw
JO1atT1ZM/Qwe7HbK8CPysY1v+QfvCBgXuFY9ydtK7GySnTuR8ksYjGV4G2R
Fyj/CMliCiJqXg8+MFjg1o0mOrkIWcAvgGVSIHGenzCIfurC7zpEIC+w1cYX
PKfhHhAhFUlYKY4+kp9PQbxk7DLJceg0Ob6135iY96w+kaLKSYFu++7aaxyk
cKL62+YLh7Aaz0USopWdWHfL+Ay1sPA5OgviW0NUy30Ojaz9u8O6ILAHwgyG
DP+7M0+XSn0AmFaHdiUZGm4CNQqNGLHmSe4SnqvIWWLa33vMmy7DUkQ1tD5Y
Ri7OqRbV3/6xWfg5ashcCPVGPp97BgYldYVGMgu6JjxjIuYb6Vw4vfKhU9cu
1/hL8k3gSO3cQn/YIhjNHaTywPsKQblBSxtYwbc4SbDeNftJ5agQFIWVG76o
S7xlTiT5pjndonsEhSt7EBMmZpVY8Ev7I6+AsJDuuCLmx9UdWtgTzmhasz93
DRhv1gVfeAFSyJuzertGS7tm0K1LbmWDmMH+r1UqBlrt1mLGfTNPLAVWW13L
DvZiZymehbxW3IWxSslxs7u+UnhR+FkKfLJgDgs42lFxEEKzP88y83TClN6E
T9bsrreq3AwO5jPZofTPnl0IAdJDjWP0QN04PaNhVgLNXLFbG67jpm9cxvEH
pAUtfLWGWhx8wloe2ndwQ4Q+YAo8zF6Fe487vTYFTexaMvI8Qbwb4eM3QMqt
On3BuV/hJHE85CyVQLquxu7VwlqN6d0IRfznKwO7yt4LyMF8a/08joj4ebwg
r1XkTSaLCyJ+iFyd0rZq4ETXixOo8X34CdOPTnZHG8s8kEoi5JBTAdX7JbOs
hj22Xi2Ud008FIrwjtoSaz5RTydgGQuTSMOROl20rEdFSOw95WqAC94DnRCy
6x+9LXx+IAvnpYQiGLoGWXuw0ZUDXnNP/bHokNqBH2o1XdQ4NrlakujL8zts
wK8ztvoON33B1TAjU4tXPyjfHe5Nt64/GdXxdB1jXVdsX1P4Z7HkHcfYZJdg
JHTAt72EWmP5tb6h+0dhQ7GlMGTZ9rTVIgPIx4dVR2i4ZzZPBVbCh4xL7c8+
9Jef/M43B5Yw9JYf7JLG9Rk/2WQuUIPQNNO9YyDz51ERy0WNIkqkjRyHQ9oE
bvoaDFOPABwwzHWvX7Pfi12NvW+jOjrzDEwRwNnq019piFw1k3GDreoqhuUX
xiRULOC21HRmIXcbVfwmdg/WjH+TDFOgQDQD5vEmSdqzvU2xjOmvxAqRu3tl
oVDZTw766CfsBZG+aG8+KQXabeazH3xMZ4RRjvT9VEAcVmOcnqUlJ57KpfDY
fdk6AVu4HGHGZwcmP/PTsV5iYEXI/5bGK9ZvhVzb31G/SiJ/i4rRPSRx1Q+x
tCXL+ZUxwxGTVzGk8tkFTShH2F3vr7Q0y7hWtY02Qno6ZdSkLOWtnQv88uVx
Qc/0MAJfzv6yr6mCNxpwY1H2bAMX1B8pQNsqv+IBS/m+dyCzgV7kbHX99Hkk
v5LcVoTCjNV3mtaaYWfHOZAnWTyK6f+HpInhmYn6vkdAxzZCIshOftZOnIdr
J7rn1X0rz9WHKYWoUqYJRRbl4uTUR/e8lEQY3TgfGj0U7oCjcj6m9ajw7Gej
SNcQHzTLP2J2esNQFZPeNnOQneN7at2TFxJNFJ0eeyQJDwzfsgJ3Gv7KxpjF
wblHA7oSTvbn5M09BR3+YnZgR8x3fh3u6b8hjnr4b7HKEQxyl33Mp9us3CtG
ztEGlKbfrWNOx8QtWtlFA0lO0SEQnAzMfVQsVP+dcPHDclgYm3b76jxEgG5U
2jGduFNisV3rUd5HLoZauU24H2mgeQVXoDA0uSX4Up2GTgrA/nCDJZfYK8/z
seWYSu0RXar5Ou+MVuoGmP+oAlRUHSxsHhGQ47q72AfL3ZsGM+5NucLq7l+A
pmecYbc1XwSHyGWxoyQnvWnq6Azz+pW+JQMnjCuHvLWdtDZcReKYPvDbxCdK
6ZXrqqzgyVz664xLw74rRLCmM1Sp05zW8D0knkLRsugIcPE776tbihXoXk1h
tou9dgUhjgXYO5xm0v7rcJxlKqOFyxKHCz3E3TV9Mvr8mzSb7ElrgZLHEYYT
TpvjBKi28Y+pbdBH5b/MTKOYf23xNv3yq30EdcCAzsfhZE5uAux2Fa73efgR
lrhdYoEUg960eCFNrKeeyHaqRusS4XPohK2OgzsWfTgMkyuJohCnOWDwOTJT
7M46ut6JvRjunhtIhGOAAGF+xRXV78E2dNcmpjFC0Q88+WTzlBGmJl/KfBOf
xey+owKylanS3qMOFZ+DurVfqA0THl0kJioPL6dpg+9zYVVyRG4w4C8oIeOm
awaoFp+foOPPSY7wGITexHUCIsyz45lOHBCSIWSBUEeF8+ypNfe7WPPHVzTD
05iUKzFooyU/bqNz8UPkvmqv1Dp1ndkcm1rpBvagg4xMJQELFOAktUGol6Mw
QKMeGt+bPzLkWLNylfxOaxeL+SHCfkd4nRfi0PJau7rzygiOWqd07nUInvFS
uA3rCdDXFyGQ84amgR6ZGwD/r/84LRM8G8h6ZniZutb9WblivSW4emDXoRIm
LjOHSfCuQJzDU18Lb4d/fwWwUovTOBo0iFMGlEANrttBZPti5SOH26JoSwN2
dQVqpS8J80H5XzQfMxSi+0M7bFkwN4a67TSPsyqm7GkszNyWqd0xE+5RZtQd
qr0ug4lbeW8v9QSQj5HoMiS9QEJyiQLzhyJo+06JfQV+23i5z0yVg0KpkZc7
47KCAVpeXIhD6cVRut1NjdGew65s9eZz5SNY+C3tETfdPrbiqB2LQ7pEkyUK
yExy+UJlwrSkc5LZx2ezj2MgGa2WT2oCK9l334sB8D566ezA96MNkODZvwGs
hWKvH08Iu9qKJls7R6vT0AVUOtq66L0Qzn5zUL6BAxliI82RG3lSFf/nXdcc
kOOcZb4ELtfChoNyhxcEgGeDmCFmBvHupx94ixPtWmAADItvGDeB7d+r6stk
sYXnV9UxlyToynehHZXoINrNJrvkuYHTXKObwm5PV6uxsTGdYt0ZchSz40VT
+vi0Z5p4lF2Zk8gtbCowPokjgeXzhKrFc8f7ko850EVuG1zyrK2pVCe4O9M7
CsPh4TmPioWgtoJkUGFUuCx8L8EtN6zDTOlgsmQuOWPRWGp1DXUD1sfAavUG
lNydAygC3j7Uva1pgo1azsCMIDb+X8yebbCJ8lu7VqFsV/KOGRLtDrBvh9JT
FeFBt9XBxAVzrvuXzwoXb0BEaZ8aT/UeaqFMQa/ZLTx4rM9nsaK5zdrHx9zD
bx918VYTtFN1+OKZIuJBqKIoP77q23ojP0A+V8+MAyYdCOtduBiN7h6mMl3Z
GkXzjjmXujelQFroB1a4Cn5qQkuwebA87c9Ne18MXM2MeAyf9uVuXhhmiM+G
8dRjrd960XKpfrMaOqBJAu3x87PAlinw0+BEiF+BNG46cdyd56C7uecuUKwq
r4iulM3w2Kpcg005M71bUFC5mQzDh0LTSrDC9o3v/2Pnk6qUtjHc/BGc2/YS
hDUmrY2DJhlmkfvT1KNtl8p82Eez3xs8WuHF8gJzOEH9ncn8PulxmxbNalHv
IpjDagws3CYB9+v5O5kpCsAjwDMSIv4Va4u/K+jy3ARoV8xCVg7pUiHS/BHm
9myIZrPyoNkDHn6RylYYigHSfepOI+mNO1fpvQz4vWxZOgztQ7ec5Kh8LwGP
1Ay9r0nHKkVo6mer0ivK/pdAdl5kH2kzdD82kVaBQAxv8xC+htlhQVrUqvcU
uR5yk5egc+RznYtr7+QQFFf1j8PhBXevpnW3+v3L+z8lVMDSYlGPhtPNiDaB
sdthppumPLPMMiNg2wwQalkeD548YXaDPLuCgRKADL50Ww2x1rhhG5q5BLx7
pSPAZWYNF+7mw6ZSGyqMLf9b6uuVPbfaLyRzQZBPI1wyeZUcIvp/BK6gcw3n
90IUz6uRe3oYou8QVoRq+CVado/8W0ldBtjQl70eW+I9z4MFnw+BwZvKJwtg
XEO4UHdbmR4RWd/KaJ2R9/uxWj4C56zIMXbprqaMtmr/mytvf+atQrai+CjE
BoZY2VsE8OZrRXYnV1Gxytqj8RkvXzdVVE29E24ip5nJFlmFW5U2qOyMGZUg
02CcLPZgwt3TI4BbrdNTzjryviDHFqXm1316hkUK5k6oSifsd9bM0QLVYTE7
PADfUW/7WfEzCqwmQ0m91LrZ0BUZC1/pbCSAS8jQokllx4hDGv+Jee5bp4ft
0mC9iJ37/PzXYoAbuAYRJqGl3kLW3hqqrTFYEA63r9QYss7+4WHeM/VR9Y5f
JdJ/BC/uufJc8d4jj4UFYLDNVQctPSwV1Cd5JVzvmRC5W5lRlctQSsUhhxfL
C7CYOxHATpk5VCKyBMqJNl5Y+rtmtADmfEipUaKstKaCzA+BYRMUmFaGBhld
9nU1Kcgkm2akOwRpQtLXGgnw3TfJkq7an58z1XDJJqOpyTVqSgwBnOSrRDFx
rdW2MduUuToJ7TvzwheqDlillk3UrMbcJLRmhRUZvY+ndzDJPKLcld8U3gp2
ZnKUu2UlZrcbf/LduQBJTrkUgRSrOSPUMIGxDzDF1NmhGcu3fpEIiPRCarpk
jxM3fBnQA9/dzDBHTrHWD5PMZ6ibMsHqA0IboVqrbCrtCHo14R9ykVtlLL7v
57LY1AKs1LbC4/ypyhDlG895piO1yg7Gok5FYDB1Y7Ij062Y1/eQSMZGOeEB
6uURyaPd2z0ckmQ63ECUW7wz1XwS5jsgqwKXG0JTILCwwIYPkLNHuvkysS+R
+1iHJdmURVXHK2sY6NYbfmYCHCoyQAzI2KI3W8hIQM5vdDc3qqsns/wEfvx1
LSx3hhF8YOfBUgSK11Plw7WoKgJYrxdZibKn98izFSK3s5vKgmbwDCRGinWi
yqaaSImHdfVFkq2GyP1y4y8xUGT9zXHDJs1wDBLnXb39RXv1mHmBT3d6pCO9
7/sFGNrR69hhJb+024F1ZjevN5AsDA/uM1DZlCZsva6rFIEZrO8K66gRk3kZ
ePQwIQ2XdCZgbHVwdbJY6AlzuKjoJrBIJeQnl+PEhAtUhZAw8Kr9me7VmFHH
ASNmtFtoBRsvvHbo2xy4YVUUdNWd/hQi+cOpCeHeUzrBv909wYvAywHjmjV+
BS3Us9EcMMn4bv/T2M2pFpVR/JSh3EKzlzpql2dyHMikONIDnXlVJZAYkgW2
AEM9HBNxNQEbOx5gDsmwc5hSWzESZtvnpgGn4HnNVmkfoa719jhUN2u5j84V
WJVlKwNUeC+Yhec3UYlvXjSnepzN0PJ4wUsTCvlxWtd09m5+iJV3HXUWDJXH
Whjr9u6oh3Kp10UtCwgityw/ArhnlKFhUU85izDWF6vBf3rnA4Vi1LAb0juv
kkzXJt0lcyfNDkKZAsB0zFVBjDmz/C6YS7ARl6ID0prHJyUWCl9exPYDh5Qp
3tOzWCPBd9i+VrRH88JimdoWHvVchMsQAvvp2OyQsKkDlkYnYyFTepRhTPOj
bNW3Xpes1T2pTLNkwXL93wUMx0Lf8pfIFYKsY2YTH/wncL4JckaqoRyfVG/M
fbhJI4RTu2Qlt5eZubMgI4O1ljNli6q+wDJNmMfX7wBPR1Rpaekf1hyaJaEM
IZvdKtJa7om5usiwS4Qhi6Sp+omnT9eChdUr2/G7i4x7T7iTrv6bPAr+niRg
CLYsZ+om8EN49aJznR5XW1S1A4jdIUnQUjiTeLJ+WWOOuzAfiUeqb83H7i/6
Fqmz5V4nvV2yRDbYhza3eXgzz+dlBRECTnhNrlphp4B05D0BYhBA2rCD2Qib
xOEnBbDSxvrVUefIDj49hiCmU+wsNTP4lYv0emIPMoBooHPgXygUiG+NVfsj
GR4NTYQM5RM66YAUoqstyhzw+kzqwjdsp3fn1zIWLZq0k8LDBST5LdbQpxob
DKrXtK479Q8d9Wrdrq8yriYlhtoq6JvN6l4ZflGlc9zs6VbaJ69Es00g12o5
WYTlT2m+2D2wYY8CJr9GVirX4xLyE4Qv1nc0Romy5rpXXwe5Dtqm/iXssISj
5S+ihn0gwkZi27fAWezeEQj51ydJyna1gp2MaKQEqMkK6UCln/eXR/xUke0z
PN+rCk08xOs4RDSyJ2t1S2ljHlFsbUF6+gkH0+v3JtAOy4YiTFSfwrYqi+LW
BPErXlduld2oK9OD57pivS89FNEv8b8/x5eGLAaH8V2oVFB0BV8vpVAq0f8V
JQbcup8S5w7AlbUAiV4D46GouUWxHOW9MUowJqvaonATqHhXPrDWd+YTRJxY
v85AsfVDZ6TOjW8ISRjyxnvPehDkbOIOPZzjbFtsC7Ew0JhGYsvPCFSyQEhh
d2yMlGSUXnwsEPOF6w8tIGf3busPpmfpxhGi3t2m42VpCZoyTA5jm49YvZjM
o1yChyyMmfZPNH5VeJ8jjLlzLqJ4s1wGdM773c8I3xjBSRR3sSVvO86aXIeB
an0Ro/Zsqh8TWiRPUAg8t9o2FvwVvF9F3zR7ISdVSg2k+3A/oekrdM7fGZf+
oU3rUC95zSdL5ZMNsu7MmbbAlg6cH8iG7/b/G8iSc+VtrNszp8ECS1/Eebzo
/9AGUmSUfZ8hLEUcc4lc3uNFW6I0GdHA5cXHxBNy/3WnRH1cg4GNDt05AQx9
p5oUhgYDbq8kWvdkRFxfkOEoSi9tPEVPk+TV7Uh6zfYT9bIoHGuInPoV7PHY
ObaIN/tk47ClUeHW1cNug2glY/VjEkgqSgThOcn7USIgUHnzcKRaCY8+KUUe
gGs5fd58iWAPFMceCLBpK9H4mn44chWj1c0G/cb9/Tp7NSXxUuxEMwvfuEtm
bryN40pMoI7gQSE+gPCSkIEOoveQ/TDfJern+3ca0LN1NgRiHjWQcCzTAGMF
P71fnW8k8Ho/B6rUwWoNC65JrDPFHDdYaA2zX+dteFAPtYiZPjj50SiAajO5
r3uOhE33gfHPVsG6gD6RTRHSgor3iTRflptEbNbGxTicyGloK634FPwMPW8s
W1qkEuIPItOGG9qGjoEC9cH0QVUO3KHKEdYc1CkEdIa3UnAno9pU2mC5Z3XZ
PCj6m9kq2kQljII+9yFjIePvlQnQVgaFxe3rSRQINfS8yJg7DqzDlxYWPD7+
OBjmLORtZuxjHZ72/weish7M+s2RG5arD38cWpOdNpC1LV++T2XGKS6NFIyG
Pu+mCoYNL82dottimwx3J49HeETBOdgcxSgU9f9yknKGPtQlvfVo+zxTw765
jik4t/IC1c9lFcGIsmyB92FxYiYT0sdQcHu8cGngV06eWBSEyfzhp2EUUKrc
MoxVcIcNzyC+vdBkUwmPoxSQqtAJlN/5rnRCCMCjB3s/NIC7T2Kmwibkg/kb
Cdasp0wWzSUywo9OVM9b+s+DIaLXn+J2TqI94dl31FefRcgg/2pSXwrghTK7
2AdvgQwDjiEy4zhVZodvPjsNZJJyuYTtKB/m8Nzk+xnsJcwm0KvKX1KnCDCs
w4uhChxZyyj4leDFQA1EGX8fWpo5I0Jq2v2zJJjNrYjv2d1vioAYvAjpvjdA
6xxh/tQ6bG3OdPCI0UTCjimCIJOWznwrJ72lXecnIbCDOninHCdGLvyj7U4K
yAjYF6yOf+qb2zg1vi8uAPho1bCCkdPYHBLPVfhdCyxglvsRI42hqTEJSlFb
viDIOg2z+1oDN+fK8WW6+r4LuGieGmzK6IXN3xrg8i0eH3Nd51juSeZSz0Mi
TZ/18/95QhZxI34GRojpyaaCqCkyD9z4wV5N/egME1FtvLDcZQ1JczN7ZRy/
MazRXZHX5Ad3BM2bUJWFpHcVG1IzdAiVWZNusuuPZGW9xTr2tsXA/9YjwAph
YiHDVlnME0mDFdTazwTtcpMblOdyONGi2sHtqA/JMlqQsyIanoR5bIqC2nUW
Ub3rM8HKvQKuDClMFA6+95zBfLHqAeVwIEFxoNNJI9RfELFl9YSL0saZQ09I
IWSHP4S6+j4wVe3N813sOFJwXX6s2O8gfyiFEapPKSSFqKsVRXnCP9r2D5+2
fyMsQncd0QWY0PrbPdoVYFIq+je4IVYmrfeSVV7c6d7t8d6FUuxhdK+IznsL
JLOBYNZxDyTNhOexjH8H+Fyy+Qx/nPXfVgJvqQ+h6w1rwERY+Eubjcep0xUW
X0fKIu1UO51xHB7ODycAxRK7JEyCxAtW3wWwcF2O0zS1XlpiPrOVW1LiB1kj
TTrtZZDMdvqr9ZXH/dmiLFqlgVYDKnMcA8h2+vqNfiOw+V4qJ0TWyY/O/dDY
gh7C+Hz82ddGaEPfv4V1uXSkab4HHl6CNpqeUaaubjDh789f/xBBej+b6ivj
yxDDVeyFnjipqlf3WhMVJEfaxDIqZmNRIzmwL5AtTZmp3H/hNac8Qr6jng6T
8byf0OlaBX6KXAQxmX9poMy49UEsMNUJG4GwMlfhWoJB390ggnCPPozq2tyA
mcGLlT3iVNv+Q/tenwO550xbFAlzPbaZGiVWUzB/++hEcIjc+Sy+gs6eU4JB
we7nhjqvCl4KQpQkM94vOeC3eWnmRiHghM0Aynv5txhJm9CcOEQ1D5P5TLH3
loM4ACs9PUIHTa4Ozm/LLXWD6XNMU2q2ewRN+YgiARASe0H/8mOevgGkwCwo
hh+bFrSxAZsfVmC9Hrkxkj66TA0gsFN1wbCIdygseeLyZ/Ni5lHg5uO1My0x
kQ9cTYvXgMGzp50R4YcTvbCcucWTk5doBcloWllqqEDnQ3qOTDoC7dg2u7Gb
3LmkwVinCu9nM+yTtuSUQaGqcawRk9vculdtk5eAiiB2tmEUhyl4v83DHNyY
c010VlLtNXCm8xS9B3F7YvP2lsfXn54HfVwQJkDhxsnnp4bhyt5ifTEKz648
EvpgEcoym1i/07QXbjSaPU9oeUzPMRC88i2gEEPmjWjxYZQaCyQN88zpeQ3F
uhSY8S0pO0ZOGbLXMR27iPmIkpOMc/6I5Ybrxdp6kIKuRDG21Mz4cumtC+8q
qnYlMVHvs0z8l66Bvlul4XD791DiiOZJdTXUZu4+ANAvzTas3UrhEIuUMPbQ
mFHX2tdlnKHdNMj8fJKDhcfGXE6q1v7ZbC5tskDhwDjOmGWmyuxTnDemelbw
ZdnJTCMn87evWTUNKw58f9drYpTk/vLvObSeqKuK+k0PGw9uLMCX8bNLpVzv
bqqWkGVJXrQdrxyt6vfZUl+d2VdVF3YHvyyVPm4jwxDv8D/wQWQOD43pE9QX
j+E+HUchbABXoHwFis6Fwm4twkv1vraJp9HcZu3lT7msp/vmbq/GM4b2uyEX
pg5FCcMiSzYs2Dh8O2Q7ijdKTRGG4c4Yj33eqUSTs4LrvLC1/l5itfZyjLW/
H+ZB4v5DGXElAKwNOmYJ5Sodtqq8wCTLcdocUm+zSTfFTN8pRejfQ8Ij8GYi
gjYzqwTe8/SD70puFoNq7bxDE3VidLjbH8ycIJgRiJK1SUneUTrgLub/KGiH
M6DylEZJXALeaBU+gQkBSJkbqZdpvSlJI+WfQzlX4a5KexnC3bXqk7J1Dvzk
Hup4e5maHcIDy2wZP5V6sQOazvT5ANZxv6LYB3hl8DuPCtd8dCJrlkoaVTyd
w0i7VKmtmx3cuA2FwJBi2Ute+h216uoMSuHpRFgKw9WdpZRLfXWpTmVQPnFD
r9Z24h9ECn0VvMbj6+M98Ho7ZlR0pkZCLWLPqOtGUDZ8rFKqjCRhKDj+kL5y
C+FaNKOECDXWOyIx/djWWrnFFeVpuXz8yX3vG7D8HhLjaS6z+dEgm4Olu1ZC
wJEcE5lH6obC6hw+myoyryYTAtbxm+zVI1sECYIr4+xs9OJsPrliJ6ZcOdFh
T5IIa+vQoidm38uOkBAGtf9rKsUIH/ObYjZdU+v0WM4UYIvdAIxbkPdpB8uw
dkiTvSt58oYfAcKjWN4rGyjUm447BlruFzmOSaBYCIEULAClJhtwishWXBwb
aJZE8DaxhgvjzoaLgyf6HhBA6qNxxj9rMvmnJ2U+JvYmfLAFdUKbAt+0tLCH
lBw8Xo+fQe4+4ktC40kgazeqm4lhtT7qfzVAqwrAKJq8ubXFe/lC1oexknGH
EirGD6rOg5rhkujVplqRfCpYBQLC8GP+up/Uojw+vZGCizqusb5MNRb26PcX
4Th5TL+SfJNlsDMdmllUcwU+mvdqN6NSvqWPnAVLgNHoV2oPB8MJnSF4j3Gt
fAlw0ID7n3CeM1WBseUJHlCYmR4O8JsU80nqq6G/XKCU+CjxCuTiAuuMkWQq
6GU5ejfALpmruXtvtPODZBHMD83MwSe+7B4UanmAgLBerf9kju+yrkCcgtvC
g1mE+wcvb3VJycWm9x0F7MW81goMhoNPd1+0wuJqRcLuiXE98AFjAfR6l+I8
eO2Cvy1VmZE6VMVf40otrDWarJpHlWAR2FVV8L8TFu4tb+vztqC1Wb08c/n6
GPRx6bCXXfPD+Z8Py8ZFBYOIOEbwX6vIiDWqcNZg2cjH57q6oIz/kUkp5aQb
cY//Ln4IbxGO4LD5PCyAzepX1vD/SXQWn45r2nBPUK6H1G1rMhFgs9JXTwzu
calB+7mNMqMobqErXGRoQjzYxk374YhhFUhsTldtC8rbbfTcY4eT6uelrbHW
MT+yiJkhPO2LVhFv0piXrmKIQRADdMEcnVdLe+frcU1nBaL7Wfj8TnrPwhn7
EyVZGD/xLlsyAVM2CIClSZyGytgy6vc9VmRNfPx1PG8P3cXfZzGGKPObK+Hc
eAiU2HAS7yCU8Mgx94CKYLZ9h2uZy+AWY8pVqb1NkZ7ExApsu9QPFASr4WKs
U2dE1HLxRjMjFraF54LEcyB5TjXPIuYOhWMvKQTKw4q6MMuKuMGG1BtvE5Lo
k/3nxKKqxJes9Z1vfEzZnEx684LUojwtXelQbYO0V39Yso5Ln4BAEDSzt+kC
wEuuDNSa+sme46Bih75MJ5+x919+tfJaZphi3MH3gRFi882tNZivv77HXbmR
plFT5Of3PPsjswyQJQVzo49RXsmLAGtiSH13MW3B6Fj8ctZdfMMrWIVzfUk/
Y29fGdlS7rb1Vm8frgj1EL0ksdyxv01I6z52C3l+0opt+UgrrHoFu8X9oJZ0
lmABbYL2tkbng1VhC4Whvlw9a/h+YWP3s9HOKQgj3L1zSU+BaiuqtNAPQO9E
NPlofR7n+T7/39r8cQOV+3AE54aeaWnvETyifiYY3DD8VrlHn2fnfqWWSI58
GRPCCzh6iILn9+uk4zRiodSwAlwXh4EN6zusg4dHsGsvW7Djzu7VmgvjRvFx
xGLIuXco2lCNGxT34oD0N2mpKNyslBItqDPzks8Jv8OxAPjVeokj9aPvCoLC
GvPIh3pKruwvRaNNgV3Fj4VnY5dM2KloGM88TNZBSOBOpmInjYPNjPPLOaTY
QWAr4ZAHBudD3DJqvSewmL/dwwTL29lrr5rRr4U5343zwOvoWOyNfpV0woVu
zry3opm27WUVBGfHx5svIYdqHvtFfmKQpXekvHoHm9P4Xf1IgC2lDZwml9Gz
W0xSB4o+G2+nU9jZe38wRALuMfbpbypm//hxIUoczwpLIvo1HhwtRk60rmJN
JiO9uDKBmgDF1F7/uFY8Ds1lXPuCXI++QcyKn9Y17AfoEVyveVGsNmSRNJ2C
ZREraU1I/ddci8bMHnUJ871ZqNK90Gq0gY1/kQrOyM/k/k+/J5nsJKNnTAiv
LkkstsPNYDFidnlo5JfsVdfiTV/xhM49OfjLrIU9U6cQuDWN96O1VfmMGcCd
8h0b2WYflGwNVBj36Awxeryo5PVFYUb16XX4HLaUpMq9bUACYvxx8b4D3q98
fqEpY0+SPs2QqENjrfl23pEJv/2Q2ZPtokL27kP3PnAJWLKERWyfUL4nHY7x
j2lFwsYmvr5JNEGwyGSzWxUf0JBcRf2Lql3mxUItGuh9Ue5CKJ50QgDg0Wxh
6nWoEGHr1DNQq3nMtmMVRXs+5yQ8Hy55ga82i2P4KkoXlATNm3n2EV8/liIx
/i9cfRxjzJgTLyJGH4TmEOXoQwaasLf4ALS+rGIpmA7q5Hn+1ABfx1HvHOr6
vZXMrtyn3eFVinIDaW6BPs4LVFilvTtTkamn7he7DOKSkl8scNa3xUWteIuL
weMjVrl4mALTTN/SlYYpn/9LNER/qe5BjSp3MDJcpRk0dNta5PETxpqk12iN
Veigie3EqR1D/ofNR+l2+rhrYRTWhOOp/JAlqqBsu63afRyOUg+eO0QEBGng
+e2vLVq5KOEpFezR97ZtvMTt8ySVvIA29BAkcq6Hb9U49wZUgN73ucIaTECO
i3ucFiLnz2oV5vnZU5F7uh06bqfEBZcEdIyI8xap6Vu2NwawWpJIqlfvbT7f
L7XZjIrLOcaFWnJ9a9uKUthIhMMCT2E5Rle0CCUF/i/OBhIPbsxj0A3iOV9N
gv2bgFnhLN0qONdzawc6UhrtYPwpPqule0GQzzySWBY+M+sW3XhAJPBVGT2c
7hHHJt5p4ZJKTsHXvFzxZHNwSUjNsAiZOLGvtj2+ebcKhOhB3b9zdj+mFf/+
X5gU43NTARQciUOHmzZuWXSPgYymTF4elXMLIqQ8BOFKBnwjXPCvS7Sg3BtL
3MATlVyc3PbmIgsWVKvBUO47MBwRNnoWKBaSmmFe6Uz+sDC4+XgnayUxkCYb
dOHytVvjIUG6r01AhXRXeqhjQ0FpY+1dWxW7Ybg4UREWTO4reUxUzHfZs9Zc
KO6nRJpJXmIF6JvsKLAEUIMNod39dEHTlas1jxjdk8YR/tWBCJeFPksvjuGW
w2TRlEUnBvTviXxyRd0KFnfWtHvHHlQ6sdGeAfTnLb8nWB3+LyoyN2xbUgXN
yJeG+OKgWGvHAF1MtbdYzz/kGI+/Mtkan5a2XTTfgalR31QG4pFZGq0sfd/l
ryliJQXQGrFJaqAgqyYPXnISCHr6PZoXr9u5q1P3pFYeA4DOXS4qawq+sLMU
94nTa7PoAyyMxk/Q8tUZbccwAzBbRyvKBRnM2iU7xFNQhXDl9N44ZILpReK7
t7fOwPmN1CjqpiLQUKkHMSV9WSyO7X5PfQw1Zhodwbh1JaEV9lbSRMKzzgi2
36nmUxSGh3CBHCTj6P2bAwTE2jwH0p0fn2OdUksS/xn/3trx1kwCCId2caMl
CI1p5GTMosZmzskcKGOr9gVZgTVZEKOoIz9j4l68yJdHYAfptW/G6hKioezw
fne27lcZM2Ivbe5oYiEFJAzEXfnQJuzi7q+zSiFsEW5SNV72ZBLH7kKfyCG0
pdhQo+dd4wrl5tZDv4C80BTsgl2P/miCwpC7w+bvw3wzSQ3l+B9c83N/NCpK
wqt81uAAiaHyVZklKT3o4G1qvrqluJiebC1yr/2P7lGhc563IccUApATgQOA
FSbpPcEm3xdvfEazAlYh0HL+Umc8+TYrPLXXm7R7FVJeoRrriSbVH7BzoVC9
prTV6mxx98QV5ORkRgJuZTjq5gtJbRlWZu3QeSk89LIfp1Qj9hFgmkFK+r+c
aZY9SVdC5eEIwdJ+I7DIEwi21eNYJ3KrZxmBXE6V7yEhsnemwH0oyzJrz/Pp
5LWR2Rd2N+Gc+jmWYzXkSZqI1Izp7aqOzNYobS1LJgoAfWbiA8Resxj0LJtj
G5OVdyi6mEis3jQUJYJVyX08+NFkgabhnXLNYjE7Z5AfFkve8eZSXUobm3Z9
F620LiTJOaqdRnbYivSSXK9yQ6k/f7s75mKrVKxEdT+OqYL5sLRxfcQa/P4E
ub/3tHHxvNYzXrF5h6xBCUMObdf9fi6ZhOUuZPUeuD7pFMeNEvHIc73uQX81
pO5uABTdXwJMyn3S0cN6QHlS633y5I+6Li2fhICcUTDwXCy0F4I8un13nPnz
sMjeg/wuzWeTDSTH6dasqoSK/BYljVk6bCWfzU4RWExaR/H9kySOrDcPFUYH
klzu4ZQW0sp9bDvzpkAlpJ5JVZ9wKRMV/w/FanItwDTg7eXCeYllb58uY1Jq
I7eGyY8Q3T0zQY8CR+27jgrnzaM8H8Nv8v4WU97PQBRo2/vaUgiIrciEc3to
5nZeTcO9H7QP2Euw15HxOG3vLt3eXc20aalan3gRX+wjW0Et7xl1XCsuVq2L
t2MKVAt6XPYrBmKTVuD1cMAj8cka0MnWsGOn/TQbqYptMwlmqRjUnN4Dg26d
NrGsP9oTWq+phxHGdsSVZhJoUIIsVuh+6ovmA4Zk26aEfgMY4Ua/f9zNrxdk
03SbnkFW16+RTlAKaWimMgRjrWnUnmcQ41lturCtcFcxr3fx/dq9/DSP96fe
VHM+BBF/Ol6rmhav3yyz25/HY04zzXj01MhwEXIdqUGgz3qg3IGcdnq/psh5
ahh6kZkkAeomMiFzgSTJGRaOKHSStcOKZAC7hXuuOK2O0dWdq0QgfOnMfeYc
8wcZSC3p6tfsKKvbh7J3tYvO6U1JWV0DslycURa6cfZWjPJAB1u9JBUwvtw7
tKYOCe8p4g6PEFowgeSplC204BRe+XVCTHJMqpLVd3ZFugdieWFl9FWO8mw3
DISF2ayqKHL3YsvyOYOdfwY26iNBqltItkGoo1zRQsDUqm87XQQiikhhKGD9
+19II+lLCU3PN9bXKj+MukuyjvJCTKU8M2jlR7Uuf5jqzH/s3gEOCrjWOEHH
nKS4g9YMx3aniFJvNFT5wQYGTIO2bQKJ2u+alGsrAQ5AIdBy+IS0GOxfdDMt
Ciwu1AORNc0fTJw+d5HViyfRCd0zLe6A74/Hxg+/hfLiVpUuIB09DaQRQFS4
HBGM5uL43gsIC8yU3zRqs8RnQuuA1tZ6aRCG0ckR+cdaso3FH8vjTi8QCU++
WtrjrEajJgrMe3V8OYGFfHSabt4ey3OiUbU0Wm+rUk0srBF4ReXz6Sb0MUrC
EBPO+/cmC29QB4fM70J629NfKAJj/H49VxA4cJIffslRY4SA8xb05V71t/VT
+Tu8A+gfTg/P91Kejk7qCs1/cMFuYd8uspxLSJYBRX/oI7yanz7m+vW9ZwyS
qrgl6bPsfKfH0XJXLTjUwuLKfWlcMh6cjZBuSaRjnSpmvqhQfq+xbrR8MFRF
E264YxhYdTFnxnaKXL+TAfnBVnfk3keBDPj3tAJWnNX6tSCiqLwAXO8F/OUp
dFUjk+myoLjjOi91W23cQLHBrTpUeEeM8r8E+L0C45G98pRkYm8ESdDX8JJh
fo4Igk3q6dvdJBqG2+dE22my4kqzuI0CqZW45Xi01XBfTI1n1WNKVrlUB0D2
Ge9T+5YGGAerx27lNV90dkKOv5bbPLYh8sn766glG41DOD8b3HYVdlI+4FXu
remiBJWpvIXxHpgS6JI5xBa1sKoe9ZEfj0aAKvjYSrWT9/fkqdHtAvgjmoJP
6wnlejr4lDwIBrobiYF11ZhwXUsTzvm8T+rc1iJnpAo0qSlKptPlRz7p6wXV
BhtfmEqeWBkYIp4B5u0FYQwNCY+UjUGx6hEcZU3wyBaprbrzF03+oCyaP95n
uhdbzQGoz7/IBocZijII7f6qSWDmYnbVnlfC0kf4SFx1Id0vMjMUyGmOp0ma
P3vkiSwsDdvBdW1YzkI3xfUFjr1aNQbHAzLLeUYwFP+p1/UfxNYcuvedTVl5
mCd3LuCUf0hSuFYocykRF1PUauCZZBoKuzeh2c/dT8tGo8vsb0Z9K7dR8Eis
fBESSFVnD7ABFvR32DJlbo7HvHi0BrC8+T8BxZjoYf7Kwe3sVU3voRgjxbrF
kvq4thg1pHR8s79POCGErHckGLh7NKranwlH2PK2qInEBtNvNQLMGJV2ufq1
5Uihgx+zRJvxqPjdNWfo/H7V5DCTJOXn6J+I3TQ7NqOlx4t5Uarn/UnYuSs9
nXeqgak4SYYt+4T4JGcwt0PcgJOk447rOu8G4vkUzefzmzheHHM9+BkC2W+t
MDSPFBfdmMU75nAFR+Xm4uCnCWNyP74cZjWLcdyauQS/l2ZR0y5WUdacrb/3
mTn6i37XSFmmybkX7xkcYW4SLYFs06LpzoVLWot/uvE5Osg5sD8EM9htIbSI
Sn6LoeuRWZrDiBVMpUPOOX3YPBQ8COr6vgJVoEtg0cfGI4PLFMi8UCwlCLMi
DnXHNDl+xqxj3NSzBFtpBvKLumfSKQnjYNTxa2//TcQfJgiivSIR+Expsocp
zhv3092N4svdhXr/Q991GsUBWxPxLaUyVQiu91gJb1FTIlXLoqFSpp/fdGBV
0wl8TCSdJt8hvBxuvsKGgSfz3/4bB9w7XdxKQ+rZB6zTqtj2Z5IXmHWFcKUy
C7ACstX98MErAURukaEv/UOTqdnF7/mS44o8vdcu/Zv1kMngzOlJLTAkzqjx
VNKcbZpfkTIOaVsxp67ZyWmroMHBacVz9tT1yUIps4OFv5Q2DbAHJQzXJmU0
ZpUj4luGwrj8qxDPFwKF95/8DuniJum6uJ8ki+sK7Ey34bzwxN/Np+WmJ5vo
REwYl0TBaeX4MJzzrwAA5Fp/oNKNxlab82zCF/XCWZpxG25EWlpj89nQO7kI
o3nTtkXY1ZFhexOF31+XLQr2+wPvXV4bbt1hytJnGd2gIbr0aMLcdVBkKME4
ROMfggSpGE+nR+KH5K23X2hq2Pne575dIiYqFn06Hv/9hf4EardRtkeK8QFn
6UjKd8xVfqJg58TT8Qqxx3pleCoHNRvTrQn+1bB4WT8LfON7ARaeGsVgCWgi
zplYt2LmQ3W1aRTe142WnBsKUdhjsxS/Ww337BnsGLyeSc6Lu83znr1HLCcj
EBSashuha7sGisMtX67hXwC+WND7OWShbcAFBpdps3zwpMOfkUt0ZfWO2MXV
r+0s8RuzEk5zRFBOmJN/Z9IMIvcxV8jaID8YH0oEDjlHNhchbSkbT9G930U8
M7Xlsi0bKQ+Yi1Wv0TkDvC0zgAzYbR+zSdq2yoEJ7c7W7ubCZ4ZWkqNY7qyT
WgbzKHaxGSBklZA23zyfdk4lTre2FsEQayGYq2jVCmdUVvGlY3nY1wM7HAXv
wZFRWhps08PLSQ3KI1VubQ8rekdx00wuW5A1Gl1wKyg1m5s5wUfkglBfZsd6
Firy7ygNS+xUhDEr//KeNB5pepOGRoNOt3XzBkCG9FZHGxrG41aT2nwceyRL
/+8x2z6JGR3RwKKD7+CWsH+YeoFoXjOF26BCOcKlm+xQd3U6DvWIKM3ycs4S
1Fpi0ZBxHpgCjrPsyE4Db7yBOtVUYszzzggYNawwz0m7NWIpTQK1dI1npr5t
auf5JT77Lf3HyLSLvygFBNZDKGwrS2h7jFtqIH9SjS9xJoR95cCOev8/mYaO
4vlmMIZ7ooC4gShgb0kKV4bfxHCy/I9WXMUs39zyB+yXJm/zmHfoKw7tufFn
yrHXe8gQk9zMa7X6DmvWqVLXJy3AZy+ag691d+OvIsCY9R5s17/EP62wEAV8
LoCjV1xLb2QvIqYMoD7avjrHxaFk3wyEPtKRxYJFYyaYmAGko3/nm69sk3Rm
4xQ7oOCNhxVJpW+4Bof9ggS2M2wnzWPUecUfkOBq+3JXcI1uW75qitKue+zX
NOuwpHuKW4Hu/liYhABLT91JVhkvlcmGwVniq5rphCgkf/8N2wqhi4JZVbGt
E5PdODpBBmWxSiAhPDjfB61gSbzLlPx8WdjnF8Ny35q4iHNrwmBSHq/HTnJ1
kOnYBwRPj02y0d3c4aRqFbCpmKRn/ZzEIEnc7DO5yjI0lzJUBmO/xs+ZrEBg
Xieff58AUrtytLCB5336RXyOw5nDBzptjc7evnUI0dTACz2R6aoAlYv3Z105
ppVLmxeVQQWcUFSYmIsToUuTeXbjz0ucYd8sstjJ0bYjtCF/jiOO8zXAMQGc
QnveN//9pADhPInzVtRHNtlh0Uvjl+CyBiW0a8t7vEn7o903aJHwUsHRv2DC
fdyIwCKYnipG7n/QPgIIdaT/p3Fw+kHgAHckm4rHj1WaTsIZuN5wrSJMMyAb
fILimllYREVtULWEiGOnSFmXQvCvqjsEr7/qFVUwYihNRqhD0oukdWL8Oyxw
zrN2zRNPROwMon4el9BPwipjdOV7Vn/kalq4hMWER4qNJS0XvKeRATIb3DAq
+ewBbIP6AsAiBlSyUjJ9Tn5ULqEh99Lhwd6EzUTs5wg2TRHf2vKHemSpLeBW
9cxHIQM4YdzWTmUyQ/CD43sDNqiUisfD0BpQYqNipOmMfAYvfZQGWamTCMWS
W3Z1yXeuy4wlZB+JDcFqO4KZJH+5kS+3oGBADbSNAQf2ac7TVxN/hfEyddZL
QdlLfj5CysQekkyPo6RfZTePDmNiJJcsclFn3t7ZHc6zxDeZCrAkd3N8KrZ3
3tH17s/HTdbRg93+zyz2NWvlRo5VlVQ7NkMDaTrMBWQ/iqEe3FeCw3CF8wfe
hsRsn/UJksTMuQF3YnAfCHvSrlPoFtUQE9ZpT11i39tw+Hwz2qLREWrckJs8
Gz/CHpJZ8HkLqHNGLrHoFerH1qQDsjmFwxltQwQQIeFEm6df9ygzykrAmPI2
Pwleqb3lzTxXgpGKgjjyqjWSn8sKvwQG5EtIhZwuczHZyxSHZDkmQn/IVBkv
UKlGEHLn7bX+W3RltMtc/vq4Fh9An6krn6SPeS1XJ1d0x22AMubtFiWz8Jlo
YpRINOm7mYlJx1Eyx5VK9Lf9FCgbYv1nGf/O8IQDVPvos2V8qq1Wf+6PC8R1
XmxwApSzVGM+heWMxw0YsheU8R9129aQIq6/juMDZGkoRn/XehFWmxevPxoM
ZHHvKp7y1B3WzMGVeEClevnD7QCYtTkosO+pDklafAzmxmOQj6gKM2+OVDpH
/NhXtQBLpYLVmyEndWIyYJGqPxfrk8gkRWTq4toNzfxbfhSVdxvUn83kuFY9
32jHNtpaQFn3W7o+rOCgrt2aAbFTH/ndYoSMSkzdvdUcewB0xV7RV4VI5yBF
0uUWxJNL37uweXj9uOGOKhYFQxEYvwQbG3PuLJoQGIPujP2tV1c5NQFfx63Q
/btn+bRXofiU1oNMHIoqQaWJ/ufWlqpvimV3LUl/GJz1WrvcBRn+VpfNKRPU
vOukfCpva5f8lp3tE2lfxrioP5ed7Tu2dRWt1rI9sE5eB9WRDo/zxbpLFdqz
uA5lX62//cDvHEumFq8kV4BAmzynVMaMQ/gILMAyRzQ0WbEts8NTOSXWJHJ5
0KWjd2OtdeCPQwNygzc4njQVyU21nNs8yQF6EuvTTdMI3x8o2rRDJhqlNlKD
cwhICMEb/S6m/LsKyuMv5Crq9XPzmBevN5RzEfVqC8bw/pq0feGTpGkVJ4P9
zefazpYa+PMxKoNIG5663DKUyzoaLOA9zCKFW7JNCQwr0PdjUJc808AP2U23
L48U1fhb37Ap4NF2l1IUsga+5CzsYvW0LX/vFO8UEsSuowujVVL+6624kVlk
72wdsrLNVHPpZ24ovHP45ptCeALk7WCMakTOwZwySygZMdGwhXJ/T2kwBEOC
eS0WlEkhYO1QgY9qEBoDyAIwbbN7jJGEvMtIETKuJskOiBoGZSoN1yjsnh8+
RWBIRN/ujtOAVyOYe1AAM8NLqFn4yZVN1uKRB7YYceSxlZjjfp3D2TB6cz5I
X887SVMUbSA5Fg/U3g7GfneimMA04Djufgb2GbqUAo0NrrBX2Ccdm+TpMBlB
Prphx2dtZVWuciRe6pNh8r/PUo6Yn43vTZIUG/jwuMmaF1W2pY+Ld7/hxlEw
nMiOSPYFvuavTzycPCKgNu9JSlAVSbsH8Ibt+OXpQZhvh80cHpWoHosr1XcG
iUmkDrhJ+16luLJ9PF18MlB3Vs5+gRO9PDgjUz91XtVgcgnHiiPukkOuFEtr
a4QXJ1Y8iq9dRZT4MG6DMlGlAUVpWxLhb8/VQczTkbn2VokfxgpsdxIo9Jd1
vhw8J6FcOAydci4eADpn0SBt75Ac4Ff7afEA9vianztnSLo0YTQIgllRjheb
GpSHb6o2pbyJHLBSSaR1Xyk9DfDHt2rzce2wH3yxpYZiOoQDrnHf8aZljpJm
VxEhEhE1aBVcOstODtq8RuzM4Oa3eRU834nEH2JsREZl/WgnzyG/5i6fdTIP
iIfAEqec2or3qnGflELDnhWPiddZgPSNnZ1L/MHMIejOBm60JeR9a2ZLJdeD
m9twWMbau6iSyAU+FzcXAdIsM3Vk0iiqcmU/DelrUXx+B6s54I0b0hRahkka
KXEAhXhNbw8R3Dm0LzxEhQuJniaOzU6610LvKjKVjEdkeP7XMN8CNm0eBXST
Kb7X1oeITG2LxF1/P14dYyoTK5RVS8uqh8lozhqcXi/KJxF2/gNhEXoNdqgA
adh7p3yfgFZzcLoEPDy1VXK4skXIlXHHXlyA0E9jZXwvtrwgQMyLERw+fNjG
8XiWXwk5nS3Q0EMGihf54mn/lYB6y1YZ4VUU5Lm3J/MEX3fLxAkIncQ2Jt5I
xSs0fpDAUg59AwZqf9v9DB0WTlIegh4WCujoMb0IJeveVOASvHS7PDLOZCFm
8ortW9uvEVIqLgOrfaKZ66vp/yBDzR5M/RHl050GUjrqG1dEaF1FAuE0o721
1TKZid7E5czxmVJOCAOn21cOXXqe+WPtimffuIP9WTuNxqY0JxmcxS1s4Wm9
c5FuqBFvXgcrn3HnchvHEPa+9hGZtSVlMSWMPuphYj2zuWCAVCp3CbZdySZy
qEN/HvqBMhvHn2nLJh3Ipp6TU6rDX/vN92WGSdRi7qXgNlrtar1m6/zFY2sV
ByoVCGtqyE4G2uVG/ji5cvvpmQ1SVKJ8cZBQoQzdefK3xcFDHtsyVsJS+tzG
6MCQZuogisnzG5rstp8M3uji9H4lBZBs3kbdjMbiqg3UrLm2KwVe1NuWsR7L
qcruy3pPrSlbsLiKwoJXDvGezRnhhzY5mWnd6HFO1lG8fh4h8uW33jhAF+mA
+4xn5Xv4yoGU5o5141PBVpUo37nMXx52XT/x/3OfM58oY/3xSO1Il+arSRjV
FmETeyX59Y3r+7ioafB0l3uNbYbQOZWvSKrnM+PaIdJBmOTLaumNUfkhHCgS
0yOFUvcCGmehWSWnMoAKbKBVLuV6utUyszF+8xfvXq2LeZYAx8V/4sUb/kjZ
EbCVDx+c+kwsWHuejm6MjOW9T+bbO6Vq0AvQ3zAZ+BVUzcLBCYClBvaSBhKR
cKQjZa4BbeOA36lutLdrtEdfNsXcP9OsmGlHW+Q34GMbD61skWFqe8+Uhrmc
fmP3it5rO+g8QlShaiTmUXmV6xLaVqVI9TlHeqtSynTFD71nGkMU7RYRlzNq
9N1WbqcrLnXjb+zVUpmq9DThp2hEyKXYCDgzzuFKQZJNL6EOR72Uddtfec2/
b1PbEuOAwLf+V9dP0MicE+0RjulOfJIKj9NnvG0hDf4LBy99l1o90MzGuJ3U
4O091hfcrsQ6ktQu87CTq4uGaQgqXFdexcqZ20k+PD3cs6h4byzAgh+UUPjl
zVe0BSr+/+m+pCxIGyq9kBjSI2YAOA7r8ZNXY2xefwkpTCL8vnjFmiWa/YIh
anrBf6xNbNq/H2S0FBE94EV9K50MvJO8559FLcXd1tL7unyuHFd/VMvENdWw
nk/RjZiLiTTxp6aF5V0jiEEGRzGvGCPLqdel0ZfFKbd29IdSbyJVnrWReT52
JeJwgADfRQ2ZgcRIRvEe5X5fDsvvx/DlOuiqcznTujcHssHo7R4brRUl4zgy
cfHu8v5nqhZtCNxE46/SYdr9Kch8OSxkne9J2NxQdwR6aUec8PTrBhcGcDzl
XH2GBsprDIiKKE/3Koyq3NvJRLF8aHFBxbJ8A/eDZh7iKHWOxBmJQJ67n3aQ
WUiwSN63X5NVRi7lYgSRMxrVxSUlw/KqVSccr5+HyXLgugavIfroNQp0tzMD
AQ0VIQkjIHoBFuClUr0aG1D2fePJs8NY3j2puNHPlDduy3VK9dhF+w+i/LTI
GFvUeQ2zoxhhklQQhT0aK/HtWxEoDc9Chg892ml1nxR29YgDojHeiX4jtz//
EimJppUfMuDhisg5DBij/YqoH6vB7bEe7nBkBYUebGSFeI5nmsPwnnir3RKA
DkwyDujalEY54GG5/EeHOf7esNkdaOMydm/o+AFdJ+1EGR5QGsyH0Bttogep
kZ+HCYT/3kRRO3i5vyhTZRR+P0wPeUyqn5VY7HISkGgOXVa/V9hxqRdzlA00
cp2sdq6stym6flmaGGY/EZ105RwKWMePUA4oJ1fDbOYcIPuFqg7btV+hvDjQ
ijr4NioxKtSW5BoSFtfssVL2Q/1B8Kr/ioKiswcBw1JP43KS1BbsiVSamXV8
VYm9PjKxXh9Cbs0TF/eqcH/ttoMCuU1unkqnAF5u+0CD0hQiauJO87ZAb/2m
WNIL6hjTKzinoHwsC41DZFhntK9kF2QILl9IDeM0rJHGl40/owQA19DqpT+e
+N7M2p2DnS6w2d7Maz/eejGxqZfWgySYdH8eCFduG/XCYzaB3rmKmsuxBJ9b
d/2PuyJDeHVQRdSKr7LvFNQrjaOCIaH8MRvRtF5Gk9Z+0r8S68/KhhnByBpx
AUTWy/CgWimFkXeagJRJ43FoeWymS8Qa9t2nMzwdSQ5kik/kOotuordCbQBA
q107HgVbIdM8hXqe04iUQ/e3YfGTzZ8fKTj/iC9Kmw0xNe75R+wEi8eXs25h
0NdfqurG9OaQzcDLxkGPJykV/q69HwdtfRq0BOML4BRC15YZ4lYOcbhsETWf
B5fZhlVQo0Jp7KcfeDY1Y5lNsFxkRHCZ+GmI73kZpt4PaRiAPli97uWThkxE
GhIX2pEm8hI3ohNhR5cl4YwFYdwb0utuFtXLm46ikaK5rVT74EeGjTcp0zIh
KixcfbU6hVBvtcd8/50ojulR4IexazqL4gJbNVxKuDovoD3qYNQdPtHQFJbK
J8MqhalDj0eWt8OZdZavZx9SwwHudFCgiAif5Y2d4++uMwxHpazt18hM1InH
7r5Ppjo6b3PK3nmi3zncXOd+/dY9PoUL3UP56VNmpWnMUJYToDDm0/JMqQ/Y
1DuEXVayS5kO4D42NEgJsNr+5Ofs0lS45RPmp2U2Dmy8HOXu34uOTpbfxWq2
6zC/mbbnzJp5d43qw5uo6J3iDdLvQa7vhDuGBFGQF48jq18E/4kaK/NPNLCW
0iGVdifLurQwAkyl3JE6kqoy+uZF43csfzJH6iwWArh95C7RF4RNzkhKex00
zf5cNMyOFcqc0XBHA6vGugEJIvw/ALvpyHF+zawvaV+kapMiLjiGNoPkIi/r
KIghiEnFaKLz5OlwQnVCXuKO/vjzXLLFIfaArLv94UBJO406wKB7+2IkxsZA
/NtU9F1AXtxZPWzLwmuxAAtzhky0JSp+v3PX8B64iZY9SRturCMsOP54KFfl
cyckcuRbI2/D1eP1EtdLavRQehdZNwHJciioSmEeHQh6Rb9Kw2tDOXVgxcVh
U/NhfOt87KAxGsgPwD6LCJurOPShY3yXnXNwAaHuJBsg/106yXU5rP5ozF3s
64XHHMFSo2RScnPPPi0pCBXIUnupWnydJ4WfoL8cc3rPaSfoYG9t0G5pvNwg
J5OW2uRvC111di1o+1NV0M0Y5GvfzjuSD3fFlkrNB44h25xQIi8ocAhnvGGB
y/QyC7dI34XLABy0pUv5ra3nm7X1tOwWWec+zT6mCdo+4iw+iszORfNAe6jz
LaSM8acDzL7IdysEDUWVSokVmp6Jw3loonu70DCQF2+Fwe6wX07rz3f34PQD
9asKZCb9bl7CRbwRJiPGsGuIxKpt9ESmkIo27u1RTIdYWsZXYCTqwtnkC5d9
wPZZpVzNkF6/urhynyIuoTxdrBSeBIKlznR7dJUN28dUtQGEG1Bzi57Tl11T
VoHofWFhTFe9nCu47atN8TpR6X2SfOMyoRgTXcdGsHgv5CJTqMrwrxgaDr/f
TULv0jYi9KsSo2I4o1nVHCHwzJxDd5dqL9BBmEvWPBuaqk4399It7p4aj8lG
Lgt8yZ2hhglP3sXCCqvAw66tA8BVt02wt/rhaeugqtJH1DCkuAhunq3C2Xrf
a4Gmugj5GiJlCsvTC3dQSnBq/YWQOx3RKOosuITasOLqHxLaus9qLMLAOYyl
FAD5oHO/MadvzreVM94fWp/aG1zYhTWTdnLVWZHKbqJDo4Zh1UHDtS1ZhB/Z
mz3PLHuH6B6MfTfrkD9njmk/FXYzRtGaEGYgMb8WGQ8Wn9Yk29UaIlHP5bwt
5//5lze8NTUsUNerXpI1FoD3XDwwvgDgaiVkjjSYDh/YnLFSbQwOYt64Lo1F
RbPklX110rpfzZJ+mjLwh4MvztD8C4kW/km07qRsRQHv0S9HoRKea6zct5Rx
C+COCtK+oQcFXcpSKFaOSYVm1MLel553L88YUNXVJlP0vObYZUdvQiejperI
MBtg4gVhigeBDWkkG359hdfTzkrEk8upMvPWlV4vL3WfMd1Qcy7GnbZSk45t
yBW19AC1OEm11VTOxt5ZSNO2Z9PvE7Eq9z5klJe+k6bDWqlI65K/gNYnR6Ga
ODbVEZ5y+sjFLFgu3UhCtUy0RHYYWChc0Thm9PzqhUxWgH5xFYBtdkyAV2LG
V2egLVUVcDxKQSglC3biCEToSEpt9D4cqvKRwUtb4K4roeKhMbO1mXyGcS9y
CD+nYTadKZNYBfKTe2xLtgKYiBlIw2jPzfsDufBA2/HMyfme8crfy73y58ls
5iX82PBHWiA/py4MnwKntqmF0dirchcdlg9A58BbpCu02+EdEMwRr5OYt0Rv
NV/9HotGhM95Df3WFpZ9fMBQXsQvTBdsP11wg41DYbpbjHIRzXxRgynEKidO
ZdZmBsp7qf9WN0a5OiM1DDODgKM/gNr+ZTRPSiMAEiPR8fBybLpwGbcASJP+
ZNaW9j+e3ukfuWZ/Oxo3Gy/I4L6T/O/XY4oZ486aFl7UaIL5jRC1sLDCLLI3
sgG846EkDeWy6R8a7ozcufq3CBaRgC7SPoyY1DWhZqUWMOweP7vJdOebi0rh
YUbO4nmSNYeGPKSDYgQl/flu3yNSDUlbACyAdoPPvX7/Y/geYuOI95p5Sybr
NBO50FVckni6EYU4jfZ6XO95J+/HKScLbI/u1Tx8zPEJY7mj4MYA93jXToQc
E60gn0KHNWbF+kSlX8yxJJBnneHyvDpzVWJ+hmgVKp65lPndYuXMRMGQfAAt
RDuNMxUP5dFwhX+qhxejazrh2jbSCck5MViBi8ajABH+RLO2bkTyoU0S/1b9
mofe+V73WPUCb7aLTmydncf6DUzhqS1vLE2Z9x6/vM07HUnmrKBUGnHq1z3I
YSn5ZiaaEz6Iju+5ZTpAIFuQRIRsN0eVw214rgkM/3ygKG6dQXmzRqDsGKfb
O53CmkLWUmGIO0u+szUxBGZ3RTjnB3PfhJ9oN7ibnIFw2mWCwAMrsUiOTdth
bJO3aIYOvdrPTBIDX2MgkdhtBSCDVEBuGHiV/c+EC6OObXXTBsd4r/tVCWq6
FL2yni7+IQgVikQk4hAUlf2qxUR1U8BeObfm629ZVK0ZlPyqzdrrAvUp6NZF
xd3TxtJ1/NGSv7g7yDwPFs0B1bDeNabnyN/KQm1jAQj7VGOfTiIFJEwMIpDE
TW1oGBgdc4nsgp2dJxZ5qYPptWbbXHRVWmmlJSqp7BnX+sGvMhUUzhtMbfOE
rXHMcHSaI32Le+VTUHG7hrW6Ghc6O5gS5wh/klC7eGOp5ICO5MMxWvfQoFEz
3958CgCqPxT35sEz2NoP9WGxA7ef09Saa+fWEJXWoyUcLkGbQOjUCGTxkQbL
lfJKNfR9b3iYDyMeN0qBG7P2kTEJhtI5D2+8Ble8T5jhj5/m0eS5QniNxX1G
EzcsN42pihtJ7eMfJH3vcY6omWp0GRgrmKFXHna3hG8Tr8mPMxXW78DzzExF
hRyIwupur7QA3LCZx0BClUK9knY0HzAwaZBiniFoMnCMX8JSDR3Lo4lKIiky
PSwMI1fU573psJwP3Cf79W9/aZQc5nHvBZppPurO4hYL+BpeIhafqTrMkJ2U
MXLd/Hd1wrPVK23tMqyIWxVcuZbZganmr0cFabfvuefIzYsicyIEpqAqcIdI
F7bqR3MiWYJwlWxs3ftVi+BjCp1LlQMleoOwa2bx2cXTPdE20CyWOUqeAPi/
XSQ/h0RztZ9ExvG6z0snm+OVbCf9H6E7G8NGtrrt7Wq1Fr3ENo2fkOG1rqnw
xJxpE2EpVWsBSop9eBUMwIhFZHcNmDYAA2Gvf8/tGOUNNbgmYfSgBUPQwLt2
Kbv6plHJMKgTL17MVo714V20s1RU7h5oivHk3i5avC5Jc7VcNzLea9PHt9Lu
n7FEQh91xmmB1FW0PcmZzbKKzY0eQQkqW0daRPu9oZ5meIeZHVjBJKaQq8/V
7rImgPQ51QCePxYcH7io/yr/LQGDJ2dr9ci98esrll/szhhejjmWUhOI7bFB
w4tHJ6ea/PButdXlrhow8U9tOAIrAB1009tDMQAq9dJqGypdO36NbWFXPsBM
xeLB0YzFS9pODLbMXydTRxC4rgRTUwb7ZPUVCl9JSz0n2w9XQufpGREriHwH
zFmUBCVWd+uyTt8OWAxA5x5KS7mgUiKVIgi8TQpH/m7Aeg0Xk45Flq71/6/3
9zB1YLd2aYR9PBDESEy29SHU/FIK6qnJycRO3xdWTOCVVWpXgJ/TIpCv1mkH
/mfhl7ZmqyhRma4kCdulb/Xnni+OnAN1FssCIIadpX5IRLUO8i5lQWCZVUvL
SOMpWMJI/PrShxDaZLpZt7E9JwDIoDSJti1ysfVioc11ghZh5wlfq3IkpDv+
NS4SK+/ZZnSGD9xAHTtvy5UdUhFEYKv3FoDwZd71mqNbQDuIJZrN/JMs2x9X
kRwtdluAL6GAaQ1dtAZCa00/GsDsB9AB0EGoYzskMdB2oqJycZJg6fRrum+w
IxnmnBPxIE+x4vMNkPO9VU9N5YDQ2RsPvoLXD5eJiRMNInpSLE0+6zi7oeWa
6knbM7ZwnmosyOePG2GuF6bwmZBTMnhRYAzs9hhOG8vZHcrR5B59C1ixkUTY
0Mh3hgrfKx08pUUqZwQ38Vfs6lyQNyJtXWnBdibaogT6SPtM+AFHyGbUbET0
xqoi8wAjGQ0QiH3ubFoHMyKaLxP1elt5flqWkvxF8Z27eCX9b5rBJnIAbjTs
7VtRkqfmpDU928tDv3VMJA29F9gtLfqFaHnfcrmy+fME367R98Q/Nie2rIAt
6MPqaJvnYus/0r54bvBuYqltnpbhgknb6Fufh+i9YqJ5QL6lVD//SFpE0r2J
qkLIKMp6ItoBGNzxPKmKX44t82yW9CaFKaL0CyrxNtRUIoWZlCyBcr8nS8Gh
qqvOqNEu2bWktGL4mpGEdkDlqFrpqR13nMC8S5/EPbjJbaXkuyK/1w4CaE28
j8LUKWHCkDK1/lUcJ55QEEgCEGH6lLDUzCDZiOo37pknb7xdfwCVUF+KpjYN
xA4o1/QXakbFB54/KNMqVuK7LAeFzhxdBQhi40K71woDdaTx7OpTk08KnrYR
fTKPc9O3xkPjwHeB3h6SsIPPM4wtXkQBGk6o4UDbnsCbM7mvxZrrHdbP6eLG
PdzOaDP2UXHC4kY3ElFhGvOwloNZCHFtMr70LEUXcPKga57QvFsn1U6Lzjp2
4iojQnbQp4epSW6mCi76O7RzXFnmLuI4dDeHWItfh5sbUwXv7DuBgYIe1DXj
QLGzRL3ilrBtMer2E17GMxTRxn2pGPvEJSgj0CkMYySf6+nILIcQgmVLdS9v
2fWdyWTMc4Yw0/1inOnj4XRrASsi2d5nHt+gX6bmXk7f2QOA3yqUldGgBZjU
X8pmAokt9BAKVaciFPNrnP9SjzuKMTTtOV+Eo93dw8hD5wMfJAFJEkZy9c1Z
V/wzQyA2gUBOhkPG96F16GJGrgcch+8v3u02a0RZH29lXkB5Lzx9zNA97/s7
hsIxokhzADR4X14PzUeUjTyh1ZaAWqUG3wSxqIwwaeAl/aflDdKqFf8ALB5+
zUgzpszqfdNWtCh4CZ+EP6oCq0W1+6ICKsaliR4vlPRQkGKqF1KU2IKjvNbI
Trl6uCmTaHzPd/LL+5qizVmCJP9JXQP/mP/gvWnZL7VyJhSyxEm6X0tvk/2k
AKgwgKa2YaJQLxnayrW83Aj/Yso2Z/02X/T1UvsOQcZJU9qxpxdfXInX47eY
L2ukhs20MErfvUBX/r/0WdRE7E/PhdYYGafbYaT2rs2mpho3gY6FnLGpObtw
Hbz0C3ywEUe4mYaYF32Hj798oo85BJjggS335fb6mmgRJ/XXuOIRHYzMVrTY
30fMJGF0Rqm48n6m9UVmHFAbh9twwYvqKRFGhNVpmsrYkyt3JSvXsXHNXDzV
Ft2cl3l2tNzNgq99JZFF+mNZtI7aXxSEufGcAtf5dTG7006amqNiw91lZwzV
k6A0Ut7EB29pYcFeLLs3XeUbH3sI3xddm8F7SE7uPx+i7G0xtKPkJHgbMNOI
i1WubA4IYkxYTlXRA4rxP7Jnzps+cdl+LMagmGBgSFZSoC1k5EEj+SzhfEIn
9n/Msm7s4nz1k+cLizktHe80ArfPkZp23G7vM1k1YWAcGFpTsKcGM4QurjbP
jrgWUhNDAiLN3xThj/ZX74aqeaVbH/kwgMSjLbduJ69aZuT2t8MUGrp+QrWw
seT/AWPvrNl6avkUc/11beBJoYTFkLAaVHxEKIQ45Ne3HNKZVcYEt6jP9FDj
kDIVPzwXPnlR7ITYeFif760bpSFz8dZkvzrQi/90RQnZr2Db5IMZtXSIeta5
ldmnFwbrgxYQwKpj0uJ8OH7Tj+15k7G+I14tdLQj5t7MDrOsTQQaq91Lhm6I
tPKGrLR46iRv4ahQvingz6j0PeZSaIJ9hNJn3PVE76ixPnBA2dosYe+Em/fZ
XJIYg5ysX9AjjypyM+bQy0b376nh7DJhYHUFZ/K+LaHn47/evJrXvb77E+z/
lSkPL84ykMzHZDR4FLf10Kffxr1w13Nl33Wb1ie7p61ARgwYw+CFkaHgXI74
oT6CmOJW9jpyPY51Jxq0+MbFPAnlzYgqI5UEuG2jo4XKD5q4Q4o0EX/6k3+q
sbiSfI5MAnempt6NpiD/puJb7vfH223Z9oz9lvbEIgM0f+86ljXb/oBQHGRy
HKIyPtEO9cTgWEsIzvhDG7GlHS/Ou6Ym/W7hK0YCU+C+PqnGSBKJgmMcZ9H3
WdaT4xUKZfmoWIR5iNsezKJySftBqaH35qCq/Z/NFXs8LYAwaPqyk602wihV
7KejYVnBz4lmVxpzap+AEjyA6TVxZynwmEWH0/AuE3Iv+BK0sb0jE0SCuY7F
UwDKkw8DSBg4WLUeCnIUnKs1jZ2LccLwe84w41Y7IaerepLOXFnHZvCs+GaB
FAEd4aTMEN3CxtCAehVNrQKwESp1PoLsGi6KG1lqL/F8wh4UpiDe4Gu8gkMO
y1R7PcckVd8VuAoQz3C4/EqADHJ6zo3YvDt+Y4Zw2D0d+WpgaM1HtqJWo9Fs
evRdMnLFjQkn2uEmHOp1FFM2y3HDWe84UsghHeGCR7Eems8uKylBvYcr+BmE
IB0NZnz54oTnBAAVjqiofUQ1NdP21QuFKd8+fY7fa/s4xGgWgfyrBitunDEo
XAVD2eGMVTfZc8H75QnJgRGMISUkawo5f7arlgxK2b/hOJNQOBOLDecx+OEZ
AR2do2gbQ3O7OouQbA7OspSd5oa8Ycf8dGMkloXlhK9KXK8/mmItdOvAlBlO
63t149sXdd8xpuK3Fm1vFX/KW1ViBR3K9U0QjG3XX8VJl7dLPhW+Mzy1eSTc
rq2K15OjNmbksh+Uk1VeJroQ2yYcPH3XhnjC+dZTqsd/hNOoxFf2rkEX3rWp
n5QR4u7BhWveosfal/p387ItmNg/gx1SvOasJif5MhhWZZBaeTVK9Xv67fzG
B3Rf2+WQJFKnijIENERBefeXB897ToJhs5x0C7NqX9410SkYXxTjV6djcldQ
elqj+54LUSxAXxvP73AiAKv3bQqrfnAEnldSuvsSZJWYKFrpVKhEb5d9uYx5
3BhY1ui1ZKnWCwdoPRaFcKNY423/x3nHvrIRVEAXmDh+iESURnsF0Z+uhkq6
DOKI9mCaINLsyp+sDygLgSyC5UEelxrSzg6j+D1tQkvvrATM44YhNjJluVoN
xVvr+vC4LR19YLRRukCeF763lpNDJWXQ4L/pI9WWZorjveQD2gn7HIzzg70J
w055i4Hd6sF2Trd36GWfq07nMKBZDKhaukzx51wjuDC2RX1gm5Zpbh5GzE1/
WsHDv/TF8emmvfWMlXzl1EEHpY0JJWz+vxrVL0WJkc/vCz2OXAhrenUBM0fk
TOEDbSYZWNj4rMsuA86daO9slBNKpsXM9PDxFWaWs0slXagQ+pC2jTTTzglN
NG+k2F9H4mlw1LsHZWtiabTl6NsKTaxJU8sCoECelHMgCx4gWTuZEYpjwMWi
Fe/O3VKeXYrhlrkLPo/f4A4xkB3SRHjFtgadmI+3hR0hiNWmU6US3CFQccit
Y6zLBsRmlMLO0ZuWpmjRgEouytseKRVS2dIlh1EcY66MEdockivGjPpAFegJ
VUlh6I4VrsHOEDD36s/v7fr+9EOyxeEWpfRruqwvRNvlp8oxSEdBmMo7bdCs
IY/JdYUXkROPnOWmU+aBIVfQzki+S384n/yP1Qveuqk1d5H/AvCDWQiI46oI
+298CR57XNOrDSVx+foxVt+iDfA0ocrg5EeQHCf4nlSd4ss/rpV15jfBhKUK
UWCxoD8+KfNm1UbSdPzfW+ViWlT9z0QQZwLy95jVskb3tAbJLP0hPqEo3b/g
nKnRfZfmBDKJjWxz1cOlxCgavQJhiRYLq0MdoENCHJyyN4eamOfmvXBWBJqv
FUZiJodnN2MxTLLGTq//cECguh9xr0Ie8d8CiMWfKbSTCkNyhEt670ZxYTZo
1eyecEmlTZIAaiTYCDA3oSRjXWVM4x1wO3JJlKAc5gPf1TlYSM7RZUKt0734
TSkGctYzesELZFqMYbdZ0eide7DU/fF6Q1uSKp1UKPrH3MxvByuFoBHK20cA
xPJFIKBgAnLIMyGJyFghoq/NcjfbKDrqcdwA3G/Lv4naPWphirRweW/ngDwv
VX11WdxjzT23sOFqWpff5s4wc9ROPpBm/fN1FKJtl+SpwxLPVIRbml9UROje
Vl19LUoYSOOX7b6JyYPguEMkO3IUUVyPRU0cz355cnd0lDlhfYUOHd8WV5x3
wzkcyeNMMM1+L/44S19sxUNM/RtEz3SKkxEifzRWM3yMejOn+QNRtaJpQt/L
wBcW0mtGGhYHYGar1qaAvyphbH+2W2GIfHa7KGn2Ri5TBBYHVVvTb9Sfwb4Z
GYQ9TGmGZIYIAVgqdRl1hAbIjIXZj61ORWX4sFz5mu0xvz2wSU2b/CtokrNv
o4nga/jNmli8Q45pkTTmc+J4AU8QyN6nDbxDYAIGrv8gW5XLHPTnBqA2iZtR
r48cOiryJ453lwVAKLMVgEuvjyp+EMQapza0AidZFaFkhQ7lEv4tFExojmFZ
9NHdL7X3e3J534Hgpfkv+G25bHUYI0qAaC4AZ7/7sP1vZuV+MmzF7RX2loNV
SqPnbvRenNREjWMOkBHyCzlhSsJrxbhjcT2IsEop8DGIhcvKsIUXIYv1T1HG
H/x0iKhPv4PHxwVdYrrsJfhepqmloe1lNSPHrlOnFm6vjrXZ/t7GiRJmJRpN
4aZ6M8O7lslOHZK/pmT13WnUErfk6TcaaYrubl2G0K9nx6z2Zb3fwT/iW9t7
WN0swY6fDT+0cSn5hRJKUiLl+U4GB6Mk+vbPEBczXZp9Yi2Mzvbf7ZkgzcvP
G8Emw4a62TRUpsUOOndJMc4WOMzXw1i6V6hEHq3JGrr1qOYkXcUYmgDAsid8
f1F56Ion2SdlU9w02LrTna4lqgI7ldChsd/7SisxS7FYt4aqymuCeyHpVoUj
tYv1AjAAgNX/8caFf3OXIfO9/yVRAnHqVnPacLIX3eERaDV2rHmBEklpuECB
U3O+L6lhWDvqxELDfpxbK5xeGHft2GrBhPtzNq7Ic/Jcfu/gsHtqYRRkAwQ3
9nktuW5l6IteUnmtxZeajSw0Mcchlykjc8ltVcydR6Aeq1+3dV4XdGwCd1K7
smkBxA3E5VkpYkm0xDAa3Wpk0VEYHgM6CTc0lp8Fo4DWpBhCLJWrCi7Z7oGi
kCwloXzlaJmBpLAgAsNQdONHiWWUtl6whctTA5P5ovtlNlpkNA5Ay6yNFXxz
WRgJLsTvBjB1lG7wA4Vvz+e7f9ZKO5zgCpgtbr4FR5P4DAgq1ndXIWn6XXLq
f6I3hi3Cu3CRy1OAId07eVVjzdWa+skqxsk7DPETy5O72kaX0Mu3A6X1LAnd
qCesEVa49hPQkhS2zV6ye4Fh9rSXV+BqorX0ALdBjWN+gbJ5nSqKYySyFzK5
/TDW2IDnzoAWzJITrcGN9uiBAN/ccF9q826ZH6j6a4zkovk98qUzpWjqQzA4
QpVjoxmjYTAP0HQAtS0xddC4q9s28L4Uu5kc8g3COcev7HWE70VinYaV8C1g
WI1nSdLcEGqRtaE9tjUWc2AzaVC2VgYJUYOSzQkffATDcleobJcuwVvaA9Bh
FtAKEY+3Sqh5pf5arsX0LMk3Y9+cqJkAp//jWD4kaQ9sQkbeAU3wmBu02Ha/
xrpKGI8krmPFfCllrMx/XlxlGutEZgl91Kh0sR2r/cS0B7+/2yfFvzVCePcs
enBj3hxRvGeunxRdmVNRSJH6IQKhAAH5mQv1/T1yoymLOOiwnn3BWUjFSyqt
qdz6T63SUT2Z0PkX+zMu9uJshkyR4DMehrl63B9u6j3rB6s6FVmkYwO7JqcB
YPGPW/9QeAhTpVDAa31yLcXDTvPsXwYZa+/sWCvM4qkPGgcn5m1ItMopIHPJ
i6KGMOqYHcQStWRCtQ0EjzX94j7BobDoHeo3VIpDi/EEnnNx/cpYLGDaSMHj
ygfbcCTgUOMS3FcfKky4G7Xm3UkVkmNMlkI859NkF1XfHqo/OCYd1u4nd+af
Cv1YGS1ef7FxfkLB8Stbf620m5mdNWv1zTSucNtsv56MZ+6naooTLru/R+Oj
AcBRcd6wOYyge8q6rFUEz5RYz21Wm7KxOymm5TXeBgErgJKIZsMgq/4sUApc
XyrE3FhDSnpaX9Teo0qj5+RVtchX8NWoWDsvfHF8bVOyBlieRxE/XD8JkjK/
hkcR3qRD4EiVtx/PZg9b4UlXFc8P9sWW5BkabfR8nDxeU6i24lckvkmI1HgB
8ZGIWMVY624SiKz6CbPRyQuOArJhl1eR3MC8EJJYHRXXPHageD8Y/snGSHN4
7hqSQ+AlPJMTxDIWR4KMVCD+ZZHFbtmuzCGF/R+oq4ehvibImScrd2q+YGLg
BaQl1MughQdzMsGiMFoBDoIeKpGAXaMsEtCXm3pLgpoP6H/Kr1qlAwAAQgcJ
322aYG5oos6usb90w+uQnHauovZNnvzP9hm36zLGD84W9pdT/lBRnFYECjEy
qnS9AnctAzz2rvghGCblSItmZzpujFGCBNWZU/CajihLQ7YG/yycZvPFjJG6
K4BdmrMespmmtqKAsvRhewGA0Fk0jEA+cJxLuVQ6ksvMpqfFBlzZem40IGyL
KUm27jwapJYoryErxFAZAN5bYIL6xCP1OQXC6+wzy/XNVcrjrwHS54tYV//T
w1J2jvHF9vyi8KZeiSK9YCKVoptm3rF721jiz0yldIG9Ip/n38hD6if/rQdm
Xjta7MuHWNEeZVTDlZFkOqJt4y2reaH+nPVrphAIelw2zUoz7RSF3KVxYQ6T
wM/HlIlaUnNvyUnzIwOspVXjU/nOS6QHqVIFUbOY+vN83/5tR3vz0maQLXgr
xhZjpSjB1nVaSe9dXpOovuxCq6b8CwRYbFMA42xWSHw9VCMkKN/9YxBHed0F
AYp0RavB/D4LF8StkgtZkZdvo1HhjckenTCytbovj1UlpWWH8mijU8fGt7B3
ChJC1iXatQfXYNg5A957ACz5H3UIEJZcGJXlWEaOq/o4PosrcCg3r9B4U1ue
cNVoppsCGFJWF6+gdAoISDGXVXe6B6pQNGA17KAnDFU4nJ/bkqhAhDwT0cwZ
Owmo9OhdYoyE2m2+vriK3iVCdp8Lc+na847CWS1W7lfScAx/104cAHGha38U
BpD2+yftbiCFWovtN6ecH6vo3bkKpyS6idBKT4uZJFwbr2R+8PcAj39P6+Xh
raYLgi9jjVvFpZOQxzvMmtj0W3Ef2ZcJt3s/3R0iRIdoVKCxkUdge/bH8sj6
4ojsNjU2ANagV8vNoSyX0K9pHOqyo5qNGYyV9KVwfap2P9rxO0bUWhZ27QQq
hRYU5lshpDCVIQfLCxXYTnmTFywPgjOL/ZkNHjLrsseJVfjRKf+FbFcMcPcv
ZBYIaTRjyy2an9fJ2Vvh/jK+hgTj1CynI45I9DRDN+kZtA+XPoOX8IeF4ygt
xc8objyY/ZmID4iLOjcwzZEFwO/e+tpabbS9f67Ty6TCCbO+EkmYV5oks1NW
+4mQ7hgbGe39+fnqDZI+BM5Xdmq/hafocf8BBK9ZmDEhR7ifvXZtu0uTOP/+
RRBQZ6i7hkbZ+buGEm8mGPG+hbp7+0AkSYDgHY2ywsnFqCb/34jEKJQU1SR3
wky0IKUZc8+wKFIsm3fWxlt2N+4r1W1BB69qL9LPmfHiDvF1zLy/KjQ671cy
5Gl8NLxCtDkdLH6VHJ6+ybehJIXbfCa7bDhcfLGQgq44d1CMFd5arqhNYzrP
uCRCfQBGsTGqAyJPV489v57HgmqMs/F+MRWFaJymSXmH72DUS7/DlR7asdS/
KH1eP0zQslNEzMt/jOmLTIqW4VbmVvxquIQHtYokxcTkubVfmz73Kbz0Mm4A
NJxNdk590i51lwphRi41PLGFUVhYUFamN5MI+u0Dp6Ok5/cZiQGtX5Fsuh5k
gQNS99XZZclOeDWSfit3WbuWGFCC4Yfhy+K+Znrvie0Jfgs8NOXivkHlQeJB
VudQc+zzDFg4EwAJzEt1GuH3SGQ17nsloZRmM2M5BIxksYVsYGWzjotBzuwY
mqgwPQBVinTwGkqgqTisBR5RLdQ1EX261h396G4M6S+N2j2mAubJfcr/T2IS
8krMZBl8CZffjoMxFhJ0zzvXP5E7t3Gom8nein6wvfgOqvozOEm2cRdrcz1O
w/KZ2HEDFI/0utZQT1mE9p5aecmJrcrvzFn2pK1119aa1U7SwXvfH+eQbOcS
ORY1XIx9wwkCa01LdD4ZSrrCT+qExa3UXsZVy/zO6AzXWcvnA2yFpm05uwIm
iSwZsGpKALUce7lrnLGDmA4saMG/2RGjpBqvqkKb2EfhLV3Zf5NhF02oUlj9
nhEg0dCIOy+fzfuYLgdyp/wLa+kXAuY5hmKgeaFLWnBoqThUWT/1UbtQ2VAU
U4HG4QXmoDU4jeO4AzZIpawjGlqyuAwwYTBw0jK5LZUxnjltw7rpUPK7ALDT
XlPTFMuBpRWiBX3Mo90Y4lnQUWp3KtzhxkX87fxgwPsDVwjYhs9ng2z4z9fM
ziYURgbaMTioQ91WqgGP/3qeKukGbyDh+/loodaZU6IXCiDdoWhuHagwB4AF
Pqpm5XFsK01mB5D0wTKQRUK1o5HNYxKo9Y/ePJevRJuehPqe7sD6EnMUH/NP
Fuz+6UNG6v3awIMb4l7p7NmXwt/Hacu1602cJDISJfDqI+SIu6yNoUYIOXly
gm/KFEXbO+k45/30/nurSBPNLP0ZEY5ivDScVZVm9X7nRYO1g8dSQhBClK62
4QhKJgFB0hwDalGf3jQlonVQxFfI9PrbEb7FG3IZAhKY57ATaHtaz6oq0EJh
ins9Oz7bFAOKiI5M3UdcVRf/x3YibFbzVcYel3n4FphGswzSivwEfIFNbGjL
h0J1awzrjVQoi1SrmNeJLcIsmaDePn165SyTq819SiwVeV36jjtnC47Ptz0c
AMy5ZBXCMK7SnvVIEa3Oa4Tkt8810kf8jbnoc+gRmiVi62z9jrAN0CtvxvvR
Fg4Ic6Bz21WmnpHV9sz2DTTAo29qdiCeoE0KY4miRam8EbXb3C18dqV1BDiw
If1/1Kgl1sSULnNYwW+XrP4BYHXZcWMEtJ2G+jVMKlMV2MSVgQ8JhCdYyFEd
Rnvd07xuHt5UIyd4uLR8SorOGtrbOhQb1LnZKr2cgCpWKllP9XpiZM8sIbGB
/wSzObgZoInBUVQJntwXygsSUHQMom8d/fVc0NOFw38trdpQtHRObaDCsRbI
fqXUAaj7aYnoNBv84s8xWpRYP+PnIph9IvG7XB/+Gvn9Ce5WRtCzdVEer4Ih
MRIPmMtpDWsiwjlq5o4cDZbxvrrcrnNrO9yj54WxGzE0EXl29/hGcxKH3Y4P
oaNE/pcXl1xCj9lZXXAeTosjTw0DWWpKqMs2OZh9TavhST89yd0b4tucDrXq
Jm60sWGFyV39i3qkMEQ6ZSdnovui5k09xRk/mKFwsi+CO1PGJJrQv72DsK67
gg3j79EawqIMGZCbZoLRxDWW8xBLYfq9+PVddajZijboV7kMLfuXRRxD+zAA
sDQXxIQYHmXXWnG+gmnLQDcbgs4PverLeZuBip4PL8050yNiDUDwkzssVD2N
CssCyD/dMcCEAmXSEixrCphBSYDPmYjci0onG/W4GVeESxJ/mCZlqRseLFt6
XL16L9I9oZNyq+pL9c8X8Qp6eG0JKNqnIt3I253fwFNzGnTE7xZTfqkywRSL
qtsGuE436UsSn5htfRCj9oAgsMh/zhjzuucdDNltH2DX5VA506q4xnMxSZdH
n0HQjQ2/Kra6bMP3YJf4iKstPHXccDi2o0SO4HdDDnYTJIuFCRgC9n/kfUdH
XLj/xQTUs/Y075Bky1J9n+XcJJgdk01TiXhkWu1h9N3cK90lQ1aXqBkCR924
y/0ixIXDhtUer5JHdMfBqIhlpQo7mve0QoPwnK195ag7Pq9dTjv+DZ+TayIg
i0rk3xlBLAIe9QaDjVrVl1M4GFW8piAuiRd2Fa1MpdPyMoWG+Yxq1dbxCMcN
SbDA7+zS93hhQ4Oy9XwjeNbB+H8EhEFFMWo1wtMBuRi6lhKOax0XuG/q0q+2
HEZnssVYn6SM1rN+NCdC5nsFO/klMNXLgfw+zRJ34Tgkhe/YPKLTR7VyfqwX
8l48QKxeP4CqyqYLK7wQXVurDBKEWTQ8HMrfw0MyXN4oeqDoUYLb7ObRR2Ep
0V1D1mMg/j7KmTD2PAjt5zklcaVqLt46nrB0P1ForeN++DG9yh1UZwAFe9dH
LXcnG7Gmx9At8DfHhN8moa+YTvYOx5n4/VU3JlseY7MuxSd6s6vdc7bI33Gn
FfC9ZSdS5HkUr6hRvMKew3L/wMkKwdsC/qKMKdTGl+KyxSWwWoV4ib+JrInB
jAoQcoIxqjOg9zW5Dw6eNauQH0OulSG++Kxr+a+AyMJSaJnsP4lJs9mBYIwP
jwRDKePMHqVgHfQYNMKO7eKnl33itgAT7fXZt8Hu5VuSBZyYszdV7kfRhyvX
Vm9Fpik9v7yA6LPfcGfAbTjsODkp1AIqI/caw3gk8QFFd32k6pKOoC3jYPGa
IthNNx7iZnf2MuEDAIPdkTmuF69K1JHEj0WkzJRXnA0ndqtz9LRuHSeH8xPJ
mjtuxb6ZA6ai9hs9Vvp52kWn2JGIPWxw/QQdDirz8cm2SGuOpw5aHBrf+Xzc
i1NfvIkgrZadE+8/XJbC51lx8WOg6uQQbZI6TBBoeMmovQTCFywVLdvtkYPj
nF2ybMi/kT9G8W9eRLCc8qV+ut3owMrPpoP0RUgNems/9ECevllspsnMENTb
nh/dhZjXzj/sH+GPral7v35/oS91XW4oP37MABTnds0pv3477f4JVpdp5JQC
F6J7we/IrC475O2wOQSCuSybHZNHKZadzN9Av8BZbuV1HoZsGxaztBo0tGbb
nA7XSF/Yww98D5P+S477et+SFH/g+vNqHRweC63J0krWd7SKwBDLYOtsNq+p
mAtKQr6pn6YX0KU03YOm6ml0KO/G/4SlnIvpevd5z9AN4nWnU7szkPV0a03C
yf+vKVcCHLUHil+SXHEq1P/xGDaWSv/aS/he7dKc3spj0LTljvpUCFjIMoQR
PkbYYz/0YTFlj7WHcw84/UD17YfTEa8LghrIK10P4FZFg/LIwAaDw0JpuNUm
5IRn4WsIebz/UP8Qn72K1uCv/qDJSxmZaODfs0H4fwxhrwNTwy0l1P4l5tPJ
mj/KczOrOcqCONHWCvLYC5gr6DUsVYVqNoWvHqKbBzwDRiKdyypVw9unIWqM
iygIkz+HPrWFTRdcrnEL3w1SLSkckqWxlH8i7mnXewVfRVgSpvtPomJw8Tmr
2l9AVg3OMDkrR9WrZilZ+bXJg7F3W82jopzkG2lHSZ1LHSLm4yqCs66e4DS+
2MvRD6r3kcQoRa52uNAToo71qSLYI5lA0PorilDm0rL1wjk0Zug8RYiau5Cc
d719nYUpVnFGM71a+z5yTm/NH10NTRIlGOzDqzYot0PuQB81Cna2ftjuZWUF
wOWny1hiAglViQS2pIN0dKAk2GCsnLXXkJNn0S29iB/IC9TpULPR/ZZxEb4m
C63ZIuI7IT8FLDS0tvYVNKktyHt9O7N7xkHnP0sEbiSkS/HiMeJZNCb/7zvB
aXGW4ttFnZPS+S9lcqs/WIe1c/w8E44NAbjCcKn/g/2CFRlKzM7DRPc15Ehc
lR6lMsfYOhPiXNJRSwU+KM60mumGQepCss2spdvnOCkmIVW6sIdCLdxeK4Dv
kjvgmHYYFyMCqqLEmen0K25b8gAcQXDT5mqSPfTcDoQVVGs9r8PvAVDoCCXf
g0sJ+voy/GlXzXoxU6qBuEsmvrjQJLwL7kxkgoFG9HsL/7wJi2ThH9r1sNFf
lXKRR5Cgiz0njChZ7CDZrIwD5Ni/26Emq8XTwnGkQSK/UyGshrBIMqGz088d
e+sTUhEWMjkUwSlb5Pzw315VUtzxcMkYbs4pyScbYBJ+vdTh/DkyXa5sDWFP
WwlEX2ifW0HTjIeKF6HEdGGhloSIHDpKMH1Lit04KIPFGIt4Jn7sc1kxPmkx
WoKUTgvDN1Pi+DFgEdB6sFBmjiFI4KbUuZ2fM9URadP2SqERt+cvFsvPEYIw
ptL4/kb4FXNI1ftkJ7KQW38u6bIz3BMJDlZf05xX+mhdlsfcez4ongL4nwf/
ZiAo8noWu+AAoZi48jnN0T8NeAUkYtm885SGYY340OnSCVT4asYefPQRXYbk
UP5fbJ/RevGJrSDctquNrRRgi0R9M2RtC+q+HArDfmn6Aj5J+Sta6bTLkRtj
CmZ2CwjzLjLvZ0BNH0t3ocn/vTyUactlyDUKv0pICfwOCl9cw1Vxd3Nbxsk8
lMMl/8Z/oYnxvKwdFmGp5zymiDQPGIzLPoZWlEvgosb7WxKWdq02NxsIeBI0
u8DW9DumWOJZ5MiL8u1fvLjb5+8Mlp1F/UJb3kL39kkNtZxxyknjUtW476EV
GvKCj5A29uaWb9r3C/RvLUAU3EVsnMSSkh2ovMzDy+I2yO0EYhfCK/UOcDE7
Be6Q9ZKX0qTBBPwl5WtwlBlj7OcFPfgWUsIDuzvWQRmENFkuGDuXZcqhlMJQ
1p2Xil0KSPN+uYVsj3g+VBUk8mCHFQd89f7jcqyJlW49JXtbAL11xTj4XqhV
XUEDPY8GT44clp3seE3rZJuspekdQpPaHV5+7PzvxJ1QKDbp2Qw4Wq2cE7/0
vQZkoWqx0hoqc5xYOUPhxoXsHK7cAXth+FYQ8yVNZ1L/jTGTvda51JJgzxPJ
GsNyTKmmpAUV0iFVBtA6Sm2YccZiz70EIFDa+7L2V2Rc995j4DWUfocqSyQb
DhEEveelLx7fnTcWMmhDP3ovCyaEIwPpI8x/9MxceTKlH74+qUL3/ZoWtqrU
Z0d7LwzfFCcMOOZqGQDoaqal3QnU41gjQ66EkL9mNR19KWpUdVUCfKXZ3QTz
PeJemZnbQH8aannLXBD5gxn3s+DTostX37ArwecQtHEPfa/64gNleU/sPNr2
KrdubeITduszizLtFXjwYCnyJWPiBWxd+5LlnEOR2oSBmEvG0Ew1oFxn6Dz5
Oy7FQgm73QTEeEb8w+1xKg0SvWoy0fDffoe8OqQNgtFyxEOk8yuNLqJ1tZot
okHGEyiCdQVc9G+WYotFucVpGCr2cyQlh+Jx+3A6lBLkMdWHrgT1tEcqYrgE
SvtWGcfJnvVvLqQqGF4mAYdu3XQoeJUI07hy+wHhsmU4jB1Q/vasruqlegsR
IbG1iLeKKw9aCWOM19M8goFd2S9wzKdVHOeYFt6kS7/ZRJvL5ri4bRlPbGK3
ASH5liOV7nRjdvS/bJ4Umq/uwjd9iBvQ9rgbZ0XGT99G7uUECw9kTQpyAB+Z
duwlkWciqE+cWKRPxW1JrooB4gBu4LQHO3iVkerOEoWdQdnCmU7RP8I+RUcl
ytJI6TKihuB7WFbvQiBLGrpi+S+0yttqaXWJ74zMMrKql2paDMLuH7jGG0Dj
DAYLU40JgLNeXY/rRfQDRmjbTg9RcPBwYCHi5knJWgRf56Gip1cfdrkMdbq5
DTVpL8iOcF/hjl3fcAbZLi2RtwB45QDVFxMcX+AOjqoxqYdYk5jtSMDQUdew
9ES4FMYHBNuSpbxIL/o+CovCpqdR4RKNoTtQJSgG0hIotbMrGzgiekJFxdgv
S/tDGEvFKiL0Q/IZhPSvYD9vyS2/Nf6pVFhBvBMrjNdpZaRYBod35OSaz5zE
SEnEpxlxZXETMgauLwnxEAAC7nK7vCwCM2h55pQ9kR1dJaZoOifrv8UBr5lJ
oyzn29hdCMa49Q6AiMj2xcdREHkyfN5N2DUPg7v/WoaB9D7mc1XSTgDEuH29
CIKEqyuCyeaPdEXtWW++4f8YWrIYNMmbEjfSmoP+yRLuXIC+flVbGKFWYrB8
utO3X0dggBjayxj/XSyIludQ7c7n7kUqDItl2oI2696ghMNBlQPFPvp2k/gW
8f6hIUmL+XuaZ1jmT5+q4flc6OQqS4wwqAD/1H7KOHWhw/zZFmqdFZ8A7w/Y
VtTiWV0tdWI4B8pjcYEoVcCOOvRdrbVoR6+/TM1Mrp90Cs5udCbi193dQKJx
MIQd2I8EqSBjHiqKQvlwtst2kTgxK6L5tX4M0vILdEK0IVLRwjsnnOBt7e6C
3uwrwP3NJ2nKoXXGKudGeITLBabUc+EUnw4qAQujgK8L4iiFOWUFzHWCvxJj
ms3BK58zNzF9CWoRIz12Qey4my6FezjoCvEaQe6Ch5d+5q1PheCrZPDwmKMq
6fq4GGHGHmkAUbz/Tb8414q3414k/pK26f1yDCG/SN8q221NnFE8A46dUmK5
xYXNYeUR3mnwJEO6UzJTrzQYLqxlFXRKdqM8thaPNuaOCOU/hmRdxjgL0Bkc
Lx05DYP2wFQW8uC9OEVC61lJ+UDbpF5bqn1G2xVoc7K5NGNssM30o3+uWPes
WLltVP07NcQPic/FsdpVW3b1jJOst39rvc4Uy5h00bFXb5ixHINVUjmowzaz
GusM96xC8IIaY3q+eVEhS9p4PKZdruAGIMocnC44du7AhiO92usjeBn5KF29
AgZ6ItlDQdxTs2PIK+iJa6qnqpOMY43MOlk7tsjxtqeBYFfr9mMw+cmqUgn+
gZz3EvIszm19nLHV8cc3DR0mW3NCDS22Uo6mmIfxZlLkN6Mi1i4Ce/N7JPb0
aBNSS4AxHSRi4WbJM8aEhkADj4tLjlFrglVg/nid+KwhbaNxHkERigZJSiMe
5hvf9mPoERXaVPaHb3a3T8c8no4+gKyJeOHkn9dYb7X2ap7q126cWp2UN3ZW
+qHbgyB5H8V+URWeXBNrs5slQCnpSjGe2pWuq2KqJaXnaNwjPjK2ArxPfHWb
r8ztrm7chasAwbv0ac88lLJcDnAg2ASljr8FJIxnXD5i6JCtxQ15IR+GOpEa
bsG/2HTpUyW6Ye851RTF4hPnisFPhuBC4jpg9cZWrWtcji0BhVJKPBxUXfmc
qgZB5w9mISO13VyDLb+8z2etBtH9qmWPQKEfgvM/oquuju+6knTUcWHV4K8R
YNxgbWCKQL/i7r9MOsxirwk3b7512AxYZViYDrM8aNX9gL1RwvMAK4inQBbP
MdG4fm8sHXnqbD11hcb/YWs3O13mZcHJkZvSyAm08cZJZQicu5hcm4wwx0wG
UV0M8dgQQ0lmS+UBJuS3WE2dyYCjycTnWceLKvro+Uqa4ZmYgzJSRrRacGXF
rO7K5I4znbMURC2QH2RjdAQTbnPlKIDN7KpoEADxlgifdsNmjQmzp2TqAFAW
ZkbjLUlle36uaS6OEouzu63omoeoP6F0QhMALFNu3hhjmz27rDQ/ovPipo/b
t3PMAEF54yfOhwYs0UXEJKwN2kTHoeH8Q+7JzYD2A51ciTBkUyIc6uySzvb7
w+42LXDk9ZOGbrcbQ8fAvR+F5fK+8Z30/jDTBo0nlfrUrBpDm+GrHjGZUlxm
GTf9Awybg5ZpSA9wUDHpNQGgGIl2SUADX4CqbX+T5UhSeDW1Hk9ufTDWeOm/
19H6BmSjo/9OTHjB745Qd/HCD5PbPFy979aytrVaBytjmGG1/SEY63eILeAT
WJLbOGXa99GwfdRae36HADVjoYo/bBdIe9Jd1EKrGR0PRRDcvd5iAjuD+Hv2
05tC54U1RwmPT34j34v0FnbDmr9/TyYXBON1VjmKBcX70ODNTgkdDx+B2FO3
b8X+8bJD5taBPpojKQ0SX2q7vQntDRiAv52xU3QgJX12qAQNy7Qyve0dv48C
VBEcRt8n6BCMRzwGcZvAePj+Ahkl7+KXIk6ldSIEbiSFX8cRUsrW3iWAmLTb
gHyQw+5EZQXkIFmC6zZxPbvjhMJUqeEi1F0MggQBV/WZy/76WqGIgNnvPl6L
lwGN69VC/juCPuKkDbm8bIKtRKt34LevnsgaRjY0nAH3QHdBGiiV42p5k3pz
Entveo7TfZh+kCBF+4vgsQ4/50EiaJ2O8Qst4+fz8O53ZgJozKXfFa/rGcVy
JrOnrEXlYN0Hfy4mFjdCJo0YGqN7kOoo007hXowqx9aBaizs5CvguhZH56Fl
0G2N4+bqbyA9YLKbeF7SPPHzuItulxAG+WCXTJN33P4oaKJ8c0tZTzGAxbhA
Ormck5nhiM7elh/m6TKWEnZulVmgoqM1Aym4OqLXayOYJoNHfsxzIBMaPR+K
+mzVIetz1zlKSls91Tp9TYIT6E9pa+K1v8IpyKAPWEa6bfuOigb80BvYg6bC
PaPOKbVLzpMy65sAPv/zwqX5+T9x8v/Pqkje92Wt723GoTLmx+CfgXOefoZk
oAIOa4dEvqtITry08SRuHgPBqS+OHIirNswwdU5rCmvcb25TZAPxoTezorRC
5BKvptygIodEOEhxBG1WcC9W3mKmhCZiOd7rDh8OyKuaxjBs4iS9vmogC3q2
HhXHoXgjO0fO+0Pgg6mzeT+w0yHm4h8/0Zh+sb/0iJYM4G6Cml4+LvqDWENK
iRcb+SOCvJvR7O3J8qffyirOthBwNDpyWUVjSrtKZLfNRIMILdkQS24szYBr
Gf6n1q/L/kI3kLE2ubRCvaO3YWs24hsvmggUoG2Lz874yb4ygVB3mTZd0ZPw
l2JIJ/t3DZX8eobEcdb07JF0ROHo+9PYzVcc+DEZ3LFUjS+8C7yo6xOubjZr
Wbt2FUvTASCthJ4gJk7cPsFVrkv4YyYTVCYbHKAJYEYrvIPKL1VnWow0ypZ2
fzzY/b3RiPKroGFClQZLkfSI3Rf73IermY174VicsQ6gkKojAGWb9gz9UDn1
/u/VMx/B2DPpr+GlRPUI30IcmSKpKbjwW1L4d9rJffgRcou7R9/yJJxjeBzW
2lNisDVtU6zv05ac/yWMUsok+V0RwtjzdVi6cnqUJlcVvwEh0NKj1/nPf4jk
2/KBJ9gMprXmxm1GHmwid5ByFw+us/726r95LxCQDQhlcQVotxthLj7ooCO4
xDUMN+oG7Uj6fwH7XFjyx2j0oCcl5kRije2LwJYihpEKJfTo+B99kkFZqTrn
EHDt+vuPB86yHPokkpQjYTJZgYOxIR7s1ZK5eUgI9DG+qHxARrT+u4Z92uTY
PZIXnK4jsQ1DAHWa1nApesGjcVtxKyUtntCkoMDQtb4LDa+6rFp1NjWys0e5
6gIoAVJQCLoG47M1SSjbdinIBaerr287mKXBHm0u5HuVXW12RtzvIk+Nm4EK
72k6l6BNkS2VErvqbP8dxcD/p4+g9fgc+oOYo0v3t0jhcz2tw0bdZyMswxQ3
MgBOb/mmoNBvEu8nLt4Zc4Qf3Zc0j5V0xHX9h2GUEwBRKj3Kq/6fdeSQPQVc
TmS518a/gi7Q6M+ppn8CIFDGxTdUAN2eqfLu4JZrJ/v2XacpSqq4J6tPJbVF
gpKxDewbTtZXutQDyPOxFwDe8Wc7N/QkphhV9qGhFWG2l314s0D6wTaxVv9R
qcm9NBCojEcgnUtr/NZaBboMkB3gvFgye8IZtXHGNJRcBSretLhunYyi2wrV
k6bMP+zEyUmJ8mP3E5KW6/dv6IjCy+6KzKpzY4REgCBpyvVsAs7EAaZvWUGB
DdipIZy/YZRn+eG955rhm00bdM8FnDTLLyCjo5Sbkhe15+eVNbwfAXSnB1o2
X+ny5jm2BrxIqO9BExS+R4wPFZQYX0v3WS65r6sOEmKO2W6lMla8WmTu+5QU
E97fn6IHB9NN5tlndorfu1SUYGnsrVKBlNkEWv/Tfd34nRFfxLRHyDoI5aLL
tIDz/9x1zb6WFIhrbm+ZcXbDw99tGblbu2VWZkRN08F8jih2mErso6mWYYK2
OT/K3JSa7DU8jgv1dNyRV2KIbqSlW91jXgck+v1YLPqR14RWykmZPbtssWfs
UrsCOyMgsqpXgqenOIPomGWF3V5hS1W3Gy8rs5sjPXdn9AiWQQWXuQU0QMPa
Zq7PxIQSt+1bSCky+AiSUG6becsEgFSMYvbzOpCdtbynB4VfbDHS8JzoQCwX
VERg3uRafjPSTkv8JPg3rSreOhPOGE/bIJ2jNkF129l2PlwZksmJ+ltaZvEf
FqxxPVkDx45nfQykUd/IlQmdMoNOT3J2qAi/MrWwcbb+PAobuNA7fUEnQj4b
M/TnawqQeIcbVsegOoxtWUYC6kMLffU3nJYmyxF2EYdic6T3QdF9LcRV5pj0
NzeviZeJy/JIkqQGnCbq2GYK8qOHCEpgOEHyTaPgeqc8Z/AAUXAUb0oNE9s8
a1RWXrP+DTi429wOfpphIAbKXZ2MC+z/llZxh2FJMmy7RLowr2bPGuhRa1Yi
i6jGDfph6Ddng7H3WGkarVTKhTP79mRhurmp+sl7Defv3z4uHB92S92PKISj
1ZjyC+72R4d/c4DE2BWCL9aNx0Namj2fTD5C1fthyJjFJXRVa9eZqnTISUqj
Ev7SudcXdJ355Wmky4svrnn98py1DTdTPJ8DJy8YZMN4TMZwoFoIv+V748KR
NEsnl529U1xMepd/fARpJRHlSMqWc+XbCge67D6eBS+GOxAQrNWeg+D26kLU
pOQvRjA1W4AhEpFz4gfmGfc33V55jFiWpr50e/f8YH2zwA9hQ3WZR94gxqwg
RGLw8hweiwvTlkOjekk3fhGdZxnjEKM30jvPGRfemtVeqHwHirMUrMAkBzOT
s0qbN6fwMm19v1WT0agqHxWPBdgBtrK3cHGIDkdKE90s7/EXa3An9SmGtkAs
kpqnNxxqaz7iFSKWWBiBiwLU8GO0FIA3oYKucAX+seBBPI/IqJx3r0WK1yro
AjYmwPyMpGzcumMl0U8+0DFa3fDU/AAgBrlYadSOXYyWvu3783+mO93Ym5he
CmJK82FyxG+RWWWVFMxxvcMQ7P5/zhUFVbdHHopBXKeCmqHodyjWfkSYcDU+
lhbrQlThC90H7rzCMIgWtz2S2+o/lcDW7WTAFoT7yumBl//ZzlxWw97DmuvV
CHXz5QhFU6CyUX/3qM/yl3vgc7OvWtEYnMPWYP0WQO9fqFJOWkRnGKRHyBQt
qH6b+TAI1FnSU4nyl8yP9wC4CEjQ1rRL9wB8mPGvkZwRK0EME95HLiOWcu3L
kTV67jHg85w46Q71MXcarUppxpGq9Oi1aNosO1ZD3/CO6FTTiC9kowF4Kock
VcsTaSYbZmDDBjWCl2xIzxRaJn8Uw68k2PcLwoBV5eeheRm4ePQdIjudzmRI
8CEdEmbPybmOHrN5BELIUba8NwaYcmxlRCljLVq/5FVGjHxYlbfJcR+evf8t
XnsKS8XM83V93orVMEhs5bAlXDOfdwMHKtJHv258Rk3MPpKWY5nVqf5tAylL
Xf1GiJ7bJLCq4QrSR39DexOFT7+DvHBGk5f+gxllX8K7wKf0KOZzi8NLfi+n
M8rKlzoAbjOTU2S0hrxsOy8Ng9H/Xv8QCJjI6iUeJdHXz0NFA3vGKMyWGrf7
ihh4JLp+gaBxFsC4NWC1erz4SS7FIzEXppIaFhCoj0F6B6q/Ok0v8BExA9VH
Egt02dUgrUECI598DhUfvuNriJFCzKAO/IL9nNmJOf/8NCCuwD+zSY1rq9rP
Xx7PSlRLbpuIy/ywqx8CoFgaTfOYVUzp62K/fJl+PKDMgx2vxUwj/6M4j8Ww
n+V7w8eNSzhcw43BTkeEGNXEdv7sHznhL0IfemkCEI4WKsHxBz0x1/lRiijV
wDYtGCXyvFnzFU89y9pjf24NRJmZ4oRCtv+oLl8mmf/rvAnXpjqwL7rfP5tC
7Jhq0yTOf3Qvaom9Ojvk9349swvFTCh4lTcRans0ZS8sON5yLH3+MjNh8Jzr
viN6I+OuFEMMIfU2QhePOcQU+4XpK4mRKA7H+6hLxx9eJOfJluYh032uvegu
TSFwt5LhIBCuMw/2ZHYms34MBcowZlvXkK0eNgNB5MzlX6XoEO5ebNLsxm2M
o8gQIpEOXuqm9i1lA6CBZxVnRz7aJKBzAr8ffycKnPjxCuLKSshZ8H+2mS+4
Avi9b6jFKKJ4LY/cUbeXK23lQ6TjEpsDILYwcNtHxaFfhCY1Hcjm658bQkGh
FrBhX0g1Bj15RL6NlMI/8QMAIhuD7HSa29mVnwhZpqONT9qfEvEJC6AtN9X/
66JJmQv84Ll4r3lBjCYMVJDo9pofLmmPC1x8K1z1u0BJE94X1s6pxH87RZyo
7/D3lZ/k3kevjW2q5KLFD5EOsxQriLBrqbIH/RRSgDWQAnIinLGTnw6pc9Lz
t6ICQNJxdpGtnlkEX2BOnhYfvju+dlBPMIkPJXXOT1lboEqx3FMaJpvc8aFW
h/CqVwb7eKBM2wT34UDUIan8RK8HmP7z+j+5CbNxvsWGs2FG8mLi9zfzQoXX
HxNHdwiB5JidjyEqYBGeoyuE6GQKDd9xm2J5E/FzUuZEDPor9K8EgmUY50u3
t9AZDtvzrrdbKGugCPpHMJBaep1V6t3iB0bqTs+iGgShr6sYwtrPU+XDkauW
8U0OIXvjgB7YL20TmTGNL0Z+5tbOBshfCrnE1T0SZyZSSsCzl49rVXPH6cep
3BQ0Kn051KFLAWX0BJJxVBu/sUqVZ1JO6M+Xa8rSQ0PIreu5TtIpdu9eSGCy
D1oUFz61oMaEeym9gEtftkikDTnnwaDZunW6M1NGbDBbXSgLJj02/WXYg14j
OyEni5kIV68/TiwQQMpkuocUPlRTD5EmG4hGjB3Qvgo/M3IRU1iG4KhKLz76
+GBArpkwDfKBEXSKT7qweMuZy3LzCmBozbaGj1I6r8bW1bIgTHcsGJyJL3Su
cw+lgsSVKDDHNwwGJckSR0nom5vht6cZS5NHFVIBDBtprC3BV25khnmAHxsp
r2rdT7FQ36jXo6RgvJeFGNbFUkyFc/ICusfT9O/FJYcJHbguGKLwllxNV0Ka
vS2lYGdBCTOEmt5ol2/Iu07Q7bMBgxk+5ihYTHtMvWoNqswRCZmFv+kjFoEb
puU4+N9cOUIaPZkLNbyfKgaXKZbJ61ZWhJbLzRrF/JqVMM0C3tl1Kt+isOio
16GmQLYdyLCryDhEiE9Wklv6R9YhHKcDEYxAoSrkxppGr8OcJGMdgheV6b9l
l0J109YGyKtOJJ+nJeFB+NVTWexCYUkg0fjSTWDHeIHpbars8cHaFrhgY/BZ
h0WgLOfsNyOWMmX4v4QnHgXDB8H6MWwmSg4kjCyZW90jCfWHJl8xbU/lxPgs
SMtTdgId0PxXV76eolPSxZVnQGRWNyevK/a6jGrBungdf5n4Ve5fOOVvdm2w
+w4OpkSj76saezXALP4mzYRJbtc5bZlXllWttPizQh0AvCzV9kuR4lQe0x+k
9Tvhy7ii3LlPbVDGiWlQRAKb9O0ArIQQPSCFv420q5+viimf5YJX1OKqc2pE
wfY5YcyoUFGRxFWlV9pJqgcVz9kciiMilMR7DGxrUrrorIjN/BZG8c9/dn4/
4zh8Pk15awOKJshs6y60y8c5GMQghET7UQCmjEhcpk6vLB3jDNSa3o4BioHq
h+J/ZNxHkST7tY4Nx/d/7kvw5Igi7bgx3+jYsHznTiWywJ9kNC3rsOynGTyE
eanMykxH+jP612QAFQfmZUGGvGFez/lUTSWldhioVf1/slEMScV6R4m7Cl5K
yqT/sDSY6BV2Kdtibqh6ZBG/X4DfZt9AHpGS6DhARY5Vdmap32mb2wHCDVQG
t23XVU4OxkmBh2WZxgFfpI7/2euC8+G5E9Q92G4rHv1VNtmndW7IIi/BBU78
6UNrDM5S9DIcyC7WFetZavXs5579VetRr6Bgtp57GZo0BWMfkmunA9WJqFRR
YStSKmaEreSTkSMJ92N9kBq0/n07BNcYxQJ4jDRZ8Th51geJecwge7+v1OTf
RnIUKunENqhyFTxMbUOMzvOonQa0jE6jfosJkLe+G0M68/B6kPecNLflQ/2m
nTUJq/lpgs1aUJJEE9BKoC77ZemAUh/aUHk/yShCLN20XNiqZ8SU5emDAeha
FDRoja64n6t36jYny+xrEVh6FZILMlux1E0s6OkQr3Nykaex+ryYqUIAApNP
Y/hjyl+CyVJYNqzFRCXSBI4Rxyf4wNmyyo184BdgoQFxCtzi0PSQ+SmxXqF+
+YbDolo/iqTH2xXQ130beqdj78X3glm+GOE+pwzzehqcxTl8Zffxsl95J8na
wD7W//yYQtK/oJVaN2iLp1SpHnWRp0/pyB2tR8EZhPtRBaQlx21c8+x1D0wj
boL+hzh+1Ygkc+3RSSQTuOchdjROqa5giaFVgB/RjAJoocgRCmla2Rg44RfO
MZl/Iruq4M51GzUOHKgVEtsAyaEf3h5wu03Ve8uCjJ007TurhGJVT7Yyy4J2
TbbCIwNImbYveD4z9sjmr7jsPhPWfUS+Tw/qknMZon+ijypwLXVXSe4g1D+R
QEG1J8RUpOJU0RpCo6SIq1kmQHBuqF29E0dVIyKPMEyVLTj9pApgpPSrg+KP
A1xl2XcPUwu8HJcLkL1RwF/fQY9C1cD5VFiR5ja0EpS/bfULcBa/B/0yG5zb
fUowiaQeiEadTi0jiEeXebzHuslZ/8H50KcP7VadNeWmkh2wwt1aNXl44Lwr
U38n4jE7OoNGoZhLRC/+QJj6UVxriSVXKA8aXW9/g9SfBHp0mOcZ2+LfsKsH
rXh74VRGqMabxemkCtS15V+qSJPQW8kdd7GNEcAARqP6Id91GNMTmU1AgqJ1
Fqj1Z1RihrEiad13mUcQ1f9wK+60mFIma0cX1wfccaggQXJ5X9vSQaOFpNtx
ey6czyEXPF66Azku5B3ePhRnSJGd6ohYP/TijeuDIprZfCbViQAKhTYmz/T3
snoxl1Tnd3f6QmKuBIHpovhm0xZS1YQX7kGI1qu5ezZB9Yt2kLbLHn8pgfg8
I59TJPcAYC2k454pXAGedTZ/QxHdnpQIswSe+AXsKFGj01mfX/rewvy9MB95
7nGmKub8Dib1DZTvQ3Si2Q8wbQGISw1DOYjG6f+q7kGAvLDLbeihAerAKYL2
Rk8xh6k10jY7+BrlgC4slNdMOzbSKeNXF+Bq4wER2MLgcRT/nBVt0bYbDUwY
a+5wfzZl3/mBcoaRWz/Md17zltocQb60yAQXEbTuxvsN4d1bEGCW1cFPsBwB
7ywJmkkzbp1GOEflJkfKOm+QHkPqzhRa796gSiIngZPqfQhMZVJLK8yUcF0p
94pwmUzcG0NVBB1GgOddf864EZLyMnRtAtJmNng7RcLo3hyFXnRW60am7OkC
2cX+LhtoapWoZZOQcHxiMGhqomKgUeVChgs+yQvOGqibcVFE24nfJUysIi0u
jSwH9aHft388WTXOQ/0pCrV2kYXnxNRIfRS7jQWonVRycSzPPE0cRhw+++5A
8QK1NSCPbsO0/sNu3uGpcMQwbgTfkFwwttfLDZAqeNqkBKqN70iPf9B5L8rY
bbxwo8do9QdampQAallczjQcrFs1V+ch1XalxNJ/yLyK5Ul9EHEY8bFux+Wi
hDahkPpwk4T3E8XxprwjN6KOUyGUkyCJpnZBzX4dKeQYOHa/IcC1i12yhgyF
V7w/anCF4OdiChaL5af6std96ZhgYs2yIQVVjbNSb7tUFx2/bp80TmgHptyv
5hsES618RSGyey5V3r8YJrTQGW+zvfH6iqe+TIyKdL23KQXcdmrGGOsSFZm7
7os4NLMBoyIwVH8nXOEwT1ixI1VfTjby23+ALJsxDYGSPGhs0kqLbiQt2UgA
SrabiAPIEEtPcr01ESUxmBYFbShVDq3vNQPs5zOehF6AhPl+RFeH99bkzI0w
Xbl0t3tk1lXTSyJ5WKHGq/Lcrx72SpWupTuP0zpGwNs7ThaAKX0hLh5dvjiB
VmtZHdzvyxh3v7muKeSCz3ftQsHqACOkS8b0iRRTNJviD644E4x3UIDCHXU6
fDSHkdGlv157oUqF3y2WDM3E5TLCYRneVU14aGm4AMVU0WDaOzRLuB2xV6up
oTTP0OS21yyAWMELvbO0ztpp1mFNjn+Z/lLaZq0BEhLZ7oM7VXmhJwcBGo++
DJNv7DjJoO+oNlFIF1JBYWUMFyNNDOLdxRvy1AK+faPUlRi7jpuJRRT6H6BX
vWPkmJLSDcBwG+Kn/xI338YPIyRQkyn6yUhcogI4MV+x6S+4lLRl3/ZfZVeH
2ZdmgSCz7Oidj7jDR3o+2ks/Ypo6TMAGGPWsNy7voaNAnYq3v3U3WJl+/oBu
Pk044gi9ODsJOX7ZpC/dHthIGC+yTJMgHenYQCVXrHQhooXE7JK1qnG/isgP
9jmJHkpabkUHi90Cb19yKmImP3dq0pryZt3vys9g8f7C0onkHZYLD5zt2YhS
RmR5hbpItvK+xW6gcULWMfOTx6VtbYxJViY/Dqo91WPAdPMK9o/fD+0phB2H
U7F1iSmPiGr0L6/wVyPibfGHnY8UimfzfeqZIYKQ+bWUld+Ivq7rpT3u2OP8
+cS2cc3vq7PIiZaSD106wGEJMvh6KUmCtH/4fWqlY/lMOm541R6ZEvAKL6xL
Ctrnv68H7jHN9OTzfKxJ/ECOKbmIcJm8gIHzUzjUBJK5P4nrO+nYk1TU5lvu
opVzGQYHQdycHxQGDrlCixkTk7PpcaSsCnFHafS5Jg09PHi7blofCsFyQnUv
8q8e+dZgAtu7cIsX30aQDFOqXuSL3H9Co9YH+1uel8RxasewCnp5AmQ87K3m
yIWz2mO6kh13zu1BD/sjmyA1ik0jRdM5sZX1OUMCkDWwEJjsHYV22wbYZVxM
6ZdCHdPCY+l0R/2reQUeUdpkukJjC7poF/z3s/eCr7HbLrWDYN1rUW1yqOqs
cYp7c6K3ihl7LQEGRFlBHSp3JtMcdm9RbYndFU+/AxrWqdfwNExlkC2kqRSZ
tnhEsbcap0NPPU4IXAd/y7rWw45DEfCGBP3RmUlHaKUlsgmsbIJWzdzig9yy
2pxSXSUiNPy7oDbVGYFI5+kiD8GN7rVajUzlYlGc7nadG22yJsKnK8/KXuiZ
y1YAN93X1MQSxRrrNmBbHahj9/exNKIbifipL/gg9vybSlMxYoKuKCzE3dW6
i37yEkEm/9hUdtme6hGgvom6d4hnCUgm69g7PG+maYeBdJDhDehgL2Xa+9Jo
0Q66kLEIBCR2LcQvyhh7KkDDkSDwJi30vQHeFR0r3Mug/XmWOiI36bMnf1oz
xPogGgJ4Yokbn2y9QwtvCLH55lBWdAQI7GK9ScvJEuRNAGxT3qQ9mRjW/Ddj
VvYg3tjYl4hJW5a4JM2ny/fH37BqrrUdzHRRT53JdYC2I1rUCZmQAywBhHdO
eSW/WySy+ftkNMWLrMb5b4h6KR4gRjV5/cXDB8jK+It9Lfpcr+JBQ68+6Sgu
pg7m1s/Rcp5ekYrx/K/YxKHL8EX78cBYeA38okRUuju2uAEkBnHLD5N4r9VB
/xtwjGKzvNDoPC3sXhyxo9gt06bmrtziJnwRYKE7rNjAuuDOvlvimuIZ1nrl
dL5YnmXz0AdzIU2Dx6uxtPa34XBEzI91k/OQ7sA7eoaSwjygThgPuP/+5ii1
8YkDNbHowJNPXhpx3QxIBCdmI0IANCBpua2g0Kmj5dWQzJWVb7zfTCcK1FSB
R0ZMNGXmrbpuL9FK8S4TQ0llswRmrOgtMacYEDRp4eetLDwTp7Xx2WxQ9kgN
bFzSAO4LCEyv/i2anHhKNGIga0BDRmRgUOlZoj9reWZq0RgpmvMvkQbSVqhg
uJ4rOY1c8olFAnD2t6Ko0iA+By3+v6O16Ic/xR40RUBy23l0+81nO2xX+iPW
0mMssfcMr1P5xnjTNJLCQRWD8HsGjjr1agDBVNi7SKtpU7z++iuW/ctKl1Wi
n2cIJwZ2Hy+g9j409guukeA+RfCzRBpTvx7pWPC5Aklu/3D6cszK0+cdDsE3
R8Ld5grv49j9Vy5LoaSuBeR79H1aJ1IADj1ed5XnjMHYm/BpUiuaeZg25k+G
stuXTIRm1++q/X1s0iHXY7PI4T4+2C9CkoGIFGUgzZ/F+Zn1KApn2X+B5lYp
ZHZRmcaYjXF63cpa4LX47CRy4WhwAXjbe09aNG+5EXbZ6n//YauaVGj5pTuK
3zmUYdu2os3qvSKvMNeDW1o4+u0FTm3NXNqXUksXUjXnKbuipxMmFVbd+GYs
emFrjr60TwYa1UO27Ca/NPkaAYFD+7vVwGwxf5xryd7A/+zCMj0fsqSxMUOo
hebjA6FJlVe9uhgGBBdc/f2KhSs5A0slh4uDuBdvFuip44ZH6UwqHAKZx/Cb
fQ2uuhlJudDU7Jkv2arPqBpLKG8ibcYX97WiFVoUEgqsIV5c/3GYpAkQXnwM
jcNoHQiw9AVHWA2+FIBiS9xqeQEvJbXtbPmVbLu+dk5WQrQsXjyp78e09XrE
hNVWiWQ9fGRnU6MI8zV7bvm8tkMbHyM6OIS7Gx/OQc9Ql/zeJHDkZtGPvxTU
2OpgbtN8cFPRjtbpTuDAmoQ2XWlVO6LwctVY3l/FkVclN+lfV6/VV+V9G1VT
xD8Nzc3SAHuCkkd9d0ScXvI5mEHCWiJFPBfXFZ3Eyiqb+LoJBbA892UPTm37
97lLZh4PD82eitGCDjsOyCiSUC4YDezC9LSXh8mhenkks+0gi6qUPCeP2tB+
Oyh9dekrUF/PkQcFVPqirHBeBzMzDR8UPVS45/WfVUiuPOL91B1bNxLzyo0a
HSH3VCd5COm5oksCoDOi0Fs5Q5dpmKPXaNmPunnxUCxeZC4NTv0BTTMzLM2L
hu4eLtBEkSEVGzzYWEo2ScsApBVLP+rG+YZw9GdyqMO7RAeDcUuRRgBZx+44
sIM/7ZPJ+Ld5y7zRJB3AkrkXFnUapSa59o124u665pSWaKsPAJ0j5JKckNF9
Dcov33wr0qhPU8RTAhJZR+vCnT0kTdo3aktKbuI4iqiVvzKdq7wjHcaKFBw/
/CVXNxaPNJWoGjFl4LxhxWXN95tVrY75NmMHKqYgGlCgY3QIoHMJCAVACvZr
9roHyvgpn/iSQzVDAyLw29vh2O0z7DTwgH278z7PitEZ1skpc5ZLpH00/xpu
xaGF9rSn/Epv7f6piC7KbEU9CzywZdmHZDZSUosYJnXLonC9L7MhEBFIc662
gerjmzSo5A4S6prjh9EsTEElHJW5tapK+kdfeuR+lynY/e/2cadc5gDyA1V0
66HNDB1r7p55EzPGsKO3erjI6BcQq+p38yx7dgW+eOWJK3gesXurOhkz7PbQ
D5aLOwBKtpjDKjq/FgAZB1hyZS1Mcl8J621yq2DFyk8ZDc2/ikTs3rWqYkFG
x/0jz5RiNCk5fSikwZUlrl5Klk11luiFC40yJojS0tv+mPfZwnH4Qvu2qTZN
/WJ0Wu0eseza4OCRWgv6mNjwCN42gGJwrUCbOCUNoNynM8hquSHB1zRQyC5x
KaLTb9LTmrEp1YVV8seLk7DiatqPAkVjugYPAPrPcuVJl9iuBnVDSPfhhJVi
XnKffw+QGWldPl7h3mmpQsyaQ8UvwJS5KxaP1YtLsvr0sevJOtfNfmEOxQUk
j75lIdLRyqiGKWXfg5a5pIyA3phvyc3qKhPmZ13tL2keZl1hfk1y9jJXGNk2
1B/cuCAYcZ96Buer/7yB0UgFupVbQLuDsHPkaSlyZT6GjAd3tEBBGzOcZYq6
QCYM2/289ae0BsmZR5RokevvMzwDAo0Apa+5IHr6ZnTQOgbQnuEVb7el6QaN
ZPpnXIq4ZDl+Px5oiAZzAVdkm7QpcRt9y0O1m3EehEAWr/ee7g/ds7IKxIQI
eLuc7dZJBb9162/jXDAiZkxsRXErFmlLfELQORlJJy+x3AEynoBzbojVMFL9
KChg1eD0xSMPtrduRyro5YyaaHV3OczS2an+8UNBpdkAXkh6CcRxx/a7kgzU
5R0dLPz/3sSuymwQEyyjSSq65/jTAGxwYYCpYf6P30K9fbvdVPzwUKar/k1h
cAhyj8+Fg/SAtIDB+U93m/EP8qBDpa/y/Zojo/p7dQndvJte5Dexj5iA8RDI
ZyqHG9IfB5CTGMS7xb0DShW4NTEG9bvEsXQn95/9sjrDUMxlZfGeOJ9Fh5ai
HDUOgHvdtXdBjeASS6xtu88Ragyq4oR0wxM72BP6R4qqCBiM2NIUAT0NPrRc
Z2Gmb1ii/DM5LA8mvCwjiP5DLemjriWEjm/W07JZwUpVHwUppvCtQbMIOTJd
hXNsgrEDCtCbzNcbZ1XDBxK6iMEa/qQMgqfWVLWiNkmUn6H2/nj2t++R1NB8
dAkd7TlGR/HgRMcg1MJW9B1UdwgeaIhkDLJQXnXRKWncGMNM8BMZsvpFE3ON
WUFHUeZaeDsAUmx6zCUyF0K/OtWcMD3MeAzn1J8NUc/5uEFBFarQUmOtophE
DjUfZSHycOs+TWPT8ZTened9zQ6UXA4zf2qff5SDYrLbwR2LMDb2L1BGHpVm
ycGsuj7WdLuXQhd2gt+VTPv4MgYT+addDuvjERSLpgkSchSiQPE8oXkJOZ1C
fgjo66PJNG20GgpgapcVDKVOdFB1viaYspJ7tCdXaq8VeEMLb/BE8YP4MMAu
uyNo5URqqXW6WAt87XjGGQJljh+ciVq8clcmPz7abOn7AWig/GpacZvNb9Dx
gHfHFGmHojR3t3GbWG41U0IT3PuwcW/kB/EaT/AoI+CLKX9ujRyDyJLmHF/v
5uezyIy/SgmQBU7i74cgVyOZo3kY++6iHim82jDaPeqmYYkKYpmukv48+Doc
WobV6Lo7GGSeebxzaShrLeK0eiFNlqPFKJMvslcwzJ0PJeuSa6y0qFnuvTjQ
oEr0TgvEDe1IcIEyQV13mj3Phb+XPsoEiGcLe00P13AARyzGAChYBL4X8sDu
A9YaMKw0FlGRTF66BmO/Y7G16Dz4qIOpY45H276Y4D9LqcOCbSQBjieOHVZO
T2JPXMo8Caxj8CrRQT+68/3kNGpwGYIcAZlkUvqjyeaSCFnibZnOjjLGvnga
JtidjN0XXfmwv50pxR+W+mj8/K/i7IyZU5w06nyDQUELCqkB3qZRxnLS2ygp
x7fWW3vXD5Xr++o10r5aFSwEHg1OEUZr0e1bUHVbwvvzwDr1g+p8hnof/evg
NKH1szHbdKyvSAeugCRl0Pp70Wq+0cVtG/9kJQXLMbQaJvjCMSGu4sJ7AMJL
p4quwCh1HtoyWF8BcOG0/pcWS6KOFQpIt1va+eutmGBYwYiqNO/2FdE7zlBE
F/fC+iUOir4Vvu/wJeRtjGAY2qGYYgQFEbU4K/ccLDgEgVMVGq8ruHzvDBcH
T6WUhBsFIGyGdO2Akd/qriAP2vW2EWMZQizULdcHWMgMGGs0fQKI9WGCoEz4
DLcDASBXQWYKULd4ntIbHUJC9Pg80TGUBF374DTy5vfwPnsP8JSA9dAqquoO
sh4SPzQLoMT+QG3YbmstzK9iHWSXaL0rceicCM5mSqoLigJmTZrbmi3qs6SX
4YXzMkjOm+gAGg3s6Lv1Tn2cCiXfCDQcHfghBn1RswBtw5N4NrBzWB4HmsL/
GnzrMEniZItsCoMVEsD2mRge4gVoy3LiWOvQJRiZrc6p4+1iuAOkIEQpsBED
PEJAqR6vfhV5CIomEbbRkpbXP3ahi2ezJE1hOlnH2bGZopnjlHYTd8dMp1nL
Puuwqbopk7V5r6so52EXVf0Lmqzp35hHEWmzR2qo7RvzjhoDHWm4Khjgmdtg
u94oWHbAxVheKceCADfQ7Sae/Qv6MAuKiBlnDBfEbFbOU7gWjIiyazbk2DTU
BDJLfeuDinlz4OpeJPmpteNcuU0zecE0JaVbpH/qgdshmdyT/qQH5EWv0LI3
CbfXq889+smSCUlI00mltwF5Hk9cvrGhNFKtgd4DB8LZZ9Hun1gNdsF9HKQd
wI0D3/iGYOZ0lkZul82eF1/0H6Dnq/rtG3c7s/gYY/qMU8tUqEF7aVPXzNWV
9RPnMyi3m4b4fZYOBKAI94xDzUkXLO45FIgH11HJIciqZE0VdlpuP95d0Ojj
ogme8Puw+8qhVic5aX8yEVsYIdLhIFAb1m6z09py2aICrs6D/V85zuPgt7Dt
TIu+czywOoFq0Vcd4QIsfCLG/E2OsiPUr3Eld95h714aTvNc8mIqzt1TcNR8
4tcTi10MX4ZCWSPGoak0+H6F0o03OKAYuBXvuIwoht8DmLWuoaulB4h+KaSZ
zjFecRG67HfSb0VQHaTEd0f0wefsCm2ugFVu+WjLc8yo6598zXB2hNNF9DtK
Hsll/w+zSx5/OYGeB3DPhCSq8YzSl0tD6gfitGwhm/aWqwB06sgx4/j+7lEV
3ZbHpfCHZ7vXAU6hU3c3v/VpOTdB1mMgen4Dl7mmu5hA1YFrTzNQ0Lqa0JOH
I0iw3lbg0kUspLpW441sCtIFYUTKl79wOXUt4AEmuOb2Ey/9Hwue+aSwBhmL
mmllDo5+aa5ealWPuRZ43rsEJFim9vMSmbN1edzQ05MwW0V7hd6eN4uv76Z/
O3zx9nX+XcYA7AqCc28if/j3k+zS148Kx5BfpHxdA6NE7m1MeWa1QWpSL8dR
DCfxCJJktT3nhpGjrkA7R1XyLb5wa+/5VpwIjvwTALZEcg+AT5MqeWOHpMPg
arkvUx4na/zNOwvNYpFIwPi2vDEfG9YcIdX8FuhSC4ZvaDkI8TJtNLHFFPGR
dg85OtvpoMbZQPDsq7Plm+GmCqO1sA77o1YIkD2s96opL8Dmzgoq3cG82EeT
dR5mIEqG9JeeW9pS7eqiXGuyhz60xnk2mIjn25ls09pQMyNGCHzn9Oq5smOJ
czhzIJHRwqbjtKrup8RjMiZRs2gqLrkWThajlIrjgV9XZ/Gl30hHfDGZ39qS
ORbUwrL1WHxcNANC10L2rgYt/NHm04qep192bb/FhxNoEWpHML8bf13kVPBA
KRSyVpHf7cKG5yPK3ckYlmsMuQZZll3mhX0KF6bM96DJcraYW2hFFaPp2ROg
TdMSLHae1Zp7pjGznOTHN4ylf0Q1v+QHYmsVB69pWnMkmwL8W4RTIzGxPWWi
xREHdhLWKlZA6N+meqkc4BpJPEHZHB7R2UXK0D2W8xuaHjMENp8R3vlVY20+
KkhyHQaN2ULOMQugqy5BTaFGN+65z/VPSLSdT5EP7pRsm9h+j/A6NpbSU+nm
AUuYV64KjoN7dmN+l95+qKnP14mdGIMqqDYescCzEi5t33yrrJG6cpUjRv5r
ag5zi8f812MEwQMDdicjuE48FNQwZcUzCFQopN/R6ueopgpnBW3jm4JUEWJO
ohNjgyTAeY+FvX+a2UOGpAEIRVVtD8uXSnI+XDtilu3hD5v2EKWya3SAI0Gb
DHcVts2yb2jmnmJthBeY9FXLOYYEZDV3gZRY0doJsEqi+Nif5VFkEmlwKh69
WHlBLXaSTyIcNQNs8oBx4f46SBStsojX9o+UVJJa4uY0aMFudDG6t79HpTHX
VAdF9795AqQYrdeXxSEWsIafD1v2x4g+N3qVblZYO/oXpzk76R5p3dLB/NtP
FczM5eeXqIlGoKOHJPJ+5cB2J4QmohQ9J6YUjcAxHuGdLvhHnavxlxNUIwWR
TlbFSHkawgAnSSrHI9PY7ia+C07HNzePke+8YiRv3/tfY8LAeTbg6o2rWjLs
YUtd1R6Z+GwzHXTYemFLECuTOH0TRq+QSA54sSHB6+As7UO9lckcFyGvTBGt
RfiVmZnP5vLUT+CRAkW+w4PTiynLlI723IDn17J9T2IPKjn7o9CEWwTdwXxw
YmVqPSD/qGq1Ri2TaCzT+9qvPpJjOZ/eVVfbY6+H99j4z0IlnFWPliP2kYdu
rOSuengm54lkQyavV3eH+DhlQAftV+GTRuQDXbMyNDn7PbdTIF6jpzzghIP/
KocdgyicCKQyECDUxVQqacppIvJHsW2n8KhO4tdK9N/EKQl/G1f47ffCB34A
oTCttBfnu5og9RXreyZVxM2USqIzQw/+PnvlZn4kCVyMd+mGja5HDf7YeBrj
BzvXRz6GNJ69GzZ4N4Vp1ajqil762ZQVZ+87bdJvzHML8r6Hv8inkKjrtXri
ibYryGFj2V2ad1QDqTb1E/ML0XzUQBtVGcBxl2DBxeWNYnRp0gbuIb6sOrqs
Y2QESwof7iiS+bWJZYwX2FtQNOP3+B9hcZnKGao/1yJjjcftcvzqtPcFGv3d
hDOy/GFV8/OBfczp/1g7GZQyx9uYxMwRQgAitIqW0BiLOI1i1P4Gyt56+oDY
9qZVuyAynnt/cyqWEpE9Z+0RqAKl62WQkUl6XYoiaTqn1043NjN7zUnal3RO
sKSt2u1lj0x7NZtQMD9HgX2MqPHapvK0uL/ntQ7R5Azp2P+AZFveTAa9j89e
YRk5Vdek5jc+OjFiWpFulW8BV92aU73nzxcAT9c8RruSVDT9CZACW3qJH2cB
Un72/PsmwC+/dYtV/0Dh/2FqnhCABfE2iwSDNLdgAsqLC5oDdLibsQWe6H/u
MCzKZU607r5hqCtiNZIVeVV278MobETgCIv3ApKQbQjRnnh0Q2KucDaXl+U8
dQcQz2FcfTmzB8nZogT0TIv8c48VjAGIWvnCjTdVJKF48577t6MZqCnkV96J
EKwUq6ku/C9gtyrRavjE3NiEklz0WagbAe3eEhhhH4m2gyBvllA/m97SAKAl
TG9DFkqaxXlpHTTxNY+iVudUCJpWpvYoE5iAev10EhBGfdqyrVrRWwj7I/aM
8JkNkYkEZW2Rs1umXwGTswp69P2IT+z/rFVVWoGxUrCFRQIyNb87Jx4U9Ez6
n4bvOlR1An8kcRf+yhotJqI8IHVLMjdyFqSEcVADsl8MjaNhvQWPb0n6YFYN
ZTxKyakQihdoymMGSLsx8hE/Rej2z2I8BNHQ2gbYa/X6goCueWjpf4Opn8Ma
orVeWutq9nZv7l9TjOs5aC8mmm+XQhwNvneOkPDa4Tc0GHOFKPnt0+dWWO+f
xBIjYksdjciyNPO9L5ioqCADNriya6APhCmrcdLsnlXGxEroVe7y6sQE+8tL
gT0Td+3RcLG/f7p8zQ4jUlLyUF18IxTXL7Qpfp65DM9H98uekELDoUpXB9Cq
j9UPcCA/itaNFMtjbtbWWhuEqdt641nCfJ8a/oWaezHZqZqxN/HVoFA3wLkz
HS3XdGzLmRW8YZU8NwZlTVA8GW2Fu0ukn6p3iKriVfFPOg6OOlbhiYi/1GJC
Tc3HdNRht5vZ7TDiGWE2JFMJO70AdoQX7Zm6OCEHKZ/i552B9hrKeb97NZbk
ipVdpYSFJM/xMdUkanG60dk/s/pAbD+mO7D9FfMUohRZ9ElGYC4x8r+pUm5+
L7QPflhxccZ5MevHf1b6rtN9+B8sdx4NQl4C9+REcIrNIS5VaWP5Uct5ZDKr
QRZvbezS7+w2DUOXLvNCxwBdGo/dJEOruP2Uqw9I6jaifnDEl6FSEtta65pI
y+xO3UR82IOgsnZUCjfG+bl4nEVEvbNGvYqvzbQ30L6fTdjsPxinkxkY7O1g
4YpoxkBYGxjRc+EZAbFTqsaeeKmDY+6Lq5L5SPRuhXAqQWHotR5D699m0xxq
TOmZE3QgGrbwsMEEJiVlPFLfYwkI5kYGE6nTOc4HgNTC0wAHWKUj7rrQYAGp
a/zBQIC1YCO0V9O3H5yg6nKe/Rg5mqnwChLWzOrNR+GVcVnj7T9AOzjSdeJQ
pMUPpbYHw0qQ8qrI2cwo3N6n2X3hyOHqt1kLj3WKP/cWcu4XphsjGzF0ZsXU
SfyCR+AOgzKmZNUZ/byvV4AVdMHawbrDZ1cdELThlpX8fifXZZm6t38fR1LF
9J3QLwgVRgLjUb24h5B9Y0YAA3LemeplMHrpznTHuPMTNJ+YZA2eg8DMdAWa
sYErxcCit7MDmN9dBAhW77XpPjJp+s42CRYQcG6WQQwpqOIAKC4lQFypJ4uw
+5xOBccvf8BuMdiBYqN+idu7rqIIZKCo/hwlC4sHz1XNmC/xIYV8byNU4j+5
MMUULWs6FGt8KVfZfbP8RQxJs0BHkknidDsa4qWkzAmijQIHhqpNhAaSbmiU
JfpJr9q7bmVUUdsMuAX3ybJIExzvGK48IMaoLGhlosL6Xwzy/OZ2OSDNkvlq
8d2HKVIxCinGh1qTBgiEdNKYoWS2ATwylHfQv9GOiPGVdgK2YOVt/6rVXAJy
T1nJvx8oAujr7x2JFx7c5MCnFYHZ321t8w2fitEYersjEj1vXYB8iZHW/a35
xn3Nk2ycGPopEEDaR4VkXxRAgDmgWEi3Z9iuY1QXmVziU2KeDhhWs0YHEiI3
sCYBuB2pE4F6/3RZPmpRWzHRwB/hT+c3CAxa+lvkyfkYln2Fro+Ww5YhR/hb
5LmovipFA6Hn8fHCX/ZeFLALI6YvVCCf1BlfFj193OSLpofJHQIHJJFwfrgg
J728G3dJJF0Y1bdLNFMchq7e5CUh50WaynYSXvK2vaRw7s1uJRI1V14RtQ56
bBHMqACJ2VE1Zq5OY9e6+rb3QgyuAfLxqM8W83x29rNdkV0M+V25aDEW8ztI
PhPN43iLrQo8HAWo7gOiD2Hy38Fg89+7C3GSvwRMPeomdBGael5uneKHONOk
YS1mReTioVIXUztb4J61ap6apT4tPG6m+Ki/63Tr0bEcHBx4XqT0ZSgVuTQb
6QsWBRXgtqGn4TbqKGHtqpP0c/6bQ8Sw0sp1b7SUw9PNzZkFW9fy9eiyY+rV
GqP+V2Nu7xq7iOJ527ZHzvoT03mrIhGn/B6mX4zYuBc4Ou83wFB1yWslWSPW
EZWUjJKyJChkTDmHZbBtW/83WTXDfaDn2EYQMuwVonatVHMXOuSefX7IDmqs
6XQu2moQhbpFsmFfVQU7bTolFxPWzoKp16nzjkPAANi6EmzO6hKLaV2cX/Qy
ygu7G+jLmIyuvw7xQnDczRWef1eeEFxAN2d15TEUTRYM6mqQL0Rp4kOIGIuu
mOqcas5qPj7+zwHWa3oRmFHNJLsMgbJ8nlX7RidVrFE4w4WR0ROCbhBRDzC5
EtbJd7g2D5RkQTUA1vt9mpqbPIhVgt5EWuETOhQS0h7s6+xroNFgiYyyI7CA
WvOrX026wC4C85wlgkNVz8ZHdMq9+JZFX+RUD+GgUYgtqbhEZhcaNoEYvGDI
RqQtpBWdkQswUUKfn16UeCINqY0WYusjPmcLdR6Nj450Zem6WkL9Yv7Rd42v
8EXl7FAeerI0OooSQLoCt9aVPDtKzzljdPkLGNDETmpBRzQXzjkVuKvzawXl
he2MwnUvUjaVCub25zIg/uhgdLQrIoeNwZPwpiUfHv2WvDssyv3O5Bwxxr2Z
uSOx6bXqqOTc0RIsQ+x6sxMivazbLb9uadJ1nHx9GjPUCJkKpS6YQ6pwnB+x
/8dKoDqZSxGPdkol0gb9z185fYtTk/FYNN/kY3hR+JsEIh8Jt0sVLHGtu92I
Q2EziPadXcFqUUXQCyx9Y+cZhGgYdVO7Yqsdl5CyOjK8sEzlz2VKQ/wLWHoD
qzclAdbrzQaZfIKLTPViBkx8cI+IfJp4Wx2231u8ZVKQKYqNuF81YyoF8cLI
vrQnbBcgcj1DLI6xNYCSlrUlbfBR5wMJKweNrLIBKBMj4TYxt4Ol11yOdxtW
lqg+NaqI6AygmQg+PxZX+dU/GXpMkXBpRL5SFRpH3NAJzugKJkGdbbO9fUUF
wUA7vTCUqADn/WfmwmNXYWxpR/OS5S/B5tnTDtg/ky3BkaY/mJiHazE0k8+2
E3qNSU+TDPd7yUPAIW72wVoWcy4n8KCyVtHXw1u1pTW40lX5bgAGLG/SELao
AzPT7J6iIFA5CZ0hRFv39azZVkzitGZTrzDF8Voc2Xo9hLSORjzEwAdod3J8
+LKn0rumW9zgMIIpTM6OjRKh6w9YDHJbEzwGLFBA6KzoJtLb5JfTwJb5CQQv
2KSZ+0jFKcZQ+s/Gi2sH0qHfd64GEY/6KejLPmWKoIvcIEAQSL14PWQnS1sy
Inq1+LzFxKUrwR1p+Bn1p4KE4ib+sKDZuKv9Fr205ivAGc+Lrr8oAZdh4qeT
2Bf1tSkzOA9U5o9nRfyQ3zsuN30pJqyEsYL3VsZ0yoOT56OQ6tyXgIBTdFua
D6cAHMOuRSPS7qVhXo+4+uY0fE35hkJKCA5XfS1ReRG/t8WABWJDydmtjUGC
td37Q2eUUab0rIe4Dg+cqXRPi8JBWGtMRZyPKyEQ8m4KeHDY5XFkoaHxzj0M
YtMHXk8OgIkTl92njixN0R8J32eyf/yFrJCGNX5lmIlhMEs9Ri16W3pujAJ1
GYIYty6GGL/LPhI18We0WURKskxgEAtPJoUteos42rGlnq8/nEe+NHhj+Fyp
VQURPCdUhyn3lOFFIrMqA8yhSbWvvpYyEdke3k/AtURsVw3qqhS4zeDSibLG
4bwb67Fb+br4cFwlD8vzboB0Ny+2tKMTrn4CWZBHSRDZmxv5rGnI4t4Kh2h4
KYvMIH82wme3imcxXCtZ6dPNQbY2mqvLuMCidlLe71UujIErBHCqdWCPXdMq
uT/UwFtodG7cDDNSCTZ7rg6MV1wlrPLDU6Axrksa1yHEfEodLxOSSDVt354I
AwSKw6I+OPgyM0ABflescBK/fYBwZWeStqr0zaLVduHXMr89ysdkvi+j8BIY
IROmRWhGrB7S91jHO6iNg7/j6C4US7Vly3Os+rOn0ZPyro3n2s7OOE4/BsWo
Gq4fTXjRpUSTIwkbXMmFdB3sVa6zPKSNsjr/nO17Db6Cg7Db6v7SQBwe8vws
pLu6Kp9BbABvP5wfIpXQuvhnYX0i+Ne7nxgPYDJ8igzojrNmerU19+lMhbJL
OU6bxJhlgKtPdFiazkhyazjJHdqvDhWXEn9m5detpCALZwvOENesvwM/gFqn
mo065bakG0PGrpaXpojlUu0NxDmlgDNxUiab/uhyXYTwcVXY3Y5B4vuu2Ggi
Uyow4l2ABv9oJgJQ7L60bupbcVD/yeV9g63NmdbRQ3vQ9+IqTI6IN6+7HdwJ
7r6ArKBU227tGUXDOy4QpN8GkJQOnS68PmW0MNqEOlkXKay5PoNNEUpWvv4w
3Sz82b2n1itZQ7aWcdaMPifCOJxDCpZ+W3yVhcQp2FQW7U/yZI7yYPI5ou33
0GlS7XA46zZgfmwaLCpLpXPQVd+kzw7H33ND2pUWJC18zZhrEEIpHRMQ/qal
UpMWRVWXnJ/ldmwal1dR67g7yZVoZc9wvfGgYRWoZKFRjKTXY+aF4wa7uECI
EaHFey+nGaFH1KVsSQAUfH5W+7TXSOpWkKyUTg/qdd2x2KQIKUWzoWUaCrLi
vHVwrjmDvn86RbJkFub1c31dtxLs9e9qubR/IBpaXcDNOtuU1RE0PANjbSkq
LsWtevYJb6JeGakpcDzJ9W29ZfAZ9f6CG4shAV0dSG3crj2U3r/Pv7uQM2QY
SEetJnsdnsa+yQ5WWvWaqAe+lJwpmoeD8nhiy0swvu6Gf0Fae55mDPimBI4I
O1RdSTr8DGWAyNcMY9ZhhhMqabwhNXGsURtSzgw9ubrGctqDB//GowE5Y0o6
cJVPAhPAB8Lv7YOFV3UHHzizhFxNKeS68ZQDZMSMg3jUF66/+a+mGW5HWrg8
iom8nwruTlA1/tZW80NQd29AvkVVCYCY+FLO6iDoHl+FQc6X+GbqMmC71+zq
qoakKczD+ChSPtI4dNOJBw49vjlqIMmmqND7rGhYbURgsL7Z3gldYaGHaTCc
PQ813+M2ADrrM3EJ+pSnViop3ewR94Tr12MaI1VdYkbsBrPeS5+j+3vLv6S5
5BJQVO1AHr1p2xCpyxIz9or/f9iT5xHq0DC4xLWjqD4y6cSz0HQWicEoI7fl
Y66Nb8+jsROkr2Zv+Xv3y53mXvqGwZNy7YWqbOqrcwK+sD9nqN/57xF40eSM
yMLXl0MnLLxp4cmkgXbukaTQt75VoAiWvAa5VxvFUmZD6nv2MfOff8yb1QER
5Y1rvWT96HBDXUCaW7oVSt4ooQ+eHEchn5QtcsqRnV0gAeL5eyVtnoqaUv/6
K3/JT2ye9/6zf5URxQM8cD/O2QvvIx1wfwfYEtoCgztkfzJPB1CTYUa5Bgxd
IUcWP6ZmcpFclrs4FkFgQVw4ic3Me3/2kGMX/0mrYId7BS1PEyby+CVBVHKo
LKXcHNhWb5xTeASSloP2Ht8Lf+bBP9CJh+jdOFqrqM8689Kf9rLI+VTdd8o2
Pvti3siLZAx0SdJ8zIJviD3diCaVvhBfavn48ht1QznjkhigNS2PyuhYFO5b
qNhvr2SwdsJJY0WZr1stQBluJovOrbRXDwgtgjOs5Snbu8nZH9YuER9x3vaD
nJWE53RL/dNDyF3GMI7CYnbzVTUQ66OOwnxSOPgT5AjYJVsFtgMEWKLPHHLZ
GcXjMyR2+IOItxKSeqP+hocjWRI9JdkmaotR/Ma2dSbSUfjHdmY6IGOL0w5s
EVsp8Me9kcoePqCXLjCCztLIkFKFsuFoPWQPSrGnYYRI3IJxad9OYzXwoNgI
kYw0NnzMmZQ5nlVC5pjJFUVT4vE/fyRuEhmX4T7+jJ7qhyY5Ty82+fZVgFix
sa9VOVbjCkxo2Jt81jK1pS9AvWjqSdws7mde2r45J9Zo5+GuuqgcbN18nnsd
G0M4jrhYXBF3iM2TD4yUPM2wzKTxtwMZncQIUrY5h33FEvwslxDvhrwf6MGo
rXZBI9kf+KFhuVdPtBNCDTLpV9RqWv/83rvPrmlLjVSqF/fwtUOvTru8H5gi
Xytz1nGOH4gkM5KCuqNbTFemcNHlslBkvsS91Qw3OPOb2lPMah2xol/PbyYQ
SSyd+gpYlZ3diwm+hVe2OMgADlbU9KBrW7lORTc1uAsnfwvnGKev/oT5bpMF
zPdT/UvMq1HsGI8yxPbtCYibcckPdDQSzuOX4YFkTWkq7HwDLo8zOPwaVN9Q
33ZpFZzONO+xbR+K0J+6HlCid6OVOL9ufy6vF/xthzXPoCd0xVnmmmMFcrB+
A9akHVISxAlLSswvfwASbKUa6ofsVdRUMJwEGtp2qtSJQeLPr7a6J99DBzbi
fkSWObEM8WRBmUH7ZNcwa6m3LJWeSsuBXz/oQ5OLdnrh4dKoiRT21u5mTz/a
QDFYGnVjI/NxFHY1GGP5W0QrW8omgh099j4IyEV/1h7rHpMO7vMkt75RH6Md
e0XaEVPtvD58AISXflwmqVAB2HtSWylKk7w24RLjO1DlfC5JGUv5sdanYH01
L7guGc61GKm9naiozjU4R1L+YEQ/R2fUOraFQ1ftL1RIW88n0bYVTrJZCDI9
0IshtiI9Jwb+4zO7HjBxz3r35bFW3T501JWj5M5kiq+7XAOtDLhuz4qG+skL
Dy0jYyj+zspl5eAN1Pfs3fQZN7ZudbrYgTMlEQmcxTMCCcUnWGAEOOgdkust
UEz66488uRIdAFLuKm/5CbjUXvua9h/ORyCcxH0TRGsJlU9kmLk7JvZAqYbe
H58VHVYuQnRFKHL3x5LysKrDsWx74ZmkbdxNofvWkEvQSGAg7CLl8ZNl4Fsa
GurVJd2E0mMgcTf1Unz9VytddMgfJmSxYCFCOreSNSqSyvB/8akBjFE2ofWp
3KnLyENUqhAmO+Z0zkRCqWnNE5xXXe2j8L81jMBXoBao6+Vdo3ztEU1byxen
yBIqZa4aPgr4YMgJd8bqK6826YYYzhyIVeorCB1MMdJ1Ljg8/JC1Dgu6SRRq
GSF7ebHjo3BEN2F3oKIP9psPh0Ele0xsjXFjq0tcej/um1oL+tFmjMT+C7Z9
hFNB0ykYq3u3iurlDGvGB+y/w1wPnhZ9hl2OYxgLM6nRs88JZWw3X1wI/EoS
pmZTujFPH0XYte9ZyLiKYaPVmH3e27k/fOhqugg0Isi5fR9vMv8JxbImCo8K
NZVa8qdN+DoGi5BMmnXRg3SEEEY0+cIKQvXUaPEzbNpZb4ykrKFrB2C1kHim
/tHH8bUot7mRmd9NBAsrHWKJn1Er4Lhu2DAaYDZCd0QF8iCMf+JPHLYqlrcN
Sa69ShFcYOwRuNj7G45rx6aeNfc7usk4wi7YSZ3N6SffKi7djeTN7QyENKyz
poeGxZqk54K2evHX2jcPhMWpmaesTRGn3Sxua6mKAsHCPaQQ4a0shenZgk8X
kZNcgnXLINMMilbosnENouYslTVPvOJNzykzDLi7WHIkdfYHt3HPersyYV4b
oIGHGWhKXWRZ3z7uvNIRbfRlzgr2nCqT5aKdAdAvBgap4yl7/ryni5TNlL7K
3DVkYdhKR1MxBE4IlYz0sK+oc7kk0VmWMyRFExfy4eKtVG1r4R8tZu1vQMcG
7gyn1yz1tIWkaznnW7av9D4WtNjExidRYaOLOvW3HLyG1baxk0UwuN4zowSg
ukehmEJ50sD+Hpbld2fh9SinJjvwQkmzmTfQsq3qsp1nPazW7Vw5jwsg156X
fz7z4hM6+j3DoMHEDFjAxiCxbWz9u+IBb3OkXGAZAPuo2MUlg3v4aM7u8cO9
IO2PBzc880JjI9tMOU3v80sbAUl1alUCVjaUvpibkzHw9nNuTCrCL/A7pYoh
VaAvyOs4z9P+G0PmqkXc0eMxOU0V7p+2btBw0QjgyTn9AyRJLvJFk8F3CNN9
tPuTAcTmt9aKAnssJ47ZNPvB2y0kxJZTZATsIBOGWB8e0PPA3O84u2e+AYLx
muGheIIKzfgTop77Sq9fR6pSZ/NgbE/+Q/BW/psrEWrFkRJs7Ax0GZ10XKso
5D/yiTtlqL4FsLsUZkReckRFcCueJwi/aKbgfEWI/FSvvrM6d/Zc+4lgPHTq
5zQBNqVwFx4xDDkyX96x+XF6Mi/1ukrtRP9Le1pHwjuCaScqV6J6+4L5DktH
cr6p3i4xkYN7bUh1XrFoCOE+UJD9sLga7lkK49QQDKFFQNsubZJFgMBt+Jc7
iIorfSOmea/REASTzmns893sCj0eXYy/C3h/0y4qmK0E/kRTLN4Mdjc014fj
S5c3rvPVZW/0H3U6StfCbaKsMuqas2SOqY+iL/EJE+MgWaFeptIbdd8JdRNk
eD/8jUqMEix530H6AI01R+5TAgiL+e6Jft7apMQ43/bb2Y9dIfOH0ltIEO1b
5aC3Rxq4HEuPPef0XJTlBTtdI1l3wPtNq5SHJamd7Uv6melz1lHGRW82DRtO
n3pDdB1eiCPiDvgoI7qETJHfg6zgEmUtkJI598UIC5f7RCBZILB36bt22JJ9
2jf8QQbe0Rug1zyXZDM/OAwNwC693AJSJPRSf/jaO6QmXK8ZtPavvDXS8KKM
W6d6DnKa+9VDfc3hmo4/qQRDAhfO73k/5J3Bx5APSE3mFZho9ZCy53tfmgar
j4W6l337Z3KepMJjG8mW2YB2MbXMduI4DzhaKrWU7o7jVfTHm0Yq0sdEcHxp
UNUtVPHTo3UbX0S/UKwx6iZx6HAXMiR2VwEYk8ea59WG1c0MdIdDojBTCQBI
zCBCZSdVHn3ujoBz3xTPgTz92yxTD/+1TlYwWFOw+oxE4rH/NM0LyVdq8Z76
lYyP0ySc364i9f8yWG/Cybf9kUEutntKWPSAeghDUDjAVY8EKEj7deWEH0oa
7eCWTdY6lp+nfjYK9dRvJbcyxBo4W4BlwmiYy3v3Z+yj0hSOcyyJsAMZa7Ao
JcQS2IR9MG9Tq2ZEc5tkdZwQ08VWbFyXPfA4+Qpk1a12V+XsudjumdJqaSHs
baRpIzK9/UKEmIkwLUEdgm6c7EPStKhUfQ8EuUrPvGoUbAvRoG3joPrDQIUt
q3Pi2e4Z7oY/ysMjOyY1qWlEAgLeVUIJjy5WWq3vn1c7GJbWe20UIGD6+jUa
MJ5o4AkqYm9y0O7/+P2D32gzQRcewfSAr+TMWHyGiNO7beU7NiczLy1I93lC
yfOj56gURryCxbz2nu1V2YBdxUA+0USiRwDX2D8YZetxSZ6y6w9BgQCcdAcn
g/4ZqaGFvybRb2hK7zQehgu02T0Dj8rXDQrVRJIlHy8jknmZFcC2doEXJPUA
N1JiUKsssESRtWRqozT7PLOSBMs6bj/K9Ul4OWua3BIJyZp9dGh2iTEKMmmJ
L0uszKzfZV9wFZKhNh7t2OdfS8x6uPmiY5ySzwrxzyEkaklLsZbYvBXP/QH5
DFEfMfiBWes2bBCYVCf2u97m5xmNE+mrOuqcrhnQxYeQ3YR5UqNucbpAvSwi
rj35ntrH4hBxy7C4j2Duc+O9iHhSo98LDOKJMnZwhJQUsJiwUTecbugVxu0m
dC2Aws4AX3vTSNOc3AS9WTGsytJ77fRZsPR2p74SITX/drSj/T0QenqEbz0t
E+A6o68lUNlQPyhDud0AL5X6gEhMKoVkdZl15FjfDNMjvNXXV4y9lGq5MZJx
cS+NZPynO5qnwAj4G0KuOUoAcuduhOymCEFmrT5+Pi+asJ/PMDLP/C+DxGok
ychzUmbSHxyfr5qmC1W2nhEJoZ7EqUYmnxzYZ4Qr5/iUUfwk6HXrCjKrUi3j
BjpON++JhvQ6ZTE0pVXMKa9PtXWmHEl+t9npbphthneHc/82+mozymAD4lkr
wQG3hd4QnwsfI7jwQED/Xz9/zylV4qu4C2jv2XvEoGAW+DtwT8BH+Ef06FKG
kyoLB3jpP7tEia6sdeCbW89HmFDszHPhtkSw5AwLwxA2qDnE7uf3dznD6lBD
H4Pvd93ne2u4lfPMjVMupj+jCfisKYjorLKoLRnDrMbQoMr39Lfui+BIo0B1
Thfl84msXj7sn5dRcVsjIX80tZJ4olQGLOZNVhyL7C1rI8L60KqIAlss0DXM
qrHyihNs7Q38cxygj/HMT8oShBYrN0LyEZMc5uR1cFDUIyOI16S48htvdFDx
m18s32TAUgutNcIbyCcV2mSMPfREZujw6dzjSWeAMKzSaMszH+beMsiwSBKA
nXS7XxWORd7BXeTZXgHAspOq5KrNtPqGuVMFq+MV3bJd1BXgGNX7a8wlrpxc
4IlIPTqxq2fTk/+SEU/Zbx9hbWy0DByhPPrgqx8xeqqs0KuegCoxdtBRm7aj
0ymSDkap0GUE0nkj5F71JDNoMHVM2IYldOOD+GfrUqDbQTSUdaGXu4Hr6wxJ
Z97sxIsYBUcY/9gyrTBoP9hYBsAt82Nsr2zpWSXSdfirWIdnCFJl8HI/+Y4p
ufHVJCJnb/NX8LRF2UPokYsWFBaO5hehlNzC1rbJHYHYInDN3q/yJ3FgpcLE
1AFaM1Y+AwdrsPv5LFjs5fs+zvsM7QGBlcdko8jSrZcywhASCkbznbYKLI7Z
2ZlHGRKcDIugKiZQa7nsaglBqViXuvMUYhKPy3FSPnrtyWGPHcJ3JeEZSpf8
YfK/VGZS/hrDT/AADzxuzVJ0odRZlXvdzwu9cJMyK3TVfTaZoMwqrUtsqUw/
WFmyGFpXXo9yD6UKFVECJVaeZbFB2JjTAFTHK/elCgTWlyhPhCt9r6Q5hpKW
nYe9g1dPt6xRuaV3do0OQ3AAg3U9Kj1ZyENhxgJ3Ue9EXTiQ+aoDtbrSc/WC
CWEgUBSvgE20/h0w3grat8lTWMehU83LAlUkGKvm4sA43iDZnSROb8rvuJJX
82quoPuoPVqkqf4Yf9cKCnJMUoassP3BsSjFnZFSr3hrX+iL5F17FttRcAnx
oV6jq7TsiJQO0wkE4xO7GW0XnLfvalSY64I8B0ZLHRKyHHkeB0FlBEkiuxAr
IanvklYKZmqBLFFwEZ6DU4qeebXQ035VsAAzLtpCiwbg7253oW3X7ZwksUH+
HAE6IgLCHnD6pSChXaHK3QkqOA+eGvx6f8WmtRQOx0YlkrWBVUSINxZ13P3p
fUqeYlYq84YWEg5VUxYzDAy+3imvuCunvxV22xH9Srayd2snE8PnuZe8/FrW
U9la1AR0Y8pYO74hvyzD4gz5GiIyYoiv/RTMq6JDtcR39FbjdaLy+TT6wpBW
WUaEfvu7+UWDBcGY4fM095IlhxMyBhna9OntFrSzSK9dHZk+MbU3FQeY0bHF
QIj6iFeJMeaa79ZowHuZNJLG3scgPdiuH9bKj8YO49T9mSK9RZS/7JCqLCvj
hLaK5NwxGgMI09Yu3lLNDK7ESe3Jt4+j3je4JDsUIdaFNLKzhXurBkrFECo3
QhieQLt+mKtdb04jcyj7AG/CVqWcMcqiGERKAMi7x0oDqfx7bVw2EFv6g5Bg
SwuH+q8xIPur3vsl9rXMkqxvJaqqkwCSzL0O5yFFRNqXrRJ9DY7p+8iiQL7x
avvdObd2Ch6p5jgjl1BmCYbuBvAx0mLVPsjgMjDSqScwvVvJYO0cuicJcCyk
Tb9/Vkgl3Z2gk0Fi64fXTFWC81Jji6ibtl2FfU/Y0BPx1fQrRzo+4ATlTLs3
5lE4tZLZeeymtUiwdyzsiVEJKUxNQvOH+4SGthbiCUv7auKa1Ho2dGBjHIgn
H8RYfgnYRXFVRaV8z7+i6u/3rPp8eSPJIibfEQMJfdKFeQbLXHhvhbpUq8UF
z6MAD4aJqV1XbNWtziqq82z9KECJIaVNQqO1TePIoerGolUJnre6cmhAVFnX
rTQ4unNMMSFaKZYhjVwCqaS1wXsngoXfHK6Sg5ecfjyMY29dErvPcXb6tjR2
yI0tmgmvJQEzjurEQMu9ka1tkK2PKM19WMWFiRtwy+iWZmcsH2n8UmNrbrSZ
ZiVyDZQ5dEbjdlscTDAiWRyRI4jFfxgqkwJ1bSX0rF4ok9jebpL+XyYNGsR9
D3EhbCGaK17xiIuiFLANDqtN510EqFvkBeJHsUbaomfghSkwN2vb1NoBwbQ8
ec6NcZmF9hgK8g/18HhYljjwPXiR03N/clnWSOLV8+QyKnjXlS2TvOg6Q0Tc
LOnh61yKiWIPXR55r2HRjloITC7wAlWm/UkkQNgWua5wlefxaxIB6sWqVj5+
lAW8uIcTBKJ4o27lVdEhKlyfqcozmIox8OrkuXCK9qoTMjCAVGlHdjlQXkRz
J5fu+/vhQ9l3V9zhR4YpUWUFowgexe2WrIFp5dtabadq4beWjHpYZjdVCbC3
S0DjW+PQI2N0+9cUwB+CZ1IWIyqy5Mz24A1M6bdyTVCvP02k75HY6LOepkBF
OLpLfLNe/o2ibGt7G9lukGJvSStYHS5chvk+z0Aiwsmjn4GJOax2lj96euvc
EDxpSnk2/frnHm7vVEGC4Iy+Gk2GjhqXt00SWMwWVt0m4CQ1A0ZRk/ttjeZ4
q2mFSkOgs8LSJHQZvdrNDzJLayMzs4xvK92f7VSYmHymp551Shnn8UOpCzKS
QyGHYqUsC9J/YD/7uhY1fTvP14EXTl8YhmLH4xO8AZl0l2kTUSJD1jRyaYvt
FL4WSujNYHYm3Uhr8zfofq9APgaTYli+jJb3fdmVxz0dyTkSGG4JcS+1NSvz
WHWBe6W0eFJVM6QPRQgvAUgSbtR5tSlV5HBnmuN+zkM0eSV/7/5Qnt9ByuQz
cKQSIvU8Rt2ECskGSH6o4pCixtlpzhLVz4pn66iuXhZufiuwY5kKtmESlTSi
jFQZRY1XgTLtcPU1BHHaCOAB9M6CB8oyQWfpb6uACZKtV3b6hD/peN/iK5dA
KyCaGvyMIvFDeg6iPpjjGce6qvEVzl22nWtRy2/z7lj55mOF+K8FKjMRwbaJ
bRnbDZkoobTX2qKtoeC940rGWZ6e97OvburAqllXfGG+BBlKVYt/JR5L7+uj
PO87Zv4EcCnvpXkDHRwYKCCn8+DCFC+GfVQyQckzkR9wwPEKohW3SNdTOJIt
FCUZXNYyRLFNflYSkUaNGM6MDso/zJQGzsbBAhTImTWJRMqo86XdrcVp09h1
arrfft9omtwwpcv57yOuLwEOCGSKg71P63kXV8VNEzGjqgQuD33XWUlPQJc1
K0l6VjodSho8KNTYnKnkasIrHs32kH/ak/ICwms5AZfdCJTIYTW0AKXZz/2G
SvWcEdQfkjO2hcX1o/gOX11CJbsTJqdiisqoVQKtFy/A7vXfFA69g4GYmnbg
mll0Cr+Dwgfl+8q57+6TAqOXNJY+TP6XnDaA44ZHpVgDJRwypFlqrl5vD/a3
unlKy/eCJBVAm6/gaK/BI00TIosfjA/11Vca5elJZvCTUqKPv2xvs1HWXpXg
tAUassqnpYWKXW4GQ99mZp0QS1U/XGWV+UYV32zK72TAp5hy8v3lQ8UAbtp1
XMlNXXpxqnnz0Uhucd5mn7/H4XQaeN/nC+F579pSA0XVMexiu58Hhb3/Lbcq
hGat6Rdzl1/rz0Em8iOJryn4keqECRrubxqY9SNWCUW1i7+/stQFwyZvbv1C
GNJLQop3URSpGLeb0RLzoetCN6JXaLbV5pgMKkfOw6q3Rm2Q1FcRddXF3LDn
H6IE9iOJOvsC+sCFY5oqdFwN0qZ+e+xM/aGBk3T8fEOvYY61MEtxUEd8qVfJ
pMXGxS25xoXLaD1kcHCPV75c5L4AjtBCG2faCmlcy+OYOUyKKjH0wFAvmITt
qkozYCjVj26ZZHZ6JDsnUX/mU2N9wNfcQ01Iv1+adR7swPlhNEOcbeFeATRq
q/841s40LYdQZlTI+bUF+FgQoY5XMtRQwFq9bgwtNuhdh03CZGP6V00EGqbP
zXWe741ENMcYYM+mOfKjVC7WNu1dnkd5NhYgFNsLqYCZxmRHT1xWVSKU00Rp
Hkv6ffwH8BZpzqoXT2SU/44HdcaNhwXA0uGrQIhco4mxUXLWjKdgOUlDM0dO
vPi/6YTOmLJATQb4rha86xPGXC6fLnI2CL1FaYn3G7LRXuV1H1vXhlvbVctV
YkjtjObzy0MO8tojIYWNixldC14CZbAuk+ujXcuBoKdGVtSZugDAE9bOHL0f
nr4MunKnY3D8AkgcwpjrDTOYOfJkINRt3TyXUtzi+7RXca/AR9XxICqTNtW8
4AcDFTv/+2l3U5ULgRj8myXgRPxeH98bKbSCVAkRmLVbmPZ81eAsstdqNQcB
219dVVJWLIq5Hdb1F+F2jrARw8NM4mkaZ9AJ4luLdMdogXbGNyHwOfLheqlH
E2HYCGyQl8ZDI3cTwiw/+6DEJqouIT1vZ9DvwV6D4+2+2wIjPJvTsExFl5tv
npzIAUTbbawQp5JcJo5EW2TBS75FPazcpjrWNbxNTXCh0QmVH+UyoxO4DjM3
f4T9FkEI60XPr87NHw0rFrqqVyFST4e1kZqtqNvu5Qt/ZcugkSLrSJp7Lor+
sphLcHXoX5tRQkq+zoGBucJn70yeQljZ+Q0R6d7GvL3XmX+U5z+SuWNkOlWu
dumzmgjkQIHaQMM89cVxsEQ2bGcDPsYZ0sqKnBZLoSZf5KY2sjSBwUfHcaTR
jqyvCLNuS9Sfyny5S4WKVfNsyQVD+rP9l6iJw6G0tiHv5fK1PkOu3BzAGGTo
snHXKSme0tuerGEHTe0273PyoZstKFcYDubRe/DT1hdIHmb2+K9wEKbMNY8F
mBUwn1yt93h3Mrr+/W8qQix+UXZyAt2Qv7ATzgFnaZ0xn57AMDPqb+D4EfzK
sQo8VhoW9gkJ1sLN/w35HfRpyfIspyLP3lb9zjpALRD0cDCXjbinWLrgdTxj
TqG/cZbli2HeY0BBMchvOFYLeoFVl6vxcIurXa9oN2yMdFOP+QSnsaNqvXC9
elkLg4D4KgPGXl4s+Nc+KvtegIbUnxJZz4Ptyv+msis/op6KDb8MxNolbc1j
vg8b0DQl0MGmfN1jCHGAFhCFAweAE8nyimql3NeYgswe3rWUbMyYXbub4+4Q
FnnOA8BsvmHs3wxekm1/TYBU1t8x5Ko7M2hGo0+/Y+cGf8fRuffSM2/JMocU
QOIdrL2Lf/O0T0WgfEOIx87y0m4mEB/gLZAD2USRtJuU2r1fHPTl/krl4b7B
+0clpH8vvJb3XBCJvWfhcSLC4k1gw8C2e/yQi8lr8z+14dhmxB7RUT8Ww1mF
54dhiQzyhRG+ZaTzYp9AqJ8Z+3VPdy741TKlXmQ9G7Cuzi/LXc0DIl237gIW
BHdLQmcnNILYYBLF6eCbEpfstLNTCfTfFV8HBlAyPqIry2feHNTUOQysplIJ
8YUJH3yluO4B3Uy1LK4Cq1b/ivUo3OrR2239viTtAJ8dt1SAgKjVEJq9pb24
j0TEXxLZ1FbIdH8GZhYcj5KX8UfEfzX4fu9XXQyVbIyr/RKzBLXbuvYVBmm+
wzBws6R4meUX/8Bv3qrryV7UU582LFmRGPjXJleJ8abTOEi+11VVfLvHrZqT
Rs7Djhs2MmyaLYWHtsVS4nr7iwgcWU84uBhMb8tMr5y0r1650GtXeLRmjtZF
/JJv9AKcRcN4XaslF+FJ66jTPVaod2UDxxNIfnIgYp48+czmxQpfnLiD1W6d
0N6Kl3nvFcCTe1GtJaYeHnRth1zHQsjYRVFjcLoXbOmqcym8aimXCiy0EeN6
/vAbzKEusvKZXzvYmewd4K/rNugqaEMDtTNSXqGGxBqyqY3Z4qISzOJqcO2h
lG88eFWZPUohGhYses4cGO6ROWtY16AnMIMAm6Ert3X3JVLfRY+rE55uUwyy
XatYMzCDmhbXa3jF/toxk9so627Zplx4PnTKgidAQ2+M+5txp1E9ru/XyU0F
1v0ZjsH65MXF1KmXMozYN/tXrtgeOkcAskDd9mejY3uJTIlpl1oskFpkFU4S
43XBguabQH+QiheThlHHxDhoNsjvNHK1gZwgQQEoEsEnTBghSeESXtrqFTbO
NQRRzuJbOE77bdiz/2UDm9WfoaA7uP+abQtD1rclXGABEM8kZg9xjxaJ8iEI
Ma5IGo3W1R4r/hxlaYZ31dKe5rGwTVQcSBfpQFlzzt5NjH1UBMEe/tMffBUq
X84RvD4QJElFlxyd4TXty3uMwn6cL+FNFsBSuiwpVpzagYjxfWnNqA9VcMaA
uRUKa0nyeargI/Mf+IVB8kJqiaj94S2d0zZmxcIWkbhtwIuu9XD27sSti2lT
b0cd+mvqmb/HULaPnoNA1mgrTyVYMUiqBiMka6EnM4fMfI8msGcMoZtEB3AK
ILbO9G7DKVYnLAoEGjK0IMzwxQ5s57ZTepSKyoAfm1mgivG13KJuOv3kh6LK
eOUTVJbCuLzilI5PKQTIY8JNGlqUqD4LiPNqbtu4SqpI3Cip6fgPArSjqWbT
lh3pR7mmULRXZitIgivgoGTI1XjdsCAndLoTTN3m0j8NKHzCNibYpqesRnqE
Idgw87ujFGGatxHidSypRs4CHzJFSlRdldtH052l9v0LoRqoN8/QqW6H8T/z
hXlk0++HLubIxTeMyybHle4PtNsOcLYcZGgpQHLTeacB/Ctc0hQQd1a9GLUN
vYuRPKp/jXF3aYfrvV18epdXgqPkoa3NZvPJVOaDUSJWs672jxNsfIyX7wTv
MVMhLlP+bFq+AoJzv4JcH5ipeT5VWER5sKzY7+ZrgeuDjAb7J8YxJ3WPeGSd
vAJ85+jsOE1sbuXBajNFbdV37+WHrfBIXAFlWtqhJTHOApugYLzQN+o8Hkyw
e0B3hrUKqmVd7C/rpuh266SsrRVEgcdjzcNoLsSX48kdzvbzOzNHQrosv4kS
sk0GgAZXeR+FaKNzTwDnXO+dCnii17u/g0WtFuNoW5cl78dmCeADB6o47Tse
sJPP7Q5MowCq3xPPZKd3LKo5GywfjmfspPf8Cd6hG5rX6KoU6edI3UYJZTXZ
3I1HAWrr76SluJLJjN4JoRYUCAZTETtBLft6z9DRouuT88/mMj+G5Csr0mFr
5I3vkqxKkus4exToSc4vKD/Rt2jJhn6ZMzRzK4CUza8wrGw38/dg6+jJYqEd
kFthBWPxzY10iA9FFfxXLCs3KQc18y51vBN0VjbZraPx7ul4C2RTtEqau1ko
msb2iZhm1PNAzdkHFVej7xttQaQgeoFnmtag34Xfh+vXkDUEwtd7Qmy+R/nM
t4PpmFovTH179QkrTuAQNKISC0FeXrVCMZgbF2duSFg/ss8vPIfEcXUIpIHv
Uvd9QrYgsc7IKSVbq3/1XbFcqbii5RhoKkDoaQ+7VpEBv4gb4dApk7TuBCnQ
x3xTdKLh5nvLtBP1z9cmaDfxYDy8LNH7lM7qfv1ybR7nK4kxD121VNHx0ZT3
FX9TzRRN5qv7a3m4gPsFLK8aHLVlILNyXPEXmZctTTvyEx2/cxABbj8wytZP
Z3mKG75eAzAaqftZp/Si0oA5xYPqLlKwSTq/HVux+nfjnBy4y51w0xZ2xSdu
bsRgS/9GDqCctFM/D6b0MciyznupuCWBfYunfoNMJa8KbR8UgmF+MHeMa5/b
50xVW5RSZ4kys1urtFTJcH/bkqYkMVKUctqlsP4JAsaVzAW6QB41YGdX0WaJ
COE4GuDSATnZas4U1+bso6U6MU9nmwSEslvp8/wTY+0heuOjW9l3ribQy+id
hsCyjf4T7tcofVf+aGVbRx9BLEhmYPqSjH09QXwXmVPk7osaaEgHkP59mpgL
kO5wpv/osxQh2XCpb1DiYIJ8y/6+9Y0N0KyTm+5lKDf3YgSloX6pTkJvtleY
cMamv9oPmQvK1P6d/UQWkUY97zrkN7NXsp2votlrWdi+58YWAGY0GCM1lnxu
PdRqeShlVyGfBP9yzt9SFT6C52hp1yJYx9OLCowuoCnno42pK4q0f1hQnZzt
BTq7gBMnmSo8ur38NYGMfZbQkW7k5aPz3EyQG465eyaeJ6UQUzs+8XVtZQsX
Z1lf0fjQmihAS083uf0Wyvas0HbihHKQupD70crh/w/W7M+JqDbH9H2i+zTl
SzMquDctZQsmKukyqaS9zRLn5mczr4jO5agKa7n+dJwGujUvvCutTMVo0fHU
vSZRxVh471er6iI5H9fLTygwQZISo8IyntnriYWMDLArBHM7L0Fb57q+I06l
XSGhtyF6GVkGtEBCF++5RJCFFo63fuEbS34TjwmfdJC366pD9f6HSJhgi71B
FKsqnqU37pJre110pfu1aI7WoO8xEEo5vE62B7CDf5W+OR5abKoGXgFPOuZi
ovHj7iRvWNdQW8GXhmO/Tf2iKyaH2gyw+S6+4pQFH87p185f3iWN3TOPFch9
rjpWcXtkahYW5Vh8jene2R7hTzGfuT8lyAOYJ5acnX31iklr8O0YE9O18qfq
AOItV5yugDy9t/YzNuZ+OVNqEXcCb1KwhF/Hbqi1TYjNHqDytStXpytKv7Xm
6ItPvTSNqycEPr4iYxZ0B3uXDyuy+6+0i5xpDICQaSGJQC/+DvwR65Zstij3
y1qhV1GwpX572wltUiJuSckODFFgBrOG32XuP5zGrc2w1ZLlEabHrMH6kHVj
pZtyJFwkj1Fmq71nnSmNJwqRfrzTOhKtii8vje5OR1fI19Z3RV91gB3lbi3J
CNUVj/XzYLUAl3g7hSsAIYbsBjRiLlZrODRaotsWu5KLVroY3M9rcrlaYmUZ
0fHwURPthsG3INzDygkXzxCR/9dsMJRmyH8TZX2+JcYYfDvS8cwm3jhtEoWX
njsuzP3n3OfyQD420F9KXSVK1LlZGf/ZoBINXRYtqo4s2IJSvTJwuLf1KEiQ
zhQ0+saH/XC4YmNlSFF1nK0dfT3x+fCtFDn27n3a+/bVCIA4faQYbjVKd/tQ
1xP1nArPCUf+AJfo86UBPCw44EXqE+lFjt1xrnVV+QJr/46qLqVa3ZnysZyW
jNqrXNf9htmN1GFsmBewwdwEb1akM0bL9egqDH/j2Taj8m6vDGOT+s+xYPBu
BK9wTP8rxa8URA2mkb9Fo5j3rvppUECwSgTu6KSg719L8lqnm+j/0o1i8EUb
tCUTwcN1cg46GQF0hqfCS5jjej5GNssQtD6OrMMzaCv0WnlK3PJQFZubTJmS
cxDLR0zYte1mL1jr3OSZh8qGrUdcDoel6qn8ZTOD+OPYwfuaMlTtAv/YZnhH
vmbJgceptvZhP+YBHcRKIXivjq3fD+5RNiiiCdhoy6eJs1fiEOufcw5MrxiO
CZDxzL2L0BvP6ZD44jyhcjtPv57IpxSXcYKwKFPYV4yR27HU+eFFym1sl1Qp
+6TidWDYujnP9DAuOJuVsaqvFHzOXbwkZXPwMqGv1BJUaIwdLA5Q514qHWnn
TBIlUs3vb0qQ1sGcHQqk7kiP8ISl2BvF9EeAja9hyouCvkvgP2Nz/O59R5PT
1LV/v3DzdOeIgN5Rmey0fdrR3mCoYdlNHubix9VqWf4cN51080bslOjjq9/5
qM+8XglHCFWxU8kb+z9TMsQ2sovEC2zYVQtJIjhayCtCVJP4R78UZIUbtedK
OzDwhJ3gyakMEl4f/KFVH81+oXIOZSCt74Smq/3EvqyTuqlyTXy2rqEXGrzS
ywCSemmsRfRIq/8fLNQyh996gOPxKu2z+vkPiHmAwdRQWNgkFfb6t0izF/3l
shkBE4Oe1N8Cb/T0EH6ODV35j7yXp+sucIJzr+Y1wB7fMKG1rUliXhOJeal4
Wm02/zby4Rn/bvuHpdZQ9YDIq3It+0aXG19Dpj6VSZfKsV+tzWWWy3AZPeBC
hwwBDeGLoaPesxyYZnOB/3Mi0WlXVf/Bf2yYtKAnGi4eIATlJsohsLISzr+v
AEVtqd9r9hMq4jBRZrfXSP8Izvi2j3DXPXfEbVW3AZaXCCL283UKZI4ecRq7
0bLxlGBpm5FyN5YRR5ezEkCYCyH65Xff+aEC2+r/daiN+hm/B6kBoxRQX21Q
CeCVtj1Q75L5FbViqNrE0ApCzlQtszi5ktYzJ1ptmOv/U3ZT0VEtHt5A+GGH
lOuPtBItOHc8x5qhXOt12VIvd0tl1UUeNmH4ZNYESWIIG5Lty1kAAShomx8X
jI99ju9eOMfaEXQ9D0dIMloJNEMdmfhrmuYHNp4QN+p74kJG7FnVWb2eMAQ7
l/glP1SDs9VmoP1SeMTDDvmaHxt6bQKcmxKe41ZRzE0DD//R4ha1JmyprAD6
y418lvyOuZMURPOyq4VacXrjnAb1RePEGwwf89NrfmUlJSDxOmrktFj/c6JW
6rkx7cQ/CiCsF3rBHpU3GnPrpofaF5JVsCYMEf0ll0Fn7HeHrd/g2UteZGnf
loy2FzBlRUVKnSPfb/WLfsxH7LUJuxBPFTUrmAIb2igBJxVLJJjWMWnnzkVm
6dgQ8jJjcL4CQ95XFHMAOn+sdBK1L+pW2HMpcKSPlSDW206edIs1CvgdHWTg
Q3V7uPANvol8FGGvllzP1Eqnil7WvXr9skg5SZg97ZvJ31HtTog152uuJGJs
zRGQz24fe8ttoPhw/sTOlsN6wHX6x7KM2ViTqoQl+fo3q0bhCE/s7RPqDzNy
eIjzKrjJggZICPDeDf16MRedZJYJ4Rw+eH7JLhLS5LbKxsBfuXaEBIS+A0YP
Z0VnjyezZQYkJnFtndKh1+YLGObkjqgkeut3I1xM51aR2ZZ66IKFhMw9VvHc
avJia+zPI1MD701GJz7jNB3phCyyrhrk259M7Ny8SKVaDEBOruf4mKDRssF4
ZjIXaodPFg2KJXFiHpb6EBppnU7hW+JwJqZC8N+x+7WSPW5oDO/encv3UnBt
N/rfIQ9wDnCqqUHY+Hql3Pl0fzRWbltaMQyfDVP17KMCtDdT9jpX2iXQD/AH
VeGkzGd00KQxSzhzOVb4sfikNX2/L2IFy5l2s2p1MelaJGqj6hmXA+BC4nrw
HHF4r6uH3uvCG7CNXk1rZEO5Jp78CnKcQYuIhA/Xbbddjeb8IeFoakWHiFfS
iBLPlKg8m6J4zBTCaSo4A4x7ZT62LZ0bb55g4nMm+J238VwbFm3l6m/fLxtK
cu7Fs0ToRP/9u6YUaXUb1OZFoWBT1D5Z0H0bAV8Jc+WplVtVKCkT4l+ozBkH
8Uou5YBjZSd3FfX7j21l2G+e15eXRlRidwoOVywqQO8mms7nKZbk7N32JBn9
ftcKhfKPEadweZ2s5KL+yueAJqSR0iEigwv0NkFzR6IXaL3bI4vU+Q6kzUPV
WFdEnnM/8pW8iw5atwDEVe1KmmPOsGqRR8rrHEYXaP0XyU/WobV6UXvKPD+f
zHci+0q87+1yrg5+qyEr8+aQLNk9C6S7T/7QlqKduq6r1r0In/sExMLm0hri
v/B4MXlo97GDxISHHaJqFh793pNbE50AeABK7SZLtjkLqrgkrrz7FCpIaG51
XMHkFvFC34saPZ/kWToULvbSMfT2hwpYXP9sUVnt7SKhWVQjFEZiSFof2avt
cMLsQ+qPlFN5sqpQE9V72+hbfKHf5kaik7rYu8Wj0fHc/ksBZ2fjlCvp2BZX
zQFMZuMmeRW4fSyJSyzxNF/hq1kHG10zbQsSCcmySYdxDg1SFNH0WUuIYkgV
nVqvKAj4K7zDn7NPiCqSuDdn8huC5fcBq0t37dpeY4wncUg1cJbDzTI+k6Bk
R2z1Gsyh/wYeC0xw9SRD91PhrQNR+0t++B2bnvTmUWExPat5FaWlI1YZhusm
GZ7n6kPzh1sErbeU83StcrZkq/TSm/dtfZ+euNbDeCOt3wndxb1N6VAFSbyj
AOP/ru6oJTRwSbTrI7v2m8XVOdA0UNdkjixtR8KcEaI5Py6rYaPR63DA0ON3
YB3B9/coJ5u7+FpbVJUk/lBAj/hhCey0wRrdPuZDMbHpVi6GVOlwL+nToeOU
GPXwY7YS81OUW0aK8tkdIJkx9JC+NT6vz4pa0RGCFhAts8R4/r+HBIGlMzaZ
pi98M9qoWdy3LeBz4uIOGzq5MTbON57Ucg5lNHb/Hsn6b8n4es+kLtB/Ml+R
rP5JK7UIQPG+ZYRWnP0st7pJvJ3Rscy34EYISlFm5nw/EQ0ex1k4TsWDmuSy
QQtDEPi6DwicX61zn4dTb2v2lE2CNYQKdQYSf0GTCjP61zcQvwi3IDrZMo5M
D8loPoMASG1uLTJ93/7XH2dA+MXkftWFjReH0himd2Lny86s4UugcWYj1wGX
I7AwQODJJpLMlI5Xtzrk/FBTvVM+gxwD4Hm6SrlhzcSTDH/+WU4NOTNuF9zX
kL7epSOcUBPsqwgCswdibK2cI6p6qS7JxRYn1EQiYTAtRgUmkkP0FvuFrwDp
rUv2dG9vtfSOn7JB29GLmVuZ6HV2dDxOe4zodgGUG3OjilvQ0AIXqk4i6WJY
96qVwa9fCRXUjFnoSUvrZe7mXihBAwZ5VwK4dmNHmmw8RNHtCUQrojfe8Ehf
AAkV6uXLOLcuVYMDFKDrg/DHr1f3SRQGusbywx5XfrvM9ZUg1Sv/5Fdk57oS
WeAVRID3amVb4bT2kY9M9QMJ/OoSISXdju4U9vspgm6bk4QZ6vXVDaeUv2kn
34CNewVLA1wKpv6q3WbfJuW7ywFTqF4AbkFcsBnjhjp/H4MLXie6tYpsVH8k
q+l5CIcf14Ole3vYGwpXCGdVvOCx6e0m1IZH1sOz3AXXBnHwgTv/YJ0Vgywb
KUHlfLd9GF+5P3biV52Gbe9O+z24sXi+2ORedr3b3hQeRGC3wDqHAIKSzlnU
s7PLLbzNH6K3Z621ZBcelDslK9eMgMjF46+79qFnDlqfzrJjgS9JaY2CTOaD
qVb4dzgkDlC0Pzz/xHD9kynlnuO3rZtUYpF68Bh7rNwOFgS6vZciINbNwF+X
hJYjTU2H08SfdJfI+7nVstvdMkC5VBa6l+Y0AEkez8eEEkO0OEBLVGYbc8G8
JGYUPYb3ERnzky9Jy+kNhyOHZkNLlZnmnzUEjDZD0msLhrrvU41Dskmxvcw/
VIVvFORI96Lq+zUl3G4I9NaLyjcxJy6YRrrTkoPDzN7jfVKe4VqwOKqEXOd+
3b8Hx81eokupLY1bYbGNZlU/khOxXZgqEDcRjG3hQAenyAZUr6R+Ncpf9GtB
OR0DFahmKVBkvyuOV/xAk9xr49EGWAfDqkrjtMsYLgKQHhjlDCY7NVt4AnVu
KUZijGI6iFy75OLgtKoGVmvR1crPZ3GI9Lhr/jQg1CFdlCSR/AeVuy5a8nat
YAqR2+dWTAUEXojMHZu0yV8N0254OcPo8zvJywVyyLu4fMSvCPcQrtKM5nLB
rTJGcNq79/meuwft5ccqhRpiQuKxLD5egYNEpNMGsGqlEjWD6kTNWnIGBTJs
jMu3sdR+ZywoU8heCMdor3xhUr1TSyD8CdpA4guvP2w5QfeYj8oaZVUd0zJc
7urkOUbdJ7TjAGUJ5JOJ7QoPmZ4oYkHc0zDWyuSpIprYiAqFDSFDaivSoan+
PNEid9b5AHneOePjDfSB/KcMTJviVw+tWREgrAOuZwMLNRli9BzOO8W5N+Zh
C8dKIdTJ4NXbZy4BlRZhHxkoamDiFJIHQHyyIJecc+v3IGlSlg0fMuj5Jgrk
u4ZsQOH7F+ToQIb40a1DOBOJoLCp7kE4xqM8AXI5OxnSSaPJ0npu694ZY2dv
PcuRE7iP6T6rtZd0OQZfL54nXLJ74YFtaVzu+50Bi7UHCMGAnYINNtkOqzxk
UgwDw4JWGlIMqOHbYU2dXQ87pKvwjzzVOZq6/DMJYzcDTm9vwgdZyRdTZkg6
8npIFEPpbq6Qi/aXFrLa0Mso3y7SQ7iCyxKCug+uqJDVBYNkVnRuQGXB9ZA8
/+7jUhfURW4VQ9tvr6RFY0Ewg8Joc6dghBBr5iJwBhEzc/igK8t4ykftblNn
g+BF0MhXxuKfzMkW9l3EdIbdAuZetKwNmWCw5uvLeAVoEv5xt/+60p+rQBVC
xU8gBy7vUw3q4OIiB6HKuIZ9pQEQVF/G9nBcBxEIzKxZHKfJh0q4t+JX6wUY
cx5K1yhHGZAJTA8IJwbUzic6m5gxkARu7+C6Z/JLw1K4H+Xqqo02YbdpvIep
HEs6ip4fYuc5jWzJUaoQ/aDNL796+cpdcOAnsqdERko2sE/v3DcK5NFrJF8f
E2UYfhSYfUnFHvclDsBOAbgQew2aaAyyMOv53W/Z4l5dvhSJNrBNLkXL0PlJ
Zu9S4H1KoUnZjW9D9DCKeoVKTSiTGtgkXa08oO2Q25wXGdgT7yfn4rX5byZJ
1CcqG0SmKGAkF9z8KdB7h6Fw8wsFJgyN5FkPgUQBtc7Y1u49sNKXPFbmY3sD
+kx6vAN1gh4Tf3WvPyR7sRRoNFyeW0BW9PfG7MKlrzoLdU0xOAzYCgJ68QMf
PB5Nld8GaGe7TRQ+K8YYwiuc0CQaqxE498O7aaaq0PanZVJ0frVLNTWbhF1N
1SfXyhni/krVJlZAlZu6cgucsPy/kWlD1z2Ur5JXOrsXhd5hBBYmkAM/ZLh4
05kXMRXYO8obEilHDlE3RqbqgSwO7BN8dKpG7iCp87iHkgE+BGOg5ivoT7ea
EL0My0wCLEwWzizjA2dTwRaMxVeJa8VQKZwAeH5WlE1k5+Qe0p/YnLhkxqcH
xiiozRH9lKnZ+GnFln5GpcWp+a2sU49zrpQzzlKFxmabm1eIgmUhoGlSWw9R
l439E86VJdftlCjXtoIy+F4L0/0+cEQ+wCWp5npkQiSGULewYIEPTZVbLBva
hnsLNaGV6DCiTQiN7nigTsMYaqwUhsiVfziUYRx0OgdjUp2Khhxky6/vLF7o
6tL+wy0+1gajSkOZy2e985pzu+YVih3XLFlAvwRZa1qSMHE91eJRXD7juQCH
wJpYLN1yDv1Yc+dJdn3HR+ssd4TysSCeeCK4PlwmEapqG3xnwwFiLbtx02mJ
+ZsUyHRqZh8GIxR2VN8ZoQvAEmBw5WaC8ODj9ushJcmo1bK92MkCVz6tLOUS
ILOf2ZU3c3meP8dTFUmkPFukN4AKFncvY7qqqOM8yuZilhpNpE1JkEZp8SHS
Om5BOyJyRZxZLl6AAtnw02ZIby1ov7ZTEHYPdAYvh8ShtTm8HwdjXS+BgZvf
aMeWzsiHttEtljaeNpGQK08AT1VohIGH7KwXwaI5pP0jQdLkndxG+V1FG4zs
QIHRv32/JbgHEL9NNIiaUm5WXTX97qWQACszdP46vS74+M3yMUKuPP1Ctusl
7cfEJj7dTGkef5DPal/rQWVbaI10OAG3LKT2dQ8L+EAFxoaxiNMeSyEINkrO
bDwMQMz/qfLrhz4NGnz3xhEx1n1Rocn+zMcTVxJN6YVLwpyHLUlCkSCg8HCy
2Te3ulzS0OF5impDJ7FZ0UNLzvvN8QoxrETB/mfky191a1JDr0i5IpzoQVCm
sSrxYIwV8WY2rOX5KEB0zGTb2hCnwIITAWkuEdk+4Lo2VuIYjRsMJibp6gzs
wfUhuij0+JwMcfg2Wimv7EGelpDAWDK6sAxVJC0QC1BUXhCV/DR1/iDJ8tFl
ztAMJqUzzGiOnCgyGtviE0b4pY2eo1g6pp3xW61xEk6GQu22Owj5jHGSVCzT
c+FLxrwFpSRh+qKcvH1FAP/eqlnqDCFiPLP01YwGfsGpxXvXOaRHFxc72tQN
B+XelrXtVUXk4CeThIMirwdbLpGvjP2zNAeMg8NhvFuW/c6G1H9euaeLsH4K
+NShXaN6fDK82NxyF37y6iRNq1MPKYk7EIxtesrrFT0TEpDrSi++ZaCw1d0t
YqfcF2Wh2F7pf4GIgZQT2l+ZMHKCAfTiWDbeO2JMaa98s3bYDL/2AcWic8Or
dYmf7IO9t9Qa1MSVRYytk3296P6XcKYQ9olOFf2BbNQ/OH11OOydvh+jEu5G
HJ4YCPYBTp+JHE3qOdUK/ZoMu+KT/KYpFZ/6Try75M0f/6PDRiI2sIyLdFyb
IuRPdagIjzXmdTizpcUEhOfoKF9O5AxRdgd1+JRxbL6JCec9V2JtVOQgh/Mr
hvwyAwbLlbSEJr5kP+sE/0cKrKPWjVcYiogq+BZJfURKHaHehA653w3r3hqq
tnDs44eNuXs+11JqrTR44ChPH87zP008QCbuvbHZ4QojWRFKx/Y7pzbue7t2
+Ts+RPitxwzjBpfgsa6cAYymCqfoYkD1QZzIFbZJ94ZOV1xh7NaYvxDuVTBe
WYvT4kfM/H91pCoI+ije3S4EiFQIb/YTzHrUwrqRmK7hDOmwKhnjDWdJEzQJ
2+VkkrW5Qp4TFDqBvRTIx9Cgh8KhvBRzbBGNz8jmaJM/5lxhFdz/n/TEGGEJ
2wc7lu8xMNzsH4H1IGh+z8KIHHGTuf6KocXHyVRmO9z2QEJHOQxuMhboFypu
8DJNQpHEYZLfIr9a4ceIEsJgLSom43NUQly+QwowV38k/2UqdlF3NJehfwte
uIhfnIh6s2eNFRjPh2khOonlMHhz3Tv3Tw1XX9H6Bfeg6PpiEFrHL8PfsvwS
uwHS6XEWlqJy0hamEro9eUH7OtPTV7Gx3K4ej6hcoHFjLll30aUzuiX61OOx
yutljobCQ2Vdg8yAOCZwUXuTKDGs+sNz8um5WOJi/x+ROYWXLaa/7schzwgu
CT3PQZmaj+s7wVPoMCbzsgaadlLU4QzPGDX992LJxWnIQ+7wP0a7YD3abG9t
FYN9S7OF/Trm8p36feyaxa1WWZrtDRFjYPE6TDMTMokpKvEaWTDPEeCeZ9Kr
NGb4hxAOHRkCvzKPYmxF8OCqULNxTdPP7REXIHrJxcP1ki/fSAbD0GMiCxSs
loO3B+jYQ4+mRkD76Zt3CDQtsTX7nJxwEyCDZJEjY1KuM+jwAoSc3xZa0OIm
Ylj2qIR93CWL4A/FzlzJWkBaTGWfOBoWOYwzOG0+PT7AC6izAW2bwrkg/ZJs
ODwRAPh52wZhukVY4omZ/6kGXZJl+NxnnHSpw+/tM1d+wSj+iCOxTBly6L/D
k/M/dWK+sZBSmX8UvUA50y8X9RmXoIEg8ZFueK3Uzq2oXTf5m19nyeVe9Yd2
R5K5x9fyPJVTH79/Yu9Gj2MbE51k1sZsRms6YBWFSwNjEELN7UYQxF9icUxA
F4U/4Df48PTeenMWkF5CAuzv/XrF28ehjHlxkbd3oPTgEnMDTuZ1/uWcjzIC
8sqPbxd7IriUEzQTeUaz+gOdFvWBnAa7ANMjjTczEQW32cylcOr8a40DKWYX
mPP8vgNvv/reKLqTu1R+QV/Me2avTzjqccmN7P1T7//51JAAINYHGi1rUBNZ
wfVidEusCfjiMIz5cvBzDaOaCXUFz8cNDQo1j8XJw51RIi1C/1wwdiGvc/QO
irNlTln/5VDrVVvPebzUVFGoC/4/1ANy5G9X9ygChjfxLB2vbbV8J/7PICG7
VgsbiTqMRlt1ye0HxFZwdgtEybzsNUQ6BTiLeB10C873Z3dWlxYN/F5yO+ec
JdPU/EjTghzxefQWJ4nMYcGnSfaA5wzn5v76QtwxBqhNsCv2ybWfL/V1APJu
epvBxj7vfd/wwKZn8UfsQbRNfnWAwPqXywuQDZTBjZopy/NHyee3rh5OHQzv
ZeGTRvlivTF6Tf18dqJAxB9fXZbEGWcTbY+apyYEmTimk2u+Q1M5yzyCLzBu
msWhnqLFreE5sWBs11H7fIeNaljGKv5dyIJRmkLxrXG9AT9AEsQFWhfD4NVo
cvT/vAm2U1nClaeUHRMc7+7VhfJu4GpH5guVSuDZVMX/slUOAQ6Yw93jLqAg
dQtsKKhBQFaHbsHQlvUS5MVg2SvuYLv0IHnOU88an1p2hNACCXi93Im8N9ZV
UR05m4GyT1Oy3RZbIE5I1Tf6Px0rcUzxfti4G7BQjiYpH5Ch3ER4QT+KU3YP
y0kwicETOQDoFxHOvARE/Psvz0bHVPLOmZG+oWyvik+8CPnI8wu1AHlyYxuN
Wd+0ijSc/KLVaIfS3PhUiWpEAFZp5vOONR+oilhfnRQhTsFqLGDrfHlC8X7K
WKkgQX+qqHlHitMyxTwd3aw5dn3rgHbsUEfuJJwgEK0sz4dzts632v43dyny
nmz8OUL9m2/NshKqMpnb1rVeF8t1mJTYOdyNTBVFULPsLhW6ppq0grEo7XNZ
TQqYnysTsNX7OEKXCHv7fk4uzK0YoQa+eFBcnleHbPDqg10nJS/jQljBM2DX
N/YuocSakNRILvYvfVAyE7kEmybTrUKvDH3VmLtyZChKLQPcfpiMrxtwaeHN
F0JPcpfN7PnOKwornjLmIMhJaCIIkm2E/SWfd6Hfaif1rV4zLHpfPEit+ypR
y8A75fcak/piPwv2n+pXk+vFpNUMcNYd8sWPQb4NB5r5kjGG5WqKeKfThGCg
KFOZJ5S7IBz63dXpO8cNZJcA5jJ5GvT51+OhvvLrXlz0U1W/KmOcBH3Fg7rZ
BBubiDUeAbW0OtQRVzaAV76BNZ+tTvw4yxPKPnKLEIOEt8w5yXn8hmsctSmM
UJRV7AxtydUJB4TmFRFXs8r62o1FvcW5Wk+EGgG3zNHKDAFsLmUVvgvuMemi
/SPnPiVxwO+5+MPA//jk8Rtn/cGhedmEi0Im2nVyv1LHPc7TEu9AiXCxcBpd
V5wn7PhHoheRtoyqNCwM9fwSdUwqCcVWpNkic/4Mpxkb4KKH/w6zi7RW2d5e
e185bxJ2P2757qnHmqZdDd6YVLZHHaazc8SQPYT7B9lw+isjUnPlPkTCQm+2
7/crfu56lTgEFlmSK9y1KNZiPDY7jfHd6R/rMhAbDvchwjfOrPpaBuF+r34/
pC7G2Q5EnR5TYiJNBb/GxVkpjNG6ir2F5v/7Azl3VEAA/muzFnRs7uORThEB
/4aw5F1b13uas833da91xLgd8kGww0g2IDCJndxyMaentTfd8kOC2dIJy9hi
zWWQrWvQJh5P+g/iunJju7YgnfHa2iiqICxrYVHWyWRwALustZjuqLt23UXs
HrGU0ycPKzl1Tqno+r04sfXntFm0stq0xdUp5oTuORexFJSaTl/EqknADn3O
hiJHU+ZXIwEYhOcfqPhDXh+tnY6i80F2Cd7lrCaT4ZijUaC9UtKP/nFQ8xqO
6YfK/2L/DdS6R7ktiKlAy42PqQxHG/5CcxOa4UDJi0cWs8kmgSHINw7G9CuK
Y2sWFtlz3zJsqQ5wcasgrcpVHIdnCUirZdB+fquNyhDlUGcV9ZauS5CIPvs5
KcP0aT0mCeMC40bZI7089gnpIAD3aJQAa6GtOYN+9UYOS5iKZZjWhkxVNLEh
D8tMeN84HDHepURN6V3vRyUUY84DKQx95nzaYU/wKuFDAAlc1J/5q7Mvpnaa
AXhVbT7wUNiidY6XeGe3bY2Pot+NLKINIVmQWjYBzt2D57moxJAGc6pI/9mQ
wg3YoHkjVNh9ZDjNYEsU8RC1nOMvOKYt+hV1rM006olE9vvdpKuSb6bNvC+O
xYcrTgsN65RLlLrupVgKJjiGRkPrZBw9wIFGBhzHT/3PYVtb0IStD3tu4GKj
R5O7BTMD4OTMkZVJokT6iABxFq8FKSaLLzvnKPOlb1pKOgLzO3Pd7+bKRja8
X48ZF52W+fzL9n6v6dXswahUnszOf0SVLox64gJdW4b5162VWZpBYFPG6hbV
1xzjFCDN2PIBfIw9Nw5Wb7kSupS++muaybE99aQJVskTPsMdt5GzBQh3CnM2
yJeHLBiAAijj67ycVWqIGl1lgcstNsYPLh8MMDfypwV0D4yRHhojJh4jRBOY
d+h7zjyq70HOO39G2WQ3ot1JzqYOtjCGBv1pNV9J4kAQ2Y+n5dcXBVnIyQDU
ALuWxaaSzyZJn6moUfV3rihv6mLrBArdMwix6Vthqq2x+tb24hGaK9ChDDmL
KaA+C7ofinUhEV6vRlBkSKX0Dl9ZVW4WNmkEPgr9PjpG3xazuU7Cec+I5IJ4
QzrX9f9aM3WXZQF7zHp8T/AreE9gWcOe59mM2gZeHi25ylAdYn4wUn5bY7Wo
xnzL/2E2CPEZcfgOY+4EUjUGoH3W9um0hj2Zb82VUogDvmDflmaUfEGpn1uX
uQHfcAfzMdq+Qpxbq9YLoNTjJfY5wBd800DJ3UYD4J0tPONfZJk/FoWyA9Td
DSXZKV1TQc43uSGZkPY/cEmWZSEnx56iBO0uaFt5xpsfDoiyyVuXGTYq9iCU
QJerzY4DMTZ3L2nOsdzQbR+8OQ6sul7LBNtuy9SdDUxzlN9KAGMQCoNgU9cS
gibOx2qEaJVTqHV0HOY0ZKilJ3ToTfuFVUBK7PVSuZc7If+YDIWKUM98pHWu
vgqTJcrl+eenkaFoCb0geYPcR3EfMstuNrNcqCmk3al0ZJEFFVoU783j3tei
pZ4wCrtrPjQKsLFIQuB/6hXWpZOedkGlVQo7XJIklblCfOwROFR/5Je6gp/y
oXvepkF9jh5Mb957EeUFf5MDmz834wn0QZzHwRohw4gm17UCpZN+S7YUrlPt
/UBc1GUuD1YzmWeYksQHDA9R+LfqQWxj7yg/D5ZrBLHXB4BniuJuBDgfAi6B
bonkmer+MVN6PSbc4RQXjBSHcPNVArIIo6YVOOKJs/EUZjz05XIcOzgjfh67
FplUyeqVtNIKfes7el06zAa3Ql/rOC6GMqygC2kVQRqCbh/+1vZ5BC3WWA4p
GnGt2OA8j32O5qb8v5Ljd6PTeizeKz4J0Pyh+M1EGWPvUncrYGrmMsGwN+sO
nhnpb0rDOFGJGsRHSZguGn9Ww1UiE8bMctUVvv9txkUa5AQOOcz59XrU8Nc8
DF5rhZejhvCzwxLXmKIIytMV03cgk2RPyDqe5c1ImwwbfHNrbK4D9XP7UpQk
5DtFAZZfHKzJgDKb85VecMMUBuIdf/Tjx+H//bbFRmwbVuyucMxpxPFYm0PR
CrfPKAMqgux9uHexTsERz2druCOuky5W+hMHTXitFDkLFuuProBmTknSvvLJ
qYgxqq1Viw2jqCl4rI0TMQzOSIm1JTFyvXKQ2Whks0v5zgCTQV2s+3kEOXFX
Q8woREr8lzOUbdlA7dE/U3kwtaoG5oGcgxgIMkgwwzpu+dBdyX7Bw21iQ8z/
3FE7eToU4TpQcdwrJx4BpXiAkzBqE6vBcuQvMTm7ntJAxA5zeSRtzwCn70UD
7V9kNRaZlWkXNyE9CZl6vw1uuuq3iei3Wpp4GdCpUEA2TCvFRVbYru6jCO3i
9wxGZl22TIq7SiOs1DMLA0nsQfUHTvnSWTAfGVLKiV+blpNBmouPC2/76Mte
SiN3ICSSaZ/9qXhHnCtAqbFNFcObXHGzHj8uY0fxeyCiu9fy8i5Ey1y+XrCZ
WOeyEHvc+tsH9FWi2anhhQJaU0/D6fJ03lYklE7WqUcIVeayHaHekDHb+qo/
pBz6Dq0RbDKiU5QQfSBHcihFRecl65/cjlnxleM2EkdIBjC9WqzOjczCAjpA
3nhfytd3PMUcs7joBBCfhIkdJjPF2L0837J/zyKv9vRptBS/K4q+nEuuLsOc
sXFJ2Z7+p7As2TbTL7tGPM9OjBhgvqqiwIRbVCcvBk90q0NiimLVjtNat0Z8
1FN091OGw29buWfcmIZfUZqY4qI+kQY3C4zdMXbfCJ4VjN35C+tk2SFD0FgF
QmwkswmrTNAVf1j046Mh9I4neFiVerfqVGPm591jXYKa5znEx79+krBx3fya
LZAzf7DD1/vmo5ZBM8tntlTIlGgBbwFGpg4CD+qO6LpNrVhlXXmmm6XBh4Ng
iI2asdxYU82Who/LPz7NddLQspVURuYKV3XMAIq7Kpz9+FEQ7BF43kDKfqCv
roRdd8L+D7dID45t0Spm4iu5vYTG0K1zPrM86fXpVAv+oe3jWa9yQzCRQigf
96Y9FPEOiMii1CI+SJF7OvD0eB5U+2yhSL7MjKJw5UtilL2/EbqpDJMTMszE
sCGISJPVUe7LXfkdmmlJdpoGEix0OAayvJiPZuVKiXvopbJJ4aLHiLM5ib2a
VdZAR6H2t6ZGTJR+YUjNiV1y+32FTyYkwXO4fheUqdxsXjmFPzjnXbQhrMFg
WieFUgWJxIa9RBljmeCx9e/FddFWPlx4XPpZexZzB2ze7Gv42j0HtRmF72UC
qVve9+3tKqCuM8PNmxAmBVT4A+CtPr/ps4xAvvs7cdmDha/1sIa4q9Znk0en
I6Dr1Byi67o6NnQ4SmEETQ9fF8rUqShUcQCsm6Myb5kKcJni2d95TyaE1r17
mTnUePsDyOEW2aaxNsSNFWUgpLu4jnVCvJGIxRncKzb34NUA3+sLDrwK87wD
LT9kTep92eUzxiKWd/cM3i1nu6n8DBCPSIEs27u5Dd+9toZrME4QSfAAOwDe
lIFw8tiU4xZV8hPcPTz1OcfF8+5URIBpQLwtuHz6iZfmi8Ee0z4BJHsxz8S2
5VwMJTmKOtebDKVJlECg3yt+erh3L7Llt31ie1oVcQKQPYugIP3zNL4pJhCm
+BYCiAFcpecJ85f8eLrIEeQAGTXvvgh3ChbE2XELb6oFxkdk92odp5mSgkGY
UPT30Tc7jGqm+tOOP9R0r1ZrjI3+ngB98OceNchJYnsTXSX0ZhW4G7ASf1Tp
1nuo1oZDeSvq2tGCLkamyoVA7uJ4585oTg8h3kpZvhXGz81tycL6rxM70tn+
TyhY7eNvGgi/rj8P7n0kkNOW00CGvrrXDpZJFW8QR4mE2rumk33xwAp6Y3VE
mojJ4lMlT5lle9B9wDWqGZ9GTtRU5HJqyv3kqIa69g9vWVWxLmVVBz6t/cnh
oHOpWCmIRR1bZa61bIoRNJx7RHVWPj1Qq+9n+BY2KXFGOYFv5Yt7jIY7sRxj
RxwEj4JKCYyV3YtJYh+QMPXto55Z30fErXEXlIcmli0Pj8oPiDobJ1u7PiJA
oSBYY/OxQ1MJKAoJg2lyLVRCYZr9kZm8Dcv39tfaNm5n7kqgqhkFC2sARMzx
P2x3DvH6GAWOEmKO7JSKpWrlR5XsduNyJQst1qKrnGLJBoqv6ejKC9hh1eQs
kWgaE587Xj49/VntGiPSkxFYRaYPd2BtsKKc8jvbfG6KEpobi+f4Y0hus2Tc
uxt7oJ6rfx7UOwGIW1a6lRKWCdQSmg4lCP7Jh+OaxollD5mSI8HSJtQwcPpp
2l4ZNHwpjfpZ4E8XEuizE1otY8MCw411YnPm+Y8akcJMyD2rP3TjXjpboF7K
USM0mrJvkm+8CgdrfDzvzmcu60sFuzixEO94wcrn/3YlsBPu3ZMdxw3dP4UI
/bqs0S2NkfwP3qKC6bS4qhQg3UJg/iyNMb6N5ADq7iSNLhd3h2Mz7nMsinyc
6xpaCXX17f5SCJ1ZyYnDWqCHmKZfBKsTIIBhiy6IucS/Ne18W/Sfw40y0ALU
5kVEDloHiIYrQuplUN852Mt+2mNGAt0rfspJzIQC7nOumQ0s7+SdrZ9aYwBP
xG9KQejPZ6Y8HgFvFj3q8Vrkqy876LFVQz53yaux6ParMHEfaPhKfFrcyHFd
sERd2f5oY0nhPUAKoSCqgxnL136FaWtnMaQOfnu+8taCYjMXe+zedl+b/OMx
GcSmzUxafpmRjEowF1N2wyL4RnDS9bqlHkIKu7CjB5IE2pWlFDHS92Ij7gT3
wKPktKMxs2sdK/Ov/93hyunJEymmG1eTU16bRPLmFm7yte/PEB6ss4vvshh5
EVd53vhJKQ1bGKPRSVPdsxha4xFpoc6qtYy/wH4iGN3CmT6DHYifKw8YHdWH
wNtanzuXClp/s2pUh7P5cfe+NCeKtnmPpLSVDqZCRNRNgK1/3fggDx/2Xo1w
r5IjlCCyJX4oOMCT80IUFpJSvB+pYnOvi5rbvUL4uW7dIo1mk/Pe5MDB9Ojh
l3QrWKnABu2M6A6j8QxCX9zoT5r5ulIdlgYKjTTBSAloW8uI+4OV2Ckka7yy
ZsUJ1BhAglpGq3i4XmeDdAvlJuOOqhi7EGenHeLNF0Vz/h5FmJQ3Zv7CL9zu
UcjkN4FtY5e7OBGbUvbRSENtjME9Z8kUfr7IpWkgODuUFMhkm9fbaFIQmSiM
ZuXeJv2JMAg0SevMS51S+2WmuhqHBk+9JHXbt7PcyRh6pDimL2hC/3HoT4nt
IsahhOEOsfrWIyGu7SLaNnwYpmEr+/+a+CaOYuAO65GQm2AksB+IRErUngUL
B/7Pu9kflxi1gvxiLVlNFNVJIYnOcFHZO10BjJ5Xa1QdeH+gjW0Qz22I3oPn
vnZxCOK3OruSnL9apeXigWPRaqSVVFpzMaVkS/PSMTYz4TUmMY+xYo8w1kGF
u9/PdM3ZxjbFE9yx0AvSjS8xS+ETU8felpp1XXcR1mL4V2aBaNRgiDcsairf
VsqLkpcFmvrRCCeMuTLtZhDJ7mCOUtaH4yDzGXkJPWE3yOBgHT5GL5RqDZFQ
v+Trt2RGpa+vdLWJAvNlGsGm9PHOe0mTnHFZ0pBp1kHexjWWpA7H3JdbtP/U
g1jLKkhzy3ZPcm1L6wK0GfRhO/RVk1w+0CvSZdSKivVkgbipVgHYjj74winL
nNBaXQK9b+TeeTa3OkJZmzU7Z0RydDZo5tBf3L6CvV4Na2BX1v5Jp3UamO4L
2TkBUj4fzzmqau5yZhJDGR6xJGsvuhT5C2x83gSItRtkd2vHaOTu+xexRY4m
WiKp7mImjPF+ZruyNtPCy8cZqLLv5PFA2+xCaBGDIKPnVcIYeehRj8r8NIqs
NcVkYqAyYKss4/CcyAn+LnL+E0bHfJSoK99fcH2uettgGL2/JOF4KEiknv9K
ux0I+2G5d8srBr9Mjuomnv4SCE5KpAFYswrCTP+/u5++166qGJGzG+qjZc1H
OmyCTVwvehrhHJxqvYsOzaQ0kTFSZ5GY7Kh7CGnxxrPjFK7cKamDDtQQAVNO
A8LDTHOYVu/SpOtWAdvdZzlv5GICBcPyv536l3aiXzE367dZonWRuL0wgVzN
dmLdlZu6aQpJW004wvSL0xhnq1UER+nnElQGkYSVZ8F2LrWa6bSlcImNd5gA
nbP5vP+UisLqClcQvMrkzdK4CvGYnOPKQh8HL7gU9Qxsu9HIjicowOAWhBuz
hohZk4bipRD7h5TlvYx5ntMXf7PtLqi6CwCA+xWZtGM9aB2YiswtYaOoYTFu
grKTwBr3SRorR0t49SIJMsoczagImO57aO6LYnNHR1jC9aaRfbrvAoIXRMk5
Dpk26bo5FLSngEtBHrQ7HDkQIJjuMsSfxrHep/QYFxhpcBeYh46FLPI2hzGr
QFZQOvQJWMck13R+2KMdN4pKx6FLRPYm2jL7WzkpUXDd3UQOqDHL6kaU7Tg8
bGuRCyRAU1fd7octz9Iodt/3RVvXQtjptSDx7RkGXAAQ3pw+TVKOCrYnnRQg
YlHyrTUhHs3jciCVMRq7c/sSS1/KJDUBxgpWcO0b0oODV7yoebmOGZ+Pdep2
/AWGyzs7rFhTLAdDSK/HxwjxUhD3//O7CGDWtBQXXWPkikflLtMmFM0CCtjZ
xTrkLIqhX42RQRd4IFmEtYOTiPOMsI21EwezBTPIYy15KPHAiKdN9sRgbdMB
5DXS9FE1zcVceaYH4e7Aq8IwpcYvF4gbqpGLFjxZh75NhoyqmPjBlICycd/x
QIOQt+UilVM38wcFOSBvJdgGInKijKWvXuNBjhqI+GFfTZzVsvMQc4t/ABFk
KH1aIH1v46aVXnbS8WDy4BeXpuPsGWM2tTPY8lXydv903oM+OVRqrqte0CUK
Z5NI5xj+P+6/0FwvDWcJBccGheZY6MWZigTqkwkAyDEX1QyS5efz/OqXZdB7
BQzqX4pXYUMJlOM3BX0etArHJuUQ+AGrLPSR0/t9/9VCQHqyA8NVNS4sA1nX
Jy/sFZk8Kwtcvkr1A4Ko4jxdbaXYWcIK0IWPw1N1EPh8UdfNuUbCmDGcosOE
Sh3+cJTCm+qr8yoi4+Zw3Fq3xbn4fqIy9rWxsc91JKlhV0OTV75SpeMbaPLX
83AMi+LOfR74kirdQ4ifN7Y3Z1p4xmPTCnval/G5GP2KUJlatwCc0ype3ev5
5Aceoc7JJcCL7PQ1jAGgggyqtrWtGfDJvYu8L5lP76YFUn5M/ldkup36c0AN
bRIn6H4eGu5I2yGCJNM/js5GYEZGi0mI2yGTys0V/QR94CJ2RLTi3PwCO6JM
Unjud3mk2fwXJd4USIvX7V87yZIw76Ld3Dpu17T/apBljJe1T4ilrzPEfLX3
JWbtuOWEiaN3NC3xc0MDCEUbdkDKJanIVXqXN1KlDD1mfx+I7Lc3OeW9OdZb
ew7n27FyydeQLf71lZlhsvLCW2VqXXbMQv0YH7P5Qy2jpCwhCSAjhMEcEmnV
kd0s6zBQ+yuj+W20MbFQDk+dtf5i5uMY77oT4lCybzMG8zA4r6gyYPYWmrld
U9dwyo83TfDJA6kZd2Bt7yzB5/WTkLqmh8vGTb8ArxfwPlRSOwHr60AReVt5
zbLplQCFVHu+cpM69cGy1GJiN1t81f4D44bethjooG3QXxnbAUBdN/sIMm8q
YWetxezaHmJDaH1tdWErpYlVI9jReQv8a+52dlGZqkde0+PfUPjYJC+Baubi
3adEYTN5j3ok3Y0MinlmtIQuYVFwwkOWABSpNSUzOCDU7R9kn3YipK9gARQ/
LBRo6WfqkR/CyTssUwC0Naycjpn9nUtnj/yBX9VZWL9oXAgJtfbFgBycMSam
4goeVAtGnLHzeiw0xh0h/IfUxgqHcLBEYz16rwq4HfQ5NTJogXVxWTvMrlN5
o7wiUA0sTHqYYOgAgjx1hanBdxevEknaYukEPrNXDtmXlm8LNy0JkPnXl8om
YXG/SFltg+6tfVZjHIUrvwFK+7myN7gAc+MNZTD6fGPsZt7kciy1dxxVNkI1
wTFo0RQ995mRaiw1I7vQWq9X/WQNpu5R1Sy7C09MLJholaBeOybWFnrx3oVg
wZlkFmniOXw7tDzB/2FUAxjeJ3w7KiIsnxQLoypKaKWOdtnZnozXotw5aDUi
tLPwxnFWd2NGITdikMJs2PBTA23k8wbrhuMtfNixLzOhcS+GW5Q9htR08eAZ
D8DhSMJc9rSK6iDHpE1J7ZJkl6Lcg9oOA6wYwlVOy8DlGSMhmJPdn0HsZ4PT
Kgm5Lfm7QxK29cN2djkrrg9W4K/+cjtl/BlAL5adGq98i8jhyZ7WGQdR00QK
srQBuu2SKjujQmOgvZPF23bvj0cGHZVmPVZM8+0UvRJgbXbeq/Uz7M6Tlrcc
NCyAJLjD1RuAEjQ+Xqwn/OGuqLyuyIRTYFyuVZiEZQ5nRtDXUoGQNtNLWy6h
/PXmpMBOW8q8gdbIj6QamuknWdsR6THrKE9kOjfU0sOjF0wp3A4X/5uHtiE4
bAlzdABHySx9giWYS1dOdnNw591Sk8yl1Escm+Zz79OVIQyPLn2pDc+M41tL
mgO2G1FC0uVmvlm4o3m+KIYppWsvsXE6JyKD4qM5+q4fydkFjyKS1Zjh52ir
W1Qi+yvri3PcYK4HHw/EHBBGgFARp59C9SqxkaEECC7cn76SKQ4huaH7NtyN
FA1OxNUo5rwENcpv7j8UOVqGwWg0wHoufNZJ7x5FRshVJMWyxQPPI2HwvmQa
t17cFlOkKOZ1+rSLtSwCus/PMlDS3P3/R7CESgCHOacw1Pi3vTSR7heVy4E0
iRQsqFKD979hkuWVxq04mpRDMQYba6SkcI1ZQjqLQSTHhfxGpQ2hw4wyBytv
dfU6PX4xYEbCpeMuymtC/OkBmHFnMoU0yroJWDEHu0F5jL9dDXOzW/QwKrsj
TL5572yNItpDu2KE/Fv0+Vtt/crfLwi/vxQfENseWrIQHZ9F95w/yti3uTTB
02bpgBwCG119txiu2Etx1tqks9zXJex2CvXsB0JdjTPnuJtK67gBYBjyoOrz
chl2BaeI3X3Ru+KtW2zcO2ti27f3RmI3eRZiizW0iJzLbXYuDyavdksY6AtJ
CH6gMrFXdXv+GviJWzEjLWJnxApBUqc9c9pr2KYS/EgpbF9M/I4l+GcWKpA6
zG/YhV+Z8WvXhe1HGVLC0hi2cr5yKZjx5z2BOVhn9WAweORg0g169GLOou6u
SPyguBhFx1Ood31+xkpu2LBkj/Fald4XMBnltBD+xIXQSb479Jt0iTpF/Cde
mYsTvQT958QNsN7Dh0g6DesUC4zGPQF0pQgcScUojxIrZkN8ZANllILopzva
toGbr+edUP9gchCH/N/YjoUnbFBB1/aH/ZA9P+HEUtWS1ULpUz5OHMEnYnNs
Bg1lYj7yip9HoiRXxtZOA0HwvzrlOcyKiFHeoZoZcYHhgqaNYS4e0QB0AsF4
Scnl1zahM3r9YwRp/fToEOUF1WA2hwHMjFKZczHBzh7jHIscFSOdKL4J2Yke
yjpnsS2n+DZNmIsYEDVnjqPt5BNM2lJHIbseaexfFxJ7LL+xvv7Wv96gTRuT
fG28+Ug/773WsorUTlN2HOiPst9/8ZOntXJwg+AB/sO7YuV3pyuLYA+PoKQb
qtv/5HMeQkvwO/3bV3zFjKGfC4OV6VjK/JT+j3+QIrf/L3yJ4v2quiD9Z5Z4
kCmU/t3shzdkKu9pTjhYKhvlExyWPpuoMPzjJbue1iEYg1i8/Yd+Oh9wfXRU
c7V7txk+Nfd/ajIMDZyMtDUfGstH80vaVNiYh2JglfVivIHgqYs8KYj+Gt6M
LyoAOA2cj/l0qsyPb88+o9zEdzQ5DymH7cW3IBCm0U1787/BMs5SLI3BFUYx
7GdSORqYuHpXuAu131zt0Pn0OyjwYZzDAKEssvd1AfvZazDzvRLN5ji8mbGh
fh4HI+/ywzZwAX2DY+vGmNJg/DtKotHX0Y5/KIpdnLvfVEa70Do41Xh+rgC/
dTea/Zbwg+qjagk3XYZz7btlLs3ZNlFCJebFytuchxpUkoP65zRV2PX+4FIY
0hBfwsWIUHZ/jYYyxyehDA99CFJpMkANDx40K7+g/eVAf/OlxiAS2Ri6UXve
j3JEuIQgsr2u7dUi4fYXLZv0nzS95eOD66ZXP9cU8NrzcikginMhnD4ZqBv1
JW5N3twv9W+8//pSe7HKBFhdMc6bCnney/KZIxoztMn26/utM+JaTh6xNtpE
ue6Z1LkVWh7qFRfgLvU0HBW3h7MGLUuHy2YYIcMbA3ldF43PSJydb/UYnikh
j2PSpsXbnjXSh+muW7IFVTbsvSiJ5ioPAIvPMgDp6G20J7cP05FPRg9dpUAt
+nIpuLkeoseLprEv7jGpjys1BRtYA/tAbZVeZm8Hu779pwoky1icJlgTXvCm
VR7iIJ6Dy4KbCAvIQA3ZV4/SMF1SMc6KP7MzRLqqUsMptY+/z93T9fy8zihE
0DwecAVki7zFEeX3Hfu2g6cvmeqCwZP8OutPgWR5o5qy9Pimq1PCHIETzUxv
cL01f4jzAdT9V3Vdrj+QqwQTcx6l0UIVwctLPO1c4jcLO2uCmkiVSagjAnn7
jAM9OPolAJjzU/o0mFjqgpf7qmreCQ3uI9jQkziidREk/Gx48tT+FqvttzLE
YctyHRte0OuqSY/uv5qZAs/nWvZkvAIAMbPMr4NU+A8TtWQYaHj9CUc+lbPu
Qu+6U8yvdx4Bjey17MucZkuecyFQXny1xnd2mSOWhzNAXFvmbGxPXgqYJ93j
hDapC288Ryz7QDGZwfXB++xPrBHI5pmBAKxrZ/lcpbyHlIqU/fyH0A/aKEeT
V9LBOGu/NOdmhPg1L0R0UAE2NoI90UjY68G6e38WniomZCY7LAtOubcq5cXa
gVbKzsmby9GL1K5RXQENVg2PCRl68jGMKqZ0JCVWiI/KYpjkZf7k52XJX5LE
GmIOF0dl/Pq5McrqpX9U9F2qIqzaIWHay9rOkCJ1s1e6+YJVMEFq0+knWcid
/FfNUBhRBNG/rcuD0CJ1UV9539NRnH803e5baAnxS8CvzIOqG2qAXuhOpg+S
IgZA8unLN6FPQyIiD+Hiyrpbc4Y6obegRDn8KlJ2b+rU02yvnwLdXDpy3nR2
e6pguWCNcywWf3qv6mpKu+8w2GXBHw5oeaVo4d/ltsIdAdfE9Zko1YQ8syGm
EzSUuJVTyULe2iu+CbKBB/dT450A/YprHkvr0SyQdVYUnuM1PGAYo4smbRDd
0Uf8kYVyUDKt8mKjoTHqBIOEbfi2y/4q946fLLJz70pOkzTMWg8FLIw/KUlk
w1Z/RJuvfPMB62bFljL9SESr0zFddOP9UoSINn6VrTRjW2wFfsQQpCpUCAeM
mJRtC0fxPSxhU4GXteVzFd3hQ9mGYZuetEEM8HGUbrfWfJjtGfG/2HhkBk6N
4/GCRrjPMt60ZabbV8az+aesu6pogpzzztauCTf1XONt23lSGuEVtbuhvTFl
rUNzN4kWaoLkD3m2kf7HiM86U8wVl74cbv4a879GXKvUp0ly1b8PYaFixZIf
b2d0iJKsdjBzV533P5tmOY+b/nrRpr07aJ9kjdP+RLDKvTFNx309QkB5QBZ0
QD3Y8u7oomBlmy6FaAZwDVhGc+psk1WTeptVTq8yeY0iQx9RTf5+HYman2Hq
gfbB6wmVELA7dXAFCA3sL50atGTl3ZXr3n6dCWVSktxQeu52iN0ZpHC9sYC/
heZirVQEJPcSfrZHNlZRxP0OliofhL9529YBzQ517QgItVAn/FH2GRrFb3Tn
CXG3W7AOqP0LJoMhmz5kr5a32HsG5xPqiF3SRPfytz0rBJJaFUMZcVoHEoP4
QPQQHXFG29rwH7RawziDS6Cmqzk7y4bUasU60WCzrsde9ZXnACI/HDJpBHhO
o1u5bwEzNLGF8CxMyvCz5t8WDFTdFtIM/hySkgouLl0tGyuoSrkKENgSOJ8+
U4zkqraS3/ShXQ8Med4Q5feUELqLzJlOMO9Xd2AMCXKGgddvnA2aSYyV8oqj
gI7bCOZPPWvJgmsFYwVKtTbOqIz5dDrXwqbXgGftQBubEyGO639PCwlbpnDr
4boCAdcgqxUyHuizhQ4oVwZcUr54INpGFnDO0gSJ/t3RVs1zBIeqqNUv/jEJ
7sqk3XsMjYc/9xtB42SFWw1mfsK7jI6UZV6ReihqE/ybmeYFiErkTah+rhba
0Xq2LKrxaRuSQDh6eMVuEArlrThJsYOOZ9J7AMNhNy1VSHlnWS27TpnJvRDV
KMT+suhLXpyg8MjlqtQdxUNUsTGuhMqsq9UjMCw/3T81sGGOeRBmw4nFfvAP
fMjlHuPKFXqPgbmq/+YesKaCYRIDaeI23r5drrHzjNa+oCBTG65lLBtrJZOK
MiRqRCqsrTnvRUAUIRRaV2eAUTLl+EnVBy+DTPMWDQPYvNmyRsGeEAcxLJfx
rl95io6Kgzq7og03cEc66gKcX3ZKcMLgN6/8jf+s5t7vvwBO7uXxfWFfz6Hm
RkXLvqiyHV6GB3kae4QAZ6XJTP99d1LJhTN/kklx/MzmYxr9OkhXB7+iX5Q1
mbEN2YTbZZUtLks5k5ftaTAQbI3GoLxadVboaUeuVl9SUxLDTTwKuCOpp1qC
TlRD0GPwIiy6Rc7pxFQQrfuaOPQcPvFK1T5lSLfwqRfmPE1ya/27YNhy196K
fS4A4ONGL1l5/Oee5j3TvyPryRg3m+ps7Bv1k5aUcGIGakFZ/gwmtmLTl4CV
zPz/QcVjCg1V6Dr+feMa1KbvoCfC5czLl2LgdznWVJn0awReOnqIjYS8rB2B
i93YI/qbc+ZmHf34b4MV9XfCcaatBvu5bNyMyDzngf2jOeiuA9qx7+6I0UY8
HbdHYp4z+1XZqsmfkhr93T4Uz1ZsWARH229iHmCvQAWO3Gw7Op1u34q8Xdst
pe6Wa71Zb9kigUQkRWpXKKBDxp+lPPM0h4AwRbPAxyb7k4hA0W818QZZL536
dIV1OElDPjvwRPUckMBVheSbiqGyUxM5Mra7ZircBFRuSUMH81a92k8hSK5V
7kV0tSN+Rw2hX41WZYcEHCcwgHuk7FnXd1cUQm2PcjMlk1GFVFE4kSnfr7D5
tV7EdbtUUek9+Kh8wB5L2FKjLyw5mfzOWwZ0I1RIkk+a18e0loYAyijm4BDA
xDS/HafkRs0M9R06f3dqNINIov/0xOGPDilRpnU9HATynwFFk/dkqkmzmuP1
c10R4JuoJIvmQCU8YRFeOCcFH1C33VRkLt5yoAMIVrqy89/n+1IjROIdDkA2
7/QzIa2Hg9a9QEoiY7vQTnKjz3QQMYG7TZSmD0VgmNI7IjLR8rNIzyemZoCm
kN7hTvoy/7oo21eb4uMPEz06DXuw/0zLhG/isF+sYPTE7cKaRKOW4c49kcqH
wigCRQ2eJXDkG8mCHkQsw5eSg3mgHELcXsKT3H9Jjxr8l/IR698C2DpytFn2
QAGk6td9qX3GQaRBICsQC7Unx6EWmHJvyqlA9LFOc45kKydG5DMM+tN1qFrZ
AzFE3mtx8n0YD32Wbt8pdfpHxn97XJdfrNgIZPHgFAPr3l7BVZEZ2JsVmh3n
2QTkbnmuezlIaAJ/R4ScY9GHbNBu/TC4yJZJc6WgvURWWbty4Fu6VoQ814Ir
AOALGwtPzaojvwxe6PnIDw1SWQ8DLJCIu7Jw2N+xqyZ2qGS7cpvt2tVqy8F7
aVKXN9VSXmQy19lSsAMg8J68028KG/A91LwxDC8umFZuoH0fdkvdPXmpYcWT
POMvizmGZ9H6GfghpA+pD6Y1CpBPb0pjfgWsbRgSAadWzRm2SdyX1K7zr2ip
iFf8MF3lyrNpkuXtaarOTfNSe4ligl6RROA8j5qkZNz0BdnZ1bSGo2RSPlF4
3NrCfhSURXUYSioD+/VbKJ1oJ5A6/0qjtgpqoL55Nm0c6ooLxvK7QeiLdiLL
S5gA9fEawqsLv5hlKdbbqAmk8daZjitsxC0AjHnjL1+lZNS+I9ALgKcW16qD
NIhuJbKhrSuAMAvkx6ClRY22Ad5qgWjXlfSvvm9b8P0WcwVtcd4W1BCuCmA9
5i3GsJkAbBVnia+Jr50mPFiKas1m4Mzu4TLXv+RIRTA2emhm2wfnQuWJJuhR
D7Jemtlvp+3y7S9FfXq4gYMRGC4LqXq7Nb+stOuzo5VMFqnDn/1HBniZEp7q
mQa3PrODDUUGlEyC3EF5w8rIcqEWFwmiyeXErHSQMR/4sYE/izwjtDo8JlMr
LB1it9kv4YZ+ggZ1f44XMVSzyCw/VuYJfIm1Ko1qp5QgNV8OtGAZQ69rr6du
4gTTEYlECqsu1njmVf6uENSn4tDbTlg9OsBluJ0OYnJaPxTPv2Sp8u/z3jbE
k4I8oIH594rRjEhe0ks9Hofoyzh3e9h8Z8t5t31zQuE6MALYlEM5KnjW9rPe
Nbz59xyMDjdPOXl3n6rpyytXPJDZO0Lxr4rw1w0qVR9RlsALZrDGmCpCEJz+
Z9TfR9xP9c/2Hs7AzwaUWUEaHm+toldl1IuK7B+nj3XKuXmmR6RqrOoBoDZj
a1+m10VGj6x0JdSIC2aDM8kjo+BJ6krJzmKcYcutcP9FbiUiaDPPc+Ronw3m
ilqz5HsuSgYB06foFd2h3Ow7QIOJt6OYPRsc3oHjkLGQFNgY/ulAYfm9ifFg
7OvQyxcae15Uhx8Q6cUKl/9mwy1ayjz+az75MUkYMrEkFoCRmNYoQgbNUM31
tDoyrXsBcGknpUEVgRgvGxWzgjO7UrQjtsxOTKqvgelQ3dLzLQ4QIIU1LYyo
TJJ+WZVLrhAiZqwpHe6vSQQs2MDMQpMc9oqqf0+Jq8L/gunRAvxoVDYcQFKL
j5Zu218i43cPoH3MQItvxiJey8zhiJ9kkRSEI58xjeo5vcNsLhfBxbA3zaqI
UCee5LMjwq76a5wsNCcvAHjtO68HZx5Gz3euJHY01OnwyBAzrRVDGF29m4ni
BMin6vUjSt/6KfLzbz9jYNo+74c+QSgVUl9eo32SZoNM3Th5DrXfJ0vf3qwq
gDbhkZJUaDixNmrTovZ3kFKKEz4Z+zL0CNifMWFeXFluWNlCjy5PqOwfBwDp
3R6srBVIHQddZsSFJtgAo1Mng/yriYMXdSguH+euZ/z1FJNL256Ihur6LCnM
d5geB2D/SCgDF7Hhw4a2WIlmogJZ0pfVtXHOb3ivQOIFMGp0ufWj1SgRaoxN
mpXgRJZeY5NXzy58KikJC6mTKBqcBlgR9pEpafbTaqdqO2/fnSE/e7EX3b8P
gKpy/S6PAri+/nLn8xTE1fYfbLs4ybcM0yjI398TI3JjoQdP1kfla5XlAm7p
7bf5GE1Ks5Dm1EPrZ/TTNrqsHuPwHT4JUt5/n/WTj55b/hh7ggw037RNYADR
TpwFYEW4NG5q36T47sgZt0DOichNSlxLielm6ZBoe5Ha2RtKf+mUfedYVFtC
wNBXjJXn78ZuYhZZctdUXdEHeamjfnqOwjSdVcmdwZOMiJlCxF/BfSJAe+6O
ejuoxbPpDoaLbvJ0I8RR5fW2KBGgnQj6mKs7M0mQdRwMMSkK47yXeGwP918s
zWhaf/Z1wHAAldkni9ff82ndVPc+d2s7+ssuvLuWxiJkONg3MeDWBqtZjWib
N2FhRKhv6gteboL8vPDLy04R3lcURzI909FH6g3zqd24ZdvkDdc3OhB00kF1
PYiAjd/BYlfHkgQqGKv+cf+9RKEiX63Cjzr6qIQJ1/BwtnqGchuO3eTgug+T
o8YK6k5HOf4vZpOXAu3E9k2KTTOT7qyKF066KMZhcto8txQdO1iPlQTs1APv
7r6o2VLUkb8ZRPdv63Ha6YKJnoPUb5ECi1UsX0fATwLIiD0q8Jy3yMq7/UCd
1H8SD0W8fx9qsGoIbJG8snDal/35gs2M8+vxlYpM96ZN14edjbvqQpoIJ1Y6
8nIt3CU5qjZ67SkBBrq1UOKT7tWMytIASxLa7MAIDVTRnXyN7B2bXtnwOOXt
iiopvSutZnn6IHZQ0uNYS3qoCMGz9dT3+38WXQxo0A27p1spw2G2ZCZsk5Fd
OAFiD40HCKOL0TuOP41DGvMRiMkGdUjw5bprmB9z9EKcr7ZYCr0SpTIrg795
alDQzoJCfcp0FCFAx0UP6qXCRl1rf+LSIpj91l95LwLrJWF64/aNGc44p1EU
nqf4KcRYPC1tle/BwE8CzghS2IrfNDjMVvYKy5QEHnmm19NaNqBw5P8Mk5Jl
eB4PrxBRwWu/Jt43xkdvsZSv2f6MHMmoJo8Pk4G8hN1SryPrheKmVKzN2KFE
UtAZCLM1W7g47XegmB3qFZdWUlL+OnnIWmEQWhdRretHK5GGhFq2PSSD+5kN
SIAPN58Gpdu6wfqcpxn78zdw0Nab+ODzzuhefbvR357sBHy7wCefDBxEXe6l
LSTx4Bp4GXTxL+WjBIDcz56tPyqCECEqe86SS7CdfluRKPNFMx3/iB7YFOOe
HHUx2t5Hj4G+sKZkIZePZ+aHxl2V9rSP/Tos0DOOpP+UpsJYgW7kJBPOkjLy
DyPp5QcWxSMDw1qKhBcwUYF3Sino4ez44MG719GSlthS3eLfc44TrwCGptlo
ZV9wVYzxHuRzsdUsoADbPK+7N26bYqf2xTZDRDGV2DHFbN260IuLTwSYcDZq
TgoXAcK7wHyBfyzdVVN9EPYUL9sxDdIPI2d5lu9quXgYxmgKglZSAW+Q3gVs
lUUfySm26Y99fhSvhag4ntx3qGbJjjtCzENc5EzM4IepyiyZ1GAYCdzHMQrW
J5uEFphjmMPgjMSkeStkmnk6esmWLUc2Y3KEC9zBRlwb16Jtpc6Qs5XHK9FR
xBZC/tkDcPNIQnf8uEkXMLghVGiB80n94syMWF+wQn+XjyTtNiv7NXbFua7p
L8xbe9omKtkbrLx43z1rkMjuPYl8W+TZKIAlfArScUwJpcAG2yoYh0Gol8g9
R0q8TYh1L7ADIUL+tv6d1zkTQs/ozGcs/nDoRNz1BSTJTk0DMEk+6jUdzOGq
1FzHMuT02ykHE/CK4CsRANg7KpePFZQmxerjzu2/ZfNmU0A5+qUYIaT1C87A
HccIycbLMOY/mU/ZRm39vjRrUbQanY5x2qVz1edi54cpqlLiX73mvQz5bQM7
X/orRYGvVfKyEnqkSwMBxRcVnDA/5N9bU5iu1BxgbPI/8D1WR2ELzqLPRylI
vjsuJt/IdcvsAB4I032MXF0jtgaQScWSHFa6mWcedp6EQA5dGwPCLOlp/lrr
SsWr+Ehxti85O8x9QKwf8t3hYUz8LJDXLbr7TANopN05pV5A6SrbGXTz8aNZ
H7R+xjThfwumG6mg1mtZIK2CMlwIiDTIR0FeE+NCyrOzLBLRH2gV7i2hMzIe
Mzo19W+OysGg85jP9+iaNc5sRDUQ+oiOF0QT0uS3SmEqONoQyYfvXIbXV4+A
7iHtAmtmEvXbf16K4ddQM4EVo6ffWxlIthN6Y/0uQVNh93RnPQs1pCDPSyg/
9L+e63vxJpmxbXYQNM0k8oW95MftlOgcwh52ZYhxTrHNuM7Tkfna/68Ez6PY
Vt4LWB6Wm89LxVN257Gbjeq3mduEQT6D8W6KI4NdQz+MUj7E0amxOGU4R0uy
Re10vMV4zRY+fpCrVSpPRS/eYAxt5L4ZZK+G2CRRz11OJqQ0ImnB3JtskdhV
0xnAnD34kKJDLBIxFd+shfsdY1E40nD0PBrU80fyMJbmoHWCXPI+UQky0MtU
cF9U79EuSkqpmH8XU2V+7alnIe95aKqE7qWrgGw+H7UQ7c5AK3NRgEKCi5aV
cqaOP5RHGMOxBCjXHKR3dTgqFOjmg/vWfcu+PoHgpcCOz5ZCYqgsdB78cQC1
jzlqzjbmQ+uAiU3S4PLR6o64FdQEB/7Ih4z7PDIJzeF1j2IB4P1J36tagm5V
Nd2UUuhY24WTEbx9vxYpctt61wL/KslhwRC9O3MOFE0MMiv/dAjLs+P6jTOE
z50xfpOCpz25MQ9OR0/A7GxSXwAkpcHSkLJBJ1PvfzXmG1pQ79OyYsIkhDiZ
IzCEdC0pw2hff6c6js8Mh4DCJXQjVnA7kF4O+DL5GueLjkRXBLB94QJN1oD8
4oz9ItKTzGnq0mW9f7I7yE7OByBZkZHIEIQz0zuSCZ7AVH534VPbCzyM6u2L
H9EjXfPPGmMGWMjFVt61SkPbjDj+DJMVmE5+QWq26hDWUDgEA5dOoh+MwUt1
o1Css+DPj4Y/9Y35AGAg3Amt5h6yHixZ/guKFLLYCNg54kk5yQIHWCbvmC/x
jV4OW11BmpMnFvF5rlsKpM5UiTKiCwL9GjulttU/00IuZZ9IOoTYFXvtIQSE
IgCh+BTOwe5ooHwXRBC1vV/AvfDXzxP4wH9f6qP1wxiWX2l/dP/rOXNXYIwG
fPEWXQi/YaANRK3jAEyIIhUEw7FWMx+5kM0N4Apl0SeaCtqYj3cMER3RzoPl
X3f7gDb9DIVobyGUhiiH7bKqKDmOMvptOQvDPpnIjE0uLVkDG1oYV/W6Zem8
DasZPrwTh8l/OUoTgjVLNdNGtHobhCoQuloQdVXskuW+dMz54wQn+B+bB52C
m3XBZJvg8+yE9gBMOUl0iR6OphR1PBk439c3d0hlU+Df7ren/pzAWZVOHcOn
J/N9lRw+B63dr7rwePrjltxl0dFtai3TJBPyhSXp4e9Z71ljhmKvMCknIQUT
vF9BrytgV8+fFYM4HQQx9frq+dhdbuXY7GASAvaFEJeILyNx7h+EFQcXMe1L
RCxX70l83w1dySDYmwl8ek+RvZnN1oxH0zoZo7wMxvjQfYj05gZsUepf2dIF
ThzOKcvHQJecawxmvdGecIy9aDSZnc9xMNMINjzxFGXMmHbpvzR9UjeLeq2K
jd12hhgEbTwojAAvqmIGbtM+k3LdhOB9Dnr6zpxYDd7n8yhT1R+ksjtXPHkF
K0zFEj3BIYpBVGtY3cklkEEHSj0gaG6DSvisq+/ZR82e14jdJVUj5brr6+GW
DlBuCqu4dyTLith9GZ19Tn0yr51J9krSwfRW/2tIdvyZgqaGkGizJipYJWyH
0qfXE3GfL+WnbP0VMPjDaz1hNM9hRO7PxY2uGSgrfXBbpAHqqct2YeRY8q8H
ITzjqwf9LfsDrYYlXRIxtzLGZAH8hTzjoT4FoCVJ6+jfC2xsLHTba6B6d/D+
10YK/0FTt3sCfI7OALXH1DHaz1YleyuoeKx7xD6K+Pqi65UEFqZBnPw9IfRY
Dw2gkG8xuwrWkqiKKLhLiZIuGdHXv84dzvn5v180Vpyht9Y9HZ/euQufHRxg
0/CZLu3EPvrwR6VHNgZ30/UH5zvvu2lI6Qh5qf08ORDgplbBL2U1jhXaGxPV
IZVX+ONd7Cm3TqH5u4D70y33MNsDSi0P2b9TbDCVJx35VIggiwgOAwkul4ua
dx9eClvD06ohi+lD6nSH5ZMbe6WcblN79KAj8vgVfSMtgeBdDKZwORokOa+V
EA+5r5risIsxOhJj8YQJ0trujO2gaGfiYnc4g01lmOYFV3xIMpuPhsujKfFD
nNUtm+3NRZ+Zl6MK06S/TE1yqszG0vRzOvqRWsguNq2f4ihnI28zVXTUnD9/
tkCFK9koQg1diZilNZovbm2ro2DQsiGKQGLBpFp1BUJCK4+CuzKZlAUWLJPT
yJDPGllswNR7D5sT/fTDjsb6HNWm+bKOJrq/D22ifDC2EKhvAuQka9bAJjMF
T6JP4rtsisf1J008X95SwCZJRoudqoHMm+eKAXFFzchzRlkgv3grP+kvBLKG
9ehk54pASjJSWXbAaJKenUVSTeg0nO8PHAIgA0W9r6RlDZzxSfY6ssgTfTIq
Qdsey0qkQHX13+7KqhoMO2Nfh8L6J0BARfyIWtNd7XgRWH1m62j+/gKNYMah
EJFEb4KdzRAWB3xF2wIGO2qGELkv1TjdRGsrxo83pTrPKwPXtP8pZNCIegMh
15pnwQOZHwm00pcRHYQJQ4ABqz1LmjCeMPm5e/5f016Cw05oU8xSy49f5j0q
AORaoXB+o5HHLZd97x9dMQwXLgfjU5Mf6kab5cAIl+ieQJJy59wJUUAC64E6
mDEZMyVIuDBpA2+xZ8ENSp2P5uHWO+bNK7NNDR28EGBOdf/pf+v9zth+9zto
i/Gvkd3UHuWREwq9zq9LqmzBDszy4141BwEWy2xe4l4MoosdxsTfjht+IX1c
zBDtDrBGAMKcaPI+CuBk+Tz8QmGqRT5E7AvVu1ZNNSnXXC98BTDVGtaVXJb7
+GeQxV7SaBJ5r5c04NTKyq7QkeINDOvpDvXjCASt3YWUSutV/HWiRHnCMOE9
8xwmCGOLj6gO6YVGgmezctw9fXa9YC3UyA70OgBsoSTse2Q4va2jiwQpgbLG
Ltg0HmEAhWx9u96wSgZctXkQ8rkqqckTLSaHKUstBUKMbc2muUmTQEPatT74
NDBwjuG0FUyj7HeV/18x8xyM39ufLfJ+Cb9JLXfT/iPE89PrEBWxDdpOg4HA
eMbwgm2hCp4JJRfRIW9ZbwAFtr4Dz8/11ruw/4gZ2MwjXcmnHh9fQhVUAJcE
7HTvMbXhI+hkWNybw7seneCcV8TsO8sffVqQ4uM6ggLGcdRK3qaQEpvFdw59
VGf0T/UQm6qWT+nFftC4hTFLo6COld8qgFXl3KgblvuOC87m4SjqD3cVisVT
02DOjoH/110GfYI/8gvpPRxCAcwawbXtOBr5mIEUyWUCxkS+eYYlQVja+z49
A50fz2Qvs2Damr53uLMPguK0WaIxpPs3DHITgnVEQvOV/5h4DhQw7GUy5XQ0
YWuvWxJ0J+T9YGiFgl2NXDcRuF7kJ92FaLVymakGoPHM5nUAlZ9v8Of1p4nY
D1JPmFXKO0WvOQYPihG1PNjA2aXqhNtKQNa+fJB5w4WxtLkyERhxJnzWVUU+
f6g0rQg7nPU6fzlFwXXsScEFjMG0c7TB/d4ZfnwTagsV4/JVn5UY3AutDZdr
ZFUsbvuQM3h7Eni85W1TBAbcTGLrxiQzfDSlIVvMe+eI2q8GZi0PNbRfQf9S
gmKa1qipRJIs+WJJ/FCCydyT0Cz3wvA62d8ODaFFknTDmic8NA9f7hXUaBlG
dUyhuC55Lg4clZBWrc6T3NtOtuQpL7EEw7nDBW6BzPbxH9OIc83C9BFyImQe
45jCHFyOlQVL7nGU4v0sMw9uvGbkbLxu5+Yss4p8tz0ihr+NUj9ExzI8BY1K
YW0JFEEJyd84fprb5v+5IPEzTbxluiFSEt1+L+n8OUxFrcnqVm37tToGqZBj
WULG9hLAdziGPoX2cBUldP5Eq64IT5Io/LDf7claZHwK3uDnjQt4nOEzgUHX
fDsug+3jVLxI6dUh8OTQTUIycmTvRo9hczaHQQubaZqyQ7Chz2dX4RmmdPZj
2759pJlcxzVr/YsN1eph7Lcsg+rWZyLkcW3b5/G+cXncTm3DbJXz6EGilUdG
iBaEbw17Ul7zyTPHRSrWxXSML3HZST0QGp0MjATpIQ13PSkJS4JLPyZ8WYVF
bnvs6YAkId672spHOtsN3bJt0GlBGqj4MP16uAdbvlkildfwvduJSO7dOgHo
XRt5OAKcch0FRRbtvWQVO16HevpVYXp6npFHXn+qsewAC2O6zvoE07AYx3uX
UmD6nh9jg3wSNUhfp2nIL/9dINntIg7OpSuiQQgFbK/WA0Rwd++72LrURDtw
nKdONOnm1CGHy/Vr2SyhLWs8qEoSXCXrSKazR+YCmlMYng9e35M/gusYbjI0
dUJRonQHzwenGYFRed8yah1QNASRYdyA8PvaZb2/EHf9bggBIC1kHkG5ukea
vQncktLNzzi7GxMjhrPeh5cXEiiCJzZCUU8k/Yx0OuZ32/jWKah0qYOkpQwF
JQ7k6M4vYozFh3V/wWaUdsXuzWNZDWTF3rYfQKQk0XPAMyy844eKLbTDN2Lw
vKuEFHrNMImqBIamoWmjdPJw3vPP9qevpwqqExTGR5HjlK9cnQxF9xQIYETr
Abj1Gv8sruj2Q/7VHFBE3KKTSIi956rPBFH/3vlSMbMXI1rz//SVKW65oY1z
86DXGA7h6QBAceeKRtXyPl2v+Uz4yIOs2QUMe7j2ayhwPo21t10p/RV0y4P4
uHMgXna2433+5um8gsTDu6F0TPIqxaNd60+2qli8yENdz3ZW1xWKBvbIBfJK
/FGGuY6FdsdaOcYmHNHEK8Rz5TWIk/H+aki+6u41Rjz3GZ+haJv17HcsVqS1
N0ea0ssS1+eYPtCLx91cHSfx73cS6ozFLSeLg6Ov1rXNVmNIiIKSqifmhZ2r
QpezYK5swx+BC365DO82/YLJs4CNu+Tw1j/ce2c53Zmqu4S5+kBvno/93HJF
BWQEaGZq5tWTre3UIgYcGLvDqtVNf5o8OcmxHt1RtClmFEq8d/1pibVvDuIU
xN60smaHeOT6naT2bWF7ANg9yOI2TasgF56RQeb5n3HI9ws1QaYWMhbrZtx+
u6nAqp6Ub9BAtIDGWMs8dRkDghpjyT3hAp4Jy3wExCILDocEs9yS4BYoJBuB
RcqjYg95nqSnGks9GtXaB93iw286YNyJICFTIMbtwWZN3Cj+FK5h5LjS2waM
/iGZFpXq32Hy5vrjbggJbrgXx9apO5ZJVgT4a8xmd9MnnvC3nqH13znAxNBk
5t2u8Ax7FQjnwqoeUv+V5eV5Bd9SxgbZgizeIzdecQooV212liuTMx+OXa6X
uLuHBUptxDGbGu7qjj13pdFuPi0bTzjTkDZHJm5H9/WTicbKDDS8ch3rRvNU
R4Cx1XVuPaE+YaR83tKjQmKgAI7wIy73uLhcODWKNMQ9fORVl5BI+q7iIIEO
E6W/dhAR/aCd2Q1rS3+hcjn8ptXREzmhA3S4wNcPRYhzu/9UGIXIILer7bFt
wr+XdZz07tGj4CZOW5npbFzaxI8lzedUAgsmTofZoVxhXE9jqFkwCTcVscb6
wGDmAhKLpTaYDEl2W2K5lqDw/Bqhlsr6tY+6etKiwhPYs7o79kIgljikQdBD
xFAMhvntZrx8lDTchilHF3zQ1RnCi5SJCSUii8wJWRQfGUMRRpcnGDRbpayO
pGtXSI7C/kvf83iEQitfAGz7MOcCgL6FvB5mYAr+e4SJIUlnHd1cX4nAfx1I
9boTJCedLOiXGuiYUlZDprj263hHwE7OL7FW1vRpzORPeLTpuaRlJVlHs1tx
sL2YcnBQ+M+ne23OzLCqLpybHUluX54i0zfCVCQYgESXyjj4g+mOGh2neQ0z
bg0tBWO4XriuOtQW0/g4FxGwtEE0hr1HA36HKZ8v5Oa99ifC5f+3cGrcavNP
/wUU8ShMouCtj2BYa23Jki+9tTwH1QJOuzPOZAJSSMJ5ixRdKsqHt75ogw2Q
/SSmwMevsAGKYzo5MbsClavOPEzkeaFyO3luA7BoZ80hjoYcooWrzUzVBLVZ
dnPdL/hWWVpN45aWoGqhK2mc0QzowW6dC3FHNk4ZRnWfVFaPD3Qmr0ZCHEzs
CUvmHIY+r5FFIvo40pzDd7LlZYOOx4jc32IBRyHzNQ4+Uyq8nxIfSf0eFcZy
h15bVndJiTVEkG1leFS7NLFryTlKdih23Cs1uiIowuSDVOLoGXH4NUz0WmMF
q/H6F2OunPfnOnYE09pHleZcB/v7klazm38J5FYt8dpr+dZzqKQ9duaJM5A5
ce5WnQZ361Wz6S2Qx5K1GxW9nZ/MX+eaVSMSml1hb55dBbiH8qidyCEUUkzb
mwRa/lwGHCRldg7AqqsRujvGngN9GAl4N0E9eQXKhfpR7n1Z0zO4kvKN8KPS
us2VlcvRw+qEdumkSIStFvwNMcul7hSdjUZ/IdFEtY8eIApjz6gQwg+NICxA
cyXCMQ1s3AWpdAAe2ixBH4sEU3X1x48i+YnWmhT0rFDP6eiFNWqLKzx7Crxw
5ZYmwKKlzgKBzzI09ZVJZrX86LnsHh+HQ/IKVYEyWb1BxJYfWyvOJGVXgLBs
Fq2TlFBY3UMuSHaKAO3S9ZmcouqEFe6YD7JsJ2Tlemdc3EzbvUZJAXA+3vYn
dTjSwfd2XZnC8ebgrCKtaszUE2OXxo3Mw2SdSYrlziCLXKdcuXbB3wkQ0HkJ
gb2sAz8gB1LBhKlURJhDz7JusmroUE+2nuPONvCV44827yjgm9ba0thP9434
HygV77XSTZ4csDzWzxiM7wc3EXXNlV7BWb/mBhaV8hWZfftJWLffOyCk/fLY
fmbbnqXV+ktbwJbXaHrxZPl30aqK13OPzazIcUbUJ6r+KNgkjb8PaEr9uJ85
8LBNYjeAvy+3axS5QYzwBP9pkNu6/FQC9xE2T94Hwctd6wXWcZTlSyOH8Z9H
4CdZj652fknjVgOuRNnayP7nfeADWifSYoUtftzWFp4rtzs92sDfPi0J2Tvo
2q1oIzbdMs8E2EDRSsjXiJsaU01Mp+/CSrcODRHr7TCH7KM2Kx2QS/w9pNTt
DBO1m/FR09eBaR+qj7EPA1LLFZtE7Tb73rc75452X8Z8TZ0BfcKVB+RJx96f
cTEvy+IZwvx7/4PKa9nVSo7UimsFMWxQFlzABjFt6qdh1DbRM7YDK+/s8mTt
fkV2wQZaHcOwQT+HdEfSm3X0aM2elIL1xZIRGIhfJveCuZEUkyXinu/T+orc
3RgRw46FSxeF83ePMUM6w95WgzlqFwrYcLGP6ZB30ZHkMDjaGcotGFgSHDkZ
8iDbrC9LOXnjTICNrUZ3By9UNQ3REE16fSGEw/rqQ5aXXyrLeYDvukgZK4iH
aDuyM3TaozweVRRN0VTq9ZCYcXOsiX2Gml8rus6TceLDtmeaGBzpcOJvqOBf
geD7Vhw8GlWIGoTyZUIjqlakd8loynmb5y2mwMYM1ENK9EqqJgFpNz4z9Qwt
9b+ek+JH/ARA9rvdZuj6q3KR3FH2ow4vLKaXYdohoN55ypNOTjiza8aa+SAD
vdMQIOoNhmz8/T8QXvI0HQ+zgFOgg4nkbCVAkK222QIVB77/ZLBo5omf4+ST
YEF/yh4w4BCbgOmJHqK18IqP1F4wb2NzukO/OGMmVq3/j0pk9NpiRQI69SgB
VAoNpgrcD2vnqZEd/SbQGa+kjnKfkJy2DwJ4VlqsjGyim/qoCHCGCOos20FE
IRFIogeVHc8fufd8CRVc/JefGEETfFFhJnM+wMW9DZ+by4i3gVEHVoyLrsqQ
jml5UMhZI1ZnE2yIXwEdqqngTo6tebzHGo03knhRUtZif8THZ2V43ya6/nDh
Jgs4rkyMkExrvHKUm5mwqnHOXCZ9quO6drV5ccmrQv5BVObfLwXzkyhC31dd
R3qCEo4fwKBcyvYi1QBWnPJduKmCBfTRaTNZpTzGbvFujvcUkL8xkzLHCUgE
8Jx0S0KeN3d4Ew2sYHVQyHksM4IBJZNrJ7ceghj3FzG/FXzYQDLFkHteUpWm
AocUpp8SLZLeEoBPht0ZjlpXp2RDnkPHAFCKo2QJwc31cVoQCYPdLOT61N1x
0fLQMyxnHfOZgEpceePCR4tXlxfXLY2je5PVgSdE0O3PqJ4NuRurq7/jgU/A
zQyq0vDuXo8wCEe8SO4BbtdCn0GjdoZ91rG6Y8TocqbVGrmWNkL/uvngOnFm
tOOC4bUtD8OoC6xGPACke65QXZNFfEbcl4ow84sTb9YOP3ozGhm5tRisaGHB
iwo7gdSgVdZI01EsFQGQgE7QbWIyCbwOmakTlk9N7y/VJVXBISANDkKvQQWp
W4jOfTOVw1K7CHdKB5qXwrBKeZjd0qGBqfVZfTWgH+B7ta4QI5tKE1FfdvYa
QcKTSwJsnc1fkTFBCQNptBc5bImu7FI4Qq9av0M6+zChRfkuKCVNAFprNTbg
Cyb8j8XRXxF+mh3Jm37LZhTa8I9lh2++u3I2UttqMkDyWZqT9kCXpmAM8InM
LT91Qu5YJZH3yfIkR8jXd8XUKANHCa7Zn+8KiW2FkEl4Y/KA95seBXD8b1mi
SHsGX/aeGu2oA5QbM2w8dEQ1SqH795CSkiRb1cuMiOWHdZLq10ki6QyrMvWY
FOVShspqXislezzyOm8c9DWPlbqJ1a4wt19aemciQ5+dBNhCAmDrx+YKGI6K
XPVTDpqLd7Z8SjSm+Xs0qYax8bl99kqZsQmWhtcmf5EvY6cDOQnruEJDsYXX
N11Frl5746yka1RXG5aSzO+N0H97mRcHyedKSbU4VMosiCPMVwUpYKuo/6Rs
Soh0V01PZjW5xuFfNdFZe/tCFTZOMTERkxnDNukyokLBDXM+bKQLWbO4BeOJ
ZRNM++FcBCY4J3KGu8g1tO3RqolFSr82bo45sLzcSbs1usx72VCBNe2rF07Z
zs64Jex8BBL3Ki88GiXgMCjHTly3PX9prk+JptynpRbxOodqpl+0vhX+kko+
4R/UDZlkYSs/29yPXPZZjw2scvld5Xqa4ejXdPjYJvv9vxqyqKy3E1in42MM
nF97EETpRxIothw+L6SdFTu6plnOKg2N1mYYokLG+gzn8MSw2r2CEs4L/qpe
YkWFCyH2UVITSDy1ylRBOJwrHtt6VfyS1uTBIz8QqC4XkrClxuyStPI9FF/L
4OZVp3IQdtVWJ6yEDePbYIhj2TAHQc4MfU+WjcTCv/nQp9LyUdJFjH0awa0n
qUfEvbsuP3550Zb/2jOhnHoPJMq6p30CFij102NvTEQ5hrNLhI3GCE1aZikm
Z3dDUoerwaKBIUKh39kSxUS7Sm1QC/3ii3QC3JMCVRrQ8Gzk4cWneSYwm1rP
+55XikDIVtKv7AmaDfIm3OZHUKY+EXr+x6dDP7CruitMDLI51kSIVQicSF3Y
4SZvVlcF4S8pdQUwt6MzOs25zdP4ebiFRZqZxdEgU5JOKQTkFfNb2lmlPWW5
4VuhcZtCb/3ENE3qbjRoLbzAhueGCrgow8OR+k6UtdRTPzD225yt4Z6GeOe3
hSD1T/FcK1sBlfuUXc43tCNo6W5CxrARkH394o/gexcT8yMGog+vTqSJG2Gq
38Ttb+4D/Hf/Aadr7po1K9GIrPvufTFmLSnjMcZz5kgfwKc5iKXQIHvc4Smx
jUp0GFGCdApl0VS1sOucYz35Ea049KBmQzs7zVB+UxkKD/MqnDWpGbRLBWIC
6cDuE8utZrdEzLPLve2Lz+3SrcJxLa1NUBiMA5E2d8yDr5jK8Yqf3aBcVMDE
Yi+qiv4z88ffOTclc7qLeAooxLD6iT51caqzfJgZF9/k2ZfoSwR5XTBitGMy
7F8WAojHOWuhT7fiZX9BcJynQEe55EzBDVY9/ub6gXcMStYUcD5IYisp1Ywv
wYkLmNO3w8hDkc3DyzwCmLF5WviVxI9qqKofl/I5nQbXLw1l5tagAWN1xWel
xRyerwd/zI6mp11wXrc98EMT0v0JZj2sKGgfGXidewo29PEcZSPn7zGv+K7B
QuBwCHj+GhH8TySD19LiGhkCwe529TRlDB+H5dyxJXkqAFg3alJ2HOsQ8RXT
SED8ZBrH0BxgsNluIMHvYVfePkXVKEVRgKpPYitwWM2pxDcKfK5sDjfALTsE
Fa2/avvUTNK1Ia9Vy4fjV4qPpvE/rnGdcRDKf7qoldIR1wiLDEDTSGWYmc04
WTE9PJeMGKruG5IAkzXD2B4ukNewgt7+VIRFISTDasE6v9CXuBfvytJFjpNj
rwO2fjKFZByOh6OPIDKb1RSs/93lUxHUkxOdxV06R6eSgP+90j0be/TmqGy0
viZ9+GoBrDyn22LuU6mxS4FglUhNo4c+16wrnfxhhlMD5bjs+n2QhdH1sVf2
qmSsFAYR2zlt/cYAOk4yKgCWSEujtb2mN6mKYllbRtkbg8JfIbuaYqkCgpa2
EB9jMs9vNlTd7rZDYouAlGMKIlgRVUl4Q4X6cAdO89LzItCtD+OF0R/auU8W
iQgK1TbRHN18UyF2sndSQbGdgJt2BjTG+ekbfOsLTsLxZUNCucmDmIxzAVGR
GcLFZ35vCu7i0g/AoDwMjuxhTEhngMkQePjVlUal6YxhxYD+36pqCj/exFVD
xNLUVCPFXubNpLyiKo+OXyyEkWh/NCk9Dje3wlbON9V1ke5CrDJAzlTSgFv4
vdxNI1xNJaB94AMPm5ydMaYkva2PQ+5BCDrtjZhTxfUsDjmL9Yx4WkN63xrX
ZnFwRprppfLy7FNOReHQSBFro+dc6WfydrPgj0XJ5OcSr5LPLC2M8VeN+62A
O/uLNVfSngLWmpCUlaxAtHGtGGPh1fr/9e20AhCKTX5gRUkC/lMMJq2dK593
kCMj7d6ejTW5hWTm8iMKGyHDt03aFfkh5+CHfQA8/15QLngY75t0Ioajn8do
kDTq+A9nwcAvUs3ebYe7gCyOotTX7cRW+AuCEWqv9GGhn4i2oakbGsy/lvjq
p/1bcyHB/4G0tYb4sTxiVq7DhU7HrMNn28Lq1IIaJv1TlyZK1YSn1e6+79WB
gj8j6hJwADcRbNXl4Qv/sSucQZjLEJPTlXGUQiL0noV9HlINIlB2lzQw+ywx
mWJBUjzVfRSdIdDIrdJ6pMy/nFiaHuzuYCknbsrZKfrVutmqjlvV5ycY10VL
kgkhitHUzOE8Yu1aO14KhMrL59zNq6SGqx4ORTbf1T5Q9MYgjDX6TKdIqF/N
f4r+5ZKJIkYP2NQE9847OWVxszblv0tWEw3vZXO9cKS4vcKOQOVoNtt1SbVX
KZY2UQmIM9LP8yulfZMgFU+HUP1C3HvrCzjWhpyTi3fLLwWUSd54W9JzMZqh
Pw/QjhLx9NFhCKPUT+MXmqJq8dd6oQI3JG0kpDzzg9Yn7k0aFkdo3c/hrrc/
vLq09DwrI2JqYetPjbaW/X9BnOhGnJNCd/M+5PQpd3UVQ4ky5x3JE3I7tssz
PtkxA8PBfJNj5jXypdB//KtLqpQxRMnoaGZNTx7R3GQkORZ2jDV5WNlrIcvY
uxfqKin026CKFNJJicZzpdRiMq1xSyLGzLdcJoZAJDA+X6j5ufwsTMM1kyFG
auURS+jeJvVUWRdef+dOOOsiTh/cLFT7njImDOxtxDoRuDMUBPyAIgSvXS2U
Cvpg4u26qxOrHk12iHkSw1VQjRtRw1yAERD5y+Pxe4Mek5CNUmGux1Qs8H0/
rXzTrc9J4fbKaY7XRYknYZHJn4JHsxNjLIQirRytRXPDEzzxkaemnGkXL4Aw
ooV7pj5p1hd7lT/dXSa1OjxLSlUQ4nor7CcD5rSsdC4inqvVKQeqt2N9DhqE
S8sk7XfgnW0Vm1Do6EQ7ZousxIiYJ5O5M2ajkTxYvvrf3mG9L5DV75kn7a3G
k6sDkp6CfNU23rsmmF4S1J7TB3+L0jnMjnNTTAwYpGhMVw48S90MRBC9uw2Q
18P3iiRvMq06bZ0A6Z5dloTqyaBA57Jg1kySDGcUTifVyiUxyeFzFSXrxwTw
DjRy6CAjp9rmXbQuUyXEGtLq3rjNavdH8o78/yrDv2ZYttg0NfMxyqKFcivI
DIkjyPuziosCfSxputKtrY2Pm20KPbORqVUbgQ7mxB8XkLZ4zd1Cck8jddWo
9e6ewJunsXJDlU69/hb2vJO0pgqQHmkLDN56TJJgTT3TlWRKCGbbq/TOUQ+L
gl4Rx8dynvA9kth1l8c/FU3/RIzrGvFuEhdZ6xQAhqfetUCx6h5006B0JPA8
g3551UrFKv29RmA3UCOiACDs8uRTlXuo8tnfc3UCrIP/d1+vQSd3deUHObTR
ovooiuU11q8RQtf7jBpoq9myLN/EY6WMMUfAxlqY+kvUK/pi+KL2mUFIrpvj
eWpvd9JEonxuWGAf0/kY9fARdysSKuypE8hIRtqHVYEJ+TwMTNO5iTmu63Ew
YCNkn4HX4XU7VDmKUCWIeIpGDwt/jNaGBHw2jmVgX13QC08w7b+nU/AWmM4V
qWpn5gaW7M4fmfe78XpyMfx280bJ2sEaOcX1ZqdM8QOXiqemTlvH0zMRqZkz
8EOrZHhyEpHVHtwhb3l8wrLd1ssX3lw/j44QvDbzqafJ3gBhfAvSV9mbds4m
zyZ9M+dh6i3MskS7DeByf97m4H+g8NhRlmkAIAmiHWv+tRddc62liN+ULkgl
ZymABHvUa/W08gSNs088LkrNWXud5MZv8H6GEYMD3ab1Tlvwkstz9J1dHZkO
7JCtCXkGivz/tzRSqOJPTwkKLuuvzo7LkUFZc1Q9pVlxcHSfWuov0SfdnfRj
hAC7efW1X9rJWPH8mnD8wOkiOtIvaCgk6MSfvDje7b80uONPGVDp8jrrt3gb
gSfrPcQZ0uhJxUY1OvWic1cxyKDDfeDqi+tWFMtofNhAi8e2rST56k1UqbuG
BJY5L03BFB1LPiydOBDERlfmpUA/Qtxu68xggSYf3uD/vf9QVO9JOzo3CRVR
w+VRywiXJCTgPxgMev7dtxNRCU7l6oFGQFBD/1tJvKb8OEs+/RH30V2Wp8tc
7EyvwOesy9p8BJ4Q4jO+UvaqIDw5/PpI5w+P0Ga77Xc3O9EY11dCCoVukvXb
cHwGDVqng+fKvldJH8DuCbmOMrhJ6MuXrRXbxhqZhd0TVAB5ilQrFt7+ss7C
0OxbBjLqZjWbtt2PpocQ039PISGyXSQ1Z1XqwTG64d9JPbRcimukC0HNl9vA
EeSPl//DQZn/sGHqullqVxuW5jsOxtvEc0wXdD0ZgTqswYfVpNitgDCrpexb
HfqGgKACXhLe5dsDQUyRTv9xJdrH4k47pqVYo29J56zrbAYxuNBq/qR65lo1
CRYzhUzUOynPZ8bIh8xqhZef9CDP3BVRhadgqeboAB0nNTYKRPzkyQ9SHn6w
o0tIphl4rYHc88x849rpxoukkxIq7vrzKX3qltOIMUvF6riItFMTY+PdWcAY
15ryU3F+Gze5BkWR/TdswzjfDLx9o2+UdEobPDjy/1UK6hAl1HGl9j5AUnM3
QNpgQDaJI2vhyqLXE6mRA0jTEXan9ETkRcS0Kis5IOr/qEY8watG9ajcT7o1
E0gCJiUGpfWaE5ORhwmthqbDRrBUi1ycNxtZyb8YwRg8tQUgMs1emFcnVA1U
Qlk4ypwDOekeKXNbEfXs1ysCEuBAfvX1ZutiO/S+xS3W+CnJqk497LITaSGx
XtsFgj0KzPwtpHXkO7hfG0hBdk24YobcBgHTwNfuwCAOspyYeGvbKT0tg10H
fTYBNGT1d/3ki8Pc8+rENlSrfrjvTHgGOikB21R1zSZQUjMBNK+x9Uw6iuKK
ktdE/ypp4uG2gudP64/1WD7Pdx6P8FbOgZ2zyyhV/abfevhqfg4ywj9NA5Xp
cl4uuHNUUmXoTnU2qHcx1WbFkbmngOTaqnYrNr5QlA0jWIi2Y62iOLRx4bGU
IAt1hHCk92vu6q3PwtOqeGhntcbY5mkzNZV54JvA0DEVBCeH+YlAQP4ElmNc
k+wFpghCgu0i+BkON+7r0BPcJqSxs3MLRQjXZU6aMHXWWTh2KaWh41VHXOtq
g4TJiiOe8v+Huf6WOxKCUaVUytlzc1w3cBIyqRufawUv+wVGBq2xYp8maCAG
N2wUi0nQhPqMqc022U4Z+mko49fjjr1eEMiLdBXdUY4qPhYTFe5PLZS7dMpH
x0z0LF5IrIDJigrGXCaYxbz5gKSIYln/U4bN1aqgNRxGTG7B55FtT7adMMPC
uWrCoJwv5mcbRMDRZOSwF70Mtcay1bthcrQIWmIVRbANrnkxkX3F07E8oYrC
2Sl4Jud66SXlfjsH47wDNG7GZkeP3mbg1r9tEtwqYpGskTItopQFHpoDArJe
mkJ9wM9akeQdCnbxXciybQliJZC96/8f3Qc8Tw0xKkqDfbyRfLGxQ+Nf+IgD
EIJ2kt3cIiQtd3WqkSEc9BLGpkbbLtuLnCKEkyA/FdpPcj6jvq+FY4WTECdM
F0ING3OQBFX40cOEbYavFh08fkeJUHl09l+jLic99oo031zCVprm17PpeCwT
gk7ymSXKEBpfIC4wlhfbdvFsb9JtqdA+idi4oQ5GSVDLbJ2wTosuOxkU3ZbS
iYwvoTasdc5PawCTFf63r+KyyGdR6KWQ3OPzyJ8/UkrPlOg8OXfXG8VPFxr0
TVIZ+DGnwik/PHPjsaQY5667qC0+GkC+tgVZKWMu97QYMteJbK3hvxI8+IIF
Q8DuNTjlW5hbfPiBhh572XMqEOLbZ8QpwNuE3e+Z7wWm5yCeTR/pXpWUB5oz
EQ2hvI16D1NMqTyZ8V9ca6ATDc6PHEGl4WeZUA15thlmrC3ii+1NfbOSVERS
jwZAyIU6se00LZD53SjJCLkd80n5i2zLDqiTVYgSrFcfgq1TEwRua9P+w2Mm
G27ROCQbEvAHhYkaOCEVp3gsMl8t49TYoCH04NS5XH1MoR2/lCe7S85UqzDV
PenY1rtlOg9IyTeF6GR96ImUT6lNmdEwctTf1/5oIzj/0YSEi1FAuXYIabJ6
0hM5sULnY56wB0fl7m3oYmWcfidnl3+1vWS94Jjei9Ae6hDw/UHktmfRwt0A
GlSYeTHneDuOIREYQwE/VDHMARrSNJcDicZGUwhbJmNDtYx3naF23w59Pe+h
u9D3ndct+Ebp9lQlHsO5kC1Vm0wVOpgW6Vac/5gJXp/+TMu2K+7TyPlue2Vr
vBpTxSQzAHvue7eblAIqcD9SIe9zVXuDv6jbhGgAVkRwfz4AgSsCqqyGCHpy
qrqKXFRjzYaI0CKpK+E6KjiipVEbA7Tuc8PrfIPTYBofYAYXe0wZE9zbtXDA
4tPglOQGXpB2cKQQtY/RZVZA4eOXJXBJi5nSC4CZ2MfsAsG4Sy4s/j1++ntz
rJrRWYemE6JbrVi6cXldDZZGmmKRIJ26/JvZyEypdj40mqs37g54/oZcM9wG
fz7FjuhaRjVAzTLtsUZJCb+TIvxUxyxyZ9EDTgbRs4i9FFpnK179OdMy97sR
77jR9ypV+1Q27gdgbzL6l+JZ+5Rrvb0cZHGygIn3JN1tzEJGWrr62WKCLiNM
OmyWzvqR63OrtlGUenas6M4fHloTrP8oEjofpBsAYUJkysFg6a5aha0VQvGE
RCgIrVXqMxNbkEUkO8N+Gw07/orFEXe1QSKn9FntmMQBStl7PXjSQkVsbnVQ
50uDvH3ITdGxEFUotU/wNRFFPUB3SDEqAjWQHz52uOGI5ulcRLoTGtaeD6qG
NIxRTyDSEMSBb2umOY9vqeJBLyHnJ9a7AXeob8foxN5jtNJRS5PhrS8wHxih
O7+FWkZp00h3LVacLdCVzyjrfQXlRKYjqxxW6/pIBtu8npeB9AJoeAt7M/Sa
C3MUe8Xo7OgwzrrdsWhAtPurjop14U+va16z5RU/YHEJf3qVtFEWYMo5dlzo
xqFYOiutTkOjXtWijwxHxNdx2Q269ES8klGZK5EWbUPq1EsDosl+flJFeuYR
oDju8pqBGqZyH8RK4Eqr2qQgQ87Oeqmg3RQMU7cbXWePz4ojS+yUH2H7oOUw
JNanD7c/aB14MXqq34SL1qQvl7EO27L9WrbA71FEdl+onL+Gc7zZB8+quWcU
C4S+riVNXBEeJjq3QZcp4IB9ZghY7yIVjiI+IAwAMkVbPRn9+1h3rQQzi+en
E4EvbUa+tb3jRwxSPCTMtC4m2KCv+aJRtKbi3HU2Nsi9Y4X2xz8DIZw/CVVk
0XfoMhlB/U8loDncexhXEdUCsSXiN6zu03jVnyeRvdNZo1hryh9HUdgufVLQ
d2qCqS3fsfLgVfBUy0jF2LHJNTii1yh+jJbvBjd35QpkB4tn/5Ls1VrNNW1v
qYO2BmFus5iN8qP/XhVFVuxBNfIEiYZUzSejmPJcIhH9zZqWWHiIKTRc22OC
SJMN9YZTFgxu/10nz9xER0M6braA9UBOH4VGayJSD7kz7X7WjOv/3doHeK/B
oOBTVoEQgDQrg1dBFn62E5g/oE4Hvi7diSbKRRIyfWDfcUAPYfD8/eJqIQCv
LBGJGP6ul1PIWs7m4/niCfr6MAWO5lD8bPtAYv5zZoHcVjHA1ULbSKO6xYU+
b0OUjx7x7Rqz1DB9uWVNx4NgxZlez0pB2wQth13/c2pr+pJ6/X4eEFhWJEz3
lDIoEh+i+D7atcEejs4QmOXdLIHtBN5BWNOQUwssNGU+miICOE0H4U6RQ3c0
jobMSKXGaIqO+e5E9oeZP0Yp+QO8nIPZp+4WfiAXJnNb2TGZBVuEzKdKENPi
uqataD1YiMk5QncyJr1MiUCViNh/o5dEl/c6dcjjmGWJaEkzi9w4uEJqd7HW
H6RVyxk2Z6Z+m2cldJBPPy1RxBkywBKKeF7Vge2Lj3EdmzlXpf5MVCQ3iI+W
IcgzQH5JNn50z69BOSaUxvsMBz4p62W2ePzcKdaAKkpfsZ/ae4auXDiH0GhQ
3EPf748bKFArlyIm0HhovBYIzQMgplE/dP6Rqo4yILbsKt2Jch5dCkYBPmpk
Om2Iqe8fRz2SEb2ThIXV2nC/j0zUu9yE9cB4QD38OjHW+w6eQvR8/2fB93Fj
OdRtTQ3c8z/6TNLbv6XPZbVmAsHvTXbTr/Uur1COLH1/5lN1a0Ur4LJep04A
3XZMc46m8RQLF9MC9T3jR41jkIq+vjKAZJPtTP7Dpk/j9vhJNKvF4n8khuO0
JTPqgobIQB019szGLYmppDDI7IfCV7Fk1laTthzDY3CIi2Dox/X1Dc21BBBp
UX7mFqiKSKfG2IJAtOCeN2SwS3uTOn7QSvZBuH/mnCpZrYw1XdgC3q0HynxP
N9ilpW998ZhJzCDOuW7oL9esIZ+jK4tMcg+JM4tLTfd0IVsOlPZx5FTA7u0R
IAidD29Zdx9/7xrxvGfBq/9x8NSGB9Bb1PFCz+vBJMFQyR6imHarDCatUTlb
salZQZcnP9hSs0jOJiTK5COtiB0QSr/k0D5cT5gSNKYg/uEP6+R+21zwN/sX
yXaO22FaqHohLE4tkgJnFq0F3l5E3fajeVBXfwX0Vib6KKKOLJEyXQC0Kw9r
+QQoVOF0wgEEANVj4Vwl8I9eS+B2cnzCUBc2ieXgF0mzoCejJn9DGNCcUT/Y
mdofGiUWmh9cg9yQL1Wna7+mgI4GAGePw0U7ryxLqIygN2A1M0G/JcS4fMcd
MINUScfDXRdHp8SMRh3olNouKyfOx6m7M+WZ65bkQLmleu20HPvtkV16FGVs
JXyb4yTmy8VfyulNqdku8VHV0ABkCS/MF0Vw30fvPGdmwWW0URFZCZKn7Ex/
hVfzi/+pFIfPAFA/98ONHi511ynVtqCxHi6cJALLmpiav5JHkAteXsPGTrpa
VosUa7jOZ8fzFJmjxk6QBZgB4Fpgsuf3iS8g/mJtEHdx37Mkk7AdW+28N9Vy
hxXVr0nAelTmEqF3sUixSLwsbWlJZlIMDDIdp8mJmklEx8EVAfc3fON9LoIu
ff2hHwuFgSV59yQ3HHTF+31IdAOY2qzqZGgpVVmUS+sdgt4XhwjCHouCphhL
BIiyDGtwnfDgofMYTTeTc7aP9sojrnF0w9MoNn1nkmw9Ln2LKzMCVn6RuWev
TA6o0glsmb5So0lp1N/6SJixmMtjtL0L+OaSBEH0hfWaYl98Nox4q2SZfn4P
vAD6UC/acCjPJi5DPm7MnDFP/fIM7GIP2puOexeP8JvrSUU6cL5EQTme25E2
aDlP33dLXlbb4ARNQeWSDd4gJhMkdor0Z9rLpzzf6rI36DQxUM5Oo/8V2taP
dVWc1bYUl/oJWEu9hLy3ivH9bWlmQwSel40tLFraUn/78w+r8osAFprU92wl
W68zAeN9BzZkyVIGM8faRci50SGxg234K/v0GagRVxmn8c/9P1qtB2gQ+ugQ
5xFOAgxRhJykt9t3Q5Y7Arj8ZCAnsHVVJIF1//MxZJ34f7D07/DVJ3yfrvVB
XunCEGkKXS2lW/F190wFZfwq4ypdkpbYYDYex+7RPhGR8dKuUzWSE9ynqceh
tFEgqTOW/GctwK6G2zuXheLOYCwJB0g0HTSOtlsIobcZBlr4F932wZ5j1PVD
kQVI6NTAa8Gx1eSnD/jw7pqFC2wJEccYA9RS3EDrpktP2KefARJvZJ9OXtzV
nM/L5pLxa7D1GA2d7MXNrCQknmdXHqeQPDUIgQirEpgtScjFC52TndvlD4gl
Dr76PrGvWkD7Nt8e9deYXwM2iJkWmmBh4UBSFmdfKSdv83hNKcWdX4F/TCbA
yALstkXz9jWr7le3RRjxyiYHrsecT0z02A5qCXU7lFgF4NHexAUe8BsUY+7u
jqvdaPM8CEhRgVQAzXmgDvfwARRNh8hhv8DaB3nT+u8xfvzrzM5aODRj1+Ef
TG7l2NNaCwuq9PLzgS3Kdd51Bgq0V2KvHjHZ/ApB+zPPBXUPR5fMnuKaCLz8
aAtB6l2/qtXAjY/xdsYMiLUXwLFWsWIEDtVN3laRwUTJ9bE9T6BNwbE5UJJN
oVx7BcpP6dA6JIKPh4iCB2plVgXAP0VFy/zg9ohBOHKJYtB+npZWWN86mPDg
2F2+tIgt0EuAwl+lZ3ewzGKxC8CWq0N0QoNGc7RMAwxl70j2znKJIf9Tw2Ev
kbidOVx5jotQU045Q/1+kJaX/t+qCnrMAUwb10VTkG2t3zKpXkfnVXSq0it9
GFyXYksIMaVPg7Pgb3zgHGpWPDMLhvNOPnRHU7U3AJAJYpPFtrSqQbX7xxK/
EAxMe9SwuR1nqhQESPkaQPzrG6a4O40j760XeLQtTpZHpWBLG9lBIrC7o6Ya
nhOjmdDNEyLDhl+q8/S1Z+E79PvJVnrQXJ8L8M28BooognuGxBOkJNQ0syQf
ZhkSojzzWLbuYvNRUY+MZHo1rBozElkNixsKRCrixPgE/00IqlmLv05d/OxN
t4/eR6G5xzmFqLl1yQchSoJ5EOZAMSp1w1iAXMZ2AdClDXlkp3EIdUaGkkP4
fYW8l6E+tebQOUecTJpQDc9hgH3bJdmR3FU/oZ45zX8rI92XDoZfs2Pn0q0+
/6AVCz/KsCa9kKVe1KUMfAC+LGxrkaulsiMYHZHl7rUNcq/cDRUKAKE+0ixK
f7oLfmz5YJ8goypF8MXLpfh3WWqDMoVatoUtfdykLGdLaCbCiRNnlvCf+fXZ
LOzIMU/T9Z7MgQ7pZeQaPdApLOktZq00ekjQLwM94bVygsmA0y9wtCI2QWaV
79tiisE9YQuf2ue4sCwsuARGbzi7zu7g24vAmHmMWVejpuE7Vh5dJDrBVIuj
RCdECsYyDmlbHUU614mQEwfSLTE5Dk3EBJ/EZLoXp2AYLE3T/40In62AaBlp
oFOTbSS6/GrrQz6UUeG4cogGt0SF+AOm52IWbIuLAzU+R5Jbp2SHSCU6AqrX
gJsvkl5GY7XINGNn/rz5Q2sKw6LmeQxk+sey7QbXGipX8AHdfMJfXSBQAMDZ
dvCkMiqvtEk2SkP0C3Qs23MMK6jS+cgYuHabpC1Ivg1w4mcrQkUWdhHPK6yk
HHb2oW2pGfysmRugX6Gft4XYhB2KW0n5+vl95X8CrUrCkFrE8tBa+GKqkmgi
0rwlsKzO3brytuD4GI3wdQ3JMgjGswg6m1XMgDh0YGQeq9rSL+7R6UFfmB+k
3YXN0IuzpASZn4TqOlL52zQKRjfhUu8Kfx/OMPx7uybF61/aw0sNpI+KDNBM
5Nq2PLtJL8wF4UAhSuhRU8EGrGwgN5xSvp9mxtmvreNXl7HgNXkX6EfE2GGE
nBVXi7k4r4NwTijNNKhAbKAEuE8+EZKQpkWJhNLv5Z3phbYRQ/RC4PMSqrUi
s/11N7sjUP0J58ed540Vi44zvWbKnxYcWVqTxVSuBtXZ26zu+3hwc76edukB
zWk7nrtcZTS0/iiKgkZgAfzj3hNPy6bhqUO9zNea/X+V16YmggnRe5Dqy3Ne
h3O6Y2WKii3OYqHPOUqLljoLO2meU82VigXLukiSMNG3eQgBtAJ5e0KY7uVn
DSBABLNKYLC16wecQB55WhXQR7q4hNaXqLFtNqfgeFjozAmghJdfZtqga0Ax
aS6DLzaGK9CZg8jum/C+JyfrbMrb6iLUs3le5u9hCiAlgDwO6z1POl3Or7fg
71M3IlmryWzSyRFe2dALBr2JnOavuegO2kTonIChrEQf1aPjbeBZLDepOarp
4oQ3pLa3QSZEQJzOEOQ3sKhmlG39fDGJoAtaMUW0Hq6Lz2l8jKLzQbMidODZ
iFnh8brSqFEzoHaOe29wGJqqkwszRyc4ZRsWZWBNenOmqFTJXR8+SpGCPdZL
l93LlGY2cvDhL8yW3NvnF0AsPZ+WOEx56Fmp3bIi2jlYefdDr2vC0o6v3TxL
oRtdptz29cRdfeA3MN56Eq0oxJuJCrQh2zgk+BclL/2a2a6/AuIgTut6BCdi
+bJRepG8qkhZUVwdrHdUOr2kJezK7+oM8UYBv9bx1XagK+3m305GpCFZKJAj
Wn8GxyPKG0BgqCSbMRE5ZT+6IHcac+ingDJUV3j2LLAjaOWC5J7XUMDZr5ZC
S8MNJu5wKwQs6hv44gilJiGegd3N4RpUGv6eHkYWvn8SSYMp4slhbZxLACb9
MoasOms5RvzZovDneBlS9yfhM8KqOAm/01mEYxvwkuvgihGmP+WZqtEKbr+5
auKjmE3cRfHeDpDTjC8/lzfrNvZfZ611Y84pLccf5uloHaftz6E4oISm7Aqt
adESXIWxUusPe83eE1+1i23+OctK6git+dTL7hyPALQdIgsYSCeHlpuqTOAm
tMh8koJBpK2tjhHtGcGwX5qUD0LMzSojgh5CbMXWvCcPZRQ/o/dl1SapCXOD
KsBBhXCGjpLjhDHNQNDkW7pEio+EHAkg3A46fulZ2FoC1wInFNBrWDwiX4dq
dpns0ovMQJANrYKSZvlOxnLR0BeL/Cir6TCor9zivm5/sInqadtwPm15zl2H
+f2+imh8/fSI7zhfrn/n5Sg8tCGl0FKM7cPjAKx0lWn2vTu5dV0UNIyZ51By
FCDxsUNR+lrNbXH1JeT9OtU/Ltz7umuSYCCrYGB8hixZ5O3JX4DCc/lqhK0x
pNeHefBrDNx41xWfOgYEgHjH5btGyi0bKflDbPS7spL91dW1k6VJ8VnZnGQW
+Ss8VR+sGrCeiSzwb65dskp6ZPpfxRUqxtKiedabrmrhjeSUt7+c7LCelQXa
LvXg9HjSvzcd+285n6gu+/czh0QRLRTmbIPhM5rysqsvWU4fUVdXpMGzzTma
yzlbtiTiUtVi8xZCb3xkRz5DkcPKNbIJ7j/SlHXEw7FUbo6u+Fr5juOZZosI
loFqDTQCAnEB84lg8GrsgP1bjD0YNX4oKOVmnI+qNBotnh4vTBF9VM5aiQ9t
NB63vgzeGQl96bCjyLQ1GqxnXuWc6w5eQZSVP5i712SvQ0k0PmfW1DzKWZww
CeRDbZaj/HhY7508OGoOT1I/QQByHjih+WnjW0s7Zr8r5GPwhorXt1ChStJZ
uEgvqhhDG1mKdex4CfyF4ydc/5Iq/ZwPnTM4JKEk5Ho6ZnM7mpDXxI4zUVHg
RHEKtUNh5XmW8G+Z53jv1c8J3qfKfQT9OOIA0EdhsWAjDtkItfNWT5+cF1qT
Ad9XzpMOySOhfPaEHhDHv1v4HIw1rQM2OhvBaeXhQwnG3z/y3PZaBCN2SaFI
2o4bhbvMDOUsgFwiwWLFo0n8Ev2ZZO1APe6/MEXImnWDz2BfbY/6NGL4DHcX
M53xg3rTBIBfS1U4I/z40Jqt2AoyOhd5ofW0IJFxk2AhCklxQ6dK+joP5nEb
+Nk+iCLvO+d52yodXc+P6DUffCDDrgGtmidNRXE1GtpnxM92pmVtQjz7naPi
swiIHcwaXYqVbTaVzqMCgDU9MAdMvGbSIJa47LXKgQ+2d3FLrev9T9FmXJ38
02HHjefuVXreZpvR056CiZNTeWWL14QKD4NjGNYxl+yIESZBaERR+e1EqSq4
06VhQup3FC06jRls+wl9Jamuwej2ra9ihoi351xbqmP/h+zIWGCc9223l9kb
GwlE0luYcfLbCE4L5DiSf5uk3yVFkCGBFxWoV0sH8WCiRnAkf7xkUWM6n1DN
FavsjiZ09wR9fJZIipAM6xsyd5AsEJbJlzjxqvH+LUBPH5yJWtfgvH6A+fLj
pBKuhN18W4w5tvazjtdvj0+ObtqPzvaIQElLJjYXt48eL47bXvLpm+mOGss5
MCf6i86g9LUi7nh7TLUQ71Eok+gvw7NAq1yPX5EwSjjkemnmupyic02aXB4f
Jl7z0rN2wmJI7GOeR82B7z8Tetl0sfgI1E7zH6mRcmKArujEvsUwnaAvvD1J
5XUe/Kzpl3xbAvTQRB4B443sqqwZklTD2t9IxUn/jotuinASTmPDS8vdsECW
WaGB+h/737+vPUC7i+zDB0mjdxdZrp7UQ4gHBpYSswpNLRc65rbt0X1eKQ8g
nRhZbxihjhajIaEGU9FBMz+qVRcv7DQ6iGHZUVjMlspYuU6vjkqSp1P8mRbc
JgPXdVX+e/tOlNVGF+syuEnykCr1Lv1P44YxkekVvKlNzqJNnTeHsUqNJL1d
TyNWNtYoknB10X9zgxhnBQKpPxIUITpQmKIMQC5xfUBnqqzPRN+RcITBWSat
VzegqbHQLXUE/yqMdL1okacbtbvvx9V1Tzw0d6Ak3o7Csa7mMnnwfF4JWi5V
3eg2WABjHxa8YlHhTgqQuj+jUVcuCBsqi02l/gSJ0dyZHX5sx8SruHKIQ30G
KkXioyF1xhF12H2P3mw352wg3XZyWGik1kTNkYx2duoZgo3hiNALpEB7e8Mf
o1PyW1DHqTT/Jj8In5oNDNDdNdBAbjJ1vyRZWbu80s61Mf5yIjvp534qqmQ9
ESKiKKJ52/upEDotDFnhElsHoZK1bAcnbbAwGjmlOLv77cN6jaGE4qK9HthV
/t1X6vZcGadFCr5FypCLTnZAoI+87aI3UbmNx4utfEsxfQCTikKPTMU8y9Bu
+JppS6+/3tkRR/cxF3WOotS1Rj21EFJdj6NteoFJKSZ9q53bLtC0xGy9vmv8
r//1+C4VfEcZ4r9v2CROlnWm5JabtsNd4SOHXBb3yxxbN47q7OPViQCb8F1l
4rSitlLcEEIjIyK8i9NZTbjg1k10buwlHh76I7iVYA68XNfrvSuZgUP3Z4u9
tdLTNkcuEYlxOcRJ/n54if7KXHu4lx1rwzZJCHtvIw6bo3s91Q92quc5o892
3BvRp8MkIZ5yitekoiLM3jicfU32609tuD+5jkZ892dSRoFnxkvliTe6Nacl
0T+8j5z2H9Mm/puy4FqpAE4xRpuVL+h75kF2SYUYOd9Gck4U+RkGxbKpiGyv
mNfzeCqQFF7HtWJPc1ceCli9fZLfY/IegivYDKLNpYVlinXTmKQcTkWf1BVr
RSplFSVuXPhEZdWfgmtu1fprU+RZtGhSTa2VWhQImNcypeBAs3Ty1EtreKZM
PudrxOHkeNGsqP7cwEOznQXI7e1HaHLyZv3aw6HUrknrgO553+Cl1oWmKE68
63DLcDBbQteMsnuJ8RyxY3wVgPGnH+vNxK8tSWNJQdKiLV88K1zbRmn8EDM8
8a9RxS7qOARiRV5voOQLjpUEC78NsDTV/g0Cc5BPpsK163RDrvFTO2Zk9S9a
z8ajOVN/DfCt76M2sic4qBuegKjuzSogoS8yyBRY9SPqegb3iv+IKwjFJ7nV
0lSMUERjiJxUdaK2kKn1wlePYVkj2vAee13hq6vFe4ZUWsQ5qUpi99NXVi9d
Lrl83hUJfW/syfyT0fVAIaW5AAGs7xnTire/X5Zr8gMrL5CxGKDiLb+cR5oL
Je754POnT5f216iMRUQ5andpK6kj34Xcb/6L71+W31Y/hi7kPtRhVfVzB+mx
FYtkXy4HDBOp7iMZcjm94zORS/dDD6QfF/40dXi2quAimxDFFkDI/UyKBmqu
qmql+ibrcBvV6HCEfEdsz54dfVNXFX5GQNAy7K/I+9Zb/Fc2H9JU1N0b96iJ
2K5dYxZp9tVLaRD0ya1Xfn0MAovlnN7LxYF8G4cls8bhuAj892EsqVa8UzZ3
tzDH/5A2esRgLgHA5ZBY0dLvg5f/Rvb+fsrLQ9z8hfeLoRKIdcJ0ExR0t5tP
i7NcZdTh/Ci5cNMz4w1U5vVhnPVOd6N3xzrOjnbG6Yrs0cgdhbUGIs6/zw2A
cOPAbc3hQ7siVejy87cXpg2yIrdXSqrq/RukRzcKnbnyzBk3vvNjlOQJCswM
5+fQLu+qmrZ8j8oBLXbco3QESMHu8AFvm6VRuClqxgIGar6FXyCv2MxxC+Ep
wSLrnfW0JGaaXMh/fa/IrC1IMj8if4y7CMhy3SB6V/Muc/9d3SISK8RtnvNH
m3IvNrf+M2oZDwf8GM1+Yr4X1QdLtqWWKMoMx51hHfncD4bW2TcyvSKBIPVN
ANVZz9Lz/jzX9S59jtHdlHnY6uCz4Lw/Esjx1UhtSR022f6HM6Cczom7ImcY
pU2Y6zWH/Bu/t6rWrgQkSLJXvt6szXkmczqNu4o1vIcooJVZhc+TVaO7y0/z
WOBZ/fsGmjuJG+XUgkP7Fc6v7tgGS0ptIYCBUseEz3IUqhEgWHWPu4/mSY+P
44RO2rzrc+NMoncfZ96ZEH9HmXe8vvnoD4gHkFkqwpONBHCWqhG13nx5nIuU
qEok80aNhDKi+Ki7N5508/d1mMUlXFjb9VOLc5NvEaqyCm9Wyo1BRWOhtwZ4
JzTpQuYUpQofN1EVXcA4jpfmHZ6Jq+ClnCwgo8F+Plrs1+I9KYPtQOIOgxFd
ycbUXDk+UtFoFfFpo6TI+EDkfkpQq1IM510Vir4uEeAg6YZ9h8ZFyGVWADuT
KbiBx996uDn5TZ6sp9xldYLB/zS8IqE9XtBwS8p5dQMRLVR/GAt61R7tKuRW
n3AcMXCrqiZdHmynmAwevTsXngLpI9jLRZJmVwF0lPkvbIl7NuMeEAUGPV7h
2ZvfDlQXQRXvRnGJPo+uYtKOFKfZoq4Y9DgTIoC0I88PsK/9kOb9U5Y9PCKB
/DKm1FGMj2IReoKlb7Qf/Lo2TwPFqcwMIv+da1SRFDCkvjwUD82T+eAK6KfP
T5oPOP5dhNo7kPpjshVtBwKh5FivxrBhNWLOPOOQf+azmI22d1xidEhjngB6
Ap23vEMmvmzPjChBEPN1mH/4BmQEVZxTfjXt7rKAIaveRlTRMr3PNLUzpUGz
wsrXVSCcXPrGB3ch5Nvk5MEGhpohpDyWwnnY6vcPuLr4aYqa+xOzD96Y5jKv
wjUwlIVArXBmE7aOnoOUZ1RGmcgBGNZRgJRwgmDaq1gpWOqg66MqvDkDnIyP
DAvbiccxN6nauR7uhv2VRxrOhNqtAACswoQECbykPmjlEeV0ZUX+JmNLXPu6
fWHGI/i041/HTF+rbHfe0pnBvqfZR/AnVS9xCnPRB8SdkZOlfrNqmSnuQjBk
ht/bPtowE4CnU+iVM2xlPS5nCPMMNZE2rmjUOKaobY1itkFXPHRu+ZTtkdj3
MyLd6Uw0dZvYrFv7EfMBkFLrdNIiOUMZj8LWqdcJZ+BQObRYlih6odRMzX3C
orn9mAYXgENJhmVfH737/go+xh28HQrd2ovFxWnowvLhFyGlUeaRR5bwQ4JW
oJNrhK+HM4aYbrKGJBaRbuHbWCk3ZTdwBYgYKO3IZz3sdkMJItcf6kgG0ctt
7cBpTKUtT5Jl1saWnmNGa2f6V7sz863kFj6WQb7rznZ7vhd0mzsbATNsVHkx
gyoDJ+FEKZopGuaVb3HVdxi8VNOFz/kfjrINeZNFJ2wg5Gux4Kb1KRvFPCRN
ICaHfUca2IbEl7Os7Y0ccMr6THbDq1uqG2tKTNDvho9IIwFV+0mM42QHM4/8
HlBNq4tGpzUa2m8e/5Lxn7OSaPiRd8Vmw13z08M6NhEe/zKlbDUizVin0ZHR
7b8+XvqFXnTJ97R2Cg+lrUsh5VQR5sZhTnVIj5Bo236G/f1cslRNdR+MqfUJ
49IxZR8KEicToAIqBO7mG5RU2llTJgtsAYzxH2tEFGGq/Y7sPU+krtd3A8nK
tqt4OJiFW8418zEmfaCGQVUok88otrjFy3C2hXyb9SS9xAWNdQZ3eit0PNV/
GUUYPpftKAESi3+sznhEleazat3eojoFHYq6jFevZxC5d3bGKCQ27pt787Y6
CkmnK7LTMvUcFYegqVyIjleNPnyGb4kW0yBHXDugA5P4Tan6jQ0V4km5/Nkn
NUAKbiX8BMqw0stHy4MexIfAiKb0Rdx3nzFywrPW+evvnLWRBVRrIxBx2O33
ZUU9/yjW5Yh87yjiJgaKwQTxJIEXgjCBpKoy5fk5YMfRnBaVGbUZzvXrWAUc
/AEJtC2AA72TQUgzSuloimlkn3d492Y4IhSkp1dL9hAm5zwGXCJJ8BVYcGcg
8HOX0woWyr2d7c387oPZPRflY3NvJrF3YV3z+7XOZsbt3jIcvDHchx/kP1UP
zOxC79UC2stAY0pbo5BvEYX2Cs76gRWuYDCj9Z3GzSYE3bbDBwReK7WyhEYE
4/+n1O9zLQvjdM/IcRoeTyg1xeFCKJKHg/J124iZaw95reAK21fxjTCSr9BU
qjsNkINpH9SGXu1plTQobIbPkh/l9YTd0yEQNnTToxechIzafcCe6FsUeCXp
naYaqJyeUIzufah6sS1tg8G6ZOPwmKudBTXZZCBds0kreh0WtwhcqqcKPaNa
F8r1J756WRdMsjixmZc3duN8FuiOUhGxRT8wamqc3XcbcX7uir4V3F9cQ0Ne
IPrW6GfgtV7/Hc+zvJy/2HiTyfYY3e5nOxrsOliQ+wj8E8lQGno/Cbk5/dzK
3PaFjItVYlB/EpAfSXlroMdR9DvdT5XZFT9BQyq+SzrNFsOllqgokNRA26rW
DqmpQOXSWVY/NEh9h/7Ukd3RR9dBsIsI5sH3BZFGyId/HQ3qQwoYBCirRmms
88ygMqVFbh90rPoiHI+XI9rEbO+piG78YF7QV9pbhjg4kCtpp9VAwaAgLDuC
N4DMlXYMxpyOnk2A5NOLuydJQ7/KCTGjPRmjbaCV/16EhzamPuBBmwxgoTI+
I2j0z2kXWPWwxrOKkTnJLOrKldgWVbz6ScispdiYsHP4Wo064uPmTegDKtnJ
KgvPvybTB1W7atmNVZbH9uZnep2qaJX2Zg03e21Oek/JY5A8Ia84Ss43juZ1
V31Uq/e6HcrHDTxf7LBS0kcwzBlQtEMd2gub/2Xj7sEpyjH0YCgbRakPs9Jf
ZE+bwEHCn2NI1m50LajiGDo+7Bi+qJ6qB+fgrDnaJcca4umcZ00g1EXkH9g+
QccFM07dPLSnUkMCTz+YsmeeKtU7JYIxcmyKtF7QMP6gDKxxhxNlQJ3q03QP
yD6MBLKFcV8yv4TPrnhka3xjYOmuRdJkhMFDMjfXtj2CEiAqIlaWmBbInqDy
z+yk3mqy5WDB444M3cJvDqjCnRUgLdbUzCpcFtI1V92FE8L3UVAVmOOgBEsS
NHohmqeTdgurCkNYZ61EtbBuxPyeSC2Wck106EuiUTQrm43Zto96ofKaGQPC
JJyeWvkisgwRbNG8skb9XsIILQmuLm+hmu1w5/J/FLjmGtfc6uW8ZWA7+SE3
I4Pgy1Z/vDxXjKQQWWVwnLp4JTkeKyi13B6n6GcyXTXgHrTmvHtbBIMGEwwG
tJeAFUkXjpHpT5YKBoV0MYBczFzj8oP/WyfOopR7+ox+7Kv1j2jrJZ3NcwIV
/gqFDbk7HvIXppmf4F4Xo3fq2vIldp7Xg/1TInBrZ6oMGdix5zp4mKffj6GL
978cjssBOK3F/yiLP9nyQ+odq7KsO+c/96DmAis58CJcT3KiuP5nSS7KW+lQ
AqtApehph/rTsMR7dqfDuaQEUXS1cAlANPrIt7T6WagZ5xdSREOze9HbpbB3
jvKejjPTPXYtCrqY1/ZUgKLAay/arX0EuCv1DlywH0ncqvWVlobK3B8PUK9W
3E5tkR3B38u5IvEriVaiUHoUhJ42M649tBis70UfNi2Qgrqikn7IgTPUAmPB
lOwbb5XhVbuREt/nNFpmqUyw5maMVQaIKPz4BNzT7ws2LcQhJrMcpw9EgQoc
FljFo/v/8IFbIcZwoOC2PzoBZh9kmN2nQz2a0pJ77RiIjsbVySUmMlOaXqWn
Xr5+QLZJoDUciGg9GekBAckaQdz54Bh2w/d950IWYIGzmeyeMhIvEAOqHb5F
DRSOnFz4vW5tGLiLYdaHwus5x2KwkRw5lR1UGwMxCDJoiJPvbENJPKlu+3z0
huoy4L8YEVItxCdWhXn0nsZGXaKHWbMg/6dS2sSmNYuOPp5b3d5z7NlSzvsT
yy3vIHfEjXM8YejpR+R2/o9GlzQQr+RxjNLjSK+LlEWcS1Kh5SkV1my3Ib4k
OEjazJd/0E0KQkqDPaEu7rR/h1AF6S4xjw1vGeiQ7OzU7OIdyRdutoJSto68
g5YGbQV2mEwGYTXfoeqbBSI9NDWdqUUwpqRaj7yBS6zo7uML4HbS1WmM/gau
kl3wTUi9RLf38GgnCe+cNIwBC91TPsL5wJeHgAC2H1GKnMDAXSLrDmEAwJwy
eNkVk0FeDtboqKhTaH0PHTQ6NyymHRR2F7Jt/88rB7TlHS/Qa2JbkhHGJ6Xk
A45POI8xQj1Nts3fqzE/CI2u3auGqx4L4zXO2ZuN2i/qydO40YEvwRVgC57d
pduL4yrhSL4dzkGMBhHNGy4n+87ijndXPl4J/qSMfXbP4OJHnBy2S+4efUvo
LSekSvGq+l1XoiqZ++XojjdLFxFy6SqxthX2SLuDlsmTgH3rjgHhXSGZf42s
rxGxUY/FwfvMwSCSxQsF1+rJVs9cHZTGrvXTuv+PwWxmPe5sVPYBRKLdm9T1
53HPFeKxRm2UCTxrTaI+3WvVqv4P/0SpZ34e89PVmJZMGFFQQ2fRtBSciGWI
8VOmey2u9L5o5YM/OpShG2NCz4HfM0W/v2ZHEa6p49fLTFbfJPaXbJT+1SsA
F3gcEBDLARcYrehcnXiBlu5CU0hxx6NjfGSDtLV6475HnWDR67GAI2JLIn+l
BjBoVLlVDMiJ62HxSBhuKg1roX8kOPxdP+IaBtD0IxHAQ+kuoIUk28wq+zEQ
yT6dk+DIqPpy1XkYpsWLypc56Q0QmMESrC8/pj0gbDkaNzgyDIWl/yAuNENw
PZerJKvNyfkDs++nZ1avnMGGX8ZQDZw2CAEBC3cYLnx7/G04Rm3wMag9wt/c
0YrjgzMvnTXBWdsInZKId4edYtRc26BPSfYpGlFbx1Sk77kAKQkjEJrjXDsz
a9LiuadE1rYKMHUfEm6l9KqBcGfMQ6YQa4ALlyjHz9G9USePQ+U8MZIlm7+I
v0clm8seKJhW55zh8AJxDS2vPvXRNPE6vSIy+xqx3WLrwv/goJgKaCY6PDmM
8hwhRKc7TayE0HrdOy+1FYNg9NeRd8YlmcAGL+/hiqRpi5EJ5qJxSsgl3qsT
KZVBs7Vc69jzWBxNiFQ6WJEtkKQGzgJPKQstavx8R7B+ZS5nkLr7xu6yD+G8
4bXFEQWoxREujLobjNjGzn0hZsMUhUfYydFLB5za48NyUXByzoP7jAWYIc6H
QsmOrGvETqCfhoOd42dfFoG+SOfJ5xyR9nFcv4mjjM5G1AuaWA+WajXDt6tF
ND+arLlcF9OirsLvXHA85AeU2O8vk1y1am0crFTZhp4Bri5u3N3Ra/IhB9o1
d6cDGXD0EnDq+hWH45Tjv/+UFOP1pyJxMsMv6VxmNz4xz7f45JgEL0zXO0u6
+GB7GsO1XX7cGuxSENLh70wmwlugWQ7MUjLdA4qJ/vAcxgWjJdrhQ5mYHrqA
amYYvSbbPvu9VUNjGfKStigudFOYPbsDHCMS6Go4OUaLj0iFBx6D6qp1/Tlw
KxyHTfq1gQsab01rmxXOV1vj/TxNOgrcDHl/aS5YTWeaBROZZAzLkpZP6f6n
tpo0bl4kLr7aKkOv8pfunr3/X4JDShcZdXC8SjIEG7bSK6EgQ5beWALeiguZ
AJolx2/b7fBdHFviyJi+bqumqKGTCHlwibgyFZAy85tiDGZYFGCYwvkkHNvm
/CEtbD0V2mEaaNG035qBA5+2SFbzl8wVE+qp+6f77Mr2YKa7/b5wM7AFG96v
GtS2s00KpXoqslX+NkSJRL1z26k7UUwNgejHRP2inr5vshbohwX0r2uuHdc/
hGIbt469HWXar8RsH53FXv86g0HnogpHUJ8v/bbctIcjnTHRVeoE6eSxCGrX
L+uUqAXVQXeTYhR86W3fw3JzoOOSYWVWqRQmcSzftFkj2P7JLQbxKd0JKpAj
QQebrjEypf65zLenCy145M7835NeWv4odkw6wt40HApEIPpwcIP0E7oOsaDn
4MeBO1ti6iOCxetrAChrechUIbLF56WjHKMmTwUZY99mlQVp6srcr9kYIGnq
10oFTE+c6FxGYywnY9jp//WRF0oinXau8QS6gf9odi6H390jDZURQow9nqpc
5r4PrnNd6OyjzJgYiVniSw/8xOi5+rpXsPX2hXoxKJwIMGmdILX0YqGw9tt7
NhJYaFBGwS27HyZffW59Ad3ddd+s4lryMHPHk0XlS5P1tPsLT5nsJTpBUxEi
zSj1FIxab4RWUGGHdcMOYsQeNXQFc9GTQMK227oALDqK6Uy4VaA4lD0QWNiY
35hIELrv91cc8LTMtj/P85SM5qWXq1kdW5f5C78NlXo+KLWMt7BsSVebADVf
o9B4AYhlu6k3+3c7AuSBZMOTzEDnce+bo6kKQSE3qQ5qm/bPHNbdEFqCvLto
z31yqPJNXUA9tGNoYHyle9AMNsonoyp2o9FtRxrsoYQpqYq8Pac2wrk3JStu
H6HhQpPKCfX8EAmYToVcM7G2PM6dXgUtP8+1n/lRKQF4lJ24eZAbHX1+u41i
xeF0HPhfT1esHgJDfUAC2b0HulQzh+I5uXkH1VzsRfYU7h0eBpKKZSqCI4Sv
RF4xxF3kaUPBryWmT9tVKadnC55qQ/yH4+Di8fW3UAlUsvKDOxsvkHFEd2Cl
A7ZKczM5SNBaHmdaut1gv+0aZFuZK1of00E9P93UiCpzgY8xp+qvP3XbcVpl
8Mw3YB7E8mbXRtWkR3wx2rG4C0SmrM3eImqUtwQ+WLp2t4C6ff/5Wwd2assh
gVRG99feS/GN/YEeLETZ3sjEHmBwCfLuCqUqtjGQYviSq2Rb9Db3ijtfBuuY
/8naccI6Xuk3pf/uA2LYzWuybcHKGrj8iF1C9UhtP/LtHly+OAyn7eRZ6KMv
dNGvWcIbF5sNh5zHkVdFoCSNsFJ5GRWj72lD2ofW3jDN7xF0mMetmHUpUImL
Hx+7hvm9r9ZbKWvABQdj60VRNNdSogRUCQpi8DV640s1AntkSr2reHymRW5l
52bxA0uV53byCxG+1xDOrgpeBVnln4Q04qtkjtEVqLsc85cd430FnXEuwcOT
S/APQD8Uv5MTPCWsxmWifQLNtcdfUAbIj8cuttPerCik39bsGXZBkzIcaL7e
LYqNJWyO19kFzSrKAeHw9ozXBX2P4BcrU6jmGAAjV0oa2vNO9Ww2wWuxoYlj
ADQ7XxjYqhoGWhRx8QXR5OLGsAO9JQB2vitzViX0I+IhmoCze/KhJf554rIx
uBR94iEjlNb4KCs+UpfSiyimOJje0SY3o1Qcsxsl7qcra/Ja/8z101HRhM+k
slJGsNLtekO94zXMbz1e7UIEN1Py3GtXYzwph6JT5Qg+f3nmPIz4HAqTb5nZ
evplVDWX/RxZc77B97W+oMFkZ0c6zjSRsdaQB5Bqii6FctVvw0sAOXsDZK8h
ctb+tuR+6/j/ymSz9WuD7b6BG6EJGJuYvdZBh7DXzcRwz8DjIEk8oVZD9+34
zCl66IRn7uSBTQruQ3kQs+EaxK2UOqXQHTfAkv4M8lVWPivNIEw3A03EU1/p
dl1TiIUm6MF4YXCip0SMR24d1EqLE32hcWsG7/yJQ/nOsgK+MWq57MVd1EDP
Oue2kEgyApSohKDmJMq0WJ9jjxGXtrbtG//y8qeyGcmxhQSFBu/ghSRE0uP7
WXxiH8n84fifAEJe4yw3KX+V5JlyzjFsFKvxL7mq+O73Gkre5EaHLbX1WPTg
fmSqLA6tUPloT+MRrXfiX6RQwzHi3QDKsCwPoS+eIXqgAnpMT7awUn3oplRc
8f0NFo5X43648Ek/JzY8GLeKR5CkqPeWTMoBy7sps0ki9ourZHnFVtSeQemw
IhXVs8mE2CleS1jrJDwjxbHvxiSMp4AS4oItWp2MHEdnLwqqnHUKkvKp52CR
UEAIugmHej7KkrS1/q9YOrNBDzpWlrZDYZ9PMvQi+QLiU/d/Krsmhncn2qtm
0XSl9pZZxJbYQ3zm5au1iZgqonukwFeNq2r7n5WHj1f0BwHMI3Rh3h22rNwO
gZ5JFgupsmW6pfJKzWp7Nb7GSfVmNUt+zG6cv4wjNR4LZNBeJ+7Gv3utePIO
MZAKRYTVyOgpij6RBIXE3su6Eli7TxpgYy1vJVuy83klk6qU44M5I4O3lNGE
KzbztlzYKQldBRkbmrL/hg4Zjj4+TCqdis1U5e++wHmHeKB7CNktceohn6fq
vk30sWAG8/X/mkz6j8US27oUlBYm93r+qn2g32Xki7qI0a2VEwAPV7jS1Ckx
qbPjATKsVr5wmLcE4Z1paNvEUXSZbTU31L2lQ+emgpzKdlmgO3BYuaO0a/zC
DnopwFqUAhB/OUn1GFYXHD1GlC4b2h2F9bS5QJiuZuTxt5feT7bnASBBLigN
v4xxXG4RAF0Gy1aSEW1pLb2nZ8OwfZIvg8RBK5ui4WbgVDo6/nm89L+x1926
U2MOFL1D2SddzhnLmXrfOvDROcwaLeQiYGzOqFlj8UHw62jbVfCltVVUwZ8d
PmpD4iXwHZjBLKbx/w2ZHCOuHkQRcqBBk7pEnrqB6PLjbpvT7X/UlFjMgymN
AyTUluemf/5LvwvUOn7rO6GBs0LRdNCtWsVgg4KmFsr9byYd1WlX5Fkx99L5
Y3Fvg6P9JSx/yKi44fCD1K/XXfnsksmZ3jnOBHVtRl7xNeLxjPMiclVFh1Mm
uIZlqOOcfiAcc3tPB3TBNt6djcKG99EUUvYHvRCG5qU0zeYhZhqy7ESucQ43
SCSpVKxEb+CxfUyXRePzPE0WKuLXPlGLSYYy/3EtNR2PRpSOowKb+s9lLH45
MufrlzAe1YUeJzPaA8jMU0c83D3ZnCiBVPS8LrDxiqjFNzO+JA06lLwgtZT2
rZxml+0OBzYAC1BZkFP7eerfxtp2lIfY9PIf14KVVKGd7yKmzTvZbnXN6LK1
d0AHMy3ztWdrHcG1Jd48+VVk6HLUqeXO1AVJCYpg8a8peppjsK+z+ggQZ5KC
Iih8fSNyeLlu9M51yDmC0KzSqQLtRslOPVtenohWA3rIyaixOcrrq3vtDyfk
Do8EwYC/P8axRmmtEm7uUcWqlo+K2MEbMJAXPjGpw6aV5EMKbJ9fQMvmcNcD
HkLc54X5Exm8eEs9+NVjuTT1eAHXoLK1B94J/heXIQ2QvX6wlgWn4JC+G9s7
eqoWT+aMj0/DkoCNzqa6Wao++Wly3jFiIZY7sHY89Ak4S24+lcHVB00oQ/xo
Dh4vZHMBzfODdsHTzbI3+PMWrcYRnyGmTFL7LeLdqmXL+e6S0yp3WSQdqx8/
qWNgaRkY4WNiYQ7tKQgTKosyKg/PJo5EHOrsMpgkUlAEJvdHxsKr8NKJz2yD
Syuq9t3j+RffPcQJTfkX73yFWbrRRe7Zu+c8wO/FbQGEo4wN1SiEDdvCF5pj
LnmjwZtkHmkzsbMWe/PdlLVcVg1zod/JkcMDBYtO0FiLPmKvir2NFQ3t/K+G
NI8W4EunAEn2EBttPNSOV1bV+p5keNH6Ui+D46zAPuACmhdr52FLRPsHNvbE
NDr7Hdy5d6w9xUqLQHY2rjNol2NlsmBKchMLnlpYJuUXyr930P60GYcUEVLi
juMTGYH9ziltG27OwFZGCIoz6mdsCB3rC8wx+IyHrhKENkZbyhsqWP/4z6nY
mLntBWrWeoVPhBZCL67O2B2zPswaazHzxJ6alNs3fYUxKz5neqbh+mEmOZVf
z3KAnXAZYq5Wmj5w1rG6P5mVTGQPpBbzB/vikZjZseiJzT5kKDUXVgUf2IMw
0KgWGlwuu6aOQF2IBfv2Px8gYjlYE95Bu1S34II2ZLYHPhBdGhrGG5h78j6k
5jR/UhWpP+Too2v/RqDviEeq2/EBzTZifpDGhUmD0uPSMIdi7bFtGj9IsabW
8agwK9exQuS2QXtgZ+5VKXEvbB1UO4RvxMq4GTvxpo3xH/ESbNfmkuxsagiS
nwLZVegGbJVwhC/IQIq/3jFXAFG0qrNQJDIJ/lnx1sWuIGrcYQbcXzmFTs/U
Z+Y8qGnhE57vTYaUKOMTS0Y/7+NKgBcVYr7vWVdLJEmAZHHdsjCbpodKGxEC
cyIUv8jK9C94+B6EYDJuNS0waMWH8QnZJ3INTtaFlZkMpvpSD1SXbX6oiXuy
n256BNZ8WuhudkFsAUFBcZSlwUYs7FWMJBU399YcL4Q5AsyPDjnoTFzDx6iU
x9RH5YT3Ba44GhkBVmK+fAc+7Dk12VDoz7nW+7nydhq1HMryvzjqhsYSXvRD
pubIGO8oqFh+O2rL1vUM7H9Up7ygY77SCrcsD4Ce/5x3YPMROorh9INYPnq2
Acc1FebkH8D83fFY3wTNy3i71VFkZI3cQWRAUF0M3FaNtqifJz+/atXUbYIy
tuquShrX6otSsb2v+02jiKSL40GTyczLHuQF8X2sdxAGqUjVnPoenYXcjYg1
wmzWaL5D0GXiHQXNOOLM4uzE/6t0eS1GEylPKsbooStx04tlNh4HKcBAxsF2
amZ03YWCAdBV/siTNenitdx6BzSXRKDE0INVbJVO0XsDsu/i9EasJfUn4lRI
/wusu5o8kSlaepWgt9CGtV/u44FKvYNJ5t0/m5xnuWJQxY1uiAZFRyLok6UO
rBzdOlvupuEOheeIN6YtwAga5jGz+aB4HybAIdGFoS8Bbgw/e0q/3OggWdMU
Mzh/pqabxkfiXrOzo+kRyWetqCUUTExCBDRjjZ5BPL4g15FuhZJ2p6+db1jy
1VG21EKStlCog8O12hOh8xcLgVJG5wIpBi834RjPgjPaSH08Z4GAkg5U1pd5
aHNJRSZzLehJc7X8U91wEu9UCWdwlT7iUQ9bPzsiR9YTpuLBa5ZlJ0b94kVr
jUK5XDAKxnElnNMk4ecqYWbswN3Jm/tUstv6bKONdyMzyv7RFI17BpLzu9PX
7KY28qW0hb2Emds8QtxN+Cq4NwAJMr2w6Xc3bf+WhLgoXNV54+ftOUfYbjVd
0OalvSaY0rrt5KZNCq9P0PVOsJb12cLGCSxGcMflxqbJLxGFWb+z7j5H7vlt
/gHG3QFqILW9psdVQK4YaJFG9pwA8B8OCXPytEg+dGOObV3XSbwUfmbqmauN
YxUPflIpCqq/3H1dpVjURS48CmfcFB4xGEneIwRveytQJuSaMTYxhf71pzNO
C4DCUG2T0uQQ4kO4HwTM6F36cS9MOT58wZVpWezqsPwySLQ9gdGy4AxqqCpx
9DUXJExPGbTzNfGe7sTLj1MpLwtETKwnKveZRqjIu+ds4SNAAR8i22pnQal0
rySa4AxhU98Pf/qeXTl68PXPg0PcsP4zS26o4wWMfrtfAlfWe0tRL7KHNCnF
TaubLf1cHkKkz5lFvJ7LJ39YKEhycDoqO5wHO17TEylleamXQ2XVKEd794mu
/yj0Gs+iA5jgQuyCztZN6GYPLbhZBoulQS28K/Ju3WD47wxoHEdPAdWVuX4T
xuaKEw21JkYcWsRivjE3eZUSIuu2BX9rriMREhO8229Ma2TcMtyViZtEQI9K
LdgzLydz0fBgxV1JfHLaSKo3LJNZKQxneIdIfHd0MN867dTrvhrYQfXs3lh5
hcTPMuF8l/zt33mMmz1xn93ofTS3H9jE+bocDIh1ixUVpAvuj5vm2JiiQK9z
O4UynSj2AI7xSKqW7DC+7KAgM5yQf+G2HIY6SWbRDvI+iagq9CRdO3WtLe/T
Zh+Oi0aY9MSP4JYQA4dL75Js7/2czhB7ib1IDUc6I3ymNkkRnnvttrWq+7t8
3ozX38qpjZMAFY8LxJhSLQkxCzvBxu14ipy29ngNAM86W4ltzHmdsd9fIhxw
lE5sdLsZjBvl6srcjJ6QjNqKoYA6hoQgnVHAE0PHocA2hgY6Lb3lytDRKwUv
6sKTCZOmVYHByUV4EisXek7eIEGYHgLNLfRL/CW1wZ3WiXr6tcFcUMq+zf7I
lyZPWDdzrrYuCdRNITgMF/7ja+kvWXFi5zsaBAD7P1SddPxSbFEgSmhYHJ1O
IMP6u3/hBrj3DKMk/3c6rejiFJnh5lJ3JGXlnZyGl20t8GvDglDmSHGD0A4d
4VKyJI1nwdpiueItvGiEraImZGyvJbBV3jpHHb9iqbf/rIh0GopZyaLqA2md
ltTSdCVGkcKJkIWa7gJDGaBnZFOsb5CdPiZN6GabpHn7JvM2BvM8z/hqYUuF
WxszdB0AeVh8oEn7voHj7+zcJXwE1/Pm4Vvb2EoMZl9Y73HODJGUEE7UalVN
EqxIZ7vURAnRS+g5e1P42hhlDdLAUduLucziUmDGfi0DoEiXbEfkfUVi7cAa
p4GDiZ+xGU7yKzNyeM1WjcjKWd6NjqXnCIbNlgujgpcbPobkLkPPTReft4UP
JfNxkCuU5Gt6xn7eQVlRoWzmk5a3N2EymCV9Yt3Rirr6occGPugwvTfqRCU6
SepZnmsUD+GNUnWkUs14L+4WWdZR/QEjZZiSKkzxY2BJhXpS6gp3S7rw4kw+
vwDOIg4gYjzmqrvOzrTBG0LT3VkMITTQg57scCZOgPCUlJTPmeMGNFNqNxG4
IPI5YTAktYaRbT8e4MfhkjVkUnkbiLHdNRacKhMUQ4Rz9bgYfEytoQwrX5+r
NnvNdRIxI0tYoBmM5gLhCvFAY5IeLjjgpApyV28Zatr1BuWsxKE6KRv1gxgf
vDbYMH2U7G33u77vO9EmekLUV4nyaGYZrzaBS5JedQqDtKfQR7CTeCCoXELM
id7F0F1jZSXh/hQHZoGpw3uIcsbBZLexAzy8yJqib3uoWEmAe4CPH5g3aWvh
38WgpZ+KyffeV+FHhHTgViEKyStGCfYxuY5ud57nr9X3AWlIyOXMdNuDWMLW
2J2PT4mu97uYLNsOqDph4aCRrweWOuFiTTVyjOa/wZWWpF1s2gJuLBog47pS
n+JNY7wWCjFJ2lw3hGKL5Q1cdX7gFLAi4Iu4RjSS1MIwxAgkfHQRDi3Hw7RU
CbZ8RdDlatwFvFZdb7ICVHA86VpfqSmMh1/Diz3Mq/Xafl+gLT79O734oKny
8s5K+gH1A5weWzpIBW7/NXbJzBE7IArCfXRac//ur1mzaYtpccQp7c4bCAXN
GYGLjhp+FzbOapSgQtRpm2wYjeLBGuRjDzQLjeXDkMVIpw8Y6MOjUPD9eR7e
PZ2OMgsLOgk6dvFL8r4a3HqFC14+og/7labU22bbJj5/RFxB4wGYuZ+HprM4
TGITP/hZGnbKIrY8qjuJk8//oQgDhnXarsVuG1DW1KmCWLih3mEc7+qck1Kc
OBlhyUyjKT4Pzc7BvHRD7fHVUcZCS2MlKyT+ihFCZpQUj0S+J3p+UQPq35pp
ZQWOibTF4bbd1Rwhy9bBG57HiGVre6ArQq/aWwDyV5x5Eyz0Yjlelemk2XsT
uksW9+7/pXa0RRFISKhEgHmOPqIf3zEDHms6DbJ630fm4pRR6pEiSmUv/AZt
lZFr5tQoNyFHM9lX/L4IsJl2Bc2W6ViTv5FYZcHtemNNEQKPxUL4nn8edKWS
9Y1DIp7/DQ9k/p5aNMJV8+JXaiNcraE8MHTeiggiLMTS2z/5K+HUCjIBWjOr
RdUXKVixt6smXS3EmTii+jo5xlehW2rtU2/N/PKENe8l5Py2pJmupE67RWHm
EUF4WWTNaj1/qFdlrUs9E5YEHIGS4OPlKVh4KNtNpesStWn6S/VmrzUCLimy
xIaSPvkG1X2P50YwUL41eTDo18F+8UDaTLkjwn5m/020oE4YbwIBFhzbuX6Z
6VIIG2tyhA5KGjtJaHVPAxdUVwBtvthGojiUPgm5O4L8qboFOGN2lZkzf1u3
pV38vcWuDBPJVxkARrYFZ/7q+P+Qw9ZY3RvJ1vo5Fg7gySZz4tcfvAngIXpv
ZmkqRdMIf11DleOCiz/JRrv2jrcypnFHBK0tTCS+sd2ydTFRrNJMxzkgLbat
qA+Dvq08FDMwKqT1oq0xUHzDPuep64uOJkYypJwyRjnOQy06uCL3IZ58C20A
uxKAcYATa9qpBhFhvUjp1mTvIP9I91yO9+Fh2DC+tDBZa3eSdp15OdtpPGLH
NwEyTan3Y/7ORQUSXeXAW5uUIbv7imae6AM64nx+bZ2g8zY5f33VOPWsXtqn
OOl7ETxgZgpI17QjqNq9lAy1dbLDVgDX/OzRdAOtLbH1rBflkVc3kM1agW91
G/yYmyDDLS/IPXa6LvHUgSlhjSuGCekrv30J9IOwurU4/FxFlC3sfRk2p3vc
n5wOp0LVG1cgANu8qyRyqxCMR+Htzo3vzcB+eJF4YGaAW8voH9C2ep63vaM2
AbAquA+MZRSG/20q3twnMYpqBDPnee1BfkqqBJ0w2l357XQsvYgtJHpvF0Fl
ysj3aIQb6OcWlwbjRmQCBfNfvGWlt0pLf/L2yki1ZvWUIWj9YOlu8KuZ+ibv
0vEtN1eP+KSKvudbu2vfY6cSfS0g0N8321cSKFF4nrck/2X++xJhWIhBvV3k
vPAlxg+evbZeQiyxWMu6IXzvXqUDC67AKDhQX86T4OFUQ8qgrSnSCmMlXZ7Q
HePccBcWUw05eZXSIrlnFl6uac+xtHQ31jlbI2iEOaQ6NcEOR10Ev9AyrQ60
BqUOcqkyC1ZlC11v2kb+/F1gZm4sawaLQ2/JMZyjYXPYbcKdh8czrXU6cQ6D
a5+97BPQW3dNsv5NTpouRJM2XN/D/sGVCUznDXl/G6LM6KmDLxWH7VrUQPPU
cYD1J78ro8Nv0rVbGrOol+J61aQ6X3Kriz8rYaiot3J9QPcqyDyPfLLCxcfn
Y32p0vNclIDFE/jzrCMwc9pDtKEt17PQTE3KgDVRV3mYOOT0xW+vDGygvUwT
DlwpmdN3k3h5Vmnkez9rqsNwd0xGskwg7F/FWfZoaLVXx/M/e6+6Joh4Wult
RdX6lENYzULl2YIhdNbFm04zVDi8JvAo/5wid2DannFcJcXOHR6a+5+R//U/
YMfH9yAzHAdGRDZF2mOKK2L+gEhL031nOtcAEwrgiLYai4ru4slPb0NpK6jK
h8GTb7xqWyU0sqDrLNP2qpLmhdMXGQFjoI03QgFC7kCbofNgmcazyhAG9Zxv
fdSktW3pm064Ed5p3iDwLSMSMSqfOwKi9T3HOrxhOpf1P3CHnLpstOLmxa2s
sTO+wgUh1h/C3McPebh37OMiKIgcRSesqgN7Gz5XymAWKD+qAVjbMeiKcM3W
1nbWE2M8DxKrgClZL4HOIKWx4S7b+JgfjgL3KSVS1q1nF3bbQVBvjUlZ/dEP
2bjvH267K+N8FJBhWhHeSqRYNyq0wUa44Nf/YArS75LfCu3UVj8oEYxGXS16
UoxglgI3nQirRJIxqvj7efMvALbN0DuSus3C1+N5WHfFcYuCN45TcLdKAwlJ
YZvXwAMFTVDMOKgF/uGjO8BFQH4IfsMc0+/balLzZ3BAoQwILkggIKtNA1YX
HD5ps0ltTGx6Sw+xTEdotW2mThFiKh72gxu3FNMO9LfcAXdz9zbt3oa6zM0H
KDujoPQHb682HnJ2Hy1g/LIPcPAINzJt3SpsfbXcaZtAuZgxJTXpqC5aRpa/
IyZYIBwNaZ2ykAd7nhxtuWIJx1rib94rviCVehK+BqV6INgyoN+8wiP8eE5R
whTGVG9dT0T2KbH74eZtF/JVV/22j+1wOPBQNhbWhhufo25BCIjDcmuOWe6C
ICpO89v2s8EjQCARpLO/wTrYtSCzv31P0tsmLKfCjF6UiI2u7pyikZSbI1Vg
7gd29xqPxjsN4KnwCuh5/NoxjKpCpCu5BGBRXWdoo4QsllcMWPBQwsrFkskJ
67VCpNukAFutn9lbsDYV2PY2Eph0mO5Wz9op6VdBgpkZ6sgoIEMOanmM8q0b
ynL8zB6SO5tEjP4rGW3CqNwfdKkXSSFb7DqzFp7oSSZac9+4JjXWxk6un5XI
w0heRbj5wgBGgzmkevpPSveV3h08vjTs0ez8vTd6Z6QnweLM3/VBC4x5iWU7
cyZHPFqV6ovYVMYKaG4PXbLvoWf5HzleBpnd1VFS2zxUwA3U43TTwT8Tv84S
xMq+K56H7BLoC8dIXtadvyG4R4R2lZTu9R+dZhgak5GS41gzSN0ORXnddo8U
p2jSn+zRzn8QXt81YDZ0hfGUqLzxoPcubq/MaJkU76gKjYI/Lp87xxQl8+S2
vtuzGMmsHuI8dbjnBYJMC2Z+fVE09tqfd9I9114x6ONm0LVm0KQMxb4W/83k
m3IBQDwF/6aC5xbKomBiAbpZAYGOWAebSe8BX5IuTRUpqWKFjcq6cKK5b6jH
IXGdTLE274wi4cyqqg3AHNqPiQLZSXuVq3dvUQAEvDTTdsAi/gx0KYEOOKNZ
aMGYlWyAHalX5K6nzl9kTW/vFEfhMmkF57ElISxdvFJSdf1moDteqaml3sr1
NvV7ilWxZOip0yB/gjmu9pw4iSOEL4TgXAL1MYWUMdoUNYelxy9bJona0NNX
38bay0wd4epELM/2RLU3+rgQ/JUVJrVj3EF8+mvZGK0kD37nPoJX6MYLQhQg
soZSSi9rEJsoznzPMQr5F4yNw1Tq9GcO3HQOzqzmaig4ZauAHc2G3BVvnmJN
vBNbiV5PYgj9nLYtEGebRcWQB3yvwmaVNS1qH1hKd8eQMAW89AjWTzPxiQEo
lJLHUPT0TQzZdcZCez0Z2Cq4HwFXxdOKPxfi/LdBKJQIAD7VLm3hA3S59qoi
ynYLym5X8q7LqcbtMS9W3Jdx5612saGy4YeHJjFbrSFw2vFaLGKlwDQouD2A
GULwr0W4t7EID/xzZ2NGit+n4+6J6Hip6hZmThv2KcU4I9H9Jm+3/i+tYCr4
4OWZ7rPyZWL7l3CqwSdtGxrw8hMti8mpAo08paS7gTaBtu9rwmO+7CaQ4+y4
5k2vVTkxydVEltli/kQVnL4KN3MzwO0S9zLyDU09IX11svGpEURtPOWP4RJg
NoL/ZTTW7DJGaBcWpPxaDSd3pt2KvvF0EWk8Er/ONJLbMvRP/WLnQOiiC0E0
7DDAklMY6pa/t61EpiVIDFTON/6KTvXexp28kTmzM+1g+SI8yBit6Ikgq68+
2yz94PxkS8Y6PejP2NCPzcuZM+2F4CIstpGd5NEPOdeVFFFB4qhbidVaWk83
znNoPr38fDQw5YqSBIAiwFTlp2/59W/6Y31ETodyQ62BiczLpPPWTu0UyRcQ
nV+125+RskeJ2p0YzW4ePVFVeGk8D1g9Y6q9ZvSq1LjNrQ2UrLVp/wjRYYNj
njzmjFCQfpA/fnJQmBIPiIuTBpUs+t974CpFkFOfuFA/B9Q8VW8XwKiAmMu6
c+0wOuoa9Kt1mwJi4YFziH/LzpmFj2MibdZlMvo+4ezStXcb4ra/8LwxMK+8
ij38s16FGE0zaRmh1irqcn3R117R4KxHC4ITuPpwh6Kl8q54SdBRh9JGDKyK
vwC9o1qDvqoemJ4D83Uvyui4JwYyg1TM//hlU9EbTazION6mOkMCDzErWexK
IlV+rsk3vAj1nA92S+dzMFrk8hD2r927pquhduttJJ0OQMEzBX6W+3Od7fol
p9+bnSreapr0YygcomehAkj+qdv6qzTQyP+QmrtvmsQA5dryW7umYzzsCbBE
Rs95FSV0quaaM3KLAJ9LZnq18Q3AjhI6BtcOpzrwOIaB1MsMHLeqLz4zL518
zyLhHRd6NGgEqY0/6x0RQQZROvFmUcFUVFHN6PwdseQV6MutYZ3SObCACcmH
iv0vneR/OX1IrB0fVyuFsxB930Xaj82RU1yGiG73qOrGHF7boHjKif/u3IkD
SzC2MrjWkdLtkscFGG/mt33tW6fFAvYMqmDCQ0CLmtc8v5NiiDCxdTqdD+k1
If7ujYNPOpgXA9bUjQuCnkoT0nwZkh5E4U2nLwNXW03W+luNW8i2+C7LC8Sx
Dlyu+LOvUj6mMN+oj5ZIX8fiJQ5ai/zyA50TROUvee4f9fGdPwqAizNfEHME
1NMdob7MKI7y74uxjLrliMtU2DrPmcFaIav/JtWAdYL7ODOnWMDuNfXq/dUS
ZZUltFrMiyKd1rCBSs6miUMb2rs1BJJaBa7b1ORaZm7HmvMnvHBWiAvMfShA
j2tEDZlJ6HMXKi5bAcYtqM0+KlO0D4X19ZoJuewVa8v35FVJ8DXFjO8MHzKc
/idHxn8YdOaZsJ2GPgPzMqph2tLnNq6orh/006W+ZBYslG6tWdz91AMoR2O5
xJo5B76D8IMPg3kFGs4roLDuObIHaJpRuRq11AoM1ZzMj36JD1/qIIlzcZ5z
vuCXLaNyLtOM/xD/nn8S1yYU1KmGDZCwR2jqIiJc1DsBTo0UUTxEjlaqI5zr
J8X3Rzpt69sTJ3DPGVZ+fzPQK/hhhK089rt2Nr2lGMFOIJYQQLdywFhc0OXP
EUEVDGhTAn7fvKGC/y6YiMunY575jQgE4U8OCodbfnelwuzvzQDig9BogUW5
fkzQQvL+4X/1W8lGUWKmJrqm7HLrYVkgBa/xNQ/XfqBAmyKo3DS7GLtdmfsp
o8PKsZ9Nw9PrhdVLszLQA+3i+O0M9l7mTMKCfmN0G07RsnFO3ocs3ZNSPCdT
suIlHXKgbudPrvhgU9lzg3l1PltCKjdn3NBjB7/zYLciMdi3EIVMXIT/zVRy
jj+TS4R+9itHJxpWFax3JQsyQdnKWEfLAd8/nxdN+ePQBKQO6W6VkK+LSjp9
n0re91z5Ya06mny5iJdqTBUrUVZkQCO3Is/AHpNbIKJJUBVdlEOoFp+RPO2W
5bOpZWSy7eVO2sj+flafAN58HQBZU2pQQsApPw347u2WB/Olx15OJceUNL5d
dkgJ1RK2KK4n+wxPCSNYCvBO5Uaj/xWavHenvgSa9krzAAVuRgkZCujScETj
8a/tZhy9dI1kAeqjKxDr4NUHlrWFOx27Cd29zc/hx+0osVPkqg29jNucdIus
zGG404VPzn1ha1l6l3urBu9zhDeQS3S0zUzX/gJRHJvtTUwtahfL+6bngsAb
3xVPjkcdB2XMEWu9nM2tTYJ03ntpu2v+KWiLzlxvQUbJEVTxeJ6vXtO1rw09
lc9uoNRe0ScET7cgCs+YnY1ErgRxkCQL/uvad1+ywm7/8hLhT7nr2u7i09Ng
uX9Yb4Cdl5as416ykvqj1c5TwfG6s6RcoMstkz9gwPjf225iyAJlLue87+0x
K0g2Sc+zXrg3GmSDHiYIo3LhDQwPA0yxWYWUOX2JL2wsAynT53QT/TWDr/ET
FcCJGmfbsmJOrTWIRXfdRfiDB9jIPpjK1RICXBqY9g3cPuvCerUcNrrjAaRD
BNJL12KHgbxkJtvKY8Zvs0LnSxAnvvqWTnVEte+prwT2uRdAJaTZVfHzWMKl
PiGSrSjokQV+suUklUHdoTFF8tfZ51xGtSkk1i2pgGHCD6R+Po3fzAR3RvV8
FsdqMB/bMrMgfhrFFUgoUz0g7/HAtTVKhWX3MsCwqNkUtfF4b5C/69izGpt8
GTNtVCL+SApJkhWLTBx9OzOWcDkeuhdWHp1MzcljGqqFLd685ZdidgsAhHzW
DiDqBkyqAOQXQVaztxzGvKGpemZPTZ7rJ025aPplOYxJnBFrss7DxBCprji4
wZPcrLiM4mCkRMkYwhvlcWbNG0tDqluYNXB7VqxXWII8vbNRrAbrzoFXPpQc
eBOo+JT3utF2DMQyxP0eb9OC0gsCvdxVp8P0hc/RDDOMxdmcFBm25cD+DKfd
4qKcU03kiY04yq5U+Ot4lzLeUmnX2FHOdgHtKTxbFpmT4wWT0boQtJQT/PYd
giZPF6ldX6usLxGOvuTrADWbB7sVurOJaKTLOn/D0+FETNTaoVTgnS/MhBVC
KC6ZYR0aouEe7sxTO+YpxwUvu7o/Jm4xRsfkUG86ZWfqc+Ryt6zocbFiGBgr
BbhDnljeE94offc1RfSsGRFrNkA+k+8Gr3nHCnC1MpnEsV82srRoOuNCDH5q
8MsbolzfI7Pyvb0zcbgVaoG0XsbUgokv15u+TqZqs5tRVM3pCf5pFxBL3nHY
pLnnjOjFmg2n3C682JSo5qzPkRhX859m+Q/qLDWnaRiJIjT4+bQ/tpliy8E3
zH6FhNbcL7E1Odx42pyjz9DV9c3G5Q31cHXwFmGzqUpRr8rDAqXdOgc6oc4l
6ZToW0dtwfMhEhT94813T3S1lCOxw6hV7YTvRiDRHEiAvrP+kUASY1NoFGdG
VE6Jxt3NRMcEkCSbe/iV8iVEGw/bCHTQb7jUyIPvJDOPspiJr3CBbw316OLb
bVZU+/x6sGMafcsGD2l7VBmNJRGjxMyvfeJs13+bWKxsgZkfLc0KrDAdqNuZ
kt0VN3En5aiiLMnAlCvBb9efD1U40tgisuPci9jq/Wrmef3EfwDhhuoT/EqI
UpcfbjDNgxNelOnuTPKiNpTWhyBJrDqEoFeIrpZ7Afefdj2KsOVz6xrg6Sja
7YksasgdVehldNzRVIObZKFqIRpieOGxu+fiNiHwdNWeGlrrJrTq2BmtzLhS
96WMksxOSFVs1enJjwEtnHJr2CJK5zefG6AmWaYlSo6w2eqnoxcbJL96WQ2c
s0ggGAVdsTDCnwCIO6u2AwTvwX+usY2H92DxXBbQDOz76RqSi44md9/ruVxP
EwFh5k7kQBUJx04wdqRLUhAkNz6hvsvnTn9NIF0/WnKJ6Js+REZdClgsiAkw
HIkbpYi8NxcWsRLsjhcoQycFAbIDA/F54e/N5d+PypstWa7NxM611hhkSS9a
mp/erVSbQVkNkhLbBGFMzL8pl/DxSvjBQqDB9CSul9rStLMkBD5J1l6zHsk3
X5CkbcNMCyoL+RQfI4em+Jjky4gfMcsrL1sCNyjj4QPRiSfODs7Vqb7Q1bL6
og9DnENVipbOvgx0RjGInPDOtN+wOvzjiuSzBSAYVc7/Br2xgRYXuP70SE38
puZ+cX9hKDEadY+QZgkN09oogZi0u6wOxhrvg87nDSC4fu45w3+DxIdS6HS+
MpjvEfStUbNPhyUoy10zhAzcuCrbLLijKuByouAs88cmiOSI/YxypsjOyTQX
Jc+OMzYpDNyX+APsgjt/SPMU/0LVNPuQ8Md/oUCPGG9GbFG8mOKd7u5aJwTL
9Sey1UbBjzM627wPtLcb0+cBuXcIs3KfbmMpvq5iKYzYCoRY8v/qRfxtlNZA
AgbyJctHtLrP2AmuAIBnET/mglRHnLahW/epBv9opCUtm9wEuZfJN5b/U39l
Mlo4sTis+uzYXZZszQ7SQd+Mg+aPOp2OvH56T6KY0X4RxLJRRSCtUmrrbqxF
mQxxlZ8x3SZ/w3T1LWkmQ7baBBREqbTGvD+bK+gQNd8/bEc0oTwXxtkiDYi1
7o1npXrXEZ9NWO4HNvrMpnuSDTsto0sC3a9TnZJCH8zaaw2mTek4PoFkQdhY
YNRIt4I1nVDym/a1x6ylqCGu/v0Yu4ygTzW8kANgkZXkRx99d8LeZONJuPhz
6nISV6+o53eRaZWAUwIP5olWakC+PRU13o51l7NQFpnCqgMkDTubAOPEbxEs
R9U5l9EUldMsOuaOF0k9A/uBukfSdOyuqitLwoJHvWI8yF8MOBhviAj0RQqy
8398fmTuXWNonFc8HVVmqd2zBS7OdkEZN805fDNQSXc47qmfIiBAgQxbqalj
v3RstOTzhREiQRqJYYBn4AXfaVAtFZtV2cHIVKI2ZO62Yfzzf58mzhEiggU+
FGxxB8vzCvkveoxctkDZjT2SUEQCFKJ8Mf0jUxXMPQsY7+GrBA5IsqpxQ8k5
gcyi+axhCyZ9recNB9glJdCKd2SKuWv5pnOrBn1PAbCSSTZr7x2SW/kqB9/r
phmiTMsThWq9s1wXdtXTB9P/R7W1+2CzfMOwDw5qXBV9nDFAwa71yAf+NeFR
fYlIbyRpWagWkiimvgohNHZNn1V0ADepsoNaGULkB4iLjJoS3e/DLAWK1Oad
aE4Z8AcYqpVodejFZ0gzJoqpCUbj4AVa2lngwTGLVX0fXlXaGfCc/o0CkgIp
oGUbQLiXArehmbekzG9UF5NR7h2YJMdt7Wy/ntkv6DC29Dfx51XA8x8eRt94
DZflRBBPiW8svaGG2mnRsmb4zu4oGQfeVrirnB55NpyI/WsNkjvOp371Yx59
zJKz+751cCZgqzhJUFQRn3jg0vYbAYilNZfAlE79gNoIT/do9cAi4EzMzMYE
SyTJucB7s+mALAD8TjumfHtupJbCHNs9lz5foUH6XPmCKEtBYaZX6q0baifp
lPfAThn5biPy0M8pTa4RYgeFoBf2qgOK1MJBUslPIweeguI9oQ24jbesKQjt
6Y9py1fYdn4UsVV3kWam4B4P/Z8xj5voqR1SB/747ot9NJsyrIQU6sN9xWxw
Q24YiSFxWr65Bv1tO46BtwUeJ2ga2IhGMDOpdc29Pm6wN6humev0MgCN5Fb1
ei5nWLxhCKAK1rjvAySWnUyAo+plkXI3+Hi5TXhUMlCFmdjm8kxyahiyB0Ur
Crnty36NuJpOrA4p5fjazWYidYSkxcXSs8mcKsT/79aogJRQkiPKfFVnz9iu
a4IQS6I1P+CjxxdQTkDYRFS9X1061tVbDFzOH5aRXRxgC1eAWISczj6rl38r
n3EIiYdfmri5yHlQWEvVGtPDLLl3XHSOTh4Ux3ixOvnEOCHNjMkJFJ1JPqxB
wnICZAcgtRMVt+JjkaDQnxPn2Yik4K4cwT/bevzoQga0E92yzB1r5nAil6Ew
B1AXrwnomavVQM3fm0ZaOnFqxbxtaQb4DrQbOgxTF9tMJ5ECjBNDhrbP3HOK
8Ya2T3gm/UFvGI86igYKrI7qID9D1zVWulWz/VsBW4TN5+/vnJqYInFfvZ9U
pZI2521de1D4BZ+B1qTgmdu4R1KIkcIkBV1Zd+pD0LvgRSBTstxdnf9Nblen
ous/d24VdF2uXVT4rGNSMOgMBcDGEJ34jlY6CtCqefybTXa/Dt0UxUi+U2xL
fkFT2zRnYwX8Ic4K2XzkctV66cyAAqIVoGC6JsA+uCkWKN3zIKgpE33uIwWG
dOIoXACrjoBuzx8wTZyTDYy5o3mvo9soA4KBqrtx+DYJOpVKm2C5h/gWimf4
je1WAbNrPB9lgjpPqKhnmbrMCveW3NP/zKqVF2gXQGjCooRpZnw62qs+hD8a
ZHl8TPvhswsjR1zT0hRrmDz/lYwTHXCuPCOAdecHo6ahT5UG4YD1NFOe8uBd
8LWLrBd0ZeCQ7EL426S23/G0ee47GV6XH+GLgepMM/ZwjjHUBZmWBoBizHQN
W2fVfpjRKnyWEWrNKf0XfT2j4JkTGcIi6sS3ixRgSnVwq3MP8453+sxlTblQ
FtztsW8t6w6fhFLICRaF+cG3Su2KhNYxcrT4Du+xdncfFrBvVClJkxM9zImB
haR34DqiXVob4DLD6kFXFDJ+jTKeDlcS9re+itVr+OtanXDxR7BvayjdV7Ka
XAaiy9HITrrsUd7NBR+HiRHwliJo5ufwNmoBqqy0oAh3tf1S0bw3DvdYZ/Oe
l0EN/XrCLRymB34cK7Soz9IU+AUJmfzd3zjr9h2Od+TY1o/6CqoyI8mFY+aB
9WkDhGcpbGc+V+ge2c6B0KSQ+1wdr/733bjOaLBy1R//i9VrOUEzyRUeoMWB
W3EKFVOl6zP8vqRkIqIZlfNZOoEHvJgdwwgR7IJ97rMmIKlv2ey6fJtN8Ewg
DiGLmeLEoSFwCg/WYRxSjFJExIN0pJI7V4iPlwKdkDQ3XHIPe8AhV55i+ArX
4++GS77TC/zW7LIpAfmbxa3xYwyeoSQobJ+KvEdIMG8QWdTbqG3K+qhFy7ON
vA5hN6fz3PJFGA0GxwRyEzoMBtNrtveLoopJW4sSMfu7fYjUhe7cd7BqtfBe
TxOMdoIVk5cGOvHYeTta8hVRCtASur0ViWVs4jGvdDNWvDAwoG8zsJZxCPpT
E1gZKQtn9RGcex6tEc3o9kjLsDCTAHeViO5razR3S4DGa3nbdtE9DEaJiPhj
3Prq3IyR3T5ME+Ge+WHM74LKDsE9ySlbItOcFalQzn8uCNbnVIOWUZ75rQH6
guXwnGXgj9KQvxp6ixb+i3HYGXI1Wc6nuDzwSul3Yyiuqdrst6ThndJgcOhR
dD90mns9JrnPwgPSPKrv570VSI7fMYivYrx/DCIl9sGAAX6gsCXwBOPMcDrH
BjJNYO4FSyyFrI7u7R5kKDz1++3S6ePwNE0wx1Ry3L21WoupoJaFslknZFI9
xBxpGjOnEUXIxW879f+Lpd9H38Vg7kWZ8zJVqGMYKSob36YQZxqd7dgYN1BS
umgdu+Xr37w/0iOXFvPZlh7XISTK2nU7EM4jwvYKYZFfPKD6JV/zvqWsP/XI
9Z2F3vNDHGMUlEYSGq7R1iAo5o25dG63VzCNzqXuhzX2Sge7kj2Ny4ok5iug
8qOAjW+EyrEnUjA7+J6wTpfsFBIujHkFhhqCxZ/RFvbhSEVTPQejWNUrApl9
Kjr4+zOQIehNAHllFK8QN4EYq2K/sR4wBSo2wFBJw65xsvFSRbbDrhpy5d9c
TrOBk5blbRgtm8Sb3CL4l7hbTcSkITDvV6/QxS9jBIP6FM2fW5A2RukDHr7c
nvp5MlGLcCEHZn3sh9gg4E8p55Vy1ciXGUf8+q3pY3pHqKskK2h1iqaeO/pz
pHthUs5aWkR8raHFwBHEZVDdFV0f1HbR5YwMIlssc7U1SBlTe9MT93Bsc8LP
v9fJirwr1DswFJ1XF0GFGdY4ASU9VUhM0wix/TKxnVdjS/5RISYsYNtiYWEm
Yy+jiuoPXk842P75wMEXxbG2DYlDVesOhnSjtC7CPH6ojaVXNSV00jbH0WV8
XtXb7K2/BJY5aZMdxinluEzGQVO8FyfxiSCHzEvdFOz6ogYSS0vlVbBvyjw0
tOLis00hT2SGCsYi2j4sXdNWjmxUPpPrpM+6Gcs+n9uwsul/Uc5h+D1yi2V2
tttR9qY4S7fnBm6yo3t2/lMgX+uWy14qmOiYthRcOYvHKIUAkV7KnYy8OeI3
0DFrRXrWI3YxDR8F/9ucA1IxDu2cv5phxZvhFDGNbYWGvrFglXNDn4jtZODC
nk3zsgoNoUNYjowobp2e4LWU1QQaIhYl6AObMcuLJrI7P0lEVU1o8eJbXq4e
3M+0m3UONj98B1oaB3mMCUaKMRhch0oq2lbY3Zvijeg6wPTkOipz7KNb2hss
z1MqEZnFxzzX0hHv+HQco/jw9JCdtC1rVFCnWHjxGgMy/sd7eXQDc3WAOcQj
FU02nEvJb2jAzahCzgGoJb5m1hHnCVUMyemHCR9YXLtpFLVQSYONPOBDvmVn
G+ICjcxYI7CjS/mlKcf+IbSOrbL1bL1LoLbk8JpSX6uCyQLVe+DQH5prW6W0
7z3bJgHdKZwvwDOJW9Eq1S0Qhb75aUkDROsUl4Wrzx9OxMGWAAxmyISjD2Hn
4beFdsCWl05yBIvqpi8UTLk3zQwk4F5W1Q5qeHMsgoTzLDMs1VLXxopMUQ1D
C0viE2GNZ+ICHxgjUr5d2vTMLo2lE3R7HrKtTF8HWcVPWQxcdUGrPpjuCuQ0
dw3KI+iwZOf1OcHYoYFp257hi38M2cPMO+i2OOlNuh2W+VXbEzaTAPK35BGm
heeQDg2Ie/KNeCpv1Wf4ESR/v3PVpLbW9q+hLSDiWDPWXt5iHZFmb07H8VQy
9DExmeJUlNe5aMAJnCudk6nifcvSF3/fvjunRHLVfuLQxdIlQqjmWL32fzJK
UIejghcVMoBZc6dKlOFnIVgWQrLfCrYChtSC0l9RBT63SbgC1bKJWAUSbrUR
j/A25LMx0xohpMMiSwE1+9Y9zPTEEUeNMMIqz/6HsTbmULIpS2sECcBg0+eU
4WQkRw+Y785uZ4yVTxUjxgi9yE+LZ6D+4UxKgiby3HrtZm2ow19GSChesoH/
XdtCqaWqVGR28VTrV07mzIPcYbax11T9iFS3ZwT4t4Q6nP4ujrlSFaSrz3YN
UPbUYf6OTfAkRe6y4hX4vhBD9NX3XJR+sSYP/hyQb1yb4nc/UizlSJDdvuea
NS1d3XAzaUOezfeB2FZVVQ3RWlUbOiWSmSdbMm9Olb9i5glVoDq0ekguUuPR
Ca6WXRtv32GirDWTcYCIXSmu/LPqLKDvhSXeZdoVPFcfStu/4Prmfz7D8ahF
pD4yt5pAUOB+3F0gmRZMZsri3lxCSWtKXdmv2J40KtnancV0M0P12Rz7YTiK
MUVlkoE3E2YJLPIO7mtJU5d5C+uN3uYhJYJ4eT1znvmybbcSSwGjNLenNjVa
hGOC/oa+xU5XDUfahJ8/VXRllyLwPKmPmRTpulWy/4uCRZyWJJocKVx0ffB6
fprdBRClI2jH0+hbewPR9XGaaAHuOSSrLH1PtpeNA9EKO1+W55rc7rzahs1h
LgZEz6g9eUZns3NG7pxR09WE58p8TjrYA6Iolxbai1EY9hp2Y58JQ1p3w7IV
tBv0ll1Dsyc8x3dL9k4ixL8Sfxgm6h0Nvnc18grucnieBEpjSP1vytT+KiHH
3ikQQPAgau0s9v9845Lper8SRUVOd3YivCACcnTIa2wY3zdALVGDdEOWpM+/
GzfhgxALdppkKqlIcStvfA0IH22NeVEwVVGRa5X/TEdOc2WNC0v21Zj9Icex
Cj8tCa0tAkxiLk2QbYaks4AO9aQy/Dso9lKPdkiOxu1+oAbaZk9dB2LBpeQ+
FOOwfUXzLhidOD7lRh+x+L8C/QF/m5ufQFI+caGfTk1APsWAAXHIn73DVkox
7SYFKXlTSXzTDHwZHNKNtd6c4EfVkp6bJL86PW/9F8zPcrA8SwILBc1+eQFL
1UYZVh2uQDARnmnDC/QyTN7ZhrBPByjXwEo3M1eyY87pW0gin40NH6M9S4La
o/SS6ms4J0YCE9q4GdKEkLam+Bk+nrQ1+rQfBuCJUH4Q8r8gPreN2ZV8VTVG
NGT246k/J2ONrsprjtRvwgtqacnUJKN933vrm4V8K17CWJyzEm7ed/8tt8On
GLFZsMReXpRif/31k14gjDUWS2O6ODXB399V3WTSTKrD+lvFBxw+0aYuN6NT
KUwI8DkKXw6dEeQm1WztHa6IpQM42ijo6qqvz+EFNvQSMtajsVDKyx1EIlgp
6QO8tgV1JNUQtW7lN5nq4wW5SsF+2EwFAY8JvsB/sEQLBX+Q1x7qa7gbxcDY
KmxPXHUIoCYgZZ1aca0DOtBgqvChr2u0YGlzuF4nO/umYVuGMlmsTTl23tkN
0Nc3QSIjo4Oa3j/P32xg0WMtdIBWuKW5nEepU5UcexHi9C9NfJr3QGWnMCD0
alqSxQ7xBoa6c2UsmDXNGrHFfOMjRxZjtLz2CgGidfhNI9ovWE0vYo9pvv2w
wsVhOpy8CWPOft+R+RkeiLP//RLKV8/dLv2ILw8rgbs+R8RLDjc2i4dSeG4J
JzCo/PH6JooqMT/LJfU+58V0qFftxT4ArNS9Ko6+5OOWrdOV6NJTBn+Ng+Vj
LJt6tSdeQuR0lIHrE+DzF6GN7ExgYhs9UNB9LrKkjjNieRqxCXzLXBN4jDSH
O/Rdc+4zA3LGoifvgVUJpSp8MayjPSkbe/8drZjgzkrY7P5w5e8eq/HCiOVL
y5q4n1gFGkseqh7Oy6aFSWJGCUAcsgDUJm7nCVmseU2Sg9Nzwc7soUBEoTCE
yD4tQT/vJc+NDFJqbkSLvccr3+Yme8z6Rr4l5htASVFRNjUsEF1uaNHAc+Oe
VB8d+STKHmY9WStjuPL0RYU5EpcFFR1KBoMKnp5/e3++MtnN90098Kwla64q
EB6NOSXH14SXsyiYvOGDl2t8WAEz92VW/1QQdxw6R4X3WyN2wizlKnZJbS3g
nILsYnrKknlCe7gaAcQqLdhre9lZoyEoGutwsrt/ESmL3U1Xdk7tzzZMYcMO
43O8+6zyAjLZpjjXRpZB1Xqm7AW9H+nVD6z6FxdGHqPXWh6POCVKqR/1H9MH
okAnW4/DHMa9J897fS60VLJ9zhtCirC4nZ2VqY/m2SsRCNmekBOfxHW/extp
PntrXOr+zin8CojIYRFFjj5vAtbcoxvThvnHObDY7MRT3FeFrs6F8O3AwgOM
PIpY2ZM6PyuJgm1LApEdEeVGgBRai8naHRgk3GIOgCxT0DOPMwrpAKeX1wOx
wtuiTnzkb7PFRtzLjx5V7haoG1B1eHp1Gm3hoebyRK25MmSUNzYB4sQFxlwL
fpL0Cqr/E/jIW951jk+RxH+v96v8LQywGw9NmaqACluFMjLMMYZHExgNOcRu
n6woXBIlWPWWe2g80LHb0053RSqDDJ+QhURuyDaz08X8vDX/c4oyKfaNEQwF
F5xmqiu9kOkIvNt6JsLOLGxdSABIjjon8CrOkvovTQ614StMEmtWeYqqJ8Yy
0NE6aA0guL6RsskgsBg14nBj2g7r/Q6Ue9q0G/+kZOq5SoMrL5eQnHT6b+hk
96DZGHzaA2n9re/2grklbLOSD46qBQc6w9pieV/pPpZPrnFPDUiNNwB3AGmV
iEwL1P+dkRLks6XQZecR4y1wZ0ccK+bg1wpk7FusBS49jf5NZRzAXafJFqsV
BRpoOpIryqXg8yw8CG9d35nY7db34rFf7MpZ6vuGDDa0TbTfwnwfXShYgeIb
M71UAnbusDmEgd78O+dA5GGfe59l58ERVfYN3ZCuzsswutT93BrMwMMok2RK
qbl9WZUvUub0vwmTJJNWI3rXH3V8lyxW7G7Imw8bYk85zjSPPu/NlYubYmMW
Kxd9V9vRczJ807SeEPrUWRKD16J8ZiqSugbRr0liDJvBW+kWQFqGl+pCZECN
tQIQkEn/o3Sj95spRAImUoyYWSKcJjGyLVOn8mjGledIOE2tdCW+Vs+FTKEy
6IoLErZOphT0+h502zh8+TG/9mofFfDlRXIzZ+Q0hTBXK3nI/qkiYI/K3Qli
5fbpZ2zm3JAK8PUqPGMSnLV07isFqUdAvbVR4MvrHJZ3zbOOzsC9SObKAIPH
dZuNng9rinMzDniTfDTEgL2nGZSaTynJk+FJLAQO/BOaYto13MYhxualYEmJ
eP7CViMtaire0OyUjntWc9G/x2NhbFSaSlAl7tGWuZRKUA+IDo0mvU+xKgey
5KWgPCQV3DsG1MaC7PYTFXrpmED5v/8F+nTjoD5rFhjpdtYR82ecZ1VZpojQ
KEUdFebxOY1f4teIMaxyAGYzUAI1iHXppjViwSFKjkz75yVmcwzGNlAd+9tM
eFWfjrIZYCCvFk3LH73thfKZSSrbI8o2zNXCvWixI9yvJhqFoUorXaq3FRIj
uBu/AySCJS1HNv+5sk/+tOr9HVJNi3YFwLeRXaFw9D+hDqCBdXXgwQ0XsCgj
62o2TNEpiX+iaL0DXB8pUBnhxM4IzJnZHIoVk7wRo8JLtpyzNm67qrnYmTsg
JOPjJPThTV08Z6cHs/A320uY07eUCSxWsyy+1Mh8egUQo3iIEMpLl9yoy0kt
+eHBFGw+E/3EKxZrsJ9+mt5Ull/TZbgMC1M/wNoBTGOfhZWDoe3h6n+Fsb70
GAuuFOkoz6SMJW6r5x6e6Ce+1PweDe9v9MekBKDJ2M5du6Ds7irdqf3G0bpr
qEpKhUAJOYvaq2VgFZ32/8rhu1bl8f+51Dj2qpfZDZjNBtIFR/nw0W08sdZo
8Xr4mZ6OYky3tvg0iqS2I9ySX3MFKpl+BQQ+TPH/SFCxOSSleWKFeE7lBBa7
dX8xbIAE5UGrTZtaHV+Tdynia10VaEjZTZhxbYJbfQvWXmHwbqOZb6AYfWxR
ZDqQDqIEEkVrY6TslwhsvD+kCLICyFHa/fAI7SD50rXxJpB6Jw8Vvgwhn9wS
FVEJhCYLBG4i3QmCem2UvMxpb6S/SoKufEnuyq8wRpit20Q6OC5akGVMRSB2
NUu10M9IBcqvGR5bzL4ZPvXYS5HQybDAeYyUxi1s+FZde91kYDrQmJ2ueaiZ
eleafcwjSeexhdIEWbLw/n9QQgEzJRd2qizAJm1wY8SZ7lG2AuOJLT1Kb04r
o/Mt3R4de7Jq+wPYccWaKJYvvfnzLdylpOEinyPmFTPGyqAgICFgk0qfe0at
XUEeeqgyo55BtU1SvxjUgyzNw0j9RHFjhILQqBJkgLBZpl4KzUffkO9pUJ7x
dKlahyHJaSQiBzMfCd42W5bCpbVsX4IxRSHUZ+islYxw0mgWqWmmnpOGxZxy
QIFhQg0bbvSfK9se4PERSCHEw9SlM4CAYJplAuuEXz4efu05wJ5ljmm7aPHs
bnlE7kpm0hlGsGmfkT3Qvg80vl7ki+Z0G7NXuCYL4V7zl6bWDYoi03SuH0MY
1X5nVMnB4QsjkZA0zT3TLXgvHRkZr9LuYpXpN+OwjdwmcDrWgforTugS3O9a
UxWflrdjHTR/x9uJdRJT13HgO8DBcIyFrFewQVvV6ZDJDJY/bygSszxAWWW6
sKAABfRpfg8pjRs2fS2Qv2PvXVfV6axo1T5XpTq8RTRXgyC/uSHTW9rFwoRw
hKvUiU1YL1gGS/LO4bWg2p8SrtVYn4rCTmuyeyS8Bfry38M/eTl6BdO6zNGq
BwJ/X+axKUvkAQkH6EvuWoyAc3Ge9MJg+CUsYC7qKYEqw8UD8YE2zFyfFHiH
D031F5RE1aJZ8OsHic3mpgR0FoXDAafVVXjtIDaPE+tvm/VE3mbgiSSKl8xK
a5lP4lH47hFfKE3y4DivkM4iA0Y9RO7hkXln+alomhVt06wgOttHAWioOUJS
XL4RU1gbRg/5fpiWOojfbJxp3fYU7vGUlUhAJmujgxlGU5l7LGrmHiWKzasx
ble/SyiVHaxv4fOtMITQYga4+Ph87KFjofjfTHYgU3q5fimP9wTK2vbCHlq5
7lRN4ze4Z8NfLVnW8TiLJ3r4htB7gcgikejcbIj8XlUPQyMNT7+eQgHCXSZ0
LDempH/pK9NRUaIGLSXsByC4vOU0MCUfiIxcvY8cEEt8wIxOCcxpdExh6/5c
VEUCOSrqiJtpgYo22sSBdhUDMyHnq9qdn/MRoLvCDmDpI7XGVVywge3lMfWt
uv8HQ/X+4S+EN/vnc1vHKj5sm2gcnJGTrR06fSDIgWTw7BE3oS1/qOR9rZxc
LglYVhmFh7UNpIqrs+IT5hxq85LPIbT+UyKOSBjVPZb2G6v947hpmdYiyizs
2MNW4PTasV9/Yneknr8n22X81neaFNU7hJtL4tGXogfR5rzWLDK2jP1HxPSv
eDG0FeK32AGs2BVsS4JAkUy03/kIKosmNGUcgoVboIU+Um4apKqF17UezE+z
2fcTZq7h5GAKVrYV26rkVsTILjtJnvJ7/i3/XaQdlzDg/CgKL3CwVZoHoteW
nZqYsJFYZnePncD2/R76257AGyYa/k7GkQkqQK5pVhoh6H1py6eAz+X92WHS
wIicAjw9NNB6QeykPMHa2Uex1/oDInfKGKnPJaPD2DFiRX9p/K+0ORXv0LYJ
DKLHx/NZ4YXdVNFPh61dLR8SPWHS+rt4cp2dM9pa/3vqgBBc9ehdD/Lyk3bm
ZMBo1dwVkEROvl3Uk8ahntnwTP4y93v4rb1zcP1BKgPJO2nHl4v9OynXYc2t
8kYsH25LNSppOdcCg8DpUbJGg57QfxSHOhPaho+k9YDb1GmjmfngAu5X78Ay
SvUNIsMKF0ScG2VCN7j8pmL8cY6yKIDggxrjueq/W9mlc63kRQsIW3lNzI6B
95n8po20FXe+pyYZO3u4bgzyiXnDOChFKVVcdvEpv+Q3ZsAAPhFwCv1oxSIl
pvAHROSjtWE7CikPAE44bU8gQgJucdRjasxVs4pHixwUxh7gly4RkP0ZdhPV
8VsDQv3DAQ/Em5Dkh3Iw6icIz6TqLREDWSKQtuiL3cD8hdHhBran3ipJvo2z
JZUDu2FWSgyxJ2kFOXs1/Ov/v0UCdyVBBqteEUynyj2Z2H+5LvwNHSKlnq3K
oVDmpWTqYrk7oQxyz9uGP+FDz1DnFe2ErYP3O/3vXy9ndRpA9XVM+BeSxPzS
MHk1Y6WD3ySh8x+jVMXEJVz0oxo3PyQaXw3X0zyt+CQDPeZVxQxmV8seqHgQ
wax6yp9WTBJ3U+WxGx+73gcCNW1DYtRJwKcCRvw5DHT79E8/x96GmiI4sbSH
y/tesRKSFXOAAGGmnfGY8fSvRLVZueC5wjNgwJ9L4mbL0WpA4Jk25A23baot
H/NNNfua9Y6GNTBVV9kK110elyxy4ng+bDS8M64OxILsh584AllKsNgQ3Aqj
KiXdyZLZ/UeIot+HyEGA4fcmxcVkkUpS40JkBVnpS5bKbVgF1q307DZEVCNi
lbiJ4YwxmfLzcmrl3cOGxziCj5SRkuTUENXo8ONY/QeHRAOYPu3qtmbhQF+f
cW0hiDD9I7qGAJNrbEO1WXis0xgeyIF4lbA5W0HDvilSZ/L5Po07W1jLJXKi
RvQW0rTnbVBgWlXm+EZqHf//D7bl1llgQpu3rvg8SIH9vS+/diyUUQR9x/o5
h2t5PRRspHegvx80PjHqwXglSPJChUZCmziRpKmcBLNui3M0ukKzdewQ7rdK
6jvc8vnebjiTwfm1BBZJrHlTxK63fBHiW+iIp+WRf757Qxp8VjU+DrUE9JD+
A/3nLpC0HTAmWs4RvSjtYgU6wzNUVI7Z4tCbu6dJGsZMF9aHspZ4ToYgIaxs
dwRw9vDNV/g8rYdtMdtqQERBYc+qXm2cpaE26lUjV/dd18G5hN4XFnZtAjqe
iH2pyX15sqq+oUBvuD3exuSYZb1wVQZmGThGS3g9y3l3xuilQCGpedpGqN1P
eF84MTu4d3hIt5Qv86z6517F/uf9cF67BzoytJkYXWSiwJVFWDrmZY7SKE9x
+JJMnzX31kE5WkhwLl3uJQuQRKqWBsIV4ZCgNAezSelkiDgwsV6yV0Yfbmz2
QdgiWwLPtiOycuyPm/S4RNCPAuTnkvYedqL1KQaNS6eFl4dM+UtswhCvwap7
yCgEgvrx5T9miwQrgJC/6QtZLBRZ3H/xwBZrVsc+0eWBOVGg6o65zd5TYFIy
PuyrsuTroyQlhHrULPkBnHREUHEt+PPrs7s2teVFFSehSgTGLeh6UPnSZB+c
BtMxE6Ls5A4mCSxbU7bSCAOYeyxGmYUuigwqe2qpC+m+vGXrNNkZ0PF+Ov0G
1qQM2crwQCLWINM2l2Z0apFne8j+8q0ieCUt4qXgvnevyEnIr81cmXfkhGkx
l2IlwAzu0JJRdd7vDBF2qoEtq9bTp29NEnz/8MuOQHp7T4RZpF3MQAIPIAwy
Xj7+b4jGiDtHgU+ohLHv353hxlJga7ozj1KjZZ8uTujkxso/jBmbpp1hqbZK
+Ttu/d2BCmgsqZPnVlfddj7nhFCJidnWo4z01DeUd/dzAHnQfKsI2XeiWc/Y
479rmJsSF/RF70DNf6HFRX8KFcCom/zkwWw8KUA9MVKvSemYznJVrataybVl
AKZhJgCj8VSgu+Dcb5etnj8HXD+zNKAPnqDO8glCnygSVrHaiCznrUidjuYw
IFB25JnJAqDdy94fsCzIFVcgf1pyRZOYDHHU/6ucVtr8wjfwMJsyREpTxwBq
CscLqpgLnf78zjzHd00rLIiTW+7N7PmiS17ndUZo/3rHKlgG32Rl9UTaBoji
GNY+uzwQ78+U0OiRVa2awaTcdV9N+/D1SBUBCbRDABH227+MslhV7nq8lHxc
d2lzMI12C3LrjMYdHD/tdWtcCbMNLMtzPOeIV8xdDEEnLrX0OeUabD7keKPu
REWbz1b7UrrS+9O0ktVRPb/5xQsSCGArwl2WSC+zwQ6sobNhZbB4LdS75z3d
ntCNqPF3DXILqRg4DnAXYPLu+lOb1nHVL/wKCBj7qeoGNN6bMNW8/WX5YTwx
JChK6VfvI+osVMKZgdZmWSRCJbYPgAStc3sl8ErAavuR4c/d3qdTZvo2s2ft
XPoeNVVF4pKA5zeAhc486E6KlEk6dowpyd99lH4PPfDWmfHLbbVR8RaW2HlM
GYmdRoKTJIohsaP0i4SwPzpNtZX5qf0rBBcXt52DCmiSefjbpWNbhModg4Ul
ryaGvkQdeslZYFQ2WUAn6FR52g7RnGtUqqV2JwzN0KCe4YzAdTo5miJBSso7
30fwG7BAHD27vd90wQKPwilGK0mdZbwon4OfPgZl3c7DcVlra7hP+VSxRjCY
/Z9k6ZtbWv0UtHj2GG/koLAm5EhHl/PEsRr2w930fPOYvndKYv/QoT3xcWO+
HagCj6qY2Nc5akK+y+QRuhXRMJ1PMCyocSBsKiZPC3kyhgZ9iAPrItIjYC20
lQSrsqDj85MkhC24HbK6KcEScsOA+gGqY6wCWmEX8bq9f6Lym+ovq1LKbEMb
nrFnIcqplDHzgK5cTwQEuEOaFVrXHo3twg1awDVbmuU04/WBRgc6pImdsHK/
atu2v3lWH0goWpJyikU6OS3Tna29btlp2hCkoM5tlxPF1/ytanOv6AEkhfVB
GnRl3jyb4ppE+48bNOB7YOyT4GswSNvf7AIOlC3pTkD2NsfYIrEd54wBu2ZF
Jg/g1OUQ8EHCnwHTabBEHVelqiA1t2TdvhaNkjGFua0oDh7IkVrsNl1wj+W0
KZePrvpphJCP8FZZ3nFfawGpEYochrMWknrLcBg18Gz3bdN94udqTJV1NWof
pwhcvj0HLVBj6m2mBmhQXceL5j2FU+7G490O5b5j7eN2UIpl4WizkDRrQS7x
DYEXEFDZz22qObnc06a/FRCOo91fuYatGd2Cpjr0CKhUmE5Y7kpLNPaTv1sk
Z1aWSKdZVcz2N8JV4ZyEeTfBPOGu7odx7mFKAQV3qzgrsLvvzmxUd3FVElbi
q6qujIHIAiuycK4B7M+mwWqqUgG0iV6V/vKgwEwtCBCqI0JU5obr5sZIs0Bs
qwEYbf0b2RZVIqTQRU5Qk+zNMF9dQs30wFp0pitohYE65ExSKJwlD0Vp4oXo
/FPVREdDOGdHLm0vtlO1a7UL0p/AYoLsN4anTf/BFMM5EFZlMSWtCp2ZdT0G
xuRD1aqr9ESpURNb/nOADw/5OnAmH3OFozKkUlzReUsVSuhUdfr6uKyy4xQm
YSi7VY5cCgDvgBpBSNHugMutSGhgT7ehGx7SlSLCeazYq8DzomVOhnEJQSE/
x9BmH9GR8evuJpzLc6+CmbWj1qER9dL7qD5ehug2sDzXQhiRiPpqEB87vgSy
3fX9GtAKkrWff8C98Zb2fG0x1MdTAWSg7AYzMNGj5QyMZ1NeYnl5kjflrRZ1
MJb4AlKs2iF/PDRGKW9ErUrH8R25KRsaAxF4ofRpNRjbtwGUGwXNmM/kTjjr
DTgIKHHwOvaXg4eQwojgbwTamBiCIugZcL0CZHxScR14NxPjx35Io06HjKR0
R5rCKvhRE8urjFPad1vf4VXHxcymJ1xVktREliafYPgq4vifuZEW6XtNEp0/
hMb76TzV89uj23D4KTSrH1USv5fDWsTtNhWwmCjvS0COFxx7jAIjaaeR/t6h
onfexKYryeoUrVwsFvI9LEY7mrcbApc0yBMQCrtXBD79UDPpz2yFGxco5G55
nTb04Kbk44s6V0xtZaHLBEUy13hVX52D0Y1ULleyu9GWVuQGBKRszZg/m6Kk
MyLSCeQSMFPGiY09Xvcf0v5Kaj2oTJihFcX0W6+b7dV4Al7ZYeLYv+G+QLvM
ou8qjtt070OX9pL3NiAZ3qa7axrSEFDJ4x6iJhOke2U0EpnuGm00q48fVEvJ
aO3bmpVjjRYhcbdK0gekVJgbNwBxw2nnTq7Vl2WNU49j5ajvRui6RNh8SATr
RY4mMh218V+L9UIwzvzYKCefQf58Rd7B10pJfn8hc/F9X5EP7u39LZwtm4Zu
ZzhVsEHpMz9AbMG7YWyYg8MhnDRmsu1LHr26BTkIx5VKmoUodCTUHlIuAj24
zm7GpA2wloONtGOtaJXMBAkmj4/+6hrGL0aXa2DXMKJv/9rEfRItpyCZ9TJ9
oTUzmCDebWo5CsN0Q0JmFrp3rUP0gLEJWSiI8fl3dDeO9LiCq7oP+dqOVAAv
PIlfA1HYh1H6g+jKK9lEqHVLW44KB++6S2ggjLE0RgXUR1eqyS7ScGM+KR11
kc3oBMP7FlL63NAqoWEHQqIkQfahokCzRGzDntG7pPV4THyj8lVHIFnGCSdQ
vSdAP0Vs4h4iwboi4ahthux9VuA9dZM6z3TR4osi13qSBz0iDn4JRymNGBRf
9DKpwoPvPYfqMV0utFg18T1WBnGVYZ+yZLJXFuTCqDzQRYWpz1WDjQjKUmel
ux/+tHjyXGk1MgQn7qHAw7leiXKT8YCg/CoNB2WRbpCCp3OEA2/Z3IA+RLMs
xRdGWBfZ/WKRZVNxtLlNMWxlijA7qg7vEZ/2JiwH3o6jw1hiJ5zsYUg3UIRo
7SbwoeneUEvFM8xYR38dwdDNLVbTV4KaDnbZu5rEmN7i43RTuM04z3XeRgA0
Nima/sOrteuW5HZVdgvH2iRwsNMStJsO/1kYQT3lOpTIQcO6t1XY9QfGpfVP
i+ManhCMH4DC+jHjFkCKIszDmRdnZuYUGX9evZH2tx52/o9hjLOKlPiqZeEk
oHQvFvLDkIlQchatmwoGtNz0JhhXjmdKx98KixdeaHGIwvbnVhNupvM3nZGa
XGv3rE2fQ4/ewluOHrHpNPv3uWJ9BGSUDWeaWlo8TvOCQbVD+by/6Gda8RvN
FhuBFIDHdVWGBoLe0fNfCv0jGQnVlKgVf/CJLrnGmE+pjeCqVhYniO37Xq1V
tSUWW2DbfSuykyUvryjWransl4YRB0jI9ERcf3+lNrf+GQNcp7kH9H/SfnAP
t8Pm+xQ160UQCYMI/w1VakcSwX5+gfWyYpnrIHQBcywurEqAb7URc2mKc/PJ
gbuZ6F8nMKfS0gtFNd/9VBHHlShAxVPAd7AX28JDwRO8Af74/S5USOm+UIfj
I3bdlQRmx35IgHXn8BNizKZkT7TK9EO9ig7T+qxCC2lmtyb9dwbdqI1XkOYZ
BKTX9k67AxDD69ckt/OUmzCsNIfT4iOK6dKZeBpZAR7Ymgs3MmxNERw6McxZ
/M+w/xKYDdjB8plCymcb6HBy7mGwWdC1L4XC9NI/IjVLy/HGEqj15gVihSbW
SNOaKvbH8s15BXtqxEteodqa1bPQdGLxg3DgAkHhq+E3IEQjtfKW1fBMmCQU
QxNY+pfxwex1RB/xj1O+0bgnYTKcBEP+WxU6GNVevYkDq0e16tolA3NvN96w
AKbIVTMZcW9J4bQjbzBf85T0DJlEAafquB3esG8Swex0t7UfuBBnCVXRvLmR
izr+B0m64+2zjfsyIGJwedDTqJWyH67H9m2XFFJ3tYnk1k0QW3qVR9eenLBi
sIB2ENBYnyn9n+RiBQ92UiGOhSVqjaPTUDapOA0EjfA/0sokGqQcv50VraSC
B+dNJBR3iVZJlTPdDK+KEKcB9krHh15XZK37VPIzmDSMxhsHVMNXFQ90fV7+
W8MAhtXbjF4F+KB+RcNXhAQK/jIitm7IKSRe7N9tH+h9t2QL+1GSb6U3UX6+
rHogg3ElHQK/5NCtChss/8adK/qe9ovhib2l8law4rmNFEi9ActLWg6aUn38
heXFWtGDR9rOlXlf7HGGkfmNErAZTi2WmYoOM/xj9Bq9Hhzr6CQWkaRxe4XC
iMD7MXgbqziDM+jOmMJm3LC6ygcfjRdSx/Tj5kMfF9Flz2XBKpiKt7UKTKPj
ufXPVaZZZJssm/qSEAgw6iXpcvxvvaeDmAFAtavy7cb/5AkEBT++dKGw48pj
D3NrLuIaBU4hN6U16pKkmmrR49K5jXxhxN834HkDJYaJMdgur5pfOSijASvH
dapbeMxw00vhL44Mxah8nr/2BjQspgasy7Zkn1LUdK47rvzDlY62c8Uyu9w3
WzLVSyFqcfDyaJwJ4/Vf5sNBkn5Ti3EQUBTWG6WA0fsGVKo3n0tfEa2I1q8r
NvqRbX6YKygYR9QzZwq/HTA8WrifNO0rdoV6/P8p+Obo5hOCINO3ueLsos7A
yO6tjIRf7zmfwOo94HTlhcOdFCyimrldU1cnbvVqe/xLGSoHrfZuEE4Jb8sT
DrRcl9zX0soamGct1VIYewnXXdk3CZs7hcu2p9UXyn9pfbN2JHXbCsm507L+
4vS+kitm9oOJdRM4swZDOauSuCSXDfb1HkzX5OLcYIcIjrU3Y2T3K4ocXyKM
CXpx37HyRGO7Zz6ZIfUmgTHSeQmNN/TIh/OvehZq+TN6CUByRL/AoyWjy+vr
PTZuVGTFA8iVSofrM00Jr9ueOGHsrkkSJXubr4lzIENqJL4s5qRrgI8hs2oE
VRBS1tewr3orf1KPxMju6+lt4qLBOQPhvtBHFtHwgnksHWDbbe4LG3Z0OUeY
RE7IbF90SrO9Q4Of96EECY0/4Ynrfp5cPyT8/kLDGy7drda2o/nGAs7K0GYU
gxFl6MAFWFZd7DReCd8rk+llnUxBb+di6AOVHFpHDkigGIkSbktGtyWhEn20
o3osHR2+Y7yokpMbYviUUM1Lnx6/iQIvjw+jGwGIZPfpHzn6RBzf2FBBWsyQ
/zL+81+E/ykpBdoFo/IXJ3fkr7KqChEVJi466vt5zM8zKS+Dqe0jSNkBrgXQ
Zzy4nWYmypsOKrJKp3E3is4SlmDGl9OCtzY9aIV20VL1lfUPyqK4pivscvM8
1NFDjVpXBFuMScNWtOicFXzI+wG9Weq3pW+xBkm46oyMdjb4LYt+zrrgqNbg
uCBVdokS5pIatNfx/Ny2kd8YPecdVEwMtJYcLBYCfufaqALqQHmCkT6arjhr
hWI/uNtGzsQlOfYBvChNS9leqH7iQzSqggvEDha7r7HBkeiTjPgeIh+rkJzv
xWbWV7yj6XwM8E7kEJHvqMtzMFIuu6iIxYoDorWti0sBtJub3zLIY4E7MwkI
HfbCDX53fkyck4JaA6487b+xbnwhtR633OkP3hbFBVY37tDxtQpXn3+AzkTJ
XzcZvquYrDYQMzswPWB7RkRquxiUjTXhfpn3sgIoBgtyeWuTKVQ2ly5U0RV2
Y7VRO6XTiaaeF4sSD8coJjmI5l+6sA8eiN2wVNEjiCWrOalVrSk9fq7+1HDw
rId56GFBXvwbGwlWP7JBNMUGU1iKoXFhoN1Dmj81JNjOBrUtAJS4n4VfVL07
8FWH19uEW/f19JtVWn2Phew5rb4yuhgkPvIjF2h0yFVyySwzFk09L8ukm2Fw
ZklSNTYdrhYd7qkjSKnAw4GhHnrMToxi4TAezC/gfvVGg4D3kCguxoBTVI0X
z73xeWLd92WdbV/aGglUtbvJZSetaQeKOF0Vp08uaG4YzpNwHEDCvOnADVo4
05vcAVO+m/nW6zK1cylhikMSgRQfe6mgv9s42qhOw9cEZnZvRpBNV42X21zP
hdqt/M93qGNb+EMjDi115jBKkqHqzDxyw7MRlQeskbfZIKPGmZ+OZp2I9RuO
bK58u9+RerLvCyy1dio+reUURuHOEPnH5e1q43+9ZVmfT0vsoDVzYmlTj0/1
z+JapMg63VH5zsOqR2iOfkVescpWSGAUS0A89a3hY4VG3iv7RZrzREjbztcV
mF94Uf6jxQQ3o3/il1bJsJQ4S7WE0Ct4qzT2VxyXWHotiV2txY/tqMyI94J0
lIGPxakVL3QBSr8zV5+57fbbhteEJviZka3F2+lVv3d+ccfLhjCoSfDH3cMr
MpFTHdnHTJCgW5eQiQq68gzB7wmPvkM74pLucCjZFYO9t92P7uWg1xj8tNhx
hMEPs7vpjymHpnwiDjUP8zy/utLKdKY1cxt2YZPlvA6MEiMvc/kowQ0tAtiE
5WgvV4T1vxzBD1SoflYGC2fAx/7QnEORduOHafPJlQ3gewpFSbhnkJ9rNIj9
RwlpMTwZvt9fSn+OrCsz3aENBpGokDjFpNLZ7Ivq6mo2SYqk6A5u/bJBjX0t
VTKKxmUzBiFldYQY/WIA7DM6Wbr52i0S9evcCvfEEQ2MakrG0JHUlZYJy1AF
Gdt+e/ta9ljt1IA8VmbpYemz4SaPwUEHh0rgWf++P8HTyAZ0KDGHvmym5K86
oa5P1lDtCDkSRQfLo90g2tWVwcGy+o9pXx+B6Ispf1J3ip/9t1FZGIihAjvj
U1mYhCUteKPzugTtAIBM08AM+EHDXTf+XX53HMQeTboygY6stumckGuNL2PU
FiAUw8CNcq/LfdRJERTmMcNqGys0S2lMHNqoyU/adpGxeQhMbXvEfWnAa+kF
faQIygNj56Bx0X22MWbICZ2+w+V/sXZ8UOPHOuag2xxo0UoeSR9dAocSTyro
7YgO+5cVpoIWlx8wNKRlj364nivXgXEK4nMqrxR0pVnkdWc1DW7GoxD0u/IB
C+sai7VXWKsYM5hYoiyso78tZ+LKPgd4rz+aN0llNwmbRP4FIMKA3zEucCUa
KQkFIGdL9KJ0WKBhxMShlyHBEFDbAs7PCW/gU3eOdB6l32844TaW94GRHNBx
a2Y+6pMvkfOJUuhH/JHU5g1PNX/j6tUU3277ouOChqL2fq8jB0TF1Ua18OcJ
rk0mjEnLVj1zy2Kp0tn4RrjfLRngZUmDiqPQOxYALoTK8g6jtyi96OyQz4V4
8tKZ+4eW/0QkqtTchvL1Rh2KDUFcLHh9NAL7Znt4DoXnQwBPD5docrOj+xlJ
bE8ySFum41cJAp1d1aLKvMwZ9WWpR1Ei9+Rz1AKc99UjJC/6GOWK3J1izXKo
eszGbEtxfB+d0YLPxr3AFOrtderyoRAJzRRde1r9nL9I+Z8/85tRdg/mBpLr
LbsemjoztZ1Wdkh1HFyR+N5q+c+Z/oIHe4El1qSoaUuCk2pYSYpsZ9HvNjoK
pViy12HXNgC9KpbEMPwJ1eOdAtajvosKA8Cwk2JF18NCRDHODDv6iHX5bRNs
WgHCZymfUGOfy4aPtG9RNLc/Qr69a6Ogc9vDzAYzRJDOLDovGo3V+tHCigPe
WP80EzY4ObbIh7K/kYYfIHcKd9P9ktIURtll7x3VknPb9Wg0IWf5VZ0coD2I
iAlD4YazFkyIy0yfWwXhH7ZtjN+K+Egj2WBzPliGK6OSbIoHezOR333yGns2
a7zC1DN2SiiU9gs7JgjReAv6nPoqKmKcsu+mzgKD4FoZIh2vNJTqC2edJjs3
c0tA97urfDP1tCQNi5UmuPs2ZRd7GSNQxu/F5dwGo3td1AgrJWCqae99HcHv
2kbnUo09ZjMgNio3ehknQLZEE5FslbeqvAK7sk9WxyaHvAudlRIul+xS8Mep
ChMlWign0Ko177yKQ4jvA9+xqZBY6urhsA4b6QcTiWKMEY9PeWZ4gkHEWbEL
IEekb8GJnxJTUljmjlYb/haI0SCYpYdmazJxvHS5xtGCYaVplKYEDhUUp9r5
TJ1zJIjhu7/uFnDSuTpUASAVzv2nGq3bzSB2WEP/xEB4KINafzOfBPBhQ7mQ
8Jl3V8P+pCsaPsg5vnqWeQiyGMfXUlePESSUM6W+OxZ8oIu1qDvCGIeGspo5
3qL7p8TsYD4JT6hLHXqmPtlIRmTL6tghpg0eU5IWaC26QawoW11vhgIkpFYg
88KHSBRn4REax0sTA5KaXFDz2h6TpRCd95qPws5C2cY4kKLJqsDIFb1ryhO2
qo0xTBAAQAAMtv40PO4MlHejHfdrtIO9VtlZC3ojEGv8Ezfzzp4s2uGh/IWk
Vn1L6+NVQZOpHNPxYoiArNb/qrCCuXduQ7LdccBtI0Lp6Inm39A/42Ge31Wc
Wx4kbcLQuEkhkAFAbzld7SoEOdZuLZcyNcvPKrBJQifpdLcLsDv08FgdG6Cv
zZPn9DTvSWhjpvkV9OH6m2h+BEbQ5lKeMiOwxnw/VLzuVIqhAWt/dRPJtlED
XDmXl1kLSa6ySidHn++3qiGlys7t5VvETd2qXgwLKEm9qXXWOZodtsOpfMPl
m0UE7i5VuWhBH2Iln7IctJW0GlEC2ojcCQtgCUfX4YsObKfEOFqRgRGD/srO
gTYXnKX83t0fNSSur5kfEfMbmGnmkugQF1Fnjvo4B1em8JsAq10wDJllwDyS
ueH9dWGdUctnEaBexr0fVobPNRxFKGGlfkVmRzOn7OzJNqKShvqHwG9DGwil
gtoSL9GuPQUq+Mg8TKo93DaD7s8aKhe6ncpkZnTzPhGHUphQduDPAOt8qGTg
h9CjXDfyytcCun4npWMD1sUwEOU05CBx2U8iZlcs0etjVuEqg2laaeKkqXbt
gzvFEsH9eeBybCiInNfmVfqe9KkcEYTt1rlMwEnWMq/5X2pjwTtrjOOKAGLQ
TVfKQrLxcBcQP6znoQK96EDe4SMfD7H3r5E2O7mGYV0p6GtSafHL4P92j4jr
WhrC+xwmsep/xW+4btPj6iOaZe9XFCcdjE+xFXZ92oQusUyrUpmq1xgpwsrp
j+80UUrLXWDhxEERoKwJYTe+zUDhOuTRAI9UlcVjO6G5sim3G33zItlDgybs
hrpuAM1M4suwyDj9FGOlXowNDOIvJMmOCAdS0GYW+GAP9UQUMITsxjQxjxfE
AGwCA5iO6TedLeWGX1yt+aq8x6I1QE9U+a09nGxr40ApDgTn56UqU8hpxofy
a9oDldXQocBcyw74+zbYk4EC/nMPugXlGPepR9jpMqLQcMhcL9co3klO9DP/
eMXbzGyAbMKY23QGkeR/8dY1DxC6kYOIQmmND40kKRItKUjdlN3JukD59xk5
/ibkSBLeuJtnvrtEjWuEqlo1lp1m3Tv7Jhp5C1E+7GYBLdTLPHpDXJ/6LLVS
yNBgruyy0jfaBKbFihFQTe5XrQuqqSaDaR4UAPj2HKOIA2oV1lcs0ElqXia0
yBa/BFpyhw6QCaswcVXJyMrGkPsMztiH7cFmhD10oGZiV3Au7qbkGPbNAf8s
mvqqd/JwQDQdP09tz64uccrnpvpscT/QScb4dX62byYBd3ek9sdnwDvF6SGW
mJ3jJVdQI2uFGmJlMvOjfA8KnGVR325snE84HIGld2pUdiaAXmPVCZBjFqDc
1bjX5vwl7cPiMxvPK8gXn23GsNkGosArQlmpl4HBf21vG8Mlpg3ABs5ad2Iu
pu7INjMDL8Q0opaIKH+ihud8Ah3h1YYpHdh1doeZXfrDV+4qDuW3Vz5SpVks
n28UbwFrom3/cNbj+E2X7aI4HGDp6xKVeo/+CF6ReVHB0DSm3zaYx5DSUkfq
GcQUnzK+OmSvB/EedSC4lgzWp0X/kguWrGQ5xv7sk8SJlE5HhD4EdvwLUxBk
peEL/dznNyLZsdXxL3g2o4gw1jBQ91gii9oYyV4BPS7YvpRfBe+E49WSzFKT
r6FVHTADrXd5Q2wQMWHrFUd9QstxSRe9ZX16nLjlcpi3GrOxsO5aOPmRi5KF
aD2a4dq5HKsIDa4iQmPDqcSGMsvv0ZqbKAmTpKN9+ePqWtDN39TayzHPGamO
r+mMfBZqZwdJ5kwQCm7C1aZRkZ8wntvpWy/UV9T50YSMGO1VbIKTrdj7mBQc
N9AOm/+DflrdgTMaZe7eoYeP/O3DykOB3TaTbuEluPx5zHwfgUS9uMaeTvvc
Ogfcoa2nmEgmmUY5417REzcMrN0p/D4q5DL/+901nPXAlU8Grg2he77CQm5y
daCpFqTtKTSkMR13u8iQG+X/LetfBo/QkcHTxGJUk834TBky+tKID/7xj1GK
LSHQaNVHejVZSH31JVekVnuLXq4FBp6g1chBSJms7i1Uw9eSlrgOmXfRy+ho
E1A/RH2jp6INvKPvcOio7gX1hNzQX2xigRphxUqtYoTyh5o6a5mivCWTWF9Y
DIzIybdD0T6qF9Xwf+akQuUXgEoMAkjCvJvvGu1mz8IQJdBmIjWKiFd3Ab6h
kghpq+eryt2zE9NR/IJ3XAeDYb51KqMrrTe+TLx2H8rCbSo9VbtTMwFzJUYw
qqjHq0VfqzIdBD0PCiY9finyYYF2Ha5XAmKFnOAehEBECyY/sGp0B0GQfGsH
fqy9bDaF1y2mFWxFxqChwrZWm2bhKaTATnY/Frg+e3Aw/PwtV1eVAxwWXnKL
SEW0dlL8Efj/Guj/3FL/TJyXHc+oz5clpHXSE/QkRi3iiRBO9fwLK7liIS4t
6Kh2fDEhMkpdA/S0WtnIFYXUzsaRKCsy1Ok44CbW3ryPLfWYOCn4spkDCO2Q
6Kmb9S4OxJ3luQw9myKsC3ZMQ3SFr3q+dCoxa2P/wHjzzugduMkbaReqOOmY
Fx9pjQskT7RPRUyJd8JQIaCyWGYDRtmk8AFTatpjMxY5amBiWJ0ZzJknTalZ
Zd/iXal9+vHEGtxdiNROlY6bEVvEpV0b5UTJlInZOlx8lVX/TEhDf4hvv/Fs
S6QeawQVZLZN5v2gcininRP7EHkS2rPMR2TrV5H5JQLFxX/3M60qBYO0H61c
OPMOt1QB8skO9EhfvYZut5G54CbooQeXLHe6SQ3N6PYUHO0qN0+XneNF7lp+
GL5TY82DJhB8BPWxfOV/O15oFKqhHeySY4P1wKZt9xP90N5/u3QBGFJacfoR
knd0dXSnlIWrHzJwxfyfgUkVilbm5oZ8xxh+/YkEOm08vDlfHVUZk49+92Nc
i1lLbF04z9GCaDINyYwAAyVUJAF6Ypgv3o5TO3MlVRBbw6W222L2z3N/rzDN
1Z9YLdW6bVYy3sdqcRxFaU3ux0zvubd0EQP73Ft9awKtCvObg0zYwEqo1Czq
mixtPxTAb4pWIIXoOKniObRxBPE8LjvUYqUVwgXQrTv1086bkK2J69Ur4oQ0
Bwa/5+NBJglJ/KuOwtDhJbpYQNePY4HSGHRBmBVdqxPhfeNR3CFtcPTICEwp
jazboMzsnCRQ7mBZsWYn9mtFNFlHJbG83NbiYV5Hu3tbUleb+zzmMV3cur42
0Q1/8bc2I8+vEH9EB1IO041VM/CmN3NzA/ac73rPi5vTDWyD5J8uNWeN8MEj
HCFnjQeGVoesMjJ5N4LdR2lS9c1qprXHilc4Ss4p+PT74GSzJUUhqwii6k2Z
rE2HkEdi7AxnQIuHZbyaKiB7Cdk5Ym4EPar/RWiuCnzwyquZB1rnSIvDODeQ
He/kmV6fwvWVgnDCJ/tVfdMHCO1il54S+cmn04fXQBuYzQh48xbSP7ve66D6
CT/gjp1zQudd2k8Gt070elsGqxa/ERzKrGARsKDArXiD5J13JHQz3cKaoc5b
uNYXjyuJNgWUmla3AZR7L4AEMWWou3Nyjn1gZc1IYlztAZvyQStfc5QlI0Hi
8Fo88sSFs1SyiPZxFIjAizytaoXdKWfUprCUKj8fG0YTS5iHd4qEr0DyM9u/
DCb8hSmTJqfmO/FsU/FIL69Yy7J0EnPpoaKTZZdu7whyPQ5Y89qvy5Zy68h4
Shqx2hzpGe1uKZ+gOjMV707n90DltX3zHapzwfq+jLENe2qK/S1M4zJvhzba
Fj/e9Y6IKeXopLF6u2vrKnvMu6Gf+AONa7/r4cbcJP5njroEiyLiddzCP/Nd
D2+ERfz/YV8zh/K9pXVKjRHjeQxFFL+nHpXqCV3xDhqL7tal4KVzW9TS6cqk
oB4d1cM02lFv7f2beXFzSxZqW1a3mPhR38VXkldjsI8L7MkZsgIBbcBiu2Mk
cI5YdmWlfAZO9qgWGMYcj2R+PCJs1RCjoGe0E5sjJNKyE7FwB/sq513D+NBt
JwdLe7pJNqf3r64q9hIpR/0r+R5Y8BUpvPLSImvIWyOyc/Dfqes5xPWtRMYF
2x97UC5gGB3fZOWQ+eYhx/gVTdZYR4PpytY7p4wLUkITVEOLsbXaC7+OJPsy
vcx2PewRrkYa1UUW0VNKI+jfAf+YNnuE0Oh0BbL1DKxCHg0Oh5Ba4OJ+jQvh
fWcebYKBY3Q8mm2pIFjpeUpiNbpaoZcIbcAy6if2g8xXreLNmk0FI/LYntZi
8fYtqEuX7G4M7MZkx+q5AaTDRRTrUWt3BoaLpSTlObZjahjZfiXizBkJKtdX
9447ByAEPp+PTxLK8g1M8UMc2rqWox6/c/SgfAJd39Cymh/WSnF1FC6y+raR
W9d035D8nbApHQiNRAeebwEqPh2MBVsDWqbWzwAOWo+p/TdG6rlAECzo8ps0
rdegvfVkYVTP8zeZC/lk+WbdeXm9/rZTC9F0ZUJttQbEKRQ9CR8QmwWAyH6L
J+KpM8DF8B4UBGJNel29/32tfk8N47obIMMzfcQei7E9WtSrTAt+DD80eXxr
BJ8q/F6bhnp/FqCWO0rJLuyNP3R5odAn9x0/4ty4zniNM2qEwWaxFjv7Rpry
IdObgf9xleLSnqDd9OwXDIuEsb1HmHHZBnyfBlFzzfbbkBCPh/l+cxTrwG27
+6iRC4cptkb/EoPR73A9xJkmUmIkdqm7Gq7PtNiOFBEtcUr6Tlnn7Rs8ojDj
L4VA9Z0p4v8fZOIoVPwdUTWtiaf3pYSsoPd06ZN5s0Kqd3SY7C8rWO2fHW/Y
o2BlVJhMOvMldBIy0fHEDrfiYfwYMPLQD/FpD4upfEMhrB2x98x/jh9cgLM9
yxhTGHZOSOv8P8vgXj7+O7WSofBz5OPjIM7dWjpp2XkxygevNPbN0EnGkDJl
TSHz9C/CO3dPMSQURxZ9HWDorJicA9rl+XjFOZHFdQfAnYUeuX9KV4BK7vnv
rtJRSl68fFBeZwdujmndkWbUdRKFKk1ePY8svFZDOrmCotfSlkeBBqUSV2qr
7SC3U9XDXoVN2zQ0YEgfriSgLTH0CZ08V6csHLEE2vvFp/BaoA+LIRqu3JBi
gzeBU7g9w1mWs80Ivc1EwhXdxKl7MeyH5lqgA+9vtf6rdufLgE49gA7BH2yC
Vuaih327pZLHGosOGs6eIgtYkqrEP/EgMqMWNS8cE8roicIpDYryV2o2YKAF
RndRzAk+857FP9RZjURkNZd/GqNduZamU+S9jejnPV26uCEYy+NhtjZ7+1tE
tG1kLeyFSN27mrT3sFYhaaFrX07cvEy3KcQ2AlBaynnqGDf9xIpetNiVHNom
6ZLKNa7GMdASy6VHBd28WpIViT1+XHopaZJenKoEEOSqm19hAVz//Qz17Ccv
q7nvIL4T7ng61gYXvh7SwbSGTxMzfIWZC1jZjRQOwpthMDGy4tRkbvgLFuti
p5gnwa0GkYMkd7/03zUYUiMphvg6cTkQL1rXel5chekXcBYHfY27YKju4jZl
0nYH7j4wLxg3j4ysaiKPt8yqBRwCBEF/jLMsWsYQHWAA0t/4byLKdrJNeMMb
gVUjcRJPHWb9m7gHL4Vq+MR0wihRYi1g6iss7UiyrL0zwKNr89iEAQdrutMb
mC+oVXW/sEvY6W/7FdmUQ6+70lnHLZaCRHGTblXpoR5Nbdxc7toKzp8AMEZx
NU/A6jyxWcpVDbs+HNhQ6TDlZb+kPhw+PNiATDt9tX4CTgAzMeCDL4XJYq5f
hjMI+xgLT0kDmCgb3dIzPe0tCVUrNW6iakGxqneY66SmaVNpZ8dEjoNkjbmr
hxnWivAGagQFHPNT4bVBjo2eha8Sn8ISFmP/ZuMVB1AwAPD+IAv6A+1iS44S
o8IMwmPbVCDXBXqcgkehpIIhUlHy5h6suqUtQmlquAQQJtnv2t/HrwrYjNEu
8IFr/QTDgNT9d4+fUqbEPbOCC8kj2ACFxv4xNkKzLog6Jt3X2s7F2vwDH9Bq
sZ2a6NZPsIUP6dXU8ZRmr350uj/aQ164/LWIF3LZ+oYA5H5wQtd37nJwZVqm
TGPcPvsifbTSyXs+njkYy7p8xCFYeTTI07xfvjSH5ADq+wnXUJpf5m11W2Vw
eJ0xrLjVGYJ3q4W/Dd93Pi6iajk5nq9xq9ApLK8tzROJUVJ8MbtxMkRDr8C1
96bIsqqN7jE9m1KbKIQd0HfIER4U/DKL1CxhvkZCgLZXoJn1+l0N/ZcoXZ6N
JlS5EnkWYdV0DT1f2K6+TxQVmLnBDvEI2WmqX48byLbs0LWcqd5gHGCHBBOt
52DsxePIzIBwN/U9m8Zbhr7b/O9Fyyn2tj+AB7+aR9Y0DRQQ/HpuaUg61jUE
o1pq46Myj8FvKmzZlNqHfqDbQgWT/8jfHgtdmLY4JbzTimCtcJHBjnni7Qtl
KQd4JaDauT3JsVDU+ZWyTj1hpzMErHoIFNOzj27ULB5bIGUSpqETZSw8NT1Q
55erDA8WHI0wFFgd+oEJGs1AdYKVz/ACiV4wSmzCucK4WeqnKxe/vHpqqFU3
yNK9Ns61/qhZQqmWt9e22F6f4yauqkzwn+yHGVZB0/WHSn0q5d4YBxCAFDQg
XMugc7aBwHqrRAJIyyodr13optqErOEXobACfEMbB83HMquPYpvZV7bjb75C
+BNo3JlAu9ZWmpzgX0EIa5orhAXV/iB5QNVyjaBu4FhdTzpU4eYtIH0ZmKN+
dRqFG/H5u4MCSATAjpB7KziRD0dlVKzQW5wVw+3oFiijNQzcm2gnWFmafW+C
+cd54pt4aw1gu1bJo6Bju9SY7c3haIh7H5oCfzE2wStxwnSzKWiOx/b8Zh5r
tW2XpPvD5s3K9bvFFC5vlZX8WRaurK+AhGNmsVxJTIl2oCNxdVJlcn/2UaEQ
jChUXnML80qktmnb+s54lyK1lKpbtZRWQ0tdnTQa819IZp4e+TzLpKXky0rg
zOPiIleA/ifT2DO+uM9IDu/dV+hR2Xcs2sGQ2Sg7VT2IWlgG2w77phX/ozVl
OMEBha30L1c8cHL/yLEEBYcQsycuETD+KfY5yfoXsz/Kwc6R1yUrFf/0ru1l
T2fc92+/NN+G5VdPPlxevTab1CeBUsu5qqJIuDldiIwEUCv9IylbhWsysR7t
WyiLzO0+MCHE5tJXU0wZzBIcCVLAiFziwaIiTOhMhIJeHaJNRAMtZCpoClCH
nLMQerxr4mb0V6pVfSPU2DJ5UsRHBRBGnq8JeKcDw6+F/rEV+8FoXK+4H8aA
yo5EwExnXN0NyUDk84EI3Q+uqvEZ6hujIggujBELRlovvH93iAWGwaREwuXu
0bVcuo8iaAsvxZwZCumcd8CcFMYB4UkHD8RcddRjQbB1zW4XB59SlJ5fqpUj
tR3GWR0bNwJCELFsWQxiRdKfVRioFqu7yVTvxaFPH3rS5OekzM7mGM9fzRc3
sh/c6U98fNeiIEoY80V42X3SCOAW4q+hEVfpxeTD1TbaaM51xlg0SiTo81vK
R1ISRZtwy8QHunXMZsZ6+xl91x5kZzEkF4feuOnf5VZIDqAc7XTn5f3yVjXB
rgvTqLxaSvw33mfZoW4Pe1mHUV59iTu/rRLYkIMqP2fsS967iY9MHNAIsri9
GQqJvp0UGzL5tPGwFkXSHmxKResgWoO2eHtq0JG91H0a0MPum/0O58zPBJUh
YG6BKLBjDKBbB0ZscXfruYhVuQni76rsxyLo6aS9Wd0/7Dkv8HnABB5gKDwm
rcHEHeqgR6ksyY8IXIPMrBNKKrOEZ9vjWW1tBwTxwD50C7yYHGR8GkHswwBA
GbVB6WWjX/qSL0S2ypxgLsE3Q45gTNe73ApPlZWpAZMLMr9y1Gg3UI1YE+Q5
sozI9MsN+fS58hzu6+1vbcXmmilFvFp4+Y4jCRLtQJNBDLkfbblttYcYLBcb
IrezvT+zJiMHx2av/MELuCFybb+SROsWclFkhmBNYyMHscrKevD4ckltDvEA
+s72dSf9qK2jHDxRjHEPhOhB1tiKJyFEp8e5l2vJ4xKZ7cWdmIVcm2QJ9VKR
ul/N0xSMR7P0Jg4qDlIteVxFDoiCm8W7RPEu0gonrf3WqUfM1skZYi5WcaBg
+RcEkonvZ6B82S1M2vh6KOs2VJStwmvyAb3aZBrnU9cY53/cAZUxQ0Uoq26C
o/AfS+KvbTonCa/C7vNR1V650UGCbyRGtHJd98qwVJaOOHvsNE5+vzjIwg2S
A7PsU01Z3APlufYNK95z8LrhTJX/7Od6AN9XuUqewgNnrJm20ks7JmA7vIvN
tDNXP/uL01oYDkMgt5rflQ904XryfemQUcw9ifIN2cDrD5ax0FuUT78jhqmG
XexgT/thEmFnwzNkX9ISLJvbD4VYGuZn1cMBEnR8rEJnGOqH/vibDfbJjo7c
tcMhArrhV6C2k5VPAPVqw7ZnxSlLepmYpTEP5P3073Lir2qArMkUhXIIz0oF
Fo7O+5vULKCRA54xLlLJELRdnixbEql1/OBqOhc3//p2DUqBECyE4wO1/DV0
rVI9/1a3tGKDD7XqpM03rfT7AgJ3NbkwCY5qiTBraOEHBWM4J6pBm2yWOEOo
8WnJOfWXa2+N6oRSYVFhldLrREFQWuVRqI/HuippGwQlcYvLCPeLeBmvUuMh
5wwldipkeRk+Xs/yykABML6RIS3XBghKwwaVlJaHiM+WsHpwMcOh9fqm8di6
OkZPC3vHoeLKArLyjVw8qmVaY7ePynNgjp4vnnSkzvKfJucpcoi+kOok44nF
OjnrwWLaIf64/5gZHdQbYkIPVzfqYi0Kb2Y1vDbFfzYri17Oa2IcTkioa/1j
Nt1yyj6Jh9WQHhwWWd2RddGqJAezKxNMKcDC/F3eZ0Py5mSBsrKYp3Mp2ErX
PkoZCY1nAETncqKIFc0DRQcDg9H8FEowyUFu758apgJ82pmfnGOJF6IYE5Qf
snfWawkIfmuk1lXe65bd+f6bcmWvMjKwG1XCIzVjUxtdHo9neyPzWh7PoXT/
blv99Y4MPwq7DE1Shjy9beHj1bB26SpyhD6HjK3M6zhoHYHUIH2ViTNzpLYw
MO8ZKvnUNzP8dHdr07dp+fc8OGXKb+AiyXnrlXMs4tswwzs/QKaZupkGt37a
eJY96gEDtHHKEQ43t53UrBfw1t6HK4Lc10i0UpCmWj12hNnQepDghKOUtFbT
PQKywAK1WCNUTwNWF+7KRHkQjcdJjxalxS5a2UJ5R4O47yPKn2wEkBi4vBkE
XsD+BAuiL597k/3vZNYTp+39xsJjVy2Uhc3aOSm9F04L8nj8S/MzMgZgIbc/
1Ewg0kdmDqK0m082t6Eb5QhkrdmNe65BhRbnJ3+X4r+lf+s7aaSmtpi1aBhW
ra0b5kyHY6c+KaCsgMZvOw1dAqNBfcmgoeCfmcdd9OqTdlogVx1U1fk+QzhT
OdZ5DAMgEeLTTxRPKXk14XVJwYoeYYpDdI3fgyRq/mHJ31ZZwDlKFXxXYpp7
BvN0RqQjLWFfHmgbtylmw/13TscBnrMxxCbpnR5o25pWQmQZKTtFMBTyApPE
KQc90eUisM2ut9Vnj3+5BZj0ULyJqCujYpnDnREV1Yrxg9oMi6HbwnnYr2+J
WzITzEtSEnZm2POyqv68kdxhP0YOpoMMkZzPulWa2ySqKTto79tF0eZJ4yPJ
fBkpnQlWTNT0/uRFI3eQI2qzThPFOwavLpi89+W+u9EHtbkvh5+0znrYyiju
I8PTu8o4RVs1GnT5ugla+ncwdN+XY2X9TOaFiZllDwLULlItrndTfrIBuKqH
vDXZrH6jWjRtXPxSQ150Cld8Qo08kq2nwR1tfM5En9Ie6QdC8DILfY+FfAhW
oELIMbb1tvP+k8tYbDZ/idhHvvvn/VdcF0KAAJ0oJBrq3gksF15YX8bCBUic
9G69PlkVLJVQDZ+xRY+GxWlwX+VIi9VYfCh/Clqu7G4mt2sK6Nz+8cWkPLdu
Xnq3nOHQCuNUtsbcmHaC0IalckViKls+fXCDeLk3IcBeesm9eIsQ7DCg7VCK
BICe7M/113lt2+DMbe3mzuCTcUov9Cbexa64XKSqwQtA3kHZ1UkcDAFhb9fO
jtARoCwqVdSruE8Hkg97zjWEQxZiICdiq2CjmfpWgWLz4QJtx8upEhqZIkEg
mQCswV8J5GFxBQZ7crnibshRHHWK1UVK498f7DME5osgwNPOIGv+e4zWjlwP
VGeuHYWWvrtXM79fLy+yTm2in2wsvdFhzmWGwsFwwVtQ4pjJC8J86gjAD4uy
HVl+hePZzwcL02iyG4vsOT34io7kUf88MvmW9IgV2MLrZTGbOZd2U6NgtYq8
nAvRMRQ0MBXzZLRvL7kGc42iq09F5GU1305Wrv6/Yyut2R+Sz52XVKOs7cKU
oWT6+Qacn9mXFcsLaUWDZOGWSELZiR05K7reaSFcP3n2aHPTBaz29yeTEch7
cLxwrtEedZxlAIoCG7wjC1ML2z9iP4Jp/aw2VGgKWtfRMn5f8/SblcQdYeQ+
PkrnLNhFOVS15O+bk/iByIMINf3Bn2ulDUAwOhBz9MBDOFkF+GUGkxzmDjRD
jtw6lehvIU0M/xzCAWGX7gjKcJlT1pathQ0POSGpsqNxCJmkTm2OBF5iu7ei
F32OEAh6NE26v01IqPBBbx+TlbrOXW4xsQATbnT4+EYST1lcTM4Pp53IQlth
dNyC7iUPYfxXzahEgcpvu3ZUdODlnZeym/ctmp66sLXZyHj9MlsFrO5pUkIB
pP1X1KkByP6EIGMHaCfVyRFeI1x6k43WNveZu4iK2s9iKjnCEywiP+d4mMnA
RDFxcwzKzCHpOrzXZKlSXrOGxlSxwL+pz7svKkDpa/ibS48t3dPMZCsjDjGh
s+lq65HD38w47OK/mHze00sAcekihdm2Gh/gM9AoEL7k6nnNG56LD5FAqVVr
Z2U46KPoopXwCexcB0B9dscXJLRcjdkmM6FPNC7x9cfSEFO/kAgFx3K7/xkz
VnLzwWZ7JXdKRIdeo0fiEuf6Rkxn0VDP2jb3YqE+CtqrlM7Jd+0FuZjBz5L8
JqBksPFc2nDXxCXO+DyVxXT56R2+oCFhp4tyXgJNIwGv5U/OEE/YftG7kfsc
aoGziq+fTe5GPaNVO1bI/EURPDBsbU8yC1ClgLGHEc1nwVt6MViENTPtlWnl
z6hLremwdyOpIgljCnv6xZbpXtDjvmPct8DiCnWF12tX65fXkeuzfTKAjD9Z
Rh/2lYpukZECtfJxTZewAz8x08jvmwnmK3bM8oVkRGkwOR1xYkucufcvLBp6
bOQMQy1mgPshLcScU2Z4fZVL9lPhwR1y9ZENBHQC2Uj/8tD1H3l2OhZnOkeB
gVpJlLxJG9MdLZuJe/GtXlOR+WajbnlVZ0eND/SNFUI//bPovTypFHp/DfZB
Cab4/lsvhDHt8qrUdCxTT57TRozCc0QDdyzT/Up1c4YcvvkIP0mi1KajczLc
OUAuOIpUbPKAFxErLM5cRrRW92v6e5vrhnXF1ItZQ2nB/xEbp0FDQEKYB/jg
9K5w2Gmmgt5zAQA6ubE6XUsGLaPZ5EYjUACqkzFaMrrKWHbqIqsZvqqMfOAB
8JdH+z0gxFemG0d8JxY7oaBSmARYoWkjgVb1N1jFR9qkduLuogUhP7M3VT2h
AcxpihmUqWjgLH7x9iHSq9fDFOFvO8Xh0an/Q9F+RyE+OlqVdhCjdMuPa0xH
iFkGn8I8BKnaxUsNIU/lPwX9MQqDIlzS2lUsuCShOhMYSNzA1WsJyC3YGtxq
3sSX9fFEW+54capZOOsmXUINUQWRw+Hlsepw5kOyjuBeTs4Ezzh2TUMd/9DR
bAY2RGqmQCpro4MRGjOOUk0hWvErCKtUNho6+WqzqYOIKyndy4nLEUAySc4G
h9oiQIaUZP8SB+ZhrcOxsjugFWu6MZ2I+lJxyf9WGLE/UxE9iskqFRAJWq16
hSC7s4pydVPipzt3IPUCIZYMs1TxGw1C+rtA7mbTtLk1gooRNA9hdXEAHkQD
DYmEHhAnMbk0pM/Sn00ZI1551+FRFZDkx0GXGEPDQ6g6MoTon8c2P+rRvyDn
5Hmug3hr8yQSJedSXjH57kPQR+g3Lu56r8blZ2O4JgBkIZb4Svf/OGO/MIh/
4RnO04buHuvAUGmZugsuxna5JYN9IbsAkR7Wrmvy/JJru8xTOmP2SkMHveX+
JMdcBtkA+XnlSYReOeseAnOKB7d6T4eJRZ28jLjhO9cvn0/ieqG6WQme/kik
Yip8ZidHJEBjnDVp/zP3r9LpbtnnvlVoiw8QP4D1Wg2Hf5XCiPWmODHmeGm4
TuY0N+ol7buKZRwRcp7kwuYYd+6N/IeDPMnbyvJLK6TqzHPS4Jy14Hil5K4P
SOeAEUdAF3a4zalszWY3nRr22CFbE0liJU/um2QTWRL8jRF+taDfiE80QRlf
zm7l/ie+Qnf1uZZzMauLrpEzX5I6aa/+GOOdm5/omdfAmg5llwKIRDS/IiEt
BCiebNey64NsPNa5hQCSmuXo+mYWWOcPMeUA7Gf/ff3V8o+Fj0VxDedWMiE1
jPEVnbtwDkt9okinvFuWvZswpqPjE4v38+BJINeJjqVqQh28Q354KXWUSJuF
wiqwYANfRAGkkuR4k0XhhZ0wWSbVjQm0Z0BT8lN4hlapQHhffOW4Qb29/CAa
aXI0igaCRA0PcvflB26Cif5tQYQYjMMTGMSUrd77+sWu7K7tOdvT2nQOoRTF
2y+VA7h1YkjPZL+VWXyJYrl54RKyY3qgXg+KEKswixKQA1QskZmXKx18j3Nn
t2Jxb0uMxJI0410I0hxhV6YlIopmFJnz5xSnandyxE6b50Cd1ON3yjAoNaeA
fAzN051DB0+dWPv7AmHDUC+YZuAK/hILejo9E7D296sQ2QO1IziMFSwyTiU4
G2AxMo/oGOXgbxT+wXgxHAanvGCeaHOEjG2OBWjmGHVltuYuA94cMw131681
d7tGTCAF2OlKfHTQO4RGRX2bcHTU3Y4AN5Ztddw1kqUxPBQsWviAg8oka+x8
65qYyAJF3H1dCDo4C3BQ6ETvt7zWnNqCY8ctxyeMkI6BvVmVYYyzep1LswSq
wTEWWYE2HT0sD7FyuoReWbqojmJdH+zUrkfhxtdr113ctcS8Gynb3GfaE+cf
XD3LS8Ux+1kAYVLyCtnD8zGkMZJyvmzsOceNs5MOEjABSs4hQvUncoRz1bVQ
HMPP2FGqJlXbo4N31LE6825l0mf86/+XvQbOy++2h+eet8Cce4zG30rYbz8t
YgZrpAAGCkv3unW6iSmandOWctUxTC2ueQ3YX0bvbcUanC3rN1UKYcCRD4Yz
fjgzpxJPvdYtlSUDK7hAl43zPD8Y3LIA363QkCRsHIrHpaKip+Y3nacrG7lj
DA8O+OSU1AU57tHUz1OhczRlVhblC2gyzICIv0vofr8bQvV1TXLfii2JCkPL
s6yPizZcPj5kOjYqOGvYypTo9JKDWd9Bp3HzjBD0R04ikWX0Od6PNaaJQm+Y
ehnpF2woLwIucFFXEI4rR4wC4ZgxWG03ewsUU/wJnYCwvHkcVi8H2kSpov+7
qLVzOETrepftiBF/928G/IMofNriM74R9nrhq9QVEmzC1UKRpE4BXhGenU+/
Di0pOpsR1TatnIFQwd+3ZcFPxdCs/Tl+9NsDMyW/4rb6x5ddYHjoveFk60Bc
iR3QfnhMAvK+jahfwBcnCpvyiws6Dzwm4WjQaKXUYOPgTIqGDba+7DLXqdpN
pKRF90xYzEQTGkNDIUm6UMHmEK1EeUy1ZksW12dXh5rayo4Hcer/fsxtQeOL
h0Xixe3ojVay3lzxAZXi3XrRZbsc65sPUGFfI/ehnrSW1i7/Xq1qCKiZPilx
dNtwfonfpFPaX+cpU48MYYtqjhlkYtPP1/k0KWGOTNTH0YYUC/whvTGQBHgM
X9lJeSGV4C6mDHUBBoTLPdgT3K75E7c95d5GLtq2xd8HCWvKOzaUmiBq6Uvs
N2euNb1wGjfCMIx5oWYwxBRyFyamAeywTnd3rJcD+UPllkcPImG1kIxob47K
VzdBsDRwF+JWSCKG8gSVvDC9uhG98VeRH+fj1ui/hqV1M5pT+a+U97LsjSgE
Gt1fxRqvMlvjU4yGMo3DYmbw92sh9sv0TdLL4sYAC48TLJ1df+WIKIw0Harr
b/3eMMcVK//ZsB1RwC9dGyH9iqP8suu9N7YRw3Q/cXDMIo2eufQ4+GfiuzsU
ROuPI1gaiqxhIwWXffpG51B+xMcpQOmtNZVf3wLJoUl2xi15r9+FaX8LZar4
ioL4CycxOX7S6OIbj9UO7p73ElD9tVYeYvQ3VKavKrXtbZGzjbnr4rpZtH4k
qe9q3RRDVy5U9v8wA1LmV8itNo73+tj91NGV7XKnjcQECoRKp57uUoV1NTL1
L3D6tO3z8AH9M1Uc2EHalyXBwL38HBIsxr00BJq8vWUzvIUsv/F7fLpzmK7r
hbuHoNj9S9qQaBzGCIR3dxGEe+s9mwKNHXdVMoGoBz7zWcThgSiyr6CCKUxa
8Q4pb/SFtr6cjXbjqhC6GUEEr328Q2kwW9xnC3hdD5LU3oJrjFTBIxP6h3Tq
wLGnU0IDX/+o5zYC90xCKkoZRkn2Qzq1J9x067Yl1NKPzSpxTPXDhVHNm/ZG
qyT07+KhD14EX68A6gjpFhX5jAxN57nUgQsPeHgx7/uF4aUJGmCbfPY+CUAJ
KOq5VQny1ZKOgZ8RdbOAbzAfcD7LrlnVhKF1OI2AKO73vOHDobPRo8H35idG
is/o3EZY3SOpbs7n/GhRWBhCX1HoRwanfpIXRZviVn+AoB4zbdAHaYZzKi8c
jD49DAmH6kExyHqbTr5vu/YK/CuSLjSv4TKdc6CBaDuZJTChyOxt5eY+pUTl
ftZSYTGqg22wOrFdzO05lAon/GIlOkBx8DGTPMma4AvTunTcHXGqqSmywPuk
5If69nRagYpTmqs1WiZPd1fmeXO2Nm+OX5kDBeyFOuF/j/+ND/qFV6AxaTvO
bGil05IhbAk6ZLr0dxakiNOJRX95v85nIpVYEZh6vJtgNI8CNIMx729GSl5j
H8r53Vv4IfNniaWHRPezmiib6sP0xNzHVtLadAQ0neWsedrOBoJ0YVkhB3Rd
6ZO57bEGMGNMCcnocpW6Nz5v9Xz3tQuBLGFf7sIPMmh/MNQ6MaG12Sq9JjLc
vOvCmvnX66bpqkdpaYpCWyktKgvxHwwe2ZcRQzE0zGuFAIT9mkOkAy0o+3OP
z+DDDROzzJp0xz4eQZbGDI8mgbjB9JU5cgX6kugY8db8m9yaIY7xdZwGM3bi
3QVpcloH9Whiadqv+8g3/g6BvWLZL6iHWPmfDw5hZW1NN7pam8cuLZJxuQv1
bPHw4dvhNyzZfZ0tlNKXUw3xAO74MfK8E1dXefHQZ0n8UWsqpeyPlaKKWXOr
JohHowrLTJa1OUnvKmxJYvS05/itdyegmja4LiRDFRnpWdm9gMHB+hEua8o2
C40y+XdAVCgIpYUWrFF6QXvNYzb6QRYP3U9Er+x37yvXHsqV+oa9S6LxcwSf
F1rmCUQviWn9Q+5b10oq3WGjgmeRXZjXBZDiBCKMMYm3iPwyvILJ3ZFUvKYt
Y5p/EFnpXJe7eX+0LEDU7Mh4vbjL/QUeCudMJ5J1yQQAHr9hE8Ig6uQ8HlVI
AlACFIY2rJ6N1mOuZfCKUqsZGpwDtHvMV+ntMZhAjhBt1ALyuwSbXX42hOik
mBYd2VzWP38hWpkSS45K2XdBFQdCTYAtlvNbxhYgGp8avztd9xQwlQFCudk7
7/wMo5a/AcP++KtOWSz8icaCMJDc1F6qEKLCZkU/k5b8OuCVH9FaDsmTlhVB
C8ibtIHOgtpbSxY1Dp9FPWzS7jXL0TMVGaKgVT1N3uGxQ1NwO0GKWfH0XiGr
NcJxEAwrjAn5jmOvWdLnc1x57s/PgtcTtbqSi1eX0bxhEvFY2SDFmEow9+DS
/p19KzS1LtDn25KAR3NPyawN9TPAw7G2qZ60wMYkrFoh4yHwfI/k3nLXaC9+
6CpueI9fKsomm/PReeo8J+Io2nefCIqAe1OsmrD4qQMlemq53GS53FJwlgsq
e38Jo7OyEOSUENGycQD1CTUqKtawCUz7eY4fBGuqQ/yLusIr9h1ru8EUTscm
rfb08qrt0DjoyDSIpYd51KfSSMUxNzl4lqSf3u2LgYCHa3zheKmkAKanwdsW
/8CYtZ0AOlQWYnQ1Izg0TNaipXOEwPcHIy17UgwNOu6tNst5dGI9BaGBUyfg
dWtMQFw2DGdqGitwyl2K1VvQwLAN4+jlx1LW9uho5TSrxXK52kkpq+/ZO4l7
uAleln9+92CqyyuznE82WbBPnqomgFaSUoXD+27VaveFPqC9lAaKUsobQ3TN
CSzVql+3Bqq1zTQ2ORoQLfbNI6vnqUoqKcwNYOWrYobGVVd4GVX0fdtbCR3A
Gn+fpw9t3c21+yXfduogKCWDJf98iVLvgRj5fuubGJXY97ogD6yfbvnYQAOx
Z5xDh4sSlFDbYpkTrpqT7RmWphosGxwmQi2NiIdLaMpcyNTWFWsbWrWOWi4l
Czwgr8gv8s+88rnRs1Yu0bGxkBChlWIkfQ91qojJv+zsQcPFNwR/SmI37Pzd
yX71bbukL9sVPeQ+3KEqfGEXxlKqe16BwNPm5Sv3/G4zarzIJ97dO4xzif7T
5m8aCVZVgKqeUwnzUhk3D2IdKuLlBEWH5OFgoWxbkWrYUxStYN5toZ8KKdZN
PWcap9DPaSHw/twxGY3IZ7ovjLsZSorVnjgS7qpI8SeuVWeG4IiOHDcuwduJ
AoCqGV+nx8OKtWbjEmTbu5LKB2TQdx8pHcPBC2ngfZrJfTGEVB7HhL2WoT/p
EC8S7zdLg0iuaolI2ymI7qWLyudp2bK/IvGrqSmGkqR7sVJjCm6pLE7pva+9
DtHOAiNlZVy4i3B+RlYyBvzUmrxEq1GQzTIFPux+KlDM9koyM9IN0l29mt7W
DIt4e7bf7ZiLemwzvRh7jXtFWTnK2zaopyRmAMMm0Jtw8DAqF2zY8tBNrFqW
V4AZEoK5ettrnFs51osZk2bnnx/oY1GSCdIFzczQ0M/pf7bP8sAeMVdnzkmS
KsKdPJB9dxshVRabwo27MQApKOmrRR0s1+2Nkiut/hTGMorsvFaCwteS/1GL
eu5OP5MrI1FUuUWEZuiz6NNGSqDe2bEVagNaQ+1RsLP3p2+wy5/XCcysMby0
maLPz/QHRGTMcjIO2YL2YEB3BHhLHeOVie2tqnyXY5I2UT2JGxpVTqfK/J0V
IYhM4C7YhRqQJBSZa70bRUgJZ5OdJoh+w16nbT+LsXXCzslFmUZWq1SzZm0d
aV+TErX4ydiWb/eXlz0qIUf0PUThwFGi6vkuVvirJXR3FY7LI/pPWkgGmTD9
8sV8XUdawttKoijE9P1WceMVE48NFwlsEkvb1VN9DylUsF85rE3rVVW2NNnr
yhzsQXDDOBHAF/SlfSa2ra4dzrV0gHHQveYTKC0FLNfVN8R3pCv9YlzlZUyA
x854berj21f7RpHWRQDhrSGW3MPDOhNNKHrl3YeAxuLZ7yXGxrsbVjeRoI7U
Uneb/a4wceMWdfk5+iRQUm/Hvyzfe4WrSzvnXpX5CaKw1p5hImFp8CJ2tfiv
ie990vyy/SQvtCjVIS+JCq+yaYPCZBJOIah/SF0QeiAd5kteoMVM4nP50A+8
azRDwT6dRv40w599ncyBHlZ8B5b+D6VEPDgZGAR5ixRkmw7VgtCpg84JHNmL
lyvx12H0YAUFxoJCxDjMBJilnBYsTINaI/jo9aZG5w0ZaAUhBDP8uvp9knBi
YW273iR43sPBqDXaCOTvO6EaRRH08w0/iuzwcb8Snn9nA9Mt1pVBHAul3ccI
FykEkS1FlBoRF128XbYnaieWi+owmHW6RXg6e6KiIGuRTOIrVpIaUA9dtf5P
u1sfXTkQBl8IOiiI2SEvcOtT8b5rMKuUwS6deQR1aPA7oqz3XfrB7C2E1/zP
9WCkUxgGEBBDf16qglDW1gJflGpMpyGJ6ZZ/unnul7igQ4OAoyEe6o+KTSIt
QFADerbYcnvF74Ac4OxR/6j0AP49HeuzB8cNmUzWJrzjDbJNa3GkkrL01x2R
S2o49NTk8UbOR9kiek+rIsf7Pc2S/dDEYCLFlBV50KeOL/TVBdp7a84WUTYp
5u2XFTF+8VfvwELM+LjJeQx5TTdY3XpnxUc5FcIxt6m/FIOit4UAVyUr6Ulv
x9xeJBphoSc79feQ1fL8DH730siRZXXaJUy9p4expwtr6eWPEn27rUq5+p9Y
MYo2YjUV2wFXzlWHi8iKbUw6kl7BDZPk5Q2pVkVwtO+rTjjivvvYkGYqcS46
2qtX/xnLzxyZz0UUc1/ii7by3lwVOOWEoy8I8Rls+MeqCX+03Q7z/qv3qFgp
mzmAp+sKqhCuAku/PPj478Lsg+8eWLviqgtQBGz6Wf1B1X6uqNSYZ7Cl51Wr
aYq4Lccwt5PKiXOiaqYT8DngCyx3lGy8D7NG5TbWDV8Bplj99WYmj4cFxVNx
JbSvGsknr+z8eTCQJEsjRAsCWw1w6Mfk9eZlvJRKSZnw9LQuYqvYsZlXdJBY
f/aDETKdQRhnveZH83Ui/q3z+F1ZyVO7cge9OGKejAHSFtSYuJstVVraCFV7
Gik+dgDH6shykc9vg8MOcF8ERukcPTvxyOwkhtomjt+tNt0A4Gvj882OHpwy
/ADUY9WZdCtD8ztwvJ5oSz1ET/trHuc8J+bmAFhSalTbW0w5GwMl3ZV2wlJi
kJhf6+BfOm1+4nuJcVJfI2Gt8MefmwAJjBhZVhJxfBISv86cYfLBmL1CKkFJ
EAoMIUMl5HVmrGTbJGvoenVIS1okkx5nLe8v7PfjyQsTmeMkLhVMX9oF2Wtr
ZoaEzRL/jrFG9XgTkjAZ5V7wdX2IRgsF/Uu3Bvrt+AjNtrN8Iy+shvN1wuvx
i8Tlf5oCbfCnByTSRWWrb9P4lP+mnjjicNFC3Zkzd+C4b3MyjvDwPuaSH44i
v8czqR0/hvNF/11QfSuG0zNGf6Geq/8GCOKrUeAWqAe1cmBDtqR95eRoLP4H
tFP2qNRsJbXrDvBp/mp8HKvQ/bVxo+r+tA1fRT+V4q3gyv4jlmRiXPxWiER+
I9pIQA6lQLg/qPzzPeg4zCDmJ7Cd7phyfSyv+umP3EsH22pOmwlA7bLbxBNE
D46tSVtlfubDC7kWlwj4F4Lg8cY5gPeDmr2dP2JB41uxPAupNOM/bfON3Fzl
6ufGxx3GkAjQpcCLbgAXJzn48rf4VIcAeDJbj4CCFc2OpsJkR2Xk+AziwauF
jGKl8/zvi/957spYiVuWr9XDsybfOgnx5m5iRhR3GHy5/mI9KRzyY0EuIz3o
Nu4TtpaFmueuJGvNfjUSM1SK9keSBU+SWkHMHqnnfpSYU82MSEz9WhotKcaJ
+ciEwdPu21V4xkAtSZ7m++FCmAmFvISjvIMsiZ9T1dgehCh+9HbSR3xVwCdD
0JdT1+fR+DDZ74+H/FrADNITnKEwf1OXiv/RcBgsmHK77ApjjDEweL6t/xMG
vDai2/6tgNnRnRSY/5up0tor87DkoLhiAud9n1OTJiYX+JaJEuoQKZ2L9KE8
WziPi1BvTTovOIgr9gUPDPhsL33EDSdFTXc9rqyHv356nwqUM3wUNQl+LHsq
mXguLVXp/DJHNQK9nSchsuYZz1PFZODqq/6dlaN5xzob2jAtu1F02MOP/HRg
bYyBbQhPKiHifmXzDbRA09OoFKeuE4cylaAOKXkTO6RssSo4SDDSiDF+A8ou
b4YncB7BvRGZGPjpWkOpR6gznJjpumU4C3ZIcvYVnJ/cLRQaq6CNeAh1wvGa
Pna+wz8L/I0m40u7E+HP+whAHuuT3fVQUUKL4PVfm9lmo0wN1ghG8nJhXYK9
pCMxK5poYIOn+jFrmQA9rd+frfS8gaPBukjV9TnCCVkMDHVSEAydxSXRvAoh
l1SFgfmB/WRubzkIeyulxAi4iPN+mtkOTBByszIzQkS4Oeo1hrhAcz5mu31r
hjWIsMf9SqYtD9u1SrpyNhWitIj6HlZPxlA+YA2r7zfHPF7kleVNjw/wNFpY
nS7jerlySu6URzcXhuNVbkLePjSnizWzn/aD5HfiYVc3oIqzupSW4l3O6mLG
7/VlCo/PiLy+wbEmNI5aVGy+pUGbaCSyIy642V9xDr3pAfeY4k/1bWPbuVSD
3UtcIdnd1UfoqfNYJ6OrSGfHUmfyBiI2Fc2Imgah9TOfl7Z7A0YjEtg5UoFB
fV0DR7VPAYEJhSJtyXkK6IF5bvYLvHJQHT4YpRQLnJD+ySMf8wR93exlbXGD
QIDgvfMseKsw0Wzwwun86uA0EfiII2O4vw3iLhAXj3Hnw5CQD4AIaunOTHzY
nvsRO8MU5bXx+3zi6nCys8Gy1NTCJIPjOOa5pWo6XqWua6hse7nw6mJOIY5Y
rsX9xVf4imG70IcXBRZcEk1UEYGZlLWzrgztRB4Mxf7l0T2EUDJkNnZkmkQM
2W/bw01KZWDbfxqF4s2cYrjUbSewOKDLjCgJd8cxC1YbA3mcPXPq5lTq/HZ5
NWKc/AuqCFovcUCFO6Qeldfx/guSTzMmzBNWPEvTYzrpOJK8aSwwm1OpOSao
wVNayKq6w7X+Ecyt1DOw/1IChT+sgSVj802WlFfcUq5ZW2NZw9QbAiLFxLr6
uTFsRghCqrLJwelf0dw81nTuysbs8Crw7UHYs9Ebkl/2DUmBd0uV26FjCizq
6CXxydeggRwFxxZl0OyjTtN1oQhUuvqUOZ1UucW00xUkmT4J+P7+bpRQz18v
uy8hpAofzQcY8DBMzRATFVSXwOLoWHCHp7MW/557zel8mPuyGhqrae9kO8XB
JYs83vECja/AApsuxT55XEWmYlOYtvXiOHst4ZlE4JuFdtVNqUnEIpnSMf0w
g/yHUv6x41VNpAlGT/MvK/7B/+frl329JKYOUFnpC+mQbhHJ5u4OHoF6BoLn
XJY3IW74U/7vWD7J7nbuMrLx41iwu5bFbBOvDF2xHyjqpR/JoCNnKlKEx/OB
275ZhABjYPU2QQp5YZPBWOWlaoUTKL8vwlC9OwmcT6ZOeFXTni07U4Gx0Bve
sbng13nXgt4ymB8uJBbFMkhLFFPLldyH74Vw1oPk/6BnUZsftFbofXstNcmM
7suSzLvoWE7SpsDICJg6nxaTMbxQKu1GxA6znV14Y9ck86nJt0088yCmL6vD
Xeap9jMAZjUXHSDRUvmXV4Clu4xO8/VuuLgCNymrLfFSCLBe1JGKUecG3wI1
fYOQyNaDkpq5k11RwXjBotBC2RYQeAbeVh3rBAJv/NU4wSKN67Zy/WNxTi5M
6thFJnwBqDH0RXgJalJIutgRIfWn1i8qXTC6psnhz825CNLxYndWnp3DnqL7
JI+QrqWr1qpcGiIKXUlrKkZ+9i+XitCGIBTAOLnYZMvTNgCoBQ7m+20LIekH
fBRUk8TtlEG/Xf8aD2CAXFdxWFYC0RKC6bYqQmLvacAsqj0ukf4sh3UgCYGT
4naTL1yXFMWND0SxvlCkTpjEzCZAOY7emJppPm7LVZk+shwxaySrFEwbHpa5
CVL7vt0Sw2nKdMvGAd5exNfL/vtL5EKQBojPIarUZ4v0BwYhxeK6XiFaROK7
TibkgURElAFddwy/qDSdSgGHl4zAhcxPMiqMrn4oD7ZIPfoJ9TrOtoy0A4y8
jnbTp8fK0+8fk2ey/5bwDUvCJYnd4DL7huhg6tA+xgZbgs+Mudyh6MFXYrfR
ZZynHUZ+bQFQ6NIlfFj3qWHLW/UUyifjjcQUiqKOi1l37mjew25hc1jIpx08
63b7/MgUlWVBt9gXfXsg0IwSpBtkaQwpY0tqdh1/7KQ2ZQDwBivMITHiB3H6
6n9JkG75uoDbwjjgpABPnB3ExjQRuk1qS6JmCc+ym95eL4k0SCYx+DEsA/Ox
PrCPXYg6oGA9NmBi0UxjQGkTjkknPCGoZwAHsGxc7+oudZWEzaaFwQT0tIFf
HWixU1uBnvCeQiCcXfCxph4+otdyCYUE348bNBLuK4NNOLBjGm4cAEjTO8WZ
VlktCiR6z7gwM4RBvapsBmuqXJA7C5gID44f5BG2eW/y0mFD3vWnpEIgBHfF
7VUdqmVNCeB7htU6rzglizAW7eqrctIdEJDS/nYS5jHpkXAr4N+pk7mCgHs2
Ey2C+ZyLmmxeOreOdqY5myX39AjsweHRCSgb64TmXEdCYE6IxMJVRgjC+I67
2/MZsNrWxUkXi2OqNKkK2pZXOtqC7dga9mZhEW1zM9n9YduN8m6/IezYe/uL
DyxBfce+pKMZCahvepkGB+/75uQOHZXiArORW87e7cFyLdHHGmRtIzC5PpyZ
AdRv2zbG2TNsd2KgFfcsPerVabkFbT1TdsZRMqqvDAT3cnDRRjUaYDUeDuTA
RJhOBeV+anSIIOocZ3roYdxwpSa3AruJcIgsKLNHG4d7X/EkA3Pr4oTveldI
RYtwTvaMLZOy4fyJNKswoYfxCx17kKV3NqFmgUvJ3LgtExEUi+w4JUI3k7E4
qsS8tGqtuqyRftWZ4pv9Ll0qkUy1kv1McU5SKFH2N+bvp1GaYioDg2uxQtAi
7zqJDeBHCvBRe9TAF4dKtNAWNWPDkEBCvfzczIHP9yNp2y9uOcANJ0AdpH+p
ye4KPA8eA1LNgyzWCtjLE0DVxDJ6lBHibpqvM87Q+fzRGulovu4pGfMzbhxX
GbBgbQrOAfWxHFup4907icmJaj0D4AK6/tR+nOu8WFTlavHw0Ue4iePhzUWC
DeUkHECIQ5sYHz0/N8Xxrldm00yMAxjaUXJfR2k/x2724WDWyxO9pxsbzX9c
qdUgrFwcPieOD8vD0X1iYYWmyB6634uy7u+YVnT2nVt+ZandgAPy/moBs8BH
GHHNIV2/gtL4nKa+Xl37phMf3rQ5w9XALMVm7tr3AoO/r1xjhOEEDwiByRpP
NMbBQCCR3Wy9OolJiO8M1xuQC3anYiaP5Iyu03IQyHFA4akD+tgNYrj6S6hY
dCx3HGJL1Zr5yqmc24dycP5ZizkvcdaldL7cuzR0UMSXTxPdO8rZ7/LnSo4H
iVe6mX79oZ/GqmEdAF+5XDAVA60kIvqbpkIbe76I+ePwD5OANYh5qM5PF0fP
Fi4VcHZoPnR/jQY7ynPorcgulfpuv6YlhiHFvA5om+HS+2JMZBlUlIDBD6W1
LgZrHATOkXCi6Vwytizqc6K+lktAPNKF6Dzj89LABWXe7vTpRCLsnNX+OTux
/k/GVIoXs4DSonHOdn20Ly9DbD7zuMU8gSJb8ITFbr7+Puzd/Mfn5kvBRIdE
RN1uMCClxpjfQ9zv4CFbCFkiYOugh08jNJ/CO1sfVQB5QlWP8piwI5IeJMCN
8xzNytR+DOfY9OnTffwAkLJPMlFKhbpqibXFwLNrDX201rmT1sacbKX0tTj5
b56Y4vyQOXiXhlmg/qHiLHUqzjjl74Ztm+vgIBIBdAvoRPZpQaJrWPFufxSH
kTQrCkNz9Ld33EzkzsHNs0kYOjah8iCUrsQHRyYQ/W6UbDX+tgq1WMjTMRaf
miqc7GnfkjG4+f8DascgnzSmCP953KqMrpV2DqhbIhJBqMTySMOXl50rEGfT
WCpjLQ8qLPhdrrz6iA735bR3XovrXxg8y5hkSK7FFKjesLfNBGPaEm7L3b6T
Ca1Ogz7SzPTEOnJlUcYTESBwkvZUKBTA4U/NB96n3oc/YRCRB0Q9qvi1W0lK
4Y2Dw8+PAo24cFX9cclbwlnLvISJPTrlFbAjm3ZC6jOEzPS8L2a4zPhEWcHG
s59KirsBbk6Dd6sAQl2Idblz1D3/bo9a3GOA3OJ5DUzZeUJKfcL8An1J8zh9
+7shIs9oVqRNDhAGCdOAk55JIy1nUF4zQE122qzQsaB51ZnpLj610vua9jzn
PHdoeMZ+zdfR2KaCW4xphk8tvfXHdpEXJ5oy/Fo4b8FM3MXoyqc1wtBlhlOg
HhMNO/nmQrTvhONr54uB/PAu0S7ZzR9yZMm1IaoNLnZKzSz6qngn4C3+GgD0
mWpNk3KanLDRnzLNKT1LLnCiuYRAiXZ88DvZqPYWucXNlgHe1TIlxUz3ToSp
E7UF8Kxr2LBjKOv96LhnOlEF5FCKMS8Si3CY9TTUsNFxsXnedqbs26D7BDLH
Evr45YIG9g6Xkxie15kW533gRAtu6rKyG5hkzJKTjJYVB0z7r23/BmGHHPap
jtw7gGicsbV0Dkt54l+naXehNkY/f1o2bt86uZQChrltX655Tv5Xh/lL3Dvq
PCK5De8juuwWcFhR/mytbMEOhNLP2YQ9H8jRhsBlNTsQVnajwGa9KXcadrCQ
x4koXjUtiTZ0TbiGTJZ55C+uVpMQzPu2qf066wEv/7Qjthgb8NMQayxuLoTW
OPUM1r+4clgZSTbXnZC9rn5C+kWbtHuyVFWmHXugj2d6pDZ8MeBXEHcGKuJJ
UL1nBkAg2LvtYKFg7+BPbJhkSi9qXsDk4MogKxesYwpuU0/qXmTnT3zaUlsx
GxuZ0SLEVUM6u5edKlzRnZm8lEC3OgnwxeMzzyzyRIMVmiBq3Gwc2nUMDvns
RxmOQc0373Bd1AlsKIGFvCXFE6XddyaVjDK67hHKdrjrMWoZNI+V67ix1YtF
xkBAAtYsI5qPXvKx29LZDxCOBAskmIbqILzZS385IQTn27Gl1QtWJDA/wH1R
vi1AlQXJbb8TnM7kkr80tJWZctOswxH7Er+JlARn2futRKxSatLcneYsBLnz
osl1LAHdfb4sdaZkvEKr9gwSr24BvfcRVy/quhQf1obTebAVmxD2eaiUjIC9
9LmOi3uMoNYp6YgZ0I4UXKU91oTw8rdaB/JTNvphDbSOeYY/P9lQt1d87AIW
te2iRc2qLT6huc5QKTeIMbm/yHTUa8pkivr8IYSTGR6TylkthoBaInPgGzz0
TYVEvSKlg8drxQERM672NEF7Wjmm6+WANPfCNW2kxQPlyV5emZV24o52smti
WcgCv54ew9qF9EOPuKzd+0i0w/BwAFDxR/mxXmV1TYNxO1DfStUerL5IFdaY
+trHzpgYky+3eYGHIXyFa0Pg8RsmMz+8nf9zfk9IGrXvnfVtP0zaSr47tYd6
64Ae1hnd+lNXPnixSFWdXuOpPNf190Q6ghIExzedeLwVYJnmehIAfIk9jT5S
F8a2SoQCrZw3Ao2/JuAtlgeo3VpVu8omr7jQ5BivZITuOkNjVKUfRDWluVtR
XQbMBxpu9LRs0H5ttjz7OrhudF0zmgEXB7VaJaVRDt27bbLyyTzOsZisqfFD
hZVRz8XpMLSbUcRtQKjO8tDGADZyLBXNiOASARO9xIwIzH0L6Le0d6I06/A4
vCwS4VxPCfndbTXBF2qkbojNj7Wd5deBTYyS08yzty+doZKVV0o7pvyJQJCU
Ljzh5vZyCg0ynhWwf3eI8RDZMOctAysa4oQeC0lINmDjUjXdv8/dF6v9UoE+
2wHpxkiBjOQSTGlgp3fPWb4a7DmtCFqzGpoCFnQ2dEsh7MHNSpVeQaYeI0xG
Mj90KpHMaQvidKm1uBPJQe0FeF9LX4ipC8ztlmLdQNQdidrvquJzknqRLKZg
+kJrlXjMETIZQBUVa6IZxBYAYWFWdawLdMLlWv98w86s9Lddy0NaFVw5TKrZ
aOPCloZcEmwxIKx2GBsSd49Saj7hYpZ+t8obL4v9sC9ot+3UAvz7kLiafCeG
XNdS+XCjvlowPA5RE+ljVe8kzSCV4hAcTrkOqvPOyJxri7FS++CdIvhdAk7X
3rPQmGOSOImJNwQ1AP8SXpBxZrSfaeFONv62fP67oZqguMScRMfykEBW7pSx
0n6vH1gPmr1QPhwxuJGWtbWmzZF/iy19EmnSEemA4S6ZeeCamxsPDm3g1Yok
T9wbhYP6ztsfv/VY4TvCKO6u9uSag1RZFA4feNRWI5BTR2y4fI7ZqzFFNyX5
a+e70+lmGRthj9/NSVRuhkqxttzsYqg/ot/kiBfyO+LxlBSOLoIh3n/PF9ci
iyR1Mx0SAbJ4Bn70CIh9H97+149enlqN29S9j98FZpAwSzS7t+Em4jmUCqnY
vsp1JjIwX6C+1H1lJsVfrWKa1mxu5nFJcNoVz06ARZ6kyJUo0ghYaGMqv7wm
rpX65BufmwAnmWWaOrFfot0hOuzHUk255v4mP0vVKKP8CgUdKN/kCye8hz+j
egUSQWqW/nIK6jqUODcjuLn9tBNupKFd5nGO0ZltNgsX5rTd25oz7izfqbvX
pI8PE7RhMer7uDfcBDAXx75XhHbID1vv94sDQvUtWmlr1GaG97sg4C1hJqAE
ZKcw65FMrIN5TMz4JutOBp6m2v59cyZGItIM04/VLhS2t6jSfcNiSto5V4Jy
vnV84jA8SNdu8aCeLJYyzNd39Npso9JoG2BdOxGekCw6hdgATa2WEQr0mF6r
WC7p6bk3P18xShUnaNyiWhx1cfvMKyUXcU3oCEkdagPCgI5mi7aQaEKqaHvr
pBsmjPQEFF0DD76LkYE83PPHTVf0PlbAIMTM2giUKsmD4Y+CY604nmGIfTfI
mWy6dU50DK/d77BNml6yPgRA38T9LpDq+SoyLzhsQx+67gXUpw5UN291NArS
454z494fa2YGUeghcpFYRK+sBRRN7RnTC+cSD/Ik3AY5WAiQrAT/rdDSZeT+
HbW6kvmBf1jA/4getZcsn5Eud0xdV0Yao0g05hebTjBQZtOQpgNUPFX0AAwG
1FOeNcNTYgoCtPgquPHrelUguqu/mIPZNM11bgmYaMpyKmFw7k8fme8ln7BQ
nCA9VgWGGUv3G8X3pIj3xFexgQb3I5w4PXQSrbKGf3NRqtZJoLGzwWRigPap
FhQFfb/SkRjntIO//xs34uYk/FbEeVhg+7lyTc9g96yYnzECdB3cdbSAFziz
CCDLmBrs5A6aN/slvHKvhb0PZ3+lSv4bx8HP2O1Rr0X1QKEig7ta1L2g7tks
bd7eicSAvUVL8Tp5Z9IBU+doY8hjjabiNN4B4ZFkPqtIiMN70aiF/jh3bkts
DXAXfIaxyjLt1LWhCPBe4SgikSx4M4PMxOrG+kdVFLy4OAnCpeRmUFds01ME
5sGlZOr9pLYvGtarxUWFkdcLzOSRoTW5v07RvxJdhhf1ida34bS8GsAi89RY
fpYrB5T+U6FC6O0XxNiWoaFNFtOSphNxOY1Fh1KXp4+5gnq/0eFi3UXBsyzp
hzdR0LOnZPsC9k6ybyB+TmnJmBMNB/weVJTKyRgYAoCCsunxQ/+dJs8RxQzq
xPgRBykNqJQtBL2JF2fSkwLXdqw2Lmobt5sDMH3HWd2//YQF4nF+Giz1MEwd
691TUkPUYKyMWSaQNopRHMyQcWbyAxhYLJgW7U3xO24Z7239lHPt2mLd2yK2
W3JpRShn6Di4zI53HToGApuCZ4ztOrCpIVI5hq5xaVOwvfKRe67cC7L4Pter
UJFH7OXpCswb86CB/flszs4ZTgNk1LYFyKdlIFR3pw5NQQK7Qx/eJaBg6coo
DNjkxeXmjsclcIv1QIqon1wfXI/fFQPa2YW8zSWlX4l+txgPSnHcGlpAmNQA
aZdpne6am1dLrDFWb8S4lyVzqvpjUHscAJvBzZ3damFjfxRnmYtnvxZLiYd9
dYkb+zo7q0d7qnj1CqPkCXD36VbHQ/jJJMt2jceOE7lm1OMj3A00DiVuiUm8
CDF0n3vzziVBtZ9GeNLGoxp7E8pXI1n4LQ3gW6pSuiV2wNd+rhpIbRYe2ocH
uz6eLAsjfsBkcBe/7J+B5pYtHxZYIJkywJPncLn0+nPdG4FtMlMw1QHgxbLF
C7BgaR5jinvmb3hE/CvBt5SajMRNvq4/y/9JnYxsPuxpzfVAWGufDf9HzZQm
WajdmiKagWFz3YOQAZHlANnyF3isK+rhD7QzE5VnHhdrxlEbj2tc2zOhrv18
iGv/+2TBJNBtaHJAd7kngY/VMPSr+a6ZjWNVPJgTZGcNG7Kp0iDGIK580Ynm
yvPlvsResjdEMyQ5z5nFi0guqAGFljSCHQ7k/xxbL1jxL5lrOMld8B/VQtV8
02wmKtxReTy3gGymJKkTYDjieYenOxf+RXiFDrftnyuuUKSUSxzB6UfFbyXD
0OYDwnERT+/JRcSYbbaZ2FJls6Fqq3KS7QdbsYBjT+M2EOvnxqtkbkgsWuCv
6MvQ4i92nUI5mxKDrRXy4w2rWKjdnPwvGgouFCHB/NPGRLJrxJ0PrPTgJj9P
xBqR8UL3+6wYA9e1fRNO0IFyXy5Ljop8+E+MZblXPIX9binlbMyTmti+JrU4
qkWjlJOgj57VeXfQaCi8KA/aoPkv88TfV+QWG0fTX/itBUxuKWl8kJA/JZn4
63vD3wz8FkEei7nf9Eumvq88N4Ldwv/pGSetz3kXZCKy6drAxRDbDsriiF24
Bao7xxKn8NGJBGgrjxmJ7OaCYp+C6iesnVmf+4oLDBXdWg7fLzQHD/w0Uqzs
VC/hpV3RA+vgFhp7Y1bDk0iW4B9feO+OZDo8rWWHUqb1x+MVmUVekNO05BTN
JVBpGs6Z9NjslJVwnv8nscFKuZlpLKnc/FMSxwstAKbwldr2z20A8DC80s3l
+pXDI9UuxCLSmAf0Uiyo6aal33TX6qyIyVlEd38ITF9mOxuG7dC73mdAnb13
KaWlfH42oPuEaqhBufUYb35fAh3m3Ivf24wqe5QVqIqHJjIQ2K1L+4es83UL
daqpjgLfIGnbGqMI3JrkpOrGCbEGWzjXgrodLy6W4PS+XQxB0fEflKa/Udbx
PEG4JqLbIvnX02yNxRrHsE7kCeh3bhVxdFdRsbY3AG5CKMLaJIqEmPnqTcGI
j1H+DdxBlK4ZV1Ei+OGIKDgAV650KGbfmOCVPMwK9U3z2dtLexnol6rJs5i6
2l5EpnDuKWvtoU+jZa5G8Hnuiqr8AgWYNHLWI87FulUuGCF8BiqQWYvLJZxz
nLehSZPX4cnep9kVnoZxOpg1l/A6EL/qSQPj/guY93kLzcbzD725rDkyN18c
8PDDu+h7AlT57OmG2PEnzfXefdb0Ta4m9oxNx8p7IApZQ+A4UfL1vLLIRQdY
qonJwrZipIpuzgI/7840BPJJT4rAJGkNv1KTAW2ZFzxuH3NnuQLujGBNMwI6
QS3KcnWkYRhGe7XM7FPZkAI/mtWuUxnx0aWA/+MNnusLSk48BcJTg8EBJR6x
8EAvSghE64a8QQ8w5fWTqadAcmSr9kc1w2pM0D9tZ9Wqnljkq1tBMPT4GaCH
oPC+HRjwZUKTrlFejXlgVYFGBml8xDJbAuTo1j4SBGjnh2yvglxxqg1PFjCl
5gAc1S0Abvy7sYuJ+nVpguNZSoZsaNeS2bKqjF6OET4ootDxP8s/hJBZ7AsV
QBwZT7MTpTG9+JqZsYoRidpY1VGzzVt4aYSJYCWCxr2vVxkg6YXX6PH4yqsT
J74R0Zp2H+hKz2sRBD/O+a9LpVO3D5rkSbhYzEQpJSeeB7ff/kC6V2PzN/6S
ioUjD9whHq1dCBd8GwsX1p7DhzB2qHyMHIom5NJYwXGzy9egBUaOHxP7crXH
o/YJfDKb/ZeyVlGSMr5OamNau/B279lqN7JszACkq9emeXY6Gu7IgddWkXiJ
4xfFjHrkAXmegVE2em08rVxI2ImlJwdwkwMwgh/+KqroWRcKzRuln4qu9pAt
GE9eVIkYxBwvP+RAXSL27vKAEcYKVORLerfcFvBIgeivPfdYtiP+v8+fjY1W
HjsUvS2vBjzD8gM9lCh56PqMLHQsRU1sC/sWRP7EWI/tFIrim5sY+7Ojeyez
gTwhgReeCweVdiTAiZYAm5UVma8bwNavlV4cMUzWkcMwC0H1FrBRQDcAGy+w
SYZpoy8LYdL/pCUwL+mXxrLrCLZDPm6BwiWXg2zIva7SC47b0xxC7zqwGHyb
+4ci951k70dplsl1YMu0NVv//v3YzDjb85sn/RCsPFFdrqDPIgdX/7dWwsgA
JxcrEmC5KPil5wZpHI9/ZHsVifJc7TQ14DLQtyI6cTqmxe3IOKGi/zueGZ+A
GpFPsMCq2pQBRa9OxiTPA/OuiJ8lSSoYlmuMfo2TNPRROJ3v8yceMoerZWeP
NhqvI+J+PtMIMg9zR6cWjR1sfMlLiFpu1VErhP/W8zRz0rqe6rDbs9J6uKK7
y5fSTLMvrqnCANRKPlAQEqyQpT+MH0wlzQTNIVP8rBAoylFdXKcLeSoHOSjc
+i9sEqikuTYJq6L5VYAYO2unOr/yC9KwYqX/or++sCVgLoClmxis0nno/fyE
FCb2Veq8JqIVxylO4jt9L92rT7pqL3/jtE1Erj2i2kwsIJuKUXEn49lunJf8
mVGJ54XVPZPFP2Mf6B/35B/xQz1IEMzIq2k3Oh5Q/YWAtl+qUtIFAeCyd+xm
MHBVF6mb5GY9MbFBlU555wztmuHDkvlCZ1em0/CTWH48qmZ6HsC59x8Pwhca
J71Di5hHTiVBjUCKNS5v3Rlm7IgP90YTjXaWPTqFbljfVBFN+MZOxpmsnkiO
Mc2rE6iueEzH0pswGDcrhLxMGhFFoDAoMrK+fz/TGRDYBWrdcoUhM0ayPmcs
XwvHG7bgyxN1mnjthh+SK0zUg6iv15yiSdbl9vMSK3Q2tveshLOTV3/QXOMT
OznW2CWcQU+sH7g1HmkZQJL+X7LiXoX4XggwF8FL2mvqZSm390NdUx9bBzpF
U/Tzw4bW5ro6jfax/hiknwTWvbq21jW7NGZ487vQvd5UiDGIPwlglWHzx2FT
/LquOlDfKwpRfSoCTVo3rmOa6VWjOmjNKDrCyZH1rqvhkj5KpmMtkBOR0/A/
u0C+dJgwhDqEz6doGFSnaLw2RVc4XV+paYxqK419F+jG9qqyCO0MojpMOHG2
GQww8SdMfK/lud+Dbe+t0lfGxwVHV+/aV4ZYaXt2e6mOxGeBKyws4l7lkI+W
MwIWcODgAKzLf1keCLGtYswHn27W/65ut0R0P7ghLePaahrg40cTRRPnhAYP
pmbYqHh0q/LDfdN5xhvZ6RZXr+SNUecIcXpVNr1fxUbOKKwXvwzgEQRAZSGs
vAftqD1Km31XhNs7SL6NYKFIVSk8tEmBips/bYH1qUbFhiT/xjZYMrBW7qTW
7S487B/6WHRczYcpjvuU5ZFkNqz+WRKO5E05DMwMCsjy0ZeneDhCVITV/CXk
TFHO8IQS9C43HGcoFlJP6ux+b36O0TwjnGlOxF3IGHesV4F7YrDlcCfd7c3T
yZqlPvftiAFbRzVYIAM9/Jtt9ZKprDOjmI9qnwSYM7zmfvLLj5KRnLYXERbP
oRjlMOR5qMgA9l8TqRpx5tfS1U8vy7/MFAxQWK4JvxAR7i7GkHPtrw2hJqlG
HZ7s6bZp39oMyRqR0pjloomuJvWLm8a/sD5gNxr9jc8lmWsjzPb27h3VqOLk
e12NVHys96OPiydC8trqVcGCFlbgyLQL2T5hiI7iFotrcBBqgRksbMK/LQ/b
asepq7MH7nrRaRZLlkqq8Z4Cuwp/kb1zqYQ7DYnQ5jyPJu+PFkoYtUrROZyI
udb+VGphSYsCUP7UCd4vDyS+A/5dW1uV/DvnM6IBW1UwHzibi7loMTeFh8D8
x52Cy4UkLUqJlNzm8ULDmCeKCNazqh+sboE9fF5aHy/CG0WoysrHprHlvAFP
DYsxhSZri4lKJGuUuT6b50Hclvfpkch4GPQlViyUSgfieyPXc9k4VPibvXo7
a6CTiBEvxRfxbBm4dP3836ebFNG5syho3Un16bECv4hm98ejjC3IIPy7sQnd
HYhyl8CPH+JLrh8otGoGMBIbn8oVwl+hsJMSv7EFBgBTPUYnNiG218czvvL9
dqvG1A18sWpNkPV+5gyeuKRRbNTEvGNMXHpns7g2xfTcJEfjgNOwBLQU/gwH
5Wh9T9qrFzmawFcf7Mh2jTxvARV5S5qn7xTCh6QTuMPsOG7VJ0E5zYP9hP7O
oVU6EvuY+j+dM6FpK9+smwe492tMgFVNxSaHLcyJ/7ueiyL0fGyrDvrTcbQ3
yM/rQwWpvaYpXi5aEFOJT2yi8+kwecbU2Bv7cEChx2dhQzKYFPpGP+/JJyIu
RAvRY02HtkFvBbp1jFEEVzU8n/fuRbVPpAtNbCev4zgGQcSZ1FUYS1AHO/yx
SqSRTWoEk5SwtHDKcvAO3whC896CdbTW73lRc/DdK4Ll2qoUIk9o5vZMhzdu
ddsJYocuNetImoIq3xCD+wyJOSAv8UwYtF7GpUvyZq0eK/wBoM97e0Bb3V2P
uJNAoJtYEx+hHy30+huMnN3QKU3XP4KyH7hJDZEQ1q/nwyvHPSo0OKvb1VGe
HH+I5twwIcKUPRjMVAcE8OXh/Vn6OHnzYWIrNYrmVBKr63pP4OLjLRlvk7vz
w3YIxah4LrOOptBO7RnhZ9qXHawbSzJ3HxocNtg+g27xA9QKlh7gsgdaraJo
VPuoXRaX6H+x5wL3XTNyfweigQdpkpv/g3/Bk9NiNYqKQin4Iq1jq1fDq8Ye
ynf8sxYp5N0VmjaMD6pO0u0CdxeFl7BDMinZnvDTb344ZdZ0qd1o1AmeYkE+
Nt93FdI4+dMg51bJSbpImm0XhyBri2eKShybRP3sjnAD2EEACXGXMGGEhHnO
5dMwkWuWgn2QgsPx8nqUgIX+RRqp9JHj2b3wA8ncojhFdzNNfCUV+sLX9rk9
gYMoH/PT8tPBM1/tgF2M8hh238/e91okMGAhMpVZohtlQHS2/29tSn0Pz2N0
hcJG4dSBpmFMkGMLkaXI2I0bqQjxaeKhQenI9lxTpprPQIcF3t+6F1qLQneY
FgZLqq+k2C2Hij92nDIX0hVDfE4P/wohiN4KrleM2MWmT/jxUkGJdYIqGurh
Rxf5OtEr60bBOFUptOFTaqkddiLobqmURKKfjjoPPkFrB+DwqNiHjnc8MeXj
1MSoT5jX2/Q8WnRrXXbmb4YSYbzEcvwi8Rq2PGR+VjVaYTXDi5yrcVvj+/Fo
H0uvabt6n+sOxV6eRzN7zJNLT0t8u9TEaolgs59ULwlAERq5zxFAl1kfoWJT
NS40vMI5LD7HUkOEvP6JDa/yi89OG5tG6OV4kMmEzAlDm3WAFdZoo8cbsCwW
q3rzCSznB4PG3S/d7P0aPRyzHcQyQ505Fe3+/bnt2/+D6zAZOSw4zAQnhi1g
a4lvLYlQ71mQ7vC0FpyygY9lkNkPKlU20cGtuYsF6QWHXHn5SsjCIZrl2Clq
4FqX8bXLX6GNzW+x5hBETViAdwYyy+XyYN11SjCpXh/QLkG5ne73WpF0lpUe
eIcmC7bqVjt0diTbjsCQ2udstvxOYOocWiL4Sl4aNQHwlgxJzhA2Hj5VVApo
WF+mlx2Qih6Xci7conL9hjGlhXEx+a4BP+wCJwzSYVdbJHZVOBoOeJM4U2qK
GsaxNcqn9CC9DCT9Fs6Dwbp4lopWKQKz/Zy+3qN120j+j2SzMiqvlA15G1Ye
urLKP7DaxFzT5SDIGXJnHdLr8tc8jPZesw4YGkz/HqYOIMBo7O8fcOfYk2G4
xXYMxh20SaWWxbl9uPhItsieibpgb4IGU7g1ICmXgQe+RO6iSzgtf5bh6ilQ
mKGoYVWuux4AkCAQ1wCyRt78vvGxZ4t8C6p+LDMoO0FLtLrZxJxORBMn1B9K
grOcONbWQK+fIzXDxkLkoH6qNoQSI6Xuodn5AhfXtx3xj3eoBiQf1/J1PduK
OV6FueFwM0I5QQnpTaFbdbn1lU97u2k7YP9SnOgsVmVPOOj/LYPgpdFsLrTe
AnuNqWw/MnAjW6HEGbDppIejnaM0wkJIrJAl9bGqDhkczHSCLCBz31pYQcTw
85MYfWf42pfpXZPJL0TDMTO/Rk/vnQd66yN4VPBA5CSH5Me5gPiN6h8rs2+3
SvsTcWmPSgCad3tVUfi2eOWItg5E2SHlDCmXLUlrrLJ8IZ3OmOuoCAcCQgTR
XquyGn6mMlSzMzDOfmoCtCnCpqeztArFnbPWIpewnhKI6MLS9w7mpeIWAMqC
EPfC3JqjvMSMW75cS4zOYyIQwt7sbXAmYztElRg/hFJJp9hAkHQY/aQY8802
JRsyRk2LIOChQTbx9oUsvnKbscBHVMT1QCHyAVK7TtDfvp65C3F+7kEYqphk
yCUwd/NgtTQgti547Og5ORJwxf6gTCIZGCEHsKpO1BCOGRyXHwN/9VxDAJib
7MSi4LCG631X7GNTnSc5M3tF/FAltdCCKkPPlxiyobzoV7o9I/HEJlhAVD+P
xCQn92UjMHmxzD6UWcHBYAFbpEwGuWCaSfR2N9UqXLFBjReztd9vtdoCOoSx
jY06riSyik9bl8kCdqYSZXUEKOdLTs3tLC1Tc7Ea1ZgYGoBUO5jJ0EHBCaln
xIeEecMOmR76VDBuw6cG0O7BMU1ZSFx2TeF2FZZqM6+/vLcWzOhyIbDi72Kl
PUj0sHIpSLDGtkPkalOs2rgDoz1Scdz9rInZmR/w7w6sqOkVsUNKI3zE+NTf
IW6vk1U7N/vayL/0mP6pJMRrxZvlz9PdY3kj64E1pDfdFOpLyg+Q/LB3LL96
PSJyEZDZC8bFZ9C72I1JG6ptF5b9szIKrkKfJMtlS6Y4ZUtYKxeeKAxgBoKI
PyU55ZwWsdmKXLOpObG5T+NdPLsmnMZvX+cyueui9DLYUncmuA86ZM34ayVq
3XAKtUL6q+shhVkzd328hzn+lTOT0T7JUmDZp8Mz3uwIaxnHxj53ahyxAOfO
Sws3kXjyZ2XgGFIYUFX/EAfR3iaMmNizsQaxo7R/DzPOR1rtsC30rJ/dopT/
FQBWql47Ktav0j/jqiqoOFksSH3gW/cATq/8d1Gfda1MWKzzd/waDzkNufMo
qNcYFVxsaLjYt+IH6Qx5IS5dvaryBmIT8J7oT7eXvvBMuBzJsJDIIj8afnRK
AA5XXVzMjkhlC9ecd7s7NiMuzKObNF32aFSyvqvXzaws55HRDOLdpfGNqpqo
KGrCpj5wOoBOuREgR1GrhLjBsH00vzseaSQvHfaLICvoTRJQeFkl0Jbk0uyL
rptaoooqnFQ/tG28XgCLwzy1swVq5MAzSmzpp7KiG8ZoUgSHKNqh8Thm0grR
oSblJFeOi8Z6al6+w82T18H2d4fmzecHKV6ZjF4590StowI/T0Noem8hz1fS
T4CFzUBk8mHvvSK0gdfXwlDmfSVkqqpc10Nwzalw63ljIJFREM0lKFpapG8d
Rpnr94BhqHxqCfjDEGc2wLJj5CFCxmeU+yPH9PEethGb5cBjcZSfsrQ4mzx2
JC4byU08A4PK280xEhFLcQdY2ETBKCJ2ev/QY+FKyGXJi3DaDljLiKiAZwrt
gurf38K7Z7V2NjTO43Hev+uW5oCyM8JzW0Qm3DLj9oQMsCloVmbb6jfYf6Oj
Um8+pEar3vnCTcjaYixhT2hLMUrW7smPJHZE3QQV2k1QGhv/Kbf9Eynv9x+z
OTLm+2hefuG6H9GW1mJTBu47dTar41MnwwFqsxjVzqVNu/oZzXB/1Emf66Dk
RcEj+F8jiq/Msgs6Klc1bKRwcjz8l3NywYsTVaR42Vw3m/XAHTEkljq2S+GN
ksfGIvUwlcAY1osvL+0EOAZUXKszxT6RPTSYuTVEyaQePRRxKerHtbZi7Dqm
3CAM0fgnqrZGOxFctWn1oQ4MyNNRCm8+dGOhd9sfQ5IN4ZYT6+WnaikqDsV5
2sl0IjXT7DfoSaduLjYvqR0PC8v3OesKEw09K5bTk3USHhAoCxt+9zRwW1U/
y59pb5BSKm9NUWJEk5VCxtmKs3y6dWfuinnPHqkSd660yyliI9IYGClIZM5B
dWuYsTf/CqP1POQn46otaAdC+NoQr6w1iqFOcorJ2yzJJUuZuisRIqxKD5kj
s+Bp9gbqt8gs85xrkOXTcFDfuczrOy/tqLykyn4G7Ww5PJ1RfWEKOvM5NTDT
Y7ZXduV4HL1VLpjvONb9yU892M7451NDZuSBiwVZML57a00m1HYaPu2mlbOc
YOvXyEJEpsjrkb8o7W+DyIO2Jy7BtARR6N2nwGBZNHKK/G443sAbNQc+rozi
LjIg3HTh/sDxe+J7PgeVkF1b3fOCiTZg0Ba0QFvWwGwvUhvDSJU8B21UVW6F
6Svk2UQiIDDnEQFeNAvcqfXfp+zKU5Oe6uF08XMOPXaqJtYi212SsNP48UnX
LlSG6VirFUzPDHaUVT8TYM5oteOscfEiqpnNEovcB9fY86BiQwIYI/ny3eyB
TFUhdNSfhA8kGZKoKFgF63XoiKQv4t3+7MHLLch0RPUFQYQkhI0w6ID5Im/X
G1UyhcIgu+7VOSCczf2CbMnbCyNdKTc09WGFGIhSjjdEBH1fgjT1ciQdZnSV
o1o3Y3qfRiklVxc1G3OYe0qjDplN/+o+3PBzYwBzEVRsyiaHO/QB8N0dRDs7
D6oPFZp8o36uWfiCG/RzYz5tY+t2IUxgXof/4CNS73VqUsglxfF9Wmy4FQA/
0+1RTdiLbtJNHQTtkh7i4yLFP/l1/TE2xmcQfYhClwrdlL+dqoC/JaBk36OL
9FoxdekbVJyDzMKa8V95jBw20Z6cZo9/G+Q4jKjqsvgo0X/gUAMycpLRDpun
D6cso2pB5LzRr9RRWPPZ1rNFV9Qn4f6zfI7KfZ4dqTjJhgeAOcIBWyDbisZ9
xbL+kTb1oNlRHN3+8r019IGX199e4TRWhKhLm6ZLefbqgKYYDQPDaGLMGn1d
PTfjdA4WqFzD+KS9Lv/aWOrABfhSmRF4WoqjBpUGRxI6b+deNWL7Ed7ibSOo
CDZ2peHh9lmtP91cpaZYar4xcZihUVBljLO1Hh1OlQCxBGP8Qh/KtevPTLLc
PgetXrhermzjWq88kPoqysyFtpETogPv1kS+LsX/4kqzoDwn5oJsBtJkpTlG
/RHQKjitbiOEZTKIqvfpwe0gA1E+jTXis9cBpA3XXmhK00Fx8v9NDt9Oll4x
aB5rbJbd9AAIhUhxSSYJvNjLvzaA8g7qKcGw89/mOkK47syXN9v+t6uJwIJJ
lDlr7KcZgxYhRT+HGvTSOtTdMg+ykTwG5yc28nu4mcLS4MBcSjwwv39lRC3s
lxAhUidP+F8hrUNJbn2ob9F0qB4gGpDBUZB/GMzyXAUoZueAOMkjwR3/48Jb
NMpuVFle9kLDehbbQz9FKVk6e/znEOGIcABG9niljDt26kiWCngW9VClRfEF
fqJ3UwIvienlkO5y21tzjl+GzS0ZIVG8g5uuNpK2biC/F5tJzCx0F6M8JPo2
p86GRHrQsrH5hMjSzlT3yY6jaTXix8tn3G/QaLi9e4e3PdwxCb5/GbSwrcaE
OeVGL2LU0P+lEwJ9nJsyBKYJ+2fPUC+sOwRRESYF4+0cd1SejCVibmyu+l2r
8QGqzifGYSfAVpD4bJQjo4NEIre7dObaXT63Mt511r+GsRuzXWjCMh4Sx7yF
ITH8sIKgv4td8RTOkdmhfRm8YTqY2WCW7mQCOe2R8kw7QvvdqWcNKUgZfLdv
IkhX2uongYl73Ciu2EDCoJCzQG/dKG3b0gbPpIA9qXH5Sqo++AQn1y++JcHz
UurwtDTkNZacrCykvNaHkNyuJoW07kRpdA0czysLB1S89cbx/gVqZrXWVNeD
fD6oC0m7EjCtNBYe1FQwzKBOUcqG5ENZmJ8Mvem2JYGiBZSB2XI0syDuIZ4r
hIbWPGfZga0qDXub2sy+PB9/dtyv9OCHFvSjbFL0gdU9CU2JvPjtUj2o8WKO
MC9W47IqujkwLC2Zzy8sExNxs8U63pO0Jh2B5XygBsLM2BqjCoI/vcTNGl5O
Izd5NHCHDFis6rKS/UFe15TTfwRJKSjcPJDv5UcLNpVpRl5eqKc/uM4lHITW
M8qTLM6b+Mbt4A7pk+4eaNq0iucCjuEH95uG17fN0VQ+2dXVcZblhDc+XU1N
pJGlwZ7pfLfu+NFa7ICMYNlReTlRqoM9UHa/s73qhW0VjkV1t/zZV1NZBHju
NpqiuIuVCMbCUhissLrghcrVb7I0Y/67yYj4DXfl9mFR1VdvCoy4rUELf9Dm
tVRNXrSgex2vfxfwMlufwHizprpMRorpOjuB6ad9Xwv9Fb2licfvVUANsXc9
EJk+WdE9OTy3WZEnGODvRqZ1XcS1IiYMZ9oJDYmzBCjj0sGrHDCi+1sMeDaA
dWzT/e3sFNhMg1+okgVWU8rx+LDcDS0mraonXi11Y0lqc1qaXrRj+0PDV+h2
kX9dcSqmN4SnUhceZfiDhYvgQVYFDAPEQagbbnCm1Hi8Smy3OYVgGwc6uHp5
Clw6nRH/nHkv50zoQeWsJLS7jLENQXzHLRtKdd6ducvVI4StDMUKkK+NgTnx
4twWV69TQ1/ABgPlp3ifGGPkKBHhEKGzDV2WfryHyM2gBRfS7UDzPkRey7k8
buA3keO2mIWVtRCwmYDSMzP74F1WKPYN2acxwUkwC70rrxoJScwrH1iVgjnA
fP7EP7vXp71G2fgvMeu+gT45QrbotO5Lqf0fL9SO0e2onxLHJ5dXZ6612PId
a4d87oGA83QC31RDrQCWEKa2wb7djnprKkpOaHvfQ1uOrO7FpFD+lhjiZ3nX
xuOCBc4E+GVAY0hYe898EuB5eFvkxZgWVQC1LsSNLGXCcmdrmhIRLkrPJ5bX
bFyfA0UQ9Lsny4dvDI0SiUYuGZYdO3NSNHovPoIEkxQTWbYmghhwQJV4mIjC
9ZNYu4b6xE40QZ4ZB0eHGvVe1V6DNW+5eQt77KYqm5D2jkpZb+5p7UXvljE8
PQeSCNR1ouK/3FYxwAfftV/Gx4D0DUllpSRz7PZ4J4st2Ie1wAvrSumz59YO
ofZ9cTmkQS13v+Sn3ofz+o4OdvmrSudpPRxYgT15oS3rZ3WxqqSMeq8haMdg
rgfD3ufDy/FR0m5q3oD8wHdSE8f9StE7GvLF/10V+bytTIr8h6D2m3DcB6P5
J2lZj0Wwa4d8AMwD1cfuSqRpoKSdd1fb25d5Kk9e/87FacHSM/fL2/y07QUH
LpYglTUfoJ0vAIkOZiU4hs0g/53MwuuMiJu8LIvksXqb+D3OjrVRA1dMVUR3
9ahsjAtEm8dP8pJIB2vqPjHBvqhFk/8l9WOwZPauIewCePudSawNM91IFw+p
DcEOPbII8Nj6CFF4DSqFEnPGwj1ZsUN1YKPW2nQwP1Z9GlcMS1s0LhHVk6lQ
CYxWDxeXUAjmbKd2j8V6ohoN7pCoXLyh+Vm/uGA3bGXwp4rJ1fI/gxzUWey1
iQrBsiOi36lV4yzm4Xc6b7V6vPeNtTMzAkE0Y0QhTWfgru108QvRVDosadjT
AJfTjwXiMrNyIefNMbHtBtmUJ9jwdJlAf8kHpfFabp0U1VfmkRUPGSy95Ysg
2kuScrw50CYX40qWWIbLj+wmbjubxyHfLXRSTPvprnFEnkayvdu7LPkF0Zdu
QZ5HAH+XE15yRNSZBVZXv+SSZSjvLF9FuVw5BTqynM4fo4Rbu2nkrjTzTpti
bUGWVWF6Xm1hYnfXchhjv1iGM2UrdPF/zSlZoVt1Rg42jpig6s3JPEwMkBg+
/x5N5csDOdi225Jqr5h+tdJStAIqk3O0PvEhiBVJV7dfPonJxNjcXBy6qY4C
VsYbTOOftu9MsqjlwdXVqkPvG8f6KNwfwpHljPW2Q/tUThvWSAuLilf/l14V
B0xuTZ5PByW7FZEwumc6dkYKlznKhHZmC9pQcUQWQKDlSpgtSGfMIotxiYjq
cTyoYLLYj5aqh/CGIpHI+8CyTu4wY9SPj3JUKvZk9p3lkJINhF/2RZmSPNbD
Eq523uJ9HYJH6Bb0e1lKWvS5TrLQgWA6VVqIGXhj+cz6ub9dZtYatow6FmKI
KSo2MI6LNhdEWJRZxF7vGxueiH7QbGR6qtfekYC671aokjbFqN5NnWVs5MhQ
ocWQQNINdtaiVUs7seJuiZERGbThMr5X/JoqKeJVenzlhXPhlANUSKPBfnDS
hRQ9Dv/kfG+AXyQWOKeyW8JHHEfLXLCWLXScO4v69lzNtop+urzMSYiQk6f0
T28Yj36eAGJ7hPMAQwdF09f4SBBNe0RYezATnI+01Kn9OQgJ5X/3L5+NoaIf
P4ANpyLrZi5MadwtFncO/JZDBxPLgHcpoFVvaG0nI85NGAL2hp3CQh4GVcI0
VvBBzLayKye5K4K42/4i8zMj149dAYjY3KppFgMCmp8AWhv4LhcsJztB+1BH
OG9+xqtiWNWp/3HskAyiu8g1xF3CaNfjcVkee64H0loZy9dhPTlKAvreaZt7
izGxHOfdbMZ2iEQMKnwLr5ElOY+cn2BlcM6eAkUrFSlJLWOmHtMfB4dZhjLO
MuVpEI5Rrd0J8040UEBlJZlrTHA8wfhRcXw7pw39ROPOOLbFCVOG/vuuMcTl
p9b8W8oympUomntS9i2OMreWh9hgdMkW+pR8jopDE5Ar2xW9wXtdcJ3nPq/0
tpEaJN8nanSX3opZsUJXqLlDPJvvB1Ge/x83i0yiKb7ls4zS72irMkVjS4DF
ks+OHgVEAwN0ilQPqx++yJPcanhpziTDn/odluhwcQDnD1hQrFBIfnE0MF6m
hSMllFeYoniJZQJNvwZGHZQHqt73ylTgTUoykYBoQzqN99Zcu2BXchmGb+bk
PsY49SdkHsiecdbsDGyZ0cm+MTcCnvEKcz6AGn06yc29TIneruX200lfBLNX
WG/B4J7tcekSAPpCn+zovDML/pXlqf2/epUIIDCacfmSnCis0ayIXsMqKZas
wH9/1UQDrljJgfr8fZJVkGKzM6vf0clCzhyVesFusXyWu0+j87RfCmu96FWl
zu+bDnlJNbdBa8dV3vgRGBYoG+FRiklWU6QswG8Dha3NExla2buzckyz9HjN
oU5l+igzCIn4GxwJPdvLEcg/mCDpOlqcoCUSSrcdTFHvqzkyBMAo1qHvR4ts
Skg4WF2gUq0Fs91MEcnYV1Z/SQ3VA1fiqoFC5aWtQ5jUY3ctBQ5dEUDiJovR
4xNfBs9RLnAaFXemn9yC/co2UK/uwQA/r63yPF6ywDi2Q62toG2ikT8NmbMl
PXws8aZn3ZCaQ0t9I/CdKZhJ/KGz8mLW4jC893xln/z+eQWyZET8I/PWSFy2
yOC2wjiQaC9EtknK/SOhJeB19dT5exmYOFWBlWwiL2ksya98A5uyts3s/NmW
iaD3+bl4hJo7h9Gpiagufbaj1WVo7ujhWVRc0YcJlDafD5Q1thTnUUX9sMOV
p/F4kfP8Tye/t0O3qF1y007cToKeYpow7Vf7vGBEEn9m8qmPEaDGtX8l7UxW
lGCjOqmXSUjQ8VJFJFpuk3YTeNDXmuxcHdS9/vPsIjCmJIGkoNyXPApbpo18
O15m2yPZiWgkDUdFeoOhZpFblsDPggDRKhPCSyBHRstFwUjXYunVFbXajW5i
OzxXo7M09+snZflpHy6FE293JJZ8S5/JwgaKromJlqHxx4pib/p59g0mHEbH
y3nrl1KD0BuYDPTw/ysl7UQbRwOowzVSPvP2In/qfuCZH7zDVRrJwqfdL0YA
DTk/KAaClEpJ7jXyPIvN/GY3mfXb45VvPf/HbaGcUHMK11soPOZUJJ5dDDR6
jPVVGJFz0h7K4jh0evrhVRXmAXRr1Z1e6h1xMjEpYxWadyI19hYuz8LlIrBC
a0ACcsjq2n/y84E2MVLAbNq7hNAEE9Sx9fknujmmynmVz0Fa0l5SFobc0O2m
kdi8JC3AVAYQ5XpmgiY857AA90mJ7Ru2381GvOLtUeAhXl0s181jSg+Ef9Ze
PDbrwwrU4P9ns2wVSGfhoythVSRdgy4Jf7lNr2XtrK4HUP15ZDOKg4tPEx5r
+AwSChla0tcc9ER7B+6bcENZEeuXt/NLyreWz2rP0HbTW0JBaB+vSN+bJsJ2
g7cyTkaYeiiANBYs1YjqUnSvDyhf+Nm16LyPG1s5KuyhJyGvZaAlwwtUf5Ib
D3ahzu+PXwG5JeuELB6REUyV0d0kZqjiMLACOjBAXtiuHZBf+jnaxx9mllm0
Jb8cQpdjpuAdGGDe7O7Z83mLJAB6EoE+2qfCB+o0sj4wpAsVDqBdL6GtWLfz
Ne9SoB5b4obd0KX/Lt80B6a9Vq9FTOA7P0ntBFM6/vSkLWwFfhaseDwq84ej
DOLendc3rNeCVbZbyYY4lO6DHJ2ycM/fTiw9enHPBphhpSvw2EZzp1Yv0VRh
kglRd5CCuvLK6SEMueR32fQyEDNPs130hMIlzZd6NjJFjsNxJ/qXnewOQ/N8
JnkrruG9fEBVcqet5L+hY47Lv0IkXxkLL9TQ2smBDJ4gHe7fkgUI0AKcKeG/
FY0xjRG6yDiifNNaK8XXoVyJPDl7Yd4txg5C2i7lmP/O7LoByq9r/TmXllw2
sgzZ58Lvc4X0t7pru7NN9pbvI0zGibvGB4eIEZmYiueTk0fKw/w0fLTNo0UF
LuTAjsSUGj9YRWs2D54qo3Yr+H7y2X4ZBlZzpAzvncAU6hI3Drj/5er6uaTz
NZJNE92SjO9+5bE16OIRKGL8+KuSx7gQexd9G6HRA0pjpR+rsfF0EHbOvjlU
/el1TWAffmmxkX/ajBAcWe8hOvm9aKdR/HhNdIYSXdUvzDHA48yEHCBiPETY
qLnFVQEl1aLZqUFVAUBRxeyfOt91kNFRlGTZb9JCG3n1tQ8/WhOC3B2obQU3
QhcJtcq1eVTkM4fgiQbKHnqKbHTZNZC+kuScYV9UU4+WOtaWrCQTue/Kr4z5
x6GAr+VyetAirGN+fpCFLnwln6LM6hO2pdUypLF2tGL+m19znd2rhlQ4vP31
u3U9xqQO6h2ARtwLU0rViVx5Sg769VB7MGfdODxZEcJshpYz4nLa1Q6vTEZq
GhtFpSy/WXmt9PvcfdCT9FMb++dekLycHpH536qi10TE8g7GypWojAZwCrqK
i6OlYI1pe6p/dl10Rr6HyxBYCfdqtgmt/1AyLh8CF187zOeiKqMv6tDbK3xP
aOwgloSewtvVirQFC7BeBU2uTrq06GdHuilnZT3dEvLbotL90rKyQ2W+Bha8
5ZlFxlBYs25977J7ssPnH0iNBardAojp0NZ1BzjIaMfYkTzwN3IBdmA+CP7P
JtNzkGI14qbyNFWRw2nETCXsVKzG3uxld2Wd44rO7zL+7aB3rBDBinYI4pqg
Mj8yhL3osyjCxnpUyNv7NHQ2brn10fzBCe6UuWxjY2Ae+U1j+8+ghrlOe1IL
f+iEWyGac26gddcFwNBuWLX0qdHseg7rF+tOFSK/1nhaJOjDtnZWb+zymAD0
RxGuWppgAevSe6p7nenpLHCHTCjGzuwQwZvDD0PzloysAMCa+PA+DyUaQX71
RwCkR3ITfJqyAhY9jvAPtCcnijvMR1SjJlBLGDoGAYqWZ1AB1bN79zvuCIAN
LqrvIjOvxORfPmyQRtVN/kuT/ZOJL201Irdp1t5u14kMwUkDHLt5VgxsAa00
9WosysbeTpcKTe627cnFUUkFYEADizZahXHj/JO6KfuxPNPGPGIO0BZ/9J5D
kMJuGSeDqYgi5E3KoDDjgD27tkNrDy5o5hTwsxAADQFikRSqLoWKXHWUjuCd
7i2eK9WS86FYz2JB502rsDcLuN7lRZ0+wJ8/s428B6rSG0QLuk+GPnEx8UAZ
cGCN6e9znQoCrjbybwG8MrPLCo65Z3jP7NIC7f8wg7DtR10nU63C5cONgWvG
J56lQmIVkZxtRZW+xwNkj0RaUFMvzZ2RLwqxxV/HilgatK/Tf5IX6Z+qsBTt
57UQphJs8SCefRj/HlHbFvS24bP21evCEHuhVoOnUIaKSMxocK1dRywi6GXX
FcJWpqnYwMOLNLKFUiMkXi8VQT1ZDA4ekA35wxNEibYEkeFXWa2XaQnFD+5F
/lTIs40utDOHSGEBT8TLGMPkFNdES9RkhJni6UU1bHDoizwTCo6+lLAcsIBy
GzKT1aHYg6G70Z8zRFYbwNZ85Hg+J7AgyEKV+syZjg81h9WgQOw/0MPoYBit
Z7SbX9UmSqRycgMKcJWRLZGHKJezEGCDWSpoz9jUn0nfnLMQNcl086+ePpim
uRi8BoDd+t//wT7jZ473Mr2TGNMz2xpXSsmMifwdlczsrj0S8hGdHBiYoTxI
sKbHzH/Y2+oOOfknM6LFR6mQsq23HQ7VGI43Lh8B+mfn2iqzdIi9b1R8zl7s
1ush7FGkp3ukZfSWF+c1OBZwJ3GDxaQs0sGQmwP+zu7s8dBBAhH0R8AGxEae
p0lUNaDPk8ih7y5Xi+68+xrwUh23VBJDJyA+w+Mb8eRR57Fma+4KruqCUfSe
qqcoMj3DfRbcoN+5O7Y8gZJvoqWWLH6QYPL5kxXchGhDZSSYM02tvk7Lhjys
Tl+oG8lKBp4GrvugVtHgCus4qciSfhyqa4j3oN0hLGBXORUeRnLPluNHrSXx
iyq/I4rI/XFYwWEmWVw8J1fzmjYTaSZHAhsACtNKpQptgP+XKXFyocWyaGGo
6rc84WJQtWBc2gZ1poWw8lkDk1HEZZajl/3bAfNrPQsTSVZFXD9uLiWJemfV
lFGzuUBoX8OBmF8rsZE2kgV1njqeU2DEGlTM2dK9bxxw/waBV4VTiIdN+WYV
fJTQRZLeEwf3YJqDFR8KmRQJZ5myeKcvej8+yU3HSH2j5QxegHaVTTwbnZKm
/loPh3WZqzRcyyY4q3cHWXp6wm5aYHhB89l6ACF+KMpCmnWsEZ7ScoPWt+Nc
iphKKSM/DodBloAiUqFrGJketb+CFwLfn/77PFAo9bm33W5t7PC91SSI14Zj
1KQADYEG+lPL/TWbur/DqqXF7RUn2VaOqLOOEqOOD+u2AWjjVUSChYrpRKVC
TZ9CGAbYkFR39DNnzITFdbjvd9sjMPjXjEhL3IbaMld8UOut6Lp5A4ewXLxg
pJA2ylG4Hj71pofUO7NHgjKZGJKukWvN2BIl4v0WHvFaojEK3hOFR/xR84lK
FVDZ8mXmaL49EI0Q5D3dPqUsw52cxR6r9NT9LFN1o0KcZdVOYK0Buna/2pkF
DT7cE4HgM2pHkKgUsbjko5r0n99ArnBzYb8ZYKgDS7wx7VombhZ9zowvXv/Q
jRZJli5WhKBmC+nC3GVS21/11ZOLdTWTmBZr7URySdxP2beFHBy+SdQ/YuZs
eqgkb87OnoSmVpDj9W0zzAd2X+75wy7TYzfzQmM44FjqGYIaRM3AKCMhx/Mb
rWRGO/k7kf0JH8B5mBUolB+JYgZksFBrWqQZgLOs4VFmW5XchEqIMGDMtnjk
YMcEmaiFGVywrU8C8FmeWL3yY8Vj/c/ro5tZd7cdvN6yKqOoLBJgrI1ingUh
h05uuM9rhO6BC/gs/oRtSrULwliEzJKpQ/Z1zOsavf/tNS9jqY+7z8ihJycB
i8lHyG22Xed4F/h1c17gOzMfPxuOOkBBp5ukC/DHo7uTyq/lby4ZOQegnWI8
Ce0hGzGdEYFCN1CGD1NlQVFL/fbfAvqITl7IMrbIkedeLdiAOwZ0nx9TtQMe
bjWM7Fy651hXTMOIpiMbVokJ5TvA6DFUv1UMZUUt3j1Ble+E6yXNOxsuchYI
GmLgFxUJNTlaETg1WpBGAq0kHhQD76DVf0OQbC21XDXcKX9zzFMmF5gYuc9B
JwlaecvpO807Yo3OEOoA102+asc3+cxL+PVlYg20UvW0qBVOODU2YEH2IDeT
TWkBxylvNY8SqwS0wQb4Jmh7+Ngw359vOQ3GVEhoNNLcYpma+HNyx7lVkLqN
fyPCuWVhram5LJbYq5mm3+lyacAlflZLSqAnghdhNDzL5p9bGkH+V7THEXno
QLCeTT6mBtdGwVGW6kO6he01peAcOeOzHOaBC3iUf1eZOwuHy6ypaQb8JixX
917FR5RoVDxqlJrwQhfeEk69msWDPssyp9FAQLigPov7ijhCXOlbDgcZsiH1
cQtXlGmry6C4pW6HwHQmTCjfi9CPJb3eUXtHy1UpC/JpY7nlD6Hk9Pb8gyXf
/vLCgAVSSN/2s9fLNIRYgOK8kQ0N3Z70FhTekVPpwUJjvnyUnD5qZ72+O9LO
CHC4MPHLqwEaoLPWBzb9Y6O6fUkMHmAc4KkfoJRseknzhxIGx9OcYks6Z6Wd
ngKvbMkuH9J7chsI/LuBsoIeCJ/OPDY6P4FJGZJOpeqE1aln6WpYUKVj9hRL
wt04+M9WM6PtxOkCZ++VRI8eBiWDIDFFZuknFY3ogGuBWphbsfI1LSjSToXu
BbRvdGivKjLyJAIYwll2VJGvDhGtPDiVmgNd37uUCJtrDf4c+ZF/R/20iK8y
mzxRj4VBZV8+iAxxQBzJMT8PL4ErYLmp5HN5+BK0/5FexBvqezMsWYWXDLJB
RCwqETNUvoVbLCVZKXPHpruqNyidj23n13n/9A2jjL8TUEX1P/dm8ocgTDDB
w8O8h/4O0gTGMemIBN/JPtA9owGlDTF0zXKawszowOYNu4h2xNU/OTs58OV2
eUgnmEMYeBr2K4toW1oDM7GxpcDZ41QlLyeRFfDL8gklglP9/gkM6s7CBkSx
7V28m/kQHUARmZOjcjvkMrEv0svwBN8K9lgRdWfFpJhlJ2aRQAvgx7woNxiL
XifGQ2SxZkKWtBj1SDPm2QKb66BH9g6LzvQzgKOLFMOA01ef/W3aAj3IiWDP
4hBwr2s5z/mKqEF8nQVAM/cW9JneieQmNrzCk34XDpfMwUAUxdPA2iYkLlYx
tO0g1b9hD/dyWRoyu7mB/jlqPrn2vk1QIA1t+cLAzLmDsiZMQBUqgMnZwvkF
bX5NJtGhJIeYyn9TOnIBOKpBR8/pdd65l0vdKMpMEhklcCDCSXs/au2porM8
J9qmASiM/Hhxrh8x7gVNmJciS1hfXEg+Ee+IXbB/bFJ5mscrjfGdfCE4CSDD
2Cs6A9PT1jpFtadG+b6rlo9O1oEJOwqxxWdGKgQVQ0RVogc/e8IXSIH5QJ2u
VbDxLTvlLIJDONxApy5k0ybAkJBLekiJDxUdFdwkAQGHiSBiaDQ8BCFMK+f7
K2Fq0Iwl3N1kBW/u4XHaYLo6M+StQb7KUYtL34r/a8iPEh4fpw7Q3ZXQycUZ
vUPdVNE/HtrN7BvDQKU/F+fsVl+swct3gL34ObflVTDbaPNFuC2FKQAGlJYY
3a41ctLIgq+VSQBPTKS3XsUkudMOIxR5kmfeyjoWPogf1GcbnBZbEyqcJhT9
7DO6YlhDa2WNffz+uk7XAnj3QIof1HOSJpFFsloFpPWXbjxo/ed71Zt36KOc
svRhs+5vwOROoxhzQJGWTX63HsmYrXwex85E0LI5yakd7DyY4vWuKv6ltV5d
HoLxWZm9zXa/oCuwdAnSNUcW7PGZEMinMxMaI/0GFCOAGgincol9GcJIwWJT
diI/p2tR77HgYK+SRHGF1smg165uO/LY/lb8Rmid/bKBJwNlPY/IlKEFUKmo
8PdkXgD+1ystIygv1xtWMnjl2Gbl+VPMUjegf72rUNzTh/F/s9BwclHAZpF/
nIzPmIiOGl36yt8e1/s2De7pESe6vPxNn2bjGG/nIHwSnOwsteUKvqkri6Tk
OrygSnUd+Hkg+2DnLKsZF3xOWFZ/9tvElaT6itWR5vO8RR9toI6kAfL3P5U6
R/hKpPio0cLuArC1Os0dEcenMa4+RKGTkpqb4lUg7wgj4dYXjfLIzFXtr1CW
pgium9gGeePD1I24VSI03rAb4oPgyLRxld9i2JFjkvrWop6lSCwkBeCugvah
f0uSD6+eGeEAeLliIxmAuepBm82pBPjHSW05hQ1/vP48ADfKy0vKLbj4i9cx
8Xz3dH2HUbwymMOh/lvz26yIV0bganLjSa8ETRm7D5SHYLbtPsxdECN1Ai5s
/wGbkCt3W3Db7mvz9+byEphzwJZq1tUtK97XVLUPLdIW1O8UvdizdSWWcFz3
hntdA/37nRZYkynVH1Ebq6Zn1U8bRLzO9xMvIbchnZgoTvIRBSIoCN0AZ/hq
xl2d+yf0VmgKK1yJpjcQrRasU7rmr+B2YB+dFOx4VIPOkkQhTYeiGI7kYJZj
HwOIMPf1Jzz8QfgSW3Nm7mttZZ8aIYYPKL/CFQgx7uTTtlLnlO4I5pEEtSQv
wQxWbk1Zo7lm1cabaCEzkFHah3VoOZSe/FYFQfnF/ziBqYaJ4Z79i+YWHytx
1+K9IcDfjc++Mu5mScD67nga9giFmMe3tknUgqXLWdKimjB7xQG0ySYK+bD0
lXnHw/lKcFTX3oiXLYQxEsTVrXK6uQY53/HlXEjvJQGku1rndxc+u4jfaqM/
FFrZJnTXRPO93SB8kEljCRLxlKYIOHKAon/nfJKmNW3pSkrCVKnDFclF9bxW
aPCW7ECU23xcZ0/KatXzU1oatiG6fN/thkseS3217dkoLgitbFC+n5n+6uYl
9VdJtS9x3AJqnWR4KTJ3FOi8xuktNtlEpJN2elFnd5b3djncA2kWaBLx5BPA
tk/3vNAQLNn6ju6M9O6lXNhqnC/TE5Jsiw3lrTRLY1oi/GTLjmt+dQZUF3Ty
HMQoQUscspa/3VgFH4IER+CpOUobzF5+scHNIJ6I9nxBSdPj1iP/Ji4SAeLT
pUnUgVlKRW50K3EEgqDkRz2T5YiWgFNYKFiOSj1Pqw/IfkbZLNW7L+Hr8DsY
HFFw7c2SBdXNLicjvhVtApoYWzEVOQs1pDK4JKDtZT1sLYMArLVohEjZTaWy
LA/9nHa6uUPCPMOle6ZJHHTweOmyQlHIpmrrj/gSrFfHIjcJwblQjbvAkjbp
p3Wsd6H5XMdcGCiWiewj48U6fpUzsjXDeO0Di7P1K9u2EVJwXSn0cJJpWKrN
WiQUH0zE14UgWP0HKVA3/ramkeX9aTPcKT6mzStj0zoyoLyO2Wyei8VN+3Zk
Au4oTlCeV7fWo3jjIxADx9BkQ0mPZzw+h5ERWINmfOkilC41DLPB77fOrH7Q
yXcQdmF3HITdk7yTMWsgI24DjI+Ze5nIwG7kpEhb4U3SFNesnoihzeE8GH4M
04X5ZeSkp6Z0wYv52N53qdWulF6kPxrkCv2fY9GrnQ+DSStZixLeYVAXX5E1
YtkBmIsT3xR8m5UXlIkmvYR6azXQg9e0XOpi1vuSjYx5ctLn0/JQDSd/tqMB
axSedaaj3B1yQUbww5Wh39pRJEXeC4Y7wq4nJlYishzeYIrotCauAZoaxFSh
k82lBIvH1MK9YcFev0Lac5/JX0ZwRaNmT8kWnchI24INltEYLISit97yoPKG
kmzLqfLEUIusb9dCla0E1vuR32KzoprfIvKsMmkbW1hjeEsbpYviq7fDfukl
a+DCuK4FL3Gz/O+QCPTIt6KclGZxiGxHVN+g4su4i9isYQ56G3qI5FZlIc2c
bVoV99sLOOR0C7jk1Au1HoA5rDCJIVeGUv2gDFtRH5AeaedXpz/UX5/A0DH+
WaknD/3Sj1q6iYml9hB6O1rZNVzIbESyZacb2RstxjIpJ04E4KZBLtwF4zIz
Xl7IEjtEU3nnOJk+y5FOICpEEJrkd41fubZvduAvMxZajedWKbH2es83DaqV
j6vRtsuNo5xCOZnVdeblFjiVU4b/+du4yr46h91SY8S7/tWktqjbNmFwFSrW
uDvu26YxB7TJlXBuuyfOMx7hxPfoHmZxUDtBZ91bVaKSu89uphBTIQoVDKqh
v9UjNldTSNXGjtZsn+LtyzRC8qMsshrnS2pf5JeHT0ackMa8t7OccrzEBOsd
dOIRI8kDLxjn6D2K4KobrsGmfPI56ZVKBouKLlkgvduUGecAa+AmQIRmMigl
9esGVgqvPQsepN19r9ZgIwqmELEGgiZnhYifrfEbwonu/5LznxzR9DWZZwYL
vLBj8hGOVBkG/kTfde7rK0Rr8ZHQiORSC4sXUPFeJIcRPKHBBS3aXIw2Idti
XtBrJajb5neju3HbqDXhkngaiaLegbA8BbkXY+QYWpczRB9/MD94wbURazBe
tnqH4CfQ+RuX1jEV2bsoi9i/Qvv16gBq8Xx6Lvoziv61LO2Pocn3ax/npXFc
vUwZjARXBunxjhGjj4yEeraMuPDf2cFrTbNmAan/7wFXdWU28pfwPFY8xlwv
obgZpbu2+TiqsjgJ9tDEVUQxPUCenRqHCTICYUwa4qyWVFsVzs8Ka3kytbvm
XtAJVzZRHrS+cBWNUdrD6aGWGJ74jmuB9xV7L7CQYsG8M2iraJBR0cxwclwk
WYkVkXhbAz/SgeMP9RI96AwezqetkUDX8OZWj+XZjSb85iPwumPb4O7LYO2T
q1rFO9LhgJ8LER9hx6jjnF3v7h0UwzOge5TKPMdbAtqbYm91eaBwJ2HR1bll
Idd29vQrj9nJvzYHAF93QbHVfwlPnpWQBrEaxQcDwB2jmWYnFukTBZlPD5cE
/plNaxL2zAzn0RaukSStPkYGZKigU84CJVWbOe7MVFRnZRtLfL2ioJK+hoJ+
PboGfirb8Uoi/0wT9mTVna3kuw5eEGthgOX+JjjeZOfWV3g2tLscCx1m2fT+
zhLSuOMWmhcBT/Vw8alEbDyw9uF6Ue5phzDFLRb8D3nEuPauthfZRJZ3lolK
ipCz6IZyBHmGvINfMfGsd+FCaDCpkDC2jksNsynswyTst3+xv+k1r3xy6aEv
NIcps+p3mfAxBAJDPzwATUaTxT0ux7eC7AzvZzZAQTjGdxeSEQw9icZJE3eF
RzVII6+RUc8HX0YgS4Vd26a1xYqLySmOGs3hAetbCfOOUKhk+iVOIPmW8FQm
7N1ugZwVs0tlgQPWB+iN0lf1YWiap79LZdyobryCXhg/tkEFiInvfD9Xprxy
YLPkgnRZ6/KmtXOPU/byCCvDNFIljXG/tWoI9stlZFX18uHt3uToch1Xrxw5
vxKHkIcJRfT5qrDDkLnjMbnuIkoVv0T7hBJbdVHeshHd1HJM6NH1kpgejuMk
4CVqVsUheOUhj8fa1UliG3l/riHJ1hhNhQfK12WDXGzeVOa3TWWPNYEuDuLI
jueOZHv4lUnKgVsw22iweiYXQyDdYQjGLl1VVMhBq5BmwAESBZZpPtW+kRHA
Vr6GM+v6H0ig5gy3ghGL3cg8Pr6WZQwtZd3aTtdsOLZGRBnRNeg7FGQTPsYH
Cl8+xQRUKnkoNoPK7jI+slZWTIheJ5XMNRhMziqnr1RzLf9DL/Oqx32+qoKM
7hmhsUBgTsbXKgNXSoC0Z5kFstdzaCKxs+BbYfBgcqVB1L9SZqpyPDFOt7ZH
D2jXlLW3HdsmHk1IsGSpgkPNRlUayu+Guxt+r3Zb7U1n3Qt288uSjX6Drc5l
yGEmS2zcJRWzVABM11IcPdTtb4/EMUw8CnHNBubzw+oemqVYRm49ofTVstRc
XycEKPFC5PcjBVgoaLM0cpbcKGjZFnUMPug5NKDn+EoIn/m+VOjrfschHs5I
tQ7GqZ5ZHCV+YrVv9e8Vits5zpVX3CdofFy/MhM8/3uFXdGkGbzFRhnpQaE7
v6dKz10LWL0BYCihmRbWD9THwwImEd66mlETyhjdiqWHMQvVt7ZzSBm87O/U
8E/LsRGi+2BMBIGQGKdxyAZUEgPiM8OA45xGa2+8x6MMBiINxClHv+yZsvDj
un9se4/sdGaYSMNK7pSiHt47zq6n9cRJJ8wIvnpOoPRWDQDoa6lmOxMHq9xz
RyoyRKWa6IHAGVG5cTuA8grrR1SfXdPjVSPHljMuA0nwPlFR/WGaze3btnu1
ecQCQsxz17bYLLm519mWUcDZjjArOBCQskD0nIn62Ei1qYt6tGmQOV1nBfO1
VJGFMkf9QyPxCSQSdBecPlBkMY1dSCGFkvLvwteBaiDrYAhPbt8FehDPDpNk
teppbhDzZ/TGhMejRKwY6zCbqPMbY03SVzsB9C/wccORFu4kxQBLvgmFT9f0
NphYw6YEpX6h49pWWdzlcsIbT5KmLgCwlon4gyqrt2FSk+2kBnEt5Zhms6fw
3TE3T2NwaEIlnPrcWU/MSvMhb7QaczrzYzoNgFhExIS7lG+CpDWSQ9a8DMRZ
/9Qo9hpHbpgJSs7WJezbujeM5yFrSonhzNCbR7HlKtzZE0KJ5nlFt0QsVBkB
XxYNMS87kO4sb5bhAMhB1qmD/ilOtk5kqxuSxla/NLd8HXvzVvZc6n6rDGUl
MGcdnlar2b7Av65nY8z9jyys3rj3rRAO3MpIpRKNnMcUaST59dul7mYBc1Hn
QQUJudic1aG5yX58SiGHlmYAPMD85gXbt0EH6CuR5RXLXrbhDAYF4T6JUROK
GKEAw7nDfOIwMsvJJq7JHACl0Y/Ojt6fUm5H7voMnc50k74pNI/TuyTSqP7j
i0v8M69zF/zm/VftS3i904IjSecv5PHlnmlqoBMKUAOgxEbpQh6kGIp7rFX0
ibW5H99GDRz+O990JsP6Ss0DxGN5yPcwnYtePph9gtvMjho4zPLNErSmUbAk
jjBlu6DpW4+PjcaWv6ghrCzllrOzqGeFG/XvSfJOahUt66PLFUryP54hfYW5
irm44RFaDYiSN/iJJUzBqNWY6MsxhEnes05CHUOlPQ+Ag7Jm7D231ICjp2JC
/PJULwoq2IfyHaU0XwlJjAxhi/olHq1gZn/GJI7332Tt+hgAjw4YzgEQj8hV
kI2cz8+GtlJwl4OX8Wi4agFq4XDmw2x2orHsLZ9nBNN1f9S7j4XZnNYDZx/Q
5fm5Bfsa5iZm2joMJ1qCY2INrTo1eCgEcNFLpMgwfmlN/Np7FvriRz5ARQKg
qK076XdQzJ8U4fgjZB3rcn9W7yc5j2IWg6sQlwhDkiko+mix2xuz4Hj6uyo5
A72TXv4w1e31GIN5Wlxdhzkh0c5xt8rvWOaFTJ5Nk2WHCMcDOlymEM0fyhVV
6u3+PMIESLXMV6T3M13llgCv7PFdFSqXvwQUkLpwjxDE+is59PzCVdYrXxrz
wLvdCAcMXMl6wqnQcPNyFGTbvFTLf8DFOxm4blozR2YPE9smQhs21KI4IXvl
bpDVCHPwz+LDDZSVTzRWTxYTpij6vytcSYYpohQldxNv6HXR7pcuw1CgP9Uw
9ujQlaBqL9/0TdlwIu/utBXEJjgroRyWrmetKuAIVjrTLmenNzmdDAbnC9m0
A1IKTiGk6m3tRFzyL6V7rqRpezgTTgeOyxIrAM6dehSPtHeqLeC2cqkx3GBb
j4cQi4eMDT9gITxJokSk2r1VnqIS0VaAJxMr3dRLtq7zHoE648IyaZiDlG8X
P1e1an1mAmETrYjDO37cMdxTJbYlq42iRUeKE5N95nTHiwKz1YvNDHMVvydl
g4Vae6v0++2WwQMrgs3I1b1ijBDRURwyAna20MhOIYLGy+20sVFfC3eGEES0
s73UWmK/fy9mZejN/eiigpbS/6k2xwkqxjAiAC2LmR+26EW8Gqt4JgUCx5zu
1fXtu/6240BUku/25XsqC4MHaO+Ve+Gei2ejF20vLvg5e5Q7sWBerjq12Eme
pS9uM3kyxtV7pPmAgr2o4yocLJkDjI9ucSfXt41kKjFM9/JVwHkSsV2O7HIp
dcZO79IqY0keL7xwkQYZsIHk/TcZWFpzoU5MP/5195ZwEb9ZzcrZTclv7heQ
rrKRQ2Psg/dk2mXCzlgRKGMQySNu/bCV/L2ZVG/N7aJExsoeKrtdrKA47bHt
TPbL7owxkt5Pm2QiHVAxoKe2w7qqWT+R16ChVze+kJf+IdtM2f95mnv3fIte
oh+8UvE6fFry1hEdvFZM5a7JPIBYtZdcb4L6obz917nbiGgfQMSyjxCxFyzi
yy8yAzw8gDcjeEzkwmJX7I65sn8wfbHnAOkQjpHKIqhtrYakxiZfkpIfyNd4
qGxG7AL40VIeCaAEKM/WPRp8G0lvoDNAQPIrXZjDqvik3jqwjmeboWIk3cuc
kfhoYjGrB4HJAJXv5T1glMbZShFZXkO4/EBVwY2ClCch09gdx+vbbDiZX98U
6jnh8xcWVgDWXi45/vasmNjN7T8BcY6wMvwws7VJHugc/38naHpxfkn/Lzu/
TAiMJj7Xx1Ep3gO8V1Lb/Q3HbuR60cv5tZJvvdiMMBmlSDZuO9RJGFAOYziV
3X8ffNsAaMwvi6zaggLSp9uS1Ngs8M8upR10jBx7zfzFgPQsdu7qn2er5Ng2
CCBh0YoC/OO+01l46JCggmMFa/vOcZtzmLqwGyCdbV8z70BqyQ5S8dWBlb9I
mO8ZGxJjlpFIs9LjUePnBPdXeI8t/ViMivWGT/iyquczgFj+SJgzj3RknlpK
joOb0MQuWIWvJlixqew1Vet0e3aIYe2MkKqZ+62QEGSz1JNyyJNSWlKGBejb
hnjNuji1Dv5rNTMHXifI0Oe7THnmFmdTY1VZc8fegpCgB8LJxHo6IiqLIJRa
OaMW4+HrZOVF6Pd9Js9eP4++M8BXZMa8Meu70a4T91aePgo9/wW++k87w3yS
BRux2vJKHubcKJbJLRgBMzrO72HIWtpyoRPWgp96VYJDgI0BT3Picp9iwVw3
JIPE/5CbX1Hj8MpsKAffxPmBvWPDzgvaO1CHm3jeoXLySfPFeR9ibyW9d4LP
qiAiTC7Ul/RfJnYzDIWbT+hlrYZkkGIAdB3JLvSWKPUnSAqE99H1SK+AnOo7
utwwDxoUAAKONU/ulGj99E7469Ez4CZM5MTJdkEH4RDlze891lATf6CPS5zn
tQZwSog4xljG1PdEHjL1wk8cQtGo0po/cdX7FJVIgdu15gf1H1hRmVpC9m3I
pYVtKlZsnLcymlbene+QWyfeh8/bOTcKyIazWjHwxYZbwNxSvK7nuK+By4pw
2l1n7uokxmSuOfo4YSDElUV9l7chOveifIOpHEXHIs71FHc29XTjzeVxmSMs
3JBJdzzK90dmXoIcFgTz5RPjhhdZMFQvLdmPccJd2Z2WV8S+6bdeuP6AdhrX
mI3rmiSR2y5HSxPNGwyKAEPouJIamsVfsTHi2++pvf5EK5N+YUCqflIkofTx
4iVy+1zlXkeDPBZEEecyuEBHmj6QhOCDZkSfVxIE55Rq2ATw9BFWf683a/QI
t7eVOTtkOsb6odVEODoUbW8RRMFUxc+cYv6euYsV6Qearyap1Yh0qgU+MZ4C
OgbQf8UYdYZSA2YuygIeanE1C7KZFlXpCiMv09CnkRWTxhStSjiHtYCew3AS
E7sydRpIMleTa8wujZWvYnYieAFIEymcP3bMj1rAMUDllvP7+QQOJHwDnJ1n
FbRX5nqTHQWh8FE9WftoicF5e9Q6VF0L88PFdghBYeEc57OVJrJibwPZsPTj
glV45qAQwsX00W/PT4TbY6kV/D18a0+hMutDOeIuyknbpu7AXCApbHqGWOjz
fouPFu8KDZpGGrmskRKkDUmzX6KvQ5+3o6FdLcg+wo4ncAIVimVm9MQ/DMAf
yAqUMxGDaC3uPv+V/8Hmf6Rr8vL9vsbZEIAf/u9ikYchUTROPcH94hWkwySX
60TwygZFlYW9j2e1FqOBzZlmC4zG1jMGgkzYo39ZqAIFDqm7AT5WIlFOxxA2
ee7z73786dY0yqSy/T16BfMc4gjaNZTZzvZg23MrkQQwi39bvBKwh59jd0LN
Dkswcayo4CweKO8mnVBaQz2m81urZukiWDE9MXOp+uAKuLL4j7hTaO4M/LDW
pU5ZB30JOOT/+9OmCqiMPKXQYbwhD46Rir4c438ket5WxzYVXOOWczZcKPqn
0wZMxVkNQnrORLLOO24E5x306zw/EgjrGiDsrIKeZoZ2fP2T+gKnX4qjURUn
O68/BIjEj1R+D0sswToID90Pb6ZHrmJIDLx+zvCUi8NhR3wdODr8bzbEIU+W
LAABXCR9c9Iak/v1WsPhfJ4rAZZsmDe/7MYA+DS5Y6c+0BOzu3QljkEkPDu8
DcdXm/QAjnueKbymkeSs2SQyzKFv2pH7PT7iBck7Zl5XsIvMq+tIfBar1kie
ve2Y4O0VpWPq6+nJc6pNR68GjB5YKIj3/oSfqVkd/tdWzWj/R5HI7yY4aBqi
QXb01zNzYxtCYk0QnS8CzdgyiGX0FEsiVA1ZUPqm1T068Pu5WHjualO7uZIh
M1ewMs2gWT1DlhE+WObok9GW9ct1TZT3KzX25HUn9fdABJdeX8mkOXdAvYQY
mP/7Omi8nDR0CUfv5Kn0K1ivLSKutG2gDjC7drYDTJszJIXIyUD0BOhYq5ek
vhwjC4Qoeaut9ScFKFYebYMWvYsNmzxMf21l1A+4NSDV6rqso49RXUuJ2l8F
fqAwhVK0OaDDDENAhvfS1Os2ZIjWcwXyLbJVy7MUbbW4klD3Vy3dSy4eWCqi
XoFZmLKlaONEdRLqUt4wYl1SDfYlS1R5M4BTAUb0Fy9A3kwOq4GiCwGkzRNL
arzHgPCSH2SqK1u0JREVtqrqvlDGggLLBsrb3Ply0s/76I/4Dz5eegyTuF2K
MV3UahnBqMztyQNEm4u/NWWxBNNTqc4CMqanjkDSKBJWXG+a2anyU5X67FYV
mGgUlr33y5bBN6Hi/d0/1lfiHpi6n02GqpibtKVXojXmtJUT8zS1GoeE+TmW
Cur3Szngejv/w5ZANMXqci4t4GFfL46gMoynXfLAtvkGIMcIpdI8hIy+DvkP
TvfyXDO2eBoeQL8960aw8yrVmo3TuPf0oaIJtN9sFd5maO7s42pD6DECY2u+
mdL74FyCgssjsGhvX6dw6qQ+iIjnDlRqDflLN3EC/cutR2GmI8yz8Iz/uHV9
0yfPVzSNBdGbLz7WFIW04nVS1me8/ZSgr+YLXdvMN6mBQxEzxNpzOHB4UG7F
K0nC0APpD2XullQg9EuYIqbaNi6u4qOeIMpccT+nxqS2VsJfxxXRYkHg9UW1
M1ojsk1dncQNIb/oEdG5gcBTjnArPCNGV3I6+y/mUGmehMuffmFaOmG/dWww
eKd11t5x0mWwLylXFsuu3jX2LHMrZRn5DlmRQmRD60Zb+LJ5HeYlxN8cBNTg
LnSHtBprZWDUIqJPsxsvSntSlmmV0qRYQRq+in/3AxJxRUYh1YQo7+I70deo
0HswfoLxShmmp1pZcTy3b+U8wKB8Fxx+3eonNqdD3TZtJ+mH+PdfBV08TV/S
UwFf0L984Iwa7Wc0hGAW40MY9zExC1XuRES9yXMfAbGJjXw85kSUkDJke46o
+xsn1MWoeN8eVDaGHIEGxpUAUvNkklaevQbwutLYVL/XNap/vXdzCZwRm3ZZ
4zbFlMyr6VBz1ZXXLSwaeqGWWGES57kD36XfBgegJy3wqO+KqP+zb2G5Nilb
5xGFBOFBoFpoI0bh/5AFu9fEzLO0o+agTC9s/bATdYz6s54LUuhWupVHLa8Y
RXAgDBPOq0heKLSETOJqvG6NA3B4fBg4ayEw0UlywCFgpThS0nacjNxh29vc
XpuFMDV6iIJzLABukPYoO+AE3VPM2607ANnU44s7X93+5GQCCyxISii8C3M8
CkvM7wFrN2sliq8bdar3mRjFyYA0kJ0NGizY/MFv5BnqjFIAt5pX+fIFSfUJ
PhM1aP/cbJYg1V5VBq5dZwA/wQPbO3eEdkjTPnqhE/C4mwrGNgyUWijCYSj7
u4OtJCOC22TJtyeXxKi3vIbPg6wCveqhYT4y4ID9pxbpem/pqB2Tjb+LqgFx
G+ujEfGc+pY11SxoICG4UC0MuH/5u2P9ploMK3oBHeGF3NgyDApq7k1VXKX+
0GaYchjYubmVuoHFebPaEE1AsdJAuKtGZwm9XqVJ8h5uUy2Gb2dG4I7m1bqj
6Qyix40UORrzDzo6sqn6gLMU1phL8ZL13e2uBkN8GdIpuB2Ds37oD/nebepv
Jn1oaBnt3dcu4VNcLeaFSGvIXcP7FMOqkDbZgQ5dfb3N0xXWTMDilbNoLbNi
Z7vzBI3O47uyDIX/tK+uzDGPcPUC5LqMgOgATvHkHueiA7VVrhGk7CHRzewQ
eg5MfF3EYLHE+GLjQkV9OrxZqQAPQwQ9lUH/kxLW9BUmQ7I0H0Gcox6mVDXB
afYm0hV1P23cKLqXXr47qHw0hUuB/XRZAKXhKvLXRB5FqAm7stSmZJOqjhK2
+Qxcbkqmdm/ozfFf9Wy/lj/EJkdAD2JaGf+9WOnu9orNkAzUPNa5ldc8PNpP
/mtF7W4jU+B5HP53HEB8Rw/N8OklayXn4YqoM8ngcNT021/2NzjS2JtL/pRg
3Eg12C2ACfDumL2Caj1W6vHVngV+Zis32g6yU4sIQCQMa4Rd/VUXwJENmwcl
Sdwo+uDb+Cr2uKPY3Dqd/xyqPt22TQCwqKAD5yhmBZSHdcuWMA4/bKEWJYQh
7abPEiS6SuJEUvtY2yFpReKDk68g3hQyv6OHJaFlvlp8W1HndCyH6ChzVbA6
4BLvWsu8i5av871Wch6Nn3OGkIh2SCVQURXzxvZ4XN8pve2zm6ead8Sa9tVg
7kW6Q/FCLpQ6JRMvAOeuCPeBdmL/Pm04oVM+G87IxqsPWfuf83M8uqXI1SEf
IMTtMLJcZvBYIbjRhs6GKCrRnlZJPo4c6bXQ3PhnOZAQK6U6XnUWXuqOzkWJ
t8cUmIV1bbU5K0HHsMf7nICy1ISz6Xn1/cRxavCfrPiyUCzg1NhPDx4Z4MDM
EziVTDByxYyhToH3zMjp1Ufc+/nyG0T/XBeM3r2VfdLqRSxdRRRwI/jcZUle
u03H4jkCnL637BX20ZKQOjcBNzhvQ6QqSo5t1Yr3tkVXkXxcAq58OhqL4Vu0
S4O0PTYvkMjTEsbKiiGqYkr83eh3eEVihCeov2Nfao6fQ6vkw9HtGbH6adan
/9I0H7SbaeSQEylyGWdbt17S5BPk5HUxJ9rTaKshoytgU3lZM7o2fx/Sn2kH
g+6fSuvikg9nl8ejx3W2liJQfdbcS7hCrTLUox9c+hLTSRLo6v+2K2eRfSma
ucoHUIqMAQ9JwjdKMUqquCP2fgLr89RuRBlxvPUJdDXvXuGEfNmUXZRQufp1
BLvmPPGyqyRyblLRKzt7aTNmRGwZjmbXAxPtvX0oV+Pka5qauZaVxh2II4iU
+YD5TpKYqfMJcJzRe4T61oK+LyPUT5CSr3uv5CBe0jfOnYUfmm4w+nMvLmwi
3iA6v4EV9G6xkjLkBrWTl8jLhGkH7MzxVY7eoQKfhTF0fsi4m6Qt9TZbWCKF
fEzHL0GogvbahwrTpXb2J15SYDXnoKkJ04rNQ2sUj0j0ZYGGOssWUE/1RW3t
T+hwyDCMBiTTt+wXP0+TGMTfh3wMnNG0uNS2t3SZ7tAa0Nff52Z6a2s0j9TE
io7VUB445gzTeNMEjlgKfjhediqEla3GWT3x0QijqfzFBJd0+Kb2DOScrara
EPdToymTZN9hh3ws3x6Wry1lyvbp7DUj41vGhL9C9cku3GnEgfaeWN47G4UZ
4bda3CkUrBazKPUpvB6CkubUGagi8Kevqy2FyErXWGihS5npuykSFa5AsU0t
UpnQNsrPC1aAT9fDPx4bRZjKmsi5L5QmA5IMSvxxVYGBHZvFmMDui+HlsBXg
f2UzTV+BwdRB8lareNR+t+4WfmG6G9of9pyfD2/BuA2bWBHX6l60rVtF4SZ1
AIaZxhhdg5p4FslYjW2zNZy69ACyjwnktn+GN/vFpasy/cIpKo5PvFOuEKJN
RJjCOkZ/3skMJSxznBlgZsGtsbhPWFv1eK0m1Q7SPRZHqtHlB/JPUp7VDb/o
3w9qANvOY/f8Pqt9SRKCS/VNaJcMB6uoEbFThnBnnhdnsmsLwlF6uYs+fgU0
iamG6v3gHebpwJhxHQfCkQAlPKBd7NSH5Toz/oRKHvLHUipjmljBNso2jKKb
ZOy2I/vPlvCM5joZFwk9e/QbttosBsPzADwrgjLY03q8n+hrnlQkHSsaY5N0
75KQM3ApSeaz45RPXs7NQLowgRYTS6g/RMFWKgPNccE8rBTjavCunqMC0a6t
Fpqr3V2dKqGOvemTYjdR7oUR0Oux20/6bGz4borjhewGzg91rYE0OGNzP/8N
aNkTNF7r/Wd4PH71YAtL/ifeNSb4jqn0uLI38poItXQGAqBC3rKmlP3hr5Bo
lF4e9aN6U56F11ZTNLjzAKw1ttLDOc3Xc9jquDygDwgAJgCewo3JuuHHNZLE
hFpHTPS/gH/2DGQKgB4MX+7YekF1dMeryzMe4A88swIvitTzoDWkXfFSNhDV
hNXNX806Tpp9urb0YOCKDnlf+1OCxn3uuoIuGxfBRqIrn+9fh7S3IJZpHlUG
dQApiGdosmroDFWGRJ9EFJsE2rQZ2bDnU9ETgNbyOxbBIEd6PR3q18KFBX2u
Jq/TttGEchQX6tlyapSbfmxYfHU5EL04JqDXKpiN5tMPuCGQFeswz/XgsdQG
J+ONjwqBcPcJy1QicjBWl6O9i8JD3B3E7f/xnBBJmAvzIaqVK6S6wL+xgrx8
kHYCNZhcyfHJDAwbQzhEUoWxkGFUhL0EK3T5Vxy8Ej0zLzDAZOrEZwtcRZ0l
Usv2thjQyjfI27NAKKNjhL1fs9P/jwC7us8hPxH9n1teYtnJnVTnGRLzylcO
Gf5WbMHnoFw1J9/WwF/9fITP8Cwy0nlLn0UMxhnpk2fV0S4RA6M5alQkASiK
Pd1/8guvZNy4Er6TsZNiyD6yZucxPa/3viVtU/jr3AqQkMRu3z7pFpdt9dMu
o+D8w/2U/v+gBolrfJiqavlku6Z8UoG6G+cnhuWo3qbUvPDFdWzLUZK1/3Q4
RUT6Eglo3mHKK4PFtzFVy5yg+/N58weZoC2X0C0lSai2LZzIHF0M5nmXHzzh
sp0RM7ZPj+A64PvmEdI9E04ngEwwzyCHWR5kMJoRgokHLlVOJWgcXq/6ebeA
c5y74h+aAGAzaEcChV4OE/9mn0Gsun/JkwuwEVVd/V0HSDpAysEyRLv8T1LX
Oz31WwpV2qnVJN0WrIcehrKRuYipYQBvg7XhDMsbf3ILFGH5V8PlUtAS/d0+
jq1Vpa6CeghqOwfhzSBxQM3Bcg9h6Ja2fXlHaqYlzb+q0sNKCMBK2y0D9+JV
/QTkpYE4lYwsmCRjP+t+957C8iiyMvs+nwsinIs7QvkCx+XYDDMgQ/mbLzLC
qmt5uasbDcAbIy9oqttL6JQBCx2HLnnil3imsBgCbJzY+tABQQuVyi+DmRzX
5USx25sNTf2cClETBUF3AsAZUushuErDIyPOJc1Q03nuS1/OphynTCDSD/D3
cxk9mYyhCW+JVtn6SatA/r6922YcPUa16aECjuiS6O2BfdHFeHC/ZqSiHdNl
RSomS1IAf4xVumx3MgLyftpCOHIL/yLR86ZIeGJO5MIg0w9sa6IHrShic14i
/H+pMg/3LOv678QoOq1TjJw4uXQPxZtnv+XCL4Wl7ViNQsdrftNGp2jdj23x
9xHLOtprGyrJ5MC2J6S5/nD8iXw9Pxkm8yF+zOgN4CW8l1unN1oIeU0fWG5V
y/TGjKp+e6t5KLyEdfW5d7GUtEmjzQ6AIM+LumoaNLsBFzJ/csOdNlCBF2Kt
hzR20meVWkhx6VKPcCJ5TbaLkwkwOPe9x1d72L5slSwY1kWdiY3kBKUbNEMo
+pOp8aBYK3LqNhfcCr6a2xfFBirFO9rXhV6K5mqVm/kKiYuyY6/YCsBM2alH
oqPVhxsrdua9S8MeJYXyuD6PWp/+uVsUQIQq4VdexU3BZkeuuISRyzB0q5YZ
3SeePxqkKDSXp18VZk/ct15Hp7NUScRfiZCpQsXE25z8Fk9YzjLXIWqfNPL/
EvmHAcf9wJYNvNIg9FEswHis0Vx0OnKTiAZZgVCJzMzElf2OmI7SfuhZn6Id
4sne7UpNYyQno8NnJuhlsZ7dPfJ2FuQgO2muExLd/dRXBoHhN7JTgDJTx9oU
OkA03mLDfV2IG1r8LgIx05117/JAOBedVzHjFZv3Kmbu71CEtM4/5sOtHNsz
ouG1AHbaET3NnEB3fuHE3aP5xxTTbxYnyY9Qp/abuIhjpLzXQoaLJjamV5/G
Bj0jQr/PSI6C6Gp+zs+p47ZJ7s0BvsvH7vm7J9LnjeqeYU7puIZWWbBx02LB
Y84xsuv+JvxgEylTto0A3jx0Jufn3OG9qV4BSEGS2j9XNw1rwRvkjyoM5dzA
x1FiM9/WJWW8RwWyAeDilcBPtVJ0DWTU/Z7EORJdwI8kn5DoXgOpDcrdahyz
T2D/EZlYbF/8xhP4jiQ7zTIQkwYWlKaff4txO5MFi3h7owQfnhCWVfNWWFGx
iBjqBjGqIEgzo0cz/ihAu/2yP8MkCJcAfjm2SYA8iA1jWPXsbSomXxjXiZBU
WeQDbLXzVQDatdkabUaAS4lW41baLoiXIlRHMp61L0uyBfJugw9rOwWHgrhp
/r7DmgTNYAIIRTXOQWjUTO37hbt7vhp0058wUMuNQ8sR6z1RWdfECQfTJcl8
l/epjV18vMeaDbLmJkfM143NX/h1KpIr9K1jLYBTmZBj2Rq0rv+tZvvEZo8p
0QJXIF2yqp2bUijB1BtaEh/LFaAWIoZAufG+AyfTSK3UfJh4cjiebr+ycNne
bluOQ/juIaQcdmUP1F25KGWrd2R6VZa8PrvPBVstaI2HXempF/rB8M1Ijt25
55RBZxNIr69oWTfmAbzy7mzH+f+hoKP22HOG9Q7c/rqeiv+fz/va5twqil/X
Ttaw1Ew4LPJU2JmcWYa/jWHlY5eRaWQxqYSwaNrWNNB8Uc3SRuv+oSHosYjF
Stut+JmwHF+LFAbrP6AC7w/vxF4JpFiC0/98l1Me5SEzF7c+vlHSdGNt8U5M
Y7sJ/hfBb4GG5kx7yAuo15zztz651Knvik1VTbKGRitm/YRjW6ncHd7m1hQJ
qYgmqd7ug8P1l/ryOSK7JS7e3C9QGg7eK4lVWOC4e9psgNX0muPGZ1hMjM7k
L7L0abTlkCwob8PrFghMUn/2fgXn4zL7du4XfYReI9d9M2J1gVRHon0fdzru
dyefcq/SqJmRMH4eaHOP4aqqLrX8jpw/FNWktsCSnbT7LWBJMC4AEjUfbLnK
tp0eUL6ToxtJdD5zG436yITwFhm87SP37dPcZ3SxGEXy7kuwYIDADum5eOHp
bNyYUxpPinne7oaJvoVegYSM5Kd3IRX5LGAafXqJwJSlrAGtiWUbfKwu6DmB
nOXNILFGALdA51ARuKaN8RmpmYqSlK9JXVxyUoixDKQrS1lH7wRBHgwCrhdE
m8oGlwxPPVCTYJzxxpnU3O7eOtHy0L9MDUae7Yt8J2/im3NPbbUmA+1P3a8I
srLVmiYctd4BxBvOIsG+SNIiCxl7digt6QafxlY8HkG5hbHBN4LQwLtQxtsj
FmYFYAv8BOpo0Wi6qWJD/D1nWEjtjS+vNPbSisu4XAcnnBvHZDh2VCGZK+Mb
ovzoYZZmFxGV1WCQSmntOE0C/65R5VEuKQX6Ya+Y8TTbjmjSWpAfKnucQH4o
71msp5njvLLGc8z3zVxNx/SmYRXZcZ6L+dzuSmx9slo2YenEKwHnixPww8iY
szqfNylLqBR6IzdsTAUM04Bet0kLVQadGX2Uajx9SD8fquVWmaE77UMn6/J8
dEFlKXmLyRud+vKKp0CLdlP1Q9+F9KIz2b5jGTJo5jy1Jb6+9wlFqCbW4yIV
iPXmtb4yNeY+wwGf3n/fXpTyi2ipPiw4JsFYwjheqP0fzP/2QNO26qkv1Ci2
4r2aKfA0HWPO7EQ51e3Ez5KZ0U6LIblMH+0el2qXZVTVqbmKsC+DP5jSZr3O
RIjVOwKKO9w58pgYGWGUBSGMdzCugs9lNZpCMtezSRzu4qhpXy7o7kdifDiH
Sw4sjRgHJCblP72iOgTBCK43y3I7HjKj1Ro/yQT501kfQlTeiTlucBoh0TbS
s9dbo1DsT9HQwHOhHV6UdeiqE80rr53HtTg4ioo91HXOFCi0oo1taN1fqI4h
SoBBoM08oJdgltDGbmA2SnmBilUNHWAMFt0ImytJmVHk1w/f0iNkV2lAeQly
JviuYqt14V1NTqQTm2Fd/GYxvBf2yKDh2xGNvzkJEyFHRTC5IU6LliMEjkCN
5pxuV9ug6q2bCDwJ8IAvcgrEZ0WJsTbp2Cp0BfjTzXi8z5kRcUiZ/hAm9FiW
afq5H7Be9wHeOFIPhMSCzTZoBj5s8GHO9/vVJQYHezmwFID0o1lwaUjW9g3T
Yoy2V8QfFwltYzFB3xKO50DSPtQ87Ug6MHUbGwZF4PJeVv1Kxd1pQPsW0503
bmg5R4MEXE/0/DQ9COdqwcSjlvUWpsO8SkLOq7u3k0zMK+TIZ+xY+S9UKDNb
kyruZPk0rdFRVdOzqKfY0jEs3nXtJblrlikreus/EZUYqzxSgcKs3JvWiaGc
RgDXChLXqsVKkKi0i65jfkaOqy0pQL8/Sp/PYdpXctaGgd4qBAaD4o8tRAse
/OY2TEZ+IFI2TrUuYoyuaGy14FaINd6388XRvpewMzKRE1A1wyNKM1nSOhqo
HqagHdp06bhwbK38h3xd64F+QU45EaBtaFwdJA2acytWlYlAqoP8//h5nAdq
+epiR0TcUaI/X2Y8buqVNfNdKYFOBaGN3lgLuF1FqfpH3bhJ+Bg9mKwBNPeQ
k6GEwbkE3vi9r5EiZlwT7hQp32Srr+1s4SE7wiXdpRmf+VFKPtpuOTjVsrIq
LM42ErrMuStd75KD7bBkBLMHeY8SVjjojfEmIO26cMRJ5YNEJ6y5mNNZD+C/
9T+fble6ModHYfVi7ZQejcXy2+rS0NMcVc82RU/zx0zGUKiwndyFSxKSnkkc
MHjr1xlBwUyUXi18ndCec3gN54SjQulKb8H2YEahYcBipsCsHbfH+2JJ+dQu
Xi0gXOdDKF9tjWowoyhKj9UJ7Q/D8LhrdfVjPIITrzxWXORwB5DIG3UpSMBZ
vYVubZ6P9xYhOzVCReElnUzWprJP8sUV4v2GtI7U1QxFw7lCx47J3hSv1U25
4Z/UeyF836bYdwQqt2iA8772Equr/UpmIFHmqyIGy+2/Pxwqx7n3SHGYKpUU
Shh8i22GH8LuN0zNOLMvBy3avijlAKe/8OjSRFTvkISL7khw1wGF5qnwuGkl
MXdvyuXdt04xTVlOwsAsF/9GFx/AaKrj1U5EUPiLFrrhfs0jI/z4w0RoUcCY
RMxi84IXYfu3chTx+slpj0gdxtVtF9kyPxPDjQqExThUIWfs7RyKShK/aqwD
qcQkmfUn3BYxUPIHTVks6WHGTyg2GYgrOMc8o3/r86gPlZFdqQ0uywbQBqsz
oM2TVPL3aj307AHw1Q4YrZju8ZM+/+WhNNBC5DmEHBJuRa18iE+A4fP86dWi
gbp2T3INW6LD46d0mdJ6hIFbyJFEo1/ql5WVx70qpXhs4bxZYVe8fpHSJo1t
rCJuuzZyH/tCGJdI9lrQ8ThcFP+DJojrOf7OKCsLWI0gaUzflNVaJrO4A7py
UfmVRD9HL2C7Z7SWDZa0pAr557jaimKphbz900JX1sB+uNlh4l1OGVLwfpJm
jMoI5wqyYef3Y2MY9fTh2itkhSm5iVzF4tL2GclX7zKRNLxbzUR5hFFEZZcx
CIFNvHzgTOclRy5iaUKlkhvRlZlRHdoZHXByElOQPk6q590ut4PCrgPwWyMG
+hI5IsPj7g6BxC2UqqQ/E9v4hVPisrIbFL0txCz+HakLMPX+hwJs3ZsCPfmY
c5DwcToWK0qjsf/IDERjXztvmyS/Sx74Rg03KBFtbath8cSAm8zqXA9kiyx4
U24FjQ33CwoceGNM1jkOQMT/k64r7qaAo/u5TBHlgmh4MRNfMjIeMIidzEUl
ZSeWZg6850cQR87gbzlmFDRXS7g9TXMzkKbDKt4FNRmYNT8T/OU6maUgkSKh
Dy4yAGvHmBBcnp+mjaKbg2GpRsjLlUASMrSLNvsNWJoxn27qJjhD9kUvdBOD
YOv34sP2YmDkewSJfqMq0FVHCBsZME2ZMta9suys4WLg5NUGVci3zWnH2/Rz
L9H27gdfQY7v90vgLD0KcanshnHmQSNznm3ujayyvw/0ZHrPJ8ufW/XMMtNV
eY8HZKZg6DgdxF8mkqM0UzWcMCUgYsWM6WiUgHfyKiUzGlBJdDUMzYevUvkJ
MXrXv0wdDhh6ePoMcCvdwx0UWPZjr213XsOrobeOWRS+B5Tl9yG7Hag0HSNl
sZc7wyUn4JHcDpt81w5BUF1Rndtqm3PfqhJrmNNENgCNCibAuHqG0StbCGiZ
iQKk7daGWP3ufen1U5CQKxzLsF1miTFr/MZiNCFE8vlFgPkg7RYepGRgPVPC
dL24eBa2Rp1MnJrnQtFUet3CC5ugVLi7qNMxn6H8o8dO5bXl65mQHxOYE6on
Hv2Rte1fOiwezagKhxqjBj4rwFvW8SDHkpkGcZTStuJskV1p4EISC8muk/93
B94KVZyJ2q4uLjY8gFD10edZPPfVMlx5HoPeVgRh1kiE4qyThHuburmWw2js
Ut+X2cL+9UQG88PWIKrQFfyy9uQVZiGR0/QS6VKFA9iVmwXu8vYMNwQeAQ6U
LpQ++ad8l/DdX+Aofn50JzdQZcp753nGM3ENq6DJRD1oOLnTq1jM+pB4FtX0
ERngB9dV2n9NYZbKjVgRkY/nPoLDzaWK3SpzIvfvSEw1KDld5oOKxuL0C7NH
WcejEtu8ncq8qJhIzr5Kbbi96K1TVSskwB3DFam6h77vKNrPhlNSNpY0zYBT
PwQbsv8qEQT6Zva40occ8sGmpY6mwAVa8IIRfclX+1Kh4I6WQNYH2HoqcQOR
GCp5Hl193vkkYTECfKVEbCCcO7y6a69Nwy3S1D59ydeuZ+bmt6Z6zrMsUspz
lAqDTgvt+aGqmd2Y+BU20x6TUqGqh673TGVy3sKMmJ32FexcLRvCkjk8sNgA
BMS4B76dmT+7J1B+ZYHJMkUlb5zRvXcP0HtnU3FqPDUjy8Ar4kEOTNJ0xYVN
mZN/emK8lBs7tCeeqbensqettAC5NohMXCBpVJYzwNE1o7uW5bj3sWEOpAsG
tHBydQXBZ4MHT5r3v+/u7HDQJJH0ddQFBbD0QZdeMZLWGmrdf47GEIyHLc2n
Yv0dZ1r38fGYyw856QmQtOW3o2NK+Yo5hmsGW7y2FxMLYN7vrrgRui4LmtPA
ULxl56EURRw+8KttVOjW8hrXk+UG7awBSLvk844DTRyxyZ2M1gMgc7fPL3a5
mvg932oyzMrlQS1Tyg9I1qSeRpcCxtu8j1mESzbFEsUkBzY55rxP82p1f2zt
ka1w2yV7r/fnbghJvGWeXTMW989txeWmFXd6+DH4VKyHLCsMKVUqeP1plEKW
UzF2XZldFo+GqMeTPP0bfqi9BTN2AxViNEuvLXoUkwKFA9LHsveP8vBxHKC7
aJnqETXOMikBHfv51LYjxEg6U+6Wo+ROTk6DuP/0P4O+XTwO3ZXJqbHCFvN8
b6Jr8ZUoTGE7f/IdRQJXpu7pEwUp+N0vqV3NiqWMqvEoEZSwJefUFy17I5Gc
D3mAgQZ5CCS07Bnt9nCNbC1BLYHfKYYKYK29V5ZC2gLarlmVg6y2ht2ANA3+
VhgFaTiZyG4NhMLOZ9VFO9wZYawBQIXj6mfkdYioX6FCVW0RTYDjczxdjYkF
anZPwkl6J9MMGBugVqQcyVaod+/PpNWNLIBwq/jyqCGbDTF3N+z8meenCuuK
cP4mHWxltjAHlGPdFOc1Ol6xD5p7nPhevonsRtFbcShkWnQxRCi52mFA35Qx
SfcMMTTrvBshPv/RAiEbQ55ZQUF8fTCrV9TKmUCUiLt5dPtSZP5KwVXnY1hJ
zjRQ/wmczB4vYlYgN15OAfQOhBCt/Rsdk63IaZGFZXKDzBgrSLQCVmbxGf1C
jKADz1jkf6q/JsYsvRXzswWf0vJlYnmB2lUGycjajPYTAqu4cpXPVJHM6m91
/ljEwkkSFrS8x0jeMNSKYtCDCAHbYm8y9VnSubAhDs4rTxUeOC2mhHUquuYX
Z34Cr8tpINJN8X4KIAkhtjoP5hDSwmPaXbvOCTfMPEHZ/Gduov9v7BFmGA+s
3g2fiWWMJ7uyDIUjFaAQwHMSixDpx0i9yM6tvaAhfpzSe3DhYHjQlbCOsCU4
dzzRN5BjmCGCWUbrNSJSkfmQ4fdkgQ9qZZPIKIJH2q731sTdCMF8Jg1GFEcI
Nblv0tNgEOKeY5j2GeTeFmcXZ5u6D7IMPNjUiGX23SA8WVAubysySagFtBm+
Iw35G+DgXpK5wttoJUmnkRdjEnEF0arj2mc0NB8lyDnQps9imuJzik6kY+wd
Bc62AvU/aKb6quXoTaOPAcqQjnbNAC+Tz17GvG6IBxiohoC92AhTtBGGTs19
aOYWOhfOTqCp87JJqHNYg/3lb0guf3038kUS5FRhG9Z1WTLIDlBhpgxSSqCC
hVoXdsKpZ0bYMNVmdk/801GJQ5TBWObcmIlnaX+b4PYcK6hcl37gz+RoFo1J
fdOc6T2C1O1SdMULavPxAVjnLbxTQDLWlmV0KmrU830b2zjITr/+tmHxnmie
xVXsl+JafJvLtHGem/7jhJIPTMDLRLA5ONaidUwYSXdBCaZA0B+uar6rYa8N
EZfmJN1vKDxK5tENRJSV83YvolnuMvUcDDI8LiBQO5sBBYIX1gaeqUHiOZ1V
uHravlSSPg5IahnWq7Pd74OLeNxOD0VHl96/bFpJ/hU1v2cruwk68lbaOxBJ
dHwg8xqDW9KLsnq7tk4sKh5JOx/V2hlb5G4zQfV21pciZ14HEmsAOiItmGai
Ijyv59yx/rdCAUbVSW+V3AqD1DtMVsq3htXYiAu8+vgC2/jsSyeGSx4EuXXJ
48t9HtO6oZ3/sqFUoNtEELH01j/NBhLuoqxRMpA4bP4qrkgnaMaoVOnB90+o
iR+L0zzQxXqADKZSMlyfv31zgChJwLCgz29LcLswb+GnJ36ic+e+OMKTAFEs
yJjh07Wa376/fgq97iCXsjS/QWrqvqCNSjIAhyCbrmcbws9SFTDs86m9vSOk
VU9qYkqZqun7LEjqLYRMdcPnSvkb6Chopw82OtsTyZOaSi9YgHpSmAlGknZJ
QTEdfGT5XCRIIWTZilE+XDgEfKyqWsQmqDi8pqd0DsQPADOoFjUxllqfzxe3
tl42ZBZpZwHJnvkBRUEzgVmpYRxAF7C5RMUVsrq9DkcxJrGYFRm8jGCOp8cK
xu/CIlEr8W93aaVbxC6nFTFbwuskW1kKLxXJ7LtiLyF4vmgBpoIbT6NTKKsT
SJ/GU4HedKi2jW3e5uT8I7/IpdRp2kXsC316juwR4KS1gZCysBlroytfrkc9
QClipuoZ7FhYSy00ty7Sf5TAo6OMhn+Iks6p5aO1f4VDADOxzIplq0N1amxT
MIdLQ/7SGDrPjRLvFt2D6agu6iNf4bZv4Td+bueWlVj7Z5RqwGyr1Ol3vdBH
04t8uCvyPpEETOQ1aeDDUQIwg+1Gh6Y7ylPoD8rwTqeX9AxenXOTlCZxFxC3
+siNOKcHw2Zu8SeZ9ZKkR7cIloD9SpHcZ+OqbZaDEsxgudxRx4rY4CP0QD9l
wJRnDq1F1/Z+Aqve5a2rnE4fubkAgMWXs8Hp39qaQhy0ZWRJR9ccvmlFrlR/
XDmSlSRfDCVby9TCAToe7rcZ9uyA4tMHETTwHKl4+s4Hf5s6U49wdEWH7mTy
550XE/1mOdR2feep+f/FUT1Zw3FIpX81+NbPr5TzyJCciuSsMHF8K2OrTSCV
QWdWRqjKqUiidjTPK2OKJPoxEtftrMmxHweiOSHN/TqGWGEu4caCe1OsoplY
xETf4hjxrT+GBQDtymy4XZsbWexIK5tvsWz1xtQ+Q0xTkY+5jbD4ENGUA1SA
wslYfiw87IysUuXzoVu9Iqi4FdhhvEZHLFXHslw83TCZOoFJ5QvRaLx53+w4
wh88AcplfDQ3tHfc0lIkZZC6j2z4Z+XU2BnotACPDJiVlDvmQllQcjm5once
/pKgyJpLnNOmZk2I4k6hW13nT+RwBWHNks9xSW4u9XsLTtsGaUbpYcTvnjn6
lngVD8K5PSCDK9OHViBTeW/JVHslkTtOq7BUd5uiUry7Ddyh5kigF9NaPHhP
JNSis7fsFfxfoM1o9W7+yOOxRlqMZT4FcDNcapdS8dDeoHPL1rc3d0v2W8t+
+Pf1nJ8PQFN++IXhwNpfKk4/dMNubDHCx0gnVQzaWux6hKYIY0JvI1pGcCWg
ET1qD8mHXmJQQo2RgLQnGbEdSj5XOk2OuuVQ+Y0+v5CqXvlV2PkFXAptOqTc
3Bv4c53i8Um8enazW+7kOnxVa5blFSQHjsDu29/WQfkXNT1OE0v5jTzQpe5j
hOOn34t9XZu+fq+LaE3HbA4sQiLhKCWQ7cD+GfLHRH2MOC2uj/If5yfrC8ID
cvpt4D3zzt09XEGybLm16XFZdDY4erCS1YE0zUaatgH7O2RsiPVYdBNi2rHf
03152Zpk1H5PQ29zvuRpvqEyQWgzcTg+p0fCx25XRs/U1C4/dNhGOdXi065Q
Tf8oCrFk0GsKALQI7/eYlLmsPiJk0wkw73RuWY/nZNR5R6Bm4vYg/QwCkzTn
cqEegBI0ySndFOxJFf4TJCdBnjcaqRwUpfManE+I0ssEycYVC7TXLKvdZ2ME
hnTMpjo4a3RpYr0UlK4TqEuUXLTo2u6/8uCvYMy2aiVr79X1PwcEWVuiAbnz
+yTHVdyW7LCCHp93MnyeIIsZJ+YI4E7xGIZ4w7zAXadqWwR5yNIq/KKfN54D
YHtaeh5mdOykImyM5H/nrhUipZmaq2shvDEhaO7VFbBoY06INHFsmMpxl1tK
qXONwKFglY994d1LYXLm6fdP20ZIoYJERO9BK3I48vmuPBYtRZ/DQHJ3suyD
f466xUcLiBgm1VIGFuTr+yIlI8W5wlKO7tkFDkIiWXKOhrE2n2rxN9hv+w1C
lblE+gxAfGYfFWcc0VrU8XzxAnM2iSG+uiqu2E9tYr2vspLJj7EoCFWUfkcI
jKSi3ufQnRgQHVmdeN0iYvx25S50KmuI3DKHHfIbqVIxIFq/L3Nd0+dTUCyD
AXGMi1C8UZ5C75Oaxtob9p/ljV4k0Owe9xPViAFSgibAdD08LTQMZbnwk+G2
W3MlbRjkZ3313Gme8Hkp3+DZYph9WnSsKUx7H025BKMJKqjSi6BG2rVrmU2O
AT1O4p9uPMwbwrWLPdSL7Kc5ypy10knOf5I1zFBGjmy2C1afIsJ7TxYhkJmw
fjnjycPPsPIl1w8DfmLOFRPTxvb7NNLshNY6WId0lvHxA8ulpHb+dv3y/IBC
VjEEoOGqQLJqrcV91uFMhABx5Sed3kjXhQgl9KkygHE8/9lA1kpMMTcQWeG/
ReguzKLYoUKVLnXRBdzE9r3vK0egZPBTtMGUO81yY0sCoPSKxCgyVMPMvnCx
PO4SLc9SkOtPdCRElAWO092bsvkkmeFMcRizCP0C1kZLIa1EM0uZr57JkaFB
QIu6dkCKP8hcy9nQk49cJK5weqSUxv/5oMSzRhSNFxIsBOlSlYXAVxsQHugt
rZIpicCC4Exh75PAbY9MWv/hWYQbda7NhRjisbbHDf6Xh6LF1tSNSLmpaqT5
vqChDMMgAl+DWZh2JlNDp7SplB97pXcdr1M1+SJzWT0TbA1JtOyjSDVU/HB8
SeGBNGjZdOGoC9hXhAnAHF/AjNB70qJvZkDKmCw53ogJbIdTiREmP3ZvDWBh
YJWg9QIoQLeTyCGgiqAmCB0ikZjjAuPZrBpBFa4zygnGEoAZNSa6RHzjHiJF
sxKPp7hMbdi08USPBK1QBGakzm/B22dBEIWv9oHR/00rRPRuwCh3cmNjVK5X
PInpcQIoBMxwZ8U8dldKsmXOrQDebUNZAbOUocOYXNs/3LDWP2ncaQeu8W7Y
cgRoqIT/fIP9it8+UuBpRntEHL9yNKJW+eDATcU9i4/UvK85A0QXf08GSZGM
UekrQeB8WCxQm1Jaomr6GYNnJTxaATHKvG+60P1AkOUcJqjxJuZ5E3FKACDP
MIUdkByiALUcshyDWg5ZMfScvgr9p7KQtdzJKH24jO84IwFRshXLKkdzYhmy
yYg1rTYXzMx9rJ+wO1jzg/6zGaC3jE+fulYJhokm5Hhkn0s5ULV75qLXc9wP
KooCrUvR0oEmn1nDonZu5yfxsqQEHopH6IEHTEidpTphG/dGzPfz/pawYmGf
IchcK3g8cnsAODUU3WiTUYgel65MlXEUQXFwgvueil/uOX57HkS8vgwi7pOI
Z9OM9tavKs5/lk6h+H4DbrOlT6gGyEMqArZe0F7iqD3ifIRW2DF7ZxeRyk5W
4kpMCAYIfgoBRl62HNEfUJDSXLeOsA+5M85y/RsgHqw0sTWencUdpxV0C06v
/L0SS/eyd/+1eZ0nEu/WhBqxbykzxT+dniRishUl6iLVovHHUKIsIrbum/EP
yho5ptvt6K+mbVR1XXuUtqM9gnFDKLfV3EsMMuxxKXubWRmLG3gLvuFeGg/o
YIqRJwx7wX3ADBuLIk3OxbQq/pHMXpjveRuWhe4FsfMo/Te0oPg5YpGT1nWR
3GbNEcIxUmfD7kH7C8c+xLfOGdvlzbAKvosRgKlOnbbuMMHC9kqN1xtSlHVu
vFb7Rd6mGKKHXRDIVR53W9JIWR1pEuwl7X2gAGNazhB2Pu1SI9EPijzCO1Ve
yg5QC8ZZBddlnBv1FAZUHx3jcZb3h+EtNIxj4n46Svgj4fXloD/paOsNi5TO
cmPUeSP3C19GmJEQUYrrII2T6Sxu8ZWB4L95m+dmztBGVcuUhj9YHTnxc7Dr
rCbUuRnjfu6tISrNR7TcM8zaUTuK28yl1k7DPaXX4MravB/ro/Mzi9YhGz+h
hLxVZtrRrotE5LR8vRiUOAPB4DCwzP0gPqy4lJAzh60HheU3MDeKBopg/YEP
+vuRTVcQbsudv056+PZbz9cklfGZG8JOGPiybYITqijjPWemrj2nlsoa1EEM
6d6Fyx5ZRSfz51GzA4vfyKk0FGxjoGuo/rpawKsS+u3VnjOgGA98CIQu6358
2qDH9abPHwwpiMSF9v9ku0O5HY5MCAgge5vE/GxRPA7cJhZslkaztfxuWL/A
J1JoUHqvuIO66cX7M+8zPYi81lH7kPfEyHLwPK8U/+cd2GlJCok5/yjpIgr1
Jlt0Vfu4MLV1Bbljkh1VS7ihi4D00Jc6vAbLecp/IWsTg9nmN1yIzzSgrRnz
nU9iqgC51hXWL2lw03ans/0cX4eIMjkKcaZjG56td3zcoXV5/6IwjtkkCBu5
LfElelF5J5ZDyaxrk7jhzaRsopvFAlraP9YIlhmRA0yvof/Qi7CBGH9n4TCA
rkjN9MVH1YDcgMb+F9Ghc4PHlzY5cfk45fgnwvhUWEpI2RRzQOKBLo8lRooo
HGiF0ZsnyI6IGR4klVmpvwfOln44O0eT+EZRMgKD2TV4i/dR5G6mESfVZ7ii
oUGmDKPtOWM/MCDK7MiHXA5REIrBzAoLYA/VxP/BWJOfCnhc/LrSqMECVB4R
kg5frkBzK9lxTc5tJBaoiLfdj520GmzcdmzW4VG+j3lGPc/cJ0F8BqkYo4AO
ip7sj18vRwHQzynMIk6SCJNGuoa0V4pOwcIKdep2kqEWMnruaFE/zhk2lhuy
Ms9KIudIKCv+9PwZrZS2qXAMneoXS5ldD+TBtEUg5bTzGy+5PcA/hNUWR3fp
9Z+8Ckp4YA1617+F84fheuFiwIIIm7FrV+gkl3Mc2ovKiGUfcEhlnpzc1JeU
LXB19qbhL548l6h4bfEC6G+hj4eBzSKvNYlw4mjoZaPXk2QkRz6OFs8GZUxL
v5BQxM3GJmH+/iX7v8uVeQ5cgSq0pLHEYh8Jr88IaaT8Dzn7zLQl1aYs33TY
2qBCyr9+zUR7lgjHhWgU3Ug55pDNtxmtcLFiCfCCCWwvGpXn1Pd37nckXGgw
zMoR0PNPybaU4L5JKnCUyO6j1K+SNF0ZYh7rOpSt7BFKEWKidkDjD8JWNT8n
kMsw6gqWu0Ft4Ar/7yNLh3FizvpoUOR4N3uAQFVLWVGySms3jMQ8lOvIBC1k
Yf1depE12aQiO0QcvQ12gaJcopx2fcL5lbmrBxDztTmVWh1GPAogWQzcMETN
1KZ78SNrv19jhDuBk2qE+WMDqk/dYKyUiaiKPdfHrEc4T1YGGWm81N81bB6O
Emo6t45i3jKK9NMI2BCg/JalTRymDzNsr9wLmva2djfgAr1xVuj3dGP8aJnK
2CohkVmM65rNKcVj2PM8qVRElYYE4/VfqR+DdiWEMvGHohibw8aMVYiMbW2l
znTsR0Bk4P2Xxi+nBExy6PLVqhUOtzxz8qObodS6MncTT12JmY7JYRg0mBQQ
9z3q3pBmQ38qlkDTSkOBae3I7zFuiiwvBdrxCFo5jS/XI1DeOXMY5jiUn/kb
NkwbjtPr7koUehG6T5lIYEe/rGE85sx3EhU/A7w9CIl8LEEViirVvkkewVeV
tMzZUOfheV9TzyQozpvCT3V58r+X7oajeuSK6lYOCUs/a0GMsnS2+xsMOWTT
9PNtB/YJuA79pO/iQK1O4WLRzccAxrK3wEjUjo3PIEQtvKQ4XinF0ncgLzx7
/3pnkUYP8DQvLqRrdReJSwYgVCqDRZ0khLgYzzM1DxZQCC8xW8KEv7A46wjp
pYfYKHP7Ay0neOT3SYOENJ4y02dPJjP+WfnAo6Cx7nHXgPLmuTtZlZeHVU7Z
gQXTcNuaLeIMY1c67fngzjXcKCIZfuZh2cuiKMqoWzvCcav/QSx1q3NlE0JH
kxQ3DMkJu6JaTiO40U2A9hftKJG1CObLhbpKWKwq3kS2vPJz2VsGDw9cpBTV
D1f2sriR/kJYlqGJL8Z/sC+i6EdOS+Mbn9gAo5OTLgde9i8f+NuJ2bfuf95i
u7n2BnijbFs2LfcYjWYLnXMJ69oy8qayoaowmbpL+kqYcKokJBz3wCu4JNMq
e2LOVFEQKKnHOtSY0BMmjOYjPKbHdyTyUmmqUigSOeSxQjMOHIzgvExEbyZ5
3NlwEIEfCwi5m8kyp8WmbOR0XfjbQnMxdduhMsMwkn0KbDXOZ+E76fPT5M+n
xEnmfmHYEz677zBZDI7SaenUCpxcMzh1nY7UnN2YAJKFVQvLasUKS2a+hqDM
T8qk28eEorSxdWqD7QJvaO9o7f+LSQHAqS7kP7lYfRP0pzyjgyH3GQEzTU4V
+y2BH3CPkJtW/CdOPOntBvhZc5cmTkkLCXzsi8C5VsGnOwHQFdaurTXPbZAa
HYoh60SNnaMyDWAbSXh5RTrHXaW3t1J/abCCuUORJgfnC5DJ9sCJDumW2VH7
v9znlJDxfxFYNotgO6euWbQBcBfRl0HYNWXHpTsiLO9C6eIrgiVUapullePS
NkogZljBrooGVr+M9ENopZHgG/sxIsv/HFURSC3UTOKh4R/3cQCj+XFnt3cs
T8AtFqqThXzpA1hXSRiIYEXjvjwyZKqd/4UYGup23gKze8RnapgcAdMeh7lM
EcARdN3To0vum+QIlSbIVnzkbsc36hUGIek7xSQyWPw02eMP1b1+wXl5T9Nq
QTpe0gktgz7ujPlukJAe1AkGGRzXyY+K1zmFncjtz6znCJ0rNmLfYlXvRBB1
7NZT0nRUQrpJSRmrmUVfegwjBPmfZXyXGy5kSOH3leJFlT6+NW03COJZl14d
pFzKoEkg99T0RCYya/wk/rWirq6QL20IJ+jvAY2lJOYsWm5kAQQ9nmtjRFE1
JcIOthtnp3Sol8REc7e1+BPwmS4+fvnedIuWhGpR5aOHQ4UXWE2/vogsyxkX
EropBPAwwyZ1rr7Au1dIaiHXOgorXe4vD+QxT9DTs/02EpCoE/FDMD9M+0+l
HCLxECHEB6WxeY+d0OVV3yihZ9OogCfM98zM8Sh9OGgRtSNIVUkFxMsmmWGY
0ITa+E8eX/CReJnbY3fijwyn+oPIVVWtk7jTUSC6uQTZkr4Yy1w1zBUR7NFv
A4aLN0GtvNlfX2TqI2aY7OBDlG4QAPsWGyASQcOu6wbaH9N5iSkxs1hYYI4E
LnWdRQ87z1Mi+pcbgdZAYGXvGff0ExCEudoq+4RjCmZsj+62pbPo1Vi8Ss6r
nd95htSKI9YvftI+ytijTbJOhoxQYn8vDcjFMC90m4uNf5Hj39rDGvdv2URe
FI+SAS4yB7hToxCnlEtClo2K/6NZL0UtaaHkIhPNqrut8FT/2ApVpzAWfU5p
LIGNeFchI8cNTuEMxLsVLixkvHzkjCzG4XMZe9t7NT9tetuA4THcUj1/5U+H
zo9OTW0eihg9Zt6It3pUvsmvgOSQCKPUcAII/j/++YU7rm7IsmkP032GafLU
Lf211wJGKSxTrttPLxjjlRP1nIRi29lgrIi807g9AiPUjtf+II3PPcWZLVIe
UPw9poV/wlEnIGsk5kgYTRwdggKXKTstMJfLLSLETJf+6Ad34H+drSm71/pO
basNfR4T4F04mgKJF1C6eA2MCj8nrfzaFEDdGJOUl88NwWPAtdqmJSxn8hYE
kiGSGCSnYHl6DKrWbs3io7w5pE+ymnqAQ0s5lqiVfZrA7AjJE/BifBy6aN2i
JnwakIrh9fb5IWTdc8zX0Uwdt6VDFo0y8VqgLXDrDRj/FlWqbL/WeQ3SfN/G
npAdYqJy6kedGSsu7dul+Mb7csQ6IA2uSrLN8iBAk1FgECHs0I3y1DP3ogxY
+cl0FygSAvxGYCycp/0STQ/eokHIaXBXKUTa2vmsHk/trd4kFB7Sld5sZSk4
XAVSSspPDnI2pgGsdouHt/Y8EN6bLPOZ7tdWsHJ9BMZWbX8FzZYhnHEgszdT
6NLBV/579ZZAxs9k7Z+mEh1JaSOCnj33t3KjHjfeE4y7ah7Iz3Lm6T2s7kiO
qfBdxTut4In3knoqWi/YslidmUKP+C21E8uLHaFZQ7ysI6KlnuD1272vc5kK
iigyMRUGywyPOYAk0g66TooXPMNTk3vashD5w6FgSqUWSi1H5Sq8kxUAd/So
v9BiQZm9d+qUI6NL/xpUCo0rN0vHLjJ+fYinJ1GiL8YGIHRul65UQC3xntGA
BUkKNVZqUyP2oETyd2EaNy0zbextKAl72odeOC013vcgfvV7C3jvuhcg/Lou
0GHGo/XT2K9yk4PUL5Ez+8TYumr2E9bFqPinpx+J49CQXsEx5pgRFPRIRffk
UpQLYzQWuF+7liHI6Y5ZSFExSPQlvNA2bs6ApgFo37OSZyemTLwS3lEhaF26
aSgokykkyLjsYK4mEnPn6xln25z8uS9Wi5L7cFC6TMhmqiDX/xSwCUdvlMty
U4oR9NErRLV7frRHIT+VW8Q33m/iSkVwKN3bXTcebz+37RX9uoFwl07i82EZ
gKV3rOLxU9k30GZo2m44tYZsT7w95S8JTggY5Vt1qjtWR35Z7qGFWaGbAk/4
LPBwcOBKqraoXMZrr0wqc9LCvt8lgtu1tWBAYQml7905oF4ivW6wRUEAK3vW
93pAQKsSFXBjEVus0bi9yWik55ns1U84+ofMc4Hjv/+Vcjag7CUKn/5z11dc
eRL4Rc4NbiHsjwWtQz5tFZ7y1SlMGuWvjhoQXENGHbKtve6mf4YyPkZE9o+d
ljWLHag1saD8TODYQaQ6IXTCpWzZFoF1sD4ksJPQpvjRr1c3d5K2I8g6E1J1
S88qqQZZe+n5kGeOUZuBn1utDNBerNkRnCq7hcbTU2QMEDQskkjTQWf2nH+I
br2wHShRLHNkGIMda+7pYudiuShn/fIoBtNQ+0sUiTeRY8Jx+ZYfzCE3+YAQ
FF0Zntwo0nWYesHV75T8wkSiUQ6rjA6e5r5i6rtSzecbaCm3biQYGObzH6Tg
56CKERKL+Vg/B/LRuBoxYAa6NYUJcpDZDWeoQA6v55I76W8uexGQOffMRPJq
0ay21JZc6NBIEcrY4XRLUP40wA0CNdlX35ci7Cc5GEP0PLmkZPWbI0bXNqtd
mOhOQ5PDTwsPwZsbtgX38PR2kN2RrbUr9g29hwNZV1ZMELx4yP0B2SAs2PVJ
7Z437kSmZ0aPXvcjO017Ytim21UKl0boM2GTsbozLqeAiN5XaRbUUY3aWZ/e
9wi6cXhyqc5Nwu2WCStgFb83VEhmGAz5NEWrgNhi7IQ+bPfTa2IGFA8aR6wM
987gVn2bwoOyKGO5qqX+rRoZ5ntuaNvQzORfoP9GGXrUcr5LIDEIP8mZA0wJ
8rOOA/gzrc0bNENlslB0MQLxx+QqaEE4sqXPKpkVFlnYqcFiT0/RCWiJtNm/
g0JWX1V6Qxcum8TZbQwctTGhEBQa6N+DKiRy6BVTYLOyvjVzgaYrQoQ9NLuk
qWZLSJL+LgNFa2T+1bIv3RWWTRlN02Yr71AJ8nvmI9rg3XD764EDFbK//wLY
NeCKtMkiGEbdffQJontXrF5n6wHafr6Uu3Ge+16qJkjgRnOUenWj22sqvmMS
alk20/6xonisqN1yQzrAXoamEzJA67IBb/zthW3aV4zH9rMLOJDK0f5Es84p
73Wdc2g85oIkfsvgQsQHjnpc+i70BccoS/wpYXtl7WVzKwwzrc12+mU31RKW
dHCNxbd4i5zaymJYcDrNuSgACHfyA2BE4kS4qoPofFwwSnvcdCwJbFFhjq8B
5SNB8ihebS4RUukyZZl2doBNopYWkQO9qdtMmjKYxytPe4gh0YYgTk1KMvVC
7YkuaikA7kqHhwJwBoI/lZZn05ugLgjDN00B61kxgdQVYKxj0BfIpaNSMB2Q
PFXzgE+0ku6AEZFjJDjLBYy+QwOFKu9ExpOL8AIqHr7aQcPR63F+KMsM0tIQ
P0qapVgsIr0ZcMQTiV7atLGOxuyY+EHGRGgE0MekKNf73mALzeczoSsAK9b0
YvUrmJdln/L2lX83PBXi4IhPJgX6rvDTdRrnjlX+/llRFb7hxfaw5RoCCN4C
o61a7ZWaVJULCvuqh1MJPKT93AKBhzFkTUeQz/ZPkdxzPsveRXxeSMk9fmX6
qfGUhdEnSihObHP70aCL5PQne9v46kkLUOwGyah5oYsmssDH/WrqKtLL/Ac9
b0Hskp3PNKSYhyabZzSz5mHWL1AQqGLtv6kdR7+VP/ghXc4pX+uMOATTq/tk
vOhg6mcKZmfhvU0MP92XA7f0tlQKvIKpvc/PFMB3JDftg6V35p+GuMjvhdaY
WgtPBqQMJuDaV8RSuQH11GKniuWlpN4aP8LCiWaOjhrAOw7JHlV6DzEhn6OO
4XiPGkCGeRlcnPJYQ3uwWnpw8DfKUtxHSMYgosR/ThkUzfPN5n7ER/LG9hLy
CttaPz1LyN1QUlhTZkuwbMTwYD4gHbfl7fXYHTq5fixd/31boIMpJShHA8PJ
SbaAimCaWIrUm6iUl2Ideh+zxCjpc0+3gadXoWBJbOJZf7WmnlJ8vz3tcBuw
rseJGnqnT6qUMaIPvP7zmB1fY7w4o7LzEPP1Ec50luzoIOhnRE1mVlv621ON
s3/+dbglNf9g7ew10yP6V+worlbZ2s5QsJINorFVKnbZ8EzYoW+aE4oRiWpP
Q406oz6pE76Om4TKTKSFD+zbsD784HFchQ2+sZOGORB9pA45hZvpFD/8diFY
LFTCmaGOcsvQHOBes3geSVbb+k1F8RMDLTLOsZMCVlRMfelvGJSERLPpajxs
H27TKT2uEMMBi6dnGAWco4TWpsV8jlKq0P55IxhhTOchrqTkDRuTjz2LZS3+
77mPb7UeRH760XKTXjy1+Okeg+mtS9rlAI7qGcVeLIlkCMjXZU8pg1/4ra8A
t+cN4QpC743qO8v8giu6s5wvLU3mB45meMWQHpQYYr6yLGsB9qoODosRn9Kn
J9R2q+bk88eem1t5nyrnEm+XRaeUwXaOZTXWYlgrcxFUoxN3szTvSRduMYV6
DBtF9RX7JQ0Gp7n/Qaux3xwxoeenTvexh4lBeRpvjSqPey4o600HSyp4BAUs
lARiWEnw+MvEEwREWEQC94sQirPfr8yIPzHgpCefSHpKc8MYANrHwfof8Xoq
z453ZXVfl1OYm84Pc3ue9QmMGs0MJkhc8BeecFee9IFwg+oEYs4PnYXcvEF/
/BACG9iV8p4dpEzGLeSCGnJzXJIT7zHjGa9zPta+h7YBZYbsGAy66iO25KzL
vx49UOApdXyJLTTYikpP/zuNEOtP5nooRkFQmubweP3DnKPHABHkAN7eRyg2
++68RMY8Ou8dp2WiBeFEBuG4s8oxVF3HMuHh35SeY8iM60K44+AWq7S3kTyn
+kHCwpGEVf9BIUYzqC2qoyyTZlDNor+3O2ilE8cg2yDKB4PxqSGQMIWLpbEM
NHrC/TJq/EY/Z1z2tLX+ndAbfwQnqZHKRzhdBmJ5/czcyEQTHFMHtFfX3X09
1xKGB/EG7Oy2Kg8Wr9RFM7D4QnXYMYiZXW8V+qYJ6x58IN5rizKon2zFe1St
cYm40Ttt+njCccHlH1ZSCnjFdzRcO4FVWCVU0uP1jZre/WzinrBueaVh/oAv
vpYVqjRTgGq9XSiHHqrDN/Z8/8lCY506Rxk0cgb64oPLyIkPbrKeYdFGJWAl
5KQkJ5Q/gczlxfoz7nzVpUNXMq4R5ki81nNgVFMqfL4KRbppVJcBf8WQBmZA
jIIgsHCyra8V294Q7Ln5buGlJ3m+CBreIPiTKb5AV6gW7WjrCniFJTyBByP2
u+UWNK5lRUItxa8Wa+IlgO2tkqF9W6GPZE4VF76jQPR929wT5qXat4aDywYZ
G4/X7mxPbuSZMwW1XAajkRDW4LmrZHiXm0/Vrvj43q8ascBhlCm9++dTY30H
gFFZmb2Pfgd3285QqZiKgjA9uvJWuOBKS3XdIpIXto7rzeTvQg3IDriW7/4X
+Kp5HKsBgSfMpiiF6g9tQPJivAXG3eLLVDPYSvaYEjKhVbVh/KkHHjC3TB5M
OfFHSX0sHqnnmsa9C2iMmKJzSn8j74NBYaDoo7XflMC3RfaC+IYkvZU1jG/1
ewsmPZeKsW9FwHUyCfBXAt2fBDPz6RzMbLOq47AzdKEpovEuyJo1QbBH9mp9
jubRPKEXagmBV343ale0BM2+ltpkz/7AuDxSGBg7kLc0GZbQz/lMuFj3QMvW
Aakcv1AtgXGbxaoQ5B9422e189V00OKeneFLvo7yJwPLSuWXs9RBlTzDf5vd
7bzzK6kJMaeSiG5aMAAcCxwaaNwz6Zwy9UKOHM51KWxqtyLSXnf7+6zPbozi
3g9OCCVNhM2dmpsxM4A91HUuzAPRUEyk/VAAdiGIiOh57/9Ixst8iOnsTTWL
6r66UmSPTo0WXNWB8/Zydite3K/zdnYBzXgdUMZjx6xROpfEiLXNtpsHDLD1
vscWpKYF48Qv83uEMjwpPL5ppS0ugHcI6tuGxQXJ5Cffarx4Q17REj2xKfQ9
RFH6PAyFCzF8TkbVpTIbLX8rupSENCzF8ba/r/lCwopcXtvZqmozc/EftWMJ
2LjVzeD+drh1ewO7sGyaJa7PNy0DhcByptwmv4NwHJV3xy+OZTH7b+Xd4JQz
tI8FeRMJb+LrU0cDoiGaSvNtiKNmAt1STiJeIgntFISbMegdgu1LwTZAWA9h
MeRLp2A+cA6m1FBKjGbGH/mQg1mnaSE+XQNRNE3eFdzxxDtAb4oFAf6jggQV
g8YLvRsXZi+rE2UCqdxMZMEj6qh7An0iRmJYWsFRApF2thsX3wsqL7UDHvim
10a0eaRhBmlfCJLnioCoRRdnUBIgRc5cGcvFcM7ijE9cuSO5+DmTXLl1+2rE
taTDWFnY21zPjkaHUBYCCjyN6yI2eReg7xqeNCBxfTKOzUWWqdWdN9bvUkEO
EXrZYmQ0ou4C4CfEznRyB8diX1zt6+iQkZWe1fGaq1YAC/Vl1ss4R2vefDEC
5fqv2s5xH8pYuFuwrciwtYOm9Qn+O0mYVo42xxX3cNBTs6K5Ge5zwSwAxzO5
Id1qKpyy0y0IsueMuBowAPkIQtN0FSr+d3sG+E1uYKOfcEABGpT4n8yG4CNX
SLiiBamtjEk+J5YYB1tj2jvtnRi1H8g+FDuWpPx7FxyZTPtcW1tpWw8Vvl+C
I1fOFu+FuO+kF+o3oaSkowlCo91fwtnQaSMgR2xdFzllx0sdnyzd9ZS2UZ79
B7/RRiDpHCPqPPKHl3RTewvkbJRAvsDBFXqNzziQpi+/TnvNiyYdvyqRHdTl
ZAirefhqf//NsSfdEMUrzXZFDAXo5Z3PWifZ5NWdIBdr820icvQEofgG2liZ
bC+kC4baQQPz8+9z7ZRTN2mHjjAIqfyc7tvoK07Kr9JYIIoBmYykzlyXDZSs
r3HLTCb87qbSkJvrXpevvPAG6kdbs6KEXOsVPVGEBXESWjloq8J5Thr513em
ValebbUBYfOUVtGbYtRHUBEh9bZwWSbJqSPnG7WEgrMwP3JOpSZbDq4pCKNS
A9vMdejKJXg1ayWvUaxfbqxbPxskgoJKycxftYmC/JajeUVxkeTn3K/iQDJr
2ErKpVoZEnxkjRYr1J5piG88RB7qp6ExPWggyQFQFTDRS6MUgR38zmMcTWl6
tisr7+I3Z1eX5cxrJylHTX5pBPOS5MMYm17HFIo5xmvazAC/8V8YEhFbFlE7
m5Mg+2Xbs34yncRRKPRO734ty+my4WfgA4jAsVUnVK28VX7LakRAGgFIXEgB
0sPid4VaiJm2bqXlm/aStNcNv0Yw6Pgfk74KhdVhbq3S5a7kDRYHd3fepyDK
Y6u+hQmKIYZQEbDBodnmZHJV5pTm77GmehEYuDz9AmUWJga+8mWg21wpTQ3P
p+47+imcMtI+hV4bXabq/DWjkKFp83Z+NguTrGONuz0FdeDuyIymIQ4KcARs
6QtpK+2Zsdf3kHMgNGBzhKQDlx+2qFsH/ki5qKNY3mXkzJw3Oqc4jtx5V2uv
3Ro1I+uW3NIlbD6FuHNtM3hlWyok7cf+jTbEHDXbpAoMYDhFy9jQWJvdM5R4
6A4MX23/Y/8QkP7Yy/62XIrhtVewz8rx/HwI8J0jCF5EcEpamyC/jogoS0OJ
9Vv8nav+zgQJBP61A0Vxpi4hfh1RuqEcrt3WPkHxywe4AGNJ7NH5664cGmhu
/3z7WC98wpf539qovABowwv+kUF/LXN2xw9xAlYoPcpmqO/Dhme+cjFhjqHj
mIZlrXnI8r/96q26ZtVADlepP9JGrvt70xixXtd/mRdVYTg/y6bebfDw3GVs
w0/BCjMRvJrFb2JbGB/So6h0Gx0b/hA1eFTEJbdv515J3WQq4wsJK/5luk/g
Om2pkGS8uQL5/CO5NqufLEBhUWlXIVY+cOncGkSzjGe8SHBNnuv+Z0UyvEmr
roKCWjysDJkYNvuVdP5OZjJsH04oVzRCbKq3K0qZbIxxum/hThfsKhChEl5S
vngkjawvTThJr7d3w/tiTpu/wjDIws/QmpKI3nfUznvePmKLDiEnz8emabRm
WmqtXImi2V8u4fMNbjnRBWLyDkZyk6zteUn6cAT3FGlm23A/ozSzaFqJ9nQE
R+qhdffpQx9OSWwXovIk7V/zadM5PHQi1jmhAx52abaNghL3fOQaEjFNLSM0
6YIMOV5XwrhqAxK0VQYj0x5qnDh9OjxYWNXUHWUeGhYYmpfN2FA4eT50omO5
gRquGGXdMWX2WFDcNqMcEdm36bPF4xIRU615srDKj42wFVimNC6BKQ5c/ZiT
VazQyoTNJoRG6Q/RluHCx7cis/DCkLVlAkum/Go0E71guKK31TnWqrqJFgoI
hSnsrOysriNfj5pMEtyX2hdDGIOfo3LknK1rr5RAe2bRTdLQgteSopDGvzzc
tXw3hUSExGFB/0XPq3MTWXnMfu6Ydx2x24dQAP2BNTIG/r5sTlHQAMb0NFRd
QVbuu+FmQ+GhtJ2OALCRbRljNo+NkuFgaftBnVELATA4NdO0cxaf2t5pApPH
HasKbP32kjrw9y1SzEGgAxZoguY8pTtTZURaQYbRBxXF2YTA9mcD0hXSINMf
0OOkN4YlZ43DRcg8EN3cF8iqZMGq6ya73h4A9B+vm7ApINvhxkOWMTEU08CR
ksM74jETHSVFuQL+q71GxrdJovpVql9jmczYYNwE7F6CcavgOHH5iY765qJ5
loFT4oMGML6i5mPGvslHi7tdxy4WeKW7m2ZJh0Mc75fxmEuCH/rv+DG0mKIC
Told62qCDP+mz1uVexHabwJePNNX3mZT1P1IL+hAZ+avnumZqQ+62RJ7I8WZ
vXY9nCNuqkdHZ5uChX8OG9B5MMBBomNzgQicjGYak+HBNHT7djTNdliqIzog
xYhnu40XlajtOdU3IapniK/flJg94SNPBXaX0OkX4NbeKbvwUJrE+REd1ZSb
/Eg5k8he5KAo2L4KmZo7EKPOjL3u8l6ruaY3y5ApZbSoR3gSLtYnP+vHAs0K
hg5L48dGd5D3BgpsyzGxavFqEjVrvM3asKFnO757DA+0e/SRMgsINb4/sRnT
PKjNrEaN1Yd5hDpYwapt7tdd1zmzcjSKER1cQaURADXtARuIAQ9S/c+6GEw0
ZqrRwPKzjwBpyJdjHu8naBXnvqn/8govJhP0eDKwILwTF/Y6MrIfubmYT5Ac
FwrBk951+BuPXeiQU+/yabRD9x1bXPx2IqTVpHPlPjb0CKQUwLyLLe7h+fCG
8O8LV2SdFKKD4Q150Gs9cQDj6bUVvY93dUN4297x9t/z2jUfbl/TiUiT2xkb
E+xhMShAhiumu64JtwzDatPFw9Pjnce1b3PQaY5O325ELlqsFgyKNh7+d/P5
RUXG6nhZc5aHRqm+j8nGOWFT5i4Jf2FwlAvIPDCjcc9JmzEDYa/EbMlLvmfK
E1B+rY4hLou7zZP34688232TDLo5TwqrXGBQhTle8+r9G2VSpCInIrvOt3QP
ZD/4/cuLJ89dHXtP2A1wzU8UAL4bZTDfrS3Kzp2ZsKV8f20W5DBlAWrF69gg
bdGFhz/GzXa8M8I5rnMN789wq/mQkYpaQgYOPZ5eBhe8R/iuLC1Aq6pfzKAf
8T3PTjhyN0ZJ6ooJZMro0ggqFBl+pjykM8YidWOZyT7EPJz8DvgZhXT1Gniw
7ckPGuLWGg8vP431QvIkFA8tCuSpLTYPIBbvaePPKDqYmkgucKEpN/LHjCRW
XQJhDmv8rUnTFPpVOP/Cjck/FRqPEZhXiSykJnos2SIqJ42Wtb92ZezEPVRg
wgup1N2p1Z1DgAr9l690dzYZlu23Yl0BS68uZzteSvKC7GI+yShgHJzNgS/2
P5Uqs/i5MZAEvqgSX4bXk0Ba0boaPhtOWXkY7yUxPRBqemf31urg7lr+cwmw
6lRGhwsjQeqtfi+0vqV9rceJCWvOSBZZglDclZi2MsF9og9xwC4DjIkltrzF
vwU7T+LxOG2haLsOWJDo/zaT/Ei5zEuPP2+s2h2LKAv2RV9hvWL6iMUyTCmT
hSo3FaB7yYNfXKgMopRBjPDdm8FUTGwrMxrWC1wFgR43pCLpzgpFS3Na+yup
ApjVmmzTjE/v539WFUmPZ7mEca3ouIHdQro+R5UoJm3ayd9aXoLITVHPORSU
7V8Oik1qGa1gsfFFz7/IJNPUtvsle0+e4Qri7BICEuyWCRcPjZev2M0A5Ey6
owNOPuZqSxqsrL+S7DfQFltQUcvQb5UdCXU/UvY3zK7Rbb2zE2Qk1N9r0mpy
ov1zkeZLRoSw1M1z4mnrAy7e5JrMa4S8DR3INJISVeiINEfuKj77VPxlhES0
kq29GqRP/0sVAcHSESm2gZZhfZUhCdMMLrDW9uIwb3ehK/2ELmtrCK2gTb+Q
SAyhChmwTT2q3X45iXU0LOczIw9cmQX5Rq5dPZxz+UHGPe9sFDRpRoflvFrY
32VLmyCACTDuXrbBHmip+2MAYhkglnZvyrwAt/72pDqZ/WzsyWx6JrRe3+Ju
KDj3EwkzXq68z32FaSwTIBbh0dDnE6ITlyy5FQYyE4azuVQM4LKqC+ZNU8hp
bhE1lKoxePBIo0iy2x16oOLstKiQ+GASOXMFhumf751eANsQcJgEJiiLL9l7
wEdQX7ipeL9ffEW8huy7EVWlSs9vXggoHJZH8KIMo8Itks/TEka+mkccGr9w
plaYWuMqRewR5sfJlR9KaUtps6WDNe02SJUNN0/FYr+sAPeTQde6E6zLp0/L
az4DLUvdIyaA9/GiGVGAdPaQ9J4f0BE/aMRzNzACP6hkNNERsr8/Arh+FZ/s
OjlMKpPB3Dym8ly5N0SaJwgno4iMP2BTlubP1W0MEBQAVjGRT5o5651KmySo
JWYYnWtFxFQLGyz/7ZJiIC8cypbxLe75OGtM+Ig/i+X2fKvkD6D1RA8oGNSK
4B/1D/gwQWI7DGQ1+2jt5zhM2v9DrqeGERMum2hASN1AH23UjVo8XMir4Fv9
vW2YCCvuy4yIWzFtC75W0Ebpwnv9Mmqw2/6g5EaXWk3rVog1Gc3pkogn4rmZ
wc6rcTU8urZxyV5D2cCK5H/81CtPuzdb3G8JQnkSWyCLdsZEYh8jxnxr0qEe
v65roAKE6RCLiz5p2yLphJWZJapYplLlf29s73Fv5UtFCUJYvlEJ82qe5CTb
Ym5p0V5x9TBizY0xH5bEA+Mkkp+xWevGLinW3nrUX3QI5kV5rGnFpm23DUdL
qqsAfg0B4hs9mjckHtz9ZLavGZitaLB4s6RhU2pOE6/RvFe5seEBP/22wF/4
URz4z3jkJpolfRbGs+exEYQ0cl1vcTtea6E6+FI914xLpR3Aw+63r3cnbD/b
KBDTnwMEozOfNU+agI0jT3oghRzsEWFjCSVEy/7HqfYTrioL7TA1SGPUdqF9
Go+bKRVTeKRlr1yUOvwViv/jwG/yfiNEH6iO6XbtPqQCl31Ouub+6kUFjtJD
LXLSJ8PMZS8z7o4J08r+UKyKa5lt8rxxJgaenzQ83ZYcJAWNCQnVkj2LDEyw
zw3N4tTgPJv+pLo6UYfaKB9LWCtYM9WaKrh3xACTRlITmoCvuRTTP/wVaFyR
uPj3pWxflNFRTHcdy880iv3rw3GuPHrs7qkUdGt67yCYuqXixWSEns7rPHMT
IZC5rYBMxrVDU1yuiJZ0+LK5zZJWnSla2qkb1xtsiFTCtxz+oKY8R5nKVAk7
mjhn3WpjfO+H27fNKkn3CYVTbNhR9McYonCV1E6d+GNM/hho8HZxHhqARIrh
lpiO48vfDmf4JhEz661u9BXAn//uIQ+6dVT5TB0RAGB5ZM3irdXVHzEvfaWI
SXxSqo7FDnVKVo22xnGdP78jBHZbcajuSphM3TOHYHWUyKN6niqkqtckNghH
hjfLsl94Oowtts2u/j8HsZexwLe8w4JCcAjKEgAIfIDlpGVL5roFKuPORJ6d
Wb1qOPy2YMomfwXtoRfvb6Q+EJM2IJO1nrD+Q9fwRUfSmlhhPyyAYTa74CXN
pqaWZNUOPKrAXJXh6dBYqoz7sOS1MD5/AKwDoeIlMwZcgJJ96KuUCQZRP6kS
ycP1uKrxFtIQdrFLUJaKmsk2hpBIkmEz9+Wejxfh3aRcY8VgYVMUmUiYTYeg
wziop4zKtPE46lEP5H2WzpUX1wLmBmtGBCpOaRslPKUqYBhYeE5PsTpUSuJO
4zSf+Jwm5e3AUEwb3BbGHULY+cN7u1rJnUOHMEvDW7BVN5c3bVUQrtFDEWjA
P/isOa9KUzM1w7hToEfJcGzorw4645HvdpM8q6lvCzBvLvnaxB44nyb5vPnM
23cwrvdaBTwXq7DAtGbVuwyyB0VtXOaQM9+qFOuwllUC4446611k3HJdnYfg
BwHuQg/bt0W9bTpweXQplRXGTBNtbzQnvlS68eLzywrVz1MISONnsZk6DLAf
/nUvR7WsiLXOThGr5rYcMyy0pw+MFJn+H2D1FKwNslhPh8JU9XFZjL9TTQL2
K/PEfnpLzcW6IWG42KB48+AyVee4VcVaiTMMNSq/7Chboj5nKcglRpKzCbcp
M9wGfCKDxdA8zQZTOGliwPkN/zgg+lbqgAYAOxOYctRTGI28+CEDVP7Om0Ts
EuBav5sZku1k69UvnqMs574f4sn3ZrsX39r9CDV3KxwxASxjD4fYymc3fH5X
HdbvS8G63Q9pOU/8RX6aJqtLd0awv8vbt15nLDOKl5x1b4GKueoFsqB2wqr+
Pe9AWM4PuFy4oH+Ql8QEV6AmSj5esnqQgkSLYiBaFY5ilnPXkvk6Bzthhuoa
C/Q+sWd2TlOd1M3rsRVJgS1SGXW6Z5HFMRr6hzdX/I3n5OtWYITYpzXbIV6u
M4/4JC7JVDsbvYDNJN7MOryRGFcgcnMrJDFGY5HPtUyXBIJCMwx9QlmrcctE
bO2FYDG6vH69VqDLE7nr1Xu1/OrbK2f4S9XKnIiEdFzdqIjEBpWdg5exHQ0l
CzGTqYbwUoGHfzrfT49Ivp8mmXutBtFMJR3PfUGSHq20y08mbqfSNdCYaIQw
6EUjs0T8/j3Gs47NlTWvQBx7kmeJxS987ZjNsNazjRNDZqbFTT9URJS0OKhS
F2vj4A2xXr6Peh3W6TiUXXZjclL0jJcrI7Y7slOoyfKz4NgXyTjSj7/iTkkb
2I/Ie/R6Rim0xvj5DfMTnJXlxlxmEcvFEyKh4Jcw1bTYfvzzdQIYCfJ09Pwc
5uoRpkkzYbHxquwbwmpe++k7r/siGECk5MEUlX85BZVe1yilvsqFbHqkZ5Zh
Jxk/5ERZeLvERbcTt7KCz0+O9ZNaGgjJu2m2XM0yNQ5+tfkf9MGGDD+OaBsJ
2bfFJOesWhAegaokzHozHCbpgry3D+RihtgrI+bZGpdwecgfNfRClzwDOaMF
/1/3p4CTTEUr5QVJW0HLKtpBXAjfKY66ZwpQJqz66t5lmi56iKXPiiF5sGXf
L+MzcpiY//zC9Rc60Re8j7ICeMafNhu9P3l25zXwGIfNpiF+Z4vGDXlwn+yM
e2Kb6+ciOh7MFGbqQ+GXvtKRkNxkOJTCNvMtG/1S5RQ49cG/1L8Vi+JyNx32
ess829uuXA5IZA1rF8FCon5hka2vYtcNpJYWmcEMfS8LeVmwhy2vBXyMmwFa
MZOlQVzL9RpI+DZgd5xkkyZsk+4g/I1Wr6DU5a99ypbdeJ4MzuXtYpEAoByr
A5w6QPQ7No+YIwGZ59+IIctoIrUD5t/zVfKl42grkqfJAhR48mpNebOQrp4/
E9tJW+Ijku89TFf7d3BrWYq2iSPK7LJ+HWFQrfcPBqZmdH46Z5Af5wmqmsTP
Z2UTFQ6ikit1LbHy2f8uP2Gvx6NzGOhjCXqC1gIRPJWzvYyUqt9GugpLk7cS
Ti/YePyx+xKdYJ8j3DVZt6kK4TywyGORQFQVdi3MHILoIeJJjlE2MLxIdAfE
3Xnol8NI6b9pwTTww5WZjxj6gMwm39dO7Mn0AvWP7nO8j1ynH30GNFkGm2Fa
5i/vm98thIwrDyZKU2Cn5aoRFHNJJbIUL5kVGNt8pBoSUxCJjOOxuUH9GXS+
Ndh4mibsG3dwyw8AopUq/MzpuzNNo/jIapA6qbuNk2NuR+sm5etEJTcJIT7U
LFePy3XNh5zB7uLmQfK05M4b+uN+uXhFUKU/ZipLfi1qw6txv3iz8ZoRAM+r
pvZpBcNaWdRNgVxkMXazPVa2POP5PalaEVsoR8kmKOobiOV42t+E4BIMwPFl
0kchFF4uThuCm16suIGhJUFnzLDEw78bVhljozAgcVHbFNGc/37ZIC606sml
FeG4NpBacRwf95d1wogub4CiEax1Uw3Up+gctbk7VVsj3/2JclE++uoQFw2y
RMxsP1zCxISodRxNT+s294ZztZJPaAgSqAT8m9XHSmHEQkALLApQ85bAjLlA
R4ZO+ajpVdDPBm5+A2BJxYAPiZrhHpkspXTQ9qiDfOoyfUihP7giucOcORHn
gQvXeHNdvbpgOLLMaMooBjzYlmZN4viKZQsIE/94DYWN1NRYLHSOALBj13Ym
hEtPO26iMI4I85Jcq3oRWQz0msqsZsgT9u0GFm4JujTqg8y/WTcKO9kjKi2X
IAIGS72SsHr+b7U2ldeo96J6Wii7r5DUEsnSPNqRlnF8mpevISQkwhw4iAlV
ANaSygIFnvvpzkCL8hzUEuHHelf8+qj76U4T8NiTWtbHMgk8VnHaTmBfT+ZP
6z3gfTiUIOz52xqBLhoUhCSSDP6kWldyxFI/aUcqV/yCtXxNAWKCcN++0z9u
s1aHqblWR3tQ/39w+TQIAi91WNQv1SqDITjAAXEAQpKtETwO1w+Y0Prib0/I
CJe2vU9CEoEJlvutVk5wBMfw6E9/Y6t9HrdY5WbOGYH9Cx1aAmf6xia7khwZ
SrZ8qjIbs2ObyJlGSJJXPGDQoYoV9N7E6vwnWXnvihdMXvY2XaLWzNKh8aSY
Gpe23xsefAdf/aMXK5YPpoAc/0KkB36Q+2H1hxYoY2pY24m8CHRikPS+NeEX
hDdbB/+zdlgHzMubNCNhLJFYJk5e7H4ZxXiHk6PderdDSsJllXidaX6tuicF
r9UL2kMmIWUyCqyKN1RxSh6suYBbkPGYMhrsqCzAHLYreRbfRwsgG5Rg2WUq
D6EhCdTO10Bvt3xs3F0EpMnVpp9aZYe1ruMxQo8cvNR73339nhg1er8czzOa
CTIEM6ZzhEouytIzFNNb2GQ9WPJf9OQgHY9zJPAIC3YqX+9aEf0DLx3yulzU
fkEGbW52eYiCGIzaqS9AzFhvizQ2gC+0D96aOkRYiQtOdUZNk11q9A8yktME
CtJvaoOOwWSIZGns8cQjSu4A12+MtN1lDx1kK+IqmZeV1D/SHm/4OILQ4fWd
lgQomF2NrgUN7Pxpst4/abxk/qjVqySHQ4j2DCYAodzcDygjMYpv6c7q+zfX
QT9PbHi0kiRkk7DiCGIn+a5tYRUQM/2Kdlg9SVRF65rlckK11MhsRTBWYfcq
Pef0VtJulnjtDgyUfryRsMEUbb4SIyA7SPf4F03PWY+dAVa8gEphvi0e8ODK
TKov7vCJK7ZLe44T8NEVbFe4lrVN3qwvEia9JXgPjxI4KfSkOoLCtHwqNJsC
iYsEWw9tYSgARVYqxA3hbDrh41OFDrk0VRaUlT16pqsDstmLXY5i6D4AFG9r
xq/9MEgsxUA/YT8nCpbul9W10BOVZ/aqAclov3QaLtbJrb1+EMMW612UNF41
R2jDXgC3coiEqONRUWFvfVbiAMuAM5y+krR7EsF+qyy0YHEqT8nvP/6aZyUW
2vrhJei1LDFDOCAk0YjodJYlBUmzmusUaGdOX8TCuMj2onqUqeBqTSPUotko
jBR+qgTYfwhUu6bFKYKzjtftieE6LYM6nZCDgaDpJEAWH/4DfrN52u1kMyMX
c/6nStrJQEP4prx+fNHrm/JuJ4fGH2cQrwIxcIiXwzLkA8f+yemgwxm30qTz
8SzDTawr/M70Tp47IXHBvUki94tXa6VU0RprV4juCaxgv4cS3Uxorn8BEj1V
FpETH7MYz4tSRJ3aPXzlnAQ7WAuWjDO7tAgggeG7q1B33jSMipVgq0NG/8T9
2qvQnufQhx29+TMkcS5yMZU9gCP16mL8sozuC/zn/mqpV1DcnghDSFyzMqFg
albHR08OvMwpWjrovT5tQokpDioIWqU4uTdQWk15vsHyu1nchl8NSq0T/wIB
1XSM+k5FF7Fk1++fZTzTaWi/bhooUatHcfqMUpEynUdzGOnNjcLYKrnYTYh7
YMioDP8iaASYerjXIS48Sz3LMfT0gQgTtXIx4S+gqzwLs5D6GVK4gpXSWzsA
iCLaszjaRCMobaUwBita5mQEHKq3vELNcvXjQCmRBFUy35edED+bB60sboMR
6bc1wZzVNwYpOe7oAy+dLyCQ8rfCXQ+RhJ2SJQWcW5Z1lAm13I5XHghu91Hy
Ww0swaT2KaPkHETibkeKcv923DY//FnScK7QEzixRBQbA3/0gvsAe9BrV746
/n16q+iCpanjtVtTmFhEuwn2pJJUdVOmTZiU6nZ+467c3IPJ1q54sSqAawA3
pH3b90cesDZLrT4H3n8/UJ7/Ss6EZF6k/CqaLlYN1ZBvVcBzhZBaawnO5Y4W
nXATMiqKVCfLHUtJx7nKMLhsJy8dKPJXqUur/tClklCxHfinLaCb7/r2xU49
q6BJX1zZYyzLpJJLzdUvvtJC11Ac+xSLxTTbRzCC/CPusUmpP+KyaOj9GNhu
5hllyVn0Y6ULXfIICVRncCfYQDKv+h5mpmBI5ECuPMAUhwVIgxHk7GIscxxq
CR+v5EOT0pvyhJCJO6r6OPb1TAaEDdSG3KvRK14E59nVEbriziGdJ6vP76Yw
LNxQJCGNCmcITbo+wrWStspHOIkMrWud/W07hcQ8aoYfBxvUk+AnBcYhf09R
y0PvV9Kf6ZnNxtom1aw04CipuRVY4vMLU40HHq8lMj0rFRcoQsfAcFS7QGPX
ww7/gXsRcMvmQL6lBjnB7esUGDSq1jzRSznVc3lfbS1NpBpbCtcam8kOjes/
fcRKE41aU44ShtnpCah2FKGNFjzSIsPXGusHIjV6e1XLmbx9M7af7hPtTve0
QthQdId+rXK4gOyDLdZlMJ93VxU+iQyHAjeyYH1UlEqahkb8rY/dsb0if1Us
s9e/nRMZ4M++DSCgPefI86eoWaIOG8MNyib0NWBQF+tZAiW+3E/k7vug9B8/
si9Je3mUj1KoLkQKtarizuSj5kxGDVlUKB91BPY/Szqtfn7N3EkSWvRAqFUr
nT7oOXol5vTxgG3Wb1hgn3li6rjFkj5y5PBNyAJiYYcxakfANCxiHEAy0Tq7
f2XSTR5UDtuvf5LQlo+PCC/yS5FMLmCO/qmk4eINJWMx+5d9MKeMchkVtK5d
4OwszMDpvfY6cZix+99Vxm8H6dHwqBkYKI94gnFZJOiuZJC+aNocLpZ/dPrR
dEzOo0h0yK333VV/KXijgA+sApRMTYDnNn7dHtQjceLLUAYcO7KDBGGshK7W
weQNsBjFh08hGu6OPEkxyYbaH+cVyKtRoD85HeD+MgDNt9DGgljBxFlOxDej
zIA43sgCzA42fPuiD8RnttSIqt6truXQ5Ku9LjRw/SapFVNdIAZWzjVMCaFb
4R2T4gQQpgqFxiTNx9/qHUuiywBn7b8BJiEgy7pKYIEEJMhAymzoDpFkCGPz
+zR81OLTBR8LbrejuebugVv8U5LcrisiDp4S20EFj3WrdVg3MK5dH8r3gCP9
u4clfi9UIcRbYHE33k5/pWalLpbVPYBWpeoTjTO7DGOj1Vz/uk0wQ9G31xdk
EZcAIHjOz2p6MS86IUZ+uvmNNS05b5SQ9i4mkcFGqvLSBBBAP5hYVgMypy3r
YJYv5TFdf/CeGJPysQKstwNmlHV4BF8FSgGaGvZ45Tiz7+NzgmKpgY/Lrt+N
3jV35a4B/flS4W50/awjv8eXXqgvu/hy6Bpk44PAGxJGq9fO0UhGJmfL5dj2
Nkz3+gqSoMAgMnW6Pj2Ob429LC0HCr7UIaza79hzcGEAeJV+yCH1Re5mHOYI
2Mpw+ltr1F2uayhah/rkOrIGXe16gjH4U4gE2sbVPpCt92iy/dBjboKHwh9j
A6WqSU+MBH8drTSMjirp7kGTqJZlggLB1DekhyBfiWSTePSaonpMLoTB3+Eq
NLmMqnCG+rS63TkCCxy/FmnZO89o0BZ/jtd8E96JYjnUjqVKM2fjuZNyjYA0
FRI04SsZ9TCj0luwyMmL+Zi5ol/JhnmLAr7bejlK3plhS5OZ1nToSvEOEXfN
Zh5Eo/4ORxrx8D2AnK+fwEfHpNiSS+6iW5CMP11zHrAcp6c75jXX1s1vZVBQ
21B6zX+wYj4Jqs4YsB7tW8Wy++CJQVv/D5hlCT3Pc0j4pVk2whftRnWToG++
RDmF3vhEjtckbunrYbGBa8uuUM/yLkDqi3WQfV2LcuCHm/prl3bh34j6Bc3S
43aHpUIWUgQ8txcNOPZl2YgFMPSb1qwm4ZAEVL4Hz219VwHLdEX9ojz8Rekw
GKmsA3pfaEKijQU0zHHfIxMN92es7Jaevh5iU/YzsVH8H19by6cPKXwunzvB
79MUBTvy6BOwM69v7zg3J5pGmw+vI7jyRN/PqBYKJZ4iggxT8Os1qYqChMTc
8L8Q7q2ow1rXqttDfIGf8RRzKZyiDjoLqs8TrxS7CvF39RaHmSjqrSQRls8b
8URpZqnPgIgk1q48E39htb58MKgHWX7yaOFeyT9KYMS1xOMk0WLlBy7lP4BV
6gBfs8l/pvA5UBT74vTvtBQvBMbtHVG7mZ4cUwelSS2eSZdZRM/apRn1ktVJ
Wy0wgMSKYgrPhlsx+Y68kwnIjM22Eo1F5t9iJVTBA54Rd1KOl8sr857qnLC8
faT2Z/OeYnxY8VkHgbUFe4vOhdu47Xbqc0pb1QxTDPRMQPf83pYU7LqmhQ+d
3myBZ2YLyGq68AC6J0ytvQKg1/6rRwR6TcLGkaLkKu8HFp0HOFGLNcUx7MZg
1PESHisQa72cvLfFpC9AHOK2rO41dRsSnbkJhDppzcpgxETFlMq/AKnvscnu
A22m3UnJ38Dg1BN7WpcIWKkO98sjMtQ1SOGp5eVJN5pM7lp3zeifggVaPFgt
81iXmdgCo1exIq0dPOLCI8LZu/olkS2cbkdUIO23BYn8ykEZZjOcmJrog2R9
eN1rEK+MA33btdpjINru32FTAUR59lbUdKEb8F1vKTuYb6Kl1UyK2o+MsRhh
ImFxhf0SKRhVeASiF4pxAA+wQPcTLq3busLXR+/MF7EormS8Bid4pe6aogOr
CClI4yghTkdPYXmqueUak2qkffulysO+dRo7aSCx5dZ2Qkl0cYWqlnnjVx9x
oM70zZ7em91x3phGDw/X12tU19yACZU+ydsdzo51iLfidMjT6zQcIRl/gQDu
fgptieqShOXFu0uTZo0EjgA3CGTNxnWy3FkCsAnfAW+peYhJQjNHf45kWWZe
wp9BL6qfIuknopSfxgg2bHaEi1JH0tKUqSK5RjYYbKZejQMd0+Led59yWxD4
jahKaFHMMuvTc4JJlqHXcjL6tL8ErFf/ebe24t7qJGCRT2L3283fTlezFpFh
gJcEAoWSMzuYDop3nVpBm8bjORCqH+0mFsKJXetcNv9EtUxjRkraVRiJ/98K
FJrJpfQUwxaqchqK+4Po7iA9do/zh00luXzlwMTcNMHaLB+GLkfsSmsPm8oD
NkgMPn0azczrgqcT/aJ4AbsEKvqSy5goNmx1I08A8OpDdtJNxrTXHPbVLNZQ
3JWi1bNDjV2cv2Ln2JNNSj3Gtm7Je/BzMA0STE0c9NsUlncq4LcHFZc/0UlN
7FpNdblKzGWf7oQMpNSNEdsYZquYixsRBpXLyQh0CVMd4G5uhS0BlX3jTQBU
uskYvLoUr4vnvISLJ2qOOdSSJfDFlGMyDdYrpSETdHgCicyaP/SypeCDP0Go
ZS49jt1AmN2I6H9DaAgOKNjZZJkU1q/2kwh52PE1ojvNusdEec1l6L9XNHew
3g9QcXNJMHOcbg54yaUCe8gGknwwEwjFT5Bs9lAMrjVxGbLx8Drxxo+7Wsjl
EG7QQp2tSelP9ml5VsltWMJdU3xMaRVP3s+ZfOKdJvzHxfJfd5V29bOtOTuM
rf0XEnApeUG3wHYff0GJTiqJtFky72Ra+vgxSLxg9jbYQ5bSfk4+URUGCNxm
XHvZPfSObLYTLQX+imYtp3zek+/iTTYIKN2O+P1n/LepVwZzUHHsSsfXdq+U
ng7oYckFW8fFPuqCOMtW/+Soeu725Cpc6qtfB8vf7o4BqjThNevE4eVBeO33
k0Ep/T2Wlq5vDjBTQFnfRQD2upqGTsyZuuhXxuI/gIyaIBhVd7G4gO8IoUEG
b+vt+QrZXZZKtaEsx2Zi0A4ZtJBtNpwiK1bUJOl7yRpFBRL/awmMNnTJp0fO
LblqmVfcNp2iw3ZborWuPbl0L6PKaOp27bsceocrbbZKP8heZ7IrcGM+5R+N
MjdeyTXKMct0aYFwXcGONdaqxznfhcj2o80xhYOm8IeLyCiiMg0TVq1vxm75
2ZwtwY7Ck+KZNoyT2VDHYAd34nWGy2ZaTsr8HtjFTopwpxzqfxHBj0tcMul9
T3c5DpnMOEtkGQIcw/MGwfSDO+QJpYdqHG0lNyO3kwU2uUf0+jc1hFkoUiBw
20leSg/B/5cbSuCerzKiG6fR6yqI88N/+Kw6MBTJnHDBLNS4yY3o4rtZAsgm
6dBu7B/fz3Dtwy1vU5SJBht8LEtm/EmalSCQDj48bnJZmYn4kryIdS4+LL5i
JRrHBvn5SRqFIOblT7pLfL16pDviPgScWB+bQ+EqK0s/qpbr/DJgunRwfqxO
uXsm3Eu67neSDe+yI+6zvsMkf07WJQ/vxJSuykOJTVdG0DTvrY+UMHqq8kOe
St/EISc2zDQJyGUvHD6lnEMjH/kWQaGUFHBwzZTPWkWPOgqdSAIjyt6tiDlm
ygPrkwYEHHTbI5fwcOaCHAEeshnN3S9JnxH6BfpX6A12guPqXymuFiaq8Abl
kNwfMIKtKs3QPl0uXpxDkQpzHjGRLhPTEiScuGl9ESwJm06D437z28XAQjb0
isSRdTyvJB9+5T6iiX8v5tYYWgklGg7KhsGpZe41YGIVdLHjCGaf7g1deaYz
bcow+bfr0h2VeqxKTsF2HjceYSeDq/aXoMC7zqE9uWGYhMHSH2ERZKewc1dS
BiKn9qoDhR/oCAp6cOIdI4xmGahxAZEpJtAtAuK6A1OYasucTU3Ohh/ZTp2b
HT0hEr7NBy8fL+lFOj/XFATJWzCWspN+izVuxCQULzz3LPH3J8xt0vS1ZsBj
7yYKxouBbu22K9RHfflp0cw4PCUxBTU12ztggn32FZgYJdkpF6drfRtk9lIy
zd49CSv5BL6mXdxLdDrf3ktGT00JPnleEhr8ti5ag0RJOfkbhhtms1fO5zEz
92oUDqd+S26CeZmRin9MGSqwpKqC7THGaK6tRDRIR92lrgbzsIu0IU0H3sKp
32+JwXH+90Xt/Gkc0scGMoQVA5oReClY54FODrmsYXBl51LiZV1u2bmLX3x5
ambieDebYCi3odWc2Dr8s6Wwp+tfCoU78vkXZQVC//H5SqSIvpcVylvxUjQI
81vaC2EB8sBlWn1mcUlnIbXq7EXxNit+JTxWsI3YvsOhXWUyi95Wx2n+pQMO
Hya1WlGLQJUrCn1S9ouQr+qRI6pKSl8vbStOsWa4CFQke6l0s5d6VUGfnfPT
jCV3O3nSup1iqlDma8gfD2LjDsiAUV1CjHqG/qfstANU4schLM/34yFI4qsz
Fu8e1EdRLJmzQdHcT1gsggUySqYrlj5RRNtkpHmhsHrDbX1A6A5CbHOIc/VU
XJAnAi6uP8jP4EF5CllUIQwu8+N/A/8vL5DJ9xTpP/Joft98Vm+HjmMzyQy+
m1bsApN7m43n9u/UrRbvcAC7hDxjIvgAlSDruFzRHZ8NCjuPyTjr5D/RCYxj
8Wrv7dVfjJmPFTq17kFSgLCzZ7ZTNuqmzDTLZ7Vsz0rKBec0zB1jnEEf47e0
rfA5N06Qh2ocVHl6/pbs0QbQLiOTMgpYsFq7SEAC8eQ/ZFkwNu/tfDLlWOkI
lVznGkGHx9+TTp/rppTF2mh2Q6IE5Mjfs5Ins9++TMFKC/ER1V9Xd/P7IHjJ
dQ92sWKSOV6hXAZBu4Sdjib+rtqLvEUGp50yqaK+fp31H0f/DAlRg+F8V0VX
k15dIvFNBZEO21j9sMdNAYbrV/NWBD9hZmSW+jE3WUOqf5xMSBcrU/EcX00C
4ubpXv4mqRkXiviGT/7Nj6mFvenG3MGUGQ1u7HpBE2iG+IOdI4DOLhVlIxPB
4MJ7uppeMCQ8knebGigsf65aSL/2O9gPUaiOrvLlKh5Y5qeAZhzargDkdotP
g+RZpAveve7DyCVbHY6QaFs5oe/7Vx8Ir53/71CD1rZ07cqfmwalBhH2jO6b
OVvIbUmkgcdJlZNCT4G9iN2DgJVG++nkwiPLv6jp6zLfw21geFkOZq7OrAwq
UQiWRWVlfBKK9DDrPnfZVFNEZS4VpdEGKAfkaEcUADqz6387d4/P1KIWwCrV
0FS2MyBms9kwbopQTE8Vhk1uhQykFnTKN3gDL+1E2ORl5OjscnatYfJN6ttg
JLznp+hX5M9Q7c3kBdJv5g1uRwz0DIlrP5vkV959GpRX535FQSAE/9LaUcPG
a9oUdVIHBPeN+UHfC52pFvXxhhwbVKLbDH8v2J9I+Z+vdq5k8b2SJoqRfqaC
IOPQqEXB09OoSYQdYt5eWuPuv/uJWngr73D+idQAV8/AYnfJTiVbo+pSYbJ3
slqc42cU5KE0PTtAhQ+lBbjnvm390XmV2IKnGZyfGP2e5/GM2EKIgDcfedJC
sc2XX75QfOjmkCJDEnTDykHC/dS77x6hAMP9zhbbf9TxGP9TBVnI4VyOa5tc
FxNxZNlW3ed6FMuNNu0kaCgzIoCoNGtGevtm2vMGnAG/Doo3VJWcpHKQ1Jg+
jqgN5TBggecvSAEDe+iVNy2+2S4/IZ0+S8ZeaKPVPZvc+Vq8KD9PG0rfSCU7
Be96+/yzpuPFp1a+cB2kpUjbtPrcUTgRjaKSiAJdP1NiR/Y+yFQHmf6+WZF5
smkATixLEvPajA2JULY0kQ1mC+WjDMMDKV8sjl4WEqgqotfermzmIxYzkkGJ
OCF442mGx9JB9mCc5aCdqAQjz9YwyqNEyGCzEwAt9E+gSb2PqW31tIc+1Wdq
gozX5mhNcp6OhOXce0IF3zGBN2lIoE0Db7vlFgMa7Xx3Vv2G2jeFZvKw51DJ
Hy37WO1mYQtHgfEMD98b0X9Ze2A5lQ3AG4WkIopINaKpM+D+jtRp96piFhoS
ZlYPkBxUSL/pA3++b8sdtmCAqlkbr8nePh3pGBWMCP80kipFMNRZm2W7Q2qO
pkcpQaXEVPYKD1sYMpFp/fGz1WCji9T/FMwaC3jguLB69PmXfggyaILZacmX
CjqjBumGU5Ys4vOh1y5Wd3VWMcC8+4EkfZnb0NhyV2Al34A0vJo5+VqQTYWE
9VEFRmpROAy/aqDo7dQcp2fybiVmTzF+p1c5qCZv7YzCyL5qGqm49U2JiBXo
8UjMIkRBq4G7gHXy28AsMUYP3VcMEnj7YtyPu24q0B6wvlgtBlHBLJ5GXL00
xN49Kz5fWZZLtZUEIs0nn2Wis8yDOahpXYK7peGw6bOmH1LYCAVilztPfvMy
ioyr48VBMB2w/QA1sX74mD66fOTET+J4UdBlk9FBMlenSKQmps8qhtOwihv2
OUUfLHi9dJZ4OcaY+kj8Y05qkXah83GmvQyE5sSeZ6fN+mFj5dZQ39azvP5r
vMFSGoQ79ObTrqD+PiLzmYRo4ah7jNUqxVn1EKOCZseu3wPtFXON6u4H2kma
ORYkVGchG15t0PTXfps1k80TTnXD5ffovPv4Y/03hwgWS4IkTDk94wfbbfEB
CHtMlsrdERdwlrBJ87DNlonditropi2lT5P5oqUwu+RDx6Gvo2YNkRkrQalS
uRG7cjOYYsSp3k45wAIj3yuG1yQ+hOCSAF2f56i6ITT1P0KSnFd3S5Nw3M+a
dx1wAywBiEPqR77J6lNiVmiwMx6H5qFMMz+OJfHhVsEjBzsdJxTdaoRqr69y
HOCwA4PQPcpm7rQC3r+aXBvBUJNdkPiEKcP3k1Cc+zzkQsTe9NCaCM1Y3hHc
5QJgfAWs+208ZQciVQ7ngkWfxxA8AncAdRj8Cloaro+KSwckiDTgYYGhScLj
0IWfB6lOM8LWoF3zbPBYhTUtHRa3+Mqq3sds6LXfbY2RQlKh7O3SwSvTXhV7
3XX7heMtUVKwyWbcJ3nR7uLi9s6eVzcAWXMwfxAk3xXFcK+7+F82XQRJrYye
pHEzrXP120SYOyyRZfDMW+xbM3igSVTs1zRyfsk8z83RKr3JhbMjO6QG2I9u
GuXWoj0GlfaKpsU4gastIEOK/aokjPTj/OYBh+11IhPMNcLlezuLzoVv5Boj
dwHEg9OeXJ9UUEV5yCGELLn50yiQ5TfSrYfWanUVtOS4itBX8ZNahEccTPwZ
FQByFrYwNNaLUZ12WP79PIn6xmlaMOJ+Lq6T1VshfYqLO8dxLnYf0dk3XbMb
teQ3P7fUkjLz+4YfCy9yBxVFDiviLRtPRKCMiOugkeZUH0Xko0NExY0JZWxG
pJJBGuQ6vt7RNkVH1M8nCi0K35AhZd042+5FqIChGnHZq215Wp+amfpnjA6l
9M3VSl9JOH4VoH3vr5qpqbsVgRq8oX+d0T6rA6xjGLdXQD746j5+L1RHXPYq
E4Mi3wIEjjMG3sTK904mPA2FX+ejRN3HhH+7+OhoTjmxQuffmPTTiXoe68t9
Hdvu2WXTGWioTU4jEpdlQKcim/DVPNwI3ykrluOOzph0IR93yS2OxJkZVVBF
sJ5WxerwW/0By/0IYkhbC/Q5g8ldmopq4gPxlXSAbyn/+uUzd8SUU3EglV2y
PEqzvrLvzkQFYkcRrffhOyyyqpiLYFhCg2HooSs+ZgUvM5mQnKj5a7IR8+Or
rdwZug227dZ8Gfvu6qa73knSzbOUVjPatHORVytCGFkz1cemXK2jN5d/yQXK
1TgDMW/OG2dLbBKkXM5abf5yxc/u0+a23Xz2YEMBI1RWLAg1nJJhrvhjMR43
9Qly+DDmi+mo2FHmepf3+q0cTmmI/WohZdYsB1SA5Cz7zmpLKbaIAbEZjseN
3egzOhIO+oNRiIrIBdD3SPPFjMz/xr+FiennwjXZkd8iMfCxL9wP983pLxhq
lP4pM5F2WVt/OOQR/XH4WDc0u5G9O8vvUXONHYlBJc3b22Dla5SBPndLSgj/
zwWlLmyf7pOyC4YHJqJx/Z1eVy1x/+PK0BkuwtahWXeImPLe/FjW043BkDzN
tfOFKeiyzGHeiqoe1zs7vwWGjswwEllXK35IhruYnDkWVP1WARZyKIzR5UNh
5YqjRt1+rZs2WUXILDePe0SCDOH9aXrfbGYQmwMlZo4/1RxBEQP2UHEEBr1a
ZgBD9yInlzjklYqeeUk4ks2HJ/j2pWtU/YyX/fAx4X1fhLuio0slSfo17WQ3
XsNnRYfBPkMb6eM8gMdXXGqofDCa3BtDEBjgqtwJ52F17A8olWGtjQjJzpkG
3w6OYC1x0Gsp5grvLPpXANeEpj5EqOZRkfNccGNGoLVGiXRTckQadyw13c3x
e40nOe38rVRQLXDgSPZ1swxKDdX8lGndB/NxODOv9T0zol5jnZ0HpH/tQ8GZ
rJ3pUX6QgQ3isesGCXILCEynXGwvD5gXqpucRr5/nPgWEVL8P1rFRHfq5ppx
Rh/CqJz9GhTwxUX5n5Eo2r25xhCs6Y6j8idi/BdnufDdFhNGWxBa+rjMh9NO
yw5jZ+2WyN6hcKjILtblm1AmUDRdBMUpjj/T1cO7Zw+hM3IcbCnzyxqDoR06
Xgx9KBi6rWwSA4L1Zpizvi+MgPL+PMvkr9X4RULsQgzwnHTBpmG0ZFMkXAWE
/zli54oHD0EYYiZkSaC2nI0wE4nztaScFA9zwlJvZzkcW+Gt08CcZcetwuyy
9mDx5RzGkNXjSCntS70o3hDLQsDPAUD6JB7GkC9pqPBiBtSUYtcHnvUxd8Yo
KbHOFYR1ZTtsu4U0RBRN+/ZBzMGcGLWiEYy7QjRdCaqNSlV8Br/u4PBgFYOd
mKyb3OXhPRv3Y7tmxsQbxIlt3JJbuPp8dGCkUoCFgCDMN2ofkt0YeRtF+ip2
+yxRsFyIe9UN2QhT75TKzBdMyA7+L35DnIJ6d+uT/KRRglHgAeplwzq/Sbso
HmBF5hgHHLaSGcry6meAI1vXZCWNR3IQ6qs4vGnBQSiWxXWDvqwnjA/81oFl
Bgsn2WyIuC2qgnu851DzwhXeb+95bHZ5mcJJYTdfznELdZk5RJgPfuTwqdGf
gAAuFhs1b1W52qoHqSVcSaz+kHB/jt3/aRlf3aHVQlK0zo21x9+Ys4n/4CPk
Kbnk2uc7hQ5LyvA25YKlZXftI1dDpupU9doDoJpovowR0K4N3Gqueq43eYUB
447nv/qWumb5W/nBsij4wS6ZV38JdC8Mb4TGII4Uvec1iwOCzzLz8zK0yR6/
Nv4vYn2O6etrRVM2m2p068LKSvOcXz1d2zW711vDDtzW4bJeCgP9Oj9yNtpz
L85hjtAw1OCVt20HpVn31tq+teCYulmCjGuvZMPDUaxiiAVV1qXLTVngO3wA
PUeXai0M1JYSHy5ZK1BScvrEnbkb7Yaeg0auYDmnIuWb6tMxUASozSxI7e1G
47GoRNTxlVfMWSYZ36tg6HpCpa5AWe0xEhg6+NwV4szlmhNHDVbSyAEy0DJQ
yrjsqxchI4ba/M/MO3WG/Mzn2zxglxLb15I5KJvfv4Oy4L+effbWuYaFRb0M
VvEcyo/xHq83CXHNm7JG+7nnhOYxktD/qzM2CMMEMruSPyerjP0oDyq769X+
GH7iqzambEoWyIQ1qogAuFXbVWBWELeiNz0j/XoD+f4khHd5FcRISyEOP20U
NXjg5e9p2llUXWl0gpyiqyyk3jbSNSjcWuzEbrA2zu1XwlS62FeNypRzwypi
CMnduwD9qNyiEGeX0wwaYU/dIlKMnDWDfxw4XCQXBrDbW3UkpQGhjIHbEp2b
1HQKBsghhVWy62NFC0MTkdNpzM/a1Yon361IxjEGmQWlNW7mKgTm4q/PEB/b
3NJF/aVyiKVvvWeZ18X0BKhXcWh2hfteMrQtL9TmdkjRir3CJSFaiJw7TeUe
N1/wTJpwxj4EckPuZBhdr9aqmmn1sByPFqVjQkq+IhNxvXGUZNvvrnCMcxhT
hXGmMVAXcxk2yjaLPgKQtfnz7oRin74PQNJKYmpl1KQmAFbPVAm/G02CT0ZJ
lxSnqsalRIGduojtxcrfKrNcCBrU3w2NTG2Qb4iwCPW/yJt9xnbAlA0B7irz
QuEHzp3EjXHX53JE032XUMEPSo1J0Asd2+ZDXyZ5wko5au2yNER4yaBr/wgi
XdkuT36bSMtoi2A/0SeiEBN2v1GoTavtOaRfUoRdQkFWID/MsnWOihhGi2UA
vTGYQfym41+TuCbZmxCGK/3TgVKpx/BK0fnUym6fd5kMZEAxtaQyCj7eRGh9
6dIM7w/Nqhn3jfFcpr5L/lOx9mkO+W/LCjYmImU+hrYYz4yqcgodQvXfrDGX
0rgGr56x94DPGB4RwiBWU12KEuvWMG1aa2OlSdC1pMzzu3PUiaI4Xd2boz6w
JJ3e1lXd23bydFD1lE8n0jLrAJd+tyHCf9HycQOtv3HyllKWE5rL/7gi1Ois
GcWA2wQBt86Qxp8tUFXJbi+qFLq+f7NNAUuY+zkW/QdjdFx17j2KISDW6p6f
PvUSmDVVLW/O5nRfq1u1RKYNbfAgxelQEGs0ToELXTbPwQOW9iSPVTAgt7Oc
aZ93GTdOM94ffAnEAErV9CgqKVSZpPrlluBIc8LMfeJAgL/UXAaldt4yKz/v
Unsvvz4bRXi3RH1r1uI36Qsyn8Yoq3+se6K7mjDHd4QZqBJhPeGT6MY4VzS+
+pYcvVvN+ee96Q82duwPX7MzzFtm4IV6ZYNG4Cx4+UreoKWbg5lE3+wEKkYa
6p2MowO81tWdbRFJGZbWwbqBigJ9Epp6PqCbLmmimz9xS3z799PmWvZ7HUNR
OKOR0ZJ8GManzxoGpRYey5ZvwhtS+R1s4RZtdMDxiYBU4FQQqMVesiloSuQA
S/ahS5znDwkliilbSLXltlChHqe35fktVsmss9rF/YmbX8nFfzS3bHFDUmR+
tP5tsbtwBJnW64p4j27OlJSkh2zQj9xxidjH95lLd0i1hIcRe7gt+vv3Qobn
AnRFkuKlcBeLJD1wLCcFlqDiN6jyWsQUbpoLBdwWS3m+GkTrg1f2fWwJadGT
F+AcUmIlJ1fucfQcLzhH9bVOluDflJRZv57YJLGYqqVESzyuI5SFeO2ntGGd
pd8AFIe28GithdRTKjI64C/GFCddsoSBziViV8xBRgLWdTGj5SetFwyw8YuX
lD8P1z8UQCwkRwO/kCstXjLhWBk5hPj9e5IqBonym4gbpkV/plmF+4qUi8IV
KYRAYJYPTli3Wnq903aH/0r2kGeiH/owwNoC0HadFT+JpvZXELgZBhp9M3td
8qYBQ5R8+UElaRUT2qZ5hdszABa5UoVOtRP6LswJNbAyYg8ZZF21b8R7IgKW
WaPVWrVtg43HbF/BgN5kFDboeLt9JhLSZCXX+jbP9DN5+BptXFO6UlkZ6IMA
AGUbeC8SgEZbEZoqxYGk3cJ1SKTbHrMsv08OBh2hWhzxzIHccFAP+8hB5b6q
HgfnXyQg4/lfXnv+M0ipC+uZlI4smb2eS6pNRNhLhvvaBCQ3ubnG4ogvTtws
Q+0UTwe2TUoO06KlO5hWqDKHgPyLHlWelJV3vwKo6awtxvmuRGXLYAXrXy8g
jG25S7wrf8Kn0o+7YRKlxoO2u3bnqCokLvJb4aD6UbSbg67mtkwulPzQZ84k
MD0W6N3so7vpS0MDh7T4OTo7emgTdjnW6xsB+1z1rtKTyQ3Vqy1+KHAlPiqB
glxDjLWTJEQQmialM015azOvTpDq4+n0w942sFZTwHs3USghwF8j1rlBdaXu
f+Thr0/rK5iYJ7jwu3n5VwbkDHutyLiACSq2PJIvRtk4zswwOImgvC6IvdwR
VQCfiMfyCXBRa5YBI+Nu2f5N6Bx0pkyQrp012AYULTvpH5kdXNjJN+x0utq3
cPPEKd1+3KO53l7LSvihAUuFBNdPALCOhm1lR4M/8PAs9erR7hCLVZbEQPwA
QupI17wI0Q+fO6BROJCqD1py7wv0OXuHGrCIZG4R0qPT8oHCD3sn9/S8pupm
xTHeFYK9yqQhR8Yr1jqqiTsdfHAr9OgL07Qj+GIRsyLyzm9yrYDXMhlw0p/F
LSdVWxt7tdUn9hRH+uZDIATO2btXlXdVIEnCyPd1jAVHRlz77WXqJhOoKzFC
A1wbyLYh8he3I2MgmGb7hQjxIpX3pp0qKn3jW/V2m++NFROkslZQAoUZuNam
FViV9ljdRqK8dL7wLvwKklmO6Pxbz7o34RwZ1enYYL2DUEALp7KI/hGSWZhJ
j/MiPgSCcxbU3i27CscTg67M3M1WxpkiuFKHmXKOQwOPMyQOFWbndWk/P7Zy
aSXSvHxtHlijbvUsQCVeG6aQQoCBWjQ0ev1WZAa5N9iDLH328f21ns3M5H6n
uAOkdS4w5NbG2NSQ+1a7IZ3TxUg4xneBVXEzhztW2ZE6lhI4/TN22uwnipG5
9NIsFJfgoWpLzv2+HHU1ZrumQ4gln3K51/sM/ZHZJjYeiXScXdarysT0ojJe
b3LdS0c+Y31GcBlZzCO2bNaqgxn477UuWmJ0YDlASdXgpk4FgS6x0IGr5WRn
B7zTcoBmApMh3G9k/oq/TDLvGn0hYm40ZyIFOHpqpgiG6X6YTlFt2w1YF/7L
OFdCgUP1DnBu34l0degxb814Jfkjy1V1n5wcFBtR00ln3ZfWR5gR3EpHbb6P
TtMeHhREC+mg9pGW5j57sg65QI6BFNH9ZB4JanagxJ4CMiqiFSSqeCmOTt2N
kDjrxlfVxmj26ciSDY5KRq5Epg/K+OeNhhD6kFOYqR33f4SLlXeIEsAgiwC6
hlzzcaFf2dRJK06uj3Ej3XbjFDF7RjSUaLxFW7bSZQ88ViNg8ItyHaGt6Fho
8VdHBt2EXwuaCPrKfiIjAEjvkpMi899rf3WwoqeOyefrU7GA8ej1CwJpsonF
JDOZsNjoqezN8c9+7gl8VNVWm42JAgDXJeys2TEcR5duHhCJ8vigyhfwCrGt
Nhd4heD7G7JmqHWjmIE82rUuNUthKdWRaRtZQVUFq+Vokfq6rgxLZv6arQVC
dgw6FgMnE525hz0eFMtIrGXSszw6c72MfSkwc+rqK6J+SqqffzSyChtX58GX
hTr0qhiRUthrlMZnfkcQ+DFhLkCHzMu/I6ewuLpNsE/2k1/QPBNKWBk/BDun
JLCtJ8Egw9uWTR10039mIBeKobt7zUXkukooYBmCQn4s54r07/6QXnYgsAT6
pSbk3AYUgPQ00/lwDts1Qqk/o1BxDCK6nomxbolgRJbMTNlHgrGoHJAwQeXI
MVlnzTEKmp1lCCWeguwDjGn3pz45ZpHaM9qTbw31PLQjm3i/scdOlnkMV2PS
TiSgijVLIiL5urJvVgg3wVnsIy6QwX9zk0w0MA/XIPymVQk038b3XI+Hv8+w
tDyhX2wSUKNQRNd+9tX4BCoZE6JKgETcnVqEGn/HCJqbjnep0OTEp4fGj7yg
F5tBkQIJrgkoTAsehjc4+tVO14I2qzck1zWU7l34OE9pcH9V4iehNzFHjB5g
+5CFVdmoUvk7gOil5dWIQc+6mJzxYeODS0K/bAMuF2mMZs2SVGktAtGisTWF
8uziw4LR0R3RHYgNiONKZXnukjlaEmhEkk/r8PJ1kxUZpjyPWdUqsIHX6WlM
UfylEjM+tQOrxe1H0wVkH/Ajv6pkDj2UvWU7zuOeSYWmwsy272f0prQdggIZ
MZ+Q08Svqcz2tvn5tcAYNjF4CSDI0LdH29673WpUYLTeEUsDYz81fyWeSx1O
O1MefZbuRn7oSuRoqfTVVCsu/7acsrxbqbu041Ul22fqyvJuAeKLX5rA2x5y
3K9QxI8ez7W4P64b4ir7lyhkyS/aOosI/O3eKJm+SB1OLhSNO4uDu6M4kvNf
rtk4qBmk3GU0P8l2G5kZzsUZX+QeiarD/zHEn19/qprvMe+zCIcfKfCidFJA
SzJESbh2MMhDZJFVTT8HVWU4DQjF5n4Ij+unYA5HRGXtNFqedmjXR80RSa1b
LqG67p4uuT7mllDBHO+xP0A10eS1FzmjOsK1EMvE1ktqqLyaImqCpJcVhRMv
oNwjVLdq0sZ28WkRKHawxdjMxuDXDt0PR0GEwRkPAbJwjIP508+TSuKn8mPc
+oux2/dTGl94PZG2OFkUPDBsp236HxmM6/Oi4MWOAQYMDSEKvI4+PP33Tb4L
rbx/oRbk770qPQzFInXvLNRNMtl8wviEoH+gch6zoSDsWNxZZjBzFrXWKKNV
p8RaGs+G7PQJOhdgYxIn/zAf31vHLfXlkKNnUO44cnTLsz+sFeAt7ajh72rK
oSeXyrI5DVShtTjFBEIqgd2GylnjWczMzODNQ0fDXl0LCUg/+myalWo8ywX2
yMcHyHVmw6yKe91tnaIugJ1LuN36cZqhlMjv0qlwDaGgHhfYs06a7bOnPQSs
4E4mDJYtUMmEZj3alMhjusNxH+5d2Taa0UhuJahL80XRWMy6uyZC5Hjo720w
Ac1qr+FYohzP8HGFgOaAPWgoXZTCsn3w1kuFqWaGKn/mYfGGfX5fH4ZemZ4e
EHAuvu7MZ6MhqjEBTh+VuPbLT+VXxgngUXb6DmfQ6koyPut4EbBsumOuA/MY
tHRMnzmrQVX9rP6JG1b5V73PU7HZKclVpXD60D07cHgriFB1q3vfa7tTuaz7
hedZ0lLfBvD8jufvPFA4nrViFqlGQPQKh8FxKQBsc3hFGMBXCTEthEmYVnZQ
V2jiebxS62RWPDO18AyrTg+xSyVmT2lsAvCm1fSU0qk2E1ivjlJ0xWtmDj05
mmCA1sb9eKmCisyNcGXLwodt/FnbW0o3jm6rLnV8XlRb/U3d4ZP2VdRNL0tK
/PMpJdAK1TxKXxymSk1OJTQP1sJ9J3ui4x7wdEKfPqDxQfgBGbMQ5/U24pU8
3dUHK06GnKglDo+D7rdqhK7EkxjiE7LBp/pFIY56SgC5HJNARb7Uh/7Bu6N6
qPh/QGQAM9cmLgqzPT6e995HMaIk69VHa2w1F3zAmBOsBx/EjrZOmujy81c0
k46omRIm+l2oKe/6Mwl3TMmbrc9K1eUCsu6+93d3d1Wa/aApeOTT7krqQ5pd
wJ2cTikAN6SHJAj9g4j5h+Pwc0LO7DZ2xu9J0c9G6PjTAM5cMjoZigSIZZZA
SoJZ4Yu6nor9eGTv9U9R8ChC/L8E3XTeKu9rrwvVmBCLtOjzm3B/H8DEIFH0
beZuTmU6GW4Eljw0W44xhY87Xwlw/v9iVKKSMDt69GHJn1fq7XD1zOsiEWKT
n1fn4cqsnRi4IkyDIhnMNcBx+ArD4OjoZ0dg6rIft8CZN5ZPe5EoBwn/dBtA
hqjCxXC7BcN5ZAy8ZhtelrIMD8RY6/yvu0aPbyAiGD3SvvL4gNGYc+eZ6H9T
DuoDNwkaGY31kjR7B6ff22ACbUggfZvpzE2d5p9mlinosRNvu/FTUAouTi/z
nfbvQ7of8iv5B1FbcFk8Cie/A3n/MbPF3dkUpksknfknrekMtBE5Ae3TLyBQ
qQnB4zjsukRSFxaFDsuudEBznkM2eNkHK3pgLTLiTxMrrhTi1iBM/6oP7x0e
hCjFlkYtkTXNpBp4yyIqVmBu/6gCuMl313LdUp3HxHLWOqy/M/i4XVG/n6UK
0gdH/pK9GyIMnr2VLYB02DixXWAto2eETEdEsuM/8B57lk0HgWr/VdqJaXJ3
Av2WWqluxTVbe85efs4wBL3EZSIAISTvH7PxWD9FdmLWFm+vfjy5M3A86lMZ
FBV6XsunSFl38utyLTIbyMN6WToY0NNgJlIOJg3YuIIEynCcCv93k4VwbFv5
HOVFKfHXDM8ux/qBcUchwOYItrt5X9zLYYQMmFFiuRwNU5JJ46qek7Uek8K4
yC72reJ5RZQC+HrwLG1tcNm3pWsrHqx1HdfqYoCQr+ifW9ur9BJrLINWhlUi
5xls+B5oB2bx1DMDrByRDX9OUM+nIJXFLHL6DlFrt4CxyvdCbBJ+IURAZamd
73tIarhVciSKUfA4JtU8TwnSMgIBQaa4BhHCRhbqLKZVloli7cO6o7FOawAJ
w2LVK4v7mInLPociqU5LQJ2C8Lk8ZjiDuWtYU/f8089ajiTDqziAxLI8LqHl
foVf0tEMZ8CMVhmLQQjoNwU4tr5Cz8lxCa3lgLTMv48TVHA5vhRyi3Guh5cj
pP5VUkK6QYEc/FzpngBAHlaexcoBVjXHNlL7jszsk3K5fDbC4e7CPRzTHQVz
AEjpdVVhH0CGzIMkEOXa4K/huMZ9wKVhToGbUbQ48UhbVVZ7yGDyED+xPNWF
7Q8/f/bJLIiTP/e1DC17uzMx573zEoYTAJsOUwVzhtE+vZkhaBULeYUb5RX9
gHUvXVjXfQ5IM7+ssAjEHvyfNtGC1FGacKhFnolAR6CB7tnKt0MS5Suk1aI9
+6xCAP3xT3WHeeambYY3lGpldAGZY4FTLlN3MYCAYgMp02dsuuRn7rcqrXu4
n0becOpPkUmJ130/wXfz2auSNfea40GpAFRtlUYHCTM4dVypp/hw6CbgZTlJ
cNBU+GNbeZMm47aIt6M/Svdb0Yulm9GeRyt3HViFV8/4M/MF5Tj5NcNa0JgI
OiG/iGCjGy9Bh4d/qObjiCaCNAgmgWPAAULoVD9Vn4jmG5RsUu9ggUfDOM3H
rBy32uhaLFEd4wkg1uEK2AWLrSW4uxkkizwWz8PeAMMdPuzsh6jnWtrpnp2J
SrVGJ1ZWMUuS6HOU2SW9dOeSQnjApm5xqWTham3866tBn9EICUL8ZOXXKZyv
LWSzM05zosizZAAVtjeUrlqnQUfKRxfhZqwTE9srlTiY4S3WeTVtAf2vK+Gd
GWv6m00Uv+rJvLyVwcEWoIM0hWl3akizw4gNmlBDU/93a514Z9BGK6uWAxC6
gvpuadn+YDHdNDPa5vJUWrzw6cT8/AmrbIy37ftAdapq78ql+erF9RjaBk2T
m0Chq2QEXSjdNIBE8MlXrLFzf84W1ZGXcch9s35WfS//Nzn/KJ/MlTMpF8Ql
Fh0f8Ky0PWaTRNw+2NtCBSf4dQV9BsQeIumyj6kVzsHfsMQzrv662mt5FpZo
CKngKBchNp1ePTFQCSE4O+BHtRpgNdmmBQD7AZ3qT2KUbpgB+HxM4N3ppEYu
q/T/4ZHGC+TTTGyhmMkCDQ5iqZ/zYdQq1oeUu3wotmi2JfM8LwKe3FCbtE9F
+sKA2qpsd/ZK48V0XeIvscuIQm8aRetLoXEAcIig20csjpFi74WLfIfHb/Ne
WA+cESfl6eVHc80R6Uc0ltgfannKlLF3J338tEViMDHhoGzbhyft+0owu10l
MV5qHk9V8GGuMvrGyARgti1LubC8oUZoBrMjOj7g/Vt6fZgOicUZX2XYBzUj
Mdc6GiS3TLIpCIsH4w/RB76QhvjqN22Bo8aq9o0e7UVKi+pmzuy9sefUvTwq
XD2oHB4/pZGEm3VEH2E/YTVGyPJb767PtDnQRDnU6gP5XtHcVQ9eSpMQ5cUf
fm/cFGTWNlQ3SSITE0yqTQt5t/yg/o/qZXW3ZWNLbIAM6DNMStQrXfK2cYdV
lTAX7nRrNamD2ZORwrMkqc/nPs+W5juAfO1QAZRv5E+Es2Urpp0BMwsOpLh/
Y/oK/3N8Khoh0HZTcb7cCrR6PsnC8FlvwZWCfxgN8FenngXjXjO0DLMpuJDN
bWRy0bkTaya24mjIqS6OcqhihBiYcC1nMGP4m1ZQ5J+dSU9o3X1CvrGqI4hR
OumKNN+a44Ecgrl3GUZeAmKmSJdgIaOX7Lu0ZG1ZgMA2j+dY5jmLzhcz8sn1
P7tC3mtnOb+L5CITp5nNUDS9SkLI5SlvPL7vbOeq3HR5FFAqJygZBzJLqArZ
ePLMqsd9n/ajgj6zzefKEV4chcL2olA6NeGTTaUrzD1dgUUyx+Ni10h88ty0
pH89pp9HPHJYf5UfxY7yNYUrdPtUrJs2I2yoZN9SSuNQktdP4O1I7+wOhrKQ
gII+UIrBDONFGwyvIgHATa1t2FuyH2iCPb0MHF3VEL0DFBrv7p78Ty48QFpY
9ycRInRErW8ea843b+CYJpcwenM//0eo8GowKNeuNUGlFoyeRq6EJLdTiGvi
xZfDKhmm9g42Bxcdm6kfl7R9BqpygcmFaDfK0l6RXmdgSTAzgTKUEYwkoDQk
41tt3uPhu+CaI5G+13KBSkub+0so98mXN/0Gg4wU9TWzMZCar4FLvH9sRL8F
t0aeDNnrZJ+KjppujL7hHPa1Yzjvw/ChqpwHD6xVS9ZjBl0R8JM8xv5qw6LO
CvudTMhkqHUFzULzQHTEtBCPsQOLah5KPHLAjquAJ6AuP6HsqHv135IsXcVH
iMLaznxoDnp4QeIyxN6bWGPtvURvlIeSbGxze6r/XF/YfR5mSj/VAYBT6PGr
iwppyom7B81RM56XviJhtTM1hnIoL+Ub71HIFg6jmbWPiiKIzEVxYVW1uzpR
WDRRWtA2W3cbS4BGWrcisbYRDWxbjEqg6Trqg/XnGu9wGPS+lWpBzzXbBmWA
RCr8Dsi/TRLENRgst+xqV3czsIdcjlvo8BXreO/h4C5gnylii1AP2tZ9Qaec
ZibTxzPiQfLL6wo7CTxxOOPhGMoSzeEM1zOkFC+W3UJNN8CSfxoOvV6pDIAq
5cnp3msWzgoADVjVVmfuAP6EhxYggQNqEKXQHLe3zOeXadJrgRM6qzhwRU0J
z2bZeLdWgDGN39z7GWUuC3islxYZj5S/eZ8E5xBk0XlNOMybkGCO6ecsOi+s
AhGFPyO0VQvUj+4cydkruRFIDwKhwM9KHOBGmudlbap8XKTnq2EU++jWXFIv
S3nSZpJKvz/H+JwdnPIONlb5ky4D/bHzti5EGD0l8p548N1dWplAm+aWItGX
Oxb7bQWeJnzVj7ToXZrGtog1aMhRt5m2vmJLonUeo6b11LYPX2gOh88sSSVD
2cRA83hpNg6U9w889QJ7OgoCPTHXQQsd/ruEQTfPdHL4k2OCyHcESr6KjrIh
IFzU/FUDdnwPce4Dt49QjT41QC1ycBk3604UHRwWWHte3xdrzd81Ajbhlj1H
7/u3mf84q0jUnZQfSqQfcyCn1jC5zwwijjzgdwgrcxwPRK2en7sPirdR0Hco
JGB4JJqGt69ItNNPx7PU9IqVMoM1Bs2G9Wudx7qIpsJFRFP9aBwNvrzv1miE
dofRDNv70GTniS1nXeqlrMYprK2LNNb3b6acc5EsuE5iOfUUa42v9yXyrzQ8
0EjajzXhaUma1ej5C7emWsK4+Q17pb6o1KnpQ2SJEKhJzHK3RmGOpbtRHNnV
DYNtbuomn99dlSI33XHRKdU/UR2lsBeAlZ7aDuOdacCDmMX5cwyePPuoimqG
RP+j7VuG3P+h+hFvQiWaQAptZp4uM9rl8ETvtplqD9OSPu953ankOxTWNwgj
v1RHVanyCoYKAqceyerlc69HFBV3/yuSZDxgCmWrj//4PTJQVojdSPRMEzvb
bp9AIt5aQDt6JaFeAAnKZ7QK5lM1Wucn7byzcJOvxm4oWjcEHscCszXZKayv
IF8iMZvOUKRTTFqfpI4siXiP14EsuCO8HYO6ZCtjhLttXjTTnieLkQ8sOlGS
M1AlUPP5Q8z1tNg64SivGmCCYf6E7hcLnmZ1OzVQSU/vnJKEiQLKWKdtAiRm
piyTQFmBr4tqnoMttNEKCV7a7d+6IPabPz2MfZzZ3X/Wp9OYzLg1i0pcEHD3
Vwpa/CbFkyEngR4o5thltCDFihHmSgiHRxizRZwQGus7X+Tp3mE0vJAcu8Pj
qG3voZ/xI7I3fnPLbP60D/PnxDwsLEQD+f/ro2Y6GiB0CSgzxMB4nZrlJZY2
biXI48ZWP6pPYF/eb3dKuIqj7qbJgJx8bQB0AE1M+gUuw/+YYT1Tg7mBVxsG
QBSZ96CK2MVAGm2R3UEGBDNnL/74iWhQvtRP9hRZE9SO9dQBZzhhpJHijIPt
uvUZ8AOM9YL8YB1PZ5wfx5Prlnpbk1t0uxlUJ4PLxjQLmmWPhI/SHJTIoTQh
f8k7cs9y1G+Qq9P5bs0CpgTZJDzMnu0Y0wl7dBzS5NoVLXDTTkI6VzB9Zg/9
7XclusTuz6UX1MxXY4vS3wUGC7mZU9N1/z5A9ajB+DzMbz89nA37xq+nJbXD
6NzQ033fZOLX9ivaZC7d9ci0hwlTWcpJg3AjiCqsJdWLtFX8mo1Wy9EI+3Qb
dNZOXB2vr7ToO+lqY76zbOP7OG7VTiM4X3BkfUZaEvYUW4RnNGBrvHYOc1u0
2d3e/h7mqrBu1MW+RccYJzXih0xT7QjS6mLLjD2fvAa3GNsfBYIVn+5ZDKfG
CgxF5OMysSPixZAhwoJ9D7kMYvLpxTJ+fgS2p7h0P9sqRt8Zkw5CMJ1sv0lu
i6F9WyFBMZRF93dVvK58J3K8I/pR3D99uvyW1oX/ctkvXq2Wm8dwI6DKt5/y
687MNS/l9Y6tNUN90AUsWF7vSN1aYR0o3VvDfujKJZeqHNmbkeoQ1iVfKjHn
jyqROL9a1FlXKnq+KC8u7GAE+FjHC3+zXQMsNZH/I8yOdaXALSnoD/y/mDVZ
3tIElXS7kqYn4ui0+U4RmGFbifKXFFZq/wEIOJAeo6oVXwp/dR4GpSjLyKCk
nuJTA4VR5X1C82NMyTm2dKlkb0zQ6bZ6tGpKyyZCh319ORTq3ToKOzyZDQtT
h5h1RtFMYy2EYjTSx5qnh74zPnxfDDovqXNYzj5RC5gRUpvuG9jGKyyMt9/B
Mx66u6Op73aPEqiUoz8ZYpk8WYItnozg2FoWPg6VQeKlBvGummlCHyF+DC1m
2O+jQfP57TRaICYvaYaOR+uvasiHuDbax9Z8XmEK/pQFSmT77l+mKfKmwAwq
nfWK1fLCWMGYyOx+0cKWLGhskg80KFuFsg9DhPHEwV7+mX1rVQyXkT1PToji
A6iWH5ivrQzmH4jt+XwDPPpvnDnzj2FlQEs4y++bCMySPbYAT/pS6ga+JBDe
BlQg+WHOKkQ+pfus3Sm7FOc2yVKA1LudO//zieoV45uiqBSd+dmMYkD/504l
ASHLwLdn943bSm0haw9dFN0QR9Sw5zJSu01U9fN2kdI9N682jK1wM8X7b9GT
RP5lrluW1Au1/Xd+mEZELFarw6oW2NnFOwO0T81i4MlkY3ZAbj2VUYRHiCjQ
JMMqIlgQl+/2Hlckk+SjQfISWG7oFZydBjJ8LYnL68oAMrgl6NlnmYvzQW9y
hfGjr0TFShcd8HHqn2Bv+hvooSyJwZNUTqmn3+NiE20QVGeZBf/UtBZVCwnR
C0M4b7hqbUTAA02s55hUCU8ewx66ruZj/7DG+mQmTbTf0i+wYPm0/f0VYtJT
pqTsXcLrC+6S+PsTTMIKPValtOjtYZyv+pcBmypBbkXF1Wpez7u/dUwl/b9t
lZ0h1quLZjMrE8pcD+kJuB4H18Vkn+y0B503S7nWyNAvFFzK1NZgXF0OnLU4
S0UNsq/y4zLriTgXGXwOtzKPNT9BYHAkIbN4P9KmEY3tY5wXkK+a+q6hV5K6
AbJbCUsd2ojlLXDqd9D0rbXJK1ML6/6U4flewyJA1bzNFRl2Q8HjuA+S5S58
kb7sVKP/8MC8nA/l9phRGCmd9O1mB5stUDaOWXgJrpkdPued9gSu19NjHRD0
QDMemZmohxaUonrtw4/YYwdcicsu9BZcoaz991W/f4UubLLUnwJkOGdRQ01k
7vUO0IbkXcS99WX4kW0VJ0gaOwYaC/0e3Jd3UChFvidqtoYBTjZTZrz2ZSwV
vcKeiQbVJ0qus5YOwPoCdL1GgsgvmpatY2eE1fRiCeKKOvNtd1GyjKFHoBho
8UO3pVU344VYlLdf4ZvJm5/o3dz4b8rLirwMf9eh1EbEUtqvdsVIFUBEOj9q
EXxiLp/dlJPZCr30KZqbCK6KqJQLJSj6tj8a7XHlE4A5j9ALwJL0qFmxVpqW
dxX2M57ZtCafqQbDLyme7qKCOJDqz39xWB9BqZkh2WrNXErroDTZheh54xjX
xzyBdEX4CiIq424gA1Ry4BknuG6z3gMkLvpQNmbRS9jWBRgpx/187BAQCkdv
Z13mOBBc6jDFjtLDC3bnkdkswAUOwqgX050dQXCU0ub8N7TVX5ZpRbkBSJZ4
YiO65EXCKlxGBugVd7GyvAJ8crSCMvkovwU++oPzXSzv31A0hLp8/g+jXJZ1
7i9KBSSxRnGMXF46WruEWM/VuELLROGSxdSmgVvtF9friGp0HXHuCcznMn0E
CNEH53Hfa/cQlDLzP1NxNz6vIzir8nW4TyPiSi/FzIXsTgJlkcs5tIUnO1O3
Rr8gY2ib1CGMDMeZxLJBSBOVuuECgWOqY0NvkShLZwgj0jMEMlFuoP80c3QU
wN/ulZ9HGq/VYzcet2yk+L5XcJdxX8mUzIKn2p6VbZ9R3qMZI54NTMYAVnJS
RyB6qj+mpetqLYIirUqG71uZYTZcJup8GXKXPPn0hK8kAsm8OyM79+Xm7hBq
zpGd5OOovAKN/AyERdZRC86cni/pddEUhytYoaBHpF57ICQQ4LzCimG4YB7a
4f59JtFCUATyB0E1qMpEdgOb1AZJlSgEmVKRInai966BcEsqypANCE2FM9UC
FP0sCi7/lO/VT5KzR8+bOy5nUKGKnkLqhBRNoxqcdBZJF9l1qfopVCc7FhwY
Tb6hJOMqeR956S3XgsBl4FVdI5CtGFM1YOfx4JUCINe9cZF1gyIiPFbIi1n7
4s5NWQsJMOwWXM16CJWECB0mioxgfxzek0OnKz9qB37WApJe8z4WYZqJkyqH
el1Nz6+POSGW/0fo9C0qnYe7WW2mY7b6hNOnr95VchmutXEhlY3wMbsAY/dh
OyP0n4bUpymeKLP0BMdp8R/OHupNHTgi4/MF9VS/RhsJaxMTnJ9MpQkth/0y
i22wjXJwc31cjswyRvpj009eN6yAcgi1dVhXuM4v3nMOQyfewZwz5l5oMo2Q
H/oDJh6aSmP8OHYM7VIMEYAhRbwDKQ+GxHTgCNXttE9aqYHPLe5FdiZ6qY5B
h5No4biltHyJLyrh6UURnUGtsNgy+e46rB+BRLLFLNNDnvroEBXHGprOpqQp
jmzas/3r1M694qeT281fV2cJMfl1OC9q+UqiwPR5jn+Jd04CQtUJBd0Uz3mA
CHXrATppl3lUm/HjxmTUsc3zK+487Sm61hpqsFUyRXH5Ovq8JzPg1MfsWgoj
9f6/05foqG/hHn//eg3laSNbRcNxSVsj4xI/fxIOytyItBpeS9TW/M46pyXd
+vdnbKN24E97TMfR5M8xihcWQBT4oTnQKtR5e9bQF4JquUmLDeY8DFJO7h5d
wx1dClqReikAOKa4wM0h093wJldLt6whUgLTNQjS2zuxAHey1CyW8xhKpwD9
Qxoni793lezUWSW3x/ZXjj5mB/FBb2CaNtYQNKkBdUG6yFfF5ME1irCQ7m51
m4zuRHGZTrWgDXq6FjC+QzOyR9H3j9E7hwTO+jU8cRAQj3JIr3UK01qOG2OF
GSOMnl+7y1odSmCQcgovvn0Kv0o7VboGW8X2JMMF8oV5ZhiwqEYIYit7Dmu3
0xq9Nf+EdynQnDZkInXJTfBpV1p6XpqPlqFz5oNDq0voE2/9yptEIIbGOYoQ
1Xc4O8qfGtQGDayGeunGAkpKKp47y0aAdxewhFABaC+zAgA4m2Y4chmW+zR8
2IpPjvlwhrC9PxiUk4X0LwM4sbSSg8a1FF7oG67+X8lstZ7xstDRxLwoJinh
PbTuI5zKyfecor8xmvb13ShfJkYWM5+nNrXvrAo5KJcST8HJeLj4PePvuusR
HNPMqujpn4naIzKFl7xCsGAdMvXP42GAA9QrO9kxkhmH0JsccOeLJw4t6XRM
9IrM2ybNh9zrjem4uac4EZz+wIyKsPUCGuZxk+6GVHlM2AvvRrPiAVxk4hTK
qL8+iDTFw1m6ebaecnBRGbWOC8Y0z3sjfXD9OjMOyN8nIH2m71T3ONM+oktU
/z+po449o2Ez1glWAljOc6TdkvwMqM8YrYR1AaVOVq9klybAgNdbaU/EzEqI
mwlRdc+8lSLgqUa2Lq6q/W+5GEnf0x9a6Pc+CXuJGiAT2JgMICm3qYrm8/B5
1WR7H6t+eUhZY7zbgFw0fEXwz0tyvJyNJ8Oy4diSUmQTzZM42SCOyLQN7wXg
W69OS4HqYcVPk9hDQgyFDKT7VLZ7x0DVjuVho3gpg3AV5Nir/kH1LcFkmxyX
X+XBAiZhaHUaEyoRi6yZ16hF8l8Dnu23CLPT6e0dRmRj6TE9JECkowbLDG7V
0yrTJIeCZNePxckxtu6bTsc3HEqeF8Wdd/P2uQbEKy2XB7aoeTD//OAeU3K1
W5SqnmLXzrGrt0mKNT7KEa4ZXe+5SvKx4O/IC4dyXoudqyFTVSovO2wSvHQa
YSiJdaFqLjc1jtbUGsfVJ0E4a7e+Oa/4djSKJqR1ADrEp7yWRFnxfr7Vh/hv
TK3uk9GEzOVLCwxJrzTs8sARwPv0tLFAmnYWiEjCdW5QKRh/jlTUvAXXMNql
P6zJEILiM/ANcMij2sQqMaoCgwWy2cWBda+86pob+2N74zcnIsdBLAk5xLET
7vT6rFIv3wUky7naJ0IliU4PeW9y4yN3Ukq1paASgtgrvvEeRVa3Dwj6epZ8
lTZbtMylpzB+B//Av9BEOVZ21sOVAIGAJKK8odjaF3+nyWgZ/0vYUoNUmwKs
rGGweFg8EdSmANVP9jbgqvxYunqgo+ftK5P2DwisrvtSfBE4nt7674y64Oah
h+RtzOqKaQc/NQMSZPuas/VckRtM2k7Y6Edlz7I8uokbL07GvubUvihxOZd3
BZkad0JB6XJRsh7KCgsN1/1y/K4LHVXRmhdplF0LsWcp01JkhKAxzeyV0Jf7
5E1T3qy1+vE9TtheW2Rau0zY4MzaV0a8YfA+S4YvnSrBni/pIoyVyn35zLTM
Bdws0rv3W03tNZXqtMQG641oFGA9yJvfdHyIwEZHUjuE07Yugq3Df2Gwm/bc
NRsbGH6KIHocVHmukW3zF0NF9og0l5rme1NhvVe8chyZFzbvW6IN5plk2/yH
iirT8bOVzCq0y37MkABEpJ7aE9NCFg7FepyfA2UaGHWRjDQXSDCqZkhZvv0W
TXfMSBoaVTXtcRHBFZogR7vU5A8peEwExDJfP8ImeC2BGjuuML1yk01ny4vL
1Yni7g1GzJHSywI3YaFQsyUXzJgCod2Bl9OjnUA210Jmf0GaQolh5yieEnqH
txm/mVbBCAzSYI7RqzWI+3ei9nag0510RFWBAT0e5vCmIzmN00pNuBoloRrq
cvfcbEeO6mf1zKDIvrg66LEidfYChZDaticy9djbFLdEO/wW5IODlzRcRIzF
7rKVhVGXqg/AA+ivhllMLWSdjG+1k+XtQnup3hx7U3RL4nqMCgXV5KplfYL+
vGvY4gDj5aPnZro9ukHE7o4/QB6MBcuzuiaOPrqwOqjoOZEh7R2VIeiF497+
ma3eRdKEoxXhUwzgBOdV3KOD+A3PPT7SJDAI7WAqg2oODQfQJPDTwJzuTzRn
sk0Feqsc5AH6lOhQ3Q8HxRBjedUzztGCasRp01KSfl9PoqS84whUfI5R+apR
3iwMwgRT64NX4Irb/0vGzT6cjc441otvrlszxsornFEa1Yl6HDketXZHR2EY
SoZ+ThPfxAGgqzry9fy8iOkQPIcoXqqogCo6ZnnWddV9TNw5VIg/HBavLIQp
1o0pNWqCga3EjsbwMlDnTS8zYeayDNxVlOPsqcucCMVHPcaSTRVpFYWBH9/q
ESx4KqM6MAAYk8dMbn3e+lI5N6ZYpYRW4sE2D3bKT2paBJZZ77Bwye6K5wjc
tmJ0MdxGj8FnUe84VEj8SH7lKOcfooCES6Rlinyo4V5zvE3WfbeF5sxeM2YJ
0x9fUGIqzIi+X6FlvcWHkRSbR9QeAb6gzMp+tCaLn1FXrh86ykHHfeaITraL
Mx95a/EXhDKSGfJXRP5XHMRf621pfbq0Xffd/I1S/eISdmFyqQPFb1LMb1C0
23fvaWt3JMgK+eHYRIBKRuIkhla3tIoayhcPYeQG8aQMVGDmm3omAnUB5cWG
i6hO96FshKRH0VtN21BpieUyNVD94gzbzthMHSzRHbZH+uphnMQW4GvxlBgB
qvOP6IK1Sn1+KsQyqQ6Ji9vyqIvbm73WdlB1sf6ArRt95Z1kCf3KSKTj5p6z
CVu7GNZAOhMDbtPXnmRNpjkgKKscMQkLq7NU3ZODvdJNeUPz71oX45rwhdw9
hnhhK5O6LRnCgjGyTTenziARtjuz59qVzuUA1IcRuyotaYtQyclLguAwyPNn
lEe5YQ6CSFB48yA2upqk3GGvIZFeWOxHlXqwHs1x0ASoaH4kLCS2YdypYqox
haak8VO+IzFEWIq4lk9wbUhzlNx4Vk9f1qfS9v9NLvxrfQ4/CXIkU0/qxQwI
VOaNq9yXUiGYbAwDKD5vCH70LFzk1C1/FGaolrTqU2io6dIpXLAEZQfleeTe
TxG3H81qqZxuw42u3/Q7fD/hpzEvBei5XUFT8xQ7N+GD6BfrbdEINEaPVlPb
dJBwOx1eEACcMuruXMyvO2xDX9VwKfrNz03hhrt9DdKqZFYxusTRA+4tQqXO
s/e2XbO1dSqts7OWVCoW0blCEZL0Eia85j6rvJNfOD3mEDZfiY72NZ90Qnr1
RZ8Nz4W6ogjEdEIGeYkQi/WDhRx70zg+prHwlC8dtcAnDg1fa6kpsoAgvpMb
J0YYojywWRzktTui+oZyQbUMJkH/0+LU0YvFtQNGCIDsZu9NJQ3MtDZ2zQVm
SQz54YV8tSSlamxe6F0OxT7Ip0ErgNBe3vAXexjmbASRUcNxgd/eqCx4J6Dm
M220nmxQ+hbyd7xBymBj2S7so6ouyYYRb84gbqcVcgc4KxbYxX6NWUqI7Cf+
y8Yx6oZfMHkS6bp4LuPs4N+6Nt9ctBr251lFWMYymc/UnYZ8F9hqlfr/tte5
k1WLCxPwz3lVBG0u93Nw0NQWGWfQqk5DfT7KZufyS7HjutloGjrXQTwoDA4M
kxqaHJjGfUYJYzW/TrCc2THYSE6fGaRGd8TBe5xjGv4PI9XwJIIXo3AsM7Dm
FLZ46plA2t00u/6NtaeZXYitWz9sVandin928SaEBPmjZqui/XcPkoK+kutd
Yb12zhbmL4FBhIH3dyKgXTW68jtpnWCLuTs/qP3vfTZg5CUQ36FgTisMi2lG
DZ7rU796yp/GoIzFKhevEmfdmjnhi9fmoXQFp5twqz7Eppbc3feLR1wtQDe/
nPMXBNicHkWM+ZKm5jzlQoe9+DdT54ILzCC5Sbxkmd0ULz+7kfY8b2BT1Z7v
E/sThnyFO0C9zMZ9Gsgr3YHD78kqeok/SkVl6+c24uSvS6TkeQXxMpGZG0B3
FDurhlRXs45osxzVOw2x1knw4ryS225z1eUuEtDeQJ14WUEl5ujwr+eKVxDh
fQykvLQ7YjbQZfJcM3EUQ1RfwO8faPLz1cO2aQ6X1GZ40Mwazktm4jfquPRV
V4zuc6m0wF5j6dg/ITAWBJuGehR2VooQBuGO6rTCvnnnIfo6TLvqrJHwh0qs
O9gqkL/iRzts3VJsEoi/gRX8zFaL8AMb6iGZtvoQfURMakOqoaxl7DP/sD64
8W8sDa9Fehkr972VpORtozmp3XrYXpTgBebjSZqB/JF36L3uS/885MpxP3pD
/gijfNwcbDSt54N2Pi3QOH2n7Q3NC1nPdG+RisC1lk28pfxtOdu1aww4XQq6
Xft6TS0HVHuBqgBfdtxmDSU7bk+FGIoI5nMbs2u7sQtqtYPyX+E+Y3oN5G3E
e3vxguKBvx1UXND5r+NVhGN/HakbzbJHj2orlsL3/7hT8jhbX0Gd7z0PwXCi
hF1+p6uDgng6sHud4nu6m77mprEcv2GkyBEaOndlMF+X5iAOgEjTvppzuNHj
6xTJSqsGUOuc+6POrsIr2ha7QDRcw9wdJlwjwBPlu3y/C9/p7bR2zHB0g12e
ReCibAUroRB6RKPyWVyNvq1rGTPnSbKZbAIKwQFoPkn4ieAVbLxONGNd4InR
ELdX8TLStPFAn+BCj+eQ4CxIpGtvzGISEWr/arMDtkfOuB/qIr8mzQU5tBwo
Q+rq9o86Bmi33LtP5IMp+/NVfyMWCJ4/mOM6gQ3IKTMZ4avNQqxpADrNH/Cx
VX1HnynrVPtkv1/viXNxKCAQCX1uVG5Fzo4leFPGuKRisskULV70AHHUTR8q
6ZxmftXpy21b6Xxq1DpSBmvcl0m5zlliknLY05/Z3eB/ilEuJ6y/KcB0+Kl/
EwPIL/QVUdZ2xRdxnl045tXGTT083iMxbUjS1WUgH4fgftNH3AXpmd2w4hl/
o1EfFORd6tLL1FP8ERJMvAEozBQA5/GIzECKUk6RmG/133/UTp/BoWoUivq5
eZylwk/ghSe7TGPRWXn+ODWnIa+JMJLCIZKqNPqrdhh92nXJQO6XPDjETAvo
NLe47NYNCX1rl4zNWf7ncjRgPMs42aiu6mxOtwYKzy0jPgaLsuM7u1Rz1gUI
KgEGgk9MFOVOCe5D2un4+Qg4+Q1AmgJqKhYs+g1AmtU5PIsAmfH3FghtO2DG
1p7/PovNYdMQal6YgnB2OQhKTydUwcMr58aTQ/fxF6AqYGP/W2zmsU3Z2wNA
x8dTpgPlZbcgUE2N1WCoPcHj17tYtPlSl4dv/p/Fvz55B+SIl4c7pxrn0qQh
RExHyq24YMWGK0022ZdDKEZ5p4LxaYoXEv6vyEzmiUgGXzZHkefUpKR2lKRq
hZj5iz979D22VRHdwFpf/AhQhiXJcXvpy5svmkEqdEU5IQsCXsFJ0EqXU0MS
yZ5/UoDyi57MEghUPcUw58YE22qQXxVVYcaEw9e6CIuGB1YqQkD2xFOBAc1I
ek7NkwzPfjVACMQcnj8DUI2TgnS/X1BWjER2kBjuzUaLzPKFioCYjXKKQzy6
fEcVUzVyYQiobZheSTNbYpNKHx4USxl9I+kusZVfy0fEn3IbZH5dsEpZGX/N
kJT3dJg+0q3ihzn4i8Tw4PeFo6jX8HTznZZSPzq7V15/U7nDlixLbytulOG0
yVMVdx6rBa6RaqcE5VbhiZquL65WQ6fLP5HOrH+TlqcoWz7VcNTLYSTTlo0u
xoe1arbXonw3mDbSNOdIRZ5KNuJehoFtlcnkjDVDJszfqISxHR9wVs2X3yYV
CYs8AYYIKkXuUMAiFGDzgl+tx0XS2mL6grdUkhCTAgshmS9xvRibS8agev/z
mVwg3frh6SXKsl/buFR9VSDvUBzs3RA/jBcPAODqyU6URo2rYMcDTOLwb7NH
hxdFncxauC4y0Hg/S4MGJAcX3Oij4PyJ5j8fg4QsXoH/qttKFKGWdKisQYPc
pnuap1oSUMiiw0JYYy3KS+ymm5/2o4wvCs9esxlPAVNebZm6CeGhNQ3eVRr7
aIgiOms2u5KtmXcnbBQFWkybq9VZuiu9k3I0Ow5VyEhJRDRWKyGK0pUNXbIZ
YyeugqIsvkOwfKJTv4IDvoPq8S6Y7QPyPfN05ATFpA87oddgu4PwKkfM671J
OGKddRptY/Un2hHzv/oF4An8RR1brnT+Jvtj4X7QNWMSwu6iyvYfsSegS8Ph
mRzN8IEZIpCG7xoWP91o6eCTMCDvE5sa19VTv3LAkLOMZPbLFikZrty5z974
ciqDMJx5vfTet12NXkW9hJQFS8dcEPY3KyfcIsKVx0jpPwo+rNet0aqcy6cZ
k3je/9xcWiK25A9GISSwhHq4mcnbChvghTbm/2DsEtXtgFuCHwdcS0iUmxz7
T/hK27uNVlAxUgqqrBpL23nYJcv0Q45YRtHsr/tiO2WWgNKRBV/YwbZzrDSx
AaYqw4Eea6LGL97wiaGjY6Ixo6EmIO2GscLtUwIdDOlHfbRb3Bd3v2G6ihbP
56KCx3Ex7U39euHhH1cLgFuEH5hMb4KK9LrDi4hjTa0jiWeFCN1n/DKmVi2H
PsdhsE9/Sbl/It8cHCvAfAaAb7PzOJVajehJJ42X6bsOndHlDLMRLDBNT8CX
i4QgLov9dGCXBRZA85axBBLcd1EQr48TKW495ecQLVULM/m5VitWPBZ9he1E
p4tvImZxAkSBk53OV/x3DJCFnv0nAW3qfmgPg+ADVFF+TvNkYYbGKH24OVac
DKZmAz1TiWGOaRK9zICzaB3CaSB+Ljhkwo5KYqZ5zaiUM0Yvuo/EELcyk2c7
FjdLY4CUK1vq9yy7oR6Wfv/oCC+uezc6CyFUC/LOKnCD9erl1TywPxWHXOwI
P2nMtzm0wHqaxvh+OIgZAa4q2fwvwFLitvEa8lVqFRwnwQCzMyGufCShkp06
I9tIgP7YNtcmrCD+Mxc6HqGClGmckoyXpSXV8//X/btuIGEpUx0sh4xGxBdk
j20miEBN1NytG9Af6zPzGPp4gVpKHaiO2rrfHI+xmZ1kc6RGzyVbnlYwC2Y1
P+vcEaV8xLhEK/r25pmNN5dTnjvirk1FEJqheMCqbPU+PTj+36mXMH3c7YXG
fSP52p6heS3lhFD0u9mic02xS2WmoleE1kHv2iMQlim7XzK4HiVbh71q2Y6V
WnTzgo8T3+mCW/Eazd//nOVT08qdSyzLn96p4a0iezSkDPq8KdT25SwBfL2a
IL9hHJ6U6miX3kNQtRXgK58NIF/2qSc1+ojvhkRUVPY8Go+rqmuJ6+6PJE9k
w1sFwaV+MHczvYhIIBKmldTkU77iLeCvcoSlN+rkJuyWaEOknD0hKURvEg9m
jIGgzYOf8nOjPIjYxSPOxv+sHOWUekrLI2isH7M4fsymucHbUU5RHU4hxKk6
H9HvrunUrjOmJYfDSBDc0nzRdA0WLNiocQrVQfiNaCAVHDCBomxagUQZI9UW
xseImCbrYnsuBXq6RnTAW5eZypcUbsK8w8bpBhc15d57BYIyuuWUW8q1iMld
mLh754Z3Fcz0Ae0SIUhFWr7AS3VLglbW3eO2SCGHytfnDFjLQ5Ge9JfJiJx3
kVxl0CAE27bPicMQdK81JbjGil48gEMOWmhapM741sv4d2dZQvXwanka8drz
97iqMY/APvDmzEsmAB9eIUmavyTRqBe9Oh0fAyfEaQZq6GWEnbtlEXDwRZH5
uCWulxInx6+izDAlrejUHohdYctu7SvKVB1DZ7zCUYAJGdOQGx75zgpzraVv
dKc/F2a2hmx1FhBs7AaTaLmTqtfWaNWWxbmSpWscyF6MoFBTBtWhLaCEdrZ8
5xAsi1OuKuxaolGa2j9myL9SpvmYGcRv0Y1XorrNa4mmlNJP05tgULaSydWx
91fzQrFxrV6aS39IQ3L8UZrIS+eVVHd/Ji/lChwzZWjSsTE2W04WybcReAq6
ZixNnMAzjC12uh/cSKeaAiX31y3grhhfg+98hx5VJKj2y8tQp2eDm2Ikfm75
IUrKVdiP5OMCAiHq4oYWs+RllaVmXdkMT5bYeB3EajeaZik3+88VnRNBd8Y7
nrjPIo8ZNi8kfe1yD6j5kn3cPOxEpDIL8XRPj6MdJoX5zFuPrO9QyTtInc9v
mqh09ZUaG6UZiKRvbXLe4wcuqa8NUVyiwSj1l8HHc08zK15aDccA4UPuh2XI
97ew64334AXauweamyOBKyyzuvB9zmjt3P4N96IrW8FhJrRLG2NoPaZh0DSq
a1UiTKvylVjJNcF7/p5SaF9VgWo+92JBpeXy0Ins05Z4h+9BHQmltTuD9bXV
7WVCL/iW1IPjsf8+3Jkj1117Uab2UpjnIqm9YMShGR9DiCkJ4vX9cSX/ft44
4X1G4V1drteGGUiXazSSRt94m8S3IBfwt//qoW64lizLVYW7Tn79Yt2HJfv0
RTdmEb2IxFpw2R+Ytoi7dK+aOrhB5tDrGQUipajo0sZUeHj1r9qaHbBI6aF5
1KyIGxn+r4OQioCrh7L8h96CZKvMWFdSRQgfAct1E/iUPs2tBp1fCydiEyy9
7QzcYryLGv9NnCd/hjW5ysVs8vhUTPLLR39ewK27f2HYkciHv3dNMcqENfoK
XV1RiCEj3jDPIPUfNAkASUe+8hPKhwyKTW8sYZ/AC0qV4UQlex2VQvA6W568
L29MlwLIVN7cj+wczZbHp+U8bimrGituXWd6TGRMV11It4svCHLsECsh5o3J
oOiZ1HbGrs4VvdmFbmkFtp6qnM0HwhfxntE4l7dDHblhj2I8MhlJcDihsphC
NY66WO/Fxiavib+jQYB5zy2faPTLIYuBCSRU6dhNFypdSK6Unyghr1fQb1Pi
fsbljI3u78qmmLt9X/u9dztirkPcQ69Rxe59U8HGH7+ZNII+JzmwBu5/W3x7
s8E42gbfv6qFsXM3ukg+wUqNif5nnIH5e9cSRV/RZGHrLhqIK2X0VdhbYFbh
i9GkelUOk+09uZmbV/cAz9jS1Rs4zjKwR+BDDtdebiIccFT26/HS7CG1Bj+5
lJh6WqzG7C6tbLjWR2nvsRUSiK2ewZw6jbIaGiIjPGsAUBs84HhUo5VlSWOA
fgxLcxBWbrkLbKPeMhyAaDmBCKNUc8qgtFzcJ4XLzIQFo37HYu7E7Jz4xLe+
ThvOOaPp9aC95D5TLAVI0R5I5LpMOmzytsOErNOKKzXlizlHDuZQDqhmokLS
WiKbZAmV0vg8yCamVcKrJTpnoiQpOKq9F/zSVKj8puHrYrMW4wOlDl3EX3iv
t6/ZVCsGCSy+7aVJUYbv675DvkwDpX2CCct1Ivb6VYlZ77/bEgGPrbZUBoGj
jL+DJ7VKKKTqmrg1r9O2EhbBT7jlaPq31SGytxGR0VIJOMOV6pqvtsDKFB1t
SDVrkIVFdGwQ7mN3KxTXGHx6z1DPBnRnWSiVWp9fClvllJhSXmzZ1c0gl8kE
WDnZb7K2m5Cp4VGj8mcyj+a2DwG0eqAB4of0P5VZAlbgbfPCDk+1or7YV2zR
xf2k6JXAzjr+gMZ0/lSojHVKCP5EUMx/LOp7VscgIa6bdDRpL4ZdmnX1sliV
Ft6g//4H4nMONNEUcEDdZ4ViQymLc0Yb4UpvYYgI+j8aafT3BExCEEdXYyDw
0scKoCAwNW/EuF1yOtQbdAp7Xxv3or5448FQzrw0oNVoFT6/zM7qy4J3eG4J
9YgSK8AZgg0s/TFyhZwPU7T1gtsBNtgzl2acuJDmlnnmTFlAOokh7dGxAofw
3skAlwsIowMpo2qqWzWIolCw7SgetYrv5kBzCinSczTe6Qko6ZoLLpwfde+0
2pxMzEhy2+KRe2CAhusGjCHe8I6ZAykWXTRkDAB3xLGMeH1fN3iD+5OL49uk
Qz7nmeJOH2WqqErhRUcyaAgL8U+dCwSPVSGnC0cPb45T5B3I8hYDZOO8HG41
xRKjZOXQnqMGpfvWdiVr7jIpqyRD0bKP7P6x5tappzHOylnkIMKweyIRYnSk
kM1jnRp0Ua0WFBmr+DPOVlR3ExdjQXsY2Pa7UtHFHatW9oiG/zwNyoi7CD6j
XfM1ICklNjNZNZsIeW9tddlcIWXcrTiUBgHuVgY0ip03fL5fdhRw7obbtr90
qltvxuUEUwl5KrHT/GqLFmpDV9ozJsh68KVl9erXCrV/vyI1Vyny/WCjR5KN
lCOg898faNTOz0bmbnrdQYwDN4dVQCZ+APFNNE12fsMMQTLkieERHb+IL/Yb
s8aPTh/tZdjMofqgHg8E6qY7YmhAMjCa1u93JlMzQr3uzFZIar7P+aOH1c0t
1qkUyjxzPpuo/L5ZUvkHIv+37fanAW3+YXXXcDa8LfixFXuMFwVmgPGbGbVN
U+OcrtuubD5wwM9/E5VH2gbvQpH+H3m6YK2KskLqPq45Xo3/rQusUN2YWrcF
L8Ia17TIYW/Q1oyp0Vh/HbFFb3Rh2KaqX+DpftEPMjMDX6m5D/okx4iw8agY
bQoG8klpQhsLII+XU/qE+TA0xmIGtRLsOQsLiZhAOa/q8e6uO3v29CKisYWr
WuE6x9stjaBdekFGI4cHlSyNNHaV0sQAtY3di2ovM+VK7PatTZCSEK5Vbdch
CtM9hdRqza+8LMEDvJpoS60RO8dj/bUDc6RI7SI8A64+UJpICzurERm3z4+c
HFkAUjd6axhPyDMPuy7xZFWCbp4H2DuDEj1o7qnfQvO//MI9xL6F3VVwjHZw
ZEUVLOQnX7DVI6YYhd4USJ5MIe13XMsWJQs5GhAOZlXjF3UTolL0EoafG5ga
fMnnkpvxVoa+z1HANDEwokOiKVnJdb85Gt5cW7wRCSI7XcN6pGXdrAJc+7ng
WfplZEH3ocztbht5OYoDa57SbU+0zBAm0NXI+n+bKWIZW4Zr3tjZMfTsmQMO
YFLFEWeB4RcasqkoHDYQjc4YKH2ch2nLkq1+wTM+Td2JJ4AEETfmPv6leF/v
y1M/aOOaPZozPKJxoNfi53xVc62/UXViSTqghOqPLS0CKKlPtd2S+jf4dfep
9FjkbrFhUIg/3c27uhD+YlBR651ErQV97s6e7A7/nrv9nFT5ii7Mu2I5nmK+
z5AXkzVmNQxtaQ+JqYdwvAuRPspCKv6NzT5C7Wm8O4cWMtyBdt9bbtMBeghR
39ZfRItHfUYxxFi9Hv2AZf3z1HT7NtZkgMWJkwbMY8DDflE48ipQOvw6I+yP
u2RwLCd2fVIZCfJwllNkx+G8bc70jOGyGMngWfFJlAE6TjuFV7ZMUlmqFSgP
mhQ1jNtMj82iHy9ohSUGEknIIK5ajY0nzO4gbxAtOTquuhDBfvI4IjBM/4+U
Hfvng9lQqwjZk+Kp2mLSdXj2I8GCeoM8ao8IkUnf/jUx+hOHK0VsvRGZsm0w
0bBBiabpxYOhfqHCcjAhvlc6DTdFE1xxj9a51yAMRr94JjQD7ShhK/N4ISgc
v2bx/LsJ9xqxDkkMzT/z+gQelTZd7Vbk+LLiMgt1M4COYd9wtM0bJGxN7oCL
UZVlIU6tXR/qOt1b0V+HN2Br1HgGUlQBNxIpXq/rlmyj2RGYo1Rs/DS54B5w
prNNEIzLWzCkSF/9QJ3ef53QbzurbF5Ve7U/Ty9Yv1uQ9RaVuSq1+0MJ7lfv
PaqeKVMP3sLyIh8Vi4XIaJRPWfxZOH6vFM4yRLJ8B/C4Wqs43DTVvIQcWfj9
/uQNIKfUzNlRYGCr83gk9O23wyr6VS7WM7HTWipuE6YQHokvgMGv/7zmSaZ/
amBeJh/0TuF0lFm7ehe9mVtKqH57T8F9sYtMPONjzYQS8emBfJ8eGpWT2xH9
E170vRlq9FBf28xvQj8vxBeoW1ctMUukdE/HJaNS/hG8F2CDKy6XrhRVxyk0
63SFoTtmVjS1wLpn0kDivZ74vCe/qIju9hids+C0fm2kt8MKX9xXjRe27WqM
QjIjRpZGt+IUl+cNuU5b/FwKfFfgh/bKXKFwCRiK9wusLaeAVNoyhrDWuexK
wu8tN9q5w5cgADLMj/8po9tgpKKAgiJxJOzFU/ozb3dnX/EqocjP2J6eJjhN
OtxiyHdEyQvYn8SStFEy6thECQPmhMFmwBLleddWVWGBS5m8aGJoT0nvqU9R
keILr1DQmqEnAC/G8SpC5iP7KDqduX3RmVplMjGKKFy/3jghjZiCncOkRsym
JZis1omhVrRu3PaFLM3ohv/46P9N5I3FZmfCa1SM/r2q9o5TUBSDu3gbjAIy
1l9WM/zfxlR5WeNSeQlPi2OrLQrFKIXZpBbCSQQYBh/dncPzNkDTeQ6lYqKH
icJVfdQi9f/eXJt4lCQhiqRP4hkUojsG6YQ1bD2abxUNAuTRnetsAHHeFQ31
Q1uJON23kAjLMHq/e1bMk9Y68Hc+vvej75tl4i/EoPsAnfzLbvixx/Re/oKM
sVJurWzwii7iLDBMBbbQcDPfCLB1ScqdXmogswt4g9qp++1yc0AIRs9TXcYq
/Y8vIdYgnqJNEkkJf6mpXnvc+cSnHI5rhrAQfy9t0kbThGYOiSnCNl1UizQw
+LR31lud5F9Y7PiQKlLcGz7NW690pGPdqSnEz/uCxT+HzG3iGQZRrJSjF1lf
Rq8xh7S7ZcHMQlCMAF9JeDtLzHEnG4hR0DXN7Sik2MfgATR2t/oyY0B8JwOe
S06aUN1PjTFcQyYL81EnW/RxDafZNS0BOD2mJt/UArDKSe/6HLPfzaI6X7M9
QGPF5qetzxgYacjMmHf+c18YgItNNxEItj8u8+1r/lq/K/wNl6kOynJNhws4
tEEwS25nWrg3y2h77OflNGrdlSq9WH/QefSzh1cOBIYV2ubQq86wBxEBn+Ak
vfzsC0JiDidch7bfQMRcmhDsYeyoIoCSfRXWA06Y5I00uADzE6Ixg8T+ZHC4
Q8YjMBuzJ7yA/LBsnQxFPrpf4mLLltw5mDwNXr7n7bjCT+9rtCAtvwy4kwP8
UE87WDdODeG8h6NgcSblRc1q3VmYPpFj+/JlzbalJ9LVCMRaa/ualwZeYSWu
v4gEtkzggZNGCwDICivzLfdHtvwCT3lmokxEkL2SMZQdLhgeV5c3IBHws8GJ
hdDpG74xYDKRYM+kASsrBTCEgmRglpHsMdQfDQvPZS4RUbWYyHRxPzVdD3jY
RV0EI6TdndsOTssB9fTkcBRMyWrNvTSePDEoyxGFnHv2fb7DjBIwevfehkAD
G071FFsZg5wBzXpIfqW6/q6SqoSSC/jwovZlUm+lfa+WWvvTFS09LWc06fBw
tCn3pirucGRY1adZ64UiA+W6CHFXxQJKmEJtZTd/9JLUIsvPbqb9VCoByl6S
fCX8VEiShBLnQzbWJ/zI8FzibREO3FuHYCj2RzY+r2/lKR52wyFQYQmtmjJz
UHPC1BY0wGB3tkYi4OIFiLP6Al6qY+o+Fy0VhRNOEGBniIl7pWPiubXqH1Af
SNtQVcUHRUaPYSA23vjjYwgJySG1+iRUXRUsYsKN4hlY1mt8B8z81qg2qqw6
kuO/dvYjTuhkhVEPiQ5i8itCRCrbf9oZKd1ni/xrnBRTiLpm1yvbBuWcJLEm
Lz7enttoYonprcNj0iZEhG9WQsdyL3IQsX6+uTx+2a5I2HKSmpBxBL9nNNPW
W/eaNHfhbqtOPrCHmTS9FxIhaGk652SNSBfm19xBqqbSO4YwPb8Da5kZ0AOi
fFvhb07RVn26lzY2Qy0nHskDAk18a4RthIdCwFxl841HmDgqte6DTYs8Vjsa
paxcIkaMaAAuVnqrCqmCPnHOFvxCAno6i8hUDq4eI551PkSBPjlG4tgvAQy6
WMUzi0l1hyyws/QWmgFBplcBXNNWirJGaa23Z59WHH+ec8RgK/GqzYJ6uP2T
mndPQJnRLLKeODwBq3JZshrNB7rCEu8Rqh1Pafo+eaabnRmuE0mOVucbO4El
wjgF24ibAHszImKrT4XObc6hWh5cG4uRpTQz6vsHpIfKLq33Mr2c5gBYxeC3
4RKQxVrFGUou+f7uYljTqBg2HJwff+goN0KVFiYEUoDfCLwEIiISNjb/WLZf
Yw2AT145OXHWYu5pE/xkBN7jmTCDOxOi/yGVMJ7qO83m/Lt3gVOb8TnMI1Bd
KHpeUMMGUXtqp7VqW63NJxpu2LwtqylGl9Ueb3yJIbEEiBIIgCvYxIpf8EWs
h0iaL8Q5fW4q7RSHliJvwB2j4Dzk15wwJTbFNlIF6+fz61OOqcXc/la5a+Ae
IiRz4jxObsyS4tuL9zsa9KpUq3haafHaUNc+1yxEWATSN2fUqpBT+8O3LSSq
spvi9HxvBIIJUydk2OcDZLF0QwdR05wEf35Ao7k5xYVwjzt+d5RL+Mx6rn9J
MH1VeoIYb9Kez3OP+QxjPSAnBP1RFaZbf0G+AcsxkZPu6pkOBFnzA/JGJrJU
QZWA+DGNyNhWo06oLTb41W6s04nlWBZ95jB+o+2lMEzBTZQBc7GBtR9H4msL
KN7R5WW/L3y5gH4UxHmEnd1rwcTlWeyB7Powvqn1HkxuSe3pF5B9gPsGhsJc
fIqW+9IjgKMGeVFxmCbUA00ZB3Fj8BpJamnbolq+/oAXzmg3Ywj9QHxH1qDd
pSBaZR7iVCEvo7zh78Mx+sOmYZ/4zrdT/YxMowBVJr514DO9vy9jX+FoDZwv
rEHinrY9faxYbM5ADNCwyjzYMdQQKo+eAB7ksNIwgbZKWEMTDhoc+XjBOkZD
kt0+3mKYorSnnrX5KQQq1Illk+ZmOifZrHzhXs+5orpg7K2ygodax6zeAyCy
/Hu1mWSj4L7MavgpwHldwT+DrnPerdoVFzRsFV2ZP8hTQCDNQG/1ppbN7olL
0AypZfgHZGLotqHFucPDlH2fXuho58IRmDgkLGbcxXxIkfQMAres7SV1Mwlh
wuvtpKZoBjNta0XtJTXgNZAlOV1eyL/e/CX8QF//0a7DtWG7GTKnwhrr9Js+
KSGdDiJvWlHp9FA8UXsINTA9ShKg5u0LrdYxl+xd5DrGvXsLntgvzAp1893H
YgA2OYBn+2XPcaBZ5+4BDI5Ql2hkkCzGfkLbh5p1C43dU1/eH12Lj4SuKPTo
3b86WqoGNcg+i4HXsdpbZjGBqWxHH9LT7i4X+sELseWUbqTlzRfISz+vQxEz
aLJSF6lHfA+44FtxrQUrKZ6jg9nzw/Q9PnwvDAyYXhrRQkas4bHMIvaYM4hc
2Fu7+tEYF5tVUsUmA/bq0VGVzemQycHvMeC+bcSG4AMt6KcYraCL61i3Bcib
SZYSEddV9+ac1e93NqO4T1O5CcFdb1r5pwYNKdX85XFhhvNdLwT18LRIHd3e
wWBeJY0Cqu0knDHgdbSeaEVOpZCFkiQ63otz4NpKvZvIH13TICts7cKaSjuE
iTn1AguqVpi7ijQjZGfqemOjD9D987zBurX86VauHWK9YUShuMYYZmHq7jhM
eRMK2r73WyKy9OFJcSDh2txVDmkDL6lnIYjneWxSqBwCBuWB3bpu7/aD41lK
0a10tpp2UWTy0yYV8hgq68mqFUStXvj+yvvdUol6MzjStLmPo9LTG7QuaQKO
RnHsQqS6GmMo011LsPMmH7b3P+mci6VFlSZrIAAxOaN3uXcBXyK/lAfayShP
E+HeRIiVrr7a10A8qnBBgPFnXw57DJWoVGB783F6tX8TC0bZ/bry2K6qENYb
aWwj1ZD4ofa+bbv84wBXOvL/nfTTrW8ldbWIRONvxG9qBRj8PUHcztLl6OLD
W3D0emU4wuZ5IogZNeB+9i6N6TA1bR9K2MGgTBZZRxvzhSmyciwXxUy7jcDn
bxgpf4Z4Khj7dWlVNNt1c3IV3KBTtLkvpoTiGT5949gdq1COOwFLJyZaEdet
ooJiS5107SpByg6/p8iqviHtFZUY+3695YnMbpXUHJGgtl6C+RACwSSWkKEj
zA2WnznVzwqGYlmTWgnibcpVAwMWmmM4MNrnpeka0zQPNmuINe7XoIpKhPdr
U7NJfqAMFNlK8UxqadIR6vwgxz7X+wLabGNoIrY7+CeIOOv61azLLFl7835j
j9N+J2G0avz8ctfjUeh4L5B3jyEXs8NP6MZQ+ucqAp45+N63aexWNf1rFqdo
6o9AYJMsf1vWSZ7E0AawRB44zx0OAFeJ8DJTQM0ZBne3rqLZu0ddnx14gAnD
Jb2CKFJ1dLNKP/ll1q/A8lzR436TZwI5qKUsnqnvMs4u8vpprvqb5I06mjsS
6f8Myf2Cs6BCozWLLfrxJWORBLDMsBp4YoWyQmbt0dSNSqX91r8LWBx5PNUY
lDk65BeJ55a1dadeBrGG8cOoDyRVLLwgN3z20PjYpHsimox7G4pDOHs+34oz
zZJRkmWWy1Bh7yw68IrHjXU9yEHPdRb7k/uFDD2eLpKKASTskY5nxlwhvp3k
z0j5/MbE1xDcNA/rwB0R1zsShorSI6woqHJNr2RrEA4h+D0ulMn/xGUSZMpw
4i0DlVUc/WNLAx+ETc2oGUMmzQ4ngFgqF5JAHXm9O0DPqhQ8Xa3YrByBFUCv
Fs7KeJFoqqIybvDpdwVW3uUOPg+ORfVLTRyWQvjp/zGDng6zfHunbXO10kri
4JWfMx/QOHzRsSrUeb5kEZ3CZb1I6BXfV/HEt0MD35xbCDJxWn2CZE3t39s4
JREE3agCZbM/DKh7RO9XptlIMktS0KCUJEz7gwrZSeSKJ2gM7ypbS5SfzFwd
whn44bTk4HDw+EdzG+Uyf9ba+8tMqspDeMes/9AnILnWDe4hsMYyGgmjhKlp
N7oZVkw+WOAxLRUhVsX2eWnq/3A5PidtnG05K2jBNux8MilYMqtN+11fCiMq
taQri/PnLBko95Y9K9ehy1KQYlXDO3SXGk+366ZR0s+R3G42DV3nNFWcj03D
McmR6qNLuo9afdA6IylvpK9gqXGL1TZ/YnC+DW8svFiv3V/mCQaXw+BXKUvT
JD0RxQvGxtL/K60By66kXkkbiqUrbQnDeH0jk1Vb3NjtBXHfdy0CTAR8ZbOJ
waWDdyYkV7vD1uRuyssyr8fbZiuIx26ex0Ftb2CNOzkIffgb6Y0ppMrL7fto
A16EqFH8oQ4soAwm0cYLXylbVPFbPaFDpVKG17ibpm4hGXALqo4pBl9yLvae
BRa+CoiwUL4kg1RBKNooXFl0IAVZFDeuj3nvhkYB+0klGaGF8jnn7GQfodst
8dRMZjM7FG1D+Glx26tzIkyh8yHY7PLnCGCL+vkYcDE4Y5Xwu4sxYnwybdqn
ut20WhKtjGlvME9fn1snSunJpN4iGwKX4TbY/Nh3vWDGCsBkaL2eqyA/dep9
+7QSMNYrDtmD1EuBDkjACZseeeXG/WveWMklj9T2Z9odUrA1lvVJcdgcWWce
xndgBMQspYyO0mw0o9RShveKfnGYqovGWaJghzusRH+txl/eMLj0DLrRyDkF
VQuEExchVefH9/lnHaR+Ks0ztTDs2O65KgPrp2Fp7FdlO1ykaKH77QHFDUoO
NcdofdTwTNwFT010RFdZrdUXDATncJbHKbdt4FtpMBIUef8zRXO8WFnnNHMV
osffqToTeG7wLYUb7hv0DvT+Zq6xD11+Dakjg9wvBB+Q0YdrfnIhF8qqjLXZ
NKq1UVyLOOpHh26drVFlagtioENjHSmh6XNYRUfvniRb5Tm5HShqBR3u+mGP
KLR5pxHno6ytXW7CwSkonSMoOqkr4cz4AfNp3qHRzCEvsSpDPju5F9vUZfUk
3b91MNVwkQ/uXz9HvHM/hg0ohC9EbOwU/uH9lgOyHtBlhyceYeYuigcNECsc
ixkdbbpogQRNeB57U168PC48m917U+NYDYT8fsB4BatCtC08lxUOZIjgnvro
IFVRBuBomaPDA4/befVedk34VsYH/+qn/dHbfflYtBlJyUWGtewPyQkDNglz
iy4AXSjvYbIP9cLx/IKnC9yZkU8wak1GRokB77RJK/MDcMMb71kx5JE9T0m2
h9c1bTq7U+tZXswcRUE/Dq2TpiPJpRBLA/nKTLZUMG3ovye/2TKNV0LL/kAH
sW0B9QvvGcGYHsQ0ma45KdGTQpRRi9FShZ+xY+ZDYN54su2DsPwQBV/YC7o2
7MDkuIJ3GOZY3uz0alYmM1/+bqREGK6bF7+XXQK7blMNDiCIYrSzHNljAQjG
HgirOS6jDO/PAy7uwOdUdyADzDO30cj+WjY7eRIOtAFszi+lCvfZoflGPD+F
lWTpAUd9nZxIfMr4R2WP5JTwgfiVtjqL36hoxfbedjBRqmXUZR1o73bFovpp
ach839t4KRqlzpZAxdAvsgFChNLboUCRx6Zj5Qj3xZO9ZXhysDBeVRj+Hz1t
inGHGDNnIwPWOTJwES3R07JOiy8kDHpW3KaGhLfPyvBt/tWJu6bxh5Sw+x50
33bIE9LOupOR3YoqEZWQPu/+seaJO8bsyX1UwMwbP27yBxMoKD6pTXiOlVh9
msidGPcKvxP5720meItyJl1W5Bdzmx0clGGQYw4aoeyD8Gr0wyxE4lWFEEkZ
WxKzCXhUNLpAghH7mEAKoWv0qQM5zw6HbXGb6NEwAq/nGENbaVzLDYjFFTpp
xO9bbQLBC7yHRHyBVROEKbyfBXoCBlC3hwbXcnuYl3bISe9qnhjc56Svf7N1
zg40gjznGKXow1Ry4ZAHVsZJTQ69PNchOq/xADm36D9cJNXnxKD27W+FQkqu
biYYhP1+OfYyigPLoFN6BgNgunbZMIZqOoafHPOj+yvDZWZK+jARWOKzbM3y
98sMFZq86jsTLG38GChd+3/pOQsmh9xGZnROtuQYciLyJrhRZftnS9uN+zh5
MaLDdt9+4b+vkNj/TMx7EOD0/anksiIMEWtu0vUURtNBX3u6YXpCcYVhhzOX
llCcwH8uibfPkICHbau1q3A8pTFO3ksdGkA5hwwz2lRcwBAgXcIHm5fYCjOs
BP/DnN+/f4nfx3kF8jIxoHohXyhUM1k0/OdsouBPjScU4pvTT0A1UTJap4L+
OVsZmgpnwUjUxxTkgRkrEqRKqRBviI5p7aSIgnSmS66cr5bVBL4/t/mpKTMj
bYeD6ai8Tazi5e52/WB9XJmYXIYzqk36Z5iRZBh++aqMh8noVdL1m88kIjrP
CHreluJhwl41KawKjmu2WFuW77xH8wZJMI2/XwbpLv4P81VWKCWlh9CbPtVq
j2hxerqtzFA7O4evBmKsQKx2FPIc1NNEkyp7nF7DVl+udd+MvW7graVSokdH
BYkuo3wDZL5SnG0SXscaDbmoBsN9fb1jsAaG3LCeBFDOBMJXz00js1mCZZYw
AmSc3GN5HwpEv8MhOSlyA2JIqBksxJEO0ukd0WgNa6qxDRMWhGNQMbv8BU9v
tQU/izShgiQOhIRpazapJiJrja7+irf2P3rGhgra8uz5nH1BKw4JSenakYG4
9tkEK14qn6i4Sm5Ph+sMtrgYppawxgtjRbCKzXo+8AEYeU8KsV1RGQzd6pJQ
DwNvOdQx2IcS9pGV025+Si8Mb8LmtCuDQka8kyiyBJdnLUGeAgv9eYwJBM1m
BvOg18F5QPLD/fpXYBLgoQYhTYCNdloKxil8uG9Ywcfn5iAjjbAoE5nFBEZS
kJYwJxUdU7360fi/7JywnW3l14+9D6PYifKbIbi8ENIC11iW5dh3WHcF2oXv
lE7cQspnJ+Ks/kydQMzMbegDo5oF0KT1jFe7liukCE1Jv4kO98HL0klCZlmj
DCpyQK/G0ae3HIixFZo518o1EyA1VBwd9MbNiie+ePRISdHRtysHHzLxOAaV
28e03Tx4uaxfoatrEvfWgW6oBH/5iYLc8MlQATd3urxJsOPp1WZNvF01pgxF
39L6RBj2GcEq/SolVgeP1HY1WMhNVRNi/yL5i3z9uPMwLo3g9GzDISx/RdOW
YkF8ZX84JWYx2OZOWT/MVCxExuZJjvcdBs+jNVkiP2TXCYrspeYK/UQPwkUX
Na1ddp0PqjLEpLN0DlNs2afvHdV3eLcTM3zIEUIyP8vz+5a+aBjZDLJ4HwDu
NYhWR8MBDwbgh/XKZLb3AZRB1ynwimXDnjyv+ay4EXqDh8FREWCTZEr8PtKC
JphLRKQGoPSmsDD0ZvU/+xEL5zakKepAvelqBwf83WyHjoB5vO94dtJ8hbtf
HCVV6LNUEAqC2EOsmBW1Phb0qUeSzaGZ3wrgNGiiZjjlWPCuTMNOOKd6cPmp
Nmiy2TR0bIBvjNz29G+HheTXifigqQ93lKzbCeCk0gH6rArwC6hj8m4fVW5A
fw0w+5fn88ir2IDdDspZzk7e1/+7OCBQCDm7neaVhgUlQF+ADy4l0l4I1hI/
ob3BNFk6ETON9fuGAXh0HOKRX/ZKLQxYrGslTOFOP+3PiRpPpECGmLtY90dh
EBC9KsF7bi4o6gC0XzOJkqhEltlvfwRVrPeaw7Gp6QdjI29o98SzJVkXDW+h
2jQrYs7ngdJ2O/UWkwnbO5k/jL3aBihi2rKKAn6TWoTzSWoaIxgkwlqhqyOw
1FNRsAWcLHiYWwtxPMsmGuzKzlV39D48THNyZDtjPKHcTITeok1DJkH9w46S
Sxl7yiLsGF1uO25v+fU8vdpIL9EFqUag2d5BwAEyeL2ree63LRhoXkmUcuiV
R4V7BcyuluaoOBC7nw4/S1V/bU8u/9uI1/6u8X9p5mp0ILQWIdBNYNLjW8f9
JZq/AT97/PKRQ7bq0h9VA35jNSnCe6osJWCCNHnX7KkzkzNn8N3KMXIkI0ix
YNxKPeil8Fa5tFk7u6l0LJq8Mtjnk/TkbazHTVHwC1+vDfpBl7jImgNecD9X
uUB2Uj0Xd6/i95U3gnsUMbmsKHXS9kNEu1iJfY6Fnr2KdvLlJXOKf2sZ6oMy
g6vyDe37ztu702FY4wflRMrOErSoiLApFcCebrs6Jrp/z3HyhbbBSiaVtSSB
uC/yfx7QXmzDJ6yO9tPzb9stkKC/OUrSLNRq8kftg8CbEIbNXhfNkvhbkbNE
TeVesnhSHiFfoE3QXGhRQODYJaezbZRjYOvl5cXribpaE4oT3vph+5AyMDQz
tlP8zq5zV9nXejz844nhWS6sv1TYqwqxCk9+LCJYEYhixdxYS6lD6Uw+ojfA
q2zy+530Usx4w4u47mSErFf9LJLGaNymkQscTgRVhCip5uVPZerLHtXrq/ZB
1NUCbo3spPLFYxyP1RbABpT4xOtkdSRiX6qxKOlY5r1xROkjnOAQKRa7k43Z
Z08+2q1qr6NWstQl1NeqOsK6hfOSBgUOXu75lcWOXWr9jszOyzfyQISYYouy
v+3zShB1VG8APXCjGoCyA3uWFKDb4aKscpXS8NRfBfun9rXmCmgPQIV6mLsz
Vxn49q3018LeJ1c8SEd87HLtpLIqyud8rRM/nDkGNQgQQZy7mVFuQdLQTd0R
ALhTpAP/cgQfWZak78goAu4R5k3wXLWhHZKksaeRRaiRJKo8J7OrRWYy/nyH
KK4OdO9tq6H3KMHEq0QBi2qXJu4tctSB5sx6yTp8F2vjl0KhLvJHNxMCVYeG
CKt1RzgJdLdlGu8qJWw2bxQ2bEKveF//rSK3aFk6pNwAv5CBO1WXvjKTi/lZ
6H+H2QknIfHisxrl74VCDtwADvrOTWcyA+BRvLs3qLE9/+LPt6a/KM0CQQM7
YEpU1FhhBVae4OWhcOAuJvNqu+OCegqEovw5lR4F9Gop4Qf+JCT25N9NsjHz
Fc+qtxScCELbJV/Br23uXkEzzAOX8mgyxPjLPZDTGYE8KL8ibOsYQqFgmS4c
y8fZD0GQF6QmTFtmuLTsBEozrLxB9O4EDkhHhI3VbkarRW6ygS8bsOQV+Lyu
SdmZpzHQNOh0YX6B/ERp//WU1Dbt9D0jvtVirnyi7+dODDqqo+wTYIIK2bek
6wD77KOrbIeltMhTKLUOSJMWt+ssComEOaZ1OySDKSywrqx0QfST0iSXllsZ
XjIw91w69XBtwr7Zmo0tARHxiDr5nEd6U1nPjC6EXW2DBZaArCx62BCRmKXR
H0O59h98A4KYnOSF6XSvDVH9m0CqocSW5Wwx1Bhx7Iumqjbb45ggCmG3w+SU
8zj2y0IEK0B44S8v7OPph1OhfPDRK6YDvfXqEZ829HTSQ3C1BW1lFBO0wh+E
Rx8r4KhHGGB/D5mj0jmgWhDH4vCYui5MC6O8/EnFyStGCJAjM/ygPlfjWvza
y3WEgYNkr8wpCWRlmRDrUIWxVIIP/H9D6QIfEx5apqBFkeRmtdXm3PmcIh2i
QPkUZ1V6xF2S3C73clwYdsNxJxN/gK0gHxNENXAW8y5vXGk3qeqb9MLf20oY
ZXUla33zJ/s+9CvuClcYzGktC6zkPWaIMCvVmmCzsKpojt38EAdWADQAGfUt
1YR6d+/ceOL6mFrtLF5klx/4NZtIFlIinXnhiFV+9Uuye9s7j28GmlNgc8cD
TXz2nMA/SbtBz5ukBbRw7gy0zOTU/YbE1U8F+yDeBPBZSXgp89UsEukrBfe0
tz8vusERhJ6b/ltF6OfXHK/wcLiqAwZ4G4uSwurVN/Lmnvvl+1DIPS+Y4Klw
NAzvz8/npLX2tDQt4qDNrz0A19bkNTMFmtfRXBmDuPKWtwULIlVNPPJ7z1HM
aU2TD14E2Pmnf7hMxxRk9TaxkNFe0MyIyKas5zwBg2N9VXbnIltgBcTX8IX4
NXURN3elriugeBdpHrE9j4pWXvY5NWrUzY60vCBNekJYlaSSx55gWbIVYClv
UY+KkHnv+QedDZPv3Sp1o6rxRji/NjCtwVpmT/YjjqdgLFFDH2lr6D6vxWeZ
AS0WGj3A2GvTRfSEMu+9PAwzSmThLk3H3hV2YVoMMjJ9a/7i2aYNwpp+Z21i
SzBDIapSjmTQoWjUa5rpfnvPDJwBM082BYLEuVXR14YyVo2a3A2F7R4eI++1
VUKeMwlxtJIMcZbk8nvVjDuWANgzg9vMi9h1GCAjbjyh2XOrp8/b7t0hyb3d
uEa58ap0TBo05djmfnnCs7AEKzxEFfJlONm7YBEk3zetzDCPNBxoYj7kOejz
nl7TbPNm68nKSS93+zCMHhjstBnAEMg0EuoFhxBADLbtr1MpTEYuYQA/kSAh
mYKbC0LxJNG30zaxGC1ipqFWiElkrMkkxOuy7jG7YT+2N7ITHrXxEMV9LO7a
KY9sNv08wEWnmfgf172X+d+YeEzGurD/zOj5cLoxhFeD7qh61s5St16WOpi3
VHC7nVYq3310bekAigwcgsjgYGxkIEJHCTnvF3tn6+ZgLX1llRtDg8ALk4xv
iSRXk7d5YhliKjGGa7kt86cyZuSQpD9IybAV4Vp1TuwJNyCjuhb+/l6uYXLS
T84PV6Br4iIt9S9D+vMuSbT3TRs43FIKrrGHQMyZoOCmDoHw25zK2V9/XP6E
N38kkimPkGN80pS/7lfse8/EoosVGVK7Gl1WfsUsjgpubTWqAhs/dPa7xS6f
GFitcVoVGyxkMaYeZ8X0i8ydGjmyaoojtPWk1Zcu0Xtg1GJ9IVWyCQv3xXwu
7PxZ4/094NQjEWhgG/8IdUrgrCYQ+MOq687XfKh2jWDtU0ROoBOP1jf9mEQc
WuqXNVqnORo/mTy+plyRBjDcEh2T1l6AcwIxpKwo/rjrWWqdeRlr9P/tt9Xi
UY3SGo7S0g+FTL+SkYBeSsTQOKku+S0YD3pH/0+CdN/1DWrSuy59+WcpyI+x
ZQsHMY+XayteXdhOtjUZYJCRZ801wXVEN0pM3rBnj89H4q8jxgEA8+xCrz60
S6nvzjM1h8dq9ltLO6p+06J86hCf4NCTVSTR9N+d0E/CpsLuFiobq0gJ3pVs
WjCdERHA2uxoaD78Oubo+7aUMdP6188yLnAGIQwG1PRwaduBr1pszcZVSTm3
OLDLeUvWvnb+n0GN5u0V7xswA1jaSKULd82M6PHUt/FnysdWMVPfDD2H7LEh
b9BDxxuZRFpqv6DEmzbaCafFEtfZVjWKoGv/u4aul8Wtu55z26MeFeeDwoPe
YuaDHsBKM03cExa7F5FscO0Sopfpoapfy32cXt/h4b5OwzwSwr29KjBGUVFr
rJUxjLFqt+s1bpkK5THOY9NwXWmONJ3mkcTq0Fh7gkxVkNy71WTWCEwZjJqA
ZreiYpJiEA0gCOcOc8KmyJpCwZFK4ckknQTmPCcEmPEFYpehGOagh3FUpvbv
d0DKTY+bkzU6ayfwozJLK6IwtY7eOtxYKGrpRLA8MNGvVrJuC/7Ji7z2Bak8
hHDNSWUuJftV3veN0O8JMCREXxMRPLUDe/NKaDKoLZLQ9n1YsPswt4RXxkdV
eqV0HWxqMTesHMJAQJwjQ60A1A86lVyew2wz1O9WgqFE1y04GvjAJnpkadKw
cWlKlKzBXp1c8Oth0VZ+1/KDFG8bRU7bnxo6vP5j4JN3CV9MoNdIuEZoh2WL
l0y1+AfbLFfhG0aqq5Trl0oTz+PYj3wUJd4oDqPdAJuwoWp7VA56NHNhnyWw
dEXg6IxCDya6XuLfYRqoMeYfIyqNnYLrARcCFqbafcoZkxyQUAWMcMeyFS2M
naCOnoRIlQXczZQ+XNMIT1ud5RwamJdEKPGVH9QadCGQQopnNjvUPnRpx0n1
QcZipqCQuFzr7lk3z/Gw/5S6QG/oapHz5x2XwNtpBbZu6dAvFlQh6VFcfibk
IkMhb5lDPerOkwVeBrDxEAj03+u3Ul5b3hLtw51muICsDiN8AruVxirJ3jcW
bGsQ7HPnNKraRBbEcpP9IALEgsh5c69PfFzu0YD90ObbKEqo+cvISIiPoLTc
34L37gCTUF6qB6wcFYNgpyqew6VR5pAlN4rTX0qncebje76aDtX6YRp392nC
yat3av+2NwO4jMvREMZaWv6WKMu1xmbAkUwX/d+VCFlYj4VNIPWKlqlThdWO
gitDaZwuO55lKYZRbuCbgzx85snteA42ty1ykC/Osk3asklBPIBoPF5MMZyw
RjO6p/7vKheQH/ipc8/nNtlHafcQ5MTxWHodeWFSO09m1TDoc6t81fuA8m1e
byrVzt7ee4K8J+kREuO4z+kx2MOlSS1Mw8aWJGABWPfb6JAxt1ziHzAbrO2E
/7+o6NfhUZYi7+MrNxjVL4DRVVnZ55d4z3kSaVy/n8tOkihQ3XBe4H6vdsLM
U/h5gMWQY3lpid2e5cH+/jAUlTo2KnXdo0/7SiY3zn6pPzhHp3Mym+J9el8q
/1HyJ91+T4s0HuiuayGFperKKbrBUgQ8bda1zeTT8idBgXczuzSycPA6xcv3
fCxUP4CWqRgUxQHo4obokztEmKkwoKjc+ocKZL2IbpV6WIg7Ptb+iCf7s1xP
8TCe7VZYnX1DrcvVYZNed/kAMIZklio6Kczu8sWbdZPUs3rdrpRkiWT4TZqv
haBSE/QvgMOt8vOwjf8S/mVKp3pLACGLcyfItdrxsZcIlEwcXKPx+lnki3i9
TuNRuEy1j5NkaEe6wZTrmwmGhcGmiROYq5nOSl/0j95n7NAKfzA8bUb+nAV9
9bfI21lukRaY7l/TG1Thl4eHngOIsCj1kaewbhG1eufdEdsmHsLEn4U6mmTe
Inv5DwXv80/x3mit6mOunCSuP5YgLEqC+BQuL8aqRr0vWQ6Wf5WhhwJwmW4y
31oFgeYGsJwLQpYRoz9xZglufAfw8lmoEPZ9ATdS4dpBPVjwIQZ6kbDrsSbL
UT9N/HmCebmBBhHHsEXzn37mYrfXerxE/akqndD7INRdt1SRAV+QRh51Go9D
z+1eseWQdyCMND3qfKpIaLDR2dPZlkRicMym/LbMLt43JGsmaNW2OkGVV+sS
AIz9uFWk2nnA0cmGLBfO5IH37SwKDvadviaDrxMPC/VUn5raSr4v/oWUFQ9M
7kTygVM1MQhy4QJT7sEpzaOs6MXXVXCM3+LkP/HB2zEwg4FbO5qEHpx7dIEJ
LAAmvHUzN1fRu5MJLAwHhOsx/K81l/rL9PSy/zXTUam5vIAEyc6OQMHcijPz
A7H8KQhXJKlRFXd9ZVgwIgS8U7QlYcXSBzzRsRrtsYUefBFKxSqV/V2bwo1h
Le3AUUIUh2eMfiksmYXMkPGGz71reZecke+JZdXlQfZCizh2BYEmx7nSfgTN
i1DYE2k5rIAKoVz+SolVbf3i8y8kfFoaOVZTCpQsDhUNUp573VtW1KIONWdw
Kols8YWtHhBeEkR7ftQ/ZyJurWlQrgaMVgO00Xq1p1kpsSKFnwUuc2I42rBj
qSAJKfsbopYOXsxmYROQ5taFUA9Len0feam6gaAk4ecOOz6sVlSXcpnhv9EF
80B8VbGBibj8EAkbYSGuMqd56MjvOc6xqvxH9+fPxF+U0rqTrd3ZO0Ng1VZW
zUK0WOSKTQCWXSwr3ftca3taX5NVI6zgx31n7hxnKFzmIm9jU4xDObYKq3Qz
yvLUvAq/ztY5/M8DchNTj5algQzpfyCt+bcQz02vVPbJU7qMvTzyyfoHwM/s
Z4sRk5UghbKPzHkrpXpc/PDfgj7U0x+fslczSS7dO3MxpRudmnuGNianedEk
CUhw5xU1iTZ7fpLPLXICIpOlSUK7szwNw9s9jXllynvFbNB/piecPoxjIfiQ
8WrLnXAmIA73Ef2tljIuVOeK/8hP5kH6Xh90Q5g+QAgdFXkUtwJqu7hBd6hX
C9hf0vI05uCNbwJiu8Z2GvaayCqRYx54TZUYzbzftbYqh+bqT5Id+NamE2Kc
lcA7DGvMHD8bKbotdjf7MpRN1stMHiMKBlHQ6SMc5Y7uk4aZ0i2QV/ucn5ok
YWiKIw+ro0jiooWoi/8EHPu0yARblmK/ooeQbxQwuIHHCYkriC8hFLsSfF0s
Kakc7ghHdpgEPzXktZW0q5CzRFOrDYQaXnWGA9tvvQfHsgeCeufVtKEsbb5L
KdPThBlwcWxfdo9TbPr8tJCbowhpS+ohkbehLeegZJFqueulWuZirHOmUN0U
8wNEREoWxvAn3zoQIHz5aCsuEjPy2ogn0mCxvGHzSDvYDJYoro9pTOkn2OlD
xObJYpFYIkCGwDee/KrhmovMfxEsxquS7dkNNARJudAE6GS60NVAkVXXGmeW
rcOyVmWaZ94rk0d7AV8O8wNvlhy1WX7iGsmjiRNUW1vUvycjOafOlwGPR537
/aDyKZ/SeY1xTlpF8Y1qBtT6BmvEGANaMl6E6ULsL6S+OaTBWIIb98FlwSIQ
NCcS8dCi0aZrZmCquqMrqtAt7/cKPRM6UwqmZx5yhb4O6p6bYeSD5j2YoaN8
9LMUNDa8F9stHiTZPlLHX/Kh6+j06DCxevCWF2cd6f/LP8AO2f/50lRZjtJM
4eoWQI67h0j8ZePBmO6Mo+sWrY8/xQp7OfbQN+WgnYvNuuCBe6aeriCAlLDm
JueqWLKcEzDBRmzatyCkFJyf4dxxpmN7KQHMofUuAZVhsDTkrNEGU+fatvsR
SDxee0Z076rZkx3Z79XUrX83i6vxvgH7yse8Qo75AwklmPdkHmM72XBJOh0w
8KSRbtgr35VSvY5W0VBC4EJBCx8IJDZn5dR7UMNfdfMT9+dNbp3QaaQH3qpB
YCAzQaDU2m7vOb0CHgRdnelUdQDKUZTsEcg1LRefVBYYfGHQI00fZWWmyxZo
mITb1644vCQJsdx3CfrYtjFR+f4AiT9fUjmAZBu50cD1JWa+DR09j6ZEi/46
sLd94ywAvYLlT9vNH1CkZc7n5T0HVLoSMjAlKMEUEPZynblNVM9i9pThQP0k
dNKg+LZgYC5jPlNQaLtNVFCmqqjWXz8dlxxCxTdbJ91EmobxNQHJKVC7CenM
JCvnHyJtCYYvk31QO+KbFyh2cGp065b5KZl4MWo3YZGoFj2X7rQPV583rjMq
PVdBnzbNfLWq8xiAca6GCtbghzUBADZSIez3lK+HyP2ZvMDp0EPzf0q2wPXj
7x5GXFiweWov5Z5coKi5Bg373DBkHFkdn0Ob1z71TyxY2B8ZIpn9D1bbubtH
AHW1u2WUU0RiPLQ4celbRDd7gA0mqibjCN+aF/uqU/l9BX0WnK4DgZN7fCW0
OZ6q/tswfTVeFyhYGmlDSo1UhAIa/KYyOsAy+BaKZ5PosiT6q76KyKhY/dHc
3eGCSXpF63WIGJI0T6PnDI8tpqUh9oM+XLyGlXJDNaNfn4WWP0jxFgiTKHGQ
ZGAL6UUTC7Kx8RoifWLMQGs+7odZmpzMVLr978v3EftwcTtY6ggYNlx5bMgv
A4JiMAQt2fPt4hDqRBX85Rw0OFkXE6FV3IdAfFIyIg7CY/6bFnmrwxo+1WI8
0wasTguEZ+tFQiYB4MKeZFmrKwtByB/Tprxi3jbcsNhRS0Ebs1JOFemd2Hf7
ZfgNht+qFn3T8hamlUlmhw7pnsBOqBvwulDIM4llOiqleYB+e9HM+HaGSKpQ
G7IPpMfRMSclyBQVawtxtV77eW42UEMHzAvWH2OBJf+mHQklTnU0l9LO4G1d
HiLa9/5kLIto1lk0jH4WMqE64x7EZJ5cGsNjzhXgBBUl19w6GdsYxr3ZXIDL
Z10hWuVTaR1q/5r3vPoOZEo3umIlerPw26frYLNjkX5JfVIUiuhEbBTVW4Ow
yT0vE2jbPXMnzwnKPia+byRFosvvadXyQ+YHcExbmP2hop6F1GhHOOPOiLSH
MKHKvgGDo2ujucdx2ARaD9di7Vo5f343FU1i1OLO+jiwV4PxdLcxKmGnqDiv
mqilIpDhmTf3mDtpdq7TCMvIb5xi6gXbN9u9DNk84RbssMIHi+DCnMU0gZ3T
FaNzh26/7UxQAAWaagm3hDSU51vPn8/1HTvKbbA/Ry0TGMDKhviBl43drS0M
7oYa+5YOly3gI5DUzsHCub1WY/3L/0jGQEbULeVmpOn4/inRa9MPv2o4OfG2
4I+JMel4gJLyIRZAv2lgVIIp7sVfCaCFr0HhRL+SLZ+PRHCMtAxU5PUhT3hR
QytHdtFiu33mh8FXbsC4yjegxfYLibIIPxIlYzIOF3xpzcSVBA+lsukh+E0S
vmeZppGpU2E/zMvjLtSbBP9hrPNBu2s2zBV/sLvsuvbhodeRvMdx670rB98O
ZT2ZL9mqsQBc+wGiWDnyQ3MYV/MM6AgPSJbaXBFl+C82q4MvPMO/a6N+O7EO
q2hTM2t5NeqhVnUPpLnEtH8pp1QSIdttgib3JrSOdeUbWS9lQSP/LRLRdjEi
9lUDBAuYcvAlSnZzZk93TXGEDbQENA0x9ANsZLSWuqoK7LAIVd+sCDE2MhGy
SYWWp95HIem6If9A0oOwb3TlhYNJv68/bggpw5XpMWTA215q+cCT7yjf3/Sv
V/0FNVBtn0qng+2hiSOmc8J78JEZVdIoozf7Gf44p2VggkuIeJoE7Cu7qIYv
c5HpZd7CmndSqDJ9LuSoWTb6DUis3csSDllUM8RzdcOpOBz9IgZIA7Zup2r2
LxpwDLCrGjzcvBLEr3TYiOCriRl1h/3RXUhQG6mOF5R+eKmbNHptimYU5FRP
nLBdcjcahhL1a/s7VFblXP+zZyp1wbXNGNhzWqyKdCLD8/pROfIlQmqybiHM
/jT7m19FZrYWlkrRjhykmPN+dMS/2ZC3SSKX4ZyJCAfE5ESh5UdzcEfA8qri
7cmna64cHfgtex18jD6FBCM9uziLCq+bLSlFj1Cx5sHXVeWYWutr1uAbvhQI
hBsk88Biyt6uZ1YN3ZndgrrMQrBcwONB5xdkG3ZknTd5mCmwvYa44hAqLoam
H+7WxOPNzfIUbZ2ZaV6NFoxh6hPIJNuyg+ZfKtIPdvaDTaam3zymCNEiCsXt
PePbOWnxEtC9zodPxWYpLnXes0C+BXxMDhmBBmKvyj/Ou+3S3sy8wnsZ7rfk
APqitixozppyFbjwUTCYrK7FEYms2fcZ9MGggh8bpVFa/BtG+hEQwms3pfYI
fYD9NslBaSBcDt1J9lC/XFt84VoVDiTzxQc47Mf4/A0Uim2kV9dxfHJ1TeM5
4IVP65ueLb7OQoSeediA+/GgfbtEPWjt1AJ0XMFz1irmkEOJhuT3WqILJZ7Q
oLFWtpdjAoOS8EFTRLYJgkW6cWnSmwF2wevD0JMKaqwNtSzs+8vB0FynsAXh
HVWlz2VfA29iiyy1Be7QaqUrta1QLA4e567UzWXqOwazaLQ290DyjPn/NiAK
D5ABHOdMtcvnOXo1gXm01EVmJyl5G77u6b5Uf/V9OdES06B4sghsUcF0N8jm
jUc8uwHv079VblKNePhNzQw8LWaipXJ6obrzkRRYEnCDxtjbARCyHkKwHWqq
GlgN89vu3JOR2YAfUOMy+cM0SoNM6PqZZQDbUhCc6Ikth1+TV4AOTpwdx55/
2DnUZ5rTodhbV1KXq0or71JFAdUy1j0dO+KYuRKPZgUI1RQo8APMzNNg7Pfo
8xfM73+R8zUKcAmmq3uYw56OmZ5cn84/h9aidUlm6JFGQ/KXlvwWeExd2ffn
RIFVSHcJTq8jPSPcA0gba+y/DBWJW+jcxhL/YbUK1j7rJOoWTdRdYzkuaEtX
OdOPmZ6c7Q3rmnZlGqgY6kHM1FLrhkmJ2XnMR+iRdEc7802hWbV0GUGjwCGM
ytGPByjKTj7maSMRFnd7PjehHIcDfifqsU9oHtEM3unjoETGxpTWDSeGd3mX
lxkoPww1xAa5cT1wd6W+/kwym9rLCY+9xV2I79ScWLftN4GMcs0+cNAqKwqf
AWnW4RpZkCG+J+ybOz2NgVEo0SOZntAPNexQYtzeqVcXDPuvepM8VyUaAJOq
wsg/ll2tROq13T+RnZX+vgp9/kJrmWAazopQ0s7AjCiWeQLvDlljMryMFBiQ
igBTJdDoTJfTstsy4UZ20ZRfOUe+Owy+uUICDZfoSUqwFys/IdL0bBzLGmDV
pvEmwD3yRpkOdYXSqrZQZ6+1d/9PK3Zq6wE9mryleoXMdV/tO86TPidtmMV5
JkkelfVjJnJdl1Eb2O9Qqc8jkkRvcOXqZBuNQhvJz/JwQvuO0SSX5YdSGVXp
jw12xGgGqMIk/tMmNGHOt3RhGB98sOcdSA7HSTW6z9gB/gb5WYxoQYfjPuy9
x/6FfcCEkmCdZ10qOCXKyVExr5hJ+sjWBfaZIxp7qHmjJfDq8Gp/LdGhLXoG
7ts/cix0Q2k8MxCMvHQUhMzNvlX3vyH+tjfNUgV9jAlmh2EDg6GG/zybN0cF
PtjRAEDahwwbReeeiPVPxpdhgG3+jfxE40DAdgK/87Rfya55DZ/Ws5eyirVv
woRgQzwJyivPdCuAkf08Y6AO5dIvq2De3qrWMDxtfDG9IoF3OD98AS6KQ3nR
PXS6tc7UhFBaBZt4RWGqcUFN+mIcqHm4BxpLvq+Ma1tBNECzQKeajupY7Hwi
Hj5fJII82K5oPatI0x6h3NfYPvOv8wpga8DWApdK9kh3qaPI9m8cMP7p94mk
8FzRTdh9AEhE3wMqEGy1fxQLanwGAtz1PVcZp6W9BItmlan9gnLmQrGiZRTH
CuIMAqfhGjG7B5uKX4FNJRUzXve1oRgjKIZjGH4Q9vrIZYxKa/jWLnXkJbM1
qT/XfxB4RFwCbnT8IGc5hzimQ2Q51+k6Q2+4KeTbFyYtRaN5CEsDEqXzZXii
IVWXGs57ebXsF7NrYvsLifWLfRXZBZxMem9rdkagJFNsYHhfbzlwdMExkRea
hy0mCXPa4Y7y7jdSVryezkPdnw09NYAnoCILv3Pkj+TApqWYq/JxbJoMSZBZ
ZQhcGpssPOkXIRaguzXRL0xaL7ejoxj46KqUWBu9yHWD4A3+8HDUeet0Mrkt
DIwUqnXsVpRdvh5VLwA9v3S6HSUB5DFogCsjI2fFa3nCoQeQnQADfn61lZW2
iSFxhTlPCN6E2et3Xntui80FZkyho2a5EfKJID47aIxa4Zy7LOV2cmUmK4VF
TXiBaQBCf8HEqUN5gvLV6VClNAMe74QiN7rQLyEFe48ht/KqoGt3LWToTiun
3hJ3gGrUdaX7M/sJQWGPSwbaY/Ua7newAqVcf16YJJbz0bQTCND58kxQH+kJ
SaBL+Ds1yhtvu0KVdsU2MUpjJBChHYC/2nGx1HOHuNBR/0JAq794nsVwWq2T
s49M1FxjiCAU9KAS0HZbMEncj1r1C+0ipL6i7BBqVh/+k3AU16eoigUZbi85
lhBxqWSWoeILYkGifzk/B8rqyu2o0YI0+GDX0NBE8Wi78iwUfvQXv9TlI/7Z
BVOb828Wo2aJGkErHbJsngng81VA59GenRTytdv9oYwPonOKNu5I/MfJuOwi
uqbDtH2qFFXTcQ9s2YH3WSQLLYW9vvBr+JapTFV5OBD8M+MXJ8YNfGrPaZEw
XqsxWCWvXz13FfSXfxl8L4ys1nHwzE0SskqsRLso+Ke2hRpYUGUGrHl48ZNW
kldWZvLOntKhkvbQZaRv2OlFnw8n3uNzVAReOnVy6hop7hRTZU+/eU1VvZ5c
ztD+40vFnfgMxPLenaLVCcz4veqQSYPLWMKsqjl7IKUFMASFuaMTLC/j26SQ
62flvN8g846cEzvea45m/zPLR3C8A/hN1D2nZHd0IjuMcd+DBYKKUfNg833L
3gJr7SQTsZFFt7MQWUIpB0A2vBMZicHHk82GereYv0nlG4ujJ9m5Qe1EfMAH
ptGRLN37T8H9fVppH1NR8ojTbzySBdwfDsXiLkkFLWvIepmI9LrIi6B0OrGb
lppTZS2LEJc/dBa6MUfSF2bwGShkbjTdbkvPab1pQ8IKr9Hy4OYaS1+lj9gJ
VttjU5jUCu8bEwbos+xy1pN5+nq+ZiZN62z+FhpZvh+aiIV0ZtCNfYUuyldg
1ZMRQC3VS+vERIrT7HPvCKQh72fj0nf51JnazRwQigrqoSd3yLy3DETcw2Lp
Mxacb1LDaCkDwDTEg/AWzolGrITrutgRd0ZTVHSFtJKsPza+PWjubWjFGGnC
5TN/d0E9Elxi86blIFrQtAMGAC2e8jTYl+I8Hq9sCIKLXIPJqRIFUU4kzgBw
W1SMVExUpLUJjtqz2O4iLYB8qNJ6oTRgSjX8jtTI5CvElvHGk+38Lr2h/rk/
a9fYB3wU/hTpIOlwCJ7lmT7lVoItrvzEEuPkguTwlNvIXbmpI+nekkxmv37c
TBSMjbKh5UMGUEmUxgM/bi4L5v5MTDyNf85bYNFH5bE3a6gUOthbJIU33wSt
/ugQ9tuyioeOaTO/ZNEybRbO/hdpDCasgn+spyzirkoMbBmBMEV2OOj1RIS6
5293jWCd7nm5jH8FkWRyc0oo/R739eWVNIkufljn3tHZpw6DPxDV/4CjrpuN
/CfqQkKfeCFnVQU5cAgoUO+/HNHfm5vhE6gqQXQ8OMzGvc//+J5XrAm1XOQm
ggHJGF/tegS34jagBiCVBh0im6DBklACd/cNWSxZhH/ZdPQLBeJar6OOuARa
GOWwVsRhkOkfXiqCgq7978M1QN/rmosYVQ7xBScFXBV1TIfaQ/e2JQYx1N54
z1MGYxRMxZnCUS5UWBfX9QimYLOGS+I0GWNDVB/yV1o9lq9bPCZ2kMq+YqBI
uWWARiWFc/W/5P+Kr+xDikq0Doyel0fXeZ+Xa5ZpDWSqO1MAtpcOYoI+GSbH
xr3rq3jMc8w+7MuCEngG6dX4hTaTT6YFNGGjBOpWCTJ2grxZYi2CH6toMxS1
R4Nd8oW+n3Lmvp7vJoquz0fI7kWCSE7ypKOz8VuX5VriScawVv2f/DfS1mji
V8VQswnwcL+vAkIfLTsJYjPlZf0fG99Zbf9ZzW5FvOsP/s+f5hEbSg5wYrDF
8EgV8y0ihr5OFnfYtAWVEaxXq7uE4rEKoffi6ZMXO6WdXOUtnqYy0Qodxbpm
oPKblFqKXX6UqyABxx6bYircmuS5xLnjed9BIyt6+A2gmiy67CriJwztWNyr
YoXP1yZtfZmGhOEtBI13qj4T9FX4nZan2kWymKVh7MG/53iWzIjnIMo6+F48
96qGUqto4c5Sdr42T+3JIWIgFpaJHEc4ZncMSFL2uxAw0APZ4eRnAYQARcuA
kX7KCHzaaBKQX0fNI+3nwWGxyvuua22xMz3MPNnYiulsTOoXN/sC/tncjQQp
2HCbsC7zAnV2N6HdfqEf+KWwaReT/Df5KGKCDWT2DjnfH5pkQmgneU9rxR2y
g5CV+MJpiq33U7g15ft6PG5uIfbn/U6Dt3g5XtsCT2F7S4vRsxpjCpzJi7mD
DkXIlFZHgYosLgrenFrDkrelLYcduHPwGe0n3EP90vvmSnM32xzAuClguuaV
X2he7pDw69pZJG/UyJkYRr4jPSJmJpmJ5HCSOuTlQA6ztorvFBCE17mwiekL
IqX69tfHKD/RjNRGzP97rf4ctPd/YUb3Ah3dV5R3gCYl4YNpLj9oCvIthQw7
/Z/QIvBvFFwt7ke122vroCCR8kTdAMU5Ee4AVCumq6tStBBpXFF0m92IB228
hG0eibsWonQqtVqkK5Y8+X7VI3qxfDjn69O8y25oIGVoqDmjLvliYDDwUuUj
WpGbwwg1HKsl3qfvhw69WPxmoezy2NyTq1et2KNBKKW0H3t/6JA0/b6xBRHT
Y9adQIl9Cy6vsfaDXdPlZbCT45SGNgscfgTGdZRqd/mEFuHPu3ydRUkG0Wld
OA/FuspDQ3Y8TcwJal+4cJE+m21BDbJjLVOY4GGWt2GXhMDUVhQiduZAePzy
Gckx6EIdPoGld32aRJGZEUPThNtFJFHMT0HiRfW9F8fRwk/7r0yVOFTRfLvU
hq+7IsW97EcOkO+atDCm0X8XqHzLwsbJWZLFruMOKIV3zSqFuqrhP4vNZbbK
CYe5+2o8wg0vYh7JOYFBZLY7dDrht+/BVTJwvsukieQrkJDnLLWDEklbBe00
MlENKi9B3BWDjiRr+mPxtw5hyFtsRD1pIfxOJi327qx1984b4ap/wq8Xhtyp
3Bc6FeKPgDx9EAoeZzsnwjHynt44Zhizr3gFFDVRSNsbl29wvbpDvj7Ug0Fv
YwATES4TQBNfp3sXN96aOpWoloO7D3/EmtVRPLo1iL68N4kIiGzusbujIwu4
9gPe74hJjqagKKtC+GEGQyB0spnen6JjUSTKAI0Jj86GLgAeivvqnE7kHN7H
6XtDa0BZ/PoxZGDx+TWwCsEJxoknfY+Se4vgDbbRO0FmawtDsCoda+8/R1kY
rAyauXANB8BETWx3AhjaU/meb7eWG0BQNgKKI5yus2NgO8ddny2moLelD++Q
Pdtl9WLsiS2tsAvbOGDkVVPd9JPVi3MSMK3Y9iTwArDTsitNd6WbapCeezdT
TRA5MXaIkPGR5J8uKoVJ5mSybeWXjpWgTNNmUPVX09vxSo/LvBwbYY52UzZx
5eaa7ShsCi8iR02W4/effxczeWL8oOSMcgk/S3J14XpwM2WMXX2nt/SomyO0
xFyVFyv/wrq8XEl5hP5fMRcc7dtrrlDq4Gp4tBnq/6we1aMDFeYTq5Qj70qR
o3Zo7jv8i2C1uJ4CwsNuWyfq0KB3sqy9nuJqo5CD4Ul5S+Qr+GMJhzv1MxPC
bcoIBENOQa8o+LwLVekBYFYdWhgU8P8Y4oWguS1P7ccfYR5YioMcwE0blwSr
gDPCx/eObF5IYi5ABIstbdGt2JuxaYil6y1XP//E3djwgnqQ1kq8xGaUGLby
0wKGAvLyA6DIliyiAlncuqGHXhVUSXyrUz/rO3w2uT7+zLkS69IOdUdS90nr
kX3y6M3mKe1rZrFJNZyXB7BE3g9PQ848kwaRHSabGKssIDMKTdMVtdeT0lZv
X4eOj0Lu+zjLqd0KoXefyVBv367JKF7uKGD2evi8n6gkc3AROCvqdghrF6Z0
xNmzQmzkkOmIF2ksBkIhb795dCS1fvHRfdFROYi+AUcc9HvApVVKVMdFqcXA
3f0e+LvK/keApkhbxPje5NDtz8kCst1vyy7igTJTCTYw2Slh+1ABdEeMx24B
sTA5Juu6ymCtOyg3u9Aeln6uuL1MwcK8OIEZVeCy/cQQah+mQk18X31OEzq1
8bhVEYzB9jfbNiXgrWG2RdO4qCyQbJIpTQeWMPrspD6yv32981xPysfkCEBW
VBM3W5CM3NskFFRAbR2QURWs5yocTzAN+ko3Qa8g5OLmGH6LYhihHHnBW/Ga
Sr7aj3ioFb5AQkPbLNGMzrt7cg85IKq4Kq+t5P093Rg0XsxAsbJP7lAsYauA
BhurJJ+QQ/DMrHT3OXubHTfZLENSRs8K9gL8/VgNbYeVJKr+JbodtFd0mMNc
nh4pbrQOuyltQnzHlaZq81etOyFMkjCcJi+mdGY+4NM5DiuF5BHBkvMej1EE
gwnlT7l9rGYlRTfWLAFi8IXNaqWrvNhFcmk92EYu1uI7IKBuy+mcpElRKnbg
498F/85ft2wHxn/bCim9BM8a0ULf4/GWOLNtFppc2FW082n+ypnl8Gx2w5S5
7x8UknJFCB5gnTXyJCSJw54zj0wjQVgZ6SX4AtG20d22Yx9/RQ/gIwMBDnQ9
Wu43S9axT5Rg45papr9PgC9gRO8gwZ2+13xBunZO3pLJhN4LYUxS5e5zHatH
3MDjAMOyUQOd7vk/vXiDvCpZ1XXFTH21Ujq3fmcvJrPiDu7DVevVWT067Tzy
WYslQxuaPvaCbOTVgo40itUlFOL392p4B4nNkYJ90hU+KK7Cs153V1pyEV8C
CQUU+RWF9O3ZnYdomEZdNyzNQLUUdDPbfpyWyPx9OcFHd5QuBD+M0i1uDK6g
1jFHXgFolJCh/crPzAms0llE3F+wSpzxIDuwF4OFW4l/LOcVU5j1o/SkR7yY
LdYU5rAUjqguWO/rJtwxtcwnm+jWCf7spE3xdAun5m949MWmEuxlhjLpeV7q
SKFH7IIoUa27qYTjBKad+LukxCcq1mriSNjua1EkhcNXc+pvWyftRN3p2S+l
Db312nyRp3ySscLkc3/JGXyWRx8mabPs4aiWKVu2yI/GtdxoZHyPXOJe+kEh
47w7puqAMOZR4BY6ORGO9nyv+SGtZrcvMbJU3vdOgyzIF5OSaYz84FPZetbW
Hr/bYB1/Z6wbuWrsIRvRe11P6GRlez25VCGXC00HX3yM+bZq7MBQZZN29noB
LvDdkmz3zxu+uEqBY7kqEUAUEA7adwlZIdwwio80yKAaqhOCgqt5nzD0L4IX
RfCMv24Kb75KFDQdG70xVoSDH56aMvbgtuM5f7wptCGZW9A0QF5RQNuLNRaJ
AWyi1zWCO4iAO949C6hcpQ6edDq/EnSSlfaeSZYzcTq+2tVlT+fUGYK5163M
l/9zEujvHZNedEfunhuxN0yD1RNJt7y4lQbS2X2sSGguBBnxYrxLazgYFduK
Ei6qt0SycSgt8XXB5hl45Vw+P1ymH9taWbv/CzR21c3iAzw7QsYsFOJgbPar
diSu1vSXqtGzOncP85JJTtkoI6scJEPX32fYQq2SjmrN5V/sZyaGJfz4qMEs
1POVE/SlZQ+WPutE1S6xc//kcs3P+SiGrcPgG05jLNDy0JVb6slq8t2S4dO3
DbkFhWF64dq8W+FMiVO67IH5tZ1k2a3rE5KW3zh/uTmIW/CHj/pK7uRyKQAd
+m/AgvPdZ4IecFPfxxggOCb/5FrbwFTSPy7h/niXPKNdyXRPzMbcXoi5kG9K
gI0hwB0RN9JzMLJw/R0R7RMrzkRfbMcggqyYjLJEP4/S3+SPVK2EoepB6TVK
siJESSE6npu8FcazGkqNjH/f10jpjylVw8dNEOIrhcO/67S4EggiEuzEjFzu
/Ub0EKsl+Gh4BS+qVsLv1GsccMGWofT7S9z7GTUBX2RF/yvWn8+rA45vw0KH
IJyWWgTZoxPGSD+4yqUPr3ilNnM4ns5fpsG6T7My3CV3HvcS/L00i2xM0OUQ
pSgFdQq96DH/OfJLzItIT3uHjNqnYkMfnpksNHid5JmT5cVVxXyOpETQsHZ5
MNemrWKt2EfqIwocpa9k4Z6F92ya9kW9FHP5C4EE8Gm+KU1KntIgzOUtDIUQ
0DGPi/29ilGnLnZTBHduLRAMdj0aPkiQCBqG76o0EPV7JnZI/SO00fjlPFXy
eVZEpBqqlsdwJDm9fe55HkMb3qsYV+Tc/GmKaGtFOh54nnzoDqwnntz26qks
Pbm7KxzQ2GSrVTKz06SBu9G8qEaf7ZWyx/Jtm4gm/o9skqOg1ZqHO/EUxtGO
mvg8Vf+hESVYr4nMUxQXH0oju1kPa0IFkQPZegvdEAqp5UI3UoeZghYXi5bz
OCYJa3HFW3r4M70V8B9QOinMFVzpuSFQNo1OL2qoGDH0Nb5K2ne/4CA45csc
S8FFv+TXnoA4k+lzJhexo/txpJMnyyFlR5nsvXSwDQyKbtnzb9xnSWEtEngZ
3vCtLDxRLHn049A0N2M8WrstelnKVWhSOFgp0oGsjfaGpsNrRnpBeLPofbiS
+cc07yNk4pak/x1b0g1Pgr1QYgv/S2RjWBrtXWsSrWsitjjWiWDQLyavpSCd
ogr2FWyAS3QwobLXWe+lten1rkSyqgrUAMHfThGk1erelbPpO2Z5RMQ8DFZF
x/x2wF4X+2pSoW87xe4a82FRyDR8rOZsCiwbQp/7fHyiwC9de19JMenj4Sp0
N2jF3Zp6eJuBKQ3cEYBmkPFXggTn3GGxY2qLC7qOB2gODT4XT6uirZ8SaNgr
eTyiIieZwFTAfIppESq+Wf5qOXzZsNN925/w1C1mQWqD0a3q3kBrQvB+/DSA
C+2UBHiC43rPUxOBiGnhUqR4WQEMEQ1ePcQ4Uzu0oyJ3SnhSiDq4AtdX0zmd
i8D3jxtaG/g0uBSAf2X6h5Ya5CFnf716rjz9S9xPbD5/u28IvK9tXGrs43g1
HBBX0qD7m4bS5qaGQG7Ma796zYPJkGSfLsHnBXF5JcL80zMkDIZsoMPJzl5J
JXTJhKPmPucxy6nroIwx+w6YkjF0BMalklachvRf5vvRRX6BEFOh0zW71fpb
u8O6sTcvWQubfNX550NmI+Oq/hRQ/b51YWtRmkWIHToKR8XJIC+JHk7UUdGQ
R03/IK8r5WcM18SZ/GJAxmXLA2K+DGMFaBZRudOvRVZu+LmNKQvLkk2sZ+hK
lgsw03SL2oi9d4tgyhULcpn2JJj82b6SVMpjjxX4RvTyqDx289AFOlM+0lNt
FCXAaYuFDJrPmAwGq8WNQ3lrFcTr74UKQ0gtqdcezW10EjDQ85OZHjFOChYC
eUU4iX2f+iiEwUyJZbhUHxQRMWGdQlM2OGcK/5y9EEun10Rzaiq53s83tety
5TA2SfdmFN2mcTODkUbEtdty/POkQyB7R2hsLxxoicYewnQFB1R/59qVboZI
2/tsSJSz/XtLMMqfqx4vNoedqm3qxeamKxV9Ul+Nr5Dp+A/VG+X4IKFxdP+w
mVdYx2Z5FcZcK4uXsjSx2atnrk0B9tlRf8X/VWuav1DBMhVHEsYqAPJFXOxx
HXzPlxPO5iz1v2VZO72qxk5KFhl6/TZFmPEi6nL/VtJtql9+kGaqBvn/zt5F
DzMynpMxcMYa0oys7LevnPpXRtStJc9BbMNNmRftEYQTDUyKGul+od+VGSzT
w2TMdqmsfKoDwTbURCBCVH/G8U0TOTV15DwbC7EebH/zlSyP++U6P8wVwSdO
Hdky6t9PyP7RS5GZBhwdEZJtP8GKoHljogTcnit3YSF6jpuL8aj0BpkEvjcD
RhTcV5TpZiaZqlqrJ1AEfVb/yKRvA+TvkImhKyxYXn5OPok1K+n5wX3G+jhl
ZQzJBYK5H0L4Do6dBki4VxWpYMwiEq8eOPJ5X6whJzNqb7cI02xfPHbVedZd
CFZc6yrFYdpw2Xl77/VxvhX8gLmk2z/0KGpRtUXzRMYq2BtxiwfniT6hjO5y
qdtzbSgMO51C63oR8ge51qz83EKWPWJhqZkPGMDE9/2AFrTwzNbwr5Uvbh87
rsuQ81nwzJLH4CEdkKnnWkj4GibsUzecORnhfXgFBTFm4kdeNe/YzfIlI9oV
GSux3NYcl8DTsO8m6uLsJvggpTjckEJt8uuo1ij1pDJMpIzmwH5EoE6ZxHRo
x2QEfzO0lcqir0hiJ6nsgYhgIZQKlAqS7jSq7ne/yMIoIHOWVZFm2imgSh/w
C/MiCJWkv8LRV5H65Mk+BVS2cAY8u3PMraIUYmzg/Ch8B9yAssKxVP9qj9Bo
2aGNWJaAcPy8MPKdxNk5c+kmIPDVjIwFs7oCLnn4wnX8VUFJhVtH7Sf+iXvY
9erLVY1kyniMMxrO6ToiNlHO7EafKVeO4ywcMnCDCkDf2gwZEF5pCs/Fb22/
WFafNNrQzYZ1g8XME3x7ie27eJjb8F4Lp+3wVWMx3N3hjqEv5iIyfUhghsVs
hX8Pe8vVe9kjZsgNVWEh236Nuikw0V2Q047AHSb36t2F0bIY5E7ndebndqyl
02wHJME9wiwTSpdQWYRza0pEyskmn6gwx3sAxYTrNrD8GrNNfRf+y6CKEVMU
TKFj3qrIBH9URXQ+QUkk0r/9+HXcMSzNIeezIFO6CvuDFhdPvZzgjMGCxXT3
RNQoVaMRrSixqfS2zSyPTc0/oJP4V148VUWkOCYfU71A2KNO3hXe749td8yN
fw6p67VeO+01jmtQoN0RB4DNldZmT4U5hIEN/pLFo3++Arrva0kcYkz/lDHs
c2KuJeGio5voMODhidDfbrRw0dC63UDPPk+n31z+DsQlBzcbEzZrNUlgOEq7
tMbF/ePoHis2kV5g2Q3p4bGgPCOLE/l6iE9ByVDSDcl1IuLrN/a0QZ3SMf44
H+5x51SOv4tsXOB8ixLYP+yfdVr7bmJdTFIwVQ75YPxY/hPU4Yn8hp/iS+uB
KWothLKN8ekmgw7uZdJyCV9tGUBTDqC9BnXeM2bHvOQSgAZo70+p7Q2hJ3+g
Go5A3MbQlYDdvsgn7PrZocwsXHz3GcnVUnl1vljFdGg41sYv2yf09Wg5Jrma
lM/ipA1HZ7ZD17SyEtlarYgQFgj4Cr5O+B5IU9EWjefFgHvFh/UYRNpKNReX
SZo/VP4Chi0fEDkbWMiYbZE2R88oGtKK1wyCWzngxidFeSxHpNMt8YN5bzCX
eT+trlntdHENoNUvh+i6D8CwtVFzGPpAjVBNvYy+vKxG6DvdZaE0sk+9C/yl
YhGuLIkDUc8aNqzHuRFIiX1PLWTPk4YUK8oBPqQ6n1+ajLmgdQFNzY8/6Svm
V9oDTKutKEIhQg7IRTtiqTWFCDCcAf9k5Xl7TUNy1o7w9MkErxlQBuVc92qQ
kp6Axjdy3WAXwVheTqR9pxsxV6LjmGohU/lO0Re2NdCqTxwbPKcGjdCHpLP/
XvEWOGZPkXAIDvcUtNL4zElfZxyNq1tJUK25kyR0GK6oqHBAw3vxqnax1aoN
012Vlg/CGyIcQjosNMKP8ez7cKXBFw3RSZ4Okv3ggUxn/sIWEeWV0vaEamlz
Zy2SDw308DcrwQKC+YBhOe2Zltcx7KyRnqmBei1F4ochVfPER+Ra1fOgoi39
0YiP1HzXFp7vhDobSyU8hCyzTN3xdC9A94+DuyRAtlELIlmgLjZYRImiSZw/
zxtygebxMZD8gETpF61WicV0c8Arko5WFWm4Lf/yMFBqnRLeSAOYrqO5VofY
y5KxXG7jaT+ZKIfCIzAXLAgJcdehOIjjJelrDn0MjZiZR3a2zw1PvsfQaELt
NCj6BjmsiWEAwtdmLw2Qm9UF04Uw86g8kKs+/nr1ALe2+sxOhTBnF1/1jRs3
GE+mie90sGUU7AUra2m4WuCXQg+DyD97jmCrKz15X669cuWG2wYl/ro2nUtX
3n28Vxq76jt8eT8slMlRkRhpW0KQrzDarc0/NwJZxcfHMtetV9oK95KC9rJd
CWtDGBf78KN0G/1vt2aMQslcawRFGQB7CqMO5TteisOUTdELEqtDnNvT5mXj
cUfDA2ZWd2VDd+vbRDvozB/u2Df6QVcEytLnZ19oEBGUjAU07cYJHK3laJAc
pYz+lqI8zcL/mZbgby8NRtX03XnrDYznSp8wl6tX2etsw+RxvKONzAJJVf8L
B+5yoqJZw9j0hwEVSgtuBt/u2bX0V9gwCw+tcttW6CvCVSMmDeLkWP2XzZEJ
hU+ghvHk2QLWPKrMKUYOsNh82eD+rx203xBgFtiWaeHlcKnhdjs/xdx/sfKq
EV9P1hjrHAnBhmmccT+LfvMXml0CRISfCu5kCffFHJZoKfViL3XaRLGKVT+x
pL/PvNzSgwuaezEojQRBzqEt8ApX0fqHflfihpBRJ+YZjPHTMl+Ct5iEwn/D
Q2qgMwKAkxdocO3pnEdDzG+b5Bvbq5o+PNFY9ave4QPB9x7gWfBfJ4B8ec5x
0x+TcsE13YwGDa78z1d29W9nhLGD4/pNrO1gkk0Ezx/otLpO7iEB0zoBM0hE
2BvdCC3jwlCQ9hOTjLXfcE1vnIFDBxgQlBRNnUWkPBOsmaahTxIUY5WGlPyR
+qEf1YI6b4HrERmTc/k6XgTpPib93HgOiwPZm0xL3Mr2oJa+cPiIQXen/7t7
vGdNfUg35ET+av0vqw5zNRoopiow3Gx0ZWKku/gj8FyTXrydT+RdPpCAUCVx
v9bP+W3Jy9smx/JrjgrqzfYaks+14npz7VGXrRb3jl/3KEwKzbGohZkoHTtI
ryE0RD7Ky6Fi/v/IlKDyVvvTbVv41Dknt+iCVbmVdZjGKHNRRgxa8JphO7Jq
HG0Dy4mvMUCLMqxmn35jO8CvhyRBXIYluAWjbn6x15/+0vTcIqbWDogG5B1A
9KriefgL/7i9puvtsFVOooz8TCwEfA4OI5SVa/eUvOZgN+bgq4bMqR9H80M3
os3gV1AVaeqf3mLezWrhDY9qGRf+UWjcYJ/cFHOSv/zQ1WxVUjX2OqvizOgc
ojr+lFVntdBBnakPqQUufA5h3vbgAXl8r68LYVA1UZV+Qu991OGj62pRu7Sx
vZes3Sc36wk7XmdhLCxapDc/F/xbO3oEV+CHg6qyEa21YqkVHS+J0wfc4v+K
bFl4J4UvanC/E9ECiLtoiqs6nOy0zLQSv09+L/7UA8Ncj4AHo1xpStaAdxYm
27ftfZXZh1O3lCtQ+AqyRtVzuvIUAXeo2fp0z2XWvBCDkPZP8kZwemVBb9qk
uMxuLZVijK2NhS0HfJzP2sFJ/dCBKlPaIpwyA6ksr+u7XD5r2uboNcJ4Bgzb
KIfuHeXidfWM9ffrnxV+BA3pi71NohBCU/9HH16ZWdN1ijYgF0ItG1Yhlqdj
7HOGxLtW3BgxmwCJBlkapEQGRjYomvRKgSHL5dtDWcsOGmOA6Wgjuj4gCQSb
AEtZuiA5kMX1q5+879T2F8IEKxIcMIlzqkC6lRrYpb0MIDIcmYRhH1JZEbLV
7u917u5MY7Ii66Fpovswk3/eQsnji10J3/CS5uDutWMjptctllbv9HibMqF+
TyUYUdZVwPuV5g4XFW+uEbgo5HY4n4IuBIQVhRVlNTb0hGdVMu0rSMqERfBo
5wBNeNsvZ+84gdRYkt8WpfS0VgdMnbfx3d/OFsY8s0dukY2Vdt1s9BZXvmud
ghO4miqHdUnFgjwT2Rb0UIA2eT7mv1IcEOz16iRtQCrlgO4dnqvwG9qGy/CC
aHOgduaW2n7eYbIohJ8RH1WNMrm7c3aWmYb1wHtISIU/UcU8vTzQ9EZjCHG3
iTSRTTCgVowu59ROGHeiSBjCDu56qa74mrPUz8Pzit7KOz5nNnTn8vPsCesi
my423BU0vGt3bIA/noooIQtBRnijWNb8+F+KeeS/NRkY5q841cbAJgZ3bxwU
FR6twDrEiBA796ju36jiJklm+gWZs8UQkM88fr3nxM+q7RoNV1DQCSQyjkCf
JdOeBvX2MWx/8rbCFos/aj0BeGZKEcCSSzIcEocYyLoU7hxGLbkyLAmQl0qo
wGH6rIicrkSbfx9ghHoIvF9YF1XAU4XtAnijKqqfeW+3c98EWFSVqgFAqIyg
ZdytexW+Q1CU7OZYYfeeGezRUHIlmoU8bIbC4tW0qs7BF+EJjInuta4N3v5F
ebs5lWcAtjTSIvlSqTYvKtwjF7xabhffx6Gd68qZsAWpY1uOTbtS4di76Chs
LXAcciVvMXfRcp4WdfNWxgK/lXbNDtJ7U2pSYBDMQsso+j9+wgHRknsrxHH4
/aSDkHXyv2VJWxyEFjL16YtE0V6JdeYq0eTkzzOhEBTYyJb2JpzcDRykOWtf
zWiM648RSXHZa2DJXWsxHt8Nnba+hyzMuTdZZKhBidyO3VR43Mubl701JJa4
RONWgQT9phhPdGvpu5O03VVAaR0TeywWf3lrYhDsJ9HdrzH2L1QWiF7qWu76
61IOlUE9ZxMWbvhhdhXQ5CpAL1r6HKHGZtTXYAAOQg6PiPKQPZMNyTv/b9DY
jO+0hYn0Qg+dU0OYbULgVBSAx20zfnf080MY8q483+rL48gV+fs5BgKWxySg
tpEppTRj92bx32+jh8GB0VOdbkYLBszr2pGRkKVJEiuq0s2ugzr5d/8QBhTq
S+10E/7RDD6xNO7YiU2vVX7eFw1b2jToYh0jtfQQWMcAPyRUULGpc5Do71O3
XaGFt78+3YqH1D2oCBVY0Zc2ehTE/gWVxtBGf1L4uB4ON1nRuBd8og62dLVq
kOKAmKM6rJcCuemLDc0n96mFZ7C/GQLt0VpaijynbhkGuvDHxQh86fY+x6si
t+XkPopLDHbeZRXN7thKnGL6l+7z96VP6RuJ6CVeJmWZXpOjp2iWdhQgudnt
N46jH5iSfOyYiPhIjVr21F/in4g1MI5QcyVPWEUOTHVDePNIklix4btg8Rac
SzrBq46ficw+2TrvgPCpvJiyDLVNlQHDLEptVE90mAwUOMmtFKhAYNW/oa7B
X6ZsgRI88QvMdxP/7DFVPWsj6QJoTy4Ig9yfV3CJy9qCHxYH2wE2JlZC5kII
Pk3goGMWgOSHk7NujeDNASXLjNRZPsuP5dAd4SIYQC1pjBNMLXFR6BtOh248
xsoPHRQeCTxSeDCPlzqbRJrkVguDjG02/JAJghzutEHFByCSSlxkP+TZ3WQy
6TmfUJQA76mSgvi1hRs48sS5puwtaBThV3D8ROcA0urKB3VLvXvGx4sPjIYM
aQGRFSQXUm48LXkgPlXqF/d13CEONLSJSslBn+g6r94n1m7qM8GPX7Saopvi
RWO8aI02NEiHHosigFofL0+vC4+VMzYVydYq96YWbPsBcIeo8XDq3enUExmW
vY72kTDVlYqinKYUNF57Ou8gVf9vhQ16nRWOIdn8LVGLONayxiVGHciDiUEp
qOmAaDfCZhPadbuMKHdOBmXHx2JvCEsDv3Djl1XPmLzQTA5CfUh8jdaX0MGx
pNS8VnmhqH4niyYqjx0TmRoNPY6vhWP/fMjm2U9txJF0jIvaGL3/TvZzhSkk
KNxbSTZG/PcDyf9eb5VHDMa9nZrPuWiA6iojp4nBCkMjqg8kpqmjRXz3bGB4
EcABiovpmMei3Xpj4Yf4atwV/8zhaoRTWxYPVLaoByR4Nh/6qErYFsVjIUZs
rhEMsTE+ZfOtDg81FdzOKwN/t496udY4MNJRGWTGZs4HRIQYSbCGO2tF+/9F
ElEie3euZiZ+49Q5Reg2laa9Cgrw7DWZGWBKqVd6+rKbrAmRBYGk3I/gC5Uu
bOz+IGAFd40BNAJmKv6uxQq07O5dsBBJ/yC/atsTDGA23lOP8pDy9CGrVGEz
+yzGGWJix1jBHJgYOVt9QQd9o7rhJHOt+N0S2fJckoU3nDhxz7ZU2aBG6NZd
9DelDoOvDss+7zz8XMd9fv9z1CIcviHz+lioHAwygObxHPCZixz1bQe0Eiwu
eJTjTivSbWYeMLkdb8hGt3xnhb73/1TPPBYf9glkboIfqviFdGkdMhll66Gt
1TN4dPJzLJz6gkOBAZcrbglgOElwzbV8Hsait19hZt2LQvJ+Ppu821/ePA+S
GoK2xZKhJ4XqYx0qXbEG+1f+Nca4qIR4E9zpWuwFjFf4muQaUTxhTu48k6oV
TpWntSM9Jjhv5uT1DWTE/llMSLUZ76SxvoD6SXiNE07uaJfDGIlhkiaKC4xF
YLRJC1tiPQ30gRqP4iMjif/hQjKt5GWy6fUIwz5QKnpYz+YQ1XjSKEZWaF7q
tY0VfXPZqfywqWqyFAVkrjMYPfeXmT487ArSbT7/ETlfvp1LTGfa4/ctQaL9
G4rA5jTjSzdxe1LsnnH+u3xKpHf0qkGe8qcBMhQePHOgRYWGczGmu5LP3gNF
ZRdv8XLa5QcVe+h4K1mu1Ltwss9d8AdGwvADAL2ot5fYYFhcOFRcImqkVEt2
3n+lhb/u7qgE8EtfklEWMW3S/frISenCnYPE7d3WFLaTAbNIBxMp95rN0TFd
DmpNqMDYB+BmoGEWnQr9cqN3TbLsul50iCCXhyCE5zMRkdAv4OnUFgnQxxUU
+7l5bPpgR74yiDYyUI6EWpm2POVM0GCw/OleCXJfKAvZSzn4djFxv6LFtlMU
BguXep0rnRFeLFKdaHV5glKYHFEB7d3Zfq/7+3dJeCI3dZRRxmC5Yb1IqIQT
aJmfE7GQnP6rjUf0DMKb+Iufe6gmPDkd4AhAUFr9v3nAISdPT7Mz3qDRqoS+
HYgn8CqXUZokkRNykfK/exj6f+WKZiY8BG80Hu1TTFXuMXSUP5AS7dc4e/GN
+1HwvQnib6dOvNQcBKW0Ao9FO0PwIMuG2H0JI89UJxgJVT5+J8pK5/GN/CvS
eW8mOdIgsuRgmmQwNAuMyi2z/t8/wE4v0+zZqSZ03t9V4ajqDDYEFkWwxzzD
oc3/alcCHhufkljDjg3BWZyp65jCduLXRpfkRIG39Y9qhWparVmADc86JOs+
Kqr5BUiEQJP7Uf0hMXsGkKmoRjx7P8ZeX241omvNUm7afpW8SjSp2H+qcKcG
wUDJTYzQob5jl8a+8hA53L95ywUESFeYSTvhT7lK3DgBuBRuazuoK1xfkiTH
IFbH7CLZBpyUTmmGFVoaXwcUtNOwgcQtKOj2+am1ylixsg6cE17DLn7jvSKJ
GZcdMy8nOi7Tmq2lz/19R56rBcmRHLkBH5m7mK3XhX5H4DSTiV6oPxorfXAO
DyWMBe6WkjXMqgsrn3AG1crYI2zS39GoILlVs3z0VKiBlYPrBu2/D8DE8RZE
Jetb1paF2IKgEk31cCyKVYNKspz7JTnLzzIZiz9El7hu4J/eDQ9Mn4WLuVC3
2zAyYyxcK10vRNOnZrGWIrtBFvrhGL4VDRGakEtsoqSNKM3gEZOjZk3xWgQ9
FWCcm+cpdJX+WRhbBEL0JtyVgSElZLN7eLkwa0mIoiXTqgatmwhVSfOoX2V3
KQpj6jprCdNHfnV6Pro2n5gavpgk1gZDMD+uG/C1RXVJerLLTATFT+bdw7lG
qolua10iZ5fY+w/m8Ql4+SYgfwuTRvwQcBJJul4hZl/vMa0Zm/BZTZ2cXN97
H8xGElDIhrBT9K2k7N8b9OhFvOtFHsKPlDlyovwc/Li6S//huqRCQspPjO1u
GPv7YFwghvxIZkWY9qAVkSVmlG+/ZF0xK+lcgZPtJGifS5kiTEfUW284j0es
YEgApiOuBx27h9LxefNueVLHqHomprZEVzrMgLiJthVfbepSZf0iPRtJTCcc
2FJ7hCbGDiHxat/oMew+pFw4NFTqGDTYrYDtq0MTf+ATEWSgVeIH4oJWO9nv
d4EuwuDzhi9+sSIKxDwNOoYJxeCMSH5PSNMMY4F90bOEEIlaT5rYM79/falD
5vqKUAMYZYtsEydl9C0QDYiiKMSn74n526TDxrcM2Jz+vDDF775upYuWmEsO
PBSdjaTFI9cXbjVlXfRFyWhX7vXXaUuKeP4C9FLpZJh64mmBkMdXCCF5Jnke
m5k/NQJ+fFGn45SjahY9DP91qIwX19GrOVNBclNFu6/dcggfqCMb1c3DgoQa
eMEzWv0j3IKyFpWWD7VEsxVZNeOmvt58jxjCd1Jcw89/N04y5WOm9mr8qSdP
7nEbsX+b5QKZ5Smbkjeaqjw1Wwg1lFboL3kvu3McwYgYb05Xc+c0oufacKj/
KqvSC6F6r4Ur0Y+fmEdpeI40raTNRFgpmsDM6768/qrxQgVouCMnYUkpXWDW
Wt0fLdupYKlVKyE5W/hZt/hyLfgHPgV9am3V9R0e9wFjqgi1ycHrvA1Dj/71
70TKpFs40naw1FvujTkB5nveqBw7FiY46BduHlK7Jo11WNkbp4QPise4Mvik
sqIzmLoTEUeH+/HCHHFOc1aYfap+hXU+onrTl1pJHJHWn+imn19EOUSQEvjO
pnBSDTUxZvFCxGjVD55VVSBvR0/ouquUL0YqOvEW9UHh09GhjRJN6UI94Fcz
eHUKn8TLLuZ6tdG9R3cOpHTamOENFLCGz5MiojOlYfzZa34KPGgYCaYgiab3
zmQKvMlcWlxkWwr4a/ZrliCiVyL9n/L3I/UYv5UCqnbulLgxUb7513Q8COp/
rdy+v7jVcP46RSmChghSn3vk1Gn0L/KjzMPNVaKDazAfTRqkpsvD+5hpNmp6
FrFEe7aXVaFRCt19Sxjnsw9WXApNGWwQb0cx2GGgbunPNI7e/hZExb+89tDv
hzTMTBwsmdhKfvuyihamy5Vlld6RZMIJ8fjzNKvbnoCei69Cex3o8sD29wpI
iQNOZD+aAhFYMwvsJKepTyP/R5Z2BHIUfOCSr4irgjd735yFnrfkQP2XpodE
A7d9etiHXUcmp8vOGthwKGmaZ8qUqoACXqzu5Ht0dszvuN5cMyyBSbrfh4fi
dmoQQoFMwqFuIaHPXgW7eQ7pYAqd/2tpClIFEgmMUk00RGoG1Y/1fe8iystf
fCzbpN2pHZqa1jtxiHFbm4o/aXoRseBSOdgdfA8y2JMHNOl+1tXkngOesMZe
ikhJKcIBFTiFxUx6wMtusWHYcs1pVM0OE2mjKUKzikpVw7dW2o4Lk3TiwCkX
UzCccCpUT2yAyZ47/UMG5rm73BjfGIijruP5ELDePTWAehF4i/sGvZpT7Sqs
xV4B+ig58TVk9+nHuRsdk9nIfyY/tO404hwrCAL9ItnNCxrcQQX+jnoVvAeY
52mZ+spJMKOMnmyxyVBCpS/dwk8Mjggy2eyZYnYoe8yJhRlJth4sS3qmNysU
+w88B8K0PCqarDKHRy+Tkvwm0UjMCmq7JSieLvNXx4yJIaFbFrV3gisy6fau
bdXsyfhs0uompIRLb9WLDCDIn3xfqBdmaaBRryiBLje0mSAWdQ4wZJeEj67+
cYv7xOvD0HUfiub8hZyb0M52LN4i7SIFh8QiBu3VAIsqgdnps8lWjf9eoWGA
av5tx4BIppc23IlQuzivxbkpSuADhdH/hb7HEXqsIbfBgytao8pIapqGfvhn
B6QTBuYqaz2U6ZvQEJNHz99ghKWuklOHdnWNiSY8362+gmZgs6wSIBsTg724
/IWvM1Vpwwt/Ov9EmEdmKkwcsbqKwGPHI04HlNQty/R7aKakUBbJKxAxURnS
+A1BUojg8thEqPQQdL1yEnYhGXpAttQAPzevfwbZfTAWaI/aUQHce9QUw/OY
V8QInAEuLyeuGJQAcj/yxO+SgepPr86u8XLR81AWy/50zI3gHsUFGj7IbQ/v
9WbqBK0DYnSLUdvoIypKnU5PH0i3+VrKZk8QLX5rq4HJnMPx3ZKnaiQQsoAh
qX6Zw1gWuBjqRI9edxCb2PxQkX1cgCSqtmZirdBEH+Rs2YM8pTUPi7ISlVKB
a5ylIZh+aS4sL1KfevGx9W2OvAG16HQpJpvHiuAow4XNQQzwgmFpNfWUrEX+
IVFWnHiq5sJ2XZ33qjzM7p0v5oMM4Y8mpv+hNzz+r+TRGUB66C6Sqj8Ibc4e
gHaOPrz0/7LKgwHG3pDXobdGOQKbgzI+dqyuOjU4l1gs7E2l4F9IkH05YVSS
8ysRJPSvP1Ai0VQAT8mJPSwWrjuHkIYlPTa4f/RmVA8auK3hv3w1iBmg3YHd
6h32q4E1+ivpiZMriDVdMhQN/YoXwaXPiVlsdsyHp05B/XhjgY7ICM+yx5Qj
CTfvJ4rDk4SLKvpMeFkltKp2XiS6XX21kyKL5fKV5P8oZvEWTtqVicXKJ4u5
LyN8EFioc6c/vAS1CodLS3tH7TyLo2xCUb71eCcpVV/UhqljGyeCNaNVb8o0
0vYYpr3fEBbrNfU4E4tTuTG6wtqoYwx3b3XjlBOEBJEh+8N/r4xBAu/0QyOz
Obhvp8aCHmJm9H1Nh5qBQ6LU2H8rgC40kmdU+noUTqMloZSffHCe+FWOQbon
dRtnFKJV3FDvn3YwT6UO7bpDDdufoRsBLHKPgv9XReaseMJ3+kONKscQGw/q
psSOdLYK3aAx/lNaSL7+qovAQmqo2h9V64dHOK5ZIdKBe1BPQ2TXhmBkGctN
DO2Tqto3lmDceBCnbO7Ma51+zRwNnoOGadyaQmOOPU3ILk+mynGt/8WUo8d7
lZvX2Bj02RQOuvJfuhpNU4K23Lkssmwh9CCnSpd4Gu/tZk49YEFeLBowkwGP
ET1UaBl2Umq2E2Wj5whluh43gTyruw7bg546g0qbWVTcAtb86LlU0ehWyqfK
PYxCp+D6V6IQiyrHPxHJ5/OahBUhcLvJbEDn52JeNiXPIaaOJ+k+SE9za7yj
3GMO5vAEEYcw3tJ9Pe0yPemR6ZMRYcz0d+FspzbYYUSCHYdQmi9mYloi45vk
pVOuVFYw+wIwwg0tYOhehRUjs8on4oNg92DnKn2RwVF1/fR/3fBPvwY58Xqk
1XZRSM00hdMggHDqQ1QW6vL8uf6qrz7Bcixj6hp/3RpU0M8G8sZMZBb5lh6m
zYArrzd5ncjzRvcE8axUKFajFDioCqWnYCr8UjDHdjrlIkwYYFaQaB0k43CO
Ccgli2gYF2np9Y/BSFWHwFBVLDk22+GAlUCYwaArryAsti8kaeK4b2ztyw5v
0B9vRHvZY00UPrMXyo2dHuiLTmLgYFo78tTGXpduFm0nQNgZ5gBuLSUgtu3S
A4S/tbvyuhE4Z6Ev+1xVrv1pWMlnvqeGGg+AXhJjJlPar30e7c4aZo3WjRTt
2SFhp1OvH82+MDZtAYGe8sDTekUJs0d90pMhJJ6Xz7vEwk4nST3Ltuxm7io4
/BHr5OMtp7P2+4OUsU5YsuAWFpb5wjJr4jxvyD1FhBOV2/vUAojurdMQ/Mfm
l0wcde75oEjnvwNMyQKKoqoVXeC7T5wtNh76I9pp65LBLnxWAGj9O+HFmeLK
Cklvup0XykJx3YGiWSc9+35Z+cztw6S6Pr/8K/AwVOPlb8gLi7r24YYBZr1c
PqB0RNL1rl11PAV1uaKf7y/IPCICKGu/unUoB/ANPX5qsGauBjEX0vbKGzEp
Ew3ygvG2J8Jf8dF/0CEVzd2aD303qnQsEMJphyTyh99rpGrCCRL7aYHflUQW
ZueJi1jSatUe72PhaJCV5r3t0JLlfzEsLUFsGVT+X8Zf9e0590XT/4IsChsJ
AkrFV9IXg59BsHmqSfYf7+yM7nw0qUhuroiS/cPMzjfidR+G1U8ZG38Ip5k0
XgcDqmWRDizQTI9TZSEICtedEzlTugyDjmCSrhnzhpyX8NoeCmlLmiwC0cWJ
+aSwduiK6FB3q93q3lKBxqDyisuBNq/4xtkYOEzW3HvMIDuKJVmW2xCjFiMi
2t+Q+XNm/p2KHBika2N9iKRqPuVaerlucEFl3oxLeuEM/qw23AYGRiuybYeT
Tst43OtuPtNBI2GNYuTWV+KKbXe1v9KJmgpk/w6bh+/VeBS3vQEniw+S9kdj
iryjtjLHUxbm3MM79fRBPfyseXr7KW5M+D21E7ZtKDN4B/DbfH2l5wELhfTv
78lYbq5XhHddNKzM2w1neBMxAgwMGNWJcfkfsueiRJooSKlOpZVaCgnEdj2U
c1dlRJ1JSUPfeR62yrpb4llKGNwHIB/1kdAiQHGP9a9Tydb65XDFIQHzCLs6
M9lZEZ8cKfVe08SCM+VDXngk6I7RQdT+a27N8Od1M7jj/q/u26hoAnHa40xq
7K1KEnm5bGdgGcmeFLHRew5tbUnsAlQed5aKVucxEjBeSI7mL8frlKDYJsB0
9l6FvORWUnhno/9Yb+TCLXQje+CEsam6x6EYZ6JqMGZmWwBDJVc/0DDljuD9
+uQ22uyd/75fgektQQz3fFPNeTmoyF0YY9Q0W3SzN1oPw5x3qsgAI5XCtoJ7
ELfs59YXf0YlSpGbov5hPZ+KMNC38/5QqB0uoemmjMs4jXd7EOv4BXEG3T1M
33gLapNqeiyhMWgFYnopXSj8NYBvlJ9jpHxDST4ucNk1KXlHFHe2U7V50QDW
AWeB+LjdzSv8BQbengq7xCipUn72O/apAqPVDVcszJ6D5kcCIq0Euo5cU0BU
qqaqxxRyjfIvah7mJ1kJOpuM4zYryrrBkLCyD9dnIHEMBQsZAOyBxpLWcjWm
oaINbll+gS01vjKkIYpe3b6jH2Yu5ZKNDuJtC8srEtbksQxWaRna7V8sukMv
MhZUfLiXRT+gbcBGjUi11XYFAC4IqjR7I6u7TXWt9JAMnQZCtyz/esHG1HK2
7eKqtt1cxC0aXyPqnwblmQJx4bKV2VSm0BqqRrI2C3MkLF1eRYja2vSxBDCq
Y7JuwnXHIAxOuKMpuK8GUwV8pX87Ky3S8MB+u9Z8jck5pRkL5tpJEcFnhrnw
yjY3rW6aa3sGPoLlkpUSU3VrcWejmwa9DbMBLwcXk6lzC3hKhUZfXIWUEoso
t2dE5FmstKzSgynDea4CpSD3SeVyOmVvpCvQmj3rxbT9HLaLcDlMDJgKCayz
VxkMel4WNzWKOptTVo99pcNJSLVvJ9q2VonemMo8C/AlHzESNeW5PcHyYLlQ
krLwXImFpkhHIQFoyzB9ujWJRx2BEZNLgVzRfIvSMbWHGwCruU+3dkjht8qF
KZLSRGuk7vIKNcKBYG0vhqyUBnQF1f1msx+Uy8U6oo8RvkFd3A4j2LsrQ/PW
WTnfY92tJE82LoY2CHWiB8pmFcBK+mcswU2495pW8MHPNZ8LsqvzfC2JowwO
qqxUNZxWqUsj/5epkoWo/MQ4Hlr8q0TEj3cLP3I+0yJBFJTGUjOPqxTjsWH5
0i62axJQQJS5YSQWSP5ZeitdKKJPYthtqFkY0Ew5vnARFFrbM0IqXzM2DjYZ
LVG6J8enNB5dH39GGH4AYKIg/Gaqt62N0mWCziGsvi3aY0nzvjGYvfPLDpkH
vYYMSHiKZn5jQu9bpwLWDl4/NlzIOcTFayXXnc6G6VcPyyCpMt4fcjwN86ez
p3gD+ZzRKLOAveErwh9dRABLiDWlcwEvLdJAx1Q3zZSZ9gxXIU8Ui6+4xOx0
yxHLN11h+pkqDxSVqzOCy49GwR5EcBH0pgJl6W5coazwtsvVlNVUtxBi0u75
VihEO4RUAf6he83F3+Btc3kof9O9Vtuml5IybU9HC5LnJH45LySYCcZzWen4
mI/B2CuNplf6WGyvrsF7QFc7pLpGHvbo7mnpJ7mk0PMvyMMY8CqKMHDrNmi8
sDII63FsWQxbu5hTiNgdx7ej38ZsT6xuwncmSM41+Xb9cfl7KaueePd3nFYi
Ae2XKdhrA5xM8YzRcHUR2pQEuCMkj3oz6rHXaJb4ghJd/W9fpB3+LF4yiFem
n5+Bp/pOcs6jN7r2P6jwVsrAoi9ippFaoHu8rzjOqjTirHF2y6SPTih9n8ub
vCyZee/Vb+VwzWOr1Lx3hXml454fjqWKa0T5Fba4pTes11Yw0aZJCMxUyquA
1Fq24rNeHNX/OTHsGTgTKaexhbNBEpbQfHFUoNBpjX30ruNLuevs793qWfpm
Lf3nJ6J8pVi/9Ak1b/iJXcvAnzd7xJvqKJDJ229KatPYXhCT0ve0lsMT2m0T
LO2mCQ9mA7rq0oNCvvQZmNOWKyVa0fB06N0e531XDRRcKw1BxwlS+rq+5t7W
2n3UBURlvUcijmKxua/wdhqhg5LBtgmFV3drL3qKZVvoADPUzfCJ/O013qV/
qf499PIDrBlWZm8P+uFqOO5osSXzz1yYqhj/GJmmb2qujojuHczXSiCHrYIT
XRn95P2m0/Xw6P7Ce2wPExk+7cfeel9z6Vsz+uVP1s42pv0PammYzt12wKJC
KYy5GISr2WGFgO4mjSENLpIMtruTrvPFIP/uJZ9/QQ+vOXNi+lCt4XgN51K0
MH2H7h+Akvh0Bsu9+lybCwPQSZNN6KGxcQiBguBvLIIidd26NFq6c5fPxoTJ
One9V7IyPRpXuPiCcDcuuQnGDlN1S/WYTFCEzwIpE4GrZT1U27a27A/+RbvW
01oehLBo40DxKCGQIrcSeWWtkCsBPFHaySRo0F4bwonfBKCqWNJEG0vWF0xC
QwNQ8oji8T7Bvj5SsW5E+y14IFtoVr6ScqBQ5BKxFX3LIYud38JI2JwTyz4B
cN//78GEcWTaow/3bE4VQoThDM+f7wl510dEeuUI26yMSgqLjzSETKqq5j69
YBdp5r9dS8zsnBR86/lWJsTp4oY1l6LxaJ8mte54wpRO9ZBAzTm2qSsypkut
z5QAhai7uQaO20u29n34G5RGGWgOJkOT6r7h2L2RRmqrtQUSUWeYWaQZulJs
xXEpYVNacmlapO6t13aDTFBz+nmti2IWZVXFt9gIACdyYs1ytSfRpnUM+2vM
8PZ+5GAwFF9yaseTX5TStVYDI55bpRd+GAlHtwqdjbNyuAoQQmRZ7SUbTWn/
q37vduEccjHiiyiZ9N8sB2RgAdInaGtiZwnwXUUE0nTk+YngGmmvNNYRLNUf
QTsa0944mXe6cEDTnDqSP5kW/kq8B1fn/zfEEIi7PwCL5WyFsS158jR1uWdS
ZJsjET+Qu3WCzod7ejmPUlM4rHFcpRjEJ4Ud4jbbN/GLXFYiOEw5/Nm9q2cB
I9qrxhhuZiuvKshg1IGwMs+iETkSN3t1JRzzEtqxBs38HzY0qZRutjaX9TNg
QGV8ef6ntY6diVYZE6TNuNohshI4Y2+N3shdT6vNBQBu0EqAc6NJ65gKcjkB
DZntVH79SJJHJVGcddKE69VrwWNP3Z7stXv4VkedK2wpxdi4taHoY925vaTH
lck+5lg8tL6UImGnSGSaCFF/pMxBM6WfJcChxld5clMDBsqWKtQV3HfMcN/M
EV8cV44jNmxSy7EMpdOCidRPSK1fftwy4voHiewf4uqFlUxTj4/u94qDzMDB
5lsEtnHQHf7BboZWPXTqjfybUWSE/Gxir9WhmOxYKgZEfMz8SdlTANGQ+Zx+
bxDGe1cJVZExKoRYgRlkMvbYRtyPlmT2wml4VqD7jTl+TP3G3GwKFDHMMSmh
d0vQK9MpJXMskkADglKIDwq4ie4ODDtNmSYNWxnEt+HrtsznJQXT9cakZ7FR
k1qbYRSHqZIxhIpRaHCEKEPqP/11pybvFQKyl+CCXphRjdvGfZPGUI5Fjr6K
czCcg7fg8EKBcFvdtrLL9gljUL2sQG/1pLESFW5Eyet5/1zGMMQvcUMCDW3d
7BSBqmK2Wq447/uExvzgnu0fDnbmtlXKI+5PosE2WYZ8ciajWNiQOQ3+ZmWw
N9lCG7I2nCdZtDBZGHX7I2fdDzUOAj9/Q4SHcPgXOKOzmzTOQ63vfVvCzCGp
QzMZ8fyDiYT/1zArtW1QvRSSWyuZzeTZY8bCsIJUYv6rPFXOzvVMtyZESjs2
YGdsIRkK0noAUV6n5mDyeWOekTXvNgURUQLZ9NW9rxlUq97QFPBTeNOZztV4
zVXoAU4ONBZQxMgHFCsFEHiTs2tvXu/qi/pEEvyHotGDPBb8GzzIGeN2L5Rc
I38rGqcL967d4e4tPnVtDdBezusBr9R3l6pIIaElQcsrKnoIIs5V3EWCA1jy
bIY2OA8BLeiseqUVEf0GF9/Yhnop8hJkSA3hXPSqXWzbLKXGq0SB9/8oYIx8
lX4KOXPGQIg3Co/vKpYgipji0AgYYXju0NxSncfTsNcZRQoUHct60Hkhecwz
yLMnq1wYUOWU9GWFIh1QOHQhTHdbQD6Y5/zyv1JgISLI6nyuc2uwU7840O0H
6SnrcKzWKHep1eaJBwqnf3vsAutIbGmqgnLFcUDp5SVp+buhhkRnSlqgMutI
0lnIZwlp1M49JUfkgUftIU12G6Xq3XEI06mJvgc6X3SrCO63Y4kCib79rtS2
0fBByVZGFVx6g82MRx+Vs6su9gb1yoqmvjZibYlCumOyxS2+KHurhDHhmtwV
RCOrYuuxGd+GLGVGC56ktQe+2aNSd6JjeGNHbCbOjdYhzvKAcPDylRYvASvF
fI9XuL01dzqIADhvkl9bgK6I4z6IGwsXRQx0cYjWCE5gZlC+evImDusKtoA5
LWXRTvOlXkDqC+KNtfKTnyJDqQT9QLSRAPoYxsvhsfvhpoYzSOOP6jS9ROQH
twPqKpl4bto7IUcc15idO//7vTFLbSbiXWZAzIMQDZUxYY1gP22rbBRA2Vjg
bjOu18YvpXBRc/I2wbwBZNkpFNWIlq+z/WCKqJ0AkjAD7CbcJahlx4kxq/qB
Ou95uWekjREFmk+FGwuOkOwzd0TJcTjsQFlQjgNW66U255Vf1KPcaSlH/fn0
FgSzc+1FPnhtMeANHfQbBZr6N0+8qoqqyGW+y7K/NqYGvNc3C/E/sJOuZHcj
4ggF7oecrAizmvSvGMS1sodsczVCBxvYAV+bQczlxqgGC3vNKIQNf1lz9zTT
2UbqoFewFQM2OW+E46vDkkWISejk/k585d5IAk9W5ruPlRItX1PSmTGiSCih
TuqXW7PrnNJbVpUQ3Eqw9NX59KlBzsItba8Py+u4b/1/FG64n99UdnrP3JUl
JiexLYvI8iZKbW97P+Di2wt2ocOWZDufmzgXStLi4x48cWitj8Qdp9lCfujz
66rAn/HZ5dKkcwdIAeZn4yqCQxZi70NYykdq4BBtbY6nekL61lCMcXrgTq/m
AOgMgMj8DcDsasGWAtjSOvzFracns8Rt3GaZJzbj52i5vYd/GTI15KixI9am
L887ZLPT75B8/e7I848QYRP7lqo2iLmg0y6XYC/hdm78YhwnhYimM7+80O8Z
Pj1VUhKGtd/h5nLXI5+qNdNUhoudW9nWnLqw9QOQdcC7gfvy4enF7KVB7CdF
S3+y9zw21xeH3N2CQGNLMN/SLh/FhdbHjjXI0ampTYOzsMvnP4wolhZZ8gWH
BNf53RXXxJnka8GU3ZPHWWNnMzPNkUxamtlLOnmAYkuqaNyWdhGoaZ50DZ1C
N2QjiquePTJaocp644qBoILx/gkBTQlIa/hzGJdw/6di5p1WT+XfwfmwaCyW
KjkVv+uhbEPdHVfwW22xpTIreXTc6HDlOuWIN2geziuv61axjE8yM7t9oOvl
iUvOuzrsiJAB4+zB7zIDbSrZ5GX4VxzoB9XW9q7fCKT6YFNzgdhbzW6RCP8r
pxhWChLbfimE9d19QmsFw09rTNKsKTCXE/RGCylGs5kcj4VpJ+D9Wz0x7vnr
BWqbdVWh3LoHD25SCUBAB21heJhDk/dLZrvCA0CgU1ggZ2B2eyQEMcim87CA
DFppXgtR1Q0ohArp8hNeGRWV+dAt2CRnugm9KkNzzlKfOukH1kuLx3blcilA
G4DGAmc1XVD3zyo79zdo3S5jnj7a7qySgpZQMmfnHD6MAn06WfVysszzdhwT
jMlrI37OJNdcDjOTNjrF3gQbIE+pBf51VvB78nDA8T5kJyzjctOZdDX01+YG
74HyORDAVRTKnpsycNWDF7n9j2KPDCgnHlPVxVUcDhCC42TyY28RSYIoRUXj
zW6O4fKgTZcuqS2We5s427LcTdHXl+iUo7TbR6MN9Beuds8e33di5i9XyPP1
64D1ZKVxxuANtZOgo2/2FHldqjNcw0aljkHgfG4NNhqpBe5tV9eXUzlwGntE
PKZKHCJpYsnJMwpKkn4Smk37Do00HoHezjUhZmthWfsS903AiKoefK+wYqxL
rUs7QOSCcf/kDrB0bD+QvduWFa874rk/O2cyFfdHf/M3pwi20i8TseHp+XWK
H04lHBM5gRp38aHVu7SD2ycRqwrraDIn14S3bkS3sOgK9XpkC8cHs4YkSthf
v+4W5pMjh90+Pgl3D2SRj2/jYuGJVAlio5v3dX8JYJjaeRCEoZ0UsAh4FprV
/imC3dzi2RTuNV55UoR44uXU8GEbaWDO4Vwfiwhhn/nDUOOTZrpM1aX+W0zk
j9DsK0y0KIzNVa2ryS3IRMUYkyLtDD9Xtojw5iRTBn9jL7YQDOAJAMKvTwom
Oj8ZqeUYEmvfcf/hShB8g8GEnIKpFkmh0NLQVAGqXlp6Yb0x5xqD4O4dpv+D
sPgtpgH9gOfhHqgrjSYVbTm0Q6BTIa7Xz7xy+Hb2YXe07D+U/DWt0AAC47LY
hLfl0wZ8qK745wZuY8ZwW2cx6iUdfkU9Yp5IiKTNxUrjfez0vIPXLKhbxhsl
1cmFo+ZYXuWvEzFtm+wV7PpeO1KXW6pyaJqjhd8xa7L9N0pq/FUlx/sl56rH
FW426KNBfo6XzXL5NV6JnG7eGXtUyL25ChwT8FZMBTSm6jFPl1WUV7V7rZ0O
rMh8LlMwbLrPcc75a7smFDpYta0bjeg744KlR6VYZLz/wnYacKCPucuB4IvW
GuuxoTfPeXmVSJ0FOFC823t73VLUIjs0VMRpghwgr5m9ytaN5rpgbuCafhG9
LKS0WWYycXzlVVWRl3pPVJ8ziOwurRwTSZMzVWcVU1+CRw4/fp2PAKS2ccQq
Q7vI7EB6OjHDGEAbUwl6Rv6d/GTfCZIGTAYdLgxJ9CykZOU+z6liIQDKGk9c
8m7zZOjjl0NF+9zQFzWMb+6KllsoFcLbFcgZEHbfzaUTODhDu950yx/EhjuE
JuzMKdjLwIXo0z6vQoFdf3j3oPXobdG1Ue8YtjucW8Ced6MSDTnZ/i5O7uBq
K1GNh9dJXyn6OxQb3pmvMHNgd0ea3lZWedj8W1lEE8nfyELVsJnyNkjtKS8L
IczDiWYDCKMh+nI8BfTTpyK6UkC4+jmonIHxGbS/IaLJKPutPa/f0ZJHdmGc
wof61VfFeV1+gM6If+tZc7igDQD4WtYWZIfCanPWmnnwlJncPFJBUT5wGQeS
ztldjnazPsixwpHeuCZP6Wt95ShZ41LRB6Zlb8Ag6tBd3PzzKMK0fleCpZhj
L983bUvnLWhcNSneEV9Q0IQNeY+6Sdg/LvvC0yP6PIJ7g2+08S5sfrPEKqjG
Fo57Xbfzt35smPZQe84W9zVDiUOmNoBbvEsvLioE8sNtNRBQ4K/jmeSnTBjS
nSSSDnAo7aMdzr5LSTW93wWYTtuwRJXU8+YHzeg8lCmT3ICNYoho/lUWh4R2
MN/aGy23Ei6l5N+7GLBjyhVycufGS5e4e5WcevLy+wsT3X9n4E2X8HEF9TCZ
Y0Tqmslrm8bMkWe9+vBZub6yEjMr8jL2X5dzPH4jSd8Pwn5RNKbjbV58cKJq
gQcC15iQnGrIRNa1d57p2fYkjSmyodyBXF3pa51mUqPYxSPdBsRJUg+2XoHM
Xm8HLr1B7PFavd2gADkwG/uu81YzNEvRBIEnLPRpJ2MQIlnkRNUf1NTJ4UG4
RALb6ZSSfRqlmfc103hCssLWAhzKx+Ii8ATtclea01pt6GfWPPPxy6wk9hZS
PuoaD5ZU1zC7v9ZpDzMWwP4Zc9xjanANbPS+x9mvT4AoEE+/aBx5Cv6G5rTY
CRPHhzeoQ8KEGT/mxfw711aZorfsJZNHBL/u+pGMKQeJgEeCw4fquXtYHVmU
KQsFNcBFbI6zHwM5V+0008B7i20159esUwt6a2xLVD10FpxBNdjtlEVOCkoC
R7GRmbhiv9WLAuHPpKkre5DiKf2VCmclqIO07iEPCmfj/pfMKpc9wUwz0bvT
V9Pcj//Tu13HlB78fVno61cnMhpzEQkVi7Ez+oUkV6sqi8INS9jfK6P04L7L
ERFg7LUlpophdvB64SUGN/NrGyOo78Mc2irs1lcOKYbazycut3F/OjR6MqkE
RWRY8ESxSUla8d2Qh84559R7bTiOky98B2nEAyO7LFK55iUsOA7PccAE0/+5
qMVqrbLSijBRfln9eS1IcTZYo373pLNJeVFJZ56HnVlm9iRTG8dMUni5GBbt
AcGR4OGC0EuGE9n/LpeTZZfVkjPdXZ6hvOv6FTajU/2NOw61JQjCvLShqLV+
DoCmjXvOMkZ//C5PuIio6kXNnSBbQLRXBHRh8JW0SBq+NJ4Zl3ZaUh9DgENc
plShtbVlwOBc7NddMcoMOFlIsPoFI59bOxW1tGVbx9pQwoifKoAGPKHtWqpi
oyVBsIIvHikvVZanc5thDFXCGxd+t8difkZfwCPCWHwIFJz83PIDW8IN7V/u
J8Y55IYI7YFmbNIckXMVs4gwMBc1Iiysj80jE6AGd62r1obeBObO3mSEfntt
oF/cbBLAS0OBDjBypG4VbY8xyfDm2Xt3O+pvFeY39OLQOhU9mqCrxyiG/o4B
Bfyg/bUhyZrrbvVxFazYRLs+JP/m8YQRtYMkHIlZxu7yCucFsSompTe8jdn1
rfin+EZ1xsc3WV/Fz4L4nj81KnjD4mufI7O8Huc6uR2VUIzAQX35FgdUsg1y
6PhILxpmRVQ3PkSoNywexzZBPHTKXZSCL2LcpgcM5qYk/vkKlWaKv2nxzvza
i+7zzCTOHAp/5h9dMg+6a+a7Eh9ZuCk1jRSd0EdTmHd5YhpyIBPnMQhM+7/1
7LOtT3cQshmCyFPQbO/4IOXcSJ8vVXm2Mmn2Nfj8bJZz/5lnNNDvJT3mX3MT
ZXGvk1SxO4NhPmslj88eC4fizKbwap5GZfeltaKyS911QccBYmHXWu5YZ5dX
zPDJy9JgsaFNIK/lgYC0M7MNDrwlM68fE9gHKKkuI4S4nYfcnoWW5+V/r2lw
zA8scQD1n2MqSrHdgOgBVh38XDFXDBFiL6iQydZdzxyS9hb7DGJj1rHl2WLf
QYE8Yxg7wDPXww45ivEqep5EfYn6kkzuqWkBVmi4x81QkToaP7KLaRhSIjDR
jfGsouvrN7mfCy6y+vW8j/vvl8AHtTbH6qlKGnrCGx6LwHpoOhRFILdjO6wO
GYlbANI2JAohdS6sY+z72a7B3V6pshofOn88BjBY36i4OQ99OhYt9+TBg/lg
RJQqLFSnvlPiGudZ74H6Wd5qpQZlpBQdA8j+H+rBdu6XfhmnCoRdVbEtsNwH
IgiZtT+lnS+3uNabTUgjFYemrzzkFr3jnHxrgdUpQf/RaLpBMum3h4dxaQuD
Z2AZhoa55InugcwEFZCQHpU5xnxh2I7u8gwDGpQZxhF+8MTeAAhTtwAkrztW
LG3C/CpP7G77xvIqDmnBmejumPGHidxOaw4wy5XCChy+TRoTt6QGTT9GpHne
K2z8rYPdr04frOQXH/thjOhvnngF3lJ+jOq7XZCN3IHtznKJNeAMdvB70ncY
fzVfjrC1mi6IlPh26rGUi+5yMM/PGFZszK0/1df4awvtzEd/aKoQeOR2U87n
gjGj3ktOpX/MZSbOymiCsVys4rHrulLCL5MdPLBPD/uxNDpBg2klED8m5BpF
Wl0SIvZAVvP0w/+oksQF7fQL6ngnrYQe6+8A8VRY6boU2z1EkT39NNogrDH5
OtU6Bn2nSShMTaDwGp5WvRux+yZjmyKcAarCcv4UclxxXGiw5p4mwoXqle8y
Y2IwGSDubtxoF/YxGrWQQC8hd52CShJ9Iq1f0OjbTCb4lqs5OZUQ0BX+KQRS
+LLfbWP05efOY6r2y9oMNtdej6XBKymlvi23kRXsqT4BzRCe7uF9AjWBW+Nw
7KyhOg4pits9QBPz9erUNvOTxweS5iuIDlpR6UljpI1SMVesV5m9GDWmEBhm
2wQGlAyZ20ybT4JdbKS3sCmePNeu3Ti0fsid1mamKjSU2b9xUDr2FQvHH+rh
JtTlvZklj6/UMAy2OGfYQNBNXd35l3bJzp4Oh7MBg1+FFkUVgrqgIEW9ncm0
cO+Jt2myPhomMjwh59FgUzBOV24xaOsV42G0LyERAJewXlzvHj95tUZNVGTM
8DSKBpqyMtUHXxbfoBTiRWTAcRTrkZ7mtRke25kiTeUKUbfAC57c/RTWbAoz
UZoGLt1AwUB6+SMs1DMyGnkpP/XSHMMBLlT7N8nsdOcgoUDVZenJeOWa+sWy
9Jk8HWJDls5KOKFbxxmrYhdYU6Tj1yP0KAvpULhPYHm9sUaaRuM+8L9fq0Hz
OW1XdKo55MOrb6rVan/stw7Z/4dUHAGSoAJStHu2Oh1y1eeIjNu3ODIAXbDh
GInUNCFTWIN7JC+m2F6+sAO/aD405OWDy/WJaZj136T69Wc0d/5t4lcs7SED
w3VeBvjCN3tjOWdow//FfyO4DzbQdc842IDOxQxqvzrfriEMZRVihxpMEGGC
D+ZxHNYCh4Q6bu1sbijIt87QCKoPw9f8W2ohNUoVpQ8BbNDMVGmsGAp6zO22
8Hpe0WldYxjf9uTa9SynGk6pXpIhYGdnerbTxTw63fbBCvGsCbxzs+VScU3S
TX7BYgn1SpESYTTia1mPNFM7TIeS0cC6u15zOvGo70AT3N06fTsJAh9a8Cjb
fwklnRcrgupzSf1Tqzd84jcom1sBDtivJcoY0AaWJlZKPacTV+jdTA0qrqzp
NIj/3vQEOjhbIrBwcvRCu1+p0ugvRJvuqy5s2DRpmIs2HK8SKrjDZfLDncd0
J/VCJapUl4f04EYt4PuUE+PFet1ETGyAOXhcHfX/2e/09V0E26qyx9TCGVXk
QiI9M9byLbC6t0m/4/ami5J8ckBxnsOsQ6VsZ3MbhQgErPPKmOOvbduIJV5x
RmGapTWFxtxj2DxsB9rJ8Y67DWBcBUHhzfZJKvlg54VpS5Ex1wfmNkIdpNSa
beTCtXfKZNN+kvLb3EhmpTQmP/1XBbwhsRRmADgRtVefUwfnZe5aFVyPSeuT
sK0Yymr/DVq/A8zDI2zsjOCAmNVMN/n2DrHTksVZvSMzwcMP9BjFzWYX80yW
kxSSAZtbrt3M+j3GDtScXZTDRb0KKhs9W9J9+rRKa6rhRCMw3uLoRrsM3zaZ
Wpb0EPS+xkD+9rNalzgNQuMjTShIjEHs7YZpJTgzk8zTDOnwZJiXthKztXzN
ppNEnGTgFIUzmSxKYS1fcVHMVO1AxbT7uFs/4dD3nOTMA4pVR5paR/LVzJ7w
uoFnfHsMEEA/9oqtCOAE89x3Op9o3Yh1pOUkRawAQ+9mJFrIQkEePpiHfHbM
aP190mzjLBmVhyWzmDV97w37XWImyuiy8t7mA/cHAMMko/C3tmfx8ASxPkiE
M0DiO3qM/qIc8wlfuNkkTcEG1NSrCdkFYS+U/hFIUN/zmYaHtc5mU+3Dx5kQ
6JsoK0SRZzTx47RUyuIWSkP2U66G/fOeyLNFIejR0gxjVJ4jFCAHSaE6esi5
3Dgb3VLILQAH9E4lks0oZJAq14NLibJLH+nfU7dyOKzkozdBRcOhbM6r2Xj/
U0k5soz7MJgt42jFc7KIu3GbQ4gTnDVQ7dHCAHrfxqpjR4zXhyoBNX1EvfeM
iBFBJoQZawrA+6uMcDbDpQk2H2806oLmz5vMLK9iVz8hoa0MNmVa0SxC7Tdb
vMnBJ2P9iRHboNGUFlsvnhy0cy+v8czaRIie1d8lM7F3nthsnCRfYjTrMvTu
WofIpEJLg126MBrq2VNNeHbaBNQ6am3CxdTHYegTOT1EFTrqZjVX6Ov/+jx7
m9SEDNtH99sfQGGesNqYqmYNW7yI9l0UC4mMYRIxvZAmGoMU+QaQKy6TrRPI
5BCKq12/s1h4SpK6rVt94HVa7hRq2+TV1OwxtIv/PoRRyyVAvx/nTUPoHh5Q
xO2YY++e5hTK3zCgWVRBp6JozE8uFDCMWCU/LWYLlNyGU7HPXZQi1bf5NcJQ
lvf36H79InfE/h0SbZvZvMggkNJcLM/ZrXkfUWiZri4+msUTjCw1ncO4LaRU
yLudhWutuO3fJdRJ9ksMvunbB6+AZ4Nr5N5LXvpBDf126x/ue7oioYrRPLGv
dYNVfO0ALac1cmwnLliAmk+QfS0kyxSn1n4v3GrJ4esiF+N59EojcOy76YXM
Ypgmgg8lpB/uTYkRFnV7iR+egdjjD23UuFokusmWTVSPTyFbmonXSvvtGkwT
fpRDDePv/O5AtHlg1YIKhsuPT2Dpg72zEGJqFamIRlOdETKdkOeMzV2T2sM1
DYdNpshoafSft8KNmhDNyva/xSwVdyPQjZGBA/TEoNOeydE3XA2v41YH3rPG
UuyXICNWPp4yImsZMFeshaAtilYFDWYMeXysbGoXOM5sthlo3SRNs59pULfQ
HBTb0kyp52+/zci+7dfwjhY05IS2UWdKbQ1/iLOqrMBc0+MB0vYsxUOiJJT9
e4KTd7Uw87urConWv6eOY72bAqZ7bEkNNfdN0dVVmhCOOli3mlxfTqnQpFyS
7UTicM/AT2qG2W8BunNsm4gmvm75ErRAlsu/hWZlImWbCX907t0KHhrO6mrC
a6SVvPmeUye6ckjvVYGCEn/vmNA1eeawq5WYZLwiUxGKlOuj7KUArRHgVAe2
UYUZzTTfbPMsRnniT/5ey00zWDv4yDJKqwKO/e0aAwQ5gjoyZhvU5MuwWLUg
4K9YGVpkRezjRPvc6XWMV1jnHguuJ9cBy9rHcy5+4+3kyBA/+znvpDMgh9Ro
3PhbsHpfWIV7bfptcwjaJZG1vin/hQl4vXZCJQ3CL/eE3C58tjiQNzd918wm
osA9TqBRrYJX13AtSYwwp90IaZPGFk9rrVTdn8g1ZxGj84Lb00cPdhhGWZ63
LktOwCJ1uOF9gK02zwvL30M9DTmDGA9JibJorVvKwkwQ2QrOdf3gVr8gyNum
qnft8soxir4BO0YbiJxe2ZzlqIMySBBe6QOdeUsi/gNu2Fy0Z42h8EaQywRT
d4ub1+HQ/AhdwT8Ad/96uVaYvIQPUFc1tXUEKducDgMGTZdpqv6l+dVv5W7Q
V1TO/nvCuJ5B1odkPot6Tty1CljPGFVisWS7jDsLZs3nf70cE0WeXg27M0TU
nkTTAKntDrBbMdrx1Kt7h15kz0mFRr9EXzKElYAGONvR56elDqkTO84hk5ne
1ruKgA3nc4Ct0XwxJ0U6CijyRfCgDHQWyskXmiCyokSpYpauKognGVocBtP2
cIqCsyC2aJMpsG87hgyWQJOoIRf1Ihmv3PDMoMDZH2BZ0/4vn1wyL0+L9mfy
k2putzeGa1/ZqmtKlV8Z5XcZsYTM95zcdDPEvo1FRTGyS9WI0Hscmo3f3I7B
uY+OmFxnAXhGcVibJfQEhBXBfqf5qWSPUQ7KwJUZAYMG3DylcXYhSf9AZhUU
ZAeqGN4D8BohgGk+B/MtKWauAeHwl82YGXoBhAswy7ZQyKt9a6QGwOtBj1VC
86kXb1vY4y/vR6FO+Vxn6SXzPjqchLhcwFnYSLBnvpQB6SMdOcSoxWSOUcMM
JRuKu9hC9uCl173FPoq4TgaAN7FPre/QJC4/HSb8+OphqnoSGQK+BV3VQGX9
o9W5z3ZMtw32RzlHeVlrTaspzcuE4OWqWte6LLES0L17QfLF50i0w8RDytSM
sfQscsQ3qiy7DCtpadQ8CVF3orfxtHgf+FTnI/kJcN3adDTzz8XflTb42UIR
d3CF4ptW860n0IErWidC9oKdp5Sc0T1GkmlKWkDI1A13eDWBTqHdsSHW5r8Q
TEqD+JJPFMn2Xnvbt20LCUdqpL55Dg/OaJHctcHTLbOcAt2virseZ0sMYqfs
WTzD9x/XBfFkQWNmVfI29wYbPrd6YUYqTAOupqjF4dE5MohyfNTn3eyKJkvq
bbkRYMgucJuxrW39rYI2g/AMG802ucfH3Ci2XfmGvd1J23aoytv351rGQEEy
JnIvqW/+h9IlJfoYGk+7Kq2XkSRcUACon9ct4P3BNonPdk6ZWo0HusW/srmh
ezFljzbFkyRipV3fnESm4Jtga+ERBTfR6GT8uwIntDogkWtvvBW8WC1EmSAZ
06HFzIIoDheb/16XW56VT1J29zyipzicGX81ODjR3pKeoxAj34N6N6lUWJ8x
p5E+xXGtzf+YlqKiYJRPGw5JYbF31LtMAYw+DGMc7zLelttdJ8s/3Ye50tEf
tiSLu5ZeMHdWDoDAM0uRCjiO+AlLr+nsTblmnZTDNTezZpOPb0xp5CJoKSe4
eaAKfc95xQ/moZj7/RuE4Nq/LAITTi4Dh+RgpWP5Y4taGjcYG8OtjL5QUWlM
fHRDykIQ/deK+pOE4ZCf9UUmW61SSPH+lOiEfEQezXCPpR6Je9u0kGRb5vR6
PqxblCZH5pE7QcPL6eLmDy2DnK1eTefEfP4XokMQGKh+JRlysLDrWSYCYlHH
IBeThFOtENousQ69QK0Lizt8p6CkmLASiiM3i7roGe6G82IgrfKGaz/k8Q4G
CsvtzXr6Md1Nn+8Lu5bo1loBECATgIN2HqOPtBll3A71A0QDsFxxKFoJyOHQ
5vtxiO24sLtOtj1nz3GUYgRF6N2fdq44uP77P75ZytfsPwWJFUiPUWiI+0Ny
Zi0LXw85cqinLBPU4cfk3DZHwtfH/Yb3vudvPNTfyYsdfgy4MyvfMm7ChcEQ
Kx/g3q30abY4VIsHo+W/RzYK+dLljBa+PWjpUH/jK/s8+hSVmmsJX4CJB9Jx
5L0iwymDaIPB5Bj3/xO+JPB+jaVurIdUIVZTTj1e1kpgKrE/tjAVnn1ymiIO
lrwe1//8F6wTugAsBKqYrDVvVEv0De7khv/eo65RvRV8tXzBKzJWKjD8UZ43
EALrHhejXwQB36486GJllmbxtsR1WAlhsnYL/LOzk6cygTlguvfxkW3376+3
2GIrfyVRM/U0lFy++boLtZvjWWZ8/AElqThyq6Ef1qnif2JwI0ce5NtTsQBt
n+g+zbIAhGJxWayyhUQ/Nz7nYLSFwVe056ynT9YxpVe5BbpBfVDHF5YPq6/7
EU+iKzTM4DJKfjeo01knsNRNCBI/R7Fjnvj7FwozbKMYIK3PdmMGi+EAT1lz
5s9LruXSKNx9JgCeq6Et06v+m76uLp8CYjLnVZJ2EM1DI7jYYJ74kNSkAwZ4
phVaM4Km+FHQHGFzOsB33VqGrFkgInbJ6ifIj11EQI0hxVUAwMl/kkRswyVj
F1WvJZWbERtbBQUXBsChZT330+3Z9KS1PwNuIcXxFFyAFYLn4PKL0+TNWpa2
R6A0n8VoS07RmL8X6h/Y0qIGd0l+lyMy+d93rFTnlct84iY6n95oOMy8mlB7
qoSiPZPNSRTWtWCZOSxV4zXXQCHVR+8eQuue92uDhsO5Vs9kF3axtXfD7e59
pu8NQcW+R4XmGSVWoT+KUJNnOeV7kAHkMiqosKRYrpVqRmWmUW9Jbjb548Pd
4KOpkqpnFFu/lKiTXqE+rsA1l+lVsAuSGE6H3xFFIKhS+/X4fvDz57q/U34F
FHDcaXK56oE/5WN1eivmYo8NOZLDT2Dhewk/MFwk7tKmb4iiaq2nvm5ellQn
uPdozWj15o5hgIbjTKXqhFyeypJiSZf+53LvDDiLBkOqegihDGikCuNFzLUq
EqxmH6DzaUMpMHag01KygJYz/w7qcUXZQ2T+POc1AucIWhubTERcQSZkwt/u
8R0XlEaMGrUH08NJ3c/pXF352XYzPlDM0Q4I3AvW2OIvb3v8aU/tTJdovHcI
HMo5A2RthymrQDi4PlYK2DDKIZg9eXwoSTvza+M1F8Wqsqbqz0lMmEki0myy
MnbYxFbOdyp/oMUA6esux7OqlspdANxhOMZIWQd7CvEGurjwa3kDULmpKU+z
SW2zWhkLtFjmCu8ndfLIcJAb0tKDkOGQd2V2uKFjWD/AkpVS3mKkzhFZPrQq
AWjMJm8kQgQtKxd2BOJn0YRZvgnB/ZM8dBVnBrCJ1ogCArMaU9YygfjZZqRt
tXte079US4K8BkLL6t9U0puZ5yXlXQ+s+8vdqeRM+v4hXgE/HN0RO2XMlISP
IdvINPZ6OK4jfw1S/wJqJ244sLwltz1MOu5CZl8fQLJBd+bXvuYHBjsiCgDH
u1f2lo6GfvOObyGppyg2rtOVa3p4Ea2gfTJnyCQ/d/sBKRBslg/N+ARs1sX5
elvCwMEzyE99F8rt/+5GTXdYxeGxbxLb7P0M05atFRmZB4czBBsI+ft0AzB/
8m3ebgwuvXWn8bkqKE8M3wPpx74SbcXh2Ko5htUyXNREqdsj8/IIg6EcjudQ
zDj29jqymMIgAU0/iFrS/mkNMWApMoWZR5v11OZ02cuX822WxMKga6MoCCvr
UlvXWw0mkxPSunZARytu8pbCfRejLU1znFKVgxC1y2wh4mnR9DGk+fjLHyqA
SkCHuFaRK4oovPGMJa/GxWxSKyo5W3iF6SM5pnWpk9qMZdj8A7QlFxZ7xm9V
SCKRLDJLKXkqXzmNUZ+AJdaBZkvQgachoMH3KlvwUMm9QLMWqNohEIRu0gRF
ckHxpW7F4wHQCdx/86/SwU3YIMJDD7pqtxHFsarM0yqR6fDfLnGWaqmVSOmO
VeuVRsV7203RvEesIS51e1/0Pv6Q2jMVDX3bTjAr7QMJb+JzFDo2ws2ztgFP
/jOIhpNjgIlG8rBnQA/H4Sl0ezDJNSMREgcJn/hLW1qPv6rhNoIKfTUzgFqd
z6hNJ2DDk9ptzpRqMxPbKLz8nJhqZ1w2UN63AviAqNVMh/nf9hOMiLi5UAdW
ZvSiNhAmIXY+fs/Wy0nJt2FNcSJe3zLKwMeI3DNZnBHnc9nhwgdH6847mHYB
n9vsHsZP+rTOtKOIBZ/WDJ65Jt1lOsSgTTlZfgWIZaZhkPXAfzSp9uNfrVe+
x8S+tmBV5PpakZd7/Ngx283lHhnWsw0O8bJA6qz6kP/WCx6kau2Y7Qc+KIij
qzO12AvSBKhlUSWBtQpMvEpMf2YyocA8bdcP5V9bHdTeI1uGj/P0meyN4Zn2
Rz20m+TTds43duzLP6Y9E1brMHIosscGjTHzFqG7F70m4vQ/cq0nuEIM+U+Q
EZSf00Tx9w2In8JGbrjWIJq77i9XpotjS7Qo6ZMcO8tMaxsCGVCuDRpR6Y6z
8AXPI2kGvf6iJgayXsBR6SiBHgXUsmyXlsmd8sKWYNWBZTXgU2d0rTJLJefS
p3kT9s+JQ1OSyV8+zbeng/pxf0yk86ekpSDVYfS+pGRGznap8wDB1jkLh0X1
z3UxrF2B+xiaK3B9zXhTvBuBW5HZ9cInuQTp2vW+nNo8TgJXkc4/fegqvTme
4WTKZjp9WvfUHmGHS/rsByjFjX7EbbJEjErraUcj8XTU7ja0zI890LNcsLD0
HJpJvjDzHgLhcx4voRox5K9pZEi5hFOBCgjXmRMQUW2VUzlAOakmpBEcOcjm
7FRNNufGhq7+s9yBC9e3Vsn8vHO4ymkuW9B9CbzcCTb6AIRn6duC0+de9b9z
cygb7qX/Pn2W4vwViZPRDP8QOsJb9IfbmZCmkQOEO9CSEZQeXRLuV3t5puc8
qYOrK6qAWaxd0cv/M3Vxz22daGIyLr+bxApREeNHqnWig3jfhdq9aEe+ypIe
bODcqBaVCcs2WOqZMYa1Fo6d5Xh8LwjbBlqZ1qiygJ+8QBLkscW5QKAmL5a3
wMiwyx5AI+VZu9YsD9E8UI5goWr3ZKRBudrXdS45r15xtSZn+CVQovCzuKGt
k1UPlugtPuyPhabUvJwhWpRcza35zCODlejRMW4JVY56V3l2LgVK4u16RZM2
+h0wVRROH4qJzsfuJG8P1SZk5s9IaxqJlVVwQuJ5FM9oVIg0h66yROeBmI3t
2mNWGUoZxFtyAfWVM7RiS1yO4NpDjFgIRnSckCb82SHMS/puLXXIEkJ7qsjZ
fgw//5nd2xJu3h0ueag5CEjah9nOGyTbnfx/ztsH7R08N/2NrL+j1+XTuN22
E/yFGCM2u4loJij3HtqPq2KmR37tVfeK1FfWLxmPlR3NHPi1PCesF138rDJH
4VD6+QHSJFcDk8BZOirWfrwyVitutN8/WSsEZK9NEpsQyBjBrDfAVxW6BTRb
98I0imA4z9e5Ia/2xzW20ip3NjufY4m27zEFC5i08LL2ksUecdvoVtKyjgkL
++U/Yl7FTRxGsiUl2xUeyUB4h33jo7JZfzlCd+caxZWTV8KvLO8E6Y8ZBzBR
yz2MPoQ+oP/R+38ZkIgzvyYtKg6UngSW/Ni+nasfKFO1L50rnlkcc1kwNlrl
mELyXyydOVWywUWneHsXsq7i6WXQr6gZhwuqkSUapaSEEDpfMxyoKtEkrdyq
RvH4gzDdm1ozv/HQN+3sLLVqnNVMu4YP2lFCOhHofML/E3lLqv/y02eWTqvu
e0U0x1a/hox9SET3IRQXvk+y/TZ+uaKcxz+sObPFIAnOJZDc/G0zdqI/hM7u
bmcKabxXFgiRfecdY1R9Qn7CgC7ihQclx2MO5TnBWnXjUKOPXecqADe+3xRB
AUZu272CVXOPcMhJlJ8EyCzUVz+KUANfgHFO9Rha20maGQZJACGDamdGULph
1hC+KzxajVHAcwr1sT7aDH+YOjmLeaemS2IzykU1ZRQRGBiRkvTO+22b5eXw
oAtzTVlOK8FHAuLwT4GwdbubJLN6ohvbFBJqttgKysAFbdh7Qr6MeJI7imGx
J+HuU8VgPAOVuvWE9rxzcgQ/6P0pZ+Tw7fhsEeHskGBnX1kkSxIBtZk1IHMi
Q8JAg6ywpK02ix1+xhMWnB+upg4adiFsNpGMnb9VMg9Cl+yPbKaO5pUpXVsT
FzQoCkEqynphUwzUcAf6UO4xLwcTx0Z7LZGTyR4Gtp0l/nl2kSl9O7alu60z
KvNgU4aLOzB4urGl6EkkZU1T5vsYaAFG+2S4Bk2XiaMniNX5Kme12KYVpbEs
Xxkvun8kn8gJIcSTQNjmvRhFwvLO9dE5BV9JpF0/Sl8sur+x6nxmcEe4wVTr
0Girrjv4G9ioLMTcT+1Q9qqbxNGgaS3fZ/3utoC042BWsLKLcj+G5anzu0na
rNRu724wXqVjtxVVYTWXYXmhYcUYnHxJQwLb8eHqQjO8vIFNnxUCf25LNnRA
8cYhYeBihNsNQIZDjZzn2NdC7HAOIUQfbK31oF+mv8QjmcX5a1fFkfjNZJc3
vTV52rdsyANPhvIdYxRrfDEGYYS3mTW/tUrOw9DxGRWZGpljsBA2jJFtxq0h
VSabMmHpkdAKDGeFO0LFhEkBBjX5LmG6t6M7q0oMRNmLGx8MjUwfB/G9wuej
xo2R1GWbCfUta9kJ+VSKRIRz5k1S4xwCtlhsIX+/Rqn0mxPVNKQDH7B/ExdI
oARqO2ZJAfHqkUHRCV24YUnds0NP2Bn0K6CJd22rxux3DoJId1war6OMA8oq
QKXzs23jon84YRL/kg2BS+krNhz2R5myBwZ9tOwm1MdzxVbA6TQmAWjDVP5E
Yoa6iv8zbuRJLIrosDxGV7kn+jFCfnJc5bM88mid7AY41LpXa7cuWOfyMQTZ
18qh37fzwBhsnIO54tr5g2VpQcZnWh+2fyyBU3Tq7b4mjeU1grdOan1F9WY+
sztWmXgujjL2TxW3UwxKk6jC6Ab4rCJzd3btzI3W8DE+I+bxg8PIVtRJSpGS
xwdLDhNe0nbZjAj21Sd8uVi3sxIVE3zR3TkvOxloE/kQXCWdxdajxftxxoR9
MLcA+GK9lWpZiXaWyFcDf5dUfrxwbEHoN2zBc9AFiSt5dDMyuQ1/2xkVrj+1
EE+AMh+7+DiwrcqhXYoVUILaY84Y3YXAynR4fKMWwYA9hJPlQS/PtmIm3Tco
rXs1Oegp1T8RBHeM7kD0lojMhRZ2MkPcCEas6XUSSVzsxFIeHSAh/M2TPN2F
WOo/T10Hufwk5cT5fis2u+iYHXfeoBuXKSbE7sF7RbRi8/+npNwX2/ztiXTL
GwmMsrpZJB0wqmlx9mDUdB04XX/Bhx0j1/ZePqiPapwC/wTImszrgRQcLtu1
WjeL7rDVs+8jKR4GWAs4y/K2h00StAYgTed98eJio+ol1YvwTIbw9SfjkBgz
j0sMckdLg5S/hV5+7DC8NlbUIypUQIae7w3xOjY5v71G5mucqi4CmCcob7OE
FofrslSul5AqSaiTOqT/aXmPBQvbzHoUkd7uZvt37wi2X4briIYPtr9xutQp
Nuhqr3ebDQrAPzWR3mwLxNnfMHR2JiAgL06IMc2rPn9677B2pg+ZZSnatUor
37ZCEBcq+UybkdqwTdYxZWadzRdA3FZ5N3biRB4QYGFUY+RCNtYMna4x8u6R
DfA3k2P+fCeCsHYwQak39mkOhzFsfxo/exoxo9cqE4eXxQKJ7bkZfuNfO+w+
41Aql6aX90HZ9j5Mtq8Wvx3rEZH4lO2uJujZYds0My1ZvMwCnPrri9aX2McF
X+3SUqO7SzYfwLPcV+cvrvJwJpxaMKpXuRVv06GpSCEB79ougIikxrNJikBA
/eGwdmORwbJm6Y3nycMH8WMuK4h5LxCxYVRAj9fL/Ye4Hiql0irGvE9mts27
0am+tWHv5Jl5rDA8t8eiUeQE/IS3MTla2kTVA08H+zKgNV6GMfWfON6zeLTd
7H23CJsJFWdTMRpOL1EracLmF0nQ+PbdygJJJJBpunyFqWp3IadxAPV+jSjq
MIh2N2P4NaSEr9YXFnT9tV0P44F4v60qeI9yNNG11L+LZngFTQ6LrvMZGV9C
2kBU4WMrZy3akE6ib+P3D+K9gykzxN3fn+ht8HVtm46e1VeDGyYnFoATT41z
svM+WzmTcMVBprn0LBbYJDmZU6/5kxdPeVeBzjVeqTEQ5SyZ6CBJ+NAUO9wS
1JHchS9tkxEizWK8nkhsbTmTWS/GECtto41FCB4gHMAqWxsltUMwInAc3QX0
mA3efzqypcIkPLgbgOjH61JdDeEoA5SI/kCLEl8vlV/l+dQfzorE++J79EfQ
r67Ltn19ADsJs9ah1hTTtAdImnfOTCH/VNuBHRbJqC8uU4lTt8fU14EFF3lS
9yrH4NdkeXIcvE6EppmTShV/G/nvS0aYgzWdJVcVbbKy5F1O9+4E56Kquncb
DHFO3JUdpIXM2SZxZ8xhi8Sz7XG1Hn+2+ykn6ywj1Pa8bAHwfVAlcutYp3uS
ccp+OUiWp+iGcfzZcftiUnHFj7QuLoRla93Z/efkUtiJ8InD12xR4OQNowe7
Hw6XrQxNhNcrcLDGII/rtbPpBWtcRVVs+KYEyf4P6Uhz7mwGfE2dAPp+TG1R
layqyK1BpKqi/gg78wdDLPre1k3G8QU+XcHIwoG25tDNJSp0j0vUnb6ulJp1
QyeNgGhOfeMJyv5CUX1ne+Zu00FK+YZTvyCojLpSw1C6US46aZim35fYUbRw
RbjYgjgvNfnBVF1AEMb9wVOmZjX+aqVYV9qUydpuwxJKoamwb/mbYrTRcviJ
3JXLGQOQ7cy/x2/HjpQTYk9+qOI6vy/Ii4Zc8kv1O//ydQ5VgcqS7bmOpZ7c
K7WtDhMDbLfcgNBvrlARQn2wJOT/qtORRxj8CaH3tOljbnTRHhMfAqBVeT9V
qXfI+irU/Ub5Hmm/NFDuhhYB7QGcNiu/Q6T6lYL6N8nEjz2Ucoby6KeQSz95
MJNRebnqm8qWolNWzVvtX1ODv2s9IKnGZ55lWvDpPffeDP3gyf5claGBX/tZ
4JD4uIhjZZBv2Ct+K77pC5wLfTtafW6LuYQrk7JWzb8prempSTtYLw5rdx7E
52VdnC0HiuxRv+0Ab0OrW/BnL14apWdUFnA/pRG2YWS9xG/MnB8m6kTaUlOX
b1KEj5vimxFdV7VDUTybVBC6JHXcPTGvmeKWICk9P4/E2BMebvtmH4IiPsnx
jN+4FZbZWEnviylHsZpVWwHcP/54SA+A4nUl6GG/d3Hez0kI8fLKYeg0WNqh
kSNz1mVgFmnpA6LrxytTo7Nc+gCTXqTOsiBwN3iyZIyWhLYpER+cCAOltIty
zM5nUJygRzJ6VzH9uyHwc1H6XtbAjWu9YeFyMcHL8PXyAijoXvxNHWg84BiY
Y+OhV9TSyJH+r9kSOxUwfGVvTQkVD0sBFaKXCZ4FaXifxIIJLuM6rZW3viZT
HE9daGnVz9jy9ZBo8qNrZI+Vm/7Q8BEfcruS+311llimlC1HRaUkEmuUcXQh
XUxLDrvryfr/oTiJKuwbR1YHUFwPNk4nOJOKoX7eyikzcveMQzZSjHfW5XEh
b3rHkKYsZ8ZZUKZ/GvvpNonBMj9dpWwVNrJf2/CVHbSaWwuCvGKfWCrsC0ht
0t8X4S6ndl4/W33Ovuvj1+FAjKhYaiIpkGjURL+U4sPazidqk/6kXby/nD0M
l+5elw2Qf6v5X5hu6sBwUvg0JWf44ge73gWNrW0p6CGXxd2a5VK66bm+/Gg5
Sjv3fgXXmCPaW4oxV/1ucBC9+b7efko85WnM/d2DPTw42xFwLDBBK0ROtVU4
CtL7muxq9bFKSVyDUnnKbVRGuxb5CbP/o5iLBVjYMsv7SE4srNx7WFZ6KN0h
kW1ca26eXUQjOTIuCioo2jZsPpQWciJzw9DllbHSX0lsWyC9DpDe4nvIv2lx
p/Jxuyz4Ppwq8dlXpKandEHeJHZsTXPHEwiWJBilVYKWD+MJJAU5myyfBhV4
CcVyKdoSPlz+kg0ZkjHncUd5RKMktdi7q8JABNk/D6A9UbSNV2YT44A8CyCR
pk4/NBS+G7Ug676zbSgVRWPYARTqLERmhOoL0H8ZoUpDZCmUluxJJQhinm1/
oJcp912ZnbYgCt8hrl0CHw2x+iucX/z27YVtxzdKMlWIVUffQTypqUkgqmPL
eDzOEJHawWMROTys10diRHHGfiOnmzF8PNOIF6SCKHqQ14ZsfYpm5a90QUYK
96P9qT9cgB9ba0wBwlUgngjpAFqW2SbiJ6o0o+fofucbtI8A3YMNb7ot4HVW
GXysJp4ahOb/CAwTQUNu7ATA45BhBEmsf2f5//MXZAGOI3ZSaIFJDNlp5pVB
QojPjKwLz0ZdAdSoAeqNmqzYT0BdIVIZ+HiPtWAm/M75n971zw2Xcv/Aios4
3Rqgg82DDnGlhf312BYxN/pteSbCPEr93j39VObcMHMP0JA0SgbI0WkgNnI+
Du7De0hrkYhPEGzh46h+KnuuLirzFEgOzAo4WUSsUEReTmDxHHq9yQoHlpE1
ymVwabP5DuODS3w5LDXmhFw4CxWj4Y+QTTNDjXHwdkXMnOJTAKr+zgAYnY27
urIG3HkxdZFmFamoXfJUzDt3bg6yj0DjhsvidN1T/ZlWF931Pdw7rxzDomph
42X9eQUfqBOEqnJrQsVTSQ86DYafu9PtnKuBQWzGHnUpt5+2rl+6pHDMAamj
DcUh0WeyH67Y9UbXXhVYtg0rLtdMkLsE0Ke56+BxLvPg34JjZu6qI/BXDTwp
CiAkGBz03WzxaASMzoP4/GctG3bJigYxwQPyURpnADP463bN0EkY2rqpvZ4p
wdvQdQfqQnHiw2/v47me6uZx+ItLet2+GgyAkQ/s2x9xLOy0uBF0P3qaPZid
66FRXjhGpFPods1qEm19CooIfFDS1l7pE9dPUGm62nlBKwPfbqMoXfL0wEJ7
hvkTPkrf9jfm3fVJSVs4YN15cfR7B6zCRspB6hzydkEDCtGT4r4pIaG6CI36
NgW5rK4Jeefx+ev9ulMFdWLdsA6JRgSbv+uGCDyyQKdQ1K3uJtOeqwX5YVDb
PgRyVEwZLfW+FVnMwLUdNHT/WX0tJqQ4z4xqLG6l8891lQzI43sFpb9eVpus
QyaP2U8ffl7A5JrzlaxR4TcRV/dPjecooxwYZV81h7OdPteL2d7EdDUG7Y8V
Tk/1lzCthD23BrUH+NuyzvdFTil3eVqbgGt3fy9Vly/LKglnOcd/srhRHNKo
6IH6xDpvwexArvN1zmwwWq2SYw/Sp5MKLJ7RJLOdDMjNY/oEjZPAjnWdbkS7
pTSN75mBDKL2e78XNO1reIFt+GaCfQbcGUBXXj9wUpnr8ayCLAuZW9eh3nIi
31UekqmcJwj4QUoIq7suoOnl65y0Zeykkfjr3Lkh/8HJd2HCt1vVEsemQ/0h
Igu/Yd97OP2dliI0HUKhIQuArkt2Gl0BeExLWKRhr7Sd4tEuJFubz3jU862h
4qicxWQX02g9JV454CZDoozTKlI3EVl6ofeWZQm4dBAvlvt2gUEmTrHDCO6o
4uqdX+RmH/zvL8FpDILPWWeGLNXI3Q0OXM1vTX5fiJ+HDYTidoHSH0pezn61
0xgUfjjzTST89vToMIiuOdzXa1iIXXYNWFqvOB3PB3fmK/EkVt4SVotkwNbE
HkidBPE8JJtMhT/ouINz0m/wPQeV7/JgH52JfjGfkQks5B2v9U65gHr6G1TT
d2jN0Yl0rVLzS1uAaLkDCVpS984B4NAZhoLCztvgGrK5UPbWLATjszEN0W6b
gnE5M4PUE15C3U5ufI8CJy9mKp/5MrqqpGBAxVjwz3QyyVis76nBVoXdpgh1
e8sEneJhnMp9ON/jKBEjpq0/BIRK0MRoyD43mPXgibBuiBgbzeEyVIcwbGLk
QEwKV9z4PGbWe/6J17MN8v/0PXYSkgFMbJIBqdrKjd7oo46jWEIlXIp6Tlx4
TJK74A1OFWp1XjmON3Hypmv22kq1m6JeB7FPwwJLxOo5wbbUqkMlR25oMsw8
kkRk58ceJB9sxmNOyCN9Gb4Y4I173S/65EWz8tiqFpdQt/7LyG6GCcCuUAfP
/7ioNuPQLIx5fteT4j63EtBDiVm7o7+VnIHT2+pwW5wY4HmYQyYcVC0JjJWn
TowyLVKHB6wtWLVbl0IEwkcDAobC0w785kXgoro4UVQ58CONXS38lPIS+0Qh
hWSwFibvXmGhHvJ/jOMO3oP/pmjuh5FKG6C19TjqYzdQjkq89gQW3cMCJ/6M
gcZzFOIB068VGho7p+acgQftK4fuvVPShflZ4M2+Kqbr5kQRfn1WpTScBdiN
/QECS3Kgu8gWkHjLlElY/igwM+p7w30VQECAspXIuNHzRfPXS2yVTFcgRNHp
eJV7gXd34ZZL4vECnomCquy+iGiWRD4pJoXoSUCPefajNqIrB4jXDUOGBfpJ
oBJ+igCbxNjsL8Xg6G150HBC2Ew8MW/XljW+24pxTis7nMJ+hSih1c5trs1z
sNHlGJcD3ujM5wcNf6cc5JnZY11B0sG0fGsGOaK4y9Cfb+ExOF5jTOSpsDCL
iLymViEOfJreavUvS4+zRpx+SSZWMllon+TtfOTnjYMFWpSm+ZFOPM47fSIl
EeoqMH+VgFhWG05uWNWvYOwejWZjcVxR4pyvkFjFza5tRpTY8DSuqlftpldI
UuTOSo6TwN3vtyZEUzUZx9CS0jQzPOCq6IriqeSBVf7vHmfGhBu+ta669vdT
tfEfy+y1HmGWmOATTDHXhlJqAJSKjnlFYVqOj3pn6aiNnylRYRIlhvRzv0m1
HwAy+nPoyDOHCuSqEtWd9Yrb+VVfFfvVQfAOrgc0zkSzwP1lTo2Y5KDbVrRH
xXBhpZtM5JOOnzNfDyZC9JC5K0tH5lECYKAGgnPxIzfnsQyhUDq3sJSeWgHL
RX5G4JZF8tBUPmuSEMmdm3zx/zd+8PqR8CzTeKfumUtu/2QZCBNsDfPohbgO
vLZndzp/MpJ1s9uC7fW6+6lnPxHis+dx/s67ZMZM+qqPWbbsUXcycDeU239B
S9kCoiAJ40LYhXEnNhnJiQ4vnGTTioMsxlQaM+cd+YIaghT97CIkBAOe++0L
gi7WoX1BGpKZavtDIFZiEFYRMFN1lV8wq6QU1ejYZs3yMpNFxdWpmiZQvsHb
lAyIo+7867Kr4SkzE5hfRfD9nFFCbShEdf3c7WHB+aBV83ZwnyEzvDDYuLZo
/9PdTeleKH4ZPAcbyNVh7J5f/Hegt7i2saLHGKhOL0dMH1SVGlxdM6Qee68t
cV//EFOr3+eTKhVlZVKrozFxRiSoUrSERXFu/VfBdtv4c4J513NPL/TGITfK
O+eiN/B/hXMKXgOtlKbJsW+bhJFlC7nEn+5pN3SgKKRGPU5E6WDoF/kniTzz
wBfcVhKSsgbgzDEMhxXF6jECnhztXpG2XPxbg70h6WBgRUxLylnJMEMs9Ob2
MYb40z7FDU6Evh9eSF1Rp96nJHd+bdo8mPEe2F2Twpi1/tuDbZimELncdWt3
xYY9P2XpCrwNOTaufOcWIWkT8NP/6Zmbaj8GdqBCcVMfa5DSCYRmfkx+64pa
3OMRaJxBiv4VSnQL0PB+8xzllRMwVK03ySSn+2GP7cByR9p6l3kJJ6Ljdfqu
InHC/d75+koUB9XPk2Fq8x0ecORu/sKyAWSHQ0Vi26jWl3egtujjis4msnvq
LIFiUWfKc3tfqTSdb/WWlgvGqb3YLh3lA8lmPS6RQAnKW/B+XM4EjlHTL5L2
QnOZKqADF09j/cta0dS6qyKcmOqhn/bQDSh7QZuTnm7DlYGE4u9ZL7Z7mbOb
klUtF3e+ah/OM3OkafcKvglgAc9VLSob/mphCDzwI6d97gnuwoEG30dJNP1t
tQ8VY//tIh+DE6bnQHf/ylewSN42+eBIBnCFvdllQBbTJjjEm0hnKqOsaI2n
7znZsHAJv2ti2Db60mtPA367WpGqSjaqs7qDW7M5lzyp9wgC63Jczt7aP1Y8
c9jcz/Kp/8XfUCoppiP4IZapXRZ0wCa7PW68pOzqni5vR3t0AVUVAlhlF8EX
5uaoWAGCey3QxNOGLS2Zbeb+VWPW6MdSMQg82CU2+rX/SIyO2Pkz11TMUcAn
SBBYDANcK2rssPfYAXdPxxYToBPzxPjs3aXYXZaBDM6jIGS9UCXXEL88VF6h
8EOH0C6EGLbQQ0B09j2Cr0qzCTzz5HF1x81M+AtT3Pe6yA65fkYpB+Fz4DFW
LgTk8OL6OJYipLQJlWDzusPRsk7jxEd02zhnSSbmLQ9WxP4a8xAKuSLK+8N4
teTq6u/ZNpHTlCiNo3uq84238U1EandknRbdLRa1Klu846lRXg4XXdXcGLUx
jylCU6kxUWfGbfCDV6dg9KMzvUXiRnDRt7AYaU7pVuwSYZp7ggzhXbVLkA3L
C7xBcLVZfF1KK6alO5b9orXYHsN83Ag+yoctIBYJnwo4DQWoWjsm7SsrDp+a
z597LevLivqdl+N/2nh6Xt+NB0cWw6/eNV2weEpME5cum2e0CcteFA9Yad9J
/Fmv2w6F6MdQdryUfsh3l0C89PufcpQCa/MS5IBuIci/ujGKrxkdwDQYWx6D
SvhMOMqduEZSneigDOpwvwtnwRAk6GUCNSLG8B6ZxOgVx8FyAzKwV7jbLsRH
2/40rTkZHt/42kPaC3XtRZnax+gOfKhKC9WfqxZJw/2aEQqgHyc9WE4TGLQc
t4bHpl3mtgDQns5RYjzfzzzPXgEsJcMkc/DvC5ygzPzBgLwmujGtfx0kKV8X
B9ImxUoeZNU4/1woPzHILrm/LqDe4pE47pusutBEEONKLEGU2juSRjQ3Ij0u
+S1x6JTLFrVBeeg2L1aMpamPaM1hQ0lMS1mAOaTDQQf/C2/fu+eP2n15sHzr
EQ919CEmbceJVTQqneIvNuqzAmiZIcllnxuoZeZXznHjEl3EFpHs3Nck8bZv
ACEsU6mMsUTniT1xgTjObVH7hBUVQdap6RTrBiN1bI2rcSTE4Noi7F6DgEzW
uHyTvRk4Km1YMST/5H2Hp9H070OyGKiJkOr1ZE1YgHip0nnH415QzT6P+YDu
PaewM1IRYOL923fATiOfHPEJMgHqhKSOSkYOPfSGs7BJUB6Lrib4PTVN6HDW
eawRwHO6Z7T9FeXWz6XEycWLrLY5ea41cn48Im9+vG+9dOePKKERP4fDlnIL
NYMwTAwEnOw6/NuNN+Cp9DbiYI1IqcWca1B3m/7k5vh0otEzoCxKEYy3wzEA
cuopyHBsuGoEQRkmwXFAqqGZkTBbYlHrxTKKimdhpbwGM7zqQHfjSPBgAvFV
2eRkBBmp+e21ned/4vvQM9IPrxA7ZMXSIDpzTJW0Va9W1bLLDmINgrJF2stI
9cmyERyF9nbebfxQsDGd2jgq65Rtr/e25u4gAHkGQlKEhTLwdZnG7HfusqI3
lQ4XWNJOhkYECG3szS3J8/jy8Ziyw8eSLgvDYsmoywSHIP3tJ5D1djhey9H/
fBOB4GAsw5LMSnVg7jwPmipa+GiFLaTljSi57BqYfS2Hp2u/DxwnnXHTGrfa
deyeakfQNf+KtIGJY6cPO53W8BxcjYRrrw3or9jDUmhICvsTMqBJMmR3ImWA
WcPPUpLIxbRwier25ih8/3zW0yKgKK8MfRT9rimgYvwXYVaggxvabMEVPWgq
FVpWNKq6qmIZb8XSfNyX3BHmrdzEih3j2rSt0kcLgqQ/8mJl0WNoHjHkYi4F
ZOR3ZDUs2oV8pjTuqBcTEDnLXxvD/E+QBtKt77xw0zsNORMHdPqnj5J0Z1ln
wVkkHwEUPtHrhfv8YsaYYxNb+++c3t2gsDlWr0T8kj7D2ZndYZaA3/GA3Bnp
LW7T4ODBKEm/a0/SzTxYz60YSUX462aHj1ki9/tI67l82n0nw5Rcpxs1Mvqx
BjnxDCssGrwkAbb0G6gHEDMGZUTBq9drG7zQmBmaQvbqrsl2mIeoZW00+yUi
48iffgagH9KqvXgTHLdgk5arXBMf11625C6bo1CEQkw4JTNINg8s/dK6F3QX
WKyg6F1emwMCX53Z7bCJ0WU3RnfTnvjezmJiW2TmG5b44fjYmdx2owfBmLuD
wGMLJwOatRACIxrbcQYgU86bH/o9obyU4Q/wfFh4IhfHIGsxcItlvTkCYH25
7uiu3GFEsH2bKgTeOUXKsJ0T3oQMHRV9+rkb44KoroZ9q3pI/rIK1yqDEFU4
uNpU8oppmZrRhl83mZxstuzedQL7F1h7fRe0dwt7JNvMGmkGsvtPMowNdKEd
jo96iLy2YWC0Sfqz3aR8lHmWkChOFKnQDoaxnICwsagtJkepwA1tbYc57UNM
o0qio50K4V765O8TrjA9LL35DywF9OwZof2q1g96nvw/wq514+amSTHlgRvm
bFLbEEfgUYIx63a6CVMhrmpBSAQISGsC8vAJGorhDm4MdqFGQyVwP6zrZD2D
83sVloNGKm248LtOW/Vgof4ffJpvS1ZrALWv2tSjKLZT/b4KsWh1hzch0EUg
mJVkyedDX4EczLrd+11IbE812aFp/FTFbVWPFtJQBQbEmf1l46oL98bhQh18
mO/ODfTlipXN2HdjVIjVdPZQeefpKyhhZwZ9jxjbkHglq/blo/YX0xZyvOcV
xx9PgeUqAcX02o7dp9ZgFZ5ZV1D5bHdDEdizydMje/PjJIFdBS6A07aJqRRT
c0tNq99yMyjQyF6dhpLDSxTZL7Uwhb3riRv7ShUOCMAQvEURjCh9WcwiE4DL
g/STob2ezyWRZpGxC3v3lu0xhV+BBP0uO7fmOv6o/CIu0Cq3vNaUx8dHeQZo
A/79n5Bv6SKQXzAXGfBFeqRK2zuxRXpYYkBaClpE3/h9RY7yvnbo6pfB5AtD
67zOtPI5zCTSdkT/1VuWv5E/+6i5gfQJD4yHR/Xk7GnX9pzqZqmGHDoYu56s
9BEfZDLs+mv55FDQj6+0/dpD/RwBPF7/zNyOs9PzVHj0Q2kEQUNsLeDlNQkU
tJ1sKdfVJaQoZDQLJXmFeDlmqE+OH9FL+JBBoinGFrMhawr6/NrtLEKtu0M3
aqDdRz1Ig7D71oIOQ0Z2Oa2wF0+MQTQsP52pmX4nvURj9QmPmdrwOtRR8FGW
o/4I/E/8s5KKzP+E0nSR2gf/rmamjyC78b7BV0iiMGbc/U3UUOnsun9X0tXN
YPF01aI65UiP9S6WIu90fWdrXZkva4TUqRhtS4kucmVKBi1c6ErnwNschn2q
vuv4VHPuGWIzH1pHkcWaW/87SgEjt2BQvG78E5xIkBYMAxUxkFDx4rQLNDe2
HgfQ6bNPNPeAThTUlYWUUVg6DFCnubGjQDQReRUVuIeRPrUvMS1yaY7vYpSR
9vYhUosyK3zYt3LQSV7ah6TKajatvA2gWJqJzWUcPnzYeeDLz9JS/2pHdn3K
KREZzbz/P46cau7baf23+sTB3hfDLG6VOdWfkkim/R8fZgJ4QV5F2exmpMzt
dn2cDEESF3572HXvWnMo+sjWbHqzhrQM00RB8uQur+4sT3+wJ9NcWPl+QBzZ
L8qbILDYE/E8aF/G/vUN2aAQGj1PbczVhFGDzpcsTKRl8v2bDnf9anVaFZ9s
kzt3xwydtP1LJbK7Nyo9g0ItH0PBuqZheow6DIgVxknwm9//zyIex4Is/+/3
dD1GP4oTMteZcXwnsmfQuSwGqKrC1Bx7f9Tq3WIimGHddByXxDxJJS2gYRrJ
X+k3cRP79BkESlGqQ/mod8ajpVMvSdhpxzNOBwQ9ydJaMxmoFJaCrYN/uutP
nuKx3KhQv2hSsjNBnoh3hjHZZvVdKe8hvL4+JnEuoIPAbWvLo14WrtNaOkTy
150JizMUVuvXbggfPFg7g+/sDqYEUNSaGblTgcaIwFITGl6h1SXVcgi7cbze
0XtplCiGr5+pnC43DF+pmqexsu3C1TouRdm5ofKJTbS541xu1Ztig+PCgMjZ
+mXwKaU8EYYCd7zqg6h7jvNqI2kEZxkK6FWFIytK9pA2/tJQ6d/a2saIhmh4
qEP/1CSsni1jWIkI3idtbhxDK7X5VjETvtz4x1MBcCzejQ6XIk8jv8cTJPJo
k9/acLpRdiKKe0rDHESoWk4gypUVlieOFtxMlWKbnimUwkAiTeS4IDCIbaP6
K4OsfuzDErJ+GxoAU+g7bfjM75lUvH0k7kw67yKm4/gXkRdq6ehjM1nmSLPe
Ep3v0RpYnq+0KGDHmMP/DhUVVjPOB8i9EChKZuiWwinLw102Q15jqpGxBsfW
tzSBcO+pNGVarwdrLSeDh9gp+jSdVnrszoriyImKKQBEoowRCAsgIHSC0sdp
q05UwsTsBlZpznxc+zfX6NNEkTaQDsFtoVkO001uA0NCbSNL0TS4xPA/6bMO
tJX+Yh27GmGYz2D609d4fhXUfIj7Ageeb9UJQS1PcLWuCTCMjrgR3s6CWo8v
BQzedgZVb3iDU2aRO4hfWWfrmzq/C9zB2/lJ7wleUkmcFZaGJGWmqt7H10v5
IhkH/tPrRcE4z3ty8rJuchk3TsAtQ5F6j9c6dW1L3tFfqv2s11TP5eE7LZ1o
CJoXQSkcSfaVufwiBnwOC7CPh8mu746Ouw7ttKLV3P5vK0v8K0VGY6HPFJ61
+9LdM/WCPI3kSGjoo3dQvgKU6BmvCni3p2ixr6p6HA/3dF9P6TsAcoQEUWHe
XVv3eTunGJbSf3actMC2NAKb3sx1ZBYwXHtcPnT5OBeci0jD3JUx/67sAGfE
XFHIokD06Hpk5Kkb8FQlGv+tN/OnQXbDvTGHnz93dse9snvi9HWOOjxik8TN
k3CP8gy8P6g/G95j6WArQUde1srA3e7DnUxw2rYiP62nOreIPhIfoboTQCSM
KGjGiq0rJPPqsDaNjJfDQCFY5YCvLLw5LloaVwaSDAzLdeSL/PSLSgS4MrM8
oq6DGrQxskN0mNiQj2zmNx+HiEYHoGQvcnai38WUh9ptFxzXFDuhS0gLEhIT
ZhwZN4j1bhzddQIhKRE7Ln1nWlticatF2yLmPfPOpEXqV4F5gdn5tajetVa9
3yCMRfLdfkugN8idNuoJvwTNVO3oHlLft+LOBZ9Im853iEfiIs2vcfl3G0gq
DNksd4lhCRbdgFO+tfS9eT+dnUe/ylcyAfUAPeJiM57jPn/hKx+dxmUSoiE1
62Ml+iUS5nBjOzv15ZYEwkvkxvf/Wf/R4AvhWxOiSfiWojj95pWkF3+4/QQf
x57S+k3Zdw8UyMnAJeVD+NwBMBbJ5A57gaJONW/JPktSmYW/B4FIDrgJR+YM
jNCSxcN2ljOLhI27093n4G8E+cHSpahr0yKvkmdnFkUZvuv4lpFT0V1m+1qT
E7KdtWE1ngkcG4YXXxsknZCHF/4uF0sSNDQPbbpZuDECwzlbTYZRIm2hlmIY
L4tur+Og2tmwj4yIsMb1Ccw/kWWvLDZk5YXWvl3yjmkyyGkqCo35PFrD6oxc
AvcIwFYzIKiNy6SKMUe//nERJS92rBdGFP5rp2TgKz872mYwM4XydWflZcC8
9r5CDxS1planEIgE3WD7UOpJB9WP5kSTCrTMHUZyT2bQL2GiNLGx4ZrYCg7n
kxC5DxiSD3JnU2QndQ/or8sXP1nRXq/+uQKT6JhWMnoRT3gN/bebisLB2tPu
Zf/gUioBAteNPTk7X374MzC4Y64z9nArTieauaRye5bOGmOB15y5V7s8lyrV
med10Tgp/KzA+rFUiLn59sc0Ypj4WdNNUvVpEE18XPgH56lLpBCBm1cGNWm2
aeKyBcEUikWk+1M/7FXDW/SAy+w9VqtfqsGbLTp/9ubZCbIW58ERxC/o3I8d
qL4cfHAEJYB7EQP4E4AaADSxatiIRP64JUSmAP7Gmaron+TEhgs69N/Vcw1l
vq2nbf0YLqbuZoIJo+S6ZScMzoTTWZoy/5BmammtYzGqiGE8mF3zUfoXb5ey
hfvD4FiCUtp1p6u3eomjoYBF/3su5+mySY82xCtLp3No8TKviLL0vuxBD2eG
P+G0F5rSeooFgfFx8ZMwx0XwV9zh3Idb3dwbkSMmh0j0no9mP99e48Iy2uU1
w1DGck0AAXIi9o3fZBoSslShFotxEPxbU8LXrO1iJ6IPbRWoON68NMDmniWU
ADMEjuifBZA221NbkYb0QasMtyBV4OHvCdCqnOFe3kDH5q2l7m12HM6Mxd8o
o1EUrDy9u4aKGJ35wdlaglyVoYO6b+XAl/qvWPwm+6o9PA35Qx4vGKYZU1hy
H60RgqzlD0kvidpdG0/9teAYTTGgxhy9ITDRY9QEDLV6nWmkVV7bBSUn4MT6
BR5oeC3ywLzcN82SUvJDCu+Auz1uZc8Zx3be3OPiMNadRNk6FweHbH3vDYRA
LQHgMuTJynwHEhKkEpZlI6nJNdDQ4Z3Kufb/3hwpShJ0bfspsftrKTagZJmi
I4xnC8cQazR7gKX1yTu39HSl1xcYTIFvKT1HFh3lEo/j5r0EE9wbu6a3dfuH
jdnmM9IltZE/5i2Dbhy1Q0qqGWVx7eVfWgGjirTosSnq5qtjCqiM06hYgXlY
NlG9BgHJ1fvMgcERefdk668g9MJOrS57EBNGyTjAhc0OaNUY/lLE0C/hXvqv
e0tEml63+sOkdB8TR3Sq9y/7hWZjgiSkchs2td+bzw2T+9L/ucwp/sCs5yfE
ioL73bM5tDZVhivjxL8dl7Lo8/4pWq00mN4ruWONtzThdr8hDQOBuRBLsmPv
zGk6wEn0IGWD5S4Tc0A/6pbr7hb3mNlU61bfoiTnEV0OJTgv4pfRxUPyV1Sd
rpQ/It3ELTuh/VZExxEs2jKp5RuHVwZIGGDDdFDXq3WnfCdQe4B8pKKsaQCV
/WrO2k+bfTpaaGuwVXZ24Sw+bYXYkLsaAlzCK4FhxuLsybafZJkb9xojJP5a
78mixmM8Kd37RB0SbB8wZMmZPbXTPHiZYpvURyBd/QjHh9UdQf27PnQec7UL
0aMDq8wtqvdILa/sbI00RfFNQNDt9jvMrRgBlBMP1Tx/nRK0lz4UfiOPhaPO
5VVkvgAnn887d6B7ENP3ewdGqK0M1HBuUTp0qjAKQxFOGvpm40j06tp+R+VN
EYR5md7sayxdp4RncYnbpzOjBnmb9XnoXQY1aitcITUc+r6iSQDuCboBRyJL
dcGrJyw+zEjPPJiEF9fU6n2A7VZnKuXUtOv7Ro/2WiUw5FtPlWYJnhtx4xFl
bG3CWBfokJ41k1veHVWfQYyMcwdq1vfpyAM/AS0JnEYVsXR7hlFi5k4qm7SX
4DOMDIZZfZR0Nu6LPw0qrGaqoSF+kTd3MjAMXwRm5DcbQEa/va6q2tr1e2AD
LQzAqpEfHAU0zFIt0iIAxW+jYD8tlLvycycVYbn8ywyKx/1q4C2/Co6W7qsY
1kr7q0T0mLCCQN+/IHaNdSD8sTJLZ+6ZwVnbSsMefchKa/usbSbEHK0hW7df
sEuowgVkQWqSrBpxjhOS55ezdxSbjY1zNprqfYM4wolwSqHEnSF7xhAxT4RZ
+2MEL9iDMROBo6VL0r5xVKb+AvJix/Q/QL/O2m88l+HcavABh9Lmd5Hz0FtH
bS4Cb30NmMvfDJtyS83YJh6VshP6+QIfl99nHjaCF8Lo6sSuxN+KsMRi4T82
VgBBHZ08zTApZJ//WluszLnv2pUJ6O6heSYDGcvG+F7x1v9yimNON5jJTMUG
JgdA3w1zjYArsjzEFXlvJqStn+KP0RNtN9v1LecEEjZI74VmGHLSQCXKSiFT
koSwLpw7oJ6D5UYBpFdErufUv+J5Hz2Eeleq0DnYQXvB2DWe227npCPjVW0N
BJcZPC9LDcpoVleuKYntQwIrvUInt0erpJvk/ClX5jeCDPysbbmthHmYckMW
s9Z54UyCV9L1WHcpSH5eZalgMQpyXlt2eJy9YhJNzxLOiorr8yGsQ0obPhfd
ZHEdqJkRRICTxGV/f7+n1DBwZi550/fOgVi7A3pWcgfxIu5uY0PGBJsF3gJ9
GooyxB/eDaK69CoZFpIMjeabi2ZDR1r1h9dDmYI/X2yjVSy2w/4OllhpDQdq
NDPntQjABbJHdDsAJIqZ6JdYx1pxdyppKlud3gi550pJ5F8Phphj5zxpriJV
Q0w90jaukzaG3k1y40d3Yku3pp+VKayB23Mn7KUtfyelFVsDsKbP4RfIE23p
P7uuP+b4QmoftMD8HKQhNrWFa/kFBWim7eh8TCoyADjM5pZ4iYyXMxILO83T
yCUWj5KLIqK2Xf19d8PdvVS9Num5Qj+QIe2tO5koGOiskZGfqxjtWXw2twv2
unNTCUctoSZHrkluIsBtPMoCfHLmp2yWaVplygRt0SwtgaoB8RT/7gGmagND
NiTWsatT5yDIgo8qRy8VvJ+W88eDrqWJrrHxjPVDaTdMuzfcfTBBXEmMIH6L
H2hsubJtzFJzV0zp9Nw7MXAI3RgGO5HGu/4UM91jOePeXnTbGm+8IhlAJqmB
AndwqBDKtLe5XvuGLu9XhuL+xPqX5czjQ4BZoDYrYUBUUr2PiGEiYLYHtl3N
q/en/g19xZCAVcg7fbCTRTpbFmn4EKhOVW7yEJRhYekVKPWZsmgxMDMmAfTh
6VTNa6MBQ25j38VlGqw80leiG6ofcgq2t0TJ7x2ADd/ihTBrxmaD1l9Rejd/
l2BQD74uyiXcuDSYo4FT4YeC+SIuPQekaV6T8tdM9ROZLRTveAoBenZ/QLap
GuLFjHsIjxZJyzNIaWBNTPQHtmavSBU6NY+Ha/ACAU537c6LMVQYy3jDbMkC
ljcVa1HK+A8ONqwf3w+3dXG3wVZ3YofmIsHPmub9tHSxPrfr0up1umyxl5N6
7F+XO00ydmdxOgO1fRlkvdANnhqhnF861WUUPgE10gJlyBPw81pJlvf7uRWG
k4NkJkMmO5xql3NLPldnqrUs8cKsn4Kp8+X7vb90y5sLiA0wNwwx91/0q5Bx
mbYXxJVkffvfeuYjjD6377vN1+Hik1Y4skodKqCwuQWlSgxanaUk75G/wesQ
hq/MGuRC2xj4mcN9LQmCH9Dfna2ve7SxjOrNYQcbs+JSrxb/AQX7PN9C+ne1
qQXSJK5HI9SORp+sn0HrvXsgZwBewgf/R6i+c1FDLpVlOP04exOfJGDf4nDO
xzFnTI9MhnGLXAsmBI++9a+YApCo6ojS4jOZM3tLJaqCttep8WPeZNPY1cGS
gHIo14Y+DZY5q4HuoJHA8UUJ0mJultnGAzpX4fh1infelAm1d2giJGNtBNuz
3RsjFcJlowgcJioKGCmD4KN4TgnsH10CAyWZTe7mjx7X0XbbVQTmgs7XqHDB
DwwpTnMe87c1HsYaX6jv3G6E6hVg1fRuOo0WNr4uh32w4ZsjjiLBWuCC+YpH
RBG0Fps9CjToU4HSEJxpGL9ru8vy8h/OcbN9WpSCB2DqFhp2pLVDK608PJOv
rJqKOs6GrqW+UbnSwRT6o7qy7q5HA0RH0jIf1hhMngK+Nc87xBY/Hlq0N/zN
IZP7BF6lJyXwKdLunvdb/HmLjIf0/fXgKbil0OBhN798owbvznY3HCy0QjJy
YN/YxJqVSWIIFl9Vf4m3ZWUx+7lWpKSAga9iJch6kAk/weik+thQJ9JsvsP7
ER6o4cvhqGocXsqF/WM9BOrN6JfAF9FcWwNhafvEFPR7JJoILDDmJCrbBPz0
dtQsUfa2GJ0mBtLGanUdJaa4j4EBYt0fuVmYe3NhYrcdReAn3dvoYsEtoy5o
bRv79DoYa71i/VO4/pLrVCjJ1gxItvQrpllPcE+lsUQ8SjxH1qwmyVPdp7Pi
fj2At8nvpYWTdnJX+a7kgHQVIAoeUvOy+eJWr+YBTnuIoEMEwMKw5JtNfi2m
fXZhYNp7xCnGuO/qhKNDAgC5m69KOoYLDaSF65pDcb2FUnt2nLLrfxiJW2Vq
qGmP/kIGf9K5gqjUnhlJ6k2V5VDZpWAAhJqEgr63lDcLWEmECIcBX1ds2wBo
OpSWsU5Y1e6P6qmsdHXWh3kmTTsoHWd56S8rGZchf7yKMg+R5gTJyFlmLY5X
ansGeXxCi6ZXPZBLMEaI7X3UzhwlpSY667m3X4qPI6TEeZhj4N+J0CLqzUa9
WnGy/4u13NlDagJKE8Lx9ZTL/iDYX44grTj2ba6ja1tjE25RROISCRMUQEn4
lleuZ7jqAu/kG4VZsT2cW4rmrMa3acwCqueY8zgiJ6c2XDkkoBzsWACvy4HM
vyykOlkiPTtqXWMfLQn20OVycAEozp2uIXMIC+7aOaqa9DVyyxQ0rUC6yN2g
986+wda/6N0W4E0tmsWTgRtJYxVY9JcIUjYHHQtX7MS5UdzSXDEwi2M9dW35
E030TF4psjBqtcSR1P4BJ4eLUaAeASpelVVXcTJeHER76yo50xxAkufS5hro
5CNWzKOviNKB3yE9JmiDmT67sXO7Xrlfknuvm2xStnFR93DJQz9qFDoJqgN9
4rcBmVbn4jPOCFnP2Gq8gjy/v6L+zsz7sXLLWHwVutUXbKxrN+FzwbTrbIeR
HvHrNeATTYiSvh/h0nUkBnZerg6VQYbvfqNlWfrzV7OWE10wegm1bKTyIKZm
8uYQ78HCtAC7K/owOnst6479QErroHjg42/IuxKxKwdtOJLUpudVHbCJ6clR
6j9YZBZPF2nvRl3C9h9LyHVvrKupFvjeNOLBpoM7ITwgi8tfMzLTZXL8sQhG
OO9Z/O4UUuIaW9I7ru/B6mAIx3z34GEYLNrIeKfefJwyOgVGE1WZu7BosviN
A4ZaK3OCIQ58rLgE8DDEs1GCim2ammYBErJVQn48aOu4OPPzsdCjAunz4XnJ
NmQVR9qmE2a8ZKrtgnqMpA+YaspsUPkZsIC+w5MIC2cv7cMVu6lzQX1VtVFJ
xCv2DmQ0Jqc6p9+NS8XCOnYReH4ACLmMy/TkqJDcncN5NDNRoN7Ac46j8xUv
CarYeURCU8+VNnt0iVgouOL9v58CSStlmiaFZ2apTIZPMo0buKU1BDVdsT2v
bQsdGo63X0StH03s9sCdJ4IFuKhUaWRzWg/8RT2jrGGkvc9uCiu3zvtOBWYA
4zaUcdWamIu1FJ322aieUzFTxgIbP3dH597TRrMKfG0hzbx7r369dGpGuxH7
VI7POG4L+X1Qe+z6Sc1BIAEcRoQIuFNv+Z+UBr86U8At1w6ZWm9GH9CX7BRw
AE4ERiWg7TCQSvnCV6miiALLo5cTX/mRcsJgY/NDYGvo2Vw2LKbUezoavPpE
Ltmr/x7DUnB8jQyHarmoyytFLYOxBQtphnVn2SaE/dpeb0dsHvJ2GQYlBb/W
dI2lT8z9pgu9ZXVXmVqM6wxAfSG3R/5Jz5jJXUk0muOe5BPwk403QCa7GUYK
sCEUIiG+QZ3oRMaCisrkUphuRBI0CHuRrIfpByGtUCaBWCEX9axWv3I9EN40
7vwJTII3iDKHEZj5diw/YGADBAEP1oOjlxbe7P2HF9tUZDy/fwzLiHjPRO7S
Kec8Y3Tw4tY9yk/CItQsufA7lnMSqumzYtKOpNBvaMlLw0We4BbOvXn8Bga7
AdaHHVDwhM5ueuDwKq33fQocXqIlwJHlsAjlKl9cRT2fdhyxiFl3/XKBgHjo
XVJNEl0XnXpnu5o+q059jeKXc2MfTkF3Ovdytw/tkcrAJ7UEif78PizR7cMN
/fAJALQLyuAYYCk4GAryefadLOqS0JZyxef9a4F6duiV3cx3fzJgOaE0VeEb
OwUXStYX0tTjItIQnm33l+g1Wwz6fBEBTPiOg8a3uVUrLKrSkLtQ6aPP4dt/
OQsFxMjPRaV82UhphW/mBb3MSObs/NVEqZuGpQr97elxPvR8zvLeQ8QKEBcw
xve5QsDHMcGBnWHmvTGMUmAKHyeeGivo6swrGxEwYBTiumfBG0O4J92nFIDc
oie6kFmOZjnKikjg1d7/88CWJETB9D+pJUyESDKkzpWIjVGFKiZAxo8blZ9Z
DATBvSEETHPoolA9nKJWXCLiiCkbIBsTQnGAfZZlteraJbSNvO8+WCFHVhc9
CFVlwUsfDyczL+FNEc801dxYWG8h+XgRaV+Nggtorn7i3KxtCcp0nRqFJPXj
Pzf32sKVgORVH6WmWlwoVT30RIkg62hk7TrHWWKShimxsMTOKFxTnuqgShvf
3Xt8Y0WfOcJRozmNapiTRNUtwZDCjNL+AbwiRWWHVtTlpOgrycOd/hnC8c+5
4f0Xv7q1K88cv6NXSUzJBrTAlGMtTByCJDz213GBfN8pU75YtwfIrfodHyYU
HspBF+ySHmShvI2w0hUJHSgMIENHNxe6ctSUPvjBSWSLIEtgoEB1CTrfwuta
eSBTLXn66ISp5n8//Hw8aJQ1FZWKMaPfK5i+ezbwcnRSrPCbmRVYkFXkSWdp
ZUeOdK13xd4weGjY0EV+KNYc8QrhA0zO9KlB1dFhzC9KlY9+X4CI3/Tnug2P
QVP8V6MqzBc5/ypVA+ZxlLaWengFrrfoshlWm1IPA8bQ7CzTg7AyXpZYbQkL
XH6Sk7Eeq/0O+1UuR6eEc0x4V3y/sOW7iwCfMZnbDyGl5UfkczFBOiowijEG
EC35QIlyUxvbatgKaFUi0pHjDBnhHeLuDeLnbs+g3KTkHfRBaAhTON7HML5b
s2z70VBXpd43EI1GZWCQ7rdSzm4QjZBCQsxR93tWjpUUhaNgePtL4UKv4wMb
ZBgT0slgs8nzrgQkHkuCoTQW9hMnmBWs8+zb11W8iKs20IphJarkQjfTTvr4
LzLCYGPSTrM3gdXLUXgGjz4jOEGiEO5z5gD0D2AH88igncOeUOhp9LRE9sMK
fwLW4PM3NP+eZNJaINR54Xt9cowXMjcPV5C2bL5jhuyH1b9C2SJ0rWLoe3Di
h6pB+Ew2Cc9Le96lestuKtDemOX0Rnek2Rka/cefKI0gD99IednKPmBR6tE/
p5cLOBoxoKFPWnn7e9USnrmg4KUwHjnC3sPL3VMTBuWwL503n5CNynPVTiIc
qhQWYZH/T075yMH6zhF6iNOvZ38GT2e12XiFABaJhoOZmZa/F4HNDjK4TQ6r
a6YI6uEQQ8/YifbMq+ESbP85lmVGGGmfxKHZ7VXg8G8f7qS3z5l38zJ5czc9
HdxU/3M435YCKgrNMp+zaVeGZFTxs8Dpk5fiMXWqo/dcZjZnemOzHTaRTS2A
3gE7CSA8B4TEyflzWZaadCyAnCzFMrEAYA3r9IRx4zM/S9bo0O0cpKmHyF+p
C/lgv1n0tHIhERtZmQHICn0sOzuMmHB2ymO3SXBrg+wvMHAvMx6Uzwx72lWU
9ldpGIPIXdVErkb917ARKxbDTgTlStVasNJ4QlsoedGHgB+wMjI8liZPdStN
/DwZzlEsXw5QWGv/IakuaNteGJA4TuYZA0A8sftu2zffsAVq4kL6jCawSp+8
AXwozf8Mehq38fggPpUsLvAjjB8fLkojoNxoDIYZg3tPWt/8JEoJsIuczCIz
nI2iduCPzuL0RrFmV1WsYjRtVoVyg2LoDMmpm5PE3sllKui5aX6ixZikmv1E
9rKVZNllL8xJRPv+mjPrXW8jqHLnJelXBkj9CJMSwswT71w7A4g+MriY5HGD
s2xv2GL8GGgSIdIEK6y9DQWkjOBdqT4b/Ni+mOGGDb29gRU6yjyoIXlrw0id
XA++4XbuU1SFljmyPzthFcMOvg6NRixs54euJoO74HIZYYu0JskDxPE2KWdf
iz08VPSKsHnUgn3deEP2epkEMioBrhnSes2eX8VskTL+z05LxLJNHKHLGeCd
eKpmZ8wRP83h7hcR7ZAfRLbtFtNxxjcTyOAAOJMTMqUf1YasGqoJAxAl+d54
9VjK1ycgt0dN+xg+D1t5fNLfTavxC5IT3SoSAOzbaIbWU6992vmpuzsuC3UW
UMQeI02Tu2FRbEoQvn0+AW8NKnI1qM1PfMfR6I8rn+zTS89EnhJZQ9gb0NtI
9+ZVvG8O6/STwQHIcTaZQtRJWNj/QqwtZvDpNlOPhTueBgK1PzD4+NyLZBk7
u1NJp8dkQgiDry84hMq6KTAV/DMpT5Ud0YEzyFJFbFWs2lue8oMpwe717JS2
V4yDfEAmYDV7Ncf3R8D7Kx4Bmm9qy0MkSLYl+J6Zcgzg7/U/GLxXmBCs5tq7
yRNDBFmeLbi8N5C5vFEaKG4JpPmSbe+SynWAcgGU1qTxsiRNuHvOVFxBWBBc
atQdsvRbpljg+kApORKXOJwXxzOtbs6nBEKKYRZTj/jlwjiAJ3gCMyWYs2cZ
T9tEXSa2zziJljtyBBVAAYLstwTN+YP5ShI7WWfPNE00WCc/qRXibfDKtjDM
92kF+j5Y/4yh4h/9vg2LlLxRt7/xPO/V6RozdBAakd8JFdRF/IcbHHq4VXjq
5W+KU1sQFyXH2iqco6bAAA5FCP4XwuhmA/y8dBBCsQpyRU/SZQiFZ8zl3q0s
iv738jEuI67aji5vNTug/KL4eY+2QtrGC3dT82mAVjiLn+7raNVZskztU6cT
L5KXgd+M0Iu8ZQIVysI2NF5HYvnAl5+B8CoK08qpP17m+eD0dhex51nAV7zK
A8+cnPTs0HvTHA/0dK/H6FrUH5yns10M7kABGBrn6A0Ff3vCHQGa0sE/Bgdm
EfzYE/TEzVoRhjaoAf+U1NBuyeRi9lOIPDb2MFsjz9eNAt4a9nHtswBADfLG
+ory8jNM6H9nH66AQAD1lGPSZsaDEdfUn9jrfRO91VC41Z6s3XaXg0k3EOSI
ozIrFTaSK0toKUvFTIno0sbSxSJyi+GBKShH3DYaHPQc5g2Q+yIn90rkDl2k
eIUfevnLaV9c45syqeM4+BALkPqkriI+41y7Pkx5S5T25sVKBzD7HDs22HbT
n3+hWIuJCb+7mCVej0NOgRARl5SeHt4Ybd0EdV5/1hvs9Id0byT+PLZruD1i
TyxtBXRZGPS5atXrJho++ZogDjjRtPFG850KHfhxkSc31ro7GsdicKx8wT2r
0FIvkqMU8w7GjYWfwXFHJOho/FbxEUJO8ceVg/3tXEhP921lpOsGJ5hYyCWM
SHWBZ8gjaavp06PjVQGTdK8paUefSJgfT2Dpcwu1gX+6blzVbki9MEGtWujI
JGScLDKwrwkJ2vvh7l7bxW9LC09oLhPSjk08eAMomwYZQpkmSX6aWCPm82/9
95Y2OkZsBO9+zduz4JGFum+ED9flo5rYWYZ2HCzY2waYostsEfcoZK3Z0agJ
bOYIKjkPJ9m8WLpzPiAl6htTH6kiXYn7hVptOvmvDFdMM+/oj8LZsGbuxcQV
6IKyIg5XnFuHTwjEtPRQNIbMq/chIuZJl2aRSfQvIZEv4Nsl/b6NG72CbKvI
ZOr+I8fhsDfRV2YS88jX1fbY19x/smO10WOXeHQmHzhfaNDgIxNZ16bhrz0U
OxY2TOPbTF9afLqns60tH68ENS/mT6XG4z38q24THzxChmf4GUvGdChhCilx
Iwy6yy+RtxNTPpjouW65m86smKZunmNQZA6kw++lex63bSbFYukB6CebPXvC
wRY/vjEz2KnbWqBQTfRUQEPBnc8HAT4ixTsjcKGhQ2bJlaXxZz2oDs/9ShYS
mhmd1l3xlG6/ZoVRsZNmmwARzi5+Zij6io5cl9ysvyBt0ffLBuwk7Vgv8HpU
N4iee8A2Je3Ypbb0bj1PSIHyc54pVdTA+fMVLXvTWpiMOOZQ17U6F2pOmp+j
hDSpT4bSMDOdQCQ+SevA4HdFA58FlvL/iVHmVBXRDYJLit7Ckw9wXDqP/+tU
3Tevk+Hp8smt5kTbT4txKCihA90cGmU26jZo1wNuy9UykJoIwUi53Ka+g3FX
pnwpUtIK3b+O7q1KuMHCKdWRAjtG/3xoEChVkJWnn1Dy7PaPufk+tpv4Ragy
EBcA6B4nemsrXUmiFofJiB5Yf8/atOj2yRBPmap0GV30+28WAExGMPk0stsh
ebPp3jZVF3mHW4++t2Fj6sjHk8aqLGKfvufl3cBoghVC/VaTDl0DjUgYIHRS
pp7xJDN6HwN/aNzvEhyxhWUMzpcp/frf5FY6SK6ZZ/T3fOo1+Lvw0YDuCDCD
1Xofc6M6NowUPILKB2cYeM3eNBaPjJQaqQ6K/yQ1T9JQnCPLqyanZrBUIpgv
ad+7TFFujBzHkKzdlsdn2KRNp3vRcQqz5JkaBJgxvjnyBcH5EPS9+51PtR/n
JR3ERJD2lIAnKY7vL3/Pjw2hrhGWidBCSsgjoh5COrUt3ubY0xVhTXVNjsOH
wb0GetoS/ohvnmRxuKRJSA4rK3cMU3X9MNPdn9yP529l0RSnET7KPmgn98Yi
7sza9hQ/kOD9sOVps0ChpcRDbQO5NwHKxDDC8TeZ6J3oK03CiRiqb4hi+Nu5
jeTOPGDMQ8KoXli0w425FrYEsIaGEIGkKhdk5d7mKLRhiAt1oXLEgiJIP2mS
O3gjYd68Jrysd+JvN19W8tUMR9rBjcVz5JtQbM5cHAg6urGjJB7VKDEEU69x
pgiFVREN5S3wPnpiIELMPHtm80GCqTPqxZpDnb4skN0nBIiGJizBkPunWVr6
iM2Te+P5DZStmBaDLZjQV/LI2/Zc0TdSkmscPjqDO7cIMrm447aPqFwzxH7D
a/xyj7k+6GWpVaEiDtbxQoMa++mBO5Ph+q0Iu0wt3kAns26Gqsr5vdqpD6Hw
/KHBaxUHvqzejwBhFEC4fCiSDXz/Rca0hHnNAUBaWDHOtZjZyh0sUe8Lcfph
v9pmmyFXL7O0rU6l8NmwOhPH6lZytaMGydlz6Iu83o2FEFabynuvGkhCc7r7
8evjffcuWEgqn75Oam6Vna8oys8xKtPiH5DdKil7ezlt+VCFI4sJu0An48Be
K2jhdWlWHnUteUUN1ai4lAA/Sp5FcAup2A6FdVWjKp6d6h8X0zwX0NoZnWHr
qHY0XK5he1gS8a9akYfYny2LEVaTiMmT+wsLA7WpFgrCFnaW3k4bXu/t6jBO
E8bSuvWBz4jPyeAPa3gtTLNBeo7/GXvMPMRb0Qnj3Gw9yyF7LaoRalvogHU3
Ihg98ufyGTv8Ab/dZ67tjVUZzSV52+XvbmVubIlA8NQhbLw8nEQBxfL3/AMS
b/DzwrZ9T2M+5iW7M2r/v/KO/aBsUn1ERFMzsbPkoL+Z9mczobqA6wIaIkny
yZg2fy+TLmufWEtjUbC+EOTtelmAuXu7nV1m/WGf6HM1gWtNpnDhshdspl18
RsSWSDVMdbqvMT8mAn7pKdUzUVsZm2YmQwtqMAwEqM72haDW82FRO9sseU+h
qozmRBAFexlGih9Bin6BN8SzdWVfedrDXNcoi23BR5581PhoOE9P20Z+6p8Z
WTEu37QYsui06shixX/Yn+8dRicaVwgpgVdUltG91kDZexLI9WUr4o2PECXe
M9hif8SiG4uXfd3yOqTdpioW+n2UbhvPNufirZmrajo+CsGhOwODAJcIWa/3
wY5D3OpI1Q2gSiGfJtmz28TKZuASaahWpPhiqjuBMaBHgR2R1cG3HFzdEIz2
5Eu5KHo+K+OxBI3Dug0AoavlAkTwn5nnzccAIzmlNuZ5nZflr0g58SL2+5cD
C0rKrOBd8iR+4nBokx6vzVlw8wReUpExv6xn4R19ZV3bNwEIIF1GwYs5Of97
WJyMFN2UfgVcE39u8w8dERRDO3HYG/6JZz0pW9sUppoOsYxRcQV1D9/d+quQ
o4cf+4dw+HzdwV9wOq7V9doiOJyXJdWpYnKo68YPz/BYiA+EtguAB2wqxS3N
8xleE5voX27IiJuIwKDEky1UUnPQjAoVKjD5vxRWdwK6BEmkv8GxWODSWffY
hokmDm8NNOg3yK4QGeOK020nx/j6iC/teEza+ASMlp1PlB3xHW4gmsSFdvb6
TgZAjOTx5sT67i7zbePuTkDA2N+dw1dcfjWiXK0lQrJcENCvwINj9g2x7O0i
rPRovj3JIun/PNe2DKdIexeW5Xu+dtGf0r11hAN01/XryabtN0t7Glo+Fivu
3aFrCa4vvACmSDzOaxlng6StnUnclmatr/svY1aFSUMnrUA4TJ8DbjbaC12L
49M28eAP+Z0AyC1ibwxqTkN8NN61r76SFW74yygvzalRmFbEJ4F3jmwpklRv
3qYzDifZlx3pJa5SdUcg5ZyW1w0urgdKrULqpDorYfFqusJFbEHYCC63PxvR
rjaNATTu8vTD/5Rea8EFjJKc+8LZ2T1vsEWjUisGprQZ+KPIPXAs9VfhcZJx
8X4lyNxJuekRWr3b84kiSgyLZbDADFMziSzUDTDqBb5Ryph81rCC0w6hMF7v
+TkuTIm12R4taErJrpwjLEFLkmq7paUSwp4+OpseZamj70+TsXgKwaGCkeNh
LTDBoKf1R7YiZTps9MOTEFVaw9928JrhKGc5WsVjAWHnCWpA+b4Ql+p7PciM
Qe1qyDS558SkI9HKGCH4soRFL8eAJSbNmSTVhTvWcF1ZkL5CBkqkL4W9KOSd
efDPfVvg6/kmh5V3mzMW0X79oIwcBo+SBKdF9qMVrlC0vHXD0WglzS2S34u9
Npi89u27eYv1TdoRkBEVRU7lUjL5nM5wAumw1VlNC8Wwl3QAPXiJ1IOlyjw2
e3hfdBbna/cnE7+LbJVDCEj2+58NE/t+JLiuQkLDTyZcQ+/hugds0A5BxS6Z
XmlozsVnrBFDJGFw6VLBrrurHf+gHPl/brT1RKhX8++tZgSowEywxS+45hsz
Mc6o1XI+12zJQZJOgSL1I3pOPu479y8MQzJVwsz/Oeiyc4iisDb/m8lh9CmN
MRvGkmqgbi+PN3XREM+ePcAw7Lrdbbo7chCh9K7xQ9jPssrZpK/fy7+LZUwt
rQ0/YcKgnhx7h+E9kLChdtWneiC1p3RIJOiKcktrOOvUmXs7sJEUEAir1X4X
ptQ87J5mner64GJ/kqpTYVSZxVstF+X/bPD9YblbNcjdDrjrn/NmqKSVvzBR
98gIkrbgDe0d27CVieR8KY/RduOkaHzDv1uuHkr/+uin1YM4hLAn3yiqrLM/
NL41xvT1N8VRtJtdIG+f1uMlEg7hdPeRbvSc5YV0EFmtMSkvqSlOvIh/lkQW
NTgooPcnQ7PukNQbI5m76TyXXZxx1auLKUN8u4ZDTDk0zKTTmiJqOkdxuQw3
SKqnva4wisBgbRMyA4YEJokgI0x56HK37yAtQTADOiE3ZlNbGpRhbzpfm+Oa
nrcBVs01BDbWgY8QyhOmo/+CPBwKZHSn3vRhOcKXhCmneddOfDBNz/Yzavbx
CHmdxB0ePaDgYADzeGzGy9z1ZKitTGP70NR7GfRMzAEM6w7VRaY6KTvF3wsR
yma68gdk4vnOtNb9+nYJxPAHHiKNUuHDL51URXT7FHrwK/Bx8wv89PjyYRcV
6c8d9UkyCbJZiPQIWIgH462CoRkIW4hJbh9/c9F4yzx948mGO7iuSF1rl2bS
7HENYDP1sProF/N32XAXcJxUBSkFOvQ3u1IOV4jgehcIbx8tCqcYJ/QhGUMv
AYzcHL3oObwBqMSj+L8SluUXLgxsrhdUcBiIkIWqOJdxrBsaVkR4sVUtz4mg
g96Li3qEmQrQiQWCuGycG+u4aVN9xoUl0YlR7Y3veUfncZrKlCIb/eZUbxdW
h/BcpL7gs+TKFQsRsbgp/+Y6Gkr5DiY3OndFaKLgHOUJRX30F1AkmfkHEgK0
G798QWdGEiyRnil23z7OZ0LYlVpMhgaJ1ngADvBXr4wpmx9C33lOuhdix2vc
NnItiDP10VFGkM/F2eD6KqAc/boisOGa9iEfq9AI5QhlQ1eWcl+yRdeU/mHj
VvO41MagOmVNa/82h4uBMePcY48Jxv1yvGmbQqWN/566XRkNdxfkaztEPR4e
KwxgfK1laz/9Ek19SaQ5v6i+5wojCskV0v8Bue33WM1OAPzj4z50p7BBGZLz
Cqh7TkaZyt/4GIS3i7toudrdMc0lVDV4a95+WR1Nrty830uQImm26HgXcZkj
7IAJETlXDFqcT3ENwly4VfIxG/0zOrBdxAKj5uQYj2EKvKY0couRpxIlvoc2
TdCDDMNGgs1SlRWBXU2K8BMAi5rRcrGYdjBLAEYE3m+X2853nQBmymL+nggj
YraAE1eY1wuK8nykRl/IWlouELgOjZJ45vsCuF1VLCzi/X/3HskM5QVtQZDY
gyll0PSyEbQwBLAMHxBFkO4GdFIro3MKBkLgE9CZdTYIqko0bNHZFU+tjCK1
KJNvClOgDm6MR0TgAdLBNRbsmJuL3ZRUEe6wo7dU2Ut0WN61iTK2dZWrOa0L
Qg4ZjXvQHNKeZu4AjEQ4xkod+0QSLcY8jGqCCHoUGmA5BJu8l1T97R2ZqME+
qlLP3GJJbOP65KYVdylOUMOzx1lIgjolSAySiHZIzdd603MNujTpr9ar3n2C
Zevy9fSEsAJx66TPhrNbbqpa/cTc54gM3UHEBA73GiT32ZYcml7UAF5Bb+mD
2yB0Jfe//6u9z+S2h6k9aOCc1SALGYa8s/zO0DrINw9CHFJDtIu2kF0rWlr4
XVAr1Z2nooaOAJaHPw48s+suAPAWSSSQKVEhYqqeEtRDUNH4rjTseF7w+YCW
Oe0K6wuj7ran/YEw4s2112fRp410y2UTq3WNwRr+/oJAtEC8TpBsBP02jGkX
9Qy3fVLdIayX9j3Po4rqxhGOrO+Q5w+2CO90Sv4Jij7azAKIJrdw2+Y816d3
afOwFBk3ikdavHyiKzxBiUM592CL78jwB5zZQJ7oHiERDp6MlhjUsmGxjkk/
Olax+O36yXzTVaGinYZNsjkaXusjXgE6KMeqvjT36zEn70T6c0uujaYSnTks
DDA9RNcscyCusVeokQJ7yzUt+I3gcTSvaIhAyLUuk4A9K0/+YtetgYfm1bHJ
0cCN1yRZs/6918w6PEIbzbvhePjwsEVYOfbBiuuuPYtHGROYWyCxFKIWlSsU
C13Xb26+jw0zQO5KbqiqBMbbVa/vorUjDyCud8bpmMjImjur3T7ydo1OCx/I
N91KiYxxeA209dLlYoGwH1vWGtKHkdLGcfNYdNewKizrVRponvsFUOvgZ8hc
jWPVI9nB1WLy9VP5S3FzmKpqvZHiUC0HY00yPu00SeqNHb3jG34O7RVjr4LX
9YiKvHMwiEm5liQqmI/SdD2MmhDOpygqlf7n1DbOhdoPHNhAn2hBRJknSSgl
SITIZIpZGjm2wNF59wCneOlsjHTiz4MuSqkDNDRB67EMYeJ6Imcp+NzwQXwI
EfYAhimH7CjDxYZo+iDJbdrTNijv8yHz5fcg5F/ZtV9tTQACG2wGQzZEGb8T
sU3FB7BwU/AHNpeUVCK4lUqSDgXcMGTPc54tXiKfw2iP/WEygiGQkfk8Z5by
SgSNNiaflIq1xl9NPj9wT4tP9sVs8QSXVR83oJi1VhtTspQtQ6U1EGQjaa7V
/OUL4R2DUu/NdZ/LeeihzbL1w/Am/OJHz5JfRlCgS0BgrH8OQZiModu/v7Zy
WEBGPb2Bw/0iixVfJm1M4O8SnwxydITqHziRxCLd8mRIy98C8trxQkrViLVT
ZwdbsF28RdShptWnsomiLpph6r78T5Y+T40RXlw/1OmD3H2hklUBQ4Vtv17u
wllI1NgWqkeF9TJFn0iJ4hcNG7RnyOC8PNQ2y3CTQo+tmU7v5UkCj1l8EFjK
Yv+AE8dfHOmYwSA/VvUaWzjX3ReKNeuzT9OjcWr3UydQyvxW3DkyWR8/hcEM
2DaY3TW+SDYl04Piu9wr8WTCuE87OqFp358Nft5TXIeocisiWfCI6Qz9OqHs
gHPGvLDMEuj/m9YjNeCDFcXsESb1ptgyGLlIWNcAZFcYxDzIj+McSvXF6fcV
1SUtx9Z5iak01srU+QkSPiwQPy2gWwgGaVdz/7npqHjDy7/NI6pDhfpnMRAi
N+loSH0RE+fsF2syb6up+IasBw9D2fg3v1pRVsEc7NiPN/wNSb8oW372NZas
FFtS2qygJBLrytC0lXb1Rzvqi+75a6kiHocf6F6CZ1AdxXH8MI0cD0V2CuyX
x4bafk4bzLy0Qx47QEsxKb2IBijr65YID3qbM684J9mahfiMC420KZoEx/PI
70IRfrel71RLNtDKCD5vipPX2GllDG1ZI1oyn6LxYVYEAKxdAq9hEAPyCFX1
VpYtARZLbmwo6sLKuRQEQtZFM6L8p1WYNcBEIY2q16vsjDSxE2GF7novNwg9
qVCQZE+AU+eu7Z/jTMxs2UlktUS//uCG7Y0Sn1qTKXWyLEKOceQ8Wu6nEe/0
20UbrRnCeJ7+Wz2MgEx8Ao4DQ6GJwIrNPLWUS8mc3TDlup9C1E8KUwUwtDbU
8cfyAwi+4LqdyQRKDivy6AhBsJt0jOo5QKk8V49dXb3e2fZBb/uMtcpDRnIf
w4+8fLCnCij4jmVQ/exqWIkjR5Hz2FjeLqKbiXL0gzPIAyn1HPxmhbwuC/t+
CmMqsRNiaRUql6Ibm+mSVUjCAhpjqfyx/BTpW+IlPcMZdlqi8MIJPcgyM5CV
JOO5X8LxI6SNGeMROMfPn0r8b2LRctDuBVANCfk5SkLjRF3e44JJpycMgHuv
dWAJMAOcsu6TqH5CKKIvjgeD63OnpbvM4oQB0k0yWmt19XnnI21/ZHJnq1QL
7CdVotgZCUxuaBHo/LWtObo4IWJ09JpoYmMT64kPvimOWt6nccj2Imo974bR
5vmHz7qvxUDnXQePzQYoq51DmDKfjCxBtL7I4M5zCOHdNOPQ/e6nVAVbuuf1
7nQgle/Nh3jHXmTIVuuo8Yl+HW/y7AUa+HpReInkbVjZOMs6BlJzsEvYOeeu
eXcvdmjHxXrrAbuF75dhvchQO92kWKvvteNDUaLdd/iuRSKueNZONop7s7jA
1S7CD0AevknHzCeRpMnsa3jvPt2JbsnEeOCW361taF15fevRhTl6KjV6IQ8n
E5poGPMajLkb+iEpwwF6oEbZZoXomE7rBHVJC6/XNWFw42aB5myX20vQJQfY
qeti9rBpDtlKnxOC50W+Gsa5njvWHADE1gA2K10+DCKCMUzRJsKdVg0KLm02
mxkICeZts8L6n4hoI572cm1dxM0l9xx4AyQUu607ktNbA7plon+TrJ+e9yR4
NE8li6/3sbWZQwcJ55cfE0d/nwRN7kP65RzaN2b/li2y29yS51Fg8iygMW1D
XLg0SnfaOFgtVL44YiKgSvf4LLGi3YH8Uue2PobWeE2fQpxoh/5HABhCPrZI
bAcM942eHfiGWGZWKocPoHXM3MQickSCI9nbyXGwznyDhfvrTYDS9oIwT0WK
IRX+Ezc0BeLx76jtr22MmG+h8F0DP8xXA7fAeHlWu0Dhw/+d0HbULT2pvF6B
6QXamePIsmFzyRSPeteaYYykQ3Dn3tAvE6QTZTeuZocLyWGt8WLlXfPnivdI
wHAOcXxnnQzz8Bt11eZi8w/KRCJdKlcCC4H33VmTE/qQB3tOokieO7tcmz+o
tXBC1KzqTvjnnEdhrGCq0AYJs7q6RJXxSkdRzugM2ugJKrh1+gLX6m1VCTrw
yCt2WU6DXgNWNVCnL2vJ7LzYY+sU5yh7A2hWTxqDnyNp8q4a6PPopj7xXJs2
MyfjbAs1N+JnUuwg+ciuCSvPcS//xEM+8eJ8g4gV9D75CcIJAPXgehNoIMcU
YGUTn47GYGDhqBKWBNUOnA1BA0B0ETiqkqeDejoM2hc2BY6W1d/3YPujlVum
c7gN40ELL7fyVg3y6eswfH3Bwgusde3qFXsKHyypnxD5vFzWavY2F737ssKx
W72SadrmnI6YITGUm5wrN13gJEsnrncfVbjwonYoGGn1Ofv9CHilkVCTezxH
mceC55SdlkYoPokqlCohRdXUZ14edqntAtZqJnpBH9QGzoGV7lWA+sbyOOqz
RhYk5r7Mk8gkGjE5mvpAkQncJhf3+9BOrhk9y1qVyNoufOqaCeum9KFTmAEP
zTYzzoDnc9pSZMCECEEDv26cw7Uy/ZXipq0uHtRdbI5tq5BEeAG6T+wym6WW
6CpEIGRF2X+gbCxZFQ3t4e8OhFYkb7hp0m4maYVrckDxFXR+qobgXlF7DR7w
tspIRfUSpV9JYLTDnAo69ssVb0lfM+n1Kz2cY6szOxjaevq5aRn8ZKlzu1ep
oJhgZUaQHhL1DKRPJFe1JA1BE26fHR9/9/mOyjYcVTEgPM8qCF7y8FcsHetG
TagJA63mGBBFzfNuSBtCkzrHJyOlT6a7MgXRYcJgpA7fw03Or09gbK00NLSL
16MOJKGa4IckmMUy05a4UuxoOCaDslFQv/Q+gY+K/zKRsyANi9WXOcStXnul
FIy/dJe2+lmgWCvVdCikL31gOpHZF6P0QobPGxN2nhQZAZkkxmRmTbbTlibp
tbsW583UWtjOCA7LlAB+QYj6S73TeUPLaFbBOTY/wQW8CV3QOYrucRU6D1NF
3zhVq66Q/r/1sC1hf/Pd77mvTSTTrTdc/7ERiGbc4mu574zDxIbDr8KxY4FI
1GbTqAPFbXNgUjev5slz1Sg4rIHmX83MZ+UD83EWgxPjT5Kt8WaV8ZWHN4NC
S/6hr+QRv8/8nfd12vldK9GnFdR0LVFZhuiu5oVleYCskLPRudPmLdksN+51
Av8X3cuReZ0e0E/h6vng9CXzEfrwYI2+aYZa+/68lplqIXAqiePiEg0Wjw5C
0MDyuD2OJZR2QZT8yKM0SYIKDPHHViNPSqiWVCaY6Qv95ImaryOzyf2Nmkqq
+6HatUcTRuPMH2OxoolUlG5NFluRWE+KolEwUZRD5bLfTNz5nAWh/O9oZlEe
3iNEmq/3PX1FmCQKEyOPlWk56SVSPBsQfBbUU7dz7S/Vxa3PSYclgNkAUsDy
R0TptxtXekVpLBNi3D2YSC7ryDQWKbylp39apSuEF0G10sIfUj+EKWwoxrCY
Ld5u6vqikIaTZ6ZD2TEHTOe/IQoDBqDTmpkjWX3sxIfYo17lX7uL4M+TazrX
wdcctLvB4QgWaj0/bf5w2xHi9Dow7UJt5livzE2qbAHFVNkwLQ9fqRMaaD8Z
Ih4w7A42vZoif8hl3NZd7RhpGuJfre/Q1d2JcdYZnMOPfzAlU3ERgw8SUJct
D88EPWQTEHjE/JqXircr22LuTKqRb4PMFJyKKfN3QSD9SRXJogmpMpZ7xISO
zW4NYMDeU7wg/YEvlMNZZWOECbk+rQi3AvvKnXEMJSqkKZJ8Dshdynqy+kWM
9qavEK8TDKEppyL3hsiOEOg6kAxbYDjqLSr85KQR7wD9h9FdO1PTUBKmIP5y
CNqV1cVBoKJiwhZy8YPrwGxusahrUHyEwrxOJ6wETLPcCm0Kle7Pvtrkw4qS
kLVn8b5DovzofYIP9peTB4nA3LoNvhRzXM1MZnjsnbnu1rutjQuO/XRXJNeu
jY2KhrvCUnPxMirvHfX92kHYBjbm0iQAFdyV/j597kD6a69UyBoosJuAj3k6
ICmLImIx8t9uK8DcdHMcoKD/Jpy9EmX3s54kXNUTD7wRDpbl3bkQk6N14Vn6
eG2RTN6fZQJbrZ1OYHvwDn3dmaoP/K+Y28qwg6WlIgQtczdpsMelBJTOOAoy
KaUzL7M74jD6tnpmfw+ZkmRHdeqo3qGHUCRj+F3f7OoM1IfRNiuZOQll572b
3A9MjwoGtzMw8YnaNWNXywY5qG/IfvxuWIae2JXgSxc8+4MQF9NbrbG9utzq
atj6wbZQlt9yoxVIc30ZvymoGEEw2t1zYFEppqSJU+hqumDI0r+9gIcYn6B7
rgC0NuqwWcR3GwuhjzaW5Q2sSWxXs9Da7ts4CTf+HpEx7vR+LB6O4GZT8SPb
gVdN56CbXX5CTrZIHiZbuiRpMj7KmKCdzbXnbJfirLR6wAvkBz4pShDaBWo3
zvNA5hijph8PvHtJfIrgDQ5kVPG8IG8HBGI03W1dDxQL9jHXb+8B/2SnfRDW
GFURhO47/lO8o7VMy2SIB3gXnM5YZYtzMKKeBr0udMbMRWPjhqUPUBoSAK7F
IbkqX2cxh9ZDk+p7++XtNnL3wbaCWz9miBLMCR5kc1wdkrgkulHTY7b1mvNS
bk6+NVH9ovwGb1AvnJZssE2x1UtOZm/n/4O5TVIdpLiihqyhY9h/zAZJORLL
pNp6ZqpJOohBoEv2cRF8OD59tyKHJiYlErHS+QghGOFuIprEPx/AS57PkThE
mklaYO/WS5Ep7xVluLA+AfysCTZnuFbE04I2FDCYbFu2qIIXGCsJhU9ObP+c
D14gGOkAG9ZnVOHtoaUf0tr/71K6yuEjeK7B/t2tyXJiNyuftlqBBHTzPCc2
GkzfC51guyrOgOrHsKSBk/pe9gjWadIseWznhiAHtwuxeFGOiBX1idK4aNsB
G+p7lzEuGzj1JuwPzI+SGZLQb8F6OLcp3uGtr80I/gDtpo1MnkdOnDwWV+fy
I4Jf+C0nRe+HppEUMnRCj4aaZR3lR5C1Bgb1zxA5ZWg0MiowhvzKyH/Hh5KG
KluTlAa+k+Rk27bW2G2Gw3qwB+IoS9dGkM9KVLqdVCO/SmF9ivyt/U9/u7Ue
UXD9farewoYG9z4U/8B+zyWKQ1ouCIhbRdSedeE+FRx45B07sh9kju4LyNNx
SU+Qcqq7ILrudTCvdw8FHtg6KX6O3icuzUkVDR/R+d5+mRyCdMDk2H+rzwKe
JD8AxpMxkLUDBsulkOu3UB9E1MiOgkwjz16JN9IUYCSX5jvs2sOQnjVIrwVC
9pQTh07a2PRiZaBQObBo2pCmVpqK3UId9vk06PlAHGbKSpE0q0KLJJXEW1dq
UMLYGBP/+Rvzj2/YBvUVAl/MFDII8m9qbQPt6G6LyMbKcfoyiSnaDDMhyW6m
X5rfaVqg2j8cpAABsDztK7RLRyxJGK7SVDzF6z3SPzmNITKq1lkUzhK+D1jI
cowexrKYE2qLzkcdldGS0xOG9gg3XflyLJADsUNPkbNiywer4BvbXI/Nx8El
/3+X6pNmNFakYVBzrLaC2YcXRDAbxDhZnHUI7kiRbOkdHAiqCX0oPqnhdgQ5
la+iJnnQe+O/qQq1AyZ3its/DuXhUllukVxmhmVtlqGCFT5cS7FHJh+GVM2o
02h0Q9g9C/IyGFu9oAH7Fn+4FkZM2ppMKaQyOdw4ZWW6tUEy8AOxnjFCvTp0
s2SNVTt5Qf5a9E0NiH1pxKprIX6QeA/DxuCQkYeyaKO1OzZjDu9mC/bEW0d5
/wd+OnPsKNN7JKexUUu9NoNNwg+9tgdbiAEsT/oJ+ghxnrnWeqTIHnm3idUc
nPlqLbdY1CmM70NnMwl1O4tszUSa4CaEk+6bTphpN8UJahOmniRrnyAn1qAP
YAt61d4z1AnWIWX/bUUZMBlreIzIfi92pj5CpRbvl6U8pt5R/GwW1op4Uddb
vsUQn3Y/+rfFslYXka7DdMJVOOieNACahqB9VS2XQdXcGAAEJBKZnKZOPiab
yDM0JRFgPRGk3ZccEUkfnT7+OtLW23t9vtw9LIg/mbgbVCDs+VjK9+h+0ubX
H6gIQBD/b0zeoCj5kDW3pyC8EiImDoUeaGQy+TsGlWWMRiJgTOp7P4lqkHiA
2wVZedAISrYb9vpPUDtS/kgayLhh5z5l8wPbHbCvOB7Mfl+j0jbUM3eTKLUC
PjvvEFAPC4DG8/apB+lcitFnM4ek/lRbQiHQox+A8R9GJB6wXSq76zSfhJek
+R2FXjZirM6MWfhAFUjceSDGPrpg1IYvVKs2Q+5C7JxSVPX0kp5cD/maSQz7
ZVlDLStkedgtyBIr4m54JF6tysbboLlfcDsv02ngoG0nlwz8oCa1Z8FaATEz
J5Kx3PFITKdttRKANnlWnNcOQDqlMYeBS19s1WJhB7IHmOueIuA94aU192ZE
0topnD+SDlN/puSm4QiuuoZ06U5eMt6ZtSXKN0I6wVC8puSHBXsxsgs6KByT
sk2BxTgm+zLVhPLg/a2fCByb/37TYfM34wRitI6D7XPd5UUVSMRxmhbPX7rJ
fkC513bHQ81ILoOtW+P39AQ5avS3IFRgRazllOTfE0HXCuhXAi/8t3bv5kLu
u8tgg8XGmxcUH0QeTl5dxtBeMUDRJtpFIV+7/Oov34vR40O7tlgG4ra3CdCe
NGH42X08UX8rOFdqCR1S3dnvgVtwyaKJysUPpHdPRbagNrZhm6UbmUZgqZac
/rlKmZpMNP4/KrnAuL+wOFv7VL3jHBcYOR+D/Ixr6xXlyuU/eoVOsc+pTbuh
SVvD52VX0Y3VK2nHpaXnlaSjL9SdQHu5nttX2HiEQV6WQfpiyt1n8Z0EKtu0
janfu9EXTWzUas0OKdaAmIjtYGXS9n6zVgpnhrc7o4FHTXXIoECS0scDKUKO
J1zPW0tSEuEDp6gyQG1UDoA6elsukI8qKTgGwhEmt2VvAGt+EfKcyhLvp7GJ
xzKXr1ed2i4TEWrjSPi8NjeFmBohffq43yQHNN2Az1Zxyqd8Py1j2GuUHLzE
n5K8OUjHH16zMRWWPk4xKNRAuXBpZJOq4YHTV24Mj1KEEfYryeo1stz99OCW
mdqoYQqXcNBFbZ+bCOQOev02K+YBoMTEl3TwlOwgLG1JqzFo3AnGBpZq3gIj
STHYcT8XQ5R2rre8S20G+uSy5e8p4SEvyjzZMcKWfLEc0dc4NNgHE055zVQu
CDKkGtJhIVilGsUjJPPES9O/4utxfe7RaFYAHgNIguBsta7GKgo8pDIT8L/t
qtMZyi7rCYz3merYBv8VlEizayVU/6GexazdVC6Puqi4HRYmAxYkJ5TMRxPK
L5ubRzuDCvkRT0pfZ+NYFq8kOGg+Wxj6dNLxIDCrHD8srRRKWV+K9B619ZI+
KXONANIelTxXIVbkKFnq2vq1ofbhob86Nw7uJeJnX160uJuKNO5914DlPrnE
cv1rHnrAaI+X27aeU7TngLmow0IvT+7lVPTDwREUqGYY/eqYgj4TbqvJXek0
r6Ff9W2ISU+84oHG/u1QQrw6QSDSF8Gf0Sz90eS6+kHtnzd4q4NCrSqp81qG
M9QW/EMIU5JiNMVgl5XD5yyWBn8FkVGJpU0JSBP2KA9VnWvE/PsnJu4ynuRP
a46d1LhGJNB0XpU7acgV6dG8YO2Q5AWLmzf/Hx4Fyf9yU/qeRCrcORr14uLY
/qZ2Ibxb/DhYc7LGGbplrSqoORgBxl/zJd2pKNJJE0HxzagCXmhO7nFii5Pg
gExWBKBy99Acun7a5VtAfLJ0fWga1K5Q/IFwBK578S1bJeAo8BucL4OTKM4u
qhJnu3+YPzQVU/kxTVSBLCgpOoJRfAfKkoZfqmze4s2jbS5B5MEqnP+vN0BJ
kadzD8IynqN+k/6sfjESIC2Cuz1zQjsi4uWlBgRQaQQh1MQZQWvZsPe/bKDs
vGS+3attM7+PfIn32ppjVT07VocVdRuaf6oI6YP7xIBscsTkE0IaXSllA2OS
bHtVG9am+j2PG3KNy1A+JjxRzqDU0fNvF9Bqt7vTMVBRl5pmVY94Wg0eIWkn
vzBnvXL4hjtHhrssKUEi/wbfx11giWATF3GjVTFif8lMzYBM/LEYzXLmUSiF
AGnh/gXmJRtepqgzZ5AHyEX0Rk8jea+Z2oPriCHSDIOralOuInIk1zkPfHgB
KxJa2MdTOq69G9KhKIFbJnKGu8aIutg1avKJFrJ5O6npMPSfYAFv3mydCnff
V2F0R434NO++IYNuOhyxSjZ1K1GtF/K2omP8ID6ZGAl1JkYNrwJNUEGaFjsf
SLkEYpWWVfQINLxZo01duiurZvhMePRA3NOyD9vm93luPIGgBC3+7HfABgO8
Jr4/SsdL7oxuMejtqVRqaxSb35Z00L3bSXqtwUtcBZx9dRS7QIewMap5snXh
sDrvIZOStGmfyFtTpWNfPtlWbiQ0GnK6EkTCHGqUd22tS9Trp+FodmGa1qLV
8a1DByoWoMwdZOXnNoWkwH7nNxG9cshSEZe8oCuWKipENxhrBlPhxobe7iu9
LXkyv6iPnLo5iYW+SfsgaRqk5RZiOPDToEx0Kh7wsElamebaZ20SOG2YrOhJ
roCqJSqU9h6FzqVi7WjQOFFkNPLwrx3rgsR2CQdYTjXgY5ohUJH7D+QwlbE5
T1djUwP03EZEDCa7MVcaVtqnKM8QHlo2zo6Qll65v+xMSW8m64CXC9b1fYT2
cihTdgh82xcFG/oaFiXORj/lIgxBz3dUK7KAKDuQLdLtLZUVvI3BsFcPKTAC
lsw7blH1WNCUiKrUE3ZyaKeoLiDcyxf+0HiS6rmJ6NCA+OlZaTozX9IcDoo6
5Hbgv1rJ42BP/k962z29dcQa89kRqyJVqMqS19jN7sviJHQt6Kw5OdHikZE3
3sCcDjYjIwS0HrkZLeRiBMgD+mPNZ6esrFEsDnsDlZ8luKwJAhKkeEGaK/R9
9XAZ3kf+9Gpp8uSM+gru8mWITDJGcuacdHr28/GKgX6ug+DKF+4urmnEVAwP
/mj++NuDUGY/+opowVvbanQdMhRSTLWHFBcScckF9cIymZlgLoLlAC2YZspj
9WbUhqwESem3Gsf5G+GPt1X755m0tyom1S9BTxIeiDEYXJxrqWSuCiCVAP2u
avdjxgwovneNtAAU4JPZ5TYAMiMytCmtCNimv16PdyUJ+V5WvgPhT0GjVUBU
UIsVR3cPytaQrntlouPF+N/n6W3QIjf+uYj77se6VJ7NxvLZBOAnaGYOc6je
uSyP7b1DcnCD89GXCrsui8qRQC2uFrlRJxg+8WCup65Oc7cfWzC9krhOS0um
/jcXwJjcBhzLVUHoGF7Jh9uEw2HkaPyUgKLqqrELnSF/UHvloKLuzK+JIPvL
jStK0XAiKpbELsgylal1+2ooEyrkl1jo+tzdxuvGxHkP2jviQtFP3mmiT3Mp
Z07C7RQFyeFmpDhc2uyvFFjbN1KkyxxSEpuX0oEMNYTqTwUKk+qlpx83NLS6
9k4QEODb1qwzo3dwY4c39H2h12zsdgHypdcAFlGJ/uhUHiwzRxSYZoaweJwp
5UAmHnpTUXEBWlZtDQtNBhos2DiZbHYhao9rhWVfLk6ohMfhEpZ4ZC+9INLw
1f6tDG7I0yUVuKCJKC3XZv7/LqyucuNXh1lz00jXhNcDgq7GzhbHOZv2DsXo
CEUiwbtx5hHT4k9rlz5b4wthOBOhkymnXGE7GmXYA8dlbmGPZ+vjPwDMuRcu
yngr7HgzeIbjf9CGI4jHDkwqKTToVtFIL3uanPDhb778FWsAyvwbeFzzbRUm
yQEU2HeO0PEL0lbmBNlldb+5b1IiOIrdPpczyL17u7R1qtWfxHUGa3Gp+UFV
iyjFiJVxRMolmSiQl9JkDUNJjXZOPoug4tc9yFhK+LFaYf4IN75U5hORXeiB
JbC9Q9hK1Kty7IFw0/zniElGTpntaaXdMBRUiY8K6o06lyHvVYpbuZCJlf2/
lhowMll7y1LeVlaHyRXdAJLzP5FesIrLEYMCwtPloUxcz6Stc4y+bktZBlVe
p5ubRP8PhgIVRJwsuX+7nRoswMm04BtpfuDFdx70rRqgBdhyXcHIeKSpT6+A
Ix2O83nS5nMMyiPy6/mVciOLpRkoHbX6Lmgz/dA15dIG06BE6TZE5wbnu1oj
nxlEsCs1LRhsceEH0tsEfbCqQTTi+ldH5PpClBO9hLsOLs7v3dCRKdfDQzNb
K1PxDQBu2+aUX0ViGd0LYhfI8Qc0TuhI6BxHuMgvH1y7zADwiGLUJR3uYyaT
UJIXZ/fptPTNckjZnT23OSj0Tcda8OY1HoC16uoQ/yxXCITXqBVGcif/syqT
HhplEzwA6UDYdAq1/jTVnRu70EtVvg6oAdtPQC5vMmQsIXOUARUzeH+l8HNp
eD9/iPZuYKrfYnJbL6Ez5QAAz7RF2Gbs4ksZaDx9REj8WvNRM/L8eVhxBmVG
7E4IayI0T4c5tFClPkyQuus5S1VsrF9js8gpBmXBMgUgdkTTIuxzu35XoXx5
SHxNa2ZUVAPFavU6DRCLUK/KIPZ2IHWvgH5DmWpLtBNcEdJEsCSjMFVjyckV
KL/LejvuWxcrJSfgEQpes7iXIKsr8nYdimDqFest836I+3yvdc81U7cM/QBU
Ul0TSyS/PYRr0GszoZ3yCFo7Lre59K1KQEzhdSoMXmB4nb7nGUyUUrhcOVLw
urG3dwtHF7g6FnakN9+vYrk6pku9jX4Dw4cue+CsC8PQuq6wllYLUfoSXXTa
dDLQ4QEWFr/gKmUG1gb52LKQnkALPZO7qfhHFZmOe++CtjRFJ+/3vMGxV4bH
ARNxl9DyCxQoGxyhcW2qr/hWom4z0tATaw2ThaQb8hNjpzawQOdLQNmrVqan
RRHv/zGPxnekN/gBnM9HbLIvdjB1XiAAJrK/Lc38LMbe61VKbt6zq+T7Yqmh
1iDpcTk/b2UdXc+VtuRV4KyOdzDBqbEqwmRi+5jPLIpPJSyZwyRltWXABsvU
eJBDkd2xAP/qsd4CIpT5opdTOV9L3fa+QZpjZKXOMIKrtee8Khj2tsb79BD2
FtDAF4yIzmbru4QoZOd0w1DYHamnxhoKcByzCVGHtcLVvAQywrVnxtN5Wcf/
y5mKtvd/tV1iXBAkJEBnZwMvP+kEKNX8Wqun1es9tF3fmGWVRzAGXRLzVXrs
SBkfS9SR+JOT8d06K4Uo0jByYv8Dl7uxZA34qH0CsaE9XM4ZnzJWq7Clw6m5
CYCTQISUtA0iHYqCnJ/4IyS/qEhcBbbwhO7tS3ukVI2F0FLc58fEsfXDSUuu
LePgeqIh2G3eKcNLlTQMxmyI5G64jEl9zMQKW8B/UYLFtukUL70ALPyTW42L
7wMvno8PJyY8DLRWeoX87mEa+DUWEgiS92R7hfvkBaeewTLFKVrcJub4DSDo
6RJpuWUtQsELajQXlL3u+nZFcLu6m70/ryi70ImgTvoAB0v3nP7bcmNrOL7l
pc/uTJTetWGalXoWzW7GTgGpk5ncuTQAmonC/wDA125jNUsAYaf6A+QLnUle
+Z7EL25eixEJf9H3ABN9j/mD0P8/ezbsGpYK7/x+HjOhUgpfzmJEOzGLXT4p
w+m1oDbAI6JyRzbQjfcTWKljxqglw7uc0FMmXmlb6iO+NZ95ySsL9+SDaRZ4
dfA4/NdWLLCixCnURlCi0JNCbb6Bk9KSfbyuJFk71FA45LaYnjjFwbJJ9QQO
2XqAWbcWMn9MLlPFol/QY/oh+NMP7q02Z0mDE7Vb6M2zDQuQDo/cjDZXA+b6
w/Pi0HEZAIAM2pKio+LTSi6IQVfu+aStcFN6Wi88iQvppJvUz9ek6TCUNSTV
9WIvIJtBU89PvyfiyzjuSYh9O6W6zchGG0u3iZdF8jDFyBM0Dv7/5iAvz5Ci
gl2ddftGZ8McaCGtm0tMsFJVwxbVYIEfCJMvner1o2U5Df7KGdhZw4EfCXWD
/vwsgev6ucpaIs6yLYp6SIlJLwPhRCLKlIo1hxbk9hawAtDH0JjrdDDflXBh
mp9JLO/gwGGhIjcUPjlY0AYXEM0RLY/A2Hy9MKf21wg93hh6jd5H74llaqVs
E9QXHqSehqjb5MuY4IGveG6rCHmbgjPhiwDp2RjtbYRk05Ad1cgUdsDj5Tk0
0S3Vu4hd3W0meUsvMk2oY5enZlTauSi7RNhm5FV1sDyUx0ZhYuFx7J8esKxe
XCY18FeITnepCPgz9wXj/WrMO5LU9vEqQEANa4s2QYFB6DyHiaVA5LJLx/JB
GBWB4ctxkHvaOa1AeVoaWGXPY4mnQjii62gyoclyRFfYVSjuhhw2zt3dR3R9
/3t6H79NEjCdAzhyFHaCXRS9MA8Pk7zBYP3x7atY+qvPaGv3GdlAyvUP+c20
u1v+0xR9ZmZ/bXX+cf1VOMBlQPQYO5DX72aas7tx9Qn3TedJipGM8mbjEg+m
92MsaxQLNwK/F15LyP7ZdKna9UJ2N426Qdto734aBTjEgAr6/RNlHy9korpm
zYjuSCRXyABC9KEWSQK89BnDOhzkU/yAlooJllmfN8SEWOVszgbYZ9PAFZtj
Qliyf6MPIKo8qiauYiVqAomSbZ3DmCRa9b5M59UXYNbXz3+dpexK2zbHhT7q
WgP6SL6VxO+E63mfT43uSiTJZ031mJ4+45dRiHf6ReqI6Wewd4dOixyafZKc
gBo3G34o73E9UeXaqGmP2H0pKq43cyu3U6qsVkArMQWvgT4UJEla6LGYw90M
N9obOWI+frFIdzENssjsh1oYFsMgHzxLid7u49F+FLmp1mp6V/tdipFfbin4
h7DLMgA/bLcnCVWM6o1N3jgmWCOtW5FK6W7dL7ha/ZGgTrvyq04qJSdz8KXd
qvAFP6Grn72rH8aZbqzekLeXUHX9eIUBk1ca9yB6MmhEfMKPnlMMzg+umxeX
aJh3t7jsGgQkCI4ycXiOLcgPNsyd350uMwEV/KmomtDqn821ba990bwGf/U8
oSZgyovanGLl7VFAzRW03cV4ygbG3MqdVtsHwPXOSiBV398TGayDuPfczlFc
2bIHG/RocMzfPsnmXPsoSk+TC8pmvFUjm5gFnGxOaiJ/L5aUzBBkCHWrey5E
A5AMz6RnHQjrR8U/6eg6+5fRKFY67UDrx3gFeDdFqUNnLOHy5TBSyGwWsCGg
wPDxr42SzmXXh16Zlabp48ygSVb6+FyLVDFz7ZrZJ4HQxIbUPdTuKSTHVa43
yxTt2wImW7Hd+6DQBuFVn5+ZGV8pgxouULMhUykeo9rTS0kP1MWkexGHS1HF
qmNwX5HDsLseygxYJZkQhDsh1grWoarSMhAKmVatnL2ufspEcnX4Xxp6JZRM
28lyuhWdnsKhIMqx9HqvLa0f54k2/P18A7yOklVw6xf4aM22nXRNawUUbB/g
T80Efx/xd6CDPbDppI1l1aBogE+3zz4ws46pS79iVtP2gHKVZt5+WzpuuRwB
t0NV/k6FGBC0BnRKXig3THg0tbCw4PupOrOP1FFLY+6NW1Ei6U5t2k/gabW5
rIK4IRj/l61lfqB4Prjn2nNmG2dj3uz474kiRKDXgroNPGgvZaSUVQ8ed3Jf
w6QN/yYjOdkvwTH2VRO0FZb9tZ3LUQETz0BfEEfx5JbSueqa/Hx+HAL0a2A4
Y01n/3NL+0sHp1Y3HdlXvtL4ho2iZWu+i/LjgOeQ3oJKwUXQuwyDVUO6MViw
2tD9+mt520JCJ2TwzN6aoMnZRoUSQjgSXn35aFqckLq+ikd47RdAVn4KKhgH
Pj29TtEJQofODDIbwsubjkp5hXvAvEhUOczmjqBRgvH77xRtwyfaocxgzcRS
DNv5gcUNiWD4ts17D1Lpl8R/COn9kPpa8mw4Up6YVH5kLmE30n7kZgwenwSw
3LDXPGQlBROYyaNIqbycYPqhKr/tHxcKy9qOCBdaNkO+rvWqHtdqfUPc3hWK
+3hQDFXq9tgVfzpa3ApsU7xFjtM8Bqra7NnOnPbmJhh38OTMoBR3hDRbUmji
jxD4jBb+Fcg8hkCLju7wx8IjSCKORd3RaN2j6h3UE8btin0oOpl0QZGSBi+S
wqY15PbNlWeicySJ5sERJISmCQCfWHG+xGw2XbomA29lXoMSNnPPzAlPLpj5
iq3q6mxe1YFqLQ3zj/5CmRpvgXisjx934J33PWU/feH/rPJl0J4bG+WgRxZN
ozgNsQu7fVWKwtS23z8sA+ueIzuGopTv4AvlnvcYVK0TuBvKH8eex0OHjDyd
r5828ZiU+z8YfLvk8kuEAzPj7xC/kvzLMPgM12vPIEHjUmtO8KEuDTC+VSA6
mfQEdlT7Tc2kTQrwgW8jHeFCw2mos2r+Sn5zjizVQ9h8snCHQ30fYg8XKfN0
vE3qQkPuIuxtL6SFvpyPTeXqEfyZx/3mAeozt8SMnampX8Vxffl5sO9hjeTl
qJqY1VX5gaQ2QhuUcjhX1Xp/LDHmGcquUOgIrraN1kjsE/o3+ioDqFBT03kX
+U1W39aXkJ5naiza3C5iL6epVFAe3rPidAodO+TTAk0AxXm/05G4fZxeDUVc
koRhmSn4Epn4dOy+uVcCXr1E1VvnjQLRvOtC2wXIar4hZRhOytLfKzBOl0Df
d7KzQSicq+B6FMc+4AKh5nDpeMxiPu8rls2k8u/eTzznovo1w2IKjfd83T7E
8QvODYCHCvnrsmskT77EotucG+igsHE0sUyTstT5UZhBOA5u2iekAJUCm8+W
Ga0NOeYfNNMnu7dvWppVTBDUhkULb3iR4p4oW0HRCn5dzjW1ctjoW6AY5NlP
8OYbr81H3Y8NVaQj11PtDXir+X86sLO3qjoDjXSXSOt0B1f9wNSKQCn+JO7+
0SdtiJbljDqLFCKiv07XuiUUVz4jztKb5wjkC3XtncV3cpsgBK+19qUuzhPN
uTI1sqed5cJ41IJWV4wZGe1C8psw/Pwyy8UzTY6NtKdmN7b1rVtC8bz0MX1n
psRzp1JcfpkPqSkmQKAipjbtaCC0jMboHSTkgzlI3jwmI1MpIdpclCekmv9o
kBeLINU+phe3Lv30GQ01VgOC1oMNrPCtYlkSbWG6OOVrLQhtrN66rJ73T9nq
v9KPxkI5H/3pCbI8ben4twWr7OZwxng9HlWGPsgx+jwkSa9t9uviN0c68RMS
XdiAXcHCJaaihe/aJPaxftasEJYty3z01Sri0/va3fVi2TFZnU4zbSYm9yQR
9QwczfGzSeY2OJ0lAD/SYPar0Bp0WjGlUaBEhAXA2QSjWptgFWhSBhU2hRRa
YMYXBfXDrd6OLaZN2k3BPy/5CSdM9CvuFoBH+pubvJ0yjfmvYcuMEC4XkMmr
wonKTQd/TVCe+incj+kVafw2juvJse5O9JFbklvR/QBvxcUngJDb8XVS8z8l
z6DqwFx8FlAIjyBP2c2oQnjCBskIhvIeS8O7AX7sRImEwL7ZebSBkUxWugE9
tLChMHt6IeC7F6kPsJyoTy1qF4oD7ltuPvH1NnE0y8nwIqixEPCpP/uU7dWC
MIVvF/O1txyTGYHFveB2fD5gTbDYTtlXToiUn4zxXQkIfIPSi9U5myd0w/Zh
sQJNrO0lR1HYfuBDI7UxsbqGal2TdkCifvy5Cmb7w/41OnoXYwGmdKjvmwBw
AEMgNe+gJ4APfVqrwTVPA7+Dbp2kbzXZ2mVFfkRvv2sTGgXnusm+FvR0Z5tr
jjqb3OjAF6jafXPrsCueJU2oOdIihmxirJdw7VxWHHs/DueK7WK+Fu/tQQJA
xXoPhmlc0hO5KYaV+2G8Cnnst+JXMMO9iBwvzkI/f3/XkUkHf8bk9nh/BFTm
7SzOcO601FTDKsfzGojpVh5WCXcErFI8Jr4A/y6NZeJVO8S0/H8TKmEIkq3N
Cj3/EnGgdBKUedt57w9F5KfJyAE70wR4hXWrM/xQSuxP5X1dPhZY2Z5Nfl3Z
1igjC20DNaqgMVOiaKT1jyt37pz/hM90vq/jtC1rSmCrjGXAQP1K7wVHifH5
LXJjCD3mcQG0tczs2nyE/WReuhaKQYXNnQ04tt4GO4fQ4h4wm4u14sYBLE2a
8kn1XAyO1Bn/8RKeE33xey7Ez0Oc+kZFdJY48p/P4uC+KOGO0NJy/LfzvJnI
Ocxv5kWJhng8PgxEurq0rBsmkapLfzQ2AEvp5eHiNNi48cdTFBc3rhlFXdr3
1LHQtyVYQ5crTNRFXLPDzcAsw6VPoEXxfI4FfE0W+Hh3Y8FDmyE1sVmRrPTZ
ubgF/W0ykQKtVF8ong79+PXgGX7Td0V9orpGCqH2jeuIVhhL8lYmrpdDGIeQ
3xHb25dNyYJTNWhomS2WyzypRA4I/zsTwqhnBRifnbZHp4ADxsR1d1Cy0+UF
6rfWsDzl/fFyDTFuzdfC0PnNUrgCRA0bIp3cOInWL3vrI1yeemWppqAD60AY
WsbQo5/JH+SXf1NbKP6ujtvl55ppQvCZUZ6TpipoSqmT/m2wq9JyNR6plvsp
rffnUdiEvXF+z8atLfBfwa1DkmtWZjW8IIjTpK/i+zbX9OF1RAg61WtDi3Yt
QwzRe6TSnHxeumj6K4jYQziebobOXPLvJFTYQnf+QNxmNeVyEkkfmWLzkyWC
a29oys9wDpBdr6RppMHtxGWOA2BjBaLPxv+n4Yr3RFUbo1T0Rp2qt+0mu+Pc
/PnsTikoCf6RiDPCRViIlcY+UlgXbXMqzxagpUfF5X9YbIpJY3Sy8EcKO4nM
fMHR2JS+kxzzwk8jc0DTGt/Fi9XNA8gf36nryND7wZezJ6/f4TJdbDKhiKGg
gBSxNQ7kyySHjNWpuAyct+ZRt+FlucC8nDDCWOAvj0VCjOEjndTeZzOc+70/
9uFHRcaRdMEWVIUfLOvohs1GGioi2y9iqufJs7vLYddM1dYCi4M7xirFB/bU
vurguQn0oZC2vHtfrYa17NCjcs84zzYAuT7zy6U7+lWvCbjvNftyPW/uOkQg
QEvFiUYQ0Wd5ztilafeFRjqBWxmoODuIAa7slGOiExPCTEekOPvMafIRqzjP
xDbdLSV3cLBiE4Z2n77bLgR5YUEW9ABWfGCAlmyOQt5QYJ0DGGwKTxbUwVgB
Xx+Ylnajvs5qCHUFnghQMvvMHH9lFNyuriLbQ7Az3nJEPvg7jabQi6BZjA09
q9WeqwTS0kZxx+5d+3sTaoDw9GvO9W8qn/EyeHllhG7avhwLmO3MwMFcy7aH
eXyJn2XOPsHstvciWt60Zhil72Y4mkotoyhL/bC1pT2Px14LXLWZD2ZgPSj8
I6RlWMQUM828kLrcXZzM3TBhyClC72ONXOIt2WPkQy38suu7FuhVqsO+TDDW
raeijWf+DwfZz9jldJYBHYWEqEOjGbfKsn/3lbS0eky4pKA30nkmkPm0cVuZ
bIfozyL47LV2rhWLrbb8JfNHPNQPM7FJdm4jT+TrYllKMs3kPmVbr0IDMCOt
4nyCePmwnLGE7/75N3zC+v4Xwsr4ol2pk6WMNY5VSn+dTCMWoIGK3plb+SQJ
Wddups27lf/iBc4fxXRtO4leXQi8XjcF9ayzx1Z+fyjgJrl48DcH2Sq5fBLI
awODn2IfT0uKUBw9xRdM1ltJZ2wNrv5P8aVvf+GxRAinXhVRt6NAxFXu+gV+
st2T5rziLgkEu7xkwKh2feW/Az7xne1HMrVX5XkopG81qYmNgP9RnonofvaU
8MOEFHTzBqMXVeZoxBy4tinOwSO7kMRnmRifRXFC0EtAym8h7LaVf5g1M0ut
iESbG9RKwmsDD5s3OkOy7NvLXfYtJY+sKA2ha1Lcxo+CfgEutSbSjIk7Zg41
0Pr+xL1hCtntHxuirBSsqx7Jjq8MMNRrSdyvkkw1ulw8y+iOIjtLLxvj01vh
vtjpP+Zt9zhPf3jDyt83byppZQypy2qKiRQbXkAYqLFuuMqNcxzJzevXSihP
Ln1JUFdYe8RvrhYsrFHHXns3vsLNsPYoZin3GjX2fyCfjEaa6u3DFMKUlm77
q4axDW2r7S3I2LtDz+vvuid2M4smYLQLlEGkRsd9ZI4Toi4u1blYpomp7qgv
XLFcAZu2aGL+c/YdfCXMbgOZOKkfPUKWnVZiNVqMgl9UC4S0NHU21eN6xuwv
S+Q5bxST9N6RKkUtrVN0bFt2zk9GIe1lQiNzbidvRTS9+DZyOfefVG9ugyXb
wR6O8BVkc8A7K6QjFECJ5y/TfLnGTHM0E/Dk7Fwf5hRfzfDGQN1PPL17GSUq
HwvwMivPLVPW9Wi31BnI9EYhZcIHeRAdU4gbZeymMXpwKuPTdLlWdTTzSqfo
5QQnhrNI6kZFRW/wIaqQA089DU2cBX3I6fnDb3WKBxQiUppUTR/GGlmqjFRB
Xc5Hua13emS1TVD8M35QvKYe9v0Gj0vzh8wOvIJPubD55pO8PADOvn8c64sb
fUjYcs+ed8MUMMr8Kdu0gwWKNAIDty8ZZzYq/GPnQAJBRTsdhaH2xLZo6FGn
o/tQkBKJg+uYISagKyXiVuXKC60J7ynN345+b/iFQf6lUvYHXfYEAz6BCuLV
mzeO7bRdvTiShTlQuaSw5NnM1Z7320y+edo9TXytZfAMh0Be14qrF6+rGCRR
mtT3/s1Fti/NdjBss+qrojJhA1Rd5YHAJW/z/JFiWkd7mBTR5uZDDWullHth
b87al9neOSaC+fFVqc38K/QDnCw/yJEf7YLWrmoMnf+qVPt6LVDBKog5JLC/
wCBBEa46uMcxuIf2OWAEaADuY+wJnX1IiIZrO0gn4MfiRsF2uI+BeGgj4LTR
QoOht7m9k2lxNtQ4pj6gRzSsENNPWPdyNxQ5h5vOvkdHheQLVTWttfX9fe5b
PBtWLyIlBaHldobI+4rucLpziWatV/S3uVYPXydJ/slX0nabKiQujv/Mgiic
1Sh6IbE9m0IgQzFhAsUqMdohI00J9SNs1QzgbUMCnh5tkwLcP2ThI5WpTiPm
1RPw9WYp4a85GTeKCYKLKBUUmsPGk5y/ES2F6vBRtrt7Itk4B103ZSqEdlLV
BfyqpNiwE8ipBdxjyZwXykHbEiN5I+6i99JsvLtHuz55/qadiwX2QhSje6zB
6Ca+6/Cl2AyDw/fO3HXKlHv3u8tw/kBb50VwCzAeOs2QSsLQ/CCdPdXYr3mX
UgTTYqg35NJtm2fREoYAful7gEdT0Qe8FkRuHE9btqK/IvPrVvLXnT8BJU7+
FfbyWnAKtcybeVn7Z0PcxGOHGdeNX6m950Fg0cmjwFGeFMmQCfsle9MGCVYj
I5bVMJWg8xkdFSMA6bUlu3g2BMkDC1/iDVnzGywRTZOylog4iSbpTFAN8eEN
FCetqQksLRNHJUpD/I+IKbAsBmCZiABmjh/P+zIklhHtFl6Yu4xd/NDSEwvQ
lVF4p5p6DoS3Vr/4dfstfSkS/svdlDvo8tqc29yhZBm1NU7tP8tWlY8deNDO
cPtAgNs+AafFmICk55P3UUdNI1sPdUbWpXLWDDdYLsJGo9kQFbaxnzQ5eSql
BBaJQe4938V3f3s4max63vnfGLQ+Bk21fPQNJrJ82njCUDWFqvu6T7McNl0l
Ol8TjZZJxdwo/7Yh7YNhigJZ6OfD2OhnhP6l/AZlCSjZEnHgHIHX8dnxeITA
ETvlME+V4HUkUO614sC3UXlaBwMm/Df7ZKF4HtYniXiHqnpN2L3ApnTXtS7A
YqXOQl24jfqV9KSDVNDl/Jl0QVqNUXlzRN+X7nD4KqUX3OTk59CcV6BOcH2w
oll5DhUhrFUlRW6SuagdO4kKroxM03AgnvlDwBxXcnv+umLllco2XcneKHj6
inzw1ukIILZLPwmQ9dRJZ0ylL9onQjV8yKDmFTsh/bevoG5yX5ofrwXYfEB1
Iza1HZcmjWi378li3rhhiZcyWHUbh7xfL/5rAyx4Kc/aVZIEM/FzvbM2FAf+
Qtk7F3G9hq02G2q2L6Qimy7GmvtjyFJYXMJCQ4IF7lq+IbV82rTyDzfNTOj0
oQACO2SglqHUN2N01spho92xxdVEIkh2gGjdAbchAOWtlT8WFe1H2HhZ+aiX
7kwiiYSdv6Rf2tAp0b4KEyV9UfQI6rERIiVDCubx/uQwOXe7x9fd31y5bg2z
SKRxUs5fZB1z0q3gz++Sls40nD/wZVeyaHuRJ/bpmiMFpoqUQ+NIYlDqpibk
kgIhBTDdevM8dx+wp36A08uDfetGE79uBX2v/3c4uESSqReNtcrc6ZCiS4je
LMnDqmrDBoynBpC0g0GczVsDUsCAgTNFJCyHM3Rl2v5JebGqosdkI0/toCWR
XZVqlhBlTAMLjaDqlFaztj5bIXYSv2ChSeWEZzxCbZWABxGGriiSLdTGtGUQ
0sQIugYFoOdE9NmBWRQtYAVtir/HjpXpPqYBVb0OpV+6a5CYiDT44/Gs2HQq
r+T+czfX/N+SGpxrl1s6f8+plnmzP9jIjDjOJhIjgatPzXSkeI7SC/vc6i/K
vdmQsRvhJZBcaWOWn2z42FuNxQh46AcByA4qRZedFQnVbLamwCGc2xe+8jSy
1SAKsCe/3P4KybeYwGDaiP/zaXon4zXsiNWPolH3UUCgBDWSKEytct/arrXx
OLZ5/+fUIgeLt2SRk8Az8avBrCAoAjti8P4F6cWeFkYLI61B/dgnI2j/wQ8F
wVpR13nHjpp76mwI/uaTTowrhSn/jIE4VR07NXkx0pQTuNi5yQikwl75RC7Q
LjJ01OKJ/BRDxqN+bIoKsWvmJnf1kcpyJAuoewn1bJ+xOh7h2EyroU1x6Nx2
rqFdUn9VX2elJzohPNKQVwF5Fx4P2MaARBetPwQ3xEYxlWxNM4IjxDod3U+Q
wJ+/zLolYpiyDzxx5KdiXj3GGAKi4XQ9Xd1Lw9+E3bocKCJoaz7dnkaH65gu
vQUN+JHB0HDiX3bxZzV+QBQI/XLngN81kAjw9HKdp9iyj4YecNkGLwnXK9Oa
76+bah7UIA8mkYVwaFmqlAnK5BDBj/bl5Asei9/uiClO84DOynKMxWuKGn8e
5WkoArIiPFuFbxyvVRD0TjZfeIgIfeZACl1evQD6JQaJtEsI9sSmuOOi14a4
TlU8rykG5lJ5EkukKPE8UMM9Tj7zpbjeo80tm1RPr8Zi7KSkU6iGDr49XmCm
p/B2Vcfpmt7oQBlGLgu44hT31JgUKGgQA++Hr9ij7zd8Fw/dmlbFQSbEsbcp
U0ugoC16tHVFN/5Ukc9VRS8fQdal2vswAOootDEn6RudBq58onD/Pq1MR9xf
F9p9Ltcp64RlVfW6IxlWOJWFel3bSmPfBZ6lQl+LCFtAypIoiFNx47yGRp1Q
9SLtcYc9OJW3uv8xhENZPU1hznKTfDKN2XVAiWOJU7NGB8kJyrmlQho4fAaS
cgxVnvzISNOaf/+fH6U2v0Fsdrk8xbYcJZk8JBjIXOWvEAZTUHzbkMW55waD
T9pVFEvR+lhdf2jGFjMxtXcLA/ZgzsLzPWULLdi/x0kBhrIcWtVd3VH1H6z0
SIlUf3CRjoh6ezpHwlqVTcJ8pLIKya+JXpc4u0eUJKeAfu08iGN8pIdoreJz
TvcNYuD7qbeyPmXG7He356RoD3O42PjuHa3wRnAnHhCN2llDdfjHejfIFL70
1wDWnvFbVd//bBleEaGtqCyrq/gfvtzTk4kI0JYnFaevnMQs9JQ3EBaWikQJ
6j7hnbPren7N05hruLKboDT+an0aaafQfrZi/mzMiSH+w2UopIDi8i0aPdXk
xko2L5s0lMETI2qRlO6UO4hzVAYfd+N1mvIW0mg9v6h/AMiH3nlKRrhcJllz
VZrX/3m9rAUT0ZOoC+mpVpUUQx/jw7Jj9Mwj0BThweJZaBJHD7nmDPS4wyYK
Kcz5NEA+P41lmnzokrTFMcJGo66x4QQu8XSLRijB2vuLhosA9e43hhCEaTec
FY0WCWKodSa4cAiPvGlHHLW+mVuehHv3dHDe9VBOsumZa4lKE59QFZHPlhfM
cwv58QWCxEpZgXKRh2reHb7K39pgn1VsR9a92AdXbiRQsr12uRfdghIbpvUh
e+dYKDazWytrBybeOOLPlBgxz+feW9z0W0iDKKIdsBAb3XfMDSEOP5h3ED9R
1eKPeUlTtiBaaoxPbWNRZaOuyjjcYS4J+pXoHwX0eYzfxHVWaW8OTBu9tfAQ
hZODrl/sYBbZTV+QUIOlRLT25v8PJ4VbC+J4P4Qif9WEBKtQG2QG/YrXA2TK
6PFu52BCM3M15QpnT2R1vVuNioY+8+EVosLw3HvqQ0tfs5v8uyPXfBlwXwq4
GdzLxBvtlBz1R9ryBTC4t7fh5FnvlAd/h0O6ZmCS8bhwTK0mCL14rY2416xh
T/892RHQE2TXGcY9yO3k9YNteO0jI216wOZgKMPvigzcmJLn95Xg/JSytZ1C
REwdRUywQlFuybIv7UX6XpHlb3GSR8XpcQ5GxNM44lGSLtoajurp5w+GwKLl
kn3LM4LbnRSvEg5DVDAYGy/nXYWucjqd/snM93hKvhET/yOQOzzv7k7wcbPe
PS1ITo9lC7qxraJxm6ksz+GqRd8ccVHXM5iy1n8Th1LL9CUdmNDBsKC7w9YH
a/dtlB/c3RytI/Qz5CTzesVh6iorAgifmKmVM3cFuid3yTCQS/ruJUmUp59R
DnYwCM+iHW350hssyR0V3PaS5kN+8ova8mJDV+u+2StFgZMczglMCYnscEci
SARpEdd+YpvbLRWGAQseblb8v3bogwE9Oac1phrsB/U6KsCxzT9lWwVLQN5W
+CiqklFHV07VmFyNBYqoroX24RQB7bJFgCNRbbe5pcM71qh1DEOVcImBaUt/
LIhJTh6rMhaV368ceelbz58vhEwNIB/EEITVbEsClZA1YbhHW8NQsAWm8WnK
6xrM6aohPlsOkRi+U1D0xQqqKH/TRD7AvVGEDoM9+DRqdcatdFHxOKTzWw4R
KD7mQNgXAJufVu2j3mtfs6PVRMHzytZwT2bDOs04S/i/EYNhqPClMDkPXyXy
zjyNR0uytCRAocAcsE6r4g51UG662ihGEOPlq0e/+aNbe1RoA1B4BY2tqPky
xUs1eq+vRapZhJg8eZrbkH3drySdkniLGXjNwdbqfMNHxQw6RiUYj4mwS46k
yt/O1olYANPlNNKmEaCDQ0i2jjIFwRerkulrpXA9clfYJd1DLxbaIkxp9as7
ynSsDItrcyNNsHuNfvMz8gPqC3PBsSmaT/NBZ+6kGdaRkELqtpKP3NpUS6qx
Dlo49vRDhLKKm4LNJlopgDaUO6lSNFY7SrtbTmZM9Nm1HY1/lmZgjx1Mhr4Z
ULlkXAYLUNCMD/CdpnH7V52ViVTtjomeurBcJNYB6tacoEQS4Qlpy+EaQZ0W
wQC+qpfAXmr8KrL58Ahsc7dm/8OP+FAecbsf6lGNiZssX0sSkKjzXeYQAg1X
6EAO1gR/ysUVVFiqd83EapdQLSA8OPXfuz4b9LFPMPsu8Rt/XL7OhhWZ3HX9
wJYcjfSdhwsH0PNtBoa65oXk9nKtKHOB7Z/Z0+leklkfjC32sLSXbu97Vlc3
V98JXNZdx5nj/v0psshplAnSio4fCTS5gK0dhr6XUSyBhgg/vdMheqoK3L0W
FAQXYMGIB4v3CdpVLfnGb93nhU4fFzjQZ13ezCe3BMCe6ROVtGoaDXbtqmTj
fkz0PQVNiS8kkY6TkLMv0d5VYfHVSEZTfhF4d5KX0Yd/xzKKeulI8Kq4CRjs
sxabOzg0UIYgIKz+ehltkSryfuwQQv+JtFTb13IDJIX7kp4gIayuv13TZ7pU
w6f1hgbCZeTVHNSlJOzIGiqmYxYL2EIeWCP5amTsD+d0hS6YvKDJ5aaj1FDK
fLkgvdhn0cyAAtw66meihnmHFlK4frzCc6F7B6gleyy1y5mou/WCujULxjJb
g4jJp440T8s12P+I1FoYKLeoy3pk69mE3xmKkxW1AQDLtcUbevkvIqnR/YTO
M0B77TcYNBOUpDpQgtrJbEPWb9NupceUAy1hARx2jbWcgToeF2v2AbvI2GeR
hE8oSrPU1gW26gZUpWew6MYYSDjuAfUyQNmIKZn//JnihFNU8/BWcuQPnlfG
GOd9r9AerQ4zk4p/RgsHLilFhRBPIo2Nw5PApbYJBZJTE5gCdHe7XR8zr5ii
ilt0HYaQevVavjPWMRRX9Yzr0lKnMVYlekcyLrtqUTnbiLHuwIc3eqBv/ltX
nZym0AlHLjdbUzBomR/2IAiCNeVyRl8tBpXKGksJmUZ5+7XSftSsMGe2FMXe
gtbqYT/krFKJsLJEk5WlYvaAOjlXUXrneOHXm2l7CrFIItJPiEPxFy/x29fD
M82UYzVdhX5gmn9WtUutJzvN6iBd0PF9oSd4jRUuDd4x2+02UZPFzz7eRHIj
ZZjX3W7aGEkNPpz3Yp/DYlZi5N0pttEQaboCSznuRSUo/fJGLmo5o25FmBK+
B8+RdfAuijU4a92QCS7mSE6IXX4oFss8sRJxvEzcNyzPW+bAM/bKyjt2wjeQ
j/g6PoPAJZGx1pL0i1mA4UljVYzRaf3oqCehQLkDCHuHmh7a0J3F87mCIihd
aoVuvsC4KZ7mJ6fPN5C1ycqP3YDJAXy97sTQY2/TnGXSnUvo+iunrrwie8WY
o/IvJFatkNop7/XfDdholRyIM/bmPXqlj5tDHJTMRZjJJ/s3+EgIZXdz1uMv
zFJI1mlD3dc8AwiE1CDtdoC7g7qrb2lzMKCkVOvkQ0wPH8vneRs5H+DTKPMr
tMEvR/m5j07JWQ7eXhXcRqVkqsu3lW4Mkze0NJZwxLv1TigOfAbQQTKpRrKo
/7bu/f0RWf4dqOBqp0Nkwr0EJ4rif03DK6IfMY92SOWSM1nqSmNmijf/ZrxT
wJCPg9J53N3/9KdJyPDnZ9o6XdgJfYjTRfbkfoJWXU+Gr+GWxs4YeWHOW1mC
CPTiRBzhdyJs8lOftBIpCggVmqVdMjCHjuII5pjp1kF+idDAqNJU0mGZrGnp
sDfKzTGLvlInS/NrjRUwGwpAydLIZAKGLe3xMOJQ+VghiTAI9pUvIHmnMY8a
WKLztzmmy5DPrdKUMPHHYDsXJMvxN7DwUEAHbSzQXwikoFZ3UDaidr/sjG/7
tDPUJEAEesP9EENWaeOIoJIieZ0J0RanbC0JkECxSinC1fbfMSNQsGbDsnpa
DooPK6smpBbDknNz5pE7owFeHqJt5WYejfUCatc2TC7tde3HC9mRSKXLq8j4
R01IAn4cnjrJsY7+2lZb+SdTSui4YU1O07IYNl2Sv5reoM+hiAwiFUN4BGs6
rb/pcNMJTliLGsvNNwvym2YAk/lSsBOkxX9wttSjC4j3KWLyt+eEd62RdB09
FsDYZgcK86KGTgxJ4Ce1TY41t5zOVIPtlYCYK276rXaDK8+D/kskdemE4jKv
N78wxBgse/e9n+AoCfdbk/z0ZOK9QrglIFooireE5L1nY5lNuCBebFtzbwzS
5ecdgbV9xyIM8ISsRZEDaz+1+N6usqcAUItvYIW0HeFT0e2bT9xTq+pTtuqP
c+Rc6RIZZnhMLB4Y7Wi10jIN2YO4lcqNb7L6NiRUzm0hvMJD7ZrB+12YjlJb
nGU7agh+r/RC/55kUEtDQT23MWARegsIaB+lgbKZTYYmV1rJTeWzzbGyZkms
5Lg9KD5pGzEbf6gFAdSGgaoCHcyHqXka1628aBxAfhY7iA1/K2+in8HvTGmZ
zyJiMP/Hsg9u+lKnYlflfCWn+yyug5oPekMm1HF3ClaxkDSpp7ileHpMB/9v
PURb1gP+f3i3T4cgmmZpaNaYkquEPwVpU+gAFpInPhWCnfc8RYdE+yQKXhA2
Xq/WRcl8ZQz0WIjXCgcNAkdE+MG3VRRiwcyHjHO0y5WNBmk6lOwN+N+PEYC6
eFTWzWt/RWFaXozOTPjucCN073NbbGybn9Oq/Dul76btYi+nxJ0aF8ougT0w
tZmO3bYaIgJ23qLZ62vkzfipai+IQ1iS08ZkvCzs+gzp8Yd/KmzYJwZTuEJG
N/bkf9lEwnyGQeeieRxhn/eJRSCQVXhc+cDvNMOmUE2JVEqYIhbPeUo4+MrS
bN5zGyUXlWgYqpgAJaxx1amkiS7oanN6/JT3YkaqA9Rn8jwsE9c2XvRO9S9Z
EJhqigZd9xQkq6v5lHsie4Y3VzC4FJEuAHyJSC6q66bottExwO8KljqR6vjP
2pYMw7Xf5p+7h4/WjdpvKkFzARGGx4cUtijeQYJfwsYrGM/hOr/Csm0P1DqW
mz9fmeVdUiFDWxVl/j3bTueaO4HNHXWsm7EePOGeehIPFoiOIsyrvfY0rAef
pQlk89oH6jYsFZpWtNHR+K5gDtCezoV+roEXjxwPVNcqc19e0Ol+36eC3nAD
RGVC05q7AmXbcbnQvstJ0ueLnEHxBn4ggbejdZBIOUYdBiojHZeDjNLjx2hk
UGgjKpjGbdClWxYtAmMOo2Y9bSXfc7hFQhgYmb4Ga5tXeJJhloWwNUMgiV1+
9sqBEO4ksHy0IAQ6y2Kh4fQ1My9oQpYauU8qmvFZv7+mqYX2ACxi3sCPloSg
ZDkUnLJ+Z02umfLZxFafWMtMOSvv/jD8qBtmV1Sy/cudr7HtrkRqnVshGRlJ
fHN6U2UzxhNnfyBVi+foS5vVnWo4cQGPh6jzloIOtkaM6V8FBBYQp8f+ih8O
wySHtcPf9wPqp1H55INUdv4Z6k154MaVRc8gSFY6tnc7jTH0TIUXR5KcVP1h
HsFNwCeCrleVsQjii2ETJ+VNNYzn9NNmf06gGp91ClMAWMH8VXFsI7LygoM1
h3lpzapBFZ6vZNbjgveHeLLSGQ0ZYmWCVMcD6S3yhjWdvfZvc3EGes1+kCx+
XrpaKsp0j3PmIi48LzUIeG3mr3UEgrpM+vb2WfoeKhyHslAaulGr5EgrUV6x
f/lsoTH3jjtl22y5MH5Jr/3i0APqgLPJPkCewU4Mxw8yum84RYz98s+QqKjL
fxIZOmm8X6TQ/haIKitcmRta5lkZ0biWm2XOTWe6cHwaRXX3p2cA0TGo+N32
eR+r7mKBakwyDNoYwrTH8C3l3OqZaWpPRTi6HErljYj7DKFERU59EOLbCT1g
hhuq9gO7UaNCW6i2yoqSSaZ+SBxxWa0c7NSBAh+B6fXsonHmmqPCoYWcwdLj
9QxRDv29gNnb/xepZC93k9Unf3aA4Q0fuR+5UsMmNu4DOe9XES5btm/jjfz8
bi1CRBCZYI1tsONRyqGk7hoJM6PZOI4Gcv8lGMBwlyiKtVmRIpKHEOvkFckQ
dP82pXdlS4+/7L1smSNcFvl11B26P4v+WQXNJ0DqikafZky6J//ylkBKcOnd
3aobiYGb1+Apwi4vNCh2YdRcjmpilwHbVJ4iq0jAjR7O7b2CI+3UDy7mcLdp
utSMJlUO1ybw8oUHa0iITswU/6lJf6JdxI3oKci2UG6OE9ylqQmtN+XM0HgI
e7o34cnDiz7TgN6RnbwiFf019s/fnDnmjHL50nTVe6NH57dPJFcYwizzm0UN
KbHj2ApT4ZAnSGOT4hsQ9z4Eg41XkBn8a9x6ea55Gsi2cYjs9AidTmvz+8N2
+z/JSikAXovNa1k9omMP0Mc/Y6Y/rz9shIjQo4HHi4vlSpDQC8y7rs72KdvR
Yc+x4u1mqAxLve6DOGDK9Gx1O69SeSwkMBiI9qfLJ/lvalS9qoPRJvrNrTbd
2FxyOaZkoG3MTObSZClBXLwN9yBCZB1JKqGWWQ8FVNNz+kB/POp4nKot0z/S
Bn1f94Jk+Gi2ASFLnFlt+epAtROKwfdHyJvpkTZxn2Iwayx0B+OwrrcuRD/4
lFVKKDK0wR8Nq3+0sZ57ohRodNxP1Y8H7kBV2wPnedUnk/pD2BsY4PzGDGgt
ty4qlsB95a+Pje4Z4ryQBiDbPLom5XxcuqXnqDA/099jwjaWA5yW6Cr+hZbF
2yB37BoPBvktgtBjBKP1M/F4nbLN1+FNQnDQjUJ86jwWoBB+NS8NCWPQIPIy
33Z6YrpP5b61fxuS0JEzV6f44kj1rvqbRoHFEFnoVulCVjNUNpn/gYvd/3dp
Q5i78d7b4hw4jUfakoOOoLTBC7Y0wvNwwBHJJYs7JV6klv3DfjrD2OoILAIL
ZNMNdKhcnkNzp7liDE9BpBMJQVOGm3neYaKVOSKxM9o/0dKpC6l9AcvT6Ato
z19UwcM7iUqx52Sd7N55R6fL56DvzXwkmZdaXteplYli8Pen+5nne0TmPoNb
qY6dFfSAICAha0kFlQftKTBK9rSo2lBcYT95zloig/HpSReKcwsfplvuW2Ke
Az/tmWbabGQx6DE/g4mE+QX+5k/ddbaPzh5HfecaOxPmdyzojwKe+C2NG3WA
HDv+u97ibJgZSv1DDUIxZfQa1ndtoa53hMwf5kAfBylXuUuZ+xtxyEQXDcnq
pS/YNePLoFDUcqCqQQjteiaSFYcno9iYNNtBTkjKf2c8WqYM8YrMaorpimxz
b7Oo2WYthugGD5bBfL0DqhMYLUZVv/O8LPzMgy1C64s6D2d65fWzxIs1ZcKD
v23nprAnA243I+gbDRBPMDQsTOJPMERaIfJKsTsJLr9N/KPYWMtxyh0z250q
DQlKvClgd9DpRLqHEfiU5xmDiuBG2J1yRzm/qBYzwTsHmLb3713V+rBaSgwA
kOFkoB+cEjlX89sGFFdPGFMPmUhE+mkASFP2CZki8KQiv6aqb01VOMhUOREV
L9rSCon1gZY3jX1VpJ2YJO7IoaJHChSxIAMu3Lof6fbc3A1L+4FAzJz8+FnF
KDq7JuHTikJihYIRDt3UZbG67nsbYyRBmQ9p4ReVPjddmZP9j3Pt7SJxAcrY
J80o8Yw5zpPgJeKJUuRvHzB5jf/BMjEWg1G3o1O/a0qSSYT/AoERNITeeOl/
DrXf/nAEKZ2H+vIuaB8F1Q/Wnwgy7zSEpkJqjotp4MJZfauomh+pXEvLySd8
K0mNL6msy41nRrFl1lB+FNvszER4FCcnbhWVDdCKgsJ0QD4x0K0Oz9R+sCIK
jGUwv2qs19hdpiDyIs9wcVCUjNgxSVhirWdiUAzMVS2GgDYEvC7SS9fmOQrp
c0LrHo0mRlEdtrj4Ce3I455NjFoufC3HUlo9+xdewewBhd4/OZGI3Ny3dmHP
uRM6QaVZCu7IhbohE0aSQpO/+KiVpTLcYb53yxXikIBN0/8A6lma7i6A99OR
4yB/gPdS0fLyLN2GtZyGluLtwr4QVUJSfQHshErsURwuRlc2o2aZH8DvT942
HWTNe1PxdL1czwNvMlLBCwegUWF5ThVncMBti3/Sc2Jp680NATjqeLfgMQHU
pVdIcVhAF267G/+mukvtGHVurxSE3Ifgv9nShx62mb24ZtRxapVEVvDexcyL
8hTU2iOWWmLnG4UgW0qdtSGnh3gY8a886iVlqjX80BJDcHDQYHgfG0MU00ns
neWsuM/URQDVrdyD+ibyJNebV4/482bTYkxtGXHhBaU/en4m11Py4Fx7jSGt
Y7h91EMN+8gYZiB9Q6lSvfrhziEQsMHq9biZ/PzqAJ8PeXPZ6j9K9jYFkKU3
aLqoJkvNYN+8B/g4e8qzHaYvNcVJHjXPr3Czn5qTlHDuATAryUwl3AUmn7dl
v6XWJ5XLVu800XsNP3KQHuO2+4Irw/F8iEEeDTXj6PpcMhJ7F8+NEIKBCFge
512czn/uvHwLaagZT6IxrulxEHaTdGwsyFGu8aLsXBxrG0PtaWRDH3t+Lka9
O56CNSaGfhzJRWvlimxNWKV0A2MXKkr3WtJ7YUAn3xwY8eb96UfeBH3uuSj3
3UzGmzMUkg7JxOikQ6Afbyov05g//SvsvP7kbn/sVn9JDjuVGuHghvRlo+Bt
nL8RmqvRgplVrM2ldGHXn56/Ci/kYSDXQG7qSSbrRvKV//M+JYBKD52jLs8V
1LYASLVlvFINg/+Wp1q+/99kRu4GfYd/Jvjiyt8ltdLuoOMTwUcWtK2KoVVy
MF96Prz7aAPNKRUZB8Tsn303dE9E9RmHkk/5JsRD7ArsLi+JFFI0JxdjmleJ
TTbslenhMIgcOiQTNWqkvI0MYhpBFdqrjXAs536eHcPIQGF6zZFlpgc56pfp
UJ/xuSNYN5MJ++2K3S9Xig0MqWEQLaej2AVW5gMHcBtPbhl7kJ7pl3a4pUQS
S5oS4LveHF3frhIQ1/yaN9gGaYLKWrg1wtkx7oRMuQXQKMGJFv11D60lxRz/
Mwaa3jdLuOw6ewkmaQk/O3cEaC20Wh2M8p9sTvt2NA+aFB3wdQyTdlirZEh6
dE7D5Frhm9RoOPfohQsa3Ygvr6PBZ0HYxHskCEwBiCEgChD5DtM+TjdWHWmF
D5Io8heC9B0miKB1NAcvlT8q8UdpQImgl2LCYo2MO1q8WnEIOYKTB6xwH4Fr
0q5OPV7FN61TwG1YlXzDhlYrynBUmdkf5cZD1W27pZpOwLTDBfNG82szFa1S
aVA6PH/n2eDFeynC1RUP6quf0ERa+tExWxfUxN8Ta4jq828DbL6eowyMTo7W
aE/ExGjEHyQEWtFjSwbnovzYHXYbW3e4j4umf5m8HYuzxQMSFGdRRP6eoMt3
cSjWnUrn8KfjIg2SaAA2NOtGoeu1KkSa5n0ePVWh+mFCQ4eHg/IrHvMzSX8Y
ArXtuLQ3oPXOVCKlU64KwE48A8IzPJBHJOs7lOqXuogpCiFe19T/kKz4++iA
DQVpj5KkeXdAc0fhIg+e4n4TbNbsyTRbUw/SPnuzVrR5UXP2i2ZqYnJ/4PQt
49B9cmGFCBIXF+vZlfgBW/bFeBnLWKVe7BbIH0CFqP1adQm14qAUVd263cIQ
gChKwNX6U2lb8QscFrz9n8gnd7ZIJymO7iPnyCagaLOao2D5Z7IEf6c94tQn
UGUaYzFsSGvwhUSE5XCddIDgT1C3xrt1mTDxAPCe6+YiNVHgDOuMZ8VOKJRP
Yco3SOyCDOXphAZSzCMYLw6ZNZmwNF72qBV3WW+kFRUEz+wB5AO3hUHpgGwF
UjYvh1hxRBh7+Z+7MDcxYVIH+op4yC55MoSNmbW5b6r59qHK1XfabD4PA1fv
XsofEhb86xx1GbkETErknyMw+yqM8LcSqLHW7sCwR99JJ3uXdhcrpOI0Zi8h
3iK26FpdIiy4NqhvKqjtBaiO1N3jb6VIEzGfmwbwkh9HOnwWNB0d2SkCCkCD
NMPSXvIK0qxVo7TQ6QzQ7RT9Ut1Fq7ya3bmDYAcxD3OvnXkCdSdt8t67GOBu
FUsbo06YZQ42X0cFPZz51l2H+gWVxFhF+8g2Q3vTq9t4fUcRl+9/mpZDNlb1
G7yVn9KG2SdUkEFz/AAlr/MdQ4vP03M9sEpbWt8g0PJJ+o0KxTztngy9OaH9
azz78wP6RoQ3cTPFPzhhS+nce9uR50oRRcHhf7zZdsxfCxyYzWtHDzlAvHI2
iz0/1Gwwmjl5wPAgST+/71BvDfFbn7G/AeateXEW997IdEBQNAPpcEDuhX2j
4/ATWHlsME5fJW0OulTJZt/27QMs4HNGYDc660OFxhE7L5qd7DP7/WOeDQ58
O1l4uGuLPE54V8Zjj2QeZy2lFvRLFTtmBgo49A9JyaABeif+dEPU8rCncJOH
Sk/zwexie5Y8Se46n1FYrCU1+qLOMKPEVlfO3h/8+FA892OmjuJRxjEJMf2v
m6wd23Er3EfuIPKXDV3zir5yu1+Wp+Grmik+KpMjej6bbHLK0et5WMKqRSZd
RVSvQVmCf2fx2qswyuGVoXePhKYCSMApgcQPmR5eDRHuUDgJoY64V+RO+b/D
RIbWsL2x+05jShzjA0sli+MUiKVjhW7yzIlS0wEbCSYKRkyxs1xODFJjDCbB
mV91Rm3mxXI6f98sl81f4nc8QSjHfauvq9hUHQUCa9NSamFYbVQXlIvhksIz
xf90zIELdKL/mrI78kcgP5JdrMQAIXVPaHOKWgxqh6mkZOZO3Zd4vLiSFJf1
bLJJYWkqLha+REy0+67dthEldxdkeKMZTwzCci+fLmOcljvyXP0CndWdFyXH
s5anJ/k3WQ3jEVGCALlVAaHws87NdQ1+vPRO9L0Xjl8VCRIVyaAY0u0P3Awq
MkVjOrEUYmTlPoo/7gOx+HLfUhI8N6djh5v/MVYnPW/7LfwKmt5ZcIz3+ybo
G7sGX+IhoX0Cb542XdmquXmUz99XZQJFGZWwGqi+pgw96DHxqXBSnI9XR48o
lhWTGkZ9KoMUsXUKWU4ZXbM02cKsIZzUPpNdb98GCpyZUmyiLmMcCA0iD8WZ
PI4l0nuJVG2544rdhEJYQ6+mM/YEtjylWO78xW7Fqo5qO2JL57iOygs36igU
lmBpw3XD5+91PMMIqYFmDrHWfMYD6aNomM01YLzsL4cZbqTpCJRLMAqEiG2U
Oe1rFlaJ/c1s78jjJAY8phPbPvDXlKqGPGD1BPAT2H1UrGiGmXITmxYqgj5q
F4K1+WI2jzoCELyQpWQmMTjvEPjaEuHdheB4MyfLMMwuieZaDdJKab1j0E5M
QJDV1/gZswp/3fDp7aGbfj63VmJx5sfrWB6aDRxekNDHMIgbXvp9R4q2cH5g
SqT+w+HkRehcPwUjs8IdlPHiQeBCece2l+ETX0hbUr5mk+wyO8s2BidZomVZ
dR6eTz0Poi/h8pWtAS6kBJScgzfRHrqZr02+lgcEeaLNMQNmvPIBGOf0U8KO
BCUCi3pfEXu5bZK2jrTrpGUGU6Ok0ByORzl6tPQF93sJi6B8T3kN2pgKDB0l
5RCL957JfJc1r1NfMsca4VuPzVxWia30oCZkf7Vx7WwjK6PWP0RM+oD5sQ1u
oe9/XquvX+MNjtLOpb1CL7XWOq+8V5bVMJRTvS5Bhw13VvEA5d87dIIVKop4
1cWTvONU5rn9fbw8V2dwXdJpeEi6fT1sEkJW40I4+dFYS4ew+1ReCL20VyqI
MTEm+PnSHXNFMR/Z59AWqz3hWqZkVyRVZ7md3nBN4fao/b4VzZZ/iDnE7TOB
0/SysrNta6rQ3UaO1DGji4A4ZfXE06NRlYWGchjGfM4lseH44E0VLw9SChjv
2ERvgS9N1RT1iDFZXp+KbLjmlvs9IkvSEPCsOCk9HCJHFPeAYqp9kWES1u4K
90shqqcsLw+gZg1RfvnzTfocmbqrarCyItFFZmgdKqnfAsxis6CqBZjc3bIc
o/YzXEhAPtd7cyxoghaRgxlDCrCaYWOTcLk2iKYPN946gqg0gt5ZVG8ZZvq3
0I2b2GHIDbJMPZTwLISy8PRuoFLmL4Xr8W4b0/bjbLB9nMxdGyycMWOtEMTI
sHNuh176RTquvCDjkdgRs2aZ4SN+xLTFae/yDNlkFLKYXuXzEXLsgV1brWLp
CTMvAloahCBLiwfsQca7OKDJoapWHMWn2ePf6obxqUJUuew4dQJuHROOyxrN
POsG+Hy1D+Zj+Ju0dmX+6XrdV6vSM7VfVkdpBuSdClXxMy7X7V+oNqhuhW6f
JTig61JDfzGQKWkQV3BfsIscLf+UOqnPQwFpFvjjl/Pccf66SmpVEZ5ASmu0
+9UPAKiNYd+KGWclmJLp9KKDAcca7eyYhqSl2zsf94aXawtNyW8NXiGArAa/
BuBQ2gwuiT9fNfD+jE3Y6cxbKp1rCm2rtVeipAKw01oP1Cy0p3PSLQIlb/sb
aJMcNDFiEWLBgHT5p//zkAeo+4LKHiN+/ACkfW2euE/zKdvpHxTTylKZIDsx
5gtp944Lnn1d2LQdTOTpb72rz39Pd9mTZSV0IBG3O4Txs9mj4TBoOPWqmXTt
9kvlAWQxiO4dr7aozLmRDtSIvZbTLw7hVPQdlsRHEBpWGOs6zSoLHkevX/Bw
59F3ro3aN/ixvo02n07uBOvKov0iuRg0kEWIZqustcYBUpQaXqWGnyR1E7tj
E4OEqUlU6H3Y8Th73gpYuaO5QzT8eTnWFCdFrYY+gMgexCwL74UVB6OuEUjO
I9CvqmqQ8YBNuuuIiZAFNeFUHJiHCVnfWA5SQmEIoUDIrBYB8sF9U5i8vlGd
34TYT5JJm9MTsqmz8gttrjGFe9CG0QZVshbLG/3jEB8R45HPmPoM1YuaMgz7
Ny/HGvJ7zhtHJVO1JCTKvllpm3dN5avFHBHY5iqr+EAQf0S5CGcnaTf4WrAC
gnX4+afCLkqwYsM4X/iriescm7U7vOddodwRv7SIWsPVxGn+f9yjHRVmsWQX
5FFZ/LS0iRztvZ91Dhbi5BHqHJ8/CsE7o3RWEF6NLvHCwmz6IaZCOacWQAmn
TxGJPoU1s5BQcG1MtQZ2pkuMwwnlL01FZS3DfGeEE/Uio1Ay05Xt2E1W+6nt
r/r/hUveaEElhKZbroc5JkYKRw/nrNqDpqzJVG2ub74acRY+yxn98RzsXU55
LTWJEFrbx6U405q3zdBoHhCeqKzTZAIQOd9kFFjY5n0hWdMYSXlCqjcr/JLy
ChS/rQjaxeDP8iMOhVnZfC/6n8wUGdkLkGPc+XzWlfQX5FTV3Qsg/u0iGfoq
zAOxLMVHgGlZFWmAQHPB5lQ5eYqzF3lOW2ff4wamPjeCGqWHWWG2EB+lx9ES
XviYTqV1XEEXNRLtfHkgx1GkmiBRJvzkgK9RgCI2/35NtpKQbVvZbBw1JZjp
Ax3VqJ//qV8yu1N5qugq6FSrH/+6PM7Nh6Jp+t7UW+XU6x8sh5C4KVpExC8L
jo5Itre7bDFJLC/Nx+RSyB3eMxmHYKoHbt/sGsI+PCpkPR7wwoYysIu9eb4U
Phb6NTBB17x5wFz4M2/i0ijjOnVG1Yqxf9dDry1JKxV7ULypxrwpHg9eS+QU
H0vbq+GoWPyJmPPZF2qvrj4kjidEv8jvE6ba5ZsPALxpjnMDgI2Sa3yxFnUE
u/Uhe/c5khXgMD/0owgMkRaapwVkhRPGTPJ5RuceuNUmEPlSKx+e1KCfPZ/U
/Tj9VSWRGg7/BG9uhrKf/QVy3H3mbZtONYcfK7yuom/jD5yFiYhoAalKgEjT
biFIyyKEP2rf7HwOFvcdGwaPhwT/RiwsPPD22ZeuiXs6sOLO5zxu8xIifx06
kdy32Z377C753tX4lg6HNzSL3sINB43LNd/Glww4GxhKu0r7NmoRJZc1lGMy
zvZPj97Vik/FyXmTDGJ9ayQgWR4H5tDmnt5/7ujbYTjwDsMuD9rK45P9J0nb
RNqr2F7r37WfNGsWGJjBGIf5fKw759VFeMIHhO0nD7+vg7dr+GW6r2JawtiU
DDmWTHVpm2iK+1fW5j+LAinil6VD+rYpW+wtVjCK1MGtDGHBdwxWMWCT7e6x
FmSfdGrJkTvw2JJIn4g6J0kGIyIqio4dj3sPR5pHJsKJIs0jm82GncnTo7KY
PIM33lAkIZHA68lgpcdfkd98T8NvPzWdfBgQeZgvRackdy01eVdIZ6lX4vC2
w7P5W2LMUhc7cOkS19HdrNCUdBfU0i+ief9PGrwyUPPdR9WFFdng2bSyz1X0
p0UgQAzrZ1kXwgz2lf5keiammaOMtHU3WirF2MeXN/IddYR9uFjOfGkSgXnw
oHQpehIDsR/gYE+I0upxrGmWbzlCCFRusbJtaIDFghMoUsAc450aEvapLG7h
Dmbh7NzkC5Ms666trvwU8lI8cpONxZlbb+JmuPAOe3DDcxa3ziZgAkd4CVM7
7nQtCMCBqLVRfmvozE9WduioHAF4RQTKCzxrVL3SqVNHg8VoDm4qxyBJLi0D
5QJNEzmgmWf4jvrrgAk308a4aZX83TFMivW0/QJk5OU9mtFz+CVkCNKIyVmr
xlKrbDy/qgErIGp6h2FQtspZ3K9JP0MSJJCc1r4UdA+JE2vRmPxepFXDLu7A
RViCZDH0Dq9kDGXAo6XnIB+GvPID/QMIFLSmhWSG/6YLL3e3xmmhmrDTQ1p1
IiAeFRk6vRUFkcz0FTasizoFmcq/1/dF/571YgwZmPlQgWVqKU0PtOX7hS7W
JmnrhmlPUfP5MovRQejdk/MJ22BEXVf9o9WKwJlb4+KZ0QXIM5lAMECVHEmC
QsmnYCnnUgfBw3InpIMkvRx3cFP4nuDOd7v6w3iJLEJjfNbK+zKCMxwc331m
6dh9G0OGtAPMo0jRYhnqSjRpD4tn3173ex6UWkjLdpdZm2/nK2Syhg59xN77
IpUL1Zq6a7A9KolOMwp6+WMOjLsJ5vF5M/DdeqDHntAHF79cMLidtdsBvb7F
BlsO+eR6N/G7Ef9PGUt3P9JSBx/Gwtv+LqdpCi95TOKCxeZp74JYeiy8S8ST
79mHZ/7uv9V/yC9u0HPKt7zaMU6f4TKBKpYVv0QF5xaLfrgIyPKS2iR1PnnU
7SOAk493eMxCY/Qvw9iEYAuiDINH5Wws5SxK8UpOLgBOga+QHz6/IaoPHmw/
9TFmYIJChNC9+0F9SDZTyjm7zv15A1yDkEOanwFK0kH7upRg5YWOqhZen1Pt
OF8uMstifDFrkmqit5hKBa1XEBjjMLjgv0KZFlcniXUk5bAaV0mWZu08CtLL
XUJ1ePoWnIJ5bmNMnaa4a3rZodMpwp8kUf/lOHriz7Nsd0Uf5pbAzvDydd5q
YOqWEnLVDpMrtsg9RJNGWj4YQvFdrShfku/Q1O8ZEQn/owiSMJYpZPGHUGr9
8NjEQtv7sPWFwqMTORzSNVnSZNuQ4LWNx6ysgaGNm/ePVC6zwLzYm7aQ0S77
8SV9nuf6IHFwZ5U3776g1Qrd1SpplWbo8gX+qT0wwOZiF4BSJd52gHr5yyud
sMHWQVdJFeQO/AgBWHCcjiBImrI6HvAOh+XfVNdhPKZQltwTNUmAFQwxBZV1
YGYsszVOfvhg/IZCZpbmQ7HG3vwS+JxeG7wmc+kBX14KLOr84Fo2g81ymk1n
GYlgDN/p/lXGuDQ32m+lOQ+RSpvz2VoHW9+sw0/wPWRvshFqHh9TaMGx7Y9s
o1N+ONJq6u3rW4HhqWMfiW+Gm5wdeNsSuuPIwRQgwPiUPllHNoVV8ev5eKPw
XV4AiUAWQfp6SIwUrDDERXRupyQu2dt45uHhjeym296hzEgc/Tkm47sueH2Q
IKXSJ5vt1H8UvYr8i8AEzgxSJNYNf1YONavly9H7SHQKxt573DkNKBsi1ggo
oULcU5C+kxNNGtSm01dZBflY/Cv/K3AK+8InuNN1EG9L0h6rXI22ld1cX/Zt
aYZDmlwlpqQtc/5P19mg+p/zdpkDfdY6w0anlGl4bI3e91JoNTMGZYfgl1Jr
JTsyA9LrvMhg1tDWSD40rpL4PxhpOUCAP+ZikirsZO7j71msK5QOYPAtMMB9
NiOAlgfonka8Z59Ea+szMNr8RTlSB1WqG3wt8CiXiRk1h2XEse1s9sf8IVtT
Qn4FeoWMmPOEMwMnUKelM/oCGjY07ensMliYtHmoAVss4swrAAx/3GQQ5d1C
1KYieO+sTZxoyh4qmX1PzsRvLru2E7ot99MZZKM3gqwLEJMvDU4DwEzdZXyh
nQkc/l/EGHL7srPbY6rzUxjs+pqy6e/E+J/uXRTWOWoMIeDoFg7V4AvPzf0E
uetDhg41upJUUOrlLOzviZfzhhZAhXh/fMK59mms5bHnbAY61CgrBJRqyc4e
a7gNgnYgpsRsYyQ4rTulssnrg/E/I5WS3y5WtpN57tYUisK/3U0qHWewXOPN
2GrQxZn92ZQIlaIpuIF/zZK88Xd/S67tBxOnpnuxQcwwC6IbKNuTj6cYNyw4
Te3G+mbNeJoReK5kKWCQTrVAvca83CwvzMU3cA+zEtBLmJTrMK/Kd6Fe8kzO
jMgvsWWQPKtacSMhKuEZ+8A5khra94P10tk9uPMn0rF8cTiA2qLNa9nfTclD
ZtOySXT9oZzb2HTGN8EJ4ycJF4YQuVvZPWIgZQrBNoa2ScDsIAamjRUjXoNu
u0Y4LGWwYpJt9wBr+HAybAPy7CnMxAEjuDpJ8SqigE+7Jx+WU+fnUab/BZuA
gowJdjwUbs4V4t5AnUpIb/qCcH90VRcs5iy34LZQFSNACNUaJugAR2SpJf5d
mLVttHTs0JJYka9Co2lx1IILbM8GiiRzuueB5iKaprJyn5Y4N9XW8FNqAPMI
+hFmjRFaBwdCxYxXSexV8yDB0AVofiB4yNc/dP5mtl64umaarM/njkh1X0T4
4XYJNB+oEhDQEF5lmyAVwxeOxr/oCCwfz7KhN+HorU9iloV5cHNH2cwJCgiT
xqWKu95tifkqhp67eK0HeYmeriSA3FM+wuT6NEYfEmNo8apbIEVu9KDssW72
zrZGb9CaeVX4aqdFHGEujroHh1v4Zftbu9Zzm9L0O09DWmY+TsQEEuyxPEpK
IoJe7dZJObQtRDXHTFgGW+hMSOgSJbUoEy6vx/mp+jfRsvQKx05OXDny7mWR
0xJDJ+LD55mqyohrsJd0kEo5MklhgVqfQ9fNNGTYaf4eVYhiisIiEo4ZhPLV
X6zw+1bEUO4pKZ6dmVwcTacFX+oeb5ayoFqoDMzS9aty6lQJ0sCdkUDO4hpx
8WoazZGbLjnFlcDe2xAF/xiqOLv244jMsyYiDrLZpP2g8KcDnsnHJpZq7BDC
4YZlNUJVGqCx4Nc579aBv09prVZyhvYGyLoQm1GctBCWndxq4DGKRi6m6tir
xrgwB1mVZI4IM+dkkkoXPebcmVW2HZQvBHM9O0PprNe3AZCNc0ZvqyQNqpJn
5HjuV6aQ8S7t/69jnMJE46yy0b3pCXBg56ouXBunmfqTKibCZXlwmn/ZN8d/
uRSLzUFC/pSIoT1d5XtYo3pNoa0vDnkyg/Er/LpOH6xITPZiyYePuKcAuWW7
vYbSAAzCSnc7dTnQJviiWsdtM4WiI6e8dp8wwolx0tpCYs5bAY9x+Q5jdzxX
9ChZ6Y8ib2gSnQ2D9TC1/r6RAz8JdZPHAoqDcahExK64rzDDjJVkqg8VwQa2
8vPnwqpHCdU5/iflxESiBxy4DBAJA/M/Uj1SgTrl1/Fs+nEEpElEf26QGzlg
WWvDk454vYJSYyLjrddUtNAt1TYCFfGnDU7yuY4hB2+eVYzsR65N71axRdGO
J45HNrQHEVn3Mx91hOFO7F4QlFxzgY3nUx1yOB3IMkr9qT3cH9QbMFFu7DDN
xpmhd7cleczx07yLwVbW98QCkWVe/WkSEAg0Ydmu0J1rIukbHX6YJMHNat8f
Ya4YppFsseO4AV4z9YOJ+iIr9FcWUrhSh2f1ydAytW17cj660lLL2kvFI3Rl
4AJqLpihcA/zi/2aEaYAu/1OeoF2JhShXeCet1ST13lxn/CNwjoOgs7EQIU5
bIGhd6iVBEdYT3xVXR+Ct7guI8xvqfIs7ieWICXqcQKwJ7sWDdd2mUSnBdP/
L9oR1O4YTT3VDEBd+0qpnY/5+mWGv2iJORIFGBoOYUb4u2tTusRrVpiirCMC
UrWrAq03nVn+3c0hCzLJrJRTud9rCcUuTu/+1ulbkTtEo4/SJuzAgk1Wv0eH
oOzngWzirGkLtkXPIuOu1v33iaOAfg4xFGWlLA/fm79szLbh2Ie04DPAIp6S
7CVBOEOthGgLGejG8rSerTFlYJXLzxl/ob2sUHLMf7j+i1Klmve7jqazDB+2
ZRf9k23fYTBi3B48Xi6RpqDlWV8CeArYzSTlmluganM3C21k4mUhOWfPKVf2
GbhtFCCZfpW6C025wXz4PhgRMyUeamd1xVRT6c0QlYd/ow6UgJSec4XznBkh
sqJ60hbOHUNVl69nY8QsLeIeQZsmEiQODOof2R0OTo9MG7iref4r3koZGmIO
gW5L0ar93c+fBMSPaJIkdcfB4f3gjEWhWKC2m/sT5LJzlAAaG+/NlNGQq//k
PT2K3JivuHOC+izgV2LpBbW/vOaPD0p2ZVbLWPrJ47XI11T50QozR56L2IIO
PN3IEbqIpijXDGwNjol39d/1U1irbeVeDjtqWhhJaidVSI9uU4Itm49dIGLW
U/Z/3OMazQu4APxhJDHH/dkpmt+90H7qAWED/2UQc9nuEk9vUGlP00yucsni
GrWrK6ytdROgyTcWAE2hDMou1B3qpe/uL+dPA8X3OueN17QGsfIalu47Pzwb
r1PD+bF2SvSehYsPoRphVRqN++lXGwAyQ5cEh8R1vnezuuJ/HA45MO0gVOTi
Jjj9i7Evp1KHoR6UzemaI2PXKAmgGHoceigkahHyACQUjl2gGaXeJBvkionM
Z6E/ovIRCJ9s4gVo+jcAqCg6g4xxTSx8zjVJ9Vl2AYLb8eN/7XNs0y9zE3eJ
p26cbC98NeJD/ikJvrg2MQgz0Ba0V94hXQiK0VM5qtm8o6h97Q9DApP+/58M
LLBOznswtWIMu1RU1CEmWzS/yChk7n0B7CqudaQPDdJFUOfznxX5U3osdoyg
OG9ieNvAdG+qvXG9/bZU1SIu5TXSQQp0lzDZdZ+ITYdcDJe3TxhohkhUGeAT
ekA7uT7YvtgR5h9zkMiwM2/x0hcSwWulxJtRR7uAdLZiUSttevonnmY0uZDc
5ilGGZ/X+T29l6qeeUTBa+r+Qe2AsElrqXYd+1nf1PzOLzFzH5qEcwL0smtb
/2htu2zswFDo6DgXyO0CuhB9nXog/yT7VdFETm08i3yuAiEXSiY0xzIiyJyc
bKztqsqDfoByYdDyPqSCd/6g54OuOkmHOufh2Ku7k6UJAZcY9/Qd4GYyBHm3
DPjL8ajfFCLqYcIDlJmOqyWsm9XeRRbSuCsjy8lHI5gDqj4EysdgjGV86ue8
or94mqEJ0sMvt768qPXWfn7qRoOi538LE1IPEitRVUfqrgd2XwJqTUGjeraC
20XewppBhKt8k//6PckoPaAQ+piqMFsjylICtGB5O2Ot0mWiOc6hN5wTEC+W
NGVei1f4+mkVE/mpzjkMPd3LFIIGaJCXvAiouqkqFkFrEP3Nh/Ab4vPsEBH2
xuk8DWot3E6UvQ3BZpVF1qksKcH9a34PUb7GVItYQ1wwF4hMV3MlvLagrNBN
G1XURMgLdzF2As9AEcWlJR+u5UGyq/UPjkXQ4hUJWVPMdWngSso8304439oi
SXkbxsLg3EZmUc546xJdDXCPwEZH0bScIR0idPTsJ6Z3pjPMyrEMFdVk1eLn
3kzx218v6Rhh7fQTgAkedN+bT7hfBVNl2E+ufcCl9hsL8D3OvVsyl155TMw3
vsNCmYDHvOW2SFjKRxe+3zfdluizHLlLPFswexGHJVYQn+7JwdawlYcGaxBN
L3qWp3l4UY8UCLWRAeOuuwqajk+VP/pYrD43zbym6b0VtWVtq9QXRRpuNXLu
AgEVklkpdEL45q9J5AdZ/hhcrlkcCI6AyCPZU86S1R6QFZGjiLzRzd7zkbxS
hkUzoczC2Z8XgslvYyx/0/zbGMzzRrhahCPM2WbYmsCfqYS3ZvRY9dEF37r8
KqLCVdtSRHDQeIAJ7Pd6uZFjGEElhGmR59USrqaI7cNYCEcp4SitUCQ1/yBD
CqZaZsRdQfUXGdA6MyhtPoiBQg7A6J4SFxrJQPtRXPx6I5jBcQdVG6hf4A5C
ASwU6l66PZQmfNPle29oAAATiUOIoz8UwSq5o4yor4inwhtLtlMnPd95nEG4
L50BI0Vl8zSW56y/oP4t5pRBa1s3D9MhgFNZRbn6MMyZo4dIq5Fv/RPz69Sg
yEwjHFPp16tfQQVxG6WPQ3YD+Ua7wJ/e46T7LLV5OrenXT88haUzxvE8Tbm7
94Tr07sQvPdBlxPUnVyMIUINRvyUYIOH9Nf6F0k4keTdd4RimZuxOZVMok4Z
TI9Zbkt9y01ORxi+ATqkPFg0ZhjhFmzUPLd8MdvAmOGkTIT87pXulY3qs1lx
a/gqMr3hitUlC+8E2hkaeL6jMgYJLU2rK9VP6l8Aaxl03mz3OmA5NoSz7WAm
kJZbQjPnWHBtQ/PYFX7HrVTMqZ2iwfl74np7bTknBqXAIoVB/hOoi8xlxqEs
/VfW1mNxo9ydjOcsY7RLXfh2ZP/dxmcw/h731cnT7TRGuwre73+MDwCeyqld
KBItJEbJ1D3UbDLIElB4nWPjJqIuZxsk75DHJqV4/09KwZlR+h9mKs3ySVE1
goDy6UQok+8BHZAGxm7zGkUBvVdSY52Yq38W5yoZ40pGJtY6QiEXHTyGC+xc
iwJCLeToHbLDeUMUPWU0tDW9JYFWE2iSXGD90RzeF9hHvh38inCG6Gr27kC3
8/rFCa0tLEqsYTKicQln+96LmN5SekjUN6E59q/wokGL9jJMCakjIVcl8zSM
zDflgwCnpl7QRLb4urUZCcqnnbjJkbIXwTpk5+sG8o9AmAodSUXHam+rYgYT
8eZ0Je+N7sU8ckErAdytXQqlWtWpVTlgEH4x01ZnJ9imwW9tBsudE8bAlm+a
FZGfsoaLr5JwWOm+EehpU+boejQJYr7mqTiblyP6VAcIs9l/PYHpjJnA9gq1
SiTfL1AOQ1VMYyweoGPdY4BGND7UVNb76bx8s5cJ/wn9DWXwJWy3ljNQqDoZ
lpcpOHVeTYKuV3s+bkVb26DNqLfokWpTnZwRfo/0qSfe7kZpDMIyRXA69HFz
9b9Vh6xYLD5iuA7IeJFcUimVvYmgKXkuSO1pXaLAjkE8LCm5IwQH8nL1PoM4
60vQ3lWDfueyOHn+CZNMWy5UU3yXWfLo8Y97s3gzha4GP2eWvJW2oqZbPtyJ
LfZpceRbGEtYtfdkmHUTfzVQF/aTPeIp49UpoUSJc/KqFMiXWiG0o/ti9zHB
OTEKWqOPXDdhTISAeunBCa9bxl66Fr3kWrepT5YsvMg/XaG3eHKcZR9Kf8vk
4NAvqYOPlmd8kKXV7gHWm3xx1RmOYw7gkLmuOWZ7bseWwPBIH5Biaq5JHzmu
Di7XL5nVBJ1/YIMhTGPYcxSv85If2fDt7jEIyddATTVNquAf4JGNkeqfWcZ6
bZbK6ggmie6Yir1sEhVBTiToZBDCopt6wqZ7Nw35S7KCF+i8DCWTPt6T0lW5
IhU5Dpds+I9CqD0kn+PDILtDq8E038u9z8w10CGz+dmdV/XnEH1dalIyfHEg
cBEGtOf+lqGsiUT7ESyskS8ZEJ9h4KTs08E7MnwYVuZwKYafXJsAM9d7kuQg
WJPnOAre2FeaOjar12UVNsirXsXYBCGaAY2V5OcocqW1WH97wN+qSQlGonD6
QN28PjyhWuIvXtbC8+Y28S1Gdf1w+aIwXjdVLLmsRDTEy2C5HrhPD8GzmCMw
khhmE8I81dY8sGmeD0wHsz1ubFy2cx4jOsmgyTWl9OkOjxOKiqEyYF2x47ND
SWYCKG33F5TaPrmnJ717EkBJFLfdYQrB4u92IgPsVcI1dr8QKSuqE2d7bK+N
hLfrAiZ/VhIkHtbFVTzaR7P7W0UuM4WmC8OyYVZdJM8h8Om5ijDLrlKFMMKw
NXqQbcHqzGum9GEqcfGKJLJA+6U3btoEBvQFbUUnlh10tQRHpH55uqG/lwbV
j0BKZRbsg94yYocRk4/4c2z4sJKqBBhWkI4Z4cWl5+wtQI3LHQpg84S/cSjA
tEf9THdBNieVTXPp4PJWkC6CNSmw9RkUmlEiZoSRa6DDpoAn5mMf58xoqCk9
XMn6W0Zep166P9yE46LMLop31NlLSJQTBL4dYRWjIXoHzPqC+qH8kuLpGg/9
6LkK/LcpDf0MMfkP60XB5rat/WZYYZ0ITHIcQgQxCgKZl5etiJb8lU7OBaQr
RWsFz2Y48opNoNZPaq3RcRWj+j63fJrwS00mdxZ5xH43ojqv8yPBmK4A67VY
uvJojRcbXBEqv1ggx2BgdnaP//Ml0fRo2JP88H9onHnzs8AheVg+UVnyCu9A
/7toXgEZmk2wHoiFbTZhhGTW/J8j3idc7FKyP4KASdxeUPG39GBjVewNgrhO
yfrBZpZ7LHVFJdVvBx5tFznOrn9h8MX/wR8I26CfiugvKFwNHgmmPI2frsAF
pG7XsPbzjsty6mPYXY2qgIBnmbxlCQ+cMFG7dnRpq/1rAo5pUgz5+AplAOlo
t3ulfqUXtP1fiZPIKpUpjdzLzOeBU42Uz9UwNXBQHa9shh/Dd9/I28fjJqeI
P23Y/JssuAIzO1q7rhMAAIPIyD+1JLOcXv8prnxarEIM6YJMr/IE8/k63Rt0
JR5s7KMtoSN+x1T4N5i96yy9vktQUYye9sec7/tQWO6q8Dcf91cj79QCbyA/
/L7j1/cmD2yU10mTNU0xNmJI3pR/JulEpI9eFHHq5v1hVwMXuOvteCEgziem
PBoGNmwwf0MuXqT2qEJnNzGyjFdZv1Q3tJjGuxNcACEZTv4jvZns2dER5eqp
/3CLFO0jcGvcP3zpkCXQE7Mp6IO5TpuECzetBkV/RgfhYNGXYAXdbtP0plbU
C3BBwq61sbiHDDMHv/UpPptyvFM43HI8eJFZOjVSEN8rVljoisLRD5Znv8Y/
A74xsjMngPPeiLkwPMSqA12p4a72/6UJJmq2q0WwX33ma9X29HUfaaLptczl
5IxMJmzeHzbR6HS7FKi3fpoK9fX9y9CTUNV/daSov2I47lUBiUUSfFOsPEp9
jc0j2dsDkGpsnXK23e2I8djDcgjjelZSK4jG/TbZUj1XUjxxREZeflQIMLwJ
8iDxQSwZFK/jPtOlAWPISWYyYXSQg+TSkpFC9z6XFYqpUhztdHR+Jk02caDy
6VCD2FE2pjjux7iI4hreMQwGFiFg8WdicDDl2lZd3bNBIDctzwBx+BMffvvY
QyfqEnaehAMHKszoWZfmNEroBx7aMbIINiCDoM0XaQsUSTOYe3f5y9hpRoo8
9XoqEg7jKSntVMSLUTqKyqPSBE0ImNgBUP/zVt9C6Rb+yYOO/aWJujoiEx/k
o/okwXKT5/QAq1UwMWuY09g6E6CIbAfvwV582oAqaIR/TnnUoUQsVh2O7j7d
dgRlHWKAEI7nkygEmjcHgjF6/1oXmTfOY2MYiG3p+ZG82RZZPy0l5QrB4CW/
t7/yT9KWUqfsb1mSz4srB1f81ORHX+v4GkqjfgpcaIqMpe4C4sp/HKgJcgBr
6SUjAqYrwtGGyFMYEMeAu6l473kCuG4m+6GhQNpUG1wiowUyyiZ7TkA93Ljd
ofbNDqpqbJM32IT2fpADyy+wj5pv0xm2+TsN0bXwCrnSzHr7qSe96hj1Qb0z
YhJBenY6RD0w34DCjPbMSG6K3+dCbKrDxfNDf8r/TqHSSZTvp89O1s4/CKA0
HhrYst7uf5qj1p7WffSQarwgUjvB6h20cVsr+TP+ZHklm+1bMSwQWyTYgKR4
7ubc99ReiRwwIlC7QVuFgDqHAz5JKS9bV9RiiKqWgNQnxQDwwgyIvU9VVCYy
NtTMPQiyh3AhnNBKRYToNfTUkB1m/gfdxkdcSYrL/vPNiAbgbXIFuRgCkPER
jK7kc1+SqP/EGLvLrdRIlsbXB7xIEeYgOI12HGR/DEKJDa/CBItVmKgPSZte
AIwtXyjzUgBDGHwez2dq6bN6sg51Cl4GD8e0q3gRej0OiPP04fpmwhOsbuke
rhCFznO5BWafAArnzneysBiaijOsGdF80AuuB9CN97hR94H04MHslSi6t91N
1FpxiZ6l1gGwaC4r1in5NMDr+L8Iw2kqKtoeWFV5pIp7s4JzWa6o7Z5X4bl8
KS8hrK6IgQmX4yVf1SYnyczBQXDeeMYBzD5qpODihAF8nzsfMFxzPnWwh87V
64PrbDkQ1AMvK5eZW1npIjW7R1Y9QHrrx9Co6Vfu5Z5601IF2LlFLJobRu+G
hk2Q2Ge7PoQxVbA/g/We/xz6KYMbUFURt0sTeDUmJHenfWMcpghAdi4uJuwC
/A+UbVmL1FUxnukc4TIsmgvZ/nJmIpJXpZiyMyoxwAdaVzy8ZZchxgdqn/Ya
6IzH354ztX9braj7++p7GbnsyEPGSFCfzRL1fPLb+bfn2sQBu9aA18O4fy40
zWzUUR/LTFx5ObHd0aOcZL5qlk0mkZaGs2IeunGcUnZgZHLZQ88u5uxsI5Oc
6r8OU6RfczObE2nYFq2FUc06NzCP3s8EVSvkj0qbEpczKjzUs6HaNkDoHwBi
+dAI8YAr4l3UQOen2UuXNw4X8JhUGo4UeP6PqvZ1Wxf28SLNW36ZfrSPnUhl
7rgCsZQw5UVl/E4Yw9SAeuJdogrNf7RWvbAMCjmTSiY41GGcAK0iFsVDvjA0
e7FBHhDjcCVhrvaKmq59P+mKbQmgDlitFMn5fjS+Wn96ZcYWTSDVuWnNCx8x
YlnSF5XwCsTWD31hIKr0PQv5OyA0RoptRWrLLlIqLQ3WUc5jhU2C99dcVnZW
uxEKI49XM2i4YZcjSDQFAc18/VqTJiRJZIVX6GKYF3cuRiKknCCDJDqJLnrm
Ge2unJqyMj1VRs8Y2mMz+JH3yFWTgjlot6KNmEFcbehb0+CRUyFXGA0RTIyP
q3+tUWO6NajXuDldvebSKGdXu9ujFsOPaSWlwl+FCvrPdFIDFKt04xb1A+19
QsgdlYIpDMO73DnTeZjJ+xn7UwEgn90KnPrd00ik9677MhAdwrzi2pDZVS3u
aPltqTLjj/TsAgUcF+DNbXUl2U32EEmmRFHVkZGNxOpSWW4dAt1g7jjMxf3Q
ITrc3/A2tp+yVMLvkGkxf9NIJX2Xs8qqRFNp9QUoLF2KQNaALVNIkzbZQuMa
hxSSWJLcuz94yn1FlUXxtZoKy+j3RKcrR8TZJZ5KvQGEJnLQDvL6d918MiXM
Jsh0HWx43Ajj9uw2oXN0ELLVWCDGIayYpydAbdWvdYXmTj+H1Ks1aFTMqfeC
8ockFX/LSquP8uP485vuMIasHC1+RcuARshQmDs6QqNNXNXZ4TnnpPgGSqV+
rnxF1/gtSa1ckqPmT2Kytb3TLa7kCbcn7kTwzXUlZBDVyTlLRZ9PM7mt+Rx6
Ckgd4IrjBV4Zt0IXSZfThOXaeaFq1q5K0O6dblJjcf0l1PQnBz9ugbta3FCP
08wsubHILwwFha7CH+N4WysJ2nGb8CcLWpm/6H1NohmGBb+c3HWoOa6ugy9i
w+VAWKmpR+HVGfhuYMAH/kgUtR4KMzjD7VQEs8p3TUUqR8pmb5c2N/Dc2owj
BYeMmqYLhaHNCw1XR2hLnFfYsokM6pRHWfH3IObLySYpmiRYwE66KjzVgElz
S/xehWtNPzfN0s6T/sm62PTkOF0ukE+HausRHIleXk8L/2TY9Bu3bdrItJDo
xr+kSlx5ZvhgDkIJCYGi7hZJaKeZ55alRPYlpUhjqB/60vjwFsGEgiBwOEnw
m+F5ZY+C/fZ9Po1VDaQFBVzBtf6Yhpgb3rqrriv9npHik9ookGjIcw3kkUzA
mdbBRqLDtMkutsAT0QrIKvK4Eq1m3L39VOP/OKTw6YXiFfJCCSr5v1eatPBA
/QqWV87m9ZUkVKZGIj6jJyuDO6UWAMm658sxRCDjfMp+6lkso0TcbiBE+7oQ
8ul8ToGqtzi/BEJ1I8YG2YkUk8bODj1i8u+6Sh16PL39/c9T7i88QnCLpetg
bFgvbTZReaOtbD5P4+yN6+tygp4TFZrQ7L+2741CaTXVN58U6PtShp07bfzx
4MobKK+968KjgCck/VHRqyyBENRN9we1LbzMC3fJV9hwci8x01vdMkpNNwVA
4rH4CW2D4WHqAUAsffKmFYM6dA1h92ENhko0pp3QK9CoACminH0vV0fEHo/t
nPu5q0Ss02rEwh3Hr56qwE+5Ep2uQZozlKeqDY56B3I6arECNywp05jXn3hL
1cJr9Hh3x6qv8aaFZ6V+mRDV9fInWvFqOpx98+4K6iGkWMmLC6MeXm7Jaaj+
8R/Ryz2gRgXvM4aNilXePaUenOlAzSrYwTi3Z/ScnscWVsZzvfOT6A+p9Aob
bgTsOnzl6vXlphTsWaBnvWD9YLiTKPN3J7iRXXEJukJokoXZZktfQDWqGPfK
1YYXc9SjoWnIBppRZiRR0gyd9/NC4BzVXECif2HW/XufjuKJPyJiI3xaeKuJ
HfeOnfsF3fZSZsPp+owO14APsHfJjWKz6V/w99cdzUtk8F5/KqWGU9HILQs/
epaNXOm0A05T1sJshyOs9mAptKG7knry0a2oPNWTD1Rs8TLfQD2O6VB7Q90+
fZgoeA0b6KB3ZAHb+XPCfKEms3D5d9a9Dyo2xIe3MBcfmhrpJiTl5jOajOY7
4yIcmWuSgI+d4LOHMMuG31gdLDxVtsM2aiR+URv5DOPNxRpQO7THsF8ss2mx
tRYLeINWV2Do625/JlUh9WUsJTI1HIRUdbNDJDx7vmR1qgk6Z+TF5/Hj61sG
0y5o02fB5+xOllVxg0jyJbLUIMRzyHfjJqHJNEhBbf7fS2iYwnX2YbJqgicd
GijgPImr2zKMIaHE8Z5ttl5J6cCZiz99lXf54tgnfaq4fRwve5mNvbVQd7Re
4VxChyOdrYGyDPOcplZizAhh5cEErHp/tNDc/YL2UCa64laEcg4UA1YygcN5
KFFZPTuAImG6cLclGwTJD8i5eLxU0HMSLl4eOMA0te6UtlQDL8iBqicT40CX
Z+ewE1JqQgjHJ0p5lnlxIrhyEG+lKu+bKNhnXX3dxu8vwHFqS6Zg9TfauIk/
OraJyIrYx8+6U20i+PQTpHvVdaqvr+xtzgY+vWSziMzbYQRBnaQL66ArzGxE
+n2ZELazR5Bcesq/UNQTvOsDipvsa3iUz1kpcrr595aJAsdOv7ZE+Z0Z+WiN
NJ3Sqn0U1pv/Ni6NgsxvzBFTyZJwvESYGtEEEEokV7qQtguIlr2tbA9ytyEq
7adhpIs2h5+RONaf0wKZK+9Ks1vQGRJOpbiTDIm7l7whP2SZ0ocS7F9wXE7q
DImcdEhGLxpUZnr+UHwJy/hknLUhUkrfIfLLnLIv23amk4dsujIEemy0h9/Y
oBcS12t6uHX/lCovH9MDQUwwdvNZLUUIlcxZhprIYlG84u0Rg9WGG2B8XIDY
6aO0VuEGs5ViP1Zm9heUQfE5R8gU6Gy1llnogKMm6Igy0+CT+pKdU/eoYXjf
ngLNAP+IJOj4fvbMxKZmvDWYreI7WHLEGmBJuqrXZBp8/m0f5rShlw83lQLb
jUEaOyCmv5NLnwifK/IEhQfl9MImfrthoY51lMuDOcEZoBIm5yoRH5VsdZyS
n2EoQCLmPleCr4Ok4It21WPgatUR4ExtRAmTAwd/i6uylEWwbCO2hTdWJ4Ow
goWBsEKGi7ex5pyLd0Iow8QsZeSXob9e8Jzo+WiLNoT0QCaX0+YtK+3hUvkF
pbe7O+zWMHDYUCUa/GBqp/2YxL6p8b46cwoPm9oTjdLQZLZhRAeqqwL1ASKI
tMl3ysnymR1KN7ePiVPrr1x6qYyBJrc06OyWjF4iuoVkIMyv+D6OVVN6pZdQ
UR2Alsd0BUqix5Az19+dlXP3o0qlRj2L3IJRKqb5py54YJTG8u9zmxIS1lmp
MICqWBgySR6yUFPBUiIAYu0kaBP+sCEuNoR65AmsCSeVyBQ810WODPrN9zMx
wYWg6+hDqGSZcshHZP/8zgLHOvYS0s79vn1aNFgOTSgLrMu30Dmy9Vu+LATl
/LLQdFCPYG3wyS26sMtelFKGR91TXCw1t1gB5O2aINnro3Qycnrvwl5DRTLI
vHkOO1d2wHTb/Xfmy31O6ZFJLaKkj/MLTzlV13caMbp4JFLqgrVYLpW2YZeS
+PjiClmSQV0lUdWjHhKETz59flPdDyP+v59gJs5IbOrkHoTHLdRZiyI3KRaQ
6frClycfUBaIy9XTD3DwIROSb3xgeq6pUXiYhJls3A/oNa0L8euSrDJnm6QG
/0O815wMl3TUWgvd4y6p8rTvKMug3U0uSd61V2Ho5Wtg7cJNXe0jGSD26RgF
tsWkAbX9SqkFv/PYFj3qrtO4UMu5c4Un30NIolfUnMkw+LqEDmh12cL3CCSQ
mVk+0tqReVY7B3D9Ptp4kg5wjZfV1m7BrncUE6rRrFfTBhmk0t23BuKS2gaQ
6dCGhRGGV4GNwritazv8qvpzwS+aswFpBxJBNKTcFS8BHguj53AtyBADiaCw
qwZqBR/RtCDBI+8pqBlv7gygQOn/RyIMv7DDHPzW4SiOFwmXoRK6Oom8JhX0
EDJGt31LwLvL3qoFzX0j83aEThvwMjwudIEjnFS1tOWVH45OP7w3xJuIH6ta
+MIuEvhgVfqL8uo5+yhEILQIbIr/uVitPTSu2bPkZ/bS+O+fv6EfpLPSklv+
KYpdBLwjPQ0n25s5lv4Sh8uXrLRNH10WTqiw5A3PjtIytKhj9JomCdH3UNF4
qOUK9jTIMdi7K/R2NLvGBZRmO0xiRlEMp/wxqGSPHX8MvlJAFfJuZ/XenK8X
F9p6oVXQgdJ+q7x0qjJOCiUnUJcuWkcJRPnkamdeV01GLzrmqKkXGGq97Q1m
d4/MxNw8O6cNGavBOssCfsgEEZGdak9DJ0+Qrmjb9TClRjXo3AOQqIrfbdAA
96E81EiLeHgkHbUd9dKfJHDkNfpcwIEZy/SrGSPwm3Mcet9760U1PS8my4bo
YsotI3YOvQfMW0zihwl8rWcNYpuFNtG2SzyNPInFNzPMcpxs+uLvN6yW9qSc
enw7WvDTZK4vm+vA2eOLHLy/abCW9tPMG9KRYClDSVZZiQ/sTNojWevbZ264
R7llqbe5EfftiH3TYOveu7kdSNgBh8PPsiJw+2i73lfYXoPP9KQ+39qlnavm
VVkza4+/q22ajfLquFHICsy69I3nBuGzb5TNHfUe814tsrf0Kq+sSNLfWnWN
tfYhRPByHDoMwULOhAnojd2iDc0M08SCpl/8tEI/7Pty01D+/61W0igeUIvl
qrproSCYEcjfqFAmVsl/03VOcgi9FLPiiSYaW5ebpNtCV207fE9pplbWfE1K
gm07YEDdvDhgb7DdBh0X3O4G0NMldPP9p1qCT8gEbrInmmFOuPkVKxQXDGHs
rCy6eP3LRT3+vj0AfOmzNcDXXo/59Tg5wek/CRO8gg2rY5sSyVCFvnHRDTc7
LqQX+bLqad57tu8dFtfSzIXaH3JXye63bWYuyEMD3q45ijyGhkSN9A5cJfQR
Tm65ujwGM0xha2cwRy5mlPDCFYspUHJ7yp8nsSxSNPLNfv6/GBnuAazio9fe
RbODoSkGL/vOEqi95tj0gf5Sta+u56jRPQHUaMwShKzweoamNB+ZhBNv5cPi
CqTwNPdExRD8o3c7MHH+QBjW0QFJqkLSdtpWas1m7VQ9eNzAK1cvwYfUf8wH
XsNGdx9E8tRCeuXpLf0qTxzXJX0D4Mf3jx59q/jtkwqaVJhS3GmxtTMpTibZ
G2GktJYTI2XUSnRLzE4CR5erC/9stlSzNq7IaPY2Ig4wgeCAuCDtH9ZVCF7+
RK1Yu12GexXlpCp6dEBruI6A+gqqr4kTBVIGW+asmtSVnjeSLfqbewIxCByq
+M+yACqV8msG56vJWP+FtsRViA9b4VbnYaMyKBUay0q1iilgp7G+S9m62G8k
r5tqRdYik3VzZT6zgBXR7FJTjiV9XvYVmGX4QSE+Mbm9JGlm2VMXZkzEfT2p
GfbCvWdQlA7BIHMGgBj5ho925jvYDvwx5bCopY22Rjw6wxu3Bb2CpHTPuZ03
4d8ErTXoP91EaK7zDoFF0M4aLS+vOxziZj59HgHo7qukR8xh34meKprcmVV+
avTmxLs9DeFVaWpkufjT9zkoFiMkCpRfKPATiQMJ9xP9FCj5YFH8U39Xzmq7
RgQ43wsKqw/CG8o+RuSW1FIZ9yy3Ehc1QIoDrE6DDCDGRSBnul2SdgCW9E6L
t9KesY1bjQrz4Hh1DTtinslmRtHOuC6RgGszRrylvFHkRffg5DuMo/pAvx6x
pLvQtUvxQNirmyFPNaXVTyy0i6WBE9vUK33CVPCkGrGi2Tg8KAFzkLWZoemp
WcTNJ/M+xQF29QGTCTu+7k5gNn3FGzXyVN255KbXpLMc3u+br2wcrztVAJVJ
W5zu6xPfk9xrKKIelVKmDketDca6oRuLYpmZawAirSWQNHeT7kLNCPGz9ZpN
gbf95bG8JZOIGTGz3nKJt7T9TX4IzBACLe+FUC3zDZ/H7JtT5aOnR5pPCeXc
37meg1QDknOgzKX2FlNA7GzKlC0NryGD6ZtbH6JUetMcHQXvfq90IMLgA68t
0UQZU7DvQ9oG4SsNrRZHZAbc0Me3cf2W0Hxv2d2YRITPndVXZ4LqACYm2wpU
xasUeTlMfwlA1Gg8W7o8KI2w1MSMNVQx90apUukx4vPKQxM3isUr7f0eNlys
rMli/QnKCD1MXFlP4wXrf6pJUv2SHQ+f5CxWaBhwmD9DVT+X/AcEO2WflE88
fBiVcqLwHV+4HJmG1nP9s6W4Eaca2mPuhUs3gDAHG9LlLidNvJfuUmIQqSXl
J21MJHm6r9DoGj6Y1WlR1HT1Ge/BreiR5SD8/V8NunCac3U742kXmZj1RQq/
pvNUoSPX1z51FYhNbTJNbYwN6P3WXerDWpiOcVAz/Cq1S2F2ozPxVCrOjcEN
gYtwv/tbh7UTgje70NVaVgQyFQE9L+/EVzgLN4djX2jID6v7WwK3j4BidxlQ
QRfSN402zMIo924TGKVC0PJWd0zg/c2r24fDqpxcrduhkhQKNuGesarppw46
XXm7IqXYvWUgBT1PCSHBipHFREcD8Kj4rlX68pH0/5Z08kszhua8dWDwnLGo
kKB7E3sFmRWa3fkTiGhQXPU2bzxZGbCgtZbsKmrNuYbQTh3RCeTfpIPS9nKi
aqElwU5Bqd63riwPGR77gY1oxre7NUh+1JpzeReSvfSatskbsbMjknGWwcRW
nuQnaRHcKgyNzKfZSv4djyc0xO22B28mewEu6O2OUh20Qs/2fOMWpWiH6r3E
4DW2KMptDrxppIzSI1ST1VtyS6/Ab6MZghvtrPGXB8aU6OQcsf3rsLL/NeFr
z6k8h8YqGurXX+hNKA9rPZOhfApKjke3cUsPMpcNb/MhNBbG3x/VWCphBVHN
okDs0H2zZY7MX+zBDWje/ewkShtV23QR6Xbn9pFQklZyPXh1y49VbkZZUEGX
oAYFxPTw1IvXvRklIE4YrVtGhop4lfwh63BMPgmVH1OzeNwkrRk6ZFPdmizI
OrgG1pCLlpZ6vjldkwz6M2QYdjEmUhcC1M+bj9YIPPzp3AIrl2p30aFqI2Os
mcwT8zIox81m+2y2Jk3rAaGMSUe/8v0HJH1jHHPrOZIRjDzPabyc6wRnckOf
MEnoVIRGomS0nS7WbQT6cC9sIPcaEMriT/QkJhkilxlVAVkhbSjVDAQ6/nS2
FavoJaMUeOAQCdwY2N5TSUUx7bGN25Ge8L/IH5X0Z1xY3o3b/wp3cATybNZi
xEEo+hbaU/SzT4RTAJwB3LIXx7RW/PxTC9zdO/HM0zmwaJfKp8sKiIWITji/
pYOq74V7X+QumNGyf+MXzaQgY79FCtbu0K6hIiY0RS3RAHpad9de0nicGki1
93LAdNYr4jWyUSJ3lXY5aKg6MotxvzCnAuQcRtVKmMtSEJN8aKJUvEWm68Bh
wbliUY2EAcSf3FrHOP5fCrFng982s7qmLPccXUlxd3neEZ8nZSEg49PoC2/P
yrm/Byx/QrxINLmtbgoiNrwju9a0qzI7VAg42tCefpAGmZNvieVaUsrYLm36
UZ9u9UKUk/oGkFsCrPUAL8or2IIn5x3yfC/wT80J7dkLq0PFUZTc1LA73V3T
dC4f3bQk5YVdfWyHh9KYP9FQhGGHXnvOsypmyhA60GFyugbJSaZ3wGRYVoJb
yOjyw3oU/Ho8HE2VEaGVoyBIG/cVx+ezWm0s1fjgR15QIf3tdepN6O9/gd7z
MCCbFAQDnujl/8C0LaOdVFYvbTaqErrNYU2qsxev7QQ2hdPkdwITzHTQm4pQ
gt1f1jKbFLAe8/LGO7pH2iSdUgvwByyLfWe93gujZ5JlugkIKU6U7ShHsEBL
Y5gg3csz74WN9Zl5jxFEXpZ9ecLGtMDTnaNm3NsTeXU0kIpiBej1qqXbXAkB
udFUxBDSTFd3S8Ob+D+108GmFcc12LkntQBWNocTQ/qa5yOxugSJNiyPhh+E
U5ienaHjgwzbQJHYI3GXRS8Y/0wgiUGk46ZuhMxHdAjxxask/91XBbSfeeqe
8effX8ww+tz+cAIdB2/YwRQVS5MdpOP0W35s3SxdJNXu2z+2NcY8V2ZihRjB
ntPdu6Zwc+pKi+x3VzLvqbJ9aqJueWn2CtGn26SzXjpewfj52rmDvuSIjlo3
mlXNOvWWZZGzP1c+sHrbiPHmo4OKd5XJdsCT+6vXOVgjhFJsOHU69CA7qiCS
e+yR6FkhYnSko3kMWzzQ+FPJFunei8I+kmoqBE+IsE3OCcdgSZNBj9N/9XQA
KDIn8nDwe0iiyZ4HpnjBaBLDtPa9fLFYoJNSzur+wuvfYMILMvkdVNJq71Vk
BBPXWPZLtgvrWmGeg8IAju/Pb+KOBejCRvhq+aWaegfJlfoz8Fsi81qpH6hg
NUuaUynkTxfgwt/W7wzMKm4yNQPO1r/59ZRIzSdhuqL6dqjxYhp/yXuMudMA
WbcolW/Pf/5akc9z2E413zyCXTKtC4+wTZyjDkTx3KiOQad5u/M7GvUuVFZr
emv0FqTvMABRvAjnzBbH7uakLTV8LWPUGDo8BAoenl/md/7FFPKCUkU/uaAL
e0goDr0hV6Q8Esn1LA8zMFmqyXHBrZrOfvP8Xz+I57j+3CdcuUsZj4O1cJ2S
Vk4ynEezrBeXQIWbWgOxPCtAIKDCoEVF2OEGj3Nk+/6zapUOGILHD+2bixBM
RLHA24Mg2m2At+OuoRVaBR1iCkaUfj7ikThSw0z/Ho1IwBE8bNAc6tqW+dSG
a49PqSSgEaOxBWTr2PVNeCTyPwVVReQkfPAoh9Tracff4DM+Uu2CFsoDuri2
rpViphOxjUjeCLq9pM53cLhcW0Aw21TqqIy3imk69ybBz8z9khS5hSSuyoxj
M6zqrgBQRBqe3ky389R7IrApXGWmXA1PY4ZT1H43lzi4Dx406c8oGQoTQidc
2aUzt7FQZnZvZYVl5acCLsKq0TQmsoO70TYwz8755WWsHnQe+17UaOYgDkUP
orpEtQOzC+h7Q1Vxtv24akYdc/c5nftN39q8HRSn6bLGYSAIosRULD79E87Z
QILBfrlH3y1U8/3xEnR9cZAd5SnTSOLBD1eLosyIYZd1IZBduxjX7aflheT5
iUJuXj9DxL9pQTq31N4Owt1T2ICtZFBwmXLpgxRbJ3A2wuhkDNdn+b7P+18K
Tt0iUy8qccOqHob2i0FtJeFO6DgA7iZ7f/ObAMbODMlvvzfi2K95oDvcvzDl
mB6ne9Y550mwFB9rK8g33pxZ0ZghesTyHJd5UrNJI4ilZ/nFzT9ZUQ3iGWTu
pAjVV3m+KZhj4QVBS6T09GAA8ASnN1krwnMvmQPRX6wLkgYIXDW0UOJxtwTK
3ybTP5UbsmhKykwUOPjJAaWZV6j0jAGuG5EDlKlbyHdWgsxRYCvEMZo0M8rt
G6NV6Xxu1eAVT+JWwZXiyKlgywEKXUVAoTxuRsABAsvcsX2gW95oYa3KSZyg
xpVe+1fBYjlCCTZP6lRmCeSmQPVUvwArSbSNjhFfgb/AaKcnmfL718FOhav0
0YxA6rxUNhf7qrRTrcmiEi5f5f31d7uTd2r7RoBkZ4+RTGZocxyOxnileG/d
e8mPw2yDknDGe5bRKXNX+YqMkCgTuFQj2IQZ2a9FfNBuH+ASL+M5Pr1iWhFH
q5oK9lBPxsn0xBlPeW2obqvSbxkmODviiUfVXmxN3yfbSpO8kYbH7g6eBZjl
f5dl2oyENOyNK+CtsL0Aqvum/ZXUmMPyQmf3Fjf2umneWhEGeoRW3gehmMjk
syQvwI+c8bX8x/G7g8TXBQ9pWzKbgTMrhk2m53jX3/J89rKq9Fp4ZBbGtFb7
iiaUH+hWOLc09aKKN86zbj4w6EE6ICCZ2BsSNbwrHSVB5/7rlquyfJWuFsnF
29DvLG/tJsv3K0dZYDJD9eIU4FHV3mb/mUPuOqmc4byHTud4asxnZ4XWEiqk
uK8oTozvkE4SUOn91m6ynpjpBXaD3vYpKlBJlDyyYuN5KGZyk0rewJhQ9FiR
fIzKOy0/O/QGoG2VCq273h2OdmbfCmxS9MrXsqR7fqeEYtxD2cTwwEzdWYMG
xBr8Pgf7xiVW4CXrgwrU0TlIyoJMbdTnl30jhlbjm7aHzrYUY1qeFF16FGVg
NjR23yYJ/eagtGMNvF8Uv4uGG1TAc2YGYDX2dBPgcKDJseBstICX04bTtxcH
4CnuW1t0VZrG5BpEL7mh1lcHL3nMuFUe4cM8B1TqbbgAQkUIXQjM88bVQZPC
eiuLF4n5+/T2B1PukFHBbh2jJ1qG1gc6Q/vi3aS8uXcBuJbKDM/v8g0ilobj
tPJXMFyEeBQ2yNdobybru47tN9VjPHC61o0236mgBwQoPGHFJ+oinAzyNFK5
ZtSG+L/AHltKfKYb6oG9t1kPm9mtwoSQJl+Fc/GHAnZp8k1oXCNUjoU1i1cj
KsbZvyJedXFuAGBqU8flZQgU2/tWk/EEDSnxUTGfoGq3L3cAgVqlaLVXBPok
wyn/Rn2FqYVwrpdaX2QH7PPzE953YewRnkgKYVpP6sjto2YgmlMyWYV6ybXS
4OGwFF5BB/ccB7pXwyR1Y60EH38hLwWKjVzKeTmbwUWSjBYO9AN3UJlyeCTa
cjnoaN20S/mU6dW4/I/QjYnl/04YTa4y5c0/1TCCFTkjR6x+cF5MQf5/HK4z
WfQS+F7Lf+Rm3VSDnWP5pTncbjz6nZWaDEQPvXM9hARt40Aeiucxrd8atRX/
I2q+MiVcrpvgEDAlIlCxAP55i6f9gZ2V08Q0CzGa1tKBpu0E7ESduIYDyNXl
hwQwRObels6awa53mQ6Ln88LqThDMPMgzVAutS10XjFIov3Bf5v4rovcN8cn
iY4W6sC57uRJnt0yXLwlfR+bsQkP17WnpgDkR6d76cB1CPt1LeeJyyNyrjdt
vuUBSUj4vFJ/R5DVhCyL+y9KEgQtm5+uWrzziygburbQQlFZmHh3yTvoLF1k
vjvYCguTbOH3Btcw/0C3+AHTxrzcjIrbR1SlumQM2+D59iKlKePYfUrivkwZ
T+6zByTk8BSfvqJAzhp+Qyhe/E2wsFQexdEA45cBO1lv9JKd4M8vlP4O59cn
FtJFL1F+ITJOrwp8Fo7sxGV+lLx3QrucRhK64E3er+c5FVfLzhMpaQn5z3o4
IEylTqtvnM19WdBQzLFrPqi2ovis37yNtdtGG4g3LWiSMkkiF/QqL9kPDzAM
2rZpA3HSv9wzeJN4J7Wi5Jy/YBwhWzae+ouaciHokSjtR2Mwmqhfot3VCocp
OMAXjML0u/S+Dd80HZdr9hzODeqAMbx+uh/lCQ/6hlW/UEf7yTgbQcytSe0E
l0pb3p6IgQgMyzxAMo4yJANZwJGwzEGZ7488rbipfYpM5n7lwCW+iY3yWxso
3TNGZbZAcAv6G/ron76LwiDYZcaibFBEMW7ix/ussA3j5k+4DAozlMY+1Cs7
aEzSea/ob9C56Hvlv1Jc/CXr3MFbOXY3dTKIpyZ87vWb8WEd6vly9Iwjfr7z
b2pYbeBNt5HUH+byZLSaIScsvR+K758svSUjhsUYatY2kx7W7gBkDYjCwXLS
Q5wpH1qJjDbLw4g5PRNSLSTLC1AJVkge8gFeBysQbxNeyzFgTC4Xy3xuDxz1
RyDTa1Avp5QyeEz1sWR0br0TMXZVM4VPcfZ3HRvXluChRX2fUX+KL1Egcsj0
DCPQaNIBUMfiEfKWPuDNs1Gpryo/HUgTCUVnaLm5CBzULYS6/3FPjiGEBzEI
9w/malOId+VsocgzgEJycueLU/vKTFOfzG6bvlS9lUnxAYdv2V07K7mkHp0O
FFqJz/I3RffvIRo2d4iZToYGvXtk6o6jPsmqj25j0LC8aI1hLZgvugxYejFY
7ESCiOy5Jgj2ILOGNIJjkvwApoKmj0EoMJm4k4je2wETULrxiRtlfy98E/Ng
vn7uSMxrETZsnpY5BmBB76MEVs7cTDqqTjyGl8OpG4bLS9Ry+Gh2h84j3TBD
GuSbYtpwwAquH12/iiQPt2+uA96n6crWgnWpUTU7rarYgh7AgUgzKnJ6oaod
G8GDM1XnBpqlJBG9SfKN/Q6Cu5kgvtu8wp38SpMR6XHwa3E3KGTyQmRfJaFf
7bLiWLdIsAWqQG8oIq5/brNCqm3jjYmWQxEHTnhZ/bX+vo5JOh6DX6wCdWah
WDxapJmrOepDDAQq/gtPKKcMB8NkLiYjz2WzKjKqSzcDPzGmtIo5lZhn4bH6
BeDwaWJmMwcqDaY3L6jXvfXLboyeQQ5LfyGPn1PQr5aVni1iuC4aGjcYZdv4
xBF9DAGGCBlXV0vFgN6bGeDXgXzxz8lU+PuE1AbkqFc0Bp2UnMGYoGmWc4XV
mBRyxXadEk4gXJOHMmoHxVfvp+BONh9RvMu0LxcrN/llR/ios8JOuCFuIpc1
hqlCfRPIy4GaoO8JYxZAldq2BUcKjyrI5an/JflNceWLQkLPiV+/UIz8GCyE
+hhdQjNTwvyMfRl8rgIhEKWhP6aZWeanquukpixyFOMR+Jc6WNqQCLRQ0+h+
HS38D29yxz/PtgerDQN9MEp1UY8cT1CPOEo9j53nbq2XQvt9w7JdVzQoSI8t
8aFhzRh6BPavT9tyPy+vh2O6Wg6LP1jLkCfnXWGdHt/Q7jcmuganlKBXFPNy
g0UI4MCJRIJmGNKcL9ndhCDYDpswlF9ZwXib9h6aSI9IDB4ge7TWm75j2ZQO
IpzBJVKsDTArI2O5bAIA8KsMJjqgmox32v8uRRTNM15QhVhwRF1NxbtP+Hk0
3IPs/cwSy5pwmR/itA5a3JhwmmHKdNJ4W35RQ9BoGToMWHki8zzzVRp+PK3S
zGXOyM4PtYGum6KgqMye2p+zIycXPhA1R4qsPJm/gkwt4S7m84euzeX0bae6
c/0FaBmaJiZPOUDdHHNfAbAcTIKW895BRnQBgWikWSidI2N0yOx9d7CtRp3/
YrHdDK0vr17BOuXsfVc97j0zlVRcSJiKSEcBX3ZG+OD0imZVNxMdsQXiD/uZ
lr97EQJQGp5cMUt2cL7eJbYXq5RZK3Ov1Uxo+EOrqXXWNSgMhRytIm+6MKL0
QXmw/D8A6+p5T+cX1SPdvbXnH9l4563capFXDCA9Q6A0cWxWiKpBTe0oktAw
nbhbHVZ847HlG/xFlf2tVQjrg8/t7dLm91dCAyV6HyAXBUq0AIVHxyF3DdO7
qRsxAkyWQqjG0ifZBZCAmD+t6z6L/MQ1K1nZmaqIBEuzktLQYz3xWCj1Fad3
/VgVbM4cPBMejzXnkqRvQNKQbJdPFtZ1ZPuJ/fakOuPVJD8YNT+zJZB8YOZe
B7j5/F9e40/RkGM474zChFr+lGdkV8IoxdvEjv2xiOdEZzHQsATTT0dUEI8n
AddVUfQjlSOe2yegH1QvUzeEmXTMNLRtGD5+IOPRfZn6S1AWjDe4f1JPr86H
4Y9SvuVs5c7Xu9THgII7yPFHdEQL+4UPtmbWJe9wnUc4Xgn0LzdOMLI/RD3W
yLeAuf88V15P6aiM5y21C3vnkwuTtUHTTNFpMQrC91mtu5I92wwWR2kOszEr
H+AE6x2/8hKFgk7oOLeqkSO2E8aHapMReIJ72umYJ2gvFEMahev/otRasJRf
AHDzZwwUom4ESTjJKNZuRPKg5VyenrnfXjPmbK/ecyEFT9Gi27xVvv9JQ9f9
L2lE4nA4CUFM+94GWlJxGGNMTE0tAzsVxciF/Y8SNk+kMJpV0UOM2EF8rCcF
uo9jtTcDzS6iSr7MCWaNMl5qxUNlft8LBSP1Plk6LH/aI+zU9l/l10wn2trs
qrNlnfvZkjQdMfZZCN4uz4sdILv32TDYJTgY80IjrnD8EQlUOw6klUg4aGXK
K+CVJI0quEZnxccWrAJwUKIcGgNs/snKRPW/yqSrtPAxe53coACge/QXuk5K
/U7MMcxoDmAYLOPc90+WxV2mm7yiec6GfwtdK68NpjrLnrzYH7nT0KcDawme
JbmD4dTzYk8TjuIXVRVZdZICm0b4N7y872Bwme9J+T30NAa2Iab5OH0kny9g
1NjOvMQNO24DP+cXWQ3dE38Mm+KSJ9OCBfvwzfhG34oNLMX7r0wKYU6ZUxTF
xSIXtH6J8AM3f0wkP7TXCzxdgWVlO/sGe+9tMOyKjk5MjCrI1Oak4YFEGevv
quS3MTfLiZ3y6fSP2vFwa0JZ1OTLfLy7dHWtyqjQ9ubVFO86WcbZrSyR99mD
SXwI2PNpFlimsxuiQI8MyPHfe6jRqPEaISND+SGEzP/I61g/64qrFz8BZKyJ
qmkuIcZ6LNwva+CU9jWNrNNeiBX1NVYutmGxE0YFf9NfyB/uUmuSNrYTLJMb
n8kqUjqnQCa/odue6jjZ0bfs82quuTwIbGALvVFC4JgTvYG9SqxOz5NjNICF
2SXHQlCw6MFWgyzOdwa1uZ/bo/KEyY/ZW/OfSVFKjPbvefMF6mSrOPvBBn+E
pCiOeqU7qiNHwgGysbKvJfktbbm6mOnqTyEzNAhuzx0k24UEseqY3wJfJpwr
GIQgPtUMWuWUSPsFA91Kfvrg8tmfqzSr4tIX5RNERHt7PtXu6hJrWY3G+mxy
Qv2JCOlX8r6e1v9JEibdc5qzqR2NVfzOk10f5+g4A2uJI1U8lW9T8D0ZpPEp
WDpGd/+EHW4vHDa1nUdfB26zZ6p1q4NT6Ww6sNRqp8J9Oq3q8hLtLUQ/rr4m
esAc+7bYZIwewqnxbKztUcUjAQDxy8SDtRcwunB9lNBgC2ZT1LhU0yU1dtvI
5waUi7l1VvQV09HeoP4TVvzvrh/RjEaQGQRCl4WWTQ3PGQzzmyQNDG1dBVJX
ksiKR/Yf8z3ec5s8GtOo6Pj2Jfs8VT4f4KaojBrOy63RA6ZLM+TYyLIXNoZs
o0UHksfOy+u6F69rdqrcI5AE4n+gJ1byl/cPexedsRk2uS0jtjIxnaCwFZi9
aXYTVgPcMqUjmi5fmhrGgWjqwgUsLKdUQ6j29A3VhOz+VM+B2wCD+P2hEMag
gekTqgGJbM16/KAOpiJTQpsh3YB9KHK03yqGMNTmj9W1qxFnw81XB3Dcfrio
bSM7W1aVnEr+hLd3PhlmH/Y6lEpk+Ib4zTUm7jni85cBot0GYgjsl2xktJMN
9fGFGV1ZrWnk9ryaYgyq8ejTHJ9IAYyiI9h2cEJx6qmPEQbMFNeFwSHY65Ci
Ja2/anU4GHT6PkFzIctE0XoyMmTRPLgBTg0ujD1v2S7qyGGMz+82VNrj3mC7
KBkLHwZUHWyjwsJcJUyVXTIfENbIljT0Q43bCv5bYoJuA1RNKZ4d0xe2HI06
CnNFSLZfmQL4TJXMJxU81z6SQCMLClrHeOkax+DvlALjuONMb90x0ZlQfVFk
WAa6gM8Z5huitWGLDCsmBIECJwwNq8W4aCv0uxzFocpIC3m7tbaD5CD69eSg
Tvb0Q9UXgpias/yk71MVaLNA01pMCee8/DpyTfNCkRrghXSrBkYzcn1I63PY
oIQ0Ob9jlznB1FH8LN865mOVvZ5Z0uVLsfu5R14LhHI48vB0dn74zlP6DY8j
wFxwsAxFFs6n6rl7lRMauzcFvfJqYMPwdK1F9LLRGBstzcygYb3+t0nkEDxV
AzercG6g87VzvntHJAtxEMzri3elVzR4ar4rVU3JKr2y64zVyC92J3daXjLW
GsbklEorfhZ7Fr1JCP9gVZ+lBMGRlchhKZS9JOmm4Ln4lcva497wHdcJKdYf
Zbz+7BF5BBy2OMH/4AflSE+ZeMiWoLxWgr8gMj2KewImoCbA87hS+JVppudE
XwiPfeEZQ2iiH5psX5SAjI95NTg34bcrQiHn+VWMbIgs3Eg98h+v2D+DlryY
neZT8lvWGIc92Wavu+6EgfnDsu11PosE0ZYD1UdQcWuwhtmOXgVIhr5dmwlr
iz+HXv9DiTj4H43IFiVR6dsXIru4Ebp6huvmZ97UEB/CdPQcokEARycqPors
mlR+KSmdJ+C9H2g74MP+GsTeJ41AK5I+nSZ5yzsHBBgcpJ5zlwi0mkHajZoY
Qv5KpqnOgCrvwBvKR2MO7nALqv33scWLpZ9yiSSt0HCZnwGqw4+BINM8YYVu
0rB3WuHf2qnT94v8rKo1n3GqCjtgMMLKB0vR8WgAVckYZxj1cKCswiGlqz6g
8JdNmtBn7EQyfRv4atyfXEsvxn8gh0yPJffIeCb+DmZxKcJJNvOefQJ5/fFG
yl9dK72ZUVmorm24HxiaQpSf7kiLNhDbTMK5UuSE0a+RWKroNU/Wa3h+rt8J
Gw3ej3Lm/us8zVDWqMYOVRGoiSl3vSiArCp+GDsywYid9KXKYuZvBCIrh0tm
Apjzu3rfNolf2Gn5yteXDS2qTp8UcZ1aOEaBcUebpiZf6NkuxfMDWOWW2STS
k3nMroGe4Jxe9NspumaZjxryW9cZX5SQkaIq5e8kKo7UCSlHWEB2NGs636WU
jz/bJVUGizkyoZwnO0JY86WzpjFExZM3uxQDkWtrf1Skzn3nucZ1+9N0+zow
6cD1CYWpuXZaZOtrnbwe9A5ygPaMcQ/AkUUA8TzIdTvimtDuLN722xPiNNGf
0l/31yDZHLNQA9C6C0B40ciUBDIYfnStRUW292LXsr+9D6rMoLD+7M610EuV
1wmRhbHKCKCEeuzkrR6/FFnA3qTnbQ4qHGjdy1fZ+MZ+j6ldIThsgT4D4BU9
dnhIZC/FrhxePQQLz93+1qZDYIVD4ukNANbRU5Cmn3qpbzU2Yqz2bqAGNUEd
4GN0HPfDpSXv/eJKstiwR4u148BresLFVOhUXK1TUnbtAFggH/MDll/0MlSJ
sArrChKbrwHwIJlmmS3LlPBvrHeFYY6GWjaG6ix7IdF1ljN+w1KOXSCZB9HK
CTI07RfUG1xh7AYEyu/lrMnjrxbLcqOdSYs/k905qkJvtsOmEi+ktmHnag5q
CY9cabIBYHJoEXfs40Mz/tnxX8BEwjOb5fo+4Q8Fp85T8GIJgV2pUjZ3c2G+
1BRtMhoFfoWu4quC6iDMmIR5FBPvRXfeG1pBFJYD00T9leha+KFSRUjKbFf1
ODJGB3ANyzaaBG5bi4Hot9YWE1BBB9lO2zQ9GhY9gMtS3knAuG3RWFiJp8FF
7zpexi0/Ik/mcsYULmw64bU0Yh9lv1w1aDJr3nBn6eyNaWPvjeNcw6hZhSTa
8aynin82sEU5ep1w5FUCWsRfUuu5GiK8lvNBIMFhdenPdM78Y7ery2HzvwN8
qFTm0cHqYn4mXGcKfFQHWmVUwSx6RMACSq4+10fu7yjxF5AavNu3Boe8oIX+
pHGWYZvVoxL/o2b3MDM8xczCgb9XmYsfEyRKoJSYwrKJemK5tNfBvHtxA8XM
BqSw+NIfrnNqwZRLYK85REkFU9P+cqXTkQdlmr8aBF63PtkW/rAlsXp3W7Gu
BikgC0AJLePbRr1ZCNoc5nkWGGxgh+yb1GtpvEzeccl7FOchkBZdVPIDv+58
sY4c4NvwmZkGdg6k9FPwzGWUfEfd1yToLMMauUsYhinCdlIKYAzU5DjWh0Nc
K+8Khm1aw3kGIV8MpiTiBX02cV40c27c3Qut9EIpdjp4fO4SdkOuq9i/Kxyn
X0WWG+4dACiPlXO3IzNfgKCEkO+NV3q1ZtPW5MeHkSI7lBiDIW7op/2aOnrv
F09ew4XSpfpv+uepaOjKVOAvZJah8wT2cqEi0RDTx+6U84hhY1Ov0s7Mopz1
JiW0fJuWIb60AFRnEJNdh/Da4JVuR7fTptN3TwlRi5vMKgk0Nb4ABLmc07Fa
NWWokaHvfeh6YtZvYf2Wn8d+jBzdpRORv8Dncb4Zxk7gJUmCGPQduxOFcULb
hRf86MToIRcI3bzSh3Yp6UiczxT7GSaLvaaVfU4CDdwqH6mqOkwrcE8Tz9di
wqA+xkZYmFt3i+fVYPCBAwfmHf9bo1cGnMN83uOXsVqqmVnuxE5Ds/76z652
2o9gM5dWupXdhwsS5hPz/ulEu6WkNpbu+dJMDTyclOU/CamMXwKUJtQIajMe
xOM6456RD1LLgWuNMJ1Ew45yBVcryw3tD49h4TiKARi/z4MzL5vr+ymP7G2e
MwBM+/uA7lzsmUkxLzN1ZiSx20qvX2ZgWzWAmVuCX4PAYyTGX5zqxOHv9zdR
e63ygeB9kwNaKHMLvRGFRY/SgSK/K4/d83n+QpI6UNk0CCXhvOCAdNBCfccB
YtmRbAkxE2nNOYEVRBf+8YrAozhuVmlUNrMDBGFjaYwkg4//CgfIsltXYAJj
xQdny97uxL0hbuv6eDeWTmN77QQeVD73BR5sY7/YnNMSwohupNo/Q47H/5Eo
4uGEcnCP7p+sM8FFM3iuOIj0ivB+YjgDXIcfNdkhU4cJ25ZqWce1Rb32yUac
kFYUzhpcQtkXg17EDLyGD7b/sQUupCoDK8gBGI6Ba2+P9+kKKzFIzUtE051w
IUGf0sx0LwNfSNz3rCWRJ6vf84LYlIAigPs/lNKDb1JgGKYXsJpRyRgFqoI2
eON2oPudkuNwEe1+MqgVC94POKWQzhzuu5JgWn6kJfw9TE83uMO0mHS4TIqs
rvXhSCuCiAJ7T6eCvH7qaNA4eUnzDQmc7ybTE51Rmn5ryOns1YMSV8jaR4G6
q4Z64Hiv5ygi6S+0vYzYh32mBOqLPVfANaOSGq5GBTdHnt8bKNL9Cwg1oako
WUGVyaKdSbS8tryny3saomRoNeGw5PVSPPdSqXxzAtRee296+LcA+o34iRgt
BuQxCkfXao0f22szCH3/ZuPdpxlxHJiGGSg6ieXVAP9/C8hb0gpmnl38HK8P
dWjlSydKiVq9W8eCD0o2HrawrY2IRNgWCRVXtXPhmgk0kn2T7oEmpsOiGuUX
3IA2lgksr601uh5qBDhV2C4/JecYQZzLpigWnmmyqBrA2ui6iLtHWKllH1z5
mosXKKPrCss6fPGUspTpj2HEiyFXupm/Y4HTIg3+YzkCwbHb1AUr6gRfAUHc
10Q96i13qAPpKG+AniILIwV24UcJ6hyW4IDmG7GZOvDqQ/qE7QQj9OpARM+e
Pfw4md9gCMVe5/eFgNgcdGxosVTbtPqBRT4a7RYQloeADkwQN+lZ1O9v+wZU
0R6hsV9pd9/22N6e58eNZ0gEeuXVLZGFWhpP2c4Fl8t2pkHqutR3Ny3hWgdL
liqVt0QWIBSI9LgJ4mZU2bfa/69ojphEbS+WUT6/2qdUcAU6cDIP6Nx2hvuV
kIpPvxtnzIyR4ZQQXCLAH2ztgtT4JiyspdFp+cTF2+ZlW1qI5VkBg/qOLulQ
wID5hoOmiJ7xzs93nWHLovkpxEQLxRsCG4jOHu8N69BEpoHXTqBiiKQ1GW5u
D/GBRe/VX1AZz4lFqfJbnVg3ymt0L4uvgcYHSEyTkeZZlF/2yiXTW6HIeVmD
Dw1wP9Mh/PHyds/iAUOSXR+HNNVNLaOrYOnwugYcLtC2oHUP5fXG5BCN6qdo
Dx7mjK0oqzJS5sy52xuBn39B3u7S8291EWaJ5zKZyPbzXVjrn7r2AR+sV+N9
DxHV3DWtYVyH3w24yX0Lgoa9M6Y0C/UzGDquTBjdNaOXoyauLt+9yITkw70q
Kdd6KraCEb8wJOE4vuihKwo/IYy9dH7+hW9UbcFiRTezxHLaqhTKSpJbvocd
dlcZeSMbSxW5B4OXkt6xMWg+YhWdq8RqC8LB5KSv+6S3e2rDUgeAgAB4tznJ
j9mn1wCEMvMRMCYoUzxxjpeSR22yg0yHq51AIrubVKgXmEG25HfrI8DKD7bn
/f6G1eSI3SsZegbvJD9QrQ+irWch4QIMlvvXeeWopKVKnwBmHLR8G9aaMgcU
ewt7QqondIBrr4F1iZLeE8u1X5khbC3k4TrOTOl4moyU1oeXF0MHu9rGQDjJ
XxCVKpFfFQueYnILXnrBgEGtqbsn0TDO0hC5P87YgBPVnYmUgSFrsLAd2W8t
Q5WbWkdK7SKuXOxOCHIn4Mc0ngWBKFfMN4WuzP6ZH/tSJCWUjGKlW5u9FLM2
JuH/kBJ4kH7Zi4f/F2RZr0qbVm3KxILRLOtsAg0Iu6ndyg6MrBmn2v+3nR2n
t8iqA1vvqYRsLLvgyEe5a1T7o54bNbiq3XLShBtfX8X0g4St86m99L2S7RW6
9uc9ZddA0WS7Tn0UgrrA4Gw4pueDK/WR39iv495tQ6TRc2yuMcORdSkaRUO6
pIWxvieMN8kSlEJCIKsMXd73/d12ju9osbeud6Jd83Xc+UtGEIGnI/BsQ05z
UaTKx5kq79IvadRS5fkQ35rE5NZ3BEmcdiVg8HMZADlkKYp2KjK9wVpdsfX0
mzBtasGuczPZFsfbQtiamxsRarA9jSEznesULhXyHDM42Re3GPAVfOCQNw9Y
q3rNrQdGI6T4ZIjOInhbiv4/I7TyMtfGR8adDOaiR3EeTbhgEXn6d663/8Hj
rc9/tTUO+F5j/yY6pYUeBXTvAR4eJgOdimjpCQs4Ekpll3QPBgFp4UbzGMNc
OQUt+zaKaY0gl3CjwLtMmM77GhRDRn40iX50jy8amgwB+fEHTLQQoWQOhCGF
aCfNfgUXcRB8wqXj7Dhn9k7w8wNiyX/S4ldbB0AGB4hW/k3aBSsOdmlcNaeZ
eoxC0KZI02GfUZW0QxtWo0x5o6YFW++4sZNeWCuBuTW4PxeP4/qBX3b1lA4y
jOLLHTPTI2h/+umrbIpjglE7QbKruufkojXadjjlLTT3JNwnSsrkkBDhxgwj
DsoYBdbdr/hCZTcZkqAVTk2stMOCcIfGZU7P2P2WN2Vh8UW6TaoFxUEN4f6j
TyywlakM7Uw6Bum7JlAWTQgZ/7DuS0T05A361Bk9LpcCa01hi6Kn4wzm/XzE
ytVHOWUBsq6rm+Aypwesz/jQInoUUiGKeebJoWMoyaMBXzWEnIhDrB++/Qab
h6E5B1hRbo8x36ttoXVTHCmnoM5z+voSKCJZKXJxXoSQSBP/mnUtbDwYe3WI
2eCHMv7uZ9jsr3mYmEKr8pKbwZBhm7I/RjHJMGQq+UFMttXSN0ULDdHXWI2c
aBqyNslyuS1LVP38ENZAqbzu3mzS3kbi6U9xzyZzS96nQ089isf0HwTkqKN2
EJ48qTR73w9q7z3Iv75qB8zW0vSrlhFXUgcTppCxEu9HEaSYvY0YxF9d5G0E
ci0rDeerTbxoc60guzJJ37Io+hJ9tebWh01oeJ+4JadaF9UxGPZpKzIq4n/u
oQ5LXayHTccrOttl+x7/mktZvrkNpf7oh573bMxQpMjaLTnnsCGYpTS4Xkuk
toGtL8yjZyqZyZsg6zgnLgyE4HRl4oushWuFWr/toXs5RfIIQdp1RFSd20hF
i+I0fsBJs09MhWhAicnZ0w1vt5Pr8mH4tJU2bVQH0RfvMZnprTXDEvEk+/Kp
+iDt+mgVuk1eQ5r90xJsmz2cqgVm4zD7QcCQYHYHUAbj/RrBC5MzFDLmsg2Y
+9ZqlEuH6bi+JBGlniWEmd9ViDSbfYSI8Xkg5jsNblXUcuG3V1uCKK4edXTY
hn3m3fFBiUq8D6df6GjZJQsEb2OAbKih1yu7kbFv7hd1Dro55IIsuIWlzt1F
X2X1MDZFkoxOLzs9LpgB39Y5duf2Yw+LXy1o5GR9DC29DtmlVodErHGrJc0H
/1c1K+2LAwBtazcNmVdz2nqvq6g+fBHkYpHQAHvKe1kxXyJcXnei24kYAngt
Wskr9JneWjAM9ML1szuzb6vAR4hq1wOZROtrt2GzqXspmKqLk3JjbqYHZplO
PdeXrZBcQjd3JXzAlRYBmLM1T3bb1FDbyT2bqtzwD/idSMx5LOa2nS+rJsdy
xTvczstIvKuub7mVAR9pdXaglfvuHu/aK9L3+kbGoXZeLXLUaMSKqM8kMprf
H7rG1Qhfyv6KGxbuoD9eAlsF0Ab8cW2o/1rweLTvQOoyeRAzKznFsqSva6DR
VdN7gBzYSFhPeo8ckGE3Gn5xOLgjmUuk3760YB1bbth2OABF2bfYFqn+S38f
v5ThAlSVmH9vSotFGMyXqSzhSOG14M+GGlpeUrO77Z7sWl0/vhIYHsQE1ejW
veBr2J6mUKa45dWQ205/BCiAC5timFjsyZJmW4/+NHJ9R4PVDOTqgAVOH/cH
U6yZNO0RxI0uMlXGWKouCLP+IA5aSr/VAFTKWDZtdXlddP+t/dzZnJejVeg0
cQgLfdmwUClTEKeogDSLW1NV8nxjwN+i2SLkpxXP/Vng1DCcdDNMtLXeymYw
ZM5iXpYKe7udTnPrr0/Pk5u1Pr6Nk07OJx4gR6W7OzfGHzyGBduKF/UiV8gh
c365eAVJJWwn2i9ZCYQSvyixYfgWxqSPp9FGTV1heKQ1M5Y0E4NATLfXPJnd
NJbVfulWfMzQG9OHKQ9qQmTn8Pj78OqydCCvTxzFmdl560soEVUTuEZcLwDb
bFLmkHkDw+9+Jnx7I5xorHTHUCsvRttM13wQ4ZWDoYXqFLOMD5xT2QWZIpOB
vicGj4PZK+1mVy2nVt/uswg3WsNwsfQ63VId4DBrSCM1RapDo1RmSavLya7z
OuPPuo6ulLjTeb7pW2euCVQ5YEd7sD5+OCGShBAIWpy2r1AacRmtMkemU1Xm
D/m5Un/Ws8cZD4vGcR33IXR8BJodXB3uNZFcnQa+VaFR/DLLxg/sZWPbnh6a
M5BRK3j8cEIusqe0SezwHOF+ZcVgUF1tnvhT95oe8wfzLm7psof5mJT4HxgD
R3xU8rZh7l0MOj863jVsyOIsPcZlNETVsN6+RVzU95sOE0GEs6E2eryp1Yqp
ohYwDnI74VFjXtxJ1bbvACDGR00CYcbdthMhwDHRoIM9pnuOCA+y4iPIdXve
I/+0fdlSEU7BM6TRPvDQNI1ofp2UYbyZDsNCR27nR+uAFPnmBaEHX/1epABy
/Z40uyhSN3Spa/7iJnz9or2vEgJFaUKF33kjm2U6HdFnkLHx7YwjfbzCoAc4
7cIaOVrCQZt4aXqE9o9F3PlgoQbC8yJZklUYfCpgl/j9KafKtJUzdZebCYn3
YIOIu4yUgEr8I/l+pXT1FHXt4vGKvJx4CRQyrwUmlHkzcdgutCB4w5wLjgqw
+hdJtDSz+g9QtiDg28W2C1HPSUs5cOHzQewhjFLmTL7pwu8yvEBJ8mDjgSju
7fUTGm4nCJoAeV/zaRU7YGm1tl2zDe6gdx7NVf6T71HYxhhw6LmN9cmQB5pG
lDu8KuKwdZwuzOqYwn96L8ClYJJAvCHIJAFZYv3DfcjYpHsIC+9e1W0hmSQl
wNC7pXT3kUHxsHxvorgPVKn2vp5J+MVDAhxbs4xZFmvmOZewXTo+UanxSDaD
DipaPFQLNm1iV7JNbs4tUoWmqMMzkYC/SlRkHCEYJc65FLbnUmXvqSyf4Ba2
p60MfdaSdtsObX3L89xnX18/nx3eo+ZhZxq5p77q6frESGu1GQ7rwbPsPERE
E0K+uswIjkI+9QjZRj84kYI7KYhaJQbbqzPUXhK9FLrFO12iVA9aYCtZiaIr
OuQIJtd7jlPse/CAIZgxIhNBi1SQK+EvM/OkzH5BtRV/0F8buOr44s5Zark5
y3/ad4/SrQcJGAcV7sAKYTdI4xk6yGhffzH8qePjLcIhWT0pMg5EVZtmbLCd
BhU7Dn5Iw1cTavAMWXCEo8dCgmI4psSb3cTNP6uEKerS0uPKLeadwnMEQbQB
M8/Lyj1TcwYwBaKbXLUMXszTsILYfEhxx67r2TU552M1WIJShvysBu8ePKWB
rBn/EbOjJNxdOKdLdCBq4Ar0hjwr/xd/KQvqNdYNKvHdoikmo34+ANgldqOj
o7ya/Z+qHWx5X9OtK0nxjDDVXOj8oeQwvEyYz3679ojaOv1nH54iCYQBBcDP
5rgDmavkr0H/uzyf4JphunYbdJeAHSdKQ/qGdakQKZkwE+tEHTTmnYy/I6Ib
i+qumL9ar030W605tME+cjN5DVTqOUG0BMNH9DV+EVxVhpuWezdv12eR59vu
YmFblMVR9WqseX+CyuDwLmKT2RAnpbiaZ/GX2Fdd+fqsP+WUmOT40yr0fiTt
wlIDQEXl9OPLlRlLOG3zroBet00BlDJKp/f3k0RvhtGXCYP4J2KOxEhwKsg9
mbv910G9BNUqG6zh4jj4BfnUr/GzO4/p43vo/flti1PxGrdxGAOB1Oe/Vqif
xtLUgF1/vE7zq+ZpIch4sP8n02vAiymO/4J/NyawczcN6+szmlKiD4deYb3O
Rg5q+A2INVjTdy9ZpiiYHTEWVVh01rARh5kAB+dz21Ty9zOZc1U0U8sS5QY5
UmrZ9Zpx6J2QShxtQh/G3hMJiIQEPsq1Y3LrKuWnXTqaou733Ygx0YMduFWZ
b6hIJLXqXLdq/rJzHL2ldnpd1BYg2hAH6fuI9jDFvJ/jOtG9Zn7huP8yTUN6
5tXgnGby1a4kYUnBlLZl+jKuKzTxpvyBbq7N2bsVmEoOxPSzDFj6NuZbn3VP
CINwj+HkZsptBuh5iNAhhIymBA5X+vOTw1ogNDS3VFuU13DVHX/1fqfE7L1E
XTtO21Dx3S/P9wIJ2cF1lLA/b6qsTv0iEnfN+afLqb8ZRvW06mRRluRMNEel
RNiwzAlga9F3jNskXWiOeSdCKGXDkwSW6sAKIWdkA6Pj3QgPZtVda7oi3odX
MnCHbuXDxpxEMGHXAmondIItZXrSO98lEuh6bKaUrakCGLzUCxDJUDn+VhBb
xdCT+jiZ/qmzeDeUcqtqOJ41gwiXYJMRVYbsmOaSN0fj+eb7YOGn/SaZiFjQ
z2Yjc/DFKE1XIWYSKeFpSmp8oyBRPik7IOeVfZTJHAc+8Tiopt83BR/+xpsp
q0bJ8w+tuEyXxPBDXf11ZjOlFseQBTTcD7LghfPmKOH5Pi05iHEzP0+46QtP
js6tNlnH9cUAq48mddNxzBc/vLzXTc51WA3MV97Ko86WLmFwSMu1bamDRR2o
Mu4yO8HzO1rLfoVXZXBWo7dIZ/G33wpyqKsLupT2C3C3AXOaiv0Vfd2qM86e
3/57w6QkQAqG836+0VlZ3kqsCSDpSh8ihwkL9CmhV/bEi3IPMDfTyJQk13m3
j+q/r7oyaLQgmL+NWBTggHx62cpSUvzEYp7Dtin39uqYD8KmQkUmwgx2GJb5
V8Sr3OGVFPw/mGZpPBuXgzcwlzrSc4HbCYVLclBnHMqFnCNIy5vfp/kQl5WH
DatqBCEl5GU4c00EwwW7UWqhCktWJJ1FP9zafXfnJdah1irYI+vzksi7MHzI
OjThq0+HVqVF3Pv4tr+P+KFnzzmshREnZSiy6n2eilMwaKZxAjl7qDw+77Wz
ZYTRu9G0rvWXiGiIAPaB0sfsEmoeXSeQ8uoLzrcwkDlTaythWl2moB6V7hPD
DeubXTGK2z1kOogKLwzQSXSaPfzE3o+IHBcnWufTKnVl+RuB4/ur+L+xdIOG
x9iLg6jgPnGvVIoW/RKNiEy/YAeqh9tOvOyY9ZNRaFQqRoE13WoVwWol+Qur
RvJrbZKYBU5isTKb44sEI6+QnuSteYYSNyLFDqokvUhqHlcKybPaiFhnOlJU
27ymDzOKJBt0SQCvAZmwFtp+YZ/7lyEnYLxASYdBQ97GuI8uN2zHd6vMCbRR
kgxsY0UgxMf5kgAxEhLiQWw6U/NOlv2psuW+SbhP7Hsw3Ae6j2ikvRVch/eU
elqmciv9bshk4SSu9ONM0MAq61t/7qu0q/eMrwWe+PuTMhR2xa39nXHTwkBj
44twP6zkSJQD+M/HpNdh+9iywrTWtvj9XGffshNjae73Wd8DEHH0nxQJxLCL
Fsi36fa85BzxbFMzPUaxIxXUZUwwNKihqYpRL5wxNte/WZTN3RbolijG1Gfo
c1JcHLq4WoCOpCpF7Lbl4dB7NHjD9d9x25TENYm7a4vt5gUT/OGU2C2Q+Jet
OjWKClZhuzE3FbDjLNgek9ULoFp08/1utbNOquQf9yIHS2ZXGE06hRHPToZB
9BF0PCY5GBo63IlBaEVXoorpvOOLXm17DZbjHsEwepvSWb9sh/du++JpOBv6
8Ii7ZWV+06MyLF+1zGWpsnj6AbNOwXknLhIBPPy3AvV01Fxkcbycf24nDG4u
kL8U5SZfT8rV2lWg4Em1HZ4ZJ2DvTAk6aBUf5Dahhz9FasdGK7G9kaGgaF8u
YhriM+wfqKRJOaJ2OpUij839f2pqB9Y5q9zPPbncJznIPgREJMRB53xGtu2O
VJUOYWJlZtr9hwnU39xlX+JYB5wwQqdIN5TnOxfzSUmsY4HF+PweqQWV7NQ0
/NOfqUy8dbEI991O4Bl05mcR8NuyfdCIEACIbSzPlYmWRVJjRsPwmmR4D17t
9UFNWE8c7mMZ5XFWqGkrt7NWL/Zyw97UUIUz3Aj7BCQ8u5gM0Umb6f2E3h7f
FAzTPk7/e2ftrW87oFGlb6abkeRnWV0J3W8DGKHxnKmvb70ddCzH//bklsSU
26CSflOAD3EaUAv9hn7bKXOFDHXnGiSNh8gSQQMwS2BPIGmYRkzDI+NNKznR
zV9K7Wxk7Sh7Ap8i/pvuPb/vQLr7hGn9p29ytPd8hbXEmoec4hdD/eyiJv4k
ZD618Cx6ietMnFQNBvQwBP/NXZj2GC+wybwRFo9Xa709LVN02aIPde5sCFdL
m8mXtA4BYqtQaxNovbwsOv04poHaq62CZM32FqThi1Uo1ccru5cHZv6HEoX1
7RWgwL5JsMhUrIbg/Effw5b/rbAZCbXpvJzxVl8ocaS0pSRyXgmIUKNANOQK
K1sCOaH24CP4pZaPXTOIV1H4KVMPz6leVwpz43NJyyqwwZWsq9Okr86OUbFw
40S4TsM8LOhqgx1H3etkynYCh+U5OOgWFOA3/mAZ584CtV7foGtCGA1yT/ym
5DRgELm/VpYWiWkwXujxzCkFbK6FfZzbQxBzTlSthpIuk5Tw+AevJdu0Mnhk
ExzrtHDka+E9nerdBxUM5z830DIdDmLTtscynxfkuHBv6uylnNKj1PoCzWBr
P79Oc6NQnFO/rsHY9Pf/5l1Hxo82btW7yroONPrxDgYXvyac8zOpth4BTM0J
CbtzV2cdEyKWwAEqppO8xQoLVenAFOimrRT8J1JcVdsxHV8z2F8YbKT5U79L
5g3ecdOFBu8yZARQMkLDeZ+AsAHkRZN0Fx1Te04jS4O6nsiT663UCjbhQ0vi
8sKXWkqQO2tJAGPfBkSxHe/VlG+zSYYpivngcQkyN9lbA5RgjzJkBY5yKfiY
BHtmYgEjBXJIHFspK8H+HFsl3d0pvxQl7zWEoMI3STv2kVsWfbvCdi3ObThR
/cGMnMBPJB8eox83kKWPdS509EnYGyWsjaQMf4/Mft74NyFAl4UmQ8Qwn+6v
c7v+ohhjVGtfcs0qpjv8nz36jl8qbisyewq4B4uQYqrCTNieaSBZTacprAhx
6xUqeh53u7ISWs/DbYSFDNa7ep7Zb80qI/sSwfT4t5uTneRE3LCwAiLygNgQ
+FB0GJT6jfo4j58e6jHQ6veKQBDHt6NMcpBJyLBc16JGPqlM7qFpLfuojUb9
/ZHiIwEMIH3oDlotnYOfIsfmEkIYLKIxNISllmcsBcWVCHcO8u1gfznVs1JC
aWbpUiRCk2HWfHXSeUGTtC0fFSOVWN3BYWmVtWR6vF5eAF3zFapUdBu2rSiX
ydtlKCg6rI+W7VcXt9Z7NjLSSs895k3VrAR7yOhCERs2i7p+8wfbDt6XIVEX
wDvZ7qm297MbP04M3Nid13rSHx0HWCveBXujIeucd/JrDtNmvGbjfDGPDolb
dflkCAMGYl93c95EKS+TnUdkPKvN9yE6wsYB12lxrU4h86NJOVpidSA4clij
3lvEkmlqGC15/QgdfCA7ySnQSz2b5EPxqHYatRTTHn6AXy0e86s5ul5ED6O6
y6lB0d5FkP4+tcAkaMpfICzfB8HdaUFr/dMM2Ch1y8leIlVOEydYCalM/2wd
i7cAuGR7NakIRffSMaMZ2eXpk26UkxWg/LZZhU9xa+FuDpADloHpgyJ2D0Ex
FuUd2F5dlrZ92+ppWjwQz2uR+zXTwnJuXePgcT1IPDKmpRMk0+LPUpmmZfbE
rKI8F1ORLgz7vgHzPZqgCtDWWrvcmOWohkq/EKrTuoald2Bd0vW9aASaNSvg
m6J4tJEciBvQN4rflAcDbJUmZAONhFnd1nqLZmeBooME6ZsLgbGB8jpf2ugw
dlq+ZxFOGCxzOpk8MHjl+OoQpgJqhvIOHfAW5zGxC01ssemkX4+JmhLBdBkP
L9Dk408jlCHqTxzJAWzt+98yCj3/Aaje+lBSQ6W+m5UMz90MEdIagc9UEjvT
VDt3LKlQ/pCLOAGDH5EWWdlRH5NW4s97jMZzTq/Zsltrm1fbbfUEa5d+oogc
pz9jT3njQ6Uvf4ZnAbMSvbMAKgTMQBA19SrgVxyf8hNc+96WW6jsU+oN2fUh
COvursq8zNtdPhYqVPQxTDKsU5zlJCKV7yJr236Zbpv6PtlGHCe/7lAMfaH4
8l+Wol/vq7Mi8+oeV1ePMcH4tDCMPN5Spy1wYwgl8eiqBbNDQIysC5Py685p
+nXdyt7j4YPg89dmCeY/jY5VX+9FIr/txWJkASP/bjs3JFpauBrB5+lY9WOR
fy6uZtPH+BL3FjOHW+1KwFobYTrWb2bZGF2WSQw1q6cTHJmZGg+GL0l53jac
Mp+++mv503CTn+4I7RgVAJBBOKDsKpAFUehAvD/LGlPJlrK2MFN8ZX5mLqmI
i59dBRY4GqaTg5v2onasQUwCchbKEImUtGKlFqgECrBYuKjA7pD9S92S3wer
nB7Lo3txXk1SxIBsPUguA4sZJX957ObEUXVAJtC/Kf30MzforFN5VBBEbICa
1Vrto2DG2/4CGy2KinHPk/H8Oe7puX+zoxGLVh4WP8wHMgSXW6Ckghi6BPSV
jO/dNsI/9Jkf9W8shPjRa6vQ0yQaXGoQmRWRxZN8I/EPPgvfV66rmnRGmomS
8xhaXVf7XvkzRP8U9Oaa3p6a58V7WXEVavZ/2J/PUgh4mhFbTvpMQMXftKzf
49W0kuCm2BsAA5A1h137ndwpiN8KAPWBdRvX0I7msvt+P+Yd9aeMfPx2uAZU
hkkGSdtOcfImXYs9WZ6USLHr8PNNim1P+z62IMamKSctlSExc1AoIm0wDTC4
38mdRKwZ5OESuJIbvlKzHTSkpfI+90uks43kqnzNVwpIxYdHQRAxOdzfPOBD
FW7JxIV29bGGovmfRlIhzSLPJm4olOXgwM55AkyNbkRMCzCAZ1hsftF/2hlK
4uI2/qkxp49WIt7Iahef4Pmca9IcU249HuyODg0WqCcwkhyyCG7TWXiEpsEU
XKX0TcLwEqhdaOyquXOh+U1BueLc0teFksib+8WW/OQl9JxbA/tmuIPJci1I
izwolwqu7Roz0QTo87Nm6OmEhji7mQF7F8pSFuHn6XsMCxuEBjRT0f8pncOe
Xhdgrdc/a/qJz3aPql7vMmUstLJzPhQk4nFLwxYJrcaYJUaQp5oJG51HNcPx
EUcxlZ2TBMPNUYyYxccRq/NV9ag9+C5mU8UmtLIZUVXNtRSNxQl9X0Q1rD0k
2hukcUMOk6UEEOQN0fUOQXYP9VXQBkM5ljAyvujyl5QUN3thGSGuYiXRd2Mx
TPiorcIh/EFyYsAX7HoH3eYQjmI/5EV4H/0vrHjg73YeDMjsdPW97qwIZqjA
YKrj4p+kVgiEuPwzwJoZTTGf9zWmx9pvkBObbMoXvlF4L/F8UcAAghx3Tm+M
9kqDNYYCD/AkPX28DJRfAtd8z+afcKmwNtZn0P1DA1HyBMbjhrEVah9ybyI1
SFJWXMg73cRGe+Fw8/cF4pPnN1CwecD7T2Uze/Jk6BD7y+wHW+UXWnpY44uD
xI9/1ekAUqAsFVhtCVzozY38MlMEUQb3DWrdUL0YjSqguutoIugm8+H5v6TN
OcibVbNjeRowm07wHAS4n1TwtpTPNdJI6FvHDauiFvnRl2TQQUbi4hs5WyEP
c3HRnimApnsH6xppBiFWXdwayBj6z6lolz48aNoAAK8N1GG6gbtDVlRMEv9f
AurLgNYPXC0XxJzimA3A+Nf4+f9yzr6/FykPE1BBZURjqCzIEK/tg6rjpTMe
NCRHD5I3hRk/Va77hbzU73KvbXE2NsVHyLqbcRt+z1XoOF9Cp5iDKy4d1mhF
KPgN19332PlQZ7s+7z8ty6MsTVBKUc+iL6ZT1JOaFmi9QdtVc/z7OAkkQ9uS
SX3yvX+Wn04HZCInjhDj7Snt5WxX/0Xe5l5col/HdC8InnUrz9a0jCOPuM0S
Sh20Ci/1CIdnvxE0SA7YwSXyCaWTHAinUkULL0nDdfqtmjG2pUIBX1T6+r7h
nxLjUHM2/9/Z8Vvy04QPoQHxMfSnMfP1Y1TJXz79mGyiMJ6pgoD6MgFgRVtf
DV/dJNmR+Xt7JBi1AqTwiBBA6qX/04Aks6YU+67/mU6644NARoxWX+vFIfIo
RG5nyi+mjXyYcw9b2F96Puls5Vn83et2zIdn34ACnY1thdfoHrUSTJMuhba3
ceDCSvccvItjXGTDlW79LmzzKu2ohyQASm0AYdKx4VXazNrPFWuRhKhfvPuO
vcXLvT3YNTcxjbuBSNIMJTlt5l3r4itB1lJpn1Ar1544/HIQbKnIJZCslLXq
pZDBjwQfLCz82fT8xLkJq80cQioxwcVBbxC+wrqZKRaXfLQlliSw6M2Uwrzh
iBUFRmMGc+JNRoK8Ufvk9fGz6WBVm6g6jDhFPpZHpyThmtgRRVP5tHhWt0Rl
tO/L2sVp9mT1Dx5TjVyxeON6WwDcIl8VRsgJWchLn8IxVo7AU8tBofOEZWXK
HlXBqQA9cOVGdaKrs+BZaSDLVULcEvzmUlYzOKhO4P6VboAGSaRUm1bqYmDx
ty7IGNSxS9RiQzvb+kfSaMBHTlGfoqQNKKbcq4MAeIeYr1rLQxRGnCrFYibX
sRM3lTYdC8LfAt/hAQLf2KzCrfF1+xKv8Fw3C+8qADdpoHoRVgoP9+4+Ice5
PzFESYu4PQsuriiQLhJS4AxEausn/ltLBu6qj6Zphq6pTpYR9Nia9VmJ5a7e
tKYFEFwwbpOpaVjT6b7vlPNGk0UdpaB9fh77yAPKesRjCcnuds7U+WY95637
0/yRp7sRJo5rjcqmETLVcP/7hOkAdgUGUWZmimEQROCK+7/wb1MFR2HhJa3l
NoaknELjcYRvZxUJUdILKXwIhM1+WblPUIXNVOUNz2bvdE+TbkXnhQ8JbqDi
o3fZjQhsH5l3Ab34xp4BbS0HcI9c/8pfPXnMajk61EnqBVTzcAYsGXbi8+Bg
eCML3v24JO17bLUSFx2wUEpXSoeEHSJfRX9m5Hirmdl3H9EGpPzN3Wiljcjw
zwFRA8qvXZqIxcDykUN0aVO4QUSpCqh3k8/QUEvC/HgHjz0hKOobOmVWc2IP
Nq137LwJLo0N/ocE8S2Q3zCNd+dPgpiHSJWw08YCDgdYIcsw9tz0NfFRbURi
cCu/EefWiIYFLOGSC3NShqQ1wxlqvbGhuwkL0xaQhOuRnytkemO8fc/B5yFQ
rew4ew9HuViA9kuSOegDTvzcNeFccCAiSdg+Q62ubmT2D+49sKGdrYXNpFIk
tgMtUNNbV1nhvzWnPIWewDlGKM0HQQaIT8mzbQn9pEcTCz19PAS9QIgr3CD3
PC4bHq9FDBitUZidZHvFN5w/cRX4/cQjoqiWr3djhuUY+iGuapLWrZF+/nfq
10LXkoy4zfmQuXzWiPYUnuWbOt3/fTzksQpWISCJUb8zgIUqmxc5RlkPOlGq
iq3smqLJxb/Nw2QEqwLE17nVh+7lJIao/vPMZmKz22tzCwlRhUypZOnbqCwu
+4eOJxgwK+q10/DGcHdfJVWu6a+jhRoCsFXKbbDaPN/GPHjBkXxfxs/Qk0ne
wv0JJvYhMtkUbmUkPcgKRXb3GjxsuXXQoN5SZd5KcPS6xHgmaaCKARhLaaij
MrOtKwCB5TrxB+5+4gal3ripTrV9ZVAj+HKUKlVg3Ruc5SlCARsCa8cnIwgc
1L3COfRA3J1ixc4bENmlzLTFgQbKQEZAfVzjFk3eQ1kGoWXmASekgLA/t4b8
5xHlYhEc+1SsLpJTY2tVDWEe9SYZ3hmwA3ql5rWiBZDXuuPRe0Q0mET4glV2
NMlD+KkQ0O8URUAco6R/4zx9JRl0ynQCV5EmmtNVKla9lO7Dk22b5qfb2OPM
Fdf8W7QhjcL3p3NqTnUrahW5qdav1rGC01vypsMUqGIQcMU98OX4GBqEoJDc
3BiKPJ5fAvUF+J95YvANybL5bL+WMLrN5q+EEUI5F4xIYDpV42twPReNXqvY
Edn3xOjM4jwaS6z166dtu4jjHVZwD62R0mq4kTromrhlEG4fnJKrcenCBvvj
uRR26cWg2TkT1tB2g0MeRkW3MMK867sDG9AxwIqr+q8beOGqqnLII/np/PGK
akZVffBdIGorZPhbu7MbneiJ8E3hTElzEagv0Nzs4130SlthSEvGDlw+KYhU
YGxlkiR1h99bJ4cW3RuvwqFxkWkXHXTqpC5AiVG1q9tP/zBAn+IKiJDoWcKQ
4JwB9Vmd3FHwAbp4ciswOFT0k8KIsSFJeNeD3wi2n78vt0iGPZWLvIV9SaoN
tCRjI0xEsiNVlUPjPnETU9VlZuQS7aEs6PjH1nS3sJK5Gmmo7SHn8cpbh9ed
UrnGGQJB9TiWJGbiZLc5pp+P3ETeJM600+wkrfzQZ6jVswnUZ/bFFCrmuU2P
uM6y0a1fAlfnh8YfKXQJS81V+f2DDovUPXM20zG0fReY4R4ckjJruvD7A6I6
ECgrCzU/aZMfSm93dYmCIafBHqBS3g4e/gVOMRh8QTFbQzDs8fvLvwekXMah
D4N/s+Dprd0vR8CYSxOwprSwc92cICg8r4sskRn2yNRP6myIMF8p+7hLPsje
XxTzPQpiQR5g2cAuAgG1DrBmSMnlFIGcira7NlenmIb/FQuCzoLvWPgK0VMM
1yDnMU14mzJFekiHCXRlSTo/SuJGewqqCvsJnN+a45dsQ22YtoXdOr+NryoS
wbKS4rpULfWa4Tu/9zMphnsLzcFOediTbl0F6Tio44pz64azrdI6TYABdlyg
CVbZmxMrKUn45hQlfhkU5l3lbKBL0wotZwneoH4mjBAQuhpoFaslvF2xSlAH
ELgzT/axU70ThG3SPU/trfD4GxKqceUVpWjHLadMhvJpGdS0gZP6Sf16Rw28
hPvq0aq2JVYnsfdqYNzT+bv5tJU9qaJWfiECbdi2LTLoA+Vi1MLwijr3fhss
jywOlTpEsR8creWBkLD4uZp/5G7F2GDgtkuFZMw7aR+SJ8eUo9ACtNtI3EDT
nmduJ29gjd+radjli/wz9yutw2W/C0hqtwAUR42kGSZNrnyNA5Uagpiy2W+Y
I4sxPjp7VeU3jeSv6/JY+p/Qu347KSCpjNyTZS4Q5CKmcmYsyAIlkSI53lon
TwioFOkp+yQuhNXC0FPxAPpzf8LMbO5s0OcifNoZtB0ckCKTVOlaDFT/7z1I
Gjr3VVpGYeLMuuFG2DfXw2f/N2t/kULieHD9nNTqxoDK4DTpLTlntG5x+3gF
ylUlYJYdT170Tz11dMiwLsXQc200oL0pDDEQuGusxjR4jZnXzRf73MILlMTr
9uQQJaVIHq51zImNSRce2TezUUV4l8AZrOpd5tkgIvqYfRkrNKjAMXHiwSBd
6l/jj3JgSd+CbIQ7KeTDk5r9/BoBnCLySq3CbG4Mfj5RNJHx356uBoTRWtvJ
kMNObfmJniO/uOrnOFinHbtG0KsjotMwojs9la2wl4VUrdXYelvBaYBS5iNA
tKg8C+HkVHpwqoGotz51fix/yvB3FfL+irsJkcFqA3Hn0ivBPb/MW3BGT+18
Zd3x2HDaGVQfYJ1Fy/dlE8DpHAgOeR9mDqRPHFFTfBiHyHwRfQi60oCbWK18
mccHuuuafvzAMeId+eYXs8UTrm6Xl1N0zceAOF0l6HWrHBsbMZGZa0g1f0YT
ll6mRbMSZJ5we+TFbAARkGSkFz1nq/HwbhyKJ5jTUjYe74l9qEF/OjJegeCu
9jDYPX+Xpm45koWLcmh71k7KxKh622ei0mtuqa7F8cwOl2E3HUux0Wt+wpDL
xGcntXoiG2NCJh9nvBxOAMRiPZMR2f5CVpLbVqeolDr8f1NdRPm+1Mtw1o6O
vzN4rcxJ7qsWEZXZtuoi9XrvXLuTN/jvw50uIx0IxOJRYgacHGfZESTjXPVT
dyRkCgwtVmp8weAEXCpwbrUaLh2F3idO87WqkJhJXZrJYDms9DnC+Gt3dMIw
YGxxCFtatK5oN1pr6jZTkEpQ7mchEF7pDRNseBjAmDlsX81WzYy4lKr7MDZp
RiPWUaByJCs1su1WLAz2r+MtshTzAmzjt6QPceTOqsn32f3uHQUH2YmCW1TU
DJss229b79mzWLWatutvvO5DVOohkC+B4Xg/qFHjTDtc2pqKqXIp+6r5JI+J
FDAZtSYbryWuLUNDeQvNuIphhUx/kqouCgfSF3BACO/GiePomM8Q5buOYL0F
5H+NS8FeoiBr44vACFKDd4q6VdR7r40YB/44oGnAG4zMlhshSESmUf7J+rsm
4BT5vL3eslgZNGNksvqeBnO7k3pY2hB+M9Um04j8a2fSHfxAwQ7wKanNE6at
GbyDX2/aPkUhsGfGARsOGvtB4QVmAzAdnhcjaHzBOIZE52ruuSuTQS4wWdWh
sYTNRtD9Mu3bmR9Y378zMvJ04m4E3vAoQ7EVa44I38BQ15HDFIDi7RdTHbXP
sukKZgCpfanXLF/mLkGOjmcPhJ2C2BP+jruvPUmpGQIguEsrwrSGnpe/8E8t
tHbD+ldW/n/5OPs21ll3+WOBB03t1XmOmzOuDCNcYvndeekySGwZifb3p1h9
kQQ8ShSW41XdtgWyVrDtMOhVtkEpj59J8Qkl6ELe+75tzaN8mOJ/sESUH3zS
tC+fJog5YkIlU7ofuyHhB3Z0j1sIaV91htYwMvqVvy2cuoGseqe7KkLZplAu
/yICDuqcqZygLI/jaoTTWjjpDorm3PXU82rAsiwxaeuI4fJ+Fv3Uc2LqkhVM
W/aX0Atf1v+fYX1l7oj9SA4GUeQtN8g1/kBOosFYO5WjXCxTpH5krqOV+VKJ
BMdFgKql6NXZiQldTA1z34uKiGoiRIeqQ0TPQeAL5hRs+8BCGAtyS31Fp7A1
vF+wPviZ5/HoburPvuoy5YDVD/0iZvNT0SHaOadhEKO3/DeXDGvEuYPhrFcP
miP195Jj8mXhSl271r0EsZZR3cfoZguOzHrrVVqIgNDp8fJKyGZkFJgGpSAF
Yg0c8XDu1BDQC7+dUxfy67ND7meeGqxvWneTh7jFvHhBPSCR9tIV7gjWL0eo
FW5MvQtDsNEUumDWCwjjef/d5GCu7tS6/VhzlpFk5MIsPnUJaiVm9jKOx2fX
ow6TostwtCzCJ1I2x39EIW+z4l0gwr29/VaXV0Fp12J4d4j+icDHuLoiKTqX
6RVxcaWUfPh8/2vFgYVWchM5p34l7W9laJNe9E4wzWfIfJO8a6bu7a9GrUWg
+CH+CHvYgELWgoc3cVHo+4kqNj1cHA71neMbwcLvzLWLDExBWmbDzt3vDcyY
ThF3Vrj01QgDBRzVo3GydDahfunY6Gis9+cH7BaczePrcKeajNZHOD5JO4fz
zf/3WUt5i+23pznm3uEHYkxPtqae08uX0NTL6ETwnSrKWeZ1/5mwOMejoaUw
riyytrWJyvwbx5XcOjHImxeWRZ+/qpjr2C+rpP2RBc/VloACw0uDkD+lsRJS
5UCZffNeXuq+MA0WupxfYWIr8IdSRTXtTlz3e9QTgCMhYhoM8bjiGMA8Q48I
K5qqGv/W7VKTzEWNEWEQ6wE1wJE4SfT/CLpXr7JzQew+nbwZyiPnM+DaOppn
pQKa+P1W+URKNM7IouyC1zHydZK66ka4KSADGGOGPC5SdlB5IfjZi+YwuGKU
/aMxLv61rFS5BEYACTBwpsjcGtlbx2HHT8tHCL6DUm3KWyA6UnbI28yIPJcn
1KrsOnLI/nddsOngK0Cfp7kOjMO0WBFDOY5ktEIoiUDCg/YB38vv6oEckpI5
keGKEQM0szpYrlJ8UJYKoM1jRHR3J7uHpX2WBkT46O6RDVu+I6rMv8Fpn5Yu
1Mws6Z0VLRlIfaSPi7tLoc9Q/audbp2piAQw6Wiu/5BBLCu7cMA6hMCCokcH
hRII65+r/NA6j4lgQ7+etpl/PeooCyoqDeWmIV2UtejzMbL/ZLU921neiczs
qtky8zPDfdqcexUJoESU4WsPjqK0LNV1qXadBP9Xa28yt2mxCIQzhCSIBTvp
1nQM99bb41YGCsIwfPuBF+0Iad5DPn8LlUk52h8RQs7wlqc//I3XtWR8zcYI
PCGFLfMQd4B04lk+DT5oNdstGI/Vgu+kA36XIwIbQWn37oGyuhpANgZPEQpY
N9pJf59kGavY3b0mucW3FJA0CmuGf4DPOihuwzyeNlxBGO+7N9/7hjT6aYbB
AdQKA+LWfhfxrtJ+tPxOKn3hGDuNQ801AP6ju6g4T0PegAidWUUW4TfyWq/A
MQz9zYPSOFkwX24GnZol2R0DH7gaJk0vWXfuhDa+UfLWqNQv0PWiodnKvyY1
jOnFgSTndUOZzCLPdMRRnykZ3LLhtmguFRHCgigfbHVuL8/9w7oPJcZvWivQ
DZjY7ZfTbHfygBHb/57LmQM4yWgCEeLuuKxGQQSmUU18Y0PRA28Hvle2UxSc
ijKjmzSE9WiZdjTH8TJaLP1yurvcjvUMfaWoKihAKwqxWLIJ+ZoGaZH9clMV
L3I94P7ffzl+NrKkz3PxRTvRsK2n/2mrMEQ+yjjvvXHIHACulA1MtpK6cH+f
5xUMXSr93SQk+I/GqAukrfSYgbt9WZ+nSUoXfZUZnj53hR6D7bCbxRIyvFUx
wEwxe3RagsZyIOs9YV9aQ4jnYJEDmSnV4fKRXbX0GTDimVk6yS5gu9QeHwLL
GSW+HNjU5LRwwNOvJ9yOOa+nTIjiNvIvAJfD+xjro3t1654V1Dz8XLzleud9
lRNGIciMQ8lJeUBLvYlaHXYkwba6oDASqjqh9cjwiFaoq5Az4NEVRsAqM6Rj
UejnNg52loeToOqNIyiOhzwmIpgC5d4BonyrxPXtvNCBVPQSQ1jmxF4CKpQB
jz+0aWR+IdqFYiPqoth6ohv7Yc4adapU8UxQjAOYwwD9tMeMroJc+qRpL8S9
VQFubMYEfMj2TYqTTu2l5NxX1Un0Nq3VM+MgeK8RmhSFZxOaB72qd0Iw+Bcu
SbaOz/VCiD3izIvImNyc1MB4rg5JyMSFoAdlshxJ9Kk3YNIiI/u9/N8VB8SA
pTbUf2LxJYZboUa/zNSViAaeRm8xPxngK1NIifdbMxMhvEAQcP7Vvpmb9WEH
HPz8BTihOtXfROXbjJa9+8H3kNh9ByAjG2PSDd9YKi2KXrFLGUo84Pt4Hbue
NcoE7iVCIa3uKMsCW4KfAZ9omvhc9S9OOMQrpBjOb4DTFtNPcmozziCXS9GR
AHnL6n3hsiIQppoVuo5y6sog+mDd6B5g0xcEHwvd4L96T2xFedWjr1XMJCMA
WwakviDBDyLecQii1xvi0gJ2HjFxDZE3wIlEqiqSAD6zQcaGxbTh/Rmg/8an
JMfBYgr1PWQpUXJCFA0W+SwLSaTV78fZ1wGW1kUQoY4/mogsms5iiFkVyeHe
wVNyltV1debBJOmt1p491hL5ImHjVOIHLrVSpsyessnKcuJ3YZ4lrqq4+2ko
N8ryXnf6Xpi+F+PQlmbHD9fJ2IRYpd/TDHVeraFnOs34I7tqHtDB5v+0EWno
WxjYZNYpGyDwsvMw9LKXEh98D6kAkaJC5l5T5KLmBvjmnYbJ0gnf0CTksiTb
RNuGdYVlwA+V333vmMRtV8WH0sx8Ek1nob7+OPwQDpAIfn2kVMxSg/mt9zTr
GOMbpiAMEWanvFERe58ZSDoL1UQwA8jTCoZnzg2UZyTNHTIO2Zv4FC9KOjW9
CoS/JvQr2fvondt1QSXgcV+AxZG9nC6+1uefIsvdhkkWq2Y+ccobSH/CDfbe
iyf3kPi9BMgdLMtLF0FhTL7greXraZ4hxef/9vvJJiz2vtNfUl+ayvPdCTD/
iVm8U1ls12Z07acEKW/8A4LozKQHu3o7cHSgHTN7FUZUaB4CuGUcIX5kBrYr
5FlkrW2YGn9ik8+F8u4nENV92Mh+xMrCUtIJ1LC7a7uK+mMz4otuppBk9SQs
+1QzpXE9XSbsVWmok+JqG7jdykQiQIiBLkt5aCw3MIPjCNIln8i5xGGpJXMk
G8rEaJgS9LMFaR2bi/4Ih5DZYY1B/arBVHu5QnM4uePCXG3PyUHJY367qYGW
r++HVqmbyXtwHP2z/Xx5WXrNLRz2mi9W6zaoKJs+CxNB72M6roGP/TbBg2mC
doTE/VRWXGScYHamhZOfwXy1VIJH2/KbKIPA8emXmUuAFra4Ppnq5QoyhnHl
wCE9T2kiGnCn4LU54/5g7cQgg9F7/NMvVIqcVnrjYZ82CJ5feA4X7vqfWGZf
vVxss/16kZerJias2/tNZrNiEDJAKCuZENkXFlr12Vxq9zMvlhLj1WTnHJ1r
M60JbGCp7J/Psb+qyi1ZvkFdbJU03S4GuMI8l8pkQ5Lb29KRd/gSobfFITTX
Xp32l0YTIh2SlrI4000gJPy8AdXjDwouHyeAzJ/kRdLCYKCJQN7l44oo9Zra
dqTuhXT6ctumJkkYsT45g+hxLhJ74F0T7hvpV6XVjsDjuvYtVUVyrRt4b4KU
fzkiSLrPSx+MzatJuQboVX6ks7ZjaFl+0+4mu7UR0w7NzCqrqa8DZrkDYQN8
9WIyaobcRNUCkA86wIvMIi1gaJkzxWfhOEH1ukzEsSTLCzGrVbeofA3F24aI
+KdxTH/KWPsHOj4Gr/dfeEL+zSnaFzxJB6sIkraBoF0XZ+ixexB6ZXxpjTPt
P75wXIP7IfpUu2wRrK/vkK43qC+PIMjEJDRntjqMIBHZ0k3Wc7Z59+FFUVS2
8rbD/PXBkxx4SRfFlp2HajFFuniAeRsU1SawtnZHtBH3j1kfUf5L0hSkba2D
SYogWxikddK6lHwbI58M5Z2j+2o8nPPkTrcJ47ST17tUdba62fZNa1usC9f2
s6KBQOqbUb6WYK4X1Z6os0zNEBPe5ZS331MBqT8FHEiROiTEixGNR9Q5/k5r
z8r2q9WZrxlsDZ9lDWc+jU0q6Z7Rop1J8vdIaaJXfR/vqXSjj/XmObrNWuoS
ZCy+SKKSsyn4A/nJzvF3UTJuQzJunnXlZ5fLTUE85pjsijPsykQTcoIzIkaX
wG4RLKrkl4/GCKJMKMy6AX0qoxHl/UY46xNzPgeDtplauyamm5DqTlfdph43
t0MYIsmkQBZcrmvh5yWVdPc21tXNrMNanOhcV5XIWJK4y+WHsQzoEwKbc3AT
PEZlL+vpIomCbWPXhtGdlgE6f17bFis7AvRuYZEgFg+BQoR2+eZuUrTg8zdq
3AkNt/GvrUklzKOSdYwoPlSpdbybelH+vi7p0O69VztiGRujDHTPbLWaroft
DdCXPlPPpBQ5kX4HVw/ScYeRAW/qie/qT0BXSlb55pMdEWHQWz2ktkm0C14t
yyA0uslF/ZUJtxTInt42kPFaN58i3bUxrYFyVpX3uaIvnZ/78vMBha5LhW5a
V9W8oxw1mUwqLdz79ULh7mLfNlAoVBHzEMKC3LQ0KmKmPUN8czSEb+ar/Od9
KjtxUOtc8WsEED/dDp2OCyLq8SyHfUtJtFTfxObjeBe/lclOZLuVCIfcPfNJ
apW+xZXsuLa54ga7R1UITZzeOZq0mEIZ1zs/qsgsWSLzICGH87RFZ7Gj7d47
pFD9TmXRE3KgDQXSCf7Rk4zVNLPHqEjfJ2EdFWsNDniB0SdBVLDRtBZULpx6
Zkh4tGpcqNYc/BryIqKs2S82RnQZWLp2UwxxheeFW4GcpnDgv8uBA+SwaFjT
zJ7Y7QcyZGoYHgIkRqr4EVX+YuX0QNLJI1z1CVzMJC+anyDCZ5D9P4c7APn/
MGxwj6yfmwptQfWfv9ULeT1vikBClHpQprJpkzhsjO1FVG7U3PFf8VYRPJ9q
2GbqiPHa1Etl4s2f+2uEjxGO7zyrO/qMH5K/FBqwnrvO5ySJZpIF9eaqxaz0
asVndt/HukaXD2lKprV2MPFYxHWCu7uHnNGVysMpTU1uqxqumb6rsSjpQc7v
1RhlVLoN+Kqswe56xV1LaiDqNZfWNnIjbghTxrEi23+Xtnu//Fnb13vM3Rdh
2k9XW/IJpjI+XPWLSZauQg+tM3iNUpr52B/OMVDrQDKbWXLtt+XpdhAii/Hf
Ai83eCU/NJPwvMb6V6H8NQa0cu4gp59q79rkjvx2L20+TQKYv7SqWVHpHmqX
/8gcI2AC+U1uGs2G6YsiAB7L9kfAkihiQ8H3wyy+6Dl+/QnwQlT+5QFbDxOJ
0d+YBF9tgCpe2kbCdd7fvjLRDz354hrlAAoPzLfuiuu1z1P1VZ4/LIEqteSx
nkTLBmranuRVQjKihmAYwkws/YnR5mJqSZuuB8Rn4d0TglNkvwEs4JJG5Gb7
oMxGfm1ZgsMuBl5wPPT+tSAAWW45ZeflUtGEmmO+u11syL6Vujk3ptrE8ts+
GztqKE7D4iwfK0s7lUglv0TNPzRsrH0ding8ThFM4eG3bcBYfm0fvSRRdDdV
tgV5RqY1dct792CLWjCp8SPcysmxlVg6HwXucKcsLi09yRj0J59uJ+0gxogE
zY5jmIZrf0jw5gMnMru+gQrNbPSy0p/zXQN4KYFC+jeXX9GcVYlARYbkH8TF
rrerhTZrYqaMLm8d3+yHpePWGhp0DXbz+oTZg3IkpPyN0JZh+bM3khik8gsq
6UBREkjyOBIOTbysDJ7zWrNVKAve+IaUeTNiAE9XfhqxOUgF1ef4NaaaTVMH
dMFGB8d4vdRAvVIAB5NgxJ2NsJ8JhXvgWeHmG/tDxj8nytnYgpriyLjeyDG1
Sy4n/wuRbVvOUli+b/bZrpmLSUv9yy5pDsqG1c4Sw2UCum7F8gh/AKJ1Ye1T
nOznDhz1oIj9Q66SQor9z2k7IWMP2fDn0bGLsBP2qYVNR2YS+NpQyBM6rEeK
9/Xv27yxZjZU5HIob4O4JcawU8FGbhLz5tW4CbVJ6btDiSK2T7J1uZUup/+Q
T/lZVAHO+AJBivcFfgQJ/6X4xaTFxpusVMUt3pfGjiueGDnbHKvZnibBn52E
TW067yrC/Z5y+jPbgnCa4nW0b+LEdp+8n5ct56uXbcB95LRgrSZHv/2XFeF9
CfDoCiMGa9zIvYTVOLmVTf4JuG722Flg1LwkZrc0YgNvxIElnBJJT1kbHNxy
gNO7StAjlQd8A/kz3xfdg2qc6GFhZIEpcLPq6haRhoO5yhBTM7R7q0l/WshO
lzoQqxH/2EK2cN70k8/i07TVwQxY5yecDJ8adDFbsIux4Rfei0QCz/Ql5H49
lnEundsDbBjG1foGmOYNhYobJlDo3URWle2CzP9hSd+Exx+mQNywKpyapiAv
SyMn0+FdmGWtXv/v7TaY3/2ciZSQnTw/5DOlWlfU77DvWhu4bFEQ6mSAJirj
IJSJmfT6eNpyNVfYz3SNwrIPITrEFJgGndI8KVTCtIIwrf4U4IJOWCTEnuYe
ZGWTl6BVgsNtrjbQMycPQnoSwVRBZlGOpuUh5q85Z78Tz/ySGLI8cU1dKAq6
nLVJtfaGrYtFZ99eyB6S2k/f+RmAC81wLipB4Wr0HOfR9PMY6McgTpzWIVmq
orLJXq/JmU8/xS1gPM6ohmCsRGeu0gKDnS8RmYL9CZ/4qbUhoOH6f6hrFF1n
2t0WgKJRnCTwVjltoOiYUdgAplFP3fNr5kLVKiEz9Q1rBznkq3uNUl+zJ1gh
37WBdaUkht66pUHJdU6WjkHA5Wvz10bRoI5OTz2S9ZCcYbvMl7FaQ/qwZY5l
hnK8conum75ELkCRHUC9v+M56AmcvzHM76AWpdDfC6Vj1ykJQiXglTD4t0PX
ambwV2pYb3N3J+CHz9Zxq18OOqTXn+nkWJ/pp0PtNAN7DFtxrOhlvX0sIqEo
9SI6NTVSZLForAjYklc9/adQYU1fHV11C8bjB6XoWunx/2YQvQdBUEWRMDOI
3zdbyFUCY/DTQQDSDRjG656FxByxVe+af+SGQWN2jIqcpVw09XEMfRDgnm5r
ypuhKsbgCxA/N+NGJSysusagAwYNGkrhoCd8tIWcjNjkqv4HZxgpWIE0w3+r
ariISEX38rfoO0+68yg7A9K3qhaSOpVRVRmZaxAjAZlRdTqVOfXSlbHMdS4I
xDb5IMO4u4cCzqhVLKab5qftptfEkmFHNwFd0TRmPbf2b4AKuxwQMCFBBUWA
uSjlIE9It5Zo64mWJ4lP0zXirZ1qIHUFNqes4kd4Ce0r8J7DIiXrjK7z3Qxa
HgY1ogvq+wK/9bkv9HYrLnvJHPaaa/iOWmmQBtKW7NncdxyKFcbB11MvrERT
AIzteeW/cCgnjgzefKrJv4eDYkLdUsed8au73S2XGXovIfD0bBCdkOTKd4GC
wyOfiabDY4uwZGrWrX17u4Jcsli3N6uoXNVRMlGAUU9L5VmAG+MfzihGxno0
YOTwkpGgZx5ShCsviZ1D3ykIB4a7rhVhwoQSt3SE5ZjyFEDkEpfkV9sUbokm
CDUL7Oq7kCYP8ErX0hVxoDd907DeUB4jOpTVqrqIjflWg6vjBzyVEo9mRanB
cdOlBQL27mXTion7Mxq/Xz+QtilUeinoNIsS+eBnBB5ualX7S/b+euPd86L2
x+L8CRdxtAKpVwh4PXQLVwzJg2QgsvqMgzXypZeoXiBOB1EdQpcV3AIgzFHf
9gofc25UUsUd2b5Zzgrok77x8q9H/J/DGxNm1LjDqxaVfDmYnEcBQ6f9A++N
jtn0PhWFwhILJ7LMjuYkHqPTjTuEk/mAnovV1X4scKj6FOZ9UWMq9lQbV2YO
Dqm90P7R7MLWsVYv09eXCydT1KTUK2D4pVbtJvCXV1Z4ZOXSnsZJm+qtO/Kn
ux1H7G8Oi7SLklau2A+NxHLQ0n9eXgWQIaO2KL/YQ2TpkJY/oysClgP+7pIX
H5kRD3ytUzy5Y5GX8fFG6nSHJAWighp2Ucocr+suCyqVXw3Q7UKg4jmqQiM2
up90ISWggAtM6nDxC2AgaAXLKel4a7QCgGC6Z5fLoaQmAvyVf7AZMFEbkfw1
qoMpi0ojPcZJeCL65goqUirp9J0kpwaPIB0D8i3VIgqT9WiyoHrq8lcLFOFT
spgNL/Ml8t0gsLLMCzNYgN13GNcazoK5G/WBcrwv3Yd0HGq5O6/EF8iIiAN1
d+d1+TUYHIeK8R4QjcbHV9oxJakNrva40oHuxHS+v/ojJUa54Ln/DxX1YvWY
VtwRpB8jeKr/G9+rsH3hCtLcvUEDR3ELLlBYVAzgdeZVTbf7nZQcZU7dlBOT
lztWqeRF6mxPvlDNMPzSKBLsPk2DAi09aGWeEn9KJqXBkDgfbRvQJeU8MH/c
OrJI9pzmopm3vTN6PvIRFu3FUKRix9RCakTy3hpGa9SRD8/y00mBtHtatiBL
3sESwOFKg/RZAE/F9ZsYkTMABTLhj99ukJKLdXCMEsbsW05upv4ncTAKI4DU
f+NQ+CeLE4Lkz/38cvtN2qof/WTN1CAjL5tTN/uYN4tKKvj36F+9tWkrgBk+
YMHHyh4DPk+8+hDoHYO5+NyPSDugg0mmFhPEySY9qTwodakOhdOFWVoWKCJr
3rTjFjtPppeHD2mQt1wlWG52OWdC1TxkbjWeL8a/aKWUmlgrAIyhWYa2N04A
u5qlbplNc+tHDWI7zJ57t3Ejs0pooGOMW6sfgqrPyuEKBthhyzJ+uvjWIuTH
U92Z1GDmkFyY/zlS9zNTX4mwkx/sC5p7iqWUe0j2PmgGQKI2li8Z+NIbI5QO
/axVcnGjmE8czDg5STSneIeiHwHLYL9sKc8fv+8fHF9OnGkSU7kFHeRW0Q56
uyWZUTX+/UEhykpO6LbXJsSBif8djFLDh44wVFdPF3iKt+j5wgiYBVK5HGgI
j4Wl2GID913PXrmxYmCB74R+5UrGw8zQHtXbYvlVNMBNas6efKPC0qmLqSyF
uWIdjZMmbJwv41WoZslI9V8eVkZAydXtNwUe5LM1sOyx2JH/xLGBDQp9nr19
PDgmw3Q/2Uph26qyGIEXRcq6csOiFx8u5/kt7ibfethMWbP8ZRtx9RYocVy/
HRImOgDQqWud0bY5oC8EFSHCyG/9X64i2R2Zzyc/5LpT86YVliswA0yai+KJ
GBvcXY9VRjcdm/HUM/h7Zougdq339b5YvI4YjMIL2UG3/yP5TSeyVN7mg2ce
rAZLhTnHl+34BCVFUcTAxjdXNruNYd4uCDaktFDyMGa14/fQMKWzrEQes4kx
FWADaTGmZiT+qIWd3lCY486siOxnx8tD4mIedfXSCFjMyS+OiCOtuCZ2SOpU
1rgWaRErtd9E/pvmdtFtlSy7iDKDNw/lw729wfa+UqYb8M8ZJQaG58HLGLvR
ecxOyjmopLQhyhnvZhd0VJoDh6PonU71XXlJojvaldWEkoMaiHuKB0a+5mD/
VS+fjWskVqTriddFfp9cDKsojHEGlVqhlrJmsOUTgTlyzN5YzWJrnH5m6Xj2
6Pn3hgiDX0paOSA5RBD6uj4ovo6slF7UqzFhAjMQUFHsqIGmGvlD6QYK0t8i
s2JboDze52RY4R1hltDUaJSwuS3IBJRpJcLYaeLFrDeLtSiU6z/S532IY/6Q
c79DcJUFM06UC5jVeWQgRndd8m//BsdBSGBZLKkfjfS8urpZRN98+YPvn6PT
Gj5d3KMmfPcWtOmmgVCnILqYaocvaju19oja/QAoFPttocE9yfzM0PU01QAJ
REY6dzVWjM8fkWcmnDVfemAsh6yvmg56171t93EYqYcwmgPpM2qhaNrvLN2M
Nb4f+m5+63XJAtiPzUe4lqMW9GPeQSEThFsGq7TtiKAsd5cj3MVIPWrmWMal
a+v87XBex/MxYjT4GJPpQQxQRu9fYm1y28OzZLtBbobAIc3yFa8b9+gk/UQX
q0T1YwpaRSpVxHTGnjNEYw+njny2zVTx6fVg5f55x8No93rKe0650oBkmZQJ
ZT02hk2OkJAmQkINXcn0A+kxPBd31apHhoLIp6zJeYaBqOG48RSgvTqTbdww
fl/qBmmMNz/FqaVg7xLK4bvCqVgSvCtMWGzbDuHJSX+pNr4iGTzMJUi1rhGv
etvVsdpbTo9pyHwvvmuXl8V8do6n1vzFMJ+qV5gq6iIzn8t3TTK3jJ0btp7m
kLoEqgmh3ugTvl6PcNbcS6UmYMr+JzOkVHqjB4fDP1xH0KF09wJICj0LKk3T
XoMuDCZvOej09CZoBByGHeAg50ayK+ui5KYOGbJyaAQ/7ZtZVDxJUbTbbKwl
DCMaQhKLjy9sT1HPeAZj5OlnR1L/q56c/C2gOJRGB9A2W9sIHIoJWi1j/sZs
WvBtimgUGkFHS2JTp76VUfYXE/EK3PkhAr+523FV7gg4UWEeSNt2KloDeY1k
igBWqs5/EfO8jy5o43YUKtDuAHYMG+TZiDhMkihIQ8ZuQzsT8ycdvEzVVTyU
lOT0zZSb9FtSQOJ4hxmUkgwe6YM/iF31NYSczp1PIn46nBWnVr0ma2vWzhfm
DXg/JcmXXipeNQtvjLzAKQOg57rn1ZS+huOgtfTsO8qoDf7KtlwPLOVS2chV
FwrqRp/dYGZCxkMtfVm9RKhoE7ngQZM7wauzceIp7M9E93u8zCtM4wGk2DBA
jc5I/dee5Tca4a4BOuJWmf9C8QYWX+l/28zns3fuj5FxAdeuOzCdPos9pXs5
M1QorSGL7yAs6PqMmkmhssgU7JUVRZsttPBcGj5NCX6XDyARWax5JbBN2/2i
nAw6P4QmHSRyJoanSjewN6aOBONg/FtaRWyPSGfEp6o1UwK2DiUuLFhcvmvY
+aHx6JSMbSUQ55+jmUt7+wb7O/rRmnA6GTZeKVZVsr6t3XyfmwZjMOqXq82S
fOoIDHHC+kXH+w2CxGuu8qYcVMf+1IuMPw+siP8GcpCCiqNIgU1LISB8NRcD
oG0jhIjWB4BJO3mn5fsoVwYG22J31lluobCiAKr6RHEIrwUfp4bYduuWbT4j
UCY533WwQzAGgCaPp6LCDDcLaRdwefd4D6KtF08ic7hOYKwToDLzHf2t5+XA
Vs4OwqrD2uG3DBmAYZWz5UELeSb4fsTF0TMy4NrueMwYQI7GCxgyYPw7d6tA
JmehOqscaAui7FgbeNTtpnodtgAM8QWU864xf870F7EtRG5S5mHlPq/yVFfw
jRHtsu+LyA/ZvHu761kC7GRuUQvW90DVClhFBmjcQOtPzDy/M7y1b4aylYTU
66rJlJ91zs0UerSaLtliDOPLPWSi/dyBWZLFYmR1ZAeUi45ctnqy0TzgqDVd
aMu15kzMNqFhVwXWUtwdkOR2M+qxeFSw+9gZNWcIfDU7QmovqctMwvp+PJbW
J46m/NTmHkFYYyI6ifRJIszMfkmip7KWEJ6SdVXOVqfgdfs/M6802rJgedlW
b4qzcumDLt73v6j3eWqxnQGqXWPlPcoAlD6wkyLsCVeophBkBXZYCg1HV8Az
N/eV79pXyB9Zf8RGamzGrZR3ex3Yu6CJZ4FhGUA3XtzvvuXni94MyzEWcjIj
1dp1Lp/kIpFAE1JYB/iUBtnycWm6sRxnwTeK2wOsd6xn7zaXVQ3n4839nTc/
mBHukyopqnQAlpPGASMjPee7M4+ir9z23R2SSoKB6n1rJyZqZcFWCnaNuS6h
MrBDmn2X8yTzHwRCKdQGEU+aAkq0yiVrpEFlncgTXFUSey7rVaH07rQgncGc
VLPh6hnDfCDqXE0PCJyOYTZC6P5VtP8PJGKn9x0YJR5o1fnRQXarXPyMj3gA
IRk0mBf5k2TZFKvUhJqU/TsjPBzSIydbzl+WEVIcKZV9+dGvKwwMb1Ye/jqe
Ur6mNXO1tUWKxnrfmM4Lqng3WRzWM4Tnvz+o508QiVPxjvEU0Z8CQgt0/NL7
om9Lk8ADp8SEAh+MoULqzsy6ELr2rWT+YdMZpjUxAM/4AOYY026xIAUGuMI+
9R9Vl9NLfarZBeLEYpfUxkurpucjvaZK03SY4N6mwlS6Q8lmfSR/NjQUAFKc
CXwveCY4ZQmPTYYD18SKIBDGcKf44Fv9kUU4JSbCBWvRhxwohl3Tj8O+cGKO
I80t9a87unsuS1W6esOFMIvZZ4j7c3GDDy0nwiXgL2Ui5g+7nqm0VsXOE7sg
watRaXk1wL+7DoGuIkp+smSHKERtE6IzXAWYsvpUVndYkJqyE3+J5GtyNxpt
l2QuUqpsYkBrQVBT/r6utGI7W2cRzkPDT9HTQlJIhlnU0UPQMM5AgvJq911U
Dpf7U/Nu54lsjiMV7NVJTD0odP6PuNs76AgsNk9kIW0pYcHAehHetIwiFDD7
FPpzsB4hDWMAxl3w1AiTjZfc3vYzI2ZfnGGc5ctnIxGM6bCxBtAuVa0Juicl
5Kmuk4BGFtvX6MvaRr4JQGaWluLdGk0USAZ9/Lb/hvAWdgBcOcc5xWsialQM
cwEkpuwkcAc7XWnLzv7wFMsacPnsCSlC9N+V1lNm3Z8HEE2ovD9kDShvUzxP
bTpGQdRX82wwqaeh2L7iwVXFJvoRM6fApZuh0jPAXlvchdaB2cNt//3tqtvh
s2J07e3j/vrEZN2Hh3d1uZg01lyoT+9jspforylfSFwA7pYsN006r6PkE9J1
C6BCwMzVwXY44XoLpU9cCggyqwHfbHAjpcOjmh2+MAlGJMb0S8VGnLreR7va
K8Ic3g9ubBLnXuQjWpRIByfg1wRsVbDHA9wlC8TCqmnh16v+V0bIIK+3H+/d
0z4T3QWFLG9WuFytUqRZSUFOMeBEbz2iffHrPkMosJEbIQXmnzhO510nYLQz
Lj9+oIC4r0IKmdwELTu3YZ+cHz8cCV9d77belTrEIzyz6VFY2NYAOIu0kg5k
RvS24XkogWH7lHp2aX8It1mBYXfXbnFOM4HKrQuhjPR2FayV9ULeGUavCu0I
Kmw5ESUw3+Iu7cCRvNSUMn/yToC/4D1lQwNcaDuGMc3DMPLRnkPgJXybfN3y
2T5PzCwe3G1ATz3px9K9YmdwT6NwABgdxdD8RLp8Vtz4PfxP9ttIm8yGRHz1
YpFlLD+OWyCuMVLiryQU1oFpbFnXT56iQvuSrLvWHHKcQACy6RsU8qP474jb
1wZJVjwSm6cdhYMGoNpnpQKzw1F4wJKg6fkK4Bylxxpc71A2D3s1w3jFxh6E
dPwvYpTdD+FJViIOc9EHqGw8hY9EN3d7Pzl98rOGOJH5V3YJ5YNVoI/wDemA
NZJR6GOtJAedTZEK7yrSmBlc/yF1dpY9wTEGjDHZ3jFKn+e8ug1qdBgn6KjG
qn6uw/HOblc5t8RgMRDcGIAxa/s0L+luUsbzaydc1bBOk0T7VeWmjTrRU3fV
srghq3HiIuuNpttC50KvSZ0i4Ld5AizdREkUwni+wKBaIeiJ1b9skEco5gF5
E2VP15e7w4lshBRO09SMbASyNUgYclB/3eDdjEUcXKyyO6whBMJ+hnyExT2f
PAz2xvIWXHy4JrV6MYLwZYjUuGzn9YnpHI2CYylYpw5bFFpj9Sg9G9KucRzt
LdKzJPSSEqEatnjSUCL0h23OFE6tG6VdNpsBvPhTlJA2e2oGlrlfBeAZNKOZ
VxWPGW0zJox4b9Aw+46AF4bkFtZcmPz08I3Epv8o6MbIIVnVgB/VzxJowmhy
tGj+EimCQTgD8SQGIRrQoNyMIUAhYKB5hQ+eqWqyy2b44duRCDNzaSkU2Eul
bwSxGyt/0pgGjJZQAFvPyPjLzIA+Ng47vI7EjHWxVgjyI4eXhB3m6VuwfQzf
iQb8e8+j4PA6lUVmJDY2/6fsyge7XbyNwK0sMDTLUOuCj8SE9agKmG2R3v9E
mFt10/YzymUWf43QuuJLsr8Rxy1MAbgv3NEvvZ8tZM1D/R+cO2CabmRTnksk
yCLG8pqUDVXntuXxpB4vihqhJBw6KKYcI0txDWe+NnIq0WTolWPZ6RToGl7D
ZGWET73AT6fCmVvXmpCmXTQruiAXWiB5wSOnq1gU3mbPCjjc1Y4Nh4HXz3fp
SvXVau9+HcIpcBfolpgQ/xRaCWltC4ZvzNCfx8BygCPgiDPHL0VHwaBovzJi
WcgOMnwE+GYow/71EqtjrcQENclr1Cw3ZGmJPwdf/ay8vKPr8B5jiyw/rSn+
LKvFwIrAkPl1/wAPgAV38Y1efYhHrW3W6FY955SfcA25nJqc22KATbissTGf
ZpwU1MejJ+rXSxrsJP+bxeskl8BrSrCuUGD7zfibTPfD49rsBNyCVx8VoC3Q
hASFkeAWdma9U5+hcORulzMSHzfXDvyfIExrtiTf9jiUPU89EhpbqQv1QCF+
hmZU9TNTIIQ+3+kSpNddpDWgU/lqJqUpTN1ddsMy4Q8n7nzlSrAFPzNpo9iB
8vZDgkbaQ8+M872WGzDxm9RfhqxV47PM33SPis7pJcK+eNQxX8pjWty7zPRb
mPt//7kayiiLzGwqA0XVvefqCjwAevAKjKezBIrrtSuZUlDRLMrbRfFCZu18
B0ONoRjj58kXv93e0Gfj4dfhkv3z97WlHsEhDMNnCJy//2Gf69Ppr0OuMG8h
YJofNl5UgkPjsdm0A+qu6++yGPTycg+JcKRVkTL/ruXrgkVyo/bxW1Nq0zc8
8DltlMVPJDmkCGULmZwhsHxQiZR8DpAA15Wb/jzuFjekftHldw8Da5q2Sc/W
ssr5Xw3DvwY3Uem309wncNpfWqhsOICqOxXDsm8X3eUZx/unAm1eNElapkNB
rj65vqAqsLWiFdrvJcD0x94HHtBNEBJEQzd8bGxSTypQ8gumr6PjrEZoEjpu
XhtoNZlTWqE/gepd67pnNXQEE2ZXjzWYT0N0vD9JJc1cwUgNMcQnbtBjRpqK
DGGI5sSwRutjcMwqskJF445vX/hnI9mfJuFwkt9j48dw4u5fw9yaKrLl2MMJ
EPzo2sAL9GhTB3UICgV09gmf/lIEU3DJYv551axLD4/EG7hDq37Zj+HgfIEK
WrDwe8+eRnpw9aIhixTfRaSVgkwBXUuMevkGL0SrGVmeDfQmaBV5Zpa7khLS
iMimZuCOSmieJRHT0wMlLlcdC8jj/YNr91y06K8rg5RVX/5tU7sZPavmpqp6
zMkBukp8IFWFdUt6QxJTgEvqG8rEta5F4gwYSMry9N7ADnZSDd97kbnkmNcR
HNi8+Py6tQ4+UstdNpnADA5zTHsH73+g1qlGejP9eq6NowE7qsyonqsAZZaM
BOePx9Q3bWfoB3CIo+obIR+YTAXH0cX2CUaj+WLCm5wY0ylb+exU5GLQDoaO
oQZFPvDqLbBpKbAEqPNSznrREmXYrM0NMSO9qctFBoIfXYct/i0sJLIkNSCc
sqS3rcpfpM88P521ZAXjk6SFBQITlXy3dxM3yVhRKYGv7X8YgN4ydefOCT9P
gyeYQ9q9UEzolU5qRvfLo8gytgzzOFb5P9IB8/3Lfj1TZFb9iRizz0OEZD8m
4ZBM3nFQwvxw4XGwINAu9H+mHbDVdCUF89eFB2LckPs9zr9lweOnzY3kJB/D
lYt4HT+jrEb6T04Ol83SGlSnvpl+uieab4LVhpkF8uRcD3v+V2UPdtdnM452
XEld6Scw/qs8ENYlcyyt/aZxsQgtCaiVqL49zfQ/+1UpoQ6Vn/xgb0/eefyh
T+sTT+bU40w6Jij2GjAVQVp5yP2JPrLrLGvPxkr77EMHQxInlNi8vs6s4zAO
JBiZ30WFJirPdG88NTouYwoNzl7Z9/2Viuf64PQiccO/vXwW7DY3cVOXjggh
6NTA+bA0SsUjSuXlpHeAZfWQYknxgE4aL7G7eOpH6m+GT4X7XResmBcj2Vkk
fRQdxTgOM9b32o5KN7Ue+uwOHxvIiOfiYEsQv1gJaSqmN9iKyCgFlpC4uVGK
e4o9hsToNfVKeGm6/FvRvQMqsg62zmSFW4FtkEclDXZ8mPYokA6oxrHLgfDL
qZO+uvMuwkKZx2QvPWxV5WCBoqAKhm2BCufTu7UDPZj/lncLQDDlbLe5OZZX
RG2UmcS0Rp4sqx+JFTRTQEaK/AhlnQC/nEL3dDuP5sZTHjDsQjlvGWZdW8Mx
jiAiP3GQ/a9Wd6TGH+COMLC+gkrKAL7XiJ4Wwth+rgUnfHHMIe78wiMzy+kV
OsmeXBLRhE7o+CdNjfu+fo6lt/BQ/CvMK+4ZbA0g9ITnhEPBzA73FN7HK2fZ
0xRqng5ev030pDEEmeztI2468hdmC138nKiWOeV1LxFaLw+8x1WQ2UMPLfdz
q7eAwvdfZLyMsPbKwhF9CMar6X9OSdV8azwvn6+UOG7TpJelV5PUGIlrH2Fe
n/WV3cmgRD4/ud/ZpkT7jfuxE0mrTjsLeW2Nvw8xYGblPaifKbjn4E43Zsy+
bwawcEqNQk9J1AKWoh8wseMux/LS47uXynKQDHIULotU0q3spQrlqGOW0O3M
DCA1P5NBfhZMk53hW8rDx1cvusFuxUep4tOEYCJqTpU8rfH+FbNAFQ7bI2HI
jXelc3t+3JMhPbPiS/MSPTEGihyLefqIfrXH6qiAFWdYOrUFPXBJB2mZw10/
Upi0fPH9XvzoUUH7T7/qohs5jQETc11nC/mXa4yfr9BWIEjVNl3luUZ3JG9W
KOgtv+MrEtyKDdaWVtPnW1oU6Dtft6i1dMuMV8qFJtAaKQllW6Ogf8sTFHes
ao3WtHaIB1brRI1NNADNsuzTUqwcTj9KYZpuEia5qgdrHhseVfYnk8a9+wED
TJPmHUOq6VX4WxIa3Z3ZVlvTGRlSn2Vc939rgsdvZ3Fz4Hj/kaXqWbBNXR8+
Yv99IgkyMI6sbfDTVfnuaTi9QXR1unhVsHPelrGEqktEDZzf+7Kk69iUgQkZ
3tbppy1yLrr4U4huJsebXkHLwNAGhDJuFOzJfw0XcxD/aOomYeJ3nWWL94ei
M3ZHVZgXgMRHMLdzOVtRtJp9qATyWu9itTYRZacI/ET4oyOqRB7ZBeOdP+VS
ZNbsHWH4IkHVVJF5HRggZ8GvU6VANv6hJWNMcoWRHzCJqAUbdXCgg4G6we4j
OovvvIdyMr0Z8I2UZ95Jg+APHd6nanyVVKD24lm+kItFvutO8vbBaSx4e8+j
ree3QdU9LzF9movI1MldeXO9vt0neFmR2/H/dAlraSG36ztZF4GlCqMi7ssR
RHTTPuWPXHQY04HGTrP933ef0pFw0FyWn0DkiWyvX1RsmPEFqMMqGQpDtO49
esOZCIenh/76m8Cu+ETKQzf5Wgouw2Jhir57mtvjeVwmSkGWkyIB8ziW+pz/
keikXhtHVQ+FujFXhXMAoSwlyVe1aJwSGMpDvxZMx/bDV3GM26oeK19k1hUU
nsREoKP0VnSujicPFixTr9CThx9FYA3h5H5XU7IIgK9LXQ0H/s/gI+gjXyd2
LmfD7Tk0tCj7Jw4uUHjolXPDh4YZ+sa8cFBQOBTfpReonEqZjoJrXsTo28tZ
IuwQS7++yuOLibquveHy0oEBl+zX4aBLJjhBN/EmgEmKlHDcRrLbiK0Y8C17
gfov59DTeE7SGFV1rbbxGqWIYwjonFLORTJkJhYw0W3jEjKoTPwpxafUmXmC
Ib1wFLQmNoUhiBZ+SFNqHJiX9nHSWowm6vU+tfwnVSK1lL3YAUV8A5TeBUhR
c2LlNJF+SNA5pxwBMWBqP93yD1YC/VRST/Ju3Tv/xK4uEMS+Tnuu0Yo8NfVr
rNxc5JsNem3ckBzAg4kt9EmcuTPOeoNtNh8cs76UBbWajwXbxDiIFl9LP3Oz
6Jmaq4ha1CkzM4SicN68EU00qc9G55fYIAfUbiYQPdtHjt1W4ScmF8K78TBm
4qZt0vgqCgE00o6+UEi493Btyl4fPIrt8HyQ1tzN87q71gDKnO6322EQ7JFc
mfeShHyzkekdxr9MEJUW/iXpwolJslE9NzPjcDB0CvtRm3IqdFGlZj0abtuA
dnoGi9iZzQR9qIbAOd7Q/wT4afzdy17JdHvja/KnlM/wdStSX0jIR0BmuJhw
1J7ewuiNZa9c6O6SPs9mYHan9Fi9w9fo5MAjXdNv/6xYDN+MXKkOG9YutR2Z
ZT8PI+ZsHEQQOLvLTM771dsF68PWRfD1P8++qNt+K3+MUTXyjJyBvu/xMTeD
tijdboQ56oD8rElsl41Byp7JSxrZ0zEc/86VNhuKbZujKVBX3kEFKl98ruzP
7V5FMmDwmEqT27kPd/lKQsBcSWbc8IZo+kisYHFzGw7BnK2tT7gKKoGzNoJA
92e+UEK9QtPimwqXGkfX1kz9VnqbrM/tNLb3U+/rf2vJdo16VopIwixRZneJ
C1RjUBEP29knhEQ74UJdjaEDUlTFn2XXC68MEe8pfshO5aSlwNhBARXXKf8p
dgebpbZ3jtSPV7QS2JvCIHwl8AAs/RZyR9MLgJvfhNGthkPsrBKU2aNacRfg
0ZHetiQYgr+Di6dsq88jmC/8QClYS1/2m0k5QnO/UJUIzMMDJGw2i+F6zsOU
dhd81IkeEdr09dltVk3stHQMlHXZmoV/C6MAG5ZwN8ex01xzni2zdEgnvutL
9dURUj9DOUUJYUjQ0JoE+ABFCZLtwDS0BOW8ScX1/rkye4OQp7bUZ1veMvVJ
xqDkbQuqATjq8ly2EgT/Oti93hbU1j+kZfafsIZnGrK6oT7zUQNskuu6EtuV
dzzIYBSjp4DpJfgJbwDsU+lQAB5eRU5l9nWoz+had5CVHYgfp6qU4RZUw/wj
PYZBqVxYGqhiwDlWTejMZ3cz4KAzM8or8ztAJ2iqD94G4ydS4hyqG+OLIt+Z
f6+SlnKyatQl8cPGT2iOUnlZXo3lVe2rAu3VB1/NgJfJScudDqXBu9Pu0wY6
a3ovKnROP8LxtbuE14NcaXIde56PjcLYqF9uIaV3WGnip9fFO5STYFMvFRTL
jGeXvN5KNcvKr6/UbOsTSRiAwBV5aNlogmmTX46RCh0fvv4seKUeLKgi4G9u
E95FeFyFtiB8ds8oImSqixvFLu1ntrNET5oZmH8iv+cWqB72B7IlNoOLFG1A
7ltNyFqED3GIMtAw9YstVWMvhyD0s6WT1PCirmwD1TEtQ+0aQzqRaazJ8DAc
a+tPirsopN6uE0+BDfQPnIV279Fis8vEnbSbqaMBQAOavuqRm8SUkUGUvLNZ
MJFrTQxZvC4bAgfrl6MpzEpGmYxTxEr9TEniVgGOM4Zw+z5A30enkotTwDel
XJOk5iQXkzSP2i7hhuIsYGFfVGcJnRWCH6VeBYFnRf7GTpG97J8eJN3wJIzD
dN4S/vKNIjJDe9ZulYz/WF0WrGrO7iQ5F0S2ayWka9YS7VbtN4XcMsgXiba2
xjYcy2gjPWlnEEV5zmy/Dtg5Oc7YFJBw8nYIHqoLwa4XBQkcjZtU9NLjWkaW
SSD1LKRPRvq5KaFQcwNEM7RQNBuZmBkS1W4Kyv96qDtI+l7pY2N/5tDbhbhv
WxQ2VwesBknVPE/V7qca4G97dabpJn8S0GhA7k8sL4H8wX26tZu0xyG9hUzG
zo40pCpBHVBOEjkE+C3Jk7v74fz6sJop51utYZ3iNWyk8nLrM7lHwU3Gweq6
Kn6PjvHb1ApY51xJM+i5Lt50BLKCon7FQxfNk3d+4RJC0UNOa/B7C8XqhVno
e1Rt/hUz/GY+z7GnqQyY/BHs2oBbQ7i1O5X3FlqsRDaVvEWJsP+XQXbOfhJn
4ZClysYbx6YlWoqD3ZcT0w8c6BX9NXcBpOibL3omlYXBvjgou/5Pa7G7t6L6
g6Emgr4ljAdh6LKPuvOhjftLB7UmlLdhiX0dAMgvkFrfU7jmjMerXZ5gH227
e6Ed9+2s64EoK95Ci7vrxj54LW/KLOdVjKVcyL7ewmeWxuJCAQNmBTpAD5ts
spqOwWvNABVLOM8EU4k/WHMN/hNeW/wKQzznOnFAhdLYkXoDOsQpe6nmJyzh
iIA2JbVpe8LCe8Jy4rx+Q1WzzG3dMVmhSJkIQttcopH+wF6FfbjEjNDD9Ggx
8yM9TF3VcN2mXbb5UiLLUiefOO0EcV3E/61vyHE74wpLTBGf2VW6ecPvxTpl
7cdbUY+NC/adebZWOiFLiKTCLPw3hU0mnQDm6vWyUZ298/ASEWc0BDsFPXRf
rBA2z4ClOPnzcxmAYVqM6qQX5D7fPI9dPRRK+SH/nK9FOqBTyqszPp4dTs99
oChxBEm5geb8R0VhP1QA/fb1Zvm+t/dsQsh6dtjcrCqkefW1feQW/YvS2kh1
S9o95dYeHULlhrragGeTJh4OhqOYnI330yuDsxgq3HcElXwpuJfiNLtEpPJu
ZHplS+/LgwXi1xkygw23gSoC1z4Os4DADjEpONiaXOhqcMCymJXj+e1/JBhG
1z0ApzRNjoPanLsFWj1jHPXZcpR9zEF9TZmEfFBTag8nyS4t4E1T/En+amVj
rPsk5ZIlSciWJf/dFv1mnMgSJHLWdXt81G4IbQqsEfoy9EU9hndwipCQjaTp
RHl/vOG4fsIMGzBI0hEaDNKWfA1BhM7zisaiw5XxrKAziwTfVZsMEN6FFflz
7n5ZMbR8qzQOx9GqNzOm41oSe3X+H5WpYVvAyiu0Go5h99nqAuY1+/AN6hVS
lN3z3iAC6jD7frb8+AhNuuvy8Oc9D6LGXUcYK6siP6jgrsFEIBhFIgxfCdRL
MK/HlsfAmMlbrVPAyN/OGuhjO8NhacVT/fVNspLmph/VThVnE8XECS7GpFCQ
WWwtZgralTOoTbWthw2mQGFHs0RASiTEuzoifCRs7HK5Rzg2maDPTkxvyYL2
1eToc8LsExdxkRD0ZLGGuT553MWASJGCkhcRtaDGG9m6AUoUqT0eAUOV8q6s
puh3gm4fqJjzfb8uIrlWGDaETwbhWRn008U7+js7STReSFbE8asV1HSLuoHl
sdCc3P5AFGkyWTqH3qVx7n+KFfUkp8rP8XVL0vuvv6SBXpXmbQBM4zXjQbvV
Lj8+onk/hi6Kf0lUvoHPWxNxo8V+w2muGEQ+IVtDuEqOSBTNBB5dlqZMwHv1
HepbViRjYNVJJsiZaapi/H6pzpwfiowg6+DsqMAz76CNBTEYOCoN0kwiDcx/
AejOs1quFZVbtZCZ/fj9L89ISwQoJopvKbF+l9fxuL3BH8sx6VcSVB8TXAi/
8XHlHOItBjPEAcXgXtYrBgmdSY4hXq/1OIaG3Zi292RsxwkehIuV3Ntm4yf8
IpOntGlT6+hCG9u1IGt+8XgaLUjVZ9e2xPyoUUUk4b9L7sy6NbzIfV1byjFk
o/D7twVHCQMeWWOZKaIa8FHLG8fG2jAIi+ZT0i4P4MGodruniRHoKt7YvW46
qPpq7aFVQFC5OKwcB4sdWMgZXmmpT3xKGHKl4KHOQ6Mm80t6XF2vRy7K7SR3
LpqID+vuG66sumdUZY67Iq47Rs4z1ReMtJcLg1MY7ujrNJ5gh7+St82Iu6Mh
kZ2YoDpdSsvuG96IYCHF53+YT+YG5Lkw1Zdww8iujgZDNxpes3eaNc6sNe9K
3D2/raXGbdiltqiCW8DoutaeSmjH/tWUPEDnbNITc0qk28YMIQ4YGtHUjRCI
21GXY8sQOmstzIruLx6XC8xhomEQ38KVJmbPHG/X0umca14DflJKBGoGz2vv
KqUcQVAI8d+eFqlXG6MzQit3MLyAqI9BzAAgVAuCue5t5Esd8HiFxgwaXebr
RS9fjMmA+0BWRxkl91BvzL54BcCDOweZCQ5xuTfGYR9BzdmJsg83mXdaFor3
SAD/lPuRo4cG3+xB0GYKsWmZwvjNNXjzizS3AR7PZ32xHxl0vN15ZifNXDEN
upRXaWmepY8adZehMmbVBh0kb05R8WADOOeFElThCXDs87bMerUD+EesfeZu
YrenP5EZlUdkKDT8YtCFAvAyFozR6o2lWbodlhJZDPsfQkjB3Zu9oP+PA44n
a+Ry+qZTmoIFXy8FdgQvKp80cug1oSBlDXhzVWBHwlQm4vXMiXPN56iPygdu
iKwY795SInXWkmkqqNqKo5V3Zh2dwF1GFAi3y+l+qJfoXzmXPCTc1Y4kRpIp
/PrIlPxTL9CMzqwE4RwUW+jvTrpAvIot/n8zEwho2/233Q+1cN9ZgIn6ZmK5
SSEFTp9lPgbINL6HmYjXJUjfpx58jssdvv979nnjkZr9OVWVzRsRWp+Vtz/q
PKabZ9U9YYtlDKacQW6BbTURlqCgtdv+Cg4pL7XGbt9mSJHiShF359/XhzxR
ebyDgO3aSZmAKu4Fqe6ra4Ik1WpDAf/cj4b66F4TfBME9Qp7xnTa8x3Jks+e
7XQOT8lU/5T0jaHFYPf6k3/jMz4Bcw1F5Nc3D5wotA8dt+JeUUXsEMQ03cSl
zaMzhx0S7zoVQulIh0X4B5LlX2S29Mbk2vT7S1LkRXnPKXFnd7AoHjM4BCmf
FIIdRYrOX0yMVvR4MXr/kgtFX5orKu9tHznAWRvtx/nkINV8RAKkKOEXNEfV
9JS9Dy4lHV8Scqy2W2Ed9DoQl4KwmPgnurbikTh5tD/ZeW7BvCxWI6Qkr4Uc
cDCgzGNwxREU5FQIHlzOgbAZ0DfZlsJqy9l86aiQ/ebUzNHQ6RL7U/Vcqi5P
7R2gLb9TghFWtRwsYUP67ppxCgU6kEO0oLjKGXyQubkddzJo0iRlQTnAib31
8uKZ9aiyw26nS4YutrysxVrr4MDisJ2C5XqQBf1pCo5+PP7n5Y2LGQF2Lh78
yYd6dZVoRYoSAWJxTC92O7qUDrSZbq+kOOIcQo29BfoipCXbKB81lXBSGBrw
xw3fD4GCue6DWTvgvyWRYQO9ZuLZLncq/EmRvP+BgjGMrpsIre+IqBPKp1pU
MpE4CQgPOoIEs93Bs2uN9p7l+pxfWIRPb+I3P8F4nEaoWIKYNNiG7PiaF1Ok
c7Uv87cVZE+whrFOporQ4pO+Si/LHnqt6OIm/JkjLty6fq9bbki4yWsv6NNG
f8hvReNsQZbm8NcPVdN+5UP09VWAT/LWhrC0HGNYH7FwknMEk5M4IVg91xBM
5WRTR+ZngCTogQvq4Qks36Q66IBbUYj5EusoDpj9X2w1lWl1B3gdKQGM3W7R
CyVVl/SlFKZVknNWnwxdASFYdX6FpwZjP3TC6/ZzCN8MWWdCpTkgovZUZuNI
lS0yK15mietZo641JqE883kEeIKEasGPv8AH+XXgIJ31BoRcxfFfO/O681zl
srS3IaGWiqgdLl8Y53zroYboIoTNNtMilFa9I3ifvtarqMvgo+seNGkSrEKw
/ZyT+MhB1Qh5HnQZd28XQ9vR/zJOofnvLnRYLxu36iEFRyBxK9yV0kLU0wMj
2Rm5fGxLaGjJNiTdnoSVouoNKxYcG2FIibSGtQof3bYFh6V03edpUsznA+Zc
5AF0Zi23WjPYwzu8JTKmdBfYiVVFTSJv06Y0aWaQc8++SfMUKgxYia62fX2m
mFivYVWbaroblRuyDZyQtZ8jyYZrnn1eN729fx0V9I2xnoTMehSrUxR39o/2
HbEzLMmWpdKeVicwJtV1FkzDMwTgNb4at/5X5pVS4u50aoVbsnGQge8vX396
gkBuDS+Vm9c1lL8IB/PiSFZkR816PYlPjWVvUwg8lGFKdHCNg9SQD4ZsbnXB
e0J6wdwlu4LfSYBsqQor7RyeUmQmr9C798hu00kBftL+XW0pcyKxL9wljhmn
WqoxKRTbN9IE/Crn8/f42H+UP+rlVK36sf6JUTJ5cyHzeOFTIYbDg5BQPRZU
xuLCkJK/segW+1sX0Q5PJ+zXxjvgcjQUixfOq9Bpbf7aSBTj40c0GyKqI0eW
RZ7f4PpkiKqlofRWp2Sd7D3pYnTqRbEvEHtcECu5/dw5bXE4YGyRdi9zGlDN
rjSIymwk4tVogf1DUaLJZYp6ScmDWSMSkD0d5B8zNmZ8mpvX8mKX6tn+Lca1
644YUxUinbvMWFBtZFvGvAvSkr+w6MJOszfD85iBi3wZ2yk4v2AgJpCxZqGi
X6RqCEGiKwDuCBjUoWfjH6kiybb5P3xQt/b9yOUR1MFDJMWgMqP4u+t3Xrhf
Ef8xlp0DPt9HrSuWo0ZX1b9tVCWmi+eDscz6X33xuuHoex3FASMIaCkhdTBg
5FX/Obqo6dSM/J2EVl1Fprjy/QG8q1k5pqoaER+YV6SfC8T29YGq3NXzKIMO
YWo1lSMLSYavabh2vsB1QlBjtuEy0VrU5Mo2ouDuH0VxdBPNtICe8/6MJ4UB
65De0WKvHIYQDbpEV6JRiG229pLxIrYjrVb+2XNy5rDv5oCqfWcllOvug5zA
40kfppcWHgzBiAPha76w2gE8D1jKKSvfda9V0mXUPPmhcNLcNbXK9rCQm2Pi
OFn0O8fletojpOv5kgPN+X7/FpbFZjMeezX2mJP8/rczi1wX9QbYVbXaPdD/
8VLcVZu4nduPpU8+X1yI/5sRoFSAeDN5S9EotasdVXUgOmcwH8s1ks4CH/0y
4GzwKLWLFr1mx6eonvXQyHqHV9Qaf+GDiGkcRaHzTg++XgdegWAVuK88faLo
cvb5grPEN1fAGC32Y+FGhBPjbxNvSdvT7nROzQkLr1SUN7y+OKvdmHTWeAvS
8hWd+OyL+icTr/GYI6mZcHvuBWkWT23TtfCPzlxNVI3Zwhsuv33k7IWCIfHn
xSn2D1aqsATVLNm+iJcZ5ytHSLWbSqyUQhQINFDxjS7Ejlfbmq6HNPNVGvjh
8EHUH9r693kAgj9yyl31ZYmbjhsDCUt+rDMmzxn9BLUGBcuEKCxu4hHY9gUZ
pC6TmXvU60wBlvcsZNXSD7Kt7oH0RvlSTaJ5CVQBPMOFVbwt+NUBFvbMCZYa
G6+qgYsQAAKTGIPxuvmGsh8wEOhW03rDqg8LuXNX1utQrTgF1KQ8XFgMBee+
HQEz/s8Zg14kQ8ADXUDcaBwuh12Ay5uNFfHiocumwVUuUkorHsQsDHF0R5Ok
Geu9mqkebanpOMjU/t2d5k3VFB3tdQE5Na+4rSz/Hn2AEuPD2g5xuPpYjWrd
D4cdnVeD1d+gACD0gXU5UP3AIbvDt7DJVt/g11GzRjB3le4MDaE4+WEtrAij
O7rZgGiRVKIjQb///ZvXyNAorNU2p53SknRRsWelFRnuXJdJishBpGbiJw8c
IAmgl/NaXcEXLKU1tih570HFIv4WXeNIE4WzzPca1QMoeYihBKvulnOXYV+R
m68m9NK6ZfqLK8FL1/WLLHg42rGGEPy25qeU7+QSLlsrx2a3Spsfm6mlNpMs
ANWKPQezLRYbj2ETtd83QK0JUC9QY4xkQo8oOUx6YNNs6nxH4J3C2VUU5aX2
2RbnXN4vvAgG56xBhjlIRhYogR/NQoLx2Z04vnzl2zf4+dm9VEpajFQJHwud
5UXKePKPWS6vbqJ/HduRprHkNqaNQ/Zt33kfm40B4V1mxkK4hZ6ySZTBRol+
DXY7Gx+zAVVRdKHc9o0W5i6sWNWUC/BBFDYqTW87lfJFmSU3Q7g+t+L+XB8y
+ndnUBJjvPi8BH34ov2h2EFGirQbLBqBKFukn9DvKAU5gmjgITsoKYh1WqwF
jKAeHTZLooHSNLRjuk1BU8ojrGCOYWLyMRRT5g0BsGHzIJgkP0vTmQsyhlcV
vbpBP/wz13RyxGz6l/tu4KubD8iYcohLXlbVAvjFNwziOm6r9upsgF3RMqjM
eMOivxnUgVr+JmydmvguN8giVp5ZHLJ8tLYLavU4btn2mCQCxSWGWRhvXuoI
IO3AUOlk+6kZyBWsm8JkVYo1gR6d7bOUix9u6nKx2+oQdRICaf1ivrJ4V/G5
wXxm1nwdsh5lb1EseAfYevikgQRc99Jh00fyVMokRGk2ACHpfQvcKywLexy6
wGfN9AxgOiIWULBd8xqQzUerTexJH4+KHQD+8FQ/wsYbNB57QmX5rhrC4wcY
XEKcYUi48xAnyXHOTxwVCWNecHgRmzJBJymBMkGU3Xj7r2vhk4gheZS3d9Nk
CZsOQWhfHfizCoawNRkkLGxlMecHoetXpz0a0buxQyst4K8cETOrSwBH5Sgu
qlaWTVOPllG6rJhmQbMOTO7wBLl6TQer3c6rvmLulKxNGCZlp8D1AhbmPA9b
Cg6Cd/ZCFjBCNRko2qCphFe261yJ//oIWb0HHEvxgOVQRolKCuZSpD9Gl9tW
NxgH9E63PRSQdSLkjZv9GEpy8Som7L9w0Q28Us/GgEnjvpTjo/wLVmSs1T7m
vrvNBmWFqJsnxTug+UPg0gMBDs27qDEnkV7b1Svr9gXmWvYIUWRevQ4KCb+b
68n56Wk53YbFGameXp7NjJMty5i0FOV3bXzByMS2JdanmT9tUOGo/KFPI3IF
grg4cgikgYrotcgrx2vLLl0sdx1oUHlbqKiLYNPtL/gmt+YYr1yfy4mfJEqe
441ZER0FfwjjL5u277m86uloccSZA7epxZZ8zGt1tngwndGjURN2Sqhx+76J
KpsgedMPS7Q9ttzupUhmDZbwMtiEO00PqsIf44NymOt1GdVYoQRfnhVsw/Q3
Mf2+YDVNaaxdBK6OPeTYySl48jdwshoHSUkXrIY9oOJWOZz4L4FYXWFDFMA1
rMXKellzC45+b+JOVouA+KvApwSKbXvt8CAOfy2gOv8pmTYfNeVIi8tpV3na
ByKosZ1XNFTTE+uQXCIR1AxiFXkE6pOdp00cX/3wG57VB6L+B6mUlg0rhlBH
ag1TB9/AGGoKTTgTlxaOLeEXjevUQuBNl9MYE9Y39g+AadmnpUJmRXv86jKs
bjN1tbS8F9SZaBCw8yIkjqEX/axV+t/rOFrRM1qjgkb7Z21tr/3KxaU6TOBg
1TJCFbhHorAqoq1nM8X6ebIwckU+f06wjOofzRCvx+CMQouDiIBiLH11sFgL
Y2PDfe+bwfrvla6FCU4BZxI74eaMq6zjlS+s9l5OuJRHud9airAFn6lbx7vS
7PFsWCUP8780S17rGida0sBhPE+kmB9iPrydXhjaMhNrzjihrL1NDuAzPCiF
43UMKzQthAo4ujfLG4352ivkT6obuNWVPAWa2KzMelCcnqjLKGkPKMxuD/Kx
dysHeeSN59VuHZacxCUG+MDDiQJEgyMOkNF38u8NHz8OvzHek849aUnGckM5
S17W7V3tft7x/BfuLzH1W4NFS7Jm5d9hNg5FWtvNIgY+HgGASMdKNXDJc/CU
Wpw+KkX8N/t6UOqLLzw59ZvWITaXBV5Ea4hFMFLi166OaHBa4W6pXAFMaw0G
tXFrABrkwYn00uxW/NzZrgKxql/TazUDZavLam+OY6FBi6VmdiavVWd/oejI
R1ggs+009EM9fl0+jZd1IbiPqNSWC61Id8/Qhub+zjgjVzDdZy267+Wpc67G
M0A8P98HfW5tKm9z9ifZ6cOv9OfjRvgLOOQoeihRtKIhbL82yWTZ1fgrBAM0
Q24IZTNx04hH8ojTp2+18mQpozAuTnNvaSoyR6z+PcvHbA5XQTJZD2ta3Yc/
pT5wsRoyVPECa5K8oCprvNqqDjsAZAkRG0YMQ60ZzzROA/nDgQwe1aL6vofO
SzTkO5KQayeJ1Mk27nxoe9pu+PKWR5l+vQMCcf98N9u4JRgzjBzyg10ieMJS
23znYo7zCrmBBeSw92EpUDzJVa1bg1XhS/LTsXAJVgD4+T8UaAgwQOm3glMS
cQxEUVQFdMhzx+eD1AxZTmKC0piIXQq1SPlObednTRe7HkwDsTTsaeTH7nls
+V/EpRjjOy3XSJos3oWP3n6wSsgtr+rLu2T9dak3BD1zGZQd0bNK5f3grK+w
kkwGOEw8CFJ+1lpCuibcj8M6J8BK2EC0YK/ze90PnexF9LQQoxeakJgePCUq
Y6nHk1wf08bHULDJhvBpOXILJOluQDt5ewHMFXQW2MD53bXYuufYldixORg+
GS5BEKlxmdcsX7C6DCQV6k3LFgHmnyGrMlPhyxIvoJH5FSNFJ/sgL4lg8zlJ
wJZqkDM1O+zc6/KaZAjpWrFzh/N06QE5bc7n634xSgynGkyAmbyPIHfmKr/+
rWFkNz3/9RxZbk04MGod0jB1QLmsl0t10RHMXTOvCi53GSN0isYQHSjFUqHo
HbLTUIq/PljEj/AitaUw2hIK8l2wJKlrUY0FUOn020F13iq4DbGAyHEiPWaW
St3Ognmw9NfYyprJnBnK0+DjTt1AMoaPZQIFoCVvmLOjNgCVZTkwc/rY22uJ
Qb4Y7RAON06rFLKam2frEa1T7MF0hpkK6YwzXGzqKhs7r4CNnopqmw4N4DP8
qMEZ03E8hYLnklcwsNj6bwzY/1NTKzqZNLkBMkpwREdQ43Q+9G3ab3JmLiVN
2rBUPKOOGB5s8vrXrgtwX4mxVeQKB4rrrBtvxsI6X0600ISHkyjDtNXVrl8p
8oY1E7P6xnYx5O9f9IluvR7qRZnEFUbri3IG04oNSScRTRdkW1lFaPNsOHgA
UfzTmymCkcBJdfaGXr5fpq/RuZqPwvRUNR3rvF9rmdfyrqdiLlX4nd/x9YhX
9dy/lD5oWB/PbMZASkm4pP6fa0ASKQoCHG4CVvjVE4NApXpPsm25eB9VAY5B
aEyy06uYT+LSag8PmW556cxUFc95y/bEMG6U0RkuatCXbiXfe86I8L07f5g5
+QX5XWd1Vm28vQv/KnSO2SBF91DD4K2fJ/y5GAbOgfLUm8+wvNIZTwOLjx4A
tsfLcYBZiAD3CLtRbmOUj4b0wlz8443b+HKwSl9g5H+GD5uBUDdVDGQsrKo6
uA2iPBcmGa6O4ZByTCVfJuiEkYmLBpksXREAlUdKnFKiSxHS9kJJX/rU+C4G
cj7FXWUqOQp/jRXawbywr9Lca1e4V5BrnmxqHzBUXhU1XKwmGKEKuYHW5Imn
HRFtqMRmB4lMNtNmowZLbn//FAdnDhvNvSK87G/OMUyUM6YQ+nafhLHoTDk1
Qqq6aM3gtS5l1ZXz1kuTBhJ9uQ2E8dSIM2kwHNj++5hTlNi53KvRfluKecyw
KYDNegt/noe8ayobo/BfN+nt9zVAcAH2E8398JwuPU3PI9SC65QOzOjiMUCO
TKqepQhK4ucIBJxmjYIWWX7XPchv/BD9cOWfULvAMyWQYnuYTTDO/OiCGFEr
tfM9QA58ljaNJ+xOdrifut2ceeuhHvQhSPmXFX6UVya9ArQg6hLHd67m4uua
8/aYB84EgFuokLZkCHeUgb2e+RaT11mFpASiK0xBkwePimRyhVBmVAEySdHV
zCVslKoKD5Vz5t5vF3li4+0cKnkBqhNDXdT3F4NWZxwGv5ny6RyTeBp+CKr9
lKwG+4aHKvlS0jj2oJePUcyDMnNxC7ioyehW5Mv0JGn2AlY3Ms1T4oy4KW4n
H7CBAVkstvNpdEmDVdNv7fe2eHgAU4Bs/dL6YBm75D/tWid/z61oiCvLupZ+
RTLDJuW09bqcuRImXqdEC4kPueRwlhlBk5kAFjgSGY8my/HZK7mAzPi4Ixhp
HJIAS9gYYThu9zGDP+bv1y5s/8X70RaEW1LldSXT8o/eTobJLfax7s9qPmp0
cW0QrJkjh4sI7kM9s+x77OR0lGePFhAevQibds7fA4PdHpDZPmm47EuBDbXG
fkze0Glm/Tol9UBB+6t2rO2RkHYNjpobGX7QYG35YK+yeya1mUoto53qDmPy
tz95yV1AdxqYThl4M9B7+fMgywuomUk7l7FMel5G4q/dMu4e00Klt0FZXPaJ
JVBTJutRby/0ad8JlkdlDlp6Hrm2cl52RfftCpH3y9rmd+gKHW3YMHL6IQn3
RVgFVzGBYcoP60YqY7RYQ+L+yHyNSFLd/XzYj0X9xwfkuyr8OniwadR1pPsW
L4BzKIxVHxLvwU4cnNT7lbjrOMy6M7R/ivUqkAO217nd9rwrxYR96AMMWTHB
OJyaZN/Vv5bD3DlrFTMhcn996559q/7ndz0u7NIjJWsFkwFQ/8JhzKFQKJY/
pN9O0pYkSMx+6e+CKgnlOBOaY5CB7qNtvGGh6kVBAzEeL9X7nkqTK/nIZ1I2
WqJr9d+EkpPCIlJ44fkExVkc3NIe7IALDhIolPr91Uf/3tjXw3+HSkxgjnpX
Ht9riWbLyFoQ8gE1VrEdwfIQzf/Gfn7yyzjS75sJp9JpfO9CUEVtVSzLxwXZ
9HICM7vzc1eNCeEeDnibIUtsPP2nlJhvusf/cwxd9uU/wvtAW6Vuc7SmJn3V
1k+GjlIXVAukLbJEo5672Yac7RsktI0SZCNOr30BWavt/0KDrv1K9AtSNxaj
zCU2NDGYd58SVhj0Hp+1OcAn3cW4PY9BRFxLpYQAmdFYKPeKN3vQV3FalX4U
uMuyzCtH7WMsbDzXUrAn8SqK8ymbYGj9eqJ/uT11d4ntcnO8TPdIWIXkHGYF
zon6PONyEa85NVCoDqZDAwxO7CTS+j/7onlmCQzdaFtpok5ISw6IKUcBZpjQ
xr9BAoN9ILnLeUNdZsxipcjWTFVu+/wWI9YD3mJXMNFdlJMzC8jNA8ZsClaJ
uMW8hjpuU1tsCHft/lUm/XnXTYk/LwWAJdlFD8Mpzq7eLRQle5+1bgBvkqq5
588Y9z0X2YgjaTmKBCtDloFApWgM3ofeqrd/sPBIr2WbxX1PkiwG5b+2eGd3
j7d5XDdyT+Egw6+vkHuWyXi65gRsSYPVmS2OaabrIcUeaz0hskcpmDn5Ts9y
maE3yGAnXhUiRVOP9Ho3b7gMEv+E4ATK9QEP+kJrAU4xsozbQr4qNB2f+JbI
sykC8d3YJ2YghMdQG+8r0fmI2oWTr11OF3w5YKlvAp+h6cs/Zfyi6uRcrC2o
M1R+ox6sLYQaG+wYwFjEVFz3O2X9h9fL9iGnE4LH0lZZVV5a52zXpVMl+fMQ
pWUOsm8USTHBDP4oIjIzLiXDSNCabOAeAH83OYzPsTXHve8Gc7UWpW/ZvQHe
9LNxkDjhvdeRTw6UlLTRDwE8iZ41FWvomKBX2bPw3W0gelkxMevauk+LPJFz
HCfPn76RPcmO73r4uOhCcd/b1ih0Z7MwgDBY7Z9kVSE9FSfpGvhEGbTiJ6y2
TJ6SLAC7yupNPfpmJZRcVlgMLx7meakiW/5K0USCLYeJAawdyh30pWmIdldu
9I1Iz8uLFjK8vOFbMSvn1kAH7iAe7pDfJcxJwNmEXJbsBoQqaucp89PjfKOM
ZVx0aFRCh45f1HZMjweLEaal0RqGVSj0KEGxzO2Fppu0JURdd9kO2BB1V/ph
wdSP4Zf4KsqtrD5NxqtCQ7KcKNFcMKweP566aXHEOE7oRZ50GtyxpcHOWzE7
1qk3RGB0nBY4DDqP65u5ee4ka2yGhDkq5bK50p2SGsod972C6CjqB/O67S93
ScW9OUfF8+A2r8n/GgZA6KMaNXQr6C9IbZR1qU6uYlo7NTgjLpzQe8Xe1uTe
uo+oPEJWKiHS8nfenBGcyCAHYnULxbj6SZrOUdTev1b/3v8G9I6R6qP8wf4S
9jfvTeB2h6luPvxe6EPV9f7mq1J6jIzkBuqNub9MFs15CJJHhxL+SVcE1giz
6U0T5S7oXvYeOUt3h79UOcV/P27T9qMAb5pVKrdl8CcwHtbXStIW3SOkjjSh
TMz+MgfCdIaQJPV8lDSsNwEGft1GOzRAugS03RyQh+WAjaZRhuXSy5uvdNlG
CTmdSrZF4XBn2e9fdz6XhH5leXJ4TUZ75uhA3g9hHMpuesaoQ7PxP3uYSUbM
nc4LZo+VsBQwDxVsBpjsk/h9gNzMAdq7rWNqKyt9eVHG9TBCA3Ab/qIvWXfw
BABP1oxmPlr9hI+pV9eJfWfJvfXhu4IC0OU3gACVGtts8KjCV//COPbTlPsq
1v7y8QuE7Y1TCztHkJKWUVsQlkC0hRKbWakUZVmWjMb34+y+UYeM9opRrmvQ
G0cVO2tjqjsHofDzwHDDHfP3ZPm/EZ0+AT7DTIbLRyP5rv47WZvdR0/K1Xv5
7yzY3kDYCF9LPzJQmG8o2eUuUccm7s0J9bxVrfsuaYhmc/ivKMQkA+oBb7yf
6/q4gU+wvWMrQaNlN7fzUMjxkXsQsN03Ckmvzf/4EOVMq7+HPdlLj7zEyXf9
hf+hVoeqsUd+lkpvRSb9P1TNGDId1Ce8udmZsT/NnsMjJgVlCx95WgwFLPzf
jqdPBW864UzUg3JUXRMF1rvLIKubVnr8RWReUugPCHNY03Pfy+rOu2gyRluI
SXghVr4w5O4fl/xOjlhIWUMF+TYz9juCcv4FR3gY+9nZ4RQEJEaCI3diNOxE
t1ImldEY+4rFV5d+Ez9YPTzzlpnDtekgyotJwUsJdy1AvGUJ7FCpe/TSFb5G
d3YxYquBvOD1MvUMs+oCjQU5vNaH2ktPGTPMv9/MVDkege4mMg277mZi8CBS
f/f+dx6+qIF3tf7QksPjIXDqn7+ZDAZmudcz7AiqaeCQs5+Q4fR6fEBdIKdD
HAYiKuKa+/p3xPoNEXD9/5t1JnLkQx4EbN3u+dmy7qczxSZFbsP/B1lgmozt
jB5OXoWNQ5JNeGhmYQmR90ZfWlVwhrTKuBMJqzP9ECuGoeu8iHVt8jEccMgy
+3FA9PH1Uha5jIFTcZR9gS4xGilPXTbaURCU2swLIzSwu4qIMnkCjv6L5HNa
M66fqZVspVe6VgMianXoGDwPIVxaM9EeyyBjMlaOeyKEowbT/9xvaGJjTL0w
BB5qeLQpr7wvlzr5hQ5DI+v6ABnTeWZBeES4oPXR9D7Y6+OAGxEGeT3ScYrR
Qi3mv5nFsFxcxWo2OlgqZH/AsmHVNk43yxye8Vxs4EGzHnopMeSMIzDnUznt
V0xfZ5NNtX0pAqGhAr7hsJ/6DkjPG6tsNjTzpmnPg8YcXWgGU4UKPNpUFA4m
EvAu3aI7lGfeMvAepdX1iqinPeYHVL/kWYkWoDrUcNZP4qbxdtO/QzaCoKyP
ZdjD0Quzp1DMFCj1iAFDkhjMQdeCBN6ov/stlEBvYEjxGNpa/Dwu5n21xTUG
6YPBbj8IZKq8zxuTQFthkx9HpY1lMzetBXoekTOYED+kM0PNJx8WjYznnQUL
iYLMuwQKLwyvNqUSwJJdXY/Z8iUvaHNPIA0pVPC3uGC7Q1d6eEy6wlb7yEVr
gdqkH7+TAkVWAGM3yJNKkSTKCG4HDPEkkkpJ3aMdfx0UGmg+LgjNUcbkbov7
eJCwrVmrd+z+ekL0vIyd453rU0OiNXDJtjmnGSzblY/5OnIVBxzHLXx22J0c
w2cRcDI/1zIZpJos6rArKv4iAx6HTDGOAp+no9jP/IoUcgszpLb2GJnwNMSR
aQ5lDuxXV2So+1WTlDurlIAaS1Mfasg9xLyrqqeJxwWPxse1K9f9JxIRWkw8
RhRmH0lHHJ5gRaf12+DysGq5KuEtowtO/ATG5I2wEf9vAGGT42aCbNVGVfxM
dI1KgY6dYCFT2elorQwPzF+ILi8cE/Ua5nrVq48AtBHdUNiqzN+OhbcW6sav
IG2uQGFy3eOvHJ19pHl0OUyR33P6/fTtk/vmQisgqc5oGZ3s8Q294zLdtvr5
/XsB0tSdHzU/t1t/vMJ6FMzO7EKE/EYdt61DQXMrP1X7FU3D2fmEczAF9Ln7
RJ4C4tKnQ5QuOdoO7xKCWgfnr1nwbsSdx5aa2m8D7YcUMpY54qxL/Jt+yjjE
5pUVSK94WenzP1fqbnqMOtivHPkQuPHJpf87Wnr8mXAETt2rG4fzZCFZ34bY
+AOz4fBl7O9VFU3ItZlDjzVe4lYOGLcJ5NlCm1rUofQUlkMWtmOc5nKj5WOZ
D1SZ634hYvZgaKglIMv6+hd//sqQnS30y/PYeVOMxwo1KVIqe+RivBmZFULK
RLJjMry7CKxHgfkNZxJrYIkyGtXdKJIU0fgQGBmvM78cr0pGb1tEle7Rkc2x
JNFa9L+K2/GzlKT2aE5quDydaGFocU464N2V5QOoyqYbwFvYkdKHFB6M7CNo
5ddNEQUjsvweDw1A3pBm1Z1JYi80immWGsu6+pvICU9r8xJoAxFCaq4e2r22
mrGHpyM5gz98TGk3CfP3fnGnZK13DCAZXd3OtAg/+30nuaoloR66r2r5hXQC
idtorrFM54jeBmKdzWODDTfOP4o8b4vQiU69L/WebK61xCuBqspghXlAda/z
sLu0DHwcb1zYsa8mjV6A/1P3mya6rn/paq/BwzEH25ZbYYtTwzoJFl3fVp3A
qBu/m3fgyFEpN+w2YRdkzWhFIxHFPSHxFFiuAWsTyAoromQTm00FHWV8GWYM
4ZqeNZB+Xd3+1SOKSCfgeqntgOtArBa0NSNR3Vi+9ffFwYhvBkvUoUf/qqD5
UOMnri4EfMDtQI7484UhVV2B+aLBVHnQVBgHGfimTQRJ3FphncqrxQOqlPWa
q9iAWO8yZ+lOcuyTdYEOstqJe+Q05nEvoXPUIYCJqScWvEfX3d2dCzcdLDwH
/HeaA2XchfuT2DgqZANwIjmpTmIta6Czw+sNWZjCa+qiCs5AYD3n/xgj5lR7
qhljaE4P0eqXu8afoKe7CXUl2PHMQN+D9IDOkpO46pqLBzM2zGrExIdAykYu
yuSaRYgDAlhUWH6z0a5rSBYByV8Yr5jtJ8QlWzlRwRJM2BUVai+0FBRFZA3x
JO2VZ7stDOCs8ehriQ/k1afVUqyAlHwpjKTQQVK5Q/xAjQC4MritPTSmvNR7
2Scmhew/kNcqa2/hEL1K9EdUdVP/ksOLiIFm8FdJil0j2fVePTciYepUidSD
oIBysRRuCFbiQQCkgkaCPjuciLC2SxaBa8h8jMAt/HuSQWU1+xyXcdn39Ep8
VI/OV8js15Gg1qNXcSoKc5AdxVw2koZWMOBA70bmofxHsBpGXHfHIkG1dhbc
FsIhaIPvkZdlj30QBVrFKZ7grx+NOY/WWsENzv/Onuy48agPrlna34BmL/hR
9Hs3Z7f2YQUXShCMf1ZtX3an+v6aH4Ziw3ayHTpAk5NNPxR2WWThs7CSpWKY
6oqkrVWni9tk8uTdinJl12jioYL+rVBXjMaBGG4/D4GvjS+AqdfeYGK0h1iY
N84bNJa97qbjvTlNzXm4kJJ/u7LVMQiLxC++OsPjdB0yhJmMCMTEW0SLRcVx
hkKde3egix00IZ0i2T9ypsCfX3WGw6GNdhUA91/ivxhO5B9pGYwUfv/Y+/yi
drNvNEu4fVt+aKFHixwDPMjHToGiNY0c+NhUWtDmqgOrg0XuSCBRsNtyGaQn
u4Pg+PoPk/oPmH3bWKy0OduBQ11+/1CqL6vmTdvZ62nbU1vUi+jfhipAy/kO
qN562H3O0GFHrkgvq0Pas02/AohJnglqJFVoDSDWBfPzxfJtW1rQOoyYMup6
t3YsPYj1uiMAMGjJ3aSYT//vgYLp4uTPVKSrZtfPHKti9Ccts/+NYQgwE8Mt
WeP12/+OaWwRKnIN6LSC2AlIiTAjqhXKegF8D3cBDXmffazEU/sHYkOEZRmt
7/J9twEyEoEHWP33WhflZRsmKt+npAD9pgJjiCZSxWihcYpSvjg73lVVyM7d
07eOpREvNUBR9xmj/cQvhvZjb8kXKB4VxdYoYU4up5U8OtDGeYu1kbkCFU8o
lJgpJnjeL1HOF5kTYQhqankaa8xgOJvPhNGu1ybLT2wcyGyXgEvsc0CeVFVG
nDQLS7NtmpOmsLbWrbgMFQsxuvNkkoXdiJcbdzmuMkWin13dUWIoTUStgEVR
Q9Dt2k0I53wXp1cJNDYati5ppVq9KeYRFRxtIR+jD9Bn8WEA+nMmHvMD1WBf
8UjRxKWA0SclwFuE35E79fDuakzbu1BMvImfMGv2jcxbnlYPQVB6aC00R4a7
Tzb0ku0A4qf3INLY0TTTXftV4rZBcUpZnfFWE7NgXzGf8joWzdirn7tqa1hx
5vlUn0wYLJ8BXOsiKEeii2i47Z4W7NMVR0cI58/TvkpFwQTDbXZXx04bCz/8
cnEeQzpG8kQC/a2FsnZUUKKxy1hhPPaB/XpxfTlWNRB5cHOGrQsEdLdceQ4D
Ge4C/AD9ngiiXdxEhvuhInWlENOOr37JQoEo8JNOEJJ+g0r7m8Oc7D72hCvs
BCpEcMYOaZE8KQYWnhGfVJyAsk6xOGutbx7jlYbyQscKGshH3ahZpTDRcsya
Nig03YY/iK/a6MsMA2IDadfMvrHzzPgIh++U4Ixs0WVYsFF1GdiF3sEOnmC8
f9DRkomrO5g4rAjGbV7iNxdS1TvEsuVPT9NFVIuhFcIQkDF2L3rHMKy1kdxT
N3cvzjuWWwg82dpvmstPUkMlT68VfP79CPDVQ8Narw093pkRObvUZEa+S8Pg
0NSVIIOn19bMlg75YsiOKNQkGdWTZrNLycrCTUq9nIZy/kDwakbVncTIUrRD
54PO50bJ5ruyOKdVtXxCdAbkA1REIdp2sJiF3XDBSmNutaKeBdaW9YyNkVvX
o1+bXkVnnRk62wnkze3AGLUP4Mf3WsMZbly7qTFuXqKZeCbJuFh7rG9dkibG
AE2Qum8kUBRvTyrzcPDIc3ufHChnMfNrS9SSAFG9PmiZ3G07lQvGwWD1MT3w
AbqTFTJjCJEzEAnrXPWrTjxZf+bGQOJpP0Bwv9GKIloUS8IyQPdYq42HKDfy
takV9x0vr9h9qyJIWFpvxvgEryFMevcUvWiI+bo1eQ8+/zLkz+3TNL7nIXOL
DBC4f+ApyFsmBUvhSsf5BnSOfpix0ceA3+st+d5yAVWb0LgWSGxgoh3TlI3l
YcV3bQjGbZMDMfQcDigMsNJMsd1Z+Ue5YzTzY1lhNxJbVtvrvefJ5yIaPs0Y
TKWQlMVcwPYRFbN67K/3pNJ14lnsp9COxBWo8PO145lY2pvhfs0Zc0ROI9OY
HLfd6VRSYGFo0BnpHBVFX7ug0OrXOOVnaYuiKTSa5SyavBEKfCo3DhCh+L3V
4iLFJEMyXsxu2cY+FVCvj1piy5vwg9Ym7bBfxb/7LXIJwgoaHP9QnIwcqk8G
gTAqUYaXh2kqdFZ8/0GTgjmIelFtbFwO2DfSjCqn3i/pCrJskSOUhLIIGSzy
/y9FKRxGbAx1cbXNOJpIXvuzolrYdJbUNirXFvZb7JUPNEtTqJfPzn0COLkM
B57ncLki9dpIH5I68DMbdbGMAONgQbZbCZMI/KuRF3NlHSxOIdSnl0e3Carx
KD192du1QRDATKrDKw5BzyIzxl5WrfBi1W8g6XTchOdZVjbFI3v6KZEXvs74
j3QVxaotywoYBSOhr6GiEZ0rbtnojtBNsz8K6huRWWVB2cRnKup6N33rE+CX
qPQaSlVRNRdRMJ+iusEUsh6vfMJllZf527LJOEcwTgFWQ37YbkKoR00D5/aa
vZeNX1ujKr+DjVDjM0JORoJDdIr+dbSWFUo6/cpRLBDZAEjUqf4nSFdzpwfm
aXZBiZaVfDJ6KDb/iK9Uk6bqHODo5TwElWg3WUapOYZnxghlkytwPg2Og3bR
E2f6qMSeaqXtUxOgijbaLI/kevvRj/ydKVcqsYBvkLbR4iLLkUAr8eEhy3vh
y72RIsW5oku+eQE7vEwWl6yOutd4lDaFdZZYp200d8yqwpEvosZQ1waoUeBI
gFRwyswVI9fbpxYZZ3IBzXQyfe1SQbaMcuOynrV8Xd2WT4heamZWROQLL7Gs
nwjnEtxoO3XcEYq75UH0b+x0XpJIc5/DmxwQp3goM1fNc6syBYB4rE00uQY/
o+rY0g6OlfEERdkWaddHJlfQLJOJVfKRHZyQDkR7fuNcuKGOMv66J5c6WLED
4UM1irRBYugvihbqWOoOtl7r6FjJ8uqUlkFOoZbSzZm/FT4RqWicQnCKZMSP
pztr4mPAkYJQePWrL/UMEOYRnP7TtPL6vl3ZpslzkRHbq7aS6zq2qlLbhcXq
LT9Ykk3rgXjocidXbBmdHtfmBjYYy6RUMeE3mzxxNlxDb3h4WHyME5no+fYR
uvJ9p0d/ee5TWqD9AcSScZ3O+L9WKlU9embEfeRIU3WVwvevJuZnjs/ddXWH
o7W5Q/o63Y0F31oPK5/wRomI9VtHFU2uCx33qU4hADNa2mPyWic+UzgOMRey
sktjQVWOk3mEM+qro5T6wzeQ+zn6x1d5S3J/QZOLs2ZioywxjZPbH5noUQIV
ehNjr3LqJSwZpG/yWWmS8QTWzk6esvyMNG0JoqJYAzg4gMZkoEIoiHwL3GR9
uslFjm6lBnIQY0o8A5x/+CTlhr3fB/T7bwEe8TL2XFaAdJxfKAlnh/CFzTMS
9z7Ckifr72SIeUchey1OvcmCLd8Lbrh+2vZwdMyEXI6t4lp0JtQ4omueUBq3
6QfWET6z/zK3LTm2/o7HGCDBx8WCRDGzCUwEfOiLbQjl4caj9efBv+ncl71W
1qBwHcZIyGW3dfLgZ4NW8hwnDn9mrZYIHQiIWq++ngCVYCII3LhrjRyu7sCS
5vJ/YNtjJDcJO+jqPmPENz+53EcljWKE4XShPV/Q++07ro/hfkaqXxSqGCZc
cXL0QSjqOnlPbuFXopZcb6FtTUxAcWxqTzCpi//EZqvHyeXM9OiaTmKdamIz
fXvbuMcd9FvYhKLYhuxRvaVmxXFktYnwLNQ1unaE9G5uKc8I2oOhsCKmrT65
j9OzRV5moC8KfnPyNbsPju+8vlsd6LL/mWg24+ABI7CQPmRRyxn5b/M+VqPY
tfj1NmzMcPJawxzFziHKYge674TUGKHI396AtRvL68tXBAAIXOiVuKyAfWJs
3tuAYslyviXbasPSg/mlNkIqzzO8LK6dGBGdu4X74dAG0yeZ6hifJBzmtF+I
1l6WXIheIvTHcf61/bbgnsqYL+rrktrBTIZbytIAaIs+6zZec4wlJ6/IX7/s
ERtJe0ddFWSj/Apec9mad0lRYgHVK1VVHIwfWZtC4/clE/HZtd2JduGzTg1D
rxEnpFfhm7Uum1s4JGY7ptIoQyAZa4/PRGdZqbPl5wCJGigMV0QaJumhaLHu
bdfMegnjlr/p2iB1hxt9+ZLCNGJG8xlwyg7pdU/3zTf9mcKOxxuWDaJ+sZtc
mCIAUOb6A841VXQMNVThifqowOXmcu3jLnCYeVEp9j1cx2TUNuvS6tgtwJqm
izSC0RfKazaXqWz3RqLcpAywJk79zKtCgNtPr9Q/VXXk+tU7UEyBA6Hjhp9+
dgijj60VWpMpzD0GTErgx23a83v5AvxNbQfAgwWYDsvdL1Q+xLSAgUjXK9D1
IGYszU9DwxNBipKl/IE/XfcFrSBUSCYaClYuZs5E/SdKf+NXpZt4oSPh10v9
Y/3di1BPP3+vHNrZxpQS6UyPbAKpnRqRUfTCsVUvX3RrZBXf6jjtvimesZUU
8etq0dDYTjBPkcS4Cv73gW0HYn0+79SXWesAvQOanTTmrFbjGX8TYuLxsGmY
u66PqfiTJ2IiGLLJf0IQkD+asppWPN6ZkuRjpAsRWp8OKy25RggZfHeHAXU4
LxAfl+4csROI+871EO6Jy7gYp/yQ1JrTdARLE2v092twfmw73sxPA/oglCO2
ja/2OCJ074oOGscrrtDAoN72dD6eF0qtNWo2/LJy0/YGq3EIq8TsUMxWpd6U
yuGUmzjxNUcZK4c6hHAMDOXloOdrtFcMelpZQg45UqnYo0uu0b2/GZx3bZQv
VfAUWgnAFAO83MZEJlzb+wEL5g2CnjMf5pe28QuH37R9APTBOlSUogSkN/zm
TVGaenQ0J8UQczp5kiUpFl0QPCNR+C2hKYXcmAHBOL5TTtRKkYY2x3hM6+yd
UN4ZasXRpkfGGtvfumMR6lz5lHNlM2mBDRHt23oEDOT1hNG7LNmd3I2gW8fo
ATbUXTsTTE5gEXsK2Kjmj2hWc6KPJ2Xiu4NIhRqlam/YbS7qSF57W1F+EUWc
dYYzTCQgdrHQ/vS60j+Hr9rndxZOSxMRf6QmqhbcW2e+wW69l1FKpOspWVvW
xjJlgEhMcET5sp3Fm5GfEzsUeg3TGeB8B2jbqLKJztvrqtgBFm8bW+Zfv21u
e515zpdDcWoMue5b2uWZEStXaefh31MaOO4M3maB0XtK5Q7Tw1zK5k9beuRc
HWXUoUPQLcmx39ZEiUjJjmMYonIQP+3uBGFR2JediyQ8Yitx34NqmuYPC6n8
DAxaUneM/nCK68pRhcykX2qlsRWtTS1bB2AGl5nQSY+W1tLnJzU4LQ9CdNyT
33B4g4TmGTwgFQhTcFMRHG8jD9FdUj42bxSBYf7ppESEHhGZA+COsLPFPMhK
ckfhAOX5Umy9B3Pu5Ytq0Fml7ZfWcFLXI9k2ziArcMNVPuMPWSxCKJalH1jZ
gPpFElRflpUO9qqoV6VKBoIobglg3nVkI5xjztZoklg3Lw+I3lzQhq4+lBF8
6vG8kjOS9/tXU2gLKLsXTEuOS0jHbv99d62IWAX7yUDGP/BP8ZiuEFByWIgk
zJX2vD6rqFcRqlkXbzofbvA2CX2Km0VC6QISly43iLwtUdoOsva/SXab+ktS
R03RtkFAjdbr4KcvX3vigfDuMDGpCn44RvjTCwNbvalRIQXdpGwaAiz9JMxZ
UFmbPep8RsR0Ban73h4dS0kA3XnPxrfWhPyhEocRV0CEK9RmhFr8PfBZgiG2
Dg6H9RikvBfDcg6wlrSNexU3SPpKijfN7zyasoY6YPm44h55k8l4i6sPr/ry
pcWOIPIa+75FM9ytH7ug8zCJP69vVloY4SIwpF66+SzQavrKvKpKcda4eU87
r80R8zQ1PpFFoX8JXZc0hD7OnFKVJv/DCpeYRzbbWWuz4EtCYgQR5PJVOrM5
wwY2acDjB5bAxFjPjtbOzw4IHtXCV3t6vpn0Txo2AtgRKp4r5EWGRWX8KWwi
FzSI/+y0rhrVs1GrodsSrL/wTwx4tkZDddfXYykq5bbNUsiNlWFRLuhJS3jP
hMTxpZOcn9IxvcTtMcfXJIoJMCdOpFT/WgPUaUxzHT9uSvqhwYQLAPo4/Xmd
ITpblpQy7UrQGSYNlRb9dAiunLTrr6XySAt+6fAE/G35wtddAboreBBxRpx7
s3yINYCAyRVLim02ZNCrYO90mff3tRKFuvEis5scVJLJ0FN7pstnuuB0yMWT
TfTRMr8LYCqrk0731ug/j8NTsexfGe7A3besEG89iEJn2pkkmWzyoDtePkOY
VBgXKURuuxGVImDl2eaQBEWaetwgxAJB8y0q4fEYhF7GhLGP8G4R5AjsDt1U
0elhXX+vQZ6HAooU8bQ8PqAlWq45JHIC9zqpejSyCeF8lzytOwa72kI/54eE
2XhpzAH0qP1nSSq7n4I/8K8783VJ4Ws8tbO0xC4GoIWeTTV6hsuV7ld8SstQ
TMxiga+w92FNKjWe6ngi7BnZWCxMdgbAwcDFDh1nQSqS76/xfb/DSby6UDS9
fCBjqWt3VAQwFEpClHKunEeC8z0rOTP41iSaqey3+2yy+eK9otxSdYoe+W7N
m6SQX3P4bm8ptR9Xy6DMSS3+purbcvXNCoYG0pyRycgLhSKIlt6JxLhgm7uG
1V/dzExjz4zI4eq11s8PREEwtChVknb1D1dfR8iNF4seqEhxLkDXm21+C98s
q6B01vFNW4whImY3wF10pV3G8d8ZVOuB8B5ybxWB5Jkje9K2ehD3dM/f/0ja
ThHW88OF22TiSmrroF3uiLK6TkomK3UdYL2PostVx/z5Ce+mHRlCe1oZpsiU
hQWvnfOqG5J4kn4jBHJLvRNs5gzQDyqgW/sdEQELWIrkGwKcfD/h6+mMYJL5
V9idNICdL4FznB7CYSUOKiBimV42sKOdeoQxcz48kwxTbCM7RZYKHjbv3Fif
YI+hFBgn7DBiHayOZdlXwnM3cygGOOy0YbZdzBOAMi8R8T6KDuqWZ4mAaA2t
QgnQxm0euKrLi6GOkjvGMxPcEhL5s3VPzrVjdTwXjKQtIgtTV9PvHpMvwJYY
Y22dsdoNOReZrpayzWdN5uJeNC3WSWq8jD70Qws7AfaFaefRlNHAEuirvj+O
AqUd6kpdqP54oPVIIa5uJ6XSFcpwS0ghZ3M1RlTvOUfYCQvgAd6uqU/1un1H
W+gJY7dCy9CpQsdhzedCTXcC1Lomz5oi5S2LQcmdrgmb57zVH5PvpQMHkOeU
u56dXxjE1v2HdhVzzPybJ4/t3ODv3dkIZKvnJ/OUWUl4Q5TfvepErNqynMji
PvW/UCpy/ShL10zJZ/h4khpsfvBfcmEJz3t3sdaoU+3SV/QkMdIL8NqnZu1E
blnzVySuYytMHkzANhoGockayAjawpekMYjtuBF8FrEtWgsUAHCP1HSq54Kb
2ijoS6rIuDntkFwiiPjgUNOCzQJQRxqKAji6xfMdhE0KSYf0lskqawVv0U/o
uDtA5dSE9X3wVf6TR6nGjmeQbrWOdRah7cbg5W3Q/nSP1c1yXqzpq+Nu6jF5
Yav69nfLIiRMDogP9bAZ3hQHEJ8y8+jOjN5YIzHeSR66oP3vxMBAcEyv2qg8
/Q/N8vZw7iSqgOUQj1V1Y88WpybFpvQgJ+NtcbI0uuGDwesxpKZ8kTBv48EG
ap0l1nOFcS2o2K1yz6mVsZD9Q8WPXfBCbJwWEG90Cjrf9jxibAqMI+z3m1c/
MR/YR/ioWRs9AwDvR2YPqQQYEnyDGZM5BLavwPjeM5cQtIgGzfQDOAaxiMBF
BURI/V+4EopP+4lbIAxDQjFj2uuN7Br9b1Q9JiYJNJu8cyLIIdeNz7j8tspJ
f508CBIXsHQRBl83ZVgit5YUvRzMn9BOTfgAlQyOu0dY1y2ZIe4t7OiIdXDT
pQbcNocvaQ5Al6FDyu+J3x1L4zlXdHkhh9JSem+eBAMzd2r7UlSsv4ayXQKJ
V9X608OwSTAyibyvQWz6UubwClE7A2It63OsKE/u/37dOOuKHL1QAc75O5DF
iRw2JRLIMFPGeT3QzVYqhabnEKeeOvxmmAevaNsJwwEJkUIGhzcdWsvKm8+Y
ef8wyLBVAdofSJ1UvLf2+f6mN+3Sj/TALem78Lw6iteS/mOXPukNVOuVk59/
9QisRRJvKkIoTCWGO2QrMwzZny00UjpLBxoEw+lE6QDH6nKgH+EviYE+0KvR
Dk8GdBWxYZD+nlJ01Fhey0NedKrs3CsNLec5wbim/rdWxh6pBs+FstXNqoTv
ucsc1NZ6jKlj5uPI4sLeTR0xA/An/qfGAq1ldHSmOGitqlgIvieVVpI8ANz9
H2zhaNEXC2t0GZFBHOqf3xuO/T1EHyctXy8EkDBMFoxyJIb/VCuPBqJB80HK
vn1QN818nyrubBrHFLJlxUglM1zAOSl4BHyrNNWgCPBj1vC6dbUuOTnDyVgO
YCr+TdvcYarMMt4RR/AIUs0rQtm95KijNniKIPMfoAA2+fk0mQQEVZPeGNWg
Mz+dYW1e83moJwUDuTcR5Vr1o7o0pcrDCrU1PEiKTX/74uLWnOMApTfLYNTO
3t30Q72BdU05x00VJQ4ROwc7ceVUA2K8GtolrZbfA2+J8Sbg4FTOuyuaCwqy
e1Tdp2GBcAtMaSXg4CoUByywUiSUMhdUsGabva+kr2So0QjYMx9Hb+KtTyob
H6hJW5odOEIgCTQGy4HvSB1RF6RtViET6OPoM632JQpBKiM+3OqVAiiNFOpn
m/FhxHudgjk6JYgnYAR1eOWsePOEH3o1JIOV8uAQkmQJ3qvaI/026ppPjjcf
VqkaGlN8f3XeCax48TL1hSTgWJjW5DrJkXG/0OTbGDXR+9AqZKOEkRoCLer7
+Ku0hnjKq170JAQ0ONeCV6pPXzLWJQvgE1m37FV/ljHy58e0rigGm4LqGqQI
JN0rLznhEsNp3qL4nN/lHg86X6fE59f802vqML/HAauGCmKyJFrutRd0I1pt
+ZK8Q0CCx6PQvsCkb2eCWwHNLO4BoqMJ5xQPHaDtP6jgCAGDOclHPM+msc73
5R+OpHLEEIpE4XF17JC0Hq0qrpVPbAJmhlr/ZrZavjLBPYIusRu5ImSYN+qM
NE3segzw6gMml7zdfU+oVZSAkW56nxkTecAjId11vlt7q0YDboWiL2NSxoRN
f7bqn3E4scNqkPeP8ePf7UC97ggSuRN6n8x4glqMOghPSFC4i1PqRun2rVJY
CzwpwBuRO+oA9gtbikaWeb2N0ocl33DrtupvYlTWTOb2CkQFYTxhoX94O5Kj
js0BmWhIjJ39NBJsOhIm6aFsSRDCbOdRLgFG4XrpIzy/Qq1O/xvtTAX7UEwL
NcTdIhaX8EKLl7Nd+y7fI9Bu7TyP80shbeB6N0Sm1yTafdjSxd9gkybZqFcF
8aP0PNQsRyuZUiz8DuhZaHuD0iwC6yz0HP9qZiyn6FQElnLJGEfKO2cwCR7K
tgUR7uAACjQqqA7Nm34fVRJX3DCtGFehpKh9fZ9Zr/sIIHlnNrWEn3+AegT8
0M1sPPWUTnse4J4/kgS9bAdMlY19UaOKSVrNrPnvrnFvMBUz19tuBTtLse74
BSSJBadLPlWpZgE3tPOccO5Ck915J5Zt3305WDcQtyIsjPn7vewfHmcFKklR
utKYghSV+QnoWbfMqGiWNeXpCeFWXBfb8HifwKyafGhZJdgD1FZxhMB9rhqY
zizLfuNfpZuUKZsca69mgAkvEl1LvuNMXTOcRM8I/O4FG4JOh1T0CKA9S4bL
ziRKPjsM9EVfNdXSeSrDlJeICl1zm6Utz9QniwegU1Cr1xCI3iXRuNVbswFO
5R0mGS6sAN0/akuTkpXtTlPYQU2YJWGADC8F0/3Q9ACQdtI7AjqX7ZQpPLBo
BMqZITQyELB9/OqyvuAwKfor9WeVMPmrkv6rvgfKOnNgS9pUJessxuQCUwpW
RGE1gLw2X/WDyhB7moxNLSxddEXvdkaMIuMOW1U9YOnwvquhrhFUpNlwW2BT
K8CuE0b8POkx7zirqGu81ClHy67Ti+oT/8xTkHwYPIhcxZfHnY7yC1R9MUPR
EZejPAInCET8moVfRmckj06KuR4KEQOTX8/ltVV9TxihwDsBTrh2HcaEfvbk
8pRiaFrzsT++vBb+rYgOJn+LYFnW0rj6dnpVzhUeFIkounmD9Kcbz5UQTbaX
+HMDf9BRvHTaeMjUGMUMs+SqHBg20YDrPcc77Ps3MCnBW0L/lNSne/RtSlMt
Q4b0Znk/f/6xhckIezao3h6pCQ2J6EUDnSWdr3/z/DJhEcn3jR1hHycP3CXb
nYXBD/z+SazFxipahcVXVlhlkT8QFwio6gTld9xdlHx4gmrlpIhNmdFUPMAh
LO5TblYZw5kwu7qO2dQmL9CE28GRiPgA7xYdYIQLIIymgKw7nYwCiWDkWJDt
2eho7/BH0a/rZxa0+dKsGPxGyXjofMSmDq10ufb4n5ePqVmuTmXEXdooDlj0
vzB6J+BQNdZy7hx4MFLE0DeRWXz5fN47uzsWJAHHGxp0IoFt+nCIiVDkvpE1
Dsx2Dwf/Y/aTB9GG6jql1tldpjXuBbkTDFbRYjJM9uW2vfAAhou1Exg88UeY
aG9KHKn+vWYZg+0pbhyJD4YGO8zcx6gEab6hTZoDf3/hpecDS1ResOKKgRtr
BFmzvS/Yz5yifmjnwz3rsoI/ePsudbr38pg2ORLk2cfGtbBMuNigOl6Dwbw1
61fuEYRPLxs7gPO1zH5Mp1v+TRlLeqHQGz0mx4rxUatxxhrj25/jwv9kn3VS
sJHcYCGXqhPgSXmnl1MHdbEGwHPJgUa3kDhbQihn1hz1Sq/RedSirG6wKeLS
xoNkASSyz+XnYAuFPnjiVdPNrg2wAGWdEUaQ9ItfF0fBAsHZADi2+RIXdkWp
LBE/DGn4vKpt2zDZeT4Tda3S+zmBwAsMAvIYTCs5sUJyxefcGuou7WkqKLef
VLOEFBNE4rUllGoeEmTujcEiH5wp+MixsJA+MRHX7953DX/pzL3DUnUfcrDl
XpGMHFRZA7tf7zpxD7/HJUC9CzPUc2neso4MvPRryQDHdSXgV+B0+wg4zOj2
8XpMkBXvyDoZEzfDLMGuLxkwU1FiPndCJDXIsyDpcK4vy00WSpQ6ssTfH7+I
AwKiT58l/m67p2JvqWuvDXNROKc+kWc0WUiPhTF4It6+F8dUfTYTI6l9WXq0
2zFCm8HrpOoyl9sHlW1F7o//a26mh5YTCOKDPlHKS92lWuS3wK7JZhqQS5Z+
RcQhZ97s9oY/CT9i5iILdUtcZKYbSIPy/RflZkoER8gPe2aDKH8xjYfU23BR
BtfM7NMAek9HchMP5q+mWxfcQ1FFc8XLWz/s0UpWxkigf7k4j/S0sMj7nGBW
r4ICbwpnShnRD5ofdhIPqFpF1sLs+DTH8UNI6IYy9UpYc+NEYFEMV/pj4iqR
vTnytXgm7xGZ6xMTXcLJUQfHt/41o/QMQO7dqOVrkr51SUlL4ys7gaN49fuO
spIL/IsKv7AhWp6H599UWhVyfoMZCyFRqHDqbV0Vvs9aucUz3EaSp+XGQ2eN
ny5YZBpLK7h2VOkNrVJwxEaK+mCOaW0096X6vBEcVui1kwvn97OUohsXQy0B
lL+uEWbMgKN0DN5Oq33kuOPPRXqxRXvCzQi3DrLDMWCh1+sSJYGg+66CZXDE
cVo/iOvI5/tdABF47wXuPbuulkGLYR2Bjm/77fOFiWx5FUPQltMefVBeUZ+l
MeIKQjAchdXBHaVq+xd7iLR/QC2ZyGvIQrnOVtCL2ocvUrBzGTGuXmQFKPWh
ip1PHIdH3TRIc937eyY0PYoZ1/OIKs56PFQO+bXskH+0ENqujkH/TVkKJuWF
aegZ8N76BPrmHnFsq3FnK0NwHFsQj5591v9N95pOTjfr2mmzebaJKEoKmJ3a
5Rq0iEH4pz0C0f4mbTbkpgzdPVD9p1DIBYhP2h0LQOzfrg3/QdBY22Rc9BQK
75ISorY4Q8tUZ6zsP6dLd6OEbDHPQfX7hV+3Qsz//6OaA7CpqWrLp+9oEex8
PuMxNmeS8sbSgMVt+vBGVyCP5Jvdh9JfofCZ3NeiIj0LQ8Wf6RvF8wRG9XUq
IhzcgJMIiAS/mMC8NeYU3grCVEJ1rIBfn8uqiVtWLKC8fBCfPXulWdFcYEA+
Knv84BpCBkchdHpyyjNwNu4Q8JrQ8OJ6us0QxJ6d0yG5DdHdabDT/tnLe6K9
Sk9GHLiLgOfLs0uMEcfjAtJzVZy4GXz0QTqg+/xoZOL2S7J11FRoXTnxFjJi
feAvnvRqgZyBSKSzUXmRSh8WPyGptKLSlzcE7kWemE0KiJx5FZ/hnkov2zCB
FtBE/dXzbJBti8lb4AjUe2vRG8SpSCZYhOIRbVgkWPziqPwQeXtBugNqfbCL
O50IHTi/ucxLTAGX1njZlkM/zZLt5XoVO/NuCtDjP6t/Hqhq/hzX8enGf91d
dF5Q6gPEQKV31DNwTciZfDxg/Vd0QdasHzhmJ/XTfYH7PMLl4fG8k2qH/gUo
YqEOmeC0+Me+PglQ3ps2LnF27pK3vXrepMZ4guSTFJ0V8Z66+LZf0CZsYvt7
n1+2N+QdSJgFByyScWTPoGM4ey00mSCTA5h4QC6mKpX26necyXTtiAVt+qF/
pEr3A6Ho1vqA8LrGIvkGKn4uZEbCwKlxHsRA/BhlfZg1zXFjPXB/WDG4UctK
33WRtE/HBhRAARVWcGuRZsYziKo61VcmBf83C+qQrPt57inYizwSVK4eN9+B
BYMEq+FbuIn4y8kagbXIN7WLb4dvrMmvFToQy3hlvZ1/+wT9eZUymtijd6SD
UWdiq9uwdhAffUPNLRFLA5zLfvFfwn0qAH2IldHyt4wg0H7Cdf76tnVt21kg
FrgUT059M01J6GpavWnVi0A6lbDFIiufAoTJ2JIdl/YELTyO4Yf+HZaiZDDJ
Wbdmp+jqS1ZYGdE/18udBydfMz4kauVX2Uk6ieVQU/lWtvP2zC7mmrcwn8kU
hOyBb7JxWwjqf1Srqjyr/zAbJyVXaTTbITUDRbHVd9bGPZboLMMdk4o47Ttw
LN/ZWZq4lbtsFqxeYRyYC+f0MJlltvsDzsZ5bxSmZ3Vd3dASZnWiHP2JEeCB
kAkrA2rutHlbIe2+t07IYm+b4rH+Djg1317AFIa76Fp43oS/SPqNUewEj2m+
XIfFqY5gT0XtY2gfOsAZ12L0ex5zQH0w+Ve8EdVvXdGNL47oz7WKvQ6CuDZX
vGp8KhcVgDx/Kv5E41BouN+LomG/cJuOFONJdQjLelCs78g09TN23tbg/D8N
Ng48urhSeu5+j8HGKwfHcO/DU55eAC0lrmqLTaf4bubE9yrelNhkwKcnNZn/
12Eoq+ruZrakkEYh8/WLMWJ5yDTkEaCnAJOL6Pn/s69YtK/bK0qyL095XMdi
5FbIsafbgvYp2FK+qMKvhqUKTM8TzQaI3Pe5rd2kcsWn7uXm69CPNnQstjMz
72mmIEEEZe+hz2xXSVzWTM1f3IUfa2i8prrmBUs+QyuMhFYGxPhylIJhFYJW
hhiyb2O8JsPVPNkIWGdEz0l9v3gEs5qn54iCTHw8f43J86Dy75/2y4v9dUae
Fvg4xyPrasIQf/T3owuNdUcI/02UOKiPVqHCeIO0S70LEVW00UcMZdF5bspb
7OaWteLGOWlGxrX9Dkv4dRUotIEcFhlg4BNeFTpHj4y/Jd8kmq/NIL/+lGDp
n6ytcdfGeE+l8T0iHk1Q9mKQaCwIoV/ade+DBV2TSdt8Y/EBcXrfnKz/X5Rh
pxEguGzyHYJ1i1mnCo+rzmoKue0tmjeS3cJ650OfalUsSBBMc9fQTaVI1Tu+
A6TUYJYaguncDNRPES6YP0eBuJzMEWNz+hq0yTawVHrwY7wMHM6QzANAHyf8
mONz1Tf64jdqdq1qLatlU79aR0D117liLNyw0OjcmfFtJwNl8YhEMdA5sZsp
6MwOa8+xCcZ3A+3P0EQTPZBPrwNT0i9oaF8O7zo9X1vdwZRFgmIb5v97sOPx
zizua136XJ+LU6pS5NbZOe2v24ZtrFTm2KA1fnERFGZhs5//5H7labLaoJcf
NE2J1AefzX0hqPFYR5hEyvhW0EPIH5RW3Z6gzbiyjIgVNMRgV9w9eRmnfknJ
Cpywyv5ojkTVz3uhfbFEED7YvYUugLE2vrw3q80+ehLalP7fdHa40H57QOEj
SeVDk1KnRo2w0AFLdHZ1WwzOhAjTM+ukgjjhW9XfXrcWvHRHf7BsY4447b0u
cyEBVtXUiCvOaeuv2zOJFqQ3HBP9pcV8bXF/t9CddrdYBAb7CFPj2Ykvo3ab
jhrDPAC8T0lZZ9u+/OISxFvIpKXp/jnqmieu0oFWzc/hAkAwXQMWEn3N6PE4
Xf1VL2DyoOMSMjRr9jbDKOvPU4SNyKWYsfNHNZxJACyqANtjn8rm4xofkN8Z
UeAqEqFv8T2wrej0wRmvM0gWTHLm3AvZrMERBTHbrdu5HyEZ85zEjUv+lVU0
pxPYH3okJFH/WAZdTLjALe6Q2MBY/+8Dc0+vg9QFmWNdrK2xcxKJNNHfNgl0
qZw8qX16Gk8OsJAP7zYlnbf3UpcGQPMZv8JClqD4spzLoxqRpuoxnYyF4mes
tXhr2phHHms5y9WHjhGOV6g6O0J8P1sij8LFzXZVi06flomuAod0yD7Xlf9o
6j2CwRZs2JCMu5GMKImbv5sELecGcGlH1u/yXALmjxXcnHMfFV9ZBZ+mKI/C
x/1729+Bf7dfUOVvEQ62opafsf8pbFLkIAQxjk5S3zOMvyhf4Ba1n+H87YDq
7x6bcZ49yK+yotAcZBABxLc15X93s3HKstWW6jUPr50zbIvL+7yEOLvfsbfo
Bp1G1s1D6LBEGdsk8hQa+f2hGrSOnvz2cuLW1G986pGMyIkHPA5jhXwnJOUY
PjjBGMSCZiga8MveeYy8tekCrH81EopGY7IySHMOnfMJbrCM6NuM31+c2Bf/
Eotrze5rxuWDIHWBc4V8nTTnYndqmN3eeYzuuSAetm6xdADk93ZXhFaad146
xkoPSv2JSCK1G95C918xm5nnihRdbNS3ulbPk19/6CSnjg2ba6ioe6y21E5W
oomgcb4JO2Jx2ES/LqtVvfYNvDT2948LuhHOcY4fRU8Rkb/JAnkimcRFHHXH
nnQ3iOFoedh0K0o+fdwfPBFus/cC2Eu1DvMVS+k1cx0VVE837gsHwOVLo/FL
UPcLzjPLZDrqI2PXFdfQGIEcBZPkUg6jknzKYbDooxmHl7vBxxtm2YLd8IcD
yEcB3kxmErESxYfjeRIG+x/U0H9JuLFuZwrVrMjTATXMldRy9XnOm6v9M1iA
AIPmG8vMOoztnMp/aaNUWehLMixUDWD/rI0rmltuGcyAS70Yc/qXNpWfzCUk
v9fT77FnS8QpwSX1BsvatA76GESiIoirwVv0LEsKtCdkgQd3jlXi5+NRnYB8
U2Zs95VzQE1gC6yaDtIXs/ay/LeXGfy1E5NBqgGyniqj6YkUbsg8cvJeFZMS
I1yOrXAp9IitotUsvnHopU8rLcBMRwmQK5jb39Xw7Pcn99zvzYrNwob5hgIu
HEjCdDbqbMah/c6V0uK+zRS4eavAwbTLur13HTeMoV9Tq9S+7X6tmiykdNs0
Suh1tb1aMR91QNur0dHp/9LuW0EZiYbWbr8m8khHY8rbvP9R5eFNTP0+JcIb
vXTV1raKt5EUHo9QZ006TYo9veOzkTp0XJQlUb9Oa3s5tao8pbDsmlvCiKXn
BvNun8A9cs7szcpZWJQaVUCAyHWNwrOIxBLj91Qz9gPvItPnq9XD1sKlLT4H
kopWQniPUiJculhu0Sin7VyXYiB1oaZPeIPkeUJ2fUa9UtXL1UvjD4Dm04z3
rmbnbvqzxp3h4hpMElmDml+LYVGdIIAo2+hElWd6sESSPbtWe/XkGPYZ50Oe
ZQphref9Y0HFk+FSoK1LDqmh3KDHbc7mNLMBEpVy1eBGIbMPVC9ogqWYMCqz
yCK9JIGU9pW3XKC85n1GgdNA8LbOe29+mRruDg9hrJhTTYLXRqo373z3xXnx
wQVe/pdO0aQvJkhLFxwAS9kovGqrLxzebKqNcnpClHwsup+dXErvyo6a2xr0
jrIR/WVGIr9KnlVOnp4ARvDyIOJT2VcI1QOrw1Loc1RE4bTZDr4QFSy1EihJ
+S7aPwenXYLSDLxYrPH5L5rSNMZKJThhgJ0dIkRNy92vz5Co4fDRvzv5wX6o
Clk1fE/sJ/F+KHfj/pcGV92xao3QAaMYtgRIymdcYUB5dsovAaqWqmAwM316
6PGvyQ+sndLzifIxAvK969Bww4KMnFX6Cox7+/2R2YM/n0hDDi1i1RdGtm34
XJfiT/L9opYVF5zlyD1aSoSYZt/Zbral+nwXcRrg5ipYxi7dWa6ZmE1LogcL
XDwJs0cC3aUWFJLi+YvPzGPBopWm5IWoXIT4apIkDxJhN4uJ7CbUNS+/jJst
/9b7Y1uUca5iiDPQQ550BtBfy/+6CGz6jdwHkvSHPbEirW8DXElt4r5Bndek
/2D5QKDj5XCB2nnElIILUGgFB0pfrOVhVKg8JOsfs5gW4lWhiwWlSqZJfYS+
8sCqACYfSmUL0rcRtHCUa4iIFPP+V4sNgc2SI/ltPrXI5IL5VFqktN9BNkRE
GM76fCecvUyto8jfqnI3bc/dKba6ewPE0GCmiOQKIOgnd2nHka3htzP5WXp+
56XwDRXQ5EMaO0gK+MydI0XVcnoI1oORxN4OVqdel3pcEdnsU1SBR1IM2Owm
ky3Rb5Ii0DB1fSUdJsCwLAPm7IEjvZMIMNJGtzOwu6pRKPSl6cp2weu68GWi
S8r48gidseEwN312zgdF6hdEIGYHNekvj/pBFzqe2ptat6ewAUbGFTJWykjy
v6xWYfXDIFX5/l+UbfXVr4josgOzdZ25LRc7mZJbqIdqvWXuQwFC6BAsuWsG
DfpOlcyy89H8SYthdm+Kb2D44E6KsbzvG117iUuVZlfj7n4bIgpfDRO5HdEN
hBBLsQA7cMAx2ZsoIZx1NI954hoX7MTqR3637E4bF/MWpX6rKlabEp1NmW0x
XN5ufK71oYF25Iua9pl3yg6tcv4arS35Zgtqh8T3v5qPXW1cJ2jDOTOxC57+
SyfhD0jUNeOmzNZ9xnszdPG18y8hK2rUUge7KTU+ykBH3nTLQjINYx/ONddc
owS+DFid+H6Xd5x5zrTOnEgFv2evSYLLW0mBiG9RFPMlcN150ObSw0HLfPGQ
2Rwaw0GeO6LtOE1QSdJsLjye2ucmM3LtJZeArV2v0668NeOGynrEugFe5luJ
RViX7HGzz7p03Q7J5boLszHS9cyIi37R3gl4UDytS9kpSFyz0UDphJKWhvu6
Cr/+oCR6927E7ou0L8Qo/yzL5G7NmThv0ceKUhoboSGmF60AhDTsQ6aKj+aY
2QpujJEdzFfwejmBxwboy+tVh1j5yyyQCeEbgnbZo51NX9z4nTzaEJJJb9J9
CM+StPXwj7U7Re9r856G2vrSOX2BEQZ191Iu/o/dtCSnOuocAeFZ/WN6u14+
8w8El5Tb2G18EeJR4Ip0MdoeWPfRN8deRTg8zYvb9i8sYyNL1W0WL6Wxvfwy
NJ6B6MpN1HARMarqhkhAktmphTIp/yplkrsOg6+ImjRcS/I2HQwU4QJuvfLG
GPpf7QecBvlwprpQK+I+ZCa9REZqG3Xu1uMNct/3DsPANNqVD7aWkEfNqiRv
+PNkJFiKuKELdgcoXFSAG4gU3EB8nSc1XPAGpHa2P6e+K/F+rp0oyn8L+XUv
t1fos8CYbuNHsFI5rR4NxM80Q9BdF5gJA+BG8T1ftIHu1aI0mzhc+hNn5y2L
AwfODF83NwnwZGJHXnU5BFccIVXjZ+mwVrkc2LIFVYOOeTC/xblhPFXaQzXV
C7eJzRB8rOOT/UgXRoYJMqhLIUMiUqZYaDdurwT3UMyaW8VQ6dB8DG0vygir
eg1hkmqEE5m6gEKm5QbCevQKvC9awumrisIBnaVOZXnZ6K6pcRWooZVthanK
OPjZxMWB8pQxGiKJ7SEmNoyX0+wX0XWIqtlI7xuK9VGqXpOHgA9coRm60hf1
se/tCf/hIUe5qS/uYxXz9CppAOJTO0r42c/St6AWi8AeChx3rtXIMnLa0FNB
Zdtm5sWoiwK/msML/i82yYlpGUFJ+1XwdUWIa+1ziRFGnTf7gYzuILSh6lI8
vCReA4v99kt8+o/DC4y1FvDvRnqpaENA45lEcjiKoZn9Qd8IRgui50zX4LQL
M2sPcJcT+fC77p9bGiYyk4RBTif0Qn0JADbaHWgkVE0HFQ6xTHVgjOWp2LRe
HuDYKtFmwncLBlPB6cWlt5514jrH4G+CTyfDFWKVavFH7zReVS/HAEo3VMV5
JD7y5zRqdOlHr87w1LE5A4M3aqs/YmeCPBSdO2TW9f7w6MSexzb1X3Hg4lKk
KRubI1khlkTUTjHXUmfm0cCV+vr1HUVkjxd0oZHmBqEfS35shGPjsI5Pb9bn
G1TWG8lvCCRSKF64K4iuXchfi8sQS7G8D2R329wlgLKq4wOMerEkqr2Q+hZB
22S4m+FLxLwAt1X7AomlaEpRza1JQ6zB2zZrFycQa4Hdfqa58Hk5YD2NAaXJ
cy1EY+J56pYH49t+t4z/60ObnYrUr96TwExm5OJM31MBs9ubzhXytWf2hhTG
2ZvuNghbFykgblF+mW8Cm029MdTfEsiHiWhFPN69TJynnKItBAL5IZA96vXl
GDghaFGtV4yFzXHm3IFpxCownGjuJz5GCd+Ncg6QfltbpOEAQiDg/lktcHnL
9azoxdLPoFECI6lKWR5icuIsb4T4rOmQj/PxzhaCBqgLKRSwSIPppXVG48Uy
xv2sZKjhYxwCwB5XZEB0XClhOcicftOOM9/QurELsxX2dcC/SC+xkN+I26ey
VFnA55+cyHwh1A+UDASV5xnvO112ANDzZniAuzIR7TJlFUZ7fC6bUSfiitMR
cmGZ+kZaPFExY4034FVRzoPNEL1sNaeaW2kUv5SQ947/BK89sWWH57Nj/oNP
yduwwJ1l57bvnp/f9rxtsUcrpgSKE6LgWE87gBC+xTARBgJlospQrA3LpOB6
c8YSbZ5uING7DKpJ5JqfASSf6o0TgwsgfHS4NN+TXyMs3TZAchdJLK63QSyy
fNDncvviBDNyU91sJcVMtFbB4j02+b3mrMiqk27ztshGOSJr/8l71gqbQEfX
wwGmtHqg5JjX/dyc5eQrBda5HPXG13x+22b46LLIoH40mq5FAXdq6F/Lr1YP
3jVb/f7lRjfZcTqc9CQwDRJValwsKLgq5gcKH1WEthCu3xvcHXCEpZero6GO
wb6uDf2oWND8cqPUbK0L/21ogs5LYi+uJR1oJ8Lmkk1LbOTvBMLBAixwAyJ2
cVPKCwf9KXR3x2rXFmxUvNJR9DF17sJJ3Jn8rl7qMW9KMYVrNv1rd5irv2VE
COJR4B7+QcAu9eY+QicFFKvGpWp2swC9o9hJM5SfKfp8HTMqrHij5lTMImF1
NFxQAkPyZ42KfQb5mYIV3TlZKRVJiCtmdrSq6kPTHhOYKmuM5JWBTxjKhZZ7
gKAfFemyb9xunZJwWkxYaWlaC59LBjbdbYJefisX9ylKA4NiX4iBxlYakLGi
1TuHwf8R6oCggzArvDJDzMuDXX2zvswq46pw+VXOx1OU8oURM1sQWlu5X5ql
SOSuUBOoNYAk05cApcTOwnEkiU/YlOP8vf/HwzRn6xDdeBnYQUlZBcQbNHfa
yXtRYK+Gphhosys2TKA3cPnmC2xxETX5QR9oQmBBAFG/7Hzys+qojJjWMVKD
YkoMtOgRXFi8essIZQyGPpCmod6BD8DQYg0T12uoL4p08Os91L55E0Nj4LAP
VXh8YZ3SkyfoD/fi7sjMUrbxsZuQ3oEbhJbUPNtwv7hqL/UZcX7jCLB7tm8r
C0YcOCsEjgSrhuCnH1tscb8tjPr/N+FDdeqW3htP8cdeXbrpjBCPH81mCHoE
drceZ5U5jrbyaCN/drid6atF9/d0mC3oqRH+zF/ucui2qXloZI5+WZrZilRp
ch2Cm24Pwg2rOXHvVrJFNlAxtnd/Q6wibhbEk9KoqHRGt0v/23MorZS+eZz1
ihTh6qAaEvdKqe3lFIk/g0eHzmIDTgj9C3SIMIn1iWEZr1FvbPhJNJ/89SB/
zZwx3EJSGuVdT5F2K4jklp8KcpWR58KbPe5kL/gq7Tn8Wb5gE9abeSeneCMj
DHcgOJbClsCORgsBTss78cbm8yFXr8ehPapwkyTG9NVjVgCsrsOVgdUfG0Op
+GvbiO/XSHGQSW6vIEo/0RtMuaclqOjewbnEdd7mz3lJkHtKZIc2CYp6T7tR
qta5rhPlDSkvQmVADsUMQolix1G7OlcmR6bUwGdsdn385IS0q8Kix/BqM1H/
nH+XscbTk56UihzqDuq09bwt0R5a1G/YoLuhpvOFq2tbN6KA/YJQpAWXe1v6
nGiKF3zOggr8E+6JK/rEKlzU3BIdsoILRyhd1g1NBiTmX/n9lcEmPBryx+YR
4Q6R0eoWZBRaJ4KDGZtxL0C+fkkwBL0e5anDAu+acnhgjSC1vYHGX2N/AEwp
FDIdZ15/OEM2WiOderbHWLqIBoP+ZvRHYkrPQK+p9u7DZye8PsoiggC6NQwn
kkKsjHYa+WyDEEafHAL1lOt4d9o4CbwZrtVfbIhXOlV6WqEP24Yo6Vl6vGG9
sq44VT4TjXKMkuuEc3HCuTWNZh8TU6RJ5yU1sZAgD62bb7iJIW9WilpOkHzt
URTmJ83kMWJsGhlnRI8MJ7mE8keUu4AYxFAGvrriRx6K9Fu//8FXvGV4PydJ
nl0o/hagtW/I3YZ43XR0kRya9jXSDT6a5FeYOpDfzZQgOIBxPYn/7ztoRweC
kPD95kE5hfTmP0ivE5LpdLhpGqIaSxHk6cW3jUKK7B2bHmzL9tuk1nIZ8Ot9
4uSSschecaxlK5aJdUrvTsOG00EhRdf7/81In+YI0kHOwuxowY1QkA0TTcDP
isYf44Qo0tSJ1wpFJ+Vyd3G/fmxra7LE3z5scfxxtS4wqR5iqIoVRtEafnEu
r/ey5ImLljR4noiMsg7OZKolmpaMC8EV8wtdTrrYsA5fR1+Y4UbvIYPwS+cf
TaRlePFaz6nNEt+OvkFHW5+I1OBuT2LNlVNZQsEE2VQIrvbM6FrE29eR0aSc
J/VfRoTDqiTvKSKi23yCauWgrFaGfclgP7/RocD4UmD0vL4jYd2Val55t64k
7h0QdJzrQoP45vZxenXssDPwcWNJ7tavHTohTwJipUgumNzcV7Er2TyFK7LG
U81wwM3+WRMYkCiVtCwJ51o9zvPO9JIr/hJ7ZBS+2nb8sB3LmdZW4UKqUwBc
nH5XfA43nUYxsnZSMKgFtbiqiBQkDWNYt5YGCWgOTKW7Y62KUZimC2EU92VU
UeliLGtHUFg7dCm9gZWRw7RM4lRMge7++Eq32fjgnZtt9oX5SVLzZPnHYfd2
YecKP1/1+3f4nmjKUFAuJiKi2gURWycS+XqJMv31h6JmUc5wA3gWfqMvUxH+
doSk1mfuqL4joTv7Sbm8QWKkXxXjwUtQcFjGC7SDAeobnClGsgGGjiR7SaYM
oEPzf0p8LwS1lvRVvK6y0LGWmCyNyAob89lJZVTWxbss/w5wJFR8/adpYwys
XUUgmCA1gwzSSmYKz9GLPdtaGiwFiPPc6kXdcIYO7Q6c6akiEgc1mq65Guis
FwoVnfF5au1z0kh5sEziwwtwjvtdkkW2OLp9YJUpSl31JXatarZhLBuoQ/Gg
zp4rVm+6Q6ms9Oou9PhHG802hBW3h+tggc5ZRwbhyXqh4N+1RCTHlnphajE3
+xHfq2yL8fW8st+bV28ssozFyEfwKZNWERiE6Ch/ZqO07rbp9ewZKasK5F7m
g2y0JV7D5z+DBwseGMQmFxMwOVwRli0Fx6LwB3ytuLDl/Vxzh8+R9m1h3r9R
tH2SZYWaC+cKCrHZVPe8KcooxsI+TX+yMbkGSjNsA+bRsE7Ek3i/bdXct9Ma
Iugbf2z46Guk+i2/R0HW41hFrZchFp+jkAnQv//+dyBIcu+Fp5yDJhJoXUNF
ffdZb/sHk9afhQIdgi1iKjIZ8LlcR6VLnRvlnnqxZQ6ByL9iKWYwN66AijKW
g7AhcqmlqR3N7Q/6qUr72MY7Q69EwNNuuH5+FMpKIU2y10ZvWSeMhPCyAmIy
Xw0iBElvxx0c7gmBfrbL4a6ACtbwq4DpXt/zXrjmyBOVM58/c1Wd0cYgi5w/
zbHcN0ygzCok9Itw3QktdsKtlAELnAYEFARwitLceM/Gt04kHgCEW9RfiZU2
fYT3Cq9WY+mAfv4oSeGMEJ7HDizq/6lL3mNNbcPo52eGDLP8p0MqB3gkFl/R
ProhuVp+Kvu2Z0sY2acNqiEE2eRaBKQM38KxQjjhgPa4bXjurUcFLl1aP2fb
nwYkj5TJdpUpCvp9QORnaudE3mWhiih1PcBB3s2UyclWbHBclHG5Q1UoIHA/
Jbr0CuKevQKmnizBce+V48OtBl5hpd9zRGTPIg5KBgN2fi4JeWzs+Akiqot9
la/TwT01lbwguymJE1+L+KPjTPrEpVRxAyRpJ1ErfcU+cegB4Akww4AMKp8q
i+kbEQtYTKdcn2Mwl+/GtID5sMbOZPWt0iuBKl714C98NiXr/YH971n7v0tU
zK+oa+8fAAQVCDB/UqsbPLkXXjkMXr4jHyEZWuU+/2AXvzvVGLTeNKVfKC3N
JNQOouAEPaaAwqGagDb25+H1UNKYPgd18NeBUropX+FUNu5WcqI3CSGhCM2V
J2z+CoDARFc8Cv1zZKxxrPzjthgWx3w2HScbsFIySt3cgujyzLZ2pzDXWjfj
PA9r6DYN/h+RMj1HQ+xocx+fTumue+umE2tbxoIhKTzPMudd0unOa7izXSyZ
N3waVXkSIM8YuLUyhqAmmp4TYH5KB9KhpPA2InFlskSodbp+9AIhq6h7SLu2
IkMpNCemirHLrleb3W8SZQ9X4GMjqOO9u64aHlJuLoqYq0GRpu+OW07q3jQM
8C6BDxEeXrCCmtWC1np5Gyzi21F0Lcspr7gWLVzzVhgxQVVwCM7DC6MWOvFD
CxEEfB7hNzEQn1ISCr238DQxymOw36cYlF0YyuEEDJxtgWpiPV4AQkPc6aqI
oOrezMpfiZ+tvSyrRZmNvDwQDewdDO+OgeJXg9znT/JIYs01Vvcq6z7tLzpv
0AGRjFSF2oI+b7l0JLI2qZR2iKlR8sDz+3tu4W4BxHtLyPigQvkFa1Z6zjMJ
L8I4/xkKllSTBv+L7TjLPEYW2gDrBUGvlRxIoEoVyEINVvzhQIDksHF50gtY
cwxrtx3MgLSnu/0zDST8qtqcpKkp0b3opMCUOy9ku+lCdEvo5155+DeWyl7C
eBfWQtBrgyu4j77/3lYnIO2TDQ/LvuTU2V5dAf5xiJSc979BJYt81xkwnrSS
fqK+EflzndKHE0R8QIc8XXeEqgsZhsa7PKIiSWUpHpkJWfkB7Pwq7sOz6CFl
3SKb1/hxDuE6XiuxNkCsHhhWuxwVGWL7hv0g7rvGeMEcLNlUTlBzgwmsdIHk
T33fMn8MCHyoz6q78Ul9e3xsob27hYo3rvtnQPePeFfq/9rXPSgR5FeXEGqd
0p2krOG+OoLmS3DXad97iIgTa6ug7tCap1N8gC3T2fTa6JMeQp85S15M6kl6
mHqmtVjzJ5j3wGb00ZThKTeEZm17zlSVUJWj8/ZX/1SVVvIwGXiItnMYbXsM
mCz1QkwUhZiKHwBCXCgxIw4EqyycMuv0lHemd+cHllhN+GtaUgqIRafhb0W2
IpmEY81jjPqTsZJ9eT2tAMQvvw8g7IckvmT/XkjSKRJefBaJSBUNn4ZlmlBp
tBPJV5qKpOcd0SgTU7SYfDOuZci738TLxFHmdSsT/6ppBWLSeJaaVPHttDEF
v/ZoUd5YnS3BxMUjaudYafAJvcZVhjpVGP5tDVA2q5mzqM+/184LQSRp62UU
4W/BMvIX8jDB7bkDRRky/43P/2BJnCCDZkXZeT6dvJHWP2z7qmc77O/gZqYM
q7lvpXpFWCFE9und1KgQQup9ELDd3giM3i27WhGmnknX2cZja5szD/Lvh9yj
ud+xY5VoM+e/3HnfFpbIm8bw33UgCKAHO5VeGqPEzsNEPawlgppLPhZGeF0u
vkJ241ehl95iJGCrnxyCaJw4JN24usNJENo9dtxwoYGkGvrIa+UmBuqHN0ZF
Q6N44/O8ys4qqOp1qge+vBFAIIqGxLyScJW08oVJDsJpaJOel55ofSsSh3J4
nhqQ/clFqnZNkeif29IZOMuiGXiBY514JtR7koL0ycUQWXIqC6k2butDi7QT
o2hiaQbzvM9LXjE71hXhhx6uexPzn+tImlWWmrwrVnRB5kaQN2LwO34RXeZq
2ak+upQZzIp00POyyJIsqij2IuiHGse1P0hOH1YQY/X6ChKw6VU8wIv1Ij4z
HjBJ3QTPZZoGizzeBym6h9DIohvvfX6Ru+LCSIliNxvvghBmFEKbj6SL3qGz
kTMGF3UtnMgH6aPObG5yqaa8NPmcHWbIRY6Dyz+6QIhuWfxr63bARHKEmac5
ZKfVg/NoMu1Jpw1GG/Az+7ez3gwyb7Vn2u2OZ5F3KE72UTLpwvSFqZCPkDB6
8ZIS3eqW8CTNvD7AT8wRhflKgYEegpZOt9O975EhRL/T5AZa+2gwu3VVGV2g
reGn0VJu7rDxk68+mSQ/Ja/pUrA6Gd/KN7zDqnzI8Z1sBZF4misFWY0Lej1G
tlzjYsa1jOACVbpO4H5dnzbZ4827c8Fs7Y3QNCw7BSsaFuvNL0JFdogN9qTD
NigymSA/g5kuRAMxTYjFxYWydvGA1cjGeez40GoXn1jZeDg5U9/p+mGHjGOc
lyNF37OJt5FQTtBKN8+T/gfLZ28X/w2Nz7eoXRLoMuJJlXcObIXrxdrJzHNH
g3vA0wopsIgqNjJlzf41ctURUNBfZ//6vwZnUzzyzx3QrRJ+jw/rmFvmjkAy
vxMGN/v+y8ElpPDfKrNzP0uHbcXz1gEKehNvupgj4J4+4w87asxBmd0iGtWr
icrIEypj4dpAfDANIMv+EQ6KwkRudSoKRRdKIeZvv9FEpiYSHSO2tGlX7kjl
+MtdvjcfuHHj9ltdCbG05tghRnxkdvNcpmQ9V59DVfQVxgSz09b68Pqrm++u
2YQmssPmUuGZ0ASqF4QjpBh5yJ2kUeT88iB8B9zzzk29wVosGr/C3bOIAMdA
3goT8f9toFhQOzqFZn1Da9+Y5SsER+5Ih8lx4ifsnCgwprU/UX8TDeibJPBb
lUkzrNbq5JE9qZFfB9zix/r89vmGMvc8t1Uofl0upMSFBRPLSmgyO0RaJlu2
TMMENGQLdkeLO32Myzukw7EECfJ33zawFcbR1d2dP2BhPoEEnXDO18ABrj/B
+/jch+imn4YFvvgUWecBTS9Qwdaji0+kt1OxtxPn1UW24xVbm9lfKKzn05k5
b8Kty/tdlcJSt9BN1jkAz49zEJbQPcyJRhXgd8eqzYBBJfvmeV1Q3RJF8LWR
yx6ZiYe6fNsJaMmPMhPGhSQt9zep+/zpGB2kF549Wg2NOpwUK5VT1DiFKfA7
Uj2mNcCt0zplcKIZvVuz5QAF7/mMgeGU7HB+SzCZ0W219NXecEe54SuYSL7R
YB1zc9czXaUD+VN/bH4Eac2GU2/BPDdB9hE427mOJW0zxilCnLKIVJRjFJhH
Cfg9q9ZULW+cgNhWucv42RenBkJMoTXjEFyPKCVCB8ag5897IDy3y+Bo3Ax8
2DlUAlRH7D+886RccjxA/H7fcWtJ19xh90sVtBfKTDhSVieQUr7gAtcoLT8E
CoHEWrWaY/ORRnNm3wzgD7N9Xfrvr9w5esQRkFL9hjxL/mBG8JZFnNlRCscw
qcCx96FKShFCZ0xX0yeYLOFJn9cd8F1T3htUS6h+b9QLk9Tm9Fy5PZIkOWQy
xwPxQYnXOMMb6FW9qbtfM5KXKC/ha7FNQFNVE+SJfyyYcMxUYfe+42DgNBN7
d0U2v2MsMpgfOXcKxHzPphO5yA/LqSL7yN84BhOTj2WTd/LRLc5eptMCo3aG
cj/+CQQj8ALez7o1D5f24a/CCIE94g293vYn2yFhzc0m3Chykw5NQG1jo5BU
mSmY6YKpgB+t/Ec7zvWJ9W7gbwIRCkhyx9kcnI3onvzN87yR0s3X3pGN7k6W
pl9wKH8DzIq2Ea2UpCK5g46U9e8FhWP/vIhnwj8UYIyDn0bdQi+LwK2xBpxf
rzd5Nu4pDuJWLI/OSBuQajKV6VPb22fwtVIWz9PZv6V8CD8SjOGsDzS0+qjy
DNl6xK9GGGreEJ+bbsjLi43Bi6oLi1GTRlQ8sQBhDhBhuhCeUjKOS6YPi0Ac
kq7pRG0QTo1GItFkHiEjogdmqPOVlDM2fuO1kLsxBvJGmeKbGNSQhWouljvn
fuJVLOF2R/yqlytiKPfpCZNN5jZsiF0MCiSGDf9GqtateVKV99Yg9nIVwf5L
w1xVXqNmDvua15NC0Zf5Qv2HnobBT3qiV0L8deE/wqYU/ItlC+ZQGXDa6NFG
yMgIi0wHlo8dLCjmkUFZexMQJKu6YYS0auC+M5bFE1T5PtWRBi9SnZUXT+sX
IZ9UhLHO4eTEhCzCks4WpwuyVoe9NCT6TztB4j5R+FT1wNrtOldALC0249Op
NcyuGXwkIqz5HVJV9vWrP8EngaOIvZJVTSiP8/Y7XE2+P5nr/pBYHRSVWOBy
P1YkHrHyh8kOL8Cio9yVRU+RAij8V8yT2c0zFbd34YIJAyKS0y53Oadzz3xP
vSxiDgNoBd/GWXq6FS/kS1f4MPhe2ev72k5Nf545wWKehF1bSYIuakLwaHpd
a0PibRtgz0APiFY4T0gteN70PELNMLKWc2K4ynEOktUFu9b8+922hBT0pnMe
u2dldgh1qT8dxHmuYMY+fnRjQHQEcGEp2f8l84+QxocYhX08CKxW7QoLl3xm
28PbClHPprJ6Sta/3OC7hUDYRy1trfGHjz7ncWY8cp8JvTYI7HJOHzCg1bS2
1dl7UoAIGRWYp51juc4Wc24tCwaJqeA7LIKravi9y2gydRBHE4+48ZmDhWe3
rInppBvPNh3yFXdAzlj4afR5JuAQZ5vXhu1hIpdbvGQ9wLiHBQiV+I01QwmG
QsVteB2ucDkt/8ACaExWrjiRayV77p827xOE9DgGLCDXebu0OpzTGLhSjqte
Y8jGr10TuTKWGmsBdQttwcEiVLGpOU43UH13CzRJ0hwZHBpWAFmsMaJ+oguf
+yikf/bzUwr0r+dMiszcRr0xFPvvIT9LTZXUdLQjDvCK8oXrz60WsAnbqsKW
fnBk0O/XJjiQ8sdO/pGpjzxcrcYn0IXpcyz9sGH5dAHGLpaP1NA9yXUxtlNa
g2nK+SDZl6fiQ63OtweIhmwuw4Ybssvo8Rawp55GYU7AaEOazsEgsR5qj2Jl
lMK25KG9Pqj/98bZeaDrsgYrbBpTpFPofp9VoYGL0QoowYD1GfdGmRUq+DEY
NYx4NQFiKM37vzIxYTsEpi5biD/pBlhEah5EYIqesp6yrYutam32lW//xTs8
F3eWU/HH/F/GHdlR9+w3NByrxAo5/8xtTr89X8VQ9688FmpV5oMoX5YWMLx5
0Wi9Cw8jWBCqvJFqg6df/OVZfd1KHOgrgV/cLZco5p/pdfwrkJ/7du/q/nYS
q38/K8M6OH5/xH6nu/U3JvIzYWh4XtjpI1VI+Mexr0+FiWQT9YKExZ+1EIDs
No8ZdHlBkVpyQI3VhoUe5yy7wyo1y6eWRcIYPvimrzaL/jvB8XMtzcn0pVyj
KLRq00ZCRkqrJiyRRbhX/n+/YCZX3YI45V4kYxz4yW+OlbuJ/BhpnK7tC7kB
nhTBvuSFmrjLCmje0jpga3Af/Sb9p2VeRzeSFU4FH7So7VcbT3p6w0f6RBpt
wd5eI6vLz1y92JSt+KPqsiUwEFSpeXXqvsnnwN6LbGHvXtsV1veahDK6j1Te
YTMg7CWvUh7bQjn3b+pwVq3/rS7WFdGOl8fswgtGNPmANwoojP641IN2RIO0
hvNj7EAKniEDOou21mkJ1hWeimOrckjc2JSisndiGRxyQGDQSmaey5NqP17j
TDn0P3MSTcqbHhkjz6TkkcCsWGNHQx4MX7d1EM2g9y6YCu/7zKcTZP6w9Nqz
InYsTAXBgT6NeJe9UCZqc8zCORyi5QLMm6NX33UsG/F2oxWUtN1rdijNg1gJ
lCbiQOoZNOg3GelLNAHw1qxY4sG68XMa5/gFJ/ckbrTM7ULmFxsCzd/XzIhG
z3tR4IAjaj7ZRLlygQkTEv0S8Jm1uXz3bL/hTXh0qA2bdCvln7QNlMvp+05n
+Bvrfi5tHNsRDMe1Uqi674HNinXpwzYB6lzcpBPYoL5XSRVf2IwTy0PITf3z
roLbv5lROGtk2o+i4Jy/acdicDCcLPh7CI7wRgK2v3t+1iVva5exfdbxyCGu
nyGivJwio5qApT8rAYc8pssm4DvwSH9WLeNp/oujm553k6SDuugFOMSU8Cq4
ZUe9BRZkHlaLHZ0FEn2XuE5+GO/fhqhucxdujaiqEgkX43AiAFgpcqr/Bd8/
SbJ5F3LLN78XXxkrhXt0x9ay5GzTm80ZgRDlehPKUhYGNBpWb6LR+PDPjfjQ
hyNv4Ww77ymQFtReB7DhkTHR30upE7uXbGHes5FV0FNbZ3qP991vCSvhr5ll
BQ6MAuR1om4X41pIyRXJGAw29e0/EJUE5Qakk3S96/emuO9omgt0SJF7Z+Ah
pkPRfxZwMtroKBuMZpIoCL7mwq13crGlzYVraG8JX8SFAkL+xXzi8UEsezrY
ZC4bQ9xPH085GPgrbz2sb1nUfs4SyzeBj9k0lKlBxmOCqbgryn3WuyDwLweH
NhfMTF5CaOezdr8cBjPZ1RPD7Kz+rZgYr71WOTxaA2Ia1gB/ED30/+DFFmG2
8dssM5OABdKrU0ILzPq3jm1whg4FU6U7VGLIdRTNdqiU4Qqq83siEb74DqH0
WtQJcPHvby0OUqAHN8sD6cGUv0aQIkhSGz6Py0pZE+uGExtU4ITOclM1B43q
fuyks9PNtiljM9BEA3b/RNBEzxMxnSfWiFZh7mvwvtEPsrE+P6e5j9XFLFWr
IGNudyW6J9UyiTMpGsWoQYBHZHaOa99VmMLppwW4E50zCmXLdRhjHsm/MbkI
uh0wCbIJCtOKrNHi9FDWOvKwqAhNxajTJiVRACzDuZY0In9Paq9mKwf4YdcB
QCnsFpk7PDb2+tbkvvvRVtgUQFr8rHvZ1oJbWIl9t6iud8ya2RRZVbeyrt5K
WW7XwAy/Lojk0wNLcAn4kwdsLnJErSGneP/uKmRbqukysPDnB/P2dcDAojnh
MVNuu8+3HPam1JE8CfTHaIHRUnKV+8AcICifOzvqnRL3BOz7hfqoNfBqSSDQ
PlFnrlK3QlrM6GvWwlmh+1letG5ZtKihlzSiZf5nKLWfJF1k1AHLHFFv5M6U
tJv22abiUrTvZmnrW8gNHgj1xB3fjMKGkVV42LoDpJJFmhMx5ujJlA2gPHcv
EMk2FZ8KjiOhXSfhU52rgiJp+1UpWSAgTARVnPnuZKq9+RVhbFqJNH92WrYC
7NZCaIzzlc247ScEk+WGD6UdXjVEquAlOJW62zdRR/Z01CIOPAwIMqVP2Z0I
uKpc98whJA4qdr9jvWRZmhVBrsBJ570E1Lb/zo0/8xi0MjIb86BFw+4CiNAU
InTXw9PNB+yXtOZ5O3u7tLFp5A8V7NYZ4wLw6K8dzTbr2zTZle+MbvK9PUx1
LhWj7gyraFFQow18du5D8j/mZgKfGKfx+We2UhHVdhjULlm9ArREcjihsSII
GAkhw/up2By5zCaSlnv6AgNajNhBMwVA4/ZMJXByk/o6KLOiCq0iyyhj2h/e
3/1VQ/8BmLpr8gnHgeywDlGB3v63Iguwxd5ZNdVCQfWy8U3+2nrJAa2x6Igo
I8IvkGTCMpCKcVwrarsL46IpeseF3rkIONLukwIOviLec+C4b1kAlywkplWJ
9TpP5WIqe6DsLC9C3++KzIQ5OJn3wl+fs/0qkyCMtWMX3A1ooi2go03L0+9G
x5Q+bI/NjKV1FbULrZaLcq35ASM4ssCXmcTFd5Ad5omTv5xgMbu3zIE2lMbq
JopHaPi84h8R0eHQCzmq2btaTacmxc5I31FM4do2DWq4wssJ2GrjJwYMvGuk
hlldxt6MTbFf8/yyXtyI1lZYm1cjL0feXCjVLY1tst3qjcKhYN9VvxzdO0Kl
GBm7Jr4dbOlmcU97LHUFXDneYxv92hLNCNfIKm/OqQJPZhUX0zC/Xd+7J56D
N08F8BNg3RygPraexvir39itftml4bWktBc9iSjU24CcFCScV8E00+TQ6DMO
zYi55j7ttRiVtjhDkPveq6r/koFCzRZBbKcMNDcvPIhETLMh5yfVhHMYHdFH
/xG8wWnipFZPjYMp7HM+q04jwzRMKeIT4fqcx/rQshXpbm7wFEyhECNMcD08
moU1ewovAmjkhH1CZVBYmL0b8tPbWLhFdCCSUGc3V93lHfuWM76sp7GRVGl5
t0Nu48KLyxUiAgXi1S7XvykplW30gmkskspTx2jLLaS3HeSI66jRDPPJ3B5z
xfEue16IKWPS489pteEzJL56t30lFpMOQHVPIwJHw0DhFL6ow2DsxwPrcF/Q
4pCZeuyjQw6ZpAZi1BLp3QKW9tyoFlvCaLkeRTkrhlNdWSrlJqSNgcEfBkHn
KZRZg7w/CNCRnbNoSHksl5Qqpe+ukTXPrA/wVoQkCxampXcz/rYH4+fT6/zu
+tlwzFyGvyD9O+OX83p6fu0/NBgvxOH7CsyFba/0XUOHOhKpNM+00/G3vS1P
+s6NUhQtR1sipUDqmQQPfFoXvGH4grGLUGPN77tP7bzfcqLRaa6//vytWewm
nXFTM5N0Qt1XODbKyxTm0pNzWc389nFOCcaH42aGyvmfsp3uSGGvjZLC4PRD
NdQ4PIE59WN9jUpSBtA24btk5j/xmB1OCcvoxhAzjTUBKCiW+/trSAf6yqCV
OC8Z8Wu+0CDXsGi+P6845DtiogT1vemaKtxtNhBxAwJwPO+cTUTSoh8jAKTu
ABYGwdlIwwJrKaptJkjLyGhvs3VGlJcwPcFGi2qQ3qeGA0SFNsJbSqYJNQf/
Q8GOQIVepMcyuF+az2Y2Rji4LGn7pNr5ACg1y93tECx5DXHqSsmhfVKOeWgZ
zezAcJWf0ZIsEBATfEC1fMR5Vr8MsYQuSS9BovEv7fiCKRYX+nJKwU6kTVoF
KFpdAyfjMUkaZoF2Zxm6KQxkn2luiedIUR6VkzSgCGrtXswqbuaFr6whWIep
4XpFCskYpaxdEkwG47q3yeuaQunzu8rShR4MjGVRrBtLf3IY06olWrIU2tfT
s7i8ylLfemEtrXf45rWc2ig5r7MiK+99nl9WY5XVS0eWbvpSBb1aCmnqNr/b
MCygq9Dv6mMPS3M2Gi3/Ic5Pk/f7DfmqIGpQ0j0dtGuVMtsxO3+J3oq8QaYm
jcbPxL9o7SsuwgNg0NJluijn7Z7AzDIRFtXi8jis+7rURS8SWZcYwEcCEMoK
uomwkGzgB7djS+0OswcfDjk0912uYW/pBweqTlpJtl/Mi5ar9W3z4E41nwNq
DWpo0+80K80bFs6qDUee7+dWj0mkzsick/HYDR9w0ZqHgunDtRh19zoZU3wC
QP0GMysaElsjJ7Gd56fwf9hzU2cjAEwggH/9BGTG+mLoTGPO2VzBgRLBJuxc
YRY5vWYPgLWMk/7NSD4GXkWJFLtJatsdBkPz+yQZ+y3UHMf+nGUNrsJUPADv
NoUxm92OmiMLA0VIfPyZ2AtXjqRdrFYZQKsyLuH6Uzd56wr08TTX1nPK1vqT
lHIIMR0rdiBOTB7l3Bd9U9Lo17hkxajB3xNeTucEeQPLah0YelNid6k+VkFA
20Sv9n7o+LeVyskxoIwx9aWhL3E7OOp5y+kcuG+6LnUnRYy94Jh+7DBjc9pI
JLU847n1MEVrTbUfUsisFz/GSEiSewiJz5yIA9LdX9w+jke89IFjISvNykDM
m1hHcKz5uk7J7ZB3WQpoY39O5Q/60TAxYgEASVUB0m37YDb7sXRBP9XgVKFp
dNspJFbl7ObSEStxpmEvI5R44FWUkLOutJ3TPTXa8ZvNY7NuQ9B7DKqzRO9c
MWENLr3OzNSMkVmY4AKxBR397u+l/WClHcUUXUWGlHm7FPJpNVSFH94fLnKK
yzm3li5YTojwj9jCqxtdcIb8QslI6pEZ+7i7cuCmcP/vMzX26sIhjUw5US2D
fEBU2ik4Tl+mjwY5XIXheUzzhyJWsgZ+eBliZn5y64olzRlkHLrw3SbJmF4L
ZuRAHzbkCsBwDhg7VA702P+hwYfhDzSI+6Cg1tFUedYUw5shUYYx8+vvvlsD
AVbl09tpg8eAZvnOTBpUTj4OBUztzF4zAk5FeH9/sluLKkk7O+jjJXZY1oo5
tRFAE9hKALQ18IlTei5DrjhAKLU+n24Qmd7gLylDv2kIYlwvVT3SnJWI+Xqh
GF1KMv8Eg3OXw5bMhGQIC9DMLH261X848bSMqlRbTe5HlK3YGGzI+eGRXUQe
vIZZZQZ5DWJf2+fw+xCFEjVB3uzP2splNaZVbQlvhEwlnKcgJi+3YnJCvds0
6kshlz3F4AqrsOmA3Yab0Q+qTSjwJ5oOd0Yc1NqVWIsALLoh812U/whCA/GR
i+oTOahZJ4heifFX+kzvDffnSMdyYOnAtUyfDE33Sks2k+uNA83zLuOg/uaR
BUCeQEL8BbqBQStzcH75Olrf1wbHXupAI/Fvu6ePiu8J0SjuK/3+nyyj60FF
yw0EKQ4Ifse/Hshue0LPtr/XwKPDLv3BCiHkdzbVN0182Yilurejdzgwt4TZ
wIkvLhFbb95LFu9tzoXcwcHXyc0U14EV6yTITjT27Mvs5bSIMhg7pOWbzSF5
SWbhLYLI0TRx+1O+u0mWcfa8a5PNi9ALkxMVa9au5TTNnXwSJeFS2wG0fgNg
Vm51TSIXBj6kJjLQTXIjo5Lo/70Wg+8ntXno2IYSduqUvGoMNGDJH5WLpkig
GIrfnRZc6irG8PNBHS9YXpVzzadzZVkx+xPf5I6JQmTFR3XeCnflKmuOdZMM
18Icejh4rTjm3ebNTexD0dPt05k7iHZxyxXG+etIIn/9VVdVGSr4yMA1QDTJ
X5UgCNltcTCc9HOBLOedWIYCriD2LGOz8f9W5FLiz4Iyw0d8hCYNKsDAqNZG
s86QknT2sLOI7OF1o2x050723KQLOcTd4d1l5tuGlZkTFXBOKH/HAUQDl53Q
KSziJFSAg8VJSkDwEgdD3jUun94ueDj0TjgZyRIp8XinitB51Ca98j9tq3BF
jNlCHqH82HkT85+19ph+gSn0WiETmu5CEy8Kp/+y39DBBZUHnE+J8GL01Osm
PF3J2y3ebax3BfvlBhTK7SF3tGAO0VZ99gntDc30luq9iIS6cW8z5ZyGXuFM
a3r1+pPREMZBttH3HTgZ/MqES0s3yQ6zm1WalVgvcnZe7z1H+K8iFz2PTbIG
wp6NKZvAWkOBs4HVrnXgdzkp5SLXbfuAhBo5uwSzQoi5BdDx8xkV0tCZGL3J
pQuMghCKjScNEOzlN9OoqPE1opl0JtNFoykt27LBdPty6zkd38abMIHLEXmw
M/RGffMptAmenMgscQT1N79inLEslsWjPpA+PeXCxhd2i15JXSh1vnI+JTA/
soTUzzG+gvETI4LeNdoSL8qLw31gULFfP4BVSm9IRDAvYn+LlcEeekMTtW0v
Yqw3ijAxdSDI+x+9VEUX9j7UsGIUlDVFyz4qqbqkjx8/TgQ0Ixx+7UZSncJx
1Fa3YqjoHUei6q9+V7uJczKOZSd6LFS7e5QHcBcUIkDOe9p84NiNwN5nptm+
41tGHpxtkt308C9b+wHsk+v20KyVfda8SS0FKD6jMUG1A0BrZ4uM8CduaS5e
PdTYO10+DuxgpyS2Nj6G8q8ovB+K8+Kc6PynKT5LtEWHyzmW8PGNBmOqsCJG
YANbOF2hDP6tjrzlQAt60IovZ3H3nRnjz3xIl1+HmDZ6gp1SDxB0RCmH9xCA
F2+aT1u7EmHYbsuo5aJ9ST2bMgD2csClLlgglSBd8xlL70gzA4YMcWVXgquI
QAATbt4Qqfvo0w1/WqBmbWbU7fO2V0syCI1zSnZvZiwYxjkqPOBLiXK6pXza
mrPuPL2fFmTW8xx8AKOW45xQZiKQ1i7EGjofn5hjKuc+UdhMDogxRCWnYRkW
sQvPhv085I07Fk6gslydporN1YPk2BD+ZQvy9X2U1oP4PKF39gyzFP9jT5/h
bEWgYJ5oyAGnjqazRz4qcWnAOPimegDGxL2jInoBaiAe3LwW5W7EeYUcG8rv
qR4opIdxruyW5mIsdGnD6iV9BQrxv2gegKZj746YEf6NX75MqP+Q8WpbHCHs
8+0bCd0WhLcUORbJTBN+Z5cfFeJE7zs9RM7hZquHzGblM7EtqCXZWr6YMpw7
ohjLylffhKSrZtr5KciGHwhZYMtP/D+J0ZhSL7aR/dF7eoAb/o4E9bwnmODd
0X2unze3UM2pVx92A/Ur0vSJ7BUWyJnnipyeoLx4EoVW0dTgAvO2hPSvPWA1
Vm81ZLyNP+TXxf6peIvGYFqfrGyAA7gQM3HF+fENLfj7qbC/hXVQM1/vGiIQ
oxVIuz71HXBzTc9+HOIIKWz22Aub1q/7caY8UaZTYkYRxHbxZuY8JJGaU4DT
m0+AnUY1sNpofwuwovLuCOOm83E6uROnjmyqfdHe5ObdoqMfIdbwQMfroLpY
tMRoIOJqlwxhunj0ctHlNnAghLgegOYNvSHvNm1zULpbdanqTxcNi0S08c6/
GPM7R4WBBaeOROBuRFGw2jEMg5MlcxGne93+KzRWL022Q4gwoMNLNgdLL5sQ
4iw8jfr0U7fKsQY05XSAeYNOq0Fzdfcg4xDovOkseqg5t+AMj0Gbye6Eyhkf
y7qNqBqpnMDqfwr1Kq8jP+/AMZRKsHcWGnP5qaW9wtNFgKO+Id3HraUAZTOM
9KolaWve2/Rxqkl6bv3USTgyCQk3f812aL3pYS2f/+vZydzTxs/rhT5vPd5i
ESqMPDnihjCQdQBxVve3Bm7sWlA1ErW2nffWnhUi4bfrp/veSsE8SxqtabYJ
skUuM03zfdcEy8ifCEnkuq/eqYgUWG2njL6WbvUO8eHwMjju8la2QMipIl/+
9bvenC3cC38VouI/shWUlytQiJr7z1ltBU0StOra4Uxjlxv13bYZbJdO6OEX
v4aEuMTcrsZlautzCov21qmbqPjQl4SIWRiAfb9hoU5e5r1DWVL4vASwXieG
qq4jxyGU/JJkFb4TnGpBgR6xX+UyOdd2YQMiM0qgfjCmz4QtJTfkI8JpKeeR
1RzO7DH6lGh9RKwpTqe06b99wwveQ9aDaM1v8Ef1LtieUuBO4xkfgXFLk3Wv
QCGwrmq2H21jtZ/XN455c8VNm1rMu9/1u5z8js/i7OrFsdJG1ZRxbKBRZBcW
pKchvGZFipV4FdsKyfY/Kcl3AdTRTOk1wXUzS1DCh7oiyookFBeBujwy1094
brl3TawGx7k6udMqpBL+m9ixcMAiKe6udU+2vWfwsPrlEkVaSbRaIpsQ77rw
U8zB0XqWHKeqg8O3gLPlTGbEhUh0vjgijoyKRuGkKwu6o5T9/cbID3T5hLI6
iUvj95BCCZO960esIrRkOfh5FhZCFFcWDfYyY+zElJHnA/wNrleY7hK+mSHZ
BBjhzgL1GAhkzA6KScq0vRoKhkrOygdrYYz0RXipJotZIxmS79cNboDV8f94
otcOuIBCG4LLJu0HQWQ93zovfNXwe3RND+xKS+/OvEui1HrUWjVZZzapP9k4
ohg36Z/BL5uTv7fkazTHx4KDxXQsy4VwPyjFduACYiToblhjBuHihLTeJeRp
7X+xVMOTdvfYXJvrGMrMUXjs9rQostDZg1D0SN7fGZiNANl4k4pTVgoYznbL
NspWiHBBL/jtazx3aSqmOJbRtLLS71eXil/gIId36lw9MdG3Vta8gTFuUglh
RVUOg3vm7U7Ae1L7fX+78hgCMrUcrooP4mblToiOg6lB3Fv9R7SNprCJacvF
yF7xTbxLJCxVTOLm2inAuC6z6WRsoestahaAneKFbbmcqTs9C9zdNbcN3ZNy
j7gRPZrGhDHwKEXcaKm49Ayh3lrQ2gN+uVOPZnb+xcyPRcz1IyER5l/ljpJm
RblusmXZiH0M2PBLvsgaFjBwO7hm9DRNeV9G0yd75ltOU2Q9B9Lnx+jHZIuh
hxohPh6ADSrsOSHMYNI1K657Gf1qBJ1LsDVAyNf5lspfuqbjwTglwd7IH+uK
norkMZr8c3O+DyATV0SF2iQUdlA2Pluw9/epltYbJIIlVVIYi3GPoJRgfyCC
vnP88wqKHpumBRLbYIkajyOFCPYVADGiRPnKgcl2WEd4V8xMERo/psyXoww+
3SrbRA74ZCg16UuUUAHGsv4B5B+5+7g6x5M5+yuU+dQZAgg5yvngH8PL3gyK
Dg9a3S7xte9cvrr0cQNXGv/DR+8j4D81WxfxO1w+F6nC3md3ugHcONk7jYT2
TbOZ6oEGwveyYgdcn4eYsdqA/PdtwHOgpnh9ZX4NwNmNuxS0+mcRzh8V66k2
BmBd4X5LtWGO5olV8VJpRdlZh2UibImpsHrce/CD2aUQfl06gVGZ/juiWhK+
utUQHSP6zN8V1fb+uaX3f8/B8fH4T/JcKrJjTaqSriPHFOM1BKcH39puMuYW
Mj7plJMtUgRxLRPDzTH9UxLUS1YaeDkrz2cI3Pz8VADX0pHaGVP6Rcv3MOzS
lZbSZHOLXfxbrJ5KMPH6LVhkrlM3ji/gfRvjzGUsM+NoNGYcgqbilR9o9zmW
FkI2KJgaayIahNEqVUy2UmskxKeWXn4mL7g7y25OH0S2C54hcudsz3N/qWoe
L7iC+AepVVi25BVYaxSGMBtscoN34ffcgM72V75sLAOSmknWR71cBe0ZK44Y
pYrLT3e6sGJDuIRy7JYwWXftJMSZL86GIWKfOk9T9peSyC+3vTgC+iN8oxqO
3V/99YoqVqdmzbmvwvTbyOeipuyC+qorUBgUQiJvTDQgfZvjnW1raZPCb0BQ
qYp7tfCOtvbMTIoS6k8HqgAqxOQQBeD0Oym5zK4RGHwI0RSc/j/v0xpFp4S/
Pmd0jxbl4d/UpiYyVTneNZPWn1EJokLqa9U15MwuHns252VcX16TyAJvz2dG
O1KxGasgk8ZDsHdkDAhZd7aS/05z3WDBsDZsx3b42CXPdqNt8arn+VsfU54A
FhFKx/3i4hXkOgqhb/vDHh1dLnbjKJK/60pnCMLPB791PSfRtJkl+EMu5lUH
1HUrqI/wnqmgVlsc5FDwSwXOS+aB0TbaFQ63VbZhL4KrdpHYs3daV+yqo/Xz
8AHpB6vW8nL43ofC2lta37zruyfj5txCkayPwkSDoiGV3MxbiXdooKZFR2vn
csW9ie6WBLpyNfF3tozrOJU4N3mqU4IA0KZAgKismMtfx9B9oiH7Q98iaaW8
ZGKDWedmnvzCx+iXkr8fMuYXGVyyhnkmT792TgndykJwBagiMmK9i44dyjwk
aYbNFRzMVL6aKmi1EpNJG6rxGQ5H6SB0wMxHHNz1OnXJhNGfKlWfZ5jsIPtm
+O/l9Yt1//gJTDntG7Am47fXqc5fjX0QDchswDeIaB9JhwVW2HgpQFLkaAuN
Dnj5jav4DV/Rsysc9IE4sajYz0y74KtXN+tHaLXMP/e/sXTCF83kkkiHTply
Dc2XXz45yv06f9TgFRkwy3le1GJQTy6lMeZ87cbRIBOJMbDpQ5nIJrZ6pG8q
Z6hmpQDt1IkmL4ldIVSYI/qW40dZG52iD2UXzHzPfHBTp2VpjE5ehEzaxR0C
8UNds82xCeh/hEQSoFoRBKGG39B0FLTWHOiKRr5z89VLU+WiwGuORBY6IPEt
SszV+s3o4rTnN1MoMui/WNglL0kNM23Mi4eRuSm1ETx9ALDiFvtvc8N3yN9c
vn1v9yiIOtNgYI0hJQVH7Qga2y+npI6zSBusBIa4FjxHAi4WQXgXb338FvNd
zqqy8qf4vdrsI/1sCdBsMQloglJYlSZb8qtI5uDHKyIAWVV3+6QvU4qSeRT6
FI5JfQ4y0bA4uS/Lv8fjsfvGzqh3ZDM3L3jErDz7qC559u/ydFo+73iPeyrJ
T4UnzRT+7aZa4clCLtdvmDqSUCJADHqC0JDi6aiQWePZ88r5utGDIZySjlfh
8TC7o8IMOCBhnkNdoedO+D3XLRoN6heUoJ0ITUgZGtkTkZwPPcn0OiSvFnI9
bnpfF3x2Xh9hivk3BGSrNdXJf/D/3eNCOipfxG0DyKOY8YFCOJmVtVSzBd1o
UPl8qpAqcP8bO66jdYbXHKOCxByLTbywbe5Vo4FvZwCp8ZoOqrUnFOf2PTNZ
Ycd3nWxWICGl8aw1zgcV5vQNCmcmV8WoYAV5dyhvza4RIG1Kf12KBSHK7H63
qWMQ2FtxtGuxN5XWIZ671pk1r2DoC/9q5QcOCKU7d6jl6OTXUC4E+m8lDol/
TKWGzdcoppwMZNzNbYVTKxxVOQxV7vx8hKssGLEw1WJn9MWILTYIuBs88apX
wfNHABpytG8HDvee4aVZNR7i4xTf1Ww9Ap+F+pUeXyTxOZRjPpnfww9wTepK
qT2wcUHV46hRY48RwHQkuF9cN0Q7aZltVhjKQCmMOLf1PochqA6NI0I9t2zK
OYSuCZohcy9WuwP09E65UEA1Fn/ADiHaUuPetaTfXolIprsRXIiwzPDfwcvf
XlhfxRx0F36ZlSDx4SfBBBYz7uJ2BpsUYwqUn+bCiEHQJtqQBRqjmlqnpiqO
H8q0Y6Tn8FkKxlfPhhq65dcMG3rpgFm99pOux77nCvGbuIXe0LWW/tRqaVzX
sp3NJryxAQRWpt90DL9USiTwkr/3cMxjzAHB+pJKlg9kKuwH8HaMG1PWX5fE
HUCgbsOtGjQo5q4zFYGfI2VPsOIRf0xiBYcam5WiWdScBqH+0Onwb2S/d+/h
0LcnHOc2jmt5zqpAhvj42YhDFrhvr+d7njjrmFzTanEu4jThgOeDwZiHFmcL
250LwuzE+z0LsTIcZC20WwH7U1PSpuNYp7LNcP4pVhM/g7qf1dzViU9TKjjp
9NWEvFpeAHizq41bn/o5P2lo2R5VmjDcg91Nz+rt6eUrjX9xbXZDq4q9eoxi
ZcFSsXnk1nR/TYY6NQHUphgOoPIEz3FxhQnHXA0U1PhFuJ8mtztDsW0INqSj
DRlWDTK1varunITP+nqVc3HMny3ftHlg0HMXiUO8VyiO0o611t7X/ktdHmc1
ukTJoQdJy7ktkFEoA4kR3FHOHbtq0udUN5XNt3ze8l7r2RtS/qtfMC+BE/Bf
0Ww5SEwuJS3lksHIYfTtQcxFNDtfj1ZWgm1McEpanyYvwof2Nb9o25TvVUSB
WFqA/cCtsKtk22ouTWF35ig/S+IInZwdAG1hSiFRgNqWuWeAPrUGgB5Ca911
rVSjHIT01SEw2vrg3Mn5YVt+jVk5GdQM4s947mcU3MlbgGoxVbgx0ifmihI9
JMQkZEzo8xNIVVc2rhcl+thbL1N08OVZb4biPttS+eNnlTeTtB62IO9NIifi
0WD7AdfMa/htiRhIudNB2VuqZVucgRbGKhkdogDvLunvR+y2xGt+ZxvTPqFQ
r0SkSLQYy8akRRjkVUYAWdnDMzZGPCdmM2zE/fZylPzJE5cVQgeHc5GuN9pB
GRV68I4N//3v0/dlnGOBGtKpGSKXiekRARV5qDyev2qSasrxBYvfBZZoKt+W
JRJ/Z3xIQHZuyu0oySHh5DUakKsJHoLgX7GxFIvFDZKMZ23l9q4oCKOv6g56
8mktRlL6UVGmoPfNN/5puEceJyUpIgRBADGAfF1HiGHtx70nUoVIDGPhbbCd
vtwTAnXtNxj+0bbzbNy4GS6nAkMnLDqJT1k5GaO7IX+HD6zU3IY31Cra9xkn
D8TBPQfH5AfQIbDro7vYpjFlSoK/lFWNtAdVFen5Q8I/xkIgN17SuePkskpH
NbY2QhXCYZ3qImqWWS1sHScbmZYQOszqEUj9wq9T9x+oEPwrYvmXldXmCYIZ
zhnupoSK1uuvqWSYKEcr/kHn5wIGIwuKhO6hj44Q28+psUmBNSyvb7v5qr2Q
zbnLVqqS0Ttra2ixb4hvxAb2tCH1OayxCpSq/c3VZtCeKTmrsPKdNdS2yZ4E
L5XeDRk20n0AR4m4yCkZXj36RSbILMWgAblUlySOVYVlHzwV2gnZ07HGsyQ8
Hmpt8JkVg98U3IdWrLH3PxjwAKjOkX9CnBoVrh4yjwoHclPhzandnl57qQHe
SS0bCz2wIVQVQobNSUDzB4BJmnWXcpySnMEvO3zzQG840WKbsRV4EBU8mIqz
LVFDUpkoKBFAe+I7sSiQGJLPRy+JOxgILESQMcoiHu4KGxGjgNQFGfyAy//C
Us1dQzxvpaAq91ol2hCx88VUfcawresO6K4dz3yRYTsh+FK89t/dPpJ952wm
z+u1x/YQcXSTLD9XoL3ZZ7Ihvi0fvzYOvQ3602OyRV7IW0LOEiAx8X8ixhK9
AhHJPnXRdGA0Yf5SiCJZuUPtERjQdfgpjKBP/8Xpe2hT/7FIzPOrnyfn+7tN
IIb6E5vqWcKO/zLHDPRKFfVOWIn61PpdhcWIHWj34Sb/81l9YZOCd5/jgkhQ
gOD62mJktIZmBivivfiJTTmx0Dztn7Z4mhE671uWcI+w14nYvYmzqf68A3pl
wsnMin2+1XnPMIyGpAS+R+UqUERHyxeJQiXltIkZP5gR66hznrRoDBYKNJ8a
FmPflIZJIwKLyNSn5gAWht76JQVRPVYsyEIe0cV+tfc6CPhFGqEGoc9/ZSdT
ZPfr9H4zMhvWs3ec5W6aAJCdd0IyJ8o7VF3kT7nSROBK2bmr1u9r3+O0Qrxq
enC1ZCVPcF837bDazYe6QO5ldLlPtQcsHOQGvrLZZRFasCqI9HJo2Z+HSfkQ
5IeSUA99W7bXkI47Q3Hr9JsB6RXtOcrDMfbgJ2OQzFJdJiAuJcZAEUcmIBo7
mctbhlXPgMNqFsDc7JjEfxUueHbmm4Y7suE8Lvad8wNJY8/Mjqhj4b0vGrcS
6rG2do6Iu9FQIMwm+RMAv2UO2hX+lAnykzeYMhyyJQXR/YBDaVjPuQ25SpTV
JLWHO7XRt453D2V1+ehNTIjur797mVfS3RyOl1OwwQ/Rl9XvjKBHaj/SJLEE
WkUK41l3X6GWFm5wlnox0J34KVTF6ttHq5Nq1wjZrPd2vIxpxhBFHxomJgkP
4dbDIryN450pR0pVt8+QQ0Om54wNU4kWDI/ysw9rvl1oprMxUmOTnp8KEiN5
Z9o9hJPuwfECgstvMV+meYEdRO3ozrbrTV1O9mqzxkGM4+PSGzzJIjl1nll7
sIo464qGwGfMgcBkea3ZONWoWw6nA4uWVRqJ7ShTY/rACV8OfdI7cQ3s2L6N
5aS7varlysgfDBds4WymbiFkuQKM0BcffQS1mu1b2tWI1eeR+Hx3inqHFtHj
b7mqjLEf4P2EQwVGGnTA1ZBQ8QeX0Va6MUvM2gRbpKPF3h7RsSjziY8n5IfU
Nw6lcVC94F50a6q+fK0aNancEXSMVWvzjMjyc9BG71GSLT6TaNOyr8hVXvR7
7rVOOd3KSvQXOVuWyxC89ZDQAVXRBbd7ch2LmnQBhE0M53pNYZysQsrozkzN
xiA2Bq/G8CzGC2w8x++HJHVEUcHsVzULzqKcOjS/DayYZK14EoiA+zPDNIDP
v4iqdRYOU4S51QkRicTB/IOuU9xCCELddUjLQUnCO0qp6sujRvr2vTp7iIcw
VmjG3sQKhBiLZs/xMP6J6dBMxvklsAgFoAJvW/u14vztROU5OUpAbMhjIDgJ
3U2rzQcBJ17t4A24fhFGUiTXsF5EAwT+6qSm/gc2Qxd9916etgvCFvxTc41i
zBkBGK2fqn+autbG2dgzKeXSod/soxsVOVOEYvS440TB53jAlZ9Yb1HO/1j5
LarsnOWwuLXVcI4uDivHwQIUw4rTN+n8FLSEJ1x+gGdaBXfyTSxiznM1tDbz
/8Ht1HVMUMOxptoC2AW2z/q7g2wmOA9QHLjS+1B0fwRb3/2/tUfMnt4qEo35
4cTJTdvN9g0JXBI+92pgJYzSXu7czt1KCZmQSKMXY8BR4f3VeTXbNmOG0xc/
kfv1WUCZKOdEFtT6V7HujxyJzJKtNUfRpbONGcAC2+aS6ZRZvfY1iR40InRM
civAbEUX5PEjvHL6SP2xvT+uVVAx+haaTIizdakl0R1yCG+HEMLYcq02AUON
7k5JQunNNZVWQoP4seD+OiRzo/V3Xyjpm63e/3zf2s27jo3TCAUZPLrkeTD1
b2QdoHPms/peeAwS05Q/cNcPPuJSZcSgmKJNqytp1ijVt3zW+KD3Del6GjpH
3Q6DR5MvwG4zi8rj7EcIDCxa8S2Qatzc2ijnR06vAYJG6/iVbIxr6sObzgnu
PqarUBZnQuqKuwQ1lDtIHFoM4G9iiL9Uofm5QIoBX6qbwPZV4POwBMI/RUmT
GFDQmFZ30suL7wgwvXrmveCdpzK7UPvsyim6r7UNF2q5d0RqYMdd+m3636ty
cNqcnbfWO1fPEuvs7JCuKI47V/ZZDmyzg2uTBQCJSgRF6emb8ylrdwCnwlin
3PWwnhffSJAPXSqKLF8VzA7gQttY9zHboXujMZ4nK2FkEM34POofCNPIqr0O
Fxh/Zi9gqXYDDPDYMGvaPeqUfUSqgiRTFwjNS98lKrpwoclKDPY8DUU9Zzke
ulc9U+ifxXeoIeTBbOp3E49uWNwtiaTCAONT3Bwp5yCRe0uQxGcGlWBT4qT9
ZEsmQQRMupafyWY13lV9+YbRFZoYudDjXDx7qnpKDEMsOcPiCtLfBqor8YDZ
Q9CRjMF5QS7XJiO+91zOIS65lmekbQoCoXvuwoQvvm2KUxKPrYKkCdIQxVYq
ucAs8GmqOgFjnKJK4EDPkWu5EoKstBchRuSjjmBGBc0nXacvo/evnIusdlzg
rCXR0VnVO7bENEL6uHPbxPpo42OWeA7mVHzpwcQPe8qbjKXpCt9pnyVlJ5FI
woxe8n7rIKuj3nzNi9MlHYlLCzEdKlqo2p5TuW7b+iO/Ivx+I9S4mT4Uvdyz
WLDc1BvZdewZSQPuGCWsFte+xzAw1LCholVvPomIoROqci7UAHZvVg1PIXz4
CGgPr4A+OmbDEfCuDMaCD5p04hgQZsBEGEpRCU741TnphKZXuEn520bi8QKe
RKcj2+dTW+4MKYeQaKhJFficOBRafPjAVL7SZaMyue5znvV3FpJ4qXj0rxK/
e/2vt0VjX53PV56ekFbl8RpSxc7ALD/1Kh9UDp1RNxuveX+tloHYJhoY/em1
m5S2Mh66j8zi/VbrJ48xZ4Qe4Qr1ETKPtWfFmy2hidtTaXezEvd4Zo5QbZ3c
oXzFqqTXIclMP7289cOvtC1eMRtMJ6Gf9PymTr+ThHEr0bUNmt7+quemV67x
s1bE36YJjVtSg7vO+bxnp8pL1IMAW9qgLDUONoYog/F7bWrOJobCiNpuPx9v
toRCOTYOzi5Amcsydmlos0UrPmU5mz2IzSnNaaghCpVUKdqrQJ/zZlR9UtO0
vw6tCCBHeWDIxggaTCotkbsHz5XEKKxLf8Z0y0zNEUNwJN1kBNzec2sA5uC2
wz9CDYfmKFuxsBIIPMestJt239l4vccIX9RAKzreoUnczJwHlnrEgPiJTBtu
M7eUzWTfkurfEdiM5mTMWaaTNnzwDPDeRg2S4oddzC8Ysr4D7LwroV3oHyav
lvFx8CyN8ujNyHI+NriGU2CcjtTmTSHIfrZ16nrOClOgAWzxKJsLCltnRt4B
y5z23/r/hkZaZK+Ko4Nv5afchK2HK1bw3B4Batk2eVM3BCmUL2xdh9UxlFPY
aU3VbKIh2ah65VNqL9CHv7KdG1lQub7v4smfa14RRxRQevfa7PbmC6yGJO1F
FKlSCWpEUdkKwGIhOiEr1hMne6WwpQDOeP3asvtzo+ZIvAmjHB8vPJEvc0EJ
NUy13bgwoZZu0wQaXSTntv1Qema7O2spu6R9Wo4Ae5Oct0vpx76tL+nKXlHS
tHe10nBbioJTrholCf3SFygLsfsgkTcJXMnr+K/2pAa1qctOk+4f6owUjbD0
Hrvrn9wdMQK7ETodisUj8qiTMDqEYb3lvq+swTsildTZQnv4xyc6CxKakysV
9+QGe3WQzjEJTdW1amh8+BAK8So2GgeSu6zKsAVgWS92YhHXTiDOPBA6UYXG
OyCsqKkhelJrKpJtP3snVdjf17Kgy/hK2LE0I2c9P8YkBKe8WM2yOJS1r9Td
83e5/NNB7dbOE6pxo/Bw+V8e6fQkUj0xZan2tjqo2r/pqrQHgH6YaOb2n9GA
ii1uyiJRkkiLDa7b9FC4HzLgXvaQrYEDCwOFGIllV6whyxQDG0sZRV4ztF3W
Wq9wPH6PMlEufgJMT9pStNNNR5be/YGa++AjJatRuSsKLDJxoleetYTXz6+w
eovlPbRveD3WQKy+0MjyVx/iobqQzgmIBZaOpA9XTFY2GMjQnm7NARYxPaz4
IDWMqzxNpFZfPgleVssuTMTQkBtZIYmuyTUPirbtiR+KUZhf2QUa4LmCAPOd
IEmXkNNfDKOAjGLBIf+B/s27QD9Y5ZgsaGbj8eaIx/0fTfgCOwn5kJGVPf5x
b3lpGC+S09oUtiHi5jaAnDUM2E/yd7PS992jt6T/Md1px1LBgjmpFfXeN8F3
7AhnMSVC4a7Oj+DngblgTrTWhQ1gRQs5aCYaVQQ+t109Pt7F/PPU7sYVThfo
GTai+qEXEGRskuljvAVmt5MUHG0c6QMTsUTcmO+odqNURpmtkGKby0sowFlJ
zy0X5mODpE8KG2u+y1q5Qs/NdeVu19hNYQubT3ztZR8i5x3hrSWjGgHGP4MY
0ajjVd+4Kbf+CwbEH0cnXyyn5wZZtIlF4LxOGuOANYGEgNxbOV/PMhSA1Pye
+CXcHCsB6sKO+34EYqbvlMChH5FNFT202LSUEM4gBCAIdz3Iq96ztC6MJFoP
O7OsStBjWF+oCXeCPPxMvsjvNv11crXEPz4oYHFG4bFCO2rnEbEwdaUXDvNt
7ng5assgeEMHCrl/0xMd8+JyGYxLll0KAwX0X510zyxfONj8m6+pvY1sGfnk
gCTysiHu+2PTC/Uaw0IxQH5D61lBhG3Kz0Z8qpWFNn87q+yf5QYQOFdxJGsU
/jpovnFXCN4AmESN91iOd/o+dzeGhu/gDpPNJjkn+OvQ9lEmwmmR5dWFV3uB
3bEU2SKmNA6fbRAuqO259P3QEuQ+v4oLIx1rf/sY6R6/v/zbqUk15Z1dEQpY
etbKp5Vagc8LYEgT0NFBqGcJmCmC8buKTZStC+pu7RqIHxWqMm8gxH9hLPoH
1JzME+I11e07jf1yDnOiA7JjcHWsCGpFGpGHi4O1R2IqlvKu5egGQMaQglJ3
j21dGlOtDMvPMeotWm01qmG8JeH9swUstPledgbFeDb9rFY5wKbin+oD0k2j
CulaPoT98NO+t80V4nsckopZ/l251lpV29eFXAUPOG04X4fMFPedKgbrDk/W
nKPXIyISkM7R8On0ezH+nZmC57WXaz+zaLDlIINe7nneC0618G0396qtvQhn
y+DHb5MpmvpKossaHtnylvHURta8eXArIVUjwM/3cY3zW84CkYrIGxHxk/tF
wcVee8cLyBkgzDGz1xI4iuOGCHQsAcj0sDSiG0XNISaQVAmrR0eWe2iKJ03v
Kz9PgQeV2bGqkile0Csfuynrx4ivZWqs7Tf3FqJIHMHOxntqBibRKjThZ12N
ip/t1tEVrkHJxH3Q7sSTsI4qPKW+T5lDXvR9IQHWQClyhAFm66BaaMC+/kcx
6cBsmczeyqDvNSWy/XG4sbAZ0mG/4GbBru2DARNqM0Pcm8EubzWCYNhjOINA
DqvAU4ALpYTCna0l5sp+goKxQgR+hR1eDiWRHXO2JOEoPUPdX8tk55siB+kt
C64nzbAQOcHF9dwwkggcchJAPIz/Vyti29I9svI5DaiHNK1Ds08gipqujzzT
OR4+oFQ5r8fvk47ilcebRfim6Ud5LxZEbgfR5uBRt03AtqgjXyZi6kfod4K5
ziG9x9vaQUnCwNNhwPvbYUbzJBhWK5UT2q90fyKgC4FVSOlTgAlBiQ6pUR4E
Ig+3Cit5whrTdwPo0uAmgt8CZcP9SKNnJy3FviqF6y3NMkjQkyxP/chbTAEI
xAUqKLM5WscvONUIXoOga/QE+74/iKYBTc8bVuIWS/YbGtCJi7t6GJCXu9pR
6fVwM7dxMDf4XLTx3wzGLsn8fcRnqgM1WzfzXN+Y1K1EoUb70hkrg6H5fXWn
zd28NfM4sazKe+ADRFU+2oNPdaIRM0WjVYcwsAvY0EM+BDVRSnpDbyUyzBcB
n+hTBsjNGP3YEfbqoNGtbG+m7sZY910k2FeVvJft2Bw4/3BcJbdrX3cKK6WF
1krqLCR/ma1OsLS7wrOVWziOamZJKz8XwZhnjCmFjA0Ou7gINgFIDIRVPMHU
DkiCHOLYD8bEfsGIXfQkeWWnVVTptVbEL9KykdxNGE1FD8AayjAyfQU4HZM0
iZwF+cbXkZOuub9X7rHafuGmY3+R/0hMt+snlAT1bCt2rVe15PTMpLGMgRey
y7oS1V2c7mRg7ZDkT/cyldFHbeuE8RnAYk1WwioyF9uw9eMBqbpeIBdDFmmK
FCW7TZM0a2BqrMOvmLcv+lrreYdgrWsHcvCR8d1x19idlojDo6ue0Hz9C0I4
mfhQeeOIFVkYITG/mDl/aUMhQ5NT/EpMTm3V5B7DI5U8ERhQEZSIIxkbWHKk
XuUKCc1q7mufA1UqalSHHFR7nOBpvOs4I/NOX8QBBde7wCGrcMiMzbTwvoSY
aBotcQ0ba3Wtf2vXYbDNeklJY8r7xqxxdCmS7ojTCV1CdsaBUpm/c6J9vKJx
3fcs4uBqJpPjdim+Zo6PtwWEg0zFr+Sz6erx4KzSC8zUFNtoSo7Q1iLa5i50
EGwVnxYzqh6JXO24rEIjmUcZXc7J+PA5T53bSxfczIIl6H7rVzYpgGQCZ5uo
wq9kw3+NkgdaT/2TEHlivk8DIJcUwXDiE9cLELuktCXsLuJti+50KCpaKcZJ
ZkfYKTJvFirofA6/uuP3edfO1SleEMgM0y2yV0P0zs5R7xdoARm70M4mptLD
t3IERY5DrCKvAZP7bfc8lfN6mz0bfIrPyhSB9tprfARAEIOzQweVK3UYxOam
a74xMFMeXyEXLyjLS690AKYgfMAs2W2FutXxmVQyytP3+eAGsq2F2DtlV2yf
JCljFT4vXG+Oi4+PBGg7Xt2Kc9jWIa1Cl+ODORcBsIT0+e+F0Yex1zsRjX0H
ezLxk18aKp5R5j9RXTp62qduPU3QlcSHyqzspFjBsHs6LmHlrvkNBCmnaGfF
tx9u5lWUn8RqQ+xsfpbnJdsL5t4fGmLiVS5uohi5cMmUcy7up95AHyB4v+dV
DhBdy2fWqIAuM2H9/qyQZncXrdiH5xhluT5HdAw+6uJtFHJKc+zIqUmtHqbo
ok5s9v3lbAyNdyTkJxhsImIvLSKQai6lHbch0oGGugBPUrrUSZjvO7UAzUj/
sMgL2mvAymU8VyIhQEXsYnUj3MonM51o9b4/Of507cJm52Ut2LUylxycfVHN
35g+BzNzRnuII+i9Fn7lCk2BINPkNUIep5iV8pPRBlrxPe9M1YLrtk7B8dGJ
DcgyUVdg2g+l7NfEqAc45ICK21vzVxZCJFN0uQWp6XaFHwbBgtuHhwz93bYf
tu7GET1uIZNGJfuDHeL3X4qe5zdxnfbwjviYh1JIafKOcQ0oUr/AA9Br3X0o
M0XfpOUqoNhG6hI+/tK9n56kf9xstt9Qk51X7YBUvDZm5SUgxznE2C+C5M2h
zVuyRBG5UIbxRrIDrdh79JB9kAiVmjeUgOro2pjo0SSOlnTj126m9kYeJsA6
go8mIJf9CDlCJX+6mZcgQta5zIRzpyZ46wsHAzM9RZEPyiP+v5PpyKQVVaYB
MfTbSiBf6o6SBUfyVIDQA2kPHR98YLCjF/wYhMnIYXjPveCgDxnuY3hLa3Ao
zzlQSbnQG3DPC4JQAZBQcd7a1yswpOtnkVLNzrpdBHfgDZzN/rUQxjpnm1n/
ShDk0K25Nr+Auwdj3cmaKksYVbuFzq1Nt27re051dI0iSGR3r2feXOH9Oxej
UlKNBnq6cvhlZKdQt/lTkig+eV72UmqLMsX6COPb0dCnAPkaI81dKvxr3+jR
9yWc5BWLyHm/aC9A1tpawHqxg7ny/IJw2em3zOLI9UbSJzO7BF2NvaNAG5Uu
T7QgvJzXtrT/pXV6J+ylf6FyL5mGJ6xqjQRbxLbjtDFfSfY3NIdXYIG67eUE
jZinnWKEv6/2pVzIOPRpvwu9M1zqLBGiB5h/ATm1dvvOlM/90BN5p0wlrSpU
lTQ9uknWoV2kQdVPnZ1qNi3c1XTXYGAdBtrZJvLMZz4LjvDju6IN8CwkXrEs
AfxXXjMzPl3OXnIlWlWaOFDXKnrRwkzRuYAr/S5u7OHr83cgYmc8A43q6tFS
YZP5JmCpIRFAFMxH1dmb/uW25ree2XgrsVdGi84y/X2QFEGZWcTskmEKH7Fg
fTyDjTdNS5xGInzQhdEqv+QE6TmaM75dmmq16CTaEqRVXrVBDydXtzdqY6Q8
2VHcDz7gtpJ3dGqjOzQFCnAxNuevWx/M3KtatNlBjnDENbKt1vlSJuKGHvKl
yoLzpHwfgOIRNwW2S7lR7RsZL/jVDouYst0zsytkWLvDsV+SqLM5grYc9bNh
/lixLIJdk3trO04a5wWxAIbTXC3VXDW33kRLW3IJmqiIk1Ki9ImGuu/Dijn7
CqXAIABUQzoFyyukkHoExrbEkO/JqD7gn/xwXQCNm1RRfOLMmVD2QWfBL63K
04n8+kURrreXCb4NbzQ+iAEyJX7e2aYT+1WqPuuB36XMr+eTSi756mXsSBwh
brHc2UouYqc63ntZbZgd3OFtsbKhthi2bs5HUCxRYw3gwQjn/P8F786k9O4C
YHPXGvE4hCn5TkzguBIkucYhnZMDx3d+Cb4I8nYmZl1Bg6airO6nfnwNCiq5
8w8XAe6jrHxIQif5cfdTkFL4teRQsh6o0NUXUdiY4GV+XY+DJ7URGMEZoOAD
11Rc+mnaMLQ5stfVfUl4cJtlEaF6aF1Nuss2o1wArSrP4NdFe/t7Nj6Oonpr
TOP4/l2P+KXEJM0pnSdQKORKcmpmRLB74h7Y09Psd649e38O/+Jquqo4SE64
DpPUNchI2CdPsx8WVoAlI8m4Pmy//0dIYDebs6/7pswmKoBYz9fDpUed48Aw
8SAbRxKxxKf5xZ/wylRUzuto9QoE/8xcJM64Y6Mh0RJ5DA9E2k19RqL09K1s
/X/KJSYTwussSYlzJozHcKrD5aH8RL3Xi6i4+LbZIui9+NyWx/ykpqFeW/n0
yOEBJoUlUQ6DGOUkzwmrOR6t5AMQg6jAjlD8JCLsbDdshd3ISHoh7+mw1kgV
rIYTUYPb8Az/TioDru33fAZPR3F0w9kPAmcAMGSNQm/83iq7JnKHfySyEDKo
UhQeAhZnNNTkUFdplzCf36FaBnrxvDRG7X00XpbgdjYWtdrNd4leSpsKrrjS
iuJjnTFT9M/Y065cLP0RJWei1ICSEvLzE296MsDjpuOPNFLB7KWM2DcRNh2Y
ZG1z2lq2OMwNrWd9qyKcpGKnp3DbGx6LucL/HE9aBODdWATd8+N0/niFHTA9
Bc3gRVwkSw7bGjt8Fg70aEg8V/IY8LQBKXFmPf/oOwxUhKvV5YeO41lTG85A
en5xXEliZR9LcrZC0DSWltIM+iSuv6bP7r/MgPjk9HFRZnu37WySqIntSY1G
Cz+qo1MLMpfEtqU6WUeBrFB2YKEGbt2U2WjLprLwUWFeY5NRg5YUBNA1/Gjw
6A3/lRM7nMwT8f+MybI3yz0zm980yqNfV82BBul47y12nf8tzHDNENftDkBb
wH4CM904ISmyj6tgzB+10rVWxNv9K91jAfoaewAq/vbbMXNniVCHZDqGGW+7
KgO7F3uSwdk+2zsUHthFbet+KXlLoL7LF27uTB1kA3aZHhCM49NY5UL8QEDQ
W0slyWFBrinoQ9uE9drg2IvYkhWjB3UmrJsEQEugNqjeEQ/akiM8/XH08THp
oEsRAHjbxwL46L1BwA73JbPI05LoZW8uERXA2giLrM25l+b3DT+dZHaw107v
4cAf+f0fuT8PHsoOrxPH0IktP1gTu8fW7gfpIaF+9wF0LZNf4AG+0s55WvFg
yo2bst/FF5XRTWiT5WVhz0+MKj1SeqL9a53A8rMqNgkDq2LN7poYONyh681k
6Wrwnbl2inwxSl9Th3ZdXUgIy220gIDlZoiZbEiLgR6mJp5PDNf3wZE95uFw
z1XnXuAEc8CDBc4842sFO5c0iln5VVnz3yDE/axHUmq0kBDMgUFAKOOkzjm1
nRIqv0yA/8MPp4xMZ/Lq92az1INtUbOIuhtKpx8YuRXR462rAytsprOqe7R4
rf6eUI/zVWQlWuowbTtmXVg9C80szeB3z2oZQNzekcEBfhKzTCH8SCyXMiQe
c0DjVgNWVG6ezkwLxeakpEKk3AOwE1A7/0yhK9gq/DecdSSOnCFIkhN149qX
i21J0v+fQp9Hc28DKM/bxCZ9Izylp3wtI2UY4KvP7uTnQ7ZzDOMTe5KZvjHf
LIserTOvglZePO84XYLh2cQKcVCR0TUZZDNnB+gJZRz8eiUjgmgy43qLoSWY
VAZ/ciIO+WloYY6A1CUKoWuQBnR8cMMKmNvmZ0OSYNKJDCJQ4xHxsIDtgWhP
bvvvKb7ob6jr7cbmjHwT9vra62o1E1nCZVBOyK9YH1ha/Hg7eTR4ZTlkjX1j
WHKxlhhCTH97chAsKwkcDAJm0xKM2FpgEm6hv1M22hEHAcf3OyPlNHIgQB5q
rOMFD4DRXRPzU/obZSaRSVJ7jh5cuiaGj0B/64YaSpp/cZfz2OagSuvrBbl9
q9oDA0bXGY618ckMkZMQ4BXXCh+CiPb1o+9sXQaYxiSjVr0b7LSRgjkvLeFz
gfcSADEBl1IXhb8RknvlwA+vG0ak2vZl5SxO63AOpmsXNpENyJ0AGaqw1hyT
gwkEvHtONtfMj+o2t4m9OHFij8s0j81gB8mBufpIhRy5DpeG61V4JpoI6L+l
NnzmErWceQu79+QuXsjpwqi5jySK0aByWL9kdbWtgZACL59lRua5fCPN+O1E
imiP265gELQ8fgZdsgegr/RvbpmmmNNjpqtJCRHdup9ZO5LeQ/nPrPUz5mC5
oE5IYmFDI+eQw6cCVcdo+2fjJH60PnSC/nwqIQYfnkSdaWDf6R3Y3Q8AIgyi
PU4ZTHJhEl5rr4aSvC50Gs8zLRwLdNJi9X8dmmZeTl/EVzeAOLolWY0QIODa
R8LpBKd83y7791HjdiJcI2MLOi20/p6PAS/5xkHyCIQseBZIcHknt5lFtp5Y
rqtWK9PEG4YnCJeWEhjkky3jEqZgi0iYF32OXCtKThvt5MiGvwd9aiySQ4Jd
cXeLve3HzZW4yfbD03ATFH5P0ZjtXmj49aF4MCuk9VpI3NlCGqUCcjxIvvcy
EL5jWz3GZIhL4AXW0tx5m8nwHwnVCXlSov42hyCalnoCc0wb0maDitM+8Jp6
UHzK+vpwSwgwiqvy+0kWPCxN7/NAcf6+4IsC+0Wr9Z+ffw97prFyXfdrY00P
MvG/3loafFeCbtK7ncNkhvwoAqxnANWJGMf+AoH6hBXcppylujeIYMYMdGTM
MBlxlfkPwz3i0pr12VtG38jZDPz/PEqskv0sIsTK+itmkjO91aQZgwkkV9+a
KNBzoVbVms7KNVoh4o+uI5cLoCa+OLyGoXJ1pNCWH2RHFUPTHoVCNG1tCVPA
VCcLQ1t+TJ4QGM4ufwvdnSiZMpImsGjiSQUv4FRbpUccyl3RWv+FFFqynKnS
Vx0R46xhE3RnrmAKz0ijPjU0CAEpb1U6yEIT46vFKy6xvbW1use8PX4zDwE1
tGb5T6apN/SkHhSkDSYE4NJQipqOnOkAQC3YNQTUN++0Q+6VsqOkn2HQT3o0
Ucol0TgnsSlk2mUOp+37VcSnLLb5JdKKy7fERJX2eOPWHNvIjUWQAwbbvBm/
kN1ffxT9dz9nW15dhPy+hIVXXDq0TEI+/Xd6SRbFNn03cQ5VRmwuMEpTrlmw
tH4u//sOmWsLJpPyvTTCV+AGi5Oi8u5BiSWND1baxu7fRtPFIlJx7UAVKmDQ
CDHiQwsxNWBDaZeBYgj6HtVQ8m3S1kcy7B8E6uiDGzlS0Jumj9oo5+dKSTX3
sau3aweIpxEWjhehq5A92d9DEQ4mts7oqfZsWNVsOKkjJBFoW7ir6tkm6o7J
W7Du0W7mvMeVk1ATtTW1pa8EZWgfARvtaSgA5VO4xU/AlSaZIFFf986C8ICo
i30ZV+FeXRHP9Im3bi16KTyGTHoPurDZcdMxtJ3mHnPJWjOfG4I0Z73sOGLL
VNHT3nLb6Jtlk/bSa2M5KjuPI5uADNRuXvubpmB8znltQedxgevV6SxwdHoy
Cl6Ry9sZQgpeeCTRfPXRwww+3ZePQoVe8GStd+P6T1XidzFceMnIHeMl+ob/
1LYdwYnnaD0JycmgTVtcPz7ku4G4yrW/m7gW/WriNZYWUXBCIrWSqbqOZJbs
Ey2tLTrvpMvDYcjA/kRuiQ0IWEs7yD817dJ45DCYZkCWv7Z2bXniMW7GxZiT
KayP0ZZ0Nr+5bf/d1jZ5hF6LbWD34ziOmThNeeA2nv+RH59gkNpIeazJJs2z
zuqorgD9q/sNoO2lPC6ohFFwH382uJ2KIsbskxM+T/y2Cyx1eBNBdV35CU1M
Evr6e+c4LYOhso/k3MMvGKALofztRK1Q2LxF0Kfqfwt1wEQrQ04W2fN4oHZJ
yEaiI68mV6b5YB9USpRL0SsMJKk5KCh0YKEzdUH9aQMTQuEhN/bP949HafR+
o+SUg40ZzrlnfcaiUlHtMr/BqzyvPt2atVf1qoPR1l0a283T6ajSpAEi9tRT
DRXXQeDx1zw0fnR9tCbS6qg+ONMO8hvt7+BRs50saolWcppnyPTn2yK7luod
HKdGnoGZKP1t6VeJX8Chm4EEK74e18vYvU+Yqh93x9ypMwXuzwHdOdRb3PLU
+FXhz7GrdB7I7uAJARC5DC6jbuVVmFfZijyk3GDu5dIAypagjCN5knfqAbZn
kOUeloOVjXZ8N/Fhd/YvT7K3SNWQArnZY0Br3iCkvaeMk62FGP3Kt+BCFWlI
J8V19s3vUtFfk/F5/jIItOBxs3DABZXpeWBUamnKOtk3xb6OcvlP+SN1u1J+
H8sQM6OddEmtD4syYv9xbOJv1iTNAL6NMKWWYK2fq9PbFLPMYA1Cu7HVvaic
VmnVj6XK8CJbuStg9Lq3eiufCWIUBCcbnTbUogWxP+jJ/MVn2N2qdza/1a2N
ahGXdeCeOiMqbwaPCT/b0P6E3UAR2sF+WGg3PUItoHK2nVKtKNbAFW/SsE6v
U3FbUZtc5v+mxHGIxCxqFsJCYKWxMzNX+itEJ58VOS3+7g+7FwSCsb59vKtQ
H+37TSiE/CX6B2Zd1U7ZnUaIePDTK9gYI27S97jUBo8UqjACzp6xl5ZlGywN
S6XgKmvDGCRBg5ss1SByA8RCqvEmAUhAizZrT6cYq3wbk2VxM4lSGLKVIWny
1Sxc9PHCSnImudeNnNHovZNXdBsXmvFBrPoYxoXcIvap0z567cFl/dXHFLoJ
oquEqJKFQL4R3hBuJIkD096Y9zBdPOvhwdZqMSoPUe2Z+MFCz/gsJPJ92DYx
4vRakt1q/KVryuy3BItpclI2J1sBTCZInGDT+cnEv1ezUDyT7/yVIbgFJclw
pLhi7N1OkCtv2j+E19ES1xSJT29dvM6By15c5ZnVFmFag4jGeCDtfr4qPKQ2
RxxKeOIa76tJYscSS8K1BgUMDYio0suge5Mr1mN7qF4rl54m8JSaOwB/27bL
RtCa7b8xwe07bmhmCeS0cQEWrhIFL5NeF5R1b3s8YaVv0Ds3Z7D1Ayk1itk5
0aNROsjBOzw/EnpEVqj2lkABI4QYq5F9owj8nmbxg1OF4soOFLIV7L5uBNCc
s05Z1lVZ0a7ftudQWVzmj6530iCzG8tqX2eixrXmrQQwiB0S2lSfzIoJJr7e
i1ZUacy+nvsH3Elp3OWm8WvjNxLufy3pIuXmXQyqWQkaGx/ZOXaRWxFpVsj+
4lMY8Y3V2BqynoD6vMHeCRqzj9WmHX5LtFILtjO/qHV/xRTvxy++stuaYrLv
lnscjhtvnReEimLSvk7OuaEZyphJddROKD2jTDb00JvJ4qVDT8OTP3lgopyy
5Oy9bhoHzlHzA/Lp++UOY5qrD58Sp8DB3A5FVEdPYhdP6LsB1dC1WhSnh84m
X6ZsLLr/AI4egL6UKm97tfLsYXTwJO93E1iEYLBZLZMGapSREtJ4fJh992T6
EhBg7Ayop58SexuVB4+/9GhGIpjB3x4TaaCEjlGZnE9pxPrXTyJZ2rT0Gmgb
GQfIvenDAByb2tHT9psCnPnGNJnstqeg+5h5j8Mef9J12Now9d5t/ZPzVmRf
AF5rt4bqYLwig5PsKXfln6yULg9zFRKnWYGmOsQc2MUcHp8W3gq3B+ZaeiqO
aJ2Sss5QZ5ar6N9Rjf8NDoRPcjCA+zukHDN/iZCQ3PGAgQaKKZcPIv773ta5
jbMOsyqStjRxdWggsqIFY2TwrmCQ6AMBzgrdVtRQkOCcvD6YfQ4Scc6zN6RZ
ciYnjJT5x5uGOI3yD7p2gyHuRJqy+UwHgPYBT1zVxSPFShdP2Z2FeqVpPQzG
aB/b8GtS9Ld6TX5ooWNLc75+tUFKk1r4oaRq/P2KdxY4G5y1taC8kHPanwCX
0/rsceDnGgZfbCPex/TMqC8Hc/hnPTgHg/anVYhJwzIkcv+G7XHPWjEjw9bp
bKRBPpeyIro5Mx62lus9pxhMcCxOIuVFOmrMKlX6kAUU9CnvZfdUliKbYK3l
cVaamEB1+7n1OvXTh3C5ZMXngEl5BPOZTrDp2wxQjy3IsSK0fwD8lfM+MFwd
cxO9isTWD25LF9KonmRWjDt3yAcSoXj5DA/SIQIomxRcC7CIsah4N5z3sYuw
/fKpWgwn8LBFufbh9x6Ae6tvt9XJHkcuA863xvNokGDK6/kciQ63dnOhXtGS
hXJ0dsHdM7pPd941CroXXuKamLRraIvjbrcvKDca0GiJBKmLdT1woeZllZPF
7Hz1u5V9kXuA/tqj0/VagcpCkEEFMFPlIpq7Fk7Dt/M0W6FFUohEKDLGOE6z
1FAb24NkYKje/7o9KZpKwBOgPhnMa/rsE7hCO5wZj+lcNgkpTdipCAgS8mRB
wDB2Hr2xYtVp9O52HQ+ZydOhoed80/Gy2g1XucYw5kUWr7QYoKMUZiCWBOEo
PhMixtY2yqD6OtWKXup4nZ/WEbIb+WwoEsm/V4lhjRZIkUzkn2noeOiMO2ee
XE2nx/lQnUmbdiTuU/OAGhjqUpdHlU5akfO7b2RXpR8RrCN5O6es307Fk0wu
e4TMSHYDcK0Mp7jboJbu1DlH4ai3TtXSqa2wHBAqEBpBVFcIXTK9j3E6rMZB
9jdnLPkxOs9xPjKKpfLPPUMArZu56HCnW/miEGWhplF2q4facQgs3Zr2t+ai
TwfmBera1XFUH85qE1wRNsKfss5LGHCbjnzyKgMNTfI0Pv8gvatQlgV54yje
ECDMTmhnJFoVz+JpZr/ecJTYCfdaCtRxwURuJGnTRh6YOm6RWeaDk+bAs0f2
qF0fD6OY+UZyA8aEXxZizsBMoAaqYKgOqDPRSTcA7XRVGGeFsv2XKAf6j1ZX
XTa0hk4ux6H6DrRKgsOtXYVegP4wYM0eiJG0twZDOHHwO7j91DaEM1mMlKLX
BKUVQ0p1ddtx6BbfLKW3xifkH/XCfAhL/xdIOn7ejUIc1MyEyObqBETw/A1d
9198VZuHPP1nbhMSjrdYoVQn+j20yC71FW2XI7ymfSSrvMeL2HhysOmCCEzX
3SgS16UzYL8C44O9uBddbUZlcHoBM/KeozFEax2+JZm29vzPr0DuOy+XbCgE
Ol/3Kr90c9SZ4XdJqNyKv57PRxA/3gQ84MUWAq6P/glafq5NSFt5eCJF4Rdn
5UMXeRbPGwN0ILieYaLXwN8BIHgIDnCUYGArm4tgfDE92OPpgGBfq6FhGISJ
Ffq8ibtwA+VvHQ8Tk1jp95grn6Eafvknd0IkJlKURHIvLuewDvtmTlg1g6pS
0rxX6X5LsahLVcrzl+RF2wt/m+ltDCQSg4f8bsjTr7DnyWITAV0z7R0uoH6j
+JTh6Go1yj/lYSZ/BBPqjGZrK9iLaV/ECy4KFrTH6PSDwlgG8RzEmxpIAwfs
gPV9K1JFm1IO92LTWU5mEEwSKizg58ehW9MZECi3dwqJfKuOkmrLsdnuxvUK
xFyJNZynCb73gSib8e9wGWCr2ar6n9TUlHgwLTAcAFcHEi3lzxJ6EIxFH344
THMeWmRYRGpvFJ7gfyuLwPCn6YLKPCcEgRWL4YURdusdUBsNX4M9FUIbApw+
wDyELKssvf0rkBCrrV7JH4X+VZ9j36SdnRAOvOSVuwAA+WEaAiHn4fVD8RsH
kftYSM+Oc5LPnQhkk7dxvEd4pkq1N7Hv7WXATON12vn9WaS8yBJLIcYF/VEg
7tUETupQmTtUfm8GC6iVfwfgz6solcav5vya85bgOcVTHuD78nJE+bleZ0uS
ooPFe/C6+DFf5k7vEgxjtB1qkeXtMLX6z2zaO41HJ/dq/xtAi3sMR6oung4U
QrBnGXelSkGz/Cb6J5slNHU8GWQWH7g5LSJWbtVRmf0YSla73xrmDtxVBQ4N
LtXxbl2PX25Z2qy01Etl8PtAyqREpXCtEGO7cg8/4F4QOmvHs5plcHG+Gbuy
OcIh6bj/aB67Ml2GQTQsaSQIpzME1r003JUT+5s51eM8iHyKNlv/li6RLeYp
Q8USfKuPHIv7l4K+kLWbpvKrpZ7Qetm0EuqdR9EculRaqiqSYuOev0ZjJ1+k
dWich23zat8kZdAxoZN6eRoqti/BcE5wQcHtVb7FdYv49UqfOQCjfj6iU2CO
8DZp6rDX9kKtm3pHziB1OLMO5/rsvlksnWNS/Iy1hZG8YwVu9ri6+n6JepVn
x9/uFjp3SYuTH9pPRw3fBa3v+kTFhZen1JsUSnt8oZ4dsKdDkJ0OGYk12z7G
2Z3YUtzyFsEeRMVy/rAWF5pGKOmhkAQiQRkB236h90HIEkvaBUbramDrGE0B
nvN7e2Dxmn6si2k7H0bX+cqT76+Y4VeZ/PQUjbds4aEH2tJOGLPTTURI93IE
wjA93wB3MqEVGofHFcXRiocqiybjpZ3ydCnJzKudv92yVR+CPycUVw3/2+gp
EoLxgnZks8NVtgkh/rp+q3vxXxbvO+4zbWLmwgFwCH6FNQGFi4i/gL4/SB/o
LuvpScnb6ZtZ1SMepIooLKx8t+tfI/hv4MdorCbyL3DJCu1irn12qDDs7CTY
He5VxnRCOHWwwQN+gjHsERcuKdblPMxsLoFIinuNDsM6O9mCLJ5ntHkvCGz7
uOT8Ae+MS9Gf9SUu3EUhi6ii7I7/MXaKwdi1xpCe9me4ANThzUtySn6gyGvj
ktt+cNSuKnhbDmpN8wd6oh5VqP3khv16XDkwXgDjlZQ40p8g/uE1n3+gHJ6n
mAECl3cP7137O7b/Wr/d1rqaX3/Ji6TyeTTRtiUCh02giboCWd7TYpZ9JQNJ
0UKfm172MrLBimNXwQyIkduhhGKhRkY37oxfXOfxHqIQkL+MjLO9dF9dhe9n
WgX6mFe38Xp8Uz3c5joqtI0Djm30NknfYA/tsI3S2BFZxqQsAes+J4R5v9nK
Bjm6PJgL7Lz87LDmF8HOa7QoVt201l/WYEzFFYZKqcAuxikAAvsHRC1n7pjI
GNoqIRGdvXH6XNf1URFsXziKiYmj/+7PAF8SaAtm9DzE49J/UvhgsbOWBWEZ
9p2rl3XSLI7pWmt7AGPLAONRAxODIFXIf95vXeUDa4pQn+GYc4xdDgBL0fXu
A0pVtK5AwwUx1ICgEUvH2tVk2BqLqUzdZmBCCalRl8ng7HphicPkgUByQsrq
ggxhMVzIJR9eBYTWGK6nvPdJCChIWIquSxwpvzkDRlfAua8e1gRIpcqWO+c+
UanTern8an/sr5XwJsLcNkkQSEH6eZR/rNedyXK3rTMhn/zi/UPsZWk4YMlM
YTkTMCbN9cKDeqzpojg/CuVqDkfQfLl+OU0elbmx+kr0P/G2fTLW1NBKDSgu
tVij9e6eeufm3maSp8gRLr/wWDxsnPeyg+FVQhbUq4HZ75XXOwRkZfDGoKrc
7yTGm+tVSA3XbuinTpvgadHWAvom+EtVXr0IxTx1M9PgqLcAmqX8WlsaOnbU
LWHJCyyBlACPuZdLpS4ZhLJ8R4ezQ6axuHc2E8/hmZL7VoqVEKILMZXYRD34
ek5cSM/T/uS9JINmjAj5los1ws16A0fSFZP60kYy7KX9nmN9HyyUeeRSo6UX
JUM5deD54vRgBj/XBXNC3GP1hOhVuZAlWPlROG40q+bOFCXSK68w880Ae3nH
RgqriRPjUW7o8KqewBmLrvabvUpvUiJQRMW8ye4S2CACWg63ts5LlwTVZZHT
wBUyLT3uwDNex4IxAtJd+oaM5SpK5HOBSqFOXd89o4M8NheiVsPGW4a2B1hQ
s2n+F/lt6991XbIQLMZlcfBj0KShulfltemeKR6vRpFSUs/YHZPuz24+xdnN
hN8WwUg33JW5oRz5ZlOi+V647JX13D9khlQ/JhM5ZVpZbSZlres5XS5f122B
IgZpEceVgKqC1uQSO+FC4pbqiz9nwsRFcaPognoAB4dMs1cWWaqKK+ibwPuO
/IVVVlyiXsNOkppkKjUtQkuquiD9o52+Tl0xk2CyiEhQ5pmHernQ5n/w65F1
bM4DquyvYqhBTWK1cZ2VD7cGr+qnP6YDaMFI/evhQmSUgJtsgqVQqPsV8SpP
W1Y0mg/neRkyNFzBJ+se1o9OqAWACTin0UQK4okPgTmSFkO6Iewr4mCBcS8p
gPkKleE1TWSSmE2qQd5nQ0VjnePAZ50owNcLX+E1RRvJb8y+O9duNqGt+fdV
I6r4JPSofFkZr6hojbQmgpSwK9XfWqwfXFfkYiJmUyH/jowjtLxH/0NMn16Q
/yRURKeLD6uzDYQJzrXPhfrxFjFWt6ssbmpops/ZiL6LYikryW/nDmO1Gkc6
APTQoq+w86tHl0SOZNAmhD5dAEIUzAm0lu/DIkDHQj3nZ7xn2CGVmAd7fdUw
IdrdMELZxpqza2jvfiq8+CeAr8LeB8HPAADMtpYQ8Yhf7rDpExOQbOZ+kmI7
oTsfbthUes3aQ274D0h/DS+AwWVpE+Jijttx2pF8hkTZ/Fgl/8lU/QuJvfW+
c4EQR2I+b+kZ2/4qbVPf1ySw4PIGFZGRd3SNhk+gtkBX+Chx3GaCR/hY20hL
r/YRPTJfIxPZbh6QFDaYjE93Ve0bvNdWS4Ae0gzyEMU9MsHtHxdzhsKbUMfg
PHCAP3UYDVdOAFJdXARyS7E0f3cX4yQno/HLxm84G6oiTKDYEfajPfdZSo3T
KO7OGdBWZZMNedZvY8z6kYceOSj2o54gniXkCgzbPLHLOZA5RXe5OYRZcD+x
jdXC5gE34OCuqfApsuZxCtN7f7wjxFcqZ4NMdEiBXLSTA7NMZKgiwc4/PYFU
BiT/f+ygRnyW6RWmpqBTz5BLayn2DdrRVV7SyH/GORA3tU9nzathV6cgjKAa
1udLDTZT7ijNfuwdFszpsQnueaHyYVNszym0g0Z624aSZdRsthosqcr0x1Gi
IYSZCBC18P6tGbkQ5MI9aYxhtD5ngfhEKlmvI9GoqxsoMj0Nr1JzW2rmNDoT
PEmRY6dlwHdTxNpgzQNgHgwvk0mKrfznkhhj1ireKnoo1HWQHnkKdIPwqJQf
4RAYC+BjoNXsTtwtlaCDEirzr4ezPUA0uTv+Q7K/z61RD1yitYuw1ONc+IDS
tF85+i3LnzJcMJEe0SyoUIU7WbBxjGQoruAWODYo20blJNm1JARAYTdQzazH
fYO8RHL4JWilkQYeAbz3B4FBJDEnDKMwpFL4qsNeLiUNRBmU1xJZbZbQgaxb
WDjV1+a91gevr+F+b02UaGhClgUWhN+TFyzQEwOiFPjF7Ik0kSzkSNOqLFYx
0y3YOng9OO8hLJvlA6G8zG5QlbJoEoizdtCICeelDS2c0tfqvfMz/wQE7kwp
KQDHEhXq9i9TSw6v/L4kcFbz746kQmkPi5PEYGjj8ZOnCx3NOsCn0+M7IuwB
vUTf3egCDfL5XhrtXht5M6lateuIFJsGNYJpyD3Zp9dGKynEqPo7b+RmcKaw
LKdt5WctcMUE5aeTmYpQGJgHDWHqXqcuTZuATeBj/wdjtSE6oZy4EAaerTqR
fLNTcm31sOyuQx27nApPVAWnJhOFyqeJMbW6mJaUQFcDNbvx88KrjUDBH8U6
z92LgNZuUiLi4leNRkf6o+S9x1Txju1MUFBtzt5r19mYTDv1QhfOXD5fxNlW
fSiaupPUaV6ouQvt7MaC6e9b9LWicUNgfVRETSml2Yoq2puKidhqC7/hAk2S
qvCORP/5FhlVYvFFa2gRuvXtsXrkf1Q2ag7wGSEqCXtdzn0Lu6k5hROg2zJ5
YxfpmY5CVX1XEZgxZQt54g8U0tLSjYqwE5LZLPnttgfyAgwoh3QaubZDjopH
Qnc+06clFCyi/IROn4b7SpgWF9+F6Ol0UBJi4znGe1q1i+I2N/SL2KYVGUzT
Fn5IXmDCgBtS3s3db6ZJpHNWez4f0gOtzYG4fo/0ZE12vIaMjSd56yrc1LYq
wya8j3IbkfCDRa1nuPRkhYEUJZxt9hG6+wWw4l3zjxm3h54GoMHX7hljQUsg
YTJyOF2XSYlHc1/UYkV4LNV2WWkhQb4bGlDHJUF19QX+yLvNc8E47Of4AKHz
VZcd7OX9j/lB6QSSPsW70sKqcK/tCAHNwJNupRNeEVMUnACFdF4y++iBwu9x
KOpZS+Xgj2pjjHOzlISuPFODGcAGOm2a1XUVqL1sjo3AoUc11aXvPMJvDppu
3hp/S8q1tJsAQugOiKF8EpFlr7HsmnVsg0Xx3vz6ZlEbu1DLIzGlLNsOPg5B
xzDtdO1RYVsv7KWGfp2ZQlvgbZHYZmXpFrzLOiALPJ9VSarO80RpSQC2SG+i
8mYagcOZz+95XByyJzLNiUMqvtum5EOsI3JhEqYMCej1Bwo9AoAU3bcHbxlA
iTtRuoY4uyvONwoRIatr166B352EItmMeGUK937jMw4TxLeda1xoCFNkPX5c
QbVvs8LyVE/JU5fSV+uQTG5pIVCaNwZ9c6JLSJHzCKfBL8lSd+YUih33y5ca
CyyTMTK0ir4gcQ8ULGR6wXHtHOFI1H3MB5PC2/6Y3bKJDamm35e6Ee64NO/j
K3qp6yTXsNye8Ot9ZPZtROiHmRFB6dBycOkwA+EHW+kq5LdF2SwFwsG9vWDv
qzKiq/lcIjfkHwRFmufHQqO8feBl62ToEbQ58X9qhSMU2/vj78N41bCCPNfk
eS2fSvojNJz43jTL5gUdL1Bbmmq4Z/6Vt0HZjGIhLC/5gLWC4n7TBR0X9ifh
wqkIU2oUoKLNh4ywERWwgO0qgp3Y2vTM+IZtbO7zT6kHhw31hvmXAwMp7Jy2
U/tkma939h7i93ea8yxjq2X4eJxqbRr+TIl7AMe6y3Xuw6zZVEfurovbwmu7
VDII3TyLY/ZDyZF8Z91KdWf/eJsNyblnyR8sLuR6rF/GpxP9ZfNFml/xFwbQ
tvMzyYqCfK312KOhu0Blae/UZWugipquIbzCaBFPgrJ3F63WTKurMRKlDs7h
1Xg04H9klnCZUPZfR9ZJ9k1HreGmXZ9pmzHynY5M+3htHb6MznRhlr0AV8/8
1bLUrrnX9kN63JXlFYDIx8pI8I1LOe+1H18TcMsit7Y1CTF300L03DG29Bij
9DUB/z60lmIXAezIJCBWhjLPs9bpfxV7OhPmz+RaoDhoSDaur1RhMGYk+kgr
sJJPAm+qTDwMcJsNp8MuU/3E/iSQ5flre7nwbqYf0tX0uHEbBlIA/u/2OE8j
A4ZaTEGDadheqiyW1BxSEicP2mDI+HEzZ/HmgSd6I5YLTYtrWNjOYxD7Mq3j
pDWDcpja1p+zd1x00ymr7DL96UAv4iZdIoEkIdNfKodYlxmtnNpRg9UQwPJD
6PZSpQrGibAiWhd84y+WG8hj3qNgf7DnhzCUCDyAGyS6bLAxkfqkILvIGhTO
WTzH/cCBsxIgCogRBUdIrOfMOcIm9TsEz3RH022oAZ06XZS7jI9FT0nlURU1
1DA01CJ6cnaJLCAZGLxm9vPP1amSdlwgnAEofoDCpCb1YSS8s2LRczsTq9pA
xdbDQKPmyGl9hKpjyshoK1diw77gVdz4BuUrgAdBAiaHa0NaKX3brCkiZ1Ub
jeEiGlGjx72vn/4rpfD+I5sScR5fhkB05KFIqqA8WzjqIH5X067ZNUhHnk5q
iQc0dR0lngtd0qkY/R4UUSvmVWL3ejdVKWZDmeS+WA3BAAA2DkAD90J2C4k2
xbPG3wpjREhd3g2USyYLqMCU2Ly/zjSXy+cF6smd+4JuRe3nhrbryzXnv9bV
XN0R2j84orIw46i8qBRA8IZI//XsrWjMkv5H+1Hpcjm77twbzV+bACnmPBfq
fY22bh1cKNBosg8S5LX96I66ife+e+g1XHLJpPZf9kDdtYSODY6bNsb4klJ/
4uPnuR52uOph1HNtD9fcZPzFIYAOdhEjSBmAWpcTLP4R7TkMiFkNcrVRcjZw
Ck9Prw+wGkbQ/+HuAbs8RWkyH3VhpRtGC6Y2CMpeA4tE6NV6yJ22G/h1wBEZ
yuYsoYdEA8TO1ed6ZElZPi1uP1GyYkzDXqHENHThD1a1kpISKeqYgkj2eQiY
HP5F0+Pc7fDhY6dcQyzotsi0CoSWefzq578HAwkkF7no8w+E0mdDWnFIbMlf
073B+FBj17juWgCXmp/NPTZGwyed4mBdraocUEnmSnp72vmzacymxVmE4sDw
OnjT9ZWX5aepPS0IdBqDgXKEbQN3U9CrMsF2DDzJ9DPw9s/0LnXvSYYPpXNM
K9m1VtNlH8qlpiscvSUsMcfLPlKd5inaFoBnK/8BDW9q3q0qkLjRbcf0dcoh
k6Xbr5Hoi5Pmk6hvIFBNHVwHcr+r5mKJpCjSZEQXWoUwnyXvvqHNl1O/li/7
BZWIZ+g35odH3KLQCgy4bxzTlavkGCuakmVUbas0X4Z6Ra/UVjPyWljfldXN
RtLF3tT31YE4urq8GmNwAB/PLlRBWEfsVDkrGdi10xroNUEZ7EkJ18ZL7xAg
aelSFGSiXso8OL1Y6Cb/pcq20v4Af6QGCAyoHhTWe4w7VN9PiZg9yh+nBRuQ
LouNK1Bk48ehbnPUwuQ0+aWGw60+47l2V9Nj1oLKpigqHpdCkEmBH6CEscwH
epw6IdV2wxbgVJzOknT+A69aRM+59IS8D+EFehEP8Lb4qo8RE1VIp1UCqlKO
fJbCMyyT3mlyyg7GvlpxC2paLVyTThoFQXlHg9zG/M0IvhO/qdOQWw8eC44F
7+t+Ss3uDZKpYzXyX/lt2cDAGh5GAZXh9UHkC9uYEx8a42uDyS08pwaC/MJO
yOTaleLBPO6RSKDit1Tlu0su1sMwUhTnHKFL0z7ziKx+9Q89k7RR/eVZTKb2
id7Z+uG7BUaToAZ04fa9dRfWodZyABVdEY72ARHKTZT9GendTrwFCFkdbcJt
J8OipAFhKqq+YVOr6h9vy76my8c19EI02BywEwMOHm97mkw0Wd1I+fnADlMg
O/2C5FuzCgtxiMeMpfEvzsOxvOn+f7C2H9M9Xuye6y6MH49/yP1tTyuh1fm1
+3kedMCBXjoPIBuY5V0dJFzNjg2t+/1WrghlBa5pABa4wJWuGuOasN+ecSi3
0++8DmYibFo9SEhLYiTqp+wQvVt2Z1HJTUHDO/KR602CgeuikvWICqLOnJdP
KEsyN+j89IxVbO6C3IcwnygCuWku6M5Xy8WCzfGwyt5oG4CghKEuc6/8MMzl
/EUfxgI+yOlH0Jp+gY975dGw4gLn9003qn2D+5/tlrAZfiAqG1dJZFo/CDs1
npdFJglZbN6Xa0s7BTCnIdOzOKG/0ygG2nrRxRTxmJhoQEUPR6rqbUcfIjXK
jD7LK9/fnxBT8KlLux+eIj8CPMhkNMVkxdEOrI88lGVmbNdXN7P72+I95ubB
uwFt7uoUOFf+ItbaFkaLWOR+tLehZ9hp2t5HavL2HW112c/fMcUTsQJi9/AQ
DC2QUUiwBe8gzkQYQD6fDfD7NLhArCQ4bhfH4SkoOteF9tmJXfz7/ColWKdK
Boz2xLtXDHUcy/mp25F4zrECiOl7I4wBzXInz/ZlGkpJrgEeIDjtH9sNoI4s
qjo8WZ3vH5IxHVc1iu1HzhP3JOgrvRUmCtzq0Ky98m42Dh9bPCuBk/Spa/v5
K2Qz+WfEPpyM58EJJFgPHWaTts7SaFM7bcrM7hRzT7ZWOSfwpwEq/o/W7Fc8
mmC862QMlY+O2IRAeDPQq5d2ym1Na2e7vIxgpB9dtU7Lid/IYNVgaYMB1LxY
/K8r2l463ySXmCAXHwC3Fk6UHF6iE4LB6iSS4KqxIuSOs5hHj6rPAa7SK/D4
9zlw0O6OOl8skMpHBLnKBtKc2GeQhlTy/iM50XzHww4OFGAJaWIYItQlGMlj
FCNTJ4PGEzYstYoWGvEP6Pur+ewCpM0YAGQaxGNjN5ctWxTdDSN01UjH5Jif
i5BbklAVVBwZ/q3MNFAXd/0pkiDlLzz8PcDDrfLdeTRZcVStW8UEMlV1TH0k
gLleWrapzrRqIZTZBgHU8EKXm1atXlvcPeMgiHgDVgQOqOyIg4nxivrJ+a+z
aqKgFXA+4sCey8/kVp/x9RUvPKSuD8I2bQNO7vcbcxzABINt4xFlwIbdR7Tq
PATbE2DBCLZcYxVYTggXfcHZR2w2sDN3JxYXz12whf+vBrbhxpgus+I0bkPL
1NXmEJyUzzIrUB5YfXsLIFocCMsgut+Uv6QppKd4IHFuQSDiXz/C9eDMusws
t9yo+D8PWBiDXU7GwHoMBHBbbARzEhd16ao87SExrZGjom26AvFS3r3u0+wB
efqrSJI+4KXZkzZ40WlKEFxj9f+8zbg1doYxfXfSbtKdKlgErSHeSBnvMbdJ
W70xtF9EFHEG9wyWtsORGRyp8/Jw5YMYJOkCxDuxBcsoZUO7trW3hOi9EY40
fn3jjMgmsEnV9DNU3kw3aff1l9V/vcOdUPNbzZIwrbRQxJZYdj6j3Z3V5SjE
G9U6NgzXSmV8ZalaDQrTHXoKB9oFU4gLjS+lLZZmsjSlQo7lG+mdM9w8cyS3
W1FskQO/oV/6qkYUJxYv0Ym/8oT5NkPQY+0Soa0p42jt56UPRIXf3z3keVCB
sBFY8O0zlM19TyGRktVqFAjOwhvWMBEdohUza78VhytkBBIEktw6HNQIZz0O
SNU56IEU84pyov7ynFYxFS9jCRynrCmy3RK6mpp3N29pyyMhmV7E7fDUETXC
et56NVdyul5uIs1iZl01J9igzk+ioTwyf/r+Fj7eOlDkur0fyVfTT2GfmwAS
ptkUVFQahYF/Hhe0Ipcd4W1S9OFh39F1TrR2CVVT/IYSgUd4c9m1LcFQOj5v
cOrZdt3QpXBFS2dHl1j27p7/o6AellWcza4SA0Gva/hyACQqQrFv8F4fPJsE
DOD1WuyqVhNW/TN7qjhV7pyX/LU8rKsgvN8twL2LLw7oCL3T1pch0/OqVePB
j8g1/I+PdPZjkENEn7av8iIlcPGE+njycXOkrNKJjViJ9TiARPxNaeTdNr32
MEgjhtKAHzHWbbhZV7YtoaaUdbYo41aOqaLwLlFSbk5Zc20ToO6VJvejm49m
Rn8ph0YDbdQTU8KJiP6Sx0wAdcS2DDk4ND3nchrEQ9cj5ePKAQk7Id43DMMx
bPFfQe0MQt7GvxPmofDru/hBWNONMWKMwRhIsxx3Vdml1d4O+qFSte0+pg9R
VShc+sO8irYPvns9wJqOFwo5uomYDqKjPl6HT6BxMh6EyfCW3UMGtfnUzRXc
yhSslKnG6SvuZUYNbywlF6ymsESIM78csUtJyzrloUsyaq3qsBIWVLb3uR/I
5sHjSfEqnenfeqU4BUrbZHJgIN+6H3bzQcXjpCevOAFqQ4o5yWrFMXC4IGLt
1maqrMhoz0Iwk/ITIFJKTIMUcYIcYJfgdUaXOG32cqU77DWqumhoFBD2Ghf2
IXlB0gi79fW8XZKwlHOQvtYomXi9IQRy2UfC/avYL7GQYXC9rn+syUdf42oW
QNqA0cVIOR+4kCnpkWKmVN1FsN7xy95N/i17H8fbvw0MQO1fZw+sns3NQZvX
eeiwjFjrDZjB7VnjNIZIhGyV9QH3Rls+iZt6YHmfHflAsc2xnpqiUHu8bKru
CkWEv/zq+gOCfoGbZ/iGjaf0gdZCZzbeE/kO0R8oXxukqtCUfNIi3JdPnUjY
YucsCe2lb6mB9OJuMsfrMGQ/ArIJBK4F1qIl0+JpxAxBwVWZlHqnFDmXXYU2
R/Zz9ilZ5xW+ivn+oVyFywby1FHvoZ+hHqFfGT22DCrXIE+dGJFUgeY841Mf
dWXSrNWis/h1SdWsOuOZ7N5OwOYV9kiY/yVOyur0Dx9eoJbDfwzFRDBUfi4/
2+dw0DOUGXUvZmldCJ6KhL5K1GrKDMPGMWtW8BU3MEwOtHExuuMpVjKHw2k+
v2PAXEPrerMJrlZO65UdR/t7uB7oBf3cxfP8nrAZ7as9OvcP64nygYHRvGRz
LepWETWLWEuXXGYnJaerSt/y0X7xZtbveG9E+RUpWBfzXmcMI59rM7L1t6Bh
3vPpdzL7uUSUJrgMy9i+083jhmtLAIRrv2IRhBt54ZFPSy5Cj/G4gaZPjGdA
z17c2u9BOyV2cQKp9ZdVyzH0I+Nesl6omgSzGdgJFO5rei3igBouZ4Dij0zC
/3Brm8bqKxW4StZB14wsyjvCdykwNQBjIMD7l9TLcHwlZeFQI7khTMN/eo7A
lfwJdu5UgdcjUXKFAnQCektRNivjejBSEGYI+qqNp/LszoTICoriapDnAgqD
306ln9nAi4ZWtiAcVFaJhQQGT5UEWx8AjSu5/7Stnvv3LZhxt2KITNDJZmK0
yV+0WCeEgJ4U2ZXAuQNo8dyC9Wg/oDJCLlIC73fnVTYv3TFoBZRDtciWMAM4
der1LZLaGNb2Ia5vdhXeHbx/a2JFrtqDUA2uKIdLaPw0VmWPzjm8vylC2R5M
fk87wVHbMGwdoxK9h0wkyqGF0cJ3ZC+l0A3SOjXo3bktRpmQiz7tDOX6NwDQ
DiEVrp/KmiyIPAnESX2XhUwcdH4TMcoEYkh7s720a3F28ewSWfMTBECh6iyT
8I2jc+VHfsM+pRkaSX2Ay/XbDEK8Wm3d9Vzj5mHU2gZkzKjxEi4wLtvANYEC
dikhJfLlVSN8U0GfAHIZX74RF5Q4+lhvZ2h5/8iHXz1AinXRB+KJoH8ZtOWB
Zln/p6WCGwjnI8x0q3Crj2USxu6BE1n9ypi+hSXZZpWWWHn0Mdj1y3XHiuTR
muA4e+zJjKr/7kNJ6pviWcJ39Neq3Ft4pSGXNxtmpqKCqO2fDbnOUnbKWSN9
CcfEeomrwQH0MUPVoxXpetoD19ryf97c1D30013l7ZnHXchOiPR9VITUgfNN
L3baKiWnOG0voeeC7LwbsCncqrBjIwu+5BsJVUm6JQ9uafaCHvxD5DYDjbmk
IjaJtC9QjGgNmfMOZBOl94rWkHFad24utLBby5PJd/ZdaxbjlRLelYhRO3sv
S1CaqibCqR4csNVgZJ4uO8vHdDssVKBItCn/1xt0jp4+6nbkgD7P48RSyPAk
ddCYx1uh/qA8jQLozVJL1tt45Tf1sep6uhWMrrny/AiN4YxoKxbswVlNSFpJ
HxGe2MYSLnDxs2ievs142ZNlvOe3ffBu0NU4gzxyGOp8x2QXLaaPhUuMxstq
yX4opc8lpL12syjRzLYg7KmaZCBispMJKUnV/vSNxSSK119SPuakVj5fQVAx
CBdveEs9BmxOsDdPb5LQqeEHeTwa3nSuxO2hm7AZSyc0J3OhOlKPW0wdZVeD
OaS/bKBbsCSIhai9Ln1l6EZ6Rc2/wsFqnu63RZYoGbfoxQfxfB6qL+TqpDIQ
Do93D5vyRz527tmgIO1IpBiRzK/Fvh9tmvUhHZCGaRe/hKMu1qOIx4SfQO9M
0MDAcqc79qRdF7m5/XrnH49RHQo79a4MU5oIQNk5GthKKgLA++qDSmQIhRYU
p/FmoRG2eGkF5O1sYKuJ955PiHYPIFYwKpGoC/v7NDFBtTWO0jpCU38N2rph
MPImzv3le59RSJQfdBpW21nGE2Oogzf+wKPe+SMO6kkWw+rc0JsOafWyggRR
XMu1hPhGD8rFmHnaXWuDaKWciy27YE3p04lfTJ0+XUHiZ4Shisu4YWcThv0E
55oh8nrPY7hNjosQBZqhDECvok5Mm4NM0VQWIU0QiojeHdmMtl58Z4d683sr
TxQrRP6U6ZrZET03JxzN+UF2F0tSUxB2Ni3bKb7ttMkQJTYTMxJOU6mQdGgo
sFW5JyJ5KXttnUeDYHgGKMw1C55HG/bV+3rTWHPBou4lVUiHtPz3Ip95mBnT
xUSiory/uR/c2GZ6Lg88+thGTkvXwOUKaGUAT3kSYBgxCBMvH0K3UMKr/7Vx
L6w3Kjed/NW5fAuOaKt1TNJxjr+oAx70mOZl/hghu/Om/g96qYPkso64Hglq
zp5kiLAaU8ItseAVKEES09KZ7djYAs1N8TLS5I7+V70+WXTbQibDo9chIDMw
2mkhJ23jXpHl1+IYTQAAZzDvR1pYfr5mGAZn0Kjrd/qzOGLIIWCpEPRwKAdO
tkfC93SPzw8Yyj8MQ9YdCJF62SPanDRLTJmjrjewEGgE/tKEhC4yEMtWqq8t
pSZAIFJ0ortIIDYbVfmQoXSoMDrK96buAtgJA8l3UBcljg85pDlH110hueqo
vdzd2eRutMkn0eyS5eKMeGx/fMC0stL120YWbaphTJocf6OwoNR2fXZFjd1f
xt6496zv/aUdSOLYwT9365C4LR/aYGwz8FRRqVzmKBCX3yT4eRAq/6Rei+8z
31SppKfEcRAvC1RPC1OIOhr9l2LesUFdc6rQWwZde9SuSvyR1UqYXYu2vFx0
HwZRBXIItkqkydDq1z1JeHwakqZyHTCdfMPOLgRF37TZX5nO63mVNxttUIF9
bSjm31gMN2s5lW2oNj4wPxHlXr8LWYI97Uwm5NeDjj65+uAmzMngCCUt5nnJ
wxUPSTqj2QJnSGuQZrGTakKFJ9DJxa7qQfE8yVbCfp2ipZOTBVrGAn2IBb59
CAg268z/h4hL3AIKhF+0Y+ezRRUGNG6I8pcQ3Gn4yoxEktmryZ1dbiHzFAHg
bizvOT8KitY8Pf1W0JN/03GXejFsPkJ09F8z9GsYWGxadDriG30NoLqfY6aR
vLl2Ra1efm8Jdu9kAFAitzHRt3MEAL8VRiY574smJo3aEvCO386GD4QoIt9r
XD3NM3gEY0XInKTzbxS/cXx8maU4SC4l4BrVNzmOP1lWOFhWKbYU8UPoKmV/
tdzv7HIqB0TuivG1GpfHtI6QP+kEbq9EWQtMUie5v9n/yCXo4T0sd03/gZWV
jkkujVD6ZcVwjse1WAhx9L1DxPZACxHTCNa4vxdC6dP/itJWfz9wZM8DMivs
ktE7k8P+DKifCcfCBR64b8sndH4GDqS5AHJvI0jjapQU9ebu9cdEhY2Jyh5Q
aDuyJFtqJQh4b5e/YTAMudR13EDEUng1iSBkpt9ZM3gOKir9x3X3J/crDgrd
UUhD8D5qu50JUUlf3fGfMX9W4wjgWh40DN2kAH0syf4EtmiU4falpRe8T15H
XbYPvgYvMO6Wa341iayT8NxcKmU+QGKUo2qrGYgP6AlDNkf7Ot0nSOFSk2KH
4YSGB49F3kK83fgPT5u2W5oSvwnrhdFZ1g2Ps3GvfNiTxU+tXcuiVwa+mpTD
wLxGY+78VgIzqV5XTPCn0q4GwwURlOJ7UN8Go27OTd4gsRLbqaa9e3BjuTiY
V754zImzkpkkSzTz8ufuUHxnHYLYeVVw2jKqLXqgfC7WAV5/38Eu3z0Y7hVa
t/HsQBz439M0EZ71t8tnBgdamzRUgw2hXjoSPWhX3AUtXl4yY4Kj5i8KNSK8
EM6pijBMb25v4xr21kXE30fMorB/Vqya4MAs1+6vdJ+SXL4C+E6aOr5kng+J
O5J4uFDYV62oe6nEo1Sucp6Zsf7U9SwG+mwB2dH0AwU/XYicgj4mPYm7Klc0
aV9y292fjsU125RWjoVOI52gIYohMZSCA3Vcn9Sj2iviQj8Wzkqe5I29mPcK
9YcDDS+dXqWpR3PCbqQF6TV9lLfO2eDYIJK9aPN/T5TEfEDMQUBtbJSab/6f
IYQeOvPDieWfTSEd8dnZXkRF7WHAf1ythY0QoiY6vzQ9rnzAEjqIiJxgpF44
+Mzow/egCpO6VjLNN0q6RZM49jX5mZFQTfZMewYzyXBgEd+PWYLh+z/Uwq7O
aPPmshJUrtjGYCLA0q3BMStq7TEHL0zgu10EqxPEwR0mOMzZWM24+B21O3ru
lp3dqpbhmjzStIBLsJibOgFShyGgMtWFzR1z7PkhWsca6Y9J6DKJ4j/E0bQM
3FVHDdVsf2mhxjanghUGLy08V/wxsGS/xe85M8Zl/iQkuT6lQqXk9mxjBiwZ
y/ZXtDsTGAvaOQe60VRn1zVoJZOMU8XH9jHjZs7eHvJho0pazJv7Mg4CjZZC
i/Nt1IIIs3eq/y8DJN+DVtyH60oSUMYtM+KlEEOL6oLyFKKmDbWyuGH2KBce
SWIiJ8jOBQHdcYzm4rJxntuOwD9QCM36z3kbFLgrU+CY7UmeOrRWhsrbwC8M
KXjw3Sr/oqJwhGGA1vA36+E3F5XdHJaKM0tYECMXaoJ/eCj/3xsg7tBzZ7/g
Xk6DuSK1yJMQufYV94oWDh3U7rEmw6uYvWsnBGqP+g0XZVSJs8OwjsGmpytG
MR4hWOGlmaw6uVnMF0Es2K08WvXiA6Mk7EaNYxsqdGfsZUfatcbQwP7iOZy2
CvnRe7XUY121lb+eKhjF+ywWqKgA5OyZoKkMX0I9xfjmnxXcAAOA88BURFWw
ljTbNtJbPpsNJBcvVcZldtzdW/0TVLY6rBxZ+wK/SugZsaXc5VjfKxajCt1T
mNZC04V3ZExITYnmspIg8QtWQaXft+dbw6kUQWKHNsEoyE8oI53XnmrZMVf+
HbZ3cseKM8q3eO9QX6+Bb3VvOSh4q+u8As1CTUXmamX+8C4rsZBKXARYikX1
myTyTRZdwOKdclJfxyPupfwcQCHFzJX/VXIXJW479zkcpDlUFY+5nmyP1Zgm
sMPQtobzIy5sa9txLTO2FrwDb/glzdpANDBoP4SJxf51F5Gj0ZFs8AdremnD
Y50S+G/a03kU93DR7DsxA/I1PJ848jL7weM5rezP35MsBu35cepkZ4PgN5Wy
AH34KpJDWliZmNCqZw9jnq8oD/uN4epZndI/GfbpxloPABdn9xmvpj7Dtr5Z
KSTPJ5rZQGOy6IwEAWUpqkE6tMSB3y1xGLuTEVubBl/ErshkABzYFWhHnl5k
rebh5nCLc+MWhwQsn+u9F4vKpRcn8x8yO+WHme/wIyokgws2CalBt5lnjoYz
FvhEzimwUEdKXMwBGDxDjQVAtjwTHIVdG9exeSNWf8EtGsAbui0QBA5kgkhm
+wmyZATEAlfLlePFYazMviOWPeSY87XUuHXqTlxnuufQ4aoCMkBpdKpBWUou
XrIne2qkoMOg6hHMivGvardtZnTw7XxhyEgBvZhpwEuWXex5VG4u/riaIiOX
Ya4QTI8XLJBNin/OCwFmS1K+/F+jouVZiPKf4/xk7OhcFHfFHjCN/YmqScKz
00LexBT67dIqqdCR02UDWQTLwkgU0h6ULGEozYV6dHluyEx071HT23u+Vp56
4oiUsMWfg2tQW+02luSD9ip4L4skDRqemAApUrkM1tBgdsYYvFzIMe3jDm7F
JK3W5jf6SmZeM8TyuAdC5G9ANYGjEGDtE5nWKgIfILWpAK6g5Ox3snBHyl4N
e01pxoD3SLLjxHblXkRXCLoRriM4EU2MryDepRGj8U7WITNkaerttMBz679b
ojnMfdLrxfFeEKQfYeVx4wjcRoOQ4RpzQUGtwSS3xOa4Kt4khT8goV98V3nx
JFqx5uK27XDqqFtXWol9i6qBQ2F6B7qCZLn56+xA/JRyAhMXnuu2pBIWmdzf
hf5VOi7EdFFsTRxtaoyT+5pX9l2s/45yEjoom3svNpdudPG1p60wOtK1664S
J/yD1imRPofk7SeX6+MiykcS3bTf99hG3ql6b8QnWvkmHyb11H48LTGnbxL2
PR8w4BJKcoc4sy1zzxapRYItnhEgkQ7NPi5ztlU2Tda2yInhc9HeyDCTwl9Q
ApMnQ2oJU8kCOtSygkNri3LDRTvLpjKOKetCBb8/WlQ5ZYw2C0LDJKTrWv7l
86NtsCG5k6gDK7qW2h43tkZiS7DrNE59JvxY9AMtDqw3WpQ4jby4Nm6xoDnR
C2ay7lohNRinJka1ROy+ZOH4LkR4uQ/R3w4MbTQeH3kqZesF+0+sczUD6XMh
NbQV9KbelRHwaszmK4QJ2WI5hwGDD/w+12FVARnhYVf0mRalsWz02SBRuAsW
lAHR2vVQBVUi2Lw+maXysF+eFMTSDE0IP5Vg35O0/8RXGZXdBHCHQFpwAKbT
tDFwJHvBh9nHOKzdbBVynR6WV2BE02P71KVz3q7Ht745YlKFrDvw7rIyE9jD
fwgOu2mRmuGaQU99LNA9PL4LoWF+OysyxhhFQwNrKZDQrxUh3QXit9BUbu4u
q5LrqtWxf3W4ZULOIz0owLD5aZKifW2rHLPrB27UvdtW3ONC3wChAjKhjg0q
FcMutI+oDlXf1FRyn4yQbjoO1Mb9d4O1XUiZxxxZtZCbC2cyjBRORBZTHxwf
cPk4ZmqEGDtsc7k5Vec9h0AHPmJqZhBJiiTvRG23wA/mi8dBDRZbaDKJ471U
M//5wzx4F4OrdpwIUbjcH66M8ZZAtmkHO2Ph0/8GnyzUroJmcOJdb1cD1pRa
PHv9X87M87dLCIpFpCNrQLliQqZfAeeFbVYBU3V6etH26HSUHnPhWPcD91F+
1kLfNcvE5WFX2EOpLCOjoAtk7wvc/tb92I883zbQSi1VIKIzbp1+4FDrUxK9
O4++rOxJCG+F2a8MGMrXyrMLeOFUOnyPdsputwH92R089mlWRlmuhh46IMTR
5Fq7jmTy1xXUa5wEceBukm6C6JGIev8Zb5DLYyxjT5THl04QRmHwRDRx9X7Q
AsZxpwbvKrM5iL+wU6m+4EtNUdlNB6S4KZdCQhmgq57y85WoZ5tYjpNpT0pJ
LDByWfcvkHrtGyj9dIo+jJez74k1GaxQu/746W91Uwk97dDvZDQliKbJ0RC1
f1ybGIYim0IsdUFdbyOv2iMH1HrzncqxoWjni6BAnozoOH1mFKjnjhHZ+QYe
LXm1I9bdXDpknh+FTKfZpvTtJDDmUDAr3kW6AQhCjMq64mKmZQpuwFBsqEob
gOT2/AiNgMxguxb4eiRtPTrGuTAD63va7Q1imZ+5CgKewMuUiOVWW0NnGM81
KZ0KOHi4XxUSwSfffvKgoOOKj7l1Il1ckVXfbtmtd63Susqa7iikU24XcY2z
TINEofwSaiJs/1NQ+TC6tDWx2lhXxmnw+ixDT27MquYNKDNdHUHwDyNUmGrt
0oblDK65wSnW5JIMtuiqJJ5z8yzMaQli/G8t/5acMlzPuImCUHNKfjE06q/I
7NwaqF+MEcfGKlZWZMc/hR/n9FArCUK9xH+lgIezKC7FaTpUb8c+ag97tXnT
10/iQJXm8izDl/nkdjChAOsjJSCSwaQUT8TEz0wHUP+kgug7Iiviv9uXoLYG
S2jfKtRk16N9L9v6j2hpJTwWpW9221s1SPCA0PNUIkPY+JyBEgMMOAhkmr0l
ccrmPWlmnD8T+1GYyn5DT+v2W6RahKrj2yLRNHFQMlMw1uPTdhN4768RPbuT
SN/4Ux8na0zIrY1uT7a6ODOhaZvggxHV4WpO3HhpNJR6ZchtEL1htwWDWTqk
/cy4cJU4f08Hr820ueW+FLegFXK48zRzJqKIE+adwpIPGWPySpgZVnszceSF
4QInFSkCVugFrHACTdVF0nGsRWcf0LiFqO58AM/rwLrSky1FtG4/gnQqq4zx
qZmFvcUF4S182KzswZcZmF2qEMrjNQQooODDa2UwktmKXEtZMF5AWerjK7HA
zIx9wnNdqtrbrmpzWR9SOtLvCYGZo24Bgv3oZkV25ZgV/RiTN8IuT2H0nHbm
ZDZ04cMjMxiuifHzrYOl8t0B3GiN+P+vZNSHES+ElOzxwoSrkVVjaiSPkQAN
pIUUyWxHcsPGQRjg/jQP3k/qySoz9jfOz30AXsK9vaFH7Ht0qUZJuFTU656y
CCntOE/cgO8P9t98n3Iw8/HRxe9MnJmMdvQBDOieZVMAJaGO9pZGInGPjqOp
gEW6t36DWYDyKLvIfJ5XSTooDtiYwyTeHQY/EzjkXu8WGC6Z+3Ah5KLqESvi
ngqxX4B+yH88Q5Ug6QJ+lUlecRK/8qg12v73a9XDdeilikSkhVJb8NcBMKNB
PWkLivVX2sZj6N+FkcuWTCLpU901thWUFHXU1u6mdeaE8E5ujgPEHjTIwc3Z
Ek/MWJcBtwCneiHw/dLVe5Z4HijgYqJRuPneE4BIvu5wQtZUJ5OjVjB6Z8nT
tbCzfG23nicWIepfZ+KTNfx60MlNM/3RGFUHws2NiUqEa+8hnnLWuek+/Gxm
xTnuEIkVNjb7pGA0iHLkQmPHHL2Lz7i8XQ9tYJj05oawIMT1DooUpPASt4eN
qezIrsxF/zalip5kmdaK48k6FjVGXBddZtTyVb+BwZ7WvVEQkkrL5bhAVoTt
F/c5jkIa9nJ73EUScwwr1k5YA9J+l7JDQAZrDttqQWa6SCeiVFvqM/M3MmNA
9INsq7OrLDlh4ToCi02UdtjUREwW7NfIYg9LQrOLn1QJl0NmVYTy/P6FUI88
LZVK+eOZJg4Qq13fe7GaC6f24y1VuFjZ44JMRA7Kb2TCEq4ze6s/2zpolRzK
B6wKoWo5AHMJf2rwOLHDK98If92BHcJRDyF50x/LjZk/oQTi8Y4BJLXzOItF
BO81srh+VmMX7c6+xhDLCEh44d1tXgjXhpLlkKWARc4GL9QSmBTwQd51+0Ga
0QbLdiyoa3FtCoVZ5KoRvyIWoTQA8WHgnVxloiXBx/GiYiiAyoVmCkXhZNlN
wa2LkNdqB8Et6KWayInQdubHFwo7BDZ+wyyhYEsHlBeqIJowo3ujVT/NZLoI
rJuxC2CWPhokfkhrRCZXvisZ7/WQ8JUYs8CrQGzL3/BmmJyp23qjv4qc2YaW
ufF8oW6hGK8XwtzVwGOvQyHXe/MYGcgRccKbsv888GHK92MMar2scK717iy7
CM0IspLGb0pS//t6IHbKkQ/kub1+No2+bre7nsVVL2d6ZXzUKn2iZupPXpl2
IWDTHpWhknOgpQF8F6zfIAmd3IvdyT4jfxCtYrZxcK2hAYm7MNnBF+MNm2nG
NxpCrmgaw01WA+aC2voE3jSqEdbj5xIkKMmxnhadY/Ojt084/nDQYB0Kbnx+
VAJhzitTMYUt9kUh3ndgG4yujenE6CrtOlb2EGc1KKPONmi3hwX/NgSF0SJ+
74xZ7mHop0JqGNFJu3PO+i556veojDaxOCeqzKNBReq//vB2AXfJFQlVYGwQ
j41L7aL7eacSG7n3gaGqyvTfZB/dAmprBuTEZJU/Kches5cGjKEyIy7Qs/Lo
Pj13xOUvuOYQvsFZPh/yU3+uoTkgzqhhYWl431G00s9IFgsxqO/O1ibcu/VU
0BWKKa/9pH2RQjaU8oWfb4yaMhahfV9uaR6cVzl67eVwaha5DFwJw7cM4hbL
nJ7rDuusYB4uqoxL0rMTkNpaX1yz39xxj/b2MyunDtqyGd94u/CWQsetMxsD
Hf0umjez36PvYBClLem/tqa/H7VOxc1OYL1ZPlZ5hfXreca9Z3w7YbDzStAg
tBC/nbkeJ2T3Ngf1bxt5DgPc20a4qwX+L1IAGhs8CsCrVgPgbbmoihkaZ5rm
R3azVGkCYdodgvwKUhmfJhKpiiR+LnzT9LK52BxP5W0OznSDN5p8/Zqk9SGQ
JB4etqHcxsFknY1rQ1fZfbIAxbnrcPCcmYROwycNhvsdKhhUeOkSRJJNKV7G
akUYCywozPF8WZrWT0agFYJIviY0aatQKzlNywEQoi17syuBqr+nm62mwEXX
rYFRaRoml97L9xVhkC3GkIdVIsPc7fykN8XdZiT4/06QvlDbE9Mn6ROdnQHH
x8L00WwU0ODLc9k5qxgASDnSrAFUyp3UA6yG2w+Z4wg2splaxx4Ce6/blGOW
zzkdvYarFHmk5eY1NzgI6H62gYUiSiAhY7BI8wpkvMdUZpBLElwKbLV26B2H
offL5zqASjguyT0M3Q1lCRNWsf03Z/rjN9NDY2QPQGaHfhHK2ItkSHhF7dFC
E3wKPBLvaTuH2VBGe7qOk7+Xmwq6lsB6D7nGEUY4lAdcu76Amx7mSkQ3Nz+m
AX4tJXzOF5y3v8kMIa6LeRtaxUdNkpZ2XcCZ0XY3/dg/Cq4zBt1yWIp0N6Sy
IQhida8Ll/C16PBAQC+XLeeSIYRSelYq6Ara9Css8Xbf70i86kEx7k0+zA8T
QgyyTP0B91AzG1zn/SlsePCN7BeXGJNLQI0nu1VVJ+SATokI4s7/fau0BXo3
C5GIsfK8LtpkZ7fLw+I5vewYEcHxSC76ekvHBwdWpw2xroszK6vicE6aUoWC
9Jns8WaOcYrjzT3gATbNYSGgiW+MD3Wa9dei2Xhx2XlAZyjDxVYDUVYV5xDY
3kdzFdDrZ3GsO3Aiitfbk+0o4zvcmDFqrSjwbU/W8oKImTEIaJsTlKN9VVUt
OjJBcn8azVt02L99RxmsJuMEKiEKmXyWur1lGH9fFqRmmYjAES54yEmbtMJ5
dknnTOFVGAzXYzy1urdJQHLoHPDim0yGSitVE3TCGTnD9KO1S5fvw13vkYLD
FQMe6krMtVg3onBX5j37KUo+7q8vtyn64+nns+HpW6borHQm8ZH5r0nS/+Sf
2Tnj1mfoQehl9nGbivRBeBRWsB+fsO81bJvRYtg33YTKHFBTLsRi/rKlo4h3
nnlQDYY5f5O8DwEeZGV5hRpbU/vw2hxo6VYi23PEk3z1F5w17Y3btLS6jcB2
aX9b3rfyQgTWxTNchAwDXixDe8I1P0gdyjGuioL0pekPy6nwknNSogcljgbz
7Csg5G34zL4ucNy78HEeKhZT5nLlE3MDyrPQjeyFsZXk96f+XJ/reA/vbnmP
UkvlgsC0h25xPokftpGKy+skn/3vAhmY508eVrpDAcaHDYZFbsc9CThV87tk
uGRVStNo87Clpsf9Kd7dvH2prgde3ZWjhDjPWOoUxa2yGFeR8QjbmHgATGGg
C+F96mhwrlWNvalqoz2XvB+SnN4Hy2R7tfYBlWVbh5XHrYmvhy+g1uG0TI7A
6H6S9LxjdFTRKuILJdFfC1wqOOkVqVf8obtskn1ZiAXp97QvKwjnUJc/Vvyw
XNWAAQ0ptgR/rftUOicTpev8c0UVtN83/Lv6tBQsThWFbOv32NukmyhYIx35
+JmOfX1s5OYe1cidFz92D9JAo8+q4nj+Z9CVxqmCY757/B5jZYx5soxLeT+6
FJTsFHVSghQx4wDwd+nKgy9tj1aVn4vMXlZfAHDOB5tvdaGQNHdlNU44gT0Q
+ct+YD+KfOSE17/ZyMpnMP9aeA7zBV9b4u8oF6QPhrCO8ah1peMmCsB2kTTt
XIWU+vtaBlhhPbtHhtgTJCo2D0PMcIKEU+V2WAmS16YhaG0z6ylVge43H2d2
v+4xCnlSJMPbMDxoqcHZ/CxNoRVdmgHp7zcIL+tUo5kYKWn3iHP96EFwJYG8
0lxgULCdSXz30RwEkv2I25ZZ6oUi9QZ3M4WtfWdzBnIApCM5WgZx7QRMe2MW
l71Q649ytyRZ5XL9PBQUnk+sZpUvJ5h/mtMK8lAWM48icv1nO4U3QtxiUCkO
QB4a7f6/h2Se+vn5AUqzdPuW23b9NehPsvXNqZ7vuqxY8FH0MmyVq9Y1AdIK
qeg/2SFRYnyfBgwWuvFKpESUgHfExnxAjXhnO/81UlpAN0u7I4FQVj+Zt7zJ
enzy/ov0yXN9Ts7K0Fx9oxMa6TBm9e65ZrryrC5kgWKOXcqnwQUrFIeFq3AV
pZGVV88SUOM+eybSGYoMP+ZaPTljdFDjEfeU2Dbi7nUb+uAwQyFFvxOL6AYs
VrVbMmq5YWb05k7TiS92Ij9vrlpxXbIpf6tSsBVjyzCqiJL2k45l2RPr9fN+
Q6OzNlPwuFDMO002zw/CqQJM7YIBy9QbH3nvZVzWlcLHC6rA1EG2G8cPwhCr
jHp+nGz435pMV4zximmRMMSARKcK+naBCIUqmOA5gMV8S/slmeuxUY6MG7X8
AHyFgxNzCnxb8v9vBuU/SuxPBQ/bTjpj8odPVuf6/RWW1EwizcL6ste803bE
pdyU9RwB00tfFQ0WByv4nYEyO1Y+svo//fvhDSbHNFd0SgnCRET4asyyIMHf
5aipGGr8DaeQujXe5OWEHz7PnEziCYuqC0SjhT3XIYV3K4SeKYIkPHL5TQIP
upOjadqy/JE1ZwD90d27BGwrdifLauVQFK0GvCq5MI0Us4yS0hfVN89djb7p
BOYUfUH4ohaCBh5a9CTjPPBMcO9Z/0rBHa1BgBNv6sNXOgBZFLAIkcVpYM3s
DzXqkn4wnUj/hB7r73zqI3EgJM1P0ksWANabEp4WVC95Xsg/5mA5mcWu09QD
4wHHkg0493P6bbQ3OArZEqz/aIKW8uBw3Twf/ZJFFHTnyBWa16j5I3z4lnJ/
2JhKPsKqLvRj6EX9T5nxMEwavpBuC77UZao8q6TWQO4htiV8SWNNT6CoDcsY
dHr/uVjylBnjN5Z+4R6KKzaGw2rlXxGwFeGnsr2BpEZ64dmLrbWVud1GBGEE
9/8oEu+swSHcyh6P0bd2yctdfbYDct+hrvZL2ZPw3RiYvKn21pRLYeYYrSmW
UXGX9qg667OcKc/Je8x28RtdBO6u7L788miEvC4wDRwy2mX4nD2QLIwLh8Fz
Q1o+ythhJsQHAKr075FrMHzhd0P7dOIBLhZ4r0BWaPXPYj/wDOdrEbe6IK1x
spjRXZqHynvAt1XjZy8LtuVgQHuIDuyYTL561O5mztrsm/FocF/WEUWfFEdJ
a8rpg4wqKWROrDgyRz+I656LHQJWi54YjOmXbokURL0NdFhzSD6vdbVCu9Zg
LC+rt60kRl5J0k2ahYs/gCf2ui8u1t/qvC8+PAUkmNvcJ3DVbmdqmaMmEODj
BjqkfBnCD/JHuKepdBkAGx2zY/nZtVfoytgLfGmLyyLZnWvC8u8K6hO5tQfq
WQ9PUTq/fZYkPVY/WzYuZ9oaHAoOFqx0IvmzL1l3wosuwtXw2dAhdvFRQYc3
/6xVphV2NPqwVLgPzfxRQ94vLpenlmu6lnRku9elq0H6h0bL/cVPdMOOESdM
JpQ7U2FL5EkJ5hST/zIfNjuWKqJkjDfxcv00hGYLe+AMQMkciWtHvO0wLX0S
t5MMPdA4aNn9n06Dq4h2oz8yp+BDzoFt1O786QzU8ULMBntaOZ4Zaczwcq23
r91q2mu9chtD5BV3e+5xLXaAol55ePMivw2QXwOEeUEkXd4Om4cIOKo/wLhb
9vlAhf/AEsq3qDd+8kn7bcZQJDq/K9BqGTtRC8wHYt8xObm05zq7EltrdkSa
2Rh7xdmSPciEMB+LdT5smeC7M24hzhDuqqfttQjLC8RvaNvF1o/nXdtgxC5U
duO2uyZZNnrs+fKzURLVDrVWMkkp4AzfsTh8BdZxL7gEElaS6+zwdgSC27Jb
iqQ6ay4Zwh4BOFmIFBvr39TLUdCEzzxc9tBLKb5bp5wJTe4WXGrYLZ04xJf0
6H6TioTkRNu96pUUS16xMd70gx7V/BF/9ekr1ikW9li+SqcwwcU5QpPKURQA
ub0Eehb9ncOqCubhADAvHmf73p3BDb+m7IVxwjeqbpdJ2PncfRZ4MvY3cOOZ
vTWhAjHFDCF/Pwp/m4QV2hYHGKfuqAoV7Z70p4UOu3G2kR2oUeSxWAlf8Hu9
DkdIva1bNLAhCmqRo7fmkLur2YjWlOqIZyWm1HjoPMdouLHby76AA5e7umgz
1DNdl2Br/nvclSRDG5rbtpZU6ymgn8WVc3/fMTSe4fR8i//q1YTld5AFBqNN
QOUR5USHjFaMtEQUzgzkmEDeneq7a8JYMrcKIHhzPG5Tqb1n+GfbhahZXqJ+
z5OVotseCzWcw2PTwVrn1TZ4XfIQQXzCwZi99DFYF31oWJuENts2daqC3dkO
jx+3lX2DutIHNyELWHz++gtt6pLF3rMwgCXO4jyykyVg1GOOpQ2bZmbK4W6N
y/NEmQf/O6gNnREYpZefrl9tLKrlOd4ZmfBYTByhJL6BZlsaXoIZNhoLQ0+t
PYuKeLX1Xjowr77zabbzXvxa8d0KgdF30PWJfZUvcDZM09RniVZqa2CN2cDJ
cmEmNF+BIfEn5Yjz+VF05wL1KDAYScHMP1jgWIFl/y74PeRA2vo4KJLtzrii
74um+dwXiCw1rC5uZW/QexH3736pxRfT5p4cURIaCNAPbh1lddoouG4jgvOJ
SClA08eZhEWOhOM38O8hfZQNd1ZCC/kp8G/qV+JUZWiB3qatTFJFrIdSfcbw
yavCzVP2wLW8oJehJ1I2LHWh53NfBIZj17spBj+cWtm14fs3DNJZn48Z8DKD
h7rEJ/7ozaG3tIueHbz/KKoe3Xp2PxOHzrW7taz4tsCweeubdPF9Rpj/TMzp
NVHzE6juLMJMevHogTMBUQHHySyJ9nBRSUOhXdtZGcz2cBC/fmVf+V9hy5DZ
xWtws6twBeaKkellxWYT98LxWam99v50HU45l/R/cxXNHzyT5DBxh6NVzXIu
OPb4caHqm6Awals5kJr+6DFtKCw95l7usjcjYA+M5Utq9BVV1FPuebZSQ5vI
uzN1NQSgkD6JDA2d0ELaC9T89z9sop/yYhkTSJFbe5BffGFSjRnADrvc0kkD
L4/l6ohuDHDHsY0whI6yhRhl6xUqWQrt87j6KH3rtTXJsDPgXLEf799CIAdw
BOiifYlDMlnEUzm0MTcMFp4nP+bfHVqdvQZt/y+4X/TaUpE3rQ2L7I0H4LQF
OwPzPxcC2byelekAk49cfof61K2crXMDVzLWsE4VQLJWEE+D2mXaE+ZzUxaS
EU3mbgQesvVinV1ksrlZpEXPQHRWoUUsWna5MLpABUDU/fPNoWPLA8GUxOe7
+RVJbXp1VkCUkS9AWXL9Ypono4TEOIuzaSHM60TyGj5ddYZz9ovMA/6bh/RH
WkUOvVLKtc6hMF5iAOckaUbGR8YCHnabdsuGrexSCEk13l7DK1WzHJQ7IO64
+pxaV1/s3AtEgXQmPTWbCMEsVm16u07jMOvZJnMsEgefjRmzFJxeYMGgGpZn
bxIXWQywji9EzkfxuFY12jinWnGh7sGCmxfhqhlyIjBAjYbSH+l/yAtBgMZ5
k7iLeh7XyjBdbOXP2ElX6MkXUvFjLpl7p65FE7wzlSKojXgSU03pyhfmT3Po
aO+ek8OJH6+SUvSEvggrXOCaKIZ/PMYatLECR+6Fe1sOeFeGvMrAcoRaT6iB
Sn9AYMYPxhxCd38YQHvQJJ9AZuoavqbxq37Dk9SremCwEqhMzQxrMgT0BKY0
4M9th80JsZCi4HEFcnR5QdMkRrvUVO6Exro6pabI3S8A7YfGHlfeKj1X2kK6
NDmcb2JBaHCJ9XhV/5L4TnCbJsRe9Ma92ALEPQnsjPoUBVaiOmZvnT0M9HCs
JFAdpGVZGCE8kegY+PA9V1L+EsX87t0PgTk4X/NVIX4qYL/46HXcc8U7FG4a
6PiHFwgQTKsBb9rY8dIL9NAzF5I3p3uXqUaO2XQFxVggQNGH4U7r6DeSs8Mo
ULOWm6YY9juPOYzkMJRIz1HysyK1sOVWgot4xzsTvycq9esLcPYQuJ1sgYMm
/1zsZIurp7rQBwnE03qGRyuCERb427fusErHItYFq/ynE7w2w/LnJxmcrQ9u
d30OvnoKuGzvLGftd64+7XfI9bM4eshR/CQcVlqR1yDVVeCXaf7rO+kpFgmQ
74+TaYC44afk/wrIlgnNp7vtjNkubZGmV9B5dBsVWz3yEQA2AL87jDlheux9
XNpMq0m8vCHQLWwVbveJ1+DAmMcQrgTLniUvFmshAntmMFSwaPE0Q31PkHK4
/VIu10IvsyT+eIzQih40okZcZeS2ZGGfJkDdLEpAywNFdBaxX62J9RgAGxBm
sts5Qf54dsrhoCF236GJHvnLtLv9tQLs5crZX67OB/t0VQ2W7qcGkvLzihwy
LG+mn6SdGQXJXcke2PTDur1l2lu4tebnyRwSFz+hCwqPTd+V3j1YZgjIl5TH
VyL526QYf3F23JxxipDBSvc0P/Baps4Z1i9MsyPxZuVTUc47GEM/tFat9Z3w
v41r2ppzERbC9EHXxEGgCVJkky7VO2ou1O7XctDrOZUc+TfForZucUzbiYbH
ExzmqktJ3tBF8kFzOZ4GGOj4p4oUiJVVUp+XULyvi0J33PwPoIoxBFDMHVsH
cO8erkOQFZ21MfsKe86MrKdL3qDYeqj6bH7y6kTvwz/CdvApXYwFYfde0qKr
3EZQ/CaIEnSu5LU7BmQcII8woENfRmrAJWi0/JB1pg5p5UJEF6aTPULim37q
rbjd6MzMNOglqCaUTUCKu0b1msQeAuMC1EuKDvUiADs7i9U2QOVPI+Q37d1G
Tc0KLZRvhmDpkpO6L9FIKWQ2vIWSralZ9APHb6b+IC7onyBrkoyp4tv10amF
2+Vr33KX2NTx9tnzN66Mar/KAgD40Xz8mK/e5DNSg5rMWwN7BRffopTfaSAb
U4EOwxUuaopJdljePTONmw63va4ucsZLOdprjZLoyKvkOgmHmZNFmbhgXUcj
REWB8X3PxrvVVugd3hmilN+5iw4eBaEf8Cw88//tyCtaVwMQKcn0Mesz4lB3
UbMv363APyjfhU/KVouIG7E0h+zFmRXb44RhHAoYGy6nevtGELtQXNsk2zvf
tl4kpJb6YFlrm4H3F+Io3Dh4aAou5U8Guy26uAZBEwDjaibS5HQ8i2doqF5n
MkszraeTbQnDcScOkciC5eGaQF1uD2H9SGZOpn/xCSGI+X5mHirXZKW/OL8r
G09l2CWC0bsDr4sguwm6rJahXIpJKdl7WzDT5dt6qAVy+m+nOPNRhn395y5e
RXe5ab3ROzll6HzUyBilYkl2aPU1dKaZxtXR+w9rGT0fxa7nEwNPfpTFEbKu
Q8xC6Y9qugqT7/jIi+Krtpo9hRJB/0Lv8861Ov9ruwKmMFQ8X/ddvQimLGbH
XA24pw5zbuKNl+rFPS3FMiSuF2EwyKKU07uZQPxhJHQ9EhbfJJTbdn+//jJQ
5nkq4NQYr+17h6EAWphCvUvEpXQhGxFXI8BTUMUn9+EDquuZvzOzMMCExKSb
bZA/Vp03ZWNkW5IjYD1qjcmxH4WBpqr5U4P0PRijuPGVJvG6vRM1dAjkrGTz
hGiBybpGFpdBxpu2YBd8t3RXDjoOhp+UQb9a1V3lcnmaqFv90Kt0Kw/C8Z6K
U9vY2nQPXCz4aWlLbkq6BUvLQGlCOgbDP178VwLGncmENyrIHwSc4aHMSPw/
EaVGuKAfGqnONJsa2+M6GTzaRPeFd6iAgpSpaxPzFyXW8C0AVEx+1SBOAPDj
CyYV9aR0xpf+a0blKyyfpOxrlhjjIS1KeS5HTugSEBfK3Yj/KKyVZm8J0ucD
P1dR21uMla5Lfo65pWrxzgAo5y4q3aJBDPaRp6PQlBUo9yFP9inuG92XOQiW
1gxkz32cfaka+htXFVX2kNjPIZsPEzpxmlgwmKJXhBUnMBN2yxDNY5f6OR+w
2RBwRdvQt5WCt6f/smq+Nm3Ik7Fj1ZGqNjcC1qwFsnG4MpR/8MpPrDm2UscI
+4Rc7FafP547W6Ej1IYFgjvO0kLou0gC4INQIaJWGrq8RnJoW+FPTchx2FC9
yUa6JBHyIaXV+NsaC0hFkoNwxGzDG72RLltt30uUfRn/FHeNhb5OOlcujEBK
8j55gMjgVT8x/EmPwHxCmevyiULwwIEzISd3tLHmazfa7iF9FRUpz3RfMg8d
GgsUOkIhZxmK2PeEqfZWDXLrTKdPvu3Yxn4EIpozRJRIO9DUL8ytc517K4qe
o2vfAHHTBOdSbGMlgcCvRsdXB5VmT87kRaDV0s94yTd35xae9cFHY7LQua2H
qN0xksY/lFllGyQML/7UVmFIZ2YwKLCwC+K17dcSYViR9OXecNQ9+5Rh+PZW
+EgoYmSQLlcHrwo0xUK37yf0TPbAQ6K060FB7a9tt6WRtsU6RQfinHfX1oqV
bYlJs6jEYyzNTgCV5cY73b8xx+Y25MuMdLg7y1YGHPEgA7/JYJWnLG/12ZbL
GDxOKvl+od7VqYG7MXBkK6CaYD3SqdpVjbzt8C22/UOhWW4mbdyau6Wz50uS
0nX5p2bOP9AND2/+IeViBvKQZi8Vbisdvww0NZg9Nc7rzGSONHUXhIiZ/0Vm
FwKlTiHcQw3msSv4hIjNlcfiu5yuLDWe8cJXcdIUaH6pBuEfRsFS5OqvBdN7
+P6DkwiMXdqUkkgb8ltPUxWs4WfEXthKteujVnnDu1zOil8XzMrvtbT00j/P
oLDMrBAcbaX/FXSwd/F7t116evXosuzU/UC2+bq/Yf8+p0FkRDfC8eWoQ24p
omcjLFmM9jiSNtnjOcuIHZoRq1la5WO3UvnDXQy1xA1OVuIltc/z7R0XPcSZ
aHyupMguBGgxtPVwZgCKqVeSs18atyMsqslZvj4S6c2P49Yf4gMhIg7j3bbr
qhQh6/WAcPKRvUMU8Dx9olhEoBMgau1gOXDzbk6TgfHR+IJRujNCTrCzHo0U
nzFGIvR+9SduKlP4hBfqH/pbCKgCfNa4T0+uGxpgDTRmc8lqsr7SqoIwkmoH
/Sc+7L25Eo0YcdqUAfSDLg7hyYBOQfsK23Cro71usYGLR3D1x58pMxDYUeoR
pSL/jje1h6Di/XnMRCOswYv4k5UX9txgcYZHHknIw1hirgwzx3kEWocqOlKe
3BWAVTfyQERYypl7PxtchmQUpExRA1p8IJUb+sgB6qcpL+kWpuEt31YQpkPv
WGvd4k7fiIHzuPntnfxc3IkGjD+SIyRV+W8RUPnw+uxvrL7iC9rMjXbPgRuT
aj2O0Ov0VnpELfa4/jcVHzx/4dnn0nh9phEnJ3NYgz2VYVKYSA2JID4KqPDt
ngVy2PI6y6MFLsQSA2cNuSjg1XSatF1h9OrAVqf4UieO6fluY+pQ9g78L0rp
tJxxS3NWV/n3ryyrzlnwOR4undNnOb8xblDBiA/JC3J4YOuwqoR2Z50G+Yls
oK/7+WFb71U5vJIdwp56a1n5Ep+oJba1Wew0KussTu4vb2lJ+ljdcG5dPwZH
HOuJHltGNsW9SM+gcinYHGV1qh84irjwB0uO5cDww5jvckkMbvPY6SU0qzSu
q97MRhxb7N2OjPADwqJE9wbK5lchg6c4qDnnwe3tpwfyCEN+y6NLfWbZjeai
ULM8hTN/1qvUjTINiBHGt2ecXdVDZjalQadB21uTCkuzAORaf4XnFPn0qdM/
sJPDN4Gwmk1GhEaKYsEiTIHL3IaB5qFLsipSN3W6KzdNvVJ3jUGULmfixMU3
/ds9A6r366WpipHQRDFK9TiqrbJkNO7xYw9bCwuTpLmEXCRFy5f3KXOBF9qW
UGCaYbSH/62codjjuCC7Wj5sIVlD9wtBUE5A4+IPli55Gx7/fcOTycTNlOqr
wcmT0IlviJoQxQ/du88GP4wzWskZjt2d1UPnZkg7NWZgGVWomEpNMDCEYkTD
dTbCdjOdjuExp4Su/N9mrltxZAS+L7NBjNSMrZ8ncIusDbCeDa2leynwW+e+
YB63AVbsc5EL8YCu82QH583sjssrNKjZhluIdfwSu+pVD59QFhnQdXCfXMv6
pl0nhxENmGBJqrY3ysfJlWOAN/1gkJkr9ZxUdAYM3/k8vCwa1q+3FgzGtlN2
YcpmGSmC4vrW34jHI6DimLQLhhV0W6Qd6mU+d+UF377j7u+UlJuQ+dJGZ9j/
I6dHWAnLLbMze6peURwQJbQ8iLsUg3SNK/CUrW/ZvMe3sb/oM3aoSV7Qpy54
paaptLGCGKNitYmyI6MFPT+IJzho+2xhf9QQ5ck6rwQtYGqsj2wxw8Y2OvxR
8P7ArvUCDP1K8z/UEHCqceSxYYotD369hvwf2BEAWTRmSflYAQEiIrvHyB00
Lni7vUszZadi4CiY/+r3Ks4zS1gbc3m/6QOvxIoJSqyR3b4kDzNk3K4kdLP3
AVlpCQ24GaF3WTr6C7IBDHPtGVIKhNc/iKrWpIlbabT3QbzFR3JhzhfSS3I8
ZAvzsuIkCV8+/nhcwQtUr+n8omOYS7bgOhbV7i9p1sjcCpCXR1bIM5uCK06c
9/TPiAyJe3t4fQ5rrPkhuQ1Fe7UFj+qcdA0QGleQiFze01elGIHGJKjbAwWo
Q+qSfHNQMecjizN2V6i4iejaul9amk6PdT94waUdqVD04GnnWXPoeo4jvLwf
9jaApcI45LUAydeIdihJzcxPZYcPQhMFmc0MxUQ11XyCWNAFnHmPEIT7E5CX
c3nOFnjRJ4cjIiLQXbnzS332DaUzIeEtWCJzJUxHM+8XqiNtQXci5vTDmwzo
If058AUBg/RSHE0SLfveLtadgmAOTU/isx6Ue+SVmnGulWyI9FvKfvgN+kWU
i1wQzkuf7pZ2O/E7WYBjbHDqHXd0749zlMbomWc+nweq9FjTVt7429qq4K+W
a+Hi9GAUO6k9HYuYCndTv1MwM+4gCjhjQS7wgypipdUBdE1RKPyKcvj724H4
SjWzSA/veQkRxU/bJ6gn8Wr3mJ5UGqumSnSVRtuMvpoEa2ihsqwxr/0BWX5E
zUpqq6KeBUP/JfGb8Pe6DPv4Rz9PJPhCYQ+eEADmoSXoVFKA/iS+0Wk5o3gZ
c06Yq1x+O5BJPLNEAuswSRLXffNX5eJ5kNK5pPnLDkAmn7huFftvAzCblIk9
BUw4bfV0YJ3jiztZmQAAv+xBUsky474QpB1p+Zx0IvFklyRzFrVT67pjoUqb
Js/Ro+zsEPlQfe99Cf8Ivpn2oB0eE4DdjYBer51097Dce1+Ao3eNxcyv2OIy
/FK5HLaa/JhUn4+OYdlYxwGn7vWQdUeznqwSWc3ZTEHpl/FNu2D4RSHzGTj9
p/60vya7EYkxE+YxPB8fK/H9uXN9cgWnD1ueid3ljs1qWi4GuRiw7slBqsL+
rTaSJ2cIF+HIBQpXez8Z5WgHRTkDP/xzhqn24Rf+qUekqzUX99v/aeapwAid
laTK73CE35GHuajkYAzzAdEDuoBHXhDo5VTFGvzpmbxI9ed1DYR2xgJ5KneS
XmUEJCOiWV1KltVsbZc6Jo6G5s51zojmUbrJOFBY9CdxBO2+z9KyY+M8+RUm
Q0zn84kEAyhLE2PIH+GJJVUOwBLBkshiWXbKAXATi1scP3w2q2B6c52p8LP+
JY6hB9Wck62PCRpTCqV/Hg8koZPWJ2LMbBqfjRG7Fi3getTQoSH9sZ7h/bCu
ut7w2tsrqHQMz2nM+2QngPJnoFj63PIsdzY20tKcasOdTuwinY5Kg4kzlzQC
LIQDV4G8cwyDi2iic7MvhSouOaOReob5a5Rg6zt1KTs+b2ubyrqS6cZvUMyQ
jp00Nc5A421Sge15yBeoTQWfSVBU66ePHffsVsYQebht38J90UY/3X8an+gc
L93wkxfUlvMLAIKUOhsZZF80eIw8BGlMFHGin8dxkSkxpyeNmEUAQJZc8Ha5
ADklZPtl6mYkL5xSoyc6lJCb/DszXbd3W0oFlKHUKMKgr/caX73oBpUht5kH
G1mEivDDMW7WvRCv++Vjuv+IMIPeCijCBqf1YgBo2XT2GZTLOYAsFDLx/zHY
IPWuO5gUqO6qXRNA8O98a9SsAZX+Ecv9fvezZ4Nqp2JjcGMT30xE6Bqla+Gw
Nyo7NIECDpke1mnjBWWN5nBwwyBXLLTnkkmvxhqET0tbZrJWI77KUKaV69ZZ
4EWVWqCiHD5j2a51c76AYz0Y4DvjbScOV2pkcx2s70Ey56MUr99vzT3ORqRY
b8Xtg4T8+RAbuZJVuESpLlZ6SBaoKfNXyfhdRhBBlc4UpwunyKIKgnd+EiPJ
Myk9Ehd78B566u02zafo5kUYAwfID5Jur7uoLMvKTCnYgDj6gY4dPG6OAxmn
8R8MOn4N5kIBu8DlNHqxV6ZyD26DmvCiClPuMKHOjqWKAoxlY10JSNcZTf1U
X3W9p0ZPRlyAfEwhAh3r7Lz9wLi7WRKNuGkGBGmORuULmhUZt/bLPoqqhbZa
r2cvgtcCjXJUa0T3mqxCuNHbxkvLyVimBsiR95bT54SA8sk799Oh0KUK5PSx
vnRSQ0m5iLwIM/AdWfnnMaP9CdoxotdM339xuD8wazkUcL0Yqsxcz1w1z6dw
1VEFitGd/bhw+Wf9eJLMQKSGAI9qzG2335T9Fc/L6aPHeX186ZqGt5xH7WEv
hJZ1IvLRt2PBeGGwLFnkAdEkRxThKogOkNcEZZyMw5E422OW3DGUkkpKzxmS
jQ4/CYKED15juMUMide9MU6IBnDnIpw+DU7dY60ERKowYxwnWRAOaIPdlzg1
7rhv7ZtaG+Ox86VUE3o2ZKDDIo//4gptEoqjKlLh/o+gpu04zri8L5BEbJdZ
3s8gEVsoSDJOJ/MkBizgaMkRrPziWlsde+r+H/opOwEk4g4IGqB/X2ARbjIH
8vCXLZPwzos5k8lq7GQrmz2CJbrFMM8lFqMI/ZdQCc2uXII0zkG8Bj8w++Vl
vXHAfTXzXqu2O8KBAz92nCi/pEnl98dkdBdDJ6CVtmV4zsUnpbgTN86AQA7P
1Kg+lgr6ZSrddg8CFsI1ZNl5Dtoo+gNHDfW1qQar/mMZm2dL9f1dGusBlTHc
wYMEZgWCW8oawCzmeUvIzvqJIvJ8rqKgN2hUFoUoxBDj3kRFTJPLE9DL9Agg
ax0qwNSiQkor56VbzHqh2tY2M94zKolmbSl3k24OG7UdOuYpUAA41+ZUca/7
ioBK/9qgqhPTwo5upGGF0IcTYCAwPgMoZb3x69VZ8CsjdV3KZj4TLybuh+lA
nrPFokF/vua/oPez9S+vmtNf2IJUN22bt8oPXw7wnpFBVBKrpDn6kYdmPo6r
vjm6SQUe7/FoEO47Bv4ooOcmQo5fu92dIKrhfmlWT6gPCxeNpjqCFP6QpPes
UCwIHxZGU+BXTh+RgqKMgSuhnsDsZPTvPvE0GxWaSE6fQrNWCBZVfV3F2Gmy
OwWc7ADI0T9WuEwTmvv3EG/yve6O+ykEgM0koeuE0aIhR8YRN1Ys9jBydiLi
T5a8UnG6hKf9UX4dqSC/f4lr9lOpZTTi0bUW44qrmY1o76zDRrKw4YPMd6Eo
zsrn+90DW6+1CRT7HoVS98FNYLI5RXWB4MfnxOn8ZLJhZ9P3MSxmn3lXzkHW
1tYR7vAokX7eaHhbkRjAkntw81pWYbeXZkyFExEXnWmG6zmrHyVvcVHe0thL
nEpcEu2+Gpoo8ypi7B31MJn+CJuxEmyxmYgu82JxZGClP8NKZHIgYURNYorY
3fond8zRcAN41A/eNhgL6YSVp1iUVRXE3bdCvK5Gzppu8O9a7H632cTXfwRS
QcZY1Evhfu4XsxYrYhCWoy1zNoyQDOmOwOgpW5eo6KHxY4rTDqQn1AM23Sfh
EMjYQu75VbXvOoOm94JVjMcnT6LT5ay9ZSM3Rs4ybCuxcKXpglO9G8YPbmTx
mfCazRcJrqtvzZXB81A5gPznmJ/Hxom3vIyTreez84ZRusNN9mMKHAPoW0xO
fNnPMQLbbV4dq9GDXAOK193OyiKPy96bmBi7XkROgJC75X+QHmnR82+YMXk5
Zs8TlvRfU2tHSh4dv2HxDccKqTIMKYOxpmpefheuD9KHwuL0Ec2OP5Y+loHr
56W9F2KjRQMKRRGeG6HyhJR+dqyNTqrPc9pS7GhWmzznwRXSaa9AG5g1R3lc
2A7BFcjIJ0lzzuZVexs3SX74JOUMaewdLwQaNWJ2Y8yiluZVgidb0FiXhWjo
a6RGudG+xTQB+Nyo72Mezox32ggzJsZZPWlB3iwDvFFmjW83Tqld4hrx1I0h
Tqj6AJNJNAj2vipfXfgZwKvDqmt+R+RhYD0Ykj1RcGdtGUXzKXUVE9TZGy5/
+sLsqkB1JrCtYD7+JVn/tAZ9OL9dwtRzJn8KazEKJzP28oUM29BDrDOzX7t6
zq1bkS8JuK+e9m/7ZZ5hae4Sb/EvMhQLJD4t4OCET4TE6c7xupG8Y1PkFq2b
/GQKQ1CP54klQUwk9xzYD0DuRMhRk2lKzuH76Y/JyZYb94FZ1QTx3oP4fFqM
UtA/iVpR7FXsL715Jw3WUU+1Nq3dxfojHqrBJ1QpEhjo/VbusD7CuX3+kc7X
Fl/XA5CDCXOxUcwlmFS3BI+T9w7ln0wWwrmfiHyitZZpbDcqJ0UowDgYT937
hqHMFpc/YyQgxmTtCZaFaVV6l/ncE83HK6T9s8RcpI1d+xzRq2OPpMhvxxU0
Rurg0PkuSM0eEXWOOs5HlGkphfpMAD6BROyX7M5p0asLSGWPdPtdMddtSbRZ
5DkEw5tJJNvloNTfr7aaweKvcmWZ7L2f2pujp6YC8G/ZxXHJeMlYj9kp2ELJ
hEgVZ2OvdCGEoIkSX+/EDlHFt4EKB3vvVLRYpqipwDYATxeSF0tUrqfU9zXq
/Z4nlp39t8vzhAK5p6I1zrBC1UN4qf0qotwCJUNE4POoqaR2ailG+B6THAdK
7/YNKV+x9ito3PGBjJSzFZpEaTaebc0xHl9KZfNJkU9h89JFfbxJDWiLn3/3
kYTWxC96B5xRuFqg4Mlz1SlJe2rTvkO0Xb6me1BGIs03Wi82EQICbIBPjwJZ
dKHoPdmGix8v603uw4kLXwfPrryZ+Wq4ulVzidE1h+NdGufNl9LBHcqm+a0E
U+y/1P1RgfWkjkC1fXFyywuZEmN7IpiRGiLzAr5t4/8AHEwPcBKYHY9pLMTT
3VJM+eiNlVnGEwAxD1tHXpkgiEraFc7YxOMZMzj88BrihJSLn/KsDrG6bWkr
ETsqwVTS8S2DbzEZigZgYbcdA4g8t78mz8qnMS1lnVr0aNmLHNaOOsXSs276
ZFGlqhgXhmQgwPvEzEIa5O5IqMmB+C4IVPdG3x7ahd8/PTODgNgpXTOMOi6s
l9q0HUwI4uxAmPvgqaOrhYpayeHi16sIcJ1oCCqVoZouO3LaHuLjOJ/vMVoy
WTxdsQZ8iDI0naoeWJoVa0QS/PgpbYfLssDobumNuMAKrb9L2mmH2JCg4sEz
pO0Q4L3FRpaU6VWhMZPJSZU8v4V9MlsEcfoNLt6Pv52gY3/fesjVcRFqEfKY
bp5sjHaio1b01kadFePG+IJnue+XdZzhZX07T7sXmJ6xfTGPy8qIIXu+I+XY
OY0XxTheAC2IgqRD4z3spoXTct6BB9mgKGwZF3JSwSimyG/2xAv5IZhiGPPT
MS2yW5bnMajsUnw1yh4IrTmCtOqI5r1G9p9qiBfzMilRtDgRWZzyHwNMzTbb
isIr4VEhph7gvXLgMHWhkKgKeuV0jxcYZgms1PTbawItqhmbfRr+EOul1VjZ
5sq4epPUnOBBnrjfkKHllHHGT8MNONyLyvuUHUzkPkbGbuIDy+i2DQ2b41EU
ydT4CYB/3kxbqGbxdvWsfC6Gm0XtcjLClITkLrPmRyrSksat2Jgi1BYOP467
fnlHlxV0MAHwg/ilfdgrUkPkOvSSkHur3h1lcXZ4IeN8Zac9z2Ubqjph//mY
NjUFXN4m3KDCKvHEzRJ1Urb50AjFoExvMmCjCHCa7y1f53r+GWHlJHdnCCHu
0Zp41el/PBwHcN/x7lG6OdhvZxMIBbjckP3mseWgI49jBTzcCybt+wZdIPbG
X+8tWw1e2ukHIaJrbLLlxQ+zskULQtQRNNHzqnI+u8B/YoZm7qLNsEtUD/im
HLmUC89y5XMh6m4F748pAzTWusZG6U+7vME+Ola3MhSUTWh+HgcZ6/W/oiXs
XTPAa7OANiPe4Ci4AWUZcn2pt122w7erXdAgokHSgqp6AWKWEbt34ozHcyf/
vLTwchah5EmsQlaCzq+iHSgHLpc1uz7xbaQvGw7luF4R7hA6lnIQ7ObmgS86
zSZgr2g8HyFozxlrqfuQvl8LHI9Wd3ZxkD0dv0Kn4Xke3BOqxuPNhinddHed
wtRFxnT6gBd147+HEMtxkOULikEiCsXRK2bEmR/xCx0LUYWOKINgDT/4n9Gy
eQjTGLwoGBPYm5FfPFUL/RDF28jmc2+2A1Hlt8N5pF5MkDMOclUXjgDcRd/A
dMjH9vFMWl3rHMCbsh9lXMdeBoqUlGslmjr/hsjBSeUSNOCcqBScMBSGyW/y
dch/1Lz9qyZ1zFFW1Cxib//4RXgrML0nJwhDMetMy+i/SHxSjIOCGkFipXw9
ndR3GQSaS8LRp6Hi3kuZm1rvKLZHKiacq06dQ/jzquYugpVS6odNMSn9Xr+f
oUT9ACTyXq39rkpJUAedHT66AR2lf1pYhylkxu4h3YHPNMQFs7gZIEPlnzI4
EC3inaKs6W0xznELQnDGSl5b99BnD630TNVO1/2K5bGhS8kLowmuUPHHVumt
XMo3Y+CNsE9o23lbkn399NJIytbHNTu0VVAPZAlKMAObW0elmt4K1M92DpUy
UB0gvjVjJ4SfEZWljp+MOxAK2XoPtP1kU9xiRSHZL7Hm2aAhKzaGf5DShgMO
cIH36eHu0uXHFDXMdHl+H6CfHX5zhRtgEGhqN8PCxLZBZmPYxk++mXXnn99C
6Fi+j7daprlL8RMLXY8fAQBbEd5cnyECmbOSj0kjRIpjEQe6exPLwG07tSOz
Y7MYtBRX/8iSmX9jbTYe3d3Em/Or7OpSAJVhrEiS6DDqNC7AgndQ9b/LgWF4
uoGL7lq0+ao9hzrZlpw0hfU3wOWq9l+4DkzWjXE29a09Q0PuQtX0a4xmxhyK
VS8ky7oWu4NCriR9TDeT1laAj8c89F3PmLsOiemiV8rti1xXdXRh2OQg3tG3
0CA2IzSlRD/XihSkeG17WxeLh5c5v87hPQ363AW9v6S6oZG3V8xE4aEN9MXx
qwuLgtrxu/GdUmkh3XFB1Mysh+e5AAz89irgkCbfpxVZrEr6aG8tbeIGICXo
PCtOZDilOdC530PZ1gECZOqZAy7Xz9LAWkt85u8uIuPnGqorzupTPJr9tjRj
wcMuF8tJcZYH0demRtsg72gZIhDuYjLlmZqh5GMYoPMgYfuOOGc2FjKwWh+C
hBYCbSIVzOcJDkWEXhao5M9eyQIzhpN3OWqaeTEH29bXXMgc6cNm596xc/gL
jQTEvl5fuE+2ZpRbDpHX0b5mm078jv6VYLHlSdkVfo3EHzhjJjGFRZayJXHW
E7azCmFSPchRhP0QlAL9dWHdQ2r5qwraOzmh16KXLkmR5iH+RC6g1S4OCYop
SttLS832vgbeZkKvDeQ8tJVEebOFzuSAXjyuhQzBAOGB9q/+AQ3x7CBEJHXW
BolhH0KFBDCVnhF2C46CtkAEH4xyODdYYs1QrkVvkOjquOumBAIc/6NNRGkM
R+udSGsHnx2MXriWu7AsJRgrmwSm0605lpKTVxpeUU1XrvjGEWORb4Vn8YDx
FzKm8Dfj96pxkCxE8cFi0ZJzzxPlbAuRMTHUWWcS5VcAeV+Pxk6RSfiJa3vC
crRT+IgE1dW3+phr0A0tSPrwtbiFiz5y8EGx7aNh8Nglm9Ey15mT9oAbp4Wy
3DWWHLmhp3G5gE8txyt9to6hiJWYWBZEPDY+Ekh8wTCN7v/peVGMk5pdKkXx
oJDzQzaamMBqebucCGIwbnbYneicH13dveQN5dZBwSF56+GUIwy//bPZe+ED
zWa/V4KzxeQNzCA83XWb2NC3fPw+dQ0KLEkw5ev4mEYvJhwKwUBZwsEW/pJg
SkJdjkrbnrsZcgOeyUYnqahiVEdIJ+jzmRNS03LPzjL6iKbmDU9DQSXcET48
jleZAOt5pwCNoamoivW0og/Em7wEeVpgK4xyyv2U/OwkxkT5azrI8SLaG2yK
nu5G45UwpJze5slkd6k7JtHa5mr8KfiCRtH4tO8ZAk00zA8Pe1QelhLlMXpT
B35jLYuzwGzOAhDTSKkK4Uc7zX8VQiZ0f1GqqV/6RuRVNleJPlXBihjSP/fu
yvKP6Vceq4A5C47l8tNIVyJxB1BtJRUwb6cyNepzGM7d6qA3kqXLm4d3r8ug
AHBCEL1T5h9zmthEDDioxVwoU40+Vwg3A5XQPVG5oofAn4kKSu29ODFk1Qyb
DXEmiSbRzSQExgE7yL9h+h8roST4diDfW1XrrAhqcXkCm9Q1C8VlrmwkwMYA
NDIgjGDVMgiIRyQoCUoR3TtLl+L9PKw6VXDq7szqXeJ2J+gqiYfc5pkbnafS
fqqXA+vpQWdJu4mBfJi84+KgGB6HulX26UkOCaN+o6REWNUWHBTdkLZP/qG6
+/b3LdBjrC3mMOMsduVRaNhdz1tNsrp6DqueLDGb9gAXHvLMouf5ER/ju7a8
RdhjN2pBidzUKtcqtDbxzqHZ6H4lXITQme40f3zkXYiqTzXj1/P9NMU5yMrQ
buDY9U2v1kTWWyTSDOCpoc/R1oXPFEr2kkKnzwaq/Yrs7380upsendTK+2Z0
xtO9AtaY7dWd/kBcrcM5BpPL/jL22o3kJ0ADVeJUFv7cRhzHgKJUMjPOD+Hr
r96hk36GHsEdoCd6y7IojugUt+Fnfo2rrU1v4BzKC4+RGAxRGVuBXv43PIwO
Q6Qahcg89LcLAS7VG2nHUlAttbqwgVNiw7exlXOrIYvLSpdmlErXe0sqD+pI
LDjIWwmn36hLcpIaIMDOmWxPw77uWTfpHzgmHt5HYIZ0teN8ZR7PwsoTvbEp
3gMImvk9RIJ1QzlPZ4Dcz/w14mR1je2aIStz3ctvsCLe0CEQazsDfha1T7iA
hqxp4nzll2O0bLLskY0r4l//PVyGnw92fA2CMAwG6R9SQqXZ5NhVsSQaUe69
W4jYJHdmDfZQGWGMBTbXVCrCvJx8dZ5XblLrr/WhzF/5m1H8UPEYIXmoLIeD
JzT42AfkXsbWULdU/mSMdNfYYigHc1qQ/nrbVBI5NQsMhAp1pQSbHhpcQiln
Ugccm432OG+oZpTmI6yn6Do04SGOYo9+TggLuT+RSNMRLkVixgTwe74rxcn0
8N87YPeWYPxng9fpNY5ZGRW4+3I2TGejdNnAd2FKRgTIr1+gmzXBoOJjliIA
5hdqlWoHcKfihwBLWHTRfsso9HDpD+l1P54Sg+AGySQEFKi1Ayj1nZVSEBhj
yQPS8micYtXkqu3N7ZZXhrdRsd7w1Ldsj04WyNXPWO9CsQDYgkaikVKttbJA
e8fBIZRnL/evRFUnqiXPNDxoTc5eV1dad6QuLNYijPObFhOSrhAkeWYbYiYz
it1QnvaZFCWoOt6cOkaOUFIOAJpS0XjipZS0ssaJboDYNErYuEnW1vpcY4Z+
0d34zy2QY5T3f1ee0GjRHoxlH7m98UcP70hw8qztBOEs8HM5J7rBB05IEdTS
nnQbrxa3rBks5XlwMeVz/hqZma/tSgEvsTFmXrOtDAg0Foxnz4UmJ9sZiEOr
MQ7BtU2/+pWBZbi1y5hw+YtuRq9FbIv69FN6+jAPE1H0agFfkAjMpvVJXS2p
09aPDS54x6ngDpzbE6pPh3Oqu246glD175W3EMsi82fLBQx8WXaouFsLUYTJ
kKfJj2fy9uxrBDy71+piqILt1EDfw/Ok4vXhjGkN+/3uf/rLNR/2ecc/7FCB
m3Mc4S6Jq+0BFKb1EcYHw7rMQqaK4oqk7PCLkO3FrzraQ5XBAsM3Aqs72EqH
VKhCSz4cQ/kkfq1hZHJSCOkpGZl7E9RGZigPooD7wOwD1lqyYo6cKw5ME/ho
nSHRDEt4yeN8UVkqT0USyV1rJY09a+0UESLFGiTrvvQCFjmdeBJh36P6cGkJ
HtmCSmaZEQ56tBvhseEI8xzYkVPKMN7HcQeao6NDfq/AHcyiTEuA97N8/Lyf
Mw7eVkbkX3LH9RHm2fo4X5XvBCKt7Et4BGnBeCbJOL5Hm3T0NVYzQxTNy+p+
QTXI+UuPX0xjvrTqyWvnsKJ8TUNOTTPi9T4N2TkgZnOLQPLddhRIeKKqyoun
tzlgHQDKpAwZm+yy3TpL3ye2YZBMiYLP6iP7ITu1TMeMwx8MRkNa7LbqPpWh
J4UZ07JuBLcK7MzmD4qBQxhLNf0O6kR2JFx41nj+9fKTAw7uaxR9hBzWxr0I
8fVHgwFmW1whlyUZIWUxajnWep50xyxcwDCYWFUTp6pScT0jGokmhdrgIeqS
mMMqYIq0x9k42u8/P0wAjYj2E3lqP9ZMdv1wMeX2+NNrB2aAvojzjFZ3FuS3
5FDehfkoid9Cek6vS3Gif5kNoEysmKz0U8nOjUgqekTaZr3CLk8Z/7/LMs6B
bQyyta/T3dMSwiif9SjlVi2jdpFFW4zIAbwqSM0RlZ4cnTh4holyE6nE9/0r
ovBIP1vf1t89O42S17HAn4hYP8tD0BQ44PB5D45WA/YWmwD0JfNjko6jm5nT
qm5yLyV6/cUgstNgzQcX7LqskrKqTNw4T/hJpRM8IWVr8MMERV29Qct/8TDQ
Vmg82iqdznO8hlvLWqMLbB0skk2cNZiXap7RSPfzQ6Pz2jz5adXesyC1OOd1
EQeUnr0rD28DyPYuSKvzk0szPXnx5o6hFquKh7qwPx59YFDn+LjRlewT/ez0
MkK+040pdR4U6+nkyEEFgiq5J1cS5fqXahGofYETAdn0+5m1jbEaxsUT832v
iVecpjG9dXnOsvGql3NhBP/IP19ndUW42hIu4tFd8zl9f3pyTtbegdGKZzAm
N0tOTYSfJ7UWGHq4o8J8HeuGnMlKD5gi3+Ep39NbMZ+gErO4nI+ZgrmOy7Yf
o+qUaPr1qPzOGRr945uTyx6XuGzVA7PoBE+udaur1EiQmpX9A3DEtXH3Qb9d
M5glfBnYykU1xOtDd3Bv9PJ/FeEkskCwPfERIqLgwEgO86zmJFdPBV9a2EcQ
R4HSMx+D1I4hX3OKKAb01v66as8q/dD4/FlOubzHID+k253bAzZGZrM/4Cgy
7iDFnAR6h/lBjvMgjx5I2tzmIZfjMi86+ATV5wPVeE9kHuJTvMYHn/BKQJCN
8jS7nb8wjy0ION3vHFDZpFleTXzD2EsxXdrJS3LViqVqz1Q5lwm/e85JYA/n
luLNKH9BJSgnteyQZs/LVfAN/0kK5XzfJHrBJQ9p280aPZgb3ikuNvGRF+Zy
StH+43F/ZRUijNXxvQ0elKKIKo9V2veB8Bkj/wYWh79S/f7X9eFWCTxEXe+b
1uqOKfJZ1czX71+bb3qDhzbv7nV58rfAmgYeb7P805vftJ0y2Omr1XYb+ugj
gLCytTbS0iGx/suNjSCvxOxKL0fLn7mERmpRFOgBYH/OAa5ukYqDj7Kp2eRB
6GdIBUFBAq/JjiW503tOssvYd8zWodY67r6P+S+uNt9G9vWV2Gc41XGltY8U
Y0k4yWQN8uuLj+JRzpcUpQPFDZpLszxjcmxGVLh6iFx7VwRYjG0rIWpE2guI
L8jYS4VEanit+vT4OHMti4g+RUpcQrjopnm3ZXhiXev1IAnHEemQ9+nPS41d
uUl10aGvvG/uH0AYx5MbG6ePngF3XYUelQgV4a8mBh2QJAh61Jib4jwGk+Im
aG8GctTl0OkMkJ55qWDijVXWLu4Sv6WeuNDmB83pBP+8hyKWRGz3mvF4vVNd
mAeSPcA/Uky8MHivk7eZ3W1a9gCtRiKOfp4Svey8J4IaHkrZ6qQLsC0x9TFM
GNkfNNCzcOJdbELi/VqSA0UjxwFSqcN9mKAUSS593aJD7Z13huDmyeyRdinV
pPYr1gI4YFsKW8gQYR9QsCmOvTAi9MWSL/V9+zDPOigP8ZUR+cSCvYjlQw7g
7NXXY74+A342ChhnY0VTQa+3byUlM8AJQhkPM1ODlOKGULs7GVQe60T52GFo
SzNSm0olNfm5GuGWJfnZc2vspQeVbGx8IZ7zk3WtlP1CyRFnIyUrt59tFxQp
eKwawzo0Z8Ww8oWiHO/CXb6hx6dpB8a7YOt7SFbSpOEug4MafmlxnadLsjHG
241SOkJ4RrkamolTiQkY4dhHcGpBHyDlsGLmPSkaVnQULmIe9yN9r2VwYBuP
OGYwSkQsj2ZKuLJXtibJF0un1SRhpJCPaIzn4wW19lhLCmjy4TpimmyuCZxr
Ndb3oMxLHnzq/FUO5XMvtJVt1DEBxyYC2ySGfI0oSWhRgx8EvP32WSSo5Nz0
iJplJV66eFi03iU4LAXxbX9zntITMgPoLAXq1JshSfa3R4K2TAQrISZ29NZG
Zp8cqXdOj0J95/I2q3s11Ma9QKWzlo3d4dA4Jw6fHuWUySy5ToiPWAYRTyTE
a6gywmaQAe0ux+MXMCBeI6oUwe6AtVXKF/Poj2DKaXCQuUlkJtMsCJiufkCP
75GbBHkPlM5e4yZWmNBR/JnOyLM4+ZT/nKWnPeiKa08/D6ntVU6w705A6bd/
2NJpfNaCIirItQqwuPftb8SSM283aLszLU3LDnSLwZ0yaB/tNx/Zb+acsmcu
DGU7grCDyJMEnqgVRwSPkFYY1NPlykXl4MW1FLpxp+w9oHUuYEieY7TcBS6y
gi5pQMC4GXhy/rF+B8TZjt4KKJIH/wP7yyvaJ4H2BpubXG7ZwctrYZnr4TPO
NZBDXgRVzP0dcZ31xskbV8gsVbSECfmWpx27+I/K+K1b7Dkuvjdthqv59TqP
ti4P5UEZL8nn/DlQkZUlCGb7oMbP1Y4lip+bWgiIYbEL+7TyWPP5muRImYui
jbo3BkHP9g5eHgICiLO5Ai4ewOKSaDSLhOVWpx2IS2gZwdSedxQ0TtAKrFn4
y5IptMz6HFA0mTmPXZMfGE0CzYWcno13E8k7FtFJzhu1vYKx56zDFDT76bOS
Ht70ivTWbcKWCYoXsyxAQxnV7STskuA6kiznR/J5Ner0hMUx8qystfaDIYoR
+I+X97d/W7JowlUUiS4VNWU/nZUXxFHSkjAnewWqj2NNQHYLU2tjG5xG6CQ3
8NzEr/RzNU0RvEwk2FXgLyn2l8LvFkzt1ZKRmWsbhuMrBVnhiTMRAGB5/qXk
4fDF1PqWFkD8seGzLn6ibev1oGLyXtKg7pyum36PsAlO3eH6otJbmTcjNtFf
6Hrbr7Tp0NjqvWmH7VSvCSzsZY5PyXDkQ0lz5xrNm9AZdURWDQXjJX3g7rPA
kUQE5srbmiE0zijh60PflrgMdHGfpo2wfo7kzgcWoRc4DGrKDZB5BjqxLkPW
x4p8dMVBR+DWRwFIHks4UU8EWb4MNtHQ5fU095eahWLek0lUeVjZRBxiiK44
itnEWdtqmkG6DhdIYg+qRABNfvIHEMkDU+ypdfmsfpS/u1/PDzL9OPWdC5IP
cuuQwU9c1AdNcukyVPwBATH9nF9Cs6nEhYQZMSjEnEK+fbCWY3EpgpMCWimi
VPi06gM8YvPE8cnQHmqk7kBikN0LwsaSgMG/Pm9Lt/let4vQjRNJ2Sgc9+Nd
wUoD0SYY7JPdsB8wt7zBNsJz/KF3TAw7u7RYxk4CXN2l7kNUXv2JRs/Yhlcu
yil0c1kZIE8Z2avrj2P/W7pZiFlMmF0ICc+WlxXvzLGgP89M8FV+nfCr90ME
ECTQAE9IpHlyHRf9rbn6Z4uYvlrDFBlkRBeM3FD5i8Qo4iGY7Ho0+BhXqE5N
Hy7Ew3hS/oX58o5T35qb9cUWFzoDn1Jq+OTP8ubcMvjjqYOCKj5DqK6tWHSL
ZkBSzVH0oKfvoc0+wmYuVRBzu5e4+TRezVliH6kL2vM3I6TqdRHHpHKL/kkG
llMubvUJq5rgSTWpX3mB94oGcveQr8WcIL1Kb9z9qiUUAt6yxSLBdj3FMqpn
NWCO7GVgvc/F1T01H8eCKvKdWsp3BK2saIbPASZLc7Do/xJ7A1og/aGcXRqw
xTg+S6EagIHtuRDg+E5VNvtr53KejUU3OQ+56vhaBELl69h3Ah5MieGkcK+6
5vylQwPKyZCfd2V+I76xrmFlr9Ih6JJi+oBDjl92NNA8o1gVbQEGVyfQeVf8
UTuoZtHhEU6i//jwyxEHr7+yOLovzARbBR96ep77+lUm//ja3yoIXWutRLrY
8xRIN/bfbZZ96VLJk2oigPrHVUFTq0+jNvrGf2ZA3y1gDQO7CtDHpniEY8XM
CLn4iMtThOIaDB8VBBb2q1vFYvMJdKI9UfjCBvQlzwHBcaaOR8hAtwEcqMr8
ieZ8VspVLiPQmZ/pk9wlOnEfUtY5z15LM00+K9Y1jQgIaDDKAUOMeL72dz1Q
0YN7B7LlTyqBRkN8Nj5wqDsW0NoQ245rv/OpUyXTj5BE32b0JFO0xjyfewRH
Om0TXXWPIhVwtXLSqWgmnSU642+aACeti6ez2rOv5DUTZ6r5ugm+jrKWCdKA
yIMWFWhrYSppPM5nsLcWJiZFBbH1cLbx62WuvJIxl+rjIjd5eLTYB8gE07K5
oincb7EISD75E7a9Y/9Yl915igAflbTcX6rGc6hVDbx5fx5ER1dtZ4UBYDee
/ewlAqv7e5KueIwNTtdHDVOFaIeLVv7hpmSQBM0MhWf9a3Re40YK4osZxZkk
YsZbHP1rDWBgl0P+P9rQoPVDVIBDKkZq1jFyQbRWYLpMwhaEhelQmJQkCEuQ
g9SXwQiekzKT+yNX7HcT2+3Q/YgrQ1AHMNVIdDzdG9/m0rkA3cyj463lcnhF
nNTb6seoCip7LgbMv3xpdaA3shblami/26yVP6AeDogT29LuWE7TrWzCoV3v
iLgXfaD8IC95Ey0Sa0B37QdeoPW6AjjjJtBTJF2M4R+Cj8gMhwwWTWZZ/cxB
kfwZjh/OyiiIRCYLOXZJXdqd77Zu1VmeJR4hgJglcMV1vyRequOee/b/kEGR
jp0z5alYqBTu3qclSlRW3VxRmzLyErD9BDN0tmJxWhM3iXgcx8ZvtTHMT7Rw
0bamqW5LI9bGE3zrh+SWQoW3L91CRksITDIwm0FovzMy27LsRGl0lztMCwJU
37WM1TLhjFRt1nRpnnQUEPMXKMhdLP/yVUGRlk+U5QLCWmXArLJICTMz3WHZ
SICN9uCRelW/GWhKW3i8lrAcu8+UrQwvJDgKaZbK6PYdViEBHReWcyhzoXgp
NOKKegbYvPBzw5CzXYfd5fJ5ID74c0SKbxQCRYFczfrFTwvayxVCkj+6za89
+IxvcQ0US2UlREixmOxXG04JXKd7sMqOdFh1pCBeIRwnZkxmU0bn9dwrl1aB
ulc7bzz0Pv9vUdspaIsapmb0aF5s8H42d2ebA4vbJnPRWbBc2C+T4FTKAd7k
PfiYWXEtSck8PjXUrWMm5Whd6+2Eb6VP8F/9OiI8GQvy6LI+Jvn3cJ6VBabW
lqd1FuJxjtECwzinlADm+jHrIyp0OrTf35qMQNfqW+mbx3YMULOOZN5jEN8R
ZXa8QuUBVlAeAcnMiNLqltCoc3mUZyShhyUKpRx2wZ0JLuwMLSdxA4tVl7B2
auwCTvvuApjIxvdva37Q57xqb1uEThLuamMA4RDwOs9jHuds8JQT77Zit/d0
bCVzIVId6WZP6ykZmKvga+UJFGIDO+wYP2+fZtz7T4OGsJjga6Ldc+byMdC7
6GXn+3DzuQ9Q5Z+r5QDG7XUKp3+A2Xdr7WsE5UF9EBOp47uXpk/6WxQbJ8Kc
aMqdRMoVcSfPt4SLEcSzOP7WmsQqk74/yd5Xu3TLP2jlDMomLT41Og/WewIV
6hOxitePmgzEiQm0MUbLNU3ocOZl9WgRq0MDEAgiUu8QhZEx8HR5wFiXVYfK
qeETdLTOYaYQvzJxsOfR48TYDW/95A27U6ftG8yvDR8wAXs+9vkvSQhK+n4M
3Y56wA7N1GdcR6CcfgR8nr46amP2JsL26Stupi4jYVlqDrpImXlmMD1W6iKL
9YDJQdD+dITgh4yOwy/8wdAppJG0qStD5YTqM8PR3ob+UDqMVs+wWtg/e9ul
uX2gw6uhdebweHAXK1kvhU1UA1RLPGa1hIYPsq3XrlS2a6C02ZwfreyhFuY3
fPakS5VYjPOLkFr/wutTJH6YeAfzn/gQYVvOBnXOCZdu5KaXgpql5sAjfiSB
da8DXQc+DskFLoJySlZmaFJfi8vEUXXzF6kWWvkTjj3WyD+KTdxD3kpYt+6d
lIx1k99Zs43eafQD4sJkwNtnmi3yugQxIAdhYS0uwhcoCsnGNrccU9uwX/QH
S5c/is9o0mJ5h+VjBAMEDkAnpZoRZ4V2uUEZsviP5K9wyc+MeLGv1yhg3Tc5
DH8n/uZKnPhyBq/8atNrp93qzX4a1s9fyrlk8jmfcWkZqMyxIXhiBjckRwQG
Uemb5X82cVUhaNt0CZapTEN4UW+768rdUp91psSX4kv4kL1uNWErwlMlU64H
spRdaA74giKFjvA8bNRXaoAXiElb25r3LHbOxmd8mBGmo3udh8cpuoAH1fTO
bZbfrTZX/XJoVZzpJ9jVNJiXA/Rvuw0UklKp7mZLIeBXp1hqk4A+XRbmKUOg
vt1pBdEBD5Kg1jozJnHtPNweSr9g/JqJxEGoiUctQevwyiC5csDddogdOlEv
vmjZp+AVDTzmTjH0FKgIrjq3ZBdTHAPM4GTUYRXAf2HuEwg/SiesQ8FqTmLG
hY/txGguTfNqcL0uEVWkFoJ0g45rVkk5u+f99RzR2dCP3tUdWLT9r1U2e4IV
c8Kpz9hVjuQ82TGMmE13oQL18KG9kxhUDnqmFiQWgo7029PdKb02FWJTj1Wr
YdzYdJFDyGnETGA6A17fqWB3uuNWFRE2EnDTfe+CHBqIdpl0yAUMdFgfwQPU
blDqV/7F/03wqOsxL5CZfHJknz1MkAYngnryBZIWEZ/Wdx+uVwWmAMzftKTQ
VgDO6y2RQ4t7RpvoiNM+VyLYT28OW9S+yZFFsRDrO9YwDSo9JEEjE5aelyja
0RvD81c10MCgAoJ8M966fLu2q5+rrKiAXrL1Erkya8g9Eaqi2PwWDI1fOQi5
OueV7yeFrICbTsj/lGT0uaXRa0rtEmqqGdzgm+TQxu/SO6ZXR/OMlX0Cshka
Zl07LRwj7mrx8f6uK/2Piz9i+JT9M9U1XMolyGKWz6J0y/Ie3YcssZiD54Vn
pAVvK0MStgES94jbh2UkGmYtaUxQJ+r5DeSjbx8BGeeC20vMiOnS2Vhr0vWK
t3JJPfyXUlumKLcfGnbYTDMO3Dnuw9PXxkD7ksynn0lIjsAf8L95z9FY5x5+
BTEQp2CBxZLN25tN3REYZ6mzXvK1B/Fk9B3B1orBCQaldNQNoLvV6xBxWMh4
xS16CpWlU5LEPllZAW8hl79YVqYcBiZV3gs8mYAU8BBqjX+rIbcXUO1XPLLx
JwiYLRTV5jE6JPfCrRoQkd7hTzPpjiCjXE/k4AZTJ8QDRV2prYM3HXyeTW4A
capqYIKZKFdIj/bRp+rFNFtKuSHQmqhZzri+MNs7QJvGNUTLhId/KrCSQXN9
QOlC3NePZF0RIMTnYHzg++koEAmMsPhw+jIVvyxyY8uvfDPxknZZzTJ36Mmf
6P4AbPge4Jq777GI6Fm9A9UbkPl4F5amy9CBVr185oB5CMLD+iGQ1lag7E8A
oBuBkzUEqKfJUR2fqKp+9FyIHsODX/Rg8/JiCbH0GOjoy2zHZEI9tlzNZ4ha
orezY05Azb+8UqqcNnDaJK1/L2W+yw9dspuC56Z3DSwG+SfMiYMLhhgrL41m
iU3o40ZXq5UrdRad77OvTnz+T9vF7LrP/G+0N5V9d5hkAvxiWAWP/nKyUQOr
vGmDCsADzr8Rl7K9eeIy/nmtOEOLM7GMUj4hI+K+Q1lVC5cUGCKxWaHXsP17
bbwslj3u1XvA7ZZzxJeBrcn03xZdPCY2PrAWYi21b8uqDgOT5nsg0UdR9hli
8lH+heVDry7OyY9NxYJpAmCqt5Ixbyy53A2lJoIxVT1WM9n4G+Qm4r49xpUw
UAbFuZTJJK+hGyqH73PA+dm+jD0ZVBONfT5PF1drdJ7rgD2ocmcv5D7oi+oj
xd6Ubj0e5bByOl/8+1oiwUG3ROna13NEsq9x15dSrSeHvL/VELevtvBUcw3U
4xWAnmasVxkAGrEO5WqkS32rq+8pTUPtj+NcO6AT81rUlXXnEE9hJfgSLjc0
g3E7BxNxT8LrzGaAxtR5bjki0caD8lxHG+W9PegyjxL0q1zfh1iA+HF9Jehd
W5fcr/e2W0yCXNK5sCgXGaTIlL2FjxUe8q0BDnRegzvHhXk5eG/Qryvro47C
yWJpJokiZnwiEraX13aSoh/fw5998iQGx/o4E+6vsLf9crelrOchpnWcq3Zx
hnAMuXsPmTN1lBvnObU+/Zy66yAdCIsAyJhwp97AELhuRWvhyCSU3/7iBshJ
wtg/RTKtDtpLYpQ9aMl2kvqwHOvTqW/yTJRDA1n8aGtYUqj1dzhRuIdQ35MO
RNgYNzazlGRW0Ib8zsGZ4/qqXkVu1bSWKwNTF13capozenQmRd/O6unde98b
s+DMvAtCRg+FYFpvgZ8qzc83XSFne47aclXKoVflLqM6G81Jsd+XFqGI6V6W
LdSFAlctmonjZ/w1XUX5qZrk1v3113BH3VjkRnL1HIcYExsyl8t00a6bDH66
wP1EHFx6b2ROB6hriY6zYSM3wjnfTtFVDYc/Cd0HXXR9FmGvrzQGUBkNlUNj
s/cHgbroSQkJ5fKpRNBc24CjNyUfavH846gUzsoTSEwlKIObdSzhDIqtuweg
SqLaB/0jUr+VU1DdArkmtg0st8+nwyaMXfNcv+Wd0pOQsylZu1WOjXAg3teQ
hWvlITxU6vvufukQ0pOlj4soNV8BZ3pZ9v98CXKVCJOU5c1+jdcYNKiLfZt5
NlnIIwoQmR/LAgHJQAUJvVMcDgs16tDC7CmXjeDMCFYK8DsNvFleIN2H/rw/
1F4AcPuifBl0pSJICt+gee+1r9QxiGKrJBBSyxyTwv1gTmUS4//r72i22CHq
XkxW9Qh2Uj239Fj9e2ttzsTJ8bpBfMTf7B1/wr7yMIN0jTSjHGz73t3IgexI
Du5CIwnRj6IlvmI9Dr660qpoBcdvfCUYYOwHPvqWhe1L+cTwUgeh4zlph5Lv
taUbJi6x3aTrCvazwDOVprluvJV3FoX291tUUouf0Egn2Qewur+aY9JhTX1G
mQockPkG1EqtvblqL7x3jtoErMb1RzX3P84VqncW6ybW7OjfQxNHQXfojxws
m1LBn1v5lHT4j0qXOAdH8jWeA9zq3vN/+B1SiV8wTbZa+4R76cp7uAhJ7isa
2mMkuAxsd9MUz0USWsK3eOuyKxXGM5wfSOevi0fYj7AzQPhe1fSzfXDKxUKU
N+Gv3sDh0iSeatWKhh724dLkva/LC7HzeBumdcFYALOGEfwiuWZK9ZqqXbB0
sHSwNyMlN5iq9RyH6wiM8lXGvu4073qxWD3GbmeKE4qZqF4dyLpkPaCvn3rY
62tRrHsAxhw9n/d4eRYgw1N6WhT199tl19YY1iR4xkmhNnYUZcQ/GeULiiLC
Nqea0GiDoQ+IKAQM/WHSHo5FEXdpi5fq4Xk0lBnb8i5GAx3daraK/kuQanz5
+1g92Cmx+oOE7Q0Fu4l1MgagsMe1cBWq3UfWS6WOpc4OxOxGYYrVnnBVSxer
2oNQk3ukm7FET+B/l3hgc6Z07akohQ8GdsL+fp33QO/wZm9MbFW+ulHZiPk2
g8/qOg4z1cGV1YCZWcKwtvpOryaHEO3WNeTxC6InxT122nQcsgfSpL1rnQT7
5JdeBVFwUXEdX4Hya91i5lqRs2HZOxeJVqVqXSgRtIil1GsemADewB6phcQw
cURqcqQcOxsTe80BFnUlXfqoZGecGxUBG6EzedJThEOxzEJ16duNpW8NvUEi
Pm9tr6o1n/+ggZQiTYDGrUxbJ/q/53sawXepWdeFExAIhWn9kK36ZyAO5qMJ
IiLhAIIgZ2LqJZkpwHYCr1B5ieF8J1lZXxDqrPNmkDC7dXu2FtxdkJsH0D0R
EwlMPt1OE/mk8RhHneOv/sAh/9wz5Gt5a97yhs2T4KD+KWbyFiT61PfeRFK7
JdsMNQT2/HZgde9Xpggo7QHc1PqJ+vkv6vMVsmu2PI20z7bMXKuRS8opbkXJ
nGpzL/mCsS+JaSeINkLwgwVW4IjREKQS7h/up9D+Gzl3qb9pvjwR+8Ox5J2a
Ast5zhT2PLNena0wive2sJDKpAhK2cowSUJPwyY6a+cLh0Wu8HrpcRTCosWO
jf4CNscphsqqK+K+5XPHg3ItXCWNH41kx1pHepMdxVKwUCulqrJXAnwNRQ0f
s1bh+p/6YuQZCnSlbpN2PvHn0AT+W1RrAHg/02M8chHZas3OCiM1DFP0VqPt
Gi2R1QHIxWEI26Lm6frGfw+vrTEpRu4z205WxPvjmWV4jq9UjMcu/4q/LXZl
TT8zBfTJvNWcj1eHIaxl5RKgj7iaN+Ngrfekr16XH3A1n9OhLUvRxMHJtTOE
EQjb5qTRwSSN+miFYW/ZMrmK4jE1pqScJQ7Yj9AxTCIjUEibWs36vWItqUve
bTGjnWCaXGiodah/ou5wYRGZawLZWFWdd13/WtLCpnK5xDro/hr5L9+GY9iF
9H7bK9iYEm+mqwXz1Fq+N8UdManQM29GlafZFBhyMB8t9J7+dxfxSDaXL/tB
PG73BOPOiAx/aubh8Z2ykulccPkxZbTK1eLCXlKWd2fAAuuc7FWUVTRBU8l/
XhXJD+kQcP4f8JGBF21FrJ98iEIVYmvjQm6R1SA+sakhOVJuYTEp6AK9wrqZ
vYYgW/NdAZvGGX+Vk1BZFGoUSFgJ4YkwL/rbJdeQ6kSsS6c8sxzLBesHGShB
w8DU9xb8iBj3eQ0+g7E7wm1mKCvJvvGExot71XMUbpcJCi6V4FS4CEAz7ue6
F+MzMyUkahb2/Z4IAg2mDb0BIz581g+5IKEsf2OwGoMKwJvPwuJN8hf8TXDg
yfyZe/ONV4piiTTRVktKH1kmn6zgaZ0f11twv9aVm7luuIp4K88xcGCxrunK
p5Z8z6zpJMUgdQYnCv1pFBBdgts35bvP0loBdGQ5M1js+kBNgEV3wfWkx1Hs
yWj8VMfzT6lX/tbGuOB5TMugFg7zfWOeV+L+fRymnBlG6W32JHyh72y4byUD
tQkgelLW/z2Fzcp95V8YYbgYalUKt0GDZiVG6OlD08KWjox60BDNxQhfi7GK
7pqN80AxY4Ky+hMnGhQGuKeUEoVyyhOvoNMrUkuyR208tmzGPMgE8rVEYFlM
eaNjQoL/dufLYCFbO8deflaMKcbBGs7WJxBa0bw9ti1/dOqE8RLrg4gGPho9
TnDcPM6W9oecslS2EzF/Fe/8NKRcAcVj5ctaECcMbT97+Kwavuv/47Ej28fJ
3Y3G3W1GO28bdquDVUoSBf9CgLr6Up3vERntKgMoa/pGXY+cRPhmklQnq4Is
huVhpn3HIsJtjpo1T3HVYVIUMO85Um8KmWwlGdi+ZvL5iBKjTXXhQFklAMsf
Cu5Zpk1UxJc9jXocbyv/yvh2hEdCAGOG6vxZUUtoMwJ15rjyNozU9acW5pS1
hmSsSciNfG+R+29dXNtE16S9fQAWylBAatIzqc6booowSATM6AleGlXpyXvp
ENIC55ifTlpLvQVSHZ6BbTHu88BpIYfQZ5gPe+T2CIsiUtzmTk5TEBPo8MiX
nT5eul+6Jp9w65TR5ax+OuMkP7kgHo8K15HeZz1JL3LqwUtKeUC5i2A7PzHc
tyIF6GWQmam/8WPbfch2Qv+Gj8qe2RdZ7SRgRTY/O1fdpI5xilKYgmPUu57d
OZeLp6hoZIHw2lS8sZO7lDzasHNKLZ0YEfet3SboNI9Db6K9i2BvOr9tQ1o3
KEfncJM6mj6qZDGkG6fvQiWrJTMGz0rCruGhzzgdUh6TlWUs3IVY/E4X6wup
w3oigp2/PuiMVTBJwj6a84AxJ3jhnO/WeTI/FIBaVbj9T8x57WnsJldHhbvN
XX4QjT0adfX+5DUDEZlNrUjVYHTqNWE0nuKgsV/90ms/FKccst8a2yyNVuq7
FE8eSJt3p5Nm1G5p3CjKHBvVN9kccqPQSJ/+wpsRy/700NfcX4NfXE2nGP6Z
40fMYCVK7QQqyzW6t4ehCmhjOCu3VJnBLEsruERC9jE480HWMLR8SkGgsbzo
3mBXNVFUopW08moKtLIJWVCbKxIBkxNON+BRujpP9piwSM3K0OHulWd3G+FJ
maxkY0JI1hzgcvydLBL1Y+j99PrEnSWwjCc1Ou1t/WwlcLejBWqSBtOx9q11
x8omwmGicVYBzN04mOUxyspx5i9sNznF8iDXN2U7FiAb4N7Sgs2fLqUIYccC
3DoYL/W2l5ZW4er5GfWtTDviMjPr+dCzw94SnMzLidzoSRvrBD1lv2cskxdl
KgmbtPitdfxVz6Z97PMlfAVcwM5/14+A7zv7/77/VzEuIx8IZygXhfSGAgck
oXuqgJACf8n/qm5n1TtnLG0pNB7+D8E+YA3liNKnvA1t8g8ckj4UysGUZ6Gn
masfV8R+x1r4AI/9pepAy0AeGBO3D31U1U/Rc7D7MlWKAzsp1VUXE5DcsLkF
8oelAPY+eq6VK6Ey9yQeTz10FKaKqdpFM8kaCQy0GDEormyfKvL8ahtmS+wM
MzmVP5Wy7KbFoMUoRWVQtKPJgwt/A0Z0TWn96PSA+cJKe+zZVN4MlEqzk8EO
UkEDyjtcRvEXv6cWLl6cJ+hpZm7oYzCOK681CgXJOj0oaFGND4UH5i1tBjNC
KSoRo60cTbAwEy1zHgNqC0UwNe2L9scal8m6Lb0W4l7vaJ3QVkf+YE47iP30
fM26xsU+lOoLNk+At0R76XgepFVkzCVAChIokG+VC69BgvcajYLmeJ9Bg2zI
EAwKDI6KLGng+lWBVxOifF96i5zSBTKLxbKoTsRut+St8g62W82A0JGCmm2B
tty4FWz+bsN12a4/CQcFIIkPg3Csh1Srxu9ebRgf1iHGEjjxsfxAdgl1l6Fc
kwsYoTlS6U+jvogEugXs/CSmf7WKgfWWi4iI3V2M8tkILO761Gnsvi1ozRiz
KzEzXCBZvZ8nEEiRd1qnTgiXeULiUs5q0JfiAwXOmDVYCIPoLQxpfPR7rVeD
N2prBvVkLwZ54wvfwUU7pU+2BijDcSpcbmeRpLfE5KDwNvNhnKj6xzA3Ksi7
guo1ies08w1/h738ENaXwAEiUk4Aga2DEo4kpCR3C69L/ThsuzS/aRf9h54d
+IGSBCLhUBiIs8Y3tmtu1k4QKYK+5gmfJBaVjBWuYrA+ar3q1hJqqoMJ6I15
q9Z1mlnPY0kJkAMg33zbxCsWwhD96bHly51ZIKub4jSXye+RUJYrLzdgTM+J
Ft0XoYW60xHAWA6TjjkA2LqjPxM3ff7m6OTauWEaaW5XWcNTly72mW/04/pD
nUW2oBU68hvW+mI5H/sEtZ1+i2+w5OlZMgpepowd4JuU9qfI3mTbL35HeaEp
6XcbLIRDwZg9mkVTpktj4c1+oVUZ7U52OeQyMCqMsdsMB6EofjmjtFgubtYg
PHk7+olHoiXgNRSgbsaxJWup9tcr7sdaMJcdX1XbXVO2GfGeciwsZPP86sJ+
EFRbXA0r60ANVRc5jKhyaYOsgS8rOEoYiWS6tTFuZQvds5EAJ4q3dUmVsU6F
SND5TusGKA+J2xNoTnJhaToGchT9dSd3AO3IvCpHYuXaAWbnD+68t8Qvq/FI
iiyhDLuizU2+TK4ZQiDbXRMNXA3E3Pa92JP1LuJTZToMyCPZO5dh162nKRAU
Rmm/jlOpskuYkg5dWpv2CrqvWyEKywgeHQescRM9sCOQPmk+ckomY0J+sA74
bJPz6H84K+GBW5DvPfbch34nN7Fe4BxhgdH76GsrLIu4eNDIzhnzGYsBXOEL
wJR0Hj1R1o17QkDfJaNUxtg8jwoj66ztweSiuT9xz/8yRcO9pi/b0Ev1/5vJ
U7ostl2ibTf8dsE8hAfPGj8ou2Oxm6B8tJCuPVDGG4p4ZwvSqwBeVkEp/JrM
dvDH0v9lgx9CUdAyeAaoGvHVQ9VMoSzZEeg7U+gNf/a8NPn3grR0BkBE2i5h
0fbgDJOqRwU8AAaRd6hy4/MxwoJ/6P4bOYv0XgLi6Pru30Wm9t7Ne7cEGj1T
OX7Y1Hfc/xq1Bv1bsYDZq3hj8eLht/RnK6pee72FtaisR+mmaIksoC5Bi3hW
m7CjbvSQ7BMxDctUgAQleistB80nqONLs8x2DTavDQkolK5IlitHBkR43DwB
U2lsuKlevrSQbx0tLCLh5uckxHACPsmFTjWeRcO2S4AOWahzxLjucuJ39leT
jrS6OsgkStOXwyr8UUFOe/Y8buvGnffG2H3DZwQgUzgf4B5DKOdTadFuIuUA
UERtxbzzJA6eEaFRlGExMSlsnf3FAbq9DGVSk4FBZ3V2UlvLLKEJYjsZ3OqZ
qtZIMs8xrNfoodEUC3B/5vWH1PQWd+yKvoXziqByHvpB+LLk3067rCMS9WpR
Hs260xpSwiOupord2XtL7/ZjRdHk7aavLeA4t6h2lZO7GNbz7tEV8U1POyq6
irXBYd2sMUk8Hudnz4epH0r4TFQFnYoT09qvdFbMd5T9o3oFn6CfmvX62dzs
4iY8JVErbydLTGpuI9njYNn01gQGK6o8OOegYuhalYHUiuDvI6LP0Ra+NFdR
O2Pj3frRgXj+ZhHNWgHfhH2sBle+VovOTjbqB5+5/X+Iq09M1N+pBrNejY3C
lBW9DRsHJ75n4kmENcXSsKe3WPa1gTYTrlLqb61RgfjevyWYiOpJWU+A9kdJ
m8GBNjIAJH/q5tHFkY0BLyhEpEF6g0hqscntpp7FmStXZEfvr9AIlyZjbYnS
wAV4GJ5zy7NLK+OqEapL9Mf2IWDgMuBUBxfwwpt7frDIJ73pSPjp9eAqkKXF
StSOLdBUgpCAqUdHQQ9FeEgWTPUl9lVepeYQeun/sz2hKNLLssHUTQP2fmrJ
gusofPh/w5CIWuGtHIXdDO2uh8ZJO77+mzmoiCye6BD+Wtd+zweNmpTIMHH2
8vHgJKcuwD0sCUugn/7RUhteOBh8HcEQjHfaMUccneIB9Exu7aTND3ukdSlM
K33iaTTiFuYSXEPLCGHRbNKO+AGrDGG8SQzQ6z0rhzfnIK2yk08e5xmj+0ZC
IvYxAkP1fZsLiLppeOr2cC2QJXihNuO/V0IwW1d3ZpNh25xcH/tFGXEb8+AB
tZSlKDWYGkI0INW3sck9fLUlBFUybt0b54Nl1EjlukEKITCloamin/sO4dKl
dx5XEKgDJEB04Xn2uQqb6ymh9IlJaQR/VmDP0q36Iqm/Ro0L3YCyFdiKZLwQ
DrXsOsDFOmK3Hd6Ydvlxj6zOcgyqI1DyaizKLiFeXAhTlFy2HtvthQeA1nK4
Poua3dW2Z1GMYX2WgQf1S9PV1P7UCb75bjaDSSoXQnal8SU6CCcXT4yewsje
WYl78j/8/R2wAWuK8K6rnsxkx/z0Nn9s0THfHDHsZerzSCkcW05tvWVghUht
10+xEKFCpafwnq74qTNkk1pW201nVhn/ZXtEsKim6VVd8rHU+3MGnu9lG9Ja
b1RpZwdrp+5fL5hYQLLeFr/IUnih+qDBU3eqHwLIkvlAPl4ncXBgGqjRMjad
/XKRjnt4Vo0o0gF0yV2xzG1R2ZEyuomUQkCUiX3RbGLTZ9thpS1YrMPbDj48
b6ybNYSMzLBmEExHdkDV3HZ4FMwyUO5BqIXD7Cc51b5S4RqYTZeUfBdrODRt
FeO8qi3qFrMJcx0Q05IVDVjfoggFy1qTfBk+6fdL1cchUmewcjfBxGfTCvHp
H3c9uQC7QoSkkgds4nLJGsFx6E+Z8BCOstqbSSAhP2MxABDySXLJjku4CCds
H/OsaJBh1tOuYnHnUoF9e7U2fIWQBDTWyq2J7cvhnDgdtQ0u0+SpAeLOYJ9u
JtJ8h0m4FLhe6YeZE9PcP2qqDrZGb5A4tc+ZGu8urPvdsBhYlXRgpaO70lTg
wyx3HvM9YUkfWrEKIWnWZONSmEprhBJiO8k8UcpoYViq22zCR/9glRDFZJYe
e6bADM8TQcWyTStrSXGYyGw+VoZp744u1lJmiUs5xxuC/k0KvxHyivqq41bv
nvKinSSW3TSH4vRlEr7jdbmisBQ5e68YDS5V82SlA2ZqEbNw7hJazKo69mNT
XaGGSvvQSKS/iPdbIceWCU3hBQIzovM0WfjE3orgoOnltpL/mCZiEbC8FYoB
Hc21tDAleFWQ3gPyAgxWJN3L+M7EG/QNJy/qEtaOiOcIj3PFtgIrhhyDCxAN
1esa32qgehuAZ8T8tKMOF5qyQPA002iFO8cvt+m5YsLaSLkVlcWHqxLkKFFe
McietbRc/2u2uWqf/e/Zam5UCCGubSjY/vNMBDjJ9Dy8ll/lGGIiGxFTEA48
L1Vmw7inIQw6zjEt45kbp3XAJqCWODUE3nNVklMo7tByqjn1wZMs3ubR71yY
ht2XDvPcQOWlMUA70taawqAA22XiYb5XdehLnqW3mVrKOxMfIyWepgx0i4IS
GQe6tCM9Fd4Qm5BdEIhNgQpT3ehdeBflqAoQENmvAIsUfK8YqnYxh8IRxZuR
wbkSqfYdrx/EgeVUNguWlX++4oqQY4FNUPYWIgRAbEVU8sWkXf0Tw4T+MSuR
QySfZJBZGs054FbaBJUMTon/DoUGlX8JtUe2QDjgj1j/u9p8WZFDOHDrmpda
HqdL9vEmS/T/IIIrRr3pdLFKn2rz+jAhmI5Qh9E/8HIqqgjIE49ncrq4wV+F
Xh5dlh/3QVm4AXIC+BKfuBQ24TIwVJPQE84T3nC2Mx6dwqrLKGpCv4R5fHrj
bRxnRufXEAIdMkcak8ZFycDZVIJSWFTfPgP8yfXbwhcJ8oGyLSRKy3wtYYc8
QDJlIIurQYBtnRxjq+QmrArOFeDmeX5CpWRe4kFCIGoHu6PS+tjW5xhTX/e+
z+/A/E3j95G5U8N1aDUxDZBWHA7IOn9QCMKNwJ+V3a4yJXXv69isZYLBoCyq
YALyOMkD5Xsc8tnPTSx9/9i71y4UAdT0DHQp20pH86nmupTALHNIEuV8xWBq
tZ6T/Vi2GOiIFe6Rau+idlEXyYh5g6FqsXE7zmc8eKU7l8BOtvqt7iq9XM0v
i37H6R766CS7Hqk0zURJI4cm1RM1aGv3r9KbIsHg5UTR8nkOy5TIBgeuhGxo
D6KbTnhxvu8jMUyDnAUvjy/saBKaRSvoup0JcBFkhFzh4hE5TmmibxnEeAFl
3AWWAJ1wADYpvFRaUAzHDj9w3KiThQozNtun254BSZG+qMQK72ZLzQ/pzUI+
gFbIqeN0zhhoHPYs1KY6WMvFbw57F4h9QMvpKFAKmpfIiZIsxN0Sgo9knbh5
FRdHxf1LWv3EhlGanEVXjIDaCEdiNchozpqOPX12clNu3hmQ4mDqB9LEI1bT
s7PhUsSxyMjVrrhP4AM3/nz3ETo3ZteFF/h5F4nKaVr8VYI1JHZuvtrN1L6L
cC8nhQ+Vnhnn5H9uo6A5PFT/MQfH4shdV3lDDyhzbIyZpuF9VKjZeXkkSzxx
X4f5vYYfDBnBpw+J3ATLsJFj/NnzLrAGNffn0bQ+bYaU+pxJeouy0kdraBIf
v7o5EhrKXd7ZASjSyZSaJfgZwfyErOeGjERFSfxjVFIkCu0x0UIs7Fu1fsL/
4Tc5zB/vQyo0p/YtfOu+INPaXK1SeB67mHiesC/qDe0luMO98XnCHkVGBq6c
mIgF5NdpthYlXpXmHHicaODs2EHFnm9hGYX4xrYcx5Rp2iGPIvkK5jj04hYJ
SZ+Lyg/xG4KKlQ0kS/9ztMVFHSF8/cjAj3D1TYijf2+vp8PB4e2Yw6TLyRwo
MFWC7i5Uw14yiuiiJI41wWW0EB883tzGMfCRfUm7lDxO0suR4A2zPFGONdVb
NfRhB+4QmLtwRKzrr60RvWTFgv6ypKNTyvrccvU/88ris/9UI5cSu8nWfdtz
oEy0WYJwdGH4KQuEPrLYXalSSvbW/Z+JqI2koLYd5ipG8rcq/Ec6/R6iH19w
hR15sIhGsqIyw52yPnse2N9gt9kc2asf7NamGEqO3JwIpJDH4tBxziEw7Uft
VSS4dHPwduynNNMXWB0snmTElpLHiYL9wI+Lc1azuX86SGH/7eZubM8JoiNJ
uRL83vjELC2z6cME75+Abhtk9nT5AtcufpNWY0k4nFt9wbCb9Vssut+QieEs
u6Ix9+6SqMXRy5Tj/VoALt1CmD+APrNvLQdZ6krZl1DuAybHlsLy2eRVH3wO
OjnfOWKHkMEFuqXqT5cTw5gR/m2mdeiLw32dfbv7yB0JHkBKGFweny3fy6TC
/JxHG8lupb7I1FE0RbY1H3WiOnhtmMoieq/W8LheKz2yu/lxQF5cT+otqBLR
noQSm78IYjYiv5DBK5r55G78onch8Zn1dWt+qURoNCqMGHXYG7EnHGrwF3gs
PkxEVppicQbVv0DWK56wmQrqbNuS60xOfnsTMZCL853fwGDrid4NmIJMFTk3
WiKxeEbqaDG24BrEyBRzOmqJmQM5up8bo+eJZJuTv5BTeLDGabjv7UNxdrVT
5qks7RieOEfVHQDQP7zPzPpITWcre6ihUaMP7XrzkZjQCDBbGq/04aCByKqv
pvNWejFzry3tDpjZYeACq9R9z5z5qyPnRXQZhaH/8H7VNFXwJ2TFRJDCnlo7
I3Mk2/rp04K7a1xPgftH2eAxUbQ+YVUu4OY6JPDnam4wxTHb0T0GNfcg0I4/
Z2tny7pSMpjff84LK2o2NGJP0DM1Z/dLh1Hk7I3ghRjaGM0QzME01pEHnGP7
IcGU9hJBW8D8gS998+jBH7iA08qoZmblUBSrX/7/g3SeiuqwxuW2oVisPdIG
wlzrVIxjNSX/nSn6b8qY/urIB4ubxn9E9sofNafcsVst3yCiuN/Wr9ZKo6K1
QJOuVi7AKSsNlle0Drgf5fRg4v2PWPrGbwmv7rSdEg3WfiW/6bo28SWrOylQ
LThd8Zier9XnFqrY5lkvfp+i+K32OJRR5hdIGZxkGZT7ZQgxhpzeF5AvtGAM
NtP04exrobQiJMbJZ2q/nTnTdzKhCK4ttX3b49yWndq7u6uMsxOwPMGARJET
vVXO93zqFtzslGWQGLZuNyZ4fdtWFAQjJSyib1wRoT/mzLvV5H3kpzGURxK6
4G++oyx1W83ztHVWvcm29rg11yJBzcn1sXbTzp0yl0h8JFl69HR1JX+2Q+GY
4PiqlvCmRnarW9ZnY9+PWFYGOUROXpUs8UzTCwJh1zSi72KmtlVuQQcCNz3p
QG4jwytPLRRgA4ES5cDHN6fWQ3yUt5ArUGwtrEsiv8CN9j6bFyyuc/COiElf
oXmpZWQKyhzzfwPbAwtlCuG+7GfZV84GMiOBiDA2GaGOjzQcUuSS+QTg7Trx
2itDTKt0TKm7YOmi3ZW0wFUWoqTcW3vNZCfCiv/GI76EYe6BkwAFs6ySSK4X
Jr9MDzzvJb9ZkpEODDGrAJpeVdkDhvR0YhNGpn0jUSJm2tL8Ztfi7kfOf6OJ
+O/fX0cRU1O6fVBQP+aoVWqDmXRssVwLEzbl1Dx6mWXk9tg5Tj8BmXXRz3v1
+RTkGYMVJF7AzvhhYQVMNmvGhhTYhZ7tjXI2BmIf17p1YEO1bwFt/dXFsYB1
neYeouYl4uq0FvuVsAmItp4XDfcVcXjEVSJE8ScA1woWcG/ed9HrKm/5CNLf
zFQOdZDZYCiDirsclkVKoGOZnpaNERsebASRsFasTTifaksF49IVJyHoj5XY
Qm/Qm9LPqzHdoKazGTpXlybo/f3nleHfDiwimIkjtJxmPPDb4g77ZsYT6uCc
OUA5B3DOzd5tpyOrouGP5IgqPovY+TH9aYctcXpZO3ZhoTGftrvB2LSgG/3J
b4e1pLFesVPirWfWtqKMeLzJOwQhifTHPm+KMUnGI+/Q+xQcIzNDerNCwm40
v2MUxjdQs7dWcrUNs8uUik1HwUKfgR3J7r85bpn2oNbY4kBGXLS22nSud14B
1xlOiZrMzU6RjDkbJNOjauZWJVsExEOExcobyKq7yD5FKpi6VPoPKfnhn5sC
V3MwD5NaoC5Fqg9v1QDGImX41/pa9XW+z9XW6hyvSarg8ZgvPlTl+4hJz8/B
Xvz/mNvs5A9eVAUK5svqK4D2EaFj+j4OAduRcYQaPsOcI7DCTt4XKk2fo6pC
znKzfUp9K539Y9O8lYG7eo5QkshuFcWbCQevcv6F9TO3om+i3IlR95o/Z6dO
unEm0gZTkNRd9mNk4DSzhXahUwHY+Cka/MYe+lN8VVOIOmebNBGQB6m0Pd0Q
s2uVfVjQGWz2Vyy4yJxK6HG57aqs2125ExETpNYJce93tP0vGjzHuFq429/E
ZVQsESP9pztvXtuTpibZ2VoB6tBWLiEaB8hK5El4E6NLN9G+pCy5HkLF9AiN
t/S+Q3SHtaxANtI65cHSp+Kji1vDOmlfX1ZOKV7W2O9/FxZ5Rq2NVSaB5YnE
XtRof+OUcRtTB7xdyzE+XvEznqiJ0J36P0ct3TrHNcpsYXwQO8y+i6cW888d
VWGZt4R2n/EEO0hbN8TL5zh06rG3UQJ74c/V51HflZBqFWyEofRhSfcKsW6f
dJkQyM5ZUiO+4+Yr3kdq+NJjVKQqDLEC9vXoqoVuwqR7qfmoMGyY+R9rqLlM
2iggFT0eXcjUdEEHKjci5BdWju9Wm+g0vgC+TAsGnL4kp/rGUh3loqpKUayl
/t2WW3mVbH7AX3fIjKioPb2BXMpNf6qCHYVverOSCSiQgW6RJlHKKO+kug9b
cAKcAoW93DmljceM6q8r6A1rqb39MOkLyq27iYxhpDjMF/SjuJI7c8boNPhb
I3FzYTYpyjYheiac5JCUtSU/0Tbe62mRN8imd/+KMJ1fzvmrJ+r2qtWMH07p
4clXONw6SQD5hiIlGPGO5UQuEeoaNviS+D9he3drHQPgyo4IgsSo1K5S9psi
TOprKWmKCGywHOQhpKhyi78XyAoYTB+7A29zb5Egbc/A2QoBWcCNT2ktblrf
66AM5cbwgqd5IMvkbf/ZnkOLzludbffup8sJc0tfDum3QQ80GxMAVJBmxH+/
4rMhdbVc5WtMrfvojHafJYNyPRxpAbXDIdq6HpWNpZCRYGAwuDOEWBpv/nwU
0vfHqP3Z87JiwKjeU5NLQcDHZm6w29LQD9x9wOjusLztnBF4bpGJUJMUI3Ws
RTwAC05AyvE3Bs8qZh0fOEgq3RP0iInKRg7SjpXNQDnJMyvIXas7XyDoKOp2
cGF1bMeR5QMk7AJ47pOi6TB9s0i+zLMTEvad4jUiBW6KBQ3M5TUnDEkL6rDQ
gwThGocUNvq5R/oW/AYkh5jjG1yoQeW/L61XgzQI6VXsT2zwjTGOtAm/RJ+t
xIp7Sq4PxrC/mTtzQNzt7YecVyrkeDD3KqMbjT7aIrNobQ5lwIoWQCJpk3QT
/a/X1lbtYhCOM/wuutcyXL+NrlQsHoRyOWmUiR7YiabbYxyfklCzMfn01zmQ
YxObf2dXioL5izSh5p1U9ZsK5JIBeQsBwC4Z8HdtE4ut2B+ta0mkdWVqHBG7
71RQikSOUGRai74Nnjq6QH6tS0BwgNAbshjN7NxEFEBfqnRLqD8M3WOAxM2l
hYxv6iRRf4n7hUDjEwqLQl6eJSerlCi9bA0YOnFKVH+Iu0Bj5f4k7tr4n/qb
tFBse2BaxDlCa1mi5lAUfijaC/2fpNG0/NPc+d9A/s337iJAOQUcwHDZvq2b
4CzW2Enb9CGSW1oChsCJ7igKEfLXgF6/nFs1H/xY4swnPGPhlLbjmrOz2GGn
MKJAmqwJ3XRZ35tndTMOq0q/tT3jE5XLoKbLFgWzqcbSRwF1tnnQYb6grT5f
o2ip5qd6lerZl7QRkNiieShXE060nau2vmXQpOGUaM+mbZynkP7eu2umTcW1
2WgIqp6nUfyBfouvKI/sj27eNz3eJIHdLcRQlL9LpW6gkdAFHmehsJAnK3BJ
QiTBwWYqatvODYLoUxTRZwLvK9Vqepg2ZhAqBzdMRbR+tEp5sDb/TaeXxflE
jxVbp42bw2cL5z53HxURHZdPi1Z7BoPPHB44UCFZeQUHp+TK1ZI4OmdDOrGO
X32pVlbh1BMREa7x3CVOL0mVPVIuQ2C7dftgTLOyDngoojrbNiKuFqJ16sCX
k9yp17R9vd7b2XM6bbRhQ0MHIbBudtl+1s5RSV7tXY2u0oXPD9CQcKQV6M3l
nhsdbq7pxWdS29vWi6OUrhEtbAA/MzIGF4Q31+jcHYA+di+ZKWsr8PtsuXHk
B6KmAcHsO28Fqa7RHyXAD5hsQBeig40Cs/1yFb2HdDWdwmEG7L+NcHRyFWpW
UWscTNIt426Mxr5wrmb9jzoUibNZAUX66MWru9ar12fPd7XudnTgD1tnYsoj
ovdHSBh5gokc4eAWtMISB7uqZQyCZY2FMwlh9fha0EoOtxepFdSh9h8iIMvx
ocptLX6cLr84r+8ueiKA7dn4dZ36lGYM55+mS2W7292OIBULi8cFf2JHjbv8
6kGSTuw2196m25Zwx6iVz+Zj6nsRaRqkP6hmQFE+moryi9j9F0ZS/kwD0oyJ
Ww85bK41hi+yCckOGcYM/N8erEEB7LeMiG1pQH5/LzEEZBL5gnm7k8Yp1tm3
6ekisDabpp59PguqX6tFPOQNu5K4R4VgDBbQoyaKVBZggjy/+NMiN3NCYQ4A
xakXmBOXx3QPUHXw5qVKjkO4EHC0reVwEaG8Tip6iNidVJNlsk/AlnsYmjPf
Rxt/P3GLn2A4zfGp2cXPTH+NPSGW1WPopWR9Sj3+GGFs+BIb6Bq19sLlGHoN
z6cbcczfF2ORoIb9RsckwI9CMyKUT8E//awQNoIJ2RvV3X2XAJE/vipByBw6
3ZW8QC6CpLS7yDeeb1Bxi/kWFglT1S2l+CtfbxGKdQYeYGG53+5q1i1HLu0X
q9zDKHdK5Po8F9aP7sd7cK0cC3A5U7d1XDr21myiw7OYwd+D6wGa+ggS+HYe
D/bMzOcXU6DRBQT1qO6L6Uc/ockzbr5KKVzQ3EgckT5arvhU4sDJWds8Zuyj
EqD6D34M5jNsqAvNV9gIjTE8I+9FQSx/ih/tRLn1Iz7Vc4a13rdPcu20UCU9
SQ2x3kA33xcS0vkWdMB+KxYSydv0x699dE0ytRMbDZPt3EKgp4oJL+z2eKtr
mX/027uCmWZXG33+DNjd5Bb+1zyQkCFYS83Ums3hvOKchXtCr7DP9uOCteA6
S9aw/kGX1O3Oig+n1SZlzCs/NE4hw5ODxEGNBKA2p+ZvucuZKlSlp8zedOcT
nm5FYTuFFF+/PwDOQc3onNc5snLNZoRWpbovOv05n1T89ESwZCBFPaXyBp9W
/mcZ3H7Hr1aMwi7whHzPnW1IeYi6iYauIN1hO/kA1PDR/l2AZWo4/o1mMPcY
otroN3rEjr4tCHdeI55ZDp4mBxfPb/tYDXEajE6/Vx0vQtD1/MexBtWY0ts1
I+sLxTp9lM1aGg2bFb/wHR9vsCF5a+UeNWdAj3Ky9Id00awi2Pp0q8UgwO53
hQI7DB81D+EY091qSPX/16uJys834tAZNBTP7b19MVLy6RNS703ctadI97wh
Iy9JYPox7Zd6C7noePLGd0HH8ZQpoCm+qrNnHTHMXqxkDtMAC9BuN001+Xjz
B5pZ8QuXwCFj6kn0vu9EBsamPNYsR4hYsjzckoV+NQxMC1hVZrETdYj3DaPN
Y3Aa3RvHVLdOEWmR8huepIuD/kB3aq3G0z/x2gLzWkuuETguDQCZAifnsSJd
BaV3ullRMsv86lHi6yrqzOHhQ+4UzSkqWcgFrCF5FbbTrH61BBdIyD2LEG2i
00RNlTJIdP1hFgUmBhV1F0/wPNyz7ypmUOvaogTLknrlI/8hB4MCvkLWaK8o
R6XB9+Wt9haG+RXUrZn3ijajDEx+i9SR66onmHo3hOZ9++LdNB35A5Y1tvLK
HPo0UcfU78zX1xXVcU6esPYwVGxQBhNFnK74hOtM6kqYOvxi6hKuk1i4QkIQ
hAlgQeIbSW2j98+Rkijp+DgJ3sMeaUyaUO6d9FUdkSeOvYHp/2nnjxgQTjB3
LwxDMeCPfAbBBFjrA4+7m1sla9lgHrIImINCOM0U5otO8purSyLYmEaAbz/P
9bt+XY8qVnNr6MKmURujQjjjN8vfh8atWhzs3B4RDK/2q/7NnOGcegi9YlfM
47yeS+Ug2gAxLygX91Knj1XSK/Z79TCU8WNVHEF+Aey1a3C99WT+DaTUtNsq
u1PreDRf2RK/vn1dbAIPqugIC+6Ig9xjBm100tCFP3CqBm5dlvSrssbqWK89
P8UQd5DjC0AvgK5wQ58lCU7p5RFPknNpiWtk2UyHfHVgSObmCLN5FbiNxWk6
PAgsgjSL6180uUPH2I8qurErK7cHzz8362xfFMvMbHG8x5AarkDOcfkFwlRT
hyRIrRX5QrX6t78YfCO+Jqol3DLuDMsitMmZ8j4EDQGzbPWej0CuWBfpDhSr
lhyfmcF6Ovb7J9n7j1jBQ1fdUoS/JXu0WE/1z8mB9l6bRB+wQEa2UvQKpiVK
bbqsTBgzjocsfQgyofFT43pmMfpaYiizDgJtGEH/qglYuQ45jvpA/FztWSSa
yWlRZNqx+T82rLpZ/j5vZyPALWpaxbGKdrILFHoYClIwkPhFVsa4I3kfHWcj
4sBVwWPfwjIzAoKrWcBeKAfa4CGAFzybjSukAz4QU18Mo2eR7S6N8g+ncr+d
/eitlyYST9HkC8HNl2J6KYLg+cUTqHjunBEckljWhZsjNql6XxSCkjiNqdS3
2HcfLvw28bELO13qsvxC1H58ymVPhslgxKLOjKbbz44A/jBE+oekQX69ReFv
bNf0Btyd691SyL5eJO93ZbKd2JZYfkTqPBqh20XcykQ49XPFrZYfK+j+vfUI
3uydukWcKKP9o215hJXoIgUz1tTBIHPB6C8+WBiQXLIghTsWrAqKl0gdhqK4
wPUFTEoPuSQfaisjzaoEwpHcHglr0aeJPN0BVCbIhhWv733Oe2ZbYQ9SZkSk
xeoxHUE7uaPc3cE6hFv3Vr82KtAW+/Ez3k9M0QnEHdH61XdIlCa7ShTg89q1
gc9jtTUjUSKuKpxgTWyvVnpXVnSWJrpf80xV77wv9hoXZlco24NA2GDp7DPG
1Y3WsDqQQ7+wGy8Vt9glLgAJMnFDegnh0S3PRNspU1vDJSodeMwV3iGuCuWc
kBJxuvYTfaZK7QljYfeqqrlixKdMnIMKljbntOlvCdT3B3DsafMKgQeqvye1
gLH3t2mT99dLy9zXtTtrjJPAk6PhmgnjHjbGprukXTZwFkIA70BzTViQJ9GB
qS/Ik/KdkM3rNah0Tz67e02aHWvM240sk1SOQSGIOCvR9HMTffkAZFxG3VBW
vckq43jaxoQ93MiGoeWZ6TwzldLPn5GYywiZk4xp1wKjLFkiaN1/puHQwHnx
5TFWg+nQSDNT/fimADFk80Mws8OxkcaTHvuAvIPHrahANqDx3PnWSyfZG0UV
3dzgc48EVyJkhCZ3ztafCf/G9uNsNvqDSKlhehIEAUMLsKd81YHH/TvyFLwk
YMbASO1lEHS8JcUUdXA40khxUE9/y5mEJO6eid0PbxmonztdGkJDM1xtRNLz
AlEyZC8wXKT6uzLHqjFp2FoxmaFPmnL0eHm3zr/pq4jyIHAABqbOocZuZF2/
hcve0YfYClu81MUQQP/JpoBotP0D7EvqqUW58jSbPaJnlQt1fKZT9yKOkXXS
BPIu7tE931oGjXfIt9SAS1d+efbIXqn6zF6hF5bZWqkwEVrVNAgt/SpZrF4X
ZY+eJISQ5FcrLc90a/p6SajxxPHwCPjmZQv0uYI15PHwJcDRhJ78TNd8F4K6
cquAc1HWlXMZVZTvHQPxXre359MfL20EomeN2Au41xhqn9GxG3ts9o/bUC//
kM4D1xfnbqwguc8aB5T7eSfjDrXbFrel7JEu0gYLOsWhg2mNvsAjRSbd0UlW
b9R3RHsaXlw1FOstqNW7hS77m8HhiNRI889/UmM0Z7SwqiOFVwU/ThFdsYgv
JMqsDZH1QcsaRSdmjCBO+q8D3zixdYTFWarIH0a0XVsLbHvkhFA8Dq306zoY
QrGdacgcSoHK9Eb5rTCOGAgZI8nYz4fHyK8Ik8iXu1uoXzhgAKnS/1NvTm6S
05keREEKomUKAIwCcbY2b2C0X9xkU5gjQLQJM2niJtfpWqzOm3UdfYSmaaJ6
+0v1G3vA7RB0fQjxjPVUDPY8vtieK52ja173FI8zfKk+QUjMrJfOdSKFoEBs
vMtbc91dBOnx9/UfgLRGxEMnGPRExqmW6ihcpcXcC95CLLEQIsIEukAYothY
SzlpqHcZDkjvXHB7+AGaUvAxPiLbELZoSxAgAnFPY8SAZaJod/8MbV6OVjh9
dOOgLZjihbFk42btAjdN4wv1lZQjUDwVH36sh4sUfoZOCzpRpGo7Ltmo6QoU
HBRpF5D4BznuyWYYfvD70ajh7oUy/GjCNz/uas1TVlFnEePKUCgMCJw1xne0
vNxf/Gy6KnWbWwNJ3eH3/9Q5bYf2NC/H1ERufXUFTng7EN+pXoDi1LP2AyDK
A7ygCNTtoLkXggso6GFmKwDQPJbfOd+CQrrLSMWR/2S32swJ/zxw8TmbW6VO
SqGUV3BGE4RsoksTiSE1a8ek9UNwF4Dpab+Pic0oWH9LVpiLtkSWv3cNl4RM
KX5Cesv78qg9wr+yaa+LRmvvr9B0uzi4qWkMf2qwdtdvoafU5fzZEfQXOq5S
WB3UfdtDa7iQfwqi0pZRHDvBsE+SswFWiaB5Lv+ImGr/VVO3IUacqcN9Sq9C
jrtHGct9bC7diPptwLcrx+BX6lgn2uuMKZL5T1Bo5Zw6Hf7GKpQEdAn+ySNu
rGhp9rLK0Q5NH0pmhyrV5xV5zRdFyw1QG+fJFR4+oBNjPmjA73yhCQvWNV6J
lsbRcq0v1nG7xZFelQzc7iCbIgaxF3t0r1wdt7wu2l/Edz3UkQ+WYL9q3XQq
2Aa9hn4TwfLWG9C174hl/cWrQjpm7alP2yCkdCP1GZ0og1SroPHiKAKJIjVQ
NKw/DE9bqiD4AhL0qg2xSW9JRw6yQhkhVj1zQG/7leWMqh6gij3/zduyArZl
AfrzefUwwIlpArVNfiPoveVDvPga7mIevanK8ROOOOKxrKZ7yTAJrCV5/9zl
VvP6rB/0Q0ZV9Q4rPQYb1Eiv+C87YftS8M8GvaozVCd1ploc+W8/WOfCyf7K
zlg2IviPxBY8I7kdkRTQr4AlvozyN887KJeY1LjRWiUnaoofXK6QsYZUHOch
JOJcLBJmSteM++S4oufKcTwKs13J6AG9GiU3i7BaD1ryVbAGZbc1WOKguL/G
8fLUbbpMZHwAIC8M7IYpg3hXcChFXc/2ea/Oz2Evrl0HntKs5DtIf77695a3
6Dzj5+mQTOAuV2ItgkgjfgLrxgquDEtM3Rxl5qGjLDX4OFadmaAwTFjt06Vs
4LckvMhrr6u5x/OTNumr4W4vME+RX8ck47d5I6XjtJb8K5SldUA07IUk1kTR
8mEFRoxBLrE/PRvmre6rWvpoZ8Eq21IRvplc0ji9bhMW3RvylHAUD5okyDwU
InHdau3KjKTUg/ca9x77lPeTAIZDvp41fFI52vZe7/VS3yx9orgUAOQPHU2D
8Tk2TA8CejsysrBLeyqGzCPgSoi+6ylsO8Eg2GqqDyBTdU25UVxmzkoO4evJ
vmAFXvHcMCGMbEt25IiW+O2CW6cnilfj1FXRnqRSmPvPVbCpPYMlOK1jvIcO
PlbW4oXHH9rGZVoeBTa6SxkJmJYBNxIclMz36cbA7Sm3nkMpm9F+X/VzdjcE
oASkq8pjk6Pa2j42FQTDcBVjZ22/7ZnHMEFEH8pjTWllbh9oVhSP4Zuj2PaY
cPCkqQNX98vv3Y7VOzSz9jbcPCq5KJQPRnlox3gKYJ7v6qW1k88+mSE7Z5Q9
qepreOP2SwGwLzR5NU/zf+pJi7GVK/g4M6lr6wkkaFevrAPZQayTJBHwWhY7
INBXwJJPvFItns5EBpa27qK/t/t3iBHAcSFctoe1QXIStbOg2N1Xj8++Lg37
Up0o/Pp9aNRYeoXQUyClgStcIdeDWpM4r8X+yVKZLmsvDx7Rk6EOEyWFWGWL
cVTFEZNdsRIMkTF+huE/dNE5DBulTpdw7YiRmmgiKuz0WMyiOyDB+HPaoXSq
MV6kMnPHsXQzh+WkMWnlZV88Tm99aYs5neBHVBFp6v2Er9BL2imhqgBnvZBX
0BqoPzJ9zZ0Rf774wu7FOt5InpsiJ3ZCR7BMx1oBexyduW7dE+jJODdL1HqH
PevRAT9wp9vNG6qGvBWFwyhsfDeTBwCoobQ08HOk5fXqZG6TFLaxYAakS1hK
q05WOf6JoMycVG/gR8R0pQMJB/Oh1lbMTWHnfIztoR7XuXdUvSJr+ABPkm5j
NiCQ3teDmiwcey7yijzozaAMElpE/Kpci07rFKcJ5KifedW3T0qj7HqsHnD3
GycttXL+dGMGwcpx0qhgaB1n1V1+wSDEnMZq72ayZNbAjRqZVnqGeE6P9R7W
HgZojVFfuGYIuqJ6SiQVyQ1UHA74bRamuqeqhR/vw+vvRx32nYHm0JYmjWFv
A2Ue32HhRW+N2Xk9o/w0XLJjU+egKfkKcBCqk5lRO4zmKTB7QiFFiVwlxGYr
rjp7PUu5OTxyZDD06SOs4HPvpgwqXd7woKVxzV6CtSKLxAt2jFEH84qjpvFN
H/RVlhB6oWk0UHxELMS7UEOYuMoM6hZdqZLKEC6xOa0bXx2Fa/WyNzpFPEPl
eO37WCaPX26/ZDf418s5rixtWmqVqwh+Ta3YJwvNz8sTgeni3Ajm3X9DaaqQ
+S4Hgu4zInQY+mOTfIl/k5vIcT7gIB7HSEi1Pb+myuPpFPqStd5nHUlssfV8
KD4ojpxTP9AyPqpHO2g5PXPQgHjXcyArtoaPMQYaGTbnBXKGYPKfIME1MFfR
LMMDmoD15jlbEvZNdpTh7BTgKGlhXpuAuzfku4m4kOAJnIDMCX8XeOYWGKpo
5QeAcc4M1SAfyeg7JgFcXJUM2G5PVZ67it1wNGH8vNTw4qSJ7SWZguDAWlxa
JVnO1HjX4MRfgSMkkDsX/GlBWAgPwSr+se+UDbJ5vyIDsoz7oe8gxS/qrczt
yCIfTblikJ8QDyPWeGnaOgPqWlXmz/aZBBHJNwkluTx4Ni1KPolRo/zp1RjS
F9EZswfcUcpkG+lirn0oeGnnVUoepXDJAKcxBwhpZ35oF8PiV0Xw6UP6C7x/
K03ufvA7atrr+lUMwCQoE4eGlwFFToRmbEDjWEICejFGRAg+HGFYlSoYL/zD
Rx9kDVGofDvUZ00AnPsIo6Wl409XCftKqnX6Kri16gkTWUL0mE/g5WJ99Q3j
TKW0jPOGN+ka5yXfYFn02IvNTG3lUcsdJgd9NZ+J2uXZ6OISVzFhjjorWRRB
bazmDzhK+7uxRntDNFEC9GZX8j0U1oUc4xh2/mIVh/9HOPxWxHA7UK0palyH
nE/8wPrT7Y+BfRVY9H9khUJBYgKQ6xdiguyaEQkQpvi4MEsCr0DloaEzsUic
zZRBbejhnB18mZ9ppPL2UOR3TqvH7xDu0IcEKocruLCGczBCg7DICaZQ5Ivx
OSr1xK4jU6GMjXlYh94/rSRNoJDG3CiG4dsKGmsWKn7eZJoOacbW6L7WROto
L4ojAjAwxdweUd5HM8EX0aAbKIlqokoxg/FgStC+tLtgFNgh/7ezfHW02PvM
0yd2V9z+ODDKrSIMUXbLCrt+tJVTbOZLiNOqSJ3466o873c0Mm7WSnq/Vb3V
+zEfGk2F/nmiCUF5iD5j6pzWXoLMUXF7DwwncgrGGbI298O7jr5I2cz++1xy
igyP4VP6aze6rbi4lJ2/ufBhrON6ClLDDWi6R0r02rqUHXOi68E1EVNMt2N9
LwGby+mv48qs/+Q4PBk0zTem/mPbW57QuKS/fA3cstHn6evjUWfxOXVTH1Xy
xs8R50oSQvZng3Bs42cufMc3+JfQ9ew4IMFbTKNAn0+GQBKXruZPiLRYrcEO
nP6IFCqtG6BS9Jssx7who9ni+o4VVn+XiPcXENGOv2pOM1a3DayqNKvzHCvk
PBHfLPEZqkgaj2wUQA680LKM+DYPU0C7zWh4IdWR0+u6g39rVaIvAzANVuau
4CdpSwZzbqazrepyVsKTnwwgkPsN8cav5CokVtO68juitSrjkZoAAzjYtYqb
knKYqYSfN7OfJuAE+TcinJW9UNdu86eN4XCLdT6usj74lAIzRDXPw6sb0e7E
frfaMaMjP+sWp0eanVJ7f1P1+2hDUmbeh1cBaDl9lZDaAeZSTW+8dxtpTkPq
mIkKN/aBW1M/1wTXSLsMwOXsvzjEEwYR8v2kQnhkhwdR2Y/HcXWqoYNzoLeN
GRtdbDTyw3Q3K72MkYSbnztjuCuF/lUXpZdAoxyycTK67xycqGGtSCeDAvhz
bFJ3FoFH32O6gDIy8z9cLqLYOUj3nAZnLjo0Z2lGcIZy/NFXcVr7Vn5fnp1n
THRr4cE+toxlaU+hnNMf6nBWZRoIvV9iTBOpx2RnlPMdRGhzzuad/0V9z2k6
6l6YFXYgzzMjDXiQVqq0nZ6zG60lGGsz8O5+Ee4ncxWM9zh/cNoHXiDvXewY
KkPNflHoYfL/W5FaGtdsCTZ92CXGlVTQTY5XI3ovZenHKcegk6FwExzdVffm
/zo9mTwtUz9w2m3Y4BlK9S2Gt7C9JLR3bBIQCS8zcE4LR4GiFFiH6MdZGLef
B7BAwOG21qtuS7QRkS8NPCZEKG71Uxi4dCqnLfB3xLhk71V/F5ZkI476SL8g
+Bzn6ak/ZspbxhA1EqDiML3IzW3FsYOKRUeBuVS9J/cPsyhbwXfzm55nLgHo
CMsttXqXaXO591ECuIF4Sul3nMAAUlnxCeSMU6WLkAsqnbbq17dT2vXviVgW
zUr/2Lw4HabaHTP7qQ0mxfSciWrCjDC5BKNaOECAi5BoQeQ9uk2r9thLRtmJ
+2EGKS3kumBtYN7WRJg7tlvPwGcUXURWODJ3zB/iUDnLPiTM52E/2ENsky7k
+9uA9WIEeLD1oRm8orxK8K1s6g+KhzKFhwL94rrIfJcxZYDfd/VzE9f6KclK
DpDPO/73uROt7bI1pfpUwlUEGrAPeMcEgGPVJDw5sGMZbDXwLqT0wgYKoC0j
tH82R2mM+iwqk6Jlu0+wBSW1j8Ezrufm2xYupvVNYCQBqs3G9W5yiJD0rxup
yVMqQGOr3s7sqMbsv3VGU+MzW3hAaPUtqguJnhGEu4YcENrqSFdfK//eSAFV
FXpbpA+nKvDe+j/B7alPKQNnhfm8hJ+T3reErjXgBagu5EpPPwKdD9RHiYJL
1yUuiyt4c357XWuuNFVDAbxlv8ia4OIpJ+dXLwDhTB0PuKd8WIMakq5N5IEc
CiewcGAS1qGeR8CT+eF9ymAjxrp7YANHQlcOwW8H7KYjHviAbiLt+bb4rEvG
kHvzEnA4IH6lkbYdKKvH6QnPa++vQqE1z5PmhCLzIYcJnYfo78E13s5/v9UV
IVVQR8WcNH3BdmgqC3Q/ZtsJQqI7q5G7FAhLksXdH1F+rkFPky633OQiNIT9
U/LcEHkRQbDMCp5vuvVhPSBGNmM53rYwMU41SRurGeNUTpD8+lJQJVqmAuHE
O5TDvLOuGxHXH8/EdiTIex+YZKAjCKY4zce7g5H1x5TB+2JFB+hmRbjygJ+x
6mK458TLuqc68fGFtJ4rIdimX+1oF0mqrAUn1JM+f6CwvJM34dlRl0ubz6yQ
Uibi2a3eLWfZqYstt4l2qjVoKUWsoHOWwc5xbCljif7tsUQDhVv6hFYm33eg
nadpC41cIxV4NYih7IRqeR/VYRZzAm6lLdQw6/fd4olvS+tWxStnCi1mlWa2
YGDSyecNjl61u2KqVhYS8J4IDV4Yx1z+WeT08biVgko1punaBDEsF5LHIzIU
rS8hKA8138VOIWW/6/ymw7Si6CVsAQr2K/1/mkDKhmlIqGuAuiyZWy6bm2gx
1EFLp1BMPZ+D+c2YK/19tMp9aTtJLuxxGByZxvGfgTWHdLfmlmiFta7LDvug
AGm/Ppj4OXFzO+t2pqY5BeJa7V48hnVziq9Hn7/J2Z4tvj8Z2Ct7/56oTCSs
XYFxOf4wkx5dQhFVLhOWxJNHZn1JW3BuD05UVD1DwZ/Zg9m5PfmnCUN8tmCx
+bes23wh6jMOTEm4YuE6MMmT0avqpKSDwsibeejjMCnme67uDC+E33Aah/QH
e6QjjIu3vot4XdNmJPWZ10lO0S9STBw8dbGY8Sr5tvMhSi5fRC596u/sxq4U
uSwyz21uso8rbl5IfYJU0MoreqFHw4Z7zlIS5pZJgZHz0Ov50NMw7+IDkOEF
dEDmede3fAjqvHN6YPKaOcWsMmmoxpqw9pM3Z7MpeIWc88ohiixk9GJIDGAA
fYd84cwLI6mb4ZWBrKY1fxDx0FjSxIwlCPjoA33Dl0xgNmlc9QnPIyGlcJqw
RDanpDYqFdmCrkAcYPmn/Vu/NkDYgIXLQ7ZARnhe2BFT+2ZAPK4G4U8/+Vrq
ZStZQHVHRj5LNvPyk6JLMnY03vo/Z6fL2oUIMgD2Z14p8zywlWRetLVYtxGq
0B43wG0cxRmZvTwmSYtEvrfxyhISk37zmjsZykhRHvADl4qi3XqKmMNT5H5P
xRb6zcmLOqT7B/Xrwsg0b5wn+wGtk67+DymgteIUFLH2hVQTqwtqewPGrAWB
orPtsgqXfQMtrTGHUpuL4OP4l8t3ClvakhBYh+FgyI+hyQs01KVx/KB0BIVS
nMmCpBqqpUs7If4Qnfv7TWH0Zsii4aVw1LsoNZ+ce50/4uSmHcBXPgswzQsg
FZwtYf076W8WkL/OjA+zhzbRVFpY7LWTsLKDYrMYdGd3TEl+TZXFe5FNzFdM
P4GN5LWwWjStJO/iYaQJTqHn95wvaPZ+vl6UpQ8H3B1x6Pf8W86YIHYUVHAh
dUPBk+2+RvVQ66LUWsxeh6VC0LPs1ByHq5RRtyFgB4WKbr9Xp1ZibPknOXjO
jFdFGripqAiRyWuoJqb7jmBQ/uyD+JV7/IeieVP9EUhD/Y2zzrn+L+t6RhhZ
Lna1J6yZUYrlNowDsTQUIu0NUptF45R8mYxQnBjtX/sLz+0D9UBamtb06uwR
2kAC+RSAi6+HX56D/MsB8cFxvfug6+ZTgTuNIepT1C9/3d3lN2wo+6sf9Ks5
uT/dpqKwY/D61pIcZSC3D/l17jSHDlImXnDXTk6vl5r0XbFwbTYZSUNhTRd8
jhfNA/lvND/W8EceRSmBxwn43diuxim1aMcFUlZ26ZGFIP+Og9Zhm3xc3tiw
reoug+8CnE5SPEH2oY47SqHoihiGtVx2BDeo5itcCXB2YDpJ8xzWdueGjtKl
izUvQ/O1l3hOV1fzx33R3JtDYhI5AjpdW+0cTMumEeiOLYPEvQsiDfTew0hk
GPI9t9U+y+cR98TJSxm5AvNYgl4zYgpJsIBzGnmzltfTDCrlGTeOYvvbfiT6
WolruU9wKuDcbR9zGcJBTj+CC7iAYABuF7SSmHHwH1LTaYAer/ezWupm2OLe
2QbmF+5bXEy4Fjxt3CgGidgM7SA+OuxFegu19aKojPk6x1wgjuzw45wngEmu
LTNysgJnSjyLtZxlUgdPRznZFs9fXnnAniTM7D7zHEBZLLFmjNiCtpBbPMJ0
fdi9zQRwg8qns+bte00NKT8BZBEZEhACoWW6eI+5/w+zwjeJZ6tQ5zO7Flhx
LVDcjeippDUGoRe1eXKPVwQLJjzkCRX/TxdBIx0is6boZBV/7nF3mhABNnGs
PpJEVEDy3Sgt64M3RkMDSlhHq5AbjLPuPrnOtkkiAJkxDOOQSB770Wu/i0/r
ufhv7zY1ntH+flmMDKcU7YFUjRVSyDcC/aAkH4Mzqvpf9igmW4uIo5Gp2vO6
HH05wRcbavWqxfZEMgTWJO4UVSDQXY+oNERpybYvHuJoAPBq5Bp1q7+PHQWt
T7gG+FuyHP6Z+PtJlsMChs8c4VSB0mKLYWwktcdCNCFuzubtH1Cmc6B57Z1A
qv1sCFfIVlkdvDDgYXOIb4V64yE52s/D5j9xyhkkosJXEnNvuczlofCTlBOM
M4DAcMrIXRyp69zNyAVXjEgiaeISFDrrxeiHEYsobAAWxFdLsIQc6WcVRVln
jugdE5zBdPq+5sDSjhnj0wWi1GcoTvFaxSLLj+1dPjBy7Bd9me2ROuRmRQfO
NJB8XaK9opeRUJ5SuZPXYdoFsc4I3fCb5WKOtSP3ngRlog5w3w21hEtky6xD
ZVXs5T5q20AuMPOIm1HaS5ahMqKitmDpFj49T3oDYDwoONd0+l3H/9Sknyje
wwTwLiRhGxHM/ZsqSb9bmYqNoe+C3KGqsbntoO+rHDflPn9axXYsglVBu0UF
Kb5uZBXka+sGFX5MxvmwjS5/whXSAPmcnB4AqGLOk4oxbBxQGQGeFWYHkJJK
BGVn/Qhmva2s+kWPbSrUD1IXW8un6KTy7RNeS9mQB1tu71i8kZX1jvjIrTUq
1VBpzLQAGbY9rT0sqLCBjPjWkV0A5EqdAw9V0LE93+g36VNt1biNjZ5QYTnB
Jc6qdOZ+O3I0dc6eX0Yd9ZSES/iFiEr14mA/X0Euj0sTxXwTJpYY1UbQ2h85
QJ5Twoi0s795zZIWW0lDWY/gYgzMk21pdtL1g6EXiJGn/cxbVxOi7scGf6b+
gb6UGIMllj+bFClO2VCqnq77Mo+OXYEG8CZbMx1RreGfVv1J+rjmKQQDmKLx
01s0hf4OGDHD6Oz6s0lXCKB4TQl4iWW1VFS1xI+LKgKL6yXa9xy6L8qX6C8O
4abKRrmId83jr6IMiAwCyMDJGfFXqJn1N9ooI3ShUlOWUvaO95opdqKTuQAc
rId3JOt8Ce70fNAfSdwfzhO5GOTGDYbzMguEvIW/KofB8o169U6YdsfT1a1k
CW9+U5pww8Uk7CwESFZ2YAD70geEvQjMitY1iyFL6PcokuutCW5/1KYScNx6
n2ABskq+hT1kHx9eaHhaS3lZKtfOBcKqBbXm7mWll6Ity2uiXFcY1EmPp47p
Mc7Tl6BAJAyyQOqeCv5vYGmOpui/k30AoFMnrqBmdexnm73uKT7aVOXT8H+K
Iy/FcQ+5S837aw1xT3QMkUzPC7TQ3eQjPXxUkX6Lqrrsr3s3YAuY6Z24cFuK
Ar7hNvxVGoouvVD3mIdjHpYRWvwus2EjPpohjF7VfUDLeJjpoU+R2aqabpvH
NbP20tyMij+9ADq4GsUlH9k+oICQMuVXz+zAjyhIgGZzzvlb6AUkQsAxXZCy
1pVNxHWK8TQBlY3mD9muT/a3kT4x2VxLie9Ytzcb/d1t5Fv1wqerVhhyrSN+
BcUQ/p23sAu3D7xhhkwCI3q98eMwLb06XxsZ3CgNnm772uKaDmljdoLFr/5n
jIj5C7pS46ZQg2GIoBk497YrFsgxRx1+zw6K94rt9s+lTmcuT3wHzITuPuSz
+WjH41+XxDtEHnX505V+k9hZiUybeHlcfGeHi2qZzUWnt/rCkJHoYegD26V5
oRHvnloT+1g9tnip/w7gRrHluPrUsMUQ1XxjreGP3KqkcthEXEh5LrqMS/yU
LdCzkPpiX/pWCpxEBf3TXS9BMY59JncvigXI+vGYF5pn8ilru9ij/GyDa2VT
V3cnQiWnAoL3ClU/aQYiwfT7LbFbSCFUjyV8raOUzAcsqH5G1C3GbVUjWkw1
bHYPH6pwgSx6HtCyorV7HJ91ttyWre+arDYtKE9vqg1ZuFP4X83OADgzEer2
CBt5t8RwDAVGRvsJin/As3Lsctj/cRPT2XIa1P3nBhf900uHxBqpkeHDbIGn
r3fVmkyhbbjRgsrT/GgycdzvejNtOhMR9qtq3P2mYJomP7EMAx8YCvbcdx07
fNzAGoZbqSRvFbGHTnzDV5PAy/gb1tcNT2LYmBWXJZFWTyyeV5tBhS11mJB7
QC8UBDx2/clm5GTnPrSJvoPcbMcoLUZoVWNbdnyBQH2Ca6TkmOymmSz/ohDz
UpnsCwwEpePjCI94NuDCl6EW/cmS7EWzDnwB9rqu5cWYNZGBACfrxxPSmSo1
aR5avcTCI504t95iqvy+2kIBM/ltfGnZPXVRfw1SqYcCGotPkw9rEqU744Qb
50FUI7i82AVdzgOvquU4zQ42NoWhtGF9P6EwJHKW1IUzIxA4BV8GWKG65EUW
gPWjPu/RU2yBxbU2/zOcbBO8YshkkRw52DvggBwvdH4PoD0ApJJiNPuIHmaq
ln9/MpdZewJQbMd7sths+iG7ZWinfhl7O5sSUG3WDzoNmf+t0mOZZqjNkz5D
5fTIFrCMmDbHMg0/WGPo6gEI8xjoT+JU3aH80CbVUNV/j/teVTA+fmU/P2EY
sJTot5k5lSZ3A+nZtycCNxHI8QYQXavdubNVWLv1UVDa2QsekQDrLfRBkPid
BxOi4EVLi9WbhfTC5jXbF21MmLzqHkFqPAfHuew/jamee2qBQ4OhD3b3Cj+1
RvOCO8m+nFj7fCuL3Zx3SpzgRg4+m4wOoIXXH4beZ6nNckHnVGpZAHsXr+N9
4c08S1ZEr9ietkUI5QTXVCpRcmsHEibJKuK/OQltamHVSrxjouRIzjQUZ6oH
kZ2mL4utf5taZq5TP/IL8bRHkn1/r1/mUbdZmCWwASHpfKtZdx7oouCj/f3p
TcIDnXiHSLtRmgqgb3uH6a8vt2pcAP+z2BR+y7wdXq71Un9/DNWSolfwsesy
fn1Ozc/XjPNgTjISp8O3vAz3qUN9EekeUmvnDtD0VhL74nQSO55ICYtI75UB
Ca9KsfxgwlNe4hMPILHdy/GamAf1lrK5C0c2wnUfk2WxrVWxUWgn/qpckxwj
nbALMf611g3m3eh45Pa9da7CPhyGw9ilX+j8uW1UzG8p7GU/wTErX7wnbBiM
ix0o7ny7Wy+3YQTKAS8ESxGc5SASHDkyGoEgChxkieTfy+CR5erGXVhfG2Pe
Fqb85vwfBlxJlBPmBb6ZB/eKGcBjNwRHjWrtU/BzE04DOK+c6BKR1jCXo70Y
xiAXnTEvZ4C/Vk3f5shyxY1HVfjZTEF4Jqpxtp6zWKp7Hs4UI5l0jic8CaDr
YX4DfQ/1mF63qjIMBwhBuHbOiUa+w6OCnwhCKApCDnA2Vnahen+xR/x4sCg6
399xrQ91vuIA4/EZx4/yrqFvuKjR1oJ8v04ex5JIGjFAjbkBoxAjac2h9MYA
6czvwRZpl20JuvuKdRnq6N3jrmlCRKc96kY46gXcXmUMBXleVXDj8TLDez81
GkQlllBCLDOHquqZsePPRJFajxcTXYJvBREeDssepMAixElUxTGATDW761LX
IIiSYEBN03h64BjOZdavzwRf1spcXzOPy9NE8YAPpNiUp6ayrhEXAhMSd37J
GqBZF9FfDOr3/Y3Dap4acQAinO39F3NVAvc8QQFBU4PI7DDdvBdrajn6ppE+
6j5sXFtlJWxkTwTyW5/3qBDRrFahAI4qa6G39d3FCF4nyUEGgeGnlCXs8DzT
0fO0cd3y2wgulFdiJRi+VFPt27kfzj4MurONVp4gAsZ8oCRgmPMxVNUzj9Mw
x/LgvK5m5Hk/tn3qUviK6vkiIq8EyoXpeYhl+pAslfyzyLnlFdtFIEO6DROq
78US8G6UfmWxUe8aTlJhXZapr/7uvS/kr+uobVgBruaFsZR+4sh99Tk6UgZ2
PVz+QY8H/YmZLb5HbLAre4teAK/VaWB9OWu4VSXtgfCyOh0yZVE/LAMWuj3V
xvEz2eIhAwp7DtKglmZYNv+eoPhQBMo+Pi/2JINpwcDM9TEHJYbLoXrmEV06
e5qiLQcLfXSCEiKC8d6vH0ED22Ix9eQf2m9m/t9nE2GcS3/dZ+BryRlTS+Pk
bnbR4eqV3VV2QGXrnKuv9s4rMFUtxaAVp6NbcaR8kpSXLn3VQ+yDD3MXsqkV
CsFp86dyzfoFgbdt+wFks/hvEpySfsPukYbOKIBcLvD3spRJP31p/lKMXdHT
WPHcQzl93yR5bTvDM26MtrJtmfn+kL1Cdhj2OddLw1CE5L1TLejzNSgDOo3P
/4MeY5sOJlCiCUWB1Fgv5r5RxMfsyN/5VlhJ1gUpeXTLU03Sf94NrYVZNL9K
D9Eh4nM82d/h4sK1Ci3JSXd/mH+FcCvx6V/wKEukVw/AGK9e4MKRNRrmkyMn
F1wZHhiYIPfWlxbkjzzOLgdqxb87wm3ualOv1zMKKJUhQBkovtsCW1gLjRrG
kpooEq6RD7qL7eIW0CDy5Yyb7vaXplQIemwPEvq103HBbIWJXmjMGwEH80bq
UrytKUSSzTOa6ex5zQxqvEczPwFmnUaP1CfHbWgDxSykP2/t/KlYOdtz33NL
+D7G/7zAitES0YIBMOvBPFK81BDwgN/vN5BnCGuc1K7suy+Ctc8jq4RhfLbk
gjh26xpVwcXJ8gxmbGLrTE6jIAutZgdnZnecWZicSUFWCf0StZr6/0zJQrBV
9GKvNbHjo/+dCJTPf87tSHBgUxTQ5/yCKfn+2bSgj0CNglGnDWww2Q4rqxNO
Mfp4lwZKWYzw9Rvv2cL3ZWRvP1gEidEUPPJfdZUQcSLA7QyCcK51mN97mvek
ABarPSjxuvFUwg5MQo6UVkVhXgHHqrWNUxzqEnLPdfhPDZFer+1zoc8cZxGa
q/8gQNq7sWE17FUP6p+dj+t3MlT8aujMhchgr1hcPLfWLwa1TDQkg5eZlWLn
ZUnB7bJKDvM62/2LFq4WNTGVwpMkxmLY4jJEbLFDlycvrqt7Y8IZoGn+1a/Z
W5Txqt8IXN8kLSmzbWn/eWJpkxLSlNhExRgEstnMVzjRbptWWb5SQDIZyEh/
ZTavC5CU9ZZhaqWe9We2qIxyFT6GzOVD1F70TWcpeiRV9alrHrv+OtthY2qM
SOq4HJIj9hbb5NhHWf54WlmhETEQjQUo4s5WDlum9KHOrcRFohZNguGmYasV
Q7Gj0O1/OlATCXQEzeqxaAtI3pfQUPFKnoECEm10mpvB0xGZfvr/3t4tmXtu
H+Jm/dRwS42MwIBg2nqL87hCjywiKeE+X2no598YpvIt5WWTeRcbFDYRFjbN
TxpDgdN71ciSp2G7S//qF6ZeFwOJmLlco3UcZTEQMo3v30epJ+c4dFPaowBR
f4KLjYWBeryU3S7JVD2nvZvjfjfm/npR4dMNVTrDIa1b7mXBa7531kymEa1C
T4oh0FEzPp3Iu6OQFgnX1riX+kaf3MLm9pZgl7GjEwZT9nVCvISu2HLgKUUI
wJsah/2B+w8wkAfMwTgyzLnq2KqSA+5itbVq1QIIwpAIJbeKbgSvGVK6RFkm
dA+A6gu21b+5aIJItMwkh6mHxoZVXIHfNgvAQRPi/wbrlnr6y30Qpt80Wn/6
23gltZnHhNkYCotp8efcE1pEkteb7BONr5fiIgzw6vfwNLPI9ZpZUrJpU/GT
DOpjunsLK+kdMd3XufWsP02McVBD/7BGekigKokYEInCm9qjVpX7WC8URJIX
t0RHSMoRuYr7k5xE1DSA6Qh29Z+o0N6z2Vk6InRedd9bnYF8FHK//dpHfgkH
6+X/3X1CGoY3D/qhtNn2JG3ItuRJ2cvdgHfdgU4u7X+MtdHBY6SBxR4Q0r10
9nyUuunub6IM0/ZrgmHUlCHIii5JNfmsTPMVmeFvbLzFmxFq/Vff4vYiG/j6
ArUPeqZ9+5NqI0qxyyogXCEsao2KwQSALt3sO24OMnS6qu8Hr7Lt63uHbYcM
EISOVLpnSdtwSVsbVGLyycDnDiquvT/f3K4Iv0IpOn6WLneiEL09Z+WPeq27
u1Mqk1SSqGlXnZGk2nHFnhdJefu3XFg8G03pfpWjZGZjPsw4Rh9+TZ7JhEuz
26ftAaq4Z7CIsRtrrAXFvhibb+sExR1FZpoqbEpcA/UK106wg2Pig8hhT+3C
QchQTMUntUwjisq0IkU+uBKc7yCVnC7AfK9qucsyrnSPHUh6x+GNrnmnkTXP
GD0NnQA4L+FgHNBoXorEh+DVDvZDeyuXK84hjMsmX9sLDHH1LDhzO852+LX5
5xyJ99dpQdMtb8eawqgl2c4sHdpUFcvO7vS/ED7MHFv99y/3ovlFsN38Ds9D
w/LrvCpv3sfpcteEVTbQyR/G9nWkPlOgWvMMjeqSAnIyi468UggoAuXFfN1P
uMZTgNg93AYLrGWvh1KX7QyKpgJBFKyZgM8Y9od3CC/31TnJk3SN4s+XnPHm
Hhcs7Or54H5nTAKQa/kq5lGawh7CS4yQm7ZifEpbVDXkV4CBDXT77nglhukn
+ngkgDnJNDQ+ir+0qgg32XmC5UdKs7PS25ul0QhCAB02nfGFcMQWrrT/JydC
B5b1ATNdn0sF8lO9QJOrzpwg9c/kYnBMgoqggGVT+SgztnVS7E9+YCCy/lXV
QOFew84itlWZTI7P4SWWYASNAxbTRQKUJyd3jYt6ftRMaCoqg1brRKPitRQY
taIIbkvAvcL4FkjlKyeQPb1WzQrbd+puZ60jjomC6C2L+dvUSVipQsXRxCaf
mECH3lsJwtw9Njqf675Kxs9pSFEectbLO/VXwJQGyMrkzuy/ux2yiEoYGAFQ
Q8fEY5JeCiImcn8GflR+RrYDM2OSmfCwnL3DKdbZ1xYRiL5LWSOVcmzbu/BK
XdX2J1M8EIWOdWo0skNATYlozW2HGr92Q9GbTrRL0ht9Ib2ejQjvnzHQ/fdb
S86eunxEndxsriVKm0Sox9g3tSuhjlOkToX97Wex17VNMFajxhlv8+fTKjZH
v6XpBW8KOmHyGh4AyBJ5nuTcse58Edja6b4Z3W8fHIL5pzY4+v+kALS38AID
tyE5p6kERhpdnwPpXc6dm2d+1r1VBE5p0gLNp+ocWwp+1574SFGFKGe/W2UD
4tl5TLpF5NRcT10eUq9FQMASm6aggb3SWVJjKhr55I1d50AWvgLR9by6yBrH
Bhyqb6LkaZESzyMTySqjOvSK6VAm25DBpU4GwlCUSO4SghO0jCdm1Psk8VLr
xp0RXDDqIafZaHvdUyas2L8hoXLtM4/rZyC9otn4kiVv98Y1VE0TdDaE5nHY
2Ztt7pAuc8RT4urq9Gfdkis82IWgUi9NmnYtDIRTPmKU+r24zrVptwg3ldJO
v+uGrFsI/lfVTlE+swOAHjZXj4co9ssEqLHl504bI87yFH4fs10ukk3Qh0F0
sXF+GuAPxX/pVsyzj89pqo42CzAuL2EUCW8moxkbUZvnvk0z6zn5F40YTkte
CH2iVcy2GDDcCG3X/XLovT9/GVsK1/nQAQUE7DF6zLCKpu9IgfSFk3XjjsCh
3Fi2afT0j1jowBZcPHaAZCUdpDXRXVf7Cvz5GSdWcbAiOaDwWr8ztLhnFRxv
9UjkNiBEjGnNOfjLbx5P2dsO3xFCRYoA2ujdF1PZwv//8zrxAcQxSRztx+1H
a2AtgtiEmyHU2pH0QBMkTuaCbPdgLEuM90vlg4idkc9f41pH5dMttwz3IQVh
tr5FPG/rwFUs+KAslv5qYngsqoucq7mfj8yOhU5NNj0D57i54BKIOcQJ3/gR
MoJx2kdZAqpUfiyDOgVuRya8g1HrGzbXX25mwTk9g1Sj+wGg7gaB1lpQOOTV
0Klc3ZC0FLdnlc8Bq860wF+kvpSJJKOuAxX2iS7wlkXURraT1a1lxod7lLMW
pT/80bRrjYJNag3Kx9kGHdo/Yc49jcpkanQVOeZjH5M1VBzvG8uCo+DrQhBb
jNrjJsuU/8q7ZFC0lX0E2nxzsE8cmEud0Atcmg253KOXNZb/pDXUA+Ef5g+h
22EnVECtOp2CYtc1y6Fd6lWDElUEuZfqJpse4LFI2KYrCQSPewa7Gzq8CjGw
pvtqfGaQkyK183bKHQy2LC3PE5LWk93O0DHKhZ4to8bgV5wVw0KL46Iw7ma9
HBec5mvWyuaz0KsZIt9DMDxx+CUriGA8HHt/pKR6bzdR/buaB1E2tNn60i6/
DDzPK93vKGBMvPnvmiuZZppaL1dt1HM5tD3kJMsnWECa1nnrMQVUYTBL5kxL
KEGztAbhvNVB2Z/46G8/VZtlabzejb9jC5tP+O8HD5EzQ2khKNcg7OObdrqt
UvocjBaC2zdA2L/e8RjoMTS/irNNpmaubksXVSNsxAus50g/SiBeBy2JJQl/
G4+kaHHG0IaMHE/yNdm3SGajGDlFCeEJm0VUnWSoITWvevDpNIibzpInEa5M
rqyYtbf9sq4iPRptGITQTTvAHNn5n0BqvabsC+8MetjQ4QsTs3gLuklpserV
EtrqvaOPEU7zE3Uiv6Q+HI3Sv1xQnfFWRC1oQDRM4ywS2uHNrnbW50ZTvzYa
psdUUBy6K6q2rJQHySiL09/k0CSHN8gsJb8Wwf6kRzKknrZvJfLDn+X8TkIV
voGygtmik8jv7TWVxyk/fBIfTB/lPFl/n74Wl55IKw+DBu6GsNOr+O2OjbWd
p/YdF/pno365B13nezmEM8tqeOb9+6yPlcaInJlBMXjC2JAQzOfMUYEpXhE3
RcHigDpEd8FjRPQOAfoREZEHyO5jGKCVN4ob1WO3FgVngestTaAVA5pJZ3B/
Po5ZndJrEOc+Hwo286tMb4WrtNBQj44ZQn7dqyiRSdj6FbcjBF5DgX2CxzKj
0OcfD8oZChKM+b9s3qfozb5LI2v6qCb1pfCqngt1NP5ZY5LuLp1qVQecIPl6
7Nq6qcN2aCPVLg55czubx3lylGEXb/bnOOOLFYjXgh0uh/g+AYAcYLmTxSnl
omgLPcTp7xevy1YXTg/989gzbdf3/lgijGbuU0W1KKIhgZ2sYU7C38AnGzw9
EZesnGThT9vMWqcNfqe15JD6fB9OwUXSWQL2S1ZPScQi/kMr1FKvhz8K9Ans
cgwM+/J+GTqUhgMrvet2VJWqqHc+GqNtkjpKgHj4Hq5KKfdB3MaxAWAJpGkS
DIqBUJbsB9Wr77woN5C3wed48b81joAzXWRXwUYUXalT4cIvCQihAzhEXxTz
KQ0S3hbNsrn/yB4jPC8+IBlOLEYhpQeKtnTgRsqp/TngGX1oKKuKbPabp6Jc
R8js/rliDqJLnUD/TezyE9/pHbROu6Z54CYkZFeE0cwlBimYcDr8SZB1S2Zj
mx5RRR2m1CE8emy0rqaPVFnkDu0LiHzXCF2NxtOum7sR8nOCYYabthUguew0
QzCvQe4zujctVLFhn7xAUQTOXlSynTCnsoFC0L1Uvw8lzxrdLqr2AkCg59o6
/F811s2pg1wcWZ3vHMBEauPpLNXRikl9q9pSpHsvVORoXiAAE9cp49nypkDj
RrbRdKbSsqhCv8XTeyb5d0ZicKVk9wxAtsUsqFR8dngq+oncORSaNrlJ8LYq
biuwHfX2z3O0jvS0fBjeOWicroWRKlbgMKCPYNPg+QVAgJLwwtZhOka9LlIh
2Y9i9Jdj2dGrHBJ1FcOQ+0PYXio/b7kQV+XIlfa5qz5WAPsVzPiLLnhp5aEc
qajU07OLOOZx0ntqfTfGM2mX4MuHf3dfZ37pv2bBTnod9hyCrIwiuBT9INTK
nBWV5fQaRAJnJPsg281rxuK4uB+iux/7SRbycMURsCLwM5Lgul2ZMOkcNcBa
8sEMOo5W1KkRFp6JV7TE/5NQxYPPR8oOssr7rceGSEkQnibgbG8KlZGgcKSU
pYuBvTSK4aWavaD0l8wUl2WqR49CT7taVIBCIbJqx74IIYA8kjSEkmDZb03z
8CMSkepdBsVgBcMJ5sEjOAyqIeqV5J3Vp0y1YmkdwuQmN1NkhRscDKweIwoW
5L3PzkKIvJWvlkug2S79W3HX+ECHfGqDAm9nhenu2X2SmGQfdXvPXdSXezEd
AVCVmIeuUmA5xMAEpsLEVE1v6jwCVYeQkz/caiYI08kqJo6c6m5xDBpo1+Iz
yQGC00+3O8moAuf9QX4Yh9L1fffiBe5xacvliU0flfIhRZU3zJoeyzW9gWhr
9FYXq6cHjeOCGZN3ci2xa5MxpSrcyK3KktQk8MGYWsbZ9i1wKACIyRCtatXP
5g0AznExgQGcUcXiKRYkoXSoWB8dbl7dHXEzBi0R1ujUibt3hq72GWDwTI0D
dgovPT6ECRXAX2813Tz7fUwmlsrMvwYjxTKn4qddGJkxChCqAfyFxKl9O+Nk
JjVkn6oUmWDib+nnrWsOVYsqNeicMAke6KIKtcCqEjFWJrZoV0cM0f7ViRdM
VBdrFJoHCIwPziSpdee2yyDR8IBZMfegmXZJ68qNE6Q4efZbfKfyjQhDxRWp
aRE6h7MBJsKGvk9SJtgrtOiq6tKfr72FVJpWIj0IawLdyM9fM/+nToBUEF5+
/6GnIhs3qVKLOCuc80lNFCWlGf5/ehIiSGt3p4xxkGhdDh+34rQ3GWpWlLBM
sdinOsIErtCRNz8yaHLOObOcsaJxIiiJhMS+seGLtlaunNP+SpeGrIxawrJh
tbPLADKSEZuvwvMDQRsDntEQ+HBXSvLn8uBkmZqPf5K6YCxNRhmZOtmXVeve
slrhS1Mg2zGO8oK7p9vYHJi+fGrt8e6n/NWulcS9ZTaSi/4hytxGBnNjrhOs
vI+C0eRY+gJAAJCfAiINAUG+SYieMVxf0B3CUSPDUd+ERxxo+VKXOiI33BIv
0ZRsMmNZxufzKH1YtEx4+f6SwyqvHw7DxwMGCVy+LpWqwsGg8BdyQ+oyWM8O
7igPro5kRkzxxPGqQVh7kD0YaAzifafz1WzbsNVWdH3+efAWDHc+NBlEZirD
kwiPaHsZ5sPLsDxSH7V3pHrm0BvBOXOOg2lCBjtX/gplO9R555wyEYigraIk
0Ev+MjUMsVMz3+7QrQLkUDQKT2OLUrsOmLxXu+rmlySr4NMXaUvGEFGpvPoY
Jtubkk8lkEm64mqGxmriVGB9yFnh1qfJ3G+qDR9tyoI3CRgG2AbVts4ARaNI
6B5hsSAVTzXM2XNeTlP9vf7X9XPhhTfZnTZWuaY3uaNNX0gYpPyVq8WhGrq6
PI5OEnDdBcViuzBEyzPR7oM9aQGsveu0DLn4nbKDizD9B8lgeRE2ggcPDhXi
Cz7IML4fZO1v/a1AHuQVBipAv1BjBRkLTSp/Kco6t46rvEAJweln8JshT+y5
a38I0oAN7Im65EvHnPo+/hLGxbS920ejQgCD2x0DlDofMqMzM+prMv6niIS8
tMAhqz2gUfmjSb4AyQHdnGqy6KvHAHHo0Y9u07ByG4LjJGSAVywv6N8JW0X8
na8vOoCv9RQOgo1UyiwMQRc5Cc4ZWgyr7L7bEz3UBEnEFovHlB71JZK7CnxO
kZMlkvz5kHI89P+Juhv3DH36jKVcY3UbRE62gU6H5AMRCp85wjAmIg5fgavY
m7jYEhni7bJwG7QoEub4O5busj2tsQHQOJQxQRcceMFquqPOrlGW3YTyQcQ0
MynoVOK+PoxhzX9V/TsupZvpXw/SWlzWBc0gB86Jl0Eu8szOnYjevFBQQThg
UWLjD49A5ZE7cfdNjVyOi2bpqNMhNuYeIIrZam//IjCcemU9rFoEt5OmfDHZ
1PoNKdMdzqEoq5+J+ZTwmgklQkst36s+6OkBzuFyOb76v5vrRVUVWgTk1ej6
+5Er14dC2x1a9L89W1kCdYhDb3/xQkQkw7kfWe5fLLCONj5dyJc5IBhSzir/
kdOX8nThxv4xiU1E0bZTXI18i3Au1syrl9a+IXl8xDBYoXR24qrf5hqC4Tgx
g+QlHzySt5hPIh/EqiOkurErGBdtQ7ISxv3Nxn6xm0UsoXtLJtCSQTfkyfvz
DIB7kFbuYmwD/5NkeVRpgjy6KT5WW88NSqUqeH32nCcemOkbnrwLT6ZYkPoN
6nzsGOHofYQNg8Xq57sWH0ul+22zmoVMxyPZsyIzyadL/iRgIrUEKz5jyWob
Ios51nBm+/yPbuaSH1SJKQbzwSOyMiDlMgVmGCSPi2CPto1d3E6l6hVw08IA
iqk64gTx5yV8q1lhVA7UJ3XyULE+x+HdyUFQvVeIwm7VDKhSYe7TH51CkWOB
yyICopseUOh17KHprg7ws/4P2aDEh/iG0SXWE5LYjEn3qIunY+rb3qoq5h+X
aJQpVm4eaYIacuxnoMm+GOGaWTtNmUcNKh5hqzvJ8i6NM+ezh+KCbXBpxn18
8u1JdtsEhWfWAMIwsEb7omtOH+VHPwGpTUOxWAlyVTcC5k/486zZR+Fijxnv
1KwkKARjZSW3UxTX0sik6EVrsHZXBqV7duNJYdkQM/r8DEnEBzmwd6w9fsN2
fu3pt2L8O0LLvb0hrv+ydj/wHC/Pm2CAVFcyjUTp2e5qBdwbvx2O+TtjPKaW
Pp2go+FkVySZLrrQ7PDNPEiJSSxEMXa7RahBkgGOXSUfAZVQgD/VOxl9wbY3
8VbQ2PV8/60HQNf1VCTY2yU1PKULxHW4gUjcJ9kgEX7BwCEN0L6Iecm3Ykfp
XrtOF4IP0aPpN5XxZkatBJkwF/8DUZAa7wrllDswfo6Y40K6By++/drepay1
7KiE84aUQCHrgAcR3fV9ZvIArv/ovr3tkZB7eC8YoKojYA6qMpDIBmAATGFR
n4nPcJ7DmjFtY9rHnBzH+cySrziYjA1NYUouiK1lE6tgAKx3sPHykLLE5hhR
L8Q8HpzGc3fxEvYQJRZGaql7GTXBqD/pmuXPaK5CaiCeL0L7rBsHKodYZh0j
4scDxRmMSmfREY5nHmjyeKrFMIOSu17KIQr709EvXIQs++x3A3osvUjYyMyk
ycbDCJLRWYIHE/yAZ9MF7N14lSPvEivJfK7/rM5WLvhLM5iVETjQi4ZQGxWY
3/CKzDOX1Cs7W0Dgj8pX/Ux1SXTGjVW2cTbo4/dZ40/CEiNLvvqn/YVKra2o
mjkltjjMqxnbzpQdeSI3CHXrC7I9/TXQgkukbWUvJ9MYZUPBNq+2yuQZEY9j
DAIXKmBVKlA2ycQtlguGwo4P9z9Kh0Wd8q/Ijlc4YM2Cxc0Vh0XJA+sDuXsM
z7FgyiwwnBvrgQLD9Og9u1Ke/1M7laMaTu2Kamzakev0buIh15KUeDyWK49b
q8Jmr/aDJCveE28tYphrBLSayvQ7pFlRXRmZ4Es7cBJsudUQdH7+U9WF+ArJ
RUZCAmvy/H6khWES9A8qS1qZfeXgT0mIftIW8+EgnWwTIdNEnkKbdiNUJ3tI
W7IieU5FZhc8vuBZCCrSHuPlOEmHffMOqXK5UjHYcv2DDD8RWqc6EiuNhOEv
HUzdeUGBWDVTYMBrkY9Wjt+/uZ4Mbu6WqocCvFvX7oNr8KaUmiO6svmHyrYy
ZXkrH5FFNkS8wdTCjFi7ldhRfNceryo82IgifMH/kkTS35kka5MZ116YPd/d
5rFCUKcxoBp6KiaTMfCiaVGIBBzBSI3jdW74NvBiQKvBnozYc0TwUEn7PtNc
KHtF/jjoHf+L+Qwq3+UfQHwMx5lNYE5D8Qa8l+f0kE9q1j82c9YG3lBxahh3
B9PD0t2nMRBz0yF1G46Po8Bewc06Qr4drQYvVes2nJKuDmYjbl4+h6QI4PFw
pPUF5naUQsBUAKVsoxFPziXv9y0LjKXPm0PMy1abbo3ARkjOJ/D1y6C0ncfI
H86k8XNu/qQQvpl9oSNvsJdWYZkAzYPcg6g73iQYETdrUBgxIXxywWMFXJ0v
SKq3YOZ+jr5rW2sFsoVVBmbUDGXSci0ir7DGEP6HVTuz8MEYf2wcfAxp1+Ss
9TbixSBQFTSmAzr5KrUCxNEpGEepj+/4Z6xMgb1bPVxcUWcfIPvsOHdDYjek
up4v37dglVxjkzrxXUw6D3EPSeyekhSkJy+jyUPAoeld1RMZ4i18Bbx1LgLG
3JMLwTQJgiP/WTy4U2N8GB7Mn8DTj+spAUGQYzvqbxugb4409VatleVjgpCy
MqO9vcfnfAs1PdIrEbU9ypJCuy4x0roSVL+JVl/V2Z8kjbr3PgqJaiwajgZU
oFRrFUrMZp8NPA5SxPHlwttRf3hfpnhqssXk87iKN+vq6P2n5oOFs04NmSdG
jihqxrl1A4LG5Yr+hvAN8nJPEcgFUP8DqdAA5uEGgEYAW906WRKSHy75a6BK
DGp5l77xLUop+M6Oca+r8lvn4c1PpX93gRsyIHWbgUCqh3k9iQs6ZdfnbJ5b
VSRC4+M028YEgjgo/MdlKXiQ8iDw8jB08+9nHKooFuqti7NagIyFPeKAmxqC
/M/iSTfGzdq53iZTwgU0ockIOzo+JU1LeTBOb7crsaKrp2TPrVFjV+z64JSF
CaA7g+1dfShbVFsoxO3g9JzA6YqOjXDBDRFQl+4+GWX1gb0nF5aivSptkW3u
RbL1jv4S9wEi/jLgRQpsPWhZNr0tDug3z1tkdBUgZBX4XSkaQ+VdCHUa0HfS
WpHL1wcXCWubl9+qKO2JmVpOKtEK3HtBExbgdceL41n7/eZBTMsIjMkt5QZF
UWz3I+5eddq9NUQCk06SELwS1akCPDEk+aKFNCveILr/cQq8ycbHW9KoLbsw
4JnmWmKpCzaoFjEFEY52yPa6NH1vr57cNVMYv3RsCWJiMGRbfgAkfuaG+U8a
uBrJX/QgSkO1IxmF9hN7mfj03TZ8Hyu7FsmNanOQpVFYqIbI1mlye83CYSWt
eI5Z1XwKNtVk50nZHNiYw3nM7LOdSyTOtRe2I+yFWW+TfBd6tI4W/9UPsi1b
Dx54UZtpsrAf2HAzSA9D4sdvW+8qQfZMnUKxbpf23W53Gd8E/u29EJhDxV8l
n+mlV2+a+FhWXuYIDirDwBjuANXK8oQXD13pNAb3iwPXySlinOJWQiPO5ry7
nc7/F1pI/CJm64qU9cqI3nQK8cLljF81o3dcNe7UpXFb5LhexCbtyQYsQXbm
CMDLXvPt8+lB/SdC7aKDC3a6iSWJmDy5B8p4okJFfAYILLEs6kcQ+aVGBZ3f
IZkLunNdaJWhXn1//3z/lqyLVdaC63lzUtnLtWFTIg3JToU43kMABSQVFsxE
oAPNpDsUaFjfL7DbmXoWHGzMeyTkdHtaaPMJL2lcr5AEPF9XT4sVVVDHUEjz
cmuGT3C30oglkjVu8jJpxNMkVzTEaUCFIBRks1OtO4FM2JWuLK1ngjtx4vzR
dc+/Xj5TpxmV2KIRUP4mZ8JIr0EEzJYasrIoVeHRrOMdeNSkxudGzx6F00eI
byO0PEsphq6eyiun5FJiZKhkzMmGd6dZaF1NCr3GyVAxRPKc4uHhqFMP/8Op
xPwE/x9wdKWz47ZN2S0tdpYPTk8jKGy8efF1IGhwdTIMEnkazH2MsLyyDXZ9
5GuRyaI3V0nF+9ZBZ84bZy+H9+CuRSYXp+8i7xP0rM8WrT+Vb4Jftn7uSHYu
hbjPBwnG4KvX5z27vmo4NwcgxVVB/9mq8D2fd/TVaDApCV1kDj3r0oqcHioC
xOQ9ed5jPVQd7VWw3OsBC2CbtsISG2EC2lupF4WeZIhthqND1ADsR1Kh1j8y
LIs3AVV0U8+nWIXbXTuEGF5eF5t+li+KhfeKUWGDdJQ7Acy2uSTJgf4YLb/y
qsdzWFWcl4czqWS1fM0OZcNkSFstAIcMV/AS8Qe8CtKvs8Y04JNH+hdvRZra
f39UIYVRd7xE8a+cyWY5rQ/wZGWTBKq0OvqwuTw13gUtYAUprl+uyT29XxH/
Sn0mnmsyiqzE12rx/L+jnqIiLjise8JJVuwF0k484p92TjfArU/o4y5g/LwH
Xpaul6VCNfT6C5fmG7M7yMR1TT4IN/iC7GTawieyhGeMNOjrqpUn8AIRL7zj
vzObLAzzKKhNPTWRU7I63unjjZLeZjZ9T5kWW0/tntwf4CGhK7yqTxTzq/84
Aje37wmom8ZOWIPS1HvZciAz0YsDUwTSA2hbdJVL3phFjsaQnrqN4OIGf86j
9AUGQ+ohBgF9I63x2SFst32fS78dO/FPdH/td/kBsrMMUNCb6d2Q50tNmnsa
Dzngsija0f13Q3cGdilrHIL7AyaiSon733fpVBhBCGYr/4SWi76P+/iBoDWv
HCc7A74guQ27uuEg4OjyT8NQEGZ6QOhCU7LZJxwYUcXAQPZcqW2gEPi/hhwf
0Fi5Kx3plueOjSrMYKxIzlGdQfXNL972omcDJD62Y2R1iYJiV9i/6o0JRlgc
bQV2tiJuERSngGJS4OvAHoKazr9R3n1OK/j+18m3PQ37PS6WrWYoianNAoO/
QDWKMYUxpYasvSErl8gqJDQnM65B0Yf8dOEANSDHxXaeiG8FOhSUC9hvCuf2
wAVw5eqMhEY1lmMghO0JTWqY3c/ijRgJlZ2+dwBUvxRgOqn5ta1vNaL9eI5T
c+xWyp+p9DkhCzEh3WJ8cODtvh74wthg1hdF2d+9PERGrxu2ZPVLqU3B4Mk4
0SWVDafA6DQxCyHz2oweuzFQL/BGZYqxvVdVCp1kIuBkJNjfCxeiejQRyzSJ
oSuv91C6M9YW5MeGyHY+EICHGs1wHkW4YEd7tqFlDYreLjbzt59FUC9m6j8H
ootxaqbPpgzr0qTMiIK4PUXYLpbfsdCwfApamFfQ5tmCwyEwa5Aqy4txbwwG
xnubsRAdMk6jlVHXn6rg3LrICpjBYtZEHssWklFsxSfxuGtW36CLUplp7CiD
5uu4RmDUyqbK5gF7V3hSe5Ck/CxtAASXrauhivYNUJQMb6iC1Q8PvnPi/Ii3
Lx/WyGufkrBi0SzYSUxUfa7cfMcsaQiNpsNYrv4i0aYazSEaGMnTCpc3VFKT
majQwk1Udw/ydsPqacJaaKze4Umtcgs2Tvl0IYjFptgVnAuSx1367cAwjdSa
wQj8k+MH2DjuuMnLSKYJG7SNNFpzfmCgt7EDBW9fUBxf3R+FYanbtOb9k1+O
5EhRud6EfWikPx/BdLLGALUVSxJVip1lblpIzINCTMITWcfhApbJDNwqpevt
7UXlwyJB+zbwYqyxzBpUXUjDU4QugwhYohekzLX/ZwAcam9xyUFfRtpDiXEQ
o2FhsGTjqK741V3nHOx863zxypAur0KNl+/Eqd7ltPzQAAdRMQYagwbQHLpn
za4rdH/bGIUlVtC5mp4XGe073cDHbkXTRLfN0hyyiHCXgSY8fls3D6PxdjfJ
9tdMlRfpxAQoGr4vLHJ6/e3hPZhwXPONT0xnQ6hwoSI3xlLftwoSzFTvX+Qg
6Vjni+kZP7SULU+gMMLcyr+9GSU51DR3AXAITruOH9MI7NF0q6nh0+m39MyZ
6hINBWZA1fdDSrx1vQLL2JwPR0vOXDP84Mlzm7yGfEZRt0O/QaJ4Z9fHLVvO
bM3EpSVhsAXdCW6fXh+9k+TB26OMsm3GRemS+cWvSTy+Oi7aR89B2mvKJ7Ru
lN+6j9REcEKb2Dwqnpn1Ai4sYAky7YO1vc139NPbFFOkTmWthOjWnPIPEFtJ
h52YGMf7SVdaA6n4/fViES7YA9oc5KHEeDIe6xVkqpH01klGiQLBOEBpIYsv
8GpaE1fL+8YjVtbkyA6Emfs+XsMhB48AORPaF9ICvylRyBgWeDmt4z1k/xhG
3HEaTMuvTy6N3bVK1Pkc1L4rj36qBmodIoXUwTiiH/3rw3sz/tkG6ohovc8t
g/o4Fg61qZ8UogmuUHTCc5yi2lE84TCDT4EvoYZxCDZQngvCIsX5aHp2vvgh
WCZcBxZiW0rF3WR0CP++1HDq4NMh8OwOD2nNkl4O8lf+9H2K6G19hhglSQh+
3Rf8TmGvlVGGJAFeIWAKhl80yw/kpcBAvZKxpNLYpblsECV/fsbHlaw62mJt
LPoW72v884dbxL0j2+S29qZMkcf7QFwO3GcS86xcAIIUqxnTMdhpsFN/EeST
Al1KXsRvXW+FPNLkP+2EbV6OYeyxt7f+83JqAW0MB/t44oUbF9cL9hEqjTX5
prbELvJag+z1qDw/RWgQomfk9/wsb3xzfXNxYXMkDnyOZOEq1fYBYFq2Mqfu
5naKLCoAhvKQxYDp9gj6PDtRwi4KXsZNU9yf+i3sGtTQ85ty8Ki88kk4Yu4p
ALjp56QqzbJwsfmvGODIsyVnfQVHKiL76eK6qRQZD/u0rxIp/xH8QD3lU1V1
Pw0tgDzvGdfriGhKqxb38wnFRUXpIKx/UfijjsGPYGMuM8zEquoE4v7JDA+i
bsEakdaC11gWsM7YB7RkSswyxSjCQ4M//B+ZH1bE5jK2dCGqFasAQeHcwfST
YC9nDA5ciXAY2O86+GlCdSY3cyrp86OzAq8U63/tC7NdpLERY007CLw0S2cv
SqKFMBm8kOzOOHDEVNb9zzoPkOkR713KvNVYZkyHz/dbJcZov9pfooPdu587
SYuqmNZ4MeyU+5XzoMIj03lmbcfVvfvKnZM86RR4RyfzuwpHf8g47yyQTVpw
ObzaM8eli7W5UcsmFk20W+eQjR1rOo74UB30v/v6z/xZffNuCtxGgq3gDvsN
i1WL3kVr7nIlizLjT9CZl7mZBWylwREoImkvPDIy3p4Ves/S4cEBTOogz1p6
sF3k9KuWBUCWrg+hbWg/R3vhU5Z//h03qNo99pepoJYYbUFNPc/m+Wt3nlnA
mAb2mpG8O+NVRj2iAtvF/PlEKKOVF21jFN/C5CLr45GHtLBukgPkRXTM88Cn
syz6DampcxgGVENo7Kn4SniQawGwmpSElGCCV/bh30/XZ31jY3tWZNTLKc6B
j9oOyWtBC5yUD5NjWYllgEwhqDOkn3AVVfepCRpjlhFsOcKLS86djRwaZcKy
zMF3mwjnQEhVSooG/jAGCIF0dZsnWt3WB9UOwPIt9zTlbUYIq17RY2btYuqJ
fyEeoM0miUPwBAxHrZbAwBpA9Eb49/W1Ddzj+HRaYxahl5qBxNbk8WIMGErX
nkE131LNdJgc4uysODSEPBW1Bq5Ho17CBJvCB0fRnzcJrikOQnbBTHcvAuul
+Z/PJ9ON7uuwO7Lq8T0ebohva7ZULfr6lr2++Ih8QVBzwEuHqW0+qSD0erzJ
Yea9OOghUDRzqly1YI+u2GV33naJhTsqfZBLtitHrw3zCSPYw+bhbCLIm766
pN9MvqAANUg1GnXZTREDSfV7lyZytIauYoQx1T0wmxoXJ+WWL4bRPjn65jTv
oRNe555kMXqcYvRkWxzEYg6YFjWxJH8zOx4tSBqNzoXVoparP6QHn2uW6A8u
dCn+yZUCV6QyS93M53/emRFjJvW01+kMN/S1G7EN6uFTXPpxip4uE2+JUlac
CVBchRJAJUZSiYYQ0b2Bx+emNbvNbzEdUr9mKGEOTi+qngO0M0PpIoJrmM9B
Ca72SIU3I5ywDEUxSHA7y/nZTwcz0G7CuLPJrtTNL87N53MIFwLhvlrRrBfJ
6nOgPKDQ16rVW1vTMLGitNS8dildQbCb6xcV6N6xZ+EV9eSJCWasaHoEB6XC
6ctPJBuwRMIVdxLxdqmfkx4qsFl1HW1MHTv9Z6DCqxQkcpKj6XGvWxvgrRaX
ce3/j0uuhQx3/NA6Rek2Nu7p89PDYLYwSj9YdGEInPVp841EsiQaNskVBduR
8nRD7tY7Icio8nRGCQBDPOMIOz/sFzA2M2BIctS1X+DG0bqvDvuMRs9QNqop
7jFlR1JTiWowBulOiy55g+CuAG5aKp8kmdVfiEwQaphzz8Qt34vL3q1IbXru
wPWv/3daMvSRItGXHppFW0SK8UcKgf+14/ACI5jwLx7hrL2k97t8Xj0hNQ8H
359HEdNRbN2O6bp2wVH4fCv2b/zMEpkHNZfQNRQtfule+qLKqUvz3fUilM6a
Lok6FOwe2+P5RBjsyr0amZrc9yLb4qA5EOBGNebMBjhm2RrMCwPotB+uMLov
SVPUtfRXxsJF2TPLmETzLB94aVNN/UL8VwCDnYIPgpVQgXPlERIJww4owIE/
hYKo1h/sVfJDIrRHNLiihLmZlgZ8eAKhamZHqsZqXxcRcVKR9oU1poko2z1X
0V2ks/i1QAFygGL2faQgv8nAVhyLnk4dQF4bi/60MvIHbhE4oIIwkiGeaa+4
z+IEVw5JUZ3/JsCgcfuxJu1vnvBVwUEZwiLIYtfqqlUaG5dB9GOox5JdrjSB
SORZYYaVTunqtNcd0OyyUAP3wyiujC4d05avGVQ+Qw2LPKqLNTrCzj/++b4t
/5m5j/SHuW3EagMFcoP4IOWZeFkOSTfDqBlONWlBzQCPpE9002Hd4AUTdRE6
3IBR3kAJi6uOgg1gVhuGM8YOvKJpbDaE65vVQnPHKQypazs0zS3I5rOOx24m
OKoP5zmvURsjUh6ELEmChdr/oiTliEMXrEWI072YkfS2+9sE3T4HrubZ7Tm0
pSD5V3c/yj/SRM28RCdn/vJ42anP7KGMc8nmWM8te5LnehykFb02YQXLoeVm
FF8K9ceL1iTRMzbtgiJ79eLm/7C0AofGCoSHlDq2YcfacBusU+LellpKCTTO
TRxTARjWmMqpspGDB1r9H3+R2USgKjrF/vRvG30S++g4tdtN7n5KLuQ8QDSC
sVNNvMWJhd4+T677taJGLFWGTqsa7ysICwhVftgXmehE4eY4rAVXajGu0fy1
+unfHbLqSDr5SXpaWRW5+k3XM7aq+7w0v7r3GekT6I/EN7d0AYCXS1u2GUzW
5HhB2GCoqX4bErs9qfy2lwbOm8he7RiYjEro1BILYqdFA+tr0bTcsWov5z96
nm9LyRHX1wFuOKu/fO7fX1zYDLrL5EFJfaD/PtpRvmadvBwKLtoQ5iuEEAO4
ou2bV7iJIoBSMatFs1LnRPBBPLanylleeFlM8lMdOhgZwEvZ/cAqFNCM54+u
JGW5tszcccspsqAMocukKz5qEK189Ia8JCkd6UPMnY5BpP9qUzEQVA7FuyJa
ed6TGkKOQ1SvmXqsRVIWq6hXZy4jYy5s9VObTA/eu4mGki2tUcEqBJpNLVfd
s2GtuUqMwk2iG8n8sBlfGBnN1AjAgouDjceDG4tVdgaONNlCEEWOuXNz3BT2
eY7HKh+3siDWJtw+RhBUv/BJkn8asmf4Kuvq69eacFEeem6L1BQRlBc2gzU2
k6OiglKbpVna/X5FfusFHU9dd/Kp0GYPUj6WqWE8ngOuBBhs8VJwhLsk51ca
1fNbCiSYq9q2xhlXkHjPAcjpH0rO0pguXMoi1UyIgRiMnEC6Z8oZArv2vtCI
6NeKbONJuAjxydBlAIUZCSj84OZcULY5b6ik7LFu8JOjRi1n0O7dH1PHa06C
lfrOvCWqw1vXxZeo3hBnVJGpIYgVHwQQ5RxbL3quoE5adRd7AVYgwUvMcsOf
LOnjlWlAeY/5u6718/AIEmjEkSXV61kqrqIEIvwXXWtyXTvQYcc8omaRUYLP
v7zhoRHp8dAeKsQ0LxM7nGbzHOI9j2F41OxpWW90TwWebV/JcRbBrGiJ546N
JtqV2v4dfX9c+Tx73HqFMYnN2u/CkvKXK6lF/UhFPeBHsjAy6qRb2jGFwMMa
AyVmx8sauggj7/1KWIEDfJKJOC6FiGUK8irMKX4W5qe61fZR7KqlwKreVf40
7Glgu3gYezh2fExLYW5HHC/Rs4VZuELNr7aPIAjjrq5TAnQMyaajrTO0eoX3
VquAr9RT4Rup+d7LiK65YQtbJKg4bqZr4v/W8n64ZcbHcnu2M0nH4oVpsT3x
zFb4N2SIrjygAVJXqNeru5RehGVNjRZ5Merq7XS1GRjVBHslQbBXm2AHktCA
pjiv0U2QLiH7WTyXz+QANyQm7JzYjpdBKZdP+hjFx72pTvZIkUk2Rm570/1M
Gso6h4vxjgcSaWdNMjmXfQQHYqOFCce5Cj5GgJigFXvE5TynmLcs9/yQNdDW
63L837xdIW9/9/XWE9nJd83hJSgJxeVnFFf3PpQ2H7KGa4zLoQtdY90CvWoV
a3YZV198c6vvW5POczRc7OYHDW43qXYtB4F1prikJZTW/DGvT0HAp8Javd27
FR9ztxrum3gj2KomCkrc476qpIV4TCc/JkVAaMT/tBWxXBgknl3agIvtYC2l
gy84WYkWnHXLkenW7LP2M2y0XMxR2vdSu7FYwQ0cJE3lxvwVCDzIUUDBDcUP
tDx7+d6/bu57wKmDCDU4xn6WhQzLzcvgJFD5kK2M2U9y2so0LNzHBHWy4A1g
1iU/usxGJPLw38e31NM+Y4L4wlA7tht8qnYNGX5bXXUqbXsGTcFRZLa9l0Ce
UIUUX4Hfd4yHUkN3BZgMkmEegeo5iadd5C8rPohmqHuHFc5bOEME8hpWX8xp
4wwsQOX6b6jweAaHRMH+nNe4BzaBx0WWs0IbtCAhsOdkCAqZXXPlpioPgE4Q
dLYFl9erfhzoVRj2UCIX23rBGLksS2mePulnvydnlgGa+kC38MJyiABwMDV2
y7oECYgOK6j+ZwvBMQ0S0JpYjhLz+7E8pJ9jnLjzukM1PthN4t1qGV0f5+4u
MMH1bboXuOIukUMOlpvOyWeoRF9f0VIxw048RITOe2PHYOxGuwoykpXHs84F
bJJIqPaqy0Z0Wv7D4mShchP5+6A9GWYLMV0NIzRiJ+eGJUxbzrjbSJHkdWTr
vMgptYGuh4LQuQZTkdmY4jjxUMyiTAxnbqo2TxKJNgUDzB7n5soHwuNoCzAd
lwBprqFkE2I6PQb1xdRcehdy2vExcaOy6w7j/El00fi5BnsyT3iyA7mUNXUd
kaolfLuO4R5bqlh50nQThHpzQaIyEe9Wyz5DtW9b2i5qw8Adl4yBO7I6K7qz
zyHv1km7vI7YY1vdrl9NDm0IuyPf1cLvF0hLguZqyykaY4buzcwVDgI7EUN7
mNLrwsMFoLhCMTwbJEv06VM1yjd5pWBlaP5533K1rowNauIqRGjHy6Ejuaz/
46hnbDwt5FkpZCDp+S30208ER3Ue0X7dM5Kh0it/S1QQAIaOSaJZ1rHnwj9g
iG/3syAxqJGrnVxi8TGg9MnjXcY13oa2WH9kUZ0bu1FGjugdtQxgSPI4VEOm
2Y48dBr/O3qkqRR4bxLrYW2V+14StIc2ljn1HXmdXsPuLbBLEKj1GJm6k9dD
wxMG3ewTqOgEiE3FTpzK1ry75xb5aEmrYEnh0x97Hh4k5cR2ES2jVodg31kt
r9aWT0PLq9LpnrW/PVtUGfus31hlzNvpsyMFa5DlZ+EOnEa14MnjCj1sX+cN
voCUdGUi7/KsSAnUCzj43xLk3u5ZkGcOmj4LVbpqbeI9/l0AvXEZ1QA9HOAw
gljQweCTYueNeYGw5ihVyofb5IXBVo7+P6ih6CcCvXkxJFQ7wSE85IMaO559
3LjmNG9RyX4+mw/OszY26iif/OFS7wH+Y8kHnDAYolJqZvWM+R4QztfHjcCs
2TrOqSpBQhfGbWrM4ARdC/esWwNMXteUvVaKNf/anM471/xM0N/Ca7WA3Vn5
rCvV5pd2GVpOOfch4VBb/8eK254kEbCF9h5szLPHqEsB+0f+vTAycfAyl6Ba
yqMyjmHz5HNzJIKNJmS+gbaFqHOLmhw060oLgBqrdZMyWwC6UH6x9qxz/9Mt
xTF/Omd8SDUe4hWYZXpqEiwi+XLzePWq2ApHx6HHMBH9AwXADcGgFqUZpLCt
KtXmyeEuP/AaygMS1l/AY0vIT23SofW5nrezkNv5RwlcilSbnHfCk5sGptsj
E5IhZwOh8wMP+4r8Gi29MjBCDf3ZNMqjgneiyz6P9MsmzvvAqYyeKtHY/dsk
tOMj7TVF206WFST+SMcBNH/BNgT4mPtN6cvQhs1ViNEFdUca1CXpMjp/X8mn
0Wh5RoDOtbdTqLC5E9TmM4Fot+nbJzZqKxk40XSnnQN2a01KBW4hrM4s9TIh
0z7g6xAvOfmiziWrc7SLyCNdCnABHNEcsqZ58iwuAQ62fJObCkzgIDuiCUIY
GpLsIPhhNfOpx24q51avtL67Z2/fv4Jo42ZjrjNPt1j5byB+n6P9xTdxr59L
f6RQtS8XHAWP+J+pcaAreAY3mXlWL1b32uNgF6Jvr8WkqOMpq+zlSHuV7WeA
xDdI8ikaAcJCkhI4uS9gmJH0H2/nOzWL7tqLHamsvNTbGTPei/LOO3GKlexd
HnuETYVLod6trZTwieehqrnm1uQEPme3NUgOvi6no9n+YLHlnneDlqx9rrDa
E1137kevoUTiHtgoDsm5Z/9c6Myde1Hr8BjsbB+K9RVVRgGjItX7s8W1rtGd
O2AMvt1ByVI+uEJdLH7szXMfXAJVCojK/VQxGKNkrCpQMuu756cyfuFeFtFI
HisuJrnIWGcycUL3HD1PmeQtYU+K+GvheqWmHNlb0pK5lt1h0ec45cSlYb5i
7A2Uz3AVqrYdCE7w/J3O5eKNlCqjnWe1aNCQ7xMDbOtXsrm0eR8Kosske1BC
numwk8/JgDxwMQ6ULdTHucU7s7egHwaLO00XYSxObJpmryMChKsRPyqElArc
Zn0n6Hs8V0rGTcfNdDzLiMTKZVyksq/b1ZlrYmNz7spH7jJdE53reOdqiHmE
+023eucBo8G95bLYYFYXR+BQq6BzXuHAYKbcYNSPOxkFH9/4mupafdijIJYz
yCdoOyBInjmoOjJzsZGZzQU1Pk0Z7l8Q+h6RKj4RzgQfbQ+9EzGHahOYrfSu
zeCNy8yBW+rJMjMKoICazAJfVT7EmS1nFp42p0HWlFv77n+sOToJgja4jyOF
bhPVZzrrNpw8oJcDSFeb+oW2yGH1HdmXYEPMCIWnjDMVJQKlYNjxjUi33COt
GvnlgDzg+eXLEQL/FrUIvpQkJpz0nanlgU0hNf0hWvbxKXAgjotfKi7wZhbK
wl3TieQmY5mxWUg+J9YPi3GzwgbiqmMb3trv3VSHksLjJxrZPDtBiOCeiqY7
AaZ3Ekmccj1/gYMcwsmwGPCc24g/EylxS/++sEUA7ALaV9Tl4Y7M2CcCNou8
1fiW+N5M8uof/XBbzXqbTjKbAhDGOfC1/QtuHjsG7HM4W/x8iwTXuf2wDAkG
9BtseHsV13OmnM0CVlVC0XQq5lBJNtK5QVJtDoljQLpn3IAQ6RgAxmcP+/jN
UnBmHm40+fLwWqAi7eUjF/Zxp1veIzQTSlVpLp3GFAZ76lRohnb/YpA+115a
aPcSCIXDmnPYfzXTCgLBeLT54eXHAOXR/kUmwxfnMD3V3QtbBdzNie9UkubR
GirtKkXRDtyrE32OIBkkbeLztnv9jntAeTAywbeeyrXSSNzZbiWueG4NUTFr
4lChxkEyVl7jU6NqFI2TVGDgk/+v7yjAl6/Vtv16/nsb9FTb61RwNwR6v2t5
cak1s3VMszqMdwuLzIoI20+q8EYGfwKgBhH4sQLGwlHkesJ6ZqfJOx2EJZbC
0Mv6Kt2gyCFTsGmP+bMcdy8HwXM6RARaHSgCmPdWeKCy0FBIhbjCZ4HZ9snr
uyiPmzPFgC3FOoMdXkB+QeeyFQAuUhpIQj41F+CSoDCcxp58NTuOHJa2JPWg
JmZfeUbhDnyYOdGd5YzjScdYZJJX8hPOUMtuh53cNxp0LoqHKq/6crVYK+93
v8BSi5rFl3EcrdeFJgWo0zCBx4LCwXewfSIOCCZ+Uy/LHQ3myG6qRGINy12t
1hr5RJbuLfWoOSo6R7AotkpF7l8YyTlHfdOdhsoGJNw1MKDHXfRTjzyxKmq7
G7HpIduosTh5YGFh80f5QCXtZTeuIdlGaC/IDEs0XOnM0hyC9x6uFXJrbobY
XLAFhg+N0XXOwNMywNS9RxeKALcFS3lgqX5n4qWRh+ukWTIYuFYaI6TW36px
8mS/WdG7n7rLmFEN29bu0s9L5Uyq6N6dZrNLHaSxhsir3pOg0Z6raIN1TcC4
Z4JqZrfuCwFo01s6c3fKqz7dZ1nrhaSGBzYCU4MYWJsE5zhBgj2nkEWp0HvA
OxX0Xa+5YFD6PNOvIYI68v6VttiNek9axAiUcC7McrnfLpsICk9o6Uo+x46H
atKqekJj0ZNxAgHRanPYofTmZjErQ4NsVeN88837fvp8Jk0/PJc/2quMM6pe
+eLC2TO0dgiqgl3TosdXklToLf7rKcyEQjwOZpMiH8A2YMu11JWi+a8veN59
GYjNN6E0f7EV/4FM3pf39YTthj7WRFzksy34VZUf1OKJGSnIH6l91h9hsWpz
8R5o6AkC0yCJNBNjz5Zy1cyNfAJFsJM1yIz2ez+pkTlSziCV39cMZkZa/g+x
ZkkcAUk5DfTX4i6V/CNAPYE4bcQbrLMF6EYyBHz6FWfQIZSB/pLFPmb7bzJR
h3gJyV8RC1o9aN+dYC39icHtbetsOOjcu68+8XYbXwSYJ8Oof04sqH6xqXD8
EKRzRgX84KoLsnUclSBpfp0Wl3zhuavUr1qWvf8NxJ+eG5Ylgae8OFSF8MER
m86XVWoUiOrdS/u0s93pCDpSeLtHaQO7rVuV3yE5v0wDNS3rf13gIMfMX3Wx
bDIvjYSdzIhAJfk0gTRuhgbd5wHPa4TmKXvLkBfegfhu1JtQfDoGuPiYzGlA
dcWjJ0ejESTCLC8j4IqanW2UJIwj79FqyGbQ/CdlsbQao9SudWkSE5C9fcVx
6zfqzbvqgCtCvwnX7tnlC0nFVKRkiPBfBVdEsWtr+UlWAc1I9jMnKXWm1pYH
022gfpIie/chjd/3blVMPhNOMUxEc/WB9azn+K5FNwSmcsXIdENbrQOkyfG7
ms2rBO9JfERAPd4ZN3Nuc8zmh0kkT7109X/ktDRdWYehUOrGUog3DOZSYbGJ
5bip2bS7eu4OMVt2cqosngxzB22MldKxRTcBiTNb0OaWGks5AOACr1RzpSHl
PN9+ot1YWr7qK4m83KvG/DBBVrNVq+uDxnQXXDWQlwqoyghk087acLh+eC6Q
scpSP1UvGYVVqkBqaFY2iGsoLTNBDawOuJ+A/bBNX6UAJYv1woAU38hcMrfq
BO+b5daI0lUtZMRrtDMny4G6HxSv3i17tI0PX1ZzVvS9mwEEF1AD7a+Bgsva
it+Q1Ijvq3X7OjfscZCChlYrpeG39g38B0PhV2+QTeSWPaK81SPfk2xgGCHZ
dXEwEz9F3LGYNxfIdt33w0AKTwQ/GcYYAaOVdTDpQQmmmiQSQwP0uEqDIXr6
DOcjZRN9DW5BU6/w6LfRpgv3ek/cPbQgoWG2CPr4cR6Rz+47NMIDNpsQlX2l
iT9EEqSVBY+BuN/kobXRtBaIKt6VzO7q4KgcNbbqAQaNhi747arXQjsAhcZZ
SodvxVQzq3RkHwpR0JljACVaHWrWw3PgDdatWHR/rkpMtOWxCqBPuSqNPDrS
ih7b9y9VmWP16oqQefgC8xLxF9VyqcgO4axHw6eP/e0X7EoCxuH4mjOF5+lI
lhZAUDGlrcvsKKo1Rrcn4VMTENMMZyVZh1kZVfhNoctQ/iXUMoIloUOKhwwH
vOZ37yc4YZj5xWQEoRDV3zyeAEW1EyF6EzxZLzUwnKLMpRZf9qxa5bsgDw8E
pn7hBfs09alwh5eNKs0V9mCLsZzedmjzjDEkQl/AVTaBL8wBJf16a/b1aBwK
40jkmg5j4ra71pnlfJbPYCOOKFmRlBO5XENsy9BfqqQSdHi+ES9A5qM00y0s
AwdrJRRGW/NQktYK0+m6rOieWNFGNbTSd7F6+xqEg4Qn0ePgVJTYMppvrGSq
6RYzqpy8tkVQrKKvTvzS9kPAGBK6UgQ+fCV1KK88BvxvDpgRb44v8yqTvEEk
ta0KLkwlfZbYuybAmsgoGBzx7jxIJ9vs8rxOXVEwugVSATqHt0JAifK/9YQS
V3MzVRWd0/VUvqYp9sQxAYmSrBenNorHuYr1xa9W8g6XkXKQnVF31Lz1Kt8F
IRlhykFrO3oq186Ei+grSQDvO7HHr6KFU6ND65jXkV5p6X6QJeZVzO/WkTTR
yMEBTcqX0H9cdj4GDPs8M3I1IR7pqq3/j2368LaeZmfzXegyTi3BKMBWVNk3
YDXCQ7mygpSj4w7ZniK1A7aBcVYvwI17gD7vETySS20YDCGJsjpvQeedYLVi
GT/Mebf+P96ouZmfMbv+e9xvf5FKxZpd0iRYQaHe3Fn6Zb/3spaRQZ2cbAd9
e6DRK/npsItUHjkIevb52X4d7gotuLD2LNUyQczRtPZ4VxdMKstlO9z51EOU
lu+A6kWr/ydvGMSx4EOejvwWF5ZplR8K2MYI+YhFozI4Co2jsyJyx2GT4Xod
uYD7WytO+fLBWUUyPznzjwynxk3x1CxAWynoX8gpClGV1KAXrUzxyOpz33gD
gFNY+azawb0EF6jdJ6tZmA8FwHM2X/PsDbtTCEyJ5DsR2HR2glka4cbQ7BZX
UwXpceQdTIdqhzRAkN7YUz+5uKSJBQJaq4CUFql7Kd6a1gUf0YwfyINzSqt7
hKhxivqnwAU0zIvcVSYsmQaxqXLRgb2Zz4qxnzsTO/NOGPU5faBpbccpCS88
ct2S5ZSlMmN+HTlEF3b5/OaHP+kVsdQmrxSgbpzhFLc30kLYWMDqCjkR7fiU
pCQ1rSGSMgsKSAOTBvZ2s9f1qMqMjaLzsEz/h4FLmfS9QfPZR1xykJ9ybJG7
CWbt7jX85+61ilgfJqRa7F7/UznwgG3FgWGdFrrNZnq0fGXLBjH2FBuWLh4K
T2MLerFYOTqwFp9twkFUBarjejU3uvXjP1sC6eGhMYsaadb3cN4nrORJMKRm
ovVapUchKR1E+9nzxWB/+3T1xkGDuM1rwFJr98at86qZ9fUKQoj9kUvCmngW
WqfoBuB9gcCwUkLAWAevmDF2jzhgTszFSmMjOzmtnGHdSN+AxfrDohoxZgF5
LQJ1PqvAWHzosOvcTJ6mLEmiYuOBA80z5jhZarkW//Iag+b7AieVWJ42U1LN
ohN55ypekBj/jRKJ3t+HaDkcxEVX43m+8lA6ekhqV27xOPdX4/dNVcxzPSnN
0Z9Y8BIaOFfVltpE3nNQfD0dWOTeU/NC8wLwueRp0WtwEvW0iVuQgme2eloH
NmTHpD1yA5wCCjJitQiHBqwpAEnpLtUdZzNWh3s1OI8EH5OIPtPWg4Ei1i0x
KEUaFFQLQQFgBNZ7zRBvTjtJDZK//P97uMRtOeeURccGz/XT/JXsC1qpo7xd
LRGntOeC6ZR9gTa1fcSJ4Ubjeiw7aNtKsxKiQCrXV9t2JpZaOu6z/Hs5CJ8J
G6+q9V+57HaBz9Df13379A+jsiNp9DEdu1wMGEkPHfiXpRoHp8W1K+yKICZ1
TzxlZ5FkwcvRNqal6Np6na94dvqm6Tzi/Ab0/Kmbb1hlCqM/b25sXgk6lWrl
HICdcAIv7MAct2/yqrecQ9h5qPwe8kpv+ZQl5jnO37a47Q9lhAtb+8PO1F39
JOjcUWax3OxaDuJ0fsofkZL3iIHWJ4+m2G/ftsjGpRnkxaHEx/40lS4ekIpy
7A2hENpmPzOda8sHTYwVzTp+FnjgIdXhpqu3Lt6LJk/j6/NL9+fseG+EIH/W
qxLF6hEjzcRtLJiJ64RkbeQKVeBISuvd5FUDd5aYAZNxTNZOhG11vA6JIFBD
0G4gE0CJDfvV3Tyfev03lZfFdWkTf/YSuHfRdxcbyy94+Pc/XV0KD7Uy1peO
NCQOrArmWAnPUe9Qme+qesmyrxzAalFiZV2i3fvLFUX0DGNK6QFifrPcrhNQ
sYQqlswIxx2H6V6Yo3nRHR+Lip7jWc0eiR+2eycix9ygksKSQUDpYzURe2HS
v06irtCCLIJCgS6lgU8+DQ1uKcrBG9VC2K7UEMo+U9yAGhP6KxvpM5FofGAA
cDjDQqQgLbqTCnIhE1R6DGyFog1NLLHJhyqyZeMNXTTswECnahw8G0EL5hAR
ZtTuKPvAQZ8OlHCzE25mUTQB1i0qSEShN0DTBqUSWsmE2MYjmj8kL9ItvZVj
gYoZ4egg0IRVQGZnidAYUy1wg6ZsraGym5f/G/+icg3rAaDjJbHaA24/sbNQ
Ij4LQKStb9Rx5caK7OO3UX4SRqFRCL/zsIt5cqaVEA3Kp5ewuGoHZFfQQREE
/awPRs4nt2sBIXVYYoYpgnjChpC2UXOTgwUoNypspNx8NQMQuPNAGGLw5EO+
7FYNnCDE+yRqxe/CukE44aH+mYQyu8SnwXb5xC3XbyIEm50NuWqrVRX9KVDs
faMc0tbwRaa+0qz7Eeu8PWiQaBZejWYOFDQOoG4tBH25uopfqFsz3ZaFpN+V
M4OCxDa5y9NlcRofgF5TXIL2IqX0zE5yyiBWD6Kc4EW1GHeFDKz2VPAjWanB
pSsG3jdAvaxVilwhP9U2mDGVdk0a2yO3aju63b07qPBMzCYjrLYIHfmeR0wV
jHc7YzTK/QhxIvorwmcCkzb7DHAuehT4hciM+cw21ej9OtDCnZ6vxewE/G/M
zTENlDgpYXh1OnT4OcG+RLFUV2x/gX1O0xJ1boWHWeyCjrnxNTm1J4ycrOHH
JcLi9XCxIy3Uk1n2QZrZpSmfV0xIPnZA4I7F9CHZvJ/F8RM2v5DFBARgnDkY
DmrD/2JAZRdI4vcnfIrlnYanSvKsOvFAF2wxXAJMWKey8Dj1p7kCgVooCLrR
rQkqWNZBQ8OzQhU+hOHaIoILJjTRHZHWfcfA3tck2Ma8ZldTV6DhgEYSqUd9
BkaDIWB/QGGHWqRtGDEddXDYYaporJDGP5LhsRPxJ+hEXjEFeRnfhiMgmuGs
mWPpDpugOZVjYkBTvtouUdBxp77YpX5bh4B2sQasuV46gFleCtOYIxJkj85K
UbxOR1pF5iwWKm/BRVEBo7FyuhWCeJ0TO29e4xZNDs0+wDjCW0xO/tDSaLvE
lnSlQgA/ooBTT9XEHr4c/36LssXWcbKuC+DEp5Dajs3+U3aydN4cWXjDNH8A
W7QB8Su3Sgn62CEvyG6uErGk/yUQVdFt4Bd/qCPsVUeztPQcsHeRowGL9p+U
1A+6sWyR1+kxiWPdg2VMun9u9pyeQ7YDpCCovIdC4y+IjeFIdf08kRd0oG8i
7cRQP09wesSaPzzH5sU+L0s2piw2yMjfVvA1u3ly5ninIMK6Tm90yhRBz2ps
3vtDahzLOjUyg2rhZLe43YqZbq4sAGSlx4NqmYd1vBg/l1J2Y8xP8R9ucyuz
IfzJfDa9vtGyrw0H61oNKUUjDS4YLeAAEibHGXrnPmRSoVzCuOombxSrK1Zm
MiK46A3XQLEqmZ121mZZZDOqB0sKRX5Ifwa/sSWv8DlhrK3gbdcT9zQuRVJl
BIhZNx9T6rTFSQem9YAn7Lk+UiBN2VpRaXahiEojzRaZCViFnRJC4nH5lWL6
NeGtckveRn6OnhyA0RgrmDSZe6gqg8u9/b9UuWKaMNPZeKo7kVCSHG/0U85r
SfPKc+UcNtRjjKWI4f7kkpo65yWyngJwJvie3O0ukFd92PlOf3SKSe4xv4Nf
4Xxv2A+HO08qqUyl6QzcgRloNivDeYj5f/zPplfrowf5ivgbk2nPFyGkF04o
QqGA7V8H+f4fsrehMSDZIKx3Rqj15xL9krBV1NBLsFgNd9V5Dwli87lUI8Ia
ZEoFp4vgS8BaVFeZQiWHUVtgmhugVJjABXIPxu24Wu6Q+tmOuMU31AxacQQs
aU2wMTEuLfETDaj3jtWMv15vmCXTqlLpRF3NyUvysmsXX0RhBhUqE8dkKxxq
YtQl/WS0ye4YjVpFZF57mPJ6XR3EgmQB/w5WYg6j8HmJH//z6GQRxUJ6yLZl
LbWnJBcSf3UlTMXyge42JktL7wxTyYn6BILCM5bMGs/62df7a6AsWXCFMwuD
htjDA7KM2Sr9G6pwcHiFHrURYTLxWN20HRzSTFaWdzQLRAb/eIqNmGx4jQJy
BhcVAefS9TPMCfH6X6k6w9OOS3B9Ulo4l3RKY/lUvzr5O8UQkxo3QIMx1aje
zHXKFhL/qShxN9yMiXGvWz/nY59DZEei3VS0G6QeEFYgiYzvH4eI+ymxlXF6
0nnoFDlhaIFMQtX9zNyhv+5PqIh4irrUJndK+wRUx+925LulrlV/xQZcQOLW
lLoMnpa9v/4fSRd4vxxW7vyZgnLY7tttzFnwyV9eUhUdONDcbu5p7jWRPY0K
EPQLZMqTaSc6jGuAN4xZ7WRbN4bIUUQ4sPrallmyxFwNFjC/wsjTUryXfkTX
XL33Yt7gc5ulwJFdsSVEDGzCjlINKB3Ko2U78j+Pk885FBdG2aL9GCW2fm5/
sXTgPx/A0TllYnqPZ1EGFnhWEYNI1igbJsQUYoUXePtbAZfXcEUO2FsaCUwJ
oOGEBYRp5OXyGMlBO8FHsVk+Sn2QXJ37caRBr5E3N80ruXVMVPu1MBFGizYz
0DRj9WM5ysCQz7uDuBdj+3LNdXFuGgHO+QdIa3v3FUvZ782FHyBk51uGE7KI
JOJI9tBwcBsypHrjZJdP3bdwUpbVtEICzJ8rcnXHa2gEzpP6O9NdPgshjhXL
uPH1ZWInM/NKmg1HuddaDFFu+pyUAWpKa1nd/t7iVB7NSTykvgPiNGHdVC3T
e6yvC7jR2OivhcAehuxCvUdQg8FTeka2BAGh7fm+oZiXZUsFM6KBRftDV4hH
otsPr9LlbfH2rGSo+Qf0d64YtDXTu6umJrWGGVShymAFQaYdXc8Gv8MxQEwR
gQCiR6rEAdSd03TlnCRM/NcqUULHXu08EznbXwnB2US6H7Ub0LDg5uRjJYXK
THiE0GMTwK+WC03EK1HFX/NI1MswuscJc688K8c7F5wvf6obsX9pfLGsT6Iz
igVHGnTi/VHwzHZ5fU+oL05l301NNF4CKOyZs9xXbpSHAWW2xRF0h0lufjDd
ctCqb+TxmOY8pCF/sv5cGecd1yOJAmL1skoHzZXYV8UEJ83g07b/n6NXD7Vo
boV9z1+nOtFjLflk735t56JUW2xHvxMKPsWj/nSseVdTx8mOIbeT3LrSOuwh
8brv6pIUCuui3cE5kd+HCAQB87r55sVnNr39jGnpCV8L4De81TrNkKsCk3ub
ggK4+nUyJhAM+hl0nnc6rLROl6/HKaoLdzn/q5hN5zqQk9MrOCDQxeXja0Pk
NI0wMjULjBg5Cuuva06A3Rk8NWGle5W4EUFV/V98/XvrGhlJPQW+Gt6tUI4W
Xpo2AOx4Sqtys4nd08jtQAGbd/ie9tXLf1BmPldnfXpmO+7pCiFacNKERQB1
TGQFw2US2KP8QW+w+1S/UOa5r8DhN2YZ+zEypc7SBChuYFH//KJiHrwn54Ys
fZttj4tkBV5tOQCtirZW56+Xi8qlzkipH+DENtQgcR2SEm9aOXqX4sYXrmoy
mMFc6iRHUvRq5i7lvwBIu+uYzadAoP188yB+4sr89o8lbo8NY4sLeTUwM5Bf
TwDS8J9jmLYil/3sXhzlTQsYgmrWpjbNzn3YDqIOMnlomuZDsH+ATwvWTHz/
8JzvYo54t9DkOR6Y5RlWn/hX0upyuiEBHXwjT3ed4UOCbp2UwPvjdRrwxx11
5rPSNoHywl78VJPCVgeIznpgubMJnkuiGZqJxXtADSoENPyqJcHVpciBR3SC
yz/0o6YBysUFXH6c746nsguupE0IzzzBtZeOaHl/IalZb8mgG2ABMqsEyrnC
n9Chw9AjzOkXMdngSs832gp7XeWXVClbbswSmfLhpCkKLJ/Zm/g5I4SImS53
X+kr3zIdgiVlbW2UKPGc1feiQ64bFW7RodT9IyoyRZZqsFw5ecuE8sZx/RLo
NGhVXR3AH8cBQNKq0yES/z3n3ACsJORGUBs99XJwvFwE1sELYHnNdJF2pvpb
FNtOqd3IYrDUSQy7ZmKdopqmbxMALGf3n+J3/k5Ocb4qhzV7Oq59OlfEjMq+
qodDClzOT4W3jn7XjTEyUEINVKm4liCS22llG31GDKHAeOSrDGJa2Db/C0el
tt40oScBrHBaGSBlSu7x+3nAIfzK3dqgZ5qekeV/Dq6XpzhrJ9/5Ykh6CvZd
aRVbgVHi1SdGuvh+yG7CBA9H8u7qr/9fO6+LIqG9A8btVqAVWB4IP4BuMqoU
bd03jtcPPyIE0ST9XrbM48WH/bhoWJNRf3DYqqk0htma4poAaBISPtGvHgjf
t9IXaZx38jPZt9fYwZxhtO1ZSE79//1lDPMZriKlQdrRPJRNb788RpD2hRh0
c1KG7KvFoUarr05zWTpFUqZ7JMHCfs3zzNFz20j6VTaqVDVOAZYI5EkZU4W3
W4hqoOFENRxO7eaK4GnUJKzZi5S+dTk685NU/s/YlIGYZ1voPB1+fzzm3IlH
vIMZ1byvg3gKNV+UN/HV5IenBBUONTMiyHcsFSEA8bDSVjHQ7BCcrxE08qX0
AwYfISgzjwAaO+4PGp9qzs94+jVqHFkekOx9YoDcciUIs7OssXvUi1wkbx6c
p2vnqwuQ4kE/Mug0y+a6b4vFV/+MvWzl7knvcKeIEQE7c4LpEXFIFq3rYrEI
V/K0MeYMGGATMKhG1PX+jCSZrvMD2C7E7sV/4vLmGRHYSef7z1iXonTW0H2S
619qssEMJ61XVqdMulpit0YI+wIrGTyUtj0nja7wwD672H34KyIBrns5kT9n
0Ud2ijFdtCDbN8XPtR1CLPpK1DhD2ndXFe87CZiO434cBamDwid2j1g7qPrr
bU3+P9DvJW/ieUSc1/CoxnvvUa2PDRpBbjQcMIHyVest93+osF+WZwM0zHXn
eZZxphGP+iCOyP7PZ3gz/2U3nVozOJKVnVZ0j+tT4lblbOBEDzR7GmRj6Gez
Yqtn+tU8ChDdAosIleYrgLyJrFfCTGwhB9uUy+mMJjVvT7AmKr+eGiK2bcSy
DGLpdeh+3cAtPa6fmxFYoFxmGJKe7hG11pAkGwH500tkuqSE9hunH5Ck3BwJ
KZ7uwltm36bkrCbAS/19QjyGiRECiWJstli25KOPJZff9LdO4bHh8d4ClN0i
/ETrM+F4G8p1qcDN/FrmoCPvF6cq/Wh3fueviUSyxQENMfjsKA+ZZd/nsrNn
67sKbcLE9S1oz7eo2MT2hkX6X0AMxiGYnZ0/K9vvOGyEHUchOBHFOgUKQgoq
gO53rFer9hUYXk+uFn9pbvPS50BU4urp+dbu93uXmFM7wSRaAXzRHSKrEfGD
LDY6Fcd4lOccl0XSRKeGaXNPfCA0sVzKgoJ3ObqfaVkGDuH1DrLEGSaY0rn9
SMsUtLhYeUtMgMdJ6sG163YVlM6RHhQv0Mu2rDTyTqJXbzYEtGkEvA+f5mb9
cYZGf48tJ3iVHqDvh6m6aJ4chLg+HIenxwSqSV0xH9D+DEaiAqFQUldm1Hia
fHxLgzwG+4Up+T1L0iAkYzkJhV4KvUYAb4OfQDZ3qcRIRcCIF3qXU2yhaaqq
TWSgfdBv98FaQ12U0egmpPvXnh/5dn3EH7QXhS+GaiPPFt5RQJmGlio+aUdp
FtaXIjgrdtw1xThSgKnpdjLL53hX5jh0KD/FhYevlHoo4OyxdW+Gr1514oil
F8DWmzJMGdSyoRWo8Ui1nvdTIc2kzRavLJuwU89JsZWEzGHfVBBohiI3zbDQ
9OTn5fZZnKMc3MyAXHBpUI37zxp24QJWqw31JGnrnwLfB3QZWTMN4WUdgD+O
vNQ4EieL15CWfkJspcgeA8iKHAmqQMJBa6JGDwKOhIN/NIApVbv1NHn8uZsp
9WPG4/qM5nFqht/Wpv7RUrZmXJB0bAuP6fn7jo0ZbJANvQ4iW0rGuAAhvqKF
yKR3czryG3QFvojHgkczx9ZvoiEFby4fNqEFWLCoPBX02WagGgnVuo4q2PXq
oX+3h0kqM8Z5PphEfAYop2sVqkiWCTzwiAz/HVr0ew6fOFsubBChRT4ZCKsE
0IVgdD4dh/40L/vojyD/8nywMPx4NfeRClErlwY9z0nRGKhinofOC3hDh7iD
wVmnGTO1yawg8M7dIyafwVHpVyo5GbQRe1TCvgU3QVttMFrEFkRbghzA0NyY
zqQ0zIAU2cmdnv2AhGRsnmka8OlOsqXhzxkc1E8TwQDygu75LDPaJCMU4gje
Cju7t8UxJLCxOI/qpnop4VTQUpLnIhnMCHmC2rU5cAgzza9jdv8Yc9AvAMxq
Ur5Bf3IJqAUB5tA7aGLU3p2F1ZWdrLbP2lGbsFaGWK8ynDceFDa2/ZOdkHzs
dT4o4ZVDXqyP4lG0Ul5r+t4ICy1oQinQXkr4z9acPcjbgrk5aabvfw20+vDq
wOQT6MaOBxRHG6T4wIEJHxX4vuVDYxePLzIa0xLc1jl5UCUDs9aLQuujUGiP
EdXBNYeEwtbkJDXf/j5Vix7DKPW8JDGXakW2cFQ+7ii9C0owGVEcBs9egvJA
E2vZbK1aI3mTip5E/hY8SATkDuHXddNMcqUhY0ngaY3ot3HtrsaxBxF0oHPH
waoKB5ko4jvxiAlbQJkNi4Il6EkN5W+L8MwjhsZIuxOrojJbeUy+s3V5mpeJ
qi2ShErX1fTTLJDCwX6g973iCqDPv/57LrPvUNwmDmd47mNEEAnGq6KCMQdp
R8TU2xJIAY8iC/HhVQEc5wjzngkW8NAZgut5OLx1wSVhBl+IT2345IyL/hxs
HJLEQS2EU570spTCvLxR+KtrY5SlqznK8jDBpYP82vZLsEudaqn9le2to55W
E835YER+ZSlvJRlk8wDKbGwIa4McaWcS33Gkwz+HxyADSooq+WSPT8eZtBDg
XvzWi5wv/HJeXjUnw0FezNlJn/XZLY08bSlhEv7CUOF+JBvy3DwvexoLnoTz
Qtx/6qIEEaIBX3tA+eNLUnLWR5PINU5qEPC82hdtDCiaq5usPIKTzrVm7E9B
Ywq94PMsbzMh3gCAioX/gR2Y+k+CYZHQo+kquTaLF7c5vMUW66nGyY9ekZlS
2weQ2FHtzNWtYjxgXyuxt0zjKQ88N9sPI6w4HkD5CY0SXXY9VNGAdgZV2aXQ
Lm8zXC2QmNLeGee4lRbvbe8YLtgg18XNw2bV6BsEa8FvAHFpM9s5ixYuHMT6
ocTuBd5BzvW2PUYNmERAoyhfxgyUU0RIAF/zmuHFOHnIWb2VY9cyZp50yLcK
iQ0xw53Qquz/40yvZY7XvtEfCD41QreLnpS7qqYteREdxIkyNesLNJiTyzXk
pfpbFZ0obgWo5hVVfarCvswUQqNstkQRmDQl8TfyN7FuZn3gZMLubacw2Al3
Q6L7kO+3p7v3wWRV7Yor3oHQVXoQC7ORYWevmEEkHb/GKflBh/8X7gHgswDC
9HrgZuFk8Gnx/fZGkTjYX/4NcaAjak5xT6kPEcHm81bfagL5G5HXQfNvGM+X
xqaJUV6a44GjHNbQGcXS52PpZrBtoXfZixxQB5/MSk0SUQwBbs7gr1BaqzcK
rTLG6xA+feSaR0pndtABVZJG7d+nNJ9akuCQv1E0g6ArLzEpFLnBUcxD7Dsw
DeskQqimxOllEMhvBveCS+UWOoUoAFKBF5ojqoFXAlcq4sKpTyu1V0ymXYST
ulysi6E0FO3HazpknJbB/l5zSS/2qYYHBFFPRAZCMZTWk+x/d/oT8w9RgGeG
LveiDpForaPWB1dpuX4R95KTTSbMtx/GFXrawXOWFbyzfZD/ak7+tqdcFePM
cu8mgHoifST/mAq/j2QwYp+/5M4mZHi4i0J8s9mzV70u4epcBNaLehJyKPxc
4+wejrQIiw1vgpEpcolnJhQbg804BSOiVbB6fQNASrJJOJ6PR2bkyfrgAiG5
waEIIg3o+wNMvT8zncr2wjlDM3jHYZyZ1uzRsKw5/uAMmqcGF0fpBY27umiv
QNZyJkvPR8zEswTSOqhrHB12WZpng8Cb9fSBGOftLT2PC8/7VmR7D28M66Eh
1+Wu3jPwm+OjaFvmHyoWMFgGxkkiqaF6TAIDQAv86CO0EsKyJCdHFvPNQ1o3
hjUuKZH3LaycTqvTtXQ0ocvKhZGyXMBa444lF1Gefm3gTqXkiy/duOWkDKbi
We1RBm9Da70rfCg01nyd0CXAUOjfaeIFzpVQ4OK67nRnRp2nUfbeuQrYzuSy
EH/GUyrdsYQ6jecRqEEJF71QpK7l03c8xWEPJcvfmHODqwXENqjX422Z4eG9
69wqXt/jU2YuqWk+bLjkrO8aMXLqxmgKwY3Fwrq2eyx6/N0FhzotPBt5VkdQ
aJSaGAtrSwtOPvO1Tpcarb3G5buhJyDHunM793+qf3HkfGofmalQ263kivwf
N0Z95xc5I1F2vxk5UzuLvHwesCEGeXRBRgDSNy/TNPujclJxKcbJ18IY8B8Q
FFS4lH9N/h34mqAnfGMkDaRx280QMQB1mOB58LxQE7lKOaExDYZ8d93lYjcI
2JFh3SEzDmf4bD0703RMPqbihABuYi+8jxsveT1oZZ47dfvmsUk1C9Nn1vFE
tMg1RuYP6S5bQzJxc0ZlLjbtw2mthMjnOU6TlvvB24VK5h38BHd8YXOmgTjb
ltdhO9MJzP6OeMYDNom1SioOi3WBPGCXdXlm5KVyNyQt417jNutZziFryO8z
g10Ev3tpnONYdmupyIWAriqhESdwvgAiHd10axaXjIZfJ+A16X4yQDUTFKQa
0lQWVcxC6A8jWWSNk0s0mprgPqVZAwmHSZopaw+la82HaHHVmreb9cre6NUF
hZSoWyxAJW/hXu7kzOJHk3ifSBTDoAhILFrBEJccXBt9tiR6+9BAKiRwc+To
oMgjCEpCzbjJ5j18IXGhaJFbM3+LwxZJyvz5ymgpm7mkfraOcSg6qPyydMs8
tGDU4Rwk1CvnooorItnHlLQF6LMS3mS+3Svfmn++BSSig3nGjvBn6XJrBdAY
MLLGQUeEoBBUWtt7TEwbgl0VCF9i0kLJ3pofmHLrRJh9uydoROnitS5Q6YKP
tJFPL0CmYr1dhxdUpS/5se9HVuiRiNi4prt2WpPxk29W6GLaUvV6WHuNCJiH
15+kgmFhRAsYbvQRgNq/iVzjpGqGjNpGz33idr/HYkeMzvdcZr/Aaiy9X89Z
XamtlT5q96MhOyJIB2J/MmnXWHwI2Cq2rXHEMTFmFJddGcTT8RDyvtj3mabZ
ONPxiT1ISw6t0L7r5OIVNv7siK2wdq19iXBxWAh7/8hjMlcep10S2lqbCeF7
kb0LUxQ/mU6qGYtRffgkANVnDb+dIG7mzZeyl4zeE82ooQUjXxli2qsQyH1x
lU/gtwyMAXYS0fkDzTIjtabw5sGl5b5elvHKkZh9jYxruiBllH5A4tH/tbxz
qk2Po5wO75czkOLH4qaZ8Kfxt1UFV9NpBgFNWUJoY8v7yZ5OKZ9xzBx8rlBn
xEtohh+Cx0U9hPo0kYqCvynPmLHeD+81hxeUdhZWgk0lRWTOhVkpWGnI7HKP
Ud1fvL6xTsw/DkPDlRxTHlciL6C6M6Ix32Nmr5XPJnlrGDXCrEcE5rZTYjGs
aeJxgHEZGh6V3owP1vEmH4dHVH9ddBnliD0dNXF+kA9yYWbUDoHQF6zaP09l
EY8glb7T/CKDY8JwHeoQJAxUHMkB9VVUseSZNEupSf1ox4/+crkcgWMoovSf
Sfy/G6KLW82Mv+m7zqoMcjQe5RJOMglvoYf9kpZAwXfBUSOprk2rZsvOCw2L
DCVV0xXNkzZR6f8LQTiyN8t06ZdN4CBHLFyn5Nwpz1zvrN3/zgIu6i7a2J4W
81q1V1T2KaVd0SKvvH6Ptw0UFCecAHqRjO0RZlz0dRu3MocSi94xT5GpASd5
dpSkPRTpai8ICzX1LtBeg4SruA1Rpv3Dyivlo8nIjBWp0QN9V0ptLNPcstf4
7+764+HIzc60wBiy4Pc10MBxQkXhHO0PTvPp00F0xWyTAlC/Gkih0PxVEPZ6
DeZWtMxexzPewg9k3WPO17UISyzYLNC3ysqTbQgXnrruOkhgUglwXT54V6S1
B3claxKv0Ui2v5LRobPDlfAKHuzZVXJHEtFIuS3Qa3PPKy8jGtv/xDfB1CID
igMCFI0e8Nr4RgP4O4Y0Pfsupxi1sDcBEGPF/jT6T0WwEyywHjvBCBTYKomE
Y63j2zMZ4y0IF0pkbGggkQE/gL1DTIaUSLS12TUFtpWHjrZ+RH2ukwGgyrcH
rntgj6z0e6ONRD/RTGTm8yJrOtrbOnyNU1TTbDwcXAunWYAi8Q5rfdxwm/6e
Zv43O6dwA9drJnMFKk95vWJTgxjhZzn8NVTqFsQuMcmJn81bJpxhJNZmUZLJ
YLOIAKlt8sbCSwPu3WxKJnq4FnaXi6W3LUjPGXhdDcvqei2N07Ae3cSlPEnV
i2V9dN7KTOuvkdkWOUaKhfTeWAn05zWLPdy7eSGnDcu/gkgpyaQGtbXnvaxG
uhBoH43PAr76ngr3QB1asIqn+BnPWM6oelNWUP051UfwYzzTiIX6ZXjd0ibK
vrmm5kuKrplJ5MnaaRH3zex6v6aN37wtILBtOzgNH3GESHktcDoGmFs4vK5m
THv7eh2q3qBJ0CjnjA1rpkoWgr8MSMkBBt9JmRb8riCu09MWHwCJXBdrUelP
ICSY9iAqcPDNCI0LwbnE0a7WAeD6ohCRXbGWRruOGFlyUyYK8HTtZ7NyMYrd
wgbtNYbKpS4I9IOsYfkBC7WKsynwKsIE3MnCwUQDlzABsAFsvIhoeH2KIq0d
j5prezbky4MomhZZcypQjzS+i2dqw9E+svlP98e1nZdU7CjaoRD/4jVK/vsX
cJCLz9+a3YzyC1JJ9C2S+LlVz63LFJqfF5i8zsFq0oGt1+FiZFvIdb2M3ZDn
2OTa2Sk8WciVdxfgnCmrFtNjG2So722Fsvb95XVFzInmEQsM5ghzhjFcSBjl
vMYu5tEwHYWiOwpfh8lYtUUpulpqZ3LOnhmaAOBTxQ44+cvYO4PxttmrgjwH
IzS4RUpxg0zTnr8kTtVb84H2VRQd+tJTztw2VjEEHxrcVrybODhfEyH4kI8z
l3QQLFOOx/Yrq6Vqp4SYuEZCQ3YIRhfdx36r1kdKzQFZ3azcB3z2NmvdvQTX
RXKAWaWD79+Bu50sudUEBtfTqqUkCHMhvKJ53FmeL7JEyUx1HV2T/7JeLyjM
PfGgkJdbMezYWENM1hE1BsdUqcTFUPIYulOYNp0lJPve0Dh0EqcWVF/oO63Y
wb9crGJ99W3B1sNi1SdRYNvEAObfVCQM3BwrfFCYTGvxX7kcDUFCvEsXbFKF
WWY54xpUJ24nV8/Hfpaqofav3c4QOquJjNSzs9ma3suGzY4Q3DJxPssFwq08
5IfJkCodTSa4ofxY87ABc512JuY4mPQEVEiOd+yL/qofWuBg9OY84KwhAp+P
/OknLavpyrCK93KxVBkz0ve4sNlfYn1CUttij7aQzB9K+C2m0DY8DjvVykz0
YyhOWRm/x0KgmjYapnrECblrgwKBYWBAzsOBF1ZXDeAhy7YlETFlVOnoPlBt
Agc5jBKJgc/ksDBAmNeWtzHKH3yX9Oi+eM9UJz+mA0awTdXJeLb5KBtn9ERx
znyWVUNk+apjCEhCCJS/kBEuopAurMvaFJmtu8NPHTX0aOzVlocyYQxMhB35
Ef3eaEEVvebD8Jc3b5D6KHbc34N7Gl5bhp8/kn5WL6JrT5ALw4NrGIOFG6Vs
VUyse3FukOpC6os2HriXrrmuVpIIKhPXfZy+4qLcGLh1NkKT6VDhA5OiMR0Q
gtkJPJnZ8D9GF56oZ4UxUNhRT0ge5u7imaqS1FNoAhjagLUhWBoHJUW0eGEr
sJGwPtUYelxB0ZyRfB7xtM+/0blwDW7EZxcPRmav+Yr5p94+e2Nu9aRDUdh5
ViCHEucAP8Q/vpEGL3yssWrKkGzOt/nOqgvmiD91ip9xaH9X7XuK2+0VCFHb
isSZihTm/yaK1BuxIg/8EnXAIIpbDwt0mmBWSG3KIQj56XqXwL57piAcTrq7
EPRz6xG63FWe/i4p3mwdWFu1btgdJEvu0n7/EytLkYAuLOeWixHIdrAmKOmb
EELH8kXfn11pEo5B+tXeKWilyjwt5O85gZ+9rPr1CDZdxlbmTS7P7NYT+7y9
l8rPvWvmrxgzIr1hPWnJcV/TSVZSJCt9+U7VspQyBX4KaycmEoIQOZramIaJ
kidgUxe00xan05eq5yWMGdrb697jfmu4Avkjc2bQgHTjh1Zvk86yiCHiYiYN
UU3JOg0lvGKU2d96v3ipJDbmzn8Q26/896XUB/41zwJkSMj3nqIgGgnuVzm3
1T7jV0L6gun77YNptkDKpDAfda3EpJI7PtXUvrK4JyM8M9EvSVV9A8jASWjA
l65k5mI6Ub17uIrWZndYSuv3M7OCNwh5jDqN5FYBwC4toDXYSEuCbLA+WBkM
6du0qi9KMm6IAG/3hUkGtf5JL7wWT64xsg0nWUIFu9mzssvendtxs1yTyCrL
GQIVnXA9CRsBDdmfDX4Sb0zzkcPhMhBTvUFf0rzRRpAqCQjNL5rd1fUKxxTJ
jAOGaa2yUI/L6StZKm2wUSL8ozH0nRpj+/Wx/INHdlBx17N0LT9/De6+YbNc
IVpVqydZDWvpWqwlovKK1Cck2vx/Q4O5SPdI4di0LiTP3avUoU35olC3M0Iq
AAwXmd79OHuISo2G6iCpFwDZqgc9rVTnTbGxaOM7oMeImvktsDGcR9Rv5pAs
d/WNUSYYGgY3ODX5l6V/jswkQFueICfRlclpbsb+i5qdi8pNwXSKM++vyu6u
P8+0abz+WUVLuGUR4X/sCgdEITJdP4XE+TDS+M6xHJUPynDuRu97r6InNzqA
N7dJmQUk3IZk713AxS3I66RFBI5c8ik9zAXnh2ahr4gKMcWO0t0TxdI0OAVF
I3Km1FnDMZ48k6gnsCaGFNv4VBy/EhiebwT1ydatFPbFBLfF4ZPI8IZ4YMXl
tb8qBkJz5AsPXzC8HCBHaIRoV5k7nhVZoVOiGxlvBDZS4ZwWKWw9q573rNtL
pjHX3DXML+w1Zw09Y0ltWFWQtwTxZXOIbGkhu3bbT3+FsYHrtkpjhrtg78sh
C/wpNUQ1tHrFCneIOLC/STEnLALc6MO9hqj6pV/RxqwlEUo0cQOSuWevuJZq
2k9EIX1KiCwQrv31sRVhYzVRezoc7F61oIolSEaN0GjuYkvBnkrcr6/ASKAh
1Us3MT02o6lEqyKcGRo9rhESEKzcDWSQzlYdGXFAZumDCEF6bkei6S2xSw6L
QggmtXd/dy3BBgK1GcG3YNSzylhC4fz0pjcI2zy0Pyp+HAKdaBf4B6Wxv+xi
TKlRED3RVRhHbxLQddbiESr2ly6vDi6y4l4Xw0c/QC/JkU+bq9uw5Ydq2PVd
Z+3o4RZB7DDoBwmj0WPkEPFkKWxBCeU0vtY9n6EAtfNtOFrE7an5dGpWHayk
5KDKBruMo03UTU8Doh0CHNuNvDk4HqPYuLqW/z0B5UqSRE+exVfd0Qs5iZKT
Og2ufkXVS0eve4rP9gSwKtvD4V0Sk0qkMj0qiMFWo1ZRqmOyMjzIAHRpNrxM
+0a2fpE3Y7txduaGnKQyyJ7r+rGL7mTYzuNYNgcH5tIrJFWTX7mf+fxpCqZP
Es4k/sHNGFUpa7WN6ZF25H8iCTj59IkATsjjgxkjgTVLB6NNrdesgow4MBw9
uDGf0F5cQ6DM+GWqVw0K07ocYtcJMqF1TfFVJ1EeHV5RRYpJB9M0PgWjC5i3
8THMjV6hpceGLTKa27uri8mBhP6mgwWRX8HMIpxxg2vJmqgHsvhCeD3TZ0Ea
f0yZ2udAN0042K2cYhDQREN8lZBldHtjfKiFi6OGL7XTuECFDV5TLgziaHkY
lzeNwXPKkue4TcCogzePkKfsBRFDI1zZYMRBCaU6fKsN9Jfd61FbeoUPonaQ
1f2qgb+QufUW0bHTp7KFRDfom8aS1ow378Q/VMTaIZHOXYgd/NVpkT7Rph2F
bA0hwKhw+cxOZ9xZqQNKKBEwNLnJp4QpKWn96YH02jskT8hbu1fE1eEJNCBd
uTQFf35DYouxULs94esRcrt0WqIrxIgJSQZZCChjtM1Mwi1tk17DLcmE9abK
wgBiaJ7pCyhfNosDvIRD6xUeNp2HeuwnYITdC3x7PNsSJo1SoWUw8KmC+WZX
lZJ8jTr0qumbmgh3ujcE99RXSB2JekEbMwik7NWc5QkU7R6mMJfStKcWfJZP
BnEaYlyK1XZVF6I6vgkFPYeMj7K0mlfqu7naHJi0rlfBRdUwlAOKoVSSPfjA
ynYKIul6V0SRhegNpfZDMQxGWaLlOqCKeTn/K4LVwtAdkJe6Hoq4fWCHfDnw
bMmf0j40SZ7R2UljWlaj2LENG7pcNt+RZ+U+0WImaEsR0nNa4JGRq68WBbzx
PAiNYhmdkpN8iojFzc9IfPRFKz2rTNOcGjlCW9ztWgUdoHXTGVAl468Mnzs3
jR3E36c9++ZZ9tn6QiNpTD4MlUmDLrXPLGEABrWhP3ZHS44r1nSGHmiqZXSj
65wHN2bZKmQfAh4jYhoVHm1IqBYeg9r0aA1emGdj9mgwJH2oPbTmiBOByvly
IEnAek2OedkfwketFh7wZ3ExI7WVC3C/BOkjs2kKAPqxMfwCITHH66hDIIKZ
+45gOds/57PhkvrXMMYUC3zRhyazbT22NN3VIWbqaZLcKTzuZcP5OsCJQuBx
F+h3V8C+u1/GeGTBlfxqYaw/TOfAc8DOcAM1oJo1skfX8TB2euarJLyAIfys
1SqyiBNI2T2HCPtZZHqpfHvCpvrb14KF70mK7c4fdAcNDH4I3oGaX4oUPSa3
CAILNeLv+cDVw62ZvPSG6kf9jo1sBnCI7Q91nvVryopgSerwmsVhxyddkxUW
qrI5QKTJpIhGI2NXK/VMge5mvBqQDurSEQVAt63NHfyQVJLUdE/ng9vpJOd1
mY2SE/F0AslQ1NQuuTJ9UMtCBIrCMbTMJuSKVxSeeL1pex8Xv+E5BNGsKc3B
koS6zq/pENwgrtNNbcNSkFA2JAM/CzZ1Y+hho9Ioc6hfpj0Lxu1eE1/bPCBn
X4kVB7OVR/YDNHdSwwZCffsAaSihdDcpKtbEtgmdbgwxHEbpOMyZMEJYCxZK
6zC8rlTXYG0oq6GPbtKWW2y1AwnjHEjWniiaNs/34DOIFSqfHwgGQFCnIznR
K+bHhe/kpQ9xk4Kk/PeNxSG4A/8IEotZYGc/Cy4H2QYisaZAQw/aV4noXiQd
SX3Y7lQGTh9+Kw+7gn87+MT8NLoawSUyfqTNGXt1Sbmh7sA+2s4G9mYXiyoI
OPYNyOvB7ceicz5C8VnB0hcNzln1HHAxu/bKoXSrk0j1jnwUgWk0p8dZayF7
7X4BpKehaHB2PaGLZJUkFM3vW3tjqrzm5sL98EFaERuih1x8y0ECR6fepmZ4
jGb+4svxaT1INa7JRZ7DvVBtRM8s8JE+gQ2R7dndWTIEWOwpupU4eTjFIzlj
HKA+XKr/MHdkHsy/WtVchIn1mJSgMlMn6e240bQ7V/nfEDJ41OqqsZv9xm2R
hvpVGZJvgVaO0wOP//BLgMnQ5HqRCwHQUN2yq8BnDAC/600GkmH5Ttvo8S1S
VsejWudqhvDcN28Ii0B0Ghi15/gZ7y/Xcds6qDZOD6wHrble6MOWpB5FT8Gv
3h9GFrYv9oO2WEM8OqF05wEI+89D8W028dj80bFOCrP2QEpvqRgfHEm0ckbV
h5Zth2ML0fUNN5I5n3tfjVsukCkvGYJ+jMO90Tru3/MKWT3VhlqKIsJbaH+B
sxo0g1uormg6CaRTn4wlAiF+P2j6K5NG4rUEoSsP7c2d4bx5Cu09FIf1AoG3
xTF5IR3RpVfUA6CpG6lSGnauhOljNdXas8oBGh8hdfUTrfTzA7W2YJ3lBZwk
jJhRz1B7M8TTfYbPM241ulPxbhSZOnV7X15OnD/tCV8KB1uIZbfzPAwGuRhb
FwB3g0ak7zKpfFbil+G2THrGpdqo2tEYeQooILnpHdtB+ApX5RBZalHp8ccb
ffTpn0WxcvEOdJIpMoQ9sMpeUD+83NpAazswBCA/EVsY0/KNrEOboG3MflnU
alabBFwAidNwrx4Y/4vZ01T+om87o3FNekd81EBkc79rIqWmQjyhyf/0VgPA
560IaBB3epxCeYiNddgceu7G7yyXbsxpHMZ0P/cQt0fsNpl8XShV7dgafTZA
O/JO9w19P0Y56EipzljuAENwhw2BKrHMcV+dXhGautbZut18bpQ+d67iEmX+
cQhZQtuMi87QJxtSJ4GSKE2J1rFPtl5D1o+WctyM5Tu8PQ3oyEonIsRMcBB7
+YpV+9HtrA0pFHSYnUZ7oIy2Jm83yGnwqc5pLSMxA7sg7j7E/9emReauZtPA
pmw77mK2qO+0w6cnFasHZ0wBbgRRt7Jv3PAZKG7SdObpTDtVVgr+k1u9pE8S
nqcsra63vEPvNFv5/KP0PzwAmPNKN0e1A2Qvyuv/5UvLb+JZn7EePPl5YiKR
zyCqRZwMC/AkeYq4aOD6Y7KXbMOgFYmM0kL+GLqzlcrbiuTEE7P6UJeSbFrU
Dl1IFdDSDqPCSXRCboVp2MPBD7Mf8xNQNvepliJyLlq4Ejh4T0kyy+LOMIyw
glyrPrlIFPpTcB3TQomULTmDu40ilPAZJZLXhSUSgo/88jD1y79ZSg1mENDV
cWmJY1JR7NXYM8n9vjYPDjqBruu5RT3/eEq4Mfvvf40J/wpz4+gOm5e0OlGu
omkbjGUGRkGQHD77TBEszrlTeOm8S6Ic1i2R8WZhg5XuMQs4XLz3Z3dgJwWH
GT9D/0j0ieq82Q64Az+2nZ7lOxrOSptULgK1yuZAPBOLLh8KYMAY4fpOvWrK
lw223tW3NdzeRy4bGx9SidgW8skG6YFYOrRtd+Rpryd7sIKFFMuCAfgTmqH4
7/0JBtSgbRrMigZc2NzrS0vRWrE9n1fYJly7uhsuHEhczF3nGTdtEGCcKJly
h7IbkuLsdGD8ecCU2CzuqcZFLGOMITh8pZ9P8ba0LUV16QIA9fPmN6WbJQmU
x2MC8B9n32Gnogw4ftqyhlhqWkdoXhMt74QBuSlzetWoUQYVp0VZUkC0UAIZ
imrSyPFup5lHDs3w9StiSACJLOoHMRU2+CKkCjhHMnuN2MsZzKkfpA+0Xbe9
OzE4TRA9S4Y7bGHx6DJG4zn69JQgYIIPzpuwwrj8ly6TVe7fDR5zYkFdkdR+
y+3qDc0Ejbd0mg4ufZZRsiE7qNtVUPK2CxbLKbOk+8p5YLxaZzG+/uftr6M+
daBxR7J9OuS2A1c7HnZhbl692+0KM2JV4pjS+lNyF2x1OIW0tArI3fxduYZq
4LcamcBN19sVpdtJjjBgRkpePTtZsGpf1FhArdNP1Ah8vkmwK5xzWanjajFk
/Ii9GzuGjxFlUn/TIUR+WFPxP0n/IBw+f3MUGL/7yVnMiDLqGfr/MJtb+kie
l8Gs6JlDhlU1k/gOcoD5L2zDyN0YE1vkZM62wWvqKLtAINM/3bsGkZWz1i8s
W4MrdyIaXFjKN78WgUSutVsOYDnxAHTI2y5S8Oeqk07ER/RxZjr4IC/n4IHP
f3z/AIViCoJMzRDvJvDGKRQ+WEWlUM0MPjVmqlaHTTLY5IgkHUUElsVHlzZA
77LjB3Z/5H01K820b1rgUN7McLRHrebb0+w0djT3SrORk1w/mmcxjuLw67lZ
O12G7MeMaYtlC9t2Al3cb25AhkEKxgpKvYA+JqTRvM+imOtRvlDLQaBCdJcW
h0B+/g95Qb0egTCiRv+ytwixCN4K9dZTirEETVZvCaGr2C4TcZjZDg4iE5pD
f1tIhcQ5GYy76IfuWj5IjSPwzutE8PBJiOt2h65peFPY9i8GUyQ3gHw80aGh
kjbP/sBz+LbsBjjNZTzdqdb13S9DyMe7ZTO+E7UV4ea1NoP1PEoMiMVQR+Tp
YZGaUTc3hxJJR61KGO6UxFa2+GfIs+XpSTebf+sxxBXlAqjMJ4UYy/bTWj/d
QssPQu3/x4SF6GEZTNGhD0XSOQwo5KoVFxvHFmQgvXSqupy3xybtOMJTnnwN
l2l4LLcTwBdUI920M3Dw7APL9K/gHVzrm5zTP4TMKGEfIN2gq/TsrW6LJ05B
ALVKg52IvDFMLYy1gYUca/Zp0eKQZyYl9cgiMhVOHtICzp7tTrKl5SxP8eyz
sC1m76aWJyMNHRlXV01Xrox/VYSfNW/H4Zvgq3tKXjMbGitoox/QVeI6CPZy
slPHRPyW/oYQElUjD8etG09eOF/CcGaw+gLN6cKD9QMiKZ4C0NRejt88164V
7sok1swvYFRS26zJUhU31261+dib7JrHX6JVLqkregxrFODMcp7UOe01AOLv
vaXpCFmxJEE/jk3TCAVOTsdAsR5UAiJ2FxmVKgFt17oDcRNhDXBMRnXX70n1
3CT7fzkvgV45TWmdt6/XVwU5GVCJ7HymtpUVw1HUIp1eWPeRvKKdGsgkWegJ
g7WoTp4H9Nwx7Pz/2U23QTad6lq3aWPhvQL/0RGv20uYxSaz+G6cdbLP8QSE
8hdFoMH1qO6wXCJiK4H6f+bm1kY2fGOZEqXHY5xUw4hnN7Gh/Hr592T0i7rc
enHC7jRQ4Y8CWYqdLfdPS2knkAzm9fTnHPQAz8PH9B6a9klluh3dvBMKeOwT
05cP7ELiAL0IHqc1iLUeB0eoCQvv51IqMOSEwvpNJurux72HwO+DnTY8QFFd
+N+M36CHz2LoUJZdBLbc0DU/qEoAFpq9578H5nB6q0YcJAvklJQBiVgVbY45
lp59MUmh0fp40xAce36k3siZ9ODtTyaZ6tx8ZhJsycqWZk01h2tqQ/15GUIQ
YI6c+XofGnbEr9MHQjgeFlKXSxhk2wFrWGOVWd0d8OCg+pJ+z2nTEDx/0cEy
VASfIvCzQ4Iu/lc8A+m7Nyi8N2U9LRvCN+PfJnj5QnbCS5BBq+DBVTJjrSuR
bNFYhRTVKzlAqFrkPNHNoSIzAYMUZ/J6sEpuq4KvO/UwlmTutd2DjHnxDkpf
aqMceXfKKoONVxcgULM7sMUDk6evBd+bEiItC8e+Hexv3sASFJdpoBWYHr2v
Njtx8C40+goKej91dbAVuyY3/xP9edrLCEH8JXxO7gh083Pr+lIRxnzv/Phl
lVMQOCNy6KI3TEQUhiiaocq1iH/YW/d8M7rVRqYcbXsOZVAo3zlcrStSew7S
c4UI3gSUoo1dUzGciRWFeerV30BBjg0GIy3Y/9r4AwPreBdyNHZX+dS8BRkG
7EuGsgzKgUKMejQ/foCyQ+ulQAG+g2N5aCvosxIgnvN8qoROjWxz/7iUtD7W
EFUfeF1JAupXRUWPnsvSx/k/8+Xq0WljSXjS5dEVm9ZhOjnc14oUWhjh+dX2
Vb2yF6LFHzib74T9jVFSZKCpb2he1ie78jUAXOblQxLijp/6deeGnOWLyYSh
sZCJnf3k6xm1ARWuM3rf2TUzljKUzWvFzuKiGc9qUCN+ZcjaQr+L1GEOBdiA
CSV5dSl0qHONz7gCp1qdxPsYa8WwEtFVVeJvyi80jifvO6ruxb4xRbZuB2sF
75hCoxxOyFfX1NfGpS0ss19AeF6dKZxJulU1FIdjmhkQnMMfe7fdRKwtHX4J
t31tSSgBWeKLLQBIvLFrTPVXZHhgWLfMUlt0WrQxnwPpDGex/EbI72lbljrl
8DwnjItsmP0Qi51DswHpvbkm3upsiInKfrd56SQ0Jqby+AUZk5o5HXBiZbhZ
X7dZR8d9+OziBb38e2v4Q2RH875Kd2BgARSEnMKUZdp3VA0H0dLFo4xr3Wbh
o7mTe9SWHsvIOs5mjiolFG0/MhM9iQXaotUcVCNxQUIKC9wbL443rWWsLD/G
FkR3y51lgKGXuHBdGnxlTKlZborVzr0U8s611D6A0nrsWlTwgFVaFstDRdS+
Cvj78jf9jM/N8uNrl9okQQ45NYUPL1Q7dviRZov9sr3i6sf5EQ7x+tpEVqMK
IWYrrGiPZZfNDUwgekZrIFCKUAaYNhj1G+UHo4iyfHdt03Yfa2D4k4yJbzVq
3eGLKZoEX6u1pOVgfuiGb1SNklq8tLqu0Wg9YhksS7HoQf5s2KwaIA9MMvk4
4a4TeuOwYbA6TVTjUD8AFeV/bMRQGYilJIcQoyfzPUIDBn4Mr9XI+arsthaW
dLNT8KL+hVcPhz8fMcyn9ZjGDwBqHfq7aDnyQD3f+20IYZPH8/LPDB8HF52S
nhyubPAQDKpwpmXCcJTzWHiK+7QaNiMT8Lsl/HhBX6ZdBMRUMdVuH6/qnrfi
1ZFX/z2tquplHexVH8/dWtBOfk7UweuvNjuGeAcBDRPPtqbds3ANTK+fD+wL
sXFFdbF+sGrt7gr21XiPYSXFX5B5Cdb3ZTw5Bkl6jACiLKrK3AnkhstXuaK0
CbiyfAXMvaDC3tViQe0Xs/qBeDBq9kWvh1GpSgbjQ7eVM3USWlFCrXk0Yg6n
1ah295Tq9kVkFrGyZ98gLJSIHYTySM2W20RUffj/o8jqzcbCM6q743XGRPC8
UjQrYjlWrpLDJ/aW9Go14IhhieV3RpDpm1VRoA9qlGdG0sdgcMqD7DL3FfWz
QENNzoWx91DzlRZjPl+Vf3NWVPkZ3rjVgGvXeFzvLw5AF95fR/P+KHuiaYi5
ZfCsWSrBKMPUb7w8uDLY5K/C4bph29h0NI0HMppRS+uXPtq6R/7f5JIyOgZn
ajxpb5PUxfSgpiMoke9dIZvn/yIUnp/7/BkpvGbxZUmQ61HHz39+834RrNbq
t02bathq+d8Gn9velr7bO+yV6M0HSPJl2yxLHN9WgwIrPu8F7ucigJVfGrBF
kTVJrin8EydQu9nGS5R13ag51gQcswj6/yS5TEI6MCZVe8KRMPaZDQdSUWCY
Nns3kPHV04o2VH5iW1VSfMM1fv2xXMHZumbGZ9QduGWUgOAq2voRTOgHaXNY
F/ko+xyFvplipuREh6FvcKuJg8fMi7jw9GJnUwUBwoJuHgPLBSJHtAFAeH09
T34ATeBAciIvwWJ7xPiUWN63oo1/p9GFtgZh0j5NYjt900hQGOg95Kzpesi+
ymWbIs1FDXjypXQYJPEQ5hdTl1xGqoIR/Oh2jTPnrxWuw7kryzii46SNo9WU
Kl7898/rN8I2N1obg1exn6+XHV5hOoO4RleaeTppk6NpQEScaopPbtg+aPF8
o35IEHvxyxGyUkG1CK9LvckUkQBQCxwRLg9YePC8Qcz8e2Z7aUcumsHnze1o
SdcG+J3Z8ngP5AlOP7F/ETg7LDe0NOvLt4fn9yafduIBjy3oeBjTD5KcOoKd
tT9yO6f4vla4FpPbF4FQ3AIltPJfuqixkhk6Dz29FNBcXf7qAFAonUMGNQ9o
UrsKbAlP0D/yaAJ547bh+tFWccCMDT/8z3wpWf8Ar6swynoDByQtHxV0uJWm
UwajA+w6w1KyTRAV8oiVMk5dE3fMu1AxYLYLYLwQK8qRcD16Ls7i4zDSU87I
toW3Kc+JmRqaCMWk9PQPOoGC1Ycgwy8miiyK5lj17PGbAqETnPaT2z71xsjz
0CarsieJj5YRIHpL4DDxx7PxU08IJVG+Js/VWw8/TI9gU6nJ5pjo9cGbETZS
wR6zQwku8ui/lA6PZ4tFCRbw6cMK7kB9qSEKuc0TMmUS7gbG0n2XwD0LO1jD
xcOofezGXl8pqtO0CiGJ2HRwioekt2q+u4wABF+W+nEKatKRzQuStTv1iE30
KnVtRkYh5A5kGi3HJ3vjmLZYN4FXzmzMPqmeVbdyjx/NvKF2etXQ+n6VAAls
ZKmB7Et1xnCDK1yy+bjnMmkvD3dLYTTo/g5b0acAAmeKCyuijvqgjN/MHjDz
Rhlgi3gIGtxCqNjFkGvnxqIKsFsowU4ElBIs2ub0BECdWh8ZAzhvIwUC5chg
XGBbBSyZomibNLZViolNZipiFYeBOKGuWRwnsd6Ls6o6rpsCgfIsKf43q5GB
CrVv4c7J5alVE802SbRrAUDfjanttJskFlFU/JpyThI4dJnI2lmClfU+dOza
y35fE9EFqIOKsQWcc88xceZuN8itv/Ez4hqtShPl/PU/JcByZHGWlCXxCiYP
vxfra7ELT4jHMvssrFeg75eMWzaIw1Z/cruHHdBx5igzo5G8sHU0hCm21rA2
4XhMInUdlVBglSOpfPGS02aeH+T4okQ+AlXoUUTT/z1FzKu4tZWjxgyopw5+
CvNJftoeLzLbkhKDe6mPZrl4O/ZNE0KCo8omB+Zlhs+cfImw0KlBtc8UefKI
HVdyGvAR6iK0+e0cziz1wR2SVwiHXMP/svD/zj1upGCoNyWdDwm3OVc2egEP
s8mhHGwayFuQZF3ztvh5UwU+nDLzMWgBPEppf27W1MgtWxWgZ2FwwI6HzsPu
WcutOa/x3rqYrsg0e97CwHkeV8RNm9AvNQiuNSrxIQ4mXjXX5aYGAqHXijTr
pmyLnE3brzUW6Yb77uLcqoCTgWyhlvPQvBrpbN41ewAFa6TfnRASEZXQBMFx
cCFGVPjVx5xB7Ut0lxiCZpgtyCl930CHRyx4ZH3xTTMCC/RnK+7/C0WCQFV4
tHPamrcYLy/bvJ5MunuFWYiLRhzJPwtMzPD7nNQKH+6XCheK4m9GDcSg3xPf
9iGd2F7DoHwBm1bQHdvRguHVnH9cym0eOkhIz8M2k6EO5tClVF6KdLWHW0m0
FfxJxiY1Gi1h9gpaXm6x/zUqQecNtiwA9P7QUcOxzjbdqvYt9GGqzfOmZAV4
KlXB7a26Fv0lj1iOPEbc25urWDrbPOFwLJz4JmKlnksgR9M0+WYCwiTd63Cx
zvtcOl5+O+nSWJRZWiVrcHgZA4qg2cHNLfgc9FldmoR//f4yk63oVZPo7ugJ
beNgrOTDhJlA4vzSEj8/qGFkSc41ruoGqXl2IVzC4Ys0qZj4hkUXPEatqbFx
5eW7OHSpjTSYmCF6VyRbpzr61RE7jGwJ/9y8tlk/ZY4udLe8ei2JNGO0CELk
9MhRT+kYWmVnzf/0WfSASC0Ivoam2crT941pE7WOMc1l9/M4OubDOeBrZO/X
JIFz14O0PnQSx0k18JVua67rMmCUs8I7yizZXYYBljj2uix4kDHdZ2O7ncKE
9BelVOalTAgoc2LsBvNBCgfsNtqCEfC9T3dxFugnQ53HWN15dvnvX2Vjdbkt
1QxsykZFUKZJli/BW5I78voIw8VnG1/f7ElzjkYP4T5ByjcGXhLgxJHzZbMX
kT+ng0C+u9F9HZbTevG3aBJJt0xm1ocj/F1xgbLH4UeKkbbX9Crsl8pDFrBs
UCtQ6XNHFHCUSVPYChxVRPHWlKj2InI47yu6ELI+9bDC6BEgOCZdUh83LTel
EyjsRiTjy1gWTTJh+KdwYd7miUqkpW6v+uyE4O/WfL9PNTmXWVWj09b4S+o2
CS/F+Xx5PL6QtaP9MpUlCqXMRUZL5UNxSC0/B/6KQ5UpHnA+OA96by+9dYO3
Ieipxje7vxbkrvvyQB90L8+FTlegAM04mwgyAHRG+LBxNllE8peR3VDt0QNw
+a6/WBSWCXREwhI/kIkNLwzVjTGYLEHdF0HWHvdKgjK35KE/3G8utuDnzy0q
UkkGwJcTiN3rnin2uRi0bBMUt2HqcfnGdBvkxSz9j3zbhzFLZ4/0LGHNXMYI
cm8oPRPP2rvRG7fog7wEEDhh5Bu+u78sefBxhC0FTMB1sd51kD0HxPNWQccb
jGfIl490yYkbueZtBv3vZD5KNhXGGIbbeSdjCEAKhKdQeow8CN+23e40RXG6
NJ8jGFKQu6/votGmA+EIweuHtkuM2xu66+pH9Fv2Owc/tIXouoHhxdxQfkbU
FQJe1M74jFBDmE3TQGzeykIgwzvkuh63E/MfmLXUrToNvcTTLJACIiFsGpfr
olN5trqjz5LtUzv05Zqya13RVpsCA0G4A+GuEAj8f1LdCc0B2gJRLFdeLzeQ
ETLZO4Two5M4Js6BOiyB+pyJKOviaHKUuzte3C3ToPCvj9NBOqDM0levJUw0
Dr8DNDvaxzjRjurFBSqDrlIYLf+9v2oq3ewNazi2ff3n6DZM6DGZi/b2l9UB
l1Gmk7bxip1wrsLFazQtS2ER88qWnKuqtKw7u2lgHLDycJbsFalsYBIehOeQ
Z3Q/CDtg7Ll8gXYsUz6uP1trP5No9prm3cVrvWk3UHktd6EuJTZSmrJVxcrZ
ZDdVqmh8/bAMsReGumA+D51A8gWW+TeqvOTvRy4oLVBG3fScf7U6pjIwfCBi
BbFAe00PfEqVCSk5KEaNDTzPNDJkj898kHtS67t8LWHqVD7jrTc58ufnGb0L
SfvlxhYpyY4aJtbqOEGREAYkY7gj6pqkX+RQiBVVYzBPXR3MrfgSzP9Fr4C0
hiq9rgPIj9ou9KlSFvKaO+oFZ6O5e9Yqy8jN7Lro8rN+3Q8zt1v6BXCZxSST
TU6HOKwSLe2vYo4EQ2tRoOQDoKHm50VA6h+T8I7zjazcM4YJm05NOj8U5YHy
Pm9a2aukNJpquDhr93YzKBNbxNOvJrhBFIuy1EprP9gJvIuslOJJeSZi87YW
phe57wgBtlJuMdE1vnzhktTPNKpJYza1ugyojE9lnF47dGoRvYLrYsaRDnK9
OsZ0rQ45RxkID/cFF00nDle1i2Duc/dq6rSOo2asNYoxBB6e4S4oArqzeWI9
Qn56BKZUS0Eb+EwuP4K9y6+PyT8ESzI2GxgUzGqxaoY3+EPBua4rIHHfDrl7
tmgClBepTXVCERWI52NXGFKf9XEgD9T/MsCO56+dLlbgEoSTXWiyna6XqWb7
Emq60vPVry+jYN6Mdmhawf5VYRtXXA1MEamD1ySY7yh8VAuO3u21UDRkbD6L
9c2w6t7VzFQZsck1l/+ON15yVnfbnJwZ5AWlcYg/0lN8KNqP63Yi6eHVRIJT
YsL/VucdlW1wou1daNuJfR3KOX3wDCdwx8JdRCb4rxjOjpHYpXUHhtu5apgG
jZAXwDF0l0Sb0J2K8k8m4JR/RTYd3sMbqkJysuakAkSOTyaP6ioZ5+w87cD7
2XLP3aEkWbI+ufZk02hod/Ry6YlG5TbESbbqH2fEKC2/Bb47jYHcGKWJpATl
1GBUswkF8S82Nnj6rUDfGW+FQAnO9Lq9PmdE6cBOxMuqtBaY5pLaUtBMuuH2
KWopojzEVUeE0GACwyUn+RNvHoB3fhTzwgULRIp5XprgOgrNbiDPv0SwkPSZ
FsjLnpVPaWiq/jsFQVMn26gkjLCWbnW+0jdKzF261X3IlfPKBQESbwbXulI4
vbq0TjVnkHF4A/RdNQQc9alIWbQTQ/ByhmZxTmVR4U48s6JcuwY5r7xNF+KU
mVb0RgpKtpvCXnAjIhOYnKNkWdlpUIvXVkQkt3SJ07hhXK182fEUoe/bUHwh
499KVHb4H7eOgcfk2EdzOQmGyjzcq1glSgUZt4d/buFLkvsQsBC7+aRPvImE
uMhTR31oR5oZuBqSv9iKwZAZol0/kp3sJWhH901v6Ny1Wp9UVA4/xP3XovEt
NWIwUg5Ue0x5LuM+Di18TIjfYoU/avk9a8C/EwOT062Mod2HiPpG2ObN5FHY
nD/IX7iuN0WHQxR9pB6xk1qKePtW+ZZJaBXxWkkjlpzaH46XGxI9I3o63qtr
XXeKFB0uu79VkJ6f09mVwdM/buOqFOWBUsEdYIE7CfHrm4YtSuSXluMSRMnf
zqBm6pR9aB6jtrPTU5lDJp2k+ygLeHaaiiQAvGacg0KsphsduMYbQrGpnBpk
7zC4TN6+puCtmHqxbjo9ov9ygNVkwzdnJRM5m6OJQvb6fdj5tlWB6P1RkWDR
w4GeYXxXY1KnTxIyGmYlah4AlD+7CtyiTcnL2UUmH3sKojBqDu1smT/5nxd/
e7HTBUkiNuA7BsHAEk3nHIpZzjlRHSlF1XdwxUQRSZRwaoMj7V0PdE93/i7H
EdxepJNb4xr29a1Bva4mGVoxBt6pD2c/dCrxw6mDIyEzLFMMVxXc0zSRHoFn
AXtn6fFJA0/PtViP8TgZlfjV2EU9Gvc67ZH83vDa/oUc+DIKubxKD0D5tdA5
vM+UUr2ShBFEFltICw3avPG0rwNx0uE/AiqH8MGww7VGAnCF3FCLlMRUe+s4
DiwyYYihBFKnB7dZp002gXzPIcY8QonojKH+kyAf97dlmYaHLvPU5DyRkhvF
btPlKqErCS9L/u6g2Z5dGpsuZO/poJoBHqx3gX2iSFaRlj3IWbf3EucQxtfW
uoVCcPRK+13o5kjrHUp86+tehIiQrLQhsy7u3m/M4EksUGgn4rWPJnDL/T+d
mZ5qh//r+dE3UjTFR8dXmOYFvdh4LzkXLXMzulKQsqRJ0DUTW6R1w6FMck/P
hH7C3LKpwIZFx8DoYS22jcclaD/X8DO83nuaqhPJN0x4BWNGwqFEvca4DN14
/UVGwe5Whg129SRwDFwMvrOyPZezQP3E+onVLQ/Ure/hZ14UjKumJtoZb2vk
qIBedB2pYsylQpkPrNWEdDlBTWq98XAdqUgqUCMXhFgyNf9kZU+/yU7y4o4f
UlxwKDx10egTxV/8ttfWAiQjHENG+155DMoPghEF49QGwelU++836Qh/6t8L
LVj9FWtbbwcTiSduzY8+Joyr1RY7AuHzKwTYzc+W31hCJ1dd/YH2+DOWzdLv
gZRCK0YMElVw3s6Im1d93b53MXLUXxNdmOZECYm0UwD/0q9+A183Lu9nmu0f
+cczfA8hxYD6CqYqbrqdpag4Dq31Kqzzg+7PcT3gzxVGfnPHkcqDPErkREwf
/0+d4FxvYmEbFyvQ1BxcVzTvm3DzEnUfUaFmILmaudQOqsaZMMrtge557Ovf
nUvNWpKnGvWVaqfz4yNZJJkTXInBiyEbjIs/WKN6NzhO+tQHMO41l4j7I5wT
o1p6RnDdjY3QYGJ/jiIIZbApGuafW8BF2uBfMQoVhU8TI+Bo77+BzXrod81V
EBrat9euWpU1OcO3pygc1WYbN5QlbUyW1Y/MPAjShjyQB3GqaNvTYwkd9ygK
YdVsI9BBhISUky2dauWzn+W5s9sDuDPK00/Pful9Pg6v+5KxabIQCqFxaVX8
8uU19kWXNVDCNc+9KCUqCWWYcOC6dVNF4HNa7Gb8oFn09f3MI95fZRKodsTW
VNXriys+GyykJUkVv09VtsMIfIpwIMqvspZH5N+OOUeJjKF5xTyIB8txH3aL
PxLdxBeK0TmTjLhagaaMHhRz//flOo14ovq5sk30cV5ZJBEFQRtETuvY4cqH
ldBslB6SCd5HyO+JXvr8Xu6Lu+RMlBvyMpbVAmrFE9ffgWzjqexuDfolm1sX
vomO/fhhun9A5QqGyNKTExHmeSU304hRM6t7ksuzybsJ/E5xOKx0qIbZaCnS
gcOUq7LXdTY61FXidcbpR6rb8pnXpbz8t9nd/2VacdCmDBAh4JJTxoxhEdNi
EbQIQPdF3eoffHPsIYm5iH6FDIbV8UoBdDHiHuNId8E4+WYdjcdof3pE8/u/
MXc/rw0e6bceXOjwsYkN+Zt1Mf8YDoNPfFq87ggiRtD0rKE7sTWY+CGNf8+W
5rftqc/s/UcwT2CrXa9tDCfIRETDlNb1Es+TCK+5oMbelow3F5lxugRUIdSw
ocxGGxkmlVaS386cL8JabdQipkEL/RvWOpDfqzEaSiZkBIyXj3oYuhzp/AiU
InpNhfpLDp5g+m+Ne7kt+3gf4h7yaUbOkvUXBci/XclipMhRh/u+eCnsw7hO
Pb2ndqwSZXRMhP9z4pfUmjxJIth6e171PJQFyi8NJJw33mqiymEt9EplDy7H
t0y8YFQNLa4wOks+fFbSNpfGTLxLJoqDgzYsYSRPfkjGZ3VfzWWIkTput0BA
fe4QfnQwRGWoLYRtBHcY70t4VO4K1ODsA+89isiHcuflG1nHFdyhz+Lw6Tw8
zTixFp2rPe7DX+UiHHS+wGlzU00PGW3TMWWZBRdnhYN+ufbVKc2HoMobVR11
4n3JxwrgLN2q/g8KktRAkoA5fl9vaiCDqEjrppL5c5KZpKTnaqcG3A7NFMk1
HsmZYL2XS68cJv/FVhK6Jag5V9RmdJEoGDXyrdOhv2ajiUXMDoSPAfgBvukd
c1nK3XNH4SOw9bCDADb9Dj2gqWPLAwiKtMzmEKHn1yVvLuIuxLSuILuJpxWF
GBwSI3xcgjTXKd55MRPZ6gh1w7kQ52lVJvGXN6co81jXrBK8CxUhoDFodIzv
WWCd2pwn5o2wcQ7bCVWyMKXzsrfiK6U7dxscWIX4y2nR2FNKqynqf6l2uNKH
aQ1JJTi1CNLXQeYHtN0fv51REZ0J3IM5cfXD7Yaof2e6080dL1SktaUdvs6S
Vpm7JSug2kYJgDbWFyButyMvk8+Dkyl+GbtBnWCsfx7630YZJ0uT+PX0xhkw
N4UWsIxg2ZlGrGukpal3pxiF6Q3iPEZ3E9wlkMdWFNDdLH9aP3Z/vkPG61Xu
n0CVA9Nz/BACUqnx+tuxkKWeCAvRHIxW4kof8aeSZrjfw9oy3gW8M+4w1XA3
yWmFhPddcXmVqBUs5KKlO1GP9WooRv3+Lq84Wh6SQT6J/sIJdJfMT9go6C2U
rYSYRaNlNLTbhfDVrYyYOlLi9p5gM78gqj5T36mug9i2Vd7ftocOl1KJj9OS
pBc+levRpLzio3pJVkKELSPsllAz+M+uB1fQ3f1cooJWBRKp69Ap0bHceQuf
yuj3JKD+QW4yCMrAjJfnKtdMOXT6NLrVwYPEF8L81PDuzhYv+o6Z2dlVuFUO
e4XiomYpqWUTRVM3WrAQJin5/TMaFZrq/LUoQUd4blk2YmIteEkTBQzyNcCH
LceHUwpKqW5r6DEwp62JD661nmOToY6R+Ho8B8DFpyTwgUgJ6jG1HGT05LYU
GevRaJMgbU/RpxbblSkCtANt7Dc1EJW1kk7Carw1QDIvDTa7x5SfgrHK0mrO
io1cQ7zqMRmXOggqMGOP9X2AiW+snY1vp0p7U/L3XWfpcyR5I3el8vgiu1zc
3bOkAwZAB5rvIqlpiQ99DRax+O8dqZYglkNc7e1SFRTah5wo3+GgGIg0pT2t
aRNK4Ql3Wxa4Mj8MNXGsjnC9dtWy8sHatcGHfWC34hgs8rqBR3IinfrszxvP
fHfdi+AZfd1AhjwiKuB1orErcEFfMNaci8KIBy53bMa8fHayWEF/pl4x2khb
GSfhHcPX+T7sLUbORWyvJREjgZPCqN+kLIRXRq7Bfzj29j197QtdsMSI/3lO
TdzMwycmiCNFpOhGcrosHBxxTyot9JhfPaZyCPEOblNo1HkFN0U178/OhgRI
RuaaYvMIWixorsgM/8xWaUIybpD5c/DS7po/MvBpkwbU/DKXgx+HK1mPwe6z
e3rfJ9nSMRoViJAOaE65/IpGhjWj8SW49ZyoEkllKC90gclc1NzMEHPTVN8D
YK/1urLJuNoLQN/HhznvZBm9G0FPIpmsGAWR8pcG2hmA6vNdJ/B4nA7Vevez
iDWqdMtuzrScKUQOFE2vsUOt9sP+CUn/FlTfYRfsNWEChQ81ABNUTH00FzOK
A+aiphKPzQD33TMB7wuSMB17KK4H+kUdCWvFnXbRS77grzWrM/toKgLyYUa+
wqDcsIawlCovVqSTsQ3sfQY2BhwkBywDGBjv+fbSP/UeSpyx8H4t8cA3QU4v
ZQcf89yQ+iUWMi7ox5gfthAXjM+9TSLUBfc9Vy7gD5HZ9VvAROed6AK3Fswk
4qykjWXhs32suZwHfo72K0CDjGLiSD9cl1CwwA9wGBmo/QAtaS4+cpjelqfB
7bZdYe+OiEwIX4jn9pkvIPv3a4RTm3LPUUq5TpcUJCzmqVgaUwS2eB+LsULX
y0IJsqQcHPhpulQgGiPhhuyJVYJ5AI0QV596DlzFY25tOZPPucRT8w0dmw9e
BMqMsQgobCQ5otgT5ia2m2dAlT+810jOVmOcIlkT4ImZIDXHx3THEjiVsr/C
gAkzPIx+zeYm7v+qB81AgZtnyWwZCXcJ7IXg91Ik1NS+s9DSSJMaZDHxI0jH
vPho/819tVs1z05GNweeAQFpCXUffQ34l3w0YN1Zn2PduZslqNM+hYatSReQ
NFAuWG4k3/skCHtcYLs6LVgIU9mYsdRfmaXZFNafYRewYDV0TB1XMGSWvAFg
/v7cC9jTNhoM5hewp1qrd5CaV5QlEF3m7NBRM+Q4o0HSpH64E34aIkJscOvf
t4ECWq6dn0czLi3BTmgVpzeqAnCTfZyaVyCHLnVz9SHwQRg7R0VMBzZIQUz9
ZP3+bgpnqc02A0gSOVPZtXsj1KUo72P4Ar169yvLDzaB0enFLM12sxUx3okd
r4XsSEMV37QG1hPwAwRfLCSw8OgMgGdbKtqx/OWqk0QmoGTWarK1hj4hCWLO
kO/XMAV8HKk9HWY1nVi0DLXWF8DeIdLPs2R3uon/A6Z8rGwe7A/61BZOAwyP
hMCkB0xIQ6iMprT27TuPSXtD058GYODrwMt9pfI8ikA3mhGVE8HK6/yVskGx
ayp8jYprz0405g5YlOkIBlxJw2ayuiwV0AZvBxzUaiiZvuQ8TQVgIkK73QKL
3NY4n654hZ/GORB7H8I0pobbhrrBbjt5C9X7eUREa60llm3SPFymD0XTJOlF
PNuDwAvvdDr/oN29c5tRPXXrjXbUHPP/1wkNYx6mwOV49wcjQYjqk9LfH1q7
1znlp/22W/wiLjIlM7A8bh9iAmvF9yJwrNnCSBdE7boTy4yqaacAG+ddf2pR
XSIqCQdc/BTJ5rI378sWeDTMkk4YkRs1M+HH4cQG8uo1Ilkdog5b/IF4hDcm
JeI7sMf1EYEa+Q1h9ulSP5rivbh/HgbtyHdtY4FyvzSU9CSpK2ZojD0P94Gc
wt1GJICRTAptEtw+Je06sMgcF230oh11jeqzoiHYamwGqLHWu/zJrc5JeYtW
8ItXI73pY0qibphcGzoGLqfTVCBmpKSkwlQN4Snc6x7P+Y5TRgUxF2QZdzqV
BTLdZ6HdOMDUN3v5MKK2Fm5awJbp5LCsAPfCzttpPVs9OPo1zATQoqJA43AL
/IIyOGQWkBMmmSh9QKS+m9EKf2Rw1PeIq8852X1C8X83DX1lhB1IXyJ7RGtj
uUlR5J2Ug/g+QmbijrXuPyaj4N4J58O3F7s+cfl7itoRDLUEAj7VnaVs/VVI
PDrnOj+pGpWPVJna6dKrtDdcEbbqQBOIJnqGnu1nagTaltL+azvNFgWAmHhs
SZCZiPhimTJrGA3e8GutQAtw4ihQEh2SO7vcftjH1v6+KloQj+1W+geaN1S9
uz9HtyVQL7AXHj/MkIUe7ly30Z6ZSs+1XbDq8Bj1rWzx9X4PeTha6aRoKNjB
SZj8K6z2cuoAx3neAhNvfzJw1NeCK9YvT2GFkbK53FTBG+CGJVFn3lO+u+6J
5V954jJDeDi6oWT83nrOAhH7v9ia77+W7zSe4F2c67hXGJTPmeuZHkCLUBKP
Er/MufOF85qOhZgmAmpzy4ahJ840oGoZG48eCT8BgLRZLyr5+KF1DtYR0CZ9
6FmFf/kQ/T34FzkU5BASjEu9W00CxBReASfmaNjNHX2G9sBBV4iCVCu7MPnm
LKGipGGLVMhkW0gSJLdW5M+JdSfV4bYQV79paGW+SeY/mJKcfDgB+vL2z5el
chCWbToCHHzxjMXrJiaGppBpYsUAexGZYtlzTqJ24JV7W9dRlzjSc8NF/QyN
5Fw72QrugmWZXrJ7N2hs4vtHR/NGdxwrZsdsv+/F+k/nGVA39ytyOvHDG27q
mgAt+xZKsrGLMgxJu+HjzEjtxNK0J6I5dV3IOjoj0y5VkC+0mWn9It60XcLK
l5grqiaFrI2albVK/RVxp2GJxy6q3a5HsQ94XeuO0aPQTuDVsgbQepBXb6bO
bl0WcQ0DSXHNLcBUhm+ybjHeZJfw6Ez+besy1zgkAfz24zZzBcisc2BoXoTT
Pkbj49Zv7/HMAk/BnZKeXV3H66dMASotpxt8r1Z0bgJhm1vFtj/1IioumL08
dy1PbyrKLDTeQe7Y0pdM3FxBnWqbfPEt+6m+zGOokQL2S1wxJbQYCh+9/K1I
Zc7XQfVdrGQCSxlbF7bN1w4RnuVH448FMdeSD5i2qcxB81chPLLWTQutNKIf
1wGr66fAu8wI2hDMO/Ehza1PMiMVJXUMcZhkTwri6AhZOK26ZsAeUaAuJByY
ZBnXd0e8xJwhU/lGI95Zl92Xsj1gnOJSznn7lfgrI+6TjlSxGv9Y6xedLA2j
4NyC97dCPrYuxABhZUQAL+FPJs00plpyKUX2ZZsiS4nSAuDb/l/h3U2myNUk
HqOltm/5LN9fg41CMohiTDqTvfEF+X4GSoaj/Up0bbGv1bJhAvSZdiFLMXe3
9bkfEMDa4QTLRyl1+kAZI4KwHvd4yF/EKwZXOSKcyoJnzQqJFHx1nrZHljZ1
+MFkog3iMrg8q4xmZwBUHwftCkZDQJH7BdhFIL0VoLkmAloxrX0E/6xb60tv
sub4Hoc4tQq27y/adXzbC66rquEjiqe168iSfv6RPs/jX2AkAXj6ukBiJ+gN
P6xbMRHCKFpkrAhORR9TQ3Dc0vhuzqhArcO37SCKNAmkRR0STdVpodC7eG6e
ULh2TRf3GmbVr9kz4BqVwxKUfOufmakzoII63mhv4XXD7TgWnJvovapReH69
YH/vKnJfnqNIRVQecQteGEB1dO+nhUGM8iMAyDPJwdI95JMt2hl61/p8Ct6a
7MPf1rdEDOlWxFf+mxh0rfhe+ELJhkPQaJahlKXnhpq7kstwEKqVY+5IlHA5
Aa+0ck5qZ5ZY7+xnikS9TMB5jcHDWp0BtalItZJdHLxWHf8EOXjEN0zQf9qi
kulGEihGil3tgm8x4on4Shav7Lxm5gFlrVqfKdPoDF3ZE3In26F/Adn5x06e
BNsAPm/bveZ4rl65RU8yM4SUQ9k0vDqZStIEGePRbJp67kDwlcaik1wtMM0a
jl5pV0tZOIy4xKIrqt5emPaIjpOBvqb3CWlGyHaYSx50GkvdVPbCCB2slBRX
AdrH6Rh3rGcy1/gVCKiOHhkoAryftMRaftsH543vd9Q38oSgYrxDkQWyg9Fn
LuI8RUojJ4OWZd4JS7yUwYc48Je6aqIG07qIA/0TPl3+Vdtg0OELuTlrEcDL
eQqV+qf7t27gyja+JUVliTeVlxDgbHrZws+IXoayIKxx55gNfJuJc5o3/uEI
a+pyTJXuGz2CKb9QO2r/NpZM6kyAENcxjbtDmuV3AHmOr5IALVQayHdyg/dQ
x7mbJi4A0zygFV4AKce8S+H4+7sb7kSBuUb3ETmXoC73tjcjltwUsH48OPK6
A2wBvU9LWbBNlMELaPcU8xVzuwYKxVHRZoThv9YzGMLffXRjRMDN4QehY2Dw
j+qecbB+3QBv99cJ2IARIvxUf9c1jjRxrPMCuHq8AVkDkJf+EM3Z+c9f5e9/
a4idvVWfY54pQDOFmFV3gNH62OLnHqVCmBQLJ0bU544BZqxUW7e2Vt57NdIQ
7o2aFOYsMm4dQZe3ZfNrX0Gf6ngLjuHyuabvgKfP04WT1fhtHKciwbMesq/I
CdV25B0HwXqO30LrzGegxMtSiGkDkMO58LemA7bfi01C1+DPoMzKjsNcTnsm
kdqrxa23z6HT0S0AlPqheLqEgo+h2IX/C63/VgE4RGBSngoap0l0ZOkcEzPy
GK8r1o/7QNwN9N8z5NM/vO6LnekThafr8Zwn5hncF4t5rrtV9X8KEe8cWLMy
aIVlcojM8YB2yQyD2i6Ij5UwfQg3Qh05z0Ab6GjZK0v4LDaoATZhJI4J5hfY
mJ/+h84ydvDpbz4TguzGAm4IReH8dqaUBCCnni+nAbosWcgjTBkYDohGqa5W
5GAHad/QplDyY9Y0cRO4u5fMWSKEMVxceHpEmn+Ha/k8hrwZ9l2ERlwVku4m
6iIujbbpirNKEYqSLHWGTfCdHq7HBFQLp6Xh1GCIpzbxBMZ95E5BqC84e61k
evR/LhgFhs2ebDl9GWN0bW7k3DcJo42dpBIvzT+4ARDYAV+Skze1j/pV8eFQ
WmcidBPXPXitnpIj+zXDfwCNoE2g9N5caD28kvZgfF5zVmGWV8QMkQ2aGvWW
gRsWRxJlb+Zg+k359ODFBBu/IAwcqpVRiuUd+RQn2FMQHL5jhtETOU2EPCHL
WaFcQyr4tKqVxKUXpOhnqgVVI5yWmHSCfuzasN3Pigp9a8cpO+lEh8IDEb48
VrmaLh07Rc0rJRy/UfAP5Gk8hRifrV46UGnIwhJYXyhd6gpq8qG4A4gdUN8G
OwHOTa7gQ6auQ5tp2sW6rVrwdK3flQZ8XmSfpWxSR4bwbhwjDYqz6LTI0+CC
rY/tiU+yrFaG5AEY0aXowLV6NaYvK2z9blRszCpUYudbt40yMeyL1pnx4dN3
y6/sfiHvRWvfG+RcqZHJAVpwMZcRZg2NEXXAXf4uAvia1rbAFbjThKRVGK+G
Xj7ZLrYIOSASn513LHndpUHSR2uFfQ3KW5OzyyQSNnuM1BYRkIFv11McgpI1
RgoEs+KUNI2LWfisCFz1V3TebrH3CIL6oo8MkV0H6aC2q1AUNNJY22iNXEUn
sglg1TpGM1JLavsdtJP0lLqHy1Gosl9XC2b2EOdKNG+zN78RT/fnwY8b7jRa
hY6z+sPdzcesfRIXvURG4PMhQdrR8Mt8KFf0+v5RDlNlXXHduFkNYOLHj1p8
JgYpfeIj6aRZtmN0odJX0n1sVkzW84XR4+Gj4AB85EbOd+xpqTYYU9rohs+Q
ev8vCdIwF0vyn9osbzMCddX2bDduWH6zEvGuLwq4nQfWxg3buu0I6JBxC+NI
ILqhdKHJbhq9aWLkLlIZ73+Tm7yd9Z3kZKsUAKFEfuzDyliNLvltG/WmY0YR
hRJO9IBhTbiG8dEsM0MBB6hU07jm/slm5QY+GUQMC7IPGRjmt3Oz1/PBoSzB
BnjAQ9/rut/eFA1Uw7Y5qukIQpy0QMk6tHFihsD1GoW8/EDDLbPDgu9ubYMN
ckoioSeNXYjeDsf1KDFsv/qUk7SqsB+j6Wl8C6xyzmQGap8Nxh3eeYPoWWkc
0f+g6nf3xtx3fWFVyko5fl8xELzmaxNJCnWSpjsusp8sQpTe8VwgEo6wQrQS
FjWhb/7FOOfNOEydXmey7+DoOn7awZZU6yZEHLoPESqaNSDOeXyV0MEh3tmU
eoMwPwYs/q+yGyRuLGo3jsQdcO/eT2Wp/k2pVOLZ+jKxVzyBYl6/Y1qra1MW
bFH9NasxkgPWB05OvMU8/np6Frq4ZK8A/ghxefotApYsGaGxExIuMy5Gi7A8
RPB1sNRcjRkUdtR2AIzvyi17C9pjRCObXobrmHkVACOa/EHllNEWEpfWBPBq
6cz/ol6aTa9tAVTw18gX7GQqnWqwTfh8xxccL5bgWZNagH062KfOc0xdEoFi
1gWtCNf+QPqgWKb2eyFc/Z7ew4ZoG7tWqgrWqgqg738X9u0P4ycSiMy9/+k0
jrIbYI7TDgAT8Nu4OZ3LV9M/p09sustSBGiJ4KpCbiyvK0qbhjxIfYSt4YKG
Qy0+VTKqh7/ZopzYXMRQbw7f+FaOn7rbWDm9QRHfOqibSc8hYntlzwUbFE7p
caISRmx3KM7ugqVv2cujoM6xQ/k2MUz5ZdzlA5G5e1XJSdB+8IiBoR3OvIpt
lz/uUwSXYGmEEMTbCHyn21cYw+CkxQQ7ZO59ZdtdQer8mpWFpXK23XL3K3lx
gB3g+UEfA8HwNurOH/xQ+8Wa/RfenzaMLqQsiZzjGLQI5Z07mPCSOWsP34sT
loYacvdJKstvlR5/r6+kaPAGxuJzkvCsKsUNsf38YQJKB7iHPvo8LZFdMXI1
8x3kKfZxeWjhRTs7CLFM6sQsMMsv6kPJDoABo97h0bPJER1bzPD/PCE872+n
jJWliHZC5vjejxp8l9gWZCnVQB/f0bpWbAjTr7Iv5NIf7iYOBc8fCZHhXqna
dsik8HkF0XnHCjAC/EBjO3R/LoaB/HZDLvFY30Ecsme1njb/msAholDG9M95
m4gcCJR8rLqULFvXcpkslo65PvvN8kKMkJH7atAuDVtgmfviesT+UqNjrMKa
ZEHlnf6yT36tEO7fV0Tavo2XlfM8mlrf5e7GxTVxSaeqsXOK7V6pWqrvnKg+
9CtGq1c8mI1mEL4/0/4vZdclzQUq20NekEbYZ/g4AxnrrT4Yfo0xuwmmBU96
xR1v3d8+Wub6mV5sZRdzQcNuu19TgyTQy0z+MGZfMEN0PyVeacxY3uDhP1fg
gxA5vqiG/adNskTfojPcLQ4w7yeGvxbceVORnRQM2IJFL7jXq2RCeVSOToP6
pQECteDgQnUlr/gjOx+0LN9cSAGj2nOaZinMF/RZmmz4Yz4Cjra48DqVgfGD
XMQRaEyJA6TBA1ot90HvWwmaAg0RiJBlnU1Z2zxFjh+u5otg0NYH/zj+G/41
lKwmzyboYxCC0K9x6p6Z9/lC92QKh0CsTU0HElTNNp2L12tQGm5SgsDrGgga
6awTVzoOEtZ1eni4Qe845UGqIsWhm4Dt21MdRLnYJnRKJUtqXle3gvMT4Kzl
OIkDYARn6GnVwjvCpvTD2ntmB9EJYgH0Ydk2idg4+9i1kK2gmS7bXFzcYOg1
EhJH7s+iQ8GdXn9z276szCyUETCcw85ac2Fq488YSSc7tPNuKrimHtw6GF56
3+R0grJjbk6ZLJdtM5jW7xPLe+GypkZ93V+77omGHpGLPGtyfjBQpoTty+wW
LIMzQyxs5kX9g7FgebkSrNT9wqf4F1nHeG+TKgFW4x42Oa/PU80o/ccp7oHN
dYLQUoihyIMX1j9BBBbgC15nI9qVVpgRhoQkallNusa6MJpZWo+Zsp3etuwf
5wHUOQdLPPIXfjFF2DQchTBbEFmpT2SVo6RjjAN1aL9+rmXvE6RNC8SgcUBG
VDNKySkvf5jXLVRMzGlNsrDDauFf1sRjhacpxF0JH0BYkCy40nb1JK3PBAKd
1PQobEjYRjf6s9zJXnIcuiKY8D7KTY+wX1cd2hi7Qzce5wthJnzEP8N1zBs/
dONjqDcFG5ucFHTgmHKSgEuc0RfEAxp039wdDKHfIrzsDNw1F7kBIyOOM2TT
G4rzWhkkH/h58YSfO5pgc6R4kyREX+X8HXTHLOnpPdUbe/T9222SZchWwxCy
XHdugGHcx15JA7K9SUE6FBrKQoWomrVhYcDb8oLXL1FWzyJe2L4/Fu+j7i66
fIAduUazwwbdw8Wq3UvdoGgXDgi43fScKLc74LcSH9MayNnkE6EOSQI+27c8
vEszijL1h518ej0l+lMvP1X8tlcQWj/uAJCnlAKvIPxxxTl/qdcnF72e0eUi
ihGWR9HKioSZ4laQDZU2GoCUfP3IssuwKkhKMl1spWfZMXpYsTHJZbg/mMMZ
clkNLZIUKEIOJFATrSDUT29NgJhtSHHLPpScn1FqSADfI1jdmf/weANMmZcU
pSD7w5dkCysPaw1EfAtTThpSoKsQsLMA5OCjaKpSe70ccRdNbDga1Wrok2F1
OU0ttY6XhRi4OpnXnWSlV7Cw7KOClB6dqEs5G6GLpyJ7WFTaDbORZ0dfL4zE
CgCGTW6ldB0l7Wgfh5dUNebzz+le5yf6FbuLM7iB8HnPs+is+TYyjIyBIMUO
qWASO6VWhS/3NKSYNpy2kzWVWU7bMwqDlxyI0Gy7a1omP6CP7ahE8WfZId6m
UCmIzYCKV65rLuLeaBpxT/XHO9mvEf3iMGaLbI/MlSu0IM6/ZtK9kMvcaW2d
WfsZHnhmXEWDRCeC0gwCWoW+ZJ8OV77mGZJHJp4xNlSyR9V7kdSYXBBwcB1i
BQzBTUN19GqtxUghL3wo1Bt9DvHnIZ5toM8ImJA7cIkSJaL0gs3ZIfvncIYS
kFDlxLNYcQwXdxtDjlnO3AwNGgrB4cB3uIN7VVjT+Nx7zfWXxaqZ/2ggmThN
27JMO73ROaPcaBJLw9j3mQSNbtK82z5Gx1LlKyXsHPsnHJZNT3m8Hxq7JuBq
pXAhEe+3AeyJoIQbg/360wJYTMgTZWD6M9pZDNnDEgqyuWr6C2OTRvj9fEzA
WIyAItKA7R5RiREUNsbFcuiM5OLwoJhtNpgpzS3Aq5qblIRT2fjQpYNtqfL6
Zcf52z3osxFrYQ01FoEy0JcEbrFGf2AYd7fOKSb4iu8hRji4cvrTClx+Gjil
1hROObeLSCb7mAAQb/AH0i4N/r8m7jJASCpUcBytZlXthk5VoeeMCQVrlmz3
LOSzLc0kpVQa3QD6K1uHql/uW3Rex/HZ/fyi7CwLGsnBC7sWA343Rn2BI/YN
3AhCpE74hOpCZ6NIgDfL+ckYCRWYdpDyb0fOOkeHfm8RiXZ/+XLKfg2IMXmz
Thlt4WqfJffCOhGebzhFCLovjK7rzWciKT7NTyMNu9aObIELfQq0r9Xwo/EZ
Y6o2ZvwPUmZTetTfyIt9YjN2jIx7j5o1gyIffrI2UrYLWgYu12Xf5yrJ1mWv
8nodFEVyPH/O7KAny4ftbDZ4vcUFvAq3VNKZg5mi8BP/s2tmPKf4+GGxxOqk
JGfbhyhzyDrmuiutGe3feLeZ3pfd9CX/87Wu4gFgaRgvozbZnwErVZu5IbXa
pa/MpahZtAoG1Bc8i3WxN0X2q764oGKjD3w1VYq19iGGsOwG5n/UqcwUfETi
ldBmbUUPEySfbP3oxiIOiGvvIDCLauzHtrG6SBCKhc8tOeNveF3VKNcuSNbM
ogi702XB1Ld2wTKpKPYeiX5YUCSLafj9n1Fwe3wP41GQie4tvqGQypx69bKJ
sBo9L0I3VwCroWIUV2GuuwYy2ZZxZWl0PUQ3spr3kvhUIpYyRxLObqF7iJG8
A9hUPQWVpD6Z2eg01OgJWjlLkZS3cEsl3ShbinxsfISlBUpSsH6EBSuqLfz5
IOptzjpQkjL5bgy5AZ+rPnQDnHopMyh+9PRLcwN6IvPOWJ99OLN3ssc5HZoc
iv+Lw6v0ShPvNbZm9Rr67FKrVaJ2nlUp+Fe9ArY5O4rC7qnZNXPSZMKMYQo/
LlDbJ2Y/JfBMkhVpMPmODmycztEvTKa/erWtokyKJQlQTRpnxInf+qlCU4Sg
N1KRKQO03pjvt8EfHGBObuXqB8yZ/Q5SqXOyoRJi3HLUDuBPX5Qmq1DkaKcz
G+J5EAxUP/omxRD0hpf+cL/pYaOvRtlzR25JDO6kY937LCIUAMcTuPxKBlgm
Zc89tLCv9U9jFnHVfV5vvXMlr9D+N9Q7JTLR7ywjDBTWDIE1Ijnn52n2JCTy
tIgFyqBtT6mC9hXR/3BGdbUFQ6rU7HTHB/223zVXLQM/3SWwME9BgMOW4fjL
lSwCXCfIgWN2xYXmnKtMr2YpMihRenSvCPoFKotHRkIW/Mri8B8lw7M4AZrM
utGEOAwkvy6UHGa0wb3VVrnllyd3vI7G6np9akdalBbnc+o8xOHppoLTD6cg
X3EQhKkMgak4sFLh64cOvT7AmqlokGM9jd6aHhR19E14nL9GjItUd23Of6z0
CpHvWa9WgHg7/CztA3NqPzlAkgut5dmnJFVRLfVRmrl029A04BwV4w4HFTG1
WgmT1lq1ivjvL1fFVObBfVegRuTuzbYBjisfw2iW9JnW7vx2SlzLhLbWCser
ClCohnwYIPGy7f3BPhdhDEBYMMXh0mprZ4+lOYALM1RLtzR2OYQ5QL++wWfd
d7nZLxippDIRqPzCMpeVtV0MCMUaKVa1qzjoc45prkRZJEMrrxcRkoTlx6lh
224V9MjdFt7f1w7mw0bblGKG64O1w9WfqexB2emHLCDUHOAk3lBmNBp6iNB4
QwEfR/BPGPfhjtBMeCNm+El7bkHGlr/SwscDVKjSJb8m9OMb8Pvs4Ywgw/8I
ZwsRSAcZgXIVnZudQPBB6voL32Qs4iI0kvv0UgKLsd7e90Hr8yFJIIkmTOJE
u6PeBKXyw3GKO/ggHSpyTPyjzV06PYDLzjogZfll23/60zcycAM0+vugbG+w
AukwU7vuTRRAEQvSywRGWizzIxZAT5bRrrkp6JMunqCQh8PRSC82kxu6vBQA
Ggq69AD5VPZYP8fIoLzlTGCVQI/OWPF7/uTe4IuJegjMC95BviFXWWdPA5kp
KCwemZgbmyMqS9otCSXlILUNJFkpM4Ck6POfhcLcJJc4E+1EwNJlu/gRGD0l
pHDR8CfNwy6ANyW/8fTwuyER0i2rmP7DlKz+CahMhM7ckeMBhn4i8x3EJ8vj
buH+5owCVJnlbWkbrvDg4ExwSV4z3wo+DOgSiqNTTxbjBzdrwoVF0UhE8dSk
cugAhMIcwn0koI2qZcUTBwtQH5i9iOUFqrD28PlwZehNHPqTpU964GKJBwpC
ZVbywNa5bhIFFEJ5FZ5Pq1AQ3CEUcZMlNchhY4W69NYgWQ6nZDj/KwQdY4Qb
BMpC7GSJvmRM0HLQ1FJSB5sCFAHsRSQl4Xna4r3gjFkXhgQMMpMdOIGuMLkj
wOCZUQVBTYxoFdzz/0q/pxTfwBj8tPRhPMOAGhpfLUVaLLlsXrG4Fe65eQ63
WWTuFJnvmg/mzj7/3w4TJ9X/rqSF61uu8QD7JvwEg8YY4Fjn/6lQ92Fh6cmn
xpqqTnb7OCSTGI7+KrXcZwQfdxPG7WAZnplXodcqwAHF+XzTxv82dCdiqYKl
5JvL+j6ptlzhTQXCPPVNq2GYBI9UZx1tt/XK3sI1ufXPZJMwk2O89LnRz3dK
ROxy93v4p6fDJ58h+0Qihj2eOw8bLLTd0WI1gPvOkwMinvCcEOxDwruzMpw2
OTAPbQUK64TSP7rGCOWRSqNqifjhQglgL7Fh4hZzPx5/PDwgkj+GHeLihMSe
FtKiPAsMWKVuqI03XE2SB20LEbtg9QL7ou3WHdJjEHA7dcxAELXd9sy6uZ3A
ejFn2k44LtyWkQ6sZD+I7w8VhcMR6TE00jlAyQaOOCsaCPH00WvWylpcv3js
BX7YKylAGBCDtFqjCwaZUAVy9YpwfG1gvj+k9hrcL8KgujByy0x0omD0cBWz
NItL/Pbif49aha52kSozzMPBNNgemHRudPgSbi9AWtdFOnfYzRGZ6oK55jbG
dpa3K26i5DnFerB1VLdWHkqOQnaX2V1NjsxxaMU+AOehaAic5DA9YGHivmW6
sHIL8Zn32C8zb9FkoVtxv7z4l4FG32f871vLnFu0Z/vrrp8njKPDd04o8fRi
JsLM2mbqV2vR4hN5T1z008VqI++JTzlp/9sjoiau1EVBKqG/+0wEtejAnRHr
FjKFtSTJD7OCGCHMApfQSjP4zPhxXlDDypchtStyuVGaFACqhoalVYKtIZVu
3Fd1GiSTdE4GhhQjN+6M7R2djn5wC0N6HDZDO9Mj+rpNp/njv18QEli0tpDZ
D6yiWAGkQY7PUQrIiTnwAM6b/iBsbDFNMO+EgoBBfeykxtTjKcxwYLA+eIHG
ezMAxLOVcm2bjvMk08xHbVGLjUZUqanqLmZvmAk4Hvfht9r/WcWKf886mk2N
QZ4nBauudOtWbtWMSnLojKJPl7wQkcfGsxtmxGVfhBlikYp0qYZAPrhwxToX
f5kFB9iWW2EHFLDxbmM8wuOYcSHLbXsTqqnFaL/dXrN+4Y9W8PSDViTPfe/F
5rx2T9zYtuRPNDDjCxoyWFicSPjD6sOel1Vs2gcXxO33cQOwr2x7GgSYwb38
yu8e+iOAcYOFBcMfBE9WigYqfjEU4QLCtjyJUTmbhDi2kj76rxdK3GOSRRk6
qf3j7lgUSgH3AG1HANGDxjKIg/7+ATYagDkEchJ3Fg+FSlkUGFuYtXaIyxHt
c/2jPCtHYYeSpE0iKFk51FCXZbMzaWx4ZIj5Zpc4c9xGiztVHKff6LJDiJGZ
9s+Aj/1PYM+HIKoutOlmu10jkIlqqqj8A3pf9+obw4CuOhHJ3e7Mhm/Ebdhh
HTIU4a5fHuVoVSDqRLyLArsl8/E+XZm6wn2ednRm69BK0TAzPwz8XdvZq8p8
YLSSfL+krODfbMGQ3ZHmVUoUB74mMcKTADU2C3mr3tzIsGJ9BSywWaykMijg
5bFoUxTsAHHRJ4mzazncbvqW92O2GvPvV58upO8z5YX/5eo4s8zUoU2ncoPL
TkBXlL+rGvrrCMLkIg6u2VEx0GXjd8SNB5C3fKs4wmPyrySgZ9+dNKNo19fj
AZ0+yP48LYBAe6yTOaU6XkdhyzV1EqRDWpOGStDbn1LZAuTZTRa2/+2GiyDK
/u1sXiPLsJo44D8PDj61bH4xlzE8DURJKzcOK05haWetk5z3KHNNnhgQxjUU
itsRcibD6TtubSZnTAc7KBpOwdVFdGhgQkYCuURMK6w4cpahBmi8hAEN0AIL
+oGgQiwAduva8woYjEDp7dPoClMcC/QA7EY7/DNfWBCh+RITN/s9M87cWNtz
ZNHpSC6LnTyBrDoTa8bcQU7S7A4UtbuE3pHXA6f3b1qW2DhrULbnG9QZ+WjM
RKBonpRuMx7myAH5nCetXghoRYrNkihFN2acOGYnVIYZYEzqkTitTCccH9q4
pd5Lq2PQwkC6Tzc8L3mEYppQMPPr8CYFH+3YW51fQSuE6amwrbPyFHC8Mdqt
STXTymWG939gw5JIPY/zlN4wzohpzuKZaSsTkIWMZ/SnqQiKfHfWaVBbSNAd
aByAhSLL3M43Hw0hV+MNxengSt/oc0iJUBiK5CcwGSQinypxe0ekiuSSsneC
e8v2qn3MO1NgRQ31D98Nlca/yAa6JgLyAaVGxWtSLsG38NoGJKHaq86yMAvf
5sUeHWbIKwh8amSThEWjeLlpXTcIbpucYSfox4jQJuQiQjUHWPPzS42K0VE0
uQa4uoj4rzWDN/XwoJvQ60V+Oweo297BJa1HFSsqdCafBHyHlS1eD3GLvjx+
6QUTEeAoPYSUPKksGCSUzVKUrUePQ7TsmElO5On/K2uRXdwyCtoNnQBsBCyz
dOn1m2g+qIQvZ4QOHvy43DkTKS1rl6k+cSXbpECJq/4pIZtDqEt6Evxt9M48
B3iEHShAd4Elv59Qv6fgWgLhI3nmZV4Bmx5VOcDOlRRg6ndaSaZ0xCiajg6b
eVouRuCvnPI5nQ0Wtf8B6NJQtILNTTJKS7dDd4p854GuQ7NnsLGOWQufxxb6
yallkDENrmHeFiY2kOMLtOiV01XrexYpqyp096BsXZN9uOekVckuya8eQoJh
m/MnJXYDqbOEAAxr1oB+q8k1t9Yxc/6CX8hO9y8PyZFVBGQW/n8B0PvpIIzR
kl+InV4L4zNzB28l6HStaI5VOdFHucuM6UeOXP2OyZVSqCygdsaj6YV200tE
qeZGYHdxiqoY+dZKjtGFI9OR5Dct4zlzTQsoojgK7MACuqDSNukdVItZlUVm
RT4zkNAH8NhSUphLjs2OVmIr1o8YDHfT4c+54CBk1dhtZ3mL7xfeFCtKT1UW
wX9ubhQrfV2NOQl/PMC1WwtYOL5heGt7oy+c9a6Hz/oLypyaZ6KwaNMkve1q
VHCbqG3irDILUJ3wJNaqCBRoHGWJEXdAWPPUCijAG0yQWlB7zegFpk2Qda2m
GwKUzCVmVU8fy7VpWPKMlnWE0Kv/R9En9gtjauPkJhufdvQYCFGobTfv3qTr
6T17rC7jZVBtXbfeLSSURii2qkQKFhnrq9UOn0AMVwvuVNA+77NpxT2xqNld
REAnjCXumaoWpO24nNpaFyYS8reQkr4qFu7QuL3NRXPqsCAw7+YhPsaudrbG
aoGANsywhokNQNr1b0O3eI3lZhiaWv1YTw6+QpG5lzAeh8IJ/yzfm0uoWIZE
0opqlv1yo+ntD7sz9lquGZm8NSKDq+t81+02H/64msaCczM6FhcZWjeWj69Q
G4w4uP1hDHMi7YuPREXJe4XFyDSOfG1Jl06A0v54tAUuwd6BQbU31I4fgc09
THGXQTHKXWRDgrF2ymUNrfGbganmcP+1WbdT89s1hXSDml7t2A4xIyWRGNLp
FY9XEq0Lya1pOYWjJHrnsImRLYK5RaQizVbokvY2yRC3J2e3mYoobhQZbEQH
ds8U/Ysc6qLW/PTQeuWkgBnLG7mXDRMzsCmdUDQA9x6MVQcktKYO4YQU+nsr
j6Gw5q+RUWeszSWFDPFS3748Uc3wy+GKXJrYwh8qYLkphT5G8ryemD0ZH7S6
yD7legnhGlzljEmMicxGmJGAKBHRaJKJ2quJtjqGfHO0pLzzotBXzViLCn5i
FkBrU2ZTlYUHnaUSWPjtxGDUxwAavgII7g9h5KY8K6g21T3AwVRKiIa0+9lf
Hp7YsZivXalK5HABlCbZy1faZLu8WIH7u/zlxraa4CQfdfFTFDx2CjZ3htDk
xL2NQ7Czb0tT2WJ+uhwiwiMQ8ERPMzwYqcbzVpd0YkJs+RXdw1Ly62xPin/N
cF+rbbRmmuGmQ8ER9bHGd8jRnH1K5w4To+Gu/CSdgXZpZD9gEpPv2AZqrKFw
c6v8nDSVFHwdm7jSxzxIs4sWLzZnfmKT0sQ3wcAHk2WQUwE0hFUdCjJYH+lV
RrPQSkgy9aKaVj4tUUfLQKhfXqhsSHvNprwn7N4zZVH2T1cZG/H4hCnQTLBF
rc6YGizwuEQkbWiu+8mv+X8itIo087LtqaoiityFaAa0HijhLzLiVZr2+vIK
WPO4TNnCUZlw8vuHOhYQjG/VFVVgxCvAgzjfE86ZVe/rBYoOIp88PaNAjW0B
+RBlwFOSc2nux4jGkdw0ArsiAmnGGl/CUIz0SgLHhzrh5Nml0xOjM8mzTr4r
m3bhFD/qv/nLddT9mpSiej1lC3s1LxY24fC3LdvhLwYHArZlhlV7uixT8dob
NiNfi0opmk/7oLA3qjsS/+CNGF5S4P6AL0kizDIlE90fBHzvkwaIvkHimPk2
PSpT+dJFB8iByYBj366gDx1nbqRt1RyBdaJM+B5xnbku1KubDipPjJCFLkhT
FDNscU45f9G1ew/UsAJFdnjw+4SOi/UeLdPLUJcN7JPdg1cbxUJBhsKnBvwy
9uV4LqsyC8QY0CLOj3f9jikSmrdeo4S/MOBjBHZittOE+iIcpQ7l5jkJ5Oq8
RaKeqb1Q2p+zkFnLUSXuHxWhsl4C0qd+Udd91CiuoPUEezpbNwTdOH4+rBJG
FrCpW8mkc8v0ZoHtNDfHWpGLC3+ILSUbziNQwZse2REvf3mTLE1tgOsDGgQk
Riv8WQjZhRTSY7QLYGHXG76l6+b2HR1P4R9kVSqwFhv2PYxUb2zFJAHvZQB7
uslaslWutUmPaCvgWypkq5Gx9C5cJ1+MlXLdB9uA31mBLyUMk7dAeK1Gb8nm
VCswM8qBO0ha9DBGaCT9nwu1ow8igsEJJxepkekHoBackkmwWqFAVGIUROQw
33G4X3gmfjAoR3U0M3OVkp9RgmKuklEY+/EAtTBKKbcN6zQ6D4j4vgYt3CZ7
Oc3xKsJDU8cYGA/WIpDbmAmYA3ApqPPIHjTVlos1VkaSDC1b8/bu8NdXr1Vd
6pG6epesO7o2+dq5y2bTXcOACkPwE8+rsqxwCEcmXYsSNpbfnFgwb3UPSHhE
BsNMt4Tz+DepCF9ToX54MSMSSeYZK/pu8RyQ/06p7dIyqp00cnDRyTgjuXyB
7lK6TRTbMw42yb/5F772MrOkh4f0uTZKP0HYaahTj7NbL+70w/CjlqOcqvXR
w15DJ2Ao6MyMW9XAzOq+DWTEzSoy21xdf8Nc/FSGWnaPh6F0T10Ih7jNGi5o
1SFeIQXfthmFbjKccuz8I3O45x71ZykcniYXajhDFFVbAb33vSieZ5+zW0C7
18zt6mJUiw5CLH+IT47SmEx/J5LV5gctLqGZd6l0Cwg7ICVc8Dsmkg5URJJf
2V/k98b14yZUnSY9S+z3HV9eaPjIJSnMnZ/knNwkffQi5cns1/Wp7t9ugusv
a/ls1TA+huFOEENhb3Cgguwgkn9eQLdnDPJ335pIEznzvlt05HsjAIRGbEnD
+sgUK5Kypvs7rCOduzKLJnaRtJK9CMvD5nAfTkO2SoTs7VliPC4m4a0m6mqq
Nh1IeseR0kaMLl/3Xgfa94AyDjTPY4jdX/MXnKflGwsw7Rm08E4m5FZGsuXC
0oSi5OagDxVk4xebbinK/9BAHeK5XGJypKaBg+peZCymT61aokbyJyATg+bi
bBR4cKrtS2ISwpiuqrPh3qPsHFCBwU4I2BRKzAsrirV2iFUnmIh8Ri8QLrtV
ZGkDwR159nbQYyetiEH+XVBD+CByOia70v1zin1YXVFbitkmOXdYCsDvFoZR
lqJEIOlx3xpwjR8ZBJO3PqE3iRclxAapT9nk0BXye/PL9VZHEDts2alNw/hl
/T3qCqtMk7q2hcMZIOTh6oFjdPwmmPNL264LnWJqKyxF7Mcir4mKiylnc/Mg
B5y6xTATCRSV6qEG9AH1PS6ymz7KkoY9jwQZ6B8fHT2K0o0aI0eoMgxUQwjY
gXGz7gGg8gYXjnLa7neBm+pGuq4DOb7rWrBFip0P6/62TM9MX0SEMbZmJ57x
XKn2ZBoyAKfIZB8M0wi324nZU8KetEk3BXxzGd6dwP4MIuh/MuQCBSW2jYi3
T2lihkQH4r83mwTSIHdlQjFWZej8k1LH1/nW1XGFopYaWW3CfheHZalh3dfU
OC9+Ky+KGDccscOGpe9n+knczJwXzf76pjMqQt+3cmX9pCu8S2JInTJ0YacB
ECgirBmUWkKl9KrmXJfbL0RSvYiCciKRF5M0cPOsODQ8oEzjxiO0PP/p7vFX
OPwQu3KIbadu1SGVbgHMioCr7oil/CJuSf33eDNhJyJiKrNVrcHIDUDccvZ9
9cQIu2VSTHotAC06AjLBi2oDWkJz1f3Wx6aeoFkfWjbDYhvNIa/j/kOP7zD1
0R7+OsB8XH5yK+itFMO2diBGomapoRX1oW8ZYUVBd7fxoVeB3EVEFbMQpH3c
jg34TsItW3+Z40oH2u0Xjl+41t55/7MECN38CD1ii48h/s8NyVOJfIMRlFwc
fDoQlQHjM7dEYlcqsexHFcrD/MEnudgeCaBOg8uji6afKTvClqIrrsfG4WHE
0XLIXk/ox/HUCThlxwGZ/DhScIZJhkSHUppJ/ISCULoFw520KxHLepBIBD+z
QXn1iDOAHFXdTJsmmQlmkiy5Bb5tGBfDBvQJ+Rti2fUn/aURlsezrxNxdQlc
YIaPye87Qyk8VzIk2P5Aeu9yr49B+l9o7F1aR4YNsT1Z72IIWYwWi4c1mQtg
zRYpc/J7L1JxiTdMPJV1asRC80yApsIm+fVLgefmymay/2vrt8jH5v7IKxLm
J4AQTHfbvU2MS9w/gpJ9JdZHtkkIaq4Ka1iqtYCXNjSQLiXsiJBDYOGpend0
nhvwRORHjE80Fw0Kd+dcXy9huLC1adxb99UYQ6UEiH0HiiOqrxWvvF+QqQHf
zrZ4lkWX68Qaq/MX/LlDu1W5agJGP6ZwGatqQv3San8d87z0SHNJedfFdVfS
AH9vTvUBlb9PeVjmc57mXq0Pyc5fZnoq5KOhTyW07GB574aXbI+WLrl9ituE
l/mkRwjB7vb9TsbNVVn7zbLIVdeeay1C/9yWeqcfq6joDEFByslDUjTlLJjS
yMS3yhFTlCL4ac4o92tsBMB42C+24wyUaTI+XiuJZYGVOKDkrB/YxX8+8Q+9
7qiLmqyQF6bUXnFDruzB3ByWxrYQGj+XJ0yTGykx8RW/gckUeAYbd5Dno3ms
MLXrfsGiQqaiGlrlM6RoX1gG1hyfvAAB8C4uTu22C9/DuEFR8+ZiRxwilN3g
zzONkF7Lm8iMuPZIAPiGEDMo0ctQVGSLjsXnr5y/E36dlxzgZzvUm9iSYjXo
jO+csEsi8bwB4aknM2BJAVj9G5APlG8P22J5UxSpsZdtr07iZvUKtw01Y/O9
Q/8YNP29mc9VfgfH/QGGrbSoa5YwBC7/E3wuO2bYE69d5RrKx6UKtg1ZXvo9
EbqEAbVLdNwNlk+lTou571eKmXvWS/+NWCIumy5S9fkKn9zRzAAXgWbiXreb
G0t6nJPJcOZDuZK7q/RWUPpmfT+oTH3ZCdKoYXH5EIQrV1fvEN/g7CLSE/c9
sy8GHcVnXDubV8jyAd/8YqarEt5HzCYr0PZ4OSftQ/wrbWDtVx0FNpWCauz6
0Z5JoDGQw8645h3DUkslIzwHBGP0v9LpQXFtP1Y4ZEmLrqwEzLLljFGnk1lm
mPA6c0EJIND9r4k2IxiN900UR4RbvU1j0hUAjZ6+zoqZTBWXVyT0rJj3Nk8m
+rkkBs5h4H5n2lj+j52NHQaqk8lcMhZTwgFT86PEGAWNlQNbCX18U0g+EwRV
ueofNzyw28BteSBSUy2OH4QZkgFcN1d3wVtZ/BOZpeYgtCEix+k1gvPCzYbe
+0MtMZIFf6cOplr+uKmBIZiIx0x1mwXKGiQw44BUVC/3WFxMGhwWd/o7EHyE
UJs0FHWW35AUfQFCV/8XEH4MFc8RIdKYG2VKFlCnK+bWJyHcAmeanBaraO6W
NcDG5xjTm/f5US9osm7XYZzAv1dgBnQlmsP213vO5Mjtedn7ULqFka9T+FBK
KvT3p8FNRAiJV9eWmmTWb5fSACeL40jMUl/nylaNt2u/aE1POCbj2jdWq+If
2B4x5p+ouSXT1bxN14pVy2kaARYMdAsvPB/uaIid8uw8I63MtUzdNGLrsYDc
ywojUX8HhOzSPFZiOxkCthxR5fIFLCk6m/Id9tIG2Q6Z8mOXkgJoDujCn+4l
r90OgeDuop+2I6zBZg/533RkDsdT/JLTPH8F7yEgr13nqgQL1P4bjo1VXMv+
Oo1wjBAGn8W02ZAPBhboHSwIAsximb2E77F353T14iu9YrX34t4/T3LEWSYK
hVM+rGf4poq4Tpg9PROBwS7SI3LAzqhesrRYegMS/Q45oA7hhh8mLxenVNAN
0htszi+xDcHXucUVXdaR2BCNb/0M5hXDlhasDBgxe/+ioPXd2P4rWP5h5CGy
RYjBvvqxNXW7volGTriP3DZhfwz29NGkYQDMalABN2NkkgnYpdPH0O+vTKZ6
EzZbEpYqPDNGuDOrOPfFV/IX6if39EOMbJndFOgduDx1jx25JsEw+1t1FzyJ
C0jmLgmGj6iyVfQKu5TyXB+ricfAowHuP+BqbejhStEAlHbbNThDnI1aUDd5
Dn+jrlnqD0jJ5jLxb+bsn9OCYGN8/mt1rBZa9hAc3S2wEo+lvtsKdd3n59eT
AXYR7/usl8nZuipQueYlzBM54iDp6/3QM7vHXjq+PHRVdHqoZ3p0TX7zP6lk
EucplhTtjShb0Rxa2wO8MiKPd2lLD5tBMFprOYNvQ+FP2G/QeCrpQtrSvHQ1
ina16FJlKZ1C7WKBMMCW9QW1YALZZ6Ux25h+ss7nz3oivlZ/5Vsv7byJwb1d
XoHEPiTmlq3xfEqqvFid54wzd3UEb+jujCD/cayQPRCIG+Bc2mQm/DQ48JtK
m0etea9bjC1fgouOsvOTaYc5aUrsFFx0K2PENZUaqN0boaNkKekdNRYFzsOi
4+q0pVwWQfb7Z3coFO8bdAZtZ5WiRCJEhUyc9D5ELBf5ii0I/1rYe/DY1nbb
uZKFNtAsgWhkY6sFASSlKkjFyKZTXliWLGXP80YPf5XvIWMK3RbFdQb1ZApl
o6vSqAZ63QSvKLJ27yJcVdXU7XmELh6HBrqrhHgb8IBtov/G9bZuNL2wtx5f
e48i/kBF5mVGkvNzb61h7s8uo5w/UdlXSNC/neEs/PN0JfwmwBmB0E9QfLOl
3n9460UU1M94OPM3wv6Z2WbnJ9eNDIGH27hs6W/F3NqEJ+C3W9uvV83bxB6b
jsa49DdwvZZt5bJ0I1Yk+eGLJAqMp+lc/244wg7QSpOhbQkVLqtByewLKuJc
PVWI8DIZEXRcbX+2JbypDjwkEfkTeu5nRA4iJJn3qMinZ0i9/6nMtcZdUh+k
YFQfacko+8Bpv3DYhqnZFiX1iRqIlUHoNfRz47mH09u2feEfFOxZiZoxz/zF
ctlePbRLM3s7HtptIahdAi82WQxHEV71pRJHvVr3aPq/ZdB7F3dyqSqsXifP
eOC8T676EBE0Fp0mE6keKipeQz79zFbUgicaYf0v6G4wE2r+XaV8rr4XqJZ2
Vepuz+sGSzqGppdkVGZdVKo2kIgGeYTbB/RrdZU8TeiEGPHHoobCjrWQRabp
5obW3NdWbaiX41Gp7Jd70F5lv+pzuiyGBDVm7HOy8Llh2RxoWNzq4sN1qlqC
ZEkh4axL9Zhrrs+p3wdtAV2qHtuBX99Gjpg/mvlYqgjg288tmRbeE2vuiAZ1
EwcpoCVVLqay4+YapLFd5SGTCyCsEj7OjEHNbuBlf0Z6SJxQlNNmW69zbkvy
zDi4CXuT9J1zqVMXovyURu95uIix63l1LXLfiMLAVPKHDbXXfXEn3rCLDMJg
1G6IDvQ3/nge9m2TBljZhJA76eALWflc6cLoRa7Ln45mDycZozM3ivA4ySYq
4yJ9NDygIIgxFrOIK+MM94VfuldsWTt+CLdaooWz+UVZzSfaLPHjmip5YYvh
VkJc/rYsq7lPsmIX6yFFIsf6OYrHx+pSfSirfkv0bFkwE8mtbT2jAMNACcAT
ZoFvfi+/+7AOBFENiYMcRr1HClR4BW2Tydzmm/kpWB6qiC2/3BAcHIHfnpuY
gP5mLvbXVztVsazTJnXVrPeos7iU6ueOPrBEOtkypoUxsQZ9UmGs5JKvsChv
eoaAqPRkSpKlyo9gHFoHW3OBDUC6CCYh4UNLzS8HZFGpkDXDUAzIUz88QFjR
8Nf7PrS7VnFAyZn46zl5VFuTvscWVyBnyBtD8nmYDLgrvKdqM/YQK4SouBYq
bzh+GbM/Bx88UnodJ8jdECc55Kis5BRjy/AydH6Uo+Z86tNloyG6q6jl2wlK
WVNDHlA/1gA3J/2wQ8IBQ4pqbEJ5szHiChE1zO79J6GUkuKmvXrA5qeJtGhk
urTHjY+5LdnBgDDFFknpzuYZDp9zxvE+HTcrKitPWQKdeEFcR8mUD+RZzrjH
5iEPERge6vmR/HEx0PNJGuXx5fuPJ8NPTEKCYC2FpbMzeSQulQ3gsDDd/Qh1
AjqMQfX2bn1hYk+9Jj3c3sUAulxTqpHL53UrwY9XZE30cDOVdQYJHMKf+hqU
bJFpZ5gIn8gjUZibtBnrXUMyc7c73tEuoQ9HAkVwOLYXnWilteERJ2MJ6sRv
GxbnJcdNYpUe8nsDpiAsvOYMG+hVySKw7OqKfF08c76RPQrmmyEUvv08iaHJ
RJ4EfasuLBq9MeaWNr+mqKLW6ZDUz+AlyYZq2uz1fyFPWcQYCRQZi88+WMlt
NVMhkmyIYI9aeG4H+k6P2ZYOZeXvgIzn7w/Z23e1+f6fE/un+LNMvIkJAdm0
Y9alGEFpPk6cN9pp0kMFDAKWolrbp6/jh0fMeMM7wcqZFyr5a2c6wxF+dVDw
rIeGwKqgMtGmfdvRy0hvFeWfZhRVdWD7YggvWO8dcTbACYGi7AsudD0pje3H
peCjAUsnvzIHGXOw5Amr8qBHd1jfT53SBQjLDfeKF3bRNP2vda1e5EZrDARd
P2TGWWamC2oMqR4oqc0kvb7dfNCzhgBpOFW6f3X4p48F5baNfFhOsvwRM2Rd
qnQ0QshdwDO7YM7sWCY839eN0jU/pSRLThm229VISOvtxCWkN9FjXwi9wLnN
h7BrWloH8lCq1sNaFMYTmRL9VX+zm0VMpbcb/dXNmNCsLtBEmUNeCHjcDZDp
3Q9SKizjpt23sR9FI8kEKIC+C5Fdxkv8xkEA1ZSIy0VWwmI8moePQF9D6PLk
Rmm0UBVXpCn9wsK7rBgNMNYjBOtHX4RECly+5yvInMObZYgR7Khx4vWZUydo
FR5aPQlekR/3t/8gPbaobfBCkw77z1BUcTsqO4iOskzxisoQRjQySFogmk/O
URsE8wAewWCybJmTQhweUwskGwRbVzVMJzIw4TwHl5AHCaAF6J5V/RAmysQQ
D13LU5XDfjiKsrvsquMJvlloUQHBc9MM5AgwJMiVNQ2IkjBDOqok+zzZTw+b
XBb5SsrAOuwSu521/0tciBvek2mCY6qMSBotZCMm0CiT9J2WXHsiOJONtRLM
5guAU4VQ0QSLK5OQa3cUo6WoToARjRQuPg9RLCq+qxgk9SpZwwVuHdaVt160
6SFzu83qqFqCFCcroeDqJN7pcKlnIWlNUYTWULaEZ7MRxpqMDAZxnjlspERg
XcqJ7K8OVIhspcZEFq2tiMAAjJNG6iL9i1pYAe7FkDUIK7BBawXz7PnNQ2FP
eBewll6GqGQ14Gi1W+WMfGW6l41lHNtGshjqDaPR8RUKYrKbGdNRHocYq4Oa
Q0h6GrkAWz1c4qoiVTob3ku+D5lRs0j6zZm6G4f/hA8+aQlSdjLQ2CvtjUaG
HYr/ALsOzXgZXih+R6oMa7XcqJyP/KhROYGh1qOqUBahYrlkzIZpS6tItTwT
nK65RfWJR5yr/MfzJcPBtSFHNkc/xdPb4DOlyVWm9rKrlOgpntOaADlr4bZ9
NfEpe6eESt1ixxuRNymkCajdg3JUYOS2CNrN36SAgp89A80dE8o5vMi9vjgh
H+1MLg6MWIho4tMN55i6lZIjH3HB3rMqyDaERGxGueL4Ntr+fu/IiGMYL4uq
Zb+jPOrfV+L9U/rtJOlH5mjgW2GzAkHPQGf99uJwZ2Swcc/s1/JrVUjKGFbx
4piykJFdc/wjzJUB9B79ptyMVma5YSpL3zf6LoIYmhB/giTYkOWQwL5xNzV2
yp6El2gM5ld8ZdtLNg/V+w4kELREysOahdJ0otwkOoskNbA4KdSYGHcMwMei
HHta1rpFjPga/N/HiR7wSX+dX3w0Xbqa5Yw47a4wsseRtL6bWWo/4XlU8Whe
PvyG6RbAKXJOTOGAZy2y5I09DGfD4f/ZqrFnD35aJ3gAfoIfVwDttFE0CXGg
rK9WYmaUTOUmsxoRCAXZsJY1Kjh7dIwlvx1HkhUqtAqTEFKvzo+3IZ663vc5
1Z/vrnbD7nVWn3NdyItgPNutG6MSy44LaQ4VxapnyUU3Wfda5xNaQ/1zhiIl
EGCtFnJd+PSCX6EOrSCBZzZgce/j0Quf9wrdBxcBdx/G4JOyoDLVIA/TspgO
/SXN2U1wrJ9lZzgKIBiKPhqMlRczirW9+5CRwS87IWCB6fibTakj8eZDxpdr
cS5lPDC0o4I2oglfufB8LAL5JBMA7vMu0k9QPa0dICYBBTxAu2cVEI+UU0KX
1tCpOyhpGTz5feP2U31GXV/6HuPV8rR8YJax2fQh1pR3yGsLsRc3Z03tNDNZ
3uaImlJJCJ6CAKPpg5O1RVj5lXhUP4ibJFWOd4hi1dr3x+5ohHErcwfoo028
+Ehu430UyDRTa+8Re6GwNA3cRiOqI2g79/Myvgb/KkdFUCAaqm3k1BkK1r0K
l1NYwVVgdoAtq+olGMQgqgms/C2rD/IfGNHmpUpa7wcop6oxD9ELFgQLjMxf
a2Vx62RM/UgQOndLpKtKmrD+0jJvCEo0GQsNXilJtxx3A47v1HV8fZuLo1KD
/beWdEbpvIJ27FVOhsl2d8VEN+XwrMDy4StFy/7aihKNAO/zXh5C0LyasbxQ
cva9JyLEZlTp/GTpFVFQ/JJiaigm6lkOqagkzun9PIyWbtkOhFH45I19n2T8
rXQYp6K5Nv12ZjSD4MBiY4XE+9cEXsKa9akSv/6uGcpREi1xQIMp2mSfE9Au
GjXlLGo9oil577fv9jWvU2wiFZ3bxFJlD6FQVyEt6JReFH2Vlrnary6mIiBW
QLPBm5rP+QMkEl4Q0pZqNGloV1oTl6k/lPSGGZSbpU3mky1SziDAvLMZx06G
zIQR5sI0zvZf5ksn99VWBJhi0fkGODwMkFdjwSF18f3ELXBQmlKZDAKb1cMx
25Ym/jske3TehqZIvVoJXe3Ke21iYxDEQonQQIJ61XDSs2xdw0PzC817uFxK
6afW0vkwxYtqH0MfRGpJTmHZmud8akDz6nHtJNFMJ5/fsC2pIQHE2gGtzUof
O4a40hjOcwYyyeHKZml1mvfpYdT5WYp9IIfS964M4RseWLvNvmRfp1cENsAS
To2IdG752gZ0+qJrP6jFZ4cy1aNFLCadACTPOur2zoKR/HEKUC/QDrUEynLI
SOPbpNlfStsssFtLRHryvzZDvgCqiR67w8qI+2GB/z2VN4qbEpGPkkDXSjjQ
gpXkT8cPKMiZAtNHOIyqO6j/OjT6pI3MqIMdJrJKQ9lhiGDiZHgdSV4ndDCH
vdJ0kDvJbeLLznc1ICDAwmfLRMPt7ycfT8sLSWnVCWZzFnp3kqSyMzr8/hFp
iKi9ZblL4gnzCk+9nvwER5rH2AktkKIpDqi6ahAxzEDF5bC9FoCC1nuOOfZ0
GbXbq0isuotuU60zZSt/qBqcwb4shK5/kWnMyKfpnBnlfoJpQPTN+lfXnST2
LlIshpNeR9vRjqQIAdFfyRYQ8KdYwsflL362FDvdAjfKair3plWyItYt6Xrl
9bq1JvY2om+4DmNe/lHa5BSkxkbZSz130cgIbX61tlx41aAl3BTDL8/rKA4I
WB06rV+QEJzwhRVHYlIcPG6E4Ml1yIlPZGIiBScAsmOB5CUTGKmr3+8/OBen
rNggp/ExeDO7ayGTc5/LBtpxTXGshgVuRJ0V7cpNi5c+ZVAQex7bu6TGAUPq
zAYuwDCPMpEkmcRQqQwL24pxBwAAlt3GPPijD9MbHtPQx/dJuTVLqIUvDE2L
n81lQzCkcb3SsRQP38V2r14V5ydHG57YoiV0W95yIi+dP/qQ/gnBk/OMSa1O
v9T0F4aeUNJ3nHnCFeNeqiqPmlSm2cPKOzJ0v3HtmdpfSgqCEUBnuwq7F4gN
hwM3gblTDlYjz4WUUguMPypXzDXJZ5Tvs12Nw5iFv4+b7PH4qa4Sjgd9lj/3
LTYu/U+xiJeL9VbyBdY55v/FnoV/yegv4r34WUtuBx42TDBKR07OQx/XXmiP
c7MGYEXVsJqoRzZ7iQLfCyS8iCIuldfNLYOy4WBoO/DEn85mOLWc4U0+2zq+
oelpzSkfgcgn4l5cRhr+p7D3ZnkWF8TMA1WawOojIuclVekugn+31Pviipx4
7+cE7OJIadSLssxoT3mCR/U2sX85rIoNGMDa1x/14PjtcQ2xtb7SKtFYUu8A
MSt9+3MTDXyHPaQFQdH/LhkfEGdEGpJKcwr7dVrIB+49gGSF6SNsYUsUcsmn
2fRXMTAhW9hGUDO7BuqWfiFLCZqYQLtlwrCB/NFPaVAZ6+6mNbVamDF2orVw
xphubPe6TgdlHA9KbMSDnnXn16KNwL3z7ZnsGkCM6TeCpOiD7M973cUrPG7/
VBaMlozRfgiF0hCHKk1A1hgThMHhHFcxEI5pI4HtC2ylA9jjgbnICDqXg2I2
LBIxZgAbg/4zvdsk4/PAsxD2OGQkh0ukEUokDtAVMPTBUgh18RLK9BQ412dd
emQrGfB8zYsVTDiL660kQ5nAHd0/c1GoiUUEf5Rx2AVX2TSGzesGIfqHruCG
35eozshayfH5IJlT4RAVthk26ReMOGjt8lDMD7yFq7jGD4LXTX1CXewynFq7
iJiSNtCwKKWjJrRXszDxE0eIi6SCpgwqzc1Hkp2jfSpOzFbr3dmdLrqf8ZCW
tVIZ3kvTeXzMD71pQUyZs8hLUmuMSBjU8Gk5ISXQuZomxU1doaNiYCwZbdsJ
nAhhqZcU1tcGz/CDat8/M6PKhHGs8E8buqLGlUjkpX/pLt/b+t7M4T+WaOeb
OeFf5De4mTJQpsOLZHeKFpfNlLEcZl0jxmBCKQMHo+L6SAvoZuGEXumKUiYZ
iX8BYULjMva1Wkdzg+hspZLBDtejD1IoARjYiwSuMxLLHsXRN8V6w8dewoIr
8yXK++/De8fkJLfaoaifb98jLMQhfJtTSf37fpfeiUWxPeCdCVNDgVQBleJ1
OIdIfWvCx5QQqJwznnD3O/9IVWp9fpHndvFarvX1ons8XlkljY4DO9SlHdu1
P3covpiV3fKC9Oj6itwhAPy2+RjaZHGBwGPsjDgvYWtUGcl9eluCSAl4IKzb
OqDj4dv9f53CGdRGr6Y6pDwwFVf1uACVezxeX3E0x4qCWwiUQyikiVMsrBW0
0fillPgDBSgxoWWuGA07HVLqq9ZRzVHskCv7kupBkT2raD/DyuD86Ynho6rf
x8Yw8D0793Dq9kp6JOBH2fNiaYcwbTX0LrvAKg7WqzkUn5huHhGrYRZTyFww
ebJ/3kpBrmweIHknJr+uS16ivEl5dA8wFJWAv48U5lr9+faPlGtluP0/o9f+
CP9Z0kciA8hiYReZlecf4fFZUcigjZU0+uvHSTtmo99f72qPTYLPygoPq681
eXkTzJDrGcN7CDzJyZKXWd+woAmrWL/Hu9e6V/61UI6KnehIEUJbAHlCM9e9
xIsSmnt5knbOoAePWpKhMB0PfGO6Np4aLr1i8TaigWiAqZ0YrypfEctukQhM
aPPV3b+BebFVRzDE3xiVG+CI+Ag9/Ob5nBi6dZTnaaCqY+sH79fEJm3mDP7H
Xs3pKqCibtkd4VSzQwdkK+TW1ytIjLKZqwfEpUUoABPHMf5JhyLlvVOdVOyc
P1hepdYRpzFUkSETwCZ+MhsTW1yc0dohhWIvjyYBtGyrubToxLuz9jpow2sX
g8UyDmIm271B4+gjkumMVc46eO2K8qxdb8GlJHAcwZvCBz3eP+7somvgCISS
PWgv0rs5djiZzM0y7VRU6a/SOqoo9pWssWikXrVxKIhhpKolS4FvAPRX2znA
gdig9VFuSt4jHCvnRE/gEf7iaVLm6Pc5dJBS/vgRJFZnAs+x9cA2cWacwCxl
/V9jYoTpISSzLtAwQsNg1YHSgSEQ6c+ivfjh3Eto3i+SUcPi9IMG5vXIswiV
0qr9NEhfMIWUBCGuPiMAH3rJeMKLs9SaX0KrwG71fDVSGsgCR8nIONKsgjbr
mbr7MSPF+zqhYu2dGGPb3rf7e50W4xvvg8RGjpsmdd50yRm7roXTraoaPNEC
Xv1WwTOKRE+DHDiHJC+ss2WF5RBp+KH7TqcPn0syGJVKYj2zrFlP8/UBuAq4
rZJiRJyVl8DBSTOHRmRpSgHpdgP6obTk1dl6KU8fdYwkueCErDns0C6EH21T
bmzswyXZ8Bvub3LBKRHW5a+hjesmTlg6gFMNR02Er4XIoYL82DrpIbuMI7VK
Pva10JYDZXzMJbGy/gz3+KBdFXYavguK4WWlYbHK/FnVEMOlXFeju52KAxHv
1lCGU1hHwTfSGIJnZqOqMnZdb9JHSv94dx8lqWwd0nT3TillF1s1+SVk5sBo
jdpZ1X6Ovdj9OF+ebiMtA68PlCBIkzkOTrqHapsm5ifgS+dR028uDrAgN4Pw
ymiofrI/IYVhSJMF3aHBt0exyyWmqxFv/M4j1+jRm2EoQ+4XewNixLXZasQq
970NE4pzb9ca/1OvENTgJWmH68QVDf9B8Vq+oqczyDfCFu8jPFBUvvoEknaG
ItZ1tFXgvUIh297xpZ58TMQ/AK8jj6QMg4MBMEFdyc4MXAKntFa3TlsSRy36
iOXGeul0fbDK6bhbwfQx3H8TJq7jQjRouFtIiyTyPtfDt/ws261O7KUT6Hpp
8h1v58m+sM9DQnKSkLEYps4imjD/U8kzfjjBVC0Ltw5AjeT6AlfITooXNfpt
raOi5GApJFpGN/R3MZBqCar59bt6mHvg1dWZvRJW1DtVdbgbq+kIdV7LDJf/
u1RqvKjHH5XEF1Bj45Y+rH32aVd98TvgT88344DsbKRrJIPFIhEitOCxlgoZ
5sowMw5pRdYAf8uclsDnEf79aE9ylMMbBBD+CMhOuA9hQSRSY1VlN3xTPrE0
PIxignqDlGJKMplaDXec8PMeEM+RkBaDcbOqg9LZH926XS7Bs0SObvNAxKLB
tlmj6AApKU/M44AF9NWZ2EODTuJk3SE2SJqT6+3/lQqV/OL72UaHb3kl3T7f
D66r33TkmDbo5IFCb8j5dtCZl03URtP+mRr3r/kW3Bxvelirhq3chOgMuUs4
OmfRPS+MONIk0Y3A7AeLE+/tvlX59vEjhyDmA1/JxNxzq5sVyZ8RMNyrTl1g
YKc6AnRLcsCjxt2BdkgbIp9rqNR+DVvAO0DCdi+welyEOkrFrNWd1MVTyFxD
6obXBjqDIeFz1npoESaJbPJKnWPFv7OMdrrZWRtX5UHQFjgHkNxY4Skx67Gd
DoVAggJqhDk1zbcbdP0FjnlsT4cW3tI3qdXA5obcCeYmVbN/sC86S8LyxRT3
xt2PDgfegm4l42nG2XRwErRuFEsl79zBKU7BZMZl8Wb1VQ11JIhcGsF/v2LG
MRx7Zlx391lX3Lp7PchENg187zQ+h2hjag7MV53lGfCaUiiI9Aqj0okEwWa3
krKe2yvq1vOp/2b+KIj3ZsY43dChq3DtjK12GDsZ3hs51XCBCTma6cK5Q4Va
LkjN/VkSZ2Yu0pNpekozZ4OJIKAfc1ZLtOm0zy5/F2InmH86de+LicOA6NSm
z9DqmTC5n92W5skhSOoCjigMgqulEDktaGe6qEWay4KexBL/XgChWx6XXwLB
P6VccAKIuoOA3ryWpypQOoJVvv6aiHBvovICWe5ghfc52e2NcwzJvu5YLW4l
1HETw3xs/5Mif+xSJ2BJseCkTEwdc+XjBxpfrg/f8+yhWGakY9IvgdXbUzFS
7mRYxz6lWn3pO7rXLxvpWCV+kUX70D70H42ItiEFf6vjjtSDVRYbdXrCNiMx
4urkEuOb0ZQuOo8sE54XMeoAK+BVV0s3KhQ7jgs95WODTZ03tIwKb3h9iKo7
wig9Z5mtI690ofV9WQJ7KFkQqmL7+Yc9JtoLaVULJNUCP6+tSHtKgnu12AKS
mGY0CrklevFvN3vd+Z6cxCgYer3kHDjqqq31HIrVsza3qR1yjenOPFMPaJPm
M3pTrhktWHu+wKyb6YzXjc2KvxEo/0R2mDVcnCPmg4mBSt0xtrdDu8L7QwYO
WJt09zNatVaNDHQKSJZPB4/VvwtYBvgo+ox6Vou02BtMQWA4zLyFPXprz3t0
2lohqtJJR8kdE7+7f9eeW/6T6LJCR5OomF6qNGY9sLwKjnor1GtlElMvWR6t
8KnlC5AIYW7iiANoAthgLksHzxriSp070z20nEGhNeMAGRGQWL8ImEAeoKcH
QHQMvF2q6Uezzd39TpyaJom/RnnEgBzeVkoVLJo3cnEZ1MAe2ycN0P2bLl20
KTHnmaIxgm5Jek6kNF8qxTU0XwH017CjXSdVyoNalBhuaKD//+UzDXPyBWx2
uQQ7j8W5YOKp4Ol8OVBmsNfVzzqIdaOn4IhOB+3h62B1H7nLKKqYR77XDTu1
gd6Qjap7UoHy1BjV3Wdz1laXMUMkqbZTpdHCvu1s5kDGjN13LXHxpdv9hPES
ecBgcMkdY7lDcBHZqe80nFPW0coMtgWJc2ZusXzwgs3di+IGvsMJ6Qsd0mDN
+djv4y47Gfmy/eLBIi25nj12p3eTJlHjxAcT7aFgp95dMeZpR4YyJxVrbtBC
v5TJoibgAgjm3EAux6KwxWrW4Ztk0L22mcXI7BBdCJpvxyfjta2/1CDCJN0T
p7Ggtq8+tvtMphT0TEo+i725suj4ZxqlOVZD31O3Ho1UmvylllFJhGnMon/z
tHHewyXl7yzKZAv9pRf++d8I6ycMI8sg8V5yOn2rzmdYF5f29I+vjWrnxWYY
sS/ey0pOuVoUHKaZfL/xMOGLyDvlRNmq/EgktrFc7XV9xkdHJUU9D6hhXp5A
wv7iF7jd94RFbyz4A8cEVKVQIzOLSv99e/+VHzCMv6kT0up8SIXrRC65uFzl
hLIzGc/grTJzDiT9Q2j1ONKwxQDFySBXq3R9DsebtilHBer0jQUaRxrAXE13
qzkqG2KIg5GtWGQQtdBQYRNOpBWC3ULpe4CiARi9zIOSt2GRLsFgoibCX4sN
gZlqEDeOhDBiD8yD30NOxee2xenSUlAjFYIO+ukmTb/93KZ9cTgqzl2G0NfE
mNvrKD5wptjWHstPlQimgetELxhx4UI7w5DLjzl0pVaFFzgqOaMDZFf8a9YX
LCJeimFm8U4b05kSTPAGRPfeeGpdJN265qgu0PBC6FLW9mVloeHPO3u4oVOI
EjiaieB79pkg66MHefozzYcrrswqvT+wjH98UZzQz/GmiCV7gmStR8BNSUqu
7jCXMnFMiQOG3UWxDrNgXVjHWp2Ra3s9CR5gKgRIZjyTsQIbgWiYc/sRNlHK
2SJHN5thHuBwOxXNg4nyvOvgGUYC+rmU9w3MuPZUV3yInZe8thy3Q+u83Lhb
GjTzvmZmreG7dcgWMU6W3TR0ywmYR8fDvmS7xV1C88pa/UzROWjPQF2lFD33
+e1wee+Zm1xDXAjW7hxyKjvcTM8F33an2ij3w3to7rjVeZ0i2DAwfP/mivHN
073jx60avok1kyanhGDBUoQoZ8YOBI1JyCVXlk2Cs27k1yxYdVe9mYrcxaBB
5e1HpNpyKs2goTY8TlBXvgxXr9w2617AjukZFgjXH+vo2PW2h19kUMyJc72C
JuFGIO7N/CS0c9IzaFaLQtJppj7iumPq88mr5KepYP8sPdHHeKd4a91w4Tc2
fWULHRQcsKtggl5tawze5G0OlklLPDWwmuX0fMuab15M9bENybXehc5UIqXF
6oPp8Kgm1ChkR3t9jvyhR/5XRb4KtLP7Wo54zqaAbGwRsnfWC5pKcoS9XvYz
F/IGR2x/4ea9jLm36RMqSQV6BpOyTIuzqjWpdDaCOgvtSKDwC1OS8SN4U348
E6uBRHp/4L50rqfB76sLpbr8ZIdlSvw1D+WsZAD4IcoKNBk9OD7yqheRmHJi
4X8eo5Dl14VH3sMrBoprPCE7qWt1FxoouDPB/p0sQiQK573kOUxqRpzzTXpd
4DGPKR4oqyQEHtWhiR95+azvW0IHVLpVgxWjfE8gnahX7dV69KDpjL5Vgoes
zqfjGfWgasf16lj77CngCfZh38AqCUOU6CNcq95ZztXFHTlIqDum5aZ7/T8m
trQ02sBPJzdkKZHnQU/jnZL9qBDelMgL4v3lB4kEJ957UzEyO++d9X01hSeL
O2+egRMWJsJrMnWQAFQjD6yEgRelSbbC/Y7Iuh1SeCl8L4k2elSuQ/AEeCXe
O9j36WEO+IBFr2QOSn/Fz9KtzpIzq0b0lHUfMeAXhb/hPpYntwl5AeLQF4sJ
SBATbasOakiMPDqDam/vz6WeLlP1q5UNlerQRfXq70XRtkUNL+V8bjgk31Ep
rKeBLrNNKECQ5ZRfS/kpM4i8JdxE3ckErBGrp9ypT/ZI6zuQICdxDEEKYgb/
fN1ZPexn/4bSjkIPMXVSmfR64tEUSFIZkHW8VvBq/5mnQ/vR0ntb7akNxNNM
k4zERYkbpQhi2m2fag2Sobd65gZ9uWA8bkvLqBxMFz/MkmkZMIrfkzmxFaxi
cvKSF1Jk4U+8G+nFFFm+gD0kcrH75k+1LpDhN1EXxYpvOCEPhjkTd5bUWcJk
gK3vOyjNltmXe3xPGGlWzArhTFfxYUStMDvxbb8obQ0ER78LBnPMYoSCvRQA
j05TMVjwbgwFZbSWzRs/gaoFN5Aq5fC3XjJcbJXUD/LW3VAFQjA2k7pUONdw
wJ7PU4kMbDzxwUgArq//Dm0d9Dc0xzfQOWvncEl7oFiuEGsmxSAXA7taX98x
OQTo3XNa+g1uCBoRTZ11HWn2fnn2QquKhfwpSMn3PHlGOG5S9kSEvt11ih5U
bPOG5q45RqybQCK0NWf9xOWGjd/QJR2HmNl+uUOwQOnbAZ0tmqPSw/WdyNE2
wgA1tBdBfQDVtG/VFyrZVfHVFI6Oz862Cd5JlZ2NgmpXSENAmTI55g9pPG7D
e3Yf1gNJlYsf8hBehNHayV2lCqtKkbEwRO14jHHVvH0E5vag4XnO1rKqi4Da
CVMaXRiGREcGaewnGTSWDOkscFzS2WDNxRg9wwRdArFbDLSUYV+LPQKKHkbU
FGfEqIlN0r4kYWU+up6GvoL7CaN4B7VcVCdeK9OsxfS4sxL0iAqAix6RPDF4
cwqLTP54hFD4sPqQ5YcNkC/ap1NAt1gvoW0ucHiLtxJ1XETSv/RlO0yitU59
Gx8SR003YsBXLIqlDiQVmJ+oif4KXUrm9zyhtwLYarL42wY8TUutU2XIiVRQ
UpzROmy/t4xcPZKN313JexmGL8nUwSXgtpEc7bjAZFbNBpVoD0R6OumfdyV/
sI9lJG+gHBLUvxHcal0/bVzeqr5yUwfA1ElCTAd8qO8DZwgZ0Lwmw2WMvdGW
G4mlJmZ6VUG4E4bprE/VBc2+aBqw63TUwJg8qVwl9Pp9QcvR3NZMhowBHuxc
yW4bjPRKN5iEzzX7dgv1oicsdfwTBRDeUynmqgo9slH9JCxRkTL+/EhNFsB1
fChSge6K/JuDnIm9HueYzQoqBXDj45bFTObcRo9WXWvS+BShf+Xw30/6/cq1
RYpc2hJmBKU31UyTgLpodCwfiI92UtajK2DCBW3g9TcVx+phj7a3AMkaFh7D
hpIqJcjAtsMO/CqcnQFSSnLpKmQB8r8aF770uqSGn3WVzfZtWYydrAHXJ2Jd
sjfIANqDnfSzYsVJgymuIP3S5p33Y2+36huVZinaB1m/mBQr9X3wUWXkOPXb
t2nl5KuDyDI8asfFN2inuj+9OpW28jjjQjBClqn1YXtOp2Bsj39BxvYAso8a
IJyWSzP3+h0Hu2dMk2zmLvXypsP83fDf9hwJ/o1ucEaejc3vyGmQrW8lTAzD
gNLwXN8r3fDaUYpwlwectLXHf4qxQ2bVntuKLKuaRQpBW4wTZEthAAmY6sUA
Eslr8nwqPrbheIJJN7gdFINv+1hp77ffUR3g/L9CAnFp71TAekEt6gtzwSe0
MNzirqucVeh9tcqSMkfSzRRnAqcrPOoZxJlNK7qe8QX3eyxygsr/STrSwdz2
MZbLq9v15GJM1o9idlOVHqqBC96Xr4mjng5m7+1xliEIaXNyJsEh5JLMV7Jk
y6WGpyuz9Xy4Mdg53qwu5R1BOB3Y/iYR/ZoDCOQjtGLuzhd6x45gb0cpNaOc
WXmvXTLEZGgXTy+F2KL1uVLOn6a9Sb/NVyGq2prRPhYC3P0w4NzclX00l1Ap
bqAoTCIO0Tf3mQmz3fhNNTspEa8Hj/FWd9hDfp2BpCcCbG3dmM98DIgfGz2D
W8Qlj8++vsk2qwJfgT+OqUDw62jXkAxr1at0nSvaR21g5Wn9tjE2Pi3D5KHZ
NunyGphRvxQS8uw3O4J/0iGpGWNyQmPW9fRUKIExdOhpvTV13BNPpnbDnUS2
ZDCJHZEbzlMUoveETsTNtECNdJSaI6nfEYSQlayffy7LnD5UsKjiBnGWw5rn
gXm5DCzg2qt9lPBLe5I/Zw+fEivIMRWuxMX7Q3Lt0sIJsO5lfMWN48NNXL28
K/GGomKC3xLV0BITydQULFLwRw2eSvM0TcN9OljYQjljzlDjGbFVovviuMdl
OKlILHd78iX4PdFmnvdhpDFUujiI+1niRpPtXBDM2wp7Fltz3gsTr8ArXw68
y9TtAIcybomQtEUW478q8W8kxaZA3SQJaWQ+3GxXg+FnqkmAHGGqbtwPWKg9
BL8I0k4CCHBHwbKm9ObS3P8yB76ftEeoDu9+W49+k1nwqlHjgV/UrwV1d4ge
OvjEB6V5NsloYzavquBPuONqPjrQnEz3STR8BUMXNvEwhHssxQU9rAwQmkhx
qTScRVR5ZAtxIP5neH/Qados9NcgEFD4xwHdDFcVVDsQLWrDACIlg88P5yi3
EB8SxDxmJSNVYASQeBxrOOCkdzf3/yH636ZJWQZap3638PfKvKrS5RZ5egNv
VR6l021GB27gPZ8UOQyqoRVVjrGsUC0ujA+HJVeR5fzJJfZ9XPnyxhfSM0PV
sAQYSWeR4oykgn6A/zVdi1ZiS10NOZnOhOkFZ+wENNT7qpYU+ZaEqCtxZLwD
PUNcytiNCtAuX/hSLjNCkyStHi9LTVupl+5P/mNhSnOVU3AtXKvRJpIvOOfi
7s16nwTr1WLyJgkzJiqWUPwPlugwZPm29jTuCPB7Vc5sWQeJlBX0E3wAGL2D
jCX7d8ggZqtuTIjHldJpbpWIB5nK8INOY8R5UOOvKuA5PzZWA3tpJW4A8bKa
M+NLhkhx3gfdAdbcnTq5n39mK7jZhL5BPKu1pcXqm0p5+z317YsO5XzjvTDY
XcBxoS4sqjZTNq1lb/mknHscwkoZFic5SVRZh0I3Ndd/P26QrL16siID4OMG
2n8fS8pPTWYdV+YuOKIGM+iAuBjMgkWXUmDyY5BGd8Tdgy2dWJqFK5szjz9A
pmk6v8hXcO/8PXUoZCuGIGX02DD7sUfLGhF4n0jcS0eU4wPeqJx6kVsxEfH9
59+ghMcKYmWeQUbuOCI/GowxhO2bvoM9dNLtDDwZSzue9zqyktcPiFBzmZO4
2Re3fqV94jnqpZSfwHP/i6WNRixs4ecNg0Bj7MppI8V/QwEs3Qtn4EJfHBSQ
mO44GdnVqeBvPWL241XRjBJIISgrujqgeRqmuaNuWOSQ0o1twAEUnjfiT684
7Yk2BB/FdGiezqPExXBWSpZuipcj8XrI9hlE5XTJRmukI0kbY9A8ku4u0g0M
qdelbqHGzWz7fZk+QEtJ4vWsAGvyLO0HStKeWgfBkv+oBYklsavt8qjt8gN2
h8jeSNfw1o6ADy8tEPE0qxw2RV9hyYXPtxBDA1IC+bQSdxkp/Gekg/zFFDlZ
XtrBqPXQTH6SRs+KECifB3lDRqrXSXny2KRWG/pRHgxmMIxWH1hK++a/TGyO
cHuC1ElPQpscruH0la1btQde40G3YA/hEXXesd/CwX1UWCAluccFOVMHU6e8
4a+uvO3krj8zZZhj7J92iulWn/++h/fIJOSfJgcK253ZrmVkPqElTLhKry6G
RgXpdV/FQk9BV3xszoJAk4/kJxgH7vytHewMoAjrnobQZGbTvSXjsKOUWBiA
Pu6XPv3kTJQ7/1qrJCjRl9W9zXPSYgeX7nHkkyFoEcqYh79Px/EQRGw1nlAx
rBLbVY5g3oWquqsbi7vybjF1l4QjKExPnnD8hxjZgPRyXt+f6kJXAhFcai4G
kjOHw4qWJqwAPhYd3j1lFRPF/vE+AHdJhIkJFbRftCyoKYC0hZBPZrV+/+Dh
xnlJBnb6/KdkwKcEOR8FHyPlcC3Rsl6eOQ54QdTG3YnXAZSqVs3wXbH9zbcF
Jwi3u09TLH+XOn3tyxHEWfrF02arTbxaa/NIxpq9gfOygF+PLc2mtfB0vc/s
/pHNfN52Ge9vb3yq4tFnvLBGqFrrn0jzTKde7pIOPaq9QgTkP1Bqv0oU+QBU
I5a33wqf+1YVa0YQtZXzVIwSLJMXL5c1Orwyqfo9UxuBcJeTG8wxZywuUFh5
VKA3vSKIWymHCtxDlyR1d/XzXVTVF8dyYGs7RDu4DjGoxR+//pmdVrdeP6uF
M4UDQmEtBQOXblkMWn6LPpHLrDdaZhRqbUifCpnoaRM8lgeWyd83gbOVnw8B
ozAP+FLHeOD36W0nNclUt09OFlXNh1lCta55GaAa6U1ltVHQkF0V1dy7X9HU
i7zUoaXtDXREAw8q3ybUuJtpM5wI2Ap/FZW7zzNecrZvLx+LLKtG9EYHhcDP
JnHiGY5h/sOfJP8esD+tITMIvnrT5V3IGvESfi+C78vzVd1rOCtQQ5uvw6SO
hUuuCUvXqxb1bFfBgVZ7YxlXz7EuhErAvBQdY27lGm7c/BuqBy+D1fqBAN7u
4Lb/6JDe5RRy9YZkCdv6ZGEo+TfmTXf20ZM6F8LxaQfiogjpqv8UbKC/XUmc
HlCd66S1PBqOezlZ4LlTQG1/qjtH/9y///+k/pnjROp216eV4ZRfROpccmZy
Cpz+D416yQB5b7wJCHOFM5MsqikDQ5QO6/PFaQ4/9SOomBjL9IsABgZlKpXK
paGElBEDJkNcUNsiMTefgAKe7E4fC4xiACQ3yT/2HUAX6CBmRml2RNQvvDjS
ANHOtsBC+kZIbM1pslGWIZGdM4kGxTuTYzdPKMAFx/Jx/3nRippKfiE9+ob5
ITpYq/CsKTeLM5JXFLWtasxn1wm2EdtnFAtd86RntMQjPrCxEcayetp6+62Y
a1algKUpiHOYfoU8te9qiNBRidXMpXS9RW9xVLQIVvsIoE/MuTyLoHfHXxI3
mPFxDNWc1eRT7NjqZ6GtK3feNejA80yrYuf0vh2W8VXvc+KIJW/mPZlehEBK
iKth1VF7Ccw3ByodUvrpFqrwjvGj4pLuUqUaY9AhS9J6iZN3BZR/+Q+PzH6x
cILkWNgfTeRVvVxZ6mlbw6ONVddpRyZm4m2SI2EEbx95xOavNwwNRH6XwzD2
aX7R9UH+rbTbMqRFt0LyREzNDVc1nT8tWkOGf6VJUNeHDHIh22X/mE4ZvYjR
5cDOw1CDntX4wguAXwLFE7X/O4QrxxP5Tp0wbGrm3I69L1nO26PK6YtXftQW
jDU4wOFL/30TQIVmb+5CeWv4Jl4WRWLsUAdUigjYljaxh2GO8sg9kgDyDrYC
pA5vPcJEFMBERu0gWf3sLX5mij7xll2ywlAvzBIm4T6b2yPVjssStskzqE9r
o1k4Jwnk/KucwegvH2NH/7fcMwfE7DDBZigwAnfI4BJMUQR8N2Vo0Af1pQxn
xXvNAykErkAyPJ2VfNuQuoMzbnNEN4JcZej6hO8M+woHTpym79o0o6hrfjQE
ttU3vFvWSw+fugOfR7k2/JszlBmTqB5rFz69GHpjCgnjUgtyd04RFbcGfufV
VdaNMXZI6ocvRR3MhsHyxSNExW6mzw9cpTfPiWr9tPrtGkNiQ/cqMLLKF7Lx
jHuPMUqS6EN36ikAjDpVmjeJGeDoJHeLhT8lXsD3XwmostRdWHGbbG6Ajkub
jGrIljXLfNvkiZLJ4wkXOcz/MCR4mqPrlFLbHexNAbgBDJqX4977yrygZomv
bePeoUdLwntCuUQiosb2iCzWjmulf3gE8dZG0aMn8rV6dPSzd6Cb3wuQFMA8
vSVNNE/stI5bmRRorYjI3BuzbG09B+c9Oi73MAWKItgzd+ps5jcEU+6qFW21
4taVNcJdhpirv7vu++kqftlgKArXZ1VMlp1C4z9flljAmkObET5aE6ue1S7W
wskkUM79J3rZ+frLqXtXsMh1UV84No01PHfw7Lto6AQLIe+GWogpyh/drsZG
9/OWP5OrxcPEBKZwUDSvmlUVLwM3h/6ZF1JaLg/Ce/tFegGnqm/MhW2PRJsO
iN94tRXnQgR8nVa2HnUpssVtwAUnUVU+RnL+Wovo80if7+R+piOEdMvNM7c6
rvCmKItQooXStPGzHL0XJfVc4jDWiDyhRt24nM4yN7PiTBZe8Sc3xIBMqMca
oRc3oudmOPpo90mYMlVsDSn8+wNI3WdDt8T23ULg+jpLmeW5hKWy/KdlyemQ
iLxdLP9nUxwMGzeSeV343xxdnP++hVtKsI4Ljbuv+HQPBs9wRM41NEAmi+zh
+Y3M+LyeQt31Eiaw0BuALJJlkdIfXIcCcszBZM4sCFQNXoTw1EDvM+WnqoLj
WeRHFUCV9toDw0k8j1eGcogNbkv4kLJOPS1aNCZROHpYl+9AkgE/Kkns6/Lq
I6u/B+jYsYHH6HmEeIf3q3cMmG5207s2HkNpBwTTiPtwIHxjKQTjZENMQl8j
/bDEcoCZszTc63cJYZ1ZW5qUKtfiMOeAOA43rMARBSH1MdhuDoqsY2Vw1Ad5
Sdyi1zpVozvmDufABFV36+u0qTWla66W/N71z4J7TN5Te+z4oMnU6b6cRK3M
5p7lxrkrSPb1dTHbJCvcopjJvF3IdfRDYImG1OjIHrB/9233dypwlH/k0sUb
+C4twlQ/Ft6KwwxZBxZ/ygvy8d45AghxwtgNxxZeZqLCEfbyV8ztqg8y1NA0
upKwWMBlzJBUAH18BbNRByNopDZeG9AAYYLVWibrjJlvDiKTjyYPFLiEBoR+
neO1Wo8j9jYS2UFqb/OFy/oT/BKR6hOd+tq1wHCi8T9jj7eC33d55Nje9GGE
xfosXpccq+n78fv/isZHBpqVqvp1nEAa53Y/vMRHriihYrxiXio/EhinySfR
OwgcIeD3IZsb20Q3KYvskzplPccvrhlcsunvDHACrDDqMxQPal+FDOXoLbST
0fGVz//iiuE3HDQ7pUhwE5JfGwlYNK0gUcIdZOdQ6RdSEHMNAWkWq0RKbSJM
WQdqfJ8JVU9SGo9YhTsWyS1OR3fG3XcEoc5ClEM3+yidTqSQdjl1qHv6jBJo
qHp0qxAZE33FpNvPLfoeZ07FFRMKnd1rrwD7WCPVTojr/e3ERh8dcFr0HXha
4DsqKJubpYLvn4dfEUVlo3jNjXdWNVp7Tc+pPf5whAmwnuKrCPuClEbjkihS
6M4kA8KA+ht3no4OyN0vid2X726kC0wR6qbfN+SJax+fnVE8WHjZDfzqryph
HIJM7cKRXPWgPHj708rs/OQ+UXRmQP0SX7GJWW8DLp86AAUJMm41PcN4u9H5
w2yEVutq0xEGhTbHHoZegqj/F2qipfrqdAc8pm4Tlz5ucm5K3qgf9cM8FaRv
eERloprqG3FkXfiYi4+s5BxSzUj49nPURVoTQUneTth/+UMaL7U/ZOBshRxo
pCUdJ1AYiVkPQt2ZyUcaMeRWIcxgD95iLQ3ShJ0JUsDXA59U1CxJdJzKBknP
lrRWrgSKxYBk1mPgqJu46u0J/AbegKLmbVCFPpgrr6mVOMwmXLAAH5quindp
tc6ua/++ODzDgFIALsz3dd9VZCKAnXWkIZYR4cLAl021iFMr5aj7kWxZJ+ot
og/eUi43ObkEaZ9ao9z9S1taLfnuEdT8T5R8q1pldlUmi/2xb8hhTL52kWvj
iCVkC0o5u9JOeG37uMSEkp3palQeyttmq2JHvzVjKWNYwxgdZoOs/e+Wxu6J
ZXAxTlIV6+VIH0juGOY4HHTEhbpJVlTGXSWScuYbxfkY1qM3otL1l/o3I0Ea
WCxgbFl75yU8VvTcAxhRfLg9238Xbh+ngG5bn9dYgN4CVkTXfoiAqypSsmfI
dTz5Nef2k4ih23aRW9flsrY16WLL08uaUs4ksMI2lPqT6W8Pm6eERwBGCWES
ZklSytwiTWfK/Tkz8cvBM3o7RJ3QYqmJfoJTZXxxSeG566iYdAGtA2IwUQtu
rJxe9V5vzJJ+3mXEkHssPMr7MoyZDE6QCq/dJ9pZNF41Qeo9kaUpk2LC8wa+
/9zGjeYDENd3TN8TLEurkJ2XKWQnRFw2PaJlQ9OPDcGCZVq1zO5pDixRhKIV
6gR4LuGGQqBbK+dxwbcQ3mgeVtAeehElsjUx8fBa7sUmJvfSTzmQkM/8MrvL
uZN7ZfX8SA8kygmOI1+iytfBghfYm8HglSaPBp0yrh2ttcDLZ+H6KDi5wdsd
MFuh94JxJnIpRm9nWnv1RGb7I8oWHBHQrvqiS3eofTjxjDl/rU7Q0t5INLq9
SlQ0ahDms/ixG3fk6X9oO3foqvsk8bjnighnX/HZkr5JFRIdM2btF0zLVYQE
kPd4XHOym1m3qRBJUp4F/WZIteAKorIxO0z34WpArIi22S8jcCaLB3TlYcUa
7n1oLGjXEplI6OsBvtQpIsLiBBP7KiK8kOgHtSYrvond8iAnor+X+GpvWPbH
xxR0E7Mi9mOHo+GWxGqZZoxs0vhUwin+6TWvuXJ4VO2mjdhHmnk90HYw7J+T
ZLH8VOY0e59aRcd/dYpnjXvST0QLvL+qrGgzwbkG3D+oLgOMbxxkABz70b63
Ave5sFz/a9i59nc0zIg0iLmtn1sZqkOSn7IJrIGz4/wVFjkWy2s1XAWskBBw
R8iaE26tFa6rBABZNyh2vMqdhrgUYBIoK5MS9wii6+5iLvc0RwfqAwjtOwRw
qJdYfMhFAmO91QHhqwPcxC9J/OSkNUx/eBexXC0W7Ix0ELa/M78d/jh/UO+k
RBPVbOMUYoGfHhRLBYjiQQ3NYzTSyZFrhwWgQFTLHyMNQoxNFq1pjDfcgwCf
8O/DDld5tK+v2sBSSH+lo+Uyo8hwNLvfYOH5G5OlS+NhCNgsFXjDDGg1cc1a
2C4FqPVG0p1ej1vlKutqPmAeh41aAvW6AMAxKl/OOeyj8ED/gYA2we7K/U9S
x80hxngrR4A3wuNGhno48PK5plT10AXaLTxJoRPOZyxbPul/7xwvFQ5RHDFx
zBetZPIAB6wvAV4iwNW5/zw2sLkBl4+PO2enPXa3swDqUD7/pbxEjsW3tno2
ePROfQ1AeojtJlW7KLz87iA5iVUn973ul5Olr1yJtXNy0fVveC83iOLNIv20
WHBJL1JPIt7yvFxa7iLGo8TJ5/ayG2eSiMLNO+YRkw3UyPioyAy8yKUXn2Lp
hT+hvRhMwbAyA6eqfAXpiQNmA0tL+FumtGk6DAbWVXrG62zfARkaNQ37kMX5
MePLkKZmQ1P1AKaT6OACjHxf+kf3+dqUPFRFzabtRDu/w8TEZ5OLFSLk+j+0
NB8rqDW4AyNZ31gvWz9kDeLb3wsWL90v0amHkYXoTOxKhJkMMktE2P8RZcI9
L+N8DgWNX2vnnR9iDriF7muQoqlONDgGLUUBYDpdfc3W8Re33IDz31hRj188
SaZ2wfMRLRrxKxXWTGDJZHm6ytictdbdtDjudzz56S20+cTVaId0To6r7+j5
jHFOlzVPN+wMjzxPL4tdpUk3AKZbPd1Vp68jUUOyMS6uyPP77ofK22NPXVUW
jZzBtDXRCBQyLq/kWWuBL9JyTBniTwkp4EhKjO7Cp6zqjZTN7WFml6jMUpOY
ekYIRN6jCLUEtMV74M+TKnUxFqokSpAJNXBUC++sot96+fTZNB7ejj7Y2dHv
VF5ITgygTd6QK5eepcHpOsl/PzbBsJJUN5P5/5YiHEGupl2yipsMJwoc36/r
mqx2QqlY4EC71Fn/HDiHa2Avzdu5otH6zpHcXTV78sUdrGT41u8yewas6GgY
bq4to0I4CaTXwwnxITEm3trjD01dzt5ZvGzaYm3jepNjUmaZkBVWIX2qjOhZ
TXdDbv03uz8O50TsIBbiAg8K9ddZK/ShJH5gRvnZxW751gtLDFbbZiJwzAm4
KnKgfOnQ8eGSrnhP2nBXdZL4mpdoW6uFbpIa+DpeN9ZxVPnUUUhSYoJt8W1V
b3WIu4Ng38ohDepIEz7VLNCFG0db9rgpUIoSaSBxd7itSP1I1+2zkIJzhIbK
/oUUHpQbmEm0Li94Ah6qAJWWOIz0X4XhBfiQrHyoeX3jSEcM/sXYS/YhVu0V
BlbJcfdTHjYQ6rRSNyvOrsB2RC/4ZAfV1hbsgY4XxyczS9maNicLZiRDBKLF
ZML+w4Ue3pfKvcpDFUpM+92ycK94T9rUOclwW4XuYx1Bk6edluvqx7gVoiTJ
uCJweActjelL0pFxMhmguGwb8y2M018z7hVE6KwJwQwx51VsEZe2n3aDVqEv
FEcalgyYWSOGuT/JT04TnfcopYZqRhkKbFTtEYta3CQnN5j/Il7UV22zepDn
7N3PBctk+lyFLpLck0xwGODDwb7isviAnuFsiJjhTuM5vNTRm0n+L0iLAeUT
bBw+hZYTryRY8WrMXocbDcFzJO836a/EeF13XhCditHMxroZYXfLxVs6bDoD
uMd5zdYitvHiiElT0LbXBb7WpM8+kWuuTr3FsvgfdwyXxPDH5tEPQ8h/QvRU
e38RaB9ilhOvn0DKb/9ufszRX8Dw7ez8stx3of6zUI7a/P3rrezhsDtZTG9y
cI/KQc2bsV0WwKQiUlMdJ1rVCc6vWXj+I600SOfUbTiN/pKGqzCmsJaOXQ80
0o/5E/bBieDai/rLaLtQPIObgo8r6uRMTMRSH+Zkoa1vdS36t6koDkMjW/0R
D87SSO1qFVYna8dG6A85p5Zw+O28kDKg9N8G1QjXJF8Sl2rXwKXelzW1C7gN
HtlVuqrYQAYinXFWuRJaMoSxtg7NorgidTZg+FB3W2w8aMWclk29yZxFx6Dg
Mppx48O0pDdHZuYtjlUJdkleVK1wI3w4CV/ZihzH51njyql9gsVwFy3uZCbd
lJ+1UVGC0plYKL53sU8ZCMQg1jxdGtw0uOxa7Zl8tXPec//TUPsr67N8pUJj
EcJ3CgVo2XVH40bzuly4A5EtThMad3gzKUR6t0IHzgi5NkEML6Otb+ungu6v
w/zDdzcUIwmhIC+xBucBpe6kBgqp0Dj8hX0diQ4YleAaqwhRwfOFjVpC3fw8
v/g5IwjpWDy9JfTh9vihQD7MtPGC0GEZWJbgy7QW488qOjZ7BsY04tcEyaFG
G9Aw+9hUNH08c03cz/ntgQpyZ6p4FQBX2ii7W4e2+2DR+WnIk4Pwk5U2VCB1
Z2LNGCwCfaw+mtoK7FvPrNv3m9zdB/YTLs5CibqBc3fv4PyCO3fYu1xQrjZD
ApqnojiDCT5IRqL26zfbsJhEPjRB8bMd/cd6O+/VRsGsTN56bfz9GQOQI3Bm
NwIQANUc2Ied5aBbKd/9g5MRQCoP3sKJ2k2Y9KcKq4JYRy0YwsQuA6uO/29s
DHf4PoT7sXA2GQiHB1OUAo2DzfdpTl7rpnxvkj3qMy3ezbw44nXzNmMp2UfY
lJPgrKkUbSKWmqmmRWAHJg5CWKoPaPibkrNn6wm7FhuK0N+4whOdJix0HDfA
VBU7rJa3XMIQU1d6qno8IojFATHmecKI7GmT79ci5WKdNHNGAXBiwKwMPeXI
pzKJT6U9jJRySQWAIE7GEgmFvQXpLDppfmZjwAQH7Mz54rOmgBTcKRgDIwBf
ObRDC1cC/BESViEvhNuU1G9qTT0V2yar0xHkX70kNwXi+aSX+9WWjzDwnAcr
vPVa82QYfFkNoEFtVGpBlBfKgdaTov+CHCCY7+z9HlUkrBdAQA/dPMu5DEG8
f7cYmblHuwY5HidKDDUvcWD9OtgC8P9ddkdLQwlZzXH722BYyIn76qy0jd5x
f8c6lvTl5nBwcb8BzSUzfZiQv7ejAIOAvZbi+pgXdu9NZECKNmyJotmd2HLp
ffrqWLuIJ6iah9Xf/AAYNrh8LdXFHwGtaULLfiw8a2eQ4zD+uzrk9zywolTn
Bw25GwR0hAQoQSSMmb3lsAcr1bgsLkrv6ofSBURbcF6gA93zatp/V7IlgS4S
h0Pa68FpOr0Y1KH5U0xFQKNj3kfmkWSEfKScQtVtZTrs4Ql8sCfimCbU7PHa
wF26anC4302/WiY3s+6RBfUCREZxsK5SkZlgtd6BxBv+fwisZqP/Zhqu1myr
3Xhc7RA0lckSovf5Zw3fYe7q0RA8tPMAKg/H+FKHplF2ZkGOvRkOgBgeNYcZ
3aMopTaP+EQ2Omy50uMHBzn5eN5tw3bDpu9Kj3booWqKdZ3mSRg3H5Ms5jo+
oZz2VGUxLEiIX8CqcfOpKpP9QP1trPh2k+gFs3d0DIiJ42PaiasnpOA3jKnf
NQcKawEJYH5g/fpTWL4B0ovns2vbDI63RWfjjxiNWlqGd5O/oP7U2GnYKFbh
afZJiwvDO0/GhPPcSzhc0AK2i1nnBY3p8CSYeCf9BwHN/SReQ01foGGu0zlM
MDopxPWYlEiI2eEm95Y/RhNFSy8VL96sOkTrSZt9/vIdhEZE0W5sB1Im2sPt
BX4F5BJq/ol9QItU8PCc9GtYcs+N/GgkqIGpYhGbcLyM5jIXbNmlJRmRCO7G
vke783tNDPh2/mWTl2QlZ7/D3eZzM62aCEH6HFHK4vFWAx22qTH8tfPG10Wy
rmblgTDs3YMEyUZR6uhxEsPilmaHr982kr8Aw2CJZN1GRectRARH9yIKeg+2
XYlAIj3vQnK+pfJcDoUQAWDB3/OZD4CjTnC9iB/QP3Tm/fkcJt7/w1XKTnab
DaadQJniM9wgNfuXn6efFmlSHgaNx/cCeeCMwAJetuG5bCx3JFo3RVsv1JV5
oMDuL5WA9Segn4asCJIKVhwqSSE/iTmF+lXSnGgJhi1Iw8+lWGja2+TBxN7I
lJEZJGXL5Y2mHZcm9HN1JQS2jlWx7Zty3H0sYaMMsQlUXrW549xGIcnpvIat
aRX0whd9C0XdvMXleGkngqGQ1g9FbVslva3SygQIDQCxZqOQYbaJ1Ie9WuOH
6BWIdw5yC45LN8v7cKXX+NzfyoubL/w/msnPWR3i0VVm8hlR1Lqa3HMrzbjZ
J3XYokyneAUL/+lHz65YUGnDffEDlBp6nzEtL+OijvpXdvbK/voe0WbjCmqw
tv/sEu1Lj1BF53z1RYXzxSxKvpmEk/QrS1VjVX0TUDDI8fmV2tvevYGCoxPh
AOviyTxGO9+LmELhanYyl5NLC2xuafi4aUhvCpIQGVYz8yvs/NAHQNFzyBb8
fkXn07K+GYIimc0k2oLkG5VBiw2zK7p7FKsealWailtJLIuC9O7TU74A9gdq
NPsR3FqoDol1+eEuOoSumHCM3cCsGaUmzEKn3J6bgArbNo7xU73PCM+j0wku
ClAGmimhCJWZ7eY3Uedzw4pNsJ5lSkT3xYh5/53gWgSmmEvttDTRbDGx9sQ3
gAJrVFYZMXK568arY4DuWwd4ij9boc/Eh/gXs5rALMANwF7Auf5IJWrfBYMA
qAFpw1GUOwQAwl8lx5Os8RZoEvlI006XNt32qGIl8MQp77CIQBHthCg0miB4
3gaXDv1WVAFxWrDz5or0oxAusTU6R6t58+XQ1FpPMSLgn+wUSVf0TzlzeLQH
pmPb5Oos0De63bGeLnwfl9p2tjKcZttG35mC30FBySife0fLm3jeNICWBzP7
i7tJDyGXDKiHDIVPSCPrndTbuMo26DQzGO/T4hBaykkmuHvSCA7FPfAVjrdf
TUSwx2BSwTD5pOC6Ex4fo08D7IxzoSToHgIEk1Gaxquo7ItA8x5RC/cEVoyN
jMiJxly7X+L899QonhPKZzPmqwYD1GF4EdEho6J7fZaV9sMtO3NEFfEzmtGd
TY49kppJvN3z4Z/qRrtZFsms218jWdSfxAGb3VOQDrqYc2PmpV89fzyWlGrk
DdsgF7hz4z+rmhn7inHuOeL9Pk9yVAHeHiczpMQqdlH102AT0tQqnanTAGRF
cjbntALP3ksgPV2oLHzuAbPEcBX2zlQf7i/jVHk2djh9AM7AorcQoKNIQOAS
TVvnjAVNvH099UUf0ftcT2Szhvraw3b/0AjfoDMRh6cgs0R3jAllqiUSl3R6
2zRvHShfiIFH0j0Xcz3brPVXIpo0m/mIXKcMbmvYib8hfCfLv1BiAD4gZXjp
q7qTmEeev+6CfGBqacs5vS1AirCt4upN7dG571Kd/11ILoIEJDZ0rIi4soVp
mUsj5dNM36gQY0Tg+nLJdYkKuOzR0OlkTnl5qYybCae3zWY8pjxoByQaJ5sA
fLmDHqS8l1sAAzFEKx7gpnX8jyXZxgxPWRFbjPAtoyLBAZXBp1bKY9wvbMMI
m09U4Y+coSkeOFK3zNpr/50rPCThn6HsBjGwUzdefuH5f/z7tTZv5YA9m0AI
Fqwr+hYvWhWkNvAO1QKwHnvYfUa5w1o00vcwB3W7fsIPkOF0Xg3AVDZ+xE9g
UWwdhIiRERjR+mGmtTfDMYNffE4dr48XaPqWFsZT9MYD0aBEiw74D+W1EJnA
W8d22jbjoaWkvnoliuK5GMfgyZHi6G3NUCIpAtt9hDTukzCOI0AAAtA6xwms
RFyphW6rypP9Fl4mcQsHfY90dI9XrvwWEfdDfbdeffqS7oAruafQTEndrgwY
IKXCYHiKLAhfR+LuTHtDnU43nDZNJePsX0G66DjHwcefe2GDIQ5aKvbeHpP3
xERH4s28oa3tX6FaXkoeKK3rnI9/kXuVDfIf8iJ9ujgDGTOHi8g+Vdy/1x3i
s7bMsTuOLn2wKjghuQYjGR5fplkgiTYd5NCvnT93FSdrVIdt8w/Gkbc9HyAs
/QO1yE0kZCjOAoOnCgDpghX7kD1UoCqEsYeAXC1uUmvliD9VuRc651jbL8/+
QUGF7FoOzH/dKr7KqtOM81bbKlOULmj+qBTqYBqOtRBgL0YfkIPw5shvudjt
9WTmr36BBPRgI8Ik7X1fexAQ+0+gDtQULKCIl85Hom8ElP0jKmHVJgf4dOtI
QO09oNzMBfBHFsUmDPvxOCQrGepdiuDvV2U+JXefFgD71d8N21fWpNJY2lWq
Y5yuavBkQ8HiqmR0Or5NUWhZWUqZ6sCSB5Odgg+u3uscORlWAhiOK+Qy1qqu
qFvIcCwUGg+6Ouh6YifFwMWPvTewrcejBiUk7rUiFzhEhpJr+bmxUhn/b9k5
PQEqgb97fR6URzblfLagNFhLjE+NzfH0RFSCuVOjdF2xz+D/xfZ6PKAH1v35
LbgTJfT6+t5Mbj1UWyVQGV6HMGD7VTl92iv+FlyM2NJCJS0d/36+zSl/fM+o
8qhBb08bOXh1Tax+DKXCVcEp8FxeFLC2VmKX5iBeKAVrsR6w1YHcgivJoQiT
BhW1ER0hxeQenCLFGhY8VtRXSACCln96QCebwE92Wjjn2TreIA3tKZo/FGiN
zQpoAEcVi+SXcg6TkhefQsHU4c7ClyebZdK4BhahO7JhXg0Njq8J9/GEDJGi
vV9l6nBsYUGzsaeEIhJgc0M7ZbUgm3SkNZnwe6fNmrv8Z0QXPO1nlqrz3wwY
aDAsNPquYMJcn4QrjT4qjuHof2NWRGde7gOIEyJmAhAXvrQy/0r0K6aXFfVj
F/eAF3rPVD9yy5R32rp0GEdq5WPKxocL+MNYZGzw2SxgftVtwt0VHytYPNKz
pojs0jFmrhW0dT4gc36xlpVzZ8zMpzwwMmGvch4yOE8JVTSGP+1j6mEdeM+E
UHKgf6bnGIsaC90xuGHXYyQMHnnTN4AZRYti3qZsB6LT441+O3tEsYnKdoqj
MXgzBcdtPGoremjx3VAgwzMQNmABye7IIiww4UPmKZccPmox4D1yEzUdZxEj
qoDFCLlv3qzhbHMGQa64OB2ogp5w+A7XC38Aaov5bSJjRDNQqFSfvYHyLMLc
VT4LLeizqKTKrE7W5p7QIacZLJo8AcwH4UZ9xlSUi4USKLvBpA+zOFIpwhAb
fD5qr0f1fW81Jp143JmjtxdUvI1VdqzRqMKnGscTe7R7fNEcLblObLANGju8
6qA+Zkgm5ZCEcyhZv4lKFRELa3zPsFCXBJk8fqZQ7RZVwGVw9eK/VsDBhunB
gUwhobEPAzpsW5zpF7qS6sPNcB1DQPSx/C5SrvIIubQmno/RgSw4OwQQsHlQ
8JcHB8UhhnvAwNCmI1wr3YkdklxhYgwfoHRcpN5l4B9+97SMlNs2rYSZM2Ch
ZjqYAt9USuball/lGXL3QEPtVSsRgLoOGe+aQSkY1bFnkJ77I07MgRWagOSV
pGarSMH36FVp7SjlTbuOCXK2/w+0zpMDo2Y+B/ArEWxv4OceFX3PVcOQrh70
Yck7Xp2hVsAU6tsw0ZkzNHXjjYU7gMjMD4/cSbAK4uMM9971pnj5bEfljW8I
EmePNQuERilTuCpOWUzmTiXaXKMGPdyttii0lyYLa6tYkv6CXVo4EoYVtbU6
kZqAyghZyE0o5JqBQ+cvLO3kpVYEDgS7IKbYxwvxQRtgX3Ghb4l39Hgnrium
EAHcxB57oWggiT1iy/pWInZ62e0Y9rCrx/g8G1KFkrD+WgCWKn/Ii7olJpiw
r0yWWcFPhDC9AxR2f5/gFQqpr+hWHPMx+G8eCASUcIC7NEZFjGqarWDfgHVe
6xQYeJPuAlEdq6su8zKMGJuCQVIy1R8x/9Due5vO68ipTIVWRFyuEd4ZlEha
BbkQLTiXs3FRokWq3i0zML2RSGCv1IbDB4C/Wau1TuSyvNRUIHgttLzPMKqg
EukapwXTbtZxXc/5FwP6ZpcFTDvr2CRnB1kSc4VAza8PUQF4jcqrEJcty479
jE8u4XfrUEet5JrJq9gUfhQiNJRGH7ETObgIfX237hWlCD0s7B/2k/RVjTmo
gr/V3VZ/aOtgSGH1uGKLjBYXfLfZEdw9UE3AcsWpHL2vXIeD/7pgKX6YSDqq
Kw1GhoR/FQpEao+s2H/K8u5Y9SsnzFKG/gP8/arruKT0P0h3d3Irt9a5CFuU
0j/1S3jfssYeAGpn7BjYfu/a65yKHOAAUjSxuZWDqiVV4eSsJC+55IZn4STB
3l7XwSzlIvfPmXk0ZR+4dInzIdSyUgbYa4kXQTCkSlT8GMVJhad+nJ19xG+q
ZLGM8RJX/xnHfuvRO1CrzBTt6g36/xBd+SKAk7qIGh9Ma1fI3a+xc0qVN5Nq
MztXuKCQWdNimxa6SAq0dN/YvMQVmTfEPzE7NbyGlob3iBepMYaNGps/X3XG
iUFyVECn442QT7u0J8nlBZ3cR3zgtqAASduRcwnVvu2fWYyqNvdqlBU9m2hP
gu1dbeFrt6RVzANLLrHsRy4s2LzgVCoQ0bRDWsIdoepbsd3QhsuLLJ9MV/jx
VbvRuFzZ78cPwfSazFxCmo+KsHfWqFpQ8vHd+Tu81h5/xz8cdFfsPliAvQ7U
JXGSbuupk84uWdjHX0Ikc1+8j8oYCiwvfzCUHFUnB2W8xwSYKN+HPMMas7gb
63HKIaONDbhn6LMfF0xk7YsJ1ycF//l64TqEnva1FjQdQ8ElqN63oIkPj1mD
tBqoo/ktn/7z4CgSzI/iRFY5ZQvvy4KOFArlEcM1eQD7A3OT+Kc/KeQfITPb
E1S2UrcoarQPwVovdXsFcKCi+sWhUQZPvYh/SgH6NteApSHliOOMZoGexMgM
vwdcQ6KC0dVflTmJl5YZV6bSICFYS5CXHBJsKVTwHD6m6HsxNnOKSUfM0iKY
zQx+gBEMBgcq5O8102Ni7RdBz0OwN4eILT7a5i0UZu+KBuov2lJ3LVLj7KC1
3L5el7jhZ0Eghdl2uxZa3MtqBJOp2VEMCF+p0vYe5jQY5CavDZTnzvKlHXGk
4MoKxW24hZB6IbLcQGEf/eky6EfnLg4eW3UkVMUrLpSosmuPA6nN+u+nRspP
546bH2z0XM26uQOHJLt7cWbeDik8ANbMTb+694mBYIkE+rfH/Qs1oF5J0xYz
lyT1b7hzcv9M6Nx+FJ7I6bBWBvCdsmFA6asKX1sUrBhoPRGjV5W0EGMIxTQN
dx4C7LeVh7TjzF/HA2gjYirCVfgD6prlqkE65Pu50wg1tHVyJ1q2XfrxiwUz
N7wJg5EJObmF6ISstpZP4GhgPNLNZ8bBXu8VlvaJl2sApvZMGPZE4UsCWlJO
IL3w2WRUX0eujAkbtq/oZHYUXDRd9cUugyRXvhrW1u+8vkAoXovl4cQZFCVC
EHs5Ry5+acqu9Frq4TjcxzFegie7gbR44Cxu+MDIdeDWCkvKi49CW3IJkm3i
nnVqFpdICsPRd7d0ynWfrR1SHX9MpRq9gZMGw/FGEP1pfXze59/7JR5nSAXN
0DCOJTGfoJhZgys4ixPACakM0OZKLbIZBz60MRNkViFriJztldbk5bcsmjM1
sl04YHyo1HJVZQUhAj3qtzvXsmVb/N0iyexVwOl11zCN+OEM9gvyJOOxdQxj
f0KpaKWiKER3d0o8lTujb+K2CnFLtwHfeP/BQqPLx1/tQ0oTD7aMrxsrPeL7
eluesL5OAxBAgFHGrWnfgyjmFhExSFBqLAAphsg5KASOi3a6//J16iTe9tV5
y7DZltcQhaf6QvL+A466ATC6KyB32XqiBDL+N0Ff0BSIZuhGB8WaDh0KG1i8
TfL1i1+Nt5njnZnNZulwJ/IoBSExdB5Mo9x1zVD0y9dgHZpL3PZlgZY0OgsY
nOEv19qJbqDTdt+yg7X4eOsP36d4Jf59VgMIoBrq6SnyhcvK+tcqD690S/fy
knUUJfCd++BG9DfJDLASRRum4Ld6QUu/i3/XubbTAhiIltV2nZeSAtvIp7MF
xBJXnCdxWvczrrTuCU0em7QvMa9okGkF3tBSekIuYHC6b2FVFTu1R+USzCQx
msjCpFzm5WYWA0AbIkyv4g/WEf/RvOvbdRFbvOkH+CznOen22lca5DiLC7K+
QFLJOnzuzu3XLR7lvFH9EGXxOSglPCZ0oq4H1sBeQFXwFhzysn2avOkcXa7H
v06EHs1OdIEUwbSHAjeiwr04gxQBNMvX/1O3xu4s90+thS01L9f7QbXnx7vY
bFOfhU0Ct9AXddP4GosPob46lWeS1tWF+v/nh0CruTK8QxdAE+4OC5u9/Cdm
QmaFHPL4oWIilJZ6FnixfDcI8i4Ylrf0r7ziMj2y1JBvaEOuj4qXMy9MniS7
NfOTlbEJEBDeBmSctClYM/8qlK7UGgva8eNzbNsi1ZlGmzqfmVH6jRQBle8m
hItKlW7FleHOo383Cq9jAIaG5/hESWiB3kOxwD+sAFG7ubhqdvznz/ppOA9y
QLEmYUmUP7OmnwAF9OBK3RR9nbK+HZJhJttwI8brrQZ3BHIa+0UUuza/6q5l
2ZCDyEaORhYCKojfSeTp2CKqZhgPd/cSN3wY8Qe4rQY/b33xvQEirwYX/CZR
IiUbqJlZli7Xa74KNpuNBkywlO6MeB6Bx5g+fhldNNfdp6fdo8MqXER9pSiZ
3Ig3QM7g3eMddYaWsIfmJptdVE+GBIJVpX1/9v5vod5TmJDnZpC0j6Cljn1Y
b303jjhBB2jZESLoHzATkJiajgEznSvDwNHLi9wcccRoKTK9UvbCffkrBB12
X2DShzkuBetoAwA68rSyKPbV9sCFf6H84HBDfurQt3BQEq4BlqeusDu8sR9Z
XwWWCmC/0ggUhqJ+8YHDIZko6yOfLFWbDptar4HLtjz4Wzcyj/7y8BE0FGy4
xm816WKyB4ZVo2jj9881my/Vd0jH5gyrhywJ3p8Ph6t7odhjKe+6YbsX0bsI
baOjkG6IXLYn4n923WY8F4sAE9eGCvhaa7EbxALSSGBT1NEblixARfwDQZzM
FHftBCwJY4JORJ65w26pbV++m1kqHXIqclo/1clEdXi0BukAqf27VrcMpiz1
tDv4z5+PC1YI3WxGabmf1Vpn58dsZC4A2zBqUwBsw7xtn3wd9CA8k3w2zqrE
ai6GMhBD5DatihrNLcvLtHhqewCm7K4PY6O2Q/4DiBPkFEKxUTo1KPaEjr1S
ChPlghX4t0WuXX5DaV7bn1tGdJFtGK61MNP/3DFvkphSmZ1YciyPv5Y6oo5Z
dPGCwiYzf0A/kIrM7AE9EY4WTe3F2y4LqWP1eTqKHU7MTVLSZqA7egomZQ0+
b53pmVGooPTO+RR7FFBMNuABcjkCGPhGd+N5ELeiifCgeuowHm1+3kNLeRXr
mAIo6GFnD9s88jRjiLSl+PH/LDXGafmXgIdLnAOlBXMJSX5gw/xJHrUZ4cgj
CoyMMb5+0yIUJrE6OY5wt9+y7rM0FCIfuV89Phq0o/JFoW5rBhdF9nc3kVw4
hY7J/PeWW4nKZlte59cmbjyxqAcdPayYpKZhfL48StQ+1pv68i3nP7OQ8MbJ
O9YWcU4vZa7hkjDSBoGcR0EnRrkePAHsluAURwQCqpvOAnM2CX3aPjqBwStA
MtSEopvtXFAQW/mfhZYwoKaTHLKCEqLuWgn5Zn2zSurQ+JLavrqMC2hjIoms
y2lCOBmLMD8mZgtkulLN54MaKtBJozF52Y5wUj/aEmCOPu7aTudp7yIUVl5u
8bC2ziPrqOCe11cUNeU0h+rxEQFNwV4jkVUJJtuuJJiEahfrw8Gwg8jPnY8q
9R0ITIz/7vKAk5Ol1lwzhGbTYfIFz9Wff7TY1zdmXefHCZM1cSC8EvRKPz0N
gkywn1sOVhbiRtQ3k/uS4n2yomEAc3P8FJqufFKBf0/UlCpoEKzunXtmKO6i
w5v/XEkKhKGjhxyjCvWhQ9/PiWn1eJRe76poULZAiopu4+xXfVGj2RNVUKUl
VaHVE7TwR1QcVek53iPyntGpcLOWdCWlRk/dbOUi8WP9P5TsZdcXld8FGwTT
qZ8JAjQCPmffBML+R7KIb+auak9hybj7/kALp1mQ0PVGPZgxIRdwUFudh3U0
kfuVu86J8L0zYyQYsTm7uSZITJ6SvRr0W57L6yuAuajkW9vMq7hLkbyDKg8f
Z8Uu84f9bpq94CMK5QzF0N0TvGrSS4ZqfVcnQEH3aJ/dUcV/Pgebz31jgMpI
mmYwhrm/WxF7LiMvZ3QX9tFCUfXad6hwMAhuNpaQVzBSIO+K0ihKBoy6rbuq
w+6wOUmBbzz+9WLkOJJlglI00aZaPYwye4+2q6V3NU460aG+DKpXtRH5nY6L
stPtLd3qg4XYcei29UP+ZBIaIdW8qzkzMr5rf5WKXAFIWI8C8kXMkS8MtS/V
iuxALeYphjWQOidJE49WhaaFZgHkoq5SYUK0xST+/8C67GhEwrbGMdHYCwI5
LMYsrmRaTrySBx2GOxQtFlpkkTRWz0XUCrSO5TIUFR/aGz6Y9o0er22u0rud
nON7/TtqJD7wCcIzQuohSGUkiGgZGAx12QNBnXoEvng1EBGlZV8cd2MqxH9z
iF4OD8Yq7avKRtaAF/uUQOQ1FiRDeC2wKGGSXIsFHUgwwoNJS3+TfteHRHZK
zr4uf7X7IOYyNLo4IyD38esArHpOEMndWuKjbAlGDf+AyHOTE1FJjmXXc0Ji
N4eqVHQCz9d5wZ3IsJcHUYXnUYJ3g45LWXvpjN/sxMRChAmjONrXScvRIExa
NY/QiKkdUM5g0KReY5Ygl5tlQ8XQ67lfHD2k+EIPTBTWsSc4A4kTEJgGAOyY
Aq1VJAb/4ZW84r4ZHSo6ULfOMEJCLu6cmkcVy4EOAMWGM9lgGaMHvEvh3JG2
QlSMNfp8SwlJX6IJn0SPFEJ1yggF618NZEdtEQXbWAtyFBJU2lRgeCEc6xoI
Owo0sP430DJr0rJUJi6nnBIczPbNPeyJZRKU4CCWQevzlN13Qd+WGHUal5lF
nhGzMVL+QIRGyQqJIJpyfTtUUaDtXLV6ZG6x4tHJu+DlmDROGjKA/v0BmXVG
/FuSVvx4CAPzN9k6+MhgrOTstvElh7XEA4INKDmcil6NW5EswpHsrJoTP8LK
rRYMLJTVS8ZaVZRqwZXhrAWfnwZe849+MNWEh/1a8gE9FWZ9XKwjBDSpIVC2
lFF512je3otU7zAIBLmN5HYXDfN/KD721pu7/TcF2VLif1aEeMWh0tjDUfC+
Sd2i27HHp3wpDPyQxGxEPDKBX4O1OoUYcgikbQGtub5bJ6tOrJ082HIF6/lY
uRXJ1cRgNIZXA5wl2tfViU/gFZveoBC5DgBlS3HLzyHOSfd8dRFy7mmKN9Ib
Qxtnl94jVU1mncC/YkGEkV7dTa/6QIdIdEzrQ3Qi/ZfPsQ8vzuIeDVAi5JsE
2RggMjtCzAqVVMFOEo2/oewemXuJcDX0lCEsCGhS9EmEnFHFQXCFgN6SNQ4N
WvdmpM53mJkXTDw2A9ir2xGUFRO4aoS91YXqiHcmrO7QUmqAPaHhFUM61e3e
k6bwVPFbf2aaBhHrnuGIqAdVa5TGGNAQiU1v1zMBJcXYSy1e/oGNsM0GF9x7
k0uV3VHzMfM0TRHhKiY2stO3nvPxUD4cEf8++4ymrCt5wxOdBgq7holUmtcy
8ZJaO7XDQamPYud8Af19/ZV/9CaLhJBv2IivYpya8k6CCCEqBw3/F5GEIqoh
LfgkZi2cDhGJuE+tIV/GXVfCl209eNBRAGM4QIMebpOEBZ1L0wtMxE9wLwsU
XJvIhfC/bIBiZrY04vg07YLJa65FxlcfV55p4GHJKlsUc6l9BYkNyJuH94LJ
q2dn4tl48Acw+9TvcBzSqX+k+V1uXFWj9fCcUD7Kqo6djbYkyqYwPLq/0FMv
8HUQePYWqnNFkMuJSdvUcUwC1b80nQb81wn/swfiuzmOTjLg5AF0Xn6ywheJ
6RTB80wxFypkW7NTprXX3RcIWYcaXgD9FgBbbPzxjL6EWX73DefHIuiNeb0t
nI6Ab+PNI7vEb6wlECbKa5gS+0xYdlCCUXelAmXc5tUnhu6DlVExFOZwCdv0
xHiqcK0UisSkvG6E+YvcoAut8PkdBzNzCXooCKKZlHfsnPY8w6pZ0Ze9wHlm
6sUvGGb22QcEZJwSdvRwE/AsaCa+5a6WDCxz9kYGmOYrzy874ZS8NKolObcA
OaVTefvg3awMsnNsdmGtGe05Atn2qLQqe/TbXKey7r2kMDY21oUYNJooN+wG
iTEazOXI32/fHlV4+S0dNkKYaV/s1VMBBLpNoboqp00mRPFqwo0oUAqlCZwS
HDQGJFIu8eNDEKHQw5iOhgL/4t6SgH9fofgbBpr6az6fC3slTi5fd5bIR3Js
Wd9lRclMH32DDCs6fWHm/liSHL+QwJJM/csqU7dKIAqZsAfuKEi2R1g5A3Xu
Ni2CTpEhGbC7pbxR7Td+AumsDgL0GyNGfE7EgQimkT8c1XcBX0ygiCZqGbX2
nyje3J6Mu14Gwxz8MtFXIIv7hSItKj7zL+dcMSzdY2VlcyFh3AYXHjJbrWwk
F/MBcP2UiLHPYUvluiuLXq55TuiOmqASpBuRb8BE3Ch7ozxZv2cef1wvvBiz
4oDk4XeB9RPSxvUo26hBn0eYg1dfYL5I25LVPiSnVkUwVd2O+qMOqyqrZYde
dRW6bCIH8EKZ3JtJJ65mDZGroLSz1ocEJFo6dpghz2a4f/BKA2+DPBo3yym9
Rq23CEUwTszJqHQQ9y9iDNK4tQ3ebFtjVR4rnWHlFmlWUBWDKHSDWNwoGG1e
0maDik0Fa4DA/nszst1IIXl8ef9DfA5fHlFb/sstO5ckDEnzB4fzXduA+Gt8
i3DIdon1hWpIqW2bMps/oNt3pobUh2sNqzDfI3R3eImQHsxzp0NHLZ1emkaN
kMILVaE4IEEsYAv7y3hcEQ2an+Owu4/U9XJJaGPtgnil8Z0OepaDSjzwjW62
fWqeNYZ9y89cRKR4BGcR7ecQUsoScRrgxm9CWqIg7WUOUl23Vg866uci2kQD
x2Y2T9IBOsY5M/j2Q44DGyHMgU9x1n5sTq7nZrCmSNTIUZvR9JhOVew46kGe
ER/o8co9NsH+RCnT5UEd/4WOgd4Iml9tGNw5yq3Jgrwve7Zp+LCPkTxaJwhX
XubkHsfc/OnCQg9hd1zwLjbqpG3JYFZxRmtkQbZ3QSgu1QkMKLDHfdthF6eq
Hi4ey4Ang1wNrYXQRjmno8dgmBk96n0mjGd9xO0ScTW1wEDhzjsjZk6xTXO8
hbv5y6R9V4xwR//COlqabvR/TkFRBcgc5GhkoLwJe2NShAAfj5inHx98QBjn
Dyqvn3jEhChBRvo2lvmn39DANnHKmdnWGWCV1YCbZmDUGVvSNl4tDTDCmJBa
LxGEb2B2iTu2JVzwSTSwOfJdg32WMkbW8J8tiFa25WHqZwXs9dOfqB4qajCq
RS8ZZJ4DItqmafxoT9jVnCoshxNJtI0XLo+BDk0slbtJFe94VoZCJBMiN5AY
c/69O5Y7OtLvjVqNFeGkVHFn/+ePBmcH91xEeiA3mgCq8YyikWFdEq1Gae5d
sM+14bCh7SQL7JisGasSG5dmaj5RuZWVZC5QwL9DfjxWsyR6pFlmZ1S9qGsB
wOVmEOMztloYFx9AC8SOtM8mN5qspnYcV0FRlCcN1iacfa7eLrP3Fwjr85SG
t4Ue8tqM/HpOI4LnBaicgHTxOLNc+z21R9ESB5ZDHhXlXODVCVOJY8/BRk9o
n/bGz00wnl/C2tf2hkx/3dC0ePqAX6CgEJvca8wxkCTtLe7uQxTFHaex2Hff
Q6EAWFKXDjQB5WTqPArnif7ACZp3MJIqv8lrWF0NOvrZWWh97Ld5ZQY9Xk2z
yAzqCfUdVvFavmVYv7tNRy/moboocyMdkb0abx1HHTFLidQ6cQ0Mi6P6QjMr
nDn9abHjARjWij0/SmlkXcHki3pMnPG71WVXDnflEiK3XHmH1zzzJKfyboPc
T/g3gvQUFDz/ICoMquatHK5LdaFi8qaRCFoYtlMPHaQLPsV2msS0m5njo2iL
rELQzM3bZleLE8rEF82/8yOVN3W6h1BsCxveXCkVmXuBWV3Pq5/eQwA2wOIT
TtgF8vKixfWdXUpVv7wtkqfamAEFZ1gPSmKRlhMoatCV+whIJjcGP1KINMre
MuPz5QGy49juzXXalp+bEX8er5PFqOZY7TVJg2S03GVs+0SWuZdvV8tT201L
EdukdKrXTa6ww1Y2m4n/fzsK3vwYMN/tN+uKIlpCxmsXhbcptLcG4X1Hpy+u
vmLDArHFrnksgai8Uho6sW6yaDiQZZSTCP3aLvD58EhUkz2oXtv4rvyIzB+s
8iPDOR8K/KR0OkmJQ9bmBFSPzFmtu5NO46E7fC5O6vlpGJzsK6irrOSD+3wT
2ty0fwLaZ7CNkdBcFqAjYjv60RJ0eG2sgUsWCzIStRTlrK8j2QStdmfZi1FN
O34A1aVsdBs+1wvcrGjl83SS2e0fTw7QVb/RMgjK9JK4IeQszxkHlLnIMNhA
fccbpLGucuC7OcmbyDnM/tVmVIU6uGoe4G47DZ3Vrx36HiwpreQ1wjbtBea+
dsrjJfL+fpknopWw5VpOOUqDKdN1gU7q9tJeT+VFy1FKeCztcSZLLetr7wM7
jZUa6Kg9Z7wY6V2T8TVx6XWdGZD/VX4jqp2mHymrBKIrsob14I5xplB9owAt
vOzIu97/9iH84hc7bA0bmsU1qp6nOkiq4Du8XI//4toVY+D1M5qUzUnnOWG8
bzz84585pHHF3LYC0H2dDSTGL2nnuhn2xx2cCQowUMUogXlvGKcmRQz4n76M
bG7rmlwDiILMV4xNeu7T/5+SsZ3uLqi3BkWaOgEYRzgSyjFXF2v8FeUBQ51s
WO9en9/xioaIh26rLEfFtSY7E/zSNNTzV9zR/djCTsOv9AskHEZPB+y38GER
c9ccAuasILfNBLveozajDST2FBFs2LpJkMJfp2hwc5Bv6eOZOZsnSE2UwaIt
Vz1V0l95Z6HyTavF1zmIWTxdrwWSEwlp7B0OgdFlReChtQlAVfZ4M8jMnK1J
/F1IPrWGk6SrH3Psho7eZeLHD6tS6Qa94yrLOsVQyev0OJzuJUqLIZUd1uHV
XvEmAreEbpkR6DiI9B0/EOIstnKmWsXOYuO3dvKQTBEJbn/UNF1u+qAjS0Yr
rvaj5ASJjd2IX+QgLxJW4XCTyjXCSNp0cnCn59+LZYHFAgCY7i071mTUc3Cr
V9coCdqsonVo/paH6lZ5MI6mK3N5wj8AgSX2951d7Tl1OSeoLhvfmeXY1g93
QMGesyEsZH4HdWB4l46F84wAF5QDA3OWamCYVcvLzj6LG4QucMnTaKlfvtHA
V5OYCtLMut3f1bXz086Q6SaKhEguAdFTHEOPYK+M1slnh9/H8W+lP3pcsovy
R7hEyWPh1rZI11Ls+vL8k5k1EzsfZ4kpITcXnqveNOKqVOCB8H24HrERdHiH
cbr4Gmg/F+fcgIkZ802lcglpLG3xZF3vI4zDXXKkuV7j8Xtgrh+n9mcIHQtr
AatNjeh15kXsVwovjzIVVISE2N93xv+mgLqB+JML4+MUq37i5cfiES5Sie4N
sNcaqxVsNTZi/ei+sGM5fc0ym1EIN20dsdRDTZ7cHD9a8L7X7pEo60h0orN7
dY2QfLxC09OIVn+NG0vmQ7QpTr+XzsVnK9PtCQrpRlVRZvJUXqSNugsjxAh7
w8uMzxoovURCsJDsQ+gVUiosE3ZkCnOnvGkbo4+ydKHJTRtLSzhaov7yGNNy
Z6QT2xHzCzhdFOreK2BSRhBgKRrk+BxqyGJJLfOcJfPf7tP6QRZ/EdfEvshj
6QoMkHr/hF+CusdZ1rsGb8C6c0YeWGXul3M5uFbNWjfPkexs8y3ySULiis5o
n1ZiXoH/KnJAK0sIafEc2PAebYmouXA6lE5VpQExs4UTaZ7cLN5HyfGcjPDw
zvXrMmB8AugKq9Uno6ncbHooKpmtp9keuc+tbDWpFKMYJME66u1CkkoxuwPA
ZpoJhK1jXFRjl8SflvLXpFz2eVGYwQbUlqM79hh5TfC9m/0cLJEmyq97IvQA
DL5xbi4Z5Wm8/o3ZGtMqudRRa/4C2+o7Kdf62NM8aAHvvkV0tSxZwm8NXbTU
4KxzEFloh9H1P6CYi3evYcWT7VTOHblNbdsnRlrd++7xCbBP5V6YZJB49E8s
8iEXmzOF5pqE0G0ZquCUvzbxfoi6ftvy7TvB2JkZm/hD6tPjOpZkuHBsdp5o
NVYhtdCG0m/ii52gJvOw9/89qwqNhPd1Muemvf6imbfaopjUVR2LdjNcFani
h5PB+gSdyHzygBOW/NV4fYrGPllYR0TyB8pf/KNGOwenXJb1MnMDm0LUTu1X
MPiL84tQoD5bGRd6ohRVq5ZhV/AmslX4GefOGvTIOxdIPf//0y+zqFX2ePmm
PJVbJKmGb66vXjbjAguLyhhv4EKSjjSOmPmFXjKWMJ6DCU44b+sUtagaiZdg
nFzAbz1nxunKZeybMieTvbkoc6qc3dwFyRXnX6PxoEVvy2iNRGsSZpvalE9p
eu6nBXHsAqsuWkyWnWmmpNEkg1SBA3z/9vca+a595J2tdtAJX3N0QXBbV+oI
HTBWcdH2xupd5n+ILJHAZ0ugZ7i86X3veY5n/LdzHOFt25cnapqiK+I9B+7K
eFjF0LlKKj7w6Cz6j6Evqr/r5YdjepeEbueJNqSTtsWrlsnXGEJXoOBHbrYe
Ey0TzFTJgrgNbzisUIBu/l8wJQzBlKmP5rev4XURZmlzj6dOwattti4OKPuH
q37vpQ+Uqe3kTfQ0Yuu1WWuC8hypJMSspoFjuJy/Y8KQKGbjO1GUoFbvwuQS
sxWuXGQDOLLW0SeqkjMqHDIwpIr3PXRZgWwElXfCZ4rRPgXBwc6EC2K2ryRA
CIcjMNsO4/9ImuVx3n2kVVP1Gv/v2lbc5/4VjHT7+sUF6lNyW90InLI9/AI2
+7LPO4en34hCE/soUCMzr6HqxAZtcKkKf33rXUibV+nH0tW5zFjVR543Ecqx
HKGyHFmxrYdlMQKjkjI/AqdMDvYtZjD9y9lF4iNPBiZ/NfG6zvzrscM6Fuv8
FJYN8Tnj9Nkk5G+vIruSXQjl09aT2oZ4seDvLToYVtn52oj9u8tlQ5hNCs4h
eaBjRHyE62gWdIhwqERQ2kIzcEB9c1FaidbPGI3NNGxmPicqGdUdHVDD6Txt
Zky/U5OuLctdjASzxCLmUksRt139OjGiSQFlb7rL47K3t/MM6h+eT9bd4OzG
cZ6sJdcmPdEAGmg751+EPpqgdpXkWCQjbv86jTRTczqel1Bzps/nyJpzj63x
KKHbWZPFSAYq+rk+q+OcskQjStsurRS473jvFO4Aebr7EGMR+z+fCyvCMLmW
/C2TMQRqDGApixIONabZcgCwgNpGKmSmeVAf+XevKg6d4Nsi1Eu1/7mvacQB
P69Oizv7OpoAuXwvTThT2F3Q5CnXULLtv/xo3Z//FB9HVxfGYcQgq6TyTOBC
MC4HYrcJyyo5vKzCcndk/qQVtgVTf/7UZezjKqG+wyC8l3aoylfhuZWH2bY1
hKjguPuiFOgMTkt+Mv3XYxS4AEjY2Pvf5hC5A1a19sBPsA/a4T64ToxdngZX
yAYGaAKOUHHP+tNiVa22NPKnGrWDNPHB/llVNO0GVETCQBhb9ih/GqC4/jnA
G517/KbiymsHZ9A0vDWtP4qKKAyPCMtjaInkXtVo5DOOR7P/lJBm9+kqkgms
qAtLEQc7OrT+YvSMNTz4xQZkkBrFBk/kL9BSjZVR2Reot2MNHo1mJNSqrtF/
VK/9ki5C0lISkY5SZhv4COgpNv9dbbww1TiRlq4V2YjNHJWEylSf4ZavWOvq
k2TWQC+/3wxDlNyKZ3ISYngfRxSt+2hcbc8fvM1ldnFqjYmQWgdlrelfMRQ9
3CgqtRhh2lUViMecoOn6qWkC17tf+oxqENV445KAugMrJnSuledVi+5mVDis
8he6UWb24OaGyC2oo6+0HjplGS2W7/92hkBR4Ld89QAFXSsvd7fKNA0KE6LZ
0dFImKvG2Pro+XENWvkh9hg67x3/Olx8zH/w29j/JZu3jnSKlUrh2rB50597
DxKGNUirtwDHLFZhjTKNAo65D5/Md5h6y8PMXhxCL6k/SEhTSWjlD0NWImYH
fqbjMVQ8kdWxiGVissrVRN/ycX/Zs3rrHbqhIub/nox1w10ZnjcV/VMh5tON
UM8Ll7YjcfX50M9s/bZoyh/rXlkxO/7uj1FZ54zXD8y1iC0Z/gZzagaRKMvn
7rJcQUOy4LUDdW0BVzP8DVMf5HffuLMeacB5tvPK77x0vMV/9HX9iqz2o5yx
lX8sERqCpADnP/LWuQXwy5KJ7Tc4wQM8uWK3TiabCvDhOMW6kRFxjoiZ3YCb
YlIlK9FfhXf+lGSpvN+9M0DxLISVw0pLsscUfWQYunMktgYIvPP7zef4Wa2f
wurzTO+zXuYEX83cR3cVtTIgsXI2RtG2o1GymiR4f1RHN87qe0no+tQFhkKy
2lkPCnspeaKXGkR4DpEhC60mTcrDE3bb25Ye8RblAZySEG55Kz65eqegoEaa
DU5vGduqB7TzRmBpgLeGaFbK+hmVCsxCtIPV1c2QFEIlkbgtW9yBY0C0HY/V
K7lu9zCUn3nEGIjB8xxINS5M2AaP6yQ5IbTtDoxLA51ShDDLBfKLqlVfFHnV
7f6z0q+KHv+J2cqytD9sFOrX4491naIvqRrjFAXBok05kBhAbOvUD4La3ofA
RvBW4z9qSXHEvCfxwp1oA87nI9qoYd8QouzqDzrEusG8NjJxc6Xh5MalKRo5
mmoUHJKrSSyu7WPLtGX2mtJQaO0TkfoDY5wO0OAmLNICnv7XqEn40WudpMNy
ve+VVAdZSBL7Ll2SuXIqfC20lz7gdPW5/kem5JHkVU27VviNJYBPBckTq0GI
H9FVDopRfqnPvNp5ulpmAlWhBItQLFrFc7Y+7mBQoai6xyr/mldD65s0p109
UngwMWuvO4by6uiS2r5BC2WFwwTATrX/r9ggTQWE7GZsO6Ee9y1Ftig8qk6F
104YmDmzLAb/bGkIm0xORelzjGg16iF3mEfJxCwGejkThwHs9lhETuwuOJ/Z
t7a6Z+v2jf40DMnhECCR+TnYiMfMUnctDBeXLWk7rVgzEqa3oKfIhDQAVpGf
oyja7DgUYX+KLxOulWy0BV/S/rRnPPdgVq78IdznlSgcagJBmxMvFzAoREim
kMpfXoapkPQ+Qmxx4WWkbK4sy9p3m2IqPMU+BKznt5/Cdc4K6subJBaxRACW
6APCKUJU6IVY/LV5oobPcu7w2FE+BGcEEeKjnRnr+T+IjTyMO76o01UrtzfN
bjni37s7vDy0mzUGVbOu125/iBL/zHDp6yaH9iMsn9d/uHiMQ4D9FLWPxwVW
VI8p3sJZvlgPC169utESWFjvfCNOKkBIviTV9rrB5SPOgmjIP/WWnjzI39wz
Sdby8eXokr38LQKoGdjGUrZfFH5kzboDCmdLuepFf2a11HhH8Eeg9ZCK3J6B
+XHQDPPe1mrl7YKsohMyuHvD5R6nE+oCr5pMdkl1JIBAz7yIEgGWbBT2F/i/
vGS4UplDV3AkFD0Ej80mE5ofc7YcUWD8lx15kIgjv8baRIXUcm50Hrb1UggC
eiL1BGSo7+bM4KfPmvOIL7Jh429nAYPQ1sy5GDA+Uahk9lqeJFOzmd89R0QX
ZwKigiHRWtv8E17MKGpbmNxqhb0/jmJmw/Bqc4Ws8MLq6orcDPY0Zpmiz4Lr
+ZcnA+PYYio5/GpIwPS3v+pEw6u42OBN2oVAuRdkm2FFE9rDycPgra8LqJXW
IVPXbpLyG+D/pcoCVW0zCZ/PloFIrRnwbGt6z70oK2FUZ9RwOGYjrcWiRt0T
aMPVHuDyLSQT/cUR6bbfivvTLxPLU2N981XZ09XklDTwx1FnSKPGe7ytfLOJ
1QXAP9opGj5H+voRzNrqjImViPM/QB+XlsBC5J7NDOHcAG6dcHivyyE4meXc
m/Ooo2O/oP813rYHh2J3DD7+oJVxYJM+Icqp33Gb0XkNg83GDmCb15L85WMz
YHviZm/2ZNLWnxhP68Kluo8vxUBKQuk94ZXg1dTCi6AKJi1Kvui1MMBFhY3A
m4Kx8pk+wuQXZroEORoj6UEqX7yHUGiYuVqwSJlT/9fIdd1efI5vlKxnXmEA
aLa+era7e2o3jyA9TlFE9P9QTbo3IgSMRFqLrngJrKRPQnzEkjaYlKBtMr/c
0Uh5mb3/JKnv6r7RI+2Jdy0UyyHIzvJbza+ilVcSI8+pJkWts9fQA2T/4W1d
lMV04ZUqYg31EFTEMrCY3u3FDaQKNED+VN388qiSiLDmFztY2WzPf8DJUVkv
+oGYKiSuMvus7rnXVRswsm4AOUkrEtbcVCR2O1wvMTotPv+rUAg2MNxkmUgk
tfjAd8Ir7bQuqacQ0w3G40bjWnb7/h6C1qfzdBvdtQlyPdz9hOQlIWqMOrH8
/Kxq48boRfz40i/ZpbREuc3ys1Z9CXghjgwptS7MZ4riKGD7MB4DpUWC6NOw
SJeDbAIetYfMUAPvqmnaHfrBDFCF5h3GjQiAipXxVeU8dA3R1eOeIBdg1iJU
sEuzEhzzAl5Wjc6qchBY/Rk7/rwnw4KiCM3tvyAi7akM+3NnwcqbB9ttAKFm
ndWKQ7zNFiwvzHn76LBYgQcR4ofr1mJQtWFeMXFvX91LcRNqMPzKnQFkeRT/
nSqMxzYs/PDxkZNfok8UFzgNTVte6a1PKD8Lm0KDmBBn3AowNuBH+xuKCbxb
e3hhJ/DW01LljgA4xhQ5q9eIAwXyoE2sb4VzUNyDgtUk8HCyPmQF9Ba4Y2Cz
bkhmx1WtpROzjwIMvEi5V65w3mU+KBe7tkITJCqXgrxxsdMklTWDPbeU4fcj
W/Y8FMPQWqT1tEhH0QLj9F+Rl1hJhgrraVFtcMsMEmcdD7fr0TKAMtCuz0mi
HWsGFJHeGTiMDTGGfginWv7wWGClmrkZlbwZaKsomafT0b014KNBsirrpvtR
+qfWvhAlHG7lvmZjcL813kU4bYmXnxwpa1/s/Ry5aRwXUxj1ny05UTabU4zF
QBFtWP6IT7QHWOlLqWinSOtkbuQJPX3KF1lPRQN4ccJAj7+JeieNYR7JlHPu
U5z3/FPfapy0+cUGxvwWVvL5DYki0w1cfGjtz9eDo5MkdRe+HVG748k36ncp
Lra8rathDQ6DvdGv0vSaCxKovLtVpeFniZhJ64Dz953ybdFpfuAlDSCWAWVY
pGuafjOtGrEal1RS83XQQq/QUdLtfIDy8o6MN6whhzaRUUje32wLtzsZAbOD
ywYnqDFLVKdyySUuEdC/Dk2TGJ0v1YSbUJGM+8bGAGTxARBC8tLI2Me738EJ
fO8VpSvrVwHGC5l5R3d3tMyCEmKhpNVrP+h+Zjbfu9Tx8N0OFGedBQ6TlJza
eXt2xqXBcSh4cImaPpjqo26xXaCwD7b9FPMqxNoRXnmDgIovRhVB8H1cwqjY
LQDIDlkNIX2BW3VcnWIWBIl6XJBQDMHoiQXy3iSBQXqbZC8IILW4wzIKA48w
LjEiwSouWKn3s+GmAdPrlLkyXJo6dWnrfuFNPacxbo8VtTNEvqxu9xgl2uNI
ApO6HA7FuIN9PcwONO5v5JSh5O53vTiIhW+PdFz4zC+krZwf4tPJMtz0Ggeh
aAd1L1Ll0Sfn83r60LF1KdG/j4B6Jqu4kI8BzyISfNrWaTh4wjglmo5MzvfC
bpRD3ubpop2HebSPwesAm8lkp+/3hzDyn50HYLbbmx8NOaQsPZe7542wtI4G
4mw4TglkQB41S5CqRDLQx2Oik7McCQkk7m7kMFaJPIH7aFFA06B5tdArvwON
7LNMtslVaIDoSvxE4H3e5jhemH+f6VbyAybiVq2ZFQc/W9gHb19Nki7kGDtl
lnGXTCKBMfa03kT9zgvySmoQ9xNQVYP4PYnOuKOpA0MEOWiKqxf2fwbBgfxW
3OkJNwR1GQ1YQpGwrBYZhoYP7QNUuYJ+27FCUltd7zGsdXBK1Pr+ty6mkyzP
I27tt7E6EdD5L9Dl3tcQxetCCZG4y5rJ5+kGiYxlolXoSWr8dfcWPPBgSl7H
cfpfmgzTszrtH1qDkwYhKjZGzqv2cNq7YfDW1LyuhjoRX2RATu3E9Gw/WpTf
opyd5yjX0hoL4lpGdB1G/zBoLy7BRWUT3e2MBpmufRAmMTcvYS4ptpMYmJPM
jaRWOAkV7y65p6ogybnHIbZKgGXS1l46+nuHCLM7oMEKp8UTQSoYekRNkT3U
LejPAOFZMHHIE5I9nW9QE9oStYm6UEft6oDEZY6O7fQZoB57hG0RhHu2Xtnk
9UY3iUP1+PIc8X6uKXaskMKntD+diuE36+BX5u39BNKUKBoRoAbOR200eQVh
lPdUhXfb311aoDxVkE4/FdjQcgkEjMP42nvXyeM7CthoNvmoAf4c09sYXtJo
Jq+fJgyt7uMpbEP192jt63/tiACNcgxHGIb4lbGC709Yp/938ZSvtOps65Gc
pB52nDwS+ODOC2QsRero2pY4RtzbJoq0m6M1RPURILvshd/caK0ryHy402X9
We3/2Hrbd5vif6/QZDoFUJ9M8lqe8innTOCX4yINJP9LYPT11iFBfI8MZ2lo
O7t4r+1OE5jYHNUN/5PovdLSyYi5d/n0xmEpggZUkneffq1feo5cPXKypdn2
pXVo3yzK/gcnLZRNyxL8Ho3ffqcdgFpzz3R3PX5GtcNvr/i5PO4yT+5Se6gc
jY91WfGINADoZX0RyTfqiWeCih1cj6sMEkTILQ5U0XD2SGE68rM1r053JVLl
F5UjLBKBTW/LPK9lhwbM6/eX+Gzk3VY47cMnRQkiSc2hQH6HgFLr5NyyjP1J
UTKNazcwlJJfjMRm/cb0cApDDrrDZUqJmXwWpBbtuWbPtfCwy4dRm9dto2/Z
TAPnp4r5sVBicvkVnt4QZUrxWhJRRzFBoj5yimgIWHS1/Po59Ju6a+Trtx9u
1bd6ra31eNwcTNtcSQWbqkaGvnWYY/IoZex9QffRtHBad9OmvS8BvkJnxHJU
g9kBvHj3CNaz6/WpufF6Sbtis3T9zV5Y51qIbPNpdNE5sqzIIbnIstgB22Tr
mAhLWl2UFrsYZ8nyYbpOSKdoC/bvYFzNPGL8RIU2pZRryD/avDU7ByZKILgd
nbRX310pXg0wy7ftVAIDfEm6B6BO/lN6ave7iMlu35BR8C04KnYbYMB4c2im
hyH03H5kA6+bY38DptmzmX8Sf4dVIHjceDO6CgXlu8KMjK6Ot3Ks957fnzmg
tDa7IDz3gOWEnZhJPLBDxZqe/CxTkN1ufhnkef3tjIuBsAuY6Vjiv10ZmmrU
TxIhtzmBeOQGongbxP/hlIX6nEfF9FQwDo6LQiLfBzTENDITb0hmPwk+PK8y
E2ZBFYcwNpqqdZO6FAElo8tc19ws6kvII4dS5la3+Lvmx4i5J4DeJYVz9RSn
lc7MRLaKmj3cYBsFMIOdJcX/F4btzjIdmlVItYjSXyX51zzT0Z3M6Tb7Y32y
Yg4nL04TBQbmf6V/7jBZJA5CmHaORWBR5L7mQbC6C0ptCOgvSxfR8pfNoM5R
wx0/o673VN8Jcxh9r+J2vvmWiJFByatD6ADPpTRO++TYq4nwM4A7FX9IRLkg
QhB0aU43DNf4XiszQXTIw4pSqEiTe7yOGcg4aby7T1lOKV22Z/nVZjtECuQZ
AOx0DVj5USXxvkU/2QXjaL/M1qoEBAi7gG5Dgxw3zZB7WClUe2xZpKjmeKkY
jPNlphS7mdy8fVnThTkPyqEiSOu75G+IcG3UUGuVlXppMZEszOoNSiXHbc9J
9UQQOz+M2oywT2uyym6cdqSGC9wBLOPpYuLXPC5hft6cDnBSUzXmqXVRh3Jv
4rFCttccymixwKfvezOT6ZSphbxFYiGxstFFDFRh27zl00XsrYh0HXa6HYc6
wccZLX6IQIB3nsZX2pXD1nlndrUbCn113Ixlu+kX+EdZGOJyJfP3cA25d+E+
r2aMtzC1fT4K/nSz0bdXGPNa8HC3fX80+k0F2UdObdx6mxLYo/yJi5Ab6UPU
uJpm8oKh2IzEp8gYtUBtekAQ22TGEiVmds98EkZsc2RBx9z7S8blN3HNyQ9U
z5dPbb9eIKFTWmyV6Hz8Xx7PO8QfSPJNPFlb98/73yFGeFJEHAQFY2PmhB0G
D73kXmAjZnezKq2hSKBue34eOfatdgsAX3IrIkVT0kHXcfrYDioIZ/wX+8L9
xGP53E1RvFIitO3R/gxtNNX2uf+X9z8lmnvq/+cicnImQrIgX5SE+e81YVfG
LJs6Euo7+C5TYAcafFA6NsTDIa1wkXLTKVSXhAamdb08lPjH+C0IcS5KRLVB
wRLAaWBOj/BWShczTmdzkuiCHL015S0H8tfH7Mx6L0EA9p4fXXzmMEq3tXW8
DI6+Vu9N7BsoDvwe81+Q4rk5C/qHYONSc6zvWqcpt06opvYKGUZuqnvJJHC+
OlxedTvQx1c9ieoOWkCrX8UpI08XGuJt7YfoBBeAyA1D8Ub1IAFoo8UMBHaw
ThglkiiGuQl4WqkwTJ+CEAILtvaDdhdNJJfPBGyPcMls1qNl32t9CusWVr7z
hR/5pLnbulm7g7aJCkXznW3zNuR1rwldImnEySjPdHoU9KuqIRpKUmKcEkLJ
kDtjQXJ1KlD1Wddt0wdDHOx6eIYTpYwcqH8z66PkgnaNCfhAKmmSPi0sxHci
cWsK/dakeoVpl09fw8YTy8cF2kn9wkgWzSxhntU2NzWYViuZkf11Q6rZgc+x
KWJvkDX+e1iAkDzp3/Nruq09LQ0qQjO1LC9fjrkZohfybFTN/VqbLurxNjY/
blLIYpRH4AIfSszx00ZPBK7cBg370B91bcK7Gu3n/AfOEyby9VSXCA8X2Y7U
4ROVoBnj5qBzrOxRbo26FChPNsp/7VjVS3BZofi8yMoZPcveJH+uI6AvDcEw
u5g9EZVBQoH0njYAaXLbc7/1ibhatlj52x3C2WvpsChMCjLjE8r1qg8IOSul
Md9oTt0Wlks5uwVGMx1dp6iZlBxsHpbZsUOf1ZmofS7sBl9yy/1XzptZrq6b
wQQI5Hk+gqkv6n1JAi0rTG0SXHu0uJ2EkExZ0OX5oExxOKNT1k9J4lEj7usE
/RS9x4jraajwcnUN3+NNs01i+BfDl0r50uG0Q3QHnZCOfTdrE+v347bCkU1Z
eRJPNijU+ACYunSKGiKsMFraD7aKv4jvzzfu6bSoHTPHChUwc45P5fo44W9l
fuf6ea4v2jM3uQMWnLoY6mfHdt4DEvd4jsK+Oao17T/bwRvxT0YSjEDjiPe4
YnxNqRsKpXylLIg3mNtNJMbSamRmoItBo2iIk5JkfhasJpC5AZkcndI4TiuL
4SnWwR2X/J2cpUv88awmZrB8Xs85Ns0qjyqGL9g/GfqQybGaq+jY/JNWjz3M
uxqRmALuvS4yEZaJaEgWkVnBftfJg6zKMmL8gWFfFwTTzpbD00cSlpembEcd
mA/LzZj/PNEkwY2IBi2ogi52ae59JWuR3wY0EwSPGrP84i1vg7+RtLP7AstV
R5zeIrxcnmSejzP7aDewOlwZZ2zePb/XQn6GajND3t6hMQ57eG5dOCbuQqID
yxrAuZa3H1eNsm0QZEyYdIelziLPKy76vRfeNZY429YKyrw+ucSQ/feVBb+O
ys7hn/c4y3JNTEcjbSOMO5rieakYI4D3+1NVqBIkUP2RaIEyoQWYsbyjyM8o
BBIfiol8sDEw6/EF7HZSuvLJyX/DuMQb7s03IkYlSfSWJccnrfdUPYqm1Lpw
GA3CzVLygRMZHkO5prDBsR8Y5V/f/2CaWjUkHsAST/lqm18/C9iOvEOxHCjr
JrTlmuAq54yMnt0TkJMhZ80EHvA9aO92AYTL5GlkyfG1Fs80sqVLjP21cQ1Z
1i92PlJ2kFGweDu/3LqpzMo4+Mct5tR8WAPTSacFNPFsH0S/+je0tX8HQ7+x
3DVAP28gYDHhKwKWwm2KjIXBsR/3ZMaVtOHct/1e3ue30oxWKqpjj+uWg0zS
tcQdQltn6nld4JvCB3FMNQgExrX6dMtnjK1JN2QDK+hhZgHPwIMeKiLeaiHn
w/hdxLgtIS6ISI1qXoz0hpCrnKSuJ04gnYMNsmQl7DWsDVbIdwtJEIZDT2aB
Qtb5PbKzV9TqTQnVRxCvjs35ILFc2cmJrn0xEk45KNGjOvcUXcDU4CLSlDGY
Bwn7FfWEUbC880P+Ic6MaxAPoH80Va8nEDooh7iFHf9JG2ylrcado7G0xVtX
m9ZSG5pXrVZTLe80cisSgL9gL5sVypJzCLlXMyhBiut7ikWGlI3YRvF8Q/gi
RL4L4ncKjqG94twZpAycixngkD+tKkZd0GEZ5NedwRKe8X+2ieaYjnaFdiqT
sRIJm7EpEc5w6+roZuo/7uA8ZHR3EhIJXhQY1+f+bS0fKnu+SNooo87heufD
jiDgHx/iwZ63cI39AeXedjwpneYNIt/fnYUJyjxiMYmuV1Dyw78l1Z6FRUow
/Wl3DRST1KI143XIxPBMVDkF0voMUNXpz0MNXhCLHIlE9Wc71wR/RFniw22j
jb1uuH1AiAV/4lfaS4uo7D3o55k7XES2bVibDEL7f8Ec0QrnallXoA6h4tn0
Ao/D5nBjaG5Tvol+IgBCtP6r9g+9mfWcPb0ylcZH8gRg/u83CVyMR+R+imXI
DEmwrvDL3Awrv4L7yx86mg/u/nE0XKiDhFQRo4P1wohf3VLn9gCam8KUmJkY
FUktCIUiVAvnGfL/vURDx9R2KYb/vaZ/LJJdZwb5pfqgl9YyGBraQ3E35J18
0cNdzsRfKDQo2YAL32JcBKqcqCVpCBehSVbfkl0+KpBk1SomrUDUJUTFVU1i
N6urL/tTYU2y1fxkrYv5y7sG/0KOpA6ChLSHVRfz7LYLLFJvcc5Bui+3XFgZ
TKj4qhul7FlCd2FtX4WdFBjsEQiNrEWlAb6ORKJc5J/3cMVfE4Y8uS4Xdrbs
gnwMLxBZFor5ii2llUlj1kjDfeOjf0t7CNqojkJSOppwQiYctbL8Jx9VP41E
FGZNJcQPsMMHmIlsFOd+3R6sdM8igP46AHxoA/7isyGTLdDIuuRByGziY+2o
13BSyezhLyaBNn8vC4N5DLnzSCIsmI26Mg+l9BM8PMHN2us5oXwQ6oplLWKq
XHbMKd1AUYJNgXNYKPTVB+izI85xiV40BCWQgq6uMzDXxwe/fuO/4R7ba/sv
gkFZSXLChuV21yERJpCbi5LT8jAz/uXS6pqOVZpKGgu7IgzK4J1TQCq+E8ie
dr+01mNM/Py6geIh6ujxjP0NqZajdEEmcohJl7BSKrJgDNVPz2A5tqQ+NS2Q
0LyLij3t0C6C/2e+UG5U8vlmWAbZlsBqMONQQcsET2mE25Sn03/BqMUoRCD7
T/zV4vgKtUkRP1qWLSihSJLtqIlsI+p2edz0k4n5eW0mXwlaqU0u/b7DbpOC
E0VA42MUzYpF1og+azEVXdJF6c2G6/3JG8/mPE/6PKBVwP2Yba1iNpWmUfdH
vH2PUjEa9fQtRo6CrkvsYLs7zfqfTXPKX4BQaScV0fjDXti6rBHbdl6rFJyp
ox1GKaaVKDRhVLpCsoPm9k6jI3MXMZTi5zZL4kHDG9xCmyRziQ9iaWxgrbj8
RolUqDfPp6Cd7ISHOj2fAiPzQfXZ++MA519WQm3szC34QMp5G5vuUkRPhYQp
BOAcJMvcysmz2zsjHk0TcTpvz1CR6By1dWukuYUuXVw7tLml7CKIXePmBbVo
EQaAzDo0wSr88GeUEC6Q0r1LlniEi8GRElLHBwenDWtmGfNhBXHsw4JJcrH7
739LzumTMv3FsKgqTxSZhYSbanNi87K22RHbim6KKNTR4h9VKS7cWrYI7ESS
YYrFu8sf0Bs9C5QIYLf63v9thMrQHcv6zJQD/5mL/O8B1MncfR5q1iGdV+Eo
mLoBqsvopeZgHEOVsFUJuYF0ISKYVk/ZWyndxUIiMLs/osNZUH3I4w971lLf
nilTB7ChPfoKS2nVEs6WSYD4BPuPpc3O9pdw74URAvtTQ+OnMrOmBBXRIdY8
R7umB7PgQBkmv7/xo17/5V4HKY65LH+zzeeSlH/UYq9VEUC390wTIAqyXigB
RKCvmIKMrhm6u4CL9qnNi1IDQJMfv/x8qtcEAYIVQTjp4m4bTCJSho+8jMnx
tUy5q50PNslJaCjgrjpqOw8/6yKrQ73HrEylhEZ0q/Rw1ciHgz5MIl+SsWly
akkG1FsFvqz1WcJMp2Iz+4FaSBP/mufToSZTuH+D1ha8UpBPrrTGaepAA0sa
OuBCv3NePCeddmsVy1sY0PbLAkoLoLAMgbUtjqEwKhwtlp3sYKhcuHS61M68
zGrArtenzs39nu9XkPARbEkSKOwKCXhbaGZgA7OfCcPnX+V6I1WibiTQQLjy
PU7QYMwImpqtJMPyzu2eFJldsqVkLiJGq8s9SORs0LVxhX16HrSGMfz365Oq
SI5AMWwuQ0YkmnbtiercOf1gvAGKLGgwIRk1khPzcVdDvHoOJhuq1DCRUyjT
uYX2M71NW1U0YEGxR2vnNKcJdXsyTtrSP/UE1EG50BY2h9t6MHIettH2LEgU
cnIU8mquOGzrS/ltFmdAfuVEib/6Rv914WQHtpP/kcg+wO68UHY2AGdvkj28
KVJLFf6lr1LSAFlVm4c/JAxB1tawDd7c7LiuzqeYiOnBRBfHXbSen2UrHLBz
0eo7AVLxJO0UfbAGKU1Ys3qIHNe8dM3phCG3je2l8pnRrI2X9j+cg/9sFtL1
eQBy4z/p9zcepoBY6H6xzNYplo9o4CCfG5OgU3wy7h/+T37L1d5PWTMwO+NW
jG90o29Jp36KVY73SX/j703WbmEV42VJNXJ3PxrHgfZ4XSF/4WUHYLBzqqf0
PL4DiM6Rp1KIpo8y8roFFyySPRatWOB8xAszLckses6z48Mi+rJN3gWPtnwH
+QAS4aDatRJQEO96ythNXR7CkpF++AyuME/CXIgCKW7SckaB5Zn23VOT7DvD
h7mm1udwF0YXxyeGRjz0ecvmZmrsNOUeo7VoVLPgIqBbPDRU0Yk8puCHMuiH
CS3SQJU3xqksuXmqdf4rtjYFm4teWcQ4SrHw0df5G8yAtJ/opMgpzaCBY0Es
uLcD9Gzj9Bti/s5x7Xvf1jUOs9SRbLT7w5II4Z3Cz2Gk+EdqBkeODjnReaCB
bNy5NicDcXfEk6mvnekzSRPLnByx29Zlah0uD6wARh/3eN8nvqHjXyZRWPbk
99yNRm1gctObdP2TbG1sD+DKKYuEJRPVD0CDksFq64DpXHwPSBRP5byCLz5e
7jzQj80KNI/+KRDd+XjpY//WIUc7xYM8s1/fVV9JVAobehlS+GsRUhWFhiaE
HqlzZP/mZVv2zlJpUus7F9fERl9N5cSLMEVBNtjgXMK3+YutoZsqUPHvHdb6
7nregLXq+qZDsWwvoUE33y8AV9uewSEjow2ClP+LCgeQkqZuCZeGCac9YnZ0
ZDqUXqEDThcyXvSOfHUAANpFGB54zE6f9WQLphxJQMTixbfa/TgWEezzc/ih
QTQJrtE+6rQFFBnt2K7ZDQ0/0VtKR9SIf+YSQOLmJJHbTJ/p+uZNZuMC/W7p
1P15Z+hMUnitCCBhkenF+/W8iuRJiw8B+3ewGhZm0BSC91GyCfdlx1WDwaXC
v3ZNsKUJFvvrRO46AMakQ6WFuM4+YB5eoNehsmlNGir57CX27g78DOkY1y65
s8NHQ9Ux2ZfJrxQvmkoy3FUg5CRMgd9e8HvrjCSem3TwDQHtv1/KZ+/MFidw
73p854WnKeEK0XzFfXyBCbxLxKispneMVf9HZnDtOvoXmzzwXasUluTBhmPT
2DkRzGPFayjHwhrrfzkl+7IXsZ7Yqvc3SUqqrZ2Yho18DgXKEd1A+MiyG0V0
bu28zaPRNUQCbe20yVjYuZl4WLMw7F9WZQQNCM4TrQZdZ1KS1IoCE63CEQJw
GykgoLjc1iJaT+rHZ6fbBqIc9NMOmqeJUd3A99xiIqPGEJe5xEN0w1vxf53k
5VEki9s2HZklkc4m8YXzFF4Sho9kQSXOOtCWyCKADb3INPEQ1Ut71FjvNOeV
lrBPb59NJaN95qDQyHqam3hyVzN+CHkmTMzhEmPKw0SuBVaOe8d+jdQ28k0C
yMmXydxwalr6vePzKIBOmw2Lj0BaCRIXCacHZwBs0ARiJ3Bq4ZQk788LCXeP
hWNeouMLmZ+yNcnyDbbwr7Hz+mJjTy53IfrNGCdnNICTtlHzglLehNeIJMta
F0wmZgG5gz3IHEk4n5cdOz42PtXd3fj9Sd+sVqztftFn54pmJri65Qw+2q5f
64f2KxlICRcekw+nWSNsPMdEw/b9HY6CjDPNUphalIn37y3ymI/LfB/O0AZp
ivkcUeqviEU25/ECTtfajR16mEqL53+hMymtzGVwfDrILnE0h8Ul/2X9hjHH
7mchUm5dexz+NrlxF29x0dPOfELaAhrDEEmFhEg9WcvIBIhDPA15UcDuRZF/
a+1uJ2KEdR14FxyClsCqt4GDRYi4TXj8A7qUjuD/n07Pas7POxKQ9Uqh/3/B
NkduPirz/jgpzHDKkuHLAv9l/DJ/mDgRN2PRz8VtzJbgeZPdPeGD0NlBJlbZ
AYd+ruDRRQUF7Yk7LfT6Og1CIKKH8P0SFh3NYtt59agCNZA9E8ACegDXIWAF
yaBuoRVStZeY8/i9KkBstX1hjGW1RDl1kXgT4cuydbXLj/JxEJIVinhYq94D
MJEZykgGeQVTZLBOFs0VeCmlXiRXXKMLOLVDER+QEbmOQqcGemxehxHyi+96
Iw49FT1jqk5orEtHlRJC+6+7HnGqYbuQTPWp0IDDs0QDpjWZO3drA17SONX/
RKruxnVm7J0kGVkf3ynqvM+00iCVgGzQqF4/8CJFGIXPhN2KmKHHn/fYwkME
h1m17Ftavb3W/HkXLl3jfHOWD1iBYqCCBvDkch7Z8ETeNetO2t6VHpOEF8cE
fDqTChqvGsgbhvjj2w7weybST9s3soOuO4ewOfx8Ld/XyKuN31vkpIw1lRpO
3E2WUPXEtvzDTdbWBZqknyHDdMnsPZeCiYSaD2mVClbr11X36Lz1agmmnJ1b
ztbb+SGIVPgUGrZkP7VAHIMatwXPNY+zRSJyJOmUCvuBaGR2a+Y67RYHGRYD
6ForBbUaKW5gKk+RlSK+FpUCLnY5dovUQwnk0JioyKtEc/dbLfwVPXaHOssf
BNW0yQtpDjOZubR32xeXZaN7jQmM8vdub2bjPWihkW3NRV3waKKdVvsM+0yY
mUS34y2TkdL5AOM5a2NzRm/jKjeUXkZMME/sdsOQtEwUTSWuUcj+lI8y4L7Y
JnMs/g99YbV0fgRs4YrQL0t8hGagr8IpAxQXaZA0mH4sbGwTr7ABKBfkVd0h
4m1DBtmPb6KTfeTwZKtTFGvRRuYp8R1eQ/dsPV2y6wP2BJKNpt6nUrc6um4e
8Uzlyjk8FCSx3eWq5OFMVq/IB04AfW7OsWPXIXrbMxRMJYRmoCM1dHDTOwUu
75YQ8OoAjhK+1Ccsn8nlXZWGpG921+Ssn40p7Kg0Fpw6kJJo/fsRwZwo8r1S
x6PagPsUOXSm6giH92feWNoqYmUPnghxxYAfbQVHOsHVwDsc3PZx960jsUdB
D0ywj7Dm2W3Hve1DTqPr8wG8ApPTEojX/X5xYeMCh8LPVWKN6F9eZSzqThlX
OtwKkeNIJvBu6hXVcNqJi3GcH5iEba+XIfE/RbK0NzCfmq3yBK+QGGN4JnPp
BNpNnX88B7ft+EUpKBYHVZakC5Luwtxr3mZJy3H8A9UYTHepj+A4UovhQivg
eP+exJ9IJc6IMibEq5xQAPRT+XYfAPV1QogK//hYmfMxVya4IrhOEqympPqc
MQjxItiwsn0UGORCiqWl9K5/gmbROuB9Chn5/T1LzN3pgRPI8fbaHwS56j6z
SB0CeGojX6kI7kgBi810GEVN+lCY/f5OYPHxbvuzVbyvy2h23zhr2bOyk3q0
Xo5mZYMMzzBrRrL6L7I+xrEKyRitTuAt7vIMq8m1y5SYalieiNEAscw+nkB1
gJ/lVnBKp7PW+iQ/1g+LPrDGag2YYhd2tVsHzwIjvOfGcMz6Ft0rlHulZR5N
9GYx0Noty2XHxGwxwuZO2fYjIs+bwIF5uZ74FpqKCaCfujTpr78rIqKj8DGP
N8wP/Ny4PSyrMFrhlws34gKKsAepx0rG33+r8jsB4FnHQEKcTyjz02wq4tmx
6xOXZUR86KPEpyiUyhazmdDlWovmjX2/7X3DI0lb3OgB5FIRGjTDsU0tXEnx
wfsFQ4JosJ06d4acCYb7ie1XHjpUmR/2M9FCJ6wroEcB2TM/5tB0grXiCL18
VRW+r0qiEVDY7qF/w/X4awsaKxFRve6zsoEKdErOZp/IH3mI48jI8jcKeLOh
MuqM/SiYgvTmTTufVt9K/NrFXiPzNPR85V4OmdpW6U9PdLZnFS7sV1LRu/pI
67GLFYaR3g2A1vRE+RmjaZLylwKCe91lyFDXMGfZG+eH+8i4GEGf9399ZygP
dYfcaknioC4IJDwK7HfjO8DTQU0fRjyubwo+DO8Q5zm3EKiAMTBpuMvCGbrq
WQnQmNBIFHeiYXJNsmU+BAF21t9FBr3pYppvLukAEtU/OhQScFLN+K/aDSos
BITeYuzc7Ima7HILz3URp1jT6QeXskrY0QUAdS2g3RFNCJ4e+TSiRMeMNI9o
Vn/fsIEy5xAA5qDmoKtKa5yj28RpIDQNXf/+iZSSdc8FCBxJTJlu8mArCEob
otmFtoQ7ZPGhrkq0EeuTQ1eB6QYdh7JDMb+6iU9O+IRW72WKv9fR/q5VCUab
c43nS566lH059RDRKEsbsVIinX4iFGx3B0xMCBqgkeHfsDb24eoRTCUX2tAX
kDp2XEFYMXgmDeT/HpwEH6q2gAeZui6Q5Y7RSlb24ugwdkJdXNgVlyfTGv8i
Iw3BD7OjrPYWatZmltyBDy9zWgw608Wv8LHMEgK16X5FXnnr/Km0ODP71i0O
wNm1im9BkjtBh5SyUCKogKCN2MjprJ19oey9DKZLtSw5HAPtB4iaJvu10ke6
pFyYPLD2tK73CqVLg0inL2GL72iFhCU+yh6DUqy5ORz0BGZkf4O4dH2lT0BG
jDt/ICUcfLltQmoAt1FmoHO3mpfZvPB0GFttOVMjUKSnG7tSzX08oSZnoyfa
/JOX89ADZyj+UeDNPwLS1Fl0SF3jers6WdAOEIVgPkeKSawofV7FA+2BVBLP
HuHovSoKZd062hhKRcLf4b43de4zczkc0qccA+EsqUnN2s08k/CrbdzlSgFl
W7ImJQR4JVaFd3haKI0YusNw0RagqFhvEz2QISLWjv5V1a2dbI3mH2H9BGrF
NfgHGUSYvTxRrNRGVZ8GmVkDHlwPu7a+5xbrF4Tzp0wrm3lyeHJyPmSKAQn8
Pfupq2Uh5fAHJr0IKsk6CbpxWZe7o/LhuA2XA2Kf/wJoQGYu+mfy/pAsu5Xf
DVccv9AmrKIEeQm7dcmSYHYFOwR/V3CHLyRevfsoDtpCZL1fT+I5gMz8eS66
KB1ITdExqcuf3DLjwIPoM2CLloEfSoHtOSs4Jb2xUF1U0FezDpJROitPO/Qg
wdbLE61rFl+trb52rRtB6Cadej1mXV3Lg+DLXRk8wtY1JxG+yCQ4+XIiJxV9
nymzytmEG/umWKxXz9yiDmAW1FOWf82cvADtMK2FETGxI9TDEcl8S7YSEBr9
yklzoTqx0CBdQWyC4RnUYn7ZIQi+6g3+TBQocRhtXYdxV1+Az4nYczpoaJA+
5Af7XzQgsZRiNwDb6Rz/So8vTLNXRVoIvJVKpqTZMwfR2FQDMAtuLIUOpL4E
9rN2EkKWIMQ0BF/AABDz7Z7GMi0yaBT5dmjF3VtjehgqpH82mxA4Daiwjkuf
0/DRtbd8pNGU07U2puH+tCCqochKAlcyRPnlmsp9lVL9/8MsocXlMsXAs40k
mppUVweFxZ8TNpRZozP9OzowhXbVl2+k8kpFRzc0bZyrw4qMSzsaTdiiXz++
Mo5mGAkTcgW1tSV6H598Cq/VS5fWHG6+EDaPWPGkAVzL8JUzSp3ch7HyBQP9
2eI43aXOOsCP8IL72PV24mSvrJAZGfYHBCCOj86+/QvK5nfFv/Bsjmkiis1B
apYeAqKi/Y6kRvK0QU/Pqvfcszw7fgO9QwxTFBdQmXqduvPaju15Ibn/CZ87
GO+ZHi1T4uAQWus2PZl61QyBdr0HfWlSj+tzw+XUiFCVaqhsQhZ9NA6uIle0
1FznGb15Z3K9PKrsQ5jhaz5t/iiiGxqPW8ACUVu8J/9oiImDcdYfyK9zc1OI
6+IxJm+AUP7zCO4VLai6KA6Oiile8y4xKs1MB8aXDKc83v1I01w5E2TxdmmM
x6CmwL80oZkHbIK6G7zhFJc2YkXOdnVkL7jfz50tYB1yAEFaYLAuqC+XEod0
JF6NnBWFWOStH9X909v71/uyxSgTQAyOCkivb3jV+itquRWlCupNcS1tIc62
Bunbw7j2EJ6I0zaqmRUQzTE6yNFK/sx4YLi9Bw3FWrXyPZld7AdelssOqI26
l4WE6r1T1AqQXXC/QFtm11XBtLIo+161Nih0BiC6Y65bMbqsvtratfm5eTPO
xYX129tCNXc2m8Fg14svq44hUjizE7r7OgOCjVQgky716ggsqiVOz5jyLPBP
uw21rjA+ic03UPxvx6WGO1aVHkYaISF3U5NBT1bd01dVA8P770SujvQjGpiv
86/hFWprAePUAd5YG2bH/2tjocRx7kWLsRYH3PCaRd33FWp4g0EmuAaFGkx/
79JNl5s00YZT7nPEQdh+2k94MzpneRrRqFEuztHPGx/CZs6m3hv8ieskU5CA
Dg0c1Ne4WHtYKs9MAXuaxS/54jI1qLM6snyUoll2edmqgI6XdOT4FF0ada1z
IhCn4ShAZg1k99U1aCAuj4feIdQT3807XrS3KWL7IB9x8Cj1oS3xKZroM+8L
Ty7UK5xOveiJCmHeMTT6V1H1xYEtpEIiuGVdBisn5USEm9QuOUE45xyuScFO
FGwsUycPoG6NNw4kb+2g7qpvkDVYtt9bQeCKuxFbstT51f96viDEiQae5W6c
P/F58uyGLke1lI0AqvcxaX8+3UCEhuq/ETm3GTD1FEIoJP3iC8sXJjnFN+fE
Ikh/snhCNmjbjOmB48XP3/NUI3GFcOwgD6w0kclOy8xObwC7tSnJQ35Es40b
RKheBu53GYBzv6ykEmYAtDZWC5qELE1+cq9DoxRo5xAW6xd2BzzQW12qLj3U
FlFr/H+fCD36I5ngiPo8h2ZMnKbrZrxeWK7Uo0jblJTyj4S6VCBss+vU3Y4z
rd702sj+En18KvbI+VtgI56/QlrfSCVAqZl5CIRqqjwKL/6ceANISSg1VH98
taJvKp7CP8vjb+heg0Q0RWSdneX33efQtHWdrwcn9h+2zb5XGFobYmBJeafV
8k8J32P/BKw8VOVoN2uxnwK/2rG95vL6KYhFAr8H/at+Ijf0fGNOcWfW/iqu
V4IsbmFzJLdhssLGmlwBIDJADqMPfnhVmm0rz8V5YRxnXAAUStvcqypsTPQ3
IlQYKqeaoya8EdY1BqUIooJ91WFxAYSHtWsIER0/Zssu0TOiOr0L4BE3Geuv
/B6upug//y2Okx01F/EGGr6G1AzLkvZK3R+CcV7i6wtI+1R45SltUiplt5Es
MKNkpvk4ducvYOfjzLbC4dOffT8Yf7c93hFPcM0xKQALiPm1Me+1YA7JzMX8
MTMJxvwWl6IODpk+sNaoEm9PTYXPyNemK5vNveWzo0ecguk/dqSVxnZ//FPu
C0mSLREBgRDxQAisLoqEaHdTH1YNz/3nhKh11bOlwcuwqU6Iu03TnxIHbGUX
MSPj77Hc4jhn4xNH7L027/ooGTZBX2E52h7YOZ0jTZM+bvRtTaCIduEIARsd
YE7a7iW0y8+souuDWFf1hpW8tjNVRnkEJNUpaSoebI/ek5foaVAZh58omQJW
dWcM7RCnImAwepn8udXyyEJxWfu3ubGDAflfWcxtKLDnY7kmjNxzPzf+ZWW3
bkjHHi+bHeWMFDeAbXw1ddy11wYqdeM/kpZ+BTq1U1ckbD2EmCEiC8xdJJRz
8bqGMWBheaRuS2g0Xgd6wwu9mTYpHS0oKY5kCNhrwc3/EW2nX9P86vJRkOW6
PHltcuxyHF49xAnlMnb/FF3GZ7d8X1HYw0HKrUZRu2bwbZF2sNCxsl6EEDNJ
STi8hXPOTaz70EjH0jdpqcHTtpuqQXMLvVIk8U8OO6zBL9gqLoBOG4Fcl9lE
WilhHvBg9IwpGkj1SDTFRtlw+8bU3guuzR9FDXXwXo13fP/9kGpJtN4BbuwF
/DfStqxQ5mKAEBJWt6JBOAKfltSV0dKMOvlS5PDtSq/SRfHU6coWUTqUUBcp
x7iEghRWICdsYV1jHsyjDBu39+iSGIlena5aT+Xt1ANp8UECvZzNjORNSS3v
bhe+G+yLOoXjiWEYx3yEH9Rx1ypwDGXGfHxdtwJBkWjJfzMH/R+uQaSLUHfx
k4NmZ30NLses9tGgoH+5O7bzj0v+ntSaELmx332WnYn0WwvHzAX1JPOliC/x
M9ODXcIDAE0RucLOfjeZdbwUXBnuWVoBqzyqCpEolHRqm7ofSAfZQ4raAs1c
nYr8xrrwjThAvkW67buSJRdhtI0A+6RPRv96NX66DfWTGu3qT7EsBHcPgKrA
t6rO4aO17e0aR/GX8u95iMSE+SYg/jn6lejKJUpirN9dhoGUJ1mnwymnn9jE
enZpgePUSvI9YqKEiCJbFbDCHaHY1b/cMEFZy4XxAarspDDQc1dbKzS/s4R3
VDwfC1uSNe6t54h1LepVzcEg/p2eJkneie3iRmUos1zTNW76pS7+/Jqq2gxH
4CwBpJrd1401VJ64uxKlojN4I8Kg/sZbZzn7L9Syvuw54nr+k5DHLR1kXsXv
7HISjto4Afa7UsT7KvgInurGna7uYPs3uaxdIe2aXyaTd5d1ks74W+KvK3GK
eeZc5dsw2bB0O4NWG2rr4PUMxBJ3ziaxGQ4oNhTAIs1P9rE1EMFH9LGivmzX
FjvrDzMBczVeQjt7P0Sp6MKxFOIq9XcqUtpXd3gmFvBB9y7OJB4rtRC77U9N
QrLKSBsaiPgp72gl1Q1hJyJD8mB8mLtu435NmxCoXPyguw/4PlWFW87JsbOI
mxs9s30tp0Livsna0Vt8EfeVcts/Zi27wTzXZriQ2Y9G7RytuwVhO+ISoQ96
4JtrkAhYGiE63epoj5iAC9cMMXkVEUGUBTm6Ro9aBkhl+581UsVg6wxCBGvY
LkkQEYswCu5BAGZ1iBcIh7fMwycI1+ZNpdxkV8yUj5sg4PLWU1XiTTU7wXRj
AbVJBXVRKG5jXLuOZ2eN8oIsBLqli9AyhNE5B+H7xbvhnWipOtqzCcYCz8mS
2hYMsMgeuKpgGlH204FnOB7c1TKqucwFAnPdwRzydsfTQzlcH06OX3UembtG
grxX2kpy3fyMtNNJZHymwUJ8fGz8A5yH50P+vmRFMzPFwmf5ABR9uCKysNGL
rIRCVhOfJmqVOe5UAKyAW5Cgmy4w4Ph+XXfyBfJc6mOcGhHx+Bl0HUIXHfTK
NwP0pGxNg10J8iuu1iDSxLjYQ8KQSsAeTLi2cDNFZrxFZOJuZ7A9w+sPr/Pl
1F57Ep5NDuWWV1mC1q2xDV31jOFNH2X4YhwfqnCXCK37WuwxGDg0+HLiVru8
99KO9QK5jYTKBXepA5tdz2ziGLp9NhndrBfVRDEHPBJaDwMZjxnuKEw4Y/+v
0/ExcmZPTaJ82fCXEWX6ftUVkeBL6E9ycnMrYfnv1PSSG8i9UlnYQU2AFkEc
yiKbBNjXx+10Tl6fh1m2/yp9YqjJro/SF5nYsEYNahZWIjWQqU+A+cBLKzPT
NwsnBLExfBIjEAB7ubrIhSXE9fAXOdsRI7nWJxyKOpLv67DDfttWgQtbL+kT
MV0EiIe79TLHdsfpVRGQzAgVoKQzyvs63E4KHf/mqcYyS6yTG/ctPwNkz1y9
WlTiiN+3M/jorLt5WB/V9QvUbGFMpG4PY80wkk8fLcS77RsguZWrEUDiGhNN
L9AwPMQ16h8EG1Dhen1L/iA0AlOHYut/T1wo98Ize7IA+hA5T0JtdHh5hss8
Btb0ItZN4iKwtIjY1QlX7+q19uiDEYvEywiqY4bueab+zcd8MKraszcY0ccj
e7UJAsuByaagw+Ql42SsPu3m9QHLkIhGhoad38nsivJIhfUxF0x/HO2U0omo
9Z0tKFfzvBDQ1Z94U4jzZrWII5nhhULLQlRDztFWlomVj4i8FjH6gZevvPX7
N1yF9WNsIdp6ro2IfVfL1ehS3Ji8uAbC/coXkhDAjTvv0GuY9Eg7J94bF14+
A/GuZOHXYLHMb4dYPT80Yf0gFon4z/gdU9L4ozhpAQbBluJREtmKz5CfQPs+
RXrZRC3sNoQtkyum/Dkwb/f62zPCAahaDm2MRfX6GQgSjssZjXLLhZZjEE+C
+PJAZPQ5JP1XyCW2l8j44TiTHu4O2Km5X25E8w0+qAu95h1MaiR+TpGLtanS
sK50Ct5U6mPf6OFyQB5iP72Jry2yKkb8ZLYL6QUg/pN1diFe8196D3o4o8HV
4U9aoLeHZblGaxVWed26AIDwW8yl3jq/9NWFMdUkFpXkdFFhUaUvLwQ+a3Wf
HWZzlG3m0d17dEFX1VO0FqpB69P3Z8DjhwzEdW9TH61akOKcnMsxhczMCrFz
DIJ5A+tY1r5/N+rwAMC6XLePjrK3A1/4KdJeDRz12LSMJW27LFVK9lxHkeKP
wO2BTiMOpk1Fl2NKO8ZDMI0I5Ac4gzgL/ol7uVVOQcZjM8f/V1+nx0ek4sPg
kQtDVqLtN9RVLppP5tE86YNz1gKnuWu1zd73zEIBJDz6YHQqqUJ7IlrG3fg8
Y9nNI04caAU6GWhAA+5IM1tBN86Layqvmy0Lpw7t8b8QhkCs9y4ovfgt8mBo
iVprRpq2br1ch62W42XrmYrzc/Yd3IoTbXgN1U6TY6YQBeu45mcXsqWihqzr
lZpRy3wj/TrW/676IlpKGNij1TxGwQl1dX47SDEZNqouP+BNjbstSd0cYept
DvPDNWEfnaOZCasbGpYmBmoKJZJAzcfL3brVRoNhiMuHen5kFmJHYWMhWZDN
+aPiUkT2Pj2GGorvcfNa2sOTv0uuN6clWhN/N6xHeQCm/4kCntyjMrANWoNt
8KeqJaUAd258u4pBx/FGJ9RED9LMTK4fywkQ9+xaU9jgLRawdB53EnkBtPiN
Vc1ao/MGt/nZ3YcCXwVPotFiXj9PBPWHkrUX+065QR6FfS3F7eUS8/L+REMd
28eLBjRCDLHIFIlqyc5zDhxGX1/liapW6UZg3eeHFMDl/+XCMK+sqNFZ9gZV
1RVY4CFdGbXt8gz0fle92Znrm1f2dEa97VmCwNLkDthXUwddAWDHH6gx8yJO
VEGKyhwGNnpitFEB3MHGvlQaiVGcKK6sKi8V45JdPNmLZqKJHDLdnLOsEcSV
YJAJHcV8lM7QrFQ6LwNaN6Yg73YfF7yR1wo+j/oTEhb7qfTYnRIDGhknAeYm
yyrkCNHCjMXdD3pq1pBnteHh5LwUea3Txa+AOSFcQn9oNAoV4XJRVGwk5qIp
xLeWcSjE01MBhX9u5CZ/u0Al54mm0fQ629Rsr/k989uHuLJrPtcn3aJVYrB4
jXbIl6uS0ESi7/Sxx4NV8S0lm63EpgwTjeuIwdnpU0nlgNOIagnX4pZminrz
zMAVacugirED52KRPBwjue/bF3X7X8JlclERQOf7xui/NfeQQxxmO1KLTuRr
CiCf/KE+bP7R1znmCWdTai0ySCihIdkMMVucIjlPVgWT7jrLT9lyT+Bml0Z9
/4dLBtmDYgfFrZ3wkhZh8iGBRZYBuz2V2MwUpjxsNFE0HOhMdyV2u71plDr0
0vdNNawhES+D7UEhFKLNO4L0B2R2ajVzs72xY6Kl6/KuAFFW+LXvmr2bkP2B
2BZWsLuV/+mLyaGPOa5266BtO7LySvkvBm28u6up/JYXH2WfiCIbnnIPdArD
4EnWK/MfQTJTEQ7WXKKtmcs7cli3iXaIzMPRdZg0G3EXkJVxeHTdzfSmXkOp
Dg1TQg4+eBLhSeEU5YQyCLqde/rirfbIgr7x3OhOtd5Jb1jGhS8Iiypk66bv
EqpvK1tBQDrirtpgW13RbEKKQKlQavEU/PAF1lUNHblwFKu+T+6rstFxdV8A
Ocl1uQ6PNY/jhzh92HbyU4xEuTeGFRk27tFdTNRm2u1ZeSoqOAMBF6pvcvJP
7DC16mV1dagmBUHQ1lqBw8tiBE6KI/F3RbxNFQ3+x5PiysqkgISdqs9IqAJs
8ttnbkeU9oIg74TQ8bnpZNjPysHzSbnbB66Y69P9wf4TvHkag8HNCxC2d0PI
1xdFNoeltfyYV0BIH2bUSew0e356xczuOdXgnuJQaN5Akz5X8oGDv8Rxet7f
X5ZCah7vQ/awdtLJCirkzVITYeRL3FqqCwQaFcK9Nwn9qWeYa8Y6tya9iBiS
94CmmXfPcI9QtXOeYMxyvxNWv+cZ/iqZv9IX9edNBjdCrazQko7odQ1F5b1A
s4t6Fxr0D1bq76MzWPv+EhOFV7HSzwU42T+RbsffT84FtPeEWCzyo0Q4TtE4
GVZGK56EgY4yPWyIQow6QYkP1dJ2JknRF8IEbrQzyJhx8dYlDmmZwJKJZPs5
6gZwwzP+BOZpvqYR073wB3bDVj6kJ5oKgzUFQFv5dOShOvFS5HIvbPaH8AjO
1dja5/ilRQ3mFyWq1S2h5xFkhWswFzJobKdUZg3X0YgBKGAJRbjwBO9Iy1mG
a34asiZfiEKwzs2MI9/sF2nq1qCNKMbjUVNqswYaja61uqGIHP0eitNq2ZvN
/OVo8J9VF2gzNXUp+Vo1TJtU1dpQfACHp6uMVKNmb16rvIhWGzXhoF35aA78
fQ7sCddiGl1Y0jCCak6WwrUaTQhhQm2FPuPH3mAja+/tMn33/pFh/OFEkoix
TpzBfAhYRkfgdexBaq+4oML5Frif0Tn6rheVEs/XZ6QIIduvkioTS+ewB58G
0nZuks0HcLHhwsH9cxHfFFEU28aGj0Jah8Ik4F/mIvRk5qEUEHAVDU9CwehG
dk65irrHIvlhLvqij9eqI98PCRfwaiWq0NiCENdSF2GDJM1F0I6iyWpkqCtW
Isf2h+R2kWhB/w9Cs7GsJjUtPjvnyDQAK4mRQsCFdAB/AMJCk7cvm8EUgtj6
xLmnrdLxsEro0i7YDmr4jgbM52IxhH5AvASiwd92ICPxQVF7+9pHqEqzKxwr
6bshqSNnIXcM6oPNV8oNfZ31NZmDezDzWGQ7NHt/JxmjAzrQWFBtnf3ApjyD
8HSPCbNhTk1EXRcDGfEdYvnZjq08m4+aLpfjbP+NmbALYM/d4K5qcvc7d6gR
xsNrsAUvxP/L9i0q4yzNF4mZfreWkM74jddJ356rX83Ha9OQRUAN4sqgZD61
k5pNyGHFpYgBZxkB8uQPJ3cc8SvB5qfPa1mQzefGFkvTIjWZ9JvI3jBWREXM
l9BMHsuTvBJrCfPV6IjpSkw62flDxtbBvy8HnVO1tSk2OOJ6wxQxMkTlmghP
EVcgiV21E6uc/8rIPFrI5PiqrwtvF3qh74uoZCy4ebmO72hD+THs7M/zfaYc
j4g/wgd1JiAMdxe04jo2qDDDbU/oX1cZVEAFF6v3G7j/hSTX5Q9MnGhi7DOB
0esE9M0vgkXMYVNwn4J2LoJo9sGURz0kzTbutpgYYwm5a9cYh7vRmh4MiOO2
JoyQirdigeeOA768mwT7W1ESkQpD4Z/BiXWUAXPU2CEvz08GruLgTRTn2Fk4
yvNa7FSJQljSCvAT5KFQx1ltvZjDH6nG4YyqoBNmC7RzAYPlW4zpIWij85yl
2mKfHbT7sBL44Rsx6mUquHtUpLJQI92s8YVXoQjKqBPaVPbn53KbomBtjRgG
Zz6DEOsmzvRywF7NCxruR2nIhkpm+zKjFsgpLhlfjHd67WkJyR32AyWOelR8
5mLuk25enxELr9cG1r6ayUwO3KUjZ2qjzRzD+gL/24V83v8h4CPjIpd+PFm+
AF02Q+OBVFNFP7AN2G9kTOeaommFSKk49lXpYVTVHF3sp++JeZpOOjN8fnkY
6PvBwq4g4jxGYkYkbsY+aLPZeawHk5mRq4KZU2I6eOrxO2iH6cYjOHRHlS9Y
W7+WixFCVFBE51RFVyIFeGtSuByn3X4wssff5U+qyhIYzsOlQHL5SxbaSHFn
psHu8ezSQ82nIPf5KutVLrYPtcOAdIhXm6A1BFEF73AZ5FbCZqnjUlVks7dN
iiUgXLZKLOHwL9e2rnHG1cUbQNkqze78atDUO6P4ZeHgGtcueI38y40IynVL
hff83tymhAwBcpqSYpuUS1yQEOXyyOC+5JNsQTmCMTyhTvRgMSg9XiJ3kSlE
SCi5z05dygMRcEnL+vsBT/QTOO1cLsooKuRU45v+J4bHfNIASk4yGx1RLT3K
tWi2lMpy0kR9c6tIcZiBrcopalW+cTSjmxB4kSvU9Rl64BK15GuI2NnvP5s7
agELVpGBCU4WhijdKc0NFr65Cq8mb1UL/U1vkR0zvzQ5H2H9ZoaWb22+OtLC
uqXx6QFwDxhDwqaZ0+W+QJnowOOC280Jr9QVFuhEQZkaUV0WFneCe/f5Iv7r
M1G9oa0oJ/ry4AO8pWiX8tjaPbDulF8sqOZ7KsLuLIZSAOBliCt/PFGC0tRo
mEyIcPRjIqLMtY/VXNqzAKZ8zyTYgCUHLCdi7YYMBIWcPaUQLxmCWvGSX7aW
flqmQN8sT6Vll2OSCTySZObPmcymsh68456ciCPQx8M/FlOM0d9SghEbmsdT
LaB5qKXM8FPv7dFLdXfLPEJp32kD17DO4ft6iIE4HowAH7p7FYmc0skiTd2W
mVEnpWyrNOAS9Y9b3hXxzTUVo4uFWjKw9vefiIwIAV/hoK1JibMAnnbgZkQ8
BHsbBgadj2PzRAt4F3FozKBBUcfyoAGk+5zACf2BllBsqxwIGhTvrslYM7Vu
0faR9i6aOi+HaerFrwbt/KPvobX+x2X8Y5yYWUlkVqRTYabfLmt7WcCqUM0t
i/0Xo0YMQBjbZb7IT9PfpQ1z6hq+Z7+IqiQBBk7bXu+AxiVkoXwOI7PZ3Urs
GEhZ3x79vim8UzJwtTKPznEB6DutqXwt5c+kIZuxR5qAGva6zxROKelOGhjF
yCGEjwPa8s2K2ykA+TILSDiTx7tT/vO5rnL4gWWjsX6gopFlBbqgGvrnlV9W
2J3QyYMgipHj5XuoHXjOcN88tXVrDmpK9s9c5GRgJo02/87XpMl+9tf4+Nu2
/gEnq6q2p1N3JzA/dSJWvsFy1hPBxkcLyFQLOWJ6gghtYt+qjypkpG37nNhn
YOhdnkRVnYVNMd9/55y/SuC4f6E2/71ZfLJLArMPXbc2KEK+hQmgK/LriBpX
TWXi4NV7CcR4iinhF0eLLSdDCIaoWQmwg3/+PfYH/v1a26vqNTD3s1xpppiS
K9bpsjuz8/rzKZS5+VujgEVbpEqJaaOiN7XBdsuoR3cP6Tti1KZOZZz31L6l
hpwBYSjoKvNcEiM60PQEq8UfMGHJyvqSySY8G8BusouT+jH5pQvsXtOXYWFc
MZg2sfdPvyGTyw8JVs5pntx7i4yyBNA1eDiK962E65GYUEJqjekGRmQj++6e
PhlKnzCB8MfaxQVVqZ5HTDT/o51hreMj66eZYDhokgVsetlowu9I4krMLEkE
b/eWaTIbUOtwEpihlYviCI+K/K1K68/hVxDwwxkM+EmsyFtAEEjJg0ccL7T5
V6L8uY31XZwhp7QrMNnL9aM4gfALdqP0CYpVeMniOKJfPi1jmhe4B7cIkvv8
Jdmrx9lM+EfRLxax3GlWWuml5A9k1e6DeK5cm8IoFjGcT1NGDiNOtRX4cUbW
wpwhmkfUlR08V4lzFYeuKKM6OfntZMxiTuOsSV6PLXGUGEpZEZwroAtZe+x4
dyFTutGcBMaNGNECbq4Se8gCWVNHdl0ZLju3MaQT6gWULnnl84rSVQXf5sxA
8ub1xE1eA6AhIOtbJqqhHjYl3juHSq9z0Gg4OSx2Z7MqXpodreMMbB3dn2fS
OKb7IdcfdXOe5eJ9pmOuml2quJxcUun6HTYemfJfUJW6edq4I0uxTILrw3is
AkoyUQw/h+kjuRM0H4oGIpRyiQ5PKLtFXhuhFekdwZz2pLVvXsEEzWh03kIh
UChLptjTj5VvhaRsBlcGbLZ/HdQuNVAkTR2to762iIi2yQxIQGFNazPLwEGc
mXvEVFUhV3efwDA1MuQi87eMenL7YEtWbfxXXnbCsSsvsGHeOtbgl2yvZ9GH
noN9sQhDv/hovmUPy4D21f7+zEwpbW8o8VRbBgNBQ2iyybA4kJueAdTMzRci
RDw5mDE04uz3MlCjXZI93ySWpHLLi7U/du3Yg5nIArXpklseHE8u3Tb1yTdg
F2ht4Yuxb0gKlcb0iYcYsnMhuJ+8O5BcQncLMaPCf6AbV69rRSFLODjvMVmk
Tf1Y25wKXfIXPnlWMQ+L3eeKfkicQN/qwU8oTvWkpiNkXda6Mo5hmpSYwc4C
1qKQkMI1XURAbRFxSJ2/hQ2SKOAo5ExwaaXRyFmGyyJIzApAozgRmxPqTodl
6zwsPXgEVycr3dQ8g2br+wd+cb9F+n3BE1joLTrRed3PZukQy+EBZRoTO3QJ
zFpu1V4/W8kVvCepRtRW/hLVQRyd4LTER0Cp4I7+3iy8UqFAPMFS6Yb2u6K8
kG4nJ4R99mHY83vM4FUh+VR56ygofNE9zHN5qUuz1UKTlGwlzwRNQXvKmPyS
N79uxFVgd+weWA9tagtfrt6qp5mzSf89WMGZQNOzINImJobUX1Nju7djiMLu
2xohqjDby3IdX9r0ocUut1m3XQjpEoMxVBz3xzHPeXW0nfdDVLO3NWEU0Viz
kpR1v7OsSS+xmkf6eDXHrnKYtZa2DgLnb0ogqkhUfNGGBwjt2ZhJMZdEMjdP
J6mFaGL0a8HsASrWwS1JYFgLh3WfB31B2se+MyaUPXfnVChrlkjzGfeKF3UY
/+qaDMP3aLLq0b1ESQ1Zu9FHfd2LqtoOP1Tm1vECOHtzTHEHuy5qEGISF9NX
ELvBlo2joIRx/jrlddqM3xC5mr51IRh9Sqmj9PgczaBRUFK7KMEBTJXPcA3L
i2W5tTk6+3f2dHSXgCneCDaxF815ju+R0eApK5OBzuZ6yk4ixGxCdsf0TOQM
qO4tcyQEI8q3/7KLPAhYxogHbWpOZNNBGhRBW6XZpN9i+tfMBnSmh1GYmifU
K4sDaUJQsTsY1ER8ESr0Rhtyz5IQNbKGp7gcRJUFOWvzU24KHE2AxWI66XH7
KHwDiX+YwSIi/9s7dJAnxuiva10+Jn96eouSOrATxazuTXzJxjOXUO81/LNx
nEeOXi+9rlLlWtEU/TOUN5PkWVyPZ2k5cPuy7cnRATjvSX8EuItxBxNCTinh
t7FGQu+51I5GhGV4PUSrhwnBCSYJ+0bpPAb1K7LIIfvRF5v4Y3x4AJIY/srV
YKOH50bP1b9/oZnkapR5tCCn19uBvD6JDLMZAA67LcyPil1a+M1GuUQwoG66
Ik0GF0mXUQJj1HUmuIA1487V7XcWHqkVEjiCDMZ7QZRy4RgoERlcRHsF36n0
euYpiHMVBkufhQX+BPzffLBfd2WRToQvIZh/Q4MoW5vX2FWja1b+8Q9rH1/Y
TC0HQf0urrDS6sbY4o8/jfPW9brIRJ74dVDyJKACzLhy3HikbDslGeg/9B/H
yUDY9sWIa7ZI0Vp7q7UrXi0/BiGJA9vxxMDlknHv87YRNlfUKHGG1M2j38FB
6BO+eUfPaYul59NIXGSOhsv46FP7lbREkO5CI6UhkkuFkts2rtp/xX5qlkv0
PCNa9sq+keN4w3eiM0ir1ACklDILqmquh1r9a/U8opwDHGEsoyLBZPAIHJVm
lFJFhkPe3DVQtMJ+aw9p6tfjIT1GsAber9UMjbaHJ1Muf7QLgPQF49FQ3mF6
s0Dg3KG/48nV/9NbV6TY1WkzH5bypcJOEhNGDdwEdEOiVkACc4gPyFJbiK7d
WAEmh0Emecep5nA8nJbCzKJ2N3D7umGqjyozD5WwdTZXOUIXcLSKFYZw+ZfU
TbdcpDcTjIF2SJqdw5PfTKFrQPgk4Q0BAKxNe4Se9XI8gV4BABn9+uKAOfbI
Ol2opqqHFa4VylkUqNZFtqG2Gyk6lnKWZVlICHiN+tr3DJWZv5rc0agJjoSV
AIW1UqCVh6Oe6ynspqLgazV9WYIsbc6EsruYnrVoRNFg9/DGe4VM1P0+JEPT
z9PBtkJjvkfcwCvevDrpziNUEZjxUmVyYxbrJaRhuBEnFyFF6n5Ht6Tlb8Af
IlVBDdvFb461PPUqZFS8eFgx2UWSP/g9ug/CJ6mytLdyn5zQi27C4vNz1pp8
JQCYfO9d5HysAq4RpQ78HZx9egvo5AbMnj+ZZXNkDfMNK6AYDwHX5l+xFFUV
uMOGIHzRYBkT94HcPTJSflyV8j+ElJ+CbwOkKDzYxACOwB61TEb7pABsBV93
9nMrIZKmNbqJxDwWi11s8iQtNtyJe+A89A0T+iaKsGGa2eK9ZwzDYeibJsJ2
hZcfgz5UAPv3RlZSgKqN72VA2eWzTgYJELpqAvjjMZkRweYVu8ucwNavONcd
7oQSLZMEuaDVbX7sE6w4Nq1rSe06O6n3U6ijLUYoo6hfaS8L3j24QMpmGdZC
xKymLh/IR43LFcpJcza+uuX9v9ml4L2IcHPQR8mJNgBjKR1JRlZgVMTRbIGd
28bckSJgzHcyrGEiw4x/8yYp2+YT1PCrxpABd6UMnt0CWmqvXwIJUqbPT9M8
mxcU8IIio+OyYiqKwN0hqOC6lneuxSFlTsMR/8u81qtFha2HEtW2BL+f3cA6
4ppqxIkV0/1JG8SRvlu3o5+D0IL7NbMS0koR1HsOIfkE/VChxDg7ls2Lh69t
cv3ebhZmD1rXjxzK8UxMIg3FXP1IpumY556dY7FoQKBHRu2rstYs3KwK+4oE
8JmNLSkJXcp903jr1xmt1FTWmtAbWBDpPYoWW7McnwAxmQggf9hQw/Vh/Uag
J4s5qZWiWDvyOq2gy0TRzVtlYWkTaucJCsMfWRfskvcVSuW1xp9hUZTXbBiR
vHlND6ENDT7Q9cQixLSHEUfEBF3gbegZ3CrPOtcYor2NJRHfBiLrZCfM9RNv
bmHOf+om7RQwM8IsYpBqBYztmvXMEnoxiJkjoJHMtKCK/+gYBMOA16dDT4IB
hE5aJ7DfCOk+mFMRPygPc+1Yw+niLKHl87MiGRhXpyV/y911p0NcTePYgKPn
5sKyTd58lGI6WJ7TRlSGcppnvJ12OI95vQiD+3ZdgzjfBMg3wLFCu7qgAiHq
brtg8nUE2oiQDB18KwmG700KI/65d5NlsZ5JZSp8P02Vkag8oqbdk8JlsOxl
udjv6gwOK4tVgOeyCZYa0Klw8oY1eQl1/qaGfHSNneD2nU8EYFrqv00CyvHx
/tMk+23u6VRGVkarqudaFqls2o7DaJvWF0BWDleY71VUSFiYo4h2PR6lgCos
2tA6wZ7/mh/uhINTQXcxg3kETUSHGk2J4MyFQp48QSghOGpOfqSc8OnWCzml
R6PYbXPIkSuxNq5j+5IOgrEw9eHSQy1lTX4fE1EepUiKVtk6le56+YSp994A
b+xlNXo3wFpfJrVjymq/SPnIguH0eGExxbS4uuwPIr7itKKL6MEobGPKUYKb
e3f/J7yVRGcGcaD8Soih6fPj41/K0zJw27CjSg8X+9XwPm4Q2OYBL/E0PQoX
pl91fOfmFhwHcdBlINqnBzrdC1tJ/Tyz9AcfCTEnJnC9hQtSqbYel8rT0ZT3
pEHGEZdSuREPsVdzzIJkfCutmUFqPPMCodoegZKeIGLh4iGMsy7s6j6lf9tW
tIQ8MnO9wYLNzrnL/S/akHAmNl1etFikf7XNfFNHrzcYXdpR8OQxcRo4Axea
/5mfziRdz/jQXuwEJ442JXP5/n1J6WQas+SGrImqOjQMi1upki9h0cTxnqV7
ztzHsbeTEDauxwvUGqodeiW/aiF4Dk+X1KvQ9L0bpQnEQUQAxaGE3kzo+u4z
Wvu3uup2lJoUyH4gI/6U3CQZHM5cdpscyvWCAmVm8puyF88YxPlrlGXClKof
TjwWSquo7keAcirq5HWRX7A0/8XJb1A/m6N+e5uDGD65oYOWivwTnJ7BD2cd
RaO4Uqe5NU2Pqo9NcvV9iI39HeAmRH7shdhF3JHbl7bFI4s3JWLtfiEyYJe4
6aCK0leFUeU57rgwLgATgCmxHHLDuQbV41tairvNhd6plNIOOYzzBTFF0FE5
mq9BQS5xn6J1NvVQlkrkQcq1upsXQCG7FkK3XZ5CfAOvuS/UPnWg4z5FUh0v
rNa5kOOZhhEQtKPEZyPm4E2RNeqomfQp9RCV1u5O2JBrjF5CzA121stLN6F9
ejQuGZYyTi4k4da30WFsFMp8qG8R2dp1oKpoUrX5MYZ5NHa8qAgQ6geua8rB
bvFELo2tjaw0BRYFTENm2l4C1ATMa7RBB1jvpV5PdHxRDf8EtNcGnZAehysJ
LgYL4spYY8zRTzhagyG618Q8C0wit2kGQGqLnnmJqXeUFoOx0GehyXBtCetc
TkxPggKPpMqBbldRnsfG7IKxqEmaMhVHZ43xXHoZ8mHt5Ri1t/ufWGJpFb0e
l91B/b1kYYncERKgS8falNhOStr5Q8rYY1hA3EyTaGumFWEGzJp8aMwPwEjP
f9LLTEej2GKbIrNOjcQ+GKP3DN8Sv85o2uWxnRPhQ3wRZAjC1Xg16Fs6hMyo
/lqIc8hs/jO2dovgo1HHILvtG9wLJloLmKxceglDqCpGW9Z0FtAMlMvIfmN5
t8bEu55cEiuSqGNFiad80t3guEyC7/jFgZlLgzlHjyeNwd2iFY1AcUtndw2F
y3XwwvFFWVf2fAqh0uckXnRlrQLXNLHhv1W8QBYw/Aot5ypRvaU7NHpctfds
XzYxZL+iKQ7jLzfPdQD/0lv2GFDwokOCQLr25Q8dnPwUR2X/3qdX1nQi+37d
sgEbsKWM244d/EmM51yKbdadQlVXgmYGVVuj+4+bOGTjsVhFE9gdC0SwZXC8
LH9j8US0PrZZmk++0ah8nc6YClCKBugUPJ5Ayma6zc9ovsiKn6+Rv+Ica3eR
0+O7KgFdfWxfJ9OmUEqM3XrMx/skFuOgOc5frN9WNSq+fVvLZWx0PRYTrr9H
eXxBwERKdWvkTb7iRzWPY3UZpuCXk1wifqEfMfx8c9Z9XwJOpHgQKUCvAptf
RnypfL69AGT0SrONtc09n9nykLKIsa7JT8BBzubZZFAIKNCkO5EaLmKSXLIQ
GJcrlEYwq5pOns51OOBCtvKm+nPTrYw8aTIcVmOKjGwCt2EFmI9dOpTNgVvl
TNBWfZzEcBCNisOFsyCy41SGABsRwiKeFMhBEzx5bCgUNtYRbGH22aWpgTPz
BVxql80FNP2BVVSr/CImq2TCFtfu6LAvXzKrrv6dse43iPC6JJ8frs++7kTz
TNR3bCcN014QdNovPyB+9FxZez0L2w+c4/XLuH3k1GpZ80sjdl5dN219I7Ur
P/Vqms/j9L1i1qwOQapVnmKh0w1ZCPmQL4NOSIjbZ9Mez7MDoJcRKKlmyCKh
UwBueQ8/IyIYEsZSdLYQOLq41TAG++yp93if6Tl559f0y9feYoRIgAPuZKyd
Cn3+n4hrU7K8HEmOHBGmhGsW6iaBoVCVTFwY+nmTLujOjsXfjVG53rCL0F4E
39nLfVPsn1SBf5D2YpUOJrvjBBiuJXZgaM1UuPP1giu8TJENAN/K6M6Sj9Wj
oCzeQ61vNJFvv6nmArS3JjogxOII10KLlVq+JbbOuRtR9pH7YIWuto2cuVTj
H4HPp781pRjvvbXS1qr+yEAePNec0O6pGC7QP5vDrmsF0vs8/BfsPXP1sZhV
TlwWSjhm0W6BM1UclZx+baL+yq93YFI5SmtDwz3NKe/3uIalFu/vU2vgMOJu
6ZqpV8uTJhxLS/LlvH0Lh42vunFjB5el7Fr+DSFQuWnFoqbizQ8C78nHMrlW
BDYO2oiEr4e+k+kI8GOnQU8n6iEP/obWmaCFYcQBqFiUeuQd7O+iTMgdYaYY
knmdtUhC7yZp5lVSlgYn2yIfzuvlSipvLiANcZy7t+GFu920ZCDxX2yNHi8h
qh2t2O4ocQ4NtufVQQNcsAqS1pbHcJ8nEouqRCC/AEWsGyp6vNYfK6SLmI2Q
vQCkzEj8Fjyj2fedqQf6zbO4Jt/eLvsYoKB+fJvo1vcUqcL0M8ey/JrS8Tpa
3BzCE/rUeqfsnTtGIC0taI/cyGFGYBGCRcE5rPSi8lFxrhy91m2SGArIWIqK
VKYDRUu+iy+SEdcwE73lbaDx1wuHTy14Q9doXYp47bKRnf+I0jsUS6VtfSH1
gaXlDiyk5vN7xShE/bzN2+IYpS0tYw17yzO2wl/hBcBedswPz3xBDNZMx7hM
ONg/fhM8RQtVTYviL+/ZU6BE8N7KblE+FngFOeVsDklzBqXdgpGh5U9/AS9A
k/bg7h6UyLyNkjzgSjd26dFfdaXE0o/CQslX8L3cGaAkvOaaJxfJI8qF9rtX
t3ODVryzYqDneUhApCLPlkzCUesNCw9U9fcYSVOkOMraOH9F0gl6Y6++0/0u
yrXUygGdR91gtm657Rxp+iA0JT8z/YtNbiZReZtxo34JUnpcY5kFwiSisHUM
i6DsObksyvn/ZosocYStB8/ixdInCD6JSST6S2toJ0f5tI2cZAsfM9k3fpb6
yp5dVfYkyeiq7KpRZPSO+1Ti7X6EiXz7bb1fuvJOFm9lv3k1GuYV4/PgUiyf
S4WQD3LpBzJVp2kuflYob4zHFHzqVr9y1G2m+dOHX3V7qq6M2l7BIszveQ7I
nMonN/0pSr0bCnHnOIF/pf3WdYvakmSrbqabc+BnrjKwnjx8SO8/T0iBBGB3
jldedl2lF0Sexa75+UvvDhI+HpamhI9Dh8YywcSFL39/fM3lv5skczzyDNre
+beiytsmYCu/kU9+Viwz5hgftSUe8E+HKHps+3ej/Qk9ITq9h+RntHZRx7KD
UfMw4KBFVOcXC+QSJmOU4llQAftI1J4LyaWmtKim1B+e6tn7vKAy1zP6U+55
6xLHLlV1AMsRWhuQlSC2b6sKLHlkIlRnR9gZdoBZws3ivHdSFjMuCUdhjYa+
96vARZ7grwugYpvVsvTqvJuLxm2dqZXLjXkll3Psmk8Xir6754nPhfGw3cHS
/D6kmXGvOLLihgi+gJvbDPJ8zsQgsCS5BMHZSwidN8ixd/NhkvZ1nM2CJpnS
6Ml2hzEoVksNxxA0yLCyXNw0eX04XO9DedAFMi1ksIkrBK+3mnqycmM24KrP
rd+JXI3Z7a21Z8U5T0zdB3AOHzkClKyGsQxHpAIEMYrKiYvDftxGc17Tvv6M
xnWcNEGdghQdgyRzP+Gd+YhYRRmHRY2JHgIzVT4xAERzgJySIXWCCi7QFVHV
9JJu/8khYUzkficsvQY0u2Lf8FGtlASSiQnNvXq5PYQ7A9tEF5PtQHMgsPw2
FED2bfIEWiYQH3ATgHVb7wT5o83S+yykIVCZiaKQ3tT3r/naE9BmBlrnvX2J
onezonh+QiNi/Vh4IPAix76nkium69/WZbiFfMIe0qlczEJ42pDEGdJiTbc9
RBgQFOstiQ3t6BQtgJX5UT6NOP45y7ssa3Z8beTTFd1MLGtlOQs6wRC425tN
8C7Yw4p2DQNF3+G4hqldA36eMj/jiL2BXj3j+43NIiTYFR6hWTyDHTV7Vly8
yIBKX0N455q5I/NEP8KLZ3Qw6e+CzfkePUqm0uBjvkBcTDMgTehy7Oz9SGTC
GPlG8EIYc5ZBW6Q72FRgafcbL26xyE1WySlc7Bb8UGxoMmtyiUQEQcULMTGo
yVMR4ZiuQQtitisKQg2F1sUQNnFSdRowzYlQwOzQhP0CyQi7v66uTJUuFL2y
fwIike7fwnuxur5o0q9/kJcVw3ohL6k+FjpNAh6PwDsU5XEE/AFwi+h34u9O
G8rdCQvZ51/juX2eYGXmNVUMUhtdz6m8lEGMCClFhHOuiXov6top/3sWHPH5
iDxpjR+M5JorzRRzYfl6MWjxYv+p/893HXLegOG0zJbDEKDbqTeqTgkLo0uw
lBwA2fsmzXQrHdXy638Fa3x7SgQf3Pw4D7SSCSpOVut1nHiXbA01mptR5g6S
aHQP6+pk8oeEymkneYhSkxFCv8qZR2pE0lpF+lBnvvQxDt/bPKB/8cAnncvl
PZMISSV6ryCLmJcNVVHklM5RCC9IYMzLIBr3uGK7gGFJZfuQN/iGiEzDtrhc
4ccvzAgGSa0UHW5rLTjJxhI9pbPwaRg60vT2ZZLPH2PfSRpPJRzfvRhhaEvX
fS5yAquXP8WZGuRYQw5rkWGbrfv7O4nmTpnEf+JZk0k5H7ToWhPTLoweAK6f
UfJteniVpd/zU5uCWosAIL/gVe/I0dKPZ0twL3kyIxS/Q8iaza1XxLPD+Uzq
uSf7x0HiW17WTyDCSySocH6Ivaoz4fXNt8K4NXrGMwzkjR8xB/luR2QJNbi7
iMpvq+N0B/fovykfJ1BhSJWCUb3pwRCuaHcLZiWhW6Ow2Q0CV98gWUVGd6OJ
r87VZ3KmIbgODlNyLsoYg5YGQ4iNYW+OMrfLCFs3BFl8+4XUFX3XEXJDBEM6
s/5oRPpO2be21t958IqxZpROATKfGmVwjJTfRfkvbeXkSrHodjcGKpDuz4Jf
A1HSMQGh1SwV0bjlVk3uF7klXWAV86FCPXcCM05Z3bAy/wz5bk+5rX7//UzD
hOX4QyK3ApHOzNPeXXr2pzjES08dZkkjbGiEG76A04+1QX03FL3X41jTuhzs
yW6SQU0eXULZfXilU7IDiYsh+pJ8hYRmVrlQn6GXEK3Hrc0EeacOV/6qpY5u
65fGJsSNn0+/KNDV6Oyix3jfWz2fqELvnlPH2ovZSfbRtfZzqbuCbv1abaZO
QLMuW7XSV12/pXMqkAXqa+00MwpMlEEKeQrhPq2EdkdMZ9vKTxXo+W6rOBdc
FGsOcHFpbV3l0An74SJtjUnKVg1GaWgCyJrhvmzYTIKL0Vv/8TbQThYYcuwi
MUZWxmFaaGkQeu8KKSYoKUrYXz+QGDLoNPYIT+X+kcQdva9t1i/UQUWL5aeI
iXwYcWHm7AO/1sVZ6v6yTlNuwcvZ9jDFSHNvnSJof43JT2o5bNB7Dr0V2xrT
Y6dwhlqI3mq8EGh3oPfNNh0baSGAPbHlHKNbPBVD3IcvC34kcv0yR4ZAAIB6
v4M+EKMVc2itWnEqAw0ckTXi/jK0satSNhVbGblxTRkBbZo1jYvsPbJy3A+j
r1X7jTXX6lueCMPXFZTtjobI7nlth7x9CSFYDG5uB3AuzWVQXaAQYs741rO3
Ww2wIAPBEMO+hjHlSTCb7w+SjK0aGV1b0rUPlAqSIls+as/bi+cNqRwlZTC4
9w09RO2hTW+yOuQVTkdSXr0aFPMkCpHJlWYIU1zGPldl8zqvSUGWRRmwxMvd
HHhZlsg1R52wE8anXs9xt7Hs8zl6WwCAI6r/QtlhZyo4dtnFare9do5+6vzi
ncjuxL1eo/oNOMcdQNSpS28Dvqib6EV5JcL8pkXuHWOjHfojYO+kjWpI2CP8
pkCOuOHwswHs/UXI2XVw+iNdNNBdCUP/yL6jPB2GJyMryoFi72DXJy7PuRBU
w2K3RxI+PgwdNxF+QRsD+W0tJrBYszR5b72O6SLA0IUAyqMFTlC0LAGtXkw6
vYoI/TzTMKkuGydB2XqbvmEJxgFR+iMIzsL+3coZir7dHZYe2IHZsMmCBn+1
ge6LxQxaDcMBlZjbQpilyoeWbZyY40tQoMGWw471Y2ko4MCehVUlP9tDk6dP
MVPfFD8OkkPdg1aUMNwiyVIL0qFvksocajz/j0s8Z9WONAXiZP8gQVYLfaOC
vGNZjsPei2vqCrjXiJpUvc531gat6WUe3RND2xWrh8PNJQS9bZ1BlQR2wZNp
tYIXn798IqDyX1bGw/IyvLK98q7kJ9VeR67Rt7wgaqGPtJ97JUzUCm4Nq+Lk
9y/3SQWnared2XxNbEA8MVBbm3OLJIatk1VYylGkdamYJg6yo6yOtzqoj7Bi
gEGmEb+87TbjoW0EyhPXj+Gox2UJJZgbn0VRGWHbHHicR5C5sYRbwlURoWai
3AOors70qTOvX1MkcKj/VD1/lWwb4/SCcL6J7wHd3RRIpat/BJW7eA6RdsBB
Oc6IuerRAZ0FrpNX/e+PTPL+PL80pl27DK8/ZDscsBYF3mL9Ry9lJbNmsREH
7Ckjq9STOySELdXIwu/tr+8w6CwDIf40rQDLcLepoJ0THaPpGWTBQPyW36k+
xJ5ytpXZ6TMa/+1KHYtDFajGXGTuq2P2JK88MeiLgoN/s5g/GGfK71nbvF3p
8Ld/e9+ICzwYQffP1OIxgaQdt2D+ve+pMtbnlyS9Z8BC9uMYIRyquFo5ZwOF
kwYqBftsWbf7TumVNreTUdjn4TDlcUA1zJXsPQ3EJ4/TZHUKeJr/hGswVMo2
1wmpXjtpp3zmQHLqXWKC39MSQE+4PBQFvkd1gIXC9ADUxY+V9vRN2qTOYZ01
3HHxEkwPZV3EYhcps8jSmiLfmIffQcxIM/cAGKb0TxuH6ZCXL82XtlzziLnG
qGLV/NCepn0s0T3d5JcbE7+6Cs2ZCblp7TvRR0UZVDNWzxYYqp+tKN1zS494
5nrMMSwiF7V8g5YmkePOeyCw+GSOmyJG702/d0RagD4Zp2C3oY5t2czFuVwI
2JngMvQnFtoQkdHIb9w+0AGg8YxS1WHJSSXCLsPvF+fE8k1RPiaLsgUWJKdQ
nKiYuBor6WoKqqjQMOyj5MaqSHaXzIDwqEggQT2YtMioDTo2y0NxKfcN8WtK
KcWv/QQT7uHSThQNv9PrkyYcPHK97gKfXhLV6eNzX60+oTNncAuOmBaMQ6q8
CHKWXcOpkz1ZTggqP7yhAtQjSHhPduvFLFbSdf20xgw4Aoabd4xkVgbqQIVz
qyBBD4kuZcX84RpjVoSH9/1vELmqZR02AMvhb7IdppfMolKQx0bcYjK1zggM
U0BNxO/Pwusk64Yhc5DSwIIn6RfPOqWMaULl156Akom6YSDDNDXokcyUc1/6
XThcOL23hadWgrRGOHY0OddFNZIR1hD5GuRfN7N+tJCLvPOIv8jEkK6hzpU6
9XQOUrICIW4izAydzKiSPuSA8tuwXT7kt1XU0Iw8dtCnTU3A06I17mtPWEbl
zvQxas7YnB459Wa7/rDzLe/Zh7r2IZeyjQgtMKoyA8OseJRVQzL+l6HiuaIr
8xil+g1LHvuI2IbiX5PhREFrXVi+hkQH3IePZhtjx+uMa/fJeU/UFT8zI+Jt
rjg0IpamNtxlQy6r84n8e4HhtBoCSwud03ao0e46pL11mDDpY+rCIzxeX/8Q
WPIcq09pQMP6cttybEbKePWrTIOJn09p/0DvsWGrRbRyGZrgJZ+VgOVAYUzW
PqBM9NnG/El5FRNlYxgsDLr5ZXlzNlwEQ6KUIpgdzwOldaSkby6wuLNUE/9M
ZqHhKNabC5E0LBOruv9t7K/xYHp+6LBt9T5Tde4PKxV7Em5Yd9r0z0X0F5IC
FxW803XbYIya/OUWcWn8ZcmGqiGX5dzTH4mOVgzXx3KbgLWkY9qVPDD54VkX
p4sSSTr9d5FS2FXtjEKpVFu7dtcLj3xReml0P2aKiE3TL6pFvmzd2hzDDfAi
Z2RKpl5dGWDmC0R0cAuvbAUr8XeeuCAvUfvDwAO0pDphs2Ccy0GppFGbnubD
iafG3U7Yr5zIf/IJacsCar9QAVbsJAlJJK6dig7Ve2Wuvh/a4VgINI724lxs
vVKtRkCsrJ9fWO2BJ+olsaLxGBFCO+jvU942rFbNsJLzyR9o+rd/fDPrtV4V
1bPA1Y2gJtwwbT0IxsSGNUz/WXLyf4EA4q2/z9ztOnLbvT58CGaoNmFzDBXB
dwjQGBaQz2VbIUH/MNgL21ez+NxAvitwoG7F+ilJ4Dg83qFVhFXIn/GRmmLN
mpvwLrjyYnhaxaM1MptGBae1l7lfa/TY+UmAOa7cIIOTjeR+fK4x/JNubXhl
K4JXr0+LLI33hrvYf7BbWJuBAPFkIq/2F+UoUipaTID6JQxN6UYNf37D+XRz
rf5hctweVxs2aU0B41A9/fVFbguGKj+s0bayPPuRRnyCr/BoaDnOfIOCVhxa
NZLpqk8YVyn6fzxyKTDP/q5Toe48wS/a3L+L7WP9mWmxD8+zsf5gy6UKGzJj
ZNF0vkTIXP8yH4YOTpktTbGY219G5hFoffM/GAlmW1iWWT2X2xKgxFrcA/o9
TUHxByRrzbiKCsvfLd1YbQGrodSAKEH4M7sXJvIbWDtYgUzd7OIeWZChL4OV
5CpUIvAb7jzU29LRuveZ27pOAoP3rYVhbbJj1/wYfsB62ZKcKo7BpqBmk4Zg
A3ZJ9QaXOKjoJ8docqWF6qjMNoouhjZSe3wkCjk5RAMv52R/SGuiOdIu87ld
5KGGnYy3EYXAC4hJw07llY8YjO9TmSrKL62ps4dvXYz6DgBZLobk3wWRH5ED
Dso2w+TcXuusKTqxEzhLb8KK7sDNhitysZkElJIF3fRk8OoJK1TuIE2JHRRI
D+CbiiXYLVjsKDruM+ZMT51U/M7iIJVz9YpqzbLkQ7UCytAb7k15RIClxWnq
QKTXvFLoQeE8L1m7OCIa0iOFgJpFJZXe+GIawd9x9Pn+YoqYVoa7tscvH2y1
LmP4LprDW5ekYsqndJcPJfzP3PJo+owRYcE9M+kDq2wpzxtKzTUlW7rCHQDU
tBmA0O83zHIdXXXzfF1mXFPrvDU9Afld286v7wOjP0ux8BmTwPLQQkUefnB4
Gp1DDt0MxO29NEkB5hkWQX/J7wKhSFBIqs+2IQC0WJGPJquAzRr3tRacNaTc
6zmUIHqwN6qmRfdlmOzIQ+EozBY1OFbN6ecHr2s1D50Y+CoTo5EWmS5+6oQA
GVoGTso1xt99odnWv2wyPXIY+zkLBVKSw2vF0whEomIcUvHM9C2rXpNpNhyW
BtJ+S5HpvAP36oDnN/EGT6DFx4RyhSia1A0deXkpOP9dMuemkSTvBwYufM3H
2AQblUyWylFmaYZYiSqF2halxZ/WzuVHB2d1pUJTv+r04xrA5IhJYB7aHS8x
w35wh8ZGrNLh4lK3SMsKBe6XP+BJUQbED79Pd3RGKag4F8Og6vEpU/bvUNVe
z7gpxJaP8fghGuo9EUBMx9aptDq5r+vHdcfx8TSsDpWkUr/8z5sZs8ST9D1t
GgDYfq28wKYBoPb58uZjlAMA9WpL/ILHUKYiUAxDS5ZXw/2CKzeIX6cESgPE
iKbx1IikX0x4ECuDW7QR61zazzgxnJzrfQbbZaPh3fcSJo5TuYJdW2CZfrSV
MzK+Ax3euxgC/0xh0YZBWDPDOKKXP5dwSVv/S4oxWEU4jm91QcOKFaSsYCk4
vYvNz4lD4RqQK+IavWqphGd69CejWJral/Y8sQ1W/Wlli7PAOeVmWp7cUSFM
1WrEHE2mP+eWPVwQYQeyWTEUn3f5A+mhO/Y0pwETJwQ2GG+k8oi9GpjQAEs0
OdnrEx82auZQBmq9vAblzsAp+15HCabC8uPi0YiizRxeVQDd9S11nXCZ+8Vm
p8X+DLT36D1NlDsZFigKzzwehbewqr3LvWhCIMFyHToWkLSCPj6R3ydBMLFU
mXK2Qv5g92eLMtQ/+mWkSEMGYW0yOssJsl+D+9AOyeCerkHDOjZ7VubP0olC
tWj8q8+Efn8Oju5VmaSRJrPbENnNyEOzCH7RMsiiAo3a+uLOA5S0VZONUbZ9
l6Y+QIvW0IJ00rZC2DCpzP4fpFWGRKLX4bFadWkBMAHNwRxDPed9IaGs+PiY
MUk84OFbbUwGQ1dufv42FqCuHuyP6FQNWdWLa6NQwlauorAmG8x1XV/RG7lH
2oON7EcD1hdhsIIRjmzAr4zuxdTyKjMZVdJUSJ79Tu+4BIN1K/SlgpjWyC0K
5BYlO6K8DcjeeM7jajKcvcU2FxmLTzpqmSVaGqwlhfRLm7uhn3holsS2TLrE
OcU6BC3rmjmZo8eWeO4bKiMn5NOA1ISmLHgkIXHC8PEuc8ou190z3fV7huOv
UZta0VQqlhrDB3whiVR0HXtXRVcWxbJ6/nmGd5p3B2bfDyZD0VkWs6mB6muQ
BP1qyMapeAyjUi7KydpetywRHWEE48lBIgaunzkyMuE5KrFBA1H52qEeuE9y
pZdJJhwMHw2yQiHmKqEuJwqMhQHWLzFGSYzVGdQjMT6m1Tw0wYyMmSezWPgG
EE8pX8zrke2q0qAbVWBuUZxt/GmIBmkMyL6tWI+Vqo5TPQoKJHYXYFjNAEdf
zRH/g/w5zOrz6MHK+uX1l8faYmq890r7nw3VGX8stMJ2qVdvzJtcz/lqYLLF
6OHN7jkJcUv5S63PgOVH2pD+xdYN08N6Zx2T0ZlkHypCUFKW6G5e/qFpztpA
WvRfCYXEcZLdpUkXvzT+uOGxaZad43InX22cMLqhAjIM/ppCW+ci8lkE1+2z
UiIIyGDQWl5CxQywhVTRloOg179hbtLY6ktqMY5E9KDLUDvyy8gRhgwnxVz/
rYL1KSpccCJqR9EX2a7QEPoCr0fvYaTQH2gApRJ3xhwK1WpNslLiPkVTTorq
r8nvwgTTFVApoVGWJnprndgkElEiFQLkK7bflgUn8zcY4wrbQwvqvPn/wXq7
DmVHAGUkCK50yQySgxdzEkHrzEADkdETFCzWK6PXrm+BGzRDVflUMBWWOFjL
C2jFSoTBOaUSXgNbjUGAqvsO7HujCg1taEUIcrfqmRP7wOl0ux8CnCSoFz7n
eYDewXpO0tG6yciAm48K3sHFgVPk9rDLC6oCbwIwcMF7tvb8Xjf2eXVy6l/h
Arpn1f2dncnv0Jvz9HiXhKLhnJ4qyt+TZztV74L3uFWsHqVWD3WzHnz5vUMQ
6KZBFZIMCh07ViJDchihXeiSHgl5BKloth9liB5dhVecLcquegAthzd4s5MO
rI3hnDySfeREoAx/0TnoSmPCc0xom36VgA/bpjHttVgXobYbgG+eZeQci2dl
x4lMAwFNGRhIMZP1omQzfNTmn6DjGXf/B1Yb1w2T/oqvO5ZwSS1ZNVJs5GWg
3x3ld99Ttc7jtmVsJg2AJL5Nzuv1Sd+Rwz3D9LhLuWK3puTak3AntZJKBGVt
HGtPyDuKNstUM/+ZKZjOWIGMya3cqsUvNW+IDQlHkidj2PMPP88Cvq6kF4Y3
VXC95O3EP1BFT/tzr/w/giSJy1pNZii/E/KlycfuHDfZimZW7GQKyUpQ36fO
2GZ706G6wkLecbMEP/DYe42TZmXlKtmd8FBLIEJouCnoM1q6ixGJMwlHuepx
eQojD/JtGl6qfLUFszywGCCSRBWZ5SVz3tr6ryduvrzOirQYuOv5tIt8SpFK
9BLLrJL0XAcMF6WDoBbOEVE6UZXYJRbvKTAUuIdZHV6igAU5RAKQkXDG9eup
qWVJiauOtrg/60GODRMLZUjrTx+Xn9Yl98wdEC11Aa61D4V3ticCdeYwEYur
AWbfhGpRM8VyeZlNPjEKWXX6FX4HazW+OoiFXZfOLim0OqhMeMCcxlXmeiC0
4+WER0Xg4pJpRpDTERl3G5X3zoaRc70tRm+c30poarQbYQj8hLNuZ/GrEC5H
vqKdTl+jYFmiqw9qz5ErWMt8A2U5zWL212AdGYd+n90Hl2Mz3ZZKW+1dhqPa
nbcBRfVMgIldvy6QooqiCt0kM8dgCz0wq1SlHgQXJbZ6HGtqkiLPSTib3mBz
/ZCThgas6ayG9UB65NHzk9y5RVFI4joB0osZR4X7IX+AfdF8WNP3oGDXAe5z
aAY1ZhgmaPqGcT8VhyGP5sS3TCZwzIHQEEdKhrg85+b5ZbxmZdHrB6Oxa2d8
iRLZT46dmePHZlTm93lhx+yW+sd50vFmijcivU4Xevjwvu15AD5byrzXHgJ5
0wK96hZ5Ebujs/dwTSqSBc+f97I0N33UKVb86Wqpjf7Eqw8Cn4ZjlFUMmXiJ
D7zjwQkR3hMIgIJzcaE3iVMgYrMPkttHrCI5uhuT9eo1D3atgGWqLW6vyTXm
EHVLNTfZpKK/F1u4U7j6cU0lWD8ks4TURVz44jYf9vElIJ9bhtxbhUpSjW22
1HncXRvvaewkdR9KjjcKZmgdX4Rpqv+arefhLfcj2er30G5DR/hHv5+VLmAB
of5TZlhhW/wwntRZFJNMwSB9ACuIWkQVLQrIaz7OT73nco7KFV/rD2EjD6zu
Pkt/nIam1kcvw4JVgAhXDO4UKpdOoKJjHpwJItazEhuNBeKAwYSAs39JMeJl
a4i9kTEdfLBS0+l1l2S02xKBiDI8eP+XzWfux48JAM6GgmKnG5D7McEmRNb5
cVBlKL4TtgK7CDCWb057gVxxOAoDpnFfNoKfEtiLglh02CrCtQJ+XBqICOce
Zx6m/dY8nt5R1WStduRQEBW2SoIqQOeyaSCqH8CDD6QN+e+z5sCOHB5MBWmW
8pzAJ+Adm07G6h/p+gJ0BYV/k+TbNbsgA/AVU9VXAjIY0KFvdwaQI1Fb6Bpg
z7BzVfCRZeMQ5Hsm31lf6pk4r33okJysWJLkaLB17f16iYSbq39lqslBnMS1
Gai5Jqvke3SCR/lrxuWn7LSDVm1I2QV582Rb1CeqnOPH4PW0hfV0C8of0bQC
grPeCd7HvwGuV2e50bYvNXyq6fAg0Tvh+Ba57TMx6d3We3eO6zN2A5DJNuFk
5G0dN9q09vmJ6H2jiH/Iehw4AtDRJ+4nww79ENvzNlISVFmK+1OfOIHX1FUI
HTau5ehyhIBLw7P+htwO+wDxjY7c74mIBhQ2xGerImF58Kn+YP5lkr/EdE1r
t1V01y9RHqyHvyoZn32DLKXNETB6AnLNSFGu7URgLp2LAlUrOaj4SxvmtlFf
qTvMZfav1RRKugKL4Aw1by35Ev21x/tddUVsI6+oK485Tl96zgIXHLrlpNIW
dMxqouIRi0B+jhQFu4BGglHn0hpiKubRPyLN+l0LCKg5WiLrtuYw2e8rhLj3
GUUcw4L6YTPktuSLNPRf9HO8wz8JQfkk8shc/aK5Quo5YvcKkOCDkNTivy/5
ZIwSxW8WV0MV3azoZp1p9DdIwpi2e4eUSZ4dLza1kMOJVjL1qlj2IO1HPV74
PGRlVujfs1dpR4CNfm3Kyj+QxARupeh72XkPzMmJP+UEjwwtQFE/ZXDKeEk9
tijKGOLq7N9xpLIrHxoaJIFswiEVg+6UQ2JMJX0V6Uc/OiIcw1cCBO6I3raZ
bEh0aGlGfUEhm245UqKF32LuFiiPnL0rOir8RZWEzApMorbV/sQFXfoTMnD7
bt7Zey3FBoB//hNtbuk39Ek5VkpNBIpNM3OJbbKQV87+pbNKqBMumH99IIfF
8dKOr33WJdJpak+1b3QqbjvsRCA37F1EOpGltxNGfPNtzZyA22EKMqAlakFU
UxMIEym3aDhOfId7+tON1X3NpuOtcOVIaaXrlC1amxNPWsLaw//6HTbnn7RS
nMsm8CGlaiDdjti/uQubuTSB2AGiIM1OrsACafg9aZ827pVGH3j+50LcLUhn
OLzgs+BePTDDXdNnzffW1lV5KscOSD82/B/zMhRliJJpYBIXnkVoTqglHh7R
OjTFO+whf+RwY3eLnZ8KEGDenF6/UtUD7yTcccBGAzRtnM+8ysSBhIHk/sCq
Czi35tr4/vxtHJGCdkl+N+sl8HDUWQGABRJJFRVTCg+K9encXYjNurHR4rxd
oA+Vd11z3HrfgoUEDluLhz3twSWel9Kv55oSmjgVr+MoLlq7ChiobklsUrtY
lPqcFTyy2owfS65pMFGpotIq7BKRyCkxqM0bHm+p3C7XApH77cYKJIg1np10
dHL13HOWrDXvInHEYAHeIAQ+dahtbIMxmTcMDeU7CQaTUhQl301gO1nFPmqo
zAuuAGT+gIFVz1gF3qPaQ2bE//YQsFe/dkx+JIf11ajxIb8cVQS3khrTZl1a
HqukNwTdJTh+YIfQ/GthZNEDqlX5bvbByoOAMXFtkGM4sKEPPdNTDXOHGlK/
fCpArUW1OK6nyJiulyHDSFtJVfYR6burShkZdtN7/srLPw7zaMXDahumuNQ8
hizrif/6RnQR0k3CmRr7zdlkpbJvH6XqdjjUGwuvXUCdHV6yhGk2zCVeezPi
SkMTqncM1+/7+9s6x6q8Fq28Q0w8rau3+33nd5mIVGO0Eatlty8ncAKeCJb/
ToU0rwLDZTqRJfPB4ZuI3FdcbuI780F3pbY5X3jpvMYm2/ia4fl7L6yvY4FU
hzY2ea5x0O87c/XBjfpag9dsW1CE9dyggTnEihjbPt5B62kZQdGqeKx6H0Gj
I3yeKgsHN0r9FJScy6lpRWB7EmoAfuYOs5J0DWhnF9O0q22oHNmtFeqUbADZ
4Aa+HhGLN5iR1x9BeklK/6gZFxSI6am31g3CmhFuYSgmSpIZikiY+szj9/ET
s5qULogKSCC9iDdvJcNFqXc8cLr+582g5Nn+zLSHMoARR9eDva+L/LvB93Kb
7XBHmDnnKk35AjiXKEdvqEwJ3yTXB9eXTJc6NsxI9WjAhmrIyWRfw2sQIgNQ
REgmCsTs2JBonn/53BBG5ZtDuReezLSaNUFVm3DyrPGJjUTBxsKitav/m6Tq
1HJ/iYEWWhGET9aQCaXV9NgikZxTQyjWwdNjN4gbeADifepKClt0E6lVTh9K
wdY7DuhusiebWUpgxyTKALfN8eEk9i2JsbPkeasR/sBSd8NLes8NTItLZ2ht
DqBCv/3HHmQcSOIT0bG4lO8+Nh7ZezO2c0kufQ+JmuCTZPlDCAR8IG4Ornjg
29zFrUR1W+5wFR1otNFQWyv4Au/lbdnB5TPwQmEmD1DvFhoYdGMR6FXaE37J
aIv8b1CbqNSNfRoq/pO9og0c/vPt1GVaRePUInafKkFzNTkziATQ00tqeh90
H0Tt4eZsqVGdrswsg6gs43E2geWxFJb4ztqQc3CSyJCBIav+als0Pw7jPh1m
Qhc1J6527WTqt7nHzmPbIx7IU/mAqCErA4IXUxdJRZAVZ8F8cSQ4sdy0w+65
hRswGNjGEGg0wOH3jEGttL3rQJYf9rfD6lBrpIbGlc0vqNRWmzv2ytrskOnl
Pn9NjZqRi58i7uafc8tkRAKJ4M6F/B37hYmV+uowY/nMlXng9MnPOEUOrl4u
6hgZTT4/trdQB7r4AhoSG8XTDPPI90yahLL8NnSrOCkR9abeHcaGRbp06pU0
jH/F8GB979FlMIXjYEMnljpoXao0WvzwQF8CpfJdVNT10AS8J/Ra7jQJS5ms
HnapRPPlKtJJ96SgGxIE3XCvv88iyEXatvaPf17ygHJIfAonjHGfTBzdjKys
IwAaNgU3iANPq4hbJWrOBi0UjfxHE8JUGiCQkP/NO6pvAgGdmtR+qOthfvn6
vIzankJU2W8KHrD8xw6GJWuLzO20DRGDgbi/JmqLEuOWh28ZO+BrOte/Qqnr
AXDOlydUrji2GPy/A0hesiJfYodEW0bGTfZaTD54imhoiFlwBMXr42c5B4Oj
9rxe2oUG2poDBxfFUhRTUFqhJtu8Q9La2y59p/rSLe8y5xxXEON2yjlfUGLp
EFUmBFFNq7wllbZvUvXRArcjtzHj+6RFwui5obDHjCF+/owDGeNwfNKHWS6N
OGyg892XilQGmU2+Kar5LGF21hJm595IsKOF/yNKl/JJSzVHxYXbzHGLijWS
2QlO/vedyOM6KjHHRYXRt3vB9TXW7ke6t9keHwQgF+z8RlPuGheYfv5xX1ph
6Q0mV+UY6xVtMCf0exG6IsyNtsdYjH9Sbt1XvUD07fYZ8WbTR7DcNpNrJ83W
4uEnwjaMk4WqhQuEGLucI37SjRdiaIsosH7jeYAGz60hvZqE/G41inCZ2Gha
c/H7td26umxLfgK5L5hD9Arfru9X9IccwAseadyCkpBUVmXoiZ1/mKXJER0X
DX9Fr88fe/aNN1nFOxnrda6Jg0mEoFCVu5PIjpR58h6VobDwdjqVvGu4fFf3
mVn0brssJ0QE6bdVkepSfXngU9ReAJhEfykzZ51bssot5vbBKX68reDnWysj
NPNrwmz/7CLPE0c2SKbfKuz++LbT1d5BzIaJJ+ISJY4BzLrhEwtl/1I2NOyS
83Cxu8RQQbwUJ77mL6t3ggD2hFcqC4/6kaAQD7Mx1TVyv3fyUOXT9xBxVtxR
12sm5IhTwyf1zdcOikJCQ1/LRp4G2HxSPYlPVm9RiuFSSd0Szrec3EatUGqi
1ZqCpH2didX5fWZtJmao+RVI19toLdvpDh1lHENJlW8yXBwOorshGymCIt7V
KAQwZSEPPb9xZR/XAuKogMV79jY3sMivfHo5zxbon54vnZT7AvJ8rQBca4Lc
63/DJQjqAjzIGPRRWAn4X74Ixk4dt8MxndjvxpQ+Ux2hSvF6rOI34EVw7sEb
7fEawdOMDSaYiS6vSC5cZS4tauIg8N0J38mA2K9VGWqpSeIrgfpQyjCKrh02
pHqwDjo3IoTt2PIX9PPUL4MeSctiko6aTAJthNvuo5JcWP5hEbtEvep3aw+7
aTCM0dptra8DDSVnTU50r2Jc5S/QcsDDNXQrXJ0zdMCUDXPSAWDI1bFSb0iK
PoQisJSsOTHlACbxBtLGbemI2l9Z0I77taUqdOfxCl50+R0Cqra2VxWktpjW
E7ud87rV2AY5RvIVdlkxcaBOm+P4iT2zR2pIL0DKZMbHnOjUaLepuZCluCds
Nsm2ow6ep0JiUw8YPI3xX/4cIdRJC4+nvwml+RiUejdqaFrnAHGUjb7kSG/o
bh/uK24wJ3IqHfZKefwYCfVbI+6qsexvmwUQRt73bCGrw+GBWeTkxqvn4LHs
1fUFhzWyF6P7x9En06neoD9q1k9PLVrKBglku6sRkDehdvgfsyWQV1RBxeJH
+zjIlBfUOo+HU0IufxHgtaQB1tMcEYt9A0bxUmaRLLW8i2hyCOukC2KKmOZL
+E+aiemGoVsjx1K8v6rU4FNSKL0WCi2bnqTj+qiezpM+LgzNfxKsrHM4BxU9
fgMqvks5FAY6FuWFw0uDo/O8NR3IEdjA6pe1s58NiWT1AWj1jRil+/QQCwyw
w6iJtXJolvtGwwolwg1ovg8LQjSHn5oec08kI2xHwh0+lq7i/8J273GUUyq3
QJu65Bdjyo/dW4hdOit9Vzq8aAwGlGLqs5/YYs1lZFHq9YM/4N2ZceltiCLX
vm7+D0ZN1Eka29ojJkgTDM6t1VuTx2cT/A3ys8cnI5vZInLzd+YartdCCCoG
e1jE05Lexb0/mWHCvFo+hmUkNBga+JsxkRFQ1i6VyD6ai4ANK8MNzqHnOYJi
l4vYyli38WeZVg3hm993LZpXVnrJrgzoVa1N1uvtE7LLa8STurKA2sWyQ3y1
F/7ibmgz7fIzuAzuw1ONKOTiLaz1QILTuVrkfLd3U9TKkHwV4DTD+ChmPKeu
VkEkGsvOC1R++QvOhQnu3ncv3pXg38SRoaUQ40WvsX2EOP2AX8mNp8ADijbd
0vqx8L1K95ediLM53uEAbjJSnLF0TRX1TQvwBynFoZ+DI3Bm7FPMbY8wC5rw
5vDTJt9zKWjs6knF1+t0ujEpyTb9wcdkyIjhyE2v5mre6IaIhsjxN3GHp7Vf
8W9QDWHDdqOtWUGbQIHSWzPZBPYzWCRHp4xGGtDu1SaVjM7O2LPIAcGJyiYz
qALXRV8N2SaBhDSw72cfX2Fpk7BpEf/rpW32OgqaWdX+G6TYlEv9MpEJJSaO
taKtmrl6BpE8Gk3y/E8A83q0aYkJ2NptDMnud+Jk3sOg/PLzKAmFOlbq76CM
oFQhFAI08ArOn99298PNzyVuuQ7ATdRlgJn6EZyxnWEhF8eEoIT7QEJMLQJT
iTvb2+upXzeHiKrRJ8o5DqaCY4R1hwLISqE1mMV4YY/976uLUaxcli7HwbD4
BlH5tH/Wai9rV+I0tnn+pEO9OU9+gQVzWisFT6or+XYyG8qK9eNOIojt3U8k
O7owwSuh+D/t+LqQgsdcGcSLw4XVfGn7kbiYFAmaZyW+tK5A/3NphNKtOMwp
f3O63PlryN5sQ80hbGmLXqgM7EBuBSVMPjRYzVUahh2QD9TcrMMThrLxS4qj
TYoXWZ0jZUIdXxmw0irJccy2mxweMaGCxveQ/exnzFk028QAaN6EDgX9G3Px
96h1LPVISyPdNtu6+2ms5GhKLgpCVUmSaXujOhdCn43FGP3s8IPOezMTY6fs
OBbqCcsUEr6WRex1TsJOX5TBGpK1BItwjJsn5tGXVdRzuvyTI2l3pLxv99bO
rGdkvPvVAWZ1C2vBVYiXKfcEJXU729arhD6CTc5edXxBYz0Y4R8Y9GsbsIzZ
vEilqsjcrxR87yOumfF+jJe8N59qF1ahscs5uJMzUJjaRBDr31aMWLtyVCQy
h3IkIpn4mhGi1KKtWIzdLfcMoDjcVSkqsgaEJCvF6gBlqqgrj87BEFXIl2/Z
NrXa/F0QuhHLaC7BBlT6thwCKh08tfg7dqoOmx64tST6iU557yUmBa3xdNmr
wwYoXMON4xj2stMmG93UcmKKuldt9nC1BQX7DLAv4XP99SJjajn8FMYTCfYt
gJ7YQVjrY7zRPgUow2ErTVpgJ7Q/Cc+lUUx3r6vjX0mrEtWBSiy+bA+Fm4SR
MmCjezwYrnbrw77rNuSOYb8MPiLStzNb4UDb7+zxLBZDWdMNGfKqXEuZFOzr
SZChfeT6EfnnPSsp8DuQRPg5q4UiZ7zMPbLhYzkxU7vBOEzrfaNmmuqxzMI/
foalmvk28WC3eu5enM9CxAVje3iDOf5fU/VwZKtqn26JHtyC1rK9eCalpqID
RGxAdayePtt6fTgRqIZT52/HDTIKtpd0TWXjvDkmEF3MTvOF7t35I14M87cR
BOFmEScqTFlS1d/nmqspV+e5gWq0NP4uo7Li2zv2GJD6qvteVOFCu3k37de0
0Yi8+z1VFIsE3otn2dfXhMnyJMMg8jO/mkOwxbZ9WEdGSA+x+Jc7Krstku6w
qyiFyJHLH2ex8Kldew9T6PZFVkTVziqNM9Nq5txfm/BqdjyiOPM863lvApg9
VBt6A/t8j1zPdgknDi6BcNZoenqH77U9xFxQFDR8ItPTI8MR3dmLc/LBzLBW
wb+KE2LTE5jX9fWyEK7ZQI+XMeGpwlUZOdx6acBGg69qFdXUZ+doILPJNDDo
mw2d80nFRiGQHDv9Ty5uYCRdE1gXcCXbXTYR43yB9PHPGnzeDL6OhxnaGBs5
XWQVvQbzscT9mIQhfcTRlKub/ySsZg2QTEaaMMJKU+2x7LdEKqe5rFpKA7Mg
VyW+QsZ8DOKZhWuCQfeXKO5/Mf7oihlIH+Tkn+W0/u1VizjZT/W2kzMrtDbr
9ViUaGwiXvWZlRkAQLQ9T0twyPrHgMzZPOjbr+TKkn2Po15uH3Qy5CquKb3N
H8wne5XMIJNXBnz/qhOjVcqZ5eXckw84S3UEY7C35NeX0mwwCxk8TJ8IELpU
Nc0MsXN+gAxNClmpyCCkG2DsSBq9ktIVtE0FW5w2OKB3D2NX89/9Gmg+TAtf
/RDI6q++J53xgTUgZHJ26X2AWWeOBAEHLhOd+S0F9kl1Vi7Sq2CAKEQ3+pHi
JfIoR2LX3Jwhg60+cbos22Uwm8XM4lMveNzC3yGEy1sj+C9iYmm5MBAaiwVw
jDQ6BgU+Vj+bwPb2eo3aJeImWu7txJw8lcLuP1+MDwpY4nyVnNus2d9u2vx1
ZpTUYJYwB0H8RLPtMopEwvue5XgziSevAbsgWSIl5ovTpIO1N1H34N3+Sgv6
GnAIRMUCIvy27Ks7kzdfhqbxXiGdCnLxsqOXSH8+wPdNeV8g/tC4pXJUHWh0
uANi56mk2N4VeJePoJ2S5kazH+ZlMVYKTi+AYFUY7DV8CcbIDrLXAeJtyTrM
adIJjxmj4ZHwlMHRljvbX0Gi1g446+QJqKx0oYtLSms1a5fH4CVurlSIuVLE
/HiqF/Zt/HatEMNuvSNh6bpXwS5NPPnHAZ29kdY5dcCRyXbTXgvt9CcNf5ak
Rrt/tTtXhtuD56Zvox+7Od6qMHNP9hT4mQWduOd9wKi6nG9aMd2+CIO1hLpX
Vgy2iHm9VAKRiwV1EbyMhbHVmRrO0LwAQz5QHc367CE33qfY4wEsmv4gaB7W
VbMD2M6md0fqQyqglX7ZHbIQJ7YluEN2w2wUQdMFEeSiTBvoTUujUTEOHT5h
uDb7TuJ02WjpRkJSjPYrPJx++WJOET6+GtDg2WEMqVuhbApPLDFdvX5tPDSi
Hm1GAtUnu8k89lT4l3hCwS8IWoruvQqcS2/bk1a5091WaeEsykZrQ/y0gKLW
NwPilUpC//LSmC9FTMr9juwGtWsZVWeRQYeWYrGMNidMwaCabbaDXKRHREYL
kMKW5nScUmtB12UBTrL1WqU53yA6Vn1a54lUM5HIL7znF0YsRKOJeSRCZ5oy
vUT+nS+E4uIxkbPkwD821kgBaPGmQW3L9wmlscHsyVCT+Shdg5w25nWBqh/n
dZMzhd6qR6zMDsHeCsXgjOC/jFcz3vvP8nCwqOyR3kwU04ap8MqCoCR2P99A
pRG3RXaR3eWNZNVjiN1+4QeaT5bhMvaT9BRmkpyBKQ+dOuvikdgT32gQI3fh
rHj4FSLGGKqTVMxUZR48g1iI/ITSG0hJciAWKY669Hpjiq2M2eDiO2Uym5+U
TiRPFZqc2+x24edRwLQhamO9zHZAAOYXIY0UFZYFl/hb4+uwlddiJvNFSYwd
9fZVQhbnpT9s4Be9qfET+bkPlw368etg1kJNcnd37690ocEfkdUp80Nv1tc1
hCSsQKzZoPymrFLS20MPLM9rIha7KFBrDZQexYHDRxOS3n3i4hvCFqHQZE+M
Ps3wskUTmqyavZnuRoXQPx0M2f7pfN3hgcb3qogjXQ9v7rON3EcAKAbsAcLX
7ia3EGpYH/ZHFMlk61IaaNeUSHUVpS89IzPRlsklj3IMQeuPN+4vBa11u3qQ
YI558sfnvWxJ5R8BvvWuXErG3M2/yXUPcdHi/EFxMsx5g+KlefdI5hUxA12i
lhQmteTaeRo+v+El4z0r/IXKmqOmz4JI7HrnZKofmTS0P6s+VX1oOq0tLJt3
kkhUiIzbgv3KRyHP2PRc6+4p1e3QXrm9oFRTHthKZkkZ1Fd97A7/a0YFG5zj
IVkVlv4CxNCBP6mI3dc8klno9q1Z8n3O43quUNI+6P+U/wPu40haTvdcap2m
GA7Owf3LviwgqXKQ0CGf/M1eggRGUXvFwb3QV3yJJFoKEwFULJoHFqRwFPJV
tyMM1wnDCC8y9yseCqMoeD0K5XhvNnkWIpeC8k2tfpoT40F/ODoYuBQUe7hL
vxOyxQqtcmlHvOx7Qho7JTmaErWOp+Ffnmu/zyQU3MBZBhZfGOlsprR7nzLV
2CHvhAepR+BzjJDJJX4FnZZAKuO/03QsGLINuhSJ6epEQ46hrLViKo77kuXw
bNCQBpzhxyOG+U0RRiQVbySdGEBp6XmagkoxbnakpgqpmdaNIF4OKNXk71aE
cQjHk9wWv+eneKdOo6TdKFRA3unAUM5VEIPCYuWCKKPm4wM7N5YEB77opGyD
i8Uz55VRZLwsykFA/gSKS1UAb4dFv+SGEOvbIBtClpywDmGuKffDPtNXZTeD
k6wj/xY+b4tEcrTElkGG2zMQAUwPGy8RJWb07QElr326xOJIujaJVPYQWPyP
TZN376t2RyhXWZ4ORMkiPWbHUhTwU0YgVQcLUSCbAH2QZeVAhr3IGro6c53a
pW0DN4mfF/RKKbUkqLm2dVVycglZB6fxq+DpzmZvXN34+BqEjMVflEe4ssc0
DelosVdXyG02NK/4p4ntDv7GyYhkAODsv+6P65YOl0AD0TyC8IvvYORypGc7
mlsbDwAN2inc+qxcLKiH0fxM/VE0+1vexORuAiVjl7aZr8SpVKm35tP2MrJ6
9jeIAvA/SWK90EphtAftee5ioM2leMYabZurvFytT/BWOzNDA17BDkv+uCNE
ziMMnymARplKoDHTpCeKVczMxKWYuYLHyuM+FDVlbTQiOFR8Kjg8QIW88qMk
mHxIpTzMMo588LVzP62Pzy99/Uaym9aS7Azk7Ncys32TyjyWjTV+K6is1vqd
0DdAvSKmicpYE2ejItW4BgShcGWE6Kgk6GV6q9ttOOg1BG/0y6+0Cq24iRSx
uYVOpc9bIyGo4pr+0KHUxRH3pvSQ9pPHvRwooncwd0uH+A/HDbMRMTWeuZB2
my//HNhQWb0kB9DxBhN0MtoesAK9c2b7ebiPZ54YxFUHLWctL2bXsnKJ3AII
WBInLLjosepKERNGYa/ZSEEI0jx/ywlDMQ7fbjq+ghiKBSoBhzig81vIzqjH
AIlbSxQhwOmJLbmlhsvDxaxkZfIhfpfQqGF5lfZFWEwne39O+Wrw25GB55jx
mc4AyDkTJfTsgay+l2kF42ZJfGIC1fVcDazkrXz/Md0V6mCUjxf7DSgLSk6a
sdygI7DsyK6j0I/4H/ME+5CP0mzxsqJi+yxuh7wVnR9YsDcmI9W+Cy9TgZY6
RQ4uk7t1Pom+jQF6ScJxA8+Zuv+4k677DMv5c9/B/5Sc9N+JMzCcXnYb3GFE
bm98Fpi/lxaqyp/GUCO+JSnQE0IKJNH2qZohLeV703io2dmczT145bFT4ZJM
YJ4sQ7KqTTR6ZglF7eAhbOl/JcTxNdQVoWE3Ep3ZdNUQ9Iljt6L7ZVfkLil5
abx3zHCs1kLtjUMeeY9cKBH3PmZJvb97EWsfRE85J4PyxdyAyXVfgcuzm3rp
hJ1tt0vqlVvLSwXKUU90+cvq0lB606VIKHcT8P7GZTAz/axwfHNVMEieR45u
mBRk4vx/yptG99GYC9Fh0XzBksUB4JECwsTx6zrim5nAAM7xmDanTjGM44VQ
jJTJheSQ5ypKM0ut34auELeExFlu6k8sU+GT7CDVHbcmxK2laI3rYkDyabWr
G62ghYH9360nUfDsHK9awmtlp3djeXf5qCItrL05/uzHidwXmFeHeFHaaadP
aUkLvb/MmygvCceCvesPDDWNP/1zxYtRpS7X2ahtbcMTjMdgmg+aprXT3gLK
KKkIFrsM1nvfgW2MP2ZhkCGECZkb/UOzp/R2wma7EX9bQDF8/Sf3ptvKOFCH
xzc91cPH6r4qV8EL4JbIv/tfgqn8viYCDtETJe+NU2VzBtQsplgTU5lhxmr5
qynv2mI5bL/Y3nqJCT/GVc9+sZKk+8j+eMspZLmwYs95s60otHFcw2MZk4GZ
Pe/atS63L7gxRxuUU+9xqxV84BBJB5+lcFy3P1DC2IZexi45EeqL5BebcYvW
EoZxxD52NXNiXB23dnIPapW3Iwm3OD/IxhCxIRjKDzSaXy341ApGGu77evR0
Zonfsv+5z2RcWliXZdf0bu0ROYPXAAB1X5mY4Obz8ZH4q0uIQOVxbDIXQrli
iz/Ejcfh6ClQ+JWmXPYwaFPZ3Cumm5J1qVDgeI6HJCyXL+sQrJ+H2uEvC9Um
yCpjrWfw3DnC83JykFJRdsI54QY0wJKTpQ2s7LDivPT5QPpbW0Ag6XTe2o0C
PyHLR/KCwJwPXglb/IHSQWLl+z4AxYyQepGm3pJCsPwY+uzinyRlfSlDqmsj
R4X2jlzwNIZFyT4UuzerY4MrG/ZqwjYTfjy6/Yjp/Lb9H9MHrbNQ0KqG7hoi
eOoPOxGVKFUECXlOON6it16JqWVu4xEIgAM2hWx70++3JhLaaqbDtFFnVXva
14YfjGsD+rI8JAIKZf5hRNWYs4l49Pq5a4byvqAN8b2nuhUI4Kg9JWnQ1Fq1
VJXjRu81DEMZlVsFUNGBK9KOJJ314GfuZiPz1CThWcAn0v+3CXnAVp83d9kj
hfSWgcuARj2jjrajidmF/JnQsBhkxk2CVJe6WpMDPK9j27m6ajo7fj1GBqHK
p1qz+KmoFivq8Z1cqQCyf8kAB6IvG6Eji6geLABaW6V2pBJB1XyKPTaGuLxz
iEw5evkhwYwgPQSlZm7o9kYK6Cduiqps8XfNTC8PzCk009f8ImNeYynKRoRw
fT3cbPSOoHNhY3v9+naKOx+6Uckm34/37RFXtFqfj7tFj6/M/osbrfjA10Lu
3l+1Wi6WRxv2Rpr63QBdDKZFrveY6g0q3LgrkmFl6JXLFuoPaSNV3/s9y/GW
yPITcXXVqBs4+fplrJJ5L7i1plEQCosuxiBCjlQNOxesuDXEbo6QwYr4VxkK
Bochz1tCQFLyg0l/Pl+NJ2CquxKJB78OEj8+kzZtcW/Yys3zezJd+ywiifN5
pEW1g7c45VTKWGowgdNO0npXlFeioQ0w07eO9VECNNQ5WsgYHKGtuFXqsseo
UO2Wxhhj+inkFrFrh5qqL7f6YK6Ij41LRhfF5kcFkQoWPQY5sCT+hXFwFZw/
KkBrPEDg0lTD9J4ETmk1CKiOLM2L6X2UU3dEYAnyOzfe7D5RVyEzlXLBAqx7
J9zN5wF5V3q7jfGXW1L4jqdJ3OEujivsY/RxUa/rcPBFroIyGLDb1T94shBS
EPKm1btARHxs9ea0waBojOFzT/sEPFqDpvt5haU9SknXcH39v6b0W+uOSclc
FnNk5dizEkOQDYMxcv2s+Zl8GTYL1SVcmDG0NAX5uHvb4atQXn1AfVnusCs3
SK2GwlLf6A/jgxttYCMMV+eHjmiJRba8s8wAoAgzx+rc7hI3LgymqVc/TzTu
LGkNDeTDhTu/9ip/xCl09QBc5JWTrK2kvl1YBoG9leYaKci4F5GFzHS/waKc
ATg9SKpwRG1B8G0ogSsbwIV+u0i/xtRpeK5PxOgEq9O4qMPaJfCAiBbvyYeo
HgKimiyCOWP2NBafZ681Te/3OdpVT7Syj1DNAtHA0YGTHFS69d3SJN9j69g3
jEGSXmVZ6IVFtgwyQ2Yqv87u69kb0eAEG8W4VuLEEBt94y+/QvwtJ3YyV1Vx
MCkqdWIwh5wenkbsIsL2SXUs+0rtK/1KQ00CfcS5VHzwbdEI/TnQgxqewWmB
vlHhxGa/7o5PYer2u/Andvi8WDp57PJdqYxUu6zxewYNkT8XIWrKaYF17S87
Uhg3eFHq99jK80reGzdmmyr3uzS9syu95Vwhecn0KwMcxiGgEJ9FYyYRB02W
5wmwRTKBYlWYikPYpI4gyclLeq0qcn70rQw9gZjofreEhxHTFnln/Xi7cHA4
YvzN/bquSqwk3C+GaI5eNJOoFaqyU6VxzjiswK99Y5p11S9xFDJy+QXAq2pQ
BVfziq7uNZNvSGb3NAhxLm3TETz7J/eeE0nmP3CJBIgQPb1WteK7uFedlDxQ
2W57rnKm7cAeHtEjNIh6+lYeblatcXgrotwVc4lyxoeFuAmST4iA03TcFFiI
sgzVQ2L0VI7SW6NyptBakGScgnyd5sVwWrc7eDHrggEuYah1OmUiLMmkzdYw
SOcG3CvhmS0sdEo5E74keU35mnI0NzrFu6A2NBNwx2R1JZIk0+x7zmRBDDfZ
tqs/a6F/KqQR2ggzVAat/p9Ff6P1VX5PXDfbMlXpcjuymRHoVhBXJcoJ7RsT
E+t+89a4zP/G0rsmhUxMEqDI0DUYBoxuYF68bekI4Mqjfg81vCI8LsJwfnzD
WR57ZgVWUySTFMTI5earAzRI1jsJRNT+XVh6Ky1XCRd2Qu32lCwdU1D1E3bn
cGhQ/mBtJdFrXykco8o7pFvpFh0jXfy9zNK4ZYIgWORXX0KD6Mw7K9MvIxgm
qojqyLW9nbRNzE/sUQUv7BmwvJzoBeofB/p1nPWX/Yv4bBsRckxLZ2pA1CJe
I8s7wA4JdK3f/v38CAeGyJzvMmauH55KBRLIOY3zaT38AiLcojEXsBOl/gbL
yggcVr2KmKG2MEsY4Ii8MWJzpznNTyzK4QRe6s6UZkIDp6jVrv3K2PImQ/3c
n22hDUMHEqHS4/aSI+VfT3sxO5U/nxVTogAWLokDZ4dLhCp9aYIiH4hvDkYv
55uF9gyRUB077CAJT/KkGvipSxLTFINcZxBtRbp08Q+RSzacf9Par7qecbId
r/ZVYpSek2R1zTuwQupTQKKN0BNZKVuCKzu2Ipej/FpTIWNz8hDxyExaBJIe
8KVDVANh+uJVVWRkmjNAqDJVJs3ElmBS3AJ876xXe0Sv1H73/Fs60ZmDuryc
al1mleRyZiNZPu0WzRNEQACD1AQWjyitRoZmf7ob5KV5cICcQodgnTu9JbHy
fogtoiU9k9vjI2yWXMPs7P6kmtrlEUTYWOmLHXSSvCIw1fwc2NpvINdZA97h
2rUFIb/GjisAdP1mUT1StyQ0/G1/nMjDOb0BEXayYBfcJeBdSRC2i+3HhSQP
ZRpIpq9oEuQO9XXMDR4puYIoPdKl7gmPnO3KJZMCtBK+EwWuQcTBNa5caZMD
6FpLtuAJauDWrGGDPUINlIgAt54AxnUwyiIYdIts0eYE84hUo4pONneXyoxh
xWZVDbjTsczu/MzYbD6WNbHib3OGHzq9PPLkFFSCBFeWeEps86J3s5ur5qRY
rL1YCwS3/qNOtZmgm9A6zHsr17LgNW1w1vKchsB0R6B68D+iq/GWMGno/mbY
0PF0IsoPkt5D3kH/nv4dnkoY2zEOe8AL+rHn5BizZ+2V89sMrlG7Mzpe02b4
Pj6iUQJyvdhuN1OT2ml8wP09aXCU0tMYYB9G9BvMaF3GzWQ/eG1SYLNWlJWD
85JgCGwdETDPuG4Ned+4LvCa1ql6K0Hv3vwAXpkVJRf4J105S3v6CCffw11Q
DC0pKKUp+5Gp340u/hC+Hs80fppvmaSz5DN3xx4YJqlmH+iNs5uLFK3iBrKu
85bV8VfErGxNk38NCtJ8yIlqhFoouRSZtkKrrs+RkibLJPyKKm3UYe/J7mGt
NpfXKJm0pwH/QneJYTbC96KJOJZW8Mb/3TNgbZataiYMZ2dtD//txE4J1nRE
IHRPYIuLZxzAnlMU8/5/fyuMwaN4IcKYRsU1Vh0zOXDfdA6MIAJnOvKHwiCk
BC78dXFXEkjGyhVXWZ99MiuBO0QIYXcO2WcPgH8ZPFPxzgMi1gZI2RUsqQ35
g2BMaRNBHWllzjHD7jQSfqD4bqsd+dYZuDljY/OPDsIVOl9NJthriLM5Ib+V
wn/PCf43D9LsMyqUUPFyVmOrvtc4veUor85k0eH74AwK3of+hYTqn9yOpu3L
VOjwCvUIBjXUpw+4Htu5OpkryEykfe45a8bNF1sOM0qO/o2490tNo7aoF8Hu
zUY656oMmqGH/3nS1OD645ywtrZnaRTBd3qk0TOuPYM1+AngTLZZjCbANoea
k4zmhtrO0citN0HkJuGZ8tdyYX0oyzdD0nA4qJKGk0jJy/Can4+01P8s98vv
2ev+Pg0yzHOeINOMu5ASHxsYmu9Oh1mrGMefAR2iFMPdV+uiemHlsrHYzp1O
7cJN6QtTr/bMC0N1Up2+v8QOxA72vZQUYrU7NGeBKwdSN0RaH7JWU8WZwbSE
Zn/RMTfZX1FfoYG5hoP2ugF/I5yHjTJ0+omGtL0XGa7n8EwX3dKeXls/Vbdl
6hpO9G5QA0EABZl9Du5qHeDI7x7aCuj9p2cubI1/0G4eSwXupWFW1t0piqUG
5cb9npeKD0q6hUKD3TONTbehKvTf34CuWyfr1LVGdAPNrx1cMYns0bGaqvRT
3uQ5xeQZEJnsd93anPqR0/BYEWf/ebOpOldj50RpZUDukhq92o15mQ3Y2NOe
+XCJv8G54J0L9d6Hzdg3jH8vN2R3G6/ejQouGcLTWIbbaUvVDsEeAsEdxzkk
oLdIg81YxUKlT7ri/dG5NUetIzdUS9SMrA0UuteQEuPI1CEY0ZoXL4zdNntq
O7CJkS86HRbwtU5rzA2Atmu4JrRwb8Ee7zEzlJHSFKIVOmpQ9m96mhP0OUQz
GqYlAx1KI6witQjx7SECeH+l/DBxqQtogUQXETf37WXQHc2qfm4TBiN0EwDW
4LZHwEGdbAmkCRF0y6n/6Pqq/PIP2VGPrO/PA/xwKX4ZkzJiGAG8H+4LxhnW
QIq5sN1qdCZMc54RYMXP5YhNA+PX2ZpqmyYMNXqgPvSIQByHDJ8dAqykvZ1a
SkHnRzkwsHF/joJHdtNHhcUvRkjJCAFqs8kytPiE5ysRb4c6wBVg62+rxDzJ
QmxirlfAdNLpczzm2uIZ5yBVwuV0JItAFMjRDs2yynC7iDPk7Nn91NatrCpx
xXaC2+f81cRjCR2Az/m1XIDVTnXTTSrkcHDssHijIqUe3IeFC/MvW5SJ3wiO
R3fgsawUb3NUM0bvkV8mvxvfPLsPbuBXhhEP5CRzrAfmxw6jnqKNMXn/HE24
h4NJkGD2ba/uG1NVdX0gYamJPz3LDkx8SrucPM6Njqhj2eEzYxDqOX+PAv2Z
/312NQgAjPrzucqTnk1ozoJyQurG+nGquCNpQglobGREP8efV+bo1Sw2kwVb
SvDriwkcFZzgwsCvqPPoHnpcTJMEWeBwKoR7f74gvDvEgZnTwl0kby47RugA
z+PnB3H4fSqnMU3hhfA0ilPuw6cKfZVXYQFooguYx8HdzmhTsgTyl3Na1NCz
7mb6VrTzpknxLXBrHbLd3JAOqbZTY514MeFEWI4Aqp3gje4P83vSz13sXzMm
qRVFnEX5VoRmx06zGYeLEolIiZMrDiL1+hYk/bc+NUXHccFMm15+HfXUVAwP
WZcx7m3LPM54C2Wu4H2l0IhHRcraLKvQiJDxN6a7pHkUIQVIyEo7s1+MFpt4
zGMmuTGN038QiVGtJej7CJtKzAJxsFRfpqM79hBEk73r7enEIESQVOuJzgqq
kpjDK5V3QSwberyF5wH/l8bIyEireOkDQhXPnohOfANz3p+7Mo4Jxk78JRrv
L1MhUOIGLRmVfpC468LJv7DcYUu4vST/bQqbJ9b29EalWWCTCTuS08s2Fpm6
xOm56QVjiGKUIvil1XO87pmaUbdYVFznNA8Ixuxj2dru1X135kxvUU8RzmZa
FDCAIsBtA8U1gKwOGIVUV8W5AlYPMCtEUobA0Fiy4HhiBkBdjb5QTNYCF6Lo
x5s4VwH9kgoNy0CpsQMH23FTur73yJBXe8DRid4OYxJgzds3tV2DzeuW1BXa
oVTqCeNLoVqgFWItc5h4OXzR7wHE08GO0cwUZLqSEd1MEuJ/LBjOQ4KPN2vE
UNbIG7YhIFB/GKtWP7F7DyH8rX/yEmBYeurgyOHliWrvD8RQHU0UdCqwm3at
K3cWuQjVmegTwHTlOFyrHNyT06MrKwyPkoF3LPjDjuoSSnezujxYU+2WiH1i
7oPh1Z6nakv+PWhrFpMpShOWjJ2thHrexVRU4jecSjdgBNWFOAGAhB0XNzFD
93IIHc4xzOAS2L1d/QGb5uZUP0NvXsqvlSzcI7g3vMcCx8AAaWXUVdijRaru
6A+MXhimpcook+Mo4xt8bhNVOoxTGviLPh8Zu1AjbNVw3rMlrE9VG6IEKNal
z376cUANpgKicCkluRCgQLeN10PpdS02nsohdWLh/7GQAZk9Q7MgdPoY4pMO
BQCnYQsfNHl9O/NTUyUyb1VefawJaIfwbcW8slk5YJ8iVFu7uEnTqCdx5WCB
3iptOnOw75+Uf+HgW7i9VYtEKYvaJDcdPXqo2NxVDwo/EC9hGphqir3nn2tt
GpTBmbYKOZv3Btx9vQXguZ0RK0lMtbsuxhJEeUP0kYCXnKA5nMMADAtav7UG
NhVOPfsN2EsMr4a7fLOk+eAXvtk8fzM9Ykwhigyu1+rq26Up5Wwka5adAL5Z
sSK8FORQw/xkZua3D0CzbOYyuKXvVS9heoQWVTjmwMHPWTTVXCBHK1JVQxyM
GOZcM2L4+5ZAU8iq8HLEkCerrVjAFkxNIjCJVQQVPHk2gicRJgv9f67pVRzo
9aOHwqHPBMZiacga+hRFWgdcOIWoPJmd0z/KuKmRLBdOLGiLbCpbYAvdSEEy
TCwPXvG1gHNzpU2ptu6l+VmD7/mIg+1E9AS5CW8dbn7UPgwaCa88xPpB99Bu
Y7HwgHhiInX6ycSnIOa89uG51fr1v67ECZpf98Aby7ab269My3FREzr2zpLr
UslayjOvPuy8Xj11UlIKa7ru4IjA7+WZnciBzV/RDfh460xpV7+5/avordvS
KZDs8eTbJWyW3HNWwz+bL16Zy1gh2vBVg9geQYzDbdyQwYsnyG6p1YBT51og
A+VFdVHlA0bUPMw1sykdG9cGygarRa4LLXRkSEdvkV9TGjVplaV18jIjZjiL
49Hvl/X9l2j1ZwKK7pxMB3TPtDvSBiltZyM0vD/4l3Q61V3lN7WhbNLxESQN
g+o3MsUHdxPo8tc0kNZ17H/TIzPm7tygomuPKQ/gGNOwISBsq/L9M67KQfIp
62rdQIS3M9xXxezjHReHzfWxanvpyvt6f6/zqudEkJ3apDZFx2c1ILefTjEH
7KvrPtCAVACyCdX3gkbCELIzCmqlv89G5PAoouhvewTwQJqNcYm5ql47sTD5
WGiRKKp14l67onXd6foPTXKyVDdUFLcRhsylJaWGoxeAd607noUenS+cLOk3
PMQlQhgQtom+/vTlCGa7zbIO0sqFfyMU+SwT9nflKmrpPQd3blDtABqaNN92
lB0vRpY7G/fiAsKPyPN4bScy1WRkVEJQIOX3RnhjEAxV4KpiRiZLGmmRb4xi
M71XtrZu3F9OqGjuu6hab052G/MhLQdg0cg9hlmT+XS3Tjyi0D+/wpLgyVPe
sCQX/y7a/3D/VY6fv5+5K6/j6g1EyxMNVyQN2u0Uw3HJy0xjyWDsQRQmQE4e
vfwT1fIFGzCOGR1WPHCPKScLOOTLAM47WhC/wEciLJyTjkuha8pwz188jdEk
pzZt0QH8y31UMXLsVJDC1e9LRMNcIq0oUetdfQrnAzHjr9UXeKEnzC5rsuOt
mmg+Qb6A5pfq8iiMXJ6c9MGE+GgHu7/Hm8Gd4dYaawztBvHmuYuVq3BXQqv4
dTRiLRae8ls/EaVHqduHixaMm2qYvieWaPxsxLmrTBUu2f2gG6ObX+rZjXGF
fuVfZmyzHPtBnqSXJ6JcucuwSk5DnMu1kVdWxXr8JySmTFhiwj/PTQjrJZ24
4rWJFYruKnKyWS0DikmedPpecNyv95oLN5c+WSmCbEqW5PyArFRaaN4C1PxE
OLlvmUsTUyBPxEF6/bO7Kzwz+z9acPCD6//NgYi1ZXkAdn1ST5IMGby74UBo
Pups5oLX/xJ0+AM7grNOLDARB/7jy7WPpVG4If4THHpNCayR89E1XGQfK4UJ
HuOU/kZd4dnIUU3fj2LmHYEWxdNalWJcWGHqmeSa7kYbsUu/4ngNG/cclF6L
58x/In4ndxZ7Em5Uhf1cBn6j7Hm4r1eDN4Q1jvHlmkAgXTaQRFEuaAEiy6sK
fBiubECJO5Ux+k0dIiTA5FYQsMESZUsSFGcvY/UXV3Q5QxJSMUL/D+OoBr9N
1bujSu2HSlZFH6udtuDISXu91emA32eErvNsFu1j9Fnm8nIB586E7AG+qx5s
LnOEcsgoYwrAFSjPrVHenQC0y4g9Rb4JkJBoW3ZJ8j/M1yYcAgT5gVdpI6GJ
1XQhHk3jcQHOQZ1uM797BzskUr2D+8NZp/GrZgatgVI7Qe8rj4UH7pJkE7Ms
qJWJikP8QqTAwFQKJp1hk8j79DZj9rEZ8SgKPxzAdHbMPt8srHPBOUY8W4Dt
mO2mBOO2P08PpCsgeMpYnkF5oSb/9E7GVDkjTjsKj8KTAj56KM1jY3YcIiGK
VSou2Srbs87lbWjbBasiq6d8fYNUzXC8ycxCLx9lpLO66uXa66pjJPThO2/r
O3Uta2J7XaRBEZDqyZRWNKZfMXYIFVDdUTj5xcyea/+Zak8/fvzs0rtNmZRv
ubTU2DJXGv6QcjYjUenjl5or//cPPIbTXsCJ631zPmghyIOimUoGBxwh84gf
Kv+Py0hqXeS1RTWep9hINSoEdTFAKhLcMc2Oyvo1TZ7hRd9GNBPPkaeiTkpD
uj3IUFEmNn2kdM+rbOxWoLxtdYVWBnA0hisL1keYcozG5DierECrQ8uXCUY9
YdHmdiGd9POqZOITT5Ed9weuYGdXHQfXuYCT3faJU7J0DvDw0bm3CemulJeu
1Ll3yCHCOnxXMUvC87oVOuVPBlKDcsbb2VDhcgfo8+QxJPZPcMwkw//SOdOu
qEaJUPf/TeScD53FayMey6ufYmeSnm3BA4wvrZUja1iYAKjAKp8OaCeUXUrf
1whEVsjqhtWA0fztbHKuFpsOja+qZJmfW6KFxK59McpiU03QXvvzIRvtAdo3
3XeFebon6+9lS5AEygYc2zMZsVW6C77Q3pigxkWuy/H2QU76iT8YK4GY5rEE
Ures+/rma5Ni8ATktdlh6t9P9HNk21tsM37LNP/LUbMAjXBy2aAwjRJj/2Os
KmP23sZPog1jrsMv2GHacd7EPJ+OtJkt3uPsYkv9slgNb3hThrqmF9q254El
39sQm2VNYrlLTd6gELh4O4OraWu+IayvAFl+ng2avxi7m5PbVmzRPdNge2qo
S5ypgMZVegUc8eAuwZdtwN9lNda5n5nBr9WT1Qr9TB8V3XNGaHvOTZP2uptn
9bRlrHUGc+7Xg/seaS7snOoONwzqNgptrFcnb4U1dNcOJrHsIxxuvmD9k2J7
qeAxpANpIS8NF1g1ODdCOYw7OJGoCSlHxaRUvhH4OdjsAceGr3EqgJgRhwc4
/5dIPksSa4SZTwAxmRDg6as874gQXd8tXfTXUQ9RQwVrVF3ZK4GaBJkczZFd
StNmuDvOgk8qBdX0DcHTCpgC0afFvlbhLmqzTy8mKczecWfqVsdT46C0CcEO
Gsro28p1faqisFk5BVA5tz3JXczSm5XqQDEdXHhCBsa/Jwcnao/0HHFi18EG
tfbHWIlPo5TnRI7i/tb/vULDR++mJMPFDS0ZQqJMPZ1eQ/0CXZ2qH3zVskKt
SU/3AN8GgTjS/XnQV8waC28H4pLq4s/qcFhNAahbXeU69xJppHDxuj2/LBI5
jE+Bca0RIHIkRfbAkv2OhgImL779cz0oSQapEbSs3rguaXiQxIFvO8zgB2Zy
OvaSbc7ejBOY1tAdUmspj69YhyrAH2FdmJy/ppajVBQ1iRjpwhnRMoYyGPAV
Q/aOaQs6+Yd/VKa1weAgwHvnDc9vtAktS1REPhucVSMYxOfgBMHQUZMlITzp
DwmWj/ZBsdiPpN6R/6R4ZYy+gRBeaUgR0Nto5pR4zfBPeoNwRc4t9qSLz2wA
aFV6BcqujQQ9j4wreUn/N1ei433g/CC5lxAw4HcA7sU+5M1ypm7O6B1QGhPT
w0TeqRH4RlVmrsSLxO15J7cICsZzrDN5l4cXw3lWYxk/JiKIsdSPQEbeCrh5
UCoDpHpiKum4kCL4eJy3TmpazxbrEgrpzVLZF347DDcPjxTZB8S0G7HBm6qD
6X95N4yprL8olD45tVs5H2hqq2DdgRsJwV3zWmG+mZllMLHH4mRrsaLmi6S0
sUHiFMRDVE2PyV8es2vrjxxivk39RmDx0vu1eDeRrrap+H72aHf9Gj5IoNFl
+XBRYpKGSRWWpibhJMVETkM6mkFJV9uGYJ+2RNvNl3Q41CLShx7A85Tu+GsG
75ZC+58G3KG48mlUAv+ODnqcJoOV4nt76HoVDqpdCZeR+OWqYUNiX6Z+af41
FpeaG7LV8UF6iSsEj21pPDeBZcV4uKUb3d6yXYPZkoBHnmGGsYRMLL8Yka/q
Ood3YhpXM3ZH3rO43bnZEFvHNrYJGtXpOiReg9tWeC3W8k5J2zts5tGwDvhK
SIHjJZXjiqsMCh6v0lY08hgmsqDRe30xQF9pqYlyGE6FOEiGnimZ8qxCdRXD
7G2CYTkPlFd2IDoe1oqTBHpLrkxgeCS5FdfGQFYSnes1rQ9YrEQu0XhZSt09
hSS7NGQVwXlCfKxZ5rO++c2RB6phVlUZRoAts28dF+CEjJevmXUpfWeV1UDA
8RUZZQzWCXbi9REAdgCS8f6jOSg743iXV7ZJPAbt7upirfvcCHNOJ1jaeruB
xTsfHA9qsm3jLUObbAPkgxZcVbu5DT10h2gHufK1rNQoy43G4ijVtF7htgnx
ZAkvZNpDqFVdNPjhLyaZCTuSmX36YZ44znZhJQZK6T1Wi0UL1djfiKx3GfAw
mqIHGD0eEotpv0dFNfs/dOZxgKDUB7eFktRGADkcgZR7W5bnaIcmRSu1/xfv
atBjhpFoWiYJKsyza0exQzswkB/BM/KgVaBN35DZYaRomYuLSIBMFK9Y5NV9
lwyEBwgPGT67/v61FDfEWE4KZ887JUX+4vcU3o3X8ECO6ZZ7TJnIMrf6PmcZ
MjcC4GRRCPzDqxc4qI6GE570UT7hjy9GVb+bFOelrrJgNBGTvZeScPppNyVT
YgdIJdYLA75nOfWJhVrwriiDAsyADNeGFIG/tfKorus0BxA3JHQJ8YvyryKq
rESZvSu41m/PWQC6UXWcY8ONNtLkV7tUdJl0TzVCmOAI2hAg6W9CXTc0bjuy
hVj9aZ6ThtW8RDn0I/J9oLLpxeT401FbWSyt7meuGfdFPq2CYUPIV2NiBnfd
Hbt+Mwds6TsJNNdWpHjyPDtys0advAP2yZIbynIzEcLqQrDRFis4Ii1X+WyT
bZaNTAQ4RqGmhnMVQUkPF7ms2k2hRt8A3pFGreyAPNGrHOSl5zvwDfrayF3D
4vrfQ96SIcc6LRQ4nYm7O6YNiZ2i1p8/tsE936Lo8kglXvEGkWK2IbfSuZY1
Josj07y3Np92fvahj+vXB3fcSdlqYKCphXg6VnKajMFLA0QYgaUptlWdJrC4
gp7KOd/sippgs7yvyiEuUP1zAOSeDAnzDhVIyDi+j+bpnUHdlSmUqZN5sDSM
SO/FR7cYkZgdjOm96L+4QYLsfl/jNU8A1zLDRSIlfrh0+bLsqFlT7mBTZDaM
RVIxXoopSe0oL5BCy7r5XPAUwwout4NMdIAOWj9otm24njpIIiqIOpT3vhnR
i9NlhdsUvyTeUCn1j3ulq+1ovoMWKrrHRsBQG5/zMoHpPpRDH8bbXFscDNPz
8n0hdOkUAbxK/iPDoumgbukBBXNHvpfZ/PncmjgVYh0CvJEsyfe8Wow0G5R4
dbAvVA/x736jciEqhQizDtw1jyeODB0vdSSVOVreyaSCI5wKA2Mllh5WYcZ0
lo8qFCsxr8bhSureUCoFf70aB/PFYDG8ZXq5lx2MXo1BHdS/5uW/+47Xm1Qu
KKhEqAD6xA+gRvZGhg7YJIuWirv6ggdlyDq10Mz42OOuBE6VYWPphvgqOo3/
2zWG8sWeiVKUy9CX8EU8JvSPWvHyFWqqSgyLxQ9JFUqZkhmZPe0F/ymdPKy8
qZ3+X4ZUHOXfMZ7SJ9nuuv9Nh2JjQb+Wjb9JvMqmJdo4ctzXvmgjesxJ0Ptw
H17N/q6pGXgJpga3pAAZztcsupLvQG/yEsVmfSGo0vYjfQc/5M6bfvrq1wO3
Feg+cgZ+Okqq921RBlr6yY1tBIo2RKAOwJEfLu29yHZGpA3adKHY6ZKkxrGl
wyPMCaGNwJS5AJIr37S8L0PbwYswSZMu36bnuWeKo6oIiT04oznjO5iid+Hj
8EpHS/A1aCJhzwx5DJZRxU7YdsuXtjLLWpnXgYrtme31Ln8lt8SUb7olg4yT
Bj0Pod/uFxbB0DQOQ49osxI1pLV9opIxOULWfkP5JQRIW44VNsvyoP2dTKb6
2t+qUSImPTV6BlDft4OUYdNXEA5uIXGcBOuWCZFYTLQwhodX9l8US8GIeExG
s2HI1JU+fxzePn9PH/43Q8ijMbE5hgeIHzh7zgq7C2xSOiXbP51SPE5YURAb
G9lmWyPi/KpCmvIM05XD+QDnotHDPHn8EM309oBVNUWCGB/baSAD1Y/h/8Wu
kXlLNItVMv7QfsHgMqDt9Lxsi5C85eHyxHU9Eo0X2a/ewfR69sUsQMLzjpLd
63CJLt/a8otxgUXkq6ZlJ7azpe6S3UVUdro7eho5esiIbha+Gif3VYlznFZY
yHcpIclL9O363NgfmQ0b6noAsaCafmbyKutRD9XaPPqCd1/DriJH0HQWunnU
LTtrwX2s9qgxSQgM/vSy3r5bZccEJOPgrb2jX1AXHWnCgBnqd3h88HMD+GEw
QXCq8NpQdJ5umtRP3pzFjlt85Su3cP3oQ760OnxFRxhunWhLns3BgaXG58eE
1YQESW+a0CUxamvdm1/HXeKG+S3i/PF43SfdZWwDu35TAEELTfqs/mLsaPB/
LwcQH3kPJrvUwYbZfgitwWIUVwhmYP/6wuBlVjrmBcbIrmDm9xE7mF9wy+Tk
lOTsZLBFqOda1hlK9j1ZDbg32lbhl/57BAJXcpS1X0M0/oTObDVAni3MsddT
uIjGJQCgHhSd4r5vxjD60d5hywBAqxybn9WPKQxL70BhHO4wr+0e8VwD7Ckj
/IoZRx93I1y+LsfVTPWoX2Ip+xZ8iPg4fJSb+ntgdv+3BIgij1Cas1onXnuI
M3sJaqZKBPfhi0zYE0TvERU44xMqk5Wq2jsqNG4szD4kusa1D9AoJWY4qCAy
biB3Ofq7sDNct96WaM8eIiLkntuAJXV1dcuaSmk7bovMqyV5g/CrgJLHPVPT
SnGkPFzwEhrtSSPfHHSx/MRzWwMEnDF70LM4YCp+ohd8WtB4jB+t5UWLxDzi
vOtdA46QEU4HN2GF4Fx+LQHr/P79YiEhSzOwXKfQGA52M/iJV8OKSf4OjF1t
WyGbYbuy8LTsW+F5p1PvL6VZstNlvrWf/7RS7MvKqWKZSAUtFlQa2dERA+dH
42U2pysb8YFggl1XVS7db6HPTfI+mcdu5r/u3Svs5tW26SKGfeCvk8eIpl2V
XzUp32L7rXZh6LEI4+YBRJVl1aLy+t1WBMNbC7LXGGurQSh8rE3IY2D8saL6
FdC05jB90oAAmrRa5qc1qfSW6MNORhQC9godeE4+zm60ej4Y4WP5bMAygMen
btrlpJbBX13PSWHOfFjmQnBRkVSuQZgxB9ZAlsDPynhfWLDSsUdvX9V0DH+6
wIbbXMWm3G2iGMlHJgM0WzxqtkY4PXF2nib1zVfgc/fgoH7BligTZQ8f2XbE
plwKu6MtwMjclqIlo+97ga61XP7ZNWlKTxHFcJUdqIKSIT0tBu6PPiZU6VSl
fAMGzc+0XwnsDfZJ051QLdEXO8WpWJu7K0VjVHuSciUGRfw3OJ/wosJClNpU
Xc0cAxxP66JnimanJMuu+wd0SNJ6bYwmlxbciJ+frVCKRgYNprqItsWKXmWe
6ueRfZke0cciuc+eROQr5eH5YAy+LoIda5Vie5sCkzWvI7VAkxguELaJqqtW
HXQNELfGsLu4gwpvJkLrXMP1TkKX4Dqlp6rc4L0Qmr8RtX3SW66PVAa+4r66
j6kp2OIUoykEGlXN86oaXR2qFz2y/YhLuTe7gUiAKP8ZHyt/p3wW8pwUAdgO
ZEU8M9+Oba+vvcy+6wN7ScT94peCF+Bnv7GP0OTQI/+8Nv5NqjOpp4rZ+3Be
EP3EqKpS6WxER2TQb1oSinRi9bokL80QgeC9EaLo5/yVIDPWSCVWb4mNWu5j
ldF8bjkxoXjbUmCTU/kJw8VLt6nCJKPcljbdvVxexlKjj4QcBdXWWDaNXU5J
E/ZoCRwIxhp1QQ9n7L1iD3CQsq9kICCGh/PXt0PFwrQYy/c2I2E6cyZAYw8u
dR2a6gMcrRzvgXKOxfqkCMMhomvQTJubXs8Qv+sFgqL3wb91WttD+zvOTJIu
f8Y7u6PRfRDNa/G5wDw+Krx8fjCPobJAXuPVRSEvm0KwC69+Zy43/OaFwSiz
rMY2OcEeziiGgaTjGrO3vXphZmn9uiN+LWd5HLFKgwixoc3l6o9ryFavJP0K
IgcZKVkjx7Wi4zl7Q73iyaT8V6Up2GnFg6kdwxHN5Er42QEp7KsMLxiFnQsc
zjhMMhWkocHHoep594xuxv4BWtwL/M8TUnLGBlEehmOhJiHEBkdGjQhwtSiK
m74vsra8YKGSilOhmPVfXfR1B/KcnxM5qHTjiBzNhbAeALAj8W6BQPg0lSzz
+Wc4+N4NyVZ+aMSlHNAqvcluq+ebP4z2TQaky8aEhrS+YqZDLC1rScJwXq9U
p9Re3uB9Hv0RrxqGXHKeixwA89K6n405ZiCc1WPO4K7olS04Xn0I7B18o25d
SA2JXo4IoCy3oQcz0vU5W66nFazwLI2sDZ66BP9RrL7alAWWQgN2c1hhJTFf
VjUSmkGtZzXjUIFRi38Kz8kATWVqmRhQCnB0XBXYoSnVXZbXO7c0Owdw3Btj
b0Pf6o20sm2K7T2AaVP+H9fPViReAjNNoBSNTFFKgib6nzcFHrqaAUK3DsKx
jEny6pSzoxN+a6qZsMcSi1hD/HS3oBWD1b5uonm9UmijPHifNAQhxU5iJnPA
U7YTVmN0hEMZIGlaQvkoH2GiGRQt8TKD2HpmLOINV3VEm0U8S6dQUbvW81s0
uW2Ab8Da5PXzUXdQWnU46h+QdDhvV/hNRlGPKuztr1kivI7Me0z7EfEIIsoS
/JzU9hbU993t38lLVLdRxpmK2yO3kXiHSkLOKk4+hDhJ0gbxoOwN2MGRo8OD
+1/7oeXg5zyK5+/3EL+Kp6vqWpY5zncf9b2jR/9+R4d0Tnjvu9pQdXRvkKa7
M1qqFBHCgt2E4ovtF6Po0MApEX7JzHZWdfo6kcDfOGkjwIdyc3+qeDAXO5o4
KUwewtquRqR0uxpBnTllCKoHxqJBPFSsKIeS2nxnP9S1yVPekgVCvsUEHFOR
HGJMJQAqw3QaZkvUXXRelik2P/e+r5VXUiiqimq2+88qlQAcxuwxJGicg8X1
kEa0MLCWkAtHz3GYT1+p7vAez55zG3JAAUROgGdyonRR8MZkXqMQ4bm29I9l
SoaZohS6Y0mSBNFKjf7Cjt7HoIghYT5912VfnAXOFd2yn507JeT1nHSSz9FK
qHlofULTOwBFpy5tOeJ+BkvxKHm1mdwbagUAmDqFd/xUN8WQqxU9d9IweNCI
Avpw2VRdlAetAO6B0HHWcDNNhcE8jDpmPvtLenYwhjWFEVyziPI9I/Tujx82
EufbWxA+Fnz6jkSztq4HFZET+RlvnQjxDU1Vivcb7eobMOE3aUTg1YLpJtyc
CvJODmUm7xclC1npLCLuCbe53H7L+FAOFwfyZcLF2FBbRqw8o8sdyqwmcI2d
G0mhXa20RZ0oW7rVA7RG+6yziPoPVse7HK+LNrS+0yyxKqbvy5F3RPP2hEzB
5bNpsVSgs2bmOiT2+3LYipC0jmZk76PRRvwhLCMcuRPvh6Rpld9XL6ZFYH6t
3s25hnlIGmam/NVMuVWLjmQZaz1MiaSDUSsg2k+NwMtvLTrUVzaeDKudhd89
sMwQtmoRmPC8q+ltucYS+ZV8QMdM3M1cSBKbPtmw7E3iJlgOg9ujiv1bZvAQ
UnCnIlKhk3TN73VXMdkykDvVDfdc7ETss7Dy1iV9H8puAJClv5UBbs7Ur5uS
53LUysmJAVTmRViKg7AZpg7+lI1PyStPSrtRnessAujyTsy8eO/RqFLEwKRz
3CuaI6TK8aqLhhESrT7FD1wvaDE8oqTvOuwtfxEcjmVxSBv4+7uxozifZ6hR
qUqJysnIdoxnZwWeehhrnYmpyiPR0b7YF5lFTzaZzshM5uMTL4KrpqGcwZ3w
V3fmbWWFPZ2Fn9438CVEegmM+VZtYDQQeJKa1UMBO6qSE7VuTc5TP5egMVdk
dy7g97+8/QrCy5Gno5zx2br6UnPR+7orcFKW0fCeLNh2RyU7iFy6pq22faav
ft6ciX1aoZolrU7v2YBhDDzt8YWtBif7C8HNa8+2vyYrBryVZfY4rODA3j36
Xw9YmcKc8nG4hXfj39JGQFn/+4A9qs7XZPiqvKbgZUtPVydZcT02392h0K/R
fypGPtqmR/8sx0rQZTv3ykdbA/Xfck+NmTnCn2YXVbsOvzlXdnwiN2gMaQ/x
6JCNbU37WzRX1po917jJNkh1KjGN28b73pvaUyNpxn861kr7Rz5RGLASCUVM
Y7AWwGosr3jzixNo8p/dFnJwmlBtEvDB+4DZ6QTiIN47nqXDrL4UWbhtwhs7
syfJOML3SM18wVBsy3WoyQMawGQuoyMP8qAOI307hWxb4v/km9l0vYvgN6bh
CMpzveWf5b9Vf6nNoSfR88C5gx6Q3WPVJaPUhNAEiY4r5QV3C8kXZkOQTElB
mJsmNGox4a8mqLFzXIS44EU44MURDCF2seAF+j/vGaImHsgPJekAiKMJKYpe
bnm/501qD/t04iL+cNCr2q7fMI2yXtr4HQcMMIhZcKf7FQlWCoiOu08yQkja
rpT5kealRFdiX5C/YX4yrSUY/N3jnVOiLCkMcEAoKHscR8Flq2gzoOrHBsIC
1bJWmmMeEZHnwTIui/z24t/iDx78AZOl+G1+IS1FuXnx4HvGKZs+K/pfqjlK
+RSunz+GVGHxJ3plNF7nCGd5cLOYNGbAkKq7cym0AIJon+GlczY1euYK8TQf
7/wKl+Uwgj+AfMgxsse9Y8IjIi7Zddl1CFwYVlKLQUfyEhIWIh2lFzRkCX5d
jwjMKG82yT8GhSwdOO2CD7ICVlq+VGScxC+w30QSGwvtR5ZpbWJwIxE/lZ5d
DuvEScNk6KAG0LllBHEEKrSyp4csFb+l6aJxk6aWy0+zbsEAUW/EjS32c6v+
G1shbU63oKDwYaEveht+HC9Dngpruy9E1agLO/kEg/5aC21gbt16//4EnOKX
ndZUIV7/qIKVAuIW7dS83XJObWmAkwZZSy5e/HCky4BNU8x1IVDE8KWsBBVP
qtAWdEVdsTQX/GwrcmzzmxAOgkMYDZZHDQUessioyh0wl50C/1xoOzXX6B28
UARntFZwr0z5j3If6Rolc8MYtMH0j+w8PEQI0NR7Rxoxx6i59VmFgTpyvZmc
PDmE472/ZiZZJm463cSQArcDhppr4J/cR1G51F1o0wKQ97DMV32xNhnFoWQd
o+/kq35xkblkA1WX9URLDiPxP1ykfN84X+3ZcTltFAiKQ5NjWBlR8wALir/H
GmQrc8BQP5IDUypDxSJu0Jnl+ljDofpir/FkaN4akqB6BTaZKv8PVb+IMmmm
VSBPOicS4AD+a/fcc6qZ40z7LlsEREu1ubWmKt89++j2BrtjHiHfxXKy3oEJ
Tf9wmcsvq3KnDZt2VJirs0VP/2i7STyz99/mijOmGb2HimFUrWC39YHYqKlm
U2XsdxDtG5ax2inBgfYQcyf95yky/9UTNFo+xdSCPiyge5J1W1EI29jhUN0U
luJeHo/ybd9g/J4xbUUUdyLsIlQevKzuJ8U+JK6Zdhb+lQDj+XzPx+bHBmah
q09NBVXBk0ap8ljh4tyuNCX/+v8X20sO0J5kdssnY/mvqE9aMQLtIkxOpKdN
d3TDe594Q6xmSVmRS2qZy7CPvbB5aumPZp2A4QZEYvb48koG8vXOXNiTyZJS
Bt+7kkxv9BsYCLrkfno30J2xd8WRgyBNd0/i0BScFg0yqNnhku3mk2czORj7
0J+GWvATIjYOWoOIHipONezf5K3enYB11Bwvz4WvHNmW6zSY7vwkXz99pmQM
PY9LuXZXbwjBzibdPEapLAFS8zqKP+Clq9IgUiGyHlrFm6UY3tKJ9lVPFEGD
HOkXUV/av69rBAaYAX347yLxzKxGOaDjpOS+rj8e15opI+INOa4QELwNaAfx
oI36uFz6yJg7+41VJkCtIVb3WgwApPX8qPqAMYFomLL85HwZ8CFH3wcV/SwX
pmHshwbE3LOq7uvH5mevVKwcV9ktV2fuhHft93nYEOItjWjZB/SQlqJincQA
004XCEAHLyFzrGVeVaiAu/td2RbJo9zWGQwV7ruwPtvIScHcoH0TsKokyh7L
3J+uvimRCYjUdVcg58I++ikRNqFmPFvefH7ALQJCZmrDGzMqbNZ6POopaLX/
6ibvUoFC4IPMAu9KmJeuG8dWwL9CRMNoTJCtHZyDBpPK7OcA75T+yXTzY+tq
Qg+1f4kFwpg77NkR7Un5MXW0bkxUDQXV0ipX514HeuHYHM5Qk0ZyMWaxEZUT
Gd+SZ/QsER2Lox1Yr03mQfX84/e7d98BsPfTKA5U0JwfU1Qv76k2xdr1M44G
CCtVvwOmgbUS08w8P985SHcLPDVLfFFgEJfQpkaDujvIQgbjIU5+UWZ/JD0h
6xFYf4EDqpVw2ukg26K4JCeQL8G5vG52aRkT3AT8C4hnYfTL+ClErrSeuBin
Z19Uth9zWBMPhpM4UaePn4irdI4vwWhCLVdfdIFQVNnro+FjH1lFirj2b5X9
H/hOpP0HST2FoLYcrhpon+qgjoaXhesiDUYA9pafuAa9H5e8WIPfgAJx1Uly
g1Y1oNuQMPhPa+odtpQmNMJ53nEghj+IJqueR9vtgfBP03zqybpTEqphua64
elykQZpqgVBFwXNvINGsPfwpxFn7qZsD2mwlfn86zFF1YB/HHTPNriLdY3GK
jEtvQzYwZ1anvMN8QOazCOOztR0BKJ004LXR0fEwE92SCEdQdeod6ETM86cd
qavd3SA5ruJ6kJLHzpl/eZNUJMfavc0hkmyfvs6BfOo+fB3hskViNspos8VU
ILLnj08qVXGmSPHFVDPeosAjSy7LWg2CJ2y2t4LkDn7+o1kd61hCz0gqz2BF
625NGReNNvutp/RyQ107Hj9OUby3AhIhIKMyeHJ7T0YvUC7u7B+fuoywTXcO
q05AY0dM2MqO7WCECxwB7fPKO96i/hCJkdiF0HzpPQiVzREoLRVx8K3AzA0U
UrG4OplKyU2J2TbYJrNzp5kKEcQMTPTWoOuqjhenw4OOdCFUMr0e4DIYt5SA
wwpXlaOif00WOpynzI+xkaC3KzOojuXOHTY7i1f0luG4Lg4OEsKkvosG9IpH
KgHTpX15HCWvJpL7mYQ25SenvCgw6PEWgaujIimQCVKA3cl7L48JLkP7HsFH
U+1kbp5LazG0xsb2OSSE5iJ1sm6lpq3Zh/6mVoKUjmwyWcmnuzlIWcKCdi5u
ixqxOrGU/pguibLX4LIl0iH0j8vrtN9KCes0a/uzNY9X59DD7+oi8USm+urq
IaqbTy9+TxhKX9+sJSrz1Ag17smvVPteD4LD+V8Nmbvv6upGbJIzsogDHNuy
O944OHxXJEq43erVOgwfdI9kmjEA9U38k/9TIhAB6Qj0J3vBxguF71JxTDXK
fZ5YpCrsSX8AUtypj7QIWru0g0fX6Dx3axRcRr9Qf/Ue6ipprWWu0+sSmo9p
PnHKirr4lf48h+mSOL3qx5/skqhXsF/3kTSiJ4P06G12FGJXwIJ82aeOPeRH
6p5/Y+cRO319feXL+i5ED4GCwKjH+/AheaJmnEPramgydP3ZkD3SozHJgcFi
bDoSAZ5p8TjLPDdxyoqc+DXXSgN58WWGTnsbQIW4X/yXpzC21n3hnTeJPaaX
j0yxsSHaDpn6ci6r4RLiqkOb8dkNx6NbGrBFijMpC2oXm0HGv4vYItdwE2Kd
0EkxW4JOtPiAsYi0yZXQUEZX0Rm1w59pC+0EioELuLkustFf2YMXZ2khuxo3
5zsRx/BtNC67Vo06Rf7rpKFtAPP3kVl+Q2IzUu00KILIvxznU+xAQ7UJCzRr
YV+pksykA6+dfO8fLbbuFdUzvdqxkKzVDdux3CH/HBQ7+HdFiS65XIsZhC+0
0sZOURKAiVy3T5Ep2L94svrRT1ssHkRZOiSju0jVZyNWABNIIFr3/JkzCLQm
2VE1YTO9ICYkaeVxe7FQJaAgs1FLQNLVVPkOPT6JACSXb28OkTUKKjoOflmC
YNs03h1MsXNwawqXxZxo1TIGguBydknKUocUnDadfb0dNXmAAJHYWALNwJGH
7cPdky0Q+e5+4MVPiqSrn0d/EaZKmOCKHqNJeWzaqEN+WkZJHf0oXTcCUhoH
AX6ifiXX74dlDyrXwRUK2/8h6KiaSXj+U7Q2Od/PCX52qcd5rZ4CR8ulqqq0
sszW1sgpBx+Dzvi+JMV51o3BXX2gbIuk59q47jQO9qAdDK5wIRIL6NH0dJf7
FUYkHJoacORuqSM02pRXYfWwpXtorNW8gaXSwDrkUWtl24U1GGQWgWLVvbti
nZat/BEg2OXNPCj88P3GofmwFvELjva7iHHHiFOgEMK/DO9FLjuX0qbl508b
1pFryMW14hssf9K1Ty2jqjI50x0Y18Z0+Wsgou/ds3TuFV9MhzPtYSqjEEQV
oYqRgS8iNUVRr5wf0JOEeApU7lbGkqKUVigSrh0VjKoecpELPDEXU/RNtQdU
eDCviAhoQQCQwVA1ISVB+YNWyKThOdSZR8AdjVt1K9hf6e6ZJygFRPlxX33D
/Cr+4U7wB4EdLRkG4MrizS/Ij5Sy0DsyRBEV0Tap1fYdEGnAx+VrBrU2dADz
4yLjq3eJfNHmvzAt+yd+JP935KSKiCKyaLxYhwbP5ukvV+ysyjoT7GdlwVr6
qPXAmPltpRc0UVKmxrWaSJYf0yfF42aAhJh0CT0Dc6ZdAAZvs1qn13gWs72I
f6rgnf1QROqz1HSX/YFmyQrLHK+iNzCdADvrWqQ9xtdT9A4zD76ArSYMIsWO
+tS9rkF5xEjkSJi9O+P+QZXLVyWkcCBIw/oBYB1Rxeaas/OKcRmMQVBPrXFk
M+WB4V1ekrFjWaMI/mKdXWMCAgVujgKukCROcC/uEERo5Ls0OLfgI6On/uXa
6MdypKR7z9i38iAZSFEhtgHs+9B58BpVA3cxHS7bnAb5Kfw0Sm3+uBxHnEIA
RHjJ57Dve77yhrfeuII6evzDWAVsIo6NxFZ4aAxKyjL/Q7TtbcJfuhlviTVw
2vtz+KZvx7k6WF0cSYVKoHOCp7rtqb5CutVr2eHiGbbaKLBVbGk2JnktkFob
W5pCVdgJp51mRQpSjoVhBkoHraTvND8QHhVXmXqQ6kWLESfmedzGbCWbtN/O
p/58TqwO/erjZHPoVbZLr+KRA1XTWCvorJ/Tz+ev8ixTwr6VR65M0dkhjYqk
pntF8CgYqHCfh92IVAPNnnzIHYtAoBvZln2f9Ob2+HHljUZtxEK0t5PnZILh
K7yiuGsor36b6LVGxvIuh+w4k95He8t4MrprHLdxMhqE8PJOBTuZTevSjiPz
1TgpoNkkXjg/TAUvdABjcX3lKHTMJqwwpjEnLC5t08NALwezFK0478k0Hc71
VyOT3f39nk2IJPDkn9lAGPSOLe4ZBmwozZdok2SkkBQnVjwCh07H6edgd8IH
1CG9ErbTsKaIlmgf5gFxvIVDeHR6wQdRB8xR+o09pyneCGbGabC5gtgQcH49
x7m8ZOLxRky05jW0qnroidqK7iCqHeVAKc8bJoaTfp6Jo8OvJCighKLI/Qqi
aAKg2k+9EFap+Tko9UUQ4qhNxgcyQ8hm3yf1H3MO1SGqlV4TXRBTqQjACTTo
TH5Sz51RdFutpJEFX7KblpkJQCiYFL46K1w8BYVt+L4kL6E2eO9XgpIA8yQH
W/8nsvsUiYDAYtHPwZI/zfOxBQAyfxdXxGU2aQEtTjCT7t/5GEzAfzBQHQb0
1becE/OHLpq+EAT2zZLURfhMoeuSFLkRXZcLsVuRuxfrPQEYhOIY4lUnSngl
4eEfurMWqggb2jHUpJtSw75B03nBt8UK61l9BXgOtkNtcrG1+fFjbAtrmp+/
O+dEp6FYMaP+JFGTbzhI+QwMJVECOvk4N9fhzE5WKF1Qx5Y6vUvOWVtpj7tG
XwuKluwY+hs8B5VtC+9x2+pvP6c9u3dmpFe8DRsaokoHlwHsWM3d0ic6R4OY
dgZRe7yGbq/z++6HE7dr4axsoj/cAiMD5FGdJWIWDMevS6M1L+596bzYzIK0
xUshOzk85QOm1hb7pmw0DZpv+V8is0grPjHJbyupSILzkfCuhLofbM/805sd
vrFWnnpj6D9+03DpuftepyPOIpfdaBSFDca0CMQNuR2YFUKfIL/RlnbKANWJ
GjLoG8i5XQmYtXCn7H3Ln3xaU4up5mBIKOVS0uHJKK7ge0vub1Lg10jgQ1hy
ABwBWbTHfpSLF7Nlj/4GksDvtEaOrJVQRqrgFybS8nLpnke3tyRwjXVgQEIh
r/+9ZSNFUvWkKGyU4Y2CMh29r9Gf6nYXpRlBOCpNl7Hhrio+u2wNQpAq54J5
AiRX42ljRkCfk+kESdFk6nlSbJGLehs0Btc429MIDq4HPCMdjxui7gOM68IO
hsdS3HzDPw76fDcI4MjlAXmP8uoh/75uFniWvrfJdQ9dB9q7rM8DQ3CR2YMn
HipZAnLdIJdJZyqgqcPEh53j+UCxONvKn44fmB57VSDJZLgbtqUfwHM3NWda
OWpve6Hd+mM3KNXzwa3c6/GIwGppsI3sG/yoFNKBRNXH8nIvLOGd1S/Vfm1L
3LNFPlG+eVUpeI5cKtnx0P4jZOjObFMs3AVvz3if0T9fDsNoAQMEweGaXR4s
gr8puQlyGMRiV7VTsyQ1MWvmpHo/RWW5XpwD/+t8AENR0tFUWTcLp6CsE/Kc
T5O2ezFtuznAFkiv7snNQEltfEWlf5y4j9CZgOnH9KpZyfwd9FEjJalJzRp5
zuO734u+IulLzmHwIe8pEOier0EOdL9XX5xEhbM81hDopIZ/fOdVpbTjgcaE
3XitFOJrxpy83YEm4qZyqWQ86l6HmeMnVub3fBJRbJStGJ9vJXQga54J7L24
yR4c+2tL7rLrUUTq3P14yuh7L7AV2J+26PgO+myLhJYH5y2ORLHEDfRh4gfj
YtjhENwVVcw8LPnOnv+it6kOOhLRT3b0zS2t4MTGRHU+RFQggu2xOpryi66X
ThLAuphegEPgEBwOc1Y/lAdisV5/qqNt0brVotOv9GgPZkSm4lsIkTReiz74
Mygbler11CmTAivVXfyVVt4dXt9pbP5ug48U50fb0xtfr0sgc+kPl0Px5Rge
XucLTih3BR6kg9Cyt/+TFStCGcHN1Q3ipgcH/7rcjoVJ9g/cMwvkS1gMzQ+I
1OUuYg9WOIjGKxjhPVw5PZC/68iDfecTEdQ5lOobJvQh5iaukvvVLfMaXoFZ
5fV9/9MzvUS+23xCSVzVRIiYHN80SSPwjbpAIVYHi7UnV9bJz+z1+gZcSqxR
CHuISQLyztgknGfmJlqXNkMqsLpNAR1A0exIUbAYpg0bMfdU28T1Y7g9uITB
ODP95dR9kUyEmUgRQJ4f/jygqOf200j2UUH+4kVgIe5mqabcCoDCbhcmbda6
OAqE/NoIlI4+J+KtzdPZRoxJFcvugq2XwvgPw3Z05jy/Q9O7Fz0pNuh4MkCj
0GLsDCSAKF4YQiPYI6C+dwz9yFmBPZnxQtjZF1IZ39aI/iHrWatYuV2/2lNM
edjsM1Hb9dO5A7CFlzzK0hQG3m1lOWu0UqoqwjIbaol5uSONwkPutdgpWe5g
gu0eJSnok3SSKZi6rmDO439VbzAsfqkovR0UA1OAeWdG/pwvo7bJkGVT1kPq
aCeC/5LiNlsHVqM8Ru4lgDcuKk+5tftl7BNCtI9qmwkhd/alvJ77spGcM/jJ
3BV80s6pkbaYY8e9d9HCXjD5f0TY2iszhASb5ceD41nxaj/YkAwyT35J/uD2
9moIf6H9NthTXPXPrCANlaPA6si4PcS8ujCiFeDbt2hHNKDDz7oa9U7FeyBm
mZyuOdKeFyQHj4EnPZWUKyV5ApkbT443C+0LILMR3fnODx5MsI14ok9r35T/
1S9979n7+VQKWb2pnb4guYkBOMgPd/u7l0WfYhVLjMUhr3dIxcO2A0m8/vav
EMP31+CP8STrlaVsqOUtjmh0g9IqBBf5gqS6QNS6Ap4bAQgVHEbb5IIVSWCL
FH5+jqZJ7JsEXac43sy40usCYIie+6glCPmWAe2oeR/i1Iz0DmfQ0EepGnvL
aSYTS4h4u9NXQBrVoRvgV6T3H69jZV/qbyLvMnLZQp0v1sRjBmtojf921jtw
zVpJWiIPWB5KE8P/Nuf5X5TMiKyhJkcvRO70HIYTMwf/CucJ98igqnKMfd2P
/nDOIobsz7Ih6TMQntinCOT/E+Kx0x1RNppnQMP7CtzJ5ytX8WSDYrI4O+xx
/x8P863jka4FfYpHzjbhqe+/am5QO/R7ukgK5kvjJb9p1X4LO/wJ72ETfSqK
WfHj5LQ30ajNOmm1SlfV0cW8B0mv79b2Eip9q56yM3CoOFfr7ngRA5FgHnGq
vA/LN+AiaxxoxpXiYL9Ad667omue2gF/0K/SeusE1SBcrEZDPAGBJvVGpbH1
1h65bVxebiRsCrAUkgCkFrY5vwk/izVWWZ+it7Rfgz2mi7X4DEwtSOoX9tOe
VJfp8YasM9/0mKCLRxOAsns5RSOkzrB0KkaAqL0lM++8OPm8GV5SKkQIn6Yr
/D12hvqnmFkdVp7/6Mj3ECEeLjJUE1DzZGufxhOOxcOBfW1FCl8DgwQWWiwL
PtmmoVU82ibyqSijjzMWx/Wz7aJr8Y0E1zd7p9Apl5Ter8W/MTLzFYwcW7Fq
RYwWkfpf25OiEOIxpq3igJyQ7XNj/yZMzJWI7knwmJzntU/zRek5CU93bc5i
tgshurlwyYitS7yr7VUVYXSuKIutVgo6haiec+vJ5pfZZ4+oUic1zmX4qYYg
PkW9btDhS/yanWiXS+JgSbsLlY+q/m3NkMlz2z32+l3dQCtrjvM10zO5KKWo
DGr+onHmyDpLwZnebhVFUxXv92Xna3ZElvjclJgsHH/yMhZ/ylCRajFGzbvp
Pz9urpppM9hfxnDlH2PADxKUutamholAK4CoeLL9bebC+aTUj6UZVZAY7ioJ
cLNkeVMcFVLDT1E3tosEzIt4HpPwBN+beiZK0he/csr4hOTkVKzGYvrhTjto
CtEtfn/K+BR52+QTIE2RoMzCW+raDWe7hOuRhe58/y8TJHqy0o/FsDYU8/5M
cvLCuFmXJBVHYhhNs4S+AofYRdn1VD8gwpjixLTmZK9Rl+40Pr4x9aTf6yk7
vYQ+2/nHvoe3mI+cxCRUoWwWjp5DnPT20f4JKOabZgEnCzoMTjgwlgdaIZvD
hp0kjBfpQJqhBFuDMXvzggZBFnb47jVz2jd4ZjNBt9lG+/U9Gvp70rZiSDzo
hI7MpwgSdLnF2vWQoDrdSgbQCad8J44niS24DQe+FfVPDm5PatWQM0MiQEcc
bBZ6uUAAabkD/3eQ8nOK4cz4ISzpeqseymAm6Kzhw7t1/+tjt8TrYHP/fXr4
jQFEfDYqUzCtF9CyHuXWXZYYHu5GOFH7OCmddvaU+T54flO7T9kHZ8wYZgQO
Y+uf2I7NqFeRazRW5I7BC4bgzB7GBVw24gxTM8UDuEnMzQ0PG5QR4wtJormk
v9XTJrJtNQVl8vn1mmbJaIuCcLys7hhd+4AOvAUKjKWuqVZ0aEVRhd9oATUl
u548Jb9xlOBFtA1xuv83CmOrNuR52Oll4d3fogAcYDfxIQTKEUEe1ETeaFLM
VFOdYPA68T5w4aSdvXBuhPrJWDGS/oa/PKF48ZkhMhg31/7i0tNgrbw+W1+S
zI2lFLmTD4eWwzDAj/Zm9lyhqst5UWgz83DxTBx5DeWEE3RrtfPN250kix0A
WfFWOwn9NP4qqLzekgR5kVax4wvJxowvnihFmLUBZmR7NDG25mQJi3AQjnRA
4eKf9lyrKA1aT5W4AU5YXxEOL1oNslFDj7s088T6UkyOjNz+Qg7MTzbgAGPq
5LCPVYbi7ZJ6nbCm6CahlUueEtIw/A2iIRbvThQNrYzqWfbZf+O2t4PeylRz
18GsJNJpahkIwCMJ23NmKf+SFkReen/Ab1Iv80TIxzlPQpeSUSYPt8kSYAKa
7P4EKXZJJJ6Wftsy5mFfOYfm9I391WbPswNhDLRPcTsX//0SF985QI8E63Bi
/qKLCC55HaTvYoy+EMUQheMXD5l7RmvrDMPRBCFx7V1Hr8FA8G5BQjSiPDH3
ZKBo7IYAG89QtntVHR32AWRJVUfRouIXCTpGvQtUBnXPzcbxmIZU+WUrJrMi
WJIMUJZI9ZDFFyM5i8JO3PpahSrfJvks+xyUsuF9uDVHeh5+3PsXgQNbarIQ
TSlbJ4F4F6tTOlIO98EMv/hCmzbKrtlz8JgQ0pqgzR2pgXd/xy67kzI9HYCC
5a9iD3DjsNj+59Idw55ss3hUmK6Gmec0EBECfVudA1Zy5axUn19eQU85dYC2
03hC4tYovD10GfX3YB6xcTSRBV7nWm97h27AYJagur8GeG0aiGkfwFWzBbN2
YmIJ1K3uPtT9cfyzLQDqyzskzwB8m/AxJa9pWxTDFtWq6T5MyP56C5Ga+740
cn6BYGPEjVlMToSoBFuKG+qr6gbXDufaSiJDy2Y0fvDrkRWpFXB5RJeU7vCX
4eUYAnuYs1R+kk1XeYAkFa8pKFy6ze1VynlrsegSLfzA1ZNqc9GGO20xwU5u
deHBe2hla1Q9HqSnj/yUg4yeQryKonc4o5Du4nSuIoaQPGFpOg60llCI0NCM
QtLCTKplTllIJmOqCKuDLax9IG9rwjiTSHz6dZPsmtj7yTrSJvq61napn9D6
ounfuwcO/dP96nKlL7IH5npLAo+UcLGlczRMvCXKfKc6l8TBvqCGPgsXlidI
cHsde4K94ITDfryxn73c2XYzGNNW2rvZBOHAs4dbcG3usWGyOMmSgRj/kXYv
Ri3R4TuvX/scB9U4v4grk8hJUW9jJyfswFrKESA39h/ZCrjY5DY8xoweruzl
Y/o8ANf5MdFP9VVOmbLW1iwuuBGNaIna7j7g5suRclr/YpyDkfQki4rtqdBJ
ot0jx5Zz1+fb6DRFVne2B8yMEJVGS0O4NH0Gsl64emSqxbgHlc5hcLRZ7xzn
q/hy1dkokm2q4nXZGPoNl9QQGDKwJZ8IQgWNmkSsjb5AEe0pMHbCKNj/9707
TR+wLWqS3HpVYJ8iaVnrQl6VWbq1aD9MVOLvqt6IjQ9U0KRfwGvUAxeBTa6e
XTyasi98HeX4yQPMfbmpF3zML2BcTZiWi84lesF1COW7f2I7JfF0UQLSv9si
bmRElOjqPAF/oPq9FnxjnwdbguuTaM5E/h02laSB3ixPQPDEZff7iPmx6bj4
MFNNMJvyfVA/nW52+ky5lpxnYA9GiG5ZrWCfdyasBV9yrUMkdV9VwZOU+zTD
NkhCZ9S+3AnZY5G0Sk02wBS3lV+TW7HY1/AuOo+PuQcl8EfNZwHW6sv8GMZO
OtfBc3kjX7NToB1Nhc0j4j87LTg6GHkmmsY+S5L81+h9K2rrJwGak3yzrix7
tqn+XCebfZiYcw77qAa7rr6Q5hW2DNWbKIp8xt07shOtONkdPtVVMbT8UtOJ
xdrKDo5UlarcO6phzagxYdJVYSniBe+wkATSrRA55Tw3b6hSiwHtOrGG7abd
v0T87RnMSbMW9jEv2/z8AeKK7nSU+4e0QONmn+/PMu2jCN7ANP6CzPhJutrn
vDtf0qOg691G7NbQpME3hOKaXzPwoNPOfZ05NjQfUGKGfJnn+U5ETI3QlZyT
V0fdCd0rgLbIM+Px6LP8AbaBidPszsvJ67y7bD9Dz8q1nVNzV5OJfCRlmEKA
W5F+pPEQLa4K7XmevA9YwI2HvgD+NP7i2Ui1GkY4zX8Nsj2BI1Fuu7ISudUv
koLcQKkGM6GuRCtM5SSTXRprqMqz0GLXoCXkFxAnPg0D8TbF5oRRN9qGDBJl
xntyxuVBM6cc061Co+u7dOZEWlDje0+aSzVVBL+4urxDULc016V1Ec57tHxv
plcU71WQM+COXBtAp16/E7h/stvG80ZYIGzuWRMEtoOudfFJb6kX71zbIKWK
pJwffzf0NqtitC7rDwCg3dv7lVw3hJzMCIsOjpU/p9EnVoBxLI8yhdd+aaGb
U7bpFrVGwyrOfPC+hIvmR/nAHbOIKV23IML74SVtgVXFbeirPo57h+DiVZmD
SFi4j8Yr0tEy5+z2R1cITM8urc8z4A1WfNBF7LcAJqGWgYy3A3JeUR3puElN
VJb+A0JGVgu4fUIrccuBOyue5lhyt4ErtBQ0RJGPEdzUaSeb04UQfUUwODeb
Cc9t0BXNI6sbVaxWPbIH1B6F9UEdH8njXF2RviqI0R/Tn7KqRIgMc6Yxg+ow
0XpoXwdaQ2S8qyOx2jQwZrGv54P//tE6Dwf6yRy6fX8Q4dzSPWtqd3olQkaD
T5I3H9aMR60SMMQBMk5mUU1PWxV6T3pmTivM94zVh3ze6EDAo59QtKqjVFjC
c59Ur3ioUlSQROKelIbNvdpD9kiWIbVP6dGW/t/X6CbnqKpA/vcUgSSpGHCH
FmLfaW8f2AOFbX28fmD3FomsRhOdqDwTOH1+0v+KFKEsxZ0LUqu4tjLQZX4m
Cab6+O2ROmJGJR1mWIvuj+YNAARX02b0q3+3vIjgHzC+0/njIRz3F9EWG6gE
3FUENeqFVmrQfpmKA10mu1T2UQpfIZD/epopWsUsu21ehVZNKu8Sbhz0Las0
dIH3kdi5Quo2yQKnlj1NHCaYdPug9sSUGruITmLH8grrBSKucJ2qeGhKVgXl
IHlJXVzdCwmc5CXQvOicJ+ucb8CEIob6nBSt258gsnTltrufFEvMWRfHeo7I
QFg+hPmDOt9LoGNzaASnCxLgFdxPY3dQWPk1BP3/GnrYazosNg6IxWt4UqJB
mb5p2urnb24qcFZaKaKfSIrUXp5aK+Ypv50iRWMJR+26+JutXGQmay6vK0ZN
OW5mXIoIFOdMD/3np4qiV/kjqmPGZB5NVZzQ+DU7nBcdK4hdRLe7qbmEnGlS
USv/nERgIxw3qr90yp8O2vMMXZ5F1DtF8S0g+2wjnRbKhAPd2b6RBGQ3J3zX
4z85LVedgXM8Hb72f3LnJzcRL1F1LLAXmsXoVy7vGMyBZah1rOi+esLi8NMi
4NaHL3S4/s4GEOgwZj3YdkMbcczSJBzxVOVuwTKLp7gOcWM+cQqVp35IN2rN
jbo6zOw71zW4PQ63L021ctbRao2WEKGdJ9N2Yu5tC3Z6HR6XKsf2djmYe68w
X3wgMTtAGlwS3V+EZcOCXcECjHxQzT27elt61ZAtPGEflws5nUx0dSDRFKDY
ZXCsZZ+xwZCfOdbcnlM1QKqVtHxN2wJuLmoAjgDGz7UT0JCHJl4BOoxdgqXp
qPfld6kMVqZX5K4CPULVdTuUG3AU9AHM4EVvIrJggfoC2UotUtB8iHm6WMTf
gU7jMmXIOOmpFEJlT8f3FMi49NUj3gLdK2OBydnBKb74mVwzBhcEFtqPO5kV
xSOUTls2frW8ALTo1Hj5HXg+usq8SgTMlcEh6CYnpda+/NZzV5TT9RIHD7zS
RXp/RK83rgozESmkCr7vhEx5smIfSO/7LEm9EHS4INfpGJVdFWNKvBI2uDrT
dGtB1ZkHULDvutoCDhyhkqxg/Ueug1bEremIDL2phA6xs4tVqQ6eGXwWi/gU
/Sx5z4pMcz3ewIteo9NMYwSvJV3yV1GZV0vppEUKyLWvjp41Lf0I73abXu9G
dems8TjuB+JJPaPZ778tzfJYntG3o2SNxT8P6p4eSYaOSfURXtEIBJnBkqkE
ZGHymdBF9eWYduuumj6laCxxkd3xMBqmaEdufiYTxxIJudvg8SIEOcVbFkAs
zoYzeh+GL73RW73xfiDbJeRl4XKS1FrFsdZXoWKLwYK4PQW7q+hP1x5IWgA/
6dpH926pqMjks/4nKcKTLA0zvyk9Ix4TT6Kddf+EVf6UXCtKbUBzKRroC+o7
N3QVV9i8FQstdDKChsg0I0fxsqmU2T5Vx8Q+7SKFmRzhNobZNy5QWod1rGu+
kONqaly/fxzQE8ajpykBzjgLqbT/Po7gtf9x8Jtmn0Bppd0rPQROj0p5vr8V
RcXsQyqdKYzhlsB4pXgVrYhpR94Y2uiFzEgU7EMjfreYTKv3DFIAXeteAh3D
2a3LjPFANb8MXRpizDwjzYt85WuNPneyapcPQnz5HiohmUenqHiZC0anRKpr
Jn/dObZIQNGp22paQ4CVUUcYFsHJ8YS9xLIZcO+xVYdnxpymx4vUOriEhmrX
Mais2KtTsUKTdraFTyqTRRtdc2VT7R1h0hVp0KcoyQ+czpCjW/G20akOF6KS
M6LGXuefrfV6tzqpLuLYp5R45OP/sKTPA02V2NoKQnT4QI2JKCaCu7RcDI2t
yMlrFZwncvvEIk2XmEob1JYdhBHuD9foi48nhJg1Qaz6qRpCHx3vz022ka/G
VhOf8/ePMpogwNZniK8RfR+EKbY/RBPOM8b1xtaCFJSHo46mekeBB0mpXWgn
446/WoW8/jFjafUaOfA2oLpB79GFgn8gg05HjXGi+YjkM6sOFywBG7dwuNOK
cEhH9ma05rZgS+aVV7/tIrSfDb1edPzK9NcQefQtIDl+JnLhDStOAnhZOnMV
mCBJw0nxVZq6FGi8Rp86xXpe9ck+cy9/RPX7mciGAle5iSFYUY+mYcn29rUw
JJVMXal8oB6BMpaL8tivTXUEV6birb+O3S72LIwIIlAGtQMzUg9Ex+Q31UZE
VcupT+OU7piorXrAL+KX4LLXMqptIBJ6sueqOfa7c0nlmmnHOwh0VwOh270W
C1JjpNU8RDT+kgX8/fZuTxAAHxkg15ha9yw3oWEWrquFRpaWX9WcOCIuNUna
jkYGskg2cG0JzEWD7rHRxQ/Lvg5xnsxB6VIeZm3WPq/vPVryVllh6ybdQbfq
7fxK7gBnr2Ihhj7PFPjE0OtlH3lb04ieUutT8JOuDPGSE83k1/BMIiBIIt1m
M0EXsGQqzbWqHEmwzYQIMECRb+KxlbXYZmWifOcNe7QCsL/dmAGgWBjO0dY5
9l0uQ7r1aZs86GK3w4HyoDr/ujIG3FqjcKd3D4mctvNsKdMVf8yneX4gshzt
ZtsRgfO0Gst/dItFxDFGbSUoee9x9YT5blpHWEQWWPI44vkzgFHSR0yo3WSt
ZhQVx85ToRgSd4H6cx8sy1rshtDY93AGhw0/Zi062yGiptE0GqJOF9EPgmUr
VyFJJWz5hQsVdqQr2ZYkPpSqRLas4BSEeiKU3cfvjnuY1xqrkCjthMxzVp5P
6m0sPjJy/uEtTOsiEBagEIp7aQFZaUL4vPzO6IJ3WMLPrK/iSoUuAOTWsX/n
9L/3EnQXONLm8gTiBwkYcARgVO88Ji9svHUTZNUjberB3+hEF/mhuSbowZBE
dqoTgiHaHbZ3uTdoMg2uSKTQc9grnPOHMwOZ1jjwUWVY6YmzZeQsmfntPyyE
XrD3/GUTp0dS0tUqqFVJ04kox913VaQQR4beMhKI6X7O3rLHHCo3AoPacnWD
/bSDWtvbrm7ZU/iE5QWJWe5aGtc6ZueQsi5cP/2cLLB2ObW44BD8mKpQ2u6W
6DV2/dlXqMk4aYFXaqkhiQG5Q1jNnhklbcz5RZPp0nVAaDjMFlUrWSKZH9oK
UGRRnCZVMSqmTOHvP4VgvvBkeVTzgBS5/nev2PcVVfOjd+clh6DMiAhVeINF
Z8YcFvKzOdV1rbqlyIKX6DPLmd9NlsGEiXPDpEqlhaXtsb8N1ttGZ4ueMJaU
VfYpgvZHA1Ya8xWfobMs6M7SdoS8XCcxUJ7SrkfQTBfjezHjOfcj9KWKoC3G
d/IS5V1rlaLpHAC8D6Yi3aLAScwceWCi1g0kzqL3eyjDpbqHvNcXz9bQPyzN
GgBPQPOOmm5pWGBlZLpgakU1VINC3SIfjJHrDS/bqbVD4W/x5GvefgbJ7Ljn
VC5pe3HAq/48t0AFO+TsMofeDb6tH9qakp/lbrbL+qaXfRZuQqDnaqKNin0C
vLaj2HW8684Ex9ediN+g8bGdHG2R8YpCPxPGTt91O65cYmeCFxlb1WznJWST
V3BBN+D0J1oWpBQLa6O+GdeQ9XmvMXitsNbJsLvwLnkKSNG9J7iX538I+wXc
UuX2FavvBFfcYPNhsBdTYxhRBmRA5gS34zqp4O3J02Q/N6xdr7hdUoURm70H
XFyDgQ1/Aonl+ACSY2QX05U224ciSrv6K8a+GnDioODcrpNLADoOKYCNokW0
NwiXOXs1XNqfOHucgcyyMhsCoHV3D8KUtqNePb0hkgWyG7Pa2uvSrGqxmRzG
gK+UWESGbq9d/eV44BQvuoSxc6+P+LB/9Wte/PIADFEYI/sBIZjfmCwARoft
GFBS166wHznpbgvY+37PJkCH7ijv2dAogGeahCSVyoCzJ4S8BRLeIPtB8ySP
vy7ey5mjNNnSLsXT18cQI6Pf9y8taKs8fL9r63c2IpdYKSUUOAlEhr1O/NCB
FjKnvch/ZnTgo4ZJomg1XwO5GgFf2JWV/3W7XIyJ3AgfcoSPiI6flLItIk+i
ZeRAQwDN/5c685fgz7F+D2nXBclD3mVSb7WBUx+lUlIRZNxUCKBs85M1OeRI
DxFu95/CpP1rcOwmnv5tEt4FWPbWN2V+23IN/8cD32MFm13EYFCCKEEHoXbn
p5BPSgKUWZKaPSO8luq+Iv+bJK05CJcG1ZL//I814xLOmsreGc1tHzLJjRbk
G3awrh/Rax+Vk6uzj880BXKs3+mreIKWsN6ZISRagWYrGjGyLO9pzHu12vyD
6DchKjkOPE8s0HzYs8q2uLho2wcKDqkzXlivZwbD5FGbvPV8pO9yivdghzKs
aTvIvyc5T9uvCPn6KAM6q3mNXqSE3JcVjNGkt4AzPgmnegWc8SD639bKRA2L
dHrhO1wo/5TZ8sMbHcFnzA+z8cp0avPHf4K7qxUcxN2Psb/3LUq+XGBeoPct
pcdMl8pDa5fvxy2DsFmwq1obJGl+/CFn3cxPrZEEwVNb4d0wX8nSrNZpAbqQ
7EMHeM8+9BjupxT/hH3aascAXL9mBwaTMXJjuJtn3c8ADzAACb8txGwJ7KjY
QC3wqjesWUIjA1Mu44VrW9jBqD3+DTEcxR4ra7VMA4EEhq1n8iIx047EJ5Ve
+wdmftizWsvxKBp0rAtbMkXeGpx0S00J7fTbPotDtVRgbb/4kM2XAV4BJWpY
/eT3KIR9E98ALzzvk0mqc4AwURl0j4c1mGahYnrmaqfHZypgPJS92n4PB2Bg
SIBpoch5tfk5E3iG6PQR5E/B4PC+soHSGb0vNvpsap8BNRRB978a5keqY5F5
BophFmC0q1trllA1hiawOytvtwy2GwjaQyYfjL8WqsDZ2Io83n02PAqU2VMX
s9PpIvdn3FSor9qQ2EbdI07Zai0u76Swk17LiEZjGLYJsLBOu8Wj0hp7ETBq
jzZvG1OVWjNMC7HQGpBupp8Xo2Zgtla6Xk2YpadE7L0oJzHT42gJTPZResaf
NoBosVJT/D7Hz/CmATPiFAtp4Ej3ZrESYTUtY5mkFOebWgQp5vDEMFot5EGa
q1+NRPhDdQP0A9OjWOdeeYfKaCmI/4vvYRHFxPwIR9Tr6DH5xF6xuNhsAI0W
FPU6czPZtbx/1/+dNIRJoJLJZe5JcQHZz2OcQfOmLj8GEq51M8xXSRNkBMG9
/E3gsmtfwdDhIkLzhg8/HDp6y35J+5ddlxz7PVM8+VpDSesyLH1+V6ZXtPoc
O8ePE07/GsT+6/F6WhgTl5/xU5FtymwpcpAhRw2YGilrIBt82UOeG5NmSFkc
iWl/0LPsHZMdD0gNcL0/d6P1ka0c1bQ4j029aeySoM5hfn+/Oh3Xq7Ud5/wa
9eQ4HB7ZTS6t3mkQmCkDWk+azMVAvFjTqleajTFNKCdPtRCRwxCSQAZnbqxn
GQW2CWyuc8SHL9xULHdHq4jVfqeIut1SyfD66VLTvwNAktj3nbTLHQ88U7qQ
kHbQest/0l7OtTIUjRLY+nqfB0YbVJwjlvODRx6tRA3WsFjYRPHh2BcVi/Sh
qmvlMVjypiwzdZVo5Z+wZDAglu94RtrU/U9gy/tdkWrP3E7QfgJJumoshHvG
H6MwjJwXbOchqYP3iwk/KhSXC2XHPj14aPIfA5/Ih4tls8CfAXWVYmRnBef0
5DGOv40V6pTl/kz57LvDK1Cl/Mr8zMO+iax7NxDVXbRpS7W4J6FsS/Jc46Gc
Rz+3lgS/42RH4YJEPw7gYJk1GaaR+gVQBnxTTIAFZdi10jY4nQuiKRNQUXpz
84AlkfyWlc5furCN5UbmQPJ9a8kmimqLLDlBkIhpwX9TkaqOCOsDVgGnK+7a
BuAD+031G2Zek5k4C5qAPTcidBHykb5Hon6mFMORQOVRx7k3S/j0PseWfXH1
b7N8ucM+aIBBpVIkVIn7NxEnE8J2ZQCl5Xi/yVOgHwbMgSkaBtpL2D5KAlv2
WaoGTibDAGxSxetQ+Bgp0w92waQHt/1c5NXHQ6f5hCdKSThGqISf7awPRwuW
rEdA5jxglGCKKFKjwRQQjdPiTEi654XaxFN6nuYJAnUuxz8O1lORutoU3Ch0
zRhVTOpm/CU4w1eJ7t6mcBR24FPiXXLpkPU6aBj23YM1VmxuyK9znCWPegi1
q6x7eBKsD+IfwUxcE5DNyWQyBz2zrTzIkcvFq4CK9HK+8AYLNpoe0hfjygFc
XYpMRX2GW7MLhjXCi+tRmkRLg6NeyFca8XLZJjRP1l2kyMbyzu2c/1hgzt2a
z2CyLUrbvAlMf+6IJ935kxTWOAfNzmWtfimxUgrA40qIrTTT3wBOkdlkth/K
ew18m/B6bPWsnCkennKzhN2SqQlclNsU1DaQBWN+SDRx9UkdHqY1tKImSNxz
Kff34iol4unNhKcifwZSPAXZ5zMPlmpWjCHck9XPbAeYvI8zqEd8b/mrxheD
P+v0+rMTxg8UxYd/ZkLOYR2K8QxjsvBD0KV7r+LpdXNI7UwDDX7lJ08J4mJP
FvGpTDOx/dgeGXBsiEzW7nnP7wo1w3XCXSz+Ftyy5pTQnu76Uf13RydukPUZ
TZ79qv3Idhf7BXNypDxFSQFZAVUVX1Z7AHbnvpCaC5MliXOmWysxUvQRQqty
OG3w1GLIsPNaygTxQEgvescfMQbynyamaG9bcxqFZbOeMdXmyB/0oIHTutsF
kp0EHmrQosJScJVKNOfUld575StH05RoZv5jatdDOrJ0QQ0wiVgbHZdruUiE
MLDYU43XKuJRp0ZqAhr0cSFZxz9pV2UuPPuvVxu15pK1lTedh3q3Z1kRVCWk
tBbSsHSYUudkJfcawWhFwdGnLmixDF8LEl/sHTLzneMajJJkimMsP0OURDTA
N55cj3c2t6Fpkb4KgCo93hb3Q2wHBFJMMmZBXRDSBQjp0PXzlYsx3G8s8WUr
8sg8pjd8n7azPCGZNN6DihBS7M7IZkUFQn1CYhzAPr2lJ7vw24AgoKKYUPe6
GSV5x3Gg4DsZDmZUwDpHQzaJTjjKIC0fCK4XEwqppHJaTSqWevfA3AYFqLr3
uDU7xr+RK5QzNPXmJm5m2DJnsNgUs+ZywU4o1aan5t39O9/ITtl5SybFbA72
E7JL2wRKcSPka3an/uJJAgTvvozY+/uLlaDDw0mXd8wlBR/+C+10cEHXbaYL
T8qaxkR5agF2cehtI2xnz6RQElINmaKPoy/g3Xp1CeuaPBgyu5W2+DR7iieS
0wN81YrNP6vCkEJDkmDt6A5sgP+KX/n8R5XSdUBbg3ihwXigMwRglQkYdNuf
Kw7Gr1arU2swA94ZIyJjwPzmCB3MvQP7JtWXKgL/WMt3GSe3zNzQS5WWvytN
xQqSPG5grpbvEGLaQUDMM+wlXCADJNfavywbHAaTwBppn785Qu6gI8n+1eCK
IBoSf7BByjpThu4AzStwlb0NOqNVJl1wdW5uLg0JIC34jZ+3OKYd+IqJoaNh
DIw6u+DNuifhm/PWfVRWBn+9jeuKLu0sPBNEVABmENJ4ZnnKRrze3ne040hi
hwSu2Y7xgL2/D69y8lLKR5WpQroV6wsxrG8mteQGPN+ooPMLs9+m+WQl7p/J
GEiDSQXKB6MCpM5itD/W2SY6vF/FOgKiM9tvj0i4EglOVz9XKTmsz+8TzinB
PNUwIF+R4u3SjV89kYsxqh3Wp89LoOu9A/vVS8M/2Ixh06jkQOiC20Yc0vJ0
G+B/qMTae+BeekmlJX8qLD30SI+kcIPyJZchRuB1gbsJshEx9oIoX4RJXgvJ
168UXoXZNe5g2XAn5dFyFAEb44sixmV7125F7rf1fvKg2xJ+3rS1CslxwEb5
Lir5QVad3DXqXWqc/2FjfbjkaqpO1IJeBfI19b9Ca+z3TuperYhrsu+MWega
q6cYo8Jc8Z7XskgvnhNDDxhkAz0Hh3iOAAc7PdBl2U9SuXVuuS0kEdu6nOPN
agvBsKpdBwltLG8KvbZ3QEeS6AmLqxyIt2cwSTPuO7zDLCRpKWoEuL4a6Ssk
3W0OSj+CtfItgFxe/emYS1+bka/3lamdaMOkKEP8gKHtN/7GzzYOGx2kTNSA
JQ3o39JNgt0dM5L9HhCFwDCYTc7t9blruOG1zFWJfx0evEWxHjd4ZjH1shaC
6bI+5C1aRA9iXk9AZjpipCPtsVHVUSXwBhw1JdzTSyxWhIch7XfBsDrshFxe
eMTUny1wVpuCb5Ux/j8APTtw7DbJ7udrdYVXMPUBVIt59rV1SPT2sK4TfB8j
0wcI7EA1UZnokwIksGkSV6rbLfciWbbBT4dIG+BGZ2UFkLwgCQTGQrbGD1Mx
IC39QvnmGLavDQTYzS1MRgm4fJTzTSZSqJJck7SCIvPJLA8frcWcREhMiK+k
CyD4AUtUz2naXu2dWb6/lcuUF+04vF9vW/teV3dNJLUmGpwbVCpRRqGIBYNU
MpnG76DI4ew5t+U9FyvLUl3w+7xvocamvUd+TQKAz4IE8BbhcTwt+tWhynBx
79gg6pAbFVSGY1cd+ZhPArX0JwC3UYpSiGCCALNjl71tkeXBoEkI8sj9cayy
zfSYx8OT+kL0MCe+Uhaq4IwSk4A3P3B6sbW5nQ5PnHWzs+jIHqHFo4Mk8sNV
79lmw5TASo86KIWthE7st5SRYt0HadCuJejtFbSBUudEEFdWRrv9yDMQoPkY
Z46RQI9FLkVmK3VrMgpUudNeoglraPEpBMXOkBdlq2sK1dEMVLEvG934tfNS
LFkm2IwreWyo+xIA9C3WqhBiGTBjZgVVr8Aj53x4+JKSzSerbVtfojDknMFj
xPc/tgg/taSxFzBwiizq2b4Lm8fc47vIzdlMsaufu8bRcxqXrzuZWHsoyDas
ol9pUzUHNukD8PP4FLwysZCR7UrrZU7ezjRgM/ABgnipAUBWwUzGYqhjAvD3
adn8mRU1t3iLppSzU1SfnGrhGLRmFvyJjJ/fyj48mgZJBbsDXk9X9q8YAKae
JeKiTHaY9MrP6W0en+uTML22Rqxto1DJcz/xQqAFykmASv8GTLkJ7NQkrq55
wpGm0/yt5DP3V5BOQ7aZEk1MEI7EzGAAupc5oJJw9+zsv9regixP/frhTYNh
RVqiOFOC30wgseNULFcgJXGDl2o6H2SUrgaHJ7XQ+G6QWfmGyLUH0Z40pG5T
zBXAvfQQUyjVDSYRKkEUJV0iJh4B0grFW/6o57hgDzncLrcex+fvcu0/kw3I
4TZ/UEm8DBoC+2SY8TZ2oS4ughVq16MW4mHEgS5YYbDacihvbzn7LTn/CWOo
IZvEJlYqVkGOUcOIoAiyWepGAoS/sTHmf9JSlXMMIBOBztybw1StA07K+qRP
tgOxEBbx/l0NqDYkM3Xu3IKyKkt+qjHKsXzRFznTN0O0h7qxhWAkik58fm/u
q8Teglos+11uwYzKqim7vc5/mmNTVOqo8mTQJLjdYX0YzltLYpWEUR+ur6qF
ccLgTpZpfVd7vrblMQ0aty/e/38X6ytzMfbwnbjnwJUf7ZctNJ1cjYU4YOJS
4eNbhq1sjCT3CTsYqa83WLbDrR8Skk8AC8NQck4ArGzORdX5nzxz55yUivRu
vyqwH+juukz6q+ZoGGO7SotNsbm4ggiYHDiOA3TaL4tvhG/4b0zfZHSsr7gC
l9WdgrLLaT231eiyRcTMcFg1ZQhITC8Qcy5D0Ic9ublEnhSSqCIN5EssPV76
f2U/NEWdGUfwf9aN78FATdWtZb9CoNIr7WaiyPQh2UUDrrY4XXJ/3fpXxEtj
8XCNGiIBFf1slrdRjrl4sJVjQmaz8qUcyDY8PzO5KN8MHEpBWEfGT6M8hip3
IesUVBLTIvv/f08v7507pUWcZCiXt3nUrKSull6nu+4Ns/vFhEjCCj8RuPf9
2qbKgLjVl2lUxeAqy7w/SUASAhMjGqD99rdNXvRPl+dpVobWqgFsfCa/5U3x
0tVQXbb1cN/hdGQgVnUCdniKsSvD6kCHxK8YVKVzMYT7jl2vJJFhYfClnAf+
pOZX8psPieyOr6nRLNK37EURrjtk83q2z4gEt810I9PiwkZQ3uRY+NHEBwMT
O+aOf+HBdHGdUb+ZlJQ5wUTfBtU3tlezUjpyD2hgPwQXo7kT+Pd87TCyY5CV
x1/XWq/cfgJyIkCYnevyWm9RGzCzTVUghiqP0OCbcutHzkfUPbSIThJfixK4
s1KawJYP87prLNKEElhgZ1mygbvQMJgfT5tcopM6yPSsywNZuWXq7W9HG6SM
29/Pz6HcmrE7ZmQqiNOoAo1U9yqEib99WZmYcCYxOooRb/O76E9esrh9xB9I
rHzw/0kbPeOSXMWqCPPsRHcfegEUPitbnVBkPhSkUL8M3AbPYWKWmYtOsMWg
9oMlL/dgy+9POhEE1UlImmQI/PBpK/LpqISCAg5nEEricFeA7LAkEJQ2Eevm
n9wrpTcJ6h2Hi/2dvoRcjbfJTZSiRRbqvZScsLlL+3jkWl5g1HmNNhMZ4c5M
Ub1VVQdjwwkOcjVtYjfEYLn9+sojFAlHHiIxqu7D9nqk74qc9Qf0/qC0Ed6V
SJoP/sQ1c4vhkhOrd4zd6gSWtF+j77zbdAYLR73hprtu3TTPoNm1da5AHGYV
sENae8e7YqeJpbhxTC5xq4dBsKSi9v2SJT2sTM5L2DVgdkJ5N9a7+wGU/n1v
Ud7nw/tpSQkgDU0CIMdEf1ZYmUEfWmSraIPpkc1iUN1oznZ+okOc3LbcyPK+
oPLHOR3q0TcUhDH7keIeJOb8iHzw8QNk1Q3KR+9HjCFZRcOJoHLg7oAJuQFr
UkDpZj6jbDCHCtK4aXYfT3Gz1gHkyzX9DW9JVJtAFvqA/uGqSZwFPWIZIhtB
e+X3iD5m3zeRk5zW/3lC1SSoTXEsEiVm77ODXW6GK1RUgY1jSFhkQzfMuADJ
2WTPwfg9pc9QrVZx+BUELxHOCUItwTT/xIQfcQYu7dFbAnEV1f/+Z796bzQV
rMmfP/sKlXBa0sAc0f3Uyb8YXfkiFG2X800RvuWBKp8y+W88iFG4bP10rsmK
MgWS4xMjz7zt1iGnSF44M5XP0MS8aIDKWHJPbBz/5Yu4YQ4nyUoal09L+VXh
aDV9MQxbLRAmZxSaGVgDSf9gUzzYnqnEntkGMHR/pGNq2BxWizVzhlHfxh9w
8BePC7Q1DSkjbxsMIhyGRFGyCo9xJF6z3AJqEiBGsw7CnLpMh7unTHnTTCwV
S+//c5WdzeDO4Prj7MiwxBK9P52q0ALpgqW5GVy2eKooLd1EtEDYnxLlfyN7
u3mWQuSpdVc790bmNOz5RqHkkTN2I8Mqq/muB5IRKmezi5lkQeQpJIv92rBu
n6kWfpmBD7jyqs1pxdF7kuS3G4TDtgHKJ3sadF0pwWhbcz/KhLRgQBbFHrDk
AKC8vjTVK+HUYz8AXkQV4qSVNFUiwZMBLdbgimY7bBnq9GXYeKa5T2/zd367
f8wJNoblR3Kp0GnKx1laq9HebW3kWthyZp4DFZ6NvXLKGWeGKSy7HYZ537JY
0uGf/2f3K8ZqQXu2apE9vuuhvNuzQJKQ8zZ3QEG0mUNcJURrs04jTn3m0zQP
vtZyex8XNkUr2oz222BQANFDgMyFjblV8OspUXKFOjyDVZIK+FLvzgGfplPf
CpEpEfv+qfWFFRR2PVT98AMAPbnIvUfAEJawAzV9s2JE0oRZR+PNXBriIvzi
Zia5xbIqAi3hxZJaPeQ0oymJS1WVZXAkhHNUZr3aWuLo50SDQN5weYUDxloY
RhFvA4epcIfjH33jQX7jUe10A8S9HvJluV2BGS9UTBbN8VJD7UzS+aewgYKJ
ynAo1OPeRt3eTwJ/rROnKElY385S1RHPSpNc0hq6GKkjYSh9IpvKdBDijP+O
PEvrwQ+in+8vLUSECm2uVGhdN0n8xdzZpjIWPt7SQ51MFwCThVgxW0h8RA+z
Tp+ZzEdSpS3m/a5MD+pCg6QdUoy3ABqTXbosMlJZBtf0VQU64aXz+I32qVP4
1gJisE/7IjLsYmGHMNCge51JA0K5HZmfDUxByKDE96X/OB4jg8wEIkzeKRaA
xftrXO+fhOh46/nRXmgTzcIoKiI+qjMoEV2NtTckIhChq+uU663u1CJaBSdi
Lws+zaAZ0sgfKP5FawxqoKXEd4hisCXY+aakXGflTBg/G/d/rpbsedgQZXg5
ZRxXonTR7xZ3l2mBubBWgo8E/JKY0kL5YTLPHgb0eyZVUeZYyTimXfDPsfEC
/WQXSsdPwuzeDoQf7dE+lhHTRhl3ogs0ahUHfyj9ldIbulL/RbLMNByBtpCs
RcMZFmVwSiIqEKqQ+oAZMoxuBqAZ0H8E/3a1TP/XqPXs0bfeF3QcfONdeqLV
AClRLKD05u9pe0llrWTVG0TFhLwK9pwv7ELL/4j2kJJKOfJcMthTtShEuva5
LmftPhQrQtbDufVibtJ9lv53btEGG9JqK7TxLelVTOmHfPvEo4OHXG1v/vPG
IyBXmaRCVmG2xC69kMmB5T6E+AnbTBlM0ocO4Yys0S38R9dpYAPOCYGx+4ry
Gl/CI7QWOzIaNaIHu/AkSFIdu5bCFA1EXEzQhd3YRZ3t52YLSfDOxBGbQMnr
5KMnLiE9tN9UUSE+hxGQbT5D8TDWJbCHPekTjJBsRYNUC9LAnnxzhEcv5j3w
RdrUI8Z+w3OIkMSCzzInXUnAr7eE7pn8Oh7cuIvrPqzCnozdxNT3E6kCUJ5W
/bJblaWdKdrFrP+BQFReQw9Spw0QNLTUUiKOiiaU6J0r3Tayg0qtbTFzq7eG
SZE1EutAfpma9Pz8Mzk4PsRUz3oQr53CmvycUeOnnRC+rRiJ6gPez0frubNH
568ymKnlwf7muQRrEZfXMxuU48vdt826NbVGHRU0DDCDYHA2qDBHqTzcvkz3
EGL4/3st1J31pU3OfsXHqNZ1k+AdE794AjVLCMdszuJNBNpePDmob3saiRmR
hRrKEeOoAnPUgu/NgAN/5l3brFVZIwSt6n/Z63CvuNWZRg60ZXgyXwcSQU97
7oSZ/j88XwTcniY/y+iTDed4AGQPDrDJJSzZIp2cMjaIFGblX5nhQe70Fe69
yjh6XdrRPcZFpPGFW/gbzQVYkm48Dx0i8nq078/K4AQmIAV96A53RVkN40EN
hUbWx+9XO0yUsBGAWdqgRbdgY7bEr1WNEwp4Ohyr0w6IoMZlXfjy4idFVZcB
LGOsqxhMUijEfxrG5K51FbyDq2875ABpZqJnkNBI9Zd6MO1STWr0oIbocJyl
Krm0X6iKoTgw/KvBWazi3FBos5ZtCWpa05hxwWQlQLbDUjaC3OyQLiDlZPZG
IEpPediE8734Zd/4r9NTSS+g2QM6lYU0aNWGnc+lCF4AwkiWOC9BXQz3dYd7
gPzz311hYpzcG2/XR4yBaXQYyr6X5H0Fei9xlGRUk4PlnqggIWh8NhZQ1A/u
JPjEGNGIw9L4OSyDUdJRTehEYWrWWUNiIDx51A3sIqTcHmgONaMFy4rLZ+6n
vB5niX3764YscHJ5LKcpjN5r1BSHXfRS/qD3Rhl/lbOJ1yO2Sbdr6jhNwXx8
/9SfBC8NR9EtD+l+tAIo4s7b5V8kxJEYs4zOUYRjT61jGLzfNubaoynftdWZ
Af6gZGZxhiO7zwam398GwbJJcCADqtZqk4yuSCzFJF/r5Rm6Rbq31v4077dA
hkftiUqFzwPbe3EIoGUfPAqT7UYhR4q4O4aNJKrsqa5wza0Kv8kzKK/Bx2lH
TsOjmEVfUtvgvfSkIMXWNqejRr4HQnbDVG0RK/SLEurWGEoRI6V6osktveDw
5BvlvNY1b7A0rYdOwXtkysHpoTxSEWNoPKw+fDRl3OZHOWs07EZ6ocqPt+wr
POMzGyMCew0cb7GkXS3EptIZJ2EeryQ53zsAUEQoVSM++soSww4St+qMp8nj
AyndfSOi1FbS4h/WIYSdMBz8hdk435xYBqIrs/OWOmZrDIuQVCt4/ffikw8B
m8tFZa2/r/AEwv9WjIkAy7z4d/+7FlDErrDVp7iSTw8vSz/l3wwdpLW5IEu4
CD7LA9CfCXwybhd1qpZq3h33zpMlrxDQhzYfkJZlJdUVOHZQ0lKfa809mjyU
NlQjtr8lApW6LUjM7kJ5vOhaN6lEhrlIVg0t+gtiY6zPra0jofH+yQMqSYl+
i7mAPP90K45OJgywlXkzV2/rc4Sf4gTH61kBZPDNZm6d0se4UPwwT4Z0BXYV
EWHqlv+FzFnWY1Y8Lu8LWh2Sb587CMudjQxZodxhN+sIbENptNVQgkRk/zIr
l60yTaNC0Yttef+s68ANresbC8WVeGllax3rtljo0Aj+7UdiZMNbLE5U2o1q
d/xRcRjzanz3OnV4aVeMnu0agfkpUPeElSJoiApGg2GkhFWDAZiTJMMWCga4
ojOjjwkh2DtIjKxX9+C4yRg2i2GQsL6GZLjY6uE1dqP8vbcW2DZdnv3Kgvx6
bcdhTZm0d4u2w7LzbK3YdN/kX7PJFIB76rSsSkhPbeassEkubSU7KUE1/kcf
JQvnTPo52XBMAgx3VPBN8O/n4Q/cTpjEPbAL7w2tLUFf6o74FwkL/g1Dki3J
W5Mu9s3nEBjNA5aiwB+0VBX5NdGHHaSwZNFQZ55CAPEHdYVyeWuh/vvzUl4v
D8umeVXq+F8SWjNuHSPGiPVuCJK9jun1gZE7rDsfpoIr6+5GGmxOtIII25oI
xVhD7XM+kx32QTPFIrPIo48BBLhYaXkhmZyodOMzhb6fuzl3PCo0bP1+49A+
dkKz9WTYh8U2Kw/BBvWYYUAWv4YSe/0f3dIDFHQeT866UaANcALMGoqjgbuY
eM4nyaeWuRFIpZJ8Y/KBqFU/0N+mUqCz9pCc24u6OOIxlrEAWhJStAKgw4ND
gMx8rNKga2zgxMtJd79X9AdE1l6UASEsVMAF0qHceZBL9ABO0SA2xxF3jT/y
QPTR2praR7k0IeTqgOAnOH1Sz/FczkkkG6M4gYNbTia88TSnFIECD3SVtW3E
NSD6acwYi1tYMz0OkvJgX+y7mMk/8qAvUHGOCaGcZUt2Sie7+RWdoKx9z7Rq
oJAw2LT1p0FI++ORuqw1muUza3Kv27p612H5wLREcFa9OH1TNuxMTABL/oam
owEPg/Pf2xISeL4exaWNwDGlwDbM34zVdGgqj3ZA2rmIQZv0maWL3CY9z174
GtuMacJgchmV7xg6s6AmDFKycQUtin/ljgoRS0icBGcAFijoVg0yij4k9dc6
EgmS2Vr5ZWt/pS1V/CZhOSWMrZJ5SxKEwq1sBuCFO+9XxeulLBE+4RQwemi9
dvq+i9Jk+0jEMelbMEsQ8z4uuBtrvvz5o56jgth21l7iJZJXwvxJC/4vve+j
i7OMXZqowgHRXugjUO0k0wsHJep+2gBRRGCD6cxKu4ok49lSWr+moZ/8NbPh
1/hcXkkG2JC8ed/9Kl5REJqQ4QT1HWIE+yrH0rpup0r9nAy7lEueiuL/Tlhk
cN9Nk6eXXITMQxayfoiiThQYHL1ZEvA2FKKhVptHvSuRvdHbwSf+ga6Hm6HN
5RUv7Jghbg/LjIAsbgxuJ3kNEhT76K4ir7tAaPM8DZKeanmLhG76c/E/Pvpq
gGemGLh4xFBYabCll+iiE5JYSRyjtjttc0MCWFxp3DmNIqtsP7M6trSlyCHS
/BiYTQzWfNa8X5aZ15l0kRfUCSXhe9lqo3rgI3oOltglJt54lN7iz9NmH8e9
+cY6bTY7Bjwj3/i+cH/zq/gsJJFk6aDBS6EocR+juV+FvrFAm+mqlqBjhdVz
ue67dYhdIgZSgTnT0txpehhyHW7acxPAun6RXDM13ihbCk+bKMWFmCl/Ysuu
pfKJVsFPZBg0U1kg6z0GJaZt5PceUmo4sxxoNTSeaSzjxieKJc6V9Ql8bxv7
KdXasojto1NimwoEuRkoeCE4VI0bU5DnKlrZUe5kTrKehjEL0Wm0vi5rkOp5
DJzwylftTYFFOEmPvP/kalhv92OBdwr6khNL6pPFZNGW9s8qqOO2UAYvQz1T
XkvpAyi9ubmCGjlmAzQtzmi+7XqCoKUmmrSxHzAWUmc6/+lDcRUqBIbznZd7
SGIFP8sKR/ObuIQJmo5bL1lmrkQg7j1ZL+H+HK5/y9AhkxhrFy3FFPomxBf2
rfIYz7OZ72DSN6sPbozkoqaAjFwTTlT5yLSzYSVNdKNoms0uCzWep6ue0qIo
DIz67pFMWlsD2fa623wvAFJGOSKvg6NEvQfcPqHUE3LBvfGpFsFdOpjulddW
AM2NdJdUj+KP4go3yB81cf61zRkFbKEcGaL2Ytuavtb81w6SIM7ODOsUbGem
oY1tF7rigrwTeKM1RILKy7cdGPxH8+8tQzMCQN7GDhHqzW7GOUbAv6INuESN
YNbmHAMWjAdZtrU3GiQvJfZgCw973SeiBfmXkGvIGG7j8UkjP9uyaW4J0Osb
0hzyLUcbyews4t/ElGVy+dVI/uOt+a/HE1EP2vIzeTNuHLvkYAwA1uA3VGh2
RtKIgQoSawAv1Yt71rWNeGJIQBRDUaMNKA8My+ZRMnclzvyr4LG4PGyuRzIk
D2K/M517X+bLG00EetgRUpVCKwn+n/+3otoAeJxNc0jU/XbndKQLc2k6QXgM
M0VClTVjfmLuVLYUQ5w+6afr+drfya2G5mJ05p/raJgTbekQe9XgKRSP5vCf
nZxtbWVqfsmzfq/5jx1VlFecxzvhd3VUzQFAVZmxGrXOuyDKidABZN+Tce/W
t1I8CbPMSMZf7dH+Cs28SIDKg12NThgVbtduYJC1JxBbIB+r0Y4mdyb5OW47
CBMImgtrSfYpLBlT3JEbNCq73j3YFF83C4F32tHiafsJ2WbMXUZA1xbpjk36
dEZNwIjS/B3o4vRu/8btol8jEGDz5319FbbeSXXtaceXixjmK3ZBpB6Kp8OO
pNlPWjKlR6TogjNRYGwR+7vU4yYdKU7aDJ3+Thgb4HmIcEy4Kpk0JoPm6v0y
QlAsctIaUCNMQ3RP0Ep3QeK/0wV6qnxG5CEw8ydRr7y7kXSWUolnrr/aNhHQ
V7XJsZR3igjOGITuSDYwBH7JM520x1LeV2JvUITy9wvc53wHPsCCpLSOPUbq
B0G+nN6Cl432SxA/wyJoQe3JHK2JeWq7SQa7nYHRFejb83oo6Y2ZUNpoGc8w
zlt0FtoJ9IsVVAXzjT2eHi6xvHYkLTpMphQ38XJwtCCBQS6bXFNpkB8Be7Wc
Xc1Wki0XdSeJ71mZQLW821vN5tLDsElb0yGqYAxcUX32i21eJmPdbzfFxj1e
WGRgdy+bm7N2WRhMtjPLEHuOLLYyu2cu5iOhZbIn2rUyRW81SNZza8eUJA3S
mhzpIYTdptJgbI50rk9DeTYfbM/VmRHAHBKoRcOWaWJRW8jhObI6OjaKD75d
vSv7K7DuVU1ToHgYrG1ohruwxjmHTFZdxl4MrInkOKPKa7HgkBlOzhnCq5z3
lAOYGbSAWXd6MUCkWh8VNBuDz5XKpamKQOkyzm/yLwFoIi63u7nBFF4mXIu5
XPFHv0f1FeK/8fe66KJJTcAe9DOLJXTwKa2aE2YsIYjTQHJFUQtinV7wq0bI
yjg922jcNLXI2AWEXumIdylmmVUcomc1ZFoQbdc9rf4xsVcTW9bw2dzx0dSh
pchTs2zzhFSA86VOA+KGiTWe7LnxJIhD8il2NMqx5beB3fTF6+R4YZv3ujRe
rU63MKJlGFdQbTjDuIpoppr9yjHMV0Fb+QddUAwvaDhkOnaItHkPs651lkTs
xL4wUB5X8Arl3IkXLhYnQ8XE3vt2IjYB25BwMgfsbV+yed3ZOsBRgb8WMIgV
4qV+rn0WEhpzqmL32/6kiu5OUmTtGowK16JrAp3FH/+922pD6AwkBlhk5GtF
buTVI8IBzJLX4VHXmwUsWmwjOHuM59Bqtjl8s8ASQgxy1fTnYayax+ASiyR4
RBeRSRUGClzwqoR/AoiGwBEl91modwUuTfbh9I54tUP3HmQ8mmwqR7r+6Lw1
4Pj/pVX81C407La8FPpNCpnvTfDCoU+TjDSJRwbIU8qbvwkEKyjz5XsC1QpS
AIXhAzDISUGfc4oxN7jEmi8A9vcm5cVbPbNOPICz8aU4YxXb55XTEimGRb8m
11pYNLy1E2OHOVXMd/BLNIvNmEz2SF2Afd4EtVmJV7Q/YSnzcy/U9YH5ejsy
UF7KApdt/zlkax6/NjELyT8oivyeVO4iYDVbjkwIrDlNuKTenTVF/rmaDYtz
Kgg/mI5q/2Bspr6a6qjP0H2O8IXewdFYTQKaBi2bIFEHcHPZBREBvsqFPp73
wyIgrSPvkSEksK/Xpc1nkv919k51ijJyztC07E25kdAJxOgzB5YCDUZRzriw
Z/BWmfcp5ooEQsMEAQ8OG4VeqvR+2s2inD/3D+NgcsyRSqAEspi0KWALQtXa
pEwNGSJ1CUyVI7J9Z7XE4sWsV2LESxGZwNloJ+Q4iCQDjMpf0vMvJqJ7KLSo
05JPOxn8fsXiq5tXSGafZ77Fn3oz0EihdkUDsERthz2rxfl2L8wlvqRuXKfS
9OprVc6k8rZ17E9NOqjfBzhm3l0LhcYfKbBE1c0XBXchtVB4ZZ1IrsfdG2Ve
zz1lwS/qaYazxyRqPYihFHgdBtYopyKCrq9dXzxSSX1tka42Q1qwD5sn53vh
0ZpE+f6IvAKauKtqJFYG0+OwGDMbmaDZi+M1u8rnDSrHCfRdZB/manLngvHD
OGghB56DQ7Yn2AGIEdBeUPnvud02EpdX0YInvdvZo+LwFrXlbOBzya3n4Ysb
sVEpzz31fQVWme/s48JMv1en1NxTMhhChu9bif2fmRZd55e89QlbCMPaH4bb
UP6Lr7axoAjQq5U6r3ZR4XNFQqdbLq56orpFJeEnZY7HBVZEOwp38EV/Y5UG
3v276bbK6zdzXD3eJ8rtVUsYNuccZPadkg0bmYoux6MO/2HUG9zOc+HKyIfK
XRNCdPvcDhPCcmGl7Z4aIfIfNg5lIoWTLDV9pIwNIYK6KrwwlSBkts4JosMu
VWx/IQ7wcstZhRKzVV+AwZvkwqQK6KmSSpQn557OyQY8EpT84fSygzScD2xb
FdictQ15rTddwUeYfKmM8nRCOFO9zz1lry7xh5PSarGx2YYEjEQLsolEpW38
VvqHeb2bMcJeSmZLlwrNKpVPZiQEMyYhps69oADqqNABBzR+W8eO1SlKVSX+
jUiSF3IFk5s3pTW1Af6KUgRXQNsNNQyjUD2ls4aJ1iI8C+7rJsItGcP07xtw
dQ2wVdsLtrUzGY4yl+t9SHHshNo+i8bQnRY9Wnp3XqJMHsiqQWJzMi4vAWMC
+Y9ngIluGsDfNPYmuv1Q3uSiZJvIPyihomqEZ7RBE1bM6FqtFPjyALG9Al5Z
OFfZgp1voAIs0tpa935vU+UDRYH8AJYD6QARWBgwVA4WqV37v6GFTNDLo2PX
KQqxft3GGuVcF8h66BxBopBY0A6t9TUB8xcWk/IKoUeE1yQa15/JvEmWBDda
zPPJJg+qg1JHK5Cstn9WD0H89lhIv99OIlEUxHxrdcfMgdWWH0WGhPEmm1ss
3A18PIUYLCMYmO5HKnG9cScxr6c8/JDvmsG1Sf9ZdGfyZybIEIZqfwnBmOMR
aI3qCw9oxCvugd/jI/gzX20sscKjB/9/vWe4E0qlcYzV1sMmD5ryV8p7j1hM
hLVhDDOAFswPhnXa9LC2fE5/8aCP+fZJ/1k3TCzmn6Chz9Vwvse7tW1a9dhc
cSCWoPVtBbAsLQC7hjdUzPY3IxPktRnrcU9gERd93v8zty2Su9xLWm+QVavv
A24M95RLg+9I3xLK5oRtHrvPHGlGZa5BB1SLLJtSKcXw3zeUKlgAdBGRcaJ7
ZM4BYKveYEK6FHOcHZTBf9TThl8WybGh179mmDOSnyb4+0BI7qVNUbm7QqBJ
dVLMM09tXs8la7Fjj/oeRRLBPE2BeIJBlS2GgWrRtGMBNencen7nEEusYY2p
BuoWuLL7B5R1kEy2n5MDHN2ZqikrirKLBPu32LfO8UTcgnbvwbBf339nLMhG
+mieOx1QGqC/Hr5IQ9uklqFfPv4cjcOwn+3ShNHrS3sQ2BX3PAVqZkPEBHp1
yIoB6XJvHeCKQK6NZC9Ve1v0z+18HEFv6IlUf08FbHWARysjRnrPO4KZHKd9
Oech4i20GEsKKG7U0dyz49POHx5rBgZGxO5RCgZL5m+uPZSqNBK6JWk0GDsb
3EV5JKL5pJDY/eTI5NiUwAWAS9at5isuXwItNbYWXvoJ2QPcaAuLxf/2EwAL
xgGVP4r+5231m26erohU/LxxWr5/s7olLOTibYLPVq4DQT6okQdu9G7hYW2C
+5hJI4yMkzS3nm8LI1FxMY+p6VbM5LvhnGqn/MLsfQLe3QpJXLiK7xBFYxZE
HHH+WdYpZYevZdYG6eemZku83OqfkpVJ2rP6rSPNRbYGj8wc06IjmOqndlXY
ATYwEzD1szMaEENsSh/dKigczLPQfEk6sNoniIVYMMuMygTuAshRJZ1HrqeQ
liJZgNKdbIMAbvyrYpg+Fnv8FYQGTYgVJ65ItyLFEWVzWJA/1Fauv+sUen2x
fngqc3+lPML0oOoknLIjIeRK4bI9cIPMP6uAMMvwF1D2QrPrPesoW+okDcan
3j5Uh1trwMTmcMby94RzcSVi/qfbqGA88SfjjJeYNhLwHb3CasVqtPGhWNAt
9oTem+70vlp+4C1eIeSWFfq9Tv5KEVC+xM53YEZUoN22GoM6FGf2qSC13SKe
t2EKLkHUubqHaDV44WiSC9r3Jzfkp9/5vpSfX0HpjjRaPoBr03L7fDZDKPvn
Bb6EgJ+H87MIjTRsIkdt8IXDtAB/scaomdXfsI4nqASCJHgptvQS/afOx/Er
5v+h5ahPJ0wkD33FWIIfUfXTO81cLzdKUZEPqMilY8ci/4A/Xufxr0QOEPWP
3ZdX1n/63486RUs36TndKNxNty6LF9TGiCP3mmAnhqBYzd3PRiXVMXbPA9RV
ko5ZnsHxqsIIDreCazP7Q+PSLuCgKW7UCxecssg4ScCMIYAaH9C5cBNgR/DM
nscEUB5jkSQ+wnOy4nSflw+woZAVAd0FuDj069o27Z7FdllJ43ONCtep1Vec
iQ9atUuxzsGxUlFrl0DpPxme7/mipkQiOQvKTBoV83br9alGYiO0SLO0hHmq
/f1kod/0PbxZkwMKLy9qksJbppip4V26wmwPyAWrQoe9xtoS3sNOmhcRI59e
xUZP+VW4Mwhjcs+AcU+InIUhwhXyl20KodLK9Yu+iM/awfLXulyrVXrSDTt8
9KexmCLypygkQkubf3WX9Sl5ndO/Bv3No3bJZn2PpC33wtAwZMhc1LblAZ/c
YYqUjzET3gl5RNJXfpEbWjlPXIkJU4we/53rNJMBOoPOumTBxG2dwbnCgoXx
VG3BaaitkiHIISjaxRyE52mHV0ev4vB5Fvfqx1CsfFvnu+qpjX7A/fvEOQNE
5LFlGSveT/jvFgncnAXcf9HncROtYSaXesP0BpsHG3mucrNWlUqSHArrvTnC
5AfadFGHz+O8xd4vwJfklCm5oiSi+rT0zFqrwivt/iSfM6/KIRr5JIl8FYEM
45l1piQHG4Xm0OYDFN3wuyE/3wO8+7QoF1Qc6n3bTq7gxPZPj4O75J86cxyr
u+rNNTsbx1MTcc3KFcM+xtkyULRnouqTL+y7S2Hke6aR+T/WhkhrW3oUz7dW
+EJ2Gj7Ub1L0A/YuyqhwtxhDAhmp4OZDd7Pdg9FgKSmIqgv1sR8de2hJOeAg
GTQzVE5PHvr7VMa2C1Fo6TZAWJL81PKlTyrgB6ygK3jlL6EMeIk7tBecDHSE
YFCxPT31rsSRICD5pz3j57CaZkyKXqBIqlVrJgjG7P9zYy982TF/CY+3eu/f
HTaEhEpD5e8qgKwNg2VQ9qS5lctR1A5VQRl8z+u6JoRBILSdy+uZcr/eKnuT
96WV8+qdI98GyRx8XFonQvwp9xU2QjpINUyCZv6lSmEZ3WhgU2+8zL8L2Kvp
AG0f2kgHpcPBzlttahHYu7W4ggOcO/MUzVCRz7EalsxLtQLZEiXZ2hZ4+3rL
uc23/X+EO9b+IiL1GnjiYCLDiqREi1uWRKD34vnyiPgIyiu5enDOYnHyhyc1
3Bc+hZ+xZSRNFINkH1BrlEPBbMtVEdfy8w2iU+7U0xzvFYqeztTOO791OfBY
EvG+czyDz4fHwUqrAYDSwkMHq5K/lN2jYnKyVCar5i2dHoCM2FTZFajc80iQ
dF1kYW3sr0bRhpHBi3g7L7D9Bf5Jh0PitwOLC2HWAT2OcTdxb/xuYPCaXibi
ZPoJ5IvpZDNNmSC1sOYb8t3RL0OBBFwRZLhq5stBVOiEYcHEgsVmD6LRFUjJ
GWzvuvDDPTy2W5pI5C1b2bitJVUJYtyYCvQv1UcSCh/5C2aYFLebY8aUsWSd
uSvXVG1ovOP0H8kDVp+f7BJR+RDtPDcpizl/wkGo3ZCrjx3ZNZDCatU+JxCF
ZKHtFumiIUKxhTji0qHdPQmjMxiH4LKc4Mp8XbxIEBTGqylzH15dG3+u25wp
3UprtCCZ68EnlkQayCD9ZiypT1ze/SjFdcG8+TQbbdSameQNCPAlpuNP8gJp
elIsp5SqemRwWGrwUE/MN9two/JUkLnvSC0SJmjR8G6Tjfx4YpwZyEB95vMr
nDr6xJ41f71UfO8U/zcZiEx8tEkAEJNWG4vyRCFeAqGKFUwZLNHgu0ebUHwR
Aum9jibWqFiEG3Z0R7V8hF6Q6IvsjZi9OD9/901Rut4vctl7Wn+tYaIOz6T4
a/9lj5smnL0tdolm8OWZrwNnpl8oyTvu/gA/N/Dom2KUb8H66RowvDvX037Y
TbXk0LdIQy/4pjumlg9NnAsiXio/os4ipW/QHjDTUxcThzgO68gUAgFFNa3S
oIviZiXJwMIieTo/e9SA4aTYBlXo/iYiAJMpkEIVfb7Dg/fq+3VnVDFoaEKB
XkXcSIo9PCVF+7zj+UJNZwIN50mubRvjhJZkKwW+WsLwX+uG7C++EBckcHYt
x+Iq4+N9g+Zwv20Pp50StqRgVInvvyGKJ/Bcd6EP7R6mZl2h3uZxYy/o3ZPt
iQKzpiT5qjYIiIHhfkTJZKqNeU557g96qgonFpPvMJxRotKc8M3PJilCWEGm
tZl774d3kVGmzO+HAuNEkncWUA8ZgKGXjiu113mch67bFZFL7txHaJJ00SSc
xnUwu6arZ+hzqSjCOJtrJNTkEZvYMtfLqB6JWKfN6AyuNCzAWWuyynFOmAap
1frVn6bTrgNJpFkYcayDQu2AAaVmp3prB1AmrCWMJQjcPu57rH1S7zKonCyU
hYwY4xKWxI0x4uL//6U0bQQCP1GKMRYMq+9XXUuDfyVCuN2QYcntw2WoU1yX
2rF6vQPzPDj1G3gd/n1YZgB1s56tnTAMJHfXohMwwuRL1Eqmdd58iH8sCdQO
qTCCBL+OHmBRsOwSj75nquKHkVwjhqWCUlU8qx4tzHNuhtbDW+kUm25FVvBu
/r0374npzsPe2bgh5BD/a60YFYE1G6izm70IuEE/bo0Y4sh+83NtaL21zN4d
qPkDc++7l7xuv4B3lt/mopjTvPAhruVco40njw0huVXkLPuOtEUzVQJvuCTn
fy7e/oq4CrfsDAJsz4ccYDI/c1tXGOaxqXogEp0P/MW2YCwA1rsyV998u1W4
rjB+xWn+alBhet10NvdBGPyC/sLb/hIg5StaZ2P+Zonk/5Fi4cBXT8JlaLzA
62nmaZxE4O1XNhZJbOMsV716jI5RvlehVjccVSWCzVEUTuBB2BywHy58vhVv
4Ntx/g3JB2osNUVBUwERD/ThNClzqA2Rui5hGhCUVZrIC5x5uTk9vVTuGLTB
i5XLoitmrnceHvAYuDgN0EHp2KUIIq1rGTtjGhzRlh5HCNggHdny8Ot9eRrB
ZpAhZgsJCbhrVb6swQp6IDCJzDMy1eDV/4N+BwWvyoSsGS8s4vuimRW3liDx
0kdeFromkXKvd8sIe1v7Guol76pRKidNnQWeqBW8SSGWbB97KFZq862ugR3/
IcEbIIILzATi2I1JLctauHCRQH7K8q9mO/kkGjO488v3rlt8pNU4p4xuH5QJ
llvX9106l3/is0z9sHb8UgFD3Pe0r+e/meYbwNmOHjrZ3kjwjT1GbWq4Ov1G
5K9WTh2TbyCInugsWQ+peu+cf2wgdAaE5EGpv6IivKR0ncHrjbPfNy2rdms9
TVsE+6QvJ8K7HUXvGoy39/zW2YKWM83q9vako+RCbIY0LmdzbB9m1gz/i1dr
Hmc0rXk1g769JAWFeooZTT/TAe+UFi9er+ov7Kekb7bWK5Fot0HdXlMBGSim
cB7RcvFFzDq+30SMfoU3qy9e3GTyu49NjHgU1kiEFZZN9uj1wsF8wskUtjdi
qBb9L6YA9NUUS3DuUGe6kgzkq/fEkV/DSSt9ywIk1Yvwg2vIEUCsND49WgUb
YExuwe+4vcGrGnk529Wsa11+a/sPe/LONZqUl9ynnU8H0FDv+Zv2cHtdGexd
kFKY/gokMYEwQYY78ImfojCJU/FrEZ3SvRBl3ADxP9fd1yuTrMlNpuk3J5OB
kUJ8+T7nQ2VpGrojOdzy3iGJ2Qo7+i0TM+bL2xt/9VMO0ov750L9iQyVe6IV
MpafbZpg0H5qQwp9TzDCgrmTREmTmCeyDnAR4mI0pMNBj/q5h5OMULJNNrmq
1KikTq/Sgp+yhd+cBnvNcdx8zMupNldUCDuJSGtoKaYIq1b1pkInnWd0SIoy
mygmUIrkE6gA/EhjVECg7+plvB68G7VFSXCI9CMl/O/yxuX6P/OjYXnwAoOO
/izWkdoaopaTodGRbM/9WiO37C6ucFq4edICtHHPU0ttjSfB0wJic4lUI3Xq
Zs2odOiColkkc+wayWhYrXnAXV0wX4DkoNrZW0KR/j1ByyZXrY7pfttpUeyF
Nckmx+qq+b4O5lGwkTESkYwxnpfbqZx4UPc/d6ozzgdAo+SELj7UiSPuhx5i
Qr9De6+k5/LTTDCUg+dzhTcGs/UmY78n1AhVSrHIjQ1gzdIezXB+kGkeaUr0
QNN9w0NIGqOtOUCCcyAvozJcGLUkqde03diTt4zTCyAlTAbT6I5wrxa29tRD
RgAqTLpNNIsw0p13dKvRe3hjwemcIKeHoMpZ1zvkTwM66d7GUg6ZNJHaJ9dn
JBzg4qub2sfxIt5nVkxQ6oVQHfNqxv+XuJYdlm6VzJdazIfcG2YhaJ6xt25g
uZd78ipf47qRL+7sl9hc92W0WE8oxVqgFCHdmtyanIAaJhJcylpz/xuK7+JS
jVTuFZHcx5M8ZztLQCiDP9JxxIdeuJeV5+Z3OH3aJq6kui8OlzPcjI7goBO9
N5hFsFfP+goIxQIBwAGUITOD0K7mENNMEsH90OOIVvaWo6KgeJrdYsUXBmxh
B/hMcIcbA1ES2N8/seQH8i8nqyfDCr/42KzSIKr1eGgHDgSK+sj22zS40jA5
hN2D+URbKdIDc727vv5daM1KzvK8d4wEmpox563BED3cnL79+gbt2IIWThSr
oyU8CMsync1E2UTUC4i9sQSSLYKEDVweWPexLE5OwTKzEAM7+GMVuvc82OVt
Pxt16Et/xXFLNa5XY6IReFlw5yHrPjdhdiBJxJgdl/HBPPFZc6ZICQfl9Vcd
MIhYq6rmVM6F0dwszbk7iMjjNZztFGZrGm6tsibx/J/90f5VobvWEKsSPVKO
fwuqjpU9b02EqfsCqteHsCsUCGidpW9JjBd0eqxk1vpk9DYESqs+mhgkoicv
SnKddFpQvaC5bazE7KzO/lpcwrjMh5HbZX6YZB9Zcu1LApTzrLTHqZadw7ZB
tYaXjoyI5vMLN7y+uJ13TGBXIyTmjEN7pzXplwF8g7x//nqhViwW+dycjVP+
jme8MIftN1NlBpeqO9uZMs/3x4dOqX/rA0HcrKQVoH3OHYDlBdjnvZsyt4g1
WSpWYkhLoyGMocTwEt0fqk2szetjRmKfjIvNKQvwRuBMYwy+pRyvpMDOyc8F
Nkk2ISJIzEmSCU2N+X6oIBGsTalGQ82zSzeHEfoRuExoe6ZxxsNtBayJRWMx
SelPWyt2p/nUw+hacmR6mooX97FD6i8nTrXkzTW9CntxOvVhvN91kixOVKcI
NLr0HGD8htkn2uHLy2Aq2w8xRB6BzqL2OPp4+bWLBjpO/LrKeEDGpzSChu7W
+K682b9HLdWwB6zlIMliY1wq6shuX4/g2EaO56gGgkkB1MtU0eVleqgZytiu
ykSISqEEzTf+Wwhgzd1xndy7ouWMnmPkew0UUvNuXhToHDVMMDDbM/eYtQ6d
zLCkCk+OqLHk6wKuBiiAn6KA3s1wjRzN8wn/FQcqF73nfwbHG6fR02K3cKdA
v7H60pCR2oIkbgrS3ORp0HqLsxfDs2WZoxzCxIrTU74IpYh87s2yi64QjzZF
wRxrejItaZHW7bBOcGRbtkPAYF3rSx6A8mB9iz3tF0bYsGYQY0kUQ/awIvZv
ceBGKb80SK/MRas7xA2AQ6QN7Ajq+6p4QnNOID+RpnzOqfH7nJC6gqupApav
gHXdXqj7snIVLR+28JZ+IHGJTR/iMLfE8x3CZFDC0QiCV7DlTtLqbAu5HTaZ
BV4uaFRzNAQl92NzF3bBVrzfAIHmhLeA7NBqAce4re/OMQ/8rsspspvgUo5u
LHJB4MmkdWhWfTkVQZ75nP1tqNA8Nv8FAIpHDUKC4PEN9cUhrkniYWb9Ovwn
A8CmRq8N6NgqGUqICqM51j3PLmyIWv9ORnnL7MlP6H9u8u9q6estJIYtW1B7
EqHu9Z3mPp7Zh726UeQaM1ftupWDFNiFKjH4K5RQ0QZuSmEEOzzF1YO1TBtV
xEoWgM8pIMZrUkyuz3QRBP3hAzTLWSt+IwHl5j+zESKUvkVhkz/pMmbmjhnA
kLasAPY5QrpxeUDtzxdBzNj4GwyGfkqx9B47/7u4YevzPdK4BVXtiGncrNel
ZEa8o9SNTxParn2DmfxSYxV+5ksTPMn8fkmPrJul6wR/SiAkqyaIzDP+xUsX
8f6o3ewR+aSry3gmHgmWBicZwlaqGsCpt2FwD1srXLBWwj0UpHUnA/zpaHlz
U7sBP0jl3BB06Eqjv9MUPXL0UixGrBGIlvkaja7dQPCg4NDtOUx9iu8iCf7P
MDfiiKrZ1VGE8XoTUTT+aMfx11IQpBJhUr2X6cNrn0fWccSQolXl0LNQsHyr
qqYEvOmEAK2OrqeGZkTFa3W/1ecosfkHrHoERQtDNaC0jDp+Rty8Y8VGE8jj
7zT8NIlYWjIonpgaHukhiSUIXKj7gMuqQCKr/Uj8fw2QGeS7+AymIb1G5/4N
0Qwf52tov5PxqZ/nVJuZQXUN72bK1tSld2eUrFerKq3HRA4xYtewuL2axOmF
wLJUwdm/mktnPNrbifWmWl/WHyrP/8HLBYx3VPNLIpe8BKYeTVUuLBA9zgRQ
qOzgXq6sjNsd5x3wVwCoa+pgg+8Iwl6lv+u3EVTCx+DKPv9PCXIY1onD3VPj
40Ob6Vdmz6bTVkIQgQANBaRd/7A0LkB3p4MTwQU8cR0WO0P2obW6hoqOLgGl
AZ4dB1HnVQjmZ1VjJv6XUHrgOQAp5UxkQ+y3muEcxeGmVX0bqNnK38Pxcv2c
qYkAl0AXdV/9B+H9a0J5jeGhap/MGQsRSGhrvL2z4kYBIP9y+kwQVPgSoaQ5
kOHi4NOF+BcgrZN9WX4nOVvQDLzs+pNNdeiwT9MAQRzjceSAiWbpGa4JAq4M
cxW0w0nz8568CysxqZazxbTPOBnBscC10MVp5H6GynOvUZFhOUoRVTaIvdmi
vtGK452jKctztsmZMyEnOeRPNwsiYsT2lbAODY4N7KBd/lz+7kvKoQ9Ri6BH
QPRaZigll2UnzVY+aQmxeSEpp/BdjUg7Z3CnzQB/b/DvdUdQigty/rKU7gob
rLqQtVjBbG7e0BNQgwIqdzAcqaBGr8/w1AhYuo3kWIB+N2OWlBc8x26PtyIz
MrpeaBzYRf3vaiLSPxHOXMjWPvX00BuKvi2mYH6Ta1YRhD0PiziRnyTqxjvI
PrNBJwWKJy4A9iHMnXPT48ZzLKhFkImerUxpoxfQenF3GK4BUcNeHKoqw7md
4xzatgLxapwolVXYfGPJ1ow0DDkIooOU9ggqCp0o8DkaoTF2h4jn0RYsmIMN
9yFE/Grguyumv16cCHCOu9XCpk6h0ux9/wnpGZ1g/NnLwKToc0E5UsUgr8gO
zW+WzfDSHW26aOhrE5OxIYcjJO8J9bvMiotiqg5P0YMJj+VytcaE5Arm0G1F
1TcNLFw/54O2jGOsOdXuoRojzCqNfS+KtwoQWf8UVFqhSDwKI4NPPp/1UTpj
Z1iiVV2DbHy9g4h5QLiokQe72u2BxA2woDznUR2XJeBvqNn2zn92tLNx4BSF
uXo9Ms+oJrz5EEZFG3QYCQiP6V5r8CQijhbNKzTmqxwkyFypaa9vQ9BKDG98
7EB577IiT7e0E7A/tkzt+3Ggvwpm8u8Goj4d9lt6ajRCRzMTupt7wsdzxeoA
gwBE0G8DVCIrtsEvoTKSjDABFAEG8VzWFzkugdV79YOqcQmV2XFfY+MzfpdW
H5WOfiO7On5TKf+Jj3xIWY2nlGZKekherT5saaJhrkLa2VGq/KLAV8/V2TK2
WXvsv3pMfeuG5CpaTY8PWdPnx1hYAo5ei+fUEk5HCaS5rWbcaBR8z9ww5tui
Z7ydgBDSyZyEBpR+GgHavkXQS4zZh+m50pnLPjP6J39hI3tGTP9eD9HDj3es
GkliPOo3TaqCcJD1dpuc2mlEZnUfc3+USJ50SUQLdiv5QVth8H/OW544WHwB
tNI7Q1A6JDcnHjTEYVxtW4Y1Y83auXskrPagPzTTBayXk5GJXtqFHmimdvZB
Q+T7RPluAXvoS2JbZlPFtWCAnE45cpHO6sa/kggoKAdUvfSnthcb3atk0Gxs
PSk9CLBEr62XVY7BHhuRLSuh1jJfhYoH6kg95Uh3YHtHl49RRtggQicnfC4v
eOsSq8uu6WuaaGIO9Y0yKhpShwBcvBh5WWxjd2Q9t60gjsAecMd8V3+07cp2
VJ7aCjVGJwduRw2SehdsoNBLbXDN+FI15/yvLr7752ooMrX7m0NpDUvYxL+L
3OIjnXs2EJ0YeCvW2DRsXffuhZTHIAKBRwPlapnFpUB0NMrvswWmsx3TV4cy
/KlPBZbtMa2g7DhWNn3SSy1510nx28pFJA8uWMoJ4N7gvq7OAVXP+reyArpr
Us6wb+p+JbHYtLIscaNO/OodK4g+i9nSA3lc9Fjkm6GnoatAYBc5a25biHvh
DxDKrz8tDvMTkeyccBGf8cqwtz26zU4n0GZUdjQtjeyZNG40fRD0eG47boGJ
yNN9/ZLjC8kmPXVq9xW0sFFlG7sjLU6RNorZIIt+1eabam+usuEQSoqU/MEI
/5vDoK/b5DHg39LU9BBg5DWIkWVmx/NZz5wwdM8ncJaDAmJDp5nLpaNIr1oK
kbKIf+GPSCXEAplQuMaEYNf9kG1MEff7t13DeOud6FkBx6hdUPzMJbMOlomO
ATvqhfi0dlYuEtVUztT/JxdVubM/QDa3Hq4kJT+HZ0JaOTHnJJLNbDxs8kha
sCQBJiVtFlKKG4DpRAJFR+0tHDBp8LLw3+1urtBvuFvYC37yscYxMzoNE/rN
VNvdikGNe8JHc8qBx21l2rU56/vEv3a7hs+OhYC7E0LAHAAczeyN+1ia6xSE
xGk/JvXmwv0Alzx8KxwWlyEZYQ/9mqVRh6GvbZ44UYL0aYHausnWmd7hng2U
v1L+Iniu3uboYSnhNnoNftpWWfTsV39tFhx4Z26RaT+y9xGg22/pB0IuCadT
eMy8zNOT1n+knfhkalyK96UMvzYpZSjZDswr4oD/aY25jT23X3RW+xM5W+9l
OsIR1mmCzYptvtc0JYfGaH6MyDF1K+2eiaoXrxQTGWkHfGbAxMcoGA5bD5c4
PDN3O1QEL3tN8TCgqhq+PzPhx3cH71XcU0aPptDnhSgQeFYPGyIXD/3YS3Zg
dAizE9c75eH3C13VM3d3VVvaORlzwMhhjy36yEo/ki9zbhdQQ4jflX5SkBRH
6WloigvZ2kmlABiLQ9QWl4cfGstzMvPEz96P2TUO13tq5HQKQAdZGEz0bagv
e7DqkUAxV/scPFZKlehMgJhd9mJTbv/YJzyhRVaffb5fh7wJNW8bThv4/5Fc
85Vlm4XVhQCVyckmynuLIujtF8eSQFRqiGTpIO5YykSTB+I35H774+pzJ48I
dPFo0Jh+K6j0ZeL400Ny5rIVp6L43vbGoTcYhsobn9PvKc2182eh3GNxr1DQ
CwHHMlOIXQ6WLVLePgx8R9FJZ3f9I+6EzAknnbsU0EfGwaGrISON/Y3Qo12M
RkCYq1KISZQKCV3L5D88Fy4aTSfyrn7m5E9lorba1kosM+9a1fTLQ2lskVZT
vZN6phoD4Vja5xTVKie4wdUMUdgc1XKsuAoWtafWxjK9OOjPMGSrJXBIeOm9
Xyqeymh6kOMiaPTE0ASgi7lREFaX6MaGz1oiZGsAm3PoA/4sUpsmqwmM/Pcy
JjNhMIICTftPK+mx7z+GyLE1oxyvw8udjCK9zpzOZlXhPrMs/NnD29AYXnv4
ihXp8JbXF3umgp2Ot1eN6bT8H5VA/0mS01833DRq+xsh2zwImCtyIwEyBeNL
W49cW8w77f1HVaFbW3rGy1vpsvhmNSDuE20S6SRVdY2cM2NADlWC9ro6xe/6
hQTLPtJT4gL+BBUbt1Ob4oGGhWB0ywpDeQ2VYDrR2V/M4hEw+Z4CQcZE5DIo
XYmCxo8HBGIDs0udzQuLUmMrRqgHbIjdiAAqYOJ4beoewTciucclSDWaDg8t
jjdnVnJfop+Lgn6Elgx14v6xz4zRaHkZVYZg+qYC/AkuOdiTu5Bk32Uuu0p5
XcdGVGiN1n/Yfq20sYOJxA5Z4rKss6w/S4mc/Auo8X8/UXqzYS3CAZN4KnL5
y7uyF/M0AaqSzuNWEJgj1zqOyrjmv/GV0aZ7EwhAhL95Gf+e715dGnabiScg
mBFtUH29RIVvyS/uc3Ko0OKf81+1k33QxymccrBh3xdd/TrzvIVBZrRYTUp9
/Gt6MhW/q074Fhir1EbGW0Mmt3tiCKvcvTYZ0Zb2hHaK3D4SsYnGRjirh48T
tjJ/oMevgXr8FmEq9SDGxSF5H74vOyQ8zS3ilYwmQPf8TUrFxXYwyP1h/qVQ
inZPfrnLqtcH+lD9mhThQkdazjuk1abuq3U76FHhcfOWtMRHysCz8IF/RfAr
QK3JfWxoY3pVeUeUNdrgu01s6oiKbw4pgu3H6/kbx9hhFxEYWGVqP+VOu26+
SXZe4abZwr7dPrDv6tmvVU1VAMQbWvj5SueL8ZEQZJUMdEXEGShfljG78aQI
4GoxyJhyQmwS4epW1KOdmUhGmLQ4x2mhUXPlzBumnTvw7k3KZl/XdQQA1c5i
lztqbcPAPMmp8OEcT1OhHMZ6jS9Um5QYaLPWQQB2MSZyNIfuCQjKaoSPDRPO
bxRemAdb+v9zOD8hdbbvuJ++1umdCuWOUOyw2zlpZXtvBa4M2u0y/YNePQDE
G3I9gqu4tPsmNbyFFnn0dNSzUJt7+a9SeJW0SzXoaaMkciKJRJlhKFJB2Izh
1E24I3jDF7MTf7k2iGGFSpBjo5tIPh+XrCZmT2TvyTwD/PWRU2xfkmnn4epI
VBQDh3KqNr5TXm5iq0IXWlIVt1Ik4JuTA5m7oRZZEK+suSBFyqKN5P9NMJaT
a7Fup3zJwJ8e4ZG+TliKO/pkm6RK1f1sci9hQ78/ZG5FQyhxf59Sif3FeT6U
ENQEQbVrf0RUpRbuDRJW3GOWAgf2Hgdyf6Jp9QIUQWKeg+1At3JyXNVtwnbH
hZJxQw7O5fm4u/VfbagA/cxuS2kS1hBmS2gMAM3xagKJFkLPnG6DeYagzm/N
30p8GQBl24JBy4rkgR1lBlQOkzTaBWnMCqLkE63AF4+Zpzd+itnUarB/8KKz
4zbXx1H4sXA1OvI50b3GyfDL6mYlGrImvaS3Z/HKQUaxClHbX/hfs1x5xKoq
TuM2HFZyy2abJv4+GpC4+foOBVwL7G3w78t55+WSp6CuJylNDaw2Nvg220K3
+DwNZFgtEkkSmhtPz+Yd7F76KOifWX96DPQcNA1Wp3XKh6EU8T+N2Q76LiAt
pmWUSkjbIo3jCeiy8dkI4SO1ZSr2wkUf+CboSKhbT4BljNaO4bieIGG3XFw8
7Npu3grpLpi7RwoQn1K7/gfu44Yhb4OobkYY6WixwYndAJ+MucNqhSSmKzvK
fSJL96Qg+EozaVKjPygepKASqGa7CIoEravN+3msYkjAjN39YfAUjo6e8j9P
gI89ZgYKyiX+v46GKzFJNgCmT504tCuSd0Cps7xsj27K8CfmCCdg+xRgAjp0
RfNnXNcr3yRGe4DrE1Kpa8klrVWc7DTAfFSn82b13RTBJY2K6LrRmLB0Wsqx
cOSe6BCw3ck+nu77Kne6LaCnL0xd2B9g9paE4PjAy0GzsqmjoiSyHeU+CSvs
83UDmR7S6MOjw2zsxwi5zVPcw0aTUtz8k27/mhK3XLEdZBrk/rhJDyL8OYMq
HS8beL9j9AmBsL/WlmmjM13H0wwmhK53FG67LolAwiOZv4M+DwzNqqQ6ALR9
PcarzzeIX9IMSN/9+YaAJpCnF+U07dLDr+3ojQOeg+sd/4F5biqeB0MelPMx
BU1i+zNYSBYZYimI3TvWRqF9tD4or1smhDx8zrVmG3UkabyBZvG+u70RIk42
UqOcvvmj4QZvAxJqHow0XswKMGDOougJfqsoHKE4SNDpyMzpdlgYolv+O1eq
q7WBviFaLdxXDhfLQYRK2DUfsXyXFhlmIm0c6FpeJnKACGJEfd6mrL8G1SxT
O9QAibWwuFgF6V6N4vdNI5i9SeW82A/XahYJ+46M67La0i8uWNd9IqbQJbsg
27J3VTCd19eAezJON+rK6CdtsEScX5U9xd18ZU5liQsoAMjBg8MLj/gM9azb
s65qbJQm+OD0xG3mN9JzuuNIWvu0RVSA8rkzJGZOoYrS5cl/vCsnhoQcCYu4
+4Bw6A/gCMNzVaS+rUlRfRxAmQB/7XYAk5xQIjLjbsSNYewPgxp6Rj8l8BZd
QE/48tyr4ge+Un2Sdj1NC4JOPEuFrVmNIJIdEabOzRnog8ybeRAERQBaLZRO
JR9NhXOvJiJswLBGkzBEKUoysu2oUt1rj6lXmTDXSeAwG++T5H7/ETgLKhdC
qQ0QNIqA7ARJGN17RULOoDrkt8VelcMT84dylDgTIzFNwxiL/2c0xc315H8+
SIk+L8kifSNS+B6RKMf3MAhixeNSh+PTnoN+GEQPh8tjH6yAQiLaW5quqXsi
Ktp75j+NdZH/0SNkSLPWXOfjmdt/cglLQWjRg8oNzVxY1CIgcCCcpBBPnyQQ
XGze2AwhZpnMM+7/XNA3dObO/yBKagCu/Fwy1qSmlBCkXvodlCLh90DXiHnw
ewc2yt0KggPC1zxXBZtCNamjGFBzbVSjPv2scvSA4PG4Arw2R8tZeF+GpQDd
dGjU+tSUbiZNaL2qJ6MM0zgPdyNidlSocrdV++39XZxPgyHZRmtEvH8n8gWx
f3YrMBiHqsHs6kS5np0DvEylGo9tUWfdSkL0nMGcgKRv3nMXg8C/gxX6CarL
NjbNIclgsNl2ihqQJEY7NXOHBAyiwwG+KXLQKGFRaL8HaLgjtlXbKQ5gais1
pHBZE7PFTgPke74tSWBFJASJeMc+UsV6SZI2BcYPbnST8IuuFcjWXSNs5eRR
3UqpH+6crH5qyjYh8Lq6PIjJIYBbJlpN5dZ/T89bRAmk5Vbfh8jFE2b9ww21
gfAiPEEo3HVRF1vIeodyTED2515/dkqsd4HY8LPj3J4BSfWmiogaftgNxbxF
pixCI+q78p9+KjV2oTvxgPWCR/E47cXvUGwKkUwRIyXwa48WqZj8E2phTeKl
w8ktrBdOIhFd3lESlc8RZhS0p8bfcPexZDoaPcl3qtlxYFGAKdj+85IuJ3MR
AfH8ohOusuPnBpYOVb0+5GLizlmukzQ9FIZSGrmlW2tkLPE6YvGka40Exg/o
QFJ+nwEtQEIHKl5KDPRxe6tFMxMChsrjaZxRPqEng484AAOE7mpZU0biaUmQ
3Un7/ZskWh8FWPYQ9zgEIG195XxoyvISnSxdNc2WxZIVnnldgkohKlkEgws4
SiPq+pTOre9qWnVgpKF95N2yemZdN2PYCqfU+QKlMP2bos5qxLbhyJFlUOts
yqIafB4wurWaBEbQ2g3G7MdckcXAeLgm+0f/q1iZxLKmG7EcbIjrodNRqGhr
MXrOY1y40r+Gd8QU//Xh8eFlxCd7QQZMy4z/NGhsJAJFp8Ei5FCSAxNkYN6b
LQvb+wSnKQDeIRUCQOsdN2hl1UPDFKEZumrkiIWe7msh/d8v1Sm028zO9ava
PNIQOqgvu4lujco6xUc/O4NgHkGgC04x9bfj3wFQjryI9iQVuktepZ6Dxoyc
8OdRsuZfq2KMF6+PEREMKA/v7VHtcOvZmE8kHDp7uz+QDkWrmyBYY5XjHypW
ZVAKaHGzVW8GpbyAOHkch/lRXAZNk8OdKedqYZfSjhUCDgTTVbAaDyIOGHLD
f2ct9XqXQyPOXnQUbhTYfOC9QnGvBHj7AVV68RiXgYPDALGRwDLt2NfqYZ/E
GadnMYKsOuPWDBJrMjveHD2kp8NtTRzhNvRfpQqy9IehZFkuwcRgDdaFtX/A
0w6vTt+ggRFjrUgn/Samm0+qL0svT/KBavDwntsg4Jk+Gfism5my09DNHHuN
80LVvvdBFYHeyFAUAvCvb8I7MPed82lKjSZQxCwfOv7OVSlzbwPZxrgomtDG
eVw2Js6xiBp95WfM+iR8gDl+0ysLtYQN+fHIhiLToKNmPZO3xTomuctq5nug
vYHlky9edRx1tlGBt6/ANEuQMlGa/nV0OxQbAzcwTsbD9N6XxUUaUk+K/iok
SYi2QVoMbHQEsEMmjo5pT/V5Zg13rza74eB8mo/6Mi1s/n8uZB6I8WMasr0Z
XtP0gn6J9cNS00XTmjsdZs8Af0Ghiz1JS/+7mB5LUY2w3EtP88gpByIOrEN7
XdtjjGqXbTYAa31TRTKCRGl9DkfZC6bpQmtjk5stuKMOor69cDs3LSKcEeOJ
QCu0tcr8jxBtAWPsC0B3maL2Cg/kYcy7xEC+wit+k5lD8wv18SjTIY/NL80S
cSL6rC4lmTcYcG13y6eA1W0bclrDsWK5gbaCNhNxy8+1qVmYOXy5XfLuabrd
AubEXrTImvXIG+/KnOCRs87kJvBFCbzkacTyWj6e/emcmhHIja9X6iqOBcKG
aCa0bTa9G6DZW/zCaggiPnmHv2C/xgHi8kyPRAQjiaoniCO0o9KqV6WAxHw4
x0RUkpO22NMYsBTkGM6OwvcAH0hXgEN5YPy72EW3puQEmWQRkS8vy2+knrM+
cTg7dTONVugldayDJAzx5wfkp24PXUcB67XS7Kifpp16NccsM0ZBKi6KtzXy
lXR6P+UOvDDegUCEDJ8e+FQ2M8SnKH/5ou14cGBEje0/9UWPNwo+xa7K0UVj
1Xr1LOfsVNjVPqePakqtVSjXApiye2+AhGUxJOFPgVQSxP2WlHh1QNHmRgew
2/hmKf1UNfMMPt/zrxqsWdfUcL/O86B9Pr0mH8K+QJD0eSuwfSlXXdUaAzxS
XNDKPRZQDDzb1aWvWsVaNWtD9UxP3BWxM8/mpLIXxGNEY4gtxy2n73SVwSpV
OtMDfbDwd70MUmLHtEaTZPw94PMZNofGgtqkOTH2ciqQVVa/Cf2rM+BWP5Wk
z0T3BqBLpkSoGxhKy5gyozwMWQYby1KENKZhHXcmo453iwl8dhk7Lg5Uktyc
OmOB7zmujk/NmDSD/zR9f0Cl91aGNbZV4fTyQKp1LVQkUzKkPwIC735dMOD/
tOG/fjdrqwz57uyBB30fQRzpoWwljKSBgaKvApUGDjutMDqbupy9WjY+LCOi
q+rJ1hH18UdkfKupHO51MfruJrA1XRC80xfQSrtKmjLpQ6IzV9mcDBYKR/LB
m7VYPEuYvhOouuGCmBMxjod0pQe6y6xfkG9FzQ+d1r6bCPU1uJ9qeNSkwD0h
r/zcgk0YZs5g0YDvmSGoZODf/RTH4VDOdsq0n1vrZIr1FIqxWCbpsHJsUIwe
s9B5OEIvStMJMCUwkWNOD7lLNq+KozPczOHQ//gLp92zYRtlz7rxwtDaYHTd
Oeb48hdL0Kr7RIXJVqSBlfri7X6dZXc7SEqeAgu2hCnWUFVhgLB02Xi7DYZk
8FSjYiwkF1CMh4ugBBCt2ku8G3kLQglotdudF7UTHkpP0/XdpGAgTSAa2slG
uFpzFTA3OWrvygtEJkccu+HtIJb+YY0UJd/FT5P9mmcWnW8k37xmp853DNBq
fcFxMjfvGBpNzRqi+3l2XvyK24Mk/MwrDSAorp7eq6d5HIVjuertNHOlw5m6
rqN4sGuaJF7in8CU3EiAALIbjWxGmxlhvAZNM+VMYEWpvhzeCff1emhbRGy0
eyOM50yLfBfImuWHeAvlGQbGor8MmEafGzFBi6E4UMd74f2G1QP1nPmGyc5l
+vzgTveDvjec+jMnFWpp+T6vIO9PfwzwKnXO+n3urrlLNyS6F/dbWTKxHJiX
14Nwr4y7TQpAVyuwYKr2h+pP9Y03uVYrxFHadFvjaZqzze+4tWFCU6gCT125
V5immG5w9PP2zkstJ7iMzIxHzlsMB47ekli7zxzl54rpOa8PDKdJUP40pLOb
paD3C952sG20e9xg2nZ8tD71gzwxGJpMkB1EmZKN2wR9mQxgGFgnvKg9CipU
gPXeE4hcAION1U/w7HMlAq/019tb+MntwtT89Q3OOHcsMwFQhRP5fCnAgjZC
80LQoBYrAw0y0vMTo7fqFYXvcI9PaAN6Nlqf00saLilRE2L/TisZG+xpCt6z
HVHxkCNALQPnHFklXybp8DakdaqdvLQtnaYUPAQhTzY9djE5asSb9BKEWdHE
PnuKjJqiru2fphJ1TnqkZhRUUY0iKwLhU6YkjhykDBUreuNEwZ7X6rjfttph
+azC057JazutQUOW9jByAh3kOPh2Xr0P225GPCeihfvZoMxaotFaWNF2DzFA
LyFzTM8XSwFrNm3ceDniMHubyoaybFadCkcplvSGDRLjyLkRj3tkjexHuK9I
H/r2xAXN5kukELBlYKBptYCzsXZUGqOC12peMXbmT4qVVPtoLbJy8BR9Dmjw
8h5kW90orPR+QQLJp6we9qMiOPSIpiEz/wz/i558ls1l3irLMd7Q+UxCtzJ1
bJ3/ZiUoOodMSnYVJKjp9caaIvNrTahWB03QmbzYP8lZLbIRJawN6mtS7FRY
uSJY8W3ScW5SaY29HavY15ocil8VsyL+Jt8UwR/ui2//IZVlbvk4Wa0pg73f
pVvFzSKuJwBbmgJCyTudtOg+5qk/NPuNMpwI/3x0owCPIGzgYizeni9YNuzP
mo40etoP+Rpd8JGNzxFTVCeJ2OhqnRx9oA6mnPMc8SiBHdfL/Sc4CnzHFMMw
eCgDyUet6Rh7u7aXzjnUKhEXdiNESb4m95ajr+nTMPAnyh7YzB2+xQ/yZzmp
mjCQfq6W2OAvShKbk0Uu2IM63R1fMxdpVo6ZGFjMfeF/oL2tAzVx9aN/selL
ZMuHAP9gwqubNK6xOzRtzTBIJ+Z7JluFuWQHcxgXSwskS0g7dLfPdD7agaxC
KqevIaGsWsB2HCFxmIvmsHIzFGo70soUj6/xydvQ4ckLFiCCrnKwQC6KZtCc
zaZxM495cW9x8JfzYVsOdL8AqFT3E2dMRpSDnUAfOkkNVDlcYB+64qr34Kg8
1KbQMOxaKQiTY9t2ZZKzSuqqdhn2ADIZ4T8ieMX5qv4qGqhCUOfLoLO9F1ei
8DwDLSeskoi8xstoJkcVzrqixhxDc86m20H+b3xFj0+qNHBr8XVqroaDO3S6
ZnkF2h6yYhxic5pmbUOZXPclzKNvmeetorbPFJyc9KYDP+pUlU6bMxCzEuqa
8S8cvlEisJZhM3YFp4+Ui34hPzNc1nqaPZ1N6/g4siAEWChe//5BoLMAXWWO
IZEoGma715vqrAoHp0vYXhXexckCfh6/mo4xIK6zZAd7VvmE9pyDBDEnZCjN
MgRNaG8OM4eSQaS2ERIIHASconJZxZbrInslasX1f1Dr8RS6c5JzdbbQfKmh
+wKW6VYtc1JwTEbcbyX+2aXkCuqwk5Rc6OPUZxUkcGoUQw3pXD6gbbFYFcHo
sfHDzxZXN/sXckxIFiy2NCjTIgGu3CnAwhiyjYaZopHB5tOdWRXKSUwngnhk
E20sbk7Sd3sRCBJmgq59hPOEdxvIWIIC+xDeeg7khEi1IqrnqwfOMTVNFI1P
BvQqYNM+AO41KgkJmEYaNzkaSLis9dJnmbEg30JUOKohR+lKX3tUZqwx2m4G
7LSswbh9UOFYVdTD5f7UYkrvYpYxOnqW/r3SCEOV2NXPyjvSKWOQkDsJEOUb
EKUOSJv5sZ1Jd6er5b9DPj/hxaq+teUqcYAlEcdDp8bT3E5ts2Zh+KhueyrW
7njmsxRFRp9oNBDeDtAYmttx/oKWMQXXJwTEfzeBKsxlO2lI5i/4H4ddbk/w
OBh4SiUkhQ7dNz4Vl6xhI88PklfoNYJPlA9OV1HSbUxacDo2/4NnikeS+SnG
iozaJ8vywmZZz86/ePOt1r9eW+UQ7o6PuAxxbTe5bJg0AjAHMdc7ePdp8wcu
n+dkOSTY9DmLK3bgkzKn8Q3IykyX/9zuh7sMNxCg8HEO9WtaUOTeuHCoNPQP
CCmkcQKV3O4UJBlC+4V2wxIxnbZzOAei2h3rD+rSai3bv7O53koDr6iN1uJa
IDIkdwHml3yz52Anu8TTihWDi7iFZ1RUf6ESgEgR7/cp5ziI935pt1Y58cHJ
T1RsX/2C1/k9MrGVLzIPxmfczC4N0XR0tv7YOx6eh/W5t71zrtAPraoh4HBv
94Y/w39uiTIUYezOB9ME15nBz4IGpYI5J3dhQ54pnf5CFw1/bkmxPXA7ySw/
X+S2Ci8gw39PSqGETFRkSKXoskNanwn2NMfDUzY6TMFNf6yiPgufSN/momfo
8fT7hAw+sy+fo70TN5EkvLD0Lw41Y/zGxPT7EMa8mZbsFvuc2Q3SsftHnqYX
ZxfmwEiw7/3/ZoMVLsjmu3q3GCVTDLCFbgizi7MsJ1euhkJcC/xsqdWJ92E4
bqfeHiBDms8mmmSRW0acL3ERa74FL0j7CgmudOgZrjGgGs42SfIWQ7ry1CRm
o44sCsmV0XwIBEge2pAAcFFXH1l+qhQfuzKPkL48gyr+l86LuLcsktym7JuZ
a4716N4y8I5iRKtZxYtmPYYBOmLOqTZbpSQ69gtq/W1XxnD3Hmv0P8JawLFE
sGYhOcFJg4uRaeD/D2D9AwjiINncLG2Wki91gs4yFYvqMh9g2Ds52S5kIxcD
bP6N4NZqsNCVvOYfJ42vKPwBqRkgz1EzVhdxqEVF+RLdPRe/rKjWwFIMglu1
4gS571csaDe/1KEb46s3kN3dpSJJig7eTBdCHG7w9dYPiV/4bTPt+2noNEwJ
3oPpeN853uqi4FjMJ//avYZIotrqfXpYUO6zLOFnUbYttwmX6UYoYQSn0un8
cht5jHRyoA09EHSu13vERdCWoSEjcUgXoLe1M7f+ERbytRcwtQH2DxLHvxZ/
nyRp6P+/35+qBvOGZxbD3e/Zw7f2S63ZTJWYxIOHfakfQo/lmBRI8ImHVaGN
INn5Qxg6zIyNhedFv7yaXfarG2Jp8vVA5nAHhYWfoa4NLto2gP9oFejzWzU+
9qTBJgpOi26OtWLQpZzACqCVcQ63A/cWbbG4zadMnknME/mY5cM5XvughLWq
MraEcKXJZsPh1zl2nGCMOkJEssZo9Pi/230mf/uPq5AymAOWVXx0c/Q42IV+
s8PtcbZC2eYMXWZVLofIifQJgJ00wprWA98H9waJ126f3CzV2DgF1juD6vtB
GH4Uzj0CiVDKImblPs3I+4fCVfjLJhBxbkYV7xEU/mcVzNqQH69/REwYFmBm
RXeeP1XyAIfLoI12XthA+9hML6xQVWnZYE5oE+awcpdpwB/+6CJdRPQD/Zmg
0sVoQbfVM2GIqUtfUsZr0v1s3SFpvVklNRSvuKUGfmSYDb79eF2wAyMJHs5z
WWaMtr+qXW7zgfgXLnuEpCGxSq4xFn8CHFnzIZVyGidnFcasl4j9nJb2m/Mu
KjfmLRdhm2+QATvyLCi2HjJoj6Azcl9iPCyRI0oxm096JPRvP9Nfza7EP3yj
Ix5JEobkxA7c1mvWRGkbHeBglgQhOwZOkn5ibDXvajMHO64UJC82rk5PjMg/
+3NdCeEQHcWp2G63GhK5PWiM8JwAuwAFFIMdFmS9YGMhtqeXVeY+B7xSFka1
R/VWrHuqE3W2ao42XVNLcB5hR4amBfPLSPEadtA/Zq8Q0Inhg9x0JFiFbPrU
A5KZie2oFeKf9qKLJl9o4GwcEy136sL6BR91+47MUYUeZa8ikitY0L+UyXvZ
pstGix6LPbnoWszhKGxNEda/uJu84NbWq8Qea1BMfhxEdVcfZu8x8EBPSQSN
b2ZOzS0XdzhQoHvaqz8MU7+IOl5/+QDEf6ESVdaaf7QlOs54/tAoE7yC5KXi
C1vUlt5+zPMl6SNMcnXIkCPSxkfH7DjCX/VshyGX0nGgeqOj+/Z6RPjYgyVX
5jMr3i2fwtMGprW0eudB+5HkXrd3zdESHeHzX+FSOXquuB7MlqW5wTAUd4Bb
OvmnhFYKqPWPi3glXDXhMDDI4reKMPfVVUT2c7d7KaPTConCjnBQDHPjAKuR
vzO+xKj0CrR9RBEatLfDSR3iCIPxA7woDX6J5MmJRaFMl0jHR6T7/Xb54DuX
FXyY+bGvIopNHemubDVstvw5WgNdUK1cUy48LZFCL9Dkws70xbTUy8vADPVj
+qG9mGOiuOlviTojuZ5P4gwVt3/Ve4dn0Btr08ZXve1kxaG0XdOIpAI4P1Nt
0XLshnjVcu4tuQoc31pPCVw1pTDJpltdfdLxqq1zLRw65PRe+ZQx013d4JwJ
7o30B4E3k7Bxgh6+WMPqVlXlk5yAklph29uZUZyd3WQSMUf3WJIXd4wvmAQ/
3lJdNsnAop2oIq+usPAsjyiHES6Bwm4kxGSpt9huVGnEhtdffo/6R+vGyfnJ
W/5mcYw2I+8CDplq3eD8O/60s38EjLMX50tu4XFcL7PRi7lMZGblSYVkuINJ
wwLBZYw1jAgF5YMsswufgkxx1DvAATH3YVv9nOGe5hKJIQbF3rrGjW3TaZgQ
CwY2tekfmh3wAe9/b/A8oXouNRrWhSyfaaeWOdfJI9Y0Hm/qG5ogfKM+EjaX
FYBLa+Co28diUzyrpvohHqR0nUUcQEnNkgqobETfpg+wYlNTIzsYfFR4bw7a
qIw7WDC3CMX2rj89tqH0pAVg7mnaLqU1PhMgP6Ijy5RM8RXsFMmRRFd2/Pfi
FPRaPtGsWI1Idr7Wblz55RBw0Sp+nISORmOBjAuOG4agZFgYt9RbkgUs+ahC
AVYISdPjgY/wfBrUm0ZLBhC3XPR2gLmpisfcD4MUg6/2IwUZRRvErvyQkwFO
VKoQ4jrUCNTsUcBuN0p+47QzPWmtS5hRfvxNtkiXkKOdNlGRRtwRli+sx0Cs
mbr4c7WhWm9mDtuwz5me2roPCV4nFfp8Wd3GbmUZjRCsdVrPcYyXPCfMnBOa
xqTvpi/kvTywPOo1Waj2AB6zjw/wN8MkzlRFob0fF6FJRkI4oWZ1RW3u8E0p
ImXewmCQ4WFmemHvNoTnXP4TCE10ruIK8oGsDpmMmfCyzJMkaczVmXOmVies
UouclDaAzp8GIzmn/5CsQh4vESUsY9RQhHhrNBzO+pZqnQ8kmgk9hpUbuWys
EvnIY0zWsyWRjhq1MYWORnR8Hf0u1/uuEwM3mODy7wyJvL6wWyPLVZAi9js5
3Cr6gTI9Fr3Bvdu3r8pA+a8r/F7k35o/gn0DggG+HipTkhttUfz1Yph5ZB3A
d358Ku+ec6p3sY0xZTZPaMtV/Z0f+CT9ypXNBt01DfoXw6yJzwNX1SDzvgdC
i45Wy8VVTizYG6A1poIFXVIG4PKTkGKF3wtUIifjm/xkGyJ2Z+YByyoaQ7IV
mB2AvZBpZM/kz+ux0YVor9gKPtC27ullgjP4Za6RGU9N8ObmPT57AlpZdooP
A3QEvrL3eY8ag5tQIBZv47wbQNoU87PPP+Uk2h0OYCc70/B9FLEPZs+WyR7B
OU1es1v1Qmkve69JrI0JjhEozyC6iBj1mZpND/1pVRjfCPosiGSl3cuXdZfG
vUsqq7U4haxBAbXTvmFyDUMOJJ2m2FeFH2+vIMExL5cfFJwf/sM1FNgS7wyi
s/yiDRiwb/R/CyHSELYcxw0TacoogdwDbImK8zvYfMLUSgwUzMH1oQ+lHpBk
B0HRnZEQN76aYQncVTswlfzqDHX45DqwV8rSnveO/wmpCDZyMWWb1ZJfDKeC
H8DeJPyM/ZzwBlDYkM+MAJcF2jefF9jKr4P6MeHoPjRRrsdORums5zfPrsVg
IIrRcg4F6FTlxDGSbIcD7+e+rJitzF4V33CNLYVOhiNovW4uVPMJoztcHjG1
osIUzR9tU6nXUv7eTtSZIAzLkkpqduhwbvNPgJQFKaxu8NI2u/6eUvCzhkiV
OnNZ1Q65wjAJW8KBMyfdcxW3IgqvEDq1nrCLXMQLkeGkbuBrlgXrKL5GXtrl
PZvkaKSoMysjTFLjH9vmuzvW+4UFgZDTxX8uUfd9PjT6eEr9nAUjtxApeFGM
wYtWA2yXfvSw7cGVhvzeNDmg4SCImxhU2KAvj3N8DgWwrq5zd4v7zXESJ3WM
/2+IXEGnX7ICK/Ab0IKcDCAh/NJrE2X0daibHgDod8z1BmC8Zh0YL+ifhNHu
EzgF+sx804K82vzxTnoDjlrGrp1gvZQ/ufTNXbNtDKmuQuibEQ8RLet0v8sd
KpSg+ZkCZuCugjY2yONhcId16OXKfKd4hQJo5xQ6J7uAW0Y+GTEIdd0Oqi8k
/3x7ieZW0lN+q34hRChbedxbgfCfmUqoLR6tnGiQWPC4/dVQ1ctF+YAbCicG
exxO/LgqbYGG871pYTm+WkUkaiE8D367jxh+9bFQbz5iNVFBCznojiPMEMmJ
B30h3lBbrGAiO8I2n/QzPfKsywuIbczC4N3z5lxfly0fp1AB5frzmT5o5lX+
kKhB4GpPu08dycq5E70vlGZbiYOO3dJYdXR07LiOOg3cl9W70mq/CZgFSTNL
sjRWmE/XfmjcbR5F6ZX/UY5A4qk3C+WFyajT3ta/ow7UzVkf5kBDpkTfxpkL
lglPmeo57OJwulY8VRAgMW23+vOMV3TlTSAj1W2x1E6Grlc2Ux2VeoPpdaJs
aNp1/3spkweHi32BjUaM23TbZX+5PctH4xKPtlWK1HhfOzvL4wfw8RERIloW
V0OB9OAxhmB4ORstud0Wh7ClUcFbzj5wawru7kE5sj39INVN8ETr6Ke4PDJo
CQbL0K64F/dj1o7TdHjZETXbMIpDb1PY7laOM8lKtPZgJM/x/DBmvkMOZDrS
qA+dFPm/yqXMCVTWj/iG01lOJoKNSJih0ra+0V3nWNotjeqVAEFgzU8PTEBE
GBpDFf3HJn0q0ZPC3RCc6qNL/kFtrUa4EebmEe49pc12+8mIDN7Tbzdk60fd
U9XM1MQ6vuusUn1Obsmig65K4Dp2eBMfFAh+syc5kfc70oVyptvEmmq13186
5QocSa9CVYFXTcTtz3vxOOw8AoHnFkfAl9trp7aki0wzwO/Riau9afKv0S8d
ocNfFzvbgRC0GgDOXRYzNQGIrYuQjYVKTcIdElPj88PuctZT9TDQ5aEiYPNq
CMvktFQEpLujhAuhQGzp47/jcCm0aFkRgfYT2h5VJ8wyRJy4Xra2us/dMrE9
I751VKJvSAXqSLxripCkM/PdIlmB8tCyN48MWl/Sk9labxJilNZPhB3btaLj
QX1vWIj8lYtFTbLKQlLogeVBMr9Po5dOBiDVdreynQkWZVGS2JqQL8vUwKPo
ovLE35Q+6QpTc6j6Q/PLXz+xYzTUdC1rU9CsMcvxbbZUWEAoDOpzWCfFKYD8
VkQo0N6cf5HGPVpp3uI/D9QK4oWi81ye4uG2SWD4cmb1+fxkv7sjTR/Clbqe
+D+C/KACdRtThbEnaaHH+6454Xxj1v1EB9im76ol9htU+T9T9r+f8ZB2+t6t
BJr6NGT3KmnAqAmY5QaRdQ/aJu7jRyFmmVg9c+nA+To1w/u43ws/b/sSp5AK
lc8GOoe/sSR6rXidi5DW9lhPkErLOK61WJfpEZ6eduHoUeVpgiYjRiaz7kZd
qW06hPim9YXXC9sIjPlhCfHrAQJAC55svXKG8cCg8pIgvjY82SWPt9z+z8tL
dQ/5UGZrHDLTvJSfiQikFNQmAyX/NAVzu024eE+lh5oUGnlPm0f91MGioxBV
kP0l4eHtlgbGflwIftEu4eByeQW44MDNnPGUEG5/rk8KiGX0KJiekQ4vooy6
VqNtDrsNAWn4Tz+PHl6nn1b9h1LQIbisn23d/qm3MvQaA6XrI4ra9T1XhY6o
FMs69tUb5IVgDvosk4Ak2jD+OhbSJwIaM4QbLLExyihtktZJZUzgJB+hA4yr
m3uJ/cNnVPbbJWC/s8d2AhEWlXPLyYsvSJbO4PHXhMiP7czU/0BhSJSKidD6
DVxdBz5tvt7bxwGUj1i7I8FdDTMb3jcJyeJcZ2taJpjcOk3cbUfCk73JwagL
ca9dmeH/QlW4CilO6xyGdf5BctVCcm9m9EUTmB0vPw9HTyqlDINHnaHeHzFW
dgmUfN9t6DOChod+kY164djLkkEyS6OIGIE6OnkHY1poEJ91jp//jdpW5GSm
9mAC6LtH3Rnzv4peJZkUatfB9H0JLk/B1lbIdSHWY9hhNV+ZbqRt/IDxJysU
C7hCMm0Ah6hQR8Vo15kQ/hCgrEHdFDi9Y/GlM/xMODMF3wlZCg9gGJLjjrwR
4ZJctowjo+Vh2MKAsRC3Nl5KmZPsQ+2DrpaE3UVigoDhWI5XNGWhqdyDFO+Z
Lzo79WVd6Ndx7+dVYbwclq0tX6nv967XxV1hP2EHw7BpgiKkxm5XbWf/HWj8
KOgf59JV7s2YvWHlFDfS6sQPW1dVoc+ZkprrcthN2onZhzGBK5nrh6ktXaCI
nVRPPOczChe+Yb16LZvZrdMQTaWHv+ZsnowWQTqxu+GhxGE6KpDhUwfLnLeC
ZE3TxFXMO4fdpMR0UXUcWTm8BKvqgEnrwQ00b5r/1p38nOy5mConva93Vof4
ZbcMNwI3+oxLAG7ueGZNNkZW+qjIg5sb7osBwSdwg1Z0nrTMpu973KKgFHt5
+ZAlgF5YFB6DTG6MRSO/93i91TjAnakNf3VnxGoROYSmOiGvvw1R2WFHsQa0
oXJw/CK6ARU7Mk9m949eac/WCM4fBdoEKzMy7p5wXDIrfmTQ24hjac5YAT6E
WgQ7lBHh56VD9BynzRDdQ6obtMeiIPB9hvbKqpcC4WhyRANH+lR4tIQ61ddC
86TX8+KSA0vwSpvvTF9Upp5Ez7v0s0x5TdLKOnL1cvW8kvvMfufENjH+QGFt
2dfrlDhCagIQdRRvn0CzKTRKae0MNxVX4Vy/yf8ILaqT8835+tRZKq2yLMks
jfD2lgwptjbqNM4Fl641mRTXefCyEeFaphC7Ry5hogr/GFW5YfaPrjNa3Pjt
ptdAKr+10x7y7V677hb/VR7Cg+cybQoLczTyoi7VZzRO1bCQOD3kBEObDGe/
qOhPNsg22srK1gvhedOo26yNAnGBZ5OTkA5P0nC9xnqGC+lLRibovJH9raws
GLj2msvtmPAvhmNSWgPU/2wM6AOL9JRoyXGFSZVsgn4VeCdrOctTQUoACQYY
Yj3fL1CndQkFe2VuMQhS4ube0+5XeSmt+KCc8z3YBoPz7nxUQjR8xeoPK71f
aleunHYfrd/agU14RHPEbVjhOCCYojyrUWif7jPeEkwX0GsHervcF6yYHtxb
JpFHkv7c4952CBnsFM3zeyKn1QRIYelMQJV4zwPhxkHgteKJPgqeNRNwwZcd
wysuYeZTe2UHtJqaBdqj6PdKF0Vd6INPns4km3RSZiP9gw+UwM9XLFNWrtgz
JZkvc3kyAJbNPK5h/P1TtklC6dqqh8f2DlqNtITFl+FsBxgrjFlIyRKet084
dTULWmqmEWW6SAu+MycFrPEkVFjmEsrvIY/wQaNNGwGDjft/RjWJsVluIAdA
uYn3+aXwc7imVlaCi2NhNANCWLV/mnmwgbVRftSIgVJFZ/mqLWgPS8wGWwou
inJ0s0dXx0eNK/j7SEJ0u+LNe33qh+YhoYhy6kti5mAGCAAiAqEZQaEmb4Qg
fIedkuzEvH3sSP1qNeLncFPwydd62mgHjqoQEff6BPfaryZaA2decNOGNCBs
HN9XmiVUxl3CLFrjAOby8dMuIwUW/AHQwR69h7/HRrHhiAeXBoOGYFpDewBJ
eXYrbLMkhUoNOQJ7omN84k9tSkdZ5afATAgp3NUL6H1ONdkAXlSIIWfUobVM
6AWrORI0QmsxjiS5Pmzlq5BRyqgbMAQicTHyVJlu9nSOh+R63agE6iOM+5B+
EbX7EF79FIWqOAD8kFg1cxL/79vWME8Q4jSXpQdTXyu7+f352PNzMVMJUHZk
6ULJ4vqcsWNjpOQS75HYgbvZ5BR13qGlnRs8nyLbXaqMYm6QndIRaefxFgix
bJwPAr6goIB92ekrwn3sYXJ2sIs0mD/phWo1IH4kntX+ozzwSo65o0SjcIRX
vbTLSZOE9JekJb7kvZjEb0qRFZUHXfmy7ZI2mKoFatLrIxSXq0/Tx5oO2la1
lNUWf7ibDHjDqeyM5gRkeVzcoMpRakfRnMdOO9zkeHyObjrIjZeve6gdZxoh
xnCi8Py0GanQ1XAqjzS8QzM65S/eU0IiF/Pdg+dsEv894yyF5xTY+s/+ALps
CIfPl+Y9SijTvADkA5hhybBClKwjNDpBG43pJGIlDuPq85Kw9ICSoCa5iJ+e
2efkgc+p3lZ3Mm+TkmnMGW3yxWGtfbyNjvvgkC5dr0FnslWTx4pYRDUSufKF
cNORYGVCxvvq2uyj6ZVTtxaD8pmnXxol3YSv3fIswmFEzGvtti9OcEFfufEC
6ZCN/2YJJ61eD0U4Ac+f83bX201YloD3p2Fg0bEsp4LB74MU219DpD/KHMB/
MJy8gOu/DNzgzYoIvqrgx/CO5UXj/IjrctOyHD3hqUoubwWgpb+gX/qu/Jr8
2ZjCgTizKChglvm10wDuI1SEhZ34z2vjSj6fp0t8LxkEQlYycAT2DqryVa9o
vYoBfQoFx/FspKQU5UJHTPq+7X8eOFDUKWY5l9b9qmICcfZPKiSdgsvD6Mns
8anDSw62WZt13yQAOOtUeyiscej1+4z1I5JHi7NSMO1STUB3NbwalEaMmW3R
T+pavLigQ0XoO1CgfuHffLKnHpHEh7C5sKgOhYSWeldpjb2ePv1mMuDp859T
hAB6OcK1TPAft7OAYM7lkyMdoofJxsuleeQI4VR3jbW3iWk/rOzyjB/BJuMD
tmSpIMcwey5I/eaTKjklwlS14SzLf+KVdnnxJT4ZG7bF+dgIZkUXgbFRDJLY
I8P3ZBuNtziWDiXGwuGiTB0ord7jRb5+PcMIG+qf+HGyOYeGK2InaDq8lTH2
ZznXtTVjkaaSH9j6CI9prODJWXJuzJ9af33A9hCnlpotZYB3eCGnOtGc96nH
OiIFxDOa0/RVr/W7+/oNHBMC33siAiPZPxf3ocW37qn/auzdJHAhLEqSuFnv
5n+YTo54JyyBckbj7L4SP2lE6HCDzrVCNBdZYY5ZFGvrZbVgSQ0UgHr6/kG8
h1NYkRK3DY2QUDzs+TxGR7P3s0281MkjtdCHXnKhsxs+UY8AItYHRIjl0fga
Hv6WruoK+0/WSBzTmNhU1SnzIKv/bZg7Ax/ZRj6B5mxyhYruw8OkrgJAVIYS
t1sKpqMI8UvBwTnD8MjWM4wXGKtn2eXrC+3Vo7M8vy0JcQAfnmstqZGdujHO
sz8GeU1i+8AFt9g9YnGLpI3IfXXYxBxF0Zm7I7ZrQFUTgRGRh+no5PB9ZJ8R
IVwCErdDP8DAooqkjAU4YQunvaxvkjVDUgw6iegj1hpqxmV+uRQleeItXvJH
9ZT9J8+Lj/2ijg9sJX3wRFHthCwpP/Ev38vm7CYvd9K80dqcKsUtgAfhhAUp
TsSgRSlwWxRR4vKX/M8dQ0lyQ4TS+ju2QMvcmcTT0PVK8AL6cCWjgQIyopF8
AWrUVZhVy+H4H+ibzUP4XcrCm2zKEXiMyQy1SzQegf/C16XrhIlLzQAqiovQ
Eif2uf3XYPl07+n3zuYS/HPPiR3AB4WamtBZuWhWpmrM4FBpcfJ/luxyL4XM
nbdNTRIkA2xtoUSjl2/LnzfDcMrXCV9k19PYTiZOrOfIjYMNAosnTTC39IZ9
TEHm702SP1D05JWZUwC1+FjyuSj2W5kF2o0M3QzrjOau17a+3hlvgZ7Awhgb
3pZsyxo1eKpWWnbtuMqmCj4YfLGanKCSsIy7HVSwBbRjh2qHp9rOD4JSfSsN
8XPHkDkMhk6xAl4HP773IqbyLY6v/fltB4qXORQQ2zQJVWq1PhI7SFTvuuh5
LIbIqRjROlLwwQbysh1HeB/oDFX9gRoUQ+/xF21hDtBQrzr9pIim6cblFpS3
IHbXvUIe2vLkJRQzFKgkK9euS8W33X3JKhJe+nFbqQIe9XcGldbU/zKZAmLL
t7abdY+NYWqdRLNshyxCrnKSMpeyAJ6eBYjXEmgZ7ehMmjNYopveW54peWZn
1icOEuVBAt+ZjwFpsvlD705+5hrOXQ5qpGfLBeKf4MKMzQwyYcTl/faAr2Yv
16hcrh9V//oKzEZrQuOh3ORDup1dJ3FcN2dOoSIqU1EtKujj3dq1FE6kkxME
IYbOvlSvhnRqR5Y6xW++5T5/ZsfqYhHU0VjqlISXY5t+ubi5cL3MlLUD74iI
TN0aIO2x3ip0a3Mtt346YgjgMIqSPX1rDlU3RxLZFkU2vauvKhZw7oX5NLLU
nK8Z437TrndRgl5cu+4Le2IioePfbewVng7foKScZaAWKsd1UJD6+0cWhMN2
VxRziR6BURQn/P4nmHHOekGI4oxYDjMZy/pBr7XPBboHuP84AkA8c2gWKfQ6
JeEm1kRrFzWZN8cG+aL5siDYaHK2WCgOYIqRf9SznmRd7UDwOxorU0YKk3oS
Uv1wMnx42AP5wlyrl+YSeyFEE+HqnJ7gyIGV1/YJm98vdNKsyyfmCgX2nIHT
tAScBjO4xJgmlOTx1nZE1/uEGOaQDScy+yfxxpSNky+0+m3aJPWenobRON5T
mUXt2jY1iTIIJyHQJS/69zg9WVJN9WxIdcrWfDNy6GaOagtOakhKCsnGvv0Q
XXJOXQJE9vlRYvND0IXMswAzszPjwdtLCWz6gTRmSJrrKwEWgZ1D6dSjpUXb
5X/AnnMpC83ddF6Yoik5X0uDKnTxD9yWj6DdrLIAR4vMbETbdkUXnrBc917n
NHE+Ey2h+9hNr0+FdPJQ3QN/2EBGVFg2lsypu3ytxmnrvDEJYTRIhJq2x24m
wiM40fDGz+lyPO/4Oru1VvofuBNseenjfjjHVKeb0jxrHBfz39MGuIBUO4Hg
ERwWyhLhqea2/n4rmRzjPA2CtNUzCtKN3aePtGFTorvcUSO+Q6IwjYRrgFql
LWP19MMoUg0xCK1TASXS5msHQMVPR4fofSmLMd0LsF1Hzm1UTxdr9HU2CL1D
XO5FXEaLNSVxkIr0ZltiT3TyhGjKSohMIyP9D8x/k2xF3GdaUQVyIH1MKA1h
1GCMpJP9y5cOik5PwldnxhJRc+Oyi8xhwo/Y7qTcYx6EbiPCVtJT3BNnpjMA
GOt0xMdNv5s5z11IdRx9CfI61XU1WZix2mXz5wGjfB2W6+eU23B2NShfjURo
1uyx9OJCPqF1vULqAlvGe5og+65O9UP2WzfUJdIFyKxXyy0DsfYJ5ie3+TaE
GQanTX9KIakAp8kLlPkGyRBVMU7e5objOgM68SCLWAlmB15cMvDaY6mE3lE3
N4wLMEck7cDsd6mdeGKUJXaQ7k6ecOxOhoLRul4qh1j7EuhDIYKNOSU3HI72
ZEZ3k4i/h6t7k1RC37lNVeB+HKE5E2tmPse4Hnc4qYaTaykkWLXyxTjYtnrm
3CriEvh4M00IwJiH5bv7QT1fug/S2OgqO9LKW5Xr8+LKWUN1CJmZSxXni1R/
Gy939hom1RDUMxhAX7c845SsEv+OoS9idIvdG5HRKMTquePJwS3d96B8W39H
CI37++y8Os0JaaDzYTfRYEFEYq+ILiMhxNnX2PVUU0VQCW22+r9GMgPk5WTj
bzm3UoM5cvoqFD/k+HCt489bFhMpgyrm83SpF5Jt6Ce/48t+kmwt30CUp2WZ
Pi1jYj2cQ+2RZXNU34LExJzc6C9/KA3CCj9btMLwpVqdM0oSMosrY953i6rv
nj8H5Ta8vetDHSvOPnvco30OBhsDpj75d7ggVQO0kPWO6rWOVGV1G+fs1Miz
4ib11NtJdm2RMdYBAKwxa0t/fh7FyDjBmpML3C1iWwABsVyfHXLtLHM3d2l4
cyuCr3KQOn05XoIn8ns76+gPayERy5QOKA5teN4vrphdIVA2ptg+SYNuAh7n
XN9/rFbSfDkN+yczJ8d/wxGbeugYh9EJnvrcJP0O1XvNzWOJAwDTVD25/DX8
zyOYfuSprTFBme4C5Gsn3EH5vHd2bEt6PJ5BS1gaD1p3mDq9u0rxfjgBqoq4
r9yd4fkD6IEbE5irGb5/QABYewd/o2I1yEp9NWBIbV6hCKr1LI2/znJU9+EK
WPVwu+pDZ7y5MxmeJRWw7qolI+QZSpO2a6Rt5YpwC65UDtZpmUpfmdgCYfWj
d+2x/yHBlX1rqjcKbI6HS3whehgjz4Soqj1BwOdwN3Ff5hmFRg5/DhNFT2BS
XMBdvUnoaiLKH+4HNKj0Bwry/XzqVae8sZnyizJB4+kKfsg4Og6ucCYysnVQ
K8QAo1n2+N3EEXXu9sIZSxUw8BOBqus7QU7u1UbrZqnWSIGl0CYMEE0kEhM6
YPxPWWhJ5gH4/tceYHUl1jI9MKK/z0IzNytj4AULDai6Oy8MHlIOoKiwDF1u
GSsyEVf/aIJ/o6xt4qKRO5U9daD8njyYkoBckluxqzjMTmQ/AuvlVEi69MWc
a9sN0gmgsLGRx+Z+hbPrf9K5sP1FqugSC4O8zWgb/JQ/it4eHMxqh1M6yhpF
vR20NYo6Riqm0lgOeQOhl/Esf6e1GUOLaUzUtq3Fb/CO4gw4AT+sG7MOMZy7
ZcFau7pqHSOVHIbXI42ZK7YQ2BiZT6ekjpfbIcV/2Z39UTksEUgRcJ0FYX0a
Hp27LPxBb0ysuCTWemFSCQcx2HV7E+oFiwqCl58Ur08NqLbn+4WWeIy52HC6
q724geR4dVhxSccHJj4dWXJdFSWVcbnjNuN+xff3g5nyRTaAO3k0f91wV2Wc
j2KbSST/1YdARSV90LnByNppVY3eHa1t3Y8OMps54Dtuvmr14efwz/HiuDGn
gpxDDvnhaj3RH+C982SbpGax14vO+qJF8okftcBpYR8VgKSEfcoUHY4QUi+a
qZa7pyicmX91VEC+nLAXSPfn4p3qR6u5yor9qvMNblYT1xh82imYnLVidWlI
okzFrklwFYep7Vsih+VAo88fB6RZPO8aDwC07h8hcwpDNcpqPaZai4HBW5yV
5lQahGUizfWfccVP873YtgByJ0DtYrA2b6aOX5nl8a79xTcncFEE1gPp40BQ
mShdJkX1/lo8nYPr6NHjCorDhPUF42AiewvCate+gD46XUuJdCYwrZXlI5ul
BsLQB0CuXOVzfbZJHgr64ZwpkJVL/Hhx1Ba9ocMPzN+B4BthjQJnA8w18YKR
ekLDZ4paRh69Ith3P+KJyUoAbKFWE9f/NmUg2lxnN9UNIaZ2HKR4NfW0AI69
SygQWch88+YwrUOAhjkntts/n+zgalXUGzM2HrXzlqxzHDEhkn5ziiUjMjGE
qG7nwb6keQ4F1ZTMXuSWS0ohP3ST7S20sdv2SuFBosVr+pZ9PLt0CsfJnmUx
Iy3jwNodDbfpW0MPMxEMxHbuMlR9o3ApiaQhMs07H9ZZ/ZDyC6Gu+r6Z6Qoj
0SO8JKbVK18gNzgUy82ewDwFqSe81s7n42+ZcVhXvAiM7N9mW+tjfNlWYJDV
HlRRaczyvH/ayngjpUJGyjm3E72PPTznFYfH+KetWwr1m+/nm3XgcZB47FwD
GC08NqqCKiYwaNcCeSOBx5w2fbSRhY7BVAiWmbPIXjjKo5FuFstQfzdSuLzF
1cBKTk3xn6znP8e9aTek8Frw3R26BCWV0yCT0CyknbSg7u41Fw+ZaFglqlRV
bnALq3bfK3LBgu3Tf22IVOeTHLlFwVzBCXFPZh+FDDjocymdKe/SOiGVO7dQ
IWdY9f6XFsAc+RQF05ZOeVaEXQyZE6sjX2HhKk5Jc+AxGF0V5/SEKKflh/ft
s4fGHSC7LG19NvLxMBqya27Cy4fOTGiVlmk8xYhVvjdC3LBIpgj9ihNKYWD/
NJuZ4x3OIqg++deFJgK9AvZcHkahwwVHnWgGqzqoeMumLS373BxtuWd7V05W
visG2kz61sx/R/g/DECuo2VvikaPJj0WVLPQHvhvx7ZvdeuQTb6rJZdwqH+y
Wxplfdg0IGW7269VCwggdSS1LKP6q75MTqRme+QqEXa/iH3wol/3/X74u0l/
jGswW0KL54Dmp1SNWOF1L7/MxWn7T4oYVK2b8/IHPcJpI2jjc/pHMZliuYi+
gh+61Tz7nlPAmY+rxJ8OCAbluX2pgZmSdFdgGAuFajzlOLTuKZDJlK/d9kz8
juaN8jdHX7aSY5kCirwe0pUXqU8RalkGjGQHSYXLjV86HXEcVcqsNVhdKPUh
/PYtG42A1iPKAWll4HB7XB+LLuDPbbyGFroRaXOs93WPyiJSdGJcac2r2G6D
m8NDiUYmVYMFa0iSmu8MUogoQ6ThRyjlgNUXMV8j3yBNp47CJy/aRngllT3N
CIUKqSBPx9GEiY/GIAxe9K7EKfWK85HB4PZySzH7onIOhjVubpagtrFaSBQ6
CL8qEyYuY8DQfh8pGCASLqC7S5eTunJso6nmX3JAAAHaSbcyei4q25Yy468Q
ge2IAUIMQM/B0/EmhyR6gqEJxss6zVoJULh6SrF/biLM8FXW1SM/BZT9gwlw
qoJPDNlUZtunhx+TT3TRVv0Oya3iXm6IY2nzclk2GkqNLxWq1PZmOGzzCVFT
GBiwVsjKLw+tWGpTyW5ZoXVqISR12s2DpyNCTJfFU+nExVeF7HRci6CuHp/F
hRd/+hEQ9A4cZB2xeuiMCC1bsy1mE7JBva8q4cKDQlSjm197W76/Cj8r6rmK
8JisGLhwJfq/F7s3OXb0TOS5zXBBxGjxm6JTN2+W7CbDCs5weDBAB/uIVIdL
RaZSDIMxvzhAVZlJJhIEfryv4mjK/WW/9AoUbP25F4qdbZ9dVrM/wFKaQdjS
EwQkH/g6l6Mq+mwdo9xFeRR1Y7Ww6Pnh7JiSKaTO6h4x6/aJaSGVN/P7FuzH
Gn4D02YyZvCmxSVVamTgI8rbdqvjFZQ8M+aYV2okTTxL8fGhQ/vBEStiApoG
SdSs5tEOKX+Vmpdhk83/XivtVjlObSg9lgqtFR/OOwvT/8mKcr9mt+swh4F5
UWCba68kBFqzMqGr54g9fQwiMlMuh4FrR2W6IPLDAhvOfwKvdrI3XW3GWxaZ
/FUkgmNeBx+LI54+Niu3V9OMzTZTt5Dsz6f5uh3pHuy7QPQYcVV9unKjkyQq
mYsxldBGzoDsBUF4Z+lFaS1VF3ZdP9acZc5shDyZlqrZWPtX8liQsKZKe+AK
BFSr19BkzXjB5RE0loerWWGXWgAP3D13c6FGjal7C7TE6VfgGjj6EbSa8c4O
o6GF76XcpAFHjNwTh2/j/Wzm2BY+1fzLwxtuu8wpCH2DrsZMRKM2pgvCGgjW
J5fdSWKtf5Dw4DY/I332ogYHbt2oa7QiFkuQQGCgeP1aBw4S73MwpJRdA6Uk
utbl79FvfJ6Xr9YsHj5XS8hQk1y9SGqE+XX2Z7jOJQVXo9r76CNYafqfmpZb
dBmAylPPDPYYeCccmyxqw7W/mJf2rGdeCjtaXg40w3/pKyUwLHK65vLuY20q
VsGA7969ZyBX8+N0zSYU6kpFVnAmpkNZZAMdMxRDD/5u72+00MRzPeqysxU3
YaR7z1u0bJOFiIVqq7UL3iniuyC6Q8VnK0wK+E3tzHntvVxhEXFfw3+BuqZI
sNe4pPBliFWnWzi4PyZ4Ninm/nNz+23hrdBkj8utC8v3KEpIpdfbuP4D1/7Q
5mN03/2cE5mMcxKDrd4NZheDp0S0WdnEgO+qJlkBqGfP4BYxlkAg0TvjwLUm
00pgpUTS3Ef9fEUA9jA19PsEcVyMad/9416OBvHc0yfra2Po/gGAXZ6kMI97
Cb957yTgK9RsJa61BSJIWlbeY7m6RpkTvpGPWYD26w8pzgC3jVDp5WeRVITd
g8NxALQeDfmHAoFUpDmsZoLxuJp+B/P8FSXEi7lb+xjAcJpLAj0NUjSmBulm
trV8cAb/Y8bHO7jrWtSVC+bqEOXUhlMq9UUevkmWxhRLF0kRk4SRf2S2W04G
iFdHslpN3Q+SSZ4eQwHCr75GLjIIib5l4IBghDF7s+8hJ45H7xPCtb7jdnXb
o/lJGwEQGkzbBJMmWBdehyBu6UAKRZ8po7HDIQyFIeaPlwDzOs8myI1V74j2
cyp7ZX+4VDFA2Q8lwmQT1bJd/Y1SUxZ3uciCBl+vZBT86gebO3IpKtBmQmC/
l8aUkB9beJE5F8QBavFp/9wzEk2drbset+FfEXQgiQs51uULg67SOYhCasB4
I4dcC1v2oX5SzXh2buJDOSg3EmtdnDhT5OHX2ji+5/M4QN9Ea396Iq+unciV
6DzMr4vdudRwVQr8b1hussPeFz5jCPafhewZX/pc18aqtTfqgbFO3Q/y1+KF
ZtEkTnHel0oQO8qhyjh3eLyl8Q1rXiD3GqIky6riwvFkL/gyKsqrL8TfU/BZ
jqhUnUyTO20CRe+u56Dh9zZeBccKuENRp7xoTZBSBVIZp330Rp/nYy+2QnP9
xsjmbc7wF/hDco2EPiH0d6hT2U0ewxXf/0OTZICajKYIw0+9nL8XwWpGLmk7
zct8FHqXCgpavMLJA6k/CAZwaeCQBhv3dam9NrtUhe0Gj+aBLvz3D/r0O7nD
TPMucOoE+vWJzTkh8+nd1HGOWecaNDGJo5zAEFgeWgk0bVLYCzh23ZlfAnrm
vWSGpeWMlj/hzAjQHiEW33W4qO2Sezc1BSV9cWkQhkGXCTA3nunCVdoTfo/V
TqXSDzW0ajvIQc1E6yEUQH7Y9/yidkvTHn9ObtiQTImbn1QuVbGOKQkbV1ju
wS6aAjqXCJhg+6IQXxcDD4MlZUEp/y1cu6gLKgktjk3wIEJeMFdKsnwaFXt1
4Tj53D+FA+5pxJ3PXpc/oJoREd04oH2HuDiPdbAhpFdKLHRwdpsgp481eA1c
o3zi6392GcdkvHgRMKeDKVo2Cc4pJbelVSkNdLBc0X9qvD5QqA+oZNbtw8ab
00jYrw3l4bqMD9NBlr1BedK4oslN1ne0vigqPvHKtUM+MAcdjykIFgepE+d1
kW+WPNE2Mkt0pSR60X3euFu5YKzbc0sX5xE+lsHUEsa4MIXxTZiInw5Pl0/F
ZFd6uf9Uhy8o9BBaeADt4NNcMgBbLoYl9+gEaZy9Xs6QGM5ZScMOu3CvO19Z
NM/q2+nEpClkTYolRlxTVEVISowQ9rwtp29rfpkq0u3NCo+AGLYN5yrXa1EX
N35aK1YiWps1kbukPFh7OuAY3tzZ33zl3GNFKk91m013zbsQN/A9Rh8lOR12
FxDfFNGwOyUNyxcV1wT2UKbPVrHMqAmJ98Yp1uMq7VdJIHvubt+YhPiFjfKc
BH8KK4834Dv0zF1d4dm3ZvzZQEiO55scZSq0fMVJuS1XRBr5aePrsPZltm5F
TXBoxq8zwDIdp5gT5cpvrE+RLdvIJirbNew4ZBRz22HTmVA6TNrSOssFnfmv
ia9OOVX9arQy8gOGK7wjnytyPZMOVRGy5kt+b2tOfVfTwAC6Js6lh5Amkj7l
yOghBfoZ/GoWMgG2Im3BHmD9zXQCOPDLppr+O+WUd0MYOzdE86WOgo1Xpna6
kdmvKanaErZC4OMvUz3wruk2RJtgCGwOgJNgI5J0X89gEc6O/xGRYTsRGxV/
NBCwwSnwkMmPlsJwmwBlh0yAF9BJ1av0FFwDyTaIeSjKuth7VLEzpHOnHELj
mgrgIDsSNsbWh4FolfaedAKHUOgsw2uliQVF7jPrQIGAdcFBcxpKEshxU9As
6MN3m3yy1q0YoxP++Hb5RgrjS9JRQ5MdKnK82/NEK3+nwLwT3VpOspZ6V8vp
Y/F3UZsuwv/xoMqMI2UjEyHwoyeJmRbbnhcncsROaBzjM/Gws1oAbpBIZj5i
mSQIfRydX8KP5B9+9GyQvB89i2Ptf7eJkva2byraKWJZkmbbanQlNFNa2nrZ
53d/KMt7ZSowEN6ROuc1fbIIAEGTX55a0GgqBDF6x3HnVIbhxkK2VnT1ii1n
+EN1M2YzQW+a3QaJ7OsknN3Og1aHGLs+nS5FAvujxUnEvBD2oorxN79jSSmj
1S57QNLxIOlBIZIMuG9mV6e8XqQ+2GnN29h1udW51LNnVJzaacUOnwCeQiLj
nBPg74QthSYSFfHbB/bpNmcmol8xjD96fJVLuNsDU/Hr8pPd5GucURNuJNio
lgxqt84XJYaoS9C8fhlCm1BB0B+QmMSCMnbltLormSOxhctwa35LkA43l43p
+9cCVB/+cmaYK/9f5olEcKFE9nefoetx0ouCTOE1e81KkZITEP83fNe0pf9i
bbmpWCOU8bCfRBbSUDw7yuWcamCx3ldBKNd7m+P7qE0aBoDwXDbnoNOb3kha
D0SdShHMDz+J35xVAnX9HBm+scuyxm/G9VPxWI5S2PgcMcXKQ/qmVRYLF2gG
39gsnG4T9ekSi6v44K2DxRKX8ZSlclRi4dEotAldAxj/dn5NrFCkgmXqc/zK
yDhyVTWFQu+/Ox34bJ9vp8jdjNU0sFRykRUwBwBMtJ5R7imtV1HyFirgpU6r
6sSgx1q0dEeRGv7pqdPZXRH+DJNLSdERsdbVQOm85K9V3EAlZd6QTTT95xc8
yDL37nsQp26fVy7XKv6hg7mYt7HR92tLQ0SiPwgu8NJgEylne3kQf/YzQKhA
qH4xBlTJbJ5ebsxz6JPgKbph8LXrJ6TJpIxj5v06sMljPLVULoZsHOqYVLgj
ouaTug7RCYNlJeIJ/a6MO/oxoEWiZvIF5vpuxAY+lVMtRw+BVfPyuYmMZ7yU
Vfb4oIlKsSzrGe2BBU2uv/a5uQCAJsRyMtWi9TUH7Td1HyDDnESJmg8FLaNv
C9URIdrvgFvyf3+T1RC9v0+cOgWSL4f16xC3BIkPvm8HYiSVcezIP+VQiBQO
LI2C4dGHwQUiI4jjQQU8GDBhEVRrPYnMl4ujla4zxlMI79Nx1UhOVEC8b/A5
WuIlDnSbAqc2YpfGjS1WsKOWVi++5Yam7KxrKYrciV8TfqRnHHXf9cBAWkEr
2uL5Rg2ASHCv1JY8pru8dg3/lPSYMHxpENmIFfHseJMvv9dRf7Paxy5BhXhw
RkNaMky5i6Twf0hqFauLtO5AY3BP/3Omc6Mu7blJrXo97gF3COmt+YwqpK6i
W22W7EKhpC9LBYlagGT8kfZYJ8MjNFlNOFP32P/+kaLXVyyG8/I+7xng8RSg
hIhXweppQNzYVII/jRkvQ6wYcM8olwudl7i0sLOBNy2fN4MfSqE38nSxHW6v
ft+mDFCFrfHelvdtYOwqR/UBuCSd/Vgnwat7O/vzjTbOdc8DM3pIc5aUGG9p
d9XNDpAIiGxtw2iUdq2QuII15gbJ5giuacKFw2x8ittQrkRKfPlBXH0nKqQa
KTJkTM+971FbQMeb9rbd81bvNVwSXY/Jz5lK4G2YNQiCKsAH/EULCrNeXf6G
A20IqoyjN2mRP7zvXSq8JjxcYNyRB1gmQXRQyXsUekWXaNxykj8yNOZaCWkX
x+x9ccIRLr/V7WDX8Zvs0QWAuwnVDiFTjwDL/V7NS6BPwUhVFJqVODENeEhK
hIYIwfEHaahhx9PdR5K0s4cqGDNdTmcDg45ifZqxaFgy0kqXt0mI8bwb7+Nq
QleesLxPvV11xPHF7TQsPcVb3AT4SKWLYGIPkClYL+iK/Ev1/DGDgAyVttwi
OU+RVOIhILT99YxRGk0H1ku4OYUZaJ9yBRbRg6dz0ovL8KXNhkcUHSeg/5TX
zgXlkyr9im3T7TZ3diSpo2F/buG7KPaikxKD3ZFgvITEzYygoLwOp7C5oHdI
5YphZ5JUhUwPGNfL34a2LaUgCjL4dq8WTdW3szWt/GKGmEtED81Db/Svxt03
5xHfP7Ncr/P7l9dUTDsZQAZfD3IMqh9ZPtATWHJCbD4b1O7h+amrCKngrWli
qJRkKAQz/39wHnUlOZo5gKh/NcjpggZtF+A4xRjAd36eFYCrOg1CHUHfZC6C
m+04d+1jaFd7nNICsd4A3FVcg6rzsRYlyFFbu8QvHm+jzjqoDqSDILwWf2cL
BmvN4DPZkuJj4yaLUiFhlYrbZob5Vk3GKdmvYdpFsXo9DpM4029juIpmTTnI
FAWe6YMx/SDeAJ0gj7FwLKlrgYnW8L6T0frvYWpwG1DWVhOa4JetMOLzLDZ8
OMCwiQLQ87mpcvrFBuqi+e20enoxPK7yUjFlE2fMApSEzFnSyUc3xEfLuo4Z
wyDEbRX7HXTBkYujhLKHQeKlt0mEWHmKQS6W36x24o7VDitUYYz4P8RW6Q3Q
SX/gsGBdiOxI6YDNzOsZAQOKX8v6aBaMo3VSKIq4ce2Z7SSfMlTsv8D5nWW9
wVmSVISIlHjfiWYgv846KHM1mK5lIM7APsOoVmk0zys++2XG+xfkJ9+BDlil
E7BHtH4NNeq3ngZBTDBmtpru68swNceJr9sGHZykIJIdrGGZawKQ+f7VtZEu
6Ro/kSkHgTI4f5B61LEu2G7MJhPh+09974l4w5SadLyHz8z8Izp6pgI0+AID
jxZzH1K7Bz9HFmzKCbqTQDpcMLPupABzBRGTuUJx9xuveSOVrfxJIu2/3wha
n8vXGZ2fJ9e4yNv8HK1IfJlG3Hg+P4B2JcAwsa0q9vAa5fF1OLSJDW4tQ7oV
X9lb8jP6plWhJoBCOqpHGkslqUoTdVaUzArQZGywt6Uq4ZUSac1xP8TuW2m+
U5eS4IXJWTpDZXKSS+sA64pAI27ylQmie28ApShQLiIo8oVNcEmhPH1Zw/WF
L4TwuKAhdoguLtgOlf4NayBR9jiVDhw8EzAEhMXt/P2S3N4DfpFwyDpthkQt
VE5g3AgwSrwTw3mtntrTde4XTZKjOwQO97bqqofQNk1Cw+jENC3RC26Fc2Vd
ycIPztTBK282fRZHZvqcgpQyJApZeZ2xuR2smVw+s6zgvietVh8l5kAZTFYd
daoom7KJ7jdN0g2cLrGR3lICrrEcjR0Ay6Ix4jI2T/sJjWCiFN4zNjGq4kB0
F9to44W1Su0J1oBHUa7mXi3vylrZfAjm89TNla8ES4WyHC8TjSvFoki4hjXx
fs/nVOhejbNUQtDzWE9AodcZenQtFqCxcJCamQOD5dZy67BBG89+OyTBtkvO
4dHVipe3bQugJyjfwE5YBhxk0N/T8pChmvpVqrzfYC0/9D+gr/eL328FyHB0
4csO0Rrc9Py9KuM7rvPL8n5gnna+LMv503lFGqM2gq/Lnfk88m3AXwlDf68x
2+Lu3SrHTCiIU47KImV8dcqLS2H0MDdYNgLm5BCylW7vj5rLlo9vV9qcuUeC
gszSWI/z/62mUrIofoWt3pOUhiuRTobq+AaNrw64XBDYmFxMgfQgayMpXi6m
Y1zRSv5nmDWCKb+q2XpxVUFINed7p5/TV+irRiAGkr3bbadB1591jKKJi1CR
YEg1DOhWxRk0xIVrYG5pgPLJ27g/5SHjVKH0i/jd0EEKlHoGpCU2JL5ZveEr
EQyN14Q64QdVG9J72s2b1+iu1xYPYCaovGiZaWpMTyefo82VMVmwGS9uZwO6
an0MzB3bJRlbimJhwksNa9Z6wV0gs0rxHljsdI29GgyEMxuzNdW0AfoIRmnW
TroKar99nnJh1Y3O2V2UD/2Vg/mtrE0/P9oaNjuLz95xqaan1yWw56f9EQ8L
t/zR0mY9MUfElSo6qa8OixXlfPFKJalXZstZzbWWllkVt/Rff7X3LX0yVvuj
lKttyDDVAwTQQ/BSM6tq4nx7K7hkus8j5xtqY1APdCRzbxT6fH9gSftPpWmm
MvdQI6agn5gJxWsvR3hYow+seA3QGpCaSlxgR3oLPxeHhyha4NGeZ7UGleS+
G5M3lIR3y/KKfuNv48NuVm2y6Lc024B623G3ZUuvYYK7nkkuX40ZpL8x7tzW
em2OpR+mCZ8+DSmPnrOpKxAeZ1Pw0AK1orOqomIMAAkwBGcMHXB4RWdE3zNI
E3rKXk1tXvofEO8fVqN00+lgzJuK1XxhboVAOk64hTW4d2vngRLPg5PWTnIm
Pxh8OTFaknyQ6Bpn59bsDs/oBon2YwS4Ncw0RGhPqssHbzuYDHr9Y19TsPkL
Qod4RLGK7aI6mK0A5NKeU2XgDvtzKuyeYK0+F0zDptF3gMizzF1XZZrcTozM
Yw8lr3WGD13exyMlWjw+p49H8Bas/8vqNbEkHZzvQW+A37se0y20jBqWWEnO
Sw/CpDfo2ApQyWeIEqOj2kCE95qAFJF+n2zILl4IVv/iLXuH588eu5u2tiDi
kTfjZLBQavnYvkicTsOAQ+6JWrZ/P2EJyzTD275FmtxYf8nWFQL/8n0Re0vl
cWG9oi7EQ/lmE42/wyAlxHdXJx7HmsO6U9SMJOEOPfO/Gnkc38cbk5avHPLs
rlVa9KaCqHNgsyMn+m7/YB2FaH6kpMjFp/x7YKXr3Ny6yc0D1646TV2Y0Ndu
405zwOi2NDJqoEXjf4BYzhimFE1uoimUTCO4gshC43aYPbdDNpPDzQa9A+pW
xny1L8xRTJIX4bhUpIpAh648jqF4fH2VQYMkxTa6zT6P7JbP+5+6oZJ1F3lH
ctNPyxP8OlKGn1hQX3HqDq+6od3Q05BW1tlZp2s5zwpgv3u7ij3O4DX0WXQp
8MwAE4ExcxSMKYrIrs3jGIxtZNoTTiXltrVAn+PZw5LxOlcdC5Iz9GnXEwaL
PS2KOYXfnMUHEVZ0GkM7zTvl/yJ1FQobj+fDFIASzgivaWJaGFYdYhjnCp+P
zHx3QvgEltmiJTCf+oG0yn+RK6Coa9L/DNOrqX6GCFUjwSMGyAOWRYV/pqDc
fA6pO5Cuput8XEQaLDewXhDli4RRcg7YFa7gg7InyXcwvdahB4A/jvkV4Skp
ESRrzzIPmFNSYcG+tnfqVUUuqschIf848Bl61g3YNXXmToiJ41XLh5GMvwrG
pniIRkvzeJyc+SkfJYxOee0ZGuEhLlBTbqjYdORVo9H7tKdZkS/EMaI7ryEN
D5bqYNuADnGxsIZIvY+jrLZyNqJ8JbdYY4IBUPm4MX2NrN3CxlD5X4t9Qf10
lYxiY2Wc3nUBzmLqrtyMlSe94Aci1cG3tsKj8N5vlrXfosQ39tsOb8KeZLxO
VqfQJkwvsxMLU+2zkyRctStWi5uKarogM4mePMciyoLGUS8NhZ5P/UqopSMk
BDDjT+h9v024pa/IPkZWpxhcplRh5Ws5EQexce5SSxaBATZR1XSF0HNiH5EW
7+5HGNMDU8fHaXurnb1lPU4PHhkZRcZZOfjS6DiAr/Z6QVeZRbzzPtk3Wmuj
+1JxFaT39KVLeFNRdpbWHPwTT+v7VEegD91iIOcwQwGWhbhxPvAikHx22yCx
11KGqF8ol9Ma/zHHF2oceUZb/xNa7togOn1lmSunkQZaMleBJimGQIjnf1oL
HFAi05yu1q5KrpF8sOeSid5OrCbfHYLyszfBE0fvQuv4ysCLTFUSbMvDFb1b
q4gKKwEvzpHNYpGqYpKsWe8t7gUlnV0qKitgon4XF7hcrcSfkouwVtnAI17e
RtupZGThM6AQMy1k2FvBqVCBZoc0sQN3XR3AAwp1BJiCdWdptNEbRpts6vkD
+aoO0+3fKJCXLhT7NA5NCQ8D883oU1LjNp0mJCd0nA5DYdRuU0Me9iu8EGdX
e2S40fUhizsCpfBIW40iH3ryCFfQwGSsr/ihMt25ctYFcJxGSsPQ63R5WeGr
meElAwJ0p5T6x5TRrHRxbL+on5t9f7p8s5r/yuDcHnWulCm5Vepn6VrS16He
9ktBMVIUnI7Wy9d/7IxrIt1ubDsydfKfqVtgxHbHVvefGjyibrNB5+muPLKl
cAcx9ufyxkl6KvjyH4rH5ed0XmAcIuhouJK8/AWigDbz79/z9PwBl7vsEDsF
orTQodKznYPLyUrvsalB0Yy+S+x3nVTyJh/3DJYCOvucGeupisAQRHBkmpZJ
Xr7HmwqYrwbeb1afgSRfKxyHlhXCgM5yCNPcFKwnGtBE9uOXB164WxLZA/IX
wrzJGtZw5shgfYoDzukZh585rciS5BLChkBm2otR+SZfLT3Ks1Ye5U5YJGG3
xwXlIAv+Txo3x3coZPN46M70jr+7hyyDsyPNB1Xry8tURml2sfWeuqRkmGe7
7Ia9KP8SDj34XpItyAcfWeXV9uETbOAl2Sg8U1V+ML0Mt3tjweYBibCocKp+
WPlLphAiP24uWb2t1DvEyzZdMbEfMSlYWHNBob5uEwBJgr8QAzHYnOjfY/h7
9RXCKqY63HdzIvI9D3Ux0VSnNEs5Bj7AliBgACuyPZcswq/WhQ6ydPWABtDA
ZjDCTogaElHyrnlGgwjjGm5LOzbVFdhSxbDBOz/m08ObQITHQ3B7eRo8CfGF
sMvrL1bI7HkVUpR9cxR+6eCs/zRsyQcQBLsNEhDey31OnVj6v7jsmA6MPJeR
G5/7PawyBVh1Sy4AGyCm1t9//CvguSBrw2iL3eyaO7lUatzdYthdoCZCILKU
1VnkrUvQ/3JLUVZNvGKwDT7XZ3FDh0H7Tjn2ClunVlHMZx9koDHe3Tpqfb1F
rnubh5ht9pVylxX86LJP3zSwbyLx57qoKnQ5BAilOYZ6cp4DaHu2G3fixdzM
3499nq6kmWBKk5CsjyxLUdeeHJYESbbzHT4uk1uI3BvCwUCnezlQaBxm2Mf/
zmcZdQ36oMWdfUr0F2Ln3IuzbPIFXucg2j9Aw7Dnxja2xjsDyWLfwMBXe3X+
H/IMnu+FdQr3oYz6Y6/pN5tDybO6GWL91aQKdH8F9yx2As+ljfvZwCwE28pg
VSrWuvSKmUcLuo7H9EXWUnunqcdCP3jWH+XT1Pz//EOnWsqsvg1ItGUlCmxW
/WTJ3Vo7WykSdRnHWwFIde4H0jl7FM09OEAJLlk2vna9zpzRervvlhIB+Vc1
pLB80toLx4K36A7U4cB7abfqI9IvD6AcFXRY8KrYF1jfS1sGjQECfHfx8wjg
jnyt14qjgh3SddlDTdcIjIuEyy15QkKKpQgMvmKWXgCWm3PahBkLULbXuro+
t8nvCG6/NUC71UAGL/5eIC3w08TYl5hyX/CwvXWuJNEb02ZhtdtQOZ6S9hAK
hq3Eov+Cm6ihh3RelXm9MQ6ues7Aqxfvj5ebTuiC73e5T+52aACoqggF9H5r
SFZZl2HQrTSG5KuK1Wac7vHlnHqmAEk+X/eGXWllJ2JzYGMIn4jFLop0+4lJ
XIPcIQOqY0VmhYpQlepsOzknFpUysJkX8BGcCs8ObFB2OrOMNSiyYr+ZjZIo
vm0pftIxVVY4ReHtNlRaoM1R3+Ly6gOcLcSlyfmRqm+nUcaDw/5MHKG93wIn
u3+ZCHZdRqE5lyUCSQSD50aY+y027rEB4FhaWMiEF10PkuOw87hcn3zYTunc
J6uqFxDNKnty7UjokigAUNhGd/1q5HUuDaiqPghLIrZ+DxKWES/zQGJ5nOaj
hZzNgW5aCNnLIoEjKF0lIZz/GgJbtB0BWHqVsTponmEMlD60S1cArQRfjaeD
zBFpjW6psdIBxjmsqE51EzJBqXt1adJjQ8F+u8m0mYiTzFHp9HS4t+npypRC
dutLErFxZl7sdsidHAwyQX4lDexWmezxH2UvFokIU8z0Kx6D/GKy6HRtI3It
2BamisQKigW4bi38zEEenYYYRaUM+Nqx3pv0fU3Gk91tE9LAaSsBRF+NduXb
QEz9NIRts6utAcfV3EF6ZAvpKixCZ4IvadL1xLacDdgyxU3gFyr0w8XKy2t4
+XOIrVsaOx73AQq1IBAX9r7BqkaXI4xaXxh5wGJtp/hHN/JGev8HQDBGoYAn
XRBv/s1IV4LmjKBnqwQBiFbkUSvqDYDz90ebJCEdScuciLJJsv7YR4JowTQF
zl7Tibpf68dLefT7jUNQYS+WFX89ZmjjzXfZlwkemGXeAOVkwwQTos/iUiGi
PwTqzY/3RN0Yy9BTAQ4BwMekAKmS1h6CqGRHbH7vhQY94DCHiqLl5Eyd37Ie
SUeYTBMc99YpsYq9XrsDEzN4H+4UqstMrckdHNhAoVPxyv+B/VV7HIkuvmVc
TUBUnSqYQ/rFyRcvM1VMFdkiSQTqUb1jRaofqSzcsiY4HgrkiVzO506UxgE4
+Jq5x6qzlLkxD3od9pvqk7F6zAJYJ6un6d22tYpcd+E2tEQD7hleiMGBaB7r
JjtxIrKg7QSENOIhnwoHT5y0WiY+uLxNGOJSwV56ICNRUFJ2K4pvF+mGP1jO
k6lVU/o8eEH2iq6gIylWXF8xTBbzGcy7rtDRXhNQFVdpTdc2XxyrSzuHoR4y
D7RMDAsrNJCqeKr9+ZEp5iAMepS+wAIu9lU6VMmCw73SrJTIQ7MW8zut+rCJ
AF4f7dNLlPQfvu1S8eGQO4iBJ3F0RUioS7lbAYOmy4o0kqvIgj6leLS6FQsc
k4Ff0gTJm0n81+OBbVQLBTO5+lvMCzTGHLZ9AReqBeitgd6hAjanlWsBIpg1
K6CIzX5R/x99PV/zSi5l5gRO9y63DEbpwSWS4hLoxqe41u6JJT9WqUFKuEmx
81VtS2htk0apuCv1oRYK/7yisIymutfT4hQRTveYQQesrOEgKwFbdV9KDQk7
MRemvVXkhmKw9Dg6Bd4IhewfIPPlTONKfBYM8y1qDuMJhfEsH/x8T3H9jixN
OMONrz+o1Hs3FDXfkeBPDgyXDDisvPAiHt8n1YxTq8ZOx1Ua8Pkxj19yLFiP
Ql9tjf1yr5eWIR7t/SKUu8HB2laOLYqZ3o8g1xodkU+JSaklvGYfDT1SmvYF
Fh6EOeKsCMDOJtBbqZ1vVi2qCwyDAR1vKxjl6yi7EGxCLZhxoGQwhVwXmPjS
7INV4Rp9rgY8GmwViuV3yq9a8CpDGr+BVhK9D06kkeNo9nu44Qf2RqBqZx40
ZMGgdAHZOqvGxOFAARwRdbcFV82XbfDzbweWvMnRmd4qsJ1R3umZGzvo5aTU
jKpMkPanBBBH4QSmNedB9sSL5r3rS4oeJ8gXU05uyULTr9ffErUJi+4DnEQ3
1PPUqaaABaH6EtqbLiz4WYQRA+HPp4flBHEORSII8/fB744gZEjQ1XWifb8j
Xcx4i0Uprf/cjzvQUWrdhR68ZSwkpQzJGgukBpAoLCng9GDlPVQgvyB/SZBd
a7X8SVsA9eSQLQgTjgBohJTqtbm62hgrMt2V6XypOWGJ2hy4tnWJDqeq2PaS
V9Cj4uoXCGkV0mgxtJxwmVnwgKTSAB6Zw5MCSJ8dtQLR9gD+gHZkzEkQvyUG
PATC47XvqvuD74AISOnybTWGnhzEaWZJjemMDTxjpGndbgCnhn29+KBJFFZD
N8tQtCFSALF7nxh5LKG7R2mM50sLOb2pSrPDYhww+63U1qYJkpOlIPMkFzsY
EgCELRCWktkSDLLiZv8PUjgRhH26mQzwjcTYzWDrhiZW/Jrzg927GMZ1r6E+
dc9tyP/9JOiHHMGyB2I11XSXT0xNqsx8GsxNJPGAZOYvYe2iFuTW1lWWUStm
SVuT7vlhmekVoCfnQKcKzbd2f5hRNt8e0i+5IJW2clccVtRoL+PLWRXhUh4A
Jbb8qdp22jfpMlwBbGa2407qkcJhS+5Hd1D8N058ADN/klfnTeXDO5Rs3LH7
m3Gu9NzkM/RhiFN55XqYijTnteuW2u5KmXzr7OxSwvMmLebIjgrbZMQWxWIC
ATp3GdujSq+UD0MqZVOAasDDouhkmrFQHqDpwj4InV7xAAhbwPGYoUWP/uVe
3UXo3pK/AkIKcJgsqE/HCkp972vouhDUNoNQfAsgAkb/F7F8IFaC+QwaI633
iv4vDEJEm8BPtxtEGbPU0j52CeAx48r4/Dh0WdicBWfdIkfGcbL9pbllOPze
wupj8rjQ30UNWn/Fx2UQ2d6JG2B54VeC2DPNgoVsKf8215G5LfIrAJ1nGQk7
7XfqC2IVySxq7Voz0RJ62v/2lk+GtCEU+mw4na8vl2iURH1RDn9IMnXuRN6Q
5NZjn1P9Uaq8EcyPgA0DsyXRHy5XGpER5NgavfqslcVAWQAw0RLmMtwM0Dop
T8/Ra8RLRsnn//WRn3DSn609KzjYe84nC6R966no2xwGLxYtecvocJT9zDOF
cPFanKR3sw/0RGYgt1vfwCej/JEorfSxWCGPc4RBvc77ElkDjePOG9XbGDX7
rz0zsUISsHTq+O6ghzRIWS4t8LpWBP7Bza1LGKuNmfQrxSc5j1s1dPtBb7aL
wo0gEWgun8fIBi9IieHJvVMarx/EpOx0AymusLbix/izZ7vTRYDAaXHVt8ky
6olyJ1wgn61K8fl0E2m8derueAxdApO4M9/FSAMxSmkZ9p1XaEvw/jiuCGfR
9z//K3XIzURptCZSXA/OFoSbFBJdqnNKao5z5EUhViIsYn3++kLO9g2llBfq
ZME0EOQZsGMEl3NHsA3ENsqzgifFOfEQPbdbb6csdrfNy2vfS+e4B1jIk7OP
4qVSMf2j1yxeja5muMxBMxRo0CGC4/l+w0KqSSdgBmuPKZGV9wQ0LkIwRHXr
a2ga24bxCBilXf6HyBhlUZTzTAGcYC5uaSF9uOXak0WZajfjI6mMR2rZ099i
Ri3AkmNYjLZgs5s/ZEAeqkz355wckLigY1tHH9tGTm6htxg72iOKxpHIK/8F
dNzkjW7Pcs41FlGplsyLl+eXfn4NJIx3h184gd/sqWqGSvQjBQqa9iil+dn0
HpXReTjgHSVTL3AzOC2yXZdbmfCKPHOiwZPivGP8gZZcJy9xe2nMwKWE5yIK
ItKI7pH92sJbHglyJQ5BoTyYnwKPEzINMuVjeS17U88jN9symBgMECBr7Zle
qHPFxK1DXhZtWyhyFUSZ22I8GL8pGO24Wf9WI8MyPdhDh9CeA6BaQy1oarSf
z5pOec676eaOx1gGNR0EcDBki3ovw19OnF3TPLBQN7U6ORSRlHgGNnjOuZUm
n8eZOa1zTiarypwQ1hSh6eT79JkoFT9QbY5boqZYsYrgG06GYag1e6FAjqhM
ZKgvXMeJFmFl4pvK7CYYQMt1AQJ/DyXne3JbvRBSsOyQLcEOVMCApSEw1RSN
5J3OnhN1Qbdj2OnXlVzeVYtnfky9iUkRu90CZeNfhowUs/+FB6YMkQJrl5p3
O+Os1XJLOwxUCb9aPNiupdfsuy7Wr5GTAI86bLtp6mmU6vV41aE7JCcVKTGx
Ob7523sVldPodtwwzH3TDxHhbZEsdebRL55z7jm75/UTd5wBQADHQNG4py2N
CC4US9r+gOe+OSWjBTbdsSzk+9AO1r9nqubRkLqE0dkVnLXFTan7txDnDd0b
kh1zV/3LERQjcOZWR0oQcOIPvtRxiqlroWZ9yu+9kBuHEugBopRsBJldq/vS
CF4cGtsC/buC8brvj+wN/ooNF0MXcrbXGNvbt/i+V5zsXjBrmXyFi5WS/FK4
3NnGaFNwBgtHkbuEUMYRnv74D9+P1WS0ICo/TdIFiC9MSPiVwk5Vd31Y49xz
6MgZUCnyKN1AiJqqqfFBx9yeJeGPJn7JA0Ky87YAEcHY5WSaVubC/fKG3tx+
DuKVfRJedTtj7RrH6SV8HbdlowwjFcJsVaRvW5ha72rndn5KmqZkw8vL2J/w
yVdS7lURJOlvK06bB3aMPBcUOlYWLEAB1H/7R/7SLqbhd655tPsQnv6ZGeyu
/LsPMkhY0iCjK2FeTe6Xu1trbrMXLZmo2NP4yU496WP1LPmPBC/W9BMbCt8H
g/SlhQ6bCK5YKpSX1ZglDygA1yTdi24VakEGjWTXVKazANOeuDYeD+UoOsga
j8b/M0/Vezgfb9x64bU6sHR1kP5jxmf0LnpN3kfjHaq0KAOpRKMw5xvP05wY
EJkf3s4629Vh3eSqTCs1uzmaLJcQSO2OS6YwNtJw6GrvDUkGHvyxePd9+0Mx
uHrzKoSzoa+JzdfMnqat4B/bfN28NbmqEB9LDTTV/PgN+XX/gi8Jy2TlRV3C
z5ZeUoLeTQvb2owa1+OLSTc32cHqtmuKJlBZNfh1hLgRjFEoLQxhQOanDHqX
noJkeNMZyzSbL5AI33+PjBVdLNVc4xIZSL3So6r3ym+8MYAT4nLYdldQlOx6
mZ3t+UtW8kPfS1PUGY5QUm6BFon0YlGSE0csZIXxmHBtT0tvCVLcKu7pk4iL
3S7mSanfunOnzwP8aLkE0kQ4vVvotm/IJFZuELXGtCnsCrR+/HI7hiLL4Q+T
1h1Glzz/zdJ0D+FaYt5RrYFyMJ7r9397y2GdG4CwoDINkai3Lyl8KJEN4Apg
L8ER1GrNUyC69IkpVROKLz1Bv+3DUAV8cv653YGh4fUgfeKh/WT0vOKmYal+
991IijxZTtIOkHY9SmPx8Sdj04Br81lCRCj6d6jibFO/drZF/RWUdmulGP2n
Vs/2icrW+CgzDuLXfchA5+twPg0xuG+JytiaL7lQXa/wD/mZus1luygjLeSU
mitSQmWPF3rrByqLe1DEX8lgVPOYTCLEkZqjTVV7wEDhU9GcOrkljrGZTpqE
A29t1PeuOi3xpUlsmQcOmt8DABzTwFvKf4Pmxj4PocgpRdG4GW1RDaoC+yQ9
eU209CZkov1bx2lGWEnHbw3pWK36fVcP4YSsBe+vJioeNHswR02svq0NMmeF
+fVNJefv3pIZPWIPsrXctnuf7mdwyjcjWEGAUOyV6U6ReWVIWrIdsRxPlAc7
JUZEx1cZIXoi2QNoy/C92OsGqSMdleAGHDiP3/JFOPkdFWNH4gGCl25j4TrK
idOi6HvG2RktYmyxj6ymzK/owgWNbTGwxBmNls1Pjf6dAB3J+tYIE78Tcdkc
ZcwAJTCfYIQnTK9k0nP6S1V+m4cA5xbMSZF8IjZWpPHn1FVLpWra6fBHYVPh
BD62ktD96RJjS68H2eL+OMYaW5sMBQYVvAGTImJtX4IhMlxCL/Oa/DtnbvEa
qDemnRFhmDgi7cUFIwKElm8yDGRal1oRge7gDZ+JcrQskGkOEM5NVZHyeHWU
GncAQH2YSHaHFUkzv+vYmQPwkb2DEUYnAMYtTAlHuDJiWRzx4Jiymi59owI9
94PA3lLO8yAnrQef7gkIUdDURTUdK2SvL1nMgSECzwDuvNGeQmfrHs42lwlq
/Pd/prpdE4LLBIHFWicxJginYBAgpiIs2kJs2r5lfFE4GA39ZdEpd5RjKNmJ
yI6iZ23Y3gjJ3xZAsPNg01MvW8vAxGU3DDj96fl6/zH6ckbLJARb/irK0OyK
rmcY2GrJ+CyJXldP5nJ8iPxwrfqCRvGoZ8y6DA7v6/cBSlN1FAggKaGZyd9r
PhIsEQJ1Hk4V9fjFhuwXT0ho4y6DJiIhuJ3mkwn2bG/fUYyBHm8LJVlj3Jxq
Arg8Ufz0gecDARsRpIc+CFPUurkv4QZMWcz2dwox2y9lFEQUEfOtet+L84pp
Bku2V4Ji1kKqZwIwl4gLqo3o8EIY08L5skiU+eMoPddbRYa2/PWIrY041x1Q
h7hlfK68sJt8notNUoupTJpXlgnHNp4HnfSdiAwpVI1x3QL5ZbZlpbfeQGA7
2/FGWI73nAKR/TwehenRIEyHR4UMhufWUwxWOf4tq8BZRuhS7e4wRLR9xDcG
vbKMd+76mAf3EhdCa1IGvCyzVpqPQyzfP7oly+pE5AkVc5xVkMFzIU/p3zvs
rpAcfOiAQ1yXA9XLcKqFFn0VD1AxsmpM1HddccdYgzGyxIsMWCPswHoBV80a
B4SGUy+JUyn6ZdOkQmPv824Ogm4dUd0NnEsU//3ZKbdKw45pcuPWp/7cpgXv
NyHgClhGq9Ov66p3WVidj4c4qdVvAN/qFkU6qnG2mgcBzKNRYyawdaYPvVS6
lnC/uVyI410V8Sg5SykTaVfHj4G1nBzNImsV0wqNwBEKxhj9hgH89/hrnO6K
gCyQhi6p82lLKuQyovlJVNW3pBcTTC05sYZvsGWM5w9ucTKEf53X9LdhEDny
I0k0GG9EHzDXCrGH7uFRx095hUneBtgzM2ev87OjTdBnivZO2jPFoLbJAOG3
7Hvha56fWcnKlZ1+ZuYW+87va6+WaIB+yIskzhnqyRDxL78XPxD8N7hqpvVf
qF99l3OBMKxSL1nXk5JSeahy87MivNDfvAR0OVec7i4AKu7a0FcPomRwBuzy
IGu9+Boyzh/W3Z8exkOAvkwHsBUe1yzpClvV92kCmC098CEPHSB7V4y8/9/c
m27R4qN0QEGmSmFVzv4PUdpTQoknvOifhFEHAhR9jnHWCGELF0ezh9dOdn2r
subxRS8YtyXEM45KL3gXvc6/mBpNk7N7DuBbD8SMyznO8DGor7d+lRb05nWb
hTyxVisMznzY4PsUrdJ1vtfQ7AXQpFxN6tzawFR6XxDdNwV73TgxgublL0by
Tu8KL3+xs9xDGLXjG9FyjUAyArwWAEHtykBiTPde2VrEAXBf3e9OuNougiC0
hRWBIfmPFovTR0cXM70/I7+UQK4i1ADBe94NeU+nzJxUGeQpwXl7L8sZdkMk
4J8mfdijIyymDOMGh813hFsEHaow8/t1lO4M1y2TL9pR3WL5H9pXHGaD42BE
+qQgo/Hlqe0ubNbbx5IGcvSXplphiBFsSgIFp7Lsw/6Qx0o2NYE/8tej7c9N
l1BgWWiAfsWODans15k9hOrqsaTxCkmh0IXhpIReKqNigaygei6I/yOkXxsm
dWlK8XDmrjQx3+UPnCsPYEbfbqQWqjIMeZPbk8UrCLxuyUynCmKv14dS6DlW
65BJsUuLJYtEHEejDnTsVcHfyNYPICHIR18Yh/PA+PLv0ZbTDNwqT7/AZ18D
nQjdiX8QIwk3LxFXExVW7OI5FkH5q8SUYHqrUiINWJEyS5pVPikZw9sAB3yE
Rp63SI7yUvuVsKH4IV2CaJMsd57xDjMfOZt5HEhro/h9J/SjYeTxetuMTuHx
UoTdwNGQii9kHM+sPt0HP6FLKLs6jGvvlt6SlAFUk+p+jw0N0sofDhYOUnz5
+7EvIj1trprIREkfiJOQzY+IFPdmucGhPf6678+yqNwTbQnFzJ5YvyeuZWJE
1tcWXtAA22PZDI2aa7Kl2DGf1dUi2VXdXH8OG5+Gv3G+/HIYwc1QL+iTNIf9
Ym+K1hH/j7pgwQRKVJPNTNAz9BXB+bNsMdv7/sfMh2L7tD1Ps7TRRfD8cKjz
R5Jo8wBa0GA/o7FVpLBSnCJmbbx0LK0QkP/u1FlVQPH3TOl1maiKKymQrIbu
F7fmg6f41OKCTmv1qNacaChfuAa3ycdlbONgbVSV4V5xCr5KKATFbXOXArYS
HvFe7MpKD80ZCcGrQKW23msTCfaNPslrjsMgBXFmJau2fGFZOLGsMnPUHRb3
/CUdYvvETiJbJO/TW2Fw8yP3yE0YONYChNWn+HHrMbcZXA/7NG6I9uCg5Jrp
1suf1VHsAUilWkPrYx/h5VQt428yzc5x5BBjqga+/+rt+pH0EKtp/c2dOAGS
VmJn1tjRTAI0DQ8YWWT/5V+gUIEpvlxKhN/mV1rMqW4H+IbEzPs0dqB8fxl8
dxmR8oeLsN7co49TSiG5FEzRZ6ktqJdjemAr2NtJXXRlsQwl7OIVVJrNSrwU
SRLNCHd+DeqIgzYvunPqNkQQeYSWkIgoxTrgCklMJlwI7WoiltkD42YZABer
vEmupHKgGuub8NiJx4fY0X84uD1QoBbrvHeGKym/RQstAThAl5tHSJ77HKzZ
sccD+uBBqLz3QC5gAvKRTt+egGjb7wFxuKvhJQjIwQw/HfK6X9kHpn51kZm6
6eJ82fxa67a9yYQTAb/lQrh39xvAWHRon2cyrvXV/TfIWzh/N/pfukHVNbw7
6Szy8kcL329EVBUYJtrOM/xbMpeCRb14RUEIzw9jPY3QJUsGXu7Tv30v5oq3
+U8gYCBWpsHlfykNsAYBhdjYmSllKZ8vHydUe7PTtDm/GcuaMOxGZbN6tf8u
PyEqTeiZqPqUC4gW9N8uIj88w5dl7TPcXWrPVrFBrnz1fpM5wYPl46f8q9az
5wF1Q/e2voC0/H5kxl0U1KzYX9i4aL40SIiVrlfVDk2TMuULUP8fb4nkTXg+
ptAk6mqzrTF4UFhOAW7JWeBHcG6KZ0NUsWHkNuJhaTRuK0dVeGdPdA5NxVNI
so0263HRhoK6mKIGw+0KNCky6cvfTDn0L21oDuUtwhrVdNpHuQx8rvfdY3VL
HAVZXH6UMqQGKrhbs6wBZV8rm1VMuq0ATuOAz2xxOU3GKIcWLJQxupdSWpSn
qFX+ZLxs7fQJyfmFZ55/OrJPFLP0lrPxcOImDKJl8pN40tGt3YaoDAMgk4td
B8Jh+oxt7vAzJJTSGMtA8k3MzQqCX1p3Az6laaqi/qy2Kcr5eplF/Zj766iB
V9FERaKl+bL+lTXOuZ42Ovd4aq5lccoZ3ImYEvYqEpjMXPLByUuZaJsStMaS
vPC1HcBQUEe5oCp49KyTU7s6vXmXWE79TBB1qZzRl7zNcFN02M50GdwGsuGR
Yc/XOogERJGFxIA3kK1Xo6UVie7byY4u3BXLB/gmLlnQTGzopVDH+fl07jzV
vsg4L4AGVbw+dpdEctIKKrTmHrJ81558dDBI8IAERBq4hZGBwsGb/d+AeUQp
kV4dY3dTo9T9pmYO95ECJDY+E4rfOMxYIwMyT0vgWSeROv5Q4qcsdKiOQgSs
XH8NtcBtdidzUPHmqlk87rCuhCHGMk+TdgGoGa74LvJyNF88CqB8Q7/5BUfe
MbGhlYKU9pL8BOGOUmSAbzreZk1dWiqiXRNYwkF0ZxQ7fUEdY91WWR0Wya4W
yRFQyDVKJ4GRDCK4MUQ3383d7+djMomK8IxfXaYL09BErTiM5k7s3ZBmzc+p
k7GNhsaneXCorT0Kdi2JRsC4NzZKxZ9P7mkoG0zrswIYGQBCvxynPoUUJ/vP
ZAm2XqqiyEoknUR2xmxj1MlS5fWGaLgDT8z4Pu70BgZ7okZ3C3vtScX/sbUl
UI6mZX7YY+UkMsah2iuCjQQ2btAVPcY4HQZ4Lr3hG6DozE8GgUlR3n+SLBJq
pNSkx4YToJShqcNUeadYdZhFbJjGFGvuwboXDrbFpUqhHt1NbxhS6LIGo24S
/+dDT06/N3jyJBP1baEfUvuiW2T4+ACpcGDvNDUc6juxBkI2EO3vUsgV8KGH
PULJ9Bto7fuyeVwyZkjai9dCE5H/wrrCcG9zigYZgx/R6YJM5RnxHBeZzIb4
vfe2rYTccF0/sNqq3Awfo/vib6wOlyf3v+GG4jLD6M2jMZUOGBkfneLf2Ix0
EvRBPjUFdvEDh1XSbZnK16nrHATs22gS0PK3f3R7dF0KbxW93FkS9nwd34Hi
D2SnhGOop5A4t2NTNXqqZOpxpspRARF40nvU0Srfw+jwWdwrfMe6hiHS3GjD
wN7kyPB4uNNpIDFlokKqCoEQZcPdO4hcRb6rMP5EKhyxGsXS6ZFlT5Od7N/J
ZJn+ULEf3znPl8z9tqx5fOHrhne/AnKAE+oqKIo97Mc6TYEh3npXqFumKA+k
Fn8DpFbVqA5FoLmdpAJKJaJctVx0k1cHaat4aGBTpDYCBjpMm9C64CBjR6Xy
BfpEwwePFBqFyU+T+7e6IK5211Lw6SM8M7cbkXLId0z2yNAsSBVz+QGpIw6/
1Dm0H1T1p0wHf3xVBjpRtvVgljYhgT3AKnOmdyzmmLJzbxH+K2c3IKL4PjHf
ggpUo9+pJAjIwQ+czy55ZwYjztX5jfITbpoobPo9V5WloP+s4A1cqauBAg7J
vhYrjK6bdoK8C5xwnMmazd9YU9AKWjjNWUR6h3BZk80Ql9YbSZNT2ExVVGUg
n7CElaF8uLPlFRFm8gpnTqEYFZOiI2b/QztYA+EsRtLo+vKFcWT5m2+EWCIu
MtZ6apB7sWytFp5qDw5/bzZhNsk6URpgg8knVW1bJaJm9SWO4NKC8ap6KBYt
Dv8TKec8wEWJ71iXQ99T290nT7VogJpHSza3nq7GSqX8wmtWSEnck0dSv+xN
a2DFa708EMEm2OsFm7WPMtOcM1i2E3Z/KIgRbpKtmHxiM/XIZwsKwVMHZio6
Kioj7VX0XzIdo1fnuFtQq13d48j1RGgH7TwUzDlyBxSfes/qhQXV5/8n5RS7
c6vlcRYfH0m3KYqNPsSZNul78NOP8bZUFieY1OyqOxprhSK1su8sqK+wbgW3
5KdnPo+yUk7dxtETb14Ha5X0dN9CW+LH759rAWSjgtjod1DhwAYxoTPMkmMH
u/2fjzubuIGKrrSIRCIGFGLqJ1aaxdA5q4fH8LyvyVN00o4TbItx33ZgcTHc
d1PSoTRMJYw6XOsftncEqOqPiojQfYhGP7iMgFzKm2QpGMUPYQU4IGtNstXp
+PxK6ZyKMvsW4rBSPTEgBknkeyiRKwJ1ihNOwRmICK1HWZRddclq2eu/909w
kWeL1pkJWjmfyrSEcuymy5ZC2J1pxpCVonaQHqqA0QCser+QIsoJujFPIfvq
2hpjWhcL/3XSziHhn0yMI6FFnwIEUyER830Qkggs3msJXCIVg2e9T8djFroy
2yDGkUz24qvGIDLrOfIoeu30eQRJwmvCRsvXtRpVkoM9yQ1IruacHTHZg6Pd
LfWZhiEWxQBtycNiUfCHt+LBP+71K7nop4ZhEe5Jc0uD6Egr2KwpvUnA6d4R
6+xkReYLVX5xzV4TNRgHhqFcXZcZycWcUkTBUq7r1oukq/jf4gLweCJlZcyV
WoXMk2y39YpfLN/eFGO//PgXhlLtlDAqLfiThMshShO+15Z+cJx1Q4LTRlpy
XxGC5+q3Ik0IEAjG6OheSOOrQRpkzGyeRvl9uvIl8KBgdjNXK8ksRvIPjSAz
MsiS7XOANalkBEcHugzK9pl8IFheF2rWicR5UuSVjoEJ94C0gjV/61nqmvDB
kDUNZuJLKw2tj5weYDFaJyHQj+pJdzJixUKe464PNlWXRsTvVcYpzBtQSSpZ
LvJiC1OtzFCZY1znBNgOHOmMaMePRojleZuztYvlqzR23L5a3ZPgjJgkIGc4
GmZhJ1dQXlP5lV/xIfc5OX0pRoHZ2ihOBE3ZVN1SgJfUDL57exnMh+Qd08/S
/7Hh0GHDMpVEL00lQAREvNlmqUIVC9txSA8QgOG+uYWvfNxNUXgndNwSenSx
tfyX07DsBGz44o1YMZzCSYJ3Nq+KskUsqI6QmNKUlHQ73smGlz8kg5wB2HRm
cGjKW4YJ1Y9WFAuTCbBa+FCt+XslHzP46TYe8sdGFxVMmhOSGRDgxptZlMwR
yT5YYQqxEZW4XXvOFGlP4kQcgyxCHIlhdyNj9V+lLsS1Q8PumltI7EhkpuZs
IgeGdea5bZJXkMO/b+fiCWA3MLCmuD7jAbGH2QwLRlm8v9w11MieLbCUK0lY
/Vb6GYLHvDR3DXhQ/RvPxKEkcRfL2movh71V8ZSF0sQ2qKR2CyWiYYjaIoga
eCiY6AiduZxLc8PTtZxvSeVrxU1fdpna9vtPvI1xpWakjvNmwuj7/INTa/y/
JVw10yxxCSltZB6VHwt5QcdzfH139nqcoPks+YHuj/f5CsYzstM6/NDX49U9
DA9cf1EoHCmRo0shTzoDi20j3ooDl9Tny4CYYwZ3RHf86Z4w53/2Rz1i2ku2
QKqjovI2WNgEP3fMXhZ9+W5BClJemTt2kBZOIG+azoyunF5S3L11oP4o4wuB
tpP46e6eppKfvw7oV1Om/ra1drhSKJlVGwsOK/vGcGGe4HEx5cXWAo3NArRI
55Uc1g8n3Khn7XU0oL86JtTo5Xnh7g+04nL0cZq1SGHbbgAYD0GLPNNTYESv
esDqrA73W/L+pzSBbAjS+Dt8oVu8Jk9eXdtrCZuxW2FCEBzFBJuxa+m+4WOm
dAuUOpuJ6C/lIHj6/V86IKBKcZomeUuEdWSkTlZVSSBqvuS/bwIBAVP00Zwb
oTYslB4Lpu2OLXjgLiibEjW088BTzmeOyaffTlLCi7yZNOhLnS7v3W1Il0nR
we5y6MeFfb23Lg7g5IfLWLDqPozAEjyGlaHAdKTCjlQjvUhwtfDHxZmJ9bht
1PFRPNP1YS07KSpHPzOTT1JGDISExOocFVSgzWMC6psBju8tL/OhltI8SSEL
QQxKGsVLZ7p1EfVcjRZ+8lWvLbLJWcQXbfFHtbsV9vWbIgnEo8+fRzGxv8+a
Spp/K7RuBrUBFgk3WvUxwAm+tswSC1oKoQlyrXFy3WvJte6Fi9mVGIe/XbnF
ze15myH0hwa2A8J4wfo4IbAU5N1qptyEIucFbSyMQbeamEjIlUS2AqCVt9PH
0Jsx3VM+vghuBEq3x/JktDZGLqnLtFF6WLB75uvxjInQ6QJ20ycBqaCsvjB0
mYyDfQiNz/P8ejiR3TYUXlIUz8/HoKiEvkuSzvVYCuu1HNOXLk77ez90pEa2
aHfgEHIDJ52+bTDxtRpWSdxP2E6NQ244ag96/g0mxhkhb3UWeiB7ytDYIiHf
oVdRfjBSKG8YtdSRL3AhEMTklhSSgXWJ0mv6H46GA34uEZOOQSmUJpOZ652r
Mdr+2GVzTcH1HhqHYQeH1hLMr69GysEbSoWWFUzrTqC3ExEX/SWASqBtrLY2
7UcZLImDuQoyFAOw0yZrpBJqr64dzp+goQMYhWGNKUmK/I2BvDM2zNY5IZrY
HPY4YEM1foLoo4PXgsbX7ShhWUdg9PEWqmmqqiJbV+FGA/7+ARGFuedpGNim
MfUW1/hrWyZcmC57GKNhONb3N9bw/LSb0yGs4ZmF4roiwLhmnQTAT1QhCD1k
d5oMzyYu8R2pi50aCDi7OsEh7041wDGGIg8IxE+Qp2IbEgfYHD8XO3PQiq49
vXF5pjtz/c3b/6GNVMGL8mvJ0HcCTMwYAHvI4baFnfV5ExnUF7HLsb91zZlo
/ZmhzXthFL23HmyeqnKbC9UmsRQRPjBHIS+6fB6ll4rbugLgPPRc/NaMhTcB
WGcZJlrn+jCsrlb3IpsMlYoPB0NJjL2hTXIBDkLOaM0TnHDmu0fZH0AflkKe
9VkTpMI3piIY0zWAKhBJB2oRbHzudpuU9x2YE4/HXpSaWtYQQUyZ9TjIj6/v
KJO0jhW6C44KjagAqEp9FHMF2cKDXw6sxHNmC9FykJTpyuLP7DJ1F3nBn0fl
cRIHVHN/D8OeEQSg9LAmn5VY/IogIQYNhR8yse02iWXs3Gb/r1zpDV7uaCos
BvGw5w7ytezb08VwSuZh2HIReOKyzwT894YFI/EYT+CcrTABwfHekfSRemPy
+bgpPo+OSffcltSALVSsKC1WsxxHoJCC6R1zu5ljmjG5+0QczitImSmFs7OW
7Bk/IupoJcmZ4pvL78DVpJoD8YLnf916IURsmLpf4PhuNel1DEbSQPFZWx6t
2EmEIm3yw9o9u1cZaTb2c6fdGdQBxgEp5HIq0/QGw7WOHwrXFeGrx1Ufh4Gw
sWZLpkuyGxq++nV56JP7piqXia4JNMN2sWJ5yKcNf+t/w/x+ar8uRTFOeivd
MwiQ4fgb2WuAk4BopAVSN6fiY8AgDFPOVjvlPuynmwmYnK78dePDWOQLXDLU
jNMRKV77R6gnd0r75N4j2tHN5UmqshSEW0J5zPzI8OBsWZvu2vfnwECjMYNX
EwPnpOTXcm90v9URkkTizy8CMDOg2gl3qli8FrOh+S7pd6y3wq2fdTHKa/Xz
KUbkmkdFH96W58sEW6UqTJhSeFIryJX2GpXy5skR8SyggddkmoLrLf2N+u/m
OHoGb4a9rKLyKctlDzB1G31y1efb/xGLCnYkVSdw/QuwlqM5tzgGfnIFMslb
zufTunHZPrq3tSUtmeen5jmLmg+Jhg1nmYcu54EnEScDhf+edMaEWOEF2bak
jGQPgNTt61irSqbAL3kxrlh797UWQOOqQphNdB+iHuxgAixH8qyxNLJIVP0g
7BAon3/69mA6XXozk8vX4M2FqQWbY19/AqXhElZRQh5UKBovQL+/Qaw2dt4g
fMXsCoLu37pOK3glwFWl+TQfbNno7vbH19xLGLgyZrQxme/bNj4apE1UlKF1
2j/OpC3kVRC5ANYhhQBQ9HvgOBKmm9bcOWsVZzjY6aecLLJaj6KEgezLXh8K
Zq//VUGFtJ6vNorkB8E14MifwxX5N8cBXyIzItJvoPwboQ+pfM3gDCNlaix5
H0d0UKeDyHCsZ2gHw/0HEuBnS7dU2LvASbXuDXx/YRfwLLbRfFZrMZsoOnlt
di0JW/h6p7hJNdTzmKFnBhYHDpOQnT+p0x1tT6zFpB+TTXvQNqqwZGGIOKcG
wCEDSP8I+ZxnCoixCSliyaY0xlCLQuyBUEJe8OA95I6VgU4qPBhuZIqskv+y
a0ZBk/LgtKKZNosgKiEhsbGPF5x4nk2wBWMD3+qviJ8nDVn+JAoM7Yx69WVI
Xa4etC7KRjQfAkmCO4yQgyfn32uSNRsEeAkMVP5ruiWdBjkJ/ps3Nq4YGwjh
Zf2EqOGCMFRzXPbOunZASIc/gJOWVv4UVRXk0xMcUEjb7rylQSzd7QguuuIW
ROaE3WUI+ZYCTfX71kKQDMI7TKX55fDUZV//vUUEk6vB4DKkfFl7Y32b9Twx
DVKXGw9sGT6mvQ28KOiYC9+GRr0/F5f/aY1bEr65PQVN8ezD+U0ZgxdiKVnX
w0bbM9QS3HI2TYi4zsA4rHt0nnKjkaVy9cAR33cbfMabPMYzyzUkvTtcY5oV
IdEQF1clZcTnIiICa7rMfykOVmJHBfOMvPToxjBf26ZbBHcuK/OIXqhqWy/0
Ul9RHRTD2VlwWzlFFrEc3Viu87ZastSOaH4f7gwtyJGx3eXKn5tFN3m+mbxp
7MR4oj+IjAzG6T5TNlP4nO5Ucuobt6/r42cAf8IglkINWLlq8rL+maYfrfXo
ACjxxxnhlh0tYpDnVFZ7Ss/7GQyI3oSdYtpmjwrV8C5e3nGdsi3NFXq2cxVC
xTFmIbX06hw35FzyMkp7zs37EYibzH1FGdM3XqlnqAbWbFfzfMQwexNT545y
ssiSlXLYeyobM1gzj/f8KnYP/8GLZxpwAwY60rwn+aJ5ewItMm8Nyd/BUbMS
pCMGQ6ejQ20PR9QL2DDu9mkNe9A21FsJbaOq7u1gkNhBFvif/McJ2jmRL5vs
RT5gs+ZN8XMX+qJjj1da7t7BQiztdgw+1DjBqOAZOy3hvdr1BuX1lPWb5cIB
Qt2EJMeE4u5UJG45L1aBug6S+ObkUg0nohetrBVcuRBbRTPV4fQKyjBGRKds
dpIoqz5WdwCmf0stkzcPeIyhxYy4+e62c4fYlzE+Nmxmu2Y9bKxyOe/4dfZt
8AIfxnkGX9Xy1Jxh+S++Ga7cCecvUEaJmlLTdfSFHLFZllAe6fPcER4YvDvq
FmTXrzv0WScv2v4JSeR+qPxrk6TjM8rceetNfd2irlS1JVs9G9RQty6kFUvc
6dKnaz04Uh294FR0g+aO966efanIObTBeKMIBuO1zNhqaYaAQfEwK1lo6YmG
EpHJL+8Y1SDYyRz+QeyGUWvL+zXohW3IsllZjBbygwB7A97D6oyt4zSsq2AS
tcnwmBjScXIIqiPBnpRcp49NoEJVQGYJHFfYiwy9XRWU30CLt9z6wqzSA7K1
zx+kFIMG4rjHrjmpe/cwn4sLehG8eI3C755xDVOZ3rJI/S3OlmwsgB02EIRm
dQThfFwjrGO7obdg06tMnoidH5iseLko0MGz6AFJ1REDKP7lw+BWUg+BumSF
dtdnObop1Z+kc5rzcxfvmIpNrcIhVrbU2PrndtKk+Anw0P9GxT1RoJCMHnFo
QB5o5jFawQ6KYCthI3vOJ2NZJL8If2hVZVA+vEjloEy/SPml13N++uYDIFrZ
pxbw7yxBJBe23jvpe+2jKXAX6m4ydIzalttVUv6cds2k+C3qrMlShreBYO/J
XKD5mNUEd3KZH7zxk/tsTBgDMsJUfycPXN6PmieIJGpbuTwWO23pMIIyVZvq
8mUu6+PR/wHS0oSJekYkEkT+8NU79E7YLdY0tJ7jrzCEZD8flc5ToAjuqtxJ
sw46YXVwZzBOhQ4bJctzCB5DfjnPa5K0f1LLO6hB3MoyffljhnqdCfaDJhfL
YHVktZtAQcwiV70fSlF0h/ueIze0pHhnQ7M7CsR0+VFVtEq+m4iP/9RfZMyG
GpT6lpHmgopmh0/FNaiI8eIlCrlAwNL1SSaEzzr/EbPPV/HR5Bj9+hofNlpB
X4JY7R9egDpOz28yHyOBzokkLW3uJEFUwFCBNry8nfjCq4Ql52SbD+Dz21GB
5u3wnsZJmImKTBeDTnKrsTp5tcNYeB2P6Ej+nMv5NF6Uv/fdZt+Vu8K5boA/
WxQHIDfxE5xLWbeUZkSE7s7GhWekRtn7wrJ3KpKojz0Y2CYDWRXpYvvEcqfE
ROpKCHbxP49UWDlAUDQcT9A/9YJi7J3e3Xj531Xs2lGuZUQqG07Jx9D2CmGY
YHseeu4CEwb/3K9YW2g9P0Hh4ykcehmNEdH2CJ3/QCOaNl20pPBYMvqYnH3A
MgV72iYgmQRP4RzmfrloRC51P6pgGqfLFm2pYGNvFavubVZsHoCi34IpT9WW
9xpGGM1Z0zKHSQ7/N/tISc5kZgzHnlfhXJn/31hlGAYF8107Ao/HFtE/g44j
QLTeixQBKTIAxvOf+DUTWVFANqzG8iVaWM5mEdh9Bnbi4f0SbArCPl/uSFMV
bXKD4VBcEtjuIMLiDiCvMnnOdc5mKRQmmkgVnctA1tK6x7xdq1HrNm4iON3X
T6lz1POUB83fIdJR3uBuD169/ljNKVeo2Uxx91Vfmrr1PNV56T04XoRDEHQv
Qsgl2EH/bbjA6588/xmD/bsAAphWrGHCz8p+GcGpO+MzzD+Z+O5WkKoRhBdi
ONdlHlTwMbp4E5gALKYWyt6C27g/bPTABEenThosFSX1HbGt2FuWa1YylaWG
o5vPjssT5HYXDAsc5sP4c3G97AqWdb4w8/4qp9Ys+ipcs6RSXSjVzr/76vIy
/NS5G4BDjFsyqX+0bGpdA6sMRR55ppZ0YcDPf+OLU+Pp4XMmrKcHzMwE6GJi
qhbzag3jmaZSdv3WHjY3Tmj8yye1dE4HuvOIzlDJRF9mM4z6kSwZRaPqH/WL
nXFHeB9H1KR4Ywli9HPeMCMJ77jEOXfJw5MmwAP6vFLj4p0ozVgmlPiHUXvT
n4tAqr3Zy73HxNTnEN3o+bzWKdZ+WhjH7Ml5/UIPDHq7d7yG+fWl0l+wr7yL
3fs7LturI01fAZH9X5AQcAbJ92B2KEYhbc24F9k/SsOqqnN6bA6N0PBZvyHC
t4ZF7TU6lNclrKvL7uBp1NQ52j5ND8RkqM8W25il/fiaYK25wVhfuNdEaumX
uAfg+Q3ZyXnLvXr55fHeWrfoHWMZEkAdLjVkZ5ryTCESjBAzNJFWlyM8lfmm
hrrndpATIrETNjzu8JIeSOUf6ctelFdweUN3rEaGjqOIy3PU+BeS8DgbuMwP
8VOb3fC8zdtlyJEGhQK8HB/H5v1saHetnIKwN3nxKqibyw7KP0ZOOBm4/J/K
uvNlOP6AHmbqpLGB/VKOGy+oVJi9pNLojea8BJbeSxlu+1X/Kw1f+fHSFy9w
KohOR0ntVX2fKPjnBj8jB9OmHgEuSvB3f6Xk5ciqBM9yVrUa+4CSiV2eOSJk
e23fufVuxPPNHTeOFPpNonryoHE+nNtKneCpdDmI4W71qMDzikAw9TJOEkQM
glFLnhc15OrkWnli7ZlmXsxLLT81payH2sUybSwkbPSe0aWu+T5H/Q2OsW24
TngDX8hQ65eKDGvC3HGeM/3o7MeFjG6ybuh8EJkmrXzRdSQiSNtwYoc8BfDp
W24rQS3hSqVk8SEvDwjqhp/iAk5Lgsy4eyddVMAi5sJER4lgq8+F1T7coKu0
XF0gC2Ix1aesUbvS+y4Jvn+pjfVrhq4LDiJ38XkkNmaYEmF84z1KYDOe2Bs2
MzVG5gOd/NmOim+WGWdPlJyEFn6KK+ho/7DoVgrw5nFblasRpo8cfAZgb4Ep
h0EXHCSmY9gClqNGRMvh0lpaO+L2ou+Oueszjp85iPYfALQevNuPwZ5wa2rv
W/oE9nWjpt3mA1xLHNCayflfBFKvVirLTXY3ZPzCLjR3+ldOJKeNVh3KrWMv
NMMXNiaLbwF+BQoQH4Sp7m0S2ayzecyVARe5B0D6GqAi949XJcMk0I7vX2/G
4MafaGJUZH/2DUpqaWXSRB9B3NHoaeJuHD2NT0mb506u5djoEQtP+9vPDK+5
6ykq5/dWxN4XN0v4OdYdh5LA3FtX94UIsImByhrkA1/XcOx9bsSgX3VeZsdN
xYlaRewSsix7Bc+z0e29ZGp+/YY4TvQjrAo5Z03Vwk3TLk8fVnVVVIY6wOVb
ReOSMMPwDBF2YBpGgsA4+gH7h9VRyk6FbGZixYG0zcLS8gSJsPuYP8ofDzgq
gL+xgsy3VVOnd3upth2Q/6lWhHMIQQkQXhO/bYDTJOX2zMgu+GI0HSr81Arz
ngiTXJVV9UMsNBA/lVfODCT7fPU6IzwP78HFysMMSgKjBC6S0h30GtZMgm/Q
ygmiZWDYjxXBJjRHB5UKf3t+7MdqZ2vfKnedNmI7hmokradUtWsxQMzYROD2
DHo9hmfAJdn2epaAk6LUnx6QOqFDxJwzxIIt+lmrYRFWeLCGRj0tGdfc6h0a
EnMsLzqPyrdciqqX+ssgL9F4mwdo65GzNTKFJr9NIsggjfqEg1lH5H140Xuo
L+FeHRqQnM0pcQ/pGVi4mvZ8/PJL7EBU5hU3uf7sg6u/FNcRQZQI2y3JGGce
7mMfHIx3kqdkEL9TUVXcropQ9CVkAKBCDKbz5c67FjCwyT2Ox4sfwnNXyrdk
yaZoqT0IdKiuDQsU+F87JZh/pPFad6rgDRsiTABWLnx7uS+K+8SxdQUoeq7h
vSK4bRWDEwWBlcAOnRA6kWJhtEPAl/sBTKanZ3TjzFUpU87gL2HH7GCpXY8W
/zpv0yfqvmVoj6Tw1Ye9Ow/HtPzVKPUtzyagv/dUWaj/1dE38CJqH+3kqI72
a8LoscH1NMUzCX5TFuKueXDYBv83ifEBQtigyZGyRkl8kEQvkZNrJJz+5CkD
BFCDDPEzo906TyzuEFehrP+cYflvz/E12M+7g3WeyW/Px4COo53I1EfZmSeA
kcTEyIfiye62PEcZhYZ3bqltNCrX3f2Ct4asVIBf/OUlXHDN+pRxab+SMEeW
Rg1ZVcXhQeZ92zM/fhwBTiXJPTIfqmliAtvajwPUu5ObmFd5vcJyI+C5w1x0
//McTgUj9nzD5jym3SZ0VQBTuUohH7Z89hpgPwvA8LcssLiWixbj2Tykvezj
BpbMVi/jYTJ86iecDont5n+xVcxFgxPN50RqEJW6QVC1LaRMGi908yJNIkSn
OSZWntNNBPkDEyO+9h+TPhK0fQH8n5rvD+CbliV4wds3pyNGa9nn7EmXWvXR
K/9xY+RraKTym1uU7phC5YCH5vgQgorgG5c2aakp70KK8/r6yHDVH8TMZz1Y
9fuJbXlUbw5KDoqOVE+k92/yDiY+fzDeLiAnHeL7PP3BJNCejBDckDYTqTv0
O1kViWL2DfQuFqlVfQAzXULhhcdZ1dJzXhnj0CiPQmufK5gjgIc4wuh7w2Fj
EwF/+mbAE4xso+5LoW8UgLMVQ+ey9IT8raH8yyytglDQsAOxo7UEmXdqn/bs
J8wL/kYIibT0FvPL7FsUzOZ90+P1+298ZUf19XXsYYFBrWXeuvMp411oyju/
GCT1NsILNg4y2/TAfCtDahxrBXtiMGtpeSwdXgTE0Kyo6OOCSNnOoudXF1cN
W2KrjvnMqGynyXtIQegSss98w3IfK9SC9ghTJPSP5xyCcszsWQEWxxyi4OjD
mNcnfZyG6rMlWEofNpHHbr3S1CKmxB6IraezmNyQZ8VBmuIYU2kx/PsiYpXp
W6pB2Esu7gUlMhVG1eibQ4QR8WjNELlrP3h3CDNjhU/EFE+Jllrryjag0QtR
khq94rrvUv+Q9hFxVA0s/DP/nj5hoB4WODwD9eH1IM10iMKdyH5A2crgKoUC
ljsOjdaNIcjeFVf4HHetrWY6oMu626ln3ZtuFGEnPN8PA6I/e5WNbyi94jo+
wQdW+sFqY98FfhgFy1pwNQevLH6F2BRjIjKaxNO9OH26K2aHkyd69hsAgtVl
Nter79jKhg96PBgN/JLThcemmBhCkua0ScJXPza470PvPb65X18VQ4cmteFp
xtzxEPgOFdBSZDYMNbl6Ur6LTjw+S7HolEp3hlbr/NlRlu6uLa4OdptmAjix
C7akiPyGy2pJskws+Lu+ZKGQXB9r95p2ukkdrTjXrd+7sv1XjN9+IY3Luyvx
BxhK9InL6F3gDDgj1HKXxRgLgXZC+8Liqjz8UslAWimT/eUtIR0LMjse+Ynk
Jid8RgbAgCC++ILV6NzS2aW1qaZvA5wDHcTbD/OJYE297TvVkUUFyXwVM0u7
qzGd2LIWADU0VlDt89QR9QHoT7PgDhcX97Mal84nQfB3Tq49pVNbMfDBvKET
nId7Wt+a6L1i/ViqG6UBn7sx5JSMkzu15t/jLkgTIXx7mQXHNhL2a7Cbixy2
dLsYLU4K8bg10+fQl77nOhP1BiK9DFFOPIYzojLIbxJW8xXlk49RQtk9wMnR
c4glrTDPvm90HpndIMT1u3roiHqSWg+det+QWiihMypcL7hHAT7hJNAy71ek
/wXihVGFfDsNStTgQZ+7k12hy80cDGNoP0azTmCuV4COkgi9GVZnaK5Bslp6
fxnxrE2Jrzri7mv13XB1daI8JsCN9/jX/fCyf/ptelwFN3lHBlZHtRMBkX4e
3ThwNFeGBoXJelvFBNshY0+ajCKBycOroVS+ACSZued/2wK/LSyDaXWeLlSM
GakMXgBI8JQ9ZL5QdYtLGSikTd9f06aed4B/ytIXzdQR29Agx+u9kSh82XMC
2Anw8ikUFsWtmvOdN6GVhdwboVaEtFdCm2hl67+4/yJqXfQNC3mQV1sK9QRg
lE58KKEevIIB/RU2MItXf0H9jYt/ZA9zvwFPbMLnf5/m2xYoyMMpxTrTvQ6D
TRRAW8tbqBcuAQ8aEB9Dur8lwwJsxE7efjO2m9KngBQIltzMN+0CSLovxxTT
GTPY4xSNVyBPGzB4dcByCjIyRbrqAurDzZ/cLIDqetMBmCWZV15IpStEIrip
ABTqVV1Z9ZE2ZHc+Bhs3fMqV866fx6mNejuvRsJWVG//6Q2eHLpyTmPUVwuW
sGz0NtJXc0NarECybGq/PZxFPNeMInA+OAUSNUOvvALtVNt1tn2LZDu4riHY
DGq1GSndwSF85tWiMAKXC1TDjbVeXSEolZn/Ems0oyH5Wsfbg8o2isHHsBEt
oCL+LEa+0+qVK0eGVrfyH8kVBRIzDco4lrs/X0NxhCLUgmwbnY9XQEGABQX2
3HzohKXUzzbOx2SfYiT5U1GTxh27Rr590lJmFo6CQyNIPzXmUaxsWM3ilcFY
bffzKtkr17JQCztb4DzxvwZdJK4u1I40QsAkbAs42jD58x2fobtjfPV/9UNL
QX7pSX3Xs3f0ifu1Dux5WknnwltmbsH2oTyfa3RePZWOlpfqaBWZD3/TcX9K
PABBFhuBfKaQZeiEdT9OKJ5pbaO/2XIqjc7k5iDoTN+6nxlmyjo93zwmhl2L
oEQzgujseibETy8Sp6ygrztpWZL44xVb8gjwICIvsxDkvuifbBAGABEFVyHT
9F1tq7+1Nwzx0XjCCooBMQsK3B8TIJ4p7Kd+aB2DByOyvpijKRHEaajhN+PD
FhAs9igXFxJUua1ef3hu8JxkaxaZvDcb+sF64of7pP9ChFykVuajLD/JMv6d
fwlN72jxPzySYhWw63vZqUccviSKdv1O38beSp379fTVoLcNiH4A52IZnGZX
JdQ1HjaLUu+0Alj+OzA+FftPFlhulQEkCh6sgiynlxOiRPworrJ5tVM31l+J
O6WK9c4IU+6ZD9SzMCV4w0zpJoVLW1qLYFxfGyzEj589yIxEq88TXiYqk4zi
nob1TvgrkvIpUJzhchiai/dK0szN9Y4AMY1ukVIo/6BIqJ4LyESMfaWDlU2O
1EzJS3BNTISYbOt/jkOkfF/gSIii9TgCdkyYu9u7FPOboruQo8j1PWqZEBle
myx2veldhz9fvTCeq0aBztd4Fz96E+YlPXM7wlI5+RmBdN1cJosIKzSvkYdq
qR5OHPQeX9eZeljkhyaYRWGrUwvVUYddQaDowPyqX3I6adpeR9MSLEs/6+qg
9OBvhQX1iHTB+21aCFat6Ao39BgCZ+hoDwmDTnWYw+81CxFq8U/aYdmUq072
YjozPFfKl87/33AjihS8u/Di5J0q/bEzsM6cMvQBopI8O0Pet1UsPXbTt/rh
6cq1l1LPcrnb5D8YoE11moiu14yjaWv1ZHZPCx9VKHpo2UoQwR9E7KWLBY3z
f4PN8BOFmPdaeXf4DKJe5mgJR8/huHjGWJGT9JZBwZ1G9g890/gxU4cjmeTb
4I8N8cX8pn/nBU6Aqk+L6+4zkj5llTu/lUyLYWYGnS5bSt4HTcsxyqcz3kXo
GAlHHdnTpJhGNWA6NzliAld7zltyN8UwtjXoYKilTsC1DpFbORK5O99lHmhQ
njwPPn/oFWfmC8+drHNkc+VQgY2Mi8hdf+v05c2juVLyLL1JVVG4/Oo34Ua5
6MeCOdHkVKgxLGDag+DK8mIQ7aqZDzHTi7leLqb+rBwBfwK+iHuddgjbyya4
NGcdR2lnidMAM6tjVMT6+Wql/TtpYszVA87nrvlyTd7ggfNCUF0DR7q0JcTM
deiI59yQ40mspTwoWMfKVvtinDII/xuKKGAEYz5RulmOB3KJbulEehVnwW8e
0HO9v3sUY9izkvtXzsR60W1OYnH9hFtkJiRVBum710b/UjbScLBE8nGGr6oK
SRlPu1qtYgp5x3YZHNwsqI57SxjJx/LgvdSv6m36OwyvHJ7xxpDDejdleWe3
nErMdNXY9lILJRLQH2V6HIkeZocwpz1AGBm+TS7B4xKIleOGcxeA5Xx5fY1Z
KFG8wezLayIAYlSYi7m/V6DxkeTJpBW+0FdQ+uWMxej+57Lc2kt6NSyQ84WS
r3E/gdOCISFXvjQQvl6dIdOb+gBx9oijcurdKTTHJWYpCaAtnIT16GiADxre
4MM5tbdV98TS1yDlSyXz5q7jmXswAY4i8roOHz8RYvKl6YQ2VScTJHuDYyeu
1G7jvdl3fdAU50mmNQUbkzsJNS9PE41S/hEFdjUscuV6qpABKLrDJS1rV+/x
lrl5OYqeyOP/dWIdyPa0LTAVamaeIpA+/eUpmKvLLEMm1+H/w6hT6SAAnC43
D8r1mF/ent0uXTC2Ky8d5ohXYB5bWNbBRA9imV2kxEKlFm+CIRn5FLRBuVqR
Jm5tCFLjV3BPL5vfrpEfc2XaWvQvblLMIDmTxIS38dq+/KO2Xo7JOl3+QKL/
q8dD/QE3ADoSBIALqHxrpzGYqYoAVuX3XvvOg0uVVHUzsICj+T+8iGBFNO3O
jy2B/fjO7xK3XaKlHAeVFaeZZyNxElcBqraf+PC2JhNFlTyYbDyHLNHoKmBp
23ExZ3JfitKSu3C1bAqgxVGg2HAvW1vQMcfQheodR4K+38pu5X8CX0bXYeDV
0Uxx33kdtAtTp9yeTDwlkWpfBmcuDrVmpsZewsJ7Ep3w2nTrWP1zUtFjoR+5
V95db8s9M/iTZdkUdwk2sq+amLKVMqWR1Ptv854fvvE8uOCQn6ZV1/NsWUon
QnM6EUnhZ4OcOEsAiXorwYp5rLxmG13rr8ZY7wFAJX9mMTnXxuus7NSPDpro
Nd5b7+8YA51T0t7WMZ2azdlfcrUoKTQscC3iRBTGj5Z23oEKIEUasOjgN058
gdyY6KhC5K0d0+LMqgrdKuPO1ycVDrqVcJM6k2m8hMowgHjV5WMRQDSOpKxa
1gvy8PZNeVyll2m3SQdJ9pcOhVB+dxORmcF+1sA2wj8MzagFf/dnf4G1ItBl
SBvCNaeNnFoDNryveETzCSfO7EojUGZh7p+Qi0I611TP143TCCU2uqjdeeuq
dH4NRxmJsRrHOU7GwnCHhXyZdljzGE2sAHJ/0DWVwjKD090k1vLcQVwfKRKV
wIOQAUfo1YaW7hhE0CIlXQLr5lPZHAH0yB6+8ATFbieu6qshAOh5u7dp4WZI
RXoHOKbkbYqedPkqQkvB2T6tgbQe6HonrKr8MlhTkS5dsSLnoQ4NMJX+ul55
9L9h/TcViOgV/WQlBiPiWNQFVFavesbu0sayK2WAr7bW/irhVMydTG41keoh
LOK6EhpaErygMSpgyoNm1z3Ks0zqXzveU1/cUOS9w6AnX14Ntev0EekzjVgr
B1mz2yI7w7yLH159qEd6WZvFvxN/DkEFEDPA9ELQJTfXWxY8X4INFSZTk3v0
CMo6xwr3hiWu4HQhCICj3VA2X+ESF2IWR00WtY+jF6E9kkhDIKGig72fIqBq
x5h4cxeCxhe5Y7pLks2Ez4RanQGWvyhVpJIKSu351dhkOfw7zI9qRQi8bnwb
GNaZPiTJOta0RZ9cQvt/WF5ssqP6vHGwXfTAOPfLvJZHBQN6Gx7Rd8dZhJHk
mnY+cGVmwHPxyNv2xoLgiNc039TjH31y9ZKi21kWjnCbgRx7QM8IYX/lJwNM
gbc4/kpFjDwsK8iDTlZxbjaYx8pxRJOXAqkP6kR/s+4c74OFe7L1xzm4PY0v
HGECyAJwJt9d4A6U55esfBogY/tLxnZn6B8lorQABHj/0Sql+GAW1ph9qIP7
8w0PjqVGpqhcH98/uQZ8N/3kpxQ+BuuFG4ctqc8LaI1bYjdZKyQzKlhxKzmZ
V+sEnfcISrwEqZQ/SGpnYj5RPuSSYCnvhoyFeYYoAOaH1wN6dfSGvUHnuwpO
LX1BJ3jOqXHjCjeRj8EITIC8EWQcC0bKtOZyb438y3PY9tqbc8H5uGgBAN3b
iv73FnqDswktc/4IRqJ5rGx+WQysF31nszxaIoGL1WCiUeWKl7LLYi8gFjht
wqEuAqQa9qEf9VgA3pkSnliBQk2snhyC4PwlIomyOkaZEu7jw5o7XJjJiL65
oCuLwSKOn2LARJeXpg3dGG5BzMVWIJz4M8YonmtmoOhXRcsGO33vLBa4NUid
PcYQQYUw4jN9fp01gCxS2roTSMagGGF9o2DwSTyZ8hMBhWdZ4buvRot00Adc
vndikqCP67BaQj7HyaKkvhdNISelU6KCnE+ukEtcIAbBKTSwSg+NGmOdRNd6
u3+WzFjKpcnRH+1HOAyaPmmwUMgSoZO76+Ij+80/PVOJtrrhoX5Ik5KVkD53
+bKikk24vxDudQ1GPMgZ5cJd/1vbzT6LuL+mGBAS2Dn/5/WiABMALydP3xL2
3GcEUF4iYPNvatsXkCXjetZZEFjxfO+OwiYm/wV6+cEdsyHg/6qNcTF3i3pq
sfUp6NOnA3mw+wSDK8UDzRriJ8N5s1rfSrCpEDRWP3+oQL40woOjkZagZIbW
HkiabU46yq02XFqIzp2PEkJ0ZfCCDCnyCHqROg/QNw4s+HkfT90xLB5NK1Sw
4bHJtnQyqh+rts64lBJAYJmY2umAtFGhH9XYBooMEedBu6xbVcZ/EM6o7wvF
V/0K31ww0tTVtT9xuRdtNFDZxyDKtFh8Gk02MqXrGA9gu1Sh42vkJ6j3z7d/
9LtyXSTjagxtshsYFUyeg0q1ALwd2huLq/aVjYdjvuUwccojNcvsn19mKhFh
Yoqk3pb01rqaCwjr4USLyp1kw8Y8q1gA+RMTo4eLz9T63kAfewYQXoDLjoXB
YqwM/uGjWvEx4qVEtHtF7cKqhamWTkGj+VGHar4NUIMmADDLB/QSbxJWH114
Q4i8hR511zIfvMdxTV4HSwJXKrSUhemLlu8BCNeE63zehKU8LL6gg/zKO2+e
Exs9Y/qr7U7VKKe6JA1W2244vUrzi17bHgtQXhVxn3RT/hPc90l9ouBR1qVY
iojHdfB/vBKqAjHmMH9AaipDb23amrZhP2hwzl+JrGS9A5TqMu+ErzVCxCu9
jNcg0KRiKj0ViFY35YTT4lpJGPFyZUJPdeJOvz7A9RYDbUQHjYgcfSstZtDL
MXcKHG0k2B07KjMw+ABQJB+676V3C7sDeA0OrmsB0vi+ORlDV+vcwSyvOg0M
gAHBa3UsO6WJyZUceIMM6gYqWWhgHAIytYxstTplMAIgkjqU8zYIRBwBx2Lg
xIeqerKjvbiqI0JJxWpJlSVkT/aYrGBm97gwMG/dT8yU/tzEbD/wHJ4BxBes
QWKWQPO6nIJjlHAyJCavVNQTksQa/Jj7VRYzssjPHSR2skaCr7YAFnbVQ64D
QhP+iczkp+aZHSovFQZehFgHCSRz70cBhcVBzmxAWCC+vjmWsPwhVMMIBWlR
mjU5Ac3wkyqyFbA5gGwbq3LQ6bMRslqLpWiV/3+OsG8lupZF7K5qnIesnGkk
UmQdN8TGwtOOG+cQ5NLc8XW+R5gjq4/vweiylr0XsToMR5jK9pHLxgULHP+Y
NJOav99ftkWZAkVsCXPu12sNPNpQfJX+KQtcS5wpK2es7iU7BlsqEYHXTWmh
MxS2UG9n7ZO/bCfDY8TcnKeAgctDNh1bJVA/OGN2YGlpboYt2tl9Vhu92pQG
ebgc5HPKnPZjtMGVxJFWu3px5Q8Jpk39fo9ZfdLL3BKErn2K4N1UBGix1ht/
RS+SM/XaGG+slWX1ydmFFOwK+FnibicYtBOa7kqsruok5a/jLFXrU46YAm5u
dx4w3MRSIcDn5rjIwjt2rqQggEh6S64f5uF3jkIqH6WpShm9AXbjD++YniOM
w1TO9sCaRfEK83wON7wzvhAAeKjYZv4tSu7RTAnZxBmkbUIllDmshMlspvqn
SZHJJxgEW0xjlZFwhUMul0XEtI7y8DyY1E3ami/6KNaaqVlsALc3N3VGrw+j
8tSiuFDHkU6yI8etbVQp6G/zjPvwoXc2aG9yI0owKoYVMQW5L6aiY+8linOR
0KZIDgPqtPQY+1R4TIci8S7VyFQ92mJrIwyS/8sAlaUZmeNVHWdDk+39iP8I
Tf5TeZTLkSninkIYyNcOGhZ/VbsDQimA/u+TAeeq4JWhREnMth02vb5IEToo
HiYO4Twg6pnGzpuFrnS/PGbeczLJALCDRBPTobg4fieSWxaFwNBPII/MMfqA
O/xKAu1RCZQ15+Wgio6GosDBjdxfZTvhTyg4tSx2g/tHVAGwmWBPAH4MbGZN
CdGnFP9kbafZT6y2qX5a8HmHIOZAx94bqhzyHUj8eBTBRoB2UEqNf5cm4mfI
7JeVv0Do97n9DLLiNkJLZuFPi0S1/HwbIwd2ZF0EeiRag4rLPPEBzxmbMaGs
O4UchmhQlFCafb8tt5n4hw8iz4muJ7egHB6Zc+jyO70rKNcVX7Hg+tjDyVw7
51t1M2R18iEuW3qDvNlQtZbvtAg6fGYqvb0+1+UCgJyzD7AhPbWI2Et8UxgB
5pxqpMJc70iY9YhMEpKCiP1F78s3omQ2AlhySIBeg+WH3aqrA+B6bpZ8mmuQ
k8ZD5mfow0Dk24TlDxNSN3tKoHne4k4E76zcLMc1i33vuxgjnP5KXGul3N0m
AzzINSAUnUXjdOTGQt1dx1J7+QNOaukk0q5wZScysl1tuiAkfMGHfs/pA4tE
luZ/smpp4L2msH4JkhUy5EvqmjdJ9er0+bdgFUreJhbSLV8U+U5WTtUN/X7l
B/4ImcWCkLq7tikYs+eBr5iVdZTCuaxkHdhmE5uElEHhgczQfuGbyAgFkowN
OUtRwvhnI3OvwEaTUQpiSAjWACmbOludHAg5BV8rPa7S7E1ssZxdD0RFLO1x
3euLYJNiwo3hk6Os5iITAiX6OL5e3MfK+1GhBXMUcDaAdby2Gjn/79X2q0o7
imehQJ8X/7m5BG9lG+65f7ihQmJTdBz37arVzbKeY0T5JmMYD/TBlOtUsT9P
IiEuQ/O7yNdBcT8lvjhcsvmy9aRQKlmPhYBL8/M+0oB1pRnx3d2qpjqKLLrs
yj9T5GQH9u0CQ7hGWUoTvDqc6PnO12Tp4FWqaFVcGFv79rek9JrEuUKH1VKY
xVUfBj3A6xmF41z1gcQaGaxlX8Tq17yjcCRjfiVsFt6bK/wsRY2Z9H97dPBt
E+kzwu/ECQvCpEj0+gXJofliSyvSX5CquRTkmOHIhWAiKQHuRY6jQdEPIUU1
54z+zteJgUgwFOXqJUGV3QgT7MDiByzpnf5paq5gQ1G/1K70EmwCpJYAf7yX
B7OM4AXp4PP4TeK/Nfr9ecUJ/U/MZnBI/B2MhyiormQzWTcs0P9dMoyjOrut
UBdqsZo2BYNhe0xwu5DjWUkfTLlalfb6wC6zIgWsy6Gx0bP2J2yQq3y2z824
xDLxJFzkV6K4olP3PsB9mq4RAgpCqIo0NMgFmCwNOlUG8Jso1bZMNPq3w3Fc
EgIhpkp0boWGWprwxgV9Pi+KfqTo2mCgpaLhaLR7vfbEk4UZTRJdC4XvA7qT
4gmjdEdjmlsPLqRvopBS18ZaAjMe+fiGbcK/wXPgMmQvFjBmkT+DOckcVRBH
dRZPNwhGSmhA5EgkPlwGlDX/jHgXKyr0kpo3xoZYa6rc7NkeNupbUQTci9Dy
L5MYCTulhQ1ly+xZeJNolIRTdMhGVPD/QrBoRUDKEZjstueEeEDgqf+FAOpC
WHUBc4UrKUeN0ll8v1twvvFS3USM2jDuP0YGcHAyhaTTx0DX0V3fRopsmokB
klP2p9wesrg6oChwyTxK3uFR29HCCGZ36CZGFYOaXdR9KHjJoGj42TM/EYVd
vSvEWIGwxPImhqtXrfgjfZ5EYj+HXpv/nKS+zFU67sKup5r9AibCgPlGVty5
PF6zb8WdZKgo5sTDqe8KYRcwFVOm2Osh4DsVxGi1/nAUsF+mnjHCKxL76Zo+
XiZ45sqU2IXEyKuniu4WVwSVUSExKh1BL6ycSwnK0tsn4ycnCsQNbYAc+dRV
SWv8XcldJEopWM/ftStKtpr8eswpYrv7eAmS/Jh+c1DpWPJiuv66vJvcPeCp
k+XaLWCI6264wTYql8fQwXTPVPMqmrH3DKuHCHTAe0pDakpRxZXFzTbqRkdm
8XKqOSgnB2HeRGIysWr7K9Klw+jBVFZhASHUD5yWvStj53Th++7hO5wU7wG0
Kuo2N0/oLGeEQrbdIPqiEYwQsnQ5wRpnY/w8+TplZFPH/Ltk0QGOq0yobeH8
4dMglQgCYpYeNHXGYR2V37aSHB8l7CjSx7UCl8QODD/VUTXqzo+O1sNedKGy
vRZ9XseMSNRt0Y1a66BRIqvtf9BP/l8XP5MsGqRkOCX5Bfmi1dFdf70BLyiJ
V8zLwOswKwkm7+aOex3KG/qwB4lUmbNs+gc4cZeP1/IyyPiLLwka2UwvY+tC
XqRT76dNEwQmTI7YjEh5TWTQ8tEViUyTC+T5UCflX1mt0ZQ+NF9UPjrtHPrj
WFDXMVQhnBndyhetagZEwNguFQmCYUQT/hvB1SZyd/Yulq3QjsxRslDstsks
9JhPtG7yDInd5qSIzfRUMyPtA0db//eLv1HknDtXXrYcjCLy6u6Mf4ZC3p54
PpsycZvBNUxhUYCTzwlfbWh456Dh6Pi5VGmn7pFOf6qiBGJFKF7E5S4xNuR9
B7BrCR6i4M35YVm27OB8ksmTNN/B9Dqv1h9aRpHr2OihKquotDVYyeZ+txYU
+l5A7IDYMZXCD5xfcEh4iIBtk1ClvGR5Qij2laYn69YjYXh+gAj2EwTIEZik
6AjwjWYg5AFlyi3/9R1djRpmy2QEdRvGEVRpuxe/I33WjVR2WYjZxRhsbSr9
CeP3MHobXdcN27hGuS82W2T9C892wgQ/nqtxkEpNukRkIgOLg3rIME62U8ws
GO1diS8zT8H1C425PL7E3d+c0ylY/y33sQoMQBaJdzQwJbwJuMC+eVXi6miE
YujYjrJJzfc4rXItUFAdbDJPEqd3lae8MpyAO972znxxnoz+cYEGKkIybQ24
0rzX1y0jqF1JUSZYHY4Z/bEsVF6b9RRpZ8Gn3cFUMusJWSBIze+pHcVWZwHJ
EIbZAdnHEXxiz866LqhNUH9xP3cnBvR1xFajhAZGEdPcgpSHybHhSGZtC0U1
Yn0TGApCd5ADJPjg83h1itviz8YRwXJzX6cRWDmzeO01JpewTj1ksqWNgL5P
mF78oJZ0qYnGJ5EcYD9guPLcz8/RQmhJHiPkgJ+McrYgYvGQ2YoQ1PZgM+e5
xgmBVEzoUeqyWVWvhMhI7gLU6UJc9i1AIkFr88VotALif1QR27rgfeq7AVGV
xNYg12xdne20y1zwOqPCY0zwF2G2EbdcrACdQuBIEshLqL6Si8Tr2mlA/5xQ
mO4FxD30iGPavDHR6XadWLxH9raSSftSjcUk9CedqcoJnmPiHsj3gxNcttac
C7dSg8MQU0bLJPLh3CCVPyiauwThxAGUMUBkdIQMipPAd7k1tWqrlfqko4FH
gzHmhQy41Htfjkai5Pr4CqvwodeML3MFNZd0uoFG8X0N2jdThvOgs2trPcrZ
RgfmqrmyeKKKpcREPOoLTVO+8eQmLYhU5KfCrgIcDF2GySuLQKjBYIjgo1g6
V42iaYM8kNDlEtj4P4VF15yrF2TSEteWjMroD59udEN1hbk5bUafKqVYEx75
oqhnEsYaz81+kcrPL06tDQfybGQrYVCisW/ySviLL5PvxzCfFeCVfHrnk9kW
zBidtIDJ1bUzS7Bd8tYgvkaJkytGN7xobyIx/CfThg/EEHnrQ2UoR1o0/392
+JO6EQLIqOw7OJv6SEvstUAT5uC5RvLtpmQuUZN2kPJe/7ALLQUiMa3cZW7R
30bd/SEFa48eMFPhJIQe2DjI0WQb8/P5XimHPsbHhnFIeKuOC8xc5pFdr6Mr
m8qyDN6nh+FAJJkk8dOpYr+rZXKURfodUxyzdun9+dHJSPD6TvfX2cMg5wxm
EB2qi9wDRqweYHKSbfrznFKZPehxQW8Ta+LYgG57mPMdox8JAxvsedeUCNoZ
z4rnE0QhHlmE5PEftMU6vOQFE1KBbBsnsrRMpCPRh60xmcWhADpjt2SjfFDl
TTM89r61nU+1g5x5zoZy14ZWywxNEdzglEK+5BUQkM3xwGdag7QWTeRlDnsu
o9qlmj83GpuZz9waous4Qdz6ePkKMqkRuOl79ZfaQTbi+vrQntnqq3Rg7ND8
a3gU6aE43AFm8viehKYnDpBB5EFMkzo3CnHVI9jijO7DQwNKQ1yTYgYPiZej
765mEika+jcpjwYTJ8nx+PgAhyoK61DdxepLRCPRKZkPt49PhQ5XMsNz9ptW
zD0wUZiBMqCZmoyR+PrnJVArSox5yfKPYX+b3ChkowZyRdRh3tCRyx/Iyn+t
T7ynQPykE9GTuUPPyVVwVX0XVNkp8Acl4a+jDhWO3ALFuRyMxMRj2LpzdKbc
NXyOoSQe/4Hoq18MlBhPgblmDSSUorTmaHZUkp5WQmoina12bKNmHeQStiYr
pbhNww0Hsb2qIR8oYs8r86dAbaUgEKpMXm1TcC3nZL0f70TSH3/yE7SdgXER
nB7KDgsy7XIfnRcRGhk0qEySqwBiJBunpCsDytFVqxquDuStMCeGARMfckMT
X22nzY5P8bk+6j7CXY7TGL8GCuV5eTtZp6IndOMos7jc0kQnIeOvxrhg/5rQ
jhq/m2Nvdgq0Zo3x7AChnXSqLTtYIK18ESOGKQD4VigfBiQ4VAvskS0zTide
za1qvMO4g4r+OwL87dAVuTm5YyMEWFagVdBTCQeZvXTgDJmuk4KmpFrRw0cv
FDuW20MqJozmV5zdFPNgXKYJCrEpMidVkWf32DvBul7B3W5VpdEAgnI/NSpY
FIuq5tUeX3F7jzE3KktZoh9MAA3PQI3JWoLQbDkt+V7OmFe2MXXrYUaBXVXr
XhHzfOgqED0kAw6VHN67w71vc0jiuecqpBT61j85GN9C15xVlPXBz8CSsevT
Pd7pbCBJfQEcjhZZqucXkO4WVcaxp/WhBJyV9RMgg0AAuDe37vhx9npfDhT1
XwccQdESkyqf6cH9woXMnxIvk5M9JgFugdUP+C8SyZGy3+dPz0FT1vwt/gfP
QRQRoI9JNWK6LOImm7GuYeTlixodYLc6Q2r70/XbeGTRk8vlP9sMh8T2s1HY
8z/wOv9zaI6LGuGLx4ZQqqYm7kNux8bKFI1TqKWm4OIk7bQ7sbuSoPf0jl8J
mTgIyG0/TiIUD48uR9aF4pZEOaZEgWe+08b/HcqnPTSYGrsIUyIo7IK0f1T0
84X/pAdn5jj0ZOaOd2VjvG2ua0/M/jGlzcvISCN3PCB3K8/6bYrB9awvbBjP
DktnHqlthik9qNVCfHy1XAYyJmRq2f6VDuawFYo2uv5hTpAGG7EswwGtNbHu
qRNrcP3j+x3FQ/skOR6kxx0fZM71ZlBJnyI2+J7tL6ace3Pg+YjXzWc5QcOh
f4qDRhdqKAlw+Y9LQ5LpISSg/YjepYfSNXApm0/IM+bxGRkvoy17e1sk0lpT
nwbszv0O9zxNOaflFtiIxSzcVz7NB/NuZgY2A1s9vh9Ga6yJuX96zVeLLTJW
NxMVZWEwa6r6jc4UtwVfSDdMgK8fwOX54e1VQegOyNNU4WNL6Qs2AA8ykWGF
H9wniC90pNeSsFGRtbna/qIE9wVP6s3GLczsr8HgT+EsGQ2ihculJe0+fk9j
ClpUZDiMQt+XTAMoRz/jrsb403J2gGUZUuqQXMpz/ZE5nbl7LxR1HhX22sX2
JaLQGmltX8GlAp1N31LEp0yXRPNgZ2EecB4RtGGM8YI7dhBcEB3S3ieFgtBd
cuS46zAy7J5KfV0VtOT+soUWUmr8+EiTGZSUqSmZwX1WRcYkaf0FemXRtMTw
dQaxZQWAKI1viq0fv6MXJloYrj/iXwEcveVUYBzQvi+Fz61nLF8AJ36Dq9FD
6Z0Cb4LkBosqE8MP0CHoK9x9e2/RT+hb2khLD/E+Wncv/xQSdElYULUCrIgE
qdbdsvHdfh/Ca8hSiYZtHFleb8JgseHGVLR5XwmtJheOog7cSTLYiP0TUrxh
DK0gVEBoJ48TtUFTF3JEVyH3kFB4vyTkirgFSqWVWHgkXf5DGT2i4ZKIpTet
3exELSS4EQWHWHSDlkUIAyUYsXAsWU7MEK3k5oMHKwVhzyMmTVAMMBWk1cmU
Exewgje2L43m65Fqe+9lHDwUAta3lO5sTrp/cvqqe9kQpaR5q9dlhRGOo8Be
jjJj8VVysppSS7sfnkc4itUW/hvAPu8eGItFrEgDXLsjDaxGoMk7Yzvg1E7R
BftacECyReznh6G83qeOCj71LL89hWfzNCjIccufmRgg/37w5fefJ06iOQeI
1WD9a56GExGZnsH4xJ3Ei5NR7yAbrBHrrTSsUvTVKk6ktBWSzlk2opHMgLLf
QgMTb8J0FPt1rDNF9JDaupRXEBOTWCgF5FBo5/uia4yHRPaqax8ho1+4DUsO
1uN8ooI4TEeQiz8UTDVbpE2NvUv7huC8Bw5YonU1XTl1CLvbQtYQE/1PgqkC
7TlCGf1A+P6FVV87ccCMYGzF1FqYfy2fYZ0LZZcp5Ii0igJrgKBm7jK+ezv9
Lg8DxACa1W0RATJJ9U77XONUUTda/SXaaFkXkeqljkb+FMISsCBtiWRsvKg6
PMDrotpBbA8+Zqn5IvT07OtWX3JMUueCgy/0EhqRI+4Rb3BuiuYGwvMTZRlh
R7rjdGQYakjYnbgKFmOIxuayXQZT7HkTubCN9h51NhYEiIFGNI9TR72Qe//i
URVgSZOg4LJkW1i8W1AfItqXGcy9rhTKR3ouQIg5ZlM6Z9hm+sBTYYtP0wsO
hsr1IpBY5xqIrNzK+AjNHtpWGiACzUJ9RfVBCXyeXKL+CnMn6mjEiJ3o3crB
ea7SACSu7zc2A+ojgrbRS+35ZxdkGxZ6borFAH1oQ0YIsrWXgBdcyZWkYqpR
nGAPXMxhinO6Dliz+k6DjIV2HorSzSbbKuPKtptLxHlH9ersRfk8lpHJKYhx
SEQVEuHTuDKRtfuHyXoqrBj6ybvYx+fCX+2+X8BGAuyJtJhxSI/ZDvF9a9Cd
tPD2j7e4Qu0Dy5qp1L+dQq4sbCEG82P/oQ4XVp9aWxlW9wd5CIx3fEf1K/vk
BtVzX/1nQ4ecllIJdVfk8xnb/Z/SURZrFTf8yGKjQzqUW+hEdoRg+VelYCe6
Y0qMci3EDF5xawz5JJqtuIEJ0hP3MeGELXup9GxzhU7BeXt8u4JVQcee9cvk
EuerDdz5uBDOMZSBekgGfr5W6EE2Ykj/vdDnDiFXEa/Lddi/Nr1LnQTt+Bzy
Ks2s75u1HW8yJjEQ5rP7aowRl8JOG2Tw9e5BNC5cecuBM4iwOB5xvkD4A/O2
oG+XnAE18xBD1lGrLzoIGxqECcHRanQ+kyiiTDdIKBfxEmMchkkAYlEzIDT3
y3hFjeHihUsGrkZDIHIHSVIvUsmCucTPPPn3uA1dXBZO1MhmO1XWuEFzmLPy
YzCMWKIE6n9BGcoTIkF4pQcZNYlPA0BBrrkqlBtgysxMyU5wKGDTJJyLWtpy
yH1pzPPlipwGMJyOuyooHkNHxy4L4gJb9jdz85kLSYSNGL/i4XOM4f3bLRAJ
M3EhXKy7bqx5WTkScQsD/ubcuB7zvgHaNCfEiN4KlDZyfQXIwjcYJ6ljB8q2
4wyNzbs4TU4ouHRPCelXur79/EkXK0YKkWYR2wPieSzFccMuJDU41USJmvQ3
42FC8CmNnkYwGDhVfYT0EPDoY6RcwEvth3oc+rtZdkL7DUYe3XuBFxTuduLA
1+oQItvr5R92XTQElSos3GOwZV4JyBQY5wlzBZLlwKmy70R3V/op+O+ZzubJ
ZcD1X7QxDGJ8Id3/TjjhGoaNUtklTQVsiewYP8inUl/Ujygedarvq/zCbiSn
/VLBG3oK7iExoNQCfMkDy4t5ynkVVZ9+HKF2sPcTjamsiYn9N5L8r/T763ed
PhvSDovcL5tHalqIYSaibke1M0CgpgEJEemrJ3IKov60Wr03Bjf0psc/FZqS
JbabFjHuwDRCEt9+vzpfq4tUwaNLHyZDapTYbcXnDzO5ftGCM7tUdTwKlNNo
1Fev31bD/aARaTNCCY28MAgtQFdL30/+36jgGiEu73dZjns4n2XMVAUYOv8K
V3BmTiuAIhZePFW8RUyzGtUcjZrQoNO5FqurS3VhyoDR0yt74te6CAtn49zm
tSi1jzirTvhlwqg1yuYv5A2zjEhKr4Uq7UZnmXrokSvzc4P3VMMsZFQlce0m
M5VVvWoY4m2XboZkoWgAmCYzoo50jpeHHEXiH4efGzlz5HKfKBSuazC2ITkc
sxxE7oFsFQ8801vU/dkHdItYWbTJjodKfUywifpTj8WXcjvJ+H1ltPgC9PkO
Gb6J7TjM3tdaoJTXCkUA1qR2U1ZLNGP3fY+gq9NA5QaKgcs9Lahlodsu4e/e
4KkLx30RN4bHuNrrDdEc3lQOxvg0R2dEFlyQFJx5WtHKvVOyRpmIsSEE4mfL
Bb4LxlYerSf/H3XA9MO64/B17G/qfkBHzVxrZkqATrM59zWYv7fcfkIXxNT+
fe7iPcsvlbs2GLYe1Td1zW5TEM0aCr0OqbwHq3PqbRuy0+g8dY45icVNZ0eF
FTrrcdnIB6AOa3bfff3ZgKXmhcRraQXbHNl/7v5yT1KJRyprRjZEkGAC1wXP
mBWH1ukubrSCeiJWW60cnPX25KIcNzdZwe5RsLhUKXdUORGSnV2Zay9ioqN/
AyZKhe6lxbubg2vuFT1Gc4vqbjW365LCcv8CtjJkMCY7k3cwpKhibTMiKlMS
MmTnGVsNaLC9KgG/DaP5oXU8EJbo8AWlV6pbdUP1+atQqiA/wQ4vlf6CPPEO
iKnT3c0dqZ2vNZ50J3QtZiCo7is7S50Rq7rxE61YK5JCVhRGHvZxWuTGdcBE
nEVzDTBqC0NnIxOj6Vittfy/zNNdcCvzH4bMPg6Ga4gIMCEy7z+ikXZMG9EX
dXm6tBKAotz1VXkuPyczDHjUiwIxiurE7iZYyPaz0j60JB4KsuZaRf7Rne8/
rzhxznERxCKjpBrdAFSndQcRwo70wRpSFKwvnGYRoMTj4jJfc3YZPjmAcLJC
m6KXI0AtYBwcUjG9ncDHU4evfSR77WZzQtAz7RhbsZsSprCt96+lKLCkZ0Uq
lfcLL3wX/9rro62UDZtMnCp1hSnaPacSM1cwOUaF5Hxkbic2+RsXKK0HWjhZ
Yy+nOL46kpKSQjWB+1vFjlOgztQhsqVfis1dgkY/SVdRdCADF7dtCD/xYwt/
WimPW2jgJkKjjkOn2A9SdU9QN5pN4iY3BUI7f57LlrGi/fPBKb8ICTZj57Gm
2cRc3UbkTXkGDYE59M9PpuO/w2lce6eOA4YF+4x5yBK9f6/BD9ydcmhFeyn5
dIA+0py7yJZEcNazbYwn9r34CpyQMzCYQPRgxD3OqrsssPE/6pai69EhI5nv
Hck/HS2XR8XM9NyHOvfKdMGQ2vJP++6Rz/U4+c84zJG9DbxwsLFEarWFGRt9
Mqd/QsflqfhJ7T5fN0fYBv5e7583j5Kewja2e0Daa2EmmY0bnZgPWEDUKsFF
PEKLmZ5gKhr0bDA/bxpdwwDAu44D/rOYfYNkSim4AMnKWOp0DXtfsFtKygTf
68UcEVImQdQDBxrVuNqfpXhWQKRr1rjunT+yNCnSdN/UiU74XaJ1ULNER+oO
KaINcrjLce7Xodhzkr6uEKZp1ch0lruxn6uIDYnq2SPuT3FK+LGQ/xcYIwb6
ITTyz3CICJBgER3WGfxjDzokwZKFNHDT1g02Usjob+yxLilAiE9aB5hVGioG
0Grn5TZD4koXQ5XA6iKRZr3KxErSUBUY+SIBBjAPPWY5tmLzjLJ0QDkYYgde
NZBO9gljrGlAKZG5Gh8nD424vslSrqHKX3nkIOpwe57UpBlsMqDJWxGAAwzx
vHT6sge/N8jAevbogtdN4WtHIdnUfKcFNE6R/Tls4uuuS9KZWmbO2fhHLEog
MmgmcJ8rUlqpG427KGBg7qonCyN3OKrtVm02neQBkGNG45heev0WPT0E3RPX
GyoAMKpxsr03+Ov4zTrWAfRCWGTNbm762XQpSL+60I+GxCBCl9D1rNA3mu5k
lC11vTu8j8Q+y/2U3KelQKOf5U0hYzuIgrSdLA5of1AvLmbUMc/5euJcum2W
Li1Dm1bsBv7g5qkh0xPC085Lb4IvDLyfY+1WbvzYg1q7GBNQQDYGH2NWepTI
+MoinDU1ePAeR6/fNCM7Z9ueuYbGViWGBkVuHmab3AeWp4fuVH4ro592w8sd
3qSz/ivwP3KeRXeT5DqfOIALU/pl5wfYGhv/fqi+h/D9pONRHzv5LOojXFdT
JVbzX7relDfpL7987tuV9WupWfZS4dVe/TlLJXA1w/BiTOkKAbVjOOCALpwJ
gYEKmkF2+Fljkk+wW4biGl7SPGJ55iF2d0Lw92QgJmrpU7KviDJ8BLqx6ALT
ni7DEuP7Xogjjy0nYVsOpbZtSvVeTKymT6Pzrg5utRI8/E76FoO1oZ5r5Z2J
xEmfrCTCWOuLHtDQucrerlV1PWT/VZGf0AKuoZ+YKVKvreaBpyzO3mPMbw+P
bbxIbc3ZHdkEziLM0YcaOA5V6q524tfpKMhGW9baTOsVC0wGKF8B3sH/A9JQ
JR/VK6BoFAlkS9QK7gt2e/4+LgHywGTmu2b/uqtN/+1QEuGAHioBM/hxyphq
qCSx3wV8ek7mAYNyViOtSOM6eLa8ufm/sQ4l0bIl99n+YCmfkbDTbKg2Dq+z
0YAPH9bReIwoGcyH3sjl3mFGvad+HQishvD2Ab3FCmRXujZ6ndEE6pE/xDvB
ZVoGkiF5go79ucG5J5Bs0Qct8vQl1SGOXR9cnpkpHxUwSeLzGprfNtyWTce5
1TqWjD8zjpYaKhGp2heJrwbKrx6WfQZmZ3izlFvlZf55SKua44pWs0rmr8UA
/MGsmwOPAKwqxKwzR76sd6cflBGnaJKTUeZxW9w6OeQ2LqoDbrSTCpwJCy0m
v3EHG8p7mvFSFPxAz3/Zcf0b3umXbxVGkz8k08nb8HQdb17518bvbu+XW98k
xKgVoiMTS3l/TxcVyYYVSu33L+QguYOgirBzJtndtjaz25UfXNV/ogOtMw1W
5a2ywOZPi11gUD+aPDRdqTbIY055sz9qtQORFRSLUyUdfdjML6Q/8gQw64/9
oz0+e5I1W6x3Mm/AoglctElKWsgQKvbBhp8w2br5B33yWUrfpcdvGShSl361
kuDymYpJnfh7ooJQS0EHpRvqxRwqPqY/4iRjq5XjkF5xFmQa7sTvqII6K9u+
24GL7tP+rW0lsXC3D2qdvZdybAd/ynIIr2ANqvlU2qUIt+he1S8VvTGHk8pe
DCkIxTQHwdRi+VNCbn7qv9TPJThoBypCLreSQT8uxADe8F9vTmYOG/RAYwFy
yRXhKTZvCees/T0bRivgVAPauXQeJTJAhSIJ7OIGGJIOFYWG0MQegAM1RCCJ
gtOJ/VpwFz+b5U0zy1gYDVQqEXKevUkCpXiswxAWkgiwKuO6fP0YC/M5j6XM
62x0EMqPxEy96mjcuWucVzVs2oAgPzC+HAOXRM7XiHo9lwUaJFwqvu7Ohsy8
D5peo8x4umX12vlZkYnd/VLKy6CxCifu83xuJGqupiKaujqE8fQnY7/eBSjU
IPgyqGPHIEUjZ9Yr45/P0Uc8KqonLmxpVJYIMSzM2dESeo2OMsRixozGwlog
EBv57TvJUv2m7N52gnXxTCtqyLSimmgKbLysy/bcwpoHDoNHa+waTaTs4K2k
HlHRSo+ZZdSo9hjeIC4KM80x4EHrpXj90JKqeH2C2tzCBM21eyQ5H9BFNOeK
pEqXa6c1CCN9WYm40LwLU747+pLg/J9U0W0j/ciOU8FoeeL1qdWp1cS8qIqJ
P5nsEAd3WrTTDRvpALZXjLAeX5MP+yWoVbbdxFAZl0dIS108NkQ+7eASDVsX
uZRltwKqm10mWqipEaJf49lNftkSlDCyHj600ADmogAc4D2H2SMhb8Cp8T9F
6ac4Q58C1K2SvwaLKvZqq4DKCoJRhpR/kEuXSMmAy6gYNbA7yYmgyrPe0QrW
4C0WL5yqHlCPOZhPqOpXJqvdQCqOsqD/1WevbjroMqhq0I/6ZPHL23TevN+1
1L+qDvGSJLqiTSNgFlBTAHIS0kaC8uAaF1ZkzcaKllIQOXjxazAey0CtM5BU
OyGdUfshnTbr1WxK/i2dKF5wsbRilk3eq6V4qb/uRc7CCKngIDOmU6ZBNhhz
doXjCE+sCNvbkDH3XNV6MQn83ZImefl6obpSH3q8ogbJj0SK7K1udGThvN0x
4X2uGO5OHZC/YUuZuG3QcIaHuc5DRRnB90Qsf2t38IPvox4Ih51ubizbcqwT
RaUONgUPFXgsekTCepiwG/rUrrR1TeTL5wiMNxU7Tvaje6zElkYTDuliVPsn
fvmdX/20gJ+i6mHNbd2yXEr4E6G/YFS4t4SjylPnxofCTsOGZOR5/voi5dfA
PBjYLmbcg6LkN5/6C3BrWqhe6Jlp/XTj85QtRT2XYY/NZ1RZoUQ8L92aawIB
HAeqLP7CdfqFFfUH9KoTXhT1r8NWp/qxKeyjLivH1px9BjE8rRTxCHOufSBv
mMdfWW/eJw6AqScbvI/G/YPXr1xZKu1GMwPWcrZczsUFWCNsYCWCidVhyoZF
xdmax3LjfFykmDuqA1jMDxhbvqiJpSSKFFSJ+2Csi7PhEqU1LIVPhD7ZtsFN
KVrCmSb+iWIVKaPmbxuJXO93T4eDJ8TdDXj0m6aPrvwQf9zSXYrGycweNd3w
p2CcMHyG05h+bX1/uB13yK2vPCO5gBy0OpxDkXrj62sU5uxrLOUEQEt8/qzG
3qksrhqnfaD7QFibTYgFPNwIPSLFNo0wN+YFyysAa2wKieq8lmPWx5OEv4ah
EpJ3Knv+kdYTATGvEbTd4LRLC3l/yvN/XkVMLZUYWeSdp0FbEKwrEyBS+bXC
0hyUS6jyOy1wYbE+DSUKJgwuw0TKHMnWkLnLSZl+uoEjwSfDlRn5WINtP407
HaMi6l3eZmwvB85E/gh5MRFfnbg5/5yRGID49PY5DMw+9I/Ah8een/jtVvGG
QTxCuK5+vGNTD69jtNZMDXQzVmmQji+gOiHOCXQ8QfmF4G2YlHm1Jenub7Xl
omyDVXEZLRpdio2rVqBIpma+cIfjr/DdgDh86a0ECSsCFwmu4z4in7slGDqZ
ONHgh2Vv5vUTuai6Np1xMVGOJ0t/RZ55DfyX9vklGAf/YcaYzywSGVRdAQy1
LuoSWOCGMMy88ZAJSE6QL3PrV8dwZrHosxQ6x/eGo8recgTU9X3UXoxpXRNg
5GhblR6K4FmaXBMyIxeRUzOEWY548I09ehRbfDjTZLTVIn/OCQf+FpMsAWub
6pjZdjfTyRGTrq1jJPAPlxg6CBC/BJTcQH0UWYXejGemdmzrI9x4z/31FcZm
ALwZqYkaUqwZFL7rWpg8YBL6l09Eaei10Cap9X4f6EkbV6Gtts1K5B2lWjLT
yXiR0QzLBEXcUtwiyTsL3vYcH74eDpvMPYKAafcWFVkvJLBBWcbfQkEskrLf
Rx8g4YNadVfnxhL11w1VDBfv3bDZgRcp8lgvSFOYq5hQbczxiJeL8S6Q6Knd
Ys4AXAt1S/dKgu6sVsEkrPfpklK2KXUk16BKYP43NkaGb/m3jQ1twPEkC8AF
NGuyqdKwNh3/6KIrb9lReuqlpnGBWCYy19cKYGK6tYfmB6E3mlWfeQWIC0zi
+zRds3up+KYqMLQFAZY4uR3E72yjbHvKvZqEOdGxKrYPAedYdvGbyn9mafe6
39PP6JbaqyOZ9JR6uK53O43ScY663ELMmz6+o5mXT5CP9sKRy5XsGy0qij3w
ALKSi83JXVMZe/O0kJKC3+tHNZNnHtbmAeP995PJ+/cl5fLaaBydhxGfdv+L
oj0I/OqNPwn7U1po/IViOICL0h7UiZEwNonvq7fQWzZ2y5Pr7+XhKOyFRJwd
NZ8Sum4M9yPoElSEyJVFROngOyQGbFUqNN43EIzVY+lE8Ha8YRv54Tu9lH0v
FNDDE3tAcXy08DT4baWDFYuyQgZao5j/GtxutbopskMXZB8XMzJeZxEpjR0/
5PuB07filSowN1XxHyM/Q5TQk5YvdCYuTmHpuuJgTSuxmmkbfZVY8g8bDHXK
nLcY5Z/r/UnQ4f/K2yo0GdlSyzJf7jBLId5NU/2R4lWFLWtgFyAqhVKdL65z
JBi6LPWJG2uiwmCOooF3RgrcsMFnCXTtgeGL6BlHwNe9DIUyNSGVCgw5H8GN
TKs8hwGKTTtRsj7iLJG1V/m+IXX0++wcGJrK22cmUYd29FsS08k+fgtMgalb
yWh0SLuebvxyzXBESbN3mAj0PkhzE1Hqo3XN/mjuSmoDMwkkE1Mu8yZMk2NC
lnL6rngCYMa7pMTxROnXXnxZ9VQYQLZsvOvvTaVfmXGdyBoHcJ7mMZvwitMy
FIWjGzUQIMGGL+ZSF2alLXOQyA1lm9wJbh7OMvDnWA3pKmWiq0LLJqtr4mmD
A7Y0r85UynlTmPYuqvZb9k5bPYoEZMXFFKiSBpUsZIBRVksKdrg9xnb9JdGq
zsKOxv6EwJHbKzhxqxo2DvRc+9NRhFPZG7MRMsVUxhWDwU8p1J9m9yvtEP/z
33eYccDrK1wycGb7/HFTSJ1Tt+ZVV+tUe/eDBGZ8clfTsaask4T9L4l6hf6g
5GHW3hm02Yfp3pKOZxLzAHdZnfPv+1tt++guJ+Cx/sEmwIiG6kzRC9fgnxlH
aS1NcxNObkvwb7/VHg/l1G9MEg90tzdHe0Tmqw5zGduq/USgGkkCN26ZigXo
yitSuiIVhF+HtSZpwQB0Y3OIKFYVTNwe/PhvMJ/XwoXA7cqyyG2yYsuitev1
lqo5PQ9oYF5S7mMCtH5ZZUHNvBO2l5mLofjodVF/X3racEQ2c9pLzDkS1m/e
pjxsa+qK/dmKuStyvRY72fEg+TBQLV2bbfBbsJucFqPmhKkdEVbNB3q/9mBL
HcV5+HhYxoOoL4Nbx3GH4Y2e8GEKyrc4b7lRZU1g70VamVKrRFgRo7YHT5wM
oo5Ehk1bXvdwqtuDmI0u/EzBcR1zK+5Pgn+NpWqEBQz0qKmlfEMNJ1pAjgVY
3rt1mAs2QtjSHU5Wx+0NrdUctLXqYmOhe0AtszLT1N5TcPZYnh1wtLhpqly6
uXbU+SjpmxYeKhiZBqZ2elZdnvYRPZFGqMPOX2rDybAKg2GoxMp4/ODDXzyB
19hr+W/2ZtuTJFxc+j9yVC0Z++HvDhl5cB3ynfrjBnPnZ4PD5wZD73nZkwrY
b8ZEvHsJmfrMJ8IkNsv6ite6bvP4gYabyZE1L4zYWGT7xdO2HylyxrrOBABu
7YzuBdyTnk7RRohsA/HzXnpEyp3ic2MTdyieYUyxapxYrCs1tyPzcwi5sMT8
QMNsh2aO6TnJWtmNeIGW9OKflrY63v5r07MLTmXmgfXQ1INlhFf2y+HAv0Bu
ysoNcylzOY54hMwA9NYWVFN7Ilea+pInhJj5VlVF9Iy9rcL045Jjm/rTLm55
pzQrUclfyxIyxVU9PSd1wNtDbG8jlDDnAzXhhQL0ykSasTusziMgi+X9PiKa
f5CJrMItR64fCPZyl+YLwnKPqxRhB+KnvClNbNzvAO0IXXMcwyVCfQkuDpao
cKOCK5qxCTGQNBByLvI6lFFKTFc0KbrJW2s5fIMFAwz5VILVkXS33+sIn3Ne
BjsI5mwSieL5Su+VzxYmcUmlQ67/OS3ICIOKVjp10ACAlcBfoPrZsKtI1hoj
lZ3wq74zM4zPU/fdKdn7RZKyTRWPc/CNVQCQG3Z0i/9A2q+5Mm928XxWEKpg
QNp80mLhZGEOVW7pJ4ff2VotSPOPIwKq7gZMrtzcZ2cil/f9Psor6/6FJ1zN
Vw11X1mzJDsgZyDcN9Wsh7HA7aflaxoFULRNrAluRJiThoy1+uLmzryHddlf
/QmKwgSZEbKLHv0RTOBBCEuJjImG7HxmybZ7PB6UMw3otnJwmDwtw0PclH57
WetpsGekr3AhzCcNOxZHtTTlgHH1iQC+wBHzvk1E9VwAZSUVBSw2s2muj1vI
6aGbCg1Q39B2YaAGfKSz9tdJFnrD/yT7yg9jSWsA9bsSp+IXIxSBMXQO4y5r
mpJD7Mjmb1MYzialpDqdfARC3i4yJIQVt6Jq68JoIEZA9B4/PKYXB4peYR7M
aYxZwzC42Rx3TpPQWejr4yAJolcZKzlutzihHLXhupgVoYrzX6GHsRDTRUNI
Lj1C1UKTanelZzhknqRDUnMOp6u5GoZf+hB/gpOk16rL7osAGWytUzTYXs57
nImI65yMzaTPNdVQTpxlTirJ6KIV/2bApYz55AGvv+Glg11JBv3F5JX5fI1a
/KoH3suQDAYTwKD/Br3gYjqUHZFaoEb9844MmwIT2zSPEVVXpLMjeQH7urMR
cVBE8ZmaTgmCfPnhyUsGJnFNcg22jya7jfdFTwIB7FiNtBlXrIKiYUaBarLu
HDy7MA0gtPCMNpsUxbzpQWNLkAyjy2Vi8JQlsqDEr1f4AwDmj2bpyHDCDRI3
JTB+gIVi3GzetXFhvzI5fVXSDjdxCzl/X7wVjUKp1Tw3NxIx9vR8S8GqYnex
uqDbM6fwgiomrUGXEsi/IlgcLaaHRQLNePhsdkVlH6Bzf8A8OcGPEcgRRwnx
W1YBXCEQ7vNakDOUsUfT5Wai49OZGnH8gW9iaJitsuEzdYXqcxjV4pV1s21o
NWTZLO8Zx9rkcUFngMb6AAAQFFul5IO4iqFL3c2Gtumi3681xww555QlCoC0
1l+2aQOaiW15tvfz008XjxT2+71Z+t5uTqELfqATfOOflyGKDiOaaATkqrPP
VzKEYi6XLSWsylTXglr2SWrYUlScBX+gxIw+6EYu+zNoA85Dtk008BS5HpTD
YtPqK6q6z3DDc+nbA3zt84CMpdA7+Pprhp4QwmVSOnayEMpCBCnTxYvawD9r
+3fMR0ZC+lgbYDCTX78rJ7Buk4zKSIzZ4IfYX9KLmAhwBdB+8hmV0TiX88bA
dYoZGoGHtTrvdeUVldW1dBoWuZF4n3v/myUr9aAMAzAJlgZtLXltKmmz8Nvu
BFxrvlgZ7N0KwMxYhoA+47075dkhro7xqIv6aW8d8XjIMmOPBxHgt/1vWTpj
eJHH2KCtqJ+90DoyUdPAyvLluj/YhRMhG3wUV9Nv/clUPFo9X4sSdkpEgg4V
gKUEi4nZg/7kRiLDq2fr/egYvCx9e835snLtVK3s/aaI9PRWtHG0qUeH9DTi
fgPIwKXfnzmEFyyN5KZr9MiOAute3hpiG1EyndZ0MALOEtviyz2g1g+KyVJ9
t5+1b1500SMn5nv9WaTmANC/J8vNdCV7z/BC1SSFgWwKshLeSwAS58k2ZhVl
URxmsfj2P7hwrZRnE4x4sEgTLjoQZUY/B1GfN4em9swBi2hCIxmU6ARTcLkc
tO5eXwnggWgcBOxVTrJDLC493Vqg2H1y6mlxanHNQyC7VQ0wzuxkBBtZrSeD
9mxvcASibwrmrrk4jZAtw/zHkhwnK42WJNIbXXRZj4dnTvqR1KRoWnt5z85n
5cU5oKWcTrN5H+DmOzqRVSTZ8nkkdfZVTWRh2aYbjuaGBHWGjW/sAZJIchHV
dp6NEYhZbOock6VpOqTpALlOEmTK5AcjzX+m7/FGzHue2VcoVQVv9bk3z5FK
IZ/yv/RQZuBUrduqnNX42Nkn/XzBd7+ajfItIrlzHuu9OKSS5j50Wj1Vj/WI
jncoRf+C6qJRLT9mMe93P/SE2S0duP6m7RJhKUw3yco1bUDD/G2Vneq5gYuz
92z89ZW9FuQUNWIa9/5oZN5eOwI0Qw+q8O7/JuIDaX7cDy60AmJ3EeJiSm/S
26BY9sQ8wmvpxidY7JXIa8sAfKyuxsDVhNiSZ81nI9KlH93NVj5N8tabImuH
+WRmyKvIg+U7lWMUDXBtY2STZ13b0jQAZvx3xWm88wgeTf5v7jIGJyyz8Kr1
42FN4c/ENmqv9pb2SAlz8698mXfQMYt3nBLF5zNLduv6mA/LNlvJVEErfed6
WHkBbiOcPMfXSnELe0Y2NxhGux0kA3Sov3tFLQ5Ye6B2QUDpb7XXBerb0cst
vgFMImxvHiPA10w2RqJYo4RhUVYcGHZ/zZoQiwQ5tJwYmWiKWGBYUisW5suo
jciAsOVgTH6ZRFoGDdXRYM2fVlLRQAA4j/rmXF7+sL6T/I9abUHYxg0M9ckN
BEJJOaS83CEpW46wUgIuNfS2OfI2CUiSJb9WNkpC3A1k1q8rxEpuYNQ9AD02
/w38Kbpbtx/9EuLL3c0J7RDdJUVPCxgkfMuUTJeHUmquBq1tQ66B0ZMo/Kie
i0mkiUjbDylAZCi65hwAAUOZaYZ8Zt1gL/feD93RHxAMkI4UA8yANStisO5F
AalMxRHx6yT0CMLyZ4ywUHcu5h4i9H2U3V+6F2TQJbcY/lZ3AJfNMtxajJJR
hXZsP3JQiesMEBjSwJwQT53Xp5XL56Fxuf3asmW4jrBr9WiWqRYgWhYiPbq+
WY4HPJYKFTK4MVIwFm5nWmJ0N4HRLB9ufl6OPDTguvahpjpV/j4tcCRCPKRe
SFE2dU0N+S/WWV6bqQVZNouQFfTY7S+klyE4fkQnbfdWYvghFC7e2Xm5WgIp
6gs/bLMs9evnOCsUYwYxO8dkKqVrgv7LYXPX9vldSyRSkiS/hU0+2EOaLeaz
r3OqeMovP8BIVciTWiQOq6W2/eSHd/hytvS6AOE5iMlmLdYYGYwPL8cI/eO7
nHhANuz4P9z1M/sjnKwv2v1DBS+hIIryoTAIwrWv/Q/rPsn9uyFd+sgaNRyv
660SVhnv40UU551YHtrgKu7zMlcqyQ/y9qDed9ZE09/HNmiyFsjfPm1lOoUU
uzQaa/Av5MBo4X+Td/G9A0mx6iIqcqUbmUewyMhehWuIWOTVOPJu2JwM01d5
n4/QEaDtw2pAMUJs2biybFZcfG2WU4nkX/GH2WokUHVthPCklMATG+V+rZax
Fyz6vtJIrfvVL7B/PmOyN9hN2b6stMIl7qaow7AOTwaqlwq6VvGA/2cFOwg4
Vslpj8KSGkHgyPPB3eeDIdps5cSAHc8mOjMVGDzjWXZAgc4m7BIqo1WLyIxE
rWGCaN4Kz/BslUwXsq+OnjpkXWge9mGl7csbYh460u/PvgBFLjnO/ASQfCZh
yohtlP87nb1Oddonz28go8LI5+369PEtm6moiBiP3uPdPUi2aH5nrIf0lP7K
sVD8ufSbEMv4EoOwOOEGht7sxUAhbAvRgBqRlb/LVAGQ0LYdQBenYJtNwHRP
BXk1FXPagjfhxh1s/T/Dxqr8f6b5m48eVZ/aNbwpLNDlzuU+VlAIVEhT2cwB
tZW6mHwWE+3yOxzeypNETfZDRvLxeQ6Pwb1Rpttk9jaYLZcoY6PS/4wd73Y+
ZVmWHNnjrUgaHVCn0ip2LBMDCW/XI/qOhY4BAcCB9e+AS41x5W5MuePJsZlp
JfsXmnWGrAUMtinXFPkbVUxuxUDWTG8yM8+E8CIyHAswH9pjukgrQruerW8e
nezcvFfljW7meMEctCBhW2SkXxmKM32MFe7dbMAdFEGMI8SiRLC3yMXJ4Wj5
1WznDOK36nZ1LCkVOdRveJobmkdwrj5KCyL93vX3xaxH/UQ40bGeUVOYiqvR
jzuomu/fQMGRTzAoWNVAGpeChD4Jb/wjAhEAPEH7CpjUZENA+SZo7zVlRBbd
IBtg0L3acsX/KbO59v9TAPcdJ/T9EW6H/oiRlu4vJV8Djv9z6rtDNPD/xxqn
g9crwh1PwGtUIqcCFm9Vpjym+ied5jqihgvxH8B5E6mZ6ndHHRxtqrFRsCCe
SqJDWQLetGTw5SVzYln+a7/uGF5uO4UhGjtng//z3L7GtOkLimxKIPBATd88
QdJnFi92rWEea+so0SRnVVeWt6It41ZkMpEyW9LIlhHuCgnVGxofiWxZ7EeN
GChLklQzjg+ci1YQdnO8e4o6VCK/vP0MVWvxVrEWgHGcB/wQj+D9w4uVzpPQ
5PSYiz5HC3l9A2x56eUdS7QD4xbjB8ERctEOl8Lm218M7Y/55bET4iIiQHXj
nHBSZ8HPdumrGeKz2EKMclK8hvpbzdsca2mVaqRyya6xdFU0QAaEl3nowcPV
z7slqkJTEACPD2Sb+GqLAWwUv8jebz6pO5Ipt/AvOA2ZIHq6XCk7ISkIR0bq
8VO91UYGggm78wV18oNgRLAJqLGZV4XczGZwAObsTxvxbAE/PeNTS/HPAu1W
ZDtJhKy6C5wm/YEuZrd2TGASB9AqtD2RTRMunEUesptaQepJc7JWovI8PWeN
20P7+FeK0UqeCCXxLtwqVPmvBoOSPjsuyShatsk4AyM+8JXsGSxO1cLqrweN
BTpQh20dRH3pvjE5iJBvlWBovPbCmzKj9Vafu1j0WEfif5Q5X1P7JqelrviT
bN2atee3bLpsZiPq94mKO36KYerVnu/E/eYlm+HQaS0qCR1RuyeHh42skHKN
TgCOPAmr4myb3UVjpJaxzdN8Oj+kGCf48rHlfYS0EJWPxwipX8XS4+yly/nt
81LbAgoo2DYZY1FUAsMv5+EWeNZH8lFNUJAxElQu5cKBi+ExiNkL0R5KuzyB
f42MT1U+3A8DOCGVP+x+dGjO7LcR//WujrvMp8kOOhAAHcqJVa/nqKAdr82W
FVXLvS+3fT0CnCZw4jhh/0HmIiBq+qa6k/IQBktbzVtMkMcsgQsMKMgQANri
oT0CicdzPj+ljZuP2/KufH+aABIzTtO57tZuOT/j5ZaLF/xxRrKxKQGRGZGD
pVxL3dnV4Hl6GjgGp91I/sEHQwdLuf70OgjkuO0ij08o7lM+IDJ/nLh8Zi2P
EGO7bL8TxU3ujMnkc1GXtWZG0rrARZvRgUsNkhKf6lym0C/lwJttHA9EI8Ry
3hvPabXJzKJWr1WrfMJT673GLKmt2Ot02nLIrziFhy+S2kCOBIIb5t51kf1b
2IbIGn6PHtE8+L+PwwWBBJjvoxugVC0ESWNlgyi66FeMMreC7E7pFljSWkMS
kPAePaAFbT5MNA8WoJRxSWY4YG/awlOl0kDBoF1Q2Me+1YYYxtntnNhI94iU
usjJ58dhzycxZFzdHWMOyZRGwO0DHXX0DjWXerfJMRvBLkTUpUwztZkAREcj
00Kt/bIKH4V8f8xLhvgsvNBNtBENdaDTRcGb/mrqGJMYjIYjQK91zwrykkNL
31LeVtyXMWXSkbUwXqQ3ZxrQtrkjeWM9yAu3wcSPWJinJwbaKTg7eVfgHc89
d5Qui13oDoftn/cArtdHrRmNQBEk3LMQPc5SP62W5dciLQIgVI0HVap+jr9X
u78/WcuSQ/5DZuGtVW4QGws05pJzrslD3tWk3I+gTN4lJRIPDcZ+22GLNrwz
bDQrPkjAYS0JOwZdBeTF9iLUROtqZD4nJ4fM/cQgA2Tgj0DgcSNkPygHQweE
u2JtBOmJhpyLuWDD0r4B0yZvB4WK63Kwgf/vXExPq8qDA95tIhRMSYQxJVtV
77qFz6F0FKF+N8b8+eE3dQA/IuofDclJN1QL9FtXVtwielZ7F7Ewz5zyRxPR
aKSOvbG5WP+XKO09TfAdOREfKEkhdfo4eQijjOQGuLwjR+85ucPKHh7ayLgH
VUyZZ6gnqt7eaQBsQduyLqRWOUZJmrfY2HbWzFiFjGrbNp/DuJv52VLBoG/s
WmMRvUNrWmuCfkS6KJD4IKZvmgzd7YtSteTUfhQ7r4F/OMLrZQqKGPDhFOXG
+q7UARRdmp79MdEVYj8xG/FF99XEyhGMKaBl5gBEDAtWteshMsMvmZSePlJY
bAUx4RBDcVemhBKTmNCut+7/PPggMxGtqe+nHDoB7A5RjdsOu+bTX1XJG9ZF
kkgYCcNJCDsZWSWUHeOZZjIHrmjqYTR0LKVKMhjW9jfo/Yqgyh1GZkUVkC0Q
LEPi7QE7h/ODnQFoZ8lpEug1tyyMkqaMP6LfO3xDLU9m6HWJ3elA7WfSrs71
n+mG7fhEZ/st3iinO8dm5IpFbheXqxjO73ZbsZG1bf/oswqBP6+uJOcRTnGQ
wD5eiqXuBTqiMK8a1DNgQAXxUiaIaC0x2vJtWskwTc+x39tBxhoIUIdPq6t1
D2wV5r9xLGm5XsQP4Zd6SOqfKRUtchPsrmdHtBZ2xTutCddV6H8ANVdJByEr
yIymi5mDFjZUK/pyTH693Upsb+inYjnDjyzZAufxEZZSkBh1jpJMQTZwNgcB
8Cq1E9ncnWIc+aahT2PDoAaO8Z1h6l08Wwf09NcNWTwNxhhKeeiciLpee0Mq
rJE3jukZWy/5RLrctjbYtvyUvSFs8LZs/2M8FTU0gkEY7geIg8i+76C1Us0M
ZJzCB97ralKHcuVXPByJOBW9r7cNbr/krD96ZCNpWMqW+VGhQWk5Eiw7Klos
OvjmvG/HmkGxDhpGUfLJ3DzpHcgVq6+n/WDhwpeiTZ9shc7vO8wCh862MlP4
aS303mfQ86L+4mZ2Kvv/whmtzyWpu/GsNqzFwIUQMnoamt0ESRn5qkKdtUHD
Wc/czurttGMKKvKdVo8mMxZ5QoyaWvDLppu61u89+hERBFw6wFBB7Hjb24A7
59lVkxdNNJcfS2PteWWDYFe9pNECW3vbI+8q+cXtxcgerULnytQMLxH+uD8u
VzMAcKT0g+Vd1DejsZjeUv7ssQNsTn7J8IfUNxNOkG6qWvUSylkUti+MNhDY
re3oSi/2CwTvMzpQ5f6knH9/jLaG/KMcKaeHEQvA14iZY1T6wmWRMwVbdXaK
HMVyT5b2EvocAHqOoRzaiZiPN2+oOjXxTCKvhjbmginvFAiyGmkPcybzsuWj
dKhVltf89OqXHLj064hfCcNAMc4MisoL3AFIGTcPB5TdxEiDz3yKQtMnxyqh
C5mz0wfF1mw/zzs6e0W8IvgUlhHqBy1FFLPifRO5j5LAVMdVVu04E1s6Emdo
TTWiMYVsQIKdiKTOrsaOVatatNcFVpndwQjMb4SotLe+/EhkMgCncGbXkLlJ
45kN0xQZU9qQPQ7ZS/tYgQZCrPOgJErG7h7hSgCveR+5nsxxgP5pyNC6p19T
zpj22ibjSo3Djok0gUV63TOUMKrYn0iAssUnye6SDCuJt2759qIHFS2LqTyR
MoFrfCztpxZCSNrXWpGDDjmNwDfj0fcw/SUkBLzMfOjY0RX2+pWN2r7UAvoE
X0JJf/nKx8yKM/aDu6qhzacxImcehfGu3xGUxZZq83kGsKo6HK/+O6CWSZI2
NQ2unIE730LYSj3n45IgsVEt89pEZ9KqCkZKWdHSjSRUDsOf5TuvLUjlb/GJ
JzNCGSyz0rL/wkmYnulG2t62vkBjFRqMF7t0u7Qgs8j1XMRZK1scucUJANC5
SZWlEl0v+erHfmiXeqI9UdgpHGBgJivj41i7TvWZc4o1HHxfFikfTIhpg9xc
xnME3vRLy5tbIUm452V6gfL6FMT+5iTOoN9SSlXxCVxnG3BI9sumKlmdqTYV
RNVUh+yc+os6N2oCjPTZU9Qz1z1Nhm5joDJgT+23odyhub9e3mf1MKsDIMjQ
PcC3e4rILrvg3iVNqSRzwcDLtqqRr+I3qgXVm0I6BTvtGjWIUNN+JoI17Rkc
9qHnQaUpiWl46+pbSkAEmjCJeglGu8W6U/ddMuz4SxTG2Ra1aX9id+YsCk3t
r0qPUB6ilZWPuo1t9SNGp2CMlIAlR2t4TDIGvp1UuMK32SGhf2tno46T56sA
32mkWYvmvFdwenEY6MB4OJAEsF0j5xlOvUklVt/KKxwQCNSElfwJX+cIt4Yz
zJw2Cmo1Dm9k1bd7XhwwCq1klWUPjaK3UDrt+0B9hsfoSqx8MfV8OA4KJEEy
MPMrEZDbPeQxpHgkBeqbkTeTDyOcjTxJvMYdpiZAFH4kMRhv5FdM9xozwcXB
CdMeWeaslwUW3jP3f+gnGCHVw17n03uJpgOk9uiKkqiKZogglfWR5LcQHstz
dM5GP2BUoEdM/ofzHkNESsO4+uqJAadHWU7M0PW9rZEvgNJRSpFY2WonEQFu
ND9eWz10PLNc+JRlOOiJFFVA9q9kNx6mgiyurVHuiUpdI0gGUvfFujbzt3GT
OWsNgsIvfhyhHPZ1nSdkPgiU8ySx8AlT6/ufoSTDInxfo4PWPkRpQLbDcU9J
oyS+vLUIIIa3ku3ukhcpv2bmBO3A3dQhsE5CKlmfgRWt92LVq+Smu2+V37Hu
G2shVeEVVn6XtLG4ABN7hfnXK28X59/O9JzqKChRLhPlQEh68/qIV+Dq+ZUv
4j8+504cBG+3UFx0yoedyoBlbaO8y3i1v/Y9HMJSjd8xXqmLHBD96CPVt1UU
vJFaqmTIjAjzXoscF+IPwDJHW2gEodBgvA5QkkZ/oDdTa8BXaf/+Uhk4nS8t
1ffgKhjvOCcmdztISh5E9z8lTiPXHQ/y5wWuEPLbeHDR1MZ00rjjo+rIL/O5
//mfCWRox5TeCNIm4145X9Ok6Ysmlt6qDujHp6WmM3MI5Rl5Pl/P3fxmD1Wh
+0TYE1oS1shI4lkRN9lXC705FgXmZllQ64ULshHN2HwPpe6DYLGsoMQbtf5D
NBuWaFo/LiNwtwwnXWX9dipYrvLGFLAVk3DCqeUahZ+wOOIQrBiozXg7KjSM
XtytCaFzWTRRfCAkHKPxTDuQsZ6NKATg63S3OTixmId0pTCSrloaj0l+eHRE
oVMALmLdEeenYgPbWQMBl2EU/6fzJ17Ch9L+m1GQpetDDvw1RPhW3ZCS9YXJ
meDQFAq1FO8xE6kS8MGbjZ/lLTirnrcTPWZGPuyHvQNDaV6F45MKargdPJNG
Ky51PvDs4C5d9goZ0KRsn6U0w8O/WEjC+itTVVnvV1kKvXlX3+6ugePUvwZX
zhlCbr6YTqq9vMyZYa/HzuBoH2qR55hx7Q5M/enUYWRndIiZTR6b2dOhBzYw
VhG694KGRB440aQ3L2OoTUgt7Tw5vaGRyF57oFKLt0XusAshghCjAhRXMJeo
UgdcGojKPKf6p65W0y0O3286XfxnrnQacJwRTAkCDyT5nTror6Xe9kfD7yK7
egv41uTCHsgivN+oG34damBm51Nfko3Exx/PdA2QXvyAfWVPrQq82OKADrSg
DpS4vmI6Nl8Jwz+EXy308hW2niLtItBplpuCYmsNidJ7G1V7sPB+3+b8wEXZ
QPNEougS6JpooPdGV9MaEN9/6ah0erMcGd8JNu3ZFPh7OlVveN6xFQGL4NTL
EQ9w4B3GyyRdDQdpR+jgV5zXIeQ4slRzyVPcZGfeY6mQhPv16nAMHeSu+J/U
wQSOln00ZXd23ZxLF2FqVRERLOHhp3BSLF2VWI/hd8aNSJocB/OoXjEk55+5
sl7ThN+YwKjiJ2uzIYq+KspDulF0Av++Oze7peu006Us0e2DlG4nUP45HgwN
EXqE/sivI+DPbrAP3/400cUChYzCUb6ovtkVwH2nrMLicLBKARXGrIK55Qwq
1n8SZEFlLIfIFYICwGxjIAhLk5dTuztJLa7zWCHQwEBXaAZL0TJsBaJZnB/5
+/pRK04zAQNo0utyY1rTSka3AeWe74pooZMngqAtt3KYkbaafRzVuQYV9kze
4e12MddwUT2VszGgetvGNXbFHRovduhOPGtDA8D2IJv7GmGJyKcDjqKFPTH5
jqNY1G4S2QCaufLykb/yYsdXzRywzajcyMHMJyXGC8C8DUE7hXt8k3/no9r6
+mf+llYxvlHbzbbAMrsPjM8Jhje6w5OPkSKZTIutUxKKjL0WbcFV7ihE2kg2
l5gdH3HhUPlkp146zqn15LV57kyFAj8Ji3Dy/JBLaj/fF1XbDrMrOFdQ7HOG
GQhTB50Hgd/F3H3zEoeMR+bXIroD0bRP7PJW/o7hHQpPUQNAXRyAQEfyxQeF
zP25nfmK3WSXHEhRcrL52L0R5KAvNdYU7QjtWPO/dW3xttqvWdXguHZIUupZ
DmPgTeK6fTh6EM6JSZthJZSepsQr3whLnNCxPeXPQHy7rKxeCNU2D2AHAyra
JA9iOLvTPTIyIslaJYyiXpAAjzZgLXKKpwLaj+jXGr+ArCby5E8RwYlKvIlY
Fq4xoqzEinoeCx05Jahm61GnpezSOlIPPxKCzg7EVdFZv55uprQbKy5Rjvma
G1qLNdhUJlaiqG/f4+cvoAsyLlDK+Db7zqHTD6qRvRSYhNzV36lH0QFuVMmJ
4VNDykN9HgdtgktNCFCBEGU4Pa1/LaCSvCTpQrNTuRgZgXIKINFdMCZ2XxVu
Ar7qmsBYC31/Qa60tSPh89K5aps40Awp7u5x2fAcvaOf8PJiyt0t5Izm2k3q
Kgan+FggnM7IOW3K9fMCmVbRyQZd0bBIrEP7fTrTBPHoV4RphQzeVeLK3lvZ
AecLwBpR2Ps67g+5OHzvuB4htsp8MCiQmQwEgTB5/mdksU/CXS7TI2oiKA8r
FuNlGM7Ks+wWeZnE3ordj7kgpUauutFD2sPWix/KwN2eEptUuYtbjZJ0r8CX
qRWsF5vuGu86+IpZGqVQTTQu9utmBjb0wQM1lAbbmMrempQpqINi8k0ihVlZ
5yAPbM+EV1pVoxf3aJVsZc/1Y1oHOQ9cB1WlHzf69QX9G3lDS7JtBmKVQZU3
s4Y9lt9vwnJbEj4oDvqKLxznwEQu4Xzs+SbmdRGCbYStVr6Prc1vMvWJhKLA
+eguaO4xRwJQd/cV+rf7z8dSrrxBmohnL5kk96SFIeBtmlhKZADwS+YjMEjL
6m3//z2oFEiUnBR20XmxECId+eipazsmmxezaUH8uGgxLkz7vyTnPhPBzLiJ
Y185vbsJGtnizma5sBRi4XZl5SidKe4K3eCITTjf6yyeInEtsj30vNsDxJkh
xdjGsp2UOqr3Yfge0lbyVHwP7Pj6OpTXiFO/153K381WMcv3ZHn2p32m7pHA
8WptTBEJPtCvVBxTVgDAq21xKnlemZzd4v7LFiRocssrBGQfEvozrXc3qnZq
6MVnAu5eBP//sPNbgHHWXmhOumTOinLji8rewe0b0zDkn+tallS8wlT3oGYm
UCYV5Op8s8Y8zt5rDOMh0NMIZj8GBZTECeaJ6U7LLBfkT6CwrRbbiDL6+G/3
2QnPUUAr6PDnUgEGQ2HctWyS8d35Dwt3lFqClB3LeDsfJkIxcIDrAD2a4NPj
+ZL9TBNSZpFsFP1O8Cp2JM98SfHJ5u1jZBTmJ16rFCfm2iaze06ey3Lt8tPd
SNG38w6rJ20trWWKigrR/h/oQYrTyUJ1VQGhslWPsZK5MANVMJTFfvRCn7WQ
mD4wkeKKjuy1f3/OuL7dmKZ1Uqqey4DeBI9pxCXh9pQxi9Mz+KFUq4XfxqVf
aYVLftSu2XHxm1wuCmbIEsP95LR4pb8Qq4gBLbhZDnofk05FpemaYmslH3S9
RaSCE9KK6iNtGaHbILKl8UiJz1i0jt5Oh2H4NEqqzTklnE1lTBFekn4mEZzn
gyMrPRjErUyHAawIM5s1/OX7W7MFkQksSpIuU0u9vY1KcCWHXss1yKHwL5JW
57ZGlUCY19gT99ReALaop/atoksKMtbaVzRkU+yeJ4TDuLRg1gQUYln+X8Wt
39qMyqz7zeG2PX5zNzQh0HuIssC/mWN2Xl+8a4yU/dnZ3oqVwxOnSmAaEVYM
56qJni2gUuWMvynRFXKWG0cpawq5M4+ax7kc8xVjoR0HUMWGkJIuWmShgMxs
xTT4acrvhGNmlNuHdbfbVPr4/g3E184UXU4/7EotBPA329qW+0iXFSgGSuHS
OjTJq8pV/lMHNDAOpzjhbBqG6GOMknIK50wfcsrvMsDCv41vSYpnsd9RUbSu
jPrnk5Ztk2ShLtvptZh+wAku5NdUqTvwvFphm8QW4+Vx8Q0oh4Gd9jzPVj1p
R6zTRI1KPK/5FNDOSW5XqPVJtDi/MFwckvXiudN35CmxMBs0+9OBEYYcnpvc
eBUNyZj1UAk8xgJM0CS4xvicQrTMuw5ssgUZkw4oMjqT4t33/KQnr/xm7XRm
wuwv9gk2oQsViPalETT/HxUjR0sWxIXqW5w9kiji6TQEIGqWH+J3o7QKKWF1
nZdnTvZQ23n6bA3H2rzM788gLiDBabnVCD6k1jw1sMXlRqMs3fKWnWTwzNyF
uTBItjCcB+aJ25yYcs2r+H8492hmqtF3yz+Iq3uEW0lPSY87GlB1WHC0AVjb
yWSTZqxnO50xBnIcyicdb4Vr42diJQ+Z4Qpny/MzDq7j8ENqCSDFYKPqDCez
WER1ffchRbv5bXUU1khmUl2gp+HNftadeSBuaVOP4IG2QlC3AUJfxd2/3/h8
bq+4UqMy3z8APg9xslTpG4pdkhIOwE6nRDGXV1EvZ55bQCyqgMu3CzVtYRKM
3K3P0lADyjbDNoYoEhaR6ZBR17Jk5fXexMCMBddIbqGEGAOmMahhjWs2eQQL
tBaIMtowymZuNQQDTzy2bCmjK8nOne9mHnPggHJ3tmRKfTh7cntQThfm4UwB
ZtzhkwXKwwISt5OEx8wjK1m4l0Ob7rFdkoS/cVOFDvxX4D7tTLoYajsid2wB
sS/tMji2MKE9hpOX+XUznkIhBwVC5oC+AfGqW4B0+/56KJSbFF2WQQpvOG5n
AnygYqGDX3Yj1SDCyVespAqbBYyG+3J+9/IMqjd22oUk7fbH1YGJmI+Y1vys
Vfx2mqPIv1uNmgD1r6qewoD8DX7/jufujQT27Bz6YqX+4vlTGtvBDIxK2mpU
oP/kqC6JuAaWFsqNAmS6i8HLlaUkOf6aWAWKz6/F19/6C9oTO2U7oWMj2w1i
sCuGbZxAqK8yCdY78hCq/deqGgwTjczfOgY+s6JvsdhFEFTTj0/ZTE1/2TkV
zhVDFZ+9KoTq9hEWclFY+XBFZJEHmWvA84rU7nGc5W/h11HM3g0qrpUsWJYr
63SEHeDVJaneQmLq/UpwQNUOmF2zjNmPrtYKRiTPVu0ihCt8c9cpWPktDDMi
WX6cx13pfvwyxmy4SQzP/mk/blpVBT7kvQXl90MNplBF8eNuW+1pEu0E6qSZ
VYY8YVXjdWnywGGE+adJDbkJnne8Yw10AQko1uTVJlO9brC2kdMYjPnMtU/t
RfG8FsthdnUIPg0ib3lV8spHSecdoCdq/UithFnEZwbg1i0sP6Z9Sd94/auJ
7SIeaqKSTLVK6J1Mg/jSOpATE5m1/pURN6SzIw2iUp8o1Ho+yvB5sD2zv1UQ
La4I2cTNOXhSrjpklU6iCxWeNvPavBMPUGuIiq76IAXg8bUwjRsqtHBT0ck0
3yGzU6bfT52pMhEPd5Y2mK82kAM6lh1XgIAu/6299L62+kAwRFOJsghQPJOp
Ysro1zD6v6+fBqq/31dxYeHHQ615htkbKkRl3yXli53Om70Dg632i0gA1GqV
//D2l65hMtcsHGWxEJd+IuVKO+cTl2aPOL4S8mV1CINUcaA+kqGp2Q034cnn
4ytM6IbGMZ0f185Iv7u6j7kRBV0U4zKFU0LNJ1klcrt9kKFFUz/2UMm7DH5h
n88L6wg98wPT+LG/5GjGpaidLgmwXcjFn8sQoKo24tKCqn4kj+ESjPz6BeuB
mo++WYGeG+k/bnN42vwy5Uv5WjZbmZJium4uTF/sBWiVpNmH1Ixcky0Yv+C3
kjd1IMYLsrR2MKKs/RbnCcjMJHeXqKGCdSuO3x7M/HYQ844GnbAkEk63VJk6
e4kLB0PlHG6o2pZ7IJMYgB48TKP8AibbLT5MzH5K7eFK6j66+e67jqVz12gc
Y4Hc/06hfctvOofn+thEK7Q3GL3zmv8uP0nrZgq6rEYVylxXUX0zOiexJd3R
ryI/0R6d7obKxOZhbNRl94HDqYDNqsGfYsW+1hEUcdElsZf2dnDjvf5GeuP7
DVOAFo9GzmF9IAOCTzzhv2qtRSk+BqJNNLktPQqv9KPx5PpXetCIc8nWq1Ss
3GLtIbVDCdYdcx3ZW0JhSZF24LiSc6LfwnrpSPmKzrhujNX+8fXFK2KVcl/y
32WHTrcDL6AtPgbX9i/BZQNxqoN5TvKs+2AVlXKjDw01SBY8dPmH1qhrF1gi
oXEXCTPkyyZB2yxfwvB7+ZXbpXLtpQ0nuNWzXTjDXVb+dQsXgCj0ZwZlJW1Q
P16NqpVKi9qi+1qufVN2OPHYYsX6dzCjoT123r9n1wWQWq95WrODRNadKofN
WMP4QHzLeVdKbULkyO1YDDQEYtZAY45pVQkfHT7nqddJPDB79vKwv7XOoC+S
0t23WhxpfZVF4Cex4gcPekvOxC1BxZtD6+6ExWvm619PghpXmztAnt6S0dJW
g8ROWyB2fi7Hdlc5piabvyvVX5l8dGrpzl0wKb/4PPvRgvBV2siwZINbg4MH
uRPuiUVP/zpHOjc8iHwdZatSzIeS0KZDOxUxmrwP2XeySCZ4cjS/VMrPxT+G
q7z6FEAv3kMpSiYcu7YvWr+3pQ5T7xrv/y9w4H8mgsTe2Uvg3B2dC7II0Hcy
wBzfTL8vi0c0PBRsizCLgadptK+aeNoI/zBpIWeJJp3dVCbkKOV+0xIz29wO
vqCqoB4tYBcGDtiSqBi+3xMiQlGTA9Xy9J5canejEWkx0ofClKubsvS2le98
hocW8Rv2+dIlebUTQNalzHghoQZnP8Gkzht43dEu8JWWw3wODK/8bKJxQXaw
LyO6VVg9/ThPGQoWcBvTi0M6SQMCbL0zwY/4Av1xUojMxE0Ah5gGARg1GKmK
f5dMrg3qvXxVcOecQOjK44Xth5Wp+hLhB7kNby1nmwckTbQ4bCCJRmwM7nse
gMPAx20VIbYsyubMfv45uEJnffh3eNF2xdh4tIIfNuzw4h5qJuQ9cvvJZ8id
UENvmWJt4osaVSzT6CoRGdZZn2OfPdO+xhmkkn7lgMUDs8X/T0Q+UQ5yC5lk
luD10gaNt3PMvsM7zsfMG6v3JsWpxkRmNSSDSyTjJ9AJdNLZwgmEDPX5NT66
27ZMoqTxQIHrYzZe9VjpefFY0cx+BHoPVJT0RKnj7st7vQ2myjPanObTxnFO
ywPlY4hZ36Ly6X8oArkV1ekGT9fAsfC/T2wTM9Rwc8mE+F5eVr1ldvMc3pza
9zftaKZBBDoZ9CAQ4RTK5oj6nGw0hzkEDxp2/1NxD8rCO2LyiEBDU4smIob9
pgLeaF+RNJW6enMPTJztNW8hCDsh1Wpw2AfL7nSZUJr1cK7b0BBS1SfPB2Vi
PwN/exkD0b3K7Wr1UpiGn/2XhdtA5TbFxR2kHC2KPg/x8+jXd9duneecv7mB
HiRKv20qkiTYzHyLxnU7VZ8QgcbjGXtKJXoks1QD4ni5KWxoB9bWn3/RwH02
W2TwaJ/v0r14ghIcme/ZW6ES3Rcu5PXTSN2daMfHXtXhJz3pGcW/MFErMoI9
jDU1dZXDdPdowq7M7MyAY2QDtK+xqspLJIpiIa6sZTnrcWYXq9Mai60y6hsL
BApy77EY+rVnrJV2hFctK6dZ0hvybMHnR++K3LZ1LTZQrGgIWtYBWEAemni6
f2UP8EQxqXg4vofOqgWPfjZ197zPxLiIW9Oj4zSrrIXvNlbm6vRRQ7tEJPNZ
/S1iO3tOwm9HZjAz8SfAX7NjTU4fAScRxN/O+dOFvA6c16KEQ6HGfF0B+ixE
NA1GqlA0bTIslRkktp80bWs1FEIkqv/klDEscvQNfRxktw4D9GkE3k+GAm5C
Qg0NZHrBwNFr0EEwFjDjRkUuEbpO9+21XFfl5/wbBrCZswx8Ds9mOus7oT6L
mI2vtmhP5RxqsqGaLJ7meqPdowwaKjXzQ7oX1zDen3bt0ppCX2DuHkdsLXh9
MJb06IiWV72MQaCyo+NH+cv08LBQMVnzCDDUgroexosd6Ln9ikIvMzoHwspl
j8pWl7zv0PCUa4O+aKjH+XFkDviGoZpUgjoSeZWxPAPbxetC19cDV4msgEzd
g0XkB1Obtuc2VbMXXadIGFf5jpXPAWMWBHuy+wHwFKWlPpRIIrmSraQzfZwC
QfbKdb1TTu54tV/js1t4nj9jQMZU40x9TzVDLoK5vxTiUv2QpXubPYHZj3hA
14m/BdALzD49V3tWns67nEwNuGYRV7p5sgpj4E8nhxcrhly9msDYdIHNsZSc
U7gT8zqFPwn/6en8oSM3zFTOxMo5en7I8Jwwt9MVBEV/EX9VBSe2njJUvgmR
6kecZa26KaOISRPF1RvErRMb/lMcCdHBSnCZfOCBeqKCok7MycZlPQUJUmVj
zHA6EtuZ7zrWxNZZgXlxD0Tf9vZv6NG6xdklNeJVnFsMzyVnfLvxq5ROqb3w
zGSOo6WEAeQS4jefLx/VJ2rT/P079cqHn66amvcpwZ/5jW3c6E1Jx3sM54wa
Hn9BYDzmVlF5u0k9hzf/z7b3S+oJHNiLVsxOri+u5JlsXOy4qOrsJTGRQBCG
8rd8qOiKI+FnIpJ5+JTaSBpxL6dQXhiYptopPbhkAghdv09bzsz0A94ziw7G
Y78E87asDRzu28Y0r61Gb/lOo0/6YNxMqpUt3yiukr0E+uT6PfPLRY1FAsc/
bEoxV5TP6X1yFcAuxWRLaYoXJIeq+BemvYGYoYY5nvzlRVqI8jeX1BvihpJU
f/ChCNH5Z5xtt6FgHRs5hNQ781db1c2l5zdH+iySyrKYTCa1Xx2MmsROzoVz
Ctdyr1YG9WVtQrhJDNhe48v1aqmIOtp97R6nLdzrTQi94Gic8G0rCrYVlBVN
ODIy18b3S78nnUF2dk5BhsHatATly7f41ARxw5aTqkX1GylSAa4rkW+0+a/m
rI+xBnFZ53KgqqZeIrmDVbZ2gx6GNIpgOmfy74YP4uNPH33huVZrxVOAU0x8
Z30c2VoNSqSSXTmrF8BzL8oKLTLjeD+N95EiQUS3DIUhmRzAIjUqly7F81XX
bld0P4YWzLcFJfeN2HK0D3HuJHo89EwOz0iysdcbIK2Or2nP53xjLTV2qM7e
N3RQcZBrXVXDV9z9VOcKXsztXGpgpMuQ7IH/xj1gAAH5MpEoqbUCd5YOjv/E
QVzqfu4UKnoYSH1U8ZmpZZbx9TOCxdU7r3XNwrLWWuoe3ubEJsElhNbLisVX
RPwPhqOGUGYcbRTFCklrET+jkASRbSzXl8Zvsth0g+d3fqNBwGsS+cNmZ4Of
S3XW6rAj27lhRc8r5xaJtFZoi6MssUAKRkScRdZWFLXOi1G29WItZjKOESvK
VZZU+Z0S+lv1O9Hn0az1189AiDEutMaBlcWSs9/iAsWZ52OqW5drVs5YOJzR
Jp8F0RbjhLtYt/Pp0FYMaHjos53TTxS573n2dJ10Nzqz72/EZpfFn0BEtEeW
YojDJ3id7doDMBS8p4qchbv6BRBAmjDHmmq/4VxJ4+M1/QulledOa0i5KbY3
WziXrrmn4gJZ7aX5ru9RpRhvmaP26TC4/JHjX+qp0cjSmV21HBaxif+/fwD/
MaRGRXfOa/m9EIYg9ZG7WgQUrTJK/Bpj7+IAt4BjCcCb6aA35kquQGkZQMQw
rcY0whhgxCb1ZqnIIgh6fGQcyw+LtyuL2Cuepv5CsWigDNo1IVrTOj3XlGGs
+C/2xIbGfvZahFqI+LHbli2/N98FIx3dOi+OQIK81PfmvGtviHa/HY44Ojpm
M1t51F/OMp2DgemVyxjuOB+GYnUEeNz+FFxTydyer1y9LEhew8ulhPBWae/N
cD6NIOjGDHPBQqw+Xz09XZ/xai5lAKoiy25Z22F9YDpCqCIHLI/J3gRaksox
RkDZOSI/0czQDydXyGwX7FGZVEOOEes41W5H/70hYK/RZ59u/Xf1bvKTl4XT
XcgtPS/8UVT3tE/NPgBHI02pBQO6CtdYAaJF8RfrIEi+WtK4bdZEjR15T2Pe
e+RrBgYgS5UdmK/8A8+bNoIXb17hFqBglPTFOJU2P8k1stWgqkNcG6168ru3
IT2RnWMEOVMDGqnuTqT0Ww2Heoahl9ULKmIplVCC4yBU+Jdjko22EzhY5eN1
+5TTFiGObRWdNf0GH5ccK0sfIWd1kRAOi1Wb1Q7sZulzlPAXCvIsErNuSbXZ
fIxQrqAgWiq+nFHZOmJ7FYjzwY71+TBetQTaO2ptNdgvB7WaXoYuW4Syt7ZG
KuddnGkd8TbvbZna4GfpVYxVjEa98wD/nhXkzruajMJfth71axbiZTsSEGq7
ULNCIgWgNNRTytyf5An1kXX+GZk/93g9xUKSrVxh4YWV8WUqfvUG0sM6Pp9O
SN2A+92auooKNZ+hYadvMVPHrNv8fOHhT1o3ANugFp2V4jHPpZ9/HZ2bZXyQ
E3FFGp4cFj1pYiwDiZ7n3aI4lp71uRY+7mbjKGSGMhlMexOn/JWz162wNneh
w50JZhSoADg0W8kbLRrZEPcRDLuWCrRQo07krs6d1ojJlF9Ogdf2f89fyJQg
FzAzSGUFTh/GVhvBnmXoJ0DWn2KPTjoDtjWemePfCyPY87jhLZiaZCsv3QC6
NZjjwVlyPNxXG10JDiVqZxUtu3mdJBW9Bn8qaWh6FJ/rRbEV1IHbSRym5xXR
7hwPFfrVEaX2mW1TrwDO2WYQSO2d/OES+dboJH3UJ2x4SgrRbk0NOFktFdga
os1YnInX4cCHBbPVFnoDi5j5ougbOjyF1rVY7lrzCc+ypD9dXhxIz0PMUG8h
n8QUNogFA4D7c1KkqRLOTwXrUjMCkmbGEPzpd/Q0UY94RGH2JmfZO5v0wFeN
uJohCryZLpHv3uCFr2FPRF1WXCqhLlSaFt2vulaYNBmdEp9nYsCtZ9TyfvfG
KLSzO9t9Fnyb8gxw1atEwctGgL8QBJbhSRfJV+LEhCg9FqVoVn/ctc5j1xO1
s/RPM8Lnc0vl2OxgzmTJLwV4C1sQZE+rqRulGbmdavZB5qTyn7zQDa/2+6ub
skofyRa8CtqImlgpWXh/QI/Ie7cYQXgYfAEo7Q4NSfJf38ea5bc/lbW2Mu9F
veYR5H5YrfkkCBASM9GTa/Mz5Lqa/jny0yhwwvEf+xoMSIPZGMEli4GU+fn3
teHqKOUoyWIj88uOCt2Nxxh5VR+mEtwUTKHeuTG/RT9C62VcYAEmyJJ5kTvH
99iyP8RVtVrkUwnqXpNjFnTz4BauKgU8A6bCzvvte7K0cUq2veohvpWOWxO6
LuaSIdHn0M7ikqsP3gtvU8qEx1eXyTfED/2Foz3ygJcROyKrfFuqQnoQ/0Gc
na9Yr+GrcvqcMXAoNYhXDSPRWRF8E1Sh8rzMlenxVF93+G+ZNnCUh+E6YhzP
RDpSi3R+KIWqjrq8VZziXWzmAuMVRvfip6bkIIobf5ELZHYSwSh8rfWRZAGC
A3zUNaongj0Jydsq96kfoig1YtCZKGt4wMhRq8QXzZ0ea80DrnAEpfbw1TMz
RqHN6Lwtywxs5pXMbHnJ2gVLN83eOvKSD/FUHsbAXuOE7KWdJR1H4X5RyLMl
etg7h3iC5gvKxoHlppFlOGwzHXM5pQDU+xVdl767sG/OI8uELgbo6APrWG9W
wK78EOg7I/3sF5ys1tADSVnxPCYZHcphcRlyayYVwrf0gTUXBhQP/jmzLOdh
9ILrGXAIabb4ZVraaKidju67qaWwPMcadZStTiDuhZwSzMq34PyWpcn/GdHg
GeCPUG4GZXyyDHOsEaKshz9P4rAQ6lLOIs1W2hzghkKsZI7smikWjDPeCdk1
5xFmBOyf2aBLUpxLB3Dp0pAD3+kMR7YIPr9hMUL+bGmuDmR/HpWcLlseMYBQ
gB7Dd3vn2ICIHoGYfBW+3vmesfshOZoYItqdzS5u4mbUTMHbjbHA9MXUzfDF
QeSrglRQpBzI6DX3guK7ea3WuCg4bCwpvOwxLHzPuGKBTD0Hyh0fcXp6IR7L
YB1idmU22xiFAggeo346k94Roc1MRAcpFnKjOLoREpolXxhI+OPF9MT6lfgn
G8ztYeT3tYE+Ox/Zes1yO+FTZOaQc8vCKndHvuBCx1fp6XVfTwnGDfCOiGw/
5j0yJjLyCY0b3KWAi1sE0Nvp3WtTV3Fc9QyLz2cCOuCrAQKa3lHKwItn1zz/
l8kBPe+cExBuoeFotGW1V+jj/JDsgzSV8k5L6TdYKDwLfFOH5i0/KUa83ysN
BQ59pVkfRdmyPxdLnS5AWfPg5XDxcGSLCySeto2GIKSlgHb+jLRA3t09Me3V
k0mB4SEqjhSYteEVzuapzxPhd73iIpcjv3nJcZK6F6rvAniy5GtKCuOpBERz
7YTjx14x6mLSsuF/WY9tJ2MPx80+1XyhA1Sl4Re9jxVbj0sCfjKfCq9p6GdJ
pCeYMq7Xaqsqieh9Jv3NJM+ZYaYLWlayJ0UPjAjTf+RZFxkfeatT2mwMh4l9
g4240UmEAyUXrq0ykoMuGFGA7rAdSov8Cw9C4GIHCcRYVaAQPFQGDhjIeseS
ATj5wiPlkt9lcRptSCjRs/M5+F3myGh1JElBM/KmDexfVeDlPU6+LOqTyx3l
MGdkyNXA5hM7U6bnWMXdFlTy045+ee/dJqlpm0bH5qTFnEif4MXymDQBd06m
CKFh+1D5S2buUTQ9XqKZCzcUSzX0KEnki//H8j5GP3VAwdhe1Zki1jBSBXYH
zMAlLbqfH7NHl20SHtdmh53ATDM6D2Gj9MKMf5uDGvRQbJS7XrnYnJvGEANq
twGlg3DZFno9c4UVyaw5tmH7XAbadnVSo36+wiaUmMtHbzcnwTMdW3WNKpsV
Cyu4K7MS+ZIqqIOCXrthhhQrcnj1Rv/G+SZBkBiGxfRzr2/D9WEJJy0YyqHW
DV+xd4HxE9O8vS8ZBF6WSuCzG34KXtmrHRuYgeIbHeDvlghxcr9kpueLxeGE
T35JMu2pwRmN2l3qhPSioLIBrijnoNRjfiuJ4f2abd/UU3bvFWc8Ptcz4JFe
6RhqpV331lpbXG+iCfyP1r0r5QZQKjP0ndPHvQP4SQ1fhOpljC7nJ7RqWGpi
Wj52F3B/YwrHj80gp5YOPAOug30kNwNz3i3+3BzMzq6MN82d8svrxqqvXxVP
2BfJZ2CVnHA4rRdZe0hyqOo7BclwwGidofqLjmFNuu2+hxN18JQ/t4j73ZHB
fwGD2pNz/dMxWWXg6hA5Gv/bqi44gBWFELUlRKHOeZPQO1mOdHKl3AB/2TC2
nOmxow21CjJ7dsk0iQidPfW4wLDRmFG/4gIPzrBZrdP+4gm7wi8yZQu3K7wS
XNYxAx8VYpkTmzBTjfmYa8tegnmxjlyhTpzzef8PE9nYyjxCAwaACNV6Yryo
JQZat95pQDRc8WxqzgCn5QptReEItSMtEAc9H1j96NTnFUPnvZ3Mpir6kJaw
Ql2uh0V8pO5bzTr5pVYSvQvAfuggEQDUlSzUr6l7CG6CY0PknOfszLugqkr3
XGpmAW/8L+B03MgCCAzVrmWtfvSPwT5ijUfW3jgofoWU8xRJDZ2BGGu2eXQT
ArDpqSFQuAgfCbHPdMod0jFe//MNoCcAZ4fX0eEbHrK32MbStrgxPKUStKFU
PoeTN63fqvpWOWXs8pg7UC1R1zoXN9A0kpwdCo5ZpHcE5v4EXyLYQtJcLT3o
iX9JYMnWSr7oO2aN4Vh+Pi6pWLGLOSJp/VMn2E0yaHTDYoPg7u2xhcyZl323
hTSeatHQmUU4/FHGe1TxNXraNgkfrrFqDaFXToSLgR6i2HJECq1z8KklXjsk
cj2fAWzZqUKAeDsGF7OHJGw4bjwSUbsuaqvue2i9oOGg5TfF736EPMRw89pR
4NEBI2j4fyKdKqAKDiGDvg339XGADKAzNP1FFTMHFKBFb5OoSoQPOgs/9oxS
3yQzhVH8bgUZK/WFua8XqI2gBvcLqgwVXIkj9wlm1aj2bzCvu7kpXdgTbTcY
AkecWwWOQxZHX5NIq0kxLdJujqO3dydvsMBX+ZZOxAOC6GEo84wodRwmzY1b
L7uzgAUSEr7phHdPcox5dvwcNY2OOSvzMhA+Yf3rh9JDCdIJrBpZLAiy/5A9
ZUorRZ8fmIIFJvCrGH/XqqbnpWX7iRxC+Y4epPHvwm8DWXCR97US+AL3YF2K
vVC2jQxsQ9CHy9uddtkoa1zFxH75arq4y6e28stGLlkZlzLJgf2HkpXH1QB5
JQPNfM7Y7fS+VKQPnPDkvyBdl0wdlYz68pvQyVHd1nhA/gJfC4XaxgKkyNjK
8ypTV2gvvtvruC3X1XEGYrmDf50cZwRRiZijo+bNr9BLBPyKokUt5tSBQsdH
0t2QGQEti9n4TykJNi/pvK4HFODqMcN4t6/WHxwDnoT2REBbFMmJIGdiQMlM
QbZCm+M1qGp+yKGr5cvjSxa0KLiGJWP1dC1e6szUguaZCeErwVZpq+NWmqc+
x9koDo3qneTRvsQpKvlqmPOAB8213TZUw9r6MhekvDrD2TUhZOIPi+XWUXGn
QGLxJNRVmpsrjrIP50cItTQxcf62ziK5OcCy0/hOdH+TZIwypv4zrnue1SwI
FkFmPbjcFjiWV5ctIWcjYDuCNfGqA/xnvxvEjYb6elOKvfd0mPxrDdQWDdBt
/UfpZD7+f5fWgXUyGpvdpFSaCxCaoDfNAY+Q7q3wpohX6q/eRdjpnRDBt9R9
2uA7wjbWxFMRox6a6pWD6HHmQ/JE4V+Z1v0ObjySm3JjS8jJ4Hx/BOtcHBPr
gpFgUPb180JhoYeqTl9VMguhq6ogjZWnTD1nzevS9DRkuW7B/gCAynZbmODb
XkkMm3QMFjgnnhmJGBn3i9BJNWJ95mG7FiSuwPwkvxBhQBhMd1NXXwNCCLyL
C8KSeZX8mTiUx2noaEq5khVZ6ZKY8kxzEzh3mteS738jGLVv/FeTiyk1tlXc
EIFUOOObGfZNwTOGSA/IYHsF5ynTsjKTwxiwBvvz/FX4dNz9NFagImg0F5pR
TFKMQuwzakQ2hnoIjqwUt/R3tc0K1AbKIK1md2Q4gM6nNUv9+8I+uIFmFXiQ
LX0fyJSz2MSr6V+FcCE5lgwfbPnJuE8WsxOpqjyI6r2RZOZhuJgHe6EhxQtg
HxpqRRyFmJrMPf7CIhuVPA31purYxiuRpsU37wKsvigvjA1LJOA8TNdbKdhk
+AfOJGAuaSG76zJPm4NFMpyL8HGdqFWIuXLkIkh8oJjE66Zw7OAKGUT1HDUp
z5uqgx5NX177IzUjol/czdOEo4xe+bU5g6Wzj/7fYD4tVUCcXfV3lwDJmJu5
4z7aaXBAUmmTAx6NcGZKcEZzFRkrzn8qCor41CFNV34yvNR/56uJNRoH3Ac8
z0oKwJ7ZiXVuC5FjZUOnruKbthykXXe51pdeta6E9QRq5oQjfRg3D5bSJqU5
Z9fOowz7C9kFwJshnO1jzQ9OhSYrKqwoAWOKLpqhkAMu9F23TTQMt6Vljw/c
fbNBoRLY1LYhTxsulToJ7q9ciney86vBiuhKXws4vLquUqQAyzCj7GwFctiL
6AxCosjx8ZqVTj0tkUuU7hYFGOZZDcdEDYBoJ9c71KqFF2FG/uwHXtBVcz6c
/shKgXXSDNGgD9NaqrwEMKG5T/UwELRmJufUmjkPmhqFOf62/hJFpM8w2gqE
4Z3arZCwxQJ/oKNqrl9e5hI6u5A1A7gRfGR3ZgGM3thdTfv/aYRTM/dNw15K
H/m0Qbg30J9x6wH+J0IZK4S6FjbwtlQHVcvsVpWMu/D3aJf4TQOfESMJwSN4
p5lmLWPzfEftoG8yrsGckCn3A4SOG50yfH/I2HLmo9gVeHiKSjbWmXhUaslI
Xvs7TpP309tZ7KnFbbQ67JtgUHKGHHamfqU+n/j1snHrVheUPdueQZMdoni3
BQEPC0rD7Q6oZ2iiWP8zUst+1qGrwe8vasDJTTdtiEM1F4trYZK91seaSQJL
fQ72t75DlMNYJPrUErja9rY3dFBNEoJPTZVN4xHGq8gpRGsn1xWLjcnLtXPP
/XFVnI4T/dLS0HGC/jY2YZmZweiuEhucGoXI86N6inIa/o42hMW/fMgEBbWL
X3ke095R5XMQ3kbP6Q5MVxi5KZfXt7CU2gmrqnCijPdXCG4Umx2ua1K6wAPM
BDcN6NX3bQfzYma7/oeQu2u2wlvWoPTXor6DGBQZaqyeNB9cI4yAiqNRFTUk
0Xa9CWHRchKzWcHewi6iekV82DLV2clKislDGSgWtHval6lByCFU/Id0zTJ7
sFr9zj/8C//wFD84foKcqw48p0bPLF8CL/r3tlQFZbqilW6Pdk57ekVQLmJ+
6UtW4fS+HOCQ4gaWkBOMJ0Hc4U+IhasptZqiIbNPnSRu8ZrPxtIyqKCscWhT
rkZcq/DFYHxJUYmz1jKkzXDp8jDyTP5pofZvkJQpE0gz6qK4bmZRu9CnQ3HE
NrVYbzBi8r2O28gB7PZiz/4YoWi7lo/4UBj4HzIRlXjamPJQ5WyqBE1huIK3
KhOxiu9oFIyQ8BEP1rgKTfPkZQH9T0Kf70TqnPJjwvapiGsrsEwBbFlrmMr5
OX+2ptSj1Y649puSkXxhExq6TY3hvqcSe7g0uhfpc1u5XVSYVt8BMxB+iYeH
SCzKHaNNgLKZFuAzxYGDF8Al1WOdyv3eIfjdC9w6KFrs/bDZyCTJowjNbMQD
EJtt/I0hI/rx5F4mT0Wy2ivhrPD3hewsKaEUOEKEw2cCe/JXjGkN4tMpNKYS
INJzjX8zHFP/qP9CcJ64K52bH5EBsqC5RFmjjcoaIOvid0Ot9Y7kn8lippKJ
9Mgjj9lNZyc/e3xot51jw619SjiUD4amOM8toWL28tECXpcO35f9abFy+DB8
j1tvg3NcrEB85XO8elFuoHVCl/0fUIn1wtEqq+pYiTM6vtR0TU7LyNh9ptg4
gIwUUwfukpZ4SgcHBUyurig6Ziw/ACUIJ0jchYZwxaPvnYJsMTbP8QkamZ05
qSI8xcjXR69VxYAN+z1uk7w9tQNAFCKF91Acfk8WVp4CZETmXH/5rF6o6wLV
YFg8RIz9eqD0TOcWv9+dcah0usoLJ1QzNatFg2p/SnuVzEvxiqkOa4yQCpUP
VATfy2nec1Fn7g59vf94M72NOgYbHa2fJGjQlrVGIF2nTdkBiYy/dg9NAMv5
65VuZpE44j/7MkWXnp9yyglw+s5ZkE2+HHOVppmaGMCFu5cDiJZ97Et0Ip2r
Ut7c40x47CKs4rnQOPwTJhvFjm4KcwXjLLjHahkaovFsdZHW9zDpQhLQJ3XC
uIbOtKNU0K339Wmds9YVLvPVdzsH5v0EyQJeFOz5NUy4YUBvKUOYIcMB70E/
4Ons70AE/5tbx5HzoZd4O1qWpeeSTQXC/YUF8IGfXnsg0OlF7X8RdCYH3vmc
VSdY4hbFljo6Ksx2CaLtNtRlNulwQg9E6yKo1dfU4YYIsot0z+YXO/QDYKkg
iBZJBiFBzqpvy6Y2V2SsvC2eUDcgYGTEtCR4hfC6CJBNb3Pi18+1ReRlPomi
cFwkrWWQ3JJX+0k4/gs/7PCDYoN1iSXWdQjO3hjOD+Co/dvQbDMHppFzwQym
RS0R2k4T5HUf/CVzzV1niiWFYiV4dgTaaRL5iyKQvzVhWw0pgy5Xw0J2ka0g
u5yDT4BxGXgx28NclwNAfGdqn9Go2emiYIENUT3/KHGZev+APcqXyiD0TTDx
+5ns2gAPyLd0lnLwt3pha6M9N7zXcvNJf+Dg2K1uAKj6N+ltYwjcqDOrgLCc
msBJ874qnQZn3ujUwo6dBjOPTamuvnXgHnqGSH38nF51RrRh2H6TxkUlV0KI
wIOmFS8DJ7p+DeIsF0KHhUEbR4vs5IIX2wfb6dKCyk3+9GjvgiFqoTAgsvSr
oHKTkOLtUCPgxxfgLvGILhNMpwKdtivwQVRjk0dpIUYSACiXGZAAr/buLTMW
3fO04T1WVvAjWYWCnUFmNbwT99hxLtDQTPoVOZONmlEXQ1UZoV3dSHSBmb7I
d5+pxOyBLekBTC/3OnCOUCh5qIam5MMCNCqa7YvNoYnGTLexI16A3F4F69rN
5GJ9xde8AO/WA3rhM31ga3hFNtEmheFaeCt2HuDg/HbtdN3/7ZPg2+dc9Ior
Z5XGDwp2Xi7joACEDksg0eC1EotcN7XdpeJs8+HNzMc0tZX8h6Y38aM+4ehb
pwSEoptPTl1bZW57bJDgO5NvTqZ098yFygg0wyYvK3BLcTDXtUul3OhGSWdS
goNYdsbfYJguDVJbO1i27hxNx/CfLLhCET+0cSFnlauvwZTfkWeYjCfBHr3A
lbI31i+7W/cvMpo/dnJRf/VA0/HitSoRB5FuKzEaJlC2wLXDiRCPgeALJdc8
DaBC7jvs6E6ERgykMRERUBdtii+gE93LJffZ+T6hb55tGFBctXMhGSyJLia/
ubM1G/PKrFSWFv0uLZP/DCfv69qBsOIEijsQDRU9ctLK1+Kj11jYMN6iXfkq
fiC7/Hxe0IXMMmxfn16l/lJwm0bZUg4eWF5FZq1KkIcWL3UPC7p/hxqAf7t6
OnHFnvMYaZQUWCYOYldd1uMTR6w1Nnc+CSXahOHleShaNic3N+wi1zw3jsoI
wFwEvDphHYOiN0LIT1/10mryJcRGTTWTy5azDmkJVc8+mV7M21RXsrPV1PLo
dut+YhrU18yF2QKhF0/79I0S5utzSzYVm5dOFe3beIs4RMoq/0BoD/qfV/Rs
0HAqgTT3h5tkWCZ1bO9OPErA6E+e6OBF2z5+7AD/sXm28tut6SbibRFo+1Cu
1tpFd2OZkm9kfYnBGDNxXG+N7XM+oK0M0/vniI9y8Afh0dltKCd7cTKR10ci
frkD0Lr1ZAssZoTWZVzPhykpmZbKdc5C3mqGhxxotjrqxJaOT919pnBHexPX
FAYGoPJIHSofRUs3NaFviNYABNW59LjKEMT4RNVqZinbuDjrDF9ZJnBhEyhJ
q3yt6FhBgMnJFk+CN6bJvjhKSUp74ZhnD+n335BzDePiwFVhpgF6ewuSaAhR
1Ih/yT/t0OYkr4hQG01elPGNbTjw8w4iw1RVYaaa0Dt00q85ZHZTADXpdyr4
yuwfyeOUg7/RblYTRN7KgfZKgLKa0PELxq2yWjWqGBFsqaCsQ5YKsdhtIRLF
3qTrxCKl5izpjejwmKOedenj/S2pD4groePDxp1HwGTcEDNsTnC7ZvVyEijU
G4wWJdr7At71cOtIcpXmBp+y45JqXixUGiAllxYNQJYaeZGMp1j51tIpF65o
+GrthmDONfEQvsOlTNcAyIzJNX84sIKwxfQDcaNt1/x38+PoQpz3lHHSGMj3
RT39zCxKJG3KFzdcCBoHf4kbPvaNvEICZxHdgNNx04JsNL5U9+yMEVL3RKlE
N0niz9WHOxE1r/mlif5XgQIkmiAmWP7ZQ1oPcEjPni0BZp6aTAqe93zaRpXV
vVF1KdfkyofcNNpkbqBUwBodAx/Nc+3/VuQr8U3CfQUZYaD0dpoxnqSEUCp6
q6z/xxgoewLqtE3uJSytl6or/jqioavt0PXsGSwfmqmVmf/j7Mx1A+4tAtrz
ZuQPbhq3hDI6Iz4ru3cOEIsautCbhHcwDnQiZKJsj0HdTJwLuPgRf02fsh73
aiHkybUwaJKzLnn/DSIGY8Ujf9IG41Fbm1a7JfK9ZFWYIna/aElXY8Cqldjp
r0NvV1ZBG3hy0s0rYNxJliutTrKv62FfSKAeFWvnBy4AQwznJbx6mDnn7HNP
HecGTFC5ZTxW9gpGwk2ddsuFYPKwEcAq+1k+Pw4kMzofmaQZtAQ6peT0XlaW
Du49f3JV+60EmYaQU+mNzmXx4BGjSKqJ3acf9JqHciQAF4MWOBhChFBrFRJj
OAybG/PVbD9tyApdWVihusnKKOMrPxBsyj9+KQUfIF9kfF3MeF9DzAGrJZX+
HzsOj/8sD8ZQXAQWH8cCVBbOSiyxlEmo5P3s9rzlVl1UJ0HytvPx790ANwRb
rZl1QW7SIN1oeFnIvSuNW3fjTSdnD5/MWMECKWzZJRy91op0unuk6QC7nuUc
8uBsQOdsXui8eGnbBbQ8pja57surJ2D4jw/pKFqkSX+mATZ3jUL5cbLdj27F
UtpDxo//EIGcLlLlRxtUSDucjWsIIJ8rRkRhT7Ydjd4j8jH8OnUjG429g8sQ
ch7/2VpXX1Xf2lUx5EWxbKSDgXmLze5Rz2SIrDJiUt6rPqXwdjinpLg6pRDT
cS4PRTf/k8IUQxvRVmDSA3TzhoBQvT+/6ZIxjck8Cinv5PqK/WRvbyMxQ7Yl
6VzA8Nduh8+qIpZhkNe1hkpXKSCQvjJSr+fMeyOIvkiv1M9fBxNP0kMX2LCD
HczJWOsQFimgevNqV74IZYNay5SwRRMef73ywIeYKycEpIMUDsmpTZ2yci7w
kDhhV2AsfqRcmSUzsWU8FXxJDgrSX6ZVSd2sVztHSzSx2gsGbvuN1Eieb9pv
jZ1DccxvWeYQvJiJtyyc8BH3u7GM7fIS+SU8YpZ3rhIuDLYBVRj3ZXmXv+25
BSG/ia2bbjeRxZt0xj3YFxESxgFfs8/T1lL0TwQlcgxKNJpJBD+jyIOprohx
NRVx+Up+aQIRxBg54YxJ73AAjajY/HDiK62uSkky1iJpFFeIw10HLc3f88VC
t7C8uJ+5WHvY7mEokoRbvn092y+y+xqESlKak1WmZZEAtlD08wehuvZaGUJ3
h/8kDBwEyNpOnmENZ2O0Vf/TFqpBA4/rF4zbKa0CfgUv9CXUjDGTcSYhW9z8
j0NhfYPseDrAKztFMVWdAmAzh0XCpLCsCaTxxHP+rH0NMR2RY5qOdwoY9TDZ
2yB7XTXJD+OZMFDKJYrWkdVRsoAtuAg2+/timP1q4cIAPwWH5wCx/TgnCwlU
XhPX/OgltN7y5eb1T5gm+Yle5+c2uNMRLhFEUkFLE2R3w92M+1a9aXGhzoZt
Pz++fBx2AAkZN8ord0izAhRzkLPbVkWf8tmjoXNl+SExP8hLKeDzWshyFinz
DDL9aJwk0MoHi9v6xoHHq0xlTuKz2ioclR3Gy0xO0yYcz2yTvsUOqv1McEJ/
yO6k2+yCevnFkY7WwtSRpf+eG55S1Yjrqt/cNcYBlZnI43EAQ126QBVm701E
7m3AVDXvorT7RHR5Vi/E74AfMnuTWo0+M2mOa+uNGB7+VTB/IeM/2zBH71cp
R6V2cUrO3zJ/pDYNX+X2iki1EClZJ+/oeFATL6m314BhszuKCnKM2Y+JPtRE
8iRd2t2TwZajhBjT8uNY6gWtXt3lQ/k+VlSCmx1jGBWE/EuckUPQDUIfRbv8
5siAPm8UhrAp1SdT5wUD10SuullQa5k9xeGNHfjsXj+xcY2qN7fMV25Xa8Pz
qFVYCpY/qlwqwT9R2Xmnt1enPFPeCACIFGO8RoTDA9yB+KXyqgzGwO5IpuC0
+q+WIydjPe/p5lbGhjh5ed3bZUFfjHl47gzx4x/lFgA88guRBKhCVg4OfKxo
9zmLKg6mP1SJO7GW0RIXSJTDhwprgvfG718YPe6LivmvZaPJEc4QHsNvGMnu
xEyQ+icssvKiqC1KuD6vbEoq3J6vvcYlrb75opAxhBTZ+0A+I0W0yjqcStSV
CID6cmJxoDqBigEfrrxadXbnmVVEangPDIK7L5QxdnFZ6Sr5f8lCRlurtYrN
I6b6msgI58UbRlSjzgWr54N6BjUe/n10ZTpoCQb/k76gUJcg97938tZ49raL
uSyT8CQ7kut1x8Nqe47DlOFxXOmjD0TX4XZHe9bs5HKTFbNMPd57Vlh4bkcC
dqoPnVVrPhJC37ubECMhAFbQcpZSqlq64gJrqyv4YkNk3Wq16or9DeStBrXu
EdM3GiZga+QgtFrPYPCdWM4f7SxzOe5N+wBn9gMWiZboH6RaX3pi8JZQJA1m
N+1IaxzyfUcUhkATdlefsTspdh1l8XU4k8O6P+TV/irqlk6NxGUnl6BzMlcC
zQ9HBnK4+P73s4uMYKPjZOxZLLNR69+JU2EMUSNs/wDoUlXwp7PRlmhrmC8B
sxq2FBt/pf5gYOM8/xXcHnuERkKW2UFjVJIOPB1aM+w9dRJ5onwzMdNPERKk
bbuNl2X5IND01RJNKb4/NKIs+NGb6Xver7oQe0jR7mPDRF3KOc8ZcNdzd13l
9ttag4JBCTy7DiE0G2BIqJkU5PfL8nwBzbp19F8ZjftJISXN7Ztl9gVAiJTb
/I+Wa9i1hjC8H8kWZKutMgNFBnyqnfK5jwGnkqGLBMbxivQlfeTrZ9QCnE1z
ry2pbfppqrYJlR4C86Z9bpWFOEhzvYlCzQRfQXAtd8SHzizCQjJp505QY6UV
8as0m2dr8jEpOhlc4S74MA/cdIvnury0D/iOA6QNZ3eP0ums+gZKFlubHCNA
x7vmgm5wN3rDJ1xiu+oLOcoioF2Fd057LjEHOvJkBXLYjR7PO5deD+7tWbX/
urliuWPSmbVQhs2dbfvw4Ih9m2hfOk+o01L5cmFYSFn2LtsZquAWR8ot4mHM
UlDRjfGhKDzZwFX962GnuVSeRVaqT/pTR4Xp+bTXV/t0Jmf6l6maYqEoQkk/
Q59E0Ad7ALKovfPc8RzaWskdXbSihIZ60xvoEqQE3JGdadnRehM3/sJBCQfR
C9wAzBgbavgrmdhk4toZFi7/3M24z6aMxDJkrEByYHGsMc1ThAAwwJWkn4w5
nD/hItVfCSXNgbKwaBIPgUGzA0DvQ8kqv/Jw1RJO8SJt2JQU/zZRB7h5fRhw
Fnf56Gm6j+j6mk6bkm9yx6VA74J64ucS0Z1tZQ0UFRD9b9xaFJ652N4R2I/q
lqEp5ahg4Z8Vn4jrMQnhgJnoKSN+C0MXDVNzPF493CcEFN9v+4MqPVYPYUjA
F3JE3c8ttAp8ELZq3I5vmOMou0LU6luYUH8eJRNs9FezpLdriV4T2TiRo/Wa
BEXV+HiIalFIlMnLL40bGfT/bMjoZywNj4FWctW8GVRO0btUuPc5wEgNy7a8
HtZbOx102CWoDIhzI4GkkyfNwrsCx3s3+DB4Q5c6pSANOfQxj/Oh+SmVdu98
pY+BcABhankmwVe075ESt8ewV+pptT5FjFVxLI1Y0jwsrgIyl7Xs3jS05J8f
dGOekE8Atb4t4yoMEYAow1DV7VnkVVuIIafPQk0XaqOmnOJTTZRLhRtLQFqm
u9e+svpeyMkGNhRzlepwTOYzvRqofb4xIpsfb68ZpF+0xlgvKHbsfUtuwDJG
WGdn4R3Fsch57kgYG1sNLU7pcFAAdxIJPiQ9D3gaL6TPS63x0BDrNMFLQZTd
EMm3o8OOdfYhqVD8Qwjbj7I9b/osZ3XLBz67Pp+yOfo5tsg84ZkgRMuKfSzn
4GPEVT2RBX8rx/IDTBrdVasOIBDaRaROKlgwqISlItv3WIyKzSd3SQ1sK7gZ
WyQZwF/pc3FarYucbIEHmeTDiWXExW+7GhUSeqTZcGfP0m28Y0TEG/UmgThC
AUAMr59NygcOTh9lK2nRGzHftLy24S7lGJgtSEFJZiPzd+tOSzZLFpYj8yqv
PZ79W8+TTxymx8rOAP1MJhNX7FW2jUbXFYZLrQdG530/T2HLfFe3rYXze8Yd
ZleDrgkw8tkQurAxrABUxjRXg12A4VrHLpDEUDUd1FfjqUPbOJjufsvTZvtz
MIvTBB7xqjQeppUNtt61MouDxCxraLGeoZLQyCO4nHKjzaEju1B4qFi5Usly
jFQMbSNp2Rm64HwRJI5fq92fTSHLsgUNSeDpwcqHh/9HVIwc2RkkWQi843IQ
GaplGq6+sigbSJ4ZEbhm/Qx3nttZdEiGMY18SxckMR6+/IA0XYP4VTwFVpuJ
RYacGPJXb1cGGBuKArQI2RcUgqTMxNOpYoCWwfun6S98YbjG52mdjnbW4Rle
hbn9DZqjHQTfnn9Nli/aVeSwrgyyGMCvo2ksALYOGxvL3+eOhiJRm1WbbxUx
D8fRLj49n9sj7qtna+r2WdLNSrZJSPuAH01H8tPyJZ6VF5XIIo9BFn2W4f6i
LbpzZS6NDgv/4+n6gC2VoyLjoQeAwCIKGOnhiWRjZhIAWL+UFGw/4DEtv9hu
EKzZAQQsJpL8Vg3gHm0F+jucKiG2cz+lLwcukGSXqO7LGDJY/ZRMhb1Rr3Qr
7WihJlzDLK8YT7Vv7EHZx+BQzQR3YIz2lc5v9JhhC4Xf8dl3/z7DNwKPqI9I
+W/dXIKzsk/6m3BecIcRfgmc+FqzZ+CFM8vYpiFwRNCh45RJZttv2FIgKhVk
DxnuRP4HpaBNpsVloa5fWgnrMHY3x0chZN1VDeUOfNObNWG8J3vpX11Fy7k4
FCgAaRzBpjkTzxhFqF2tKJV10r1YCTz/PampgdDGXCMycYbdkZKpqOrhYRXN
i5UHrLWUXrXXxxYcxxZQiweZcRpVulfEdPiHtmM9MZDyF4r4L2ZGHr+mieHJ
JChf9YNv3c6p3gkbHr70frJDTV/5RE9VGXRiRUekNt4tLg1f0MdlkyPa0Tcv
oJJomjvtTUezEpHDewBKL5zf9wHoqZ79Vjwn2qc4Dqie4eczlczMFSckiUAN
ycW74vZ63uLUI336GCQiJAUKEFtVU1BDz5H8nouJtOZH5uvr25nhL//KrrVs
mYCgD/qTwW3/HkKUf+CuWRvzL2RTY2g07IRt8TnnMZG9KDmRM2IXyYLtQYyD
K3qdmI+SZwrrsL8/w0JjHnonxLTiY20akKN/gnqxTClQ/t37fcrW39yvwcML
BqOgxJfqumFo5Bb1KmWXdVBY8c2E2MTVtzkGBlAb2MBuGE/8RDbJqdDtZXCN
eTpdJPn/CP0DmPGRmGcv67HW2b1TD4yvFRPcmLBwgcoPlzLOL5xmyMqgwPQ1
WPOXJU2w+4y/UFRhdTs29HH9y0PHhsEscsHl7p3KXoaZHP/O2aNeIgUuUPQ3
nzuTbAKN/vcrwjzolSBkpYJsr6Uu8NLIXJuVFZbFHS5+wyZlAGls5lS//8RW
c+ntKkiqVPZ9JgGeHjHcz4CwU6NcAfxxyIPx58wlh+ITw2Soq8XnY96IN/lF
WsHQOwQbFa2E02HHJyBMlH/9ChQtfXesmkM23IswCl8pQK+I60CyD2TVJXX0
mZ15KTzyOEjqYt6yvL40Xnrfct/uswKmjNKnWbdgSrHe9CeSssVv2bHNqlgZ
nmOyXKEn3nepWWFJnO19lHRQmSMdIgjnD+pTnfquIy+Q0Ttiw7scVRGAujbP
gvAczstHK11shq4/cjKm0edZQtIj6+5l7PgLAyesCarHYISq1jMEVeu7uTN2
7wvknsRw56L2CpmX9QXCpGsz8/D6kx1Y7n+AZDbGI7JcFABkHTx+vbm2YNMN
NbI5sxhPe+FBjRLm+il7mFpN+KV1wdrxxKYRHF+CxpMS2SMyc5j7kw7uyYpG
Kv826E7rK/he0zrRQdYDqHaIzcC5x8YhpuQDI2QD47syP3fz9VZOzVBJHaKP
GIUIQwUMES2wM8ed59sSm4I/F4HvDmqexx64ofeaZ8FbqL0YiBy7EWj8Mz9X
Sqfz8A77geNxBd7hJCLmROQNoDqnOoWPDbMpiQM7De16RyFY6sNwMW7X+6KH
qFCjEZERbY5cHK4YehTwDTtqwJcrucqOvX6+bSF2XMnKgl3Qt3OqgihRi8PB
spVOCBanvcrvdeDAkHWLnk8XoK81l5GlXmyFyXgZ5NnIK6/AxT2I76S9iY54
cVtRslrXvyZw8T9P0kA3VeCAxcuf5gO1PhEElpwcqhHUwaDjxyv993ySBxQW
UUv+kqBw7xGa0FG0F75Wg9JpjNcOUWfu4jLko0f4rHRJ+x2uUX6wwnWt9v1m
14NSj047IJG9/84ofgr2PtccRVfz3TdZ6YpRx19YcMhggiTD1lUoS/108x4m
ELapw9PZg5D+LlzR5Ta8IefDyuqF41ZCpoqJH0sM+NmnHKqbvZ0t+0ugeQag
c2Kcn84ZYQ0UdWdDioDeudd0uvhDPkoVBErghC1LLxbfqAGxFJEs6ziNHS1A
Hq2tmhrJC5NC9W/wGjIj8MQCcdqi0HKzj3DNHQug7wxOzIenbAUZonY69dRN
qzbSr0+vZRJQ+6Bd+O+RmgF49DPK1yCmHwDaJJi3mQpgze289jR1yGIbR5zc
UbwttyY6Z6QfHMLat8viBQoGxNMpggtTZY8DUKJ1gG9DusFSk8Jcg1rD6i8v
hgdVNI+lHTaW4JS6ybsN2LaAGnVxxNOFPjt9ldP5bUIKHuYoSNphbb25LCMs
JkRqrfvB70ihNUtaKf19GLwEQnpv+KjQGTxwZQrx2Eg+M5/MkX0EMiU4I58d
kX+WOrmNZSS+7DSMj16pJOUAOhh2LGj+wQcjbUgGKXER4ln07Dl8zn+s86Q7
wVBkOSsAAuQMhS6jn2NplqPwGe6/ebO4nhbl76JnaSAYb6Ro+E1DynQOYlou
vYIp4S9O3JfWSYkXAj+S9e5cEsQ9WLrXGD0SsoUgcIPB8wFFex5fq9uswPvE
Nz+0N+0Fvo2I/NaxeVdc43MEtyo9r4iqgU+hRWqkHv8ScWJzYIcHLzMHzjOT
h2ni6/DSaMWVXbacQ0aiLwQFHpqImWgAI4gAZNcmEbub1LKxmmHgO/T/x09L
PbUTGC9FwNjt4SmXCjHRFhYs16TJCPAoEPt06EUURZ8Zj+sSrOPTkn/gHBbT
sxDROSvfU9bl0sKix8APqww7sgmxJenKI2GSobjDqvpisjHUoIfMEn21otx7
3dLNUmShQYvrqbez1DQSJ/XkcNptBP5KJRMrczIJi6LxWR4YMYSEI75JYqp+
+1gsO9UyUf+shsSGpfwSMd0y/MfAHIRqXLsMjK4SXkOYiCEuVmIbr5zyqSq9
GZkBVci0KT/0QWN8TgugqOp56omEAsSCcWkJ0nWxP0pXQhpviVjPliqi3y5o
BV24W41g/sY3tIPnqknUIv2pgC4nl2L18QqNliQzBGuk2vAM7qH1GpsNL7Vv
25RdcRcO91HFp7YRxJCNzF2Y23hDBveD/gTRDFaCrUoAR0Rl/TYPRhXERF0N
cdUywcv0kOevtKIYYfxLSMRV06ofCcmknEogENi1tRRmydW2vrSjM9nQsfk0
HgtVUuL18GHYOmgCvJKAUySoduZop1Uhst0bjDqt+QQyV0LDfuZOBvU2kmHh
IBWoGMjtnVWYGaYGVV14a+/y6x/KS9XPPgDQHnOZV0aJwhhKBqoS82cgoru3
Qybi+JS0C6m5AmqPYyO+eZAEhFzjkFGqbj/+oM+qmwKAbMK0lkxTgSzThqRT
O6FAFM0CCVrjCDwLH7L1ZMJCRnYbkuNBy2GOXQElu5Oo6r2I6VZPlOBSeBXs
q3VNRDsLmkKlQRl9AeoJB3SqD73/QlXKdM6LEWR5DG5zjOvKD43/ZBcpwRTf
95LMP5pjad4TqXJ6/ybfQQPJdRknKfPBT9XO/EnaxTO3sWVJ1NNF+SQVZG2P
vNFgDZJWkCUR6jwrucdD31cE58wng30nMT7PmeJzeH0kd8eHryfH9pHK2Jsk
NO21LbwOKLAzXyPbnwdnyjTdfXGjcJnWuS2mEkpIY9mtoMshAbUgNTIKRHzH
suk7yrcW0k7hfJJhpjlzMGDm7qhN2r98us+tBGRqxEoXhTQvmh/FqmZ+ipRd
PK9gxbdZhy9RRmA0h0UcQv2U3Gvjq2J1riDfDLHx35LdZtW3iCLqzeAYyUuk
3BPaMu/L4bHA8ARWYlnOK1R/ot3x/3rXqIF3e3b09cBLfMgnF6M2K+Onbf7S
Rmp0LlXj6Udu84/2LfeSW4qG4RxsUQLz62eznz/DhadR4WafMEtRgDnOcA7V
OYNk0gcKY7UnalWAExGlcmvXE0Kg1P5JipH809Pp8zhSx3Fr/8A9WXS3O8da
O+9QMqt/2jXFrVE5+SlyxFxiXmFuQvpiVFopH704ugokUhxhYERPhTz5A8Dl
F869MOjpBSch1yaQd1EbriVgZ0TE7oH5Hv38O2+Kt3Cop0RROR08714lpolB
DyHK6HAXwBZka/rYfgkxe4WmPgDKeMS5eaVY4aHvohShZ1yHsNibQaZLa4bT
qcvyDuSIyRp6hHg9kXTBIYoeiOFPEuxd93H9hP0P0voT4Y3WUe5O1DJHo/Od
ELbSrAC/NcP7NtHRZ1ndmS7Kv3pmf20QfAnkoW/TZx9wfIHB1MpQ2cjCCyg8
joXEiLDur6O9nbloKkljAJgMs6YaagTHIb4XoXlbBJ1AxdLNLn05H4xAiRzO
Qb57qvltsEXLOjBl6K68J5jIicoT+9VqU+CB6V7FfQs7eomg6l9QDwIYO2h0
8SAlPQy0SFLiJpO6EIkzP7jKXPE1P6PH603H0p9+yNVxbfc/Za2kbAH5naPA
dVxCtCQetJewGesAkeALDtMMxZVn217Og16kPy+A2SWs4zqjdRmZDDZ8zDvt
jCQxydFcAZZoKRurVULyxLv9zCoJ2T53nEzs0IfY4/RhuhfOo6c8ybLGQMqw
IV4hOJ6jv1Qc+FkZVnLLbGdGSpntq3fp7xLA/iCV3prlwNFKzl4pUwwcWFW7
i+tqJaAOdWcQgD2fu8Pf/OBQgR8c3ESVWIJtVm12tcqbvCP9tfiETNwO4bua
vEk2qgo9Yf18+h9VEdgjmRs703wS4x0kXGSwQQY687u7sNa56BQ/aIFGK4Kd
5QZtVE6lce1rXPu0WKjSmV9LSlAzi9BdWx7yWer/3RNklOPxO95W+GPrTuq9
+drH/szK0k1wfeFo8XDo2kKJWLrf+CGM4+ZlINW6R1wEnkHzXR1uAgGEN9Ts
BS1ZzqMJDG5MeDMAc75hezhKkQr42IXPkEoswZzDjOWh5bYaoAidBHyCU+GV
Pxb9IXmiaMgm3FL28oyNvt1TrtlXeicsH+3xapNe7SSDwOjWsArmIJa2KOv0
xduuRM02yJa2wbgUbrg/AGhiL/4dM4dsiOUjoAML3r2duxTDHH2BxPoGztWz
CrmsD6lXUaeB4VoXNPv0lDmyEb1pmNpSGa9AcfF3OhM9GmAH4ulMSlCEsOXh
7XDBQTjz9saY5qOffWLH4huEP2Iot0FlgSu+54jxce6wmL+uFWGSF1nea72r
QaV2iDLr0L1hbPQBetrX6WopAfPOWaWQMQDBbNTyKWDIPzTpiirGDzHyH/am
AZ60SA8oclsbGAz8efDIbx8U80kNPImDQmD01xNgfcH1s1yyYcI7T3m1c1Iq
LKy8upUV1pcbUmWplCeCl8TbHq+hCI0rod3jinTkTZcI8vJ4x407ewdXrUBz
2kWfOWV7h2eU+Vf1cCimdrwCdO5ROA14TnEQDxSFoaiNhFrS0+x9r83xzxAn
GGwmVRW5VnH/2l1YNwhZCl7aAfWk+SjbRrf3ZjhfNwcama4RsEQsc7CfCto5
Nb5fnSvEE3YUg6TmR7PCMDF5GWmJZh+qBawpDy5Vg9U78ElehRPr2aAeRPta
TpUl3L1gcoAw/v2EW+DImArMJgFeZEfl6qUyD/RgUSqU/NQTwCk0QfHazFwp
1kpVzoqWBj/B/n6IFki3K0DCfJItkM80Jm7PasY8GF8ZsgeRa7RBqPXAXI5z
MRgHDcanR0fakOBTWAcvn297vrHVtabIv4BP6/puw3rJ0GvHykhEHK7VvceN
iNSpj6RlC+TWZM3N3RRyMwJswOhgiiZB14s4kF8TNWQxPqm5wU5W+uj80En3
H2aM2gudWSjoyVtnKI1ALMv7m2D/UNZ0I0UzkwdxDvsPMpMnDMeX8pYA50i7
khOZbl+MgVh1Uo/4YDaoWQ5OCl0g+MqFhMqmhZKZoziqhd5UBemhm7wvfEyc
Kt5+QZozcKsPA+9Gy1ov90OXnZJNzWVxx5+a684ghBlTOQC4N+Mn5y5YTCYj
W25D7CRInUqNvDOx+QKJBfex6ZG+hft3hxh+Tggm4FPR2yvb2y0cuAFq/H7r
Z82WuMAzAX8aq+9jyd2TKjex7dfaHQlZzLmo+AcC0r8X/Sdh464Yq4zR5Z7e
dPN6A4v8+r1c8EI0H2oy8QunBIvrhT7vttYzU3dGAqg5tuQqEYmDpTepltoy
yAYzUWDbp1vBcdVqFZBRQKdKy6b8QqMluS2MXKaX/o3QQJg4M9eObJ05Z04E
t+xBObihlC1SuBsC5MCs+AjftgdGwOtgqHAyqcqoyU5rWHoJ2uKokWK4x7Gb
POv4l3Mo7g8DR0t+mnDhJ96AbSOBaDLfwi1vQXd1WKh4sWOTnlQRIFOeCYgY
q9wfSbGAD4wgIG2x9LqtAXFhP4y3GMU+fR+f1birtcInWhlNQrTzGr5Ity8P
agTzp/NA8n+nLlkt4X/Ykn0wqLApSeIhgjA/Wu0zzPtZMlGopFjTW6wzFb6g
opyNGuAxwrIK9wRXpzXaoT36/QT00fPtH582q/Y3Zn/XsUjZJ54c1ae2MQ9t
vICPqktKRP6M0nYhz2V3i07PgJpTDCIi0PGlf/Z7wWh2JeTM1E6k7D/WGyJQ
7BuGwHP+FUWVtiFKkntcDJDSeZo2+XQg8+6Ed4zuL/bmm2V+QLbR2GzaTezH
Aoprjl2zYo9+dEnCcpHuRa40MwQiU+gtbYB00IuGlvGZDnRNQx7FM4hWY1tV
MV3sZGyu1MDsBRFAJ0cqkqBDcb5Js2pcWDCcRpHIQyzDJvnIp6O5ldPFdpDQ
i9DQnFKzsm6HPZmAY5IHzdBuI/CvgFJThRj11+AmsAqu1vXeg1tuFuGjuV3P
YnW0M84wMN/6qItgHW1I9wWODnj+UValb+zbcgjQHYypVCcknzjr9+vYWbPj
LRTCnCOVDQNnFLPk3+dvcEDYUeWvWoMyv5ptv7KcosHdu5RczpHa+scRb2Sh
wyfoulku3u6DWLpFzOXLtjPws2D4jD1FtyOJNkGRSzHivFr7o1/DdmOGORW5
T7ou8yYRGJczD0EsLHIKn68mZYZRQnGwUNRRUb70AYabG6ybptuYgD2tz54V
wZDb69XvWpABlinG/NPq7h+Xm3nPIWt8kaxxdfsk0d9PFKLCdx9yBwKz7WTV
ZJ/IE9oKo/3DiyIqaFjNH3z5lIIsAJjqrgDOIJYf2/VsWTuXb7ki7KcytF18
fzPH9Rw0MtVL/Hs7x1CJ0isyctkoofslnFnFv5d23G+L9BUXr1Ur/2Em+GR2
UbUgbsZfOKLzlZTpqdkc+X/QffMkqD3/7QukYl753lWo7Hk08/tvMUILTgyG
iuC9EYe+f9+er+kh60P6ciAbE5+dEi9HITGjSvdgjUsZ7KI4z3buBmwTTb/7
absSDr2PwFg/D+/EYS0qO9WC9Cj39evpk1fsBIqq1xKBvTo1KJQG5QUqITE1
WA/NGMuKUkjlWGcBAeRRIyeq05ocJtO4PPnKL+7MUAsr+fAgbgaNVb2yVSa5
LJqADcZQZ0GtBcCqc0xRuK3197ie2N+nnOs8LEmUW11pzFem4we8Tf/1qRHF
qwFllNg8/2kk5qfdztHDHnOQ1CIwZCS0nHiTy2jBBgAlE+a/rJVeVlWLO95g
CcI3fTJtDS/LriQ4Lb5hBV3pSgpHmwtXkDZq90sQfPgnv2RkXf7taZvKyK1i
i/zraoSlK589I6Vtyh/kDK01sWM6BYhsmXdBDpNYsUmuUjr6PQW2l+v7Jn7i
Ypu2W3HvvPdbegSkW1mbrBxzIzKxe+kTtVLMb3K0XQTeUIyXFUcaAR6fspKy
Qzg+gfnNmzKF0gcmmJ1D+4T5nTtR1qspcvHAt6saLGVVGp85xEOqGzfzgw6Y
DzcjaV/Ri9OXpTyZGEwtBS+rMQ7pwuQqXljRp1KG9mG6YxR+PeGDvnltS0Ln
Uo5+f8QR7OUY0KUZn5xUBPMfUhgibNO8LLtZOjTdesuKjS6hgNYhzIDwBx/T
EsQVVAFpJ9CBLvtsafcebmcOZ3Ex9PzT065GgJ/gmB9LXMMP0FJea5gFaT7t
mNgZZS6yVb+DdwYnVduqf7N2FsbmLxbGATgRiRo4eyKux4/BRInXtx2X6SVF
PHaj7eI3aUxh89KA7fnSfaNTrPMaCsKA65GSTeSjE1zarCuF+1DylcAU3P9W
4cJOFO1Im5mWBzas+E/f2d1UQNQPff4HbPEf3AgjYT3l8yDYzPwekw33RLy9
D8QWCSiqCFx3TdfJ/X11uQPdxaUrIf2Q14hVFTV1BO9dIMZWQvp217dIFrkj
HrgFNqtGP7alg7l+z+YMksqJ9EuFpwELZwRIgrZtvnDp8R1QaPAPDsMEj9Fg
sjA8dEHGITcFlRYAtEab5I9MR5MeHOMQ+3VqNQilFYWvq7+0buIrcOgiWB5u
yK99/V+wcDIjf/1O6wtFV/CKMrBbTrRzesv+viPjufx24GozCuup+CD2QCEc
BPo9e6cBkP3bM3cPRBCl6uqNzGlf4zlur3cCtuSU7vEpr90ZKuW4EfTbg5jC
XY+WZXuZrxNtk/DC+ona0bTMMtTQ4csTdWXs2jPI42ZAMJUc+1tAit5Ei4QV
Iunz99YIZhpnlzf1CHHN2XXIeMFbTO5LyaQqE+xeYdou1YX53NEVJnNf9D+T
D3mWGLzrKdUOmBra6WGNJ2gMNz+nRSbMDo1Fx2dSm/K0JYvR/iTODcUIiJDn
peASwmfwVnGfF1iIU8tb2S9TrwPu1/UXTL6mv6BW2usWR+gRKOKCrI746Vpt
FrtLtYK2+v+ZSkiYmiS0DxM5lVwCaGN+oUfpaO+q55u4SlQclguXVHzvEOu9
HndWU+IZPR3xXGqbwC03aD4CwkujFXLBFmi+AWNx2QMBTcprKtA3oT4k4wiG
RpL9F/V3D+x/vytNeIGkPyKZdOiZfzSCprZMZK+U/UG7AvaXZSkskoLMf3G0
sl2L7l77r8U3bH2p6wNVd+StWa1hcFz0XEnRR63jR7gKWY+j0q+JpQgIrdhd
ngMHyA6xmcrNidHEJW8ol8sEVFC3B4+jMK+i095W5UWkMS4eTuoXXVAJNhak
oRgbFbDcDh2JlPkmBPWyRZkTTKO7MiiFMetLixqA/a6Xt5Q17rCT+omex5mN
+5RyK+D6gZNtj+b5UmOOMrPn1bKHxSvEy3YUeUVKlO2uAQDhJOnnV+LWzOTC
n5DWSq+DCYvRSu9TtopFl/V1TEwbt1F1n98DN7rVr61Z8mv8X/CdbFpVETEr
I6qMcsq+ddtGbtILFn6Ft92vxcrvEWsIGXtX2mPh1HEHNA7pr22TBrT6BQ9S
FaRdsQ0h04VRHCCJLH5Hh5zaahGh2yka21XAN02+3p1NTPPTs1EDGPjPMKg2
AQX3v5tAgIspjSaOsl/Vi93m7STcCuJnsV+PBsNaiRhzSIETergE+rg+Vtki
YZK7Mu5c8Q1C3tK21MPEeBNvh+mAd7Tg+rLfaFCnaTb0tvCqwdVr+wEY8Psi
p8Or3HGQ7aWSu3x1X5bLsGcdLADX5JAcPHpqdR2n8ttQlTFwHao/z75+tjQl
wnvSjnxd6NLL7kxtEo0hjTSWnKWM0zcMW7yfsXfTUxkXQQ2BGmBsL7ZDgdkp
1SZm0yMcQtqlS9iVIsojO9gTCjzgkMM1SWY8P7jJ/Mf84/I2IfPMCNRZYGcl
U2i9W+Vizus59MAD6Zdele2rJ7ht99siuimyBSGNUoHTtiPLCjx84aQJO+8a
r7kfaWu3DgCRYMr/1THOi2eIVdpYFzd7MpghqdoKVeHyvHf5kXCW5+VLAega
2RUDEaws+z4z8ZnDbq28aFZGBL1pej6G+/6Njpp48xFZaIEMTyodwtXe+ETt
0fIb5EVoLdRaxvtahDJbcpBck2ahhvruiqc2WJr57oYiZT+22BOXClrZmVF2
eNBC3dpzPlmsfaZ5Ew+IfwxdQxSGtXq/17g5xtov6GYUzLCujACBqOX68LMW
/Dp/faGlTMk/3DC8T7RSWkT0mAMT/HlZvpNLylQm8adFDjsgDzsdfGet/fPL
fmswk6x13BtYD6t64ozrgjB0b5IzJ0yiGmyFHqGdOemJ3AhmxI4uEESXge/j
oxG7g+3SCCj6keO84zD8vYzgIx4VmJnz3WQ9w/O7o/EGei5nFQivswnGo4Ra
E1MZ74BVIzasOxCkSD1F76i6DSRMS665zmJqz2FIS0GIfQF0KbHkSiRv8mCg
92FG4kGDYLJxQhqBsfp1QnGNGPO+Dzpz7HuYdU7+rZSddljqk+LSmwk5xFLb
gdx4VxBF0k2VOguGvUzCbTcg7vslh+4acvsSlbZtsH/eT2bwjNOzsFzmaeFo
X0wNL7+0Pf6DtARvJ8qGT0snLOZFESuSTIyd7rr91yvMMZadniYMMmGHiIHv
Pfu+7UQQJqpwZm9+rWJDE3tPTYRZ/e8M8IS4UYV1QcGbeXmS2iTqCzR4YfRt
oyXvSWVVffqapECV6fbMi6QQXeYW7lA3zPDfhg7uukjuaZCbOjSWF7zUIKeZ
QIllT8k3QqOQWdu/ZTSdC7WgXRYSICdIqwYqvNPugfxN/vHLqHdiL2+E0AyA
OC5uJ3dHM1IcHjHef932sKHXNRLxNPWA9m91r/BiJvR6JvGNipQccrPndyMM
CRd/eJh/H8d9GXIyXPU9k6AWK+GYHnIm2qB507ep+/ZQMYKBFyXkQBg6CMFX
ku+Zvs6NGXoBgU5RUIz8WLclr9+XuDVxOtcPXlbs9yNF6oV1Em+OB8CyXPHb
xtE8qugcLlJHpwu+KVlfhpji9c766pVc3Zv58yplsT16zAPqTyNGfjRyewjs
40UVwo0HLNdKA8EyXQqUZxV7Oq61c2pOq1ZPKgFNJkQkY7uKC3kBszhaEMrl
IIgcF493jrx0vx/ORl5f6GYceKUh6OPnESNS3jjHlgLw2XbAJQ8wvz4Qpbou
hPuxlp0Klo98LbRU+YLh3PK7VW5IUQsF3XW4Mh2LZPjXg+t5ZM7t9cRX35jS
RzX8lgxzKg45T/3vqCklnIgL61OJ/DKQ7dEWdzRwNoqFWpaJI7l+MNRbNWXe
lZZKC5VkOFqn1E6JoNk00ifRElR/V69SNsm3RZkk6KomonUEsP26OVB3gRhr
WscreN2rwKlnpDTaSPKmqanSWQ0vvu0S1mGxdoEj1MuyBROAQnqJV6Vm0nHb
J3oqe577Rh46Cty/3VR6baveHH7z9GO1S0KiKg+CD4/Y0sDHhEyr9JvXQE7V
BPKWBvX4Tp+fzTedXxKvO4JlW3zVYL65JXMdT1JNnXKxfEgpWLPjNdzBa2aS
tOGUK6rh51WsWBD+J3M8a/9A8nCIGEyDKbsYPvd0imG8nBepgY1WJer3RlwF
mXHjAhvfGvzhozSGUR1zoErtCe17F438GDJc61kZQUjBol63jEGLzIstT4qz
XXS1gEF/ek8u9VHWIHw2rBES0tIX14OXrGh6hPEniOcffXkDX7FQTBbUbwpn
hTIt4MmvpKRWGb1a8+6bbzg6OA35Or7abAWHukfEdPD4FYp+y9tWuWk8jSZ8
coa4i5h8z5meO7N25NDUcy4iqn+JNu/jLyu/rbDgIM0gzQ1MLyoMNc1hmVoh
YqFFS7Swti10FXh0EZxgDEHmQQav1dnBxpZBkYbS+6uPmqfYyW4Cad5G2NeF
/neJaMhpy6VyTOilK8lTSoo19LsA/tULVGaM0+E7gblXvLkVP8APTxAAvQFK
1Vum0QUHZmVOZYxDk/lGzO9HrZWNpTPReZ9kE3TE+YL8k+jvDJat14eoUi19
O98NcVkSeTk9i5y6QNyDFXHCgTx7Bdem/gV7lllA0KKkqnO9U+R94wSHa6vs
KtF3zZ8xbdUQAMXcv1rK1/fXe94g1Mjntqf9fsp1dPf80izPnbgvYdSz9gD5
VRL4TQmOFhEqmXwNsQcyFgX27R6kBWGYmDyJOTEx0HnolmU+xuz4CKm+XMGM
zyLr2aGsdafzJ3ZdWuFGlNq7PmLxsMMb3uUDF6Ic1y+iiIbXxeujq/uFL8Le
e0Ijf1+Qoo8M52mVo/DEsab621F7Eqo0FBUqqjWl9xnrWZi5b2Ub2jTlhWLR
O/3KKoccKfrWGwkL+k16iOEKrHjqEOuslzUdjMSxKzt5cCLazHqPrprIPwx+
tvMWU9IkzBRy7hgq1KQJOr8VtlopygiJ4F5inrEsuR9kCreORZrvbjy0fFEm
0Qq9Rizn90wiadBnPfQyBJ+i47+9RDjR5b1q+SUwSjO/eXNZUph9pc2WM9tR
87B84zSUZC2RTzH+CqVWMbJFRyT09F3PEmUkutYndYCL94vcI+76sXUwTCwn
j4ZZotygQRzcf9ZuVKskcMQAAunLq86+qJi757qtekE3XzWS5WdiEotWYKfz
f+nlj4kWzoSsNaRpgxw2eVuv77eNmAKysXOKkzocqOnuaXUqWYdWuER20dZ3
q32HTtmFmFljMGUPZzjD+uvl95j9LVqHk1H8heh1KyWNQ8556WfT4VkMxLIJ
ZCJ/+PPALeU3JlfetlK9t4sZgdC+LWgHuK0ghubVDk0RsJzu/9NUcO4rPmcr
6h+Y3GuYfsdAP/Q6dx9tpTgNi7p3HNuDKLQc1T5QhzkoVDqB3mTMypjJLq6D
Yo+UGPzyn43Pb/v3Vx0cZKkbjVKb+8AyFYqQZRwu9H8XyvBGayJvkQGJgC6I
gal8J60rthzudcKyu2ZtUKUnp8zO+wuBH+4lGh5syfz187ibHjGA8g1LBYOn
vjHaZmj3K0AcVXZdzzMHMhApKYDpC2gQ4xB4UWpEtZcXgyzwVEm/HlGOLl0t
zuH9o96X3vztwLMkwrxvz9pS+Rz0WVLlrW5T8+ZigopFSOhREf62b5UBEPA5
2i7hh9IdyIrqbW+Ad5GHU51LXtH+dtSPGSMwh4AhPJq1RPahOQgNetJUJi0A
viMwpsUck7PveccqYeC/8xsSPoygPaXpsRqi6n4Hs0JTqJ0JIcXJaqIEt8oP
ODDDzepizT3zbrRSxOgaU1L2D3c2915mo+ILBdOjvhpcS8ed34+ZP7mFIQOK
ARPeh3I6JlxJisHQ+N4sG9Z/W7up7dtvIrnw3XJBQhcVTkopkbU3XPrQNsJF
STe4TOF29TkAgzwBjPVQTdro73YakvNAD362h6YlDCroQw+dBc/tkNxWL8dF
Sn3avJAHdCvFcksum7dYIMTNcRaERMCHMszOCkAKNVssYVDH+pTgZ0FOxmi+
p3GLanaqU8YNCeCQFSqmkH5wUQcM1q7NxTiqffZJkynsKokdBk5V9uHznurP
FkOOuv+3aTwDiGpa2wyQ7xirPM6YCgwi1q08ywyJcx+Hcs7KwE7b8AtWGIny
EuhTOCuRgzDOkxhgqMkQT25+3KQ6Lx83/gjrdWJGx2OY9I1voncoA+9KnhD9
40SxwAcyJsMHJ4/3d9oU+1T+7iGfr2eFbujxYNAAAR2RPofpOMc6SV7GR+3g
dAKVwAGGFODT8mDPio4Z/QuVQjMOU7mBA5pofCEPQWOkyYEU49htGqwlFCpb
2mS8G/OnxyiuMiujxQDuEUKUAfhQNNM5T5m4dM3mq8y7sbeBlOFCUrlMOuph
v1Hufh5jwvOWhV55aSaZM7OET8LVRtWTHsjnYe1SkfXrhhlEI0XoPhtwun6y
7WUsQ0X1qc9OenClupkHrpfXYdCpZMsUWxCT3TnnRO49KWHP+jMGt4uVZC1j
c1j4rkiQtM5jvoL0maC+Qgs1qO/u08Eoi8NABB7XQ3j881uprTj+u9KFqsRw
tGegG0dv3/rxjOQ9TDLBdhtkzQNCPqd3DeqpcxcJjmWRh65wT4M78jXe6vvE
DOIoMk5n4sPUIuJL2kTMYMW66S5s9XWaDiJmvShRQuH7A8TtNerLNAdujOnJ
Z75wYB7l8YItoya+5WdRfmF1JuBJ2sltvseBgen763eshK3SvLEL3GRoDfIp
zmxrLzIOmsuQHsJ43WetOthpGun3f/wKIMcxLKpgYwpmPzGAtOqh2wvbaM0E
RHA95q+jXTDsQIE2aQNcle9JlUQXoZXgz1pAd6W8TdsaK8ydcAZ5a2ZPaMob
TikHPO9QfLhASVL6Vqr8i3lRQX/ZtOh8JQ+S+bEvlFgTrco31fvKX5e6oIbA
rQVNlJJvk2gGIZ1H5cczBEgk/vicBLH/3wZkNQ1LP104ncqMQqQ0h6DMYqb0
m1Z8ciTGJVVe+uq0bBhaUDHFmAFQvz5jf5/w60s9p8ZWmVZ2cZQHRf58YSuH
2g8SNLuv3pjZhA62Bv+ZYxu8Yj4PUuJysuvgtewjv+ifgEYcK+Y5UcBKqfJu
pZz3laURJFX/khjvfaj632uiTIx360QbAw4UUPEr/wKMC/mAGATsvdbBPFOg
/JWomGXKh7U2JrHqeGauayWp0sXAUXbrBg56SYQrNlVlUPUBab8mIUtpHgpE
rK/ukgxAdQzQIy3EGaUrcF5qWJkhFMv4CYWYSAPGZqLnLJgaTfdKI9Y0ckaY
+rArHuLMM0e5lapbXgw/Hg2xrxFQD2lm5fjjqukzL9s3Z7l5Yra9Z3vjLQYr
MgIv4Ne5kVLxWjoAFx6mQDL81xDWlBKudXb3d4iGUWsFKjCGeDj2kYzxMMAe
H7cOMKTkjv/709TOTyN1Py/Ul7xXogJLZx2Agnk/dAb2L/F/sLjrUobVhesO
WVJeekqKu+RcS0RK3QrtLNuFScSGeg9gTrfxUKdSdKggu8O3KbYIkyqIx1E0
wjlnyXlf6mvCqSU3FxO3ST7H3I/cqincTdgFayAz340NE1Bc20aGzMUKLSgk
Bso4kkMfcbFB6Cppnv5vyAG3z23+FXJMf48rOABl2w8C9b4/2vxqZLqePRx6
5AGjvWzVtRI5gtSBGfM4GHKhcOmGAGfOf3RW2K1VkL85tf3k0e60xMgUsaoH
w9gXkRjyFSUplBl3AkqUN90XR7EzuOGWVSTFjO86WFeSA5wVoRkR0rRFFB4M
/4aiauycTV2d+xzvDEpEFa31VnamXreKIHYqFdtDe6/f30JGaIu+VV+lX7WP
9zFuff3fn44MvITtFTyzI05xutNq5nPqJQIxkEi1KKjzP08Wsb+uexO+vZmp
Et7F+PPF1YAENbaxpdfkzkXCIVrPDtIDgGyG2FSyiwLIR4odvkQ9e4M/CIws
MvrH6UNfsmTZWA/jGYzD2WlllPt+z+SqbwD8/ey3ZQvtq//0Ete13qLSu/+2
ve3rlhGLdyjwcaC2WnuCg34mUrzwg1bHkvqPSmbGEz040k2tyTJCqgWXxinJ
NkNd6h5rqpZ1OURl05UWpcQ4TMryuPMyEoMER4B5aWlYOPZWbS/El0S2joy9
v/Ru1d6JfTa46r3G2ci4JYWXFxIOaN+mLkaHLsMgfBq4fAsggHEEdicWv0an
ocJvAhGzc2W7V/lkokOspMtp+3OP/VwnhA9u0mr5YY6I/Ybi6osjRKdfwSAv
bE/LmDTU4a8yqbXjuPZUpVrzC+wj5beowRN2jWkPzJdsTRwek1E9Q04XxP+t
wrVvoAnuXV+yHPboB7sDlh1bip/a+jTQ2xQdzNDiS3G3/XwZKZvvUzY6kB31
Y8u70QflxU9dnJdc2c/19p8vwAF68I1+eq3tplDBBk9LiXqQK5a4ynE90IIU
L7x6LBnMfZfye6YoqNkmaAPD0p+OL3G2Zv5/4p0P4zkawhgZ2/UQa+t+01oB
OQ78azCNDyFj2+44JXcKLbX/cHBp1u7nO64h5UxwMjJXOkDIflqB+4/2RmPN
xdxCGJM4i/cXv8j0AakPS4HGYWOVcnn+IGReYt2xvI5GVohRun0sSHt1Bq2W
emtggoBRVDW5FZxxM8xQYUiD9nMOLsu8CG19k/iIqbllAm8cYGxEPTux32y+
ctn6ZmhfCIdv2D8M0pmgHDmQ2HHNkY9YqysxoUzpN8mcZgjhh3j+6512a7tW
me9orcNCFsIPLp6uDIyrBuLv61Rtf1EVl2vECaHjathGYoyb7JHP5xt4IQNs
OQsdrQyOxTZsRHRelz92i3N4oyruibInwcLIKYuJbGHuo1WQUv9jvjMrj7wx
UoLftYWRjOeaV8tKVrx/XaqlEaUns/UEXgk8rtRzCtUk3jAzOrY2hSsjDH2t
8MhX5fEtsvF48Uq1FNJC2635RfbpFcAJIoGS7UWhEpNDQOIfSSDyb8XAZ54v
nYO1Se43dy7ALp99xSs5na1OBaJyPRvL2b85RZRdAX+63RhH+OKR7HCrqmhX
vs3caw1bDOVwGWHqpKnqJ6CdtlC84fe/xc8uFe/OBf3lHEd2j+IAPcZOhGTH
LpSEtPG9a/8K0WgEcIvdT0ljCwZq/mtr/nc3zB7MD+fB4tZQhZqIcVZiwlpr
pPjDHcGXxer9HrrRi64kTvroEwG8rSHNh0cRt3wnEXaso+97Pd3bC3owpyzc
Ik7U/wPrDsTwC7nxLUlvVvth7fC8HZTCoCl+lV23QG4cmnOup2E5y3i3c77C
Uk3+wBqLZ9K2r+LoeTki+GXcAQyV1y796ND7Kkdyyk1TtHyVfQ1KvGweQflo
yezJIF8Q7htntpZuk5+3TkQLV7m/KIiRJU5wWvHiutOA2HI0jqqXyTEE/wt3
XyeiP41+ebSUte7pMJ/3Yc3cnpeQI+WeKy9xwfK57dOZeTW+j356GqTgWwsu
G+vvNJ70HKsu7YpjRY3eBREi5blIPOuqJR5B9i17beFjq0Z6CwtJ2gl9rL0U
dLJQRFeeLjPIVG7jNogJa+yW9CP5R4MFPwnhhDo3QDsEYqdnUAKOvfv0iWCq
jnbPTOwGRxTlBesxplmTfWz09xaQQlBXUC6dsOBRWJwU69LlBV78Lar2nPc4
ynYUddgZqB9gqalz8aL3MPpp5QCwkXzSGaHof8LdV6apWWyDMIBniHd9zjuf
UldChON0ywPAn9my9FLXxo/uTTRK3GrTP0KlnkBrYb/FVGcSEyqTTb4qpTNf
ege8YwmMrAbQK3QeruartHqF22X7rQpXATeDiJSzUhd3UiXN+Z/X/GubdWyG
5gunPqOwwk155QeCzTW+iXeBlf3YZlo6V059e8t/YLXeByIJj72T6CSrRNFv
C6lZ5JrGvNJgTNoFwcuDmdVxybkn+t+JSDfOmvxxF/LsR4TMk/pthXpE3VfN
+wh2tr0cyzYi+h6TKDnYpAeLgAa3gH/8u9zZnkDz3dRuxR9TI+96casubcSP
Y8CTtUrilondn1mE/69FnML+TTtm4w3VX3BTzDPi2O3fa4sOpBMejBNTuSwg
/NX8ejINRFw0iVPuO05jS6vG0E9xxzo3HkBOySEfRpK684dgMnYvneaiUzmE
AurCAOZ4q1Q7Tn/wpT1DDUVDNpBPmFaz4OPc0vzh3mqrYmhAE9AdVNPqn9cy
Vn6D1/1yAJyK91YP5mvB8ro5QECzc+//556QA750CjfFY/wQGU1YhkoR5Ob3
WQJU76akQux4ohZNL+gGRs+HI2MeKzTtJb2YslxO+Co5U0JJ0EnoOUoNt2tC
utmEPpg1tll17IQFVZfrnxZ3bhf2pUPmSUqxETGYaOXymMiWkkgzbckIzQ+P
NVsGpF9Ig6Lgb0jNyIHz/Ktev4GfGxLlLXSlBHCrGLuOLb5IVKpgKOimFBJh
nZ2uUQHAba47iN3AKgt5cTGosqMQqbojDucMnLnxcI6Q0D2L03C+EYT7Cnvv
3Ig4xfQobVbAa1sA6qHw6geDpAhYZUUIlzQYgiqFm27/mz7RwrdsJYug9GIg
yiPU+p5wFp4vPGd8Y/ezAgX01fPyb9gCeiYTRCE+zxVXY29I1XSOdY1vXpGB
CoYhdLNhIg2shTS29pb4eVXww+cmI9Z+8DaE2ade/rZ2Fa+KshihcG1d2Fz5
yCaSv/YuIjG4bwVK93GNabuKQA4F5hf+NPUGMmseOcrMUZRem+jDF5iGcsZ+
4gZyh71rpKUhMMasr44ime7aB4/3U/4iQjI9105tqmCgH6ZxTErRQFB66nhJ
6xvM2rwefSCr56XyHQaUqS+1oEwMbyw5z6fsSu2U3QSI0JwUq5jBUF9mdMmy
B8vkRpCUB951dnwgkYkRAZDaBB27X0Ul4aC/l5Ac2lSd3BXbpiyr0FzuUkJg
3oiXKZZmVGlDeAVcJC7TPekr+fdY3YIimXxl3j8LTQnlusXWXsCCsufd1wYC
H+rU9cRadhKOMj/GaWybTl+kxF86opBaGcWkwcRIOth59js0pUed3OBckgD0
RUye8KMu+eedei3dvyB9HQucrQaULRB4uaaPVft59vWkI4878bP7OjS/vmJf
UNJzhcJCEebPBkv17ZKFgvyyVEEYV3OGOXzoqnyNAK+cqyRV7WP+j8cdBZ2C
iPzNsNeDDahRQ5sJWueDjwy5BQ0yUUgRgPR4o8B6TSo1NKVi3m6wZtO/R0r4
PSK+UM/kbAnpMT6qVAJ8NWIbqhQkarNCjvpZr1x5arPhWfP9TyCUsN4uScwx
KkWngj3vNpzp8rIj1s0HzMr7p0IN5/nfUvedCjtbpNAy+pG/zr0G5C4gfCfh
oMCipp8q66X5IAxK7WWp9gikZXdVnJTyJ6g6QcHn99oHwwVc4C5jIdYyM0Ct
RLzB1MRCWI/VCPXJF34FmM5qBuurD0Y/wZoaZUYrSjUqtWIGO5CD09W9ptar
Q6rbDwLoHnqxv0Pgps67LLGV4FPC7HU9U6mEFITMG061/xiCcZ9MnsuS3W20
GcBTkH4BmplxLjWURWavrIEPB6NzwIiYoN8oGsbmVvHwn6Wt6Rd+WGhftKry
Ui5PeCcyy9Or8FT3/Mb8aZBBe0YH8zFEC3w2YTMEx4Ru9RSaufIQD1QkvDNv
iHtnJKtd7XkHDJX+K5SlpvX8NYWoo2rag+BpbZ97b2XtyJEBYlcGkYy8Bo93
Pbd/hwtlykVG339AWoaE6QnT1GcX4C8XQpsdShoyHLspEORhRjR3avTyirjJ
R8d8tgz61lQoLenqpfYWsr7Eor7QiV9ebuL7lqByIk2PhWHU5pHZjp8g8tzT
7CRAQsCGS36IlA80+huaVkfqZoF3kNVjPvbq5NzZfl6o4GFf9cWS31epl+ow
Tomjrz2fv/JM7K8pWDXLz+Yv0zr4YVKMxUA4/ldmS6tHGEVGy/ViS+rK+SEh
rOA4g8Uy9L1YpV7tNdZP9IVzW5Et4v6g0IliwN78kW/kMY5vMUur8GbsT4ud
nETVl4tJSpQcAZ6iS32Oan8gtV8hun3J+lFlzC9KvmD4poyuWbhqOc/GdwDB
Kkd20YZ9XkDNj2hmdo8kXI/QXBxg5c1DNPvo/5ZVr+bJ5v5F/f8A3mSRXOTv
i1fAQiHwJH77TYS+hRV6BuK0lN210603eNTT1WgXZ2ilUOnjX2MRq0pSqlDy
meiRJvuT68I88+sa+aeEOnMcicp+z68iECCKPj8sJpVg4SMNETEwN2p+OjXT
kN6vQc41eV9v0txVQHIqyBnNz3jK2tWC+l+Nzp9jhgy1JJHC10A9DCNtOD/K
+Mee3zLmm6Xa6s7jBtL2vNr5ePGK9O1XaeYqncIj+46AHkcJD/yNbYethnJ4
w62OTeps8eqQiJfg09wDTr6tlQKZ67T953X6bbgKSRn+UQ4UiVL9trtlmi8s
J7AoBFLqaJsgN8bZnsP1Mv33wmaAqH4SeVVHS0Q8JYEowS67URFwyJpFRfdt
b8uz86pGU3/UUkSdhiBretzjhA16n1Zr6VQW0FDYPQlX8NaCBztnbev8XNMv
ukZ+KDbkOSVXknuLt+721x0BE8B3eaYB/Uhimf9hVWR7To9b+fManVZqZB8S
D2As6DwvrnMvOERLR6goK/CTzlD5VWkesNIo6Cxe1/oFC+DtJ4Larq6mjP5l
ONb9S5dw9wLz/I5L+KBDDICW0bc9G3Sbr34TL/J0cdwOwiwOGa9K4XA3JZnI
uBXB2X4B1itpmDn52xhwZkF0ExydEM4t+TAAlLhi3w1vJvIM5uvFDxnKI3Oz
C4IlX0nRuAPnmlIFnrcphq3AUVii+kZREHfjJGEtKoLalYQHJIKtgA34VA0C
mdMBKjkGDzC/IZxNmUYBQUgbMBsHzARW86ft++yB2dbwZZJPinRxjCH/wut/
V7wuS5uJU77hpMNvaraNcEKsVDcaJ0vEIO3zJ+FZL/SJ7C1ce7YCAHUIOJn5
VWCFzRRfMAAny7qmHZqw/GC10ihgleppj6XsJMaUjpOVHOOpAuN+9qC+aRCW
U8jJKudOkWu7UP8odOjOXA/xk//F5SCCh2qpwhWWOJp+ENjRPLOSCdwikQkW
yGamQE4c0/Eu3bWvNHVJV9itqyblmSh5a3juxczEITphjFDTD9w3ef0wHyaq
CXUx6+TDMVh1kziatnkqcfGBpQSnS/MNAaBytoUuL+CJJtp6aKUi2w8UhEjD
8UWMnORaivWl/xxHebowYGN5WZsU1P0XWp7ODUZC9sQtVFBibzVn9P1KR+dl
2vMgsx8dCSQg/J38zmQV7SpzwFsVR9QolW3rE+WGfBuIxNhnHdNfPtZ7995o
JpT47ukDlAvq4DiRKh7ka8vhKkOoi0Wi6YUcx6LcnIdJAumx/f5xJzal9+/j
ZmGizPE+f6IP/3u1OllHLC+7iiEJu2rZ+7MqZbuxm4AdMNI/jcmIvmTpokZ6
dDvzBApfnOsDgmFeQtX5z7XvwRDo0eGaVBPxVT+xkm1hz9gOHj4LW/NLWPLj
4efuvuLzN8NJMq2LG0/kLGC2Nyc25Iaqiv7uSHIJvcprC3ZL+MaNtnwhInSi
QaRTicMoqYx3ru0pCF+TQyWEpe1tJFDSUOshctsduOLjeMTza9LJnyEeos/c
XDHzOeMXEaNOIeyOAdGI3GogPAgV+mn3Y4Y2Rmvpznp5BkTkRaOPd8qETBF1
oaXm+0ioli2Ycl8HwvSzCuol6U1bcwfWrIN7918doRTU0LPGsNc75pp913gK
jVNP908RM6T2no+qjCPJK+M7CHOOxsvQqNA72yTLipvGLckpT1AO+qixit66
3nIJTWBKOJUXAra11yph2KZDz5cBbIH0yQijhUdT1C91/OS3GOpgs2nG8pJG
4iQ9QklMlUorOjwzNF1lNr3uq6QR8PluGTkIiiTwMZI+wPm04T6G8ZUKWsd9
7/MbvjQZ7yQMyX9ZwLrVULlpj0MPZBWC/T148z54ti4OreuiJ//7pocjDFMr
1OZT4Su1knuViTWfNX7Cc8woMvy5PNnlPnGhx32raTQU5+WxwH5g1kLvPiZq
uZ53buh37w7vI/7Ux14G1AdFjPq8KN+bdma73y+y9cmp6ZDYvmogGYx4BVeC
o/yXLpJxKcTvVJnA+CdUR768QP8dKFEuGR2x/kux4zYTn6DQ/qjexRV1nHQ5
b+6U6DgqFiuo/Qj+w5RXHVVdhVUUtGWOlcXbM3SaTY9/GmaZGHkPvRIS4+Bq
LD6ZUXM3HmdjkDLHbNFx+im8jKT2bdv3oHez5EB49n/i26OI2tmPi79ZacDQ
5rsKLZq1fDG1BNY4h6RhSItMpNYaQB5DBcJADFBv4eMmlP0DmK/cNJr7gCg2
J/vpDmYPCMb3xjIgThCRK8ud9QnopnkNI8CLL4WJVwtcWeiG9hiTyg2Dz6EB
em+MIetDvLRmkp0xKE7sIfxR/H8LB/phK7cAj9zO6OIfCZCpPejjbFYSlqim
ku2MCFhloaEJWKxCT/yM8qgYhQSV3v6mqgZuaJ1plHLIXXt+1+606cwiuJmK
rWc0S9AuEJEj+JbnvRHcei+9YwRqUeHgCtITPmFMK72GjY8fAU9urOee/dEq
fY8XLd58n+dh9R/da8rGn38S1YyMbC7Y5dRVW5MzCVr39v/z8Wv2SY4ISMC/
2c4KI+w30XpWIt6O5UTK0xRu0l94+1FFlnCSXWlqa06JAzknUMDU0xfl+Ujp
4aF4csba3qJlyVNP0oyfrWS7lYO99IyYKGb4JR3gE/Drdoxv1HYDlUaCQhIZ
uKcjoQgC0M4ZTE+HHyayIBpYSTvVW92bvCp3kikdRetwKRA/VzEu6loValKe
4m8h3L9wPdUgvfSi20Dn5zrgbCzaBcJmsultqVssybPGBShJwpNrO+otq8L+
ORdXeyp6b94fT8sHI5F3bc44bqq6xljorbz/Wi1Wi9U3UJ/COJX0itY41TjS
YVQ2X/LMOuOJrjY9rWtwK08qpBryySF3Z4IEz+Lb06OpHK+pw9COrhKQfNHC
ay8VFevG9UIT3Qvj5oAl/4fK8FTW6u4Inul6dTdfWDvSO0fGdR2CMrMPf719
Gyz1IEsCma71Srhk3XWbdgshh4l2ehnU9pCrHwWiU9gFSy4BPkL9CP5kaeKK
ygB8qIt+sb59hAXs2ySNA7MBnuqvkeXxpji/H+BQRxFwE/f1pD6VMjYzFMwF
vkLztqKeG0OImY3uwoHk26BLGwEhTyrM9jXozOTvdWAwk/7RErzPytVMUc64
OrooU6IaqinNrqlU36uSlrHdCeb+cnvFZO2fii2WyGlzp3DXpvdtH6q8uuAO
S9PDDLenYxMKohzyuqTwIpl3yYY6Oo1UAjfyE+2yQ0gfc2kM1soFCqBuIWvc
gO2cupJAsmK3vBEHjLDchuPW57eAJYkNFamOT+F9d7Yhu0byEzG/CunyakLm
Wi/UmbxkFM4Bt9Gew8Vt3Uq13f/NKkh5TKInprDBl6kuHK2CqHENcZ2YCj9t
GdVxm8qDZPaA66GHkwx7yQR6rP7RljMoBgbqLYtZK43hK90kZs0eyGsGksA0
ey6OSr49znU8JLXK0Glhy5yix/qrnd+TxxXNa+wr7CO6Q9NfQ+1nNbiVm4FD
6Pb0C4JhPjVHQnM/elPbo8qAGRKlh0xOobLEEbqfVvMSzothzyiH7WM5EZls
RBoatlBTbTvg5OW6ttbJzUVCpECUxyP+p1XZnRW5+MSxqYLQEaWHZbmJfG9z
3xS1EJcB9YO9N6OdLhCScogSbBmXrw8tFDIyJpI/IsBJ6b4vLdVG2HEZnJIW
Yi3J1xigjWAzeridpBZncuRl75VVw6rzvhIefVlXLDzMcHzZGK5ytB02120+
L7QgDNS+eRZwCeJM3HBqnJa4NDDUjQhPxp6QRo+w//gtSGIirhtw9DZn7o1d
wvFXSGLtWQ70rwo6JymA5K8RiiulWp8IZYNKQeaXkpf/2mHPR4v9iKM8bzhc
q+fQSygYBYkp9ccUvLABd+/nb0gWX9Ny7owhiS+eYVL3QnJZeksPQsqcLpo8
eoQhMomgQUWN5KpfgAUxZe1GDnafIJaCrs7iTNHKJPqV6TdiGDgiPGUW2Q8v
3DCRZ5JEGsWw1Tlxqr2+/EePe1kRTcgmiT40nQS142i8cq6XtoCI43iWmJbw
QmtVCjg8BORnqyRPw/fjAnvv8OF2Vy9AMM6+3bWopMA68x8q/0F+cpbiaHJb
c8rqBnd86PamQ0KdD7WViF/SE+1fEKyCIwPg2QFQVqnUvgpkNzUOk57fqzUI
CQ2RCwQr3irL6S5MPN0zvdXxMGJj9nY/EVIkookrpl1XulGysJGmvwYpZ5Ex
myesb4Rve1kb6SeRTEoZnf2xObm/vsHP0NH4sKi6miXuHyTWa2l/IxHbMAEe
UbDN38c6ygenKTrCEkx6QKWeYtUf1Z+zf52k4/OHhHYalxb/40uRjseCi8ua
nIPqD79Ed0DF6QzVMb+aDS//TpPW139x8tBticALVBryaCUgq19jxd8Jn+Mu
CE6Tu8UUqEMKFO8OLvKRppXDFrbQhAOPKCKD9Gs0+wVe0+bWt3Ij2hu/HBhd
GoxdV4N6r5ScCXFjARJHAIFEEQ908oU+RM/L0jZS7wF9i/2J1JzR8Gh9W03q
kOMZfYHLR8yk9f9U8/uPqAhpsCFytMngvY1kqlCTNfBXntZpZv9deQjCPcmK
4AK267UXgj70lg/duNuXoQu/7YvGU/Uf0+6H3xdV1WwYZfJn/uNord+DmslV
W7VReh4wM/vd7TC/IgPCMba8/gZEjKZ0aFoJfiBl3oWsKqAwXJ/QkFG3Ios+
h2ljz5jePbd1FhveEkFDNinAya9it+MyUX+DgKP5uY6oShi27ORtismUbv4s
rGbW4TpH6qU6+dSRn90RQ3QpKU4WkB9Zid3brdZ5GpPq5PDcxT0L72C7yCLj
8ELG60D4a+K+aSiLUM4RzY/3ZFyQNPOH3vFlsgk12diaARz5eaostw2VILDc
2NcnDgreDtmqMTVygzQZCFRlLhS+UdtmfWBySci5N4mSyBquJQh7/GRdljMU
5GO7ZmOlKEHw8WOhclxYmaOTRyTFXUxcGiBbAT8n1sr5JqwIrHyHRlkBZrPV
QJ21RTBfoR2s7CPY0gNTl2kIO3k82tC119qzBiFT6crmE2Cra0tnvYfMZ0NQ
kL4Zm/rqH1/6uif45BKllI4WXplt0W9dmqstSpLOaLnD+qF7YGVxImjNRuwC
lRaNY3ZvUOHWmRLoJIwxiuy1WrfSi/oXhzJlByl2Eq6zb18hwQ3ItwEiIVBK
A77wmbdbPbX8Vhrnh9X5pz5yK/fKkqNPIfxE9WUQWKFyYxsKrG9BsZF80ID0
cVTo3Vp6gPL/cLRHbQe+3NzygZnQr+R8ZDTbpih3jG7yURca67t0pABSXa+d
HmOm/AdBhQ3qRXdMOAIjYZzxpII3xZfKHB0Hcc7TVbfkdmnbp0fW/Of5sPhs
ErNIou7ym7X2nmgChbfOw4nAc6klC6iMNBy3ghEaaPBRI4k2sgl0bPSs9mTD
VsACqVXNvKygo8ZONUrkBpWunaYjTm+u1Jro7tqz1mCepCbu9aLulp5XG2RB
a6jugXAq5AlOS4vpfwkTJfiK5um+o/KYJmIa+HHDLtahUkv4DB8p2yTdjv0H
WXnaxY3fO/fUQI8S1XJbciWECjDi7LVvh/K+c05L3zTu1y+Ngts9CFgi3cOw
CfaOGeKJHPbEAbN/YpPoJUDlbSytzzx6ZHFHUHnYTCEIB1VE4OF5ZIal1WSF
a3/g6yjL6yWXROpLwhlGJ6fTP0IyJ4A05ZbvJvMJR+MsM/JOBG4/ZK7CfpHy
iqx0fbTglPIKlfK5CLygQbm9Hjs0bXHakGXybhu9c/UUoszVYQC0KS3ilAh7
XHaYHGvo3sZ/laS248vAHNPABVp98YAbRgMdJ8A2FsdNE7QsD7YaUDPbNE63
IAXWrWd+loaruUy5N3jBY7+K5JmQrma86l4hT2FPi2FpMqpupgz8TOJWxzCo
u57hSKQ1y3sa4tR0UZYIBVx87jMajtpuG2ESe59MoKqsk3kbLR1E01+9eX8j
NJr2jPHg2YLQ5hkfQY+c4btyOXeNdJJrvgOCqYUo9IgC42H0LTMZyWWyX11q
eb+jdjpUOfO0WAlrNLteca15dd/JdkU/1k5pAKLshynTB1i3QhwQSgj17xbh
OBfUo6vZFSJ7bSfum6RVypgC7L7w+0F4O/imLzzDDQV5UsoxabzpKa39sj4x
M1cUp509tBo1gs8Exms5nPEsnqcARGs8OLpmpg7xzsjdPFSXSsOQHiusXtZb
zINJ86Xk79Nm2b4no4uixQJI7oZ7KeSCbl0OxAhJG9kGEc6FbbY1HbVgRvQb
fQRtWuYV4UsKFSX0McAd0V6UueRyq0veAxcFSCKrZjE1mjUW9vO9ZM8FVG+g
zlOYGoOvudTWvnCv7eLerbqfKxoxgitr/LlwFbTWRfmmQFuwGVuMQAMJawno
uGWnk3UVaYSJKFF99ZRerpsIJ1XEkYDJMOK3SR8jA1JjF9rA5wbk2u+3edGd
qOW+59LNJMXA+0wVopcEdi6cy/H15KJHBAXY7f9TCPETYRG75qdEWfdCRa0T
XJv8ZOa2ovK2iK7x/KK3ScAcp4n0piKrVM1mbUFIs2F4+eNhmp4YYY7LNUKT
nrtBktjuDiz0NbBFKIy4p65by9KyenKl/xDi4GqYrlYcz3fp3ZV0L9gCb8Bm
DFwj9AVtiMlggib8u7oZx64sGrX6ArwZwbHu2qz/zvvjveb+3C+hYpMe14mX
Dwi8VZ+gJE7WfJH1tpEjqTcaXObF+C3HSgLrQhXM3DHV5UJJ8tgBiX9Mg5xG
9PpG7JdsGdALEV4OlUnITHyn3ocYPg7XBvv1Rp/SU/T4V9LdyMdgGK6+oohx
8W/mJa4NSGNZJor5r4jo6jOm6sN6xE2P28eRuZkbOaBWt95TROy2rnTGraZ4
rO7hmy/kdbhQn6U9xBXjD2A63C9BBEbjXHs6ExzQCoAj03AxuT+hTaYzUatd
l08f5Jp+qkTFAOYjXEnf4oDdv66IOyivhA8LKo0FAqKpJCQpk/pvONWGpqph
nIS1Vv+Is9X3r2GwWYp3TSZ/pD+6woY5ewZdx7NG5qjzIQ+G+DRnGStDq+rm
n6LFUUG6X0NvuQ5bIiDJsHeEnKE1E660DsijgYjjSzlPQm/W41vcZlNhcQGE
4+D+/erNHNYHULZ2EgQYUnOWOXfXcagTFBG9cwctKjRl6OSTYA9GVv/GOieq
ZhTrpJMKt0i/f6AW8kltYYHj+WbVC73ghTD+BtUIbQG+/k+B7BwFyq7C5sAG
PDa9np4fLzncX2BKSqDO2ztU6K0/JGMZdqC3u6RSeLuBqmF22NTFjjqkeHPy
OpQ4/rqIqph0IYfmKMhBAbvjB8XvpdBcKqkxHF9SkU+MEf9AHokV7xBOXm1X
RwWYrdjvOPojW2cz2FxVudX7+z8Jy7vMTqG2ymMEGGpc1XEFvWonTJFNZ6Q8
6xcHTFDnPuwomeovqUobRFqm206tR3v+JdHMqTB7Jeo+FN2tctxXdyFxihtE
wyPjI8mvb8A7Jb89mOLW+RzoUouLvJUIR4Qe8lGV66ETdn5HvfjdH/xb9G3p
qO/naoWlp7JCCFvT/DOZH5uonVRWQ3Uvh2sHvZFf+6PgXNVJychvG28V2i+9
7koEL6spyE6EJHLbBhIFyWDbV0e9g9AEaOjy15SAf1acSh5eZBPWr+Md540H
arprlPhrpb3HeY/vRJ3B7Lv7c6+PSiuWX8P9qG/vGau8WPDyq7/KVXWfryzr
84pki6lAVjnsUm50SA4/hCbDRLSAYZPKTWtmqSEMe3/ckhCNfpK0zhIVtv1k
qLxsrCm+N+xdvD9pF8bWOOlBZ1D+4pZJ9r1aJjwEi34+Q+cjDh0ZUBLRiH3R
lMBbtOtBoXKQ58omtzf5qNBHMW3CghUco1iAl59M8Mev02sJz67rcGqreaUw
oQMMhT63LlvylB+weEtx/+ofHItYsLuoOy8ryaoLuofFwIug8sOCIDnPYK9S
22CBMMeN6d2p/PJutSq6sPI97uEBJMtQLfkoUJjVEIPKVGuVY0/Km44hC4yx
fCQnpU630p0PP2CZqOhenddRxGEX1DxerF78xdzM/WauqtNH+3nmABQu4t3K
g3g2+ATujDfnHctTiKBA9sieZvO8B9HYDBtfFaifWvbmpLLxa2BPHyIywVLA
Uccm9tHmCphJYkzjn3qkXe9aOz1OH2LUbCaVg2oE4RZd8zHq+OZA//pdHTdc
wxDzLfYF7A/18TxXTYxMxZDAHM3o5Wv083TznB2ygI7xnGuIUUItwEcLm+M4
JKJAhTz354kkgpHJ+NlEas9V+rljfMHHTW7cB1BV+hsf7XBrzpQccdsVhGUo
P8xO7Gpb0jAZU2e4moY6MIai+RtIuxDFrtzi/VzjuDP4/7VWneysBZdl8Ax6
Gxg5l8q0C9Iqfh0lV15nVohWEvjzIS7SA8vSGLF5zC2WramPwfy7U7In6HuN
FEr39+wvhcPvQRt9/cJlkLm9nJTls/cJ+MJoCbB0s2szhugthFLVWxC73jdt
2iIq248oriJ+tHXH7+H8Zj9c+QYDcI8TvMDF8+q5oEoPYQzQ44rURoi7rGja
MFGmzVmO8LoawWG0tjh6wpo6MYl6f+OQwCWEoIlys2sa0HnkO+K0WZ+dup9z
5OL78ZGNaIH+tNCLGuHLri8yN21Qv9Zuv0AADfCquiWZtU2bDwnCOqVeBWfK
EcO7b1ReQkQd6OrQ2VW5j2oJkeXCt3NcwaM0e6CtDaSH7lnMqCk//uXaBnTj
5HKorcQwvAf94+/hUetqJremwAc2Gm4ZqJSC0mVvUGmlJxLIKEQKHHSY1/dl
sFqGzBQRSlwyTZVDw61+NWGCxIJHKQIp1sKf3ghQHSI2IUvfu3jeH6Ao8deO
0XGr2YdFUyKIScMZc33r7eigRUihUgEbYqGRyQy3KNDHvyS8J5OhYNb4IYAg
7yA6DWgrYt8Lhc5gMcc0KGGw1N6TQUvbHNLNPNsMIGTYuKkvCU9w+cZVs7Md
SnHfDFPxjNM2iRHy32rDLuJs1gcbOrdtnm4sSlKtQq7MvgguwXbFFV8fxQro
3ysr/DGxREW2bTxrOyif5dz5dUb0VEVp4RP5Qhb5172XoKfpIHDxXfu6D3Wi
eKUUJTlK+qDj3pCEpVxVtKmTLSSx4ax2A0tSKQCmv1JJlR5RUL2Kq1h3zEGI
pvRherscXCxspbL2E0RfCp3rtq3HZXD3fn7fufkiz2gMB0wyeSe0edvdB6WQ
txXlCi01SJXkgspElIypc7n8dfC6/gxMl3jS7EQxJ/JmOxVvcMaFOKAWue4F
SrYPUXXKed6EuvO4ARtKRZQZu9i7qVV+TuZ7u3EfoJ+DAQh/lvV3MYE91PLw
27aQTEH9VnGjKvQaVBoRKoJkwkK+cla8ZaK+4gvuw6kUzPUA9KeVGYWKHvoW
qnfboL0oijXWZjE1y1p5vV5vR6wnpHZieAAATBVLXlIhL7IgsYsl1Ln4fkpd
9BrwwMK5b22XuUaYR4bEJbnht4iuyFYNj+3ZrMhhaETljPP3slhBSMbfkLDy
1DfWJf3VutNN72BQcKoq29tH9pvrLvoSyJ1deB6B71R39YsZno+14rhIdUg5
wYbZTj2Li31GdIOBwvXG+8e+jlgpsReC++tLwF3LmD3jqUVuUwZ0Lsza3VDi
+0DUqfb10JbEFX+snCIZIC/1oEgnq0GtecXOe81uC1dSBog13svqXMhqKrr+
rXDeO0iVYw43IbarHU+/LZ3cbyVVXD6m51URJ+ZNNIRATqs15R3OIl5NwH2A
Jg8lCmioD8OsMINousM7yQ/yEVgHefBJgFA1O6x5ROPKQ7Xf2adBJ6knbNSS
jlvCMLrhKs2eOvmQaclnX4CT+ODZZVM6s3qYNnwZXzfsJVZaI3Z7U/lRDl7G
9LP7ECA2HQHaujPrV0eg1qlpCCktVLRmhgjvzdCxaio4dfX8InDed8jlCWWV
b3WhvYMovtASprZPTajrB37tzhAXGU3aBAylhoLLkw96PFo/KxUXzxnBfLgy
HPbAlgpdSd3gPII7CvUIs5p6zwDUa9UmIA4o4im/4Rfn9onL+wCPC86Kq36E
6sir+ilcg7B58UjlNXVFkoKfOF5IraMvPdSIvy+aB1K7h3/Lw9W6aepTTPo7
5ergTUDVf7RN8WWKd+4QpJnx/HXph+bNA64yDKY6lmLZonbUskEDE7ygHc7i
gYQa6Bsoou+W614Tuorqfk4VQnuEw8ZyaZaxvZU22OBmxCLt0ikhjmOpUJlV
4o/C7Lq2OzVc+mYCDAzXdIBt91AAPXttTJ0AZNBYz4f1Psm+tTvWNrkivtXV
rBrfW6GnfOXCk0qCcUIEVVBSRXj/QFEaAAc7sEcvEcXAbI+OsadB25GIQ14f
4L79PWtS6Pu16x8qUAwX2sudjUbsv08GFJOF9pL/5/YnLBW/skEAvsDRiA5m
Mt5WNu/5HU6gpnnBQFxpB7meVvEqOopU4YH4JOywxZX0CbLX1gDx1hcSWhmw
b/wvWsJ4epLA8ctjp8B2vtNzAukrrrRMTe/YYuOh0DO3eJQq86WC85uqpE9q
RrzhNLVLq5pAV6Zu7O9dHdmT7GR3Q+Q2LV09gZ2eR50B0X9KjdTquyd9FZbk
pTkap80fI5qosc7xjARLTXQbB66WLPe8NBT7tzkNi0EjkGLqAqa2j1YlnS2B
v9HpLaNM5E3uFrJaFIuKkpSxZdmnz3So2O5SjNZihRTBFxHRVei5nIeWrSrD
rvsle81ipkDNAZSPqfQh22tAkT3I5DJOSs2cPljT7hSuXTBngg6upHD+oNk8
TjTBqGTJ3woa/jvGiM6Bc4V5OnPqfYQ1kXatPmaDw92UVfQ66JeYrgbnYTzD
BT/chqq7o6TwvWFWtTk3Q9x0ezr0YFTP9OeJNNu5vBnL1AvX3YCeaO8CPGG5
aDiqOYEkdtd6OH/N7cocITQVkJTC3kgMiGqZrY8m8iAuTxuvuO0Pi6H44194
nxoPgF00WnJyG3Qtp+YeCDR4TLxMsrWVgtIOzs1b0vyydtbc3WTabG24uVE8
0XPB3FKMth6jb49vMAVrDOlBK7mM/8xVWLiDLPK0Xn+scaHJd93FaMLPEwZs
+dH51PXeY2vmpJX6rrYPdVmiXSzp8eChvYcduMDBaTZzwlKSdOyIWigwKuCL
kUAopsFuXCnLcFjG3NTKlpJodBblPZKmiaJ/Gy9QDvf4sCAZGAgwOMmjG2ii
NUolnnEYq+dO09aCspScbanPXhI0HVj5U8woaSgy0ewNpfdcby7SGSQKUFci
AkoPZmH0S6oW/AFqDh1LNG1lAtx6KJPGRULLXXQQ/WZXBBVC+b0gWFhPhq1C
XUuyUH9/8lxSUhr5rTuhoI4XdpPlHdHFNDWwLVsypn9mr+/csxfrEJpdY3fr
KHA+EB/XBbsVoT447I3Yq5tQw4fgcnLOw/2gUug77StraH3ugZHCJ9WFeita
yOZ7ekJhnLrwwXgeY7SXqh9HhilEg1MJrS41Zl3knakvG6TXpi2zkvFC42hp
RVrVQxlOPZrl92iurwupy9Ib26wUsxZ8F9V4I1uQKUVkjbC2txf1NxAw+zH0
kDNz8I+Fgk+ja2MTWolVRwtg0gbe7tSefU8aJ7fvwkBzJCd4hATlivRBUUJk
c+FQJjsih/Qcn1VJuB7ulbwAKcDoO3Fsp4BnK1Wo6qMZ2rOFwDuc7fyppeGZ
LDLH8+EFWoXpR5tEbaPk0BO3c1cnyImRAY2OViERIkVWtK9w63W0XBr+LkFr
U5oV/4ijzssXCf/WFckhuYZ6u8miMA+vEoZRnKwUlhf8+FSATBTiA9Jyun77
VRRskWJ3VKDAZFynhFydaf62EypdNZ3WcVI0oClpMbcbUnTuTB3N3LU1UcJV
/7LsHMT8Bgf2U869otpqMV5JTsE5RyzbsKDJFba03RapacpdS3UGex0KQwCr
i89eUPMBPI672Vhth4UOfjHfWWh3kW9rjC9j6RTDWzwTfgDPa0GziPha9mCB
/Y+6iZXqGYNEHrza4g77NhAY3TmqeOVsCfNlYV2bYMHoL6nzQG4fpQGz8D6Q
U8c5722HuUu3iBB4OZXMJmTPaFkE/nx0umnvQim5VraqPedRAJKJwv88Q+0C
Npv+KVcn27CUtP/UJI+zQ5H9v3OmP7FxYss+XG4UDRZ//5+JEx+EgP1tnhjF
OL7Nc1rPyBM6kIee2EXztxXvr90RLopfj2fMifsTOpAC9BxbF2NsJp+HFSA0
ekJs0pSB+qz9WHHw4z7VLhKOl90bdJYKaq2/lZTlyPMQ9Z8idaSkuZ9jTZlZ
pCOG6iQ7zik/5JmHtIpwpQ+gg/AD/Dfe/l0Xg+VILlZTPoTRbbsmZAFQGFL5
eUWwZnwKjPDdxH1q413zWFo6s8HLuA/qNSOmafbnzR+5EuKdFAPyc8bp4yrI
hprazpHsTY8dAucO4VInALjKh0S3y6A8e2fGCaRH/u+ogyW/X4T8ip78Z7n3
84jBL7wHAdLelxC6Z3Jjw1h3wayPI/d95hVz5e/YQxcsdipO8hpXVJ8cY6pL
2nRHV7MUbcRxybIWbN3+/yClPpiSc9eLc/W7jRDsMb1S4n/Q8+6z/nDyvCUA
T1VQf2Q9nWfJvIrlKX7k6b28HX+mPNf6Qyd6LZmqQwxXo7IUu4K2H57UEDEj
hTLvi3BFmco+P7D/bViIkMk/rJi0YfG+swisAI62Z354vO1vnmPf7ER4EBZY
jSl3fxU82Dtzn2lg8iUHG+sDLwzWEf6xlNykfx6IqkVldlj3wonxZy6iYZeP
PYVLaEJxTE3ZoGOcLVIA4rsiCbPWkKUUPx9UGOwg29DSnnIMbiG8wcCPePA3
wViYYeUY+ysmqZs7R0bPcRPgTmgA+7gKaLM6WBfDD4T4l0SDd7gjlnV901aR
9bZ929eC/feEDTjBwi4psT6a8nRJ2MNLu10sxBsKKI9GrfoV3CqZ5NRWcxcl
c3RKeNRBrglTLt1pAcOUVcf36DA/XG18rbSWoEUs3/LowMAhgqYMpQNXYFNq
Z5HCjO1yoNl7l/s0o85nzDdA90O988iZusj4tfeRm2oYz6tKYFdwgBdkGOlT
CkAWfPCCoxqDEyTMKFD/2SSsZb5wLRcOsVgJb7Ur9gofToEOy5DY7KO+gkpB
2LBy/35StVeTK2V2fzxf3lbU5JMdnkOaysJrkIkw77p1mM4p13Q3B0Ti4WE1
7FdHMFuMs2HplQ87/+uoGGbgfb0SceFBLb6bYEoZJ2LOr7/a7y8xWSFT2mIJ
Ew+/UULJER5UGVOedsHZdYSFFe0LwqQSBN/SytN7DEPNjlF+6KbgZiq/SgcY
4STJMlk2//6T7Yj/InISuSzc11k6hJopZ3rhUcFv5mwcBv6I8oLYEJAwdabM
T5QoP/pWxW9AdJUsDKwR42RVeWpo7n1/eZ/GpZ01OYzQ4kdmC+9v5ShuLeQY
0nDEp+A22kQ1beynkuui5jBEa30jPPHzUeTnyCeptRyaoYqsqveNr9/vzgXI
bHaUSptbD4SAb4Z+WdnrstfD2YqHnXhi30+Bz+Pf1Vhfx4qTgfVCFlRTdfNI
0IOcV7BjEv9Xrtczm0fUfprcNQsDu5R4DXIkP3l6IZf2myBKxMWReG0cdOhg
FwJMedAq8uwRfc8qrazRJLmRf0XGYcFuRdZDVI7feSG8NQ0SYnkqB3ulc/EV
c6JBMS+pGwxbqTOiZaLh2FHdVxDGZpTh9KF7N+ZCsCGHmdsURmP3dtPsiNkw
cpo0VD+gwmctmttCzj/QKJmkK/jJ42nIQctDUeJyOx8x4uNNjeHOANSZdknO
7Srz8vnQgrUj4morPSsWEhuZhorzRouKF5UvZj5PFflCEXmFxOCrjMzMdg0Z
DrpuWIPgVdY0ccs+9AM5kn9qu4Fu7kuUgJNF20bqbsU6YZ+QzbUzkVAi+fFW
lECxc2G9jeKxinEcNS6jVgfmG3OwrZ5dxDweKeUfpjInL5a1S1MYwFWqgI/U
ZLPKjTMu3yRtqa50Bzin9SGNVZdPLroFPkOL04kv6vTJxLI+FgkSHWlc3Nmx
flqHcCfBMYci0sXpkJcbxl/LOCsINBoyWVsF/AdmGm4gef+MFy8rK//wXdV4
yRgyxJCWfZo2zQjlnbgz0AK2Sx2UGmwXmUyAGG5oTLajIkunmJ5mIWZXN+yY
BGhhdaZTBIDiarysoNU8HfbNuOSDdY1vXCWAmio2SHqhFxbrx8jyAoPeSl/R
6N6Mc8waYN2495zVZMfIPOXS2YfjjNh/J4HcWJuOkouUk0IWbrBDxgV0fFsl
ZuJJYxsf6W6oU0fB6ulQ5UlLPCMhk/fSYbOf7+0jQ9DovKZKMILCYdYUjw37
oZMu9F+WPSShSVyXG64XLZ5iESYF2FtdOJ3UKfKBsARgC/nnKWjoQtmGufp0
SyS8L8eSekNktvifZGrsHIW0748EwvhXzOkY5Vav4XWuhQRR8Dcmgxy+HFuG
MyHFMqTgJ8a7+YCuLa4ZxxMC1G+f8T0eijgFz89KwO18fsTnV0iGAbBezNmF
g5W4Piz6r52HQi1HJlPUnDWpBht7gXQz4AAEGo6DYu8VFuSNK7acjYCXQbGt
J9G6SJ654KSuLgoE0MmiDswEgWtmpdRIqjxB86G5KpMZ4tMavR/0q7P4YOp5
CpyaeHNYanj8uTHIKF6XZUcVCRvl6EBB83YhlkCWiI8vpiHWQvrbYAuwQtzj
LwcsAtMXg6Vw0jTb7++EVHxNUL4o9c/Xg0JA3KacIQf/kH6dN6kFSFiIBW0t
R7Qnt7puXLB/78ORDx6Kgc9QZdGsg9UrsIpRUe+gPQl9GD3K1IPBiI+2EfPP
CA1K9GH3EociEZ3EcsfpFM9Ea6HMFdqomQxSErnmMy2kMv4hZK6IlM9fcdTr
OfVPG4w/6VmrOEVQBXTo33CQWj4NONUB8j9RSX/DO+j00e47gXMVr6Q6SsU7
a5OWJYW0+qvEnCbMoN3jQQ6Sz0cFodgQQqC14Ti7lMy3U+R6fUGnmP8U+hde
1YZaP1oy3r89xdI3awx0YkBLnU+EE37oBciZHZLZne8Pqh4ZTxhh+XHjXXrR
Xvqs06A9dyV1G3qsQ676jjtW1s13MOMS687kBqtND3yg4x7HrrXt0/QGLSN1
Ri6F0xJkgGppx1vljqk2a30liaZYzX1ND3Ae58RtSqnoXTA1U4tbBnCm/qYy
k+vLWDN+nlrPiQ2+ZT0ZWZ16NHuJAphcA0Zldm6HOsKYPHPbsprx4kmW7/PR
YQUkDlHHf6Yy2cIzlszoUq24D1NJQQQMo8XDagLeJi3kbn5vrPNQb6Rz/TYj
SR2f7B4mIWIXv8TLauhNUcRJihmFI67s5O1O/ES4rEnMVzT4V4ObZKJRULh2
R7D+lsGEdQT80e5TjUpiR+ax4k7tEBFLViaTCTCokkTvnOywCBURRVaFIZxV
diJ/4VB3wUERzwleasi/OXnCNKKtH7XlCW9iZMQImrQEtnUCD5Wnx9uPNv4U
hRYGbmy5qYMCPr/UfgPEFVwzusOza3fjV83DnGNoxNuk2zqk8X8R5xX8YxpB
sVT3JSv1gta/KQSaP9fTSPvaap9ySLdFRLoV45hSLM5Amg+5S1d76pSTwOOe
Bs1YniVrDBv70JeUzq7dqE7pmnr2z58NGAeDU1FKMonZ9LCU0IGpL6Oecbu5
gG4MjTmOd7/01EN+828vLqDXLuqTRJM4DIRM+cxrjOsry9KgIZevAui0+P8X
d3rYaDOHSQY/WF6ZtE98PfCskwtTmaTG7shRRWUDoFVBo1k38zzIyzzvX38q
6n4L4UpDikYHhJ5U7s61VilvcivByUL7ufJd/rpiRqTC6rYgIvGJq2hCK9nL
32XafMtFPa8FpCWJtDGErnDtAogHQUkbM2DPD7fCOPM1ialSg0A9Yvr5OTrc
Pux914uRicATIPrcd94kf3QhhDKV2PWr7Udv5oYMfJINgDTmb4EluWw0YcRg
LQ0jFpjCreC4NKRcu2CcxMKC0QiXE15+vah0iBz4Pe+dgtMBGuqIH75NfgNW
EhItP+6AygKnHLTuG6+Jt60JFhh+emYRJZqiaQLb3pVpKilC5WKGMLrbDDto
jGeC2TpbLXzYh25HQfsY5xK3QPo7PFi9O9/axgIfm8pYJDQr1dZHYt68aqLE
1vZrdAM/IevEsjOD3Q+xCEBmdLc+Tf9QRa83p6tuHnn+WOBs8dQFKR/ubS2A
6hKOAYt2d8aCfgpXvibHo9ghuo1/g19d/FB+opYByROwj/Vw0VVsWyqt2sFM
XDC4ibNDC8CmnrZxrzsDcF1mrvoQFORLZDG0rMbJxSyWFS7XCSYdLxsd5ePj
Nb8cT1drvdzapmoegHsjBitWETDiVBvGon96B543psAudfw6jUxCFlmHPvwE
JbiHUfHISBN2mIMML4P5XyFXknz5lGU/A3YEow0SYnFYrIsdRAQNDkMHYAhB
t7zE3pNjnC/WAie/C7CBrSEaWHac58WuR3vwB3rCC4P4HOm2KMlZul1U9dqt
bWsZIPA3Zvo0pmRzFgamPrhmngzkZw5DjaD7825o+fR3e04PjObePIGhxnoO
kE2bMmXHh9zG6faIeFMFViGMWDLZt7eNwmQecbwxMbIUTVbIz66oFiL7djsi
JOaSN5Ir1ivxKCvC2azA5MLte57EnOo5xNMRlQtPPEZc7e1oYp6Hy8Dmd6bk
2Skt/OKipptHqa3QEaMxyVKryVvqRrYYPYF11bOutMJXXN/pH+a1j1q0HGY2
NzH9ThPnCXqSXN7xDEoBh97l20jZ7axIqdMEWSn9T4YRvWs5KWFU7RGnNx9L
sJFqxmGKW9hPTjKFvbD8A9eFIyABVdpnru3MkO5JJuCJXjy2ypraiU/wqIvR
I61CftdWwIlVGWoQYDcIeaieE7xtGzVPgbqM/c+jGZVt8H/toxWwhAAe5OO8
zkIFVpCIx+NOwAVRag75BZd0LQnLklzd/Ep7glsubXeSETIbXNsm0sbIOgIr
C1G97wPjoUzfqfcoKZuxmEOOLqIdYTVwiTQwa9ngqC9JytN/Z+nkxGWS2lNe
Wzh+laAh/DtAPseTTL6U+knj9ZcKUe++J8x7YMu1VfXC211Vzoq04ycIgrYn
7jsdcYcd0yR4ZMWYPIOmScKhfyECHVD++dnPBWPbVJ+hdNvJe7+KMi9DI/1U
2CzFqmeYASpKI6kvV61i6aiaHYqxGL6RFuu5Th9HA/P8aupa+tajrCRW9lWr
UGOsfii6pJJt9RsSu/u9emAe2psDIEW2oDJIfpu8hqtDrgn3LTlgJalfDwFY
hPrHRuNHBf9DEyXc6ammO+ANbBOzNgWVMhTm8saotb0nZUKIor2OkzsVUnki
JLZRkQ50gcHWxTdiHt8Fu4Tb5yHJIHorz/FORrdaoVfpdwdU6tw2A+/IXRP1
tLQCm6qpBtvAqEfjAjxbalImA05Hpuppn1jC+AVyTy3cfWFjTCVBRV71zUVl
y4g5YMoh0lNpNUffJNavmrKZa4ICzTnMyKzRSUfZAFJ0Hdk5tgrnn9tlzK8J
9JgG5pJajdYSxQFLHANW8rqMbTsH1q3ETQZuddolQ4tHljJO0VI1UBdSyuWg
7F7YO2NA07Z3sEzSW3EOpHIu5yPUMV+Rn/bT8RPhkruDrGk43lpg6nLOUziy
r7FlgruRCIWRws1C4BTnhsSYcDngzT+ovD9jjk4qNMx3kUAdWoE3BJcEZ95l
blMY3ELgFWB5bPkNc7su7HOS8OQ/OeAGP0qrTrBckIfoi3YDpEtozkzTdz5B
Zso3gBwL43Gr3oD5/TcDf8DfHiwbi6Uh3zdm1+PffJndrALkYkfxsPDSmvia
OFlvhUCfaVYtjgYb5gHM87CJYKrErJw7WIlXY1Oj9Ei7OUigvIaEZdCZ3oW7
rkWvfRKBTioto+KrZH0mNziSsJ6UXWMFpt0xF8MSTEj/f/kmTFvjzQRdm5MX
8an4EkuNKCAkO1DZSPOlJEuSVlVce8hIBnJKj0cWMLUVJY0FX3zxtINcPfsX
k6ENLHiLPF2cl4woLXhjS2wA12AHGPk59Tr2cEthZ2EJeqvSR3uVAZ6a0+DH
UeLy9thTngGhE82OE0xqIn7k2Y2V++eS/9bNdDZxrJ0Dypz89PQlmPbJEY2D
lhMuyYKY3+Okss68nOqr23fUFUammpY/YjEyFHuXsW1q20j5MN0C1gCEEZjU
nKlmzzIe4jPQvJoz6Lvj0T1NERE4woNpnzEB5C3TLuq5pGEre+BrL4TJdeKW
WuDi9vSD/irmLo5FGxMF2sqhJYbqVP+GD3Q1GheeBIW6ckdUa+To5bBEIhA6
AITKnF6VVoUyoxMNS2DzAlQz1HVCat8XL/d958xdfb6DYtgYHIzrTlZ5qI6G
Ju9VNn5o0CrgQm9EJRHKS0QXYELrb/uiuieWoY6DnrI7b+HVDrylJ6lOBQJV
4Soyv5nKWHq0cFlVDRJSUjZkqGGvvTiXXPr9lX8IjGpRdfGNb5N2XFCHZaxy
V+td5tOiP6OhpE25yk3Na5WP6k4vnRHZZVzfPwCFGDnw3xp59ohqKLuYu3Wu
qugULof9Nma46QBXki6RfxeQbjPrbSAzsoexe3Ciy16sad6DWkX9vvrG0342
DBmYmAGYqvg8mDELbtxZZOAKd3B0BGw4lxpg6q7jvjYQWQUAfqR4OAlYfvRD
TTX4ERQZ3GWb9FK5fQWGbv1JX39Eds1NuzxYJ7z8Rgp01EhfPmOImTxi9t7K
atl9C1GyqYz8B03kb1sFZsZnWSUdkOljspWVOGMCGgWPidn41G2ad3gYzT+M
Qf2zxToO5LzWkMthj6tTLZenEwxjn5Hks1esRMWpyHKs2fO5kpjTIfVdQQg1
lWyrAv4Z6B8wCDTuhSVC/hl5eWaDRm5G9BaXX+eoeQzROGcuHiC9t8rRNk7v
iNLAuG3tFBrQ/ZiWbMpEXd/U7HzSueXCIsQcbQBGUzaNkg/Hx7CXsQ3+bRD9
1AuJIcsdu60VyAZAAlF0QGviJ0bAwxtc16ziT2wM+EARi+a6jgWspiLMaba/
upgNpvMZLu7y3AXH8ew6qHPz42lCh4XlueeVb7r2sl+0ERS2OxkNONXS0noi
pdbi1R4FtnyPVke0I3HHbKQuEcU0v05WOE4NBgi5ZnBV+5bGuQswspAmKVeE
DK1vWTQxBrrKRfszc0Usbb1Z8bCWewGM1pP7JoBWjXHNsY6v9iRhk/Vj1yx9
rSycJ3dm9E2ncfxE8D4+oEcZt/L69Zg34SR0HvQ9AJBt8ULuPOFrZ7DNz/LF
0WNe7BYi11FaeUfwd/LO+e1lsO3T2d75xM+kzrmi/iepoL9f6yTe63hpIMgR
MLunypqVEAAu78+/oydp1tDWA2JrV/Q7FI4TkEAesBC41w4XsEe3tp4bxXum
V8RIqKdooOAN/LVWzrHjRtdmW8IHFZlhOOZzW2RDUxxsuHTmSfky2NvLRpyd
SZYPY9whN3GlhIS4wDmcOVUXv6ZHYPsFjzgycKqMsRLK+qMAbHrqk3gYH8e2
6vOeAW7WardT7DeHNMmwnpkONMeGbaHV9uOq++kOVU5XYcsNRzKowh6AsrTJ
fh+cRI9A/ptw/vY8vPGjkK1536Jvt/GQsnDwIQIPS2h+kHUQ7nBbijsobazK
NBERS94OZbgB/4PhuzHDv5KSNrJPHy0v7+8AOTKBTbvdCBywBAQMD7Re2ipT
zilUpTULSse16wR6HibGwccj2d4tbSABC1QKWn4HCZ6F2uVTVSFXlhP1Ht9o
AYlWCCMQF7vRTyvxhsnA3vilMA+rFTZktkK7bEyTgwfUcWI9I6sWo1AFBda9
3NFi0h/Lv1TQnV2FSDeRliFbG/6t3KoVJ7RnDZsz8FDMgvLqrBrq+01RX7ST
E2DBojMj9YXXH9J+WmEvdwK3+IganJhtbK0wVpLA9vGisVErPatnh23ir8Dp
XHCTrqppVpOJNx3pKBNdP2tCp+vJckSyY8DDlCCdahH6sGk/VoPp2ikw8mch
D6zNmkyRXzlaSIlqKRD1lY3bzeelmHpaKnpk3TZsBZerqBuXgazV22f2AtYh
Lkc73qGI3VJmwvJ3JMUFB+j3BVrBplqy2wTeoOUjpAFVYhsob1jTVaFY5oYs
3k0UIc8trv1E33OxS+2k6gPW2jypse/dLBW3Ls+UK399/0JrHGBMD+AK02r5
BhT4bOYAqcNEx3r1yKg6pnf1JnL8EEPMRkSANo5mqlA1S5HBhbef/JwFock2
KiAa5FGWl1c2Lx6Bd3Fnp7GIWlyP7buPHxEGIYpqAKyIjFj+3F6sV5A0Seo2
blEdTMKy2e9e5EmBrgek80LGxJqWIkAF3aeOjoAEyeDOoT1a8R0xaoEGP/Bu
on1gLiTP9isUAgH/LxeXtxF0BbPJwDXsbk/yp99yOtNP4rMX1ohKMju+fJyP
JVSJwAGZH72njbAvAsaLVz9lztsMWdCepvW1Lvv7zQx/hrmIpoWb46dbsLFE
m0bUdoNOGYV2FpFjgVBOv7uDIevJa3t7yM8REF58TigF527yNzRiBnJz37ZL
TiwUpCysObSQ51ENnA/4HifSukEDLjSjBGMvXrHr28p0DpmWouCcmpuE/Iv2
JUogqXYKYqhydwYg3GvYEtMRzGa3LaENl5hmZRyQ7n2YjiTkUTFG5UhE5MNq
uOXG6GBqSQPZ8poC6wNLEJaI1ywsc/NgaN1qFmZYJgPpSg9/UBdFlxg4xX17
gARqeCwMZaXr1iEuj8dbTeDlfGhDhih+g0dMeMi3bixzo3ZPqXxv+daPynjq
6me0G/9zs1ycEgOW9DD7zMb4iqUClqkzL5/7d+4BEQykqkiXWCncCP4hMAJD
6gEuomlDnaYGNl7dqWXDF9aZOszsOhtRf0RZJVQJmkhdKJIj1yiQ02n6lyGu
sfVzd9wyReTTPYrNKxGpmh4+69UeRKSEnpo3LnEUnPVFYitHtoa8+8XVSLVh
IxaWEXVFeo7qlc5ocoO7eSfRfS242SPW3zwws3XBS5O91N3AnKVmq4jGaDAo
QUnYrgbRNsUACk8/oxjbdvYY1fL6nDpWzfvbzc/w50OAnZO/C+hawMC3oijT
3iQyuMCi6EBgjkwxpchbhyEztwoih/+c04XH68DiIGJyccixAiD7X5B63t+V
1aA55oLeddwCuwrLnJXjkBb8RrUneea4c8yLVtAhbyOy5NV/7tvxVTPQ7Zao
h0l70TXIY8tcpKU4nmxeqZqRxfVPQupEfSC5li3F4L1H2yjFB9XLe9DFX3lz
0Taxjv7XuRGz3ncT+YDS4TRx+dG54qcaZzgtKY4yk5tcZ83UaKONGvDihxKX
bS+awlL5zV2u2s2qdE0dBn//0Ypcy4nPiEbJbXHNWAOCxwn4+Fg+n6mb6zLu
9v/9RWX8QOn339tSB6NCXQYE4lFMicUpg2XOES9NN9sdW1WRWaD8dStzIa1S
iU1tYCfGIG9jOpF/QAxvCUwTx/UXV7zAJgu7+nbVoFpdKJC+Lu8PO0+hX+J5
qP8/ozVIefZ8oLm/2MqipcS8YEjxNf00FQaKqNqCBWHy04s9DWpGhGsDHZpC
54O3UkODcZIa0PnfTzMgsCRmmmIzutIRoK4xN+bTLgszNzrC89GyBwXLMNeY
NdHCPVKEtHjaQQ/0HFO6jzSW4XIVtvqiNpd/vG5tFCqKHvKO4wZPGMNUkA4k
9xADcj90zQMEYQRDt9hUVwMBiH6GD8C7+yj28ULyRslAQrWkPUw8m1LVduq4
VnS07McjRRW73jZx7y/Eldea1/saHbqBKyqJ45rSCHDN40UBRbd6vBiTnzqK
4olo/chRYLjA6hc4f7r7M8yb8KUf6+XzzZJSBerUllhu2jEYyP04XdL+/IxK
rToyJFv8FlafcR1K0hFUT8iRTfP6zA1FpV5tXI9F3d3gDkDMNZiPYD2mQkBA
FowqCX72r0I3FPd30A0ItMipv2lNgFMFW7j4BgxSUI6XoMF7SXNVl630tUce
fE3z5A2amlzPjBHMD9HuChnmn91Njon+amlxUHK3ei+GzUhvL5ievaBopYuR
lD57vArmH6/qbVoofZamwf9YNo4uZECkRYROOGK0o3SN2uEpJXeiGgmhe6gg
w3seojzHUmMRo9aqL+tllWYhATn1zzwXndxragRrmFC8kWcQpYOKU0MSotxV
52nZyyKM67AS/ndz8+jWFUt44M9wICvdgmveVwSvTiqe2xk1weZZor9QMR5o
8BRge1v7a8xbdy9D2bmXCkofalWkrL45TaSUiUYJL47U8P2hVw5gs+om15kD
pMhvOUcy+7BFbqS5WXGbztbF44t+551t2CCXt2AukPSPv+BEWhMrlIPIgtXo
tfc1eTWydFYT+sUp17oj83YNr/bt7KmzVFHOI2EZp1kG6H7NQXLK2T8DqJ2m
8AQepxErMjkUcR03HY8yn/ckMpdTooATxKGfOBq7/b1LPXEhpV7SK3+yBLuI
KUqYa+mBZs+E6+NLIqTDZWkcgqnJo4eSB2RTPd6baZaOgAxLLrgjHr7VUJVY
C2A7h5CtSIgkrCVypPzJDdjka/Qt5suTyobWjuBr9feD5eSY31JFaINF/a++
PNmFw6ZPtfHvVtT4GTdaH1vipMjQo3JnJvz/P3uleTBrJ0FF7Ug1zzM1ctWk
/+WL233SDtSafYP5nlUi5qoqe9qwkA3Fi5NB0b4V+WYys1CAOdf9c7ZbAKqQ
uGYFlPTAhIW8rIrHVqvR+esuK4O2tgtuJ3ZtP6b0GNsu/NOopYh/jsuu3Xbl
+g+/Vq+HUnprEE7cY/2VlOEhYaPox0HsKQYaihkkFdO0fN32h6/VwOifHQTG
LPhSjb+mjVuuvBOl8XJiS+lYeENlJpofE+Md3GYgrJ0AgSLry2wwdfB7xuwb
DZ49zrx1TcwLbNQ4LZvS7KpHnd9OUU4hQUAR+Q3RGoXhYtRajK7qJrUq9+fV
f85hXe1uNaoI2aaD2ohgMCF6cIHi5+2zs09N6eKVGhbl1xjUfGqCi9MLSoZZ
zOA/edOaDkj2c2jaIkxD1wIRNqJZ/Ufx7ZQplo5npZMZNoDfpz8S1QslALk5
lXja7SMHCiQ7h2U6TkyUIBZcBq6TWAuWES1JFAZoizQfx4M3vrKV/5o7TmkB
BAiGRFo4sW1ACBPGnTCZzrQ8iSBYRBkxvW8FDve3di6lbJchqrvw9U4md52E
KHiskCxOirXsK2RNiAE7dKMPaUHcnCXcPlDi6V1eYcd9ADai085eZhnF+WIS
XBAABCB+RBGkTk0rOX1rb1o/GgPaR8p4ZZpp5vFzZx3bW+ffWkT65ZdoPtuA
zbaG4r7VGNgzQOGZ7hGCvgEybvYNxTZOP8DvU/KtiHo9TnwIK63m/C67qaZV
ql+gyBzYo+zi4HbMb3lYmoaFud2xoyz4NykR7EkAFssXhLhcFUkOsueRBhyk
948UwFOTQAMklNWBgQPqtk1vtLNsJNgq1lIqfusc/MKnItrOy5c2WUlolpVA
e+x+Sltc/V3W1z5yQJE4inHL1I3pX9e2xRYFCNs5qWVtJP1Sba5ncTPSLI8n
ODPYYRsWYz3Rv0ifKut2nCZCgz/BFvhKL3mvEE0Y5Veul3L3SKYq4BkpTaGB
Ht/XE51bhxbNjw3vOp/ueJcc441XTxFtgIPCw3ShGt6B+xD4yquk3cOYaeE/
SzpEx7Lwp+DZTk0stWnEC2YI+dPGpkD60mSrxwT5eklyxta3P6e2e7+EOKkz
wsk1kN+z5YLOQ85TeetWqG2RYlk2NNm1lehVqeQZ25KQbV3XUwonF+PELKKs
klEp3F5Yl91YmISvSuQrzsCto2JNJQaXmPZ5JxjOpMP8/HOsafXZ3DG/m0GK
F/CC9sOC0n/FoMkv04QibffMEj9k562Lk9UzALYeNA5MdqMxFgwmI7H/3PHT
KVSGVLi8G2cZKWYIP3FcB0C7GoovfZiPtj7SejFyHuKR+oYcHQlFUKoA4UtB
xddrrd6Tsf5nbLk1E+jCDnHA4sRVZE01fYdteX1Qfo/xKqrs5Js4nlXLJahQ
mEPwDrENiwSW0411yEMPyI5kdxLpmeMSIp28xPWp4HRg6mDENUt2D5ktZcjF
Fc/UZbI6ONVI/0VG+J6gqplvI4cZdzEqOI9db+lysJoGHok3LZfxDx7+GPw/
wJGspswQLm5UQ0RIR1japSXoTxPoLH5tEQsZJlrW0S4k4nG/+ehk2xkylFP1
CknQFW14CeTzvOxQVmXGGD7rf/emINfEj4h2FUObYwrBkeMEC0d9lp+nhsvS
O42jpWo+mqH9AYpYBI5nhvgVLS1qnBFDrC355nzvA3zMkJhvRwuPBIZo8QVX
iQvle/ETVABavUqoorkHkB7P/5WGHirXGueMnTiNNMwQnSlXzNyZ2oQRpNt9
Z9ehrsbveJ38Tz7UcxJXpm2gQ5mhOH7gSwzYxrz2JwNzFPtO5bv/rIEdJo2Y
K6m4LtQ71P8aaUtsZ1H2sBAfTnxAyaG0XGoYSHLHpgeEzCry62fooMW9pL2Q
qNEuXF6EItnyVnJqaOjMdID1yd2X5owgBtTlhIJ+KcKh+wxt69NzrDn+bNPD
mhDHjvJt7S0iRxK6YlUGV7Jt56gjOQkYF2VsxFH+lg5YMpOXBP/Dk3y6o8/a
VnhmisT+uyu1bcYd6KStFAPuDaR+zL40ElAhPgF88IdMlYaNcAA1qEAL0mVj
lMp6tF+NfuX3FHShh29/375IRlIt9/vQ3wxLd/MB/i07eVL1hQ4BK8FlVH2Q
dxTqjfSngUxdowa2DOFJoga4eoNTD5IelJihiffOzTy5OEgqmiuqCrsx0y+U
BBsWGqyIkKXQHD6O941JI2+LBgvgMP9kpfkw/RcuYSVFK85J1/N/QsRw7zsq
bONEnnew5sqWGnh9I9Tkac0UxHEqpZwPLIyBhx6uLJdU6RC6URQC9OltM3rr
hgnKEMABtmSoAAk0HQSiwZIl8dn16ONZbPaeS90t7j3uxqbInW8umHGOoSI+
XAojW28NN7c+hJBdj0M9zRoqhJQpFPsL7JfXYFQ1GLBtL/eshCVuuOWzwKn7
eX+o+LXOQaA/YicpwvUw0oUYuE69MTiy8wLiki/iMXcUSPG2sNIh4kUQQu30
qgzgDLDPTL9iap3jf+yVCYybOpXrRYp9pPDQiA3utVCetMs7fShRsONsKiJ5
dBd6CsC1tHCPlOOUG2hJwHHKmvsfZRM2rISVM/sfyPZIZiTrLPKZWEDrIDSH
WhZd91dOcWihBFjxwp/j7LrUKe7CJcBmm4DM7ily8/h8PiuqOz0mnwkU7Jd3
QBmUfge9Izc/wZhDtx72eySolIhMZEmev8ngb0Z2PAa8ed3T5bNNg5/XwViK
/Cz9IhXiFpDqUPQEyZrCPTerFLAY02YaPyq3VVm06CtG6xSK/OzqkZg3CS1Z
ZNQWXIhlPpgEqlnNRchWtTLRb8y4uRpHug9B52RBbZZrAhtd5POpsiyAycd6
YdysJ2OXH0QiQln04hdjXwmpyacHArfvypVW9128nhQTGDzjvB99A75iCv4r
hyHP2qADEdBSTHvJDt4dywdI+f3LLXePzg4gGJ0UHFC3Mojfg2G4lIqVcUBa
wsj3YLylgKA0CEnOOO0Y7s/yxWHmUWnjPJSbowcKgVKVqsoMnALkEyZ/ZpGu
DJUhhdtmXl3XPnuLl9gthTOPo2Le3EGfibLnBNTJ9+pSB0T/e1Nk5rM+OOC5
m7sIPLjnTypedPumX8BzkuwhozKEABE+GA65z0VbEn1nqXWTtUJrH6pNC/Xp
WZ74yQNplK63Tm1C/oAWFdpE/4mDEDemNoYza2Vb3gFsqRq7Q1owpa8h2GWj
ceGz/zv9Ndz0AStC66Ax90ofZMZRe+yfWlexF2JWaFjpajQRNTsQDp6Mhlqg
1L+Xg94O0NV49I9+I9mpA913wGGTFLMI/56zGdoaGJnG1MSihf9sYAnt6C8U
uSFGZav3Fw/hBRQZoNJNhgLl/sQYu6XQqYyAvLdgDXpvTXcfMtEV+qid1XDO
gCbh7KGXUh2wW8rSerGv+CNpMbzT+12kIDUYcegFlvQymhb+SR0vGX2tChRt
IahgAl8ycuzUMQIftWudl6GDH5rZriwLeUaG2yRQbqmftS77FFNWdm1I6R24
/h29EixrRHj1vpXHS6Hm8WOGyMYk+qFPk+6C8aKTMDl8sOMPA0DVeoiWSBlQ
xvNGsmoqz5sL3KUb3bMfwOQzaPrR+7rJ1M6sK2cSYGRQM5H2xFpvw4mLGY4Y
/nO4/z3Lnz2V39FTQSzUIexQZvkttCTdJ0+aVlmsmbCJobm9IWA/xVQvPd69
n6i5Qrmvs/duvvwlKiOPLejZYnuCP92yd0XZ3k6qBYM0rMJf47PR7Y0AxW53
cc3d4rkIyUNLWhQPwtMgey5pMir57iANNQqwsse4bSRxCNpcPEcQB4GsDG0O
3FgoPxzJRuC6BTrRMhkcZxDQCsLypYOklFFBp1wR8eEpx5NqAsj59kxh0MV9
0eyqUi6brWvZdZaHeSjYLAJ+4JCG+1G/Bt3PupUKAxsPEmHIfFwFfgxsrITL
SlygRfynsqKxmI1vyIP2JbhJ+nEV6aRkhZSa1xBqpd2utUcBRF+G50v1J5pB
omQJ7EnpuLrvwjzzqS7n+D8Fuv9mXuLaeeDdoCPkJ8I8xrABYnGLq8q0y4t/
GKoLik2wL0ZugFOJFmMGng2eMdOoyFTR2pxUpufhB2EVtyKdeqwUbKXXqYjX
n+fuF7wWCw9zbbzDRRiCceTZD7SLsZSPbuwwI2G3ptcz9WPLZKmqiq3c9OdQ
i+4mpIMlgtl/FRXnJZh7ecr2k7CeXq71skb8ib+qIH6L7c24/IJenEzixdiT
7yi84bbe1li2rlqSbOVwX1TK6hTtB8RGXqRZ+qcOYvQZcaiiKxjC3u9rv7Pj
VyW4cL1DilE8YSQEOGwDBkk+KaHYUmXQwvIDE0uoaFPJsCT4eeZGud85O1ZQ
llTysKTrZvD8dyD8iZe0Xt6B5MHOK85pdRIS73uOV4SbaoZOfYF0zqhxXNeL
TgujyJAkBwUU5E2pWmA+xN3SgnONmTcYTMqthSVL2Vci8knDO3vDBJDkOM1x
A/oKQ/HGRiQWx4e1XduUeHC4IhA1ZQAuPQCZbrnLWwcJ20sMlfdEZMHjaBor
PZWJ2XvVizhsSClqkpdsOjJhGVq55TjPapT6qqd+CaQwjyaQ0dU8MsiOvIkn
PD7c/jmeuyl/fgNY8SqQ8ysBQHaCrHxHXUbWlL8x8LdoLqnX08WbMinPFP9m
uXH/KByBQsmcv8gbyIJQIDBZQV+Dl20J54jsv6ok41+oqOhn8w1Kj0pv/whG
oo4Mx31zsEfJ3T8NvlnrVhKUAWq9jjCZTnRePD7ZlXL8SjM8cbitI7B1xlJp
hrmrD9EcLTg5qcffzeu9Ln9qrK2Fkh7ogL8xbKWtIMzeJBvxRElKGOT6TQ1L
/20RhAzIoONJlRLlM4MGEPKIanXVmgt8zz9dGqxJDpIAnPyCaxJPHaHDaMEv
0wqbsc2Ez/ySS8VyOACOFxo2zJrTZmschAoMEFJSny7rCz+k9yYLL0mEmiJ7
0gLnBplcN9owYiTh0vHJSoeCrpviTItspkDm9oomgn1b4RvJ7JcBwIQXL8Hc
vxSe15elCzgRYpapaoZAZvjOwk5ngQyugCirtXljtIPK+nm68hcwsezz5vcL
qDv1KU9+vSo7ImRn5p+XXl2RSSY8w7Eh9KuQPEphaqDJOR0oP5dCQ/2RypNz
oV8NiC0S9vaBubesYooylJcsBRGdoxewB49K++7Atqmv4+V7OpAet3uW6bZ5
6IM7EccRQrJ0iXiA2ZCLaMUxsVYq4eaB8XkqXPE4V4eiHjVVUmTuz3RDTQfM
MEJu7onK+Rl9R/jnizkCug3gXQ8lCtL99IhCFhahaVGTJUMo1nFaSlK1mYjY
wJaAfHzRs1PVRXSDVwKqV57dQy3ecWI2zw+fQPGbZ3ry6WyjfX78PWiE4O2f
rjjv17vI2rhiEvhhwpaU58nsS0I4gjFAQpu4Q9Yj3/oEbzC7HzaX+oA3ee8v
2xSrUTpFoMEjCyJPeLNpR9qPXvXaw7WImmQE4kQ3Wkp2TlYHSwX4iXhxcDNS
4LfhGtyEgabz/7B7hwID9WMpsIJqTqrFKh7fCDDqDIwzYwSaYiT4Q0WMtzNa
+zfyZTWxuT/xcuRT2ljFy+quSB8P/OU8cvInbYVVr2CE8Xw4qib8oiRSXGKf
j8duoh2yJ1kMZUF6elfoRZLCzuvgfbUNBRripeV9dXoF6c9JYXwucMBl62AD
eanlKqrQ3mPEJiAtNloUb/3WwB2ZFarA2UELwgp0Hj69pTjD+eSgJkS7qBe1
RJP96vGzSAYBMDfADtTp+Ts8nklrMro7f/KZQ4WquLO1c8x60PvPd4Q/nVQv
H9tENeZLcGsX6mb/F78c9azj9ZvRhN+2Nrj8vgNWKZ3GB8e6iX8n5HYoArMw
rFQHlYY6XaSmwNJos82DLtkpR0rUAY7Lru+FWK/zfrlhZ/EXYvxRwkKVbicg
WVYVlq++V1yzP3OXFOWsGio5YTazYmrA/E/9aKxXqhNyGAxW8sPovAPFE2/E
CB7YS4wmUMIHSUCz2ASygoXJuFTivRTyD5pAHyNTKmhyEFGVat/4giHR99iU
iJugeRS1ODMi1hgk2bX4NVWlQQjVvGzgwoMTFUjBCjOY68kbK71fi4RXY/mc
UzzRHymNM6r/CDCwpn+0Xna/hQE+OQGYTkHkQItvwoaHetoIVILKcyjMQabU
Co9ev5PVJXxbssvdiZN4l86WCw3mLkgzCsOWE5EOuAFrSq+DQZpSazYvRtA8
w1HtpFEJY6NIVoIeS+Dn9P8YDNlN1F/ug9NAhC1xAy2Mb7mpRgq9M8Itj3Iz
nGq04HZRoWuciigPk4X4r3kddLeRiVnren860IlWPaV1enkPj/2qp5QDwSrC
ScOr/Q7hDTj62LMRgJVQKlPAd7Vuxni/O2Y5ydvifH0OLDYrnbDZCc6m13oz
x7PzsFdkLRapt7TUsyorNNrR3mslittyIGEG7Oc7VpxxFaTd0o9EIwLVitPl
1oFZAihZSAHu3ioULh9RYR1R5GEgboeKA3oYLtMuvg1mWiptOhQnGh4ozbLW
pCHDNTAKJe2j/qfgwWRqHmlGWG52CPN6qgOvyb+0W7RPFbfbAlpdQPLAkJga
3xbBTWrL6ndCeyUyigGOa24TrywFaVvQEKJ22hPb5L93iXMxbNL47M4d9rHM
HVK5o2cX+y+gWzs4A+l7nLoKbPzyJ/p5fJ5UU83QRr7ca7FuKh2wEP2RirxB
rFltRfpMZZPpyHbYb2b/AIJk8yjIbtAZFLqhCpZtZOzwDAyCyIjUlKHLkZnY
7EDWNwheESfb/NKrJkU/u74+r24buvZect0oKDNEexRCAyBnj08K/HINgD/H
mF71MZtt8ZtKaci5CjIbWsXam8DsfMhCfYa3op8c7V73XVvdx+ZnolKFg2DE
hUXnfSXi9Zcr2N2NIKEm4A0AK6gVQCpxJoJPp7ZKMds5GmPpby3sRC5cDUqp
LnzbvRbsul5K+dWy1PMs/yQDmPPB2Ts7VFVjhmbuADecqvYgCNqV+siRElaX
X/488TilKCnkTRUt65LPtCf6n151CIjv9VHlxC4Ta/z3f+yl/D54Nt23k/zt
Vx6G/yavwxQl5NUEB6Zm7tgX9SlzgtToJtyDe2hOg9StUvQObauCNHBg4G+e
onVk1bSSbTnhLwucTrGiHiHkKuH8sBo242H9edqARUBFw1j51Fmuke6gExMl
zXih8u/aKCF3QrNtg3DOjA36keWLzLLqylefpxnPZ9RScN9xGJ2yCnBlP+zj
MpaHhBpUtGVIrvR1antfJRZJqyaTfpoP3S6GaGgmDfVGYq6/dEIDytG5NAaj
nUWGtVG0IYb2uGsQyPmRLIDfFCCwuli9R0+LOMSFYPdzpP8haHY2E3cmkcMU
b+QY6ezFV7G4cP+hAx2u7wfEN53a2NrD4cjmRe5lycAj1gSBw8Y4Ajid0R7z
VyNG3rUdRel9CZ3rQFVqkGTryuu4lwV56cPEclluwhmhiq9MihIS4u57fdN1
c+Gvy8+r1E+QmtY9cGElIf7lcE5oehbNtAMLCYev9rgKBCU2qQUJubkatU66
I56kURJBOsjnR7tfnYBdIu/b2RK/4sxmAWyoGLxGncSw7ShuQuufNcTJGrvs
nLLuFqLkfMwG4x8d/JocPsGIsUT28pvknNEaMIUgdGz3I+F4wmlxXXx5CvoC
pb5EXUmuV+F3cjlefWV1XnekmrgUIg/jKXggUPaKqWzwJAWbemp3c7PpsbuA
RIixztHEAuBIbivX4C/N6VSRqgygRdL4RGQuTuuES1SM9jkWIEfltKB4qEnf
nDDqtoqfLniFviHWL/Kx3z9Vl3JM1z2HvTOd2Screuto2W5Q6xFsdMK3XW2C
Hy5ble7ILGzB/kAM67YQTwzJ7QtadN9MtIClryVBCyy7KvQm3BqmEqBC6Daz
GErMBrQaNEYZDBiaBa8T1CJyX/vnZbgL0Pb+NKfwRa9CPBAKejPr4msKHQaR
jUpVfQm3utHGkdf7Uunly4mjLz9fTxcFqeeSrF+K/uXx1oa+/bPJiVOBwTdc
C0uVafrXOmFaZ/I2ml19J81ePvR71al3i8LGEVPYsuPJlh7kRnore9Ue7siY
ybecztC5ise8TOtlNVFM/kUS+SRyEOo4DSQcvEjiNH05BAN5HpoL6m8o00Yj
nL9pszh/DbwuWAUfpdBvVjpJ6xNpb3o1HBqfRxflHByF7jO4DsIpzw6p6RrL
PU8eHxH33a1yMIRGl0ZuB2vj8q90pF227aYQBnGkAMq9XRZAyKBAlex2T1lk
f3d6R0hWRZx7RSEcIuL9YM7IHzv78H8Z6WTy0n/+uGFCt4rCzj+21jAymWHy
b0znPjuy2Wl+6n9McvN18pR5CRcnQnbWWcaPzJiiaHXeEOJ9/VeJVL5wh3YT
zEIKmJpMUsfj5BN5X1phBp0KoB2X8r8k5EdNqAGE52flLt86LeFbpqoCQLOK
upatiuGyclIvSDlNjJK6D9irkr/0bAVp4fwAtSRn7H+fVJMrho9b/U/AmmSA
AZUIUSTaMMh/eJAeCj28NWQlyLiEcDxhYZQVuqGYoXT15WeG6nKNMikHVvyZ
CYEqGOnjNnkjKIuxGJEsToecyWMe1KC5XDdiBLIXE+tsjw0IFaPOQlvPcTiC
Kah0jjFHph6zhwGInJoX/8QSRgp4dZNO3FEPzzE3itd10tS7f6IaY1eNlIjD
3ttI3ZOwr9D4B9JKO/AiBf8Mme90rWLeehjpb7DyWDNTHzzVMDqLZM+NX8l6
WVAos/aRyHptW6CTYA6XZJQsRBvOhs7/GluLRotSj49OnPPOLT+OCUIi0aBA
X1ph5cyUUBHNJFIYGJPzUl9umYQeU49r5ORRZwruuPLQPfsdrFRIn1fnqn86
kilL5KKNoPYWxO9dgw0RGI+7EH0oTSRf3548cw8arYfgK742CFceowNnF+WA
syv6U2shyBl69nSwZPIn6xUkDE6Qsw40lu3AmIqWgxPu4J+LDiydtTP4UBD/
d3GEAM4NBdx/d1AK070unFuutMQd+lE+PIahdwiwA7IdO3807CDOuoXz8OUU
l6Y3FuE3Px9Zd+VeXnpsW0fM4ThmCPUYew3mDifYgT5KICt9SnqnFKFfZqaY
6Cry/5DfzVVOD0eztdVtz/2D+P7MFisTeMZ41Q6E0Br0WQ08DcFS4hFvj6JD
2I7Z31Ku0PsMePdavCUEq8iB2Czc863dmRF9nmadWe2SdjjDWj5oKuETgUT+
dnbbgr2uMGfWBblVBfkCByluqI/zTE10MCsPtofwr4cgvWatx/7wPeMSnaGF
PdSDvFYPe20/i9taucHQeF3AIUs+X9c/HDKNmPuZCpA2aq+9JtgTaekSRe1s
QJvkAm1rgHwV70YCPq2VTGhhJVmfsiArDE8pMJVC1Ja2MSWpTFSK0gALrymW
mK9gf/qE5/4ssgae1sjGKw6x4NAGNiFluAhCvigVZMYHDRLKiEr4f5s2Bgks
cUcbyOVPwLdhzZQGJIv3XiyvTozI2TdrOzwFYB2bCJH07BJQKUAsYHshEY9i
Y3iiDKArUborW5s/z/OsUoBUTiJG6hj9mb8cVB/3As1PnG3EZCCAkmTeoyhZ
daXQJZmTGZ/oxO1Nnl5kTtRtOPEoB9LhVEXxRZ9pFr/aZ6ILnKFql9kspAcB
sg6Ogs7kR1JuiQOlsNQEFZ9k2xJacxy56XeyKkwiUFnvf2e5Wu3FNO5qrIQK
ZfEOgVJ9vk5VDhkV/EEk1WwjjCAuRcurv7blWHl76Cn/W/PsfzX4YAU8SHGW
1G9BShOj1LezABmojoug8Sk6IbuPrTvG6Fe4t3cWpZj4hjwBpv6jhujcfkuG
71Q4f2TINbzA6VI786rh374y5Rxr3NbO3NN456MVy+QRruyNdE0+HkGcrPOU
rNEIkS1wcrR0rj7W+ngB53hRwKKeOyYBvnkFR+Dq15Jfi8/qQ2sPUKvyTtix
KP6M/MFQdMHtd3x5tAwX/CI/PJSr7BeE0U8Vkq5MWT9LZjJ1/AsB0DHzEKiY
YH12qyHELEYNrms1RG8j09w5dcrsScTELG/3YR7wtkTBjvsLXQjEHu+02l1l
XrJnuB7yVcJQBx27s1JFeTL4I0RFWHsGXBIclwdVvXYX/vtVWj/j9ryTPaeS
YH4IHm8cS6x3sMhiU35He3yKQxjJHcja8LISuUUHK+5+wpWjSPNHRTJyaBiY
WPHWYCXOZ20LiZ6OO0ka+6Cyzx9xRtrjt4ciqDgE2K+ncGl+7MrYeaLuiFzw
scWedRnE6c/E3F0MnPDvEWy5I9OKqaf6pTLgH1fvvHe+BKLeA9KqDTzmVNjQ
eaOjPh5B6xn38nOHyNNpF4nReS3o786uTjOZg+ZsQ+8A347x9WrVTTXvmVTy
+HQuJ6keLQd11XeRodCb3Wq+wzgHOmsASD/0tFvKiuYnqvXb4qnez+V0MQ6z
EqmVFI6ucj35vFW8oQKzd4LGNd+2Yg1AnkEUsh0t7DY5rgCHn6+rBa3wrcqx
gwhjTAfxbefNc1Hvo0rjTakL7Bv7GH/f0poZdRC2AAgGStZ8nF2+Ko8ozTpN
ozuNNDspfOlMQKgbUTHXSSu9latLqdRZJmhtGFThhikZA6RHGXKFOFBd1VRT
stA+mN/g9STQkUhCno3T4oyfjNrjdYc2E8fGMIksO+a3uTTsADvr4lEhvIc7
brMeMpsv+u1UDH+kyc20zr8ALwR/1UcPPCO3Ul2Egpss9MbBvlcYFX8SS7yP
zDR1/xv/2ZgH5PgzbsBBijz0JKiFTbnjn7FEzCJ9Y/a0bJpUkdniKd4MPoB2
r/5HvUXf7LC8LxlH6sIzhLJQN9TmZJiA8Fc4vrlXkXvii7uoDSXB8rC2aIGw
/3NTMIap+ZpQryvB/LuLWn0+mtuoBC+StZFL9U4lLY7uQoTfffw87+wVwYLi
AJze4bbnk/A+y0lzvpGgcxgswZPKbS7q5fH0YC8R0hZSb+Zgxq5Nbv4fEihO
XgJFW1CGLQlEehLx7++bgCAUG984ovU2HavtDoxu8LLzB1okMSiCBc5wAmf3
ZGYuJdsxZ9ip+iG66mh8cWDTUBsTgjdpTeXJn+thfF1unVfgKxCh8yD3PnbQ
mIFXPbgaO+gx3hnZj/7wa63G0qCwIw+epFBUMk7iPAs3NCQeKdznvGAyT8c5
2Er3Dj9X20fX4dbId1dJIEVSsKAVtaQetq3o5T4c3zkBjY4JGv/A4zbiRkUD
tDaLTIuRwPT/i1FerSFj+lafLQmGZxIQZxhR926ZvgjmtPRTTjlEmtmUJVew
U64HyZQuB+VNcXFw+C20jvSkNxOh+Q8QTCkUJTwjoTZV2PglsldQepsIF5ZO
cOWZYCigKiy2dTxdT4HRKNFPikdVYLVQrYMlH/dGQn1mvK6ZzTU0Qt911sxz
4uWDQkZk7vNS07/zEnOOR8AFiQiPFBERKYacDAkbbQx0F8MoADLwYT5VJSAS
Agn++JaB0gDWFnrHXLPsAyLihuH/+f2i2lwZcie75E/M12LCXu2bv0VTYrHv
2Te7u4QLA4Ez4TkyTzB6c7eKkVpnbY68MBbeoYjzNFarGKOUYm1rAFN3ECVM
iEf8cP3eXvHud9NaZSr0ApUpj+a05wjZ+h5XC19wkxOeRjX639hEFVkvboza
PFz5CdHS5+T2DDogyICH8pvlcnANssbL305EWfSZ2NYDKpmC6q8n5L/R93ul
VNmAIe8EwM4LUOyDED22rBe8nxAQUMGUw/JSJk+cQVgFd5+ranF7YmID9exK
N0rUCeoT2Ys8vMCAkD7Fwpk68uuza7uIMdn6v8SZIFiKcygDP8DeWn2DS0mG
+VdxM01HSOF1z7nwbua+rIhyrwUEP0UiCB1HEyTBA45XcqQnJ76yj9eKOF9J
1sn1o93HlhzZMJJfkNt9vEvMSINFKnilO9fs8lkJQmbdpPRl+Grm9GUjBWmK
jYkjJNthkM0lNvp3nicay3YdiXaOIRRWp40Hy3kjgepQxkA71uGBDxl9bTd7
S+52EZnjohTiKfZGcfyGDkRgA5pEndDoc0vyOsLy/FxIHgNqoiS6Jx87E4DL
W+OHPIfvLIR9xJG8bGlshE3ZHqNzPTGRfxyK9R0lLVTMeujnaJIdE3/itzv8
/fCkVQ/0A2RuSJ8q4BR0p2B+SjmLB/b4xC99UtYCgBtMHDBtkXghEa8zJNNj
EOUxH2Qn8zT7Zbt6ITsn/InCh5OmsfXZJGI6IdPTzvZ3FFauMv7wtS/NlTbc
ccGxmC2wShuCe2uWuFld3ipWacx/TxLgp+lCE9eVgKgGlZW+FTN3TWZ7YTvh
Qx4I4RdZ/gMbii5oX5YFbNtKDqCRbpeDs677NrFKZKLuFPmclxG+e+StYR7f
vnv4OvxPj/LV6C39/QNruYl7F4wKXrd7lZp2Wp90DS6dMuiKVO5jIUNxOpJz
rG2xdBwk9jUn0kHSpgQk8aqfpogOk2pzoCIQkLeraTZ4PHJJfg3rWtPwsFQJ
6HjmRA6KS1gT24mL29kNaGEZ6jvS/NA+bDvtXiN/1vgs4aFhDPTksarCRPnb
T3i3saXqFGY8vAe9lRbYrWtKcptyKFtpVhe222Q+4bNl4ig7rKmGTiQcrNf2
1vGZpJZvPG40Df7zgB9u05MgC7GyaUUq7VZf65F7bGwuI5AassOOsS/QI1Om
zoKmFms+zpGQmi7eZZ2hUroVlmFDtEtAjhB0F+jU7XTc8q6hrbumVEk+uU7B
wMB4VD8Ts4IChxgNPIcUdqJ7FDGDVmGEyEvDUs2KpzCwmGKZJeWozfwrgugp
x/IDX6RZv7mfhU7hxvmZlGdmyIMZrAzxvzlZMe7mqCvDgiGlvS8fAqj+GDtd
4caHgBM0Wg/ttRqxiWeauGwT7yLgQzRiN4NjUIs8uqWCUJRYV4X/zkMqWuMd
ae29De3JSZV0kztMrWCQbhtYS7oQtGu3veJQLWKTTLqJt/G/zjh6np461WIt
KieWX+hYAEAwVZP8KCOuF2z1IGUBM2L11/k6r9rOzEhrXiPQNrOtpQ32SROI
GK/Cezt4FBQtYsLryAuroXDBhrYcTJ8ul0YkdRbf5Fq4jTyT3o50WJCopeJR
02LFkw5IXrwpnp9p/qZDtA7UuBplIWwSRBg5Rk3Lq2iLw4xqbshgK6mKm5HB
fdeTQRo2d1J1Dm7J+WJ2vPSMB75SsJWjmEPH6jv1tdXhpVG+91RqziyrpMU1
vLchUKeJfo5LJHCAVpSDoFi2aTP50hx1iPmG59vv4ZWrVkk4zjdz9VFLfd4Z
WoGIEa4r9OMMzN8y+1SAHLFSsgpmACLqU6D5l24A4OVFZOnA9zgxeMbrRXuC
5y2aL1lhLVjas9FDLRdlSZpGXHTb6f2ybXIV4GqX2xIeoK7eeh1pl5VdHYTE
tYUBXg01HT3sLLGyriSVzsBVbpQNWa4b/dt0NdLtwXhARxeJa8CJn62rkr4N
pKjpxYkHG0pdgLEQJrYPIrp27A4N6JjeAEhDyzOa/Cd8YRqU8ldJJ2pf3dad
ESxpbAmVNqkwzDMb9oPGRkjLJ4SNHfDOHn8TKQpdGZjENiflj9Z4tKQagjPK
pMaFR/hAbGkxp0RlwIqSrXjMtJf4K+5FrhBiepIiSIDLplQMCOYG7B/+Ljxs
U+ZZ7NZ4SUYU3ITrBE6Od5Q6Doq01bGY8PvstNLlG83wWPlB/rkclglnzgko
HRPc2KwFdCLtm1POkEhWGadGcm8KzYakUorBQKjO5K650+BoLxc74fiV2idH
msDvDz9K94Dln3RgvcJME1hFG34qmEbIRR10seuu9L1INIZPhuWiGK9eVwcQ
CzNwcFmThwQXTZi+9MrlM1+iDA6myUDmfdz3erNJp1sqg7yL0H/VGRM0X7Li
YF6wcdj9u3v23CAjqFKCdnIKiPM9UNKyghPcz8VL10K03vldifcsFKqR5UoC
yr3y5wfPRYHgTsBvjUKQ0wXKKwyfK/XzgilSQbo3gb344+GYHZVJKDBg5Yb4
nCMooh6D0Z9+N6dsFZkLD+V5mj94KFm/WVfV/j2GUVlHoHDAewAH5OQ60XMP
y4V4HpYWen8nUxb+cr1DgdGDgCXdMU1K5lr3HfeACfqHO7HGAWwD3VZcrQUJ
VuKpw5HIZuXGNaXhZ4jSoPRFD1AV+CLJHybV887mFDBNzjLXlJkDfl/LdfV7
FHcSPFMFhnyvohjvJMiAaJ/077H4vdAkJgC/gqlG+YxEtJ8QzSHTG+TMoZYp
1Fn6x3jyu4sjbc4QYZyR0ywCq57kRIlWaaS5A9QCIL4z7rzwr5wgN89MZbHw
/oJR3PHQxEKxpUG7EU0gUKVCjW1oxXAwdu2oMOtjXdGllGdF1IlHYK1eMUiN
rmyNEMyil0hQdT3SN0FgzPfcrM3bDxqNjLWMqiFv0sc7cCqLY/4YaP+vOj8r
jgJfYJ+ldjzciZyJfRBV04yeq+tBBz0lP7PMtxs1TGT1G+OMFOoCf3bb2CZE
5F1fUGV5Kf6o+dVlLoJcG+JM88id3hhMAGO7sb/KlEj1wYtc7EfedD663bDn
L1TSlREn3TTDYyuBOAuB9QdlNnjGcsUdijYBSV5V3hRJANNnReJCx6u/YCwR
z0eO0RcOq+BuuHS9PCe/msoz1ea4/Wo8XV2kkfDgcQwLmcWOLT1W0KshgXwN
8RkdTKmZu9GQPOrV0evTDCapXw11iYQoSEropExo754dE6uEw86/mvZZ/88M
akar0WfYpzWhFdZnTE5xFmqyXPT+n5xMWWZ2bVYT+X4OOwM6sRyzzrpbd0bP
aFVi7+/cknpjUtUMdlPr4WapGGWQmaStfR3ojWwN2VBhqEm/XJbjRcfQn8TS
sfCSu4ZkWuNaWVbDU18tG8QAkBFq4RYuNGMngvFlZxjYH9KFbhfm6bhUYaWa
ow4xa+uZtsKCAZMLA7zZ7nkV/meuK+Dpgb6nW4SC+cY8npXo6NKSG1DIE1am
F9nVyP+ChbEw5u3nV+BMLH3/73FlfjQ34kDPWWl/5XavCaybTtBaVbsahDvG
wl3EtErFdPKGlERC9hr0Mvd5+J+qCH1bIB8ueqAxMGH3msszzblLY3EIlfzK
A9WQdiswnGJ9kaAyyAdDAYCMcoNtzfo6vD6y3AWnQYXT7Jp0dJGW81T5buYL
3ViyuF/RyTzgRB/ApQt6tHr6bMw5BCABJntx5dBx+qVxGyidrDyYgdJ0ajhs
XkwVMlKeJDTU2MD4+PACmeWDH1PJypX2HVzNYGZDqP3RSMkWZOTU3SFPWJcj
ZokKfxORfCia3LWfBbD9XF9nJJxThrHKbQl9htHPrTyZncyqzxcVdNAQxImz
OzlpJrvy5nDQyZVlzY3YbzW22tgPvXPMuE75P0o7zEm1SMpz7Xlot78cJQEU
BwrRXKRj3xP+E6wS5+zlIHlr22Be9fnb8fRTb7oTGwK9N1nC5us1PKH8f7YR
oiwSMcU0896pZH8OthCQwPjfhSt7guYLLBPs65F90LDYi2/Eq9SX2eAgJnWs
sOWl8EyoD+IJc0fYPKEst+I6dBXHqrjP8d5hEXpSKcbL+Xu4CXHJ+rpASdda
yLd/oJNrvJJv+igjpVAUAQVNRZp48MxUOVPYIk+goU+OCwY7UG00qVU5zDyQ
al9AGqZDguxVHS4nQ//Ok32AYEI2l9fzXAdLHmEtvuhSEh4Jfuw0TfnbGunX
zVagZdIjEPvaR+RgnHXHTS6UC6CSoJZYJP49lY78l5KFhcVQjyvxjCoJhvoy
7u/XA8FXUJlM/UEpv6oGR48Fpps6Ne07U1GUWkyPm2itekyX4YR//2kX/Voj
JptT3dkIZT9TGJxI5Bv375ecCnEG4kjIcSGpMfEmx6Vs4xZWEcQXc2lcKLzD
y7T68cmwUQSr6BRS1SRDTTBfUZDVlrPD8mwH14e9CONm4RpPO6Ea46KnxVj5
7zgyMd8wPa94mrsoyqCPKKIWjheVA8tNFQ2FDVThumAEc0CsMLsRwQp0A48t
8c73TOc9XQHN99dhiwteAc4kJL9+NoiStvnGhn4nhaepyYXfYID6Lrd81SYY
sbpoNUTHCiAp/r+jJoXzM7ioFttyQAybJReYkF53vq8AVN1WUpR9vgZaCbWU
A4EAiA4QmkjcmpKMKq59i8ElEd7yYiJVsemBD+YxQEjbcdNK0qaOPOU9RZXa
bGoI1D79FrpjupkpA/HWBxRZeDn83YTY8M0GTI0tySnvOw3Xj9OonBbqhFRU
+KBzIKSy2P2JaNCg4tWvwEitoY+YD/atdmpKQCd1RmmbdJoBYp4Ofcxyn0Zb
/0iM4cig7jeSolBgKHZufR/nas77nmugriK87A6BRCSSGj/3E9A8x6G+zYw3
FoSZq/fq5LfhbD3ueMc47q3yaXP8qPWq90FBklS3zFxbs85Beomx9BSgLPeK
BvUW/hZY4Bq+gzBCtywU/D8+bz5J79AcrVHYE3R+Nm1pfbgWsfRQGl9eLtz8
dmLTN7nT4VkcUbXCLSRMoSRtY1wcUsfIZdcxUyOYnhdQn9J2hg8K60gr43y3
u9ksCcReoaSDgYVJixyAi0WQ05ZKDtoOQATBpe/RxblRyTp9Nqx3yyvR58wI
niO3kl4T6JhejdhtK7okJRsqesnXsF+KIaFBCOfJUuJxYwUaY5RwPvsT4d39
164oiFRNLYdjalSMzK5hmrQG/zBVEis9xsWgqWWmcHPANmBk1f0gTXii/ZqN
uHi8tOOKbzcQduYqo9lZqv8E5McyElCzS3Dr8srLBpoBQNgoc40My7csoHRA
UKNONy4jvfUSSzeyQCQovNXTog8apo9DciYeTNQMMUltYIiR/ZqwPj1CFDod
PURXqNEnIakaY20MlUtrNMqYEhYEWXDjvpywjP7n+K1O/94v8zq/ljRkMaM/
O3FFHgSfZl9y2H1FreJGaE5iDcOMJS63KB4RgUvL56CiesO2XL4xkzLFNCqO
kD8j7PBUVw7CBlJD+mR7mAVqXDWyGxpyn945sat6FHRkafFB9CTX+e7xyLnc
taVnuRbOMq/PHhx8Ya01pcVUYsjNP+VjkwalJmPWzXYEQMH3KiXXRshICsM0
YRbQEH2bIYpOla7G8p03ub2cyszf/s9ZTtTl6T3ItOmjrFSa9/6yNTvOvERd
8Q8rpCL3x68TiMwUJznkZ8UE7c6/p2nwkLKLmcd4y0FRLPG8o9oMf4YQmg6s
XE6b4ymKeRSAPFw5E+gGB2Ofnhdkc1voYH6evDaQahqYl3hisohYLpcRbsQQ
WIHpyBMBDxvCn/9pR7Gqm43U7qq62IwjHZosimsM+5oIIqu4nvGd3coVpzfj
aToC5qr8hhrM06KoenEtgvcX/Xsxa0Olqsh/qLt2kKU15m9UHNwKee70RHR6
kx2hpJouDPgZmS0A4+4N/3zQWXb5xF635lYUieSiBop90OeCCJfzJ6zi0Um2
vP2dUpd4+5hQ4SPCBj4t6gQ7SESNvr94dkZyW2PVV3nzABi1aDzcC+vrTP3L
t+OC8xPacb1m9j9EiOoHNJlJ5V5Ma0VsgVtcvYGPjTmOEPxaCmOeBiX8qLWy
6J7QiQTW+jxxSGScQhMjXksyX2M20lLMMDh24+XGQV+C8et/4Weuowdh8+HM
I+4phhZTSbGlPbpzrAhQln7oWIFdPAUa0Q4WOH5oMCmhdbW2sZWbhFpfKr6q
p04AJDU4/xCm1LnGos+9ubKD7U0HVi/DnR0dVe1NHfpLjg75Qr4qTCG44uvD
OEiOlrYyNdTYDWuTLjvk+bLZTjNUlIIUFReGRnL9KlCTpVzHGfetprw8jBig
tjIZnBetOg4yqZZ0kY9rMi46XB1RtKf3NSmfpzsskKMprCxwUybhT6MpOEkZ
7THsZxNhVNkMB1KBxucNI7NydWdB6S07IPyeb+PH8lC8kTr0gSu+2pQGC9EL
D4Fz04Oaq+Jra/9lt3n69dpnZN6sTHWwq2IBDETzG+6mXHezdYN35YDHjAhF
VMUuSlJhlj16jJre6gRseYy1rbJL+9LTWVIGhMvuPvCA2DoGNqu4hYcyfdOl
gFy1Zzh8TvSHQvNfBw5ty4ACoFD6RwXMQndL2l7rFBAqHmwp2EuU9p88rA9l
HbeYnozfy6VaTYJDYyg8GBBbMExN1g+c5IZGnnZ+Oa44JqTW+5urWwgKXXcD
Kwp5pqEC+2P3y5RZ68ZR9dNhv52rRbBWZvSmJVHEaoN7INUqIt5os6qjJ9bN
vaS/1MsenA3rXefkRkEFtfqKZ5VQCQx4X14UBj5ifgoNkjE5aJmS7iHhe1/v
p6PMaPCuTXicplLq5xRjW8qatoFS9oLRYh1rYamH6GF/TsvCeA53BSUWcNl2
iKrBmJ9MLB7B11RXbSt8HKd0kSvrC8XLg0fBq6mKZR3z0XNbfQ6NSQR8wI1J
ymLI23n6kiQuwtpVI1szgZJtSS+q/0QNnj40Xi1d4x6UGtNM3irDD7NT7LJf
YK7t/EvkWrQsdIRssq454pjvnEwNhV58nJOj0QnLJY5YZe/QdJopASzugNHN
Wma+9XqaJ2+13qfPNXX8RuKUreoSAXQajlJMnSwAT184A7hrZLKf0k+UnXwn
jakimZb9naLjg+MYf/VKJ3PevLunokg3Lw6kDlI/qtdXjUw97yoShno1O4a4
HaqqiRzGec/S/3b2TvVixXMvSWEPKKgfjcUxdY92kiK4SoC580EtWwBuZ1Vs
zEGeYny2zcn/KmGSC+SM0xzMG8Lb3Gw7N7+X5TXkIT3eb8utCFKWI9NIH8LY
aO5uvtC96P6GN1L2ZQoe73lYlhxMq8P4SIczHRul1yx+vo/G9s8maIopqYnt
wWMfrdfiYhNd4gTGjr+ItFS9AUAvmv5L9WZtoXDO2LcO71R7Az0MHqSD8iBU
WzQoYO436bq0aAIny/nROSZhOLTpz2Dtgm7FCWw0rIaPwE5gmKncrKu7Tsfl
qCM4NOcLlS6jc752bbrNMgLI9RAnmH0RNdF9OfuDrogb17Wz7rwxkHe2YLRn
tQz4X+5FnHeJcYBiQTkV6TL9nwZksbzgsgA4dhUo3MDCiIhvpNVbdxREGThL
Eqz/cGQll3FfZdrUCM8YTVx2jDGHIewAml7MXUG3OKYgtlgcqVJVwOP+cjKF
Hbu2SWbHQGqNxoKCPt2BxgGrVi/nI+o5wbLhve88G2SDRv4IiOc/qpi9AgoO
jV2f5HN5QgJisebvmuNuXSK7nAoiX6Ge9YvfWuug4kPDOStbA2u+Hj0rStov
KRrNVuzlFQ/lBeEs79KYqq3vLdsLEoP/mNWrpVWhSdpm0pwG3M0ZIrBPzRWa
92N4emLFjiuaAogOrFbhDGiBnNoTL1mcP0s4jwm32Rb8UdozBpnHk618qD5B
fjebg45VnbNJYgTKIADobsIKJp7JC1GIBg9buRe7U+YvLM/OmHdT5CUWwYFJ
Hg1jQPmGaCQ4kObpIpQ4PsL36js6Bcb+5vnNlTAnLEzLFh4/c0x5bCzDt9zV
zr6hTzhkO9Klvqsz4Ig7v0NNiiuYMf95T02dcULcptEiPadNiE2RlXeO2B9e
TH7yRC60fd7P3jZivD5Dk5GrzBLmoeeS72VgDQAjnHqEeCEiwB58QCW7wY88
h+pVEPoUEtFiUK3Lhe91KJJK8HL/TYqc8IAcUEIPRBsBeq/Fdxvjj8GwyNdn
yAWzv8rlgLU5wfiwXlagSnZkTBJARM4xOTM03mniBMj2i/K/AnKGny1ms6MG
qAq1K1QtYjHi6/HeKC8ZzoEtJW6HgQiqd0CBf/NBFtK/83cQydlOlGxy/nFf
Xjxzr2fCDYaaKuLB1NynSfaHsw9IdLOFTZftOf0sWUfwygf1cvT5F754J7GV
DI9x56NVJYoke9CH/Oa8W5p8q4upSI5dz3lHrHzia1XL8sRi/sCMCJgtNJ7U
C6tICqLxA8xXJhpGUw3j1ymYA4kJkNV0VG3b3wxkMXMd1WGgUIx4rTsIIy+C
3h11eVPAVPPPAG0lRzrjrK+q59D8mzTJEDoMbfEyJKUCdPCkwiz+pwnI1x+I
9cr0HEj0XLcxTJnQAcnO+WYpRyhrGi/oz8h6HBQm3Dy9+a6umj+4W0f1VkBW
2g6GVd4Wwrt4hmYFvuhIjBapKg4Tu/G/Enpj+7Admh6utchWjQpp2R7WIh27
Tarrkf/asCFY0NR5VG0NEK99lFXt+1+31WcQA7ntu8GGTgpCHYqRBAk+Aa9Q
leGzm8o7NKFF4/3gC3rhc0ZlJ1+f+fJXTkOl6DXuU1O6XCb5kKpsDUMw07Yz
fDsyGcmduPd3OcvHePQ3hdO1fVGUt4Ov1PNk/04F1AYCWmjoOTuVoKDZspDE
zgYzh8hASbNB44CzoVGXk305MU5gyZyB4CJw1gm01eNyPVC4gD5ThtE4UYsk
hN7TUSJRbCNp6DNxMxND/OSg5MmAkDJ7OaU0W5dLC70eRrXNaXIM/BKFOz4O
3eRefvsLcsXpOGbUaLlJU2/SG9GCrQSgVNeumgp06J3FfpoZadQ6/IZHuIE1
ZtD3DqjO7sIBRTKk5dh7oyzOkKWXz1creOHWdC1j+tZ1V+ROacCdFt6ssswT
KJYIqM5LmX8Tscx9EoogYEo3Jn+ZCpfmRbqIR41m52UjZHRRXGQMVIXHr082
CVuE26W+WoqKtNeMVB1ZZPtXa63gP2AiWL3W7mpEwPNVwbWXKl77o1bmtThV
oT5zK/CvxVSDGD+oPxPhsUvvxw1CvwJDxNeQUaEenyr1EXGHQHw6bJU5jgIK
15m5SGR1uSWLYzD0l7pEYLQiy6ooP97m32ogi4JHmaDf6Grv7xXLFbgMQSRL
eD1Vb8ZnGkdVIIi/h0CaoiwYrtS56JB1t3QOZcP34VPIKCn0OyRB3ZazDMAf
v8j9NNpepIdeNt/ovOT3zfT4k/CaU0qK0t60w8zIR8SAWzq78TfmY3XBv/u+
mOuY5iCigWmKaMSd50WzIxZ+gIHxcSu8mY1CPaG5mqJKq2weZ+n+fOxqqAln
VOc9KDu3VixzTzm/wInyUk8Hbfd3+LaVf5bE0TeggS9zQ9TBl2v29EogBsBm
tpwNS27oTMXcGACWwLdgaTo9ep0BAYMd84EjZn66/1NFQ5/8KiBzXXdp2zjI
YkLq6tJ3eVeuX3CWAoWHEBRNsx0qyObGN72KwiAn/yXwgtRzcp6qfa56ORDS
rdqrDhOqjqNCOMHSwoAH2ZeVRK/FClLz0DIJVqP5wA3+B0fxAAYMvWRD0S1l
Etfl2RSccFOvxNv0e01Z3D0QwJZZ8lLDAxasOpD0cCOr9TXGo/QVj+xwRpJF
qdNLZs4Fyp6UBAOz0emWEZQzEmCgYAFv1ucngSyj/ThsHbKlAcWKB5xsK56o
jE9eaiqluFdT/pyrAxrgF+gkKqU0YbeZipe1kwPhrvfm4a+lGBkmNQ6/6/zS
wXgcmTVmn/pqIp7zJ22/Fgt3YX6fSjk65MuMH55EdlToNqiSS1T3K/Jk66md
kV1T2bmefa68A8AENyRVjEzTVrXWUK4hQvrFtX+lMzobq36Pe98WR2hx8ucT
aJJtIZnBts8GKOQQXZi35JGNuWjU6hwNVP98mLESWjWdB+65bhkoJijfojK/
xsWGZb3VYb3bFIwMQmA4VoiXO/9RvtaDR0WtUC8pcXU6Zj/4gmwRT7gRzVWP
r1J9BpHMO+sSNw4NGmyVeicYH0x5rCu8CTpH0B1v58zjkK0AizyoCbDJyYCL
PMx1NVD3Seic7mI7nR9DMeT9tk34ytREWpA5kb3h14nPqX/RZZ16mr+sDHyS
/8ZSmWs8cJOAY6UOtx3vhDPrIiMQQqhwOJGRdJwfWpXNlngczrYzsve6SN4J
kMP6uSRAtlzAtYZ1JoqVU/FZMCtWqnqRQtGFt+zo3gxBkRHFM5074Kqx4hrZ
TesyK7KU5XbkuitdX4jIzdGRt/hePUHRn/n7s3lU6YSozm4djXdk7w6J0Cqq
kEztIslZ4+VSQCRqpfB70ThV0dpuNuH0qu9oLAUeGOL0+UCT+l8OnCTBUCMs
Gf89rA6Bk9OmgZPy9JIE3Fsl0X+rI7Tmbjca48X11NFp/pYCQCNMRxFyjKNw
e6fXyLcCGvh2eUal+oO7Sr88EpznhtQvWyJ37cfBTe6viRqCk5+T8YYBm9+v
WsueTD811DwBlG8t9fZ/EiGyUB7QSoZzNH7BvgHfKU4Xiz7byO9PZ9FSsCoW
eUUClWJcvw3PQNnpKH/8yB/T3Liy3Xkd82wjG7oZ6tnIZF1SJnM/kx6TwV/q
MIUh6MdKYmVb1wgnHHUFEj13arMb+rCXqxBw2KURC6Af0Np5XLz/8yvMO23G
kPGHgqwGu170wAPOrvUaf4zuBM0BcbmMbd0Cio7tF67UiNMfayrV+iSOWtPL
UoqHnE+H89XaaNtLa/BDU5ZjxXFXiogjGX7XHhnJ9WPCDeGWvtg5ddP2dUeD
RGIO22nrFv6fa/0XXZodBOpvxGakEwh97R76ENq/bWZmt0HQ62dYQ2YPBR9t
v/kut50W/q8ZMQWViqYSU2KXtOq/SQS+nLf+Rk2gq7ezKk1sNNU9dXCTnjuf
+p2S13TYt3kbwDHZNHRbZ/Nup4t8cdbeGTBEdaBrfFCghLwwzgZtbzjo6qLT
3tTN8J8pj/WqSMaNUtyz4r60UIq+1YNWlH8UFzUTCUqDGZhiEdrvH+T0OkQQ
DtPVVvJZ2TZkXsCiQbPr04DDdt8iyIIxgBA6Z/p6gdIz/eEEfMFro/QvrMTS
kZY7he5iXr6EY89Ou79qrqMOmbO/zFD+ot3a2T23InWtA2CyesU2sWKyA+Zk
sMUhN/D4tKrS05tMqKYsqiMrU+nAA70LOB7SBH14I3UTJfLITcO7JrqCfjc2
HmJ1YGhIaRhNXvl/v8mtsvh0JytuxXU89ZgwUcbjyBAUNixL7qGQH+Zn+5CJ
OUsfSL30civ24QA8vybwLnaDptUDlHImobdsTeV/zDcH4DG1uR4ekUg0RNt2
cgEsJEfcV9HmagWiGPnUZPADb0LOwHVWSESFGhCLzzNFwYCFPExn/VzPW1J4
hsfrV6n9Ub0UuGosIjiLwXAudYrJGuFzs2ywEuxYie8c/Akizsiuxn/57EuR
vArKlUqqqYcejl1SqQJrNPZci8CSW80yijYt5tXzkogRTHxn7lHLW/fhdTqA
cwdup1H2W1TGnv9EttLq/bsGI1olk9OYGF2cNSquZBbuuMVg3tEX0ENKCYwJ
ZeLzMdlObkpJmaPAYLJZ6CPFuFstHK8w+E/XIjmRF8egf1fbQS/Hz3k9AJ9V
Yr0bRr2594DjiOmSDasRS2M2TO0P988ck3f+Ao4YWkXKaQPcdgWWCX5vdwc9
RQgLe2Hw6fzr5BMhUdf7l8t9p9iS6R/HzRUhvOTiRAJZDpxCGBuHyy9do654
p12HAsylrEy4gmuGFhDtlgz9Z1qNCukbSAdfvoNIAhMG+b/6h8iBCNcvbc3w
0bMAyJBt6QAtVJUACBBUlyOu0ndE+ZKrt0BzhXegEOruCQ/Adhp0ajdesyzh
GCWSt+8yW4FbwZaCnqygtAMa8ghpFE8P0Jzuq0tM8oT08kOS0ip9TV0QLvy1
v/jCoommdLDo2/1XEXaSnFqgciWIBSWMFIv3SHRTGtJ9CZfCTr5DNXixS1bF
JAmcxYtSWSZwuADJrZAoq/Ao7N6f3NE+znWih/QGoPOJIFQpVT8IgLfat3rp
Zg+8dR0JFrzA4D2CHGDoerRRGtDaxKUfLgwTF4NTOReo4il8BDp2rhuzaioG
CKlqV+JaBGcjeCSCg4OBwGIMHC+fX8MDwkKiXD3nUXhAILuFWh/kINK9kLqy
+DP4Ys2yM6SCuDe3bxq4izw++IlK0gUkSguLdCqsqnrBQD7/ERPtqbgm20Hd
OHrIAyVgzm1KXpMZlsOhaarJ2D55B1NpDi6Y69aZ/TdalzaKxVL5YQ14Tf7x
1Ee2R3biKBOD/ziGwWYCRg/E4eUKa35s/wYiIM1UWm4Yst4Uuhw6QklO5Xui
AWItHpB0060kjujL2f2/PLLW4xe4JBMeBzzCHlfIlNSfrBrBaL0FryLO0Wsb
rcGjqhuOdeu9kgothtK0+1Cj3NFP8fYJrEf3nFWFD0QvSLyu7iew+9AnMpIK
NxdzWPMT2UlsJnb4vH4fGxKoN2bV7JkC4xHJboSSE5TRZM24HvM4oDqlJwYd
zSs8j3T0WPl8WhytHMEcjl/E2cgv5I3bL4S4kAFZKQvaZ6TR0ZAxkETcXbI2
OwNWxHHyBp3HfX9HAgI/VfQLgx/VUkbxqbLq5pOVTzWn2d5y60asJ0BcADnR
TzczsitEumyvkIaiDP5z8egT+T1Y9SmPJY/kglKUOOXx8zoEg49/X4MCydJ3
yube0iMXq6nNckRrGVx0vxPpWWjryDtT8poYvM3V82WFIAWyscBZJoRvhLfS
BYznqP5DM9HPX3y9rq8xsxbFwDSQN+3jIb06IbicU9tbZR0xVIORKmxc9n1K
RraJilYEXZhRK0otlW4MQJMaBnSeQtjlijNn4NpcizSV1pXAxWypNldRWEdK
sXmFm4Zsx5wyLgBpi5WoDsR/S0uN+lriap0dctIB72jdSFIXbwCtIw4KKwAA
3T2Hu38kGE+T8tocbb4+m32PXPWAHBKoGT7R52bX9lK1sFqsHGdtTE8Od0e9
3DcHXzOhptClE8KuHg5LRwzvzssbyjVXe2JNPyUFzpzS+yGkTpk/lHCwxFYZ
x/nLhGLNr9naSTFlSOvRS4wZsVsAalbQw3Xu8BZF73SNpyqF+SltKSmdwZrh
XebNCdHjGY2u6TIWgT4FBrJjiwnS8YSwBXlkBmtCr0eitS5mR67LjqX+abMo
WkSmD+keOkd+CZrV/EmfkXTQr7wD2yhbFFqHEZP96FqASOE/D38ULAw6udIF
wpf+NjPsEZ3mlUeSe5APz9cYD4AfdGq6EQJojziJbszn2TAHAtF3R/MkCto3
vqbCIgKaYoivFkPSefyQRj0/uTgnmXOuix+zO2AiRr5rmymPKL+FZjG4ZYpb
+P9b10TnFdP+DHFo3hoWNQaVB+bn/py4p6tIAgccytsY8gKp21ib3WfEeSpD
8o4ErN42kCbirvQf2PkCduiHb5V50SCu10rXGMsBENOZBwP9V9ZdQDTiIj99
92s6S+YoNvm8cKCHaz3EdhgY5Ie501pRqunJHmMNpizitRCNiUr5O6zZP7QE
TSqcx5WlM9iVSvXsSQwuGBOBtV1RbBt0vS+/msmYK0y5rmblLFN5iedIYAuN
ynxQHgy78zcH+bFvlhRqEJVI0Iy3oD/TAJ2lloD8sotIZjjpNjOeDW5fSvcd
bt3hbeFNGCWFYKEcoHXILh+Q5spxtMPZJ4d2VqUYxl2w/KfiD2RRAhdj4o75
/NQJ4B69ubwt5JUHWzDPHOoHo28CKKUBi8vwwkDpl9QvuC3CK/aOMlfMFY+K
txOAHF9cqFauCuXjuX1odu1rJZBcSxEFd+U0Y9wZkiM4ojlo9e/vZQuWtcXg
5alIJTstugpDL83uvc3W9+FovxIAbojC5GE4NWrr1eBSo9Og3ZIVspO3Gvwr
A9yuUotDrerzudN64qoQNHndVDKn5UAqLdDpkZAQfJvKG4K3sZeSj8yZAPVn
Dmk93ZGIPZ4ObIXklua3RI3EVM1r/jp6mjyB0YqXn1te6tz9XOE9DH3TcrYc
dEJ5eHKYmeNGA5zPjBNbbfO+/ox2DgLr0cP2Tfb+v/wIiJ79ovG9u/8YWHi2
Me2PRbRFdVQ0bQDOe6tPx0rpKqwiE7et7SJUhoqv0KBg3ZfXxJ4suGgbVO7V
txQEcXWgK+34H6bTkPPaDdYynM5fK/lcIYgM74bFM7dbuZz7//MWSV3RM/kv
IcTQfM8qs6SESYM93AoaP9yJhn8HzY7SVwIkSKEcqSxjeHIjSqbygfaT3NP3
BWvkmvKR/hWS3z1n18cr/C04QZbEMyATx7gxm/sguZgLF+euNojbHfl2fpuf
lKar1b5M1pnC1QS3r1CZ6gqGhNCgIa9aXEo6sgRPEA5v7lTLy22RJA90E2Iv
5hehmjA3z0nc48Gq6ycBvtu+QpFc08RIFvDzdZV4mWHtveZbYK//ldfSiCSi
tzfna2b/77Kf8+HDM5WOvl7xytXFkwaPFWoYXKcnIyw5PefpTAk+G08zyhrl
IBIgqmaPFQIIxDXAckoCglEfBPT1bOu9UeeRj4IS1hbN3OW5GYwG7zWon732
AGF13cinoXwBiKbXWNLDJLZ5FFmYk8+rtTj9lXjpbjNmQJL+fPhyJlZdZhEd
a7Tiki/T9QE6MW1QMoDUbqDdGIbFClbryPB5ozCsKLbS2y3TOm+fKr9PuYL3
UBJB8neueX0Mn7cacsySl1RfPQNIfHRwqYbRT75AjKzNJsz/YIjKjBoqWx4/
cfnYFNEPJsD1NID1TUsXocuGt0y80EouLDSOpuCPWn7PuD4dbXx1UKBtcPT7
37f5vFvLbeDNQspQC/OpR8L6+bWgzWYZz38eGKBrcKf9YG+pOVu0uxO2Ss+8
ktb28uwp5398LkNVeOeBTla9PXQR855710aqj2W/bQbmOyzDCxjl/jlZ0fY1
Bb1VglU9M9bC0W/m/13279ydY+xiS35vsfDItQ8XzG7RGVcFPW7LOXRwWO4z
ON0ugcnWEkDsywmGW0UBn5ElefJeAq16YM+TQvli3iB5HvWY7qqVKrjiZVtf
5Bktp4V4jUmcwK0twR5TYZOcfvFgC3QMzGWOK5wiBwA+uW5N7/xhyQv/F7kq
ZDzAUwwn74Oyr0Lo/NrrV/WWfrNWsyuFJjvVKhl1P8o43FUaUDIqB0lg4iMO
gnItqJqysIVefYeZ7oGMZn+EefOrdkL7a24wHjDpye4OcRWMdLV3mqeRIERe
TE3dTeudAeEfjmHsAUdurGD1Dc8KXgk1PTvn6fhr+IVJ54k/5dmhZfYSIpLB
k/2Yt5rjmHBZIprtBTyhe0e1+ZpUr1HXIeN/gfYW1LaqqAU6ZJukXV8cA7HF
pHaDJ9860mReBNdnV8cRhvFlkGYnBVJKXFbx4ySw0hvWx/d7stE/Xg4bhAbI
+O0guLfIpbapQFiOiwTX/qW+VSHbpY4Up9h5jz5X6EpNqs787EbBn/FGzkvV
qA1R8lrmvUTotQojJXw42zV5RT63vKcpAJo8NF266ZPUWhg+a3VVqapRw3Ce
nWdHIRX6Eh5th79VxevtsdNBD0+Jp7VPz7StwVKyaRW91gtYcgFtPRd4k2OJ
rMNvUCD/Q0krPXRYxZzNdELWywJuG+DQUBKa79dSD4v6RY4F2Gd0EqOSr3dg
WM41uSfxGkX60m4feWboSWiVrvNGOL1B4S+ngbWmPbwxUBWzuq7j09g5TuYv
mTldzkW4QWcLil6rSWQJqso7D+xLQXf7tlOCowMCGkCOV73fmgCqiJePHPDK
OVi5yHM27c4WzEJQNVoCTrAk+yn3fU2+L+zn25lj8LMyyYSLmN2JjDNdfMXi
1BTe+ih/4pDMbsdnf4m0GzIJRR8ZOZiGh5Ts6pgwLPrsXCsb65Qlza+3cY39
WyyQsgYVLmfDxWaLJcw8rz8wPcdrFy73fKsqPCVvBndkF25GGF5Pu5zAPhXR
59e7Zji8Y/ctCvaprPVzyMHZzCJrLb5ZNPLw87nz+J17BgTNWaiU0ulsWOFu
ExZsyaa7BtmLjtH8HHXmB4mijEmRdQgg2IdwZKXEft7ytEY6M9A6PiLCUsoJ
zxhFQsnryUmhBCA55i/CnituzM6KfneBupObRbgXNkMnX08ellRQCaYaws+C
H9xO5w1dsQwVHiPuiAdO26p4nQkYdNo+6QV97Ypk9gEuBKuTWVOr2C/804mH
WCchCSkdix41FN4cxwm/dUfzWVQke0sp3QOKJmvhjJwvwi8SyGGcEymGjB4A
3PlJzFU5fBaFm4UROHC5dakrNBiBG/AH4G7XG+Wj5vs2M+PWxboyrDKqUGPb
jA9Auxbq19OEttBn1Lug8ietLE7Rt9KToHpw4Oh2UpJq2qHjl7dwhY+H7ssp
6qzLn0QDwtH2w68II1eqy+v2LynQ56hPMu1V/USMhI1oZv3Y5KUNnZdx/zMq
/7Fu7xZ73hXLCjbJcd4bFF/rxHgg1Uye4FUlEZIWBocEjEy3R12Lc3Xh6cJt
f4gkwS1HnJT8MmGdIYlSD+rwgbYy9U1Vc8f2wM1yaNHNFUTMx65Hmzk08QtS
9PaYlp0QWmJ38QWfspWgIRMru25zWoYm2MrmGpG4Eg9Pds6bCEZekhRh63T7
T2nfwzjiWudfFEu+G6ZC0+r6gnl9EfsP9nfmur2JNYXPVrdak2QyeVEltX7i
dw6dtSfEsJHPdQ+iMlsAliZRJQxsTNhnALwDJx2tztGv7gZrdkGIJWXh6oNv
Yab4Dm1/Toa6TsfvTzkMUIIfI7pSShqei95OBIZvNUFqZsWCzTvlSxak0oKD
+dwsOKYaTDiUbAoqcMfgEV2/6FAN/piGsK04yMvO2nmcGvqWA7PURB2XzYH6
2KdB9IvCvFTxHY5WnZRyinFdMDettw2iRf7cqL4h6VHJfQVp2qaQ8ipSD20A
0aCxaLT3aMruI7zQhD1BEdJf+nYHKn+AUYgCp6pvXMQYQCNc5+/ubc+gOAzF
gh6dsKepIwGvxoHokZxLaDtoDAsaUvJu6IGRoHyFFfw66FqQiOY9HvfD1KN7
v1NzOvGQIwPGxLA4Vn912MUKwkwTAUUS3xqJhFpl/hyRp/gQF6KHyu/w+l7E
2kDWQp/QvIjHLhHzVtrDno793d+jVZAYGLJnECAZ2YNk3yOZocy7unGDqJgF
cjzLuwYvJfNBl/HjbQLJrQBjKfnajmPBiB6UQ1NiiwJl7fL0jFA9fIfat36a
JMAHLqPjlnwfI73Yy5KqHSeN6wl4gxBJf1nh1dITszr3B+Us2RnfxIy6/Il5
KmsA8eFJwcwBhoLPJncGac//nf/JuZwk4aoPDLqS9vT/Nu2zHdcNX479ToVG
xAo4aWN7mKyvUez6DW6jDCOqrS5DuIPKA6kl/VLx3Bds/tDwytE/+bO2Kj7l
3SNITMq/ymaN2WvY2OjqVMnEi8LGT2oQ3e+V/BIjXHdhGdpzNF6UqZGB2cNn
IPAVZrrWDrFfc1fgo2bh7Rt6CdLM6BJ8DaJfLXkhm34b6qhZjsdONSFAfAMu
seWKgc8bnqumk77olq0o10wrf9gvAhXnX+0N1YPlMMg5bxQpGzHv7DZlFuGA
Z/7tFwkSh+1Msex4lui+wgZ54EPQAcznkUIuvKSXIMvMslkRGZFatLBg4Im/
Uq/3tGIqcUhTAmmV9jH2mlkrb2iIO+oWgGZm8fNhZG8oE3Bb1oaZiR3wT99v
tKApCMWiMbiD/5VnYBpEawMux6OTNNJnJUXahBz+e6p2fdw89wI2ztOWb5w0
mp/0caCCSr1/2HUXUSCGjzKNXE36BevlHgJygHW5Fx9F9tLFi94Hq+iLz/ff
XkGXNnCFFM6SjFMUgjVEbtCJI4wIrndDYXD7VSxp+LQr6KO612MwqGifgnWH
CHS6enDsUUxNwbRzApc/voM3h6cxFkuK7QIUzUR1iKk0+CfdEWfSPQxfOxAI
PEg/d5GWYoUyucf/eCgJglwJ2kPt+9r7YZkf5wIla/352utn5pZ6EKIErsDF
6HIUoqTqkKFoL9+FuBhs2uq1QD4q0UdkDVXIYuDvLukGQf/rgyhoP7aSqKJI
ZlaBomOjqL5dOhg2gLuwQbq6p88uS2ZdOGMRXdVoU9kJaCbBfRo/bSprF9dI
PX0+/A2DyE4c3CRlvVRzV4rDO+C/p8G+DJMhlPzDiOMnJ+sFWNORllJkNgv2
nABTzEK76x/+ZocWSN2T1jucFZYahPDaCU+MKh/7WQLSjRqNlL2Mm44NmZIF
E41DmGHBpjkYtzOVfCZp8024G0jf4+8B7hBWjDd1N69qc3m0aQc1IoSo8o54
hsgR2vWg1hJbhN7hDIokLA22Xs8uwXqaYFl5xewlxFuytwlMaqVT0lE9K4pf
UoeobCPebLna1ZM/L1YUbA0iOjdzPD490i2pwezBG/JlOKOu19E02erHMMfq
YPKPx7hQ33U0rUU0aBSQxBe4LKnak/hDgJ/nYZql2R7bYVLM564zpeDIbPMt
MU9+Fjx2cCBymt3KP89BvDO0P1/idPqke4l3uo18EyWE5PbsKKFEy1is97Ll
unDMzByPBG751HztQMLXIrsjnWCzyZg9B3YUDLZOYdFea8dYvngk/oQalZ0D
RH8aBnUkKZGeCSZp2UvX6+gTMbDYnBCwlpOkkDBeoHEJF7+mqkrOYXSreGJC
iNiKGK0IxLWxch8+tR/FevN47QxH1r65gLC85RiTTgCtx0WMhYmMuuS0Fri7
77hwmWQfJU6USy+9kwShN7Jaq7ucvnzLr00GF+6Rb7eoQHWYHLw4dDswzCID
1yHWrCf8TkUIXoOMBioplmexRnb0rXK7p62F1IolIcYt3f7jvutCFUAAVxtC
PIBEsnHOIuMHoU6iNWSh31vFmjn7qpKNx85Cs2mFziPitiWuVhPrR/cqxQ1H
9C5TbWDFppleRxyk5aC2g1OgehU31sAibQSdliYmxwp/IeSCLYDuRl8OWX8W
y6emy1mjIc3HgDNiXF4mp+kTscAA9ZyHBYX3nNEOdXB3VjAIy5GyuZU0Or2q
WkkoerHPLa6ZN/Rd1GMZF+hzUQHfR/wxOntQRptFIXS5q5gHT11zvKA0tHCR
r1hW86xpS/OmSTH08YLg8WNF7KhozxOCF6tw8Ap8Rf9acvqXbx7BPw+ypLZb
cqZClTBHZpdtxEyWAsXcogVQJF7/UQQd5Z3ANzr0x0cwPOVuo3P2ZL76cNph
OiU+EjNElIfWT+TsKrzIxa2m7Hlh8e5fdue/2vSKh7je/uMTBfBqYPJjRU14
qpbIhfUl3J+fR2d22uw54FIY76ZalpZSIOup6fGZi0Av8peGqIhBabh7zHlF
5R+U6vdu1m2vkGdc+DIB+efnf3B7kaFJNS3JfIPysyRI/J7sW6BTQZfedQPD
bi6wK3qB17DftwjaV5LJwq791gyRL5h7uZkYnZ0bZe+vHpoAJQIsLWKkLrop
cmbYWnO4JxUy6PXoWKiVjxUvK6LNoKx4gj/33/LZF+TjO5KPSaEroiGqN7Zj
LBWtnpDuQ7qeBtHg0VpLr1V+MfCxrVb3HMFuiNMQOxFeu98SnL3iu1OOPa1q
GRwd/OrxR67h1NdmPKkDMtx/cQwqNE5JCOyfUyc9QgfmTWZmap0TFQOe11J4
Si7TE7yRs3E+cMdSoK1Vv6sB55x6EeJw2vF2SD6eJW7NKZHaml1XqGTvgz1O
KDy/AbLzk0ctTx1yHOEwbV5rPRFfI4X8XvQLA+BgMQJJT9vsNWnc7QY0aHr8
fYvssNbNfbthcGGPnCrIQYLHR2m4XumkTT/lVJ7amCJhFqSjPoqIgFh7Tvfs
wmdWLRFBkvMPjqiDCAphzl6LrFK2Eq+XenO9R9cchQ63sN2RS+43LModNkEL
+moX+dVDtURzv9/QvFd435DF80a2Dt5U5gJuUOEwuD6k1gQzQXwIIwHNha8D
30iEKPxN0rUFjDwKAeln29duMG60Tme5k8se5hlNdVlyhsKsVqXDHtHsLZ3f
vpkw1Jkp7tFwkgt0q8B6Sg8TFmrEGFkIkfw6c4Dj9wOMvNJk8+Tpjrm8I2DV
AGxo7ptdeP+oDXFMqfl4R7Vp9soaTtyb2tWAAjJ05u9Ibp8OgZnsW8p9p5BT
I4riQ4DBog4ZoesRIV2/UyCQBPKNPQo4DfA6oWbDphJHAM88/+ag9+VykBGv
t/w35VanK9C4elbahH4VYde5mF2CnHJSpCcZrRtT5rA6sp4eW5/GQYNxca3S
NbreUqsXFzdWFcITwMnI4he37hAQokezbIoq5HCmgDbIJBCaiGsDNKkDFnJc
93g/8LXDXD4khgFpOauIhF31EstJs6RbEc7icokX9miyQh3GMOMi4U7DrdZc
CpgPi240UJ/bAQomB+UXkJSOmjhNgqUbLcWjcZwCm+5bXIBU5nX/GcUfv4Fu
GGm38jtUDnZT2SN5MP8+05juZwTcysqw3wxskG5i2dmCYBGOTj8ar5x6M3Ew
szO7m3RxCkdXSRJhdUesQ241InmgQCWSMsR5kkRdKTH0W2QyaQid8vgV8BLg
1DV9nMccI/Hnfx+j3ePgl7HNhzqORU/RcRA0jEZBRtgFB3MXiJa24ErdDBXD
MFOporWazA9iGIAQUsX8gbkVDFz9VAhOcmCy8j1ivm5zG9rwxPoPXmDGBxtI
4dbgbpJbM7kZrFWIlR100wpWFTjagRF0eg5hJ8o4z9yqnqON5HFZmxbprR5+
2oCsn8UXhwGDbZJCsJyIhtV1/meUtrEnsJ1BMipc06mSnVSP79mipR/uRhbQ
EYvR90kNoSCLCVVIT9NeKmDmnkknO7EW408kZaQtsjnEelK/ZMuZnAKMGb83
dsj27aYW3MnP9/vyTRtvjxBP+0NcW8lPxgnopdnia+ctd3CazQ0Q+1ihiheG
dw9WJvi7c+P0ijPZY+3Lb3yy3EHyPI4TUmVIdu7Phv9VosajQjkXMTp3youg
qxpn+TR2YaVKHA2PwR4xksE4YusHjF9ILh65TgA0SEmL7ETvT6Zldxa3Pph1
PzQ7XSuXZgtZ+ZcATl4ej8eh8iw167FEwMKPVU6A6BAQPaDCK16SCS/NRsGW
d/w0dYM6NIwV/2LQ25bCBJg7CWle9NJlmh7/wkbUy4o3plPhV8fVgPnmxoGl
7w5HArcjWrV0ARKuN9LlQdCCouvFf2o2Bk0DU0bqgCUQplY7r63D71jod2XA
IZ0XlU3/99HZKF7s4HcFDPwABwvbWGfunez/zxPoNUMkd0d7CdI9EMCxYcXX
jpnS4kY6HR1NYNr3tIEjfvQuUgqe57vyrcD9L0/Cqm4JzlFa9bK2qFYxkJ82
Zc+aXaNyrgd+JF3JtyTJ9mKM5q5ufqYzWW1kG9fM/jZAMhMedd4KlIQgc41f
CnA8hMKu+Kgc1GhNNNsouuOmImcI7ddIYT5ZVkGTyEkDmVOJT7Wj/Euzemx5
3/LCdQ1BIfGwW/mHG1rRMSm6JsFrEfjMExHYbjItsUhGenH0bXbXsAVxP6BG
itI32dr+HdJaNFimbh5a56dCfLXk0v4+54Hnp48ZH/j1a1k+hPWUHGl9manu
WmKXVje3Id5v1kdDt4MvgmwixNSVMj/BJk5DRNEuaUbMtfV1IVOz6HIWICi3
OQ82pY8F5lZ2dZRGgo2tw1g5Fu9a5EfO9pBDaJDfysaR4dFldE2ERmTSgb67
rDRFAqcu6/Abn3Z6dgOYmXjvAJcfL/hp1ORrM9uWna2sBUPPhRnzXRltoQC6
4YNDdPintAVXgLC/3O32+wNkOgUc5xtXZ00Yq2ZD2e2QazKV0VM3LBUhPwuA
7p8ZSj/JoOM5plPRRIDV3Xdf9sRKHmkNtKUF8jL+nd8gGu950GlGgE7FNdZz
YFqEvHzgMRvFDGwPBE0pIJLIF4vH1+2XeR++6x7+yl18E3ys1rijcSDvZtSz
E//stpxyEJXUdgxeaeT0Td82QJfvBaAQYB1d/YZr3v0KYd/1ulzGqSlZTQ/k
e/8LNYVgEjXdH3CpTLNpDs/+MAHvhq6pT35vGR2ozf5OkOxeIeJMhN0sCdCg
qry/gGuGkDoM3KHvhqAsnf/Z0kT0tCDVV4Miey7n4gsdPwjbY+eev7gGy97O
Onl83bfnzb+SfT9/+yXfpFewFDBDJ7GyxZLwL20856K7quMIrMFIk0s258na
knVyUe3Q6UAXPQL1HizcMUZY0I7xqI0mpvE+uP+KdpOQ1vvScAHqIKJf91u1
L2gXo8INxNNOfkOyc1BYirS4zXsc5bibNCCIx3HWCH5crrTOBCYahVkpTWDD
hCcVu0SUgGaRsPn6oumslZ8JlfH3wjkJv7b3CJb1Lhd47Xu2/ql52tBeZVIK
1z7AprZet98lv0pJ/ziVa0iUBX6tjzHDGhWk6M0tfVpyYSYSsnkj3G1cty1I
b6K7hcTYwbTuKP561uHyjJF9he4uT/2lcadgBbiM81EGONGf8oepNBnWaG0S
qnGw7TExrsqsYQKbXRqLrnjo/uKH53Z8aUNGf52VS8DhWBZ7v5vdjoLM5ULz
v8N035WJYwbNBmDtYynQOSpOuDoKnyEYAiNz7/eM7h44twIIpIOpOHw9nVJV
sz5lmyzV3y9PNkPjhCEqBOGLUJo3pK2wxdfmyKOhk3UGXsiAoZC49+Q0aP0m
eizu9XY1Rw1MH4fRVOkfoTWSg7LUw97qKz+0rC6NpRzPeSU9pas1tgd2zUMu
rFMWh32c5dP+DkqpIq8HZcvDeBlQhxl6hj5qs3inXo/uIot0MP/Zo157eo8E
h1i7vsmKc5PggP2Muzwg2NhK1PvjW+97VxMRRb1XUwhp+vtFDJu4N/VwJeQ1
JC56CFQWgsFQ/Kr8wNkCaASCmlr7ZrX6Lc3E2edhoK1uy+8mjIIzRGHaePfE
VzjS6mdeH21A/Qkoc1nRuwBvQ4hU8n+7Qt92E4OZpBAi1HWH68U6hjgbPQT5
JJb2JE9xAxByaqyhux+hikmXyynQrP42WLp7eDaS4GOYfVaHcQdThZdLJlMS
5Q5nEYhMpEHKxWWVQajv/FBA2lx9oIcvtjmgMDiSuNOMZ+TAf5vdmJoISCdB
kDjB5ugoVmpK0r/9Ppu+A7SwbhuAuxbC4NgMffKdMnyHaw02OiPba6uY5SFL
/vxbSW0sp3kJu7l/aZUiOW9p1j3Eo+b3Rak+dHKCeibyNG4GrLrltEZw4I0W
6wH0ARXkoS8fC0MKzgoQIVB0YEwDOD3ooA7Mj4/6UJR35XwIHL5VkueHsNKY
gNOs+FISKBLTO4gENyVoC03DASw4G+f+iKQXrPQKorCEPZnGjt9fmI1dLR3Q
D+Fp8LZJ0BTqnN6XYJPmo+W0dSE5CjA6ZKlhgVYq9pH1eA/cJIR6cqNWew7l
5UFkFGxocT32dGdav57FFUR9N2fdu/dMkOSxxmkqmTnteSPdXmqUXOq+1lTY
NaSKz18KrH8MxlM7Lr6wPRAdIGlq8vhVQk958QMaaOiG7AqIvZe+IV8ZhkOH
b682rhIKw/LFhmKN5E+aWEV5oseSjIs5pglqqVKwjmkUT2PkeG7uVLG4yKR/
JgONW6D4lR4VCBWgTGoJz/ANbJ4TuG+ZBRJ1oJbZTnvqwyQ+zZxy7wK/vANu
COjhlqMzKoDr6b0nK9kXGk68NVbNkFIOdOsciwIYfJA58hq4/Gigkrt9w5lO
5FTkVbAnLUZL1riztWtPOWHnQegKWz7nEDbSgdGdjXJGX/dYOuN/ER9mzJ68
UtfmmFUWbS0Yx04eslTsOqPMQ5H0WrrjnkRiooY9WzNbIGyNq+VapWWfgZgJ
rKSX+Rwcmng/Yr9IOAuRx+38bIcjxS+c6cycCua2x9VK5iY6uqgTz/9WqTOq
GNguArXOZhJ2J0xdCZY2YO7d8qiVmFyrmJgqAK+gD3ENSD5zAQJQeVF6Xzc9
9uHMwwTFXk955z3IOJOo2b2FwwLTzgT7gIpdPnkL/gwLS6EXu0P9Updb5sVC
xBwSWuhFKIAaqVgkETD6D557kkZowCto7b5ePKEE3RX4z6GnXuOx27PdR6Wa
WClEabkjrwrEBGYslCtjG3TQl1b9GvvOljFjyGz3C268iorWSqEySKHAbtvq
2eQWt2b1MN7MTcUs/eR6LuLR4PPlGBoB0OOtBL1uF5V9v9FtwaED/EHdHlab
ryOQK3wLtFibA25ksrnkGmedDLn632Bf9xMI8a3wI/kXSt0pIDVGn1rU+ePj
cAu7EIjubG9gsn0TJY+nPbk0uc648rjQC29e42+SkVTlgN8cccJwjpWAjqzY
IyTWX+WnwCZ1sh8WS+VgneZ8HgsEws//mmHxpHgezVfBmoW8d6bbup2ReZrf
cvC1bwgxjqcaGqtdHEfdkWYp7uUBiezpGZt3BQIcXFr2sFzzErn9f0M+EjjI
0FzcLpTSvUUeJOs6NBj0SmwccDBOYzO00RI6Q+1WKly6tmz+58Ru0bKz0cWv
oHarXAabdcygm5XXg7N70rvkFcxcJK5MobqVb4GqwAKyvI3StuTxnUewxJQa
BbRMOatMwHtWdYOS7jzni4j/Z5404UzgxkDv4aQ70VHbQzHTJLGTUda/3bIc
SuOl8Yp1FGpnYYWFGvK/a3WCPKocickDlSyUIf9oIeKlLOAS2EUJEzwNL3i6
9LQIDNhfQ9Mu5aLhPbpQE/M+6Y+BCoauubzXeb2+1T2YddA4IJAD0duyBIKl
64GYtAfdQBRBEj0qBpLr3mUJMGljqeh+y0rwCF7efdM7oeST6nS+FuLbdPnW
Z+ZnUci2k83q3iVKKC/Oq/XdJK9SjHJAVSVUFek1ANw4F7LXSt9PbE7h50D1
k9r2avWEZnkEpYEJFubYwMtdrGbiTSWouTz0lKMnbj3bJJgyU/oabUj7t0/A
03EtDuSOxiwMpzMTeiRqyJS8ydXkCn8oVtl+PBkLhABSTpp2WW4dPRD7XWVX
A7IycCsmnijsy2Tietcw7qyJnns496Y296d0P1BBGFLJ04gz8ncQP0BWtHBw
LfLphX4pk/dHl/SoAkIz2bPRTZqD5zqTQNein31BwHNDDyy6hCdqPckNpdL4
25DG7L6JlbawyOj9rDhkYArX1fWLd2CbOyUyaY83iyZq9fj0GkE2TZI5n7TU
6ojHlGqBC/xfP2D5UrWG5Icra7mgXmrW5TRv081aEPAzdNNnQMvzGrnFBAIg
e4UBU/0mxq6g1cZIXnw01y6pViFcbB9Ih53Wk0nPZJHisuFsndeHZEJfFJTX
60btlGqRidlIQc3CiyXCWAoTGEH4wLZ4sbjuS5CYYzAPs7O4nHOFUFBfs0uy
EJ0k7q7fwgG8JhPAqUgQ987FF471yh/t1Wn0k7Z8i5cpz/1T0QLhYn97v/S5
2WUYVXbRhCT3+Og3G3DugFF5eHL/kQfNo/4ahukizcpDlnnnH0J7IqsJ7Lg0
P4iuiAMSvm7lJWT9VTsO96QjWwMVgkylcHrXatHGvarXax4VguqTPLPxhGsr
5CKPcWqEGN2QmyjcQrxokNQamaa+EhF331UnbxHvvMGNkUGFhyFhg5nQ22pq
WfjI4ZFI4w8UOqdnS7suxi2mQ+gDAEFtCQJupkJfdbgt8+87bq1c9KZkrvWg
8+rWiQHTJmldfFEfIcy9Ph7meBuhlusF/IHHtfeWXp8nwDp5XoHoasoQcpOb
fWad1cDswo79zPSikl9KkSU9Yu2vOqMJ9UsjTI6e2NVRyTkvDB57u1LHJunD
53nmItQuQ5109JC0u+F4I8c12jrwLXSghKcCMtJdOf1Q2gI5t9dhOFSjJmlq
oiqYZNBSn19wxYbhJTEKECTwZMpWS5eShyaxRLt9ItW5kW3JRBkhZQ0WPiQ/
FZuZ1aFwaD2KaZAtcZJSRbfCXkCzWXq6x8ani/gM2HpCY5JzQTlkxKyvQUyQ
L9gcUprwA+uY9hzEhaYkYW3kwJWa1MbC3Ez8YCyhNzb0HSwzlrBscMX4MLaQ
xAFO4M9wMrLzXiKWdI2V9ZTpGnANiRUgawe9ezBf+GS73BkPn3ua1NHf+xKF
mjSUE2XJJW2DNhDyz4p6xH9nQRE5Bq78uZNtT1By6tZsxMplIWx1oT3HXK6s
Sl4noVvO/NRKGtZ8nxeC04gf64jkAPyOKhlPrKscKxtpTCTUMPOl433m+hCA
jTYipfPNgkqfMPTMrc3H2eiE+fKsQ9PLG35v7s59g/G8pdLEWQNCjWpf5ZTC
mHmI8dUZcvoYQWEpVYZUKOFAJSdPjR2ZT/wk2pG4DGZTAf5IC6t+ADJgumxI
+/dEDoRJzhM4JjszkOe7JtSoUIZqAac95/KJWMOKkRYTrHMh8IXyBSsK/60C
hxhufyFEoJIj0iO9SoSQuttwBoVXruJPrsyaHESvGzOZqKnu4qzXTwlTYWfX
3WOQVLTz0oMTwV1lEeKCGhDntOPolVvls2AyEpTRlFHytEMEnILEc0l7Ezui
mhHSWpHCbmOxLx9/Zffn46To5iNWRnJzL7JPxTk2iAJ213MOwM7QoUAV23ch
BwCKm55PdknSpHNo8vEBt3tRLuHSNZg8AoQ4nbPsDHZE/DD/HlfpmxbeJeq9
3E8+UOXVPrP/f+vzZ1x/q/XfEQ6ebeCRlhLqpXpY5PiWmI+SdB4AED1aQ5SL
p3/SKw51229rtWfw02zW3NSvSd6N0pBDu1/7RuGoxdxZcDOmqeAYnJJY+L0K
PDkxxskiGr9wJ4W31ZqyE3otwsuKbBKjkrfl6roz72t/7TEwNXytn/LqSnob
bH6Gv0IOkLEgjQd6IEya8Ng7D10IbnUGiKH/DjLwiwP6c55J33JU5lbzVuvc
UpfXZBxCtTvOiA9LprGLwzZflgWBcIJZFCJJgEgOwV08Wekg2UIJk6//gMt6
xhZUx4UME1LC664nLnz3qvfOdkJUIPWiXnMCoJGIy8Ei7y0gFM3wL4ulbFCq
pDmFy/ExoATwlcm82a67EkbnD1hTH99KViU4GkPJ/N8pFsIMScmNE1zGgsEQ
MMrtJNCY8jj4+F3et3fvDpMgXz4Tuu6fiNl8/heEw51FtPI4BBPXxyEWmiWQ
WToHgcWk1giUkvg7eaIUEYGtAexE/9ynje6f7JgHhmwtxgWoricDJXozf5fS
nlAZLZIKhiKYExQKUUX9JQ1Fa9VK2ezfAQdzuivd2MWOgmTgwgmO8XXKEx9J
tgmqTh7qfBNdJdMAt8CSl+2sk0XRB+XeNID07ceHrOzGv4MR2T24IWBDiX6m
MWtBtpUUvCdQv0E/FJU7ayNujaMBvt4CGQcjNGr8MhZxk8kZU3PFS43rZMSP
EpvsxiiIgPpfJNTLsnDKK6XADLufruOzSHL7+WU2aRIBe10zsYXOVUBl2YHF
Giijvv2hgJCRQ8zliL4RyEn0d177jGdv+LHiO97zfNyJCH4zETel6v+vitDu
6RjnZL38biMXSIixedMdka7j65Z6YrIg8bjhokLlljrTz6Vabjs03jWyfr71
jJvzyR7EkaJYdjWKshsSQcoPiwl21MH6K/pZPeg5W6kf0Nno4tC/xR8VjTtx
7pia94kWaOTsjFbp09Eggx16l6lQ7F/6rzAO4l3isWsjkcG0qsi/LKIfG+S5
bQ1pF6em73NUATNLJhV4N3ry8GmSd3SiXLJnYJGurqwFH2zzYNQXHA8XV7Xl
mr1UCRnU8M9uh+HH8Xw44UqPy7YDnh23pYLaQi+ie23FlwLzPXkHd2OVW/Vg
e84lW4oFbUBfdhVgo1HHBBAJuAXHWt7KCodXNj+cxONSZv45ULyqPDEWnxj1
zitf59yI43invYmj/FkZgnj0E78Wnx5GSPRwOpCd6bXHR8Ssl+ALKG/ZifGD
CNqrHTW9Tb5aJ/sEj20OHf2WDiCj9TqQcbm42ajcFtfYUR6UUDp+VaEppVhh
OahK8ZWC+aTYF44jKvKhNXZIwiGL7bvgCS3UGy2ZKgeEVeOGDIl+NXXx53dU
utmVHcbipjfB4g2UEjIjul0QrPS2yk5VOGbxGRcONfCv35kYPQBOEuz2umgs
gtqmoqOCdeo+5l0D6k0SE1FUWqcYr4KwfXcO4m1/RExsUPuGsmh9ZxLUKpaW
iSVAuoXr9GDU469beGdS9Dmc9XlKs0cMzw3mNwsKCPTb90ufrOU9sOo7PRJ3
20BddVd+ZZinLedlH+yvv0MjtG+qbtqjHl6SahwuG/2t8o2NIiZcKZYSFjgd
+49saS+Fz66Twyqs03nzk80mer1DB6P5oF4MIWD3G8h2H2wyp59qnWqHwga9
NTBwxvF9w7vZfj0a1J+csZ0ru0HeRnxA4bqZA1qjZOa1hHeYCASZkNnszKMz
lkw2XTo9lPwDZtvSpiHH9Wbhhit2P96pKNzKIY8qxro7o8evRjpfeKhLqcmh
DieHi9uZKK5IXLfbLukN3yHm7UHFGNXEYWCMXjBRprkX2PQDUfQ6GxT52L5R
jXI46B4YxyZwBDxFamGXJljUdqJepNSAnEaqBcl3Lp8uVZnJugi6QniSVkvH
3+Lp86tDTTE1KfXoIONvZVXHpQq5sBW3o9II3tMIRfT0RY53Kx5v427w4+ms
dQe1J9s0/4W1tkAiHuDgTwFHGiBlrdiT1VF5KLXfgpRrfWS699Z7RC4cjCMC
Dc4Z+R4Ng4er3/mEPwRqFvvRe91lWuAIlvV7GSF2BDGGhnN12gfw/jV0xdsB
cXtrC/hFd0gI9rTZ4Y9T2/YFI+gWTnl7axo2NRdpcyn57FcEiSDC1mTh0KGZ
QJ+LemUbJqQubhoTTApqMM/lHbjrdMhW6ky8SKv3te5k3dUifRS2u22Zbfde
8J5HqGHIGfRst9yWnshYNfAm2Py/fr6Dr/5LGnNOWTnWnCGKZ7+SCnr0cF7/
DQg/MBvtDu4k2BRLP6dOgb2mqQJ4+hrRSUP83gRcYaJWmLfKKEQtBsFwJW8b
NwpYl9hEFS/xQu5VPvIXVr4j8yRb1wdw1zViZR2PiPrgOxVxtpkhwFsKeTUi
ZIE7L8KbRbvMZvdKVD1zHolI9YFl4NbGnkljI6xmknJumktfc7ib84nDO42m
PQrUq99Vs8yQmYSqndwgNIpHv5+fWNqTgd6AACAgz06wSf1ng/BzwneDec/t
uyJ89VTQZlBy+KNW/RGvXPOznyNe+PZ+z5HKMiFgSnNgT8lMEPLEuR+69p9Z
27AFcXyjzB6Et3aOJcoEOxuVZ9ASWQTZhSn+1lrLaHNYkCQ4/122P4x31abz
VJov7G6vd0AGgdIMQEBHH9DQPKGwdVLmS3/C0tdT6ALKVRWN1VAEwEjjckwA
BgQULC3RtAn9GRceCut4d6/fB8igKsJ6nkkLuxnKh/U8GBlAPsJ2t8TthDQT
m9K8tJJfrysa703PNeCo3f2RfpRbXWBAJgDSsppD7WqUod667OePiqoLHB4O
3ARs6asvcR8TQEJ6L+yqmA3ka2RX9HEhFRcawX81igQ6f6vgsxka4gOfJqQE
rZwN1UUmgYku1MxATbHc6ZUWLFIjKtYH8WOVOTLiibY5BiK8ZU05DtG3tPkp
5TV7WRwC8sptlF1Mu/copOD8XoUVGKbrtjdUAFPBU1DwKR3BnDt5wu1O2eWG
yt5A8d/EiPfoHAnm9V7NAupkctZ6cxZF4+RJb562mkdEoRXV2ja6t01VQFDJ
kePteboMMNLnl0MDra+dDSWdweyM3DtIn/T4nZeg4NQFiD3Jvrcfxg2qxPkE
fikDJpMb8lhYfIFXz8fOJtprOWu96rPB9OQSHdw7UfWXQTTs3R2odgIN1V4C
r93w65BT8ZBZrNmMQ1abgmAD2jrvY5uoGvayYwxFIwDF3OcJMYdzipl2JaBj
jxxtcAP3oyzM2Zo0rAN+s2dd/NNnNRdZPPHvjh9edXukSmviU3lGTINoYx1b
6ZtE++v/1DRKDi17jbu0UrYggbM57B86+S+oZwLM4bKrskaig3owClIeUo3W
hrqktylatfAvJ6KiHTznScaIFX0adIlB2Y6oExQgT/6riOlYFJdEXiWZQ8qb
URRgVkCaoU8CrQvRQ/4cMCS6nkDPBpgx9gFn2gegnwY17glEtoY2K4vpVqoe
T1NvyUitZv6a+ow19XNVgRP49ZRQmu+za6r/cGgAzGg8eWJbGanLq2MFc+lG
0iPdldq0+VpCOtEvGGrnLIAxU9rtxTKrjUwEIq/A8UzM3s5e2FXQiO8tXhha
Y/AKL5L9OBSTzXMNEodB7OmQcnSo+PSBPxLqzeOxNHJmXSzqPHDb7VD+chR/
81TlqIc1ey1OB1cf6hRc38jFIoJee2X/xNH4aVuls1Q/SoRg7gHIOja6AyQq
dBV0EolaP93zsD2kItllNSF45tTnoDREJHh/abQHXTNEyHms/TDAw7BFp44D
Yw1PbL04FhxieR74QxCrUvRnhnINl+yJvpXnZcr3qpDMcoj9kKBO7t68UeWM
DbFrbfmlogjuoITFyi/ega1ZondzS+RUtLz8bqeANyltya5j6J4EGQHvdlXI
1kG8PpeC0hn8q/EegAem6sjoS0BmRMDOtOvvn4b6RA/rauEF3MBGawysULNv
OmvZ517OMfSAtABhXvW7btcEJHN0S/ty9NU0q6XD9FQcYC3zdQTg3lq+rw9n
0aBCMdoYbCKQRB8J7GnUl2sPHnRcIOU2E5A2FwW5Kpm55YwdNYV6x6b45slw
42GSmJvFNomQ649ZTJJ5k9g5xrENAQH2cJoAkvjtyvwCAnOBgm03mpDTWLUD
flPS3xQA3az8vIeW7TVWIamRGNJ1MHIaLh8vVQvnFv//ga38PMlFOyZNBuLk
UmilCZzpZsZNE8WHPwJSh3OT6M57WY1es2dcBEZhwdusriL7dO4rXp+tOqWs
ICr2sZuoTM4U4qJZCw4hjEP8Sbm9hB4ITR1yAIJf/VBuRPYKS5BLLabNqq+r
M8Opr2HxHTnIYwSkhbAWBGyNEBVdJdq3MiRbgK9/gMamM+WLh9D+AtjJltYP
XIzXmMMut2QsDx/lRffj6BULsLoSl3RSJl0EB396mDLxr+/X0mphrXJc8Px0
lsQU3KcOpw7WzGUzqfHd3neX681qijhZ8MZ+fIqultoUurXEwNjXwu/sV8K9
MtqA/qKHxFqV47BQ43y3GzrfTFTjxOH/Ezt+wbgPb5c6mw1Mbqy8o0jhBP4p
r6btJZwzzRHb1MADxc4njLsmGUsWZzRC1bk4H1BcwqNe+xEEyro3fgJvf6FU
jFFBkZyP7mgnHhr24DRybvCHfIaPzcbtTsG6tax2Y0VrHN8lAeXVKxFtzu82
luk+uE4c7hy7LgTAN1RT78qolWo0xogbz/V9Uua4Zj2sV1BSXt16ZoeF/IZ0
oWPeeKjAe4FJntN7PIwJQdiJwXAGSrl8ELpd02Qfppkd4wE5uvNO+zWqS3f9
6qLzUnis2aaBdUbxnr6YrYc9yf9823Cr29krbgEvz2YNqbSfDfQWTlPJUXkb
p91NF9hi4YKGiKUsVl93lbtxzJpFcpKo8wym+UjIQWpmgTe0NaVBRkdWYuWc
q9SlT5ymE2QJGL7kOGU2a42Hpp5GixrwEVhCvT8tCjaIICqrJB+e+wCUduQQ
01V1myYGsO3jCzixicw9T9RriYJZkFQc39wOn+NnP6PlbAlqttm0pV0zInWi
oomTm983p8XJOXyZpbNy81XAM9VHXhujHqfzA9eCImLUlE+EJZxyT3NUq3jM
K3OuHaFRu0mV0fJBFeB0NZkNO9FbDiClnez0YAc0toWqIau8ziT0tdVNFvYL
uheds48dJOf4hSUEolnu+E77xQZwbI1BdZPbnHNQOnLADvEA5iy8DS0xUPVd
ebKXVmuwZkCDSiVy9W3MxDpANRov7qUYS9zAziPz5W9OLGnTtDMl3YOIfTSz
7cjCp5GFaCnCK88KsqMiodDgVg0DrPLu6eR6kuG29+LBEoYoNPSSHiBnNxsE
GpmCeDnquGmgKfRLvcNSUS7HO0jUlB0OdKN4Jk/JkYuiTf555FBWoRAhI4QO
nfZaMSUjVxohrAXxfF2Q3yQz8BUOujKuFUuK7oadrf6JNGuTtuSTcfdq1uxc
j5Lp7D++RZ6vzTgViH46YgpdS4Qdvbdv21kTL01k/ko6KVdAKt+RFRY6X4fi
OHd+99SnkMQ8eGvVqtUTazlm58kRZmfQEOuqSNLJnk34CZLpNClUTTGMqRXi
dz6gfciEKpbHvk3PKlQfUCElThfK8TpAzELJNYgkHpcBE3/1dlVktjmCdmnE
1m5RpTQ4CRlAoQBNraxVvU78qWQaY9CVi5XRCdMqo+wanTriGR6E4GyTtVVf
0oScORx5h/5BpGrPOCQzjW3U6DX2PfCueKJeVbCqYsySBP430KBwvDE21CC3
PbjiG4g2LXoFnnMqr7UPD6J67ZWhKQz4Hjo74oyTgmaW87w7JU1qBJNQm3Wq
bZknsTg54nKOZGCdet9jVI55zJxP6nRMaK907ETTGYL8aOpC6F2D4w8T9vuv
Ob2y836+H39QOOJLyI7gsTQlzuPR8tKEqNEtn4MhzUKZtWpq3IoAkNHzPUTJ
cehY7KRFq64nubrLP1+Wj6/uKWVp/L9h48oa82hqhpe3yx9LeSPDvtGiWJY8
1//zIOdLdh+8zT1vGor5YzL0LrVmWlJMrxGvl68a6hCMgTqE/tVBkdE3cfTV
skLyA197PZAfxtVI3EiLLjeILD5IAOc8ch9z+r/T0dof6CrCZJnlXM83oE1R
c7KPJzkBzq3w22o5oe4gBF9xDpNCEYZ/lK3RA9zamrJIsyD90txclMU/HSlA
t8p5MXBs9LULXPORJLS1cF97VqyRh3TyZZyqy/buBZW/pTKV80S+78ZhQeSm
NSkqddhmduXAV5qTSlx+XVHcnLctqW/5+D9Ub6hKXnznvcbC96xL/inB5QV3
CKRxZucxi5quXIsikChFRF97UA2Xu1/8E6dYpuSAO8b7WHUJfFst3ekp+Rwe
5SUhrXhnFylyp7rEgibLNCWFn63SMMnfT3BslbG1/liXzZsjmZ1DDF1sjbWM
CaVQUk3SuPSW6uZdqXs2tYUCjxe+elztt/rvbNxCStPOz/NVEtA1ghtlx5BS
K96zilbh5WIDzBQaq8HzPGsnnSBppbog0oaek3uKLuWYS3t2zwcRwLG561Bu
hXs1GrbMBq+nNjN7tPeyITmEDJmqjX5YHi5X2AZKEMIIxZLJSuIuTgsuFfCl
Y/8zqbYdTm/6qSTYaOustHgC2HcZCq8+Ba8MM3ZCjoWPISDjcyti72ZjkxC2
0FC+T94L6d5n5qVqPo3009YJpzV39ZpSUgYPTBzmR2aKfOebzbWh2yrY3a/M
nSmvrPR11GHvS05K6BwBLbStS1beAsthxx0s9W61SI0bx6QYXn44N1cV8jDA
0zt9+r3KKiWyYyPb1nO7FxF6hS14+z+21DctTa5Du/uURRLIP3bxQ6Bj8bxO
+Bvgh5YCb3a1dtOxEGk6eZLutdurF2OIgbQ4IFzx4U9R/ebuIrNcuAnieitX
lugTxeR4cm4ftGp2YViUuxAQRkSRZfNnaznmztAAUErYGDdwHclEnmCsBoAh
N5LgAbSSyd5sW6GDeYPhI7im6UeY1vRDwxqLCY+m5cgnrscK1eEfQfeCeCG8
ADtmUSa9AV9YAJAfgbtVBrx3m1Seka4ijG22jjAnNCM1qASDMP9P8dUuITHj
4B1pqJh/7knrDJKupDuRXEqK5ZjzcGoYYFRzWOlBqskRQBBsC9uHml8zM+Eg
tw3Z/bWT2A65aiL5v36J0WjdyJJTT+sEMNLR2XT5RrHLWH7JRNSFDiXKkaVn
MoCXKyVWfGm2aBqtdokSumkMVYuOzU21ajpSf+oYx4vlKnaTsk++8Rar/wDV
lE3gLlIvJfxnIQLfJKNSzAnUbB9jlvoYHZn5u3ZHz1owi8dwDz/oUsM8j2lR
KWkZEYdUpOPkshu0Ls8GWGDGbnaKdsudF43/a/mstULRu3aaOKTTBcdtcmoJ
IrSM+rJWwVsE6zULb1/SYqVeX9VwhTK5vHFaOGchfMVoasidYhaWYVtgbUTW
YMJWT4yUZnSdaTjlc3/IYzLqTdwO9QyNx5MVmmsTxspSFHJnbuZptIYyDF/f
trV9e0KfgE06t+QPcdh7XkLSNTkMJ8nFKjL6pY71kuf+Ux/92kbhGSWnZ9+b
dmtSZY3KYldupHeBS1p6DDQZaKTWaQpkv7tBB5f5bg6Ozj79kvzYFBgU8KUk
36VAj0CXk1K+neBtf5MEIc7RSuZBiXBwH2D5qsWl9/OATyXEIFXn1JUzspmt
BGtu6TTl1GHNZgzmlkc+sfwJe6MEftq6gf7HR0HVWcae+AVhw2xbbZsfZKPN
Svf+Cwk1bzzvGyiZIT/x8vlx58uL7eGfd0xjYG2aTELwtFx4YkXyGXc2eiUC
oUs/V9v/9EZn2dNxTa+0wkV5gNS7MLCBvw1VYrfZMZt4JwG6z3q4ljeMRFSI
5imlRUJ7YBTriANPva23C4++DmShgUO4YSEEs6Pg2YKz+dgJIrD/zjhlv04l
vnbUkU32OAOTvzAVfSND678unDVfQbDtm+rk8Lq0vk3Qrp0RWuqyC1ECEdWE
nPYqPkjtxyaIcQZB+/qPeBqo1ZPxhv3Jo7QQwndY3B7vgsCXzW1NlO9020Xm
ZH8YJz3XuAmnBwVerD9NUXJ8i1jacH6RG4UGZI93Vml955NkrjCU6hmQ+xlO
wE3KVO69ZbMFCupCY37soH1AmEtiHnPH0HC07P4iNdTJ9uQ/JfwMxPdzFXWI
A6cM7THwzqUYvKJK3PUISE6o4jExF5lrrkDX4lnaqKQYA3LdbKaWRcp7oBPD
SeNhHKF2yXA7eEv5HOlNP6i0geVIvIeLKP+xwElsRRLvIXTHjTv8h1e4FTbf
NRwGfQ1OonwZLYamKzhKyVURg5xHGBOUfOsCE2ldm6lyYW/tGzM60sb8L+sV
r5PMPtEPPJnIg0q7SUEiiYJX+Z7h8rlF/+nbBCwFpW2LDvArytjHLS4hQhzZ
Qp1a9chi9eguKfl35Rh28U/NoPNO3cTHVa3J4bJ2bfx0xggRc8x5zs0xqXbY
qf9mJCIYvbOtYfDPcr1JRriKUL35U76A0DYKZDiR3kcOPkzUJdQRAxqkzElC
iYL7YXFa28tTSybihA6dt1t1I4PPXAThBh95jjCWefggJI26DbncA7Us4LQj
RbtO0Bb+Jut8k2/fMkWkpSsh3wgO+ER0mE+tgZzhlYBytJEVy3kLC3RQ18Vf
dudNOgjKgDlnWDnaVU49jYAtoPhu6pZRUDpuWDpw+RLs1ZesMAkueC+c1S/b
/2utd1aQq918rhn63cbHWDD9zFWn4k4fAb26ySSaLFqDBkbrZJWcRoFjTTx9
RJjearx6aclLCfGD/EN7GZh4CtpTglauP/GDtgnkrMdRMyKiWihP2J+DAB2Z
cKTgZFYYpWkGj1qUwqawKQmuJA3+vkU7axeBNXgmaXgg6Oq5+C4cQRfz28Av
PFqH5Bkh1Fxw7uLygsNliGUQovjhtUlXgTU3e7IeAU/K8Rm3S/fXypvqB0Va
6hz8qTgY5aP93av76/FCzdD9JDQKnQRASXBhw52PDWzfu7kmdXYfIAFi4yEX
4HPOSGEqVxnoYoXVqGyP4ysyttT9w8uNr26Qz77fOepDbPoF/Nddt4SY8Ze8
+4oDbPiMJupAJJhJGxT6R/tbeCF+tQUoAwn/55ggM2d232YgkmshIgcaIax9
vAABBzl5uZCuaJq8j+jABhbdtquO2wukQz5017OeULaxFbVnoB2yl/Hzspw0
0OihhzA1NUDdXzR73AR9lZqr7bnKUxn5dV8A/kQftPORA7tGWFwsx3MvZTkc
Hacl6Li78WY8PB0Pc2w2FCUy9TnzXPAqhqLKs0Cw+gmROV2rbLEJyAIfVFi2
WZ2bfXzB+cma4/Rwjeo/dSI00PEpeQppqjmCJSVxt+ULoE/VaVTgqEEeUyy2
HyhMOE0G4BybZ4LEijnLHV9vAwdtgtiE+P78J/7KQzQvsqUBgec6/8cLw9i1
sExgCcVXBQ9IZJtKjOBcoN5f+TUeqdakzxRKeOvX/jdCm1jxwOSOXc+vxjZe
5w7N07w/777OjOLoMXjk6CQD/UxUxedK/81kMSsdnETuEPf8wOgUpzGKYavr
5Q90csNKs5lU7YCYlV5CGmhlUq1GLjeKEpCACYVzmnVGBXe0j6WUG+MB39Sn
d1Fe2eJIHebv36j2xGGTK207cSByVKDddjGUSOPV/CtDaN4BV5k/g/IKroIi
e0eerC5YpBSXZNi63EfLGI40Q72pnFnEt/B/gRQgh9NIwrQJ9fBXnWGYvg4+
Q0pqourLoyv0NFfFvbFKPtWvVA3uVtIlR1bm7O3pPDAyG+CHFOtKOp37Bg/8
Eh3DLXkgp2lRkf8ugfAmfQljkqfS2vBaqWgt8jbtlwYy7pOo8h+VGZxTJ5fc
opkpI+tSjeDGzXX8IaI6XKRzd3TfpnPs+eEt2JbRNo57kmYhgtnOwysXGU0D
gk/VDBEzDr1uEMvmudFKUkfzKDv0qthzA6IQf3FDhkerA9JgbmRfsiCbi3Q0
OPCOl3h0cSSIv8KkbXOtfSzwp7W5H7NXkS8R2mNKCbUJKy6oydVxjdEixbgC
8cVXR1vE8kdF/siX2L9mOdXtHKtK7xXt/6B3XAXBU7TzLPN23Jy/Dd7OutBd
NxVKH77ZGurCm1tlYVa+/Qs108ngB6tNc2PlCrfjgV9Vl2RK7EYW2p6zFUPH
jIFHkT4Bu152pOtmRiQY6L+8P9IVt8SWd18sOmjlLCp1le/QwDe0kKLYhgD8
AsMFzEKULMO6Z9nySTvmlQZSY/kKzIl/EVaZez1aHOe2Qepaf4COh30pmz2c
9W+k7hiWa2lT4FjbyQxO8PUOybqXV0me/UQHtM+AZuqGOvwk+kD5pGwi3qUL
SGHutZUpNwMJ0UzKVsxYWUmEPNBfgF0lq2PeFZHfeKAdBvn+bAkSVTDTqofP
WJGihlD+QkXGnX46+snA/yNYQssEr/CCoXFCILsSeHUENmVIZy7qTcB5WbLh
HuG6zyY/KPZRHXSGqdT84vDlo8c60dUrlA5tGCpM9yKoW63YisYvM9bciKX7
uYx9f52jCiXOC6QtQJaph3ZLvBPIV8N44s4tZNd3+T0SXjwZ+oQr0CI5Jw/P
Bzz4hnGicbH1WqGpuZHs06uy2yg3YGbxbZGX76/eF+pxy42XcL38J/Wg5Ndh
/tvQV3EI/ywEcte7evfKnDplJw/l1eWSSfhUbJicLJqbPE+/tY+bs/yAdo9U
3KdnlBqKQgHxd2ONY14Uq9sroEhRLjoisD59tHTERopiaGcNEbEbnvV6O3Fx
6iJ63pZXI9c1lf6+u7mmJJ698q/rwA69IvEiaUCqqN+L4TUmUehVbZ8+Do7K
Z8O+SRXGHS0M6CgjWn5gP1sJ27e+TMbdVpuZuULBoBILeG+5fy9rvYhYmgno
eUN4hD4KAQ76n71y5OuOQFLsdfjPRu8or/yv7o2RT+IgmZdTE0aZ8T/4W1fB
31d0htTz576BuD5objVQipHpHL+nVGZqNtrQ+SRGJ6YYP2+UQLAYzMUK3Ps8
7Q2mXWoSTFWvEcoWd/Ge04sippxKWo4l0flkajeUs3SLxpTrkrb468le4SMh
4XDACVhQYw+O3fLEccdfRvyy68C0T+VfgXUi1v0h/0WNDO6w6fAoySUIZcEX
W3ypbZCyxOJvId2xkbnN3mXbmv1pnZ8f1R24EhrxcNaIPlfGgICV7TbYlgLz
95Y3n9eNNEyiRoa2Rd4lPVQSw/XEmNdJ00ZUaakAAW5D1cNFdGW8zLTJ6W87
Ojmc7J6PMV8q8c1EG8gxwXH6VA9jaipMvqFTbC5Rhjps0NwUPQpCgwDlNhxc
El+IIVQZzl+85BQfAZOPMIOxg1PAKJtBMOvnbf51jYLhoZGEfbfvHymROljT
lghLCBXQimi51d4ViEPrgFF3I5ydkpa5Ai5CtXN3JJ2DgcCHE46lLMy/LnuZ
YcN1N+9lmGwLzvEprwXxKtWDAC3KnWqLkzqRj6Zh3U1lZc3ryMoN3KdhVjEd
GkzapgOLYGSRA956uovFyrjmBMIvCXETFOYDSGO0oQrANR3RSp5Hu/pwCwlf
spZool3yxnrc8aY9OkHxogSWTewYN104DhZuW/atPSgzQXirUOaI9qCIEl9a
TB592fn4kE8tYwUQeEOx30aER8CDhQFn/fwPyKT97ruEEb8GRG44RLJ2E0Cc
bGPhVKlVKHSBox/dRSnPnagwbiJJg972Mwgi0oLQN93cNN+kApFIxZ3sBVmL
g7Tw9D32TdsA04wMpKMg9i8RBo4lEEVSHywRDXGKQhak7pSS8tjTjnONZ6kM
YThstM1qH28sdiRI1IqlqUgTqzcMEiIv75z4LBzIGIC7bs+2XfSXBvfylgIb
ceGUfxVZs6NHqHsTU9yHzhd7qqYFrqX06uuo67lFWxYlihpAKqg6XK0RA2Hm
tSpOQaFNJSisv7YiNVBwmKFwWhkG2qp8mknlq6GY2IHLGEIQ0+McQ+XPDmMK
PWD4qMgB3bygjfcgLrwprE87dGNtyOpWXzWUIgkDQx5nMzJ9r6NHl8uiruPp
9Ov6pdOb6JUCkGUhRJZGqbj337RxH7o+ejaJdr4I5rhaJeuaXE28sVa6lcxO
7sjQtcE2BaBk3QmDTHmZYcwZ03ReILfDzmxLbpjBhCNHa56OgKGiq2cZ++5+
vE4W6SYNjm5luIzfQcNwNwXuwunIqkRS6XJKsVhdDfuuCR19k/FmVKJdWKn2
ZgwBRDtztZybOU5d9wW1mcCWSJ5vViYh2wzaD7GhLqZlqo6XnKY7LS8TK1K0
4YV7s2Y42DqtOhUWlmZkzhWonBYjQyTIrwwUY85r9xukEtATjdgVN3p24aeU
fHxCiFHlfBjHfp5eZlsha/tuWaVBWqAxsPwDmwWTTwdDXFtBfFK0tJAGLPnx
qtaC+LXWsHMy6eqrlsS21TX5f4uI84vMeayQhqUAWWzW+bBMRV9C2D6VAro3
gWHpuiXUJgjgqr+4WkFD+vScEid2IRYTKMGwj8Bu0B0njB7JtFFrS8uSOsA3
I/s1VX+H4dAK1Y1vg36oceI87w6vI4urxKBEll3OpfVG49a4P9LHAJoiZQTI
hRnT1OdsnQYQ0C/cTVF4Zsb8rC0x5tBYPTlpuONd4j2LQMcAsUK9Yc9CxXUv
RQWX0H7IHNTfmNYEwaQavAGuYuVb9HqtoPzrcdiGtDVPm1aXmxvbGsecQJwr
2xmqvC81pDlrtx+Fok9L4wZkw3J/gZx7HHhQdDzcS3zBCyJ+I6RU5oEZ5wT8
36XkRYsqhlbqHYeJgq19BJnNc29nrMR3DRaj2b9NHQgD+OVAk/cn6b7+RYoP
v5rf7htoZlvohDkstLaxhl7rOLMyNBT/NfLoToVk8pRzisto2FaUvmgZLZbD
Z2ruJozoyElNSQnx93YeTm+QEftCKdd0FvoaSjRVKPRIzqesJGnhcn7Adq3a
/QAcFB4mkVoNeWUmUviCH+eStQhU9WaOMePw7FBvihuf7sna39C+LqVoBHMN
ih67rjWUmCbfDtbezsgGGDe3fE0KgBznc0Nyk1xJ75FTarDY9BSjDKK3nznk
NvrFOEPaIqPB4LSSNPKVpxbg5o+94o6WE/0UuLFGiQ6VvbtbPrcbNNZyyjla
Z4V5kACfQB5WiAV19d5f2sf/UiTwmJ/JeIosKpmnl/K3SJJRITmHaECsoyTD
+KmE6jGr8+4KoG+HH2RGm95tAwJabRCr0LiBm5Tb73ks6CjgmJLS/OCUeFh8
IIoYAjPv0J7pDXmOSFBYI4cTwIOkTG+RGpPEd4QFQLD1VptX1jNMSKLlt9+S
ejS+HXeT1B6FcfXsKAvT6NSzSsBL/4lef4sQ2Lgiu7Qamuvpw3KQHntDMXp9
9Mu81Dvkqm8EPvj6UAC3nUClpQzJ9gZUiqy4rJAD92MJa4/k9dgNIdEgkBeq
7OdAmw7QgYoMS6x/20cEyFXWpBWRkkPIsrW/UyS0m21Cjn5JgtR2MRNz6D4F
9kBDhozUNRG6N4fBxLl521rmfiV2fkP2pN6Jsqf+aCM3UnT53YY6BAga4b8h
Z87npw88mWSZsDz+tj0ao2iP3xGCF3nqf0jLUEq4Zdqug9//jXkr32Ql5hez
LJRbM2jtCMirRLRQIgqHwk/tgSmwGWOASlAzgM8tbD2WrI4/8s7R65LaVLHf
xccAxWsELmLZ0ZkGss3SKDFUdK7dWCq8jW2oqShraRp//t++dMfUw43lIi5O
EOEWrwjTDQJ9JoIu1K/nP3ON84clsPN9OgWR8M0XLcsLBU5avuu6VMVpGBs0
LCzznVLy5NKGNr9Kq/MbWph/X87ExVEnPWYFij6QdIVlBEWBB8gyFLEya05E
o3t/RRpO0ZkCo5Sq9pKW4R6S0FXAivTq/g5R0FACvwuuSqN9C530iJ8dk7gi
dMijEukx3My7C+e9iWyuaB57kU8s2NpVA/QU31sEncJFhyqNS6ffDWvUpBGh
dOECJ+dSqCRes52DdAPYvfCM+E91++r0ZuayWFOy70pBzvt98VjEGdK6lT+n
z9u0kp4Ff4n4J+/hi9CkMrY7Nnr1db1mOzD6+FDYdnISIyB2EWDrkXA3ZAf+
NFNWbdr79Oer68nn6028+TsIgbhj3AHQnc++aB0yJh4wohHlsnSNF/iOJW3v
3ZqOr+YHrOnzhJIdm0wlrY4sE01Pu2g0PaIv3D3l8stvK3HPWiDEQ92VFFT2
jLRNkELpwSwcbdYMM/YjgZZNdN9uqdPBo4AbxW+HtdAKOtpN/TKhblhVWdpn
j6R4L1pKS9X3G/pArTK0LsfkOd38p7TOIE3O2qhnvh75/jkX9gWMyEwn3RI7
3qZaqG2bzLSyS9GIsYf+/IxytgU8gjNOwSRPz4j1KGWgv9aYiECrFiMte8b2
07AUT6dQdqTdhjsP2FRpQyzd+wkhWU4xZmy2SW9cItuUzNZSudPf1gMGsb0j
ITmBf1BkGVVHGffvdOwNyzeOPlgsBIxKcLqkhxIopsle42kTr/GUcEaxcFbH
TVi6ToSSgv6nPb+8ahP+DyU5Que4zgZPeAbi3jyih29RmQ0nQuGHgeYGXaV7
O+KsRB/FUQF1776ZPI9ffq+dZUoqpCNoVqdE2bxDMrQdGMnIFPEOaxwz2rcM
RWwavAfsawpv+L6TlPaMOF4iXUHJrVArjHNtvZF+WaSJ1T0fAB/vl5ZyBV+G
odFt4lecSQD90VYIpmnadKcfaEIIII4LKRvcOzHs2X/0/IFga+2OrKBAvg32
G3xel2SD3ETvjqtNwyu6U9rJwl8arxvXhrGKK222zIdUBRs0x8pDi5B1WYGO
fV+Z/2I/g42k+fd1bstSGWPvJVrBRhc1SpWxSYhIvW0ftuqTZm+kV5svWpFG
iKYZjNr+S93mrCf9879vmww2hcRLGTrUkLNibqeWY2rwoo2lv1Zmcu46KxSL
yyRBjgKMFs86IsItwbfKf81AA/J8uW3kUMyrWDOABixy0yAuw+VZVgcXsbvs
4lDoDC0QcXzyVvffHsCeLowPLhmJoCA4E98QXbF7yinKNi9cYNLgq1I6ECOd
zj6LguLG1klQWCKgQBKFxMDR9hlsfm+hZ6WSy+IVe+LxqAxA/l4+DFz3zB7h
IBmgkqbJ4JipiYy65qjllCG+hoNdHX2izNwRApXwvCvVh8BjWUjdoz1p81sJ
Fh80kmSxX9Mv+zy0fa/j2a3XteDmQGDQUPPWUIsarfLJrfgtxpK3Xh52U5Mb
A3/joXHVJPg3mUAfxUECmqw7pUfbTN8Tx/cu667pqgmErwS0zqAEnMYasEp+
6Xt8ujwsOcFPA9FSAYb8ZYMTUQ+tE0YHsDD1pDBAiZTZem02TMtGKxlo5lA8
5WfK4xiwd/JB8Co+uH4rSY6luI5VoqBlzawUvds3IQtoYy4rCeiSKy6kEYzI
Dlhmqk8p6M+mwwmKAK50llHe4uUl6rCz0qDns4hnBcaoCIzmL+R4yLRDuE91
vj9RtPHn3B/n9IFj58RAcRBnh4YAtXMYfa4NE78h1JJCGxF0fwbC9wWoKsmT
Fb0k2px2POQonBMN7EExA7RddyD3LO3FPA/RGoa3ZCf4Pa/AhpZKGB0mMOGv
IhS2dBNV2sP6jDz8zNuaW/AMZ6dQ3dbAvZV4sHvNvwLaqC6q4awROXYvzXV7
WuWBfDYUEM7UaNdQhl7x4B+RUce8bUYWw+GBVl2HZt8vOh4vT5QGmgYQXrmA
AqAOMuPDkEezZ1e5ey/o/DPMtFvv9Yg0ydVcOFPY/IlRZDPcRSbT+4CzQ43U
ZMPXaLqhl5VT2TcCqEg2sR0PP2R0cRY1rPqczIX0N7z4klTqz3QcLdcX9zyD
jtbop1mdIrHh5HvhnP45qhX/Rshl08fGe8bklF6Tvuwy3qaJMYUL0it0YWhX
8IX4mRLwrt5QGkGk24yTGZjs3f9ydRlNOv2UbEc3hs6iKp1KGE7XlfMLZHbS
gP+BuLbBrfATK7TcfLCjllFVmsrn476SYpTeL5oWo8SqiM/ixgVE2LnLUMNz
FklPPeyZ9+JVar58y94YGxFN4/QJ95E9eXQY5DswQQbn6VpvjSSu8i0S0D/B
m1jEZp56wnIuhpbydWHuqJtkt4UNI6Q4qu4oVjPVFmW8yN0hU3mv1rCk78tl
GYmyo68PYwnoScjxSVkheJb0R+mrULdzPKuP9ZTV4xpdgvz4kKK1sQBbLEQZ
gclnLvtii7hzmfkaBZiX902T0E6L5FzYZq9FGZvx3XtpdsR3rRCGRLGoSD+M
vXd9C6VVh5eQcJHaP+jHjTlmh5YjdeCeRXZaA1IoOrO+8IOZA2bgsszLIKdM
DoKG0KDQlOEUFZm8Qmxkwiopga41OID9/FKaDsi2Q7BRGGifu+7ngqUcc6O+
oN3sklwQUYkD9L7HyL0cH3ETxf3sZM/ALOGV2jU+6nJ8zbcYGQ8rZJ1Y3uJH
hw07wEQy2LIhlaLP/vsRG3xzWzWMz4srj3Lz30vcxXfYGQITKtV00Prue1Oc
RW3udUDFd3XLDTydSHCGcOkJlM1XmFJCoAggYFValWvxoRGbmM4Kxkp4hq12
3MwesTdz6U6NbEAcVMhrjzZHfBsG0nF+Q/77oeLgSFR0F4yxXqBKqPDraq8X
l61R2PM6OgBE4fo2QEeoUZr/C4i0mNDyt6ZZRsPyZN6w+1f0EPW54uqUgMWL
TiJZMsAH6z5i9/PRbIlFqsTjTbDpqOCulvw3767t9v+pPBWPQjKacGZMnK1M
DawO5hb1uT4iHNr/LsVR0dLYMpiFmWX6gjRKPxuG7krcYSsQ3vaKr9kl+Zh9
IEj+qSCeHofaegjWslJlY/C9hD7dssNbug0ufKMYSlRLSff4vV+tsUlg/Va6
XhntXKexv1m4yjJ5eSFmYvVrNAYEeZo5zcThAgnCv391iBE6SZYtGb2fEE3g
z27siEWebYa6U8TW544xhmCp0PuMXSd+WiveXOVKS9vHXh1JMSKoQ53/iFt1
QCDH/9XJcdAGOA5lNfw01gc5LZHMIzBQB70G1th6BDKM1m9aQnvDvYipcKkQ
i+XVQP0ijLzcmaSOnOUjF+K6GukPNNiFJQvcvZPSFbs1W/1mliltE1Xkdmdd
PYnTVrnxYrdt8AwENwrmQ2LOT+JGg6f9eVbweICphTNe76rw508RZvQsdQm3
NT7EcSfLJEqRGuHo9E6a/5kZozj69QQwAkdP8+NdA22qmeQIfa+ZefKrAqqj
3eeQ5jKCPgfx8nYTqeDfv/+hzOUEpRNkWXaUfTnASSgfPX24fPS00rsHwwdk
FT2shtRdirhsE/eqCZiz4zY3OfawI4ObnVT679lriZ4RpWwjYPBll+6A7lW1
wAP9DPC69UPoKnZlK0ehZ7K64a7w08N6mO8s4bjwEMgnl7knVAmaWyPiyP9g
UZVjBrW/t6Z0K9klB4Do/R2S/hLcDQpwO9KtSwu9YQzjxOyzCFStPkFHzM8M
cCpesTabms7Z+pMGBfC37Lt2li16S93uYoeW0T8jnCaq/aTYU3zYpCQamook
YfnDrwDEAVf5q93OFHweFCo6Tcdakr5KIe/q/7Pg0GN29J6hirVNXT8WFguk
DjtRmdDPSTalVr4WIfstuixtgbZpwKe6h0uJpdyUl0jbUbsOMbbvekkIKmdz
7IjDcQ5B+YwEHnTZEbHuhTgdGPLQ0/8u0RHsx0eeWkVkgUvbUf3q49e8LoGe
YzVD1yy69VfCQP2qHQaiKZP6m6V60NcPMyQGlCtnjNzgOrrRX9RVPLZl6kJm
NKPgKrADJGB9jZnZvKr4OZQc82tBs7tQUHKWtoIC+9UHmZFBS6idPeM334To
ZjMo6YPz+jnNm/rE8SxaWj7tZyQGeFO+DvFY8G6a5oqXepfQOUsCMLQjZuIS
69cygWFTsQSdTq4LDXvcxiXdoscOXd3jumsiVoHGHzEQHXnZsToZlxpGzmt7
Y3Zj2nxtc8qT6Lro0pUhrj53K3eC340xDcHqyxXHqh/udKe08GR9CigQsaZs
r4WDUft4lGEx/xH22cJL6vu44suTMH4hQNJPEiOl28pc3bY4c3uFWHtDZJTc
/AenqwPknA7+5AmTKBfVe7Mo3O7VOomkOlmQpYuXWklSCY4mXelH85JFo2qU
rVP5mpSjZ1FZUtdTVtHJ8d4OmaHaxLJ1ImtwFXT+84wiO7G9BYOgQt0Uayjv
IpuyPb00FaeC6kg82jS7SYUqmcrcl4jX2Z+McOT2rtv5YbO6KPX+qBF1qlVD
9aYS7P5rsX7b4oql4DDI82Fv3rx8iss2wcxCzd2K0mvxY5wvW3FcxHAU52WP
abhQnex4S3wy7gTDNVYs1dlx537/WdFXB6BuVmj14EYEyOT7yXojUXpcZGGu
nq8Oh3AWEpNlSpyOUcAzJ8moqHFMVDR7gyNWgG1GUE5fGxDz1+O1Qj9ES+sL
2uDIZfhQpNxB460m7BCU9TX58ZWmFCPFoFm18S5BbHnJAcIHGkN0N/vOqsH9
hhK04ezKrP/jurixV13OLUUhl6VOT/FgUu/tBVJczAY8XzMmMfOEOJkr1Mq8
30PUqUyy69AtjQhn9fxB3cOaLs99fYz/JPqEUGoa8sCjOXwHTvtNOp9lqRq6
1zZqVRMELTqR/+l+WiFyNLwPNxd6A41KBjzYZSfdfLaQeNSIejZHpz8RlhIN
b6G3qCL/pRJzPZolAMJTq2H00NAbs52WC+8iLlxH4ccPKkk4neq+BB2BseAM
YTCwaaHcpgzgQ7IlOS+xnCqxnMD7DB6GkVRZviE5cFvei7VVoCVBdX/TPUjN
oD78Xez166B8GD+DEwwQrX1uBN7PwyOPbK1NZijveF231Jf7uW1g367sux1D
KAOE0NP2iuqWzKrfvn7LkffjPHY/mVB29+Myty6ukPiUGtRmkJiYqB/96rez
esZsFzfRXJqodomr2tfy9S7R9d3gnAH/t4zSHX5ZEhOP2KxMGq7LkZxH9XOm
wqme+vtV+c7S0IDcSiW6MURe9nJxDjz87ch3M0dgrCJ1f0cCKyWHwpE8qKtZ
XRsTH+wOVB8YKts0SzUiaYi0EQiy9flqYZJFrA2DcHWt1gd3YSG23LtO9Bkx
aJNqWir6IiKuGFEyFNOWVrtariWJlQihqBh3MoYvAcJdYBBqQWnb8qERbANJ
dv1KQ42U4QamrcWcfbAcmRPN8FnlMNIUc0Mnter2nsCLJkhKopzDf8KX0wxa
i29Jch99rl3UltV1Ie/sMRCkY5UchdKoccldZcbLy/jCYbIfv4bF3J13w1fy
PUXgITJIIkYglrh2Kkxl6Neb8gTvq80DRXgm30ri3Oatc/09941Ol85YIcjx
ib93A/5PHpoSWl3A8dv5hDnNXINTp2vftUuR1/jGhnPEkh3tp6/dI4BNNRRk
agX4VbD2X8JzRld8HYzEGw4+HbE9E4WB/3/ehc3etjRFuOWppA4S5cdgxoMC
YZ9W9Nca3cfT1QigBE845DuW/9eoKFGpQqjvFF5JOTtqorMfKXUEQglpCcIw
erbOefAcgEaXjOdYx28hb7dR2J7lnkBrnJxgj0u1waLotjq5tFViu4ImybZI
IJMvaG7r018LSUj5GJl9EZjTDKFiPbJuMsDd1FW6RjY6ZLZhGZ5pT8zA1Qjh
qO8q4XBUV3p64FaqiNjwJ9edR+TVpRoy3L5YLs0ty6lIQZN0r75Bk4trc36I
drRdoOBOHJRSovcGt/wNTh/z2fJOuJWBseqwT51wlG8YW1qGorZsgW+nP4T5
vpRE3npf1yMU0Z1vR+HKrcHRf5Kd8PyU59QD6hcyMuAUS5aWFrcUoS6LgMTa
5SzHJKFEXRQh8BYQb3GeCAQVwId361U6/vLQi40N1+tjkxbDCm2ad/2PEfwU
V9wgqm7U6N/uFafv6DbSHBZFh8+De7UTxu8WCA6wV8pHMOe4jpjwR+nPWnhV
GHAXwFDyVijtcUvrIL0eVXDVFuKk6bZfr5Swd7zzmyrY5V1o/8u9tWpYaKW+
RMCAo5nRDM+fFLZw1JMa5Z0UvBHXlBEAnQNjagSDF2WO5nuvfmJkAef8lawT
BmkugcZKm3royA8T5g3eyvw3ZrIo8s7z3951QSbUvo7m84HHIBgEawPhg363
OhX6tc4+J/wOii/N+4I2aIXXqCGrn5DFIAmsnZQTmqX+49M8HgckdB0VBBhQ
vM6O1WkHMB8LQZVeQLqEzQk0zDU/cQM1WwksrDBF5tJrdhoHckcUO0FGcXhY
qjtFOge6zhEi2uwcCglgvmrMhl+r+5eBRAFJa08qpb5F2n6XqVcS4XTgqym0
S35p6R04yVzjdiRneF222b7dzLHWlVVsuGxkM4gRR45D2S/NWU+2s3kY5i0o
QBdC8PtaJ2FB38FEYBdM4WhNE5uPP8pLk5lWGRAXJU7yjv7+y5s1r4xSSs7l
4G/NASOK7Unik2QHFObgF4OT5fpg9BNtkiYtcrf0K7lSIlysnN/Z2YJ+UEE8
8we/NoGFj3PA4EOVQoXEB//smGwFwp8IZpn8E1BY1+uzz/42lXZb/n0oe35E
x8BZJaxqN0YakXtZIlb4Mn61gv0YZw3NN78DC1DsEx3zZFQAB6zQw0vBHNmY
7GH4KraFbTbvAwF6i2ASwTPexi4OAwwee5pcJ8EV2+nxfZ1EQwDiFBRoJwO8
YlgEOtH7ms0NZT6Ufr8ABDowcDKfohKcYADhsBFKwtqfjFY/wxPxXrJ1PmV9
SzBDol2T5sK+lFmWY2BldgrdbUjuypQ7PAtKOiLMN5K7uJlH88hqy3L8Q7Ex
kXZ1mqvraVcbRp1S0z5dvjGemHhktjjoo7hugN0wq9yW12BpH95X7ZOuOgyy
TfxYLCS680bUDELA17b/WCCqluaMF95j0Fdyj6vmaM7biTBo4nKbIWFFZozk
9zPEFKdUIYjLEYtEBA5BCSNOfApKGCMlv1gw90Cv+pWvhLep43I/JrLaT0CD
LLM+xo6Npoc/ObzTnd8rEVWX7n2YwtkIyL0/lwmjGrhpOsQhDh4Pwu44boL1
ZNKcwOFHw9itJfya9zwJ6aIwZHkHxXDEYusOQnJYLVzwryPZLsm66ir3eQLw
uESE9nYBl2FJHd1vh8Mm+iLJgvBYGt1auOnXpfCmr1tSkMK9MoB7St6wPE3/
nequS7xjolCEi9g2m64yYjQd/59X80wNIs8cxzjD9WP+xAOx0fkG1Kj9Owxv
6tD8SE471rbc1jxNwchN+QLlqjqwlI/j8hVV0nadAs9w1AMwj/OHbG5JdajX
H02ZhIxji2h+nEoF3fwU3ATlNtjL2WSERjnQNKz897I8abugaOm9eLzaCWhV
DAeCuP/vO2ewZi8hwzEik5SUThf3pu/AGyhPFBXVHqxm7fcjudajxTGVlMuy
vcIoON/mIbh9Dha4vmBmISv+3sU9rjoDwzWptO5c8jNvZgbqnq36yFOc151u
Y8LO92IvC/VQyAFD1MDEj2e1bddRsaMzVpywje7sLqrfxNt02UvW7fCwtnJA
xlpblT69KMNH+SJEzUjJpA3yacYQvEVBp1evzNecf2OkoA3X7BANn2+4/jOs
2otu4fdDmDX9kqRsv7K/h/v0E4n3vOMxrV6p5n8pwaYKqzyiKc9/hxEIXL3f
9uEDzYbSd4wxvGR8lJhkPy/lU1Q8b8qTHEm+gS1LRnrVlUFv18SSpKEv7RQN
8r6HT3PL/3XI+1dfe5/CUcFlF8lzjHpiIJ0E1XmS/hIiBD+vzAJQsHRLNJ8w
H62lJX5WDre/nivHRxlLxQCRDk+6d5LM5CneTbTVZVOz/k4B8xmT3WzOdQil
jkvvLb+oskCYXSNBjziHgxWuowZwJ8lhSu5O1cEJnQ6jDKWH/D/bOzk4W1ah
rFE28gwVsWuzjo/quY4CK6samEP2X01ity5rx3NigBH/eQ0Mc6ewqsby11QI
5ei8LSego/fanymlXuodbTuS0pfxG7SL4OZCQr0Rqb7sSIipmGNbP21Zabqn
SBBIfBQpXsUlhL67Ov72aWjxCk2+EtNv6RlgqpkTlM7W1g9EDEwPlRbQHX66
m3dJr3tKp3wa+f4XgytijsYfS5P4hA6Hw26VfcOqWOkYmvlIOSYzSdOaWnu3
LlfyZ3c2EPhdrbCsFNfRLzvuBW2J/Ze1kXiAO5waIMbZeT7dOM1KnTopIU4v
pM2Wm9FBaoVDkX1pnFiDQynUhVDM5veRAjyKdwtUKecnR5aYskMOrxtPeJJs
y0YpTboUAr5y3JBnFIiYqRMLR7p/9dZqDlyDnKmS/7qy+asBNpZ5fHnkhLfN
h+VgCTofNVT/0OiJe1dTkaZBnHn8o0AQLhKUKtS3kKpGp2PJUinm3rfNHpvz
eYoyBryFcnkYwjk9hBSJmCrTzMqkonsvuRcuD9vE9toXgS4rL5Njyl0oZ3jR
y3ANCpBzlEFRED7LjoFoqRKpNFzouuaK8L4bW8mnxv7UQZXnYe4+PQsMES7W
4T2DMW8EOm8Vw5q3zxxAE95oZFti0W0zCGdQhFMnvPPcFAL3jPaVsxmkfRRB
QmFknYbTHQfBPoh69Nx65Z2Lhq/Np8JkCDMHPK3clx53D2D1NfPeBshTaDi2
dR/yR1XLIoOZBA4d+qH+zB/VvkrCTUitbwFRNZ9wHv2qgRn1ZIELYFVI1JlD
WSsd9rQzJEFUSD3E91iMOgbKAORnRXfXSxV2ovw9YVGPLZ4Ls7jRFfRcZycR
UKNhBvO2yvunJVy3okNfoDvBKDrL0tD1LpP7M0HH0FxmPfzXrNNpktN8YpWf
Bi0gyJzu683Q9oWvKB8AuAPC8aoBESV2Qm+5PFTbURSPk2us40+mGbqq5rLr
SKE9+kBl0hvIeCMSSsNBUsje2LgubqizV6sfLFfF6XPs12mFoIBGo3tHDvS/
j96PuIQjH+KHenGzz/Z7FiCIpM4dNQRfYYaGzadDx3G+uQ5/ij0r/4U6A34x
R196SsuGBn0qx8PjsK67wP5OWYspWyh+EjWGWuq2c4Q1g6GgEpVyXJsLol40
dXxVR4UE4IA70rGXS2vTq5RIdfLmWdCpG5rSeP23qh9rf608aakb5vQodO8k
X5DYjHGNMWv/IElhYlhh5VbXNSMYCtf+0tacijdaB99YTBR2DTBzS1NTk+hY
1k75b/hf8+xT32UPXjSz1icFXaRQQg96pq4Jku7oc900rk0PurnkP/I0JyZO
xydX3DP6E8s+lYMGrMAszSPqjtmeUvfLm9AdOUDzim5jnIXpFu2HZjMeAFN+
7YhOHCqdhjo36c3wqRH+CzG9h8VOSGvS1JCTwR/2EPlCOfosT8QTe7MJ+E4M
nvYmfU6cdlO83y8orNCinwCCDOatIPvdgba/tl4OtLFE7f0awPhfAuhWunM4
/G7CTFrAQ9LdyYhhxbah2stBVDNwX2EtzFqWo8uv7K6CnnAmHfu5I/83uI9/
09bTD9nBniJCn9CPbZabX7GXhnhgAIDcdkAWUoxezg3PEMW65w6O0lGZDC29
+BXEWBVqVoYHwGhvhb0NXsYkaOMZGOgddE2HICT6XtcffMmfXgOhaLa6ZVf3
letVZJ6DmraU0xwLFFhqAJUzkC1MELkKqjMcIbVV1A9WnSZ9f1EVznWfY2V8
k+ZmzCAoEwNq0QEV/H+9BcKkYAcij5vZW1Nnrtv8WzH6NZTnjwWInE6Q4NKG
dbXwUbZW+cAN9M46z3ACSvg2fJT6DdPGUQqx8eEnlSNWlrZ4PoPjTVh25OGr
AuoBtS9KogEOLbVBxRS3Fd7nwdTXHuwXI6gPVeZVi6FTB4n3qgoMQyGevK8N
jzzaEAIN5P3BBJay0TO97FkpzQOGXLincbQa2mvRYfo/5NBdkgm1nX3r8Vji
esRBwn7wnx61tO5yZeBlsrvZ2Lc3mXZVjJMTVTVRZbnriLi0Bor6MwFHSoUa
npR2nopuVsAAnj1j28NH+m9qcJfGf5tLO2g0ikFIjdP1uXuHrq8HtOJ5kz/W
HutB67jOg85lxyF+uThoaLbCL4/quuWDYi/NUb+IdXJPdcGxrvaa5o+4x7Y4
ELJUUDH/NB39kJtlstW9JZc+CAE0qH1zhh0nKM8cU82tbCiR+/RJBdPuBTHz
8ypK7sPGHeWauHcL/Yp+p+RJDuPSLx2yGVDS1GhLYV9swgI65S8zi1ana7/9
bJEdaYZiw9v1DDxeVee5hxniqgdEO4klEpxfdSwN3oKRleuu1yWG6X2G1ZAC
jm4GtUCtaLil3/Z6SpcwVGNDNMiASAZpTmq+cAxjNx2V/FXDTmY5AY2kLgKI
Q7EV193QZy7wA4uDeer6ZWUmyHX641ho/dC8oweRld97qmcvgD5xnqDDBVih
L45Q6bpJXaXhHD+pmxv2CpDvXVD4NrAySrS7q/UYChDpLpEWcDFIuFh1uMFT
sgtTYg8JGmfueZFYFe9pYgi/nQ1/ISCi5Yj/htPAkxqyXMGqnCxSfzOl3JGW
jghNtTHXwemFWPhRvEL+7T2CBsDNPl89UN9EYtUDWUwBllJeaqBgziGAP0To
Ld3mTsjOMhZM8jsEPbYl+Hz3djwRB4O1iuBf0nqUkL2b8W1vnmS0cATgVR8F
fB1SeR9mabkBdmiIUNyef61N3psdhE0DToLQYtU1NxkyHVOlXh6H91ZyGq4J
iZVgYJiFYzw7VcnFMxLsDlbZpk88B7g1CyqiFTlLJrRfXl4NRnltRXc7s6ND
jMnP2fnoKU3+Poj7AqgxITVOtmA5ejCF111xyIUF+OagvkbbB+tKjjvwiuoO
CXfvi1XqoZbOErB1OYdD7E9IXAOl4OuPbSF4WflkRw4oTLNB5GkgpTY1POAq
uokpIP1YkSExS+6PalIckpn8mBG8Y0j6wCJOgl+fkxUus7pkLVePC9L5Qeiu
iwBWfA8AbkTgEsz2YgngNgTJuqzTtyoUZnDayEDGgQHuDh+oXz2IVvLgoGfQ
vVLaJi6evFKVOhrzkZyEvjZepzNmpnJOWHTmFwt0AHkTyp9iXdeuDPHqjq7B
4IyfkPBvlFkcI8Bnf0Yw5TunpmMN1c+dqWY+Is1uBynG24GiZV2ZlZxDWHpd
QwYmzYqK7lsfU0BZ3T/kZjBcnK8PgFKxwrbYkUHdmR+V/CRFOzyaaRv2ffmq
aRUvn9X3TaDT7HoOBhsALVqy9ZThYB5gPTejbP6z/HNQlK5jqIhoDV4JUe/z
zk4WaaemVcXpXlyL7tCn8cu2Ljl/w7qpbN7GyTT0NEgfLsP0ooDp7XGmZAND
YxpfyWN4FRNXsk7Tev2QJB4VJd/Sz3Mg3y0N/ylO5JDbPcOQ8fwYiz3lfgEZ
8IuaObIBse78kOpfKJJx/e+cBeFru7VBdjEgfPwlBTFZNbj1KmFeFDnW9Dbs
eWw1x8BwFSIxtZyCmZLTuVMmR+sh+mMW/0Zcw0lzoX/WKnuszJx2AQkYukop
D44rAtHmiRpKds2Az0NIdn93O+MtWhuaqA3BYWdGPdLYSey7gpyhIxCUUF2G
528wqhHS07TTLkJGSetXwenl5Pwd+0anTHHDE4vKA2sSjvEaqg9/0xHjyI8g
x/9ozAK+T1q2buOPON7aYI12+7h5SpWQDGnGi01lYhCfPYyVIuykw0qhs+1I
RbbvCzUt6KYqBNnyLxM0gXJ/OHFsr/VjGPXelY8oOXH39yiboKuPxGsXgu7r
Czih8Addwcbhv+gfCeZgPC8DZIlCJxW5blao2tpdx4zST52aJB/Rp7bbj4AT
VVe7dAPYBqKOyhzxC6TKWz4moShXnZYXYBuNkzY/WM1EH4iJ1+u9/SLVZWi/
g6Qi2SkiUPh1sfKt9VDSIjZjVyzG1TesbfpTpfdUfIyLGj/SVHOCYmSq6nZf
J9QmIhQ4xDXVcwF42UmDNJKh2JgEm87e4aEEVEmMcyvHGgi8JbYhrE6oBmfk
L6aiAC+YqX8qDPfUUNJnXgMZR2KhqzaONQedgm9hj6tjnqJFApVTBywMfquD
c9+un0wlrpedPDsRi8kYM+8DKLlc2SPTFBE2msZ0ZGj6lkoKz4P/7fr37seu
DaH3RnPee4PyYLFsqqSuhaynoZZx7SwFzDwEaAqfSwBrH82qVSFNT6xvC9wi
FJ9LMYIMsL9q+tx0MP5fzVLNv7eww3i8rOAlNt6IoN5arZydFrxo0b4nt1L5
msiw+HP1zGGKWXMUJ46ecDhCfW8PqFEGShnN0zhVVU/NXjoDB7kJ1WnPSZE9
Dh8jUBCwQQSqanHYOh+A02XgQIuREGadj9bMs1P/qOgYkmLT5ou6eEpRV8Vd
5gRv3MB+hYrFpjHhk1Y3a3hmfJXrKJWXyQg+nt0eA6O+zaV1p2IJXcUuTGEh
vcYYA414d3n4GTDEG00PpfXWWTMYZepSHa01Ws2LS7VS/weqc6DkeWoYbvhl
Y/uZlm29syQzU2bdlcZp6mlEZaKpDrBkjWCVE8RGLKo558+Mau5IwJtSL5fd
K0fJGik1f4Yhq+cbePZGMeHmpc7pu8Rqa3PMl94hiKBNf8Iwl/DPN53KKynw
W1DDlPoW9nwDKnactBGMX3aJAIX9Omdw0nsrx0UlG74mj5sEHzEeaZvjf43+
vwaUVwZ4g6x5mdM/MeB/p68LggB/6eyaOoyOI0CWJSTIErT23CnJqUTSmcjs
PZad6hCxf++dOEA+MqMnxk9usn2VqXGzSAwK+fmhQ+Kzr9lkRjfwRMw5B+Lc
MgeK+0a+CSqPM0BkDzuGr/aHysqvXHkyOKuAjEZ+P5mOjMMf//AOCWB2PS7S
e2gxtq2JS/oSg/b1mAvPvFGIv+0Ib2Gd2aXdcp53v27yFJp3JTWCPnZIRJ+e
lJMtMknH26OIiBWI5dn7CULF20XDGpTeKmnLaoNecKv4L4zhrjGi4NaaLYPY
AKyKZ5++ed5heYu6gCb/gKQ8/scGO7ywVDpI3FOKrr7OvWKxchGPZxyQz6/A
ITNg+hWWvonkooiNtauRmHfcTynegs67WqdL4NSExYtqlxwhQ3zJA+dsyXj3
hmr9TW8IB3oY6aVCrFwZQUpi91cVFvu71zA5IRX0W78mwxDmVMHC1Nk71xQb
NLdfkb/EQ/RdOXsuewSfiaHWu5eZAUzEsVDOv7fl4ICAMK2AueQgQan5ea+V
N+9df8BviomuPoZ2zKXGzcnXkG/SsEfkHQYp63Tn7blu73S1VekTzwt6F0Wm
RolXMd/IgigiiO+s2k0LZC+CrCtQGtygTe/DF/JuyZ3BydeRLdOJ0dpH8fE6
Zy1RdeCCjK78G/5y3zC/9wVdykFDbroXL/4a496SEFkMBN3HZAfoIOYMDBxD
/QVvugdGmPLghh7Y7VK4qfjtUSJOkN9j6m/u6ofaieeaiqyOqf3ccyfpP0Xs
AbOZVC5kr8cVK3BJf0ML5Eau/dieO8IEUZR8T2zFe6midkYeF7VcBCtJb6rK
7pGXa0FzDKSFZRIhOt4cYkr0UiaTa1eFLyfNYRxH6aF5TaaeuHwwkiGXoITh
EkAWjSaDds4P/IMupOmKu+r8SNX+sxRetGV5W3fZDQ0Mb99MgqElSs1VcCOk
/WIs4aZZS81jsL0xMvCaEYGvRrwadBRe1H3lrAstE/+dIW7O4k0YwHP1S/sY
QpiGqYEPgBQfYu7HDHFya9NAC6qZWo4mKI2da/ky11xu6KNwkNAHFPh194DV
lPBrk+7PX6Spb1qAinQdvueC7snv4hGKUuvlMuFVzFE4QaNX4MUaCC8YL+wu
oxbz/+SoTrIxwmeXpcOL1YnxPnaNwCLvo5XQzrMk+HWu/RhZgELo9YpAKGlm
QADZMYq9GgZdC9HiJwamFXsg6wzlqlZMPNesilFHGSL7qW1IkXSVag0x3+wR
bjsQj9e7ozCW6WQRGzlIDX29jgolnpJPkgo6t/mYCDgEwdnd3aA7MkAhRrrW
iweB8Scitv2GWFjWN2tZYfR2t7gtmrla9o6myZqXHNMkICeqPWglW9DwKgK5
LiZLlJbnPOC0tg1Mj2SCOK8SKO1z2GviWjqNHJ3HB4KEXxzxYo5Y2z8DtRLw
kO6qiarPfdpMWGjlcRXfpV9djoCvBL0xFq7q0Hd0QnOmscbTlH07YygrjlPx
J+uUdTPCq1OoOdq8Ker6H0DbNvPA1d+ZqtUHj6+HDwrjhVbO9QL/Njle06C+
a9g4AfLTDtV3HYaxUX8rch6hPrwNcGzL/AJo5dHWtIcB3w3i2tCXokp8lOgd
aWEH/fFecKvxmubRDzYfzPPc2SoCkq1g6W3lLcnDWHeXMAYkOJxdpv24BkOA
+zOB+gzl9aa7XF3P8rK9IWvFKDMQKf/vvaG2WRD++D5J5ogj3mh9C9E6yWvM
TMCFt7h9J/FUnEBphsDNg5DMkrUfDdrVFCqi4EoJRpTuy9nTSUwBM1XujLKk
q/uI4y/cfQ4llqfOuwMPFC67p1TS7wXIcCf5RRPSoAMiAmMmP0n+2oD0ag4C
9BXCTA7q+udpRZ8va2hllqLhF6FZOo+GpX3Q17gGEdCmyxwB8sKputnq+PRe
uoIOxBYrT2vZ53nvaLFecCrgFuLcp/GooJ3BeddjPf3/gTYtwv+zBUd9NCl8
4IadNMEv08IIvRZ+0KPK0kO5eTemJTw9Aka0ROUutJTplQgQbRh3BeGZUsGb
4QvL5gxCQOAkY6vv+gop3y6ceDaSC20sAxn48T1v6EI2hT0IxQOPF/GTlidj
TqeJzdBFOhm0mDo/Q3n01VcVWtehbA875lIuSt+qA/5HAFwUJWodm7dcyQ2C
jcot8x7sz4vd2pbu5fhvbng5u2GYjjvThmYXbhShdsEILwQo7tJrKtyH1dGo
SFgnIPZChFTgHepeirRaHsxF5bAraVy4QoAOk1BrorM76W/S26xcuUGNg65p
mxoNFX3aGaaaeA4viG6LFsVT2le4mnlAxQ2nLBG/3N7ompxPJfd2zq8u2CV0
TjxcQKY8QMD+8lujhsFLBsPK9nt5ba22iEeiSxYN8k+Fc8YbHwFZy3YceN3S
OvmsWg4b9jvJ7vmlf2r0D3F04Pu5egEQXR7IoMqHgEBQcYAL3HmFCaOxEIuc
enmt4NBJXgNC9qACkFMVkhGkoU8QIoXA9m3a3bQYS9XUB5XFtXCuitFpJ2n1
WTYQ35JefE7L/ImBuorfi3idgLhGDcTyK0WKD1xO5Qht01wdhXXMLhulq6pt
Z/ryAhYUbjYcyvXfhkL2nOH4W6i8IjUTRXjjJxIOzAV1KtIhwH36gAoIT+ox
aFNcCeLOnGvIIZgS6CvCilA4z0wtyjf30cfC+dq6TYkk0XrPdhw1KE9yCs2H
6/7ZK9or2fvt+ctxVxmbFRAjXnyXx25kyo/0Zg0lpGWyaTA4sSpcExSNIAoX
25xehWAC/UqixnwlkzWJ62svgMtGDY9W3jDFHzRsW7iLzg4OOG+R29hy50D1
/v8LHtjv3x/p4L8uMvS/jphedZVuYCXzlHUJ4CssZdXuVOqqtdaqvQ4f09Sx
5pwo1sdDVjXi4h3ocrTACENVV6r0uNQRk129Ed+Q3TYwavmPqfrzR1zJu16E
sUZZKzqKN8qgIc7/o0b4OVw2WCbpjS7ToRWDdNSEH31QtCUaOw8uWCfOlF/W
gjCUkPKIIx8RkrrmS5jE4NxA/3yYg2fZTgTKUIc8bVwpqC3Nc6aEv6OMXRic
xpjTafwHS/5QbaXM5BHwHFTwtH0PrcAJGIIMGmRFApjrONmvcO4gWzaIRY1+
iFIRkYenJcS3dxgXYt3UPV9OO1KGc4xLgDDsNZ/udXlDp9AJa6tja5plvMoO
vXRD/Rd9z+jRudsfGwkvOcfcGnpqGN9J9YK4ihVq+wdJZK4RgcBEmis+Eifz
vHgwX6gbTafiB/sAGx87yhRSIwy3LXbQeHCts09eXtqvQwSBcbCooGiYNNiO
yC6SKcv+UqYKzm/qv9vhrev6dAw/Hv3N+8m3VdSeISJmZ4bsAro3KxPwOHmE
VZVOuK/qchDAwuv6KO9WQW6VXc8DDPpHp1HcAaJXHM7NHmhIGmOobJA3EWLQ
2Hv8gmKeW4skvdfc2vWchbolJObgqcocR+1Vb+60w7h+iqrv3yLcCe1/vJHU
AyY3bEJIQxcYwKWMPy0kEh8N6fBZSd1Y7NvrkAMF7CjA4GhE/FDNuV0ergMZ
JxEWQjwoYcoGOd0pAnB6zJCYqm8kSswtNBFAte9+mVUMSKIwoG3CQe3nA4qg
+gnLREoP3xiZryJr7eWUGETCpUy9Cfyo+HpOsjtglqR9BP+lBuJYL6h3Vks6
i9Do0hjoeiYA45egsEUwvfUCq4nlBdfvMSInG4v4ubf/atgkYGx78Y2t7oYR
LdwqrXoJvT7UvFtH6wBgOqNQMlLU5Li5AyP0pUFdpmTRIxDMQ6E/m/uKf907
bsrRX39/O8v1riKSEvZZtI9xdw3XsryVI5D1AdcW7y96JhFapjAkchn+7QFM
4Rz5xS49atANaD3ai7BokcEoeeflwgseZsyyJdRfEBvlLlhZSCjcCP5O21E7
S1oVWJu3AMVpd8V+/N8eFIt9dR3v7QtyPU+MD9UbA9XKfClMIeam7B6pvlXR
Q44eDJaJgSRM1jZ6Y+A3lFYAykTBPzKycM0ZZGwv7WMAhlwNyqjSh9gc29S6
U8BdKiFudstGuzeQq0ETZpUIIN5uIBWWRbjD4SG1eRVmzT2v/DGtxM3C/3EU
qWYTm5zdQAUtxv5G79DrcKj7ikoUzG7beCW0bDvlel+GAkOVKiTggCyUtWj1
+ybaipVt6mOYSutIHrmsoF6v3P6MaUBVHgsJzNNKHBmJ1ldbC0sPkzw6VvSx
1nN8ITgNQn3sUSpMtBF5lEQ+/SPFgghF3AD/FBIY7KYaPdzSGZbpNh+DM19y
OvAK3ljXJPgu9QbtXxWiHJ9gxM2O6T2eCNMTlekBWiYZsKYPR1ihF8aORgKe
bX8Rl+M/7QE85XQFggSXmTNjdWdmG7BJlVmwoPZ5jxW89QSzGWSj3IVNjth5
oPZxwyD0axBRtfyKjd4M37MKQIBaUN9EfoMzCMwKaUFsHdE3JTNmucN7eItC
k2AbCg9YcJVsoLE5Vcz6Ba42RCFbDOMQBp+aqVSTudXx6CjtGKaLbJjR7iq0
1ynO/+bNTq5J+rP4axHL4+8MCF22djYUCJ3Mt7LyRW6YZUb+r43jTtX7avLe
7AaTePwNHNQGO05nGNMDRFJKlroyB3nnjwMau0m0dGOh3/sdWYOZBZqtjZ01
j+x9wQn8WR9/FXDEOqqi/AoXEiU6BUfnZrSG3KD3zTOU/klNnF7SvpMloU9b
CYgfZLKhjzAC7Jyv//sAkqa+Mu8F82ted8sSvY8R+HjubZMBRJOefv5CcCXW
s0GUeZL47WKMTmdoB/IvkTBu64af2ZVUwsSRLziMhSFvJziyGbxcN7PKdd0d
oZBpzzapqthbdw8WsRq3mR5kv+YUHDkcg8Z91n8NESNTJgNAbehjStieVCMZ
OvnH8ljQgTuWrD8iJqAD5YeEF+lznsa5rla9r8CjZRTlu8Rq8qd6eL8lBSiW
rUxks1GzAAR4h0hKjKpO+iTBfkBx4diW/NkSpOs5bTkJM6SYDvBOhOR3JQLh
nkaIbEgGKP4nQS1nQY+VlYIlbUpM0ntGPJYJIQ2ylQRlfOdTuHiYbvjSMaLP
TcY37tmQeANXUMispffaKcahJCl+pIbt8sbGHa8jjtN67Rcq+1oredq0hY4s
EezEV/rbZl7yaVcwiZggYk8w05dLAqSJprcxRxBZWAvx9CV4qzsXC8io4Mtd
NelbVWj0tGt9tHPxt8VChVPBKRK8XbRJ5D+9dN6TwcXJnLQ7GCYl5+A4DZA6
8tpGIFBCM9CHuyOZsrT3Fr0gkvEkV3KlLRTlBJwyTlB58Uns2BPvU1UOFQcG
Uddls5HwmMQ/h/hYZTrRR5DlLxiEQRs5MsH/pXbZ/QjzLTmsWU6M2pFIXOs3
26sw3CuLBtdaM0LHtJqWhpnys7YxIY6qhnfkYoy8fJz/dW6nQ22a26ROeSrQ
OckqFVdQ2mvcRehNIDszHdVKxN3uwcEdrSQeZH6y7xWPCsJq2K+aV2JE/Gzp
SgrDfoiHI3BudHsN8r3ePC0L8uwBDEVS7svKzin1l8dyO07Ysb/ox0W27ABF
OS9+F2R9NF1cCNyjHM4f5R+W0Q/AeRlCf4FO9b1qUGRoRm4uq6qHKLKBlzXb
uMBYCU73XDtEgxDHliHa2jdgypkw3Cfh69ytHgoIiKj70OG/u+bngcOoQfE1
1Na+/Hfwy+mB4qC5NazLJ6NrpdZNo+LBkU/eIfK5sOB4EM+ptMxXk47fUEeP
Hg7xKc1saOm7xaxNqO/oE6ATnlROPt81nOYi1N58VKZNZbNSE837Z7bZayZP
BZSgXB1NlBCAkMOr/CwVBQT+SVgCCFWsnCtxacg9W3x0KifPCCapmIIqfTDd
82jEeH6pmWnj7Lp9/pkASK84MNt1TEl/ZMuO3+yKyMnkRHzPBs9JrerakEl/
6+ntb0ZtXZeX4L0oUTNyUTAtHNyYJwuD5sk3w9mg9aQLWU8/OKrUQL+C940d
HJ+XTdVq41c6EP+KDJ4iG1bejI/p4YdpsfnRI+hlS089jw/wWhq6aLstz33z
VNElEyWzpQHSq0qh6jx1b9mjS4iEvDCjD0vDYDa1nr1XLOBqIqRp1tFQ1oCw
rSFzBYgZbMzBd8aA9vplZ7JVASiulxX9W+tDLvoDqCB4CrWIT9Hat9emzI6e
3Gns532k+vcFPSevlE1cQihBcL2ZPlQXxjV9Q/hKWyMw6v7OPgfv+G0s7oTw
WQAq1YGntd2QempHHEfK59qHCndPg0ZkrgkIKtnBa1EIjrIT6hVrI2mwcpvc
ahJ161A9WObwW5EpO7BYVyMOwx+1mJxgk16ExjEBmmugAxe1RHg1l+cQPCdO
bA9ds8heYsrmiNcuTBzHbpFZttrYaJBHWrbPNF1pvK9xOge3ucghUlWC0MtD
UgEOV5sJ78PXbpx7Hprh5HpxytSEAx/zoOyzVnXwbtP7W06bpgzSkfHe8sDH
WLDujf405LNXZUQbIcqvPxkX8FBPSohPxxVusWgdzdQUXkAWzOABWDsi2efH
fmxIKbbGE09cwWNEkquqArgjdz/rBQpsWOgvGqyIIdzwcC6LDIwZrnZS4X10
eNZfX0blDagQN46AHgZGBe3RkBjxncrIubID07k+N+x39GNMmfkdwr7eJ7u/
vj76k7y/egpkZ54Uk1Ex2jrcdVCGY3RWAL26j56SGKwc8olnZF4HqNKjNZ6Z
J9AMeItBIhYS+OaO9TFAqiGEkUsJte6ByEh46WuO/Jex9k+lynJGFjaQ32QV
LLLIvxv6HfuUbTp2ZgEUDPBYcKKY8elexm3f0vyBemDA/9vX0I+vyI6vehzL
PbDSs6CVDMYpbJTson64JD8TkXoOkAP0+5enwIFmbkNgar0iUdsWSKzGwYJC
20/IH5LQnvDkSiDqkk3EQdiOuRcpxvlQutNwWfA+Ho+6fo2fy90aXolG8BeR
Y17tvjUM1FOBH9xnzmlpsvWikW+AdIoTA4XEdsodemoVYHLmLKlc6JgpW1Xa
tKT8q/fMht5tTGVT5UAtSRRLgOf/nYzfsFa0sZeUYWGoFNPkFffR1rt7UPDF
Yf1jMRd+wiTzyQCGKsSOQ4lfAlwxzXc1jCNSjWCoQK2yC0739wdhpVGh3ELS
Xj82iEEtoVDIuDZBeHoycsFL3jJkEKo/kJ2JxiLx8PK6EbipHwbL7+KRst70
tPJIUfXCyl3gkKhTSD28L4LLgm0+BT+COfg3gsJlj4hz1ptdyh/1nzNJ/W0r
bJKcj76t1WotnZDW9wgc3LHRCwDIrieGWPQ49aC+IZq2jkK0a6x2Yo+hcNMn
9rOvQnn64ff8jKNXPMuiVIBUqfmKSArRh9VE5aqGedBeJzX4LWZFdPQIQopQ
oXmFqzkf1oWPeE3GaszL5dX6uW3lsRBegC/p3XV9MrkruFRU5yXqTxZkOGab
kbPaD3y3Gylk1rWoFxVJtOepd0GXLoYhLPQeTFmhpOMCMZkJ5VwQOhV419n3
OiHrJz9HekRmjA1joxWMYeB/TWhyfuZU6f7BzHv1W9BcQYR42RDKoqAjySBi
q8ZTjUomsvfD/PsxDnDNu/hJcUV3wT3uq83rPGYPdjhbFNUe9V8iptejrX82
BOnaxrRXo8P/pSX4ggtM+3iypH7E0+M35ymyE2QBdxtSrIfTr+o/vQni4KQw
Cya8e08q+3FAiVkLQNM1EV+zTeHp3cIoo110lvRmTpepd3MXUeTUtxXKm22r
dCddEwPDUqn75DUgX5PkL28wj6aCfu9nSN/yfm+7ycn0GMmFtGGW2Jke0KGY
bI/laqPTbxXfRmHH4WrenBcKchFbOxXiuM4G0xZCe7K/FwO14z6pjMvsixN3
JtuImG3ijYUAmlpJJ59zpTUSTSELpc7eo1YAcLALSNDyP2Ic6TC8ReJ2owTW
/VLe5Gg+hI4Z4KRl3CHAr8fuNQXWhqJM8fTvNnfCuDiXI0RgeP5VieH7GXIV
9LbPrleJxj17VXT//LlLxiiozmskd7q550BDsmOOiOiZUVieAwhIYPBp6ui1
Mgn+hNP94WboGQKdwpgd5ZkLU/xCJld7sGNWT9dVCbSjoYe+lSGPdrIsCV7C
VdTDCccby1nDQxI++//ImXYcG7A3MgLcUYzMo00/+pVJRj4n5E2bIZwWWyv5
A8LFbd6y9Bc15d0m6A87km9qBHUXGfBUaJyTThs6GdhUISn1CKh48NlQX6Lv
/3p6HLEYbcnSgf79RCe7divluJaC2HVcIJO+R5mO9MCc2xuWXSRCDqr0PyYi
1lqe6Po8epwn7gWLLckLUtELj0Y9O18dShyQD8grwhs9tX06d9JaZo18dWpN
J5uR+XrSfMBTO2lKIb/88xTLyrgkDzMAXp045kIFoeoGMDSEAAQerCoAnTpd
FBvqLW9BXSCXdDeuS5dJ6INeJg26PwTc1WO2XIQpS0gtoB+wRh/0AG0PV3Hl
WgrU4IP+C4K4xPsxpUkYN81nK1X0MAn8Wkv7c7J0hzE2181xs8HZedIqlc3U
GE+jb664I5MgKXfGMB6TzxfGakBkPh8XwyL6YjcijF0kqfZdcw8YZAxCNWjx
EQLyw3Hi6sE+ZI6wOHg/I8Ko84ZfGIt0yJdYRdBJU/zRuLvg58UbZPQDObu4
R/xmuDBaJK1tZb1FsD9yMQeBvimP/+BFbsR22ZmxHgomEOyQPJn2Uspbs6q1
U6UCZCz4yFL2hOCBe11de1GXSf05DqPFiNQEz2ICwiTR/IvNSpd1zxTtxfde
iToyftHN7gjNW3t9XPNhvLcNq7bUB06FH2kIMlFyrb+Ygo2vmDcyhFJPGakK
U5T1pvBynQg4lSt3ECKu+h+H9RIOK9OClLrZJLnd5jkHaK0MjnSCg76athzi
MQYY+O9qUk8CqFzz2Y1Vil9ZCjxUox73zDMogjLLScBIBtwOXJfV0bbb8Z7R
LXnm00miMhO0nbChUz7+z69KDK5toYZQORBuigdLo2zpwIYnPF6hz1DYCXTh
RH7CKfFQPK25qnaRkYIyGSHWYGW0P3bM+pYw2llggDG4DxowqIRGJnmZR7D+
d3FzK1t/OnQ5INeqRFMzfeU8+5f7Ji2zVan7wdCyJ2DXbEv5s8wN+j3Ok08c
Cxn/iHHbcxDhJ+ZZEl69c5nRw4mbHwJQUE8mT1kmMvSiQB+9UV+yv4b6jGyJ
7rOJGvdPlyDx2LPK2ioe6lJpwPAfqyhPtdjwlb1iv2sUZyNbY7pqX+NWmvnc
0+RVQXCzzjGpJIPgcYIgzkyNQ2cEerii9g7mpRLmvIFRPLzjbuxZJOJpbzHP
DcitqW1cQRuge872wzMVeY58rnIb89f3Vxl/+xmjv7hyJWiQumis7zHsjk+c
QBD5dpiXDir41MMPq75Y+x9EiPWz8Gqp3IA72du4v0yzOdmAcVuohCi0loAt
uaxgGCsO+aPRsYZZLrtta3jMFpeiYQGL6pUz3OAaqqWt318iaD4TJrm1iCuK
JoOmP1FVm/go64qlt3VbFRQgZYDeggQWHgg3C+MpxTk7wkxnTCNFHIkcmecz
T243SLc2lbJJTjXlFgzrvmq2Ng+8V8gQmOQ7dybdLP6D/pjB40j19MM5h4Ah
/onogiz+6s+XM4Ru0lCyUYBMpJYj3gLVYbkHWQmpBo0mlNt+GSPgC7KyKfx0
ZSlTCJLghZbJUKGrZnxsOa8kLqIN5axf2QbRGbBy8sZvWXlR4xSKXCaqFOFq
sQBhuiypa5IoY7sH/srTfQgIjTTqwLetmBEWxGeQJOmnKWf6qx8HAnEcT36e
bcWAu27itDBnKYZk8MnhZMbjzUK7Vq305CL9FRthdJqECt3UiDVQqHBpumxY
M+4IONeto+4fPeESs+tX1U2e6DmvjpEc1+H+u7xU4UuHDkyJAh6O/Gw4APWZ
YO+6ZDSfaHE5rMm1yKOrZSvPm+vNmDYZgII2cjt6yw62nRQt2yfA/Hz9f2yE
g5kmLOuWvSc0wCJAP6p5DyjChtB5mrTRFsLTjW3oR4BH9WjhRtJ1Yux+YeHj
tj3ulkCDjBrCQbNgCpBmCCl5ANIDFVeyOiTyD7Blto5arNMp0/OBICSjnPeG
0WfUbJ6avWx720wt1Ohcj0ZnDGMI0AkGC/u1sZ8h3Bu3+YqgMf1PBPVQtvs6
1h3kWh11Lg9tVKVoq8FaPrQ2dyVC4QJGOHlsznwekVccEwjEwxrrbdj+fktX
kwQK2kxNexPurwqq11aD4+kZkwFAkT+7ZeaBUVGd6njNDISb0bb0bEGXfi+l
xp37ypfTS4t40wC2a805qaCqx2kMGkeuFztTNa1yguBastq14rc4txmWdWTL
kT8Ko3u5s9w7U6TArtzSjg+Cp0WzR2r+sTTlX2ybFsb46uXKNr9SV6VRUhcU
yh7Xo5u7xbx1BMm3dwhqn+o1kBMoN82FrBUjNbREd42u0F3mB+b2xLZkNtn6
+87bbw5jwihuxwc3+D9SsUX9qWVePvFGQ+1SL7XAZTnA/Rm7jd506Xw3tO41
cJYKrES1PRJ8K91LklvzA4mo9HRqLm+7zqITI9xjbp78ucItAqapUgeYgWSa
N6pTe3VpaQr2WhSMSsiJhXzISEs90msGjz7wW5ahjYx8mnOZmbchRgRv6AVT
Ix04JG3PihG9HYFRrYjNoQAw1VQ58fzp/77Q/49q5GOp5ud893iI0f6wcVDN
y5WoElqeC7gx8cYvw/ldCTyKzFuSmWcwQ38bKOMY5JEX8Z/io8QS8d7MDwGN
QWkm1IEw33kkLbZHs6yQWWitlN+EzL5rxjiG1vPsyzShmRx51+1DL5zXWyJK
LAGiR9UB73vC0wNUse/Y2O77q08h9InKw40hqCe1iX78ujStHEQbtPIg5H2n
vCuhyd+fCf4pC7quMH6Bnt5AbCJ/5sVIMdV1vnga4ILGrCsdI0/gmwSM6FeN
oZvnrABIj/jtmBuF3nKK9Ck5IobRuqJqrvPWN2/dbo6V9qb77vzKLqOYDl8S
YVdo0EXK/9Xqz6FugBPgDMVAv/UgtqHq522LcU9CEgaMGHDhwmGFjNbi7cK4
6sooumr409ojhdKUO1S2FGyrQ5zL7Lu5ZUD80VBOPCvWinWQc0eG4MdjQcgl
wzKEijw4hVjtCK9tfnnEvcDiAmGndpfjWXoYVYfyKe/dczRgN1CJQTL9GbtL
h2QPpz5DKMn1PEXz6G1hvNmw5Az18OZ6D+ID6G0a7Vx3asDMlaWWCp6A0KFB
g46LcEGhsirGOmGulZ6r1p21I6ieEbwdICe2tH170bp6mBiuXuizSrbB++0H
6g+hXYOAoRqMpPMo684U2gdvlr/dXyxNJON0XMCkb8adusPj8DjbrpjyhDsJ
zFwf+KPj+o7dLucWHvMV+5nELwcWEKvwWkdiRnHzyhiLW+202aXlJe/znwgD
CpqoB9NQhlkdwKCVfVGXeq3oaZzOlLXbsy10EoH6NgnvOa0tV5gOX2DTW3PS
ghEFsWux4SDqQ7AOBcvm1X7Q+IPfnCTqx69eM2pQd2RgxN73H8F0PRaVToP0
UJL3vrdqqj3qrdiu0NkUfIso+JM3rVkAD3nCzGCHvDjpmJcbJegSjwjfKjZy
10gKi4VaGovsMeguiNDm5TCeg6l8ebFnNCpbXTiDW5d3AoF0pIx4Y+W6yABd
bAB7MFe4XUmQjdKyMkLd+3/EZhPf+wtABnHfrjzyHFGTjeyn4IVTTspKaNoV
HylQlmHXxlZBpVKTwGx00PVzJITa+i0LEqp+ffuu41gVvg4pISJiC691JoZX
1R5lHbCR5jhrFw8nuG19SXfH/wGAp8hn3CbncyTfuxemfibQ/9gblCzWKjWV
0bQljbQ/sSySb4FTgpnt+HyFg/tD/nj8MfvwQCgNWdcM7xmfc3l6QKfbNyTO
uHoZ1jtmoRKsNmVDtFHhRS0wIyFO9CwHgQMjO95z3eSfASZRpPMqcLg9QkUf
Wk0qUbT4t9iSsUSrQpuPzJWj8opjvq21vjXSszEBEPODoeq4bmkCisfqKcwF
ipmVgKVH8vPxPG905UysOFxQlt8PPLz7fikaNKXT1pyIFOlbm40zIk7UXKL6
1T9olkV6km6YOleQmtB9RH32euwXcA7wYqgljboNGraLYM1eX/ji4Gh3UGs3
XDdR704YSbhQ8fJ6ZVWpPntdzdik5Wy7g/6CEopJntR+QZvDPZrU3f09PMxQ
gNi75GTuQAQlKsTrkk0pSSDeZiuj3HQErZPvkY/pr62Qy7TGheiIJmhjSXbJ
YEhlPvAvs6Qc7MWChzmkkOSvrk3mZ0UFHS1Vj/r/K9os2Zg9oivSWgekJ7x8
ybrCbCJFWEiIaQ3I77amo4q/NSbhLSPuvLKF67IDzrfQfp21ng+3hcm/KlXT
Wwid12NTe5bW2rjAYCXT3rmdeNOs8h50eJ7cGkMyPL5ZQkJ3zHN1FEYHpBJc
/jxDsx+ggYOoEKtYMa3BK6GOMBvu5Ojru+wsHd0TBjZ7c9IMdlVFXfwKCP33
PV3SX7vUjH0LVmJf06xcBl9wqrlqOvCbCZKGyXGVN7MEL9mSoRgeTl2XpD8j
9U0+LmeEs8ssTd+BV+SLRZf2jbHZm1gjnbmLuOoO3O+Sv80qrawZp1c04gs4
SChi7w+gCbGBog14bHNJ/W6TrDpo0Mm0uVnomHeqQEqTn0DrNQXGiOpAws3U
T6NGLPf3XpHfyrL6UTpBuj6nk4hB1MnFYi+e4SGmeeTdYzdP5jkQRrQbBbNw
HR9E5bJTJrwdWQNuqa3nRyKtu87EJQYAi8uEqsf6Gj3HmiqVbO7YuJvAnOQI
3k511fDok6BWt4gTcLBD36AVthwxGtj+jUMyU8c09O+1u8cEbkb36Z6GzOyi
usYzT4USYOlZxT1QbK+BBZA/m1anFd3SR4nImRGBu6uHkB0vYsrqxLKj/bKb
ls7psmq5yfXmkGcOCvc84/4zzSt5eQjDUmMdbGJcyHmp9hzec8uvw6HhinTX
bqTKIwIXG6Z7m73luf9jmf0sdX1fVHQFHmCHTkAlvgT3XMBiTIMELvqpjUgw
kMEjHvWDV7TBbVh7EpB/qQgYtNzMLnU3irkvwBDjFqkv1OXt6Tq7QuSoz4Zq
0qQma5x/DWIZnWJvuzgG4OPJRgpWggFLNYLYJPlBqpgchjRMHTikB7T6g36p
j2nFGRZ+lN3yhOWdxk8SXVjVF0is5fpDLDRp6cSpxAYNmRSlWjF59a6DgsTv
PRVkFRkkbapAWt1dmtT/QvsaZ1VCoSgFaAPosSJpmhlWVZamOWqUEr38AeCA
uA2tuAkGHUTovyXlfXg4Hnq4kQEwLtI+qtA7YH0UJmoK/xY938GsObhUqcSE
bnx19noJaOzYqbArLzGKztP0hzHUxyb6BdDbNRP9ErXI7b3GSzvsuvMiApa5
O1ACvWPuEW9LQfjYDhwA6dLAaBGB7v4X1ZISojgbo2vnaUQ4NXNpGvkcvoaY
53WzZ2HuUYmveS9NjsbWInyPj9LAwYLmwu1jQ6Bow+HGZ2talpDE6aSRW9y9
yvlATUhhu9s6BUwhYS3ZQ8ynk6034zTEet/rQNMt/RO3Fq1xPwXOMr8tudC+
Gp3ZddC5mKzWlyMiEJsaNlxAX4CtY+OSRuWAZEqrjwfxBGxHvYFXKRSTZSUd
ONyTioN1Lr9wPVNWqKtBGS719Srksd9nrNxgrmEnm1jmmsZoCQX6/6C2vzlX
BODeiDjIR+4L0Es9bv3se8BTNQ8dg158d8ZAxoWAJlAzBkfXZtIHUW/6r9BR
spRq0phMoUIXuneeQ341iUN5/Eg0bcf2l23zna2nsj4ESf0qjh/H4rEwSTqY
c9sSrqh0F10U5TB7+pMtytwUpEsGstRw58JzcByI0Ea4+8XK0m1GciYjqVI8
9UUjK0JcCiSHOLfmuWNvGWe+WEsQFnDsBsCYBlBvJ9QZdgajH96A9XdOIcFV
Hf12Tcx1grIwaj9qmPQ1CDcWu51p8SLJCj2SsQe+XGH7+m1OqVKH9XDGVbOV
Mzk3nKdUQPJxosk8tSlZy/4fQ4TOMPu1+ohwlVlR/JQX9YM4fFdFRMXP8FDC
4J3UghrAboVuBxmJda4+fvZUOEmKIEsG/QHK/09whKAGKzdshy+GGNAtKXHK
5/fdHRfiVNuqE8hWVfQdlm9f3qBl04xrE+ruYOzglO7zgx4QSnjN7AsQmoQO
dnEqtGjPDztybXZSHaYhilXFKqAStXAVliMV5p9fMcSMGVgkyzIoGfHpFUut
oHvu/4EouWmLgV6gCzX2dagbaSTFCQ0RKfxjFLJnLFr8fycrkMYaTYYlWqX8
6z5aEKGUtSvg3sTJN/+0lu33/QT74EmsD6avMLB+54uwY8NmO+VMz9xM5IE+
+Wle2XfgKzr3LCm6JhRl8y1N2LJxS7dIFtqOIKJfelVgLEiiyIv36uQvKhXP
cvp8Y3NaB+nicq2JH9k1sptB9ML04OurlYitVKiDACTt0nkAjXLmf3dGeCCD
FpL/R4l4iKWr0LCTkhSDU4PN7bQZs/AZLdadpH3rd0p/C7B3faa0UozPGeDt
32+/g+iShgvrCNMKmoyGyomXROn9BMuKL7lW+6Q6poZm/Zr5yh2+Am7J/Tuz
kSJqG6lDfsYN/DtJtfxAE1lhOUmL9xry3XyoVM6uTrxJGJr6tuQTSna5waCp
jsDhzNUIQ4/lSh1+yPzjDx+gsSZaHfwTySlYPIkiKsmqiFPSOaOA42HqpqFb
Bt0NXPJGzAK4+02Hp0yU09FON9QvRL/+0ejEH3mWmxvq8AaN4y/fm1anrl2i
usJGNDZn8taAAbPTxtnGJUc2zuL9MMYAYIbgEw5P9RwEu4VMmYr4Q4QtZ00s
MYHNqnS6QzoIELU50jhwdQnpxbB7kcuAMtkUN3jYaqkIzFBHxvi5uMarBfLA
kPDcAYhxhd68Ekbb0ns6Sh/weLuUEyvAOw3tB/DM6WX2js1VOZF5nULPP5uN
SWx2ZLNCJA4vACA9myrIs+/+fsuNbH5VWjbljfqv+qSNXg7L6DTVyAB8n4yl
v9UBlG+ns05JPgGL8xurUvzZZnP2stwIXW7lAvHlPOAyOZdCdDK5rAlEJO/J
jZD31a9bGhSzdlCjqeSLmC+7c9GSafeGBV2myWoDEn0z0Wiytrdjzo5YaiCP
Z/1ByZvAoCIWCdZCmA6szx/zuq3zNuNbQgcaUmSn7BcvQkfg0I3XFOggGk2K
KvE6PDVqIuEjk7a64dZS50R/OqS1T9MS5Uv4CvRWlN6pH3w6hdnqwfgQ3h4b
SoYToJStyJv/qvDbkT9+NpMuScCELMe7FUpquXlpawFT1jJc8sus8J0Q9SpD
MaLLL3p6J/YZX3uhUWFCbywTQISdRKFhGu9uSF2ZSdcvOL48MNqYdut2o6ME
Bxjm414kyN+VBuutQ5ePT6H0BSrdg3yBznCvS5d34JD4O59Fj386UyZ5yyWC
V7CbitL1XfDD+O1TrinvE4v6hHBIJthBcNqhMDjuDeUZGjB4kKkszcK82u29
dkk8WKdBG9UYXUD1ECR/KS2nKgFcPrLlEg40VO/HFMKEcrP8+kr0EGStquUV
9mmsFccnktdbuw8n3aUM5cSG4gyjWRBPsfcb2tXZSjxzLitz5i70DhrZQvcf
hZKCaQjcLLz9DBQO0106APbr1Y4qN4ZrvAY4gXjlP1MEiJM4Ad9TExhMp7JP
GyR/+qB7rjJtkYgcm4rInpp9tsvQgM2OPFf9yxYxaCtmV4uQhCn4IoGR9Dnh
xykKqWWdN7Y8eN8fD2FxiodmCbP9oXUJBqjVZwL6yBy6VobdMIZ3vLRcD088
vTetov0ECIa7Dg2kppiG3X/Yi/YI2Q4zWyxxzyorDKUCXTVkxZF/Kap5qRbH
7+kNDXssHF+goA2WwfMPCpu48lt/xiMrbRrJv1Zcw3IdyxI62B6x2vPoUAn/
onA0xNXBGEcZ0n30zL8H0F59C5aeRoP9WYYUsHVoG/AhznR5nS2bHL7lbr+U
3zRGW3NR8yb4cXfHadXUhk7+A85aFSu5hwSXTHvOLOYTMygi/2eCBrTF7fvl
jYP04SOC6lOwLBuMYVdlUbiHxxhNFG2nnfZ49Gmkf1FVy6san+pQU9Zp1Z7a
tvRaQg42QkVEZmX9Zu17P4pjSiKK2nYHF/fY9mzjiyM8bUbnz/riRG3L/ciY
9VpkdVH6xfV7e1+YLnX3/cgnfUVU8/2Z1hmNfCZHaCfjasv9FS2gTIs1xCC1
0wcFGyWJQ231PK9IpYZFeCvM35SbH0FkkTsIys5PFeKZJzf2sDTg5IB7lren
I92MxxQRqRhQDFkh2AHIXklSxODwkFs7diHI2mRj2nxITgGuSawfuZbPa5iU
+ogPKeZaoLCaTottBhTgc+DPkqJASBeZQezzSKjEV8zSto34yYQNhoqsHRk0
WBQ5KlLGn/gfAV54hCDK7Ftto3MakEqBLNkCVyz2/fjysvs/j9oOz7ZnpXrK
wQ9lyY1FmwenWzcSD36qFDaRP35793va70mdqd/dTxzIklqDquf5BhXJ3M+/
tC4/tgRxT2QwZ6eTo4PzMMJfsMeZRhuey+sa3GEteewZobxSqIBsoO30XmMM
9RT82L/QnOrDC5gQQlm/ka4plduO+8uBqtObzc+7tLtRQHGxMJqL6f8iDukH
CVU4BJfANttElqOswRmUjpZ92FqNB4qr0OA9XR2JTcVPWiyu12OWphGwCHKG
vUVvVtOx7+l6KKAXHr6kRGs6FG/UVSvbBILhYbhpwDEpLRPND6vQ+rvod18j
MA+noENrVe66cX8djY18dywmDVB0y4J/KyKvpWkfiH19wlGyK0fuLMZ188fr
XmkaR7hnEemnSSOBiJj+8cggcRBR+5jnr+pnUobYrrG8XHFcK7L3PpWbeCJP
kQRvc8gIwr93e9SyQ2ZCqgLTj2V/L/8cbzTjVoXEMtn71jfrF3L/YRbpLIFQ
0fWdRxBAkGI3Ls9RuMeI3iaeOUe6bA94MzESYtpNOV6cz3tKpZEyLs1SB1gX
FUMQTdaE5N4R+cxYbe/d86kI3S9mz9Hf0LtNZg7NhYzfQ1GlVAmbQBbHxSxi
Tl0t1rZ5wPlwePbgrHKxNRaVvvpjs2j5eeMPSkepprkOWnf72GRIBkWz4p0E
hxO8Wv1M7r4dBlzDlh+OZFmhH9DGsj1vibjeiMVb9LWjSiA6lbsCKsf7fov8
6eQyVF/uv21Q7Bj2Y0+y+f4/UfcOgqj3B9zYkMbB0f9KcMHFLOEG+bnoZuto
twUnb4HgAq34E+w8mP1pko0OAVEAPpI3Q3yd+2DTc5hv5B1PnM9Nx0I8TG0g
DCFFAF95zLuPLBhwvv14A5fy7Js89rHNzfrGvV/ODy2nVMV3shrAl/UT5hD7
nqp4tDmQMhHrccBfVXvUneOShEoEWmoK0gkQnSsB+3kvNwhMARdSifs/xIkO
Z9cSmWMQMFNzHBcQtsUyyhhvocX9UYRegVmRSemtlPdh2xX8Y8Dstn/vbQ4q
6bDXEGCZ/Nvj12xiDLEHUz86kC2tkFOTJ7tdfpu9tZZnP5wevp/J2y8bNneb
PSe3eCZH2/kE3YLbA4lX+azt63tLRR4ktdMBrdCVWcvV0Z3UBm1A2bKQNmW1
dtA5NUfPoihlSX7p/PlLSMumomQOVTIt5k0+cZHXdDBEUltvri874WNLbeqO
5kqDTPl8HefUoq/ykXBV4hEEc5kB9kzhRLYeNIsj4TLdCsaxjNqL1idfthVc
5KkTTKzbeUkPSbam967e2Cm3FCKFM3OBcOIh69ta1l/5km0yqAbVZ/wGCqWk
NrgQD0NFDcoz0x5uUmS+6KQZFymh8rSYSsRVvxqrVkQX/37oegeKQ4Gei4Rc
/wZVv0s5UtH0WbJcdwet4flXWSeLP3hlUYaYSwM+dG+KaCw+3AJW8de+YOve
xL3Zv3S1cZ2m7e31HEN2JkmOvCm1SYExQHqZ76CzsNZa+5TKeqdVzl9zeIUA
aqk0vMXLAR0CIYAd9lZ42hti+7BuyKDcMx2/XXhYIMt6/j6/nROgYsB/g4eX
gul+AnpkMAAfuOWAmuDxM649uM8AVIkAY32ivyk+WEXF+xaGr8LbAumOb47c
rvl4AX14ae9s9ZB2UJT7OTrt2J23Y4I8tB9qq9fX7rgTqkq0IMUeg1ILyLlH
nRKlK2z32YhUrK9MJFYUt5OLfR4c5WbpMdtOHhJRjUmKyAhB+2eFEef6Sek2
CYfKzIXRNqKUBRCF87QxaAH+5LfRq4tdrBa/7HlQYUDBTUNsc9yo3HfhgT/h
i7jYow4339wEL1NRzXNCbnuTrCG6MaGSnBtuB3iK4sf6X7sw0BpAKRU3jkd8
eKG70Fa++PZNzADjCX5He2RXprHzCaG09ZIahnVkIICBKo+ToaV0QoN447FQ
6ZcB7XwnoHYIa5i5oppsHLzM/dnzeRIFRPnlZW9CQkR5HTi3JYIywc4nMEQL
OZBC73DIWiB+fPXF/wl/Kpm9oVZg5mupYTyy0UkAm2JlTX3o4HYXKaWaI3Wo
FtetTPsdhjrwpCer9TdMsbuQb+g63PqNcfMW3B2RGPy9gubLMuZeLnyFjpFq
Yii/NkOf5C+VzHJ5BjaOl/yM/yqFiw5Z40pNJrhoLt1shzY5fLsOan8vokEF
E22CdMXVwGMdrIVHWD8YsOZQEz/Nht3u7rFtU49iytzggFXCgcT2emcRPA+G
PVhuWMYJrscxoX2bSGcqJnXy3UbxkDdZQ2XbQEfVcCilCSBhBVfvDo04Y/WF
cFfUGevaQaJSJi6XrquDWo+HWh8y4Y7L1ylT0jkn2FG6WLu/S25Omq+zsJhJ
kvt0bK8nYmyk4N4y2laPYpqS+HW2OrOn6BDFSKX6ruquk+oquQIQA38x4/Ng
TAPlcJJxEVo49KqA2M50jWjkZ7cTFW0A9ckufpJ37GoRGdSQuvktopCbu3D1
d0ywgJz28jzr8L8ihWZJbQ02diBJBoD8c2PbkPevbqTj6X0NMk5emfBRRQO2
pWSf2g5AOxO3ZgIKIZHues5Z3Y41MeeCFBs6qWPufodBPHfIvok6YmstCy5/
Fik2G59BX2hIO26iESYxNpQydp/KCDny1YzzwjmqvyKlmidX4r/4aLy5D8cq
hdJthpVQIU0UWwuHADJCZ/XEue7hA1M/sUB3bcOLacdmD3DBNHzFM/AsK34i
tIMvDozheLYZL/sxhhHP02paMwoezj2frPxyyqK3RtuPpxbQtnE6xw4AgEAr
8b3ARZ1zYMRFrDV11rF9IxbEsoysUDNRftG4zIyHzv5IaiahxKF4Whvhp17k
Aa1K1n1fWk27NQn49MLz82wU6TG/sJubU3x/qt5tfMykfhLGcXdHfhcNlogv
aA/bh8YUiI8wPS2ylC99GV3ox9zKTt5WLpWf/IRN0J773UG+fjV44ExVylzD
9ooIUlVxy6rT4Jk5UjIm0cecHWgzgxugHX5Ti0kjHZ9EN6EAVjxely9g6Ohv
6Z1NKzQaKBoWVPZe/FkXqWWKawXisT2d4Q1XajcoC16hor8QLvz05GEC6GbB
qAeyjJLIyCVU9Wgav7Kzp3JUT5upVqk7TFfRvAWUR9RHJyrvGwiSJQf0T60m
ImYbsYAYpD603CYL5WMDYm5e2JaFEuF7UHf19fQRkD6PX0dfDgmxsaNi4N0D
tztGZENfwO7/UnUeLVfBXRDSEN2hWdOyf14DccSI6H1qO+ZVN5Nh3ZkEPGxe
TtW0bmtSi5kroGVsO6poQSbUsdETPx4eG0UG2lmAasOp4MSpCOrOhYpVDq81
JkKlOViU7b8eCjzl9NUiDxf3nnYAfFVwpmx6SJrL6gjP3sScH2PNt57gUfVE
SviDgo+iz1lkoZ92YwmHIcp/IxDUumr5U89OudlhQOwoqmnGI5y1PfUknKeC
4lL2I6oAmtw126Qbo89Ur/vFecsYw9jG2a5sP9hgJ1DjRCE69Zs01jQADhtk
9js8oeOIDfheca+kVSAeChSs61xgfb0tRAJL86Oi45emUpu+bsd9a4+F9kLN
4sAZPJsLVJYJmhFzayzzpe/dzbdDJc/RPg2xH8fNjzmk5HvjUHfmv27soFTv
g4ekzOj40ik2LOtvxRQb4Z2gm4x8qKjzyXj8/F8PQKrQH1XRwjUsVu0tsSZZ
ys1HpJ6ahRxFssDKgl4bbFjH9cS+1OnW+lPyz7oDM/Bj3U0ljh1lgjRGTXGe
wgLwoTgWSD6vHXoqQFi5mB5w9ybhexuQV8Ypp9lbxmT9M1E2Qbpm4mLtHa3B
OSDnLCH7QxyDq6aEcR5gtLfnxBbNRjR9Ftr2XDVr2TuqOEgrGv5Ka85Q6L/L
+b6RbsQV/lisrMAorjxZazF/tqqRPKHHbqztOSD6Z7PpIPRH4gkXBxNjNXqH
cIwdUuNdIOLjbgifLYULpylRczNTUPDWa5OWBoKSYhhC6HyBtnfw9xzMhU66
FlEoRkuwmsC0K6hYAEtN0xT2lWzbRCigz00xFUhz6wJxjVgKy0E4fNjS2b4j
OxkQUsP+s4KPq9+K+BLQNQud/HfzP7d/QyosDZcUqMIojhKB7R83kiEkW42o
3JF7QwBYctvl529VkFre0YW51xFcjM99fxGTy/0ecsloA/gtfBTo1F/SZ8Hv
beEf+rLuxumrxDSMD4xOG3mHClVZ83T+dXY54E881dB3UTW8KppoUgUfpMEm
Ixh7zkDBV8P+3ddtT/Xx1BqJaltwjg2Pt06+ooo3hyd9vdVClC2bbHvSk3qx
/8X9+6K9AtHvyzT5t+3A/U1ceZ8FB+BQwi2hYDijNbTE/1mVSjnqQj5yXif8
vQSXtFfwIACyZ0xpvjLT1/MhnmKF7niXLQcTpvhS7tEQ+rztmyqjVOv8AeGz
e3hqjGyXEHbOKOzKCz7nMRm3OIuEub9Texqx+xgj0J3YRuKmP0pf7m11l9BK
eTEOkidWAtZhZlccWDhKmdF/fOxLsymBoBLSjwB+APhMMLizpwfq8kWKHmWw
sIE+o0iSBw3VbB1kURNcOzv7LFjPwwSnOjUPDWaXRcNmDOWTxOSFnOegjq7A
5E3AbxXxZy3g+Baf7efRfNTFDZxWcfL9pXAJRnNbt1u/SDwtz+jZyxblFBfL
TFfyUWP+N+fGj7ckYrfRNZDLYFD5+WVyoJGHGVTL9a2kDxaBCtB8oryRGIuv
DN5Q3t/q2eCWgsV4KxAxse0wMsTh+fNt5IZ4Z6VeB2z5mYS11sVlvkkVN0WW
1wYbHAz8sxGvF/TetLJwfnI5dXcxyqfzRwnaq+eeYcCK92Hl9uVSQfr6DRXy
tjF9UH99+XnLh5EhY5A9+1/xrImn1x+igFgR4Q/IrOb3ENCv4wdausBZ6QYp
KXrjKBue/7ASfu5bx30/u8O+CLgi/qyyHVHLTz9DnSWbZ27t34p85K+vvoKl
YYddhS+T3pWnyfw5rMgPyhvAL+ax3WD9aEcqrejlK3q7OcJX7VWcEjHhuFNt
9+MzTpX69eM5rYqkAYfIbQRzV8+UGetb/mL1pfDmAuIhqOj9zgBw85r50hGq
Py3TdYX3dUko66fIlb22vnWvggGP8wrnfjezlFCBy2LvUF8b+8O6jg1QbL6y
S4qv4xSWrr2M62vGSXVEbR1hGRHRMKn1hdrXC+eRqyFE6JQiMo8M0kN4NScR
YqCFY6B/08s8/RFPckcanPyChFtLOfMIXGhEz0eirT82aFKsiSkpHfsphiyD
Wi1Jlnz0dunM0OTKf1I98ck9vAPAKQXx37rwh2gpD0kUTc31VqVNb5l/125i
fePrRMRL2qwtQzOr0GAGLfnnNSNye8SlzKpOqj5dHKfrzIjCYg0pPYpuKN6D
wOhsny69wtuBpgJYRRJ3N0RadOAY9mJWf+zbn7sTG5xJrC4SKkc36NNm4O+e
/zsJLudFe+LXr0JYIqaCKP4FpQ4Dylm/d34E5OUeBT3EYbkEznq7NeJ/uN5X
IvB87GPtupzbPBUAdUzC3UevqIWkyPnTrylrZAavI5fasMVJyQ4f7uZgY7tQ
Stlrsu2essnF0VaNThzLy07EvbixxwbLH+N/p4xCNiVC5lQ5/feZHwUFX9LJ
BJnizI2pH1M/480zzGSAelvFEgsRQkLsOcfz4Qa2XEt3b1cGBfhnaCajmsXF
C3z3YDfFvz4vtS1ZRj8uITZzmiSbUNZRciyGFsnaSWiok5oTMzdzEHYzXZCX
hxBvfR+m+8cATnOLNlRwXL9UdTXdtqH8xT/GT7hR0h7c81N+UiKRqEoNESm7
V9Kww3x1caUqTr0L+XNMIpTrFm/TOdoVQtRAmiXXX2rbA1Umb58nQs8/K7Rb
GxrPNt8HOfAdsIv0L/5J9MwWTMNJQqlWo2PwNJvu7GQMIT5xaVzGtNkBeBdG
xi2ABBLhrt0zOaDNeE5c0q95U+sXqhgds2FekgVTs4+uetFoxlls3NJN1s3Q
7AyMMjdC3lP/vrzbLXG0JAzRTk54GOSMhsoyKIgr7fZxOQBmc4uM2KS0shbN
CMThnBQvzkron/Bck9aYMz6T1QTBb2yyTwXctqhi8EVHlhryPotr4VPENKvD
z3HRy1NuV080QHc9MbjpJYT4GHJFw2RcxJRuClWWRpFOhHrymPX02/YlA4kt
xcNQ7twp2icl5jWBFE0EHtv7H857Gggln4a+GpGmcDQM0duoj60WmKeAXqBe
2GRChPpOSfyKiVR4x3vHUVgFDeDFpuje1umBL4RTVQZGSu87sRO6LBFRMVkg
b9AnQFALg3/6sSMqtmRJF2VgnkYJmE/PKxMuXSiBDQbhF5WFOb3ajYTzqDn/
h8QgQ5nGEdmbt1ISgxwdOhwj778eTT31WGaF2U58Tj6o9GJ85RHPCz/arn1k
V+pfwjek3e58CYjB7ujkvA61ykzC030qtdXnmYnBj5zLN3a39Kigocsn5LoN
R7LMZ0h+h1/+/2+eA+97EJkd0JmJblavcpNWMEPgkmuVCXf6NdAHsF/4eP1U
IO6r5A4n85n16zoR9BJpEMJz1h2u+TiePe+ClHW0zMyQs+uB82PvvtqAIylD
Al+e/cVovgHXkI8p4QfHX9L05xi6k7qXmqBTZM6WcN6VnYtuv85t/F2Ay52M
fi7/qxkX4I/FkHrp7CXLpDuj8HxXFHp2uMmuqL1K+LK3cCsxON+ew4yNN968
XB7YNa2Stu73DaAlzdQ3Y16qtpnKGI6EgqjkzcqnkHHrY1pPzzHvVnE8YgKR
diQ4vYe7Vyt3eIa0LmvApLSlk3jVouOW3RiT2/iYmqU/RhfZ7lwDbghHvjAx
aX5IYh8+tixsUKknf6+MR6F0fELoxv2hVMQxtan232qRajhMwr+D1mEX3HCO
6uQy0cM36DYpE49ZVPwN/BuXliRMQNxhUruyUhdsxn11EASQ/BDecy9XivUi
6CEjxS7HdSfYExWZSOy8CTWDO4jeCUvNqpP8fU0JPSPoTDIl6ciakz/I3QJD
c9uoXMrdchrK0xhTFLYhduBFP0XLQqcvKneLKTE7Hc3VsG/PxzhMmMGRopr4
kWyDbQtP0q6UquUDk6UH9ROXeTBmLLD2x0KA0KJ2jf8RqjyOMEVeAZECBL3J
cVVdPW+QVX2A2Gm3bRQpo2EHWduk02gyCpNh1LT0zQSrfjZfaV6egYLCkSgc
nJ+hy2W0rTXy0PjFaVeYyDefMJM+gJzxV//BrZXf9UeCRmVxy9CMN33RIr/V
KKBJbZgalU4WIwpCsOOFxwCxSwqel9kDApIgZI9YwYhi3LJBC0XiEKK71YcN
1XUStBVI3YEpE9Tq8fgpda56LRt1ainfal/UVPxEXgo8fTOotlUdF2EnrMnZ
kQTyqIMRjYni9yU+2n1qB/pmRWkG3D+Fk4wkyjsqZIr6LDKQzB2+Ecjxk0us
fRWv2niJ9ZFkfoMcvViykTv4U0gapORoguFX1rXWQCfz43YmQApE0DR9+y/R
riRxcB9dEV0hhpbK///87DzSEkfM+5YX7gazwvWdDQmb7ETGbE39xi78v+ax
Vklqz1FHLMsUXu/j5PDH//cIr42uCWRDR9h/H5J2O9V1dKhxQsANiO0xvgO+
KHSDP70fffHTp/Cykmgush6jVHGo9mzNcC3a+/lqg+LD0xZRNX6rHnnBT1Jm
y6TP7IglX2LGxjZPMWuxEew5O7NZKh5c0uGnSnUX1B8SYKOew+ns3//p+BrY
l62eON4uDT0DuD4pIAoSky+d3kPA+G4edyoowNsT4GlXpwHCw0Dbaacm7hLr
sIQoxH0Za2NMGKv7KdmISKXO08LKKNi/ekwx5TYPkEI1UbcjorH9LOAoNTgh
m28hgkzM3u7qMP4wGsq75aIxgqJif7EzAEkOw28HS4J7e74usTIUPqm4y4cY
Xh3MrgqHxZggpHe18HqISKPCBJxVkuZA0SsZEZUD3rzDaVIa2wz+OTxYnHnh
Lzf4U6Lhs1GePX42rriYObwUA+Uu3+Q1dNrU9Yqmw5h6BazEU43M1WXL9Frx
mZNoC3efbVtNhaJKsvH4g7PamJ/kTyggIHZuER8Hx1S31s4YRdp1hS6h1ytw
LRD6mYP5akRdXKbiKGg9ntyrlA7y73BVaQhG3vnGjO2RRXJtPj1+SRJkgdD1
KvFTBO+8z0HS1NmW5GgKHJ/E5Mr+pD9eYZNOGTCdusXojCkms8tqgLn6IxXc
35oPficbBBVmT0cvGoso6A3+jRdO3ZqJkIksEzT7xsbUGtbtgnTeiKU7C78Z
iSmMmQoK1lG0mVaNY4mH0fIioO0nvzHUyZ8VM1ObdlSP12YmNeLbi7ArzEmB
xeb2S1vcONBrmp0bnjdL/W926Njhb8prxST0FRTozgH3EMgNIsPs53IF/rno
/bJa7Lerhn8al5qqUzLxR/IYDtZTGcvV94uFKdkmhqHL9EIKfmoAkTiKHgCW
wE7J02BnwPlBgpDFMERhruWW2QHyOHGMoSmmCP8JOzIppzo2T8YjFMmfEsS/
nlFH2z7C9oPffxdzy2d73ky0jyENWdCsDg8XY5ST5hsZnIFlYDLxWxjV2vHS
xcbwxxvlN/k4bKZr1H93Ro4i7rOjEW3kfFh6cSoTb7VXX+/3JC4BwzVV5Afm
QDYQ5G1cEY9ZV6OzQhw3yt7YZUop45sJJwSfqMpRgOwfucoAUMG9T3j6qLQT
icHUsLvz/53sX4ffvm62i+x8sh99JqN2EkwbgB9uQG4alaKWVgnlctU8ClCg
/7++uSwIjG6l7LUMiZn7gsPOeVPeRLuVlcg07YMkuBuv+gssnJzGc38TxqTd
+5imToum1qNe+5j8eT/wnzyrc+E0CypjeNNKgd6G0wocG0JjL5bn+6eNQ1ms
Utw1FqITneoJvw4FaG+Dt3Nk20G46jZlUQPdAXPxz+pknA06NeRKnTcTpwkc
B6dXonITK0DvVuN14obLw290CMP5jnKa9j8xDT7Eb1pV+YkMcaL6CDtJCdCO
icyKvUKDgTtcBGbkgbcCX9qNBTHUvAadlfTA237/ujRJDiCzxSnssHzbEaz3
nwpQRmlXsqE7AjbxmI616VztK2H8NIVb1D4HruhmQNxE6Ayfc2AB3yST/P9q
0U00XyQ/92aklvmls2/1B2769NSSh7REModEuOvhrcWpisGr7jmlQXeOUAGv
zqbbm0geoHaIs0xKAG3WDXb6ItHVRc+XFCkKTkHDiAfc3GSTRqiov4i816Gq
AsavNXt8PmAZ/dxSnnREorEyyJI5z9ehDF3rVqUDZg/ZZ+V1GCGoybnNyQTy
TA7Fd4GizGD2qTSVoJOa3Q90iFO9BkOaaXTv9/+D1iMzQ/iKZmzFOOj948YD
H6kq9dUk/KVec/KQRXBDqIME7CHAzuzAvaw67l5cHRwwB80Mq9Mpwa/EOoVe
vFGg4UokuRH41BWwhI+JfDaR2J//Fjtv/Am3D9Hg7r7DN4iBxUUq1OywZJjJ
Hb3IweJYU1OKeflAARKZwtS42BPwK3c70Fc28iMwgk60z0uFnqLEagI74HZH
o/2UCVG5Hln1O4FJGHYXa889jFjbTRZ5CbyjDE5udX5rOnhN1qB9VHE4gM9b
T2qoqeCM5Li+N6zHVBSFSZxKyVlZV0TZufQ5WT4m+RRwk9rkNgk0wWhRIIJ1
WjluVy+Uo6/AeS41DpjI5OQ+yfcvtewieO4jqmKZVRLUoXcaRecXdX3upstn
Yi0NesSmguj0NU2xmtTWCK0s0SVA3hLt8dR7rZSEEGEGVsCVoPnGng7DdsHO
zmUXvATHxVkje8GZhmQyBxoUTor4ZH/Qunk7rqrCt5PRKseBkAPnqzMdDorI
tG+ewdRVJ3VP4H2kaFPqEK7LIJDdQOXtJId6+ytARjscs4sS6yR/KnlAGWjK
yw4w5/BMuvKKf1nC5TCAIIjO/gDcEakSxjgTfhMdgcFBTE5IignzWYDBPMgw
Cw8PAtigt0s1lruIx5FGcluvTmwLWZ9dPeZodZU9P82uUfSUfgTHcKIds0uI
42GKrBFOxo0Sf5syHYs/9P9rtxrLFq8/Xrfqwcl8INoolwl4CU4TmOQ8r5xr
keDaTzowOe8oaBoX6i9MwcjcXLVL1NsytzhOz9BPhBzXJuTW+pkaOfNH40+s
uoMh79oR4r8m91tvxCZ9xrX1celOZk5PSOk7jHs87VsY2J2wSOEUVmJ8jVu+
2p9J8/EXqaewCPCeR4NF2brNJRmbqBFAOf0qw4SUYxlE8onynIsKRZC6fdrg
lTSghhpEvNTOOLBhgUIm++i5ve+B37WSapbXDMZeiwdtokXPSd1bcFG0jXVO
g79DC2YgkaVDrEfSoxPBmJZxVv1t6H1cWx3nPprGt9YdS50ADhHGyxdI0tNM
HaBF5d8mIU4YkUbGNtdOBLvF2RGo5mEbMbRXOR/bto+pE05OZKDi/wo1H0wc
KQp5gINWW4R+yV2V+X3otOU8YcSJTV+f7dGS1Ayg9l+XgjfU1MMQ4ZEoMYg6
TSnyxPsjGn0Aj4gIp9SKFO6IljKuyxyMMC/8hctvKp99+HDJ7S3S0XgaBLEU
EEzQca8CgSYrCgTiRBg3wQN4vwEyytH6HWMN0KNxOUMTD+7EHGuRUdJKWWT2
wUJnYP7pjFkt4YR8OxdYOQlUSgZkfWCBMhAFPq/VcnrufCNiUKGq7roYqp54
ngKEout7IDKhesk7T9xNeZQWftsPeELsm1S7IwhPdNwdrllWTDO+Umhy6DWo
+8ft0c+dv0NfG0xYYsyO5XBXF6eDRXkA5g1NUPxoJSivt8fXnMLzHqAqkyTH
xZVZA7TppFgvDWYccNxGHpERFw2TXoBE4Cyiidv2uzw1wEub1f8+XAPmVoPC
vcebFKZkeJtBp/cW86x+0Qe5AlJ/8hGjk7NhyveA8/UEftmsZZHwB9pMn/sK
nSuvtBr4wg+ZNesQApaR3x6NGDTt5BcJTgRKIiaiw17GPAwglxv2kHFhThYs
W7D8qbqEADkCYVerEA4bEvYMQ5ib7j7hF/RJYn3mQ8XxucsoIlwb9GCjlhVc
qBR/asky9m4s9sA+6upG/xkNbnewvV6w6q+DQmKwzR0R0/FDEB26InRSZNiZ
X7fzbVii1BS7mC/nxr95CcDMCeEdJxW3wefm3gvep3wwYBqvHT11iP4V/9n8
n6L3890a7aSe/nPj9RlIK2p+IDCkajD7wUs5ZjbB/l0nYrRtluluZCE9kbpG
PmLLVcYkgAoyO+9O7aJsKEOe9wFsrvr9HbgxXv+4E/Yk+gRskp8AyU6pRkVc
fUxW6+OPGHdULzu3V+hMkBtX1VuCxKl3Dpn1AdSfgv8nxt1V/4fd+v4yOedA
8y40I1Ol6tCK1xM/p3Ko75QzeMAfCGfwwWkc+OYJ+hE/nmY4x0yJilRYiyUB
4F2gDijxkQE038CPWQeGP3i4H2BvTeF+zQj6rFgPmWtB71BmRSWBFXQ/BTzQ
gsWpq5xQ0p636uZQfDE47rtfcZFqTEwhYcfRfQFwCaZzCIIui9yT5l/4dNtI
M0al8sO1+N8RFBNvTssu8vxIz6pfjOkupx3tfPM80wyxRO0SUlZwZO36xNkq
C8WYaYypdlXUd3MQKB/LEzZNs7nhUnezW4Xj430WArtiunGpAmHvTYpYRax1
3ifaq5Q9uw1W9Kdf+Rxmu2nh3zqon14pMy+1arV4IJItI/BrsbBUMXBdvR2g
AIASrJTpzK0+SxN1DmG+/UIpvDlKptbXCQk2olOYi61Pbg/h2tkEcqpVfpto
l0t5AlUb5r5aQKR728WKoKeibMHW5wSb0VIvludzpzjJPZ6Br7xpHtA0gzhH
DtIpHta+LJMgruBdMK6DIMw7FHVn8ENfnaoU/yQ7ntIrW1Vm+5xZ+nNNZCIn
r7SKrwnRTxwgQExz10aB4q8PgEliftHtqPS0+kPdrQ8HqPpZ+VPLHm5cISPh
2vfHBE2wQrfX7eYKiUeS8cMkg9eABRnpEeM1BMkvW1scdJJO0GtRKsxC1Hbp
ijN43NSWL60AYcxDn5sRjlYGmZav1uBO7UwfG03EB02cbXwhT690qnngI1mX
7+v/xmUha3LJIFaggoQGmJpLEAW07D+59tIoOX2eU0bhi7RznHlutbEdmTLj
7PEK1Cm/QEIMTp4Lp166CpTr5oV6nSHYNO/a+m2JBqpR2yU+qJ9r7+OCp5jW
HZuDQ4E1AilXwpEsSfm8aRARdiBcXnXSQi9r+EdZ25FOSfVdShm3PwlYYSEr
yxicy33+vkXUFz3OSYs6GtnjZgEa5lcyC4gqTkguJ5885qLB83I/T2kihg9z
U3S7/2zvpSV+OlHSAws+PHX0IdtGmVJA3SNNWwM6HvDNDAqlmqA01in9m8Y1
jfNP3+rAztJssbTZdbhM8Hm5dYIJfwUrz+irXsFoRYe3arbUupHMhzu6oIxd
8mdIXyHYO1QcPd9fnoNGD47ilATvlxzA8rp7UtDA7WNDQP4Dd8k76oX1q3x/
yBLoUgq9jUGMmDvlNuuC7k7v2X1ihy/zZqsTzikq3FZYXvmYByjHj+KjykVP
JFEMLJm7sEAhfsF/TOMyVlfhD5NzRD4a8/uBXwArn/sfZzP5iihp1yddAE8P
l9i4mqkJlZ1arPwjcyjQl1UnAoA5OIA6KPK6UBMA2FSXDAE85dJmRblJgN31
Pe5znLjVIYsWPQnDeHSColz9JM7YJ0WLYj1DEziVWVLnWr8kTAiYLvq6POcZ
G/rIEdYSdUv7wQeXQmnbWWKbeilwj8nQ8jaootPOvWB5ntW+rDvUX4bjh2r0
zpTDOZ0dK0WtJDDCvCNqyhX1xWkTdThLolYJO52l5F0l5rWb+CZOGvcCNHJd
Ugt4KPIkY1UGJOdS4Y+TfXTjGm7+hfpKKOa8qXHeE0y/meGLqvUPxtYMv0Ju
LQBuJ3rbYLyS4OYLThOmXJlhJC7t+Cs1OLo7Fo9e2OaH5ZwOFCZsU2YX5ncI
aB4Lb7TeAUKRNpz2Ekpuze3gH8RTjayfMV2dBmHDioho+PJ/EeWsB8j+4ho6
2Ktr2ywrsVmild6Ne7R2WzNmm6ii+8hgf/s6Qe9HsrVbu/0PblbvCezP3QES
xDbLk8sAjEg88utSuA9Fo622czLC8hF5Us2z2LdKNo+PbvJZyLTRaqd9VqIB
xsO5KIIOvmVyPF75BzDHa3G/eEVh6Vz88tUnoCTKgDJtLblKelcJFgemR5HJ
xIi/ejVlZIztyt84Ok4XGsYhXiQSxqnYyUD1xIUXRBpVbyNRIRdRudldMkKY
SbI2yoZ3sVTviJYjnR1dcnYfFZnLLFohnN62UKzppm0Y574NFVy6XhV6Kx5i
zJ1cwojKRHtAN/b+L+0/sX0n20Bky+1/UZNV1kd3UjaF4UB/lcw9UZpi+g7q
shQKD88eugTMGK4mqOPVAcEXB//H5HQDVnlPJOWCFYeoFKaaP6lbjKdgsXw5
IGoawrfp/jDY8T8q7nsNbOE5tpkuTW6oDDVqsasrrtZTA7EI8E3pmToLZTmX
409KdicCdnGE2IeyBxsMjSe3s/L7vQ5lygn5PHRabTUG1W0EnLdPxO9E5G4w
wDCcnixheuUcCyctoLAwjycuE0ZUcD0AaKuqX+gpJ/ixVIcm2eyfJkf/GYzt
rkywjeEG3dB5xDE5/CjYp5P4q9aehVcZC53yXAlWt27GzVF1v3hlaaqdU0qG
l1LPYj1LM3iePjHpTjjZAKZdWlVR8ACYxkHDu77z8WHVNnmIpJoIDpFizb/1
iJuSeSQg9iGDl/CRTnzto2opCNTmAIOwb6Cv/KklcXJedbOp3/8m5wbD8GaZ
qUXOH4bkH9OBEkbUYTb2rtxMk/l2aorrTx41uCR6zPJr87kSTDt9dlVx8XIB
C5EBd1FnAuchUKZo00Jr0cz7b35QDqBKOikJC1UuIVHZhXtqSXRcZzzGiRWp
EWoCqEyee5AmJ1F1rctrVxb5k9IHt8CGifNWdd3pJIX8hQYuoGNlrym5Eh+r
I7y5aO4frfWIrB3hlGCB9CflldeM0xMX2gzJawL+VKIt3t4njWSuvC4L0yF2
RVLhvFatD/k2CkSe4XlxxCvRdyBWfmiEOMVMsBIoHiG9xn8wIgqD08RQkU47
F/h5D3IgBZTZDkPI/DsIa/efAXF9sUcYP/Q7r/HzT97ZgOua4xvBWhx2ocen
p/XLFyRT4VVDrlqxAp5+o3e2yuDGjptepeCNXZiOEL4SE8f4LXram5QRb5w0
Ucm3CdnekCcgAhLhCC03rWmKxhEQX8ep1v8zVYs+oeLqCTlLe71qxq3hIT8l
OgK+jWkNVcdAJySIrVDYNkFeFVXJOu1XqKwXd4s0OMShzIiT9P0210Pc+8EQ
rF6oOeIgMslHCxHOwPdIf87hXesAhaK9T0yrWiLazLuAw5ZAeuTSYA7F+6vi
lpB88PAhIqci9TYWlH/tU/dX2eDN87Ns0BQOwTwjqhKbcV8NV2FIAdjr4gKd
gfaCOW2GSK0C+p1iy8JF3Iz9YWH+w6c8u4UvEUPgeFWR5TN8Ak7c3MTouSAL
xr2Zb8CJS1fYd/wJa8q/ARQUbK79/PQUYuEUlzWhroil1Vz5coUQzWaZJJIf
4kgMxG6bCaYXooWMehiPeaABRh5VDFCFj69jq3OrK+U5AxE37aM9h7FF06VC
M4KkUoh1mEPUGgD04jSjbFqXvZ5HMdbcm7+5g3CEv17IXiADkFQ0vaZ3Rxqo
SIBaC4oFmMMHXdkj9h3saqZOtQJ7d7KeLgADVepFN6TrLsujOhtbAmm/R/+n
QSd/9grqj48uLcM1kq3mS5bCEecgP9bR5uU6saHKAvPhnnzvdg0OJsFxEwH7
T2XaiqLQeJZYY7myktMmckbVGnWcUN3geYs8tVrNU7qArC4VfFApNDLGVFI1
7E+BT1tUxOjjQ4s27JWmdXbhMeOAjesxwjm4UViuvAfjlcDzcq1cvzSbz8wt
ffkvHbOUWXnL3qdn5vShIzXEvRm9UcZ+yUVSOsE2EHLjIRfzXCbp4lIIhTBP
hMF94FZXqG060LdpAU8XUZTyH92O6itPBIc2m6+SkVVqAvrp//+z5X0Dvjo1
7Cetuuk0T98pnipJ6xZm2QUUC1v4ke61J5RJRoO8M8ZuzGV98gEkWYOP5AoD
zFvNrHu/PHzQC078f1SvHkqU272EYuTNiYQc9Wohu9aZ7BELpZdsRmJDeBBf
yjGSzSRhi9JpnmC9QPPXcOXXLoUfo8AUCC1pl/AeGt4q5RyYLFXwo/btWJc6
Ruuw5b9TC6vG9pLbjpTQBtqT1dx0tpVww/a77vSZccdA9kst6OKntz2jbIDV
s7sB2zOV0SHU6c/63jbkyMZiNsUq8ja1fZePsy2chREVNSGxGb0WuZFQrbbe
A2+PXKVGdBryp7bfcK6Y0CSFnp9uHN8X74yYKbT2amiKuDH5WsutTdUi4SrN
LCseXhjiWITqITNx/EO+ShE0PJLMVB5z8ToXC3g//vOYqboxKcXTRPFWJtkk
L3tpT0n8l+ABXsMIHcFDJenneBwaYy70ROVwV2yhYPbHoJCEG7p684PF3jiq
zHfIgdlDej7ywLSmXTXse30bfTbo6YgRFvDIjD0Zo/FJQZ+QN66q3Nwt07bs
yNKjUHyzR1M7MkNY/3U+y6x2TER+a/U24yHa1aAKFJHR7Icu4ffJH8lDiZVu
1/mXci+9toTG/OFhTbU4mizE9LsDyuNiCxAIC14pwNO9G+q4eS8cebBWEoh2
hL2JWQpG8PR2wKlSwDKVk5HWf/xJc3Ml+o0klga3M+H6IKfhS8aE2uxSNf3J
KUBcD+u37ReoYRLy9Dp1FXz4jW74G5/A009A65EXhEpd/Z3LyHus/vEuMVRC
zilGgCqWoUQrmYdLXp28yYDjTNioTAZzRxWatrW2JoGtb7XOFmfBgI5JQjI1
/8OhmG7qYoHJLyLaLCfanwK4h7ARyCb67dILKpBmil2r2o9R/kf/b/JrJGHZ
BuOWgnQ59qpvwDLRHi54DIwIJM8pqFUYw/i7/xKmpfVOZ7u7FSmevyB5Db3Y
Th6gB1JQaDpqt5O9RTGH9t41oMTDoSNO9Cm4NRr/I66N/RQpMmx5dFW8JBtV
XbTklKdu6qG7efP+XBORqZCfLoD1GfwRSyO43ddw+0ToVK4FU2mOpm6QL7qC
LAunrO9jHG+Aj/3EuzhlKq8f3Ay7PKrLIpWpQ3OKZ03PLqUn+Jj3MEUwHFUP
cmoNPC3q0oxlGi2CAoeGEWsg9pmrnnF92DDs3dtfFPvbAyH2KMyxRtOtU1jm
/Og+b+m4b6nbn2/WFvCTR89LtHgWIxmEAdNVTnvFcQXjr+A+Lt2jhvG8Muyq
ww+WgRrSA15TKd67smq9DwSQidbnC2pjpb9pHamFTzqkHAdrQwdv9GA3N5Q5
mePejQ2NkAjjNDIc1DWP5N4Ke7kodT+utmrKdd33gEoTx0l/l0j+enGWiOBu
ADsevKUw+A/zhql3cvEyHmRI6XYSlJulwlvb+7ImlmW6z2vF4iIzhaK0102S
k6EMYDSm8NnIjMsmKXox7EMguMn+PmPp2z1FphbfoAia222HwuDdWZQwhBSY
kwmvqZeyUuj/WDmVLG4h/vDutUVqKTQeewPXWFs2WsvviJwFWHBiPUVVcxmy
i1y4L6+CTBW3plVm6KgKFSEuIgxsolvi2s28koD103nrIQvA1qMBM1Mh+LvU
E0/gonvJLiZBTeAtIygf5E2aJnBTRfnruo0CcFC2hyYwK+Bm+YGGkZ9KJgzI
HVNW9KxGfSExbLnb1j0b4PAjAn76uFqUxM2HXOmThSmgxQoQEvEed5H5J+UQ
hIq+2HG16oyRdog/h4MOsWL9WDayo5zTxaS/xcQ9Y14qHVmj6d4UlTUYZNVz
N/MYm/nQnQzL8730zF/cqgxH+cRfBcYquZqtYREEYonAjYuBfuQm6FtImP++
TnxTduf7D3Fb3kxMB/GtEYpnKeSXxcaKHX90b/jyX7sh6kgmYYS6yq7fFyGz
5dVRfepXc3vSmOMABibKJqUTC9HbUXixH+ii8AOvORZ4OHmmTl1ksJRJ4vBa
hci3TleloNeZicFwoAU2Goxf7pcBjnqWL20oOFemvVuZCO3+mAFg3sjKjhGU
iJmoKWR3y6Wbgmxo6VhywnhMBgb/Z90eA/HS3uOVzgH2u5qe/alv5j3176rk
B6p69Bu1oYgvCZBaVVwhC2P0PTmLAoXhuApD7Ni3gfh6Duk2WAkV5p6CWz6g
3+bgpp8Rj5iWllR3hStbo3rozR9oYra4EMzlSw0caXK/qjgg2xtGSbLwddkq
RbW2zwiCxGbF9LJxx45qGZG8VSQn3anKbcT8VIkqf2s1NPqgEgbNw+8VBVvn
J8sb4RXR5s7XLzxAtzU6lhmXzmBcFngErGf7wl4ef2ZUOzox0+zXCDtZWMr2
PY9+7IqketvUvtFYsS3wDpUwG8tl1d7JauG2nFHMWk1GKRwOgiGD9V1aHwGZ
P/+OPMgmJayUi/bGHFm5FNIytfPAr8+c6uXOfRSV2zuZCMvqhtoqqeiZoh52
hNmC/QwmRTZdqfE8wNn7Y22M/pzjfqCIj467rI3BoykfOUvvHhGv4NeLUdYQ
ER9VQM8tu2M1EKC6MDUlsSzgv/3WGQwt+SlSsoI8vxs16roMhDhrmW0fse/5
XkB9rBOTu5TYRXQrwgsUlPNyX56eD5NmFZoQBoI/jKflzX6WR/EAB8jWdQd5
OgZjRc/IEFAQ6nvBi93UGnPISdD1rBGsshVn7OZgM1cczqFkjVKVgC/ORWoB
He8PTl38Z4PYT2RawAiaT5c33QlMpk5cWruzMgZmMbw/5QLLOtg9Wom/q4Mz
Fp8K1AvSqeRSe0Qn7efnqJ9QBc0qBL/L242zFv6dKEIZB6EYuCoK2VwFynKh
KyFctIc1Zqm2JkPuehluRKvklJHsHynaIpvHDknEsBmXc4MaxiZbIFPeti6A
xmsjZqiNnF5ca7laSwaJoy7oyh3OvByqHhRglA9xVJj/KRU/0PivLDHL0E3I
q/rOXN5z+U88M0i7tcpjO01gXmGIqCEOF6/ZVEx6xDTOL1ep6Aq0q7c1NHWt
mB8qdU2UQMinatEJMZYfZG1CiCIxR/1/lfRuCIZBg13X0zlT5ivht3zKXnle
+BQCM+mxBNhfYpXW6L+MflqO5yjX9Tx43jlK7n1xU7oMIoKOmJyiYPkBvLNM
NaWs0X7a7UptlypG3ipd6ZPtxDix2bRHtLACAg64dvYNZEU59zbkZQsSLPnh
FcbCnUwEMSM4Fatu5/G66tmWFFW5l1YWBUlXk8FCsryjJ9ecxvQZhz1p13+B
bpOYFBe/IRZ1+8nN8AlppKWyPbi+iPyjrj6iFCWZLQE8npchA/HGnhNQulMs
BO4NhMcNbCmNUuA3lVh5qAJ4ujj2ujNqxShvshPb7Br66SYENFvG73gVCHDI
kAOdx9xUrpP1PBT7OErkrny46f+uFoePhMvq+7ByLnxicIUfAcCBExdJPvfS
PlAoTOOQi1p1nco0xLe3IFjhP0vK6uLiP1bDwSULOVI1X254OdbbPOoedEep
UKGrQos34XoaKOjAXrxKIl5C5GXv+My/+N2Vnv85pesvPSzHkS3SUoeNvd5Z
X0frkJqCUdW5ZasstMqQ45o+jZBfdKo0xALxIvuO1kD34ZaZPtDhUYrb5dFr
0QnvBIPskgkY700l6jTt6ki9uL2o15RiDjY1qGHknoUM3o1SNMmvaAEXA3Fq
Q1bCDvA27WQ3//Xqkl3AAw2Cy8hVxNCGOfexij4x3zX+y/lYTMYxSFvE4lQV
ZZGbTJ1GOXcXnG5Ex8o07I6EkTFasHqJLP1/yYqaUbmQgOMfp4xHPwSdbGa/
qBw085dQM0Tneig4fvVnnquq/3pwZRidVlKHzpI8WNkrHulfhV0uiwbK3x+g
3ihPSG6uxOTqzSVzXF2puY2g34FXaMtg8aEQiax3jcMQteCuyk1Gyb8N9TWY
Av2eU3wQSvSv2n45OGX539ESbXBqPnhJMhbttRqv1OYKyVlzyUbPIF+hkI93
wlkoP0EGYQ+l7Dko7vCKogYi/QnwM5Re/Ulw9Fu4nQvpvyuQArl+h1J0Il4i
WrQbBenVnEhArY6AM1huTDDhh0RIMfQiSbwodiaqkqYEg09KS456ptB4G11A
TTzmklEF1QuUNc6BR1UhffW0I0rGEl9pW3F6mO1+LEZwnBFf4DLylqE4hzos
BAzzljNg4hA7fDLBHtu62gnjuggoC4X5/Zk93S89SrIiahDz7SbSYD66DY8Q
fcdZVHev34f60xleAAMBjFJ0ukwyuTvOYmw/nrWoLbttHEC0pmZyYkZbVvcC
aopF7aDE2gs/w3ohj9e0ixb4k31iG+99v29lcL6CvM6dlO5icp+Vxv/f4xTj
YWAvYAF8K2MpBLX4fTpAk7qmvWyy87a7RCn7BJ30H3nDTpfKAEpPCTjuKiUD
RJ2UKlwlqxpj0xwiRZWKL4D1d9tmfEN1S6ucagDVe8BjguYyqgL3sn4AI7hd
ZBpD3EGmTZHDnnRm62mQbQPxXQW8kpWo1/q3KIXu5JawsD5il8shvXkmGN+A
pcFxrYPm8/aiK/nfcSFWBqUzwpKJCISSh4B/egfcyKTpbf4kHv/ZkH/t+SMv
JkPJSZ4t43d6uto9/Z1cVf4wg218TXzag38xNwLUu8OoUJxRLiCTCS3LhGRk
1c3RtHtU8QqviK7i2bvSFcAspbkWhwOCTWv+rX6sObUp1gXHW8sihlbkliX2
/vQ6On5Od8y1LtmcEnqxHIrvOsC41FQ85MtasOYKS7mgNBbEVdsp25WFSErT
fhn6e0iPB2h4vCfc0k+bcJ6pWhCM4UvzJTLUaHr0mbTTzSGZZjgd7k1opAZO
KWd779XsITIvouKswDl6+K9IDz9r+H6r8EwOKItYDq2RJk4aNdDLWJ/oJDFU
NcPw3nKKyPJH4jKNwrAhVJ7aTQ+7ozvQvNjdOaWnb8+J4fFhVmir9yMmVBrD
CpmJwnOY7KwCP8Ak6O19fuNTLB2ZyKBeA+mZM66iUglHEU1siVA05xM9Gzwy
Lw5SBWLu3xkG3YwQJhYrfRLBL8l9TOvhFC/b39RLrMJ3zXyPRevXnJpMyFd5
jK7ISt8cTntn0CCSpg8jMxwndvq4mfVUOIt3DaSQlfHafhbPkXq+I2gKoame
Qg9qvR8UAdsoANFyzo9+gVI0RNu8+orOh9Xre5Fv5a/XsfCn4R06yp7ISSLI
Nc6JneGDk7sxZKk/nVBAmCfkrkXDw14WWUZ6Eaw+wELo8LEd7NX8NcE+TMy3
PwJne+9wyuUomuU/2xAs07OF7GYDwcpLU64EP9DExu09kxW8kUdnNxizfSyG
4cHOFUtrnZloxU0bwmNRw9lQxaFs+Ybra+3lfdrEUwNr8CfURyfNU8CsQy/B
THfF6GF33TVXCcOXxYM9QKKYLDrWs7vr8Tkfu+lWuSmpdhPj51GknFXASerB
PQgITp8x/7/3eiBWxfjGk1eEMRQnOmvK2rLxOOrjZVGf/tAHBlojVMku8N8X
EYkZlt1L/pL0CwGCpb+65T2ZtStrCzMSOwISzKL/2uq2slfkrMZNtaGYMvcf
lwT/7DB15Z9yRyD56L/OiGk6Sgt8tU0be59GvP+5zmDvGL+CspaXb7Nl+9nj
9FyWEWi+QFG5fCss36U6v8vExKErO6gdcinKfphPrEyQ9ozRbkYuRYfX6VWN
56qc7BE2s5G0/mHdlsvg6/PKZhI+N1OfgKdc3OSJi4OB3e5mUtdowCIKceJz
39aevxBtHWKbsIJ0Ykx057qLFjtjVpWoKWC6YCMBw/J1xxNIrfis3Qr/9LtU
JcDDRTkgvQbYKJfcNVsDwIk06Z6zVggU0Rs/hlXawXrGGRQ/6MUCw/k6mV46
6flkD1tpHV+HWoVDiSp9bJ+1qgkTzqUhSqzqQv/P7xIFjybfUk3W01k9AwR2
5/f3Jqfa6/3xYeTyovdANd7kgja31ylimYNfKsCU+zwesVIxu2AdFRgBvOba
cqvVZAcyPSrs2RiJcS8z75utYvcjchLoSTmOBLr3sSEvX450b4dFMf6E2Zjj
mf113Rvfj0Jxuqhfr2HUWR/aOjKj/S7sw3Z8W7CwLvkd62OMKu3Y5ASmpORP
+93ql0t2feYMIZbPVvpoUjs4FDnCQd9KAC21vBIiob0TmGFW/ipB2CN7KQoy
9+L4/5T57MgqbosVkEjnJ6rEDxvBNkYTcKgOU/xJNBdnJ3AhVQOO9Pjcm20x
dU171t7bb9qzRV/aLnybx6kfiABYXHGWFwVa46L1rHSnYB1O1ZxLL94xOUCN
qWKWPmibTQAWfIiXzfi42XOUI4M/6VhXSCSjySXLCBm90SvZGj+5uPZTZcVo
d4+M2YF4OYX6n9K1p8mw6Rud/qCKL1/8IFNHuIitx+hMbAMKcEQlL3gOiOQO
tagEl7HYuwI5lo38jVuCIPFGvF8JNbLlKvuPQlCNC6KMUUSkCsrp54UvOvk/
xj2oSO+/nhauJkWDmXpDjY1ximVIMNLbImT//LvnMi4ojssfVTlAO8QWKF8r
cVqgFn+CG5lbwlHI/AytNnHGqk+vhJn1kRqMYsx29S0EhX54h3mtpmwhK+Yu
icASHU2jFOpIPyuzinLTVo3b279OH19mQ7Ef3BXZzrzXfY/x48Jsua4neqFE
3RVvjKfEj05omxJk0Bw515GfoWCkzC1PYevFEKbPHI1wsPfes+uYTwGBlRmh
FMYYwGTH0qW/KX7HdRAJRdbKVfm1mbbHcsVXPQLJtx8Q4SBF3YOO51snX/7P
WOMUd1BYZSPgQIxLjTE2bUxN+710N7iK6Py5VXs9jOTNqCst72RjI9akeWEq
kQDltIrhGVf+F1aYDrhFNUSxkNKGYno3M9/hzeJDLfstOs2iKS5YwtY7EzjC
fTL7h09G4p+wO3LNAw1//vqOR4OMeudEZidUpM8z8fOtTyKp0xr97BF40C/0
GBR0b9gcy/xeCbFF5rJ2sIDPaSFuE0npu04RnNmZTcDamc6hlTeEvtoa5axh
ZLlm7Ur3cDOYK2tc/XWhwcfeOq8JbPaFAmKcsRXDdSi/XyZsX7+Lia2QqPGZ
px9Wn5m/u1o061TIOSu4k+0P0NEHfTI3Rnr+Nku50h4SOEvT9JsVoVzegL59
XgzwgnmaCbNFVdSAhDkMW+YTlbqla3YXa3/1xDvq4y8qe3v1aEWQuXiXLVCc
rkAc1Dw8t6RHtpooBgi7hrFlr57IN6NVhPnUXUopJwm9SJCpsyoI2wJcosBM
l/vPvaD3NdaQp++qUTNPYihXPf34DvUZWrowAgAJ0ykt9y5j3bDWyHpAcjZi
mM9IkdKbxmXhNF9J4PzVEiXmSJgBtlFzKO9Xvwl//Ut7Xo4ie4Jg4XWBJPAi
Fk2vxnaFn7WvGoaBE2hoiiMmlRfrLKKVZzLqWWJpMmfr8Zm/U2IJzjrwLIBI
V5eVAXe/mC3l/e1BO91r/lzEMPuaQ2MYTBJlo97BEwxryBnmItL1FsltV9W+
WXt+VDCSFwd9YD9NR5JAMYUMKQNa43KIT/CjoyWd9APW6pTr/9VP+rBdPg/y
+EDrk+UlBqhB/jMG0PSHnMPhl6FRYD2oZcVrqjEgwpMiQTalAmySejWC4qY5
nIQNCkUc5R2ZYIy+tGfDS19+UnKmANZleCpTzC4uN9tKaY2JbfwlRvG13TCY
46AauLDhcEV+4E+pTOga/vRAYwu79+VE5jlPHHBevchucGl1z+Li4CSFD40N
sg748O42wvSyzJtXNnKA091J8Um+K7jwYZ+itVtPZ2EIeOqZDXNy5sdqvAHr
M9qLxZT1j3UKacs/fUlGHdqC+H8dWew2QxjW7brXrDLGRuGZLlo3IrZ5m9bZ
r/fId6CKM9QwQrQAm+AGXZ2d/LSfiIq0DBM2jjcfIx66StA8H7PEE8xWj1vQ
voW1WrrxnS1tvYk38N9mmk2pDEj1UMIinMCmDIPU4WRhakdl/wz4DECgNsf5
5zdEF6sy8naRozfSnQK/uvadHCSNLUX2jON4lvNlFz1pvqOcpzMym9dOXiRs
0YLsMeuiLv6zy0J8aUBS6+r/qopQlolCRPmR9EQ7X3G9IuLnNRXtp4z0/Zed
2H+KvaSzOSaHOzV321AFWd7dpcP8rztQugXukqb7Gv8Ihx9N/LGhJ/OXzsZw
6YTaGoy2uZ0UTq7mQsmRzSns+dolhU560Zcwi2FONTXru2CvDbiUnw8itSvq
W8cvyLunRmms8b6KP4t7qqHfWz+/PltBGkHXUx5wEwM3dxjPGkEPkjsoUCDe
JOmBhfQRvO8evaTw2wDH9jxaNXXyigZ3OvQwcOMQo8zusCIbxttXk7yYxk78
aCFhhQt+zPfov0adnJ2JwAP42wNyn0S52vOymxQznpn3+3Qqyy6+YM2t7db4
GFObnRw2YMDrgJtmm/IjvgC1I31KhKVYvXeNST5Ok6Zl11mGrP+zx+d9bsmB
7kIET+QJ0587v8qbThyaup3Y/kLhmjIEtLVEqNRZbKfM8bCb4/YYtFDj3VSw
LhVcJQg9Y9a5Qzn31/B5YwtGMHMfwfv6kZGvbhtW3Uws85t/fQIvMqgqHO4f
DH1k+UXiBqFPMdlV7E+TkWvQ67m0QMdf8iOAJ0A9TyzEfNyKfuCK3Hh8vX2J
5I/UBn2d6cDQiHJhMMVxhIXJkPlnT/y7+KJXen7c5kI4ReuITAgB6qj/wDRA
zZ4wEUlnJqhzHJmqkCN5HcFyeNzg/DlZa1qFIbfvneoKDSeNY+EZ+aALs6LI
j0NpR/zaEp5PK5A1fjg6YYyE8g1swiL+YpBOE90b8w6fObHOeWP91Vm1SvQg
1/ctclb29bpXkLIOszpfTsGkro1m+mxefGFMbQwywM2y88LzTCrRiVsbgcw4
UVsxWtdhTd9BALqiuBAMP1qQ8RdOvHyeX80lxjDGg2Zlb8/fesEegN9kocJG
FXM9+LfwjnWHjlw1frAAcICr3z7GX/p9P412QQMSRrlDv2XgQX3Ab2PhWZMd
2WmSLzyo80BeKau1c3TQJfp8EwnqxOosoS8H6lY8AQ0EjXNaVTufQuZv4Hvr
RV9siu7bSLE4h7u0U6hoHhIXksQ2AimFq4l2nMoOT02+7DvW4N7trqMm/xZL
mMLrBxpHguGxjfbPzqBSf+SIhKa2agrkdCzT18/eN9aJ8577GUeIp1k/0FqL
+KktgaI6SlZyQAYgyFCuVE9zKLQiO2/PebuaAoCm9RmvuEvxuaEOuajhEsR6
6fIWXbkF27yu0CxxZgC5PEDyQQr1O/1KSZ3J8rDgB0AbINhtqbpvtDK8uaSU
tYhWCY5vO6G6YHZG2r4VfKmzBYkYC0ftwumzsYDJ9pbiYvx47yhYzcfoBsAS
c3UPTcp1YfxSQrH5C1nEOvG2B8ZBlFTqUWUYHPQ04byWhFDhQ8STJEfKLjz3
43CmuefhbTP+wQ/R6DF/T0U+WJHcNhBbDKwiiEPVT6+EkkmqZWsygFMuIoEP
ybLTTnYGTop+xb7ipeeNuiXsuKLj8mrk/97yeUF2823IZT2+bz8C3erdImMR
ft10p2+QCj0ffBVVO8dXrJl5aLQq+bhyF9HdsFAFmykn5A2wH4yrgvhLFGVw
+pTnbgkk3FW2ULndiph56zbWKponH51KRCv4hFhukD+a5pokddg2eBy7SeIJ
ZWLb7l5hc7Z0JmD3WHSFYdiibjoGHD5Mm6ts2s+ACgXhtuCxIHEjuVKNukEY
tuTyRGPwlqQW7v97salD5uqQfZwrhWuTGeL368qo5uEYFgktX4THJKo+YdK/
NOCOwZrS4Qq7OKyBy2d8Ao00KarKAnt9WCCDCG1KcnON8Ba2u7HCedpVQ3tl
oG1U6WUuSmzshjeCcFenKraMFEoPG+i4NL4kP/HJXxbwd/q0qUhGZRa0MmPT
8CU2sw7ebPmLnvSZQFujzfNL2+QVhv/8dX4rSPeN2gcmA8XzQun9c3bYdF6P
b0JcOF1RWFezM4800NTxS5O/eh71JntpPCXOPG/Z9Gjc8woy2J4EE/ZIxIWN
0R35GfVKkZ/1UlRUz7a+7IOj8UDzRjZVWo2fAfHyAx94xPddgSL6HwdTvgB9
QYDG3JoAG0are1XOPG/90PL73Z4rhRR7x1hchuK67LY6+kWG2hMRB5bvQepm
Xmk3WzZ/BzW69IA+X7GraavTdy0Oq3sFkfJUCHpl0CfwadAAkW+wU/btAHic
R+i7rf419QTRPlmJYMpb7qgtliFZ78qqCgcFutBFxwatYN0iizuJOhhIEg6s
Wsr7jXAQmsZv69fdgZ/BSBo26eZQhOYSaxJZoBq/kw7XwCS0WdoWSkxuXs5M
2+adg5eDYyAJ/gCao1L/kfykvtVpndorX8kphLVxya+HCCLLtVqCWOEHyxUU
v6MIbqdQzzz1VKxiNCwjjlWw7yK/VkZMCpEZLAEctWUfCNlo91nfIMx+q18p
3WrEPQU5t0QLKdIgPuMXcu51/yOYZG2tTwD6ZqCm3e/nQVXw8cA1jJIdvhEY
obsTF66PwmalrCgNHTMcqKgvbY66Hw595VEAMWs+Tz31kHNeKIO5ZkQSaVha
3RTbR1dMxJB66UT5EHAKG9uvjDMEf0awthfEa5TNvUpNi1rQLvf2Sl51DnbO
WcK1OtMtU5ersaCM/Z67gd680Bovdea3j3VqvDwX8bocEszXSx45H0X9Qo5x
Vl6ZIhVY+BnLymRmQlD9y+Pnfd2mdRmGuMSYJg7tftRo1KDVfWhze+K0ffjJ
J4p5REtfbTU9iwmOqccIwSZ8Dec7ilUq2QRsrPM5US2Xn+fwiD5XQT0++lzn
XSh8TdZvJYGjAyxgPnejMohRrGg0P1k/93miWb88jDvfT1+9hculnF5aK42r
bMg8qq5ReJdekpWnMopIq72FNxzQ7fPJ1xBoxZAXzceCBapHhHKTWuTAEIBz
W2QrhHGNB60zKCOVGtsMV1LbnqZMbrwzGR72R8fISzbZJgSDGOSMa+tUd34u
M5g2hPfMkzhilNR2GEkKrjALhe/S1E4l6Mv+nz2noXysUt9EFhyBEE4F+3VE
3Vq/9rLtuGoscxW9EpDkORsWDoRdgN8Od9+yeP9ZYmsSVYXXWUDdNky01sWy
eYIs0ZWJwz+lxqboO8ghVoJ7OTO5OGSt3u/Rdd6p89JPaza1+lL/PGfd1GdK
YNUdycL43MBI4CumSZjl7Ug5XkT3gZLAMYIkSuS54q15WfXLpyycwpUQIqvZ
XEzRRgPAGY1BIOeLj1tbuDns9WvqlwSBvHD1Iy9eNG8dApH/MZgFe77oWEuN
AaOJL01FqjnMyMOdVcXlyZj2QEHRvuYUMhLLhDnmMfbhs7l+kSB/bW9q+0KJ
edsizZ3eGZrtS0flXhvckaNTRl5x/WOt0bbDyAiC95caBCbDnwLAofiR8qXQ
0saJSl1KDosjWk7FhC5+dJ/IBwt01HgVlbf+xg1KNuVLoXYkkqpSgpUaoSSA
sE0xswiyTxajiu07JK9gV07yew+2OltQyJgqQIuF1XcOj5aH4G9noI20K/Bm
v+PAd9DGAJ+uS4jIB0N7ty3ZqftUNJ+4HHn2yFP8daC7hXZ6ezTlYWYAwDnD
IxjptZC1m5/wTIiKzsn8oTicTyXCIK3wjNxuNaw9HHk5OO15wcqwkBnTiy+c
RHp8+7XxudityG4U5q7/6qcuA3mcUFlUoQw809+GUnsLyjoQUqLKqPN+Hx+E
IVdRvy8eUOcCzzDs533JNaHVeu7ceDoBD8NJHsgj2kxUhtmIeyNaQHcEymrJ
oSt9ZTKICFpVeOvXN1y+zcCod6tucfVqZTUwlhOkFnr4JAwoqXAew5dL80jV
sMOpu80ycHJh/gh+NVv9+szCdxrpnrolzYiaiYBjz37rn2XiFcKPjC2LNlzg
PoYfZevlQsKZBGVrbG/vEo/KGFwSE3z1Axpt+n/+j7v7/iNhoZ4A/3O7d9Xh
n1hEX7yX8xzBEKglpbAtXseqhYw+y7z8Qep1v1dhUboUoz1n+3inB/UUlrax
ZmzasBR/TkP6Me2TM91yIeFF6jWqJVE+n4FYUhXQvav7afC9XF0oyq53NfbN
RZ+B19Tp71twD7mhcaQrUWRogO54iIvyD5mv4QZjhoXwvwEetnhzn1aTXxXZ
LHYNTRJMFubZUnN9Xh4ajUPV9Rbn2CKobMjwhU1AYCGr6v/QQPD6IXpfoS3h
51ribB8EpWBwnedYj+HdDxuXcNMgwxLtcXbMluAiRpicd5dT+hLqZzi+fnqD
QN2vfKOLunnOzx678RPxFOiAvW/byTNgryNnTSQIh12YsQqVh8CxCsunZoc8
ccO3goQzSRNNrQU0NgNHSoFjYE5UOxrke/198I8rQgrpwIk7mtebqTs6l28/
q5NeeMCqJvHeGXVPf+i62vwSk6LBEPJ8dSMs3D++yV2Aiwwn66b9QaFcYdSy
xq6taoSxNrE7z8ni0YXap6WL979uR6PuL0VB7/O9gUDtRKU088gXFuwk1xtw
OxV4TVC2aC2U9IWUoFKEPSTCvDTBuBsq40v0c1x1J8/jVM2pjehh0xgi4Rl9
N59Zc3QzT5FT3cVQ0n9r+k79tA5aDLa/BqNZA7tjy20sDdN1bhDn6Mio395s
2pCT/1ToUMh2mo1XAjIl/SVcGuSI3UtRTjCiO53WX0//fIe/KgQasLIqBSRJ
OtZkXQAfIQ5gvOkuq06Chc080fZ15W0N+R3GpibPEmiAtoO9qdN+yXQbQ8de
DUqMbSkqE71lsMT6/MP21W70ouci6PXqifgQwhqhGERd4xNr71hImBlkH/gl
G7BljNIXzaz3HqwoNSofNxgHZFp1PISuJgVhLwsEQP/r/6N5HndzHFOQTrWE
2Gr4hWVV+ZurrIF1VGMCPcij1jH1fsrlFm9rq0IhTXW/TeeFgRYd4AiSUZ4Z
R5W87/obiYMMzIneZkDsVmHyMTr59iHLAE3YWUfAn0PV7uUQR4QnweS00ZQb
B7dja6uPAXpCBxmK3uEQg+JMonribuzZGyg5FJ25/GcnYSTEFLuc00VrwUb6
ZKYCMvc7hnVQn+9Uuej9lE11HwCndvFu0BByY5oL6tFMLPfHIV9nYtjjEa9P
RiP1ivUw+C8Yne2w9PMO1rDpehOFEPUXcSD3//tCA3PIgmBqFq8xYCSMfXnw
ixegrZ5QV3l2OQW1E3ZxA4i4B/DZSMmoMgmKYZzRqSkVrXKw4ERwdKoUv1Bw
sO25fsUryQ20yyh6BvO8P6s/wQsirGbc4hVJdCYHNMvvYwjsBvEePOC4zFzO
d42Zu25lMaIA18x5Qbl24bkUlHXMGflRiSADh4L9UwQbMQ0Lqqb5M4IWdXJG
8M+NmLKJXPl+2j1ITdC8iQTcsnDFsuimKFJHD1xTwaEMU24WzASiByJIToSB
ctOO3rk0JMwl4mQuQg7yiF1lb8DPBjZPjjocjBtG5QYv09DACoFuTdIuukwo
H/LQymoeTA24TQt/aPtjkwDYtZ++iRkVQK1O9IVgxx+tBdBRP97IrvAwZGBs
2paG+JWsESfKNEy/3xdm1rWVMedY0t6dPxl7SswhHazmkdG2sClQLtUpHYOB
pd9TLC70+n/y331bucue6FNRiMvu7gtcwkbYNBmaSkxYdAhdOUoFGOhFhsvH
Y1UAqPgPc7JdPtCS5kKiriCGd/CsvNX9h+JT1tXEbFvNWxGsrC+MDPeSa9oR
tUTo7FRHG5+MKdl+v3KVi5WLtqrNSzpMECrl66Vs/FaAM7EONNiHha8wBpyj
Ndtu3MIlF+plgT0fwi8DkPS2DzCIzHBj3w8Q5b327DXBolGeL7krxZ5I7oZd
LCr0nDOtv5xCyARf38Fip45XA7xO84+zdLn8qGxlntxovT/c/75FXWLIJ9aD
pjD2B383dNC9yZIbajd0HNIgNok0+1nTxkaCAgs3K/w/+P8d5zJe4eYluToX
RmM7omNGM7n3MTrgCg5dsgM8f1IbXcbgmxl9yqmDHsD4lRccMUdQ4dBgF05l
Pz6/8OkHKnbTH6NWY4rOuCYjeqffwApLAvIaVjyGk8VSdm+zFr9vSYUyz5gL
xgOObGt28v/qqAqCv7Ay4nCj42xqRKgBl9JIi+HHVxYZg/jfDpvycOrl+Tpt
uKokxBJOAJxigagomn+5Xd8NMtNAj3kVJyAEELJSin3wGToRrDaQ/YNMkSYC
QlQXENohMc2HDRYUOvjk+BdbfdXf3xIHv4m5hxRjkY6RLB/6shkp0lZoahCX
6EvGZvmKZmCioZki4yLDusgTVzUk1a5N7DTFBf0c+8po2ZDfGMPpviZHFAtU
LnkC50ZdFduPkdpcJCDglRctAGRagaOq+xe+w89TfenRupQfHlBXZHKsk0Kq
r2yMlP0DkB5LQn6XZHFkeOyjQSdHl995Sv148zgfBF+mEikKmB+QgGuaV4Kz
t7k7pOJxVaOcTJcmCA99e2ZVlNeZzW9dCttYzXPzPx7GT0ULtbSvzbW6s8BD
XauIMuneYShkGMFNeJpj3LvKYg2aKF7MkwSpjpasoEERGTblgyL3tCNKTcpZ
7iofT74zn2BqmS8O/McGybM0f/7ahdBy+5ZvI6PDUOPyOW3vci7pPYU8jVnW
j6dNojm6YyEvVp/fQKy9H0C9EblCLVGbY8tzvIxcuAZUhWiY8iYpAk9AqCWW
uMcTE8is3EZMCzuKA3Q04wP5clSmswU4ii4BK9d9W4Yn1zfgvngN/Br/0YNr
F/E39nkvAvkYkMNVe+Mfn8yaIFH04m9H8MxnM+Jbw4OQntcH0wCQqRTW5etf
tz/Gn4S+y0IEL79Bp3h6KT6LfM/rpdf01ZBzTQnkucl05vTcTJ8Dz/dtwrvl
KGNg9fvvqWIQB3oZO0J8SBeIkxIEVj6GhLIVkEyHnvu98k/Hu/ZlRng0Nc1f
YbAJsMgbp/oc67ucAWCx7Pu8QaHDZ0Q4qx66ANRDX7cYH9psb66siZOipybh
egeVtVXt6lw4IU/suwcB8sC9y+lgKITNS0xzX27IZvHgXkN0cuA1IMSWv4Nt
GgpeJ54VK1gT8xczSwEuudi7QSwzAtHsg/KDHsuHhKdupvkdQM82oOpTz/mK
10HR9JJETBu41Ez9EVnzcZofuvgxb530YclRWBcTIfnp6BgJfHGd+FT/XtB9
EU+Al9I2CoQVNEqFjx+NzpPeMIhRBgP9Pug5XDxcdeIQDaQDhBtPcalt0GY7
M4Ujs1IeCIM36u5KDyhmMZtmuGVM+U5gUivNzJgbPKQayYBJUja8G3EaJvCd
Afge4ydasuQnhjsexV5AA4wxodYRzDDt46yVABvuECBZLiWu6a8GM4gclMVz
XNRemSq5GxCIH9UNwQRBBooRDhl2j125i2pX8orkaTxg6I5UB57GNS6qqWKg
9f/wOsC2/rE87G4zkAUCFaPq8q2TTcKEG5Hhng3ixIcwjfW8J4lYI2XfO1OC
0LHr+2/rAqWGzNjFY6Gz3LKIsf2R05l1dl/a6MEA0Oq6rXi3GLXC39yDoovK
KTNgq0IPlDeuXt/VKYehTmetv/t5+IywK0pDgBvg+/qgCw4M9sgc07LaLbFg
zzbR/DsrpFaW3KaA6b5fJB3UUOmIj7F9pWqfA6SJuviWuwven/3+nagshppr
AgXH7mbj5GaSNso1ezaCjImSS49C2bWl+La6kAI2VJ80sYJL7sKQgH87pHqj
tccWYSzXJNMlnigw8tuBTc7HKWUDy/IcYdP1tIjZnrqFQO/qtZLuN/7Nl+/W
rrGLbXRfn8BlJI0SanPqT45WMemma8sCkNKBKD3uelOWEALUSgZULoQWQerX
1MfvE3QJl9/4HME4Ak2204c10HcBvJqNVN4oErDfXDhewjciv/S/CP8McL1x
+qGP7gwf34NRVK4VrXy6532SlCXsG2VK4mDbKbqxbLNsgTaaLmeb6SkhQFW+
uQCpfej5+NvnA1yqc9r1gREVvKr06JD10DZGI3xjAyY3Zonvb5yrHPJ373NE
GCKU0ysnbvwJhtL/XSttFBko7LDdjeZrewv3Cl+kqFmRdbnD8ZwATCnHbgCA
ncOo79oMyoH3uFjhqaPQ7lCL49uyZJ8ZHHDqSySFzXTfZjSTedxhJvRjfDve
SFLZ9K7re5TRFhQIg8bZMWBs5Vvlsd1Xs4ZuuoRxAybViuvMDmofbVIDVVrB
vv5o0UiKiypvwfQSdBnUQxCWjXdsRaoTaIvKHc3DgB9OenobgzqcH4wcgus5
sHHwYPXkcj02hzZt4oB5wnqbSkUjP9O+jWUZUT9GxulQkq+sDyPC3d+DKGQL
0+m33TnSo2F2jBwFefCEackMMUa5gu7c8keUX0cjzGlz9serCI7X4MuWGJLi
R4op1lxG/baGCWxnj0hU7VoMMmxIihsdJCSOchny8n3Z+OnmLVFhnhCE0V0t
kHFYRcrfkAptyvuBITayHiYFgdUXGGIla2qt48S1UYVOR8pk4ev8/bFg9RoB
1PWBVzXLccdI84ZwfFGvs9hwYyS42WVxrG34gYlz0QdlM2g0Gi9sG0JoS/x4
6hIdGhf7TuGriKqhZFxzmpPtxsCn3cN9kZu2pwdjR9aLtH8WTrtQ609mTDC9
eovF6J3U1zH9YCCES3h1d/FJLcdTCVHCneHMp53SHsDCSH0p8Ir861H36O0H
2trlPOOnytKvBKE0ftF3pvJmMvOKZBEbaCM5IljFKaM45lZ2Wn1PnHmjHYmN
Ksc060CPqZL+8dR0LwslsPuuNQ58o+vnvuenT50NYJ3nxLid80LuEkp7JVYL
YrkqiT/A9DPbEHJMNdPZNK0A33VpuYG6RJpJOtjQSSkbOW7Ca20C0lXK1tU8
MwDsTgdUbHzd54O29Mqd/e0efsnVRYGYU+PFgKSWy2GTulhS94RyKFyxip+q
MeWe8THeH4pjqEXPF11n/z0iJmZZoTYJQ1IRS0nYcp5g7bK92JTwtVRTHzrZ
OpHLiJTBX/uWfVTHkqrMaV0JHFr12goRa/50lxQwGs4aiyAIkAsDzK36aGAl
llBNcjGi+u2q1iGXLYSd1iY/PG8lNSmN0oqOzkECnXpB9ZdswQ7+EWhFkwQJ
1pfUb+HFrgMmd/GtmwkiMQ7xwHazobmf7JpBqbx6LZLBI01wIHGoGwEQVTq7
6YyOTP/rVsDxe1r2qEoL86vqMcvql8PUpxuMxPb18WqKk5Z+cL/goU1olukf
UqlIovdH27RCrAuMH1nkr40fJuiyP2C4lrlCZ94veL0GPopDZuP39crYS0UZ
Wsc1My6S3VUxxDURI/krHnOxhKbZLKuD4hfKCE5i2hL4y5Tc1PqSLt8qH6Wn
koFqPgUQSTi/BEtlCNzjkyCPedkdl60XLMp7gZH5+G1jDPQhUBccSFnD7LeB
ilrs0ahRIPQdwqvbJ5WqNgTwf2yskmCRFumxqjBn45637yWwKN9hnHA3Pji7
NjkEgP4ioPI+MySlA180BLSbUorcA2VKVOttRWDeufSgKYpOeadUmPSp5kqf
Ev89jS/eAof/P9sL8DTggdI52cpIsjSk5EkYwvCwUvpnjOP6TXX5I0Xg0OJL
35JauSssKSBhqkAmujSIYT5c5CsEBHcfaNZA+6zAnJ2R00HTPItkLhf50tK/
FgQltrwTyjDltLZMxhkAw/wIGptEf3n3NH8pteWutmmERYuKGwaNo1OI4YY0
NgbEFjtReS5h9WtvaKdzR/4yFe0D5UEG2/fnzUaUE+mN4FwhHdlOTEgCFoqi
8lotJUPu53y/kWJlU7doH8z2IsnlVStDJQxXYf+Y/6f1WPc+OX8/x6l1mkal
aATP60HcRqNC8ThpmWEuUA05g5DI/1n9uyTc3GSSQZTpx6MjfHO0v28cOk1T
xKlYEnACbxasTA6TAh4it5pOhUmdn21eL/g5iB5N1Nb5LloQuFae+0Kuh0N3
pRMC4GmcqMygs9IcGOd9Hy1oxtot3RhGBYGqn8ccsLLFL+WjBMZjx4tcM0Z3
V58Xg3/tsPh6WNAcXcyzA138d1di0KQJPP7LsbYplOAljfHiipuMz1GFRBrv
5IC/OPgu1ywasOARY/58Hvk/KxPW56FAB/2pIwPuRwVALhDOGnrrl8LwfxFb
2BHPlkOo4DlAhXZKJv9xxiuIKMThA3aCSZj8FAnAnkG5vybffO2Bp6f7DyFg
egHNoZ6j85xQJsV6qclTLrlFYEQz07AwnkESZMqbizWSo3Wf8vQkZ+xdglG0
az+6NbYPfpoCPHpWtiVmh5jUOmI42lMG3OwoHqsKag51KFNCPmpZ0wvtRNLN
jZKBULOVjj10qFavLrXis8Te6qdS2VZkzCUoB3StlH8PGTN0aufgxFNh4q5j
hmsc9JLhg+iZBUfSPLt/tMG57L9DCR25P6d12Zu2lSD8NFu0WR/cjLmagpQG
PqV4WRjPmu0OJEvv9PIhl8F/k02huroj2QOJ7gnzbqmFsYoF5nszCiYXFIAd
tfSemQJZ1F2V1eijg1PjR99ZcRcPSgTQn94adnroV2enavoO49faXYWoCMfo
J9qg6nLjSzwtGDbGT4msdwqryzHt0IYJXk8bIivVgUg3M7Hor8dzhB6+ELmN
FNMZ2kIgW/FoqNKo0w4xtKAi+oghP2Wbu6SuXopYIwCtfIogrBDHwW8EtVmS
P63vFo2nRuXU7nsAsbpKGdQz9Rbecp7Ot/MyCm27CgpI9DYNwvZ9eNq30wMx
p8QsBNFTHpPf1E9G0PVtfIhT2S1ERQ/AcY5yUB05yOExFGkycT9RZQZndBUs
CKNtMtRE1ShreSaJnkIYkuHfDsW1B6sn6KQApfT+bGyqPkivJ7HL3VTmynjy
xjgluh1U6XXCmHsWBp5iqWR8wo5I1cFhxccvmfgP7/Z6piTsxqkhHgqZ8s0O
AD5+BDM+vHcdFNP8E16MxTbQMwCcVwwCtVeYx1GCjYCBjmjf7q/oF/Hpzhb9
QgbJpqWlBYR80E1pwBCgSscyQYnblbyzWcq37chHsQSgs54oH3B4TVdTgazN
iomlq1lQ8+Z9IJmoaprV/H1q6/iR10tbl2LSUzVH4HZSpKSpVCRtWtUBg4ZK
nZ9XXK4dJTTTylxEHsjeBnvnq2hxJNPmZ/QmFVU8csWKVbk9a+mLrWBohSQn
3iYS2XdAYF8MOTOPTfvq6e9176pRGN8r3oIocb7vmT6M3LaHkAap5Zd/AOPV
++e2D8KPWC10GNz2aLIzWRjRZNm60LeAtmdPZi6FM+O8vFAi7bFQRlKDR/KI
TnUmRA1Ect3tH3jXnEKYuFWcOQ1FKE4jeFAfFAHX3RK1fBos2Ct6jbmhlFBd
+zjwoE9+7NvldCR+vBWX8YdVzEW2IRfGHMXGhRheZT2HMRH7/vQHaM8NeHUl
x8cozGGOj5qDDQUhO0SJbgFs31V848KpIorzDfk/gmYu52yZpFp27R8k68u/
e01AlSCdvw0U+AZhZvr1h0z6CwcDaMnjuDjnCosZ4gC0qIMF6jJUsF2z1JXq
Y9GWGSLngMkTt81tk3Kl4oc4oqcP74N4M0udbesyL0ilcPf0pZyBq9lp/tQ+
h9KPAuYNpB5aIP9Y1yzheDbkH5T8xREeai3SYC3EI/JjzCW6CCDvw/Tm9fzh
/Kww44gyIbnSU8Pg+L5tZjXq6YHJ2UiZaExtuAkqyWcMV1UaZYkDYS64szTZ
JJRKV6FjyBI7rWqkNR4BzZFv1TXFbCxKySYD8e2DxGB2tBFbHhlkt55AStc0
VPRMmhDkLMiEn62+49QXFi0I9kezh+fN6wBaUgTFuqWoSnBET3d3PMW9tAAN
koWiL2PbGCmT/zwfh0I+wtC7Kf81CrWOvuRCxn3vjDQxWqV++GZ8+a+X1Ax9
jASKmUchj1BWed8l9zmM5bmFyHu6iXteSQ20PoasIjm0hvMPqEtOidLFGmcz
4/X9C2eQxzBXAhIKjeKYGRjLMfs9tzlBw6jUO/t10ppdPGeHc0mityVrRniu
Om+PsMjoG4aqMvLdmi5adEJZ1S0I8JszmiRHpwco3WA1Kpvnoh0N+DcKBPEO
zAuI5LDjEhh1u5HalAMT+hJ0aLoWzaqNU0nmZvoSM9eIxZcIYnpghQbipY5E
q33cJttljN2/A6TEkpj+BwDNfe+zHSsSg8pJQozVj2g911Z0WhXxGRoP4rnI
syBdxGQdg7Tt9/GlW/tf0JKKEv5k6qbeeNvtSvDEbR4lE22tOXb4sWYMEzC/
DKmfIjIMNt8lQmhRn0/FbPMFO/nRoSnnkGiYu6Y8V857LV72+n4A/3O3l3hc
nQpAjlV2Nc5W2Xr8xI4mfoiq3upYASKf22S/2dh7jva1AnjWJgwldPdH2p5o
GeHsuj6SIOqx5g9AwXFZA7jKUggnD7AENMsltM/JWfGxdonsV19NsPSOtERi
+1VKyqHo+TnGtCcjGPTKzkHBz69MciQSLCPSnCfr/lQZLs9KiDyGenepz8n9
OwvbNRBtVf2A9wWBS7h2nh+49Nlc6VIRtK9Ns86JIQ+MZOmsqIx6cwooC1UP
EDjRDO+7+H5TQlmxHcqhNTiCo7GgOWgMfxAMvF9GRxg4Crh/Pf0nFf9ATqC/
bZGJ7EGE5aOFMJ07Ydm/AhTAniHDDxgCQHQ7DVc54cGubdB0Qyk34wLf1AEb
f4jVbaZsqoFwcnG08mvLgbO2QIquVBwg3IZbQRA5H0P0Z1QP/ayu1dDaGyW0
PujTaUhH6i+3sEKieZRTXOwxgSBU0f5aTXU9WBA0Eoz2M6UjUTrMGuRBaHO+
udbCj2hRx1FyVYDJ8BH4wD7q71h8C6LesjsFLNQ6VXE2et2i1O3buJQNFVDb
IGZE2hZTvUMaJKKKcVPXZq7urA6gIXs+CCGtcORW9FNArlrQG/wnpqaGlCHz
olUWgThvhCbNVD/dduPi28nBURjPPHIhmmlbnFGvhfGX4yGGYZY+TSV7kR0b
7K3YJEy+OOrHyDTgnZ+2YyKGCVokw+i4eTJAR/6QhFVDQCuuTvJ+G/7J+e+/
Ort1h+0zSs72UlFKF/aJaPSw6C4gfzJAjU0bMQDJyPUbVsSniW30wKLo0MQR
K4uebgIIYFAdlp+vt81spUkNqFfKh/nodjsdLt+8ym2412jMGFNxRxEyLPKx
pkiAODpl4XFhy1Lr1e913mzfyEFsA8HvTFFHD2SxN9/J4GoWELfwsVdoGLTy
LJN/UOu2UwvDoiFwMvW/ftkGnEkBed2yjGp4r76iLUT5Bzj6KBpfKkO0e7jK
JAziPOcvC+Htw06wJXUj+tlN7WypIK85qYYEcDlIYQ+PAWmVkJDzGR3dqvQR
JPIxDGpE3aZ21GsostTr8XFeWdE+vRx2ixnGMQ00cqZwGlRZo1zUoW7woMjJ
/mAGhCZwitJjy6sqITFLrDH1wZWca5NIIOTgq/p+cf1BK+6xMdJZCNR9KDrO
ySTivEuW//TZOaQFwwUopYTUCB/PJ+ERG6iNhWDK7iHI3VPAzjGEIPDgs6aA
jIzWAIC+FNQiHg2X48ozz2l6dnqW40prwe6pCJq+m4ENChj8geh6WMEMSP1C
NZf/+/dpnbhtiMmBHhTaGyjxy5dBCTp7mFGNihQXYSgWcrWb1RM4j+dHqzDa
C1JTQEFul6Ua8FXZecBIZlBIYKcRMIKaj2p9ZMf0su40W6J3+hGceTWmeSBP
kID6Df7cHYnIpK772x1Lki3HRwoVeg5yh9dQ4dh5Tb6hlToAcbCzBtWtT4b1
PPTQIAnXmeQvX4XZELHQI7xmvq0ndhyeJFplNHwOHs0JX3g3yxFtfY49RtD/
hyoO9kYa5VEOffLX6a4apWurdycFMJYtHSFAK6tFGcM3mLoAy0CrnfxYRRCX
KhQ90SVNwXjzgaVh4UZ9Vsv8moXoqAAHiSL3JJ37FHi+e6MldzpSPmpnEAcW
WuNznQ67reuapU56fmKunaJzzOc2JCmU6GHUAVl4QRb7SNAuw3sBGnYiAhUr
l7PtMziIXVUJzZBU9EalnvurTBMnyU1jI57PXSbihHCVnIbq7WEN/gCDwhvo
dyfjIg+VC9xF00n1gvpHHUibXAJeGnZXv744ctVDyp4lEP4FSkC1Je+51C3j
Vsit4/+jhbmvTIElAD2eS9V7Obi1GtdZ7Okq+EaeDlyUktqJuqXeTCzJDN0p
qJLqHrrIB7oHTek+i9q3sWYBRMtcIJy9BwlUwQGgMf1sYrO93muj8NYRHNrV
eXNerBI5lPJjalwEwFTtz8CdLD59dVL2fJ6yiSPGSf95sLrylW8uH40boqdF
VphPm1lpisZcPWQesWhPQ2qDTmKN+5Wa7l1VaC8IH8dJboF2aQQEZVziHfSU
RWwlCuYvk3BQ2ahTFKOlbBfBXHWTNfgSBTOE+Nfpw+GvrFu3yHQelciyblSy
kHfAAywhjT6yI7Rf/BG6UPJm+NX8n3Z5oBKMWTwenMg2mzOK54u0DWfoXzcZ
PnA/TbJwkkM/YqHs6YIDrlJl5SINdbfZr3fF3XLovdPddsr5F4s9bUvjDqfq
HT98rLmTXwEg7lQIxopsudsqU+5Wd06K/zRpMnjFH8IhrkogWUQILxn/vDq7
DCbICqOdu8fymP/gQWz7m9mcBKJ8ALrvWcAU2jWMlzknkVG1R3ZljtFBc6MO
49XJjNVBtfSaGRFtfOqBiv9S2O2Qy1vgyL+z8ht+T+lxeRXLAqgsxCxVJb0i
E0sKEztrcfVLewm6dVDB0EDZEwd2wbxCd5Qs7RyGyCuRFXEQPS72aalW24g5
6FI3xA7lNapGhBCrsuGYwEPQKIh/NdgbhvBrTLSGc5CbNryB+wIt2iIGAHrL
szT35kdmfv6rxAYpa+H4hhyR3eRcR8G7Dr/XoFc/BbiVRKIwiUP04WKKabWJ
PtyDNAMNaRW93VWorxYZIKqfquUMo7nfwx5Z8AhdT54qRkEaa4+PXSnowOrG
f0z/zGDZPwE+BXxP9+gzeJjy4WciINS2Qze+wLMY4METPD01hOYv8mLGRj6V
9Se48Ah8na8oz7lrbFjCVDwg92inC8K7CMLNlhBh7aEGLiFqzYuU8Ix51ffT
rh0jzqVCkCEVnS8gdW3vkQf3cf+6F1NSjGyXRI8UZXxuNBBz0UTHDsjElaSb
A66cHAkRbB0jnlFhi3OcQuDgWpDh17hVHx6sZPWEFJp3KlLRJhSCEyM3jp4r
AW+ejSFEbdv9jpdDIpIl9NbVeI8tW0pYJ5iBUztnKlf5y794Iit3UUZKjLKy
z4XKxupIuO36dg+qCfwmbam7ruU0lGOdQfgOYb6daDJBmmFcp14idIcBngkI
x0NjRQFBIx6eqG0M0GlvT/lbq6F83Ug/AgF8QN1684v7PdMdB8g0XlyCFwdC
DB04FmQfyC6nE2eB1DP6dUPD59GjSl08DAced/VPZAc06ZJhLGygNGnOJ2xK
vMfzHsmMmfZuEOQxmB5aLfkmszSEH0lLIAXFeUp23NnO3JYOXaUDj3Z5LRNs
RnSrygrenxtLcmYwfJMyflV5L3Lg6LS8DgkpqF7cwIM0SmiO74kQlWeptmmW
lxMZdVnQT0KNMa2NjSQtfyFi2F6TZJOyDAKxH5DSNjGESBge4vt+ShsPJfhh
gDfJf7q7G4A15d3NSVLmcJQgqvsWLjlZGfDoLKlIIZ5Hc1ydb93+kGh68g7E
hkyJnGHcuSjs5TYBHpFYQcsFh9+4zQdxzehg+KLGp/Sxh24+fojxARmKhyGK
B7TJbxjZ8hu23WZxYgk3FIKcMx4f4+EnD0htpZ2Dugqiczy7OTQnx5PPgju+
gKMsZe3Upp98hzRZG8O8gy6XafKtI5P+/Nh09un48JOmbz2BGN0xOb2EnXy0
RSegk8h3f93vFWYbB28Tf5P6VsPCdrNbmFO7fU4XQnZNOXqaF3KazkQN0VPQ
uag1ejY7O0So2g8MPsdUG9zNrsOqExkvyo5OuN0fg3nF6qQq8Iywxns4phVz
nG90+HVpzfrv5YYofhSk3PkZqflCakzKssNChAehJkE8HOVJyJWP2SudLbOq
vSqKeX7RAhfdzu4en6W20Wk0e1JE09k1rTVL55UW6VMpMFaavy0jdf+frH2k
7IHJZSX3f0DTtbGrgdmdEatM9wYvslXDLJp66UgfuCOaFcIouRUfL9sisDHj
nvxNYUyAgmpTZ9k2XtdjDNI5Ez5ih4ELKdEHjhYMvj6Any8p6sX7CXc9ZT5G
/Aknsq9CbdSojdqhJP7GKMjUDtXWJRnQGiI+MDpoz53BCP348XfTj2wUtQlF
1wv96CPwrgDa6fayO6EFadKcCrAbH2v9KWR18VGq5WkY1HGlDPBgo4lusLgX
k+vMfE1iO0YqJAYFp7OriSp/oYBjyluYTMO+xbaQpFOf/qFUCH2HVfcJGYr7
0bT7Qpl7NXa2jOvkQUJ3Hcmf+DkpMJpX5e8SYgQY+oHUAekB/q7HAo1s4/6/
mVPTDB6tih5S7KKDh7i0Pon8km0YduQGkVHe8UN0pN7FlxY5142wqaXvwuSZ
ZdH6CWJrD7+82BtTbg7djOuuybYm6gEKyb8dIf/+SskAQyyrh3GihQ1pjMHn
eUE7n8hhv/cctRNuEtaB/j0yclX5zlAaYHKzeyMxRCfmVptzbV0hZ8TfC1QD
o3mcGvQDBfI+h03sMyTTGh4zLAMlZL/YCxxxwn0XO6i96yd7ogTjD7Po1OBf
90NTICnqNPczqVY2/i7WLBg4k4WEUKSwnFO2MJ98MH6rcbZDiqxYsg6RdTwQ
qSqj9B47z8HhXJ5+hZnBwWQT/6YNLpFBY11xUAEzZVmXLWlvR433Q7kd1g1i
ern328r41FCR6kDYeqRMKSy0vWf2svExy8RjXS4N0zYwJuKBpLnZrGF1//Xr
2te2t8uNs30Vm+MqvCFmyv9wPPW5BBdoGiG4UuOPjN3KQGIi+IMoE01rm2MF
8L/MaH96MOFtVFGOCJPM8rqpawxyURyPo6/yxQ1cxDMiCcDYMUgK4wrhPpBb
K6u0YamNufPQww08ICKKxWenlCB5xiFw9Mat7IYxuYnBwNMAZ2DpnWiqgI+q
WFJuAHd9ZOFNsCvSkSXQXrm+hcT6D49IcFh+mIghqVid6qbBt1dyEr/MF28Y
JkF6aC1JImXfEDl4aQXYOAvAtrwjzqwactpuMPSKrsH0UMrc9+jLcuvnE3JU
QIRR2aY5PsPdzhZu0vIEEMHBET/f+xjusJ2cXZbJKQ7/1G1a5N53+UWuPEXw
DGp/EMYzHf/Q1SokvGGuo1ekQrO2YXgVxgn99rrFB9S+7m7hmFEmNq4JNC5q
KeHHzg6wvcCtf5KDwYF8UhKbjwuM2RGQkktzEgeF3rZRV5CnMGe7O8BzJKJo
tnryzS3STFFGAT5jQrzKoGsYo3XsUhYszzOV1abksaYcSK3Kj8goeL7JouOT
Se4g6rv2N7EVvKepAB0yeSEezSzSP1PWePVRW+Qu1sdIgpLTB8QZ6LWY8dlc
qFVxkedpkV33DBNGDPw2GWH6ho41IFPVzZTYtx2jQUBMO+NnAAsOPydzPPhw
PN9CdjwMFxc+RKDiu+96GfgA1QSx9CUY3YVEP3klJX4UB+O0JK0WBRKI0+Xu
NUXrP2kkcoXbYBlsNVX7CqfE+HnTTTBW51vMH2etm5BcCcfr3iuEWAes3fQt
H7FeRsYHVez6w5ISl4kiUdKwBdB7LkzPpsZIVNuTu1yCcYNToli3Pjhos5HV
g9/hQ+GZprJ9sUF6sumQyib65n8Mx80OddrxvXcPIi930y8ZjoHzB4xZRYRJ
lf/rOoG16ZtcJk66vKPod6kOic4vCwr+SbkK1mzIv4c6mUNodvusuloCcKY7
w0G7KYbPKQClyp/BEe1GCfCvmooL8s2ePIWFvkZg70Yzu17SZRhUcqPgfLMQ
RCHydH+p6IzMXu2mhu3OQ8240VdHbEhmJP1DNT2CLEr1Pdwr+Oi7fiCjfQ0k
VGkeNaJG/N9+bg+mbYxDfaTYBJis9W6DcMSJncPROHosCqdndjl3cakAuEFz
H+Vju3J4pz4DhvwJNjxZFkAesMqZ2RxSprQ1bLdnov1xCL7BU8Kok4uMm9Yg
QLG7BWsoJD4q34wb4CSTJxSe553g9eBFjz1coMHhyzd7i5z9JBS+LEfkcfKE
WdcY5L8MXdTlYRR9+hyg42uKo0NmLGN6qjCKdYS7tRwySdrjG1IFUW8jCYNO
Ot3uJHt8hWuTD/7rem3qG69L9mTsSezn8OoC0OdIXUNG5LV09r6AcKPog8Av
8o/O03MKqXAVHjUx5/yeXCxmayM4DpT3co4SKfwDA6fQiSyTXQRbL41TtiNi
ODXiMJ/zo22k1YZbgR9uBJ7yPfsI7/hssNCWSCxm1BGZchcCveqM4ZhoX6Fi
FIwSMRluVg4or6Cjl+qulhY4c/IluaJrRBGw+9O6hIQK5Xadhosz+4FFwsFs
KjnI9m8kLoXTXicpalSK4YbmJ/Q/xrULX2PNFOtWXPmU0qbP/zXtXPsOiFki
DFfVBSKE0u74CDMpnaQX/TT9hoDEi9XW6kJ9joKoNU6r0HhBiA/PFF4PpaKM
siFlrfxeFVbod/3/i2rHrCXaOR5dLRu1NjEmUVfzf+BUlZA4t6H6VcQ4TLvm
J5hnNG7NB4so2Mise9O7Mg+jM7jfTy5LW/YYFljz4PhaObG835S5dT5AhIhT
rBRO6PFmUdAoeFggEs0VCeKm1L4FI5abnnZT+G21M30g21YrAQiOTZhbVShW
+Qp6tmPnWTn1WTlB0XQklKkY7EEQi7Q2yOwIi4U3sCRRAnzkAC5UFY+Bwkm0
hvgxgIrD1OW+XjrPbr2eEjpLFYjDl75rcTqbt96hi1DJwAtWEy+L53scWiov
ucl5RDavOXBSd+UvXozOJJaUDKEK9XeR79kHFsjAbk7d3BOpuEV/eo65nCEx
HGZP+2RphPXrDeVRbH0s/sX9q5wrzMsFSvcNBcdeCKUlpgxg3fXJJHjbqyWL
auFTq4pg9vCSqlNDOPv5VhUVxZagdCAVIwu11VmQ3LVUYxDpYU5uiohMvlIJ
7sMjLyR5yqXo1beJRHUm/i07ZLyIoQk3yUvaVTmV8nKynpE39opTgx9dZ79O
RW7k647dKPkB0uhkd3nh2q2cCd2MINFJsa6rZjONik6VQnyebmBg10xfYvY8
GyFTZ23swwCUK+OE0pjaVxJlCg5XxVVeKYZcnrV/pTc6kANqEAZL/DTdq0Ba
jcS1GkpE8Z/+KwQJKQBEjAbI3XaiYKKTuV6xf0+JFGKVFtGVlzttR3v2G5DO
BKlgDIWUlREtLL14A+i9QPt9IUN5xm9ywjc/4F9g3Lt/EZAuc6chQS9Uu0Q1
tr1e/TnkXTn9mxT3ZzRbK+sQtDyFR4NFb9fpMyzT1r7+0EhCHVq3yjYOb7yn
lQKljXyTDFp2Cf0yAN9iAbGe1l6jHeDzvn4WcTVKAfCJGGfqn4KanMVglEpm
psYfs1WmTxtHoN6R1pP1qq0TwYb5kmYMvpHu01bd8O7E3pRHZ+eLWBtH0JYg
lnmwFzN5YTucfoRjCXl8sxSQKpjeMoXHZGUb+6peElBOrO6LS0SFC9yzQQGN
KSyhND2EJSeHKQpYNwTXveYG1XuDP1FrHLrtBMXyjJ/REY72YYpnlflko6+E
aqDqcvo4RaJNNCjl+nQc1dH6PO+C7n9W4wr7KFImB+kT5aeI5jL8vbE9XdoI
Z7u8AQ4sYLe9KL5CixHzSObtFtUswPoeZlLaja/Qxbkrh0XMHL3yc3/ylr5r
ZwvNnv/OgdS36XMUG77zZ190PTUXTaFBhOzULY3RJuKPqlyqoVoPW4mNyzO5
j991H1jMwaeMHSPc4t7kTmI4xELgUA2A5Z7JCrBgo0AUZVtVQ7I/O6AHrsWf
vaxj/+EkfeQkyRHAjsPHh6rQu1+KLNmCOu1GKeVPw6QULN7lfHoAPlb0kvD9
91H8YOdQUFxW6MY5zl1l2oDr2V+5hMWgjWJvzy7ev54J/cYf3BMi4s8APHqa
ts+uUIXUy9h8XMzKQmO2NK9qYltkUWYR3DJOXBQLLLcIXm3/NyNefN0TP8Aw
Sk2CkHKHrPB5j+QsP1EZ2KKPwLFHF/6pGXDjGckPdcHkac4B7+bzpZeaeBMw
lkcRL/DRrYr+t8Ykx1zHc8dx5btde1/hUrbkpvtCqaNDUgIQOZztTpUyHfOj
wsbA4Udz0JNFbQihSZ/a4MZLnd51RgpCNMnde8cuYE6LHCdST4G5ZpVGAGwt
iPUqD4n3BmYQB3GQ7JVDOqFxeQKFQw7FYuWF9lhpY8T2jX95/+ktsXJyYjYQ
gQnf7FHFBmbwxb1pNdbUum7oTpbkCxmXswu8e3czZ6OQxaTS9e8ATLSrsf8x
+AiGMcPsrTY9GmVp0jgHjvXAG1b7b/6CpQlB+Le+x1j5K5zt1NmGDGYH+9cC
4ZCFUxklHXTuPEWjr5RYeU9u985soDgi3WvRl/XuptjwAqkQt84ruftdso6q
YeyQvd2N8LHeVDG5TxbLEU2BnC/cLUVGQJtqSnMLk9V8VwfaKGmv6bWKqWaF
7rVke+P0jO3f70OzGS/mBoCJl5F9lDalreAVCAlDtGMwpMZ2mHFfMG6qbooK
SXQIdK9f6FXakvGuDzunMyNrmk1nDk1Z/FIaZgwPpgYr6C5QWra6Rrt01qQ0
Me7LiUQMzn7vXLNk9MvfWhhFT8VjSEYJ2PIsiYun3A2KpQCYa3c2yFSBtgmf
JAvzobhomb0CAUpTqPBGvfenCJwdPqZSgcIvz3mKZifQSK/tuNc5YD9WUQ4B
qOjQr+BTqsZ7k1D4rr9q8kqx5TjPpu8uL3SgcPZhP7wSkrrC8kHSOv9gq7te
bPuxIxK4BtcXRMTuB8oa/n/S0y/B9AXpUCLMt0aHzzGezmmMOVbpvE9kQfDH
LkgpovkhBPX04+zCGQZWq7VKpfRXutBZje8GXgEqwlLmedjxETOeMnPOEH9o
jLbMI+ktqWrkc8DhStTmJDguvm4lG8+Z3z0SVkQH3jqUVT2R/JF/2kt5aCj7
4IdeIIolF+OYT2qu4qPWlKbCFkkK0I1eOy5/7HcGZNCngotLXIIpGW8Onbbf
DHMxZ5e/P14zXbjqTqWPc12VglbFNCJKcPw/UYCXN1fUCYgY12ziq5G5kOIO
UpJ/8Ahaid+Fi6erKfjOt3WCcCd3J8xdenv9mgwVmYiuanDLBLABk1qKAa+4
RV3kyy4o+FaMzNARJ/A6fy+OhcLhp0+kq90YJpKYF9O6fkxw1lnHKoNYCyxi
487ukYkkFPLg+Ajp2yWAXrozo4WCJ0fiXj7n24fhkEbhtHYJ3idpAHCJeZE6
FOnH2HmPQYAgzPil2D8iC+zHYhHc+XS0Czu+N/MjI0GMhwk660blGYwSUY6+
NJBVcdMo3CNZ6QtDhXJsU9IfYOlzSF/9dQ2u3f460kotz+v3cnaXwo0VYWBr
o7IKbgukqBxV+XNtJ84SJARP6IJc2UR8DJQYme4acRJ3fm8qfK6JqjtiDHoA
rPPc9zA8gAPVlnidK+8NrOKrO568j5lxZ8YSF6OZ6hArlvQf0E3EXNHjG2rr
vavJSI/rLC1w97GbZoJBEcm8WXYQHkkHVY8AX2+ifD3ZENbiIY+nz5wl+XpZ
8heWf+Peq7y8mgCNsQik8iH6jvvVvz6rP/LF+aqUIP9AYrwHEhyoMhHzUd8j
JTz1F8xAWZLyhNOu1Rl9e4DB0JeNJ317d/L6w5ZX51xk2CwLN6UWULhWtANj
6z75uGiOxI3aMGX9isgeokSDBJeqHOtCyxxQKljNF3N62Rmbx3otSU+JE24a
cwrj9K1UjoqE2bO3exxx8vljZJLxtKlNAZ7Vp+iMVLMbvI67mfYpmTNpY6DA
QINFcGaNTsF6giDLBDeJMm+fmWgiHDlOv6I+iWxTcgVvw+76ml65suqkLDOE
j1IVf9Lfc7Z3THUOiQROFs5+v0ns2L8z+2eZIvhqYomOz/vakPXoqWseBcUk
AG38pdZdGwQ0JDROlvhYhILmxgprDtfvkR8Ak82W8iCq9Kb/eSLCTNjMYLWM
59Xh/eO6uSJ1SbvcDcZ5PlaUdI0VTWQ8al1zMHYgIWvDqyQeRxqLbTdeVCcv
ZXgu0M1x9MygXcXEQWBiGmzhWkXBhMai7kv0P8Y6r5FRHmW0LHpDC2EyNTEa
EX6fLnNrRhrjK/+qPO2gycx4mYj6iglVIPHBjSm9rUlw2ZZZfBov5dNH4okr
j/oiXT4q9qdKNSYBxSR8pHBa5ztCw7tiyPYlrLdh9sNCu7PLu7jczpToIOPb
+TDxWxfjV3XagLXSIVbN0n50yo8CUxRstje1V7W9K712J4z+wTXiwJ5cgN3T
1xKEZvqf3VYnXIxCtODZfb4WkeWecxODis4Gi5HbO4tDY6vdoadnXQlkYOyd
VbXmIsX4A1VLm6o6bWZmfk4lHc3YqIq4hizVmO94rgc3Ss2AtcMePgATbBO+
6wuh/1UzcdAKzuxYEFQwZA/RvxP/jzQNVJDR8pvToHnCe8ZkOIuCZs/ETXAK
39w/nbcpQMOCme5MKHAu90l73VDjQYnzX8E2XOkw8TCvEom4Nb8zYrhdpFUg
9VgMFfZHM+dEvKbjv6XQ/YhI3zuyBXBCKDqHIaNm6Zv0Tgp0aHcRsOHVltH9
9oiB63ZMIEQ5TiRniqUcemlNgWzLVvXw1D8HE6IYcw7gdo4Ms6C0FvY+T+SX
V7OxCqGY9CadNoJuOwlEtTOM4TTweMKOn7Q11ipA0uJd6wdZ4lkdzMmsry5e
+BcFmlOhKlU94NnrC/uOSUwR99PkzNLJofKKXESnc+btmBYkWcnp1j7FhMCH
ZPlxnISVPCT1mvmnSwpEQ+OBA0czv8byRjw8Xn89JONyc1StiYUxaVJWl48u
dQ6JnJ5UYfHnW10Ie2FfnnT8MqIHX5YIhpFvCEKTrP7+Ffirw7b4X6+Rjv00
JWKj+xXjHOhE+ICBwiwNqHnEIl+RZrxqBXHnLhGnBRgihCr6tX+Muz5upRfX
cfTlUWryc+6aM8FMgUs9XkF4ybdLyGsAJLPRx32PbJa71TO7s7+KqcWn6WC+
91lXIKaeo4ZzVqa+aFb+niWUxulRJWeZAdcEczbndWL7VmS8S/gchctI50bA
6jTC71fh8Zq11zbpiMZcDZA8Fygl5dOsK57jz4S/bo4S+wT79SI+dV22O3om
MGlzIZ1xdyrJxh1hz+THj1BmxM8zBUezB2OpqNfon/P1UV5B49ZhXIdAwtrP
zhtbhm8nXiXdrxuBEwI17N9XosfqoXnpC4m02T88xmnyUkIyfwE0F4J7hJjM
06pFj8q71rbCaDJhFXevlakY+7TcEZfjlhx4svZjDvQLhEBaMQhmzAo1CJt4
JvP0HROqTr462MTds8snZZqmgcl+ULVaqdEPxk0WI1+8py4iw9KhKlUeUIcn
FtmpbS1mhVXjM8oPF8zmJw4Aqn8lgei6+D6KfxdclMoR39XZ5JAX2cHQPXiR
L/9V/J/08Dr9VEG3NODC5b8AbdEFb9WUCM/C1y9MNDOlSGveEi0wnmDvmIDF
NZVqMxlhB8Y4hjolROGjDEnfk7kaLIPERXtZ12YgO9Asu1M4L/5cRVEtZCSv
Lj/t6W6gBTTQaLgNFUPcFJcGeO47JJJT2bJrfoqmWPCscDa8noE5odoQMilT
OftOeBxnQLPKKIp4Jc6RwXPQaxNdTaUfoSRyBIZIz0Fyo6M+3nCDdsjQfIcS
ZzK2Z0+Omldz0ppkVC3HlfuiVw6r+qP3K4H4YARsUftwzP37TCdqPWWc7Er/
GvywltdamRkHRrqaVnd6sVjZf1Ac6w+Is+tGr1Or83oVrb2T2xEATkC2QogA
qGgktTOgTjAX7xtq+ksvkuz2OSaSWWj4TRuWoUs0INCp/Yms8yI2SBVwoWYd
ei4c21jJ7z1VscAsTAPUlK+3CYHrbD7Nb4O7SOGQ2XVnI5nqWHfw9iZH1v5v
ay6GzLlzYLoeJ5YiYUUgRKS3rWKpqTfGq7I/zayFTcLIXiTGmTRXqc5dEmK+
Z+LAQCtkk79AuN+h3RSJ8vJ5jU56ErGoU3S1TcBbrW2n76BJswt2NVq4ooK0
J3BBDbP2zNG5PYHyv8prMSzI/FVsway1MA0z6/1uIsBjJXdl0A7eRCIXNX8f
g5EOd6kYHbfYSQqqc7bP9v01z52qgavGimkYuUz21XY1wOA0/TJTv/hegTBc
CMX3Xkk0Tm4Bg9YMu92WxTqCWTYrk9XJpAlDkBWdNBhSHP6Kv0hyeAuOVLqf
Pnhpy+w5HqCJVSyle4691Uj83P2DFga4KQTrYQVFrAq1oTUV1QwxIcXlHfLi
kVBS4OpIpGGWw8r8enwvxcBvc+WTJykUa1VEbAEJ1InIy4TGTp6gJCYr88un
T76IgGi0vU9JOKHJLAvhlJ4dNxHlMj+6l3QRTqM6ZsccztgbErbggCCDvtcD
LvWWRgGo9aNj655AvKZTJ88GaIJWkoyvJ9OamxQBLR6V3S4a4v0nLnqMsEnP
8aJUpQH+C2ZBjY7ahsIUt+t/YWNzoFM3D+7j+XFHvrS3LnQaIa5nkOUJoKGS
4hiGq1dcqJWZQSQJCg3cjQ3hbqY2n7do3HVXC3BRtkxvQMhIPsg+CgClO4M4
NnK3IM1ZluQZ8WMMtfBdgZHQD6tOg9f/tM6vj1O6/bfEYwUwUxs1qvdZ9ZJy
EnBO3YX8/Rkk3NfvkKtbFlsq5D2Fte9BKEoUa+nI0ikrxJLqLfYBzUiYB5VK
VU/TVcXcke+CQGKEG2qVTj+a6H1cMa1m2q/Mbs4bSDK500w9ks55A+aIvVRX
jM4YsvJtHs4nzAZkPqanB1lc4/XVVXUm8gkH+I5z0PEnowGynlG9GZND5HTM
yXS7+EbjpWhaLRVET3juNg0MWoXDdXoNuLzHhGMnJBy4j0FfSsUC3nAIz/VB
aSkzQl49/pkhV67KxCAH6zMnpxJNgeYINgadM4ycCFvUyW3bAYCfALJC6vXs
2BbIavSCRKQ7R+6basoCe0JSjuZmoN4nVy/tpuN+SsN92WzalT2AjHiNYG4K
nFMegDHf1zZ+VeGN8QdIUvyWZuaiTkebRGGZtxqaOt4s2aq7Moi/JTO8bPNf
/bdWN7mRgYU4Yk7AXJajJrGU0PiOWAOiYdfhx8JuL0EDt6+YIkZtNpcpd5Sn
BD3ewdJR8q5UteDo4TS6TOg2otto7LjaMBSAJYFjofLurGCps/eyeyJtaiFt
DzfR24dgrlgfTyDydt6S0H4i/rZodsyDwsZAQnTS0xWwmgGKcss0ZEyJ8lFc
5vRY2V+OH/QMLc5lwzUKa9EVjvfXWqNz4vbpk5DsMo0bBXnqsmuYgtwb7NcK
SnXoE6so1rq1x7uujFBKr5lDw2Z4A6bqBVsi8Ayrf51oKzRkY/rY031yT2Z/
Kd+A+vf2Wvm+6y3MhXNX6B3MtORv0c2Ql6dLLLD3I/cpjmgtw4DaTHrz+azR
TZqiC80Snbx3sXRGuZtCJHS0wIc5olEyOZVwCMHwWUPqI5Ltu7/0TylAls01
Mpp1AxSZ710MLaHpfn3tmXe9Wlb/IXvGGpAwfGHOsFy5IZQ6sUY9Acw11vQl
bFfx4ux8qja1AfbJEqV2dOwldC/fj+y3Ab8h7J9ac9yemYiq8WKI0Ga81oQD
2UZJA/fcDBD7Qt6cAbAZyC2hJYIgb6ELrPEMvDr6e6Ll2lZbfOTrxWUudqg2
rIn1tpRVIHA+37tGer8JYdfSzmYIDsJYqRmZTAcEnCY9li+OPE+dxz0vA6C1
976+wcjeIALkRDxaK9qXrBA+m+KJ+722HYXXLThp6pphGA93c7r4pMtaN3vI
frqAlDu6iszk5VkmlrNj52WqH5j7oLtF1YOLMG5uNylFIoMtSLeAKy1jMzAr
L1xZtig5TsPHavvBMx8xdxkrbwpuh1+6nGwpp+RU9tvy8fF+kkeyM/LeyfVx
TfF3XOVPoshlFgThr5OpRh4teNPyrzQWyR3L2riLpdFNMUQkQTMlC5osnd5e
95Oqy3LP9Q6md9hrRbP+sqMy7qQwS7VU3yYAGYqI444E5oIJ1ojfh1Hp5Mx8
T6Rd8SgMq2PF8C923X+zdPasN7Cnwd9jkxEl2bUPcZ+nzudnnyUY4XEhbkRe
gkDDulrVipbslGDCRkIIWCPbJdauH40RqQeP4aop1bT9jNkjt6+K1WARZeJi
52Z/aX7T0yOJVHRmUnSPxa1nlD/wTGPcS5ZWNgozsViTAggW+BYvRW98I+pK
c1weUs+pr6SBcdnbfE2wDBECMwi9UPIzVVr2wUBKM3jh8IlJWFeBmpbRlpgk
VycZO1pOlxoAc6qVr/1pq6tHblHmvTbc7hDh8znHzywG+HUP3jtsDkNdGiwa
i8462tOVDKsbuUjX6Av7799HtLiTAKjexF9XxKHgup9RdOfzCbwPlVZcchVP
3dDFgS51bw1kZJB0JAT5NSLncYwVy2f6XyQanilhm/qly728NiTNtnc0VzzS
qxyAB0v1T+4uvqyJE0Un2H6uQ26BMCcvrR4qePrqK6sTefc9WI0PiooZK546
PWkco3VWtxB5i+IVwAh/qrDzaWEc5DCNz+sJ3LqZMDnk0/N5iYBlL0zbQRjL
C/MtUMObdxAd97wv2abqqTQWwHfNMcwhzvTZhCfOmGU5a4L0tXHYgx9z6kuU
8/EVmuw9OzTWiBvHvgfEIfAg0LHBk5MiUP7jJ6wO6AnXzb/LzuJb2QI0X/+4
Mo9hhEjbE7s4pxbxzkX8j4CO05zCYz5aAduVbee4fFltaJOGvb6lEmksfOCv
qsHB4ylVVQ7u8wm/KrLG4oMDcFd7bQWyogblTkEU+TWbq5XwrtKGibm9cYl4
UXiDErCt3ZQz8fGT4m4ey4J3LSOSIYxA0Q3t4NWV/BLgARybbSzCoIKPLrVc
kbTXwFbWPbq1OetQt5bBYcPOUcVMgsJa/Av8wAM2sF5qH2Dw/5QzPEIJWQ97
yFUzGq1/S8Mfl4gcfT1+U8uZhVvNKEwqlZ3TU7zFimCY+fK3Tmcv62a+4x6V
Quj/eq8cER+KVeT80fGHJYAjGLj6AHdNPCnudG6M0lomllLWFyNTlH4gaOHC
+sSTuMuO1T7aDvLoUWgAsfaB4EjC3KgO7c6tbDz7YQOscbu7Hmtz3Ljnd+Vx
bkVX8gO3hQNYvGpHBFqP2a2OnWyTaLFJwkuSJN/VGIur8aWB3Ts2UqzrdDD/
745qsQbtTYdp9KBd9n91UsCeuVidOWgc5X+aD5B3Xnb0IlS24JGVB6wd4Obd
z803CAGa2YaFYPlcvROnyNhvgnnVnbwHLMkrEF9Vzttx1sJHMh0aE+1ZILEL
DeSIcJ8fQH55CLngSovx9DZ9H5Jfb3fnxgo3xYyEgUQAjRt1UsMKULIv6Bo3
YDeKwOkMe+LiE2El0MEm7u3Kl5/S99NDyNzWLxCe5u8vLkDTEjkZFvVQzAxB
+BYxhDcAy1lf60bTdGCOQ+DZj2yQVhoQENnA6V8rfDuECIHGOeIvtnsesPoG
5uEFnCPZHqUmKgikYsLD39lIVmc7Oe835prY2eoRlUEiWc2ZJmKUQwfdxC3U
UXcnJFfveCyO8EhdydeB19CYdy2WaPYE3/Cc2lCtupjrMz2Lhff5uB0vQaoN
0xAufZ9y+OO9wDdcX7tQjzzjQABsROsr7Jhx44pRsLOTDX7ZUs08sTbqckLY
o1dEYX+UKCF2upN31L4U2fm/HC91LCquYXmIT9fAUBw09TDZq6ToyWCzLjcz
RMYEeKw/HHC/ElvkQKPmNZZuJ07OBkMNsoheGmU+MotC81TyND6tF1SI0CKq
1RLymD641j6UsoveGTizcUM91dDnDzyJV0KJd8mxqeydi9M6+/Wgf7t6D4Og
xtp67PKeZJjeFMtX9yWYp0CoSb0OVXaXOhvjkdrC85PY1U9I2dcUgd5nmXlv
9F4H1FcaHkE+Mg7WBK0nv6fVTy5QLB5Fteq6LVF7dkPZWW/7HW0j3R7GVc9M
m0PFcgv4FYHEEuUuHZiTjj9gxeTd2GQ/KQvUtJELP+Nd+UYSJD4GR5VW4cDf
+g1aWk3id+NFOLfx9fIieq9xFo5GoUwzMOfZ3GJd09HM4Y+JcOO70Hrd20mU
tEYK0b6YX2bJVzwrlACiDI+MAmkQy8qsqMmEhBK5lLEfLtKO7s1Uo9/nZsgB
0RSXcH5plqmQzPGVhQoRckA76w7a2XGmxAMjKv1WU6vrIbPRV42a7sIymB4C
eUJqmqqY66jaVEY8J5z7hR1npr8CCJt6w6YWsVqlZrbV1BlaeCXWWl0WJB47
q9plyyZyYQ/QO7kXz54MuHB5LGTWuSxoRXJsCAEs186igb/9nPIYE+gnDiYk
EmzfbNaUKUWRtpTqaoMaFsQpFrWrczLLiAd3Fv2CjB5qiotBSqa5hS+o0fK7
w5Gemh7U2GUgeo9Uam5kzAA7BTKsorG1AfHOZtHj+gSVU3Li3fmYbEY8mJAh
XdPRupu2yzzL6MR+PrH9GKAKghMFqaUX+HkBqrFSx744Y5R4H/3iGAqSKE2w
HyPy+atLth6eE6YyJgkWo/oBRRt22ur+Z9djtH4p3qk4ZmDKPq6543Qb5cO3
AYkWvRdpPOWWGtJebU3h7fpuE+0cl1ax9Jy/foWJLJSW5KKTQcsx0mhZvX24
K6dQFE6zb0tI9NgFLTfdeCd4yLUWtTKR8Dyl6XC8yZe6qWUkYkC7wLtdE04A
CCcdErqd08UOJLpcJASjCotrXfyBDUr+YyMHt1CKa5sW85OskfiXKe+EYr1C
cvT/rie4FM4+QhKRFFD67i82pQNvGg1FhxDMaSgTnl5cwflcAh56IKTrGTma
HxG/wLEIB5KOpwk7iGwTDN6IPsE5li+/Obk2KZObXzGVXuq+ZLeh0WmOaix8
1Wqu+Wb4YsrZg5dDSXcKQfxhVMIXGZMuuVpEcGL0w4d/VWriZnmaE1RKaaS0
OYSx0SGbLZbIMoplwVhiU65rgvUmGOxTQ3P6GIn8IxZw+4PLm5Kc27p/Z9Ax
UBlvrr8ekZPgWAxhqfUVjc6F4hKv155T5NgjyFHpPWffGDibAaAPm4hekAlk
lwB755apFZpu/VL2TaOihhq0ujQ0UEFWF+lFtyxgPFhPEvD2ApYGB6nNvrIr
y2+nQQB+N2/Vq4SUp8CduXwlwNLUD6kE0PQ4B89nhCVxB63CE9ai2Vj3dpHr
2cvY+T5jlHTS5ffXaw/f7cMHNGtZHddgi+nhiLh0A4Cat16rNi2Wvtwj64mw
Vx4etUudkmxQi4rtKDnJhlHQ3o4d077CsoL0JnGfVBRXT3nIMb2tz9mKSDgD
vGKRDM1mQzBj5Qnmz/Y3sUt96YVjNwvqGfUPwgw5bM0vYMjKp2vOYgQ3mnOI
u+aGIp3Wa+SX90SdMIpasTrLxQ/3+QIWzSZdXFZg2gk386Qw5ORw4oulDHAx
5qHJT04nJlXJTg2RLp9Z+L/R/eHCqmHG4jbvfDsCWARzMEpf23NMirGeivJG
276hFeJ1Xmwws5Zl81DdolWngrr6dvzV21MHwADL+LhY2QDXxc+9FUudLPWF
Ou37nFW91foYtTijHV5qPpvcr8ntnXezhg4TbExibz7h/IFUyW81iVyO28mR
pC6L9U37L114AYHYBk2yDzFHH0Mb3Fi0tF3QArSOMoRC2An+ct3BSMcbEvUA
hRfzKbVcWD6U3zSoPHI2eXVBmBIjEfDCA8SiiksWK4Rcn2cP/i34Nsjz2ffe
jaMkuEMZ9BhHNdhAcV2Y0y/DCpfvHZGniLK5nRQe8EwtgrnPSPh7r2nrr/qh
H8VN4cmiG5upYr00nF6bSvS2XFOmd0HZp8Vg2iTu7lfHmGIstzCBDzHAGcVo
i2Px0G0KTG6DPF2ztlj7R6XlyXqsH+v6NSGSR5E3e9LiaQOE1PVn5kEWfIZy
EEkCCFl2OgqC8enrcMq802jCAcyT27MgyVkI2XbmMad22Jc0Ph4UtE0rQI76
OUJbN1d/9tI1CuTVgquRcZuG1/D0UocPd4U9Ev/Q/suKDAyQKTTUN0JDZLt2
v9dKAs7ummWFiEd+nqqdtNMKD3+k6I8olZk+TeVopSz/V+nKOV9eLP23fFW8
V6CHKmRA6Nd4jKgVqGYUF1fSyjXdD546phJTDaaorL5hceIYulwzuE4L+RX+
41AHz3Gy2vrwMzXaH0vHPIkAekiPnUIQCCQ8A8K5rYhU9vsyjz2eJ+5qYUNw
vRbhyFxUd5GnzhXYcP6XWm+HhxNO2WEnoX0TOomPD4s48cUaj024SZTwzgB0
6eN49YiKAET0zGcESCY+2XpR+2AROrOntGkkivy8bwIi0oawatL+6SXasofx
J3VvIh638l8iWBj1LYAI5vKhqIkvuBbIBaTOHXkA6Ojo54quTbdcf5+yju5w
XOoMEvDFmC4OLEv/bwZ3QeZXRurgj5sIq8S2CjW/ra7PkR9RUcW+tHG6i7Ux
oLQX/M6NoaIN5WKJfhTRFb17W4fe8w7JQBN6ZBHFNZryicTTUpVS/4N0Yusf
A3sofam3UHWj89LH0xxDYdhH0clKqdasn+W7mUr2xU3i5Zs3W59Y/XWaL7aT
QuS4+yb3Gru7ERK8Qmz4H/ZEtHlEnfXWsWtbzremKWxtz9DalEStONL6c7np
zaUytoDlxHdlzB9Lp98vFhgV+3r/5jyLRuFB8LO3aJ6mz4jN5WBLGHDiMQwM
BYaJddSQNPLCE+866Wh3/LF49Blmnai7OYeEzl7zlDxKVKeeMMuMIVrVjkdy
joOPXhBrZbwmmjSLxej1b/ai4OI4hm0CtbMa7s5+qKDAwsIRBN9b5tHjtTdp
Fphy5FlhOstj/yMCz5tPGFyjUxgIzHJIuva/3VolXmx2FmosStphHG9uEa3g
YgjVXEQdLmXTlSSSd/Ygd0cvQhDYX/jcRwG9n8KzsWisJTAFl30860UDnQ7x
yeJV+FjkZcS7s4wXuxtI2pajDMcRnJZmbzxhjl1LiBPLROXsd029cUt0tHYW
D19N67H6ZSJdHW3A24WR10DMfj3Vjo4w+Ijcgx72nB40IIrS8Xiw6mf7jBW1
nZFaiQr9GXSY9n9jhLl3Tv7Bb8vzbVXUjy6/TeM/gTWl6J7onoKK1EvfS3a7
XneOqqrlec9IfyduV/kIoWYMHpozwIe//2MadbIznTR4g8zf5G1R01VQOADX
AdrIKGXoPAch4hPun2JSUzxo++gFckEAvFJuCMcClYGrJyCM7BLDsZwDuRUG
ugcHB/ux43ItGAWcj/FDxOZ/blzFfcvxlJ7ZghvHvZwtOv3Fq0RpKIoVGFIG
aL2FsDxrhPJJx22wnYYOWPNEUrP7e0rCZkdrwtxYO8q7c45ZTAbZa9qyqEt2
o9sDvkjJL1RMp/2IkU0ybi0VZvvJ7edLrqHXohCWEWpRLtkCCNYd1BJYjcuL
q+l6vBimTLEl3iR3mTl1+NZYu1rRdJA+5/LIwX2BSfMpRHHC1LNvVlbq/XlL
8l6AAzeaJ5rAYDcRibbFSJhFMcD2q2Zjw7eilSdUHNp6lr8p06oIRgbgVz+z
wLESG4aoChkoL8fcrSQJ+c/c5VWZ1fiRCP6ztEovUNCVDvTmE8PSUBAVpPwT
CL2/OIXgdQhEznjRn/4o/0DT/3GGK1aLwssW/WxRXkRZ2LJJ2wHQ9VcrrAiL
s2aSKtexML0+gBztZmkPo4dGvmuZ2+xGeYz+jTT5hPB+ZgvRhYL1R/wdhPrU
ctE6kmko9hGprejtXZ4LCrV7XcUSinwgCWKs4mCaYy8VlAK6ODloKt2Vs2Js
ZU2O2XVVSjWnv+wuWvwg3y0Wdq+sX5ZjDTxV/I5gon+zeJXmFX68xyYKsd68
a4Y/xZBXfVHZq0/scvDjcPWsKXfKFDGXf7S7NHrIKhRuHT/c6LRtgEzQcjzb
g+2WrOw70wIQvs2JEyqaDttDhtuF4c4N8iYfXLORC71/CR5XA3ZzHVRbSfjh
vnYW/kuGCBKO4x8VJugBe94bC2z1if2Uz+kReirDbMp89YQl+6+8/f6yAjlD
BI9Kn2Cc4ofUOjvqUprVRzVzH1W2wqGBxMTt8xVTTcd9BiOBeqYfQ12l7az/
JN8PH5OGxap+waSv0neiK8I9TeSnjbGCxkttiAlKVyeN3tzdrz7jpWXLwonb
9BQdvnvB9k7RzlkPloAVTBlVf+bosU1sAOmioVVhCHkJ8G1/wbh4Xtl6qEoS
1FMIE114EJsk6l56Y+sB3dURXoMH717+eXTCudqGZkGFx0nQ0TQVVpt0Avxz
gcjMLunf0Pd4ChRmnjbi5jAW7DQicD+DgtgE0LOBERO2+YU9wQvXASkaAlLI
H4aSPT3mO1ukzp4HWheT2Dro9q3CY6lsIPu4qyUhyOcNHjQCuC9AgBwaPZ2e
b3z8swLnFa5nua2o7c5ib/ZaOT/P6I6Xi3QXyptl2zn8sIYKJvQiDdU50KlY
/c/v/OGUyuc1qJYmskba4K8IoDI1fMKHX9Zh1e+NDpGOVdbuAv0y7wOhi5VG
ncJJskVt6ErzirjNkKyjtPsGcoQLb9OgLfeA0a5P+MQqgBd0pLSn4DG6iX+B
TLDrRx50PJiDx0nivueu+HUEsaOetFLqfyeFqBS1tEbxPAHtrPxD3d9caZNN
8lAuwx1yWykTA1NHKGBSTGqads1EHpQ5ay7mcGeMksE4dEs1pbxHpxAFzLoS
1CdyTcVfFZJyPgmisw4pw3qD4YYOfRrWgGlLx8YK7kN8YUSeXN76I4Y+keBX
jiayZnE8tv5DIcGOa3/I1Vp+HvRyirhbBs0DndvyewIS3a1Q46CuS/yC6tOa
JwplUcwVcH99j3lJHt4jyamVPYmsZMeMpuLRA/4VXk4WfymxEqm9McdSq/O8
jzIuz7PbdheMFB8lMrpR5j4m76/EKpfHniQbkePcGaxJbPNnhR3Dqt8YJAUz
YxJaS579VgCNfmpc0E9VUxwKxDa8WPnrAH4QMTuerAjU3W8hCGOfiypWpxEI
mI1Ga0UlURjqFLLIqn8c1IeJVG11jUvzA7o3hbpK1lKzt3Z5zHkXGiMUHxmk
CzSZQaNU7cX24Zumn8kzZK14aSE6JrqlhGedEI3wJ/MU1JE3dylXUpzoZv8G
yn4JGmv24hkn10XzFS0drT/OCfOt41O9oYNsulTyx65kKOGU4/T47J0d7zvk
7lWrvYdFPYJ3TNBNkVVDli0YQaGfF8AITJb/4FLXI+c5TzV5SjHB5BiuyCqB
nAAP6YdCLIbcA0Ax4j9G4NlHuTr8bvwNu9LtlfLOEf92bITI45pj88Wt4vCf
QfJP7ko9ygwqCJqyeRvM5wtoUkwcn4a4JgZCAxONfWuy5SDxPFjBnIBO8dXW
NETKBq6Yk+bXoMPsyptIL196Xu7Ccothri7TwLzHw0LyhxiUKQzWowk6qDjG
El8L/OdVhFxTvKfiX7Cy+a5a/yGddXg6aUwthKJ0WSFBVpIB1HyP2SQ9EGjX
IXe9XpLrlBguAhOLhB591XXzMKfzVmkhNIZLpgb6j2CK54cIKAbpckFlu3UN
KDwF7F5bhbJKuoxoiXumZ+x8fYGprnduN1HadpIsSdo4ZsKHKPBbnXKdYxNo
rk9ziWb1yMyu0EBiecZGAmO00JqaalK8JNPDVOe+F/OPdNhTLqdo7FvATK0I
qLyJ5TDMFQ4kTWu+chqmvCfoaJT7Y77UYsoT2Sw3ODp2E0RsVJM2QZlOpMHX
rBvRRm4MbrsFYA1XvTV7aEktaqHTYGdeKT820daOEsQy0y8oVJoBdXX4bhPh
MhUkoHPxQft0t8fiCrHjGmknFaI/xiiugBUMCzFiBmZGQ/7WfOg4NIqkzMXz
zSS0i+FQWpbG+J3iiO6AYJpdJ8ZciRyjgOq/LKEv9BZjFeCzjgluSj6H72x9
qJIQFwIF3YUxaZdb5UxQGtpA79xjbbXRv70cW6jiWUztpfqQ7NUW3jiy1mx2
6/UtUrGnzQOz4dzNDLYs3JhJ+FhBro53uTnPJFydvuo4X074q/JLD5VtIN9C
EzxOOvLwG4x2i+c0ue6nUrx1jeTJHf3vA5mkv50LwPzehYpsGeaaWvJMMM9m
oA7o8Qd/Gqhe+Xo05KU5iEuLnAC5q0tPX8jsxE28uMqaXheewU4xB+v1FcMy
CmmePQViYUT+DELMtFqQyBMO+Wh98fuKTehkda6Se81MlRg6wrFuNsRYaO5Z
w2I+ldQb87hyswRNa3pRz0q8KrZIXGdElpTBP2q3zcQkDDtAJS5125GelniP
IfAyl7D/mT5TrTC5pgA3RJap0CnC91ZXN5jWE7HGUtXbKfdwHyU3MzaIq3df
1iwX1a0yHMvsSKuezehZBGF42kcM13Yzzmev5Z07X7fqpgqbO0yEJoGcbDAS
hyDUI+mEXG1nqtKnm8WFPVoTCHHW5qRc/MBDGLFCLYKwxPsZIeNKA3VSl2o6
nujD56QjZf9FIRLbhJHAh9TATcqV64Pt16WDzmnY8b7rTu+9AiyMaDeOqZEf
Ou+wwd51+HPLOw2c9LarGD9Tldvjm/5iPiDufBc6AvinD6xDtvnjZ1dQtRZB
XJ5wjq4B80dTI5f+FvsltwkJI7TXSVSjj7NT+40FI/9HSysDY9Yr9Nl6kZYF
oG5DYF2HS3K9qU/nJEU/R/V67ckqMIjiLWr3C75Qx4WByvHODy2w3p/m8M43
7Kv0j/R0zl4d0pTf/oG06F3RnYwwh1kU0grtG+F2CPvWmd6tz6ki0r6XZ+Z3
Bb1O+8X7Fpv6SliicNmEtGIXp72EXkcFgRNM1c6byiFl4v8nrki9WPUCsDI7
x8ucACGU/8m73KvGbQV/gMcCE6cWm2a8CcQCpRtkl/OE4WwKDsENUR4AmWMg
dEg/aajdWucfrn4+x+hWP7qyt4ahJZLgNlWSKehKI/NdnGyGr4Z/4NzYsu6o
54y6hxd/NmpYxIycw/RhPxmOmq7mBbLWqZGyDS6Df23qgT7Ns51NOd8P81Sa
iqTuCxA0g2LJK9vMLrr5KcZHUQhW/UiZ/KZr2lG2e+gGaO924YIld+U1FQcy
vW4Aw+GgPCAmOA/J0N/FWhNV8/1jtkjThJss2ZxTQ+OKeRYirGkKuBQPOwq2
plWQZM76sJzJ7tgLBSyV0I2+wC4mGe/vAMh0TanN5xSMqU+b2ODAQV7Gf3ZN
aid37MAl7Gm8KSEXaxxwhfX7CoetOChjcS0x4BTMakVtVoz3Dc2QYILTjwEo
XVeaFdJb82hnW3/VV6ttUjBcpZdq7+aWjl9ZilZNKp63U5+BmhaqOI6fUEQ/
XpjVlNgwrLds68IvrTaKywQuoYeZs0DOxwRhBja/ZohsmHOt+wiuW4ME4us9
fKapq7SJMAFV9Zh6LmglEjI9E0VE8qEnyINFlE8QsWfTCaxUU9oG1aMNwy9m
7iEnv6iaYDe3k6yqfQsqbXNob3Q77ubCA+hOzZ0gQxeLwZaRP7fmM+8Ldhhq
RSA6sU6qb0aZEtaxZ2EMV523HqCzly7h29Xl03qM50Xrg8Y8GIDChZQDSlKd
6w6nt8zMABUFwrLRhzlZB2NkXzccy4a5NcrVa12pZJ7Gua7TZxQ0eRaXpC5E
Z/rdp0NQ07PG4cztNqddZUFqK0x2oV1kGrcZ/UxwEbDq53XnpuPYTOn+VdZq
O+e4v5uk3hJ5virJL8srMQng7mtP1dGTKgiQFAI6NRt3WV7i/QvFst4if3GS
o7N4DmcBDPWk2BG6ZUE7+sq0hkscyC6UcAYM0yupGbBG6fVLfYPjhFiVbYa4
sstgo0pyKUBLiJheQYDfqg1oxozLYriU0HuYl6V2zTPVoTr96O0GCie2XLlC
CqIFrBuJWO81LkknHXNcWdzDDLler4CVG/gxEqAsEgVkQavWBYt+GgoA5HQm
KcciwFoRXIuqVHXT3RMZEvMNtpqMpICSWtsRM3CUhy0bwHwSFWFKGUqLIv0Z
zUvB7yCyymjoKe0qdkAhBxK7u99R2Fuhth1J66zXeRSU2Ia9ntCLRWt9dUUw
LgnowbafYSnw2kQuHAlxxw0/IKZjlmNQpCiJ3bbM9M4Y6uePfz2sUyo+iOl6
x1qdL4YNwH2lL+C4rRq7y9MF+0ntb0TGz+7BJIgbfbxF0jltP+Tlj1wP+2rE
/JCjzZELmejj50FrK/GuqPJZPOXDuO2fzanoucIowebryrt03rJYn2YpxwNl
eYsYB1xF3tFMS8+m0+nuMgN4vBjfVJc0gJgUETPUAJ9AkBu6bs8vTCurCkBl
T6lB15lZiYNU6p1LxmBPp3IrmEJpfQv+yr74fL7rvONgTgupFQ7DmgvDQ604
V9FPc5j6nyLO9opLCyMcz+00jebERAk5x+TXEpC0xcFc9R4yvBH6bbIDuABB
hi3hjJd9m4r7KG+z09WBNzzzS3lT5BnU3Kync8zV60ADrsbOITHU75BbgUIa
VEBftZW8q04xVqF03biJ3/vHvuXBX/P9uvZ0pTO95RqDCmcK04a9war7aKbf
uBo5YR5RjY6CGtNc+c7zdQNM7KBJnU0o3YQj0zHetTYdVAdX2do4JKPYBM0D
Dh/RL99qL4iwpUiruq4TYr6FIEO6NfJ1eJ8m9nGkXEwHwh244qE+EAwbYBZk
C/tAkOjkO2bUpWsBhiebzSJOAxzHM5anZrfD8Fb+kLYD1KuJqcljep2Ne0L4
0/0XZdGMjnty7JFDwSxoVHi3olsueqM8ZObEB7GTQrTwrYHIMdpOw9ZOzrD7
tfZUTUY26wEcKres2G9wUfsr4yNPVL/dTiFmKEHdzwLeoAxNreVhmGJZqzUa
lyCn6m8Wog3g1g8vBtj0EiNkYtUo2o5SN4/l6J0GY6WueyB3EE0RGvo5CFj+
Wr1tEBGGOXm1WX+W02CPtF+IqZ1ELG/yM3LY3hKOdevXFe1ULq0Of1aOU9Yl
JzeuE+6MmStsVmj8SLR5MYIBs71KB7yRp7L5fB9PdVQHAKLByNuNH0ZSm1eu
llb/tTvzWpWlRfqPtOEPF98KSmD/jZgl8KXMjrFtChZq5lKei2HCZUz2zwXY
ZDlwjTDJ0El+TdVWl9hKlMT/9vWHr1PrwBiKM+NQj2Yx/5sQ98iMdilqeUK8
TtHvxg3S6bla8qbK/JxiFbdKwE3Ssc3mUFHhMxCVCYqQAhAPf33MqQIXP9tL
tplltmFj4ZxC16kF4PR1+J7nrrZtvnzZJ7iVS8jbCzPjemGhivmtLyELNrsV
Vzl+Xp+8JEc1hZYjY1PvNXBPkEDMFw5qCyKTTGt1DhjZzGksMBv8+ti5nIMB
aD0AmcxYEUTp61N+LE78qzM2RU9yzzz5Y4D7NI9MyI9tWiptq8Jk6wXoWHB8
9HMHZdCCmDzsdaD30L02sedlqXDFK9AO1ZwFbIm6jVMHiGCxOi3c+UHI+cA+
nlZIPJeleaHI9EAM2uBCbpR1fMHHlKKt2umdJGdGR1aUw5eB04lVFwDNvSlX
/2qtiKfXbZF8ccQVguwl+ggEJCYL2g1xuioY5h1H9YQLOteGX7/2HWbsTrte
YfuywJQO7g5x+DBayTYkVC3d1qctBJkVbcQy1lU79FJM4Akz1YtPXCyRQIyB
tWSZlQB1Mw9go2I+KXz8YVpYjCWiEzvH4RfNf7EJJy124EbioaF8gSselsv6
zZ0qTIbyXsPNrYGc4jH+d6aB38d1OJILFT5LmaM6IsUMlVenLldRHUjzZ/m9
ePk55WncHKt/b0NAajp9PbNovpeLXOSD7lyxDfAzC1M04op1qFVNbRNkemEm
dWTSG1g0zwrk1+lqAd+5i7WvNKZ9qM8AWsgfdulF5ByI7EUcND8/IezIPZOW
xqUBF/vyE0fGNOZc+b/SuOdC1G4CsI+hi5Tm4vZG3HuSJhuJXe0lXg9Ae6+i
42OEnD1wJvBeQOq5kaUZb5G0xBwT1EpTL3PrgcZJU1XdHpo8w67XtY3tVj/D
JwNykJ9hLCoYNONQyqNDgh6bA+/7T1E2O4xK/y5VviMWSQCsoxHdTiGsg4zI
u4pXc2BsfwpVPDQPTcH83mW4viEcrOVcKLfrG9Ps3f2+8CWJOxN6aUmI6+jE
ZhHuUxfNJMoR6AvaVAzIOSda9SiXHef0EkkJc7tcj/p1Y96ASl90Syo6KCwP
0roR6XRtoI0zYeujBwugblw9qmhZ3eskR9eGQvy2Dp0f1FmWFvEPDJma1Jnq
EgYj9KkTJ8IUMhtgJ8yc7TNi2LJu6cHZ3jRAG0ZKye6Zb4rbjO6mWKpRUbjQ
TzPrNkIwviFupL+CE+c5lQl9lFXmW1w3om8d3it6P6MhEZvjCudkw+s1O3ev
2O2yHgeOKOrf6BlhXf7WcwMf6id2fZiuTTvZ/yZN6vP8QlmxMM5zD8z2Xl0v
HOCAubXeC73xX4DR09cX6QModcTeIehAI1GtoYQNlzaS5lIxKV7L7DeXcC6l
LadZVERazAklhA8RgucG1ZijalPAHiQQM/fu9HqwfKQay3rE3E2Cq0pJ+e9A
mbhS+trmYipVrRsn0VbfrE2n2yPyxTYsGJ1AC5OuSlHoG2RUpvQu/A7qA9s5
iroZmmm+IQaoIddbE/VLS1vMQosW56hB0JpkEhyJ5E9Kos082il/TXtVSgbN
WeXvzvsx0DpbepH1YxmOakSJbFRCuwj9ownNC1j/lUEwa3JFBVN8DuGRgKh1
FRmGr6eVqzF1wGSDmWAZyg5Kc99wAYzj9zyycBmKJamove84fL4UYB7NPt1j
DqnE1Iua6N6OXw5Nq/jcvf0Xl9hr60SUbgZFhshAHhAx7WV/LE78r5gVx+kn
0Nbz4ogFWVaZT/cp7GvAjRVJKlxDFFyJiNhSPl5AToRnJMprR1TZKluRrnxd
xO8d3wmIJGPOken8GcEHaU9cFGULG3726QgwnYlrZvlgaQQBqCxtHNrj6ez7
r5zk8XFqDsStdT2EEyjdMLnHlKFoTau/A74Su9ArkKuGpCITg3/EU0kK3/2a
1R/6BuMjl+DNpZb9DlGWF/odiNS1eZEpn7zMJgyRalqOJFqTUJpe3ossCcRQ
HZrFbuO0GO+Z6zssOQBxGtcngS9flUVhWq/wHU21K9fhEvHYf3quqpVD1Tm1
7pEvlXK8YUgHdxrxWNN5MSWRJjcUSp35yAsiWKy60Swyod3S4+nNpoaoyj40
RMN8ywfFGUYXPCndxY7pZ9mrGWmZlgSUofpzpXaP/0Dcl+UsRMdCF+7henjY
ERev3WSO6QyTl2DHVr1G/6N89g403vbxgEX0qn2xUXQ17cxGuri/ca/Eoh2R
8hUybAQswK6TGLM0tuGVDhAT+ED2FhOqKuKbhDsNzCVk/sh2Sb6yhGVc7Efo
eTBYZl/h1MbYRLJg4bY9i5Det36oUaTvvABIs1SGwe+/eaJAxoT9Yaw37hLO
TTuRDau612VTy65IwuXeKBnDCaoNNuwqOafjA2Mhnrzpk/INZaCZyiXwJwSz
x9yhxplJcOcpoC5A/mteum4e1gvEdeiYZXch/1gU+3EN+j1UI8N46tDi+InW
WXqNYZgk5brHwPVW4MahOLCC7BG97GrfOaX6JyVlbkyv4gGcix2yKC7G4hZU
F5rKzXDqeFqIQU2A31EUreWfVHkVFvgub5hsXznygNx57/r1t+bCndL4H3TV
GX/qMcwo71NGzBefjU/ztpONuAF1QAjT1NPhKaf3r/AphGsywFqm71V4uCY9
fHvePQp6O7XHq0Df4+BDnUtY5B7HrBWUeGwqZOVJUMl7V+W0gxuHxyJ8ch4A
0f8bA3GLdrGnIghJ0zzxux9eTVcTYJ+egREKlNt9Rzv6ZCKAOYuSwM0EQ19M
4u2Q2n9s00yUOe16ZMhNVmEFwksJd0jBqPfn0CaOwVK7gatJNR+BqLtnthWw
TDcPFkYya0XZXmw3vYEWrQ7yQPux6uWdZxNEN0pGXG0UQiWBCaIaA9VQbTec
agF5udInmfYEyICF55kl1qeKF6wKfm0nOqhbIxyzvTxhFcAjAnte99CyEGBW
QT5dFs+HMcUlg+ZtLFMGANTREmiK283U7QbZ47RZ0fVRmvmJnI9DEUfuR1H+
MdVx5Tg62K0REPuob0HLYWScNb6wU9/TVn8I6T3+GZk3n+8jVswDjZRceQye
mi0JZFZxzHktjiVdoH/gS8Po2GRlYHISyz09PMic5RTJNo7afN4wMNbJxPXr
CHcY/1vOkdqmEBDFk6ih+NXNWvV7Rj5xtQcZ0ElwBHrn8zh3XNRb4dIpr09c
wkAwDLtGVftsXkmwzoZ6MKzgCJOKsOQ4T1oxVtjPJfY7zBQ3qzEgmgEnnOfl
/DxoRNciRgPaZkfRPVbfMtrdoeNQ37LZhwY51PBcpcIdJ6o3vwzhwN2xRK4t
nqa3o0gfvalQFWxfKAcC/doCUs5+0owJCr//sqQHDcp9EyuhX8KASt30I4kV
JAQ5eWBopz2a/27Pn118EkWSQKM1w39lGA6Kn+jAw3dNbUCk4IyGDJl+1aBo
GAcF+/dFTyH2uede29fBlE4Fiuy8LfqqZXhpbJ1lcLb5Es+bs5dotqzMOUdx
p9FQ0kUK9Xe+TzMQ8Frr9dxIvJ32jBQWVwmoeisXmgbimk0C/eCWRVl1dBCE
UoxSX4fgqScZe5X3swQYLBrh+LpJ+pLhQyMG4ZxZ2y9+0ghoe45ZQjnwVanz
9dJqyotrywYVl7Jbp9avYA6ofQvkjEwkzvn+T4tNSAYYM7iSvGOpYoJpfbNN
nBN/tRcnUCCrHLWQ3eL1H/bL59c4jJ3N969EWKw4WG7NGZjAsV6OWqf2XXER
5okt/GFEvuISzuLj7ByqKdxljdsxlChh+rY1L+oA4yKTAh5J1q8+wQnlFfE/
aLEdvCcddhCJVW1r0kg0Xmp9JVtjOQuLRyM2yZNoYqVUO3eq3VkWe+g0W95j
w4ET+HNSp6zO5jP8rk9/EuDbqUFK3pWTwL/6SmJmU3CJBhcIQ0lm+0xYchlb
qTeYkb4U5G8YSeaZAnGm5kH5KETpqj35aQSyA1deSm1Ynw5ybMgj7+9YXOP/
rAvq4Xd+Mc2zrLjcy1ORV9M/T7XJa1DXORR/rgdU52bWeps/mkLM9yP6FgiP
lqUPI1zhUxH8hxhg07V8Z6dwGYwTCnd/RiNtxUDmeqJFksstt1yJm9qG3GEM
CewPqQqNFaqVTHGOYeZo9UO38FBFlOizvG9KTayKZyn4BXWboXzeiY7WczMk
jw/JSTRKPbAJxyxw17lRSAAJFSiHv3CQWdRXRhrju9DoqyvxS3HLKPVUzpGI
9p32k82sbWohyg1fkOUTb+bPKyqk9SkgKcgrUqY0KSFcmV3vjnwfrFEgKG2G
EwOKxswTAQ/QUQKRxTChKrIZJjeC8WthCFmQ4IubZdwiOMAWICxFT+NVhaJN
rrMSpse1vWRydqhsjP7HnSq1fRiXCzg2vnvMmfFWrMF/JrZIhToWy06ZaOCf
8+39nE0qEsNFk12VTFz/5hdZbc+e/13CVPWApLZrT0SZHB+hupRKsgVrVx5X
70zh0SNP05mTR1WnpInUk4FN1nnR7hDmD6ekUbSr3SDA9Amk946DNjh0mqnh
zBLnweozvLdKtuivX8idGbjiJMV24quZhvZaNz1JwXzz2KNEfsss4UnOXs22
bkfY/xkPPYXteTsjJkx090uzLFN5BpX2YJfFrbmBkyuI/gha5w46XZWbhuxI
5LnEhK/Qq7k+BdmPDGDpDU15X/2OpR8jGQmtd0BmMzCP1/MllAKQE55IdDpk
O12CHmLH1BBSrdZUWQ/tMbRhyWHE+FedR0qP6JUQ6q9ozEt7ebkhCR1bgKQo
cUjONDTlT6vS6iAGERoPk7FeQHAtT53IMYGkyOXy3Y+dXGltU3x1xl1owV6u
4YohvDd29LH9r9FYM6d/0ONGgrDoI2V3Rl8q8zqr1p+06cW6V2dXpVtT6ZCH
tXVABs6jXGqdMSLs2yFWFBQ8xRma/lUZ3/PeUWSWm7qp92ZDmKkmrUm/B6HP
BidA4/BtswIPuRYSR3nsmeJ0FqiWP8QClX10fS/3Xjizvp2yL2RiJCpf/mKZ
RbtI4JkCWL5aUoeulh3MfYkVB6dHOn89bslToRmmhdLzyzWimhjxHRtgVngL
YwI7swA9bXBlRE/hLCSINNxoH8PwoGApgvYtKdY9dDhYYvjh2B7WGHxkqUsc
7SZP/iBnjARs8BGEL9DIp343P2IXhaZYbEhOAVfrX3WgDS4scK5/bhZaJ2uu
KMfvwL/+OCnAzxfpZjIu7kbvycrSPHgfjZ3oxoAsZC4J9ygwMkt1oPlv8gx8
VaXPEjGpCi4mgmK5zySGsxNo4bEI1L8FfYJHNvzNVPB/YWgh1JzvkJw1ADA6
/jwLeh+E7H/Pvntl9l6MBEhiPrEigoK+Ev5maKL9lZtzosoS3MwtjYsoQZrd
YB/eIdDdeQX0TMZd8GcEMw0ZdfhQywNn71taMtjZ2ZdkVyAnXczaCtxwQe5W
WHGGuo/eUAgwe6usmmhSzHXzwrwFIkXRFApvF9r1jWOTFKDpK9PUewHpnTo0
XCuCnepmwOolJUsQG4GqMZ9LPIJzT/JPmSo4z/U3stcVMjx6L48Wt+J0G1Yz
5k2VqKajHqzWa7IHwrbIoJ/+aNopbrMJRlH361oEztCnc3uRQBQZTme8B+/S
Nxzoxpt25uN0pZOYRUZpvyTX23/m3eElWMJYlpqT6VjJg4GnjcBJRxT6SQNZ
ySR8urh2RMf9BeGKV9hPKRM8f4r7IJQmuT1nEZEWwPnKJjF4Gt2Krr+W59ZG
HMs2uJxxDk+nazvbgFfEFGo+2h+frKrnvhaN4KqGdIToNAvSPy12vpKEYlqM
nqNSmW2IYdVjWzHsaS6+uBoJS38Iret0qO6buD9IL+tnDHf+cHMFOHtsu8nC
GVASNA4uY8kjXM93R/n+H3GW8aCbdPf/rEBVYe6WjyCa8Zt27Zzx5YyvAC2g
cs2PMUcLZnu800r3rrDmkUpaXOzg5qj7vcWKAnB5WXnlhUACwHALsCe+NDgn
TxHTiPl1tDaeT8MqF3YUMGzL35PyWAgcNQdvAPRgJKqCdxIVcRhY3cQ7d20E
Nt9Pvf70QcbJ/Kl+o0EhwAWgFbKk2S+JMVBGxbCfwlEZJt7WZ/2Y4/O6sQ7/
d6TFlKuQKYmFv9tL1Ek8YZUEDHstqTXOTv4BX9omEMLKMUB08S8snAEcDGIj
/vMJL1IWcmlGEpTHlWwCfi8jeWLOcfeZdt5JcfZvsk5PZm0pCmIUagDV5uWr
VJgQBo0rHcSiFuvklTMVMWEG0SxvRCG0U9o+9rG6wbyVSmNC8LXZ4YMfNJre
nD3dqKlbKePKw2UyGxroy8uMSZkvPFXpYj0+RqMdZU2NjFlZZZH80gR+OlSU
TvbyYOhL7l1kck/dWWc9ptmumMsuvqY8o5rhvoFm6k1vSgbW5MaRhXw/UgVj
Gsi5wGcPQWjTaS6sHN2UR9SoTL3tjVbPT6JCdStxeFzMdYqZMwvFuayZiIXK
toI8sSRA5cJtpplTDE0RKXZ7h6rWQ9ozAYbzX+szSwQiB3dBCMf+Zpbb8kG/
3RS0WYRd5AfdjC8v/ssB4YfLbFFSQKC1eC0Z0uTb+AdGA7mPZ0a4hjzWH2/P
ktL1kWMw0LCkhpFtsKQc/AGHyHTSAN4B9fhsHb9p/foRVVyEM+qwT2dcGlB4
qqb+G83sE0P4knPnaYALAxypbhUB9XQ3xXVQuJMOsso7BjaXqzFdaka37lqS
3nett2hu53w8vcCvGBMu9qP44kHk2IrHOH5YikRBUoNgp6ntHnhYTZdFH6tf
QIYZvF0hV9fibZ3FBwKPTOC9tyc6UpI7XpF+q7LG7Il5KZknyvEqc1lqmtaG
ZG9dI01VJnXipleHI05/lxM9HnjGz2XA2SDL6pgIkWfju1vW6db5Kd7t11+l
PDR2VClrv35GphLvRd14gIqLrkWrztrttuIDKiCE71RPoV7nLs5YVAXziswG
+w7evmlUbcyYs3ElrMV/lCV87+YqLwk4ObNdG3PPoKxvE1Fosv4sgFZNYGAn
KD2LpwNjQ2QsPBXk8DS9dkXq8Q4HqrrY2Eaf7dkLtobE9KzVhu85FK0NfOLp
42qa9vtFeKfpYCsdMKzqGUsXCCxJ25fhMpz+6e8tf+bSjCJDbXQ0ef/lRdrG
WqmgfouyFxrfvMzArx3ru5ucR2+dhrHg8XedwW5D8dKGQxNJ36hcJ8zyIUPY
OcillYfgrbWAsb0w7ZTg8BIYjNowKN4F3uyVpoRvpFA7qNgQ0YZ9hf+/WKYE
4ld6t13rRmUHd0l1m6tFzc1FQITCyGKj4KsmC7QkCbyv+jv0OQkJiy6ZnJoY
4y2cyOdob17svASqenD/BtxN6zOLap8zzICAXoXgwZO5bvfsXTGBrQwPmCRA
OQKOHhhr5rA/iukwFSa5YJy9+ofLXtCGzinZD1x579b06ncjgLbQncAJK4fS
1IipFfOX6PKWBLTDVD3h3tnhUV4vW7kj/8xEV+7okCWiEKrRJKt8Ly4kpkhw
oWOkOC0vXkKhuCmX4TllUXVxesT+h6FdLYDzYe2WicIYr/L4Cw0HgnASfJgO
Fmx8KL8rveJ6hYOTI/07DL3PYKQa2ERUiWT/HRnvhHF0fVF4y/oINmfgNk6m
FhgnbKrqDiJkbb709Hslm+1NvkD7TSzqgaP8jji4pBFZ9DZApvY6SJFikoTE
gwPu6k95m/JPNF/x7Fs7LdnJL38wCLTpFi6agZ+toDQpXHsu7oAqI2JmZyCk
cSZzmm0oRV1uLOBPRv4375zJB4ZM9pe1RsBy7FYP/1kr49IVDsdG378IbE6C
mASH8P3GmlaBS5ONaOh2EF6dAycS7B/xtOResg/pvooUBmBTKMEpFWeVw6Fg
tDRWFBRJ/2TvpCsJntM/zC9q+JEbjDrwIQaSxpbfk3LPy8a1E39r2OFCla3Z
YqadDhUlfbOJCyzv7fJs/jH2HCAbfaS9DEyXkej+YPrl8/a6zh6Npgr4boP4
Fkt+kQ0vitlH/pHRUJ6cSW7mYf8+llkyzh3QYnQT9XajR+o0hxEw2YyzlN8p
i2AITi2PrDb6bSGEwdQwqRJGR9e/H4cj61MyY0ABnDaZ5M5j4Ft+cRIQYWlk
5Iwvnz3WsC4lnr/YCyTHuA08YE6/yvXdPxnycKQIQXfN2kwe8c86DBI3jbdS
3g4Xc8ogSNZm15ee6Q+aOPicGBRguHnYVsFFk8mBl2bemjUQQfz7TeWrzGLt
G4C+FmDl8eXqXxeoCxEEEgPAgzFWYKxprkntM2QxuKZxjZjCl6yE/NY+XAKp
EJIiVDMftJwnYFkfYbIo8FIf5OVsgxVyeM1TWEMmBDuNHRSQpcfwfSX2QqVu
h3NOrys5y9m37KfILqE3WdKcJIFQphiv/xCS6XJHvUrclI8puceblpTzmJYd
TfL1T7u36ru5xCp716x8lxmuppjuq9jmGg3uaEq3jyX5xtrZJV7RUUr0ilK0
3u94Zcon4hTfO6LmC5lZYJFHxiKqzhnTH29/Z5ll9Ie9jFokjkq8UD/ge7jD
kwqFxJPOoIGa+SFQDhyHcTzvYxE1NP6ZRTtyHESYvG+MMx1/tdUeAtI/bp1F
yKQBDNGudC2xVa9G9xomcHtTJA7ATItUc0AOtgMutVPmsvi+jPWWTxy4ADsM
HCZ8LA5uFGzmAR9i/xw5viE8d6/1JPL6RB8YAwjrAHaVAj1Clnh9wuHN0aBm
v8p7cruK5lmyQ2q0+TONxzhWp5u5tXULY0eJiMMehg/pQQvEBNjMfOWko6+1
45dHoU+Cd0nAKfbYbjQo9cdKCrVYsuh38eHSIYCnf2PaXdvvRZu3+J7rxF+T
FmOnHOZAfRHCICWZkcx+klcb54P0YEtkCBSJmz9MtWbgJaOl6pwQr6btxJMc
dGPlf0DzZjacuHP3Hzx4FZxlAosgKmzuini8iLhd28asY9Sgr2xdABA8eXLq
Fr8xLojl5YiV+lI275XvMpF1rBCgMPs2bIelSzrxzfIDrx9LWCyrI6Ynd9+7
O+BOLqy1n+cXPE+8gGyJUkUoBQJBFGDTyjlzb0u6XlIJBmPK+Ny2/2Bu7iVh
GGHnwwr/xLVoou2x89FevPiH0oDlHa5zR7/GU5vxRCG4BzZgvNugXTWsqBMg
gWSZJNxGjYjPJ0hMocNGEuI+mJEEkB5df692lor0+M2wqSVnZ43v+70K3bNh
vhFZarsDz0KNzOtEXBgGaWUbGuwEUGwsiDJBbmdj4stw3i9b3UKpXeiM+Dbj
0DTbK0s6/yVM9U96ReomMUaioqiCF5LQyvFtxO5IXDMq7Wa2IFH7hyclWiYp
MKgKaYRyz3xFSqzS41LB4F0Trw/cIKlQkV/yhw26+sTlj0GVK4G3LVIy5XQz
cR5y8yInZMtJw7dNbk+jMU3+4L9wmJTUncA7Iy7hOLO77p1PQz5z+B9MbHI5
Eg8RQH0+IO5uW7S2cVIkHSs2VebYNGQW9JmTG9iIGp/F2FgVQtTXqr7BVJ9v
gcSDy7RjjWHUjqU8nRa5jm5Uey0EmnCVHEfJIldCj0jr8UnI/pLC12SDNakj
RaT1LyvDMI1rAtLoCjDyNP1BSXFO4P7q6VcsGUiFv+AYxUrz6oEtHoYgwVMv
/fG0lJUV1GGe8AwTZ9e7Pa5MLCU8dQusmYE10WoVXYZ+/KB1TvoG/7B062YS
E/RnuJUTcdX7gqsYcADuukexD8LI54aqF1uHG1CNNTxrAgt7xdSfx6JaMajS
OooFUB7lxarAdE0a3hlLoAw4qoXhJTpiEFTmnQJDrNpMRCpGK6nBIWecrHMF
pyE9EkQuA6tTGuVKppbmB+OCKPJVr8olVLE5MygiHUTbfHLt7lrnRxSBlqZ7
yvOMGg8Grh/P7WB4ycIUvRQED7WQ1Xm2eSZcor0A3lFdTyH0O+RPCGFU4REy
Hyw0DSLppmHSoZy3UuaBICA/hwFjl2r2C+6XMiy8mR/JqWjDzCPAIY7X8pVq
uE6CHlGQb08BUY4BhvKvi1w8EP7zhiOoP7lpC667hWdsQ/7rh4ibtvsSPE9l
P1AuGD+hMHjAfNjahnA7/5MCYtLgf3BnzWoug6NZBysjClmY7u+CVZBj9UWH
m+X3slM0fS7+pZD3CsWzXy/0YP7/6VhgDIOcsOQCXZTrFB4TgDOY0BK1QSs0
dyM/9sn6XXCvJgC57QiZwk+IkbOzewWo9uN+/DX0oR9Z5YRqwIWocUK3H/Vc
GxNZabDhSdyIRB6zMa+MkGkZbG4z9sPgOTNodSln9U4KUWvjOX8DeogCUbkh
maDqx3Egy1pu5U3sKKdothg0xgB8B8wUqJY2XsN33/1fhR8WtWmHFQ9qv+z2
Wo2GPAty2ol8/ih3YSep1FaV3MEKYRb0VTA3wp2tbKG6PNoo2111e+2PIzaX
ivsjHwhpUnmX+SkLNRuB7nAfOytREb6WrC5uhRLedfoO+RBJ+jg51XQx55o0
LDram+u1yrGiq/9AzTUHoJ5PutcAsyZ40s/keyEm4mETAFFxEnIqPErOGTyc
wLNK5bOD2zJEPH3VZdoqmY+GpXfloQdwkEOf/Gt4+2ubdymmxpvKXQN+vLrf
MWoHq8yLrCdNbdpNn3nlM8nVrvvZKk+UKgfpkxlFxj/zOvduo+6xJpNafn8e
mLxH8zjtMD4KhXvPmUn58TLH4k0CxcGBrvchCfVKHfX2seV57s4ic1+CR3VM
cc7vHxn9lh1kE690lFmIxGRuCuUMJjOWPqomLLAY/kkSOHZ+F32FU3IIEnsp
DQMLLlAU/+asfrYaSRys/HEjplThJ/RWWswi4a/zqGlqhJ68IXmyPhcEL6L4
zooQmrITk3Iu3YsrIIKLMoGa5U3zQ7CSgun0hK/O4tA5ljHoDn1x+BCYdgE9
R9mpUbyritiKurk0DCF6al0574orfV9vqLfMZDMhBXALstE7VkdbVywLugZj
tZrCapy6nFl8YEXIPfP8no1JIQ33eWdWFBKshaBbaE3o24JWk3FNn8rgdP6p
/cheBWCOHtTRm1So1gXULHgBGFqSlYjjKZ2g1EizDZTeE6NooD3t3JYCBfpP
krDL8HbkaNwJZXov3mW7lONbhB4bXgCAhyqbD9OMCGDpq35owr8CiSPy+SzA
7Y8TYihZoL9AaB5u90HS3Hrp/XkTlRci+vU8jeZEGTcyo5EsJZL6+LNm5ku8
FvFe8BhMZ3jxg3hEEm5psYE24fTszwPq9YLq7RY4/HHQBG7Z8n7+HUJy5dkx
9bJp65oVN6kWyY5v1r+wImGwikNsLjBSDOMF3tvRZ1YNsRU3S+xX9fWY65ay
VJL1Upq0kgGK5MUMcMewZIj1QUlGfrzrx6u1PPyw0Z58V3t/Xq5TSOt56+E/
eOUtD8kNSrtWyddpFesJS5nvmqAu7UfWVvhHi/TEv1IZYzsutUAKU1UksFq7
aNopKTYN6OsCgIHh9zSbnRbmo6NROwA9AZEizog8wQx0iiTj+5uBju15mfwa
mrr3Vx/USnnqYb0PspJJK/y677LDoqLngExYvpTxKmmRFZwqit6WE3NHjRbZ
eOJ8SmZJfOzQ/SjVEJyXCjMFF8wQw5Mz/SITVcHACyyW+FgY2fofokRmKILz
8tA+X2L5yr4fRFcxWVxi+FB2nbvWpUHamJS8a8+YoEO0kQS1p100uqKAgct4
Hca7RGS6gBOo1h/xbQ74h/wVspVpVdoigwXaTWSEdZt5B5/cpRm+H00LOs2R
H8TE2UcT/J2LYeiAO1jPFEt2VWPbK5PV4MEvaEXf9obPnjmFDYsivHEyqdwC
Mb4UXcp5b5a6uAVxqyGWe+z0YWxoTq09EPoPlUGZ2p9wjcgIEQRwidZVACgF
wIRQmO0owzucA1FGTeO7jtD8tYUsL/ltxf91mUhtCPijXaxZzuhUA+4SSV1m
4pWswTJipZmOxa7iQd4DTc84ONtnAM+U2D3Krrubd54KtSgijWcQ3G8CMuai
k+X3o4YjQBL0igNpj3nKdw5vP19oXAGCGipYxPoMIPGl/LNq29vBgOS/yqeu
cTkzGG2VggrDm8C9oAELt4XRqRYb6NYWA29duPHAtb6il+9yOBJJvTGzlxsZ
5oCW+06rJIRSoqwy7UIHpwzIpS7EAqXEDWOI5neD0tyqxY7IegejmtaiDZIw
eZd6C9P1X5TVYubhK9PwqD/ulufk9awMqJROLVu0/5ZrgsLs4nl4LwHkvFco
bV87/YEuyNacfpt7NXyJLjtwZzoTSEGhPZKuxU0rK7UIMWIN61874ZZqoEoN
1IYquj2ajzKMSrwwhEU/rXPkv7euEUxw2R4z84JGOFem8d8dVE02g6YNyUMH
ylo7yTsXPwwt0WppiDehA3EcXxX2eO+Xr6xU8M5sEL+BCKZUex/QUWP462kg
KKQI6zKfH1FJuo+Y9I+057nkOXmuYTJwpVSFTteC7Hzp54wMuGxOtbzZe1S2
wEBXirnvi23iiGPljFuiRKQGtQOLVoQYdFH8nFHGb/tqg57eT9erZJbW2z8j
46RxlMTExORexoV1JL4pKQrwi0sMmfzJt9yvNdR8DYnjzwm5RRr6cOn6pfac
2moJQEW5VAN4n0EzX/3s4A1jDkUSfQpWTubJJmKjOL3FRYwg+jqhlx4haE4s
xX90MIogLs0d6IVFoSzATImxUYfedtT6VXquy9edfm3J9+EsZWFV/X3hZOmZ
6C3gTpqN/sj3/aV0D3cyyAIANUjvTWGG2oUZeoetme2I3XYOaly0dueBps2Y
hnrDeAunYDjy2ZkeK5G9D/DFHnIJcrJmuCBKKi5mBQplVWKgF0CixXpDeuL+
LZEz4nu8Pi8VJ3v2EdDnTDhBbEJ8NvcGnSXQNTube8+R2s6ufCNAJSrWRPrs
M0TB28pwLQ+bOst00GD8piKaIGoml/0Wi4wNTKG37hAFengPtZOrfDAjm7eY
XXJBCfIn3v3x9ikM55urylugEf7/7SPErJwj23KuuCtEVXDE2yaE9EAdDEX4
DlOLe/W4gg3AnBxzURGOAcg2Ear4lT0U5HdbuWIzGGxRHzxXnN2jjKVbLwqQ
/mPnFD24NJABjE+IOqEnZj1kyQyB3IBGQB7jFviPJ9bDtF8PvDDbk+JvFVqs
jEyOQ/HbxInYOtj9EArKBgZWCSdSD0b+yCr42XlcfSwLFOLMnMpIziK05kPD
Gf05JQnN8W4HMot9DUMY7N42McPCg10bAw3mMeTT0z1jsBXDts7nsBxLH1D7
azqJPeMfsZV4NTVFbag67aJ1tzDplHCEFC3KfW/2JjGgiyRzDMgaNy7GbhgV
4PlZF4WVzmdmQK6H/L0rbHyY/UqEiWvdX/AwiyB+H6nBFWL/NLuMT3Cc5LyC
TyqN63076/Uh7BIhwHfAexf8eCMpqmNAiz0FNDHqz7u0ZhmB+0SD4JYsqUCy
7knZOH2hVTBKF/xOUlO+2nyxx4ftBTtwi0yHiUakEcKeqDAGOQfTRCkkDJLn
ZFQjTWvAXLTGiyRjhSlW55XZ5oxKA6JpCYMwXbm0G1WcFOetBn9+1lJf3vpT
1Dg5mwFNozaheDgusFqLu24sOGSo6m9oyC7P17UELbLUsNfHpG4wnzEUHvRB
WBm5NaJb87VG6ecYDhivtnLxxZQGArPSOBGl3I9XQ9J+Da57aB0XnWfxGBBd
qrlLVWEkMrr1b5N8BfBt5aD1r/ho5BKh97dR93EQptVbqXZETVAVlznl5PLL
EVER1FMuat14PdfBbFwANAH7JMEKCNfOVSewMkScuTEOEFADIMhbvQJPXbCn
yKgQNDjy7XwzgkmdXULEG0CfXi3tBRgFz6Cg5tLYQKLn1ss4qzKcJjnMy9jy
S0Xm3WMxM6Pblo4bZBW2QzI2R7NRh6B9tt6Li2vV7S50DVxg8SSvf7Aiz+VE
H5ZRKy/U07k4CFq2Wb8Od65YWkQ7YilADcGXm5gRChxc3BIzRmU+BP2BjbAZ
lc4QSpd7gIdMPhAGUbRQZIW3aMy7i52jdFbomXLsjazfp/+lI6iOl7u6ulAy
AkmPYV/Rim0dRewHK98bFlWKLxJze4Zwp4r3OpBDfTD8s1GcFEmKbnFPNG6X
GKOm0c/bmd/uVCU7UTpSorzK1TuczPno+mC5vxdRQEwKIQ8aCjr6LX81AyIn
D0f5QgF+k1CQPG1OJMd0Ha5Ra7GeikqX7qLQtgze9a0sCtds1iGJuEntllBR
8SOFac+w6GsTKBMVlZyuvXghuMC20lS99zqXBn2lHtQtPyf6ISccm/X24xdJ
H1u2G5gh7n/ZmG35yMaPN4GYKEsrlVh6glweaIAB736y3yRsChAtOo97M1Hv
k530DhLKGq+pfQNrkT3fDBErXcsBOP+sh7VYNfWmiBJcFvybZ61TE1c34Pmr
ERY5eitn3oKO9KMq5wLvCEw4hHiskRjeAvClq0w+fFjSDbf113qWFMloacbu
LBwASHxs5JNb+GMuMJ+oJxmHtpR0ZAxyWKvNJ9Mj/WM8ttUpnVHFIZdtFg45
cOZmdk2T2nWh2mDE9KX33aYvhjn9+F3RoDH1rUPjh4908+gN8QM4d5nzjkow
gtjfWYLmE7mUd8AR7OZdpWhgiS/4PwRoRNiuqEyJgOprfYmSlQfGG7hOCApv
ixsKtUpDuo7zBkUU1SQRSKCPIzM6+RSh3HeRTlxiewajLhyKZmvf9468Gslo
3CrB2cJ/+8hnEhZoGjhSv1y32LFYs0NCtYnPK98wFKt2f9Dqt9X7Uac7jjFv
WTQe9nTIgZMvaiivfVhRxduQMG9MWPb37y3Vq2+HaBfj32SPcEvKq0BCIFAX
SVUVLGkAwiOHaErpsKyBosWaLixxC6gOWSd2Gw5PTy5YzilL/vfU7v22SYhp
uZyrE8IMe4FhB5WDV5Afsv2PfDw4GhmauZto3Z++lJnP63FR9pS0vdWcytzo
FE3GJyTzq4ThiNQpnmTUBFL8Ph2Jxzr+2bHmmeaxIf7mUy72e0ypjzYLtbaN
HlsTkc+BMIOb8XOypZbmbDqrZP1/4v5oDk/9ihCb3Lmw4KYXNfCCgtaHfhnK
BoWwIElOML+IfNGRLpH8lT+KBqudTJIxnwKbH8qJff2fH1ApI7D2WhjUR8s/
/W4flPh0wKG/epzXzwDXyOInomGLfS1hLWujquwgTIKygviTDIziVwdtq0Kg
MCUwqfDRdEA4+X5m2Q1JQJFzVuHFhaI7YCXfjeRuc8zZOoahoo5D8/bO93/A
dXtUXcOx23tjvB4AG8kanIBComqemz+ItNbfAMOTOM5yKEwOxCAxMQMDdP2/
CkADmRQdqJCVVbldNg2B2aAuVy9nLV1QfW9AnQ2ODD6sTF7o+6RTgDXiWhLi
jVnNBc220wf2p1QXfigqTLbhOc5iM7bEXniWyYfccWS41qbH/+NiSh5zLQun
oHaHtE3Oo9BnzQvhMrJfy8ffP+Q8e8RnAYysifXqWbWPtSJdrbmhNp8VEOly
jJ9kv3+QIiBgbFr/q2m41mUEuk/i7zZonQNAh2+b2c7vjLwBkJG9GkzEZMDJ
sOvl8C0oWHvWGVECwfzGU+XS6ZacP1p893u+QmqhuF4ryf+0LskTMCdWUyWY
A3MQQ6aHsktkEzGAkoSiaDdwXmy3PW1N9yp5ROmv26vkZ8Wpu6wuAt0OyI0+
6sKoT2b9JNA7UTLDbNlY5HaA3P0uN6wA4MwL5GtlcOfQ2JLZ1hHWtwYUgCm4
S13dtw1VzR5aHMasHIVZCGoDum1/Yq7BjtQ2U6dE3+rkAZm5zfR3ZMSsHmm7
LXUbEou9lmbmIeszcdDxjjUOmhSAID2tB8tgIjuuVwVymc1vtjhBc546wpVI
f6GAX80qAbUWFdaBtkiXMfsyYNofY+EnDGu8nbYbXpkXoasdAWXK/Ms9Hqhd
kvd3YixdaIDYaIUeszaVbUPfVB8MwmQT9spFeRgeYxbHff/PLrJE9FBhcGOp
RPMF8NOH2KbgIfpTzirRppvJZN9jHMpc7ki/9RpBCFvJaoKAMGkq6bvPn/7u
pLEdjRFvo4GbezdGkUUrqQWJyEau9rEI30/4U2vxz5XcULbW+PI612NOZY0U
lFCgOaRCqa3WSQ+VwCLkNmMI7mg54nZ5muB1l3WtpC6hFlLohFrrLdJGjE8P
/Fo/B1oXCbcIKFWhX0ilfojiv2wtsNMGxsKo0RwWdKMohXTBl35pXyORavE6
rsmjWJ3sOfXerK1OLcYa+7Fr9neqgI/QwbXJxDmLDveO+ll1oR31T9gRNGGj
M82rP3s0rLYqXIpSwMryrK6AD9Wv/GnLCeJf0I0NQZWbXBd4sQdtTVh7JORU
6g6NekJ54/08WcoB18ehJNjL4NYZODMG4RSYUiqnW3Gy8xdXiZtWNJaGbZga
6B5IRNtLfWneDXnlzpaqTKgzM+NmToNvLnnmo4+OfTiNvA39ca++B4YiosrC
IxdSxG59WjX3p/Ciqk4BdfYDhfwCciQY8dW3R/pZqwWnE0bgeBM1fjwIX9Aa
3F6h39TDeNi0vD0Zh2r+FYRftEvvqqVpDCtycHhGzGO0622uE388TmB7Mj/j
U10FYIAV6ov7XH4QTuxlBhQ9rXFpAIfDRlV9I7AqipQir8OgS9SRY7m46wTS
lhJs9JL3b6pI2kOtJdfRjM1DFeTDF55CHdl4QTaDNsTDcUyHVTq26qVOycse
m8GRwxkz7jKzPiVsjsvNEt4DjQlipkZYEUGwAepl6OmX2d14cfG3vaZ61u3b
UXcAlSJDQqoqQjYYTDTfwBK7b2XNFzR6Vnyk59ydO0f90S2hAbKnF491zk+F
K5PIbtDbfzW7aNhTJNIYRp157e83cy7YM5IpOou+HEehAcm9VIHYHsinW3rJ
9Z15jjOHYx79kLCtkU+i+dWgSeizZgItCTNy942TP5z4EcdWMzoxUctAWKr0
qdrUPRHkPcRYzoXSnTFB+HG9Qt05FP9cMHzPiAxb6lk3XLgO1h4/Y1ROgzCK
rYxF7djd8tVm3vDIaNFBcsizohiyCHt8XH3krDDW8GdZGvS8zkaL2xlYe6OZ
ozSoIiDEQlnpJAYW2rTsettgz/8f/Wh7Tll4X8J+oQEz1XnqNZdLvy8rXfr1
LFqQHtg2dUm84l93sgbqcl8HrM6q0lERCIn75J3K/bQ3ZCItwnPNTbcGRDe4
DnVNoxe57Opkm5PRRejUwdxzq6tZIHopwd1lUNXUPlamHrXu03DT9UZI6prm
SFbZgNjtPPaHnDfSLn5O35k3SREih3ubUHfOcLNax8qUI29CrOnzTiGKawGb
lbBU1GqJP3E8Tvz0QjVv658rkc/QliSgd1CXog7OE0ZX4No0QZWClicjKljZ
yAuL4lmihUuxlO9IPGXewBcY5UAR7FhqqasFAo+0+p2VKkxSRqXyW5dKe+F9
/obJqonGA63qprlvmYMYh9oijx2rRoGunrvgmqaSePWxNBavE6MTUZNuApTy
NdoJ+WChR3zzATxnhE7cjseaFgy7O0WKg8mRRDHb469Ly0R/u76GpQ1cjSz+
3cUqyEXqx91e5jyjoAzfAOdU7lyEmKMUbfHXe0rc3thEiPAnUX0DdCLseXpp
20LWfBZMMGkTmP1PnHI0/q69z4XB6ngWWfGm8Ygr9Dgde/Y64gDb7SCiPCIq
3Z1Fjmmw2oPwNSemUycYQ4sqW4OBh7FLmcuses6MFEM4Sy92ZYRY5Wf2RP8Q
3dq3r1DgiyE2cOb7ZYG78hZZhM19rmV5hICjzEs9OthaqkLi0FYfMAGWYUFd
D3HhGV0zUkiMDwnQnuCZ5GGOPlmGad/qbl8xCEHpEnrUS2YycQ4lKLGgcGGi
iwNUNM2F9PfmHPdN/1jW0JobU7pMXD/3Wp1BZ6iJD/MfdHlLFPvOVWU2gFTZ
H4jLfiy4SoTlxJ6CwJnqtxnXRFu2XDtCd8wenqxr4d9OrLryZEZdR4G0EePD
WhQ77Jxai9iIQwHc5gRh0kJ768Dh3jNfRjbm+chuqY0YJy3ej5A0J7hz/ZUa
LNvgRy0IuK1Bu6tslnNdel1Ayj8LF86E83JylEvOdIPnD6Kz0V0/kooNn9mB
qtopNcRuXiFwJbkRdRqDBUrsiC51LYUAYcHn3vsZY7t/Bwn7XJWjyMWpVbvI
EOwwXTqZdFD96mouVmeolX1MhplOtEi6vaP9/3ROCiLsw2z9QkRApmRJYx6l
7VsQ+++sBmj8GmuIqi/C2Yra0USwTFjSS+c2PIueOdzVkGLyngyUrWtlbfDb
7A3C1FLvkLQBOWHXo9FbV7vpfqWIbehPNq9WQC8usm6B774KZAZonMdCLhkY
CFk2iNVcInCbp8pkS1+tdmCNZtFJ7dKKTf320anm3jWxK+sUgBEwF++9vQUd
kLN+DFrxzcNd+GYuHCtYWSCftRq6UCjrZklQbQhNDh2Q4FcX0Xv7pRWQrMSa
opwOKfSfFJG7AIKg5KQsUydcKj74FypN+mjTIMevCRP67jnESnRvnADS2ViM
o15ux4Vzb2OGokxUgqAA5GZPvbzS+PLnWhpPyt1fM8rBe0GAY/iGNBB8PmJe
RYJb4NqX05rJtFU0Jdvntl249LnHKaoNwpUmxvK9BywE6H8CkebAqdUWr5yf
ZBKyLNNWMklOwXb4ArSUNywSradqwY6xWv47NXTMKevtZiGqWZfUADUnPx9y
+ZTMYD1FWN4DA3Mn7pSIN0tV0WpxlQJ5nVJnjss4oyUaAl06s2CZjwDe2i5c
/j6nuW43LM5QT9MAa6FkItT0/FhP/I/3YnoAtD91wNXVPhG/EFDcq2VSyDg1
kI5IQxjouMNCgrV4G9NNJsLuyXr/e+9Aw25iEhVPLitANBYQoxLeEZiQIFzQ
wJMN4SXiJWtZKe0c7guMxt6H/q9cKsz7cPk36W/poFzsd2L15Gs9YBEoGY2W
xOeNskzVrDR6+nCT4tsTuOQbcLN+eUmIzIUIjiFlfC2Ztk0Z8olgcFbXB+lO
nLjeaIqB1yBPPu24tUIzYRaV6XPFt2oxMbGpDefGcmeN8Oq+pOmcW2TjY6nM
XSti8F/aB/tJvo6SYW20nfL+YHVpFDT/gTod9vf9G78EezmHTsWiX3oBolU5
+9U0opKctKZudIAry8K1WDTOe40wEUPc51Q7HZ0/8qwBLNqKwB4pkXSxI8aW
zrrnk42UChvHPkE/8eD06/7/kG2UC8EYexySNE6QzUZqdERQla2jh86mRHLA
gV/8iu30TItzLdoHKNSwbDVRLkGSWkidpNoX3lE8jIsrK1VkWtKsykBQaDJE
R5IOiMzKbu/KeUP4dNQIMMwrd9zfXmGGzVxNYaKlFtNvk3jh/zAkngUmpx0U
ZILx1Uf3xSedr4ykAkjtnBmMyhAaJdMVQZozFHWff+fcsJfnLTOR2iMxK/QB
u33W8q/WlcHJ+nHy6mzLJBkCMqlF8z8JzGsCCi5ANEorw9RoPilTnYfeuf13
dDnwvatD7m4z34XlxQukDGqpV4ulq3foAqEH2IsYOulLw9zccjyzKZG/uSYL
wAzQfzsVVmkmedOvpoR7u1teoiA36U+YRIyi0oVTsa5PPlfCon9lG/62Icsb
om47na0pa9sXJPDpDVFyi3zDDfwX/DyeiF7WhmWi+Vn3LJrfY92lulWX6wmp
M1SA51PpgJh4GfSLhFWTofakom+4dzpl3e4SWTGnvGWRNv/Pm85S0qaGSCn3
yuBdx1aeug4u5rR+KcXYL+EbchcLH+btVaHylnI++2jLSzIWyeKwH76bU9JJ
y9VHVIR0CjFCLmJIuJIOt+1rg3wzwF4t9+5iHpb/f/SGZUeDj6pTGa8Dq/7R
A+4zTNVMsfTP8XjxptbK6KBoFgnj589JtqK7d4CWst1ZoruIEVvdvqydVL4j
5KW/ByamJYb6TI+RK7pAe/qBaTBacCfT909+Ry7QJL97vyEmEfhq0Adxi7vL
mEGKzJjvjyXBf4JSfPEcWvwGSivcoZ48Va0W5CGhs5R+rgsmt+2jqJl/5C+n
PiSxYXEYlXTTS1Y8yVdfXJrO1vsJ77eCrFIZTsH9cCMObUpqKBFbn3nwBZuL
MMCcS9DhDQ/nlW96Y2+vbZ7hiK83Xi+DXOZ+H5g9iJjphJv0WvNHUBIlLuvC
YIsK4k4bSAQ0mNzsysnoe+h+7b2vYGB1CLHnoVorFLCAthF8FK2S4SfGDB2+
sTUFma3XaObl+TCCUfx6RUl/+MCQ/+Zktf2/rNuWKZAnrb7kIM8qB0H+wBn5
Qtu7rGPIOfV89Lmkl80OHgUTB5EY6oSXhXqBr+5wUJjCzkCbV9At3NVgC6o/
cuZL7WoHwf8zqIQc9iyiAA4rFRXcn7JpYxoXuYTI0j3+d6kPpx1luXrXsoU5
gl5Jrg3OxgszzOaxGFIqJfcDRR0KNYhdUforqS6VoliGP/lIW6pJ0C+RPR2x
sHlpmwBL1m+H4TQc0UaSg2eWTtcb3BK3H+GGenjcfDo386zO8HeYDODduc8c
9MOEq/8LSikRP2VzQc+2SgHV7nIGTK4JBsoP4AS6BzSieQibjXQEr7NAS/5U
yckQS8BfMvUkAZxpMoijEeN/9iUPRtYAvfLi8CWmDbr2whajXbLhKozLYihl
hT8Agd11qNrWwBwDyzYjTzEAHmfb4ZcWptVc973Mv1HFzUjXZuObpC8VdQ0o
UH3YCqTRWQ3SBEy6AIAzhzE6z9jfqO4s+geOP30OEI6cAKD4aeASZ9ljokQZ
ZsNGvGHYkIF7ZMKWnpfTKBApKYCAd+Q59uck45lwrQ24spm8YUqq88fEnU/D
b2s2w7Qhr8xOfvjk0dpLw36Fcd24q2RSldgRW92aD5HhYxAkGmlCLS22+JBi
fslK4hIhSQAn380fNQllHaCbGO6Lb80q2hZNZHpXxwCvM9Qc7Oljpf8NOu83
EhN2b0PHvYm7SxL7Xv8URGHCNJPl4iJ2ZaZDcIoOUV8mH59Ezlf6Qc8g9z5u
V8NOq5Bp8O+LKHZAd/f6OYSxi1dw6Q+CmSnVCWsVdfVJNPKEfTGpcffMdz5n
jJ6pG3oLipZ0+Sjno7zx1aZOKhGjxPpzIa7jjZCWj0zkU0wMYCEXQExRE/Wq
47jyPaq8jqezfrJuYfg5eEA9zlCd7xIvBjm9NDIbvq07XN5frklk+JALj/B9
ISgtGlPAFW/MfI+XYCTFq45Idt8SC8NJ9Auna1bNuuriJopTSzFXYVAgoujS
Md+6b5ElZDGhIPIzz2p8pLTHpf0It5NZEhe4Rez+isWEaj15PQ4lGFIvhH8X
VwTKJV8vUfXWfwXPUYeDYTOsaXbFlnTPKWiWPvqMg33MxwekpC+8hadTmZxk
Sgb2eOA/JNzhoLx15iOE2Z+7+E0DPSX8CGQBrOLsB2603ZlHmAz9izVzx+B7
9/jtq+SvM414O0R4BpyJXxmozAAiXyoDHX4MUnBASN3arOcguyhh9ErOCyk1
sUWMZHmaXwXQMabC46d9DALjFg92TB3qJTziuASXp2ERskdKhydk1ur496L4
qABY6wdIqzJZMw7yI8UWuzOaD6rdsTRT5qgxMXWXgZ71EL/fa76kdw1xVJgG
CzKc32xNF6XM/PM3huoGkcO7kDpRYb/EOMnDeA6fWmar8wnZrm0ZUVt8POtB
iBUGsfuX+Si1tetDXmWryhHB1yj/jiQpR1pzPQmdq3Nmr2pE4bKxGHyeimQK
AbkzH2xSCSlyRF7uOrDSaQ2+5tpL23vS9Kkz3T5QnvPXIS8FbOJ+G6vy240s
dOZtMJyXqqsUuxhHZUpSD33mBdXS8ppFXSMlNeBCLN03shVfIhpdo2TZ3OCJ
5ju1oOVXdRn+vN8HUfWoMoYJxA5Bh6917QTbSSEPn+wnuk1uT7Sempa7E6cb
1EmUzaPWfPrYdvKcbmOrKe5F5DSHQLayxFJbJ7VGAza5BzPkVy4nI58t9adz
DR3XhthJy79Yj0gTGsOC5qub1xhul6cuGkL0ICwI0UVPysPRRC8odwa+LuRs
vv1WHpWuZH9GM5MX2avpqwibLJ5AjSoHmZZuqtdCchzat1Z1Rzjn+49bdMtN
/ljmyyxJvZdYLNIwTP+jz5SOjEndABNjulHE3c/X8gNA6KSRH4wuqNqs2w9U
Ix5FfiKkzzvtZ7Or55dp6E/xsmgVs06V6OAnH4P9hg2mRxucjqNsvF3r5U+7
7x1WxQ4VoJeqK4Ln4LJNCcYIavs67r1aNpmbZzfEcMY6v7dDpRNRWj4R1/ev
eOUHvznHneDBVO4VCO/Kr4yDgDKllqGvNurWQ3SinXBligOn+fcdvLQb5Nkd
ebW2VJz7ImFx5zXCt+IGcu4YfdtfzqstO73Kv1FbtrdvLqBq1f/Q5iCr0NUO
crJy82nfnus1cnQFRmlzShTLnyrNp4pUzYZZ+IY3Y7hlOYMIzEDcUixmiAIg
G7+mj/ae+Uw00YcohJuVdaGlreCbiFfYi3s9OOChLuaj4o/tFP9jkfubnFnC
a24nLUDYCjDYYNVhgDjLyvSs4KnLezcRUIfF3lF9TRHdI/ddierMC5XeQkEL
MxeATsJso9kJWQFyq8JRZNFJ7+A3XkwtLledWcAJhg70vLccSjpvTTaRK3CH
XH/NN/vZAb0K6T3de18CNgjbhTmk5XijFo9ftQ7Uf97zTfILG08mw3PZtQ+A
K6gGDzofw9GTh13gg/mNCWBSmRmwG2CjG583IIFaEQ4WduyDHKzvrt/bo09g
6OCKPAC7M2S93i6ys/odvSXFLgZPGlqi2+DXhrWwrlEPhvAb7aYBpoF+Zw7J
fvf3JbqY9jGU5vJFZuidcK+niJX6CAGla910OYjBruoxe2Uzp7zTOSyqJlIN
jbsptvLODDNpzK5m+TAVpHCM6TwluNTsv6r5nBO8fzIdXIqilVHQXF60EY5d
E7RQO27E1a/+qGJk3vp7Iswa0/V8t6H1rHSaWs+o8IL1tGrP70JyWoEJGJrq
jNDWCOM3hX6yofHM9PRyC4RxJg5rTdss+5opXBV0V9a6PRvJzEDHnwuNRhrx
lXQ/EvPwae/ZRRYV8OVcrOvMO2lWhb06WDi/MkoqXcGFu/yvYnyZpmyqdU/J
mhsNAc5naGbRIupazTZqPnilcDj7bB5OWN5f+YFr9C0rIaJ07WUafRb7x2MA
SSpsHQPhR0fZyrhqfZp8ezEdZXuMete8EgphUMevZbngoYU8pVwCYOaywIuu
Nj3B5xDQnCG8wYECIuHXFe8TnOu2WYP5Dyws16RZxY8icgMzS6dvZkaENBol
hPArWZ24D1Wv9uLwZ/yW4ZITgwsvVqPkY9ngq9URW5UrYPdGbb2wUk/qpCqk
8PVgNEASu8ACf98vJsGzG3s1jySjOyueu8WBlvMMR8ogQbvcifBhiotD1+i3
ij+ZLA5mqowyMnSJwLwfs9oBeCevEhMGz/oPZRvWOEMKMP1C2bIo1lgQ/lap
nODiba+sjXId2GpNksgoCvf0fjHzShmM4FAG2AXJ9ni5PxoedFc+sYdhh8uZ
fhGQF2wJaXTkTwlOoGu7C9P0N33VaDTMDXqhbiqTzLPM3ta8U2DKZfFnBB64
vQ10ei2yGguCNVgvaG5CAphhKNZKDC+tJZtqApgYMUTqYfj+Agy22HckiHxQ
PpPAC7TTi0wy4U2/huyH+1lKbmWqttL5YWGtkAiVz0LpwT6y00puSa/DLGA/
q96feUb9XlsfoTqiGAOZpp/ehiC2X90t0FumnLQMIEyzKbOhVhQ3uAg6mnZl
j+2/AJiYVJrXFI1pkboc4nLbcNxlq7zmj/b8YMcZHrHZgvhGfQNnh2E+xGv2
2pU1/2bXOnS7LGJ0uFdeukhyWtGVUsmqj+GtOoyYop179Eoiuuwi5OmbEhSJ
OJA7oe18Vlwpdpq2j6jVCgYK4+qP/f/ak1oGDl+CXnb+xWf7n/awrxk/zfXq
MUnIwGRYnz1brnW+5VYJhYxsTYGf2TrQqe+zEZy0mg4GsnfWdid/5rUihxHo
DEMK9rVscXX8c4PyhKnznAmpO/6y1SxA7VAh414pRaiMXYNKOQdAo0mneAhs
zg3lKcIB+WMN0ocuB/BkkoFzRSEX2dQyXJqcBjejwVBkO4uSdZ6aWigHAo0L
hCrP5zSE1qYDc3DmPpNl38rG7vy5rbAXad+UFOk70gQ5HPpoXvSMNWIjrFLn
VCEV+2aZ5WZL0VGMgLlISmdp6uA8v8ErI/9BdQUVKQU+V6meXZhz2/YNKxoB
6dOn29kBNCjL4DKGE1I9oS4SjQrmslV4juvOLvzpY70ksyPS+qJmgRzbtzBw
wRp3AVYj2ESZxFnOmdxYmas1hv31Vu6ySlcxOzElZ1EVCpHA+Qxd23FpFlND
W6t4frJzH0FXCiB8BNOdic9NKpg1O6jLHspzSpoAiAI43S40OORGPJj+pBBD
6KQRNrOCkoCDSzCnyYukdfphQ07LbjPYN6ClMYPkyvog5+wdqhciDs4vTIts
rUHUFHf0faa3Htj3Safb++XHg2HgzxCJKz2o383JfMj1qeYZbqTeIu4OHe6v
PjhRL3XDGDrqsphMls8kE2RSEKony6+FGiY6t2e0hrWhEjMVQQJfpgmqSSsY
Mc2ioij7zi3R1y8daNGXDckAJiJJM+PtGxLYvvrkboD6wZWM7oAXnvXksq9O
4y5sdG9ROft+g/eXXXdsOIoGFnFxnKG9hp+pbPY32HVU97JrJDXYDlp2Qqew
2FIXNEAVQC+p98EmW2nTwJF106VXtOJNlfyd3mqb2MeXZbTSRV5yzVt1GzNq
r2GYK40nBGq6JmeVscrIt6zODfnci2eXSHVSww3oGFRQMRG9iUTCfn+EWkeG
0l+t3IjRTloPjvrdyHS0jFduQAWacj7DqGVhIVhuNzsI5r9EU1VVLyAKuaxU
2lIBMgLI7d3ZjtzZFh3ouH0hyZZVbjelMXovbg4JviYaLusEGy6lUu19WD8S
4e98Ab/8DM9+tcTOhd30LY52J4lDNUJU4d8IM2n9PpK+gCOCF0mA71BKkUBL
r2rQHwlksEwZInm2kHTFMcW8Vk+9s8Ul4E+Ov9DZGJrMIem6I0GdvXUYuFTG
xMQSDUWMpprj0X3F7j4UfYtmELWy1jv885FvY+X1IydhzYYqCdvymPp4Fl7Y
QweOjdo7FIQkbTJ9IKadwb3umr3KtMGXl4vR5BgAQA5FAT9gjT0HZuoY6WIZ
RzLsG1VOHV5gbhinIFdmq2wZKafieNgKpWCq6wCaJB44J9LOCEeeMgMi/7oo
OfLzwCDXJj2GfHmKuyQJi4HNo4Y2uSNvxCJy3eSlgA7Ra3F1R2pVZpOKk4lJ
DhTxiMkRvIR+Ji7KDHEc8ghJgPI1U0YbkqDlADPPA0pwzo6Hsu2zhlhlGc9R
OrsGlvssDOAplJDdpq+8YAwpNbp7HiOd8twnV4rFVyARD1MO0iWKNkcWLSwe
6c7SyfHmP+qMDDx41M/uFKcXPODPk198HCO+4rsuPHwT9Esc4/Tvgw4AXhA6
X3qojBd7USTQ5hYjcFBTUmPtcRwuiQsGJ9S7nWqsNuHwIXwmg4115LQsFV9h
++B88H4hwRcPw/nwd1y4ttXhYweQA/MgCwLAPS+t16V3uxvw3TgdIzlHIEQl
wwlaaO99Cw1ruCdjcC8tM9kcm1jjyNvRXKZfJ137mE4La9HbS6NJGX6H9UAK
4/ObQUQHBVanHmfzcz2JrszacGPT7rPGLavh93+zksGFlZmL7LNvqMWkDmjb
Vs34xA6FkuFMD71syh5hTcBSTddX0dL6eYFgpeA/xih/B7ipNJYyncCOkXYi
SO8bsRWnGCHEgM32Ju7fIClckedxjty6MhQL3khA3xV9NlY/1cBjX/Iunfab
NJ+sYNUeYdrBEY1QbZjzAJv0k4MQE5n9lkUKK+RRjhlN5oDOGY/TjzK+yxJa
I83M2Iyq6kUJkVTs6YoMyMiiBi3JYowxWNCZyelgRIAECDKbMXbMSA0LNfN1
EI04bPLRmMhnZ42ANVKzc9+1nKhIhTekUeEMgkceA73e6MZ0B6YGllNSkQfi
IVy5trDFwtzdCwl4P/ZmklWPIDPBGe2ALY+YIX60CJdELyx1C3JzcTmdSSGc
k8O8qmF3w17lo8+bs/T6TI/GGDhaQYvtv7p0QnIiG4Vy8rnqH/4lP3zMWtYg
hbORzSqivlrSeiVCTjqd6xvDeuXSxsct3uaUcqy9cXF32HwwOzm/L6jB4VoV
NYH/B/+ruY/BLz9XJ+6+ZuBP25bMpr2UR4uK5PgxC6y+8RFm2DEupFU+K3Sw
G/gFSbXHJFz7Qixd0lWPOyXL30SqPQrguSPNkxyaMCCgvJZXa8UmEeKM4h8K
z88uFa2lxlF/Vdvjga/iyRY75kFc/dQ3jlrSZ5ZZb9R9V07cQFJXW0fZeL3N
RTzYQC0P0QAL6UNmRsJoF0Z+lSusSYY+Bglkuhj/q8DLEqbrgx8Th0P01M8c
Wn9xSRyFylX641EBNIKfZ7YW7zm0bgOi//AkiWvqTk7pysNsH8cReXnfjw/M
B3CULcldY4+faO93utgbNLMcYKmHNS5I8WKoWyRipaNZ5VNVdNhqlfKTgKBc
GSYWrwy2+gEScYltsvqBdJLbhSdfow0YYSA1NtkgluCd5Jd2KhO9kcUDjt0J
60Scft29llT2tv3fKvhCiSxiX7uYgDJtyhB83CxY2x3jADKoo7cbdIB/A10/
8/ZGRWhSW+TFbXrNZkEjDTKpr1N5mTkraztUiGiq5hPBEzhwTZuwIO2fG1QN
99YKOF90XzeHHytIBH/FaHz9oIgXdK2NFFd/muXhamDqHJ3rTh7RtTsNFq+P
zNQFFJ2oauQWTnToqqgyXBsMbCAAmkfpAQtTDfnu7aVwf2X7GksR6+wrtsSs
WmKqdhuk2KQPg/DZmRIH+Blj956TXNFt3yPJTcGxzHwaGnqT/dnFfb8W741y
fFBgFuYnVmmC16tPnDqMo+mFdhfKN72ammANAgzBLTA/uIeLJzPWobrUDLKN
JhMl1LqEIk0BiPiGUEIdk/eKUaF39F1srskM5xX33bYgGAkUVPlc3MWSUziS
/ycbLy1qQV6lCDLs7ZM9kZL4VA0PCxmYAcVDL+cgb2cFR/WYgvU9f33gBt1h
WIRf325LdZPEZRsGj56IoYsXSj1Bx12N9w04jkToltnm3/1s+uMETZoW8wXy
0mRR6thKs99tyhM3VkO/h3sQyVq/lJyui2zmyYBCA/6c5fyg2QL0om4pdnCd
INm7FtiIvxUJk5d7we3Mh9Z+nvpTxH9r+gPtdlQsPLg3K6EfUh162XgVqgIi
9mAC8YXZlScXZoszmkHr/3GVXo1TSzx6XbW3+IiBH/7o5RBzblKsynw1sB30
VHdRJF3IeIf0s9WsRjw09+ebuA9qyF/EG9zPOpNaP2chqGOIKOVRuDV3Ghe9
QbopDvNIJcuRXLD9HaXeLrETFNeAzrhXkYonxpp1iy+eqRUgrlGEhMuhr0Rb
nICaLCSwzg6xl+YXux1o5fnivpty+DuPKIhB7+RkLx2JYe/rBaaiof+DVxnR
IA5irmRo2lmb6YRWs24XaYiWW1FPmmSpBQG029ZisPCK/fNyrNXSoTVmvs7l
PXMIKXzWiFb5CVX/uTDQBDd9CypeR3Rb/pc3pFXp3XkqQV6Lhvl/2mqIVoDV
hqGGZaMzaBQ84YoRrNrjhVBfoTeYXe+BiVcvBwmlrVwfn037yEcDH5wwAEvY
FBgBfH71kKsNBajWG8/1ZTMOn1MvE/zDeoEA211XePj505jQf9+HhYAAIKll
1pKzeyqKVKacD1CNvz41T/k2GSEcS0Jj3sbBxVIJ0Aq/ULtWBhm3au1hEjdy
HdSFt5F04Bt1qjTgg+aDBdTQDhWjheiRWuyQCAEU3b1R22PFKiCWRmTRU6SE
98uKlbq49oa4nf9JGCJI0vDhj/xORZo/rRTdTNEDCi2XCEXml+qDg/wDuegT
CayRIH/wxcjZxV/ck4xFkYEMNyrzQRL/rGZ6MkG5clqYxnlGd2YCXA0TvrhA
sJlGr4YaFxRbqWXh4Ii1hxI0oolY/BALQZNaGBL0xZt/qn31qR+FSbv5101H
SMZ0pn9AMdpisYW/HnJCiU880dga2KBuilVIfyU3uy+a80FF5788sF5oD/EH
AfapJfkl0lsPtAibbMYr7qPHql0yU8QldAJuqaGkKlGMLNlS8iE0I7CL4KRi
bkwKCI3xAKEit6AEtXJfZNfYJtClgo6p/BawEQEeCdPOcjUajSyS9NA4vCwT
6QzvyZLZeg6G4SeYGPSzsNNruTwa2MCkMwZpoZDgJvCeG2GPjmPp2o4TT4Sz
dRtac5IjFWblphYx/Bs39IaXzV+8T38Rz36MzEBzsF4UN4nEZv2Kp7HuZLOf
bZm3n0pT3f8Ej5ECXFIxqXe2Pf45wVtrAgawreUk2y0feXEzR1iIlq3BaiBb
dNjznhWfhdvnKD7UvQl6ZZIytntkAgFYjMMmq2Z2yhg1j3m80sS7k99YtgmN
zn7vbgGPtAclQ0ss/nT1Q1Xv22ppAFAavNU/HwV1BZYpRDIxxL/ImoHd4aYL
SFzxbD8Lj5zTcIi5xa8ORQzef3uYBREEmrw2J7gI2yf/OF64FRUGcYmY/tpF
dcRcn67515h58BlWKhtHaNZIX2pN2RIYkIunW8yvHolmFmeKwZwW1hNR6WsX
5rMrWLHcPxMl98b5SPnb0LiyuEkD76k4Ucqzq7HBkDJ2Njp0Ni61K+0QrPMz
2d7ssm8cRGzpEIHZQtX3IcrQLVIq3SA8aDWlFd/0akQhMijX3CtJ1yMGdCMJ
K3AaTKScUZPTIKmxuJl/BXYqJ4QGa5sL+75SLG0wRPYeml3Z98tmEX255FQO
karCT42q02SgXqDgvD5PBgyfKorb4OSigVSYeScuFsYPwmmt2tPVz+DAQgfN
tHq6mSBMG/r2u6He/cYfOMZMHWPrfypeICibfLGRcOrNH+sVNjzkoBdtsMMF
zJ4MHkQSLr12nxrhqRRdBYNlVRS5GkXqIbzc6EYohYEo303+mr0O+5t0pYUB
J9ohJkLrOlmRgcu9ewyPnLpkpWMPSaZWClbajXqQghVb+hleGa9bE/MuqYVI
oMlYSy6sq0sjnA+KcBS/qY2w9H3c1tfzhfkeN/w/qUJ7NkFHY2pvWqYkm1ed
w515omlmCnCOSlWX91zrHJ+EXxwEpnO0Yb+egUrOXqQon3iAhXQGElkS21IE
6Z1jbJyFzQxnLtGsNys6YKfNOTsAAsEXuMYanHiSVH4fuS7f8UgGe8l6L0Uo
MxAA5hgimDx3uQY5bgZ0llNi5v5nPpyNhJBJNxEstdtiwnFvJtEj19s6gUpn
BMo6FGdZ8kyXlp3Ds5cY/6zQtpfX+JIHnwj7rbDxcPEjxa13E9pyS+tLDPTj
PwZ6jkV0XvL0c7qLOedVjK9g7an/wY4Y4Am+gqSXGKBgtcSU5/lsN9neEcfk
VocalVmwZFL0mR4ZgyzuhpOF0AYWCXiYD2MIehVtLFB5iWn5PZAHoJb8ure7
5hTKaJUvpKxgEaxsT3zxEhKY+rO/OQrzcHm3JvQLBDTowZFb5/3wGyIK4w22
hzJBPIW1dnbci/wc5UzHR+uQaad6N9IrdPvil078kFV+R/JftBJK28q9JB/C
Zjhg0m5Lkw3as63CvVDYEMMPIfwpkhnvVtp2cHrbz1bJUbIOu9l65Vhdxx3x
bTjtO8/Jk3OM+4swkXY0ExaCIMTww9WreFJS0Tb/MLkpZSfwsFKDQGmeHcFI
35QRMeIbqcN+hBgMVJ2mvM/2kPlOeaElMhCF/OZfhDfHsj0/kpSHUqzwIgyt
yWWFiG1lp1drokQYof24e/9IAb/yq6nejLhYoo6LfABGcNIWWcgG3bP8Y2AN
p/R81b646AGAw8FhYCsgVh/h8MPfpW1ci9wYv3a5+55L4oGVXOVbhTT29uhC
GB0na1/DaWyxqozZFSFOrWZ8HRdkJZUbscmB1SAjHPC6HOclwboQiw/Tl83n
rDL7RJNQ4yYNI8YQB7nOoODOGBnM4FkhDPHthiL7+ASRVnGUddm7R3hm5hxU
GGnGTE+p4fIZ8QJ2JyQy/jFX7+bTuwPOCYbe/oeZ+w2jah6XfrrUBBjhXQA4
8HkPuWA+idyCbWus/nO2I3ZYfv6xikczZ80rLpFfYt78DGb+v2ILTJJJuTXG
SHBA9oyeklqGoaJDfAeXnAnEADbh5IdORqBHBqveIovRbT11u96wrKnscx+X
Kui9SuchVlOss66/joWuG62N9T9feCj80aT9fn0DYAqwBjRs67sMIULeG9MH
N1o1J7QbiuQfFZ8wxSbuq7YNuNcsqE6f5IfYBPmpPUTLpwYQ4l9JWcgowatQ
IJd9ieXdBNwTGCfVCOOSxsflocUhazODri6/GVU5MhLxuO3jm47ZD/+30LhG
MPHfH2FdNfYkzc5hoxIudYWOyHkJyJ3uMtpO1vEo6ub9tQEO1yJeBkhpFRPI
vPWrzCJbwe07Xc6RtPnlYYCTTF+Z/YgYw7E/LDglr/txYd+BESBQFGDv8Iup
2bDMcmwBcGdY8D4QmNhTSApyg/X7OZUgtpblEsKeddZ5EvnV02Lcl87ILsLa
iVkAp4Qvch5f9f7tYz7+MNmdnkmtzmGus7CopQ00QseOh+gZyVm+LzT0UiRv
LF+nrW8ylqtgPDCDRzEjy6XHz+wpBOgMxHmc6DT2MEOpVebu1GsVBNFCZhnB
FElkytsfNZPNR7lsumLajbrptSZlAyMDU1kSCdOMpiskSOroDvP5gfTwXEZL
HbCZ3yNQkWGek0LzkSpXWnGezhbk215iYvvW4axUHJUHsuZpkGNiIY6YHw/G
75hOhnDiMWvpTWZ+QmB3gODmPqFb71Rk0vA40pU1ntWRhhd8sg3LQ5+wizgL
c/rC2Qt0cxpLCwkTbaZZwLHmkSfOZmNXbLf0lrHdHzmPMn0S/2TXJU5PXWJc
+fGdzG37wij7WXHhPXrby9MeT2og+dyw1BJKStNyEvUyxCZ3X17HGVuhH4YR
QbmEgY09gOg3/Wwby/p8FsfAv9FplOzgKzFJ/kp4EGtYUrJeUUEQrucIYYEP
eVMHuwpMK4p0LDNPJMJl+lIyXqmnU1OlpO6778OYOFFFBCgu6XiTh31Ysjlo
GWMRu0XxIaPYZxy2qaM81d/ioJKyILobkE8DhNgMncoJNps8l9FM0NIlvc/z
jX/dn6rpQMKMLKaPzFRQRU3UqFsUm71HcA01RylZ8lFSo3VAG9Y0f+Y23VSc
WKm2fch2RVQPDUhy8wJ5Od4440gV+KFndxYAXtQUvLlU1FUevsYirxWsqjOf
MhIMtBx7Oa7B5oH87T3aoeYBNQiCoPrEFZ5qJ5W/TcsQ/c3pDQ85johLHMXF
MlBPJ2FGF7l66hrIZFl63x+y7IvDWXNFChDkD0iQbOdy54L8aFkdaMxVLa+v
L1n2NE56yxMN7ixdiLUAD5wr//58rrTQ20J/zVF42TzrQqJHK7RfFdK9PrFi
JPEkMcwl6COi772jC5xfpO7xcY5HZrYWIC1FsYuCRJ+Hyy+B7hw7japGSBDf
8NMFf5m51dY7mJhYrFlvz26O6uqMPrc+n+jnaN3HiVk6xu+zt1GY4SyNrOIl
10gzUj5Fe3STMsP/c8hx74DKeCzLneNjDwTIZNKh5LVcNky1ptYXA2bvdqD9
rz75apObP0iBN/B3De/QeystTaMszjQcPDgVtLTZodB1C3Ty6Mhspa1JWp42
M2gptwQgassGaCG9xGN5wTxplTsEmZQUPuAj7FLb45R7BCNFSzs7UctFt/BI
JzDxSdklh3TU1n3I9aF31rtPvSu0NCI9yfzguP7WTjVUdgzMdDvW1ifbKEm1
WFkNAwjMHdBUxZkWGM0G6WYrgp6kILvrZqPCFGeyt6ch3SfRl2szsyum6pB9
DqBzbj/g5XBbTDvl+4qpgmpbfrUjKwNs2NAQNZEnG4JDZ31CnFqCe8VjVBju
bE4e5DQ7tmwYy43dW7PgZnQyUcbZ3oABvV1gUQiY/wJDQY0QikKP9dljXktd
bJacLLREaFkKbMNRqO2Yu3ExS3hVZPkeRhaooIwNFyaVpzQljQcdeIqh0EkB
qq1zTbpMi5UPsZEt1iX/vwYCdbD1B4Tx7WJBgBm/4dgf8zuHKhyVK3grYpQA
72P8ckRnljNVNO8D/6GVm707fb4KaidUD2HNRuWobqatMz1bd38mEPkhcstL
Y04TA3601fu/auJgXjG5GiQ/EM6hwWZy06dq8FRzyBc6Ra4gKo+c72Sbgvip
JTIag+0gprzHgr6L39YxiNxrgmap1sHGIVeMNYIjZqWc7fW9i6f1u8LeuFnW
RgDFDPUuTbHr5UloXtqYrtxJb4BFaUIjAurDoSWXdMqAK/vyf01T7POOo5up
1S/mBa4V80ZVjhKnZuxGnzH36DirN/lkfVFBe27JhjgaCy97/p534G5jF1hq
9YupmwG2r4G2uMhIrJZ7KofJwg82dCy5CvIh0nPB/LQUZpU6An/EKoxSS6sW
yU+Mco68/9/rYZTqlYlSKsogvl0m3R1U0kbEO5PjJGYBTVqv2VxbsOPhswqc
ZDM0xqjUF/v4dvwew4vuOA6FZIDZEfnF5H9tQaamtZSCKMgwExV3+kWRkxri
kfO1lE8y0DaU11RjUbC/95Um0GYHPFEgUMpqlJ3wgnOFrt6aFT8ADQh1U0y0
gzD53Z7rkM3qX4ZFAA5xzB85YqBPQ45MN1g7DPAQGUhGgz/itcyVTCUNFThs
ldum4w6KxcaQl9RLyPN5GhhV4lzsOTaASP1Gc0c5HmYPMuJZlbJ0HIFA7a5i
xY6Kja9TwObrlDWSFYM0vYh6rteCmDx4SIAXrRr7VqE5uTVjfiTUl230utMO
aOcg/NxE35Nm2AIG69w2Jlpfl2mw2jvJ6TvJIhcZ0fDb3rjH3P2E2bLqdes7
yvIiqMluHMu9M91Ynq9edrXg16cir4HoGef+GfwqZ6385DrTGWePv/A8MvfH
R3hdhWgdwNdFar3HBuPKQo5hy9yIHSQlLtvqC6uTeuDaio47bz2kSuX+aKXW
2d+TXrsMaNnO/nEIg04LNAYShIrUwHaIOnUg1BsBLH1lAJA8MMCBmQo/lSHE
utUtEVjZ5OQ3BqtznU1Mwig6lKPUPp/mq9iuP9yKnIMbnwl7SGi2kVMJ92Sm
+WSxsg2byo8kE2VGZ00uNd1qp4FYMGRBQHV0pFvGPwkVP3fq+6R33glqQped
jKnASeYVnmb7qabK4BCua5/7GG51Rq9/yTZGBFxOPiFsM4ESAfjUazdrP48b
nZcWgpd5eQoGVP5hVeRs22tUSM91kyaSTKK9MH5k3jpzZJ8Tl2RMKan3BBPr
CBrRXTJcL20vT2O3D4a58eQJDh+khOkdO61H72pNn7IG+g2qppkV2I8DendC
4GSwxZct3eMicbU1FUFWq+hjz8j0Z0iK2xXVSq8ME2eSSTkAJP0kLT9Wr7Jc
wyUj+RchiN5IL9FIbAe/SkuZTGVi++8J3RLCXeEF5wi4PR9Akdp9/0FNWIKq
1vdkTqHEdfilLchopJ8VSy+PdfBVw4is3VJXs6MoPadr0Fbn0DGD4DtQZ7wC
xgt58GEJdFMTbmRa7yUhSPNFlnx8z7uIZ2o0Vale70MxeT8W6fNYpip+XSpn
HKiKIVA+IMN52QbgWiyTaNw6slz/8qAAR8Q38sCddngQg3QUHy5an69lJ3uw
y+libtJLAtJESGsqDg/OBBTpsZMjXqztSgphZcVT0dVeQp4zDS0oQSfNWAlk
f9AfDxk+5pBcnTMPXnGPNz9RFdDN3t8U9rMRv4v3iKeO9vaEYxk2gboPtAL2
En5ViTskHDdygoK/HmGOzHXq1gwcPJOxVde8C1jPQ2K9SUIAtDE5F2J8vYuh
YnsOpDdMsK8lxI6ziRRrZ8uRxNyVwPtU6PaRLLG9mbou1I0F6jaauk/0pyPc
aVNtCrfCwdO4LC1vN3XqjYNTRIx9Gji0ZPH819m6GtI2g2y0vvL4Tr5RoYCx
8iTaYQcJXLym9ZVQRvb3wozYffkCYMB8/j39EQdxOBFxlHA47FpMAccVmVG1
7qzvAEG/XUxjMibKIOz2Ne88ubUBe85Blht8bmzKlo5z86lqDHIlFIu2rmje
GNKtuC77/aJ2lyk17DrJmVOWEExSajIkH7uhVEcyMk9pZlI2e26Y2hn74VWZ
NHndeiXTe1C6L9ln9ZaJADiSkcDUJ8UU2HxDAifpuozQLXeQbcd8dN4C0O/5
DZ9faDMKbraigYKfcBCvoXOrJoWaAacD3xb69eC0xhrS8wSyUTPnalRNl0yF
NAWx+IogFWFkG+aUPGgOQZG8FlS/p3jeZsc1LU8c5emvSWD8ewEkRy5cwLBo
mFoG9mW7K/ZuuUJ7Kb+cR1t4c6EuoH8xixLpo49BJRKaDR6PALdd6rymy2m5
jyG9/+zKWi6X4F43aoeMlqb5+TUFPwAa/eopyb4ImEtgJCSR4pNM+M/v5tgr
GFLu2Sa4uZRnfgfDSyh63NT5S1vR/NnYGFRIBWNaS6Xizv3cJV2pUkX6UB3B
rqKTXjCHgonntSqoo+SKLxWEs/z8fu3Pemx6ncoHL+NBT3AiYtyWFhtczaM9
+CNaYiUZoEsXIec/Ta0/L+fnPzoAJKsfG+KIKic8IFdyRb0/mrIA4aRw0VS6
n8e9K23F6AF8DkWW0r0qY9zZVIaOByYc8Pr5/hxuxn9PxUr7lb0x4I6dyGjY
H9AeNIN+XpQPzRjd6CnBPBs1Eeg55Gzt2kPpTiACYj3c8d/RBvxLbJLt579m
e/mpsGUQgZH+Jp8CIGSku+Ghox5ANN3lzRl+eUP6bSfNW9GIxRNS0j86vCsD
efseOjnckbHYorKiTTsC8VhD0CSDUpgymKhUmh/yceMXpWan/5hoPinJICNi
WNGsieUfwz71rb53zcm6gg84NA7tV7zOOYJD/5HVEgR9/6FlfnEdvKouYbO1
mDy4GA5LjlxaCIivV4EmryXZCo2lHQ7gTdG39O4/wPWiAw0zuyVUzI6OiHeP
ao5esYYu+mioGLzsQmVV0XcnlQhIArdE+42/9B98ekNVpu5sXPfqMADXX8xp
NsMIMK5+w0glYFXqdjynavBuhXduU6hXGUv8C3PQ/qCp6AsDebcWeqdj6kq2
Y06c9hZBukKnCXG8rIe48OpasOr+AkA+BwpQbqtecYHTUI9dRxoGXjdiPQUq
pwKH2/kd4zvHnZd6RA1FsAsXp57MRn9zDBO5rq6aO3ofTM7RCHNT/Xdel73t
NyrrEIjXh5XK6t8QFuTsm5Owt9MM/LvcK2saDWT4SN7GvHMnB6RQ3HhZTa93
d/sThZ1IUccAc0hzBG0W26sRGqmlXt0iU81kcLGrigGFGO9Inux4PH5n/iep
KJOOmKzYw1hPZq94hBWa1CZygQ6O2Zte6kxnQ6F6U0RzySPPsSH5Nrsp2cn0
fABzH4czomVJyvJNxldmgIygKO144HUWgIXM8OTgN9s/aaB7sfbEg59i7eu/
oczth5Q66WJ7FagTNkqDiVDrturSeh6MNxTWxv4w9eFcHmc0pQBj9vW5rMMV
+birowEKsDfM3ZQWwv3kGL1ID8lnoC4KfeFH6xQlikMHSzDbgO/ab3O7+48A
OfjZv4JWgiUfasY6voCJv4itqkLZVDKrS154joY70TUPrWeefMFqalxYEBmM
uVatC/X8vS0aB39IuYjAt2Ny8R2u5T8nD+beHDoAlk7Fr/hLhyJjUE3go8lm
S0KYV2DLPgQjNY2MpBitPTHtrIQ2FORoQPjr8rTSvslpyADiJ0uAwNMJe0Ry
IUJUm0i+bsSE2Wda8I52GNP/oarQVSafrcBkT9Z9BwuPJVecDytk89fumUrs
V787XK8/0EPD6FTidwYsvcB+hXJDZep5ZvBhX7HmMJejPrPOAHMG/umAjylM
uHieLJlMjFjtjerDaeXuNJ0PUvlb0ZFPKM1dkR1WfGqpDC2gmsaUBGQpffrJ
4F2gGTIHGcilbpe6HARW1aEf77ReX0lyfC0Uc0Pvg/y7nadgEgWh9V7lL//9
uEU8eLw1botiS5H9H56lJXVdXctUQVCpQpphvUVleqRkIt2pcdMAYKv83EOJ
8TeL9zHBNqIJTXkDHSMGu7ddI7Tc5LC9Yb+BkRdUCLgEsf2NaNXjAbws1sqn
jtti4HUgJyzAVkIowdcpfq7+8epJMGy3l7DhUw0feZc7HrnS4+ope9jCGcem
3LRwnyU6gtwOmzRTPhT7gHkBm36wNXeGhriECz/Ooi6ogeqoluFkqhn7WYCf
pG77TsQkgjD0NpEc9bAXAQFazYnPhkzlDpEYhTCMPUZK1urWwY38cBS9jMpx
BXzPvbTGjxyQyOv9je5fKi14EJogSE66H7mPt4m0JNm6SuTMdboTMHThPv3J
Q4c6xyiuo7tY3qT+0Q+tNwkgruh9VpL8RMWTugk6IuwSo/oXyFKE1bb39KxT
qJv7THk85M9AN1GW/mBiXlnHZSvl1CnIiZeNA0X1UtJKj6Rf423ytmW+2BC9
J4T4LY7My31ZhTK+Klh6COZzwBEu4PkWHbBwA5fQjOhRZ2CuwwAmKgPk8AZ9
S0JMsJ7F6xQQL8eQkdyQC3CD3aTJcqVfwO+tcH+RuEd2dz/NqWyjtXnkEu4+
fCh50skQFW5B4hc8ByR05i74IT3eQCzDnRyp7ld4EQMWzZMzibGxBGyNhpgr
pwJ9kBes4Mj+2zXNdRY6jXkuU3JqUsvwH98+ILla9mjLCJtueRLfKpfv++ka
p+/4WbN0dk/W/5XxtxWiAUroCSeUuyDkZYY10arCHgbQQSCTwceBnkqQjrLX
WQMtO/T0vdktQCRSIJynbnEysLD3DrJPJ9u2AUvZXC81VD8OMtM23WovS2oD
pOi6gOiWIR3sW5VdAXu31d6Kz1hsN3X+dgohbxdwmY9nFUu9u1WFu25thhOz
njSyYFZr6Exnu1C+kiUWm5H18AxJD4zJaw+0AHDwITvKlYulAG737kJB2Tox
JrIASFBWe+WbPMJauVT5WcfRlr7aBBkVHC18tGcBIj6P+m0gY5sOs/OQjJOA
/ZwSfo8ZU6Rr4aorDNm0p/i/tVebOrVqkSSTUT/1mv3RJsw2AjHWZyhGjIiY
tvqw5QpuC6raTw4cShu6CXOA1QIJy9w+b65F69ID+Jdh9atdIJpc17hJYHOv
I+uRP25XgBK+VOke/PjiC45YjDKlfjVyumz0nRJF56OgLD8DMQ89LRzc4rsj
COf41ej+jLiqkgpwFF8eGaYzLLYiMozvzlgsI9ywLmzXtyzxEf0By2xihcHS
6B/tHYelg3in3WA51J/6WYrQ2F3Qyug8vywmJkie9TpGpf0aREcLXxTk0c0B
GmXaLW/aQ7VBjJ/DVOdA4ARDucYyQVt6bNervd/DMQGliHXjQ41UAVxRWMhd
+fy4VQV1z3f+67g4eJ+GrhC544B5U8wzteTorpNwtYZzKZhXZ4wSZqFmcEsR
1ptz3N7wfAIEDfp4m8o1U2KRuQ7Ybc0imbBPxgQbFniGCGZwICTDxzisXaBt
kQIjcRCH6nCGXGZcS1qrA72UHnfcMHJgHibSlZGM6Imen6aIRUaaHOY8Ewa1
vJ9pHaOUrjYfx7cm5Xi5oD3rZfCRabZniW8fwRVNw6FSOqV80lVgNDiyI+iZ
OyfpXi9bypR2N/i7fg/ECSUNuVVMX8U35eiCzv+4LKF8k8PFZXVNHZ5cWZ/g
3FfSKUZaX/10X+QJ0zN+Gt/mtXPkr1/hedPLDZbTN+lo0+2wMFo2KBpwydzE
+Bbplxp6R74d5ewkMKR4WHmn1WCnNOI2zIBj7zSTOX/4GGAUF7xt/XxAfFTo
tQLhaSAJcPSp8V1yB8p0+CWBSBLz4YC8pK2Pw7ndOnogMCOP69cmO08LBaTQ
i1X59I+xF1/Ho/6bSVu0SWBV9jhue+c2yTmuEZwhc67Rrs5NJa9b7Vgsj5UA
HQFtsu5fNU1W0ED8VM5RPun5yLTqWu4kYyZtOTV5Kw0M77BeSQ8Y8by2uHtL
6p0ra4TvyFFVBh5WYBJizNPVyhWKm3fHAUGGrf28wwGENpZLchWOTB8HyAX4
c9mkGNXuazS+BLRsekbCLNMqK2p85qRfDmhjlpsogKtXELb4nOS+2fEVAUaL
4LkSEInLeKWmIvAUGONYXIv5O0zLExV4DbJYjvYR5JNX5PaVGFkd6kQ2y2pl
pshleW1u6prz1LfqZZ/71ZzK1reVVmN7YF5uT6AV4i6sZSOY3gpbhkoDkmZ+
Ac4pRGpqu9NEzBq4sApsXlLyDwL7IrY1Mn6Le142kbfHnIVSAbLzSsSKdt2k
97l+jOrkFWH8M91xNraj8zXKvXPfc0nsUxV3TLbBP325+TRnP9C4HaJqav8x
xgRfHBAwXYypc/lqmH+8HTo5lj3Gmvr/1YLpuvwFUcBm4ItfhRHA1j9vLW6D
6W+Tsr7XPZUqnfA5Y8hk6Xda5MhzPpnroreQHNHe2QhNmUIukXZ3j8fFjXc/
G5+6mkBdTlb+rNWwLQJ3VbDU1bUQYOdZEGj4WDMkR69HWOV+CY5N4OYi7xmb
Hdli3DM+IiWDidiBf5R5n/hcZtP0Vo1ZVbafmGR+vjoJvtwRmxAV3xCOJjr4
DqKGMj8mOqBw7AXra85MAfQaWX6pcHCT3/wBMMWU1ar6JjGcDLJCk3B1J4Zx
ybVHPZYx2XRqO5Owz8YY6cG9xf6KF3EgnIUab52DB5L34KO8qYPhZNteryJg
U8JPRmGHMPqpzq//qkidsGl/M4+TnS++cz71nfZCbtlV36MV+wi3xiLptcLF
qqsWYBzNhtybBlowiJNUFYcXy1RxxTPseqC7vCAuooQcdI6W8R0XseRVbrjB
CbLrTmbLvHAEcsvBcZ/rEH+KQPFbnhBr1waFiCFwxGp8MlbMcLeqeLOVQwT1
DFZqmHZQd5sllPhKRnZXq8qRabKAkb/iI1QDbbobXLcbYMUAY3n7+6U4UVga
c/vQNPiHoM8UkMpSiXhn3CYims1+CpdDbjqRTYN+NN1vULsqlEpeFCXYlCe1
1SuhKGI6y126S5EgBxGfdmzqyHUjJ51E3tSZrcE5vjJudP8DI2A5r3rRzKrD
kyLzyjePzDVW3M/oYr/AYv9hdbqB/rABSqXlajnrXznlY0PMWNQf2+1//S9Y
TAH2NnU8v7o0Wc3Vhd4ZuiaimBXSU76pQPhPrKx3e1GBJQ3bX2oWgPHBbMVU
1Bn1GdyiKJCDeqHZxlXa8PmI5aqhm7DPw9BN1CzWDxmk/SpBzkEEq7E8CFsI
l8TmCqOBnXjBBgYYzFm6UUJE5EJBH4WbFpuaTt6MvxjWJ0Kq60ybPPq2HT2U
m6OJvwxCoWR+wb9cs3sqpJn51SwvY3pn/C8oloFn06TGCF8QyOtw/yqHzquh
X9+v7FHgsXUJySYARqjz/AJufTt88MRCTFbMeuwfvv1/wVbGto6PN7W3Q/t8
XmHX83HqUIdSkyf5dJFHcK20IaCXWW4XDaYZjGZFZ4LGSurLvsBMJI7MpPAN
c9OpdxEtr0cYQB9otSAhaf+w4k5tvYo2bIIehN7h0iwTyG9gqSQxro/tqVFg
nTs+nAK5Yd6+STRtj0KWkZvBFoNZGP4E8ZhCz/CgOMxbRzp9exZpSkmictLT
3Gv02pB6YjQWyWm0NtRmRBZdbpyuywRHTugJ1QdA7vthfjXNiXOR4At9qj00
Z1MzNY0OFzYPVv4I6gJdzraIIVPTsIL2rlW+7y3OvgAWuWxMB9rtm91uDoKN
YaWBm2DkG1KxrT6vSOeajc5GhZGI6iold3+nSyj7kXAxykOORXMZILJHkY+/
+9Z3LLbJoBPPJmF/rmVl2nH7/DIAX9LqryGb6d58anf+aPm4TCTcUUzC54qa
4kYxO8lBl2f7ZBwMi0xIOE8fdPbS9y3uv5h0EQS+UcJ4wIa5o3pGuLwv3jCW
MD1AEtW0PtdwojJPh4Is99G5KOzrgGU76jcPdKdX6f3WliyMNbXhxmzF0+vk
rENOsj3N4rYu+SOBz9A6/8DJmXjMLVnjeGD+uTuQXGrsoDAsv/fPmKgkl4Ev
JLrKCexqf5vbUuSq7Lb9NRi7jU+r9myhqWpel7E/NEyhRQ1lelc9lw9AkLa7
2IpeP4k2YzFkUuY9xz/1MB08Dk3k0JC6UYVLzKqrpeRtVEWDCxj8mR7hu5Xp
23wWZokxNt6yIrpIn9+c3QJ5bZ8Fjec9l4eVxpKblAV9uo6yVg7T6qMESG0h
AGcKs9g3XcWR/ZWVIIREUH9ASY8l7vXZdQ2YwaTcMT4VxBdQa286/5MVQC1N
TRJUQo1i394eR5BEN7rS4MJs91aUYzh7Ob6JVAHaeQpA0FWOHC0kkibrOzEH
8Tn2RMZcqG/20muYa4UF+NPZShCpIIZ0aT9Yuw+QVzLt/U/cFpYDu55AZEOI
FhLhycC/RugPNOeQyCOiHdKy0wgQLd/o8ATaM++P7AG5MbU7WpvO1y7RXIzE
OPVneJ001rAT+bhrr+X9IxmwCkS+euowyVxY1AbKmHLc1OJ+1OKVpgeaaOcj
A1WuOEAyK7Ke3V72xRGQvC9oCG4ClXkzvaPJH5qlaMK13feswE4weMBE/cPS
buQL10yP2MbkWP0XcljSJyUVqGA/l9CyKworQXJoUbyEsidH7t5Ipy1zxuar
P1fpH8HlZRI9enrWWyCXWWu9EWKk/nkZGFQhXsFo9nt9d9NwLjaTlirq2c/D
RfIGD6ZXeIKgxA1rX0/mhhD15K+HqXW9LGFDlYtDZYz0vo8mj2mcnWOZDskF
LMT44QZxMO+rEHEE8zI/usm5Vo0ZRILxxezE0gO3b42Qv7zcWZCKJLz/Fnnk
V/4h7KOsZZcybFGlg5lUnvfuq7mvgTqwhHVnTvv/ZpdYryVrXNbnS4kmoZA3
yu2JBMCVPWwOnrriIeokYwlZyZcMBK0JA+YpWQKyh0TnK/BrXK0sJkt3GyFw
cgfA9jMakyOHU+VA/B1GmmljkX6Jr+8QhmY/vW0CItDKDlx80xFFQ38HIsED
r+QEYxXx3TGSowGGCkHyr4aCeGmpwTUKRAg7kkwD1NWaeuv2aVfVRApmBWhq
MmBeaZWR/ZHQfLLxfleEz9JTgDiUHk4tw85ip2kRRZQyHw7I8dOrbUQKe87A
pakIfrbfrTMa7fGrzDaE8tXGevUomih3OsgLfuY0KNxocq5/hCWbG9krTQWU
XBC/jFopGmJ/wNRnYidx5lo8g7OZZwU/ZWSOovsR2AnwX+HC5DNGgKIrRfgq
OIh+1I8CtkAIXEScau0cQKo5ml0LewdXI/sAsanm5bEDjdICTGb4EW9x2t4y
nrU0lVixaKXDOuCnT5AmEpUDBR7ONWoeUVfY9EIysaw/XsHNxxSVw+Nle9f2
Dmv/uFz1DOHNhGmJgRPujucNNjAvLz1f69qkFhvAy1orITtH0AtyO1maeuUN
9hs1IYnHYAA65OeJgSxawt7hX4wWEjkcc148jLXSkZ79BLd0kxAeLfMW4dKd
VWQdpJyUppn8wacNUiLEZOwVsqzeG1wY4VS+5KrCx8W3z6v7U6fInAIJwiL2
pypExI3mUQbWKvgw/EOk8p01nQzg5tECxIhM0TEAxclIaZ5lQMlyxtcHatzB
+Ycashh0XYxR8S65KlhxeQQvQ747ROld9EdOPKtqWs7gRyfIifD6HTAHwpyC
MhBvu46Yay/u/RmIXOr8AcZ7mp7mhEycGnhiwbZQsSswLkIOf9ehEYa+kBpL
Wkmd82+w6Sz/dDEGsWbqL9qxARP09nO+X+J9eOBbC+zPBp9RZdALOpjd+kMo
U1vmy7El4o2IJiYUgitN+Udj3iC5VWiienN4Ownlu0KoTAvUmgRnMx3OlTM4
MPXBo6IUfxHec9cYGp3BQvTxwXZSPYT6BDIx2V4cj5NSGVOYzu9Y+wFrKZct
yM62eewXZyW7uPVwTDo/Cs9pX40f4efdG6Xrryv1YAGK3JvLUM7Uw+BSaqc4
J+qiMDM5HRgFzpHAUAWstZQ/Hz7IwaGhR3SCO5Nt/NGk17ijhxx5w1kYQcT1
6S0Xwtnw/Khtj9nm3JMg3gVHdTONYXxYx1YY8bgWf2pQjh7Pdbxee9onW61i
wI3xHDwMshbKaquFW5Q0UMOTNX/Hte1W4Y79vBBO8yAvf20zfV7L/L0NY97Z
4cvjmwqPmgn52g1xra4HnfWkYp0QJu5J/gzLnTmYpRK1nD/ZrDN+Gn5otbNw
YsSsCKohuNSr0byx7CznWNpVrJV9NzcOTypFXVSlbqZ+R36K7y+uAGJBq0R1
xpioM+nJRo8URaR2K9I2zLfCNvZtum6q5Grmethv7Co0a4FYOn468cVcg7E2
q8YWiNCYtK2QRVWmt8Ut/DTh0V9LZvXhQ95+LTCbZdqKhn+7wr/c/1+BnlLd
YTfTb2T7TO1qisjWAbyfSu936tNiChZ+aU6cI62rCdAnKM1m3Z4++DFh4VW9
8VPbe3AIAMXkKnGa7hJEa5yySDx/qU1sXdd+pGt1/jWSUriENKYAPvhWT4oZ
H4+yjE2eSArln3hLIBCGdxhaJwzbAzKDUe+HSZNjl9yo89PFsmyQVI/2rDZA
XEs6QzjaUJAG0wObslO97vg/rl5q0LYN407T2Bs7pK/muxw3bHLe3vhhrsq1
eMpsi7muVBE/Nod1ddGZZFxCEM0kTbN1q6SDzw7cGdsTMSM+1BB5S7iCIIv0
bFeRwl5SOdpFU4C1MxjvLmTbLsslIjiDN1Bb3hHNeS8ivQbJR2rrCQLiUd3o
Ms/Ylp9yKKO4SO1m7JO4tp7kB9++n1WWoVx1X2x78hUh01eseGt7JvOtHEHO
FLGvLMIGFnPOgXid9ndPP5tfevLdJs4wWSyycGetc17XXLdrHpPwNqWeBY8c
I1uo+HEj0PBHKSVLIOv6JtgZ3RlRuyIaJAghCrK7sfaq3dbVFJJncJPgnCDS
616f/xJ1V+7oA7sbwtpB8dbFGZV5kH+a3WLklPyswoT5AKGTEu6zquXpKUr7
j+MJMbjR1Wz2louMXOmYXMmpPW4bt3EBYuuVFDyHuXLjOlHDV1rAGaIlluE2
2uS8w5KO9V3x6ukGqTY39oRnC7ie/TA/LJVqM9UrXaz415EEGZMwW0lH+UfY
jczf8SKm7rR3kPw6SJf1cR4e5EhXKPYYSljHvPYPlAG3LIAQVpXdw/AJXYX4
PZcoi83gPMJBGvSBQRrjVDCkFia8z4HRkCj2La29ZOdGgwhDmf08O+0PI3OP
V40UvfyXBX1yCc4sTdudY3fmt5E1BgRecRAQZYMUuT/z8nTWjOpGx//42eeh
u0571g1CwzK25+Jc7Yy+PmvgDIE15sFCF4ZOgcJJ71zwexyDrW1oVrWjoyM6
4gCAPuqs8uBAn6hGTs/TvchSti0YZttZ/FC7GdzuqU54V5xKOIhyLZhekmiD
RApAwow0bA2zYIKaLyXXH8Fu12Qtiu6lEoqPswfyjgnT3N22zK5uU86WClvT
yS54Poupq5o05rSHucyjEy1yTDXkdNWPhtx/D1Fnvv6CQVYGKiOegSVsZiRp
RxAH/2dqYfL5DQ1mombVspwN6GUu5nOfshudo1t0Q8HGPfGa4XWJ7AFkiyqN
tHuUkjckW3poUtzwISwX3x7oWav7QvRd4D7WkjP494KZELW97vPoA+PBz/AG
r+4OTAyXonAHfZiGN6KG/GspXOhDoDmnyveX6VFnmW0Q8C13X8XAZRjNhB4w
4xwYA54YUFEI3ip5NbOvVGuNezA7kqbJhaFAPyGFb6/CVqXZE8t+WbDbIZ/y
x9Dmdkm4vKQPkVDz1Dese1cRCBOd3MP9EWIRKLCEWziUHi19KqGiD/I+sO6o
PxyN3Yqlozu0XiBudAi8LyClxEat5G2iAX9Foc2jPMRAsLT+vsdGUDzsh9SA
5U0eqk8eGEfr/v9L02HjyPUtWlBk6iESYoPW5Y2zaerMUfTGTEcA3WddB6HZ
U43L8pg6MINg3kE7oO3rOov4/FkzQ9IziT6frzidjQIo9D5Y+3ugXoZgfOiY
Y7KJobWjt58NnxPjUtZxHrH7mviO0kh44nkrGShD545UIqF4QXmBxIl8YOBP
0yvqXrK/u+ilDXYiz1PgQxAKjm8cKd+Bnpoup3n0Q4BJxYBJczd0fbp+UY7R
EHuij4lvdmZ3uWNOidv+DQYtcnNDmZYx40w5kE73pMWI1/Dxi0eyuqvsO7i3
ScPxc18+yN/oA2oNovdWOcrXbEPXmuxmkHIxAwaFkTXqJQNzEtxWjfe7hacy
p7r5GVvwB5aczItKO3Imp7hbb7O60KfAzdHkzpK46Ia9wyiazNYFHVsWnJS3
C2gTWeiovfAIGwwKvvRqEOQ6uuJuqmHGzw3iilkf9Y3S6R6/4ZbyAbei/GSs
Jh/YoRu5Udhumxlhk11t+WoM271l+eeLHMrxXNhEec3/wEkQL15ETKeT/zor
oy6vHjPaqMwuYhjuMnT7J3LStgH3LqjOEEmUwSIw4uIe71wL68namxSxHsEF
eQ3ZZL2VInn0z9fvVxAsnTYWosqaKhsBK/XDfiez1dXguCcJe86wkzc7sUKO
/IzhjSzB+mYqYwEi7smiPmMfTxIo7VV/aZ3B9monGKrg+KTdxvDCahpUBVse
QGojD4Tr4BHgIfAyoXwOBg5RwhJZyspDGkJxzjtlSwKLO5vZXynaLSBswWt/
EW1T7ztCYxKBTbkp1kqKBRHxFNJhEIfwqS5vco2zsDndVH8TNcsGNBiNycpk
FvnMvFyJSTKxHjK0xTR+uZc2Yy6sDKtdck7GnLEYvLXmbx+/t9SYR17THFrL
e1GYIphGg51ywdWfEDEKYD/d/7DT7O+7hv79PDDtRF9rsukfbyuNPYSbrkpE
g+m3+pvaBoOzC8aGEx0eo8QC2OOkswGHnll2olvtJlJBKIcDVWMSyvOg/99/
2qWpZorcaWBRVkjafEu/6m99XkFmPrQ0OPJ16w8KbNdcE9cV9CN4n0WfSlgL
hpXxiQd3fm7YeVq5xE9GyZP237gDZxZJKDfpcrOks75CCGCVOzaEewkoUB5T
XX3VhfFSCuS0ReZ0nYa1vbophhB2R2r+FzAA9YmBRdVP2YdMFfT84g2ZBvoC
kR2bYQVOWd91LegM6dnZkvHiktJxfrZDT/q8kvCWInJtMTqbWQTVxTbkS9xp
/kBFmBgb67BqGyorqZazRXWnsOiFMrcpGv13MX6b1X4qxm+Z6ZGu1SNaw+9B
mN+AfXIWSNYJVPZz2mXE/bbGAkPMFZ0he5B/Y8ntY3tLxbMv39LO6Nl/NgUZ
+ljvHyLw4OXbYR92c6OkxRycgk8ijqDL8fFquBDcPhYglAgLcU10SGHwYrgl
7NUjhxYq7wZV30yIo/rXKUMu9/TNN/nw2GHhOJL4UqGIAPrc3k84ob2f8Pqk
gALInEehAoRVw2pxuruTO63874vYjLyIW0TnY0FAIIrJvuE5q4qwQ7x9F27m
u7gIWRGq57kzYpH1ySJHcNAlTfa34EUdgJdBip5bdRejwbtmg50giDvjJ0dz
xMdoQ9H7j/+oc2sWL9CXZmCbFVqWxotCZPeXr77IchnDsHwX8S7b1xnr6ZC+
zBGzZiEmzc19/xwN8Pl7IRN4zzeqTSegoyiesXWVNuZ+L3GaLGkiG2fcdoxw
QhPwcxCLqXeiB0eXaQe0Acua6JoAS3i+qxXG3Vl5lKYsml7spALuET0aEScN
O+VFANQ2zu0hZgjDJrzhh6ZhsQLj8+5w5c5knDxJWUHLU9hYvv1IFdRaAzpR
9IpA27TsSjgraIqSyYIxJpyGnCa8PTKVOv5mu/mlBT/sGyNJiZMvODUcEedB
Zeq8YeCtqNJbfnpU0YKIvipJAr4pnfSXWwhDAkArqJEqiZta7/P9CgiaW3ji
3kpMpO/EaO+JePnfAnCvumMrvCDfSRHG/MEXUCpQCIDUVQ6Jc3ZIrlEE/hZX
VASECPp8m5B8cIW4IDVEb2EO+1kxW9phXQhYB/jfNhr9J9P/s/c2sEDq5vKC
mTqRbyNw7UwEAgWYeWNaklGxUc55jU8H97UtVP64PcjEQX8aZMNRJuS52YBo
1dshtVgMG2SM/0AgiHya08IQVzaQ5wYujVGiNtiEyIAthP2mQTNNYccMuNU0
y9o/RLjWydQ0mTHfcWzoiHpSLEVAvIGpO6cckwPBJF12jW7VTqzUUa5EAx8C
UoSFxshgvdaTT5cKykA98QekkpEV4kvpE7C27O4b6Toon+3bfrvLwD85IlBN
MZPfC3I4I5NGqGaKM7d3bZNcLIigRHOA9EC9oqC8Os7ecs4PI34usS38nhW2
4xrQpOTC6WXoIkrA/PkMIFF1VXuX7aBe4AP616dUrMDOBdqPgw4xAGkMSc78
gy2NS8/SOa3agmcnVk8hq7MVbBK/TY4GXC5q2ZiPxRPlENA8ITJC8vUIvTVA
wyoJ6ciYkuIyxzgu2zP34VSHzww0DNE4k14xzE7QG/bJuXQV68FwnQy+/idp
5mzxaMbVANfT0hYgVZv/uB777fsCLKMYU6RgvSnYh+rk0eD0UKXQQBfL4V5p
t3BBjkUYiIkJPeqg8hwaPH6wfrjFcirVeAtXsiol3BwBNGx2TdvvJl51CzLz
qG0S713AdulhfIGeJ5KPj0gCQ64JzvrrmQ6MUKtV66YKvPYM9YAsFLQiAjf3
sZoxUpmqvQquqZmiCdTrjbs3imaYw8f+y8KHrL6ca1IyR3Xsm+1T8Jw0Am7D
QG+2dM56rW9q6tr8YQ/s8lmub7pnbtduC0x7P7ZyR2I2O7a/E+GKcjZy4pqP
gnttNu5deNPg6Li6LRbQdDYcZMi0x1dOumJLFBPSv81MXHDS2oyQZVNFe2ST
vYLmD3DvZ2jpvqfvpbFRKN07SHI6BTrjYhCWbbbNakePTLIbBt8S1RAnPyjl
eBUEusvp/uHFOsHQw/JdFzQJpUOAuzbGDQDnpPy7OiuVzfgBnKbGhkgEfv7m
J4PBJIUgMOj3T8P65bu0BiAdqgpjJ987mwc7bS1u3JYwbFo0k6Chd6kPG8LO
YdqGLB5WlxHIgS9/WCCJquDWu7SSHswtaDzK4XzMwvOIeZHuCBwUFgXQ/+P4
JuWN0tQI2kRglGqIoj+Pyd/hiK2rTF7/BpiEDBL+uanXFTYI872bYvgGncYe
4yNI4BT52f0vls4yzbnO7BJAAiQEy0sEH/lVBkQ1MrF1vpO4/W1BzcGo/xFM
BMJDnPLo9f5+M5yYe5fwsp0pLwEQvZZOCH2grUhFl4W3hfbn44b08iXOPqs7
YKwnyYRniT7YFE2stvw4e+ja1D3gsJpsQ1pWyJzxmrzshvNN6wfKSc12fRz5
0d3ztz5uoN5RK6gAHQAmddZhqw0QWDHilZ9w+SAOd/EmHhMg0vqPbCWKt+RD
Ukg3Cm6SIgwmBA9hIm1mkmqyR3BUi8huRbJTtM/Kl6b1jOcrP8fm8JPge0TD
FXcBT6jRiHv2z/txhNGI1KVoioV3gHNFzl7rWSPJ8GEeyxTImccqjJmMTdi2
pJdx0JTGx5EmjsV4yuQP1jcjvzAO/AiJRWzJkYzwxlZ0RIdrzUTmkKa7NDix
8aLYxId2LKt07DB/Y+54kyztOx4bZ6u1CopSKLJ/78+46GMN1aeL2fvgw0NS
vAFPSELwmARURDcv82c5NJSXYZcpiEn1/2WsYBBeJUVXwjRXbd5bQ55O6cZO
zJYRhxcDGujtt5G8qDTMG9A7ebpEDGW4uCWAr8Sdh2cA/WmEMENvtUIWvMCt
K3JeGROicNbS361vJYULr8DaPbbDFLPw6t78ioC5S3OAzeRmA6QdJO+us0UQ
E7K1Chm1ULSCqXDhxgUDz5nuwLZyS+6+BJgSIjnMV2s9HeLIkC2Zu3H427i6
MIak2AqLhCRBP9khd7kVeYNIWC/jgzQ0I+ebRrSl4C9QK142Ycz5jAYgZFCV
rJMqxm+YiMrEB9rmlflqQGvJGnG3WvAzNT9qsn/HOASuTk19v+WY00yHLDHq
a8pTxpoBighdQvdCnZGIpL7Ji3Acn2jErD2ASm0DbGYBy9YqlgO8DDOVxgsM
7TZk2m5N10ZzbBcP+jLZIY6te0FtY/sAzOd6XFUZo7mLYq/phAbnbsy/UnPQ
PFvD2bJbzAl72QjsC+ogVGxyN9qQ605/+or0mvlTBoVKvVi6FiHOqUC/uB/m
KWWK2X1kEAeea6jk0q5BlsSk6PFPwbeLv3qIdqFoFrCGwAy8mE6snCQJ4jcl
RXucQSZfHrYRkbYG0dvGfCScxdkUquQQug29XhVb/F2kMny5G+Luub9bLLWk
wa1bAazRqczUOkhSHvS+cnOiDeuKktknNZje5/1JpNtIXsoKdVvTsuW7UYs1
58nXZI6DUPdUn8Mvlj+6EcDNOFRtOx3jSJ0xiNIlIaQ4ayNE6qOeKWbMtfTQ
M72PHOeTs3wlHjQFQLsP03IXMb+XZG8Z1sqCGW+cqASQhOC32nm+oHjiPP9r
sAs/a8Ol6cocb78qSYNG2Jx1/qRRBzSZrQHINeu6+o4RfW47IQW56wUFPof1
9UAP5XJRl2bWdW+EJeuMPeZyjJzyLzIYmLq5J6PfZZC9D1sKrzbhDdIlw7fp
Sz3keRsUQBtghoY9nfTibuwKM7fCUI1OT8iasgYIjZf7PJBSjV1yxah8YAFn
Sx/BNdfDRttyKWbgiqnO8b9tj/vj7uJJkUoZ1w7r4OgvKXIrug3i2VYpySi2
UUOsKJ6eZhT5uHfVha2BaDq/R5nPjjR3RnFq8cnrR8+1gIySPaQB9kV+0wtT
e9c+Xks+/XU7jzD803SMgSAcw07F7FPEXTUhB1s/9KIXoIHIh8j/ENkNjsk7
eOVfjnzGNg/mg2tsqISNG+6JmZf84LIK63+GvzD27j1rIFAK7Ht3yocspqiP
c8pmgWul/bVUD8/qBuccNcH2l8hdOYegY4qLasUryUhS8daCTe+uroyKeUBj
WQ0RAdTfvJkiJS6ymX3EzClOX98lIT86etwo+TWiISuj3OC+Qeb87pzX9A62
ehxJxDzYIiLvphIHFj1op6NdUrS25QrOB2cJCZ6OYsg/BuybiyiRYpRnJzLN
kn5O1LAoRhskI7vxwUkAw4UfWAyIlPEdIjLimI1/iEMwIQZmo64FqjbokDmO
fqMk3MTrrHCh7i6D9jcje1J5IXFUL4fzX3n8zC2ny6OytqZTu4h9u25lGY4A
w1gWhGeaZZhXj31XP8ECrFSrG26xK6x0CZ0hoRxA1BykmnxeV3wjLdCsRZJG
/9XiMZ/fKt7/ZlCmLpetjvqRZ6Byh1unr9/IGEZ3JtaeLPOAc1xWzuBZPn71
A6ZsdEw7gxs9XmtWx4mIzUsYV8L/FiTr6RvBNbUkxwJcH0MTXo63T8KqaC2J
hWky1gagUfYptzrMTti96ISJxZvw1ZR9gy+HVIj+7Q4W0yHNu8vAKHpsEZ+u
gq8/xY1jrkCz4L5cMUuhJWDYqQwEt0SHze1PH2lqM8SxqBSapnqLcMA8EPTk
93BcOwnnPCd2Uk207BeVUaeSlJHPxdFxKHzNl5GVYyH625+JOT+a+QQ6NjH+
Qo/zjGrsFHQyo9Qaxrn27yApIpQGXz4oVdb2AnmH39LJZRXnNASxWivGgnGx
5M1GZ+socXGh9c0I8fOCgwqZbNhRdDEZ+DzUdHBiFWjvbOjvR5QMt+ZT6ynf
GL9xC+/7C3P+ZwdO3yWGqhnOw4qSXY5an7hj6gj1K+vy8itr2vd3NxdEtxKD
brX4kVWHwStbVp0tMGX3gu87dzMIRn0Hlj+adBtDw4f7IuQD+Npf/dkCRL6+
uOPHS4jXlmYHJDvGx1yXKCuhSf4jEHbaST8nYhbiWr4wt0VKmB5IwU/5qL9g
av83PWWxmGI7NGnBWi9DL67SLS1XzDB8M6g11vaCcgJ0hY+/LiYGu3XPu5lz
bvBBLQHe8FHcDNAuPAOPBZpm7VAIOq5iUCeaITtUknpSwdy1Xlx2ywwvtUof
QkZlYM3OMXPn4KX9IlWrS+ZW9D1NiHVig4U5e4dAzTV98NdAms4z3Mj9cW+O
Zm9lvTxzRlog94WuTwWJeYODWf9FjU15lUvBBHGdV0Lan9sI5p7gMceNVznd
HgGCnKbZCpFquhqQJJhyD6a9TcUY7xRicAkvOH+OmIyP3KOEevmXiBlUYACt
iXkZ/punOKlRcRJU5zwyjfMgMy6659g0fQDF04yVLEdbqkgGyH88EgDZOjOw
6I0Cnb7KFAOqNL0J9RE2bZfUOfYbsUYpd/G9x7v8RjTBW7zSxtEHwY+aaMc6
rZVUcC875Xqsen+z+fRqm2Vzbvdgnb+fbltLACCI4XtwuYjM4YcS7gJG09Vi
msaqns/IQhuEAVrs9gDM9zKWObEtVnXrh9jRXWg89qAhoGWCpcOTtL2aKIhH
B+h1mCxWZ+eV0aP8jaeGjj0ajTkbIC7JpRsslfSqrnLOs24MW7vGTKqWFYLv
H6Z0lng+COle5wPPYx19YYJiTJWNH5qUeJzvDZTfS1P6Am8bOKxW67Tgbc00
ZoH0qveyUGiVS3c4cGAjZpMrguu9BRswrWtLmDeZ2SYnv8hekOccCjeQMtDm
fMblQ4GSgo5TG//+2FVQnvG2TIRFBUT/63KQpaN9TLmK4QtYoe7j12JKH7ri
tq+GvR4UmoHWOgZL92mujZAdGQHkucmd/f5QlHwn6a7Ux1ni+6GcXHF7abx5
kvWrIJ75LbKiVMPaCQkw7x2p2vVW4LKB740fFm4XUSokBS/YJ98gJjyymIub
zFnfGhcmxo3hf5F/Kej+TNAaAxeUhI/EkFw8L1jZnSfwMKfkDa+BmZ1K93Pc
v2pYJJ95LDj4F2JAl/hzHTU7enQxbv4Sgy8ylBSJ99cw5Z89WlyKqaAIOPrd
TfZNKEYeGi+ZuZedJvL/gQ+BOAkgNZln7a1wzSdDbWLGYWU1eUiHLConXnlA
WA8OquU0juleS/1unP6sYQTpxQ8Kr5jpudZ+eVBUllFcU9vchrKJzw1nvSkL
MuOco1nWv2U26ZX+0RUTcw342+lLTjFeCQCL7casvxidHPIM5RKZ5YKYKB9/
veO9rZD+F0ucYvJVBOWulVBGGb0+8hQXWw0m6QGrTPyZNhzjZnXJByRecJO9
mczDYb3XhmXPeozRPP2cxe6oUeGys7r8y1HB6CJR99dnypZiaMh6rd16bdsk
jRFqkrS0sQ3CWWPH/bPRbj49ri5I2UWSKOVldwUBxmg7+INw0t+6e+EEnWVr
s3LQ696BjBjhzJBkyvj7/Smd7gxQEbYOyzetJGmFIZiZ2lz1j0sS4bMy1Hsr
Isu16tau9/gLhLLdiRH0crkzg427mTMMDXZw1S8iWB1dgh3l62rswP1O6VM6
xtjFi7ThocI8z1Jl1LN6lx/P9ZoEB0jqLe7N/rRcDvtoa59L+b2JK2kN48CX
tqN7tQT7/t6S4ZY94J/zVzCTSz4NX7nbSt+jztA5dVU0fAxb/g2rpihoOMxU
0sdCYbxqQAC2ZDxCkMUf8XXezyiJ5h+Cq6PXWkpVzVgX7nQQ8AKDWFANstTS
3z3sLILQfd6J+CL8110bE0agMBy1JlVfewx2lstKL2PThc2FWk7p+7KLOAtu
Y5lhmb/9cQIG9rQhuSQWmVPXyKSRxZyFmPEe39MEnh4LKm3aTIbYARUbEsjm
2mQck8pIU4UK0AXBp4Vzi/iTSrvwtCaC/VzPl8nQPpNel1fvav+0X3csBGO7
+zmD07JLkKOzIglFkWRohiD2/lcPvD3xRfG+h//KVwSjdj4DtEEbZm9wclf0
8m3Raiy8Iun7TjpRoopY7YwvPfLLDe+M4QLV4MmdvMtrI5ZJWb2VXvdSUVOE
FjYvaTjefF1nwW6z81lbzdgek2SAd1erEuowu/WU3X3BMsfu1KgQHeTN82Rp
Vn+UUzQzcUbR0Jhq1jyyvXeFt/te6KHvp/YV+Gurkq80IPMRwJ2PtKSgbJTG
nNUG7q2MPVylZ0XdVBZHbxCF1qbz4cJ4vShJKg76pwTSmoT8LlmND8edCmXJ
nZRPGVK9+v8ilPPK8AvfnwP1doqvws7nLuKIEvupKwZwJDCe0HhXU2mtM5Ty
UoF7ywexPcGOQj+2SW5xb3ErtdwDFXjVtkNmIu3OuIDRshGZ2dv5uxrs/6v1
84fV5XsUcvrie92/dFnWjxAB+cwbpnm2cpQ7bvWGWJMmRG/tmZQuqpH61OiY
UQ8UhwMeX4LFs2ELSmfh3l2MCp8Vb2H05/cuv3LBJok+ei7mu3KBIk1L7Jd6
ZUXyX1K9ErF883nNp/0oyDPBLPekbBEmt/porJWaEymioTh9yNJogS3FddKC
mZtTWEEHl0AubK1dy+eWqzJbPj7LtGi6BCPLYFQ2JjwIzKN62gRp60l30azz
lOnR28qv4KsVPf+D9DmsDI4cpv6qGgoApILs/PvhnnPne8vkxro6q0uX8gjd
8ojS9SS6qLDJRoBaBkZGuDJnjhqFZJG0Fo+DvhS7xlB6XCaIV387QXuR+KS7
U0zyUC70gr++s1ob8LWp+lcfsWhM6HNyfyK3syNceXLjy5ZjiShx0F7cl/o/
rO+9M0h0PkWBramKd2dApKtlCtVl7DuQi3jC3r9kKH8KRcVzdRPyk3HAHUAs
rojlPxc6PkUxZuJ7jQpPTtmMrE2W5LbMAQd/YurIZsbe0OYO1W2VmaHUuXs8
tIndMt/4GBTFuurvqnsgTvepcbsz2aHEJtwiFoijDWz5TxuA8/YnyI8jo5tV
ytuv62AWJq4Pvvlp1GVSZtLAcTE1g8z+r+dxQvYz79gk6IOp9sE20QrSerZ4
mhDiDN26atVq19cvL17GOUvQRWdN9J/0gNhZQ0YvfkPuVXJ3ftCGsOQMEAcb
826CAtdYAwK7eRi3pnaM3HMQ/vnpEHCxRB2eJz0i2BJlj9tC7mUhIY/Rkr/F
hUe1c9OcTWQSlsTmpceqoGG/XXIZ9tI8V2b/Rer4sTQJghj09D4n/n16Kn5G
4YUBPunVo5NN/Po2N3k7pFEUXTi+BMQirVEUAJ6TUH7BN/psH2hkN15VHVMS
w/tL7YYJABNuJeYxUD9XeulQqlM87lSm/kwPMuNWpOlR1mVlyk1iOh9szFhv
VLzrCymFUx+NfrL+Hqaf9uJefQcZbN71HaVg//EwqsE/SGt0r6I+I0o6Y34t
X6a5Q/4ZBO802KJZZXTNRVYkVZRFDaZ9H27FxDCPSV0jl+4jyQfk97UXxbWL
U9nuq3KnrTJE5vGEkKsUlxR3cvCaaZ5urkQ1ml+h/NuIxnQIk7DNLRHR9zO4
5r/CCamjZ/8Xg2gjq+IC0XF5XZxS0tRBrx4i4zVK7Zj7oNDnddQWZdMMRDM0
cvUoDm2RL5rymC1PBmwA6ffdqCGDRjqJQyu28FxvjB/vCf9DSfL1KkVqPRmW
+WKMCE9LHZzpZyF0ntOLHqckQ6gWSD+SfY2oTIN8QK4SeXeV8mkv0AZDX0Cc
BJEhd5N6mpYkWMmBPm8mBuJHUAbI62lvL6ka5FnLHLjtMEDGIyNIYXGl3MzT
+SbB7D+vGZHhcgtkTQcxh+C/SZZbq6f3RJ/m8nIQe3EyonY0TRuANsu3fqwk
7oUxbmEvK7WX8epCcc6nYNYceq6jIh6K68wmLx5FrMK50FXVcjsa4Ad8Qnnf
qXYofdemTRni7zvA2oJN6JLMQYY68qIdbnd4Ctzwdftj2QoWwTTNIWDlcgmL
vQ2udiFcIu0a3z/NtYVEcZRrZU35SWdbEL2IXCzk27pGza5aitnbSwbycadH
CckEYJ5mjx2dvdSrcOQa850lG+zjFuNbAJGdAFj937V6aYqeWQNn6bYm/v33
b6T9pKcF7eF0ZneqJsuFeypiEfXc0nowlw9he5CCGRy0AsH3f7BwuK367bec
bfKSrBsREOQUNk6QQE6jO87MoPrHCefxuDlwAOUlAWDBORNR42rwbd2FguVI
YLvMIVE560YJpc2DaLzQ/rnAVErlNJR5rBhSbQ7i1DBISNEt8krYANXIHpLR
vidgsbsKyZscYIuSdvSpTlXyT8euuMZBezE84DKJv5wfaLnBtT60U1jTLhRH
JhcREFr6dJSqw5WJCIiWibTXakFkj+UKhJoVxaLlh5A4zQTXhHG7Hyp5IGLv
5MfIPJ5aM+rRuUUs9x3LTuZCputhpWs7CII3apyDnT2YloOEW+7d/PUhUymU
mY9WDHuU1sWH09iUxTZQdGjbFR2YBHT/psX3YHmUhuWqqc4k1w65UIJASLsC
I3XreYKwK4c3yV17WLLt64Co9qo9C0F1cmxpyWFA8VNhaCzpdjm5k2WuouP+
qf0jrstxNQ7UIZ3R+J/l34b0hg7z5RQVkw/AzGaZP16zLz+3+QJqeh7q1gi4
oLT3DmM8+XymSS+f88FwZp6uGoXdLY9oHdArlIZP9jivT4CWiw/CL+C+GDjP
X7tiX1mpD1cwoGihjdOJ5rgnUow7txFtnkGEZn96WLK6iInSFDouRHnsq64o
JdZgBrXMj+kUE+qWgnZtSLdC51UrU096KAFELJDon9uHTbnnImsOpzC6ZxcN
rPcArb3k49VY/24O2p8Va0BXkCS2FD6Qn8li9p3GFmh8D+86NCkTch/YR4p0
GWsTXyF1EGGtBU1y/pgV7o/61dQbjtxYY596fjDR4CpRrLKyCNHLEkAJF81M
BdnI+6XEy/APTM9X+8lIi6ZERkyfTVRuNkgGIsk2pDHgp4XhES539x20k4tR
S85LkOEucBlfbA6utviJvxAR95nue06StlaKVjEHBStSzc/hVCIjfeZRUZw4
oIDCYsu3ZhSee6zCKbMW/1259Tir49r4rp4SaODzqYKEBoEhIdJFiBwEcn72
iIehqSYaHzxtWAmmDUz23A9n8dZlcOwijT2Gc+pi4AZTIbcMgI0E8K970kgU
R6WuaS861lukKLZHCZ+HppmWvm7X4OXjHU0xxikmUc1OossjMc75eJDzfV97
uuI7PW4Mvb3vqh6jrOKe+tMszNt4w68gCsG5c2lua6/y1ATncHMPYCCg43U2
la/oBTmKVnlknFpHZUAELqoBR2on1dmUnbpYGekE02WCJj8JMk+Q8QiKi8CJ
uhII0w/gvx21unwQGWiSXz3pZL+d9XjlJEHxoz8tDBTOoUSX49yQN1s+7DIA
RtqbddZVkc5kyMulaNu+9q1fXRkSwKnfrwA/dviEJjoHxTBYLug4khqbMZBc
q796o0OQKtbiVk8WJhVK3lmfX4pFCSFR0yJKYrqthWjpobl0sgGjpgpLhAD6
GTnCYMDffa5i64FpgHdD+IiaMbAYobVKB2CXSwe/8SGuIRFyTRdDbwnaK5x8
WOMiWeRBzCCrg0HGvjq6GV12lUdQPz/MkigIRqr2ELc2rbuziU20Wzxxp+lp
Wuueh+es/iK6rCe5O7C1w4Gwp0COt7oE/a8iXVk8/cqVaKAR6sMvxu1KOqzA
9RLtytNAC65xJanv3lO+oH1H9XEFUiajrRbjwTNbZFwZ1KBQFPi0h+0XbD4d
PJUvxPqikhlUBs2O5bud/j/UC9/dHsCASjXLZ0b8abAPN6JB4W/1NTlPdpo8
1J9I3PU3QUT+mlXBAeqBoNM/nSTPhPoMLexXjhnfyEfuNeuTOpzyESLwrVUf
XfR0FvdkF4ofEE4zdY1CwX9OMV3HyJYbbxTZG4pcFZ9gkIvUyR9WQz7RPWuG
M34KtJ4iRQ3bCdwRuH5RE7oxTnuIDqEMCNvWNuJBRBDZZov6rYusuU6sYMY1
sYZsbBng+oiGNN9Msyef5miAz2SkBZC9TcBMqgo56Yl85ov6EnNOGeeKeGWG
86HmQsULT8emhm99m3gXwriB4M9IBHL9iN6pnVCMzmQFSlHaJnidLKb6JRo3
nyyIdKRwspytThnhJbBp3vZGAm7pIll291hC42476/rTMFJDC3HQazEwaTrC
LqswOr1KdCvBMYze4lD0xb06HB+ErGc1b77ST7KOqk4Y8w1WmR3gk7xVibEF
0Z2OFG0ERIvDkJ/Q9T/rKmAEN9KVvRm7wPmLqpNJLqHBGopEeXvNTsk22TVx
h4rQmONr28TVLSFr73YmoDYbzD43G7oA7WifCRzG7GPRmVwBpdxzzDR9smsX
TN2pX5LG8G9edQ+3wEsUJMW5iwN6XSvY577r9QSW0XfI7k56/3SrsHlxjYBt
3NV7X1PBhb3rjLGkwp/cBY07vJxNM1XSc51Jnb50E0/Bnq1myggbio1kJK5E
zIfC3f4pzWNAIrnTmpoJsGs0NPb0Vbz24cSJc1rPyklghKLIfonYI9croKoD
xO7/kAffDateuyXufeN/HVEYvUxrvepNeoOmDISorNi6hohOTtlA9bbr8kIT
vXlRZGuKxQO0FnX0IUGY217ghrBOPqQnpJvNRq7ztIttC52Kq3o3nCxIvstQ
DK7Cth+lDMXPXL1J2WvxG0Gy7IfHTn4ImV0IatDd4oH/vvVkvJqse3VHfIJb
z5QQ1z5Sgdk+NjA33wPJGk7Ck37p5o/gC0PanPEKbCoRqrs3E2s+5PoydaTs
tV3D6mdmolHPCAlF7kcW51KMtB/9nmySakcTtvILYkmvCe4Pk6Jr7jIYcgWG
gwIsa5wzsquFuReDRupW9yhQQPElv5WMcDHKxt1Lbald56edNxQSPmtG6m4h
3l02UBfzsQjrAmEeK5EAWBDfjBl1VO1mFGr2y+vjW0yEQr3XdcTti4QUyU9H
JW9/JNgqs5nZZv9kETQmy7T7TsqswFmjm6UP0P/GF1g7qtkAoS0QhQ9QRg/u
QNQVVkpxTwKKb5+7jJN+C8ziLsP4Wzamj//MRO0NY2MNVQ9GEWFDHZw/dhwX
75h82c8V4wwUxBUJYUE0lWI5yQMU48oH8UCTrEUqqiNtGsNN/boRWu+F+EZu
zrkzvCBYcIW+KbzdteTBfLMCyIA5Ihu98DyQy7Aglo8r0YOaqZ5ga2TRFhj8
2fK+M70qWMGT3vru5FJ0295e3ncPCZHm83LDb49BjEbpxSiWwfK4vMgZD+gp
ak51Hj/hN5FYpm756KgPfQzNoJXOivQDqpLqNGm+k62yGs0Y/f77Md7vvWNC
O1RrVgLXyDROEdONlwRb052HpXyI+ovl1CabVbZp8Qox5VcI9oh/VDMM6MVO
7CJWAcde+ESiwCFEDojmVIuos+bmppEuorQAHbv985xtgsBhUzAc6bVdNx/p
YzXpLft2d3QJduxW1rK0Yf12g4xWpftF7nUQv8xCZVwfKcvA67s0l6Me1S5b
Ymu+GySujXeltLzbUEis7WWLOG8N255qLAQmL99QMYSJOsZZeO5OnegpgL+M
ZfPbji3UdyYWB1QObyvAXmKcloW6GyKunyf/axAt3OgOzLFSOGKPG3YV0G9R
n7rLKqI5myea3zMB8xlvrUUZ7Gc7lJayz5RLKJH1Mb4ZA72/Kpwenuv+PHIm
GFipbbCHOCmzW2EGN0B/DgFnig7uHr28n039Yub6Tuj7lHZsPJP29x1/t5uQ
CuXt/7xJtv8NCH2eoDAdzb+smDYEytpu2n6CrQyDMAVdGhYU35Lev5fenpme
O7nuJ/f6G12o376MEDtInoVB/UkZLq9p+SqCZZF2P3rXo0cnfNMnh6HR7W0E
1h6Np6H2dUvvKQxbrYr7SyRPAQV8pkZqa7XOB4qScpqJFpxC8nVT6m/lmzWo
sseK153jAqjwUN2hvTPX5SYz2p9yPv4xweaW6PHnTQ2bXmrXKDy4IhVAI6p2
ccFi6nFx5B33rt9TXPJqIo1RyA4XaKNNTJyA8HXKJTB8ek6bzo/HgbkaA/EN
bSWMqB44kE3EaI1hP9bfd6zLHBoFjmeJ5Pwa454fLHPOMJ9dx+Wof0HcNX9W
un2xvY4s5KKZWUSXYXTweJaKcHOOXH2ty5VhOPouecFuuNNBtXhPNBNah0J5
nn7usheSzsO3hcrJzphXGFigbknXryirlO+5r+PYgcvu4Tc9TVWJlGCDtASn
48ydCUbbyh9f/x59aa0fWC+5512f3RJvuQUN9HDeTXhqAzIG6MUMWWQhhNrA
Mxwzs8MxygYStZqWqhg7xZOlBHwKq6PvfC22DtdzMXJdGQb9ICk6qd63lJUm
ssn6a7r/R9M05AhcAkEgvqsACS8yDVU7q/qOuGBC5Dfakj/oF8TJQxv+bIUL
xfDxEqmXSp7tdpoii5R61TYCcP/WQxJYNy46AvOdLAAOYHPUi0cqggle5yg3
X0SwMzjOc+S08mGHICh6Nno6a8jwVMaN5StLAvpXG7a+GRIW+fvwxQGj8Els
m6RZl5axqZB/abY3WYS+nwKa9M76MKx7uZY2OFqiapD+t4sezBe25t0N1k3P
Dwg3YKUMCj4NysEM7NhxSal7Kx7o2sMzk46cxs3zC/vt/6qXXDA5w9K38dYQ
iciyZZp64/aDuiVAx5EeMw/L9PP+2cdq0bk0E/rAmhy8K2IyZ3NNHdFqgEOq
JkFh+nlzidFk/IViUuqvprmMPv2WR51pVKb2mebla3POFfMvg8HbDpo+gWAd
V3tdziySnihPUHNMhWGZ8YF+aem1W4Vz9a9RdrlG7YEuQSugDCPQDVe8xJPR
QmpQU8UabEvduGGx38fK77IkCgmEpFbmLUWLXFrlt6JN5Z409vhQXqEM0fxJ
tKi7jvWVCsceIJENSc88OdfguhJ5aSA8L19nt9ZbYIxoQVrlaLN+RKMfZNqR
orHDG/tnYPz9yxNH9MRGekybCxFY50kGZ8lWa65QYvvitHnv1iKZ/4u+z0hD
Ku46WUUaGJdtvKWnY77hJ1mHC8gldDcRJcXdYQdlilig6hQMCIgQ1Eom7ps+
Zu6p77EuUidBgLGsT4qMSE0UPTGrmfwZ6mhtIXI0BajCRNwRSvmTqJ1V01R2
5E3c201mu3Hk61iDxkYn3bSitKXlmULKtnu3o9MvUS74BTbh/mIW+TvGoTMD
2A3R/msnQo7fsx3UYBm8fJd8yex68AmTBARBfOFhLumLscdHDSdHcCYPoGXg
pCx8ec+AJI1mihEUnt7fRfA6h1xBSeuSYJQN7qix2qNxs8vu+uFKzcJxBT/5
0jyZYVShDyX+1fYZ1gM7EAx+KxIie0SPw2y8hKE4Ig3mKGivuP+eGXQytNJ/
3/MCLlGuuE439l0ii7L2jh2T5ahG6ZDty3YzTVHabZtTnKwGv2r6qyJ3TU2r
t8pU+yr+JpT+s+sui3NiP39kLc+HsZLQQPb923IQmPj7EpuUCdTr9Md2sSGA
hhYsPtVuoU66fR+LxqKWvSukyAsRxPJW9tkQvyMRzmsxKLrrr1RzSQnqHv0r
78ULZtflKx1vImOFrfw+G4ybjAFb0mhyjLMXwxsYT0lQpXZqKcPD4H0LMrzl
jxQcfnpBt76CcX/bm/JsnCLlIB6yhgZkV1qjX3K45GSFRGXPvU3ueBCc2NkK
h26k2fr5b2XL/Nx20misdjw6eoUMm9waligv4XbrVZsImB8fbyaw0Hmcy0cr
aR7U2QtIHs/e0xYyPqDCAZ1DtqdiiaL+1sZJPzIQHQXPW4jIKDQs3fkuzXTu
looMWrR8Bctyn68fLEEbKuaTJuUBXEWltQhq0IZjwKnPywg6hH+PGRS7t8H9
LBiVc7t76vELqWorUngqTjbWR6/GZdEgH3W6N1B3wGBqHuFHY6tfMDJLAuQq
dnzrZVP4igt88PZJE3NkTzEigQ+q3FL9Y7WfG91chIPMoOc9muZuXt3JS4AV
LcIuTx3WX+/p/9+Sij4XAl3UsSch3m7Zlm5A/SsjZiuKiEP/7MmFS+CgfYiK
50Dj1Rz+EpwFUf5J0HwgO8hableehTEpOkjLryXbUCGBkvdiNFCyf6DUn+y9
/R57sl4jLI4CFcaJBbvegGkZAexb8ftYdlsAQA+PAHOdp/9p9hOpg6b2Z9Ob
+n5M4K5CsleTR6DPd9JNYxItlKLg4ydS+eU52nQMm8sZen1l0Sr6ag26iFE+
piCMR44nJ/VwmX2/GlM8Pzyn3PBfqiifQojMlcfRwNtMV48xWhoA6fQLP98H
TUt6tka4Qug4+sAOJJP0ZzM8gS9n8aU6RlJPlKp0m4bV5ioxSanbwTTv30k9
RDCenvlFddlUvVBwjHDISPMKj24zsPcOqffAOAWaptV0iI6oZTCdahVSMbIr
095bLak+ADSBHJA6KP1XKL6uHrbeL6Iz79Cv/bZcUCjjNScz2NZjFD71JplT
gql9fn0Ny3st5fl1jmiNM0B69CAB4lNlUl7RGQqyp5maS/2Y0AtLCCdzZLkw
7KVeABFyGAziJKYInJR9hFzyHF++I1kYh6TYXxHrFQ4kTuRjtW2r/5SjDAeO
cfJn1FsFyha0GLdIm+k2pVucr+c/DDnZVJx1In2T/7B7XZFcBHBNXV6sL0x2
UgmF22xtYKRh2gKVBArlOlyRzdma+RM3QncZsrqSH32F/eV4Ha41GvQ2fcNx
8Evc3M8D+g2QK9B5PQkMKi+nTo0UDAg6VtngKYzlGri8XIOBZdfQLj09VMGk
mkw0n2Iwn5cvpiYGRlsSdmdpkPsTdh8ihf778fCINsMxsjGBzw16NipLjmzn
3atsjk8KvggACDd76hgaF8ncOlS4nMVEPDmGQvpupxQlXse1rO8AN85gQBNC
3ozmuECwUlsu8o2Mp/b0CqI++SZcvheFfubjczYxYZOERrFpGcYi6zk3wWhS
ZflZTbgMB9am9zb57oRQ/AWDgQObcvOqnyUkLk19Wu2UCyLCwA/CiQSsQ3uJ
wyfN736KzE6Q4TJEF8LKscxpyNiDXDUzgMaRiV3PxH7ucYuokA3F2A4p6OtA
1ctFqnIMxDvx+Y28Y1b9cCVuWMgWlnGAsrknpt3Popp2/ALnRi72bkI+J9tX
OeoKRYKIWuo4LMCWJ1qfX6q9tTx8GKsBoEQugIhma8BGICmRxk6I/u9GHThR
Wa4RTriLg/RAmK4GDrCNjEPmVp3oB438zkLExqOU7RuoaKaWucp+6xQzvyrx
2ayKXkdM2w0vRLSeZzW6N1XfwgSY8GbxFGbu1yqkEkuA0sthq0moUuEVaOCM
J+o+e5HyX6qXI9aKHouLH0sXJsipczzUBQ675JWogCkBuKyGEoiGsnU5wrgu
BWnVf0JmAm62SA9l4O6rzcoyAIG6b60kGJCeykx/lMh4czZBdpBcfrlC6JWk
v4KwjcCtJWRnNYX0beC4YGpscfAOp7pElVkkgnlXVVO2/52uyLeClPELTWBJ
tBUPLn/QLSO/wPjL3MsymwiaIRpmx2NTeZlWC9N3VMlZpcrOPcK4GbN1vFFF
zC1LFIxKF55n7tj+2i2l+Yd0cQofobgJglaydcf0tGU9mKqYrkPS8WSR436C
nU0LCp2cn3IVElRpCveRwqt2FP0Bk22+OujJaJ8ny5su9AiMcywY41kfZUYx
LnXEBwtFSXcrYQ/E8Ru+8DSVJ8GAFg4JUxhgTHmbPvINayI9JlcR11Qb28GM
K81iV0iY5zmxUDyip4gThekkpbrvSkirHs9a12cXR95my16yIVbsy23AGRgp
SjH56cbXcUaLNP8rDVqMGLs8IjYO09vO/W4MpKNj/g+tw+IUcAiU5cJqywmt
RGABn5hUWyUHQLN/ard/fSRtE9OYaV+PL/b4Jj55pZUn3ADXfakQGZmc92PM
Y2r9I98lhBibxiazbadYrsVdbWIFHvzZuONRfKIsw6etBZ0K+FmIMqUlAwB5
gGA/HMN0ca9pD5h2IPemAymXSZZhLH2V2liZ0I7HoEa8ec2LNzO5pO4AwPch
dGswbit11d6L1HKrJbnUTbX2fwCaSXK/Ec9WuzLvkrf3rllUcfD63hQjSpYg
xAmAbLsDWjRXvxosfHwmBGvKSK4z3y7w67AvGi8pjVYdPziwS2o7LVLPztd3
ySjaySx9Or4LjIBV2DNcXvNnyfkRjmIgZJwMtxVUJ6nTc/h+1x1KiktzqHmV
m4ZmV+XnKnIOQmWi737q4YIGFZ7m5n/C0yjwQmWr2fHvYddVFEP3ElJpaZOl
5Y1W+dsdxz+Qf26n8cN5EJztM0KKrvBWb0wFOFo2PyH/AW/KMHAx1LFRHzLg
n8oMdyPg4/roIVtF7kTuxM15Pdjy82kCY+wai1x9U+t9wWjCN+QBNmnT/dL3
bo+tQXHAVfR9LzkPbz9TZW2CPAYCPZLTd9cZLPB44uhlsvFiAovgwCMjN8XS
M8RgalbARusWjc2KxTjbzkqMRgPre9ooWYtVmGxehtdzouBG7lP0C0knU4yI
bKSTYTtoeddBAZfFgGIOrAqgSy3r65I5m0qy62ikN2MWM8Azl7avGjHY2EU5
hGcCciGpOuOgE7G77yxwj5qCIMlQbspc7+eV0K4pYRWllF3oKGKiqpVN9VdY
SRQHQhQwyR8hJ4rm9HwL4F9RBTbGdNIlF2UdXWznWHs9ILA0QmOLEKiD9DNy
tofBIuU0+NsK8FNZ1n7SNjgLy6/DA8TshcZAjjPbdofIjzTG4TsEaDoDb668
9QwVYVGW/AaMTsaLKDFUjIBSx9Uy+LQhA5+Ebwd9wm3SF9T8PpH7emfM+8kM
S6BUv/x73TTj7VhP2KDvVv4vWtCshT34KKmRDF+eG3f/rIvrCDUAgtIiTmKp
YUT1K5lay1HzGTZXsZYZhpn93OmMJBJ+fB6It/KWQFgFbRhNAzgRLDp036hy
4fbXPqXLqVjvz8UQ74FODuluWmjUZ22G6yNyM/DOJyTHOCvRvewyp8v4o3tc
K12DUVXFg8FXcEgr2x/Kkpezd64u7loQNEI+RIR4+YJw9jIlZ5ex6FU5qPLi
AUsrKw1cG6h97mMsqLK9WWNvwTUAB2/dQHzhYbaR87ewLNczGSwhbWdWnqZa
RR6XZgFkQp4pP8MmabSut88ZbSi2qXWA5aVKTYOc3ErRpaFWhEvXaCCidE9o
QWO+QkSIr3g0Rbk/AXcSBoEwsqrL0VMF8f4FpzK65RC7Xwgv78Rbcl/COmvd
S+5qw0hgyGPHQT+rKY4IgZAK3IWOy4surr1QsUHPyRki/P+KCu6oSorCS636
9VFCSkqbp0wZ7aN781H9ihjkvP+tkX7kzMnxYxy9arPW3F3yOFcCTwQrDs5i
IQHOkgilnSa5k3PlmHZAVJp6xgE0JalMWZnjYTaXGk7RgBl77T5FaphONZ6i
MYhhLjP9yfW0RvpFbRqOB9VC6YQ5l6HUAe4A8x4452ayeKmfhsn/xJ8Q7iAE
ouoD0xd//aFk1idJN/AIlbs/3moye2vpOxJ7tYUCtu+q2HclXnpbTOONlPit
MvTs6IWDau6WgyOFCR0MAKge5BdkNqrGWIp689g5hsiKaG6XNlweuweTK0bx
rLlkoxe7IMjTkZQJcgPFfDCIPQPnloRJnw1dj2a/iVMXB2ubRhYqLSMmEqbF
CJbJYlrc4dund3KMPiHEq/NKmINcJWNJbUjrhrI+VgiIU4tor/ZZJb1yU0dy
mwOsGgp3L4b+W2yz9XUuOoduYL0py3vW6I6+NKLoeQy8xUQHsOyCCZOxKr2k
A6PG3xy1hUSEcwdNNnVWpy85tTEOV3dVe2sB0+OzHei3fbIfF+0AmAmcoGRI
v7toSyDlWBhjEA9eEpIUGygK4dP3i/m5xuOK73ie4jknyHuiwCwYp7K7yz+h
GEZBHFbZY6D9CY9Gzx+ZaXyPixbBOMJYtGM0bN5wo1MMGFWJFF6n065U32xB
ikEF9itcIpznz6Jvf7U754RK0q3s36vCbDI5pDDNmPwOFWqsJHCCAFdzKgXB
Y0n8bNBdilcyiDILn9ptLHWQ0ZxfWidPND84Q5P5jRUnYrJQE2IskUDL8NyP
hhfUWf2EpluBvwr4QrZBalQKzssXEG7vT0TyjSo/LcRve+FdmxhiFGXOXTpK
DrS7CSoBz7+y/tseJVBryF5LNt16AElzXi74etUH7YjX4Qq9zHWJ9RlrfpmQ
yHD7yThgU+4xSK6zTPi5Pa1R0AUkB+fRTb+sN1H0HGMNy937J/9b4s670PY8
8Wqw3DJScRmZi+3u82I76DwzpmiHVPiiJpCDXq+1g2u0CIX3cUuSaJpv8VBz
kBS0jQ9jzuT4Bken0sh/tEMZW35B6l5WoTc1AcDgYM3deBMhJRatw12zUAbe
y3Oj36IA9Tyn0VS3yKg0LwLagUUt58P2DWA4fRfn2hET7Kmw9aIXb8lQZGbP
2DrkiIXBdFobBp5FdhblhJRGNmhg1iWpmAhXmetZlMBTDup+rybetT5DcQlu
FICQIhK0JNd+IG45C3xhA+B5YqcDC4iIhIhvF2J8zFEEDCsyT68kUCHsLl9c
jc3Dj/NkZcwm1RoGTrvu/d9VHckccNTQZ2nOwzcOsLQ7EcT00BUsVqpULP9A
A3K91uojyqQriBPpKV4YAhuVAldX71tuCQAFKVcrI2Ro/IDhU73xeKPJBbd3
qzhQ9XafBQoBgOF156/DAsH/BgZbuWW8KWHwRxfJYZT97wBt6LK5/g+Ox1sm
dfLy2lPVLzsPQHEhGryz0S75gTf+BrRCrdPPNkEVwM3hP7WgpMkOnnuUKARR
TvF58wWg4MdMoHQVTxCjjstwuXl6/z2uoylVbUlgYR7NSsKHzqL3jXwAB8Fn
RnP5DIepc+oW5Qh1dVWsENwJEq/8TNiWvvmiarDaWFTFtB9UlWvJhYgOis3u
Ikx8EPCdYxXM8WiXgy7BGpUArSXa2i6YxEQYz+WWLVVHlA6J8Wl92TddE2Cn
R9ukfEhhQ+6iGuQsYust7wULxTW0DWA9L9axF8FA6Tq05s+I70RFJm0uvnve
FzED1ktgkKGYYSD3yhSIHb2T/KNwW9Ro88l9rQwB/J6mnSm3qfpaqLB6ebco
JEoqPPKjFhTkTqhZvw3FKXQ/EaUUKM6LDQW5ouFTL7FATaNJ+5KzUTTuM9ro
WX4Pg5mfrmEzcl3GCTQ8zxgvRhdHjVwqSVgjMOywJU6TUoFkl7hup0145yI5
M6mVWUXAHyioRRBWeCtwkcX/CgDHyNLwpNnFxOp1WKFxHYSPLnR7iNdP8kPj
MTzoVzXHQT0uLOlzt0zhE+0Ur1KdqQpzYlD9cK7b1x2wsbgAlTIkoIkC+75G
58LxieQ/MqBwpdWWCAZ+Y/AR1z8WD/ogKv6sg3Vg/aiZfxpyDX/7U6ybpAYM
SSH+rRGwBmcjPqAeDBPp2jjgBoHF0GKo/TSKPpa3OFDG5Cx2k6+geeCSOSug
96CqU8MC+LTg34neG0Az6O/xcxqbACO6X95am0ZOwzSMEAABmNml9OcxuiRg
ooekS2Q9vdnx0yFT/ysYLI0bIPwOeYs07YOSqOYvFLS38k3Q9OPaYycFVDg5
UMpLN5zefVvj8aNaFYslfMEGwSEoeHOF3X072UftpU6XmemahTpjVi99zqEO
zTdeT/B5MBBFettxvoJcWJuoDo0eDMFDAlGoUOr350BP2ZxMxl2WxlPQ9pFV
XNmphQM9cl2iPFLpxCdSv+a+24yFo2RaU+BxfP43bez4lyu3Ud+eWAiVKaY0
3n2RMz7TcD3RHYmif1eOxAgmTKjMHmAWZvzem5/ZY+TTr5EgAj/eQ/IRwyG2
3kBKvH/nMyHuZCGOiMDsyLTNsiY1lBRRtql0hKLIHOAKLZfE2lY02dfGGT3X
d9ZMo9SOC25PynNcQMg0j6I0Km/LYFSiN0qSxvPlzHmzD2wPeKrmEm7hJ4OR
Q26obzfWFSDkZYkXFGCKiEE0IOj5k8g2D5Fuaa2ggEKU4l87KcnIghiMA3bc
KR3ZV6LAfNlUxRUYW0FmDK9CRTFs9rgUOUKPTNYQGfrzaEKf3dXloakaqJ6C
9htiu9C6kNnPsMbxe8+PsmmdBj7n8DkneRGB4ULclm/RtX/M9YJBSTaCU/JD
mz+5N+XwGPI/I0Rm6SwGNo2F+zat4MCiwicj4K1guw32rW6UdJsxoEEw9FR3
b2vGtjgHqADZQADUHI7LO/RdR6IeKSd5Su8CwE61xt5tEkDDU9HaHorWvbNR
e3ZKJ9FsDPtiKdZTyl6e9w3T6HieQFvRgpBbeNbqgUNMjlhP4ORGvDO33STj
o7bZy7r6E8pJAw+BmOZhx/KVcbOrFCcDilMpVTEV4imDDBYJ1Utf43SDxv4z
FaSrTtXSwCDkvhRJe3LdFG6LA7yQpGUPjgXX8mQVuqWDTKqlVFDQH1W8n6M+
rQwrRGxr/dyltbW+PJjM2aWIUQ3RqBjLQsE80vSht7It42nfZ6axTjdvyOJw
vpb2kjDCZDRgnOCDHzlwSZHAxjOSuPrk7/ZquPiiXq19DbOllDJSbkhRUdBI
T8jFpnhjp09lF7RlQG7WyPVQFpN0LMd8OpQECDq+Z91L8xPsWAhiyGbUBegW
+8rCfkbOs4xQ45na1F9pon6N81dhqyWFDS9fjrtQF48mLE3BlSRtVPWxGwGc
ENBh1rki8JW/s2LbGCbXJfroZr5h2rX371WhsknkcT1D/whIsp/8yPppmsVp
N1SX8nPoxtude/qLgHpPyveIWuGqdq7EIyo6eVZk9+vO237rXU9N0cVjTxRg
KJP4u9VaPMkuYvgkHxXHgTJZhkzhTD24Xn7LnhIojBU2jPQm9+nC1e09dxSY
4iGpV/57MMa0ofUBwxMAjUuU86NxBAh0n79sA3reHVnaatvqusGzIroNCBYl
deQg7UVrssdYW+5c/RD5JywP9x+XgyWRT2uxx2+NBoWGn8HMMcZNqBEjElX0
MSS6CZD270ZWCTfSnT9cVok2ObV288d1IVm+qwZdeJsDw/HKQi5mbrhKItMT
83lDPU8sEDaSeVYE6Aw8iFZ7PYBi65+4y1PFQfZEOdhsxmsBb+n0u80mYUqc
pGEIEJH+nbBU90mkz4a+yHLC4jApdXcLC7R4rtLp/ZSyoumqAuAwHcl+xShx
mTnfFXO2GVR3M2FV+pfC/w04uzHNuAb+IYe2XPnlg5EFb3zULL+NR2rEdyn3
Si0K8YlnSoZwPHTC1MO5lAAw0Q2CO/HT3tXTp1+9r0k2rAt+zFXud03q/qr5
EOPt4dTV/Ia7RkmFFZvUpB3AlB5OwCLkA8BYsV62SDGRFVMpZyuOjQE5gfsz
ICZc0SuZfGrF/6p2Wy/b54mP5Tqcdo8Z6Ar1ZTOyRHPMACVn+e/HipD6ADxZ
m3iRVWFOBC5TG29cEc2skghpYYxFQK3pOr9JqaVExnf+M+pw1yXgaj1ksTAR
UYYA748kOyLcyrZrAjs7Hxyk5kkC3OGaN9DoYnWe+gEpIJYSRJlaio0B5Q9R
vdxvFMaq7/V6p+8O5DP3Z5jda2y4oY5ucnkIJo6iuiLDwwhSkmAwdLqvkIJl
tYJWDenlc8+CQGOVgzUS2NrelsW6rtw+B3uZz4sgkN8OddyGYM3LhiDRKKYh
PruYMqXgQaoPSN1sgMHgFlzvFqru7Nczu0OZCbH/UJ97YrBrC5fAbaeF/0sO
5kJ7onpirkm6CLbCA+vSds7t9yaoTToByy9eUhS1RF9PkAVlCZS7bT3djZPt
yo/gAJOlzb+zrR5JVFBSJROkgYSAcwcL6pyS+XJH9SHNoJHJZyGYeI95e1sb
gW8++3JN8ogNedW1oVJof+O1/GhFpi4cBvWrTv8qrhlJlGpA1Gim7VNshBJH
XMklwXdAUwwb3+6nV+nsvUCI1IfYmwlLncoDjRVnioyHZ66Fx+oWZRB8jSEh
HZU0D9caPdTF26q4W5IR42bdBRMB+E1knk6Fn0EUovXjCY9tY6rDJyFEl7TO
ZA4Fxyr0rDwD7HN+XXVADOzdxBRSc+ttmh5JKrLlb+zbqseU8DNn/d/meLDs
GiYl56kzX43yRkrpoX5dG+lhWJQk0H3JdtjS0WaspHFiZUhGERbcylkG/WtX
UiojMWFw4F2IvWVSGxRPC3GqQOtbjku+z/EueyjygwAuTho6o3tkxXjJmMeA
9C1aqjjmVWnMej2EOw+b+d899xFyqMi3+X3Tqr1T0yMGHJihokVQaBgHoMKj
ScBsk9p4jf4djJnYehNmvqZA9S936XDGHfl9Ik/B111eb2KssjRO80+ggoc3
iILgxN01KL//HSNwPbWH2f7cUMe45ms0kaYXIYkJhCbmDxuKNem57nsIFE8j
r73iSBI4mcervZPTpc8Wg932ACtKPUh+0GNNpdNeY2ynLjtl80wSuRClrAwH
9CC49DTPZrrGoThdzuA7a7OoqYVAHGZpod0lzkKr8wa3Fa5/pvGxemFoaRvI
JlTMyYnMpneETfGvbRetuKujIT3pbvtaGTOjuZSO6Txw2KpC1mR50CiVd3uO
ZHIpAz+b+5LqmrqyjsgJedWy3SotkjouWfyfqVv+URW098W3pVM8p0Z+jZ2a
jG9q/UIJsUHo+OOPAbHXq8SDxp5hmrGenng2BL5lkgPhD9VFnrIjVZzVbovz
ioa1rxQ2+ap16vVfnNoqh0SnKTznF9ynRuEAGYcTTC/CjXjNR95aJxlREeMQ
TQiQAf0/zm0jdtkR76EHB0s/g5WsdG17c6jAMXstbyJWA37Kc8BO2ZfYhyAw
SrADmA9i7hQC5g/b4XjGKxFrKwXTQmsnHsS8QGhcMQGBelbvu30Izc4twiiE
cdYY8P+rhIwc7n04sAX8YOZP9MWQ+oQ4bcmTQSljfszG7XGTPv03qaJvMK+L
eRu8OrrXh/1pLY9ESkWLbqC68UslC/R6RhdHpLEVwrqjXlwwhPQzrB7DPike
jXY1svYVzg7xO+pPO1ZRornnhw44mdhGLXTfQPSSvDAhk7lSJiV2Widy2nVe
SJGmoygvWytOLnEPKNR0fDvD7lZbLivMD9Gpcw/KtqcUB+hkQD3k8vlQYRFG
RhA9gk9yrcLtAcPUZBkvjf5ibZaTA7IhoS5ni/cxnZDZn2TjRPHmTz1bNjRH
F9PDiwQh3P7CSEoi1WfkLRukmnChOR3x1HrIbnOy/q8e+L+ke61KwxtsRUio
P8LRFEMGxntmJlehHLWI+DcaKL45pCJKsrkLuRbK6qGNaIJhrG7iQ+Gh/bbw
H2GdaLh6Ic9q5mwL7vdCZNeYdUqH383R0gCH6f0peDq1ESjAtmYD0aM4erXB
+131blx7Sy1fFB33qHhxyoE983oXEtXLh3ccS0VsdQQT+78HDVa2veAa03dP
wY1vd8d6pC01LDolVk7921XrARFEyZXpNAQzaD7s0iPio9ldvtA/uCm87Uci
Evd1D+Srb6HK3odOB19hK+TuYe+D/orlYDt5KO/ReyoKsXQj0NrWqomRaEWc
z9+Utms+0wZ3g78xii3UeEESJDgtEm9n1B/2WgDFawmNQsWqCM9Re7SuAUBb
3QMo23tCHsLdvjXTvSGKvEILJAiJDYkrjoK++m53reoya98LgNHfkAVnUal4
1ZgyJdxR8hPNvng2j1EQxTVqluItW9PlT1t2UT7z/2yNOwtBTh0tjRZvKQGi
R1gBctGM1LC0xPlHER2He3H+yHZXlmgXT9MBImxYv2GCSaqk+I+EcYjUkHpW
kNg84eRFd1460q9dzPMRpsr5Ozm6gjWFsBoyA3jbWz4YZKv5ni15ZvGXaoeK
HRzyDRUx0gSNULY0g3KDDUwyXm+iUtaMzfWwH+YMVZmiNLzeJfZeSK0+KD4g
pHuT5+cv4KAB/bz3CaQNQaxT7hEsrA4chGBd9Og2EPVZ3Eu8mXDadbNFkgQm
rKXm7gHXV4EqkIhd01cjLH9Z9dSLKWA9kIQ7WuQOFOXEDVvPs5mGRzDeXMmo
zQNocxiZowGByf8hiiZm+5lUtcS5or0Tt6og9qyjouRZaAwAdU465PPLcook
mnbhZXVhxkRcfS9WZvaUdNmZbbbY0PzZ97xfzFPWVZsLFsKTbXWgTtoUC1dI
8BQkjY1FfFKtH7UzVlZRXYP+I2B1bJ8O8kPFPt3inH9SXU06tbPzjlDp/WQC
icj0KC+SEp+ERLEYQI56cz2qlPX7nwN+BVeZCwIUR7sLLvKoBFlItszM82Cs
PH3SIYcVEfhwnCk9ywbo69z4hbpd1ZyvPdjV79i8QsMWKO1Q2eb4Zj52vq/x
JHD5Scvgcxv1R9AhWjWNAfXnW3WFvjlqj0LN0vEp1RRO53u61xvPjNDfajrn
MsLYvmsLj4UYP8rBPYUt+4VoOOdV2GJ/HPUP6l9oQtkB0DvueFyK6I2FDp90
eSHQ3hV6sdINrDt8+fWCoTWiCyC2Mvs/Bvpz8qfe0ROMu9NuNu2vKP+vvhzR
8pRR+xOmON23tLQJXBpzSyLVPPoto5f3NP/YFY0LNbP7Fd8u68/JCbWFng+5
9OuiVdRItH7PMipD2YdXdOXIvMzTKrTbUZNwjC43JVQ6QnTbgYp6j1hoQnUz
paLLYhVs3dXI3PSF0BsKO6RrPTG3QzZbG9/SeSsPWOqSLk1jN+jz6o2nGD/s
MpiNMSWE9mGV89WNaMvZdaHB6AOBKZ3EVTLUGz+xcSQDp4EymjM5q9nwoipw
orB8eU0TbfZpvk6bP1vRYIoHE69IBWDIUpek8WfJNXcj7o6X5x8pX4RSSGQI
pRYHbEi+0AhIVsw8VrhEI/z6kAfjk/MaZ1eiHeQ7xArQRt5CTjkx7hwVfA5b
JkBUPSbhshbhV/y8PvLo7JFefLBy6e282VXPqFGXlBDNB/+qYuWHYcNY0xAe
4rZXOwxLnBtqygDKVpnDl2tmm/utlVl9aWLuHV1EBk86bZtAFtCGjMgemOAj
NVX/J0Ib5kAK1383FHu+aH3dvev3YH3wqqw3OqlyXpJtAMXBEN0dVnVvcBCF
MmlGnXHUp0qV/UyXKNMl0RomyidBX8InxPBd+1Ci5j3JB3C260QCj4waAIZc
IbZmNfrvb9OLqsAtNdCGRofUpE53A/kHaHbOP2hwTf9Ascwhiowbfrwx2iaJ
PRJ5g+bIJW47XaBQUDWDVjF5wrmtkyLn1aOuMyqk3C0OBaIQOFJbgOy4qQiJ
2MhoILlLtOtpZnKQPPsoM8/q+lJo3Yn7FKObT16MXgYv5iE5H5RUQ2V9+JNC
I8Fs/QrNFqPtnQRZhtQTrgjoA0kKaFEpAdjtjOFm+FrUbbg7nha/guLr2bFJ
x/wnXI/pKzat0ia6o0txFKcfz3GAm8FbYZ7VW9XGDIOCDf7hjIyDDOAM2DRV
4RZnJM5ueEQ0XhhYuTa9jec2h//8/IYwS/Mg64hCs1qIgK5yPRmktmWsae8b
5JMvlynj5uHqW6iOkYVJvJ+e4H2KwfiZmMMS1HY5KNdY7wuBHjCOlMm5kKyA
W/stfAYyYLS0PSO7dvSPGJn6BnMbxCSOb+oq4/2iBvoqR8np+Xalzy4tTUBo
InJMvV8Fa2WVGLHpOE65KGpiW5y6Jtvhpf0ZKQhKoZQ4y0Jy0DtquO1MVY41
4auKfQnkASG22bNNBihXdXwRVQTf/etYhFLcUgWN5pvLKdpLL3d6Kjp32eOG
vtx9p38EQ1wF3R/LEJ3LWTCrrIT15aRwp0mOc3tUHNxUTIjlBbW8XgE0ecJ+
zvAUvYXDb4z31t3RE3HAP7isZ7WW+DphqYL/4k6cLsOG1DNc3fZVnA3+YJOL
NZdwfTf4zv6rfAeGMQxgmdCAUw9B8Mq2ceAo+roDa0DPfeQlC5NqhuYP78/Q
lkv/sqskLKO3HFRNsxdimeQbwgM+ge8EFOL6Rmejf92Jczjw5sKNfQ9FBj5E
jso+51quKTP1mp4X09xPV7Q5QdBZWQk9JXAGxtWeFZHJSvIChVF1ugudkiS6
cKlxEnl4Y1xua34tMaOdYibtwpgU5YWKHfWyR30UWpwIMfuSH9hzMNp4byrP
q0j8L16gBS3TX4y0Nz/nKxCOyExSFnr6aFnMSWo/BoiWgpsN5P+uf93YZ0tJ
kOZRKIei/xP8aav8dET5bHgRdr/evxDqtttcS+qc1u04G4BPdIppmZFFLLBm
gPbQbkSa2pil4Yi1rOe9ggFcZ7+DCnao870s7xop8lobGlrdSml/ZN1CdHso
wel0Amhhczxw8bGqvDXEicvSabpeVMUJWP2v836iOfRbTTSGFrS0Yhzhoahj
Qj6/r2AaDWgbxaPZ481Np4GHrFaSEgoS9WH1JKA2Zv3lD/d1v/ZrrDu1Jt9R
UXVskxQvJn7rQBCX6CwPYccaeXZ333I3364/qO7AzNJFGa5wa5Dx2NLKM1k7
aCyIouKopa8jkJm1PKAW8h/G/vbpJ2Sd0WwMjClFL4lN2QA9s91u2hFtvtQY
E0HTO98BAtUtEscZe0vf81wZcoOhnbOOyEKIXkGHkiohZGEUcoi4yq2KLN/1
gY/9ASc82nWkyOOuaSaAa38UCQeHjHY+lFhwGazsT4s7dpgBR8zgZhYKQq53
RE2TQnOauO2XK4zHiPnLH76Y9y1AtQtodVQ3ZlyrwwxGrdFo5ypjSuqRlKmF
QSAPWLJ8sLhzRLSzjJqk1AaZNSzbFPfMCUV9PROn7TQKpUBKlkyduG3yB83k
e3Gi3OSG0kLXEKy7hbysgzffUW7mDpKri6kEOwjruEhy1kLJc1l7wTX9tR+0
aDRS6L5i7VAYdLrr36pGbcMWDDHR408B08CnkT1gkewnWSD0EHVDJJDoqVIP
V5V3EfIKLhXLER87JJdojEUWzroRJ5kPjSqrL9Qw4MLw3Edo5t6h8C3VqDxK
PEfOWWKPXRPwG2jdSaYQ/4brvHZpMjzQXzX0gFOU4IQucZRhD1RHd1Pp8wuF
VllkqTrcPdAZM2bnyVmiWYeGXZVc7inNijPTEZ1u06Ohj6TQ3W+2UaKt/mBv
StJ/kEdt5h9rWN5TTpzLwwXJCjXH4u4fHq0H/+r84bwp+nVzFCRYn24BR8zK
U3W9HlWIP8soYL6rfbtqPNNOf4ClV1xQfEsRDoVRxIPB7gkjBfPh3o+1zxFS
QHFv4zt0cU30m2imFyvwchiy6ORMz9Rb/VUqQ8JpEsvC6dwYAc3JBiS5q2A+
jziSJ6kQoDGYLj1Fjo5I+t1WtyQG/Bb2xOsdca30BpptNSqZiF0tiK3KxTxi
Ci7YdGVrUJzCq58BXhLfV7e18s46dihvOhuMSkZfaKvsNzQr/wuR12EVHL4d
MNtyOY9iA38j5/XE6Q6z18VCVragGzQKbQ5XhAIHkfqL08txnUZXzfB4tvsi
+XFdhuK62uaqDjCsk6p+7NKs7rENFvGqdzo9VjzjSkpFvhCb2MFvabIyzEw3
VtmtzA3DPAsbORxk/ReNaDNwgtqbVoIAx8/xRRunOz8kSfE9gTLDiR0uxnmw
wOChIrIFNTNh0zxDv2iWOr3U/ChceaZP++M3vRei1BMgP8y635QZfTcNuUtk
7xdwz2WHdZn19YaybvwY7zGDTE/hIOaz0nL3u314LUf9Zfd6+BgbL0NIngor
RdszOE7ABhwTbYSnjHM016R4h0rUmSmpWi7UNSnyMATK/53chFdmThfZi7GY
bD7Od4n1Z8T8RKCg21+LP2FhjHVGKIPAdl5dRng4CpnygyjQp/dnM82dc66E
7+7naqvwe+XIukVBaHdYwfmYiG3P7Qdt0rzRiCIzE3Fzs5cvEDc05ItFfehS
hUQmJdIlRSn1Y0yd+avuN5QRtTJsT8rcow/SrEFZarKkuNQqW0HyIBauXOxI
W40rUlmZoibuYW6bmnKhma2e/6Igp6XuTeZKDn2rH0roK0C6v/PbAmlqW3DB
dc4tIdqCGVtEb2L6DfzKb0Xuvf96WBLOSWeeEPEqKCNGMwHpVXBzVKQUIHL2
WmNp1uwZOW0caV4zS+DWWePMXDG9C2cAcj0gja3ukkKBz71vKxrU2YrdaRsi
piXH31S+qOdyAUdC4ZYYG0/7fBsU6BMuOWQBub5EQzDjNO5/pIlz1GVKnFJA
g+Nkutedkuqk3ADeS5y0x/tIKGscRD9KuRlEvzUvlCf3jOqKJ2S6p209AKNW
4SuAtUAPm9nRC3OQG7yjdfdjUOIPs+0VwoP8vY1DasIRV+RC8DOUkD0zGXdN
l/4cGLOys+JkXLU1YguihniJXGdogICvXE0YdOWfGK3QV/pwxKEdnYBOIhsj
Cpfi9il3Fdd5Wdnf8IKhKip8CD2czzO47goVjsminVPS9HYLAZZjGNLbAlIc
yp8YBpZvH6whtxZrg2mJ0EgWtohOQrmF+gOo005OQW3EgeWnNGKX31iKuf7d
OI5lnFXIz3AU4XsEPwhoe2h2/F8kn/uGa8FmynVwxkPeh1ZG62AV0Yo5BF3k
9Y1o+inUdZjwQxxAnggUiDZlowdVYuKMpivwVnMqqLfyw35M1RKTcZHbCLto
LxiUDIXYAlAuLbUn5z+YAFzGk3wdLVIz4uL2GMQ8YnFq3JXb/+FsxgKGZ6oO
Wel9+rtELDLa+Rd6Gm4XQwYjs+dpcfCgCtd3HlTTZJBpmccpk3ElQsHs/R0p
cDX+0/Pxm3JjENfiopizxdhotJtUvOVjkYEKcApFU0S1Gt66o2O8V8p8sIAX
MIx6pzGSKw0dED+baOjYj6iOFllCQDJL2/HBp/m4na9Hp6LXzhiKUqP9UMHM
EuCPck1nm2gU5EEl/aZREQqAe5+mPOabMa6iIDWkjv6d4YSZbyMBbB/c56Z/
RuPa2Yesscw5RyW7XFOK7lHlM2IXofC338VQe/6Rxzc7nQYj75TdklQXTl1E
h1Fb0BuRiDoIdjCKdxlcE28PnDjJGa+rNOXQX652tAYwEoW69a/p1lr40oty
VaV8NyheitmqxCB2Bq9r/VFAWsuf3xbf2TdPY6dza7+JXa8MV/gd7WF47aW+
Gw3gB1EK5Enxyt1N9COEYOCll+Gb8p7q4VGlcLd2hsDvPqwzCt9bRxkJuz/Z
rxjRy6JzF6/QlgUN8DpKsoWE0VLUTzp0b9ujYg2w6u5jnOrxtLSAYDgCHWGu
mAcOAr+WnESwqUo/8WO8bXmHW1cWfK9yMNhZOqDN7rT0zUxy+qO1UIrWeD38
l63FvJRdBPs3kIqwAmet+LKDN9mZepLNrqXqMKG8yLZGlID8Z4qK3VBYBzZZ
11ENg+zEVleXgQzccjK5cy5ud3dVSoJowlUnM7PMBB1WhnkNk1+7dUe2Ohab
q4k5CvgJy4WJuFeDWjikuU8s+RxNahiNBzFXmzUYnWwIII3GHCJO9ZTS2DyV
QO9oSF2d/XwqSvTWjexNmAlrLCq+ovgXLH981N7UR6/FGC0dQxd7FzH6IHt2
Nyr62Ytnr+Zu77T6lGlBXKSg/UieKBygPtqkvoc8IdwhZn8qhoMOVZYClxJD
4C7BLqnuwMP/n4ZN7hFo0pP3mH0H7b+yYOHzl3XS5DSwOKI+weiskKB/u8Gt
EXZPNlpAaru60dt74pme3WMZ0YUkD5PWh4WyCbMeoniNYiueuLBPGY8N11UC
sI11T0ENA2RpgGJ/dbusjaVEYBQD43u9fILtdgs9eCb/Uywge3JL0P9yLoyg
mbifNHCm2sY0NXwJRkL12zzuX+tXuo83p5/2O1jB/JyFKgOsHgCWxCWU7Q/n
9FgVgmYofDJ5zDZ/VL9NBIamb5IN3kpOL8ZRT7Opb/69Bx04BjtpKSRnVjII
Q2Q5/nwYFgZ0Ecw9y+NCVUPEn4QSJF+yzJ9S3YhxtBA1rCzkOfNe8ekbfj6x
gjePR/Hjc/D+xq6eDjhfRYxGZpFb5smklOQqYRkq38wY9wSu9j2aPFcSx2Uw
jBLPlP9xo95kL7maBQgB+a/u5vyWa2hnCvfGYvTNZpPvyW4f100B6oizPxi0
Th626wSixi4ws3M73UtqHMgVtKO/TtzUW4MN5OMleRqBVTYNomwpjFfAULn+
oGyjcypvHp8NVMqN/n1DOHRpXUmMxm7kSzoHVDL4TbptWkwMr3KRAdn5d5p+
yspAJKjd/YYWFxLCyd97nvP/EFdIbR7JASdFeMhBZ2IeALVYwjLSjxj0t442
z55X6brVJgBQbS3ez5JPUfLw4Z7t48JtljXZmZrsk+sLLqmZaF+yjBXLje1w
/k+De/omLHmS4OztWzUmjup+MxU2pRAlhnCXpPi7RERMlSmhtCycjXvqzcsC
UWHYcCesC4BYILmDL9bM3xNUQB16D4M+/0gjjYPlRAOl4dsmKklG+S6DEgWV
pUolcLSz+fhcqF1yEf91l2EDxLX6q7Y1iLcBxgP86wGDBZKKi4+Eg5HDeBTy
TOufpgqELqjKiuSkb0BN5+z50oMmdCog4R1UIxKKqC3vffAj4Cz0aqMj3QgF
YL9gtd8ICSPof5tYM3Kt+EE0VBRZ3A9jNQbicHSfnPD3wg9jCq0nY03BDIFq
G9MRNpS4YPi/Wa+14Dd8lOc3r5PwvuvVrZj+1WityNQ45vwR5Z6rohcLcQbw
vWByZfgB7H2w99oHnH7wUcTA/ESmRdVRdhTgGxODyQqqfK9zdtGoDqhoneOO
sYeTZDsyfe/6qMAYl1yCcDoxUwnOhuOL3ggJ8NJHlYJ06tNgNg2PhrsqxLn2
UVYdSCoVjM/JYBOkZWAlZ69xLqaVLm68RI1O1MLxRHHIvrMju/fJCFCv4OeE
6x9jYMstFt3KggYELVxIQ6U3JHM7EEu0e619MWGtXUnrv0VCWFFY+9D+gNr8
htdpUIrOiVpi8galSUIHslqQ4fxG2MugPpvjAM14ToERrqiFM6N6+M3M2Rz1
vPJGADcsgJgUgS0mL6Sv9bpn0hQvyF+Q2BJ1bAJl5cII6Dzr4ssmouR4i6EG
Rnjy8dMxK9a4GbC8ESkyXlfb1DViBDLtJx49cd8+EFsq2DhZ39AThWoev/zy
qqHtVxyIsfG1Bn3FeOabe/mylnxQQ4+zgBGOPo2CQ8UNr5AzoU/5uVRXfIbP
XNHdFz01dwtwbntvUD8IltyxO8NaiHgPrXHfGe+vPBWrjRk2WBTlZBz9Tp3a
h42z+RLQYZ7s9fqNNRIKiQ2h2AV7qLaDIlyZ2VhILArIGlTg0quy8qJLsU6G
hBHPsiVsYmgsx4Bzd9aIPpHpCuobKiWGLmS58OSUAM/q30FjPUW1XGkTTzmB
jVZ4LtPc9H1bnYm91eNBa27kJwnMOxtMYxHpKd60KatoBniBfXz9ZpRjM22L
5Dv+4fmRkUIYjlanppf9XxZbAQ5hOL1+x7QvHLE60Ty1PPSgrVY71klQlCyJ
uroLZC7/dvpJcWzYfmUGtqy+zcyqgx33qZxsVCP+8MLy1XRUx62CuilJJ+Dk
zXgzFQSss/CDDOFVbl/Z2glHeffOLqufaj1gFLURY6BCBUu/v7Oen9kJkhDm
7m+aQ+aNDGaR2I26aSXbnBbz3wjiZv0cE6FamZMlTvWp/Po1hThUzQO2qVTQ
62tlUuBKQ+Eprrv24dusTAuw5UQ1Y+w0wrLTbEuIEKH2EPKnXaa1CeRYkwrx
/VA5DNlmGxlmPtbxxkBbTVuRoSdGpgN6JDlRawvTqwzm752ZU9u4bNZiMdjH
0YVvd6vp5XeAMi6Xb3HYdFBBB/n+InuCMi9rmnNAsRGtMvoEQyWcKt/mbOCs
OEu3jrET7TRlx3qynA6oOn5OqfRvomvXoU7qmsn6wje1eWZp0d373DuvBcae
rX6xBAE7Q9m6h/K81U3ZcSxjbpzGKsufn3W44Cfa7Fbz0YDl0MkhSxfxrCMW
1WcFowInfQb3bzbCY9KSt3JubhX4Cp4iSH69XrKWfVimTsU52ttuLqXjgm3i
7TC0zDyHW/RCpxZKtAxNX5of7c+ehOUiu7NG8MPDxY9dfXnPCPQ5GaUSqFGU
Jff73ZHeRwoZw+bZ+qYrt8d2E0l6QRbDZNi9I/QywYGzTd02G0I8sl/Y8YVP
Dy1obs19l3tD8622KC+/h6IVs18092prKag7oPuBuIzdvR/RlCgCs18lQFPf
vcouSh7OWMm3qwriVkBFM2CqC4/TYWrRUtYaBcJV2gBjk7SXbt3ZuBje7zJA
G6crjbMKklEPUpzdUg4Ulh9LSw3LndxIGSNBCyffcUXhIZtTADbfyqWwsLsC
0P3wfDgjGEus79zjftyI+PnzZ4iKrEX9wob/fISR+xvoFCZPWMm8wzNVm9CV
gHwD+bcAbUc7/PM+34AfnX3zh49pYZ+/rrLjBXNMWzuVcDBVppneT79A4V4k
FgMirvS2YJp15mv0x2payb9EfSV2HhdS+VlYeo1Cr4bO4zYDKJG/LoD9aDU0
5dJCAEBmCy+8ypWsNAutSLdZyeZNQUsJb71yzz9BGnYOGWoXNTRFAbMhPrSI
obDgArvJflVIX9fGh/8nY53EIxlprIpo6fKi1Y8xhSu448HnTTCKH7IE+xZm
vCiDRqhSK1V6zdjdgZrEXiDmdk5pF06gCal1ZXJZzdt2itQrpg3bG3tvJNj4
VAnDgC+ZmEOA+rYyWdqmLux7aldAnuyGtdSZ4T2ag3hMZo8mZp+crH7Mg56U
uqHj8InJb8qaARlXXdmU05w+gN/8p25pRBNMC/pRxG1Tqw2Wks8atGcUkxO9
qC/+sjY5tVwvDsyi1XU2sBiDlttcoM7FgT76+nCdDqcVnTmc/ngqXl59Xcdc
V//2HXci1pXtdfP3IphZnEgFg2e8Udb6IsNFAScmoZK7popW7aK2ilBctNk0
Ui3g2ngn8s9hLB/wccVRgx9mehNpegQ3HVvyMpkVxxc9ne7LywJh3Xr3CxY+
mpp8WFVxrDYMb0xddcjWg8NBKyAekzLp0NE1m0uPlOgsgLPafDTP7eOeWVS6
T1Jy26ufMC53o2C46UhtjED5XjVeNkKNwFX1o+cu687zF5Hoz8gyMedoxA39
sBGY/CENduitS0CeczqkNHLhN1o+C74erC5Ch9T+RYtLM6TgOA7gC1mazDgW
vqgZxKi7nvJTn2HKxDJyPKLDZCwJG1OAErukAiVuNFtF6YG89BSbWsahu0bT
Iwi7oYJJy+Wrj4YVgq0mwERKGYvSmI5btyNMkP77VqsDX42UdEKO9XKGtKxx
eca0OqUx9lMX5zTXbj7ngqkK/9fPg27b+C3Vgph1WSkIMDbXUMUpww7ajuAH
1O0ZR+WKlZhZZvGIHIGYwPUJULuHmyE9bR9zYHtTOVuB9UdJSpS5ioK4fT0V
kFMhHyN9lP7Oy0HH1g86XsZNKaCHRwpv7xrE/zZ974KOrL5pIMzOzjG2TBoN
fIxAiwqWuDfrjCpdNRY5S5/+0VFel3pvFuvB9V/AbLPFX1czko5w6JbWbWyr
sMTPiuhi82dQqjGFirxZxSR225+kkVsPpdyYLcxxBv9PsXERtcie0oTg41rT
Qk9ZC04pavGG77RKvxFi20kXXS1W840+9wJV+1T5FdzhQZhZdDjGQrcv5mE7
fU6vwJyNp5valWZQINxQ+aAtujx6bRSBH+3+25w4Gg4h1iScyfpRxKLq6wYM
Q2S5+RNLx51HaHwK99VVKbS+F+FeCfTkEzX9aFLV8yTHpC95kL9sg6tRG9JM
Xe1T3cAH/saEVRShDvl4F+QIYJk6Heh5UsNQzFztVJdM46X44/B28G0S7YgX
nyNGhujtn/vTMAI/nwwsLulzXuuGETFqY6KaoiNTR9efV/SfNYfgbiqAQR4z
nx8hMsr9i1wGo2q98E4nS/XLvGRj61tD/OvU/d/M3q4YPonowCuzFWiXkVTT
lcFqbgDBiptBtoy+NDxnjisPeEXIF2xiXGpqnZoX6ISqeQT7/J0yrRWyh4Im
1L8Kr7Yrimn8HKTcK7Deskm2/6G7MO7tqhxXUx5GRLjJspzjFpZC2V36/tvw
UP40HneKyW+xxvHLGs+uw4CBP9HtJRWY81XoWRsmzMF7kJBvhWHwR3LhwfJV
oAr2pf2mB8khdK9DkLf9C4ofq9yviXmDeddVwTBuwjj3n30OMlNkwXgWLv7N
Fp5TVgDmaupsOSfpmuVjFcqmeEOeoBrnZD9BrLSTTAnkuV7NxfLNf/CcL4OP
nVrerIMn88afgYsOtjFMdLjVFSteuZ6h/D/JXcs/uKla1RD2gFIX98kbraze
kzn6hNIJ+NGbCoqgeVzvGHRRh6xWe59Tg2h9CrKjv1QC153B8/ok9b3CFFgx
QEhgqwVDV5NFzlL7us7qITd8HEHvXBXVt2e9uBEHd7XDtbIYFrB5jEX2i7Em
6RQc4dB0G0ufLijA79jjcIt4quuXGj6PRdiF/3bG9OSrlePeVMOlAbW0+QBy
PK2Y1vDAOFb9dAJ5OkrrOE82Z1IlOvs7NH80Ssgp6DBCCKa3MocbEfEAiFez
U184pfSTB35tPQahp5Ow/HdI4WVjYVFVvZBBaQWLry6Kr6uJKaLVvGZiAT7C
DJH6YPb/uf7gaJfYq2V3jYRjfr2F8Mq/9fFXS5QfjluvHUh8NuW16ZNFu/1C
rqXTQRqkZQg5s/k3HVtsMPI6HZmEG7NTyBOxbJFAviS6XtlfD2dxsNkco4Bw
gpXmYtEg6KZNz+kjZPyuJP3BDU7rP8JpNsKZyOc0Y6g31ypcYmPFMIfrM/rS
9vQeZfz7N8l0oeo43jmvtmOChIaJHhbEXWYnNrAsWv9YOh5khbceoF30+RUt
FZLn7e9BhGL2FBJoKPaXUoyNguzymIUAekpzNrkt9Usx5RhV/16c16GjN+dV
4MD97awq8WnOWSVIbHhzqWVv2OEGk6OZEVV8v6G1k5Xi3R06uiLVHt6Y4339
m4Dkn1UFW4vVGS5XHTk7XYsbvwdCDBO7pl+005X++pkNShwQbqX6EFqbgnnB
4tGRhHNguF9+CIzklkvkZygbAal8pv/u6fwROa6MmgW38Q1UshdEnCLZLEYk
1sbMDCC3ERk7TiuXqvn+i4JqpeahytT+FhEt2I6vXrSUwjkGDima5ycngMgc
rgzneS9THp5FX6oCKdzBlyR6QGnQ6MfK7yVLGm8ww1uJ2Qv/538ii/eqNcjO
U0YPPuHgw5ECuxwgjSZ+s2uChvUTu8eVzdFERhauo8+mT1cg7LbmbIbHKZnu
E9lyrkYGmMYM+DOQOJxJYcmyOOF9sqJqhIoiWgs57QhvAj7aiuQrEi8aEvo+
NHfIVgZw0fgJeP7N8Ly1YIgP9Vt/MlhsXwBsJ77cn5yb7gJxUhqwvdma/VWu
JGArEin8/1u5TrdjX6q809ZVCfd3o+vQmkf9L598Nbe3o7NYXsj4P/pnODLk
ygtjIDDw2RIGM5DAzp5FspOadGAEj6qKgpkp4VQAOXnOfIDUc/mBcTsCOT/5
cXU+pJvmr08v75MUB+qgoY0nRGid5S+kf4L04uHPIbkxNrT+pJxWTZRsefMG
30hD5qB3prJBn6r3GE53KEPAL3y6yz29I0uvc8o66p2Khjnovoa+a4L8yskh
gJu27wjH7KDCWnJxa+X1L9i05uBf+ccOk695M50iC1YWlrmjDZkB60MWg2Y7
SrumIwDT9+IoFsynVdQL1IELIRzcT0yh5iGNEhYgCTJXP0nwyBoFKXGhsyDF
/rlOpWwn0gNb8+zUw4KsFG3TOhtiJe3gwZudxCBN90x1AUqC2MmgfJBKZEvO
cL3LhJ3NvIn1mJZGfE+kES0KQQUzyp0KJvpFCEIKr+GhGmRLo0C/X0hZv6PY
v1FieUlpC4niPHMFDn1G3GQaewhE7lal9IEC8IiwaXRDuhcPmG+9flGiM0SS
QNKJuCMhvvCQ/PqXyrHInRRQx/u1gz7JBOuWdbmEbRlEAt6tEIfKy9vo8qQ1
AZ6H2UjvDWE/8M3GA2OMoetMu+HolZcjVoSVLnVoSHfMRnvT56uAAf0DD5Lp
1zCHhtzXQU0Wur2WadaPOXSClBDfG5Rvl9BTzeSXtlXTiAxUFtcNG+/NMy5D
UVLN8SX+oJkJLsGsdDKnAL3TLEntjTUCOIiWHj7xUILbPbGl5WxHEysgwYDd
jy6QCD/Qv6RJOGKjPRDuZPr5cyG7iOejLztyXxum2KXN7771Ic2ID+Liy7yg
8H4+X79w7XKtAWWkuOjPzJoHAJ9idcJc+TBXUJmPRqsddmgQlZn5oaErq/0A
H5PBAf8KnNmZnZ5NMVTEXimk4o66C4TTsxW89D70WIDhIMrdJBwnKTwwrgBG
MEoNZPOAOu9JqtJEfTt6mzNdW5KR3sHoDUZg/WxSuhvo4hwopVkV+qVKe8g6
aeAJWqRgB/FYelpNpAGITZ6N3rZqghao/8n3dtmE5Yoj2KEvko+anQwuITwI
vypBkaiyMHUoq+Nxfsk3LZozTa36Ze3P7nBuvp+FJ9VHFOoe91Zf8X3Xjt17
XC9TWpgj2eZhKRb/VR1ZfJezFQwGYJLc7cHp8HRr2K+PhT7F6LzAPcPlyLLO
ahIqlgqXSyww5shz6DVT3dR7fZwlZcbtID6g5+34aAZHr7yrzNyOphQTmdXJ
La04TR91dujRVHb+/65BQDdMKDzCy94r7x+OYakelKvJNtcOMJs/gEyHdUkr
qWf0PyY8WABRfZEovXgEEhiKmB91hQ0d/FlA99oInC5yFPvEt8PGbrh6+DDF
NTEhSusWyjjMtRLI/vknwvoFhY3nljRCJJzZk+fr73cLiwyNperIBC3c6OG4
dpprkJM2N4gIjj5VseQyJFG8PSZmZ6jcsq42R3KBkqGlT/7fEpB+R2aE71x1
BDXnic+7K9kZ9Ej4tDf3UTvQ39otMSOhqUwfPoCPqvaAcF/XJtEt/V+Eg8oq
NAW8n8VK3cc7ocdrR5SeCScyjao+Vm7y818eSnhrc0DgGNBjNuH0XrqjAuCu
gluzJ69bLRbkv2dSeupEK40sgfrZsOGyDjGXdzUXX9XcbF/AXpCw/alC7iWu
JsXq1MMO/WaJPQrN/qTFD4Vrp7WIBC5Ej/m+nfCJ5+GEJVah+uf7MDzEo8yX
30fa9ZHX2V/IzAgzuRCfCg9m4WFlw02nx4w0l4iAC+9fiQW7Mg3k9y/37Xjb
sBrxzqMEr2qblrmhyvOJevXP4JNCjqeCfqzZ69rw1oA+MZUrpcxXuOCkt/Go
KOakoZ02K3BwGvNK8ohsB9t58heKGANEAxBUHkU1gfKFPmKEW+kbprifMZa/
7gfj+e59FuThc/Mt5fs+D+Rgn1yysBHOFTTxt06ThOPiBV1lKqRYkh3qm4bu
kBfJkVpTrjSteVHPtAi1Gs13MB9F90WbndFhxcrKQqGrOrk+MzuOM90fHUeN
HmiJ2jImBGaShQ0AxXyRzjBgV1uIqVo8h0IPihZGqip2GiIVd9fwh8s/4XkI
e3QZNL+Bar/42rlTYHqCJGZAbks90WgOWrnCoGoowFeSDdAgkkrb7IYA+a4J
nzQ+7ZHZlq1YOB6S9KvSMfmL1hPaqNNsoh4vjkXhFlwsGFeNZvHQzO71n3K/
SRtRyVpkkKLA6Xw1Yb81k8Mk0wifK0aQCOCSiXQkrCkAsstSXYIpr/ZKKCTF
Mt2kVdgXvrkAoBDrQYadQCZLtrOBSPIK72bn3WTBP7o8QqnEoo7J+cFo5ARX
FjKPhi6oNmURdF6/mzDuNivLrlILUcxRbqFBXJnGoZrgeFUkJlSSRLiB5eOQ
6t2b/HM9/HdknpX69yKpwB1jtbY4XzMTxp15TV0khJqlIDiQ+JjMShVuP6si
Nv0yncUi/7qnocM/5kRWNVy4zWFrCAtjL7J7e+1GIYxQ7gA6a5fHZyH+M143
/nM0NvXQ0sfZ0vXsrK+OKvkQYkVFpQB9PFvC8WK7rQrQKNDQlEsVvH8Izn14
KCHE2aJk47InUtW43I+AJFHQsgdqSW3YBwWj7phykcug9ak8jCdLjNeQ8mvz
atw2UU131e/Jvwh+kLaAPlwbKs+xMB/Xy0QnfZuRWQn9hMhPnQshazVZE5lO
tK44jlk6hilHKg1ul5CH9Rk7bBLbHWV/COwZVXUBxQvMY374xqdKpYaN5LC6
H/SeAsutDliFkGnx5rUbvH+zxhmLZV5fQPEpA5EbBMrdNBcv0k4vXIEE77j2
4sX0DONS9MspCsBWMvQy8+lgZBDeCJBdn6aABysD+yc7h9j3LlLeXlFHEARp
VVt5WRZ9pIZZIaATfnnDjctslKk6P+KUJW9AgXsJ7qvFNQCJC2RsVaCNc+vT
EdqjcqaOwq06dxdDxdQhOU23GUcH4TAe9dXKUdtLAei8FmilS88qXPWwJrxq
2WFbavjMjFx1zXsS7DYH46youPQWZ0KWHFkZj0wPjpoMuookOL7LvsNhkQ66
6nHbBrqVmAxtoWogZCuERr2TAd1WaAFH0c8VlYoA0MZYv2q7JyDR21MguMrL
85u+QnL0KyFhigijADEylvUQ6akyhvbrgUDfX8tV+xYnzg1+yRtzOX9Cmmcd
V5urhzoDL9lmonasuItfChldjtSWoENQJMBSIdOUKnXdbGzNOjlibbfFA27T
2bkQOR9MdQmOnmPtlTJXYQ42YPKqf10SWn53RrsfMs705HBxgd6Uib15b5g8
qbrmyOjjh+OKJjVRvAbFkjwgChB0/mRbp6CW7poYQg64qV+TvxzDwcjktWE7
Hum7Z02Q0i4Wmo3dMwppIpiMqLRDCRgYTlIw4AdcEnNbAWx1/tI/aqnYwNoQ
TMsxoic9xIY5AQp2ZHSOHMrwIJjFMAqmk4IGvNCMheQ1MYD2azbqPhHc5Npm
cAokyAZAGtSndfADUYEhxcGtIgZZh0ilNqRMYNRtffUYsAatfC0+/YrafdIq
gmn0/DOuW86abW0u1y/J7cllHmyionqBUy1FkXj1uD4quR6nVFQuAZWe+Oba
/FqtDLZGl7E4ald4feGOLUcpCjThxRbuTAugkFYnSM2TvgxRKbeQ9t3j6rPq
UGQ6ENw54rljzQHE8s8HcRIdfoMzd/oD9qAWDb7KkNeFfZDkgCSVKdoYHZWn
H7R1gcEL6EXlyniPiKVfsCTvdGY4q5N8fgJ+tOr16RDTsJY4ZIUx8rOErZzJ
fMd9fAj7XyxxIVQxc9m7ZYNtTH1OYQKiGgyn0Nirhgt6AcztgL+/NVOCJ783
ZsCxDl/0QT3ij8b/evVeq0/R85x2d1Y39Y7HpVX6Sd+lA7w6nCsBMZUeuwWQ
/qWaMMFAVCiBfy+HWLjAgu2NzUTf+guX845qzh0DvWZu/06Ig3uaQUzvpC82
2pL9m8eGW82o4euP8F1FWlpiKUzinHDwtvX2GclkjEozqEf1sfVDWnFQ8Lbk
hxoqfUNIIK8QDvQggVKOl8/BLNIh4mz/r28BzG8rvmQ40u5kU0IOy/3OdBLX
0o+7mu5NWpaaq5sj8juS44bK7JE8rkVX5p5BmXz7y8FWiv/95DbmQBAMYzFX
r/3ukBcx0ir3u6GhOEDvhE/nzsS9Uu5NKBGGSQL2o8xNnBotfGQinw/pZ+pJ
zxhAv+fzHythuNwWbsoj4hMBdo6TENrg+JheBscBvF2YolNRGfhQn7KeXzza
v87P46lOW9n14uruF+g1e2+lEx3ShljmxyjcqkTY2JmCREnJvcZ6SPd+3+hq
qni5WCuB/SEMzkeCBVdejWQ3vEiO+IGEoamEG2q14cbSg4sfED49N/5F+BsT
AqrW8/0jVYM3UmTXiZ59oN2ageYnUSgRdeSx4q3eDBQIjsbXQRbhH8Ne+zbA
A2o5O2SQYkiBs4ngKr56B95/QveeXOeN6IJ1rTrcsRgVeg64EXqkME9qFfHJ
fTq7mZoS0vDdrVrZ0rWq59daI/m2jq9ufZIOqEixmYPDYindAcTyEfTf/702
tm74Od00kAig96Y3hzx022/t7/nrytp4FXtOW3v237rZtf67qMZgAwQdTIEu
VugSl79cEthiCuowSqUe33WMY7mhH6+oYQ1WiCRHsf8b5rek0Nvu1sNppimQ
kg2zteWZ1qFiPo8FE+Ouwb7zBtg2Y7Aj76UkyAByZL1zt+IG68+Pa/bFlhdG
yu4CW2Uelh/9YdQaPT2rdQ7IGe6jaqtzSMrj8xqwWGOeQoxV5DctxYQRs7rZ
LXYT6ee0oJm5SkzbgldXy4rBC/nSq2OjMar2CxVcEUMEteGkxrxg2zNIVnyf
ZzwJjQn+dCnqi7asoveKKE0MApei5nmYIzhWKIqc2rLp2kHIojEzIIYP+7Xx
4jSkVJtopcbXvSODoKJjaqLgvzz97d0tYkU96YrQiRRzd13UdOknBLzCsOjV
SevCmb7dsDq8NoYiDFVtaRsYz2Ov9l48zHxbIKswy9Se+5PnwFDanANigLFq
CnuviS6/KmRCH8v+rLJzWCxkJQ0N7sNu+5Z0GN3MYuB52Gzn55JB5iut+Q4n
gauoJBCwQVRbAq68fxTbvxb1C5txAKt2438FDnEtve5v3HJgWCnqFxzUVAdL
fl+7VBn86zXm3/py0HIYTVivy3wt6y+OiO6rexS1jYaW3LddQ4dbnW6tVFSR
Mm9v7lQ/tOzZEtCK4AFLwL8Ax19UfjspMjeLApnnSxMOTI5L/LFwLIvDU1Xh
VSzZ1Q7H7Kx/IZaTbtjLsFopG6FMfYAa/vo2ch6inHJKeNsut9cdSO4zYRpm
u+xiAUgf/rW6xluYh6Sxzm35cvlPFObRT8B+vLiWmWmI0AgslLyxwXqCnFwp
Rv0A0hpBDGxzMYahxFxDnBWIJVrfhZJfCf/jqwx9/5cdl8Y17LAHmLFflSGm
JAgHjutEFWbQnhRJ7HmhXV7j5w0y14m+hcwgkZwFwXx5WRRjv4Qn1lWMtoGU
eEIZ0i2kPbisWORbei0myNgiTFTIa85WJRG1y7mF4A0GNBnvBxTmTU0FEdwn
pMWmxu/77v5zPsmHZpNf9okT0kCy+xC2SI0M/BEqebkhVFRS9swlKpPlKETR
qfDHeriE+HrbUyumjdqry0k+1yrjrNr1iQV9TjUpjjKqCgJ5fccs2PewO+zL
lsKsg/ERCexOMHstBHspZHhuBKZUBUqb7d0FS1EXAkEjzqDi4d+axsGf6B6d
haLNpE+qo6YVnVig53R6VLHV0vNCVKd3x+txsP5awqssz1UfC8NZSJ1KNgGt
penUdV6nq/er578VdF1HsGASAYRBCOb+zfnVtV/nfySPfKhTxA+AEijyzC6S
d5aszJtPXymoGLug8PiG+BjIz4sY/pC+Nqq4LOo87XSoaZ8R6E6pL82e0DJE
vPzFVv+sEeIAbO7Dihuf1XHH8dPR/J4//HKsjQ1LoD7/THg6zw+dY20ic9fk
ItaJxgHOZeVuHg/y019/lkK6elhILWqt+VZ16irn2IwS+yoxQCEr3eyv5cfR
2SYIpwViTJxZTcOOc/kgU2g8vM7DjBZ87rgsN0bCoQE3LS6gq9ogc/MSPEUT
a9U3I56TVmpY4PCnZM0W0kHkEecCzskBFwL2hXFMfd27q0QxChxcSCEsPjt2
TX3ea1ZKhcM/zfJHPhrfzmkjI2nYrxSDR0CbvSQ/vCMLz5rgJodj00SmxKJP
XxK7R9EJV+DUU3IZNreQ79MVxZ4yS7XwhAgYBfg3AYIeWvbHMwOawP4ZLNsH
j9jXiLTpuio19ZnmhWsoonFntsigg0ntqjxU4619zZExJ7LFW6L/Q/7A4bI/
zp+Jh7e0QzV3846RJxCjIXf14VJ6Eh6MVHxpWDGOmcK8Iy0lPzySFC7X+blg
+TG+qc2bX+kPJnBrh+V1ADXSky8TCN06bGxzHn3fdjeI2W1BvOUy5vpOQXC1
za5BpRIj3tbbK7jQWFHqS90gKBitrGCTUcUom6VEpqEqacTjred90WBZYyyx
rZIkkJt73dInYEQvQ7rNPPBeCkohuRO4SYi1rzfe5v2E8sHs9HG+u5CYyVSk
9rRYTo4ZkTdbo5lwvL4xiONZb8VA7MrzYq+lTTDd2/wtMI5ok4JysmR+JGvo
5prxmg4kt3uwJaEcyN1JxB0I7J18axoco48kfR3Uv6aqkhQv5axmzYn7Vxse
XCfVEMcIoX3VZnKf9D8YO8TTUnXjRLYnv4CL6OAnV1UcFhFGfL4hqfSxppI5
9dsBE9HFdcpoCrewn+/V6MXKgpvKMkUGoXV6Yol3LrKmvuh1h68tVLrR0eGM
nWboawFqOiZnK1P8EDqCkWPLzahA9mgx+jbMT/qeVS3m+x2oMD/5PXKmmFmO
8nDkNS06WDhDW4QUVWeIoeUy78DSozFHTKI831FekYhmfuhn5XolzLvYq2jE
dcQ/FvS1DI6h1LGC6M29TFxwvNQNBWhOykAX0DeefR65iLq2q0B5yAp4uE0s
W3Sqxh5WaWcMezXxK4fb6B4ZG9PNuneKCwOsvLhzV5uHheIa6ZRxET9zYiUT
XPIJhvRUdCTdD2uCJcUSSu4XoJ5VPyjkZl6hcEq5VV5m9SnkdbMWERdk5J2y
YswP78vaKPnCfuph8Juom9M+8RRn8R7tK5fDrWsrfkKI1fVu9vFjcNXmiKu3
azAy857oyrl6v8iauWxU7lfJ3zYuysJl4Gk9hOYS/fqrk9zE3zOjeLYuxBer
9pJAjgmDsSnB0MgOBH2p/UwKGT/sDldOEPZ8vSsX15zRnBFVXfwqO2d0zhFH
JZOY5AK3b6rxbXin3Vx3TrA9CVzkfnu/9bf3WZWUf+VSpkTXzsB/M5tfzNZ6
iC0N0JfhxSDdJvHVwmxwRA8HpIjQn5ddTJhgdtNxPO+75IpCL2PX1gRv/+oM
klfsocXZZ/KcmwF8Wt/ShBKzcM8lxZj1eltMli8JjdK8htjOi30BRq7cKC0c
ugqGjuA4vCtc/QYhzSu2O0zCGpifkQ3JXua3JgsQrkFQeHpAhqFVtl3vItTF
cEl+/6hM9eCXe5GHgLcKVUFZA/9UcirrWfFsqi+tjtAFDlUN8zr6A9RRmdEt
1sxG/TEC7GH30Qv7CL+7eheSVfk9fr2ZQQHDeCLFLC5cyLET2dstJ8oCkchm
SnSTjD66cJhXG+a5NpizBuqE/770AQD1s/khIIGnxgF9T/EEG2MPR3ly1x9P
jBZplmcm20hMh1h6FcectQTsg3FWcVUcr/tV0InzjrFY85MXnD1QsAFrsCaM
x20JQF+ttA0XupeFJ5e8rdjyeAEPWOgucYIeyHKEP0Na+KHqbnwGV7ReJpUy
9FwSS46l5XAvu0mJ1/S7tMd/tbs0XTSrUJGwPp0iyE2jxxJ1mQPlApCgBB5U
GHaQqUJKak+mPBT26WmxuZWAPkT2pNmpOGLLq16h6K95+azKW/AFHihe/VnC
laJ5SXJn0uH8XQq3uasYgvEZrb+EeN1fUhNIPS4/zq2Cw5MRl0NvTIbuMNaS
gQVDjH31n4YXtyhPwePeH7Yi4YAxFTuoYQzApjOGGXAtvsNsCs/Lt7E31wfg
U33NMgsGCnMo+fv0bkqhI+rNejmBwVejn6DkiPcjnvBVflI0HfOfd1xkUqtS
Xhb833FI8utv4hMzNNj8ylBLLdaCm6Lkw/uNGnj4rfki86TWsvKqN57C5csR
OHbRIqN+6WFDao6KMMZTqHZHR5rKCjBgfgWzUsCQ7xXPVX4HnJ48i1C0TfCz
wPFN8UVjQfby4B9tGf0GjF9MG1qObpUFCzColSxmY9gZUllutKGqHREsgHcG
PF/p28x73PR9TXnhwdo7+iqmvJziQOycThd5gboXvcmis3kTZe6Rd+ROAydO
CC98in/lx5LGAl04DGhMsET21sHHWipIMp3lexFuv4p663C3CjEMGWD307X8
9K/VdcWo5LnS4KipnT3rxH06qDqLk96ewSZY7Z26WLylaWPYoeoWRLYAUic7
jSuWrDkjhGBu935Tejt6qtoG/8Tndq0ysE0EGd2nxSo23ZuWnRRU9XSkmysL
Ay/nSC7sOP27cqM2vECOpm0EH1joqKu+GmXwspiy/x4Cgp17hdkeh0ZNZd+4
NkDH1liilJ3CJahVMvzh1vBR9nWrGJoFQSYPoe743A7ZtjEffN2ixjUe5nM/
wkS/3i8wI815IE/AOLNTPwNROzDhiIrJ2qOiyo7ezIHbQ0uLKmAIaXMlswPO
wr+qp6lYIfbiUtm75oPeA5But7px3drMrAVQ6G8XI1AFI9pglcNWBng3c3UY
kTtnuGgGd0fNU/FWaiEEa5pSLp2ArVeiFF/ZSd2b7+Js41t8Ye6p+rmC9nxR
AM20Z8K9nP149tTSeuYS4Rofi7e4r2CNfYT7//GpAEHEkOqfBKZ3y5PMknGx
BTKYGpf5Qd67GL3AZVaLfDx0CajN+xvJg9OIBLbQ44eMBRjXCOeG3OsE0YuI
NddnOKYY1eviFALYvk2vQv/Uq70JDFdbsLN8bwH0hW1uGzAH1nENRCaRHy4L
X+WDd2Ue1Aam0NzaRVUevNh3OMkLuLEOW9zjkCXP+uL0QC/rgBP1gd6uXXZt
4aqPMJSRwob/nUTUzNP2J4oURUTZwLt5KyvaG9ZMm66/JT+LEEDdlv6VNySD
0OhxrG1alx0qgnwU6EnO86cgme4qUnugiLgoM3KbXenGP8U9tn3kyOFGU76T
V1HlR3erp25lNTLXBhIIcY8LLAR7xJrti5/JmLcMRvtnNpqCCu/y2mgaTNkx
fRNlfBzY1RDF9tAs8qH88SR4YfsVq3chkvwp93dJpL1tGrG32oNnK+VOLD27
z7iUjV5G2Lq8bDm7d5tRzPh3Xy9nVbMJCjhxo5GC2xCNPzhb6cI6M7uTWAN3
k1JrW+2LmOTcDfReemIQd3+cwOI2e0/rJREtLehUfSGWZjuZTs3YCPxGTROH
os6yHedATRPbMBHpRUecWWRl24o1JOCuY0PJ6kLQLLgagvKQGnqh3IIGtUM9
D6ILXT0TjWtJ8o37zdRhV5YnmYF0h9b9QSBrbjpILIg07U/hklkgyVHMRlky
GW8vIizj+3mJoXTuWOQBTfu/8pHgBjc19++Rxn9s76XHT/fG3vsK9lziZEwr
QphIspIxzE00bLIW9uYzOpJep/hm2waTDo5019iV9wbzAsbuyV/BC5JEGX7r
sm3PyT7VP2Rz3C5MBqD2kqmF0wli9alXt1diXI+dvdjcNnpLRvvgkWef+x6z
QNjY9JStfiZJPOICiS7WWP1dj4og5RrDTWlVA1gcwwynp2YQKtYdJL2NV0fL
iO/EqWvptuv/idTVyxKarW1v7+kQPfvZg3po6qU1V8G9bXDEtOp8a5DX0hUN
m1Vx/yiQcVcGArInqyd5F4y6xejKAqexVCVVGjw8vaL+iFhqYGR0hyuVd3ST
MPqUkFvgW56wbZVtJtco9wuP4tEpaUmYvKymGCkILawGwOgFigQnQZTkInFy
4aDB7CBqycscANBjaBt3nN2jhZ4cDkCnFXKmX1y49ocRMyyKk/TPFregLrIm
bFTAMtDBgQ7Y4/Ixgs56Uawh6/wpSA2LIdpfNgh3cK9oMWGlv/pZJCl+F8Dm
hgHHo9R6ubDQjDky1/POvTs96lf2TcYC1YFoq4/bIJ7pKsxw1M9ZsSVq7+I+
N/jY8ZLO52GpJNzPH2fXYEnhWA9Pn8ol053Fm/lnWqIUBxnLot0LJyZeRSNZ
/raHhtt8HsROZTtAfHho6t76ZyrXTd+6YgH/BgtYJJ4IvLBN1jfz3wrzqk9/
LHluiIk+yqva9iKNZIm0PvJyEW8XXw37K045AYXUG5Dn1Vj3JAL+w83xIxlq
+bON8MAUP+U+0YErbGZFq19yuPvsETL0PVH+dAicQkELzCpj873qg3PXthim
eCL5JZ/9N1ze6C6RTH0GEzGgiiy1ZC1DGJtEcoDvQ5fURZqfnc4S9RShI8gu
/oDCsfk0OakCcZmzvLuB+6SBARERon+MciHPr6t1LrVIHTbmsQBK1rkIVnEL
6gUyBXfr3JekLD8TqNTsonkiKsT25zMJJDmWrW72WZWqqeNeMwBOeh1UsIGk
NdBYLZYxXG48RgKSIff50L+ulxoF9aodUIpvA55sx2S+G6M4ujU+HnzNmAOG
MzP6Emntpvzagu18/16zrq010pFtVbpo/xg/GutDhSxQzPwX6XY++kYC9wOg
8CfsxCtNigfqUddvEDSsQkqi8AO4awSSh0I2pzHh81Ak84bvp/IZ8ODj6weC
aQ4FpjcV7tJS+gUIGrB3yBDMAJkxsVFoHTpko+ii9/t0bpvFlnl2YkRwSKNK
HejbO2hl7O4SlQvHeRnpOZsdv2laYXSRy/vx2RjzxfmOQ3KYwmevJmdwYw+j
SvAuaNXYDYRdkt38Wn7b/MBpzE6vXFODJdjBXwQrNZ9NDUkClwhez+K630/q
YQ9I2iOVKg+DMcQO1NrcAr6BmT9JKYOskxdprBmuEnPeQQjumM42U3xKsajQ
0nzh2rVjKtEhlu/8L/MKsSDah4+y/2EdSIWIxO57HiSpsD3VhNEXNlAgoTnO
Bdo8Nkmef78ATjMeaWM3DfdwKuShAUaXhrprqpBaQKU2GGN4L7pRsgLdoAhB
/Wbaa9pCiQeMmN5cd5YG6Yw3muKjKq38OPt5WS3MIo1tUq9xXdPY8AZTDlBn
9g+y/sHDnx181iOjT3aLYzaXJo+Tptt7oMvNSahiPSvaod5S+52N/rM0cK6M
/hZxoINAhbVr3YskiFEZkh5bFPcaTRhDt+s4b9p5lqqoElNrJ2zlXAw+bNQx
EIUWTrVD6EY7kU4+dmIAfvxQozsFjTFZT5rniVKwSv3vspz+gYPJPOc3lA6i
cFLYQrYd8lncqetRkU8DvnzOz9EjXGiig45UTuoC12aRxL3av5MCqqmA2fU8
mWn16OojjCCb2TJb/ylAa00BaL7hhGwLdfsVjen+UhTn6FoD/oBh5VNIZRxO
A/U8G2uNGd1EoTrTwrvYgGlcA9QRj1gMTXIrp9w0rkkhq9707zZTQGSEVk9C
Zts5Ioy2GuUEhuj4RAGN7Mwra6j1bGsCrURpstEnBIJwX7VoemK9ypCy00jY
PU0cy7XgQrVbvlTPmD1Lmzey6/kzyf0XUy06MxqvCHEKZMwssRWrPdMuPSF9
V9En5DI0uE2bBoWGUmWNaK/JUxHT88b1M16E8H+8uTGOrVB5Czg9ghW4hyh+
it1mtbUosNYWDZLc6+ZvUsOZZdvuKdrcJ9fE47N4FzLsrqPHGYit7/xElewm
GCT13GpBgMCjFgymd62ZBTHYAW2LtXYrCrsAbPvWx9R/tNMFEgYUi1Q3n13p
NEzVhEGmgQNjBy9+TSVUr7KB6Snhbaa9dOvCwyuPbjgw8rz4SN+cpbuMHTP9
0GrbCnmlPn1dJh+mrCD+B41L2BjGDeWYREspjjaTvTDUfc43FBZJ8wMrKuUQ
ih+fKObFwI8vGsl9Z8yaTwIwFtw2OT82b5lhnbEzaMWu0oua98iFCmyJ/OtB
IvYW5tW4xBAemN0YlYORaj7Wak9MvKSTmIYmwd3IngkukDoUePihtnV+Xy86
OFpEkQp8oiP1NntIZnqjLHeviMNQlTggam27pzgVlEyQMJhipAdIwnNpHde3
kQzsVDDCMt16vUrSiMJzn2gn6XuGkAiWPUlAFMkBTsaoQkiwJT4k4KJ8pJHw
MTYfh3b0+MfZsP0PC4J4OsI15+WqL70bnSIETJVHc01h/vuE0pA+Zry8lQIU
ty5OG2bQTovVefvZVyjqUjUBILCU9Xn3Cf4tvALH06Wb3a+EB1YV4FDOMdpE
oJQwj/LLGtgD6p5xgYesUy2YAdBJs0EaQ5Y/DhBC0AEoMPoOC8ycUDc3cp43
Y9/pVcAy6ySBZtQ1rwzju7/1GftCm8bcjNHXVCZQeTzhVwryL9J5X/WxoNH7
AedEciD5Y1Lp6F94pufITfr3G2TBkXSdU49BbV4pQjUto72VgFhuArJGVyDU
j6H22k/GCihTDZV8CKwYyW3Rpgr2kmMLPRnRZ3wM8b0FEVpA2uazVJHcEO7o
rQgOYmbwo+o3KafQoOCHcEkJ3i8nmEDH7oxt4WrbIGkfCpTN2bIDs7n5Sy4r
K0GGE0UjNFqv6YMLsrs1lMzxbCTOIFQWiIZAwx/hggZG3jvLYnZH5hJMKuQC
0UTtNAozQZVpFXbqFcyqo1hHV7eMMfluoQlotIZ+8V0Ut+wMLGcLiDDOO1WF
IPpLa79jcN1Mn/pbIm1tyAAW8lkFeHUccSefzbgilGrvMdhlkOtDicNIkotg
VZaUu9RId7UVJIAOgNWqUnCWkOVATngwJHUv3eNGs6PaTVGECUg7BJiea1ab
rGB4DZWnseqnPfIv0eIvqItZIjrF6svMklYIwV2zgpQYc49Ig7I3Cvbz9vvz
LgBBiqxR/K+NctH0KVLKmJb/LyTLTkqO+6/yQL0FcoDG89auBAOModKkpMsg
c3c6e+fbsiiR0gvl1oUutoW2LOzlp24OVn5VxZKmzA1hPT4+fqajmXQoQW0N
mIg+PIjBY7wTXAnp+N1VwmCRDAUvT0Y0BbrI8mRxGwEMSpJZFF0BxfWElu10
KsDDmj8tCGvw1E5nVvHjdrY//KJm/L2/WgnraZLpsLGkxfKzzN9/Cnn+R9oF
Hc5KhEWAOL9eUR83KRNXQlleW29/AyLTQfwoOYbWvLcPnb1DpeAXRQXoriII
1JRyAxwJo56Qgv1yAg7VZ0N6C+mcTP2IMWUkGkXwipWtg4hONxdR0PoDBMQ0
s2ZKqV3zUaGHfbFol7ztIvQ1FUr6sJd6FI8KjSTevRAx+i9Uef/5ofvqY07G
w3OAUyDKxdBImtNDdtqDtt+tuRVX/kBCvcvCk5e+QF87vVO6YooPk7+SWfxY
M/LgZbnJWaFVgD4pIcVPJ3bO9VjNVes9Jbfa+XRnVKhrSTbexiRCmAYSamm4
sa1SJ6YpyNN/RpUHMvBOyhY6eRhBdpikww4T30j4RrTUwX9AgF9QFQtKOgTO
rb6xdcGv4v0xuBNlYOY0ZT0e/F7HQfZqjMlswzRXhAOFbbcyXQ4tquA5q7Rg
ZbH6yamrm90tCFF8q82bs8NuL/773XuWbI7QhLqlQbXI+w597dx8wngNDyy6
ZQ3pr1qppo2W+2miFqJcwrnutEUZxfeDCM+JAOstCsJYRtj1GTdrTbhniTFu
e8TsQvzFJalRABbpQBA0tl/kEv6E31RG7Bh7U61Rb27y3RtF5mj8iJKAa9yU
DP8BBzfgufhSRJ6RS3exXcYZLCMctdqMy9GXdLA0FDiDe+VH6UnhpY5bMxBg
Pq4RlmGLIZsaHpLKI29BlP6rpZ/pWxo7iXni5yX3lXw4xVn+0Vz7j3iITrWX
lfWASYYVydOlqHif55wz8mgYZELloEkdnvLKMsZD86drZrpT6kyMdJTp5UB0
1OYn6EHNUyxR4R+c9brO1hVfKpOkMK0rGzjDoXQ9sQq5GhDhzxYHpn11UqEW
II4rRrzyhVcGTuJsqdLKN2+RjKVpjUNfm5Wj2oJvewAcrmMLOgo1mncZ+QKc
NKIBMs0T9l8qW49/tIVDuGWSrhLUAr18Q7SE5eXOkG5AUrKc5dl3w1o9MLv+
Y7gDF+cBfNDtl8YPk1s7XyXXSJc+nsyMeRJukWQol1wMEKV0zrYtXoxkQZ+A
65iz4zEwDV/RNBJRp2MI6wgLeuD3yyO0DEsojiHJo8DrvK1ixp7t93elJkPG
2akIUBRyfKr1+w2HOIqBld9d/lZEUzYYJE9rwZyo1XmiNFO4s+9bp3zcaOHY
RrSaJOW2xEp9teQIa7OHLYQ7H3FdQoeynORjhJkyQOEmrkonRSQEOGbrGFeS
HTVjn8nh1fOLw29zGIjNFujGZgge+SHN+CE0IoNaKnc1RfZPk1cmB/9zj2rK
N0QgOlucDqeDnkLYLAP5xTrF79uomrPhcIBkAmJV4zCtWjRauafiGpj4xqmb
wLLTMCSz9V0hro/aBUBrgz92UT3vp25hRrlKilqQkR4gUIlhOmmQnbtXa0ka
T5yQ3gTh6UDFJVMcFe8kFHQzdSc6yTAfCqyrx6AuYSiBcJm+LinCJ8DrZyDw
Tz6WmuY4eANXD3rbEDPiGXFTRIdhpSL9i7O1vXdviI5KgycJyUFyasqF8iPL
Eo+CdLG4MQtiPhBRdFGiGn2KaVd1yehhpybwVErmMNniE+ULrpaEob1YZNPl
1XZgbKntBvw7B4uAXcRcNuSxRdDVrmvBGECGs6v+0LEgffJZ670LF2SFfk2q
9ErF6wiOJ+vhtYiCOhdV7TUitqDGlQ8vwZ7K0Eb82bUYhj7ruz+aRLWcvgvj
OqDAPGs8nSbJBgf54NzRaKeoTyDi5StVNT4KpHL8XGWYpc6dGt7+jM1okL5x
ZoQClv32XdHgqzRrpIQ3q9puMDahUd1tchXm6JKitzzyoJGcVBoNhUjDs/N4
DLYgzGln8JOHD9mx6QD0R9NblsagXUXmkR4AS85KPf0RSA7q2ODM+cUg7I95
9k4an1/cXHqzd0wgZYHcXBruBRC40YYsgjjr5UMrvR/0v5pJAN5o/mjTalNQ
YvjyvpF1KTwUATf+v8mOdsUaxVbqMxzsFnoZbdDeBuLUoJQn7sQHqjwIy1WH
lLuMHedl3SCBft5dksjG1O8fsa7kIAvOTyvMy+8fXFQZVbi1DWbQ5RF3x+zo
SJVetoj44m4xDBhNNszymn9IstNB06AFE9DH9gnGGEcGblfs7QXUAzP2f2C7
se5AdpDJHQONWswXTS/ateeW1jBGD342Xp/KU4gvfUSdNWHQwmNKi2EG0Vl3
wAqxyJB6BfnsAW2I56eeZ805kMaNrWvS0ojLFN+cvuhjZaDH1Rg3Syom1cU2
KvnOXGf4UtQwXHgzNoi90Z3Vyxu3jlalGSvRn4ldUdI2R+mc414iolfqiKFy
lTaHFiokGSCDc+N7exBsDSGiMIM88NsTQDoquEPFY2oV27f8a6z3lLIAkhL1
Cdm/gW+3G1uJomeRHTHgKYwB9wTvGwdmsGQJhQxKXr/mdgXwCddzyL4h+9+R
VEcuEU2frsdeglCqDeh4UiEPpniXcVL6k9aXRGv/d+yBdOlc4sa6SlE+/cUX
Z7yyK2lNQj4ftQkMpUgThVVogocxXvMREyg4xryeGzq4uYqtfzkf53Vz2EME
z6wKnYmnBQ7RXRixsf12B1qF3OYRBgM99LYngHilA62jgHSuDoUnnCyU3afz
m8VCMo1Rm4WFhUCwaWPud2Jecl7+I4cvJnkMpUKpMLYFdo5NBV/+8Q6EKdCS
mDX81HnQZqvUgtb+zbL1d38M8JwptJYfWceXJJTrlLXz7SNPX156y2gIPo/u
CaRMESx/a1qIE/CbqNt148IPt0U/YjGYyom1G85q0p63lKPQBlQYiRGgVuO/
MuF4Ld/NnKf+6pUrZMNr20w5IvqmQz9NwRoF097xEDGduUy3baAs5vQYwMNW
aRE40naZNdEIbDFWBhgZlSDOWFDx8htYCoqZOr7cIzg8cjlaLMj97qbudVqm
Zd9WIEdGZmKSq4sbCv1pxDBfzy1Gvaaqj4MHlPQlimyd3UkKJ38AmVgH0DLB
vV9NO+uATp61MfuERYqubix/rNexAgpem4nbSqTix1ebKJIdmSl2vbjb6erH
OmPNo21zzijjasOeKSV5+fP9dIkwwKZkM7Ku0e6kvI24X81NQAig5FacPlpB
xg6mIs4ivMc9jd7jQZRP2TNsQIEqgifsdqb1L2UcgLIJWPQg/9UlxIhJeMZR
u4qscmIuV1cvpl9Jt/E+sf0JvNHXCZjkRRs3RIjKeU3bkCg4P6RjVzFC0mUv
hHAqWPcD8t21nSbVh2OcWZL92g3vMLqtdrUTyGMLFTc8tkQPkOJbzjyY4ACS
fbRZh5TP87LhxWpcvJBQ2SlpWKigB8AlL9MwWlsYwtt/eaX/zg/NxHR5txJL
N/5uTMTRHGJN396GgjO5l6qO06pNRqNzDThFHsWUFtiko76ULQQMHfQ1V5og
2CVAnxcqMX68vuWCqEYe9ouyP1OZkjYF954qJ5fNXCWkhXR76amDPIP3re+U
O8vC9f9TYn1eQCQlQ2RepKtIHFmm0MgW8g1EBQCxH7ee1bQ0oP4q4slKLsm4
Cyk6OlEV0HU59C8Qb+sKF3vnPBmcUKzA58GMXWLyH/ffB3DpbNipdSnjIb5m
sAF0+NMvrJMpjTRJkq8bwgaJrirMyiLBuQUDtw7H+P7keQHM6e0h1xqdmSPL
TuT9Vbgmhv+hBR/42mb+0MxqnCotME+vzam7KYKW0kPbl8nexpTHuC+sbwmS
tDzw+LkkXJ4X0mawTMAayiV6TH3c2jfybZJCh6yp7yALHalHS8KpJV6uAPna
Ypn5sCyRd9a0gZ6H6jchU2N60uPhw5B+3gYXlwoo/2mq+0dME9SXPmAmXW/a
Xxl9OOczrC5toZpZr0pk78mcy2wLgjl8hJQ5vOX6zYa4jWLyWbR7saDaakNr
sXp1pLryvqj0UA5z6ZqzgYaAkZ9JUswky9/VV28IhfJ4mML3ZtuNleLHiYhe
EE9G7b9xA+o+y4dH6D8/sOpp59lK2mmhXlY0GyFPCKEG7A/UAjdT5w9lVL/B
HmsjQ4YldQaN7l+ZbIRqxJ5n1uyTbf9WtSW0GpiK3nSaczUr2FdtYWFKaLQI
klsyEH+RvK45NmepXipny8XoaDf547gO+P3pjJaXQuQYG2tzfHXrmd4fJ9P4
/WccK1ONiO1VsH82IB/lmCiUz9l3DhITYyIqIzc86DUKEeDaEJLs8P8LCiaK
LEWvozINprVUIPREaxIeX7VYSKf3RU2uQ5znKfov831QClNo5IqZP+as09cm
pnzGqwLcUvYCTVYwrvCqxem1mR1I/CsBQsrXD8C6S3CE3NzKxDCJQCVt7zqG
h92GY3tEPz+S42rgN9jg03UxmOY7ScBda0ITpZE2pQWsmMtHu0VIWpD5cnlp
arNhwhUBflVBRkbcSSUIwb3KSlH69klR76jmH7qgBWKOFd7rPNHPgZwoqyt0
UfMawTiVyzlHsOzHVDdtDLNtVcSw1olRjWa3RrZF36dm/vklGTYxcnt92Luj
d5ClWNnW4C7lkcFxQcsIkkeFUvJjqeHopZ+pNy+FTLoO8crGl1ip3ddTfbLQ
ct68gTic40CndN5Db9VVGQdS/hW3dq08768L8HHw89L8hoU1QLbapaG+RxCG
icZVy8XlE7CDvSncnrhOU8mO7OnDrkRYlN3eTHJFxzv4b/RJqtAyk85B9H5v
OtzgktR/7Wwfwa621UPUmPPsdsKUISWRAk+gTnN6CjdBucQx0Bg+T0FTMK6R
uBdslJ28P95dC9xIPPKs3pCpu4u/hrtttgh9uwpr4qUkWWMblr8Y1woVp065
ogGQPlAHmQnK4krn01KWs7pR96ixKj1zbzK0OBhc0JLodfavdEcWwmFREZNc
QFLdgMCJEyS0No17+Saelk/GFgJQciqQlno/KYJCqjBJa2izkMeg+9jmHeWA
cfmz/tQP7eOb3Ag8mQh+unsaRE8E3FxUZR3PpoMWQHujRcavZoyRc9SnWRGA
DTamb0cylx15P9Cgen9cCljTHXF3mFVLtSHr9NQN4c9JSsmGxAPxP7+yATB5
NXyb4SPwIO0dW8mCNPEK6k539cBovNprAVRMNuDH6KJ22L7vtX9RYEC4BUaY
p1FDEFkwsn0G0z0NrmMcSm7D2mbJyJdlVmm6eayf9e9oPzYsftCKyxhYu2Zc
zxYt4P94CtOd6jRcF2T6DoEEk6Vy2YXCgPPNo1l5G+JPVPv6xtvJdfK7Wemy
Ueea9HFwGSps9hJIIz8+kosy/NWEpRlqPMdJKD2cW+R+fuM+c3KYwKXyXW1X
SzlrgSa302Psf498p972Y9NxR4EkDVRG7jp9+BKBLwTPJar9UVDOnrkoEC6/
FXCxXdr77rsSZxXDn8/vl5Sm4yOr1q5ikSwfi+TtFqHtb+U9nwAms9kFWdMs
xySvfNzFdi0FVvGytind9VoSW63g5NP28dSPydFSX4/H+haAOkdsGgxh9Kw5
wj0Zbhzgy6r/UX7gGYVMIsaUiXZqMF0iwe1qk/ZLuy5l6RggV0OCbGrvjqpf
mXs3DXkpVAEDwEsM+MVjn913UAzRUT6FWg857JXGlL5erD2+Iz3+LWYUn7UY
+J/9eK50DbUC+u/gC8Yd2U0ev8qbtltnsPLO1SBCoYFjOGktl+xrMAuLshA9
QgXZvYQi8DmMFr0InEpISRsm6vqz8xWMEJZmc/Wba/tXRwt9r3yqt2b/9FFE
zfVmmyocMofYbs49iXXibVNX0DDRfQ2BBP1Cc+ggFdy0XgcpB1fVnc7gdNAe
Orw5ljF4yPFMUXlYSLgUQF4zDzhEINYMJie45SoLn0FOz3vibWfKj5bzNSPK
DLL6hCMUsYs46oPuDbG/zfpOs0fsaxn+te/u9Cf2Kts8Kbd45rkbeTwCFdXD
tJ60AUecO4E2+Duo+6dBqfW0FgFvuTBp1nnHM0OiqrYg/yQFzau1R5XYAiG/
cQrqd1Ca+rbxYArOYEeCmE342HGDi3XQavB2NoRo64Fp3gSvOywKlJjedNxl
wfsdJPE4LWmei/05xnhrsIK9A/Hlg+VdDZfUz/loML0y0Ps+mh55n96/tWqY
7iqOOazjYjDUhTheM8mkEMpfs9MztEx0o7C9uDNNy00z0wff4Q6fhhoL6AxD
j2pEVgO8liJ+Vl8mel762PYTnrqBg80xuXBm2M2tmua3lOjMP2gFD3wP1SBA
5slbBkucHyUNyoVVLR0zgUdUbqFevsTQPPLKcWWdEh8HKhQ94SPnXDzQ8cLy
AGda73dzPeuek5Uo6Ud9Cp1Vb5sh6rhn8ZB0wlTuYMZcoR26OoYHbDvBUPpK
TIDbfzuIGYuVQ1tNtXVF/LYjIZ17KKXaanjM3HqO6k5BAsltDTpoK0wKVHYi
ixnpSmKR4WsF0WRscfy1N/IfPTy851qgrNyqkT1zqvZZF3oZNMq//j0WKovL
ssGkdFPWC23vRc83MhHPakpIeBTv02OOri7XVD5ZNdBfDPM9M797XEsjS5U0
iVkEbpobq+4MSHkJITfFgxWB9WR2QgvmCDLd55N/+Aosl/HA9r0TRTSbNy3t
4dtwvGxxscSE7wd6y2EPKRplc/Aa8j7XobO/fcEc6dMB+EzyWSE7nqVeIEZT
9FT+vA5Bfh5BRlgeO8pBIH4hPEBN2RF/8Xvq8klloaw/ffDYuqu9DRmav3vk
3KnLc8dwmI+fflk290EmEQNbdMHz3+VfLac1D5lWqChZhp31k3mOwFcDKCIM
V4rSjEZTHTKQwDzzFjL970S3xQhWL/hmrJHx0Y7mebwYsa4mWaCVZvud3Ou5
MXPcOVPKWuo6z9SoTcsA/Qh2M9fDxc0C6OLzAdIKs4u1B6/BPnpVsdMDFicD
BdOXggYYp1v1lg2OjApGkSfEgj3kERJYN1lGv2woD0moMNJJ8Pot4UvQ6pk9
u6XaVW6HQHvM6LnIfdmhOUwA4kFAgVJ/uFnCbycFwoRc3aR0t/UMZVhHMTlh
QRlcmx5ahWIYSWnUMrAk41FeZH80ASloZedFt7x+hD091uKoSVwPzbh5uxjv
AJu88BuQdKJBj2uqNE8+nHZ8mGizjKzaEzjLajDCYwZ6dDa0FjhHgzlum/kJ
+Tkq+LRf/raLscZEfrqhq+Ak7skel47zCFTO2/xf2ChIPDWI/EBmkLs4Qz5d
ObmusisC01BPUwtRGr7EsVfbvX7l9uNcfbV6zQJGJKj8DQzS/LV0LotgHldM
AW58pCwuUxB8ROkHkMqMkMqtGCzxcZtIqx7Hr3j0EjUJlF7oBoI28W4uKBpZ
+qmI37/Afyi2gUQvEbimO+t9V86VYeJfGYy+pvF1zxs4f+c4cvhUZZkY2zH4
tV4st41hthBQDU/II/3DlX24Vx9kGAleONgiFhEFtXR6pMptwzF80xtjO6Vt
xSC2bhn/JQQWcwkcnf/tOqxXyQ00fHF67inGDxyUkVDhtB7h/mwkmNE1Eno7
74Izq5sZS3/6r9aWzZvkPH7Ug5LJdd4mgimbpguKTfRIYNb7XNkuAUkbi6gt
rp4LVd5iWt3w1zqhS8u3/OUeiReDrRtqq4WNXFsfrJnj8OmbWfG4PPfppB13
IfN/83dOH5AYgl5S1p4pbjEMMMF7QXR7ng+/NyoPG5RQXTLFJsDyT9VmcoVO
9bV8/aZxxAcoCTOm/r+54pUA+jG/GPOl6s2jS+6hXo/xDm2f4q6H3hgu0GPD
o1eQ5XjEWo3xrIq2PCu5sViRduo7bQAs2D+e+Os7vVgyto3Xlv+f1Wl5CwC+
sjLWTSlj2adT95XBDhMy1m/ozJeH++36HsKlj7a3hncsImzIvwEHrg/++DJ4
ShSFprYnfPxxOmsInHHdSyidrPn4ptlHtF33xKt+PMrttOViQEtKtWA6rbP/
RX4cae4fWN34K1YCNtBkMY3dzJ3EalbS8FU1lwJwjlRuLjOQWe5VkVRVDv24
TB6R+QrkbN4y41P1UIrhpEhCQvKtY8oakwwUVfDsMEQCKYVOKtjtykJF/qby
Vq+3HO5xuE0/3ue8cBlJoXBDXxFeYksDsIry6m6N2P3Bc4Qj1XEZ3J1cbiL4
tYmG7Y86u/cog59+/sQT8CVErD3apQaqF1r6haGmQ14N8S2tjvaxMn1M6C5j
KiHGJxe/rCJnKNty1q1gZ38L3VP5SUe5BQx/WAciA9IRxHchOpgRQrAVvnof
zrhVoLqv36x2zvgB6K3DIQawULTUJxd4YvESGJT16pBWmFkpVWXRqUQouTO0
17PkPPvt49TwBJ/F8/GspYrqGXL/hlToS+aH9//0JhBN4uPvs+bTXMxdC5Dp
YmbG2kfddSsPWlploXpXFv6cM5dHQWqHdmZDcSCTlHqHcOcahNpH2F9JuQp7
LBBMW8QgJwMBlGwVAwPooo7/QFrVwXEdh7ZqPG+73Ft6FVx7QKH5+W6xe8eO
xAsAdGzztKFgz1m8CJStr8vy1n+oIZT9chUJih/3++FmvKZ5GjuPlNV2tQR+
QU/7u4mcosmthNdXZrZqUJNT9xbXMWsggPjNMktYLpcgslwd61AxjdubRyHk
tfs57PlcDcSFCxBuk1VriC3gRhcKlEfQt6/T5BS/YuacK83q8TwRVtom1Y5y
rkvAYknh+hyGV6DY1k+Evg8CdJv32rR5vQfgdDviIgiHsq0PBcGz3Rm+pnwd
/7kDeRSDsFOeooTPQo988cRUJP/VbYTYcRuoJQd9940hXBv802X90sw+G9fw
ztojPEuibijM+JHMgX83t0DJYko/lFO34Wzy+aBrRgN1Mxtqi4FaNAw6FZgk
xIPErxixvF95wbVNu7ZVqeoOyFWR4mUMC9WH7jKvjB9/VKLsGvV8X50JF+yr
GUL9IBzjTamSw45J3uw8gIrbtg7MgAIwOsWkNH709R662Xy2f5vw2A/cR07v
w+OIIXvrovbKPDUMY+IW2GnN8Sqsf3LXCqJmlAds5RnigqQSKiwxdGJ/ntgB
TJki3E5i9URfPcpz0/V8IZ56SlJIkEiIalj6UmdVYT2mGiiohr/ApkuDptvq
jKGkZ8dz6NniTeMHWhmQvH7C3QmQkPc0EvijCLZf619ciQYFuxeBLRCo1OmN
yJdrwJQ3DSJ6uPBqsD9Py20EwUWJrdX7y6FXY2l4fGJcerVCaEPf4RcR17UP
KE7R/Ht+9j7Xm35qGMtOsMe4EBtxDZMJc882H8MTwieuwQkUcbiwAQK/xhAs
VH/chFk9iHgOlko5BvNF/Ovzdd21WnlQblnyXO8pbp5ezgL939bJSAM4PaUO
Sx5lTAVfU0lwz9VTADKrIBy41hBtP959tX92yPv3LoGi2wd74ni9wyE9Pw0F
Np+WYveMQsjAceX/9jAOFji5trwJFnfBpM8NmhhpGxGjNjUi7W0EvsVrDJbj
hHAISWeFa3eDM2E6wmpLvtrVS/gjfzuc+KuN+JMNqXawEVnho48MyPQ5oAqz
Z84f58i6PeX4MQNZLOzPsDHQzo6188qLsxWW1Ra7g5u1uE9Ixo4iqYloTXxu
mTH/GT26ZDm9Aw3YzZcQr7oXYBx5rJ0NoPfWEE9FOWlebrBI4ac4gj7BZNqF
RBFM5mNoOQMWYAKKBwh3DvmXGw6yn0M35zDsdY+kruQQqPIZFmIHanzo+4G+
dCDVDvk54qWfp9Bb/Rz8n+aIWb9wOejJ2OWckRoeO2bwqJciZPv4ggBRwCVs
YCOKxwg91ZEEMjZ/YZ9CJXeATS3N/qkZDWllbKpteASVgFtWDMTm3fg9R46p
Dikd/RU4gcubEa0XEt1JPsvdAhmhrJOgJgnTot2IH1diPfW4ZhVi9znPyoFI
kVm3mNAru81xnmCPjmGblSVhu6VzAssTus9BIpf8FtYOA/UBT77VCvIvvP5C
3rr9YJcrdWpwCVyz4ECQqoLa9BJSZBKR6Ta2mV06CSzCzksJN1G+5HWsVAq6
fX1gHHapI+XJJWFKvmFStJV0SzMv2WgzvVesv0sa1FUCH3XMSNpky5ZxWOFk
87pGwFeF1VABUPtR6qhAL/81JuUpSmiYq4f4vTBRxh2trLbgHfshaGkPzh1e
Hx9AeDMB4aPQ/6cR2Vr90mOjOR2WEQT14tHcNAs6F7pS0VyHXNxWIGf+5zBG
40Ul9akqYrXHjr99mTZLEjmo48zLQiJ0fuvq5xoRA3I+COAPgmKm+YRAABwO
pNBppr13R5VsUAuNfr7Ps5uVrsFgHGtiDTi4lzFCZtEC/8+7YwqwpRqnL5Wp
YOk5AtRp7qyxrToWgOy4uXgRavi2LcS+fXz8QwThrmyhN3ufcfczC1zLorhW
9eTpmU/Jrg89iRWVfZvK2t/r3gkJkcWOD85LbAFK9ABRYNV+nMR4PJoP/qXb
5+auX7noXBLw1aBxKH9I5/Vgi8orSwY14Z6C2RP5TEyN8v0L5CL1wCyDkSKB
3TEB4b2AlYoP+jFyWiEdPCuCMil352TwKV0jiVBuE3YEdVwxj9m+VjqzjbtA
/bfIrha/e43T8zfrBsf09zL7CDhyA0dEqxMJTD5aQ6LLZfoGVHzoY3TEkVXt
i0PDEJo9PqdqW1hlt6/kwnxQjsKP8/s6Ti/HNFohTxbEIA0sF9ul+nDvtcCJ
yES5ikRsxFZfqQF/fw53y7azXMaSbIpJgq3mS9ogrCQaYkC4INxiFRy117Vn
lqje1TzfkxSunHBP0H2MaSrP2yAtyxI9S0Up5Q6vdWq27EoMxmNAlIWWo7x1
d7s69gkMGR0WsWFuyfCMmqkbS+B3maLmi9RrAF3UDDgLPfIJaOo8y2kw6uKf
Ak/q7EqrwbQIz5LR+nGWmv1neStKVcGnLXJ4/uBjyoABgqIPEbWEhQ4g3Hit
YLiEC7F6s8kWjtru7U4ZgkUzlhr8/Cl6KuJ6eK4RaLJZYNucEol/TK31EDfx
eCVbT6RuY1E5zzdTJdxyUb9OuitLIaMCNnSg2aCrP6wGKfjTYV9W5zNJd7AK
t2t81E7D7zS0ElRdDXvpd3rzWHGlFR1QB+AbmcR+JXQ+R5/0yPEBEplC6p+6
bxV5peEI8fnaSBKedqY3w06HtxFPcMVMQZYC1RmlIPHdt691CQcSPfx2+fQt
ad9v00J3mTdDkApjghrPOqS0wZtZFveDu8LWAHjmdvfF3JgAIOheTSCXLdvE
R6rccmFH18NF84YxMtOzgd9pKFBBXBHGv6emxoOHiKChn/RBkcwuDL0tmJQJ
3rtMX1TwqXJiTN5rqQrL7aC77bxoghI+70KLcnOARSSTazR5x48IIQuDK3h9
HFeMmdi0u//ERMGJqvYhS/v8Ug1Nre4v0ODguY1bdiJa9dZJwaFr2x/RIdzN
G2ZuLMY8wru7Bpr0Il+A5o4GgAp+dxfdVat4ia81haPlFY2ZRRCZaAbY9WMB
2b1h02pYq9+s2/0ZNWDEvjPQB5y9UBYwsYCYl5mJOCl5MevkcW7efKjQnsXo
HzSfYU9UXQx8aFp/Nw3SJ9DQeTIaWN4hNXCk/PwrBrZq3N3EzYUhtDHAaRDG
/IwJ8GDMJs770Hs0/YITo8UAMAg2+j2nxZyFiOBwMMxCJJvgety7rCnM8su2
e7qfpoJpx714xMTVLlx9M8/kAhMSKSgMVnqgyGxEEUhs1aGLyetmRPCdKdde
lT3wnmyr6qzE1qWIoBTTcKe56hsZYs1di25nomL2KegPfBFrlFLbSD+5rtzr
/qL17Q5wamhiHOY+SFg18JO8nNDZMiCg78VvodW8XuPeVVdnjOU19OUFF2Dt
e1IywHdcy70deKj4yN7jRMA8IN4emrHfAhg5qnB3L6JQ4pIti8poakXR/5W3
ZgAYegQC6VEzNXEtxOghr0tmCVwWwnPeKVqDAyndP3sy0x4SkjffE/5Yfyzd
n9yEr/UZqZDkzc+YDFBuv9PnxB9t/gfMuTDa/4c4rqqc+zBpgLgT11A7Kg6u
eV+940Z17QPn51kxnLJ0xutBjcD4wOBm5CL9hMTQxA8vj4bZokDnwcDyjYtM
dWtM+yGT+ce26rium0+E4kTJ8ntp2V/H1ykPgR3WjxznbgIIKeP8HdVcadu8
6OuKyOfKQRceS1IN/L6ZfmrGDgbOFSxMODxHzU+8WOYDe7YE9vpAe4YbcA85
7KTr6M2T+mgTBFcJ7LFYqV+dP48GNXuQW1oNoLSf221Y8MqZPYS47v88GWfB
mrZVMRiMzjPlyuDjah+NejKwos/jU61U0GvfeJroduwjlDSvtYQL5d8UAiNy
HESBapTiWVV8ZnSV/Ce3DyK9jvpYM90QqeS0YOe8IYfN1h2H5pdSHvNh+6PK
UstOxaQLLntaBHHHporwxeeDd1HBlcgkkfskpfRKqkRzCPrMJEoJ07eu0F3Y
7vwiyUB3mITfump1/x1onjphZHHNTq9JWPniiDcWvO+5LAtlfqlSiscYT3jz
dLSznRbwdlulPKzFdpDvo4iTDoTDxwKv4xaWhaRxIc6tYZoIeEz/9it7H8hL
y4+JRrw8ddW83zieBs94ATvww4/LAFf00UAN1lDjUk0vFdvprtj8mw8ghO57
QjOoRSJvIGx2scOv80FguvBOdWDQAY8yXF3oy4quM4jhBAtMUSIdKoOwM/e7
jkJZRwYiqIq0Sl5l10fHeqZuQyB4GIYGi2uS3NgQGf6VVD3yHlV1c8Mu827K
TpXr8AHe3/7zXAT89qEZGfS/RYOLXqzHtYevPOv3/RuBY8xiIG2ZhcGpXs2b
4Njy4IuMd+vDLbloCYrE48f3pdHZJdP9K/gE8Zpvp7UvfzYslJRD0FkmM8PY
vAN8vr9ZNsU8H4FNbzrszicF+ffljWETJHDKh1Afa60druA/t5TuWixGdL5d
/lQNLgVm5Ga+ly6oWxEmkgkV9Tnz5bXbHNn22FpeSODoep9WLbSAVkmP+wrK
J9PxriwaM4u0WeoTypWuevrfCzgbg7XEYBT6uOO2CRyqs7pPNA9H5m+oJ6FA
qrXNR/DV3lN/ol0hnCIl8TL4zDCSkHy0+tO9zS1qQlhzF7CmxbS/4kbPFE1V
tSe8UyCzmDmzDXFh9BfwBFeBrZfw4aPFA4XzppSl/j/1+NTzT1CUTz9VMZWA
VRmytE9txXbvB28SlvwKlXt6GTy9sSo6hJYK22e2+WgtdCtGpxG2AYqaiZQU
mQL4jM0NPLp/++j8YcPgWOxg1HZeRvkrPKsxKO4vUU/2JKd7q5G3TLtf7nW2
kDJA4Yp/wDmYuha3vw+4jJH9VUXbbtWuf/mNzKasWG6Gih26Q6AitQsURkwm
aune25Ih6osvaPQmKjngvk09jSBePYnsnSaaceKkrZQH3OT5XgWyTca8MZt1
1sU5NE1A5oJQKPkHPbVaalHIhMh0FwvRn7wgNwJvNdBn8hQJkPSnDVTvuPze
H+Ep6UgSSxubQ9BF+gJScnVbXQL2mYv1dwN9vtfwZ1qkdNAaiMj+RgfjkLZ4
XLiccRrTZui23AvsRUDbKqlqOx40mzS8EntRp+p5EvxRjvmh4inta9S3DBOv
7G2wxosIZ0N+WSFW7kag+B0cAJ1msScbB50Uhx41b5lBjIK90T3mTN+GTyvf
g9cNtivq4kglfwnEI/lCLNoyGdA+MJ5AeZ+Lo6e6BZykaRi6RpzxtUwxBGrr
mZ3b9ceK9ytJ/okHsGTtAz8EVK6En4jDiyRVgMVtWTbc3QWw2TdsRpT77jO1
a0z1Q53guPeFLpKzTmeCL1ibn+BAdfMKewJIYm3CUWaO5VlYjxvRLmuqWITc
jPibwZ9OV/prA+NIW2ZuaZAUizy7wMqrWI15GGzE8roao4oY2fzvnzuJ8FgC
r5fy1p3p2uneJfxYTk8qBJQiwKLvXpghU5zWCBXNFydT+LDKGvGy7YAtTkQb
veYjLtFvm0wn9SomzjM043fIB4K+hVnoHCtgCUU2f54bDSvcJPTUGwdLcTIF
VoPNiYpyX7/slTOqPBi/qBAspFw1IGc/sHGMxq6X+HBqxS2MZEb6/VFDBgPI
SPr5D/dRvFauQUN70EUz2BPbmj0N9gl4r4PFIKzQebQw6s+SVZxtDZ9tpd7w
mSkaKTqEMLBVP+9ogF7B8CF0HiXJbr8sHo1mot64h1wfp2bS+pX5jUf3vwyh
7J0ZcS24tO8zKtawoc+lH8VwJB+lJvZmwTgrF8I2f5ESN9ryGBaN0HIaVK0F
yfdm4buqdJ082j8S481x4b5Di4F6UWVoDzFLVaeGETpepsck4BChJNKCoWcJ
MeiXSyecjN7mFuIyrg0dDPCwCz+WfU9Ksj2nLFQCPL66OfZLE2ZYZPUOfLtY
naNdr36J9qXqJXu4n0f8gEwnBLSc9kTZ+LkWTt9lxbq1rwfPERIhaYG74o0X
INEVS5MotgTDGTyHusAib/fAIwT/ZUU3/FrZJDZgKTvsUz6nKsoDlZbSIEPN
uVDtm3QNmpdvHxoonpf5j5zwkoyX68/zNoRtBZNdh1QrgXdM1lPi5jMqSmp/
EOtp63Em1A5TRP6b12wfQzOujo3F3oBsLWmQap9G04TbTiOwnB4V3BkIUFAz
tZHu/1xAE8qb8NGvU67U1KUwL3o3kiwcjd00O5KaWcAffdsZ22u6eGzz/ohP
REd8vRWYsxJhbFZrL6D5hTqbU2lIGVU2a/3/yDryJjcVGZtZ9N9/uGgbsn/S
Q/B5cbyfQUitQ7/G2alZ1uvR9TDzezMT7dZO/0vSiNA8S8v91ukHBf/qTmLy
EFqcJxZ7CM4Nq0HfekeRJ/5VEarAZqD/g2tPjvBPXy24XhTHOX3fYzAW0eNb
3/V8AdUoSb8jlWnu/1XdxZS9Pt69tbpdF1YFgsg4/v6iMSajX2fedISM8XDA
qbJidd9yjwYbUyVzjdiXmEO/cbmUYNaBP0Rlz+9jyBGoC+5ZsECgzTiCH/cP
TrqOVsdfdIPmvvvqG/u0CVmDc7kbEOetW5FrJOluz36VP9D3nK9bNggnqx0C
iTVAyBJlA0W8Wfb6jJvE9U4AMUq7x+bEolLec6N0OF4d614lWfIyr4uXeksd
on9lrNOe1sMtG0mQi99F+MAl3VVFaYZg2HgN60v0vQee/nbHZU7A/sju3Uau
RhGDDcniqicdjSEMaXomkx1iBUl2PcVGXQLohVkYi0OA/HgRRHFcbe0C0b0r
izzTa0/WFI9Z0pPYoeGKbJ//udtZTavQSK1ifRbZuwfawHQd1RM1WPxDDPPY
jwys+STSuav1kJ9MDmr7lGi6fSEGLOcd1VkMVPc3dPVTCwcop/obl108txyg
xTS/gIEF6/b5vaALNE0SoEDjNst5iX5uIvHbwWthrcjr9M/ILw1nJ/T7Os+e
BrNuwn62+dRuyXSgnxbUxOt94oPmoXBUuvG7qxde3gmvzzns2+nP8XLcO0Uz
wPi5JRgYdZv3MIWDxJHUIaDrz/wa0vBGsxtHubXVe7+cSM77zMCRlCnszAgC
ylkjYmhk2RC4Oh8xfKVBvlaJUJcIA5xvy4dK0Jtlu2Nwn3lo9/3I+fxZkQnM
NaWBCLut/njciY5yJgEpLcmjkRrVhXYCjovJOHwwZPLzEI8QkpqWIQvrnb78
TWAuHeHU0nUmRde1hlnMgYcRItmvdL4aXsjdv6OV2Vpp8mMlm8wSrpw0zaHI
+990l1gn7KeXaSOtDQ2cu+yrwEglsRb8R3gsTtpG1Zrmjxz0bml/HBXvJfpg
3mRT4aRUjDxqlDLI+XYtlI3lZ7Q4jBbS9+26mFtW2DAcsmMMktxA+s6VKa3g
lK9wExNaoBVqzezhmtcBrvhCWeJRU5rM5HQw68fYGVJFWpw9M/VeugzD7vQE
iVpaS/UoiurzYzoURROIDyARTL4F/W4t6scwHl27HsxIToz4oCpuxXypfe1C
bkkXqBGUxKZJ938LiAM9aS+pjJC0ffccBn4swMWLkwdcr9BTT/MFjxWg9qOT
UYD9Mrit/AQp8AOqeWXdgNHIs3veGCUkW6Xbj2hW+wiIFP9o7MILv+ynjmtE
0b0MDUk4IEJyaBLiLTQugMOaPe7XWuRLvfUtqwGpzjzq9S6IBTRTVztOhLCI
M9tvryl10vn50moHFPYC/OrctcoY/s05tbqDRblHttW0nUCuLw7S/8plCrQk
oWYFovs22cSUrt4CBeNMiLydKexCJf6e5S490WOJz7MEcNZK9h+W1Ds59eC2
Tx3OhsFoke7fZ8OIb90jO7L3gV0Yaqit2LGFm5UbpqJHkbmhvOWvZRfgdXL6
yCGTb1uIWVsZkhtTAkgfZB/5VrlFi+xuKD+pnFy6YIy3pEe+1eo8aV9OPopD
8ZK6lOFXIqiLeJuo7GayGj+B8AxzujJ2gbAknrYrbeU1FJohv+CQ4LxcSLaH
jJv9nxBKCCGQGHuiprLo/K7+jo1GBgv13qd/fJZgzy+5uMX8cQ4YZ8gk8yta
XK6T9bsclEYC4PBCKP7glaRSH8jT0S2BZWf1fDO5TOq8HZDJOWMuUxCpqf9m
JA9C6nurxGReIi+mXVkyi+k0O2advJ8HkPGxrVT0smf/5rNuWGBB2oiiCnPw
SSvvSf3BBZ1ilJLajC209gtMHH7YOj4EiqdmE/bF12q4wLzODTkyZcxhOO18
jWBXVITt3FGYlDhtCMETCmzisnMeycaaYhq2koSdvUsIYANQm7uiQZPbuOHs
dJTOWZ3YY5DA9f7aXrVVA80kHfkBCijNlK7AKp5JmnmleTRooeMn5plUZlEF
Alw75+D64Ie8EirU1cOXomW6O9rq9Nbvz+SNjzMd0LR2PBiI8knu4q6bXhWS
Zzy2NzgDaCV5nPAwSKk+Z+h+yqOCwbgNl+R5zVdZt1htcZfcIFl+iIx398J8
ZwzYjGCcu+uu5ewE3auau17jeuWI4y0SUwYKNrSqclJiONXe8rBKFq3LOPJA
B2CP79AZyNVOgx18s3evFJ934ei87V7J1CjZx92Znj4hhwAl2VkvqdCBM4lp
yOK3KqHfV3eA05HL6tcBwBHrfxVj0kR+qYam0Ikvouvs4r2z8Eg1d3EpnESf
nlvsqiK3Rcgep39kj0XHg5GW6UF/TmxuKJR+rWtTXe9v5EQY5dIyxwpSys8O
pgTQPEA7kU7LHHxcMB4TParMCa03Y3EAd7y1xyGJTiSVqLJNPEQjlKCuCwI2
jD4w3N9hV8Y1Gw3vcrYgmjHWv+BI/kPl0oPTDUYC0AR7zZ/N4wBPfk2cyYno
DfFuQSZTWKwHnQm1epc08MVChXMKfvpLa2yRpOoUr/IDoi6LfYVStV4AO9cO
Lh3Qgmc2jEoG17v/0bjJWJiQvVnJ9kUONxOnkszhP4yPjbSCVa+j35OfjNQh
koOBNX7KRMczb/Lnq3uda6COJZWn6XFE3lPRkc7IHGivrydL2eqARGNOH6bl
k9Xq/k9hW6SVfokETrVLNuuHP4eDjPvnza1tWmXBD1uZyufZFMepl2EQOhG/
6CL5G2tSFdCjlI9q/atqcwyMoxiQK7GPle8JERB2WiJ9nvv/62JPni4G+x/S
3RfgS4SXicjd800n6jbJWEKwRtHUwFS3H0N8AwG2yWEkh5yg7/Vu52PvFvmq
wz00hIi312+g+3PZs5IdWhrZA3DFRYqYT7xb2yI/A0D6djfe13+20Z7+eqAb
BHoR0iGAuuQTsmIjlMWYbdHRXpfgrygfcIZoR4Ot2A9ciCKU9x43EcP3HWem
U1jKzom3dVTsWs9NwS2oKJuD05+J6ISWcXcEPLRFdPnAIBgObvwH73+CUhMW
7dTYU1KTtrAVBWIxmg+iG7Thl8NT1X2kfuTErFnkHPIzauZgegBxWPU+Fl5t
FCmQn0hDCbnxi/JQdiAXDd4JBc2gz72gfc5dB+j6I/7wbEW/RC39w5Th6gJm
ZiJCTcurkArtaeUfvZXzf2Q0+/POyXc00nI7iKjiVHaLdgl/a4TIPGN4ihaf
bLHRkiQgl9DLQChT6Dlb2uFvrRjAa6uMFzxKxzp7wyJZ4jPNO9TGlrfHCCJf
HMne7wbs+yZ2UeXzz8zgn9Q1MyqCb9Vfemzx0J//ZzFdud5u7b1kjEXDynYq
Kd1BUB+KGTOKE496UylIBkUN2gnUWdyD9S9q2qnQp8yF6czvLYaJqda9Optw
Zfzyi2xb3eYqWsl99/tt5oPXjmDuxKx3FEVLXQdWCxtU1jwQoRfofH/8VnsZ
Y6WdvIkvUREEmW4ZNZs7PLdmwtoyolIWyELyIllfRiDRknDUkd/gYpu4O5MG
gQTJcsGvx/Uc/FtsUhI8I6rHo/fiZcM2hZ93LyPZNrJJQTnH7aSDGkY9BSfs
G6qV/ZGYWynb6D7/vNUSCw7Hm8oiAiFiRYXFGdaZj2GNyXyqckus8MJloI6y
klp2ZekBfnnmvtR25/3623Owov1jbP34fUoOft7tbe2vcOvSGgzN1mdtISE1
L/4YawXt2ZhPe/1wYjfbSmWWd3SqtRGZVNE+wKdrbc6NIi0y60b6+iLs8dkz
dVnJ1kzxxq1fWbZrEFvi6O2+ooZ7mn6OguY1xXUMxNXZZIC6SFqX8q83JqXT
oyxuZx8zIL6uiN9W3r8gnfmKQnCGYBkQXj5R48WSOO4D/6TR2owSxm+xBB0O
CrWSHLCqe5PCTNG1o7PuSbUCC2u2uKqJ7u9GzTL8FOcms365s3WsYgudSsyL
wN2GiET1FOeNOobKk9zMef23LlHfglrBsRr6TDlnKgsENZrqiBaSc9Z/h5Dz
znkLdv9TxZuc45vb94VPqwNbQabr3UFxiRYqeh0C51wKattobS31f59FJElW
qwZwGWnz19hNsEhmRmQ8GBZescXuLIPsdizYA+JETbW248CdPyxeaoxZRSgy
omZWGmOcYUHrHTl+FhDHZrghfaXO1BeUO2UcOXM42wxWvY90Gwxxu6RuY6VO
7iJKppEyF4165vr8W4/8tlDXZhHLU3iGJhBz5jyIhaE3PK5lNmDwB13OPChl
1fdXLt2HsOPet+PTIRi2E5tKU9LiWq5HWg6i2l1aeinChuOK7fPdDEpRvXkY
gP3OZ/6TW+XjREOlV6s9Bop5XgqoBjwhtk5M3kbACwwB0WItUGmUzH95Smfc
6Ia4iBL58DwTKdh6qj0qPBP+M5HiJGYfZC1eWRdQJwFf1uc2jYgEi5MZw4Qf
UExRAJ11LhAjR2hjr42r9prSjRbHi4fZs5YNMgjDbw3q2k4srOnWfrKMGIXK
A5x6QSh2+aNJT8IdqNsEAzQ2yy5EgZvfwDKs2o3/aI6aGM1ir7CSirrCXW95
zObf5P+v6Ywh2WW3mwRXbfc0xMH1eNpN0cr8ApyL14hWui9Fm633r5PqOjdx
Fe9oHtOqEMVSrD/8oquaZoj35tT2EsbKq33WxJaV5D8k1/1cY20w38MVOYrh
qIsh93nPAjJ5r7vHh5EWg2qOPOfPaKB+wDQDHQNj7Jot/9sQNvavtlYVgGev
5dyno5Xo8LfWY3BV4s+e0G9g+i250ngXfrCZ9Y4j4V9//RE7rWJ6gLQwStWK
ZbyuOXy1utFf0QqwYmBLLg7T+VS03RwwGNVQY6/Dt1JAUuj5XJJEZS7ZVl5Y
qJnI+w5WxHDroeEWWuaKLGAi+ikqNkpO/KPEPwhvJjjvc8EmELvsY3EO+r9p
/NZMbhSbPEjTsuhXKukbcup0nGt4PzIWksZvR+lNeeZkmrGxzJZJD1pTMRZg
TgTYjN+6VkbeUraU/+FAmqb1WIcuRGYBgmnN+6qd5cDIj77RE5eykmXR2qgZ
wlTwE/CPW16Fx7nwka6aq4+Fu2unE9ucbxnFA54rewQ5DrKW5YhSKjdJyNCM
6sNkCHgRNGuKApBYUqgv7vk0INuZjAlLJjTMcBZ1H/uRlIU8h9Lq3Y+lqEl4
7KsPM9rRvexfoaYdp8q4n+sd47KPI4M2fzHTk5nc1otQ5nygROiInu8EHnjX
NJc/v4cB01dEExLY5EQhJIazsQgfIfsmM0VKYcxveZNy2H3ehAnGGuc7mwrG
5iOBBzKYA83tgjXDkox2AMr7gnKVF35LEmM7L2XRtClbzp4WhnRQiVqiiw3C
R0WRjsW2fvlZ4PyApzXjPlE77XVB21TjNEC0t/VkFuVOrseWAgbEQu5YY1LS
x9RblyY6GjiE6ruM/zrs2Ys/7TskpXNm00n9JTr5KMSB48lr390oQn83OBU9
0Op7AWCPxdPlMoipA+yonwgkiIOTnyLxrtow/mwbL7PZPeN+HMue/R7Kq1JL
8K6bymGDq5asq3uucFi7d+TQRMsPWA/lF+MP7ksNZO3wxmc1tTKKwkN5TWh1
x51UISx1EPWoUNxLLXOfXWYR8RXloGXZU2ndPmvgP+jw4Uif9dN+2dcAk/OS
GlQGyRRZ5KUCrE92D/XBmnDyV8E+xtarrlmfcYbOU0tpVEMhuf21p7fgasDa
/FGnEEb2abDms3eWkVpCIGS5TqatYurTvQx2PDj5xkYoF/SLYNXvi8KB50Ol
fz5wy0ZDvu1SQo1+PWUC0uP3HOF5mubQiqPTqPKDf2xx8LEyxh+QZTkvfYKh
RxlEAQPw5aargLx3DV1CL75ZTdLnxzSG2MbbEbcmyKXtLMmsT2LxcOUxzm3E
/+RVK2xYXe6xPyJNObaWPUOuonUAWHjhS01Kxn5HUCgsxov62rm/PdKaWyIs
MLOJLZAjJtNHog0QUwtyQPTAKuwUkvCXJUDfXIwnJdcAsvYe7GkkaXiWMrO6
XtW2WMIDaJl3OLtUMHgs76yMTy8rGnB4x/DDEPDjbufc4iYvnh/Unf9kwAXd
RV1zSnRbtYPjB3WDB5bomyAj3Ai+GtJD+6puIQ/HJr6TcLhlgYxxoAt/E/mL
aNv8HNk3tNX8DpiZYiAjTUhXtT6/zYxY43+LcGLjWmmjwxmnw5petBuHAocq
uD5Lhc5bRiwjayAGoKvR8QQ+NMYDVGFjlBKSK14VO7J4ARH1/xXIGTHCJKO/
gHYe+t3p91uxtJ4d6iJq0p10SYEU7ZD7MxuDaBib89UaehZZs24pfBOLSRUw
xr51c3btCV1ygao+Sc8lQ52G4jU/iN7L4/VypY6yfTlKCEvxAKtKGuoGCMX8
/Uy3VCIaWxSNd1fUC+c0TqNdwZIeVfmYIqg2ahKg7cxudRGuh7lVNmvXyVl9
Ui3HGaSa/5BcdMrcGF8bhuZ+E5vejIyX/7syv9dnF5lQEAwMXoldHHElnWgp
Ia0XhaRtS/HI3r+qIf6MRpDt9GxhuPjRA+P4EqEc8DAcKzYH6LeNC9i6pmxM
3R5KvXPlaEygYUK5ybIZMO0K5YtzRkSWCIa2WPJKDBMTEe9UVDIuJzsszxy5
tXUipYlEWRG7b4QNya7+36RGL4HAWm1f3EXXlDahcVp8M3+EZtcHFV8MfxvH
MYqMekZ+Qeulsh1VS0gkIp+O4NKcNE2itGRa4Paok6oWqQd2T4fm7LSh1SjX
ZWBDzCi+yihh0CBw2SDIXVvQ2E2IuEDr38OD59wRLri0q0LuxKdJKwyT6EQi
FMmBlmeO+UeOqjSBI1pjlg5nubzeFIwfd+0BBZLfQvGjyWJrdKRDilnA+Jal
+5ZczLQHcLbsFDM+m0oD0XubEVF+SfF2+aGdMpSfyeAqQMRTYoH7wyY9BiBs
vguvgFA7DiW9LpywlCvluNOlsnPd6UcrbWnuXgRqbQWg4ydU03Ikj9Xlpyhe
epKxSaWu5pa45ykDFP5Yyxi4sHA3AXWe8WiwgAJ9FDn10tXAuzdzFQPHOx5U
kLIL/5kFpAkW43nEW8jU1P/I1K7mvIvFy+SpEGKTscPGVFCxtkbPbh35Eyqj
WN2TOzoEC0euom+e+p+/I/vFCFOYDN6B9JliZaGvWpI0lcDkvZadxA5kaGNp
sQJGFm3RQUcDgW/g2Rpz9CQQ6DZieMS+Turvjs225OatmZbQBZCyf9hqT09j
FZHpezrIrtbC8O5VRlOak9BckPzzu36hnGqScztlzXm01B4KmXWlDnDoueWt
Rd3oNmDMWsW+XLUVB7lBX1gwDjXPTBLy5AnAUbHTHItAF8VQzxnBaJudsfx0
RIXY2hKBJBKNeFvNtj7K3O9tiES47Vcfh+62zygdYsaeqL7qt6ITpg7hOBGm
qIcNpKE2O9kGe7UZG7u/sTKogBA7PW+M7UoJPZ4rV4O3hAwDVGMImwj0qpZz
jhdQ2XLvwb//Ln7SWkbCvL6vP/Pd9YKL2RWwMOgvDAgfyH7+SQkoztvj1IAw
Y6NplmVCIt2wbeGkI3xgfncDFMetNcprw5oJ6Oe5gf8lOIi95nJdhBhuAB4t
Y1cChEXAMT4XsXgubu04TEHxDTwKTuqIqs5HKW++D469qMzv6+CFPA/cLG5P
BVvE8pB7XAqiYwuWHGuSVabC+o23iefyxMSIajynO+rTHWWkc/nYw7n6WKYx
HjHBrMXiviInAA9/XIRe4O+GVTCChl9gtf1CYgTRxkgxLkn3rjooaRZrm6B7
G2zCxBlSGh81M2fuCQ2HoV67AFjGcO+vTYabSBmN59AWmLzp9XWrxC9c9rLI
ozJ7ehDkIliD8Jpq7qKifeJ8uU0Hq6+ikomjsh4GZ6WqQRUg9mayqH23m6LZ
zafjkdIuLcqr+A3oc/GnL6MANH8WNybxMfkTGgpHoI3Jy2q0naI1YkpsbS3a
M2Xurj5ygL+hDWs9U8321Og41J6fMkyN6BDjdW9X4Wt8d3dYFbh/mt0aCoOk
bVTSIvbI4B6ga7wZPqHpopRAmSuLQz8U8zGTdPxINlDhHXX4Na4qvd1kZh5o
CE3Ay5ThHlD2WZaEeIYq94/OrGgKfB2PVxQOTRjB9nqSb6hrTgPMg4vD9m31
pprz9zbfJS1nvFV8e0bX5co5bKp0iHFhfXcEFNGVHYyVIKh8oeby0+OS5wn4
QA4VE5TtXWrcGMARfF0evQSUNzQEWgXZRmT2IOPJxQJFQA9C721SZHoqFchE
sRrMzBnkd7SqiuVQ0z9jfYfq6pbrgJn+n86aPlSvsNIa8CzYyfZSGLMfjCC3
Pfs7dBdfNFiIdBBv8eDo6cbdLgFakV+gLnXYDjoC+dF8HY73ZDihYou+3GgM
5qmvMSmRdIsHcnDIWkJAbS5H1D9QZb1/tIhH1F7sJ2Zksj2Zlv47+NrO6Bbl
6tIApSIibcB2b4jRba+MBvivcb5rlbIA0OYEQlZmiN1kMdp81TiXl7GBN666
AqbqdptDpMSH1qwMjoD1o8e1ff7HXMBN1VoqCqWJPm54GycTaPED36Yek6Wo
yfD8jA+VgGb6J1zd+FSLzXRo4gPOAzxwZ50lzN1lv8NPiWzqMFDYb68OcB4G
OBTlFdcs9O7PYxBP11hFSBB2mAhDw133Dzn4NNvoQTBlUkYsZ/arNvIh0j20
WLbeEboLTH+cUlBsVf8nDROE8dhX6Z2XApin5D9cfZ79L0Gy0et36ovctwpp
SeS8aN/J55YyLf2i/PJi3LVaM3ioME2C4PKUEGRXS66Efnel0hDGbOO4k2+l
yKoXtZ06mMlEDTM5C0Pe/WtTCcqVDG1iyr8qKvy1EO7ETu/NjlzdQkFFb+Q0
hAwnL4nMlj1zo4s4t7v1da2wxWjmtjVNaE7Fn7V/K5PONNHHC4Ajt6iCl+Bz
qR3azff74pGc381b53+FQCqCETUCxWcU6vSbx/Gu+HkKsmkSUhecclpmRvZo
uRzvlOQCOm+LsAq7Ji0gL5SsMPaJHEc2Xr2a/iJ8nY3YHQ43WVT3uPP9Qp6Z
qiXdXkua+dxb7hmJXN2ju15Q8+CbYxEa7UmD+d43Qq/CVHplol5oecx1cmIm
R/R+uGrRr84nptHUtkfqAIjwj0aeKRKUzNWSImy/jVR4wVNMFnTm3NtE2ieL
iySMr+LZ5lmJqQ9zi/FoTMHXOotUb3AB9BVcwvxxzg9bJ3MIs4dB6KrUot9+
2WEvufuzgl8YhWenASuw66lmuN9pvuxu+Vmb1NLLdugDK7/UCOGzbEF2k920
LmkyvmKaSvrh4oA8JhF80g+AssK+7jA8faMhEvWIebhMcVzmwAE3t9QTJLm9
ERn/U5AYglHUaxRlecUTViL2wTRCO2iQGIrE4G9RMy3x1yM54X8ipbghPS6r
064kaHomBphjot9IjK+ONA/Y2kxfMaPHxyt65pU7InW8Qmz61lFV4BpQarS3
3pdROlIt81rFggvvTxQx4qHKmG2EZeTenuzFjwdkZZmZhql9qEdSkiWl+5J+
fMgiS/woLlX4QAqU/J4ckrYRN/izAwbhFSzO6TPKsYbSahYJocIz/rh4jN3r
F94At3yKM4woawg+XTyzV25I3/I+yRBYhXlijYs3RtJBuoVFJ/5cQ6+e7CjH
nNGmvYaApKJBWJtllJIqQZJadz2O9VeZK7Ag1IeDsNgmN2MC4OFiShp1fJmT
s79/k6/Nip5dTRnCAY4I/fjlXgA9FOLgtBa914ZiCvLTkHB7xfvR3ATmeBEP
rKF8WDzS30BzQYe3RkkVaba5h+MzGy68dlfINpwsFQVXjt83F4//JOCwYli6
SAGoPhXVdaR+FOHf9UacA3+xwZjfvpu/toClmnFkudO81UJ9bp98CLPLr8je
gqmiEFu80niqJTqxYLUKO+cgy5hwZ2NvRTCyumXm8JMlKPf1N0oU5PVTlAkZ
lDrToXeWZWlWhhFdVJoGGDcW5iiAE85SVmx1xmfQVWjAWkbcYqnIvN/cwz0k
uP2LPSb0vwypBIDGGjkmupClDwLT36HZfy+eh8ZfSKdFOOfV02uMdMFImf7h
P7EcxH3784ReECSpeAIFgI35CNo2IHVsASzf3HE3FfBz8tp+TWiTDeYJpHMH
5DUUyLAnWBIpwOqcWxZHBPiu+H4o4iwui7kNYYwu+2C0ISrxubCoK3gGz+Oi
xDLqYpMlBCLWMjdaMl5ynduZahNq8JJ9KNmzh3UyePoZC+tGjWCw/3NGW117
fenIxbDgnPqwc+618vBk8EwIIakQeEAjh7Z+TeTPTmqnQqGVMw4cgJehDjeA
GtyN396shwDTUt8bvFKJJ6kefCZLnTxa0lP1V8HMelw/q8uNABlYyI8/6peD
MwqLp6fRYiLg/sMQ1nBUfpIEdB+GxfURavAbM5CJIdmXCetLhWNQL5JqYSr9
+XFe3aNoB+Bu81od83yby85bYn3FpvsPk7mwvD0GVlMJyUB6hNNcdx0+zN3T
zZHq+EIjn6/ouxNTFJoUoVwoB22hGvy1SJOXFybiXvH4iNyPxnP2VztYhzN/
heKm+WqwqIo/x+q3OLT7o3KIS0vhjN5lHCuql4trlMqSvokRMI+3jVV/X6Us
pJZhjAj5h/+kfr+uRhBRS5uECFG6EM9LGCjYoVlyNcCXR8R86tiEsUtGetQG
z6xc83BoEb94ArkAXb6kc1aNCsqG7/uBeAvHUNCO6ILH9glQ+9k/1GFl9yaD
W7cprCIy7S4hreNcoJKxdEO+faI/USXE1Mqwk6C0mCWNTQq50m46/BR6itQv
IVP09Z8qwzGzB3Id6pY4za5O5hjWUZNwj9/gg4bGyYtkUmALelz3P/8F5MAs
LLBK19qQTk/MP2Ad7zg6O93/A7GED12eu5umLcEsVuRGexxHiovH61+X6qV7
TAJGrNTGqkv6Hb3oJmMYBIJ9V4TzwLiRqrykpRrAWpUJs9oAXxL7ZKh0lTYS
boKurUKPgVWhJYUQUlZ6IdU3gISdBKBPq15ZVN4VreLRaR9fA/EtuDNPTvEs
MXau00YPW3QurPSDbq3pU+7QIIY9eeyWDKoPEl+n0/NGJ+2yEa1qUpwNdexL
Kp2Wosiw9si/t9SWI7cvVo2DGL4xFxZmZGkpB9GrCg75Dy6eXnacPDM00WnL
GfM6bwB0cCWkbjZVS0xr+2QcE4+mM65AYC4dA6XoU42b1C1aE5H6pGOFeyW1
MDJD/rHPkGf0lxLRT332KYXu8NclqlnDA2bUaScj0Ce97cB69vc4dT+i09vP
6+y0I53cJP2aMrxj6ZcR8ogT6KDx3kdyY4Iw3hmTKDO5Yzf9x0PqmFyuLvd0
zk5hNvIea81IJfTxdty2NFS7nSTHelUagegCsCGvMZDvcnoGKgY2afLoY298
g58rbrpa+tVeb7p33eHvenedUIHUlZqWNrTe3YqPdkV4E3gucErYWghtGd1K
hbfT4wpd0wqTSqXlfauyWx1dKhSmQoHipKalg/ZV90bVpvAS+hUenPEfsw3p
Evz5tQ+9zE543mir57+6dqIZiLTuP3vH+4DXvTqoD92o3E16q2BCfhFTUTUa
JW0M9+k8Ynsklw3RrzGSMof3o9TaZPjkKPTsnFB6320OeBaBJonuijXj41nc
aBC8BYZ/HSxtImlfaiJGOWlHzK5r6tiD32HoDKfU/mUWDfzDUWfT+a5b2Fq3
6QbD3sVYsnWfp7/6fQgSYWBlP7sP9sN4WczqYlCRp7ptwCfViu9pZVPFs7IA
5oWovBaFSAF2AweHo5YWt9GtIb0Yd/OXzVtclVgSLjeBcXcYOgclJBRuiDya
V0HV8XcAE9Ud5mQwc39c6ezllFG5Vrpj6AVlmi5my5CJaIVbzo0DltpjlSP2
2SAKeKyaBwtP+W5unheR2aczLPmn0loyuPk4aZ5K0JOp62SAapik36OfxawG
r+JOS/WpoMeGmBEOinuAoD+VzfaHTa2hTnU3ED4WL2b7IFsMLLicYh22lb7i
Y5BGiFtpwooy0hngkVzAXExKMkb1GoHxu6toHwguqCXFbVXZAkVCvLKXpa7g
asXI96KdiXcbZj/K2wea1uke08iCkW2CnwzxL+DUV+ciZY3WSIuvBqY1Hcoc
L0qL9mJiz+aBYR7vL7pBW88GwZYZv+PUq1thz0Kkus8lina81ptggzdmT+Kp
Wg3JrtRnDhhTTVi93IW//zdwn7vdOUjMIE80EgCXdp5M/JVvuLtZar8rO9Ba
KQjX+7CdYV4NFIkhGWc+DO4n8+VnCacLDf74d9gfy5+psv6bRv4/DOQfea0P
KAntCV0cgM4zDRscthtUR6U8dq8xBiJ9oSQviXnDbf0f4a4UTHdQCeLbqf62
fNq+1Athe8qjknJj+F3EPEQ/+wqCuB3E6FITHtSbZdGAPFxFaMV630Rv9Jgu
WdIrv+2kwEJ3i0jnfEz4uH6JlRyui+/f2TXySQdMHW61gmXWngVspIIzh4RS
4vVl5pv3GWJXs+lSfxWYDGBGTg61ZQDNwGdI8YG+spJ67zSQsjyFkNct8ILk
37uKBwC2kffns+XSyNQDnGlYy9t0QozTG4+a/z2Az2zi7Bvy4MYrlyD72EZx
EjRO70YZnx3aruYQ3FDK4x1ilKieOXJbPpeGaLdAkVKiNj0/t7eJRbXE2DZV
7KCd4qzlSM/f7AV0sSvI5ublQKY9t9OAzb3kcw3DrhLau1XG/jTAfnXnBykj
Je0OYIJgutKVyC+cUWugedrY0FWlbtEQlUJ9EUwqaqTs43nLH7I5PDrqgvuM
o/dH4RhkGmbuMYgv3wUfmjfL/kVf2uKl9SM+2ROS6J4SEHEuF4rKrIQY3Cgs
wfAu8/r5ukJZ4P1WnWUmHuwRThHi9bE6YZw1eCn6s4tB6BirinnXVEhoT6Mh
1JeeoS6ae6YgZTbE6oMnjQ4hpXUzedJNu/gM2ufPxqvH/c7HoUOeDOULSll5
YRGfVY9zx5mQ4kwmbDxBXCsdjDY5X9lL9br7jp3QgXA590cw7BL9vGTRZCST
kzuvRH/4tMipNDUCSgiqqZiiUM7FkYr954geFH+ud/PmCuT7zD+wiJKjDWSr
BbqbGSbNAQ2Poqfpdyj4oGRSnC0qw5qr7zgUjBW8klNTFKaiHg67imuuNSAX
KvP9Cblx0HghKf6xugrkCinr6omxXtnQzOcGtvk7Aewq74KZmmKFAJTurykU
+HeMxqF5a6EpE9MUe8wYYSJTl3OwNrPK8CkPP+UJH+k48QtBU122kChz7chf
1IF3fUkTiu8zY31zf7IMfBnumZYNTKZOGpbypSE+pFYsQNtTzBA4RUog3YHd
E+DqFnLWY4Mb080Q6hFWH3bvu2ASxFDWNRyumc4rs4kKPHRbfsyOfeRXE/SY
GycKAtXgjpaYXAjbROr8spMbU+Q1As2Cdjv+4TVqxBFjuACw6db1A8VztYEr
d1aP4ClYJ0sHwKWgLMmqhRzikIoCYMQBx8iY0FEIF8AR8PZuDMcjbWZaUbk9
Bh93SyulvrM3r6bKqQ/IlR/VAEPPjx0S/2hPEzX3oIYXsXTzDBxkoAeDBSOP
yXa7eq9lm7wWwlG65/7Znh7W7RrN8YoctWqjGGNe7qUZmmIUKvRUOJeuv+5f
blgDBLDMoFe0gTsyHB5MZvi5SIWyVaeI1+jG2n0416MP+j0UGi6K4wFooXv2
+O9W5Y9BsU0VLha3MW7DQU89JmHaDGOV8mPIzytCauTCVjr87ZOYF5b0svO3
nWhYvPPb1LVwZcXjvFfabUoBbtFFMNWm5oCYveTbm9oqMkInGS+AZ2CL8czx
txbf63JPw2uLptknLvQjFDKNp5jp+tlvt847qJto0Jn1JH7sIL1J6/ota6ct
ui8M8BQRfhBXPIKhbeND/ooXzQyB4b9dGeHD770oYfVOY0zRU5bwmTthT0Ui
+eJ/G0WJnqEbWVgsxJBoo99WTpoPJWaFs9uk9NIrit2K4nBCOTHkYdkQrK88
hqgQDawc7uRR/maU5g3L9pK++Eh+7HXzdWHdx1kEzlEIkGjtdTqFid47+UKq
YERngBZkESM/qSY1HlWx/6ZsW0mlQVSx+H9jSYfz2o7MNNHg+fT9G5YuLVU2
x0TYns46f9G1L26v7VsGcTotgSOWBrhh21Gr7mr0jdo1LGHH1w35hozr0JR8
doylm3vh3vtsnSLCgVoSmGoon+/f+q7FIZ0N8Y/21awLtDS5hmPiKCFL6DAu
GdFxgu53dw3/sXuouM5aqP679OtOwouZN3mzpVwhsW8KZ3Ec54YoTJA+XxLY
JpgONSak2iQEzRdtOOfymTagpLQqbxJLSWQZIJsgOwvAyzl/AeQ9Ode0hv9M
CEyEzndSVW+eZTk67LS0vOlzkuU/dp1uMMCvFHuA+MPmD0OVmXJcN9Lx41K+
m7lS/xNQBcEIddnXrgg5c8cIQuJVn4hkbx+ViMezTV+L8Iuv5cQKfTyTwfCz
nlIiaOBnBI6Mlynu7FjGsWgzyRjCN6kRHWVHOnk8BUiqSa0yyOtqwyR0aDK4
xf2J+dTLXymoQ8Mf707LtplAQy+8ssDaaYdwK33RWZguneUn1xDTZoVeuLyI
TD74lDmPam3hzYG3azT3w4jJp9e6/bvT1hX0yfB2ES9FPSg+ogkEEhwVhQ6l
qgq8UfwAXimfj/JztLR1kwm6tUGQO+jzjKspo6XstQX3CtFN9KXhUqQHtydS
iZBnRuLoplhOkyC6s7fqd7EXYsYsDDFPxc+aOU3FIdl/qyNk4mmOMYglkYlf
4QOSdhTJ8bMRpSuHmewHnbLDWytZScuV8kadKwVu9z0S9jrpNFJdHIJ0bNi7
42yTnJMWOu62V8fTOvbHE15zB/pXC1duZqgnX+6EDP1BRiOgNHZ45EVleH8s
tZ4IX0Pu4i9wwADlkyJ7x2M1XoxIbWeLxXtsq0TW1qAi0hLduRWU64vF5rhh
yhgqwvndx71j4yMMIhsrieNoB8jYG3+u57jCGVXA40SOtpZGpmWiVXNiXIcT
QDKw+HPPC9m66LC3K/mf9uj32Yv1ZKiD7z4bhtntssRCPbnwsqoaIMVz7k+r
kH6z+zmKojfR/rJ/m4SzsbnYga9Clq5UMsbD3d/NJJJIUP/kyQtxj/ZdTYvU
O3dRjI8yBs0v1odPMJjx/7Yn5kd2Jt26m0j0a7cr6a1Cx/0yeBTA3OdY71cg
Dlp8A6R5Yf9yBRypbPbOwuHJXFs6C5NMICLeTJ26K5RvA8MoYsrFD8bU/5SM
kE9nr0m0Ilw33GEY8oPZ+1rycGt29UopD01J978U9WCXGc88B88myMvpg3Qa
47PwKoiYAZLgxz/WPw9Bj5ZmzivlWUszkag4G0eKzNg57nG8W9GeDGRlHqWw
QuicrMovjG6/+snrtnyIjsMag72VkkQltHSlNtstlhvJI/9YL9lhOoZTFO83
zpGc2Refg2gb11KwKIkIvlqa3lEz92qKaduhAQts9PPvjLY5j6tsGU140RK4
UlwVp3e3C/Mwl9W5895thdyHIxYdtBweNeWv6lHTWsvb2TmiJhpar/J4MwMg
uxeJ13i9OB5/9ML7CIzbvp1T4kIrSWA+npBm7xh7MvXoyTSj7T3Wlz8XjcD1
ytD7TZL3HvSpeJrsWkQ9OdyiYErkIFibMr55E86UH5SuOdW5naoUIiRif9mD
VN6Yxb/Z+UFXBimC/bZgm04ATRIffdCZPJvxyvw7dtwa1r8LmoFBR3Vxtv0o
m4EtUXUvLvf23xz4SuCLc6qhCE2MeRV1AibjS54rCT8C3qbFUp6TgaGDJKd/
PiLF0uKh3xePASF8UjpMezY5cf+vyPR7qrLHE2Zjhh4xEn9o3Nry6vrrwTIr
9ruGHxei9RrSxYgcYakDS5dVWbTFDHwLrKmVcV/0SYO6+XT/cHLF61m9CDF0
XBv7abidjNKYwAku8yV966kEAmccX1oYRvplohHhEOKmNQOlnWs9Xl0GTCz9
/iGX/ohnRNiDTvMNdpZKGCsDERkFIZ/CQXTfMp+P5jW1QFvyj6r/GnVuubRU
xkP8yYLsSbrtdfnLS0bd0E33WwMjoZCom1H+O+Lpklt/7xC0RO4gdr+Ln8Lg
hYzV6xj8b/jCe3peeF34nhmKCzL8eYNGA/vhWRTqj85oJ51gDEuSAkKkGs5+
xGZ98d46dU3Q1ycOmmSpRVmJekDYfszh6blynG8nZ9dfuGUppuXkn8vLm+2h
flamLbcNHl2lIr9wc82Cod9Z8NxLeSqSLDRO4oyBCimap5evzYJYTfeAC1sF
W3OJu4zQgxwb5KS8sunaCR7zWuq5Ua2V1gdSEo92/qhz22wqIGtayYYY5hP+
Ct3LLtW0rvdzuo/MvhQ91qaAH6gyQlUnNLtGrFb7aojlRgpGajeB4tnz5tgN
q7A8EYd3viuvTUGJZJLW3x4U5vyuW+/6INP8JrHObLxQijrtn9HeX8AEdm2q
xgCl0BDL+qLloK0UTGHSoE5EmZdVB5eitWsnStm5WCecTIxHIwabU0MxIBHU
WhrRGwtQy2VieUEwGWc423yVDhT/8Q6NxIrgIv3/CeKGR+gnMVnCrrnULAAT
kfDnCU457CzK7M9UQpoPN86oKz4FizpjbK4AlTyGl0FRmbyyAVaGRtP8upGY
xW6qg32f0PwCM4TQ5XNTRfDBSJM9oYh51M0H9XfTbDKuP5eVKjUOuGCeJxX2
ZTlGX5t3B1eIsBNlX0HK2j3WpQXyJR6KA6eTbv3QcNQGNjlWaq/ld8x4EHVT
QPWR/LX/h7woVEukCLOqBhC/yPFX8Km4WYRGE3EE1hAR4VLafYzj9EUxmdGT
F6tWe3JDrbVeY7XBG2l+4CFdmxJUGUdqF0gNyYMKLx+b6rGpmmgJWPLtbzN4
RgFeD8LJjvKnsFbwBBa+fD5Nzp99BF45jARZRnZv/bE0eKuV1nbPOVRajvcM
Ig0l34X2hYmCvvtFmxvivTGEUlRlnOaxeOzRv2OqrkwwAoFZjIG0Ef3LDA23
CmRF1IvHswU6BmBLbwViP1RvCMriHztHpl/M1c9sbuqc1pJOoly0G1YelJPS
88uj/02UfdJqZmJr1vls33WbVreoaNmbXZSy9ktaHrpHyom6QzvMGt1kc69w
EPNZ7DLpIoPF6Zydg7T5c7xjeuD9YT8UbWs6tX6eQZFQKHNV8KV2ndNmlGWP
BUjmmrPpuhPk/YLSJFLn3vHXbaQSv+q0N+Airqrg3Jna6goezSDnDpopXNTa
w/zT85DfbFqJy6w944lx+3vcsBas5yyu2OEfKIDdu/n0Qjhr4grJ4y7pfon2
8RLCF1gv+Ru8dGnemC0DQ1n4nWr/bgRAQDHUCbeAOXpQEC6e780VAwHCF9FC
WQk0FqY8Q92FTMf2GonMAbflqSk98+Xi/nJKIORdbzLJ7M5g1I3C5jyoQIvM
zhZEmKoH6bow6MoRS3nt/ODhueO7ft6Dyr5kPDi9E/gfWz7ouk0KZfRpIh4e
DrUFSbKNCF44PDETj8D3ALUO/92bKb3tsbEHwb41sz7fRtyG6TjIMMykDfXv
EQIxI6jOYHdPP1XWmJxIQdEpGewyoPW0GH6KBXMAWvBtareBnleI1lj0GQIp
LeSf93qTIzp7GJAQHFRDyPPuzahRPufeAwieS+LbfHnJU1BGMDWZwE0qSqW2
TLoFggk8PRWTfj6U5WMRsoBDPplLpeM3q0mH50Gs3uJqSn+CaioZuOAcCZnp
JUGbKFZH9sMoCm8xFwF/Q8mM7sxIpr7PWoU5/7vYPdhZiA+kWlIb/xYJw8Um
7hrifiqzZBYBcHkOP0E00MGrAnHF1t/gMxXVzF3WUoTzlmy21cINVaX76ZVy
1XPsI+qZQwM31INFbje9pvcOZXbgqfD8qfQsi9KoznnaJ7tiSUm6YD+xYPHO
ozGmzHz696OO87Y5SziPyR6Wn9LwGZLrsokDaXhZ04ulitUIrphptwwBrA1x
yHqQkA3TYx4X+5qLIyKlDk7MyvW9Q1FJ0fr59mJt5DY+t9bVOrZNv372xRTA
KJKfIVukhDVc8JwWt224xIg8W4bPcDMVpuzFC7UFs/l4H//eCODswBx4d+SY
bjjQKAwuOHH77ZWEO2YRrOeUTBUgQTUpuBjbjIE106D3ZaBN3K2gZ5jAbs99
0djcHcDqBm1SOO3R2OOUw0vv0YBqBMScspdXENdGrZGBP7HaLxlT69xfe7KI
NxliVW+8CVD5WmHcorc9tWo6yEVODVle8eZJ87LbRacQtt3v6zT39khSnjVK
P1TaHEeo4yCvUjFq/2g5XBQmC4+UMwq3ZNnDL3TioTAOmngRiNMcL4P441jU
6SojK8VreKLf6nI0EOx0d+sasXmLLI+krYWiDo0CN42buHzOlkRgt0dWoWuu
wB8wIZCy+wAw38Y6e93yqu5rNeSg/xaJFs265EW6VA931LZNJo2t44dm3q0x
sJ+niL1I3pU0tyqJK92PEuiH1BVDfrjfkoZFPQybBKzXnlOWDhjPTyV3kyQh
rgIw7Mg/rvMU/5zgcPhluGvnfqG7zzG6o58RYyW8l+uSXaQCcB6ElRM+xOtJ
4M5ZFUMn2DtY8QQ1O8GIG7EJuKfqc0FcycqWaXNEyD3KZpAPvsIKrEbKgAsN
ni521AsZME+4Jvy6BEiKbgkfRQafeP8zgASu8hAmtzliZ1Fw/2SThEx0gULU
puJG4DgwMX7t6AGoEeex8pKNsPE+AoSmN9n1489ZAUvg3q5nvT4wvaQoYhYt
04q553VMBsl6+FO7x9DY91EX60MiIN7ndjvwVH2FCEbBNmxh32vYFpiQaXbN
pmyQ0uFirpA2Jciquuxwbq/fvvf8ryXdAHH9il2Ahh1vk8Y5fA6NqgHQSHNr
7ae2DQm6ufOlvqZO0nXuogxH7rVsIvCtt6+6JyYqK9UZTUT5jMqdRuWBu0sO
B8EHL2MfaiMzZyqqwrXxZa10bIrvBK1BKsxhClDdXoLW0ZN6Z6+hipxubLOu
pkm0Z1q6AHr8COed/9rriGOG6aD0/Jj2dTLgL5wy5gcFwnzGtvhsSSOu4ZnB
u8D3IgoweYGtbG+76PgYD1ZByXCg1cFpQ8aA+/CT0BI7Wn4jxWzWTV++D7Fv
AJ2RRHuVUsstKsUf03V7/Tv5X67ArPvT6Q8wTS2ayqCwal+T33mOkqOxEfnS
gB+TofAbgg2vfEe/ymCVfz3RF38w0nii7aofBWqwktWqi+GrZIpm3SPtCXgP
3oS9//WVBIK9hGN65OxSOeFJ5igb9j74HdqGUrVWy2HrD+cE+bfx8wl9OFKG
ON3lXr2NUYixO08BGRJj4E0pMTUSOeJGD5m/zYDCSxZwU7EDzqXObK2cEYcv
KrtwmdBuQXNswqi/agA2zYv2SmC2Wp6Wu59HhcwRwldGuYofw8Ldr+toYtUE
mCo0Eqc9h7HBasyQvFcQ5kEySTWt9z4zxrjnpLBZhgk7x0BoPOlYuc4ruthB
UXt5m6bO7LL6fz49r9AbYoMCs5KXHbWSowi1+8JtG3J6ivrZfXftRuDCJHpi
gXluAXnfZytzEQyRFaanJ5co9Pq571GAwEf5aJwKN+DnHrvLERfcJrNIbE5B
DRmRrhZk+i/1Rc39Q5Gt22ujWZTs0QYfXwQjZuUtdtbiQw9xA4YyBdV2d7Pa
Wz+ZBlP+9sb3N8Nv498ESN85mX2EZoxS5pwrJcA5Vz/uyXUPgstpfA957HXC
LnHnmHT7ztcV2CgnZ9sz6Gzy/aW6WQTENkJBSxyZ4DY2NE/b8AqUe9hATFWN
Av/S0SO6S9JnxE/KvyJnYptWU4OfkYgaz99xtNquiiVYlSCBF6ebisvPGEUu
4plXZELATek1BDeIL7d71oRig/GHLfudfdhpSnhPM1kTd9G7M4B+X4Dz/5HG
5vBR9AcJ8aHxy6MK3A6tz21zuZnBUe5vAiBHI8yCO3MnXc4TPlybPpEeUCzs
WhTq0joP4vB2AR1Oy5mnoJBhPmaimbCGWcxQh3Z+n4iE+KGO/Klri/4bG7eK
xu/HMm/0sp4uV4onlD7XRpwKY98w0hbHeIYCLmNDS0KH6kMIGxUpw/Jh3nkt
IhuHbq80oSbAcy+LXLzNaJsnBO5Ge975tMxqE4o7UUWSX9r9VBnsZmP1zd0h
cHyzjXN6T2oZOyUsXxgIbOk6ShmOWNif90/9SywHriKjEh/bTv4bc5HtNV5P
VRjSygbyYCo1ZWlXx9XZGjx9oaTjOP7dmQ4v720nGkbo3MnUDRGPFoGm5Zdc
6WkPPuqzoGYV3QlYg9BEIyQ3RnBGTp6PKSl8mmclWjjBezkb2jsVeeNB+YjI
F9eYQhZJL9OpYNE9P8FBNSPir488/4P5yJda3Hduuh/p2tY70EG8WJAaGyxp
utjkK9zIKuznbJWEWT4KYhtspuSHfg/i/FFQgSR2LRe5r2bslulPlPqa8/lI
avdqr9UrPwdIYuuwJzCMz1RIqkaPbTTPM7bcWAlXstxu+COy4B18BmIo6rwC
Vknit77DAofKWiBhbQIrwLRG0BtUsPnndFbShgq3I7hduA+GxAbP1eUPm1vh
2x0VvZ2Qg/+0aeS1Mrs1emEO5OIIXonDOTdaTWO5aD27kfJB7HYCdeCCbo/9
hvn/uii0cBHiSGKkZ8Fh7kxARoNDK8HdQptuRKksUsYj4pq6IaLAjkpM4QdK
ePNKK0xTTh1N3g4/Ju6Km8JtKkv0XGXZHJMouhIlNhMiJJTjdYUZ+dNb8ynK
aZo+Z0zPz37vqY+pptyglJ0JdQbk5EsXrmarB0N5mWfC+fn4/dL1T3B/7cm3
2dt6w6UkBZG3QdvStGrBkomGN5QYYXYoG+T+EFdJigpB+HvKU9c8CsysigFc
TINwDFXm9Xb76wR0BHyg55BC//rrROf+SSyMfxcM/BeZHzpX8LNBX4nf/AI5
WhPQ6S17q8Y0PP+Sf5Fr0fsikkUufshJHR7xCWnr326a4j/Oq6ykPeyZccFn
KUOh3AmkC0Pa/zA3m4PJU6EPLrhkga8hdJjmTW6lQ4igP/GgHulSYS5CCagJ
F/q7gTp8XzYT60wFBqOJtGU4vsgkjpdc9yesEvwEcFMHJSXVTFjgXGrvOigL
AhJpPPvLocxreDopDX86iKwXlou6zm33HvF3+0UlzOabxo6zchXzr4EGcIRe
0ng75Dhfevqo43N05MCXQ2dLVP5uyPuUfWspGzJmyAyI1Gx7LnZS0IG3V0Za
B02d/CJ6IZfHWrZrakRiG2R1+WFehT5vwEEMW3gCG2jhljIBH0sd1UKTC1oN
jpGgVbkoMghHBejBMDKXexn8uXRhDt+3BF7SLK2zFtP/nZH4OQEN5nxuXybh
XpbpkdHw3Dexv0w+L1tDDVud8al32yeG2jrd/iyvnNxQvZT0iLLcpoidrx4y
3z8YIYkvAkm3TiVszGohlLdcbMd3bzCA8JkhnRM3Acm7bLiB7Zr9fIMtW28Y
l4axFmq8WTZ3bn3B5xFc5bdz85XVPkaso0l52KvVzhVDl7zFLXqC89PHztCW
QaR1dErW1lWECVOiMhqndJLUkLSess/MhaGq5YI9L5zFpM7CxZscnPk3TOaK
1TPtlTCniAkx81JQ9Fp1wZK0TutbTJ7t8R0pEXDhSjX9O5wDjTZ5aXuO8KZw
dkOLw0l2WY7Zc6CDbzpZRZiFZJqOpeHLD57y25vD9le24vbxIq4lB33BM31t
8ruRQAXLYm5Wqx9wczaTTE/oyNL6gsu+xUPuqMY98mhz7UNYHEUSqKHcwBst
oSSN3n0lQoRHg4AL5RS6PJx/m7BTMgo2rxzpVf0y77x0fsG1Q2e31YXnp9XT
hrxyLv5Bx/A22YuoGjcPdb1sBjn+2IIofvm0Yk/yGaf8tMKPRZKBx6NhMKcu
Dicw2u9M+BQUpmd22u1Q/n7GJdbxy31ax1x3PeSxqjfi0rfRIrXBhraQUbHv
21RaaymfJIXfBpWRNxaXBuzJaD+xPQeuY5pvO11fypI+tM1ogArCi07MsqE1
vw7il/tmvPwWz7HguFutfWvFJR9ftstIIh3TyazBrKoYJC56GwG8TJufyX5o
d8Hk6XGrafvqDO3aNFjUrQmP/61KVl2wOvznZgMGLR21CLIgTAnIG5sn4DzI
FXfkIxaTcZPUv0pmuLXS9y2kYLViUaT7KvtzOKHxBE0krgn8H77IachkuAht
uWNSJ5ZiRgz6IefBJMD30PC+tU9G84aIpG/O4/Hlt49mHNZmLSOQChqnY3Px
0a/0YiAcZwNF/x/cr2J5kXxWIvsnbFy0Ke8ZxBxY2CXde4wGC+LczvC3gMr6
PC3OAoM0pbzypmkFUfbkIMPjfd0ZSnD9eZYFhO8N/OgJS17wnseilsVxOWs1
FurwQMQBXwueSb6Oxa7z4o2KEGtu8GcEdkr85xcUUf0iQUo1pAeP2jov7EKL
CwgyTH5ufsYNw985Toi29ndrd89I6XvPuq85eSTpvw3y14QVPpNuCfW72dhA
oWCFWiNvKgNev+YpwOCksc2BdnDXT3X2qy74Reyi+4HeI4/OzLw0jJR/ni6F
+f79Pz6bEwFOOASmjQYx/84i3KsJWaUwoyZCXCD6zIA56VvVlrl6HknE4HEQ
BqHjn4/18OvlG4bdSiXuMMuyeaVgeSKL0Jt7dJebDppiKjuCecE2aYiSXnKt
cIgFY8yKzsaG5q6MWQnv18HT4i5uaH8ce8ts+2xFUuxMdsfD7C0T8eIrFycx
0mOk8CIvSyIY0zdjUBKnGBlsQP/8c3DJAzhDwQbHr4+aDJbpRuKw89Z26xTz
aRzwd7tRoRgl2qWpcfd/bk1MRUCrAnOjsH8NGpFJWom56uoFdl2tVDeelrJx
4v247LiFADXMGrON9g/VXb083uKw1iZYl0Z23lhRXASMaX8VjgvoCmTXJG0T
TzdU5jIhZFCWqi1dy5ncAQRunVQGH93BG+L8AqbfLIzt+3IYmMs5gYZWL84D
rtEhHFN2s2DzWExaCAVnq+rOO+tW2ypiOWQfybjPSPmQpqkSj1AeTl+iPbjA
+8UJpQ1kAU6SDAvy+SaKLFgyyTaXdhJjv7TMHW5VX21JZ5OZsFkWdQQ5VxBw
hsmMvh+HTGJgJaNKreNLKD1+WwXteZAWqStUTzdKdVd6kQcPzrSs44dSt5IN
NQAOgooVFIGCqiJ6erqhnLyR6D7pohHwe5GPYlcuZkmw4VDa7L5nfA3IvpSc
iZvp5alaU10JgiotpByGG2e4kFrka7Mo686kbeIMI1R+r3xfRcMGyZUsfy1G
ibLdDq2NwAX/9O1/bFwZhunrCqsVQs/Lujf478/tn7N1NNznhC+FpEeFhlct
JwADbd+1o+Nfiu7hTznlgHpKMUbLlKkMjAo2gfQfdaQ97t4WdDlpefACBc2y
N2oUtDh+/9H1ioo4uDqu8izDreO13TPEHRyQEKdnh8jf3+VIoLsvKvMVsnZa
XMdtQWcz0BLkjTaw/iM0CkSKbsC85Z9d622TRXmW0fJSNISk744VWzv9oHDJ
BCNoVwKH2P7r75KVrBSds3B545MOngm7ihjdistNh634i7a60rfgoTv++ra3
+G0oZrZ7TY8Y0FAza0TK4femHMNfNVEAzP/hNa+orMt2f7hcHG1QjROmDABV
Hkic2KIoqWHG2cy5nY/DBabkckNZuPaJ6t7lCvQNMmHa0IdEq8wdFBXiYuFF
3ut7MU7QZWSA48QAMwf/ngud4F1q0Mq7HFho1GpfbJ75ZRtBVna7OVZUivco
rchXckvv0YfJnNdzn5ocpkjZ3YQfOyzDgiq/CaqKFcpsXJIhNpwwwPKazjl0
4Z/GiDL1YLSQpfxJJJCxjzSSW5LWiGtO/hAUG/maavZvrd9zyMgrrNAGpVK3
Ak/9mL7MdWgnytCfhD8xJVnLQ0eH+i43B5HLHRuM1vAGFehfAguy+9FMjaCj
uH5orBLSgC/XUXmJ0X8jeN30LSYzNfYPqnYJ9qr8jfC9ku02+uRVmuLv1bWf
PSJPB+MgOY/vI42BFCphMsiS+jEiXKzox86+svFpnXY3lHengnkNVylLPCMd
z4TSCzsecXoe/G2KVZCo7BQqbvPmmM6skLUE0AC/ctJVNWgt6U0pk79PJyDP
xAaKWpmbmFaYE3XKzmGtJEF1uZJRxyeQGdGH+CTVpduUl7m34FYsQwITtm9p
7chSRBXxuCbzR3/zwE0f7wyWso/PjyMsqaFZFUaXfyJOlRjJQXCvJjrS6G1o
kcOVZRABeDIiw6NAk1csp61ufDWFK5YRE22HLm5BM/pKoE+q2jnmgZpAR6v+
DMSC4CFIFk3W4LATTgxPXqjvBqkwZskUuBoxjpfGSyAiQX/AGmfSQVMpEj7I
dwvrIesbJAJ04GswASq9uePC22QHLf4M8FwC9F0xtgONh4TstuxZoFNepB/d
po/k2vTamYNmSeQ/JnGaMp2EP0+3hUVQbdSxofpqU4VzU+WoIRm8VoenpLI6
lxcAXAFBnULr78//cU9GKjxyo8zeFdxCvTFy2c/wGcGhhesdw1jEKfMkzYWl
veseDY5hpf7/TcdQOF6ZNlr48Jz2r+uJu/yqF5fWypFmtBfbUL43DVWlP4GP
hIHWKpUDeoKciWjuohbyynOYIjOp/xkVRb3F3e7YsZyCYmyItnQ4SicBociS
flmKEU+SH8XfVYj0LdJh8bUkxK/VEiNJCirlkhdUHJ4cSRt2ca2CKD30xT3I
gUWtbH/hTFw9IUbRyHACjB/kNvY+fTNdfv/AZhHeMuiqGVRhZE47aLq9xhvv
Z0AGPf9eVjcIB9Jlj5laOqxWcAxj5ea0KLhDyCeNeN0MdZ/jJL5TFwF9B4W3
DzRjGyWScPUUNP9S2DiCEAdK9qkzY+dn+RY300jQK7t4D9tYEzmqoYlxaF+T
ceJmCoqaXZTpYITALmSw3nnZS19efP1fLJVBaRHtM9GldTyV6UTvTk7GzCOf
SqOgdT9B2Insrf1liW4RmOwNWozAWVU3buEb8OKjJeAWrmrVLY+XGw7+C55g
5Vb65hsmju0hOXscZAIFZ2snLHz0J9kvtd1ctkjq+SNFJ3fOU5nQ+zGc0hpW
hzQGVwHlQYkxoeuuFchDggFzX2NEqVEn3YZpuQu7ifsf0MEBalQy6ZMxFZKB
VIqXG+VAwk/uAJB+lLOlyxBLuSQpPmX+bkgTXThvWwj09d+K5py8tJC6iaNu
qzxOUQbbuvT08F+72+QdyM6qCxTbLNMHKMTs8OVgCp7coClyS5w9P0nlRSmW
IKVsIiuw3RV9ory5q/aseUWURGL2CwQyOmGaz2+j94QZEY7kSc+5578uQlvp
RWOxTrVPwTuXrM5LQX2tcy3F5zUZ0cE0mgZ4ft3nAVT+Has5LYdkze5ms9cr
q0cI02jaschnnFV/MEr9BxK2a3QmjaWnXwUMMDYXZPpZEos8g9oPgZXNciDt
OJqqVMs0NuEgvTR0vMI4JJNFB6oEMcbQTetdnqF8sH4YweJvYw4IFU+Xt7U2
cPo73SSDgo1ki3An/S/kbu/futvhLzPcfhygKTniKA/WthmRCJ/83P40Atfz
h89VRKmXLLqphlNcd1WISWxO8+vLdo8/kDNwHIgDpco0SoMpkYN0kR8CqTQT
NXfebYaPLyWi5c5cO59GYxYaPpciOnETM7UPNEuYHPJNHbQdBvY/qcE4EkFS
kTZ5qk1aTmej+lJjGyROrmk2cMu7ZzwFI2fdrmt9mJzHAggKLJQPZ0ChxnzG
Ju7Hse1/lij87g3ehDciHKHAU30rDNnN93JT+ptD2+X0FbURU3ViIN+in661
tTGXXd6/n7EaGjWuyidu789ScCDPelbOu6uwjgNxuiBrazzOuYk33kdafWdu
BFZ7+WbEZYhpn60HM252UOwv43rNOQRSRrLIrv8yUJMLm3VwV/8b3P1c9z9y
xt/bh6SDu7rXWHyZwXdjv8co3GGFuNKffcC3Ce/6mSIiP5tuPFg+A3Rs96BK
vmzse0eyla1PG/xBAo2tkxs9zkXtKgCvxyXTpnVpJXCpPgiIdURp3HN0M60j
g6ScnTikE2Ga8i0dy4Vd0ZMlEE/3qRFjFvBHzI35in1iEGx3nXkFzd044CD0
hPSWVrCQP6n8EfFsyqH6ECSj4iLg64cFqt6YkCUJKwdzg6WuffzXCi4CrNzH
nXPdeOZSOxVxVoZUMeZ/M1sZUl7r9WMqLtElDrLq62RbtYZWcEOXbhMmMI1N
1mo4hujGwLGRtHvV+XZ91YBhNegV03gwLucR2FOZmgS++Q5a/m4JdDJnmHBg
hQscPcCuJXQH+RMRHhRGsAZ29g3zIvKDLDBlcJe4w8cndcxINB5RxhIjyugz
2aMw0Z7+5Ac0bd8+NwTRwS+xgXsWOqGf8xlQXRqUtOd4c1Dz2hnsXaa1wx//
1P4Yc2esr4cLjDEeQ9j5L56lQgVNDou0iDTn9Pa+qHLDyYxM1T15UWspnybE
/qlMsfOBvZSb6pxnlam4oi+AnydogLD01wMemYIWr9BfUm6/it6jT5UQvvJb
moDObock/AUYSvTc5AnLWm1qsvyh2r3J2tlsvCrzxgfqp+lNq8gVvLVi6nxP
6XZV6tWB62gcxZm+uHBAtezq3pFrmXps4VaFy/R+7614FBpcatOA8FfVdJ9O
vQKlKZWhsdLqc7tZjywrTzPSq8YiPJH79aqtu/p7cP22W9BVahsu5LI7TCWB
vH+BVHqDQS7XramUMqurpJ/218BL2sDdpuGe8vmopn56Y2RPiu8caTNPlGkV
pnM+nYTU2h4DIkhlRsqNwIb6FOEHezfijK+tf2351D7o274yfAw474eZHe04
NjyJjQKFZAN6gZAVTtldigVHn6E6hH99BVxU1A+6HWNuARh0WpJNTgAT43om
oGuiHwU+3HYWsLjhSP3NGqFaXlOjd1seNKMmmg6wynQHRBD90ZJTHIUiE5mE
5BfP+/nyABF7L9Osyd0ethZnheqDEpjqDwEcdbixRq6VRGB0ZH5BIiMBKXXb
uM3/2zH+C5LPkii13V2nSFFDkJxaZFX/HTBAopcTy/GjD+huiWntpsFpLkdP
5KCp1OYmRBvvtipmHWZ4q/ahY3QH8pnRdQHpAQPNzN+FRvpufs09d2sAJJjC
uO/h+5jjXZqa7PQxzv4U+XCHJxE3JHHnxVYhs8v2N9/0/BaAAm8ClydMyENS
YZqxEtqVvzy5tC81pNktoXcN2hHkO6UV+SYa8oIhic1O14SY7UxiCQVkpkvn
sldxdsf7CC0oawlnMlGtZA6A6InMzOg3nvICyfSlDi9hYcHrosfMJCactNOV
LbEDytmtEJ8dpU1Kb4zYbhtRv2HaJeh4vb14WijzkPFNckUJo5Yh0oqbTXrx
FmWEiQ6/7rmDAdeHYsQm8d7kvMxmYwvHCXa3q7kIrUCENxkHbphqDX1up7Ym
cHFEwgPaKyiZji/wb/65CkY0R5iGv7SS09Ufab6RhBSPVSPapz1IHFOv2Zv7
f4/InlI+b25vvTZ2o8PjnOWc4UUD29Y/DQWGpAXF+eQ2ZFM6fUt6OYmpRfpd
dTuU+bz2W0Hs+ESyP3ffZGosL/qtVgH1ChJT7GbuzgF1awu5qBZ5XNS2Sp7T
zyjsAeMlvA4kWDjp4petBCunFNz0YihUgY37Vb3iLlQXeCN/lzZ0pPpkqYZz
SGiQyOi6iFqYfsBzFuWn0i/DTZOx5VrfqCnVK6kgj/s10Ac4v5zdEdv/PWyx
Z6jXWzbTDKKB8AvDhCgYEZy2HcRUotFIxh4/Gn3F4sSK2rZgxme3cuWM31Iv
YOkgn05HwWi/3ndxt68GSRlonk1kOYzA9U7h+1psDPtMA+rMEK9Nyd3Q11Hx
3aqqFttKMP4i+IQ6GjSzolQyRKHG9PvzPp5pIQMJg5a0Rtc1vLjvGyK49QZL
3ySN41MTg5XWPmWFH0fEg6x7hjFpXeuvVKIbCxq1VohAzE1Qou+Yq3gB6RpS
imdWFy8/fygVKzWuTSQm0GCjSBD1nxLVrHtynwQYdLBBHWu+pCLEZh+KKRXf
2Sj5XnQA+BgJ+y8pIw+J6DArTF/aRK8FQs4JZF4/jsyHvDdV44EZW7lxOMc3
ou4CT77v0WHZ826usoe1hfrp4pUaC2qBfbD9QT4e0y6T6nwYk+BthIzBxEnl
y0v+GEEzqBVbxLzBMqHFjimGTNuQqmcyLbzwS2qw+gLtPOIciQtlhac6nwSF
UyDlyXHYv0QTI99cGtPN5AGspBwk0dfteFNiWnU1v2/orzEUIEcZLQUCEWcl
sKxm05vOaaKPgTVISu3lgI3V0thqdfoeqoARUyIqfy+zXYmajJ1GH+1Du32q
SzFtGxucujhZhZTERz6ujJn1YmXf/6sdkqnV557UOxG8HqfxPgIr8udTVQqB
fFRS0GBf5DdyqfON4JIDIkaq1Cc4WrNQ1K3kKQnX6TfIh2/GTQopID63/0Np
HZNBaNJNomrBWVFQ5mT2waqWRWwMHYiFCv6t5OgG9HjSRLqhcnj2h/7qz5/5
CxQPcAkWYMr7HKUI2e6+GF0hJFRjuzlZeHMyfpcKR1MG5ERbOWTRG2nbei04
NllASxsihvKIbGw/tgVikBQTjv1AlTZFvzpJqPi4ZKTEvNOEU2uRm5tt2rxp
xvUsyJqkgJJ4bvxgbHYBcywIl7su2aNZJtzHoVIvYi7kSGFGWyk3ohGcq5wl
gyCveOR9yPi3PH0Km8zp6hnSciF+Parjvrprfmk79ajEtnZRFox6AV4bOPUO
+hfZtkFQ8OtaPhXy1xd7/Lp38a5usnW3yo7Saf/PmRvGaOvMrzQ3PLmkVMon
uRy+bl1D1npKKFSW4Nc/gQhrTK06z9BQuBNi1yvkbxs2w+rxNxJDf4KOkZHi
nox6PeFKsazVGGOu318AztyFRVrS88nIsThArKoz+6QEk76wiQWIXsBj1r40
pyXEXBGuKJZRCu/bu5xfqJjSyGiYIw1M+hRzT3jx/jsjL7WomvW0BYYOE903
Ib7n/birjHzASeOa9IIgVN5ExU7lTEf5nuTRnQHM5GW3LhNiyf/BbkzOLpHM
aKVo/XtbZI2bKGxPh76i0qSLWrNYyUll6XD8fLeknvISsnVSQ0gLRXyqlD5b
w5iwuYFQnIxlXlMaTu7MxO2Zhj7EbU0qHc48918qYtkyhypba5KeUm4vkT7S
zVksHsucmBfxXTct1NG8aPwfljeDy6G6BtlDLwKa77cnQHR22o6io4k99WOs
rXmMRBCgXia31UdrjlBUqOH6g5jcrR1u9DIwWREMixrgIBXDVEaxq6axc70L
pJsx00UOxVvJY4rJIBSKo5wYIO+Lug31Xvs/qGjPQH8aB2RMww7C6B4X98vy
d4tOB1toNu4HqjVKyftgQa87ZThCjtctaCT34JkNl+UKxpkZ4NAFt/HkeOAo
sd+NtlVRvFZWL6M/FJy/viG9Fbs3La63dJHZ1D4WlqkCSxc0KRWwVgp6vdUF
GXIFHHZpCXOGx7xV1c7Xqn29cI+9a8Asp7flJ5DK9ETJcygGBU1Bm8cYEeb6
MwIRU5gLINsl+a5OCQpyWQMaLGLQzRgVGeWiqozW0DsPQHjfK1Qpes/Hfa/j
abkHpiwuA5pa/vCgd5x3ima1gJ5I9Mh6zcnTNnwU5XySO184vbDBGvQAE391
6V2u/PcISIiOE0E+gTXtJ6X1bEkz0/yqlo+G9qH1AwKOQxvAw2SGAfpVmNqV
iM23l/BOhsEUJZKUYCYQgIoTeew0TyEvkjCSLy03JnQYe4deMxiSqCl+mmAX
vKWFEs82fXe8EclPKjeImrDDIg+S+ODJDiywXa+tARsUQUjegUGtSS1JFqJa
GiUfybo/a3vkhMY0a/RlPUcXk4uLsGVvjQ7PY1Z7/3KuMkuhwyOTe3snBApm
CV/rfp/VSumYS2NPVncA6iBDLE/eS2vZ7xG6aG0+EM9WbxC3bmZ2tSwQO3YO
5bk7CwM/Wv9NlsiLwO3VcXCLie8j49xeAHYh+Rk8nuqdZQn/mVoEWOjhYij9
iwHm8p61whXtZHkGQ4j5Jf+luIznvru6ulgPjsfmiJZTsIuo8A4OoJwCm4+r
jhC2dYzrEdcpkaEJw/WRR72F9N/g3Zt/CY7JjPrLbM462pr1kSjiC3/iI73a
wXSEU9whvfFqewBYbeB4ZkZjPs1ULYWVEVTm9mWfIKg1haPEuMTmte/UVAXq
ivPaLgA9/bHtln24Dd7Yb4rid+KOQfjGw8Txy5ZjCRve3B8SC2WB70lRP3np
56fZEv9z2FY4A9CIgscV3inUXn6OCcDVXF2dxho5Hp4v2+cBlUgfnRncqmjX
aEfhMNxdNhpAwciaKOcFUcknw0wk3Hg5PkdtQ7bHQC2MrYPFSIMinNQkzkpE
y3eOZC1s/0drBQWWXmh5QgYvPNdx3waOtlWj/Y9EcbBW9KpZm58sPBIoFRj9
X9NwEJNwpbAI+ESLQJByUs8FU7guJQpxdmOuXdop/+rdqsaAezpze/TL+fzZ
h8xwv0iSGaM34pL7jSWpcJBdxaxe1hNVqeE8XHb2KY27z2T3W+QlUJS5EHKD
42Suzfdc2q2x1gILRFk8P9nRM/7ypjJHZ7RmoNfZIVTuJMoJGgGA4Bx9AUfL
nVtDPmKxesdljxOIew5tkG6F9ALEcKD5brxPfSGF6ShI0SiHyNLSn8p49AaH
ZZzB/pU4L0Xpye9u66rqqkwqzceoy69kNlqap+kV3LhQ8VH6p99WC3AT8rLK
zMc1BLj2rpWuGF9KVHC7VOlG9d7fJr0KeGGJvPLwlQvm1CNdRfTsdj968//S
6M6kp/92c3DK1YubFhXBK8aN8f/OI9neXPHriDX1R7mLHMBWrfhmhk0eoFef
K6qLjHdqn7krWCcGypU6f2lQiQNl2Ui7+Z3JRlri1Pjl5ZVgRMTV3DuqZv9L
0Q6n4HN5Z6ih5zIbFNhKNswnjKRofbU35y32pLTA++EHGG55Ci8wV2E9U5hs
H9OVurt8e8dLl9SedE6WdJmj8B00tSOE3Yf7IPrxj8lnI2BZj+pZBkHlWm8J
kPfAfie0+8HAHEpujjlA2t/1v+2KTO4oI9FCj6exjkQOixv/nJ4ByqXMrbr0
zd5jXC4ZVkjGBhfr6zVJ5TbxzXZsgVLBvK97LIkf9jFf/1wVpmBgH1RMkt1/
GxapsyeBlfvXHPRebijA/IoH3ZmDd3Zt7DKaVYKY3Of5EhbpUfzJbNQjEMBL
O33kg5Sh6TDfX1sVMeEb8QPs0Cfny1fMbIPTYfVTrdPkcN7YJEUHsrx5SkTc
M+lnj2w8P6uORjNnW+vT8dAEnDMMFf5E66IzujmzfKgUoLzoEKwMnlbMjdKP
0foyGC62hAgm0xknGsk+Cv1qIv8gUQJ52EaPLUfJ2m0SQJWoNUjxyMeBzYwM
CMMUmd6iaHEyR0wG57NWf1S7aSIVpY/Fbv7NST3lmNTIw4PMRsWiylEor7jU
fuYqel19g/DOQfIR889Tr9+7r13cqX9VZ+Xi9YTW/AFGaz6asHmKn/OuQ2FA
XnSvXn+SnsZMiqEYNH1GcPOw9E2kJ9SrVqGNpDx8vamqNGADUmf11ye/9yGH
ySDM0HmGc8c49BNBGBk+0Ko8uoXF7J1nb90xAQkYdJQ/QGW51IohaeaAwqqd
EylIlZNfSns6tu9KfD9/2HBq+saVfuOSV5b8uyfWA8NhvXUBPkrz+bzusSrQ
mtNsJEbQqdcKZXfO7RYFdqGLXlmHFfkADzrlfdW/KWv6lpP5PWa5k5p8rqjB
MY/6AxKq9AhsrB43ckAenpoBli+vgDNhhVLwM7rz7ipmTHxe5AJHRKwU71LZ
NT5cR4NWv+rOprAgrtIrH+14vY+8VNcs0us8AKnbhz0u3IYzU34LhhVuGo13
bVgFhgdUNnBst5E+Kkis7abdSmtwwtMFMNYUY5I+c/eFwOtwV0QQJ8WiDhnv
ujLnz2CoRiCJyve7QhHm61uwufKXwo9PlOgNph8/ra0RIGek3R9qexv6KQ8w
nOq0beveaI8sIw+HpLDpR2z38sFSncxHmeP3myVLkSlJFiba7/f1CX9AVqkV
sCS1qS0FiGKXiRSPcALEyCtrBzRj6GtI5RBhj0dqMiYpIMvNbR4OqMm5KivS
Xnp7i8RbT8yLMY5Vpg5laGSdAMpw95Isy1Q4W0MTm9q8L+xddZhcW5W2iz2F
A9nwAGIfVudfhqcm1yMLPYBQo75OkhUDBFxI6LR2ceZnEcgid93fypOhP0Au
rM7KWsIw+KO0gfZIsPbar3dO0q9Wf6v0KhPyFM430fnZUvZE0gg1r2i5vngK
8TiN/1GC1KBgUh+Zr3X8qoppwopqRL2Y6V/jyf9eLFHWQsuRW43G2qCSWntX
DDCH6WUWwaC5JPeI5ypO5Jw4Bw3xB5uQs+OhRA5uxdzjtg90tqnmI/DX5xoQ
zjR9dYN3NX/i7XYVlxJHbOy44Pu+vo8BAUR/NdRdUH5iiTfDZnt6pEC31ZIv
u1z5QrXY8lPLoD+ivAWcoI+V41UQ++KqYf2Hzwy+XMjGG49fq/gs9kTWi3eT
X5cvsk/p06l/PKXDXv1YJCzDbgg/oPq25lRCVCnsh4o0QiatDHcgDxAbA9zF
jFoG9ol6gT3qBtBgOI/bP0Vf6N1l3BZcUVs7jNIjzms2R2/Z7wVgBLQsuguI
G1348P/gpIaM4wBwoJQHRZj0zyDrHBgYh2a6vX4f6mlDl0J7WDLq29xtSwBZ
FyO5NTiH7VoYDuB3KQhk/efbAL1Y6z8VD6QlkFEgsemErvieVkyN76PtgTYf
LdHmTE3O652SL0JRVOGiCKMZfuggj7fdgzED3OsF4mhC2skmfvdufJsJuukO
RBWACH8JU+HD7tqmwuyFBkoIsS+Ev52q6GjJg15G5AErwtUyDHc1WHblYQfG
rRkQXylbpzOqcf4hohbIKlI+wx2s1pYducTRWr7+teTuN3N1bw3S9RJFPC8A
dkVX4M9BjM1hqLlmUzt6wg7W3+50fr2wZA1NZtyGgjJ1Ik/P6jVnlEBoZ2dh
9Iy7t3gjn3VaiXWGojP7/ng9hYh3lX4SVmlUafv1PHLkq0aTEywhCe5qZrAb
smSXd7NC7Rj7YtSYl1C1B9aLob3Jcbq32g3XL6AU80XsMGKnSZ2HCJfZgXRq
pZ452Bz0DEKcOfDVxnc8xWQs4cUvvDcQLvVdf507TZxUEL8hbzL/LelYCZzP
c2FgVyhTt7Ju9xHS17wWGyYqDsx2d0iiXtzcj/+jgLc3TWl7U7vexozfXsOc
mbPtgzgLKkm1cBfJK/NTfWCFErJIPPqEFMvDrTH4pJdwo6MJQKXm2aiKr2+Q
clQEjcRV0q22vCT86Cgai7r9Zg4gCv7LqmsJ3PzfUq8YhbhpNgvr51eFUZ3E
VPlRYA8leTcieaLHebZkCQ21ePKqFnYaXPTbQHovcH5Wsihc3QusjK4VvvTC
AxTV04fa7HBxAzAkCCWvpZnkNX9DTBJPQFNX8BZrJBkh/qALK+ky6gq1WKid
ZpZPA5CrxAwE0uWzfT4yeqT44RkNmKBZt2jprI+tq1U17lJDg6QQLy+RwBng
2Fjb08EEvxbHw3KnwPosBj1Aqy2LSQ8NMXdXKLeMnO8xpKn0b6xlAsyTi8oZ
6BSKAKggRp2pfPV33TOWfSP+UTiElMf2VnpRARCP8+WbVV7M4xUu6Zi6VdOE
HbVz5VZXKWHCtDlHSkkZ2SEf9G+nc44D+d4EHmJknsvgrDB5c2es0ZHCe/gy
5D3byWo57liH9WNwMcgTqRBss6eHu8/AmhMDnvHAqF2NpX9nIoS9sL61Q+pU
HsVckpRXu82VCaZL6HpTLhFDStP0Zx2MVUEaR0yGBUrCYaUo9aSWgXOlT/Zc
WCrkbWJiYDbDrnTmRIdhmzwCjnqzAxtP8D/JXzsNMTf2A6aqe/NN+0OKjuhC
o0LkSA4w7g/b474OO3rVFAys+/428uEztAgVy3TZV0nCNN3LzMaZdQ6X/UOJ
QD95ji25QYjkw+idUykPCPLEDMRtAUZB/RW7sTo5YykrOcvUIuNR4CoGDdMX
7JTbL4evTd2OHmi0Yaj5viLp5y57ZNU+Ta7s4y6rr03g2zhg0QyLcZXBXbx+
J1d71ESqKU/2SiBqqkYi5jSpKjxj38wtsUVeRcyH6T4PXHrv2KKmTw9ZfqG8
KLbLC4mqqWWR9byblX24YzVLmL2kJ9vkV2cgYqMIjjmmZFSw7q9aZVbG7UFm
vx51+FrVuhaGEXBzNyy//dYYHw/6OpmBaI/LlzqR+Zzj2NkYUn1lUSH/LrRM
XaQ5qTAPshm+PEww6o/B2JwPHhcO94r5wv62FrzUS3jwfvwjor/YhSE1SOE0
1LruAWKKMwLlPo9DiR5HF8i4wlJ/sJDzJqFJ5l76LjahNJ4daER7jtdKMHu4
9NOgBxlLyGNCKme6vjao9lT5zaRukRcwXGLuX3AOtInQwhwtr+ulhxqoWVmU
CfbsZsQ58JnDERZMquwvVntAgM36mnNunQYrR3OkTg0Zq43lvZa4ZSYNI+Ix
FIQM4G+Pv8bELhvlJ7vo8Z0AEBPSc4HKjWTF8hkK1zjPCcY2pjnOa5TOWRuJ
cI+PjK4aYxYeVXSHK40x/4/Ok2t8i+2FwmFUIsMLQcU9JdMxJGHXdId4u3Jx
4cdmKMon3wyNMSQB9wQtUzFAwFex0TjAs8X8S0leJ4pJpFZLHDgmBUlQGl40
sr6xev8F2FYbqRWqWVj7qxlU3sosMdUX05JSrr3uey363eVroiHuthp3ia/r
HEhmpZbZ1CZexqi3CZE7oRB/6oYL+jvVjWVc5b4ytvELHpXEAnggndGBGxYr
VOntMV2OCqNr9oKUKRCt+9fw3DK9pbCUtwMtQzbqo4wPbUbu8MGWJbTVObP4
rppNcp0r8C6zXDoMoFJakm67OP23f4T2z8AClEkTNaro5XpIKoS4JC/tDLmA
5UGNv+T3OYSAkvj6HCKdGWe74OYC5tP1yiPAOqktDe2xfPgRJxm/RlBIQFga
IohJo3pv3O+QI/dVl7cZj4JloI5lbX5sHsXdPJYC+H37+nza3AyaTQcOPd+c
nRhn4z9Q3en4NU6kAUrQH7yYmyU9sNZ00EZM9B/+5JnU58leuoJg+i4eBCcY
XrMYml5obpHelKuH1H6Nw8boNI+/6Kil5+6TSRxRIv6dVMOJdzGGb5nUjBa5
oacr2exV5dlBHzP3JaR/SkyeFWlc1WbzvBWrn9YKz3mA2Gd6+LtFpKL+5STc
8SIYItOoDRmFq/KfT3XnAJn6xU6mpf8pfxN5TbqNcEekRsOtm7K3JQofRSlA
rENbhhILyFdxBvNXuKqRoaI7y/yMyq5YQCd5c3QL4MUQvCTOlLJcQJxNzraY
Py/ygZflB615Stej7UW4FUyaXb+Ne+grMh9YKNNU5b+DdoBKtD0fCkK6Z0mh
O8fCr7DCr0pn5j2GJ206Lc43DufqLTtILslPfLPWIhsJEzRxwLXwqa/NEie3
qUOXMY0/DXlJx13NdwtwsG8dQeIrs/NMtmU8b6boL57Acp6gQmoMtrETIVn5
cuDxN52yJjZ/4jr1YIxZHMBKeZP3pPkOZb0W9JfsiEa9i3y9/GsuE9t37ALm
w5HChtuH5SA2bfKRMFaKRVXhwqupzb0GyG9UtTtv0DsiIGBw8DZGkKi7oTLH
DLzwv3Vq1mMG2U3L4tsdFzJbGgRrLbdo8hXV44lF+MHMrs9lGbh6zapRat9H
tsRD/BkcTYhJKEPRn1eFR+Ps6GVZtjSg8YqcrdNHa3b/kyHIG6RohjZAJzxP
o/RN+gJjM1FlfPQt1KUFGM0VAG6mTHt/MLOOui88INC2Y2HLj1lQeMTrNOYn
b2TzO6bI00OYGaiszBTWm1llM6vxDCGSp2ZXG43qpjZVXZMtNnoZ9ofW9JHz
Js4bXppXH1jEnaiG8cL9fK1/3PGnMghERFR05FaCUPifLKF8Nl1EOV7vG1XH
tCpJl5/JMJZm8id23ZalRz+VIyS4gqHbtnKLtrEjdhOmdIUpPMP2Bm1eAc9d
RDBb4TP86E26gqdRqtSxTiJksh9xBvuW5ovscKt4GBhxtcnnX5+DP9QlIxd5
6yDo12ZySqomIv86hVCbWE8xY20/0CVYfJ2jWO/XX7fmyh4orKuZfr4piYEz
x/hwbLr1ES7IGEzF7h0/IAl9ta7eJyuBrHg9VC59Wa/Wjair5pDAeyxU8Rjw
rCcEeqAesDvF8nIf66r4F8fz4nbRPABm1vWyLkHE8k/tlZPBYT0iBsn/CRiX
Td2LUKquKpFAVaIvOJQAOunq4TQd/HgyIV+lNOeY3bALJM8098HyjQFeai22
mF+OgckOJ9IPOqV/BApToAGg58jVMTEIejguDBm18YGfzMPuCJrTAwDEUhop
uHXcfUhzjll10xRnRDp7J8JrxkvAITfQnMOij//fyePGGU6OabcovU5oV3Ns
bBoWteSznH6Y420VOk6xCA4ebyR2sRnbKjHzeG1s5iCtlEu61+nb26oRrScg
buM44J1K0da14XQqp11ej5sgm1h8oTi+HcnK0k/sruP08OkhdOzJbT7ihuR2
sciQqeOKqQQEPOGT4wh7A+uuy17UWsX9HwsmXZZvsn0cCLffk8heOkB93e7u
eb39lEPfNWaEfNrxUnBuuJusPVKLYx/FXV9GAM46PPJsi2G9SgB+WQapityb
4zmqfU4ykNI7Wuq1dOFYCbxNsEN+bCQHBGYCi25jaiYq1Rxdq/230dhyWQc0
QsM9qmJDEx/hRfl4kKdO6DFYUJSc+3lLdjQ4YUYrpgrVJMnZgDppTOlmYwGC
77G0OudUZ/Px3OLtnKmP5QlM7n/AIbbdgyl9bz91z/ug5dtkB0hC/qTEi2Y5
kvGt8umahqr24MrJaoHbYeN4wiOGbV7eK4l6ZGzIv+pxef6MBQDRVNw9KuSh
RRbCZlpb9EpAvE1d1ob+6BIFAuF6vZ5Mdln95++FflRkByUQvaCGBYccA9eW
0WJLaEUKNERaKnOVjb4+TOVGoTwKemT8uixEnORwhRcJoWX3f1sAPCFF70Vf
n0KeVkY4EkUM5932EhJOCiBhUUO2Zy34I6BdwFvaL5jMt8T2hKW0VKz0LK7T
Eum4Pw1JsKHB6kZR9y0dRhWtRmKt5pAjHNPcX0kzA22EBlCsf7qeKPCGwwBl
XEUXCjw8c2/wMEYiMUj+OGH7E/cM4uzWGKDsMzUb+AYph1WrHMNbfDl4Icih
TfVV/NUhbwdz+9izsjWi2I5iif6IlFdHBx78qxBHhVPZ2T7Rr4Wt9XLOB/Jn
W4zoXE+mZh8tGEeI0MxJujdGK15Dz1R7FjUdMIh9CwgmKV3ffhqSKablR0W3
KMVFm9t/HddlWb6vXLnB9eSOWrZ5Fg73ClkYodRrO/j9SfOiJyyHwzDDEeP+
2kTO6bbJ0oMTa812NTULIT6VledVElKR/am+8f+f38DG0qA+ev2aVw/H1c5N
X5r9hirYzQKLT1aUY7bGG0yf98Ryo6vuYJnlIpDS5s9L5WhxNVOJ89dUGH0h
ZjqkV506Rmj6HGt367MGqLU1lSB1VMyhCWw5kIPRdF444cI33jxot1qLclo0
693bNA+9BE65R9sC59dINiqF0L3lypega6VUV3IKXJjbtwt33Nje0f+aekyv
aMgqnOFZWxiODWs+ZzShcEHO3PgKnPk3xVQupRmh5Jg/ATJm+HSnF3NR/VWs
ZrWieCIao+R0HqfMO0B8MPTJaMNYo8kOGfzYxK+y+0uXLCIDdCoV/UOKPxk3
KbV24AFgH2Y7R8vAlSDzmK6+95Oow/MpZzmD+Sgj93zHZ5M5ev5NUzVs6pn1
dbLf4O5qKSrJK8maL/2bR70q6s5Lkwoq9ecf5ewOILk5MfCNs+vF27NRjqr9
xMRtGMvHOAFA5i6tvkt5vSfIQqeO4DgsVSN1JMuR37njHTtrL331s2bOGkLf
Z8PYdtdsxOWBWVo3jCGdMjOU06d1aQxhhDoL6/pcBQDy7z1gG+lYWpRevrbt
PcpU35SWhVXWJF7Jfx7mpJz714cSLGfhqmPw+jFcDyiWGpQvrn65ksgiH7PA
waKxmcqj/ZxKN5gw84CfQ6F/7eP8Py0uz0oVlu0mPh+ZXAZ+yPIDB0X1mdRF
D6j2KABQ0dE9rtOmJQbNhvfEmdCP5MGhysaff/IG0CSTebWarXc4rvLIaXAN
KcSwAjr61UiQ8lT5IY4luENRnCR5WHUjHdX7lB6C+5Pe6fQNtFls8kBcQSdv
AvJw0uXQBJ8RFzCQ+PGf3GX4vrx2qyBnqjKaZGE1KLQvlNeZv3fes44gJZHD
k83zcjJZJGiyZfKH2id47D38oVB91RFre9/0WvuxiOgri2mQz0N2vxWnTrg3
Icij+SUcldHpBLbafnjv/xCMZDH1uKzDgp1Y7HaVMA3bmibjItlKUqdr70SH
23tQdARRS7ocZK2r9LQRRXCVlSrdsxzhWlCK6eak4jQYNb27uGA/CiI9Erni
TFSn+ZdiNphi2aF4YwmZniR/Obh9y/0Rf0rUmM7HC3zQCfx3HsrU+i+89ToF
HHMkI83dOYE3sCbiUGeB4q3NSYikr7VtwJnGIIbQTbKB2vo6ESXJ/ehb708h
GqQAfgsEmwIJRzx3PG3Ih7xOln/+rrT3RpN0Tn0pXZ4KHi7m0v+cXrGgVb+e
lStB0VmTHzl7GgfZtWZbIPfYmFmZl52bvEiJ157u1wQ1FRsJTeIY3939hOCF
ZETpJcIYcK24j0gu//BJ9RMemZ/K/KZIma18nmx/tLo8An+JJjvynHSZYYch
wd2vKG8nJlK3QFdykfiPJdjp/mBhZ44sDZuc7rEx09+JIp+0zccVgRNteuz8
PEyTugqmipvIYK0bBX4XB5K2dUDv6cWAxUK20gHLFJgKsvYqlPWM5z6Foi5b
JahlfJLWHScw2adVTlH260bfyuZ/yDifcCVOQaRpPC9FDuPV8JIR/JTNYdmI
y/mYGJY4aoiIWxdHfA8L0oqZ5qi3W5yfetF3efakf7GB0af0Xx/bIEIR/Vkz
erJfoQSufw7H57UtRms+p3g1Igyp67mY+pj7Zf9vmT7dLPHFCy2W7fIF5tA5
Z/DWX+SpLXix2MSvwf9ibGYW4vSz1NKnLmsjDXDT884R6+1znf406rh9USuT
90dvsIsgQ7j64CIPpGe2ZpwHqvPP+kTvPQpoDGwM9MXMsacu+wIbPDhUkRMI
9oXZkmwn+/e8admJSjtzN816MSxQf1GiDPpWIcW+tmOZAH67Jccmuv6KxIP9
qcutkvq9QB3a9wDW43drfqVFeeJYVjZ0T7AfbhEzmpMeEdI2cyrLFMst/CCI
FsH/7MP/JwbolXzxk8jiIiIXhGoUijOMDrG3be8ASXDXSBroWJb36gpRBTUd
lupbafIfdtln0sKLrnrUN+1F1a3QvJ3uWJQBGdWrHrLJL28BoxCkAwDQpCbJ
BzTDaiT5V10+pIA+O33JWk/XUdIWTv+j5YWWyRVQfGMyaElHIeSPi8I26IL/
GNOGZYXbYiWVwKbwZfj4B/H6EhMaLJ1TFdlJ4ThhZkbyNf+tPDPJ+mwmh1FZ
4OiODIll59YZLyZP2dr/nNy3yG7DvXB8IM6xEfGiPWSFDedSROydGZxRkpLw
sVdLhNT1SZyUFoODrd3684ByxIiDKuyCYdRf5GWlGg1kSo66pXNn/hfJo4aR
HcHX4igZnfwcX5hx6KiPKu6TuRW9RfnL19u5LZFz1zuURiTC7VZG7fBgfRk3
kLR4H0IB/ZcBPHYIszcq+YNW2OSK3nN/LD0vzx4uboR7hdjXshoocQnW4s+S
TmrGUafBBGJoJl1ckacnwPvjMDngwT+7s0oacDsgrxO+3YABFPbGwgm9UF+u
vrF+gH//N8g7XXwCvbCnte3cNLuSLsCiW0Z+G0KvCRrpiIUlbMfUORMEZEiz
AdHjfctZhZ/j2XW/pVrM8IzdYy0QKqq7N8k9ZWx236wxOJLqTOkv6LSQ2eSs
2+Cf+hZeySBVMutsR/cOes5Mnw+XdxGd2p4a2EUUQRL0rQzXewuYB2xymRMX
2PVThwgyXpkd2Z2OB3abZK/h/i0djwnz/DGSMManVwdx0lJuRy7oxoGD3CAS
3y525DtqO+/T7uUcFkGEnknvNJ4ZxcO0zasC4vDb4C5nY7TUrj0F9bfi0d7F
QfVJ4fGXsdkqkt3hMOlm/a10Fw4xo2Q04kV+yaPe724kfjgfaygn7ANpSGar
SOM3GkXdzjRRQ5Uio23Eya7uWh0eaTTTtk8MIdsxQgkOBM6JAnKJ7W6PTnwL
dRZAjc2PtgwPyHhUezsb+9FTPQzyVgZpKG7dbXTdwPrf1I9C+grWGY5GNDTp
PuLkNIsOOh3TwHb2mF7hwlQqkbbGKrg8o0n/W6tsYs+WHlgzsuQK8hWD5I2x
BLKj/2PUhCcVFWsB5IJj/2uHx8HyleYOkDB6hSQiB/XjJiwCtqfWXDXPPUhT
ATNqDswqbYkaGbzfct5RKsSOq/Q/sY9GROBso/h8Fi1bVSbjXI1oTWYhBI9s
5IdazVGjeZtZCTCmO0aBde+a2UDBz+6s+a+/CUSQdhdKXH0d5QWETIdMi80z
VuMAdQ56FPj03wFoKj9B/TZtrPsBD85uUYwmgjaEi/T3vWTTmQgBIuYMOrQP
1Fl4dMLWAzY2SKpo96l49x8K8h6rrPF4TYwK2jOHuYMWzQkyyRUEm9qjvpg/
5MUIRmuRS9TbJDeyC6J3Y7/wRoxAwNfrgOl3grEsbPuchHby9Ra0bh8bIC3N
u58UKDTaN1NWLBCiYMGKLKRVoZPdjFOWDmwJCKu9s8TNAEdIL99ZFaYuI2X1
y7myYl6cEZXenhQLREIHjYt9Jus+icIbDGGBiX0g3jaZEVcGcXbMo8IAZ9Gh
QeGlSZ2pBZ/LzwSAHvsNNsxzlmIIABovTX/48naf9oJnqW78Q2o29G3TZOL0
nRvbi/T5mV/ogAezdms55mcNrurnZVzI//rpgM4NLa8huq2lF2a3wrZXoYZT
47NsPkS19g37VN04b2A+yNEztk1/9ELmiwl5TodE6xmnznfY+zJC5CLWmvwl
A4bsIdhJe4oXf6D7Zs5ZxGZ3uNMDG9XyT5kdlswjOjVf8FUBqtr0eiA1s/HT
H298b4w4eQYx5kzxD8CaEYSv3yX8IZIdcqjrkbzpXtVZP4ZVUUIFWvH5ARbS
K8RESYqSekXnxxzow4lsGvkoIQkcagvpKood0ScP/X+N06EzAM2QqHtoXjwr
Z3chn3KBA8VwHAAPknDkrqezN8K39ZwqwjEDCUrlRMMEbtLifE9Jn72Xe/on
3cPbMOk72IAt5rr/6JfHu9tIVFXAGw5iEN8Y65q4PyORohSboWVCHPqV5SS4
G3wOt33SVbG0Vtkk5r6r5Hu4WF2n8mkqhSXF/24N5eguGNWmV35s4eB9pFYO
xP877UErDCrCOfC/xNjK0/Lj/Nfru4xU2Vqiw/3d/AcbGvBHM1hGPh9Fs5XY
sBpoTha9CmV+1CO5UD9OLafvcg5NfkA3f0eYwvRCUwJUWIG/bYXCBbuFPQD7
lpGne4Hq3TzIWAVbZOKacd+8kaQHej2ggjuNCnwGRdIbE85Gk8wfmz9UrgF7
ezB/uVMuPz+F+mP2RwhzBDuHRz0Wf975n4CrUFd+GdLX5eDsqVFB9Xej5Jdz
pHYrkwDn+BtKB3hqfJhbMUyP0N6GV+6Y/T0aeAuwIV7RGb1jNh92ae43baom
GxZFKjxY/ezflI+XV0xyNpI/OtabinKm2my9+I8/lFF2JwVQ6fevGfNv4PHq
uCY7/OKkPyiJig3tvpxCfd66DnZSXv7ZNqEm9GT1sdDXZbTsoqSpeShsF0Xn
Ru/vOp7fKIWEq+ieHPVbp12ZcrCR/4fKs1bqLlnoYw1U6sXSvbPIYdgdlIwQ
7K/K++FGiEj/IhrdkX2KjPFiWVpPB1IO+UExXsmFnG2XNyJBkhKRdKSE7WLU
ACAWw331o6wMUAJyyMH8uYCKzEc3+RE63bgxhQN9v5BVk39Lg6n+TUqlke8c
ZaFCakjY6LXKRxpcCHq1Fx2WWOqHwL3yXqgfkN1FfvQML1KuHcV5rXEVBdTU
DA/ms62GuAYJ+3EnI+HdEuYN+KUeno3+x/R7MTe3Bs6rylp4qysV8JNJiVlB
R1+zuzrlMMU2tss+MFhf4q+bmM8XiHdHiKJ8QW2OJzASzfq/a5FFO7nI37Fe
X9uWpo9kRCfjyVoZtbfK2V5ge68Gt9FEnG8Idp6qvNNbUti096DePWXokgFM
lGpjltSio97p7nKHjBfZ3uGa/N7iotba5eEQs840hadQfMza/7cAOnshcX5x
OachdW+pcJH/wBSprKx7FFTTpXnY2T4DiqODMXJELMIZCVGkqbQwEmXduPH/
h9Bbvth5tLcYsVdJL4m2YbZKMtkcHwlzRJL701olCh5v/b1ZKUDY72FTYjHi
A8eQw1/Xki8eE4Gvmmox+dUUgKikv7gT9RrypmquE3KcUWKKL8+d6R76GPN7
FpMqfoH3kzvCBtizTAmNmASRdQvsqA9XNltJ7Eyn69u46EbM+7plDvBR0NHr
z4J11yiha/0bvxdv1yBnjqG9HDIn8HR+ULwCoZU61+DvvtmteLzIr862j631
eIJdMdV/wsaLP11/u8MciI3OB5jIHqT1M00ED82UCGEtLygZf196F/QCmD24
2VieSjzVkDsPcfZi8QwxEIiviB4J7LAkzNFDCGUNQuZprMUuBSihf81LASEX
WwIujm3DuBAyCKkoP8REcjh2c48eMUPhD/DMs1DBA1h7ik6HtrUToK78NvfU
sm1rnm169sbX2i0otdkVhu1PqvKICzcrjRzpgm8O+V19TZe6Bn6mRQWKzOz6
SYo8yNc7q6yqHXgzWJw8VjygI4FWizDJRlr9fIS/yaGNuU6bOoKQKoQmj1Xg
mSGC9M32O00yZwf7CHWbg6HVoJrcaMEBumAIODLu4OBuvHwvzySVjQrmtLLs
YndgPjWMotygNqQ3d5p/DZC2GbnwbUkWgg2/XqIfPcCHUe2iFFf7quyWmjPI
qIQEJ3fGRhIDV9xlaS1yzY+EKGw2takl1l+pfjsQ1ScKWh/jl4RO28/mEqag
qUgraBcTkeCIaegGbTo+x6brXlx6rUaAtUP8V6IYzL/LbL9MbZQgYplNIOwC
bzprhstwgOvrcwYnBb9SIp4ki5J4szs/rAfqpFPAVic/AC3Bu2oh+XDrYw/f
8Mk5uOYxPL96SECcXeeo26QdAS+t82qqTVaq+FqsCudHnSyqbw7stZUTffAq
bNdV6UlCOqt+/IODNwVo1LlNHiHZWLhciwZCDBhTZGkOdJxAS24s+XIlq1so
VUqZY2vvTuqHt40S5X0cYQSlrDQQBGrKWaxfls7iX21c0pOKcBUGzcxD1kuR
5hzg1jqYztl5TpZdotjsfrB0W3ddzjjP1Uz6Jhh7vOdZhik7YT0fRP+8A6Gp
u3QWU43BDsSH5JTtF+zb8lb8ia4lHxrTM8MPeiAlVBiJjXjZdU5CJw01Kt94
ShPCjD7F5SvOJCSPq6TaVfJlpSSulFWqoEGl5WjknxL9YCLrF3T+LaiZ5810
F9CiZG7swQWnlsVh/L1g66FtI9XUnxve8IDjevenYsJleE092QPnlGb0AMwU
pSxtLH0cPpeF5uVleifm+WLPvkmU2tVlNRdWy+olrtA2EMw9omKlpM+INeo6
F9m92vO5v9oBw78VD5MyrJg1PD+z4FnyD3RhEcVeZW2xGq5jtfwoBY5Wc4m2
b1puMe9GWmngiJw7muDUFHutVZXSuUvRWcd/PMebQcVg63mkUP9kD9zrGxw1
WHQtW6PigJ21+ujk+vt+AyCetj7lYXgm270dvL5A0yyebUtCmOY95MXJ5nFY
yRsuK7a/LlT3xTi2alg9XLw9daOfulVwNHJlp9unwQ+kElD6haQVfNcPkRfq
sadRTd1SjeZnApTeE631QqOfoFIMF22j1Wdblfno4RQNMnt93W4qgUjTEdFC
gY2HRosASk9q9i6O/1J/HqN33hlLCQeHm/Kwpul23pnDXlLKOd3izj7uKpNN
6FTYdNN12uB2jKOk4waYzT/MmEpMUaMZRA/YByxANWECGy0ai6Uh2RpwbcjV
GzFpbsyMsTh1qp3BNWCflCubbxsbICVbMxnEmpP7d/INoShlRUcDzuE5oOD/
CGw3aHASDw1zNWKHRyYff/ZyK4grL4vf4Wgh2NWZzFT5pfNVcPSKJCIMhOar
cyMipUbZKIXxmdudAdeTtuCOtny0mQDlWdFfucdz+3rQdlN236/vOOgmAcEK
zvTtM2W8Ki5no/GYLukfFRk9FdBD9GvqrLoI9gDuxEEQU/Vd95OZSTQmIbKb
WoHUHifH2yoQuBHrhwvWakyA0lnOohc1NzKwTUaMu29H7x7O/Q68kHzL0p6K
M324A7NQKW47I9qiVrHXft/hQWejQjNVMsj2Afn7A0Esboq8PipeXlbjitDr
vGDwRUjJWrZlCplb/0cQjw/xVBZz0i7ZBrYAIsu5Fgi0ooM36xoF68FPt1kO
pW2hGrqu8uc3wbnUkHz7LrWvyO37lLK7oaRCOCz+0n5536gKl9TFK849vqKN
QS24vbKAF9QrKwUusE67lXmOc3BywShqNKZ+uZi9O3HlC6PjK7wjZaozCaU7
zsqzphTR5sIt8pFbdhTYKW/ybW/1qx/TK25gqQN6nGQCOxVeBOdWguRkhjrp
5PLbkMuT6JMpOznzG8EZfxERBL1m/vmX170uAyRxtcx2uKMbM+dgn6UOzdcN
3iYrf7jwtjitak76CzxXRMFI9oskoPO66+8XPA0iB6MYmP8Y/naxfLkAHjYp
zMPmWq17apHOvEkhqVbNXjvM9adHOVZiJDPpPJPC1SS2w5Duyp1Oww1HnDLq
T1BCNkjDBv+Lk09gO8nljfpKwEtgANgoqEhNvG2py52CLy9W4SCqXuKqGd8G
AHyLRQBhIX4p7D8erW2VkA17TyZ9ES9McV7uoQYZNekQnC0lIyYFKJ3zoTeZ
etsKUAwyePv58DqNzFIj4ZILLbZcjuqNuPVze+EB/1DaJYrAdyyuMTbAhwkf
vH2fVXUc4iXIcELhXZdBq7q7DlYX2uY3DHsIzrMZ1JPptthiskYf3FI2w8tm
tw4dzxyDQn6bUYFa/zPCFU8BPYgPya7e6/T2pDRTU9eRpbLSxE6DPHx2vCzv
mcjM6ABkLGRj0wth0kSrn6S/iHiZvm352RCAvSUg0jkeHJtlUhwTnsxGTmVb
WY5SdRFJedKaC6NSYvXCYvB0Aus0gZOlhxwPbCoNehxWAN2p61YEY3dtQ+jr
UbWgiAF9OCpHvRqcaUEUojAkvz7/H7Wr6exyIwvy7Dnh5ockouz3Zhfjvc6w
eN/CHTWTFjb1veyetcEtRD+Omly3Q2V0hoHQtgj2F85x3lIXq/TJwiH+VSaX
/G8VUuOWngEGCQdVElsqyluRTpCHc+Bcc36uNcNsNMao5wNDq9GillIjHAXR
wDnTDgn+KZICBZpJescenxMgwozoy21Hfot8JgWQwBAEJzyz8sICrsRqYmE6
/oj6O5okXxjwO474umoOoCDdHyF6kK/L4ofsJSSWGDVBObs79gMiaWOmQMDs
5SR6jCXS0/bwVyNOyhkZMnXCt4uSCrd1hn6PAjJzgX2a2P8a8237CRiDa9de
N+tNnEex5w38CDfZMoZDUMBRPDOMr21n4I79gX9FAK3gAoM99u5BFC6kLaXP
fw0d/Jw2Lb4GpiOsmyUYww8t0AZUit/BctZeV52hKljPM3vP4/39qFE3hJmS
HGCePPn8B3EqykUuKAsVWfMVP5E8Pc1nw8z7/15jab7hPD1uWB1SE/re8gNU
5KgolycaFMRWieapnxBk5Opbk28Oo68nNDn9JhoRUsuXyG2aA7258xHDr1pG
FG7k3qxku71mgd8sNfc4qCdy6XiYGrTtUw4kAknavM4MBADumBSvvTvzA4+K
PEMMsGsIZAlR9SZQjsudQEWIO6ayq6owZc5aihOI3/gANc+E2G/fusKFKSAU
bXNkzMW1VvXxSZLzgGDSHzuoLmc5C/j0FUPf8tNe6wDcX6W2jD72o+0+Hhcu
d8aw8vByRSFCEMkUisbkHz32h6U3m6EjPszkEfhZaOWFpXL+DtH6/fZ1kmbn
nceduWXD4bE5YRmwlIy1ulitfLEWcdbXRyorHMr5PVojDxp0qmNoQa8wUA99
zgY0SMDfVga0zFCmqrIoX4C0QQ+sS4IvqKXafKgCY4Aey3zwywXbsd4qFxzX
iwD3rX7m6oCrP8Q6cJXVRU1BIlu5s1bgpKx7a2vaIx08FCxf1MJgF8eS3ap5
DdhasZEe0+KoApe51aYp3M64sjjhKHaCqa87zUTHTi8ZlCK2SY2u+0s3+AyJ
iITq/GaMGGfTEFV7zgMM/l9cWROvBoav7KDKc3ehbhBbAZ4DvYnofCkHCOhp
UHw+EJoRFPQDZZuzV9tW3PYniWf3nXh7tlo+2SmhSeKoH8dMoP3bmz/JKFRp
HKkYPCfODSuxxFP5erisNEm6RKcdLsd7SrmOT9QV5ukCK86IQAFcVVpG8ctG
Fq0x0ThNGXGQ75+xlHukiEe1369no/EmWdMuOwaGlNjKXqibAUPJ5/aTCaIt
JxoHYlqdTKS5Wg7E4GxAKojEwin09lJpA7uuYru7W7Y3KhM2MSpFAjtxVYac
oM+BYhOS0PwGRlJvPFPBzOQLMvk90xhps/tvai6aMjHPHJtuzoz9YN2xz8cs
1YVtXl1WzfT9D8eNr2gd9ar/m9ZPtns5KEWZAreQ1KIJUufBw+LRgyL6saYc
I13EcRY02qApbE1N7+WXGeeOjmLA49mlEQ4GzUVWYUABpgJNSsPILGtVo9mY
1V4hSRXERPyianH/j33GxgyKW73h6t/Cg+wgRAaCFQSjOsYGt71aS8zojUKO
vTAgzbdM5z+X8TOumZwSJuiPcmeubdHgyZ37iCheqSvHYk02zeSBNrELQaiw
vA9SGlL+JgD0tXcLxE5z08cPJt/Mv5mKaNoW5c0Qx8PidHG07c4hlhm/6l5T
9qQBzOdx8nTBy+PXsRF8Tv3yosgW4ZtTHWFSD0F/rNVl2sUd9DtPf4wQk0Mo
v4OPUReabxqh+BDIOzTvVJe/yBoPDT2iVwOmJIBegkU2lYScq+q20Ml8rP+g
HwkXG8vrB5Tpi1Et46CKQIP+o6M45FC4XWwWWMBuBnmgcA34Dx1g+9/kHQ0X
LcmdmKAJac85m8Fq1IcYI2JJ2RZ/JohptNp8k+0AnuFczBcsAeAk1dI+UuaS
aOVdvtQYohHY28ixhiP+huqQNminW6HT1PbEJmzv0/Yw9nrOiXDmhjVYuu88
HVIzL4eNMRiFju0DtXkuHhsZvrVQ/R3UY6sYSmrS4viiEwOXUselLz6KApLW
23n31gzNn/Ss28uv1lfac0Nx7IAUj2kOOAuRXemU7/b0Lrvo9ql4Y/N/52D2
GEeos7PLRfJ5QILgk664s0qJAV5fOp1VUwq/PPkC0O+pfGWCBpv7rwHY7a45
ajjCETB//CQL8UjEMr3T3tbVIAZbPFPJkrVUyKwkvPlGSIy9Kdn+ukKNEmRo
RSvmqJjsZVFrJ1u8JeaE5juXQ5XQOYT5/AYczy7AX9TbV1wEOSwuwpnuTE9x
mAgyZKDFkravc47dpXxAJHoHitjr8GOlkLOd8wjFZoMQk15FQUWFXZKRdfMh
ze1rJrKTMje27OVWNxCDtkyHkFJbkcwETI3ZZrSRGHfvvDtYMAVgeoVdVJD4
D92qyA/hqqR6HDExtzAXa10Xxz+Zdp7xtlKikexRQ1XfsYZUVwaOXzZFIrdg
TYkxAOFaaW5SBkWjp6T2onOR+BYIAlUs8I3Abjp8ozEPyng8tCtMt875Hnzf
/Jz6dIK0gJNiw67yMhawULpxuLgXdePOl1UsYIiirZVyg6mwHY+kQMJ790qu
n7vrF2BrO66HV4AZLhT0hvZzZjRIw6IKtzQ+AKKxb3Yo6b7CylYv1IyXgzna
RNZ3KA+ZXLEuFWBFxtwhnOOGUAQnMUZQ6Q7BZ6+EMvpZ3/PSUNnpR+cIoE9Z
8xDvyYedtBBRV3eElRXdZXu9grglPsGWYvxhByxR/qmLYPFvEcRSqOt7/cgc
h4ylLA5vh9jOr3osXPLejKQWRoK46+0dOZn2EgCSq4MA7Rb3Fs54IgMJcjCz
8wPFeLDu/sI+Lfmych8nE8aXcyEoimhGGdrGHcebYmhLbjLU4UWz5FOGm0vN
Je3BWK4/+ZkVKZkEawaZjvuQuWC/ERNcZ++hyMboHH59N3MFfXr591tV/K5m
bjwHsxgm2hvsq9TBNydQerhXnQXPSl7Ptvs6OTuwgHrA5OM6a0pZDvKZ+c5Y
0MoeLB3qgR/3+g6M9lIoeYyBRPDieNgfd7RnTqUcqp2VE3NbCQei0B5EnKrJ
c+dP9iJr6AhEHZ14+c4RcVpo5tVgH/8fogMRouepOJSE0LO8nBLzWKFQdAvF
QRZMZ//2bmvyxGZkyunGXuDOlmae3e/Jv+sJp4gKQSqbUOXLMqGesKwe8UPG
OOo1KBfZa5HBjPUX5kknFCNryQBe4+LEZPH4YJoxTXTZmiKFDbCsFGJmlHy1
ksKTbpK4oI5GpLegeH2ZpWTjZMnDYTHTOhlO4DeNHFFg/1YKovkMZtjC7GJQ
pCy3DHE60/HM5t8I0Z5/lZpe5t1Hwg/2NJ+QG1WCC8G/EOS0iAynZKPmIDx2
QV8t6n6a+Ou0e7t4BmcYP/QfYaFf+KtOXIwssGgp6C0BKv6k+arnn0zOlsk3
T3IKDEsJSRpSiaquUR+fPl5Ii2mAx3f8TUlIUN3EGvTPMcKU56KCsIFaoNcV
hgbVWWCu2kX2Z1FgSpb2YBG9FbY+jpD429Sh6ptj68LgCQUAfKDqY7zX7CwK
Oq2a12ndfeR9X22JBXdn+UdUNaG1pUs+lgEzRiUBzzozWOLzLmAeUlYzDV5N
slkORyXgw4e97+TcCw/D7YIkhgJjgznwV6g621GmOd+6bopNJAxvEhZt+ljk
bz1tjcpRDWog3MB2cnCU142xr2B/6OYlgkLFnrWB09k/hYpUFHaVlnl5gJEo
BCKSvBKfeSF598IhDlU8B2x/f2VGkHXJzoo/T9wEMU+ZxL6vmf95LddIINXB
d6OAM9l6VzFSdcvjLagGyvYRqq/vPBPQ/euWukt21NgrynLUN8dMyp76Rs4f
FbgXWIoV5EoYOfZjDzdmD8m+sOaE9GdAse9ONo9U4DsZ+GmK97gN4XGYPhv2
6S35Gfw0sMX+e5yLvUj7Gi9FF/+jTtggRbhIrsZdgHhf7DGP2jAeXqru9oYH
zdzV0gxPhA1S3oEurDtjaVpKeLAmyU/0rScqC10FHUcdF+anT0Gca6iqNX/l
n1+MaE12lmfn+zd1HUrp8DjTigmULKGsLZCtqY5GpYUoMzfGWw4A4kQaxp9P
9+Hm/TXnXrC5v3VIhn6Kjz0jdGfZeingwFShYG7fiFsQBl6xgjZjuwgWKsdO
6rKs+OklLkx4qIfRvL/QU99vh2L6otVd9CBJvjmRyNL2L9wf9izhQ99e+8WF
/kSwSdd7SLRH/hk8mLO6r+scdfHrKseeGSnHUj7A5peUreGPvDvJKFyiI4jn
kM61d4eCZNdLQZsu+HUB91ers5K/T/Gwwy3ScqFiZ7M1tuaAdQ+LI26WHN2D
WBu5nCMB97Z3r+VE/Z8PeZMusJOxtgRGSGq8oNVlPpURTCYJy9aunvDh4Ed9
t8sTysTO+BnIHrkwrWpgYFk6zGxNqYMEkXP2Fr4RuE7NXVDPl0eFUL3Da9b3
wJp0ySc4+BZkIIpyQBAoCPI6DTt7oazYzNPdEIQDAb82WBJZ6VgoPOs5ZBfU
O/PMbRxd51CjEQ6kzmwE12bIMukvdQUdvu1BBvpAUWOlLNkqA+xEejPO0lYw
mVBoqsQnhIntleWhkFAwcsBWp0SkOiN73JvvA0sxR/1jZIJHs1Uvqgoi1cnK
gVCLo079Oe3pCtY0xcE0Z7dwKQN2CggfboylcoO6DzeZAK1ZhiigMfsxpAyU
NWavjHlmv5gSD1s5taBa9QRSCP+sxKz/0BHo2wXDfWAFWgw+WNQpk0TvK82R
03kWrfqrpfBPK2Br8Ak+cDUm7YB8zgIQucrosdgtbZGfuGqY/b3kAHL0FVLO
ef/kwO2C1UFW03o9707QKD0Vp5fpq1EjthW/tPFEU7psu/LcQgG9OqVFOnOP
adkD/pVzHbDVx3M47lnrCJx6iu20MpceslNW5N0olZupNI7aJXAkj8vbuXaX
XXwNUUcwRtI4cCJv3Mur+6j5K49LUdEXFfoJqd8QiSnNjNyacE7SCRNH81eV
ni9p+2kfAV8aIkOivZGyM1oZRDrDMLkcZczpn7bu33kxTSI6dFm4IUl3f5ey
s0FwYLYbzTKnh92UyRdMTQVphC5wo7mtT3VZpFcklbNxjhcsrk794hw667Vc
VQ9tWrsJCL4QHg9i6HG4+8P18GPjC2jhEM1fQmVECP1FhcwscfndL+SzgcBA
jk++k5b8fj/LcNift664Sz8EekFOAdJEPFVywk5j6KLvI4rhi/8OiI8kNw5A
rZR/vsKIY6Z4LLt/IWd00TlgmqsMcx+8MxkruemIIdRbW507XNK3lllQWblD
RhPffG2Ye4UvE5ul/ThgnAvH3p5CV7sDq4YP0Oa4UXuwT/xqwzoTGPsiHjDk
wTfyIgEInDxm3Wacm288b4j3+JVM+gR0XA8JEv/2COqqmhcEOZoYNSWvqXCp
249XHpCbbH/+nvTV5YipxG51oNFKhLlU+pM0aG/kVdoFoI4B9QsEbBg5jIIp
1NynqBLvYiYcCniAdsqUMxhJon75HEPzoHBoiIz133HCillQl7qidc81clWx
tw6b8HnRg/RGNGkHJzTJ9m9SHvpNBeJQhzDNGPMHFwfBgOkN68lCozPrS//+
6HzoSZ1rirMW3kP6BZWcBhgM79cm857O3GaQjoBSSgf1vgSsYVu/a2S89HlA
zG1RB467qXwXBHd0DUVVx4k+wMyvjkyqtvi3p8PLHrXwBa4sHHvIOVxBrIzy
t2WpUbeQWLgoLKj7HyvxsTmpoaVIISCzyj70m2g5KvKeLNzWg8FzpKUSAois
eKoDNkSip6V6xI8Z6trXMIChPuv7INhYhCcRatPPw6uLZkjAEen8PJ96OrB4
LBOi1Ha+/sYGVb6LJXAeSRfg8PMfgNTjE+1Vdz/vvLKxsmz+aVMM21Xrquaj
GJapm66ab7v8XwJOoYHS678rZsEu9LwMB+mSnZ+RvQDpoaM/ixNsyVV441L9
8uB0v3pIp1oZ9/3pPzMQYGAf6H3JbQd7WD4lVBRVemmv1DjoT/dPdB3LMiPF
oScHHDSb6uJ05S0Yu62LOUh7BD+z76QAuQcShGmSGEwiJ4J3jO1SjuLnl91P
IExy+xjc6o2uSqVTsQYWINFE4opn9XzG8aF7DRyHFKMJ57a42W5iz8Xc6Sa/
bssG60dkyeXsPp5YjYJqpXFggPT7EkOU9H/ZnlKQVC8RA+KgUCAmpnT0SWEs
ZWrmo8CJxaO4kZBxStzakwZqEWKpP/V5zII4ZrOgHAJ1Y7I1zcmUu3ZRvwt0
YkvOMIrz53qnnIoQ6tSFoPhLX5AfwplCkQTQDAJrp3zYMuSBO6LI6l1Gq6q1
dk3f41vr5Lw15QHdPKkft+mYf+h7gs4VBhcHPcLzHmiYIIMlImHu3WMqlSyT
qKq+NF/nE9VLQ87iykcS7tsBF009Cw+C5f9hPb14Tutact6C9xpQe0FcuIAL
V35/wtIpjZOFBIl7tLVuNAG38YRfw9s3/AUHrtFAkHQy8cX0K509ppk6rrDo
VQfgLrNnWXvQw+U7kovk1d1N+hGpGTB1smU6uVRNaKjCgiHY/eoJxt87fq+4
8SUi5GfG1hi+hEkwMd64jukm5RBlZaNDVZIbr3XdGOo4yn1KQ4k8TPqNDuuB
wZX+iJk05CHrq3lFcn3mfNnpU7Wj+qojTj58oxN4R3OMgQszUV8W/L/m8/f0
GCwpUCY7YxRBf5ER0Sbc78FH6ULp1AZ6B7PlcABJXPW31apBiDAlt5ZT2Cxm
WTdjLMPCNVmpzm21Agy5m7Czvl6fSjgaZswYEi6OexBgzXaTXDKZbJm4OTTU
KVe+QUGRJIx6JDrQ+mLPupBMH0q2wY2n7ceJYertNXSkGJ59BMQlDzJhM/JW
cK0Xx1iSZp23LIWpmNX2saZozAS49QFZbXgoIwhTXjE281d5xOOMlEiaJozK
aInH7cFo8KKicOV/jehV1XXs/gnI0UAGPcZv+qM0RcxvBHquNp0WoL2PETpz
1O0RGFY8W+MV/G5brzZqfg6gC5kOV67rBTrQHNpDjchPhEmurJxV2UWcu6vr
WKtBQYdGTk/p7MZhlxS05/jRMnsE0y+gJ8X+0MfTn5eZhvtVllr7ROTQn/2z
pYcDfG2+C0Bi8GkegK75bSHHYeQFRug9Q50ZNzQ5TlVlwIQPQ+++WeTTatm+
HxGpPr2Ldk0AB3H4WEoCjtTq3Y59chmabg5edrQdCVHoZ60Yt34huxXgq5Yv
UnHFEVyQZpDKIEOU2JZkjAex/AnUHkRIqJX+XUJdC4kjU3MXXg7d51vlfJIm
ZVuCUN57WFtl1JjiMBpfb6nhkaX3ZtJA6Bkqs1/xS+Di3cy30/POMUxTh1k6
CLOu9Cwmkw2wEuSUH2uCPRBK1QvPKWmk4ciIuvVLeAceOyQX9/kp96O5s20+
pFc2yVbfMokn9teUKUQmkIGnjyVsUT3s45IWGWRKRU/1dsslKvJJTjcNBn2o
S75b1I9ey/Ly8EJfsZL/GnyDaivkFNr8Qf/S4hBHBpoEajescgeG1ATJ1MxX
TwPa/UDie3cOxVCgJukp25m+AYX5+MU0Tds0C6ZmdTfgXBdqqXHf9Nr5rJZI
fCeNw8dvhTTBkw039kymGck00DdYCDkyY3JgnXzqaijAFjsYyV2cpa7/RPfh
3nhz/oldYyMBy/W6eN4eieZIzMHCksfJz0GKxTAIG17QravScCwleddlDJlZ
cLh1IG5jXXBkPOFc5qA6Las1kYAaSOKUi0vD1PSMeDpp0Yv0c9qlz25J1+nL
8FFagWxyGIvh0HBP9DGK9yJ0LH9RAF4u8bDgjv4GdfpINcDgr2MpWygWx0yk
t8YXzcv0Ddz8ETKS+bY03ihBDE+BgDuV71XVoCrSY9SBJcLIE2P9UMrzvi1n
aCD5hiI5Nc6HrbxBjX6epoH/1QBl3LaAmM9lK5qKH3gAgQexMNcxCgtmDrPX
Zr7uCeJ2e6+LvfUrB/rtnbSSnELoNG2ZdMEVhgr+bqgrA8AiP8rfmiqAVLT4
d3ODmXcHl8GWw144YpiD9k6YrCYhip4ZOwz7jpjScz9LJWTVwkkBUcY2qw+B
d33osz3WZ0XeveGrEP1N3gdcek7jqJB4vgCAtt3+cG8gL/N4nzAmbdRC+xpE
vDkJUtxzlhtBbJNJuB5Ju72eHXAPdfhbNq2nRIs5i5t2FNnEQj8TZeTyEI7P
tasgCvEsFFfi0s3tBohddDoOelpmTq/eFAHpsuBfTaELsrUXu3CZcp02lyZx
8zEeQuWuiQs51dSKcVLYKZK8BxXnIAmI/EzmkM1x+QNjnPpTqKJ8+yW1v1m4
U7NBPtVCKkHe/LrF72oodUo0QCXdu4Cin06pqgE5ZDtjKj4gPKf0J5cPjyRF
ieyd11y7+iMHv3cExfq4vkDmMKWfxSsinBRVXA4CFZ+/VMIfrGbYWs6GiUti
sVNUU73STq5EQFNafF1LfM1eDx80AzZUsX6u0G8gnxS34ShL0aLx+W+2WNVu
oPlvvP1ue7J6qQkjnNa0DmzZeG7+FE7TkI1kyHpuGr57vW7aCyyLcSStfTyg
wLx86uxNMDM/OLCFb6dJrAA6VTvhgsSDX0Johyvss0z5nvAsjA1WwklUx2nf
wfLPoaoX7LtmaHEOPYc3627xDuMJRCcB5JBakHKLuUShVzZvFwEsPQeVuxib
dHjVaoXbPS5KxzhAP0rqurSlcumaU9Doa/1pZR59yIlxTmBkv/U8bmS8BiAl
MaeVairZ6GAGUYm7dcT+I8TKapA771M7iovrIokGcD+PKEtARmvFoIMQNnNw
hNTx6Y3TaCjGFlzrczJq8gRuaOT5hgxCfu2M0ItoMza5pAVR2xLzG/IshLi+
0i5pho3FnfRTVLI6/8nFkyGzrY5rXZkICWNHk1Ku9blujhpPoQu7aCk/tQxm
LINvmNKrWbrfiE1p54rW2vBQfe8MpM7Y+x9lG284QzKJGYa6854fYz4EodWv
u5nJtTqRhfmFexzapqNiNNk6j83Z7VE/CXIO+J7DZo8j8NFWU8qGvJiYkdeq
MeQlpIrQFJ2syTWXVbr4WCARUMjvszix0M0/cxa77gLjMG2BfqyR8AacDhzX
0lr9gWRaO5nac1aocrnAMy9jZOLAMvU7EN+bcW3CygYkWa4gKpWO/w2iC/n3
sWj6qfsaJP31Ae5e4dj6InWP973Om8TDgo4TvaDw3hNqQOupjbSosIgRlFHW
QIYGe5PeWfn0TZKvmoo1GcqhEuL3XS8SaSMspGA7nCo0xrSIpdAWJfxZegXN
zOa/C9qOFvHq/q5pnOC87ABNMDOH1YVmO08EEoT3TNLRlrCKkBG91uUpe8rB
s2XqJeqV9jU3QOtLlM4KN+ePh4cJy8i1COIf5goUrnih0EU1jVblm2cEBq6V
r5OsmUVEj0fWqE0OuHZH1Vx7m0iZnUOafcmga2jAh02njkceQIWRtjIYtCPx
jXpw0Rhz95hwvsI1L4ifgrZ/9V8LTbCIaqVi895UEsoJ3O/M8TZ5IQJq/RYw
ZDuRKybgHfRHMKjaOShlYY/YIOC5uZ/tFXl5XvKCPK4Rope5/sqwipyOPaJx
OudS8ehEJnQcOOvWqZ4FhNodS50PU6AEEGYNDa9jr3LP4gC6WSONph/yNbv1
3ItQWCHp3Qv2KBipeaJZk+LRyGJwPnvG+N50Ilnf+kojb0XtZ+rLfKKndV5q
x0iV+i26eIPMnu7W33GK4xhLAsxBKS3xw419BHgRu2jcadWHyW4KKKppanwt
03MAtep0BdiA4tIA+m6rAORTUAZUP8UNOcG86s1BsC/nO+jQmrWTpRtZp8zs
PD2s+IVku5mQWBEUARdPjekJAsM9bAiMjFyhNxn0Op6+v+pRte6YywMbD+Ox
s31xoRatbAjGZEoVgo8BpF+a5W355/Q9MPEX6tnt64PuD7YjXnIp6VoxSS5o
Hqoa97g2zzFJPkaKSmQ//yWhl9xYX/y8Lmhw5SQvZu1z6jQSL+wme+1L0e1s
9mEaE/lQ9TI2XARneTog01T7MlNOkwg9bBv7DZp5mDf8ysObBfMPRTPekfBA
xX22YjYUO0VbfIdNwm0UbXo1r5Hz0EjhdtRDZ/5zuXY14fqpRBkuHxLGJWBH
Z0eoWySYJ9WDEUx3l8Hca927p3dbjyslimdd/vjs+BV/saSfdOsM12kvVP+d
U7/V9mGFE5Ewv4Pi1RdkoHJWJt08E/geKZjfdL/OVljeWz5J7RNlRnpXYyYO
JP5hMK99kF6I4hnXyB0t19n2axlY2sSglXRo+vSj5U68ePa2uJfI150h1g7k
aA68fTMhkx4jBj7S/yn4FQ0dTjPhI0QaM5RIXcMhpH0UGRdL3737jy0qQKVO
KrE0uocIsPANzwdk1f/xp5Fw6p6e8Jdv/fZs20pifyTjoSFbHboR5fSHWHvI
FSAyRBt6PsHxyYmZSktkHj5Y2ZOYW3XRPF0JXvT8jb7+NtYxuqJplVk/H4Nn
srC7hAhM9fODTRKrWh63k3b7Ikj3qA4ty5FGHNyRxuG5XGetUF8ZK+6xEBpq
mHwxkCAQ8SfdbnKQdLZF9fIhksTajp9B/PqgIz25ivWXf0O3u5G/j6PQEVyN
mtObZfpodlQpGX7vOh9KcDp7MuwbRoNiv76VUycdTbjM2r1uYCi7DioOd84J
7gNH8Q8V0KUfmK7tzVL8dMFbOhEJZw9b/IIIMuVwFNl4yGnWFQ9pPYQiL2va
EW6PTA1Gjr/kB8NusRqt2XVOz957ot9QgVJSfSUufIBkYQyZIwNeJz06umfi
rY9aVuKnGCp9QKwrP1BwVBlqdwpX2T+2wGRN+J5pJqGjvx/uVhGTJ8rfFBnt
vjrsyW/HcMpNUmM1Bw5z2edbiFBu9ky3DvxYjHEAXG8XSxRlfptFunX8QGag
qCI22HF96K9vydIdhsTLBYdltOiC0uPsz+DMWg8tzdZcJSy4SwOO8z2SCNHv
64JCa7Y/KiPD3quLpVcVjrQ3FgSGEnMVAwFWA8Xwne/OUmTAwZqe5SBc7yWk
+HAcshYnuLDoxCw/Znr7eft2YLw5Rr5q6ZChA1WsPZQ9pZYWk6TMZ3TWaCTq
CXYhCo4y4VpI24uJXhNc1FzeCYyxLosQ9Ve0GYjc/yBBk/dK2FSpGasiH8Eo
0OrCTBHMZNz0IqJk7fo0/d3AJzJB8OwycRHKyqqMV0M68EwWqzlA95ADMw+i
6vmKxXPOPdazXLwP9NgWDuxXnvtunj5PyplJHktBDwBn8mMORGSXbe0y0JIP
zxZClaIzSg6Lcq5lh41ziETYUYblK//A2sDm3f8HRmA6ZGi+gtmYPmL3sd0X
ZvRSatmrHyVDWj8GD3V48KXB+xJHbvoNjL0UP1zPAW65YaVnyqqBq159fI/p
vK+XNKaz8ELbQz2E8y0iof42+IGwoO/yUNhikxuxNYfOOsHPAuP/SLvO8JJ2
X45QoxKZRf4yZfzDGNkrGdVwAPyMpdvtE/xYizJ4rzuFybtNIQnyrRfjyHM7
4kZGIpBmAD4X96usoLNBVO5sBU2bIvqruuEzXMtOiIpz7sPQBjRB24c/8P6J
OJ7yPWHSBe206bfCrvE47ufgdMwIUMTMjQE5PeLOK95v2aBu2RA6pbr4ZW2X
9iglhoDawf+M15c9pnosW4ctEevCYv8tWyYNfIHKLs6AiODvam9meK8u5t36
4HZJjg4Exe0rL6Z5FSjKrW8oHONN7s4HnIBJwFtGp/ZaFMy2rzdus0Kc1nJk
mmrt8q0v0woNgEbxUPva0Xn4Mk86IbT5kmK8/iL3J9LjKEJ+oXG8qsB7DcLL
hYHtJJn5W4QzMSnbHwG7gdI5MMQ2ZkRFKbMaY28u1cnltFYA1bfqW2uTEfox
y1N8gbgmfB5+Jr6IjFCRU9ynEMTxtSLWI2JdvrHJlOl0xo4TDXNYZsiXLFRl
ybPXmROHXoklqGUd2x+sIve/FEhENG3v9o4YjHyYEEzpBZt0+gF3suyn/ZI1
vJ0XuK+bVilBYYYwC7h4VFGe8Wp61oCDPLe2qXaKYrnO0MRoABRWz12piajj
Ut2v/uIIIAmevUUWFcN7fNhZouDgOiVaGswC+dxjQo58Eq8dijmJNuoqCruP
bmr566w56WDIcpt4VcWnDL8gzwQGgcCUIrPRKEO3BMZZHRNnDk8SKAkPJ6av
DaE4fYMLiDj/Of2moQj4pR/7sUcM7MVWd6dltbQ4DOjUTNi0CBkspP5CwKP2
Sm3lcyKOaKvRDeeiBY6fuXX9z/RA7F9kCuyI01C8zZQMyVKcz7SgUrDfaqBA
uHYJWLzfPmeh/xZm20q8ViXQHVS6CBs9JmaI82AqRJifQQxS/cbe08Iqhuvb
oL4m+G7TFt3P+M+Jf7qHcWP++/Pt3+WBGRumm7IrM/C1aavzXXpXECz08Vgy
XlYxsrEFQTnE1JFBy+jqaDl9QJcZPfIBjIILDUePDsTmDUS28BW3+Btmzdv1
NI6MfW8DDTUgpLAjrfRi25oiWwDbABLzG3GtIlzIYMX5+Wn+Thez5jcEY7S6
z+UNotsRbZPZ4HCEH5wCBgCwTPdet7OJk4ARcTCe7h6gOhgPe4eW7u/gAgn8
Pt5Iy6PmHjxivffarZ+FBDPJ4ZrqHQCME/rb3PPoR/+GBiyhaBINIlY4sAdZ
/4skcpyoulC+N7XKT8IKNOh2OeKgJvrxqV3zu4aXV9jdU8blIe8sXRZS2Lxs
I9G/PHLOt0W3I4KWc8wgf8tROaNrnTd5ug7jr8Vfq7Bm3NCchbpZqzd1Eh1b
kSKnb7SxpQ/ObppRicNcBMjmGqdPGzEvg0r2wO0lDhVuioA9y5i4QALys0YK
sNiw/Ui8IzyHyP45+7SzbJpRWwU8fV6wj1qG/X0IzD3gPctEkFM6brsJY3cP
nTNcXibi8zoeoS5i7RitF6bS5z6skUn1KGq3GBA7Pz1ygY5y/aqrZztvF7Fe
ubjpccf5wlBc6qt9Vm6nEnsIHaYxMaI61cBSPWhOY4/ADNwFXnmUq6L/r3B/
D/TpbQaIsjAUE+Kw8Wa0GSSapD9eUJ/bTfkQ0xfXCEZv2fgyQkjkoGe2faPI
Fyk1/pEPdW8qed3j0gJvcWq2F1SQoEnqqcHUUaiRkeGw0ZE9n5udHDjI3jSc
hnLropSjWy7/1bvGJuktycaB1UMyziZ2CtiN3+KJ6Fv9LS2Z71SEHCKWxolL
9O+9+U5g1trSjtCEatvL8O2DuFEizMVqSrXmh5OZAsK79IBbsW7Q6Le+hIb6
9LaoBjyGPi0zgtaPgG66wdAC4w1AK2Mvi7+2YeX2zWUDlOxvQmTtnTdpiTM0
r8WGQ3SE7wMnohZI5owEsX90sfiB8FwwlMcNxDA3t2NfwKQgeRwOBBmcPtSC
t1oLjJSwCjxkRguihGsqS1cOH4jrOPFfSBUGuHLj61Y5wNzwAVTSIZU08XJf
MNPRQzWlh+5uVpcWLxWkxYaKPu6cma5SYycCVc/r4wgHjyTRrs1aSdPYLLwB
8qpGkQSh/EQ9qrxZ0HCRRPr+69iAG4fBcMkjj2cF3bewFrwJlsYxeZKxfd/C
FVHYUFsYjTuLDZf8OVtsjixvpS6vatmtVnfANKh10JB0J39XoDyzlRq7p0Oo
IrHpgPsWKyEUcEJJvcPX4vtrHI+72Q5sduacEfNu7pZ7Nt69Cg0e2V3D6tWb
tkQ6ngRqQ1Mqy2UUB/Gl2E0na7w0uuNXX6y59NyuHQkkMGkKyZparbIAAJYu
4HheHCJ8Ht/hQP6/aRqjAGRjRCBvX0zIlyVcSwIrf9bvcdMAfgMIQIh7uHgB
WM6y8AOcO8ylZy3gbF2BukYHdz8DNz2Bdd1GF5rOuyFQWZw59Nx669tyTXBE
lcURNBf5FxrecHq/uO/wyDb8u9eobVs8vxk1P3/7IzR8VpqKwx5ZcHsI9aKB
eo3QJc+LP0SjDuQKzme6ZnrAzNbpdm2qCnRA+GMZVdLZSkDp5toMKHLsshs7
bpHEpujDoBQmJMKCvfbowhyAtQmMWBeiBJEcKWeNoDMSJOxzQ7ha2+kqbzNj
SpC+Peuno8VFyiAqp5nmr7ocuOaahdMT25qJ1X4ohLGWTdBJ2PwZpzKJqCRg
hvc17ljh0MhYQTVXYW9Bi3b2p2Gt5tRXBQ79d9DGarjYyYR5Fn1en3klnCtS
vVKMeOe7knjplYZUjGdOcg5qsbqnH820w+q++bVLM58ZO2O2ZO+YxKuvV5P6
8fZUwmFFH7WBDXiLEsKYjBpXtkD8CkGf/ZRLqInInXchRyi/JMeQrEgWTryT
ky2qZEM2p/cNDeBH0jO5R97HGne4ZRyAR2rV2uC4mYmt1oZ+P+AxLoEG1T5q
6wfmc+6DNWo+jrNVWMJJBg6BXNfdJK23Sa9aCcLHUPE4AHA6fLhvVRmKic20
DwVsShGtnlZMGNBxeFOMljOAnS664/k7vIVeIRbtXJOTVB8Va4ODR9ydt4XW
NcxYLB/CjHg5IiYjFEfd+jD1giVZMSA4il7nQVHagrMlZPwCtpYGVLPGdQmE
ykqIBMV4SX1ve7TcIOp7z1oi9HZQnL2fXQCgKXrTy7s+CG7e9wIvzaEG0p85
LR7TADuuVYU8XUhasjWJbSMS/njUwDeJkN6VGgV4DbQm5rg+ycGmYFpNSkj9
4IyPMoDGOp6yc9+OK5a7t2xVCEmTSMA7MpFdBjpCOUtK/s0pN2qzUK7/o0wt
5/w4hUiy/RXPbfskUy+plgSl2r3zabqp0fN+hjsAPcGA2eAhK/996h7jxTx2
7h9doT+Szo+dnGJ0Ihw5E81/T8KzhYv55ffI5OR8GrN+bskZNaVj2Jg+2h/R
mR7Z5tIwz+B9v9eDrzIxLzdUmWkSHTXRRTopqD208KEIS5JPRQN4gYztX5Rn
RvNf86+LlSR51vzHeI9Ip3fDYNqo8Vhbdv6lwl7ONAXkiR+Kpoqv5ulhh/vL
kUD98mh3QD3qQC1agEclXXOkQPl7xwIJVtSc2dvzA0r8CxfXNUPqBmAYZkSu
DWowIJ6ersQa28WkOHnJkIEKwENsHMEOghUykBL5EoxyevRCgJR/Pj7XRJub
qvffezX2V8uqM66tgVpuaFOdefGR5Yvnj58Aq/Wj7vNaMRTch3QfV+Mukvqy
9vXRk8auzO7XFoofmCuZ7ZVejSTIbnDfSLJzUTKZzMkUDMR4GfL09ZCW4f0s
8vPzzH6YNyY01anSJH4052ATfYJ83OZHNw5mpePMU0ENo15r5Yf/q8ekRzr2
2tbtrxMjHTHkTG6kNrfxQJSQNMjf6hNg9BmkdxinDPudl7lDJfAbdbofPaKb
cugc4H1gphH5CR4upOJXeVYkfzglSn5W30MM33tanS7iP6KDxEMGakmjISA1
/GElUcxHrs0OAktVDh6Hq8uLY+O6U+waqCE8LOPMHYXiFJZcr0DHgpai0Eg4
q/CnFZjNjxtIpu7lsMAJpOcHN7XTf+aVaCrkmQ93S4uUvaZiTwwjupMlcZ/r
JUK+4jlInnuO02d09ftwmb+34sRQSI1G+RiacP6afoNb7Z744j63TKHfqd9T
w56qoHIin5Sq+tRLYa1T5Dk16YyPRYUULd/NJk/GTKmXiN0M3A664xGabK93
18eZIRkvvPA251DQUtOnpUeFiQHZZU++dmkooPecgyqghQFtyPuayLoTlNK4
8PR36EVkE6kK1hWVvmVlqRRmzWJL+0tqoM2rC0W0KqTEqoo+RwG5KDPi1bi3
ih41O/wpbFewSo/eS1mCCijKbHA99QZbK61TG11o8vbvbl9GaEdBQYQSYrMB
8Xq3O78MEfGOjjFU1vKz8AF2vcv59705lliu1p/vycU3xUeiez2rA0NBb5WI
v2554ct5MXn/E160Ci8/QxDpZ2aOBrtSj6pMVOPWyNAo8pkJ4590H966EDbQ
FPR/09sYlpV4V/OkXewDO40Rxvwj0oOJ/41aOUkNU4IvVrMcnAP3d6WQ79l7
ueTe0TWwyyceYseJZMbfFBH24XtrcSka1dd5GLzB9adwovrp22HBe40ygz25
5CtsQPZ3m7Y9rjnbFs6d/tc6a2WChVeePbHTT1yhXgfraS/s6J+rywxqiw+4
dWB0+tuN+vCkRhnmEqAv8H7n/ZD/SjoJcnWFTLaljhDaNUQkBug1aLfd7Qiy
YcLG3vt3x+FQ6WD8ZjUU4oC/cNBINAvwAIqpFrRl7CQDShLcMNr+DU3pLVke
PLw9M7POmtZuylFaXg73N8sp8NV5uiGRglXXiE+tIkWHA1UKMypSJ3tPwUNL
2J/OtbKmQ8WJaR23GAqavsjG9+ecNMDBTWZcnJTPrv9dPjP4w29/5wN/J2sU
dLDOMTg9WNrNRF267WNGwOij6fRwDeWptv7mBRpkwlmjjh366NsHMiLG3PzY
Is2eLAsXoef294hiColL9gtDMY2AuZGnFTlpKCMeQtHflpDbC571CXFDpYG4
Qaz6B+q7Fr19QnVDn47qe4/914Eb/E9f0yIBSYj6rI0BCStYTG4NRGNaAVLO
Ap5L3nIhTz3l+wTRZfOckKbqTVFF05pIX0cLOkyecpiNAIKbio2qSdmTAsyu
UDPWd66BwaBW7T/DFR2xG8DBF3PQf8gyqldNvMXxVyoz7mBhDKUaaoEIkVzH
0BPU6THblgKU488L9uVuYiiV/26d7Ur8UQqhpkuxUrfGh2U/Uz4be4Fxdz6b
Nnvu1sOIr59O17YgtS/gbLyX/0XFVUwgr0SeyKatss8hlFsOH+6jJyN5+zrJ
xqFClW3bdVc0N/6xb0M/jgU9HdPQfmNnlL6nytCMPCAQjMnzpqD1PhjytKWo
8EHNq9hkcoSXiCUQomvz7kdm7FLkDmjwU1ODNxN+yfo8XCiJlNdsECHM0Rey
ucVw8+R8SS08T8aQ6oFzFRTOu1J/5pKYyZwnQse7N0dN+75lca79aMe5bTPO
PtzcJbK0lpYd37pjyKZF1PrEIoOuvrfe3pfbx0flHXTjjzuPgDEJklCk0+fO
xGWYMlF2Q6VIjXjrTtsnE8aaXfxRSAejw5r2IbQpIDr7Hh3kMq6qps110ikZ
h2sDS+lPvqZy7y4jBoiGscDd6Kpte+MtoaASbp6rED+7LL1Ht4z0suikJRPt
xYBYJNGOThVfimMl+ZytODNjj0yidiyCQ1GnXj+gnuce90DQVrXFoaLmlwT1
U6iTKWNoRc+9ZBVbEGVKYxJ+0qrY1GEjQn2/mkor+MxQBxEPX6Zlsn5NjegU
bzk5Ny9YLb+1Zt7jAk5N7Lb3LsMQJRrzOjXaO5OAggzFEBg5z6mqdoJdTpR9
4oqavMwax+xfjDhmDYC81NNbcRfczOyd7bbn6fXpZYZmmLpBQsd87+d9SN9Z
rZutuNf9Km1g3O6u28EIXDhLxWhsZg8NPbfh3ZmPxIm+l+cjApCaaUsMs5i7
XgVMk1nJa5Bn+URbBrXX4xSuDFOnHgE2239IPfH1XSqjgHIULj10jx4DkwpH
MJA58i1/ZM0q+fOKj8gMFQkhb+ZQTJTRPCGOSIgyBWAdufTdIauYoQxyEI1D
/PkpId1pySupg5G8drZ9RP2xYT1PY8H6+n6TrILe6CKrYVPeiqwL8zhVlMxr
fMLyoZkf57XydTKqJUYxBcu20VcIB34v/bFWx5RBzS9YGjocduKccfknfIPy
XdFP95u2nsqYn2f8TMxx51jePH1NR2wgbWHdRIeuxk+ZKaa/Wrr3fESlH0vs
pTzj6AdXmI2Afwv1C3CgOBP0Z+RFvMNqtw8LZZ1wVsiwbNhjUNIVtsVhk0dS
T0GKW6QIyMtlxCLS+smThuGko7ZEkdOCmPx5kqrEUCThSiLwxSEevodeL8+G
eT8VgR/1KsKkivfB4/ERdXVyJzsCjZirJd64GapT5XwLxSZbgQ37ZoeDHio4
6yNH10oJD3U0Q4afkkLWrmitMzDaTvTudEbb2IpzHgFJaaQ0kMoq6ULmJAUW
NQ6BIU+buxPmeXe8SvWUhj23+k08ZMp+Zu+vVAAECu6N3Np6FJ3uOB/xhDSS
EoL5kIZw3NK6/KurZekQzghG3X3WQ05u0FCJbPj7ctpyC7bxnm7gQIBueQ10
+p7ppndnjrfXO3MiKvij2d5Jx6uHxm4/kWUaqnzqP81Mw/fex628NQXNWOvb
hu5Y8hI7krZ4ps8BRefcO1F2FLQPMpU2VJ8TkxsdrvwAaNeKerCneK+erUYt
zTlI4tWk1lzhF2d9Dfmv5Y3NNNzrlXFgFfxjZY/jw02GzMAhPHwC3UUi49XE
2+O8s9vuchcgB/6R0rFjDz+AJG2xK0ihANgxX1R/8MHrJDwiaG+By3qoDpOy
yK2DfZtxvR+wRmz+aRUPBIJYKKI3cyjSfD49o8iv5+nP3PnFwIOdU69bjYaJ
o0cHPbsJWDUI7HrkfBlh3mwsucF3/JpUiqvLmX79VYYvJVAaxAmFDyUGFdkJ
wUM/QU2BEddyYFXsfB/a4WlKzo77rFhh0aiSvT+rDex5XQbHOGYw68HxK7pV
G9+SzDDWjKX4nPjwQOCwa4Npaw57EOsSTDOGUSm8y2Hsmo2yhKHG6fidLS9R
bGx0MfMjSjrPUnxh9yeJy3gmklVzuGeCcoigIOb0V2/ZpXQqGRva9hkn7W4I
G2lzfauq9j4eBdei7pCB5LbhEkfLzl+81ucb+27m8iAFmcimQKbH1SeQMkAl
LEb+2AE5DKAPEZpQgKjaJn9nOF+EkB7XPI2jvTxLz6qDDmHtx7WWgmmmkcAf
ARWzloTcwjLFUQIEDHXHth+YkutRvp+ObgoGIsU+1n6QnUwZMFhqnTF5l3/9
rBJrG1TPJMAaqNRlBSR0r2NK0UbKQ1ZiVY6J8PrQbozX8CszzJ+IFyu6nH3x
87+iyWZ+szt3tcrVcO0mno7EJsdM7BLqjVx58/f3IEYy5ztTpiVl9+tZsBRj
v6Y79uGqE1RSmPwy/UL3lNLP9DgBCC2FGfjUBTa/Ci847tgU3SHqf9rjAGlj
N+TcR9J+1B6XWNYS9fWMHNHC5itwTTZJodKpz2tRzUKlS4SE45ANjllLayRk
r8zp5ILWkOz53hms1Xkp1/44MAivY9NTwWcPygaUIPoYdiIKZZvecC0jjgWy
ZIG463PMnkWe2/zV7lzUvErx6uLb0584YLIXDq5+YK7Sh047TV1m6vNvizZW
mg6ywsv0WohbycHlobtu1PcFczJmrUVFiDszYM8txzusgMXHeMGGDuYiIFXP
cS/SvfRPTTxv30YwU9e6/lrSwhhVLt/v8eKSBoITECEMzFO/KalF1twG7OtL
/uNQ88JF53HpeJcUVVou8VzRslhuQWdDQ6PHxTn/GOanCLHg30suoNzLJFU/
Y3yu5gFW+mR8uGOMoR+2B0+cqqIszZe41FFxsw4iWesCPuCX2vUfbpLzhDcB
9sBLMbNfK9AlgtYsDPuotivPQn6c26RSsxLtVEWnucu0GV7wrWnaAYRZL7B2
pGCx72Xqz0WSHmz9D5DqQnd/DtmUFyzIzSV6FI2sB7AyYoiDfgT+jHcTKm84
tjMgfEDtF2K89SzZj8MYW5ZHThB5U1dh6cvKdKkpm1EdDJFDjOHecX3MtlI7
G+/jDCuRwVf1Jm1q9R3XsQNAP6UZ653Z9w1PqmiuRXfmEQeARQxfXLi3L+IV
62gE4e7kIWzwny5/PfRsxtjl2BrASnMOhbVxIzM8cPWhtxmW6mc1BtUC+chI
VVLGPV1iMte6tmz6420jWI+5+kaWPB8bbcNuAGxENY96jsq81q5BSz8KTNUH
mTjCw6o17muPDyxfDAmB6KUFVwqr8Sc28RlkJZaf7oRjXOdMZ8NgBf17YwKn
XDktGDhVUkM3dolboo+irWEdvKn6Q9cQC+wV7296fNyIkYYNNBQ2oCx2BpOa
NPIPz5cqiQBYNuN+Xz+zcO5TJtlycEpa696g4Gh/dBDiJ+5+jR9Zgsxntk8c
82xyxQ+h1osuYm4BmILsWx+sUKCB6PTi3R3G1AcnqHi8j1i9z7u2ZlaQ2+Pn
De7nKMSpYxngxv3H0OaQIvt+YQPEHEY6+GjSUiytYykIJ9bxh0fF+3Yus5N+
DZXu09mkM1bzSHnUHdDcnt59RSMQr/9Lnj7m27hVzuVeUsOUsHGqzTslRM4z
wEfLryM3N7hDz+hZthBL/JNuUZr3Vm3C1pR2XtMQ5+81iH+s1hAytca9EnE8
SyvGgAPUrnuSZC8pUGRuoAAymcYbItqI8wNo6fsLo7tBVh+DY8z9lMi5H2Fe
RVODqv0qYCGqOv8a/jUCt0xp0RyFlHUnGjw6OyZqsgzZ/ZILTOaGOF20fJ2+
2xt6weU8cV0+sOI8YSnG0t4MkWD5/OCyYaJm5JfqfqizbcwRsm0/AGodkgo2
hu3zG+hSwJTsQf6tff1mpsUHa1W1BeqMNAve5R8sRZoa0yYRbvN9w434zC9H
oU0RyucRnvbLkX5Z2Kzf6Q4gSrbnvkTdDKdsK5C+PGOqRqGIF5+G5OnrVvaY
Jddhj+cnBDePfVgZANuSKRnXvuLXWkuP7xHHXxXSC/mwAWpdiMMatBH/l6eX
LO0v1FVcQx/reiw3W4v3KCSo7pt9iVdyFwG84ENxKHVYXQZEilDvilNkrfkR
PlsNtXJSvXgwRALIxAoF5/giHNRa7f36oKCt6sA6sqtjMQaj20pn2ba1+voE
PubtpPYcmF8Oy393I/aYc1VdDd/58GHdcRN2eXGaq5S8klifkB/Y8f5dIl3f
IHB2d5yJmLbNv/QEIOYNjEz/0EKHb2WlVQ1KRPmzjlw2wthQL6KQ34TxNBfi
ZPo0orIS+M3rGT6nXLx711uqpglofTev7OydkWZPFg966vJpxPMHj3CWsolz
oJu2hixKfNyjYOqcmxtN3KMP7mzm1PQwddzYFrX3Psd1MDOrpq/7Y4zJESUb
ktnZcWXHvkW+9IjfGC1I65F+THKdWY9ZpDoqgL0zvHTunpRWj+keOVHFXMQ6
TNpx1xhBT7U+MMWFexP/BAg4VUacEQswqidaiN4p/2pKkcmmVG793I8UmRF7
XH1voM9Zxa++frygdebcEh2BiVdwc1ysHhxe0Hl9MrXYEtHglKPXeOVHNrpr
aULSvGeoppGt2oF82noCS7fM22qMpqvI/uNdBZkz2LQM/pKAKK5r1lf2qRSx
jINvWmiYdFVPtjrDG+WTM9y4QkZeXC6rZxi6Xc4plrofMjSYJ+oZJ532IT0C
pZ7OaRKeXKISrlD6pvZNyimG5Tg7WJL66Qedhj6DFN6jxRqJ7pZLGZMNxWZC
xsPuFadtAMyoUliQKMQWpck2mBLANt9zp8bRR9H+zyJFPB1kUnucK31ipYmY
eFZQuMUu1zzNHDcEjXy3rYafPxp8975lpCPN7ZbsreIWa1994opEM6d87KyV
EhkKPPv4hpne1svTzuOiYY3fqo2El5JxYdsiVCzrtABskAnKXRRLEzdofsmw
i56GZV8pcUlB/Ew1FIzBJrPJPBA4bZeZi4i0Ab4/+3Hwp+HS0CzW9J/nXdn6
ZoDHhkb9WxjfmZMjdYj2z/xr9HCqllLGJio2MppRqMN2eh8CEJMB1cMith7z
8AFWDhfeOr8DZWiNtpyFR51BMsIXpsuIlzbAb+Fb8HJVj9EbeW3yGCpnE+SH
zcYynU60GJOYaRbMaOnacj1yOVy88r45ZFKK1AY3aNF+/SqumF0qiHOWrFQs
mpE8LmfvsugcaoCfcuAP+KVDJksh06K/NexLRG7fqWe91yDLMk0T0R17WXQ0
qBF1kKR6562DrrB7sVD7KYyDgMR84kd1+EfYkzGBnV6C1C96eXXOELlYKIKE
O0ZkQIYpO3ZPsA1xpEJTGpEoEp55EmwL2b8tEEA35pRva2Eftukn5DFYKGox
o+sH4bicYo249af0izROfPcg4MVx8cIC/kuFdtUhkhriTYA3d3EFDxb36qZm
+myZUOgFhK9YKDs7W14KYPgp3piOzdFSWvqN4UWD+fiEIK6M3MnYKGqRd9Hz
/OsiOXVtUoZoalzwb5ND43CiUdax3FxUhtZuyzsYZQ++TMntMK7nYd8Ae/mb
FEAhwSipzti+8Kzr0z4Uu9bfe/30ebpLwq+naJ9ZIzQ4RcwBR5Hxu2Fs7pjy
cKhyz0/hPKmHmfgp7+t6yMhSQlz4cCkiuefE7AcT9jC0H4unVvXXV4xYAdr5
KtisWIlvCQR3BPW4lTvo2LUqkeceO1I3ul+4HmvibbjqwfrncmjcHyAi57VK
Mqh/Nsn4kXTWifSWzV0rxM1gnzL1hQXfZ8jGD9aEecmuqenoweNxs77GyrwF
v4fl+cPRdl5aZP0rhdfep23QXmUNWbWz+7ofj+gUf10ZNvzP/Tna0HBGqzvR
Xoqn+jHDCEHJo9iQDKfgQbq9Fguno96ZNXfc5HyeCm6wFMUhFeX0SEQHCWun
43mrGgntQ76BlC8riXzfWS30uvHZSFw0AFFCugyfVdKFc+8VDFGxnMuZdJi6
VUGDGwPVEC11JcOfM34GotRZbNrJPgC1pkSc8q9VnL/Yjfao2EzkWTkMVcC2
35YKNS9b2J8BvqJfS8jFvMVEyvk/yQKhJRTVQdJU3OT9zzv1DHpd5zc0Q60o
UpPa9/rimwg7tFHT0SZ5rP0tcE0gM7OqUAMSfo7dsFJBT/n3bBzV4n/biEVi
l3b5WCYMnB8y6/pShKO1i+2kLSzDwBoosowxKN+assluu7yr1OxhkU0lGb2u
nU7uxeg02+mQmFVBKzgA9bfecFh/pge9Q66KlW3vDESOGt2pmPR7PklQpzJ+
LN/Ycm575KGMJi0Dyqf4+7IWGSozSjMcdSSxho0Grk2Aw6gTs7toyvB13ojo
uNCk7YHnJUzurCqo0fV9mEliUobr3IYzvgOD3sQ0TRb+8A1uINEYwxYoOIpH
CYPOUOFb4FtjzaBoYDtYGlZbwid/cB3DpFP6ChforrzQffcm6JHCkued5luF
9e5KvtLc6NWOU2AldGGwEXsF5/QaKtctQTyXbIFL8x+m7qLfYNN1Nu8RWt3h
qNgz0dWW9eclRDOYpFbR1yYtMqTNvcFkd6qPGShXkLurksabjOYCJTFMuDIh
JuMklJHTIiUQh43ukhwmAWAXB5qOmqgUfxB/PoWDi1OWKSd115btRx6YKu4I
9KvsqeXR5rzA815QDge4oUfYDzy/qeZKp0poTiNISNVN0wVwSeRJeJg9Q48d
RSXvijMf66/LimCqNO991t6716YXl1TtR4FKPOjT4F+22Ss9Y/1E6xJXRO1m
NuyFWTScZk2Z/0zi3f3WU20wL4lla2Xy6fC2Too3jYoYRWpjAPvMWnxRsscl
VtMIZBMEOD5TZMb9CkyffLnEKn7xjPrRaeI2b18423OSRZqhWh75v13b1x+l
iyk+cK2PymuNUe7UR5jKMipU8Bnzrle3vwD+FbFO2fuzzPhQ2uDU/xi/F8SW
o3G8FeOv3PA/HU6/PjB5uuww9l59JhfNyO2jB/yIbUy60brf43B6aTCtLHIm
AXuoHjontTnTPAeA6zTweQR/rcSXZ/pED+4j5jTG0rX+yF3RIJhgt1BL1v+0
nWW3VAYpyP4Z+oCHHZzpkihw2gux2fjUg223BEjoQZ6Ao7rp5EH10FdNUch6
hjXbUDRogcSZU/USXaQcJPZth1aLR3KWA/vu+UxRiHFojqaFfSIWyjYHwUDE
YRFi56c02GNEKBbs6DKB4A6NuIhBhhbGwEft7kCWmMh5NO14tAC9/Xm0Qaaj
9wdDieDwN2n6VFMUFRjl6ST/HIhLGsq/0ZFsddDvAZDxqW+g2/ylhGXxj2ZY
7iknAFKnE1fkrgrR8Ow002XgmnyFb40l3UNYO9lxy+xCiQ4PmBfuUcacb+oY
AetQfFNtYGurHIqRKMsYnWxlqyH43KrRwmRMmD7KYHR6IQNdAtb9nPUC6Ljd
Hk7bqMPsDHiA1miKuvwmVIkgvXa29LRMa7FGKgIu/p6DBU6RF91cgttt9UAy
IsL9igX18MjNbboYJBeSB/uIhcV5JZjTmt4247VXG6pEx2nsvRalVTxkmX6W
j/lwrGgN/4LRLK+bSXCV+Qth+0ylUTF2X0vZqFrZN1mKc4+7Cpn1iLdC2geq
K5MSjj0M20KtOUuelaGyxrSwVA+Gt4mUfuZrqCxszyRDr0cv3dNy6Gzyjo2a
zVDvBxibsk1cMaKOq9cH6wnMU1qRiuh2zoY1uQlsaqB5hrDob2XgSXUFInfK
yWRl0z4JENlxCqGBV/jGxf3OSLKUi2/0VUkO3VXamO9HhKXEwOyzllUL6hNP
DZdZ8TS+YFJQ/c4CS4/pwJpT4jnnyKHpewnkpTw5Y/hN7oC0pYIlQT47PTLz
fU69SOYvwIbcDbrcFd5w6+NfL2RDDBpyvnOCwBOBOisyaIHtEtLxVYk1pvtM
zQkENgYXEF7HH05Arn3Eq6VvXjOnsaSqdWVV5swUmR0ziRQN9Q/XuSqoUQcB
xocCNxDI4+aEgax6NXrTj+i+dNXKIHst/JMpIg3lGwEcTYNcayJmEgKkBALH
BHXXYciOqkrC6BEJcGW7TZgrm3WxQBiIj/r68MP8opHk+0HQhv2NjjlkpkG5
blhq/GQkQEWGHAvhWGy+ugu5125ZLXY9B7MEpDvoPa04WgGCFnnYS6FDAs1I
3IJPTe2th1Qd7j6G4J7U6iyyerHHFntcjQN34Dbbib2p0ATirPJqDyMW5S8K
B2yAbgtW94ZRYJ2NMCPTh0spIRo6EDjhPpe/IkfrAEG9v2e77NBH2xRsOpaX
SquhjDlAf9Aw/01mmNuXyCZqkRP3wwE33KORWVvY9rjjdm/3UZeEgQsEmVs9
rG4JlEUU7OI3lSoX+kgglxmxbXQBzh1QQ3rESZ1O2d9/QzROq4D+qUBMqKJd
jktUJmOCIiQVN76XFtVUNEPWUd4aDf0hmDiEC/+H5sFbaaYfoV0ZzkEUj2sq
uuqyaOtAVV+2U0+3RdSTEpg17goESXy7UM9k96u+9XZsoFO58EL8MXdL4Thw
pvIloFkUL8g2LDZaiq2vSCJaZKDrgLpM3+W34MZvVgVSoQHJvTAGR4Ixj3k+
oGG+ef9cH7FxmU/KD2E7jycmPD/aWoS4/DgPtYjWOsluyH6Nn980xESDpU8O
A26tg/SFJevDqFbftTpVNR7RxGv8ITHdaGu1Fa9Tn5FqfgUdDtq7lsyj8Xwu
CJqZ0itOnGl7iajfYYErTKvDBkYFiDslZVW0LOwItn0kTF5VK4AGg2mOvIMe
uhqAIpygGGmJRQcnGqWzs3A/9MWMR8sJCSh9Rj+hril6Q5TlIJ6qnWe2MAfV
2yk2iU2l6MZR+AEplLuwqW0jn37J8cNDNoa8pklVt2P3aPAaN4Iz/yKKakQa
1ecgib1u1nJYuoLjyT3Q/xpIa0Ec6G2HHSwJ2wgnbo3QzWWb03XTDwNM08Gs
223Fs9/lGRIE6teyhU9UI1txnsVB1TkQpFz0NkzaW58O3wr8HTBUyOHWHy5j
TIewSABVFLArUsvTaMRmPRbQS9BFDDBafskSW3smdWjWDQDBiQ4hLG+Jj7DC
xetzDluqvR+qyKxzEHM8va/vyts+no7emyGH8getMQh3rL9t0HCgcAuCOeUr
iIG2VJsshx67Q1fCMGh/cH/eo8C+j0icj2bxE2T1BKU8qjBWIpN1vO34KZTU
ePdlkFcQALTJdjHSO0t7JrXsc2UWg0FmS9Nz4l5kwpDVN6SJyteiCMlQ3P3j
waI/YkVG1zJBkQ0alm4fbWE+En0e5m0MubrC7AZV5s3pr0FNgQXe5owpHJY1
kv3AE72ueRbrc+ZnG445Pmx5GxXke79jkVWKM8oLkL998Pic26l+fon1/DdG
wUX/Ta2Hd1hDrNJmvBFXa+8qioTxtp/CWQCEOvfBjBPYowruiiVcB6icWwIK
qGFiyj0yACG5n3hr0TKpOmV0sxSZ6GLDZ8u3xPGGidhJYsVFazdNYj/gP8+F
+UT8FvsR/mySwfj16Uwm15kTD9n5tYlJHDZv9NeYlEeblB87uqZyqdGJE6Mk
6QCzjY8VDGqs/jWJsBGIV6idYwb+jGGrP73qACtDKzH3SgNO6kxXYFJ3BINb
EKDA3RaS45Jk+S6368uv09oPLdp2FiS96uxEpoNQwcTwpGIckDfjhICoyZCJ
wWex1XqcMuhP6QgoLiVkIwUchRAX15jYwDbkIcAPHkUtcSYikwLiL/sqPZDV
tyeMG/dFSjSAkj+/9mPUhj9nhRhp9z9sTbcdVqLW6PTqC9Ia/S4+GpXk86LZ
eh3lgX1a7FzUghOJne44KKFF6euQc9YIn+7ri2b9Uw8dGug54bjAKowl9flE
4sVS76oMNRM6XXwJAR7BjsYoFFhTgMs/Hot/WwNb1ajLXdPrUOfdsjSrPLrs
R9ZeD0I/+JfT2Vq2bpUbbOTVFiWlqOoDwaJN02W33t6Y3Hdjqq5gkQfnCRyX
6TLPOP2JaWDTMVMNi/DMwz0UikcnPHdIfDQRH97pT8vZGLXjxn0oie+tHC5y
J1U2taPn5+UjXoEL+dCSQb5WDjtXKv9BhXZ0uvIqmnt0kaCv5L0KTxubiK6r
e3ZDQecuNoXa97OvECkkhcJAMon6DXKTxVQdTumhXhPHijCnLOL7TgETmbqi
d523SR1/2+LRpKyuuCguK6wNlbRSeVNBTq+IeFEhmRfVLpsHAlBY3qxANele
cq86GFT/12FSWIM+uTlG+JMaAQQ2n07a0Ka1o75qqaMTtoXI/VGDXw44XENa
pd11NmD8gbhEEO96pSMfBLek+6PDxHwwyreLF9cLduX/6N4o42wUuiQ5K0Yi
cIrWLrk9xHe8/2ZeE6ZStLqQ3DltV3ZG0c/rqgD2VKT5b/Ik5uW7zGYQ8BUG
QrJY9Hfql/iSlGW23ibF09ZrsWhkb8+j3GL804RDSJjpgSDVVjEIJXIN1guK
2fT2m9etQ7A/HxTzr/dld4Iz0uV56bamQ8h2OzSXJZILaSXlnLjZIjhy2UNJ
bF1ZFg5poizikhEn2eFvEPDKXdqhrDNzUHNw64uxiM6f1JmeK8LGCPh19Evi
nXoCRzzDwaSF875qwnmZlLNDW1x9jKcKyI2hhvpvSeKhet/We4MSAROo1Yc8
zhjgy1S1u61tXcQNvYDBsd0IM3gMHds2j6uTSyOACHLU3y4fckCwy1fk31sv
bZlTUTW9UvGraKJcM84801OPSUmj3mlhEYS3VKVZTll8wmZPgxLmofawSZhL
X+n89wTcOBgbDGunwAC7DZuKnxzDQyEUdi0H6uDL5vw1P3c9ZILM+TNrDGTA
RKDSdBf8bKaV1R1zKFZgyvKjAvrwFY1C/r6eLJzlwlqKB9gNgO4mRSog/VKC
JAFufWQLoRY+Qtn5Fc8B5IAM0Ed0soOGjDFsGfCU8sPIk17z2qEl/AIC3Xl8
AVPU90sN0CkMyAGQtqcaFtbBAyHCvzj9SMSLgjLVZIK/S86iu4VvO9HOVyTB
UeT72t0BmNkjMLniinvgZPVlKM4Y0O65rYk9WTj+Wsm+8XfsrAnvr/uAf36a
41amhtDX/eu5CMMVPlL3htSU8VPRoW/52YR7lFZe7lKJG6osomdz4pgIiPWU
fuoTSxR9he8eoYPmJT0vdh0tEhaOdNzwIHxal0q64TCRQqnf77dCMmxqD6Nx
rji0+RP4QsMqyWRt+QIBfGKLzls1MQAsC8SD2RNnV6g1sf/9pxCtSw3YSwQR
iOQqBnnfWW/b4t9l5YO9tVL0xrS37WQXScDW4bmVkUGb9Un92rUhxH8pua3k
P6V1VJTI6Gy/40Nnx3f7+cs8RoHV3MgkcZfgX8t6x1I110kV2ZuiUxTDW2oW
3lZWq33WNUQ1YFWIF/KFiBK1Oh0kAPjfGARieqyy9TFWZmATLjhVtYw0bwJF
fWNxdU+yQ5ga0wuKiXRl0flj2NIsVxFN7x2XF/sQXFdWdlwub35mLbh0+p2B
jO4h+/YCDycpqwoE6p4LCGbrkneYGbpKJKXH2hiRheBYlLr2mk6HkZT9lM1C
3rUGFhcylruSp1jF+Bnj9q814uXkxAk7CsK/S2f1QVS2VKBA1T83rgbTSImT
3+bLG9x4RmnBbATyCrpPIBC8+x4OP4DRq+zSQ4lHw3FLlX760xaE9zEEkFtd
TRnMkH20tztIzV+w7DVkzr5il95NPaNzLhQxOGhPl+p0ck3loBOLhKwk+PBw
cSqtE52XynG9YlqBW1dGjkHVhDd0Hp/sR65WTtqgLApEMRqN+GdbEftNSxeQ
5CBjtR0uP67/DotkwuUi0n1FeEqeY2bSG91pseNotw6UwSKxlhx8TIZiXs9q
dgK3zPzsYxRool8C72Jgh/1QgJMtZEyctEkyH2BHqswq4ucPi0avClxt5cjE
PCfZngkUeMIcz/2zPbaxXo+x5xYDcgy1qp/rwXNGelkf77b0cyBCcj6w4Cul
pS3yDSa4/Yf9mSbKY3ImeElW9jppgPrBylkUZPiHoBHx9VVM0jL2PQtjwilo
w42H04yOJGr9szT1lgKfPVLAegxfgcWPVaRiRJk+2MXR/ylXCg/LSS7Plljy
oJDgp71+7ez65wj0M+Aiw2NjVnXnn75CTT6ZM21xbMtWMoTC4MdHiYKF4KVT
Gs/Ws0fZloY9um5ukINwUTSAOH52xVrgavXVN+tm7QINwuQL9lOYJb1xdYgn
jMohbA8Xkhkg92M4OrgnFgVdm6K/ybqOBtQSbCMhbgbAFPqp802PTaDLs0ui
LEJyl3Ystldp3dY14GE2tQQ2X5RheylG1JwqtBW8JwbNI8e3A6WbPwqjALFL
tqNsjXYpttYzWU/oM4efGpcj+OOprACCdPNvrUgR3V2js8lUB/2478ROJHK3
6IvKCSAC2WJPUl32xsGiMGxyr6zo2VH4Z/5tmkDMmLzQUNe+PmPXCu8Dyjqo
WnPEWnhs6stc0QKzERgjrXYCPNKIw59wMHuPZYTGuBzllBY5AqcftC9lw7Hy
bNj7odW4Ftcnb9XLM7WVs/lZiDlOKfGqfQFXbAC3k58Xs1Diew/EOwModmJk
nLnVjyoiUwXQbMYL+OKudjI7sZQGgT45xom8PsB7WA7G8aIe0/JB7wcvMNlY
RSisivUIUATi2EpcSNl/2KPpGhF41iHXBoUW25IDhr16IOxLExGpIWQP8k11
2DQRCNWEcshSWSOIw++xmYEfKaALCRg/jOwHv3vVXqtiy1Hi+KYgeClZp13M
w/6ES5uOj+jpMBE5CVZnhE3s4SfaB3j+Kdko4OzWNXS4j3UMU0Z3OctemK2b
08fBYkHDlucLuWsQWwBEtlyZSfEnmFCqX3ia4kWVFITTj9dgX3z9gSRutHQF
ESfah4fRFK0EHe0teP6PwNcGpGUUqx3hsVrA8U1GsuvnC5r0TI4AfXK+GgnN
eJmD8gSU1+YM4t49kH9ohpL630Eak+6y/Rbw6xzOAD9DjmMOIROd1fAZuNSf
knhccEokmht9koeqTU5zkZaTSs1PrFBajzcwBinURs4VyvxUKyUuSfjrUltI
JniA+XWSZULObUh5eYK7B2iEUGuyFqL+cZN1YrN2HimMLOjwUHxRkGcCN4Rl
xALuJm9xxYY+3DU1bQj3UcJ8EusEAB0hLq9vduGQDfbRhzNmZfjnB8VupG3k
WVYXKczf4kh+9TBv9wsEiFLQ9NZHHMWTLCwsBoaHDDiu/NpzkglPZbL4ga3V
bObcLOHwY/S2JLKEZcTxaWl6WF+cTbV9uEuMROqBZA6NWJtONU+aSD5Htu4B
mbUYBaYpLMIR6asxf+q5bpNtNUR0WQPSF7XNDNUFzzgg9xmg2HBxhrXf2AhZ
QOThl+0QufW/GfYDyHyM/rP9bf5u6YxJKqpPeaIDK72s/zDbzSp8AdKUVpXm
Z+ktB/1jPAzijm4czUUtmuZW8ZVGNpPxs3n9fEN/vcOrYDwWiZK6XiwMtjyZ
ULwPO5jDDafeNGzYPkrgQi8wiSVsxaHjPe+r0Yplca0oIYUWAh+L0CKWNSL0
AnZrcJdyOs5CFRwX0um/6AvkSyd04YEGmDCm1k1JYCjIG33HmgccvSvjgV6h
GAgGL1GRCH+BnKonuU8H3tYbtDpgTsxno2/vqUoSObR1g+j78T7K/eUUn2hd
XpwH3UDm7UJHXaYVn2iEXDtWDkDA6vUnNMezbH08/i7VbkIz9mSgUxTLJ/R/
sm2pYdN1y3XtNUvQPacjV6BHm98XgJR9bkYxXUl6jMnMEA4pSRLQkZzjErzS
+gHbAll6wzr9d9YDSIG+QKRVhVFMqlygeBQJa9S0o/Hiel33pYL0hm+bq+/A
RCDXHWoNDXzksMjVL7yLgMU+MtBfQBXRT+TW9m9qYjXdwuGBVrdsjIXoMxGh
N0eiNQ0R8X7N5tA89Lq1U5fp0HA6HrMWsDG0QFm87TB2gZLwRTWwUaT0cX38
C50MjAkGKaFRlegRphGd/oqU2a1pQ0GLcn6mMT83YfNNH3ODCsr42qTN6gro
jjEl/RtHk5MLvk0PUC8xWFpxPljI0icpK9PO6ZpJ0L2ktCjAwcb5w7PlmqQ+
ktDboOjPq7CrVVEyKaD7/OJmGREKXdEdxaP7NGbAMzy4JbHRI4G9VdcrHbLg
Wec0b+QQgyTQU2Ok+3hfEBul88Y3IhPcy0S4/x0mGjdnX+aQRR5h9BkFzUGi
xIiGPQkaoCBO+lEMUXH/kyj0SgsOqTy7DVfWMyequHwhoUojtIjDfkdHfLau
Sp9eN7SxVrl0e0CBe7K2PEmP6wiI93cwKEVKeVOxVA6l6P8TczzVjCK3KQVC
WZNcEWSkBSLOe292zbCasa31VYLvatC1Zqji4lLNqeIVbKgUoXv0eFADzvw8
ueT+HhNXBDps6vZRiKw8k0i+DhKPMnWaigsWo2aacqqslE1uuBL2y8Ov63N4
i9RQRatGSGnK9tL8YKoAfoBLt6iQNvRNDGTEWyulzYwFC+cnyBb7d40CLxO2
Uongq83JI32gmSm0Kn0+3VoprJpFg1e6U2EMLkS4NVc4S6A+twcKlhuxO7Xr
3e+PSUMD4Pdl+gyRtiUPMQHhavnBivQEkeI+AMRLtB6kbKNw91lGX0jviQy5
ozefwh3ZscvGKslMlXDUV3MS6siC/jTugxQN56CeisTBl7220zLl66i32WM+
tbWBxKzQ454CYpfyoGi37ctKfY8n2OiHRRL6fVkBfFPdyLzIcAqvGcl9mLlW
FB7OxBOTUUUO4eYmS5CClxo8eFJOE2pC5WraDPIkgv1L9L3TEjwdWHbOEsJa
9HzthI4/jUN4+1603B/z55/YG+kSRPX03iVJTGOAFWNETn26RnLvI0nAPLK9
G7OtQWQHuwK7fM7nqOy1eljRYUhDzUACDT9HJ3XYM7VbSUMMDFUeQccg+4Hl
7bFh6nKOSc6cANX4xlDgIxYjkyyO9eJn0qII8aE6Fejka9k4utM5Xb2podSV
UZQn+Fp+J5YkQ00OiZ0MB13mTGld4sRhwnv1P+qYiSPLHupVhxHeq6mS50Pd
Lax376PZZrjdfI5FYJmh0+DMj4y4Z8BR2zSFf9kdsXDsjeb+NWqOcrfN+5CG
zmjVxlsV1VrD5+7J+SqHYooG/HonUetTntHHsTvZrz0DavAZHQ9GlmOtGQqp
N9FxhbWEocVne9uW/DzG1rh21l3dNiEguEYsr2mIhn4YjCqt76XY6iI2cfNK
XaWzoJOfygERzdvC2BqrBdiw+3Y39QK7Ik+oYFPazfmz8dfwI0kCK8UQk9ec
8lUZRlc6+ThAcxX64toyneKzXL6JxpITDuIw6jTr4snQSfK4nT8NuuQR/EJT
p7QzCsy+3dv+eaoOxkiO0yIUKNizW+U4hAks3Gg7jidg0GCHqBCd7UGYzCRX
AJVVNlbEIujR5gIffEPteOiGKxSwUED68PXUG/6pzhaLiXXJTMDyrtuB0oAP
cCrcCBCkPtXdXhyXoWqj81gA4JMCWxoxvu4y3jkLb0moHZsRbLc62Lm28OiY
sbwjTswixBmV4yugeeMaEebGKPpkUaVYAFuTUSUTBP3lIFxZ0bc6G2FVWLN/
gZfHYLuZvq83/VUQgnAi+TxWegrYZW1a/HVEsvBGCfVvJtEHGTWsv7Oe9kxE
QrZXxfU9Q24KTNo3nWcWnL82yq8IEd0nIgV/rnY087mbNAfU0o5WCviwQ3co
E6T6CKuk954O7Zc5QQQv7F6ucH03Z9qqnfIth/3Fl21qUnu/Zf8pcP//JNbZ
Eh2HCZKpWfPhfnbR6wY+/KiaLZLpfZYrTvzF1pMdzCvSPs9sQslbSvlul6iU
A2ZyGCnowhY1P5vwTWr4bRAiJGdqUZUfbjoi+KqH+CjIQAMtPwwZfxLhR9PK
jUF3jrPdXduwsWD97s/GjgPr22w3K798l+6G/ciWtB3V3S+KbECZOboDrVM6
FRdZg8u0o5zJjMdLJBhsFNwvgWJ5IgAPXGahiaFUnbHKFiCB7ot4PeqS1FnH
qX6A+glCGr2JY/kgh99LRsi0PuPDLRlRCwr8Dm26uQ43EbqzoX3mEissf4G5
xJUqINgW87X3CGWPFK+dzzHoTkOSbSDUlBqGAuAl4t40MQovkr9SUg+8XaF0
Mnx264tWMbmxjn+O9v/9sNVLwtIJjsTEXRv7lEFWvO+JKLxVWmKEeqLW357O
LWKZp9Vj+GOQbzS6eIbmmcde2KYb+iHgOulQXFKnBYzjbtF08r36oPvLmuF7
xrvj+QMW6C5phN8jWe08sFxOn8UNSnLlpZMlf4b3dvwGJc/OgyirPVPKXPfY
R37W9KKw/ufcVzSKGB0ogDrIpqcwfdfQO+opFaIGp2TzgP4yMX5c8juDxrsW
iRcucTkcLEc87+2sOtU+cpO53iRuXYQ9KVPlbozN8GVXMY7JGQCd8/dWjTWG
GhJLsdXna5Y8StpVmeUVf6qQov1QL08sOih2JBe3GF/b5PswgNhJkNOsykuP
27lRWLjOE7rof3Lj6HcMRNmRHc9bWLSqybI/4Zf1KYzyVPwBfHbuvjVihd4F
keeTdDA9JSlJW48NBIoYP9BkLVYZp+oqV293S9AmRvbApRJLrfN42HNZ/iNP
KGIw4SN+pjtWu7nTPS1eKDdZqVkaYVnK0ZGonjIlSsit20yhcEEBXiwcl15w
3/1yIM6/Fz8cqCWYiJIPr4CyfKqzl/ixFRZ5PAl6F5QSSnM2fI6OZE3M3RhB
ANmZbbIu+GCyKFXq5Mk+SjFnSZnENggiSqECEcefdfkFGspDejc+Bf9oveHR
CZ98nd1iSuf9Tu2WMOTdY2I1abv1EFySC6VqTMwuOfjmYYYsAAuW5Q69ohdF
CB7KhdfFjmB0r6LdN0BFugIdiSnHMql+8PioVQ8tQoGj8uWBcibwhlev04AF
eK7Xotz9YTkrSMudXi/HMDyYe3tHwraIhrHLcvIea82fKVmUIrhr7tFfJQIh
UASlDKm2i895KK6wQjR31laU6A+P1jaYfHZDxkYLsZBaPBv8xF2cvhhsT5+4
pj48gbhdj7Hy6uOoJYBDuJoMjtKdCkWM+A1r/ubxboBl5dA+VZIMqdR41GGA
yn2iZIGYDneHSqGFkOrRkYyAtEiN8xuMBHiqYVfYedC3Aejea1lDMESsNtsf
XcOUCHLzSrQwfEB4o2eNdZehKoOivsJTQ/lC5VsNzvV4OhjGATxN7UXN9V+s
uIMtaihLnGsslgaCcLniw/ATwMfqC6qMpmrma3wzDzGg/xyQO53TbjgaSDM+
JnVHXKplMFxo0GuZNf5YRTANcv+jiTOyXmPgEBzijIXQQz5z2IXFrSr8Ft7E
DSGGysgUxpDt2gyGjkweyqMpdQuYEDElk3eBqlniCdJIHnQ+kRpgW70T5N9Y
lENZJu6Q4+NuJ28F4ItMnKUqSCqP/HWFVNZEBmHi4O3TmajRbdgGkyO5lNx/
nKamXMcF9VjWABS737NAzMVplBByn4DAejEawP6ORmwMDhOlL82OhVnguBxg
GHCiPOdIy/X3o/LmI42eHuF0uy8RC4FbTYDwihspfytGfRHFm0sjChb4zSot
R9rG5KBtsGhuJ18YubWpzQ6VsrkhrqF4gxLatrhfp+w944ACY1ooqGL1AUZB
rIJysKFDdg8DgNaJEfHViGD9cijGBzulssV97I2yUhIVm6OAuRnJcZrA4YbV
4z+vL1TWI18nmBACwulLsmigwZe2q2dGY2U9CbAu5JjfwFE8GjOtsW9gMieo
qXYNlEkuEuZjoKKIkY6xafxsw8UeBBUNEvmrqB3UY4QoHY0o4gKA9NRgYuz0
1pTBERs3ELKCVnUPJIhE5mpCkSTu7rdhy3alw+iDchy1xXldJwyxeYDs/wKV
Uz1strB224foS1N0PTbCjIel5MUXzi7Hn2DVERCmGiADaKRis6ZYL2Zs+uJP
0Xfz3EOr+fO02U1Fn+GgJ3vq7TbDpVGxO1DxSILgXS3qXfmJioQGhn8Jf3mw
PrC/u6ZHXpVfX1gY4oSf0wrJOEB2irGUFeowbwbJfFJLt/HesoL1B5VyY9O6
TU9g6LVJ3Wea0TmW2T3PCo6/YMUynoIGc995+oSnLwN8t47WtKk4b9dr1mjJ
Vmc+zy+MdMa1fO7o3/nAdAEC5mcQyTi9ntPE8K3OmSMmtvYa6Jd2Nm5VxS5E
SJGl1OROMprUQpreBy/MhdhsjkuwxWsG1fqu8JM6PB85AnRuLgEQQnZtMiKg
jjzOYeDSIjCBGxK9bb0Bslsske7ZWPtzalNzGxQOFCu0LG/E7hdu1rdShdcY
cxwi89uBaMSKlXEUiUvaUqOfAvzdv7T7KP0YlLVa30F3t4sAPbrMPJy1VicL
y/rrZD1Su4uOwslg3Ahg0VtPbwG2BC98sbH7WaXI5WSNOaM8wBTs9QvU44M+
yOJSSBHVCdWVqcUMJLceNJML0BRE37H3Z1ZTTWMhaxugkMQO6vBqL4XGQuv4
PxsQxvSsmWRjWCT8gO5frYBwp4ORz+fpmIkjxJ6emMEDeLnW0r3d6Lj/Vtej
Fh1T0yqhboEUp/u2RexfD2059CwtyjwldNdKAZV/9nhGsEqqg3hTPyEi44Vo
WjT6bUEj6gRD2O464/k5gj2bSs2cgYSSf7uBgKjtcEspRBNuE/ndi1neYQUu
4z8KQCG47hM51qV4yyuKrSS8iAK0mZVMngLc/gi7xabmSMIAW/79mgIOWegf
pxvFjgHRNc1S1Rw6o7N6S4hUz6pRZaxzQFRaNA2HKQJbnKFaD3R/WUHxNf7M
RcNe3tnZLhyL28iPt3Nyet9jcE6Z/PA6BgZj6rUKVcNDH7K56KdVIVjh9Gcb
RDLQMBDIG16D8OETvpWjYKzQYn4KAJB+lfcmy+dfq8XYfL77iusc3dbXvJzM
8yQFsAWLZuRZqi+qLQ0uvhgYTMrzsoA6jMn8crXOcbiJxO0Vaf0jBlfHW0Ge
F6A0q//kCCdPRJAdPvtP9gQ5mC7LVjbNH46Z9WkXtfXye4oSJ/cdj9J9GmPR
mhUX99h6XZU2HFqjdXkk8YtGtk6NiYt0e5UNxaooBsPUZs8nQuFmFmFZkAbE
lPfFUXYd8c6MomtahR3NkQBjURVX3ZGqX013hbmgWXCItOLumd5A0MDnTl1i
DNbP2aBVry5nPNwk9cBwMjdVHJqVpMfgGh3NPRTl4cEZP9mTUwBMEpNvzvTH
SQA1mVLj+vJefBTBMT8DChM9l7tPI7y75gToDqI13GQl56CRIzwdCMA06vF0
3SK8n6IyuCpGXUbCaQ4CGwyjbAaCUG+aOWJVQUbsIXY/2Y4Yot7wqTeDDXs1
ZB6MKhjC1QoEEAoyOzncaCit4ouA97Uk/mKtqoRXuAoojevojRU1O+xFwhKO
sgGFeJXt63zvogk17tPWrCFj9Gju3z8xsVNAUGrbO0p5qLXblTA0egiTK3u5
AfVCjTKkf1nYba415ykj2LEKsIrjxnh/vQ4A+dI3Uz/MWssL6zx2WaGiO3/a
lz/Yq+I3blzClqjelMVRuZqg/tJurJgNkxf5f1YXocarvtiJQxBqsXP7T2Tw
XdN3uHkMJOuXN+vBm8TAYrcZwk/5x0fjkGhR+SK+kOXMv0ur3grP2NDPB621
Hs4cV9IdTgHsnfEcwCyWvFq3tIvLTBd0O9nJwuREWkt2JrJrw8moX8U13Tet
ob+46YrSiMc1oM1aY5fvyPcB9GbBxyFH7Er4I79DuQmM36OqRezp8HYyF7ch
dRInxQFM0FwZrsj2R6vEKahcoKd1y5GdgraPQbbRh2EYkP6VXSTIHfaFvsIj
r7/VlaZ/1W/uabKUbn+UaEWhvq6BELWBwYPm7xXHY6yEjS+FHXH6Q67yD+fE
gxcme4VuBrDghUtLKBLuGokhrk9ashDnju1WPCAvdpw78J3DEE/0duoNJvBT
cUUkDa0wcNPL+2UweKYEeam6CmpIrES36OiDWdihUgnF682NnOmMU5GBq2Ir
Nd6+G1chyQyQUq3qN7MYV8VGoqD9J2xKXCCTUjNTUr9lEjqGu3kRkrTIGV2c
aOUlaTnu/JRKmJDvb8+NS6+rbk06LfAoV66F3EGJPjTlii24gg19meorTl3c
M1gVMpi65dt5jvqpE+zHDcKncTOz8c9V3DKi8JjPV2J5jOcuPKTHSATSc5gt
nqLhsGxXFctYPxBicAuK3mQGOopfWuVndw6wvacIu7gd9BwfFitIjYvjtXLx
pT5fQYy3SqDDN+hAYGRN1182DMy+VvOGLQNzjyX7xYJkVFVqV3VmMrXa4v3t
r7HtgQa294p83u7ejkJMGomQCabwHwIvNqO+fghUTzIn9Suz5V33S2KgoXGD
Ii6HQazTeLNeJ0cYTFdVsxwXH5bJpqG8909iSO6o/HyF2gQYYF0aDOdIf2Mp
MCZCPpdAWlb5H1Q3lDgjtQ2A1TEPTTgL5Ut5UWdwCjx+2mezArOAjLe/3nx/
xB3um/3Fq9sGufTo9FEKeZad0cPfLKkgbheJLjSElTonxGvA9cciebDfHfAo
U0W1TYSFIkBDsKCyBu0kHk3bCMwmYjDlmWazWq52jOuB/aKGlyBITZk3FAX5
5Z8ps+WPP7cWhWeETBmeK9C37Qdu/Nvx7/Dz0aDqTpd2xN610I7A1UotFu2Y
mMz5nqa2k0rUVxigw0lMSMaosV5V4P9eq4oEpW6Uiq4SCxemnb4cu5gf09Pq
KwgNq3n70h5p9cm319IpzgHKAuvKVVj1mTux7DWDiArjOuIYltrMwWGgCF0K
+UpSm+EigrdeusWyv/fbx6SoMZLQOqf7/2ZIE0R/sKSQaByeN4RW+Bd9yHNg
b91ToZysf4nRyKh4yUmArdzW1PpFXJA761uYnghYlgM2jAfn4OSQlWctlegI
Oudr9st3v4QjPYUIb6fA6jYqYodwIZrrJTXW08nx31jsyHQ/fnguySt2x4Oy
FGY6fhLMfONdOTxFEMj8cSbHB8GJibaeyv2DcIi/7rSOEpmPkNI9rR8K91W3
3xVhEc0Ke0iAuSDXOeCWjtdMx+r4OvTDFHwv7ySiTTQgL5rWPnBWbaVKWM+3
gN38iNWblITWn7jwD+2Gp2yK9yY3h9LWMSAZtjmXYX2+1pd2k2zKFc4Vn5bx
SpcYjgvSK/M9SgMCl4LBY1aPkJbuWl9gIPnT7ARfsL2K6QYfxjP7b+ehbDpE
2Rm1fin+pRoxt+rmeR38HBGbYf9CJcguY7/Q9ItTbw0wuWoW2BnBc7PTq6Dk
fVm7wSAiKSYPHEQVCk/0MJnI8muQgZxJgNV5DYYrk/SOEk9DP+wML85QbDZ3
v29p8ucPgXin7oUeuooDC5k2j/aLyoYRQg+ET8cfIflDSmLKD5zXk7sw02nf
ukXTuMud7Uj5JhbE5jAcKT1WE+HN+TDt6T5KanrYjdI+5FvF9DcpRb8qZ3k9
Ui4UkVE+ASFpMzH7GdjOVwupcpVq8jn3GlP8zNpMx3O2jXt9fHxsnxD32/+S
rnngIuquff9BJelCndHqvahf8/kTVwSa/e4I6G9yzUdhNkWC66oJlzRYnLlJ
QthW2mAbttDlYWmfNOaaPeE36A27jq3XF3iZZDUSE0e74sCTpFIDlSucpwGe
+HMtJI9ZZ4vkCvd9mYfpmFDMSlfEekpjR+EI9q9jhqTJWedzjBHu0OY2ch+M
ullPQ0pJ/pvOshE4woNmLB3IHVJoBGUct3+eqPUe3Td79H/D1VRdiJfx+Pu7
+tQhbhwZ0JwzK1NZY1bDjETM+YNesalJW08p4cJOgycnCifTrdGBmIjd4OFE
9s4pQgCD9g4dEi1n+9aS+TSumfQ2eEIsWD37duXLLAjFBPm6CjpuJHEXgYR5
D1yv8p2Uthq8YPxUniRm3Py5q9JWBxUK8c1oY0gq5ijHLkNPV5vi/QYd+WbB
4nbL2XlYOo3ladNxXp2bZsQpWRrbt3nZKxkl3Lf9g5dBJysL8eSMq55/Jrju
Uc7NT+toJ1PhyqYKx4GsLpdCn6dCEGE+6ESqpSf+mf2Xav4k0y+siU2AhqH2
g4k4OYOOB2oLew/+j2SDlMlTFrMtnjraW4o4mNvKef04I91L+nSF1o5NBtK1
i6Kq2YPBZO8MA2w3mHeY2bSybytMhNgAeKjTBzPATOgg7nctnBBDqC3bYXnF
zvw1waa10/XaafjqfZxI7odI+TL/BQVyJn+SEVkPponrmyv/aboczJg6jC/5
Qryy67m8wBPGgUa0U+Ghyg0GzQQP0advC3j1HK0uIGx6pN4wJS9mG3ztxj/j
1yOmM90PbtBlKKKtmtjSHFEVAA6AKYdxjtqpTsnFdM0kXttsuTU45U7o1LQH
GhIOskb51/k5zf1cQrPpUij6FhVb3DnNVgW0urrumkmVGTqX/2aJNOYVIlT7
eH3120IjrpmOA1VTbh1v5n7N6jiXGR6SXw9AujsR2IjUQ1JgjkrWooQbZilJ
oqBnvbol4T7KceAdDa2VGjW0wu/Dfw1jp1Pk91SNfIVgyZBhBpOMluQPYnoP
bB2ReziZj/vlCZWhbtDj58VEIEDmhZVVuUzGmAH1ne6sJ5YkNKJ2n7sGjoii
kAP8763GkmkAbW1d5TdvA9TbKFqt1aaBOmi5Ke1StlhOooWL2NyX4FvKpI5q
LmV0kJ4p2ECXJKTEoUTn9GxdC+bRmrMyX1RHjxMr21Asz6S+Crwg1pXkbTFj
ws9/AilzG5KdXIDcTE6QzD9d32XQc7tWbUzT6ye9iIu3aovVq1kHLJez88wZ
9ewqXcrPWb9JHRbS6ejExS0rsV5YvCPdPmnUPjARefRWgtSCXCawOalIvEXy
n7CYngl8OSShC00P7chLf+MoXsG9JWy+T6d/zzTMYOypzB794WyPBHfVFuZG
T6qAcUWDBB6IwRYPPB4SYmkProRctSeQGuPt2kKzJxbOGgd+phosg9ADkCH+
63YAIB/K29yhoU2YhMX/qSZ7Q4sc5XWKKUrLF7jksL+1RwXjvNbxWRXSp1R3
lRwFVuGT/buS5OPTp0r1d8xrYDP3UBR/IIIosXHD31SEudHE3B4yhvrgFbu9
OHenfMX9z4jfbE+LB4W/jP8RJBLEyxUXEg6zE5xhDV1VJqBQo3VB+3CBKcDH
LsMcgeIPphBV2xMWf9ulqsG5aga/LYY/3opGrsHfOVgO7MGzm+OsPzb+eIfW
hQEDbaAydJj50EZaLuzoyZiS7QIpVeWX0s215hSxNsQMNi16YD6DtunDEmjm
n33PJkBTkBdT9Gywjli0ZQAtP9xL0PEt3jVLeQ/nzLY4Fdw3iavArac+hJks
nY87TLvOQU1v9Vl4QZg4kEqHvM5/PDoLM++AFAKEL6JtLSYVIPpj1KJQWmwG
Fl43AnRyXrDt3GhGnH0pl6uS+ckBqVjl6Ogun66f+bYpKSA39i/uHoUg2n7G
jLnw8psN/Z0BHh5E7iLTODvYjbuRZsfEzIqUCpQxzRrUwDHoUIo9ZJVP6BEg
zX/3hxil3bwes38MA/J1iXNH996KyLrptICWpwi9beMPFluv6TB5dtRLbpNe
kCXHGk9ch769ULzJyTzPxGGRKge/XRxN+k5fZDz2ci1W2wrFrMnhCE+u9mN/
th2qiq01DRmREPTaGDRzK15Hx3SPYlWKqQVtFEUANmf0o+Fs7+w25/+cxfUe
t0Vl46aUNjSqqey5z0K8tXsffpUS/so/rwiaoywqojxiYk+JhpGZ2gMKGS4M
kMZXJ/J87gw9MJxo0uEfUJaQ0pEunx8PJjZIuTBSDmxrAzLVffkrqVXoxD46
7Ly92cTpy6Ov5tVnK2e1iY2klX6L5CvTjT6bZAAVZ2MPRMZd9UZcCD7ikqEW
ewIkSGyV83B8q7Mw8Z8nBloy9bxr4hNIqYR4fYHbFwLCKq9fqtguj5ci19zd
nFO4c6TqVE9il9SAKL1MHOUcxUit6zeHsArmkTfM7zLCsDTvR+uCc9rdOQ5a
uBrcVVaucDgE8sPir+PC8WcDiC/KnGILq1GORhFIwj988j0tu2TFKHsNlpfw
xQNBeOkQQR3Gd2U+xBZn8V8I4rAnQMdanwWy2GJlPTPjk9IBb1mehK+F2caW
vHOugL4KqfbSOVo7GvHW0kCmKshNlREy7XMKpEFDDVIuiMFMDzCgxIEhSmLa
ClHDjzWzUNM9ojcY9CtxWYKJcIhktMSx9eTq9rNt2okziPjUzw7ZYKwVJcQZ
j5q1yIMDkuQ9r02jS7ahmaPol8Egz6KrWsXA9M2XaV//W2ckk8GuZGzlr7Rd
VNL+UKF8DJkyux9Rqo4FTRPLKlBfVDASobAA4v+k5Bs8Gj1v12gFhpOJm2BK
LhHw0Bk/gCBl7z/mDvJ+8IYObJ88v5dqCodpEVCWMq/3w9Zda4COPcHP7beb
1aDpDbuQ9JQRbvE3E6UkRVUm3IhWJg99i245lYqc/plM0iN2v/B6QFhxfsV0
tWHTHVnR1ZLyLKNg7vL9qTqxKDXHtUvTf7ZWpQZKzZBBbMr7JLg0p51FEIb/
vGv9miGlg7pTOhkImqLhsesBdu3AQUZsIElim7m2+J0JGindQV/Q0r8BZ84Z
zTXMLcvFSnfv/AOOm1ZEpLyjDGuri42lPK3nN/jnRHBJDwZeN3jeP5OzBGlF
EwWyAzm7xQrqRKIvdyDIVyNs+qNt0mXMrYHwJ3kFMXMStzkiPh7JyQx2fUpq
HidSlXrwuP4O/h31wqlbXrZtn3dSUmwhYBTn3YsMIIgdr7HAZ/aN+K2aB0iX
MEdIwmNxyaiyLu5gPfM4tMbeRMSeT99oIUILVyqhoJpD4mk4mRYWjz4HOCYM
yxJJ5scEfCPuTiHcjJHTvbMFHrtLng4R/Xe6ZgPMn9pelOY9RaGtUheOZbEi
VM1hlg1NEFf+I4csNz9o+Y53nvUkct76xaPzSfB3O1apZ0Ur9oRuc3rT/mNZ
Q2lrpP2KSgQ8KkfDMOMeV6NQdQD3dCKkdequeJpfOvP/PVd1frDjLidAvoKa
k50iqcvQr03smShW+kU6paOnaVxRlgVTQ7OIzLWinTz7l0ICpmLo30pdRGTp
paf6s/VQS9ooLtwCYh3saGDX5CHquR0bl+uIXcE/xzTsj25+JTQHJXJ26dR0
W61kf0l/f8i7y9gVp4nwHIqGLDaR8TbiSChc1elxNa0Lv8laDglMVZUnanCR
gsTziD/qqCNbZn3rdHTbde3ygwGX88McqmP46WlLy8PTs2OIojcFzWlVCyan
EdIFsFGAKFhk3DPAn+g8fq6P+jccDFv8ojWPpsj2UeRSgC6MbiRRcLZLuIwN
hot+a36t2SVy+D8g0ZYKW6+YOIawMcpgsb1oHvEf6WftmoKIhLwsFEGFLpe9
0XuoEZh2XbaIgU05evxgyvshhOx6akdXyFIWM4cc6HkIp/to4299Uu/6u3ck
WFKpteoj9VXfpqjS+xAq52RZxgX666oVGkp4hJC0JrHTWYReFHZ018RutIzk
+ofJYuKQ/6mHEUeoH4S7S1b8TLGK9EgurgGOlL/xQuk+EOsFKuZsKJOAq20X
ZQNrMTHegACuUhNFYWlQzsda11atyZXn8txAyPboF4jTJzprYfR/xDBeqK/5
SX8qPYDLqWUF7HEEVM3245RcIMoSPh10Tin5lNqcvYh84AL/00aiEmkV7m4R
S3PvjgCANsI+E6mUOLsWt9ioMypzGN3rMI5Q8adklhycEu8SYI5cbhK/m2Iv
HkuQLEU3A/sl2uTPVUGaPnpIfVJYAda/Y+OtYM/aLCgD9LSZrr6jJkmLkM1F
HrZsmNR5G04DspHe1CQPxrIA9l4+HEjGpOmicsCPiiOUpswF0VEIwettDQuf
lKzDeAaXOOku4TUrRDOcKPfKcKpYlB8yt1KkvEELtl1uJht5wcNdlYmdOfSQ
lxw5zmEbX7gmwbT44sbk4EA4/F7tBY/0Y8xI2nUJB3QJzs1GHYKJ66JP0PDB
o9QPG4lC56YDA5UkohcsLJlv+ryVkKFiMVchYxCH6QyVhWGSJ03tL9k/Qqd3
5PPYnHruQWiyhVnSkKx7mT4KkiWElAHrKb5BlbfvHeMf55mwa80pjkn8zsz8
SnE2JYlIoyecZt4v9V+43qmpt4mReBcQYeMtf249sDchMIIcaKE/tKfEPunh
NmB2aewATNZnPnncAyQKRUHfcHwxINN5dZS1+vktP8xGbuLhc7FYWvLiiyzS
UvzGMcNFDMdjzEcDYU2U+ZjiCIVezJQA7F58UnbzlqwHqhiGjGVYvW6xYF7y
5l0d1OGoHpYnBf99Vel5vjehOpEy/7VrGGMnQHfI7s4GdyP97iuB7E5Fq/h7
jqhXLZfYtDqbVWMgmItX6IczTBO5pKryk60UyfsXZOjf72hG56kjSj3Xqj+F
t7tf4JlUp1qlpGXHk/3bsMvN1QQ/Sl6VhltbdoT7c44VtfUx0yqDM/0eNbvD
MuGeL8rU4Em7XjZaeiLeezyKFjd8NMsaWmK7GTLUPIV7hj5Ga5CzwgmTaFqh
kLrmnQm9NkUkv0P1bppIlREPJfI2Lp697CC4x4bEONb/QY4+2yypUJxjvFyY
PddHtqvgVnN2r2ALlZa4ySnMWfaw8GCtFN82g7p0zZ/wsAHLGVeIYfzqbjH1
Bsri7JNC4fI/U2kDINok5Sf6KHDmylG0wmtLcBKqX9B/ZLH/j8qGIFZ8pnAC
ar5YzLhiomaQeH62cfeBRX1tKmLMgrnqdRgirXl0RV1J0wA/TvuydhFK9jWo
G8xfxn+hH+sa/bUtOJqaPPe1s++pB5ZqIHEWad9lOrF4f9ncCeAhYD/JE09o
Da9xOoNyioa5YFk+b/UVYrliC+3oWrUxTUeqUVGI+fDBPXTEWBwSXzNeU6aP
YCx08CjhjLgTt4sC8876TONLCnYWnL/J9kSG0QhWAFShYFOCP2eL1RKjMPcu
HCRaHgMZL8eS6QW46pEVFDvCRdQCCe4jjDUufB3DJwIDyDaKWL/6FqiYWqqp
WEq08e6NJJRo4Y4+7IdEo6/A4M5HVMWn0oCEs+ju0ZMs/TBfJSwsnQt/QVzZ
iovYXefmYnnaM4neUE342kJnU8BUqUr/bBr9JP/e5upXAm0y5XDd+OckS2Cr
cJqOs7kuTTUfXRpAVdoTS6CphS056og35Vj1Se52QDAj5rDJQFq2Y1Q6Itka
gD7P/hmWXYGXXeOhlOYAhgNCsICH8uALoDqWAov4rkCdBrFMoJZppWF6G4Ot
D7bpjhTm4NjnTR7Zc6D8qmrjeydroHT3rFLE1DggWcr+V3fDyugLEk2ikJAr
QJWmTRLa8djG+qPRqRuGDimtwQKWqAW9b0Rr0F1phC0mM5+HQod685PmgMb8
YYk6NgEFjHQNMnInWvNxWgTSD0rRVXkG0JpNAXKop1WbWrw/61eaVDT6wYtS
awmRW5IaUGBtd0NkOxBTD70hbYQDsWbqub/006h9a+7kD5FysFW+HrBQEoiM
3L6kJDK61i295wRFqemRmZBCDtmq21uKtDztM9kO1yGWOF6ztvIUZSiMg3Jq
+u7R4AmdS5R0iJa1xfpZYRS3F6DLKswSue1oZ9XRFqg0U96pj5vUvuw6tgZ5
IeqRgJc2kU2/GRy9L4CNzEKtMdbXHPB2lXHGDk31GhNhqvA2gjm8fxioN4ph
1y35GuQbQr19hgpOWdsjQJg370vHtk94146UZgN+oUnAJDKVVcG7qA+0VqK4
roO4jfoeRKd9xk02wC+Qh98+hqiSDc2CmNC18vDRrLIi8WC58eEpnGIFc4+x
iKlCxqJ8enctvCnAanFaYwXeblVR+nxhLoI2gD7gXBv+Z04/mtgnFQvbsykj
hi3zD8ffnNlm+krCL7fCUXtEGVjHtjQtS7zGhYJSSm8gzRIo80BX8taLjGV0
D38MRNmNsQGhl9Ih2jxmlWWN8J5tYbx3c9jSWyChaImomu4+HbeGBu3bExkE
ExFj6obV7RD/TGkZDcv/acEMnj5PxuBX4lu4HLgmthu60P4BsHshj1jv5EJm
XA3lFGnOgjLBnOMRY0y3OD6/iiUE2q9HebbtM7UyYTres10s8/MId0vtMkUk
2E2kRuZ190ZNn0M64+GwolqtdkZ44Tv+NgOESlqY/k/tRC77nyhE9EZWRT4w
V5pcuyc4uBZ1ps+PSI6ZxHNOrPHAIirUvhW8yE2VNV5Kr4pf4vBniGqn2VZv
VitMhmYqS8kW47NK7aC26d8hsOAb5PvLzxuKqUPpNapresYEt7bfD7RC72Rc
surLqrKgdfA/TZ7WUttlSBD/FVcir3Goo29sI0PV20anbiRd/tO7pj04H+Fh
cmFmMoCz5onZ40dA923uw05Finp/ID1FWczlcdoPlyjHOt+lUy0Nz8cJlUnm
3V9YzqLqM/oMN5BSmk2sO/CQLVLiteQGmYjwOMuTB327AnzZAc6PDC1CX27o
iUymyk3Yxd3lAc+V608yQOxyDr13Lzo/98GPLEElZLoNSe0mIJrzCuvL1zhu
/xXQZxYojVyrkt55mPRyPK1dlvzGzvNKxok6RwfxGYIM4xSwhihxhetnuEU1
xUt/35nQxgPM1WoegSPJzXv3rFeT/5p9TT4oaaQkmEMAO+WurVcFlVtBwSS2
oOPz4879w9NSSqPIg2Xb4Kl2FM1w8UevBAbXhZZdkHohv8Uv2hZjuAJYmE8R
HmOzHqEVcZ3R4fp1h77K/AWC2Nmhkab9LSMyO59iJYN/9N4G/xlwUJDo045t
oPhYW0A1aqdpSiM2+aJXjJo4os9qSFklbhw/5rpanlFLf5wJoWaFw8+pOIDz
uCfsYAKaWt/ZvzSJOhIwqfGo6zswTSalNx6tE0+06kbyWbjuq0qu976sanu2
U4BXRmLM5R5PEtz3u/uPibZbVVVAD3yoTCx0HHqVEi8ISIvmOHrq7KHjkSEI
WCnx69tujLWfWZPB48pLrGgNwkbk7OcQ0FqdexDSds68blJFA+I4ofvc6Kan
SrL6QELy2OBK5TD7VWFNYFDRNwGvQrnQHnh5V6HxBYdmXRYyAd7Xq8yLunkr
bRvh9pE8lJLzBmtPEG5769wJ3igv4Zg/iS9l16rtgEFgwrgiKgRCTLJiQ7eS
txjB57PmUVfKP+EOMl2HOOpnXGgJbRCUNL1JzEQgiQ5XYDHZifotWBj/ema6
uMy95L0ci/TJmPJXyjK47LabPuqxy7KZvx8FSlTlGwXpBLqFJT5rRE6h0dQ/
c+fpRQMdnPbpLLPFhz7ZhHFLzCpLSKiaotBrkWgN0W9adzPmKBERVcK5oz6c
uAMmSx/Az9A7nObLmLOqkaXzXP+r1p9Aj8r/b3KqCLfszD3q03BytpaO4VSH
clbIzzQ2RVuJSnoxkWk8+/ToguFlutb+LhXaAvwm8TBSyukwk1WmyVDTpmmD
BaPiaB58sMyShHmgxC7OyKuP0+yxxJE13LwNbUsf1B3FX1XZGAiAKIyyzdGg
gJIm2dW/G7gqGIamHS3WAhhU25j3qJG9RvVi5UxJSZcNLq0UCLq+sszStmx3
l7vZPA0wRXLffZLIVOsOoQaeKD3tPfY1ahUkqHQpe7ej7RaKWlCZO2j66QN3
AZdcFnXsGZ3LDQEYKcxXiKy0y8V0EvR4Y7TaKPfIlZ/qUBIysgOo2VQrZh5u
aSief3VEYrVgbk1JIzldFHKoPsgMZB2tWk61u5kptYcf1bvinHqMh3ZQ9+Gj
jIOvzh5z+w8qYP5HoTvHWIg2Z0q8QOmOxhFRdBHZDEzUERUx3qZ+sS2qEmPa
T0NK5xQOrE4mNlFdQF+sCDubnaEc7Pjimzt3CO9BhQiGTJYGsXzg1ERES/V+
D5YkEtr6QtLQ+R7MR38ezStBzZiq8nqwnHwimuD8USdRxb3TF3sxMekaW6OC
bE6BHAoqgUNWFUz62QT189zwm3GPlduFUjoZZe7a0qyPJaZHHF9TbBeOyujs
M/Zo8zAk82mvcW49mnMsWA1BDpQwk9m+2RQEDJBdVV2z0eBmGcnunxpwcJqQ
wlMI1twx2q2h7OVAf6FkbEtqeHlIYXqx7wuJriDmTBiQ5HAhPb2BUK/d9ywk
cRbvzorOPr3TjlGHoxD1jcwaCPQ2hlWDrQTfnTyKjOojJAnIXiHcH9pnKmEj
PeZQuaSED0jiFGUCaesXfu+x5EGEUb68uZTyr5VL690TlL+p80SIIuM2sq3L
g3eOcwCXGrQPLi/78WJUqbAX0GL192LfcjoHqIQAvzN6AkesHDqfPxLLtuh4
Jp3JZLNlddZuznU9m9rOqDuzdN1aoODyqjEs3PntKB/wWMdk1bqCIU4ofe/9
wKF+qW3Hl3W2l0YujbGmbmxb8mh/ConyE+m0n10YcYdfmaLuacmPxg1Lh6Qe
pPft6Gr3J7ayzKzrdX87BK2bkZhQ3v7/Yh629iMbb5ItZWBn9Hx6yLZitWsG
K798KAUV1y5Cv8q5II+pnAAzwttD51k8OMsDIuZFeCp9rxvld2q2DR4NQpB+
TOAmqqo0UWZbz0Ljw7ENMvz6+Xu8gpTU+yGLYz0Z3fnnvap+P0zaMzuLrgpy
5xsVrPpkp3TKlwMRu3rpOIoqOkMmYA2aBZ5SANSW9ux2TZbUdVrGhK2KNq1j
T2PDwtsidWdm52q9sLpiLRDt3R91NReqwn4epSII/tTh+2chE94tcQlDOUmW
k7mpKwrrMO7ZQW3ICJoVhAOnIFO2srCtZLpTdMjC8AyDn++D1rZy85OPJV3/
2pEYKqfgag8cmtojBSRNruAXnkhJN6NpWe86r3vWHP7zqnzijpWYIlqAs6K7
EHirvarAe+/UCNSOQuY/BdG3ED6IJ8OpxRpjGMo3C89299qHD0wO+DsOCtT7
Gc18R2uNLZOBsD8eOzsyltxTG4UgUfZIrdfz11UuQHaU4AXPaje7oDRdpNvB
O1jcIGj9fusl50foimTlrV7LBYGKLHGnCk/uRMJxMGtAbcvqY+QgIG9A339n
ZpRYn/DTTYy3Aa1Q9fpX08w0GZq5xgSBIwpRkG6590ezqYU4R5/PW2buKqXY
bXaeRHyGJ6WxEy1IpXy7Gz6Q5xZzLEW2UQ0jyHvEZxqCDH+nXOUyJHsL0/hk
t38cl7PenjwKwHWu0p4M8vjhJBdgXmSG7+3H7D8sa2+ZV7oIPhuSwnYOPrJR
HwHOHRS/g61mbm2A3MDW9NC6T7QSfGQlk7T0G/jLOj75svO/Ezj+KFs0hqfY
wO7qHP8ey9PsEXcC9MUDdPnEcGxpMHVZrpFAAuPia0keWH1RZWEcn5Gz5V8m
k2FR9Z9z5GCp4FTk1IXCevOnSvNiiTpCtX6caGF8ZW8gsu6eRFJpfLjUL5fH
dSIGttvUeXxmAfG4Vyc8sIsWDv4ChzF62DlragAtH351ivQVS/CZi3KIsqIT
7FWR7b4uOdbv7jrDPk1+NH6ybTxujCyDBZlz3gkVqxKJP7bO/y8WLXIe1h10
qwgpqupgSZeeKIPCUuocbRVMsyp0l4ZUMMcSEoOoe1N1ID3KyErR/q4xgh1k
INGCo+C8S2vPLlFUptCf1CVELxo5yfoaY1iOGBGOIW8+UAlO7mvmyE2t99DQ
WCGOa+RXOY+GClrTrtt+6JtqyUDJvLenHLHvBm2kNzj2uiRmvQjzNs5dWcTJ
w8J4T7nSE0Xum6wFwLvmjH6IP0kUqHXyP7oXo0MHkatTnkkC7zQzkd5sXut4
aqKuzbgeafzaRuOl/HrdgcOHNW/NSViz2bT0Y7H0n0vcnzEFcp/bc8Nws7ZN
CzqPcHWT/cwz8UNYOKp9Gf7pOhR5azlwJ2p4vHULHxIdGujF0FTnWTMiWnae
Pppn6e3/LZn3uuArz1bYr3HWUtl6JiX+0mXKYBm1mU05rxwayWrRYvd0255n
VV7MTFSWzzmNieIyE1QZyvbz6nNJe1L29ae9HHHiLdzImYYXJUFGdvr7/gK1
XY4Kq1Qd6yEAJ6VgvsuagOWls5KL0B2e8X2TkNdRFc38fTCd+scjC88nRix1
cQNDgm0eZk7/pK0mkgbaseUkqN2LvF9QGMaMQo+6bRwtRRNkEc6mmd6uHBVZ
fdQ1PWprc2A9vukAUDDpBgo2d/6jgD0AMEdEvRW+YRyfOJnlNS8FHMkFMG9d
rdvVEvjZ93NsFRal0KodQbGr4z22gOs7H14Bfl5B32ncy6A/SfrRjTenfquB
dE+JTQwvLEQksxFgWYilBY98UdqVdwIxGbDW60nCUQEZi/Ua+BhhnaUkW8ii
rX8tCZAwH7h+cOVh+gFvVzJhAgsM+dXSLxK2JrfBWOdg+JyDc7s2rqg77Bns
NtH+/3i8vBxmrbduA3R1Bjp5a6fLnjcDTxSBge/5yRmFAtto4ZwC+AE9zxef
pZAXIIX4mABfnGrY2sJHCvFJ904tD+rN6TcvgCy+gHl7br9+uLoqWv62mDnL
+jfn8z+UZM0uSLZKvTvRl/eO6L0XBLNSPpLMKEUHUCrixlxFKVTbqdN2Y8eq
JyqdsyzozSyUdz5MzsW0ZRlT1U8IB/4yGJ7rQyM9werO6kY5HrpccvzVNywB
kjcWXuUXmrvRYJlBWYQvwPgdxT/Xkm8uTLM1OuVmiZBF1oY23EEYYlpJogN8
fItPEzpguqoK3JNWy5xaLJEZCbKLmrs1kpQfFbNbesu7moM62vSk1kIKCRVz
7PmjhhdROyK4lQZa1Vg77OVrs7WtnuszB0F7J4x61udSgyioC5kS21EeWiI5
Aah3HfqS3Q/lohVVUp0k+RREEZ8uAInxXjui2VV6jqdEh4XC4TTESdbAf2St
+hTXF75gJsQPdZ5TDOkJ+DQRYFte2EQdmPjvGUlRiyhTdqFyfOr8pLsEiTYL
EBI+aepxV/zXm5++xEIZh1u47ijdOSwDaA80AbeNe2BmErj6nRDddMXjxyVa
kNH0l2n5x8fhRCkRITkvflB4Hmdk4V5lQB/ziVHnpZ6GPvr2OArqIjxCpSxO
TZjYkjw/xW6Cfw0jdhszjiOkv1fVeiDXLNDXLfz5C2G7yaQEJEk5so6tVpJA
d4ksBr443N7SQImFfFHUvXJMn0kOr/8PtXOIC454hOARq2fcC9l2K5gNkLny
KmvuwVibm2MYEGet55DHDv7YfCP9NYz50wu1Kr3I5zUJPGGz2/X03Eq2+YUV
s5ZiTdqxySmETdqJkzJXgm/LhpNH9+EhZagoButoCoXp9U1Vg7HVbsOesdUW
Wjv2qGKK3rxYuQ2mKoo2YsR+LU38Kl8/wN6OfnsOp1doVLPpLwefaMVUo7lf
+o+H7u6BWFM/51tdPz7KNIImR5aKD7CHbAp6ORTM8D3xkM4CwWNHd8+98Ax1
HbM/+vt8lmKqVHz6fqX3SR09Tnxol1G+yQ23LNTLcq48dm6Wd+b2yt3biguQ
aEJcZW5OpqCMnKTkvrXihH5m+HmSn4lEFF1k5s6rBJonpDJSRraNnnIaU89h
01VwpEnrqW9EAKW+5Wcwso4mQGDCGYoXveq8OBxhjnPHw/eaH56N5tVA3/6K
49NKVuxebN46Xg7ICfnl3ikJvOtdhUee3aSN/cEp0bT4+k+9Cw69yMs2oZjv
/bt+Y/sXGl6fiOYeAL1VjyLFOTWNICbr3XSpeaUzgO9dXUoL/6RhaIyFdFkr
7/dH7tXVdemlGXtsYtbCYU2MDO1XVNSVBTEGs/iS88SVjyABoysuHdQ7xj7t
Iw8ji5FyXlJ1Lz2Y4PAURiH2s7A/aDKbmtEqpJVndZ3mX4Lxob0UAglTkXD0
/kcavyu8A0mxZbgS8hN89/0QzfSn5HOlGm77eoaCZ1KAiZv6/4sjGhfGfcee
CNyLJneO1oZijtU2S0xpcF+oxwGlYP3Ib6G9Rk5fvWZbv0igqK4GhTkNrKsZ
NgaLu6U8Je3jRh8Phh7vtD60/9L2smUsNKTGvJs9EMrDQcXtrjTEWPMdhXFn
yk+kDIIj2XHrsZHMBj6mF5kUeGJ6dv6m6G5LmX6+Kg/ven+ARFA2WjTj6oyE
gxAdRMeli7Nyjm/gjhIjMTsbVIIQFIgwVIzLhFRKul47DLArxT0pRDVrFYLm
Xc7bU+S13mchnhLDneP1u7kksdtBtxuEVO1XgIcg/4t1F1Qv0RDOghJWjiwp
+6OC6a8kU3Jer5LBR3cdfPw2RYilG7RUWj94G/yNDzkuGZ05I3MMAIB8Odo2
jS02SVeW2Ix6AJ6j/kgUlqZ5s1pGjXQgdznLp7DIWSLAI9NBk0/zjvA5lVZY
F9MOBHUPwopLVslKhd/jMbrNd+Jk7yPIO16FItKy2p4hbUQLwXAGvU0WqoQo
QLLHu74jknVlDs9ZHCYoLGc+0aqNFTn9ZVueW6hRuMdoMTWG1/hDL4KnAMvl
WYbW7wsqlVsAswIlbKiCqX/0gJnf/Uxl9ROrVkOTj1NsTSZgD2ARKGYGsCC1
W9pz39txd1zEMv40aX5XNLGnGs4c5s+7jPwwPmAOCbJ18Vj2vHa4afrfX+Lu
RFbIq1vhTAm38o/ED8xPwFNHjtG2hZHZHils1+zv8cF1Ge1911Q/Sc4baUhF
Qj0BJKX1XCZKaXiimxHUW2PAUIAfn8KnZ10pwUMmUFR7oOThFdr+55zh7kcw
nhnDqb744Ls4R5evlIuZ2nc7iSB7hk9QTkvAQUAer6aOcQ89qzlsrlu1oZJ7
mcMlIVDZ+OYWDHwWPFarFb5M+pZxbKb2uaM9gHsjs1m+RmRNbdk3MvfrxHN6
Z57YxQvZ/N+wjwt+1GVeii/14ataGM37iIXnd9qqW83GoTPQiIcT5e9vZ5fe
9mPCMVf30ShEz7GQTKnwtnsXnpHJdZGd+EZ+WLxlzpMQHnjDIl5bDix36/lg
t+MqRmWldKUjTWkJrV1ncsjRwCupn6s136P6NbgBALW5jhLFQHJaaJKDZU6d
1D4tgLwVzQRJOkzsGIHnY+AWSaO4tVwx/CM9p2dPCNE+VbGW2NZrDEkeYoiD
Bn/sTg5LKFqDh9Pbv+aCHVQJHWIgu2JkUD9st9oVsDVPXP/oYeLYJo5J15o7
DtRFRJvCrOLUKf+7gfj7/r1ozGqLfyA5WY5STas2zdNAlAeCifOvbtlKAx6N
sznLvyw2o86UfT8BtcjXB8CDqouAVKiA1/j28PrA2ziy81wCprTRpZGPP7l6
e/3eTzFihpW0hsDidNKFatiYfrYOGC73yvSTkIwdp+zsB+XIQS2mwDjH429n
I73r46nEvUWn7ytBVT8iI3ZpMVPjDv9IFQYmW0/dOkH3YZuODkNxWjlhFlxq
WXYxhfnfZyv76/OWClxmIgMog0jCsDCuSpAdmRrHvALosWzfOi3HRsiIeryo
QmqPVSPSUCDg6wPOQqEelWe9m7m0M09RlDfbggX7BoK08sG+Lw/hmjMZRrXr
hktftKzAk2aXtrfDdQUWIQ0X1rJhSrnnbgaGP/UfImQW5kD8t5m6bS3YfVie
0xqWqymsABUO+VPicOFGdnkM+Xf1H+/DwOY3CxY6u1ssT57h1crKs+A6dMV2
fXjvUSR0jb/S1OFaEUh1vTY77m1BkKxNLG39soJZEU5yGdgc9F0e3DZkvhs4
yPHRuDD0iMvG5IC3G3oCUCp6BqmsiJB7/+BDEyWK6A8YcIZ7qjQkhvL9N4he
ziWWtNU+4/KLzPMVcKu0htYpSl9/JL++2jeSvXolLCtLq/vfgLdEf0roU/Sb
+VyLNQjVLtZX4QV7r/YDMOhL5fYiV4ZLgea9DwSKW68qYxa4VcoJlUiWaebl
e0ia3ltCz8DeWAEL4aySuZYBUsz871ak+dtnIzZyWQbL/A76oYbE23piOHQ4
ybukxeGndEH08oWS7Ftydh5QpOsZkEbu9w8dmMGfaJCHhfvNvlUxUm1TJtPe
pKosjEeAviZ3W4dkANmUvc/PYHL3GpmhtD7ackNSjdsLOI/YIdqbPApNgP9J
J0XBHSUTvAzCEDCpWIp7XNJZU4CbfTXICUjKdCjHtT2TEcG74M53fKXpaKPl
MPNmnWU3lc+S++W/HCo0ZiPkU2Yo0TG12vaVqgWXWptcUwSl5qyeBbv+QeEu
c0fL0mqFgQljF+e0qIKbynfhfamudW7YFaWERD+yLmbB8Xy+LXE0kS/HwJaO
ob/YAkxjHhaFPJ+VWMi40neMip1PzVcCQE7/AGXeJaa+31hrsB4JFQ4Z+Ic4
iVw/iU9213svKUrdMKC95IVwDsezSUB+wOnthBms83xEHlXSly9nMHYVMEcN
3ON0cYCszWKsfdVPjMmWubuJsPzrl1HrG7QY2x284l6mBIBZ/sZ0cd51g6fo
x2pWpDqGAvsSMuP4Meyki3OTeANtHciVPk9vy1OXObBgOwNRF+sP+s4j+VYg
YKcLr5giysCIpF3fW26Pj1tCxr+i6s51obNeIXf0W4wLgTNG2fO0khzqaTCs
YwKqupzeeOcz0xTD7IQbUqaoKI4jplImZqaumn5VB7oX6fqTp5349nTE6o0n
bDEMik5pxFPTtR93YGMMb8QmRnzt7jj/nyV9sAVtkO3olOSXXdWrFtnlLT9n
NsP8AkGZIBeF0Cx0LBW2vHcwzZMDGKf/KWmVw5B8YbrqllqLX8Vf6wVk4cee
IsZzPtVSH8aHNQ4Yz3jJJBotMr90ggKP5bvubpM7eJGWVknHgUmuJSSDVfV0
aRjimi5DMWt3zrIscjx/kyzrOAxMXwd+NKXU7DsB0+J/cgi7IaL97TVbtVi+
QMMoPzcdXzekDY4oNnbdA9Grj/I6vWRTsVtDaoTX9rTVX5tOI3ROt/l19bnp
V8qqACkmjT7Acs0YaY64Bz5o6/eVEsGXvnvx2xxaFtjBXAAliYuAC5K+vUhz
R94OtnkMcx9DJd5NfQ/pRW2ZaC/LYvw8i05YYgahgj4W3t141dgOfU/WzdjU
mwTtnvLW2XIGshb2Qg7qjYgrEPTVEbt1R9OsSgxBRHoupC9HR8NXdc3o//Gr
bDs5nFto0loMyqKIZLkUwazmSYebXuCRYKCZ1bOyUJ9+sDn96MxtXhSgoPJx
mZYrdh5vLJ7lBs1rZN6LvNnraeLl0VAa16OCO46JrhSN+kRRjaYfYFSLpFyr
1KcU9PjSO7t2O6/Ql3IAVU0kJ75AQo9VQie6OToPQeaQn5P/qvvWD7ZFwwNl
Z91nb2bAIRjqReqyoU4GXOSjge3famTuejn//YF4aVObqt7mxGbVL/9kd/Es
q8l3jc+VZNnWHsvnUSZU1/V9DI/4/xZUnVlT8RYXtbu/TmaK5WmyP9UQ/mtw
y4LmsslJv2YEhK+Qf4rT3DkoZLgjwo/ihOmuQw1fH2Bl0CZnq12ynRjqNSoc
dDwjF2l7ElgURMT1YjD+Zqqk89VHYcEjzf+zPDNtpyB2f4KbjXZgkOKEcx1J
+8/9VlZ5ZhjTAilJuNu78BBDRD37Rd29cBRV6Wt7GkigfV5r9rBmB56eH1WJ
HWR4UI2KIp32l6dCkiFz8f2V2TcdJPmj0tfZhYbqYNMLZ7WJ4d8FoU6orZCS
Eo45kZvZttX1c6rPUitgFpHAJJNtB6bWtImyDkqRgdsCHUG0Wq/a4oXeQwWs
LRa2JmxLwYI/AwcNDqA/VlU7RoAENqyQ7V9szkKcaz4rVfLenA2TzGYsuad+
Bv7IWl8wmKjAejTTnQAFZ9x0z7EsrEP0yUK3Emcdtjd1y5oVpnjKCxvT1mdK
+djSD9mmNx+tjHKxU4/otiQpeLbTRS3fEuCB+xr8mqJCYpdPM8qBhDDxWZOJ
kuFUGWz0ryGiJ1pW0dpdv1nIUdNDdnKaYnQMSjCYNzncPmqqcLZVJNiDXvqY
4kSDYwSIXbXaLxLxgyBCiUwxhMmE18bJxs+r2ZOkGbOnPMFnhkCoKblv0Htn
RUp1YMgvBjIfHjF6HbGrC0QQM6/550nhuI0ZRP+yOM4E7NuW8CtzGKG+jH7Q
XvVaI0kZAnTbTy2glLxGGfIoRhFa82lUIHyR3bRsXh1QLYskAfjGvey3/U5B
Eav4/zH+YP7TFWG04Z4FTYu6pe/bLlZQo1NiuidKrWmNqmT6pHH740nyOJlE
kcnbIv7EHT1iq8MJkFcNdtkR0deFRk6TJwXsPUrO140++mOC2O+SPbyv5kN6
0MH26WIH/CKLpYcJqNiyPwEXEfTdHVMWghY2GGcIARuL5lrMziYIaJsuQ69W
r6El/WeL4H0CrVn3s3eBOM4emheVDdAtec6b1wigE3/mMwl80v/QPQR+h1Sn
HdRCoYEXB7ivs+Y7PxHCu/iQmyksp7lVyBHJGtqvCK/CUJxNLFGsH1yhYRcE
/d2EqhMuHe868jObSQIMNBwrqCbRHTH0Vel9nPS/LgQhsU5RxRbJOQ3GvnBt
VJ4XbcOliNOJ2aKuV3zLLdIm/xTaIVfYXN5M+hkKi07OJ2P4r/8CxXK/ZItu
IHvdkjCIhLfaepBWg8lKO+/s+nZqEwURkLrp9MR5vMuUMQb7+w3+8jMIJb+b
4VhKxOPYrz3HOdN9UKHLy0ekb/7DItc78abI6YwxG7Y/zhCtvo/fHMHaStT2
G2w8B7pXgBFtpKH5PZVeJjfVaIC2uOMxiMCTCDZPuMHAnLXnUV/X6S3YNsRH
2LcAfK4LhDWe/c8sSnYtFWmRv+ORkJSfN67uG4kCRQkgGwUxTJIMDZRIxGvj
UNYEHdhqTtQ+RWd9JwkL9eqLQQNT3ZLaN0qjRCrBl/tI27NA34hJa0DOVnQh
Tbwcu6iwqAlZ6pmlxyw8xA5Uuf7OHCmfd4Ec/LfFGvLJRsw5OkuvC0HHrKip
luaiuHpAZGQflayPIvsaI+i8RqO2yb0WYQ+/rWPULG8JmCs8DpFDtFuOwhHo
dOEMg1S9ziCVjLltEz4jj8jni808CS0MGgcDlXBYQ+aOhLSQQO0DP0wst0px
gR3i06CHPdzq0zwOCkAR0D0GgyG8Et72j+/23kBwmb34+XwDtkA+pE/F9Rcn
drFHv8zq8V8EGrf+8AZVzAywBiPn4Gd8276DQvcBpvwJXwqJyRsMqINFMAB3
eVgklNUqMhkTPmb2r8e2AgAXCMFFljLCEJRHe5CMfu/2gZHBdz0EzvHG1XUW
W0wrGGMPvAiFVkrCzPffW+T5sMEbQjU46O4XsgREWWNJciUDkMJGlr+LIXmp
83cl2co2W8xqGQuOZX38KGQTeOKfn3bB5tNIrw2yhBihudBba7H2BOO+1PdW
T++ANJB5NqXlha1jvIKfFjgBL0RzdLwMycOz6nKrxSwsSL5UeEcPLpQUcoj5
oGuWO1rKApid+BgHgog7NSxwSAqoEPPPXOChkG7nmRVrVK3p2iXwHfchk22m
/K4cGHcdaLE9hGf9WZZhsgWcY5le4FO/ndKlq6O1cnfUoHRh0rzXGBkQ3Hu2
rDL3nPMH3GrxuIRTzcvKsJcnV/7Q4jAx/iumi+sEqI3oa9QEt1AAilkgtFU5
JA7DMBP5uZY8tNotSzf9FHuDZvRHs7OPypvF5I4nKnXtqi3kXgwLvQ/1tcmK
6fAgESDepZUGzx0rFbXDQKDPFxkLiGzopQddv1EsDyGzzZwTMRwy9Ptn5pWI
065sYdW8bWJkJ7zqHZUk6rpSa0UQ5BNpVK5sToqRHMd2TKrDn5luvGPKKnHK
e0wBrrBPI/ZnwmGjLqQNv8JKYOn/7fSN49MYPjhkNKLC8IEEyIQU8F9XzMYk
DwIylE48LWHLUeKTcEA6g9sMOyYdtOtBI/4a8dUTBEd9uu/fGTFiUOq8uJnk
1SlpXCn5i2M7A4+wCfa0kOXB5GkRmEIftLqnHCWwZqBj5AbbZuob2zfmbymT
I2WXcqRBnlAKB2aH5LMDVPstb7nuMGF6EZoikz1u/17VlDnwuopbwwcUlpX5
Ezf6NnMYLKwpX/d6leI6iRNYa+oLFMLEn7klnmba7STtG91zo54qQKOPASHP
/+1bkP2lEx/mQHCiHdP6FisDwX6+5hxX2K+YtgMvbyK+ARSy/ReHA+8rxDz4
mwOxx4+M7r3xnvEQm5WP5GCY1m/aEyPYODunsyx5cVkN9va/akPBigt3/AS+
TpeSdRZ62KrPTqHKRTVKxQoLV8Ni+r7QMQK+oX4v4UTOOgp1NAUf9XMzc7Uo
iIbdj6SQKbGwC/4QGchmVWT5QmELTQMg5kigd2+lfsx6qbo4HJOVXtaF02H6
y70ylziL7Yirc27ITtFjGyTY7gnXIaEgaeLCubLHkKSWiGTpPVzkqXoexLhm
pGSdqVPn6WBXqDcsM0NmVtYCZrsGHci6UzBsGes/GCTPU/cUFo5Ru9b2OwZ1
FqEhuAOKrKr/wOKwwYOQ9tzerfsGivNXtZPELt40+z0VPO7H9bwd8QdTcif6
QCsCqEA/MbRj1IDeH2W/9wAC9W/CfX1Qr4nQstB8pujsusiB5E+UqDFgkcYC
8ySJ7D6uFVG5mZ+2lTtei4xg9anVnjStHB3OsiRK5XLDHJVK2qWUPd6lNmsC
PZnRVRokgzNsm13uaZGTxS3j6h3YZnEb0XdE3/2wUbG91ZJ8IuliHD9uviII
HvFYv15vWdblEmuETqMslI9OXm7KxgpR+oblh6sAip1vt0tQPNt6wAjRRhAl
oMGoyFDXeZDnzLS8+3W+b0d7A7jbq6m+LHTMHa8kYrR8WqAafq71yj6ZhfO9
z+W/a1BEJUC8+npFZ8Bsi+n4O8lKdRSlIl0WeIuxN+dH/g27yWdeEcPZiW72
CFO5FoIYbKA/BetNJ++oDuKVzLNP/S9IrHlnC57YRRfjvgIQqrkTw6h1KShs
gxOSZV6IMdMAqCCtQhmOJ3WKd1CVHQvJtO5vYart4Zc2CF/NQSAOQr+NTpE5
HPwZ5qpZME8wNYy5ccIWv/vXs+2XYqonJif9AfoIzC3MKFHiRHf9XwjczKUG
45HxEzYq5BikYBrad4Hzt/lQPjAERDsGXJCfIKG1LpHWxWuPM/yfOXCZPpaH
jH18ghFDsrh8mIPyM63Ik6PQxaHRxfsSHLd6/h0ET+k2GAR6D87ATBXSAiha
sruthBZAFHxl7JTJMsxy0Mbq76TtKiLasFdPy9vfxMxNQA8etzKaz1cstc7U
HlLXEp9GkznBmD0+yHNBeV/65pe+sNoCn+VgEyXXiJ7vFB/9dKAK/lzMphNr
rzBj2OJ5k5Bl8TWkLe7ts7eFQXhePzkHpS6t4g0wQGMiaDvYb77p0Jwtrwq3
+c3p+DU0SglqM7YSx3BmWITWNKB6MGofO9Z3Aq2+RKn9BKRTFnjP5z82okSP
/eqs3ZijoMFGaftLsqcTvlpII7jBMu7v7qECRSlIVcu6S+E5Ucsh6uA/ByhP
KoXOIq1RHpMijMlMMJJjKYXsTxZmIqZYKbnJkqkKOVbrsgWkbtjns/sk6Fb6
+5LwFhf5vmBWjrJLG1gYHjoCTtNEpO/4qweFHbRKi+nC1eJ4En2M4c+OVBOt
OsQumaXwNjSN3cesb8RWAopTIx8odHQJ8sAbmM5ZWsjqLL7b1txdKi9Ucx+y
Y2tC/AUb6lcoamAcsFN6ipB96J6PfWY9H4fkqCgvPIUfnc47FLuGOE1pKWwP
RhXXnu92AzieSnB4paqcwc9vjALYCZxrt4CIpfshuNevlNdKUx+TkGhMuYmA
JLBsuBYVDeShtMBAjNem/P5/ff08cOzEIOE21w6tpf5+SwWiyFuRGDnqLwoZ
Jtc1e3v96KPCHGttSNn7miilQ1OMA9FSRKTp5xsfIu9kzFsxfhi0SSc8H3U0
oYoZPBYmwvU7M8jG/DOL9bOacAJtM6JNk7AtHzXARPB4q0v6fkASExLyI0+7
iE9edxkWPYjv8Ec5MmYRquZo17yjncwPWd89yv7/L/TUl4QFhiYdF/A61BnK
nR4xcfgnF+vwGCBF8vZkAFsCZrLXugu3pJPyYWs7PuSK+iC3FBlSbggjF7cC
pEUnvjrbp7hpC5F45TvrDHiVTc3qW27lslOUcWdz5z/h1g8f1c3RtjH+ROdr
OWX9a+EAe9Cc4YnlIIeEq3tWN6+F6vDj3xaFtWP2RHmhBwGEbwIJEHxHh1Rc
vBR+OFUREjBuvfJd9mIPjIAAHEIuLPQm7C+BkokV7WrXFjcYTqlaEiY6/Vpg
u5WERzGPZQCtBJPfY7e1YZjyKGXLTKKQsL7K+nGH7kgeXhbCTtRB8mh8vsfT
i/15aBSqoY8BsovL6Q4q7Ga0U6mRlxwjBWS9VFSYJUlsmY9kIupc+HQbzLEO
gRCWFL7WfBP7TS9MGbxKJWfLKQ65Pwq+SfeKlQknheXp04HAdIRzJyy3LANz
AHonBDD08g6tJDNtFrTMjZ4Qg4EDRo/bPCHP8/6ZH9+KRGGA/6GhbcOXYwzm
mFb4LIwCZm8+pNdiKoEmLpmk0xuXv0Wn8YGq3otQFEOyZXYDgZvnTC/x08j+
bGQyYrm4P0N6RlzQIbKovpSh4c+jdCeFXBex31CcVCeRknqZUbm75+CTFaVu
BIVabYeoIy1ztISgsQMFRVBKoggLoxAQC5jBROJpFBVI3oQ02hrNWutNSzXj
Yq/a8VN+u1NIi7PDOn6b5EShz3CQCSy/pXa80gMtFiXc4mpf3VdsMHg7bHQi
kNfjW/9tEx1is3SDWiyMtY71ikECzzlPjkKaSdLS5JUNFNg0JPYgSJZwl834
cBb3K1LLX9/GXtXhdxdFFzyAAdSLHo4vdMiN9AC+aWQCmnDT16yBwnDDtk49
XOqBrnkMLTUPlZletr4b32Gv+aWnT7dZehzHYC4ydYKGg7P4vdKoRBZ/Ug/q
ceO3vrYOmigoji5/iGKtSIu7x2bHgALyOt8pVGnwZRlFX2sJKaf1ADzPfveK
DebHx48bwwVzr/Gj2WLCFjrwSeO29tp0MXaCRqKfcB2VPdJiU5sdwqitaynM
KJqCCBSc8s7KY82EYOErwLAGoyF0gJtkd9Ejd6GvnAQ/eWE2zA9FsYYaRLeG
K4GY8f006BwMr9YgiJFYO2ODFAlETv8Qj5RmjqX6imdNIowL7lif5hI1DwD9
RAhiSsrZb9exxBF+vqSr6PrKfqAey8qD790BQb4S2U4Phao3j+MoQLKnkY1R
D0M+bxKLpF6Dtqh629Dpt6Woo5eiy+CbtbcwZu2+2UQ6JS2KGAiyPovLiA+Y
I52Z/aL+w4qDn1K2oXIp0NNi23EryKR5K9hqtQttz9C3US+Uz68tqljyKpY9
ZsEPHm0e1tc2VumfJs7mfqE9m2V2xrE/yXMgmSFBF4DUQEAuWM7sJ3yVWVDb
/SUg2w89ItboglSwGGgWbA+WRKODU7E9RVmTWjWyDMHj5svv0PD6IDSwuVTm
VzhcDwdGVjhTvi1alojzVXPj+xp64U9PEwVrxFJZuh26YnEg1YI480355leo
D0bwK327vCqkktwaDOtNtrcBwBPI6ffzlIZZPrGT/gmxKy0Sz18QRx4girMH
KCHE77jCMiAZwiTOuViEJLUFpKkESXhKgFVGx+YZzch1OqSstGOCboAO81XU
D1mkCbd2Aad6An9oyfmdzr/Cik4zd0ipKOG/RehxzCVYKa5B2q+OFHpvXDD8
8uO1R+7xv4y56NwSiOmR7dvWFzKp+drEvW9nyiEVPp9a6CWD4UGd73mzfoDM
42MAYiIArmgZ00DG/xqViISWg5OxGHxqJcEU5s1e7hEbaLXgyr3r1OIOlF37
i3P76vwxdFGYb3xIy61IjRvWzkRBm9nsuTq8Lq+xuCJ1SY3sRF2zqF5KF2m5
U3WFfrB7pzgrjerzNAd7NsT2dM1DBD6QVibtohAJ2W0IKRAWIi7mMfig0pWQ
Cgbk5cWwMP5+VnIp4VOitEiO0dIwuKsHIGJby8pH/Xrdx9M6VJkn4RO35spl
fGM29RiGgX/9XX5dClR1Mah6jaeMFdUjEuObNMhKbnNAmyBozgspXw4o8HuO
/d5OhqFGm0FXNhE282E2fKDAtj/6q3Jdr9uPoRrHHaKH7JjV6k8heYsSx2nJ
c0/YKmunYG6Klw2goViWtS9EhlGkrLblHFTXhzH9lX6TLIccqFAISrrr9ElW
ExQbXoPxmshcGbLyBTXPDhaWDenh1Y//T/AaYccYbaJ41mWiWp0EWcBukp2R
bLhCMz1RzAO/VCoYakGG7xkS+oj1miQKZwlTmhrENDdzV16JXbe7yhtQAmfz
y0lMNGWIqTmzu5o9vRQbhqnlPMckBZK0G6P1F9RSPc4syIFVqTus2hQ42tIY
5H6bvwNoni//OdNsBv+qBMW0KoGLQu7jhYn8igL5ULKT5XLjKLzfI4cNoFKw
xVatj+0iTkA3btZtrgIG8v0zRyRtpxuLvEaAZxepdYrIRldZV26zZSv7X/aC
/Ns02/IXE/N3jZHbuK6nkSuyEgadR9tkKGFlFWs52P5KS7DmtQnjraLSS0Lh
L9fAB3qb+VIJkZCrhMNIooRxa+QEXJPc00DQMaDufmTYIkXxOkR57bi0RnKf
PJvkVLIc2urg2JstSHbuIP7H//LLhOjFOWG5sTTgYDMiEfK8dkE7HBNhLB+d
9DXOkvAl3j8/y6avOzBBOhO1OwbVz3rZVKuNAhW8iFplQ5o03HGz45BbxbSS
fFv4djgCwLtOFj+W5aiqDxAZ5OMXgpx8fHqRkPgwI+TsYYpkxRwIxSApe0ZB
0gp3p+oTP9OVUfMUyhAgspjMg8x/75a+lkk45Bt6q/YhIpVTT8SCUcSmAq60
O8v7ooKZ3JCQXzIvgpYKmH7GAEQhQckU5y2hZv9jZWIzGuZV/SFhCPfVabiA
UAuS1KT4o2NQeJeK99mMrPMlDv88v5xTOVQEOAPk20WjjiJfvZvYOjAH09o4
3Ka3wMigw4D2Lxug12mwjy5j/gnxq8Jx2NOqHiy7dSfiXezqmnqZnShJksCR
Pus9QRmrZ0EpjqcSdKR9fZIS4xOMb5f7EBN2QyXzZhfmNH1XPSOMts9arnuV
djGP/Rodb64l7WMas77EUdxGjHy6rV0bbrdvTkyKoYkwHaiS2Ucl5IBfLPHC
37L/C6wx06Yxan4xaTkRLuTOSxIT4pYzn9FdVbIyGT9hIYl6gEu1b9Y9kTbH
c68eWzMWm9lxw3c8TgYzzQxzMa8i0+W7tRdCM+BQ123dSrSP8FXdaf+h6geW
Wax+414Rapo5GxLrdyOeGbDUBB2kXIyOpJ0AnQeSpJz1D9v0kACqG5C9NCy0
stxVe5zFLnmN8/rYOBsQ2HK/xgPBdexAZcy8MJhj3CZoyr/Ws/OxuoQNG+vr
DBBWwHLdYEqw/5ohq7jC7dgTiX9L8OjYF5RVtG1Z0KI6YMmgsEi9RIEmF75u
t73lukvxYX/zPlGHiqHXEYggsGqHKrKAgAF2Jx7u3OtgjbP3AnjDWO2d27X6
a6pKw1H683N9wqGihgIIxcPYgrGNRi/m7OkyqJri5KUCZLrzsO9uIMEGiPla
UMdRWPiOtRmpmoBNGy2QLom2N0ZQzAA31TL175Fosl8PMfmetJUmW5O1p/Uq
FJU18Iga+6y14wXENd4jWoby86nEJes7cV8pE2y0DoO5+MLfANqWc4Yu/EDa
m1WJC/k/+nxgkWRPFxG2kq8tF5c65LNMyLBZUoGC9FTuF67FtzJDcjxpySsX
kbAQGS9WWHl/zN8ywszcZVDaBab8XHypKqK35RBKej22FItZB6CLIMtWlKQF
QR4RN/lpsZEBf3Ej4iEfNoTpz0Xu8zOGXsLNsg6mf6XOD0IjWQ9i5+Mh3JMq
C7w/Op5hG4UJI+fua4UZ4jNdXypSdunaITIfxvevy4M1mTYn6iOLCcgE0tMl
qqH0/JjynoFDABqcYYDjXJeXWi9GQtbF1HXXHfcEnXszceIHMjgt3JdWzR6L
r6QAktB73UtK7WAx5+DKJBdE66nwYqsTb3eXCWLo6xD7PZlg0hL2nvqUlMWc
RV3f30b3EaXYWV5pi49hStWUWLM/dz+v73L1x6/MVyeX9rbQylphr3KK8otl
2ixudvOrQxD5AmPGTg1YyEe65p5xmXq8FARA4EqXvttOQxpQMFpG6FrOXUMh
MLH0oijxQhMMY7W15EHxfbLWSR5n56LJYzixN8QhAL0TKKOTUkSxi1mUE/iI
kIwuvJjj66z37qHvUxeFfrX+maaeing9w3x2T+xIJrzGTV36aGhXZt3XVFHM
XDHGuJGVDbHkF2a3LPaBtkOOjd2uI4tiLDsooAiIvYraKpD/uOVt87PZ6ErU
prbGqii6HaxbpqrCskQvaDk121nuRGJ2lNplSXA5LJCLSQdH2G1Oq/tQxpdT
I8nPqLHL3ptHfxYMlW5S7oF8wYrOQB/aqQB4HKorjUCfhXjMYKvYZSO2ie3p
kHUyGm2W3tIN2ko/Kb8l015yrM1YCPqkwmGL8j9PXOamerLjqT+rbTVPyY6A
zlcAwp/2R7dFEAAUEQBnMrQfTLKwT30NM24SHPKYOTGPzUcwr0JNyTINMs6X
6JJ1lF9O68lTTBBZKNav+Li9iTSzxmOK+2lZW/RRiKyQwLahSTLQDyzXiAiu
xJoojnzEHcMpe/qP6xIfxJJUyiMjg/D5Q8bi/BX0+KLI83+lXttfQsx1Ot3b
jr084HWWvHs3eAARq5dLtK7rDKrHa6c+15rO5Ifjr2HQ9DxYYwmJo5mugxx5
RW7o5ymoefLUx2xDLNj9XT8pwdZ//iV/SV+50O8NE4gPhqVEtV6X4Y3Df1ed
IHKUR6pYEPzcCws8vK0SnRdb0LVeWaItlqtzu4MJtCPF5RbifUmGIyGiSJtr
qIEH3+qkc1kZmx/wwBwYEJePl+NTK9+DvaCu0JOXq+eVJ1Tc1EObvk9jrNCx
Dq3QzpJQCMJZ+N67pQQb1o1PG8PRim935IO4UckdLHkcprb5+IJxzaortwDn
lxtAZZBRnyh6QLnELvjeihh3QJcNPUQ0WyCN5u9vTSKI625eqDcMXJnMVAOo
yC7C0WMoWW8Oc9kBRBnQZJnZKlbt1HZcvQmZ6kpoY7MGNbbANCsWFCQU7Y1i
8dF7Y2Xy6A7J9uFRio2wyVNonQJokSgBUoaSvev9NZ4X74aOzTgZ4h1S+hX/
u/KX3kcHtbX2wPJZOGdjCoNoA5dDvv3NgCSG4xZt5wN7tWsGQCXeB9aHhe4k
23RtutrbhR8aZfKnvqvIl6GKbRX4SujHcVaNQkbS8hqrq46gK5AK98xDywcX
JobTCzFA6Xk8hNq2e2dXgzC5XfY/fZ7PjrtrhU45jN16aoJjwIsnup+O/+7o
ZGWWWaBmpCTFuYnUC7JPphha2VJWxoB43Jbt7bZFYbWPecn1zj+1f8AHJkul
/G6TfFm3sHJlFbfBv+BTHnfazRCg4RFZYdKYkCSuVsTQAOsacqa9MSiD86zO
cC4ZKY05okJCiWEL2NrqAtZeJ5qAIP4Y+gN7l1luw3VIgSeOw7f79FkNZrYZ
ona2wLZAS6AF4eHQrmL2kDbVvFqJGSa4vuJrpsb/eE4btnbXIgv7iyMyZJX+
H2yNeyAhc2A/nfhcWjwANxY2z7KI3yCRpJyuFdpoH/eNOEDaUkkSBTtt5QHR
9jSCixg+hEjXniFPnP7QXQq6UG4lJVtOqZTjf2n7YVv5ghlUHdUD74jM3FOW
jQr+3PaveuDLnA8Kk7qo0Yda0zxI//z73GLQbUB8J816UcNY9weAz0g071ca
X8/3NlO4JVjsmNrX6J8it7nk4o9BxIA1kJ2/4M40rQrhER6qRnAlsR6ZUF6D
UcPRVJe9CJGp0I9cBaBeleRe4AZjspqGqQfZy2RbM7wPbEIDuF7VAKQuiLer
RXX7jXoAKmN1HfnSy1YbJduQdySyDPr2ulv+u1dBiTtmgSYNBJMt7Qb6Kwj7
yI9qENwbL9lGgClKTKsak5FrpgI1RVZNIEgsR39wPs4KxQ3QES5K1NZg2XlZ
/xasLJMtIyyiRZ9tTItRbdbz6Is90z7mW30lWZbWk/BTO8aaX5OksDd/CcJo
pISu2dOwUJGGNaD1WjFlHNOJ9J1fsP8ppk9QSi9JewFsRzgdopx5dUCDEBR0
piUxryVZjlWCJhrhPsF5rxd203Z7ZjipDR45BMhUdo5PLCXzEGrfW+ZYT7Tb
BD6XImwJY36kqw6xQv9km8bGwbK7AjKLKqwVD2g8GyMsz8MM0ngy2n4Y3Vv2
wpL92tJpzLzViYl3iu36vE1w17NLBcby5YLckSGJo5X3r9uX0HjNnB2789DS
sieto0ac0XMBLA31g/stahQAdKY4nInxamt0nzOLegoTTB2f768V5IGqCc24
pXRQgzVQXSrFq6+GGC9wLNJgGbtB7YYu6Kc9AtpA9sR208HEdlqA37FnblGe
rihtFtxNpYFwX7pvS5MkXN0DbhUuUPlDAmjl8DIKJZtmWCR2feis5VcmZI5r
jsldjBVvpyAjsfYdPe4EDXCr0fKiVJ+iaEeK358igLvIyRxHKP9Crg72OtuT
t/eZKCHyZeffSltNDjVFsFx8KCno/9of3TKuuohvLAOlxuKLPDnmLm+rwPPf
0ItD5sLcI0THoJaIfiocYFDPaSqpo1eLJhGuD32s/83U8RqKVtDJGVnYs82I
Et+fGDUo5fLAc+pZx2AAs/GUy3s/T7NqoaHR04DsHqaYPCnKEUJz5LOnxOB6
7KDFKrT0NoffZqpIncNRuiAW/0N0RS1A/auLsGGw++ofjWmdk5McY4fHzeqD
FAHHh8wR0AJ0y5XDdN8dTRSiSaqEROpacQKN9Pz5vf18i6c4PvUdjaxj43Y9
3cnX8N3hqUSeVeHNl9HFM7OdKIDduyPtz3M7ZdpFYBf26DStaStclVw49SYm
ZeHeeUJV34siv/pp1Ty+v43LLQa1iPM0TxRh8kyp7hmlvWQKOgph0nDeatwa
WtGtEHhMPFKYJH5Te79e0eBHH9kTvrTGh/z6nRGYu2mYgo3/gfUjgOrR6L7i
jmK8vZbeWukHyvHIA3BMeTyT/9+DELLbdF89xAFGeJ1Rx9y8PaW4b1qZWQin
9Xz2NgW3eovHwDDkLQ7akWPDBA7gEqbM++onr7bab2abXT3WAXE7ymWDcoK/
iEoW08N+S4yvs5k83qGyqhRqJJF5gj2il5GYjlTo8LDEFahqNVI2nrvo1pXU
JxxNV7HeRg/aD7jF2SajmHq1QVHWnbsw6kIDtGHPs03VfpG9h8aQPYg0KUrt
h5UajsXzNYx+fUf27txDttV++wO0b1exg00nMLJfJ9FEa3TQFxDE3S0+YwNN
0rEV1C4SdFZLIOBvZz8RMLXk83UVYBQyAI1+AFZtMnjnaqk3Dp6VWViHnHE7
15TinbhvETuSzLKIUb1OKOfzV8oYx7Ni5FTQRhhEkGww3yt+URGgBew64iM9
X4ixgI3hShK72CBeZSeZyv2TQBjuT/sDiAadRbtpKfEAmgZgGyH9q/JcTW8j
fRINL8T/wTcsVSMH7UveCFbNycD+O0QnzHk8kJ/jaudeyY+qVv3fTTFrLbpH
a7imnPdbsKHuBiBdFlgfLQNwY6widVWn95gSducM/mxYr0y6wwJk4Gpa8aju
hgZA9uyH40OiSecwWkxEWM8UJSNV1vr8NLVtN22yfh9hLzoLHHC7g2atSo/w
c4QNpvBotHBg5CoR6FoHMLuxDUiaTjxVS81Vd4uayAGmJnQgwEX02HqjLZWe
yhEsskZPd0LB0W8VyvSaO2Nz7aYdW9Dz14utcop2Ny2idk5VHHxTd2lfFJJb
2vnJ2Xl/40I/i/hGsW+XlooMGNPmIoLcrRYnvkwCVwdma33rjdDLvQRNp58n
gxHaTjzQfusesrnsTI+lsU3sIsP85Pn6zolvKZ4PiagwRpB5wuH/FlezjMAn
kMWo+hpwp5pqwB1xZDuv1XfUx1IMPJdody40pqFEhTGPt4SyFhvkHVqvXzkf
pSVJez1L54UT3rmqe/CA0pF5lMJ0yB3jsNiTuwTW5niyQL/cEhOyX2m48HF2
6RUkZEpm0n3fv2l68LWQHyKCZ5oINms0xyPaOJBp6HTZECC+XCH4ToxtsUlH
m8cTaP5xEkPblNm7PlZS9njisxZYk8mVGt6ni8LB00eMCpgOcDY2QREQSr41
TWyBI0FfPcO1I1uFf0I9kl5ej9SyHAnn4dDjunCml0uYirwZEzuwi1TQ2WHH
zBYae6/tBbWfqmpK6FKSK6f+KsfHxZX6PTBLSdVakJ+iJ8xCgsb1DeXbDlAC
RegcCIcsef5sX4CCsnvgKlh7sL5Y0KuMPaswhEhofvzkYvf2iPhaZYgVBuad
gGGvqCi3VMnhH1gpYbEZkWciF+k1USjP+lK1uIqc83IQsB5LW79B19w1nlRi
ZveQRiPHeOv5keImY8VP8eyGpd2jhkKw7TiTmSoOjgXCcI/2ae6UAr5XU6BB
np6OtG0xLHjM3b4ilUARSw60Dt6rhHpoDFD1y9O/CfyUiE/OfxMvcRn85ta0
HZ5TOHc8XOGZtfMzmVp5KK9SypNTMFgskODJcYxcBitCMFpOAhE/TpiIkEwQ
CsHUQtdoa/yNUfUXNijIs/unF8HaowlEmXI7g/sy8y/DXnCImsLzdYRBL0K6
FOKnyJH36c8uVgDNs0eHvDPVx92nYdB3nBdMkq4iwScdIkJzJk5tDAznFo0X
6+oCbXiMrImH7r3C9AHnmWtS4XZohDF2c7M2jOxCus3Q/ddWkzvTo4tWQRpC
9+ihM3TXgYzkWyJtDOVDWOOdy83110pMFC3e0Tbw5xs775CeQSwTtWhUgcbM
z/PTzFZmn58UMGApjz0McV+jlfgr3IAAHY4Sz1KocYf7TxPGklLNxA1LWVyX
iRCqdlZhSvbh45LxSkbob26caJxIC52Q5KuFgy5tQ868HdVeqr/uo7ubnm8w
cAKeAr7zSNs+sqD8y+34kdH5BeobnW07UnO9EnSBUiNXtJbAJstn0OGDssFy
3AiTtFwv9LlEiag287Uf1uxMax8TUVGmPs2GmEjA70GQNKwEtt5sZyGUp783
UKJ+YTAZtYSWdCNhjb3mfhdD2KkRfrJZYRaA3ajtIZo3l0ovKXg/OXxX45Lr
cNlhkC7WA++VllDRKZuElGdJss1rovWIrkxYoeIQHRSjf36dEicX28TC9c/L
O5Eroj/5uFYJFe8ECCrM+qUXRxUaqPW3PzxBpYbGOg0Ul0/oENv4BC/fjo52
kM8210PV8+r1qlnfELC3AKcQlnrKp5gFTZD8l+obBqD9bjN9P73uFY9mOD+g
Y6VEtId+1MaTL4E7ahjkDXQvStZR9bkMMw+d1bkv/tKqwgmI2AGH2YzybxTZ
oVeUqa4KHlKJYSs5AbrvMu6Wfnh6xgzOsIamixr6+TUDHZWtTWTdGNS65S5y
H60bPNcglCPQEJ215zYEaM3Xw/LDZt4Z1ZGNZuKveiIYOMQrAIBn9APlE03m
WdetlkhTie3WTgWF6EZCdSGOOn3/J6LHc24RfcrYSLrdMg73CJmhs/1qVZN+
Kj4nU629DiL1KRFi2cYu/W3eusyVU4YJu4wmjEa/6mBn5sB9q8HFEeQeZG3b
/d2QzlYU2L1gkpBpTtkANfJ8RsWnzz2B75rL8OYZKetVSdif3Ca4ABSvF5T7
unZ+ofgTr5QBx3Aay95X52ofNvYtBSo5kZutdKsRpFqZsN1U1XRMdk/YjCYZ
VN/1zYFAmJU7nIS/FQ211D4GvBMskIx7BcBaYekD0eoFGtJQ36emPNfJQzyz
tRlu95BbK47a6ZcvYwwdljTLyjjCGatUxry2vNSbMDlneBXe68MBpLzIK+Zt
uUOP5ZNdQMixFj/Tas21pOob/YKbfwVx19FiqxMAs4SL9GJrPSk20i3MCELT
Lc+6ToIDAdCZfCjj5J6A7ZxlDzLD5qjGRi+aYQ/HmjqHi+H2GViYS/5iExG+
TMY1oUNDoy8s/E8oIwfkIATItwcNzbKppLoJyH+mwP5V/RzcxQlYyu1pNi3D
q9kqkX3G9VYaXJc9PADuTTInvNKy8XnT6kWIYmtrhGfi3h0xn7pmI3H6ZOmW
1OAK3I6yQSTUpjq6rDbFVRQTzT3DvM30WhuRut0fupMSs0R61wnc51fGlzx5
h9mlBKPyzEkRVjXjTTD4vlUC75TnREJ9GNFH5oiKBwRPqrCr/zQPuLl0GwZd
COJI+iug33Gq3/UP00kyWHHlY732N41wIxbLuxUK0d9/y3To9FAlmEXgRZmI
D30civwUpQwqnSns5O51rtIvEi6Sv6d+uXZEEUUCN+qoFkMYlA12/Cw6F0An
xDC3cvvbE3M28pyazB7Ji4JdauP7LlAi5rU8fI5U9RXLfs+Yqh9ci11bDhho
X6uHXHO5VHE+10AarkQnKFCWpFmR9gHu+GVoM5qZzvn4tvpg7TFz5St6Q9Bt
VYOdUOkK9EmaY7m4BF4hx9SCFV1HDA9d85suTxw80eTu+gbTjvumGTyZ6lAI
szn9REsMVjcrd1s1iDTxX9xV/hgNUkj4eNhexDVOUsrEbPNkHlrHvYfHoNty
CJd0GamfIxZWzAh2UoMB1qlrgAXTkSQBbwh0BrKvboTt+AF0TSHv8NRt8jf7
Tik7ujBC9DrjWYvdB+HO6n+dPavMp06Ir6FyaZn5VEodJg8VX5zNWVyRI+MP
4tuIWg6BYDsUliuvDTflk2+2rHpiqqHyF1pCoq8ajk4e7o3ygoBBlfL3bEJ+
8kb1vJmexOMdfFy1ctHF5l3YV0u0ENza2n6RIC2Mre/ss4QiakrOb8qq/Esd
atE1EiTRSbRrI3RBZHYjZ4jDlFtarWxDx8IOM8U4dS649dTDs/jExsWy3E/L
Yd3/zErGhssi86I5qSxIpAgy5aZOw7bbBfq6bfCV7rsfES9jOQ1pFLZCxgDM
/tT5636I7VFBMZdfP6pzJbLzGnvMKJtkM08xYwgudgJvWX9jOuKvPQflEzRg
BJAK8mN9deMSzx2yVH+B3fyMFl6so3JRsmsNqDJH579deQlViJ4yxvBcri8n
HYfFrSiZ8YRUmTDClxHEwO4G5T467/uRdVOxk2beWzQyF2Al/L5PhTdI36SN
3bOHSvsWgRXFS4VG/Vzsoyl5rpeHuXaryawwMFo4eCvP34j9Wfva8qKuocKQ
46T5bJOsL6FEQc7kX8rPFCiiDn8RQ6XCYXi6CgikZXXRTA1l3eQ6WN+smnga
6ZHwQCGtpL9XhHK6hYjn+WkZC/JzkPEqGrcFNZ7Chn8XEEW97fl0O1H6Qdr8
cOGCbHtUjBe8HIu9NTHc+noYW8MN4aK+Td8NpU4i5R0LUOzzXWFKOn3d0koX
IwWL6zpErvFpXXSu4Zelnx7kuTyCqpbalhMfy4V2mjnGbmsKlJGgVR0ky1MY
+kfl3VKujW3vdXwhg1ZXfYgVc+3pFwP/9+UYzte8tJ9OruPivva3cCs9Zca0
vPsi87IqoUb5dIPZbCXfdRiuetmhLgyyZ1WFgzhjE4Uq67vHgt8v0l+9O7mH
gUVd04ZIKCCmnzpSvaDepb1Mbh6j70PEhniIWblpy1k66QGs4KbhMwE5yGlN
yWNJzCqiEBlqncWP9PitXBlx4bTWUuBou1G38UOBnh75C9Hfo5pzQWAUHEIl
1/YAlgRjIxEaMOGvkLiYNziMMdpDW3X+jh7zf3F20nTSyus/yP+gXXeG6F4u
7t+Mz/5qScTW/AIj4mR8gzgXki39BLo0MXkYbe9ibJkZ/0EYrms0jly80PEs
Mi1gtnVkBZzJnCHx3xw0eapxhQNRubW0+vqsbMwgADlEaY5P5YLg3jlPs3Id
wwmxNDIPDeRHHlU3WbeZ7MOg0qars8ZbF3i+QnfkdwatHbllIS/cae7ploU8
EojBbktU9ApGGt3e2mHN/3e9KYwXvLWbnRl3BVIWwdeZQboC2vm1ZraEt0SC
lCGHUjwAHM5nGYfd1Po7Ted4z7pJnGF6kFqy7zt0jCO4IT94ov5BR3mmYvIJ
/HQyCrNdy1qYQq986ck8OX7BJhpho7HbvtY1XpL7UFPJdAlni4YjShOHsftO
VZXMWtFiaCuBbP26FwoCd9jTR2Qh3q5/t48MXIEsyL+uWIv4rGxamPgKOMIE
XMXKBGgydyWAnL7vM3HfZRS3CkaEY6xiuySx0QgYE14lBu2zSMf1Us0OxDoR
mPZysFMMcquYf3jL1qtAT/I/ExeOtXgQ2fW4tXv/azDJPXDSnQmRHd+KDxV5
Y5eyCRiQ5WLkRE6Nvmd5tKh5qjvDjCWfV6SzGs/rlqVY3oA33McQBPLoRZ6E
9elcw+yhc5EfRwLBmAHbs7/2XQqJWTDPYVOFa+Qf58+66wT0uINx00Qfy93b
lGyPaiGbqDQtZvOtQ5UkJgKZjxCqkTLae8gR+5+k4euOTRpNzFNOKt6XvNOf
WYJLkIrw/msJgfQpRfohAq1erDiex3YqyhRJY8BIz6dlT04Jt3T2W1SVXKT5
q0+Uh+dY7vK68eMQ6I54rI1kp9+LXBVFV0ANqcSPAgfdBNdQJQ695kFl0OLv
rgDoQL909miBgzL8SxNPXp2RB7MEte+/SuclgNj01vHo+fgUAyDVp7nVyNzl
4zZcIsGQEOgL2SbQcACEJo3+n7i/DNkeTBgs8nQtzOIrp6KHCGXhd0umhbKy
lz+ztMkrOVeCzPWn9Q4J8mUmhWYm8VOp1Grd0SzLZB+B73EgX7HLZxehujAZ
w+ng4oq5gUGqq1D9CF2He/E+KaLMUjm6NM3OPj1bNDzoPc3VoaFLOct5Sa0o
u1wUI0uNuyXOBAzrpyik/KVlUYjKW+DPKB4axGLkKtT/t+lWIX4VM9BE6Q9F
QU2udiLmJbBi5kKC80ediG1cx14BEeObUcLQAEF/JElwExDdMUj1cNfbb2KB
Qk0fmY0tKvM8HS/HGuOYpuuMNWk0Pg53zUp1DkhVyWtjuGFyysLuDlnA+GMR
Z+YhKmZSyS3kcfVv7wHDGsuDaws8s+TVYouiN48vXcVJt6zdgdyOC1QUctyX
QU6aasWLKoUvm3gDyL6VF54JCeDFjd9DtLiUcTd5Ly08PLXBg5nKO27RioQ3
7pDNMicIDPygShpoXbnGpQYYAiI24TGyAnTMTI43ZpnpG4cXGJpbPOA4sXAH
2EHoO6PK3B+gUzCyLlxps9/v/4PfSV1X+gB8hUax1lWTPUyjjOVU/gEyfBxY
IeRyU3YogCe3oKSVIIxDshQGH/P4WYWWClojNPWFzTymj3isyBScmsk6PAj2
oQvedKFsWZdUCY155f3ps1viRwKHgh+R/Pr2ZMpS21KH5FLWesQI6is5JllF
mRoVp4VZBpqkB3wAQQNdIMJQjI7YD/TvrqoqhJVP6LXOxFEjS/+yuppx76oa
TRk9ZMABqqlCIPLL2kyTEV+RtN1mbgYL/b6SEombik3ZKpD5at+b2XNZ5PA1
+tuHDbsZEMOQIeqHbhTJhf28iHtSVzV/c9iT93YCrmD43bVYhhi5lpQHq9dl
HI0iopCzJZQLwo91MzRq/A95/8T5hNflcMugA9jMWIkFbPYIKYKzxHIiv1d4
CydqfQ7k1iGCxlhNnc87gWkMssMwTSw9aHlN/o7Zq5nZ+QxB5JhspS2RzDlt
FcGt8tOW0zjk/weQCU4nlD5yATcqLOUT3X03bbxlcnjPMHrZ40YCAaLlqXqp
K3u6Xl6pjfZlKo4WGiDAS8HWVtnbjZaWz014v8h9ZhL+mCRGNUig2Ny6xumt
aCA2Bejm3LUsfrYQnXnLoRJIulD7tQwwW0xOyIppfHUmSX2qLsC+as3RH3jo
GRqF7krOg0XgYDm3i5PCgr0zAZuw93npeuHMoIWVOmYx0hgBuCG9RPXzU6S/
LD88TYEBPZcKKe+3S0U75tzf478R9gAYIgwa1utAxK1EDa4lsZQPqbdbJ4OW
uLuaes7OLrrfXMUNQVCqXgyoRkbXrGepn+2cybjeNx0emzBC+qHk3bSKSbat
sY08bHHdkHdeFQEinGOcYKEdgbD/QRaBV/wsssra41TpHisgpuxu04VlDcai
r9dyAF964sy5YEfn6KqvmBkDB52rCqbZ2dZBP4hei33wceHdFxypbdDBZW0m
DrJ2yAhS3eF+jGMJAkUgMAljwR+RxEl30YZrcfCqvvE/hCJo0ZUO+Ne80AIp
WJwojOwA7vLhnIAwXh55hlv8LLJFDO+QmpGVTThknexWlk8XqL4fQa0aCPe5
5vQvd5VP15ZAve2dWtF4cMmbWPKSYeLQvGaiNq3vi59cB/ljNUhqjS9l20yU
a0gYIkT9xPVsJnZ+qUB/NDGjEklAXOfpuf5FOFL9WtDDABcOabceeGOWOVaG
bjCFV1kEQpDb/mT0GPosbmWB2Xo9aDW2GydCcbgqGNDRVlKBdupA20KEIyON
JCKrrEl4h53C1SzkdRi2p7RmSo8d7GPZjUgqjonmdx9ugRjbTHPOPzFSKcXM
X1AI8MVEdLsTpsJOnXI6Lbi5nLYdmmSyidgpfX4vz7zeCBXfTK1LQgLqDMWw
+1oMVAj9nQHT3hHKuMvBmJgC+F2PR//mcXq//hvxSt5vcciy4g1KmwGmJEBL
c6qJHf8AInuzKBS/tbwjyKkaiOtJzdjZwZeSlfNwGGcWx9GDnPuwJ01WjCuA
gjg8SZwwwccKGYm0jNbxGTIGxB0NPDYZq5kSP3jkXCOB+TFqvP8R2BDp+9Rp
7AEWl0aYDTfzBYzFkLoq1aLjC9WkFtxGgUv/0MfkGnmaS5z4rA8/7obae+0W
CR5v4/P6XiE7xgl/+vi77tJ7hrQox389WshJfW/WudvmU2FXQ7t6XE40kcuU
90UrrmMcVSWSAGzdX4god1O9Ie5aNHxBaBTfTogJFk/RItU3528Lhiw1tyZg
1dPPTVmYSG+IkLFUqZPvxviPwtNlO6PyLcnrLYtaARFh+y6i8i0Z2ogaVkvZ
5gCrRiUhisBa8h/0twYaszWncomyb5cB85HrqyPKCkfdtcbK3KUH399ulVC7
Cz6QgHon+xSnwjC1eBAwPJzqgH/Eqr0Yo5PGaoIRxYE7wsdQGEgii/cq14M/
vbIP/OQEsKkfLU1w3N+YWI5Lz7fcBn8B1ZLlLMDrZ3Ext9R9HA+xWjIj+m1V
aSZpLr/IN18qQEmmtTX/8INPDK+Ddgf0PdjYCSdPvYUuIvaxJ8XEG8rj6BRL
JhsGtYEerbZMbTHsj1azSJ2bix/16PeA0Ty6LwHZi0AfL6ZuZ6hxhsRk9fC/
13GlP7zvf5dsUC250v6wV5Awox87s4eDFFsS0r3p8qKuUjk3EyY51HIKHHJw
B+GALlWtIuxGtkX7m2GYku6/Zo7pHNSRLG1MmwXemIqzyK+2vRBEwmP6omNl
aEF0mYIwwiANCkyRyXDJOmNfDZtm+o/NyZRcTKcYMrAgR8O6+fQVp1Mi3jHM
LnF/SuF9og/3MQuQ22o0uqOcPYJBk42p/+U39ez6lBFqxCTl4chmMTRfjvv9
TS/HV4VG1XpcjfytZAVoy2xQspnco0J0glNNhbqDaG8CChkWyfC1htU6SUox
qGvLO7WKPnNDXbKqTeKAdoeVPJCCYHxkK1wJRCQ+SjhCLBrjBjPVBy4XTLZT
VTjZjnieAvLu+yWjQcyp6u4fWrzuQ+Me8pkHLWQWrbDWlPboSNiC2ijsSexu
qPEXVgPonPbwoSZd8+32hsHExcbE+gYRHA2qwGgx/P1KcbhaFOgy2j64uSaq
d31bTXO/aLOIiCkBIlQvnpq9GhwQ1cMySR2nUjUbILTuNREGjd0KHZY16WOu
8sF7nWB9FXVa8Bi9QWEqtrUzejFzZcq/l5BRRBiu+TL0ZVbwBlKjp2CylU9i
BwfzA+Fvw1/JTbZBZbO39QqEW9Zgm9zTkOovJXBQSlk9EUoErnykIGT023R/
0nm/WTzzrUlRZjHHdKpF9jEmvHBl4s1T/rKkn3g4f6GrMrPwWHxaK6HQhDQN
XJ2QV3iWMFR2vYFr8KjxrsIukDrpwWbEsu5BW42XS/ZnptK4WMP0tjFoc2L6
8ip1yUOR7/+RiD5QPWjQV1F1oDbzDL/7usya4D6gc0if4EhvMmaBi5uCk4S7
ypu/zHj7Tc2Ah8/vTRCWEkgQtcrZMMIYGPUoYrnFteZ0JGH/+jMSX77eyfl0
08EKSb+kbsKnu9c0wcYhkLP9IF/y5N4Au6GBIXlSMp5KLIKzbsCERHr2T0Uj
MAJ9qW9Vwb3wJy2TAXcf2z2K2eHvjKC/CzZSXlbwzAyz3QdfmYkc+uWurYd5
lJxVzC+l126JOeQLgl3KjtyY7swkK87x6I3/2kUHqo31Ghnr1s+b5UIr4a0p
GOYONCb6aYVs7fTDZ/ASZsgUp5IqcCa3O/OXzV9ZCOoks/FOK5zJ8aduT7yL
b3B/n4BMimxJy/mN8z4KkClzikOyF5cWFhukWNLP2mRkkne4T5WxQgRSJK2Q
CTKKS3zXzJRoWr+phRW8AXHJlZUN5NruNhenwV/j4ZST+S8SzCTDDKjCTJJM
5nKlAHwJfNZqVQNG27YW/iFCfW9f8JaKHMzJBSKnb/rnzFnWlEx8/xvnYl96
nXuSbMIjmOY1uMBHJt7/o8ECgwg17gHxy2h74RC0FlApI7G2DObpmQZnc0KR
wndPDXLTTYNe8Z/Z74v3drQNElBV25zEeRKD+UWmLJ+lTx4sWMFU/QlumK6l
SGBKEdEjvTWUBS5ucMoIMTq2v5pK4CYzv2tWFbqPY/0a8jDKGp23VpytZB38
esNgKkCDfdNKE4X6eKvYxaqZfVtE9bUJU0o3fi4xRy8bF9sTp4t01YaFbh/H
o18hgVQfpAGzKQsM11VWkVjCWNcAPTe93BeUjlA5A7T3AiVOHZOaRLpkOCpX
mHaCkZHEDCJZLJ7ZIwJCCiXVIxAH5RM1BXE29BYWZjtuPCmc5uQpM2nSZ1Pp
K9XRpFvJtLKzoOaW2DATLydIVahuaC3YwKyGzhi9mdK6rUXDfXo3WvPFsBC7
5XYNfZK7cOvpgcvfI7zY9D/KHP51jJeeqcQ3c2GXxFRo285YjWhoBpwHrv5C
CJS1Q8b5hkzzVCZo+V4GbAg6IK9VKI7ymPGFNcqR3ju8WvNk5ltxzxpJh1XQ
8guXZrKavdlzJAawR1gYXFWLdi+6SF77KulzdG+q9oB/M+6BRb8LM60Giiv0
YFz3vVyo+sOnQm3XX5HWao9g0BHj1/DD1fPyBnMszsZd2UM0bfDK82xYaEdz
ZF0PuRgqAO3z2hk2XH75Enyn/8SX2bXyIqoNEhAABnDG42HkE3eseBEptppw
EQrjERSUtS37DhX3Fwx4L7iW966G6B+p+xJmjKQNqbFChYriKBVqg8pcVvtm
CL/3VlIcLFQwTrNxfM0XWSjpYXXZ6TgDKS2/EpdS+Mx+K4ns9ewFtSWMrwEY
FPECckIAODsYV9jPAdwXGQWc0Xtkdv7uBw5pHwo97pdwC93DRTAG8K8tZnWK
YiT0DihDsahehBGZJ3WjeBs7cxRKkWozcoGTAlktkrWxsk7xsGsTsx0BjNHj
ygyNqjB5fopAFJTXuL7HSv4V0RntcQIog9RXTfg9oSAESvzFxv912G7xbZOu
3rpAHN/JanDJMzlI4S0f/pOGMylLKbYHnYIvwU299s7n6GqB7mlo0h4EpTqh
kWCgHpHDCFGwMLj28D02SL1xAgBlIrgPbydFB+wmNYBkWa3R1Z02vnizvM2O
OH+W4I+a0zdU0rvOMB8KeifDeLkUwnWCFmfngO8hlzuNc9YPIaJ0jhy5CxOi
xt720lbl6AQ73kpvcfJmbrPCniuw8g1hBMMDl3DpylF8ZMKk90518TY3YoQX
1waWs29H632/tkZFSBU+6EkRhz9vWBoHD+LrRevt5k+Fz50Z6ju8XU/wK2K0
lvNtfonqUgMsWo5D6fS7LnCIjFtxQPLKvfzQBdj/jfaZzLGNWnB1w8vm77wS
87eH36sFRDRTOwxJOxJ9ccAL8ndE006mEib4yaMRt0B4SOt3kQbbdYT2+THT
dV/+AQUr3g8I/P4iclVcZKPi3TVa0zSNlVIWWL+VVbJVCuGG87ertimyScZ0
actv75C/J83LgdrWs7jpjWY5fjfIxlntJXfnXF5iqcc7p5otb/dYT6Z+pbLs
r7TZJxAdlmCbVVr3lJZMfUAhwPzDzK69LEWJFGlS0l4gwoa/RmPrM+FGkw7R
0cNDSIYbD2QxswlxYD2aBsUGnxeKKgG8krAazO4Bbk+XFtHRYVAPcHXLeTej
h/7nTgTbo4Qn5JILfoJPuCyzirgiT0SN9FyEbGZJg63Bq116bmLuHA3L4jlQ
82i8hl8rT+fDlXvrT6I6bi/rcUsxmQFfGN7gXHa2bvkB4QPVtKEgFi+hlcT+
SLyEPQck4MkOoeJvGjL10tW+wgF9gw/sOFQNrw26bNBjNYbQvszuj1P+VD9W
n0pin00BoRWKBCQMeV5wWF+0aMvYzINAptZ12QgFhnaWOLme6Jo9ZZBEybuG
EgGLJdz1fd78zvflCdh8wcmVjIqvqJaJvDVfKOTTEZrhQLDJjMGgWsXH3Cc8
cB303l6WqWBUvWuqOxI9WCSXLdLRLxI+tbj6aFdR0rJanmYrCHnzRZxbAcUs
ENHZOwlSiOt6AMDUso/+ypZ/V8qe7trmvxuSXmSjPHCex2y+iB23t3NgVbNM
7mmH/1Zx9YidURnL+JJ2kosUzKjPzmJOEa7lfy5ZoToKDD+E0jibCwdaQ/vs
L+sy7AHm6y5nfvf138hieCJs2J5LluI4zJ5VdI6auAPYzDEqUSwfYsNrBE0n
ZhV/3GewH35A49KhwdAApq33obA1P+PLvBIpSn0ql2FXEaonwlX8QxVYSeSO
V5lSGjtbRdgG7lZsMEEdEieK/Uqt32rwilkVqVcJkIXHC+XMrFGV8zx94xcF
b5gJiAZxDmzWLGUrJqayNqcj/DRm9X0RPEG/G84v75Kb24qC8PrYcdCFXBLS
PwY135ew3+aSmxKKA4vZn1eL4eIPnrN6szPlcpS3TYQp+n9krF/tqFy3Ndjm
MH+MnIGM2hr2snzM8ugdta8tQOFU898WYNKKUGU+JmizCcvD/uENZyOiiaRD
+Jsd0YByJe1no3g42AVylWzjjEiiA2DynE18HLjVvcFuVTPGnYSaEZomyil5
A8pPCS2dyHVSbUKGE0+fOAed/1X/kYnPAaQgV/QJbnMurMZ6G7BIxR73uO1Z
f3q6dHAzI5UFGVymwbGKMx/p/eXhOBuWCmmMjajzXqvDjju9+PrsaF6lB47S
fSkPM2GA9xrwgxn8vmK1sxwtC52xIEJluP0WYGMfDP2Bl5Jk5CvfxuL44GUr
9l8vSk8JM3FnjDmhv7O1x6ruFsxtzqPZqzZMRp+G2lSEKxGxnbon1/NHq0sw
WNe37geHe5GmH/lfrVQrKvdejNjPE/rWGXsgYSCtm4KhBPY35rdAGpD1tNtr
+yeKZbphzLIvJnijnSHOapYrzoxAbf7y/2Cy3N6uGOOP8LJa/DMqm5sIfUpq
EXamBRO5EHEV3pktNnhZ6pEJNeg5NCAyKUQvQCTAZ1mHRAB/44LbVzq6Bkom
OK58GzzbebKkLgwfq4/emxDqUNE5Ot6ZI+9pSciWs5HXsTmsXQhPFqbrJN94
wrbEj/SSD7SdEToSyg7XSwKhDyrDNpOUzdquEFn4KdlicwADmWS7ajPSutH2
HJj44UJ95hEJ4VZtjtXr99xAckSWeDeSYYJPF6QA0UmHint8eeNkJxr9QgRH
/t8Sraqkz/pXIDWJDhlYVHf60EITgYlicSV9b5VI9GMAwTR0uMrGJ8c3vwx+
JGLBL4WuKZdXx8tvlvbsWQLO5DCZLDK/F2/p6oD+4FMk8X88wSb35Jz2C62u
I1xQoMv+mva3WtOXCSAgVDEwhl9wIlcykIEai79JIqxr24bbdbpkDc/3TxVt
h65AacRxN4DSeZBrJiHnjb58q1fOs2r6wLls8WqPqrxHO+VfB0Y0FBrLgFFg
evQV+Rpfs7XuFP9iYzN0+ZXKO6cy4tA9lQVbgvwp+Vn6zzf/g34+WqPYMY2o
LikRJsNpuiRo3K7exfv0FtKqW7unvfyPF/SuYG1ZpwcabwYE0/6vTJk1jF51
K4A0zW7boxrV5YsKB2owN99TKuf4GvIPf/dL/7whWgkuUml54mwDzdoJ6Po7
KtBq6pmWHVZvHMlamAZ6x923nF2qKOwsUt2qPh2mK6yoEzohVLxDT3ZW9v12
7T7NXv4Mw4J5j+bhr5ipkpH5VztYNKvTP3QrRfLQVG/GcAgac6GMl1A1V/9Z
YCpG2aviLVtf6JlWmw4ImGpnotrdxJJ7kB0dHU22bWEtkctWbgjhksc1M7WL
5lhhJP1o0lMy4p+IIP3Htppis15yAezbUFM+bwNceg/VJDqqHTlS/G5o+vUn
ZHjPbLP0RaVSY1i8Pu7ZmuC+wrukQTRtHTOJNEL2s6khi0WuTwPQqGkHAYTp
xUeGeLf+POJ0ri0YGN8fjR8v6IqtEZV5ozrHZHZ9vIHBgBJOwCWbZtRYqAsU
HG1hKGcog6Dnu+rtXUginlqkGrzGZ82LBllBzbb5FuCIx9Zld10Ms6nHWSGB
ON82wC/wKGFYv+tA9oUo1PvtSo1vSPYUagKbNyhulBtALJhY46I64NoP9tGz
RdNBuYuGFbrfK0zI12M+i4ORbX8PTkvpk/Z0me6zU4t/XDcDzbTVZCbsX4i0
mhW35MoZfd5GXaCjuKfr/HRbKWx6cteBe3P4u4VmjOBczKEfdIrHQv7eF18k
+kaJiEhISf6vieK7xIwJcNTRrY/QMy09OPKnnzj5hYnf24NwPWJBOvAcmahO
Fd2aMhEicDwAfWNSCAWr5J9bWMrvtMwBRwSEi52pmZVjE7f/sXqUPe83yury
oc+jABm8FIEVEvYdL5XUx6RcS45fVG5U8tazBse21hNaGpngsqFI4rPPFdTp
cHWO6StqIy8HYO+5APl0cI/5cILMvP8pAGvTQSAco0dHChXtL3CtPRu3bRq5
BfU/ZMEINGUvx9YtWx09RfpFVhtw3Hk5j2yVOT1TThjAKnG1mDrBwpWrSZ92
RWFeH3M+VieBOR/5gWT7Gt7tP1GixpjqyP1E7yBxmmNEgMwrFwLm7AvqP4AL
es+2ZhtGj5B8CYoC/Fu6z3DuduEWJgern8JYT0WMBs5HzFnf7dC9f6vO0L4f
y9utUsCPLV1rGBari9m23n3gcRSs5e0hDCuKjq2luu/UCgOwL0TwmhTwCp97
3IhEh9/zaBJ9+y1TbidNxQWBHF2L45tSwjmwGBsnHFlT3uCGc5Mzdm99JF6L
jRvSpca2/J/kCJ1oygCrLIbGEG6n0XT91G7Uq9/yx6NFfOhbM3PCmQL51kSY
Onn4nT1JcL6QwmTTo+2J0UBB0W4uVYPlUmYBYp/sYY5DU1ZPwOMMsqhPCmcv
tbKl+QeUZ1uC0ZPlf+CYnghAwewigMXs9d5G+QCzgZmW+mNzIZkFMQiZ1152
oNL2XQZf+fGzTjmYLJ/o1N1DHkZsijXcB2u+i0ABo35BP2CLSGu3ihoQ0gz6
P2hAjwHcTwYEFL3bDo64YVk3kyfpxvUJX0+3tTHHaLU3GHptCGhu9m8w+/M1
/ClJWJSz/rQR68CnLCrBZt/z+w7LILI/xDD3C1aM16y15LBOog0TPTG2Udzz
/K3ZPLvi4svlUEPTKarhF/e8HRgsQPMo+08cKYdRCzsW6wAz1qrXqU2F4Qk+
5gJTQvQ4yVmxPKq3jkpf8aZ3aEk8cXeECRbrgwkPIjORJtVwjA8lDednZpHX
eerQ/YKRP9qRu6I3DuAzeKvLRdDMg28xBrlwhF9KIBv5mSMzB4lJ0xH2UAGi
F6jrcoLtSYxmlPyGHnbdgkwqvXFDpQVbL50BWhvnJnrOIwhU2ZqHBues8yKw
HdM0OQ0j2gD769Ga5qee7npoaNtHjdmD0V6/1aI4Lq/9nuQvk+rMhVesRqDw
yphNpP41EGVgtUNGfrdQ8VDoLZumXikcM6BVK9qZv2xIFsPAVja3sM7CZDDH
GiYTKVMsLyRcY1tozC55g/t3g2Ap68jYz9Vd+SJyMyg8WVq8LEDWL7pk1Ofx
V53Bbxa+MGDl4KeZoXPh8YmtEuPqgijKiCfH/tHBYuBgSZOAgLX0dxxeHgx/
zeItVGF65OIqI1vkLOcXJbPrx/WYXhwS2f9z88toTe0SJ4R/ZAAwN+No4Jnr
1oTDcDjBF91Li/gWaQKIpKZgrLW6MRK/4erAq365eMY8DZktVLSpwI3mo+TF
Zzt22IdEJW0jn0g3AcJaiqY0UsizWNRNxZhp70XH5lR1R/hnIt+GHbo0ZyCd
KTH6+z6DsIjG4qQ0DcCP1mA6Ho9OoM59f97t1Z67/h7g0dixEGn3gKQvZvJ+
0dG8Vw0qOSY2cKf8cQIPq4YMLvY60H2iB65fH7Ro/GpG4HXn9YCJ11jubvS8
5fV9ao1+nwFmjXbAHsW4yxCOKteGo8tN6QpLSspmCYimFWSRdXrt4S1jjx1i
20Sgah3uZYDK2+idgvKExmX0mRsHuRXfIVBBQBiM/a98VYp66uYNBylWFPwv
D1Y7tgFiUyo8ZVf0KJ3p6Ef3peun1kiMatWooAMebQQb1EfuiJ7djh3mG79H
edFm0m9gPHxCAoVrFyLNhdcXqQ6umOtx3GHarEtAHC12t+pepu2yijxcRfld
24hhsq3NmxpCPRu6C3PZ+zb7RTArAqWQ3SOKIpCQr0K76jBjzGHzVTQ9Ukng
nW/dhAfidZ5g1uCrSkNOq271muzkRYiiSJRFlhw79Qe0n8lZArKtrx39njdx
/YNnwcPuzqwtrLoq1Qvxf1Rd3j8V7C9UtJEa8wKXIdzzCb1+3hZ3uJ7c7LEf
H7nTMlIncbBn14W4F0aq7kYIcO3WSW6oTD1WbdmZzV50kF9s4bjWMq9+wa3A
1omQyQczfpsU/RRTMNVKVE7JehHaIpCP3Nr/Xtr0RhXw3x1nUppeVChgm2WS
/pBKyihplDZVZyx+0Ea+FKX3Z46ps5vWcBoiJmcWPQ0b1Qb15+9LJ/EpWX9d
w/5AdilEyoHBnLByyLL7WEcZ0uhsbd9KaI7ArHzWaxsIx8aXLifXbMg0Zhqp
HZRxEva7YIoaYOfN1+tU6AryADaQcJPjsY6lFhU1/1umtVAEnPrkYG4PKJMe
UhJC8e+yTziSAZzrb0P0z/QGI15UOsm9USs6HZ2VhvqFtLcYzz93DNWcBRYZ
/sOuVabdR+JgdvoXaKB46kBf6nQuQJEyUYUwDQUSUO3pAXtiVo+sQjF9aCMl
DmvETuP48DrS+f4zjh+si9qo5+PitpT2/2/1nRk2O9ZQAkgHR9AfvS/c7Zrw
fc4ZJuJAUSKJ2Hc+wx5i+60SIe/IkrX0PS4CW83ur+6vpc0c5nM70B8SBRFQ
jzU7QZEJDy2QV/eUg5N5PoN+yQ580RN1ZY8orEDHWTAqYxOlDSiu5qwIw4aj
5pRwRmya0XKrZeS/Noh/84gj2AxzrmVCKt7c6MeWfGGTeW4nNVXn9sf5ymXZ
9nlFbqFkHKk95DS5JL6sg5xhV2XujbW5Z/bMSLnlBB0UrWnx2QrXmEXgykFi
yjJqhwq3DX9X9nI2KDgVukJhZ1dMtyl7cD3ABtcyyGLC9NOao5brI26kyFtV
1U5LdzFpkjhOQNdoDDhmIV/ZqVz8Z85N+QY1TXR1C+OQe2tKn1cg72bt5Nmc
L62M6lOkWTbSgDHVyYvJLUT4ShUipZASKHpbSBHchlKm+hv5U9UNvtPC3qBh
8Vz0SaljUVjAzC76i0HLZP/uVnj+Z67u3pFDDIDRr+PLHGS+OnNB1GHRHE12
PAmveE81aqxmGahEntA6UkztoEP5S2KIebECDKveUn2TeHntOda4Gqejs2Gl
KedQDpCnuvB1EzW5yebr2D2wLybX0nLWMEbfB+knzJqEtekzbM1UpVOykTAy
T6kuOBzD7O6wdZ1p6ygSaQ95uYakr43lsx+yvfpaILZNeyDgh6G6MktdLCzY
DT1SQgDJWPcjfEj62hIQrbrYFE2FVt3FeUdHJo/7KWqznam7LFqoTT/Gw5hx
0M9/L+0AzAM/W93dOMLcG0N+IlXJYxZSTMRtY+eHZhqpTh/tf6ri4NF+r0fB
BwxWuoI/+kghwByaK8MeHscYcQ+XnK60MkN/RjBLky/Lb2edBMQVtKXbfWrs
kQys6ZeviJdKO+Tgcf6fkKKUUa72VC+fsLITSXM0gneoNz5ihFLHTD/nIr1E
2AR3QeYy5ZQgSOzIorLeNlJN3LA/jc6OpfdKd7cfPbnOOBeM6bkR4HfXNWyb
FLgtUk8EfetAhaH4Ew53qUR9IqWqnzwrNEgqMebCpL9SJ+cfYFB213RKhFWl
1iGZ5vcMFd5F0TNpDrSJwK/Cvwqm/t56j2XuhvurOqN4mQLE/W0eOQuO76ol
3WfEh9vQY7t4JS+iIhHCnREuf0KSKMmM9RHuRWK0novVnYNmT8ePe+YlZ3PX
wx3kkbbaduJndnxygR0iC5SosjhtRPH62udh12GfZIr1BoinIlTFYov6/Obc
BcjhVUliVDxgVMrUPtlNWoLribtaa2KTd+/GxEKfinp9a+mHDERNS2rFatVl
cS8H6IaM8GdFIxHqN7Jp1YR3uOB+jOlFjdPRqcmirbF2oev1mUXAsgNfj/YY
jwchveiy029pBjPJMRRbU/SJ9gv5KXgyWALWloLwkwGIhN/ynBOHvIN+HDXn
x2o2EuSZ3Y5SgkVf393cCzZU+K4RCU+JY9uw2E9Eg/SRrieHDd6fPi1slk19
NwTduZoU/blz56HVRPiFC8zJYrBbyz46O+n5LXYn6d0gpNbgllBFYAqdmT2h
hrSyBElWHn2L/qOfSyvHXgAhuOZpVvK0lh48K9RARllUL6gkADuiLcmrfdgh
pIriyXG90RWiHcwGsqUrpE6wrubRx4eMmL567WNmiM0WGmKyyHnPm/g6VG+q
9WaxsqJ8EJyjTc7ftXUYc+4ENH6kdOnSTDdctqfvED0P3hQVReyhpTHNBH2/
EqsnLpv89tVYTIKD2AJ55DjmJsAWdm91EdsSwOURMty/dDkH8lUAWRVvDv0I
jaeLVu08FYfUJhM0oYalGzihL4w44A/0/DBuUhmFIed6kZoIzHOYpHgKHfG7
vmMDOu0pdRGQKXdadGxO9gt0eRqMDdWPzaOK/ygUAKfT4DVOjeqx4dpJR4KJ
YEXfBoJadBKYhFFjLmFRs1DHWNNt7VFEvd8640v/lPgDWiYaO5juZGuNKQAO
2hnBJiou6p3OF8Js6gm8b0B7cIVhKGwYqeHZQT7e39T8oltccodKkk5KQD24
Xry2fR7Ximg5DxILcahLIYB/5Hea1r+v9GOIdT22/F8Kwjmb/8FTFkgg4ShO
6M63dOJ3bxN6iDDRtSe4TLNXTbvmwWcA0b2A/e2Hl1tICLPvwtXdM/rZf+Zg
SwF2nLt3pRL8jc/uY9iMtgRyGE0ZqmxtANcE+veVZkKB+/3XWCIEP1FCWAiO
rq8zue4rb9BZlqTdEAFfX6rZOtvisWj9IShgbJPZRLt+a/fI6mjQYnzLfdcR
am+tsDwyvv0dEZRLUX5JNlHMPpG4fpXb+F50hYbirCFMv3HYcV+ekHRfIxdT
8cfAIF1Fec5K1DLJ6IX4P8kA5atlkawO5+glt79XH2NQ9XPWNKJlwNG6Pwag
o6IkruY1uhYNuWmGzcpuBx9ZlPbI68MazjFAE49o9kfIGyZ8PlDv/Z8hSg0n
nFeu4321OEaptaT+rBIitwHrEbycAG6GFgr7Kj0uMqXKtEcgGrAkVFfXJ63+
sMOfoI05X9T2GsEuoP4h8ioaaJrRAHuHa3nr1SoZglmNzUMHMR2VeG+WXswg
dPnwzW81wW8IGHymNKWO2NEr2lpBTGlF4n1nXd7TAaMKcMYVMGNp+i+6XM5B
/jn5CUeHbefzneyoqdCYvqKISeSPnBfrLPh0xIVb41LK2qgsrgD7GHxQYecJ
usPltqFuk2YedR81NZ/zOJi8XcleoJdcYsMTQ+3e/ABK9ibaBBJiKaPQQlfl
CGNuX3lI2faRBKYi4hGulerWPOz82uiI/y0uSTj+azLsAF0sGO68ef6xeasN
l50GzZMRmdTmKJkzu2RhMbxO8/YKPW2hJ3pW4Ntnitz/YDmsSek7usUMvzmb
zYkHCALvX4QwaNXwxcgDrRCfk2VEeuzK2+4E/ubnUCe3KSRQiKyPeqz2cslI
gy8AV5/aN7zacJBECUWaAuGTJkWu5lnN52930wZ3oniAjvV6lsNX/1OqEZNh
lSKBs/btm/qYbfqsr9yOdMpTDo0hpg8OspYHDlLLqcGVPZ63ow7dU/fQ3HTJ
RX8r+/1hveQHiBqbVMd45CtczwfwivtPXpBDQvEX7f9LSTN8/P6PhhTUGFN/
KbJHu3Ko0z2BKIfQCzXqIMq/rBq8808Uf2rDmYxhiGeFYty++02eiVQQmpR9
2X+pnsuCR/34/YDUn3Ztxk1wrHEI3jQrjkVUcOpVULuko27ws9M8YjtNQHIv
oQ6v2EDGmAPl6GfMxKTJwtq53SRDtgAtIk99dwvJ/C4U4rjNFlb1XCGrMWG0
bOVNHdRO0wN62RpZIXWdHvU2WDtxblBrLA6f1liIkrbF2WVhKsCaEeqVZH3g
rtsfCty5OI7WHDTwRZBeUBVs9sKF6p2GN5xisRgpe/bCnYrsq4vNKQt9Xg1R
TFDW+BQHsGuHF0dZy4+A+Fw+UjKUj90iaPGkH+uFTtA0iDmMLg4+Y7Mu97hl
/pDSHesuPh5NbqYBtQjYyJq4KGHlXM5SlcgrwS0bHFF2XKGLcfY0nRfPNczY
8XPbkvnAgJAXD9qx8N0vQsPkYJG2rwLjw4DhLxH7hHQ0lPJ3OOG8XZNL4xxi
YUr2gwCfSrf4bdF/1BhhVpMjAOo6UyKp61yx24mAQHmkLqUKBNC8L7ZN2spT
HP9Ckv+XgAqbzHfzvdHWehk5ObG8QIPEJxWldoeA+dGFHSKzcheQd3XGzeDW
rNeeZENonh6bYNraa2XeOPqBYQxe37UB14JDimHgEQgsrhqfFmj+2zX4j5px
XmQMcK1aZG4zXjCADkU2Sqxovi2cQM2Kex3N2ZWAF32OquGPD2/W8Wt5NopI
jYLj6pSikgLEBQwEmQobLPpvV0AX2xMyruF8nijpP9cTqogd4EF4+0CVvjvO
vYwNy5iCnu8qVuwuVdgeVx6fFi59Ila32EEcPshA65KWuKEOy+Yb7Y0MK84j
Q6umGNYnVuUhTBMrQZAGcNV+zawwumMXdtboQ4Eixv7YUu8HdTepDFUPU+Ik
ISYMK/bNVZkke+llS+kY1RjCTiM09JJgTDJlGzem/Z5iEn5McIW3QDYfJxI/
l+v8HKUfCn847/u1z6u65yLvcl/VCChA1nEeVY65ZhjZyOjwPQ+Ks2qldpxW
2ULI5Zax9qQvj1xlx5JnXBV0QSLHXfSg5HQK9Q0bYOoYAezIH2JntyCoUycH
uTgjiBOufBzCbZSOad7NvAaevNzLVF1O5ymnJ96jJ0+vwBEPmbF1aO/9hYkV
lQUUYEY0W9wmosD0+UwTRWCfozafaD+c9I1aQ7VZqbwVm7s1mxao2MIc2nI0
D433/cQCeDDy6iOFXMPS//zR2d07vWwq0iHBkVjn7VxtW4UI6VDSQUhLnT9v
ajIOCGMxWiIYhWfKeHApmeI+TPgTO3+MOmqCi060p6t3qnXvk4xk5v0G45fh
Wtaub3cqHROa60iXYUvqyiNc0kk9w4hDBeoTDPzYpR43/dNr7CvUJA/MAgrW
cAZQKGY/maD4kYoxCaMMWCWzU4oKR+6+4s6FJt0R9ltgYezgxdX8yrEsRO4w
AqExdkg21NcvuI7RDb8BFaPF6HwPhq6VW1bT4j63cZejxsApg6GXa5WV/wKw
FN1uGTW9oRHPCpleSlAHA6JrOXjgOHr5GS5NxgE9RUXReArL1S2sQFGfCRJ8
dyuC2w7wxdUNXe5l7ZjzY9z0NT4t/wcwwoW11bsO/rUOw43KZs00rpM2Q3xy
yllYJoTp7/Uinyi8I2f66dC2no7tpJ+E7C5TTONXChRZOoJD5TisXSSZ2VTM
Dw09qdaDn0xqtQnaQ7go0iHwOlEsKQgcIJl5ZU2eLRox72PUJFe/gqY+W/WB
HlWA7ru6/Lcm6tsqH/gePOPr3P2bMzCWjIlCuFJjmQBZ6ukvoEZjMu1rDx+s
JekeJaRjlQ7JrMNeMPi9bslt2qQRdtQXuVWlUA/QSyNDk8uQCLT54vluTkpW
Vpox57uPQkC0mveMS9cWcHuwuoB8hTqvQm2w/PxayNTGWWkyFcClz4SCahnZ
znFWIFXYJaKzkF2cUQZXqEzdBG6FKcK8+2zBA/4PQsg7UVIW5V8AHjRiO07p
cQMS3DJtHFsy9++mc+/qKtLI/NeQ0Vs7+S051hMcxb6V7p6bQcfR08hgEUu4
hnD6bKX2oMG29oOmyHZ70OPm5EjOn1J1JBWErIIURZcTSybnC0tnMm9UHpuL
+mPN6NXbM6Jen1AaglhIaVTqVhRuK9gzzhgEua3V/7a6wSYhjW4F7Vgy2dyD
gHNlFIq3GwipSoUR1XwcqJQiSAIbjjyEi9ghZiMXHP8mu2Lcj5KAYpaPqzeY
BPIHald3q15njnqN7zif0geR6jolkuK9VYZSt/+fusSxH5UncT+Yd5K1qHnk
n/OoXDD6Kyd4XAmDqqaSj+TqUIyV5tiUVbpWi4prDAuBUm/iTDjsaYQmuB8Z
uh3rVNRdiLBTwReo2DCcvBZTZZIRPwPpN9GwWqBXLUA58mr6p3aDmLlbstDT
ijNk+7S+LVKA7xMMO2+b/WrN/yx/4joLYME6JfmGAjQawi3cirOwQjtseweI
z5YJfA6nhyEKasI824BoH3La3txB3ZNjMP1nkM6FPz3x7YApSlhwzklnUWl9
e7+4Xx88VR3ncB4rvVNRGV+X/z5kfTLL4uXqhEbfTFosmlMeGPGlnHFRPQxw
O0DBEnSmi5Ysqfq197OPRmE0Ov1BWKq5ZiwSc287z8Ev9/i26swwtuUGw3Dr
y3nrgd/+g1XcG/n8mNtDKjDxGRHIvKHjGuYSVKMp2GXgTmKELyBi5DQrE0g1
ZPOzIfe+N+Hn0P2Jlw9di7QxCQi2u9lp8BJfv4wl3ByzX1ztw/Nw+fZyhxp6
bqOnZhWTfCiiMftDuhJmCpMVm5EDiI/B75BjCdc9b/VSc8F8QzivkTku0Ue/
2zj5Hj4Cd3QWUdsqbuP4HuTkDBAIPylTj4lI8VWRplLBtoyjtm3/LLwEa4rs
3qkHjRcgBWhavBBz+88/Z35QAEP17SdhXhwgEsoVsgW7yTIPXXPNmZzyMhZa
4grT9goo3dArzA0PvHwt0GXjw3VfcJMvqsL6X2ulQnoZY3recukbhMw6Cp0V
T5T0fbgMwaNOcEH9WlortCoLmuULJuWDaC80u3BczbbK11qKoceMcSFOlOQq
luuMXZQHjFGOEoRwoPKAO8MdR2MrF2UtY2duzaBK6YR9irc9n4LXWiFsqRwm
QdQsjus4x2dqxeDb56X8NxDF1+xaqN6aQmTFOG83uEjFIGfJGreuT6LgFcEu
NjjSpIFDiOgxuQIDJlHHfPUKcoYMuLtddXsNKqLD+30R+N+saAvFu7C987sC
rCcRbnQWl7kLrg5h8S9ztU+hH2cqJR+rZ8MsD49ceCtkrSOQehnXKZ4icV2V
PLMnJzBRduwqEZ+srZgNvlBksyy0kCMw6PdMV/2228gvaRYj0HZ+8tlEgAmZ
c6FxnGZFy+QHl1iTUVDxhSEkee4PZqug+oPDPw9pgtbNDM64wiTrbc6LiUwD
YUDU7pVJi6YlXJER+xgaTSpfNxblqw8Zn+Pa+6t6i6pd91HYvttSGMGRlKxs
/fnaR/o/v4gA3hVe71KftfYkf8o3it1E5lRHhpXvpLv7PsqX0Bdncrukp/BR
BlvXElFmIH1kft9tHT+fjSJ1mEfxFJ47ZsyFFs19IUY/aWbZqwHojmYHs97S
GSJnx7rkXOYPYJq9YTDZ1Wh08HbsePtnn7ks6jx8UpHUfSScmVqpMItzbGJ4
gHgh/a6E9wPffiCSZeOP8Vmkq5sEbS1btLzOuuykVUi4n0POsGltyoSxl0tk
89qK9LYImP8B3AbwGniRO4RMBsBE7CsJabntiWQrfiLQb6Rl86wDpZpJqkL6
mp/U7Jyoar0jwD5WSbfnzSFL6oz5FErIZ4krIOp46EpyTFeoGVWU0HfaiSJy
t92SVOKbJhCadK+NckSdsiBOXIRS686o7fSDQgv7zUGphuq4exrjb+Yj23tV
Ml5tm6KOpGky78EVC0UAEBVdc6dk54+nrbBA4zluJBY1JV838E3H6XOd9eMO
Z2ka3r6B9Hbj0esfSTbh/tP3Nv50PuM0wKXE0gcibow7YVNGYV4Obuaaxcar
HUDqdf7bd9d48TJ2EUdYoiFpzVsYomVfAww301HyNcYhupehpp4PJ5sfZ2fe
wOVR2dpU8WdwhwoID7V+AgaRNy2Iag2Tdvnpy8fWlByABeAVJIAr+ADxXEY/
g/KgAyE8W9JVX2nttD6KcO+ZUjEM/9Wk4xyYovN7BDQgcZwHZRWC3H83Fwff
NEY5rL9xljOoxrgJCY7rw5/sNFOQ0PuxHWMwCbdNFCyBfOzFIHIU3BQ2Vuoq
novpHSzzcSB7QDNW1k4WotZwVQjI3wfYaIDzllGVk5O5L+8CwoIbuNC0egMH
09+jBeV7p7ZPjb9F3PfdDG/RKxOXVdxKnoIChRxLFhhZN25BIy3uax2XQHYl
44Lo2IlstYIuG2rIVEnlX7KUvVYFvXnp4WvLuTCWQ+3VyxUa6ChjlYGtL/1K
iMhH78zr6mgHII0IPb0txqU/lEVhZ/HjSr+eLQdw/Hj39SYKpW9few+BIiyw
hF+QzCjliKlKwWcfr+iEYLhlNa6mYMAy8gWfqOAQKgRQLwQKpz+zzDKl5/i1
weRnQcvLw3MCWYbaptOsyuSUrMhLuYJVPq0BeZQTQ/3TlbHEzm3FmpWYifpZ
3FV+4SZ9x5hBUuaKOnmJIQo4lynNa2m3WypEIUlZnCg8apLk2bqyljCsJguW
NJtPXa8GU3opDYSMYf5WRPV51iLrf5XMHDukyhAuulHXpNafxaQ0D+p5WpPc
pZVTdmpeuj7O5+HyG3XGYOIP55caRgAvnzvLagNRbAqZnf52DbJxPqxnoO5i
gkyBH8Gjt2yZ546/G5baa1rPiTG9eS8mJkegZd1FJ0aV7ep4tIND+JOh8Tt1
ow/xHSrCbjkkIx4FVIIHGdT7PzQ2JS+kVsUhaCWpd1YooKL+AVp9AGGNH7JQ
Qb7a16yCL1Tyc3cT82HwgahI8rQB8fUngo6tmtYtv0lMlPK/O+TcIo8ziOfW
t6PcTiTnGQXnLUeEHLkODvBRWBTHq+bCLQCoP6KOxF/ABYtfx0TOQFdEZ6/5
Yg5H39Nx4OlfrrXftanycnc+VvRrqJjMbG/wMso3G7Yrm9vQcHQC5LbFzS+c
neFT/Z9/cvZ+C9h5uC3A1V5jd28O44aaHXuc1O2MD/Kl+pqxSxTzkJhHPvTu
02Efv7zbmZZ0PHctQ1+Igm8RaAk8mCSOYsIGSx4C/0FaFnjJ5Kubni0Vow8w
WMVpyGGtdx7xKNH85iHqgYOcY27zTQpjtM9poVpJ932CGlypFeFDu84AHDtX
l8U7byZdwyY65E0ZLkbONssGRsVvp2RpykPCzLqUp0Fef5qHyjUiMKlNyqsR
kej8itPQB8SVocWAjtiC6SYd34fFUPHIo7DsylZsZFCuy08JPkUwwVKv4/f5
gIL94elQWyccuutPcuml8FPCU1rhe4mQEKXtVEVkYeXR/KBDklUw/9ZLx0uj
7XuTUXAOZh01ET8Q39CIcDWNCBolKJXsMN3wuvIAzHt5/i1SbSzNV93qLYi3
0iCJ+NhVuuWvHLqUpGnBsLCiyUQEd6lAZLDWnFl0cQRpUowKs18n/9Lg/O0N
RslEtBKXbf0/KtlX6gKY5U7UngQTRzqCl7+m85eeFVGrFk6t7Vs+yUfCBIUK
o/zQgUdU+CWmJaODQazu1Ow9IbSIvmmn8jyv+bOWp0k9HBL9mG3DHIvwRyth
slJNulSlGf5L1FTJUdwpG4F5WgTiowjLvntcWdKRcG1SBfudCU16U/X6MKbQ
HKWO1OSEEkBEGv3kuLBdoNz+OG6ZzhRliGnndfzpFGJ2ltrwsvHFva/vRhS2
zSgXw9EL0RxT+XNfDgqswtBUaSNApYrJ8ZXgduRPexLmde7q1PwjnvatlVi0
hGDd4XOhvp1XD5R5URjLSjGtXOtfrk5W6pPImcsMtcWKzbfwx18f/FuuXHqz
U9qVQV4OOXdB+bYF5Ez6T6UxWmQwCYJS66EA03v0pQfFlNfZtIvbwHInYjLR
jqn8WGM25i98AyYEWsP4a86mwZQF6y2Q3fjO16JCdTOFBcHpNctRDhO6YMCN
jvFbuX4OHU50n3PcsSRLol95A/MCcQrSaEnT/yApRnvgkIVtVE/uwprvf35O
JZuZANyGeO9c7LjLxY0k9tlRod2a/ukI0OUe/iVlwETSjcRIzLhcIykzamn6
T6m6I4Irlg5VT1xdOC6GTZRJBu2EU+AVlmO6Fkn/QirKRx2tGCgnsGHAapnB
nDIE/RUhmmJH9JCxmBMeEg8oZEACpzfa//CJq5npN/sec5m4FMmNIG7nRLrn
QPv8UTjlhZ5j+bSWqip7G0E0LMqGpwQie4bK9NMscP9n1aBzRmFOH8YxxPGj
hD6p4wEoG3g0/ido/xqK4p34uOB/ewk4555Yf+kC/vv2SvU2QxehrxDuNjda
5rWf2olx2YPLx15C9/4iVC/6B6+5yQlkySljk13BcxzudfM43ead2SFbO0V+
chhjRWGkP+Kartp+VUIe+ls5kJ1QaoaBQo1QcERs+GzO9vmLsmKIkp6auPA8
cwhqX2J25tC+fsIAlGte7l7fzwqdkBWb7TIFGSj11hRWz6KDLbdkTWUm6gPe
9OROLD3R5tcyWt7YhRl9CbAW0JI+ZIqfp2mmWSuSwBGMP/CTwJtOjsuMDvl8
8jCcRPMfDnVGyCi0HsxWn0WxXF6w2iUCsOVauMLAFuzvBbDGX2iigMlFT6lR
QLkZI3+4fW1kinxazWN2VHpflY/nUY2rKN+QcstlS0iv3KI5emDw0oiAx08e
t8CpbCOK2OkRrhrJW3/zcNMsB0/O3qa/SKpQ1eAvxh6OxKzhhPVFsRHwfIHB
ELYaD5cEzx+GibU+6ee0YMCeUYa82oH92GLvMXwR0QWb1NZVcCDAPNFC4527
MmAQSIk38MhuTWArTUjmL6/uHecCh4jOsIYP5PP9sMhNNymyxfgs8M4DF/A1
ej1eRGiEapaC3bfMApCSyfXsoqUSsHx9b2Odhf/a8201n9Ehvlj0k+CtVwPL
0lnkXje0jLjSTX1Yjzdg7dJ1ue8CoOuQW4IlkM+CIqnfsrZAe0Cyq5JrHNlz
GY5PFygq3RYb0olutzFU15sZLjB1g7srhOzdTe3SX5N4Vye1KFr1tz6bMNma
woLK1UYdiw76sOtLW869lEXdjgPLGcp0XfIsc/d3SDGYpyLJa/jdgt7uC0vB
y5o9smjTCKjyaZWgZpwtbbprUdOqSXZjTAuzgb3IZKWN25a/RZ9sd8nGDEP9
N6r/1ucXoJUdY2gFM3PdGFU4TD9PqwUb2D5r1qjTl2ANuNFbVEdlIk1UruYq
YMZN7Oak1FOVeHMi/zHJV83QKQNFM1v4hWkig/oh1FRo0qCtB+Rw0u6eo5GV
m7bKaKJfnH6xCoqoQelK4W3iYGlIEZSQ2B2CkQdVTcYYm2CrXtgps8/uLnv2
EiELzAg/rdGHafP/mAGLZtUpoNaDGTkNkr/PTuRmcgunt9sQnc2htoP/7TkI
B2JBXf7TqSqcw2ZTiu4y6kmYtPnNgAjUofoVI7DawzBftTQNc/PoNK+X4eks
z3+oie8AFrisFotT5LgBaY/czwBaRAO4/hQYUCeAlpPTUtMfKgViToTF/u9x
cSHXURVejRfWbamAP6RvaG7nui0ALxGaCHXlo9GDEt1tsQHw+v3bvdPAsV5o
Z04uMSfTm66GqNLbc17g32DQf7MAtrHDZ5+nHDhgbSx/sCPNz+wmpbPiCwAi
fZrYM4tDFyWU4U46xMBjQGgwu28PU9UCC2xAu55uZdeQXgeCH45fpKfhlooc
jpF5r9Qca2GdZtjSyXCiJ7mlCYnFrsNYwbzq74VPieHrftIphhdmRGOxM9Ij
YIQQyL/P/bfxDd+KcPB+noCIt2lTa2ZOd3nRRMlYQufblqJRKo7nAdxpKCG3
gefrBoJ4IkOUMbY+fy/18raBow8MqNsiEbrngWLJ+RvA+dBLru1KC9fLnflB
WwmPgQh7Iy0+XhDf2UjEbvDU0/VheT5HTg5RJ/HBv/UYu8fLbsLNEWk6c6Y8
qgcr/Vcdf2oG/CNiAIMZv9b6AoTYj8kJ6PaIpaCZRqRsDMG/LlQs1FmfcKMF
EHWHRmgl0j2zChejgCRbE9cCL/I72K781jcZ959lHzsSwLOLp3+BZ0Zi6kc8
B+z81MlDiJfh83wJTayPuXLWNNJgYaucD1bQEht6n554logMErimCVezXsdb
YFZ5K9zgtDp2tHGzvZgHEF/kVmwDhm4nI8BszqHCwy5M2StJeJYg8U+sqUhR
6okpiOg4eA3fLOtAmsgX0jcoP3FTTcogOkSoVjxAJ2FU0jgw0Z6tyEa7q8fS
XkcQiZXtEE9yZff3hfw1lbrprwJr3vpTk9/7X4HcP15jOG7Quxidx6HlhR4h
MsYwRvXinRSNyZsMvsYi7/Y2kzGxu1yMXpgdmtXwd6kHCXMpbZGkicIgFrEr
F9oA2fsDzUFuPjnUV4vX6n+MMSSftoePnZ7U3qOWa9ObIf7AgkLYT5i89tfO
TAG+graaVZ3y3veInvhfBYml9arJo+xHb4pUq4LA8NOx/mI7QJ9iAQMzhWT8
OZIX9ZVltwtCtwb5uSSVWEjI3lSqMZjOaMO2adMKn/1Gh2nN2EocOAFZSg4r
jITr1plBSJ8WyMHF3QtGCSUgeqyDZgxa/MNDTl6/Pe1US5dg2CMXYm5A/FBf
rU7wGmc6SrPthOIR+cK/oTgzMmeyB+mi4vjgjf5VoKOZm1CnnRZkRh6e1qI9
GVuMgisk/KZZfRyuIk6M2KRv2hagFRTPbBhZUrnJBArP7Hff3HdDYKIIR6rS
yG7kjL7i9+uCQ41KyPNUjwXLvU8IvrUGDiAr0NKrCvBD/Rrh59kA7NoXf0Ob
W9nFzs97ahdnjWdEls55Ep4Ne6h1/z3PYG0kCNIiee1kSylCvscxvMDFV/ol
iY35K/n1hkywh2jm/a+6O8lT4lIJ1uq3Zgfwm2NKBKohWImDIbdFiuYg9Rn8
m/hBH6zcrDqcW/KbWYblcdXV5hwYBBvA7cJWTMAD9p0D4pmTX8FN2My79hpg
tIr6ZPD0yFFS0pACAMRdnCgviSBo0/+WDQ6yLdhuWX8Wy6u4TH5lCTD3Rlcq
beOJ2TdlqXkQXVYrt3Gp2DDM7OOGGslnUrc/Z1LDF6x9nQ52ldSNwlTaxo6E
vsfGQXkQ2m6wW8cKNjtuMq7EKDeX9MrQhDG1gGEy0AvFJegdfY64OW0baNTK
6ZHOM8Vvk+IeNEY/Gza75gx8I4sMoA4a3t3V5VrtOAk+8PKDbKD43z+rMj/5
emj2CoKr/AIlNcyUaV1fSN8R4mRx/N70v9NFqRcuFeNPf5QjOZ1L14f/LMUO
+7slBjQsuQ6nBO+uUEV0FzD6v1cUmWoZCFTiScPNKhP1sGwlipjk8Moq4RKn
oGUjFrSF3YL7LlDn5UGcOUUgi/WSWPWTjVS3azF9cAbkncmMyxX8qVx+X+0h
SPP1Tkabb8BoIJwNN2U0f2Kd7S/gBMJiZfHTTeHYOWrlqX5jW2Fz6YKFIgyp
NYb3gG7gXRPZU9ONFNvWAJxnu6R1MV8LeAR5gOmhdXp4jHL0xlX1LUYCWN/s
fDKq67tii43mmXXrPeXNLxwhG+73eWAhFeeZh229upezrhnY78sMQ0/5KG8F
TtFlxV8iDjo96qR8mqmIaAqTKtdcu2YzAC+dMmaE2fTLWVjuFHdy2DCWkbrC
n8PXhRNw9CCgXLcPhHLlber8nh5/25aLR3udqhtymBbn87PGM6/OGdi2CLcU
UsUh9Zh8Zj+LIQqMkCYtL8aTM0xFzlqF4vErftMArn1+cF/5DUeyAEFwNEOS
wTOo5uQSDl8u99DGlHHCdZT3CK5642AzePinl741CcEz/faY3mw+i6GbM5c7
nFll/WhlXzR1980eY4C6hkbrEK6CX+sq5/3lofl5eUAJRFhF4rMVRxag7WOs
c6ZF6Fu0tjeymlK7WEepaOCUHeNB2o0fy4HuiOnDTNrx9bON3WTFIePxSuRo
QP6o/Pb9QyF7S/mIHaJ2uK4crtbCSaHKDvanoMLrA6uwJ+mqlcqN6MiHg8Hr
MmguVMHJ5Nhb60ACJRWdAaKkwF3oczd3Qczg0QK0ZSZOAeh3zrpd3s0bUo7U
vbRjL+vDWat1x/IROuZ0A8IbOiALMPmIIdZKQfkeh9pxSHQWG6u8zX4G7Hn2
jrEruIX2SEILNoM0ewK74uGs0+7s/qZkRnvy4kVXmQ+bLLBC3RC1xAO85BLQ
ZvC8b8qPacQs4mKAOWupAEcxINoV/siQzSKmerKNRt94U1h4q/SOVNZ30Do8
D6f8118+YhCCr0Na59jgD4kjqVhBgXy9H3s2ihaL+Z2Tr+lwERbH9EwgBL1G
YkjY8JYDxIuxg+8946a792AllFtEIfz2Uh6P2eRld+g87kOjn1LNI5Jl6ym6
3yXy+IHFcfBjA/kMwnmC8O8BbJogLSB9SbY16XC2P7ifxrKz139n1JjNOaDh
Z8RTsNdP0CevyiGDLK4A8o8Onlp7zACJBQ2Wk4BF4R+KOPOOtr/mXj7d+Dep
oTQgfudrOMKWR+xCOXGhFUnJ14toGSlzRK68IvmLdlyZxHvlcbOi68hntBtx
Yv6c53NkHaZjbkFzi5QFX7+Q3DD+DW6DeEfzEX4KZQXYfT+e1UjrrSg8C5Q3
oZTEB2O4hbbiyU7zGEPLVEl62ODBMU/iKDOOKtnE64rmGI1YzPnq7VChIWI7
PWUgHNsegQP8y+A4U1mvhrC1iSJh64PDmslAZQYq8WXRzZUf80Nxd4/a0mVN
IlJPURdg8hGXFP67iAn2gPX0hpKepnoM1Ur+KuIcm2R6zTC6zxF1D3vEXBn2
4kbXAwIUB/6cTNYT4lnDSnrHQM3lDm6MmNkigWhTGnjef4HK/9PHH34Y5UgK
j/siQJ4LKTmzBncyZ+8xwJkOKVqRh/tVV9e+saV1IZ9QCvijOLdNlEbXhsOm
NBk2gvkIwcSqTdfNyGHXGuYw9b/KApQhbFTbh9sQNDYWaaimnKvpQrEHH/4p
DdCwligEfeCuiVY2K+DvyE3VNuNuVbrPxixTq+v4bhgGQAZJEYGi/DEbLGEO
umBzE2mGvKE6usAVBMzaBfh+ubC5B8eRSDkfreOZIuXqHTL2tDkXx3TD1OXt
GbCVJQjVknT6iWL5vTtoObw4USewbnJm/qQe3tjRiZhKgPZdu2OzpNwzNYt2
ys7D2IJkHEMb8NEDLnyGkCFENGmhY2U8A0ofFT+viReni1YEb2ghaZE2kVEN
ZXW+Trunr7/L8UoL3nADpwsouHSvFLaNq0Izf0ewyfA9ahzC+X6KMDIaS2JL
00gmUvyQcB/bwU3U/TlEyEOAiawrUPUSInkdFjx6/mz57T+08QJ+YXo0wGlP
JUt8j96qzyv4zqJ1calcVnBj2zQ6HP48wXpOnizsM+OKSNj26kJXGX0u9AHZ
31GaLMusr2Jkih8FIWB1WICgq3kS3mpPdH9zWtSdD8IpQq8u2DUiq8EQgbDA
euIfJ9a0I0yei66S3eMgDphFNixfZP4uKov8FZkZLUIuDI4tFSivfvC7APrU
rk44qDwZ8mAdsL7EAZKXBqUkyEqDYXEZ7AcYxM71A3jwMXW2upJL9B7BAMv0
w22nwHC5l3J3XEsj+4l08te9Od3WHB7eix+JcjYNn9mtdZhbD1YjX/cNU1LU
22Udb2FOS+UI4+LJzJ41gFSh7qRhDslbY6FNVznuBJH55N43yrrjhimSfxpJ
H3wGgT+F1mA8UNbGswOF75Wx2V6eJDfrf6kePHlZ0MvfHhw7HRIMovg18e5s
vZqfLSx3fQJNFkwOGQ9XaQkZJYv2wXzX605cs3bSkvmjon24rPn1fwm5OgeM
df9ZptqBuddLzpAi5XwlAWDKqnWuPCDeU/OkP3J57TDGbaopcGkwhc+I18Z4
FOu1/oKS4HL0zJEmNBUk6pf1463isj7dVnkHj8f9jh4f0suMSv7jqAY4Hfkg
iZeUPBQ1bG1aHinJWLaI4Be7kD5qnugeuFOp9wszE5fIjikIOV5VEuPolQTN
J8kUbj2+WgbR+zHmikV7zWlW1REGzQDlRffN0BH/uKZtuxlhIieum93DXPw8
NreaaRB3MWMJ4ZKqlF1iB9VG9DCBy521F+u3D/lNJRaP4tFO3VWQ9mZGO1nG
cB/yGX7BCmiqWrZtkvpGb83MxiaJZWkQqdmZt0GPodrNqF1MgaI8/Tdn1bnN
9L843gjt861pXonxrLNLxvvKwXLhERMtr/1nxDTN3+AVWMslSfJx89oU9VTv
vmbW20I+RhHVs8xVn6Tb2FUCqC82B2AhQ6l88zeHKRRLtppdeuvV827oz35b
SppT/NyUTKqNsriMONyfU1wDCcViw+9xlCNPdIHeJRB3i3gmGUaCk5JQPx1J
ujgDlV0NzH/2wlN8PjkQmIBS4sIbS5CjjDoXiU/zqCaEG8Pp1qaBYi5CUMjJ
SDygi5Qn5cX4hXX4C6iutQvE8DqqGa/fYDB/MEJvHA61gUjFkwLbl2qtKt1j
8tfMqVIC5jivtTQM3iIgjU88aPtWFPReZv3Sk7WXumV9WmGiljbzyDY/ZdKy
KRIxlNUkh42Ub5T0kkrPRLQZBx9a7DfpHQ/cwflpeeQxqH6wAcqKp4D+yTib
LBtKAlfhZTNy02kZXpWR6sP0WzMCsAP0Mtd55ICbTM5S4jkeFGkMoRFMj5Qa
PD3kHFJLF4gnRjs98ufocXqobMQrwfhcmhmcLlNfZFA8E3rZMPjHWI3WgmtU
ENJVYnZ7dsbb1PRY759Mb8N3ygFUCTWwCTldI+qK/9+9EYBEjclYyzZGLRuT
1+FPxedew1Skc2/ukFTwcZGZbPyjKBO+Kopyc4S8sh0cBe3Jy9bj9XOYPD8z
RCOX5ssraq/meHcmdWXetKuM7eUnEqxS5nI2dDWEdfd0zrQznwLR68tbpZcc
huUOloTHx1g3YhiEmLyAOzymuScxpWpEFw02zsd2SW1nSQFCWTUkmVtt0gAh
9I0ytHxRaVIkW5y7Yc3qVthECVd4Vnv3+iNtUioBKlI3x2cV8ltFalasVHBj
MWOUC3shUtTbVkMYt5WfaBKdH7NgphBtRTNMQWjixxtXmrGIvUeURyptu05h
1JP+LblUfcPlxY24Z6jmDV49YC967XltqIGp4lKnKTrluqYIm5YQj1MSJBRc
SOgg7qVqmoDhACAVSFNDzom0bjJyUin+50X98sgcWW+dQk18bVR9D6Ke4lFm
49LSVbAbxQ6ZHW+N/Mlr+Y+5t6BCaJKc5+dKQhkNdSwGM/MfxumWK4hvmBca
rpJDjoGx9AQMasTrMrjsusHKx2h13mexJeBZZPtWC0dZmvalm5Hy0iRHm6Gp
13BKTwgWc3/2/uEKl7Ga3Ys9Q3un5EvCoOCR2w3dzknlQMPZ1WEw3pg3nl45
WgXMlcpFk9e+RmYWEPGHKAf+6PwZT+iXQ2J39eLWYIk19Xk2gAK+GMUy+4j0
uin9H9phXMOCe9RBVu1dcexm3AnyU950pe18CLrLFXcXS/iS7Ub5TGNr3Yvc
9A6d2Ysb7I4tD0VAHBmziUVGrn2JrtSMH6D4gVdefEE+Kqlq2YvEam4NxIVx
O763f8NCgxoy2mW3JMwpugSdivqUPE2EqzBBTrVb/XO6kc552Xsiom9yWM+4
xDjLafF+hEScdQAGbS6D6ZMTpEEvOrKKSpQ0awqO07zXii838IOBgNrGElnL
WsmddaK7xPKxnIu8Au63O4ZKJ27V3M2DnvCdPkXaA5/trErhNw9IcHpMP3Qv
nOuycDkLM4zevzLwLLZ8luEAvRLHaiW9ziwpRDExD9TvYRaIFot1SQvwVhgX
PKPhp98z9vY9I44h07mdKYthEfCBwmSvAZ0wHPW9FOwVIqnxjYz0qzvsKhO2
eho2rZufrAMz7SzrXV9DBVu9TL0KZEV7lxQD+1O40psfun7+TVKPsIidbBjT
u4LuxP8uW//su7U1sjUzCUcL/R/efQYuqkZ/WoMkSRhxgLpuolf+lI4TUotE
yUOjwrI9ZYN8rqH44N2gz3Jm9sBODY/+AebEEaG70tsoSUPBfyP1DUiCUq5W
IyG7TzD3FVcbeeC9p2dW7BZXXs2JFeg0J2q1Hic8lOglh2Iegh07YH1nx7wP
1q3v7srODyeTKJZZ5H54LkcCtTu95/0BLvQer5NiLnZfhc48syCyJ0LT1zcx
ESgf81vTeWttCwmqlRMkKjs/NseZUdsfBK7qWYlAVJloFFiShFEWpHBU8cta
vCsCACMh1+wbfQyGDFHLk+AJdSqi6jEl8/DSzGw66qxRRwqprJsShMRtuFYt
emjpSgOBogMaMAJdq/V/p+df7B6VLOqQW5g5CEpYnU0kpnkfFiNFX5SiHazR
APgOBCoQg4eH296RqXav1G/Z2ZfWj6cqlM3R/TEG3phPmqnvoKvzvuksTZBM
QpTHYux2ARO//BR95KPjKxxzZjIf3cqcVTCbZTpiPIvIL/mFfgSO4klCxh07
r+Fs5OLZA5T8yS/1g5PsUgfHGJZKvZw5+wHu1YcbhAm9QH5afrvR2BXWN/R1
NvYaHrtBJOkgvj/4p5oOjznSurx/of8qp/ssuTMkpKFDssA1VsO8g02ANTaM
gtmA4+yZfg1LgIZ9eMZPyxytjHGWySmkupQ2EEW3ff7Kh6+EX0wfROBjtolL
GJzy1fMoVrVpeh6dyuwnyqwCA+5Bwgu3OmqhTVliVwN2Yyu6D0ZYGWNw3K1d
CzjnVMcW0LjPxb8Lyl5wZEdAzR4YBTaumJHEzcEtL2pxsFSM2fjuqU5RhdKN
w0VfrOVJ2KMBeDOLU9bLD7LNfo8EWfxCl3sOzzufPIFSNnt5jBwq0EhLSlDp
rY92MLH/sVqOzqZhemqPArEbKuiaPnHOlsJoZbD3BshRoiTTkQIcGdfAmXCN
YkojCf3osE7VqIrdi9xF5Exla1gy4Ifp8qvzTfYXAqlHnU2B/azcQI+0WFEg
2rc1hCblfm7T5kJCvPYvC7ERGt5SDp/R4pdaXJoSk6IWmJshZCGo1OxoeqG+
/ZUlZ00YC7WeDqGeuO4yOM7B8TqiV9lR0rxuyLHHEl/Y90gr8GtnOHSY9ajG
KSkRtwj7sLdVf2v4J4nEDGY1+wdon+Fu+t/boN6AhQCCNfAzCCuPOWHm/o4q
EySvwZ9HUR+X0MHtDnpSzrQOLlArgl3WrHIUviMeSdxR7zLMEHsQbRS/7lh0
tGkfRvtJUvoJYDp/ylsybzO0UZN/anWe5UGF0oANUTK0xe2Eyn4Z+z4Ia7Kq
ehjjuEE1Xd0gZsh1+OFU6ciZcwulOBRiyGSkxohNQhLTDTBpzH8OnasPonBv
aYzOmcs9L+idVIsW8idmr/l40Jg3PMp8vLq+UjQcELykejGFv/wBOPWyZhuR
h/1HyQYbcBYDXWD09b7fh34czrUWcFsRCgRJQ/X8b/Dj30TYwq4ms+z1LnV6
ylY8Zf416YKWhB3RJ7Mj4g6V+KL8zveo3SjadylKk0lN4ctme4IA0JZRFWAb
EHT/jjCm7kb1L/M/hRBtlDZeohX5DEAU8oYcYBnwjDEpDaPKJSUxpxvtCKWC
tlEBnLO0Pm4e1VIiq/7yfYe33tMF0lNVYlFY+6z8G8I9cbiJ8auWX0Hh0sT6
nVeDrHqMzUHXcm3J05Yglj/bIMQRd98nGRZClQhbJxJSwvL+ywklBNeFr0MW
jouCBN4wzDxnUB+PeGEEil46XFE8/vTWtfS+J0ZWvVsKI03kLthiLK/b5EKz
MuDmJPz2nsu3aIC4g3e1PsazWYGxaYV/L3N1eS2K5gvQvi9eygqEz6GULKZ6
MOF2DBDsHjSriQWFKS7cQf1vbC7R5dSjPMDuJ+WKcKuOKUKrOAZlH7BcwQFd
i/WApeg3PHcgA7S5jGeztBK62/Tj1D3RVKQgSuPcvuOfmdcr0OZ5lRGGXNCv
n58MQmgbNEOYkTBtCVqZ9YEpiUiD/V3x2znYnVujSBJpF7GB4vuKQP19HxFs
YdXE9Gg/DkcODINpZeOfjjP1ZGuzrl5vvVAAPp4lhVHuOuMBlFbGOrW3K6MP
PRm936aeJYq24axnk/P8lFYxer/b1WB0DCTaS+wg41vYitKG2H4Ln47GpwCN
TtDIFJx7KLWccby99+hUmOvRhUKsgJ+XCj0hPsVKu+yUgOL78ZM5tLYzwGB/
tIWmTfdeH4AisaDby/R+FiqTOUcQF+vWgUqjYGPYRPNzrQi4hHuEls+bbSMt
hbUXZY1jRDu7fkTs+SnFjYmRvxa/I303KCzBhuhPi09Np6ZbZqhkafBC3Zoj
GDB96ZgS+aJ8q3jT2hju/4SVKm28Z2YtKEA3ZRPYgTj5CMkudSVwGlMGaOYA
GNoOLrm2FUYiMVhxx4kQ5mkVh3m0eTomYUx2PaTr5MmsrsBlRANwZ1c9KCga
IFGS1eQ9ft8WuNVRh/k3Jlmmvqd+qtEz0fMsZFxSO7mayhBLzUkyANPjEXWr
FfcFlGYbf4hF5wAj7NvgFlEpQvrZu+/HS2nNfZAGPQL2EAvk3BSFovrHudUc
EHRrWUlxwDueMA2dFptfygCW3aRpRtZdxDQCBRtecC8XDz9kqonQLtcqKT2+
DWfN3cAyg2ulHPgepq5p7MYLondtdO6xm7cbr8jIhGXojkF+oKzzHKnA+joD
9cpZ5joHKSbySLzX0vM0C72iPPMtIwmnIIs61LUPF4qXv/nk/hRHj2thTZoK
M+CoZUk9DUjHcMNsBkkqEbt6MXwhduEeAXdXLCfdaXYsX2ByNvrJbLu+huTb
sZsujPhVkVa43VmITlzbbtrCFSfwuA8ffYungNGJD4Hmff7MQhESszNc9q1V
Z0OeZq/8qooLl/mYGJf5EeFEycWiOdcGdT29L3guAP8kJt1t4w90MjFwYqTq
U02fu/dwIp+jEq3Zg9wK8S5UUKhZ0DQ7x/4Dt7oelnTKPse9Orfn9nNup7rV
2JlOHiGXrJPhhPh/Txs9w4OeRur82pmk2TeaqR2EDVWGYB9sTu6ogJ4rUczp
kY6N5JPFQiNI4GbFwBo3GGudA0ne83RUtORrLnPqDVM8eGvWnC28KTV+kuxX
r0YsU0dD1YZBJ2vpiIIxKQybYjzZ15lbqCxZ1Q0yCoE55qK2MXoh0j6CqU0x
IcyLv7+sY5/vuvn4ch+k0rD45HbGi2l+kMMeY1KnYPY9eQ+/I8FZrwoge6tJ
Zr2tjGWs0r1j9bgmRuXcw9t74Q50xPQdmkehWCHhD5cW5di7cD+SLSXurWWC
z/GiEDldBVBiCNIQ9ZXJKw77ONrGFXJCEK/NB8LW9170okya9FcvVegQe2ZT
Vu/G59/SM8gbe/7qBF2maJtEKanYtxnfg9SWiuQDV+X6OgJEThGp/IMf4tae
QYtuC9jC1KOyLQlz670QqedqeXTVguqgdQEjhF5n1BT2A4AZFvIBGTXlNcm1
mL4Iv8nv3MnEVslq4sTzxErXDb7366Tgk07FWGAsvGwnMYhFmIKcLB24POIS
7Sc4PIc1gfcwQU+zVVw1VUGZW6NiHXmKJlTeT7OMo0noHF4GptDdkKJQ612I
Kw2BxicX9iT/t2CXpkSXCigJ0LurQbGg9dccoVm0EvaEe8jqguhVoyrf1Vg2
a/JCrChCg8akOrQiahI7DXx4TtCurX8axltr178b8dy/K3wwfp9SXcS5JzZ6
rUJEkPReqUIg65whlEBL774x9+N+kTKWTb9UIgFO79/HTzjIlfN9O1eE+D/s
2v6bSHo+FnQ+Op2WHxlzKz8/mkOIZ27Z4oYxRfz06E0PC1VvXL//Jpfn0Tf7
AAkoUHk73EuJjuPCAFynPENbt4kmkBjEdlTTMOeuwoKWRYBKuf4YSWmjab8i
/ycg09rdH+sW5IdTo84oYHvsNyJuNwoVB1M3gQJa8Gr0ZN5BQRxZ0UKO7XRp
pXbIHUJUc4ztlW/Z3UFAhqlArwmqVSmnPqVc057WRo2prG9IwWT9GnxWy5Cg
QV5PydBhOcxdakS1mcNTc4BMqVtY8Mfwx8H18idk87xHwy5uj5FFA/zMQxw8
bhxi9l32Kuy6VefsSHYzO+NBSfa2RyoywRcFCXCxEX8gGQkSdM33Bx0/TQDI
npSofYsYV/v8D78zYHE3llfBVfH6+SRraWuVzqSpYqGBbK+z/+8dg7svVrZQ
rfAXofcQ3f5CiTVDvxxectL6hVkKd3Ctjlulb+TL20tWOG3cl4NZ5NFVZtBO
b0+q4tMJFeXJc6LknNZAw0NjPTlwpHgTkbLUybYo7E4KCQkiozDcdD9GxzeD
g8knpHUj/NEHgliP3Kj9g+SIHTq0nP51DqHqk+kkFF1m1W43JV7EocVgW4qe
NQX6jRBQLryYvvVDBhadu5lpSWcm6F8z5F9INeS9vNqQAubK6WyLR5AmYu4O
kd8R9CsRWXKv050hBaIuyl75eFcDst3lEdsOJ0ymObvwGq3flmDET7kglf2P
O31YrChWPl2HPkw38tf13PxXhh/qZvK1q0bHBnDy/lBgxA/jnnsPNKZfPxIn
WiA5q2gxrIj4ABku+5YWLyYG5Ig5jGRtz1CPTivQnYk2roCMIH8fV+kvYaCP
I/s3KtrHsqqYmAzgBWMWFYnomBbuqYoENjhSV8DKQB9nx9u8FRcaxPpY50wD
mOukvUsYJDYJoPxuCAow+RPwFZ7ITS19jF1jhvYcdvic6pdR66LXQA6wDXN5
5th/d4PtVW9q5oDeAsTMl+7YrW9mRvIiU5EjX9LLqkvaZWAbMbYtyZ6ZNh1J
1TvgznnhUjVeXGYBGCtYBMwJdiwvUbtf1WRzG1p6iyB97b1aljcICQ8A+Lzn
Uvrk5HNtnh+7d7ln4YcjMr530XsxLZphAsO8EbytdhfdySofRsWSDn5kmgsR
chOwCwV7NsfpiwxRIhU59IxUF3ZmWIAtp5iJTkIpuHvX9TimxHMufd7G1513
rckbuxlPkZ/wfVqo5lesPUEC1uTn9OeznwRj6ZKHJKeUb35mEHlMQjcGlmGB
C/p5zKwT68NU/gxE6xuJrev5txOwLtZiBkfcgtpz2DbW3Q6iCNADKJGYur36
BAbtustM6zlj5TS0BDhB6zO1tP0lOzN6TBw/OJS/aXSPKXFbfXM8R2M4qMcB
6sL67uAy+wiT/pFOuhNdSIZSq/f84dQWmhF1RoZm9ApEuAbfsFsDZpOpMbYD
nBLwjOJ1j+tHKU7DnQ2fVyRjuBkBbdiLNGPSKMtORQYstePF4SMdIw0co/Tp
tbPFHYjoerNXWHvY2n8IUV4clsi3m1Opqtbp2uTEPktlXUm9+5XMvwQP6Pdv
eyYeh2ZAywOlsqkcUHWlH5ZUfkCm8Xzl1h4kjwpXw9ksaDk8QyY650AiIhR+
V6DNKsZYRCcgRjiBoU4+PdWTjOrXmSJ+LVPkbA6Hqe2I7U7+369YXIq6Q8pO
JEpm8vcwubleNqyz4j2LvCCt0j5B0eFs5owR2Hmfvg4UZYZK/kvKcUpfmaqV
gWIE11en8lcSTvNlloxpgNYyYx2QVrh3gHp5OE97JXVOVVs6XbDbc6fUEtuq
bCSZU20b0aRufdbU+n7sf4+9GSA6l4t1MMAEIaSoGMLU/esBBDgStYG/oJ8M
Mi7g9jnBo25KeAoyqaesdFtzLbezu7np60nRi/gQGw9eITuHFGPZbI8yWs4n
5yYkkO+ub5eg03nGgdQ5Ue/8nOJPqK44vZOY8ld7EmqLSZ4BOkN+z3QsmcnB
LYT9z/kQ6CTm9dQ89CDNjsYT0skSqCzWDy2xQd1wVb9pprJigrjD4dHWRRYv
HR3g1/SzMAS6TTvqSa38FppOBWml3tdfdV4rH3iLzLHL9RmvlVlDUEZz/e4d
Q/sduVPGAIpPHstjbEmWcdL8mFDcoa0n891xkMIIwUi7mBBNHbwdVsmeiCz5
zxAJ141IpT1/pu46m0RheGxoyOYx17d0ye470H8S6Vk0mqr4yTNkC8GAa6ap
5ZJCG0wZ/rqsTyZDGyNs5sTv5jHSm2828c13YFdGC+SiRIQvW2/SOeffikhx
pJNb0VMsPx8j3xcB7ubtQy+0Omxt2WpVuTf0tHXGwkJUXcaO0GLyznAMFNWw
ILeX8jkU0gQlHFKwdK07fkVYO46d0hLdJpCH+q8wKiJK67rZjrzjfUBkDXjn
M83GeZrtkYVaKnjN/rRTEFlZaCGI2TGSbo4X/PMonIr3L4CMordPFQ7bVdWN
f1UyMKmoIgbxuusPjWsAF23//ZM189EUfxGickBBd6doC44tMzr94X2OlyPg
8CfNm+c921iRzwoAlMVTQ+8dK2vQVfhdJWLYgIoG9bvDyZ+wB1DJp/UQbgrP
WDV+C2S8eP782+FLWGTolPoivVTVaP4ZCYSREn1HJQN1uZlD8cOItUFlAwqJ
RreR/J/W1UZVqUFed8SE0WIu9CiSlJDahPe4odzxrcCepvpb/glb/qovLxtJ
CKRaSlZgJpNbT/CQzJwtll32JQSZ5S+6k0v40Hifkc9BG+ScLGaYK0jxMryk
5vW+61dDjzRo0u2JRP3pstVTw7odPGzFpx8zEP4Qevn28n/t+hvxDFrBw+g3
UoorCCnQnDSzM8+Hp4lCyCX/jRx4Vxniwt/6ab3iGHs8437COeCk59sHp1YX
2zI4tph0MyTuJ0Vz/uo7Qf6bVw1HnXg8ywcrzFZF1bpq2CKXsqvDUQljVEsl
mk6SzBMgEAPwNorMsTG2l8B+q/dRKDgyZBA3C1Y+rSAJn7ctpIhEUzEHJo83
rXEnsYWtfa3Hqelt9AV/7o2NtxQYPU77I3SOd5S//btRaXUtkbPzJuwVVhrk
s9Sqof6BMmsKa89IGvdQVBB058StOUKwHF6SmUD0mkfl2Csok7emiDGHCVqt
IdYwt0dEMbwVN7E5x7ivy5RTAgKEbF2ug+h4ItZwJxUUHRp90qIk01bVEDXu
y9MBTvtJd4b64P9qzRw24f9prQOSpK3poyP0VedW5i6pM7KbKKPvNff5RvjT
guyuowFITO/XO/Xm/HQlnRaCCcZgogiwDreKOqNmYq5jL58SAH3O9GZuxDCp
m9HIjyK6ehzF8qBuvqKi1MGNOX9HmzwoRlUFdSIjATzWlsLe9xPUYUMIGxT6
TWzcyxS3yiMSHMWAH6ET1KWsB4k1z7nYn5+Y9QhK1QEnrwM9ple64DJ5iERC
EgrxAd+aXBCAMbMkzEm0yiJEyya8DyahTrnxjFJFyWtQbhXRYMzXn7VmAjiE
yda4wNVsQeUL5MzvH/6jwEKqWQSC9zvdFYv8X6AGfxQJNjTiYOhU0y2yg7bp
zC+Oha+bxijwj/6L0ZsFNNTMmodQMHZSxtTXDGLpoD0rwmNwGQdBt5pPK932
3PbzMePTQ8KqwJ7SSyzPJix33nsH5nbYFV3Mybiv6ibFv0t7VtRShh494vxM
Fj+JvdyTe709WUVM9Omdc6aUcn33sU43Hi+/VEA9suU4NtY4Rgj83ssX0luu
Ly/ntSXFVymiCsA9pICxqCwNvZUjqbCP4Ph+UxRwxWvJAuNOGUfo4tox6Mx6
XfYguS8mvWGhQfgRGiHGQSc7HshNLOPJo+WeLIP+Y7npXPjj7nASfS4JqWV9
yaHMCtKS/Onc9QEz3qKrOotu2m1ir3IHcHTGh35gp3NIDYm8qK8+t4fj+c2O
uUwtNLLyuyZpUM8HhXvt1rvCdFYfUE4vFT3oLwjUrMexYNTaCkTMvMhdpjoH
nVTmBLsP7A/4+3FqdIbGEP8sYmqhq6vCxIZ/ZtPk1kbI65vX0CZtKfxFJVib
Fc15RQa+ArZ6kK3mkKD/Yxlht2P7zaVP4h3GGsbRaxB95DuFUbjFQlk3PM9w
ioeALT0k5i7+O4/aw4IwceuqvoA8Kc84AnyC686XbAXRZ3EamgilN0rc+o9g
stzjA0l9MQ6WvZSMN8Ww2WdKwmZu9y+8xNPCB8+ZyApIKTwSps5nuuxpYiRI
YU8vPjhovHEiq/GpsVU798Ja9ybJ0WQPdIK1AoaO5sDiXkXPL5CZPBq61KMO
OSs94/0XM/vHgp3Avif2tocunLYHb6PsPUyAYpcdEjWi1Y5fBd5OUaXTmM8L
6zNTnNw7uXZhEJge0q5oBgDDCT9IaT73MQmikLCjlqWHY6/Im1FsJBQ86Vjo
MTJvh2lEkO2FK5nIoRzokVunMARxcDoDLsFtBJEIwkfqDf7/Bokp5f6cX3yu
2ms/Kl0uTuC9lHnR6yKNBX05hqd9vHL24wz9YFOo/jmefGY2F7GikNSFZHSj
q8hXSKTcXIyfHtvqahEUwSCVMHHdpL73Ye6wqIOcU+fb2b2Cb/nlA8wa6Z4A
iMgZ7tvIiGcX8h+YiRC6Fri6583sE4vbWKEopixWNj58QF+4fN5eGoQq1D6+
3GL4akZveQQGlJx5TT16l9P249ebgMQQ2QTF4zbI78gh7uBayqfGrFzX7JO/
VhKlWBUNGJ0SXx5aNoFuLyv8WRQTSXQiIxPtXX/+gqQOCcmFBkVzO96WYYA/
U7zW9RIsl0A/NOQs1vMDKfdPi9a0E0xiOHOhYRZ1r4nO6DD1Xmr4N0O/2tZ9
oCVMR9Gosl7jdusQTtY2RzUzuVvYcNKav3aM9AO9JHyC8o4sW90uZFzjM6e0
vShZeONpibnBgvPAdSPXe2+ptPkTbGWEC7EWE8HosgEkGRsVAT9Ip/Y+Ky1u
7Y4wnmQdt2QIPWtPKGmJzbxApN0LCIx5EPQP/3Y+bj01GHcDU9lYEki6a2bo
weI6uw8A1iDpCPUc4ZNz15K5pB/SA10KAkF38bRfI9deLZm1Pqs7jE8lEza3
+aGPQP9wDFYp55LDBR6NOwKyAO6MfO1KZRxrV5eH+AfCssPqE07EOGCMyp3d
RdID7gu48uuB1FV8UTsWtFMLTcPSQFFx/f0l/HvlMAuYZJrlWofAqDR7sAe8
lekHg6105hAK679WUoSE8P2c3pcA5SCXnHnvdhXj2NUlLs9xOEfj/LsBTnRC
Bj7fae5F/D8PhW501BdEIggMQYcCHaI9LbqoVgtrvuVJgoSUBLlSeVigG+KF
K8dkVOanGCCszHGoJcG5XSGVOB/jyNZJr5mqeB15SOn1ZTa5iy39C5WQNYEt
QvppNHOSTd2JL3xXDCfI96gY1S+lM+NbMx7c4sI2nwsO6yA/rFF04SaQKm1Z
gXHvz++Tezq/GfrFvx5Fvwedo9DEP3ppuunqeAExuxQD/aZRCxEn0xzE+SjY
N01PXbkEPd1D1mA1xl3PaNgIl8E6L6YIC/4KsEi5Mtq3HmLCBkwFp5u4wFHF
vgh/QNsba++45rL+kUCK4EI92s3Wz2DdnaCiW+VPT05cuUILJNnwBLj5k3+D
y/1mkOYoAWupO0p20lSoLIxJ+RiT2Rha3mjkcrb+iFQvS/1kh5ijwkEjG0AZ
oitCMScgphNrBcr1LGM/BW/Bc4km8ZRL+AdNDFeRTZ4anQ7tc5rLx9VebsqZ
uKtR1LivnAPrhnNz76+yY27D7T15fEGlB3lNkl7tzMJiBQC58wJKYaZElZNz
nkEH0olcqwr23DJeCx0CRXZZmLPK2F/UMyX9z3qwWT6qJeqq5T0qvhQUcuMn
SFW+wSACcWKtINszp2/t5kKQ5vcpH8cjNJI2y+ku+2eUiqOJ3U66JZknwa38
HX8YCJ94bDpQeZvGuW2EX+YzQWGDTeNGtRd2pMdifmiIYpj1klinN1QZ+6Fd
I0zR7FpfbX65Igo6f8OK5HhaGSTnP4Vh2pid8wVmiGX98/YIwWYohjqauKvV
x/318Z5S9G0ar078mjctaEWnMUlKBqPkWGsk3rM+UamI6MgjC9qQhZM7tBxD
LQglgX9B7ONndMkERY3ui1FyZbXfAPsMl1VlTwjHOmeVbvCgG+ayhDy3vaLA
ZC6XSEYvvDQvTDbqCWsHrAMbc16/CtKnijWwss5Eu6DaD3P4O0Hnof6/KFKc
aPuYGgxr2JYc1xcxNkdI08FNgyIWHVhSsry/NmsW1DMCU9pJCi52w+7O7wm0
Y9VM6IsRRq4EXBd76zoBgDVQg0nppH2FX2x67bzxB6nuCqdogUlIjdk2EZLh
A/eMhkzWK3vzW9Nxu9aRTsTSMKwuGSqez5sabCa5AJCp9TmjZAF1QlCTq1pZ
8hYz3cTZra4YapftT+sbjE+ovOz0HBIDSl/0wjNj2T5o9yXWZhS3OxQKWRwf
DeXBbdzRQVvadW/IhNlFXIjy1jt4OH8ivGqm0DOpjYVNUXu15bkoSfGjAv9K
Jv8B0m1/rl/c301NYk8XLVgfsB1wCuAvodqiorABlsfk3AlMMtb0+hI2/Vne
oNd/ZUlcPs+4xOXeBKQ49ZK3I8vKT+B5ocnQLMJqFDEt7PpbG9+t/a+MwRov
B/JBLPsbJarRnlXT9aTUzujOKyd8Og5JIA7Q/u7/GIZ7P7bxBoUL6W97aiJG
srsRLnJq4JAG0D+47B05L6YLnRU+jBEVv+sF3PvcOD2E7xg/c7NZ01gBf0i7
n1Hspc3HzZJxgukkoN2Hcum8hCr8IlyBEakK0QPIYTuAT0pJS+80WUvB33mX
Zrbl1d9pTOTGCFdjOvQi1w+PhX8W2efjf21x+0ivQg5Rtq60twvBXCwphNB9
jJJDp8QhzqUBMnpJROyJsI3OwFs20z4EDcra9o18QPybNtLTSDYvYqPSDSCK
/JQxb7ugKnE9GhrBBxT6LGy4dqsaOydHot0jEcN9bUzRDxobRk+IyPjJ/JFv
+3B9SocDL3sf2YBDRfTZ5mbEj8dcl5sLg9bZEUVfwnL4Ud9DhPNOLphbz0pb
yjqNSxcq2CgjwlW28ygLFUvR8tDTQSd4E8VFvOO7Iz+YzpgnjzL8J0io4Wi1
o8PGhCFHgzAdqhooFhE0kEMLGxIxaDHnBbURjXbpX1vXYajxo0nL/1RZn8aq
pzU2YpNYCS4FhldGVFuDi3qUTnA8iQac8sXV5GHUBdmKOVI4l71IZPxp9973
nRJIBXNxsMGoFaa5iNEbD/x5Xlr6VUxqs1gh82Z0ezaDEm/Zcwa730RudtqS
/HlH+JEBFqwCMLdG+EkwoKbbilt2DInEMBPpk7sok6WsQPPpTtPKOo5qOrkV
6wi1t+Jaf4R8TFE2uYwEtP8Afu1PsXZmt7zCANzETOOmYxVY9Obu9Y60VT2G
FCrptFYHimpWoZ7zTEhwsbqs3MCN+n5j/TN1IYx+Q7lpEig4uSaCOzvupNOw
5f1kARx8b+mD+PBVFkPqSns0fw0u/IJKCSmeU69jlcLBcHZ5/e/TIYXkHg6c
6BvBNUctHcApQrKvK2x1BrZs61FS82ODo4DGHqm1NsRXmMn7Wqw9MiPaRWne
yrFNLoPTbrHoBq8/wiMcGkPHYFPzSCVd1FVOXIVXMV5oJzvEnhcEEw+cxqTw
VSH5gNiaZhmbyDh0BjCC2yf/RS+/phZnbW4h/RwxOiuYIuTr8tQHVgTu1c9P
BczjzIqajFHCd59pXye/R8JdJ/rj49S+5dWYnJk1uCovTRDW6gk3qFyBO3W5
Wqx8IfWOfsuCY0/cTnXcM8hwN6VOsXvIjWWFGIFtJLxmNGrz+jz5R0VjEGwG
5ZGdcYan/1WMr/V+H7yx/6Q8kK7DCKKgwgIoqahK2JCiRDVMIO7CMr5XfeOg
W4h6kgblzVWNdmJsc3HgS7YSW41nIMQKCtKMDegy4e+inJGHriIIDCG2lqSv
i7EoBbLwABmF7GMD7JM2h/dDCudgvOxdSY1f2OETaXaJKEfBOrahvSLO2SYW
qN4fk8OmpFUfZ1j6qlBTqg/3cBCoW7k+8yPXZtGgdfu/HtP/68pu+MboSBpE
R44xOatKTYCiPkB2lGR5KHF7VWas6MOXoQpjKzUT+poirGsh6x+MYRo2nTsq
FKfaussDGmXZB+QM7vLgmRXdkUn38c768th+QKof7oIj8oMbV3ZT+AAtWCV9
DngG2vlmviEXYsxgNn4kd3+lwdrBq1jokmWsuy51Qyh8s36saSA42xNqwLhm
bObhJyBPDnw3wrjB6NVbhjzDJcM/T/bGvS1I+nodBnEvK8XjekhzWthUfAvR
tz5FAxXsPO5PnP1b8UPRFcR8i+HOjn2ZxAQILO/pLq/slHGvGfzCEBxBoKgl
3a3SMgOYB1ImZyfeF6pFO6VlBoVWtXibgBvVHEIoqx8kUUBWYV3i6jH9GlJL
ARHJ8xGNvsiSgX4u0xW6P00cT76/uyoEHtwognbhwYgg0C58j15Rz+7qO7TQ
CpTJNEWAsvXo3RLCi6bjbzRnFK1+mBdMDFDW1D0fy8QWnpYjSIM37uuF7wjL
IBcPlT6wLQMotC+/BAVDB5XY3fEKbPYgq3BytK0wxD3A0jlTD/J5yB0GusQy
4sDq0taQ5ELYSdU+4bV6BRSEzxcEOkp9FUlev1zJHcCjSR+cUADRKyYudNpV
n4ZOFbZhyWGvfPtPMAB/zBnSwqFgegJ5bMdBo0eZXsJKXzhZsSyXKRAaPUIF
cS+HFqzTwSPG8gSxB4Bc3K1PvEdy9YthM4VnR496TLB2Kofzz4p43z0oHLTP
jGs88A4PUUWrWWuGzrYv+Z8GjbshFxYZG/2YW3qsY5VXL7+uC/CXWSQeV3f+
NctDzUtib1oUShGfuIvtUxbFAWoB81z75FgJyl0Tk8I/fpCCNC/g1h0Rh0eB
l2bwSr9QV5Vt3aI9yBg6LeX/IDXBCb8Bgs3fx6OXJJLarGV5DA8/zaQU12R3
Erkbld+ou/iqijkdVdj+m8QMWcyrszErUPTWHIbQP/Ai8pZ/w0lyWEALE4CW
ZbpE3PYrAdJyU6L/dBRV7VtN5oQyKi9dsqRQQ3/fvOwcz5umJh+oRuvnSamg
HWtF3yI4yV5EzbUH4l5zGs4Vc5vJTZFQNGKjJz7e5pEDegmJzj2S7BdOxTqP
4CYjcvgVLUScD+Sj89x74DT8n5gdFXGocLVTkLpyRBP+Cyi44/RoFwiPcfgL
Oqucti4jDP5HfQTOfZGLU+mWuwe7RU+XlAeGGA2t/RUlA1MSgHNauIl98cOL
OxJi1yneEqfZQQvHkEviTxrGnbMplOBNHJ98WPCWHJOv8oUvpa7sfuXEkaXV
QUfoLpbYmtAY3QUcz8YczqPX0O8UF4eUBFodnaz+EdwopTQW9jHrXIBvd/mG
qOb3tlmlJymt46bVhLv9TofW/xEC87ZZFervjobK1XzckF71ViuCcA1mZp/U
RtGoUjChFr8IIviNXUUMcFark+h4lOoFflhcjtGJLpFdGk0UrWEEp4DHAzWL
ypkAZ/Gr9YG21v8rJLQRbI4hV6gOnWV06IPiJ+2qhQ1NLTlEvadL3qW8dAor
QUVHQxIedc6AdBCoJBN0GM6AxvJgpRQ7bI3/ELg4Ix5CghLx+e326lMqcd+8
GYdPrF4RNXYeuGKshc+QLVJ0YqEsHx0HI3g78P1Y7cY9lVQrAjVA+2Om7YKK
yIiptVoCamcUcZ6IVQC7K1nCltsTTstuFk5P3ZOPPd2HU5Ce2+fYnMfNjnQi
YIrvU1AgoC53AzLRUYKuncGQT4ookR8o0jR7CkltZh5Utbr7BJWHe87Mcv4s
cgxa+8GfZIRTvOE9b/P9rfnl/EVr0d3yaxXNU8+yVr1O8cLnep4IZrcub/4F
si3ItTPG2SFJh5+PD9F6Rqps07x0QT1vnFWW7J6YVk4a/Pqi3DjKEHMaVubU
fIiJw6ipJ62HJGU4BF3QqO/994PIyxt/9ssD+Ca40jVlGUwNLrkPXrE3vJdB
t5qWvz2f7QnTuewwsm6IofUMhla1487PsupLpXTSjzWvdA+cjVPjPXkMC5XP
UYFyxQixVFvwfMXmbc6/VYkQR4EmP2pgSwEvSMw/7uPZc60+qKUkK4Mc9l9g
+jftI2eQAvCPwwwRcOae6aTtTCaQsLx+C5vwdkleV2FjK7nr4aHA3D0UhZQt
/c39KPvbWwLI5V5tU54yJvksyrTm8yZe5/C9AIMqtcQrI/V81Rrlj3+A+EKv
JVvYF1jMASdugp9vZW2yxEEbNxv3C+OFAxQ0jvzGzyYyXNQahlv8eihjx++t
AHfrru6DSfX6M5m7Ktpa5R90T/hOqv6HvsHvRS6V0b31qswlqsk/lu6OYcvR
ZsREXrlvogT3Lpc1845hilLzCYSrsUBWuJvQ/0bnJ0IOEXsS16zhGslVxfCb
Y4rmxygpPMD7Wx7pa6Psfqh9yNf2fGmCM1PDXviP05gLjdnZ91IalPz9JJRz
yGdugxL4VbmuxdHw3ya2fIh3NEHURzB3e6D5WMP2YeN1ykh+RYdlEtb9evtF
AvYOQLXHSOgKVZsqRB2/tbp2JVrgNT8FpR3zG5Xbh6cIl2fa5VyZWsG3J70J
J9ntQL4lzAYJrRmJ24a2kDktlpifpXoxu3IIU6gZgg5v6ykfEqPQ7/X52GWo
3zPh3wwX41V4Wh7VrJzZpHl8X6emE+dzN7PGZyRASWm8lzAXgOt8QeVOmmxQ
fP0WNsDX3KwCHrAHc0I+35XSkM32kS+rFUfjJURe4eE7ykJB5Huh7/C+lof6
6GFTlvff6ngtZNe+eMjn9q1OZRfexcWyyO1yF9+Y6+pD3QHq9GPpuQmEzgQ4
ssg3ByLvkgMG0RhpquQtqUdGmM6Me911aZVJtV5G+KrRrToEGlPtkOgjraJW
6SBMbGOJfB/NziJKAHiRYfspQUN8ISLI7U/1J0L4W0gFY/F9gZozCIoY5t16
THTqlN1YaIQuQSwCxozGVZRxN2fulUBW95kgejeuSZZN1ZTDCc7QtsfSpIWt
Us8g491o0H+C+7yMkhTcfM2sWVR+TS686vGtgLQ9jSSa/JR4kbC/Tp1E/S2O
W/gfe4rDhsjmVSO3r9uuLrXnuaOLuKzdOcQwVAwiERQHhpaX8ZYESNNDXODM
J9r5aOBqdYgf2W5OzB2iQ+ikKiRCTSpyyplLiTpOj3uuzEzGZQssI2/z+97w
F7djbCovXdD7HyDpLc8AhZdr45qkzSnFsOiOhFelzYF/gFHCjJvEY5J2/H6/
WuEkHPOlKAXb41kavV0EJF1jk3O18jYAfzVhH95jHeuNLF6N928UbgNXWc+T
4lhX9o5vn7Xx1i6qZ8qcCzcW1cJ4wACUiYbJWmFGkvjHvu3onDWt0HTbt0pY
sS22oosSuY/EKQizcLa2JP+8aVLwz3ZybYh1TQm4coqPiZW9fmYX4ANUeKlV
ke/2xcr50wOfHE5O8fRfyBLdaBKqH7VZRS6/CQBCph+xFZd0k6OU5dITLV/M
BZ9HBIDzH4Bc/c1ooARXTCXwOx1/HzaYsOAOXYrsLtXiGTlIuF4HP3yy/qi1
EqSj8u6+8wpeW6X/DUs0c/rRC1+bozuuLNgzFsuWuS5V7j06NItIH5L3me9Q
d1n+KA8MG6S6OvNQZeTq6qnAhatRuTtGDTt2EeL0BhlWt6GeA8onZNIW94XI
+LA8mNI2vUYM9bxzm8chTTAHzJ/klmqL1JyXSf2mbiKA7ggc9qdlCa+gPGQ5
Kq/b8jO2j3EsI+p2ze4ptHL46z13Yw7cxjY0TNClaA+X+gOEdFA/zlRKhx7d
2ELBdIGOZcfE54fni0/9jiign3Ux6+MppG+o9jXw6M8ot/ZHQ90CqyAKTLDA
wdsxHFY+B/0hb167I3cl6HH6LoPlTsDSzUxQGPRqCTVNs0bg4ibdd5QNpfJS
UnLy6zjQIfohYMzxnCia4Xcw9wiBnUVPD13hJP7fc1SJrd04hiPk9mEE/IHM
iF3BZpRLloG79Y6Erb4RC8doUH5435tRvIqUz5yybEg5szYRbiK7jP+nMFy1
HBqxJpsdbHXt114tNT3VR5+ANL0j69EvHfl5wwi2JUkGCqV4pduymGl3QVnG
hhQ935ZYSc0PXHr+J+cSpd8u7idJe1YvNIDlaV3cxKWKb9PTRtcFeLjCKwA+
rO3t2Az70WOGBT89wcWM2d4Vp6mu3zcney4rRXM7cyiiMWu8G6i5dnL+3z94
3XNtnRPXK15S1+NO1ly5NEU0itVJt32FeNsKmRBmefnGoFYcNpvlGhhXMq92
OFHSt3iMZCX77QVvWPRuTmGnH/m8xYKhwKSSdOLiWxam0m0x7ZxnDn6N9rx9
DVuhlhTvBQLQeNcLxlGf3r6BDfrPR5lRvDs8lzltSdTIr6i34gM3M3F1zmiz
1lfIyrOsHuL7/bDq/M8HUP6TLb6fpS7VShVtbYAYQxjTE8sGM/u5iKgo8gz/
ZJLFA7sDdry1TbR5h2Ni0E/wE4fixbYj2IzMuJ1nZEpVe2nQltDKnXPkPAIC
t9B2ZQ68DgKGhxY9JLlg8+e6AJSbJfx+b1Qwsq2M2h3d+Q4nCDmRyJu0mdkb
htiTOq+CJ8u9GK1+NSxHTC64SeyF1cXRPK+zVT/IZBG3ITrt9YSvLs21DAxK
kufbHIo4RWB80V/8LyjGARiSyS0U+lGBvEGupB92DCmfpc0EOWZ6OGH3UqTJ
YaQidIw13FArFIG8OKDxVpcVn6FtUWLn9FsnuUpft14aqUB9GftHiFa78TWu
VURZeGl5whTx40KgDGYcapNqOfnGFJW2nXkhq6YfJMtEWCyOP7OoH/6o4jK8
0s5s2ejU2P2+vVS+rlOB9HGkGKmZUumqIANjJuiNRSLI5lV9qBV9YuI0VkUC
+VTMQeGjhRrpE3ASutF6F8kwcDm2l0OKZCWDlvdV5QSpLCXHsejLUctLmb0/
lkEn3eAySBzl32MUpbKr+dZr6lmsiaGvQTi3fK5J5JUk1qTU5E93ZXjfWZvB
sLb1/3IrluErqEdOVcHWAzO2nr+jyqoF2m14pENyVi/XnK78CVqu2kct5qhz
Gjkq5Af1b9VcouwJSwWKGocOSsQIV+d+IW4JXxD9AgKV5mJDTbfZm6Ws7WE6
OdGoPlaK3MVLBqKJ1ikP0lu323G+ayBd7WG17f6VYZ1g6xPjK10KHnHYSK+J
24A1kmJJFchLauV6i5EtHecN6DFvvIM6WZTRefi/Tt7NXk5D5CB1u4Pt6rJQ
6xQEZVEc/Urk4J2C23X7hgu72ClgNdYI5eNlbRQIi4zAWUD72Pmq3Qlwh4sG
5a9jx8j22FP0c0HxVzRn+C5JR4XCj2BzCy/hJV5pBb2Zr9Mr1Q6Fsahi1TgB
ctDeo+hHQcIrVVvFs4O63u3EwmWsT8XTlsL0BQ2z9dapjzBQHnqMa3pF2GLE
DQdAQeukkq0f/PpWcXEE78jav4xWVCCD/a5PaNhVybGl0+zGh+kBt0mKAtDr
mX7LwjhHOHwPyQOZhj8oSwj27ynA6x7SidYJu0rxg/yk5/zQhJQIQxWmDTS0
x8L38+UU2eHT2+sUdw4+RRM4WVNLgvOKAZcRiicuyc1APSPUEPuAlKLtSkD2
uunHVfPkCPlMcZL+qPeo7m0ecZIAdYkdvPJhusRGxV8vKWwujuXUS7ToDVzr
lBPT62culy9OgIW9Yhg7GzdNyoBcIf+1XYyItbWur5pBQhntX5cuU7nG8Ash
Kn/+leZNqS7kPOJ4Dd5UWAtfi4zuAT8+pgrSX09Fltxh14f+gyPX3ie7ASli
D2hDxfP/D5s1Bs9sx/Opu0u7oUmqMpA5QhjnXzHaqf90ZLOpBBzh9FQj2tuP
SPdTpARxZVY83ZZCTWFmXosWttIz3YFOoqZOL0Ps3WwDoHDhWjkfrW20Lvo4
VMSm8MD1S/8Eq0FRieA+XBsmoc6UQAhCwHQIlk5aMSrrDOrVcajQxkUqdciL
VFfWWRrR8Pk0RWw9LuFF4WSyn3WuRX+vsB00UzGQ5kGvessG2kBhskmNpkmP
Z5sSuxdzk4msAKTNI69+8Akf7mDQ2XrGfxiljR4bHhPb0l5EO2L915lZb7Dt
Zapn6qpAfqjCt68z6ggaJWjTajhbBkmqgssmH7ydLe9gSZf8B9PIsUj/AyLJ
QmYHJzCwoaZwwwtQZ2LvzUc8+Xw0LHai2lD6eQcpirnPHXbx+xWfCfusHsNA
KYGwpBvurykLfosbSM9hryMKbVHKYpluhyuCxViTgXBnJt/Hi4IkwAG4BdwA
lDnEvCejqy8sx9hxYbMcl59+GeV7NOOHJgxxFPSEsO7fpgV0ImxOyN1/PK8a
y4eDiCUr8l+zGWMBXO0yDOIETm0blhtVfwXqq53vKBANeT9Jca3iGigx72mk
lM4XcwjxfjdLXOi1/rGQwc2r+aMY3KmUhMA/f5MN1yo2vKfsoxcUiHNo316w
UJlHrNOY1TskxdusdHGBA5CIOxQMOlcE9UWYh3vgQCNhAXMbzrpQBAnXOQiv
GiOdqdFFDwMCcdBLuNQzmi6mNUuJIoi6MYhl7Q6KKmytuADhlqTDJe4qo7cm
oxBiUaXcwAG9A1vwusaz6XyfBNOwDGUmxMxdj46xMscQCYBrRQ5/ngkvIsmn
yWJopdiCf5pGS5deeQREE673b0SLf1TGAzklbxoas0PUtQdg9AxOxGWShfpL
UOTtNk69St+bVJqLzj/3k3HmFv2+9RPJBDQvME00M2D5Yl72XeLtbaGplhhJ
l6/Nwp+N7L/ijdaoMynBPWjiPwLr4Qlwy3E4GTeaVpr+WGUs0EwBOt8/TnSX
0OyJc+/JOiSazUdrANlNaUh30bPxllFuBpOhNUKcoabrLY6MoEYBcZJLxrby
I6YD1ig+rv2067fZHxsoXNcRlrLIkYy5YB8HB4sxOzmxL5EDg5S0/kyVZF8z
TwkM+M+DO6GVou8PXt0DitWbzosDN8764/qcbW3aF4nrBS9+Itrf31LPVoY3
jFzVmn9Dn9+JdRQRPWEZcPunSC6cW4yQwvx/gxw1EseDdff1N9pz0er39EVB
5TeFZNP1fuO8ep9lrL2/t+xZdjr+9QxgMUoBYWm5akK5XitLf0Gw22XAan+a
lRiKN0icTiNqVwXJzoZLK59pTk5GO7GvYaOxD7YuAtYRHq078EdvEuNImgEA
neYNGOnrgvefrxWNtp0tIQ9ZXGr49z3CdKUvGtDjmQu2xfh8cTYWAX+f277o
NuQrpdIvXOvJ4sE6pcm3dFHhIAUXL0jA4csPYLfF0j4ieKEXtsMviLIDpwmr
wDJ+knVAQ6DA4sh3X9clnOkOaiYAGapKjpb0AwNbacKce66YCuAjRXlrmUxZ
YJN0jIwpUTDsbtSNLdOZZBfy3SO08zp9s3VoJnZUUiSpbRbBtZ40rUqPPj30
si0yD4uRDtMA+t4K85LPZU0iO+o+wtrM2Pa2V2TVLsW/G0eymPK/YF2p69bv
k7ve4Ykd9ZPqwmhHDFTciWudb8I7SKk5DWSxV0tq2p0x9MG/jS7MdnW55Zx4
ap/EmEYUN7gl7NqDePyVMjXNW5YH9OrIBkbr7rPkOP2qtJ0CtM5QY62cnPc3
uMeqIj+jIWKAahdF6lQDfLG7M3BLjOYCzS3FqLx/X1MQDdNio4iIGtmyowO/
WspnxoqhkFUr0yWxJtKn/HVCJsvsYL+fqJvG8niBqPnxX/WDX3CqcGCHL0QQ
b/t+1QKgyvuJPnw4YUkH1WR+DGBXpg0GpaU+RSW5nq+lrYFHf9ixCwalMtQq
lUn8sZ36cGAQwpzqNAeYLS3IHXkSqa3nStqAPM7xkK5UluU46JZNfAeYbyQ+
1kdADAabM7PJZaKO6ezsilUlK8Y8OjRqeSVtARGKnw6HkECQNq/usvHyGTLA
xTJe0KK7fKllaXGkmP5WlHSjDzKOoJPqutaTGWMWNlDq4jtyF8MScOgpmQ24
UOWdY/zdAWlXD9F1Sbn178VpuwFMUBfXL5BUstXMnNhhkKwxBRZ2dOzOcpXc
Y5ZhTFeVtLtLIrtsEC0esZ+0gH7FspmlPrnEP47Htl2npKeQSR8d2wiPph5W
gbMwHUABwKc8KudDu+/x2VnrEVKQVJeBgpIYQPTMVTuXS4FwWFlSZQKcu4Mm
cG5u/d2INWh1r57AdLoYy84MPFu1anRyDWb/gZ+igAh7dZ9qP11lNX0cuOeq
Ba30Ezwo7onnE86fisAmgarCbSmY0fbHr7pgfKi82RAONr1jqOJBYEjnO///
AzF7ChlGaBOUnLcl7pcZ6jEP8HbB/AWY6U3rTIAvMT0AYjoGLPsFy7wqNMXF
E2qMeguuZ8AmmXBRzg5i/hla/dsI5qLvLxPOFNUsfHPh2cA56idaSGrYRFZN
dgeCrudI7Wmc1tM9HZGkSUPgInKm5rWEpMLoQJOHviIxgNu8N+ELOFEwA25T
QboEdfSdjJoLKKCsAsSs/ch6S8O65yYWl33Av5ASliPw1cdHxFwZRYWveYqL
MDpVutcGcegL0cLjfLEmUPVEQfxzr/aPS8PwSQs8RFjnB8coJk9Flsvyl/hK
AeHZR/5ACzogphaC14LPzmHT5Pa9oe0H2kF2e37oxRP0amXIlFcX8d2vRTFq
Fr4Nx8CE49jGSr/3vFHDw5Fp33LXqA4hvZExGaxT/bzxwSlI8PqlZ3Ig+7p3
Pza1NBnuXNxF2niLMzaCn+1SVR6woRTD8jFdDU5QtITIegjwQKO2KGqShwtO
5GwB5Fqo5Ib6t21ygTD/PTgfwHKdYU7qRvxV9D2oF7vzDwZuqwvpOgU0zgLi
jTvUno0fX2noYk3QG7rZvWz/0QPIZ/mxcH2S+XA5PJumQuX597ufhdYPsK9u
CG/ugHsp7x/0PIIyki3eHi2dqxJHtdYhIR1nEvLBUtEON6ViYP4y1gckfGSs
PNMU5DvOM30u3zf4p9vsDPYU9q0igKeZzEUpFy8pth0yuE3mZDZICTK9EyxN
YVf52xiSZP+t4jRiY1pEkt5REpkDWA16u1lG0+v1J05qfW0kXMz78hh2mfhq
EiPeOzrGZnWK3wiFz68Hw+GCl/n3pjWskJx8RAuBoStC1ftMy8G3mPtnpuzy
gnDhlgTBV7wpCKXtm+YZwHMGbS2u0N4v2M4NIpN1GlByAvXf84mNuuqlyYq/
4G0sJOMBrcvctE0pUko8jttOu1vDwiusBEoviaryNwEteQx40Vl3rZiDPTd2
gDSi0wuNVuPzUCiv1sS2jU5ne7am+xCVwk/EF1KewLjMnwT1BHvgMBMpnssL
0gofiEsE/IlocIbJ48sZItohkZx1gXOXmV8BBhWzYrZe3X7N2CwzKk6zDS+d
lFrGwrHJUf3z77ixjBhU2KQqyTylcy9a5uyDd63jvLBFswGerbxB68UeJCbD
cWqeJ/VTL7fhrH4IvjiExI2kGWB28ZLqZvc48UNwRPNU7kn/fImc8k2j1vKi
WjIVoU+Fuk7OTTSpZprPDSdyhTiT6yPl1m+NT+YmWMkChSsaQeQyw/bPaM73
9Wb4rJUa2/a8Nc86HS9E3O9A9g6fDOmyb5G/KAOyWa1xicQafW0SrWyNIFn6
aj1RlyqUSEhYGuiXpM3USNPOQFHHrAYt/GvEuBDt8BBtI5xjXfWqJI+9tGy1
tv9a183SHgKYN+sCVzBZlj4OayqG9eh0TtrfqUYLQfVbeBeMlsd9WJ0SEwGg
C9pRpmOJQLAwYaaHtAUspJlGb6FXgWGDDD0gi5895bcbF/69wQp3oZOQIrj8
Z9SocOupXZ4iVsRcU77matT2TX5aED5jHiK8ZDOobt4so6y3Qy2GaQfgrOAB
g2viALqLvojfB4tWVBOIXOEfWtPM/3iYaTiyjsU8tItqDyp0/Dzd8IpTQw97
ZhJA0/F69xmvd8DKAW/zR2svUslULXxLmDlLmUUf5H8lJxSXje6LULHfEKlf
snsb3OTECIeq0T9TXDXSUN/VL5VxqAoHyeIA6oK3c7pHg2790MvuJjOQLy4w
uMOPF34tVeHnVm0oODJX/FD6LL41tMBBEvG0ecUjWF6SKXJaK/jqBCISiY28
F0EbtKTnST2OSF2MAxExfuaf7Mx6a9nNp8Guum0EegFOfvURz1QCWJlwax/E
ThJNNxZCH6RnxSUTaqBzNCr3A4DpOrq1lWtVfMIqr810xstKGMTHsw3RLsjQ
/XxLAjbKP6HK1KL5dxlBNm6UOryfWuq4RoZFNCMlUoYLNydZVXEFcog/c4KW
JhDiKuY2h7hxOiRviF9Clk3FVAwaQxkeR0ICy6xe3xtTsoIM/hbpc8xiYdQB
KUuX2kKaPsRO1SsGZjXTA3pt+JZrPG4S9WxbeBdWCegUl0D1hKBuQeXHSDn7
Q2tKxS2Q9rbgAOqqg6qnlxT/AX2E91WEck2Gxuu+VyOWCcAx1TlvQt0fscyF
plMx8zvxitQ0OMzNK+nCeBHK+hYU26w53I+86nMUN7/l7+TJyqjTLS5THsRk
JD1mm218+xauVEbSda2VWwQu78+CHNqp1bPiVj1CYQiZqqvGxPWIZVNS3jEO
PuWdByMBhWZwfRYjSXZZ89Vla01u5JkLWd+SRtZAx81txAayNqoEQBkONROg
8/Z9cZqQkzuNkBUMtaAjyQ5Ca4aBlBh/xoftvI1DwrMVN2nIlXW7n7ZJRFG5
+Ve0hs2b/CwPFFydltzze1S4xf3TwEYqWYYU2HLgBk/A0grTxJMbhTT9CWht
986a2JTYwPxOQVUr+4dImiDymWLCD2ADVyyBmkphkB1iYScJ3r5u0geROaMt
WcNavwuv0ARjpVpH0ZovLWkhsh0GKJfGYjcpKjOQd0ZZIx8HA0oq/NCrIzvz
HhmqOn941c61ovANJE56E3F1DaUKSQlTNCflTn1EVeSAngx4A77Cwc5hHGTu
1pTZlUWNNngY0h/i4Oe1qb4nnEbtiiGX1mLYy4IX3Fuu1BD9QaduNQwx2q+Z
vm9D1oZTsrl8+ZEV01ODExDJ+Hl8/hlsJDnk0gbplaIAuo2m1aagA/4KzUAj
u35tDGvZSDo4KF5lXKjFkp2K6BT8n2+t2OGRh04kD7K04Cl9ZXgEuunijOCf
2JML46ZkmhNcmS5Txe0SSE3X8jpGCxNzTEYo+bVcEfRJCPuTqx2IqUjkvSvh
m33TUs4Duak76SjWcHPrESkxaTwDcRX0g+VYr9jOM/YEQQhZRTYfbkyKVcFo
BmMolIGZa5tJbG5e0rZpBdck6CXt8NDcrTgDzarNpKY/dkFMJ9Dd6iwk7BFi
3N/k/OzOWXDN2VR7/ong7DXZX/b3nWi6RHBmzjgLPX7ASEKdjffAfSfX2+Kn
EOeB3jrUpEPrp9IXZA5OouygzaYFEllADQMwkiMetOXlNTk4RZnyt/1a2en0
fUD/BjIEXCzHDSG6gTmG01XaI5SZ40dteMmlvHAMFLIdWd5nv+XUCaxdQMTZ
wiyQQE5RKcHa5U0yogZA6Iand0iny7K+6Mr2B6s1Pu/FHM/Gprs9q8wVy6+C
lDcfCNkktxRYxvL9Rw8g/115ie4y6MpOTLQbbleYo1T9mRyFfxuESurj9BAz
unRhYLHlz+yPfmInjAbU+Wwl5tjGKk1izdv0n2ojDeaseS2UPzyGF3jgOvaK
6o9HeQYx6GfZF6PrUcoxhmdL9KbQFlMEGlepZFKUPQwtA266hyjQ55m6B3C6
RzTM97hM2Eg1KcIWU6pgVnA1KU4cuNG7DtiRmzgQieew75keH2+FM+RZC0iv
8pupzytl0U94ZCAqfJBDzDGB29v+WtwMuSYviZRfW60CxvETOHkz6yDg9ckm
dq+ZpYN/j9G8NeBl8DUG9TXCMpxHpGPq0zVRRrbSozSGrUKiHBXMn9GkUBaW
g4O5fHcfrnNR9kgS+oLbwk8TfnRF6gBIjCxXXpoSWUQl/EGasELHl3BcdDFD
W9DsWssYelyJxeMEn6uoyVSIvbn1hTV4n+YKNjEipFIkQ2Kh7OAfHnePzv4z
gbbENHxHzrgMqplmO7ZtZOJ8QNgsCgDLsxKDiX7lQ5aae8QdWKEs6xlYO1CB
5axl6O6EEyJRntVfyg6sOocSMkVrWpgr7sXOTDvhmqVil36p4LrCHR4bx3gv
9fJEZg0gewaokfLmPYyR2FHByNzTF+lF5JYka5j+leVK1lENO27pQOW3HDgC
IafabXxkkFZrSQafzpm55vw89yM20HZL/CnOdY/AJxq49/3lzWrDJj0DsKBM
jCavcg9uGdQkDxPJfuw1gEj0BVBvWVsdIr894x882XCn2vAHeTCJl6rdjnz9
Qyp0BREI+czmJgefy03nr1ZHlnnVUjTdBdDijGmcvhz/bm5zuhT16YVQPqV7
8BgGS54wsmoUDk13T903cjvZy1aJkDfYbaFB2clS8RdOuugI2tQN/LtIbwk6
YLaCQLaeWRiigsHpctheoQ5BednvUXfqtxLsOHKn26lS5l0Az5r0ga2h18IY
nxXKR/0GRhkywEtsrY1dirpaiuqG0x1Cep1furC7ySMq+237ipGNIfJBhhnl
Yi+yP9Xfp6ShDtfp0NNiS5m1Cqp9KFE0WzuvvqNGskso65IdlHEwWeNM99vf
bJN772mLWkPvq5i0qXgouo0HhE8X1inafItrmepaseS9qoqzoprMHm1TQg5y
t2m9q+91eg3UymjILDP8nHUWKH8V+kOxwSBkSuO5wQCIVwDJUQWXPZVckK0f
yrJ75MtAc/PV5L9OxNcNNT45QvIE+9hyLMB9Ehg5IK3Qr/38lffvCN5P3tL9
5rgUQ5sLg3Sbqh8CZ+nonnosU4r53OjKJuA8g2DavwwPQaZxOXhQRGYcHwGV
BshDplGBcYdwfh3mz6eQfE+0RTM2Zn0jqApYeJZfepSno7vUH0RxRSQOl8x4
01c9bCrfU+EBIXI1zL/smJjm2EC58tQlxtOmxFsbnlTrOJASyqSCmnd7RiWx
/2divt3b5Wy6hx1p2LZebcNHF6CzHjvA6WYfQtbn7za1S3Rw2kiDBDHmYj+4
9v/xB1aPELhrdM5uWGyWnvZ1mRA85dMHOBtHNG3NPLp22MBCh+LKNUuUcPd7
hpQ4TcJe93+qDWA6b8N6NcV57TJ0ZPy2TVkzVKDuLz3jNP5iTtZkY5SK/NYG
yMnH0mcKlr25nkiDO9hfHJ0z3FXexMaw7T4pycykCNphFerx1PjP3msGRECR
ji2QW7IRlsgQgpZySS0O+Tn79MPQdtHQNupe5ZIDipYMBuH0Doz0z6K4iaSQ
mW2YdYwGBvV6eC2O8BChAvva1tvJSZqxhxMgSGHFsZ5l5RlTplQdzO9zSCqg
ebXtdc9sObAGBaFgYpJ0Q4H2jSI3fAWi4okeu0PQzZhoGJluoeNeluIn8zMY
yGuqkXScGec43ix7lKxCGRs52mGWMcYa/TfbR20gnGGThPVaAw26iU/W3PZW
NGUKfJQ/lCE6ig/kV1rXLkMrOiSssleO3ONzRXTwjxclrEp2HrBNqRthlnja
diy+1j4dFgoRsrlBIrNw9VIG8iFd5Lu0lf3q1txzqOORg+DB9VMZr7Ri/rLA
rM3iYOcGv7QxXYTqrqAwKTnbDIcW7SreOYcYfhvJqypdo+sAyILGURT1G4Dk
IcjupMZQRAzPeet9xG+eYoeinl2rfvV7PdMKUc9tvtfJTQiOo4uirnQnc8A6
G9/6GZU74lh1ZqfwPUnbdkQXm6OOE3TetjiVPlz9WOUfJ/m/pO+r4+rb2Jmr
ixQSRct51ID7ZloOHb67Ex+oHu2yOGXc65NH4besLrT+t2CO4imvAJCLt77d
oD7bDzqE8fX0tXrDDb1PZX3UUAagy8LNm75SUjIZ4YXttmDO0W+ioHA4l1ld
uji5rXryzGngGRYcOFgVHkWgfbPa758BJeQ1xS5QItKI8vt8WFDE58Kj5AUQ
8bNUIcQOzLaxWg175Zefg3zLAcfQbQPJkUVFt51sCZWvKWq7pYBcyt1bGoHb
9p7vmvzZl60Zjigmi3xETJ+NXjjwbgJRClkLABpD7Il9jiybUkxSjVuhiZkX
+UhNc4ot1yTbbY7JZi+11euFDVBziyOxbbUeK9dNhpVAQNeX/7GXo0ik1zix
7+9BV/PDFGYskZJlY+jhz333sX3Dy0UobHgTZL+nh48Qnl/SufOxrwUxw2VK
1ePSsDfXrltz9yHiSCFnikG/zExlkffzee3yeK5wTcbLijqzQexPsJ2u56E6
5bDjgfz46CHD/6NgAJxNQXcsi7Q47fvcXDcy+6TaQ57PxDaURl1niqK2L4Yu
OIgMN0mBRwaed/cdJxD1fxFRBAGRE6/ayVum1MEuXsyOj3aE1bVdYXr59JmF
Vy3mBqDstihadfWQOhlEwxIEPEJPTWuCRCgXgJJMUFkxNEb8HVirndHu/xW8
FxIBQ1FhwfxUNl/pARcaNTYNTN/0tGHUl3JUGNo9K10W+gB6jRTE7tgIk6tC
8Daag94EbioNx6VMgnIyYCUE6u/uW5nONG9Vd57I4r7zae/t8wxkHozEl5It
ZpP6MK0yzzffDgq8RbIKUfWyZsPYZLPx9doqv2bWzy6cciRQkSX0DdyAMfcs
0H3r6jLhBkfntkWE2R55nTqyYnkqCIw/KdLCy1BSKBCOhH3sr06GZh7zqXo1
HKMmiagoLNZR0H9EdEJnS4jfgFUiBDC/1xG3hVFBzQbAPLFAStYnvIr9weJl
6n0klrQyi9k8CCEXj19/UafjchgyRWkiHOf/MFEKmuXVmdTDzqXrX09O2V6L
37wea9YtETbq5GvI32OtABgt8Qp8nuyqj/YnVSVAvvazs+aqEQ4dgYL7F0Db
OfxYXkr2xhs6zakF9SZBj5DRURw5f29qhRIqBET0kkcj7LPebbBS0ymTcMTM
YlR7rWR0xtBJ4hQPXemT9TJZxNu58P/ep9iwylDtTIuGgdJmBTWcVY+wlNJI
ukVnKN69Sq9Hf1dK0yJHuMsvHf93f+9xAi29J7Am90sX9DvJuHSQbhjpX8Aw
ajhodwtoXKVB0yCgVC9SminaG80b99wgLiQi23J8TNM3DpQdKmvchdjfUs0u
+pRbRhPJ19Y3I/SllpflM9yb1SyPi7iZFNjcZxYlZBjexcng2HU9iA8YgKjW
5jCE2FUvgznmEwtNLsVYvHVtXJXoudVj3jJ2kdzZLSy06UnNKQWaimBwN/Un
f6Bk3spsPol240K0S3ixuuvbGsLojsKSRE2tLxSk/L2NFzMlKVccUdBun0ka
ovmQ09WXl1fywhvuh0eeDVOHe6gYalz6Mp0z46WXk1lpQ5CJXEwRtO4OecxK
Uxv3DQbDHjJXKq+sp1SukfjjYJDHFrryDF1bzdlKOjN9z6VkSzgfBap3W8YB
j3gMCnkpojsVt4xN51NgiZNjn6LvVT9wGizyO4jr6VFRUEr9EU/kS1DbpqYX
QrpQV3q0Hp9zHF85lpMCLNbNg4boPfdHZVdqu9GizS/247RZfI/WLPl+avaJ
j/t1EHaXfLdDMoYF+MA9BcFPrkPDNuHmBt7HkXOJJXzTmLsVUoAotDrZIi39
RXR0YQSFNsC0uN540tbMKItqeLNrWfv9vqhrd401BM3anxxhjLI8Jp3FsPYI
8NL7RhEdk5mgc3TYdFOOEInIrR5pEoWfc1DNjRIBztT2dq/QohyxmQISK0Pn
CBXjWBU8vCW/ghlihUg/2m9b5/PU9r88/axxQ5aAhnRD0yHdSSoNXgJD/pJb
kwagU5fA2j42ylJOYjK/wo/KaOju76g+zz4o9oyXcpkidsEHWqL6NXVZTSO7
rKUR+RmTc7LlmOWhcbAOHeSE3AWMhEadWThEAWaPWeao73Bw9sCiUbRsb7zV
3RG4FdqHlJuEP/D7tiKOjcxipOjBnkthXEZ/hVe3KMM+Exc4YRVk8eCe6569
sXLNy9/wLp0zQBMvnwZz/4e1+2qMU9Ftw59iKInItXjVDsnI1uFpX2izcfg7
6FvknC4zDh41iSRdy5rsJLlKr/It5xV2IG3WmukUk6fByLH2AFLK1CIV4otc
E4QLjalwM779MrJWYlpX6C2yXCmcuD13iHmdfxl2TtmBEZkqc3rfDKcmC1Sr
O8V4neN6Z2qiBfig6I1Wiak+lM0eywRPJRQzm6wx/+h/Z5bKhuuizgrBX1BZ
RK3NMTGPg2C9MlqchZDazZ+G6NcTK0aw/qxDDQMjc1EUJqOy7ZvwPs+R/6FB
kYRLA/oYT0TDbczjDChSBCwuDYYkw1eRyG4BeavTdsDN5IKksqe4Zs3dlw7E
aH4cpAKbq0CkVooUMbsObH9nSQeEdecpwtDjrwuFYbjqbBc/CIjfJOqTcFUs
vbAVyblsLHksRiPG+gxatoRNcbz8XOrfTAS33hciDlTNFseQ77VwyqNy+Kce
F7PriyA/zWezhxB4as7i5ZiGF4WU4K5KFG3b5c/UmLjMnUPGUdwMQjTCWVRe
S0zxezlKWye1e1uoPN45X6eK/XiRwnG7vLPZGv03052OPeTAhdOQTJN3QT4n
kthojUIcuD8LxIUacB/AQTt4flbTk4QCQDW9sTSWHAOd+l8EKfcBcuAzkPle
a5oXxyB4RF5UIiW5bvIuNE6iWT0j187BMLyZzVXmH4xQ3cbY03VW18CXAlaa
r1YL6Y+OxiqJ3hMJ+uInuT+hGZ7bxTf3NHr641QxxET6K0ZSxNr5wV/Q6EV7
GQD+hMCiizUZnqAhfeCZBXlqVbQI7oh4RvTpNkqKekN1BoP5o4/JmVjEO8fq
f2d1bA9F3G3uIygDupyDZ8Z86numEuYBoq07DCmVFOj2L4lGOYaY6NLlC7DZ
90/JXzKsRYCy/+lH4zh2GJZKRbHCtBPaUPqXsSJbsCsRarlll+9p2Ep2waef
zB2QPA+IPKP4aU1dI1CRs5h17LdxGqiey/UWsW0mnkzGDDT5HrMgc11LjbNc
GnAeDwrqc8nOzyHNVkoZE2UTaj6Qb8eRmVPcUWrIgOmW6LAqz1KTpMNh42aQ
/iRiKmAn+rcVZ8JqB6KSxTrd9v8wID0aLXF6KLgXuOpsnWwwQAr7lVHBOGIZ
IOosHQ8/XV43tzsu0y9P/hM5Ksq8cwonJG4KsI3EIlpcz6oA7hjr7CUc8sqN
2rH+ZANZ7aSmlidLOZcgHrZ4MuORD5qcVnRkJEZnSEpwPGdHFl+ZGOgaUel9
BIRiyoUhp0qHc8XqhhKqE+XbRToeAXwur+hvJUJ8QsylMysmCwyOAxLDoEW2
m5PE9icCbxg7ss1JvbItdbCMaQ1fBKYVmBYnIuHX2b+e79tBDHxPc5kIJ50a
/nMSPtqOPyfYPr5P+PyKxXW8eeGquwkk6O4FKN6JyqFuyfVOUsF+y3wi5dUI
3Un6fvVS2ay2U9lboRJYwH25JqYFOMSRk/rTWeoxTfG07uwGaUBHYZUBN5I5
mf44slXPanJZSl20rPT+iAUZIHK34ec9Vhd4a7KIQeCnpSXLfTkN1npsK+5i
uo+wE5hNUOE9gj5L05IKmrHKl1FNrSFrB9Dh5awqSIUuVfNXKDTGxXT9Nv4H
fqvwKi0JCqzcrMpcLuBuYQHSlBfTPM1sSS78s6PRQmp/+73krGJjYAiSI5+h
A8ZSM6K97wd/p/LSYu9iXqvm3iuctpItHNbaRi6MrRHMHdZ8898IdmCe+Bxp
LK9xz61Tg9X7R6pHxdoXArvwJil7NnT63tcG4aTbDd8cD5HXrn2SEhtAOZE6
KJ27TxibjcYl/ltIHHy1HNpm4Mq14eOzFAxkKDiYmPNRuKDWmLikZHaihiLq
yL+MyFMaLMGRO6bVMgLlCGSOnOIMb69KZG1ymlLlA1pBvKsMhHTZnXVNceP5
RsEsBiqBsTNZ4/E/5djr7kU4nNrC9FivKWJ5sYqKiYaV0jarK2VmJkFCrNNb
JIqrEiFr6q/w3Qla1mE8XNOhOOrypGc+LeA1f+q3XyrlADFZE9CdCWiGSMDp
g8SXgTbrqprC4oWrm+CY1uN6y2I6QaVuLMyfC/dKuC+ejo852SatMCU9ePTP
KOlFdGx1yrCYkZZMh+fStqn5vReUmgd3kxlWiEWxHxV+dRzboGRmHGnOi9oV
PX8uM/37/ph4YLGIgLYAvAFrDx+Slv2h5MJb9fON/VV1DblLTCab7gmzHfuD
L62uer8CdA2eMYFdIoG71OkJSR/DOr9ktDYZC26XxjWRUSYzozBMirK47t8b
TjgcfTw6aomBclV/5Njxq9DO5VVd1maXuYU2LaMeuxXS2iSPOVpDlUCkHIzE
M81i16MMXV43/eMTpGE16au2J5nDZYg5Bqzf1aymiH38OtiDolk9tevjuDOs
3I2KM+UAcUaUzrnTJE81+Vlq1Tvu/yBlqXp9/q7v7e3w5TTl5pFcJL55WqzQ
/jCXFxxE7/HG8KZXF5De2nhdQC07jA7JyIIDWeo6rIsS3HSGNFSQDlTlFiBt
5WMtcCckzhoyx3TJlvbcU/c8V74rp4RGZlwYp4oHr4fRyrcty6kzp/LlBEw4
BjqZDuZrzNBbT7EK7O2RuisvGQrYsttijDbAg2QvrCpUWQPcOd+Cu0uoDh2f
FDSqeUfzrGfftc5yQpUXSNqAXC/Ktxk6yrbyTrNjm8qsERL+SABnb8r4cBm6
X9SXeHytNW4B0FeXGMZuVA2Z/Rwdxz+lDomXK12r+VWpneAunY1aQzuDbH/D
/+aRRbIGpCH5n5E4tEs280cDpy3db79rrcePIoBpYhdkGw6GlwGQ2u4JzlwT
H0dnoL1g7Yq/jcvqJDmg88xh8BtmrJhWyyp2u4z+295rEx0zYPcqoMAPlMqr
5lpnAHHRjl4eomuvEpQEG3kGfG1XyOFhLqr4oGL3gSGuZPOiDagYZG4P+qCP
DnDY1gS7e9h1uPDstrVZLIuUqsOgfZFUigmOtdfrgRiqLR9DcU7V/LeSQsvH
O9XP6ByuAZ5vVKptKoTRO1cEwlx8cemliEP3cMYGC1DPP8FXUApK2uHaaxrF
lO+EjAVGaTR8kDksFo1ZRiLlH/v/pFXINDhmH708D9day/ifV0wRZ6QD+9X9
DW3PhhlpP2sg+rHoOOdQGbPWJDd4kZ/CD0I11kbPUzpojPrw47B48C+oQ5XE
XFnLJEjxP5inogPLhVuqn1hkZuIel1+sD3VaubFIQqma1r6yhg07UzyiFIQ5
6yydvoX2fEdv53VmfLn1OWCa2MVsYF7DoDOuGi3o3v/mD83e9pNII0zDN57/
UFF9UMce8Jz4CYS8oFK7FLWj1jVIHLSoQAjiHKPRCjyUC+Z/bIjJ3N4YKpk9
IHdSff0/l/oGdulgTbq1G1yc37S5abW9l01iz/UtwkWqV+E2aig9v/vX3+AT
ETRXJGtUyodBuxxrDn/m0ez+F4jWUgq8ek+zdUeZ68Ip1deVaIqVvDoDcdvL
YytmHvxvpLU/GNenx2yk9/hwaG1G60S9/uRjd+HeRT1y20E1abkrf7X9jqpm
O7NunOJ41kkCXiPWiF/4GhYBd+4qlsE0p80K2cE2VyVUCzsj7bH/YhsF/rI/
oLm0SaY1AlTffuF2dBjmC9pxT/oujmPAkHeaBkr9Y1/cykUv0S22QYD0IUOs
q42Pne+WanOUl4p7ilZpBp0/EbF4K0wrvM9c0FgHDtciAO4tb1uz+vt/OkaY
IcTyNiRnRfdGlRry/osuztBXIFdKacfVDFFRsoO1rCeefa/9G4uteJKHWPVr
hiGmZpMuz/wYvYK5QgAKGbROEhKpjh1aQqhE/6jYq269pEV+4O2IPsR104+M
2nXo4oZ0SEHPA5OPXN5vWzE5baxVna2HhyopVMV14KRfNIWzcKHIhyCJhHLl
sx8klqg0EGuINUbP+v7CldqKrG5/z2sjw3PY4qlr5tFi+Abpcn1uZ6i1PJTY
oN4K9ds8XoUvSWs/QxFNBPQTO2q+/mqOykmg+PELtie6GYMHjfRhWV0VqpvO
ZTf6zt/wuXsGg4zrR2uI24aFrp5whL+UvM4osMWN+tr8FWcH0UwP4fycd1T2
cTQDwchpS5XxzR8+7GCRL4LkGA1zA5mtIXhrY9++Ipz+JyhRo+PyYdxdYxJm
2zDu9DKcZtEg6O6YTfnmRzRTPYBRX/M8Y+I1Hx+MVeLUrU7BYRtWsDDV7vYF
hddtkCzIFzzxOHPUszM2DqhbATHAYhkXZudAjEHKaNIQ3GVE8gFSLMs8qumB
24xVm24AhBXWXSX9L2QzW0CIuVR91MgeMTUaHSQSXC49I+wS4BxOuQvUFgPj
SbtwWuklk8W2h2/5POKux+a7w8rmabBke5Hwq1UoNnGweyByEQ/LDcJXX9WB
RfVfgXYCJnhm+FB1J9Bg58bdOuSMoqjxHnypHNvKluGh7s7elf6TsecyOrnr
TUGOfa98xavlOrJn36X6AnETl9orSnKgQM4Qdjad9WuYCszLBzo9qEf9kKI6
1osFaLrBI64OPXMH805/S4dGaBI/4jTrYGeg06t38BZPcMKiacdGiFwWYth7
xLdyp3ncPV+6kmwQev6niGD+4zyNWXKSxAQbVEGZ8cRw5uiiCNxdiuUThidy
BTsUx/xP2aVJ+CdTaiAQfDxkXdot55pd22u0C4rAN/opKfpX+RUYOougddmZ
X9nuRll4I9RXgDkZCd6D/ni0v7jvRf7eXCs2vXvyd7FxtFzxy1l3X31oAehO
cyJo8oD4eIyahffeSFnZ5SrgppvS9a6VLqAD2ScOLxiYEOwe2c4hqFrfMuEc
z4PDB3KzSQ4WimUg7RCde/YJhmZ/Kn32GBZ35m1QNMGA5XA0PnSn260jgQWP
Ve0nlsQgFdpjWxiac77B4hqa9ajIifhNsCdvztzJV4pEGbyt8jGyJ/90LRhQ
cxb64nJ7xM8veI0tZ2zx/vtLd7XETGw4BXGSg0Rw2cdDOmD5++fZnXv/4Jnp
GgY3pBtTNdOuTqXK9uD114+AMVqrtFfNeS/TTt9w3pqcV7+Bfu14C4yRcx1l
5dvAZnvtG+57j3o9Qe+I2XmHgqTlAJw2l/SJkLs/TGN5lelOwuIXNWkY2aTI
+t/TrLXJdkWQpcoOaBZrDcic1RAEzVVYpUnOJfXooekCKzcWNTix9/qlcnn8
tVNfzLokzTu6Y/CoeZIGsTRLFaRpR40EqPRs6AOA2YT13sSe5+eeQ2CvMQNL
rCwR8Lmbekj3lFg9m8Lg8LTfXZBVVTQ0TAoeyZtRR8YXWWrz8EOTlxTt7+sI
wm+1DQtzBMn8GChMbUf2EpUguTSmla/d8lo1W4GvuLXdUTq0lWIeDKvMVVu5
cgEPSFw7xJMXsmuMnO2RGyPlysbsDqj8mIAnQnCWUVDHNkBhRZwa47hOxvcl
cwGH7kAjai2dzeIgEBeOXiSWYkMc1kxTf5hzn05pScIwmssSyRxfJ+1VcHIA
EEsgCyJ2y7t4rY5IeXxyTMoEApHlijEKzB9NBq3vxgbaDOxkAl94kLf+q2SC
MFKxUZY9IxkroHX/dT0YBABxcYqlbq3It0q7CX07SrS4lmGEF+Did6DRLZzZ
lG0Y/3Jr85BnYlL/U+3EriGh18C+kcvxsmYacjWszVJSm8x78LCjtZnfRgBF
Go+JbWRlpYgi+gXF8BFOyTnmz0D3mC3+mdk92vjeOTT+P74OMFNdFh3iTB36
+2Rvo+S54oZuDf0qG3PEp5TjIj0akZQalfHu8sQHsfISh4L8iBRffnf1QZzY
XB0yEtttrI/V6xa7T6wrY6zQ/t/0q4lBjfSX0yZrU2Y8OquxmvNzrBRCYRgl
rs5/bWnswVilaip4CtS3peFs0fXsBt+1J1ZSorLoaaZDDNo47ty/mbl3+QZa
D+C0QaJwpaFqDlKWE/xbFRM3Kgs+aA8YgIuMZyvWOk4wFHE5FEgOZr4/5Sqh
EjkH1tgKKGlBwXDKFalCL69ElOtpgporQYr5OnnRnMt0MuXNfqzpzc3fd1sV
SEJ2mwN7bRwNIBdQLeDfH9lpytyE7KDHSttQwW19+jedFpoJ4R0xKMuGVhdX
ZTEvwk8u+yBSg88NCinH1ygqNZF7YMy2UQ32PBJBH3oJZ5MYckDmrJ+oucjk
0rJfEtPs3WxR7oN+CiDhIh//o7x9m4VkbgjvMT1LeNvv5TbO7SCH3JIayhvG
GqJ31506iRPSSuA6k+0ZHaS2XP6O5YxGuWffa+bxmMOPApwMferjVePBTuzh
W3LAoLKdl7ZXTY1SUO94gqLmAvw5fEreymmJHDaKUMnMdiR5+2+T59MBT/lD
KnPOAuvXC0l7q47xZZmKu1F6z5pEf6vaKLlmBJFp2+YMlYq2pOc8OE+JBjeC
J+4CLHisneMXALzqIbbDUCckbNaJwoohmbZpS7bcNvfSp8rCop10H2GXZE2X
D4yJd+3zgTK/pCcChOu4+AlQ3o/nk0e0M5B2t49nnkHxPQ4gqy9UQWRDg8I4
uwSO8Rq2T3q727/IHi1XQfGOzoQkZ92/ntWtLdwqWy5TlpdfVwp5jN84UD1t
BAcaYOZroeKwoZq/YjV09Gd7SLmr1eKUHIk2bIzDQ11386iJl2KxBLpqHlyw
qS2bADIO1auJT3h2Prh7aqoUCOSF+eWO98BJhCNatE0P/YPu5ojQN/z9Q0Jd
LrpuIBb+q+6jc2Mm7nCOiexPs8TP0xVmTnXbn/0pSXSJsc6+pillKyjWJ6bT
d+580zcabXLShq4EpsiDxhuHmeK+/FfswzIIdnylGKl9BoawPpoaIBu8tyzb
f5pmX10my282mGpMoNGeFTYw7D2jdyZS0Xq8U4v5IRN+4bMLeBf8C+h3KBr4
tRTXPAUFr1SGvs7wq4ulVEc0qX3XmvjI00rHwJLdQ2tm0BVlF+GeewLpjPil
YYkdN8VE0ml+iis1FADZBQiwDNUXd7jeJqDHEpQmWTv6cL2Qi0Zdjlvi78IO
p/YJklieRfzBMf52dzROkaYFuzhVEQvTLQgIBQERgyiQHBhuiRqsQuu3SI5W
szmpQEkVvfZ+BPVeV8Ne53u81MNURo7u6SVp1eNQHzmHk+MxCKqPgQcYSJyc
z+7Izs1lKt4wj+METK0uA4uQeTf/bLwb5A/+Tie1xOOR2vekZQjGQXXojZL/
Ft/QNbnm18bd11cbB2GG7XRAFe+IKghD/y7sRuATUV9TuTWcMeSYUzSA+aqT
N1mTtejPmz1oi6sPnS65tg3ru301DgVW7dWUB7Hj4Mg/X1ikxqv5UBMxPztK
NPZpPJmwkDULsqi3FRFGoqzdpqHspdSBjGgufbwGvC6xjh1v/Pbee4GR8YKI
R8+pEcS1qTip/0JG/Ekt9i8aHSmB+zY4Tv8q7UPsGggsiyzFmGRqYpSSZGG/
EnmLOGDPBf1TGbPe5/ZJUVz+USnXuhvzgq7o9Vl3MLCBbuImvk4FVnaG5if5
g4g6LPCM4s8YguR25WrvnF/qZvraJXE31Z2hljeKKkJ7vOc72eCamIvKThST
mXzeBXjUtCzdI5X7Vo13BmrJCVPkRY5oRpRCpDdSrkHWURBY9QBCJznLqmWm
1rANXhAdS6JfavIylN728Fv6PXoshCgeUGmRRsg2+TOYcG89TRHRb1qGNVpL
tZHVPyV1We+MirQbc6Vp3Yja4nl+JH/flRemTskZzurJBkSbtKkxUzFMJXwg
GQfd/8GDBo1uXI1YBNrefls0NGGlwfp3S4U8BdmchfpcOCF9xhxY9xCDxMP5
zf1wDwCWzh8yav/zXBTA5Wac6Nfyzkrwk405CDRJYHbhGY+bLfr65SWmu8gq
Au5g5W007kXeClk84db75xqftchGaOKr3ljXGK64aBJCE4RavHDmDaljp5U7
BYfTey2nAPTF9xmv9gFGtzKXdSF/IPmz20kSG29FhxYECDk7cKhJ0U90b8YE
9/ITt93+BxqYCif5IEioC+7SdWFpCgh9hBQKZMZPOrDP9fVy7AeiuhluCUY5
kOWmyycWZZkqVzld1vdvvF7r11OrBnMWAKd0PKBNYEdt/4If2jKbZ9O1VFnE
Rj/VR/wmBSKSystFv9Ibg3mzRKOqp1yuiLlS3GTslEsxiWHxDAVvf9xgncor
X/zbheEux/wlrOwtguTYrf2W5628aGtpHwq1cRuZCBi3/LUYujGZxDWkvVrd
GlfcD/EloSkiOn72g0R8td1TnT1AyZk8k7NyrSBz9RT27mRnWXO3vF9de5ml
fTfeEKejZagcd1hwJNWGR1v69MDAiC2yxeQw04D+Z4F+hG9TYYyJ52yNoBH2
k62OZgX/cf+xq2Sp2Ae3h4L8dnxnK+jYhLr0hSU7ux1VXsyD47wthZxgqJzr
KlgaPw+YsbLi0NsGu4tyteUzcFHnhG1Tqqydgtq/+2RG0KI5TOlKdoIlUoIF
SmKHrPrOyCAJ2ripYHUqYKMQ9exV65adWEFPjSJ96Kryr42mkiMxEhLwWEYf
Yh/n2hPzSgpQTjSvttiPJRrwUDAjQGa1B5bb5Z1ICWLiS0fTSuUwDgnMMd2y
7OpKdWZ+BJ6ZqtxT852PI7ir7xQfQNGkXcNlRLGqTIu6gKpV1tziVXqY9Qeb
eRDia7ieuWuxSWLDlv/OVGx9DPfLuVxp+eoQQPeQZDkzkUBFr0VSVAx/sw1q
4YOfZ5YpWTNCkniAEwq4LLvRzIdKrAvqsbZJrwPD3GpxsiUnDpjlVrdmkDBG
naRK3MuM4REDzDnkOyOOjrOiG3rH5PNWEnPfTwU5KEzBRixch064L4U2ynF9
Ztmw3gzCpoH6vjnyGzaEawyI7gObeeMX1DcGGFNawvZIMAy1TEImdd1vA/Wo
C+2gN45Gy4tBqZ/8DzGcomt5+NyNQk9sBVv7GzB09ur1IXbiYg4DleTnEvh3
KhdADK3MA8mGzvqHQm1TqG1/iQHsTysVXjaNVEUfzhW/RbdKB/mvLdBCKHbf
cADOWvi46KRgl7EV18pfNW707/CLI/zsfXZxyvvP/syErflEhS0OiAQZqyyO
KY/NmfOLMtZdjn9+NlPyQtmxqJeNKADQjoqBghBgm4ejKGVzVJfeQuRcnbqK
SuVoE1yLGxk0ZbMR0Vtvnu6bncRDHyLsW2sSdJD5VkhjumyPsvJRAAsurNox
Xd3l9goJZ17q4KsR/MwZeW4KcyKmq3EmgBaEaExmi2h/2qzxnX2pMjQ8VAHe
e6Z5hsuhS1r597ZMWsRtlB6vvBVq32vpxeAaSr/RuTc2B/A1ZBuIl3w8Kx0j
wtocZzvV1GZ//gFQ9TfYJjgZE70VpARaaMX4Lj25h+Q5vZtKl3PkFILUT4VM
gAFkRRR0s47vWr9f5hxMga7OQjhtSNSsxTUaF7yaoZgzEXmPzcem0alhBfB+
LqPyLr0rvOAjKTBQffy/S523lTTTAsIsvtJbpwVFE8CraYzV8HSJKM/F96GA
g80oqjET93d8xfsE5pJ3fPvoiSkW4P0OwR/0O9ujA7dn26jTvdYCcoV3oC20
x3QySTg5vrYFYC/ui+onh4rpSwbDf5CclbI4fxRK+pBGqKb/2fX38ISNT4An
fn3M2DsVIN6ZrSv0LUop7kTAh8X1dqqz8h+xgDyCo82gpyKP4WTj7FbFglAr
ItnUkCjIp8dxSnGPpqqDWdLFdm7p153QQ6VzO+KpzhVcmp1u4pgpNIeJyIMG
t1I4X4q/A5w+XlG2Ym28Jv+Z8Xm8kvW9/88Ff69+8fGQBK28Kgd/YJIVy8bg
yqCpQc9I//3nF4pM0Gc5qqUt+WUtCuV9U9XbFn5PYGdXp+gpHE1X1Z3EFZ0+
o5MVTqjI20iVKd7waAi+oKLI4ZKJWZe3blEwq6xYzfIs4IosdAGOiQXdmSGw
XHtJZ5FquG6KVUrWAzrvOVL+tsM9AhdsVOtFh30kUpySAw+Z1e4ud6Hp7/tC
OmkuIyYxxUN+MLVEOUF6sZpLdPl/Bg73yu1+sTsl2kk+g8uOtQX4YQTyCP8U
AaUeF05nYvzyF9pXnGU+aK5G2pAjdU+fVaKS8gM1W4qEtXZWH20WFGIxll2I
SYYky2Kl+Fh567m/xP5iB1oBnSNoAimxe6qAx2cRKiHH7NCgKSbNmNe9lVwB
6MG/TLIJBwmLAfocFgKfJPtnoHnh0VnHMJAlIf8FQnPkIOjKd/9Ps5UZHocF
5uuvQTSHMNCiYcm5M7JiigC8VFIK/rjoN5CFKgISwFG9Qua6dKWvf7S6HdII
V9fr/elq03+MIyt1uMNCPVCuGWro3Aq9aCzvZS2ObCocOLaj3SAtqu70c8qG
h82O8DAjAK5MDvgonmpRiU2QRlTvTJ3kiRGaDbkjmctAQpb08bjC/t/az4J5
9YHz1Uwp8K15tuo/sjMnHyCpPnxi8Wp5R1jKvkg0FWrnSPp54fjtaNVkdDi1
o7PfaeS7FGEXZ8KJeateusTVN6Gt13YXgnn+1dHC7fS3BHBkANfZt+vHFtEZ
bES0pfyEzrOqSdL9s2B1njSM3dHEQu3QgO3V8U8xEAACx1IKawiuc4Mk3SAo
xV/SqpV0UIemaeDcXO+btgrjIoWfLy3R51SBoDQWkLmQnx7vptF8Pb+ullyY
EAW7qdamSHNVX2Vyeah2ZH9jiG0w3vKdMdwVPHeLgg37elieeW+bgnUixnIs
ENy5yyifCy2NpO4oMNAGqUewnhirJiOodDEV3Tyxy7k+t48hBBV0zvx2KTY5
D41rKxFKYM8SxBNAaV75rUZKbP3vHTY1lpWA5gWMQwP+wQ29BEkGmWKFM7Vo
Uq4A7Lmiyc0ynnGg7sw1kfCoAwf07Jh4muqYEvdj9UmOzro0oPUBM/K1numc
kgvH73UH475HYEPmoG41GNltz7U5Bd+3brUe+zrREm6YS09+NeEdEotPdDxU
dmHZMFfnEFY6ZQQll9PFinLJuCuXg9irfFpdqzubcZZp4v328XR03Jd8QH8R
xJ5sJCZBr1Ja09PdNBS4Lk9Hx8kdq0S85rQjK72Ct4gMduhWcqeWkX49nOOf
cxs8yO+Rn/qZobwa49F+xGMG48C+UpWVkXFTlXasdMpiJhLx7+Mt4u7oWhps
HdYRlaJmib8TCNwcmYO9X+OxgNDMomfWiWsk/boup2787RzVay/f8HWJ1ZGB
t3gMrfRvi7lJFwiok9w5K23T7aChdAzwzjqBHtsGUwg8qKnEHs8y5K5qvBof
r8Am7RX3z6MyGzfnm0vwDD14rQDsr9825erCkSux6BgA9gJsuyvNcPu5GozR
yRMruyYxTWDPH0iRwAFqidnDOyiNucRm9pVM1sqmdzqJH+llmEt/qWNYwgdg
HVuSw1y6IQAaQQ/KryWBWVrTSsPKf+OVrpINvoymmMZGjWHXlOYstbIBE8pZ
5wSPVyBB/FcxY594moD768HmtZmoPvb9CpQ7m6bKSCEU1DAAEsX0bml+HnZL
uAfLHNsZAi54dZwaHXGW4THHoap2+PCRnvy9b9sxBXJ3uHhnqkpR763NZn33
6brjuAv7Ow5nd9dlBAajO/c9ctX0RW1YwduOzVG5tOyP89mkAVi2qARshZTu
pxA1VVYL2JfnlNZWQbTQveGBC05K9uSnu6DqJ7MNi65qCSodwe04zyIFBBad
OISn35jVnJh1zmnTboiLMK9DCPj3sHQy/481HUpj8WsL7N6eV29Z4W31Wuxb
hcb2f8R4aty+fFlcv1uhRhGBA2X5/y+/ceO/tdx29XFl9CfzXps9ljgtO9RE
pVBGA8/yYQX/D93rUoNzdpWz16MFfBUq+uCAjn82w++aRX0BYzQFIsCMLvPk
ZRb/kc8p8M3eDFKyxsEOBBXhwSZRwDIZ6/jcl882Z6o1kLiF/SqQj9SBvWM1
dpKKgQywq4TLR2UMIgUB5dP9coMqoYcLJ9lCmCmNQPrJD9aUUUcXPx/C4H3d
iMI3CfjfrA6jqxsoZbf4wSQzEcUtlS4uV4YFKjMkkAQQBOcpcSj0O3GRTDl/
YOqUgDtmkzYQ6Puxa3OrxRdaGmBUhhWy9vLMs9I5lQpvkFsE3FuOcpJ9T8pC
nIsgJFojbkR3naTahyDyCMiOzcZxd45CYYCuEwVsnXdjYtHwm79LgI9ionur
8AMGhlNTL21/cW55LUPvwDCElvEQI0OXPHAvkM7e2VSzB1HCqqeQDcykQzd1
o9aBlDOf+UPruhma9YwHl1QxGet1pzPH7yHvyPulguCo2gku7dKi1OgDVp8N
4un3eiEb8005NqOBtnQxgcXYktHE1xjO2kLz0j3gKYshwzT6EFhoCAHzq1he
dXmKPqQwQP4mjZvIrEztrplgSTXOmDMftoJoXQXSGmofFtPmnbElyy1thSEd
WVq8jHQBuacWSlvNoUxM/lAnhHmUzigRMf3NO2JIgmwpBEAdql3s2p9n9xaD
H4+HPZu5iFR89qWdpaUbgKz5vxR1AWrS/3ITsxll9rysEAKojwXmrt4qeoq3
YSIHtnh4//IxhpPxEToksf/3XoUIGr1AYe+oqBVSVgOL4uiklzl0Ykwz5H4s
aIl/rOMy4nRdEA0BYTd/jlUg1s5t54Rm6Ouw6cO3yRTkN+lbndxRyYmxL7Ly
ILZ9TDtSvOB0cnvLm5vBFpMRigWZgMWUi82ESZqB3aIR9jK1YQFPzxyveFHw
iU1FZL+V2jo1akmhkJDGUzvuA5yuZd7QhVMi7qmBcoJHj3Dtzesap54G0yxN
/QdIS8KLDvmVoMiUpZQrc4ih26eYsD1pjMDQoFeVbgzMsrCmVonbf4fQowNf
NATTbBJoO9zcd9lopaCXG+/ba+C/moFsc6xmssNYVUR0tPpBKdMvO9eAVPEL
5ylB+N6edTRaJmW8Q4SLaZtTYPn61ko9Z+UjR/hKej3hSbNV2lQRglr4N406
07zkFpJro/JL3SlS661FmradFO+hWvQ+CU6gKdnI8zjv86GVmbfGw62aa1lW
sB3l0XdDAnbGxqPt/iJN+Ol0XuAuoAU6PffxHsQ4Dn7yTW9kB0PSKR4WkK45
UmHKXDWG1PoMZh+j1qsqUSAVg8Auc2M1oCk6NwHFKFrqpNP9jGimNcrMw9ay
3CJtOCU6uL+OMM+kHldsNwWETDEA3x0mXNmwGAXN6vUtLxP2xYrXsp8hNpc5
zViKBIUdsEE/jegAtDj31KELU4be16eosyNibP5RrARQBk7BYyRCK1TM4/YK
bRCmQ8ybTfAr87A6QCfdRqwOhXHHmmX/elxMQ1Vpc3ZM+rWnMdenXZhoV23q
mT0MqVyN6IXgALNNSJ7kdbawBoTU3dOSCZV2I1HWdUCzWVa6MgaMSer+PBrd
XGQsXn5UOsiiFPjHUTeUqGSBTGCMJGKudLWqsliDTK6m6drJ9Sjh+G9lN3jo
l6VKer7wQfQF0hgJT7wZJO/90oGyNFqJMI6yzM7Mb4Xe6IMqMv99EQzuAOFU
3LOyBv7nvLyn2FvCKfNqoZSbyYgmy6AiBpaDxhyWLuEloPtTUWWpOuDlGVw/
a99dgvj+Y6p9koz87BGY9f5WR7BbupA6hedmX5TATx0L/c+jNlPdzGZXVU6K
CLE28u1StPOZpQSL4XjBKbd65+p9a2jVRn7UVB7AC9Bv7PehZbUKGLRrpoRe
LbtsHOsSKF4EZZce/jFY1xEJJtZ49xu1OX4m3UqRSH3INN69k8tCLdXqhpiS
QRdYesAOLPcrWqIiU5e+L8GLz1uzbjxP2GbffcGNlvkqBk0CAfKTBaxTP0b7
XMKmZaVkBag8buBRVyyEjR3yrrEkvqCiU1OS8RBXY2Z4zOJQXbdPv/bpuOvV
re6jTyFPD1GRDBofZcfbZwj78t2sKmyNc60JroqNkkR9TJFTmPKwepAFHGMF
3e29hTqn1VaocwXN8xlpeWg/SkfJb2ppIUpEM8eI6z5RLlMu3muOr6PaG9mI
RdbOskIq1dmhEswNIZLOycCYDdyrtaf2Kgr17/VOYCp6nq/dpqO9WtuoUL2j
TA2zKS9EOe399hPxqqCf6yyussKBZtjvmFgw32WTmbm3WatnN9uuDASTOK9q
hI7mBzfk8kvjDLNiEGmB/YlUipvtOQ7Z1g6yqWtGNPLkBmy6UxV92bA2qxr+
u5HMoNUSsP1bK6TTCZKQOQXW8XGc45T6Of/HyvVW3VJFuYjLyAOZLR2Gru4C
MOndW6eOE3ElVtnq2bmrOdMC1H0fr83/5pxdB9TjLrKbLlURPBMDA/juFQwT
CMc+/TnSaoMyw5u7KT7OL2jM94YArmgCbvRIi+NnsIa77ZTJFNlbrtV7P/jt
UrdP87huDmHkLXQ4GaISPbVnKTqOcFHGXc2TtGPm11DA4AnexIgKUSwtHS5Z
a49HCtat8V2EcdcLazlhx18FoRYGckbTV1i//TIJ6R8JyGg4roCT2yEpaAg6
tgJ3fiMFkgg3b5Vp0e90VmTtnH8ewaJ+y7/YxnLg90EaSKOBufHknY4Aov2w
x6SIjjUQumTPyw2Jg0OGiTQKciaM3czHdY8dXifxkDvREVMvAo+cOuXYt2zh
qMgn3E3HoomvcxVpf+LAsw5VVpKKWnsx95eeHsqDh8MmFinowCDTAZ6cu9Tk
mdxMhcZGrYJ03740XqSssC0RbspmPxeAJ3FK2bzZCU/RMI/Dl3ZUeUeBuTot
kNEWeoqo+UqU5FDFUqQca2pJbxoSFaOburaG1ecGyFbglZwP0YmL1XyYGob+
34xjLh+muWhCG0cBtP/BfaLUOkrR7ZGCmyi2i0znTa+S9EcapNgsthoXnOqB
bKZL1XhGd2MprqB1os93T0vroURbKC8bRvCczF2hR8R5VhbXhA/uy+BkBkgF
l7txbeLc5Q4gs07WWwtG1KbdU7Fo0/wjLw0pHcwb0d89pl0EzjPt73OBD3CH
1p6Ue6O1BrfMUbj1kL2nPTIKhAk77/QGRne90vVSjzJ6sRw5b3cILABHlZEA
tktKbkuxJJilD6F9cZbYCJWCAievWkp0PNT3ZmpynGg+jUcIDJzQxrMOZ1gq
1M2H0uiYMVYlutFb9lXjoN6Wz9UUyzZAu7yvzaq/31p2u8NvXsrx/H1aWOWH
oP9nN011w7bvgSfBVdGTWZclBRGZsHi3qGwYp+C8cVfNZW5QmWlHSQb1W0Fl
+nooLLkwNKwptQarPwJFvQzlyJCEVPESISpIgBOxUVh7Q511J39WBvLOyuuO
8ELKkS6hLhtHY+u9P/5sf/it3WFkyYdHUsmdidG+Ak8r5w4kDN8dUutY2bki
oCf6OSsOijD1fan74e0OvOJL/PBoMA6fQGmkLnNssfdoDkUH3dgpMsv2DMYd
+jcv7x8nKyZRqAOUXavYKvFLp6yydbDBC6xe3jRBIFP+ipFRVmbCJiK6tuHt
eytc3hMfeGsDyZOAX+uKRHgK/ipsNXiCgaC1XSjiGI0NNdnO83sZmsoXbW6O
/Rob7cuRyXqQ2jeut5yeVxLj/2kRxhunOodX0UKYSPNHSd+jpR1sJV73ldH8
QHYBNq5WSoNcPoAQ5HdWIC0hBoQxPhNIhfjtelFyNJcDrVqjrumiQx8XIE1o
IX28goYan6+mf88tyblaheRnye170tdZnIeUf1KW4QsuQCuxoRmcrlghsq2H
Uzxtu/ZMpiD1YVJM4u5giaTcyarsHOiWlJNqxDx4s/3XaXncqhO/m6kDMfrM
mCy5glAeNQG/TnkJbWKBVl4IPzve7hvq8k+H5AqSlYiUNZIfXX7hfExDn7Lu
RgA5BgQCVDBqr1zKMhUbSfe+2jgTkYPpZZPUAa6mz/+vexxNu7wDsACEtQoT
9Kz2e6M9H27aAAE7Vy5PtHiEdkhrwqO8qwfq0bs7ZI1aBkE3Dex4ybGvzRLl
cL3NPR6y7rpFrmWi2R0KoSZJrTp/Apx+NRUUxqsn1sX3IS6PBdagTf3v415H
lZt+fhPqX3kpNII620XsSr0rjuqkqFcZ04QMHqoBKFkEGNdIt9KKzOSyCMBN
kCGlqPq4g9YwFiS4SiP9cFxuAbaQtWKC+NS05xd4vdwYZNYWeZf/Gv5fjY8u
UVqu6Xa+qITmXkSS5zLdVjPJZ/j4CZmG2tM600qFX551+aZpmqUwtTXROjIK
enjvJwasa4Cq9PlgzF+W5F8xWaEO2H3eV68Z9AaGo9fgS4K8pVV7nGneOfCh
pBIJYnoUncqeeIRAzKf8hLwHAg/jPbt7awE4gKWOGb/sk8TnrgVi0pFGBFZb
F4nhUvcM3FiIk5vjx4ASsyUMpmpPWqIhJOH2F1Wc1ypLFqb2t5Pj2jw7EQAw
CwM6ZgrblY9Fsl1ygWIOtta6zWJ4oUKIUjTr099gvU+JXWfdqVNS4ThZZTGA
OIOQWSmkAor8HCiRsiRfCyRk9RZi1XYe/QonWXXw7QgeiVpg7/h/9H/e4TAI
d8836owoIWWzDnw1lEW8QfFKTXYYPvog1UU0uhKs0BGL+v/A3RfJljdQAkIa
n2tKVSc3XLFyfavyigt/wyA1JRpZPx3+M/rMsXxc067hKqzmGUsiEt5Q4OZb
x4bdojXMBoOUoLM5HYaMRdj1mUUMHByZuUbhK7QWs2NX2EvlWJSyUmbwJN5D
nLDFzT21O+NohGzt4NifeicU58XGRGmTtymmsr1PoBv3C8iWrA/6X6YlO8eV
l1EB0irDqB/BcuqcI1ag3LjBQq/V10yaJke0DCCx59kptLMMPHVplMUVjAhQ
HKLkDPFOKfNTAhh8o21xBF+ReL7G9W2DGXx9C+56raYx6HDka6GmRUUEalH/
SspMuNWsCN0a777u6+f/znpnVXKlQ+HzfXmdvRGrVu9l4mPJbcWxuUdnyJZB
VP8bJZrNMWqtL+vZL24fh9YoU1vrn3Ym96h1tCifsbS4dhlXh0z/UJqL8QMc
7GCMy7bJLQsyIBSZOVsuhdmN/xN4NLR8vZcBKC1s/VRseT7tH73qBsaNhCRu
RO8mTOm9HEvupYOvKkhmsovfuNjSFk8X1FC3WR6pxp353oueRUfaIJp02U1L
9tVCnpmV72OIOYm2HJs58Zm2EocmEfa9ymvpgpx6c3qfR/ndjnuqbygwyBfR
LNpP5OHZU7u7PozD8ziSWgnTPZ4jY5+dNIzXUmd32WmvQj7eorfP6dAG3iNr
ymhZjv9jYu8bR7QM9aceLbfwap/2cVIuF4yHYd/7blXlzoRII2dpPIaEzOqS
bG0ZOHvFtFH4OPJu4HCWnGKHm3/wfqOtbHV3qlPvoBN3JuzAyCj7n3vrve9W
qqSDiBJJUShjy/Vw09NyfnOfYuEXTX4EIwx4HPswoB+x7UjR17fieibr0+Nv
2MME0e1HNKPGMWZnt6PF7Y7nPJi7LqcbUuAwfB+G6M/9dk8aLmSg3iAwCTU1
79uvQzyUdiv2HXARA6Ugn/0xjUV/vHVnq2TjvmyucYUM2a10EKNED6nqakl3
VawQF4atDyktFKdgaop/Sn0B6wR4Ad812Es/Po7oLshqht9nMUdpeArbcOie
nbcj53UgrHhFQYjj1EyPyuTH7xgA3HKGpMThcoSB6LwHt62tVbg//KWPeA4q
WEollYzTa7v/E18C7foyc68/pW9vYKUVHFCjREwx/N3VUXz70xf1ZK2vTQtF
sZ5Jk0pMmsQRdB0DiWHq2ub2fENUr+34M61xk/lSJ+0MnYJyXFIPCqDVhEZw
L8lJAuOD/7OAuHr0iB7kWZfOgl0E5CH+s/t+UYB6FY7jlBin25TelJRBxIxW
h4i1gS6OXWvpsyfjapDrbHotMIxl6MG1soIe/Z0dhBIF5qWnx9sU5Ex6qQ3H
XJxejNJ67T49Ra/mj12pCpJqx+sjEhYEXbKLv8HXMQJPC/8uJ7m5k7TUdIKL
tbpd4BlcYXnyQ1NxBYe2ekDMAxU4ZHvYDJC+foLbmaXfAcBY0ZkKcsaHuljH
7DI8jLmwD9Wyy5VhPiV9zxylFmTbUOEtnAjpkSfCRR891CLTOaE3wUqt0YOb
+r9iIs6L95u2vDetMhDJZPuVM1wq/Id/KIsvF3HCkQxMbjJg2RxA3BroX8Y6
L04HdPXfnO0jqBqiA966Wx4jZjbYrMemFi+uT3TSOnMjwPgAFSGoB3n5fLCI
kOOpkmdgnYPfLEzD5BvZq/TGFedS0EuIA6vC2BluZ1fOA+tKkB/lkBJ3hmG5
9vMfauqzQFcomPi02Dhvu58y2ABSnhkZbHTpKvg4FUwSsUSKOdxKQJWorpoK
jvgw9LPoE3svbBjvPKsZygSq6/Qr5O9a6oC/bTZTz2whyPh40UgI8KbQ65c1
mZ7JSCaVWIECd6U1QgwepdsVwlvksbuAFJb2xr2r9D3pbx/NA3IBaF0MDdRY
yIQkl6vTRPxvMhCwgTB9XDiCa9kEAd8fhJ4famSEKKZ6pp5R33714GCt952P
O93iMF8Skgjn6bKCqgexG683EmOqZxb5FejuzFUx3fC1Zx73AwcyGc20op4g
6a+Ifcyk3zo2pc6PfFnU4sX41rN1cy5XxRr2DSg7zfHPFDaYwRGVVs6gZjdR
KiWgNyPU/Fsjo2pleyypXHTcnCOrmtm+fuBJJxeYuerUPUuR5m+YfvGQnEDY
4bYHr+BtKGQBgeX7PE0UPs2/aFZYpADWWws/s/eCvA42CahrRQ1/pQ1ViEFU
RSDw9Qf6FhvxCWRh7ONugEyUx5mmNnNhIag/0HvhAq+oYDsKIY88hiv9jJ7E
Hk+EiigWlOblLqf/2G/NyxX78Htb4Y0cL2l3ZAUv5BNalIygew4sQ0DAS2GM
KfATyCZQTzAnJ+PritQuxskis6fHveIn+m8OQ396KESxKtSepvC1Nn+Lr9TT
2cCvmckVFJT/YG6ve+2krHb+/ewo1ASmCwJ7S1nx0Q2YoksaKQYifP7QG7Rc
V5sz0PxTPYB67RVdb3hyJusDt/r//O8K3Why12A7VQEhM7KSXMIiTCQ+pKCd
cYaknCHend/bzItrhHU3o8GVIpR7ncQ/wmQuvhG0+XxLhZUrMfgdqUd3q0dA
KtK3JU+4qClHlMjqaOm721lON/DA7UxcvQGza5rJAlmfwd1hM2AxXrzypVKo
GY1nKLP+XY9OBfSpzow8JeyeM+V9v1BYPsY/VaUytVfVXMK4aMUIQ3tVVap7
YvPWi4q1AAd4QrEhjoBDi7wTgxt4/mn5ZcT1KTbxGEiomsm10Et58remUVNc
8lwqjFclfKWsJeN7XaQsd3Fq8pfqXrJ6F6l38Vbx+iyIn5NndelPmp9lQpip
UIu+uQ2+1CX3cYwclyTXoua5eSaxSRmBvFOcdAejyo42l32bbmoHdXJQazQQ
JWmfQoKkwY2RhFgdICiQMpVKL38U+0wtnd1eB8u2+C8aF7sG0CrMFzhituKU
G4laS5xEpXksSdKHdtvAiHyxM+91TyK295tXL96S7muOTwMZYdZUqHFTcuWz
iNHSh28WCtpgPFtLL1aahtOvsJRygZd8c5wycmXUms6Bz4qtzFk9BMnxYh5q
skAv3Ns57N7CcsbihpQhraJuoZVXwwlrU1lyt1cLg+cQYuK2BIF16VeErZ3M
8qz5RpbaFI5jPZaHPVWhJbidUKSNCMV7WoEE3PNldihQlzwnVGlgAlTjE1k9
Xx6eRvCL09wzajxbFjiGIgHEmgEoBLTCgpkkaCzxBlwfsPMNwxXbz/6RbnCn
i+QPQIWevmDM1cMV4f3uUF4Yd2IkqCKCliRzpo6PHvIlJtCddd+CuzNqJxgr
FCtRxcusYIXkoYlN2Ktk6IRH2Au0Cudb2WoQwigvzowC9i0eHydL3Y4CuZtU
4Mb8T0T6h/hG0C8DedguzgAPp5Ds4PeAwIsP1jF8FiT4HrfD8jXdIt79tLuc
n7O6QSnaEvGGyDN4i9KyqvbVFqUS7dH+72H1Nh+G2hpBvXNqWeoMUrYruQ90
XXOW4gBlwe/rEGE/jrWrbAhwkDIkfMQZE9GGt52uns94NWm0Yfa3hhUDiPlf
3xEwyayo6l8RTzoUIXBADQFjAJI9mXA5f+EF0yDW/5N3TjGoWP4OGJI+1MAf
8J4h2dwaFh7z2kUWXSgfEL5F4OqKZJaJNUmBqyl9zTs8Xkr81jNypMD+7Dyl
1zNpeU6dGLc81RAHa1neDya36kNHzY4CiIiLS2ZKd7EyhXBNg3toln/I2tCO
wP3N/WEDSzaXpou3ZTFnJ2noVK4QILZ31Qln2nHddgAtwI7dem568I4ywzVx
ZHeZOAfWKZoNFo5X7v4No0fWAteDJbrESWeJzCHN7sZ+fDJZhe7FZ+HP1Tzq
bhpGA9gFdu5wyNjVjXgDzJ2kXLkY6ui9R5OkmmUrtls1drPDeibcFG75sygL
Jt4S7b37xf427UNoaHDzIFwZQft0//NeNu7MIvinLAR2lWMIBLAj+8NuM6Jb
WtRNGgfq6ip8LHW/ib240EGVkNLaR/GRbVr7gJINI/l+MurhTp1WcaK1/Web
qWly6bd8hBo00+qU+AOhexOFNQuvh4UaIu7HmFcy8gKiIT5ExCi4508CPLXw
O7crdtVQO7x4Fr0CU4VkAudGMJBEXDp4wQ0hcqkQpV+PQiGMDOzYbNH/N7k5
1g+GlrCr9bkySv849D3LXDFVqMmWkyOPnx9mpcVCvxqn75BZwLAatwopWodY
Mb63Rb4eCq99qifzfmFnRJjUgeizFR3y2lChddbO8umagjym1cBHMMbShy4o
6AG/O18rd2A+ElGfifqzgQF1X87rbKT2LtE479UdUo3HlQcfUZoIE1e2Rxw8
8gwBN6ZMfYWBuYxb9J7zmofgjPZFsJvng/WVTetQU++1RsUKt1rxYvnXGQVu
GHKE6Cie0LtD/BZIPa7DtDZv4wEdUep0hbYV85C01yQdEisWVGhKUriruZDp
PW+prwl1lq9r+I/7Jyfb/d7Y5LwdElr/6Eybsl+OpWbxLu39lJz/81vUzSCg
YBl6ZtWVm7w+fTiSIhQOfIqETlyFef7yXYOMPTJ5KO1yMb+9ai72PSN6TnDz
3a+oV9i47YxqGLhfLvkojsX38hInLYQ/B9VHv0+px+zPEGnGEAs+bvE9TD1e
6aGQd57m/K6424I+KRxViaL77djruAEN57cFwVM8HnnkUySw0RnKcCl55iHk
GO9tCfaBi7x7F5keCX1+QMBo7/4fQBoh4Alt/xnR46cIpQDzhH1zxvpqmJKI
foda9yqsi3KfUzsSgkwx04/HaBhFRlTjzPBS6O8m4tmqSZfjHrPoDcEUPjkj
+SUfgkKLuvDWY4rQJ4wgzx7unWY3S4VW6UxavdMNvrQ5wr/yMwpvoCB4ZVw0
S9W37RMDrwMTpWHFuVTTA23SacsoboBhvuCBMezqoOYAzFuxJ0XfY3yRQCjM
1trBG7F3smfNbQ3kh3GnG8PiqIEkXmv4kEv5Qo99iJcI+S32TkDTqitVZOyz
OjJ2PFZ4Sn0hx7Tf3NYETOyxKt8PAAFwLFMPDfcyOw0fqhHuQEZATBfEa2aB
olkRsuWkB8scOPRikfbNKU8smQRrk+8snqxfXdmSrbHirC3I2k6aMhHlYMmY
p7JaBqJcMqTUmf2cyjxzUQESuLrmQPL8JaLS6zjxKWrXUm7RvNQe1FT8NSme
umbNXf8p86DV4+lhA11uHTqSHwaGpwKnOQxr9pJh9jCD4QXp61IkUWSiIO3E
R08++UwAyU6+nuXH5x11c2i4S54+vDS29mmcdL67MGivqagvTrBNuyDxyEc2
/wUDSXwZvRnAQt20grT5wxIM0w8sFh/guNERX++v0lbGGCjyiIkH4gQUKOhl
RevjN2/OVCu+3Uo/X0HQJ8/4R0BFx1IyAI0tfKMuqrGN4qD0QfJJzOvSfGaY
sOqn//keqd/JLZjvUp3g1e3r0hzPomOoKPsv8T9nZ1Kij6Q2MTQENUghgSYz
piOcGALlgspIQSyX0PG1WuEuRDn433LcaojI/XvzQUip7h8U7CzyTi8SPmv+
AmP+kAxlGB9+vOoEgzz1+te17BxYoPeieRnOH059GFfzGspH2rCxdP4QVw5h
VX2x402JWbSaETO0VoZ6GNEB6Zbwn/5nRpv1fc4pOLyYeTRcB1doqtMqNg1b
Qnnp3PSMw0O4kiou29cTpPwWsn+zNvVyV/adU0Is8SHrCJdcZDdrYUE+69fE
HJiEEKIgJZbtOsGaSIjou4nXkYEx8zrWXT8e+ktRkRbZESfDMmJxycUBmSaX
BqmkmudD+XZaodSFi0cKE6c6d2FwAIo6Pad7kpT4Ze1VRBc2cYpqitfQovgK
yODGRoZsbCvmyDQewqtJbU3Kz3QG65okP0tZNXzwVdyYfgGqQZbntluQd6Cz
TW7yGgOM04G0p4GYq4H99QgQaRvsQieJZIO4l4/BHqEEpqluJbO1x/bnWZY9
mBplQ1po9yTcfrgXncbDoE+BceZ0J/7cusiOz9TSOfZBYzgk390N66H6WJUh
tt0pmeh0QR5leMyaL9P3k8IpRX3ZUUvJLzROje1lXLoStHzLyNZ0KfMOVgSR
6DSFyll07ogihA4xoRklsXT6ttavADn2RMV6Kr98cJkwHjTHBCBKrGu0ey8H
AmpSz+9o2rAhLA5QlCWNhKGsxBFAX7B1gZRtIYzSb3hX578K4SwZIWFKO7ey
RttGH0X/9sQOCm3BQLRAFWIjadrnZJgv2xXCndcsb77/0c/rJpoPBnrbua6K
Ea2cEk5iFOQJMV9BCmOd3+GMUx1cBo7L2c6DKpoiubU3qLGkFWFH/yNX34e2
vuEQMGwhjpY0Q46YSiAYpg7q6VR7JlAaN91QexXSFfzcga959j3vUcbNtoAZ
VJ+9dqIoJHqoUu/1AlRswmWrpjGBzf7SRGIGDKjbdpYeHOeOZs7NIS4MOTrT
9YnkL6n6Fclm5dD+YIfGkdoYKiVEe2PLfjySvsQQQgSE9oIsKRFCmKO26RyH
mSoXeczWLe62jgv9Oj1raqHqqV2e564WLOc9hmxuCkpW2Tc3g7R4ejTFwoYr
svRp+IR52E0RYELHAoTQp0XcwNgxEDVKib3u6fgpv6PTsyx8CZFizdYMDMP2
Y/09xRapEswWdqFyIIzh+JTM1HXyvHh/mSvzSTMGI2rZLsf7TyCanAKzE2lj
T31BO3cBXWp+TuGqXmVX+WN95juszj1COFg1w8PWs0hmUw2Py/K3wDKyfWfS
TfClZauOiH1X+3lH2TVzr9bajCuz402xW8bznHeIP0y1b5MxapTtV05gaPdG
1btUiPmwWZnRFatWQiabDOfzKgClytWiXpufmsSSBPymQ2CmRRpf4Gey1w7n
5A+ubhW7EXMVFBfanOiEGhWEzetP3fe857meGxpAi4XAlbg5CHkM14zbSsmD
ya9vwDpwHA8zvaloEEpW1XMXLk98i7mqWp2xfAs1k8PV2k15P93KkO+1Sz9Q
xLSov9GhsAEzwUEaRtbALjUU2cHOmunmL88eirQ+ShdYZnhi1B9t/4L/GnAA
p1hdTK7dThyNlu9//ZWclDEGAvoronRzJ0vOxxZDP95IxF+iMabzpS1BA5YR
Inr7vFnckwoxftzNJmPPOSUp49vkxNC1ql3fqk2eN4bed411YF9IO+UV+o1P
JNRu6iha3WwrdF26bHiLzItQX74g8SnjXjFroxHlegkcU/gHRLAdDL8niDc0
C6Js/gn/oFp4CIUqPpTTe7a0FGVxviIAVkRw5R0WnJzsNqW/GbsWzx788qTo
u9t8j3tBtXn28pMK8OFFC/01VEg1jpVNDA0sTmCl4RImy55DUrnQWoCMNIIc
ERrR1Jvs00DkqhKpPgefIQ/WBX3Zr/wdKHnmTbKC+rj01Ca3tsb8ocWzHG97
dqTaOePmnpd3lGF6hQpoF5z8uYBeZT3lOBbuBhO+BWvB36HNIfrGTvhMsqPK
XesT+Baggy0wSFMoePnnOjDzaaHi4rgOvIo/bhevYWDuXFc6hcyyFqXH/3kq
ULTqUnvSdHjzHDgtJnW67uz8VdSC9aonJYj4GDzxP08qAAQkbWs62N18FVAL
dyfjhep78LC/nnCM9n2knC6Ohun0a21H0xWF6O56alUIYxOfW05/cOLY6NjU
HQ2BVEsFqVaTntEyvLcgUU+zezvPJ4SZMZTCg9Utk62assmg+fK/IdtlhxL3
2flh/JE6L7pqAhnRqiJ6CB56GjS5HTYeNE/CP5OnwAyvRByEIf/BTZwJkWOx
BGhO4sFgjPfoC6nBtAC35ZhiLRgfDJTBcTqupyueGpxmMypR3Y8pFOAs044g
NkzBWt/5Zg+G8q+8nxHmFUt4XKbCzXhOltqlCMg2jKScpMcjuRdiU56anJAU
qUhzJutOPx0Q0pgDasr7q9hNkiIePiKG7oPpQC7hgIImH+VFBjrUOO1XNS/Q
IhkATFoGvZI3fZD+X7rsql9E7hk83sL7w+q4AiXey/Hgzr6JNgKxPFs4aVbL
2QwTq/FkHql7fZ/Kmmc5RyJMbMmCwga41UTBKNYMeq+5rRicSI57pg213C00
oKUZEHSEUPWOzYjzx5zbJlBm6wAAUGkCNHkz/pefepBYDUL25s4Fhs9bnrFZ
m4MUVoxxELKTI5oKG5tUfvPi1wvkYFTC658ckqvaGDcsy9DA5rDLXm0FDSOf
4Uvb6y8qiVTp3mQ9MkCfnvRQrtplSGr/bSmFqTkcmQWb8tRICwr46meWqN5r
bnSM8eMJMXbYi77prIAlC9T1QCbW2wWFZWH6U1iMdfM+5YCSd63vkudtMvPk
DYhOxwOcS2sImN1Xbjk4qjmKwEP9RYS+RGDjTKehRUVuGCn6bomKBQbAbFKh
3W+lz3RMRm7VgkU8bd/uskj2gfLTiHqVu2Yf2rfFtbB7Luae2Hsf8nd8lxV1
21IJ/1zUol18r5hOzs9TFLOsnOIw7qeSnPznxeEqoMP70+/2qhOWTIVp0p3L
XciRjFwRbUty4RJIStZoMIIXM0dW1AlIV3A8uv/qdYJqpmCqlT5E/58lKhLq
PBb681ClW7P2oiZB31VKd8J98KXvj7WJbNiQqLEmbo5Ph+ZGiuMHyY3k2L/r
EfsQ4MPJkp2ygueaatJWpm20XSYPGJrTyt0R3mPpSaK2gPztwSbo1KreaEtB
pOsP7uRLne6q+bAYarL7pZiTQSoAmgrSz0gLjAscByz3bvGUxJG2eg538LCu
4F1swHy58N1nYq7di2oOUFYF2yJBNp3ZPR5oxPDTrK2JTV7ZQ3uCgrzHFtFI
oGZzl6jSKFAPW7UkGw89fK5UKhmn62LBVNAGltCfdeoqOgmIinmHELgTboaN
BXBsxeJjGKAxwaMeRxxOJhhhnDCfaqUo0Y+xyXOb12jwzNAQV33deV7bh4Do
VkkGr/GfL412Ze+1MP8EE7yYOotenPx5L8ybC8QPq6qKSZnQLaOhclbC0F5N
xyHSp9Xxd5FW9IpmMkFl9ws9LIo8PlvxAflagnEYcMrhWo/LipINXieSFlbB
5512eKMpLrnirmG1RhP5dqBNtBiBfajQD5QZynDolySl5NWasZpXhsc/UQbe
kIsoGfdrzSR8nQi8qM46dZ13Aa6l+2I3kuF8wdSDJt0aNvqb99fSKX9PqNJ2
3PlJ4ACXE1QswlZINURixSZ8f6vuqaIxTDzie7/HlkGKdQf+qdN+828D+Y79
DAmrQU2RzM6fj6Kf2a+K0h0vBdRfp4w3ceLmWaKaA9NZwVuxezpFxUnQE+t1
9dsiZucti/Nv7KADBWI0l5P9Z6FLvPk7BLwYD+i3dCwnAAbvhA8rrxGlQO9X
vNM8ROMAGa3uRB7cdt5St2Hopim3FBurhM+u10OKoArEdUhJJ/AX02IHJMBB
2Wt+ybgtpMjiJ64GxsLaMU8YDwBESS9tVTM2u5Hyiywp3RckufVbOM0cWIqe
AKCYVqBbAqe5q9jQQkR4/hFj4hmRpVU2y/hdzMYkALsWdXacB0vZfU/uwazN
zQDP5aPCpXFRnXUZ6vrPmeTR0iisXwpWyprK3Na6pGEYD+WdE8KNPzUtvb0R
dk8gb8uZ9HbYxee+iplYvbBbmx2pfMzZk6BH0DtWvdjxL4ovKH2m8MkCyTpU
PvgvDeuSOhLetTaE7NeW1ux3FtzNHx5in7hfvEKQXX1YJ+b5m+WS6EiIe/i+
PQQfaT7b5e23rP0YDE6V78Sikb6syEC4rexxeREpdIf685h95RVtI8wg7ICB
+8B0YVcTwuwsT2uNHmy7vUdgl6ncSEtSFi+UOVF5obP8OSD1bD3Z/OffNNOl
gFMaOPOxH8oV/zgxhdMRKUaDYpS9NVCfmDyofVkuW/wRNZe07h6VEd3VBEVx
/K0TqbkexsR14yooqD929TBRO7FVdCfV9Qx9FXxrR5TDp8Mpj551GQcdyMoZ
nL5dzqSuliakH0/ZblNOTmJ9btOtdhM1gn5AIB7OFQO83Tf0hej0Pyisj8rl
AcJ1BgaVJdmRDhE/QbpqdtfhOsWeoMNX6xWTDQvcvVOfv1+WF5a999SjAUSy
MARURFTVWLmLHXy8lRNb0NnquaiWZGaynoORswbuXvZC00hCQN5V4CdDtUwe
O49uL/gcAQNIuuH0q7K1UXFUZuQzaXHnyoP7ZjMxTtwlH/oCon3BCg+IpV9J
HK7g//j+JAg0vb516zlIemmtfK9qFyAOrzWTCRc+3vhRWh8slCVCOCzMIGHO
ejrPcL/i8tjpWVDwxVSDfaDc2GpkSBec5YB3BcgYWtVTAU4QpOvGZGYqkXrU
Mjlqpy6BK87tqCrYY6TvCBYc/tmjBVuUF92my7h6CJ6V9BDxHOfTLSYyw78q
1BZXH4OvAiqyKH24Eo1hEszUDuPva8RoxLbzeVXQSJEacRvsjSyh+m7cH58t
BG4E46nrSUZeyypnLCuXeqMWydCaoIdB58E5Q8+4yDrt4zUFJfRaovUNQ4PT
HTPFK82TVDrCIshn7tOpw/J7goqPw434IN9Bs/QFL1bHFwk2jIVjedJ1O5eZ
+sfRwxSQn15bQZyXuz85Tvh/6QyKTlHjyUJp41VRWWSEyH8JEPJMlkyg6pM8
WJYYjT/xPXuVQH5IdJYOUk4Z9Gdm1aOZRBRAEXW5oQ2rK+iZ1uu1h8YubZOG
6WVNcbO5xnxE+cfVqKV+5zis/GoL4CJtRQf7/yjj3eDXqB+YVJTkE4UcbzbK
iaRThaOkox2U9SpcivTCXBXXQo+RtjSJNZb5UO/FGCQRym594rubBrJdMiGN
Dk8zH+IX6JI7B7GyMp5uQneLTQZF0t2r4lHlg0sxnKPHoh430vQ9y19oiJbG
bqsRc81EJKMOKCEnAzHG0VJ57h4FEzTNbt3sBD0xKhNIujKL+WAB0S61Yt1B
PWCogRpV2b6l6s8ItHPWLji4LPdbRO8Jl9/+jCoqUyt6bcI27pNAqQNi57Jq
QVnLq8aPJ7A5mUEX/kQ6Y49kH0vHdAJi16GKbNuVURHOHnrRe25QEHEA1OD5
kSFYjzIBbmfIe0vdX2W7HdkNHO2+ROsA/5xr9MxTUfiBIz6TRee3A/rqsQ+f
iXDCgqs7QxTI+QmSJdrjA2gXUNIDiRVvIT9YuzYSm46fRl1eIzVyqLdCUdXX
Ie6WArwOenVrdgXsN8iCOFrntS18Y4miuAV6ytbUM42ICf4mVtAHW7+7P+Y4
cXaNeK5uMwX94gGGeFQblOdMysMyydaZu5ihYvThwXddYAhDv4CMbJTWnGWb
HiTMHxVjj+Zs6UYXoZSJq5ed8H3zBJdj66Kq3IGuLRKYXzcnF5ksnQb6ZlZG
PeGKmcr/EKRuPH6S3ZcJug83o2yKdjC3a0/h/yiMn18A8/hgFTUTab5SZBQs
BX1S3ByHGoKJQf6R5CBQObBIrZ8ZwmkOlSdSh+o/CPTWY7L7yeOa72Vg6d0f
3YdSbi2AA80hTO0tlMjxZt9+axzwt5Owh7jsWs2nP7i7cpp9syjmGWyDb+yI
n+zBluBbcXlKsdt8Kk6L7Wc34fEwwshsWYSvbOON7UCOIkLG7BeBX6tdv1J4
nhK8s0CftS4rwIwpsprAJn7hLYvFCnvCZhOTlrv1983fiSWM4K8366nTpQ7o
wvByTGZpYhvRddMxSxwSTUPqsXalehuOnAN4L9S5h787o4iK8nFmlXfpDtr5
OSVWiB+ktQquiqnQ6idyDG8adm22H9tmYdZY4jiRTFVBMNrmMWt3caYsIiJs
qKAGNDHheGOSsIY0+lPWJnpPzrJhFLac4JIH6E3ezUHVavSyXGBDHQp7ry+N
xNPupcwgGkpQa1b7sIRTyRF4eYaqymBHEoxFzg8jJwQB2W93NCN297H8JlnY
eK2UP6b8JKFpmOLFPOyG7UY94m1jyBXwrqAAJc4SVIcSjTuuk6D6P3rZCJCb
Re16HZ4GoQEt8UfN2N58wN4jXIS2g9C9u9pGtOMzj/QnIcn+ZwLDDEQGtvU4
PJZS0Mvn9qWBO/8ggM4ZQhwPRs5zVAcb2DH4ol5G+LXNmmhB25/VDCpLMNBZ
tDDZhya8RN9o5t6cF3dO5q3ytaVdSOkkEp6eXI2AGrV6TLnV3IIGrt+0hRJo
DV+OaN0BWPPDpTU17uRa20Vkmm33Oj5hgQkgOZsLjqZOEu5IUJU0EyPUyhO+
TH0PKqXbD6WxLLFWF3FlZHAynnxkNiyrSg4zfbJrPk6DhC9y+bS57CmpJuar
eXdwlVvv2EGN7lkn1SfNkKWuaMkyQ3aLnWIu6L9MLwhSFr3uaeses/mYE89O
n6pr6sbOAnQeNc3gcPvwKebL7mMGrCtxviwBvj6ot3AWc9uPAXo3Z3HjngSp
awP8LyzTebWD4uBv/ZQlCEFPOtITGqmwHu6q0O9bxwNeHDPJQPOR6BEWPlKh
jETwF4nrsKnL7YulDpLxuq/cZ1iJZ8FBNRJs2sbFmEf3S5xbwmFS8TfdBbJU
mNaubxmdn/+eCloNFp1J6oZUoMJKXMsRqDmMMftDt8GNaLPSoNT1DNVKdsjb
x/7WXaQkoDmAYt94PRakqs4RrM/CKrebKzuKYQYyaXK8Woe45TQ0G0aNG6l5
2G7PgSOUGftLRtKq7d/Vfzio9dqbek7f3gZJPpi/zyRr1zSCLthiWIzCRpuk
7nQm8RYegDqLjDA26vBV4vg8z52QPiJojkYYNO0M84qyUiclAKv8T/nwtBrw
wftCdQFtx+DkSBnQTlLL3mnfZ/HU0oFA7O7UNoe9qZQO0TEb5Vrv+UHxJ5QX
tdGaeYCCmH/CualYGmXRgmzUlVUBGiPmFV54621hkjfCoyX84Iv1oZBxU9E8
uk2VLx9JiYBDbUxQgZGiXjV31WWVwDc+EirX2cmbuhFkFaLqkYc59lTM7ZB5
DxgqDoAuErj9QT9NL2Quroug+zMWcodu6JEH0WoGEXQWhXawcwTdfHpqRW3p
W9N69cfevJ3ip6gJA6MElRx41NTMcNw7CUex9ZDyr85XA0HqC5vKDjanQeKC
V91FqairCMuv0Q+nOCgwvMFaqcMrS6gkEyjPvh/hv9P6mY2Zf2SZLPsZj/6R
pAK5Jv1PhlZb/YXXZr8x01uLIxavQkm8aerRu5Zf4mfx8mwI7V4FTxnWcJ7V
vvhM0N/YCXHmx/YGQTR/NFdpQooUjTBACSJzwp+k0SfXQXWJZTQmoxxbiyEa
NMfH0XabFy43NSRXqqFN0tna78gIWOChMaDTIgUDdlSuEEjMumpaTsWWVvUm
xLYiJsJODPetitlBrFgy5lUdgxa/KSw8G3fGbFK+iGaY6bPDsStC16dsQ5by
h0arvlfbibbYXE3IAaCoVw6AahFqaaC/qeuyFhGoiCieLhdioKJ47jZKBwGb
lIEZusaqWj5lA9e/KlHzmIlqCecbVlmm9xqrALbNL7Qg5K3num9dp/Fh+vBX
ou2/xfRGEZ2UM4gcXdrLZ1tx0Gtm/l76iNtbBRIJ6aMjngHhGqdYYh+0ehfw
sdogECuCHLAWVK75dQa+k4koDlSDxYjjal51v7L0zJus/GsPsLNVmQaWzT9s
ocWgfMnpgY6Ht0tytd0IMXPXC3/T2c8ErVZtgv+3moop2oGFP52hFYgnyAL0
ya1yA5iruR2NZGNelzcldCgNDGP4YKIy+4g+88lAGwpqWfsHWprMqCauwWOQ
wRy3NnW/inB1sKuYAELR4U1b/olwJiZtJ47BaGEBcPmtr1PxUrNFk9yTiwpZ
FSCIYqstqWZ5XLzIxxitcZEC94yBbmwKq2++l+bji42HcxTq2gaJWc3wGZnh
EnGI3yk8GxifU/wtg3/V/hBQzjFDnFpo4CC8q9Fp9TDuUHB3rx7FR+hjg3K8
VuRZVmUA3rJ52ucpaM4bS+HPvyXKvXxMHghOmLPL0lUZmYmxgDPxGxkbChOo
CwewgIZF7j6R4m7kkbEOpDM/m7e3DPfz4IliFy5A/PRC+Yztt1xJcB6hoJvp
yS+UTlP2T8+Dk4Tl+keMSEm74LbJhOJuGX9MuNR9gccYMFtO1MFPruaGFvyO
GfwsN8+zct4DmDpzqwZJx/tl+BhFOV4qrbNfm78tpdA026s1xbdx3xkSH4fz
dMa1I+xJxtoJw2mSBLkVax+lvxRhjf72dEZHf5gkKGtoSdeiFwWmc+SBqInS
VtJk89nQobQeFGahwgGGv2RFf5qlkubV1MASR1vS2YGYmYC42WfNqQiNqSL/
4n38kd2aSiRNFwcdbMDwQWTMxMA5unHHuL7ka6SuDcpW0lDI8fhzOG0d1rGb
hBnNW5uAMQEiSJ8j7rRXPFDvuflilYzZw1ac/EYKhky7P7/HCHJLqzEdgLic
/xTWPRbSUrkGDkxRtIbN1ycS4KKQ3T8splwL27us+SnfDVgO3MyhOUXdBWJO
B0VjjHJTVdaL4qzWn/gv+YOC/yuqZjrD7Wi4LNCZK/yhxBoua2/CJOJcTv3S
mJYzJmoq5SM/bduSkEbYB4e0W81+Y+s4THTgzCZqY7zzCHwOv+mn1VSw4R5e
Fwq9wso/64trr1eikIebsqMPsHV+w/nIdkPrzp6TtBefb9wXqA6OmofKHvUa
0Yp5/FUhisoJKw2TdR4cZ+aAQfUUo6C622KvGKONW3jX+EiaQ5aQcjnPL8Fn
k76d9O8YGwENDUtC4R3vQ0g+fW3Qc3tCvUSm+ubW8HzlKAJ6q3DkvKWSpGG6
BoDdmWyLwdtPbyOE0M50NoRu2Y7lcW9Ih37fMBr8qPexWOBCrQVtrFI2rdz9
n5blAn+0dRUvT04JZSLWQ0u5fIUQvKovJoer7igipxnPZ/4n1MoFEUQ60Fm2
HhrXy1jaBTcJbxOhoHlhVy3x5Rc3QxTD/gAsmnpY2wjPWqLtZuZufgbJdMgw
MHO7aj5Y/3qVCdYweSqJmftCmh2gbTV9yAEoj8Tw6GHpIg9FxzPostQji23D
IMEff7k7FOXDlGZBsODpzEDxnFDefeN4rIBdbnmvinDoFTA8daIyHvYciB3E
ayzmpw/7jOY1b9vwhz8WRyrgTWqQz39vK+SVhIcjADRRT64LBi8T4qbK8xHM
97x/d1YlIJSQcSa/qHZm/tYGA56+l5Bx2MvZMo2w9xZhgGO98n7zkGPxuPj5
5/F4VTNLbz5fL37l+6xuZupV/+xBqFVcDtYbLFs20eRUrKxYS9bN7dyxCc6N
Yxl2RC2G8eHVi6HrwcZLGsTo1akAJCUWvZZjhOBunGHQaf9HcIvJIDpCr+nP
9X4EU6YmtoFSWFko9eSVhTDXRBPpeFezCrc97TNzhpBm6EBdIHH72TeH0c7k
+5+qFJp5U1xE6imh3oegojmPjHym75Ed7bqrfSz+V5TP0BQQtkx25RUtUNx5
tLbaxtf0v3gNbBgGQTBrknkh7P/j4zhEI2Y7zS/AmeKP0tt7gnx6BQQQIeER
MJ/YhkH/a/EZiqeA1E47N89Gi/3tqb+b3je4ZiGYfuTmWkgiEl++gukzbefw
MBqv5x5drQQERmbJO5YTt9oozOLQKT+V8IJ/juMzfQjPHfVCNVD+nId2U28r
oW2X2IsO99s+ymT6YJoUl+phVzCknYKG1E3pzYL26QfmujrQgCQlSHdH3exc
chA81NV2+s0F2r/etQKQ2Q70iA6elHsMTbizaJDyL8evV74gn3ddy8U18rOd
oZSFt2TWgflJlUH+2+b/rliIRXLSAJTxrjfPa1IKNQfUm1lUkK86MOuMOXQF
ZWPw6CgDXz5Bnz1TBSUkPC0aioyvvBGMa2Xywx3GFtXvDD2D4Lyt9YBXRFoa
d9V1zwzC76UArww0UC3s1lPYUwKabh2YjBEbIeY8TMyVZvspkfez4DFRANFC
Os7QFSEz1sCAuLOFhSRGQpgyQ9vICavjmL14NpxeNxe4DazUncGKnskJ7N9N
YMNAqK11xN/8H/EoZvBUpaSSPrYDmGnO5TBkcbnjakoXyKJtsRtm2zCgzOLZ
na868BSFma1dB1pvSUehfoCJM/aKH8R4LIr7ks9r+xTMHQZ9RPIu1mDzZIvp
Yn/Kt1Pm7QTBf+T5jioSVYpCgbO7fNX0sAf8gqNetIaZ9K/G8wd60AzBLz5G
fDoGvzzgteNThm+kZOLX6wSOuQqll+eO+ZogqukRhGJ4+O6u7CTz/y25L3QO
BGdxaxCSICvjRG8M7UVJafiMpcCyPhrW0Zod1k9ub//aCD/aSbCgpExpmFx6
8TGht/xhCLOYlH0qN5zXv8mtJ7QV4HRgu05pGo0ZNXG0vXAFwjfX2WYdGlzj
owM25zXvzOe2E3RF3oKdtLcb3HZ0DiUpvsKwxBPVeiga+4KtmipZ/9kCTohN
ty4sNPGcgNPbE/XlBMb7S3TG/lcZQBjKG3GkZNm1Fvao2SDWqfoKGaa4EZnx
7ToDJDUyUDcHT1QaAu+X0VD5UQ5pKGUfnd680rtLi/om7pm3fYxCP6/xWThv
xUp78mnbzMawmZhYrrnL+2RtcHAKXdKlWNhYrvpOjo2bi+lh2X+NyuK5aBGQ
MEXaw+h2dvFCxptHQFVQ3G2m7P2H4/zDdkxC/clP6pydL/RPx70vwyAEzbAY
CjTHWzSn+x8XxQpcVNrfFB1NvoZV8LZWKVjlYqtDjXKTcU8JK3eaafYRlTyF
oZynRv+fHT2VDzm0oPo2y0Xv5NPNXdCjjAd4JYves6tPc8b+5AhCR5jel1zz
sRLVB3lmvnFe2cisPOWjczgoW8u+ctDXEMwla7KQxhOgVM0Tfp3GiVqjLvSB
6N55PWvQBhCmpKpnWDEKZKIL2ZfvE78FISofn+BMq494tLiivAyn4HJLu/2V
UxoyN+Uumkx1x/OeWTqDoqEm0l4A9kQZImuL9z+Bxfnea8L/60i9SpPN/5ju
prOvL5rqSQUMyxUCCFoMjZqe/gouolvvIkIvfTX7/MK2Q9EEfglRGCJL/Bei
FkNc5/fk5khSoCcrX0xHQXvR9bKpogh6alXv4D8B91bxUWTBO49GU692IAuJ
FgGGzN7NA3OySxIKFVLWR/0c/PqbvNi5f8hCucmS22dL2EJrzO+2SqgoLGaE
6OTvC5ZAAfpHvq9RRCToEnDBlnrZDs2ZKfHrH0MPME0uIRickbQxxFsmqiJe
w0DoTBjIuJ8zZhJpnEH+ebo4cWFJk5FPYVWrV3npqZqJLdSClXTRjdJNQi3B
7rAeZHYKoP0vwDWuabJWsc+sxTpiLEBLDCq2+MZWEvxBq481OulXWwgOZQsm
e5zs7VQefCach0x624pth8/DGhQMO4fIRJ+75HOjwGhXGhjQq/2sLePvwRti
zlk7j06ebSDvIQf0uaXoi+8701jBSpb/8Tj6iOvrwzgFKQqNUhngX6H4iGbc
upqtJnHuiEX851rmxuATwkwo/S2No/UCyZKmKElFvqDgUKKtnEXEFlaYE2oS
rddlc5TDQ7k1FJHVdo5nXb/63ruIr0IzGYfyVMP75GWuFEG2ubX0oJvXWN1R
G0yjcwrpy8GXY3APLSgvhTmH/TEdnVga7yVKF373aeKdRP9OUpDX7xPsSWfR
+joqRxyyRZEt5NJ3GnoA+YG9BbBgv9A25+zru6kLGJkQWFtVvdWaJ1LGP0BM
anpmGRmlKrNeJUaxKKpXSsikahM5bWpMqYvvz56C6veBWsifFvKscCD6G2jg
+QHTCmPEOkOCxtms2WgRbJBTXbeNJN4hH2l4LCl53vKx3xMsrKte2EybbI91
3wiVLUI+Zm6QJKIJER8WvUILeg0gI9n6CYESwajsAvw2LO3TjJwIcgSy+G6+
QFBoQluacs5TP0YSs7u1QTicLEGC3AXXGeGLj6yMFYmtxT3ujmBVPYKkqBtT
67s2YR4QpMUOtV9FeP2S/AFhLZFA+leS977ro7hpUltzR8JaKh7X31GHeDQC
pL2ohuq1jRMFiSQwpN5+plOiBoeh4qPG1NPJy1VgJANc2f0v6T3mQbWPfRtB
UhkPxHdPI+43DYBZT2aAxAc28yX+h0nYfe4Xs01QpbMgcjaU2krvkd6C5X0I
O8L3KYTO1mYYXXiPjknFQ+DAw3TJOngUKoBRAf0W1BM0e7m1epfXwjFyxvvq
He3VybKLr/S72KwGdCvEitHO0N9sHFAemNr0ZUzGqDU0f1mQ29Og8wTyPL4y
gfAqTHM8F53N3luTNYLiEw4iLeuYSQ3M9ZZyjFFu4OxP2WMELAdFC+Xx5qzK
m6XBdQ8rUr2DbrHXp6r6bn0IbuRC8zIGCrRxHLB+poYup8tLv5NyDlIEzrJC
a6JOF4N0izYej78HN5+nEWJZxiQV/lp/hV4mh3H0g/+9AljoxkW2mg2LWeja
TrmHAp7XbP8Rt1sC7kczYDct0FzsQZle+1crNIVfQsEqDmQXaiNbFC0bxL3d
lvlx8vmdwpMwZBb+60Q5xV9Z3oagzVmlB2POZzIGpMNn8UJxZp5gZpaUtF7R
BzHhuF3rdzdE5YK+PAHA2bAy6pIvoxd8XKT4SHndTTGVElZvkaFncv6Cu4MU
HlppCOHZeeABrBl7qhMem53sNoVH6nVyLe2GFmtuOAV2orDSjcSiTEfihQsJ
dsO7jo+W4tA39PSwKDYl+j20UVmtt7Tb9RgF6OuPHe60Ksg7vGR5RiTLFRCX
Wr5otZiaUJrVx5Af65raa7ZTGqm7d2VNST8AQLr66f9Eo27tmv3zafmIahR9
viMg9EpbLqVfdyQeFzntiU38+qC7OVedcHFdEnDKtMF4Ji/OWxRM+fxZq02W
M8QCW2+Xlhwmm2zjxv1uMh0fAev6IdLpycCkYlmb/XkQpHehip5lDalr3vWA
MYHyWz76R1Q1yRMz/ckkKQuPwcKvpmuglFFK8d44s61Feqe2YVxWHfAgMetM
aC+a8RPkZm0CeRAFyvQZwgG/8pnEU47wZZmxxb9+m4mdvglo47DMrMBiSYtE
QeeqoWzE11lsq0Kf9J/A6WwSWXg3LyjuTkhgwnnmvtVVgnfD6CLiAJB9CfRK
db7ucm2GzJbeJlTbHYV49S40spC/de/7R3rVKkYcYnfL+c9omCjVozs8N801
hzWxzh29xrdhiTj5lQxDtXFXHYxE22+5XiC915k2MKGiewDMQw4HFqrk8iq2
vmAb+2Kgk+7Tn09vVKeoh0KZb9O2zyKIu7prtmw/j5mWgvkKUDO/OB5uUjpf
NV21r1M+wkBlRxbzewnsNDmJxOffsw38YWVDode80H5JRFkmD634yoZ7XiiO
gcTHdODjx5SHv9GUQqxj1bpLyIztTaQl9q1sljk56PjxmWgE6jKENzkLk2JY
zxxlvQ6SQrkZR7QqN6yvPzdqBHhdIdqDFKyRcxhF4VgEH1sEooOVVkjDFAql
PJ4qhp58ZZ+y8oAyxoAxyTcWwaPDSOIH8r4ZW7XN77glurGO45dzDlgKar4i
Oy5XVd530QATai9Bn0vzYn+Wv/revIWLE4yKKeQKkNmvIzRZ9AnTaPlwZHH8
o5miu4xoj6tGl02DVTcjZYosEz7TjQNau6uK16gg5I+Lt1C0hmBzy+Slas/l
TbDm6P3Qj6qvPcc3VLVFQWsokSJphbgXw2YCPqlCJggfn1kGmBmRPWdxcmn1
Tg8BSnfrXS9+q7jzfRUkjBkwHggandloQjhA2CvjyDDsOjo+59CCVTktLJqr
QdWwWZCgEU5Gja0lpemrhh7vRnGmS9Q45hwAew5LKlS3q8kMa59xk58e+WuH
cwk14aCPwxDgiAepF1lF3zby1Zh4FsLL2HCxnAMSU2ZisJUPqgTgeocIpbfu
5VeZRftG0h6cLaSZiwmaJZ/M+t2Sh84C7oEki3xxlaoZXsTSDdjQYIjrJk1f
rsqTatDkmG+TRY+aai5ajFmjaobQNqfDOZcCEWFvKkZ5bJsG3qrZFO0ohJGH
UxWx3tWwqvclGbFRMKTF+XOKGfnMLtNxwOSK0f6e2lC7dG/l5rJwwbKb8x3H
jHqz/Fx507MH7x67MMDBHZ4lOTvvxxl3QmM3gxAPnFbX+2L1PBMMiAdOfmqv
CFiLUf5DyFw4ufOT5FNFLqiRhYFjU8oMLUbXjm8pUEe1O7dSfz5bzWyEw399
WZus0IeIpUvodTGLRq7zONj5JErUrmkBl7RgnK+MSz/fmwBatBgnOURnGftB
J9Vek6W5Hxn9EXyGRqph9R5A14ZzZ7UPcrPba4X8oBTGTCqVWwi8dPTdjHzP
UfZQYBPsHnJDYAbCbLgNo4kWTie1Jc5pG6uKExT3uZi2hkd5VThAiGCvTM8k
4IThFpwODrB0dZ20nJse6xRW66IQymYyvMbl8DqqPT3R1V5kDyA0qjxV0WUu
oJ5fgAZABOj4wcltNxz3TG/9Pgco6fPtxgVuZLNcqDX/Oq/6TRNqO2By8Hph
6CPY292918Y8ziohSUdU1DgnaQ1I2IvS5+zaFXzSwqPwn5zhv2aypHHn45T/
/sS6NTYKfGJUz7pKvAYp5n33NkSV0gujw8OwbvDpJb8/wz4OQdivdabZUj4S
HkTbAX3cxbJ3witOMRSw2cH+fgKMbV2FxVJNxxTONHDpzwx1u5GUUhN4kOmg
4V9v5xWC3hfBvgA4v7qeYXlCIC/mrMr8Mhw6FTCRtGnD8myA0iy5EvYnNXK0
4xVTv+uBgm/yg1Vf80smwetma/1fe4ek40R4pKhgsAsK+K2+8Xtt435AaW2P
ffD2sw1nvb6jmpu2I16yxygjn8UFidN0GxtrJVWaRP0xo39aqJXEo5dNY5qF
kXOj+9FFZXzZnyZiwbb+opJKPStwnPTNJvAUvjCy+XWGBxn4K9qt/RA6FIuy
6I8sN2zJoWrwKrrTb7C4CkirOgnEmYoV/GH4jEUwYEDoKM821c0M57tYFw2k
n+CqNcrxZr6hGNpk49a2yzFrMaKX67yDi2QX8f+rEENBL6xKvvwTzmIcEUNb
rZrLJAaf3LJfuz2gx/SyNLT2AKg4haP0xYQGOlx50K04B3obojJHgJjkmah0
oqNBAh55a7x+65oDgj32kVEw8bllg2MADeMTBPJ2yskJUW4mgv0Thut6y1gL
nlVvPQ1AWSuV/ARzuL+o9RVpKNRfxGvI5qtFST10C53NJvwmrTZFw9j6s460
3UwR5+d+fv4ICYmBRNqj3JthQO/v26EIBk2JJc04dxpH7ceGyZ0YGHjwLYjZ
dUdHYSMNhOsfvYJVXEyD/SHsW06BlytMvdTfSA6tJzPHVECG4GAKgU3gzVkT
g4n2bX39n6+qAPsD+k8qepRbTKHEUxnkW2ExTD9iGzfBcUaLqCXH8rQFvXPz
lvMYxjqIyglKa0wj/xmfDlMq+wIyDmDGJELRc5bVO1C1kMoEsEzeKOoZyGxt
1UhW4STofu6O8YHtZVjzSemJiyYideFulQshQ44Mb48vqoIxozeuF1e+3ebo
M6dJCzfuTt1wzp6mhYH1rgylxutK6gQigje+hIOz4mHa/f6aMwwmIXrfybNf
UJvSohCLv/3OIzkpr1JHhGsYhYWDhVlaBgozEh58UdtrhkEWAiap4DJanoRK
C7VjcMORPS93YwOLE76RZmlG6dwoCUVrkunzHJlgJBMg1pLJtiY6itX+8fzJ
XYoPdzHA5uSHm56hpBcJUvTEalWFZnaPzW4L3c1tfXVdmyeQ5uHlTMYjAzGn
2qjjOpiLRhHnejKvlWXCfd1bqMKp2FmMNkIDymYhUKcGDd5pxJtwSGgrfTO0
Mv/NWmwbalzOF1yzZtdkysMMzXSdD6kqe2f+RNOcYwVg9H5u+2Eb25fiCuzS
hRtINX+pSmVIlGU51L348RngjIjkQ0gxsmFnhJw+K6Yd1sGWuAagz9VhLB+M
tCXmvj0uLyfQ8QR9dPanUxWaTcB4bxJeeN+JDzrhiIVuKs6wQtClOx8CATCK
xwkxcWY4LzcPUt65qyUPAiUBJQ7/jGCWERItjJNtgWB/wFVqSem7vQAvIjCD
wTjBRpSqOQJro/UP0p3Y66TXnmzwYtnPZxY4RSIvEfczIZHtwkISr8TLK8+M
OANmx0jx7e2rTGd4yllpa0ECfxdmTsifBwZ2M8f90yA1dCABsgHiR9z6L2g5
3bmY7hu1ApIRpTQzYY9JSPNc5gRldK3wULQZ86DU0f/KvT8XJe+SgWBJS1/b
ieMRWxhgXkvR5HQP2o+sDbL/x5ceOAJ38uBFQeB1hLp0gxYHTqwDdObK6PiQ
95+GFBClSwxTXWWWCCB6C1cxAYpOdjF8czlVL9lxB5LBLMzt0lRAwSEATTwr
5oiUtH/DkQMQpj7TKqFIiutLz2+22V+ZXxQDP/omtLTwU4ia0ShFk/IUPa1G
gU+9pUlrY7fbNU8Ci/QS9ATBo1W7JtozOEx5Ryj82Zt5SwAx4EsZzNAz7qs8
vwPfn3vlfVvi6YWkwZkP+UmLgNVF2V0w3n/z379b6qQ6PgDc+HbiX3S5E9zB
o5mmw3GYo/7YsN8JGtk2ZdfR8pGTUbnu4K58vq5ntMaZOT9OtjlHjT0/YUEe
4V489vQs/+MwF8uyHQBImu+Mauu9x82fDkOIyggTTcHzbKT2AuVMHXJYDsKT
lYFecS89CdyOpb9aNWzwmqHWjg/jnLnL3c0rmhtRE6W7OjIVOrYSKC6N8c//
Acl3/eIsgNbjK4oGgqrPXchOFCPdPriJ1sOi/FkdApCweB3gfNaPAtTWVkhJ
QGDzQg+OoXbo+bh38rFD9w9UfBh0jerzf2e2iaNGWEy0zxOvWYZ4SCtgV4IC
TNzoA/St7aQJfvViTJ1+Lr4Qr+x+TE9zp6o1ouv3Rf+DcDoAFP2F3G+duqes
2ndYfxAOaG5FVtjt/VcRYcBlHjz3cAZI2P+VxEfxRbk2CKR/jtsL7ninZcjJ
oZWFyieIoFeWHSoh8osQnXETGBBqNQlzoGoR8rVQGzUAymMqRVG7INDe0D3B
z+4NoBQBrfihyjT58hcrVkfpFt48/8nu30IZdDFsQc0shJRXz3CHx2AXxzNe
xx4NJR5tYjp+qhHFtRLMmWJGHJ9WA4n6UXlDqQ3EodZbwg2bG4la9I8IKBIf
WZvohUp1mCjFoUU2Lyl0aY3zmESpROMbC7TddHslqUc8Je5QadH8SW3/Djw6
xX5p2zYOZseBRJTDjUHnYa1vGPQZz3+VLbJV0wb59Biiq+bdmEHzL5HW+4Vg
CHyHIDQ29WbbEvrUQl/3ncswA9Zugx2DF+aV0vzqtIa7dIvhiPUzS20Szm4A
d8Bv2+6sjXYA0UkVSDN/Eq5sR8iRSjlAqNRsJx4yJ7hSxAuHbwHwtaO8w7iw
0LuhrlwAwRMYpvuuNPQiti1Q1sHZnRed0NV3rMeCVzoss5+IAjKSCAtpM8bj
Vf5mPi2S6eFRBERJYb6kCYA0EDKLDqA5thQTfYc5hlhrUU1hIHj0O//F0a8+
efJRcgnPLOUfHE/VcQ88z5BTDddO/DqeIee1stTa8kXLu9JtSxvbzDiWGBEE
8DoWhyf86DB9BExrQPK3A6cLoPEBk+ynG35lWa6QP38EWt+Jvl4jdaTXVgje
A3fu9HV99hRL0pXcH861LNYDY+qi4RTFxCFDG6GF8fHtiGfTfX/4odg7tpWP
1a6udVDtMpxRziolT8BFD1JVH9/7KNH0iypfvrJLnQiUlIM7bJnk8L5qD9qG
xbZgsiQKwTyQmJUoCPYTlq4TkdzMja4Qs+DbkBHPNHxoqxQ36rqvbYLhljxw
6mn/Dq5DJFZW+DjZKur8tHNjNVZTDe/8yMl1H5RTJJqowuSjc7p+M2+OqElr
9bmlcGIDhU6q8nqbD7n9MgkHXX6mW0CMK132CJAfLHV2VfB6rmiLgohgzmqB
/XtvDz5aEPp4EofWtOWmOdIEow63hlcJ6PyHzAenja8cBkQtFJlwFgDvjF9d
dhS8jm+Wgh/yg1ju04ZvEJzr1UB4nfSy7o6UEK/Hh8SKCgTiFqsAay923R+N
Y2uw+jE4iex3ZuTefZmmfoh+0IlOB1KgV+aYNBsd0u6o9QftkYYjVFTsLTBb
XyxjPCVaDqsh4iy9z2dsxPthbK9TWS2J/T+SAGaNV9c3dhGdD833oT3L2Ud9
RpKOYTPnMDn6GCkXl7RyRvWfKmYJU9YgFgzMveGW9Rn+XSAe0R5yOqLIW50Z
TVsKji+Vjntajxz0lHeshIv8E2g60xOCa4nIGdkY3ouqFGDVfS4GpTy46GPr
jlNQgbvg66zMZNOJHt4WR7Lgy8jaE1Ipjl+sk26vkkaYtksEl8Z9gMG0T5sq
un5jLsRwwy3zvJr7mkCYwmUtpl6CYa5QMdhCUL96X14mMDgC9xbnA/bTPa3V
gq2yqHC0E28J0VAlVC0YmLo9KFpRJYX27Zjsvwd7NkK+7XNkEr2LDZH763fI
rUriz6NiNuGuDSXZMxtcp8goMo6aGar4rd1MDYcSqKFPgUFun68Au4qv36ra
NudkoI7cftVWs8zHW8TtgLGQHMbbuBzsczikAC7m+W1S0SX7y1hBPYQaQQaV
bTTrkoTZJlPMb4V8HyY5LrYBqo3qKBPuYPz5ajUXD7YMw+TxNrF20a+J6bO3
ynRh7PF50YPz9t3Si1wj01xxfsULgRm0gvvcLLruXKYmGe+zGDKgN8edbuZT
p0f6ZhCpVfutOOJTvz8gyFXGZPG0Skh3GjpydjVZpIKBALmc3qCTTSkB1SxC
rsJ412RpMl0d95lF6fZvrO70HeBx7UNmBotRi7Vr9asp5YYhVlC8T6I9Ca1v
i5RmtIRr6BL46mVCRF9USrbQkF0pAA3SFYGRHEsYQP7iJvAPoSQakLCoL/Tu
fGaRjg34w6bRjLowH1lLUuLIK5j1m+M70fApFfO3UtDt/o23lK1gG+xcLwOq
Ol+4EaRRl0GClkzu0CE9lIi7WXXO4mxu1Xc9uVW0nZil3dnpNAYEfSdFzxgc
EO3TppLT3a4Kck/O9j3CEsx6XXSsSiXySJ1qwc/CEe897Lp7eJibGmsdHcf2
3Pk4YXvOyIJy1N3z3H8zz8O7uykkMc7Iy+6KHV/nwxJdLqbEEGP+REqbGCAk
swmSkPDxxbQ78xqeOp6z0nNByAe0UOdFDj/5bw8kzSMsEurjwjoDCFWtgbBv
zyS4BWyIZo8PscqesZGY59+2G0CZtUNQMNTR0+kqgq3lBGHA1cM+pC3skQqr
mlzaoyflWMegLdB8V9aToRQgiygq+m/NhtW/Pd5dCHWVptCF/udwfWs4gDVE
ibnOOFupJfDD29ILz46Ou8MGP0rmXN6lTfFOGSHQ5Ms3raPzAe67kOgA8TVL
SX965jl5sSHkKFyGnP2xfp5eEJkDL/Fw9jpNl/Me0MpRTe8TGGY7nGrkHAC8
f1Ti/Phuj7tbrUGjb+y58F6zERfaQiT2ny1+JEtSyd7R3nn0Mgcj9s9U3Qjk
JicV7P4zFa9+hfKb+vpbL8Lqo3jCp9NCY7ADRxxPlV4NCP0ayCJ8MDKxlfng
+PVMYVOd0/3crhXGOAxGsHFuX13cg+wfKytk2fJP7cTfRi4/m/H1FVMRBRKv
qhS1kjZ2c54RUsUo0FgvzGUyXgQkdzo+Yt+JzHT21cZt6H8qbrRzjU8k4UN+
eelK86ZGDVIyBySG0OgUPdMHw72RMgNbPTm0AgpADkVazmmjgnDyNkVpKgpt
ythD7pw+WrjR5EdXyjqcDSSyfnU9E+pk8AtSkBKJ0JdnV3bxiMwdl5NKGK9A
seaXgR6sOIK4WLDsIYVZ4SuBYnr/8AeVChxH94m0i+3NlZRdmrPiBGk0iIP6
nVVQC6rTWYi+YPA5H+mzSyu4nEqaqnndM8Bl1csnLWoslenjL15BRHXycGgK
/NmOqe+QqrKfYltwiHgR7X44A0m4p1ZvpleNQrB8IDmYuwScQog5VaaquhcY
fy0FM/cM5fG3xAMvY1IREbdL6RA2Xi6Au4UwEFdxzyoNHQSezqw2ktHtnxWj
xnOQsPACq+yLwXdIoclQjYIB7PA9Xma2v1/GoHW44CylCaECqAxSeYLSlZxz
d5eBd1HAiZxk3DTDTCizfeuPpI2aJJuKtnLzm+kQ6NLyWfkgKidEnzNnwMmF
nyLgnuTI9QREWhbgSpkYPP8+KPK9j18HbVqFt+zuYRtO9bVpSRqwWYqeRhJk
AELr6lkcDxPCOyf1YGK578IfGhccZ4sGQnL6n905FIJ+FNBD+U4urUQdTgIW
Z7MKG7Bd+re8/Vzv67LyEcptjXlYM20utNdr9viyrzS+3NWGcupoqwLxhdL7
gvj2i5GNncW79sPPyWJBoki7IcXAFtAviCPT+06ec4yqW8q5R1iduhvrtkNe
OdF4d0Qvih3WBbDbelcb5z5Y1Xe/ZfSGCszPEh5k4hq/VTzgkGJ9AtgvuHUN
J9X/Qd4zIU472h+Imy1VxqiP+o8z0WFyIHme7Fitn1TU+ynsG4ccq9xYXa4I
4pdGUUnIqoQSxDHMUwxW6vG8eCFgOtnjGKs7tbRuJ5UQzbgFnXCpsd+qvjlJ
294v4Fn0uTLOJdoNr25qoTjs+YME+0EvP1fX8kEc9r3/SG/XLCzj6YKFMQtf
pzDziT5O16LspfKJcmwW2ppb3oQT9mUah5y58HPvK75yRGfxwDJSOdOxtOF1
L+lCV61ua2licdM1944KI8hFQesSbqNTPvDRE4tDS9XqsvDWfonUKLJW04tE
GcpvWZFX7caT58CnP11/Ws1NRRsZxNUGDsgzXeiAVRRyONcSb7nzKOr5OHvS
ImiyY2Ftb2/fMBr7vRul1djuSrD/C7J6oQ4d4VApCa6o0Y5SNt7RJTGBz/Vi
yz+D5fA1zNhfilSHknjRSlugYogn2iTwNjE1JQE84ofzrFRtvGgLn/68dYqW
ySOrtL+mh1RTR7db0ri9jRRTceVpfAvu0of4K2Lc4cQ8SxoIH81VLm3npKoT
YNxd4kOPmvp92/CnEtb8w5Q+IbNpeqNDeeigBw5WxrZnQOtBJUhTG5nEfpvM
4o65cPqFBfQhP59bR+N2mHpfCAEZcJBV7AL8n2SxP6OWw4PyUSC4mWZplTDw
G5akLLKPD/WvGqJIH5tuW80WxK2Mh7u2YuCsp+42n4nJwpG2KjIqiOjP1arx
oPCQraz+SwQ6oC6AtT3x1k5pFAvKQKZmS0XICHfvgIiAMo7sA0aKHdfsAJyc
/plZ2pQW5ZshFOLGdGYeEaoSGSF3VHxF85OXX9QD6Gl1RCMnG5DTkM0fumdF
AHbUWZ6ogdqCfG/af41uhHwSyBIrWKce5nHHMHRDFlpWyz6y72yByaVjkkaq
yR4idmgDyllx/RpWQpMoALfzbuewUIDDKOXA6YPGjdKXZvcvLI0W9RmAdKk1
Ag3X8x+ZKybmikWB5E7qRkMkKqA4GiFsgXoblU8y8nzCjqnoouYdzmJb/oG4
iBS+cndj4LAK+SwJKYCfHSJS2bSLwfYtufUtHx8kcmbhLYz1GSWPrFEZJX2D
shH8iq1PYGuGyhuyz0Zm6+oiFHRL15KacgNIRWmK7xNGbLBHkj+wldY4HJS5
6SkXoMmGzpvk62M/DGhWUQjfPXWZJ7K1FICuyPrDSPYe7KZrZwOzSt+vlhLu
VKaxZ91Uo3avvKMzmRLWVUwaz1kiLkLDPT/TvAkI3WXgYCxljTpjEISUfOWr
TaNxiYAXw0/RCh5BXzfdI+Y9HlQLuOljGJCFctoVuYX+/cOMR9kpF+xqk7aS
zx6aodTGftzjZBTrofCocj+bUlqzvUQ6ylZbhEHxO0QQ/IghYdCyczM1Yq2U
wYO/7COPG379ANv6bsgAsZ/XuZEQjSSNiz1sOW5hTq0uAqS5diOTm1u0Q3gV
HupK6v66KZhV1+zvchn13ypVhKtdhQ4PMj0NuhL8/rscsK5rDTPpigmH2G71
PE27pmWux0HLcnW9z+Ohu2dPnSP7fPA92PPqYdG/brFmH9ZfiR50B29RUH7z
OehFPWN5Z93kiu94UnQ85TcyhulMcEvw2t9ePxcuh5nCGugt0amr5Waf8FFz
kSRmbRezDB1zPJBdVUGrGgT3aZN9ioTJnQ/LsgqrDmea8pF7m3tNYm6glVWx
EhscqS/IunF1t4cfrgSg/zIyfU7ScRxSZ1MH3VcphlXw40/O33tE5DKsCZxr
G5SbDOVTzukAVabjimThrejPDO7K/V2PLB+GUwL67zBMzcMOdTxLa3s5g2YI
Z4rLpfkc+pGaVHjEzV77015HAMyfz+xp7G7NUYYAvqLW81DDAu3CAw7rlkt0
2wLQKpYhXKQcBoKNSe+9FbE8fAfX4sseupzd1UHyyKtu15l1qQa/1TddaSO8
5bwFVhTvU/YYOCMPNt5Y0NkNFLNwS4unL36MqJHIgV6nGt/K/KJ2zL4PYlPV
Eg3DegjstIbkzOvD74So+9r92KhhUMpPsQ4qqQMG/5GcQj9DidPfbDMqGwIr
softr0XFNspepHtp+q9e4Q+Yk5VVTfno+CNrX5Fk1pBNv0v9rJ24xEQ3YSLd
7OIh/xu7aHZO/1B9QUc+5Dobpu1RrXmUrRfWBvlG2y98i/J4J1dlP9d4KFmQ
evzmBKX3FNypJIU2OaSJKlCU82GQxpUlQH15m3mTzVK1+6TAdss3PsAs34MA
XywDTPvpnbOTiOJi2SG5MAfVmtA8ZJGDgej3yfkmgzmPH3dkcAQ+GPTZHhmI
HndUE3vdDJzItfEz0SGv8RimlHfd46j5g7fHK1Qfoxpw/3+xahUXvDroL646
A8RGzikivyvcJycuMcDpiyYFF8jCs2zEU3l8zctDlHtIXn08ZZ9kW/g7de9d
fgwa9K5myGN5TOM9EXgmIRhF1JsxzLN/oGvSPJEUAvqzS4ltS3HtpCJkBjEb
KpI02dBjgcX/4byuakKy/tav81XY/hMQkGV9Qx3hgIOYWhVlqNDBP2Mii/Yu
Tn49AK7BIZeLloIux2CcPBkdrZZviSfrWFA/qcoRs0lLcdm6rcuaroLoDgJV
abCs6KP7Yj43KYmVQGTWOtB1xefIK4mCyiGMdMa9Mi8/sbcEKY+iFaglnYyf
SmwLF4W4Z25S0aUIvXacR0bVzWYWwTPbF4RXg6EAQWi6nbZJCpn1mEJtCreX
MDylBT7laoN3ZqEApxyHc6bxUrd8ZaVz0/EQIVK99mRlmLLWzfUCcP5crxn7
1GRAVzdmQg+r3GU6NYLUOjP2qj/K38DzwS/VXcpg6XGGNJOZNumwueSsteYj
x/PEIdC42XgW931EmG7UMEvUG6FT0WxIXu/fQ3DelL4p4VvudviabP9bNemL
az0L0kdstJLWiFZ2LzQQBEcIWIrG+h90XE2mnD9Iw2Uldo7tL/QZ++ubbvrx
qpnuLRqEcbKx+uz4eYw2XetTFnV/cwEBlljejiyYfz8bvs8omd9eq9+Gr00I
k1d4m/a+yR25wVHBLgWRGrv8QTCOecX+2FDJbn5PTMDahHs53XE3CmgJj4cM
j7PVSmbGtsxUxsMHUiTX3tHwzQV5WY0+lclA8+txq8gYN6S1bEnUd4Ng8JqP
T88bBdzllJs8skx/F/3e4thsoOoM0uqtpfykblvqeBCHFTWrEqHD2cEh3khc
I89NKp7DZlK+CuZASGX4MB0Gfvvq5tn6zmaUuxxb7KEWpfjbdVB+s+DffTkf
ZyKcod32CTJw56vUc7SwXHaog6tRk3DjGbJ8ClOJqJf64yoejIin/e0RpHjt
bEkNFwofJ7YU5yb2I2GG9LirAM23vTkbWE+JHnVVyvfsbTh3mFmXK9KyzT5E
W+PwLE96ri40/MZMvmaRubQa0NkmSBJV6KxB9ymSYQTVtS29emX/BatehNZb
qZ7ig8g0mMO69mNs2CNTYppdMBhOyU/PtUtig5WWTphr++h9cB179S2fz7eu
ruFIguC9Bn4aebBgZzvVGhuGaWxXDaM0AaDgYDteF0GdcrX+ElJDIZn2niIl
NpHeS+Om4z+ODciCcvjOOPux6cT9ZWEJPkrfd+mnh8hIyfVxBRYe0qY4dBI2
fkZWxm2/HoO7SP/HhWehZNiMXcvVMsayumRxUgQIHIdeMYWOFVbfLYVLVGBm
qIJ4+YdWTuOeOXIrlfUcw9e7BnQ6OzdDfjAmKO8Fc0s5JardxY97KHuNZo1t
LFWylk0/zmbq+c+0NPZbDMDeVfGjpUCfeZ1qTjqk/V061XD09bCQZI/8FRCb
t6CcdjmSWJpBowS1UAG78F6Ihr60I2hXiy/5G2q4z1nsw+gIfEXdXcjit/sC
7rpeyUrFUSsiLC51URsgwilScIwKGY7q9fxeuXloICjSxAFcqQaQadgdOVWa
K1vnc+UaSmGd/I33KZBT58VsnOJF5AZBHVimTOyuU6xSjjZc76/4GWn/NBAn
ayQU1L/1vBvat/8PmeOhEdi51VWBsrKB/idFaEzuVQ8WdHStdFDsBZWPDMHY
81Y1E+PAS91CX+hblZQkUT1t16dkUfVJhQFxqOCeI6KeY1XyU9ITAM2t41tm
h/bqXL0IxvMchn00dsCTdHOgGKdqdjndi9zPsEv14iS9aMz1u/NTTiQiXysN
a0J3X3LKAutk3yo6szgJx1EJUDcClToaHevkIK2MoWPPTzRutwtAgrJS3r8p
oOFPENps6bvZrhVl/kke3NuMWZMSQ7yX7SDNrdxwvbuKnI7w19KT5YmuOsCP
5QimnZ7yLSmXged+Bmme/xSJq/F2vh/Cvq6ccCo4zHJjJ4ZuFgBK99yRF7Cp
a+/z8vkM4ygIAxwPAKlYGaAE+rwEbe+OWcYaNZTSe58n6GI7kLtWXf/QNaIr
QSEngp4C8dm9CQj+EURxGw2WrfrmwSsLOE+DGfZA0rW/PhU8CKi+L4fjc/ok
/lrXybbNh/R+T4UoaDLFamPcl+v0ZucXc0IEpA6P3Vu19ZbjQsHVfyAeiNCy
Bi7umKNu48tlfr2mcNtE4AE3BA8JGbS1Wo50vj/8PTUSu9284ArHWtGhEtMW
vwI1pLvZ+Gm2DKEYXSgSqSrT3gbH+E9lox33gPOgK2hUC3snK5aKCyuJEW3v
zhrQB0aGrbCFCkIkFJym+m2/npAb27XBjoJw9bt2UmpKENJgbLI/NfKhvNgp
Z2LNNmMpequ8fsn9gbBQvCDewBJFgKKqcO2bMwW/JLeR9yaxDXJXQFNhY6ug
VjdCp1KsoWsIts1ZEYWQf8PPmXPGSi9bArUSw4pv2HysGWTCrWisFP0euu7X
+9vDwIgJYVjfA81pb+hIfJnkHm6itbpk+6/jV3/a+AIbL/N46S0N5FSrvsAr
N3PRxWkTtkphTug2+u6gxVh84wknL97hef29+wljvg1B//MByp5N2ooW3Laa
Ndr8daD2VK40Icz6jITOvS2gz4dZ38if7FQzJW9hIPt/fgVWj6FIJccQttWN
3zvn0DRMsKmgpS1eNxeTByZOtxNL9DnQzh1IbtR3J6l4FX+W9d6tdEU4VSHL
yhV8o7Glg/2DRWhAy0hEkhF4qLC2EC5sC+PkjORRgPYfoW+f8hyILnI6PSWO
ObEOwv2fMLp6ekGwGOzyarZf7nrCsDoDRJRSVVg+w9HQ1/rbSXRXs5RSdJuN
dsxgjfmcwjZeookCSofOuPg2f+dEGPk5ZezBiQNHpC4+s2RGnEhgedbLks+X
tcfBxbV1d01+qAUz1LnRqafwbnF3Kj1FpV2kQ1XRhVWsbAN5qU1WBpHnNTFf
W99TGK6Rph/y0hG6ua5ll7Ayr8+vZjxTnDBSsUiIUa2sn8AghzA08+aR7ZqB
jRoIAZX+6e4ahtCRqO3vyjAAMt3nYF8/sm9I561RKrY6StS2BTuc/fdBc6hw
Ve3eKV90MRvSIGX1XIb9wE+RZMy+Kduco7BVKfBosijx3qGM7Jfabhx9DE3U
R4FkR7gdbmlTqp6ZtqJOwy1k6hW/buIFuihJcbRyHqDtBeb6wKBwJONzBuGE
SJu1qhjz0mEYQephVjLXWu7gxq12/EvWmeI3ru2JWgcJiDjMP/fLJRippv0G
hHnqRXzEzqpdLyFRiVBnpGdZBz4CR7I12mG3FWJUPzfRVSP+0NIijz2SxrHf
Rg2HKoscBg5DlruJS/RNfE7Yjxy3XpkEGDGfl4V+3rvZyPGP1p0ob5a+HXcp
zV7wbrbXY5Ix2+BMzS5DPoU+uhYWTaG0tcZyphmZ4vrNI7yflhCLXktvwt9T
uAnVGXUke2EsupIkZGh13cLYMsg01dfrK9xDUfGbUZPyPg3q8YIMmsyEjxSG
yYo+Qc8AekL8Jh1EwWs3y+sCIl8xaBJclt2K1sEREoNItwtz9nYMzOGWHeny
UD43XHDW0COWpgc/TWJwUfVzH00F2NtWlUZY2o9aL83WFmGSkbNMH9V6my8p
07NiOPFm/EGW5ZJimJn0W4vYWIzFeu41JcDBPZqX8NloG7fYutOmvlDmJff2
s0U9N46jSkm23L6nvJ4kOqqBKjw5GJhYbG/bH0hRGqpS92jM8aThAeS+E/kW
V2+Rgqm6r0P3Ocge7+PgcQTk2OBmmemchnKps5oEzIArCMp5f1L2kdfRurD5
JZrIByNO08Qo5bcaDVBrmQSvIA0OZnHk8QWHVHxPGFgE73Qi1o5DjPmHGcES
7P7o6dz+qI3ZgZ1tvY5SbEg1k9eW25ASrHRlumCZU1DyK7ffrslTGQzGpjL5
+kUKQdwlgXW4aMjo2GshM7L2tv4zEUOzTeNPFm1rtmi7VHDdMfGeLvRWNVh2
G3I5HQTqofiQHOsnJp33a81wsHTWtKKaswUnFcR+f3WoYLC9YuXaP24e7vBe
+PIs2Rh+FKU7tmVmxVW4Yy10eeYbGLCuo1bP59/tJMpg9SdNZedCC2WB5CoP
fi8JJSp8hxe1UkQGn2r5g46bMJ3cU7dh1WALJWZqC/LXBo5CYwCdjJ3ZRdqX
0wzA14wZ2aF1JW8GOIdw/alPj5+aOc0mw8gW9evg6auGNBm+zh7MtRkUvC6F
e7/350f3KRnDVOF8b6gnV4xCSXQJy0eRHPVpCkyKknrn1xt3p/A/FnhN2akx
y8OeSkqTbyqfHMoEs7qTl9ZockduU2+jEoKVX4Y4+5LdNU/ct6nV4yaM3BST
xija05HQRhYCiT8aGD6tpZWCCi7vkMgWNt6WxCUR4YPSmnOVUZyow+GgAe/M
TJDZniSypWvr6D5cJjvHD3RueNBndVxRe1Flg1T6CPnouMzm64/xYR/GBf6T
E2vhJooypynRT/nLJxuFwdFL7DVxtO1v5/L9c1WxV3MS8btv0cNOtIoW94ak
OO+2XlYj8TbwU5YVp6+OQmbSflm171+SeD+GxG10QB9PZrLJWrcBUEGYsHnu
42IWnwkOvISIJVF4e8N2bC/nkQflWQEBxzmiKPm5d1ITSCzVtAlHsAU+eTVi
k5yFfb8cGlD3helkiqtA+qxa0Cy/p/pmp5cUvYXjKOWi9jTDgL7FiYSv1BxY
FKBhktxF7Nd7R0yxxvXEmW3bk2QDUYbQReDWh/A/VB/++Us0og9UFiWCIdZX
nywjOtHEqCl2z/SkzUC0/oIA5oNu/F6z5oU6y2uOWDHTot2N1qp31/V/7lGF
eMm+0yN1MwmjHifG4lSCWy1/BhRNam5Z+gd6zOvteMXpHhhnzsHzbm54InsJ
gQA3qzrLd2tcLJMLsh9pjDsc1nXjVcjNitymy2RmVOnol3lVeiHJneaLnckk
bdNwMZLCGnt8qmfXJSHZATMN02BVh0b3O10giAHtvGQV++TZ8D7rNcZaaj3U
ZLuWgutHcujpPf5SYAOTXCNwnkZvjGyyBU1eLtpLygQunnKzIbpEcQkOg5KC
00n2DoY/PJqFHYjVTfuXOTM+SJcCoDe+xKQuRRQvgPVXHzw9NbNQsjhW+wYp
Dn62ZNERi0CAUHjgg5PC4RvSmK+Aj3k185/w+Clj9/o1E3tRQuA/BpPmtsb7
NoatJNZGnLn2rbVD7mYePhOd0ythFoyaM6rRDNePMRgLVibXLnFq7fXOkswT
v80/KlNf3O9tS60PzOnJDrFkafSglnGXghNc/jXhTyjsciDZM+mMx58GKrNa
3vH0n0obd66UgCz7YWK+rCB1DiEhD0MAM3gHoRG8O4/6a6QXtOoIofGlE3/r
MLdW7HcyiKuqMNzc/LYUxVueEjQ6vsy2wvgFov8UQc1kcJte9it+QUvviI5r
e8h7mcvuTMYjPVRko2KUjNTHnU86TnjkESkBWG8aGQdRMEim54I8XYyyNR8Z
nEILb22mgjKFOWca/C+kMZktUoLzkB77JLE6ppRcXW2l7ob17Fx3W5N+1z4u
KHhmnG6bg8CyrY610SEJhRW8xHAvxgp/oCUP4tkZwcLLd1URkIoVpbXON4Jw
ONG9H67Z9qRoESwV3H9bS+8PMEN/tLFr9nBkH+IlDPFE4NrNBkecjGe8TrEm
MTN+rCQBBr0Qbxi3LZ4RbdoN8YfIhzrlsPSJmxkQFUG2OzdDlj5mN5dEmLxK
9tStyr6vl97uLmX5usvo4CAaSIrmw354BUF5EDFVhuqyb8yTxUGsSo7zBDPj
0PTiRSlsvNAdSgmAD+7nqPyhzTkLgpjgNzA+4is6xxKhq3x3iYWuA2OfDkPu
b6zvd0Pbu052hum8lgkxeFuYnbEUF1EYAnJ6GIH+909Dbnusi6c6t4RMOpjb
Cby8m7965pzVjn1iSHxZ5baStZdc7v1aYrk3ysyyW19eXOWty9Gj/ok2rbEv
e3tZWNRPO3GZZW2Ji2UGgKOrCNJI1e1H98tuMQDQlZVLfIVJCcY/2UZIlod4
IjR9p/S7h1zwdOuOiCSSxP4hZJQUn4WHLbya4a5J8jVyWtHzwuBBIE/se6ut
YMHdhN6WEmmbUbhFhXinu53QbGEwixZHnraEpVPMrrZzCvCTsMywqIZg9Z5Y
49D1Y895WQS/aXCL9bX3jm+O/cxNsUjBPSFsKubIel+XvROxNNd0hhf+sFe/
F7hLw0v8tiA4lG4Wqoev4dxtaAz9/YVHoA1rIoN0UF7lAKIJrMkNJ3g1ApJD
qRm99WX6wwr+BOGym3K473aG7Dosfsa9snORqHj0zus5v1sw14nO17IOlbE/
GLkBvrhaJ3I+RtU7Lx0FgWMUsZXDcoaRhr8rx9pVaa5NfGIjZvewagUEDbkh
TSkc09rwr5Boir9KW9uUt0YtIJbcveMQcQhD5+oURAOCRnT25PUyfuk53lJm
Umt5KhPEu9JtpLTp1HhJZ24BEu5GlK2UEuO4rJSv+QIUCpRIb+3NoQ5H+lgP
V6Ic2OxQ2R3wIVnWTgTAiWpXqN4sf7r9CDqnCkQQl3rVyv8DbMUoA74NlLPa
hcjBxsQr0DLYQ9XFlSx0Z7z2Esl+MlXK1oIozpJtuOEVvCgwEjrHknd0RUMb
B/OWa6BowgYIWqCaV///Oz66suytUCpnf9zwl92WjmQWnbwysWXFb98l3qNk
0g7hjbanys+EAgOl609/86gp7Xe5nSB35UQvgykZYlNncSakuXZInrOsJQvb
Xc5RXSigvDbyXvHEg1Nmwk4HUxlfuPVU5hrk0LVZfq29WNdFeXx/VTmz9XSK
OT2HvoQmUZjT7aw87SJMHJHJncSPPtPH4Nivr59kNx1exKP8HXhAs/gUOF4q
Pnu3KZtDv8o/I68i5+sDYedlStMNMOnmhkcML3llhIOc5KaD6Da6oOz6ZpZB
BzdPBo2kGxhwyKLIFvBTKkrpvj1Ie42iZp1PxwxhTJ+CDg4nhk0Ke9decjDI
jfhPdWtUe7Yp5Vj8nv/WOcK+g1OxvTp2PqKqSwrGQ8IyWcsXLBsyhcUozUjV
QeyJiWvKNUpNW+Ihw4lfda8jAEav995ZmfCBrmUzuEOja7a/7NfhiUVKr8At
YKBuqUhqP/+jhfqy0vYdKB+4XFpG0XC7m/XC6CaLPfENssU/vZfemnumq5ty
18V7I7rN++jeOWwtNb13lOEYevpJcX36Ahey1ohDrG7h2bM7Z7aW0n/ne134
xAp+pk5S/x51g4gHxrJV+FpvjsaRckjK+drJoMgTTcCT+ntIf2MXAmem4KWS
9T3k2XHDYNZvwNmylSDESTMSw5fRjdMt3Nn8Gnrr3wRjWYl9cXoyiiJ0YvYt
EbdNInKGLeKYnDoWcGt9/igFHg/ES9vPLWpV52OuyAwLpXKAAZpDKt6t0suE
zCErQoM3ZGLSb/bFQzBg1KEdw7TseHul/VDGHt3PXNkFuDpDsLagBdg6SysO
0vhsrRPSIfNRP9eDhZ5Mah12qGn8kfYyg0XhjemQtW2W6YYK+xEypV5X/Oi9
LWV+PsHVqZ4iZB6pmgNc/5mWSU4gHXLiWktNk5jyJjr8Qus/9P7nHxvy2UzM
mlaF7wWB1vG/zn3UkycAgsvQSExZpqHcXjvzJRk9EuyWvakxCiisLG5jZkWM
jA5vXNFbjk7TyRqgEBzmD/TOThDgNRlQZoFmTkAxyL2qhtZW1iqMnZwC/Koe
FlsC9tp2HREHlgeIJzQ4Q8KYrlAK3a0U+//fAQomgvWQGCzCfRuFaCVJORjj
3jI+HgVk0WCm1b44NTAgYrfkG9pV5xALyDRTn9qWszg+RtvYmnABwNkGWOnh
dhtWPNyLLLAe8Rtk3WMzsv2JikFJcY9YRrOR4rnbBDnInVCGJI0wgVmyI662
+lL9exdO17Wh4f9KAPO+lOKcc+qAsieF0MccyQN6WCqDUBlCNEFXI2Ir54Rt
1qZNfgAwhCrPW+vV/P8X+l6LauPupqvfkQoWhMXtO6Wwb9T73++p4ev+GmZl
+lTwfbnWeZQl8tfQc7jHTc8jkjxGUmVNTkMUSGuUtPW+vjjYs3eX9Zj2N2BK
q51XEHOnhHVdWmwuIj19rMQKZGJ/OeIfZgXpUMY8eGL+ZyPW4FGbl7y4Rn5L
7z2NlEcWT9483ljYBWidLqn0VcRcSM2StmtyEk4d/KVHj2KKzVhYYG0sXnYQ
4t92ShKO50yPLv9jh7yMyqQ/6+u0d1351OrlibDgN2xm5lzrDkX+zRbCjmoc
jLr43GPZbYra4k2D2NKKjJG7E+srNu4AKQF3tqX+HfrdQEmvPx9qr+KdPKTa
eW0CpCrPh7sBZ9lARZj6izjh1LK+wQyGIou6Us+1+vU0mxL7ZnkAjuFKLema
O4pUFHwOtrIlKQMErgNYN/WaEHxiZj2pV2Ln0WYsGwfPyqKV3IbAvicAgwsX
nPc2blcslG8+o3gDSu7QAwhTUI3IZ9P+jaqVTmZFBNfoI55LfvkKtZ8Xxiw1
iUm2+86SurJVyELSdGhH+K4K0apsOAIRGtyzTIhajUUucnMTzA1Ng8tTpApv
jL+kEWf+9itn1MbjmuzCK0jG+oyzBvGEVVCxvbaMGDkPYuFjZ/L+0jRa8niX
iwf3hkOc6yfZEUfuHClnlXd4VMfSKqsXH/smo6O19BxSRjSUbVw2yswc0Ps5
RhfA32A+gn3sfrR6+KZRBWZDTPWgcuebx6BhIuZRJMJfq2EQpyn+s39aQevC
zLtuuFoLKKnQnmYIYT661Lkv3k4BJbVzrzLxxlzke0GzmrtldJC+T2BreF1S
trJRcqVDutL/ZlxTKCf9VmH6BsZdij7GVn0iwie4IVUrxh4wUJFHdgM/Zsd2
mMdVCzHxdGB/uoa3PepSCiuJU3UyH+cg7nOAZ/H/LYIjE9J1qZvt10fHem2d
Mkzd3isgtcJuyT7fuc3Phw8U/N1sJcVH2Llho1g7MqVmpdQOAG9NVUEPsYEN
LyOw4TS9Bw8U/UPTKD6gN5iX0swHRwWEQImuLBKDucWJg3sIAIlPbkyJ+Rl2
LsZktRo82eQKuFq/8Am7BJfsAGtTGZRzrYwgfXSvzKsh6105lmbyQ8QtF6o8
flkXhSMvp1raccgVmEOojo6c9d8YokBIRaJzlOqVQvwL4m3KPzp/oI3nqiv0
C61pOPJ2UhxQR4fVvpvwpBi7VKMDY8em4HtV4/w59d1SMmLAD2aTMMafojIg
AxLkxD3tVscmda+lUA2FQRe27UrBjYidIQPAOTVO8uZvGOyfXs9tiglQVwNn
UEqO+/qWCjKo8enm1kdxq4b9Z5gG57kalcfcEbPGdDfvXAWNM2xcQGZVQ8r5
5jIWXKoG+Um61AIh2uky8No48N07B5QgIp1OYAqxM7GVD9AZZNUWKxAI1CVV
daoMmjHPlQRyqsgiI5y3jJS56g9XqsQGUwt+yvNfFSISFcsGlr4OtloRT6OY
Q8GrBgmecNZQkLKyE5l0l+/upntfa6F4Kc+xrKCp42oXiVeTnddHlsEWt1nh
G9TsSd54ZOOtMqWC6At6PVv0AwFrKYhLCCFsM/Zr8+0KN+ZDkQ4SqvZrDREM
B7cOHDxgv5q8cuEDvrkS/tbrWv5PCfEI6hp1E2kNrV0sT4OL2vbpV2MevRf+
/KX3vVnuNqGKwCcZtViCV3vMCx/2iAUC24B+h3Mylk1bvHReblZ8QKnPNxeP
I50zAslA5rzFFymMSmPr1lGEeG20MxoCp1btR8PLiGOPsRQaxgxK0HJPUKJI
VBgmIvm5qrNlNrGqp1lK43vKTQV13ZQlwLG+4NuQ/PgaZdlCdW1EmEPVL3wD
fnX7OGo4C4488L8P/6EA/Gu81oBCRsi7qBnQpT8vXiGoB3MANFIWgH2aA8mM
gtE/bmmIL8mz38Pqz31gq3mCAOUQ6AmrkPevn+t85ro1UX53wgxagJzTwC0W
pUlpvv7HzB2+sI5WAAckl32WuVYhxQryAFaqkW6EoY3acf/L3TmEcbsBbC3c
bMXdTx5UV1S3jo/t/qk7bt0DtPl6yhYu8gUy8tvFPJbK69rK23SmWlcsvGjg
Gr8h2V6T1wv93Gb0Fxg0q9Z/pTpiPLA664Xia6phbMN0WZdxWMRc8L1SJWh0
wajtLYVlIplBH6Mrz++XCeQVSD52nB8jdf2Y3wyRIAM+VO0VyB18xw34x+e9
2kVA1ax+4Gcqta8GrTcaZgm86opp9LCX9XclZcDB5SJ9mXgw9W1XnkMswR2B
pTCqvq1q22+9gl9OJAl9nRZTaihQGXPIDyRIZB3ECPhQHmG1asw0BT/fAHRs
Hw7xCc4xtGRp7W6FqFZP8/W2DtDkUueYvZdhmYPp6VeXnE9m/UveLDJCHyXO
PoR6ZYALY+6/dWrGA8iCVtEd9LhKBN2qeRBIexYWCYKfKckRmcEovMdwfkdi
gXiTi/gqeGbz67U5/FRQjL59GD7q8WEMjyaPMiIfw/PXqiMXtt69a01XcNoB
P1PkM6pD7PySulpGDcjUYQf5minMKy4AgPzB/fmo1F17btqOySfH1p2q2SHY
XZDQHJJE7ImBrLuo9FDCxhQtTFrD4ZTKOGM5H1t0vfC3R7H1BVymfMWQshXx
sfKROyDmK6S05MeVzP0bfmoX4BlqHugH0tfzjjCtcPJmFWe2Q8kCMCxkYBWA
50tmuAAUOMnBbJjS0kTCJtYOrV9Hf+aSlcE6tHs0ORjrIMTUtADk9+9gNlhF
7xEcQlKxqgNis1aJ7Rr3y7ueITkYbNtaMP/wNL0Qcn2PsD5rVKzDLANhL17p
/VDm6VD52u9WkOz7Q1pOhdb7/4N7VymyPPr72YSQmS6oX7kyXefMozgp5z3J
6FLpyrMiUD5h9Feyc+iYkLT/psg2R22XU62PoK7ENrGkIyt3YpJYwaCDzcTJ
UOywn0FhcJ7lWDgh4zqSXjOXu6mbxkOtVimsVc3n+tBE34sNQl71Id672qFp
YoxV1H9NbDGCxIf67GaifLfq4JDCAiRVrdWORYlyOXfyDhWrikL3GigqJfTJ
6ndaKcFlv0cLpuSfQP0rYXSXYLyLGHcbpStkvoc9LZhLtG/q6U8LPZI0qagA
um1qGxNVlAbOxHZnTvV6C7MXqwoSbqOjXH8HeE0f1jY8wHauKWQPYmSOO82L
0g95X/cDvLLNZ7TgKUuRTBt4uKC9xdbnQlcze7uT/MdN+uDAbAsAgqB7V496
7h5SqODwVDMNwxmGYmCOL6QkaR6toUIJeVrTyqkcr16QmnB+wHwkZfG5zP0g
i4CLCLb15yj+MuWt2A2TL4hvbHy1YNxtweTcMeqMu2MklfYmQ/EUkdUKAMGj
pqE8Rx/oE93ZG4Wo2YVKpVLEUbGMY4zxpSBxLYKVCYSJ+PDAhp2p6XsOW/nG
daNwCwoUwPF1Okxu28o3cJrZ0JQnjKvVaUxIE0g3I6HLJXhAnSMVhk/HxeJO
urzkYHcuS+h9R0vEvdtcZTlfE/qqiif2F3PIIQXw4PAwMd4lQgrbZqBrmxPw
A2xoN004+mJfasJD0zwdsXPAkwDDPueCQKUDWvz5xgDvDAWBgGfhBtEIQ+v1
gjPcmrzqtukzm+v2XyfR6N16d6J/J3l6VsOd7HbRdalaDJprkth7yl0R3dNH
OccCQpq3uq3UM8bwBC5FXOmOb3A74/lPZaWRduLnXoZS2NcR4G5naV5BXbx/
mdo+f8u/lFdWlQk9IckS4csMlvDZz14st8ErSvQi9TzDg75D8xcsgGgKoQFU
pxUJpXiZucv/kuPpOtYiK3/jCR4R820jSI74LeXrXnv6WVMacCh6BcXGjdCL
F73neBhsQGTkoTgDqU6vAS8Bt0uIJWa0x90CNJbZtfclQ78fmolXOMT4Rw/i
APYOdR9a8gQ4aO8CudMH7l0IAQDIEv2XW8VmV9S1Am80KW8Xp+KMoEZ+eYmY
U8lv8hO4aKNKKcUQFmQXWz3yRMWG8o0qzfwjVwE9rhYc4bdTSkvi/B58KI9R
j6ZK9xxzUzsgXbfcCvvX9hc+Dp0C0nJs2YuswKmeuvbMu1jJM3uf+xCI3vDX
aeA/9z8KUoUtX8VQ+OLotOkwpkf+n3SKYmiwRnyCLmweDq8eumCGVcTDFVp0
q5K2FXIHuDN8V7dNbxtQaWbh1b6YPEw6R6BDkat4RBoZWZIeJm7o2DzwJadb
b+kD+EhT6hl8bi6h9S7y1IXcoCIsp7SQLBHqK43CX/RLrprWT0GmP3s6Z0TO
LKDhx/WEffqNceZKq1cmaCXoa80iW6V8LaThCB1tKfrTFoqO/7JGe94mh7w+
VGv4G+5kkt4qpAgvAMVgppECKTCWzR9/6RnISCTxQzmvj8lVbBmTswTuchsV
SygIx6/hSlYrxZDPb5BhefV1iSkHD5ERqrxe9jyIY2vxtUnxJSgB2oNHRS59
564tOH9kBnJmqf/90n/1xOYqrgGkwyd/4Gyi7F4VMjDnQotbxN2TVmryWega
15VN1cK2Wlh185esbvbGJqrhXKRTdLzA+qPhE8XiJyXTn6z/FhpIE81ZMLL/
BxbLftTkvBrd3wacktAA/2l6m/lxr8zy6eTmZLzFz6/82q6rxOtP9ErfCOyJ
aLPZlF7Seaf8wkyqzuNQJeH4sJcoWP4QufmpPUqGf7NyQnOe8DuMXg4/QYhB
OpFBeNQ1figFLsSVh+ou4uPdt6YX9YnO8JEMF8s3NRir2HP59NW/UhIUbgSn
VpcEYyrWmvpI0wTvwoRvQupc2XV1V1lTg7N50E/UMlmLFuZQiE4KHU0gNqub
ZP8pz82tD96XsqhCfHFYvp9USZRPemb8qVfosLhABby5cxWztUdsADmRe/Br
Ql2bskJD3sunhtkdTEwPn1KdSAI0IrhPpQsoSnbgNAaq2EVkbll814h+6R6M
0lMJo6R8pZcLO5aSJTmMG4MV+8DDxjRwk5E+/66ZqA0b2EgMpih46f5d6Tn4
Yc7y2fAMHqOdKIoWSyVtkOfKlO/kUDtVft9EnwJmk61gGIg9Cgvuj0R0kQVH
itOeEhDZRt4+qVmYEDCAG4cVZESjeYn8GEOjGLuJIvkoepBcivnxs33weact
C82i14sOmqKi2DRHMotCE5yuvSAEEiwUhfwbenlGvcQ96LeVW6u8zUjaXV3B
saawWQ6PLNN4S5LwgDA8VQvmfMcpA8/5P4uYfy+l+BYpSJJMFUM8z5LNMQQw
OdZUVDK3wOG50cqQBkDt0OMA8TaSZkvwuC1Sag09WcmJhi+lBwOWmPgyc328
eWRLQ1kz06jKEdrGv+5Zp54yjLasHoTYW6Fk6GfapAPE8xEn8yZeFXsZ2nBm
aJmXF7+hWrnZwT7RpU3DESNrmXeKs3KhZDYj432bnb491f0076nvpri6dqQB
ly2hY9ZX/FFJb9VVzpOR3Dsdaw3tE0EyXqGhKfg6JJu/qQEAwNC2Pof0f6+Q
StvsIXfBMm5gyU6njZpgZpQHz1ETsZGIhwjys5TZQLIPTemR7hA3DIVV7tp6
8Yowt0nOmJRPsco9z1fIfi2kZekjY4J/3kG1U1ZS0qgEUOceDI3DHbp9PEof
YfIRwHENQPuJbh7BsBpmMGruM1bDdZBg17aCIfQciGuDXOhtFjBj1mhx23G5
DDq3vyZgNvHXIBCJF6rhDbZaWV4w0brxBp34Rb+rTCwHnQC06ofRetfSI09j
Ym3nkQ+8RqJP247kBFHD9Ns0XntCWW82Yk8NeEZuEetKn+IyFT6m6q2vX2pq
Cbx1zewwAMGL6h3jKqQOxYq8qxj/91fLEXmzx8CmwmkrRtyKvC6jT02M9aLv
xwoe9g2qAGrxUBJT+viLx9Ueph6e2qIhYuza0l0e7dNvxhzToJuupbF/tWE/
ydyYeUn/vc68pSH+/RA2tGgB8jHo5h/xEK4mA08Ci7HZdsiS3nqFtAj3BMtN
9IDqzq5/dDkbHjEP/6NIcna/CookyPyViZ0Azsf9o8rSaFI51v6nKrmHLYS5
QbW5wHo890w95m8vF3YJHckQ4B87DY9a4Vvdi4yLDm/K7JHlkKi5RlflRMF+
amhKOZCczX5xEzGADm07eaRoPGOkU4vaaA2RKW+nWx4JgB3l9PbPoCDolTVj
OqAP5SG5iMAcM/rhU+DR83L9pAJ7bXLQfkUCoQxIaxHolI5Adc1wxZo2HJfa
lDul61qTpDvlg0EfKViVVvS0t3jtvlfCitWBWLluIg+M4NyC7vECt3LiQl0L
kYx/TjuxbreD3ZUUlRjpQ8U7lFwdSfu4bkiMImCakB4X9AthEilgGGAdMQcd
ivaN8D7n/rSq2V+hj28G+njz8fQjFJjEUZa8qKgObY2mAsdrevW7jh0Ctt5t
gLDiZrZ+TSR5bCwVMhpNopSRKpNIK9XstiVZ6WtoqGVvWeQ13Ps/wr85+miB
WIk/sdFHqm9H37M17Rxn5m1Nw/A1EzNgUpx6mDPYdNtqXjjO57L2ow7R2TsR
d0VS+P640Uxgd4lgKPVLwrNdImekF/RLwQIQRJBDTd40RzpErMfpF2687QyS
Ui+TSbjz+KleX+aqaN8DMFWIqSmZ/HIQ1n7WfrbrKckQBcTSj1O6aE0gJVHW
UsTmcZCO26CQKGA/JhDOUoUpx1lds4zzemj2kWhC8Ba6sjRkHsWYNCi+yYz0
jQqVGLO2cpbfy8zce7IMAeY3k7lPuFRNzcjLWyr1yEFiUvI1wCwDXpri0boC
s6yyDeZdEokSgBD+WrIPc4rNIhSBXMp99CpQZdW2dV089QTJ2KKkwl0nYiGn
lza7KlmzAxIZeaPSpSOioYs2bBi7n/4umn3aYvg6w99r1BGD+pjXsh648tsE
BbY/epfgWJfn6IkXyVyIXrD9b7FLoEhip5/adxuhgoHjPLZKVFJyNL1gudpT
itVYvmVcS5RLwdVFZLBCnAEGFUqSLRxByB7sfdFd6OK/TkNQfCRahRghHLgd
71wOFWsn/+JQOSTKatMbKqk+/J8HQB4vEhYs5vmtNIqtuO0/mcr71EKvPET7
hghLr1G/vu06Mcf11Va4MpS1hniVWJr7yGFV80MK+OOgLh7B3mv/B1SRMZHJ
LqZZhrQYzbKEpHY+oTM+tOE3h4y/WJRVr8SuVTaFz5SnAZ7nXNEA13mj+zy7
R14VJ6abg2P1xPppclcidmJ/XZ87+myS1LMjCXI7hikWPCRKESPdPOyqZcfc
+vEWwEtcvxejymgRkxc5tCQJJKfaqF3WaA2FtWCSrBf49N7kzZSFUcpgVe+1
1zR9BVITtS/7yFZdfFt3tHCENa2TLmV/6Apnu+JfKALjvppIHoDO57J7C4HK
I6GTbz1N88MbuGq+tfsd3iNzx4FtajHt275TJEuZQTVE9GrY2FZxuB0/6ybq
cahvR01T4eSIaHo2xh4zDSJtL3mwJgXQaxvoY2fzBh9P7q9DR/58s6xp/+1N
P7SXDq/YQ1hzoKkoxYL0/l6RR7ThVOQ4/LpHEQDEri25rqzcPTNiwXfGSRs6
Vr1RsRg4oBrmFk3Q1lkKU0ZSq+Mjyc5iqRX2SdJltBlsMm2YPAI4c8HvQQUM
quQ8jDbeBnYNsKTXMmgfPW+KIyVOFvXBTy1dvqOg5jRFKG427JH3fK7IVheB
ZSOJUHOcpEk/+noHgqbK0NyNVA2qlTfGYq7JLpw/tBTPmb6ygyvbW2cXVeco
jijFNa0zSUcM0GXq6RTakxD1BPe8GEYH3ZFpHa9xdzd7niHkAAAC/bygU7WC
xxt5fJbinL3ZqJqb0K71M9pF7bz4bK+jodITyybeWNZkq+kl6hXRoZhxdANZ
YhaWHBI3QZdT1anHkd7h6RXVh2PYFdP9rHTXeegi1QsIOO00tKnFypuxei/+
XXD3YDhGLA2wd8jNJsBG+Ir9LwvFHBPCPisE7rQCNHJYKmdPm6gzDC2v3Vin
x7KlzzZp3BIqxBaBnT1t7nZ60VDC3PKDxKzd6FJ6f71XNkdw/xStPFTWXRfK
4lYjCvwXYjN4RKnM77o2UTWgk48335pHIs2yu2wYIbeWE2kxfATc8cxwxnbj
6OTpQgDXNQvorlfwPtZkX1i8cwfCoyz3L5QyjotLAwwThZO9TBzkiX51fwxR
Zkv4WcaLr6BYCl+Au6XxWGP8vwLNce8KZhaLO+uc7M7gW+8reHkMbjhIFRh3
y2E3zYxGHiuVRlzUO5KRAxVgeMEaWhsvma5rSQh3pJqNfgFSZveed4vBpQgE
wBs7JFfTowwGW3cDc3yqdiHmx7bg7liys4lthmiRRecOHqxAlDuU94N8n7c6
uwf3Vsi3pj09i46L+IbO5HmczUasm5mBPvoSDKYP3MkDkR3EjinFFDpbXWSV
oDm+f8lUR+PyK/v5RjTQ4gK1f79n4J5HWKwIaaXLysUxe6+8J7pem1XIQPNA
kD2z0gqmw60+/ajOTqiawnnySYE9r73uGECKh1PcF+TLCjw6ErGO7H83EVAE
TKPAhfBUpWV3Va+Sxf74ltm4NfbLbYoaZo1Trrht+/mcqwcj0xKGDPVi6k4Z
mSj4NKeRmMIQesryFrNwkzfX+ZsrepYLb446oQwYhk12Jc/jfqdYB10nFlN8
65eMD2jK+EsoLbaz7c10B1WUyc/28X2nOK61XCjidu+ypf4fQXrQ3iro7nwI
Om5mUm94J/Z/P9kfWYZyTlAk6iLv8hnpdQyMlkEDWyj/E6IKxsHTTm/aA+RF
5/62MbBgm5xJvHJQY7tTcXHA4qsnKNnhXNm/+K5EdDTnzNraoAlq6JglV1t2
AFNVbc6nclCk3Ec5t3Q/cf4s8GHdkOL9l/IPolztnq5e0k3bjXWyU61BeX21
DoF5JmpdLFnjq+AlulhIU6pSSNM7c+VClYn+aMmzxqqdbojpqOChTNU0670Y
vItEuy0OVr58crpUYLXPBtZK0oVqXmrlJrVRRagESPwD8wnC/66I0aAGCieP
xFgN9/cz17q8gHhhiwugKCwNQOXIextYpfDkUMpnfM3HZAdAnb2794cc9cyL
+SgpEnebqTCdhhvnd9VKD1Bixpe6UWNqet4s+EaQrZyRTo/BIuVNA9R7IAV3
a3kErYTCvT4UFUeADs7zFpNRIIXns7ywaj2vYPJQ0cjlrv83HwWxbFlzlHI1
UGtX8SmhTDsnUD8l6g1uk4BZOWHk4Va6SvWyLssf1zxwaaQntqBcnVJLA0p4
eB6xHlT8JGxis/Cg1mBRSu/Q8nbUDUfex+Yxw4iitkzLnu4E3lJiKLwGcd9u
6MPaAeRRCtkC95vuuRr5/cEwnCQIGaok/EYOPstqhzB8ilvd2K9ll91Bdt9D
afBFS4JmxIeljrtA9ofZxSO8OftT2O+xdR6rJkzHozADC2q0matyeFUSEbIf
ZYv3s/jW9r/r+P7rHkAsknabaexWjhokWxLxUH4nP34+MmnobEO4D4Ha0umo
ayaKaXudTLYSOldWRK4NGaiHH5upERCdME5ZhqDIEQe9G2SVnG4E9kX0SOQo
sZAlYUVn2dzpHFmxXb1ubTJpRKtBENyIZK0f8n0Dh7v8t01WNPe0t2a9Ng9e
267esnf7AjKnQrbROaOGIs9Z2dE77W6KPI5t7LDPMtqeglXfXWuDkCh/CRqy
ymLOIA8fPku+L//d+Lm8md4FCIAEPtBolLbdByrYHzdJ12HAfVAGmi8MN/MK
hjnTlPMVo1OW9bY832NZoI/WfTZl5H2esYu5jl0uxC1AVTdXnZhNqTxOmdw/
vm7MXe3shkyD5cMJVmEWPw5vOj9DIKZW9O3yMH51ymCSnhqBnoVbOFHTsAxP
HtVLAgtHPTmmAj0LwEtn2Doub8hwJ1e5GG4WkFzmahMav769vYl/dcmYTnJP
DsFbeznGIvKE8+UzWS1rISBHFhyYbDtEb0j6wBPILBE4uzZF6dYIwCEnOuIN
cRPddtXaso7qoSWMGxMAXQYoau/w/VLYjCyOQj+ITm5MMviEm5rX9KCTO370
w8Iw6faNAy7OtqfjHejlsvFC7LixeJhZndwqBVK6V6NrZkpvzKkouYOt+AH8
Zq7hxlh3YiQ+f4HdKD3EfDK3w7dlIfSu5RHvt3LVrxXmsWrugyhoIfHTn1LY
trIRUMYqQpAfjXgV2DBEOykLeu+9X43amsBZuH4GkpclVSQhyel8dIm+sni/
a4iGfnrcVi/Q3Zst3a5h9ojMh24c1TUiQvaxaf8cw6bqPEd0J2lNjpmQqyPK
jkbhw2NKCxypgGRQolL9lUp8nlFwjoDd9WHFUF2MNGqhjHW3K7GyVkJqdGWI
8/vFWRkaSr/+Zmift6Fnc9OVjbk3GaOQOMJNxlyoTdAkU7uLc/6T+onIPjuW
85+6opbAFNmzPBCZncJYXObTuyeWBiuJ+Vmrf4D/0FJm5A2rhEJRIUu7De6j
FErX6Jc6LMmV0/dpptxq8PjQQNuXArsDmyJJV88UxMKOVzYeAGv8xLfjVEdl
Kba40NmX/+vamjGUzcErgx5xaUTCL0RW+18vtOtnNIxlC0zeLdRYDVXW91AC
sqOI8AQDKN933twoFL+kPkanoxciM+ARRh2kUxwttzPbxm0+2rN3F+iVmvoE
wfQhpJJyzmXQ4aPqChP4F2z0SsfkQMqrOc3aYDdd2BRSQXRts/ewBJ3hSvlX
tVF3JAPv5SBdc6jOUTx+kuOHMt7qfqdLTFVmqDvPg1zycdEBIRDXfsUWXT31
2kku3AJA8ug9ik0ic6OTysZtM3PkF78x5VicvKKTAJoW7ap1eN17pdcVsezX
X7SBEq83cdGe/JKcYUvXG1Z+/WvkpeN99/Xp9Zs/B1G4jo8F/o8Hhgs7afXZ
hwoezDZU1ODtd3nGhNiF4iJs1hC1gHFagdqhBzamWbPMf0YY05wYTb3yCKvR
5wwu+FKNzFFqqierAwLIV5tZD+jC+OcV5uSepidJGUskzn5ebXG1FRkm7n9i
ojOqWb7Sl8bTG53UkbQJoH+q4zflwoH88IYuN4YbTHyT4wzGpvriHnG903vF
jZgA97nTyZN845ZUgx/2K1Wmm1KrfXgjtkemisHOi7B6Fk55TmYsxGjinRTe
gLRRXXTavqO7JfKfBhilbZ2+th6uvdZ6/6eSRW5aaO5evoX9cn2rqV17HHSs
11wraVa5QvjyaJmS1XHrOIfHrkU/SsiGlG/5kwkdeKkH03cSgxkIbNpjC2wM
yOg9+3xneIeNNxMtNQaRZbRq0Wa5mJtfTX+RlSnCqkqpT5ntrarDX6Nf5nqw
NIihiiEyyStGWshhzLI+jglTpKLurMbwTvFKCrpmSNk1ezHhcbiee2Rq5hGN
QIqI8AEAHRfnCwfroSaJotQXqwiOs5yZQDbzic+mzj+gIoSQEWkBvGql4jw8
89m4G7x+dE5UMCz4JPQ5quZehTmtw6wybEYU8/eSHaGOmMoHj0SnB6a3MPQR
vlDGcs2/9oARDtLoysfbnP8dYTOGzv0zJibfKxMc/i+llbBZqTk+3augfZ42
gKn0TXFm54hrBVVOFK8tra2d9iDetO/6H9hgq53RhgEYw3GiZdyavxIBxg+l
wi8UDjElb+1dDhQJAicLoctn1am6cpeVchfh1wrJEKUaykJqJmNHyc4QA2oa
mwK4QILnNqd68r9R2VNOOPBzToHZEJMKwHko5aISQSf1EHDeEetBeSrSGzXu
Rqnl4Q8/t2krlBY9n21n9frtC1i0e7r77NtT+6BcaBroLnCKYPEtIHlO4irs
Gt09aMuiOFEylN83+5m9nvS5rIrgjf2zkaRF5URxu9RSk+hTFrimPAL+O2fT
L/wVMu2aYoSf81HiEemz5JZRRGtgf3NuPAidMXMBcsgigEGx1btqLSmprZgY
XKL8oIVXbfyQ2QNsE4MKgOCs7mlZMdKtF7vEJh+YYinbHFw/j2RxGxa/TX/A
n2DLDP26pgX1gQQ4vu57nonvwfwL5mPe37wpJRmTEa1Nagk3xHQ8wOpPooYj
xz1XQsxy6cAizRxTFtEjXdERNwWpp8mtgcD6Xsvz6AYjyhyuKMiD12mECRc0
Eo/YBns8ETYW6mF3+lowYzYSqksYw7LbwTtZY0LuYXd2z3z9MYZdO8cWjfZ6
mBzcvcPe90NOOapyjHH9sVxBF4Krz1yIR++2AKNIVhJhp43zBd7YIUI7/ZxN
y0x/hq792/NdO21wxmcXMnoL02cTnX1P1dwkPTmFzyuWCNHcwGb4WVFFSqMV
hArxyL8ZGF+l2n+KxW+/B5gEhQXxqDrzqGQDaTpEas5NqHV01cDBB/d05aJp
n+xouWE90GE4fxbJaMMVZm6agIzg0SIyGtqt6LX8UFOUwSMO/GWUlJxbp0G/
zrW2vbspezHG6dJErcIfalSmKqrCLFwSHZ+kMjC37d5/053lp4X9U01MDDEs
jb7Le8W8G5Te1QsaNVlGZdOIaW7imJzEgnj+UirBBaFSUa7MOTu5vVFHD9Gx
5XsFitnHJBuO6KP5Oe0bPFrRZKm4iZfrGJOYnCVITHlRMMIkks3DEvmPWzv0
508N5FyMk/YLu+AyW+SJuyEiHhcdMlzV9gn+FNeiQe7g6sB71V6qWVc4YXjs
VEzPbOlpO1cpXCzYELXrxzuK2RUekp7upqOW0kp8yYJx7cHzERyJOeU0xVnY
0MBtBZEFHICiZ65Qm1YqeFe872GyBrjVK19yMoc4d4Jh+i8pfT0jMjPEdW9G
Zr8XkQgiai4vxh+Hw+BrZH5YLZV/GcjEbb27geFZ+m3G+lQm8ZjQu6hewI+C
b9UVkdcY5igHmxIeo2Y/Gzk5+8l7YqrvaqMmO095N7SHHuFKY4Vy8MT06DuO
3II43JEHQqDsknuO1WUFjgflFI4K122xqkmWQ+hPLAMyCJo0z8DNF6Tv3/X4
Z/RGssI0SFLuwPlO+K7d9L0qae0lf5mC0lLtgez7rpeDyoG5YE1vCHgrzBtB
XOtLK4Gx2K0dUrZe4fa7ew/Kl3oS8CAzIvt20UOAlN0HqGevvMnX7H2Nb5Zt
+pcTXtWrxRx2gA5Yzux0KoE4qxlZE/eWP1mgY4lFfqBgSqOk6yOSSxCXxydm
hH3DapiXLhAD3aMN1CC+PySr+h60vcxck8VhagA7Gg1OuRjqMT+0QS+5T2pi
qAd57CDRtes1dgFdL3sEQq+IhzRRpoX5abdJ3rYJY3+pWgUC1DuKOiIIl0P3
lvt/mr/O7H5F8NUMRjoT3MbzDUsy7qkwWjsHQHB4eX/6Lerr6lGE2bR5d87U
FxSXs9T/kFxnnemWWq87+0nGnEDKjsQsCJcHIiFVK0493Q38yKhoUNwHQ+pO
KbPY/COPRLuQXrmbKoVVI5XQUTrI6BAaV2a6920d69bFxCOseqqfbGGGp04N
Rib6iNflvLVqBxZxBlv+9k+Uv3O1INLfREZNoimmd0TGKX69AfnyYINgsibr
YqRiHmG/oJ7G+f/5gTAzLJ5jzXrK7TPbdoHyizqXTCrnQXHpGyl/z2iKFW5i
vPRwZd+bWzsW0blFvEEe/t5ln/XYGEY5oHHFEZ5jnPg5VYg05dfi6lkTt+lB
LP9xzbY2f+f1b97uGpp7zAYSUE2+swCYWdyQBCy3shnehZ/dLy2le99y03Hd
j1F31JT634GTbNdjWvEgVbnc0gjGCDRjyeoolaPO1lHw4ndXpQdT8wSJIEiN
5BRTLryjUzkob1sSGLMBUJFRilQhc0hnC+pX8q9wxzCCJ+Vpv+zMGF15MRZ1
XELJMmTiM+8WlpW2zUlsnlLoz1FbLQLUkLXhs+Dy2lHnA5qQnWjxqZGE1p04
0LI6kQzHsUrYAWrHjJdzoE9Em3DEgEpuRb5b1perKoF0Z0AyrIgT2KjYUqlY
aBr20ejMaeKI3oR8stusWklj/b7t/ZlaWQnMKX8HHUJ/HWwKvVKd2YlyxHxN
IWkLBz5vhwLE/F1snKIHGURFFidQdbb20pdHi6KbQeCkdlmXFlTEawMMsxHO
tV3/2Tb/P43diE1QQtjUBbtkBYDCWvOoa92/AdlkShqzxtly9Zbljt/vYiTz
nV9Q2lvaBttLiDr8enCrrtFm+CA2PniZUE+uo7Ywog4R4I+zrGGQ3ld3kbio
qCLpyvb2v6mInRNPJO6bRXdmHm/95S2XmtNkmQfNz+ISARINvjgbKyamShag
lh9FUkGIUhOwnnNh9lZMzv8hEgmiSBPQMd6/3hk2eW6o+H7TX97d03fPqc4E
KboqzgRRnmkMVXBkdnly2Lqxljd6R0ROEiYJKG3CgHf25TeJdQ+s9bLPwdEC
n1QJ7q/A5CQ1xwQ3cnkcCtdkpCbZARDhOKJ32us5tPishrKzxoh5DxcXuXZP
D7cW/SO5mfs82fHhY3q2sXj7FzWn59717acZC9u+A7RgZzrfIrMkT5Fs2+C7
SDMnLHf3yRKACFLXrWw1FiHOuJ0EsrsKU5eSrHcWBWXGZe9qrIDWpckZJ0yX
JSt8E+zMW71A0Jj0IHpDtTY2KubD2yXFYwkXIJwxgLO2G9hIAFdNQwlYCNM5
cLlTdez9wsNBFvZm21k40D7cv+vJSFqhkjsjPGPDr997810C+mg1KW2GTLut
4uOWsuz5fT6OeRGFPFi75tf2ZqKJxCxxeFZVTdY3mpUGfbPR5HX87piadX6k
NeJv/oYNmDQZwt8UZ8Kas72gfgSwERs9itNfJoeIC4gs9grBc9rXVmaK2Ru0
7+imNO+FoPyd1nh4tS0L3nyipm087/UHkvfXa9JNAkBUdj0HGeZnHokQ0XIL
ZlmQcu3gcXdX8YdFQv/89/BRLMEQBWgU940YeZDhxx9CYkJeLF3VLyUz7Kw5
sIfVPK4gNJIY8nAaEB2L0luNP95EEl+zU1YxRAudL8gS5deZeEHKQugsMo4T
PYPCMh79/1hOxUEnEYLBS9kX7KESAgt5cilwx1ejzzgHXD9m7s9Eq0vHmETZ
Kt7ntkSbMQ+W0NslexwBBNew8y1Yl5DM4l67AVZAQTAL6dFc4NZxSIo6Kp8q
plJJW59NI4fROi9dz5I56XMJNUhhlgbXQIEyNK6BAFQThSoZxX0jlvcupFm/
LdU7C0Qj0IN6vV1gjgoORYv0jsroozqz3mKumAo3wr+fydjmt9W+K2fkMXAx
WR3RPkEnBssNv3cZCUilH2nhNl5fkg+qkrJosrhVLJ5P9kVB/FvW3Vc6Zg6f
iNPpCtpHhGLFAHf1OXrVimDEcX2/x9iLXG/sioYDAZAXLKofJdl+XsVUEoko
Fk/tsdmHYJTL4Z4IpZx6q1q/KXfNnnTmXXzybuV/t7DBi0J1Gf0sFHxB2WYj
bn2t8Sx//eK/QNSa5NSJZ1ZPewwNoNETWk4svzTH8PTQSgr7VsmCazGtqOqC
WiCsS6iNfIKqgz6wwOpQihSdG8ynoKxw0/NHDJiyt6V9WDTk4g4ZxLKRDJk0
9uzhFzJoiEXHDlrYsf2HhprMiPgnB7EULJvSU6sqOJJfy73H639ICqKwsa7e
iq17DGkyTEj3cwegOFSyhFWxYmpLluqr3ZQnEoU+KXCn7XqRa0BBWoqCGKWE
vpngAOJolkZD5buuU9IDdiHTibIvhNw4gYXdZo9C8SLCCdLNADlInclqfM0i
tAXwVtvVGT5VnnOI+drAGpvFOFGOHZS0TGMRTsvDji5X/KJKzLIiTMRefaGS
tOSWEz10EFBo8aAoyHnLnypd0hiqoSYzkcPg48T01dC0Qg73pnuwzgCV9s1A
CXAQz66xgOMJ9xRHNVuGiPXSKxhFZo4ww2ENglOKMOKz2/mav1MMJIqbhEsQ
EZHOKPuLn7nwHR/XPZOyghBgB+pnoVCrelnDW7FOs8SBrg6ngZjfu3jEFkvf
7o6ZzETteWE/5F9CqSy8N15gkWbNgA1pHe/E3JsB37vJANnLJTMly2ZqxBu4
3IV3bgricvuTKdnoxRgHP5RCvdhPMInY+MTfFSw4nOoMUNNOornvEAdR6VMN
4falK6+SQF3HOYrqmGyWwk8wnBkC5eyNbOJirj0gpuL3qw/aAdz5R6Bt20Gk
2Qi5lJASPqY0L4JF4FVnyEZ/bDQO7sOw9prhx8haEhLgOkvIj9ViW+tVfBnv
LacONRf+0HHksP8VCer2pb3g1rISBq3kdm+SSc9KoHSvghyerrWxlhBIpZGY
1rAdnriPoIskgT+rNJaKX98UQyyw49x12FUke1ljrs7AJf9ZR41JAUBfHPij
I+QUxS2D09MtddZ9H51BLdbPuE39PhFCeniTukqi9tyR+Tq4fL4hkY/eY0ah
aM/p/aZ9rhbqzHQnTHiaXNKdqQ/TEsK7t2wBMRw45OuMNnO1IEwfOK2gl7pG
+gEdcI5WUsWiLUZtO2IVNrN+niKXsrtVrYml25ruGYYGT1F/hrMEReNjkB2y
4dLgLClCHYwqOM3U67iKXoOBXs9YExztbIIbIEhssWVolTk19Ld3Qjuxl/Jg
4+QW8yBTi2h6k/1gIbx7h/M7C2+Cem1llP/gifNe0IfZlFxDtPuzaWPQNdp1
T0+S54F8hA8lsFcrGEJZmy7WwWXWygU7V6qE4fW1jnke8fSJl4UDOvo6XME5
qfbVXQhMy7loiN5Ht8ibynGdYQP2XBaMXnEQryjtTT7v/Rd28xJhHFQ6kfdk
HTYAHcP1lg5hb8GzVMEMsumHqi229SgWdrsQ/DL+lsAT5Ko3/e4V3DmvBZiM
0DPIR4Aw2Cq05kFxLt31iGnRE2/oSGVK4b78aeqjUIJO6Ppzkxvdtr/UNpAP
eyTVYdhhLLvQeeoS4ywnh1/JUJjaTWJxjmZrGQWMb2kxxRPxQAgFNQ6pQ5DM
No9NFBlNtTRGiMGPeDJGvktwN4yMT4jWhN5alEhhSzpajrPXj6lb+mnajB9+
TlknBlHnaeTLoy6HZhz45WaS1yjyNy6Gn4VGvkD5UpkVnVf3KsFyxwCMJzbU
9h8ZEXwkFRpMlvMR4Ai0BtOi6kKEzqSMpjHu0Oh1nfwYs+BCorslsd7woqFy
d2CSKmWFOLHCnpVWIbF0sX4JhSyvaU+AIKNZrBcjrvvI2pfMjsM5aHZyVHQX
4IIFKfRLev7g8P5hwgy9mZuSiBhjZ6Azsj0JPajWx81pE9488i4dBNmvOyhd
jUOj6ty3W8dPSTTyDzqNTkCa57Mf1oZINBut1/jMdh7/EoFMaM7z2d+fx88n
WqHdi0pmQWj8vsxJoIxc3TGnx4velsQYVBf7HHiRNtzNLbNKPOeuFyk3n9or
7SoTB52FS0tVcas2JHSU0I9TrZxtgKNm7EuwoI9iDIJKN9cxgd+ys/d2XSjJ
n7Plu1b9zCQpuKsOTsr3+WnCoU6YxVjsCfsuZKKxd0SWVeSh7zXlQLjDWtYC
OAfSOrfTeOVGIQR25Azud2h8FdQMgEiOYKB3p3NRuKZrfOf0k32L2TfrwPzH
thw1TmSQxeEGVKCCX/d9WmI2Yajcv8cHzsnIX+r5tElkkAFvmf1cQilkCFvy
ZBGyd83pBY1IU7egctczbbJa+FYJSggXnGg4BKbmp6pyoXa5CMdj+0ZgvjW2
pqj90oTtHPKHlHNjo7eb1GiAWxUnGqkVCHo3tRfEMLpUvqxIAdDNv3kq5JEZ
3rmTVxBFicZlsBTGl+3CKFE996U94vQxAJyptyWynoqocfMRIoCa4prm853/
xkV5gZKnhP/PYX9jCZ2G+zVVuERGPAtj/FggN0YAMdvSTNKOdlLK9/wNTv+z
fSogp9yxq6Y1GpoKh7K6M78DSVDjIPp45ok5fJFTjD//OcpbgzBoviX7pm3y
gIViD384EvDOGZy8Mc/IfiPBcBI7BIqeh03JhxAC8low3HvcqWl1CpnqcK2o
ZSA3UxrdjA1INyGE83Swp3n/tTx/wDkLFXKaJVAnzY0Vuo6uTZes0Unsc/M5
DxmwlzWTvuIVIO+5hJr1THWgxN2GeJm4SWPb0SvQKi8ltjEEhA5A+SW3a+Fg
L7pLsa4+DVCazoSELjE3jwTSZBhoRxleYO8zB6oaIFFTWJlUmjD+37TNKj6g
qw9yunwqSIwBpJ73ut3pL5Y+k0cUSfgu+NC86hmhW6Gv9XkYV87SBR3QfRFe
C2pJ3LNjlsKHxSdd4UEkta+zHQqEutje3VKWCaxf7FH2C45S72/IYZ8p3+Iz
F7qV4peu0CtMBnS4NiD2MlRF0/JSfivkQw01XOhp1g2NZWa0wwLIVlbHQugd
Bdof6FWCXrwk/o9HSbH0vWR7v8DUnBbnOgkEyql/Bc2mFON/DUbOYmWUfts1
tUg0iDCpjiNclby8LHq71NQBm184WHWtKlRbIAI8nkESvBokYKKji6sWMjql
CNte4PnaMHEx8PkPTDvW8GYXiZeEMYCuQZn3FKkzxXj7tmm/O6wLbn1E0XWG
h5mZlfm/ryH4XWGVh7LOyRtiglCF1Ekkzw0P8AwvI9VqmtzeviN8BUxc4WQe
aUeb+zgsn6DM1/ZmdcdMXTYGZnkpbKovRwi5bWfM6pdO4hKzTq++Q0UP6J3Y
ePRyivnzsVKDUVnExJIV18EgpjSL94Fl6u8TCDUBpr+u33FlolAc96VN31Br
DMtn4t9kcmBqJZX14u/baZv3h1O/3wkTYB1/RqKjEwm9uCzwFSAIZZSiQk2v
HNWl08v/PZDuvAAMWi3SMgnqQadKNnzNuoFVXP+0wdcSGdK72+K6rzLnjDDR
JQFbda3wTTV2DIQ8WBcbSjk3hpqiLpANWIkTnfULtoro66DwWnYmiaKsHbtS
58nKWXVMVtmzvvJMVNrf+5e06cYW/Zla4nl2Eabdg2jo6G64yjDrpMQOywgZ
eXSO5A6qqk4+k8LiNvdM6ulOiIbl/XrrECJ+fts4Rkb2hvs7DlbbWqCApJmI
yLbzfcO7zr4CsRi4OsQxx79BWgaIQVzeSmIDhTnzNd8fNzgHw0BHMmoW5kaH
uyTmY1tmSHnTparsf4BGQ7TeJA63RziVp1/ZruaEPnSFmX1us4UFi0G5aZeR
4YgsQebBOsnIpMBU5Ac8Qzo/BIuYCkx4T9/lnscAHUmSKOYFZf9fSoVmHyG0
kIGQD53M6oFb8/Yxxzb6AsP7f079NATdxkQw/q3uq1jq9D39g6j5Y211tKV0
nkPiLdMXLC+0IcfD8lBXywGWC9K1UhYmX9zFlDQPBfW0G3D2N63Yxywzm90F
GEjZemimECDuDZlsCvpvAR2OLw7fBIAC/tak06KgMBFRHChzu6vzOSzzgni9
JgFLLB8ivb2n4gAjWMcLRzAqoko+XgLixTJ15/efiAasY49KwYoeXn7ZxNw5
8wxh5iXacveXgu9Qhv9rcTlxHFbQGqeqHtwpOB5XWDMA1U5EaHeD+0sb1/Di
rzhBEe8i/RGeOWD1xDbCKnaNQrsgyWE1L35GeLNX5ghA1wI5LlECnpbXSaqw
qulpSLDfdYpvmzdZALw8Ahd7u+7fmxPugXDxqSHQuk7JzG6aHbDKuPde5g32
fu+xDpKBoFA39VrGUaaTV2Rl48Hbi9sGj2AZaBbt1dl4scot6KzGW3lSVD88
j30Kt9mijtJiO2gk+oLbRBXMoCeVQ6kZ3bDhG5EvpnShWjBgS4Zs9L6u8t5C
hxctmlkVtn7o8qiSvVJ7e5CxULWjed+haL3I0cLmPKZ8fVkPed9wkwuQ2EfU
TCaaHdIJpscCCNDWijZeJ0NtjzQyO8YvMVFlHmDh4TMC1i4mYR9qOJQa+qeR
f8fSXKDsPvVWk1YEWRjOWv9fLb9gwcZf0N3VjTRVTVZvjUQK6JmCUG/LPZBX
dSgxpt7YHmHN/q1vO5cPyENAkQhoy4ttwyLxuWOv79ndKVpAQxurC4kTQB9p
I0hV+ubcoVlg0SD44hJHn8J0tiWhdlcwGS7NlSASIT78RV5XZ0lduaBNrjUZ
S39TcfvKrq4OJyTgqN3WY3asA5pbbW5O4Z1wxPRPFrO6XF9gBqbwlOGh11OU
lkEFGA4jxdnqW0nz2C5oUwQnoy2vcjsf9ceha9Xx2g76EwehCNu2S6JHiHnh
pRGkQRAjfPVe4GlrU55IAv+COQy1eoGh5MlCOoxoZF1ZU+cdKul/wZSIEra8
l1PzGNVNbx9WQIHFKdmhH1KUDS1iVF64tUOUglu/DCnmdNNFLZ2Fxh0gUZow
J9HUJETpZsbTsoU4FHnk0BN6ajA6LgGlkOMQZywCd6rwguKmwGwDUa99VEdM
nd/kPguhwRGy62M6LZN+QX0sCku1kCUXA0KhMfVrwqvKfCGSPfnU6amcl4xs
RXEKFakpKK4rVR0hodqW6PzU33zTzzsehoqGaB99NpedGDVwAcw6CrQZ8o7U
3uS8/nB9U0I+srLLfOMY3kA0b1WZX8ZOmO7VGkMQduU9B6PAh0GvjHt77pOe
efhIgsdPySmXWwWpQGaHrXDcUokpSSQkMPJFDLayAK/6sEOZdLutw7pGdT6c
Xard05kUmzRu/TkDZQ9aQ7kyLqqIHlRt1Pmkwbz2fi9RxTBA7CTuhCi+qzP8
NkUiT4GnMEh2YN+XWxVBdi+VAexp9SR8BxWsq7JCLFwy3gEhe8TyclSqy1sY
cxOGTgEBNyKmmMOBQQSKmtOHa8PId6zt3M4rqe2DlS9k0JttaJSl0gSMxYE4
xrhcc+Gb36vpRPBuFJaJqLgaMYiR/0ILl6y8oJRkPlmRX+YtEudykn2Nr3gi
lCqe29WDB7GErskXZoysG1eZxTJujBbAZBbXN7WSXS7ufWH86jrgfKLfqP0D
wxyjD37qMHtXjkyrH9ePmh4PsusJvdoYeeOHVrc6f8PwXSEOCqrFwc1RTHUy
m2Asj6S2ZNnBNxDzx+MBMbXs+a52CXUELg5VrtW9Gu3ejx/UPuKF2ALfb0V9
jOhkP93+lPvl+xFtQC4WKsUeiG2fCwO2f9jQG7Fx+XMixFwOAkzb/4rpfueD
kkIXsx38t7re1gPZhw3oOLfRLOZMrdplSph9Ml5joQI37GETQOfPy2a0/bV5
8HwHFpxvXrw1oKkDDU24qzownHWPQIVjtPfmLaCDCMWUBgtQ4aZp74W31MH1
A/LajoyIqmGn90PLJfRlepYHJvUad7bVDkt85v0uvrVL6CzJJjS8hgOv8Nas
rwEYqHUbO68fWyvf52LqYH8X/KwBzDBqzIwZux2KsOngjdvBEiIfM+hedT99
oabmw00q/yjLDEQbdZq7UFxneKj2R/FsilJ2GtVX/EYqvdjTcJg5e2z3IqpN
Hp8vUisb3QMhtChma1XABetohwvztXZhPKniJsdnBm3t0WJu7xc+bIKPfdBP
XZLkI2dv6eyYus1H8SfqG8M6J3L3rjPon2fXYZTS553EBDhwkvyXMbGBtHLP
b6gOBt2AioJ2tylb8CvZoHDsAwBX09ql5VQ6b7VCsrqrM3Mthgkq73OD9JZ6
M5l3dfAa9+4SOWZma3r7O5tQg3W3hRjPb9az118XG4svO3Zr/+D/lCItyXww
dg13Hh10lczXEln5nuioK2gW2VXa40Bpnfvx2Z0f1p2pbC3ssHRgyo/V7T+S
cncw8kUNsqQCmhtY2HLEw2Y+QuVfz71MY1BmiEGy2xuPPdpHx9kFuy/d2TQv
9oB/Xufkl5lcCJBO6WTktb7/jaIhJcurBprX9oAnJFrwDP4zAWpXLbn4tAy5
sOA8+6y/nJXSUFGUBscqcYa+6g2H67BTJcBDWstLWO+IZ04buUHpLmFytw3u
/dhjpgzZiNNUEbW+4mca4rPKN6l4qyx7vgZIIQcuw0t+QwVYdjU1C+FIDAPB
AU3BaB7rYtvdgvjlWFxayIVsw0Ty+XSIB8WOHRbf3/oIWbOxptb92TaWrYc7
ZLdB4mEKtzp+mtfO8cy2yKae8QUWvecKBkkp+GmldGhOTMWh6F/wTZ+IQHKF
dIOYcyZhUJvRQurQoKtq3e/j4O1TLMvVUSzgLtFNH79GLehwUwgVBkr6qEVF
YLQZib3+67vSx7xHS9RYOkE3n3RjwjdOVTbxty8JpobGoVkQUkl3E2P20cxm
2kyLj2B+Qq6pGdJnjvZ8QleJ19OmJrBZdZBX3iGcoeVLvKCT05PtHR5FaXT9
YcuoSY6CKl4E4pGZJdRnuvf5Q4oMLNZYoR2aPxvmC3VrUof0ua8R0v/nUiGS
jgnug5J3CnfuayQk4gGhIiU5O/htiNhoRh2FIR++GVBJzPQiGiZhbbJYPYhV
9rTfSPbBdX0ix3aOOpfwGZ7eyCwV3w/Nw+4DAzzGz0K+PULY5KizoSOLxIuw
h2QwdY+eKIaNrNj4xfzWCM03Y9QMNc+ehSElnreCnwFwPY0cd0t/+cDliAdF
eLblVEzYLvXSZVYhy7l90Ku9llebKr6qXyPliza3gkfRwa/6w3t25IfPpi7D
SFJ0EMMNXXKxsV/KUM6ial6weRFF9ZvjzL0cPpNnJitI9WIXKpJ2xOSZfEur
WEQzGR+vr5VzXMS1aXbT4udcb3gqo8ti2HO1SrbqIoosYVcizGVDMYAGz6Io
yqa+DYHgHTJmxMm5mTt0hAC2jFqlcZt1U/fQpu+Q8Bd3u4dFEXisMB8dQvOM
19rLKjVIt7IAb5j6YcxvNDNKGFz3ezfaiuZfT4SbNb67ZYyhlC87Ud4Kg78y
0oGwOEftNaM/NEkO425XCRcFTglgxComotOwgT2PaJr4MO5ExGuYRjMjddAr
YibySo8V7iUBseuv7YNHTTTJbG6fuGwOJcqJbL14g2avDoq2oSz0zYbe+aPB
7cHeru1sIw0C56yiixfvhulVOO3QaPAIcU+gkyN2wiYFYJ5+DQvtYklfkStR
4Zc5dAPENduC7es4QPvcJLf70sdCxWeMd9uuBgC1JBmIFzhxfLW89vZHO5I7
Fno62DTutDt1ggHnCsSrjtpxpnOEJaSqOrAsHqBAz40hzFc3BVQBbsEWRmAK
GsWVB0eua2bQtOjBLpGIdMwbiaaTG+XwlyP6m0m2uOW0JYTgl8BeohVLy3p8
BT8xiVBeI9EUkW2nFUbx3zdl4rMsTO/JFFv/pIohPWNQzTmSFIltO3g3Xsl3
S/0aDKmJijyd9Nle/uQzNA3zfIsX4V0aMGEwX3FVD89qU0vkGXjb+3I9X997
rstvCvH6SzsHalLZkGbpDJHoqicAD9J1UZyg1E6jmsEpl6mx/Y4l6EBQHx0O
qbGQN1MC1a57CKAW4NObFS4vy/X2YAHBpAhoIRqLXtuWR3GA/6oq4JLxJWSS
jaStq9d97X++rMJoRLiCMWtZVqoMh8blk/CofzUvC/WtZFG7ime9txUE4iZX
Y29ZlAY8mHg8sewExM0+pPvM5dBgvfJ+2XYsFPZKrtJzcWkMsbe2zvnoFvpp
Q0KeuEWgKCMWGotplTRyoqztj0vVTOFLhDsT1yVVVPUEMlwviVCWvvK3Role
y8qSqULVsKos5K5mHr3eybG1+jPZTvyKTz7flQAO61Z2p857YrjAKmivgurZ
y+QziRs+xz5P9zWE4IfwyCr45OQf3D//4KgYDC+0VcCAXtAAKbpm+F6t9ait
ms3nGd1n5MyDo9sgq7OnI0OTKfSorPeihsISJPRT/VM2JkghG58Ox6/ZocXe
UCHPYfzICQJWDuHLT2lb+ycZyfMRZx4m0DuHlxZEe0eZ+O4TIY17+AO9YRtG
OCENJL2nj5FpDvz2QbvWg56vh0dEeeJcPL+vzDU3yVA4Tz164QgC9Y0hJTpq
1i+SQO9wZSBzB7JZ/6kWE998TXbxy5Gr+MTFySv8NsVqCvdgxuYSgDv/iUoA
213Viu7IBYAdCwWv3/oTGrxLmSGCsPYbf+SL9ETPqtXy73Uv9qZ7elXc5Y0i
8MwEpMCavGsV78zeQnf96Ime3zO78dTr6+8DuZz3txqCVIqPEiOQhxyK8a0K
D9d7MYZJvRsi9H3AaJAu19dGD4hTOTGzU8m9KrFiHLpBPdlZW5RVpU0mH/ka
66Tp386lbWi18N1kRp3FAxYvJy8938yslpVZXHysCqlbSBRw41ylsaOoUIWn
hVi817YsAdHKSQRjiisYz7CpbHJLB614TIAg3AHC0eP+9oufFHUZ1E4uJ9Xp
vzloPOInLHgFu/OEcpNJAh1UjPMabhWeeOaGEhrpHqRpwPYl+iDjnYWugnZo
QRheWz77yDCEw0wzu3w0sS7Vjm26R7fS73t5mXobZ7n3hSkPh/OgEvXRWmQU
PUq1d2+k15ac0jhRV7tfdBX5H+FoIW5zBHKDHyhNV0+r4YCTI+egcDEWiJPC
ale89f5dltdFXb7xik8Qi270e5SRWNTQ7rmk2wlAHJOg7GQjTKAlWUKI6Liz
OMZaHSyyyEmA8xFOSLR2Pj342Dthy7nNPS/dqU/+dJWXBZfGd5MDp4l8so1Q
/n78BRlcxZndNXq2hbv6QGq5hAachcJYEUTly6grkL+DeqrxueJUP0+g2r39
KGdx+uyr/rIeILUwc2SOWAeG/6QJYL0N03GTSnojfD3zop26Qg8KKjgvtX88
qWfFmHSP+GbF8B/8E5+VcgzxAeScmIP1UFfbt8ls+CwsnlggYZA99T7YPt6C
U+t6VMPGfqj87v9vK7+SNtIv+ge59HSXZX4SFnamGCOubPN8cFM9lCB6TwM/
c33px7wE+4Ch7G7O0AFAvffYjV2U/vLLbmyP33+L/u/QULEcqqslvJfs14Jm
2AKx/DrY7kZm0wIeTpUpnAY7a9ClMhz+XVnqUGzpAFZF0EGypa3cq6/bPx/0
uYhJr/FVUcxane1avs6Y8Kly6c3ih5VTzKPJRG3CtbDTJA/PtGS4DZIfsfh+
2FqE39umlFSwkKL5T8twwHxcDF5R5FO5AwqeJDS0W/9HCoK1pA8HYhErp5yZ
AUEDPhGgqMZPCK80T6RhD7kFCHtJJfdMnrZf29/KsCvEwXqibmkRUuikpf5t
EFNHYbqlcsMYc4zMFCVA116Bc6CJgTjl5hnMoYdaD2hBauSOMJIsTRjel2Uk
8KvDOH5M3XepkK0aEOCUBQYcQ1lazhOZdLugIGZTNGZ3MKTBCQnU6qf38U1k
Q0C5fVyXoQcvSZswnkvtjHIrOOo59VIc348h3KO22YS1Uqa40f3H3y7e7t1/
xMNP+KnWt7qN4Ry7Go84YXFdkXq9caLMnvRQYPzhy4JEamJIIxtl+j0mqGja
IOlZn73UPnm3SfQMfQTedqLs0/lcHk6cmdA4lLleGqfGzIEboagqX8QtSpuW
/6qWIZLqmdo/wSZLkLKZJjnCXaDPXRu3BQPtec7kZXDmXy6H6zXM33b4iZtz
OONXweWHQFVf4BUJ2LIZxIdY6ViWn2Jub+LNobKeNqpAO/YJ83mBbqRrzs16
JZM7p9DgA0KOYtebukeYMDz2XSUrJB1ouaKCRGFZaxbY90GhTAXeT2W+09dZ
JR8efc21wfSTYmhjMkq3n4Yhut/FX6ecGI6HFvCfwEBurlNAiLC8aaL7YA8c
4VZdNG9uwcq6I6DqLYBmwNaw/ojdFByIOj1QxYx6Agvr7lYZ4kfnGYo6sWgM
X2pN5daGh8wZNN4zzfQ5jGqBtWGCqXMgONbNNqgzdXfa6kkHfLrkkrmS2FoV
VE9dlOm4uQgA2Kd9YqCOb/tx4eJGdIhHfML81ZtW/8osyi0u1BtNJlq2/k+y
eeZOtK7knHlGrDdWR+IzIArDlds2WpvRBddpFI7257NZL+PSqoz6m2bkrJnJ
J8/JnLYPBDBWZ0ItbLvHt/UBuSlTfhvdnfoVjr7kJffmjyrsPWv6IdZsIE1U
a0Gsl1C7X07C2/6l9vClrBxrWdr6Ua3LZnBtkky9+sN29WjwBxUSfM7S4PDN
YKN+jt7PKmg9G4y5tC5ay2bbqzohntjdzbBjDoDoqeXZRnnq37RN5lbcheXN
ihCfCb/zzyqo29k+X0M2B1niip4WbNm8La3CQUnbBfkN4Y3CcbgyPtjDbWVq
jGVyZ9Vd4d+HIM4JPLO69NUMstz0eJ8r48+Ow99wCPZFCgzHrzFIF9Y4jzZQ
OxgVAfi38mVzmUkms+UGAC6b0e0q7wVZ/4dwvrjI25JmNb3uuzNGantfyuzA
OlB5eS2M+og+twUBijPT02P56Ln9rCrVsW8Uh3gccTy7ZdOvjtBrZ3yYCA8R
+MSTe5IKB86pw6/qyCN3Vkq38/GFQkUPbpURZkai3dLgdP9vlO/Sx8S1Cfki
BCqzSZYePl/VGSAH6wu8J6LEceVbVoSWufpIsG9vQOipca2M1OIXRs1fiEVi
NrIdd28TATC/ARUHvK42KgVLx7Ir+vdIs4OpN4A3rUmo0zQ60tyjm33VW+uT
k58lGeMo/8qhqyiwz7FaJrlHgqpMiRemGUStp87y1dqCIu8H2T5v7dzo9zKz
aS19e0sXc/zFTaCnBicMRGfYZElnnr+UZnhEz8ApyIbPXNIoVvdOzRyDuk+M
VU0hjkvVw5s0CswmsFlpOvcjrL1qyLaVgpEqxzuwiCq3UrPML26tkQRe4vaQ
og+JRe09QfX55jWhD81g4uVDb4E/Ojv7Aw4uEHbqE3iQgxQkOIFW0+PNEG7y
QJ4eH5Py7Rup6GbvPww57vcCSAdZuqL9bdWDLbxEHGFqpfb+VvdWtAo8bTY3
em9vFUDj3uD21P4cor2+mXZ5K9dJLK1A03HavyJBnrv+DqnF2IG8NLYv524Z
jaZKkBhc0tCySvaGePnzsquBzgNHRwOTVaRTM2TO6dykVhjzW6gw7DtwImj9
7ZFGDe+2qLxOGqG3mEDTdRjn2C6yyqwzza1wgry/+t9vLcgZzkCLXT6CWjEm
+Ga28DubgTlY7rImL4sZ3nQGFexphR6mW0sHVyLMtNWTD2grSc+9dgfrom7C
QJv+He21LH2Yj4FHso8HcVqxpYGpY+pQXybsUl5MFCPQI3WRf1V2AkLZ1y1N
ptlYPMOoLeGPyqN7/D4qWmEMFI0A+rAHFqlg54s3FK8R64SOtS4U6PJoY6dX
9Tr7HE6g/k8cd1+9JY1Aq2gfOa/7TTpgH7oza8Nm2clb9DN7KaojV07oLhB2
ci6b9YYwOY0gQehqpZQjt9uK7frqOlXy1sDo1wgZb0ne06ihl/CX433NkwaD
GzC40GXJnOmYGCD+XPBdx70rnnMkZtFVXji95ViZpscjyTEYEgHYwN70w3Rx
r048GFFS38vBjkVv0lFEKGGTp2vZSMMy6Y9fT+0cSZh2TBb2xv8ogx8QhheK
O9TLZ6Qs3hk5KpFkKs47lGwcbTNfQ4B4zBu1edNLBAJiiEuaNXevFNnW3Lvq
4qNuQ5YF6YZleJsD/OFBZgcPajfUNTi2Nx6bgO9+rkPHb/VCr5l6v3HjL0Uv
TxJZoMvSrL26zjiDwWWTpBMP9aY47TcKMJDRiBOkCs6jkclFCygFSHsnDgIP
By3nIcM1drpy8k/ccUTmSqz3OZbRuhLvfMPVbjRJlqxFHXQn8kHFRyG2saGC
9Xm7PfHcnrbE+vBgjw3SfZI7M19QCz9MgR5+0cMSw02jZP+xEids1jkn8tbb
wtLkw/d/m2JUjKPDa1nr/M1n/I2572nfawQkyDc676tYdZNEQZVCtpvgLl9Z
jge+CHd3JaRxpIVJKVLFSGJWmS0ib3xbmmq/AQC/xZ2L5D3uvSxS7fX6jqLX
6v+WTgQQs8qxRrfoefIGPS++4bY4Q3H5TjMU48jr7Awva+Il2zwJNYBnDWmC
3/R2YIqlFL30C9XNaNb64UP8UZvKo0TBsHyb28PawYVEIqiOvKlWWn9BGtOS
6T0X6cQxbrlbvB1gdtFmiMmbcQOSM1kg39W87cRYOBUFQNaOpsfbCY9RcvC1
Rk9HlEXEsbkl92KI/tWtp3+y2gLllcb87feZ6P4d2kSEtNViejHuAEje1b0s
ePBiA2fv28hu9uOj0WHKerEEN6G/FTSx7FJzRc+HS+MdgawQ6eEPjZgThFyZ
VaP+T2saLaew9w9UHSwaAZMkMT3twguCn2HT3RFaH5mKJwZsl2+ZgLmkGigb
jAEWr3ut9TmYJV9hTAfJCphnAJaFx6w/RCLwoS1sCmbh3VGFqG67VHJO7lZD
8kVkbubkclrRsgBB3hGTGaw4KVCusbMbw8ivgiA8KMJJQBY0/RBgcnDtmBFo
DefoneARO6SUaBqc8m5yayHDqfBYqAxoSDQLd4NwEuEWGLi8I5vYCEt32g3z
gPF+OlCS8FQT05e2ZoagmR6nvsrv8rV+z41uM8YZT0M/nqtP/Fr7dExKTvuk
MauU88TPwAOa9NF3DNG3NcwOoi0GvH0FBWPC1IW/rAWHbmNjWfm7ohQhMwNh
TEqAm/rbCDEjirFzsOr3l2D/mxNNaHxG00LzWfF2kmeNQjQF0z1OkXfM2Qc9
7Eqfy3axKuhR1FAD1Iasvnb1M7AycWwFp96xacJ9YGTVtpbPVRJq5VzkBFxo
AN+JAQ9GC5p7oNvU7Mh/tCVcwAlW/yBwAkzFymDnny0O4aAeM0UHfTVpUfCK
bp1W0xjeWzjgW82rB4vVsWQ5EWZvlfZKJ3aciWdLlLjtmJzEAIPO2L2S6Ol+
y8wyOjm8JtR1EfL5u1JgvGfgYCaWN7lo1TSrgWqlA+y/OGezs2WXOb0dwRyz
R9tyveT9I49LnCKyKOylriUJbG4aKld45SqvTA4YCNKOy2nFtnZQeeHvbwwp
iGHdA5UzEX1eyQHBTNHdBM6wmXORnDYnq6aWA88M7B3qfH2scwYlAWS3cBAC
VPH4qHicFbLGns4zCOa0o7ZLSvGT2eoXKA2tnZQHHAoQzKHsWhkCHeKjDGfU
P1GMwutquba+VDQOKbR/gkHCcbIHA/++YxZKeIiwfA+e6L+NkfChH48Gwoyn
sxwa6l20/iCBO9FnR83rAYHMA6IP62ltI2AtRQamODSrrnRBKV1rUc+JAX74
0sbNKhCzMuqN7UUxOKC8KyAWbLKCh/RsLDZessUKZ2/lY28fIubk7tcKN5t/
cEKM8N0jtOFRPesGDmBBCjrxCIoe8y95tdHDGdaW3WSh4obxZrjv0J1A6guP
C4YoofzbNYYuoUiQ957J2XKSqt/ZvjLO+donWtXM8z8vZ8U71rijmirRuy3o
ppFUcWWMPDGfkwaydRdhcGgUZXJDXnen50ZG9t11T70/XStCaUZ8NHl1DmoI
aZiaMYSNJhYmZexsjkfVuDVOiS3864r+A0b22ZQmK6AizNG5gNKtVB/nafUL
psNjmf/5Os5fcH4jbVnaSraE5uAMv5gWN5GruHWfUq5aPtqLVefmWpgRyPFT
ugJcjeSbFn2mLblLKfXlZVcd15kY5IEWF3B/4fpy1dCzk0gkZTyV5a8LdxQf
Esjtt6idkVmUF80eo4hzDz4wPlotPQg+XJAn3G06CMz2ihJNqNg/SNIXQyTU
cS8ce9LP6Vu1nrxP40p5iks0NZ80YCSuhSNSLeEZVBD5rcnpkc8qV/D+Nk7/
KoYfSnDvaRzV5EbkW4ng0GrY1DOb/oA6KZBgMKTLHwbvyGdVjlOKs9B8cyYY
++F8P1ITkq4sBksmdP8hkc1pP9mMxnAgSla9dShjNeCFrig6IuINoSR5ehxW
MQIE2ertvlBzfwiQ1gThPaS4+spPGAm5kvoj5FPqeOnxLc3cD8rzLYNqLzm3
Q2PgwE+IBgpD0E4gX8BbGV3DDgvbFgeTKbGYM/QpwACEZlZoYT6PE6Qi3psl
e5o8s1OcIo7cTm71L4lbSmy1M4OrNgNPWGGKJewV4I3NKvCljn0GvIt8t+BH
Z2tPBy/foUMi7VsGXMkD5vgSoSENkMJXSt0KdTqlVrm4k0WX4JgmtX9Gd6JJ
4LfDXzUNhzaMlVTc2RgjUlie2dyfkyH3rJkn5oIMGuhdx47fE85G6pQBZfvF
PgXmHIfoI4OBxFg6nMAPcGigTzEEDmSk1g9epE/Csv3yGowCKeZax2lhqubo
/kE0Ccl+JgybxsAizmfeDtSwbemrD2Alrte/DvzDvBwICJxk2bGejo3FkkWa
j9lbp0yO/oNaX1sgF601NzKgbx7ebsOeIdKWoQiFN/HqKmIs5iR4E3bpHaYp
KVg6X3KnZN40kmcIe50Ea/JvkrQglP6EThvdUHRukgnemWTZhIQv7OnFAIcp
sQ8CEMAsOTm3xOv+0A2E+HxmZMEmt01OV9+B82tH4a62trOySBNyJRxQPS3+
hhcngI7kv2vAR4yO66EUVCzgvfb0xma8uyV9FQmWJ78PXAc/6SxdR/EAhV7C
Oc/l8CtEp0NCKkewrqQQqCvsUkgrqyWlYNDOMNhpKQXBnV2mA0F+r0jqnd7m
/WvglBaPRSzEvXKoX6YSYYbgoOT+22LAHvAGxrtZkf0iF6WPlNoRDCfryN7S
mfMnjhZziF3SbCdAy9Ixd1FtNfToWJnJVhdSjXV+U1v3OjqfjcHT8bB+O6f7
wE+UO/JXuXqOtAsao0pHY8K53MT49r43CAgg64bqNhbsPuUVKo/kSVh7cO/W
pcDfE4G3I5U/SdvsSZHM+pcEr0F003Q5WUdiQEXg7FosUd4v971v4W59MBDI
ZHztVRrHh58cslBhBxkT+/aZ1fFW7J+oC5nFlTJK9uVmwreFMsOm4uO2h8oA
4toErLq/olOUkQjWjcTmT18j4yfQYes5XHvy1SjS5I/z1QGsEUAml8Lj3gjT
oBpISLXaUZtWIR8w00Be6yBzqZ8s4QJWuGJmJ52z4MCgjgb/BueeBJ+mDG4e
pG+KojI8MvwW9uVbft06jsqedXbuxmEDCC6v90bsTRiwwYrkmP4cTPPbo83P
S2VQqnUdA6xKCy5lgSbq2dJj8f8v8l3YR5sBh0RL8I8c4PFPU+CNEv7m3n/d
5XgkK++GHP/6eNXDXV2EJzzd3XIRqWKsI25JrZ9zh/YKVxH5ER7KA0f/Ati/
yFMM7fnz6EkT0RbAfrJArzRKNLo25h6GR6KblMrm03Ici16Haq3JFUkCY6dz
TPmpNP/u17ZC+VbqM2wyskDreYRbm+0cqwwbnLIEAHTbVgoxPjoyrd5X8hcP
OZOEjufJLAB0zMbJ39IRVbgo+sSlMEYje0z3QrY+SiFjaixiwkqmfufYipQ3
A9MMj6Campzi0hirOtFUKJ8nmw32nX5DXgIJiWHCwrcYG7ZhFZ1SqcyhIDDD
J8QJqaBNzAztXuBR6HQPfKtChYwzSA6itTaMlsrwBMaq+GMB/+4g8v9npswp
aEoOdPbgv0TG8l8+22BxyXsOWzrBCiMW2iz7RlikNS95UokecasgjOTbBgsl
V1z3rO/zJ7E7kSHtVzc85EojueS/SdRZHBg53+QiULYI4a65AexKtK+B7aVV
IbCRH9K9ga8irJV72yJQOb2Kqr418pjkVtAbhfudG3NGXm9sxUfs7ogHze3C
BbqRlNbapWg7q1YdxwKZyWmOyY1jYjVyfIRlVxAnzjiu/GwtbhoOVHgKgDR9
Qv9VwY2paCyShmgMaRAlSQbVFmj5ZzQdyNeEN+SSsEma88D7XqTFmZ4rCKXY
4EwDNVMD0g5Du1zxyXMFIsBSwunYccuuKp1j5d+JWXH+3mk92KDEtXumu8Oi
J8GCQ2+Y7zpytzr6ft8zkJ6lSE/d1NGzG6qBpL67fX+HBGYgrpdgh6h9ikPW
bQqeiPyElradT6HA6SAl6hFkOYJyDk5cBNBOqOd7uTcHMevf1tlEnjt0Yqi+
DovcsyxdqwpXcsAr0bffwIdpqfyEXsGpQmV9+UVLB2w2TlPfxU0SIf3nf/XY
9H/YqUXY/0kPbCMfqKbjrSn2EzgMKJ9MwEcOGv4s3tUYLdQfcQAhsYwObzmh
lOr2twy5kKOQeWlMdZCHtlfAaQV8h8F7oR8Tqxgl70JWjWO5B5DXoyetxjjm
orcghQIhiA1GRgLSUmnbAYrHEXa0FHFGwVJAix1nee0YxfCWAa3IDpjMEsi3
oGUAQaUVlgFG2ZCdYimJqUTkYxNjjCpRaxaWS0JG89WCgiuWTK74xLFy9dL9
pwfqerpIdymWdFytMj+n1b91dsujr+d1B+yJCZ9OBxowUmU4VygvoWJ/Wcqp
BjdKy9b1etb2k6ZgdVgPkenYdQlQujXv56rsmdiEZmiYV8QehsQbbUkeC1DB
UDmiBTl5akLNEc9f6cWGucBi7s45e3rlXuNhh8fFQ4eST2tUvZc2Qif7iwOu
3yOYXVSbLWJv2MS0svpMUG4AC0AgjTk5Y6PYL9J9Ct1Bea1fbI90Lm7usVJo
M6Ot4xVMyTiqybqL/LkedW/cb0izPg6EkwU/3M+cTxdQRvuEM/uTcemYtD3g
8Uq38WEZOYySOBetpzrCKHI/FAeHCsxEnG9/jpxU+jQhSFmdflDboi3BDsn5
JWF6+d0ZUGMH3KONPNg7rNXcCGwOGqMKKRk5+HdyfPiniyPvBPGXBGRsKwDq
ToHmuqcw0C32L9A4oR3UNJwyZUFXUa4Teye46r0FSbeB7rNCdyKJirzq43YS
Bv9ljCSXekiVSDj+A3X4Vek4oxy8qugrLZrFN2B2N3rIx6vrg5V7Z3651xgY
QMPYILN6Z4f9aPPVeVpfw9n7kEWUBQNYsKGzvmYQ7ttfnAMeUPP6xfGYQW/u
00gu4twvTv/AJI3mj2RJCHs3w1moeWc+h0EkQi7DPglZ3rOZrd44FmNqeRzW
grwFIee6qycLDRinPTRJw/6cqID+nlAZDmPDXTdp6u5UCBhU6DzazGlPKd+r
yZ54DdetnmpCjYmh7vg7Srp4haij0dQLMqmtCaq/UgiK48Va9PV/x0K4G967
BpERTO24GLyYAlRXi9+iV2G0NfMWpQJdfYENM8z/RpY6/rvEwOMj0hEqskbK
mEdvWrn+uQYqDvQwbBgykYxECpV0sds2TDECvjGRMMnBxcs+88DuWxBdMfFB
DGB2RZVEE0g8tea0zlIXDNS96gnHWv5kRozO3BMtV6y1Djqi+1tnq1dJM/ze
jeYh5D5ABamVZiWteyVXjtEMZCzqj/zdZ/NNWHM2oayp5rK2E07kJyekL+R5
Ni9ldBv4vdpkbQJPG1JrvxGJn845hPA0cDEVfQp8PyyDeEpHuYfyMy1bp2wI
EUa3JNo9SQLCuOngSVBqnK2bKm4/KdvJUtDXzcMFdxbNuVswyYX1IsoAvd25
7TZ9JGVijC+RFbXvN5L+L3UVKheLD01Mj6LaiMBAXzDSbatzAfrkgQRFxowS
WDkJn6xTsIPDQSYZ3yQxNq3Cat7zQfvd4calE89xa4ONxlHfnsKBn0sK6CRJ
31rHKY6AOv920xBt2jXtPbfLsgJTkqWsPkIbSU/RWInjAgF9v2ad2flUH0hv
XE/0EQkBY946KopFRijU08mQ0Lr/n357ZetCzB+gr40iKjpBALM4FyO+Nt5t
VeYwoQG/jW2qE2mfqAsAYmrKDIqSdBa9fFKwVRENSGDterW+zr4e2AkkbVQt
/VVuozdoKnzt3stg7lIMV4PRjRWHPg5Z0XT1wwz3I7LPCxVZ7BDONgf1AUwu
Gw3yhnC8SYAu+O8wSOz1T074UeEX2d3P6BpwIHO+fRBgSsofQLq/eOblnLF5
iPwDrtNbxnjRlElPdXHn+sb/+h3l9cN6ksuwS48uEufO34Kg+C9yZKRmyE8W
DR/lKGbX+SNy5x6ADlF8rdFADMOJYxLkJfbaN8xZ1W25hSCsq16CAGU6t0dX
RN42PosRl09bqADtKFXJM0hrYAZkqIAIY0EvT8WIfsCKBHHqkjwf1YaSgczj
Iwy3EPE+dJtMfCrBOmiV/eSmIpw5tVOJ5ziD5+Eb8q4m/o/OLw3wHFnhu+Gy
BAYCuUJJ0wp+D9kbw3vuypG+RYmN9jKfauf3I6PpYGzvcGM0RHZyb8yHQmRZ
rO65/k6sta7s8/wkdqt7tHaAy6Rnne5PwanCL3NQoURzenO2OhDeuQJFrNtm
QJsER+w+lw4rsiL/Ry/CKWspR0GKJ+v5Akkt6jM/VSyG/5J/+mv0mOWJnggZ
C3/oc5ZE0X49+hu5/Aanw2MuE1KcqBAordK7dy5huCNZwR3SNw80RyHH3HOt
Db7xqtthiKXEl1gbDXL+OON6Nnvob+Wm/JuWiUNj+/KnwOOLR6uQprt8rQuN
NBy9BO9ao6qW18ayVbKwWpQ0x1OQozf4Rr2iYTQKDqgtCiMORLfbAsiC4N4S
z9xUomiXF6aJNbgcM8SHYmNOgrALBpV5Iu7wxlXHptoea2lV2Ca+6nCWauKy
fd62S/5DMYLb/GEMm7rHqxAGKZo/YHKL8sG1LwYRuQkqWKJhRnih/N21gX+p
5TJka+h0yzx2C7hD7pSDU0WlFKaRcebeHUHbjAE0l4f0us46rhF+JgAhoTAm
uVQn4He5+A8tnqVuuVYy0NQVzinEYrQjVvbJml0h9G+nOzzS5BNoq1DOdS7f
w6tgYbVmxMK+MmE21npCv0fqD3Esu1hPgWvZaAZpqW+1ykRvk7cvQLeTXPPX
Kj4i3Y63Hs7FGXiNnOGk15gNDFytKQdiXEMWWxIiTEjSr2yyFGTeT+Ltlopb
06RB/tfSYd5QMbn82xp7Kgkjh6mtpdOgwMI9VJg0kmOxTIOr7RnTIv3aX1Kc
oKNsX17+RyzjdH7i/XAB11poCFKBFCI4BTDDdUUWc10jqkBXBZClclvY42Tf
zv9drRm1Q7c35U6ujCb/Jrl5noK9MjzB1lxHgBOLd0PWd8bW5SdIg/QtjwS4
KShdE6FcZ7oLFR0qBVxr4fx2TFetvagT/sMdw/3kKKF9K6XHZnR7vl6tXVAb
4k8tvuo/g/w71Pg6x/d2bo6kb5N6K2h536HenTG79VVEYtfimcNVV5jYyBIl
CdmOvPbRH7mpyjyy5NOKIzGtoDYNPqKw81DqGsltwkKvKUYtA1/iWLXQvhec
EIsF8vbrQpMspGyUAEi0XblDHREcOXEiumiNTcDawvuxQloP/KInnv+j4yta
iodamRSF/zv8Igu+XLAhdliQS3iYB8vSIhrIVqXVRO7dD8JJRfYxQVc/pX6f
q6SRwsoWUagyFNutGkbw0oaMjbFql9Vo5OMpWGTRLluJIdTT2M8ttVjuAOqS
NYwiC5R82stYrJp8e4o/GJsEBWP4o8nNhQYWGb4ZTijjKgpSMh5Nj0pkYRib
9F4pwJ9qDetTRN98z/vva1zZFvs8gkO/Rc0oKjd59Rk5AUVXYlYrVtqhhaxW
lfG7G7ailFgrjEeeFFdgglwvICk8QBggz4M3FTYOHvVHdKDRt3vssziQ/r36
6NVTX3oTk93JaP/2ykNT9hID4r5D99tVGPYN2S0PwmZGc7e5ucZ7IgJHwrhf
8gTymIJK+HWbfoo78zpfNg1gjH1JA0RcBMXoxHU35oWefSp0BRfF/RjOkKLR
dnQlZifiF0ZMGGp0+Y2KG0f/t6ndW6nMV0/5HR5xSLLgplizwMzbT2wGtoEH
uKA/JcZQNUoDBinFLrtNAs41HPbi7O8NghN65bSS8haWYbpGtbdvieIuspSe
WmwMF91ckqPAfn5dbOeP7UB/SKy3ZF7fNehjNuGSDztlTSpfjXE8PYLTFpUJ
Y0impV5ZnOh482JAd7uCempLNB9lSOcmO339+aTzwnznQt/2Yz5j1MsTO2Qf
n0QaBugzAg8NuhheWvKXGk/f8z8svpAz5LzUrj/Rl0OeX9mIpWasVjBn6Up2
hynB922x5Gtm1LG4Z8DQPxvEHSFBU1YN0v+/a9cRdzkdyNfL15tSJ0o1caZe
jIDzc4IytOWX76Fr6iQ7Vt4pxquJ+qSu0T682zb0HYpjy5cKX4lvf6fDir1T
TgGnv6RSXqsjLB1VGZfdvbLuN1piCIzqQeFmT22WsEhEDawkA4dDL+NX8lfB
B1OQs+2pN6TPYrHm9n6N/W0Co7CYvuigZUF/xF78ACXWYnLpZL3kzq6yf8on
k5G+Y+/2REAhjW3JKB0NMMFcY6yh3/RmxcXpZ9EQN873be1I7WoCIkSjAZzD
LqhjyO3WpoOhiEUogQ4T/hSG/T+Qck2n9lZyotb5IBENHvhldczOBf3P1fZK
NfNawuq+7toI0jC9WHzcAH+fC8EIz2s+tZCheQ3ulAgiPpGVZBN3VjG53nLs
MaXa0LPRBf070Ndcs7GGOVth5PvVBPlefb3cFNoM1Wtzmy3kYVSoWA6kTvFa
y7wD2Xkw8tCHZDodzSuoVlBqplH/7XZLsWkzMDc5ab8HOx22vk1r0tr6SI79
4I+7TbTeuL5BTCrcA2FGmXeudxr2QBkBc+vYEJv2AZrVIQeo36nzgGumbMnZ
lkZh7oX1PHi+3CCdLymzlVZhEJMRBxc4KS0AvgBPkHKCKtY+CbhrWo3iCWYO
pohPnmCodw18L0fQBtwFkHLSBjl8+H01Yo+EBcbWdnYXSHu8j5HnVcV79dFb
0Rf8jB4EQbpAZXPojmhty2f6G4EKi4/rioep2rtFD+3/dR3J3JaS/Raq1UKs
LH3hunTiLIy8cMNnCg+g0Pocl/a/yfg9ksn0ZL+xteL+F7WtQ26hFOdJ0SIF
ikaJ3XPrW8bSBBR9TOtX5zS3erzG4HfQHGQnbSQF4Yt3OxBSTHzF0uZhYKLL
RiViXuk9Yl6uyVPxgynf+RZq5EweEI2QY5xYNcBa0c5R1KIpTl5nlwv+r0IR
RBIz0O9Wd7ywLWHklCJ26qR8jvQ3eOichyJklaXs7x+SCGa6dImVv6AT2hM2
lMHFK1htUUJVWfDOKv3E3tmCro5JalADbmYCJteFzNTNeCCwloreLfU7tpWl
F+uFJh9RqE/PpGf4fkM3MXaG6wpeC752Sp1nNw7eWEse14selLWK8MbcfY40
j0BykDOOkou/Ji806sUxLSrkfEZMa4JpxwMiAdp9+rI/tmPhBPBpllNqy1eA
tKtwoDRxKZ6Myccj7UUKJ8D8jnROucTJsyOohJKfeogZw0uBH0HXq5lszk8l
byQUWyQ32Zq8f3wB2kj+38fe1Bb17wqgD8HD2Z9Ukwl5RifGh7hrYS7ySZwA
QXnqhQSoplDnzX9PMCRPypcyyBq4L5nL3XYRHTtlnHQYkvCz2A5fg66E6mRt
Vn/aRSipJCErclH9v7JYOzkIcw8xzvfmUPtGnFwG83Izps/QENVVg4/opxED
iYS8o66QsNDcdkJxP/6yefjvCcixjpzKemju4Xf1xk1swjMTzvCLRiclqSdK
qWeNrzoLsDhEI/yddIsyRcs1Sftuhrqt2UkNqJJxeRKBKwDXba8xhEdLrcfE
laTvaPnhsBkoyfsoYdDZkWviWeU20auxHrb59BZw0sc0Fh9Mw2IxchRD1eeb
5lIGt6BD8uznKPiiinuX1yhzS76dHjWs0o+/QOaFXH0UXFOnwZLpbTISrun7
UR7lJpaUwHVh9uMx44J1JNujxOGQ7ovpG7Zk1f6+2laMF2NfQKTfJ8/6uZ35
4NZ83JJDYdriTQY2be7+Uvgtj3ie1sbbSKFRMFbZLtHra36A2/LfvBEDUF2a
VydycRYRlet+r5oi0JDT6PQp/z/hsjGY0r+Eo+Loci7AyfKT614JWQwJ8UMe
wlOHOMUGsTWKlmyFwshm4/YY1Pa+RvwEsYPfCOlFS6MmPuBCwxe7r1vA5DGs
7byPa53aXxZvghANkZbll4hGwi2q1NvOswBJWzkWp35IonvUzH8Rf+YN7zj3
srpoFFDIdzZHPgtnQwrEbxz0zotO0yTp4oISJO1Fk92prxu8GzSq4Tm5LzuQ
FrYU9bmhYNHbLdF66e/Xx6k20MtgSxfx1whg/ABLnheDrFZqocZrb1fvfanI
v4gLqnq7cMseQpcYfV/tSmnS5VPvcNKIerCkLpjozLIUrDGmaTCxlx9InGke
YPkmxSW2C/KBRDHsYRpTvfsXBQPObw5ZAgXTZoHiaqyZyMcYUzLdV9dJQj0y
jBOGoPSmmS6+iJ0t9OfpP+Ra5orSomKIH2c2WM13MnqVjtQ1ExeVWlPsf1E+
1dIt6OAb8Vos2nkibyfdIEVD9MgHcCRD1YNrIkrwgnPark3KFcBWF07f3Zv9
DAjWiAXaX38JK1D6QCTizvDqMPhQhKufyoJkY8Vk9fwKvCCCjlbXkJBj3IgP
y2YlT/eBLibUF1Neo2KPa0r4haCbPZSn8IZPjaAAoA9HbuodilEBeoMqV8TZ
UiRWpN7sT0a46ku83Deb3nDObhXdEQg3yFHbFm4vDsb78YN/JOWkJ16GB21k
Q4WuraX9wSSaxBGtJ5hZgqodXV6XKAGtoaCB3HbEXa/ysfOmapgPZp0+5+8a
SofnxXBow3EgsNfjs0UGnA1rjh3MRPDGpyft42eeDPyC7LhPV26c5rjNSAKA
Sn8cozvmCJxTD9CvBTnqMidNiAzFdvb1oQXnu6NUB4zmHnpPud2/0wbPFTdU
hVbZjEqXF/Q2lij+hMxzQrdWwmmFFjEdPPnPbsFzOl72/H9+l8BGtIStpnzN
TDUuGdDB4iA0c6ZW6eHtWWA+NECB2sua9apKxtKNMhmv+Uww76mo/GnrAJQa
Twy7/YWurxbexpm0XNg+7oh+ygfmKqQGojGpMBoMBv3skHQTC61RdOhrq1uA
9RldkPVQYPS1RcuGuGNcMeneL72n+GmVY8cEpjitT1KwEobR2QlrhsLUVIk4
fF1PUdbGBtTBMNyGYEj8+sggcABZf6N6KN3gdvr4iohPJKToZRreTiIPwe46
4g2upwdZz8ofyX9Cd8mtT8NzvqyjznM3DhRp3KVZN109DczYd+q09OLl6WQK
4tDg+onaUIF2WFjdGQPiLfjNeqSXxTGDkW9Jf6aOzzB04MSjM3sIdSxbBlIo
ihN0ZEAQmUFYNbzdOpQfCG6IpB8m8pguermkP+wEpi3R46eRrZ58DHD61PAl
ks0X2w8GiUCudeyyJDlB8MGyZsJD5EIwAZlQGnC/o8B+iymKP74vKElQE5uB
N5MKtnGuUJ4SnpULyb0K5rW4iGYwlJVLP6NtYeKq4/r1fFdEQnOXd8MGxKZ3
ecPi5ATJCaogPCQFima7Zfba016D3YBQBaryE6GPHMEivSSk1EgzvblXz3oD
kgfISJWfAzV58bZOpzdXxx+190aodMoELPlJ8i0fSLoyzZAqy1LpADsX8mBp
tsVNebY40XfGHuVmKe4zaYyhe4fK30ezIz7eTcpxX4wZ7hvNgrdzjdOW7m4O
HRJajNWv5s6XWiP21YX42nN6PRjfHXFLxTNUULierRrklWjA3QKuvn7CTWCp
Hc1nRAjGm4JetLC2TB2wZMsbgBgPIcMR/7Mfh5zUrTCYhfxojYmeLz4Zvo3H
vvMeDfMqFCO9q8OzecleUhi1k2O7h4EJzaf5yyfK2junoiqqZbA9N3ciR6p1
Eh9eF+HynaFmZOdwvs4EsSy+j2n0hdWR6Q45Qymx1UlMT/TnJANrnK+Pcp2B
aySYNytjMZyB94jZou//5Mr+6VX64PhATb4/duCPA7zeDjeVCYqVf4GkEvU/
wGa23p7k0wBO/WlrfV+QPeaSnxKv1Sh8cdpGjyqDKyDxU2zPd+SDCXXWSaaR
G8hH/XyKjP2Ohx1uzw2FdgZbJ+g5CO4ti0qPRynMDXa1iInjhsOOn+lNofD8
22t0D0Um8Im5cRGDn1uj9CdG9kCL3kPh5APiwmLxL7KZ+dq7kmfTaEou9iQq
t/ZkOjVorSMdmh/45V6gaScT2nlQmEpRsiHxEOMTs/6cO0AK/yNYZouE2xWq
Un5WQ9tvzKK3bHKfvHrzHRnlXS/w5gBB+TmNFZbmQh1AndVagCh0gUK4G5l+
tQ1jwWpxlkskLfNAFAUL6klRSfogqnQueDUGdnyiCM+nw2WQT0s7p6aAi2IU
Gi7VdYJH12v4/h5b03i/fOuI1EP0LctgG4ug0/Jdeo9Dao5fxxPnAUXIfNUz
96HlOHi2VuGtPHAKpHo9eqWVKa6pRXelTKk/fMpWFfUN62W2u80EtaweAxIl
2EoEnXUiJGhZ23cTQd0wRECQW8Xxj/5wcHv9vmxgCOYzh9bbCoV+MPCtp3PV
NSD1hpAzPg1WwDnQka5p/h2MS78Itwg6kB/KE2/f6d8SfF448Y1b/uffjsPZ
oUrw7M8v5CiYZTsUY+oZJLuqNv1Rh2YBkfDQXQ0yBCrABFy0QNsKXN+ErhQE
ikeEgQ0zKFd2qevW2/Y1YTKL2SmhX5ZXQopP+VROSfMBIrsBc/3YM5+dSI6c
nYHWCxu3KXfTXjcQRSXqNCEafnLdPSRlk0Yvxsedr0hYb4VvV/EYGiqLJhIa
t2Yhw8A3DbvS0B6BSjuP4jXE5vx0mohBwybIZ7cE0N1TjNlGjNqnELJY+BBk
z+YWTks+bk/gng/I5J64j3bSXitRqbam4lbWgx8j1vWsxDVSc1HUOMym9TwI
7oCLyi91cTSz0gGSM+S6LscltKB6j/sPNVz82i4KSS9mR2gLWC9PZJlBUFzC
Ei9T0AA5ZDCIyb+xZItSBRhMAAmhA7J3oeNafMp0zwtQCE4iogZN1iUfASQF
jW1/aGF0mqqa/JPmyAmVvOEyNgWDTTqZfOkoUUm0n7lVsukve+vcEZ7xtBTx
M0dTXqCuVtQZDjuh4edBV2lnnte7eXv4b0jY7YCNMmoNzlGyyOxv5YYFdw1e
q57RUl5YoUjHtjEQjnRzXADWVCu3pKB/RsdB2FIQb7USUS8qSMd2rR9kr5gQ
2pBwjI511GqbFtQZmWR4qwWVEMKS/vtt8YhrJg2LdOQ4AD++DtpnRFpb1zbZ
6oTd2N3D2Q/pflLEA88MyLGm1wvW3H+WliR+3DYtU3UcYyY6XUDux1YkfMqJ
xOGZIiiTMkCgXwzHmys9rNtRKaoVhGlyr9KJ9+NW6u8wi6Ze55HO8YmugR4I
EQvTSAVOqczw1h7LEnKrhNBxCOwZUq2JD4kiVwswGjZ+JCkne68BzxMaI1TT
Xemm5uyqT++E1tbqbLlUwLGXelsXaMZbsWrENBnVLTLz3tg9IGu1YEEAwbEb
/o0MSlvcveGyyfoF8+H9CRlv4l1e0LhuUc6JpjkkycipQqbAImrxRShFm+r+
uxQFP3UQi3lsSftbSTCcXd/up2Z48JcswOGGt8ZVLZzM+29nk/AbAy7KVrXt
vaUoo9aL4Aa0Ymqi9k6dx7z6aUWW1SFGLhzze0hTSa/OfS1bfGeRuK90fB9S
DZZvdEyWDRpJiL07J3eY2WxEEij9vvg+CIoNAQRmYhHEJ9B+dfav2nkOtrkm
/776hcobQQBcKVrcKYbtccAbw/LNO28AS6G1tz+zliBPTN3Y+ktJJY0uxDLp
2/SFzgIy1nvjbDF4Dg71x9uTO8TytOSm4goUAjD9DpqcwKCTLm8T3aaCqCCs
jF4BCmOmWdXzoZLZ9rTQm5CGy7e6+ygUl4cjnKJEAsAfdG8fL+XJ2vfHkFwc
i630723vNlEjHggYdhMiQ9hf5a75XoiBcEJO/VTpkaIze4sGH7zU+JXEBce5
Ym65dN74wpebkmjiv7WmQeBLucmH54xbuMvv5aKDHS2fTT8fV+IwZSrbMYJc
IPzgV0/8L36ljLEJzzYx5NaMj+lEb8pZ3usv6Ev/A7qH7+4NXV46Znnx2cwZ
/nr4Yxw3CwuenGapHeUqIIXFEmWCiOmghK4tkDHnTJdlBnQhQsl57UtksdBR
PqrmHERZ70h/Y/mgTA8wSaSTyg+je4QZX5s0xhYHhL3VBCNMoC6WE4CjADnO
4Tt2UYT5dV6jFa8cn22um+Tci5KSOneIukGOX/pyjotp5mA2hheyXxTnRIUa
QAxgdcBv535mLtItAv7CX+Q3H5h0LqPxKBT1k0tUm698E/dt1Uae0sL2IEEj
X5ypFbIX7maPPgd8P54Dx646a59RVE39CtaigEQYd4PPuv8xulZa/0TtEVTb
fsTLgKq8KAiJQtLKlSrINpb0ZMKXmKfRHWcf/e7t+HIhUu3RgVf89Lpp8V1m
A6B91AyZ/i/qmGkA4ugDP0VOzSgzVygTIBRu9WXAOqlZUO0gdPf0C/DhrL3I
sQkg3GFyYjFXqah3D3nBgjMl3etLUlbGF04D3EiuKETdSOvXInpChxek1Wt9
OPyolnz2zu+9T/kBIVs97hBfYjudohEskr7RBuG/927wdWQ1dTh65Y7iqnXI
SCjJtqbub2QmpTHedvxbpeDoGDsf5f2t3NIFDyaSNweyiKdH6suJJ1+zBlP/
f3Gi4KJn0XGyJO/m58whUo9PsuYpzU1C3+YU+Y3CubXo/pxBMRyzv2quyiSQ
sgwyhH6qwGgX/EB0JZDYEq33A6iAcQM330KW3+HQ/9Fs2yBktHsO5XmEi+C2
+8Yu7oOgwvsQm/YhnIxqeLbP6EBNz1ZAPy5hv3JjqsfE+7720Lop87MW/4tn
0dC1bxPQpfG5tcUsfW0tYai08OV30YywsreJmLni2NVjBpvyelDR2iUYfJg/
yBiW598MinIbMm+MlpecYOdKxnJ2VKTm12omquYEOMthfVepzs8Oc1yE6V0P
KnQiW4ESu5Oupzl/9a4sA4FTGnPApKEP0cR6jmklbRdW6+pkpSHmH03VfWR6
/SVRqcPOqIeqBtYKbaRMOr6Ixqebj/h1o7Bu70fFWOhylF0YLno5/O2WBkqA
Ojq9lo46uZaPSjdS3Bnsm3tmaKrF3X6aiVkm5eKtq0/p6+mO/vi5US9Rujkt
H6oPD8mp7JQyAb3+B1P2s4x6X5+hqmgxaJKW5qg9a7/C8RRWTLSn4Ab4Zrri
CBSB5KR41lBAD/fwdMFyeYqnXkHo9bhGlM3cQ4XpuDelG5ZI2Xnojugw0kKc
IIbBwhCFlhr3/zWv2xqg9hvm/VfIakyRVwHyBovvLP7/YRNt9JWphB4mirww
ttJAWjeMPToNLrEHPUkBvmbx8uuNWzS36aLgVm1WEV1fhqUCKSy4EkMDbdqM
v19mSTd5/78o2ltLbJ8LjdMOGJvT60Gtwyrq1BHjaFbv4MOQY4CRQGr6sA9Q
lXBouJbylxOyo0NKnhypoT53AbDcrFASXhrt4SnJqfF5KtW562fONzXuzcSZ
Cz0/rjgAzUUYsMN2z1/UUO6dCPMEYs+q6jjuIyL1Vz7Ipi3JW4eigzXEce9K
DqRYIB1jOdjIlUuZnT8Z3MV8E4m7goUURp8xQleBcLi+XKUyp9gpJAArT7YK
X722iFANd8dMgoGa3L79sfDi0WaYM5TERQArCVve/Am/cTAEwJ1JilQZxiAa
CXUrzNgTwpby9B6/D80ZOTVBIwXOvlZhRDgh7/xhAofmwVnXsXurElBSpDGN
eGapTTOpJYR/YlsGADUxLVlGZkHC2gBl3L6TJw3k/CTP/drwkGHcBIRB2NLy
tBtdWy65qlhjhxWMhcr0faZevV5ROzQi3MMunNZoaY7oAVkbxBIIvRv+7MzN
F/I3o4vqWxMrkC7QO15o07XbZQ7eVNuCLeyA89C0kZwTTzawQIkuHfwWusuM
ejjajCpEmQCXjk78C53wq3RN9xR0PnqfuGvv8C54E81EKahuCEiKgC42jLFg
6asqYTHRyhVe8raCPOBTQG7WnOjEhQQBaO7Wy0mNNBx1CanZ9qS6Jwp7GwIc
6pr9RZhJDSQ8cQqJSNJ1FVOES6lgIMVsSR6dZk2ecPTIQB+Z4RCgna62ewSI
GxwCG4yNviMPRoXwN4u9Xeas3kqQrj5BwNSJc/mNtEz2VzR177oteHRtKSVl
IXAKvvxUFyng/8gev/WoLm6SGa7Y7/B/FAXJKFrvTg3dgojPrXf8SoXK0n3O
U0O/xhg1PvO3TGp+MG5TyKhiu36Iuj8rfvrpNQq2Pr/tfe51ZHXpvv3sJeti
D42yiYw6fe0ZPabcGkT9X9tD3k/lzo2cVYvQfNQab0AHP00l4Kz6Kr/PlN8+
WM5dJB3uGVUK4l+T7uwIHdQI/L1k4o40U1hu616fpNYvdScmEe1BfbRyMvjy
ULS8k+fbsU6jOnMfyConh/ZlbyJJGEo4dORli6PO/ZNyQrdGkquIQ/Gof+0B
G8R6CsJzLHB8gL8gjl+wqpoKetUUbvtETi5u6VeNBkL6utraJk06EumD7jcl
GLUp+/PrjmbYmU+/lg70AQOGq9N0wkC9aKZjGclRomTt/cc9eGSLfQKdOrbL
m7DwzZVIP1y42N93AJizW7C5FprwCVWYi4zHqKdUvqmI7WdK2ekcfcWl7cLY
XxYxp3gfauW1+sjFquQWPmZBRQZW03NWKYS0Y9kR59oNMoa88xZbOjIOIzMW
XAMVq9/65jZubf+c+OzylMcCQoXuG0n+JJ/yJrCHGyTW4BfM0RqMnJl84K53
wCkTLhJh3rx1rsOmx1wINDUW1xVW+HxzYoFLNSfbpd3j4MyjIZtBbNz5gYVz
93oXw16fhJ8lA57Th0+9QbAe3rcAPu3jbVRfqLOAt09nuMAFBYqq5BznJDnz
r3KCZMl/l0KNKvd0QZzTQg+7st8dEXLX+DcbXe5g1ySNld/JRonC7omNFkUh
5y9Vn9WA7K7Ce3TjrXKmOFO8VQ/DdBOEexOOZQaWK03z3K1iJiyTqQqzwJMh
Rp9K8Xqh9LQWN79DpWSm+toBLckSSmCxU49qWcFL277kMY37LaCie6mBf9fy
DW+Ba4co6aW1w2OovuAHtCFyJCt/cexdnGVTVO6yRL2w+HWn7fau/zollWgW
mPvBzL+0GZzj4YTHdIyxIctGSTsEzyWjmZlJFI0SgOHThW888z6dR1GkZY6t
EsZ4mgHR9fusviOBZZtEUH8hqwKE4zyrtUcJC1uhh814us7FkPTrA7Llusht
hG6f98ohjZfPREC+eJimmr9xpktT+LoSUIliCyRLy9/8+3OgOeAPJ6GS+jy7
ykQq/zt0RNKQTUOX5zKTA+pzLWoFfq/XTSgVdP3htsrphbtuDd0/F7e5w2zF
N0yZfT8eTI+AH44iKxsIYSq6XpmeygCHAMWYPzmOoeaEnLHUAwtF1JWcq0Gd
/6UYsNWlk8A+2cL0raF+Z5qGfHNDc6wjmmDpYJqhlFkmeuxJXyBF9cE9Zy/m
bCUUeuP+3F+cZHunBusW3YRzMWdvcLAeSVbfJ/sKw52rHwUAfEDW6fCm9ztb
oufHsuRXvwFCtnXgFuVs3bajVGnJyJ5jM2dx9hcxbD4A/nhRB9kWb2P6mTGV
GA1qemhfiJq6Synki9sy7V2Mz+MyUTHRzF+bSZ2dh8vMofxiVsBbF1OUnUA2
P1+Lr/0EZWmFyupz5mhgtvHRx0pAqUEuMk6AtkQpujC97DdW1zrF65Y+1NLd
I0cGfGjTbfaZlqJhHo9SaVgyqaPS7q6sRfMvl6vH5sp9zPoAzpESlG7Uw+O8
Zpl8bBOWMEKezZpVRGr9smdNk/JYjw9zmT+FK2yVfpz7Lgvxk4exf77hQVaQ
J8zCrWlPfSpbgrKaapKD8p1iJcpdYm8QoOcrHv9o/mrI4xBRGj3PgPOeqa4/
ilQiClPGfapHpAGeHQ53c8ouaNsmMHBhaqbjXx2hAXNQUzl1JMsscNBUFCtG
CQ6rCY/FFpYXzWUimnuA9HZD940lvnxCuwipVHGrD+/6n6yyC8x24/MxMB4X
JFogXp89tD8Tieau4sVSGYOnRmzwZMWe2JGxbdwLkHfI07/yUyIiukS/W+BF
AwM9GFGVsUxpXqgmIVKpkGa5Fk7CgBEukvI7/KE5jzMyVFmTr7D32B2Jkc/4
rR/qwgqMd9QUA/dygSDpUprDXpjXeOy0sJB/rZ3Ea2dMOa0N4miVY8xZ4BF3
swXy95DuTa6phGCFwf1o2eq+lrmPfK7728mnmQnWOdkOongk/IuZE9W3AEmI
iXkv/fY9adxZ+3VKhdz8sDefqO01hyIkjUng1hVtRzW7RSqrULkFiIKP09Y3
Ok/EJt5IOdphJA6dM6JM5MFxeOgeMc9DU0q0SthLdEBDrX8OJDez02gOzM98
+hbmLTglbZcnGlp88XM6adY4FbIrH3ODypaLUF0GI9rBSg5nO+/KvcQCz2SZ
byNqICMmQYo1/TTHFGdZgntoP+5VCqVAYbgShYjegYjYwZcuhDYt+yioASnD
aF+XEnoK6UaOMndl1GfFRHuqtwV1SR9AY4VWZD0Hrxrm5PJIjX4hdC7A+P/o
TCGJdtQK+/lOuTpu/AqMcRHbI50xw6hLWGwl4SMfaXLPo/B4awVYelPBz5YC
KfnjhkeP6jbMnGzO4uyve6RS5KU8sXSCVfexvVy7e71TYdZ4K0gBScM5wW10
xGuvXvZqycuAd7Z+1Jku85n7Igt14Op1iv6B2p/oiLogEGB3T8io1p4qrkJs
I8UrfsvJ4QtYD0P4a/Jal0UhIjrzxqK3piijfce/TScQZ6LPCfLQYshvSK70
BWScQE2t5WgejO0kkT3UkScHmJ924ZmQpqefzxbzu6FA9Tj1VtvTPDkzI4EN
5zcAK5Nmocs2QZm328kyZYTgkhVbJ/0zW2D+atuvk9rhwHAJE6FHebRfqztY
HR+lxawlO5H+RgcimYOwz3NUxgMkQrDqO0feck5ksV61N7R4MC0+7c24E4d6
i0U6xGZKyvzJ6DOH2gxskqvoVStseJ3I6xKIU7WcdNW/gMI5ZLraawL15KSt
/KPcpUY8welVsfwAXZCAVR7zXOVID/RP9qRa5gPajR7W5bfP2YipZSHHdBuj
LIxevCPjaVwTvbq9qPNFpXJpnJ1gkU1lJWi5PlD6+BpSt1/oeS3muEwlDTvA
a8qLXtAncvJ9UhVzCN11beJoSEzCOcPhaRaMmuj0c0YvqT6ErOMTgfh1Ca+Q
9uWBKgXYefIILowqrmJoW1AMZrcJLjJEzLUrcyY81vU9gnaChBJXuClnEBHv
//l4L6gWk9Ui4esJoAFiA8IjNYn6Fbyspg+OAoVAf2AbsRCX+u3BrgBRn52w
l19CGxqwrZPu596yAoIi5/jfq27qzTToCGgs9N6eixGjJzOnr0ewVs3siPbz
vQuQOoGrkhlY4iB6wFAsZHXrM4DKp+faQ/7t+9KYD7Uv3bypzGTg0YBTkh/V
8/XHc/1RoU5JJKxU7Vyv0pjc/0ibSUH8BAdVttU59rIu9jb/eU9VHOu3TM6G
Tp78ccJf6WI2S1faXYqsN6zpUrX92qhDLVe+Ya2RDSZlWgRN2h7xJOewXlbe
mtYzFLjGgSZWyTcd+rtOT7wdPLXnfuPQoWlYVdgeWUUMIJkmrLjAvTKwwv0x
cyU0b9Vt4Mgs5A5wSDxD1AYj4AWYCCQrn0+vFl5ii2bYKV9t0jQZx8MJ/DhF
OQTJFykFfcFbShmRvp32XuixnkQyA/tYMyN1yC1LJDE31LKC/rhrC6i+4Y5u
hxK3863M9xZrtzit0Euju0gEmwQPkthGxdEAMgsyDnPiv3DRype5i0/svjDC
Nwtsu7kbTQu0FzaGDESyM3yqaFNYIqh5GgmpVUS2r3UXL4tDRxciVLEJuS8X
32tJ1bBbyhaCfTTowWDD2ll5Wa3RITY/sgZySSiY8l09Ii9TjTMXWVQZ1vxD
mtEUo9yWHJ7zGCO8w0LUXFKnBzyQhNrzAcvj0YCRfR3vuhdS9OuDj0eW7Ny/
XbaBNzP53OLyDLK97t1twAs6bEK/wrm2UFLnOg79iJm8dwiAZhwyAioZOILU
2/L+Iv5wCRlCGWm22hoYSkYs83KLUKJ1YFmFpLJuS5YInTCHtpjcSEzIePd2
f8jTmU6q8IbbgqZ+N5Ct+QCHT9R0WQEv1bFEi54OlOK7Z3+z5pvAmOjvf68C
M1hH934usi86Gbrj3UK4hmLzwS/vnE3P+uzez7KSqeaikI01wAluWCyV5s6h
pzkZfaWDC7KPifswHZ8Bxq9SljIV/fHPBmivf2Nl9QOcvo1W4Sqj5yUdkV9k
p6QdtyLykBPWMy3sPeJar0Okm6XwNA+h2XBz6heKzy0CX/+sIpd5LRoEQUru
91yxW8fC+NktQgLwd/W9J2zf+MX0pbwLa2BSpmMFz8aR00EM87NV2y9bKtON
hNPbYBsCZVFQHoIvgJvO92K9FPIR+Epdu0PVg8XqqO2iV/qanpQlpd+pEowS
Us16n3Ad3o5gP+7V+1MgSHMUTB7nYwiroCbzt3jo8OJNf1iD8s3jEv6uaPPE
WAkbPN4kbrFc+aiPW934LKitLvUGHr9zvuxtSCqGiAq0Kdx3NxR4OdFfZ6dq
PUDgdsQ5HAL0i4or80YleXXhkntKbhi/RwfF5bPIJQ6aJ+pFNOmvDm0HsDlg
rFEgBMNSJcc/f0+O1sahDPnGzCnF9UZ304pmE0bONXywWIWZpJOMCiWztOGG
jhRIVp56vCUaI34KBWhNWl4i5oJZrmQDWEAcJCU+RT/mj1wEF8OKqJyqEPlF
6ZA6TeCI/NDyM8l4rHjV2JK3yC5iJKkS+E3RlkOSdWUlZKrzhv6EG3NnkFQ/
Xm7PL90Oukqj9IRfxt5tpW2aOoih4Iiiud6MKEWjZzmwB9KRscB7vwB44w5/
h3h4EYxrRZiowUcdEa24qJt5TV7n2AWHUwC57suEQsVoYeZiekDLwjcDYaPt
ncaMjY5hWGIfygjVPWhfm6ufNlQQIpT06uO5WoPDtA/P93qfsVU54TvcdM75
zVBIbD1bCWrW5KRC3iqTBYUHa9RJAGou/NjLAE+aARFQgRM8WYND/kwT1wMA
2s8/V9MQ+Yd1uP2myc2EF0i0mrXB9QbWnwJCeQ0LKCcXqkhLMSl/dS5Z6Jt0
odBCP2czZCrR50cZnbuLbspKwuZdolaArxSyLrOMBnDCfRllnGnzFySLF4Pv
9vFT3ajyIBbFK+PXElIIse1XovJiLw8SfatEWmMZFmtdrmhzz67UckhjfaOQ
vbCgFduUpqPMjM5rPPZWbgSbkR1mklGP0LhRP6xtVsdMGSX49UEiT1oLhGFe
MedwSTrKMWa2Zp3L7jcYLH2zoTM/XO6ngnwz1Yfc/n1ad38f/CSQrgVcyqAX
XlNg+a2niyeVga7wX5yVVrPomr6m49HHBcE7ap+oDE7u6/xuDLh88okB8pEQ
KBxxijO4RUe0JqqHidpOLjojwLdZ8gC3NYivJpw1KBoUGe2iRUu8f6Jp6zSY
yocggmMGkC1Gt2IMZ9HMOBVAeXubQzaCyNi3IDOAPHRWvbdbWNe87XfsuVTj
KBcnJIoEQGQB5GB4CVFHGYynBvsAqoQZa6YB4HulaZbKpgJT4EyrCGEgEYKO
3ySwDfXtxov71olgXWuaWCpTsT120J7aRQodogNLUGvdzJGrxKlBdF1CYCWH
cV30KskHViQVIy38GCb96Xx1QjujxMY3igtAmj6a4YQlrEk5xeJRmDxQMb+U
bARibjcUISquaivBw9BAsEAXsuMAd/3gSDsp5b88TM/3Kib9YnGXiZnWjHQq
7qblVxAVAGoGY+fwKxOItc1eQoUpzDVBsgGxamFtYNzcMKASYiWS8C2UdzrB
mtvcl+K9U4nUZPCzWCOU5MM0yBMxB+JhqGKSU7ZjekSpX7FAcDCf0wd08I+9
+JDBTHREBMUZlCoT0ZbS4kYUTtYD7FALbr/bz/npvGumVyIf3f4iJclamKqu
3QoMz9dN8Pf2te/jJzjfbeo6O4WEkNJijD7zRsyQCMjetmCiMQYTHnoQK3bB
wDpomdHOqVLUvKYPjp27sREcOHdnVAJ8S8B2ZtEqhADuLbN6IdsSkNvYmaM0
+khK9Ucd4hDYphzYVfMW4HlO/zWOfcyXgkb2ihd3wbO9ljKweZ3NiQgfD91w
q+H1dr0H9X7VpCKunzgEJ9vbeRZWaA4fFC4RBhUfbvRqDP7YDMpVzYKSRqxa
Ttk8016RTsPdJGLnjmu3HbViwkiogWIIuuuUGepVYzOYdAuHsdRidvcXMv4D
7v2+fsapbBaAb5BBmacVvY6YRaf6I2GgXWdpjLmMr/CELeyFktgw0fzr+QAg
eqWB/0Bir0kXllvoB9gfUj3gOVKUN3TnLDeVM47mdmt0B3SHjTRuzv/vol0B
mPeq2nyxsAdPZqPUHNvRUBZDoCzjH7RWibr+Q7YBIdkyZBDdrEkVAonnHfAl
st4/oTSxcVgYjnZVRQ/OV5lRqL+fPgbNTWusGWFJga9yQAOiAMHLObZnYcxV
GY37vnEXzY8aFcBB8V9i3MH2Y9L25Dpza4ik8o8UQnsLsitqvEhcFlSBsiSb
rkXS9tn17AZ+hlPdTM+ksjGHclWHAzdAg6qb8YsUMknQjIJ4Xj6Ru/H2Scqe
3arL1TVU/MxUWFbkKCD5F2tsasSlcpOPqdp1WPfyKww07wIweaQgXnpMHDuK
hAIC+ST8o52LIQ/OSbbACMri7sufoYM8G5qv6XedB4o9/5SDoRJ8aVtJKLTH
d5iR7YUW7wmNQRiDamccVQxPMMZAYqriUmN5GXJ7cVfyw8gIXHRYFxbbB0oA
zUZ56nkFKP+QDGgI7xO5MwB+vr14HotE8JfrUsUGA87i17e2g5pZrE1otA/I
XW8YPzKL7m/UGCKYDfxtZbLfPTyHL0PZ8O+wuz9UzA3ZbxVLobssuu47sPad
RAzI8cgX6sIYSz/BnjJNtJCk+CTAtegw2qoqkWn/J7LA9gktpIRt7iPTUD+N
oXYhsKFR5V4imL68vmYDxOI7omNrPevP33JJIQ3kfNsqq0r/4LgtopyG0msO
U3DbltWBPm/s3tCpSv0ghXaH+/TnXkX29OOnjF8j/QdBBY4iPgUbkD3/uuay
dk9IEjc8MteYReko8G3Wc8ziido1JgVeom4Z98BohbR2/WyOt81XrSwis6rg
knCH7vm46lcV6sNqwlTFL8l3kY0AYChbzJIGbDpzH9AJVD2DFpqYvZzE+1fC
1VL61dUZf0VjBaed4RiVMNVPu/bGjpVbbVnVeDJE7ihOBFVtWI/26SWT4XAP
Mwaj6dGYXcOydtZrAUVijbzdWvfMrtS2BnkXZMPsFl7eCS3G+3/dBOBMA0Oz
nmsuSJaxhy4BbzeXRpPQF1+9pyQ7FA0KEvJbOUMoTnUHnL5TJJ3pj5sAEUc9
om1op8/2UxTGyL1ix/sG/d7czivgPg1hluikvYnMPD+7RpqAOCkW3aZTMuEi
OjtshP6xFumankweVwju1jbeFckyPfsmAfK+rp1UD8lqc4WMcRVbSqAA6fPz
KDoyeM5tiynxcGWpOMcfNJpbTmTqGEu6bkr33iyVDQvWzXRSAUTS95Jk31BJ
4B5qvWp9SVAoS/I5iepGwuBI2S/HrXQaFAVBgslcyq65hngK9uTWvh7oSOHs
4N+ZZw/0/3PgLzfPm7AULI4WN8jOEWt8E+EZMWNFIj7eSPKJIDZrrjn6D401
vGI8bKzvYC3lJlzH3bTrO/nTfIVdEvAxiW28dH3fY0uLONoQ6LNmngM7rp6I
c7ichRUdnLsHdx4gtHKz42wNP5S/fMqC6UHcaQvAULgPickipxO0fuiQ5TGM
v71DKpSRiGSbb+WJFkLrUk3ZoPS5WFIxQWqHCf6vVFcfeb6RL8y5U2ymIia0
4BFKJkoV9qpKjfjE/muys38vNrzrZufEGCH0nWzbx+JTV6eapZUXAtK3cY+Y
BdDbhk59GkobsnFS9cLza9++2QqHAxrL3J+dEqXNugn5S9E9G5N3HDjdgmwj
Kd4LkZqirGOIijxER3F69cMZXw/2Pk6xgnRUCyGhPUfQg5tBP5smcTG4Kjx4
e9q9hnbjsRdUBQIgVDFGmFaWcc/pDxBUTqMmoAE+r85d7nY+6tQ0yJJ4Yn40
hTy5Y/n+9mweRigwLrFRF3hqtDa1ZgGcX2CedpL0zd27srlf8dfq0Kudz0jO
lBUdnsQ8gtCDhSX0bD77nS3FrIocfw8tgby4mLN1aiq4lFrIPNOFb7oAR+c2
RuUNxvmTRiuqBG1XbF1Xunrlclk+fyvAm37jahWAiRISL/MfLbkbHbniOqnY
lahbscK0ZNYMw+aq/8o/d9HkzUXilTX69ErLCYcih6F6N9rTr2XkyRNv2/nV
yVEf4aVFR3oAntuPnsY7q3Tp8wM3s9EmfN1IGEgAscjEGNa2Mi2sJXvrlFu0
95HDlT5oK1zUKgS6uSiv51jQjmQvHry+Bmv7EgRADAmA8W1/xdex5nN68BoQ
LcWIchW9EHpPuUtTbA/YpNTyX4ocZS+bknEhMzRXP44yCfhD6Ms/8b3MKYQQ
R6btrEgsncm4RRxWDpVwmEVTGuiOZAOemC8c06QoR4gBzbJN0APx9Xj7PQh5
0cZgg8KRyWn8jdBE31OdZDahLQt/4f9B6/MHU8keJAatNwq6Ycmx0l5ZJ7P/
R9XbfITu06/bJ9J3gdpoY6eR8UivxnJJnjEvbkwtkwe2QWLxxRh6uCxtl8St
4D/tSF1OGKMSx3Vph0DZVOfmXAPkDICz2wtGePbR1PTtYRLBWOWAXafsusYn
EpOrMjikARpoGhjyDH9BYS6W52cqvZnI4bWQMqiJEZ5LLuIkMj7A5XkNGDuY
1VyYM/7VYy++DVxXx3MHWFegN8c64hPfvL8ZitsxGyHENIhkxnqt0luDEccp
+c9CudVzoJQDsj7nI6q4UTww3jSoi1sDIkLGM8mN0lnhyzBbqwVhgajRpgNZ
B8SIckMkRH2bziwc/pSqEyamKBKpr8RVDqZc8hfkdkvnr7ytW10Q7ocyvfEx
bwBhlDKo83oZpVqiFLLjjZYWhZrdFQLXkzuwXiUDGwyxQSB3/u0QjWeUlIeU
6SdwkUXOASXr8dtcAVGC3ePzW0oJHByVIjfeN/VQlJ5qFKu/AizG4Sfd2B2j
aTsohzkXYQcalln3cb/93HeYi+mu4cnih0kT96YAVBOEq0VzCMToiBAPIMOD
x31Zp4FqWWhOCSMh1XjHfkZJjMzAJDEBoZWZr9Ri8gKLsBJE+SlzHhbRiZGy
ohTSp+IiihM+9UJtlalzBKf8zwNHqGFhgp6TS5CQ/FESl5b5OdH75kuHs81W
rBTIy0PytushJReWvh7RyAS/ea0SNIu5OUMCF9Qj2IqEjikNizTIOjFdJLfY
tPBOQLlbxECgBd+gsyWyyGy/93gfZGUQg+ORu/tSIBoHAAspOpJR5baBHsJZ
p88G4MxAFey8A9cGkPxvlcFVH913y5KnPX7MOiuz2vAXWtKJqehqYyCxZ4mJ
U1ahagFcTfATWieA5wAYTIHsXJfnqEJUqXgHDXdHsEvxvE/UGRWD6VxAur+t
C2473CepZyAe9co9doJndYMtsSfnAROdf+S9JSxASzykiP7wslNYJgVwiG4h
skxt9CAN//2r9dKBWG5c65PhuSB0M4yNMqbu0wE4GRBs6WzeP9UPGA/PGsZA
hEbCA2jjPmppPLAhofZuS7YjICTRdwELukmI8xrBqFh3kOzy5pZKQFnPRd7p
LJdl2uJGuT5uOvf2QRBXWiSBR3pSHndzS02v9d0aCjZDlt3/D+QHoowVnMuA
tDvj1hfz8hXpyTz2hv7fc93Sn27M+z71HyQefxaKYAHczhsw2YlIfnG4cpa/
GqanClJeFL+fwnmEKmYE+/45BeBqCvoLI/P14pOjaqu7TXIUoMQKqDKp9/Gk
CYnXtb7nwtdmk4AEvzMne7u9SPa7CX0YK8XQvAOo/B7rIQCmlwYptXMcdGDS
wyqD5bsP1Gpu1fJrv5SDjZL5wEQIsatGQNJsGgvZN0XsX0fQJlKFbzdOX3ep
S/qmhiCgFab4xoOcgPetOj4DfSy4wz3WJE9/2cddxk4sEsmQnF8IsK1JH+f2
BS8y38EmROXbM7mf6680zzMehWTnh/NuZjOr0vh2OBhLgOqlKnv+M6JDbhx6
Q9QKEqbFVP7TLbfveF7kBbtzZjLB3Nr8EO4jBtkn0SaJFTt47My2R3UBx2T2
oDijZUSNQ4ey4btj0Q/9OC8znEQ10xn9+msTmEKyD3gY+7hHUUiEFvAIfXWm
9AWkPHQez6ozHLOHocg8dUAbBuXR7wLvUAN1fG/Z8wnHiaSjEsfJST7z3ArJ
cl1mFjYe6fC7UmalQyAfKQW9za2K7czyldwy8wvk+1E3csdeqalmlMu9La6P
MeboojjINFP5/OTa4rmuSu2axC77IKQmFz3LW/cxGc/215lfTTjFtMsAD4Zj
SlibtwCqTPQaYbVjFbdUxVw522mne976ICOTNZJ4M5KmOpP9h4AMN7Zdrde+
nS7hiU7Uo6LpfR1FxwU5QWSFUWRD/H0cseBpfwhUmAuSByoZ1wO/rzyTYG1v
aeewaek6M7G2Gr5tSpwJEAuP+7FW46HTK8gY7e4BTNgXhuQLxKrUuzY0aFpt
JckLepAUJ8BmUYwMCaL3KIYDE5vxCLDTkepW3OLwerP8EjnqHA2dWgFJV2+T
cfU423cpjCDJARzLYU75uh3w708rBfeFL2AmQWk1wwgBucAEWy45ZDg7+u2f
5cepk0fDgsuQSJjRASpyNJ+no7cPl4PQYT+n3TQ4sRDn3HR8jyGIhvsAR2xF
R+g1zagpLlVE+FpwoO//iSOTPL10aZWQHepQKLQiIOJIucXRRaMz3u1T2b6X
Pk5EtxjnpSJfK9x+bL/3ehyGY8GHn2CsIATVhulK4vELNCgNfdsQztwboZgu
Pfxjv9PO5L+NvUU53ZNKoB9LMU//Fp0XIIMfy5FieJbtOMqVFr3nad9zhmGP
F47T4oYcZWY/Fw8FsuUXThcCsvUkb2D5SkW5gSIviGoUPTkWxgIjKFXeznSo
Lq0xTgC6Wm7RRcWxTYmzMQZHzUcjxDkAF9F01N6doyknMm95sGKVtPvbmn9v
VRVM5fr/4Bj70ZVqLUAc239QTyrW1VEEw4jCtyXQdaFoKq4eURn+3MuRiGjV
Qf+feAsnpHQAtOf/WN0Qg+OSREbWjKo3YD79uaVntOb6ufNV5AcHzHEOVd6r
4TGctab+nxySSupjVEIKt6UHbU7i2yky7BDPIzp/p40kz0dTSpNvXbQxRsEN
yLwsvPZx5Ud13X3HlUGlrRkwcnCi9n2vIh+vmFDkGPvYo6FhW7xfm07YhudR
yk4c9+6Er8JtNiY8TgBgv708VQ7trymVbMsEKE7v9Nx3+sLUQLIWHw21jokQ
jJHEjYAbDDApbWfcdM9Twt16Hm40xwc6cICWBW4s/J3N+XaWeBZtw/QfHnwQ
i5ysVyz+FyjEfNVUIfT++6MHvPp4QeYYdpiy/aW7ByJsRGLOI+nsQn1nSeB7
pVf1GDxIV5flvwGSV1y2i72lUan7F7DixsVtVs4KUtDomF6d1nJTmxNoh2hD
nqr9o6/kWNrsO8/xFXrNKy1G3GT/GdcR56guj6EBgmRV3WBs55DBg1zp7THE
4FRwghmI8gh4qwrbN0vfcm6lgxsRqmscEpGKTc4K9HxK1veXeLLUovO1Es1C
MMs+LyUq8nDMUc4pZ3Vp8Qyo1C5+no457/XYwpEqtICS10QUsND0xAYwrJ15
nQLGvgIbSlG2ozvKuERsQ+sx71R39yiCwvMlhh1j6VSsoXsV9qiDOi/wyyjv
kuZBpJf4XHa4kFlNogD1twARrF+Z20akekN9MooaWAKRc5xwWDLGyd9B5Oix
Da0Gd3ceQTromlXq8WsLiMDDV16e+liUgfB6E2i0q/ahZSXC3PcNBqtLQkDk
Rx1XGLQkbQQcHZQDgn621bDVbLl/BWElXZTnjK1Ccr+cwWZx6uAUK8FJcvih
eeyeiAF42WxOl/JPSO1Vt1cpQL04BO5fWMwsxFm/lTgnvaiTTc5XNT7F6meM
6z5yWu0NB3IWnGWbpsV+vBgJ+cmQxj0iTdUxdi8dDnlXu8YYokdyj7LpZb7i
RNKJZN0pJJBDO0S1X29MNIe9bBAyhfE2gGf1Gt6T1l8rXb8nY7CvgVZVTx/E
5JMt2aZn9jttwzwx2d/+INO76FcVXF23FkD2dY1wO9GcBgE2LWyJGoQC9LJ9
rTT8bN5qdAUFyqpLwoe6wblfLSrcKO4efdyhv+LDtLx8hduNNv4mCtLkq8fG
r5eBiA+G5raU1+0wKU8SXIbrITmhikCN9BCzEjE9+pDtHES3+tBd0MRdqB/3
OWQKCmyNBbDdF6FGYBAkaHgkFRfG8rJW3qHCHIksURJ+zxaMZW5fcRptEscU
c7F+1FUhctgJO5ZChg9vVSR/EyeQSUoOnzRoaE8U+Bp6t6C3v6ES3wQI+pGW
FV6TLOiBnpdBZeLUsJW5ZUlwKlQ//EK4yBLgKeUGaPJlr2We31Ff+X7Q5PHc
rtyVQb2ItlnBwc+RMQ8rYhwe34URzz7EV4VaV3cmbwXn+Qyj/QxTMJLcSjay
9lFBD38rE43vUVeUkwtJHtkwFkWUOwmBKQUmmI0IXlSGDoqZSUxQpcil0a0F
5e2AtRoXLE+q9RjZKy7ql7vAQxzdoVK2wV8HUXRXMToW+xlxUhMxBDXmTPFu
FXBVvP8HC9tk7JiDuHLnHxqdj7fFfvZX/P8w+Kv2jaxfgFcYu1wyKa3g4cbL
lb7rD2im6UOK8auM512HBZfyBEb9dpUYmU2ugo1JxRiLp1XrRdOuU55/0uAE
16VAmk/otvIiP1/DQ6P4nXQ5Q4nVXQ+H6R9gWehO9bNpYGcll92fdWEc0+Vs
W0gUn8oFoRp4D9bHPLNj38ZNNT0IInzCHuCVIItnCk8oEzJY4uqFjSVHIqMg
OVoph6R+DoZ2eKuIOm+hB5pq1vobHLqbrxpKVXJMfw0Cf2AXcEg/slcU11sL
FyFms2P6awZuLeFjOL3FgE1ODvp2dbBPCcKMW9V/Og6ientPkLyT7bHziZQe
u7UL7Qj1e3xO6J7jIkWSnuohY1Ngu21VEzA7jVozR9IGtSekWulz7jQ9wtNq
zOIPmEdYsdOZXBc7VBQHZXHi7noCxUlZ5vbAXUhir6rWfGHQKblmbMCnlKrO
SWqsX2nGaYoZB9Ne5HXHaXTAnL4ilBvws2w9wsxkMs1u9yc9h12WmU8YVbaC
y6tlahS8KeBRv1xCs3EywbOy8X5QJCBpRtPvOP1uCDgVmtNXXKv9qOVJ8zfD
J66090iEb31ueeHZXSCm3lhBPAAknWymvgCRR76JixJ6sG3xlzzOXgcQyah1
Tb6Yylr/F3FsyU1GDvWli1rJhqAAOdcsPPM7CDFWiFOi6RTnxhVwWYvgv6wS
wcuLz5gYzHbuwiVsjgsqART8nZxclV7Not5uGNj7i2KGaIwYaFJa/eCUizL/
KzEO67dDHfVxMHNp9bL3z/RDOnh5G0gMxDkzD4hN+3IOrYizQaueAe8P+boX
+AC0QBl4bA87ETYfXtl8YhDahm5taXv1Tq9F9gSVIZoUoVwIZSC224ddq8Xv
YpGrhlKfxGXNa+qOzzoqTeZNmFVonldTuT37lPi6nyE4flOhTUEUcJtDNem8
M6SU5XwKBkkNx0OYhvlgkOWFH4WVbSHQMJGGNfcJE5263pa/BDZSDdoPqWxC
bVtDqJLUd8uA73xIrTMskAaT5n+PuL5Nb8keHh8Qux8rJcD88mCdXjMWpWMe
44j9S1S2CbVLMQenT6ooAqSeq3FHX/eKTHtHHqpKrqIaY23Rn2ImZ0EFgzo7
DM9LAeIzUYVvI+NTHTVn3CvdJO7MUV4oaF59yoLjGjfdJNVbutaFlPTle3I7
MSQTbl5ZDEnVNFit/DA0p4NTZ5X5Ng8KKUlCW7wnS8tcuRinfOqhiJTbAPYE
7CgxgEBnCtuHt6grCKvSCfkg6Bg8rGyfPh59qYq0j8MIPPNeG1Xal9fUbRt2
dGCyDffjshPYQ0rR7ZmRe3Hkbs3GXa3cZKi4Aol81j7tDzMJ2KxcxdXgokB/
QGekfjgHUJ8Y9f81i39amYS/4wSgmsXhGPzthhPWw4Bxe+TTXq0ad77tol2K
8Bent2xQMMpNloX4vqwkZLDzMHeOzy9Gzfbg3aKOYn/+XpZyam+NpxDlIpWB
Yl+0JMvZAvsx6Aw7iWZQbqcFE+LLKNZc4aOpPDZhifIxBRYA25b1nE69N5Um
9rYPjBOD9HD/F1xJJ7QUUPGUqOphNFbL2MSPW1Qp5WRmHb5WBkujBHRQ3F7H
GxxqO6fyOus5pzJu47VUGmoj0DLqDwj0e85Abo5Pk0s7hL1Hgu5o0gVPrJtS
iOmnBvu8sLxJ+5Vu9tL6l757rDm2TWwkRGUPe2cTAD2SwoM/BIyULWXlOfWF
SzgoXKxbU6oZBKHK3/Wy++DuSCPntnEjon///1pFXg/0xoeeUvbLH1EOAZ3k
7x2TalcQPIRlxF6VYqulOSqExJlGT1Hu+I2d9TsARyaUs/pYa2TkqFCaZtrf
Q23Q6ggf9TmLbz2UGp9Dip7Hucj2+qUsDjAEehN/tYRmDfSQznsBkh0nGbjE
jwIrL4nRIeWbj9G2skeKXt90gtxYFIRJDpnKfyTygpnCM3dopCanV1zuBb0u
FgX425FTm8jzhYwsvpBog6QcyYGOV1wj+reUMOacH7ACWSsFl2Q+KEaCs852
Vlon1+GoPxkf4VVV9bIpXd5hZeR/nmPBrP2hpOj86MTx+iP8xNSkl3FNPxqZ
rwm+C99Fw7+WnRIIfYuqwdZNNGsGtUklWwxM+cVPM4uQRq7cakA9kO36Ze3c
/BjMIkp7hwiG0fevhhBACcA2abnKQbBYYoCtcM1Qjb5WqHOKFWkhyQFS3xBe
04XgWxK5CTU4IW2k6bfcpHY8DY1sczF6wLuibQAWhtrhxq+S37l9uIxJCqZd
pzz6fldTVRj711B0MyJVOlOn71FMI8Kc+OHGl54L/qD6CMZsiX8HQ0KKxRv+
a2/xLPj077MQJHTqChLpjkplTU5YIvjVSVYesv1e7xvWwKokHoarWi30caTv
CFnPo8HNj7+PIuB3VIXDprohsu610zwzARSfEk0SguZDrg6RquYbfQmEuAJV
LtDy+EVcjxjFaiufZo5BMIIF2Pgik6Ve+X33CpJpkudqHPa7TbHbb210kMNh
tMiocxSvoo5hSLQBn5AZml9Y/p2SX3AjZleIWD4HaLvB1zWBaKFqYq15a3dv
rgj5okvirfNxvwsUEirhNaYKtfj5VcOkxRGySaMY1DYL6Q0ZGHtRTGRydqR5
j7hZQywC5hNGSHPM6l7lPOSqf7tJq5oCBbsuIz3WVMdhi/s+8ZcZpXUWYmwU
V6/THuPkyK/RqzErXx67Zkwh45BrWu3UP/QG1h/JSDus4Ta4V5AEHW9X8wHG
jFRB55gC5HgyQOyp5Os0K7hz9dl5mZrccd6E5tLQDZQ0pldd4QMlDWaZaoQx
hdKEwEdKq8IAR9vBoT0//K6+2ZCNGy7JikWZsI0euMDWNL8gVaPXQOk7FnNP
Ha5pQXwaewPRUFw+HZuSzjsjWbdXBs6DdbTRkvMol+re5gXjMD0JkXzuAEdF
TfFw7afNnvdOImYnY1J9ig+w3luaGv/7ectx0vkKlm0tCFSRf9I0kI3QfDXj
3IS0t4/LwyFrPGxfkMyzmOfBEiMWcKnsYmsg59WJBvTnbid7YQIhzJIccj9b
j3GsiNm0BOFnjWyplOLi8Ff8MhNQNQqsnjlqKnX6QkT/ah0d1WmPeGQgQdMp
c8HZEOOyxWtBBkkLBp4eREnm7Chex8SDraLV7zgIUyWMJNIkXKsM/rsjPGS4
ZEmqPFM+X0Kwh/gNdSLizlBX8WzEgXvSpCnGimF5nxdvAAlziGlxjEm3iWBp
13x/xBhaaLd61pRHGTw24DoeOfe1f+vBzEJrGqYZ85TH6a4rYH5aJYmM2/3U
/sYcydb7x/9hLJKPDzJMtnHd1sPGzBdV0abzTUXqOzXv5GldoFL+PkuHhsCc
eeH3Yf49VKL17iEWAIiIeEQ7cKho4oYWG6Maud+pAbUpdQhZEKdQ7xwwTLAD
xDMLCl+4VypY49m++lN3ayNV1IS+r/LVT4H3ETsc7uLFmc1XhZ+OWArexgAV
Y2TJ75g/PQOeU+14MS8YAWOa7Fw1Ty2uJQjm3+MU3p+9/m2CoXzIrmj2yJmW
oZyZmcJYnUV6xgfoGIvTPXcia5naApJfWWcc6gGKwCAPQFWCjIGyTTKJojkY
jkCsLfBVqefIHL6zcmR6fOc/FaYtDClLj2Q3mPSSagZetW9iNpoZNKWuEIa0
SgWTDtbUOYuYMgCZnpzgVxdOggvJteKFmMFQiFRKI41UghYYvNpD1hI9hLtg
SX1K8hcBdwsV6tcswsYCPIGO+rFdX9GrMsLw34622WZUGWziZxkahxPjjN6O
eTU6TrmNHcD/TxAthaf17JTgUlJ+OoyH/Gg4tDuY76Ld/reeqOQhl+E1+qCz
9CrGAb8FcO0far2oZ4FoDjWwHdIt7KETJOMTm+dvMxce4Y6WwS2fP0QRIYOS
aWXjBkUX/tXOlpOguUzY4ZL7+DsV3BpVP9BHzUNB4JMKqBYA9GhWQInTl5i3
t6LFtZ/KfxvTayE+2ozVvMie9Lneh4X8DLoX3599Z4O06p9Csd+LnvHN68Wc
5hvkmZ/K9P38WKG/xwWomHFmafYvtD66kjNnY4wVJGivCxKPl6ciQ9Tsp96l
5ptiEZo+lvq8UMwF7THbg2mbJ+Da2aKQu7RQ6x2U5ve1CnZVxS8RqNWRgKB+
M7P8maBwPcNHYxQi6dQ9oPrqNnNfeIx8YQdJlvga6jsOzCXE22em+cgGpUJk
Spfnf/01yB6iy1laMkkTcFrjJYel6AynCuLbYeRpCZFyMte1QERE+TL2JQA9
FosTZ385rPqDzIeVcACY/8uXjJOmnF4JKIIgWmimMhqK0XG8CrXUWeLup3EC
j5nYi9ejAXuYrsv24Xt7k2JBqxgE97P5Wob9nbdb6v8u38Yuc3X+Gp5NTWru
SgQmmF2NZOZUWaTUCJR3DLUza+aqyXcT+lf1wO/nLxiRdfwCkysgn/dmJvVQ
BANZtT0Jr1+6ldLCEz78VlOAFmz3pixKAgFTZBl7VfjSWuwj5GfzfIyCYrki
YPIGcj6OXfH8T6dbb7vya7enFyafufiUeqo7DfNL+hhRtpkTzSYSdKqoX2/B
F1rplIhjh1Eubw++ss7vg3KKd58tRIEKSUUm36TSs1oqDQQ6RpKORu3bQ6eW
BanJUsrwPIsrLMxGNvzi/NOm66HgE+a0RnD6dvbk3t3sJnTaAFCQG/Ww5Tkx
PInddgJSFGiiC6IMkg68f6MlwoQ3ZMUAdBUyhL9aK7qpPZMFLlMoVMtC+POU
Ad7hCHwkhAaf958BUCsE7Jemy5PboISi4IbCu2a/gZ6wtkAitZYK7ux+GrLe
07vUKC4D4dkkS8kFZFLKlh/GXOA9kXjICTKahZ5uzF5UTPWlDCE1oiUcYXnt
Mak5qDFYQe41GRfDhR4+WptHUNL2+c2IzM1AoahWOH006NilawSATtsa65HU
3ag1Edy4KXtK5z+1EofGNt7fZ7gJ0y07ItTciqWBTYTeGs0r0KcerMAOr59s
XI+5bBmD6X1kgGcsASw1Kt5S0zYUWsGOjNYQcan4yFIe5FHf1OoZ2o51jK38
oemX5RPEeBOKJPxklZaUPvIKFABqTEDGphsCpc+WgjYS/knm2gxhRDt+wk/i
xsacs1I9HZTrC4VODK6ec+gCikOduYxdj+TZVgIUOShcbA4LYqh6zQNMFIZ0
UF5Z1t+lsF+8EzQdWHIDGelkDU3TL+GTZHHnYyGQeL+DT1pIrEhzdqx9+TmG
/9LxozyNTHliKEQEFzRAWel6g5XuRH/GitJKgEDPURb0MuAC2poFkGuoSRe0
HoDbTGP9L5ddeZMi3vOb7zGqJvyayLQnr9PuLjD76faeiBOQTN+8POE8BjuQ
onCN4xlw4mHqvGUEepStZxaoPCt71Ifv06SADyA7IoxELsbdef0a/rVwTht0
vL+U34pkPoC7NB0WV+dxP5so3pUmenkVoxaQ5lTpPZsZXz/UgdMNexqq3xRE
ZG6kIR/QTGQILi8Dbk7g0Ka4VDFXMNq17Fc2Fbib+8e+ubFBjNELA5EFaknW
B6fNEGqUykGtRc/7Op+FoZ6t//HSN4HnMJp8IEyagm/UPBEpCV6W4ThxpAYP
55w2AdhtDgYeFft8NN0qBAsxTqpZI+fqTtba3LNAe/wZU84x1D3e1AbKwkX1
+4qlWCGXBU6n115W7WW054p8BKnnPl6twu2JH7JHjWUf0W1JScEtD1W/FjdD
7+6ThNm38dLIYuLJIqxT/i8OdQq+c5Y16C06mpmWs/FXcb1GjTTV7hwftaCj
Uk+E4Ymq4BuGcmRiYbWnl0xOTmGQNXmTJMaVlzTuaLkl1r7YA5HXrE2sRsZ/
2HtdMGfnyZ9jWc6VoU5EyLreffA+BjduZrOFNeczmJRk1DI0Gz2/oHqGKlXQ
5LtwkUyC8xbjlNRl7ay1vscv3XIhJaL7KY4m+lN7t0FnJhe42xflsuzVusvu
NOR+N2HC9wJ+9VWnE5rlJI4rQQcrfiueDoIQUtnZcUa1bXDy87USS+9KwH+q
ccPDjWzOF9PvtP6T6e5rEAdY5piOFC80mJQeAticdcOFR0ew770gXPTAObfh
OKKa/P9L6EgcIKxmU//kvngVhs7EDV0pz6Fs9mZsAmnlGdMMrCMB1ArCBgOB
Ob87N3gJsE8rF5EOMlYcBUW66bSfmFb59hPXqPUwvW2Qhi+LsNsj4bfVid6N
hg4jGTAIzmG95Fi4vCM9VX7/ZEHb7bvZG+k39xlRjPoyXkglJ45jhZT4WjkZ
QdFRfMkebptYrOVPk1yNYWgPbmXiYDc/opiYPbtRtXterh5v9ujhwKfzu6Ig
pocxNq9SDB8pL4qjywdXhs2qTn1g17THVyKWgTEkddtLAdv2BUf4dnzvosA4
PYU7EgY8C7HRNUHxw4Oi9NicRryRNF3eNZBT6EZ377FEJ66r5DEZXbZkoTl5
FA1hDp8V3VypicWmMzSwZpOua49DdDcJmFvg1BVaRWgcRlzlCHSOkLFCucbf
C8hD2Qr3AhCWySXiAMLcsoqd++se4VwGTNokvpxBvzeYF5zNLYG50AffjcDh
/Mr+/GQ/6o5jJYdMotZTWq44H54prHWxXRYUt58HolCFBoSVu65wdmNQQsn5
jXLK/r3HK9+OwbGX98q4WZmNdkiZ6hA0dL7C7haFF5JFXCL7G8Q//mPi7SzE
FLhQC5yoX/8csKJTf1UHlbX0Hozpkr03plLKmffRGjSpA/Ro341195srdTZd
yWAxYK/Cal0Iv41vIHlunxMDkZdiwKVVXuuuZGDIysaZPeIBtKXDwI786eH2
Wgoeapszu8phnx6D8Xxc/htJnkzFtwCdCHixRsWTR4iK5McvK8m7Rzh9uSAG
pa+FfkOSUKlh0qzU16WFq5191s+OUxc4uqiCBkANmxtnSewgMcxJ1uu+2abA
y9RwP9BlV/nH/FlGMfVc74f6rG0xIACYWn70Y9+X3nUZcLMxRTLyLXJf82qP
xE9PtZkZb0ElxP0M98oa6d016KUxVVouVS33j+ItGP6gTa3bFfF2uNv8lHkd
T9RO31mVDaTwIJgI9qSeG1dTXlcsoGm5ztixnDGKKqhkejTAsbDnkq/xrn51
XNV6w/atE4QZhkL2d0RNTeNnDTDH/NtssPqe7k4fiMmfWFlMd6Z2UpTAwIv3
VYVZdE3ar9Ot9TPfxkTvDn//FbRyKvqNzjseLmf2T/OUDZp8RSWU0GbYor4u
OQNdxugNO2W0VCZRqXHqLC7m6v8CfAKX2YbI/7+XzLgHbriNDsT2T+X5sKJP
au1ToBKmcRygi8ymJTU15byzljuVnKUS3i7W266Stgna6tGBok4uIc9BYmcJ
hCduHCRsSIttNZEkjy5/YpsT47yqtCE6rvk3AeeNtEmsiDds80fYF9AJw1NT
1frR8S+Mfi9a1WdORFy4/jT53EyJj4Hb/9f8fWnkY7ZXo7AWtp3ev6XJOUU4
KtGPCBMtm5UQFy4K7xjue6xWbpSbb2JxykeABm0cvXyvlcLfksVXKsEsllCR
5BhzBiojTEe/2vn0Nhw9/t4zzUfV8Afu/DRLJs0ctUHMrVGWIIuWdyaxjTPx
vDwo6IWigYNN8dRMeM0SYSMMZ+pUkd2EpRhUSVYUDA/g4S90QDGfj0p3It5n
j4rQ3L3I1eoVyYnWNf8/comq2ruevh52pNDbTZa4HUvMgNJSD9MVpnCOaX9h
IBW2VhtMgydniyKAp+otkzeYlqMSP08vnVMKTrp61DF4LylI1g841n21o5Ly
jB5nksCudy4Ulqcw1NxIiIiqNpDCCkbJvXGXBup6Auqwr1TYAsZnZyVska20
GpXQUsEHNpJwp/ZO+N4jZwO6RcHwyNz3+HD36Hy4oaBRjjwZ0ufugzbkossM
r4otJIZ9ulyqBJ470PuojJ4Z+1Wl9izh1tjWUm8uO933V6rSr7ZHLKmzF3V8
ShMLlrstYVu4ASUj2QlA3p+1TQ8aHHY52uoReeUD3h43NeiHK+bLQI2cGN40
4kHhft000oAp04S9FRsSOb2qoYrMnbPlzWwrt1szBQRY4xPGYtnxaWjfFLAX
x/JOPAq2hbLVSTWGECAB7NzMU8JWRiXgeDsU1kNzBzt/bO46UrbzvOQ13bwd
DqsY38Jk6JNAsNvBTEhdfThAUDPvCPoAn84/Fm0Nm39zEk1b/3N7x859J5db
bctMfWtPnrJmIbrX2a7MrriwS2rhzi4K2B4XksnTtDkVrPrxhOCxGjlqV6PW
3ifggUZnBMaRztgo04JhYH01DAsv41T6Z6cPPoFUmC5CZSIhRkziZmitO8ao
XQvz93VsFT2as3SXj8bV1NyCjPWCPr/TVgv7mCQ6Dzi1g6NIkfDF/PZjMu3G
HofViznh/5PEnVMrc4ZN6mwvgF5+AUz7xodLXLJpzKXfPOjLSdBirPJRsma1
PWM0l9qjkkVrAUo9/vN/g/+Oj3OZjXY9yYkkJDDUxSYJAJSv6nQuHaniT3Jr
iMUy1kSSKn6blaKUF0VPZsROLv1Og2pQcnHEx6uZUW7PJA/phPaktYTmKWgu
diP2OroKWUBmR11M7C4/K4YGqDXWLJ167RtwacF2yyMh85HSyDTMkYwPCWK7
ilAlZsRAlhabsMO/hoEM/VJ4i/QieDRbgO+bxkMxFr3PBe0ZAqth+nYyUZVQ
VFNbi/Zx4ZhNKlSfjLdVsG+b7jRN63nX84KBOayTN//4Kat819IheWScxbwG
9JUq3dF2rTFj8MrTRLUzuHEhatlX7EcNk2VBEF95HMUAu6tPZYiP2O48ttd/
0HdugOz8C5T7s7h8X0mHw1q3CHMapkdbTIzYmw6OMmPy8+e5LqzBbwiNeuq4
S9wfkfE5JMdvdWd8aLG7eZkECdX/GZaWPUOiPqEM2n0CIjVtINrVVCjlA9dE
Hcr4oOKRyD7FJZlTipnIdO7sXnWjMksfWWI3DMchqMPj0QstnlutPbiUhymo
jPAJQDw+FSc4ZmeIpworOiSjg9aQ3UWNVyC/ZTkZB1oZ+ODCFzb5JNrrqGNW
SAh+rLERnXqTucT2kI9fsUQNhe/01iCYq/rtSZMM7hwj7w6QkmLZ4YQ/eH2F
aVIgJfMQc4SAQiHMYuOSG+RWYNUTN41RmZCD7SPDIEFKWaXheWfleRgoSdUw
QFB1wSMkEXg6VRvByK4faGNVYSkuaFoKu6/cthZzuzysFV/IJYyMxmiJzSXT
JzGzPUOOGpaAldYDuJFTUmddzKCi+5AMcu8W+HbHje5Cp1g+hbXNZmImSe4K
/5+3ziBybAb6RXwmIYyxvz+6jGwchqzDprN/FTyr0nzZPZ3xswUvYLmxDdO7
E73TGSQCaWK2D+dKVi3WGrRTdsiYQ40j99Xn7NGqjGoyc0XC5fCoguWeihOP
X4D5CfL4ZFQAgfUMhbLSArWzL7mGMLfRY/AFVZdjGUeYYsBypjn9TMmHaZUC
uz/PVujaomrEJTBDcPKLX0zUByOthdZe/myvBNz0qWYYR7+jWWq7cWT9axBR
yWcPjSClQRKPVZVpXOKw7cRbMaXrPQp7u84G8IkmXhWS3MaNBDKU4ptU2lvG
Z+oD6TQlgxbLjSMIt+t/FndERxO0eBQ8kJ5vpZMCAq38AWAAQOokgRvE7caQ
DOeJTLxs9m0yjuoMNR1O5NoA+PcutnYID1bmV4UQNlgLPkt+q91tMu8qQQE4
WGeB7oOr6rz361u7/VHFev0NyfbuGDQrPgvbEnq+RDX72mGF6MtcLCPZMR5g
2BXbeT4bafIWmQc3xE4334C6WPUQe+hSs/ZfLVBTW0zFAvc22NlKiG2xotjA
HNnPmLDMKitMWVSzh8jT13MRQsNfcZQ9KXiUHnRX/cbuHm9Ku3LRJzjqPdgJ
S5kmVLlYkKfiV9XGu9MREaE8VKzH5DQmTWVPTdviZ+fSBrf8XCCTrQJTD9UA
c2nSv3I1c6csSe86FYVa32t9M1mLUbIC2w3SQ9btaLNMLVAxCHJNCnnQboQe
fX/3mYBhf/ZweumcAPvA0O+8k6R79ve9X3NyJ/2LCJMr8CkEiK6DbzBHzkRN
nUfLCz8hCpw21iF68umdYIVYzmz+qI/x2bheidz1Zw/xq5RKlw94kb7JBcP0
ynIbCNxMvQQ9fiEHks8jO3jcJASdhtaKMjM0QzOwHt/pIgY2Kp9exjCzm76s
v3HER8mE9A2ydCibO+NXhqioUfOH4R2SLc55Jv3UHJEPja3Jteb6W4HoL6pS
HuOJ0jwLQl7JwODWKqfZNvcsar1kFhq1a59oiq9etghxC9Sc23jDVuYNlyYb
+gSwjWOKraQy0LX0pkniCTS/gQ8evpPpVxdEr9VG2++7n87GqV1pzDHT8YO4
GH63jEtN1JpvnNkbap3BoxpAePfX+lb5hGtTCWv/lta/5o5FhVrNeQ/C63nV
CYikie96TI8LqKzOyN9pRBTesPhPAbc9Kx2QmcDgG5d4erZl5sTEVyLs06xY
r4snDQ+HfmvZVMSknVYy2GuUU0tW/NPoLbgMNA0QDuvsL5UlxcqlqnV3BBHv
LagihtgvL28S2HR+2ijFoULuEaGf1Pyf87lRG6h6codKm7ZccgBoOGnrxN0J
5hEzNOgoj6bUCs4IpEsnT6hMwHlkQ6HKUjI+8zCwQRJuAOeJ/671nTlQ8Qwz
i4CBO4kTpbbtKMBrKYKUfuEXkSjcn6EDDqHqf3/dzMISJzTPqvjaLvbwPKEC
Na1EZxBDlWHAlXu3uEcv5CSIGqhbIQG1CGzRbmfwRP/HUoA0+5YoZFdaEb2D
Or58SMqJMQclavn4T5eSmYXQqWAx1MC6f5k8ByAjaT2VnLAHJynyJ9i9mmcY
4Dl3MymNSySpc6juXsKCr2iomgnzee9KbhRIWJJbq4Q9yru0GxaVR9MCtuHR
tBfQozOQfIbEOfX2Z2xUNkj4c4ajsZYB5+hoNNCvXaJId3jWnTX/R1MGEC6G
W9dt8LAxEfMkKWVYCB9w5XpqOyMkmaIs0FIbWGjOD7rgD8KZJ17TiY3y4uX7
Z5EkQHPcJ5wHfYYmxKFjhVOrX1boChNyDTph1JzqicWTLrOdUwaG02d3bs6K
JBz0myltluLkgdxI512gZa3p1WCN0EJL0SnzABPEZzeiAIa9lmK5FKuhBolZ
arBaT2yALr6LqBETzr0+9x+hopdLI7HlDFbavmOUKZ/R7LculafatZw3/xtK
6kcsWW33vOmrXpe3ACS+r+icbOkoK1XBMR/7/qBXIQvXYkvvDSCLFdfqg8CX
YqfsXEYdvMQPastBHyQwMHfmirAFKqPPohw3H/gC7rAjtG1LZY3SqddRGdEU
x6PWKypV98EE78E8Lx9t74pVRFYtokvq8XQbwyAoH93BXDx4HA7vGj2SohwP
KoqidU2A1Fo/fXStxaK4qEqo4bFjeoYeWm/rC1vgoM/j1tFs2iUZd8UAN12n
ZTP5g6g1DUPJLKBQiacH05fZwRVwrVBh12GpX+56zvzWj00YP31BSnPBcYLU
aSFcTV59vAERBEnJ4SASQiAnpM7/qMafmYzoAbgO2bI/cXHIem9aNkC1jG1/
4EbyHppdpCLXoW9hPFauun5YiWolDy5CueTzJg2ssAw4oZWJ0IcTToT4RaDo
Dv5o0N1PmwTjQsZ2FGrMVpxLNpHBcNqRPc2+rcK+LR5JVr1lzi1dtXZPi3qH
dXRkg2s+rRPIxgi9wbJVC6oOZrJOUu/u/8RvqcCOnOz5z3ib428jgR7ikrdF
MtS/Hp+JcnfyLKia1LmLWm+lB8QNphHBybK1zPkj6yT/BPb7unUL79EaG6kU
4HuvewHxw1XdkdB8s4Dwby/cw/2MekhJXHmBtrfW1tUjkAgKiYgurbEO6DD9
+WDb14WqargCQJeqUR4xrT7zbWsSgTpFNPNIggj7oA0pZU/1rCszyhfwwoYv
r2K4XoU1Rb1e85qxQytAIiNhbcIXXtRvV2ajGrQr93CLjj6cFs8c8VsGScTj
0K/iEnUqUERZ/16+qEqZYgjdSkRia8ycVidB3nAN2IQn1lBBsR+WKg9oY016
cIbP4e+XjYe68Mypiu5Idt0VEo+mFuDFHKljze5FvQ+aDU4PgmLFaw9kPuO+
jiMspdV8pQNjqAj7642B4SpQjWbEmx9vygNm+/U//ouIofY8er0NmxvW+njb
kdJBUHPBZe/8qMgp5V2TI1lyPTqL23IeKP5C5JmDzcbiSDOf6vUExhPKLZRB
60aWP4u0ydk00W08F2MFM1cFP6fbBc6bI3z8xHnKA/GhXnI9XXiVrCPJk4aj
ZCjYyfjg6TVYcMMeqvwIPmHcS5wP0qsoI52XQp0QHtYDwN0eCU3X6JZ0abc9
2Ojn+UhJn5AXt4MLD6AQdwjSkueMfcayO1IwDubTCHxiLs0yAm9b7/JL+Sgh
1O/lmG6CPtPWL8NcovlQ5sMFI9whMYJNkyll/yfSL4FK/gd4wmmkKHFnF/a4
9dljhCOBlUKBPE5YfftxmV71kDO08nAxurGF6fH8dd8XwARpFLgozJUqqpEC
/SpPP10Ik7jAFqkaLfhaoIvFcPXZM0/IovN/X/L/CMfwMK0TkJT0rNUG/OZi
ZcZ8kR59e+67O7mkmF03+m4RWFqtdN9VegeGbZLPqLRBFLr8hBqni++twQRN
pU3obFeKmbR9WozhGA0GJDRSd8kw/Uj6e9RQA8jXYJe0Msyrut5kg9fsXDAA
u35D0gN6IHm/qNZCkwZAV2jqWufZILMLJds/NBoBpbQrcFO7mBemQlKYhZCL
ninX2S3fP6BXQR5xrM6dqc21PM5Nu0WXZAeIGEnOFHBhTdaIyqElzaDHV/dK
+uBMABzMOwI0I38UDoetgx9qj+22tYyvaFCL+R7TUw76k+xSnKZciWDIm+sQ
DqHrpi21HEuh8zYnEkWiTwdD6pX6oQc1wOdUDND6kSe/KuE/Dej64iOS6t5q
uu5oegsDBroeAnGfQo61IFASMVxxcmspoHa7eaot7JzbkgUfm20AtQel6FxE
9NCwyebOk8y6t96KBk4DkO+TENvfk5ucNmWZHGP26cknGGGCDiNy1bhvp8Lr
s+KYCeYPrkRb1crOpXNn1liQ1EnOBs1QrXZEYDJw9RL7V5/blP0GwYeOshMy
4rkkFLbSj1RWQSJZ9hPDD7Z8pow7SlI8gz9vlmyYcXTpap7bVglyAXTY1NEz
UmDTkJyqisvnmJEms1tsvkqlk+n1GdSeUY/mFPTw5ew0e1ukwwYCzLsuN+8D
2DjK9ugxGDF6zFJQ8HUcPgI+mLJhS/oJUWdbxpTc8dTWl3n0razGwoQ5I+L7
XDxCoI3FUgb/O4ob5CSmncVV9q8pyernJhGh4cZSb7pnTvATzTwJCSJSj4ny
wwEskdvnpAN0YvidOZLqr9xMFb+5VyEcJl9m5sByy3AOhnIMM4FmEQg0Lh4x
Tbw3Z6Ovjo3SdzAA26XQolcF7YKsIMoO9hL8wERUABFz9OSrUgWM8SNNaBSe
tIiiooLzKAdc43qsaUhHHA5Qen9UKztF8gsITEnD0v4PXJPFDIsdB2XdM/Yi
7o4ItBl/XDcwMhohfX4qkGDiDPmINyeQ08NI6OufHPnqQbXHtQSEIDjNyX5x
l7famuGuVMxyrrSHOQTINpMiM44MkvQWWPI+yBac8VxWW1mABfGdTY5h9w1X
1qTCRNB7IC47m1S0NVuMQpjjsU2A0sad9eVBeFI0xlBFb98Qu8K53q4TOf7s
iSNsaUoiBz9py0AsnjNvl4kAvPRmKwKEPcObkcpdLgjP1ZAPhgSpC1RB2m2C
KxkVqI1SnqtazaoeVpzagTYctLdfWlTm6KOgkaPm8QSVv3PyPDophrzThUsm
Ht+LqQacKihOT6Q/Ts4clBbPC5i8OSPhleurLZy88DCHaB3nyA912lVI8xt9
li4ZnHI+KpUGa3KBf8W6LwniAv0XYPDxaBYgtQYnUAJadsUJJOLrCg4BtJ3V
2AaO/9Fe04IKbSeypo9oHlP+ZGSixzq6+XqbqgVGMcMYMtZAXyvblWXxo8Hk
v8tnyxQ+9ZzTif3w7NaJlSk1eCvoTMM7wwNEMfdmSDhZr13wv0ltE7EjRYYz
Rffw706t1SrLL3iqfyzjHwFXdSUjpFqWtwSHeT2AH5cMuf+LLQjTrJPf984F
QQ5JRWi6GeXAbyX2yfe+RFJK/yRz4maSkMdxP61+cUdzXsVxU0pCld/wcfNc
lufnFk3Rtb+1swSuVMvfdvRn882F/AsFURqLw5jpDuWdT6W/weEe7O/LaGiz
42OOjTxmviXMudeB5/TMYtSsY5k/7uufiQQD0b50t0AGIIP8mDrA/hgSgb0S
8uZkBgHnsIT+XWDkB7AxE7IRefAXJgRb2s1gW+ApQ9TNMdTKwAs+u+BSy/rv
9B4hROH/JXz6/idCrc4x5+24SIIpikLr5RkmPgTdZZHyOrhYemxDgpIiqJBv
OYBdV43eeqhK5R2jOxHWrBuymkbgIJEL7SLwsxfrVcwZKgMBdwp2UOrgw+eU
9L1xzEYdnrG9A1iN8wqMRDxEv5qSnbAh+jY0hksdYyrvkgMahaW8LR3tCGyF
us8LkImoylitKoHg8Ew9zppdLfVPC+6W6Mn5vfDRxBjyRcKSviT52hSFOEgX
TYA/NkiN3Qf7/Zbpe3XjTWc4px93DfcpTbSNnssdFMuNIYQwMgSmM0MWOuUh
OsO5pNKiW9lxpQVuKOJcCh5JYhCOv3eabHcqnuIJavpUxOuKvID+5qetDcLU
LApeTkP1yVMpmqFyikiWlhCLaeorcXhc/Ko1KFla8z6YExN3CUWL7NHgJ8dy
I7ceE6hc3LutCJYE2BNaTe0ViFSOnXsDkx4PzJwj77FAWF82zHvA0eS9Z9rE
qdUOwvq9QPu0v3r33zX/Fc0AJ6It5l+mUTtAYhVJNPow4X71kMytoFsrlHAC
eH/PHRpXJetin4ClJJUbDh2LxA7Fy73wY0CgMANVv090nmmX9y1lQEN5lw3u
+hKqpg2rHFHHbdTh9muLbeAnpdovMga9oUPA6EkqUqO/M78wrU/7uGx8/bDc
TFEbWIOrbbhLiH+bCHe5avtZZyj75nJOlnb3NeU/INtw1Armi9hmy0mGF3eQ
8R6joUP5363c3ewPMXPjIc9SOoR1+uh8xqhNN5UxxL2ESA44h6MrVY8fn7P/
MZYXXj9TKYnjWWmyp2nR+J0HNyOiZaEwdWmVLfPUeDJzJib7frmcY1re7zDT
wfzOI6OCQNQKecBvUUC0Wh0pHPcJgBIVbjqyWSMLEO++e9cCHCwdRiCa5YVh
SQmq0SdQDm/d4nZ+bJTR3CVocCn//hf454svFMdp9gSxkoBIAByyQpv9K9Q6
ZM5KI7tzkMztKVm16Cz/xs0FBrBQqAdIF2bs0n3Pm3OnDMRGUCWonuFrM+9p
rA9qqq4RwlwNgRSzduV4gSWBj3spfFl4uiIXk4KWgNbK/B56oBfdRNcjrHlo
ow6/t/NTcmEZmEbJzI+qGyYA+uCWIKVTGACnv892RrVfJMk1l9DTNvyPOsiy
Cs7GiI5inuEWIa9qi6Hsy6L8HIGaNYa4ISglF48ZLDz6uNvuKcvEZd7Z1l0d
VC9B+Ej+JK+4lw4cerXq9RS0IxQJRlNBeIZG2PP2t6zzUcH5VUbJOVu4LWua
kQNe5MMynp4vuxHM5/KA1h8D3IejoV1tjXQO316AW8/0h6Z51sVCmLD/8YJb
ZtYe4ETzUAbZ44XfFp4RZnsJ7YtioY568lSfTApRzGrS04d5zZujdHdtv5S1
gfehTzKJ0Mdq3gIR5RZlmrUnrm6JDyarwx7glJ5sBO/v6sq6OoBhjyAddk1F
DmIFZx1dnhtK781QA6YJCK4pULlIqB4nKGXziU1chiGvG902u12hckqQbU+5
Cg2Q+bYlaYzbosnzNBNfbeJtzpoGJkouX/Y6RkqtYRQqRmSArIhCobE96s+F
CHYf5Df0GST3YOP8ENd4ywryKiYU7xFqRRosCSIqKFaqMUli1fXw/MPZy99N
tik+DGH7BEKcIEShXcyuAVncJr4ojAkadpbez/cRjr/jgBx6tNGmmjxiPxTu
VBXUv/zYJr23cj6vVe0AJrhQaM9t1FS1qaILxijlA7Dxli+KV0dPN0gqA5hv
i/FdJ71wniYYAS3jzjsefPBoJWOe1a0/a2FKACSjrpax/b+YrXv8hm4dxh+w
gfmXOE2bel7k/AyK4um5BDnjZSsZdeTowV1PmeDaAxusmAEK1qdhrku8T/Ku
7+ZXBv1x73dPTvDFGZQJrfWjkGzurtOsB3DmCk96x1YjWrij7p2Y7i6cHukU
NZShblbPNQ6CoRyG40oBohg71dHWXU3OK32bGAE4ynDvuhCKu72SB6bdxuS6
jyh8j7spTOPzjxwNSHQI+2nwpB392SraRKL2g32NeZd6LgSsCE0pT4Q6pq+B
xHktA7j4C4MZWSpupCn5gFXsLJlTfiEOGzXZvDAYFEqdSKNungUO6uRuR5Yu
6oFk9qNvyrS8zADIcDSfrs1ZcchJOP+tY/yy3x9MW52AVE95fQCuddLy8RfN
GK2uM16nb5psawO3ZF4TZQi/m2VMNYT/YYGslexivTFP4+WU2Fg7Dqpmbu+/
dYMXKpI2ByY5XMLsD6FFFXD2qhfYm0/YFQQQVB5MjIfmnjzCati4dhX3F9No
/uwHDrKHiXT5L2HgHFPd/kqLFG0z1T6RCkn1WHiLywNHRLLlYeM23SNAYNUJ
QRaIlN69UEiEOxt+q+YUTvBQtGPJ9+pomkrmDZ62IEylLxifDTYAE8hwFMve
woS1LjwnzBsCHM6D5qi8qaCDQVc7ER9LgfrIwSWevKUm4GTIPw2O7xWWPhAH
tPwz0kQhTdQhMrBnEu4H9Zkw8bVhTc6jHZwpUTno10b9U72aHEN70YBIcC7f
O9B1D1lEt6CAwVsRuluCsfMDxvb1um0U8sqx+UmleHPkn9LMYryzQjut+/eZ
5N6Zs49Lu6iAPqo86rLvU6/185NgEL8TGLObSVqTfGwPdwA2YijkWX0DNWk7
YMcYQyso1aprDJR3gLAlZuQQB4BxyJ3djY0NurPM/FVrbIC2o8WI7qVPLXuk
4yNxvBYvkBq9OtlOggsiPJC9eqZsHhxCy5uJ/NC9qA2x7USsJfsqZyTpHYFg
xNa/s23+031eJbiPBvvZ+he0TcqgHGLOyhyBn+/57e+tXKoZYWZEHsRjW9Sc
0kY+rHTpEHta/oOD+9iocINhI/ytdZ8Aihoig3lQfJS/QB2vByjl6P8K5ikW
m0CcItofSyd24RXYfwvrsdOIj4JAM6hpo0gcPWokHlzPcz5rgtNf28mzZt5h
FE0hq67qxp4itoGn0HdbvJEAGcactAQBa7jTs2SOAc1a2uNf5Nc81wYwmcnD
oZI9zR9lkonQtP9+U2OCZjj/2pEoEu3yFEa9gN5QDmQC4eqp2Mb2BQYvXWw6
3YG2dWrcJaN1L0OFCRUGDGLKUw2/rHZXQEjV4lDYIwcIk4GvWQeuaxOWsGoW
t1gVt4RB7NvbizQ3+tMtQ+7ykltGKds8zCW89//lHSDEjtk0tzrPPvr9ftXe
u9PXZExu1qQre9SoJDetn06DfS6RPzsf0aYsd8pHQ5THBTN/+PLJGAhB9N7u
wIqaQiMJUKWwJ9IR9UB5ssAeGvb/2WTKUPFsJs/deC9N3K3QCNUxCTtaykxc
spyfW9qGVS2UasaenlLC4IfjAnyg6Ev/9+9alVxtTOSXEGIqjLfXjvi9TV1j
cy+dvcZNkHsnWlg/fSjcu25kmAGQv7oBy3revjLrmfm4w7huOT63pdim7Cs6
LYXYUTbSjy29/VDuCfnJFwTbVfiyvHnWi4H/XQZsYuoh8sslJw0CM8oWXKmE
UTr5sgBKVNp6/0wT1z3EGk1+Oqe11ZXrPf3uZGRc84q29wH6eiBqc3WTcZRh
YKdP6e+dSEArgv2kFb0qHRXYtIfNrh6D68dlfdTgZKTblwoL6nS0oaqQs2ns
A1L9HO8yMOPZeH8Z/ZQTpfaakkciDlVKpzIXDeVmklat+SflQ8MwP3Czleed
gpWYwcL5Xc/RZQJHrRAArSQshpg1L4yUnJTFLP4k0yT0fj1bTLTleVI72P81
I5QC+gOi17n/GecOS4I3Skptoavfd8g5giLykNtXxRQ3GO3wDEJOFithjLsM
+qoQ8X92CUg/kYQkZo6SjKGIXq9mzYhIfIHGeaJAHipxvd477AHCwBHLXCVV
ssuEFY/Jarz9HvfzKcSguieSxK1LWltqo3p+VoZwWq2jFfPOhEon8UbinIl1
ArQbYTpchypxo/BNKD2zzdbY+m93Qw5gSOcRwff+NMbmqpuSJB5hdO24S8CR
avHyUBCw4jsZ44r5jnG9ZpZS24XOnu1fYqquXmpuKRsQve7A0VUl/ZAQSEqr
eaUUNh0CqACUtwWl9CTq/iaVtC0nJ/IYDt916LDretwFuDSkaNWdPNHds/bx
xb/uSByR0UG5jYvcUCwcuc0OHLKvoEyzMKMcWMWh2kvQ1Gh/7BhiBtZrqbTZ
A++aZORi0t0waygGo2klc4m00uGI3/xym4l/uj9gKNunp5SFzMycHV/7kzaZ
qkD9h/voMV1SPhQJxVa373mqYo3fs9a6BfDKylz14T1sOYySqZZ7AORXAGbG
iJaRtPzEGpNiGTmaYnV2Sfh+9RiEuXbUnbC7VgHdxnpzOIpaBqx225WKGgL7
jWPDw6ZFKcuPk69hzhfgXqRB6PBzIFQX7yRUVDy+asqlAxGCNC4lJi3UVzyC
NoV3Wjt1yOWsjBTu0RcXKCUIRGKVfevn0nVusYmwhaAQAeSOfjPCNc2JZ+IB
eeIXgp7a8rlBKA48rBZHQGipiCHM9dEbNsyFJYghonY7x81bIEy6iGjbw2x2
Z0Cw92dE+9TKKGKbU2kPwGMingyhXzvDpYwrZAtj+ZC0gK/lNDH7+C1YILkC
9wafftsP/bodW1mK73KvveqTPchXjB5xF1+/4/slMafmgLBFCNPqqDILC0nN
Et4v2tXNqgLvF4wCFQW57xnDJwxzvhVJp0Cv2IB/Ztvlb/LvU84mz2Wl8iF2
OekMJkUpbbuhvGWWZcNINulUOO0X8b7KO+2UQVv1rGYHQn2R5gjbv0cF0/S5
T1uL+zgJXMIqRG+GatHzW3myZwInjae1t0xT44WBc05egIJhYgShNQ1tr9L/
QVnvmdoF5vPjC1o/I2FBQvKcKkukUaJXVdP9TioxG3BWekSoZWDWyCfQlJTX
Bd6DnDiYVjVMpY1QdANFTq8JLxOyMJfk8OiM5jC4y//ExGc7aq/MJlbKDLp3
0xXcLlQzfEXNdJSMaY+oL/rNwzEylh3gZTdbi27ctFiu3/7gqe8IZu9kWUod
cH8FpFoEhYbYxWY11zo7C/LOJAUpUKQILIHuxX0k67/OCRfinGS+fnZhr238
pwoTF9iPmh0BMJIO2ITGjwNj02NZfYY+RYayxQ2vTmjx9+R2k7tep+qX1riM
4rm1bUFSJjMaoMRE5FyTSZSXHQY1cp6Se7HS+n1U17JDz538M0Vu4mEPs+8B
ekyVf9ikkog3yNYbYyzB0S7fkXtah5eD+M8Ua3dHd0gkd93xLSqXNzqhGqvd
slMjg/NB3/QM2WwoFI3d0KP8PYVbL+2DgY+cORt4wmol/B7S8irtDQvpkt4r
kTv0XdrdKHCx6DbU+94qviQOhJRCYLfjRHsg7xFpwHdfMA9msRKM9BdUrIDZ
SP0BflRYBvJmaopF2CG5Hm6yO6BMBwkqm4oEvEMfnZETUFTz4ehy8lH3/KgL
6h9M2st+Gz9mP5RcA0l0FDPp4vZVzfpVn/f8mydXvYQw5p34UrGWzoG7TxH0
NWMptYShFna9m/OIInHdXTH5xWJFjP4lS0464QgLL/SGv86ulSoQUoRwIA5u
h9rXD0vYQilgMavjfjRyEaYwRRxDicz/IoIfxQJrQOGIPxZhIWtGOEaHnny4
nFyGp218o7ua4kM1uB0xWlBjA1stjukNeV5dINGkIsMaz1kEY5EC7xuVGc3U
HYRV+IayUSnEUoeOyVl4MKcCpPup50MXCMsXcypp8pm8Ma/zjGiaKnCkTpUk
Xupj6N7vYqapuv9iQ1QvXPqIN1l/mGPBOO3XZV16z+m06P83pBW6qT3YCjaQ
/FCaxzrFzNNNfbuA+nuhZQlXYEoNedLHJnqBMTUT+HO0G7qP6opYDyrMH9ue
d/VF2YMIYKYYOCusrkfc6CAtlQ5/ltMH/0PspRfNZ/U2SR6Z73CPDNUbEa/l
3tLSasiYbjPzqOGgttqoCoZUmpwQKxKhqYE9bXyQgvvK591vcYmCjoElPm0F
mPkhzYTj3lRbDZOgO6/UPf03o96k2Qo5fOZqN5Rhe6Tiog2veadGFGuqfUXh
CHr0kvcd1GTxvsHBv3QXrHGH3f9nmtix+IGtqw7WhxGy4aUf+bZf9JVNdpUD
V91WLRFl54owfpUmKhzkivuyEvQYXKFPclE0nolhiBN+RvAOkJPkCRstA6/a
ZOkp/snKonuA055aY7WR+LurEZc8DoHoAjmZiDz5+UBSOp0ogZb0VTCiwxsh
3L/C5gwBttc3JGMHWlx+FJAorBkH2DxSnumlEW1K6Kmn9x4VDbKb5Haf9HpS
vpC4O+dqaEBeAGAXE48QYWvyVixlltGUsNR90rjJmkXcIZYaKxs8PXbdrszL
VDewhXso4txv9Ni3wv+jBPNIh/D7EnZh35QjUGwBQM1aoFylEeEQ1GK6x3k6
O0SW9nBmTpYeU0+psl8My6UogJq2ghdPaCasAnmtpol46SkuUcMi9KImCi8D
h3amu9koHJvwfKzC3WBW/MlCDVT/z51qS/W8Zz4Y6PxAXKZJ+jg3w37ahmQG
nojDsUaRGMPXW7smJWwpTfADBcz7FQjDbC+zSKGIPMvCEZZjTN6QCIOTxG/A
Ob2EraOez3lzD3lUbjTG0XjrRCnkzvsqTye4wjLFqnLxli8Pr/YxyU8or1V3
gA2htV4/OBLL9LT/QRP9wGDLrdEdFdb+qOyUm4cmTxFUKFOVJ8ubgny7qVE3
9H/n1sRZDO+OfkcHjwNolYy7+8hx4KfjIp0uNS2Z4wlmJLB0USgdUmkilAKw
xtbm1PKkC8j/OtTdescU0J8FnWav1v79aktNboQSGZWRMHszWKZR+VJGFiIc
KfiOY6tMuiEFWUH8LEHuKrH1AXmvmm1gElC+62gupmDjqEoJztDDq6M5nMXX
bX7DVgZwe4B4nmc7mnFJ4QAcXNlogRuia3f8X5aZTy3OeyzSd7j8w3WOTOit
7Cx+3N7luwm/mSg/VwXw09839eaktguNU/T6jH1VjR4kp6SYOKCfWmPPliUj
l8KIdR6wMA1NsiQsPUg+aFH8JZ1DgyfWOG6jM16wuqVIOj/Gf+85/UvKLnjP
T8DA5nVBlt2177UvQOwooWFSPXZirxy3H06tH0jauatHaciEB3XJYwEyA/3q
Iecy4Pa8UNIC1/rgjpU0S0m7sBizrq6iocnwYx5y3djSxPyPDoP0s8+SzkCm
+26HnsN1yfLyP606Jm8NjaU98EEoHOe8BO+22ggli6IUc+O96WnBQhMzD9L9
rXKdF0aGypSpldiW1rYvoq1aR6XnZSlXJPA4p/2dwRX/8Br9nUmGWxfct+Y+
EY8wXc+DLGh2Tit3cK5UyyR1g1I6a1qnKC92NpEwZApuoWM2mrhWqLdNvFGi
69ow7l3cDoTWU+2BrhXdot+qXcgQpzV7x5cMw6nXQseTtoMoeIsfFCvUNAo8
g4SrLDotvxsZb3q4b2ouA5kH1XG4zxa1c0IarVheagmDU2ylsW/J2+3dCI9A
gLv6FbAHcTxJFcQ4C+wk67cOrcDEkK7cNjlA7oY2g7c4yhSHY9RwPwk3aX/h
Y8VjNvyXwrDVPWrQ826x50cvnHB4tzWGtBnpXrniUoYKlVS95K88tNXsAyxs
Ql+SpTTLMc1PtPcy4S8qwrJQEk0+MNIVeua289ymtSYPpyu14Y0P7J9Qt4NM
IKI1iiLDTyeixQ0On6fZtVOmJPzXRlJ1/pvBO5FwOIy8a34LMAgFm/X+1IvV
fm9jfZT5FBW9k6bq59GKBfXkEgfSP39jYoXRrwlDyYSb+5uc3xATtFmfesaY
FiHHlTRS2xEhOQPhYwAXC+NmODMSArUh0akRzrNeQxLdHbbJfj8TuDPzIww8
HwgSUtAnPfT5b9/cGg9kxG+Qq6Yx980VaQh+kRQrsxGawES+2W6J2kNGm84D
LMRGEAobLjiN5gVahtUly866rDYkHKd1+czHlA6e+UtATP8HHhPJZzTktbvB
zFwdN044wkpGh/AikYclEqK9YndWQGgMaHymJC40kaidhYt5/5iKIcxQ4W0t
gIhgdAW68B/iQgNyjebs8Q4hEHfsFYC7Eq58+8/wDiureSC3eJci0T1OkXIj
4afALeC+BYaVOPqLZAYqIaeoHBUgTTwDx94ShWzBCR04zmmFLle0ZeRtW4JU
CT0RkflQMxqC7kERtdBeBDcoHrAbwVz+a0lbMRtdTdUktd3sOP+z7e5NlhoY
rYkzqX7vcaJYcBAEQBfqDdkZ109mgtWdMwTArouVd0nWgMg6C5G6SUJ/4ptn
ZfCs+fRBp6/X75phgzddgivS3hpHu4vxghfc9mX6OyxKePAGTDVaiMx9ZfiR
LdiXL7kYm/GRR5WtaTvp4qcrD/5fmkK9PjQb5Gb26IUqg9F5GEvUsLiLYFPR
ue/Ecdrsrkoev6DKPv0wkAzstdUHQKKK+JAxnPkNk7ozLp5qfYOxR3jhSjWd
rmyT7Mk9mKcrCWbbB/7MXOps8qiWqy3soy25lOMbD3OFagkTLh0AtjWa1J6b
YXe3HESElx3WshUPM1usB3SKp9/ebHgL7sa1RvvMClTHbJmXi8AZ4K2JyLSD
xhQgBLfPUq8QdNpREPUxg6olht9jn28T395TcV3FjX6JPhDQasm0vKm2v5St
dsUE8Qewj772UFgBsuI+9ahVsojMB4Irn0CnnifvCRcRvki0Jsv5oH0buOrZ
GWpHjPSgXwVJt163Jp8PxcZckpLItqBETIkZ3/cpmPO56qw8cEplUHYt0xpe
awP6nAuD/HCLtS5YF8G532ulqT4gLxtAc2COiIo7s1WT9W9SVbmYmUOYJRMG
Gasb8jO8TYBySkCiR85zs4ar3B49HycSUFMKTltM6xFLP9GI49PcVUJ6MERT
uFYhWRqoSJ4jjcnr+gXCQbCpIybwGSyxBTt7g9RNl2B3/1Ae9lg4J5ggVVe/
KzC3qovYyc2JCTaintevZOZYVldt2oonFmUVC7X3ouhF4SweMOp7xxe8WzDy
V/heIsoPKye/ua/+BkvIszXQMyxMZwMoUgKMer7qxzL5pymz7TCGYAHJOP1z
mjHqD49CNYuihpX9N7f5HL/tk0wUliedyyKsJnMwXhBPVnQueL9zBd6ocS7C
vKkhN4NthOSKaKU4rG7HfogbtbsCycCcbOZu8kOXRtHKa0vIGjTXP938QRIi
0Wj6NAdlH/Dlc1e4BKUPLptM7sAIfdR6WEGHy5kF9ZI+Rav3j/oqQ7AcHBBr
qnFyB0cGyHHoanyCVD8x6YziTIp1F72s0pNUinOzyZZZkRF/AOxUkfGqQ0ao
43C2P+4pPGOjQ/b8OIFrDvzfx4/ZFYKk/WASsHiVJuGT70m7+lEXIyQImjyL
wdVTblQlS6gexUtFpFQB30f6ytmzi9inaafy4j+zsQi+KZZavYeDw3tTmhK4
9kDHnrV+zI2TwTD5PjREeNjNjD/iBLsA3nmNCoHgF7ZMU5VowfuY4gCVs9Tg
FbyM6C46DjWIKdBFaUdN24FqndFA0jLz+PFNvoEZKP7QsoPDkBBovlEnmezx
DPT7Qp9FnpkVIg00I3Uh70aE+zO6jDCyAjxvVMJTAbZpm1w0rdspxw+yqLhV
4M0TfvQXlynSqei4665TUjOXo2YZHB0NxSy2sNpxygoPFODoazT806CnrYOq
wH+EPFio4D+8l7B8papdlMVQPpNTRgtbYUl3aYuhzhiTJm+8BVi14b6N9GO4
ae+4kQSFIyktf4LxLe3R8bu06YRlkD30/P/HFdo+AMEdJhy0LVJS4mwETA9A
SMYtpH/u+/vUCsQ5Yu157p6G1tjdmAKSmv/karmbGs764cc7JduhCzeB6RtP
I5K84DYk8B+LmMlKXNdsqnvMqegTc8Zi6le/5Q9v2zzoS0EO/Zz/Gc6i9HZn
Tcpr9oBQ2414lmF5l/McUw6re1lFOo/QpMeV6N9iHB0h+A6AZCGO0nO13N20
JqESJzP66Czl+yfF1rM7EmIhgYdSf5QwJF4XdwOTQWPW/Zo1T/g63M/S+nSq
oK0gXKFvBEhFC0V6LOcHiUU7KpnD9BDfLGNc3/GJvaSqX1x7bPGhGNupKkMJ
0I56YZLbrhdQnsO2C6J43+wbmm0IzRqGeU31EfktBd989e5uExjRhITZHU6b
A+nh11teCmcSFr10I6B8pGzOYVJ7XakvvK9RDYpI9GAL0XHmqJJkMeDLQNIt
YL4NHQ1isdKL8VR5zpT6i12DlxFK4OwwXQrU0VjPxpcXvkMJHpwzGld+Ar+a
qWT63Wsi6dAFAXtIvSI7PoadXnWUfb3BXJDFKKkEggFk7BY2kiAxHXiYdZmP
1ZaZlF4xwnaAVWWFm8o36WyAZGJJ+Y9NG1oQpzrtlzevSTWLIac71pYvLjVi
fqI8NUoGnc07cf/gLEEYyM2QShUH7w6Xc+xS6zmFgXyHKri2dsQdEMMZezGm
NO1EMKri2ukANiHXsN7M2TfFdFwo+utD1iRNYgkM+5gM+8b2RX20n49JUMLl
tOHpgSLwZ5NBzGtNfLgwHh9RLGE7HHRki1OeVFp9Zvs40P8U83RcI/SVVXd5
rDSe8PW2bW1WjbOPiwjPWnAntirpbcWKqeR8j06mwE5iS9QuCrkmeBVnGqgB
9au0R5n6rIf2DAufULpDP+WJ3mMvPeAlIqOf5RpdvO81vIlwlRC95cIShy5A
0hzVG4RkwBudKesBFfl8mfnf7hfDSXBUbuSdo7oDsJ/dr8coJ+biWHtPAcg0
ksRCYkvoocHLo1JgfhP7YfBnf7UG5S3v+np96PK8syHBB4aA6FNUHLzbr0B4
9/IxTpmD38xSMJ67k20wgM5H/g4MgiVM4tqDMbVtOXGA7PcvwgP5BQM4vG8J
ZU7xsS7mRo+rzT03aM1LXZ/bHBdiNZkWGMe2IOexgFO5+SdTIFL/SZk6eXrq
/wLZL1Cl9Lb7Xp0cUQOp9ilXQaRRFl5Kf5ee8TPTe/SAwsBMZhYAnrgcvoEb
sDhDsEoOVe+VTxfnWwlMR6OmZ/X9TablQbCr1ZjkaBUQhgJ9CdI8YAtiEgn4
3sI6HTVC+GERXQ0zuVakrugUu17zfp93iA2z8tggkCvj20YEOdJwJi0Ukt3/
onP/MkgNUuCT/nmAhbK/DiUyEvKJ4DhykU6MbhkwEpW5bnhFgXRF19sWqRvG
+EN8XIRxmN6Mp2YAForwmGJaDRPSC8jm1vF+gDuNSkW+w6S50FxEQmkh0+HZ
2DeeBS/BDjmu8MDGUn5TMYazOOOTMrHtM22f59v1IqArBV3pn1vDVL86OM0H
cgSxUEUidWOSECcteA90NUtlwusG/gWAReltUQRA/v961+OQ+NLvmd3JuSNn
35izPjwEk42qqVxiY/z5VZSZqFzkjiu04zFY0b2qCi3o4ce3RFYecG248GfA
R3wfld2JfGWV2A53om6Svx2AxkNFmALxDbsTMpjHJep33QwvOymeIgT9B4YC
OTJICkoppT0fIIZlscEmauu+TC67pT8EhLZ7eW73OzU2HofDpD1gLApx9d6+
yKe5kUMNBza4221xFfgm7wFxIy7/ZdunbBhcAKzuqcHNTYgYBGlH223OIqoZ
Vqm2ksyY51XrHn12pivsJZnjWS+5FauJBSdI0O4IgTClPxzy+8lLBRWIQ+MV
QRgVh6/OY3cVaKMZpdd6m0fi9HQdOx5iQX0AVskuRzqKsDB8b7uaIuq0vVLl
VzXp3c8hbiEQ9QXTwmEWfnlJYoWH29fawGUKV/TnMtiFe30AzyO65fEQFZQ8
PzJlOxDByXueNXm3SJJCgZBFFAn1p9kte8d5FWvbXHPKxqYwYl60OEib9h58
5kvdzZtWOVtubF84cMzjQ224kRrgmThIkHRImkzI1LQYiYKEe7TgXMrUlH5s
/R5Y6uSAHTSkHKuBtQGDYDkbG1S/3E/gH0w2dszwKxWrfJV4+M8EYKQObsBZ
RAbP1wMxzmnKxUB84bN2elJBBMx/e1fOWfeotr9NewUgHJE2pYWVH/5xrfyk
YSuZwvL9OdjhMshbheHS3H1/9pcJKKwHjLBgs5LQFgD1EtLzyomqAWI7RfUM
Wmbnw+zJ9PdpzW+M957bfDhn1cvulkHsbHjVgRuUr8q7heb0NjnjLMl6DKYL
lS5qzv9YrgIS4REw5HWwHjH3rTKLt1uRmQxcU9vEQ3vH11WpIw7y7vFm40u4
DMV1ognMDeQ54mIHrBGzHb8BwvriS+oE3/OhLFywoOsg9Lx3gw9SOqxLwRPw
2em2KTLk3tOtamqYKfIlbNhbdki3cU28qhO4cH7FHJ0Px33yNysSXMRjc8OW
VwzRMdNU0Kp7UYmYSuoSkrdjb0dvIK1zFieSG93iKjD3GvH/qhCvvO47UGfK
ODishgsN02ISbq2fFLqZ8YyuOtNOY0hQWsLKmRtOaLZvNDWeSWwCPYiiQE3Q
KedsVGz+cNoU2Ve7Cy2vOtGleB4o9nDtpY/rkJemzY3oPGBcV6tF0sZwhgwj
wP83SISfZ7seGdOdPCK1CX4nhTEQEUyaZSppfEbvXvLYcbqD3ulRxvIUowOH
TgfugeEx38PTBzF5/fLNlPZ01zpdOCgLzGSrA2vyVJIOOqketQSw1yrbZPbY
Mny1NI8ji789t7cpXkXL8nzM9zqN1I4Q6KFBrKPyiIcbUkkJHlkg9SY9ogeJ
tDEbreaxCzczz4sCaDU5rXo/SEUQoBo0JW5NqiIlyXl5rltDJzkThlpS24t7
0Dhx1cH+srWV/YAqRFTpEwmdk0AxFg7ebGmXCgY5lAD7pihtwc87/tl+LqFs
7xlcFSiW2FMj11Iw/U4SgHi4kI2frMexLve/H1V+V9QU8dEZBNNLVCZG2J/k
lR8wVdz98nvRWJb9YGmIi0+ausdHkHJnQNvAH3h9WGG1EXh3Ehy3/tess3j/
aJBJrHx4M9fejCjcmkgItCi+u7S27MUKjLzanwcOe2Gt31J22Tile6iuOXlQ
iOiWiFVkGc1dfOh/GW20qSkqfk3MkRFgduHbMC0FfI6QZxUi553G9nKrE76B
lfoZxl4JdnwsEfvpRlQMBTyN53fcJH0/IEs1ZWGhe1pRmxvbKDqFW5qlE6Y5
7LjVLeArwcvQkWuMs4IxrpTPfZQ3eG4I+RTaByBpsbaAYNwjwT9/pEmOVzDs
8sRua3wz1jtLHb+FnTgM13zm+1pCIrEOEwOY3ZiJK0q3+LMUc9nNhKhTOLAb
RAzzHIVdlMJnMGMiw9T3ldqv3hO3hpVbpFXyyDUGc9iYR+cBnZLla8BGqag9
Gwkm8FOadSXZS9q40q2c2PR6jQWnS1Kf3sJc5gDqMhM7raxDakLNJPAv4czw
UCZz83lNr+OSAMvRRzQzPj4FlcCvQ11djTsE837fho3SZnCq5ajbH9Hq+Ost
uYQ/+JFys7xchI0kKp18vB1RoN47qGrovMt6MJ9PUS+kYyJaBAC7r7DBoUWp
2tud02Qa2KoVAvJ8/0ecyoceS34OMoz2ug6I7O7j8uiEduSN753M5rVNPq6h
ustg+Ug0T6/H93guQeAcblew2XuCQklFDBqPDt8vs22Jt2KaGV5ZfmevqTCQ
0MKWvr3yvoRe02RXy6t/to3TZNpRah4AS9K7gbJrQ+wVu0y/J7jJXpnxbXAG
+musGw38e/+tXLaN/Eefo4NFtZyLCsOvh7+gVD6GauVB9d7/wOC0rM4Jcw4n
L4f/DuQvzAcEu5efIZi0jkYuq185TuMEkpRkDtu2SF9Hort0t+rr8jbOZBu0
VIoOBA+CJgKIP1uaqLxkJOJkg2wS+9AHnlASi4V7lkmBeUgzv93Ghxq4SW4C
kD2695brJdTR//eFXxcgNiIDuptSVAjY46LBSypapuV8OtfM37xF4JiwTn60
JfVifYUcM4n2jausE3tBf4UmpB5wb95FcK/cOq+w2hIUoeB7jXQOaf25tFx+
6DqIPgbwBDAAcNZMI3X6iI378JFAwUjYck8UiDSMVjK+NIJmEIUMlhRPai8s
hV7VK2hfZCCtH/x8H3MF5b3v5prv2MuK6GKKtqrdoNr4IbhGSHkLGKIEPX3m
PNSFgXXKe0NsD9L686HLzkVZr4NRiiQhuVzkt/oVKSQeuLe8uNUZ4VXmEurU
F4sjxYT23VLBe2bVDYzCUinaYTeLh1KwaZ8Dzj6xAOXMXgVj8ntRJC2YfbCe
00pdO/Y99oRDF2/vWZADPJPBomx0lcuDkplHUjXgG/iftNGocMYy1scGlpQ6
ubtuhf/MKUjbZelm0xG13CqkeoM1pRbMIiolynHfq2n6m1H0Z4EBppuf61jU
0VnjZrPOUCPegcXnTFtplGfisAaBFH/h5uxrNthhCBYDiNeO/rwqZ9wVTtTf
ux69YAMUqXUZmBoLklZB7YR9+mjTZl7ANc7LAKmxYhjWS7m2ggkFyXGWZpOS
xFuwbqMgJvoWhpRXyiUamjodikrhSaHY8MbLRaTISWYyVEaCnsFJVGTyhvh8
xl0CG0zDlBIxWtfQ7ZLhWXmmfswpnQJPtXfTJFqAA9cXKFmgkD9DVy9sH81y
bMRPSt/aNycNWYC6I2Shn7vFxErw5zHvu960nscEzVweh7WpG3l3/q84AMNT
ITnvB6xffttbNQB7lHbftivByqE9m3GBW9Ru6bORmkhtvwbqac8FSlUQpMlH
EwhN30YhbrcZn+eOBZY8CcD/NYJFZj5mRDcqFPTSexBZAZV2iEI2I3y9qjyw
WJ7GjBDh7Tsm6BJK16Jp5Oic9yvHT/hmXRb5LS3LLf+Xhks6OO/qu9UUdZrQ
n1Ui4psXmC8TMNVeq6Y0p66nhzbq6UzK5hBQe+IZr3gfypbN9sv/M/qugvNO
B//raqpZtP2rnejfmTRC1MU3i//cGJozUn59eoMCm3TbKNLca3j2iheb9rEw
OfpOA2DyExr7yK3WDsD6Nze3GH/50CYI/o49KwQKKP5yEQCy3Yc8TfZw+C8B
uU+/ZqqUnyzE2dZxnvHDJnRcxsZMmMh9/5kSa2HuLRwxp1+Nvp0mXqAbvHXy
pPXDAnJtBXYfUSgkzzf3bSnfzFZWfvKeAfapWaer/x3+JBp/US30Qb0H3W+b
i30SdyEHvh/HyuTo0uwRXKQD32SHvgCnXtxKUJSAGpr6IwgJMvb00/VIVfYj
bLYgPFUhMhR5Bq9VjxDK+R8xrTMRD/ZURk+GeVQUf39aKcnSztTvVx0G+qjT
q8cM1MUlfseMPj9PtD9qHLuSAlaFdBMldGgkVb/Lgb8xxoNEYS9W9YS8MB+Q
CuxZ58VCW6pvYwbsS5RVhFpc6P7NCBY5ROv1fnJnaNg5qnUVHMxZgDj7KHPp
/MvT/gnbJJbUHfYbyz5GdBxzqfR6gdlnuRY8c6Mij49/gIwXImDFxUhr52N/
SWjllG/s6jwh8QMhD6pvSD1IwNwoMK6EC7kjoVe09siG0Xc7guoEe2o9z+48
8qvqcckMNjmGeoYWmVeWzLzjae4RHN991LMTHqPvDZG4j92xcFcD5DX4e5V8
giHl9XqChYO1yFotQ8i+PVf3iAF8uXci5fhJ+n/Bh1DtLc3vjjvfcYHEuhGd
JQiAhYDIQG7c7tWaALgydbUGKH1EENJhBNG5v8XvHACdCcp09I+l8t7SgP9D
Xs3sp3+8XieZZq7SggmBl1iUL6lNKouj+osxOY8iVYZfnF90aTRLtM0xlNVT
QPJ0d2uFhyjSctFSG3pDLGpx0iAUgds4M6DeXmOTiYApC8V1LSfwipBF3oB0
6I+txLzt72pwXh2tXDOgVXT+DfwVSpsudP9H5mUOe2dlYkWja3D5SdOBf+zS
kkG/vCWAPgv7oegtjQh8+5EAa95CQDIAEM8iiXiPzHi+q39uWdnXL9AeJvJ+
IPfEoz0/1UYbWtuslFvt7o2BNi3i8mhPti891X4zh9RYD+NR8/CjX8nmn4GX
/em+aZvEFQkmyaMkewQBdFxqG7cXgj1WRnFmru1MCTdr3JKyC8rrwzcQJSEu
oR8Cr4lUAR4FtEfQYjdlu+d15QYuNIE6zVMb3HG71XDJZ7bDuDHea4sElmtG
EHJiXu7P4WNa/FBi3eTC4hjZXbq3SNyEOyVohoeYi/88bzIKCZq0tzzzAk8x
qXyck6ced+n6S3iuVt9Lge6qMPRAluT0Ni+bJtMsXEw96hJZ/eRNF+mAJGDV
X1rHpJMuKUtG5R7u/ZD/b87S6u7iTL/yiaRks9Ks2/BcYfFQfrs9vzU7YG2O
tfs+/ha9u6+bbTHPXnygGO9Sd8ZHFCZbF0UjYp1eQrTQm0fEP0ptWcjzAvbN
Eq1ue2oFYPhxwkYyKVbt/V52ilruBJa8fSQAhnP1rg3fTkzFLaSeuZmSRq0N
Z9q4/d72LHiYQDVB01NB8Ud795MLY73BbnGmVbsfE+4Pm2BeJ6BbZenyyOan
ohG+6pgku2ehpmsijToX0/HRyNBrhnND0+V4kmMNNbtWuEGXNTCOr9Dq7agm
bYrqBgIl1w3tXFlzhdaFeqkl0xM+7MaZ8LsWSzOQvNZ/ENwhHfvR2DB9HDsd
7xy6uku7n0ZXrrAOeiHtNnWEiB8VxZS0s01dqw2sbXTnX6YRdmO3xb50NuN7
asq8SBnjkrxThW8xUI/nIp2/v8oTHuwnvi065NSzZB5f9tp9h89wGDpHQmzx
3XDlKtzkuELU+iDbOH2vrkCTPOKFL++VTbTGqNqoWxTuoiZxM5DAw383jT5l
JqnWfoQAJ0k4uxHeso3zlGo4AaJpOAMq+92CwFSkHO1/WkKZBC6xyje7cyIW
c/Nk/XS7KTDmpDJKJ9j2sVEVDkDVXCxOzZ+8l9lPv+wPRId21fARbN+VnJRG
u3qjYmilS7+PLu4wUXh7Bh+OKruTlxwdEJBwOSwor7Upvmk6cl8yJZujcMjH
CaeCvNsa67erWLHiFX9H3IYq81TagJ3ed/odQNlC0yFGE73Su7WRwGswBJHA
5Jiw8fo9G9vf8cpIu509FL+GgRnT27zIRhwcpdRXdSUpZ7qF4sGgBNSY+v4/
VwLUlS3vRzBn3stXDuW1zngnSIirXCkct0HltHn+srJNU/nXvEYKpQEyzr9n
Ii9xQZlibhYIleE6mUIl/9Ldi34MuGMtpYwAYpux8JBHy2xL0Prs3w58L7MS
IVcvHHDL1VPEWgswmUO+SIwh2VViVYnDG7DikGgV6dEh3S9bJuyNny1t/8Ee
uXJCnfUJUUS65pulbleuU/9wMA3If011Okp68lGinN8VpPc0R+/HO2Pvjk/o
oye8yNbFDlhMHqckaOlDpZRnYpo0jYAtUTV6WyZYg7frHrPRDEOs1RO5Qg5C
8Ls0E1RQDMwAKRC7AagINs5zLR4pZDQYGNgXB6Xamlt8Ogh+IqQMKeIWHuRh
3gtWzmJoGivAKPZLit2VeCkeign3l/7RiscMbZQ87GwfSa9F2ZCjNTiXEZ7E
+aZFeJ0qvYzPf+WXpz0d0s1tLLImtQbmRpyeh+xFo0gHOxwVRYZs2Q6dMgaG
Rz+dHmI5AXDL7YEY0AFNDrB3jmJTlLJ9iSDahCAmCHHehaGnVtU/hW15VYqc
8VKbDHMyBk9TtCoDstDQUfQnd28rsdOxBKbfj+ErEgRN3oo2TLxkuHp5jODc
EYEZztet6tzEi7A5DvklMdI4rJ1X4P0r/dI6yiWpQhiIHnRtovGAchdKr2D0
+ja16UZ4DXV50BUpjG3Mou1RNbF40uhG87Aw6+aSAXkmwqUI/kWe3vB9EUZc
tVz/3zv1hcW1qpMPGlsYH8dtepwseQx2hjCFO0sLtNdGWS16yMlKOu1u0H1D
Qf8RKyejtEcxUL8cE2UMHT/A3Z3Sr9uOL4mVsRkwh15gHsXALGgIR9G0brEA
sTkIDvolPnVRq4cIEH2ci4+QNvnsPtQr9kjHKmWFW2O5CjW1ZGZA6pnkosBY
GFp0HCvmlfwBe1Hvbl9W6HrMhhswPPbrILmw34dI9CEu9u7UNZELXqxz2IdN
/hLAQvCWD0Wvx9GDLpfcTd32LT1D7QrBDGHy1z/dWDkeJAZalD7DceGp9MZz
mhH3I/ZxPX+DU2fE7TqXWfx0u9/Be/Ve3T2rLYiga4nvkoU+BMIimUHt+leH
DGWwGA1fgrEvP+/ZDAn+ZMZN6j1crWhN1mScIBOkd96dodmCEoisrtYnapXW
BpGtWBvUmwsejnp4t6XXBeDhaKyGdEDRHJv792PsXrYaDkaKFSuW3iNNlHwe
pLZ5PWLtyDaPVSszpuWLhKhFW2JvsYWaMN6qqoJovrMorwqpEG0Qk8EuvYkC
cDxUUlaObTfDFeFjOabFPvfLMVCo0bjhogCTCz6Jn6eWvZiixg4IQYTyweO2
OTC/1hOhfimEY6n4i2a6KD+1BmH43NHGJnKXKEqC9cYbj0IM303f97o2Xmk2
5qoVunY+wlOdyxQeImZpp9Nh8uZJ2hcoyzGxt5dFEBcvcGMgvQuDJrSYMzil
VslYcYk4zLm6AkdV9nA8h2JrOufsByzew2Dq3cm3epE+hcwfq+6yS8Aac53e
ApGLgDu/Dmivaw4bffVMwGQiPCQkmhvV1P4Khc6/lijJS7D+0XpK1yKpMnBy
VZAHtZTNqdwFke3szaNymqU0eo85AfiRV6O3/Jhy/dtJvMTI3xqVHXISl7hg
vpuuGpJKrZL46EuGSu98EXF2DsUQToSs/Kp+g2gnnegrBM7qqa7SmCNucPwD
GVVLy8giielJspW9fCmLngi3q32tal37lDAJ0i9yjPTtja4zH25942Phopjw
hPSpUJyFv+M1FIdPUxZt84lcKqnE6+5Yxjd6W81m5PIV4pQDqPJ1k/I+0WzI
/pHwwSj5DuiNzbetfLnBJ983HXMg442bEbwqJA/rXzrCaiFZqfnOm7VWzJjt
43JY5M8WWDHF7uIUnXfSgFAl0HAq/OAcDEfh6ih/EDpVAZI8ZQQ3mKlQNhMc
BrdwKicXHhhtv4Bbw+eVFhOYllvrbcf5Fhlk7Zz+5R5OQk/k9jRrJ5SrOoyC
Bx7vJ0Uyy/NiROkSMqbn7MVWdMG/oPtIcbaBryqWfLbvKWRfx7gF5hpU5vGP
LHZYwzSuOdTaVyyRbuJzh4l8pzqWqmd61GGrzEc6J5OZBT5y1pXQWUhzTmpr
RCJbtSa8TTzTX6zsdRRuIiiAEe+R/dBDBgTjq1IVa615Uu8y5m6tidVBMICz
8RN03A+t9cDug3dIxFTudQcx6cmuk12B0ygtfNSlvpKGlJOAIhhEilIDS9Z8
n1g+4WOcPPrwKcNjzmMWdt4fxTythMSaZbYM/jO6x5SpdLZYgZO5zdjKkUg5
gvSd2G3poLFwx56PE5wy6Wbh/fQUUarY46GfonCiNkaOW/JpN+xkaTHdzx+z
LHuMZyfNXF+mLCw1RBOL7wOj7gnzVULt44ZHNHvHJ/MSS3VXzWs3jtLAKc13
smCdf38CbWfIDAR54etv73y0mFEjsnpiXFRBM1jliBbDB8m66BFhKYpAtyrR
/pidnzmBslUfXBXym8Emguf7B/SiLvmei66NAyKWD/GqpxbetzNczZlVbIvQ
hPyAkdtHmH8+S6Wapp2kYn58fQUipROm0HoFezts+VhaF5rYmaiuX6YxSOiY
bXqUKJueBlD3oaacTDWsfcb6nV9d+1bgyzloHV75uRWc711B8TYvwU3qJxWY
K1Y8nibO2lkVypK35mC75F11V+V4SIhjZXDgP2tx0lGBPoDPxtTUgeX6FFfT
GXV4Ige8ldqf+xws4UZgGUTpFOYx2qQ1I8XXKr/+CzOVItHWYJvik/jSAeQx
D6EqMFFYDgDdEmy/y+D9R+i2BgHn9hMlWT9943BLOpLgb/jUpLsqKBA0S3cL
WzOWjDHeFU6PW61VjajK1aqTm+GY6+5GZaTsm/gms091dEj551bKYVja81SJ
hXtdYrxHm8r11mKUNnkyCuYVMXbS4/v4VTWcvnlcEMQ+cIqj9f0pZ3LnSCla
IYA25hCFqAI6KVtsKWyTQAEr/7OT2kjy9sP0LNNHZ549GqyicYZxDhiqp7aK
qIWW6cJLSMgteffjGWNjgeHYKTSStfgMdvO9n0RqAmTm9FKfb1tdV71FS6nt
7HqfTvz8BXJtcmRfmcx5vcDErwaRPJrsV0e1maNPXMAd195eo8E93hec6PiY
w2tizrhJuHmIKkuK3XzJLvoisv2Rhj5n7bmw2aOPpr/tkfHG18oD07PvY79X
wmerfXO35XI9yfN1FfcS7BiShpKQaPffx6h2Fytl2a+hDwcAWZB7WHs8tW1m
v88be+Q3KuRpldoh9xuBnMZJ1FEz9fllFBCZwCLoNsKuj5l+0XGo4s68OaWQ
KJvE3JQ116cqWB0XEoyIceSgo7/k07jPG4v5tf9reD0WxmMDrusBp1dcKGET
8yZGwT63NQ8VPcaxxXexN7h1MHfeEZtTdq6qEpc2p84KUsU8V1h5+qGeg8Wz
Q4G6rYPlfJgdFDzbQ1x2LY6KxoIUxUdpqn4jyblw/T2RNtfjh03QWHte5noQ
yQx0N5GNUkO0rtFgLi9BTORearEHFmI5KVQp29likLzZVd/UYfQbpxKfkCCT
PSyO74Dsh5qdIInFCHcZRssX9ge9DZQrQgf22zUokhU13135Xzz+m3/eFKCf
yCZYq5wcZwQnmi0YOiLyLB6ET21FQywCEXzLuCjLjPrXtY2aN5VfVefOaym/
gJTIYEm3nVAroqh5BiMUuBdwiHLEoGMdGuWFQ7EsREUeaGWzc5qYNHegerP5
X7KpIlYkAEhxRnIOTtyaWqX6hJOwmfnbyDKbt+1TCXeiXjY1OLiDQHnshSlD
NrMLm0umkQ4tKci2eUYJqXan93P/bU+Ely9hY4pLOg2RHD/NxkmrpQlFt9AQ
mWqjOgCA1tdEogWuaXtVdGC/dAGkCV34T0kReAyl+KIAaURheUUsjsKuIy5g
h1YP5jgFDGBg1vH+Bqt5bZlrS/CJ8X3dPwyX7omEjgAPK7l/DbQVqXlO49Ow
+p2V+ImkoNEi4aM97fJzV0yJf/np7ss1yDYfv9NlKTtQTnkvf3nWK6aD9XMM
VrT776SNwU9JfEcoCCu6xXuprFbzxAYLzuTMPXAEfVx+ANImP982Zs9OgE3v
MtcVRx0mA7yigElntkxHsGm/Hh24r87BdMXZN+ILnlzHC8I0EvfshTohMV4n
4cXZHctvS3Ie3R1R/2OKeo9wNeSTDyiL4WiCN8jgc4cIcF2+3CQ/TQ+ROC+B
K5TspNz6j6dMpqTOIcMom/fCl4Dnefw6PtuITrjnM8lb4HDudmnU2EX7b5hY
ven70AMp8vlYNEqwYw0OrVPZH54UfCsTgybEWGeFg3/ALxQG1qsml+MwoR7g
7c+dtBnKJr3Jm93Ntj6Rpdz/iqy742Mjb63lWoM85nfjpFpMDkMDJORb/REl
eN+27j3Vwnj8gpfMe073YBiLnFXV50KHrSxzPJ5As4dxhqBJvlAgibA8o5CZ
h71Wl0nVtJJFELcL4AJIF1uULzB1X+naAZ5r1+lALNzGU4m+pPRQQrOXoq1N
kTEdkSde1Gg1VEPg6jgh+friKoh1eGL+21wW9JERmvZ+wH1yijpwdpJhW091
k47bDFI2F5NxXy5igMJnaY1+YDlQ2fWwvNyNyjCnp1K9HUBSbQp3nSGxSL6y
8ucbQ9yqD/HcdZYkdamhYvB0fWFqU1LlzMvF8ecEAa4auZYmbWERKGGkBO9d
bx7pSME7NZ2W3go3rEdx5IZOB75Z9yyFi9lFHLWKIGDEvQpDT6HJfC0Naw9d
u/xbyXNH79GgnziAAlSiscKPMnhkSAFsd5ijqT6DHieZ79U51iG5e8MQKVnH
0fhl+rBq1q2zwzwOSolEPr48brD9p4z1X0lvr0zt0IrA09H3iJQ+KS2/KVWO
8n2YAovU/E2Fr1UV9GMvmeSO4TcGGuS6bZCf78fENKijOONeOCGzW+OoQF9A
YqIj/IYzk4mR6raiAkSPndAx1VA61ArvZ6aiCLhWkaoLcmobWY6u8iP/ZxQz
Xuzj7ZTmDt4IJsVsCr3AEWfRr18H7iqtLDln+9WaJbippGFypfSmw6R6ZQux
AedSqpCx2vDivmyyUooDatnzjTlmeS4RdOwVP6NvxRLEISoSVwMUzz0MWGic
xTOYW8o4PGuhdSsJuzgFFWNF0fEiAVti9nZb5JgnIxwVEBLrQGfrQu8KSp3c
dWDf/PcIzfV66XpUFc/SV2mvpFJLRHc4rRe2Y4QnHP0UIzClVGzRYdm5tYq/
sIY9Yk8n+IBghrS1EPGngyeLxKgn3RQUH5z9krzByQJKqteLqllGcJE+fV/f
mn2yjJPuNsU3UVfPRcVxj0jn/H9iqwIVDrECzCNde4yDYflfG44yvaFbJUP/
17e6Cinm6G4+AgdootXlQPV6z/6T7tVfazxJhzLmfBbG2zdFuXtlpdLNpNgC
o35OtFcQkmTjgOaI70oUEF4AJbgcCN44rmFbSq7qfgRyD5yMEe52oamC9eVi
eEEQ3aRx7PCdgaamBYKY/NX90db+NR/U56sUMYwf6GlliFD8YS+WJ+zIrT+n
v8wrHPlzKcBCvRdy4MvENJh2B+itRVnQsmz2djTVunSpy8ECe9XcZczHqBvp
Phjr//A6Y6kQpxRyeTSDEsia2060RQF2OQf6GpmS1VXvi7NnZhq3d3xDrYVg
zUzQ9fPk2T26C9XoJaV5wGXsHAei+mOCaVd8Mz/KvQzUGUSsULeos/WMGIs0
f5alD0h8ZT8UselHdYzO0jTyrdud0pe2AqXReOayucEuGS8irDDkfNWERHNl
rlkzN/Va4SlblwL+nQma3AIotDu11P7NycvO/jYM26eyHhtTjQVHCQt8Nhdi
r6BOmfP4r4NlfBEskOe6LJu0gnOy7r721hvoNlcvXVwipJw3NIZ25ROWgml4
WRkjGN8u3p6T7GYAhYlYpJHoORW/m6+VoAZvpux71bAcVEfMGwnmYOB+uC5+
Qpjw3SSPc91qeBEK90c1vmS/wSTf5akUFY4ybEv11+6eRtBfTmo2SR9DNLcf
SYH6cTaxTCw9NqVnic/qdFTONHxJ/97WpQ5RDpuxFSnaKQMuhrb9cGbcA6My
Zp8HhZg29imbzLTI4kGd0VSlb6I+fhc9uctbm6ArOAHRoznLelN9AW26rbML
BhXgA2aQNm6zLBqmdj4U7UatjtRp0Q9kyuDIyH8ZHXJZRqS9yr0+KXMZQu56
r3QMC9ACjTSPZRJjoyOOjCmaZVK6Mqik3L2Kmno3T8bdqO0B3YiYHvLfxVQW
fiqlV2LSIhTb7XOGWPgNaCY1iYv06lgU9IGmygzUKCBCt4rSLAy63NWpjHNH
ARADJ2y1ZUPB7Lj2jFrclf2XAHp328KSaT5aXw+NfO1/wnkSEoh/fwUfGs7C
YS5Kd0GtbpxeSViBiCqIdwkyFz5MvE5Yeh0zuEQjv/WaH+Uq2sWMSTO8I00C
BgxPjTrym0h3r724/wWw/Y8kvpk/NmbVz9caEN9KyIBN0W5FJsE4LWK5WIQd
fYIH35hmzZm+/C0o6rOBF2obXkbrsNZ3+TtY9Ni3QTDhlbzztDiYKfFrPDlj
Su8exb1nYbIVtyWhtslGH3u5OYC0WBErR6x4EQxi9p2Y1vbwyApajNOICl3t
lfqRLvaU1ieMmBh0cXzSihCKprQMOOId5VokRVxOoseQR/tey0zFy8SKSvMl
ospBxN9SB9o7iKy3fwibd1ahmgPm7+LjC3q/I7Bts1StmxJ/8A6tjlTAchx0
KBFSX2l5mUYnhB1g9s6p0Pr9Zvld9OLV0Y1ODh0uhfCXwhv4aw1J/orj+zZj
V73eYHB7JQU5mzLuifv94MCgn5+Hzk9Vk1RhAKtQMKoOWDbCDzp2AukWuNBF
9/03MwxaOAB+MLR3Q7BZ839geqJqrBeljwLG1y6xIFs3NzOHjffLFXn8Olxo
CrgEklvWEII6IvihXTHHh429WY/Y0HxkeyoZYChvGJfEjDdwOfDlUieTQKMe
syDA1IC3abxpIemD8pTUGMfnG9uJLpzKH6/3RCKDtlA1YcZpIcAibN7oHNkD
WjvRqQW4tenwBu6uqYniudmsu2/kHS84Qz4CCbsSs85oATJsbbUtPoL5wbS9
7ccI0d7IZcJp8FOcFDdB4UXpyTSpQy1haRO2GlkksdThFhFXhQddOs/LLIgs
Pq79m9Br/J1Jw9jnSyb/dzP62t+E6VcTPAIEXEcjQV5GHpAysHSDnB2T5vtO
rKkimdFBkzaGBqL6LdrB2V+s9qePMIjHpqu0xIqY5LmR4BD92+AjG+f4rFWb
Ah1aRzvcJOdfzvZxiA2nFBNXtniCEK/R8G+Kh3pF06ccuS7z+NI+6D698jwb
Z9uQbry9YwYdjSb2fHEGHWgfyXkBElrg25GOytz5WozKfdR65Mo+qX4rj+3M
QBmHLvc+WPWwiNvnDYNWOmGeTZ8+BmykKshJmnzaWU6SxLLiYlpAr0TsxO49
CSHCbw2n8iSvAb6faDUw4/wCHrGmt4nFky+67vCUzAlQpbEA1YxvJuQ8WApE
KnezCKiDLo/f1ckFh/w5rAbxzFUGoXWJ0SvKtSie2Y92dtdq834hQiPtw0uj
PqrtZjo433wKtLbSZXu4aA4t112ALGi2y1a0Ef1pD4TbToFQFI4ewOv0hLua
0sSRfs0Fn03OM3GhJ2ERGqr2z2yvfHbIzcbmgsPOqJPr4n42K6G7RJWIn2ve
gtjeILIhCeWX+yefOKcvPKwDMAemaZiB1AhjJYFD8D+7SpTmwSgZ0mRFb+D0
tqy76NuH7YJMBVXEwCf0b3I69HXRpihuudRoP9aPdXEywUFHebv17lh8Q19D
DphEdlwVvQANooIo+ziVmcnprht+B0UTqCo87e9DhLcqJNsRacoq8cDZpAej
ls81XGDqo7XwHjG8pLR6KF4iBeWqDSYgKoPfcaSxgP+HhKupPsFZfADofRsy
TjSVMFvDC4dA0dt4yybh1G2XuutG3rSCHbVwmWM5QcHmFqCBi3zryD+h//LH
dFlVDGj+a9z5Qp77KLcx+Dli2n/VLDh7MmLt713XMxlk5BER8bGMQ8RzIHzX
Hm5xIrVtqMihsb2B9SWQ/gjzczh2bcs7lOZMdD/lBR8IYVBcaflPrFpIH2Sf
Txa92NQqKGL+lRKPw76XiN7XONJi9eAk4ghZy3vkgc999y4uap6Rlbnym8tk
Xyj8Xhf0evRPznQjb+G6r40Dgvb2CS8CmhnzWl8Wu1I+ciwtu8U8M8sSV/sD
CeyuRUUMzGFvFzVzzdJRu85xLRFJCbY3JML9jACPTQMPhVKTPp0bvRAixUh/
RV4T6upT6Kl3fOpPTd2D8RKGDuDnk14sZd6ipkSi9oeeZuWgl/LWVoXQfCQ0
KZ6Y4RP+C4elX8bsv3Vfq7T4jX7zaBpz0KV3chkfq7A8bXNOZZI9bHEaB5z7
P1/7N2oWILECpi++SnuwzAJKFn9srYuwFjAaouQxZwM00WjXMEYDnrOmMCi/
n+M95tDEawJAR4DRMGfvYrji0a5erx/40tykj/Kn7K1v9NhHsM61SKMdogQY
rQmjOOluqr5s0lGPBMuzxhMhTJkul6ROZ1vTP0QuNqbpG3J2vtA1BMGyM9dG
JXKJqwd2OEcfr48BqEhnd3C5KQ6U0OvopPau1macVPvwM1IEnMfssWRg5N8R
SpZXdbw/YcnUBiDC2+Y60eI2a4+Osws0j5h25WiHBRciHWzTR3w6z5MumhCB
klIsEpaSE1Us6aYIdrQSuw/eK6zplDfcNqh8xJOd/I3KBo1Ouc/4s3UVr7ql
3D1ELDsHOMsEcmdcrhBLvYvMW533nM23HR5dUMXY9zKXXTaELlo3E0egFLgP
GqjhsfHBRN9fP0z+RUf+F14tsBD8Sw43SooP+zm7xooMnz9lejgY+JMP7NyS
xb4HoeNeHs4+uSYHwQhy03/tsFuBOyHkL556L+6z0bg2mvTL1Z0a9Yhgd+HC
mAOglT1nOgyisAwPq3fwPHubKwtTEmcB/Ar/tPSwX3g+p7iWTxcVuIsf/Fla
7IFNfjf1bMqP/16KFhLbNVC/bOezoENFvWMQiIsGVecHAJg2Ne8GQF9JBlCz
y1WwKDonFSXeeE3IxW3yvxMdj1woQWsu/R/136A2pc8mn9HRcZt/GTHXUDAg
ApzvZI0lQD8lgNU+0RPzqVIHAD53GuVHZ47XJyqJ37Ja2ZS7r4+RqrA09O55
M38tk6MFxwMIHg8WDA+4KfpiSRG7jRHQdC9dvEjcb9FizD0JkWO9dvi5ICQD
JttAChOQoAW1BmlZzhrypv6O5SrPpe3c6rvM7W1Qfmc6184ucrJVq5VUVz/3
PbpIAZEvNxBQUUn5saNeRuxGlPx3V4z46pF7zyzVXiSNm4GqXaHY5ZXbvNam
svOMls2ESw4O4bVjMzOvbnDi45vAEdwpTRquE2ZaLIB/77k+F76a+q8P6ZjH
6HZmeGlBplcfQz95/16jwH9efZkx3i56y8jhMc8OzsU5HbqiEKgHl7dnkPjw
1HXe3k4dXHMlrR2j7jriSN7MfCzE+TSjRzKOXXcIDX5/02jqCFDiaZAnxsq0
+r8l3IgYmKB8b12NzgXaQMRt9HHzxFo2OQHDFmYqfOYxGCI7di+eSpN6JsOL
64Q946xJMlarNwRWADRmeYI4ShRfX1uWMMsGah4TLOYdRSvCXdQw5mtvMOEj
ClkodEsjf6xWDkhkvKHJ2XLHwNaHK5FxAnZwAj+hZPsIrHPjWG92612qH+P9
nkG0oC9Gp3S2s5LiTjd7CXdxUg7Rwwy3kGJinbiX2QNNZXilXeqoDgCvuXrq
b+55Tdkpc//BKfbkMjsmoRmA9mEqxz3MVtL1grBdvWvJo/vcYOoj2KToIWT8
vLNjvIzYcpvWsDqULFeA7M3DhQmBAakK2fPk3NgcDJpOlSlNkn2uG83l/SBi
6g6LZj78iAl2riBalSAk8eiLL0RF9SrlpA1ZWxHd52r+xecXaIB4CiyxKO9F
XIS3LnLuKU2H6jQMnxTPdsqN6kpsIHsrtvYzRVbhzffJoGDqMDOKMGI3t0BT
1T6UjdcXz+eQeFFEuYW/1+9cSALUJKkiCKFf9yKk9Z6C8yud45UBoQr5a0Rs
W/z1S9M0HTg5D5Cet91I6msYkBL51Xgqy0rYfLnl2o4F5vYx34L/4y4bCvj3
QXEN+UCKf62P7z1D+Zwfhc1Uuz+eJFLeNLQVvAu14cvSDtldWwLzxQjN/nLH
fIuelqWWbAyyIZf9PQDFDkCPdIkvObK17x0XmTiHHxUfssrPN/PNcGNKTfBz
Ev6NNlvyCK9bOw0ZPMXrcN+/KQXAh+kcbKFpnA2Fq6w+g+w96nFIi4FuJz8i
b5jrOvkUiPTasf2vzVey24fZT5EMmBV654oCOi7NgmAAHPp3HbMuia0tDyQ9
tR7DM/D0vFfGJAPhD9Ygu5raGiZVY/VvHul16DE4przwPPyPLaCelEr/DcF4
OzDv+bjcpOvYJxKSpkSloVOgUN+HxFVTrcRCKG9Mk3xXN3ygikt67r9tU8u5
fWZILC9+xbsYX41M9lcD5CVaioq5Whchz3+3PZnN8yuv2iByj8opch38XJfM
gXp9D9oLJnnn+magih4cd2/Bdz589h9qUZH9v83SPZ3GZ54rueDOvCstz78g
gVDBQ5wkbVizkhTlYL6IFcUzpnnAGWTHxqXN8CSswbCHoEFfFQ8JqVbb/xfv
cBpPkQIZbST4vUO/b/QlrQTMi0M8tWY8CrHpISdlIBbzhTqFwSHVJHWu0wy8
jA+Cerlo6l7Rhc1EO0RFBZnqnp7V8KoxpDxHz+oi8KqsG5tJj0EqxQeKsZji
P7SEWz3u/ZOzCadoFzEGn8iVa67QoZNO+1BvhP4nT4tUu19+Imj7S8ydO3o5
DNGDvgUkFvjU/kezaIohhv/HsCxR2aQ0i/NdyKIIg5D3WhBTv+CB7ujDUiQs
l/CdrZ36LU6gbKtJiklArcOjn8hk4TtOz2Il07Z/U2wz6BV6A2tiNF49MW12
5aPYCOyiGepah0hFtNN8bQKeKGMZ+lPl72sPlWVbJiwQzEpOaEyclZ8OQCkg
sD3fB33utteITMEZbBZJfLQbrlo2S3IygSSeo6dP8/Ssyia+6lfo1h1YVTqC
+V2qPqm9nNwV4AziRdtojhf2i48eIuOgkhi+e8TUUNjhAB8JT3SN6oyh4IhA
gaFLTtgvHKmsxdOOAp51thUzXseDI8gCjRMIGare0fNdFmR9cU3NTfA+zYLk
fmSoDVF4nOeGZ5LpvfmpaDhPY1IjDh9aMQ4aW8vv6RF5nzbKz6YnfrL/xy1V
54fcUdLTzqtsXESC1ae67mh8xPcZy5iPUiaVX7mOuul3Vpc/o2hOwBtjYtI+
3PD0CXXZweuSqUQwgD4TlOMpHzW2gCdLzNaAJlKlA/R9FOb1Cq0D7V2y4nwl
ZVuUbeGRervl33QRCzk/x2Rs1DbiKRJHL9QPy0J4BCVIvu4cj58cB3Mqamcw
LAYZuK74HnhTtYDSX+SeGCCFmDbEntFPDUQzJS8n0iMrW+ZfD4MBC8DrDX2P
YaOhUJztXI7EYH6SjumRIlMI/qaZxg3wzSInYUcQ7JlPs9LaqF7fCedstZII
RuGITWH196m/I3QBnM9dn6IAz1HoMKR8+yJeyxFkxDP/9ZuKt5dlct0qtbtz
5X5oSW3MK8Xf9kMezidtmri5pw0NLL8Ok1UEsCGmaH2VqRgxNtU4akkjIg9c
I8bZ89lr3LpE1/KcPr8xhAySgjAaePN9RKECfywdS+JZQnVh+N71TU2mQ1AT
UzA7oaANMlS0V8qG3rP8zKEKZpAizL/cNLmZ1AvsbGA+84o4vb4wgqTRC/yY
c5d+XyZk7zaaQ1VIy2hKzilLZbvfm5Amlt/Zde7FmPI6SX7cCAh25IYd0fFz
5zU1lRan0jM3V4ZPSi6pr+RX+zZbqodwQmNZvZ6X3UgGvqtMA3Es5rcrfew9
cjwFr4U7I7JzOgne2ZXKCjLLOCMfZJFdx4AWS4Qhdwd4Iwc0fL1qVb8e3Wgh
qW+9Hhjl9607ovHPpWn3r0AU75ysSWt3QJD71e9Ck7qFod98VwASsDtWNqo9
h48DpfDc5mMEOUpoxhhWP/c69jEKdSDQyPKjEfm/8y5XE97yau70WfE8kDVJ
lYFXtC1kVijzTHwC+bjNUghM3MkWuD9VK1edr/+tyxa79ku7SZBgJjZvmFBh
zj9GvHHm2fl7uAr4hvPxT2tAoS4KlsdnAbkFJkrQriWrjXYIimWwpRh31GW8
E4ctvATfITx6eqUflAQd7TdfDl6gK2iH9UfT2eIt0qEbXiLdAr3MTYvtluqA
mEPrH7DoJYIGXXQxzojr6NQG6ffKpeB0aY5F4Ac38S7dFUNY13qamSzbwUxk
BkiWUVNSa7diISXbBs75SAnIJRJCFqNaHFxSXtyZ1yZ+z7LlYf1xb8/6b8h/
3A7wX80Ao2D3BYwvugPrkAX/5N9T6/I8e3pkhjs2IbfNfEIGy1ekBq3zBHPT
oBrql22UHj/kkuLU0tVQCzlSJNjx0RQJMyAPlaGX1cVRQXla+9/kYJ9nQuJi
S5DMvRHJpz2AVyyg3jgy9iAZ4HR5k/3IV62DD73oZEP7s87nEwbG15lXTnZ3
DsyMkWcu/5ssZt5YU/yMc2z4mwHEmeDu/RPP13JLu5b2i7ZDQRToiMnraK10
P62fSBP1xepQl4VkfkxMEI97wr2zE80cBvh/7RUS/QtZGIVnQ3rPRf3aodUV
+4fCzAeFy0XaU0HJXRWeVUOonhBaePL6Vy3MJvK/HJw+PQ+Fv7f7nGD6ZDKV
RiPuW3sdG0Ho3U1BQtAk8HmcTs6fGi32lKiVlTnBSKmZQ4aCJZmAR0dll6rj
j6bfi9y8sxM6+z+hO+uKM2ZZdQaf0+DOfR+0yjn5JLdwpcG3S+jLimbjy4WC
M9muEXesPTian70pkCZS5UpXCJpt4CtFEC4y1oVZqxkRcV3qLZbwVHZ14+/+
X0x8k2eWYKbb8Jg7GKYDlE3U2AoqhS1zjvRxfYEwFPN0xCVPGwGyUroPo2MP
8aw0nMUHX7pi7hO3jjMrXJG6SKYOG0Ykk/umU/0oHrLYKmxFmFLIKAfwNNkM
tSm7zkh9j429Uvhjlhoihv2ED1E8PEqNqmkUrBUZWLyYZnY37ksghEJSrUfj
gWvIOBeIMDDavRmhWLyWK3DcU0kcIs38IX7p13s6i9aMRrYCb5oSGflZvIl4
Og+fBrm179DrVeo50mpS5ylAqlBFnDjesLh0gWGRy0F/QFlr/qG8MkvCn7av
ykjfS72HCLN0X0vuLV6HFjWgfKvAU5XTH6dJr2sISWxJoPsQ+XYAPh77KDMl
otrdpHtcWsrZaz4hvnBMIuDjjZTsUKkUiB8L4l5+LSb/m1K/I5X/y2n03r6i
4q4nEjP60IkXdrrnUYr6BT47aOxu4/x69T+JvOHENQCpuyOxIW1+hUAWtx0r
w3hP/l3gwHlP3z35TEBpdk/neSc5tMd4VaDI28kqfrARHIVcxhvickXJHJzq
KFx5JNxdBT6/eV4K3D8yThYI0tQVKkorO/79iGgVWMVdl3Q+letFbzoq4GbK
YZIciBYprm9VU5r1NiVuMRjv9x7E4pvtne0OiR2CSORLb4O5sV++KqULq9ZV
8aHIcb8HwOdnD9e+EsXpw3SX8cqZdsvEYOQdOF57+0F9RHH57yax7DDbnbNS
xHV26u5gkLFw+s6Ikp3QxhWVAgueARx5y/pkXISpZ43ACNY/9l7RkvaE2s2d
A/LZYEbmiJXYZxXqZK6tiyfcg7hrqfrTDv6efP0b252mYlHBkTIIkc8r0djM
TgJjI5URJeeiqJZ8VckHbkkFgeKVU/G1FjaogXW7Z+H51OCTYuf9YahMo6wT
dUZ2VWmDnDZTsyOKz3dml0O+qV6ytrVAKv0o4YFCizrL1pxY0bi1dFCHlkmz
uBbD8LO+sImBvGmzS7yIBz9d3HOktN6+I4TxYLIqWE7NwqCfIgFWmsxG+ENo
I9qs5yiaNiftj8aAqF3GGJiuqPeHL7wo3ZmGOnnBKlY1NjWY+KsafVzLZOVV
eVObmB72wGCPibSYWNGS7WWumYPPqYVOCw4SrQB3RDu2GS3CLYZ07NYNj0qL
BnZ9+3mNHjS2/yZbSKxqlpzU/bDAB2MBeiSdermOpwIn/DAnpSFSoTgyGWWZ
f2izgnJHguXDR4GIoIYpTP1+bslhxIW8ukm5AWnEzwO4rICQF0gGZKE3f2PN
G8XIvhuEoj3bYyj3Hzh1BGpeTy/v/b2YBCORs7ZETkiUHthAYlUArNOWNQ8F
DXLweUqMRcjOhK7NeXaBpWOgtAd6E4bqCy1N/4eYy7VA18Lv74ZlZFmie70y
Gz6wA/9mh6eXuZ/838QyXgeiU5pdf4XmAlS8bBLCGczBNBuTn/L51GpZQhKn
4l0VE8vLjM3g/IyK8MaWm3rjieJp1lqKm48frXX3v9rSw1/dtY0KSFTdPnqn
4F1U5ZLaply1EMP7Wj3YLRrPGBHPPO93rslu5vAIfyEzGJiBtDcDaXgw8iwu
yWo/ad3699yxl9EPGFsqXE7Ez5GVTGWgj4IKXSnWBJJMQ9q9do2XJjq4x0a0
aszs03itOEBNVBpmdBnvExxIkr8ZWH3PxbEHLZCvpIwsQI6eNy9FhTwLjwfh
XaUoJE6lvJDNFJhtDpD2vx5IA0cr49I3nVtx5gDDz6kVSbcj1Xq2JapgsGfh
xxwJAwyVWBWMOY2sy0tQtg+PHQX6Xn05dKTopVT+9uIs9hckpyoxvUZdAHnL
9T211+PiwJfqo8mV7W/bRGUY8t8K+AaD73umgHnKIQvNb+sdL77GplGm8xyI
26ug4QrlAA8/ZWC3GaYQBAJqEf5JLgGP49wpFfWVbigJS0P8XhStDqR15Omt
2fqE3vfUls9psjJC0jwJn9cZdiR2FDmRw3QYG+358EzD4VRxwE4fWZcpSaA3
nuSzXUzQ5C/WAFzCzA76FHMOjcOIVNlLZJIkczu8C8iMovcYEs60KIA2FG1X
aH797xH1LlLDbgY0oEP56YERUO0/frqz9N9jgX2ebET+E7J4/zv/R9v4Qeyd
gmaTCS/gZizU2IC3CJ94CeExRNDAtg37dwFM+8f8eDRiacHptdbnnXPYUkvU
DYhMpz5vjILW4me7ijbTFbUvhazyadsDdeWC8d09iMSn/iVm7kJJQ9M1Tc+2
i/WwPuP316Vo0ZItRYqxEEUPBlKeq8fe0X7Zr6p/oaw8xDL7xf4eaezt1wsR
R4ku4ZWBLzFh7P3hXXOBptP62Pgb4S8XMfkOdmHipmhnsf83OLRXYrutj11C
zr2fhq+vaGFvnNKH+8dxb406Nrx62zsvYfPm91rCRLy/ct0USkyuKgCYfGbG
66dApiKXthxUFI/tX5NsT7Hkjk8Rbeb6y05TWrUhjeaDlYPXUPX/IDqNPA7U
kE25kMkSWBEULF1fhhuLxWOdg5rW0Y2oshLentM6QgYRuEDS/PvRMJ51Dyzm
iwYBIH/CyWxPNp6TICLS1g26IxTDJQa/24nwJ1wVxatf/LnvGE+LVwkP1XjS
9O+P4iWzQZw18pOveWgX1TCa2vFWWko8lzBdCpBXeHeE+s/HlZtcrwjzr0LL
fjhJONDqYZEN54387WZLiFOqf3Enr5DUogYMCw/De4BtgHmA7RuPMMTlPLOM
Q7ZIKyM3QwmWHqUW5nAp/DxiWfgtClesjvDVd1NQ04SQYTM9jRKcwUd2Vrsr
/RdJ18jUSzD686fBFpRieQkiiVE7GHYBNy3n41RqJhRvUszfDzm/LU47bRbh
ZKUjnOp8f+cceNYUiv9hYHfBKwmLFB4yMGiBjv3n9ZZLN75dXP48P/DcAVhx
odsHtN92lMFBUYjocAL5QLUCp41YvlXVuR6BTEw89ZYAxt3NSV7ByufCFEth
WmhUPkiEmDTTzGbkr2aeFCMfjarClvQSA27O8DddkDPQfQUGajRzfJzqYQ5v
EJhPb3DOahRRCcgrwAiq+CiK6MeBceUKeL/BXK3WaUavmv/UtFGHZH5M16p1
wdEQ/TdX0JuH3DpVSY9+LpPgut8s7nr2XILBOuAsWyGfefZwQOP2XfS0poyQ
nQWtUgNX1SEGRavavCJO7rV7MbbQxg+tnaJHwKFsk0DoziNO8d4ducIBthIC
Axd+aHYA1RsmQNDbr6Ga8fiLiEPpeJZVwYqmSjIac+JQvw2txLoGIZjxweMH
/13zwxKw73ozRi6iuOfp6EazMqe1NVjcOkeQYYaR7KfY3r6YBgVvBIIHkAU3
V0k3jjlAzfmQt5EBtYwDAPxj7icu80ccKqFsprDhIgTUosU+HVFvabzvAC3n
hkIh7uoV9h45lWyqGu4boBVo0PBajXZg0Hajfa2P+yG8+wfFPYGiozmg/DT2
OU8Bqd7uSpXvCsQnPXqZyUKkB6vIfPwO5oQEQEbvXhUFP4ryvAn/+5YItJNU
yIj8BBxed7uWiPRTF52IyoT7lS4RbGp5mtqJm7KPgb7GeBQDwPXUhSgW2zyv
0KvvGiR6JzK2N03f9OYz48MsJfoofnt7EoGEf/NbORQRjAvDz4zOeBzeYN27
podk+NhbEeO8qIc6d82XYuelLWVjaLdJrSqxT/vukwrOYKaWehdM3Rz/KrOm
bgA+g5GdsAK/owQYdqefw3beD1mmzGKutK6gRYEfWjGRwqRBOl1DYKagCTu9
kg2wuLOwq7kXaznD0ILWJz6JvpHpZV5sF1GMCs6F4W3O7KrKYofcx8W1xek+
FsROXqXg7/C3U/xnv0OVzSw1pKHnofV0uyPrlCZEVuBAg6Fdt2JcOuYX2xOd
H14kgz/Jdq4Nwz6axh9NlGJiXASjV8yE0CESwbuWJyLejusC/SMVDoRcvfAa
jniDyf4rk3D4dpXraMjc2ZLzhcZxOJXPLGiga2K3Ml4XnK4hrb4Qkxe3FwiQ
2RkZm/OJBo6wavlyJGFOms0RhiUNzdwXIDAcBoxTCWq/F8EggmH6arH7Eri2
QxtwxCwGp5hJpIYWGsHnPsWBzHA7sjQXSd8KZsChLm3gPL5D3kTrjCc7mLNi
o5LoC37sKNmu/Lo27Jv7BVbOH8TKt0PcTWrJdpcb9Fd/LsbA7ij6bZhjT35S
s+88m54VrdRazwb9AkgHACRJNRridZio9e/dP0QFlsZzr4MVilJm7iRppZWB
AwNmfSLhIcHUpw+b0/n8EpDPKbsgeLHvn9PjUGJHwT4immD2oM+88xRtdO9f
+vMUhG6y7XVako1U3rgayrk9gzCKkNUMi3NFZS5K9cV6/IXVWzb7RozQ1EZi
Ccj9IOiKiuYKsKTr5FDdhl/pT4qwjpcJ48TN+bqXhQ7lSEPfMJ+cjQQZxdlO
QuoLvJE1JybgswVYgl0kk7Ju9te04OLmqU/CgzbR+iSJ4obkZUtcvsW09lKs
DveyzvdItQNxUQhLPtDtCjIhm/x/x8w611ERNYha2EleuC6RMwUjrsnS7lw+
1vml6OzMNhlpgjTBG0n83xm/m9fV7irbeiTMX+cTwuIZN9IBihClkRVNn6JV
O9OONzE6WNooaj2WemwejrxEvFEtvm8A7ms31gYszsuntqr7SPWS1b+L+7QD
5Sa31m9b9WXO++I/ZyCEAsSAnDGiKuUJEWYIzqVCRQvnRSNXQVUXhqhUk2KT
236dmaT7T+HHFYE650yOKn3gcVl3XuE5+TqAFTKYti+UwBH1Nl4C05FyKAFc
7eIdPV3qQot8SVV4EeU5o2KQ/Wwb6x8dRReSXsBWnHP40HV6cJpiULZA/0/e
w7O4o240AVDmc6z234vFDv0M5TIVPODdjNqSuzedfyXqhoSh0x8duNhySeDR
tk2sD1OzhVcaUFSHcxHv2zR/lEKP8u5XLqaIgXtgWC7DopJu/JX6GNLtKftp
Sgtp7uUPJtDquzwIDLc/4wfhjBYwDrbYPvMYt4InEgnsnuKV5jl+8ZjEWYZ3
6Geem3A8AqrZvwSMa71YutEFQsEGY0VMbpFUu3GOt/DGo8jhe3MNuq9IRU9Z
0bMtmuPgo+Ifg1Y+P1EB1duludoVsBm9vO2nfol6Ymjt7F8goDOVwqs9/Uwb
7xu1Onvfxah8zOD1ggIjfDFKFXUqXIUtrGga76DYIqFjTAp4t02r3MV7Mfyk
UzC0gBU9i0GblroosZPcArM9v4IpXsDtT/YCH1jxqqZh+UMfTgkS9pHjc8BY
9B1rqOHddk2Ch42MJSVP63Ivwq2kgISsPNecaaCWxOHYVimWQk9bG4OuWv5R
kzc4L74aJO7QPSQKsEEfkw7/X6cMxunA2rfmEYWvt/lLvKB5LsaLjoR7idq9
/vUE7xl98G/VUAMJFgJKHNVYoNzQYee1i2Vj4pLZzbtJuWehJKQA+UANEyhz
bdkUXRlISF43shlmw8M/j2XRclm3+KXWSJK832n5ltpoakP8OYZo5nI5a7Ml
e2jDDwHPpDrSKe/TyFABHMgdK8ee4RgfZ5DllZrFiIaQ0dxdiyPOLUAZKYQE
Z1yKJnFV/pFDkO2xKQw8jtwnt2OW4TFmAA93GLaiopxGk03w40dbytwQRVUI
hjzHQHu1AaQD/hOjld8X4174r8ge4Ifp73XJus9XkQJ870AX4x+JxKU091li
AllQP3X5qAVYOr0oMcPOKIC1oLpBmMYSKEL4Jjx3tVZamO2B9557k5oVVaka
MyTtucLKDaIWwXPoYL/mGQc23FGzX9aD/N2Z4pJAcuLf8H+HTWSx82k8xT91
Z8X2kxqMkZdPUSCcYGs72YAdGgLIKvfFBMw4v7wJm+p8CYrb2XRbAp6FRF0o
rb4NxUjuFc+mvU3YZehTVxKVKx335nVghPAQeoAJrGUdED3zO92L06ZXq4rN
fvl7NHjbDtuKQFZo8KS0n2wS/cqRiIZdsGIgnVpnjG0G/FwwyYQEgCpsJgkn
NLeIeDTitr14EHbdef3Npm+qA0Mt4VmyEIhbspXcRa1EqEOBVWVY5RwMNq4r
PYYjP1wlTjerj5+9/+ZpFAfjMtiEryRFsEld/QvRe5hjSRaQbRBogVqHBBzj
aJB8puo6UPvuCf+j01ZFtNdVpsoXxPHAnoIFdVjIOFnGDtSjNPUFNNERNKeN
olEbgKUX538QwHzlX/W7ebRDcRI4mnGsM5yvNX0//gCa4EmX8gmrO7Pbjqu0
0bUqQ8p4T02GIHZJbMU71rdF/zbPckOUqH4M5SmFNWfDYrVng/qkQ28wz29e
ZHvXMrRiVfAoiQFh02VC2iN4MJ6xJ6eR649yzQvqAZfqshRH0vBnlgpEr66W
au/c58jxeX9WmqhySpVczqE4dwSomG93CSZcIC9eZpqaGASoXNWWsW648Tpb
IznMENAytLRnoCciQIh9ogMXugLr/Ca05C7l9ghyNNaEAguJXse8kLhNU3iM
F1MWJMnQhOl1u9WQwf8781iLzlolGZ+uYRzvy4F9MxDcBzN2OjAlCRD1iTQS
oYPrMw3QzyL2JCxaacyEGCmeft3DUBlCfcPraS4zFSM8//UB0e8hzSGh+ehR
mECUat2qqgeZXBVsgOWinP0bXcKUpttgtTTacKKd8DB8HG2DlwoZYzOcDdZt
KEtpfamrc7CKRtBEJF5FVGz/ub1lmCilWo+GuzxFj5vyBGkJfONxOR+EbTSy
Iji4m/wKoyWrhKbPKcYJpa6NGbAPv29soxmLxs4FtwyUyWUvXelutqplGP/2
B0OPqoUU8UBjutiod20kMZSochzXTJaXIKJvNcAhGw4BvGvL/vPvFwIcsRhC
a5DH2o+Ohmt6XVRafoOKvYWBarDMWU9eRfxBdlV+f6b7A2+lcOXbfcSBGAxF
3i8bvzw2g4GMP52Y0ldqULRnlvZ70F2hfQj8ljkHn5wY0uHuqo0mPr1cWQFz
665k8Q4e9d3mf5myw1+jdXT8L5iDhDtYzxdQG1SyIx5gzvBBZmQT6gq8ZQsB
PTnssYvnGwoPDl70WRC4D9RrQZm7H5mWhnPsy4RQM5BhGtvnXWh9a7q2P+9z
8Tua1qioOAqJ0szhsQWyTO1p90kpFVLfUbyTHnFW7pgeLviKjUKsc9DxHbad
nqJOzlansOt8iUPTUQau4eyV0ydoPbBbYEe99nMfjOzrr+navN417IPQtpuZ
07fkwEVi0eNkZS2ouK2u1nYTKlmerMQi9VbeVLiuYXFOueC1sp7RFc3sR2Lw
JqkPeAtp4iVokEbMmZYtN8qgvxTRsyoC/RSmEU46eRzEinB1q3L3oLtcTVng
CdZteov01ew7g98hMjZVoBikl3fzh5GcDfpvcQlgkDFNAYjxrpTGJbUGki6l
tR7ZEJ7VH92uYeYr2aELTComUfab1GS5wwKprrMxo4HJ+70w8kLavaXLnym+
2wF88PNJ0eLyNQyVy+A+H+FXmGu0lgC7p/zKXcgYwIi7dq6hVOyPMf91ZlyC
lkw/nCPqne5yuRHlOsTzTreB7PTDqiOK4F7W3jRRYZ01WdQzTFhhNzrcA6MR
HMsbcVcgj9d9wLgR90u0Bd/v6Arob+I+ggaRJJHCOLx27d3cpYGpOeVEFBHQ
HSN0vY2tCfs+ItMlrzEvJFBDPiDu9euRL9oya+ch0cAF8Jsct12yhGa8zJJP
Phx3Cgm6XNndGIBP2UAA8bK+nF+ohDLy1Je/UWBZpdfQc+tZWqa1e6vX3Uai
Sqsgh5jGiToXcblIkE1FoYB4lZlUIYWxgAIMzxkzjREv8zVFXgtrk+z17xaE
JxVb9NMSsDtyMLRLqu1DY5fTvVxX83TTPH3oAm/afaYyL6lszTW+EdxF1zCo
jOLpwdeBsmBv/oT/OFV3vuT/jjc7xhZNLxQkeJ1eUiboLK2EEEI0C33bq1mc
S3cEWwSasIB2s5Z7tJvm9obIvmMevTuhR/nzVIeXZXnBz10STK+C6duwMx8r
FxQ4U9w4uJxButRetgMxa4Afu+2Ex/hEkuBtnc/F5xW6tCmtnmx9n8JnmXin
MGgpRBrqHJIfquLivXs5RVSSn+bN8blpAf5Uu9hq0pDp+zPnhgeZip6zQ98I
x00yAF010lhokPjCvkUNTtUXQ0z4dkZNc05IK50RjCIf52O1Cx14oWgGmwVG
WprltcwfzX2OBaCEaiskkxWTa//tJlWUnIwtRmo/AEshFx4BgABBbLZCWcUC
RH/S9MvYScudMNsQC7L5bxAlpTZwoTqxeBV9pwktfEUJgPF8lI9ZKNoWHpy0
ALG7JcXOVu8qTdZuR3UuGqiYseFYPMhIV9xB1++ZfYBQIBmuaMwV7bUGWOqn
gaapSgYK+43JUqb0hsxYLNQyrYNHmvv/giIsFEt3K2u62ksnjQNn8NLcT0LK
LPvYKXPQOOeMAi3tYEaYMVKk0JbizqHEkA+0eCryOvsI3gFNYhuITDyfDwHB
IMqzuQzEOBSriksOWcNtpWMaBHlj3Qvq44YU4+1oqcDbU3Zx5tyGnR4BGJOT
X8V2E4ST/rosMAFay9ZvzDe5teQnIEpOxQf+tkncVtiqdwvypC0857qub5XI
qHq+MJYP8BE84reCPA3vDQMvXnWdY+lxnLR0oDULrT//mBL2PndiLLtdKnQ6
mkbVs0HJplCNOjHrGDb7khBBIMEjTsFiA2k6GMFvcBP5ofsZZw3/LIoQSoAu
QbwNdWlbzGdXb0LGO6AyZt/injjlvMUSGiQiwAN4brKaxBosZWfRPkk2AC8Q
lPRqs6VPtj8JGM8WPhZCwrrz5DUWaSj551S8U7LmcbaGQ5y7K110Xmpd0Vpv
X9KcCxAjsssqp1iCaGhaba2yIdipBIhtpoDV61nClCsEnqqOosdD0UZoSbPO
bT4V0oS53NKSV+E6o9w+uHDpRw2yE2Zk8IgJ5xapfmLEmhz2plvNIZXnqsVn
orqMng1Qy2WqQVei1OuR+AzE4VCe2FVV9eZ+AdeBFHTuHcavRlune4qNRUTn
tXv9frMCjbfNQQ34vmWRY0V1RbrEZsgWaJLnRfsUlf40qcjTwS+4hJME9AZd
CBIY0tavjna/SxlfPbr30figX5G87EEhN9mLarvOXv4TPaeQX9Y8asN4D4Yv
t7BbzdTakzhVyx6YIekzO82hGLul7/wEST14feqSkP43iw7egWM0Xg7qGdRE
34Qlwzq2NOxf4rKgEblP3ZdKd44jRN9G+ckG4mPUp1uVJV8v5SGQ2QdBvpoS
aY/xcyma4KXUgWLGXBxGn53tRD4AIkGX/QvbcLPpYK5QrxfEoW0uOgWBjYV9
ZlE1u8KE8G7TSQxHno4q2dh/UTRxgEgqAGnLiAdcqm+oH3xpGAkec1utcG6+
Nq3Lwh7OYtPPNbmQh+2JgrfYTI4GQG1vOL7hzlWz8+VNPZnJ/6ehshznnrdx
YXBaS9vk+NqkWLhG/EQtdXGrkAtD+QnPwTowoE06ik30hEmu8CNGIrEtdIra
2PXXo57BrE8d4KcsJS15W5yAQb+n32Q5q/5RJmdfkULn3e2k+QjqzSBJvZPJ
juDAINnWNUgI2ta6ebfkS5K1jCQzyI+zMq/aR2I5TDAAGAnlCtW7UuwFpo0L
1PdlkbpkZTp9Z88KR1zVULLaI+TBnv0DJBD0E6XEc/qBV+XJOquTGtafqvSA
NaQGTHpY1BsNyAgicQGqjYP/ALn0nI4pYnDlBhMC2wFU0L5PV4Z+q1SO1teF
QzuHqBa83z/bAJlUiqtg5r1ZGZw9tSCp6DDFztzhv5I1eqxo3ytMHObUk6Mg
tuZHVjbrWGpo1D9IJJyEywnKPARBMixs3zZOFLRfj+qmWVvPJ3hOYLEOOs86
4Td/fJ/UEh7pazXAEpf1f0OUDSri6KFdPBGcJUDN9sSR/fa5VACy5entizEf
sxGdkl7kYaJl0es1Ji4Q/+7juc6Mb3J9XQMIUbyBH1nYb2hkwaHPeSKn5qJS
tfYrY0XCJEATk4ReSrOtLUv4oxpHv71Tl/J/C5Vz3H6eUOVuc72Uni1hVjpN
/CcvGAjgsb4H5cPK7/8sFI7EBZieOABcCMa+QXAuwTJyw7F6BlGOoN+cyMW8
QUTAWJnzDJzk4byVxyEtiQj/EsSGm2+QP0A1u/bOeMJe7WqmiGAKaHTtblA3
A0kWovTzmkvMggYmf7IsPmOAYjC2r4D57qV0tGDS5wTAlA/URU9iddHneceD
NHCYQ6IhetHo4flpoeke/CbDiy5DklSJjKA9o5dxwR4yoJg7s2Cmo6oM1Zyq
LuXzuiLbnanFX/riqFZH9A1FvVg6etMoagian9Dx72+sXBabSTgT1AX2SutC
blWD8OWG0+fpfZ8bUsVS2T7A8aIid3MeLh8HeXxh2SY/NNiT6wkUYzUoPYQb
I+XQmktZy0l86yriGEC593ZetlQIndZGoLxaRqc2A5sQqC/1QsY2Mx+7vmfB
EKjvSgL9cpS1LA1OzR3ROd+DPd3N0C/+Tc+oySCtRej93gL2ooz2IdAhBHBA
LIiV9JRKiTwWt4d+Ns0dR9NS0P9vDV+y5MeC2kvEsjvShX8oAy2KxYRJ3kAC
79did8fcxskQS4jl80eW78FGD2i0IHqfdIMwYgzwvq4uVoeS0grszWvzmtmy
WIWQ0mBlv0JTL5AaqmAXDrWwFhSYgY+ii6V3bY5ZFmSOlTxraurlX++Itxca
Vw5+HyBmiipOLZQVPPeBoxDLHDt0+qip9bz2XpzZ2w6dA7MefkQGriH9jMnJ
p7qjOVSz8UVfvmb3z44CV2/EpjC6WQwDUx1lSzOOKbNhdU1a/uNRWjcaREwQ
ooiPwBTNnt8Ul7eArBLcp1a9Q9gCHaLihC+3cMJ0+nHFN8zLwtKSgbyXgG6Q
Cu2r6v68RRJZRDzsXf31pKMxy/8yawBjuGI8tjpKUe0CGDZiwqUOkarvV9Fb
0CD3DyboGbi830SN2tjhtXELHwObU5108Ois2Zn7dxoDvOqnrDu5uZL4Rttv
IXarQjTTEYReOJdYFewiV67m53Izm4EW9Zqb92ekqTRLgsKM3dQ+KrqPY0AD
d8r2geaD4JCDtoZz95nrq4FQHD+bnlCniojrjUJ00wpG9NOM/jTrA0A0bQUX
Jf7x5JWS8lTMJ8Jt2zf3+WguBbV9sy85/Bk1DuPoGjcHpzvvf7XehMFDPAMq
jz3kkJnya+0ipsVxqDYHCfGFrdea3RRMeFnSYrS/P/WMfvsunM0gHZJuJGJ5
4lY/8AapV5/e8nHL0VgUPrh7FL+Qkw3TtQ2JX0cIx4geS5Jv56QJkyHLV5rw
kaCCvJYUYt/iCC58kez7N8sGokiB4SEAU1ETQnNQrUya3ahfilYNcqlQurEK
+/lvwe757pH96cvVV5zdFw3HyEJ0u0g3t0PbfHDJ30FtfGhDE3501OeTxvdZ
gZY2cYVwVt54H7eN0OOB/Bgs77FF4OzcYWH6sWim0YRUba51d8jJXjqEX0TR
2GoHj19ZmV4dylf8FvjRX6a+CFEI29BwWA5ZTijiRugEtHo8CBccVn3cYVlb
wvnM8BIwDnUBAjxKKvOGdg/8LcPirFgf1GlXayTC0HY6XFRVfIhkG3v/f6u+
23/AU7MeyoFOmyDlStPxZEmnyGdc0Yhk/f1H4NWqIAPlWTyDt7aPmjuxhnTT
xapwFp9kLFljQWQCB+NaF1dqF75mXw64pmXjmy2cUE0ySaesTH67O+z60Sqf
Oh1cn99BSZQnrriGRn0wm5Cb+yek6qngyf4S8TQkwj5scIdL1J9PBJuBL/F0
y6GGzS1TxTpa+oIQm2df6fmaqQfbzXl9wkwnu/GqG2DrWpgQK+RMip0p4UcO
AsibHtEnh9UsTUF9HHDxvqx2CAFXajh+T+nj+HJKsTyJajZpTtlMzja4GcKN
Q+/ybg2cUCjeTY1HPuOXLtSRyPeNw0vlHtlCmBhZ82dzDwOjTz8om//QNRSq
4X8vN+YNMzxZq22iGMPCIvD9pMx69SqHK342UeXvAITIQQyGCliYm3tG9Z0H
LfKyijRi4Ery1K9dxzkX8yE8UtWtJgBhvaK09tVSrsXZdj58ri2uSIoejCir
KwtjdmLxQ10uED1Gjm4fY6Bcz/RZdTGAg1jsI4TPyqETbfiNx/MRgnMB/+YD
tNrqqzYNbHnDixTyvGV+VLEMDeJxLRaPSBhnWjF7jAxZZQXqTB0DddoS02qI
jsEIGsLNNzD5yZkGHQapE+GOTrt1bgluC9gC9KG4IIkYVvOc7OapbTH1LFWf
lI8CIP5iCBIbNAomISwCfFt8f+V62OU5B/jzYvj3FlLiHoBaHijjb17Hfvzh
7Kvv3Zu85jX11Adk6CHDRKbNxi3e4g0ajLUAP/8+LOYN45bwOfyM97wtWFRX
I+gaTx8DFPBWLIsUjW3gVvUbZ5Sdmh1/8S6XkOsgrUusjzD53nHHpuqLh5g9
q3IUXka7aUWNWuxW2LNLd/cM6DryysPfRiTjLdAo6zn6PL+Qx63xpcUbE3k0
Lsj+5t99HikBTVbTryY8nE7dRenmW+UhwX2vXUKr46gaZfMDd6zir7eSOsIz
3/LL/pDzvuT+bjCArymqlB1hLC7vOsjc2cstbS0HSi50vOfeAOfKNC5Pp0h0
TFIaZBZqaXixgyjURSezWpaPz68MzByJjGgGa00+yUVLcNt8GkW749K1UeSO
Q7QdnqQZfPML56Nwm8nJOOqdEYu3upuHQdJ0Ztn0F3DeIcMP9asUcMmec9/f
avosTjimOKU0uddtC18xL1y/OcgsmLy+q0inLKUhYanXlt9XP7rp8LglpkNC
1cnI1ksJtv0CkSTV9Cjz9BIUlek3CNzUSye2kotxSGMWbhMBYFP9q6hOV9MW
JkgDZPjzbXbvRWapPRPIrlW6KOGkbc3ul1D63vIvEOe1zC/JwSZtVusnEBAm
sC55S/9TPDiI8nypF1hKNmE22NS97J4cHzjnPOYRrzeTbsrS5Y94dw5mHtr7
zuTnaxAP+GY9X4t3FY72toNttfuzXf8LmnByBhG46G4RezEEUos48Bu/TJ1h
c6zdZ4nopV10RH52ROCfNGMZlzS2ebJwtOPf4Nqar2U/DFACJTzTGboCq0as
KU12/FWM9fJea7kIr6GAPlFh+uyFrGWVDDXd63wCgd1BObTtKri3xPzdXQvv
yp5fF+67spm9o55x+vudtAvcw3m8qJcseY2pqyhJ9mKfYYQw1K7EJ8meGUaM
ojmUsWeoZPv9uSQqg5o7EAtL032BMFZXJuEsHm++/0uwe/pGnYClYv63GTdu
CLT4hso6hpKBwZNotbwFWpSWc1IbMyjhBUwf2zBbSUufw89TOAl51d8fj3q7
pNnIftAPZbMgN4z1rNnjD/Rsjg7+GRQHNLGXrVCJEADmMXvjpQae6plswQQ8
ZlnX7bN8KVUez2kjvey6d99JniBy1sxSimau+HF803vOo+/IYYt/DpSfopDK
QtktYTHJ+jUF7vusPU1KKvsfZAmCd0vHnewgFd6zanSwF4MJDqIdX5bt668Z
l4iZMy4pyT2pwAb3zsdk2qiDphfuGefUE+/KnzJVhZKEIjXYkpv+MSgZ8dpi
8DRQfyFPDAloeZ7yJ1LJj/5dIYeD/qpA0RPKWgmmANmiFg0hK6MYucbVaygg
VwHUJiWNmOmCUZ4Uv4256gp4E+OGljoFMFoyi9U8jgHhsqYIdqfQg3i5hzHr
jNQ1ulxlCTbXV6CdkOUXJpc6JpB9m8jWn8HCHmC/ClnZssgrt8xF66s066Qd
ziK4rCSnLpSTADopGPK3iIXe3PbmVUbWRnhTw64I0/Ew7EGauMJ4Hg07cCNl
IyS/O7H40/If5UWdqGhYhLutqpZLf7OamPLGEi47QIupP5UreW1vZU6Yts/u
DIZm9cQIHgGFkYhdyFtB5BggSo3UD1rPk5VEfRqCyFyMIPrXBnEraqEvejts
M7nuIgZHEmWD3NFJoxUzqRC5cwEKrKV8ZrBjR2CpkhloBur+/UrZrOy4b4dy
Rettffyqs7KTGRJor/2fAqSzzx3HnT02RLxbbquRSB522Z/hey4bN1zJk1BG
8D5NO22oCU//I/L/EK8LKuw4OExVGAXCRP9FPMMbuEi/rOxaXNLt3sK0JngJ
gbWa2nxP/x0y8l1rdK76kXvJ5k0iupStUtdvmvkPftPluCBfWTd0+aagiZxM
3br5VXbccxQpr/yPdZVGNAPREXisyX6kl6AmwZtRvz1ycjyMvitrvn2vCiKb
/tK+XTKkRRN5aaS/SzkFt1gdr2AmL/kEXhMJdsVO6nJCSQ6Zgx/sRZx2IZQB
AQL7knAf/cCLXrYhD4akOi6WH11PnZQfT9sqhjat7n8Bs7/aMkufQM77dJqT
8Z5qOAlmlBUy9m+tWb3WPLePhbZBACoyOC9y25l2p6KaTAOm768MOpJ23RVW
8r+iDGpkT19yw/TgENmxgAy9jNRVNtYb370DmSK6igs9sxRRNmcRs1fb/xTP
hlcvKYXL4373pVm8vpqkHoQR+Gr23HVssC8NtOYa1NNcBZqXE8bSSStWp24r
yeTt/YKYETRuL5b88wAvoHdR67dXhnEr9QbM7VoWkmqsiDyBCL8sVBNKZp4s
lR6Jt8Y0T5M6nUudrrG9D+0NiqMe1PCJp7eUC2l1wV4Ig+vG8zYq39+Zc4YV
PaO/h3IJwrbJNCWHMYoffUjhBKQ0yDfxvneFfROjtI+U2LMaccFoIEU4ruQ1
FgeKKATEHkjzV1NGMJHHi6aLrThbb5KYRi2ey4RbNn16p33EXDY66g1isqWq
nSj669fVOWlwtII9VPzw5ZufJ2Plj7tVQ9Bp1orWDOH1Ll7Uyx4hCb1aXQD4
eb+R7ymYw1k0YGe3NRozzFrwgboGPrRaWqoo8IZQ9Joyt3ngnP0vyqEJid2l
wVCa2DEyeYtkQB7XzLXoAlOQA+axIeEVY60b+MQ8T+GpTsJxMg8vLVtD0Zl6
7QCyThgISn4/D/E4Qus5JqHaYDoD6dA5OncgETb5Oo532GDP40/OyEJ7Dn83
sNd9sGdW+DBCULaVVyjUg5YQWKjrJXM0zWwPsI5CYD9Se/cEnjouOqn7V+/3
aaRiQNHrtDu1djb3Ha+vPZEfYD/X6aPgEB+Gx70KW9MT3XVdbpRcTy+xg+El
IBPHyiIuX/sFfV/vUpcsHlAN4AKXTqSTkzhhLY3RnXZ4Ua06yvYQWAvbvZyN
w0hJRl/NPC7hHWYq7nIPYkoDf5P9U4OWGezO3WC4XCQ+er/uB67CMrR9p5oj
uu/rWg4aK0En/ONEqVS5CAJ92tX08UGODMK/4No0vLonsyWobo1HH2BFCY8T
2qiBW0rhrMKJk2z4lrdAunuUdtF3vNO63ctERLEsrhqB8dInJCCmNkH0Sgar
drH+0vygU+2vUgcvQCg6gsfC+77yRzvZ2YO7lDwdlb1VvcBgqwYcztwb5FG/
mVihycJUmXox7xDqN0Y0u4ls34OatmRtoUVKs+vzPPtYEbtFyrRRTRJE3hYX
1oregH6aA8vbvI5JS1t4zaSo1j1e2pFkV+nD9U1Pcz6l9yDUZZwnVCiRvoPX
VpBcLQM0N2qDvZvmCkFU5MS71kXqTsetFHYPkzQUaSr1UsPbxn/H7EukIGHQ
OyYmzw9+YD2w4LYWKNBv1O9zFdXzwjVLFgJQni2+i88PMX0PzIB1CjNhLZFv
UPcMeY5DT3ydcQ1HgqdsVtVoBMr++mtsU2ob99rmfHVemMOuaqB9PqKd3V4V
icyWAMOwii+W6TS1tpacLOWCuwqwVQsw9a21XRUxZZXKYoLAQgLL5rUQF9a5
wTR0zCCcdjeIzqcI208Xk6c+gmK8ri1kH6b1nyFVS8wNbddr+q6wj/QCxwMs
HtqmaHF3UQUM/r5fPleENK0lTHSAdtlUmDcN4o99KxsCjUHpDyHMt7Bd377l
Xji92vKTs9o+/lOvZ1TcvADKyA5+Rvrpb1ea1yUqK6uF5V3bxQa2P4It0qYW
N6y/3vzwI2U9/08KgHC74i/03MW+9AJHmURnj/Ig7KJ6sXvHFeqiwBFSP5mk
HdXaH2H9wQHqEgbEO4Kd1YAYuRj0IFG2xzvTnb++vbsdFOs340c6oSOEOBrz
ZPWgLZAfm5EqJaJ6EBj3zdo+p8qwXGVEgFMY1ew9WT3nZ/1roevBBD88YsUO
0XW3iz79Qsb/pdojmXegPur/pn5oiTAGCIWBk+hexkIVYcwh/0rOP2ZA5CuL
TZD8D1ncbirweAS5PbbKI/KhEOqV9PxlOx9DxlrNgFYja4yUpLqg3deouuyk
/qxZ+XN3fK6Zljzed9F3LyXq4FktxLrRDx3fDF7ubOKn8HPCpCEdOpxgN59n
PTrTCjqDzdP7J9iHMA6noKSzZhq3PtD9yHBEOPUbkdt21kaVS6Y7zxbzbonJ
84X7a2LEy7vRuA83o2yRMLEfT0HyUnQryxnJxuT5Dma17FdhqbvPRIGilHRR
WVgod3TCV20nNfW8ddCZgmO6P5SSH/qcXGBesB9w6F4vvmrACyWSqtwpqvHK
w9Li8qD12EjX+pObumUnvbiME0pwJQ7ynbCwawmk784q6R5YCZT2NHr1G1Z1
B+MyQWQD3BHwPt9DWedlVI8laiiXJy1nSJqwZNDohtT/UIBGIEIT4pX61CFT
6pRrdt+yIS5uQeim4NxwLG+9l2504XV1Mwywz1Si+tiXQcZ4hjtm1AYvFFec
OP5BZopYCHCH0IxwMVHA4j36QqfcTLWXT2J0G+8KOUi6BjeLVW2LMj44j8hx
la35miY61ukiID8djVY9gtclnKRgq5C29AzMUAZJguQuvXNGC05YSlw/At4w
WbbHaa60DJbcPqbRTm4dA4LBCZv9mkBfZGXqYfPcNHuL+R0kdvxywmizyiun
en4xTYDryGMnT0pCWMjvOWxaDhvzpT23JhTu1Afjjx145KDo0UZ5VuTg253A
XT4CqYNed2cOUJb0/DLnMy3JAIGIen1Avo1h+sKfIIsl064I+b7cqYe7GhnE
kEnBWgeE3wGPtM01qpxRXXzEa4TtFZHv5MwqExiTblP2a+7ivMdi8kF05EQg
o3cfokzHZob30EO8+QnPtfkOws6WoDZAmDRzXdfpnjh1rVrZ0B3QdvWguatI
Q8Wp/ZD9VHgCMLf73h0Fgh4ssJPcekn2XDVs1ofng+s/ksprzv3BX+twWH2G
/+Vd5E9zruNfR9ahVRjzul+BtIWC9CcagDsGPTWDAP6/tNJPii3QYA6IxmDK
Y8Hog7xA4jgkvcM0rV0yy6AXqfSUEc1S8oF7YVIVn7oVaICdSaXL0ExQZgby
QhCrVFYF7rbhZQi4qEmYg9GpTZAlens8BEeNahT9bYoFvr7nQOpXb16oWKud
2sbZT+KLT2IwF5QGWXqNY6WJfFDTg/B6gjiLqpKsDPg987oHOWbetUZ20x13
WzXaQDfm5bD9vSSo7D/F20ZmX9yY6N6B/AdhoszyJvGkplQCwmtGEz2xodFR
9dyexkSBX8DbjteEqR2wnOI2rAeRlMWguprWW0jtbulvdysg5zr+pBA1/CSJ
JmyLfgCV9JdiSJgJyFksge3f4LuMIyyT+gbk63OjlNQay386hPpvEivAwW0U
2Z3lF+kGXGYQ8tRyNhroO8xydXXi4Qn+7LMIKfN23BKegsXD/FLyFx0Q7B5t
diW/nRdGBthZ/faTyIJ9c8E6s5F+4h5AW+rthHqi6UUr4qZH+3MzHCyTsT1l
2lWZ19QrNj8gjC4l9zz4LNJKe57yFb4P2Sj2Tl9fCHUC91pJkKQVfDGmfbom
rlSzSLejiv9zdF7cSGrwpLGwWvO81tWU70FRJon4WW4lulwVTSBXh6rDrP3G
fn7EibPrYi4xLQXfpMq06v6tmrfE2fWQ171L9K/k2/bcAc2jxUAhqSsRAoko
T3n85BoPgs/tjtys/39t49rPyjVoGqz29O5JuXBPcL3iKh8HQ6eIJwZ5AQKl
VWxh2Ykwa4UnxF9m7qYOix5Yh3GBki1JhImLgL37W8+iwB7r+TfjwQK2msBo
6rfYnuC4pNe9XwlaDFQjwWhQnT5+Baf09Vk62p2eDBarRC6FyZOVa1dX8y7J
Y3Yzx0AHqR0cbwiOSf2gWNoJ5Hi5J/icL+rZhzpSStNYbnNhKaK0lz50QIh0
WeY6wyt/fTCVYW64Y9V7u1SQI+vAUztylpaA987ich+xQlj9A73hTJmh9e9r
Figo0Zx8zf1TNArt0XrfmNYsFQIL4Yrmb6/PpWMLKevJ/Xpkj7jzQiO0wC5b
04NZI55mT025JU2fU6aLV6PLb13PWRi5anYxr1go5oHj57TGXqcyQM4coxlE
71JLiq9n9lmOk/IX7dJJNhfkkMi7qHDz/RYxUd2AOFGl2oR7i6e+ESfxNZVA
lgl4PHbporyLT+ezCKyICYRPOe9NP4L0NBqz+CSaXzVJpm40xoDblKOauH0j
sr++9lzsStUFZV7eYRVlEFPEBIHP2x64M1W5JWSq5s7aoGeemsoXPD+a5bs9
SWrKq0EgM5IrxlI4ev1ChMRaxpuh/SS0cZMkUl0ypl/CvjqqY0l1fA22igkn
ceienIGfxWGcYEnXNZStnoDFmxI5r5ajuGTA9YnmGMrOC+l13siM3C9+goz6
WKZx5jUgj5gpgX9vAoUHJmJOFlXV/Ebwrbcz3Qo1bp9I17hS5NL8cxmfeASo
z5yQPVk6ePB7vyuctG/k5rl4CB+H005A6hzcvmyxP6k99hXky2EEJXTK9UkH
hQjxe7ZlcW4L3frXE0RcT8sIrfq1ZGRdkV0yB8KP435fZksQAzWn06br6AfZ
Y55uihp0q2FUhGWo5FZo3UatoxtogZZ7SatZlyuXnQ4UHKzWjD9NdGQTMao8
ie9U6JoZv1ibwHHJqu+36hhQehvQPzDYYhej6RoDP3VM/i4ooEBghu/Pr2S+
SXaSADjvIH/s1hmiNDyBV4dm3XAtAIuhB0yRHwou1oFK5xzwZ5EcWvvjSvvV
K8+FCiyf+SjbhC2fej6Mc06EhTzxtOvC9oglzECMxmo5vigybS7O5Z6E5DpO
ArumFVZWdW+AJVfuvWvGcq23FgKtuhm0XH0PD5lDYSXvtOcRX/PtwxCQniu8
OzFnpqz7ZBBV2yofz834S3cQbImKjQHC6ZBgmqdkCHZ+dNJMYtf1EyW0XIdR
SOLHkgHTOZDheGRUlDihjso17ZCxd9ifXkArjBqkfl36ekFISqWN9oWUcqmK
ne4gj9ntAGmrZogo4/6+28ITZqgUz5USQPszqVwlwCbDNCKTPKbrS2zha2BW
EMBrSVvClpMt1U0o1VXPlKmf+9exFUzjH1fH9t29c5YaPEyzMnS8aPT8Lqrr
Hu/Kc7AqNxvf8By9WhMsC1JA3hhcNsI8WYdknkJHUzh5HUDe2XwN9Pr7Kump
i+chuT7qsqJVsHd04D6OX5uLWZNnUb2OQaPThHhWY8q3U9zXNdW/BkxByHTd
P4zy2MABbnRx0bOEut1Z6tcpLqqwhNGBlkMWAUokkL3sJAkFAB834PIFmXJp
+Tg7IMM2gRA7NHmwEDMUVsIXhpQFz8zYyXXWMrmeK2IWuVz4UXc6NBmaNw0q
x8XM6ZhDbkp2URFBxR9UNey49OreKMwyhWGbYfD+6YZjlMwVY/LvBbxsyfk3
Cxqfms4vWaRUUqY4QAuxp0PuO+Bg7ytHbaBQdcpyplWEsdGNugaw3madGnz3
PdmA45408Ms40wPDwRJcEQiCbhUmkUX5Duuw4E0dwZp3ZrDJv75Q4pYZ3Kxu
+n4ZBsFgqjQO8Y7O3yvRBJ2jEmpc69erhGNL7RoLr1vahOtsvBQ8iKSaqgoC
fvZBFKLxoGU0dncH8gWD0dmu9w4uJRu/GLwPWotxgJFlw/3zlWx917ja/WlG
X3eN3Z8tSSAoS8SDuW4Ucv14lonhCjiKcPN97paH+BYasYmaINvhUKWZHdjy
D8agW4gPkryAjIVgl9YOWrpZkJv5se1fTi3LTivYoY7gfEHlEbdl5BPOFwc/
LfIDZlpc0sC6BrPmdgrZsIJw/0tcqrv432poQPhktxwTGMmYr63pCnk54zI/
r9gqvKNXMADFB2aayznj+s8cmg2glMBgAHkGD7IYBKVL6vWSKzOt8PHxUw1h
+TgofYEGHUAOPlN3vEJ3rOLM9GcsOAs1A5eKQA7nnIk4JehU+W+wqEZRlx+t
NpomSjGNcbnaySs/Ayo5mxujpM+TLciFJZni8r3B9CYjtqEGJeKxHVkIMICj
vCUWbskDzjNuQO10+Imru7hub763LHViSYR8JquF7LLZmniG7ZPBfloxGVXB
XVa21ZanXxcVd8P1GFuqBspWxKsluIYLJKd4+40hVjDHiFAu52PhRFVT9uAJ
oAST2KoKekbkSLRjxHbm/nc/sJkOn6ONid2HlgWu0uNM7+uCPtyuF+8Tw8C/
FOS8IewNKDCexSfIhjE+g6mvYWktiz9zALf85wSA/ab2vkL1IftFzUZpGPvi
Q73b8AoiEJV8IF1g6Hk/llfeVxy7FJIsoljaVX155pYbDXa2c7f5hrIk2VPe
OMASP+GYJZUo3YLgJtV3Eu4bvz2EDJe1AYw9QekKn9+65+xFeOwkpRMC1vGd
TfxCYsqJKP1w4YM521pb95zNgelwdZ/PNUU7GBkvZdWnIkOGkY2tcUYKZQZ3
EhSzc6J4M04obO/1oV0jiQKzMHd7k8ESXuy7f9R+EFhphBJEGpyFLFMaxcJk
nEPGH7DIoNWpkkYdB9I+ZpZSSiTA076TPAINZmhtR6JcO8ei9/NjxNDQmVRa
7Ox8OdfHgoLEoZm2CoNKpNjn7drBkVHUT/UxHim7tABATZ8WpZRctyvWeRCg
fxCZIO+73Bme9MjuielOexHk7BQWV+Z481i9uDmSvXTLN1L598rIy73Ybhi9
GwPXH5S/8UXYGwRly1Uy7k11SRxGqnKttXNnPngkarKtI7ZkBpHdsQZnZPjD
TdWun8sYyh9NM2OnEwusS5QmPPBzjpnuYNNtzSwIW6G0snDMHmjb1Z69heZf
L7h7PaGKOImkiC3IbxP5PWBLX16Fula70NeccohhPglqUvptWF0QWG0mq3qu
zcPtuUjGUdOHJlw4Ni+JPgS70MU/ELEd9u80HuiaP3Bfqv4X0WPZb6+zt1He
9IDH37lunQ/Ozw7RPi7FnDJoqUsiTe7j9ekjFVdQiVcKzdky3MnuA0jHbhgn
bYV5OUWxGKRtP6xhLkRs4oun1EgWRK89TdJ0ka4U7/hmmc+cSOCVJyLpWY9N
N/FrqFBNCf3IRT84OTqB2Kai/u2C/cF0Zl98cOVy8U9VUGQQ+s+1IYp3GscL
zr4otna4HMkB8Z8jYKmuWmf59YmuO1sPVoVIraqz2+LuoqdVyNim9xBnDMb7
WzByPKki8SW3e50AFIHLlGskMD5SAE6bM06R6pLr3jzXX9sIXmzO2Ucsxzd/
WLF2j4nf7wKBsZnnzAhNH0PDNHbeY4z1c2d9dNQyL4uyKrXtF3OkGhf3hYeh
oTuP8i9TfdnKFQ3nABFXGSZ3K/Q2emcdrD17OqrhXHauD6FUBJ6vksQp9vjk
Qalumv9DGTP6xbLHdbuWlmaRa9EldKtftwjLT64yFwijlk2+h8PT+SLDEk68
xpifBqxpxMYuAi/a59ArWHZNZBloX7buaQna1lTaD095AO/IYLbNk1QO8N7f
2kt8qd1AlPcjvbpvr28MsoG2MNDkUzn5M9zmR5seh3s+OYlRQ7+5QL2DBwGa
3l2erjZLHxXPddQjmI8HGQTYm0htV7JA4dVl4qfLR/VsbywlwVZ4iwyokJwN
jCMQVAG8g3OoySUmz0RRvwcJHPnnjdRTK4N7vHImHsX1qOYztBB16P89dRPi
IbKsyVfx5l6Axl7MlXCu3xWV9cTllHaiuu6amfjFznHTe0x2CYVLGGv2Ucof
JqCZF3ffcJEjeNKFKzySHZI2n68R6f37v2HH3GUZ/olHCTJDkxp4afi1Zo5/
8Nhk3Vqc7RYnLmK2Sxded0LWvDjv7bv2cr0FXqguzf9mvJSLC5iandbPM5VZ
3GKQdE3kmWfNxuTYqND80q38pJ/mugsaFxgOKQ1rS5FU/4Xrqcx6SMuqLuy0
vYWYsOtPhgLAd1eJ4pJUUCQbHA0defvhnFFAW6eBZnerCWX4s7R+ETNWwnnH
+5fK/M/1howUnLS3kX9jnFi1eiiYlN6Qah5ARTqVnW9wxGtBBhrro/XtW4zf
ZtFpsnNTQGoYuiMD24oxPBCx4RPVw+W99j42IV8IpfVOAteQBvtcX7CYO95Y
L1TCORBr6309pB6Dsh8ukQB+1qOoKucqswYe+nQ9nbHd1qwFDFk2NtY95/Nb
bKuM+pl48ezUwECUdfYiQ/LA3mmujmO31liw00EEMJYtwiRX6ViuEr2dFSk4
EfOddRmj3iOJdkS0Ay+E4ddUfM+5n3tV7RYFdZNnbjlh01Eftf9ipg49iQat
iL5aFC+S5S8y03Gb67qyrK1Uo72UmqL/OehiG1hK5c6Z3RmhHItNiZc+wM5n
FGKGJgCb9YWHaSgUDjlQ/+tgARoCmh9a5+gv+Z8oCwRyW18sV+h+fYrCAFI3
S1IE1yr4HWiSvu2KKK3HqUyR2m9zoUOs8o8eNIRq7sqT7FEh+XhYA6f3zWtV
4KC8xRb1gNhMe6uGH8YmwOUUEw1eFz02aI7UgEdUXfEBbwFdKc2WSMdC5xo4
omblpVkuKNCKFFb0fMrD7nWxdpfS+Dwa8OuatGJ+e7vky7iiYgSUrMVQRnhr
reIwSwLyoys/A+shR7e5N/d5wo26EYOPp3owag+0jnvxYyvtWYvq1K/gURrM
ExsAcH1gTtnNi+sGMM+AEvo3W7bW/hQ8JMEAOoW9d0vNbfPSF72RA0wjw/Dp
NwioFZtLlEzSKBoQmHwyC/tS3SVveFogkzJ1Ap1C2lCP0WBEt6pHFDCwAkdb
hBe9IDxSDiuIQBW6lp5DGAIKIJB7FFBJlD1CsOC4+MztY4jOEYTeHWV1jRry
HtGLPV/ZqIsQ1MY7pd0CnO+Q+ImcexWvuVY6MdVI96xTIhqk6r8GT8Dm4bJx
+7BpoJL1wgUQddEJhp0HvZXKA7W2HbHX7CmavSO59tDYLB953eU0jEynffaw
KTvI08WlcDVGTZFdt+9cApY4N62p4xQzQH994JFjBEZ5Te/uBn9KaBTqXrgk
8mgWPwCQ9L2gP2WeWcj0hNur+j0pLFo6l2iTKpE37AyNp1Vc8k1ahMId2H3O
WqaAPjZitgCfCfCHivHfyevMMqb6HPRrn6fZTz8Tndyl5zcq7BuCCHDoo7s0
sf0fg1a+JpZdu958lhG1BXtETo1CQIkwjjPjxh0PzLO2QIRoRsdBVmMc2t6v
On/I2NPRasRDUZOf8dc1ynplvTrca2prGt5Du4TTanEzLUW1zvWrFYmp601Y
sHWzrE1olmCbymXPzypBd3ebZln7az00ADWjXHY560IM1ZkmHwiFONgDoPzF
ps2LpSkPTnArTjAKYAKJfMh98uN8X03Yk45WyDwHVEHdotSinjgOGcW6FMg0
HOid7jwOii8eHFHu7g6TNReVlV3Xk+loNPHXRNvuAIxBmLx3SXAeXScZHkLZ
psfSzBHhq3viNrLK12htYaLRRo608PaktKREtWLRXH425DtVRbyKSgng8Dvc
0yTNYOpTVYHQ/NcKe24R0vYTijtxgRK2OHhPHerSrTnO/YOIUWEgjAaERLoH
QBa+vmBp0yYZOZ/AesZOmqEzfbBSoabA4/58i8JSLhGSEuPuX27PXW8s8I+B
7GuJs1ezqYV2cV3p4XcOnGdI56lo6mRpthpVGeiL1zxzQRKpjVsV2Ntv4UfO
Ew+YmQk5V8+Lu+tjDFCAU0GpykDLyNczq/dHtUplo5pqy7jUx5ygrGy/kWaN
fBSK5TbMx21MofUfHzMkxCw1umnlNRwytkZ2H6itbXM9AYbbOMFEDU2O5KNR
WPBcyz3E/3AUbh2/11Z8RiCVHttqbSWENq/IDkWvoa8RMgJi72wEW82mSfe/
wBqyBi9icPUfqxccTPf5Y+I8cF6hT8G6lYBJGhcf5Xbb5Fh1X0sYP4jsXHL1
zK+ofYQ2slJKRj4YtNtT/pWqrVzYbowkMdpdAIGSWx9vn7Zofd/ecjyb5kk6
NmLio0BdtjzJVBo9S24QHp8Drb73ME0F6QTAQvykDMkAHN1hq1/p93cVV4n/
PORRaQqBOz62ILPKmAr0lMQaOV2HB5Wt8horwEUWPcHGJB0cBQaGyhxYXtsJ
gYklRD/U/sprSi8SaAeRi0by0OMvmFhnhXmqjoSaEJAHEiDeje3xagHGPNvo
dU20oxJZfLLW/zBCBi4eA37ZU3r/A8ySxlgFkcR9O1lTodACGIrHRMuWBtpn
PK7d6rKHA1H6JHKRHnXKpue/EhFyvUPEuOichjq3gFAbhXitbu/9RQIwbXTB
rpzOynzxORzs3S9rpKzmX6fb1zv+KnxEu9MfBKCwR8GtzA1Q1wiB6KnYhJ/v
jzI9wFk8/oY80Zt2c6K2ZseZmGfXmIkWeYWtj9/2IYAIjIsLtVdoR2kfg8D6
6+ZGubj2P3zVVyJL50qDuORFKd573t22LEI8hBKcj5tWqdiOaKsLgb2VmvOH
Et2XTUyzfmzL6wK8iE92NjHblsBMyBz/B7MTpTch7bnuAF4lx/NN+RRThBki
qig2qFoBE22mBzaMJ6LeL8mHKSKOam+ks0D6ii+2NkvDEbOyIVYSKL6f+iu4
6BOk4WYjknw2pQBpPfV+3JML+vDEemLEqwpIjuDGcp23yLIveECzErk8RN2n
TetF+MZ2AogIYymnV3RruHsUTUYL4pXEKSoFo5STsguno6CKMuDFxpugfvrJ
9s2UQYMwxxr4bOQeMU2zs90B0sUXtxJ4+l9iQ8pgTaO/++3SFtIk4INizP4w
3F83N7qcE9ucbt7JILYntXRW+6uzcTXCGDd5HdXHxPhVZ0cll+HpD3S3LN6u
i2ueeERCzBjpjlgT14Z9DqF+sxO/RdIkjycrMZh8WVdMr84j3IlxtOOeXkHE
qectcyalAPI+I50iqeQD9inc9e3Wu4Y8KJwgmAm37Ijb+fc4ORwqZXvMisu2
B1lEe/FzqqlMTVaFBJxWKlc87lQlrcZ2ZyE+KoLMj6NMvcawYBJPleYxxru+
8daQyDyn063HGK80nPttnlW9uTEFc/xetq5ZlqjHMJhJOjQj6hs5A/Qv5PxL
j77GSOyR+fksPGliyahKDyrLJJHtI86jSmf5kf+ScIvb/7SptNYksqVI67dJ
m/ePrqjXjzwfRUNddPCTwP7x/UqXRIYnSzguUXzUUHS9Izpgv5H7ub22yx2d
zZMFdIDf3P4+hMcXArEujnXYG9a4NDvCqkQ51TELOchY6tX7uxYnMXEn4+1J
dhdpBITRdiFHTRUeUb0/YXZJBoPzet+xe+aW0mPpqTAVSabwOEaI1m1XulVH
VCS0kbs3TL6FSAj1sHyNPzQKRWLlKt6uoUvmthrPvmtb4wt3vPHoG7FAtJXp
q5UgVSKhaOFYrurhbkMviBYWS4EAtEpcDcGZxp07/lejwn5x/NDsBXi1l1Zy
Bzc/MqG7ZgfRUy/Q5+wFHTZ6vFNn0YTi/ynQZKCz48SckiNpLFUhwvd//0pr
GvaW6N/fKh5uxDcpdOtYOU46pAxEg5uhXVByx2uIP43a7HlT6KmFuTCzX+vK
cIW8Z1bwEfjBEiCjRv/80HJaNCGPiphwqjjXPhVuIjZY4JFE3BtvGjOCssfu
QGZJHbryMlxDGorD146CpO0KGy83LpcCtqwXzRCpxdaJpiE4jCi27gfX3L+P
rWLa5dv38PzG4DO+3+h/LhLSzxZiPwv46YdLouF9QsxOEvHVIyJY2MNExnne
GACEJC5mkMVOBWOR5v9cism4zpIWV/wem/uq5Ql0RoIUhFBS+NRL1Gi12WHJ
8vCpmI1f0F2MXa5u8P0ntSp9WfU83aUUKbhLqBfaOXriFXM50khZv2Y/hrb7
XuT2par0qaKI+3E5HLgvQfQLwaYtuPCIFbEm49jJ4A2LdGx0kScxaeIMQ3LL
1mUIkWYlRdQeBvfVtn55WKWbZVXpDQrDrhDsDTMbGyhR4UM2nlWpKYMZ9l0m
ia7szPd2SYKBRTrIV52veh94SCWqWobPWvjVFMSofFqbN5DG+fneymE60ge/
+OmmWP4j92LtonbbIOPpCK1TYSZ5OE/rYsaQydoWxOoq3iTjUggd2QWHU9WK
LMxdSOT/IXCAU67YgQwIBqXPsJFN8JK7lHjuRbfrexoFX4Hi19ezfn6+6nLn
WTRQ/K6OzWLp7FXB9UWVJXN5s1hqtzhmCKcLjDCpazJS0kCzPdWyS5s2wdZ/
6A4I3350A8/Q3snEAnDLZ6/yU/ArQ/lmi4ITWEkD1kWoiYNdGiTLqGVF1UPo
08TCIlO/Oug3OCMKYzfnt1Ia4Cfi87olD1Pe/niPZfX8sYld8PECR6JdFtUI
NZ3b05qdtXRkxGgdeUBo6axueq1Nns98U8muj2jigxl9a3l2/okWElt1GWS9
tL7BrqruvOSylYqD2lpZHJf03z7wgbzBvPwxgLmw2BllNBKeTHYB6+mG3a2E
ljwkd1Fp5wcrg3Ul7tflIeZHHxREiLKftYWle3x0y2PKpbFh/joYNfN0EGi6
HCNvogM9x5Kur/HyQKynGkmenZ/n3piBvJCqiLxfz5fVd2CrJHLnq4rX9mfz
A15u0G9KVIUQW5lE20aDmzzrNA7As/KT5lWlnD8+ISUSu6WPCpzOt5YUAuW6
8WvM9+lck+fuL5omPUKiHKD9USsM2QQnUD56Po1t2DvwcpDNkRy7SGDiwCgv
Ps+tAdd/QNxtSsypQF9BkEHRkfCS9EONSAJiTGe8UPZGE8cSiGYJUC53d9Ey
h64hqo1snL+8m2HovAagASe8JuwKssBK3MH4LakEX7QF5DGEQkvBuAu3vfGu
qFqvekwmDjVPIDN1NZOhPhtUkwPiuQa35rois8195SL9XDcWsFy8/RDmYSRF
B812FG7g8daCecafuK9DkScpd2B8wicp0gy2K+h8HmXWZwfHHl1PDZvSiuna
yeUe5Nw7mVwNJTGYv2Ty77RyXGNOsisoPDUmpLSB+CJpRrgWbagjZ5qmRuqA
cFxuc08yaw5RU9E0NOqxUBy0Mfuvd6KWWQyF7UZNm45JU1WzH2aN3he/YK39
fHBU/E4CtNrPc1PxfMqyKvaNVzIwPw80E/oWHklS26MkRX31mj+7ygssJoRh
JPmOf9PCbhQUMTrdj1fduHQpMGBqFzBgwyry3A9Yw2wIB+xnJhvCFsTxmBH5
zOeRIbKbA9hGtSsV4bwLkdcNdCKZkD0gP1NZIV5VnxK21kBHWvwsaSMTmgHb
Q2ScbxXA1TmgKiu8ZxbbJCBu5X0N6LGWY/WI9PQo6qnfgrriD0uDQf6PeXF/
SicxJSoz7oyp56oLrEnP5krkz3gKwHuGvoScqPwYXxOQCMqWV1hvU6tSCPO7
0vYFos4AQ0huRbh4ijlzIFfDkkOHsxA4zrvszQE5OJwcwyIrRte73qcZTTSc
Ugejl3TxBCNKI3Pl0vRCxUhXpOQA3KdH4KrtgG4MB+xHcAFBDcaoi5wzsE1f
lTXm22Rx2iyg4jy+C9xPJtCiU26JbXxTrDNQT3nB/WJcZSiKTeVJVcpeRi3l
UEjhZz44W+kc2Ttlc60yAUH88kPwR92lc9RmUU11Oxw5PqDrccF/ywf0cZwJ
XE7MFuMPvArWQqjWrRzvCPMERHuRe80IPSi0su7ZKVonWub2+7hUGOkppow8
hpq6nYg8NlC2kBNfAbm+dsvcFQpuVobp0YisIZ56Z4djNRPezLZY+VV3Xu+/
j4WASDGrfrJ1DuiAjRSS3smUWSANX4YjYDT3W5ZVKOOjuGeolJ/0uAuJEDVE
Z61D350e1ruU0yttVduBjaM/La5iFOapNhMR+kY9FxgYnO2CeMZxHgKoBhuI
RRASP4g5Db2AbNjFAFdo43cE74sUAWpoc9IZiz23ekny96uZrXYIlyYSLjev
b29T0dN86oXrzf1rLz29/O7ng8WI+Lz1vBMlCB0u/KHwE6KLdMfzQk6+baKz
unD8sn/EtnxsspVtFP6tPg95LosVUcftDNqUseHgjmw0QM6smOAcN0iV2yqV
AzT5oeevJUbw/BW3e7aLguNTIKDAIbhWCXi/9bQ5CgQth1ZT7fW96XWyBxZX
b1/96tUxufSEh70TJD63/I6d/xq4F2di1MvfAzC4RGWilnQW5CAc3ZAHJyav
2T7UatXJvyCFHo+882kGgOXyiMaQ0xumrEZpLzN/ghFkbNhB3gjcIKFA8Nve
k46tS7F+DiY/SDwGjHQDQNh9s/kMo6QH44bBL4y14sOg25DJ7F/ItJhNBeqF
bpb7lnQynwdhNvz6DmUJWRv7H+O31TzSIhA5KekDvl3mRZdfNJs6XTNfqNup
EMW9IKnthw8WUll73SNPeGeF7b1eF/9NI35w7N0sbpq0wup0NW3bP1G1J7Gz
tjphcfDi4wKwfNJn6i3LE6WJLm1ntMi7bXgjIlNOhyltyubNR03J4ZqI1b/V
3cr/VUIIuqg+WJcGnScPnIpNqbubb4YG3r3sOxffh+kdV+QKHdbnC7ZpoJAi
2B+bogH9tL4JYZXVSNddp3IzbrDSpyr65aJY2sBhrYVUqz6o95Qt1GjmaXnD
QAEAIMhroYQbFEECWg51Lgmz+AWO0wiTn/jcYisXa74sNc+Q00zJZDHgCJVU
g5C3Sf1qoXR78oeV0cn1QwcZWAtieAb/YNHBCQ4HFGvQ3R6QNQEGTweHsaVh
GKQkKUY1qfb+dem5gEGSDD7jCUelPID4K15ACB+y0TOh67je/ePiGeqh562m
/eqkF2pZ/5MiVTkh/xofDc/4NIq/yTCUK3VHmKi9dkHkxni/NLxR2Y4vGWbR
ohzfI4dloNOgo8+JIpZh3Ry+irTf2H3BcOAFICQaGgNas2GJUvJALiAw/c3v
AITCOq0ZR9dtPMm4PjkCEwJWqkXo7/q0Yp3PJm/5m7C+thI6Ihr/o8qdMHBs
wAP5io36VFQc62GQQbY/pLjjjdlBXSGjg5/QDugArkVANinqSwX+uC9ifJNU
JWkbzMoGbcw+fkG7rvu3mjbAtgbg/j4muXA6gyGtukbg/WXyxd1nzJiR9ede
AYj1G9KhchhLm+i/KGfXpCFfVcncLzp6uqubvLydc/DxsCtfmB9tPNN98/eo
YbWmZYjHdVZ1eVMv07tXq6Rg9LW5NYQsFFzUvDu3hYxhaB/S+jC2Q9dVFzO1
aMS21szmANw+2auzHrhcA/U8rX6h95kGpr3Jy3pi1BUGQMjN/CAFClo9+4F0
CLHO3vH0asYJXtG0SheskHgsqTBC4kP7H7ooa054xXlvg0pJy8VyEHBoHOhz
804VsxOmZMOycAIt4+2HRniEOKPOyohqTtuayBnY7L22qN1ObPHmksZdvnF5
8Jrb0r/OXdUFfAGr9jYa9X1gGJ241YcRPodv3xd05g+VcXPV0jlrgKAqmNcI
JS407ZvdO9iwJrjBbMeu3XMARl2PXdh4EJHMmpQWBk+hU8f+oj5E/Zkw0p/p
Z8SNFVD2PDku7HUC7dluqw2oeMfY/EUA0/U55uAXpYNLNLvKWCksoEku6qG5
UGKNdX7Ef18XHe1+Mf/Swog/+3bgDBkBfi/t9xtGL3RMKWV1GueJrr8KHjs/
0S8GP5e7z1cDYi1Atjg8ha+6EZAzYO/Qso7G2xG5she4Tt6tKBz35zHnMov1
o/iMyF0Hdc+RxUAYnTanyT14TSYU0GP7pCI95n2Zx4mq+FtDuxB8w0BtExZG
QL+LTgmPzuJWZZRagqPdpv8TEpSFSsFIJYPMe9zyHRruCPT5Vj2Bu9UAcJ4q
wTOUXqqtxv0wUcwe/c0VzGctzW2UIqr1wWImk3zsPC2oz4MobLXZkBBLgf6/
n3Quds2i4wPMgqvyatmGYAeNDX+5PWCwU7O6OGJ7e7eGVaqQXjKuwKwYuEnK
AHeL7M83LXscs28ELGyesgUQdrCJd/LYm3BMyn3scdJudpCBS21K8OS+61Ns
1NeiX1GWl4RsoN2wt9xvyI0hRszMuOl/4V0AurCjUqo16Uzt1OhPoj4j4d/y
mxMsHZO5TZYfBH7A2o72K2V0GvPDhM+9XAypFqCe5iZMIu6XyE8GrWhFU0cg
ASZ04hy0eYi6z2995Ib4jagHS6CDmxypuvgacyTDRQ2DYRcKaOqOpnuyHfH9
bkJtpwAAnH/YQMSjO6EHub8shamKxHpx+PJc/L4C14rMkLyHVMmh8UvE1hfq
wJkhLlVgjg6xTarhD5H1Dvm/pteH0jZeRgwOWppzs9uwF1KcDhdtU3k7f9Ez
69Pw8lVU2uaTKzyMLD5BF+cL2W/Jx+3+5RqBOuudhsyQhuGFmDY9OgPgwjb3
JMn4wDAM30DqTytsUUxM5Ar2hY/S0bAcaQ3abMgqfeWSlcbByoQfAgrhKlZ3
LkMN7MbkTJxFmsi7tGZisKvp2A3dGqttmUSUxYTHrbf4m5CY3efoiIjF05wT
tqY1KFYLETPP6t81+D8Kzft4PFAPHSjh8a6vEvddp5U3w6+lz47IMhazWdxu
6Hczgk9R0rtv3TYDbq576uEzwXD+XRJbIK4oGSdVuS8NkrRlBTbBxFZEjOM6
WHtoiKSONqDIT3sHf0T5drYtdJ/TplAj+9vuw00utOYCbBbzAgjFb1Jup5OL
8R+Celh7aGIDVDXvQchTvFYqCWQyPYNshbJWvwyP87e6DEpHw/TQ/0n1jKuo
2/DQlnfWCzqQWLfDqHXcPbxxy2NU3oALmHkSTAPu7DxRjqEzImFFoim9zOgo
EgEosflYrdLpA0jA4+OXfdf8REuyAzTCKraD/E92n4oQSAxDzDwHGorGdDVg
xnCHbBArXsckuRCB/G5lBJtqlA2H88vOdEdfQD0/5GstdIWAQoP87+12BXzQ
POmFTtnUAr5TQCPQmoNok9iX0cjvBn0QfMHfjs9QPb6GvIY5MpdvV9y5pk9g
OrLpDtt4P+OlFRImdt3f/Nan57pxD79jl+qzCo8zVQRmGwMDuh2yRpyTbLqP
Wo/NxTb/K91kmPvfO2MqrMHrLjsy86bzU+/nk4kVXvqI774oI+JFO6k5JBnl
QNDUKXHHsYYBv67Mh69Z1CZwOOvctvl71BZamnvk5KLgrKPWlB12Z/+nyIKp
tVDh0h6d9eqNJVJBvb8C0G0hRUmz7L94/wy/Qju0gXn994zHFU+bTvye588s
qAsW6AHm0lkwmz5L1URctOO4vcnAWtSBD4VcMmp6X8KPfx/kuL5pnc4+jhvK
Xml4QBA0R/evEZn5ydM5b/wYl6fw2wkwlpN73ePWDokBlqoOgtvkmUwHXOdx
ZAinO1zymJ1yVbdEY02JvDS4PyxiasnSwDdReKbH2w7+FpDKm3Kl4WEGORW4
r4AiZFVX2Mo8ay4kk0EuUWihOY+3gfHpDlAWZfOxTuIqeC4mHGboTXYmVlQJ
0/btebL7aiD4laYpyQ16U4px42kc89THUyrONVcnH8VQK1nsUlPnbJz2Os5x
IcmvHulhqIwliae+qz5UPlAgHFard0CzSU22RO1cbUE+YB6oSVHKr3yVB41Y
LYUAvfHKpczL6HQvBtNToPdxUr3oAugon4K5jlxSkC70WPLR0rzfSQbCHAH+
k2mQW6oEQcO+Cc4jQNFTAhZGSYejy4t+OaX9RXR0hC8BmI0ggS1i/Q6t758s
6wTOKEC5L+htc9gnz+WjvP7sXHBUqmxq11o3MfGiCBf0OtKwKCjCXRyU/1cg
el0UU6YBd9+aTdseC3WD6xyYj+AttsoB2XVm0KFaEJtCtOcd8PHZWjeI/+5q
/IsfBfuBgc/jBqmtPYmWr6KCsgAaiiDI5UIZUrzoEVZO+FtEhKxUCM4PUcOz
VM89IRDNrp7yJU6TrbRTeTbYT60Z6MFUDgz9924m1n5UwLMZM1aYmCFLcGqs
MWz46j+77o+p2ZaHoRQO4Y4CrT42yfD6hFC5pT1qALfZqM/ESP3EKtGgFq1v
IQNMNiCBEKneDOxL39V8HwewcnNQfJXfSm+zDpxkANTqsd5iCmR1AYCkMxEK
CO5LZ1z15u4L24w4De9HlHjTLGrDpur2EICAQZPuN+LXZsPJVIc07F0ns9KL
Bl95mGBNAl0OAm9vr+mzxfd19CJbkVSKO4RUz4XbPKlk2dpr7MX8ID7yULjg
G1EyKxd5HtopntwXtlmOtaSZb7PJf+jbUfwWrFitLbzpqCC7yqDJN0sdQsJm
w5ws+Z6z4AoJK/10j0/54iRSuToOOMMgS69KMWTCyDLgv6ismUdOxFawfpwI
98cRHaylJxO314J0O0mVhg4VnV3R/xMg8GF+4wk7g1EI51nORYeuaBwzMpR8
QOOB52OsVzdybESWLkSCwRDYiSZLBd0xPuat3NvCx/m5ccCBJ+uSqELFEuNn
oHN2IZFV/duIbSLD5TJSbqLPut6EdL7GWmLjIGUtg7dvXWfDRLsK3TstaIPQ
9yGr4r+giXzYU8dKFeyAW+csicpWcKNF2E+YmGLLWwTtu1tFnqfcit8a1s/h
0L9ViY5Ng6eWE4u1J349jdote5rLbNQO4bL5EuDKw0iZ0v0rTfEKYI0d4+Y4
XmdjAxUuA0WibMnF6B3Tvie+XeC8z2ph9/lZohzO1T5O7x9KEOsTXOmzDksC
r9hH0cWV2wwr8chygcazHIDybVEBbBeXcAhnR7LzmDHhZ3vp0PTk9RlAb4xj
UMmppWcKnjRhmBw8AVDckzhbqnFVJO9nVOvOryuysJyz/VkRxeTPOslkgB03
00Qq6ASZSAP7FupGdasvJCBPV6Te9V4RYYWvjs5aMUGzii/GUuQnGihCnMjW
YNV8feFTUGap5Dz49JXppfdmn4c0k5GyryIy3nS52o+j4B4IlAjVyjtjXjK1
+WWZ7QpsRw94+wk2kJKaPA2Rkd1a2h0i64HLKgKAVPzLbfMFsYfKCICec4Pp
+zAOmcv8jXJpJvm3LGuqv8Y9cexmNJHdmna46Die+x5Nv8yxVQDGzpvuPWAD
rT4spBbLPJNDSVrCNHMO5Z/VjjwbTk0xYu1uLiGnCDBKHbV9LfYjrkCemwS9
UiYL6PpP3lnAi8vMAnHAX5sSXD0spehB7wPmJzxEpYn6fWTd4ReV1bycJ8Gc
q/lANqaXT0gshqtzhzEx8f3N/Rq2DT1Kya1VPa/uhmXk+r1SouQdI+Z+pnF3
7bhlTbVJPLx8b2Zkt9gAllx/HI0zl7aWnrX2HUsNfL2Liys6KvDZ3O9hbvmh
uTTu3SRVWQXRskXBeQxDwZvHEowDboQEHlj1hMOLvqjJ2s54dWNmpDkx1u+i
qc96pVk9/11XoYB7U+cDBZWojQpaEYVPtNbVbajDY3Yx0lRrARtujZozy/lQ
c/nA+9XmRb+uipLOZV6juyAucofPBTtF8z0smcdXryW5fik3R6cUOxvzsXyV
IqLRif1TqUD/Ab0sC+4RFss23a128e3/qBIP49bt1O8kjQYdWc26IU4Xg8Qw
KRMVO6lVv0aHRdYEWj0ZUENFv+ZxTchIiTRV8GMl2ehzlCynhClqHUUg81V+
OipWohg5msnuhxZbZMFvt8H9BJ3oAKgbxw8V11DSW0QC5hZT2pGnSZYdsJAu
XOyQnnaS23PodEpIyZoO268FasEfd5ZPvDXCJGMNDJ3/LLcnoECtQyZiTxmM
gtlaCp9YoV8meENV//L1bjeHyzwFZTysFClfkSO9jt+J/alEgASj1KZmWJhE
i8l3habkE+WAsZBNtWGKYlzIuHdPm0bXMkLpwlWgjJfnMCRboSSc9KUVafEl
zO2sfZBUahWthCHpnbtshYxLDb4e0wfTNZaOZP1X7GqYb9gYlJnR/j1dtDgr
sG9aT2P5g3PxF26MRyjAoIBdFtp1qoPCWFnNmyCWjhD5pyQ57Dry+ES1UrnI
u3V46sQp37M8VJ5ZC/5jfPgG+LXkmXWB/icye9UlDPjhhbcLm6jic1vv1P6u
36I+mUtm87nJMoFmaYWPHw7k5/52H8wQ944w1bNrCZnGZgaXU51IIPo7J94o
qBlAk9NjD4dI/G6TkEslXP2rnLjeMS3z8FGJsllmxhX5pJCDAaB+qIILYz3T
1Lzr9XvS9R/dX79S5iQaLAuVB6FPejqbxXoJSSxtNZaYrAFYCUoJXcrVbrvN
Jd9vBtmHbB1vjUfbeNpmLCa1Bi9xThRwkJfSWcvMTcfpGEiJRAdPp6nPjRfJ
hySPJBrMb6v9Ttlf12ygJfStGMQqk9w/n0vTDB4HkT4AjIaM1Vw79/+v+GoH
77bez7iYefLkjJv/laGnkHKf+nKwaAyXs17Vro4QDx8DAjvT7avu7+gXVBBv
1NXb6QqAwr9kjcHm5EIP61VSicgrg0GXTXoi3nvfoOCFU7xYe16ISip9v7mA
PfI3WYaz+x0JZPwPao9GC9ceX4fMRns/WJDkQv2QpUJ/AuftHq3II8HcVIyK
vcx2+MjTwv4KsFhEjsD55jKOaFu57qee2WaBiiixpv0i0xxAsn+DsODjVp/b
RGawLbsfoY3d1NG6OTd+4AHbhR3jMkZQr3uH4j5qJijpjAi4+aOxM1gZza9U
K27HgF+b2VUArLLQMDQ3V7tBfcI1eLBz31Yw6dRHMpMgJZgPlW5uG3n3kftt
430Apk2RtsdSvV9yifEUgrN9MtK/YzLSqeMAW42IaJeWsDOVTPFxAr7hW8mU
AVzJb+mL6a7KVHzH3fuxl4fN4LJIMdBFGzLwZRz+sJqmMzUO+dTFWpcccNhV
CSkT6WH0FhUl1cLITu3/7eoe3VEsZufvWXzRSCFAY24Y3E4ZQE/EPAL87e4g
lIIV1j3NAbCiQwgUQx9zLFwHPRbfoiYeDrQTm22F9SsfqsfVgp6lRsUVzHUk
EEm83BpcZ3znj/ef3JABk3+BdO/WgxqLO38KKsaxM2rwQL89ENBFiJbZx54K
wEzCrKVG4Qdj6O5MlZRIMxdFxI+QyeYiPDRIcmx9cD5DE+CfltjdRlh/znNp
sp7M7AHcj9f1MXQWplPFGhMpgJOyYNix+nK4KK0mk5cZw3R0IfyAaZAIyUWr
PqWIVuB57FfIi9pbFoa+8ZBztENubzWjYRU5d86FOGTwENUkACt+t8KPj5hI
WxBz0N2Ye4P2G4QGAyhoL3pyeUtX07/chUHRFymoQ+QB9z5EyDeUijS1ROWE
o1up8SOuxz5H6M+liQYc1nJhEVfkZnZGNJZu75bPvdwyfoKfzRK/N15F3cvz
auwse1d1bqlWoMT/e5a8YJsWKZs3l4pCrKKtNwEna9PomV4H7yXfSZi+dOOA
LdcnhD8Uw65RJSDLkTempqUNihnhBWNVRiy0ZSnYRQs0H22ngcecvSbQ5on1
YwPkCW+r8vOVqE6tpQXFNS/yXxFXK8g8kEq/+XO2G3WnkM65UOa4P4ygdCAp
6P6EuyWq9o2865DCiGqZvaz0E0bGp+h6xDGHCb2/HMyBtlHEN85gr+Mjkt9g
+u82FMeSUVahR8/7/lhZelHhSlomI1MwUhjamQcETRTjnfJ5y1tT/4T2GCJ8
t8NRvjkCzf3WNHcxh04sJZh0HeeC453UJRDDhZQY7TFshyhVCx3jkSNcAHVv
v2rt0pum39ruh73+uNgGerrpch2yCqN6MFStkyyaphULUHmInscITzg/ymVq
afwR77IZ8RKUX5+JijNP1zNIDqZrkpfznINv8m1867LGOmBw7yiafPDdbBUJ
i3ImAhIOIsnU64uM4V3peh1fC1o3s6yXSmwr6iiGMdPoeVOy8cAenx2zXF52
MxgZ0MoimBwFhAvnIt/cMns00VcP9oLPbu3m78RqIdctv7beYRrQIV0/HazF
5vXu8q0vymjNCTpB2fhdvVSQamt8eqj//1Ypb8aNVeMX7aqcCoz7gpvPW1RM
1AcsuV1yHpetPP5I0xvi0WW4C8CE4SV9hFFh2P0Muxk7dDVch9wuomifruYa
kfohhg67jSNt5ctcqf8oYj6tGIr//EmziOCNZEYZnxFKqDNi/VC6LMwUI3cJ
COtZoYjDV2t0zveXZJP7f2ic6BhHH+ZIb/moepjVquiPqE1ZmafbqSiNqNUh
b+4lfho63651GRvowgAUl2BnG1ag4FwelUtZjFznytIohC7sQHA8SEVQexSf
mYSiET9eHHyAYWl142DbfuWZ8G1LhDn60zWPL7BhMv9G5+jnyAuPvdmL1oZ1
JCfDV8B+ENIyZ/tV9uuYHQh3cubWsOEB3l4pwsuUdyKRyeZUIqYW8pRamy+b
UfrbCjZdrHEsPE3Fe2tUXXWKZRV13Ujsy0G89CjLcFIqVPA9Qb9kTw/kUMtS
GM0gzswWqREQKNK9kkWTEfl1nytRgP8yxwKOrZ3RfYg1k1rbD1P2pjepyL/v
re7A1tWrRQeInubzK8sSEbGvZ74FdNLauZS5kpVy134geC/SKltzWnWOBpKd
fqjRoaIGJ18yWI6rduG+jFNOFqR39A8pyYiqAIqJIrhWnUKMC7cRo/hASohx
bRqD5PsPbB69b2S/erOABc10aFs7YSUuNktFBHkdfdk8xcLoKN2HqhKwf3Vk
7Po86bNsaqBueG6AqboIA8mnlRGRwLFwLblkjSZlqGaqQ7FUlYIVIas9Kaup
5Nk0IfMMQT6lGcXh3TIyLUJqbthOSeYRjjhWwjfzkt3WIZLugICCpgaQAAm8
PkaZnVaRPPUpxEU9kCg2DnXV9Fh7cVtjpn80TF5Ye5qF5LzdAPPItQhdBXW5
ubBxfmfR15Z3KXckwTU4v90mhL0AwyixI82IZHJCpq3KXs95pN3nvaNqnow1
I6+o/PAzbeVR8dgA4uNR6Y8yj3GeQofNxXHk806ST4HyD78p5Z9PQstqUjXR
nfspgm586j7ThJcuiuoIOxdpQZ1ZXNmnTld/DAzBtEcuv8A7OW15Ai0et7eN
rejRT2s0H9DJaUuSqnojoMikEiuWN8pgxCgYpB80uNQC3BdFDqmD1DLQfEMg
1kEO46V85XL/bB4cZOtQO6Ftm8Lm9Knwnt28UadEpWp9zRVuoEBXOrTqBCGw
hTJMHAWw8L6RGKT5n6RZiD7lP0If/W/hLDW5/Jn8bjvDDIDCFjLlepz17Kbp
pyEBAegeeuEnAe6mIkL1Fj3BIHqH0OZi4eU88Cb9CPk4OdVqUVCutfZa+lFW
+3Hn8AWs3SCFS1aFIbF+gGhUnlO0Ztcmh7Q5KnyC1++ereYFjvvDzNefoIun
6DNwRhX93xaboRbhujo8F7qzq+Ci90bcmsgXu2PcQuF096IERmD6DdVE/nT7
J+VjBsK9MHjFmVrKUTvdbgKQr+i86S3kDQ/sMQZW/9tHE1ArxqwpP30hkcGD
CirosMV043hQgFowvqEPuPfD6lpOjQ6ORxgle9He53ccHPhrD2S7uDQjvZ85
7IIp+thuugV29CoO1WnH47co2NlEMQ+V0sD+bX7AC9JLS9wHTPzbrCPSBZxL
3XewCQztRmhkfJugtYPDGeCyFBfTvRt1OX8VVXXVFuEz/y5YdYoDeZruPhXo
eRbaBiV//OYYzPZzVDceL7c9YdJprIEBH/T3B8sUjn/uUGNXnF5RTLzfQRcE
7cGne/2ijfrXJoWkqKah52vWgTk+kMvnqfrN8wAlhxY+MzdS0FWuM5eX5qKl
d9s/TrLPd+Uc0Hz26nSihqkBpL9GMfOaMR+LoYDSk6LTLTiwuDbV4wjI2j3w
TNS/3tkn+j0w+c8BkJTHzB94dHgda0Ne5/y6Cjx3DoViQZizIjhfuJMebQ21
RVokOLzKbUlr0tmpiPFp30m/Yq8uu8n8PfWysM09TeX0fZkBVUhwr9BrOK6y
7BhkjKsrzBXCd9seDMUuLKwN6fVrTJeAw9Hd9vrtPZqQdgoHhJW4UsY7EDYD
z7/RMY+6TGJX9IlXo/8pcTcf5/at+vOplkz2ylMDfZ2eeovOT9JgWi0Fq/wK
m4R95ohC6g/4U8eMYyMqCHsPMQQwO3gqM4K83fcHhlceKV8DYN4Y2WWMS+qd
tvXRFNVY93JgdccfxyuGnCxcn61lKZNTR9VPFzDEE1wEHvqJOL6wGo4sAzUa
zM9oNjJmXOnDHrFNibAWvi3ped2Z09TrQh7FIsqQu1jBwM4H6d+O5C3HQCSo
WgoUt9j3MNs4PF7fcpfX7OLWKYGjXRvNbFH4nY92PpXxUmf/4sAPvjPyo74T
oOVn2ipKAjmYD+hsEkDyxYjWe0Z7ikx0P4XPoxY5/JFdTnChVvuVFc/Ux4w6
s532+zuQjkAHd3HbppB2duMs9XA8PiGVgJooPxEcQIIDJlYVP6jOdidaeLCa
EKjkwFvs+hsP/PI2xoEH3FMNDqgX6wQd0JTnPENrEcEWg4y+D0C9JW0vz94/
rNOS4myRb7ZdN3rNQxzwSOddTz13oGCnjM/xIGxCmeZ438wF5Lij8/9dD1Lx
GXCWUoZzUt+dqwEryfKWCaelPDqIYCpaFtHpjL0rLTy9KByusxxCwzQmVhw+
aQ7ZSb2oyj2Ov8peybzn/GzO0TgtIjlT9ZE3hpWmUoj8tn+pJj/WcCYOMYFh
HzkgdNCg59bNhxch8azlxcnLvvLv/AeTVFmxW9oXAGr+G1fKFiwgHgpGrRnU
t26TceX/fSfF6G+2Y92yRIaxIks5HKt8v/1/eL4dgLpgMWjLYd1KDlMCkDTt
9j+clh3knkl2yaXCjGTuM8L9VJtf+h/nmZ8FCP1ju4829O4DPmPbE9no9VY1
SwyFv2zkNmqzEdiTFNQrb1S7oKySbz19qRru3sfkZ/TmFBirsrF94EbQBGfG
mA38ny92ro+UeSn3Lkr1gszPE0CbaZfVxKuu+Ps2dT4sQTWOQIERKvrKV0u1
0/OW68r0B6flci5ZqYk+B9Cyi/ST+J37Q/1g6y0ocxaiSTmHHNhIbiLhcxp3
j2nwHCB9k5yIPXR0gjy7pe7t6Vap0ztb+Y6rOJZ/Eq+rfYjphkESs5xpGF7i
NuVC4nE5vinKRbvcbiritfT9jMp5gsfZyp3T0UeASQ8Rc6k10ahdnEZA7CK5
4ZXMVwp54i04dQX4BF0za8UPYtPw3gCNaQEC2qOqqIvCqqq87yMWF3rYI994
EK9M9ogXFYnFpzyeVlVw24mFZJGDJduVy8XHWnmj4QywFxUdxkRKTIBsUnRy
HH8xVqdhTrd8ybMb8RRuliuYI63TwsGHqJT6iF1jCzY70ddRvXXEoCV2Va8N
Fo+RAxd8Zr6IMwvjbOtCrmY4C88zD6XuTBs/YQYr7u1TR1GpsWLAvr1OSsSQ
5z2Q5MDf1ZMt+YtSgqyquHOQjKG+AIty2QqrxKbzfI9CQJF82CSMMXp/2k7b
HzRsHsrGVQUwuNdNwS3+9+2WzYo0rINPVOpiOhNHnXX9xz5NGmzrWdw8SI8S
D6mwFROexC9M+t8ZqvqMh6B2H0x0eT8ZisrwQL/kt6MA2aHFBWbdxiTM/5wL
RJFXHduXPjYeN5hxwSuKs6IIaJNxImxyJeEy7zcl74C2xiEhZrmvz5FAne+R
IcDECrdlrS+HTTVguRyVt3ovWOLnxlko2DIM7y54ePfhvjGOYxQPacnW9f94
0h3HJpQeOPSIvgOY/lRlwqtDbez/5MtJgQUvokBwkLQbhqg/c2RQDniR9BqC
DHU9uUKOme4IgmiUT2Js+6MSTNvRj9h0bPFlodQJLKqMc06UBr1+3v3cIf09
PYE200wBj9WEJLVCN8yo0PvoUnHCGTplFoRiosWXvUjGhANDZObsHnqdxRrb
IkvxIaduXGofc5KsbvZU4NWtU3WzKzbzMrFXHehvaZKHiSH+y0JgnShIFiDe
GrJQSMmdW7IW0oDpNw+yioyNvEHAM61fqzENXUj5zXHJdl4UWLjBKNQKraOY
YF85kO2PRij3u1sIMjJz8W50gaLL/CvDrRouZu6BlBb/rGqv6MLvQdaSrIoS
9bkVwYE5jhU6x06ZDT94RDG9ONMSEE9UcdfPN8kQ5fA9E/hurg0IB82v4pzj
Q7rPqRkaYdL2+7wZZrpoY2gel7azTWRjUepQ20uywNbDj2lQVe4IMil4JpIn
D8aSeDJSU0XnC2O2eDHezkcsZ5SlwWCopgCnJLIl8KpgfQBrDHW+4EYtyJPx
LaSwBTtcK2uAMGJlxESuLzyS/SkpS/XJgfwZ5aaiuEiKct6+iAapArgA5iqI
LhpXhEr7fHdmpV81n+5mFWvCX/xp/8vrnxEZ1Da19f2LCLUGpGYMZY7uwXTG
uPKNqn6uC3LTAcYRq4733d1aaXDtVL8MWiU8/OKrIVIr0g7dog5ymlxVGMa+
9T86vHmyR1jIRsRPUmXMm3BLkQUlzLmiKWAyRn9FYFCpTPbM+tDkwpDpahiD
cNMKFiZK7eFhFjYY6ToF+ym39673NIotk2ig/3E6KhGkotwc1IGpXajsiR0J
2W95VSJgSIJ6zGzBJK08/ptWmcQYtG5xzGPHTi8I9VFDUbHlO/W5OJHoWC0i
1Yhj3Lwp42B4orrodr2siaDU6z/DWTEUW05bc2sMZ0U2ZVxZukyJTSF+cAao
eBYc/6BFGRljdEv2yk5HT6kXVpJ0vnNH923ScT4MNYZk4MXATx0GA2RqV4yy
CdzlZqMXFKU34FksWdyDckRVDTuS/G12mORzdWZj7CSsItAQ0l35mAw+NGqQ
bDvo2wP98NAVDi3ZCfepHilyUHj9DVUZFG6cOJ1tVHSjOp3qXuAkY0CuXPve
TWy5hs0b2UZTIOFeb3yuvmABn1/fN9m4r2oodPhT4cCpENSclypZrOfysQAI
m85DqtbXQdkKYx69J6d6GZjlyu2eHLUz0uLGghqkRgFdpF1INHG7/dFWmo/Z
oSy/8z0ocgGhZDvVr+Bp+ciPVmoYBz3zT9+nE6PQlE3PWb3gX+wAMtxQjk8f
bFIDgw/hwYlM9MOyLk3o64GE9WO90eiKciZmqEXS/m3C8ruReEvCH4vPMJSb
yaOcTiOdIaL4S7HjLxa7O79e3+TN1Kh1Y+UCK/TFZSNKt7HXbfNBdaOLBCwr
RbjkioFY3rAk1zF/s3GnugSgRclBdriMY3LYdR0te9dhXWGBnuzlGCSDQ9i1
bXXSxhtK6XPAXYOSXY4bvCiiiAGxoWkGL6RSNWCkE2TQgNRdnnrsJJtwpRM0
VXhvvguYvcGc1bWVx2i9LAE6MsrT+KiRJGIq+qpcL7hgDnCqCRDSB6JY2EJN
NF13DxGOXzwArZo5yJ04zsjFMnoq7kf7yUMwU2M+2Hif6OxCWgfZrvCr+Ixf
ocC1c/TdzcBxQAElFbINqj2aoLlxq39oPw4AhE7WqgMaUu+ef0w26VmRs1BH
+J2AmttHs//PcyTnnOb32a305ZdBFJ5Vv706uTjVkyWhl6ZTqp6YWGGJAyHE
S7EsG8udsG+mvuJk5MFARD++aqMpIfn/0fO8B8hil92F/GwPD7t+kMx3WOCM
GgJx+JQCa+W7S9VlUSCtLshTDxy7hA35PSdMkhCbUwVZBNUi6aPwiZ2x66LZ
eghqzezKX3iA/l4UY18HbeOhfZ8tI4pxf/3Kli3gDs2KGMlpm2Bcao/sylKB
UiiLs5s4fwKDfGGHYRogkmIqUQxNsvI2owy06Y/TLwsT4CaOKAICZsAEKv4I
jzvigxH7miVmUgRtWrUuAZf6L4H/jZlp4JoakmY0/fQ7KkQAjrzcczoH/ju7
9Xj7hdsYxAlcLoglFjO/v8DJRApjpim8tN59su9vWDM2QCa7YbfmOzDi0kNw
/f68uxxvVRkW2Mf5HZIgStR2NsvcjJSGhu4ShaBi/6IWuwQpOY9snj0zDYaw
KuPt2+uLK0hzOpz2Tmyc2+vlYm3kbUuJCCeZzhOgs/y9NvoCsNSgfjhU5IRT
8mCwn0MZI8ZMHKpklwcT1UJHExqE2U9Xd0apcI8CvNjDzn6V1V0zIy5VFkyq
Pmmf8e7kIUUITdc/4r11nFzP3Rhn9B/8ertCltSnDtFbKmV+i9o3c9Ci5ZyI
GU1w9W74YgBlQ5K/UWvVr6g3UgAOn6Xg1yMD5nrKxHCKgQ/gTxlqm3hE5qh8
WZ5uNPvudE46bAwjANGf57MoH/VPm1qpbCHfG2oFts+6XfldIgxD5Qikxw/C
1YiXqff/7vCnj41hYDGHL7e3mUCPT3MbfpJyelNIMSVnh7JDnNnMkkb+rIp5
og16HHVHKDRJ2Y/fuRR0VAXE5ZnhI9YiClh37F1dCYBs+re16jDF+4lgTnQP
7e6RPV/VYvIZTo1HLszEU8D9EkxsTls7+sOK9PmFfN/yrLCcFvE0oaLcNxfL
QDs4hjrzHa94NxgHWWTPcl2TpC7ez3Zgr0K4dM18MM9gA1M0fxSaJn+a+tKc
0Og4OVtqC3r0kbcF1TIgBZDCAgXi9+ju6lbFXtD5R4LaZq8pbTNzHDx/voDu
Ce16HY9u9uAassjWYhhI29bDNdUs+tSQO83ILzw2YTZIrt8tSBQ46FSKEcZQ
UG+qNnSt4HnWEgqfGOVYMXWr4c0NdA6TtKKHDaDK1BfH71JjRjbtr4+SIOfC
yQ7pB4yhgqrKFZ8hDMdXxQjKI9d6V7tyka/O5C7gdQV5iE8w/zKx1a1TB0Pw
jO3KJ9Cr+mIy4RyeK0JT4I7Yv0EH7qRkC8SyP3QMHaTisNG5PUnVrTFAnrtS
irK4tVzEuIw1/Do5iG4hZZyu+LKITE4t8D1TsEokEzx0XM6eas2FqPVZP3k8
KoHbG+4UQmW8vlYHyAnvLOws2YNOsm5+dLAMgjw2dQXjFug48OUo7Hk8G2ZL
jrff3wE1V5sMnOPvah2D+yZqoe1wr70yBV4c+we751ugcV6Po9q5ETWB0rej
l4MU+SZV8aegr/TgICrek5Dw9o6iIOpMo+Sq4LWipzXJ20ASkXamgj6dECVf
da/1H432tvhT6G5i1m81203aAKPChTwTOinEFRHytjDohSUiuKBFaGourq5U
j7N4IigawUEiClnrKBb8XE4k4hmvpMQHyhFaSlIzZsKJdyPJYgEn055QHR6d
4c5QpfCLw91ANHO74FxLV1x1sPYkVyAZfHvp8RcbThEySt2+DvL6DGfMderK
sTW+40NwrqKQfEojbYdsblMqIbtQ6J2HEBjZzCGlUquwAGSXZpcsYdIygi8A
UAER3OGvQKKfETeC85yOfI4jNzkGPLymknlCiZEVBR6bIrm4ASizQKY168Kl
rXLJxp9Q6LUHTSLL+FPMAtW5n4dVROKt/5p5lO65TqKcE6LsJ+OeCJyZM7il
cWdW5bacZu6/ZxB9qiOcVC9fEHzvnFS18TAafbIifoMC0t0P/zErT3ezJmKq
rP+tkBwu/QK65sbYa3HCE4a6VNkKENBK6JtjbS47vI82V6shRluXl7ikg1C1
+wPF4faxqwgpBoQBtrqDKasuF64twYN3imbQltrLB1StgCKHqAjgYwXytMB/
hqcsmABCVM/QKU1NMOsA/ZnfHxpiO7NMHBQF0G8vo72xKb6/1ClIOs+aZ1E0
Czm7tGxTWCuD62+FhmFSxr3QM59yOJOdhyiCm9xYzBmWVely+qmTpzfoJ1S/
sxT7gHOeZ0I1OaDh1LJU60gy7cnBCM7tP4j79o/CQ3ryTH0G7Eruovjl05Q5
KOB/viNeHd/hfWd0XHGO5mwu6XxKYVHNdSE65YR14y8DIkA+zK3RSYG9y6DS
Qp2tXk9Li0drcVYG2BlRpx/l+lKkWdiP1xrKkJtFQAeJnGCgqJXveNPBw7vs
Qh9SMZHmbyGkvGlhrrClY4n6Z8UXwHPBArR61O+5IKGypDehUF5pjx52T3bz
NvK33/k5oHYBMDbh2etCQicctURmsZK4+VH/THxXnvEY6WdVSBb3t+gAFshS
9qK/Z0FbNk1GvbM74lCWiWfPpvitX92Uo87apGsbqwWvvGFDO4pAPB5Trnrq
hn0nO19IKcNn7PUDRsSaKglSw5axsi/0HsZCxGV5iK8LroFVOFTqyCcbeecU
sI8MinWf9NNWu30ZNLaHyQP2/eRsODSZ8z1dL4oPTdyXHXHu8E2O2ADvsmnX
DzV/jJYMpBqQltVxcE/74wkJy4NNzsrU0NG+edVQtOCv/4YkgE8mVLBmn/KK
k7IDEPPs3GRNrx8XKHvmxGqfgekeD40IIzai1DAUgLNCx1RYoh6xWBbJB752
24fvhKHh2v3pvo2T6ucvaYatfFZu5fq9L3AJIc1+sM2tdsyys71VnM6BTP0k
FkA4mgE7mVTnUo5BtHUBFYOMW2mbKVtDFKluzEBHimf4IH2+JyKEKxiVM6mH
npibZO5PnzdNrwPs/QNLA/eEcd54+bcaiRA6jU8TjH5ZlutTEANO2ocfHLUd
1yJ9llbX+BH0ZUi6PqTtNCe9WZ3IyfQ9vr0ZUAz0CT6hGQwhMh30fcT+mcvQ
gws/732oQ8GX1+SzoSIzr4FvrkmfqT95bZb1OiTI64xMsafxGsC0c4fv/UPP
qfPtgv9lySfPoHEDFX1YGu5+t3dHMr/TD1hevFMPUQRb/rxVs4V0MqZP2bMp
sbFb0TibEzLW7Le8MeY4seJtkBjOA2STgcDVPrmFx87rOR/83tyOe5ZJU8//
ZeYZMn/5UDIGA7LRx0oGB9Y+q33FjK49MDCNrhLSG4/cknThY6Nd5BDXKGUi
nAGxF5fBqGO+2qh5hJUOOQesKNclrwk/Hb0CkKxcEu28setTGRYN+XnqFn5P
7RwRCIuLuZsby+DAfsHsZV4LRgCqlcbPDlDjdc5WqzgsU6RH6u6oljpEL5Xp
acH2PZh40Bz1Xt7Ls+jykROLdwIuq3Akqb8Be1GlyKPP2oxc3M/q9Uu8H6A0
aVBLl+4q09fACC5M2veraiDDLH84rGPoMz5imr9w55Lt4ainoQQ+4Moh0Z01
pDZ9k1VxJqIZPYDrxQznrj7XAsxyvTSTOzD01nEFrFeIEYw6haeZOt/u/plS
1HqE+EU0hX+V/P7ZrKGaYem2Qa1XEquhIubGYmU1PHBb8d9yABfrezybQyMr
V6M2xJiZ4dPlNxAJwQpZ5oXOkP2QEFdC80wqulbVimMko2rzZXCnvszGuZgz
Zy7LQikMEM+OKbQXFMSzEV/eUBXlFp4qDetj1CoU8Ozj5AlICTuuoTLR8xtX
pq5zNBhGZWkP1FU4lN3tGCTJDAkTuUuczZyuGGO5fjXqp4zkwjoN7f/JgFVn
ipVS3jfs11W9MKnKGZu0meog4ZfZJdo55PFG+mkKn/HH1cQEthBwvQazyPQW
T9tslzTUT7r4tJAF5wbhJDml0TUI81XhbJTK5DJGyJp3euMm+40fHvGgxpaV
S4lLrr3pjlbOsG4T/Sk4H5Wg5aTSu2avbM9uMouYp7RNa9rBFRn8EBU/Z0GM
tPaYwijmy0gzbUz4zfp1y3VlSi9hINPgfiKUFXvuqTb8/cgMho8k57RDnUHi
GPd8WLWCzzWFbMERqVzG1H5n11fWygK13OB27yVzP6ox3se68hNe7Slv7z5U
hlG/cG6h6StkcZkWvZWgczTQooo10vAHcf2LKsvhH0Jakx/791U02xyFlSo+
sPYRNMZAdHUUyT0sOWHQ0yXRsoKn9Az2ctnPIxMXzvdFHKDzYllSWdaVdTCO
39lSIst5H8Btt5VoCQZuy+TXXjqLzLZ9Zhos489WJdKgswntHbEusc2nvOmH
Ys5ewu/AwHKOlyxPaoY+nIli/b65Awf5A/DGP1VcJTo8o/cnBPJpIE20iVz2
NG5mrQdjUJMdXpvZz4CRT0X4SMK76DrSXrKHFr66OzAfROFCYil8tISFS4lV
wXBEllHF+34sjSXHjX4p0+b3G/TLhm0Ly08yOl6MbAN9MZ+KN1ndtzZKOf0c
nuTVNmpT3OSo44eUxudPDcdhGLnQgYHugDo97FaswniT726J3fQXWRhDp14W
RvSKDbtAEVctmffl29T8FL3d9J4BD9EZ2jChR3kl+w940SHmUJksGTot+xYG
/pBdyMgXCR8Igat7QiY5DIpzADMN6/4Yphn4YRxEn6p1VYzfaxutQN895I9o
ulQpbRIEA6tnjuFG1E42YzCBt0sK405nkXPZ1yeyJGcN9MTQ1nYUu3oHaBTO
KCe7xvFcSVCssJQnXtdMOyC2JUgdrjUtUPUGu0SE4dFov92VcDOoI4SGFA6h
a0ebcsxbc5uBkiR4uqw7bGIV4G0KSh3kPCgnXpmh97fjIAhcNq6qQj51M/ZG
bXvdEF3HxMSlLXrW7zvPGMLceNci9AHylzw/VknXwqvDMzTm/IhALfLS7tor
LlePjas6A2Pq8JUUp6rGJdrgK9ZoPX6GLQBZYEcirWfMhaZ5j+dyTf/EPST6
znuKUCMQmQjgVv/e+IwYuBuEr1ozy6GFqL2xdXTIE720Tgyi5zbbjlv5Juq5
qVzNm+B1qPKVaEffvOVueU+utMN6vqDZDW0bx/Dp8UNvKRclW6mV1BDjRO3J
HPmZ5DvhCsvk8LHITavwSD77utpiF7UcynDYx8iwW5NERn5Drh9USrYIfNwI
2q9Fjn6CgxIBjpvnQzVR8pn90e1cvqIb4iQ30hzdkK/6mSFKCOew5amkEei8
dZPJWQw/qOICvp4Tcs8rz46JiNOr8EisDv1/7OKPaxmpBmr1340qRT1yqNGi
Wiy0eT5veAnnBiBuMe/PJoWVRga1khVdgI7BVllu5543yY112mh3d2t6ibiA
pPGINafGMNUTzGjzSBe357miMeqyWwI6xDrAUA4TsYxHqqtKURNxwMWk5/0L
yItl06bNlmNG/ehWg1pclMg9SmXwi8T4/XBiUs0GC2FheMQqiO9R4uzQf1bY
/aAIMJnpPThZoM7gjztamNOrzod+PK0X+vazeH9J1tGIMyI+j4sDDNix2uha
IbRfkz+WMLZK9aaD2aZincbkhIkQxt9zGXH9yfIF6ZsljLnKdyHRwAFAKI2U
7tOFW/FNoX6XGjYt6Q3NG6R+hDHsiQMcs1b7U3VV4mIjXFXFDgZ5RwwAnMwh
QdHt6Z8G9zfCi99Jx7GVpV01acm3XTkezOJMJbY6Ncc8X+BIWY7mZtMwrGS0
oT4DpB6KvHdNIbtO37Ezr/gU20q2GEptphTz14srbFuQFjR7AFT3MXjx90Rp
MLsuOsl5atG3sMvt+n8bSKZyf4DmAj2A+iW/O/qlWfwk29EWT0m2Sp1ekKL1
uN7LIMf1YVh98XkggCr4AVJjSCvvl3Eh5xuS/bjLIvdHGdt/w7omMqgvx26r
+pwDJlKX18gbcRze/XlYYrh5JRThMSUl+d1kPQDWgLSJrC0AsVBhxB0/gfR3
e7ojkhg4zZCIZVqLOeNjbkFbhSuDxIe9qLmXCxsoc7UPEggv89qaeWZurStI
aPxhG7XFY04vtDBSLRn3G8Y4hRZdCMwbLuICQVPGwwDeZbMvL8MxZJHNDmf8
B/AdFyQAkWco8bXgk7R1k+TB4b93jZnptTsAmgQ7zg0UIeASTnzdI6XNdVrc
J0Kj3B9m4b9EeyIca4pbaS9utMJh/GhGa8N9J5B847od7bA6PWNDEFoszWEK
s9sE23ccOKWrjYrr345Fzqj6j2pF7h0DzkgBZfj3J1L/7K+hro59C3CqPPz+
aSoAcSC5DACf82FrBcJZY3mQ+w1WBr6gQwnIy2Md7jMsV55krLFJP26YkvAW
LcbZL3n2Tg9JPGfS9qEsEpLsljC3m4Q0xBZcPKc5siJJyK47k3qAHuTm77Jf
6o9ZXlnXP7i0fWBeJbPg0APGwSh3apNA4syK5rCmvO6lwZjUWmlDCQika05M
UqwrxGCSAS9CLXRBpanA5iMEQqQtrqHj2YzM+TscN1eEg3sNOerogpSkVIvt
hFs8H4nyqvppVqbXI5RAlE5LuxZxz3/JBqmCSY6kjl9pVZIXpe4VEGD0owBi
Le7Eoqw8UFIGZ93qqhuUQDAY7s4l11Hf6X+bU1N+8eisTk9rheizAv8u0pVt
7cZGp93iKNwmPs/KrJYBE03H2ua+MHT1vVUruhhz3fjnrTfSnQN3r0vWRHUM
26yWRG/tXG6szqsv3rADcK1Qz0dAFf0ui9XM6hOBVXBnEjWE755lk6LZVogt
b1XjmzT7cDgt4y7pu/072YYxq1gyyO7L/5wzH0G6vgGlQ66mIEKDAjxol2VP
cQTpC5LRrIaH7pB7Bp15rTK1fW1CGgGtoKixiLe+fLGLPhIodxi2aN/SQv2B
u3GwpsWM9F7S0DS/8wa68dQx+CaRJGWVXwAATk4D/L9dQOJod0Di3cG6yoMc
YFa3GS+KVKxX8oE14s+FIOaSh9XN9M0A6IjkrxIVqctiFZDSxn1iY1QtM7kp
DSqWRHy9Hw9PxiUazZhnwjRCSJ2Aah0FMf0TX99rKIT41JfYSVrhUh5T0W1g
afhr7UzUK7Y9cKfA82YsBxBiHKl3slixXs65dFHQxLsiDYeDbgkIS8JWfYTh
1239Rq+PFkLinafOWXNeT0TB9tW6Hhyro3n61VSWi70WxZNkBE0aDdZJjsVx
gzrH9QNF+H6M+ffTYIUxdmy9se5PjfFZ260ajvelFfX0DNw4x2B0YA9o6u8d
DztujwNDKbwj8mMR/paGPXKUu4EHmrFXFGZziBMhRvoLqpyC3pCxtnFXGKxf
RlRTp6pKMM2g62vWmhw3J1HU+1R88++g0/9o3KCqZ+HVfq99tHIj9qJmPLIs
T/GI+TvD4zjvgvHkYbMXDg+neOygNYUSO9gZD3jhx/gCao57aBJzalIbJybi
aPIz8IgD0ENj1RB37LTS8WOj1yhEQIZU4g6sXH4gmuC0KOU6ff4D4PAhbDq+
57v2RFODBT7D4UPHEPCABJfKEodC0RYZNteBVyNwCWbM1VCM65hanjFdjvDZ
JJmNZu9zKOmFHQUKhFJ7F5KgnzXYCFMBOMyrFLnH97yJWOv095tJ2q7Lx1xR
jkLBL2wqLw8Tm0Rw7+w6b+U2teekMbk7Ekr2aV5Uno3JCgAOXi9FjqghvfFU
RMbYljPOLgIBainw/GElepPVxEcv0gkkO6HxD7uJVSq5kDkEavxY7A4hK73y
5vT0gGfXuCN2RVVumWIz054mPQUVwvXKeSjXFjhyhjL6Oe1ZGKVztq+lOnGn
ch3OUvuQhf2+myLqnGtw7ZHfXpHKBsEAP+Ba8ORZNTwXYTqHnGuAjwW5WVNn
tWQs//1dOl5qDJu+GypBJUY48f0TM2d3b0V82iOj3JAOVt9X51GMLArxX626
zEfZXkGNcPhP5wMKqLyvsxn3P7ZDlxGXaX+JdbjvTiIYrfb6Y5Ofxw8SDJma
6DN3jdCkafANsakr8lbEc4OC2bUqCWgDshpM+KaLdl5TS1hI8xQ6pKP08cM0
G399eK6ElbQZGlC9NEuDlwZyBB1tdwm7gkV+Umhktmlltkjcu/VLPKb+Q7We
APRLOsXu0ztnB1pSHjum332uwWYlVrdl1/2lNlR1TGnYHHEoVDvB4IKdVVwy
64lxRGj+Qza/fCc8Ow5ejO6gAzQLzr+d12auueNjvN5Y6GsiL7DbXe2OdX/R
sH6WaApAYaz77ZIm7541zBmdDmf29P4Cyq6fMawKh3YUC0PXjBMzrKEZVmSu
s+FpgKQbbc7UGlP1Yivwh1zWmxtio6jozSmNMrQhiaBUZG3BKS5ly7UN1CT7
KxJes40XMDvqVCDL0XveMikAX61vOI8zWRYKrQsxoqXrHMpgaTGVX7oPyeY8
BSkcFoxr27K7cjUH1FsmpynbIjHdkb+UvZ5AI95lKOCCGr5RgWDCXzpOa6/g
EHzf2pGzLrZOXJPBX4CK/YyvbSWHPDYkbt57WvYD0SxAZotX2hy4ybK0g3gY
iPiCidvghU991mtQqFcqNkGFVGui3HhNieybyotLrwQFST/l/tR7X6H1SK9S
BikF+S+jOtXrAL1bgXKy4GbC4ujlIDthdJe02+d2XThIX0gl5nCN2hiiVGmq
8/a0l5YBvvWzMEOb/VertgUiVkT+V6oJdokDMRgD18u0qsDIvIqLW7MnZwb8
phQgZv+2GZlDkH04rUFcdKDBREOB/InU5cGfgT+Ra2StfeRKAIoHu84FbAep
z+JuM09EBmfWh5bB279DWl/U7EQ7ZJ7iabjbpB6BDah5mpAodjAur2wOcWX6
rssePpMtB8yWbk+D4r5nrI99K6Rr/745mkVAql5YzNWKsFQ1usWhRviRCVhf
U22e/eNpNVZMrVhQBE3Sklm3c3o0jKN/Cz0jfs+U8jLQR1sKIb2ym7eEeBGP
725XRngkBCM/Sc10i5DD/bOD2Xi71OuOolvt9vK1lWdpPs8YVcMY0wgVBpjE
omNfmRIenPapQRVXPT1M0Nk6NIXCD/Iz6mxMnpKQ0t0zZDeXrzIe8mWu73+9
PBZr6d+ZhHHPMgzAZzCIVZjv8gz3YdkasmgOfJRc/KTXWhJs/98cKKQvQqCB
enYkcfsOL079n8G6X5+b/SLRYBhaMEtDSf7liuKbj/J5AF2oH+b9V1H1OS4/
s06mL89PgulU2jw1viSDGeV19+F/PKjiV39YcEOnDqXn3j3l/1ia6qrsvtLv
iBCZ3vXfbVApyO57mph1a+Xsp22QrzWId8s/fkcgWxNHwqKHCJ1T2QxPvDdZ
hNPrhuSq00Wd4EEt6+e1P9rtd/syhPXjl2QIZld0xt9AXZPs1pCPR2/jp54s
8DYq7L2oz08ghGZsf5ydp7RVmwzacApJscv//swhEDAosMU2fDlxmW5GZNEO
kYxpxI/CFfern4IvaqDmHA2+QCkSDFl5Z5haO0i8jHrj1TqYAsOIzGGqCHVR
IO11NFJujciWkQUE+a2BaOLDEOxVimfqULSWAXLjEyV/8dYOt6vRzzrBLHb4
MW/pYBgXr0kl0Ccv+4c0egpprMqNN+rp6ba/xoVKGuNXp0KCAHGTTMkGbdHH
XrOeokRq+3Sowi2iZ/RaMSXthJJ9Ds4GdiOOn129SLCR/1iqzErlH6r5k7mg
xUC8NCqqJfdbkidc4OlPtMo6zUNypHeJ4NL8TYKgLbZkx/FyQz+4dtmJwPJV
TGMMHWIYAiOp8oelUa0QHDoK58G5ZJKf/4pIAbbmI4QOyzWSJMGFT+xfpx5i
9Biu5mf4uJdkwxEMlYJ9iqbei70L9DGd/EPHrt/yl2Rc96dP217gOavGSUH/
kSr3O9R6sctNj7KaOzaE2kuOgOqTjlEuIYZe77YNLeeOLL4jkXJ18cZkRgQx
ViUDd+EcEa/IXAwCRYb4/qolL2HpVP+qZUGa82N1NZbFPzAuOTLWYyqiVfQi
ECX2EfejjbFSdGGUSl/upMpnHDSQWQZl9joUjA8fuZY/nLwiZzPXGoE087F1
kqkbmQcFAOENfda2rFPyb/PyfMflxqu9I9KfP95OwbT1G4G5YNVTP+N7MMir
mqJAtFHwbm37nl8BC/HJF7QkIQ6ootANk9DWJRpHhDVbpp8cpusojyFi54cO
JlJLqcEfvZJHvlCkA2bqxWRXbkjCogZhfewZS9B1oUCNDCnnOXDYnt7Yyt55
ro08vQfN4EJo2YjRA105S/owZFBAl4Df17WvPbfMX7q1RuFb02ta3W4F+z4q
qq3A6CUPTlaD7n8PGLVRifU9dQXqDcaS+KqI/UIOSd4yYrpazZWPW8Uf6MDK
BDOWXelLf7gg4i2f13V/RmQ4irh4lg27nL3t6D6EdvQWYzHcAQUcjivrRuYv
wdvITE6HcQXHJriqbavxTpR+Z8pJAzbbrUaMIYa/LD3mJNVjDT+VbkP1uXQb
cjOykIWE26EjvA+5G9zhOIugZ6ljXQW6+GypzJmVlF8/GT/UVe7cLy/m/cac
HRtaXYpd3XdDgkA3/3RwrcoxsGiXh5Q7aJRCv0kTJn0oQXjCETc8E+yWW4jY
NQYUT897M9D6AnUxZ8DTH7WFGNGbPJI5P2p1Hmmpi2iZPQKrHNQER+lQ3nAU
UbEw5xU7vGG3BYGjlwTJw7GVKMH46NAVbpLdZ4F26PLO46l5TQ77O4NLL4+j
t97U9OBams7V2MgShnA0e9nKiRmxOmp1VTCdyU+DLw4bEaOqFeEQdqDDRdeW
9L59vSbwLsPys3kM3n7P02FK5iWcvXYXJei6SMqV57ryB5EHyMAnemVXSCCz
or4GwjRnWvZtQex4WUPplJTuLe9mnp399CD7pAJwk1b9kqmnXuztBiqm+6pn
rv1lMDT3AqJ8IDG4wO7zLI30IkOdkJ6OcoqLfUBL5BDz56x1StHXbsX0l4cx
eQbWENsAMeCshZK3PBML9lUmjg94zPFKBEjw3623Rwj72pwv3fpqTCWkaQuB
e6pkjQjqjpE34iJ3jQ6LtRvCewY/tiYuQ+3mJf+uJqkSfgrOm5bfhvQPEJh8
zkpQGtSDWKXmIAu8uLvjw42BqquO9KDytwy3LZRQRUc7CvwObLNSNkk1zVvT
0sHDWolrOu/IsP80SbBPrSgdGvALcLXUaGz+pvAjKzfB4y5z438Vlscco72C
djv8RbY/a+jCnohY4HhX3QEVAKXUDzHB8rRu0E+3QJ1GwQxoNlb7gPWg732n
qqjFNj+PkgxGR3veulemKdS9jNA9DJYXxRCpeNJhMmoDmUtDi0JpxvQm1dhV
SekhmTOhxgupSx4jRO0MGb9OTXdMlfu9qRkD8r/8oO1QcAy44SKBhYwywSdo
Agn2ABek2ixAugJZkzDeCqz6eWDIa2Rxojpt9Xy6sJ22fgYxr5Gzx4CVPqZZ
M0KGKZu5bIgA6Di5vGSlcxymEBvvXJ0A4c01wYttI1XGnZBlE4r3HVhTdiNQ
FalSAlGVdplDw0BnsAeU8CXlzBUv/8otijYviEAWyVLpKMwKDPAojnGHiUnX
J+qMrD/hTvs2RXq8hlG63oGoF/RQr1yRmPIt9Nqs2YyYXUvqyVANRTAIbI+m
sEWD+Zeu91++4pfGZ2XlL7km4V/crv8+1A7fQ7tVt9ZNz+qfExkgQwZCYI7I
W+vUkYx3qpQz+/ZxVHUxx3DQhjpY6wFqjj+n9G4r+hb05WUqu32uZ9ZzbAhk
6e6FfEB7pU8SsoUCmlm7tPAN3icIFRRnKuP4pdF3u2TQtWqbbBYJ842pPjwq
PTl7Che7IxXCSsKSTqtqXdmQuwoF+WKXsB/B9qf4PTM5IzTblId/VFdVAuby
KOefWz2IfURQcuhM64hNCPvYcsa5i/qd0Dwm1aNWO3tG6HP8Enmr5NFHoBqH
VFEBmryYypuZ76O7f0SOF3B0DJAdARbEwS1zrNYw/wTv+IgZfM6ZkCiJbFal
GYG1bVJiBABs7/GsRoiZez5IT3Hu6CtUGE1UGHiGBfnhlLRm0pYe8pHYCTpc
aXtH7ULtiO+6WJiWqyf/l93fVJ4jFL8S1VfV8dOEfhaygcuP7Jyn4cl/duxD
Qr59XBmYiw83bdKfwsC+YTxiPoP+Jh0rOduAngcJXHo6WddBgDU1zfxsVGzc
zZ+50bXZy/Qg4K+BtEl9pVMzJ9qUPDShS79FsPeB/whmGLT5GYbFBdcA3tHz
FTl+5clUvrhkFo9VtwHf60AdJHgPVjX/L89WDFr6+uNlPuSclzQ4GaWR13eg
tLKLQ34oisBQO2s5DcIVt84C7z0WBcEKWwQVMoE3t3+5MxH3W2acV0hXb/Ad
2Oy0a4Z3VcFH2f7tyVmqG8Auti1u/mfBYB2SneAg6WzNFSwRdJ3EI79urTqE
rB4uvLktNhAS/3lq1sb4p16kUxegwX8idExrfX0hjE6lavTIEJrCDeoTzedS
e0iWzuxU1muD44+tcC9AE/cTu2tMYOxQJbtGYhBIn6ZqgDdpo2wAcxTP9ObF
VuRaBd+XGJEU2grhNRWzrXjA8UgJTYc/k0F0UNcTxbYLQ73oWEMm6/FoDHsX
KCI1Jq1cGW7k64D78vDBlxX2i7zGnIBQDIcvKbNYVYJSXhKnFn9/hjvqZXBt
k9ICrV1nBb3+ZtH2hrr1lc7HDPYcTFbwIgJ0BUfbCYW/+Pg7MjDlLBUs5IMq
TgN4QtEv5eosqpn5aF2eBJ5b1CjiRs/dU2bEDvWoELeBfIwDp+/SyehEIax4
Y95O4HNHPUC7uidVuBBMDc3Z6GqGIIvYCXCW3/mwJb8/nko2v5x9ZwT0ASZz
N7cMipRyEXswdg0h75Bx9ZNsZ/uHGPMt2BkxR/W8KPPYbFyWQteY0/J76XuK
UClZdAt7jnghGb80+ObKqXJaoE25hZCdqO3RMRa8dh/u+WGeJL14ou5S8gIs
Ek9/F3m509CEOcqz7bxanJTLKDqipR9OVX9b3mZcAW827dxSUxaPImAmAciD
oRkQGiIeEJKFqnmPN55mwcuNSb9UoFO2gUCl97Ez6VY/lgJ4DELrl/TjRXUP
QcAdYvx/jtnqI3GJjUblg11XkPWv6p8nhwTcvxVlyxMcw+oVbkI2p2nQ9RGh
ro+DNK012TJ11BVcuNoBlm/dRlX9Guu/fOMthY7zM/dXFfFRHC4XovBzD3/7
ItimU2gFzZUWY2mIrc44ANIkPSEFY8M8o00LD0Bu9XwHf4rS7O4AFwUyFuiw
mdL/FFnzXQgUFIVjRYNDxpdgIPEsTF0CLTbfzBhwQ8gbgqWYLxiK1zJhKeKW
On6hipPTx4NECb4OJWh5XVrPQIOfwOb/NnNB0dlRuFN+eMuuRRjy4feqZ/uD
Zp6u+8NlWak0c/0cE41QIZLQNC4qIMMWX//GwhtUEGReo5INTi7giuoQCScJ
VA20Zk/5fvCKCHJJ4Dd2IXNZc9zHxr/qbX0PbsCzgfI2keFBSS4knRnI1GO/
BH17b5UWbMHcV+1G/UNvCdOkuZdhIZN7ffqOjcXxgZCq7vVqiySgo9PgB0dW
+l6aB/u7+d8CDlC0Ntw4TeGPtp3L2Z3QEFpxhwK0eA198KVdS8JbjveOB2Es
zo1aZw/2lQU6MmyEhrC0obLqbvxEM8UYOsgOCnRZzd6pWfO62jMWS1+MDMT7
8672uwt4m2eweqfN2Fo2m49qeme5fsexKeIEabD1BuoVpE3oHSRa97BiAskL
XjODuqYAqf1T8zVPBXwu0YwgVyQgtN2whmUWj1gIYV0Z7vBcqLPetKaHbL8C
d7hkpud18dUNimVEfpjKonmqALtLFyH8MdFCCXf48VCr3nndz176PdmUpH7W
ocLPD7bN1nhdOvZ1Uexl1vdGk31W/euMgQbmxKNCr6NhkTukaixf08GeXWv/
++2uhMbpEuQJOIduZmez2KxNIotqHUbgMxme0YlCep5zXqawJ6Cp2GXJXdvA
CKPSIv2hBifxFk03x9WUaA4iMsRojhJwnIYW3x+4k908s88Po/ZZLnriC908
B2J/ZvPGr9yClHq9wEDtgTujQeJS8nslaTpTsaJuXTEWbMPQTwBWiXPMAz63
qNlsISmVCMbZs4lk5T5CkJPQsPA8Wr4TDWRXQd8CR8xr1JH3jT/8kAfanX6h
gnFIDz8y2S0VAs5IM+L1+X3GMECJxt2fAbPck9bcETGZ+q0bXVDK4eecLlgm
3Z3NboIMBd27CRN9Zkb1Cq3qB+eHuObxcuw6xyyuZmNAs2/RkZM5DYMgG/a7
ddLGuPoiyvSzdPGDSwlUCAK+Dd9rEpMXBVi8EoWRTledy/UidxMloH8oVg40
wjMhGw41tsJCn8YMVVk00D3Zey26JBx59Ofasqp24C5LKXoomI1Itf5ZZfeg
HI0izX1yfXgTzeL1FgFA6H4yC/nn4hOMRNo9KhA6MJlShWyp+dzX2Yo8D/A5
1VtJmFweBeUauLwbnU70agDQb/nEDcQ7HuB4h/EGEvrdykFupUzu/lESkUgq
OoRrxCB06DppAYvgYQlDwHSHX4+QsC4fz08iCbAFsCqW8OwoCPIHfmjNJTN7
IqqvorWk50/C32YSFTMX+csPDQxIyVV/MkcPl3klWr1HcYlb/4KonHNqZdEv
DSXQYt0kVr4+HHxsuTWBkvZHKvKVsWWayIZoMuyXXsiHqkOKHtcb9Npda37G
vUofaDxgYwspWO65nh46VSUHMEBzj1xerOHf566275TGyTUygqjzxE/UDEAO
oLy74egrkfGnnaIONL/l+OxUfXd6MQmYjTLyLkI+CWUTAV//gfsEJvm+b82+
YEyU1kqDsPSx3zLuvkRqMUV2PRtc6BQL/AjGy6VDk1dRdbC6q93WFBytgBgz
144n7tPmbkn082U4/Qd57M0OKrMowChrruffgWY4JeTaZ2WUbS+uU0m7hCQR
+207RRXh22Fp2y2fhu3eiieMX48ne4FJU8Tbj/ecCeJYrdJHYLtvwf8e3grR
oxvuq+5oKpM5WQ+7ul1JlwiOez+MuK+nLunrZkVN1EE2x/gTR6fmvR1J6YZE
0Zml9Ph621cpfGKGBvVWOs760RMtuHArQgVL2bxvNj271fF2bFQWuHy9p6i7
ifcdUlwxDYqGC2qG4hBNyV+qO7Vx8gfOsrsHZW02thK3QZkUGhJj85MESHz/
ah0tRnE2QVtdgMS6bwhg0wmYWKhjHAFE9AID5sY6gPqa0bJJc4dBxY32YXzv
EgUm9dOLVAK2SqrCyrO+6rDp2qlpAQxyKbPWKA/6ERAgBjDf0F0vviv4NVas
nAC3s+Xfk98R7qTGMo2QAMQozuB1hKg/tBESU8PN7gm8BV6OmyGTpZymqA8+
6I1pJAWKBDPOEx3jj9viDj3ZvZRtZEtZSNgPVTGN8UxuDBgu3M8y7txq8B5R
nEQwgbpejIwN0MHwq+ES7GCKW7YbYAPuLkRrDP8O8dbqdFr5nxy3Os+hUO05
S/4Mjgo6r4tFil/lfCFodfGx08bBiIw8Dy3t9t48HF3KN/XYlBGzbv/pHc4h
grghJO4lS7dxFE85Uu/MOKwPjM2iFZ8YWqvz1zuMNE2EUiCfftAHvrg3Dlsu
9Biij1ow+WUvrbpABzWupI4JW3Hz48Nroc8ZLxh5jIUnduNz0Jb4P7z2oRnH
IE2fg6LDXdUqu+Q/4fc0hIqaO4fnlEKsl6gABLIteekhLjKaTLaKxhv2XP8m
iNaWNgneysycLj2UL/TgHC8IHwV7zr499llrl6yF1OLxteOs8CPzZRjaF/lL
iBtXDi4sHNS/IukTJ56oNc44z2yDtltGjs1QUeBas6grF8xAY14IQkxal/3M
lJHpO7vUHOv3ymGXfgkuxFotklmxRaJgQIalAhBiXw8Dk6cZC9mGradBOZJu
G2kcuj4dKsnCmDG+LHv3O0M2nQ8aFgMdrjwEbBLlinBjjiFJLseHcOOVxaI+
hbo9WN0jUCqFgaoja+J5BSdePuIePw7EFx8UXs2qE0fNQOCVCychKSWJNBOe
oxm/kee2NgIWX9WKTyyCihhQa7DXeVlpv9OgS5r2/yaZrShtsuykLtdhYCvF
+XAbb62mv5d4BsgS1PiozFAQAuhwUuhcu9zrbp96lyAf4Yuas+D5cOXqMI0Q
IbnAma/xm89tI4RSyTKGPm9q1MYnbSgrfoY0UqLn2BV0yxBup3msnvgbPDqI
Ha2hhR3WRCWpQLalGiR9LoyDrbNWx4x3Zj6cFpAaImsSPDtUrQTObtBwqDt0
WnZXB69EOBsS5KKkUYkiZ2hLK3gUlU02w7EqTEcHwIbnJ2Bngr7z26C/Rjyo
2ZjvAcrXMm9fLpYqsZENFlhbeRlrmwKKtg9ISRsGvO/3uWScSD3DlqcBvPuH
O2sNwE64LWwee4RFmrjaJZYV4mNdq+pArtTPeg9m9S8YmV6LimY4MSHWlQF/
4jNYXwVolqxOiTF4Xq5Ryc67MTwVjdMG3pvcSEU7XVGUS5NmfFfUbc6OZHNV
MYLk9UO3ApBLIAc6rsWLO6Gx5/QqnafAxkD/XRAaCV6xig2CvgxtEiJUja2O
XAXN+SXN4ZF0MjQehuSpizM/xqCHhMhHbvT5dmYHdpnSjIRz+sCT8IGWXGGP
1BYuYEx0IbFLIpk960dK2oRFY+A6YbR0sjPxP1063sSU7OmuucHNzKK9BQxo
K4EeMjcugW6KI+b0uZxrbBqd2oZ5RMGrsTe8+c0j33+FfBhjSaUM6qyfWzQ5
xTDvGQKKYJT/Cc6elr2n83zBrTXAV5Hs/l44SIpLy3/XaWfuVAWI3xl4ObYi
o+onTrHYA78PXZdGJeVIm9ttgg6MYUD37edGyA4Z0VcZZ0KgZzvkf7D2juBs
GUvhjY/vVED5cvbEGug71GNg2sLVg6i9LheaZLUL0EpNcLE6+RPQpxqRZpvO
RZAgtpcw7QKRu2ScesvqRY8N+GzMaXXJ6NBHIHHz9eoCu4Cva0mXAuaAvdSW
f+J/s3w0lZngyg2IpV1Y3ZzlVltoEuTPWkwOq2XjrGHF4HobFSZmp2oW9kq8
wCaC6cqFLF8ogHs/UXnr0Wb+2RdeXH2bsAnYsWH3oTH+ijaKnGpgtEHSrHdm
VGPuLh6dIrHyAQQLJaMXlnY8gu/OMZ5JIolaTo41RP+zlKFZMwe1ws3ROft6
yIGdFe+4aQkurIP1fDYq29Jkc+Xt8ey4nMGJyoGQbzYMp2+K4RkJTikDCyJg
BtnuxrDgmXaKdCAdCCDCA2XyWxFhBQPP8kmoJqcss1+03RrT8H1uGOUf5M8b
HATlcskBlzgOpp+bteTXbpDVolqTUliHvb6uKmUJTfGVdZ6HMzJ2s0IkM6KP
tfZkvxK/HTnnn+KYHlT6MJBe4cBN2oM9WyiKFnO2UW9q5nZVySIYdAFErf/m
DeozLS28n5oCk7miMmiveIj8rQlL+y9jnyKMzHc91dsJnfyvHz+hB1Wyh5kQ
rccFp88a7w0zXhHpB6wAsXDof2/C3Edz0TRww4w9Wx9/Clag4GXl+o7H5H0Q
/kFzVzvBy+GaXeQ/nDxS7DH2Sp2FIQqXz74eQV/ZuPrZdmm5IIUQeswRen58
JgckC5K75J0ENYIpS2Jy7CQ0KTQOXCEXg5ErERgs7in73P+2fSQQBhPtPM9c
ulgtHMfUOfHi1trltL1YyhTkS/zjoAQnIj+pLHQye8LK9XdmfQJZQqo0QM0J
VaZw5L1i7yQHlAAt5u9dKaKSqre2UtAj+wd/n1POtug0fGdqjSKB9IhYYeL7
8THrWmw8Fqz/SMM4lLgIVn+mSBgN+RecT5keWck+kSiMOBsZiBX//WXp33Zy
g7F/JNSKPEEMl8AfkzbAb1coEMmpe2JhKAO+oF4mEuE43YWo2gvs7c97LO0M
3N6EKD9lqwH0P4aR0GzRGQ1EKcct0cWfAK33pNPUGSY5GDddUecpwd3nZV+o
ZG2uACLj7RBtHrJwTLsbu0Lwv2enbi+T211KybGaXSAoS9o8Jdgpe8rOzcCK
IUHqTbvXNuBRrOlZfbjPdlseEypeT5iqEbtTFQEyWxB9QupaEh8zMM2IFESk
yYASrMQ4lTu8s0OEsXKU++MTsYkvN/TQ96qcGvtIaEatPJ/uGucaz0ACKEFD
TL/Zt7+9KySHqU//kJX2/wnXVeoQCcFPq9Z+vpzlPF2oFSLsTTRfSlG14oYy
Yamx3EwT5abrdfVdYyxZG6KOZ179/IGgsDMj3HPmW7E4vzQoOCKDkhoZkZf8
pMyrzB6y7x37MBK5muA1GYoyrpm3pB9prqrDxiHvYoqTab8x1eknX4yOgGnC
WQsaQNHRSQjWsg6X1XN0XVHRwFeeHmD8xsHRkL8v0+hJtCSNRjFeZJEPOfAj
Bdq8BrLNEumq4+Xu/+R8cRYt6irkxi43tzJn/LOAEUuVbnKfsaZ43eMXApym
T9OpQQWZhRBejcKDuBUV2edWGbFZcNi5O0GcS4MQyutAmy2VoSvKDZAdMDMK
XBTaAf3ONp6l6yDJiuG8Z1PirmS0pAS+Iz9LUDPkJz3shhqEwEMnWJY4CB3a
BIQrdKm7FYRA6xiSti9gTiQ2SwOzbR4s5t0VOqE9jx/X56wrwRoCSoVJUE5l
Ejd66/AwhlocgDxs1L7Hb7L+BZr2kw1JMgRC5p+G1MUa7e6hFcqIJ8+IEsRM
aXjLGIVQNqBo03RzfKTQrdaD+O/LzPOOwN+DNhUFhiIzb53yE707kaVwyHsh
6G+Vv9Y8vz7v6fw1tYr6+Ob3QBit5dr9A7hbaiW8AFqhncbjTKn9WQe/yCEH
hFWJuHpa107govjtw6bEDfHFsUFUeTGu5F0z/Bnff1hV16IFSX7VP/enap6O
X8jGASYX92XJiEeEfcx+jX9yt+msxWxneCse4AbhWriysXJgWAIQm96aANz5
sDLdu3oPjKCgSmn5Ys80RjFg24jQVIddfiMDyQp31Lk2nWj86yt0J0ZIJux4
e9zm+Kdgnx9Gf+pvNBX5ax8XR+RPOsggigODJIkUZhuWch8aiGRu+kFxMZMF
nKpR30g0FHbFeofvJwuA9A7OhvTF4j7IabLAJm7tprcCBTrYQtSwD5YuJ2Qh
ePbI9vzAaNONQtNf7/qullOLVZYkhncpB+I1UrLmzDNxXnCGQEzhJeSU6vW7
GLnnrlB6zunmxqc5KSk77izsUbIP3XH+lJajnBbMWJcYffj2pQ9/FCSjBmaN
kw92by/ALdg83YW735TEQjeO5tC1KWUrW7AJ9bCysQqhx24j4q9N25/ztkEG
dBW/LQuv+KruIVnlviKW2wMZjJmnF7xkdbLhlz8e2KGePm+Ao7RVcYrN+Xa3
ytbGPsylaNr5lGqsH55MbFZ5k7bfobTLHEYvVN3MoCZEsSdSKxupdfgKdh9D
X5bBRcmWFddfMfoFRnzSDHpWjALWZtztOUqUgU633LOQRvsjEdZYAdg42nIL
D+HDoF6IiSa9Ei+mHWSs7n+UufXzHQRraoxepJkq868eBbRFPCtLoA8+yxfH
ylvl16dy3hKwXPN0wxiB8cS5mlaC7kAQZJz9oRZWKnQfh7UF8rmkCJcXVDGB
oa89gtJPt0N3LtrgR8wahGWbAnr17Wp0d/hVqr1hQLWdaUweXf8m0QKiHjzN
oYZcrUVSd+BGCcupI0GrWmzu2vrAhZv0cBw+YAaK0aLfbzdtjq9AstQgjTqH
oUDncJv8H2ShQscdkQj/43SOztA4kChK1FH0aEY2WPcgnMT3/9G3t5z2Ze4t
Mkb0UptHkycNODHA7WxOE3cENslvxBlB8qbRsBaXV+zvYEtC0u7Q5H9Lk9zA
IWiW/1Hx7tu0MPqpszvvBtl1L2q8v+ydTEaF3yd4U+bD8CleC6tcZ6FIgSSh
1NmzW8fyeZ96AgX6z5/SENwniep6WG1aj6voUsGDGJmPhOOtyC5iv2pakQj3
w/ey8hTXcrSyOTJBNmvBcdzr1V8V+Yta033mkCzv689fFh1scrqy2n5ZuFer
YVQxVV0SKqw29HVlnJxeDWGxx3m2Wz+GB3i777JI5PPb3UNiLECcq5j0ZwWH
zV4VQLr9zLps+usCiCEV4VPmxd/VeKrWwCvtvtjsA4KYJ0193HOJ+beS4rjM
yEi5GSa3z9wQfV4u6DH28PwzNnZ2nheBNmCOglNniLbhqADt+CUy6riOGJZQ
47d0aNUNm+UCFObWNUL2mOifAxJPoOndY2XsvZ+mpt0KwXL4HOIdFzZk5Cez
r1aA44PLhtRaBhXzkZOLvjdLwMscmyQ6FhBzBq3eZMbWq5BEKyGzbzQwaHb3
SEepuTw8yfVh1yaRMVNXluECIk6DJ4BZRQtQUoFC+/tkhtiTVTS4AZ9obS9k
p2zfrpqoNnceMweg1K/zR6mjpguxzzZbjAfEsBTQgDk5Tq1c+JGHkaUyUUnJ
ivG/9lKuGdtpS67ce3j6v5nP0wO3Jk3dcL0B0Rgo8v4qmnYZB/vVCu4y8FbL
zcOLNRXP+hWqm8oqP1Z3iNCmFwv3EnfJolZwOtlMOixMT/DeWqsRCcfXl+mR
hqNcO0pcQ1L+yBisxiJHfybj9hAKeq4jsD1z7Wg93lFDy2lXrofpMnoeCumE
rFAF5oQnb7vHOnW3j8HAA+bcC/i4jNGM7TNIEMSXDcjMJhHT5iOj5mcHGGSm
LPV1LMJDgYCGmgegg2lBGvZluUnIKyCR41kLNhwCQHgz1K1dNJS3m9RDG/tN
spYxTigDAJAhCTxOO4pwOIVd6K54ihMs1rtyRzyA28+LlAOsnlAbjHoBm18h
DFrabYb6ZG6kROuTPVQlmAtI8GAW4J8sWS2MLjY/kHH6FUKkECSznm/yJg99
kiw6C271vNAIBCrkcF3bWb0alNsjW1QGSKzvhibCGagHs/RGWeoep2gKjOlI
L/Vu+I6vVxpDw/+ldtyRuExk+ADjvQQCJzwPyOldZLa+j1mzkh6OvNPwvIDo
EVC5++foUZM4tiCq19aRuDn4xYMur8oA1qZpZXdSZCvc1Gi1I6iL8i+26yZd
wvACZXCQiZU4r1RblYtjHqHbwtccKEnumCt0TdQ7857wd2kbCvC2KjFIsgS3
j+CRXWgzP0Dp4iLCzwkFyp3vG8fu49Q6jAkppEPZcIr2T0/27kcV/QPw9zpp
s80HHJQDmSGZ+nGLB/GR8ab9vtExSUKatmgChmuA0gD43UJTbBDGzVT8yJEi
S9U3QfDp2wonTYW0O6BO04pMPEItVqJYPVOFQT/YMUXlf2zv3j1xiiWO0l3K
ATtsKcJWkUg6pPLgvbJIU4/a6v67lWnVfwoujUHoDMkdmKaUc/UoPBFRb2op
DA7w5B6qT3foIbuTHDjkeWPR8gyq4zTyu/jvKn7j8KXaJVGmbpuqghuK1WOu
C05VqoICIkp7a4fgrU88NrZtFTTvj0IsNFlVKGoOdJJkmQ5nEbxebLzV3KyF
bycKoXRAqCoNKaUV0+I0abxUhdcdXh2emFdZ7KoIYyglmqruieUnqWpPMMmw
wy/QrN8qpAj43f+v0EmTi7u+sghiSrdVGHKKrmw2d52juKAdiJibnuK+pMMv
fY/Ua1ujJ7wRiPGLwsyFE/bj13aD5QQhd5XYAUuQEvbziqUb3ExrMynZ5rj7
qZ+AuU0W1UQHdtgHr4sH3aWrIXGG6uR9P3i64Ay9+oX6A2hW7XGweBxmS6ev
20qkColIHl0aDzZFp7e2JFCn7eVsdo9JMxQgT/8ivXShsJ8pcB5zjyf+NaFh
sBxbG9hwfyLs8O+LSDAQh+7x3Hujc16g3bgYo1imGQA3txGZWRveN/rX7RNx
7kiYTNjnDsBCfH1x006gTQwIRrp5VamtyE6E4Vc/7iOrTXCps7Zs2wDxaqQN
55woPaNU+IYJ8voSWmoViKmdXlDh/yzJd5r/uIJhtYRTL1Rtpt61vdnnmEW1
MugwBq2Fpc+jTY7N1ILMExHW+iu8/NCbanozW8edw68ZZEoL8YOgY0v0RAti
BnMAjF+Y3Di/Wf7RWq6GxY9BoCwJ0vvQ1QGZhGwKNEpXpAr6MlsZowC36iXy
VBoyJZsZQCl/bUxus8nqS7CsC1WU8TaW2+GbkH9xbLGJPwG625Owvhcwsv4L
vRt/WI9L29l1hrh+Ck1ss8To25J8BaaxDQCEh+/wTiFZCmVoK/FQj8IzwYNN
y334RD/lAH08tx9l7ZuSmfmdjvXmGp1yWAravqqFmG37lRMefjttjf7gUmjW
ZLzI5qMSVKs9/yWPm3GOGa2Y/Httwmd22Q1N8fRLEAIlq06eRMPD10M+DNmM
iN0wNxY7TkY4Qu3qCoFnmagFOXvDkBuEYCpO9cHrq85ax8Ao8Hyh/rbxcAU4
QME5HGbS41hF9ah0cBc3qjGcOGV47WiF/BlmgEQ6qM0ZPA6uTzLlzYu5898X
gUQrjfADO4UjMaAztxGsU0nt44AbNZP0jBaRRt1aze4jNwz/BAaZL0QpQu6m
PdO6HhWheIaO+hy6/l8+1SOrHu03gaadWbJ1dyJUL3LPshm6QTLimCvKTnHS
eObE9EihPx2pR7EU9PoSaNH3uF++DuQ67CRw4Jg1+Wm5o002mMvAsqUnuYnc
5JRv8ewwqnKMj4a7+lAuk9L3lURLN6DaaQ+4VcLAWK7XT+MIWT+2OAOhrbJ4
QbHgOvKbHcSnQTa2jZIbkuzCXExMorAB/y7MfEc7cDgzuzS1tASawR1LGp24
bFDxYnxbIPJsbaIIlqK0KjuVpiNKs5HfEVFNv+KOm8P2MMn+/IWEZZTh8uce
OGGzflYHpDPlxHQ3MS45Qv/LlX1xbc6ZsFK/5L3i3ikiKqOCOA4dJWEP60tl
MKnLHiiJWZFeHy8Ey9h7ABF2QyQmDN3vWz230PA7ncKnoL3zFYiKns89nhUO
xy+v5EcHX/6pc5b+nmvi5Z6OQ+ia22AVLqOlkhnDV8E6EDNb/MHvLcVVj+d8
l3Bd6xxLsh92HIrpaCGKv4HQIs1KH2YkwTDFfMlCTnKmTS1j5GK6W/tgEb2n
7LYQFy+SiYAVLvdrNc0W673EXr8h/ux2vcgFgVs3KAuNkKVhnXwquh8RRCym
enV0QVNdNKjzQzbBGE67+YKvjKPM0Yk+30gtujqfDB+bDuKZQG8sTJOE727/
tJ2U3WYBiJlMMJEH7r9UVByarUOnqKb1lKnPROxVBZVKgrIWf8xPIATlLUj2
dLZ9T9Gzz+W4VDwZuFhAyUCtntCLmjGxZ/gEvqEnbIQZut6ZFQYgJeFHH3Pb
I7dyI8EHhfHEQ00RTDvb7j8B8zWgWBraNp0o1NvhPv0uHfbwpSEkIPh2fK5t
jDhKJb4dVutQ3YR4M9RutcJhss1xTqaFLZ0Z7HQ/UF47S0gMePPHXlpc8iE0
FD7sHDqU8Wzm5YvVkeHNYVXGiyow4YiQc1hfGpFCWdIkfmWT/FKWli2V1Uh0
viKoK/DgnrVLqTKGpHluEImlnJ6OXj7Jni5S2L6KsKEOMB73JciLY12qIPXo
F3B994FowKi38PsA4QMJq79tfqDz8JODC0uV27LvCdPtwOYBhrO6Ybhf3sgC
CndDUXC5pPdIku9XuLPLkyorPgF6ZM1iUEX95Np+lF+DgbXX5tKEnxDh2MMe
LUiYPwVlDgQuK6/Jix16zPlW1fXb8DjLTFosP4jaIe1Tha+pP7rcJR68FPYC
xgGdx9u7xydYRnnS1FMc5iY71/S76NfvAHaKZ7vS3h00dQR6v/WXNy7fw+PR
ys3rh7jE95eMa3G1epzwb97wyiUcc7n7BCFhEDMxtXqedMXCNEZsgHnm4Yhn
QnoMtntylrYQlvwkEn5P2N2AvylLFiEJqbid8PE83qnsIYoJMDVaSVInjn3K
6g2nevEVzhoBaPNx/4pv90SR8BzMgfPu4C88FGKQhP+QXpISoXFfmIuWfs32
dSX9T9/BH57VVFLLN+6gX2pyNbewKa8CovyfnOBW9nSI2KSPpMi4I+m8rWCP
44A4Kdly7n2AUVGT61ipKM2AlnXUCbkdECY3RcH9+0vXOXxgbn2YKjkjZ+Az
zBTVrkhO6n4G7v0Ok+tV/TgYzyGtGa5yOxgHaIur6n4UHh7FTXbgn9eZcRHu
5wvrPgknNMQ/Zv0KaYnD9XnmZssgCba3KoEmrS6iwusFwEAn0mI+glpYnZVP
KYagfNqb5bohBdTSJHgBhR+Tx65nY2yIticyURevU+LmD9phKIjygYyFJifN
rkerWU+br3TAKaOw657Sqk1UeELBHaytP7TjhaqS2MWU8UAV3FO7nlUkfRZ7
g8Jx7N3s090Z9Ulkbu3mcrp/no+dCjVYqJUCIKWvZhg57exRQ7jhwGfY/sOB
k49/fGKtaGWuigbFZk/dqGXZ2iFxs2+fV/hoghOPuTQJcdSwCL7XitfPjS8N
wm0eEDyp2M0wImi5nxlYn7cljnUpB1PG2YGy0qvsXkh5NL3nmdxrxiAfDz/Q
DoHg+d0j9MrRv953Qx90ZUCbQEvQNRl9jbO+Cla4RPnDfnUoRWa6cDtu5C3a
3CIwDvF9iSazG7rGXbXK6Iw/J4++jmtSV7YqHrLPir/jJebK1rffn4IZEj8P
YqiofXB1QIJNKHU7MwbXsDIWSPnbk4QteUGFvcpHXf5pkJih3rqXAHS1WUOJ
izdZ1xlGoqfwmFweG84LSqUlENVW6yU5DI6NtOQVFtT5kWdpeooM/G+eNn8Y
HVmmzkIIOtv9KnTuqnr/nOL/dFq6FE38ruPqAtwvBpd7XLzFs/4usgru0/Mf
376zMD4CJVM2KxIHgC54mcpk5GuqVeuRjkySDSztmJ/y39yW8dxIfw3q8kxT
IiNsztd4PP723bgiYzZCcW9L1G2U1zn+8+745oah2Q0E6CZSI14eJc6UVP75
LxTYroaNInE9WytK1ojgjikFYo3SB/EMxcYncx+Z/0H965hSEnGGlN67iBXe
LlM+t4AVy0YL6x1yC/G0+XoQGbl5PRBUTuwExCtheRFBlOgq5KOH1Q9WTVHi
FIUoXiZOskcw0NhjA+LPtoN3I1JpxAGBKSE6V3O92HAsc9Ggw3UmGR/xHI1B
Ss1B8HvKC7FoAmowRXAKBiLsRuh2/r9KpqbygCN+X80RuBAxeyPF0SqouJ6E
Zt0Q+4fhPhg3AEguqFhF+Pbgp8uLYNwGvg/93g3/PWXmHskkASYH6JeiLcfL
k5cDsnkN1sWvFlqc8Q86c4RSnt1dNoPSfXsNp2oliC3NJEypPK2HW2da+r8/
HCJVW+mD7eZh8OTvPUJBh7295i6DJ5BIVUdyErIuxnEIpmb3ME8rOIcbowzu
zbCfU0WgB4m7i5T/V1oazmBSriX8+drTIhTnTCjk9W3QAJgsg/EUBB00Xwzu
ApW/9U7+DXOsBO2sBDM1yKTIkkOWvS7P9b/KzG7UQ4Vu6pdPm7MFolBeOkM0
okMbPQeroAWNWIHu7pRdd05yi9uVPE1C1S6xC4jYtUkAHuwuR/ycztImOzq+
8ol3gwhSMio7UVzX2uDEmXc49AaLJLks25eFGXeGfXFEuCYzbcCA7EjDNCKP
zLKIvJuOH0JJ0qoCxw4vAn3xHyA5xt4VNKbDh6GbmpOwRsCBmGVjnI25G6BR
PrqIM6VvEQpsXXAJr4kPmkkTDxS5PvB/cWziBdleZ/Qlmg/+PXas56Ab7O5c
/1WxFwK3RHc+ctkojLXIg28s99BWxOm2o+cB3oncAeVgSXbwkYRDQQ1UKr6k
OMrA2yuyf2TOnAA7xO3go2F/H1hB1W0v46iTbH3OOJLIHbqVtvn4laOEV0/2
CD/pafh53Y9cVM0YUWnhCckt+JKCiyvWkx34kPh8tYQNvatEuxzFYD5PIU4Y
psYI4XtUsv6MJRT9j25eSUwWWyh6NRu2KTPSILjKRYvuL7B2Xuy6NTvf9z2+
3g2pqNE/CANVDmjiMensnbWIFL4olRqlphPY3gtLPEpUlS3KgD/dqyU9RIm+
/MrK2NYQ0y8fsbjVlEAkMEDdmeZk07UY3nyrLx5UI+aulbRpzQLkrdZbkzdT
/0IVywZk8GpSuzRjJzISPu07FoseqqP36eTti0rq0a1jEYnncxPoZ5rFKCua
HQpFnY21Z+KFJQMOwgbICZuOMEKLUhUNnwvDCdU7+wSPURto28UI0jBccdTO
1gfSXFprM70wQx6VWfF2Yk2VTejpDFSYbutSCCwBnxTn1khXL/QBhOtwMIcI
Apx54HG1W6ONd04HMQKGoCogx7GPH6faInyJDGdqQYiy7akvDqgSIe/Dd6Cw
x1pX14Zw8Bh5tgf7voHB0sQKZKDLpCKUuDFkvEozGZWiActKOsOQ50Qx33zk
7EUax6T6e4q2pftWZL893okkFQ+OAkgX2/KzieIWCez+DeAKJRiAwI4ISJj1
CexDbcuTaDMaJhqgVa5n3tdHU5AzDM6qkGsDTSkv3VJaeCe7C07CPy+/pDvi
salEd8adV4fQTm7NqQH76WI8klZb0KXbj5C2MDR/0BKAXdu2cNS8ZBecTn8V
bmNO/M7VomOv72rcDpixuoxgaIZGpaDj6Siun7YB2siq2X7A1H08CGqCb0DY
xRWH2lmn3LWR6iN8YFLkPkBU+i5/Mw6bCEL1OSZbeawitrinfXSmIXJYtNga
4XDnmXDqI1yzZqTai/rjxqFpbyEBzvUS6xWIyMOjo20RjxRXdvQyVR3isbBM
CbGDJTxuRgEsYVCwkwtWEqlHgXFuao+0hwlW1csNPBbIddNUFvgsv4jzUSi2
JlEG4L3GSnSPyW9eP0vrm8VoF07Pgobti83JPMoxPb0YhchKBffUH3vnSwv2
+6HQ5H93mvcgMfHC1AeO0nWXvc7vqg8e/m4tTEP+zz2ZgbSXieG8r+IsXFo9
/bbbuRUIZjXEwElT7g6/AqpIFVwEaSemtuXT1qRRmhV0NNrzkCWmeRjbb8ZD
77zQMI4U48gAZMZYztRw84yKuKp9A7VBpy/WwSIDnJgLhQc7AKUkVUyrIdjG
rsSzFVyTWg6NeUaPdfGGyo86WgziuII8am6sSgbQBtohtu/LciGDUaJF5vrk
q4FAWbfUeMaCTdeYesLYlUk5WJpWlzpSaK3PbZedQFdMrrkH6QriqJl/kamc
cmztI/Ez85X+XLjHW56X054D8il+1a4bk5lqeZlcC/QI1Vi3xP4F5X77vTVy
YCZw1rry6rDLM7iHnr88DayhZTItJvtBOIxFxAhxQM03Z2xX36KXhW6/VILR
d8FFUh6Gn5B5aJvJvjbufGlcdP9KId7A4ZULqnhR9zo2oniUs5US+YUFKJsO
hEgYDyvVg6Rv5g3h1qphl1PpP1kL+4A3RIkUyjTeNDrgfVczdsExxsQSX0rl
Gyrhs7vVur4IIqQP58aQf87hKyz7tsoPPU3Zokr5iTWbNq606bhU9PKuwZ9m
NxHOZMEFDxZcfvRUGVh2qsBnQb2UdsimHNgEQyKE0wz4oJ7D0QV9pJ1grhmZ
W5qLb8gKVw+ElwIw6IIDvkqaI3chqmO0f5RVOgxHZD14V0V2d6AOqWpeRoen
ynjz7DO0WSoxfVaGN6J8lCqadMBmIlCj3l5nHNA6KusQvM02QG5eZgqaSXwA
IaNUXzVDzSO+9W4UPNPxmpo4JJ+3b/wTPhowhdLjb3Bh7vQ/mS8k2510On3v
UrjeqR27+Ik29WDAKdFy1uL//NvAOSRvN8hygaYQDlYwYIOwPuf3RJrvBTUC
n21iEQkEeMPmNHuo7kvMObSQ3kus6qquU2bw9DaD/oxMcDyHh5dnjF+NV2dS
p5/Jr/Y0Wb0HH0qoMHu8Pg7RjZe10QpDHlLFvfcXX8r6ShbDN5V210NeHDwi
Ch71X8QRvSovH1Xdyd4Q4rbEjCnX7Ro6Qy3GXzGiL5o7DM9JDMn/c1l7ghOw
/SMZpI3ICX1LC3+BgXLc6HXCSTHcEMvc2nKzuU+msua6cqlynhrRmZXaORsy
OOwBq5r3Da3mgJLR0ytkwzmjnPsEuIP3/GqfcSkaZHLOHTAKrfAdoBATL8cv
oKEZUGcwHSU7Ul+BbZX0kRSnnFRIkA08+gudUKv79890ZXzdQSTSsj1l4TP7
zVE9O4C7Sbs6rBqJc0n92oLHoYL4rv5P3yuHC/rn8u47qGLj0r+YOczT5TmP
ONuphoVxE7wBYBqi//P4aIFN40fRAf5ZPt17g/fOVTeSPVxI6aoZpJtA9e6e
pMCLKzaEtSPp7kAdZtNLEpb3XECRuHRE/3G/FvX4woe9Hb/s9Bz3navpngcw
xIX2A5kCsU0jZYbWbWAs7sEpsg54IVUzPWnzy7AkhitJW/3RJJ5h0R8KPj++
ZGPUqnifWv4/s3ryXjL6t9I71P7g7FWK37jkRF0dHpsvRb5Al/Hj4P8zqvIE
iGmcX19/LHc51c1zcBYUU7m7eKwywbZjwy1RVphskWu8uBD42EaDwd+LQ1uQ
BJNJnWiGyAZ031yMaltnw6dG7bPlk4OUjhgRoNJDf3M/9h0Y/DoWB9TKlKly
bEos0R4pW68MaFWWJfxKeWKqVXjzxEpXUMY+CrUx3PFrPgw2aD6/aCTWkX8Y
BxpaasSQJ4Jn5Id8WpB6PDB4kpnQCiPanxzqI9BTMJhSAcPRwh8KkMQz9765
n0yQU7G2C7+X4DhKom7nUs3pji9XXwfeLXAu1IWK+YQxI7ZxjvxQQMMgIW88
YA7Ab+BOZQOw0Ot+O1956fbeySqLtMNHL0OnN9yMRXjIYl4Sk2BQW/d2NfJ/
/l53s8LYR4MdntSNEfka0FeMudAWD6Mux/XCdjosFsznrEUgDnVbxm0QjOwm
pif8s3N8L/W5KvYc1lBEzElUOiJNpdk+8J3zMYqE0vo2xkKhrP6SnZfwdswy
+MpuEQOipRSNtye1YTlRzpMfiXsB5XXyZ739zR31+fRX1+cYTVz8dN3QXA4L
/+wlpVqXq7MzaTjntABqpTfxlRNBBk5+tPj5wL1T9jtUSBY054ohR++wdDzw
By9hb78zYnN4QV8ESPyYokqXog/7batjSlHKyOKkUrVVGiOvC8p4x+xAZ1pB
SwiDV79G6/Yd9GnLPylKVF8mnqNccPyUA+7uqL9jOmhjhNhsrEWlQkTe2Vo3
00zKwkJiYmePtl0Yzibdcrdu8012BtLE31PNydoC51NhbfF4VswVAb/WP4lm
flnPpmNvvp8AJN+0CdxxAq9aTB23g5H4XoCOkhy1RObONiEUvkErV4faPlOP
8EtV4WHuY+8oJ6IoVSSdmtX+Qjsf5feVMSXfcOAlXfWM28Atc2nNpE+X6wNA
aEmHm+ldJXinabtsGQfCU83IYH7gv+CfAEZDqNx4ekMh6QRR+w3+9OwsOwLg
+rIjpwRlYmlnPhiDuCSFxb2r3dDM3TRHvplh091w9VUZMOE4s6NDgzZA+vqV
MIF7Xp3u5MshOmj+FM8Li4yLCZzkfR/Syw8JFAaC448HJxmG4LnNpyJcbniZ
bqUJ68kUxhJl/KbqwhYfCV5oIbgoiEq02Zjvojrz+meGPqm+0icK31Tzh4ob
kYZN0dp9aeLr3gMX+E4qBbnYaNg8y/LRivDkT+9hdD0t/BcOzbHjMXmIBN7m
2Xn1wd901HAiZbFs75apTUs6M7bTCJCpFWfWwVHPuTCv7FWyuYzcqP0Dn54P
eHRqhVhUyKz9r4ruT3aRWVbwVGI1U5JChjUmtuVWdebsEEvE9YX2SQrTKw4j
oD0wChkWjuSuPUDiCSWASGujGcfLrp0eyjuJ10dLrIFo5PEVlEY1Sa6uLGo3
iQAKTHQ+Ljbi+Sm5w62DkZw0vIAwuFj7La41bMkGBwiUo0XB+GhfhQKMG5A1
MRYLa5Ji+88UK7LYmC65Rdlz12WT6XcV4TAFVRgeJWTEpkjjeQJVyBGkqops
tVWH3fjuRokTUmIx3Sq0s/QiYoRGz5/TM3XMerARSIIbr3EghvYwQ5sWQk2s
G/LVSgf6XuSW8Z5KkiyLUy4baXG8DjTP8gALuqfb9BGOfJL9utwK+eoNU3kF
VeIJEV3BMNYZvjP16LGGKHMh6wtHnIXFvztCUCVmdwehsGtAN3sO83+TY/W3
bg24HPMWSvjhIn2vlmzt46N/xPW+Kkjx33uomRLhV3B2j1hQCWlzCIBJIQQm
q79ojvTifH8wIfM5mr7uJUNgqwGoAFiGt7nor/DOOwsuqXeNoDKgfcb9bB/o
luhamzM0zkKQh8uPp6d42clZJZKGsM52EhWnp2B837LjxPaSVnWBqfH1yNOt
wsZ7jytOYkBk7yWcWRcD5/Qb66Xwn+UGbUVY3G0SEF3VpmebAGLlH9JKQH+1
cMtBgDJJpO2TBY3Filf8WZasFdt0fc9ZXLCImYA90jKt7LlAR0a1QxqIqjtO
DzxhM0K86J/HGi3HV4AD+u9FXTcAy85Ntd9bJ3bdmpYjK3lsWwkHAPjdKQNP
TMU2R6UM05l3ws3lbRyxbU/y40i5mI0cKfORiqeaj42W+EXatRpDRZ4Js4Ke
V+hhOsfuiIxou/mRXow+pKmOR843K8CvlAAVshFtF1SCW1xNVKHqB+1SpwSi
Q6XPQJbz3S0mqiO1p4jHuHLG812m0q9EouJKFntgysf38x4utlQnW3W/qJ3J
OWVjofKlSFxzBj422BdWEe/0Y+NiXDTgsb5iqtyG95iS9H4ZjQ0hIDMsP1RB
KotdcVxe9Xm9rY9rbvJtKirRmadF4UCZkAoHA4hu6cqKanfneUwkgZG/Ri/f
xG9F3Vjx8KfoBLcpDZ/pfXFnvlRjgkLB9nIo5damKgrKAM96HArQGveYDbCX
N2nn5O6J4LmoUhKHHtApXJDLnCm8DmJs872nygCoiFfboNbjm3TxDfHmHs+H
ziHI1cZhysInXjnGVlK2XZPZwPulKzgWUFOZx1r6Nr0e/MaZOfDKPVDvf+Jn
TV1Z6U6ERd7F5Ezue6A68Zfyn0DoVKj1XBjeqEm6W7epISTuJmhyp/Sgqcpt
KVTkH7Fp+dHPTc5nwo9onbmXerwAPua1x2nd8dyFb0SmG2W9c2Dq7GG+UPvR
BsMmG8Ji1KwL1+/Dherknl0HGG01L6OLL+/+Cd65i+l9VS/acX+oVRhEdejr
KQpcDFcQRpOJOqCXK+rdHQWgr7G1PiMg+S7Zm6eZw5Ud8lsewsEDKqn7C8Mf
AUzXw545zLMu0BUc2eWM7zn8daxEKs7wv4p1Adw+YaHRzzw6yplGaXf6K/Ob
hXROTSzSWceA3Ap9Lne/bDOT7icnKQzg4vR0jiU7k7FM9EFY2fxSwbyAnYnC
N0CQdKkoM+TM20rM/GGylRAscYF62IQ+YTdE4fYqSJUXJQE68fF0e5pipR8I
0eCbcvTh6s5Bd43/BnU9ofnqhKFtJHYDvhRB26Njvq+SeGiHkav3/ePWQeuO
uPOLVO6JbTEBVDFsofZMxMjL0FmMWaPwt7hU4BROsdlTAMqwr2WElaRtZyoI
UaZzxDV+XY/RM+Zmcuy/eEICgCp7Tg9oc9oemUoqRuhQ4/NCvAf/gCg8zeyY
dnnxQ3wM71S8sP8ce0MHHrymBKjMsT32FG/2K65Q4jJFcWJ8XrVObIiNr/qy
qWj1JhBF0aobGREdTi3sPty/HFI0a/3NWZbaCzib7AqUbvH+lTIy/A8FS0Zm
zMqni85WyPlz19l5rpQk89FY2f6sGRZSmo9w50AUncwHEFcm0ME+9uDJ96AA
zi4R8JZsdHr+PeRs3439bfaU847dg5em5p6WRHiSMyzAEYSSZxh8+EPelU62
DyQKwLx+2oGbRQrEPHShJ0H8ICDPDsCwK9sR+U1JA6cWOMOu9r334m+t9su6
2XCcCBBuFYQ1b5cGUa+jcj7XFJG+z2do5YQJW2xV1GRChzkYXsJ4I+obAXmo
hCo2XMjTNfUg0KQnE46SR7/qciP1LyVN4ToxhmxeD2QCMR6rkjIN+bLuiUHH
st7pth2NolulFzu1/BP441XxRGjw8n2+6icXPFS8QJykSJnw5/WGGKp8CJR+
/rzDBo81ajH+zQNyHPDPoocmmn2p8NSiqRp6JYNuXEfWEgocv/AVwiIW5lLe
PShTVjwP8M354QPXLrGLGI4JNFlDHsLVKCixmTsGhA2LOhKXuVpQSgEYYLY/
GoSVPuH24o6ewNu6VyRgRKLwSlf7elOFIiJctd9lkMDgAYr3SigK5l8VQ4vD
4NI7mY5NpULBiyAz4YdqyutrZ3rWM0TYWi8Dr2912T8UR9qEfCLPiZkMp4ST
PJmk9c6dOHZ2Pn/on/1erZ0QSZdE04XfSrkLLl5p+0ggrn3WDmu8qqIIkv2K
oQXNxTvY9UVo6UNkmZ/c+H0Y+ZaWLeizSgnouoYLx02Dgli10dlM7hiNP9j+
am1BHcJ6/x6wzaBNSjX842m6LawePPR3K2buPtUSefg3cueURqwwb9b6ai1P
Mjky4JK8r37EV3fkAbs6qXPsNY3uvPY6ZFsQKtAS28m/O57FFI/Nly8UScYy
RwNhgVm4FrOXYq34ieR5PMwC/jea1gcj5/BjWa4dqYTmphGYAcdlWy0vAmu3
U9DqA/SrCjKZkvLQsNHf21snjxNH+OQ/nBlhBY1O7eUNa8H+V7RQthw0NUyF
oQAhtA1XDht/Nx7/g34E/PxDoIDqPmMmuE01e+LjuFnGJAx5CTUQfsIpg+Cv
jLsDV7bKpDJkzx9LMapiRgYvUfHUekLF7WD3RJzE6s1ZfvaIZvrlyJjC7r4u
o0DZVJYdsO+mKgsBKqoXSQnkgLEDsS5B8uMPkoxj5VQcEezB7ruXAKQVqmRc
xkBUU/JWoawZL6Ipa4lzfUQzFLIUHP1F0t4aV23AHqTN1OUflk8Qa9ifAX83
JrZXzI1k/DiIIk1uIxFKf16BXSNtyvZGTAhDGGHHrdBPdcrvwQA+zeO+miO5
KyXEe1fBp5F7EBwa4F+S+eKA4oCSAfygeycO2PG1dVxWrd88oOz6valrJDIG
PdOLy54UWN/415AhvVgf45AAIst62Yg0YNxh9uBk+0cD3xiqHbwqIl/tDGAm
nVtcU82X8efufnersSFHTuZ8bUY2Fe4Byg4U/mwAy6t84CY6qBeVyD56T2cN
nWKTl6ImmZI7/vTJIpyMtnA6h/bD1P+xGP1WQol9ecguqDr7ynJdPM9kt8M5
1Mwm+rGDxQjrXKyPJB1Xl4b9KPhE7qhr6B4OU5voNCC9jnlpqt3L7t5k8KpU
I8PNkp8N+QV2HHXg6LQ=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+Ep2A3R0s3ZFkxCfsy9ZBtxDMa/WpFQE5y+ID5SRUsR8+LqylybyYewpbt82bUO890Z/Mtda+Bt/PZQHpHUAoGVW9tR17NJvZ+e8Rj/JjW+9PDePwtcEWYWBKYLk/9tNp0dlCiZyGx4bwnYPLVTr6asXWcyisbSwWYbt5cUrQrnyrgEb/omALMm9lNj21pibe5pEmuu4QR463+UCR7ulL0q9VwUEYbBXiCObKPFje9Naw6MFOV7SaaNr0RIlT57lfPbf5SwvNWcMQXk+raEuM34GoaztdJ3ClShMxd2LYsJphgmDjJbUADDUadBBFhxVobg7zoI5ubCgFPk4qmeGo8Aeg+e6WesvUCFNbux9SjarHibpLnEGWdT9nLLCM6FNM2ow6n2Dp531GbS8evV9mzyE7bmryVf++4Pl9XwdKJtp+ZQ2uodwzMWp3xABNCo+9YBG5WJlHKzKA+2se5MorU6GPPYcGTWb9l59bSmnXsTNfAz7SmAgao1VclU4fu6ABAwQiK20ZPCYyetpT5XCfdF1FmD0nj9R+FXi43sVua7VA9MxR87KhBCLbZfNBrfSqUJhfoeyorn7RSEMWVDgGRW4jY7OX2nfvifpvRLh0PJYCTtxBuew3DHlh+fJYjGyN6E3h9K0GrABj3Psyv//hhAT6URRSI+hN0xOsik/OCANrGETHCJbmy9sgbvRkayM9pLRUcwnmfmRbZqjyYg2nq47AJ8eSqqOpFRu8gcNHxL07iztb3EL21vI1hJArV1ztPA86m5REJBRw4FfH3lx4cDH"
`endif