// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OYE3CeoHwNYtBwLTW63BKl1i9AiHNksAwFiY2Vu1Wv7ZF2wVdoNG2swtJ63Y
dDACvMz1qPpF0wIMQO7AdmdmpEvVtXkXQkXQ1a/Tmruypkc7ntMrf0fib1iJ
JYvKBxKO2GMGi+w9DLl62Z70Kn4XrEhNieKa2Ca3PuM/S3Kxb75oTC1wJPJi
tkt4QCwDUpkfFdRKQpgSrd84I1E12e/yRGcPEASZp/lM5r9bdNDG39S72kS6
F/KkLPAGuLL9afnCU63YVBbJzbmd8r/DwDqo9LPTm/nI3bc/irgtn5OW+fS7
gQ7es5dDMHxW2ttzvt+QgBXL2EVAXQ652bmR4fWRNQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Mt0SKgnZQRBEj7c1PiL6SxKI8vfU7617K6mLHWXZyRAkGeoqavFolseNL7oj
Bn5Kx295+KRR+BfFmygZPo+xZJ11Lw+woJGMCBtecoHspYUWTshAu0CnG2UJ
BxdZ0LrxYvWWqlnMfzmiveT5poHAjVBEoSt+Ghc3Mm9WX29JnlW70+LO/JKa
llZyZD2bO5hhztnZRkte68wGNLAa1FKSRe2FZNKwT+xGT3wzm8579iKPDblq
16pXF/b8EvOgLB5zSb2iFZOwg/KcM1Xq6CulUe/edexcq7VW/pRaKvIJOMvq
xdILo2+RCnmwmEkFn65D74MO8KcZ5m0nbl+BWLYVOQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZSiXal8nPQlH/AM7uaFXPJ7XNHCGzS+7UbmFcrm8mTOjGmkcYmFHe5Wo45BB
LP/4GZDQm8t2RXFS3wN/Hrp2C+VFCR1Nn+dZtc9qDX2MZFvaUxmmIgYHLObI
+TTZ8M+ANuGnboQnN8f/0ykc74eArcmm8QH4BgUZCZD/QUkMXFUcjJFYLKO0
jPbM7fBEuKHXJLCYs5BoYgTn0yhh8je2fTXLkPD5LCWTL7ipFR8u6gTU5sg1
yW7rGiLUwGaIPP2NIo40Y+4c1pA0clj1WusiHzJUmCnDFhKotekU1g6n41TL
dWRPgcYGxdRGsiplOQhJxvoQ7sVDuetS/iyO7XMcmg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
K9+ZYQPaCwfTWKoPv8ngW7SsuUseMVL1u+TACMeIPTJVEqXLqBwCBkavFLGP
ksn651BNz5/BlMGm3w9cIFQMCEetfH98glhMTZEdIXSinIqfELo8fGxciKd1
hgV3HY8g5dr8NDK5JGORkDw2n2aFFL77EGElemUeP8fhRDKeNvhlGezMz/BP
7ZlaQFe80UWhOQDqanZ5xdd2u84Uwxo4rZVDtC4p3CjwqIukTIDTeuYdeEGv
zRT4sJ21LdyE33IH/bSPJzcr5fxr4uO0vZfmKD5kiSnjT+oxOmT8nOcRd/3z
+QeyzJldQebcqEC37ugy/YGXr3Su/jrQ3cd8h1/htA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gsfhrV9O1j5W3yUAggWIo3Ejqvf5/IOMq2bjPzlsRHq77carhtQMQkqdDiQY
gh0/mKQIEJY0dqT91M2oiriKnbsUrA5HRaBnGEZtSmtXeHEsIzQT9Zyb4wWp
nvnKisuMlU0mEwG/08OHgTILnQejYyiub6uQk9SllAxPahLj+4Y=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
jx/8Oa31pajqo4PWCrCeC2wgyfuhWjX6If++UK8Bd9hDw8OkXqe1mWgNGKoI
Ueq2y/ipgmKQinKdM/jMdp+eRZKN/U9YR57+GOg29iLp6Bb4FnS4aTmOcEd4
tzSdOy8EFCYfknu6mW2G0zAePDS6aqFvzc3cye/iSH+48a3+3p4Hxm8X4FMe
EbqbyFIFrcpAQNS096g5I3UHDNGSk478B6xsCwjq91D/1eNM7hYtNbuZT0hY
rp3I637QDkB6BwqY4bQ5kO7+5T95iO87+thuG2RadopMFx39o0qsbFUG9yUo
jsGbFc7k4WBi8E8vaduVtnhU2Q77Zwd7VqxrRO/M9urMTZ++32hpRk1fjcjP
INCKYeI3VP0TuzCLjKDKAcaif7EJwrDp/9z9k6nig90xyasK7+juofZ61RZ+
2reG0BBMT0l6BbqY9U2BsK1mjqfASWMY4lTQ/+vKOKGtMFuDEZeL197nK+1c
Ntl6zdrnJXlnMOGHsx+x3MQCGPWAVxAG


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
M8KlqKasBYdU/+QuuoSJETmHuwId/965s0Nkh3eVNj2QSXclVB8Dbsd38CRj
QAHaxbfT7j/HLF/vGU579zahFHJ+tKhDJKIkl4MImm1SnyOhCIKq00ynY4gw
DRrq3N9mIqFuBmaXeT7KKNjOyFgALToJJ35WDw5r4pe0IO9kuwI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LjJFZDgSaQ2fE5u3tyKrW7nP+a/miF0ZOBWE8Dq+z/sZqtLQ3T+mz9W01z/Z
l+rKX8yUEA9HgljPiemrC/L+FR4QOqkUYPauXa13hknhlBGBrfl59skgyVFA
r+g5zlXHzy7T1YBDuxz505T6MPR1AssJnBgz5j4SrrU5TbY8b3g=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1312)
`pragma protect data_block
IJjiTsJrM31RoHJ2ZhNWyKjxzfSuGH8SL+RTIbf/+ejgmd/VcEPmh7B+FyzR
BSb7o2odaYLEy0ub7PYOYK3o1DGQfwomamaKyIOX0G8F82p7luwR3YYxX58x
E85S97QysAK9Nu+AukJoHZD/bq4EsC6it/aRCV8T7WXmJ1j1cE32lgWpHaBv
wuSf4BCqBb6QWFrTSGcFdAyTh0dj4/WotTUjFVs7++w8aTO08Eku0wtZMDS2
8VU//2SzKHz9X0qu9SMBAtioca9duqoy6C8zWaQvJ1N5GpWk8+TKEoUHSw9G
kmviHAE6AZ7HEJb6kh5zGQTQAVYIOKkpx0PRNUfz8f6keg7kjthJHHOiQLI0
ofZNomhv/wx5M8jDrF/I2kU8ff1/mEK0JNRHZBdzsItWAufEuntLrgeXVqMq
vEDGFdBisq68oPDNud0WOHPcnhOuLipxvOnejPHm+WnxCJP/hEO+7jZ9g4l+
qvzVvDLzcx53sYp8SKasikx39MFjXHFuNANJVRdKTU25upBz5UINcVD0tbTM
sD2YIvL4nezxlBjkC3bbc4Rdwae/YYlJfmk87FRUwp1Svxlwy3Dk/g9XjSvH
54FXhUSSsltrGRB0i51HulIkYcpffc+lKVeCdtWJ/ExKkJe4vR4vfHUJ1jLh
I5wpiUzEvhP99N3XmeyeuZQdxDxNrbKESljaj4YFhbqaRrV6VfH2BflriNrU
6AY9ucZcbuQHDNC3nybqXxFfxiYPQ/ZpHLuRp7peYVFScryv1aT743BkkOz/
V0jsU99Ak/ONNRKb/eA8BwQ4x07rmhKJMddYqjRA+N5ccfd+vgji7/F4lOJo
LSMEdmezzjWTpCEa+EMunkqGZ8xPYIzPWFaIo1c85HXTyTKwIgjgk55WeKdB
q0Tf0Vib9JgCgA75mDkaCIXZxbH8ZPzd0DrOC8yoP+/KD5fLzj2lOaDX4fu9
aFygmnnV1q849M/Wm3BwA0mf3VC9tR5pPz/xIe+tMEW/PUxve+kEsSRDZY7H
pyz3TdTZpYbSXo/kjzQBQsiwNdph1deBbUsxOh1vRd7cF0muFsrQNMPECCNh
sNR/9vhephwsLed0EJmaJLPmvxu5Crrc77DoIssRMx3SIua3uua0iqkenmyC
WIwbSe4zbWBuOc8L1Y7nrGBkgt33Uk52TdMMqQNT9LTMEy9NpNkwyFXqPsB+
OAvU2Za1atOAsJhPUY6WhMHdhMvMFHanweG9Z9mMUARCWNwejT3+6pSQvhHa
zkcQ4biM7yop0DG9BGnXrEcXoCGjpHmPXD8r6WsaCSzLTjEfQGZyOdXf2pav
Wty1zUinfvy1SHzJOmoWml7cPJQn1TUtIOu0YM7Y8y2FYjtpj6SLMyrsdUUD
PYa41V+tUkBJUGIMceX8B7eksveBhZCF5FLvfkKi6A+GmHEAGpKlEfS6xJS3
LJ2csXcy7m1KIySpkEHyRQ3sqq1uDVOVblF3du6fAIUiuqhyCclHBRwzCVyo
UN2I1j5AlSNYx+jHHguDdJ8X4c48u9BCwoPqMcEpGJMCYTeZnWV/GRskr/sT
2HgHbkBKVRfu+fiPYZxGy6VPFm9DCdrdR0WNoMEArMbv4zA8sQ8cZd6oMNF9
PiQXQ6/AGSJzFsSJfgkSBq0qd1kqsaQ0xBEmiVYgKe3PkuPidM5d+HDxUvVG
NlhGy58Ulg8rb+34Z7cdj4JvGK5sULi1/qE0CGUoy2r02MGvuDLktBCj+CJg
bFC5Qe2fjw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqckm3mrGl0/8fPDvDwWC+JUUW/asUxFungS2jrYn6R8JQMgGKHHseT477ZtKXYeFW/wLniJRVDEVn5pR7BFhJEcIKde3z0K/oP+P6gVmejEQdjJVE2+3fOFEdM3bWxCNNN8guv0OqGiYtyApXxFPKYN8rpSWg3FhiBvAOUhu7NcLLzwkxmmXAW/jwx72oyexvhfi1TdQwajG0I4wfEv1ihJl5RFwPgxofXT0r2DxizmIgdgIPXj0i/JG6JV8NbuAnqbVlvmAZ2bdAlaZV0/Gd7cNEL1M8QcaGjGXt3F4oT37FAFcLtPY1EcJmNtF92wYn2PqNe+lKoCnivVdEnlxURA6oJ6h6WKGqtAm9bFLo100efpSxcaOAEF27606e/uBtO7rD+Ef4prSGJh3pNN0sk4y8/Edvm711NLggal35Ujwnb86Durk1FiwZDFFmwvUXESfybZ7wBRscNFu3qZMNUL9vJiz//aIhrG3X4lJBMz+gZRQSLo3KDgEWaF3bpmiYi+C+3j6/nV5qIXkSMlVeyEzV4Ph2gnB9ADyToxteJXRZ2sgMbulAFdn2XD9POmuKoa7LzfxgBNYk3hHfZ54EPlyUwGup+OCAiiWPW1EQy5PLWubjox5PELRBU5iC0/KJS1v4OnQ5Z990flxlx1kT8C0mjSlji4rR8gf5JMelw7VyRmAYLOLy6UDeidkIxXzivgMJbyvteeNXImjyUC5lThb7dHiMiX9No23N9hAjHt2C8goMR7pVS25M8iv3s0vtod7xvEiyrf/lcM2cokcA9s"
`endif