// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dVM47Fs+W9fDah4ZuhAw0GNzSsXzagQsykmfLXHEH/Eu3ezS3QslQQRVfpR8
8EjOzYwj5YrtTVlh07/RVCXi8BeXKnD1XkOmKYtXXmMJFb6sbDL3TQAFjlWj
QZyM7RR0s/TG2mKzS/EHH7zDlz6Asbz007Sbvn8S5ll0wnGeNPuTlDye/l5W
iok8wWDkFHmHRB6FHo30uKf1cuu7z2q7G8k8rxftjy76OSkbtBRNSOgTXVGl
dishjy4jGKpZt3W22Oqo++4iDQQdWVvOT390PXuTjoTHG5M21vhKTSowIFH1
brnnCFB50taFFR1coq0dVQs0DfpF2sbn/1ih23YAow==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fcegyvTXgRAdDy3817wvrAUuepZ/VHLL2A/1/YxATu5ANlrRPpNf1E6pPwE7
Kah1eX6vE9FYScWZ1sDGkjGDPLqzJ5S/ZMHCzrL6/kBmkbvuSNBxRG6dK0El
lSa3r2BVI/UKn97F+RsDyiG4s22BIl5U4hyqIyPb1m4BWqnk7m0MHjYRrVuI
rCzZaNbl0xYorTT24DDoA/c3vzIL01vmxphQhZgXkSGwAkE2x7J4QC1bz8KG
jima5FZZPYcizBX9dGj6kPcjf67ppU3LNMRo/0QqEKuyO7ByM7Oq7z9NB6Yu
6V2m+SMhPzXbb+oZg5/r0ysolr+9eUn/cBevkFsy7g==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TiFCELjZuckHek+p3UoselHE7hnxGzNtAe85sCufY3hz0ztvsKqTSs1q1JcU
TIxiHCZLNDyGHPafc6VTBloYawh4Ztm77ts4k6ZaIDgAkqp5XynpJBQtltGQ
qpi1igiNFadsGHr3qFPP5a4GW5QYZ5PdBea/iTTH6iUPuvjPvY8DwUGDBD2i
Fnn7o8nElTNl03++imT3KZZpzDaWMuM/lPlpST2MdMjUz0u311nqMbZWHUgb
k+HCh235DjaT/HkrOG1ZY9KsuqpFOfAGAxpL8trZnK5zodyWg9Ld168Hncfn
Kg+MjmkSoiQ5BI68XMhdVIOq7mYBI/+P6l2UsGIN/A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UFgCq4LhJ3FJ3wJAfQDOsVSHRTehOqp4bQaMVAoIXRp13uVAwPsnj0nbD9qY
zi10Tu+lV/sF70rYpTspgoHW4eLONZ6DgCEe/0kFSACoJW6RqYnmRZFfhW04
MpEHm+nbIcvVwbic3mtrqBp6YXgPJ4zvMg1cVk4Y5sEjAMkIUA3UTOhp7bnW
GgF0F4h7+bjMlayyMHerq1i/rxJlfEyb/Kr9ve2U4/uYqnLqfLzErck9G3w2
YDn8kFhU+5AJPhgQR/zptSo1vU0+EXVA/VAL7grqYdm5momUnWxmNswaaDBB
h7vP0NKC8X42NzMOg8LFcJvZ15GSEmCAbjMmFrTQ0g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Hvm35Th5AqFafQCl3/Ug7Rjw9i0m/8WgsdYyZD1i4RnIeHuC2eIVLKLKksAe
3eV1STmx/ojEsvoo99dJGipMJxqKaSW+7kjyN+lRj4LxIsO6mkxrM+5q49ne
4nEK+7clWtdZ8BoQ877tWu1Or9zDDTpTY1Eu1Af0O5H5EJHjcWs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
epSLoShkKelYcxTLog60T6Vots6DMDK2B3bWobdSrYM/NMikb26AUDrMI4A4
skzrzLb2NU6IR2b0US7CTatmTJsj+51nUMS2829Gf9FowXjB9hHSq5YPknH+
a411BuWdrcZVgdp6yEb35b3Sknk629ClVntQQqs9pmKc48PXwbV4nA2q5Ovu
VnjqTvEQxQL1nAMIOjOzQmivfzGfDnqrtS1t2gcPb0vrY7zwDzipyLlaW9I1
UWe4/AIxwGZgEhdHrRMBCrGXmii4iLXpMzrnOkSZPE7KR7THuAAui3KceTwH
VSLYc100jdaAtGhp5PiLk4Am8i5MfgRi0cLFIlD8Ah0BckVp58oG94zR/FmC
keAauMwXk9a6lPyQ8VtQUDc22QzwawR00a52x5cmk2LkGjHzNDSExMg+v4a1
977MAi8EHoSpDsPDADlrKIeDyA2el/EAKXhCzOFNosmsDdDJP8QM22C5As81
oaoW1SWLmq9kwdLq05UiiKTVaPFWdpTa


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jvK88tGgK4r8YY0JoeM6hK+fWhYWbcNOxcoT+MmPoHNsmq4HOFiNXHkMN/iq
UIrhpx+kRFdXItqADEhyLhWIivcZF9MvJq1IJnvCIlxAyvuAoqSTgRbHw4K4
6tHkch04affCoR4WF7UHDdCYH8emuPy7IOscPBpyhwjsQfAshNo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MD7FCPL3S+aREY7GLOiZVYHX5vY5lwX56xXewflxpUsGDRYU9yAf8mvPM+CE
mAMPIa+OFneM/du2rxvJay65gg4nUGf5Km5CiOdR6XsAHRi8e3/4LEMHUbl5
YuVgcqy9Mp0oKqwUqswgLhUA/uOEMGj+1UYWXD/aBFh3K0wI7YI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 16896)
`pragma protect data_block
Nk20kviOK0uAm9xzb1cQzv0rd3zjfpCsdSg2WLBoJE2igm88EPDF+Xv5DBF/
iWqZ3DkiLIcYu6h6tocK0QIVxLicN/LFBAUsg2LQLeFR+0zJ/gZsNYYH15kY
mCfYNutngUpa3X8ZxipUGiervTln+b9FxvbwK57pDUHxv/4Ol6MovsaG64g8
cR61MpJ3zfNow6IkdvPrQYJ9BDF21TYbcFTCIKv12Q3PYQBMTmo9SiVHoTS3
dRDrhMDuqYGt7X16kmva3DWcLXUv6FTsx2dlFBdjqUFwFgJu1Vb3VZjdMj3f
NtJEx00ymetiuz/jnRs99n8rjQGyd3hJXBb5Z5pq5JoUSOGilriHb4QLzWgy
54MDY+qIgDFSwgVmHOyYuRP5f0Sd7qXlXrpWks+Da20PyhlLckgfBAosfzCf
HTk9tMedHOjMHmISdAdR/gxYGQaW4qkYm8ljenJPQcnSVXURHn7UccFtXJKn
yQR5imfGucXZ6orNYQiISLhd39zXSIMm6/Rko270wmG5lhSTWtsshTc5gLVG
1334zr0gK7as8QcJWpb7t+eK/qOghixINM9JjfLDs8U9F10ZYo97/SmksKG4
FU7FtI8xTPqOkI6YtDwM7rZNXCrsGgscLWnIHCc7lZXeXatqYCwJhvUHnHAM
WI39H8/RO5QdhTiPrYXh2hto1vBBhg/0pmX6iOxQwa8GRNsLvxzn8/g3L+qX
H8AqH8atQlCZMj9q3wmlnKxYBW2qHqKK1/lehCwtkeap2ouuhuyetSsxj1Yc
6AN9Re97Mp7UfIFYQV3WLmkKDhsTsFTeyzzAlUp9r+zBVFkn8mNOTyf1gKRf
RNCa0g5upm+QVDx+EPqDexVtUXmQywcXomRdC8J1O4kC78uC3DvcgVlUeuZz
T7S/eMUoXv6Lx7m2XWUazw/lJ6ZOBxfH7n0DO4gYpNcunVhrW1y570HmX8BR
xTOaBC/OwmisckqUp9gZiFChIPzT7kLeNjuzCrmdK3WJrC9DFz32couwl7KX
lCzxUNHv9Dxm8CznUgFVJCkfQa3fYQvz7gzMbeo4gnlraebhNgl5+zdKUSz5
thF+LFLdV65OosK7VTDF4DVuLlt55v1aRokkX+w+E6bEbqDtqv/nHmk6OAo6
Ulm2EoBcUf9Js9Pp/Xxt8MQLuAxpWNuo8Vg7YlUKWjU/WMuP/ObCpseKbLuX
tzRBD8merYK6QKc/lvgZefFloz7VcermvAw+grTi3avQrd7MuEfmO7ZBe9ba
rSxpSxS9nW2ExU3tLRU0ugBzRZoGwGD0waEPCpKlNJxywJt6v0YpDrx0Tpk2
BqsXOuIMTTnQCfYYdROKTB2vfDCemfG5HfuX432bxeLR59uxgzMFvyGkWAx6
dN8Hf23AKdsxWGNnqXgxV2a7mClPmhKt+idWCqz4vTn/voMhDF+U7b/dMv4l
/Lyy5+nxzti83vGgrCLLKYozxex/93LR7CX02WlIKI9xDLzXRHkBe6L1+J6z
MWBZR7cQX4O391aKLtL76y8vlZ1BUSZaufNCNCs5XS9IxpHiQkWT8uu6r6tI
yOKUYn36nFHW5bXuk/qCoHkLdTXIM8Q8WxTk6jPdmGdkPVP3//ldP43BpUzw
ZeBvy8AhXztJsmhIrX0aF3yICiLIZTTpM/Mj35nDyEIs7Dhv3O5mHNvRV1dg
3v24/GU+Unb9FMOaLQZ1Dl9mSQblrnM30I6oY2Su9X3UvXu1xz9ov8zXoGtW
VCliXxEg0e+lXHrUT8Fe7WQh/Y/ywh2yJqxBxVCzmjleTckD+WnxsAtC9IB/
o0EGCHlkR9wAoaQ/sy4aVLqVFfm0FQieX+kx0CtYJEBf08XKLmJus9Np9NoL
v2pNesMPs4RCwTaFgwVSd8NPMEZWLfxZTQQ14mLeLpbaS/kOYhF0GlKQcyma
CAUm8TdBTuEn7mHTBPHn49cC06KpznJZXQRRFRL1U6pqBI0GvLO2sEr/wkvx
s41MzrCf99HPD/wKBycO+lcwGy+sI384hUqcrzYu6u4lMf1oURB/8g87EhCR
/ET4pO9v5T7J/1JlsNIvwc4KUNrBXDxsTh44hA1NSVmDK1WUvG/kvdHxih6F
PMqjJtkaCpwEjoQJoo0sMi4i7pOteB51riKEEUwbi25qoPF5xfZZ0NSQUegx
XYeh8/yF393dzqpfM+XUXpKV3Fg2nYqvVas9Fd6tA1VAnLGGLtQtzvmJjXH6
HA9aT2WhcRDaQBMHr9zJOg8pk+ltp2oiwJP/Sjcl07ekRsH5UvcB5Lz2BCRz
i1LeAyaMGzDfKB2Ntk+p+BhuY0zvp7vbvN1ZKriVRlwPj1FzIjo8f0S7S1n5
/I0AWp3dnZ0AEHG66UqUztXYviiPKVwPxC/VNO1rmta6FWPnoBVzFJrA7tP8
lIfQAl8Q+wmD1/aBfdpeF/KZ0+gxpMCg/LEJWQRdme15SHn94LTFNCs7xPxw
uwh9DtnHD2LSJ+etOLYqWNFLKAZ8be+R/0NNfKQzjvNt36ywuXs6WDD3liCs
X6Z7mhA+CLu51NobqzFH67z4nL0++hBJZCK/cG2ykJUPwHCTLMwRPfFhlC3R
Gol5h/IPgGn87Orcl9nHOQQp5uqACbh7/nuniZFzrFM+wyf1Fv1R5kPDAVUJ
mr2k7f+ZG7jO8vtMdWUkhaPXXwXcISqcC6BppjI3zQp8OGDiKgID6jWHJ6w6
UKSBcY5vM0r+glKVN7letGY5IhX7KxKYQR4/hN1m8ma0MGykpDlFGw3ozvRl
ewuOaS17rDvhZaH5m4Lh0SMxXvQYGDQVMXsl1P1nuYkx9cRUTr+pNGQoJYFk
P7/UXT/ynS2zSjIWCV5L6oABd4VHLb2hsBJ8UoiG9JPkytbRurz+J3e13Q3C
2snftbmV6wlFZCzFF+JQfHsrMRpmggfAOyFrX3thSR01/AFCrMX8FXXrGEcK
UXvNYVEh5wy7D30hbERxjzfV8ta7ANiz+Nlj89D8YLVvoSax9g4sFBiesaYA
OctBvxZlasutlwU/46/Vh9QnZvOafMpOIXHC49tbpse9BjwLBml4MgPcn7Wg
EkAY9VH4wzKMl/TYG9QUdRhbNKQEit8mzfWTyeYDmuU3SL7eTn+OnRN1AcAy
LvOIX3YuKjc/8pY1dgg0xpmsNM0Dj/6yFxbSOZqtu/VjVsRBbmUen+M4n/6n
KXoClfmBp9vP0uasjnsZ1lpXx0LHWKZt+OWM5sEGB0vlpIg1ro6Kg7nMR7AQ
lPd0lVenNCWJLkbvv8h6qx9pvF49OBI86NkL6T9MgaTdkxfiFZfLC4pgC+ws
yYi3ejwdn824A0ArjbQZHO8HxpmbUDGkO+8BRqXClt5ZPsgrXVyUX7DC61kt
EVDZvtcFxIsAAFP9xokig+UfzpyO/de3AeWbUDw3ih5lg4OAFYgBIHzkGSem
LqijzTj5kpWg1TgSbJ/jlv4ZVU5I0kw2o2zXrSxcxtaTKM2tyuq4uSfsTl5f
COcMbkwQRBKX81hn0n/iIgIaA6XKcHsRDcWEg/narBvOe4Cav36+0TxgUQ1t
m005lm7PKj0rzESegbiwif9mPGn442z2+7eigPVmCdslSOFny5bir5Hgcfcp
QABkKxstE5SrZiP87bexKgXnQiqf2rNhMfR1E4CF22qpWwH/Nq3GeAKdKCit
Oe7ucXEbfJmjfMnli4IvBHy8Y4qzwOD2Da2kv/VjWX1wTtqiBL5cQFqQQZ2/
zIkmsDrj79HfgHYgpsKh0h+OnPuw7FxmLyGCKhujSDQLCTbQzQZxmkaqFtCX
hByCSP4a+wSB+2Ow0Qie519+KqWcO+a6DPtr4NItOGR3g1RpgODSZ79p7u8p
ZNsXvzFplUbHErDgPSxw1TjxWw6sf67Z9uT7yYVIhC3+szPIL+Heh2wFc/Ge
Jrl3OyAPGq7ybt/YSgVJclaICmMbRKUiHTnFFV5kQOLEIgH0TzPSwbWvl9ab
8TKkOPOSH4Af/j9OzcTGcINatd/GX2tTsIgtc1vN/jC9u9Y9q2VBT0L6eEg6
lJXhWnAGo/xG0jgB2Jw3MmI/FYzGqhw0EEJG8q5T7LZIvicOWACfR/QOooZx
t1jIDSvD/c27fGwVLMMyl26mqRsTiF75UBEGKWdpI5AJUr1YYNNVxsFJGIDI
/fNUrvb2cqYLUKQwXVbxoNusISUbSnlZF3rim0GmmCgVh1DxsdKH1jO7KurC
k8td65SW/uNY+nPUOsjoOg+p1+cIGZ1Ot0QeZc8bwoPSx7K5bAX+GEC4KsZn
gl7qvY20QlcYaFDzGEf3AAIhmX8Z0B1S+oj/oNeV+hHK2mkhz31+y0SQuvSf
Oa3vqyQxAZIeV0ZTcTMSsOhVvtsR9xRlAVjxLMCG0eGnRlbirdgASShxLxZQ
HlN5SLTGxMWr6ocyYva79y2+tnIFcPVWSxJ91k0IBW8Jkf82SEfpaFM5fPVA
Mbj2g4u6o97Yg9caap3ytGdVMLijKty45uAdOnsPnJgMgKx7E+3BG1ve4VKn
6pBsUgoawdDQbEDDcTuvmgUuAzssZPUxQgtqT8lsz+bBu4WTZSTvo890EIqu
NN0f+VVyzufWNS2Og+0fvVTIfn/MGeUqjtG9YuR2KgmlhnpsB0MYrJgbURCa
Xiu2X0kGtQebwXjzMwf2kfuAeTYPRcbACVCRQ+O24OEmC2cCGDaoKzPpmC3m
zw37MwDR8XOxDfikEjOZ9koOd3lBvtl8jeX7ccZ9qcRl/B/WljEAJAYtFNqH
A2rig9zXdCz4gdkRgWpW4Cbv2ck8g1uZh5t8Ex+SYwgYo1hfbytBUxqn+ovD
JtBs31/mOPxG/awb692s5lvLs2pkH51JJCwSl7nLToUEZ89tWQPRx2fzg5go
dS3YpIdhcJoLXPu/QLIIyLqoq5O6y3QjN7ANOFANbZCoK+2bHvFmr+A6pD2T
OjBO8WEXNMR/+RrmDqi4aMl8LR9w7eUbiLiLUBrjcGk16W4lCfw4CHaL6INp
auWDdr6sWOr0UaWGRf01zY3AdWsAcEwRP1xfYlhGyvcq7uhx2kFiezAXaAQ9
N6KhPxueH22PrmpkKibHU1jnkUWhl2OJ8caDqlu/gIOh4bi9PdgyW67riiJL
7Grt8yZEU2+VZH61pfC+VT2UVf6xICHq8hC40mQguy0IjxyFeRyLUKtKR+b4
AHqs1kyTe1alJzrwqPrz7qVqvjGv+t+TV7ing9PK8AwufHcpqY6DIGJ7KrUe
h2mp0uWGC9HNvrFt9EpZCRyAP62U4i0J14gf2OZTs3k+q9yDkNv0zwHdcu8Z
iLLgCjZD5g0HM19K2BO0/MQ1SwR9fJ/fX75YgJ4ycxn4z83dtemEiN63nYOJ
d7oeULE6LmKnm1GGES3tBQ1x8eneVEm7zXv5eJMT0wdkE6+eG/SI4dN6ENZi
8uTHCjxgDGlmUJTqkbgX1O1+nqpq7MWck2rBK2eLyL8bbm1t9aymWpyJGG6G
RHIL0/nYoO2g9087Hw5gdUiMKr2m7n7lwXUM8kZaH++Zpm0+oE8LJ8XppSwQ
Uw0pmpfT2I057pAqahcBsuEPCCY3OdPR/8cHUFw1T2bOqQh+qJtisOxyHcY+
6LzSHOmWdOxOjH+UcVvm8gRw5Gxzt+DWLK3IPZJVFAN2i/pIk4hzY8OIhcP+
M+T/SeCtM/rtibETHLfLsblWOM+0ppGWHD0Gn1mbIE+8AffGU1vcRhyL1hRX
rknXGzxgbjkoKc6kbB0REjUqNuT3wVZ69ZCfbn369TAaZNagvBvvuTmj6oQj
omZo/FYT3MXtFiuxOWHBlpZ6OVWUis2rqMlhNlxYMC54RDgpqyB6KLSkd51X
bYxAEs88TWknY80EwrhUJzZEFzVPCJCbNmybVXNnMhDLbmwN71pSLtsSWVP8
pJPVCHj2NiLmSHgeBW8OFGFGBfPhkHr2LrKMN5zMcwIwvkBPMNMWtDJTTMvw
1zDm6P8FLOBE/EIJ/SIMSsJY6NvWj9hQ55dvrd55aIEN2BAjqsIfd1J8GFop
SK9wbwbKZMPPQFTnm94/mIAioKYiwykwbLQRL4AKdM1RYAHG5FzfoEXKSnME
/fum93cgz8v53ke3125KFI7qYXFspeQmn4hn3xCmFE/f7wM0LDSMkV+UCmAn
Rg0B6Kpdqxa86O2sETDa2PjsYKCfc5DbSD0eP1GjsDRllioqN17m4DYskXcG
VcIVGibz0Ap/CDyqDeg/DXTa3WLu4j5bJqurvhCaNCV2coGrJQDkijrcEh6K
RkG71l4g/MEdgNCbwQ9so561xpCmLSckoJ899vZJNs6ptmCnnoiOuXR/w6sc
Wz92FmOu8KIwHYUzNJw4f31zKC37LTjXxaPGFmgpCtN056UyMy5HRtWzFNUg
hZjMsFcpEavn32S9EyPRR3R32C4p9CiXUHTFDzB6zCuedFHXfbHDljTjAc9r
uQvzKR8sK+AEfLdCnF7vdFEB7rvVUP+Wv2p103BpUrmmaDJvF+aWUyhRAIY4
4Vvb6QdNH/ZanLamCvh+F6B+PTHbZ52Jdt5Qp7p7SP/DYladS6L7ymq/F2uN
phNnunUNoeyia0p3KfR9AiTBuKtnyG8GC0zfkQiAEoPWW4iKLQt6oXHHt5sX
VcdNeiq7wk7Hjtkee4gHzL+FnCLVjg0/WUbT1rxcinOEFlzUF65q+Ig+L+YR
GPs2wr8903bXdw1P4b2VWBUKbdUfNvhlcve40xVG2SI9u2iRfnzFHdGzUWVE
ga5PIiIX4yf9P4G6fnS2bjpCXkn+Vts3Im+A6dfKzI4LPr8e5OJk+PniLNSO
wY1Jh/qWRsqP97AqSpqOcqCSL201MvwfFhVtTcwz9zw7qlIft0c6BOXCpwus
etpz1cf4IBblrd5cX4x1YntpamP9UPzXLJ0mIKsk8WPEKgi/1+w4Ta1AeWZ1
xkj4pH0idvuPP23661StT7Bu6as9F5GS0G2tBmPWnP729IcaSsWm/EFXTYN1
lTqV3TDT636l9zFlgEMrj2V539Y5OcmPZ7CwMaIRyX00zWOrpwT8eV/cTV2N
o6QhCYUUU6bt1ZbA80VWGUAftnGd+U1+pml9PG/k1KtnIlz3ba1RfuYnyy8L
8ALflWH0zYaUZiibuPpjUIFlkiPKPk1DmGFnLQxkSm38eVjLJuYFyVxTgofh
r5+hVbZASEcrxP7gT/xUXtL3e4IA9X7bwxgywf+iYzBbKMSsxif9nmY/dx/y
btY4AhQZVe74wvgkh2Mb4rsCjmaiWbTlRdg8eXBk0HmICP/ij5/jjVKTK54C
Marr78a2KMs1cPG9r4mWAJyjtFoZtx9VSn5qhqWTcD31LoJH/ZU6tQxvflIY
H5EgafgHuz7etjz6FnD9ql8+xSNFYMwSwfhlUhz34e7f+gdFq+Nrhj4BV2mk
aHOvutWJDnY91c8FKWy6IE3dCTjBdAKQsdO+WG6uzBHMVlKlCTtCsPzEn8VI
gwMMUaEFZtuxvuMUVp5QW1EUpV0RoauuArjpnw95o2kzJb32A4I/zH4bYtAF
APfzuvFQj9fIwFB8hXyGrDmQVkFp6GEBpe24ehtjR1dC7HcfStgzXGmMvtTB
OHA8f0e14ODBbsIR+4KNFeHvpYAMb6Kxp6W0k58taP5gpYsheOmh/uxS5Cez
jZvYFTN61H3i3YWYfkkoXL/WMWxKfjQOyzKrvCyU9OgtBmxGPKnPB5X8cSLe
gbWhOtKq4VRQHAZM6FhpD0fv4YR+JnJNSi15+iAYK3So6qiPkNMG7u3tOsGW
hlYa1DLpffFll3koyVWtUJ7RbD9CnxVuJcBkF0bl5mTomD3zMKa6ZJHeTLSv
VL+c+syVLQAqPOoo6C9wsx3h7EdZiT43lt4fvw9PoK3Bf5828T38VkeXjf6x
zHKZ7h48GgjtTTsIAsvtEvwDMD2kTg3YTknY6PyCami6N3JI3qAcM/4P7RtG
0sGmxb30iYN3AlRt2zVYGunkqlKa3NseMv+A2IJNbvmOV+sKnQz1wCsa/ndT
TDNa2HJw8X0uqpluUCb7um4xgemP6v31QADauuZZuoN7PyJR15x9E63jJZ1K
wJwgGozGZTbpaT6w8jWWfksoqv0aHuKaHJvI6JIyJljjkTWfihO4wtU+EkJf
NabO/sHx6lQ4Vv2tTg2lMpFbFMeWucUXyRsvZ8LD1EEfBPD5ecEhg2Cd0OzX
17uRLua7YWxrS+BmOPrqWHkL1VGbetLckNEvWO9wtFgRzWV/JJlgmtVSbdbY
J0NDhJyhY0MK56upFwxYBIlOF5oc6SfZWRJcAUO+k8hB3f04By2eY0oX4v2y
APd+xLo9B9ESwNTmRWLkMh/LjUdW9EBgh/GKaesHCMNe31jOeNF5o59Hav8w
xySgRkMYBJS/9PopVfYcThiDDVybJ52wPz9Y8WLBpDv9+aslvWeaWKHTxWX5
y9HWIdmrzBUAsxxr/IXK99g6mP4a+ykEh/ICP5pIPg+E6IiFOZ4ljpN4AdBQ
ByNwSCSBgcRkIvdFYOxxCXexKuZ3XCnDKsDB/T4DR1A1xc2ZW7P6DMs2nAh4
p9c3coPptYQOoah9pcphn4VG0mlo0+dCokXXqRpc8Gn91CGNCUM2vDh0Gh/M
Gcf32seJGSp+qpa0Gpm1XNHZqH7AtemYhV9yuJ2VRhGgUVv/YAqEedFyFlWa
SHFuGbCRLBHdJRzQ/1UJE7E3CtcLFyDbzaZssyaI5bjP8It9spplOqoL4gVN
AFjji786sKRdblpZ1m3VF6UgYoXIN7aJ8C8ttA0o5m2k9fO6AwjHvMhnHD6S
CtQg8S9x/gF4A7UxcWlu5Y65WfYfit4IOWN2KF/Jezt1lnV/Mtpwrn7JsVwW
662UmA5wJF6UYIq5CoOf4GEp71OeNMwQLJSYv5Cy0nkZBb0WHeWQuh5eKtj3
qJb84oF86nJw+YJnLM13mefsB5dMrhSR1GNAoVyR8eGbUbJMFayaHiaQk2DR
WQaVtBNTHwVZLzNyAwEolDgwxmRNknGNwPHuAeRBAwJvTdlRrzShHIynCeL5
gWyLNhGVtYApEsynVMTnBhDLXl05Rn2hlmepNq+6kWi5OQ+uTF4hzae5fog6
pyXWwsrhIB27ApIgc/ZTr+47BVH0bcp2wHdJub+F9oSFAHn6DoRXi0Ct/LxM
wGf5AVlPAh/ahxDBx1iv4nA1Kcpj/E484D1fV/9vnMO2PBOUcyVebzuHL3QJ
KoZwHjMtF72Kw66YiAfwDAgEoyoxur01Zq10iW04OhSMTqBVzNX54qYsxmVV
f7fQNVqoW34PLBGq9dFxv2ZgjF9n4Lm4F1nC1knVVON0VSB8lChcR499EooY
sGXyPM4iRemLbuBs1EztXwsEMAaN2aRHkHTT0ZMKQ18RKPtYzSHs6fMOS24Y
3TMUqz3KH4qra7NGys4Dlad0NMO3K4IPyv5PUO5qgDIQlHpEkVUyDWvQ0Rf8
MeF2U3tZQkVqk/4pETuu0VxPtIbZNqslTxk2yGKVEYP05/8nwg5lUKJFCs/q
azudHPmasNM8W+jL7kcH29i2th1upLxe12fJF0twNRkj1rXgeW48n5uGGvky
iv1gsjV1FQhDWtzfNWEBJ+QeBql5aS8/i6sv7deOEyuYWcj8NPoL91wVkkXP
vLCbGKHqof0tXVltyFcGHQG8R4jTMCdM41WcoOiFtfO6Fq+WGTWnXMZrlkuS
4FBLC20cknUDIj90+HrSJQrTUeix4kxk7dGmsaAI4ymiuLi3gyHu7E9yilPD
JB+c3FDfKn3so5LybAaPXdMHjKmab8f9fhM8FF/AEGtlFAKpZ5V8xasB06j8
DLrkfgonYVrPvNkQJv/ZySHkonTX0PnYAIjubJpaZiNHmJMAs316BGOwi1pg
3psY36FEKbQOF/y5TtRgsOjUCIKy4yDjqT1oPQAx95BnaNm0hQhZuMChzZ6b
mo4Ei5+RCHxG29F47zok/STKqb8BySwwKM93x1nTfqIX+cRaUhg1CsZfpmy4
OJXStxB6MNlXHh+ZNKDTsHR7zkzWpalZEiOLQNSLHhYR5OIPhE56oD/MfeWe
+ymG8QcRQqmdhc4SGzoH1BRDBAgqZ9DyZfmeI1WwAN7+ouZNlBs4jGp/DtCA
9dFK1uohMQxuUm02vnUUZyEeqkvk5eN9co5XsbWhLc0UwUaDxhYV59B0Vbrw
ZCo6VGLIdke2bliPSx2b+VEIJrXZMrHbkM79DNKRhQ38h5nPWEIC6eGLsXF0
yDkCumhJgi0sL3VBRa2nIvfekkU9GSaqqi/oXAjY/0YRBa3G+s15JqA61cFZ
Lml1kRf/vpx4JJ1vcrPvRgCuGROLjbKwgiRRIOqSOpdqlt4Y4TpuQEbu0un+
CGkOnrQSWJykYqcpAdmsHoTYtlRkLwSDFdtlCjYaFu92PsUt6Dh92/T4cjIg
8Wq55JKAmP/JTtuQPvbci04C+2qE2cfOOb19FI7hB+ygIlYYn+Li9J5DP083
UDNJJdlReLzsiImZv9lzhLzIccauiD9C3d53mS7SDmh+MHD4t50Hjl6pJwnF
HoTuIF7j/zKlTdIH984srfa/e2z4myMjEHJuAqb6kvTdKGCmd5M0F21qvmnI
eG8esmA3JIYcKdrdAcmx3mdL2M8LgAST/3ElCh/Q8FSejSGeBKiL87oBSOro
ZraqOZuP3uUNlq8UNFQdufDlKb9Q2PWjysmci4k34hYyN7XUywWaDNuthYVh
T+exammI2kZuwfp3dth5RLVNHD7M6vujiy+tjJu5zsg8QWlOYhC+BBMeT0Q8
kvTF+WJjbNRmJ5kOfAqXq2lwkvw+Javrg56rcYLiCBmjprbppgZvnayliLNq
kSKJ7YzoFxH4ithgXe6NCHRG3gnF/CnkfPTvR12FyDrUQVM3FJFApgEWDU5Q
L4o4wU/lkg1PNpC2f1qRm2MRIX3pS08d3kNL0PO8OIJJXJhIeqBWvZvVx7+d
dHakCr6SVVtThkevNe1QOiyvXKn/6e6QUCctnBJRvlJo3L8LVIt/zKpd8O6W
ZPCVAT8LF78YfhrlEYG08grxvQeSifAXB7KDu1AcArmP7mTSsaJbshUXJei7
X8hmNjOH6JRQgYS177gfk/jkW6VoeRYE0Fp/lU7H4ZP3QQFq2fw+Mx5THZu/
f6HnCSXRVfKp5Oa9lbq0RC9RQERTbngwsoNYWXpFNrrEReLqQSgh/tvP5+0j
c17ujNqoUc+w36jYkpGOCedLOzoelCgQ9bShOdOXD8swCGsB0tOSx+nYqFom
qoSBz0DeOioVnkbP7AuRjEiiQFH1UGKoqWXVBCen0x9oD88aYFA21ffi9CK+
E6jE74Tcc3Bb0JJ/YVkDZFILtABs28n6ZNcJunu0tnwSdkeUsvH5/AOZcEzj
g3K+ETG0gCfo44v2EakDuAPA74KuJn9oS5up0Qzp6jXpZFm7qJfrdCwmIHMX
ZiDA/zmbErX5U7uRy/pa6la3TmK7arJmzRDKJ+gTMAk2ZKHZCSIprhhm16+E
5psof+BPnEvSczLwbtG9TNceZJB1otmbtOXu/Onph88//6DDlCihFLMUej12
gvYW4h8GvWueL3Kq8TxCTv4TS4MvttE2FUIWn7UYUn9IBtZzGUin4XnDaaXd
5esVOFpCD90wkiKQeSMlo/3rBnZm6XsJmZ3q/KOCIjFdmEsiLSQfct/awMxa
p092FOJkx2IjCvOcvAt0mRp3myY7e7BLOv4JFIz0QKDugICJuwMaPhLKqIdR
2xvzqZq6G7VUICVZaeZj6gW7ENvAtBmxNHqH346jKClUn912K5Lnay5RAXqw
PIZndXiQRSx12LoM4rLki4cbxb9SpEI8Yz2aheblsuScFlPSVGFL1Vtt52PJ
YWlW48B8K9HXvc7Nnxa5VKxrA8Xk1ycs1FgYjmjYtcf6jz577FK8wi0dc0BU
XC/A8zBQPuUTe/UMGWlpikN4dXnEiDlAjROYpR7lksv3LQyqZuQtitIYlJ2K
WkwCnKaDJ0hiL8uuHqMgsCPGr3JhjAuDQ++YAEL2AiMlA7yg3Dr+wkeuDeBv
u6mlo2Ooevbth4k5iBctPmV9AAX4amBnqV7fjQflv4HuAqBuP6ChUm1YEjjE
X2TYxTBCaRWUSma1lRJKH16jYq6ov8bjZb9h6oZMNfRRxPwDIrLtP2EMfH24
4LQH4dJb2Ajoh9GeR67Uid+gectNKWisu/YjUf7KL4o5iO9p6gw4z5G9MhVN
tnEhITZfSX2lBDGvSP4y063dBPLGor4rCr9K0GyRP1LSFpDKfYqnG1AOluj9
zo5y8Lm1/W/sbTFkq+kSE33lI/vBExclLQgLq9LsJY4nYa17kfuDPSimxTuv
ThY6SXzBxVBpStl2T4OIBj9s3swIfiULVPc5SZm14XPAJJ4ZryDzPGISgR5z
m2DJaeXLEVRqx/O2YPJxn4Zr/dHLWn/HDAEo6yxrHPZDTrrgc9scJUvlromr
OqQHtRxGHeehV2GI1kKOspr10c6EsePCYyHU/79BXg7+Xinls5WFg9QtEO8P
7GgD28qOADb2mLihuyz/7NtHaPu5JNrJHmcpBIwhdn7LgRn/KaHMvha8gJqg
chPqCIaUB9mX6XnKCCToVPOzQquH24+zcr+Nqp2l/axZCajGy4sVJTHBzwUl
D2NDV9WiSGnxWwowgOdRx4pjgTMjvoybCXuyBN2AVoS9sxSAUxE8nKZkHBFH
7JQpvaKsgPv3zpibt+bPqO6H2Ap80ksXHcD2p9bDVKntdtyUtZ5qCcmSVLaK
Rqo4plsAJiGEADjImQLwlZGPfA88Yin39OWid7PcWKbB/x/C1b3cbI1KALT5
a026e2z1Cp6GM9GzXRVFV7NJoJTSVXwgQeDSsKETWfjnYGwf4eFJPGDetixf
M/pNJ6ksSAd4Pyk3z1h8vIlbB+EJCzW5hjImyF9QcVuzn6QNaJ5lLvaLax++
yzw0vafMIHPFhdXigNmxTt9Dyisw5aifV59jkF/yPknt1bJ6dTyjSU9SjvGU
57pBG/afUAZkXyMNyeFixJUI4vS5HPHdoK0vp8CFsJP6pBHkzUC37+YOJWSJ
/UGIl/etLo4+X0vKUtlF9VmX41c98trjVnj9oil0ca1t50TguU6U+DG3B4mR
adgR2D1Dicc5e4buMNCZvq6CT9mNzfmwU+/bdvoZNNO//ZR08BKBvMaUPNFu
DPfeJKmXqzUGASRozGuizm3oVJziaNB5yO43viorW1AQOQPcHXOthCBW03uA
ZAw5YyCRCrh2VRyLS0twyfQvx5KCxN16tl1Zdk5os4WUJbqy+WvaL+uA1oRY
sQdI6fj077YoFVayhS/JxNWJI7CEbm0pi5YoCkqrWmxSt95HBTAGCjEfvO1x
7EZqSQHzGRgdagFUY1rGf7G/qmCVBP4AHElp/5gflExnfqgOPAaVuY4kPs2s
ElZ0MQbr6sRHrHHKqJXuxGAbM1ruwxKoC0whhMMBisRkglV+fXzTVnoT3MXk
3iNHwf6i1HTg4KOaXNfQoVp67TCUtyb9908H5Q0bkO/IWCQJuDJ4pDDF/7W5
ppwn9WEflnvRo5Bso9lFTZYTDWipomF4rslmOEqjlwzRiuhk0XwSU+tRiueo
G7Jg8cYLAiozrzyRVlKN4BrrNSLoku4XvkfLqpfuGJEIbFgjT1d2xHdV2PQR
tNB/OkNu411ghmMfAnKO5f6qkV5YZBKg6gGqTZndOdnRA5sAhpOOwMq96Y+k
sg2UJjCFTNNdVTH0Umc4BeoYWqaT5+T/APt66smuW7GzEyCN2/Irm3xGEUek
/605n6OyAUR8jjg3OkL/eO9OVEEl3sKkLUQYAmIwFEEOq6o4IekYq4Pa3Smt
+ZPDfi/m2x+9J9bNLyMPkxRCK48JwSMdOexaYQ6jwFwqzxHon5SvjHSTdNGY
2/YzK8+/lncbR6Z/Hfn9Lv7U0gWiAGVPzvou8z7d5RBWp5/490GYLSxlWDUn
gtTz3JYRfu1hgEeTIp2dz/daSd6SEP26T1Xakmup1559X1YGVS/wD2vuPJNv
thz7zPjuXEMyYHtQm4SSFlhvQxJ2dTlI6nwe6kH+4ofRfOf43XFEJN83ykw1
iLKhJoiDSc2wbUDlAYH9o8mGBMxOt3x0V5RMDeDPWbIFiD37+patOcT2PJ4H
ITX6Yh1UWKqo4QWdVUrQNFts4eyueuQzh7VLWUHliIWNDD4VjeXADt7fYL4j
/EyD954wxhcAit2ZfbOMRzlI3bCbmuNtRDOMLhiq8ic1YlCvYwacHOShzumW
0kT4v06LpjH+pofOMqNrpn9eW07KbF2q/8Ao4MkzGyZGOMe7yulQv8wJgPXG
fjuakpjUgeLPBz5tiYGJuZrdGoCVncruuK7uuqpfAlTt3ufIgImFmRmhHscU
raGcazys3F+6S9d5YL6oAiFBT4E3VwuiX2OCq/Ge6M52w7+aVkU+iLem8/Y5
UPS9xBFlwCgMeFYuUjP5YpBNiXARaUyqxD1icKTPAboaFXoOFi+Jr/1rP8vd
lyq/Rva1RDScBaU9yMqhFmOhm6CnwwarTldtbDC3tBhMojWSa/fipfCBR30d
cXWi74vJChFPFr6szYb+0IAwnq8A+Zaiu2s55rfVJGlQuJc4G+hyK5DUReTK
KlMqvPgsrqffj/mMkW9Cm4y+UBKEj+wAJE2x9lrvk/KsYFgD0BrKsu2hyV2t
XaHcGT9Cd+fhVQ2WwDP4jd7m9mE8rCArN9E1OPVCjtvtwGrqTcgwb4GHkxN+
aIUKG7VPFSGCrE9mSaVI0wyIuB5H2JcFRlssj0/3rTUfgb6Qb1/Hb7/WUGt+
K60cDlfcuEkuDEhzCKwghiwBgyKWg8g/HDhDi1plYbNsr+OPCj4/dY4CeNbX
bGQwrALtZDkyIz7EzifwLP1SWeLpPrZmdinBAP95esI4muVYPSDA3orhbhoK
yeayVih4wPC6oTRxdXv3bDyeUrwdz9BQ6vCQMR7l262XKPZ9tyJtON+hOBtc
6Egf0SN3ZbwplsxMCkbC4gaxJvinDQVzTf801iibP2Qg8iA33SijSmjB8BQc
UbwZi9uj6IPCw46av6WIMs4LSjZdIFOl41YaS6yrsGHcgtGqUTDv99p4kERo
9fCavIKnBJgKOP1bhIs3AUsklTqDUDiGBnMBV43XZyuhyWNOq7jfYa2kM7l/
yzE5VpBvTMUtlXGYrrFMLOhMWTEPrJUo6wGni0E8GisrF2d+Esdh/58Jnswb
cvs68mMLJnl9uJ9Dpq04UD0otlAwWmkpFPlnRCzzhBm8BuVtfDqXs1KPUyn7
l5HBxESPXxrYFDVWghFR8Zqa+6JaPl7LiZTzcpk6vrLM5U2x7jRcqNrzqHbd
IgTcq6OFXrUHWXM/De0uR5/Y4mx/Xe1N1A3nh2M2JeZqKE1R1xwMqML+4A/Y
lmPJ1YeLPzosMyP3LT55GFbJ+Ha88oDwcDUCjQ5kL4vKXDSRh/y/1vkKGp1+
V99xmJ0LejgcE0AlMQ51BEMTW4REf+KmcX3lsO1VQGfnVkPpzN3T5Ige/EKt
wKlwA/w+z28H5GqMtJJzHR2YLLp2qj7CCFU42QMG1zL8QdnGdzKzw6LB7oQy
1aMoUMNPNnJ1ktJv+bmQ4k3nPAyYnNkbmYhoPQkQeV9j4vaJHL6wbV8OV555
W0Hc4RsVw4yB64nuQqWjNFODDtDNUUaFywBXYdS4IzWX13aQkhaQcNpH51Vk
3l49+1ftrJu1M/AGSUy8r7cnsgdhq/GHPlOCgK7KlUiTNYriUIn5H5RDvEP7
kwZMZHZBM0AR1voHpECYaCtgRLIbq0eUNchGZ7wRRGAsfVMGfhpR1lsvK6VY
TscSbK0nDhPQqNErkBBPjbpOFN41y1HRe5AonNocPUuOkFxl9WdbR1mMoxCL
PR931L71zJuKIabXkS4F7JLkZ/WTWLe2U1yl0Xq0JOfqW9fAwLB1LH1nH9wc
tbQiZ694zwImAOFg32Ibzz2HDwkHuBqjVhHsr9y3P+wg+cT6NxxN/D95N9LV
VauCgH3dOe4rPDJQBBk2hsH3uevf2ieIuqQebaKosdo1wcTcX705E6HPSy/f
AUSlhDGPpDeD4zlU733bqSYrH2ggVp3kkzDgqPY6g4znGhwshAXuxzK2iGAU
nBKPQ+T0dKJGihyjeTROfJBdk3/18Sje4jY5qY/slfdSlMRnm6eT1Y7NVXHT
Me4toojtAPjyKDANzsbhYJ8dJr95zqvJ0XMcn4qAO/XGXdP4Vm/vy47Cbe42
dHVubT1i0YivCs6GJP56JOjkIkop7pDR3Ii+EtXmEW4cyW5VK3AsXI/QGVMr
IkcuKoNF6WqQvohZuM+hw7gdlFKKRDcw19QqTMZoLxtTJ4EuuOqc0ldha2TM
T9LVjGWqDsWNYj/cVyXMvre8cGxjCakLS/2Ty43hR2rI4bwxHOyj5UTkZxFH
vXDsAq8g/oLBDYEC98TmU5mTtsfITaPixJLEzakWjm+rR2nHFU3H1S5V7kGy
Rz+vQJo18SNDMDjwje4mVgPZi0pPvQbpsO9aPL5auOKUfMvUHvecFlZsQTDS
5M2bZ/LDIqoExO5XvYCP9s+Fs04mdyoYqfy6EDJ6QdGAAQVWoKRkBYphngi4
zokTukOoGkBDC3KmBpXYmDPNboJCty9qWOfu1zU0vt4nC29Nk6W9EM9273+v
DyVsQryItzUwlg891sPMAcHiKafvmPjxOpLZz4YHsbzPjGdZG6s5LNGgHu46
GcwRu19u6szKomMiYNJnJalUjyjATY/8huR1IWphAlHP0x4MbInrjhzn1YF+
0RLSvgmUO/kRidHwr98uPpzTbBV0xrYrPe8tWfHRRWEdwfwahbM9Ni5F6tqT
pZHwZ8oz+bX5p2O+WGf5hLPaZ22Xy8Gn1KMZKQj2LQtiWHKqKERxHqMMEfkw
O4xUgKV5LwFMB0tkwsJFvo1PNFQ3wH6grdnt+Ra7Z7zF3sfGxBF/D2PCGh2P
+siCap5BNuwiEERkyK3rgLnAkOBaFK+vU/IDrhV6+yTlqhPivFPYeHA/j9iM
HZlEHyPlFjXSQV4C52D8rfRvtZYAHWF/UUPFAqYce/8Wd6yV4VAnfnCjECrx
6eoqSo6Y8dsBlSUFGVz/eGfrybiZkV4KbRw3W4cJnkD+9xrQw7FWwVqU+HjA
uyrz91P4RMxhwv+17MUO4ccUICEcUAKR9juS2l1Ky1m/iFDS8Wb+J9bbCID6
uUiEK6t+PK/6B0dv296+5qXc18Wh7j16mSBK8UZU8Mc351EbK2Qc72nnMLWW
++dT2Yd5Tp2ZcS+ZvrT5MQCJqFHAwtMTiGP7bzJ63+Nt/qLQYtmmJ6jRKRbu
ZhzJu5IOXMvSYNieBdoDWN5eH7Mcw5snCuFQJsBRg7HRk/ZWjSGoejECKE3E
J/pqR0AnQbFy59428r8Ew0sm9WDa316sFcHRSwylbjoFvH5fpWto0Cgsgx9j
D6j/cyZWTVdbISc1tf2ZoJEIkueRL5BdXDS8Cp/0NeXA8Jj7ansop8wyj+HX
eMYRx73VfKRyuKvcnfqgdV3MTo0jwoDZcTexu66pC/fpUFUAqnDXqdoLLi6H
byPEjZ7FqBuQFQBMiJ2thq1LI26kZ1axRsAYmPbQXhQg/VOhOlFZPAtOyS4c
ImPEv5t0YwR+COIdk0pHVAD66wCtVeEBum8bpsHBbW0uwQPmuza/DlKkYzQ0
u6w/OGhnR4VLYm2JHGUU5atnDRvnjwTv/OSDQ62WaEK/WRu3zjATWZlt/JOU
TUZt6Tiss11+aWJ/+9r8w3nyK3AAQ9c5WwnShenZk99ZqokDah5pild0gUiB
XnWr97Gty4A4lVRRoCFOX0vxi7/VV/mQYQy0DtTKINTG0/zb7A4IqbHywj5G
JjgfTeNFap/OG5nOIuzFpyU2gDHTUN124wX5U0qO2CIFa/Ki2T27AS2bNTEi
vNJheqoIf0BjfROBWEtxhBrOUK2dqwxhW8Zh6e+VNY1jRA6QEE9gcmZoYi+a
e1M+lz1VkLd8wyNex/x8MlynjG0vzF/elSmMah/Q5RFwFA2Fmxs0l+rwr/SL
6BMiCfa/j9zqOdMs0Mv/vQJmLta0KLtolOyCdKd1CgGVt0BAKnKId3CLeaFd
BYAGG86zPXFGmgaezcPuyfQFM0v9bkjzQTXfcFknQKFO8YVw/6SY7tAE7SQ/
zPNsu++NJZqFS/lk9aBU0yzfXuYqm4n8OSqRXhjnEKc5C28bOtpbbH1TfQOr
UTlDJH+NzAbKMPzDYjDKXDoex6MnTONCYZ1ZXZJpheXcDE9amaKAcVmUe/2Y
LgVsnKxWuRMoIbpXmYZTsd0GQZV2ICliJ/Y3zfVupga7+zB6EF2Z79gmz8Zv
nGQ0c4jXjxKZ8ziM+5XfOnF/pwnh36xfH48U2mA3HaJpthfW++XnZsuaQnzW
YYXbMILTX+/p0fOBTfbsC3NsDsqeMJihjTpbhtDUnnRsE8HEbZMA07AfthlI
JOpfqo0kd7texL4hrYiW3WPhOVoen/6wPjryQueNXZ0yd4ZbvWwxYh5X0ScS
yzvw53QMlHQgNCKBrTiGQuXd6nhK71HyoVb98YVtbaPAxgs8DWnG+e2D+gBf
8q9lqFhEai6j653sfHRvQ5mJsiahTMLiQgizoXtaANDVUZsPMH/k8fKIJX4O
ivGSrF+RErT8S+Xd2mawtNkV4LAgQ+xmtJ1usfxBAYtJj0mRfOnSAIG9V6eD
bMIJXElMQqxkriBfXTWXquhYJFNOnz2yUNvzbL9sPSgiWw2xUSVAif9mVA4p
UfdWGLbJDihIjqYtywilj6JrYqNw9eKY950zpV/3i7lyKg4vIneHSR4KnjKG
CvEZLoQhG+4UTxZmts8glhySGQlcOINij7l3i1RCo6Ax7J2j+BYZeI7q2WOb
zmLsiIomg8kirwi0TN9pCP91hNQ6VnsTnjOydufC8C0IRvo0ZGZH5pqwnMWh
MT3BmdCh++AcoMNnx/L25SeCHX0vDKNR2UgN1ygwejfdhTFL6WmDGOn8f/Vq
k+wO+LoWhtXhjHk4Uo4Uuq4CLhnWSCWMHmyf+xiHHM9A1Ki8Zeetr50sX5WW
MVAQ14w6H01jOnBAP0yv0nbHWJ9R+9CrbgB8M+p4WfvlynT0QlMIerm4YNyE
Kf0T3BWp1Uuzp1cFAw4DXtzojq9EzQMWVQq8CWpHNgWudzG6yMvu3piTsiYj
qkVm39PdpcFrkd1cW24a9/oTMkHlfalqOeXgN6JAdB3lxf0r8Pj1otJ1jyTj
Dd3u+suxdKJVUSA7+d6OwY7DR3FG+ujuM2sdbILQDcdIDjWiU8wZOrKvxtGT
96cMov0QGmHOD5ML38iUjrQiSQjlkbVB6pLWlEqKYvBHCEJ90wR7cCiHt0b1
X1yOO3cskfmkEqvOHonbMiUnvyY4zjY2TYhCj2P45y4aRGkQMbqVsmzv8WIp
fbZMth0Q13635/ovKmoWN57xj0XfZlXFyX7nWLBrjQRR3elLmczfFAsgwdtt
OkaDbtltsRo0/TuYt0W8Hequ1negiuAkCVU2HFWzyAndCkZ4hzAsjb1Ty4YZ
kB1MBRqX45RocQ/VjL3JDotrju6fOms/1nzWTMlNiLumXyOVs5XLR9HFHKUz
yE0W08yUB1zsYH1yKZZ55/0O3YE4CCwwAiU0W+skPamcSEr3AbBA45aegKeH
4E3ygDuNtzv/KW743BJO9+WEpbysHEmR4nd8J61mzQbIcErlWfBnBI6CjIi/
ib1UmfddmSX8ObK10KvWp9t+dTjdv/pG3BSnaWkqIJhy5rfe2FGdlnVHP1NV
MrNgr+2/DvgHvC+MuorWCvRg9Cgdx8ytJfJrYowHuUMq//UbCFIlQfB2YHDv
Pr+znIQnI0kCR39mykFFyV2E5P5LhYWNctxmBwOKCuD7ZhLObbuZ3Zkrr3fZ
XxUoDOxkjF6F9U4nw1c/sZoZxk2g4s0Qhc8Jeb/GuZ1fWcFItCu0d1+MpQX5
J85ixP25lMDjz+tQ1wQF03VffMWNf3ZZMWpTiTwJu/dl8tVYTRQIylXP01go
GSK1IV5p9gcIUVse8hCkHNsDLASMYvWLUXyz4xlLSmkyMUl/4TVdF3syT9eT
8C3VbBOPBBb8EMGvFR1vInf8PXCV7wPCVv3WtOgG88L6Bi4JY3zblZS+2gmO
hbJF5UKIUC9a152lPL33E5Ywa4Ti5B5r1cdOl6lkmt49N1GXVXwYoz8EdQLB
SjTivtzPzVUSaGIJUSqqn4A4niCvGtYtlnHRVzpoZTvo67zW8sgvOivbKQYd
ScD94NFUJAk76R5y7/ZlvX3eAqZLPorm54qrG1wjPwCko8faEhRP0XTMOBu5
X3t1qgn7JH3CmLplT7cjHz0VuQZIuxVEEPFOayvxBH+5x6ptRGyxI2+8UuUp
MEClj4s2yvj2eSnkyU5jxwgGw1G1dSrBLihLxU6DnZF3VtfhjrEN05zbmalY
c7vi0GimGtz5gSiQy1bf/3gXkyKjQyGf7g0hLq2OBKloM6mYviyxdSkiBVwv
9yu0bOCX3eVaOqy6ZIcjKmHECpvDwnV81Dxkzqx2ap4gB2g6AE+jTfKXY5ny
6t3C7sbm4zeAwJQ1QgHJa75mGdG+lvZaBsjXHMRWVi3P0qkVM6G8hCaBhglT
6VkYzVao1duCiajlwK2tLkDAagf7ghF88us8hiK6vyitggwAsZcvmsR2bicj
gicgcBc5bIaPsDIioS00okFxjOVnwOQErEA4ER/wXDxH3Kou7wO7XOMqDgTg
sjFJJ7ohpq0qs47CCmeHrpXdE6mv+0Klx7pXMjTpbU6LgB5x2DmivpTEGi7y
FtbLiHwpvzC+FNInYFX5/uzbzC1NpCCayOSlMobWOoW1pSAGLt7Gj4zJHW1m
lms19tqsSCZbYg3EI9TvFaouE6zLItDLexrv/2/uwt1jtn3gtluu4eYqXPzP
+7uTEocil66fdNx8Evi0iWCGQQvZyCndUoREKoBgSFkWu09x0/f6THL6+AZm
xXZOylMh7Qh0elmqH21KF3qHVDkWnmcvUQqmgDhyplz7jVIMLSjYlRt2rldT
BJ5EeoH9ulJ8enodPFIGGc7yTZzXzxErk6bo1RPGBPx6lTnNByzenV1cc+h4
IdFX8zqDhyYlR9ZMxJogDHBToi4gIPyzV1HkrXID5LqdyimcS6luxGVJX7Ca
wDqzDQnm3n8rbo9zPbArMK9P7as4AFtvi24lvrxeSxT4ghri5WsY5BOgP8Eq
u57qJRQvmlTUCP1sWgAo4zQzRXhT+/fJ60lqU6HMFU/7swkFYEpUc+EqUvpk
aJy9/Yb6ZjTP2c2qbzUxdg1iJQZs4+i/B4YOdMQh1TNg3eNcw56xaxY8JvF3
3Io1H/ELGnyjfjxRFa+I4MWYcsCjvaM1CTQc5pz/bc6nHt4QEvDxdPdJd3SY
Skj2MBOwF6GLaNC/HSXBe3M49TWvEsX3FMQOBpHNXtKxOpOM+bEnwyBbDdNx
m5ioLrsPHeWFNklFlwvwOh0W2nz1UM+/XNiFkIlT08WHDLkbxa5esTh/NGKg
VF3kgcrwXv4BBGR1hHFRsh9L5czr8LyQprdfpHeFC1LiDYsUkXT62MbPTeO+
vFJ/PuKXQU0KaFpYcQrcUr6wJ3kyvR2pJNH1mlItvEsYv/iA9kkg4KxNtaZC
up3Tv9tf4p/W57yHXVYGcqybz2HymkVt8JlNb69BsS9fjesrB5EML421+XWz
H4ghj+ZkhuEG07Cl+y+gJk8SsfZXUJJ+uH/yWvnYNSNJ6kUf3MulB3fFw38M
xK0SYQM5jOBD4jvRotuTSgyQ4Py6UAjn5I8/rxLP/atLoA1mZPSg0AxIoAa+
qt6nzgynn7x60skkB3y5Q10TzLG9nnk3sZgpIDHFotosUqgrB3pgoPnGyHfu
4svCtwmI61quZgCHpqUKzM4qz312W3Xa/QpW8wWVCT3wTAxalqFnV0VXd7YQ
Rzg2vBDdkWUHJLPsnF6f4sMKyYavkx+YCJ26cHTQf+yTfnsXh5gEy2swFRr/
A/nDvYr+YG+f31O7jW4Gtr1kGHUSjPCHnNuW8UtsvpVql8aNWH7QK6xud8dX
UqfwPmDeFtdeD7Gy4sNWfwvvVsEPex3BpGU0r/nUk4Xvq/+KYiXYhhddJQG7
znlOo/cCPsGTwIisFpGHOrPUlPK8Eo2c5VbShSrDHAhIpPUUQzmKb81NFEfj
4+gpQeHjZlT74n/jiFH9kdHja8cm7jJphUayH9JIc9kBOb1ihwACMQ0V6ib8
iBjWXHM60khbRmXuBmBJpgny28bsmP4V5c9JAQi8WUpP6UG4vN4LrsB4xU71
yjIGYaRvw5+B1a0PFwEaGvNb42ty0gJ4zYHrXqWdH16wIfTO7vMuqi4t/LPk
RobBc/gKkouoQk+qXkzyidXChMIzlOMZlwW8kYFBZlrwpizRgm+rYFyn2FtE
Xvth5eQt4AlPUxZm1mjCJhX66hJ6QqVebeZVnTVm0YpBhfjWGDfw/qRti27S
DJiACSm2r8RDU6JgA6R1FP9eXVsOYia1sd3NC29dqdioJzEgcUaGsHEIFcax
ldxHVwptvOoyzBsFt7Ei4BYV8i1E

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Kttctzi5aPKQ6vg9w+1g45z6Da0UaxXtt50QPmQzmLiVao+5Qg/yS2eSRK3c1uFoxS+G6ngDcAKHm0LGGibx4soakCOjaaRTqJmqblCXBo4qigRRJU5sOpNJWGKfxZC9LZLfFjqN04HCQ8ah5FN3P2yNU1iObRgi2dEkx758LbIsGmsSUmn36d6MTHQGWCnH/AC+2pgOY84Iul0q5eg7DNO6RSxNOih+2JmnF8szbMM93OCd6DNpiddU67ZKuD+HHtVdrZMke7QawemkMeOkYd+l/J82ScFe0w82oy3lXlwEGjRpY32+gvxfwinCXu5Y0z8Du3arIcbL1A7sCsK5d4NbS/UBqd5+feTWfvoUQUkiUEUW3VOgKHIAdnKyCqnuZcvvTpxh6TM7vxFv/zc+hDrcKOtjKkQzjK1eSUQhWkjbn3Y+aG5OE9B35AX5/CPHXGh5UtztU8vbZTm6kcl7P0sqD+ynBHP6SU0l8XoFPLq1cahRKiBE+gk/cgT2nZMWfENJGTr8y//am5EUYdEsoaT3Spqwx/ndP/dZvDhLG3t59pyOppro85pE7ny5uKU2UrczYYQZBIf8eDsaS26PuLQlsg9GsgHC79l9qlFuyF558QtbcMStMibJwGTcOLPYrNhsL7C5uo1tw3xO4EqAyP5Da3tQmPZyVgCd8qZbq3RxN06Y18deiisyuAQFd9agLf+G0pFvOU9dofOc47tSiluc0NKOnEyziLOxwhOCVXgYPIVJEQlyJxR5Qlx02q67+ZjQhhlUVxEboIWzJ9PXicGaEbFwzZOQaNA5EwBhimw83FUO1L1CLEAV9x0AKXBL+ud90KaNE9sftYuRxRXCHFX7P8fMxhhPQhktTCG3MlS0VOWMzEReUbSMoqNk0Liw2imTWFcFfqzN0i4RF1UU2/z43rLzyZupNC0gP+5NIHTPbto8LWFzjtuwhY++CQ2pMWkLpO0A96Gw+H2kqoVhvBYZkTMALB6TBIAxroLO7ba6MkSs+om4i8huEib+zRVy"
`endif