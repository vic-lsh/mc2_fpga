// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dAO8bYl6D/Cz0SaIs4jhZyGlJ6/ZP81/to7q7U/Bd/pkdLHzkbLsa6zQSUU7
s5HFM/iZk08SqcDpumb1dL2FPwpKw8062k6GenZt58DRe7X4g6mwag3Gkafu
jOj+oF9U43jsQth4/crd3xfm8GAqDuWidPzygL57bWvBXvmnDDU5f3mw0W+t
AsS0ebKXJC2MumNuhJJDIxBCo62Ka8uo1gReKuJuwi/O1o9GN0cZLje/nAIY
DhqoPBjiWORev5kXOi60cgGVCJBIyhgc9cmnbrz8v2zhpZXO3HRjKALAdBVo
hbFLh2chKFVoZ0GJFX4jbN+nxtbTTPy8xPSmLXICyw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Nc0efHQ6XSl93G/ofr2kJ7k2PCH4mazcE03Ni4H3bU2P8/WS3z8LwkguHHF6
wC5Oik/wSlMCRrkAuYcQCJR2nsvXzfkdfreP7D278AXev/5sjKGdm8ERO+iu
5WWnjGr7OAlkjmdJPdFdxzTSQz9vj4sg41K0byC0hvGs9/U4P3iaJA1oRan/
gTVNjKQhOXCGz7PFj5qIw36wgli7j7+xxYSlGHUaSTyoJzxEFFqjh8b7PV/o
NhEPB3NZ5I1EEnhn7fVCzMsSsi7xtWMaWYcT00y4V6R5PGT+zsKkphZ39d9F
3P5jXK2qxRejJfTmnMdUr9U9pSshj8rCvpJNHwTWGQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BZK6pf5XDfJ5GV4L1J4JzY2lpiRkiFYyly87LT8Y1w+izpaerFqC937CWjew
Le1P5osbFz4XrOI0Ork2WL9S7aAF0MsyQl8q8UdBhmHIUZtAIr1vty7QEh81
RrmK/WNJFg9mgi7/uKz+IK4w0XGYfqxzEEIdxzs7ItyUjuXwpcXsM0Q5DymM
6LWWnxPgH4ZAXCrAnrPTF+gpAVcI9PZzwAKKKWBF4IX18KYOys+lV7WQMaIK
zoAfFOzh1NHfbth9XZwcBXtP3nssaCd3oiuyd5BypopUVu5j0duRgFmaRbcT
fRfhvQNycuGXPA2y5a/ZLkdt2pxYiRowxZP9TbzS7A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QyNMd2sRHaOOZCLYoM/XeAODTrDJUwt2RhzIYzpJnq4+wt8taJDlfBiIEskf
9CbmACEcu1RkxbrBYm07xtPPmCO4Ntbv15hWXWSLMMVEJQmmvLTFAKw+gRSZ
E0VkAF5NtBpycJQuTtows3rdOq2DASsB8XXJAFDESOIDisBUiCaS2YH+75Rk
ap91IPe+GREJ3Al8e5+rNGgtBTozYfo0yOflZlP12a6Y7yqvqorWyfIFlwrw
A/S+3ZQ2Fv3d5MsmWUGfyatCzMMsqTat0Dcu7Guu6MTQ2BJXJs9W3QTR9M0M
KB383et1h44rSLZbBJvbxjRjoT3iJI6fF3YvJga71Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZA4PJR0KeL+URRDJhUxs7s1WVcsrRjWZQfB+gryvH2Bc4KjIzBtvtukCMFTm
MpDO68o3uHTtIljY+IuJI8eaXnEq9ZuJ/TWRCBaIj8oxQuRAX9oMuukX9o/P
JrT1UgPZEAs7zi+htEIebgDKpbd8YMfSfom5F2kQUfCulYDGK9c=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
lZIC/4cWcc6QzB7RZtHWjFY7tuoEJhrE0SUG9aDyELL3jlA+sMDEYI28rW8I
1iOtrJytJHGUw5giw5viHPF/bE2YspAU41Oxr8ujhizFUeLwhAyQ/DqB391q
q+v7j+TA+nxXnBImQfN20s+Bod5T/H+CLFh/cBDoX1kDLjpu2k/TvzDElUUd
80C8u4hLI4EuEFa+RD2RB1f8smuDeHeG1QrTLAAyHqlG2ShQXQ2IY31tEYWo
lS2LxA/a2N6/558M7sB7W7gHtgKj1RdP4kKIDyIkoMXsBz5bIhehnN7eK027
jlzwsL0+eBbe/2yh+emm5p3OTpebZ5ExAIGHnKuPVMC2KBxoHVYDqu0IglNl
TKwEnmELMSSmoRzbEY5guW0Au/L5IpUOou2UcAwPqbRdeD+D0X1e7VhigWV6
gznCEITijae6b/de1C7pPlVcPwVBRW5uzZjXe2qUh24IBuHSMTJIxDpR9HT6
xgHfkPPc+fj9cb4rT1RCMBpzaK/TNdXx


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IwR3Fh4JYpAjwc2KtNK3KkBlN7VispzJoJAvu9TXcj2xvpGQH3ZpZhGssI05
uxwOWYeeQd++KY8rUlV3avoAFQSg4/JZS+hXTf2xEFzoUFa6779ONzPv3RwB
SSYLw/5AA9n38+kK01lbPpkN+rWmENsfxQLjVCRwf2Oy9pC1o7I=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Cq3f9GU07rTMfssPR8fvt1q9wfNViMUyHieRoNDEKa4FCJpeBeyysNoXrxAv
zOOA4TTau3vHJPrqgD7Cl2XVhM0d/mXKp3KcprzhW8LPRUd+al0HAKego9kX
7oYW0jMz1YLTXc4di2ZYsueEC6VAj53nfTTGvkG8c+wPTp/eu54=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 475120)
`pragma protect data_block
B8aB1ESfnBeOembLRJ8zLpCbqlG3YwNbS91KGMOAuOWUP3DWx/xkxAgk/NC9
gOPftloIiYfKlhk+6Ttv8++CBzYbmZ7AZvh0hxNOpEn6/908FtXFhlvA2Tkv
KmN0m6EYR4mQmTto5jMtGGFHcNwIdp8qjBsNpt/mVxskTNZi45Dlh+odP4e0
rvF0xIpC+IPsw8joWTZuo72g8ajpDg5QbGJyM/0X7Cip1LZIIzlmz1nHbqqF
huVM2KBQFQgqyUnMvgKslRQPMxO9HKmQBuMUsLaQqRdZ5P9ZEodA7ApQmEw/
UCLQPmpKWJ+zm8c2fIGqMZ6tsH3xjdLfMwfuU3QFE8wOeEz9wQHx+o/9rjSt
V8TPA46kGTOQdCNVDy6c2u6Duq0F5GCrje0UoRphT8niKCkMyFdIN62pK4qa
68tWt4bOgFA6/zCPp8jXs7B17oq/M3PThUKN9EKBGTgh4So63NpPSWQj4Gz5
KYh/hFENhpPqOpWy+OZxNcFaS46yo6AgfbRqE3110Czrx7vZoPhay0JLRi4f
Zi7hR02JgHcPxa35dkv76PV7nT803INFAYo/tB/ZamhXHKL4m/rYSzzR5Wc0
FmE1AeFmqy7zc8OQPiS6XaFZ4qDRUL2MfUnm7wX6Kxgc0YS2sCgK7SqMMx/I
+F/bZyP9uRq0kK+kZh+bIMe50zdyebEhPF3UN+IiRGE/N6NVkQ0xjUSSYXW6
cieNAD0n4QL32KBZKkm0j6wKiJYRFh9Fd7UlD66keTpXIpIxnWl6b65MTYGi
zL9tkJpfcK6+Yiq68hcAVT2Q4rQOHp385vZ2Nf9+vRkjWQwglbjp53biygTw
E7hkHWRlG9QlOYI9pQnocPSaw2cfJUJ9yYmpCchuLVl+VQrDZVGDmbMs+XhA
sIngNUCD/MsMY3X9w5AyDfisVwGB+GoT2ituYX/Xwq0xWC5g8mj8w9Ix/Mp+
ybI7Tgor5nMUaJ31j/qY6Bwcu9vrvsRrqzrde5KoMF13CPU9990Jw4kUoTLD
oh64dkyKNwAaZN2M2Sbxw8dWwsesqkblbjzloPoWEJnTY72J6sAH6XD8gSAW
ZZm24e218HP8Ou9FHuR1lSxg8ChCdjDotPaSFHEudpCk9pZp/4s1Vl4fq6Zt
TZOlCyb+J3us4J1+u2L819NE40qEfPQ0soMRQE/DegcNEFTN4NapXHMO0y4E
IkKifaZMe5zGFwrJMJXpulJcX3n/w0Za47CXX+dxuPtSH3aLlM1sXzF/6CyR
rBoMm9Bs/UNgXrkCG6kJ0t1o62qA2KMrmW4Qn+7m5iHgfFyUPQ3Qee7xINIU
nf12LeHgwod3SjSOaGj8w6GIdtfEiKjXIwu5oAuQV5cqIEpVsrcPVOXaJS29
vKzuw9rfw2lOwBOSer1yAzt1K0pwcB4iOPwZ5vcj4Rh4aOjsm/1B4fvjQ7wG
GfM20PXMAngBd8FpuNdp6UjfJEc1Kt8OrjourEzZKdCJyAKSVzzG6fh2Wa1H
ys51UUkm6rRxTQgCPIF8SaJEdgVa/pNtlEB8n61wInoOSNQrp7kWAZVcx7it
V+znR5R/SaQ0VW5SeU6+QetwNt+xHzYZqqOZdldn0Iw0AbfxGPuTjAaWsAqx
9907AODtMcM4HhrgMUYA8gqtAc32Zj0RZfJJ1GCRihSq+sTxKiPVPprR7L1Q
4laK+FB9kDVGpipkfD6rh9WHJ5dweKFm4UdjB+9qYPn5VH0dXax3umoFMN1c
p3iSqVHy4c52OUIQjumhjMi9UI1VC2BdOTX3TJKPIA/VOjq3/K6Q6R0ssfVT
db6XYurjxE8Dve467+M3imzWprwGnExrvRQIAyk7uQ4yPQE9beozirgMmPWX
JrgVTgyAYIIC9knmCrjKayEAx6kmmPmsVXJZlPDGJZYNkg7QcE7aWvvQ4XXk
sG7AoMhH9SYe4zT5/PQ2lZd+AePwMN141w4YF1Ph3SdkHp+qQCRrvBSt/leu
DtjuXUXG9jlXGle+HnqRCEeqrvj05AhvM+XCSwBIE95RBcVy2EugGE2M1oKh
OUMUbo+V7jhAhWv9wmlhjBX+GIJClpMgFNKHTLV7Qpd0JUyG3J59i3Do7+la
r+6jCqh9DiUWkdKgpkiXpaYIUfQPn+Ooo5BFYwZGAcSJfyf0xKDmW873JhJI
WwcAv1SMJEMXX6RWGvaS4Rup3zt33nq7FY/DPE1yjXTfiK559wssmAtVjRlG
AfB0n4m9pMEnI6/Ad0Kh164qUK9HNeJHDduMbxj4UMVg+xRoku6R/CLfs00q
jx0wZtd28EI6y3TQT+b/lYCmJwuh1CoaDYD5IOacmsYcbXJnQ7fCmU7IBTzH
DCNh2F7NPTz2DeEtZK8h+Bxhvg2PqyJyBnjbOrHxhDJyqa0lZEOPCW/Fy/at
GJ0NDa5EkTB48hGL0rasRsRRW13ELZ7KEy9ykPa+HtbfIhtXZc9Efq/8k5UQ
KIMnJGUmdGI+sLpjrrnImZfW7Eej7LWMNmaijbPOpb/3ALjTnGPFODOxuQqx
bGpKmFXHO2XjEb4LOQ40kstVcQIYDhACcwDOyoRNnMVUOdYlb6avCguB7vDS
IDXkAieJxw5AmgkPKtjMxA3JjaiD1qS7rm/P0NNXATGM+vk5qhHPSFIkZbVx
mtMSqTrk/nT6oovjtLpEs0jm3Xnj+0CH8Ir7OMsszHuUPwY0Q5pw37weURsA
bpxf6DZdHrCdlmyczKyfXaWigmQ5xMNcV966OzBLEfhfKEgXodegJO8U1CiZ
r+TYJl/NkM2vph7Ota63rKN1t+FqqBZxyGe33npWq5VgPJm/NzD1U/7nwlZf
z/iy96vJ9g1ynnkmLpwyuY/McLq/tZh9kOaGW4e8KzVGMyN3EzsAYatuiDvD
aQZohOdF3xmQmZwhNe8DR5EcUrjemAk3vOrU+k4lgfrgOjyo2NjnlFSH3yNk
gwaYx/RKP1p3ryylDi90CfzchnKrlY2qjO9gpyyvCUV9BvJPwZtANFt86S9R
mz5vZgXo2CQ/xjyeKjUHjTkdc3ewF87FUG72NDpOvX0djH7fWBTXA2zCnwIH
nPGkM/fMVbQsdZW/cEWBy1gn1hFeLKFrlTYST5FijPN+attJ40QaQulq015N
7Uy+JBbVdmNNpKjANlMeNVuY39pDQNBGDhI4wIUoB18XGO9AX0yFUXvK5U36
NeTVntAEaUdL3wGw52D/V5xUdYaQDPZYzWFj8bt33QfyDmERgODJswVY6tGd
x63RVH6bS1ClZ0ATZpaxQzm9ps51lMaOP7gPHTn1BFfvmi0mWPFZFJICPl8A
mgKI+yry8XrKfLHiAuK4zkFUnNE1Ekfv/6uCFl+VaDFPkcFIaR4yTWYgWDzZ
DFDIplyVwP03WuZCxSv1MCQKrmU5G3Og3BOgpLnD5csK3hI/pVLgf6L/fkWz
/IN6bI2MVSoV9eVc4+HvzCl94t3+BVJe/u9uhxj2Jp1DEBSSuafs/ntqvp5A
pAfiVUuLOlx4QPaTln0MR065bAbsmB9nFAhfEiHTydEzs/sKM5UE6ypTEA7K
Jcj3WtkJxtYPYVwQQvDD8u+HUtvb4lsackx2YZOu4m5eeTDB1Oi1+UCoVtkL
jvFPfAu6D6SIqyCzZIYaTqX2+iy//BMSPNdjdJWmFo3ND11s4OL061yKTdU7
94OJOvT+PZlBTenF/GRT/cNomjMq3D4e6B8uHjDKS8p6WpK6N08jOSkyiv/c
EdLoDQft6zmGRfvJ5YrfoZ11t1mEiCoOfPdb8jnoXFkVT5+Hgu/8Sza/CqRe
8d+1ViQMRRZTaYfvb3OI0e/eKsJ3/9Jcgi4Sb+jSuFqI2Agq7rvN6yv5n7X/
H2QmvgGKZ2bAcMAsU+QPLrHRQybNe4EW5QE8sCH/d4H7P8QdaujMje1YLwPU
UeK83icBs1X4RA7Pzwki3YiKbAJTsR6oGCz45H7NwwGFQ2j5kksriy6WsThY
Sxw0cSJBwwtd58BlYzJoUvjsNuEaqjwIkF8/IlFDBsSMpzt4QEQw7/aFkDT5
l75l3JqAj+sU/ezd/3CyOpdWNa/EjJ7BMVlMsekM1/NZ2MWg6g1BNaWuU362
ddYeg6lkPW9U7+Pvzk0BhmvDmF6MjjVgSybudFdedfc5VnqorHjQJuZvoNuo
C/ZOieTGM6jjVQsExBzKyduomCZJ3UfQx5FEJDc6449TjfFBHWFn6U/7GFa5
eU+vsWS6hgBh6MPEmQU5WCiDBKsLUu2NNgb8Lje6TTrU0o/xoL2ylRvQYFxJ
oFoBETz04ppUoDufVvWbJO4G/vw1Xf8W7rkP4iEzQXEfcNL0rCNsy31HFst8
AElH8EvjMzHRk5NEYDVjG4hXO7ToaOAfkYHnHYc/haGwRMMaF5RoeNWxcBgi
MJGNf8ayPDSK9u7u16LCEQpf/r1qlATu0FND5kwX6C3Hc5xu4Wixmu6qfdNL
OhQOy6jf9yN6tPUiQtk1x5B4OfJUBSk5z9tHB5xkQaSeyGnOkh2fwnal5Lz8
cgEdycMmtE4kgcQcJHRnWGlwn+XC8HnCSMdVnXFWVqTVg8H39Byox3YNwAGK
a4171fqImdeiqvvb74e7vl36J3uWpGll/bqwuQnRZAmwcq1E1c4BCa6iwKop
FzoYqjR9JoVzTb2u1uDxigREF+Vm85kIktVC17Sn1nU3IOvcSd5xI1eO/lql
kyDZjmmyQAwuLLBFORaTfEMkcW9W0mj+vTXsDfyTohKhjeLLXu3marwfabWt
CCWT299DZP3HHTf8dlNs2gRIg3PhdpzREl+sIfBxwLARtPok67I4sI1alcX4
G/k3TlGTVkfwJHFyb9ob8NN+Z+FEk/2ehLubQ/qmTUC/E1LJJBpWcZCPirmC
rMICpnQWXgM7BxyYdQ9UVuzea6A96vev1sye/qSxIMLGYEFnmOQYgjgXJmU5
nrTVWtteROckbypgGSkQwWb6D6tcef0s8d2KwAk1ox3Hmkx7rpsM4h5xvVnA
JqZFva/ABHmuW+UKB2bMNXdTTm1XAJec+1HcvGfZEpK4eMjq6vAbRIJRHGst
ebEOK2aiZmXMjZmpVkF3c/VdwtlzWSzQ2lmPVKPZzIyF04Pf++tsRkeVf5Cl
z8oAZuM4dw1j+OZwHflRZQ+wV1x5POH3JawiWcza1eKnmSNfypSG58fT4RQC
bX0t6zKxoiHaM1iB77BUq/GU6sCabbVOay2Vd6UqaaEesoyYrwotA1lrfkbF
SdtFNDmIyz8+/E6tKAuatVsp+hdxi15pDPyaa7Os/yp5/rQchsnk7kYmdmkI
tqJzZtSAC8AZgydN3yPvp4F1WWD3A/CtbzJqtEEm5K/IJwu1J/PMxbg8/cjO
FaFUh/mHeOIpQNRH/LeTZY563eLdMgGTeU82aZhMaQmHOlwV4CcHrsVgk1xA
QwzktP0RXkr/wQLWcuI1qmXGBdYrU+dMCuUsFpXbfK6dZ2FIfAXeVtuXrVUl
7ypgjZngNdHV6xXnDmgCpRe4THTE702W+aWiu9lfP2ulpxTrfeVk94pkLYA0
oHyRaBr7bX+owR+9odmrEp+XiAeZlItbD2W85rgLAKt2zxiNTtvyAOhc9MP6
nUlulhnf8DFcG1NS9Vx1b8zv1cPOXLXVA38HL76OVlZST5G+UmBi+x5X4nRy
oqBhy7rOqfaOscb8DNIcjrenTthFUYQql3MbCkp5GhFIxT3vvvjRQZMOWxYF
1iDx6WWe4Plhah1W01/dJuAW/1u3EjmqqPrWvaJJIxHcUqyNUseXwF8wF9lL
oU1PZYbHHzXGMCoiwldlhl+nDh3ZO6O3CCtG68blfegH+HrQKeeFzbaL1Mi/
9pWCVWqmDT/h2PFrVjpAExORxhFl1prt5sNv8jfK+/VIsOEKoFCFZRm2Oj9E
cA+Qi4mN/Va6PytcItBDu3jFaKCVFYIZWp+r3AQ1saSBmJDjd1aWsGQK/4qo
Y7J7qfILBE/shaqsw7YnEp8L0lCyaJ74w4eNQuxZQGeQFQwLg9rJ2GyX3jln
w4G15knyEFn4hv19INeFhKprnRWyRsGq9swrzypIVnKZj1eRua0VjLFvqTeL
0mWBWemyrKvQm5B113lVlomFuX9Lg2yGiEgr7lYXUIQj9DRE9MK6qd/R67z0
xchUGim4FUFx9XcyHx6W9L5DlM4VnPaEsZWKM531JMQYArpmtbqQwAIQ9PS0
foLl4iSb4D4yQFAM5Byyhls1q9OxtzrJXDHJWjej2vePHM+HnC8B0nQVniyS
fsdj6svSexMahwMXPjiU1i1roUVh+rPGzUaw9L4cgNd5YGdb5cmI1D2GgPEp
BhxgxuhIlE1BQMpYlOiw1+JFfnmZC4c1ANhG9EJbZb3S9ZEU4Kp4LbriZRtG
WVy4pubLz8+eq9B39zIIH19Z3bX+1n+/iROA8qYyqQxVqW2BEl/DXsCXbI8K
XhCtbTpe/m7qkzNIzfusTi4JLv8kIb7+YEuNa6s8vXE2EVgqvblmopmUD62Z
1OwMdj3YsRpJvMLgB2IQdHFyscb33pM5+sUxZ7aZlFmma8SB6M+uYBtn3s/j
+WEC+zaeVMnv/sxtOVi8HVnypu42YoNmMqjkbsO0Is0ZGsksE54KZjv9A4C9
7Inrg787HrJlF3FiTLEXIepEj+ga21HA3uuyEgsEj6ylq71smSO1yhXvxrLl
a5TP9O+0W5O9g5jtcG7CTzD5x41qB1NTorpEwxm/EVm6gu1oGL7Z1tlr63Zt
Xhe5hLYWkQ2kFdDzB+xDcZooYqlxKKrvBHThMhWpZCBOKf4gideyzns+SJh2
g5f23xZ5qeG8Am9gPuiMVQWANQoSL5L2hLFq7mHBsPruYNxzlLEkxO9tyZT9
TE84UWpeMgPXoVdvO/C93Jitdqgn0Tp2CVtcsv9OLor7nMv+/JuOCaUfhWgG
ZFd72CRqdHpKYl8wAynIZYQ7isj4QA2BANQDpYMc9/SoZfi86qsw2uqNjchI
hDWMDM6ej5LWbeaQFvYm24IHehchqR3IWXySbiYjeYbTFgG7BjpcYPvdkC03
GzmBps/TA87Ly6Z8i5w4jr6wYQ2cSPdhd/fkreXLtzQyL6ulQho/ZJKTqr9w
ucaqhaGwhYSDis7vZB9YPERR0Dkzc6i8jVyuC9k/KPo1SGjkJ6NED2y3XyOy
2pCSrXSwVTtTUhKnqkJV8bMreu0OHQ8e/JBIjStaXuiGw8oudpkJZ3baOb8a
m2Tj3bZcuuEb6OJk6JSHG29U2QqD3ozOMxB2YSSCXsxlYaTjugrru4ZWZPCG
oGnvQI8pa5rP+elgdYJHkdEXMHCSGMatcq1znZJgCq064E5Imxg0hJEWMCp5
Q+WkmLIX6wfBdn4CME/G+7+h0m3TUmxFEWro5BX8/D9QJRFe83LFmag8afA3
LCU7MMMKfmWfGhehOXDkAGdFejcslq5tnCzRm33Ip56TS2ftU8gh+akJWTJD
wk9WURajK4D2yOcj8SI6VaFX16DmTqhalZlfQYwwnh2Fxxp5vnyKiLFMpj1z
Nbyviy5DR+pqWufTCbotznkozmLywxRDIPPHJwyI0JLxX2OxodyKX88q4V0O
cf6BRV3HQuLwgn8LdmKEt65sa5DAzqACG7IHCu8AoTHHZ1AWkmVVtfzgGhQ+
Rwsvc6F4BRJvZFpcLqtLQIb0mwbbREfTHhSGMfo9SySrSfLLpWqoo2RjsdQn
sDT8qZHn7Y2VX/oF/VOU/yURzvFJJqa0d7KRu8tXwRyrjabJ0kAXLiJ8V3zu
hgV2ghwXjw7BtlmUdRs1CNRFH3Sm7u8fhGJBvSxiD/J9dL7BIEls+7TaejAm
FLQJMb4hTc5RWAOTVTw4qMg/y4XDkziqN/y7IQVeOXWvnqnQzUV/jj9iv1u+
aqFIPIaNgjliRm5CP4nthyA3kbbts/lKDznuobBrNRiKrcPdSc9zi2pcA8PF
ZUzwnEZPIGygTaEG2yo1+5+kOkT1qpM9SnUXqe0pBUXbFFTLZ7K8/aHWb/8d
P7JjEWPFZVjiP7YdIonA6ozXVqxO4oPu8tV5zu3/wGPYCP8gel6+B5KstLMo
nvQnKKR1UzTHT4E3mqfbRYqcpmrA7oOPG7ybFOeSEMdPK2cKGRVSbQI7CfBG
NeXb7vhIU9txSAhVJLY2BWP7G6Y4LRrmTjlEiLwmbG21xyZJDau47f6QeB5R
ylk2lUMyCDAt+pvhmZ7QltCv+U4D709Qk2JApEU5Awl3yDQdYKp+uaOPLoEI
6NuTa+AgDOHPPRiHLa+dqURGb8tw08dVfHJgG0lZNTeNCdj+0vyg2so8tP2o
NvcO2E2iWKr0tYKVAmZv5ehHn7fCaa4Ub3batgTFvmbVI/j3EIgNJa5xct8W
BAA1i1jlMrxtPCfNAxtqmsDEtZF3GJg9RD7sdq3b1DOJwPFdohJQeDKYWJB1
J5WfZN5iq4YfqLigDALGJ/+3/LISbKCdHu4qSJcsCSWBGYnFSOYqGMwzIE3o
8S5njx4szxNqpo/mISAaAKtLi+oj6A5k3wj6Mru2EmFXVCfticuTl+ombSRL
XU0EFtRXs/XXD9UuFLlkNhm9VRKsAxFhJBz8Lwq+BZ4ENgd/HP+u2Kc5OhmL
0ACNXLeR64pr1Wxrbd1Nf24SwiKKTFbN5CYyvPSEX/8EF8wp9bXdLpvp/2ZW
BongCF3WGAh8DdpoLZJGizYGgW12P4/9rn98ydvn3oXRbWFccD3gM5NUI/v5
NDLhYGCESE2Q+sM9IqGWmLUm54JjElN1htTQkkzgfMLyjKCTaU4U17W+NbaP
74iFa/3tpP17LKLNn/mLSajCxRwZJHkhuLTeiruCXhHWcM5UWQWXbIcbxoET
07+Rsm+fUe9Ch7v8TK4exy3rVAixCULnI0hT5VgcDS+DoHLUeGJNeU0hc8y6
xE44z+BSZ/rEEvV5+efLY+ecpG7QneVqj64atGUPMePx7UvmLEXMys3yU/V+
0Wj4kjXGoPrzKDZRsUi3gh6k/DsLNOTj+clna9R/NgilQzQ3atMO/RY9Ra6z
St2xICl7NvmVvyBGDSIzwGCwMixL+Zw8Dn6jBMd+38ThX6EDVp3+19/VPkjZ
IpVt10xwJ0WqIub8zbiUEAE0KX4QIq36YTdUdhHSqWAvG3sdB4+5pANnakm7
z2CytU0ou/6ETsgfAt0x9t25umSpIQUw8r+R/CcZ3ycPwCwd8R1APcISqsnG
ChwYs/Ep00H5CKTIvbZX5SvhKDD13ZvW5sf2VfiP9T/Gzdmkefp+bYdgPEkb
rJhdeURD3Et2dp+LEHsKoTnblUYa5v7DWQC8d15kpUdKZsrniT7SJgav6TVc
aAsj5huTcKzzBYo2s1eEgJX1QNArUM6isrmXHzkAfDWVM312BzvNXiwU3kXE
J7y+dVId+FDhnjiaETlunc+0viQ9Swxgic978K1C0BSXBxMnEYZ18tv2VqDz
eNT7QB9W7qc4qq7saX0VUzrbMz7OA1naSB81iqGYI+eDoRcOc0X7COHrpM6N
BjC+t3NRL0iAUXmVGu3l2UzYLBoPLcTvPsAvXnZiDQYF5GbpuDkGbs0PUdKI
AJ1cxVv0BkuAopQOOxbXjC33WeciK/S2fxub8wSFQXLa/5B4h7+mT9YNjgx0
/H9HpH3zbDVP8d95UlrN/riXKb/7oLjJTNw+QuCfuu+bx58IqBDAoBBOemWs
pLEDNseqELVtloNUQtM76V76G4jefJy9Qw3wxP/NCpy/Rwimkj72ctXQIuS2
0e4CmlUKrg/8Q10dyXyM0sxRl0qzH7i7vbxt45QpoWEuFcBU50gwhWUp3RF1
clFUT9nJryCD9L6E0YsqzbYBy5Cclgg2isJ3Im0I9pQn7scLneo3E2EGsUPk
7MVHQ8fBX/C9mRA20IUYWnfb3DhifMnwVx2925ODYTcNcRWiRZHupv/bLYzK
c/N62W6QoGL83cdMaVfj7p4++EmX1EKxJU15pn7Pdt5bLG40AcH21YJqAFFI
ueuJ2wVy6pdECvzCUOHI+peUSgwQzN2rnuOavu4WegoWHKHeLUBLhIH1BJPV
L35y6PDTZEOzhNWdArhOJjV0KKFdAnALMpm9df0Y3mEhWF5wPQx/KRglDUOK
d8GKMtqH1+hJP1pvsdfOoebf9WojKSxZlP49NVQRlUqJOCRUzZAHni6WegD4
IIgnikkh1r6Ht3CgeQdJuhtiSTr+vA1Xjbs/LeElRd9bta8v2f5g7lhXb262
QcnT5ZP2Ip8CcxqelA2CYOZusWZYqe9ZGazws8RikCo23+gyuvRf7qGG5Bsm
ze36zooUMlCI3pbwWvBuGZSkZTmPGLVOG+HZY61W6NNaaheShxDJSvUxmqMM
ygst+3BFr0eskbhg8UDRJenVXHB+c/9Fz9nVFnwoa6jXLQ3mNO6+gy/tz9bQ
2IWc5YHOV7Ucgl+GrrNJWzt8G8Nf/f3QHwic9ORIaKLoDd91QdkSKL2MpIuL
XZ5YYpkVeMxaGGxEbDe9MjnJNSVggH1xG3C1AIsBi66tlOw1mre8GOSB6pXq
RmRJPrkcxRWgyx9OsnN10Hm6ZoH+Tm1i7NbSSP7nBNAe504gUIiqVqFJstl3
PeSVx3L7qdO2RbKTnpiCIizP5JIh8ZFtgC8Uno8po6IJM8ivbRJ1wxrHzndw
qhzpA7M+QaPpewwLjVHgfVGuHnQGu8d5M27JTPbZ2Iy3EPvGJLAr6o81LCSK
YBSVBQKZk9ABfwZbplDauwM0uMWQUuWaIDJ3gpftlQ8/PEB6fuXskoHHwUxV
zn5HAWV/IIrc4CTbBNcTfHTGWMpzKv0N41qxWYa/g2OBsGBEKsx3PzT1nxiI
cniYdKIwnFZNQMBfy9eWV3OeF7kqNozfSh0YnxLITYUHN/oNqwEK6Vayl/od
EhHpx71CqfYFMUlTQkPXlOSilrzDgN+VT4IQTILfM8u0O1VASnw6u4cjo90o
9BfMctcqkujfuD1LuQ7CT42Vdhm9U97wu15x2uszJnoMAcuMj4BvXOuwg/CV
r7SF1+cJb5SD83a9P/wccM0Dfaaq6xE+akJQNG4FHhm0kY9yd5ubWT+NMiEj
ljdSDmMalI2Ais7QqMS5AXYieYy/q0KyQs2darPu4dV+6xDKTQFLQHVp+g7K
PEY5PVQjSPw5jHHPTm77JJHHMGf0NLm1cG4uCXgpw7eIpZkE7hxR1lH+a8LO
ecLEPOhQTjghJJjmGihs0lb7fYpzAAZBbDXAiX8GQXhLjRkVnDthlrAiSekR
F9vOWDzpyhVEc+wS71k//pKivgE4rWuWThxBVHNg/6IbVfhxlseigBzNp1ie
+bpBAYiFi18RYO0X5eraGq4L+XB+BUavMzONyUjEkrCCeTVrfwkh91YcD2RH
3K14CeBFga8O6YiXGSnHEfvryAgjAluheGkfZW5MBzAb79VVuryvA4kZd6l+
9NGlueha5nPKoAKoLol8HVNbbyHonhjl2AtubAKiK9pDbxHO1e3TzP/uYlco
D03DPOPePyzljuuoHmnaklVwuxlNYgbMckPZx7s8enTBYUAdZjqQSdUCNIuE
UPrQ5NhZauiTZSM4z5ZgKpuwuBgdKJfbtZvX7vIxYneN/3HpnOn9S9KBIZ3R
btc1WTckPDRFDuNyABpJJSRq+431KuyqLYQGfCCsPf4b9/08voRbPP+Q2PRV
YwGN2j5jVWRJJTs4BbJHB50CE5SUDtls4bTwEFpx+qo6B1SMhwjU3Db2K+tb
IjfEYSi4ktdn5E5XwhadgwW5OHI2w7ouQd76m6pc323lThENA5CNDB3D7LFi
VZVZp48+q/AzBjJzXX/Ryaq+hF6Y/G4lzMaHHDzI54g1P3KYpsGagS2csrkX
2OHvHQS/xkwCqV4Rx/GJq2F2CuaSS3ulMI4P1ELPeWGUHgxJX9CWkYLpqQSq
2wfvJ+JJ8z5vw0GapTpe3Qc/YfTD52m5TTZ/OXxHpZGOA8XoJLf3xd+m7+7J
DpRVNKccnB8ruMdPOGVmNrL6yudeJ+Olc/IqsFO5sk+z0UIFJJ1VwTFbv5ec
WJj9o8bmbh83e/ED/hj/uHkYtBJuFtpf0MMT05ScwI6bcooq78pgieG0FYzC
TGW+eVYmZc23PHZ7v/icVErwS3rSL0uEf9N0j5uvB8eWkEcDMaVA+tH+ZBNb
gfm9BzMzl+KGiLBX66jWNL+mbWaW42loX0Ud1vnErOyVFrCqZDHfceWe6hso
WrdOnv4L7oWzoyM1K5MPyW7UkXi9AeNSOAUY5TSaw2VeN29F8O8MN/FwgmlD
UWw/26XnsvrJryvQdidFkjDWnwk+KbBfzDifj4c5c2127cSCKV6I2i8fcJDs
s9Ebxn8bMODKkAkJ5Fyy1jzI0H4HsRE82cyq4dIRA0iOsm7oYHlnaxQkv8th
MHHcLtX2bZ9ztWnKVO48FkjntuhzZsvigg3cp08Y5hHpklq7xwcVhrBbqEhi
9BAwSPPHTHOofLEHi2PDmmEeHyqKBLLkZu49kVoAKj7duROjI3iymS+/FEMr
YPC6ggPO8zTiKlgbVnPSGh0orz00CXWe1q70RXLJwFnpHVxTArNauNHmWK+V
yDnmHHT/yq1mrNcqrGmEAgA16w/LzXh+r066qXUNoAZ3f+5P5hOy14/N4gdl
pnTaGU9nYVXwvnh6AwhVpLw3WcRI2k2QtVusxoxahFmWxqlxqfq4zWIJZvsF
+5yCfiIEDzN/eOUiCYYbx6OD/pyxmlGZPvNzZy4hH3J+Vwcjyk7S9/zUfZiF
mTyqRzj4Wwb8b2sOf9RXYK0XWLkb2xTeanvus60yxw+tg+uFa0mjeT15rA2M
j9YA6ShKNlGn+663hPeoWNArOitslx1R+akRZqdcZsxwoCR2RXXZFyn8Dvjq
phqYtk3a2B2AGLDMkVur9DvU9/SixXp8Enr3vI/F3YAXZpPOumzGOLYzivF8
HB7an2rNSYquC+E4i4iLmCnYSGd/+P16Ul4IUhD/4Ux0MuA7LiXdz+XzVT2x
wwTybtmdMoFBdTjfbx7WqEsCIalcWAtkZgM+o1ybdPuXlBYd9eyBpH9VRxCL
pUT8JptMDQ5cq4Bncnr3Bu49iJfnks/kgJDGcj4l/AEVajZ/reBOaFVSbD7X
TCEqDKSl0B42tjayCXDm0egJKNvcHeSRzVGcNZuJT5PFAmG4OceOtMdef5Gz
/yI9z2TFutGDtvSDoqVVSJFXRdlDhhB9Fvhr0qaHQWz1v38rrKMgEC8sSxuO
pWNcoXMg7Qxxt1MF7lXURcAg6q2HdP182qutxmd+VWhvaqBRnnJJc9qsCuWF
JUW4kxfHQfmV9PfrE+y7WrVlaFjLn7vOJCYmlFJ+Jp9ZoE47CEytq+U0HGv8
/n13ZaAo936aUrBNPibv/CrjrEoOGQ4xMvdatSk1GE4CjQx5LMcc13g8s1sW
UO4+UVMsktvuVkAqMsLIvaY1B4xF35r0aZ5A+fpE2KDNth5O5mXj+EOqI9oI
AkGF9+fdIiZXgOT5CBb8HrOgqybwczgwZGyf7DqrvKlpKckGRHGgNP8sl62L
lSyq1xAyiKgHWyWHQv7iP3cMa3x5s4RSFRD51UPDtb4z+zff3s0AMVv9dpiN
65pBX938GZ0FbK6uhv6hq8oVS46oLpC5TadlO6IkV8qLB9FF3+43cgay1a6p
+1UCYK0jcXM36GSdNW7dJXZrq26jtsHEXUK68uJgqPb1spY34qTWBTcKX1Cc
RTWcMPFaEdbSh85KuVxLxEm+WyEdrYnyh+5tFlBf2OoMuOGRuZrt2yooWwxl
FcOyJaGEz1tBlqshk0dZ6yGrcIt0AgdaL3GA5CIL0eVpT3Yk7pAbn9BRSm1w
0htjcN3ARpepcE6SPAFSaOhebFlviaq52aqEfy0TVvYVtiHzoecy2WxptP49
HNIrXavFj8k4cReJYaW6uwzkwDPq5T1u1rP6Sov3qIQx0We5bsuhVSO+KeBa
pFmV1PRh01t8rDacpEsWsX3jBAIz5pVhnceC+kEBIR6pv1U/epW0ktI05wAi
C1+Ib7JSgACqm31LWE3EaNk7oQGhJjJ6CIOR8K2dxzJ4DjP63Lp0c90ZA8Za
cEfTsxjnTbRmD7Y1jhMOmPIU2Qd7/Q3w9FBwsGBOCjQtvKH056txL9e/7cy4
5rYnCS22VzsXsVauS2BoTKt53UmOUz/BvcJTPYY9vSiYMgmmCJgxbsqykUPz
Q6NPplmmGO5mooJiRNIEyXqQp5CdWoOXySFmfLpFtdw1vvkt+7mBGaNX1T+y
kf9eULbmbgS9BezFlCoRVYSFaaUPcPI+GywS2LcoU7ne0UW0RkEho8OsHY9L
jClYcTC+spFh8Q+nIbSdA/ZB11eQf9I6tsAbsLV6HiBaXa0YseZsec8MFXhc
kQunrjBBZBztmd6G44YVjq6EWFVmGWy85vP0yFQKILipoitKThBQY21vWeZG
t+4LEQH/u1br/zLCwihR6rgDwUs8wiy/0I7iYL2p6/bnXYUz1Y80h+1ta93F
4569Lt9qNoSuZzOmmiByE2ToT9ieXzivzUdxlkScIpGBLkjV/PeC8SLpX3MZ
NcN3fuFjvFpH07lcTQ+qlLhNPUKhO4K2WaUUx4B8hBk69vsG35yVl2kUwkKK
srhsL8j50OWxqFygjKW5kDz3nIn3LJG5yKpxV9X+PjYDkoTH1C3zOfw/Lfpu
h9LwPTjfid5msC6jD2pXb4lq6C0/BhNb52Xnbhzr4JLf/c+8HmvFczSWPsTk
ckylov1JpAUfPgldI1tJV9fQgEId/Bpjui11tIGgI8Ey/rFzVrg8bMZCtmSF
2eotueFsaTcb6HzgoG7zI5OsMlZQzGqb5BDdNsVWX61pGdgCDYhTthhe9l4q
64jH9Rd2jDd2rLFTgqIlu0vcJvxlPDqgKNsDegn2Ea+aI+vYaq/887ixsSpz
bXpozKf65tsbs2WHCxaZLbwUoU7w5MIByrjK7LLqCt4ge2RpU2LUAjD7AbJE
4FknkdsjrzGlvG3Lfn/lKOCCW9X3CEUs9RUNLcApFMMwl1IhxUG5NDav154b
eeyHvN2YVWto7QuKptEwgn8RSz062zNC+uJA7utQEoERXb/CN1NsBpYMwvQj
pIyLq24jWUOYCKyAqQ2bLTatB9Qrql67SGvlQyC/mnLVuAPNEvpxfltxX+9Z
tJM+BdmWpl5TqXuj3GlaHTpPKDR7Q0DrMElLxRh8KRi+js8nsbtwo8ZyrTbM
YkEM64UMZFJf9bDBKifDFMz9fg9QF2bmxE1Vggld6FCvnudH0iMJvtN6M4iW
CK3q37m6/LUbMJQa6MCzqiXDp04ejx8aJhzUjIheqk2wpHqUaufJ6ogwgM2H
50ScL4DrnFzgWRelQwoRS5TvmTSkZGvoBQt4cvXYsBoP0SHe9vzCV5eDPBDE
QUJ5YFC6rs+N8P1JweSNvI7JbUawnvk4oAx9htrIrvesDy3KqtlL3CX//Q0k
Yoxdtqydblc9Cz6rlpC9rzKR99JnNQhG6ixdXg5TCFIMHUF2YjMlmaI1iqUo
hdGDCw6D4ZgTOC8RYAaHB2oN1Fun2cJBEvbB11kXhG3b9uwZXEBU2qeV7cOj
gQLq4a2r+Zyl6tpBdCDsx4MUUWhGD/4zgOzX/TwQzr/1lFQAxL/kB721L+YI
lMgPngCiIhcWM8vpPlRHaCzTswRyyjLf4aeuD0pixxoEegwsLwW/1p0/Tk2F
QLcK/NqiYmooKVK3iWHmGI74nKJBH0WYQXzoS2FgldFNZB/7wPUl8gBPDZw4
dfD3Qn37cQ9F1U6K3RE/8JVtIgJMPgPUu6g3RGRs2Rv5kSU9X0tUf6cgciTA
Fhb2t7/rID9C1GibCWv0mVDghqpelqCIL7Sni35fAzaNpZNjoA+NPNtp8W1s
vPwbeDwj95GNd2g6D/1ck///wmNXmlh/YQWWj+BtTI3jRngxAh41lYBik6Rm
OQJUN8xMeWR8wdKBmOi8VIXUWvsjgMfyZ83LBUgQYODHgh0u5wCF/Vg4w/O4
3U1r9pni7r4wcuOdVRrsSEgrUtqnrj7/IcDXelGKYNAvB4lyhvc4ncvNUlr7
w+fJOtJqCvHLFRjyBgczhIPfVdRyhzMh89LYpB9F4KaMebDeshF4U/LaCxI1
7pS7iNf9ZxLAXNvT7xHeyYNuE7sTaWs7fL9r+kOxEM9nIEUStjiZI4J3B7+A
naRzfAXw4Sd/xZrGjh6ulwD7sz0lIOGkQMaQRamghtSXgDuBhcThVfTyhGvN
eq5xPkhiazFN/xg4t3e4/4KjSZvvoLKqTeAC6fDWzIYJ1P/r7RkfFpZTW6fo
W2r2ehKyZ3/AMUuHIMJfpai3LgU9n/TpAvGkZKW7vevxpdk/yco4BoKuXeyG
V3lU7kn1fTdDimZOeRBeVxylNXG4IQJg5U0Azl88kLKOCpna/u8WhYD1Spvh
9hs3ONUZs/RYuSc/2XzscO6H94/+GstfavuktJFIpwF9nsIXYwu8CgCh5Stx
7Rtn0Bv/2GKBkuJor+LGABE5WN0qRgapSbmek/kfoerAoGlHyX6uJ3VgO6AI
DLy7f0sTC6PK6k+Bq/6zYIL0OaFhPWusYhIMR6ULbve9OoexFha7SNxKAmbF
QfWEixvxsVUsLSYMEauM2vQ5L5EYcWrTOJUGLd34HrjWc3vPYxKDKQRld5Wa
eKzVvtl6aUyFlnmbYUgr9SdsjwDawKK8DOSYh5Hh/4ct7KYlrMashSWz9KBK
4gctnw1/0KCjxmyCybBpIO1Y1zg8B7XP9QYobpURE3xbqyDyan61liYho7LL
UJsjEl7EDIHklA76zp/PiR0FuTFAUmToZeRNHnfPIWKUkwOXUO/J8XYUlHU0
yKqjzmXYsMjIYq6MCx85Kvxz0RCV1u+7TKVdCYgPDRmtAlPgKGrEqGe06R8h
ISc6Ml9ovX1Y3SZHPMMcityfNIOcWX+V5bY3h9TFalef1BGpM1MPsEzVEPQX
ZB+x4iL2RWWljbYoxtudZgQnNvX65q26vlOQG0g8eKb4oRgA+rh5FEhCsmBX
OIJKPQNzeNFIqu+1QVAP/+Ku/fuyl9xMTIPavJiZBGffq4/eTK8hAaNN1oiZ
JEio7MQ4qFxOr9Jb2kocu7tIbWBF0u56Gt6JbCFCphjcU33buBpaOgMdAWbh
mtTNcNCeu0FGVJAK7uc/7645Ng8P9PIhY+SF0llxyRQA82sUa+C0t2OwUj0z
sdgBDpwsttQigziWxnekSIntINepqfcQuOfb8yhbwJGJ9aIgxMh9u1/3IMoG
VK+pXimzewT5CJNc65xwkv7rKkZv4cKX36bKkUziyqdb8Ybj0qi+0sxIqn9E
Tr5jLSYcaZytUrsLm9YeKQujkdnQqjsR0b2z97fUZh8ofBOQf5NmWRMK+N30
0Xm5h0fwtdiGXOVJqyBebad09vb1Q0xQyk6DQ74DMB4RZqFPcWNRZDByI+Eu
Iq42j1p1T3BMklNJMHihwXZYRfkAkBjnQXLf2f7vW4uP0XDrjIIosUD720UO
YpJwtQOzluGe1iRVqkczLFkhK2EUeBOhU/Bui6CiAnPX6KpKKqiu5Qe3Ns9I
Eq77xbiwposC3X7DvxuYcnCH0/ULXMt3D1FrmIfTu3P9XeiWJaX/kQIfm5m0
VbKRlZ1XMI4yX8WMvTS4ZTa9aoBmqVAT/qGIqsGZq30YGqgaAJs60lCxUc2p
qGMNXH5/FIWPx41Hpx0WEp9bhO4vr0dpj8GcnHk3L7aXvgngPu+1w+Ty4X9b
MPypYYH4JkXfVa8DejBq3jDVSTwok8MQdWrgqQ2VpK2JfG+YFa3318jOPLvJ
U1x1UKdo0CEyvFVYpzEpbUMTTiDzxD7ME2rfjWZppWPrUb85M6PgSNMcTjKo
fcXUbDSUpjCV1pnu+YdGnGxWRcRmtXK8gkhMO3JWjWNniXFjMe61GZo/kkfW
FKa26Rz53W30ZMaEKltzYTD+drl21P9R8GHFPAU8smMIuyqaa7WZ5rr/6c5Y
1DwfYuNyQgicw/DmqiAcFelfGErQurHkx8pmAMAaGVjnG2YqGiQ0TitDLRAE
uWCcTFvfZxGuliZtahZDwtR3KFEk24VCM789gHAILblPwzL/Cx8EmWI6j1Wy
jEYFv853P2Nz09fyEBnegPsVLE6668Ms48ZAa9LJjgl7abtUejhRVY7jS/HF
kFjgUvtD+7N0QuL5LESLd4kdtfcv34+29W7dFTxB8Oa4hRTa6QKQgHYRyvJ/
VHCezBCkppOo4g6si1vXlBA7YQlRXAhVxU75fjZUyyBSfNP33AoX8iDGseqE
5WMFxDZG21cTObcYfd67wE67Db8SYAZsE38SgehWqxhnvKAiP7Q7DbnW+Kqi
4PBcxBACxZqPmTkgpKXtZ2wqtPFZ1E/nDHMB//2IfAhGbpOwH11vvk2TSvCV
chQE4odE1pwg3p9qG94C0JxOnIA3NAW4OVX/pJm1yWXORXJf0YqCIGzqg2RA
/vIEtyCTD3Gp1nRqP2e9tyhxuPc0axQKGiv5yQPkMx9q7q1bLG5ynMnkwFpO
xfjqaBqBVDPIx38229F46CBsubk2Ql2rKAnW2hSfHpDHmEy3jpnfKs7Crl90
uuarUfJokh8xRH7TZ99Sh+I759ozCjLvT/PUzbZGnZZNwbhW1TiYhloYouvY
KvjL63Ye2SCEV0vf7+sVuQQ4ME55o2TeRLwwjUaG1k36ChWgmRihv3CYXxHv
0Wym8aI1sdkwyaY0P1Vpfo0Esb88u4aEgl9eOQt3IVQdM/eZAWhL4dZdR1RZ
ERi3JaditeQjE69TMFyZAsNRzdsRrE/ETFnTWyPWk8Z1w/kbgUX/hFqgmS1R
zJBQPyXXByDHq2/893pMiqBivTNENxLXFo34FANMxTz5UMCoZ9HQ0/KiU7hs
3Fu5hXiHy+MvSpOY7s0aAkuGTPdbuweTd4DT0rBmf2hPQWxO8gfqrxSkYR/W
AS/m6eyqdQKTcCUkG4AhI6OOH6jJWf2X1c/l6hEIbVInZbzSyIPm0PqulA4Y
UmJEgoREYAMYiJsJtsj2lSQ5171nz8tSFrBR9NW+tvc0ASTbRNBOKG132A3f
Ix4G1Z9xBxkWWi9jHTyI4YoVJF5bflOExyA7grlmGexbH/n8+fVtLAS/C4o0
8Kvqqu5X8KYvwYj73guHvG3gNQSlXZZO1EsKETaUO+vr/Liz2/cIzSbn2The
yYpuEzI91MYTMZX/Fg83aqytkJVpWacriLDn7EKsSEQj/54VsRSJz/KVPnp2
AvoWwxdQE7HdmY4WrsBcgvoXi/wT6tZwQF5q1pmROHmAlU/sg5YzVo/+HCgM
x7Q+HI+U6C7wZINT2cWuV8yRo23d3I/TbWG96IqSIOaxTLvTlYCo4rYrUqKM
BtPzgy+GOKnsGTpwq+HMH2VT8dx8nyymIHtz8FX0xC1jsSDaSduzooA/yx0R
eTNs2BSSDdBqzT/MiQblRPI9vQL042oiwvOLq1D3ReCSit32bQe/bJMwfmzh
tHM0720pMHvmEgYoFySAvqe/c3Sw3s25Useb3eCwzBGDgGa6sIl7n6culqca
L6YkkeFknLE1QYaI+vjKD5lE4uNBIkesFfWfH3iT96C1rW5VfQzo6v+xpR4N
vB3f9GGLJCrAVOv49chMWpaHCgbTFm0XnQLNTkGP0VtAl89SBVETgos1GriK
4CC0FXWPzpsNFdCBtwoUDVf0Q8qGdj/BxWtj9uqA4cLiLYj5+GkBSZerXgtG
5fWNrzdBiRMV2AEtfAnGrtwA4jCZsF9DMcnj2ItN5z+DQkbat1xdLbFgw2z9
04wvF7eB49xdlunClfzhVucVQklNY0uvXDZRHCn2yEV3IM9TfA4AjGgTop1o
AT3kXyV0EFoiCVZ2UBOzEAdNbl3jRjZPKA/JT0LWiN9GuH08ooiOdDxg7Bwk
r4hWTVubmZa6L4KczJb+ojUwxKxSDEl9Rvp5WSgiZYW5LemE3DAggTA4+6gD
1SKaaHK/Ga4KTI92gFBz54285i7sytmK7F5yZCexA+/KbGF/mWe6mKffbgAz
Xr3CfxJKcVHbsbpaA8Rkwd+gl/qCCn2//6S1mmr1Ss6Bkt7EZ/yyKZcEtMN9
r9UC0/63a1T3V6hfbhCiV1cQyGSS83rJFJyF+YMUJT7fqLoIJNEQ8AmFbx7A
83QZ/wG4yYp8myrn7geBKQinEDxT5rSlkDKLZMp+V0BB5S355Ywf6saLTdJE
LSt5l36J2iTKIU+l37SWKU+XE2y0NoFUM5tO+DZSBbFefsltSBNyl5klR9pi
Yo2pryZ1Bhtm+SrZ9ChFmTuVj4sJFQO7GMp7gQQRLj9lxq6fBGTLIhA1lpqg
yqtHdqngtC/nKDLtg0irznJJTqT6VqKFbhRAd8tIIsDVOovB365/PrOqnVIc
VBpf/Iev1l4GNMKhmc7Tk+5Cxf8YBmypNzYX3wr4qCIXorUQL3fbt/6ssYKm
Rp02TL4qVe8CT43vFB1qDZjIeTaq7CIzIPtS1sBXf/Hdy700vjFKpZ+9Z41a
bwt2n+9tVfQ2ZcMqkWkKzsyH7Qlg/KLdKKpRMhjyO5wPAEZW+afOHMwtdDVG
VF0J3KYQ0i6C6K4LELGHLrFPIzViMkq0KJdlqc7PriGWiMIeD/pCcz1YST9O
9moESyIlx0uyCtKIgvrbjo/qYFC/37pMpvOy/ZHfTbTyYlIx3fiv6E+S9R+b
QzCZg8RwSlmsKeKi/QfWQy5A0/Q8dL7uiQA0da23bCARQRIYQeRJLJftr9o4
uUAKjkqkGCpCMkZpM5GzfeSMmgTNfqax8Lg5MFejcWcJeja8MvKK0Vx2QFam
DbbDEG5az7LWZc6H7TE1pjWMoT5+j439gq3GjVophonJxkSEe+xZ17bvQb7a
GvnCKrqfz+M8H6sfVaqBUH6zbnUso/soMcbRCejqtpu2FoTYSPhIkhOve+8E
jXUbMZ+ef/GtTMfy42ZAT7xmP+sgAmIk9R4yUVjnq5lBRN6xl3SYqKRJ86jN
rrbbVJ3xcV2jvYIYx6EhBvkutQUFUXOOg6TsteVDKGoz/C4i8wx5AuYrcOrW
ZaauKvkMegbGZWcZ0iouym7NYyNh4LGx1sUL3MNuAQco+rF5uxgmTGbtb6Y8
IFatdqtF9yMbTvCA8gEpOzg0sJsp+QvQTHXL0+aLkpUfLD4G5VI4PRCe0h56
/rjYqTy7Wm6kTakm33hKoxH/Uf7rqvcDy/P2EDeoo6BB1xZS/8TbGRUq8HQt
PkBmA0Y9rvVJtcnhK0pNnJeFExG42YzucMnYBYYKlbGa3X633mDOMTb6PNaw
GrJqVInssEqvOeR3CimHiPB0k0NP1PZ6EKe1udNVt/RR5hzCDEh+mDSsg1zu
PpxNGvXQIZ4PlYSaizLlp+IxE/4LDdrGd2k7/xqE6ljzmy+yAmq1iOlRuBpm
Lwughs76m+ZM6LW2KEQ8lkY82UnulkX4JTNf4l4PXTFuXoBSmUSUodc8rsKs
TKXD+3Sov8d5mdfeBFhLU5W/eXbxj2TiFtprACwBpCO0pSBdNYg0u8pa9Olf
3NapKqtEKOakolbrVhtFMWrfiuIBIxgAopuC1/19XxmOUcnmtnpbvKF/+KlX
+N+I6jiD9CwC4Zgmyu3Sm5GFqboXDZqpPlWm6Kvwp6MEKh1acKJGQYmR+XQ5
kiQWoUFizuEzvWnkThZV453GwecPOekgA/85TYBWm6jnegce1SL6uM6U3aBl
HBXot6btWoFMPhaqIALzQV0QTOVzxW/7sBd5T18e0zwqCP0VBoha185NEuKy
jZZUQVBFMJOeJoh+6KErwq0j1jmyUeqFbMuLIxtiihLC+u895CvdEn/loZ74
623UBhFiwbMNFprH5R7TN32YkiXq8NMIB4kk6Wd6n0btXOBuqDov+efdQo+v
8Zy9asQF8TduIahgRN6Css3kA78hPVyHqtWh0wtDimGD33GGUY5gJNOxEgAS
6Mae/48WIDx/X2rsUjKPqFfDUULourE5+NON/m3nuKjiTy9BxXYkVaB4ECrY
eixkoKLDxL3gebdzZi559hODGh92P/69GBQZbD1X+gcb2vTjOobp6Asx28lW
2UfGZdRdGGKMN+/Rb7huHcSdVZxProj92EbUKjAj4gqaUHzfZ8tSufBmwKtr
AfkLee2xRXYdfVuXWREfHEOc22bhMlwlUXsaODXGzXWXeaJU4kQ3SJHnX5Zf
9oNc9Awpg8uLS1J1mzmvA7COz+bRA74yheTpxrkO2kiH1IE35l8uQFAY37Im
IAtFe+zvliOXfAc/sshNSxZKK33+paheYILPB4MC5zfv5oyJKDy5hIc8qiTk
Q8HWByJLySNw+p33hK53MZoDNIN4GMu23kLMakKutlTTmC3BdVo7byT3Gmit
guG2GPgvfPKPKsKBuP1/YACVReYEpQsglnmfEdbCAAVeX9gdRBhvwjfgs++V
W+g6E8TNDLfrej5SXVnLBBJ8ipIrW8H1d91NaPMl5Ak1KYkRx9CpyIMwxpiX
+6DtKMxUdUnz5rBrKQz/TozyFNUwa5lVZF+/qOqcBsi71fliJojrUE1fFh9r
ARss+fqLfEpuIJ9NxrDtXfUCbH0F6RfRsExJYfARWyUO9XGuWEC8HYGf194/
ICUNkPLwirRjg2BOoRm9rWWDQhfTCTFs8XwirtSt4A3exRTwS6RajSJtQoSp
PgMtSyjhuE13NFOi8EhwVNclieIuIvieAttehfLSLHLeJJIagRImM1SWvLD/
qwRaQ7xrUb31H2haL3hW3CuLMj38ftmCCgU3iQwlEcKcQrrHXFiAHU/pDwps
jBzdnDhxCF72hdKJaAnn8VEZs1KyJA57Yiy3xnqWEIKOWCuiQHiMityeeHDm
xAUhSe4ZqnzYNds1Yd+awaaC1H8vyjDfljKs4dZgmLjl73jmFh1qrLDU2Fr/
/it0NTTJF6Pa8dicZZ1Gt7NT3MybWRNrhtHtchxcUxymzWhrMYt80ozFWH2q
hjwfeCdyrRuO233cwaqbViE+kyLvjY1YlHFrPHnFJhVUy6gaii9Ta2M8cWg9
P2W8o6ntEI++N+6RMEgxILYYOv8JfSe3Tz8cLEVvNgcM7TA+ZF77RSuvC64X
q2/VoYwPbINwIWU0SV0iYujM06n7ZvhQ8Rd/N6l7x4xmrQ0Z1pc+XgvMN6A5
CeSZKdCsM269RgpODxoEf2X+V2sXewM4kvMuuUp7mZXZM+rS2U++6EivQVSa
+x1IqMnqkkyHFpw445rfPEWSkTHPDvAvIv4H1ue2kA82fjm9+jf8pSIDutmk
mipLYbm6nq4L8Us/Yp5h77sheAVzKdbMLGUQX4gEhuezL1ssRxGW9eNY6X6Z
ji5W+1YHv1VgZESdSmC8ELgafKpChs9Wa7BUuaTFczzCQDzl4BbxLquQzReB
kdXtGOJi7NbQDXEebEK8G/8bM3hOFgqKQiSx34vF7q6nrqBrgZFbJICfaZMn
7KnEcPEJCDVJQwO8KyJu8Yk8pHS1bVzduKLfP23uwzMpGBP5f4sqv2NChVw2
sNhAB3aQyicNYnQNBQOl3HeHc2BVk3lMscPL5aQzG4gOIFlE9viKT4+s6Ok0
q0CY9fjLXme/nllnf6OZozly7cU8Hj1Czt9YeWiwo+xM+lbRJgyz8MRueApX
MQpApaAberlY0DFvRNT0d2V0M9wVPN8nkjmvSNvyD+2IR8aIHb8CmIdM29S7
MNdvFiKjr6uYIIlP+uHU5fEhO2wX96iN1uDwnCRt2ZdYUQfNiYhsPdthAER+
ymxKWeEMkr7hlN+fxCyyp5tZnFOTDzRwgSwkon3Dp/CwTGCKDt/F1BGtQiva
z7RBjYJFtwtnRIpsqpBdlhopc4kJ7dT+rtCSGY3o7nAf1pJYJItYNJSfAhJa
e1nIqKnXIrG18e9bArTcwBEuqg9JO/4ahn/f3O72hPOJYyGO2ePYjYNfjvhw
gRt2w1kX4LemhmrV9rxCVv+bw+/4CiO/qLq9ivokRsyj+VyXpq5zMq222mcJ
2SnHR1pGoWWilfcbvWTKoYMIU56jphiSRHkgUnMt/c+riGKtvvSZLqGEaa1m
kElB4/wG2ikgt0R9J2dTAzo1MfFslUeNFSnA9STf8chX7ScD9oYOKO93/598
KdA8qFqYzhVMw2l9HReVJdctZ/t8oF6J6GJFFGKJzVNU4wclJwbW+Cnna6iM
D2m/fQ3Lyv0sZbRivVBseosralz48Mtm9FDKAqOJzcLy9vFMsz+DIzX3OEd0
yWlJ/xNv++SSQiV4D1NGjuUihVwAIZRRwzhKTkdMtMIjdyeUAvYFfGWaUygk
3OPHKbd+L/di9fuxsjojEPJueq7LU0spV67q1fAIy6poelqPZyfiSIb7RIAB
sZ0rBt/uWM4FWiGOs3bbQoP0ijVRjpjbO17Oiv8EvHSxEqD5S8KTs8+QMw1d
nsHEV8kGyq5Eh7Pcn57PftIbmmaOlcnfPQ0FpR0EobywfDlZlaK0wqCecjGe
M71MvcFkm+uulMNouYrIcjyLa8Bqz/WN9fp+frrXYV3dYe8G93ObvfUVeb4R
Qktlkqo0skqEn2OIExY126CY3azwDJziTyrqOUR60/5Rlty9yQ2Luw2NOygZ
0WqAZNaSiipB/5nvflF9oULEsqc+HN/OiW4V3/lL0K1CdNTtcSNbe8VV2dvn
Ytf2gOTfyo+7ouacfUi9bBD1Oo6ATUH54kPiRK4pzSJC9hTxm+4XpQ80OtXa
Tfc7Z3MrFi/AreMrSP1KvKdAuk0RwObPuEm4HrjTqg7m4BP/f83QcVA9ZmT9
ZHVtKMgRLX5gvKPYZ/wfLIBWk1KKiTUHDX7yYqiIaukbpna5XnTzTfFkjca2
1TtsdfevhJnUv8fKH9dje+8TgstY92hOllASXVbxPizD4fke5pezEYQGmVYN
NpOcdJ/n4MecWZmMcEzVqHtDWKLF11+9pcwyO377NDKbfpTUcWfZCdfkrq+Y
Lvacx8FjuF0FXx64R+csQMiSj+Uvm7cWYonCCwGj5xTtqhQBD757FJq8KQHF
86pEMHMplTrX0aC6ujnSPfUf/vdB8gVEZGgFLlnvlb4xZ3bzJ8+bGmU0qchy
uQ29qsBnonZqR+5+xpRG2fFD8drxznxGHpg+ecbAYWj7MZUC+PhthfEeBDVM
eW580+CyoMMOTaOIcKu/t9ViDWcZoNG9q6TMZiiANqobKBVSZZeZqHL2ZEGZ
O+3h2qHUaGgl8dwkmnUdhvGKHxyDEd34ooQxqsXgVUDNzNG5kE1ZoGOSDg+K
od+BYvczSm40QfaseyAU9z5QgbO0bko7iRZC+uMctGh/oavJEV2d+XR96iZj
sO5cqiPBBDbuZ2UUSBhq0+no7gc9RdBLQ/tu9VKBDkDnbLM4ep1vYOxSWcrh
dbbL/JbA66tgu3KZ/XbkDWZSvMVVWWH5eFv2EDPf1Ybkf0k/fHq2j3lrFQCF
9IOJco1Dhq8/XFGh5RyAzs8KVRTCZENlhnUrpSGCODKfRm7CI83PgCTuLKWQ
Vdck7d1wTeF7k5C56H5GkR1bIObWSo8uyut6bbqqaHELrFGjkUaZfttVLbyf
fMi38bkRTIJvYu2C2+uFPk1GzFMzV/+IP99BM3muTWworrT0rlEf7Nes5ldP
uNzMTUgR8wOP4k++HE0X8vuArpIzbh/bNHuk2T39HBsATuabZvkmrvZgYvgg
kROGIPO21Mpd9zFv5zhHdua8RtetojlGQwlSEW7LYsdPRxXvWVaYCe9xY5Of
UtGWIjYl5H57Tmy8K4kGtU9DisZamGuN0rXqJfq9pr34bmT2PQA6PV+Tpud5
rRfR/0VRKwOfxSKGoJS1s5nTF5D0IMbdAFhvPi8D+XC2B9VggVEjRZZO9l4m
hVpRAlIkSzOp4uVrp6rOn1K7TZHKzaSvym3kdAAUb8jYPt0wG8r97/vAlqCw
EGmmnU8kq7fM+z4flJzZAmWlz7fcyI4CaILEHAAtdpOma6PBaGo7BBcrcGZU
CFYnmZmy1hmDh3vWRHuOXDVAwzT/Wk6qYRKaBMKARkz3RjOvogIRx53MoMle
QIVMfin9g0Cco/BObrUPLoSweSPk1mL8gNUULJuMa72qiS1asFAO00bN3d8J
71zr1UNYf/hhpwkwO5J+AYHd8omnaR6nKrGJAZAELz+NC6ZC0O3YCeAPQ7VR
vt8rFcm9fPihlOioRfM6j72XWon2jAQ5DAKw6jFexboGd1z+DMfLCmsQs2dH
lstJTdpjRVVci7PVSBXm0eOtC3aByzhu0xW50EXPwneydGQduGwWbfRKxKmd
B17fnBBJj4ZzUNgLUzsFDx3BejrJ1ytBa8g5x0AlqWO1JeUp7bJ7j/zCE+zb
m9or1mibiob/FNMCh8oRbxquA22+npkPc7cNPN2F3VEsyZXGZiztqjI/LUHn
402+DTVX0MPgu4H13F1JeXO8IMdAI1AI5H5Triwf4Ya5kzOVPqWjcsTJ3n7W
M43dRyVsFWiQW2neQjmPjvrlMIE/54JvCqIrSi587fBqhdXjYp+IFl5ToWpF
KF3V68jYHq5U0K9165YaOdOIC0NJSSK9O1ZXOdWMVQRYaXFuxesHs8uAsBmw
6n7alJZ7MM6gyHLOOumYjWSl7Kc4KQPII+wQq2h3eZF2RNJfZm4rleGilmvv
E0PT/2qBQ7B6mnMFO6d2BN9aLWuahSRUZ0+m5BiuOWjaqXxGsgNP3SGgsQZy
xVLPb9B7OSc65gwglLbOWfTflr+OVOMuFYexrPYF0aMTxx8UWx5mFO51vHrM
DQmGZBeBwksC773SwZ1czYTZIqn8GgpNwgjYZsEu8SYEIYprprSFvz+UR30y
9a68DQqc/k+D+3G5eshGh6RuPlCQIAC+taP9W/9HgM1Rm1J424PUQHAzGz+c
ps1LLlbfgNaflflYegQXFqDIpXd1rLta6+s/HlwjOoMpJjxq8yXnZNfr50FJ
GLR25Jq95cXtdVoFtlG7FM6EjxE7IPn5O9fjHJrZ276KyoBLiwp5wdnPTIoU
xlMc5YxnCww3S4PLK3REMX/Q9DxcszOaJB6BgsKREzB8Kg5yt4yVhqBCeZrL
/G/FLwc4PB97cX5puvqY6ry2rjmk6HK+c8kyYJbadp2J2T5C5nQy2ldfULoh
fCCr2mscGr3fYOU+v19Bi6BZOG1+7wl4eY7u4abahMMS11/vVh49lIpBgmF+
hktuMUcrThaFpzt+wg6JWKSQdz+SCKKsxYlQKIRRwpjVJKtd8zZFuGVvsaVY
cVGcVVWQaZt1bY1Xhw5C/KfJc0b8BtyPlo08fsYwaqLjPaWM/SUO2B/nmLI+
GkmYk+kWBBh4y0SjFGjAG31r95fMzB+pvt1UabGBzC/oMYwYYOUtEpUmcvbB
teyq+bhoJFPCVWOgve+AkcgpN0RKYmYiQTf2loXpwucXgi3ypNzoU0sL/cIs
YFzKAKsgqj0fO/VBnduuPW5pX0u5tA0FfN3+nqixsxk8LeDbwJyKiKSpuiIG
1JQSlHLt7pLeohaCai8xZi7RgxRELvICYw9ykJDdfcJsc1jbOSbl0TSAjUPI
Fi/N7+RjWqafU41b2SRS7Vz842xbl7Air0oJMXsyOUfTzYWjxMVyRtimclT/
OPncJcJOYseKYwIbF8iU29lRxt2dCf6Jcg4UYLqPMZooZJPPr6sHKjZPw1eD
YxPEoDMzS30XO1kxn9oUSq5nDDg9CKR9BKTq1zNw1mFQK5gRTgOGBikkKfBV
FHnVrIZAHDxs45+ohrzkgEfQzMx8KWqAiX70FgaccZ3FD/7OKpAk4RxUwEFZ
2nc0AjG+YnrLj3d12LBqjdIQpuW3Px3XRbh9nsyKdnKCIapAZQtWx87jo798
NHfQ9PDVm8W9trz9+C0UMD9KCR11QTFWRY74bHYYjiXL2fuEunW27SeTf6dv
3GtWlYVpS5wDoh1CqXsyWBZq4TYinx+4IrfYFDq3Y3/anWEhBljWyF4Td+cF
aldv4y1NvQwyt3kZsGgZA365x3WoVTyhTJv/Ens0qUSOMJ9MXPyfNBCNtX58
X4sPdGI9zdIXlUEhu/aVBBEbyfj2MvqPbYky8XH7NJ9F8e8xlhtV6l0SD97s
ToDnbrvEUfFtUy+yVEYLA1aoyk/T9WC0fGP74NMDQ1vCud1Fv3GRrlooYKMb
4Cse7qbzTCCRrZXb6VD1uVBlLCTnSgkYQvmX06qzSHlgCIytT+wO1+v+78OT
WuXT2reBJFF8VMG0oMxcs/x+Jm5P11zFvf69EcTvt3F+W/LCrk1tsy8NtKM5
grIzkIai/9qPXTW8GVFcpaV8HUw3LcIvWUCURNP6tLpmPrscAmdmoEVk4rO0
5tOC/9lrbgAZKJSgUBn3YhPueTcv8wqon/d7xI/E50N7EAp4WxOsnI0nvG/C
o+NGvQQdy1YDNwbF6kRnZqGvedZfNOuPP+BaoGTnIdn4krYW6wu7hoxLT/1l
pIzjNzX6NhWqxSJvEV7zi/dQ4ITG1ENyt5NMFNvwtAVVLR4Nny+xCcPRQXsG
t15uLmtEweUDt3uhn47D6Rs9dR8UT5cPW/bmN27k9+x6a4R2EEIL/CIVFZI8
pI7jsIpDg9SU3Cfo6T8L8eJdz/9NMFEuwwPHdi+kEYDzsPPThmo9hu0nlul9
BP2H3i+0hYhnxZGqBApZxmCdYVNlw02ex8lx5RjC3xsfWz0+U6tp/sqs5lWT
tuB6RRj360Lc5bMhxtJ49semK+wfqO3txJ/KobETpOmQWf9SdPWLlgHHTzis
vPR7LOUklREG1CHqGuRuZyX1vNQRFPHZ2InIVtlJ8gF8d66U8HQEs+OFYLaF
GMXBuLijY6b9FE5JktqRXvhUPO+ym3blElABZlXfPUC159NHvDClTX1Kt/HF
Y38TWW2kYqOdJSSopUcxvDWGihS7LGTAErUJQyIoA60qxKtCH7wBUulnhTtb
YDdktYFkBXZ4gPo3E4JRY7VpeeUZHUTGIOcU5Qxc4lrnUudQrsldG4fPCzFU
3YdTUGk5LrE6pyppNFoKWX3vMS628S4YKvCvP/Jf1nzdPZPH+U04KJ7SyTHB
fFqkLyj0UpSXkNXytKPMvojp3G4j7FTeO9nO2UXvO9ueLkmJg3gicZfGytrk
lHpfcRBeZPb0ZMyiM+/+NW9famemEj3FSWmSfWIpLuYny+jLC02kZayGmSO8
sJwAqqcvrQKfO1vscwX9CyRKWhwO1P851mnq/hvkxMFPWqJ4l1H5cB7F5zD8
UydC+NwlQzXQ0puQgiFJr13froiXzJoZzCAs+s/m9WIbDBJsWMoPsaW31Z3B
pxNxqrUEUvW6z8R78TUFljsENfestxT8GRkb2QRw77yzOennJj7W/GuOPHUb
VRm4SqSSK53cE/qO1wDlqTRhRfdGw7f4focYfirrMmP/FrLRSSnAdSCS+dMZ
l8o0aq5zgdfPj4XOUamlb0C2++R1PJSufnRFMNJ8xF1t85lHNnQceJY1zjbL
edHNAkcfCj+AX8K8tFOps3LGBAnXt+Ns8fdtTmF0o8HQD0BuYyat1DNIj7hw
e2sSqjrV2rv/K17niynJKxlmkt/V/MXbLQqIgjV7aDJmCR7i4QbSzIKchamb
SxkgnXtaNMaFu7XYJHfXpGTvAaZ+JolIdssJfdG48Ph0RvxuDbtZ4nu3PpbC
ze2NsrTaSt6pmJxe6g6zv9S9axATwoUQ9WP+jfpmStGhS4+BId5343ksJA1a
5FmFWqI7qO4G5I59MwteM7mYYxluW4hCRVexbZduCHFaG0hkTqqntNiCtqVd
hJ0F6iFM5coFNLkaXINwNHoCXwf9xL2yJdsA/Zd6VG5MzgIDNU2P+i+u1eyQ
x8qM7Y9X4JhNxh/k3yyFdG20hH46qJLbaYoMxl63y/Q9cYS1zRDaKrbJbQ2F
OB6dTeMIvc/S7cLWAysYb1EPpiDbDHIpGIxZbJBZ5mOOX6LHw+ksPR7sBDJj
6SF894Ug4uMZSSb9GLYWsJKCSsEGm85JcawPdwqfSZqPsLyMOSGd2RA+yj59
cq7z8I/ilicqr2Eb1k+uZ6EcSa6rMA+18s7KIR4mA4+mec5azTHzFBINopyt
ctOfJbres/qlLipzaWi3k75moZkb5634rTebf2DldsFOXQs9THuYBsOFNkPP
jCCWrwNjLGNqIUVlUozqh3rT1wIwG0aD1vdlj2yWUPJGRCd6XP/sJQ32xovE
o4Qvl0LxTmdelQ+IdRkmgYF4+FrQRaxMw23wsQY4h2sp0guW5Hfp4XFx9xgY
TvIN+wad6IoQ5PTLswJtF3BsYXyn3R92mtHa+sbkZSKbB7Oo8PpXQ5mzOyfT
34127RY/FvX0cc1zxl5HREaVrYor2fRzuZWwnEzu+C9KXuswB3b3oWN/uLiF
PbwI6PHBQw+ZaIIkh4muNW7hJqflFRoi0udXVdDONvc9PRHtBeZ7b4aPscfh
/ZwP3MhRkCIHsYjuYTM5XAQ3GARpiuslWoYy9/GTuHcKEJfCiYwkVE8feBXb
7z9BtqnxLIC7K0rTGw1IrJOJkwfy+xkxoTufsWr4zXz0Lsa7xSaiwDjCAA5E
S8Q8rc3RzPvn7LvsflcYBzFaazdSEAPx6AFUJDlf8ndua2o812IsHcxUWs/V
vmcaSH4liBHcRspKARwocK7SeXklE0ykzJEkgiGagmuCe3gvLw4AeX5+RVYg
6uvmzx5OKzqPy/FOiKLhFwXsrxNSLAqiJpMSY0LI0oVbah50NlE1VJI03NYj
w2/p4SwO4rz9GSpBzc9ALxknFchhhSW6tutK8Suxp33Jf6bQN0AYk5r/hw5U
arDfdzhjIEOz59bajNjH6nQPZk4F3k5JLzAQGdGf2KWywthEQ5QGb15t/YCS
JqZTWxP1PgBunEaczawrx8ekE6/D02GUHFWmO31WxspnM/pUTkFi06kHpYM5
Fgv7X33GENRd7LybZw6Q03gxH4SDOTZi37IPOzQVZ0cWyr2xx/BdswsG5Kqa
eKB2jnqxdkkUqYZIjCFuCTBHPNRgZJRhDmNkp0c1zza7tLDdaztG+9t5Jawm
QziXUorJQ+xR3ztJOnv9NkBSMG3zQJVyey6VX6py+QRGnWUos44pT7n5BWu/
c+4s4ZmnbXf1aMWINmGd7SsX0nwN0ax/xxhVy4O22eqDunCyguvIx98Q0Dgn
kVGFPboHiRW0Un+fU2SMpPv2eqFzMzGNDeDHb0X5/uU2GgOtt7IsPXMVHmRV
bZHn/Zjdgwel4p8ix5tSxEY3ALL4V3Hy6eDqrQYDdexL/8qmgOLp0cGbbDbU
pwPpLJOCy9/+LJLN8JJxKd3oQhTxPi7zdgcccoZihcBhoWRXB3iVRzGjTil9
JQhSVhK+kTzZfbMVdxT7e4p2lz+/tdnAsa7qnyduwvm+eH4SdYswYUNYKzek
BD56DhABtMFqtQL8ArwaYrUNxoqR3ab25kuBV2Fx8XhyQ7PAcNSMxFRx65J2
sKgW6M7dgBCfEzqDSQJulI10FEF6V38YjB+LRayiuPgNtuuexKNnfqQEGEsw
ustJ9VUGoVSJKY0hfJs2iBPjlS0seOI2tX6/J7uHeJTU0Tu+d34Lg6GIOhfo
cbXlc61Nr1eHdPSkZYwu2Srwf3PEIO8QKUD/DfMRw12erTReoEF9DP47EIBp
LYKj8PW+FtC15/2v9dGcfSokx2xEP8CZ43uNKSO9sk0R6dTHV8fqRDFPzIp3
nStAzHFWwsgPJASe9qvjKeUAtcbcU8SVwKOzA7Fl4uoBbiS9s5gN0KPztbyx
C6qZ+/t5jqZtI+PaugUA66IYx/uNdJiuhpAo65/P6SrFbzpxTEOxjyupLxlD
5GiUrwEq9+zj8I9OgSy4SmruslFSWpV14XcZcriaRESooFvkhaQNFfKVSCuq
fWaIa+iAX1rksfonKOqm8/s3L/Tjnd21E/6k+jMssMSKgfV7Us2sUT5U5aJI
tzJnW76EAahLvjj99GYgm1mDZ79QeJ/geFn1InIi7ZkET/Ie7d+WgNxQoLwI
0A6w2GDKwVPABn987vypmBC+36Be+7Rb67Wy7P9aAv5kzX9ZGE9tslG5vbgq
1ZDcty52aovTbf/FqGs+SW5zwFHARCLvkj0e/l1xVqfk6viT57V98PLkH+LN
NB4UvNLJj12ozbprcSicTBCw3VjJyW/Yudg8vzgy62Dn2MVe8cT6P57tOA+t
wmLTbJb8dwrhf5jdtHD4dzVaY4yItra+UAwpM90Rp2q0xtyqfTlOCMyNMun8
Xr8Zayul4qrg2zXsmo93ZmAbiCCgLFDW72RNdT3n3sKw9HmJQ9PPZ9DFryEU
cPVxZWOV2oFeQjLEKfigmPWHbckJuQq8rlxUiG2NtthHqp8S9HqHb8RSKgIH
FlPLxDMMKT2mRLp/C4pcF1bytVRG5bixGTGrFH20CzuZlg4odYyzCZCGaCKd
Qp0nTu6otjy5XAla58Cnc4K2FkRFEhetYw3RJLlswtkSEZifgumYGVKWN5Fn
wk+PyqJe+HI6NtMk+Z5+RBJgF9ciTWWW5PJdQjwCWz/R838GMzYrxIT+uZi9
I3K5np1MtfaYYuQksUaCjataJTriemCbBvk+33coRPHQVGeIRdMeZ56Y+viw
++eYOscNOMDaU9auK94rN3CVnJusUpuetvNeRZ9qpftmqKeUpOdiYGmHBMVE
FYwzWtOby5tYmeAd7+N/Rtq35fF/raCfbwvc3BK2ULpOxqELX/ytJwIL3KsE
pZxAFIEKEoOnh8/6YzdfefDM8wer09QI4jxhFGiQ8C5TtFT4jcFCIi3ZOQnh
w+oyZzK5FJWSGODq2F/q57lnaxsRlr9JCu79ZZsTyEImVlRRvzDSTKH00ARb
ocNKn2cqyjTVPs5Em5//jP4wwKqDhhYWGLa8SkS+PIoFIV0WdFQIY6C2LLHe
X073SCYSP1xdpPDBJij0PfYynkWAgVNayKmWbfyTVoeZ9SxyXx2RCzHwVgk1
Pt9fLvTL7sD4f44cnUn31OviOetq7aB9743c5rRS62DvRYadx/4ubUbo3IWr
LJDO7NVqiKoGtzm2ONknIJuwmh09FHfFVhdNvM+GEhK+KXWz9ZctSvbpBFHz
EiZihzZYaQbITTiJXM7sM5OYesIJ4GJAmV72X1OWwNgTf+ByvR8hTmGIZlBC
nCQEMNyu+HVWA6X56PK+MGmfs18ArP7EtNoRj7+WysEE1pVptUfRB3sUDG3N
5e0UQNpp+swOn8wQJDB/odAgREH/akD+OPdB9R6yOEY11y45xEYRBCFHYPxQ
7DkLgzlPsfH06nHDqsn5si3nkIbmwG0erGiSvnOzS4qEfSDZfVvbkqtqdWzF
dKiKo3tJRFPS+yEdVjXt6ewL74HwLMsh0VeIIA33rSVeIW9GmDuiMnidSfAq
wmCau7TXzWl42WWNZ415Hug2D0HLU2kXImew8KDPj9LClhhgz46G0DBwoSez
/8d3tiQ1Er7L7KN2cDFOYCX9IgYTrwl1JkGiV03LLNg1T9dijh0mDHKyPyA5
yzxkhbXQbf/M6aRd89IICOYNfUjBlVfrFBXZu0MLACH9j3u/c1V0/BaSlVPK
3maYUkVUSAtAjYHVcxGXtfY2obUzHsWyzsoU6D22z3IlJPwxjfofOzJVATxE
3Dl7X3ikr6PCeAUEmZoQXjrBbPrIk+n9L64yyMvbGjJvTnr8XaV4MGC6NYYR
RMoqrEb2GExxoj+2qE5WQgVLP3tWKMbauEcJwX+tz3A5JqxiaTVnfxw5+cU7
9ScV8qFD9clJpq5b2kpmB5llBL8lJ1DZ7QXTX4W0ud/j477fc8iNC+tRmYcM
Q+YiWOfiniK7h4XiYiUTPDLI0HKphADQQ7qCDSwGxf7pmlJOMfzhFsmsBNo/
c9JNM0b6o9fENQbiwNqXw72lraTGmK8G2SUYne5Dh8lSHP7IX5q+AcgrP7NT
wjXMusG/zScOVvDYod/kKD4pxS0buFlgAylMXvgSdVxweNa4zdyd/rjzcwg3
ASDjxAZ5ygxLBQvb2y3110QLXGivJjOZu5yeoBK0cxDMnKtLTXDcdC2WiyC0
R+W0YkItmsCfh26IdYy9VJXUHBpx0IayzdNeJvXrI+jzCgdlD4Y7HfflO9LX
IMMt/CQBEQrxwMEhGWUU8GS5ofexr/y4Q4SAdEiRFoe/SyKoqmpes4RjLqLU
Aaru8wMr1lHWIfdwxq5h8lMg+Rw0YOfp0OdzHWhWWh0veLAGW3OapzWQEcGJ
uGsT+e3XNSrQdDrcNKEp/Yhm98nVtvdgK0MxV/2IHLpr+WE96Ackd6sV0sB+
9WR5CATjjKxklZZqZtdUhlU7M1F4SKKrE2vm0KSJSdJaIfDIof5cNLKz0Pdg
r5vSRIQSJOOS3WviiHBp/YVUNQNQ1/dFCxa4R9OTQ5shMLJGPH1x3VX7uQaT
hBT7Yp2bj6qeIP4mGMsxdUSOW2o041RPN2N53wkMKHEGqbAufrYoP8exZDAS
nrn2esMYODjMUes/fACFhd4Fhz7HE6lzAoN0lP3iASk69BYLF61ibkv7XTQ1
vAwqZ1cD1v6jditxUX0bocn0TtjUsSoAdAY1nh4S+7UcIQDlWrOeyo40JC+o
ZEywMqHhO1rJnRCuVIXH8qIPB21jxrIKxFHUl3QhtdPAGvUQoa/M2eTiavgS
qSTEfFELRWhOJi3tXmkwfpr4NrO8eJswabR0U3kKf2UKcpiwMuLskgGQfAa4
4gkRRbR/lq4CJoUttLh4Pghz98/7ABR4I0tDlfE19Yqk7nH+ZEooiaClRQm8
C0LOMFFImgKoKR7rSxoUKVRMD/kQjutDefzuEK7YpfF7o5Df7ohr8nWWSCy7
2kAey9iOam6txsMv1biEYv6xGytxZO5LMtaVAVuXBXWGklQtT340akNQdTI4
nBYy2YdPKEFD5TNcIjpn90BANEPR1OM9SzFURU7rCZcsfJyWw1q3wJF1amOn
WsOMVzq47GUfI6Wwxs9IaqJdF7MmuOdI/8CduQKR3QYdlwfu8JpPVOTodgas
bJfZFYYwTj55BOnVM9XS1iOw1SkfF8ZQHUSYjOMkqWSkdTtfIAnq7htzLkID
ff/pJl1sCKm2XF5muSWqhwS0989GwYXMBEoVRRy4AKkFPqheai3elEzbU9Kp
+UuSFyBQ6JyqczBLkCbqd5vgA3CjTN2l9HRbSJpRjw47XveWy4DWVQSg5yIJ
ptWpzmO8YoxefV7z7UNZMx4Y5YppzjxaIerYVJvXE9L4JsUllwISqIwP80T5
K+iMeZ8pmIg/wcfXj45oj4ReStS/NsCPaEzktYY5yeQqJRlxj/9QmSteORQw
6dGxt0S8LsfEYgaqPBdKWrNsxTDLERnWNP0DYU/s5T2AGtuNlISl87FiGiFU
J2NYkoIfKvGLuNv96FooVeEfa3NopVEpPgjBtI6vRJy3b/+e25u4rLZGw0JT
bj1b6hnaSCPT6Jl3u9nJjhvg8Yy6dhmW3qBdGMk6UgLQqMijVMM/2HZY4rpZ
3gyfHtTr5K8gh0riLPurs+l3vlxleXQn5fKWcfW6OnCRkED32CoEeNddj6wt
Gbhdbnr5ANJqPC10Q3aG0al0l0BvoGBjdwvfVXOYYOyoqR5h0uyvuU/uoqc4
QTePb0THj6HAvoBJ8+7whd4vlqQtPNG6cmByudtiGmL0ZsXnApTfjU/A/0wL
UbmJjT6xKXjtuRZTZmS8Q4HIcOLhYyh9lOUhStLolRIcBUOylbqXB6Uvef5G
lNh3lnsi3jAYwenW2qibZ95QSxFTB+dCREZst5uawD4LNwYATYBWZdhAIHjc
DjeSKTFCDpVaggCaqfcSVGP01WKO17z1yxKHG1bUsJ3j8wjWmzFlmCQQDU9v
qL3TmFcHJaj/sIjWBkx36bwgM3tV+ytyP4Tsg6CIuLlE563I1bYRfNZ7OESW
bGguwnxROSsoQ6L6t34q8f6Vqzbdu2XagjrXbuj43HvMx2VVeaX0bQc07uuz
enoQfSVRB5v58gKX+MuTbeZZsCdiQbkWnXYxhGU+K/8/NRh+Tac1ZBfTRT+S
EclvXcqhIb+kVnpC1h9ieiGFeTsxxEOjJleKpZUG2BvlriO39bvfKEEpimYM
FiqlbKmPXw8VPAHSqEDS3i49TS4x+EfPGNOduNM06vR2uwH2zPo6jy0Rab9k
YPVlkwj3JBlwaagxhTvOrwtkZIn6YL/eYxsZscIVuGXWn1ZRqlD5xjDpUCkb
kJ8/SDVOyMfmTVbeen04PEerTnQ4VffWStdfGjDNjsjhDDqPa55l6BDM/KKk
6C7WFpS5FrvZ6sPxAV0/PV5B/Q1oUj5QAz4kb0u+78wS/uR3m27nEwoXXmxS
8PzbYFikGRSVPu8viAhVmHEEGPJwINZ21SgGA6dMHKksQqwgo/yJil+ejrxR
79zRmVjrpr/7r50VvnnG4jPh//5nnmeZQSSEILYdl2BOC0skqBD5GYapsIBQ
u0WTLt0awVqG5DJVPjbgSlibtHHM/X7W8Gk4IMzvoa1sH8ba355GNDP72v7a
rOnBUSL0S2bsNOl9e3nz6BfPLljwRLSqDZa5O9xZGJ8CMaVoFyw9nOR4J06F
V06BrZGrkZcFe4IgYX8l42SgAptu/PHIdrsdkm0NGJYxkNeIr95E39UbhQj8
2FKuBWOdAWzD2DCvDgxXi+Ekqd1zaHyqC6a9yHfOwYAa8nTn722CtznHnIei
amQc1SmONND12UnZIdo1qe2kdbXUvDQuNYSjBQFrXFHvpgx9XR8wBWjs1sXj
oEDwZvW4L9alYUvo1w/lfhuP5NqY3vXqDEOhEoJyRp/6tl9suf3txO0K7cop
HnF86EPYYxTiUgRuPo9Eu1Qif1q4Eup5horfoo2CCH+723gGG+nSFsrKB9gA
M4aT791kiHHzAaXP2f2fJO5RR82jZGtTmhPgojFL/h7sdOD/8H9HCDP6nYJS
YQ2xz3k/QDCAEUIO/D2slqrYpeie0Rq3TMHY2AyCSqQTf3BFT6CuM7qK/bv5
M3Kd1Ww4Gff5J9T2ZtQ/TxPZhg1NYtZduZXN4qDx2gvD5lDaZTW6eAusU8DX
ev1UbMp2RXpiuQRIXR7ux0wxvUh32SNPypT0wOJb2zAUhXZ85QG5KW3GqGsz
J5sc75IGkrDzWbVFUOSHNxgm4p5ApnqG3xPPyNz7/rYJrX+VECTNBme1UqeY
R8RgUkevkA2mHwpPct8Ob9BfH48zTBALpbp8UHrAmF6iMY7X0SlAPxzIYY+t
U8fcGs+srC+7lyMhccuRsOFsHPvBvRy8fa7B1Wc6nO6mxjWwNQJ6OWDztfqU
O80fDNVQ9pMVxZkGNx3rOh3RNjs89E+XQXq+eOVOsvC7ezAEQyiysKyWyRiN
i91cghnJp72UisCWv8Mqk6a2Z5U1I6ZlNlsr8TefaOgyU+8B0xFEsifZ0c0G
hV4t4Y8JzRZMqlFat8fTJuPndg4dnFikG79C8KHQkhS31g4jBOcPGgmwZMzF
TnmABI5/+zMsX6vaNpOUigEXg+4aQQ0oyTiHJG2Zg3cpi6aSD28/fB4hrLrA
50V9QWwt4ZM41P4+5HZrZXoC7Ytzr5g4pYhtyjPo+78gZX4bsSzdERQI3RB8
r1dEu4r7S/iPZp2x5a/MxyoYOYp4Ypl7XjVe465LYlfrZBauhzmJQnIDVBMB
ViBqlz65d9axr7Dgib5PlAZsw8CTXT65UkjgpY46KIwVnmEew7dSnAdbp5p0
r2M4r3TGAWoU7FIrz9I2iOJ+YJ1tIAV0VAlOBlw2AubljQBSBxb7nMroVtJ+
qOhVQcRIgMvIQ2m/XYUpyIw0F9SCZfQQ9u5CSbTXyCcfrPwOpYLDJQeHa/L2
psAddS6uzCdX2rfNjodLSVWNmZZN0ZsGak/a9ZxZDP66ZJ1I518k6kAW1KZO
RsOrk2L0IfyOUHj6ODIQPAZrKVaSpmCC5zYIZXyY0Kg8bU/4pI2G1jpWSAPw
WC7tdvVvbfTJZjoKEXx4Va+3mFoOS6qtiEhF/PqvFv64TLswosn9thXkVqJ5
adCzoeV6R5HTQDd/XsdMfLix2rvx8/wCG1UwnDEu0TBfhfhE2FeliOTciEpN
wpmVjavOGamsfpx2up4tDakH4cOGR52/y+MCFkVjFf4kxvlJ//N/w0rUfNVh
VGSDFGtCE4/GqSnZ2PtFrqCrXmgpZwnpFOr1SsukXjZ+SopSIG+ICLF/8t82
JfHLSQO36OeCiFagVyZJyRgfyESf9kEKPcpBdWSndjjsd6zwqFR7mAIcQ4lc
vVcZ9JxOPBGBuJZBB0UuzgljS1uRk8pXBKltM0H7bf8NkyUm9p0fR7vsIWOg
ILpn30Csx5SCscrtvMR1RxulRaEv2kVkD8ENbvudfdbiQZ3jmyj6w35pt6Gt
mn6TNXwsCaLKj2pX2aAbpX3vVZC45njvgyIx3OgqwJIXNRJaX6M05qOuIMBd
h5E+hXgWFbCw0qLDtdXqeZwDS2ZzvFBNa/3FKMPmmvCRQDQXm3V03RBUY/bj
ENnx/ucxqSl0PrXtxFhb/HPpXbH1jejlHAcc+PUdpLm6AeWy/3Knu0A+KWjC
/MMaybEx7JCiVlkn3xPK2yq7e7bnqkO/hNiMa1sS0xDzLlcSALRbaAQhFIlO
ZjKSFxwtv9BrGWqN/m1FkeEFQmfY3oBS2ZfLMFgmxihG8HWxrkx/mPdqUhft
Br+6UwaBgzp63X4dLKE2w6YSm/pqXlpTyXk5S5aDhxJb0bq45MRaiLJbwV0x
OkEbqa/Ycx34BP226YtI1Pl1NUP5EEZO2Z8IUT6FvtxtySJflPB/bjNgyW/V
AJCekk65ZFNxJ8oZ0IQWwGg1Kio43Z5EuUcq1hAczn6YRI1omW/ZXxF8ZCiu
V34h+PrjzS3tgS+NxNvhpocRbcrq2ArVXU7U4ZCzdFLryvk2YsW9FxSS+eKR
cT+HNZVs4cYLKS9S5fh+Lv072wZ4CLBcUxZpjHpJ5uBrmUYc9B8UkVyX1MiQ
bApZoKckYY7F+8ug/kKRHQT/YTq9ldmJfFhzV4kpyun7g4Z2Bd+n93WBc80o
bV8wOq9NDtUCzDZ9/M4nW4Sh64pD2hA2T/UWO7u3lqxRM37jC75kcxF/BbcF
WbTSXQ7FhvGlagSc5482W42wYV4+B8xVbNa6TLrzE8BnvYE3NoPJc7j60cMD
d7RfN5BMlsyvORoRXixyQweTN4iqy0K7t/7+JVoMcJZOt2/LwHtQ+CICx5KQ
ywPqUhXfuL34Xj2TGXeuYPg0FiTQqYCve4r07dLYqYmhlyEK2cP7BnEouiPR
zp0Gso2ctQXbVqZM9Mut2YjjZMk/AaxWLJ9bPRv7bNIUYLT3V7Okd6geAYig
51gqo0+vtneC229gQlDPvoFiZp3ln3uifFO3UpMB36hvRGsYMdQvvIbdt2KP
hvPvIgCE242ps4da8gjtDgl7yrjWCBUv3dajU1zcyG+8OzY6gZweIHdCNfiz
k6vSN6iLOFAaPUPhTBMxjqh8BadhBAKITm1Fqumb1uQSRfgMgaDRygB3XNrr
wY91SRW5VkWiHILD44gXuakWHWrcITazjV3QffCFrJorKeyZD5ltOBR/9XR+
UeAhizl57YQqTqIYQ7e54MNeJIDXOESqD9HWmeTfXS2q1JCQ0re6X2GTPdyW
MxM8J6Rbw9Ujh1caCZDw6EkHbcAdyJFdvWbmPIfNb6hsB6Nrc7HjDd/2ObUt
ielWjcs+de2oU7ADlO0Tla1GkCtpxTPjtMgxxw2kRzS/6TNzaC7asIeH2/Bl
QY9Bmdfm3SkR89Rk6KhbfRYmWHnsU6vfGDrYYEQLT+v+4lbFDS6aB/Mok3HW
i6jb61X/UVX1MZQBFhbsf6N1qfv1vO1YUtqnwhGtgL33vcg5vzdyRUGYN07C
MQjw8tUeQIUqJL/huMFQRcw5YH0uulRIHYe7SMv8zm/eX6/4pz+n97JNdemP
HujsIMBFPTJkbjcpQSgK8IcuVZW0Ov8oGzR010ZPCZjvbE6o2Ko+PZMZUYd+
FQblW9HxksK48fTT/g3ctMlSrhYCVpjIeyTJBotRhBV+hbelQerCBOxWO763
0g7BHN4Fgt82F5GnN1lgpdDLxxF9YKPcrQ/LmphDWlkUp7Tcr5S+9csR8iKk
ULWmNI3qkV3XQkEJ7sZ0Qp1xEBW4qgk30G/fu7BVg2pQuntG4eOIDIe+x+oR
WB+5x7/aXiPlkrczO+GQbyK8QnNeANSc/Q8/VRd7gahKkMR+HU+KS6zRUYmv
n3z5Q4iqxip8TNev47FAYmVofpv2A/Gre63+/ohCv1XWGmHZnL2O2hqCMOHt
k77y/q1pULBYl78CXrzP5V3LDEfp4a5HEX8iwsjZTNaIcDKG1AjMJwYfah+8
lbSI/4Ui7x06UZkeVVz9G5NPFyPbv4PvkMJ5ULqS6dL8tMdpNs36OAGyAMg1
C33kxY+/lbkMNonfb29sJhdssYVvfeCt89TGPFz+tSCcF3nt+2aC3oU41Sds
hq7WtSTzQ/3uBIEb9zb3+qIkjeTJfQ4hHrprjPAa+YxlfeXFdVBXBbecmzhv
PzS15bazVldJy4SlkXw3Ak1SOOmVrJrCRT2Wxx5ci9ERT9BdKYN+JIbkirhN
psBRCGd6Hm1sYaVGCknqBPEQ/93fyGvmmedENUTnA+VpAoVKWyKAKS8cpkU7
SExh4JufZoLbLbicQkOdLCV+fn8GWPQRH4hA6fER9hWzgffJ+c1MjGU03sU8
MbN9vwnVdUA7siO5XbP9/OjYdmWqPqa4XukkuCf+I3KXfyDwtIRGNMbWWpUn
9g8Twb/jd27j3uNohMN5AR5x+/Hl0dzRZhtkp8kXOPHTmZRVFsPErHCMAu0s
Ci6cDREi8P5b1WfyxJmCmXvROXasfeUMPFisi/REy4S8jtwEFIl8neZdZqFw
r0CuV+1cwwravFCBUJKlWYsflfzXMZj74TW7yq12qYMm9H+c8BaAiWuQDm82
ArYkA7IABZeJPIiABFDb8kTbKUUvEMiZjBDKtBZH+Tq3f3LO7rHn2tgYQylE
6BFL5+dvRyGbs+mFOC2aL2VS19QZGQ6MnkcDd5GEtpLpi5Up1eenobOh3OHd
tW1mmcecV8gN47rOVDjOBzGEXiWY4Dx6iVbsIr7kyJ2uSRSr91qn0g/Ew3+s
GshARWpFo1EWZGW41UCAGS5Bwq9A7UHAkAfqOV1sNuAfzNBPyBW7wGSqCjpF
H+PBX9i5YYjuEgb3rLOuKBWm/FeBTiyDKzdnq//6SgutaRhRB4oTpai6z7Kv
w4+qp3RE7lSr9HLNMfGz3BPbn5v2geoYqyHbPYIGkHU6ZbM6fPx2MmyKQoKW
GW9INoq5weUPB/wzQjhbPMR4hF6s89zs7rEFx/Lrf1pw/2srslTN4ttlN4Ei
9IZoBS4Aihie2ihamUhFGa6gwMRlQSl6kyujRCegx5wMiNIDqpqiAhMHApM4
jJ+p/o0lTwa/gBepSXFo+sLdG0OUyuM0OPG/IJTfNdE4x88tcGSxpD3GHgsS
sLjVuxPvqfxS4dffBT46EYKVUMWvj5oKRaNqettpvvjpkAmwp0t6QBwroaJj
tUWYMQlGccqpcrlt3eCkrt7SVCfBZ12Mmtm7/IWb2AAenCnBkPtEiMBe0R6p
UqS3TSzvjSrvgCReKJs2FAXNhhuXu6aUHl+OKp6qWWTYC2atoO4p3/BT7n3j
tbJb2C0FjHEB8JcFGOjyzLdpN2bZtmmqCqF66pegt9ptx29/SdTpZesy9pLa
skfcqTYhqsYZJA5ap60kI8xwol9utCCQiH358LOpriy2XcyZcyQnhVRRqbUm
hOvh/o5LTv16CD9+hQOjVjba/6dIFTCwXX8KaNZ7cLfKQUleRSoe1itofP2D
BOx8qNuzL513Q3B3Nmtf1EhzoPOX/ZZomsDoJ+PV91kFxLcgH3b1zMdsPbRa
2MuqyCckwaLZTchN6mgvhtpa+3HPc/sfKLUxjY8XPNATh5X/UCiiU6O+NKeE
YIxofjLW0Uwf9kAwW03wHJ2t4KOoSrcFfqwUQfVQA4C20uuJdL7speFj2vDx
kMR/XPEdllP8uf32GgvzUfu2uSoVJKAJG4gsADRXRuaCH/tcL7Q+S2n1c3fl
bz9BGNqAePUMwQJ2aQj67ircOliH2+rIVZ7Bfs+5NXXBTH3CQZ5c3HvkvjaF
1+aRr5vKecGQf8QszTBFqpt3ro6kojNLC9Y7+DxoHT3v2jDMxBM5bZtO6o+w
Zxx6CS4g8IIwLqWH12O5uZxw5BoDobLbyAUI1yyoD0cspGw/HrCyj2OF2sKh
l8PHUzDIeiANjQyv5q6FN+XeRQUrfLHiUaXYKJvy2wM1UaS2R97YEmoJi87K
qY/5XkVHeVfmgQDUruq9m5bbFhUk4dRqskB/+afHikPf53tMcIQKf/9mM8L3
1T6WGM50zZhV/voNrv2tW91Jsz6hFZJiyVMuwxYu4JZz/t55+RwZ61k7wxET
LvIEWmJ73ENcfLQj7yJHtJplbKhe77P2zTP43FuQdvNpuubInSwZ+ZyNCCIY
F8PFyXp/r++CsOweOIuGd2g4nM1o6ROyu6jntMVLLzi9P3QUShBmzKun5Jeu
xsfamAK3d2ZFcJW/MISiUufefSF+8N31YYmkFxo0MA5Ci7/4Bvz689WgBcuF
Qb1/A5KrVG0ezIRnzrWHTv579DO5I0C5qMiKOFQzdG5ZtEe4gQ5pQ0RACRCy
S8b8e32gWIG7sZBRFNtUZrvT5lKuPUW73DHJ6ytBNOHCmK4mR8HySdXUmPni
CPLGfYb9VysKf4hXe4/Ipw6aD5JOgTOT9AQasqljuXB805CgY8F6fZCQHiF2
D4p2+zEnmH8bPSAp7d55FInOTrCS8yypDRqxmAEoWQd+4J9V/kCuPtWUgn15
fdxxpfo6Y5+zrDwnZ7x+GNzWNY1jBq8hI/Bll8cC7QsiO5EXA5rvgJnmuSSw
LQ5/AYDK2W9r3PKWcPwj4iZ2vOaNZMSwMyLq7BL+SOD4JD94qlUsTRAbjjOG
WUYgw2tG8o5DIDxW7WROHClfWVBclx6AtlbAe8gZxaybtCfUBrVtvPElIIl+
zhzblLJLiF3IZtBPacNJ96a4wdmjsRKv6h3Ch3ay/JeVNzRf5vhzraJ7wLWR
MvpFJkD6Hw7yfcpKyo6YHedrQsm1nwwUIzSTLlefaYNMUyxVcbqMiLVCVLl3
oo0A7RaznQ4DUKcVmxMnU+hn7g3YMQ3IVNUPKhModLkn318ipgF4t5eAtyMB
t6Ee5DkI/MfBRpZqYutlHtWlE6P6KjZOkGo+RWriPgY0Ak3Rk2TcBMQ3Mr+9
bSJyXysQuNFWdJdtuGbHtM7aiMxfo5ttetR7jlsB7Ge/8Wx94s0gP5Un6wUe
4H7NEKClRUfDJjtx/kvwwI9GgF9wSiO/Y4wNabPG08KmSLlE0h3JziO14S++
sU3XAiWE9IBrTWGixXX/yzXf4cQuUlJ2p/0onXy+nJNKLsNJw0ffm7PKGZMR
Q+1GNeBTU5yeot9M9uEtBOiKQE/jCt1x13T+p7AhKTX1HFWhergfk9HkSabC
qXNdlSi5cwZy3ywUWqBqCMOX1Ln3VfkpsK086zi/IXX0tMunO8DGOwmB1kK2
0rQIAQeaDPQVTs2S+yBNrwNMYRmrIK87zu/mIMe9+IwqwmwOAB+capw5f8pb
I5xHbU675Pn6EY7r7nBBD3LoJWwptmorLO88UFuZSdrunbxsx3dUF6Rrlakl
qC0EVUb9QAexO8lkn6pecI8bcTNvzW7rebyEbTtZy6Sdv7xWTmLHSimooQxV
EtKZU127rW1DY60mM3Kh+Cu96oaAQpzN/lFxjjbyu6hYDyPu3mCd+cz8zsqX
95dsxP51b5uJazbJf+lvz2abjuVDc21f9iaJv/LTbNKbPnIGpF1pw9v4FE3k
ZMikv0LTH+cEc3zql13+0A+ddD76iTZJ43RPF68FzYxH1H/DRBwdqAyfzvv8
5NJkCXft7FQgnQJRyqznOqRyxLdnRf7siIJFIlBhWHGS4UrZxKCHc/9O8ydo
pzpjrNK9o0D1wJwQWC63KrMWlXiycDrv0c33ztJqZSIS3+2gnGM+Z7nd3l0V
AnOLAAYCB1CMhriFFlfsGnwgZrXTXGDK0wQyYphHLD05d60Co2eFqvmOz1jF
qKqpkoKGAczCUlgMGtDeIxTcuomsZzsKcsYmW31S4BCVDykFMJ90gVrOLNL2
0lK6LNQMPa6kvbP0iBasxtLiND32Ge6pKI+59VUdD5lwJVxlhp44I5p5Uw2s
j16z+Pj/VV/Ea0O/H0zMhS3BMl0EInWxqPY3UUZNdrZvOFEbkKuH24fW+RSY
burxzRxOgf/RhBUhxOgSP6iVXntz5KEKwvcm/yauTAPrMLbzJGCrYVvENARX
jT7GjR01PRS9bhuMeTV9jGK9dG5MoZuuFZQjXJFHrOFAowzh/kJ6Q+UAdY3K
nh9UKPfkPJ2vYLlxetRvYc2SwvYebWUCCbBYPNNNmBrH5lEkZTsJHTLm4kDA
Q15D/N0HKShEtx+QpYb3vQ8DvKbgtBl3OA074a8rYmuiAxOQNPBMFYRTm+pH
tOM2KEFZj8Ex6W84GjBlFnQm0Zxa/yBatVe6rv4W2w84pl7vq8N4Y9wYRJFo
TJ3vO2cWIU4o2lejQWjqvq3D3wTPzdol2wQoSvy0lWQMd2deam2iiTLWu6IZ
TpjjXt+9ir0LD/yGNScLWRwO+GcMJAxicJJWaeQZ47Gv2uPwv2bnn/+KtLuD
hLnRlFD4+aml6aNrQlKxCpqW9Js+JxbbykYvjfqqExeQ+n2Gu3lv+RKB3oBH
A7UTaCeS7r1m9kTH75kh38EsYoVhsWaAYOExNF0twuqv5cG8S3QC8uJIVApU
izR8kMWyshFivv4kWr1s3i0fpGZcBkEwy0J5MyCwxNwd/FVNiNoRLxqqHK4r
Tstx0buUFZphfTCp/2dPnvttb1pWkLWITU46NfKWFe9b7AllGnyofRfbmttm
m7jB5uLshhuUwBFeCApL1UK7WaSu+k86aGyJ6EEvVpPOoTWZTZSF8NUq3VuE
12Yk3WnXHpdaaCgQKW5TrOrCnj6yx7jOUv89EVYHBVfipI7kmOVey3NIHOAU
SRDrHvvDsLSsf/k9wrMn66mOwvzSimHHSpmnsp7yPHksZuMStkCizUaQbfaI
0AMF2QmpWfrdPiEIViWM7uk3MmQ7IGmotZySOpAO7vTwn/yvSNOZaZyRBVCY
oUcLS5bvWVTk9m0dlyi6PRwKCKJ/JF3SOAxeZ6Cw4hJdGrbOwkGEetleiCRv
FCXemCKPfH9Hg639UJy+FZBHbIROgjorG1eCehjaWhej1i4ncYcv80uYMgHe
X8oqEPh4LUTa+/ya2OjtUMYzWf+fgnJw7YrPwCf1nXqoe38vPChFjZlWS6lx
y4NVUNsMVfWsw5mHpCf7rxIOgqptGv2xEYf0DwCWhkZbNUDDANBfYLmx05j3
4jaV0AzCmzHRCaaQW7NWq8dKLMHky3Om01asYQvHkcxjJiLPsHiYryMHuW48
ZF0cKLiqQYK20hfkumHqgCnNfJ4vHhCYF4AkyeWsqktVkQ//hCl2Ymy+93xP
ZUhTaYwfJRwUuGBz/8oLloB1yryaFw3CYuZGDZSY3r/pUC+PVXLaxXXZ7/sN
yJ+7uuvUwQH9y57bVrxZZ7EzGT2NcZwyyvOVKKWQBOF0cBlATMs5/I7BMn5r
o3rh9YN4P2u5rCzlJVLyrCiOOPplW3xGCXI7xvR7dZ+eNYgyX0/DF/pCwz6w
rscMakC10sIC/DXpC0DeTZ5FqqwP3nzlzhslH3SJR0zOC8H+3DlsKspaiUTV
45MEd1u+zW5Lfl8ph7QLeswNT48NYnnsM0MPb8NHi8OEF1czHbqkX4HQEJxl
sfmcusllnq0l1UITVmp7Tl6bZZOVOL7721c7DJzeorUB/+vO+IsCnZHigwhK
wPxSLnKzTR2t0dJeauTMMACJhXRk184iIluaYmN/GGTkisA3W7Q+oLTRHoZq
ofn8PupTCJODbWZA/jnD+hY+sP3LeT0VD63p1eoMARNOdhkUk9CB2Rziv3Gf
S0P5VFdbEm7eYlyTSBSY9mfis8ferUB05JY/vRqJqg4ClqgaKYL4EOQ4AcpG
QhgqF5TKrM6xEoFoFMNpseio0A3WGCLZRqdtxccmnL5GBE745HDTTeb7NGnp
MWwGXTow6FwECWVa93Yjxpn0GTYu3WioRYBZNatNF4z0HfRs5fCIdrXRde3X
KdTgdy8VOtLUAYu7vKnY3sLAfK2vlAFtpllV1ipaqmUQRQmf4y4uMJe1OchR
QwTtWOVY//2pIOiCHtCQ4ne2QZ9r1N/VheLYHPp9zwruLAsUOt1KsNqAxgSL
N+lW+8ecSJY9Y0XjmMcj6s1QinIXyGj0Tz+MNoSeMcWTbYwEooy/+ldVcoX/
CjtpLFes7EjhdKlx4Ke/EpIOdHK+DAUtjgRFj0FzhURqxA1ArMZkHNNEZEK3
Tblyh0fy752hlwIN4rFcSp9XaS+VQI4KoQ+aoUQtO74d315Ocf3StnipuTYi
lyxD7uMUqZRBBK0309n32StlfBe9qjt+CLkvBi4isFjdOEJgGfBqqDBo7A+T
4iD9Yv9JIX2NzYBPqZfP62RyLbwqAvp+0SbKtyI+eNayX0230OhwR/F4l1EA
7sBmJmw/P59KG0iXGGX7mfYzzFsettSVzRymnneI7x6AmsyeDK74StTm/Rgt
0EoZ5hYeD2YNJ4zsriTuJ0+JHUvrnE2kh3BhVu81WzEU7g+9ExQCDcXHwe7W
epdY6dk4IzXX2WLLzbfaSuyM52gV2tK+duGEzvfvJ9oA1omoddU4MiCJvXYn
3Kywu96MpdqiTCf8PDbZInp1lPsvZSbGSQmdJ1oseDeHw5qUnzuLuU1cFgfb
fCnES5XcwdOEj1V/EwK9AtAR8kE/yXt1G2bpkzH8SAtq9lfpRCSaDSeQklII
Y4HkH/eK/c0pJKNWQI+xOUBetNlaQ/tKS3aGXE7nP0nNw+J5b1n1jkBEu/lq
nnAA0Pd7VgbLSCBNEQcV380wNo8RFRgxOxnTKJkhD2HeD3GRYwhjJoLpJwp9
Y/ChNrODsgY1hLODa7YJsAV4AY92J75rHI1NJrUGYYGtEkjuHIm4CHUYBpK4
i56o+9UUSjogLDCmcWnqmN0miKLY5hcKVZK8a22n0sueG7Mppx5cVj7A5WqJ
912RLfQmCiI5LQHtRUywhbXCIDsrxESgXTcMrz7tevBBGav4bUEYo/blq3dM
xtpR9O5A0dv+oQHDEVyNUD3qNA3iCS1rULJx+8jCNhPMVGJewSDKCxM7c7QI
MnTlRmVfIPv6St8LxXhxyKB22xUGjmFkk2ZVrVUEj/TSxfjyqgtxgYWQOBD8
a1kF9xMjEbg9eb/JlaPKh2P27n6dFXQ4s7WKbrJ0L4VGCllBjPcVY9VXz8sw
4Fdn5x+3BueinUe67Vc3CYbARlj/DPMXFlaADUriljmxM80yeUMS3+HsTuyQ
hF8ie3apGCZi03RHgjQw0m7BxsewjvlA/O/FiMJMaz5gFadsEHiTHtRFaZoU
JdH8nNxPLiE4oe1VND2qZTqbXZyvkPHVGmgD/dD6pz2tS7VChMZ4x0N4/DgB
nDPNppZIDS6pFxdGJ+fdeCIT1W3JrPJwnWIXanwOzyR+ME03H3ayXHg7902H
6kko7lTt6XSDtbmb0GidXBMBavgfoOcskwW77gf9W8TFp5xduJTwkEUv5FMw
6XjeFBlwdwP4xyuXo36WQYqlNT005RbEZYG7y9BRbXKj6JsfVV5zVQPkoFqV
WxPQDqcU8XlV6LdfPa2cWfWd5zCFY99iW+BJ3yGXqtCQ/acVJL2psDUMNcGZ
e1Xnu2VYpNVDwqNzwv63BvSh8ICXt1fWzbVRnedksBdK0QhcXNNSqIC1j3dJ
JzaQGrxp5IZ1f059QhOB9J3HF1lBsaurPNmGDOYlUBNuIK9QCUp7RQlqlKVu
HDern8R6F0SGmiMrHw/uUF9edslEVWTt8WHTPfM1fowzsOjK4TJs7uKY8LXb
v8eodzZbgECmq19gZ2X3RdCWB6aTgFYci5sT0UXzG00zIDSepwAsNuoXpVji
y+pJa7FZMS3/RIfeJ9bffK+wlXw3OzlIY88G7bNcmKD5fEvlf3NgkIgPmyQB
1mRt27iPzJV2YtF3QXUFDLNwMIL/7wvfEFw9JTVOUaeUzYjoC1/1/YhNmEUp
n/7JXSflUfVIWnRHyY7JPgri/Tl7PgOw9aMYlGQwRZZnd9yr+OlcnbTCPyJE
QTazgQ0M/VGKqakf3UMr7Mi/FfKqOYFC31sCK2Kcse0m3T3bYGfdaef0Bsjp
VvLU+OPmbAR5PjR7+LEOkPa2wvHGkPeHk9RVmOGACER+KT4BlkJKPUrthDSC
HB0QPkZI7I7QLiXP06On5Aqa6CYMXT6yFtrzOJuF6iUtQIj7HTBSMQpjNZyq
1uDvx9/IIJij9OEHCKcapkL7f3TBZync4olaMaMHWFsCU2iI82kB5MncoefK
FjxELDBDG4r9pW3FqViGuxV4KdQ84oFTxlUawhFCg4w3HBWpMKOXU6Z3HY9O
L4RVVpJShB3Cv/Va/DDhSuMbPw3lrGZLkJU35uIZwFltWWRypcF6Kw1sTJ5V
eRZNE5jL47VbBt8xKBvDHKHi0dA77qxV5nxHWfpc/kkk1tZ+sNx/9kK4vxMt
1rNqMiTSKOdU1KN8nj/pznebsP3XNxM+v6S9Rp5ltRybNka5++pLYRwlX6q4
SDScoPeb2BBFmkMRiRW9jjtSZKv6mMOOMfinHMPJsW6a6Al8oCuNdTdiSk96
BK+3xc63SzYkoJalLjGnQ5yqBa/f9cBZMyj3VHKOkfTuDoDSnYr9xxBFsHdo
LImRasVLMD9poRZbPN7xWfqlZDdysLy+yD6yPSslYumvS4ZJuDIZ5BPrVlHA
/C/0zmfZ/qm+3S6zl/rNyeiZgFkRN2YzlcGoh6dSgc3ogMepo1Bx8WUI9bb5
dMxqWgQe8WOkPQ0GAi9IsIHzou2yfFe8xxpLrJ7Y6CIPaf1w97s+QuYB1aZy
MWA2b7XB8I71ep1ZkvodZ0AjXtLm+ZR1WmKUjH+YB1woOUh5hr5YFkOSaBnU
+vM9+v5rCuypO9yHI96bRlTTFXYYZAPhVj1PBzvgZAFMXFaLMgFLfMqDSO6x
/mUb74VVS9Eyy6vuOJXAlX0zgPI6BJic2B3CtKXP5t2/6/oHFEET2U9K+UH+
qg6ZivK3tmS05A24JNkGv3If5HZyljKvK2zesMTsujkGfsE00TSDzoJ/kAxL
7jwOB74Qr/CZnBdsf2tBgILcShnBRRdJPfoRc+QKT4FpQclRfCdTR7Jvdpi7
huP7B2yk/3/nFzuuFOFuiQDRMUpllZsSXfiEq9t4o6BbNzwRhXRCycn0h4Cw
yA29dKEU8NU7bc0MRK0aL2qhS+EllBJWZaMjBmDlHUXl9ZRu2KLwVrh0rUUz
UsoKbNNVN16Bkc1/Y16cZNF5eZTnL1DUdTqrBeLfeIjDCsayV3qkl1Q3P++b
KogBZoQjLRW2l1CpXXTB4PbdJlz6eAGgNS4EwVMPJZF1epsMI4OjGcBtY9s9
YgZ4cxJhQkJxSc5ef+WcUyrbeA8xIOShtPdkXqN3LcVZHvJ6wr/YC+B0hZ5P
/F7GSex6qRavnNTFcZnrmEDIF5WmF1C/tGzHvws2Q2VdmHOaRCNnF+laTnxR
AUb6ctMsdhwjYBb8W1TnRVSt8mQb+4X8E/IpX5o6H/z9/eK1xN6sHcY/2ygA
uIEsXarRQqqmsvU0YoByYzRMDRuavL7Tml/l7Nwklw52MuWG+V6Tto3W6B4Y
SJbJVrBDNboqPZh6leyP1kx7Cgxkm4U1ODZAEqDusjvsS4/RbNS0y8oSSLnn
NKVQUaVYeTmIIzDDTE+CqHk/lgNEXgMUJ1MTAO5EUL9whnJo4sYgibNDYKSj
EBnAPgAyQ092LglCi/VHppUqYlDiPG006f7H/SJEPbA9o/A05LiyagBBKHkZ
j8SHfNoia/TjUd3R5w9cTE/DxalsMEQ5/guIRGoD3QR8lGiV95J31xdfPd4r
4uoPO8RgiIe/gz+5HqApIDVhlLhOODly2ziUKWI7sL61UuIxdc6TFWYvXPDZ
8QYfqJZjoRyiZBH99HqpUJkJKmBrr/IDmoK8sgnF2ht0OuFNwtiEX5jDgezF
qgKqS1dP40Ymua/i4qX3p1Epi5PoKmFjI2XP+Gebxv+XGJcvBD72DrALUAi2
c8Iw3Np2j9mnKv8QEvXJe+fjY1WmbYscfZS+HwrdNjrm8Ofoz3WFz2gdNa2U
dYQx6ZqlWccyQ2O23Y3gI/3AhgtycEBDk/ql1hLqyje2XUwthunGw0c+f1v6
k6Ky0wYduFqnB4dmSiMEuDBelicZpwWQABWjiEPzH1Mny8g2VnPaqWw6ODm2
Z94gCQUQsCnTiBTfzGUb6nXWQea6dUpwM5RL/Qpgn8w7I/h5S9sxsxQ79v0S
Yknu5JcPeqljRAi7WCQXPDQRbQVTGji5gSxxVi+fQbhm73DruP84NEj2fgnH
hUvQGS3cJ4P0OMV0mk1LW8UgqPk3q32nRsiC5Ivf+sOBl+icdWArYBD78rta
a0sO/nAGq3akcqK2lmO8kc6oChcIoxbuZm3aMCxeYKEWj5lMhoj606xEAZFz
/Y8GyMpCtTWHoylKX+TyN/3QeUKqlvWtcocpe/bbwMltsMsQiPS5CfClWfR9
DSdesNB/6RhDIZwKbuL7/qsa0hRG9iLWf8YC47JONoVW7Y11WN14Vb3fz7Su
EuN91AbfLvbRnjdPHEFgKwel4rYPrrkLa84RHK8rgmKVEe77pLxrH9e/FgVF
7p2nYQGrKzpHudlK3cCPhS3McoT5UY/E/VmOP9kZsismYOlfIM1plonUnTQt
3zJqMW/9lmF1UEwPN6S/QwMUhv8oO1eb3I8/90VTHyrg8lD2UOe0UamnRmI/
JR0+tkaZEshEOfTv0BfIjTX/7nidrfh+KbLLsbdbRnRmXVfLQJFQyModdlRT
y68Lw81JwY1m2/FhvlfrcFKbjr5iJgYxN2nZNaHGZ9fRCOVOHSLFzq3+0EpX
t+y2Itj+aU25N+igs8kVCkoiB2fLU6t94OwS6JbMSuvo1RXpfXILi+r4mRCp
wuOHOW25r7YZxB3drPyjEaU5T62NABL41NHUb/7VOPt5JDsrOrPC9CrE+KiY
OoYjRSWeNZEyy5zttSjHtxWdCOdxo5V4itt/38KzbrGIq/xUVxaihKCT4foZ
L8c2p6rc1XmLWQ9DoJ9h1CTRIfMdoYu5PFT6EuNamOH5RolDji9ETayNeKPJ
NWCyLoVBRl1wM8oUe7W6EjcCDZa+7umkH/j55JhNwxXXFmA7439A3uhnssMq
1zwfiQpNOrQ4mFjzybLolP1ovuDVgQNemMuw2vzkuGz5grxCrnovXRfvmHEy
6i1MoKoe9IQwa7PMRbKidPqLxnu7yBX9TPG5vP4rk3tvCfZHpQGdkuBJJ45T
SyvMv3ug+GiQDhSbVxD0IOyvxnw1ftRmtSr+X7ReLoUw8ADrthJz/ok7ErRy
OIJ7OkrAjUUN8ruOi1rWkDQSkR4aE/OsAfJOlv4ZJTBSOD4hd4Sy8VUhcmoq
xAuzTC4KmcQMwXPdTlbsQSb3G4ltc+b6pPHVkxE7B3YawvlC5oqJR5JkAbi0
iksMVniTbWAsSy2VDqDqQUrEAekQoSXXVZzUhMLXT9At6WZJx8hcid8PBLT8
WAj/IFptlZksYHm3LaFAAzv/xiU57OvDKFG9Nc7DZlT6Vqfivf1ROS7toFIW
D87vFYABrUITsPklQDySOAJynz/VPzQ5EGhArUZUxXyknUti1ohvyo2tYHDg
/uepc1Lbfnc/XkFFUyDPmW1sGDM5kgSmbsvR68KqzJw/O3vHj48l0m+w+HbM
JxfupmAdgVloftXBEltie365RFkZgl+1+CD2kdTRlPwQofYw2fs5oCNB8TkF
m9tvSlCIhR0WxuWIG07JMKoV9e1E8EoIJwbWwIxvG+LVHuJW3CiS0n0rpYHJ
sPbXQlhyZJwRETv5v9hGZYdfdZ7Sczwed3IsmI+4D+qKE+/8ivq50xVe6DzV
nc+GUiBzoiNKMsD+ccMiuswpyx9bH8+Jc3LPF1yHNNxMRzyzeEKBqVrBPOfi
fBdYb3m3ZvfZGonDb9CXwILYBOMBu3RjWu9D4YL6m8/S3Z8Dvrc5N4f57zSk
v0S9MdLQAwVkga8W/W3UFPmgPGEiJWvHQn2Fb9lpb7xxFeLHYmc7jpaeHl7R
WmQeyMKXE/obeWPHzCp3fKMjEW6JIVfQisRQrwH+fYRfXiaCLXK4jlbr76Al
evje6QPbBSxwt+myipEGYub4mdVgP3I1smtq8CMq3YksKRVyq340+Ipfz1wy
sACxIn/1kSN3AsJ1x6Y1lTEhmOTvS/g5AkFPUJ5aM2Cigu4xBa7H69xwsrVR
ZjeuLf1x2p8SRuqSG10C+uovTumgEBgXUxJ28o+bfcNXZL61R71yn3hJX+Rg
jjMbsGuYxY1e0qr8kg7KAozSbGpEdAbad8wjVQI8JHzKFSFOIvB+QYVUidRT
uWV+r1rYkIvWDbpNJvCpsy72OqPGCyTGAuoBAKERZbTEv4+VSmNhg3N6K3Mp
2HH+yjBTfAOhfzmeDdBoxe75JN4mPES2IcCbRkk+QYnkFW6J0Dvt4AXgYdBr
kFB0Ur8r563DFgI5PCAjUO0smOes3Er4j2c6+/ajx/MlhAb39Uiti8iRSwvd
fGIeQwXHS9gd6jYiPismkghous/V4x269CY1KelsjiMBcC/zKIPIYETFwrsQ
Esz5zICixlGRpMg6nZ2KSq3zn/NBjh9mjcNazdzmhJZQVIZg+Ucjvk/EHSoJ
Uua/f//pf2tw5ZHice9pHpCEag052twNhFG4X0iMPYcazFPdtrEYpRHtbeDm
yfTongtZOcZSMsmzWg7YvW9fkdcQ6u5bS8ivV8tL+WzCNbZugv/ZpxYY60E+
JQjXwwlaflo/pgQCXPNFFkjv33M8ilrxl37x4tpeVJK49I93YDMhKsfK+Tb5
ccc1KixQZE4tHX2OhEbtHIihS/1sP5Idtd4A9czKNn/A0Fkoo91Uqa1avwHo
DF6TkDCWCorWVVbQHAFIbM/OL3BlvIaQLtHx/gcYRoFQorQIrhvpcz66O32t
Sil4nGocP4wsTN1/HSCNZIly2W9zUiFY+idsYTVIFx57Nugnj3whz8WeQ6yg
s/4wEdP/Ja3w90QxliOYdlR+HpBSAsx/xL5KiSKjKzbimEzVjP5bVBl1lkJs
hUY/nLRNyPoYHo0cO03prD3MHcS8IT75CL9bGg6DkE/iKBPiPC4OEJGp0hMi
aFrBfMkK3kXT99UO/P5IwlZC54ZGHGRSQo8Ss8K0WOnieiO+5CD9sULbL5j5
pH2GM/9IhThpavgJ+Di8L5+HbLA7u+Nep7nELQubc9CyUmbOvDZYBmkIReFY
QsqruX/B6+NA3ePDB0+AQZgPKAKs4WaaLrU5rdLmpMuRLcgdXXAs1KhlXX5U
3kU/Lv4YwwdTpU5pPZ5DssUCGthqlZREMZn9xL2/LtR858X0tPy5BfCvRgOr
K34ZEVr9U8HAA3yFqz/MJew6+eGhphX1Yni7SS/4ekuosOsRQRFLYLLHtMhh
yAsR3rBaLfdFrcwdO8xePwlTG5O2wKTN2rfe0cuc5n8ub1LC2+4zDJYOzVqG
pdA/0HbNz2ubsVnIi23Algi4NE9lNBYGTLgHvafdczdqU9pvzFx6ndurjFkk
GxtZlTrIoHUFTNAZnQHUspcyPHW6vPH2xujOquJPaQplWpaE9cIDbVkzDngu
0AsH+DFya8gnb+7j4kZGc0kR7vSLc6nnRE0eB1JyeAG456yMF2CiahLonuep
cIUDuLIP+H0UY62sznm2oSoq8IrJFc4skeClCuNrRPCJNnm/fy3ATpC3zWP5
BB0UXAXevdN9+eH3aE5Kz7BRZPd188i6gAT+j3kd68uu9Gn3878WNdK1iC6P
KawfKjggYOtPuY+9DBy/V6D2j6lI7yyNq0LcA7olINXd90nz/+h2pzNpHd7L
qi34dZ79R1/Q3fSd7uQuYL4Krrq+WyhRg5sJg3TfX5L6mv4YvgTbeK+XY/d2
hNOGCurEYuXS8pKfXxy8hNZ2JysC5VvDHVQSzHkvX/Ujb7B7UOsHPRsyJYw+
/VBGTaZ0ZuuK+oQvshGkYqzzssx20mn2b9xI1ubZFPYY1EHcl51bYR1sonWY
BbzEIXD3HCBqD52IrEx+YEzeijlE3pgwqN/e6FZKioGcadgM/FCJ/C1DGQ2D
gdCwFcP1j7pQgOd9KU8brsdyuDxUlDqoBQ5vN6P6EbbBgsD2MNIp8h33v9Ts
tubYnpamx5wqMi0m0tbktcU4fD76WUeyaRbGPPsu1OUtdyoNJFJEI5goxUNk
J2oBryICwXY5PlI6SGKQ8XU+pxhdEpSq3BhP3u6AuwEfe245+8/Jg6zKFdUN
Bg2NnUyHSkXZi5ImqawIrG9NLhJGMk+8eL9rIND0bh1+45ghdFNXMgNMeYzE
bdIlVhNYeUNiJ1YkR4Lw0tEPYNcBsjVmFwmwWlfaJQLyC5wFgkafyJqbK3PL
A4R95SO76YEbmYnjyHmTbu6XcT5WLtIXcJR5U3GsLniKQ4UO5T28ocmF8omv
CAEuAAbZ5bQBYm+o6H9Z2xrTQP76MlH+yHNwouDTRPiv32UscohedvfV6et1
dIlP25HW62BsxtK7Ul4HVKvf8zX7EWRs2SUS/fLimPWs+1tCyYehHoekde1C
O0QG8rWA+Nybcnk7QkSaZQEbImjiMk+laQUre983FBB9oajxRZPT9cAFl4GC
MCjodqSsDJjPmusOb4xVMv1293HiidqroudmQWHK0zOqiNutLNaPzDO3zLNt
BrBSk4r80On+4Il0LfeP82mwypYPAeVTiNwF1pCGPYFtyW5Sx3qWhM0HpL0p
n/u80afBCifLEAy/CRY0I6iOPeovcpKtSFO3z3X3J2aygq9buKw94mr9gPuX
Wk+Gzjp2n0WoRgUCAL9MYtavzWTAiifXqQSinGGgpAwvwvJhCoEjVlmXUcFa
7r14/uW6rcXFn2YaU8TZk1pQ7axemeQIDaVAB6PNXkiOEyrcl9UvxNL3ZbJI
14j56DXJYrO98hhcrGbEOCUC8uL3n+0c3ZKXaGFZFKLKXZljafKEn98OUj/0
Js3U9Zz6Ow2X50uoTpu1CBzYNFJCuh6wi6B8D1FjZ0fsfKEC4GlBKlg6F6Gb
coso7kWzR4BG2z8H9hA64UUy1WJkzIewbO489z0O/oGhSwsu5HOSTGRzJqdT
+ZQpMvu4qKxoJS8k5nkvPhhNE1RTCUYtkKdbhhEG9OzgAUYllnfWJSw5+qrj
p5QOU63AgAae5WsDJrafK5yE2WUabiildzlsUGiACKFdq2A1GW3IRBiFfjxn
x+bTU7GrGIs6sBWkigH4rZXj9qSDgq2IgEJnD0fRcE0phSwWWbiwtSYcl1cD
qHwgdzPpmqMuSL7I0CIlnkPlCAJZc+HfuR16hs8r1LC7bJfuKCwLvniyyuOH
va/IxdszGxqq5Sic3rBQF7KnMrjkSRVozDucHx4AEi7XiZ0XlxaT/7mGDUQb
n8tqYMXFoJvKC9IqVQD6jr9+SMjMXX/Tw8CaaB7CZQc5w03imUQNbROjQLqN
TffKNoX0iHE4SOQdyLy7yBbicCL5ylO3sf8GoDBbFd3aPDyPs5C6USAHz+o/
eBJ0OpZe2G/dzXtDOkdt3SZrhSbyqC40U96cpz+WFAlvt5CGPw5+5BnblVr6
w8Pz6vX+Fwz7P1cS8VzTZoJXveNY9A7nzpcSUZ7310dm3VSs0qKfBSaWZKgz
df8s4G3QESXROOxI/SX4nhEhVgUbK8iwTXWC1BLUe7Exq0C9vLR0JqpPmdZx
C0IQUjeANiYzrfMfEpSPxfytZ/w82CWkDsN2WKDQGJRsllqH3mNjHcvWdrDO
YPWQYayH3XhasGn0B0zSBq3hdSVHZ9Hd73dH1aZ/uYEqGNOBHEUvveV1rHa3
juSaChaNIWiy4L2KScMLRyC7RrQfUayGh98XPKp1kziNEaiWKLjxJvW4xeWv
hXg8OQlhzVyy9BBCx7dfuKbl3Ozw41gEkG4MVI9sm7dQnjnJ84r/n/w0XAry
mIkVvCfwZ/GVNEbE8x+RSynKn8adwhKKHgNasjoZV4KJf5G/Wi27C7UY78QC
MmUW23uualYj2K4kKao+ucMBzpIcuTAbBpMBI2srQqLsyavBoBVNxjTL0/wt
JbZR4a+djYw4NBtC2z9HOSApGSl9pvQQHx4QKawxD7wuriIhM7f2o7/5yZvq
XnvtHZdZmL3odvoYeNnQCHLfMyYnTbYtT+QvQs8E5D90JRljQkL6mmpWbz/E
7cG9VFX32ZAq3nAWPqdPZKhkpNQdfXPlS9B/251l4T2CXIduLezGJDZFqo6y
xj25inJZWtjvdcelLpf+TxEo9T2R9Wf53AHmg0B9CD3oiktRiHBuMWDE6nv9
MAt4U7gIUsyVm9U2AEBD8UpFhByehjN17jotSWyl42DUCp7Uiwo1LM5Y4JEX
iPi9UpwlZMr+jmTHydXuhKDqCqvgrrbyirEn4YU5tUHn8SyW8PG6HleGjpbT
cmrYuxWI3myz8kxHo7SHtXO0zaqs+HaM86WAu5iCvtjoNrf5waGwPDXKj74m
vZ5uGYBOOY8t7+c5QllySiDQAWzb6aBcnu/VDoOIskxw6nMDBqTcZFrzpUqY
gvdnUHIvFv+w/PsZK4TdGR7TDlydX6Mnoh4cEtFsjkTtH7PKaEJlHff1E8y6
X2HHB8CzqiOtWVdMImyQ7a5jQz3tf4iCqOsjxIit5XOfX6GeC4IpcDl2CwUE
82BkCtnn0qmulq01dLBVmTJN//32IJlYr1zB9WAuMq3W2RFw+TVRHMCeozyV
baac6NjWWqGR2TBH0SyM/JG35iZFUoGhunYNDnVhljEiT1TiuVWMLP7ATXqu
vNVU/w8qaUl4p3gyc0tARY0c6zcLCvpPIH5Bfosr7VuK+2Z5GS2st6ZS55oD
1IrEBIX/sSXwUgd6VAWtAGud33Lt5dluqfqACNLAPZwFBK70Kq3run0RWXae
La8d2yww7NwzHUUP+5+C6zDKid2MbAvh1LW6uKEKy4ZwGLYs0nGKOqJ9UxJX
hxMhD73um+n8BkH0eWVoKAiV3vkztnSjQncWQ6U+C45jI+7yKKiwkcEMicpV
nftE79jve6IDrlYe4J6g+8P4c9+tmm2Pf+WIYOEMjjqYBuz25O4tLSWi7wRK
2tdoAb+/eJvEfLlPG+pOmi6BpxNhESaq8a6b7XIlM060ll8i1VaE/fWW0mzs
ji1kphGAmvY276T2KVn0PNHzxjni7t4PvyYFdRp2gfJw1afQaOu8I3EGer5C
cOEIlklj3PX8AbwdYtz42Hks1dV1xn6/rPqboXB3lcAklAU9Rer6R87b4U2B
MZn65IDFyBL0EI7R4N2dTAZ6HohLp8ENXculf1Hn7TCJJdja/DhPhWaO/crS
TYJElJ/nZp506gsGCdVTgYv+PDFkwGkj740ofAZKHuMdQpU0P3HmuxifZbN6
lCPV80EkPkd6FwSiDP/z4BW5nJsxvUz8CCtUEXPXo+1/ZOQ971txvepiR0hx
FyACD48PhRtHAznFlUogSR0kKke5a2MD6tVXPKBOuobkf8rZl5BLSaQzfuXq
mIFn82WkKC5wPis31StWooqzudV0EU+BFj1SpPSnp6YxPZGzfjl0mlXf3RCu
xFzh4qskfLFW1tz6epBhdqwSVsWPkRI0qR3BS2xxTFkY7iusafCxwgJ1XUuj
BK4O0pKGIIEcG3f7MWmE9Y1RbpfXTAMCJy94Wut/AzBreKvOkRT++v2BDqBt
uHIRMwFh67NsXv8fWki7/m6s56B/FOFZElCZDny/0Q6/R8FKw1RH1Asvq140
e937H+xsLNmy9lZUHSzajPlB48Zu/oCHmOTyyUEWesreBRCNuJdvIL2HQTyA
u33/NFCgmXNjvBaT9LSsfRdFYvvzFQtxpsgeNUABNS7gumMwtxcsW6l6m3zm
0pRHBrmLGpAv4flWRVFFNDJSlYFNvw/XOM62q+XWHnu71U65cjulQIAFQu/O
gHj8wHxfqM5cnXlTEj+6iUUDzhUp43BSOPSB+Tm0EfrdvNFDM8mowwNWl05t
zD4hjdXPJ7F/c80mFA7KgXwcKfbittZVl91UXOOms1t2sr0Ius7TCInN1Aju
+AycV8e8vxzHhcA4Pf7FiCyID4XqaERXw+gx9Mga37KvoLvmn1gVont8hm52
UEuSB5dy7i2Lo/6JfdlMVAcN4FdvMBGoNqRxhB5H++Kv8fdRB6TklnsNtf+I
ySig6JMYe6M8BrEusVePOMu4PBVghvpxhUObYfYyXWcx+mOapg0fQYzTCxsZ
RSgiaMsJBo1DCj2lgsopyajv8rldZgZNobSRg9lT8tsZHuxWmtMhlhHqv953
vWfveMt1GWprx3zUQYWq8ExQZ1EhAOG11vhcWPTABtwpZTQiqf8Nr2SdB1Rv
2SLcNClbNnZ3KHNnCRXMJY8SNuNxkZrbeMjaNyZRyqC5fSI0aKiYKrt2ua68
WnIT37SaCR3+4Q7/zbQIAA1OOocQL1H++648AXSwTF9ZhH+VuHpKjzNdrewa
z7eonJog88OZ2ToSv26Bs5hLqFY0JNH/8q21iNxz6sEjlwJR/ftbNAE888D7
VMTmMJ7+Xj87ZZV0Y09yPkPABKO54uRHormDoHY+r7bBJstt8eM8PoC9gkbw
bL8jEX4Q44CUu6frA4ssxDpzo9ucBeRcUCrCp4nwLggUqlGhyaeN2S5DrXDO
fP/1AVzyK41wGKVVYlYtdcjaSXKrjHnZb79z0alZ87V10+xzPJnYzEmOCZUF
8/wIJDTST+OYrEyE96gpz114OA7ZHQUMjUwPUZzxSwVHrLHWk8EWf9vgOPeK
un46bS+oEBJlNVzDf1u0fMTURdCmuC3yZIKO1LiqmMvyAqKBbLXDlFdMXF6/
0WjymV1ReW91FjhnxBrF0kUCi5p2tG8MgeoxUOnN57PF0x/tR6ibB7nlet8b
E8iKb9luneNqhaEQKuRvzcyyBPCPjzDK+QFpUeGKVCT2YlXbtG1Cif7x6KMY
V9jWsJUGWCF9JoAe8j0s8ZrSZXyi4BHXlHJIfq39JJgJUqfNylJYjz5YbLt4
RjFe2CGc+jfO9aa3Eq5aXOdc+PQztEfA6oRuM0I/Ux+nrOAIicFWgKrlyb9S
hK6i1kLtN6G444sXpIJdcE0+jvo1OfLfys8T2mKVlpZoOmkd5CM1WH+LzGsO
fTZpTRj/mkCDu3n3Xnyx1uQ7SMJL72zMME/KHDAjEBASC99214Remm7lAbUm
e9FSNPgD9emx6tfn9wAwpKTnIH4+kIpXflBKVTN/ZuV288cizTa5j5X2gf3D
yN03tmwz9Mk6dGdJ2EgBjkPSLw4XMmnXU/FPfWj8R00Az8b7u4x4MKaZ01m7
7xZI/6vgdKtFnm0l+WUjUNHLw7G/+9WoAfQ3Uool2ftrDtu5z2JAgwX/hqMZ
EvYTh+UMB7fq8c0JmPpB4L/kEqyh3mYapeN9zI3e6Y7X2Ji9AF62uYNCCVzR
UKgwhuUh32iXfqcA9y6WFQlDY/TE0OpGoI/Uxe1Qk23PMqu0rEichJrk6M0t
qG0CBrSQTuFnw7+d/nFTPb9gEEwqDAA5KbhYx/454N1n089BnEIm7gKUhL8p
XsCAqCEf0XjoTi4dYAmM15IOoJJQP8pz+gqotkCNVqthtWs/7eXKiRnxFYSX
MNq5QpbWmMqKBCJ+jUA5L6UlJPOLqaCvaozApsKvHbcOKHn1tqjCJ57VIeud
V9M2vbtxEc99U+Z3CAQv4Udm/Y5GYMoQ4WCEqZdCNktfkN/gWe7c3R+bG5iC
wbKzIOApTgYtaAKHhlshz7+aIQRXXCjL1btuxGJLd3lKmt6741zM7ZSUqW1I
3m/YLAt7uVHWoMDS8jZ2aupZcQ5GJ23w3bZQaRk+ghpL22CnvT/3k3R3u1bH
+TQTb9q2+kdUklZZulXi8vy3K2fKwWWkz1APhyPH0G5rvlaC9JF2qvRzuVZP
yOEY7BHF6jHotIPwp45anMw7RIiyy4uxqQkicNsRqw+rZLvbP35QZaO5iDFa
4hGcQIikMHG71dXE7xzOOGvWqNR5my0aHuRNqgdz0C9YAktDDIOHVxCYmPxE
/KEAtcp6MaBqpe+HqPedQk1RVcQW5O5d6VEVD5E5AELwJdls0o/jQr+wzcu7
p/RnIA5yuZOJex/UeJYKoMEzD9rlllLN3c2NvLC+7iJvxluv5lRnghKvVKXC
lg2z5mYylkgFpax+S9uMi/ZDMRhmWza+k8/moULMJriq2YDq/Jscah6l9bjO
QFQyMNA0oxF7mgewf2Spav1tORLwECGZzuvgTtBVCFMjHnKPZ+PFUhVWSjTH
awuw5vJIj30roKXs8LB2hcIXSlsDwM9lYGjiZaWHebHvxRH/c68weTlDqHjD
si9O5EhJX96vD5ZeOXvq8MDPpJEi2NunUUELzvVgNjoU8bN7ezT/UnHc5jV8
j6pmxh3nzAw6b0Bn9WIU3pIn8oBNO/fyfkU+tQ22m4w9HStVDDwhkYP6swq+
6Gq9sWB/lyPu5gnCTqikkkxIYZvfhwtjYsrM0mNjEmlMXgJtr6P2WjzcqLpd
CkST+LEQ1FtxgLbBvmvM66zXri84XTGYWogE6yyE/24JKnJ/0AbUbTct3UWu
mJoY8rgNOPKZumZLPW2ye6/zzAU4iaNwBfNVxgtnShHPFtIFtPGq3FH9mY75
YQukXcyGXEKFITqdZ+JfJ/wSdbVLPVvmIDn241G//TeNP6TnvqUNTjLqoum9
HEjZfEo7fLwjs0Mllzj8V8T8bKOA8tUBRD62xCo2sMYvaqsrg79p8lKOcW3g
t51DrMwk1EjFWdfpCzvj2zh+cD5bDyl864JyweZ6GIm+0lGPaAbf/CBF3ee2
LYBMnB6u2lG3Lk6PV1ZciE5pZrLRojs+qZE1ZoMTV74byLLVFbGLnpYmspQo
EjtTN+2sz00TrHpOM4rWtRSMT3De0fdHWeHiMPddty8JF1JyeTg4A8vx98o1
V/5TCrB0CypiNK5915xIDfLASjiTdiRWL4laH2jZ3suTI4u816yNefdL6kNO
SvDIAu9bwH0jcR2bzmWOm1uIdcgc2aOHxRYM7+Z71ziM48yqKJo3vkF6m5aE
iw6Eph7DaY1rQgTYjpexQW2YNssQnWlXa87o4vH0ZvivgnECDckCOce7+vw9
jYDGjv0EbaKK2rXdMBIM1NwOwRnihCPVcadeuEvTpR2vX4CB7U2RuuTX+woA
v9A2Ekp46JteMNuJgu0Iv12EhtV017RJ4ZMSVtK/RKVqCbFIduj1RuwoGV2y
RJ+OqIB3EF4htOpC1E7hj0x0wMut/20DVg/EZOwBj3qgKQwDflH97NWnHToB
b6dZTbMjcp9k5aEwJrJh3p4GaYwBSdvKKQ6RjzO0islqFYMcSWCoVa1ypw+D
RNAs0CqSrEAeBi2/zvGoVTUxzLAKt7PNINos8FYPKaIP968Q4M7/2ouDQGnM
16E7Ecv98Sn6IcKS1DYI7QPZi2oY9OPcP/x8DWyS9Apf+VBs0mjAY2KTkh+e
BAUPAQeSW3u247G7c5DRS8hm3qHV3Sz4sr2Xzwps2MKPZsVy70N0xmTyg4R6
NdIo48HApuhjDBDy91iqzr0tlb1CbA48ALWqhg3wp33u7d6rhuZSpFwmJorO
vThlJtip4yjA840uLuF4JzECr4FuZJ1/AK8JC5UwTreCyGTO/vVTu/rZATmg
fk65Hgcgh8ZL65Z+AS3Qm4qWCm8IeKinAP+b/RpV3jCKvIWeb5Eefxylcdit
3bKYK2uDfVSsmm45khhqy3gtk77AXxFCKv7qyCMxamoMmmww3iKr+taFx+bF
2rgcw1WEChlTWhvJ0X8ZinssuAZpTWqa1yiqZzxPX3OGBvRSPltwRMlTjzlU
mgc2e5ydEwtHwOuym2+T2DyujiNy62/AyB30VcLwVnAR0tvYI5EgKgKkm9hG
o7m/WfkfdDEt5lQXG5U84wEJ/fZRwiZ9nLSJ6ZHAlrmv1do3bMIX+mMVQu0o
ivoYuB8T7SKA1Z0R4FaRgj2wOJnSe6nT40/1bJFMzKrLaDaMIArDtPwpYu/x
X8Z6ma6z61cFxpGHtDq75ojztnPmL102jZad+sKpb0Rc5QqIuYevkcwRb68h
b5ndklpoXrqLaOjhTsp9Sjyd5IL7vCkQkVlHlzv1o1SqbnXf2QT9ObrGHWV0
q3uChikZONuhRvTcFxo0x0udtPntKeTJqo1/ltVEPi0dkTEpCUWXf/sfc5Uw
KFhpr9LN48K/cI/cdB62GNmc31dlE0UEKrXvNt3+fY869+h81Gh5BABcpAG1
03bDkZdR+bVkORgtwOP6Yh6g+cmSpXgcfUWFlhI/PBg/ACbEp/DC5XTCcoEz
i4vhGvd03qedz1ih2ykT9OsJY0EEAV0S9IGJJdUX5njc6prW3OeoIpx8nGtQ
hOn91va9JQ2FkP/6pJbFOOSfC87cK4OYjYRMqcRoSunXcbNtHiU5qZyNgFwD
fITHooPFJvK5ENc4WHvgngxOSMj6Tip5238kcqpjuFeVdXeeQPnrkjCjcrXe
xkTkXPXCaYksy5OG0sViQBtwNbAEwl5UE5+jBmABPt78/VURcRI2paQHE//0
8spkdFiLWS/huk6TwFkVURa7UtuiAzFaiWeU3icnpene2y4lC4KDmF0WHXO3
L/95r9H2L0mPcsIDT2cmqkUtZrtO2bDuEZodIEs6na/u8XC4tOq6oX+Xlvzu
SD5ozJPG55rgj7Xt/N/svHTwuFzEgt+gujm1yARMOMriHIgHUh+wmPU2sDIT
HrvLvF7eu8h3SY4sh0NEBlopQNgkf87i+Mw07WtL7ewgQdwHe6brea6EUAGw
hG1PEbNENJRsjS6KVNvzSkfd/Nbg7PRWAx4ZpYlXqVb+Kd/9lUFClctd7Cgx
tUK9yHH3y9mvZrvksWq8WsQ+uMbPKtyBzn0SIuDm2rKXP2BKO95VN8ckh9D2
zt7S+szsJaIuEZOsgNXqJlVo5Virnrn13suxTvUpNBy9kmuRxTtWROOZ3RwG
6EuspdB9AlMQthskM/ra2FlTWtJ3dL3fMVzbAJ3egHZZHkx6PfjPM/Jw7cNW
xJrlnoLeB/U9PQvYvQD83Bc/p5BlB7vbr1eQqRV2JKNDD2tOk0zWxqNUE5uh
D/0JGMn/Vrhg1QAC5DqhcfhTz/NOkvmjqso7+qDDE7jt+qzkc0brIE1/5kS7
oM1aMHa5Uki4a6FEMVRTeL8odGRm2Xe8nqR43LbxW8lUxoqItv8viGWaZco4
AsZ2dXRevheuyAdlicP+AM2oqh9PmMw7LukPLf+ZQ7qBenxISeE44b1kIbsK
c1knsamkYDSZz5RDZfd8cvbu0ycw7EYreToKY/UFCYisLRQgc1mqWTPUCkFz
8E5n9EEWYG2+HdsnCrmk0SUi+ncaOeCf8HCSvlE0E/QXEr62UF70qeci/E6+
gEHaWFvdVwg/3cfTvkE2qRSsOOSx0zP0HXHj6TMgWYYhqgfu9YoymMm0Yd9q
fBcVfEVtl2zTuQePI2Zgcm6hkVFFusi/PbY30aReOiODjLZI/tW8bYIqE0uO
ihW8BPOhcjRbAMhTmEwpGa00uWYjrMfh5Pm0bmUgxMFQB7IgKbXjCUL2aNvA
SfHm1u/WtH+w9hOxPxd2hkMg42taCPl+4SZJ8M/uuz9K1JHwB7Ksbk5RQbE4
3TlK1QcUGfifkGQ67De7QUr0JFkgQ61EyEpSqonJu/GaOiec2Gur7yig2I9h
ZiQlntVbKQ2moJK8pspdPWeXz/cVJITPpEZHoles0HtGL7XnBlixPsTKVoIr
geQxNbajlfWnrT/eO7dWxqeRVqfN8WtR2rS2YD/lcskCm7Q/xxstqfKGLnV+
ZY2puFOo5he9yxZpAqpfFWlfb+9UrKA4abrV/Bb417vcAKgeHez+a6VgvBQl
QXoxgArLdDVe6gW6AEJHQBPQkQQXXKxp36QqQg8dLa0q3PpsPWhlZxvwmdo4
SHPQq/uesedHtP8u9/xELl4/50fi1JA/+W9dnIflEgUgbht5kEK8xdjAPcbX
4Vi4ukjvcfIvEIGkgIMEVqgPcNRUFfg0mCLuDMnv/kHvIZLkpRZ6kAD0C42N
O0OPid+Tm0vxfgKCMr52gZFb8D9p3tz6akHRz2LzcNfxSBV0FxuHpC+YiPuj
DSvIXf8yBj/XrTLgoW5V2iPl0zIPQ2IMUwvR9YWzdqi1g65245nOY/WW6f0p
IuRrL5IMcZOh8l5Kxi67HZ/Ip/XziEHIo5pgFhsINtOAJqkfBCoEWIE7diGd
QvEQvIv7vlmk2JfGfAnpTlu7EO1y9R05rq+vU7ELxY1lpTaQlPVgsgD08N8i
01PHY3l/Fq//kZBHPp7NGXA+Yw+ak8tjE4H0SSJ6km5K/eNCgSAOdnpFdjgq
bBITdBd7dxmHVD5xGXolD73TuIvivSe9VCf08Dbmz0eHKQB7YDDHeHANZYHZ
BWQ0yKQhuQHg+zVjPyuCoMYZfWlgOt1bESFI1sF28gEZzzaJel39ktHHGwiy
OplrMYvGiA8wXyoTIOWtVbRTPxhBAkJeeqG+etVeC2jFqX35UyrK0s4FLjzJ
Y1QcFh2HsRdoWBEmwPD5wiUcMbbOF47nANGqe3+qwfVE1WjrnsjcD1rZk+7x
FFSy1F+Al/1VzScXjtbrpyC7PmK3uuaY2DBEr9aZzjW7dmg371t/x/tbHpMW
pID8Bw/816NSez6tzEY/FhjfwH3zrv5eM1yI0u13agfD8ha5WdJBYgzuMu3d
feegZxIwzKuVT5owRg75Gvx+ihA3g337MmorG21XLkOTfGx6xlxxTr1sDXE6
Hei670X1zfgcnVQwrI5J2HoHiIJoElUD0eHkGSOPSBtdk7CgTzYrLt/JBfGi
Nl5iuY19OZGZO/q8sU26UwnW/K+DmGCcYxbgDoAH5a1g7/jtOewTLchqZPhj
386htiqijVJjvOAmuOYQn75IbTRLbpHZpfZnXZYojgXHi5uj/VU3qquy/3YF
WIuOaD/d8CTh2Vt/PsAE5ANIGU4DuZ7hR1v0ulAROaYBBQOr3lGZgwwmoXKZ
Ob+6jcA8cWuv1TvpjDINdgWJZzDQB0eMDKZ51228J1GxXs9vrf7O23xAPyTL
4wCsP6quqRUd/UI86qeMhlSVmz1O4moLVKlDI9LuA4dC2ECOHZjcc+PkHVg1
kyrn4D8HeQb0ujRSys9Ugc5FmQfdJgS3ksfXY5vLIgdntSsjudkfi1HEXVQm
EoaR7YKiifzATDHQy8F/7p1iWmp7OHl1vZ+P5Ed3Jna+IX6NJ3Sm7yt3Uaec
R58qbzfa5rZqMCEUSm5pS6G+jJwPETYl+mrB6KU3Xb8n5BnylbwJCYZ3UT2D
rVAXpWwPuPUiFIDrHZUzGdQRQHQumiNz1M6+ljqoEFHjZq6Ej2TVayyu9Ek9
q4jGoR8C4hC2LOfuYjhTwcfdFsNVvnEAT9B74+Rqjyx/mNeLzMqXC1N1je8/
ZQMk/CexyvQZVNY6Od5u6hIE0mzxJ7JZkzTdPPNNGLS9jSOHP+rQOEVa2l+o
V0y98QyNT1lpIDFh/ULRKY5UDjC35gi5/xT6TFP2EtegM7wS9D1Qm+nxW5Ng
rL3IxOgCARpw/giCH+vpEZT0Udao95CmvdUO6LGUbgJXQGZk+4bnjpg8bqpS
CBW0fkSHAGoYMJ/FVl9w2p4//mMiWjOZ8dgJlRP9p9bOE0WAJD2FKOxgJfE/
GbUi3Wi/epIiL5Bs9Plerzqdu9SgXkfM/+YMB/b01wcqcH908AOhNHXfTBTl
lABd8/XfNyIZFzbIQmsIqyf9VI8hsDMNtl9uYPK5uDMzPfQmM01Vag3E3MrQ
ojIILu3l5YJKgkBqY+LnN7IOJxP6By4j5uyiieCOD7mAHfVg+iEkZuN9yzZL
lwhHtYLunb6S1nEloJFS8/z88cZPNsXXlW6R/MuzEOreHHiKTB7ULcWl1uJS
NZNMYM8YZy4ovSrC5xFpN1EO9jPA/+3fTCA1OstfouQ6hUmdmGOc0GBwUnlw
oxgrpiOZc6zVy6cvNeNmmnaS1PaQgau1sOlFIqTKDxaRXfHYm9TF/frR6S8Y
VOg1hWwuMARvEFj+pYRA5wGlK2wYHqOQPtz51tYTBEzy13LcsNg0Y1wCZl2L
bTa48Pjjea+WpCSl/KoZJkl7D1AtHGF4WR39/RT0ENMTgdZBtbmF74VGwvlu
uYJIOIpwYVWlAZQFSsDxhdr6PRGCWkbHSHbREzEBwMGB3N0UbWwVJ1N0FsCF
CCZufbI/AydnrVpOC1YnMuGEyAwBkoIqNk4ehOSDOJtnLP79ag4kZMls0NGb
BO5OTLdIHY1SkkMJg/oHd5NXeWzqp1JpP4nSAJ9liaP+cVYS0nBb80b680GI
nz+VBg50NteV2eqN4XrRhEVO7W2M4eL1xczwdJb/NmFeYFe3pzdre3vzDjc8
TYE3WrjeCdXmoJ5E1MAxMqXoNU/+G62AxbenqUv9/Pmw5BEZpu50Vs8R3RWb
D7OPvnVQhhpdmTbWXwR6OR0kj0qAxMo93k8stCXJXc9vCkHe/A2rPVhQEzyy
21OH6Xg62FLe4FC/xWTNNizTax98IGrAsUEsJugwO34pvcydxllytIDkWiht
18TiVBfSUreduoQFVKsRrD69J8f6Gb1y5FFeGX0qfEo2gK31mCJg2gwc7STR
mqRMNAbrl7eIjhXnibcmGiH3BN2SJa15hCQjzwuTjpNKsNi0e6+Rhx+L1/Q8
ItMG7ZiI7GURw1uiqZ3asJ/OHTEWzCjOU6JcA2DBPo2wN12M1j996zO9zjvX
NaebjYkbMoTnDbogyVUMQuRqK6joZzWGzV+sb7jb54J55EYLD2pHA7hlQL9u
QPv71EdjA03Rhe3MDUr/q+YWOmVBQFLOm7SfJ6S6KR5i3irAPCjdoKSXo3f/
DQkKeSECamNbNj0scQnqWlX5FV++ifvzlw5Utg1uOstZ8ji+tN/DRkIwgUCH
y4c6fPy2FpKDgYaVN0HHpdIo8dl1QwuR1s7cnCHZXGgmzDCYC13mIoYr0U7A
ereV4dayz7udUYep7LiEc8S2Gsb2ZDdzggEecPXzbwXi4FsrJaHdXteHV6G0
4Bry+xss67whrbRfjt2dPmkUQd79iS8JKd2hTK61ithLpsEvdvegGwyW8RMT
bQx6yXd2pfKPBvzj/EojnUVgHEI9SC8uBn6BfxjQvraA5HgCCFxB+Yr16+Zm
1Tq2gETuaGjlFHO1ctMfjvRgX1BHMf80Ghp+VCCszo4n7r/wTgsiYw4YFux1
SZby//WPQ+9hyFqOJukttbo5RQWhYN0EEwHAsAHoXimq289zDkLzoLZLMhSK
kuc72T6trDrykn/ZUSFj6d9KMqLGjqLRVVB7fs5E411+4BzeFK4j8WDEowlx
tSsiFhoH2oAzVZ59Ll+v0ddtKR79hu0gnyAEjG0yFNdN5JBk+xDzffe6NUd/
pg/ko4ThjWNTGZU0KqO7BKVHKnnu5aA73cxAhPkRWWRfQ9DZ52O6CKbK9fP4
156SGdf9Bs1KC8j4i7ZDMHE6V1Q/MQhx9ZwdEPTgek38sdqYVOkG/FwJxxpV
kKyr6t2DP4Iyl3g7xbbw/uQZG7H00rFPlZQtUlymWZne9oRCgzOxbUGis2eu
xlbP3MCQpdqRfIRFtEdZs/K13RY8hT+mzBnptzoFFhN1jpRO8zjLs4ulsJfR
tFtknw+i8/nO1TYJuDZ8oUu3rThdPVkgufDH/f8Ikr7Gz0PCyHQBWPWCNBMl
iUedw6qTr/EyyiMn4SI4TnmRpaEp4ClQDd8pCmFKWOg9j67lo958l2qMM30C
sk/mPXTwGT40OWI854lGMI4qlSDO/9ZL7//e6dR5IrE5U7awVvVjO5sbHi1Q
2FAGgrfhiPNS3HnortFRFyAtjQDVpc8nMqsXDu/82sl9lDVqBv03x/ShcU3o
Z6YkdISGpKH/N/n38SjI3Sw/uLD9eD2j2ksLxTMSsMBtgfXyBC/H3fWKEg5G
11UJ5W9WnlzMdI2XqHrGzlCZuhjXyJnm+R212gXcRV9Cm/fGkIZnV4KrnLWY
CJlvqtOFYlNppictL5QsLcGy37sSCpBf9v9uTnrsN1VdI3kkDEyprQrYgfk2
qmViUF8ipjnQnAcehqrVKvebhEV457feAfH6F+Evj5+2Slty0Nk5BXCVgFzG
kELMRZZGTJ3n4WQfGSDz++fG7i85Bo/kIRVsQgZVzMSMNV/5Pw3RA6N64XBC
mO3BbuviOK1kQs6EIeX0mlJHK8IG4363OhxoWgPidXmknBsLjlTyfoB7/reB
1qiEZMQRh/ZNXoS0Nfol9H34pftvORBm9JS6pIExOrPBV4pj+b6rARBXIsrC
XvOiONS1AYzVJ7tycAFtbASsGpZLeX+V5bnPlj1OEEw2cgEeAbpd5sQdKTX/
ZCB4rFEoNdlnzS1MZSXPdFhtHsTrDptbu8T3txCWXBJr4aSfdEjYu0yEPo3j
F8DWjj0pJsWYFvnlPFggle5htV3e7bqRTHXmlIziO2fCi2dTU7tT7L09oDIj
NPpEAKBqXrwvqkLZVF+ztnehdXaCnmG0PfwLAr4ZeDg9eZz2kj6mCiSdlubb
BCQJ9I3DUwPYEue1nEmqKvNphQOLbwUpKnXZTxFYuYBHq4FJFZXquLX/zJKv
CIbi8NAG7X3hD9sdaaIeMax2nwbJZI3dj0ALwaA6ss6TBnODGtX47oeFFdbp
ZTCHeAYOXE9D+U2PTk055T0mIbBT7cjVsBY0IDaUU9xerH2xw5RP0Q46k7Oh
aHLxUJ1NK7gtPtFP3Eurl0lyJlG2dMwgtObOtuYnvLdjmtkQLhOlqteGB6it
zh+aPrNepwIblJ2V47p9jxYp2O2xo5GTrbNEH2z6meheap2D84nJNQy46oRF
hQE2o5gZnoqNGjNxQKOv8yUsBzGrGPuMbebmU+pqSaazvT36AT6tlhGLiDa4
KZ38xlR/YsznmCNVXQfC8/nr/ITQO4Bs+aUKoDK1/WRb7v8+fv2nLYCQ0SOu
B1bi6MKCOY/Zc2uOt/CluthZ/dB8B7igwyjldLD/lJwyO+Pa2VfFud8p7qEQ
YR69XJRRvL5MfQpiR3kVL3nnXmbX95Vdw1fOpxrOBHpgSPCZ3i5mHah/3ZyE
UZ3zb7UJpTyd6DIESu8CbPtG9zbs5l7RitWPdL7BTRTkrPWIntew0+MoAe3S
4tce/+jVSrOfAtAdHkA5jObP6WB6GbYA0PDkXAKLOhumU9oL8r4hAKnASMrf
DrQYSN93gGDhQtEhFXHnixxL8Lhp5UDhLdV3Ql7/XslZrVXvoDs/i7oeqfVE
rpNnnvjkJFO0koWszMrkJ/akQlwNBsdHpWJRM27n7K48jkQau4kqdR4rfuPl
84xOvCnIjvS87ipFrm7qKqGSMSrwSm/XcM5oiWaEYdbz7WPaIZ4wBPk1T9So
jFFW+3PugVuuAiB3CxTJHitzKEyB3d6t3jlgANUYxeZTIIIhPEgGzBt8tq8s
DEYngrJy6KCUrgUVCeKBnKnhWQ0hlPJWzsKA3e3WTl9/D+Sf+db0ZyuNjtu5
5zhJUUpxJtGrdpk3n1Cs0SF0VCY9U0Jogt+XljynYShdLOP8n85vcXK7tb+v
FpTDqoJ19n68J03TlH72RhNHGugZCkXoxLBhWM+10np6yEEYw5xyMkHMeYng
kajAUXTGZdBtsNgxfhUGQT16DiQ1xkTgAYXvQUtp3Cp7OskSPBYZtxUHwB8N
UqTHv+7zW/ZnoJUDA+02vFMGmyh/qq0M/14PXjY+cehrY5dUPA9huT1im13y
N+wNh254wZ9bBRUXoxz1av3lU2yhwzpn19O4ZUG7erx7YfvjMLRqjb8DWMaI
5+lvcIFcd13mWIy0V1kx5zqqFGrhGdRjYnDwDDhkR9OItRpof+pv7Jwg9B1F
pN2s0M73PPzhCtP2zhkNNGZyPP6SoFaam4iHlYtM/oEFykhCAdPEGvPKfeWC
FLH0RLZsdGmRgqI4jiqZnMLkLu5gxAhAr1YblOrWIeSUiFFVdxcdLgn6zrp6
dARlSD1dm5x9hYOTkPnSFnNVbxfw43YdbkT5XLLj3/Pe7vvmWtOcx1Yygvxs
IHOCUxf3rUobrPTxhHBQp2O4z6fleRxvvEq8hlUqfucnf5Pq1NntKf1ooLYS
gGdLhmjjG6Un2f3RZC1dtnTxx7leX3EvOSwLW2z8kqj541iarqGilwIoaB02
dz4LL1iyFquRsUJ/VjFe51qRCQadBtax5cir2+5H2nR4j4j6iClQLgPVsl5X
224SzqaezNrIctgfSHyxBrLur7DDuZ84pmZqyLT9wUQFXHyenDAbSF2vqKo7
jkcSjzUQ6zwQDhwkPvvaWjNf25f1EtiCSyvATXK5T1rBanWGQp48fjGF81G7
kiK3HvGsaduye1QGIX3TS8Mn36nDNExJJ9iocUeYokTpT/SQ4FHbfCK5upRm
nIyK8F14rJwVPjAk2TKCzgEWdsmv3sRVCcgiWy4Jzv8fBTsyaa96gcTzg+5e
BoFtdvkCBLHX/8MJSfhqMmRIKJUnVqHkawGpu5UgxLSmBwY9g15Mc1oTxOM+
Syc4YVwoEgrzEuYTiM+iUE1kShpbhNHw3syH86CagVQENj5u2VBsXJp7pcH+
RcFkfkWMhBDIajedIvDCbQ5ffXxweFuWC59/pcpHoTo1PRBpLLoXDWCSLWha
HzY5Qzim/B+YV3ACl8gEowdf5kvz/KlvQp0OW6y/FJgJsS9K4z4ns7VgXggZ
kTfMGTbV0D7u91V9LZxRVagPhvmzXxHx42tygR2ybWZos69b0ppap38AE3cl
sHldsHiDNxvtq2h65HKhV6kle/qQEXloL44Y9vlz3LSR1lrEKvhM/uk/sdNX
KjMR24igaiyuzhPAudrDcFJifJ0E+6Q3exM/agD2l1+hkoQ2339wVNqMmNm+
YCrCa4MLD84qU7LfB1yOOEQs7dYQtvVOIKUoOLTeH5DGsludaTMN3emE8KRE
vBGzbjmW24eU0XQMsF4mFgJwe2RHfg38YH6bJuTJab74EhBlIWV8uBp7eU8n
nB/gWHkvwtexNmKPKcSeKHO/8hpcpXz87FX0hd3GIR+016cTW1+/lv7AtKPh
mkfG3/fVkzPVPVdS3HYxGRzPgn+MXRBdyPG6nqQBDK2ROrTHIcDnj/SRw+6y
OilLaixVSqY4LKKzVU2RrHZjehXJGKLxC8YvXp3c+nJ2pC7oPm314n42HN43
xR6kxhZel9Iox0+q8TH3TyJ3uRo4oeOP5wOcMCIdSGeB06aBS3NJnvgXsIkA
sWtK4HVvPyww4srASicyJ6aHmzMAZNd7HpM7uHRBCntGQ0jncninsuazmZMx
gL6eLbaSIM+J/g0Vu9Pw+S76bdiLNBbUlFxa9uH+5rxsqefWgvjG4DL32r3E
sF7CwcfZcQjVNfaimuLTSgZd5auXGjHs5HpWk9Dpej3CsblZsYM1giTP2JFK
6EhnupW8w5B0F0Km5DPgj9F16s90JKX0xmSzCLhslKLDhf0fzCLEWOcnV9gk
IqgFs53yn+EI+3M+g1K9UuKWQcrJsRC63ML4fe0r3rF4/zEuudiYvajFSLcd
BTMg+xSHe3mi4BWxdeRRT57bfY5hoO2rP+ceRbwIUN1xtEq/HYT/3GdQK3Yh
2Gq9dVMVfd9m0qnR+QDbdiJM8+TpU8dZBfM2NJP/eSQUo3+Ft0ZTPAD+8LiF
CHDKZBw6FIBg7kX1KgSVcBCMG0B/HtfCIyG/UXlULpD9XGmVYph3if2gQn2Y
j8v3sHIw0yyKwCv/aRHykH5VnhqayzIwBnWkw3hJJ59NBYagWs5AGUHJjHbT
MIFtBDn6HBQxxUR4vNJN1krPWy9lvLd498dLBh5Q2islfHei6tYC20tUPv5N
jX5R7vvDC+AMgDH1gjT3q1qQ5ETmTqHmienuGfq397GWA44sqKqPgRZgaSR0
BOAKNIN12421bti1fIYUSOhKgtISG4d+BHI8oKN9+nrjTpvdVUj/JUBStn0M
tFUsj8HOEirXs51XIHgVe4LnI+5rtIf7iQKUtwPgfgAdJtQQZF7nAcMPR9ds
Os96DptYxGsldha/CKYsGtiaYcgRordb6cNV/0gQvVlZKD/0363fiB8DWt4p
dppahyn+jiT80FjoWr0U0fCdsCYu8S61oCNWbtYLygqFU2D3OT/a40fi3ot2
645gNkfhT/vWPCS5sBAiI132hi4cSuyv/cmRS+eJLBeApS2GSsoiXwR7cntc
0vE0ZdDSDHYEtmpYpzcgVXhTtrGh+l5q/m2Jy+o/APySbYzjPx7kqRmD9vb+
ICwom/Y4r2gaaaPsyj18MgbJ6wOJRxEM7ycnDlIsnwptzP7nmM7ejX4UTBFv
jCKdteDXWnxFfr2W8fJ0HUUy0821bsW5bKsdBnv3P7FIBoJToMozd9ES9Ohs
iL8iyCkCN1SzfljpNkXalRY+Qzm7kuOLb7WGZoNb3eKoCuH4VnFLfO6rsCfy
kLTeG92fKIojBLxs3WFYLnD9iMPlJf+Ae2+4gaIV+TlOTh6Gjj8MsmKAgUbF
pf1KAgJgkMXFJqOLdzQQPvE13jph8E3WCPiESR7tWd2qqAyBQA0qokAWVGaa
krivJNTHGbJnpNpyUc+MCLCAtcdRAR+xB7vuiRUPiUnHEqdQ5xsrByu2EdaM
3S3pB5pKlTY640v3Gpcl/DTb+kx0z1eusX96GGk0QA0nKrGFMup1ZHwOsVyd
30ivx1V6EPSbai+0wu+w89WPACGAA8c/rx6g8ieNzSX5ptbY6ib1K1d48hBM
DonTNFJZGcB6sTxG5J5KoNLo2yBmT0DXhM5j9y3v0N8Siv/ByZpjfbqY4XxT
WY0tvvgkihZnDxqFi+nNTxH+8cxZF3RPOFepJPNbrVXCoeodF3cNkRAF1L84
Z00k/hX3CsbO8gyUxR15+wseevcHloKyrmrAQIizLdGE2JZLqKbkvHuWhLbH
J/144pQiSgNtZJf0ZYj4QJyRKPCU66ai2QhVAalY2JCHzYbAMTERHrJb3k6z
R0VvbxMzzxF3/RcrK1fuwuEZfxVLeC5G/hiyxuXLPe5mRWn1xjUDl+Cq2SlE
x5cfrZATqDUF4tetB7XCg0Y+bJDOC11i/bvXWBvYgRiPCzguK7OoXFFpI5+H
bckDiiDKRX72BqijBGvkPiZcDPGU/EqU2+rNP4q+5kXpEP4/eFEPlZUNNyek
Nmx8pviz1dhea0ShWWu3Ky8aO7EshSGKb7ImN8N/95JLZGHyvOVlUgl8SakM
vuT3deWpBaCFuEs1K9aM0H9Whi6ecrxGInlZVQikUrThNRg8TwLI6NLRp+qA
zSLzWO0gK4wVw0aSPv9f/z90hvPqjZ6zJ82xr9p1eX0B7AONG6QlOjpfzvUi
l8/P5DmCMi5to5a7WzlRAfbnJRAUaDlykrFS5AD992w+4PEXDlREqj1XjZK3
SqvmDzlrDtLlMw2vN2egCPV8s5TfmVeK72cD26hGfOO1C3XzhOL5B3UpfHKo
kFq5XkrjihNJeSPCrZw/ckKMQMgPLmrmucfjgw+KQL7KbHHgWJWyNkpoAumW
/5r/tDFywX5dmubR37+0zPeyOY7u70FPj+sBkIHJAhhhmmeZExvF9j1pGaPn
JgzmOrJSEMCEVRLNjvuuT9C+xySXYqUOIwm/VPWs6nX/scxtSj1X8u3cNgnu
APvPsHcGKXmqi3BTVelpHkN19f/q2sTzCt6vf9dZD4RqKM9zd/+IS6J98yXf
HWTbuXd8ycc0w5pVc3xPTJ1I9VAH9yDHS5vdLxH4osQY5BaOZaqzbiEdh+AO
VL5akUE+7Bd5+QifpJYW6dwmkN+NJQtjfY8wRzBFDN7yE3HyDtNpz7or2pvr
BZ/cran8n3bgdlzsW/nPYIUwdbniN1bz5SPV0jAzxW9QwnMmeAtcnm+pzHw9
16fg9YK/+l2uIJT9A5zgpDzVIhvil6LXnT2W0g0Lh1jyZftQ8N4Taz9+e85l
wBSZyCO6g8xshrVyBqxm9cxbIC6BOE6UnvqzD6NR4lJFqNGNvDa7KvIOTnGJ
ZcaGlvjIuPpqn6FU3QzjB9wywg5SnztCmS+NSZ3QXNERWzYCZ9hs3D5ScCVs
VfQ9uB2tlylGvXW57+88kvh08GKoCseaTbqv99yvVIXSFUcyBrrxESUWpuxp
eaRQN/f5nl05dPyzSP/tyOdP7CdIXWVFVTpro8LyMOW4OQyrbqKa83jaaHJf
zkdN0or1cteMPMZK/a2l0V+SbFvFgvmtlVzdgxjdtCTZo9CipXfCPtuamlz4
GCE20x2XKeXXFGRu1YMe0j+NPIRwciSVtulgJJ3LvrmeGwXAc6A9Ev2RQeDh
0pcFcz43r2b83srCvU/WEfcx53pQ1AlEzqvamT6aA45v6xRxHjABXAoesiTE
fyMCrFxX7cOQ3R6F56sT3UhzoN1dfo8nZxi3okFihll2axIF/oi+xMSNa6Wh
UxCS+szvLKAB3qCAEVe1upARCY3JYUkLn+g+f2sfoWyqunnaqDCkfAWlPO4i
A4S5unF8uldWzdwaUZJZNuSWas7BdJfVfReHX0w6GWypxYHudOGjJBBe04QF
5MuAIT9Y/MkQOGYvataRKxHmIR7VcxcbEhQGizDUaHfpX72Y/Nrlx508rzyW
+dwb4ANYcpUaDMnQMtLR7eaIEfQ9EqmLXB5ZiYq10Gr33j/oZJgUnVTeT1Ys
nZNmUeaO7wvk0b7Vw6fq+Q291K1FMEcKxLSbHh7jCQ6uMY0azArkhBNexi0i
sfi3YBfJ1QUFZVdDqI7M18WAqVn3ZUiyeRLf2ska6SnO0VQK1SSCnB6N8Fpf
n7ESqEoU8Uk8ufPxTP5civkr33cqA/+Gz8FfhueH1Q7iqGdr/jybFyMH7MRh
4M5ie6WZWMqYj4GJhO78rM9Uy+HUTY+cGMRV8PvLcZnXQ8nHJ+5IA+DcvKI9
D5b1ngViHgED7iCM73pV1enAlO2nHm1+PjIWEbXbZDXI2P+lX9sDDzmTNW4W
KL5j9pgugjPnNrF7L+MxOQPn6DS3AV4/IDyIFLvrbFN8sBfM3JmEFOGZLHny
duG+3e2MRB/4773JX9NC/9f/291xldmUfjATuy1dGmawauM6eBLaBKOH2bOm
Su0fPemYP2Fgmoj1pWjGq+aIFC068JkCUaHNATFKEAfsBB17jF9KQ07jYHTS
xFm14+50Gm+BDKmpe4aCXndSdAF830dcvVU0Cax2ArAW8zb38LAm0k1CE7sm
r2WfC13enncZqusICP1P5hapTTxQwOjiPpxPJMOWVGzZVFs3YZbT64LrfOn+
FtDHlhFWs4SBdmMvICuG67LmqASw9jUDX5/WXtvh8eZ4nCMsvkOciGmuBE/E
8pVQMqNdwiP5P4kX4/a5mE06Lcq5eO2wld3ZoNIDAXXkHuen+kkxX5Cva2Lm
ClAd75Wq0ZI9PkSWE2cWftjDS9wzTlGGrOG+4kT17SBzGvFmidVzTxejA61a
TyzRTkT1m1igNoLG5L08xPU9mHuiJKEGIL8CxgC94Mu4120VjqR7//gIg9UL
TqTYuF6tKqUsZ8ZOsMRd6IGUW4LGvSXpkuz7RC0yNiLIhOLVMKll2dd5WeBr
gND/eYwbJFMvEC6ikx4BPb/UoS1dNdNYKdGdMxDtumLekCa1ibyBsLB6DLEP
Qo8XNw89/KpA2TqGMdIsEpaihyzdPjymrd0PGaEzI1S3tHiOs2b6bHsgvH/M
5hS5ND0Pwelrv18hues8oG12hn0eLtRgY2xSKToiUimt8pdlCv2w3EYQWbV6
igjMHPiz97z2Yjg4fsQpuJw8FUsK3b+V2p+iFs0DvrErnA/YUocl2kwxhjPg
eKS62FXp9XkCdY8QT8O4CmJVJNZ1oOxj6EIvuve9Thhbgeg6SnNHEgbZsWVF
lb/Bq5LTVaC6oGTiRa+wWjhzd602ccR2Ot9AOwPlt+EAa4eeW7xWBSCS0TB6
jEXYHZTU5UXoPGWnwir9eDd5yPrX1d8g7rqQwrRcuWnAWQh1qzwlREcX6MIn
boY0+MM9FORwe9SEnOogZXqNMfEIEpxUevqIrNxjYvJxfLLuomaUk/8YOZuT
NCb0bdY3dvj54giTAuizs5EXXNV+/uFAb7FSQbua+NAqVegUiW1pzK2FHbIn
2VluVNG66viyGYvi/+kFYDl81KnHSTwnxBtXteX6mcqEYr2BIE3gcpwxHhJR
H4Mokfcfc4ZosfWORbN5S2IzMah12cAiqpY81VazLpcSk3wWQVATJbRCl1rs
2jZ6630mBcn31v1cf8acxAVbxgZd1QYrmr5GwidvwLh1xDhNa+iD0D4dNddk
h73jjb2nH+yY2H6AC57sWjqOCZAaFeZLK+d/SCkI0t5pO0t+i/61Z1PR7One
v+Vwnhe4Kgptcmk8J7TTVSzuJHnOANJDwnQ/MuH+iW+t9opxzoV+M2iCxMFO
bElNaOOlR+hlt1rwOUKgAfr6/BsFR8QZlyzSqTFG8NXGPytQyIe+6y0E+T2B
vczn9M10pqIur5dfW0qtT3HWAOlqW1tw7T9q3c5x2FHA/hOJlnG/cP5OYrwe
gu3t05dK6JaO1w71CM+ulZ00sv2iU62us9WY9QKu7wd3fphGRlMFnZ6MMGhy
qthCq7yhCEPjKBXFF0Rbprk/DgaYGlanoO9AEZ8eMK5AGWjDo1PpMI5EPpxH
OIxKyLFBS+1eOqYNFyntrW4C10KoaVmDw9zQ7TtyIGJdAgvZ3b/M+bLXAJh4
rHDDP0kCl1AygHWAsj7ABD0Xng5Nfzt8v6dO5sIuw2nvKABSZ+ei+jgmoRlT
AJBGblwz04+yJIzkYM8ly6fZ2rxLsvJx2Momz4GD/thvRmguA4o1Kct1sVxM
24C0XpXgXhbNhToXzDK+6Tr9n+nB6VohRmn++vpOO9tzuv4kZznpqtmMOBwB
BBWPw2ICxWFV71AXf/YHxuLYYzERbr4NfNtkzy05g+kvwwauJAFbmuTwYyBL
G+dbb+YBWX1oz2U+gTZrtR660sSXD1szihcyZIsJkLij21WBF+/8lIpaHkxx
3mscgjZobGXQDIuHk5uLhUB/f9inH9+0/xnmv3jF3nL5OIGCojuJmZodeLun
YSIB6IcEJljG/ar3cpLXYotjh/X+pQ/JJ/4GymN6MD1G1MIqu6IbDydBiDBB
BwRkwoRwGpwVPuxJCPpbCtskr8WA8QqauaUYRDrk0EITOC7+63qZJqNHWcu5
pN+4D9g9d0uhr1vk4RIS7b1vXejCRW9Z+dBXHerq8In/ejZrvdlobHtkaaVC
+5IKCxr3zjTcZtfjl5G2hTGXux4snV5VhcnAhI6jEmNLRYRUHjV4RYGQuKJh
FUe1C5wlr5GXIW6r3RHdgRsKWz2QlRkQgTWohVYBO57t9hYJykQi6kGMRE+6
c9YrcMxrUP73SHFvuRgAgrj4E/U5uA8gMx49/EvCLV1LLoAlj0gsW8+u5k4U
+76avv43ZTOy/oIvsfL/HmoTTkEAAkDWYkma1iyEw0HNeKZUG+7ctTXu3Hit
S8tsfSQ9fwtg5Dbrwuyx0DOctn4J1WqzKnLoOaJ6AcrursR8X0+t5IurtBlC
DXwGkNYOP3Pgg1t1lnGZ4l0gXEW5wV5at/J93PUT7qcBY7ZEDK8kjvygfKTb
P07ZKwxtyNEzwKd/zIkj3bKfAJtHy4zuw9zGfM8mU2KFJZ5p0+pgPIIPUfk5
XLHAqC3UmktvFvgHIyaspL1m8eHwN52v/yqTyq/CNTbxHWHO3A5o2M9v4+4c
5Byd9dC5HLFJpYvp58/BD0IrFMJeVl9TL3PnwY8ucz/Ubx/iXMQQVk6MbmOh
jwoL3lV0wChLr9RJs8aGcwDQvOnscvHcsRc/n7racsHXynJB5OCwzZoJcWBh
mB6tmwx6004i4Fo6gGEesj8feFFswtWxgQdgVAXU7ulYUoLUME8VK78oVE4U
aXaYgB/z2ZaFCSL3fklhtmkXWlBCeADcjEMCsv+npHvPZ12ABDOXDBSQgqpx
ZEMLn+R0cq32p0a3A6d8ZWsRKZz0DmIWm2IiFz/ZARo2D6G1AIJZ2gdrz8uQ
Hi5OPfKmDbPzxDduKvVojF5mpDHoZqyxOeU7Ipd6HvqZ99V4JambdxteBqXY
WgtAx7/nWUs/Aswq+CTJMrRq6VKQ1jnH46FCISff6kfgHqW3A0y2zpyAAmGQ
7+gvSf2Vv+vgy0+dU7uO65fI6i5nCTX09HN6XtOU7zS3H8VJwGwl77MpMVRJ
ktjoI3XWVuBOh3jKaKjiBH1ov9qM0gwGTyK2Ix1TIRJ2Wo4CgaiM5lWs1HoK
DLHiPiIuUdrsQxJmagEIjutlfAmJZnTUJRmovSB1+W4WkYHoAkzq2So6Caum
Wvj/G94UfO878P8qLze0WXB4Ed2fGxfURNjpp72wPHbwGkzkiUJyGRQjwNdS
CvwU3GdLtZWJ0jVa5KIYsUVALU/VX14Fpuwsb2fZu8NQvQCKmgwDgbOpFGuo
Bl8MR5vW61o6HmfJnw7ClgPudMDaNUZSGfmwUuPVA0ohNPXIrZeWTc8Woa1z
leLhObdB1fYE4+D18PfgBpGcuteMPFPeGhNy7S6xXLEHzxYpkHc4RpfTJX3P
DurBIaVt93CYokgtTKbrDFZoSi86xKjvQ7zFCb+ZySDt6gOFsSTTtgxkYCif
GXc2ooTDcJk8HuQ2BdJwkI58d0VYGN6g9MXgsmxCm7qKq+41wAJ6CrnkZRUQ
9HuHu838C3uP6pTb+cbrJGv3LHAJYjz1BgJaoFaY6IgW8TJ9jHjPqWpFEoTn
bC0oZh5S4zSUrUYNSUX+z6I2+KoeYwKPX0ZtMYu3ZpVxbTJtV6ub6hP+/x/F
ndu6In2US3Tp6ZjkdKCLUsQNtThvkTnMrp15ezlrLWsnTamDd5dVfTM34Cee
l3HcrJdjvQHuHDN0mbH7NuvnL9h1GIagtdNiETq5OtmAgXlMuA0rTMyaDIeu
6Ddc2RUbtj9qsdf3IJ8y7CwIRPLGLsl8+CTaqKYjckuxCtazqLMOuOtS85+T
qWro04i/+auUFxOF7DRxnzCTSzY3SvzIDeTlSy2nURwQihuRZdwaZdK2wzeZ
FXHvz8AqgPb5DE+jX4lV7ZbLUaAVHCpcHz35xLD0WP7w61doAhZmUrLxFle0
rP4JzwonkXwgOfxTq6HUZINka0Xg4QQ/AWeq1ICaB7Pz1Bie4uSNHbHryi7K
SmYkCZjs+2DjoHVb6V9/UhofLKNC64G4g4zDxnF4k1JrqAcfo8RsLUpR9UT3
0XsOxIjp3TX/TuLldpb+snxhYutjeuhtI2UgHhBBRTH7cpL+7e5Cu0EWGLjU
sEszkWX9QqetMzEhsKBXdS3hAu7MQ0ieg7hRUtQLGaenhP3YqBgrgtj+4z8L
0WW1wD8lyP6apVYelPNXmwCzWt5KmwY3n18sW22EQEY4I4RPihyG5xk8t1kc
q9tNiHimd6tsKABBBkL7zIA15K2of69aSjW+vyFVCkGhS5dhGuquYNIPY9ZS
fjaaCRgkwR2q2E+xmMsBxf0aN2skQKQ2sIB8bhES/3YRNoF7nU3W27pfxPh1
ouia1THHC/Q9VZphGNz6w0pyMESnGxZ473lLs1WIf8+jbAShtDDClWuP9wpG
kqTYsGKJpwQ8eufJo+EPNi7ch5rjRvorseoQ1Xkzr7KNvjxK1W662lquS069
Hi78A06GjCiAm3us630XpGOHHEpYGsbzOSUtdPCgsV74XWPWPCnfNOcljVFU
LQr9nkH7cOfcGPpkHlITpbs3YVZR+hR5Xzqh/xvSfypJLPM+gs5tWPA/K/X7
CENOWcVh8OupQxUq/KRvoaCJZ6/VdBrn0Gp9MAWcC2OzuYVbzx14k3sRsdUP
hueUZyMkjpdJHY9yHh0qF1uYsunhWWhfP+2XU6UhX3KTE2ir34waZ4WQ4zWt
YC+cTATEufC87aDAhsx9wlJwu9lpzLMfkyS8TqNTJibeP8GDEhijuPVZstV1
Y0ZazK5Nfc2faz/9x4y/ATbL5Q7rJ4x4L2QNL5bZu2X80ccCdxyOcmYGWwAO
T/kZvLvhA0EuWCVj88XWRKh98RBe2lFFnWsGg3yZ3QbuBRV6EFllKjmv4ydn
+CxqZnfkzjw9HSgG78Z9DJBLic0ncsJeJey8rObSo9QGdKsFRhq9aTI3lg8b
g5yLBJEYEmkui6mgCYYk5K/rbTtlD52XJ+tXuL/xH2qhKzaWx9MUVWrEahRW
zr+BMdnVtnCLHgmawWuwPB2AYuFO2cClMJiEM+5RXKCS/lzoYq3oGHl8+otK
8VmLelKGQlzoIUbyg7XQVM4tScY1rZ+POlk9csYvD+ZiTWv15f4oW432xvj9
fWgqrX2vcjK3lrppwAaNBeDHttP3Lh5zcsX0uJQA2iyjuiJvziPSHm6FNPBE
9OtSRSL7Fldo4V6iszNjVC0WTv15X7SdIVxKnMDiKilG4M+9s6ztJ+H5HLpM
CNBs7B8Ffu78k8KHmknIMHV6h1k1jd0mFY1BnUb/AHUCdIAMZ21DLKcqXlJk
1N5XHui0OHhYM1Xw7TXodzMOyYCMDYMDJWxlsLXY85Qbl7biYDGLeenmZrz+
HcVIAaD4SzH+eZDnkjWZgreVgNhtVVNzR9a+5azoSA0hITbYLOI21ioFm8Na
7AKAuX6ZmOcl0kLfGjple+w6lFXhA6vKJRvtwJ6Li4vTAWTRzA3RpC77Bpwg
0U9k4w6/Q2ulXYVoUDDK4BZqzTP79Rc7nj+xw0KD7WwjgrO6z70sQbJi6XwW
r6vnmAod/3sjlHbt7waFuClh7y+tVmjwlNpI/JMx2zDmwPhXT0e039Z/E85s
nKEPXCvyd0bEWl7QopnQvUyBHbKotHUrWfVgiIwHNVxBXGSDgxPnkW4OQHRR
wrEffJIr0WDy2/M8GPP4HQIdjakAEhTAqRpoY8Fl2tfGVxam0CAAQNhWbHXr
6G8huTq+vNQq8o6eubdWCwuxeebRIoAoFX58cQ/wMZiKsM9emWgel4SC0psi
zjOeTYc6EGKpMrmT7CmPzBP3zdTEHkegDeWtDJX1OCF998KuGWf80BrcdnKS
ZvCn+NrTuRuix0cbWnZGJklrLZLDehglfDUCuIpa/OZtvfALgRkVWau0CYlr
nafz3otjb9w5szrM2gKTEsOLCOtB+AzDCzSMJyg5Cx+4MPjA8DLlfILbhpe+
0aYY2DuXsRxiDxrWk9l7OcgTxjupNK4K9yFBGKDKGgl8IHtDbj3V6deMfBeU
9TfGrUbHTz613dOJ0i2YQtGvlwDJ8X9+bc44nc0b65yYkYEBcBEVv9Ya0fh2
gSzQWKHeDK06onqICh363DLshLD5RV1fj1PA2ghx8cMHR75a6VUvoAFMmWYC
6KwMNPGag4ziBC01EA0YvdzNmg2qn49hkjrauPmPPzJSpbvQ0GnzrG968c7r
Av4hTM+n4nZWghoyWclfitT6VafgrbN4sfihL2GpQkKzc07A81oUHSoEC7Yz
BUBXG3Dz3mjFwtH+wZ0nVYCAaGDYRXTZ6s5hww1QS0+v/jRV+rZN1BDDYGt/
NbO9xZ6lpfzejHtsklp/ahgCcDl55OEvOx5aL86Jz/eWSH6TExBhx7U8VHK2
OWLhwGb43zHA2fsDCHFICavvWnCaVeMmopn7buKMqb9NVY9U1M4k3Z11EGRU
Kl3h13xTwy2XMgNSrEVlaslf1oLzJcC3ljdbulNszIjIMDO323/8QH8is3Ci
NbJtGzamNjMGMMTZieBYLy9/I/7OIcB8wiUT3efdEUfKex1QfoyDdclSxtVD
dRvaFZQCLuplv3LzQdEh83U01Pgqbw/JJUEYxYZK4GltBvJ2Dx3rOJm/rEKs
AX7+a+tpV0WmU8XrjeGSCGezEt0KVxmriQan5d0kwdhZpaOepVNL5VzthA6Y
w2ymSDhmxWHJmNZdKEpvyLGn9pztCXgPW1FIqrijpuHCpJawLkTQbOuuItdE
G7ISAYJxZiLl0i32vHYTAH6c9jJkn2cb4sFUaAVplTuakliOhesZO1LuUp/T
G7d9nk0Sf/LlC803nqMt8lxpIfC7zYDAY6brMJVw7UWJ2gGvj7I8ix0N46Gw
qQeUWLVA28hDlcm6hdkC4CRoFbA4PIRL8Fi83EbL0M9mOBKfkGBEcrBtFkXD
Rq0vNJUlMLwI6lm/jsI4XnVKwHHwRKNyAPpLJ9oQk/Ze5nBp2UJtliX6pTux
bILdZtIxgXMttT8sBVFCHB8SqIc2lauBXvzNKJDjNx23rly77z6l9CbqzR2p
9s5N4UqeZk5Un2vbissY5Y2yFtXtOPQPP7H/W4M700rFCulSIwcmlW3I0R3C
2cXpwrgk3gHc9pctDVGR0SJdzaXZeDw3gbC48P6Eg2EOMQmpyG2BLFb5OPHT
zH0Z73CbjjOW+o9tEyC5LT8GPg/3uhEMxMItMwUwaT1Cx0w0vSJbtxf1l7N/
n0inrn/R+mbOrowMF5MMF1+jkbzeQxqf/sttUnduwLcd1XLfY6DjDa+2V89e
szUnKiUeEyWJwAs/fUQNv8274VRM2+xSIKLsoXOfEJIf07MLeXg7ZYGQ1m+A
+R6Jtwha3O0lIBklYYZVLCTsAsS01G6+r1S8REqpEHf8utRrdIXZAAD8uM4F
aHHgKAXvJ6OkEr4Kc9t0j1H2pHudShzkThb53hS4rH8N1c8z/Krrg8tlAC+u
qw+o4soLmSktd1VYh3rvx29Fep0AIyLpIcYRJ3wfHq8IjwrwjVrJRF4zQLm6
+dT1o3dT7Z6Q8MYPcLM1WfaQR7IuIIfb4ogKHQuMBTa+kEGCofr9SYIxD2UF
a+R7hRNhkM8afD0j1ROm67JBkgbSlxI5tamP4Fyx+7fIFWzRT2/fhQ0LLFmi
ArNUEg2Zn3f96CVA299a929rJNmL1p+qD4i3kQoLGkDZkoZJxltnMgSNZ67a
0ggF6Y4UU/6UAheN2MR9gm8wgwYSRDtyqhrXzrI8gwbk0fPApM5ElCbWt1Zt
6jH0KoHadhINs8w8uOBoyagjCIg9W0QBum0g85GyH4oAla3OiqB1Q31gjlXx
tkKrgXWUi1axaGv3fFB3ePGsg83+nOVUYCi6biy9xPj8XAkIdiiQbVdi1vz0
7dSApP7RObi9zHSYuBQAAvdcv8DsXHaftcashonFGga1FNWzgypT1fbUdZZP
utG3XAxmFSm+/vadQD7Y5vKFvaACrdPHIdlEUwHTSpfN1hlsRSAW+0zoEtMk
QD9OfbcT868BImbIdO/dooeELJaAMcteVJazMY/z/nFaIpRzQdBYfaVm+x2N
t55sCMeD4YoTszre0Kugu2HHOh0NxtwNArOv0rEvPOAhT5uZSajhFHUDpR5g
94UzAsFttjuRLBEm5/wk9MV2lDLxPf5d0xWUOV8V8ZEfx9KIvcUZZDLvoT/W
OyrgTxvgR687kYuvTbDH0/JTPr7hLYO57L5I0z+39Q6HuHJkzf4SDqkOd+xN
7UKHclytvWHcLf2KJdW0AObiI8Vn4o5FFjJKCkfcCRdm1JXMv22nZSCE58JZ
dEne57eTk9kZswwFdp8TpNQoXH70iTLoNm/nvHezvz71hyhGGmKxMWNuHCjj
gPjRLvcjOcezYs6o4F+CVzxzN/sEOaLnGqPftB7KP72rVlbDyxnsulJQ/b42
gLtoLJlRe5T5LXzYnQ9lo5eSs8TlKIiWPfXCZ4ZOTO1vXDxf/7lisCMQ5ILQ
MoTzJooP4yk20ulCxrTk2E0R6Qp1qEUMXXzYzudXpkSRWbeMtrZ8+OsYQWMd
AkRO/2CXnVPUzLRrYiKSyFxy2vms5GvW3ISriy24KgW+JWgEkpCxsuNZG1Wi
snt9LIcqg/G4jfZTySbJioBnAKDV0kazz4NWm/lqK8HBPpc04TUiEX1huuy+
s/YLCWNS7fKmHJjQRDHPMg3bbWM0T9chgcG1MOjxVHt3IiHYZxWebmTiqqRU
wVYl5o8WRzxnMfgp2aCjNqupaSHlGO6G9WSWkBFq00cHDKrft4PHvjVH7rPb
3KRodXw0maSlSIeOB/1M9VMaFzeTisuZshbhGP4NlbJu1FbqPqFQR8qc92iL
UhbZpT7iu8ZshdlcPonrcvrhMmDJgozO7bFxazkJvnVDYSdHxPUbgzoLKiki
rDM7GZ8/sasO9mn8XVQvdBD8pUqQ/F3E8gTX/UTIfoqOcO9IK0bjOvSjVzxk
vnkMRg/2vDQYl2+m3kElVFT/s3fT4rxqzq5NvK3gJHtR76QLc8UfDdGIBtpY
8SLonXalODIi7Mp6GoXHYaOtHhV6z7abSDrTaxHuhZ+1fgfzqXHdrm0tTHnX
9vDwK0YugmNROI1hIaSNYKuyPqIIzJCtKppuHricCVWPmdP5rlgZIVoOSZM+
d8q+MqEULhA+t46sY/aaOVNnqN3i3uZRbRq9NARbXsLjPxcC0x7TOHIUWRTg
ex6kxwxziOVFOPG9aG6SZNgsCaSZN/XuGffDzCXgO+3Pxnrt2mzHe5QIIBIV
yl687SPdbvHADal0VDnak5O4pOMrOrUMMeV3tAubKSiWloS3Z6/KJ+APrr06
NJsqgJfcDIbTgkLm9Jle6kLSQA5g7oC853cWJyjvcJnY1B57HLkYFxOHtJ2v
/M9oxFwXqt3PhNHy7kRvLtFNpOgM5TtHjTQuhyHYHxhjMNLtEUJBctunhr/L
9pFs1md2O47DBuFvotlJQOYHjCF1QEFuGitlHqaQ7w1uomkGVf6sQ/DjrfXc
SZKd2k1LlJdPhOoSmjTiooSv6MSH7oKCGR5Si/oLQLf6WtouKfBaqK+aEKuQ
3XX5gxEWm80g9huc+sjULS+JUsfLsiWGRJ2DC3Az1RHkdruT4qnwDcerBNJc
Ep3MvdqaupRU1oUtTqNPXxJ51a/EBlokui+mQhrLTS3Y0CAs2p8MpOACy0Gx
ErRMTOGwueXW+OtyYoNs49xBkBEEjepMejhkAgohneBQhM3QB0jfqgYjppX7
bvZrquHPblKByT0PE1iGYYb9G9aEkYA1dJ1D4zJ9MSFnnPHBSRS9/36ZGm8Q
98WWd0bdY7kiVneb6ErNSEIkmzjdoR7NUTcZDfKi+SLa+qDZyxgmNB837u/p
Pe30a7iUwLengtVXKLbfGdVhGAWWmrNFVuipNiZIi3dhot8hlchq7vbLoEuU
LRq76keAUXNn0B8TvWKESN7pXi7pnbCeLlEodpOwnXu3XY8SjnsFdMvHpj2h
tdM8kBVFYPV9uVwtVs3aUdgf3WwamUk0BMF1ImD1OxLOCsfApp86rXZFB3qm
kSZ/asEL1Y60YR+yQNq0nN6tcxhAtMqBxKdKJftouOKfChiHc96RB16kt0jD
YO+otxmT1x4RBnoVUkf46jtL2+7PdcvUEwBfdfJzXa0GSCQVhUxOhy873clw
ivXJrCqfh6SFEYHZW3RCVNa1mLyyJKX9M1/xFdA8o+pXHpiGVZvZMnLq0/9g
Osnti0yQDOm2iSjPDhWmasIRTmfT6BXmxFkPo2LqnT/kgYul1JyojElk4B3m
XguRkYMVnZWeq9SnkgINdGxwhdWPjBAJ42e+FdbXSXRnWSAmW6/gqw/kfFt1
21m0ocp14lNPX4aq/dVn+wmN4Db0bG4WiEjcFE3F67f5tx7uG3/5eBk4E+FD
XuDAjgftfNCW/n+HlKULIMdXvcxAbLOxIFtWgr/wstbbiIYnwfUTCqPf5sMN
Cl1Dt6Csj/0/Oan+UcwqNEAS9btefG2Abh8ec5/HLjOpvmq/OqTLmkdMGXmk
Krmg43kGYL3Qxm4ZF9lX66EsOnWtKKFPesgYw8N5DtpQHONMMsBg08LDMTl3
MoiISE3JRlbZ3ESKvxJfWyHTg4roQyPAUQtN2AHmdFZSOoRBMIeqI8m80Htg
UlhnYvdiDhFw/XRuMbplnC8hni77WVWyVNQSyRv9P2nCXlEhFTXja9UNIBt+
XSnZLEZ8Eml5omzeInVNTwpiXIpE2yQaw9brgtnXUS123vgcLNicrA8c7qob
rl7wKWipa4XFy7eXD+XPpZ6d4FCBbWCFF7kmmdc/pP+54FB6tCMLe8IBCKDx
gOztJ/1xD8L7ljKMKLD8+8lwjUTbOVFZjcjRuo5kUtEwIi3duUtf5pbz1VzQ
c0Q8TgivFUQwOc7W9gBdt5+rnuJw5ttUCUDhGhxDs92P9qn0Lv8ZAy912J7l
N9paA2MIKr0Nm8ZOAxjogpX5FdRMRH+dLoOZjAw898OJCZ3umt57jr0XIGO3
YusgGmudERBS+mlqKS+niTChpkKl+vtS38C+md+DZ8RuERwZpo9AzgHYLqVd
d/4Ijyj6lbGsKkc5ujoEDmPSArclhcumwz/LCfMeeJ/qGM3KhQ20DnUvrtcH
oW9EhV5nYjjdAqmimj3Ge9XLq31eaCDwUfcAMpA0hw/BWy9V7O1BnSpTDPzY
gYQYIhZhl40RwMt7sTpHyh4WyUogB5ZlB/BTBlOKUGUgYgsZQCKC45HCyyOz
91t89Vgp6ZWfrb0mMGTCtyEbkbGSymDjKxZZc8gYP1RHuTxIw8I0KgbFJuFm
abU+79fwl8EDvWsq5IG6t1/i42S0JeJ4901tiMXxFL0ti50vQILF+W4MDMiz
PiQqFBBDeSPng23Y7xNkTuQbCI3v6Go0w4naQB0doAHCFAOgRpCtTF0OyKKK
UDMYDaMhAGS1QqPIi6FFWIa2Ks3vEzvlYtj/7LNzChgv5fkadMnjvsg1C4nD
AeKMZMqVbW/2I5jvztWLxGGSHYwJRLu7ikF1wRBPXGCgZ548gtkTIKUHKGmY
0BOS0lCTOWEotlO4RuroqnjuPN1RPSbtfk5fCm0loDNQVMwnO3AlQ/SqpvQt
rYtr87aab2nNFYuwD3DVeFsxtE+FMEsFmcf52cd2ykmxkEMG59gw2nhfAxC/
Wv0QWfJkixUQ2lrqDSSckFpI/sHw2vvyxTpDJAFQ+QWwhu5VMSc9IjsBkX7i
+022E55sEgmtstUgEC9XO9r2UXqB/nrz/EMPFx3+npPwXqwhXvtUW+hvnybF
1u0qq+DCzH1iIxD4Th3vwOCUDcfoJz5x+B6x7dqOhsDavw66IoBT1ICQw8dR
i+VRsq7zfjO76ZzDtcskKAk2MwVkW3jcXr+KFBQ3DVQCsAlqL8TUouzfd23v
Y5x0z2d1MK7LCTzXg9JgGJWMxIrQgAXW6fVGFaSaP0pg1nRxOz/Hu/U/FYs+
PwDwtB9SO7P238FJOTj0TiPYCSRCCz/OlN4drsr1Z2oINOLD9as0Ac7VkjXb
IZQ5snbtNhldGWl/cHgTbCc3lL3AkBW0+ZrEK5vsZz3JPZ8/WRnaW3qFEZJo
S/N7hKKa7KhyrBOX0rYxLWHS4lxye9F/mUYoSIKIuCp/HAhlpMhqjky69SJm
jaApuxUsEfBkZ2J7SnJO+Has+HqTuls+Z//5bQWKGpKryhjgoTv2JSxbNPTC
hxalbG1T3Z7BNuPAM4dtYGr5crtGSSzRSQcsBt226IgKQUSF9DGWDG6dOLOT
3S0VSYn3GS4JGG+lP+l9WUN5rvQUJNZaWKHhe1PBqrhCRIT/BjrI5O+rDq+A
e0f17gIqh1b9HAXR4xNyBh63u2umaK5/U7LShwA050BofFolCbz/x12MrctU
p16DR7C2W6dbmTN6D4er5e5FOUxi3DanS/QkyiG3phJulkbTLWIB2WmUxxFi
hmB02kqKGUvcOBgg3CH/cNc0NhMYsSuAEv40Nevw5NW07we4qvs0mJ82q0r+
VXuDmLx7QGTipuUkQqFTp5HFHF/cSWl69EObsJInNyluiJnG0xj4ulSodEhV
976DAC5UgTw4XWX4xb4imBz8ebiDn4EsWLZGj0U/SpWULvWdvlPmUhtw1mkQ
rIokILcjOOYIzl8aJufkZyd3/DFIjWseZPEWd0qIfl7sZ6yfayYKvRxoBYqc
hC3hOTd5MzvALNSbP7bTW96vi5iu6YXIwgsRE9mYYDKsAqo9uwdNZcXO8Quz
RAzq6Sjh+XCHKJ9ffwWAorv6Djl+vLWCKLcwDednsotP4qREi7WkNi/2O9A3
i/lese1AHRLqg78N6wEFPwytbb7Wl6mjCedUxfGAEVrt78D2s7yB2etrcM1j
IbkrMgCe7q4JclEi6JqCakajWqebI7i7yfDM07WFmBsndHUshJKb1O22tODP
W8ct2KEnvEZZKgpzOU3fhNL4M3XjBxtWbDjsCMlYY/+HQAFPCACP5+nkM8RC
ziEVHZOzNa6R0fk/k72v/A8FtCuPIHyIVnzEsZ8ecMDToiB3Pwj4SGqdMTdV
QoeJFAIi/5Uw3W8+f6tHuXW6PwNwABxsHNYCBD9a9ZpeHg1yL9cqlL76O21V
jLYn2Y3t4w/EFpG3Y1uNsbnTb0OsqZcwz1vpK1gMdWMA9CtexczgPS6q/ecC
ZaLfl4GlDOE+Gruf81vvRA3WAerceoUmllD1xOnFccBkykbCsUwOBuJUrJUZ
XEqUUmAS/N87WrNhO/KrTqJnAtKNapeaF4Ff24UGf7OCQtomn9g0pRfT0+4c
sbYFHgD+q37NAJjHl7znl4HwuvgQVt4rElmC1Udpd9NjOyAXv3MMwWlV233w
u++OUQJtaYV0QnnMR+M0Sr7iWr0TUyDtaPMIRO0WISS8sX0R6R2ZJtirbOXg
zxObUvV9c1qmVWF8wVunmWv1nebRP0pFzCZEWeVHsbHJQJEmss0IBzXmrDwM
nVqipAx6MqID2UNKDRwMprJYTu73PzKAzqAriDOIUjQuqk1mMvnUX+h4zAG2
gvvvJSdWvpkAv48omNnV56kcQc7pC4zTbg9qM5oGVrTp+2a4VlFFLXCr5uJj
4/1YN2x+IpTHKEwcKiMcz13uz4JUOV9sUYtDmrLDpnJx2xun1wY2zt9u9OIa
gCC0l4bwcl9XmhFXTAUSeQ4XYv1fHMfBf6Ly2eidN99RhXbc/9gBfS0YevJY
9ekkUEVcBH0qdHuFtqVFElOwgI0wqjQBuQWiFAQIVkha5MCl39WwZafrHLeX
IYU39iz3cPu8abZ0JeTmu78audw3wrPWJU9jlfPfR/9hdF8JYAN0nyO8QDgN
EBdtmWXsj8tbBxnN0UKFQHwVE5YPoauXG2x5H1KtAjZDV4Az5SNeA52Gsbkx
9fbfNUPZLAcqvmhZ5isbLGerLBFTd1li6ex7A9jFSxet57keTO33p7yMXGUI
MhfrLxtaKgnT5RSbrOR+UladcqhOUjDGsWc7HAXEul6CAHzcBPF6O+Mf8Ige
duCxenWQAz7L0/T1MyyNDBi0Kk3MiHv5DHGL8ve7xK3lxbr87nOYlBVxC9/0
wzdu42M4+cll996x79KSjXKQs0Yvl22WMq3Lu4W43Go0jgz3rMFCUjPW4g9+
idlTY98AvDQsOhTyxlp5SIoWrIGt86NPGKUUXL2rrycnmgEwffwzpa2I+z20
LinZygZ72a7FE6OnAN2V+L4WHppkRtMhS906GB/8TIC0xkV3gTj4Fv4HgNZ/
3ZX8pxROYP0Ukp1+51zo+kYWuwvx4JeBsZ9nRyVVdR9i/uMwx5EZkahRFwPn
Ryfs6e8a4cy/0jc6AxbhsS9ZUFO2m8KavF0po/oa27htf/gD/E8DHLFQGj5M
BmvVhz4qRbE+udztDxCjWTv1MoQQTxF2e9B/PgBawCLFZPqhLXAmoGoCt5QO
jOhfG9ZeVUPVDWl9PmD6yJQUPRaLnzJcVtE3YW+8GpLGNpG43z42F7okhCfY
PLejsz//r8Caq0nHh6EW5tNHBKk53xvOMD0bnM6ieXY383TaDSSiG6/DU8UK
AGUHC/k370SK2s+zoslytTzcVBKBsXs+AevUskl+rPZbd5OICbZ+UlI32hrV
23+BW+a/pR8NAxrPynu+QfcjzAdBRDnHRBM/sy6/l2O+zGq2t+4x/XTSfG9K
SzJ7qIgfo+YTUTea8uoSCAJgHWrCpce3RnDvDbnM7bPCNlLPrzg/hbWP4X7T
4UzjiqRnSNWNR/2/wtr+ZPhALiaOxwM7+dwH3NF2+m5T+2xIuLVFhyNftLP1
8QCi5FxcQAVBly2nWrvqXi7s+caZleKMCxpaDbljmMAVT4dtkBcEjSKnn5Be
KHXbxHrKdCEIM9P4jrKxnwgcwmNrLUNBFwC7Dvry+HLnZ+R28BGjhy44sfXN
n4XGd+3xSl4LnrjOK4OTdyJIcuT7MhPtGxc7cxI1o+6mlpixH3Dx4V22aNnZ
Dl3c8nUv/hOPhby7MTTbwy+JqmH4fyaPo1Kw2rgaI16u1FXVM7OC/ZrMazOe
InIOunzaNP+X1ZKBw1FwUglUg3BWjcik3sLQj7Si6PT3C2gmXxpZk2/QN1lo
MZqZOkMmLgMkTO28y4ZnuoBeS/uyMl6Chw+uhsfrwH4nGjAaWNNbrT81/YSP
P2JUe1xkJr5V5w1o9DOXabunMneVPt5/wCjmgw/I/m64puR8ANCONkzlOLHn
1mW/5fuqKoINuEP8OFHLtqqYJntM+WrD0RzW+f724AK0rbLItE2TwNe7mcFQ
MrYy/NdPy5CmTBsc0nBtSQsfy6ebS3l21Ngaw5KByLp6ZFpVNuMMvJQV5kWR
MGjAwnlkPO3iXBpWLo9l4AoqnD+Fnh1FiysvMeNl9xfcKw8mtvgDupb1R4fP
MoQ8WraDMsvl6Z4MYQCbm3n6wPlTBq+oRughH6DOJCgCqPpr2SBYuIldoIdP
KBbdfCWDwsUDgDDN4/q0i6AaN1GyW4IcFewYYgRjEAGbshOY9LLjIEauY6Aw
nNS9V/sBrb75ckyG2tSQe6gORkKFj9vt4VYpWGOSlyQsUhE91t1ruJ/s46dL
vto1wCk8vuK2EAeM2j7Ut0Gxi2B9xxSCN62yGpw/8Iv2/C5eb3UMYHkHnDwI
GxXq89dTQqj8vzbwCgKYVU1IYqrrRARr5FS93CG5dpCf7Dtz4fBNMwtWTfWZ
PP8kU/k4P8cWdkdyf6B5LHDBbmUPbec0MWtWM9F1D/713Y+Wx1w3Au6noYbX
A6HGHyVuBX6l5YXRAlkL/8rE+0qrijZEJj7W5t0PCMB7ocTMIkFeV6aNw6TH
cW8Xd8Lj95d1PVn5ApLiW28yCmvvis27cpfE10ZdXZGJXS26GiB1OgF3OfAw
6Ho/3FZuZ2pd1EIWKWmpxxOT8KkMvX62W7opJtNITZIwGkwutJfawOMzULG4
PTyCroxkxap3gcSmAjfd/jHAJZ85gKloPdX5NVUbTkVRU6RYc7cHCR/jFZjU
ZGksmaWBkFCS5ztpjynTuDyYiVoyBL4n2gyRJW0givcZpd+pIMGqBBlvYcaw
EI7v6P+Nm9rjHDY+J04a2R+di+ykieFNvF/MRyKH4qPn2VqDh2w8xJeEvPja
58A/vzzXfYsEE9NSEkh4n8xXUxlBLcOPSAp+NtTXbyjH6y89v6w25KYP6yNe
ssf+W+Aao6aHWXsg+YB8sLm66kE/luhMVnUsbgUxQGJCId24OEQA1JCU6Ex8
M91swYF5tJXlMy2dAcy0cfuEqWLU9d3CRXzy54Wz+roUzDvbJJY77SPe3WK8
jD5PYM5JqYOTJLjMIN62vE62F7c6p9R4Cji9v+kMoNOVhpMuuPpHtyyC1tjS
i+hViYyw6G5KKrFiFKXw6tXcjiota3rUvFpUYdQh3bn9sZAyoU8Besy2yXrf
QkOvZtCs7BW7Kdmg50UmFbqQCHGfzTxIaA8iYmm/qGlVmcbjmc5VaYvhjUwN
UmVdpSECF1JL3n2VnGeyBArfivXylqP6br86Vf8Vpnc54kCHqX6qzOFvfGKq
tY/57toJ+vKzDRPiCeYFrhv5em1PubITfJ+XIrxWUEA0BowlOF1rhkd7LRKr
NqO4M3fVGkjTRmWRwp8/AsVe4MM9K3kH8+K+81LVuR2E9cub0f80sHIYWGh+
ns+i6EJxVuvaVa+7tQSprd73Wo+R/9x6Yt7IGE0lKqiCjQ3OedWhHdktduIL
FTNl0PtP3dDhv6oXn56lv6yBeme6yHaVYh7BKlu4VlgDjO/Tts5JRPLiAP2k
BIBNur+u71WuEbDyn+K0TAHr7p96ZxYm6xE2/1ANyYLNoIERem51Si3SbUNf
lM69cEFadnf0LV7s6MeRCXvB/WwwEbXCqPlYE1Kqs8X1VolUrnR6HF9m3yvk
nfw2xPwZrIspwyjCjLPYsrW2ITmWd1se0+JvmjQF5fHeS2BNr4LJysoJodtG
ZGbIukSzVNPpUqxjDm+V5hh+/bo4trpP2GSNEx1JRyXhbmhMvwqOcr8BgD4/
XRYHXMY+QJ0IDN/+3xl2YcXyyGAEmRTdES2dH3lpubSAWF6ef3ZXKB+RC2rZ
LLN2WBM7SNVqQjN7GX/OClh74tisIAj/AqNxtGAX1pdmts0wMyyfPUP7JRIv
Zo0gAO2G9odjwwu22N+QjW6oNthfI/sf723cP91MM0wwALrDZwqCAaFXeWU2
S7OEqBFrBPb5O4sZqTtgc9OQQ2R43wRC0INRJOcDT0crhxmE2DCkIcXeaK9u
yuGzBqotEBp6T2v+XAxM1SHwaVCTDJzKcV42i2HYBFM/mn4Baryw5bqBnR0s
4+vwfX8EDV7DfQcd2TDbNfapi2kcnU7Nh9zyTaZkjb5sasLGldHB1XkUrTFz
zL/VrKCYpVlelh55GaL497BGjRvLSi1FHFgT7hwpwjr1+3K82W2pWXdKsMXf
Rk7R/hAwUndW20mu+nUykIg9m58tXiyiDDujZjlSbCqSBEKlvLGAuLEUfMF/
AeJ/+vsEk4W0T/3ESpYAxpgMeITAzB1GzR2kHUXb/kuwElRfiM5iWOyGCOMP
MFT3uc4MvczOKpPS4VGIZMhh6m0nCq/UElUAXm8vMpeJbs5uW57CBzEdSS+s
K16mhgdzhdi1vD+2MEGV35fFjuGLDccu82rUUJi32rE7G74GiXiq5uJy5lXN
GQONEj/k6MlmD3Iv2eF9wtmlFFJR0zRDnZOj8Cdvw16HsMqmlkLcy5ThARhQ
EiNMh8awMEIPkMWzmnufVJNb6NXkXzk7+LB867tp3a5/pLd0DUvF7XlQaF0W
xt4kJMu1UqdnXb6iNe+AinMJEywJOXsORGf64p5tb4iKtKNdVTrslX8M2lax
wib+SeVKvVvxqHPlTipE7ESaGLCSUQSX0qbkeXayie/YwsYeEFCy98bhdfAQ
PDRermIvam66tymCzp4fJpPsAnuPOap9U1t97H8cWSh3MrPUkOTRF3pQNeBd
ZLgVstwrtJRJ03JjOKeJTAC0wBA37/B7bttddVtEqdL2/3c9lid0E4ks8dqQ
wBqnDsa66V+phhgAQriZ1mY9pRgT8UJVIhAj12nUQHaL3vW26IAUeX4le3Rx
fqsXXHpP34aBVK9JIHlr8uY/rv0rPT/MD8djMTIdEB9SVBNLJNI+DgtI3iQZ
+AaP8bK6Yc4yA0oM3t3fd0FVynb6hhrWdNWhkCdvlGpTun7/Bf8edW6lBcFf
A3Ih6B2KAejbmD4O/WTjbRux0R4IWol5LddkTiU6xYp232BmNaQOtYI8Llxl
HexKdUcWMvVFnmxbQDDr2PjRu5DT/gKGGgaK12zmrbdpZltWuvwNps6VZswN
Sk+jI/YKr3ydrU1leVwbc4t2TMeGojjwgtXgyfL/14SZkEkFXAZX6INlMOzm
Ukh1+kwz8AYr8jG6RF7DUnxjmWyxoEA8gyGxMHTlhC9U/crFPU6GnA6pRAiA
A8bLqdQPKuXlCtrXaRBB9Lp4neOijU4JKNCRrKydYOts3MKcuZ81mvX8bPHd
venjUbP9sM8tBGnRzLZDdX4xlmv4Qf95NybRdlaGyFa1MBy2EQlNiiuHn1ca
+kdQXn/QPBAG/7w6qoTqkWMuaSYvoL9h7PezcXmks91JI87Z/NHAaaPog7x2
VLZoIFn2GRHa3JEr6MM9E0VA0XHTAo+2x8bipSEDlr8/qOO02JcoJxc5S+A+
Q4eAHOfk+wK8E/X66jFWWhdtMSdrRGiXoihZxo31ldEZfYZvoFOodwLgzhpt
aGWSSlOMX/igp+RGORqqqLFI/sMWY8j8GhXYnEtwZkerCFLg/DpPYbrAFmAF
B5BYUPri3DXL8kOA/rmaFRSXjE98av2AJ297MpzbbQgyadv2mnemq9/eKBC7
ahxZAobN59RmgrzMKga/he/EzZDsO/+Zi02h5+jVTimv0zh85SNelppGNISK
IBJu6eIboU58ynTGvhqZDlT1YHNhExDPrBhyePr2CcJN51Ufi+Odf1fCSBer
eHnyGMkNRwJ7B3eal7XDWVTfQkWTm/arM7xTHqgXTspcPqjcsA/DvAoyPgbB
k8QfVzSEQi1s4D81VJQ9sQDmMm24oqGu/MQVldpoivL+PriW9YzcV0DptUho
Qd/7kjmnfF940+lFWWS7KwOz0Fo1E6UknbD+3uIS00r32ShzgMVbmd10xTA/
0RW6O6VIvaK58Kc1fYG2XicYGVFPa9bY/B+rAQhQNRuPa9GQ5uXwRAMUUOXi
9u1317ZrVI7i7Ls6OdCwj7+VtenXbTIatedzNaIzsR9eqlcJ14UuCJORO1KL
llh0OVIFVaRax1SDWhalVSrPqzdypWhP5F304Sujwx/j2w6QK3BD+rPK5ryp
nX7TE7rE8jCqRvPv3CHKbdN3k4copNabfCQRtFkA1oCWNNsYOxvRFeE5d7Ur
s+ASJW+yMW0rocBUwcMatpGBNq4lzNju4tfjuL9slpfaFugCqvLI+4Z0FeHA
7C97SQudjvIGAjzjk+c7imwLHI2FekkR+W96KLmaiHEv98i4iDuuJJdfJPVE
mCz2ul/JAGtJB1Ox4RA7yU+bLfnyAlxpsHc5tbTc94nTgOi1W/Z0CpW4CH8D
gs7lTmJzax9gK/u7H3bQFr6/pm0p/+Mne1O0eYpy6xxMaHTmKv3sBn+DWgyi
9VtNBMo/3d6m2TsAgY3ysm1BNAWYTHU63rgNoFs/TA6xtQBPF9bKyIEUo8+l
tErI7Kvl/zDIx8sIfsWAKkWlt6zWKQYVBsvgClsLf89uI2dx76vOb4B+KahB
jgIazWirKrJ8AzRDw/rZGbfCbZ8ReFm0ULsVCYI4sOb3aNawtwKLESwb7NSd
Q9BqKYwOLIeQLsjzrwgPhCfMRjer66GcxSVH9ft2dtmXS7S0dRvySbgXjIeI
Nrs36ggUdLqGwu0zRAoDcOklX4OQjGmkmu2+mSjFFhRsJzjD1kTuQDH/BRmN
t6k30VBbE/7gRXrn/c1ut7WTpnBzAFhWyNq/ZOHy0yqzw+qDEZ+nESIIteqm
cRxPAfXju2jOsYk8K/r/t06YxdaqAz8F2CHgmuv2aQCwZ94g6y7kXblBnv4P
56O5l3v2puUPFUBdBUFVFfgzoarawW8GfaqczZ6scI8D6uBn/CE27LPJC+7K
TQR1oOpvN59Gdgvtf+ncTjJqbrVIRbrgjqoCn84wji+YJQ6RW5GfUtd9yc7D
z/h/Il0CzyoM7HSRoIdgiJvAU5b/OyRFYIXE8rNWMxYf5lspzH7j8fQMB89w
cVBVkJk0im81ROX7OARYV+P6qV+o69EabhwEohR+OjGDk47c2956mtbWV37C
k999xrU38JRn1FaFmpzon0jq7/DMj2TX7gABV5LUxmaCAdMcSfyjzUzDqkOv
YiZMl190ZF4rU6r2KdjftEyzXvgLud5fFjQ4TFBUdrYF5yssDTdRoAio1FD1
rAwRfvofZFpjjMNrzcGAn/JthTekYk/FMXwMVLZMrBUcpwlIKqQywIhWue4h
IA6J8+Lcc9INsJiYEa57NJ3A7HsZA3MauwiDcVpNxJ4o7spPxY8Qx6Hx1axI
3wPhEADP089zl/w+HFqKMC8QFBkrwjQAnDWldtLWmW6WN+hnabHumVlqG2+U
0ZzE1/XizBShTnm6ibbk+4rqTY4AM+a5KlmLVuYplxLfTwFA3Ii+kvakXo9o
zxkw5+C43+nIewoYQo4ERTqgjUo7dUyyc5NXZRv8RqTAeSbiOmz+SOub2A5l
N7tns62X/VS3L/X/PpTkoKldNOI6l+ICILevGzmVDzM0LezGTI7qZbNnb1FH
DMSJSoJzXyZ2+ULZVKwoWRoo8+YQUg8nhmJU2y+MO1EdsWkXWAl/2ZQ8DsvC
y6MP59JUkj1zr4GskkEDL7Pk1D7ouuSWE9qHUUv3yahGHuULa7qS5uI6WeFH
nWuBHISf4lnSQg2h5GFbJIUu9grbrfZNeW5Du5HOOiQrMAlWkuKKfPOTml14
NvhRMwbe9XIr2Je8hrviTUvBr6iZvEWcbxjqVBI3wAyUalrIGg8EjjxwnKVy
8tzkOKgBXnELU9XYpaQwdMOQS4rswrM4MsooXKQCJYKvUIdRnwFDJDkliGbn
LpfANDy9NNPn+JQN4Hyn0toXHok6pi371hyiil9lOvdO0gMGiQAyL88db6e7
3DdEFrOA5qn07Ld/Dwt1V1WIreADT9at92CYxtkgT4JdQZvYjxnb1LJZXCvO
cSwJ1mfyW4Dq3yIlXuquk1sfvR6id1nzWMld68zP0C5ofKB7hrfKrPbl59Ts
90u+kvG9GL82ppt2PBqMX1/cY54yEnixTJHMO4ApDwwJeaX42/tVWCR6MmH8
DChz6j8oVis2OwKAA2E3kKBzbopoWo3yVGcOY+KBsD8NVF1t+oI9q1GGtRAK
H8C/Ck5ZpdREFaKCmeBv3YhAvRx3g2I3coWlD1H1uPf6ZpCiteBTABybn8y/
TCQaDUJvnzQKtNwdWidL0LQ9CR409VpN6qvgU85RoZ+g1PLD8NtpRgrB7+gv
iA6jUtdr3hiFBnis6UOKd3DujF8OWagNkHKKfxCaIOy3XiS/tNaamRPo600O
kIvVybmsz4PC7UH0QfbHFre55ZewYLNUhWzb1nAejN2kN+1chJ0LaaQmuz1+
+JUkpK0n4xjTSmsbHZwgoeed0SgVEY3n/Olwlfnuzptu48vyo32uulW3dSqd
OO/K20/HwEATFmuzi1TDGU5sGibXATTseU+xxE5As2PlCaohJHTF+iOKr+lX
9mxnh+qfSlqMOvDtEhY/cRHe9x8VgNTW5nXEhoRgnl7RAWcTwUa1iFXIigl8
MwofOZz/4PklUgBYnmGA9UfWy7Ulbo8/xNHu90E2FzcKyK/dpFAYujlYc2IE
Zi/A2tjvG9dwaOPR/PVRABFEZGt1kybnq1BrfgosuS68bzey0J2YOBEUsS4t
WJ09OQstLRqUYOby4j8qHrUZuSNjG/iqw73yN8CzYKE1JOrF3yizEiY2SARC
dybx/ooZL9/N4vqAAOe/ni8YXIg3Q5AeeaoaoDxztD5MpFoigzhGivlzkYDk
InypUrVmBH0JL1GA4CpVlTSgYkQTrek4g9AB+9E+Oiyn8A6F2AUJhbNI7dw0
5oXrAIFIbNvVHU6XFjqsxFiy8q/L6fhJ3ExlQcdagwM5Lz/nbqddMUxmjlgv
pGUpw7Tkb2n9BV83IojLDUn9a6bjpzJ7jDa3+UjmwzDgC7xv89VZ+gJC8Tbp
xZI664HL5P2/eC9jANe+kg1PpnwpmoRhUoFWjkbtIJiKhWxNpk5ysS6EuYx3
01ZGljZ+wEiCXRHXaiW6RtpRvd+AiNOvYhrEVArknQETvDGsT1FHCG+cKTm0
umk+OeHZv2PSDlRIng9qDLr1wpk7bRZLodS1JEAX+UPsjVmeWbBhyWQA8aHv
uvJ2mBvgo5YeFB32qP4Ye+eTMDe3xsvL/RuCXxX0a4Ub7qryauvRf5KxNqH6
8hc3Ys+yi831dXqbGLq6EvjVC8mswsdE/Pc9adlH9BPiHbZ+RzSqQaBAoV3J
DZNZ8S1PSGqi37IiX9jRTI22gy75kkihhrsrAwKoHAn3XVQpeUEWVMozTTZ4
FhNv4vOxSCKOOrF3LzJsEljiWzsxS1rIsZtvZd97pjf2YguYuyeHff1/ZmHG
3ZZuHJXEwGtuczJoGVW7986/MlN0zeUhSQb8wJP01F16g4ATIMfZnhIr7Kar
XkBF5N4C90WF950PSiho1ZpgHDB+5z70RamTQaRvXfZVIs6EI0da0Y0nJVmv
AngJ8wP+seREcVabBUqJ+dquNwRK11cSiabE95yFcWKZliUoH6Ga+/T20XHM
aGKAy+SN0XGTLABoANpOxHPHeefGUsNbgeG5K+eZuwpvfI2cqhTVEqYdn2R6
/6Xi5a2C851qfDvXdiq2Ck9c12jP/MRSvF2cAVhh16eBINui6sMf1JZ1/j4c
MB0UM1tMFdEX6ZHO4eeZI0E7ILRPPNtmYqWBnzMYNExVMiFBLQtxO1dA4XBn
SK37Dc+H5Yh7LHJLGzfXyh2oYCp9wWrjKlYZ0w/+lUBi1dZPOi+fUBpgj/IH
Z5nP6biVVcXzQRugB/vgDwOFQsxUnywW4DOrmNq+oXducky0r7VJlC/a7kVw
VO26vLD6TpUMDsW9RcIK3BI32naxts2vOVBjn00kkpkHUEOqkQSy/gKStETl
hjHIBQ/Hsfacfnb50SVIUH6ekseQQBHoLRE/xWMVyBaW4EeK/V0RZMEdJ/gm
gf+x7UTbJLgXfpSvH6x8OC1WnBkDDVzqaKiH5m8YgQGfYo9anRSOK8gBueOl
xLEdrqbtBAjIa8x8q1hMmT4YJBNZnUON5f2WYt8pyX8sypxSP/rzmLxhGilq
PpdhH4vYEYfIxy0o+xs6MNI1CZh0DZSEzFCgWhMbsxWpvn4D5/LQAAC0z2Iy
UTmDm1Q0+zgEzq9NYUSUA7L5eiaUm3s5BfUVABgt6w/Dq4RcUbCyqMdxva19
BEPPcS7v0ZihEol61kRjM0pansaXafjI8Afk+UzZFaO+AhKqbdNaV5pBj7eH
M1d1+zIOd9+jtGZL3gnhaSjrrDs1wek7iV26W8xTSS/86k+Ibcfx3e2MoTgi
VRt9B3kHEcifPcoBXjM0h+cF/h0b+cgpr1MVCn+msv7TArJQaYjIJFDe/s6r
Ifj7klDopXsRZtGv+MJ9gSUolFjgBvc8APFrk0K9BED2jSFvuDdO527sGljm
sQ8yEzGTHuDtI9HOsd4PmYjWrUK+VIKUEoxyXMBM6JrX26yr/eEUWaJ3BAT9
INwpQJL1bDK+Mtu9NUVdCkBbTBWWXvZ4saUyZwhBdsOxNLjPJYiPWkoaYTw8
jMJth0SzHPQDlUMVxYRRNe4mqnvR+ZXF5gXMdiD/uhZl7pcGZbMs1vOUeh7F
wQ4ymtmTs7Arqv3qim98D13dMQg2GqYasUBZH9C+6D/r71OlkCkbuLWjn4pm
+1tIXLwJZkmK6xxgJzz130zx++nWH1e5GpoOGiy9878CzWjbykJZag7FbIlW
dMJyg7ryYjXSnYt1boTnNSOtFkzQ4pAvIqsCc8u47x9o12FVD1SfLOwJCOXu
zb/qUc4hmq2QfSfamOGU7zHjHTkzPqxZqG4bIk1UQQuU0D6OZEV7j2k8B4+u
3COQvhxw0CF7ofJ/TgDqUPMn9Qn4p2M4Fq6CWnJ7pxd1VFYC5PfMp7foU1YE
iG9/i58RPf6oFR4nz5D0XzsFY1R7iU1euFdFY2qOJVn8phoNVXmRhFFfvDZf
eetNDOYT6La342pXI0Gic8iLGfT7dzgD3ldpa1oIpcGcI+KgOBUmNHOEMsSg
8XNKUIbNzvhu2vWRktDXvHcLkcxJqkJgBuUyZoB5YwW0VJC9A6gnODIUYELq
UZuXpMPvYU/BxfT0GjJsYRQiqiWvq6e/CLg1TzGT32t53VtpH/axTAgN14jC
Za7up6QPF0a35lUPBghm3okHXyjdDFTCPATcoMpj/RNGc34IZtGmfepqHVuB
p5knvrq065HsrKwk08wYP+ID9Uu2YfPSCxnIChR+S7vs/FRIPUlrUsWEJtr2
A0nldlXp0bMkOb4W1OeGh4QgwcJTvmDciw98MAoUDwOVfNDrvPZ4p9AV4H/e
a1thzIabrrAZ7c0zxkm9B7UkMf2LUpPtk1uX3oOCkJhkQqdrbyD36g84XbJY
Hso40vjIVY/o0GCP4XaMlcFGhXw7hR9AJlkQo+2qnlL5bVVCAFULpKkxleTM
L1jf39pIffEXNNHYcE2ZLT14OeYb2haDGgL4bqI2Z7iC3jCRwv0vnqVhLULs
w+30r0HSDLdwVDdcnBi9HuzX9xToOXBJiC4toKy4wqJjCDwfXSM/vUBRGepA
WrBjIq+Z2yB1loICRqSWpJIsSqXEjJyfr4CrZ8sy56EeSf7jeqcCNR6O3zn3
y6AhuCRg3rauNETc7ySAiDfIY8vR3PZLbMu2FMblocemlA4kn7ag/1KniGp5
rkJ8Ips2h4qKVnl8w8CsqZkE+h/IUOrqOGJm1w71E2iizcoKUt20x0yr0UqV
6O0xzsU01WJEqFVTIbWa41I7cfhnazKIWa16AASiitYENrooV/epLXf3BnLb
VZeUECldXjxbCYYpM3DdiuAdo1DKFcTocu/UTbp8w5t44uC1ZfZO6buAQc3N
Ca4uOFdA0k18YMvVv0dwkEaDXbtS3te2sTO2RQaya7/3lft/JhUgq2QDFkqp
3tcvRa3LnzbwGC1xWsUWxiWmmv2ru51WkHznOT5mKI0sXAfEyfxfWN3j/Tkm
mRUUiAoD5bCoFc06qBU8aYv3M+aVR8UhsNaexn/1tBWaPbxCCbUT4MZV3v3s
cbGHrupqPLeFMsMzCA80jtVMx9QT3IPd5suOd6mmcXSSko0PakuhhPHWtjGY
lsM/O8xiJnlV11Uk+3QlIG3Olgj9/8aZBvJNT/HK9oUic9Dk7RJlE5H4ZT2w
3CJo8UoYfxtEm3DrzB8mw1dqx84lgTJOgXwaP4f5cV0Ykv4pqclIMz2czCcl
a8XZ4DmoFRPowYiVCYeVogC7LfWgKMI1sDUIdvbP2bqS6sZiHicllGR4ku2Z
mtuvbxxgNryQRC+wdztK+KgOiC3BSGcOawcB/CB8G9VqIJ1Lrw38euVzFtN/
ymtXvrG5NmmDIJQS7gGG2GeIffxZ/7hKAO7diBfkDuhMw+/O0pzCHNulCLP0
NR3QPl2VNtSoH8zx/8v3y2r/UTVGoFy4VQohrgU7fiSXnrywGK54N4m6Fjjx
Ku1lRWX/P04B7vNIbICkFWVghZK7JJ3P6Xi8gVqPV4xP2MMA5W6IK6dNBevm
P2MFN8FLZkOvqCK0G3btSmWnDqcyHQWjXYisjnzzH2pIFxY3hFFT5rn1rlZv
naXl7JWLQng4qW18lbaK5LomTVau31fPH6BlKQtX0Npwj8laz56oRGunX8WF
Ct4yt29Huq070NDWkzeGQOiJbLkn2btjptv6Dt0u0PMDqFlRmV72eFqDocA+
xMqkcdcrWdzG9ml6JpYfFBJ01YqmOLLyBH6dVgUCHKrdC5LGS9+sNAOqha+h
rtzcVPDqFwLpYNoMOpv3h3nxlLTL9xS104y37tgoSGlbqsh8130/5MkeEyc4
HxfShMx3F/g/j9UlV7WtqYXDNfAqfzaylgjYPnCgQhKSDUs9YHekOsXjQyan
nhNPCOhhImhYLnTrJREn7hize6/gxg5GxXNO1qwTmSAxEwTxasrzKSD9Afya
845OOGLrROgGtaymgSHqRkPPUKdsbN+bq6hHXzLRWfYf0j4OYbIqsce02Pm/
QJgqeAfIzwCLZAZczaFAmnZwRKtduiSDSp3wFBJnEAuVGfuNCIrBYi2pyKj7
zK9Yo5cszxjINjr5reM66jKAHTyB5u25nAjqdo0mBMS8Kn6V29MUb/8lgY2r
d3YugLPZBuJJxdgRl3b9eqigF71U+C6NQQDTb7XJAWcNaKGfdF8Ue9k2w419
0OoSI2TzUnr2HPUzdXmrJbQTcrjme+IpncFvyS1tAi4rmwq/927VYdTxKLFV
sO8Zrh4QB4grP6qtMXEr6sWE/1qQ5xm7u3Hc3sGwu895k+M3+OoTt+aZEf0D
Js0buTNCcfyO46jVD8DTRuw+xNnUuOjetWhMzPStWnssrydNwXu39Z58khXC
rluyRlgSzKWcVOaDBkVy47Um3k91WTnSgZWEpEmE+G380s2uKFR3v1U7td7t
jyOIDIdEkGA1SnWONZk6iY3G6fcbYrUlPw4uFk2/8uwpcHUoTCuBDy2DiQpF
4uowwdOBf4JHf4W4rT1onKOY5tk/vlJpkkvZos9sLJPcFh3NR/pOZgQnNul0
fhMPgz0TiWXs1T9pD6QyKyQmEfQ+TSZUkoK3wfWlPfMGn/h8uJokM5Ls3Yme
qE4OjrbrrSDyHtZBtJGwfJVyhz8GmmCNcpyBioO8ax8Ym8NJO5/vU6/x/CVm
EWM980exUrE8D9y8qz3yfYOg+TgWwUY+IHztuzA9vvjgQbc96VqIpyMaoVVi
TVJPr9lHmHH9O6N0RT+Xp9/38B7yiR4t6LfRbApdiDcNH7fOxx2pyCQH6wAK
7leU8zlTKKEd51plJfUlw8z6mNRKpwHQF8CHiZzvBn/s5Svtw7t1YsH8rcfT
k8Lpsuq44QYB5OX84/9A+EowVYsYVP6rO3biFIUGUUIa/VyQVEAJ9hkwpyQv
45XHvwCFFThCllMDceDTPLeWWWJ12CkiF3qiV2ABN7z6H3UwT29b9gRzGfZF
FDHw+nM9NIhLNvc2FFMKzjW/QRnkMjB3NxWNfh0x6y8uGhPeLNNUKcq9Ua4V
v0AEhaWHzCblLkCvNYApdNvmJQtKASjpVESF2J4yi+tiVqsuB+Ve0AU15Px0
gJh7cHYT70sKyw1BtTUbf1j+B7yvg4sSc9mB5p2fbUfet/GObwpXUFaHNfY/
y6PYYMU4S45jrrWBcjQyPL16c6FpcBw2WkahE3yu+zCKuY70b1aI+3QWM1mX
8fxqADbl8AtcOJd+aDzayvcRG7BAIFmvbjmHr5MtGeZXdz00a9ytSI6gZ04U
Hg1PwIVOFLUl3/deadYXjsyUUHn9fPmWFsYAWD7gHzswJ4AurX8tw+Zz/cp/
WMHHYapQSPYUaYe5NiKWoheYnAOkcvwjE7BOPnyWVOk0jkOpaH0R34gOAXie
aPpADZeoq4IBdBYdUeSv7HjXFE+IsbEZdhn+USaIymaOzgTS8DaFaNK0k3Mm
cXP2kiXtORTaMgPANjmcx5A6CgYufQKVEee4nwMWiU89lxvLS1R1cJnr0xjh
PO004TTnzPa0c07ObbsCRUflQ/NNitjHwLcb+WrfzScQqncRCZH2yeB+9JUU
cxZJ0n8PmUTCOlf7uevkI6tjz4UuGp8XSO0wag3t+by+LkZmaOdYUyCIT68A
wwB/COd0CKSzQBYb0tvC0iGD7Hev9oWE01MP1JIs/C/qiFnXLlYYuaQO80WL
6i6hqp0OlYQeV6lf3a1vP7PEyQvvZBWJM1nyvVARQGgXw4R/VPRgFVnouDTp
jIdK5/RPZzm7kfe+4gnOfJ3tVmbBbZU6+EwIU2E1ZDohP5XTfClipHJlTeDn
xiRumzzNHYbtSwuunIWiGIhi7qT3XgTMir/OFaCuR9GKG9TnMJvcsCddJUc0
NA0Z5nVByCnxgE+efIf+7RM5G6gniELQ9U+Rjz36LYADzEhAl0vFWUaBGqg7
Xr6vrjU5vEF3P4SlsASJaS1+R7qd/RUlVM7CGWwSvk8gT/u6JhPMkrrEVjuq
gQ6YVurPNTdY+sLHHTA6esM3cKGDbuLiBZ/7SZUvm8n9XGWQlqkRO4FIwOPP
/9wEEhd32L5qwZR/oCIGBtr/DtdZeEg4Taathv3Al13aRiA+2QCB9E9OCj6J
zJ005YLXgqf9sKSNq4Tpp1R7iNmD3lhmunP1ckMi9ePxHzxuMporGbP4zNTs
r/8klFoGsPdNNtmks71Val48ENedJ1d1HhGudS/6+AV6es0kN1ZhjGazRXTS
naAq9Vu44cYwvC31esBwZuFLX3NwqFm3N7v/dMg2sntyUnVv6uoX1V8ftEwf
wARwvWP+7Dg7zacqKslDjmOEXjbvTBbzHffmPNq6phA91twkFo/S7AypaKpD
FQRyzI5GDTHr1kX56JdOfH4m1m55LIyoLq2ke5DOGLc8gcoM7VC4J+ppOV6X
2DmveC+IAZ2NcgBsl2i+HfMPI1LzwgGFX89dy5AdpxWAiDD4hak+cD6K7UU2
u+P8lKG3nt2P/UQ3OzYBoep0hvbjs+oJd5kxX0aDvFYV8avxGC8D+fl8dtAA
c9/miMoxhVw1XHSuFXXf2Z9xmDsB7irrfUm/K5LGtXih1URuR6r/L+FbBujh
L3LBzZkgWaQVkzQASE9JHG8WTm/5Zs3kLZ0LKwhimHZrbay4dKyyIecY02Hp
jJD0+CFtSd7Rp2xy+wzapReMxV141Xzdz95sHXuiVHDYu3b15KoaMn0QDB+Y
+XL+fUf/xjXmX9Nrom3MpptWc6DcIhAPwrlmH3efx8l5cQa0nO4ySQ9gTE2O
CbH2q+jl2aNtkF1KOMYv6+fOrlS9RNWpnNM4or78SZF4jPVsvlpwLGYLhIUw
0QBWL1ZyFxR002e7SJ3SPJHeMl1IS/9YQ3o085SYH/MFF9CohXA0tq5oq3f6
AhZf5+qe3bAXSPhSif55E6Cx4Sp4AnA4NXVh7zrhwMQcAqOoPO3JUDYNCBhm
gM6dvOZ+DojqwZmoSJ6gomRKzHOx0kQSv0gOZVjZy/KbBaSUhtlvfvegEsRS
jZYxEE0f1KbZA1miUR5twohcMPMLLSCLpOjneaoyOyKFKkqE69O2KKMYZwXC
s8gNIcYz1gpLYLO6pYw0eumvgVbJVcjXZW5bTovcuXfUwLJoMvhsoncZxcR+
/tXAdkzz30AkC3/9zisbzQuzBRtb+vJbt64jWgmjjHaNewROpcFToZeCUrAd
B3Rstso2EsW5l7UppUmsm8YAFS94V61cQzPaQpAx06A8UD02p+fvbh+F53X6
yRkX1ICy7BdhQaZzOlmt1p7VZCrmBE5+XFFQ+JoF7OvyLBWSqVfgkYXoDDvj
WKVmGp3yivwKCWtY8VAzLTEpjX6SdaLA3t2pBKxTQBcbbGJq4zakwR0PP1Rq
tJjX+3rwHxaAc7FhyK1G1LpOra5Ac/6x9Yh9W79B3aYe9o41wKYj9nNoWKCz
7e8rXvuCEkQlJn+adH/xY1P4VMSHhr+LMpGDH9MMRl0reJna9J6kRhBe70yZ
0SnaYDBGbTRpf9aT/43xz4kEcSRjrdKczo925ZEUH1vy51CsAxNVNzQF0y75
XoMxeyAQ67Dnl3+z7DcYQ83LExMpRqtQJgydPR0NbVajYOgrJU4u0yvRKuef
SxYzWdZmr7wD4MjtrUmHSF+Gb5U0G4j3iQP0xHUQOQh6Nbqv+sUz9LRpMAAR
6wLtuAxftY0GQFxSlgRj/MdotVupBqsHYqLbVHA75AYV3/w+JXLaq8duZm/Z
uizInAD3WNlLxZUC5X5RdExJh2EgvwPSlNlD9NaCHxi1cDwfdIARYmbZ6uk0
tV1jF7XcT6GIpe34PVbsao9Fq7HBkzeHLaqiqcaTjTQks8Q7WphZrqKfFQY3
rSZ6GOKxQgdcrwrtoCXjy+h2uz5p86Y1U7bhB0u0E+SzDha49Io6zblKQl5b
Wd8Byy9gfGVuSFMTZNfOKk1NbYa/OXaxewtrHZu7gtjvfRcpt6xOECVqP1ng
w7d+sRmvf+lCNj6DfPJpC5rt4vNjPaN7FZQA8zruTGQBeRyV8fVl8g8WolQz
3FX7yphr8VHM+telRllHkqh/qwdmv54Lf9Cl9n7eSCBMceS0wFovcjbJQmt4
b5LhjauSan5sYT0/LQitY2OClqYLR2VHGvXgZPMkssveskG4WjRi4Ec0vZee
lozeesUT0MxQoIUNdWyoNKIHNWUmlge1/OpKcpvWbnYgpB+fMDAS960pN5hN
GZQ3VGDZhoWscauzT3PU6g14kQdcY5xcCL9sUF2OzR9/coPYt7MLmbiFluNF
4pqo744Vub3oHuttO4Cgj6/FETS94SxQWAhL99dIH76s/WaO6ubNC9zl7H8A
2zIznYq6HK2Gk+yoMj+HCdCgxMnxunmJKW6Qq9klT8i84aoHNPn9qzSDxodH
aW2vEIo+ow4CxbQGq44v6h2YwiSUrDoa5x8J0Ho08BOys3+vgE0yqgxD81y+
+Ol79/c4BIvhW+XkT2L8B87QDXEflgSPLx03BPqrquoXF7SEmL2NDdhMjK1Y
pogJCkLv9Wt2Go33I4guFpHP2yrLcyDN/DHTflqWUSOcaLDFRErIGUyNavj4
8xzqdP6yDLVAyKzZlSfW2Y5enPc5hAMIiEz5lyXTys9IhCmz69Jykcns4FLd
JcLTm72fh1sj7PMtSJb1J/t6mIatGVsAg98Xmq4EonKxhzg8GF5l79Nl67Lb
u41eGz7KZ28T3xcIRjxltcyEFSydb/s/+HpW59ImxWxz17KKiXbTmkGfxQeG
4RhvPqJ710yYnBwpe/wzTfVU2pBYXLFVtYcoWsTaD4RSjV9vW5vqsyzgDuma
7mlkHc+YOxFsoCt/OXd2EO4khohdZ2msW0Nkvv75ekSM8xhmtpxlYMHFY0i5
H68pE7L9HEH8ao7VrQQaaB6Qk1GXH4sPLdQ+rYdXWZzD1+NJPJz61LB/qhI6
/uGXyXK7DNOKaQGs2fqsSM+x6+Cv8g+qbUxULm2YIDhJ0fjN+BNOCx5GfqBR
qJeyzdPJNpeP1I56G4cgtao7UXEAUDkESLomfPSBtaL5wCUyRqQmi/HniVtX
if30j98NN++VVTISDsbPl585KKAhvclik5bHGDJDtxZ47NuQOgfIQJOlqyMU
jqlFVxc5zngxazYTX0taaga87KO0GfN5dXFDeQ8SaGZBTm4GI+HjS/U74iHk
X2VF+f1NFXosYN/lkedvJwAfVgeTxvphbO5HmhPjKOGnli0vPpRMjN2QpfYJ
r+Cck19a6/dQnVvWiwdGx8Pmahbi8ZSbsN9tlV8AwngeCp5b6N/vAlv/SUu9
LWJL1fPVNP781BwU/RwnFy5Z8rFUgpnVAQ/NnPUez52FDddv7mbi/hm3bwQg
ColoSNrDtL1Z1fqkBd4jJJ9JWYRvSovLnfe6wObfdMNsBh7bsXCdnMUp62Ug
MKSWGW0ZHzeSQODuojUeCmbxFlU4G1aSHiYC3XEr6P2VH/8RxAlVH3/79aUg
uZm8hRbbe84PI5JbVjpjctkLcFSs9U7ecc8io6YlssmY8wJWLwne86kqvhWB
z4aew5wircOOn6Xb+jP6qjgc7omtJy9UFOvGUq8EKLBGwH63hb3lOnEUj7W8
9sRyNSYO3mXVFsjIuJBHMJIiwqZ96Uiwqij8L1ab0hkIX3CuBpbJLrwZ31Cb
pA2pEdiaKw3BHFJg2/8jANriaesDCwQej58Rv9jEgqb4M8OUXYcRsJdURqsY
KOxFpeybLudEUUyUe9oSwzJaq2T8Dj2f/1qoqN/1+3eSUFhMpRF0oil5dRIE
+FvKY2iAP0mdP2W4kz3kVLoNgqsT/h3y7nWCMu9WVYuHlbe/seJptSCCrRqK
WhMVgQm5KRUlI+2aszr/VZALSRbVNhHyyEB0KfJoUMX5t5DZig4wWkENt0je
fUEapCgW64zh4cru7ky3A870Jo+Cm5UiwUTYHoXwWqwibu8iNCA9B/VQLTI3
+smTy2p6sot0q+Pynnp1cyw3OnBHLT8i3+ZwuuEjLY8VJFU+XNXgVWQDBGYJ
3U9OgCSYK/I0url9fH1HE1MkH6BbKHcNMcSy97nVzRTJby9t24uzDmDq0JXN
536Fw/xsvOZmg44WEnYrLCJE/rKiKZcW6i1eh8Gx8YKZXF7Io9FX6YdJQ5Fk
mD1KlxlPugTHL5Gh6EibbEOWfK8k/4ZGe31x3PN2aqiiyGZCCSHiiZAH0p+b
szeA//RMeYCBf35BEhVKkDJh1j5Apx0rUG4BzTOVwbY8Wb2x6sZTY39XQGOk
tAYrSPqE0QjGPs4YZBJJmyTmOLvDLRYjOY/844om4d/Di/SP9/KemWNtopga
mBH6RcK58jpv5r+LaYQgm4bEYfTHUk2/xkWBtoYcDTPwR/oR4xD0J8GHFscK
rAT3KFjqtEhmc46TavqXzsXbD2skcGWBUeVSEFPUnCodUmbf2MNaQ8U4DVSe
F/YIKcP2rEums1hzfocl3F9qfPV4jubuecP9SrkVPtStzDS3ZFeZcaWpdu2a
kyTm8wFxTgCREEfqRn+an/tAzPEqIeTIQGIsViX7MXVZueUsLk2Lhk1r1CwF
RGPZNMGC8/uQSheJdqmDHE7G94BBxejw/6MWsjY11TGYLaeHG4p5qu1d9WGP
15Oa+4GgnRH0ES+z/gv+eSAKS67AzsvHuhgBweSvj+HdqAxxbNuZLR7xY/ff
72VdLl8ATYur3zybG6f40kZ/eHFD219cF2epRt+F/3WZLxfXveT5TzAi8KCz
AdDGlrjfggYqYtd+N4mBmWv28EhuRyLu+ewRzA/2jSh7PpxEAvTvoChIMJoc
ncv0zyp6j3S5yUdE/jUHo43Rd4oakSGyLYbJLzHnwcBDhu/ouikQTJiO0GaH
VBL6+iZs8K2vEoB5Vbt0fdo8X0Qxhott0ruHGfcUu1ahvtpk8gweDPdFwJ+D
waE6Gp8XsnEvSqDQTrinUDp1fI/aKjY0Serc2MFi9uSutTdr10AI10XlAY1K
sjObsIfPpk0G2ju9QA/8RWKwu7JGAKb0jrPaeeAbmcpqy0WzG4jACCId1AP5
mDgi4acgwUuRwpJy9wn9rprTxTTSGPX2jxd/Z3coNHLEUMJ+lU+7PGMEdvNG
dElgjde8+IiB+fvDBNP0xFC2sNIzndyGHvS90dN/xeThZ7ppv8qYojWghVO1
UjWDol3CiQjmbAihgugLpcskTW/ycwM/+gP3wndrxZu0pzR/nRe7O5EWAVUr
u69Oh82oU45DUwekRgpzl+eXLx/+W4qXJTg7ZK6HHYBI5OfwhdeHzvLxD7qy
UX3tJ4BD8Ku/Vz5TmNMMWToEIyavAw6Un+fCZEavKBXDT0PlaAvDcqXIEmTs
xY6Sbhzg4E76RmEGdUvJEtp3DFWS9pMl7J/tucQjGojTb3lIiVTQ9yuB7ACb
a9qAJA1HL+Xx1J7Z8smOcIt8O748z88facDjSn3TFXb7a60gaqdw9yAOMQbr
2RXeAG5w9eBAnL2elPSCEzvszJK+F/x9w9uGqtq9LCKbJxJy3edaOJLkVBB4
9gP8kOJBQR6wMzOnWERHCmLFul7ih8ObC3MyHi9c5GGCL+l4GRaErxQ94tQB
cyDecn6aMMixKdoqu+pBwHTxrtnT0vz1fBaljRrY4kfHmADRE+LNTegOzXMu
z+ilNkr+GG8BXVougQxn2sEfXDSqSKECTpx9+qs5/AdeVRF0k1VR9wUJC+Oi
meM0Z4Q9iICD7BrVctEzve/wei+1peVTj7JRbHOv70IUe60VU+oTsTB5lB87
8cbVBuw6SYzkBITlsePxEbO6gFt3hp3FmsSAgPoebfhOlfq6mw4vVjgdryw1
TvLQ+LT2sSVZDclqOkRenWumqBkBnHaDH462xUGPMhfPs9wqj1L0sua3i9J+
UDDzVvDHPISLMWAgI73vWQtMBVCuNB6RyE86jSVb2LyPDtJb8IyPhtTz+bGV
LoOz2AC4AENlsEqRYQSpY51UmbFaIq2ADC5k/BOj6D7ZMA7YTH3mjm6BLVt8
m5g3lpmdol34wXJP/Onmib7+n8UIngTEESSKrwJrv/x4Vf4lZVYuaOM53OiO
n5FHSQslxq9t9pnxDqodg7AXAMG2xiVYOPcH4lKV7pMtzs6wOqBSmOuO5Cws
tu5r/l55/4xM2TVU9r1lagkXiXVMnCX1MRxo8koH7xC1PqRFMBa0wXJLfTn1
63MRwy+TnSo29V2ttpnqTT5QUrjiqzgwDBDThiQpqLhKX99LoL6eiopHiMEt
31AI9GZFCbiLBudwZ7WftAXwIY2KduHo4b+DL2yUthnSg0XAP1/tnVqez0Hd
zglnFFnhKsL0h32zZ5hXlfjmvdzGUdjBFtiuQZdd4ZXR7a0PVCMDNKxborZK
UUb/pJZdv1xxg/Iklnyfn0b9YwC6MorkESsVllC4fwnf4O56ci4NSM7vIE78
ioL1VKTUm2pjlAYJ+uirTn7qWwec7ukVhds+aOgFkF4xS+BLzqROZ3yq2J2D
YHjpkYthUSkIFNHdCuPvkoyDeqFkHNIQCXtATK6+hr9UMkbn40A4Qw6wLAgJ
RJA4C0jN56Kszih4uJouuOzPJi3Et6anyC5KfmPK52kYkZpZHhHu2hlRBf0i
KV2pXHpM8amAwW1qzsPWBl/j4SMRuQrgzKgp6AJTPhjbbR0DY4g7z+jW77CQ
3ZoBWFgEmFAyYAO+exzj5q8J47qorQGGWrR+zt9OMUvlMhz81HSWAPOkYr0L
MQvBTTeZ7nCZa1To5E2NBBsMEtUEZsSAEM5EdUS4iVmrLSklrbfa/QyG0Rqe
gQMyp8U0TPktJ5SrC/A9k6eJSopr26RjU6Y0lBSLWnug2ERjX5fHH8FEPXeY
wdd3F6/g1BZLwcZVFYQssv7rrsz6Zvdplt8Q6pAdg73NXHSF2t2b7KC0Z1pd
i3WiuEhUrjXkV4nDHhPUJpukB+z+ljWh5zOlRVmeyHMU+Mc5AXXpvc3Pzb2B
tHps7kYt6Gz1d2fjUOTZSlGXnfnB15+N87I2eWPU0KAhjIJU9gOwmMoUHc8w
k7M2jun2LpZlhjzxreYhGhOcLZ9ccrkLafRZUMyYeAjj4K/+Y5ePv6egrpvx
chncpLBc/EfDlkjNW6DfXuFjhPxOzsxT70Lm24P+3Rrfuh/nqSxg/NJASrMA
ydul1ItV4oFH7eXEFYeX+6hayzAmA+AuUXhKyDQVAbxc+2HwqeqD08uwIFfZ
NgaXfAI+VAueWW4Ey6N38deornripdkvDahNjTMvpReFBJaua2Qm1zN15jP4
ySWAig+Fq3CbnaCKAu6bMiUCSygFYHC2hjHCTsNjGgZBrk1X1Pa1Fa/3MHsR
qEMs0wQznLmMekSiYYPKaOOv8J4828SwvY3LtYlEHXP4Eqwb6BQztwMF1jMB
kXJlPMjtJQi1j9TYmmMTzO24L7t/tWjHReuc4XVTpoDmqpWqtkEY/iI4Z//X
gmDgmQFHpEHfePTgSX+4oXFyO/Enwr6+8lytKjWggZ3kTPomZe/iEQv3naAf
TM2QZxpg6yiuxPdXgVBL/2NBiX25Z3NrNijOiSsEvPveQ0bEWwWEadiCwkGk
1h7EZJSCnqm0u7j7rzF95khspaArI1YEU8ArOssYsoPfecz21iD4c4EN6gMH
UA6yBM7+OPcRjQ4IBozq9WHfebIEXQuxl/IcngElcC7svEqM+HOu6qHuwEgR
LdAL40l6Jbk3S0Y5ZVxY7CQzs7x8wZt8daXoaDhkLyjo5CEzuZ5Y1lFfZ4F3
id8r4ksDOMIJ8zO6gqXSRAYXuZkn5vyaFnaateiHcWjMxNUtDLkHUtIH2OEt
MqngK6KXaHCnmMVs9+t4NciXNAGmB/Y8fKPKe4rh2BrSw2/HHJj6bCASt3C2
TqJZSSVHE4+03EJy0oxiPXCuIzxZGGzrBXyOtRBDh28ndjsIJXG+ws3ViWao
5LfgO9d1yI1Ws1NDLC/j+347JDntyXSt/xdrvc6FQQSdzcrLC9lY3ZOJr2T4
sDYUdnZoIyWqgsh3eP7W4IjFB7qYcPOiOqx8v0gg7Dywa0O/zOnz06P0Q27q
6Yef2cFPi5aW+eS18BmSBPiAHm5mqAEn0wxiVsp55dByarvbNN1y0Dr1rYID
4yVZlb5pxapyqp7I0zpBrCbHjsOit9Rwww4q2Bqw+mKZN6RHCcYzL1DmKkXq
GvPFCigVPcdrhPFzAd6a1ayduv2xJC/z1L5Gqiy3JFBjdZ+OKGFell3RIJc3
Jm7/zDRpoY0HqrK0Sf83i0g71+fSumbKyUh/ltmpu1vLpTV+wiS/Xf/kQqE6
/uUNPKJGO1KOo3P7rAiAwd1HS8ErRbqT6x8sVGkq7hmX93cjnV3rQ5CQr/pe
2ma2dfvyrxGIOiBxwZmifXB/075ZkJgtMyHW+TEBzlffpbViUtY0xMh3qX5e
C5w85FV6aroHAl6bmf3upFW1qDS3dnoKu2ff3yfxnquKsEnsi4EJftyatWRH
m4UmmRDlioUC2RwzU6Gp6nhYVfDnCrDfaMbQyIJuC4uv1J+Z6VSDLVM8f6TL
4j0T9X6rEfJSY3rdOQ0QxJyYEeH/1ImLoPDLsxlf944SGA9lYNyqrGkZU3mO
PWuuzR65ZoB3Llm14jCCMY7i6Z6g61U8B7hxA3yFDKaxXHmoSeuqexSQDBt1
IHGoP5zNtCqZ2qEYp7rmSppUsJ/+xyKdns2D8Gx5pmEnntOVUznpehh+Ib4l
J64d6zgsH5aXI8UZDmxuGb7touuXhreq/RaqUawu1YubIT8atQTARgI7VDMx
ZjLyify8Ca6EC+z+ybnS6lDQ/kdq9tdlZ53D7QHrqt4HF5qd0CJW5cejqK2R
u5M55wUdyxUt18LYUt9xO7wWZyLYrqZP8kUzRyjHT1viRRA6VxD+kh98L0Vs
e0uP6Nm28Spd8OriQeDqhoUJS8VIbrzBoKodWT82VQ0HfCDbsYVhghUhMUZ8
WQW0sPqY/SPVEFPCMFIlXOMpPgcXEImUJCT4WX5EU9KELrQ8acsLYVoOvmXq
5s51ueHWni8wr++bd6cyJ1xi824weV+O8vXx7AkNGYFioc1ryDnmhx69gUBN
FdrGK7MnT4sFiKvjZctyCPR5/Bkw+yj76nwVNebHcLSG3dgfjIULWZVgEKk7
aPXSdDHTYH/tM9bQDnKAfQ3ifE6MQyl9D5pO+FuYAo18tWLPVlCBWeXZT2be
DOpxSY9jN+Zqe6TZYwFGbw32WiQS7R3EUfPtFJ/yzR+TbNQ568/KWC0FnvBc
a+QKJIuf1s3AwQYk/ljsHzrYikKnp6MiFuvfmyNZcyr/uBNtoN00Cb2jzMJl
73PIelFnBjgJ3tXXosEKEHvQtPjJP8Imt1FHG8LmnvXekdU/kx/EJjPsTu3h
MxN7xCs7noBj8WFQm4x+bb0mI6OCvEK0ghhAfLaKiANzt84nRYAaDWzvyFJo
aiG5nAnKU1oAiI+zs0yVetyCjd3CLyyJHpPS/ZKIPH8VN0pYFUKUvC6GQ83S
NQvKzwznUMiXxayKCXjA0QycIzWEoQklRZy/5P8G2IKm46GkrOcu2efCytd4
Q6vInjoiaRAeu77zo+y0k2nKDes5iZn2PCTYdqQkpfilUimfZKelo8enWzFr
4ztQy+0NWKiiEZHxIzSzcxZCmA6Cc3jYRAcArr1zhDXIY7jNOOGeDdOKUsYp
lDE0+uGmLu9GRWLxsstYYk8aj42Q45SqXBbbPBVOPBYKYXNgbQ2wAb3ZKl7D
XsOjZNBd3PE/6Z9DoYpqi5tnM4fS4h8Beei5xFaUbrT68EMYxR0dN6t7r4vb
YNf4rIwa/+oJaE1rGuD9nsTawbR52XpsWLmLawZbfkwOhf/umDYNxH56zMIB
pdIjCtydvU2gBHFvjm+SS9UaPaFO050HtOQZD+bpzRyHKbHEApjKtkBFrCyJ
iBUlg8vEjE4C0liRj0TGkPWFdf+9pJsGk3xqVnq513yPrWttzwlnImKCgxLA
h3FLUs2I0hNqhjCfsQZpq76mIRyeS/f9ONXRVY/SnSVUfXS7b4Qbh2bkUitw
CYHKItYr3ZexUGeMzM9zW82Lm2yQt844sq3Eje7TJUp00cEddJwgs5bbwGdA
tRaLakQL8yJRLTxPTiVYjxHsumx5shtX0sjU/jGE7kM2xYQJZlrqRaw1x4LY
OdbPACuKbQXrKCiXw6u5mgkR2d6VGCiq6y27XipEM1MLgINpTGNfgWQBhpe7
p223tvvg3Ii0o8pBREycrjvh7ee+unf21ESmhFCGH0MlpsgkSVCDIvhtw93s
s1JqsAnwXTukvh2h/bp3h1quFD+3ArayO40ZtdzipxBYqm0ED6li96WVmt6r
43NB/Az4wPHQs9HSQ6kr8MzXjRIljFJPwjiWXFtAUaNwhV5vP/Lj2LUQO6Ev
T8DRA6E+kNjplOLLWDV/XMbIbPl3p39yvJlzjHjCXF2iV0EZFyxSaIe+y71d
iRJqAJP4RLePVw+OG5cFvDBQvowB5U2+55UjRGLsEC4DPLoQGk8HqThqc70s
KOp8SSELCO4mowzG4plrUgruX/OmoIaU0KDP1s3uKW0dthPgwmLRd7+3+Pj7
Y0ViwK+OhcCtfNt7glvGtmvTzw0D2/W/2oEpyis5pT2z/wjyoZGIXFL6cz5o
MkD1JCikPeEYkrde1A7mkapg9SZ9rUKP5rKh8sGZPjd3cmDxwW+nUMGcwtHZ
0axqFpa9bTIibbv6PDBehVvQINkVeS7C9oX2RF7tHmEORkIRkgq5bJ8T8iqk
t4KOOdHrxn5ISQ1uQaBh70OUx6Oo4rNHA6ZAl5bw1kgaAeaFE3p4qWLS5zcq
pwIi0JgXaac5tOKX+WAWhPn4AZchSsbpUH26MiCBW8uMxYpI3E1kRkrQdtHI
jlgYupKNd9BVun+1kbVUv5J8aYgJfY1CdS8kYGuKil/dJZ71wa3i/VbmLHxx
9QeD4+JZ95dJ57VUUiqu9HtPhDuuIevRWOgt+l2NJwkidhWRc7s8Nl77w0cn
oBZRdnwfSBZZ7v0TVQ/uzyEhd7csYPdD7HDQVkJL7zPyc0BcD93hbl9ABcCq
PcKrduI8HJm25nmhKrmMqqMOyxUJA1dQDbgs/FhlH6t9nCTe5aLrGiOqVCKt
eTX8WrS69xzz7XiW/HLl/QjcyZOTkhPNzEVVxnWSptgE08/myOnH9nUUgyQQ
rTLvUlJ4EvtQREC34qWuCSQqtworAEr90PnjBqD1GGmfFrlSPSch3y4HCkpH
Dwjt3BasF79/l4VT8FirYWx5i/Z7FQgTf9F7/vVYDavotI89KQrDGeUerhe0
xZYHfKs7rpnSjkj1tbd4omvAp0U6+FZRQZra+izM+Y8iOaMJgQYr2o1LosND
9BJyxFfeNVzX3fXkVUN5yfSPv/EynUXZNWAMekOJyzel5GE5lmYnNcpjOLVo
r3lzchbnKaIEkyhX9SgXdtDh92wMqQ+SY9l0Xpyq+m7lDuI8Ig4lh0FuUg+a
+EPt1GczaxtmsqZRKjJdWsnqk+lQlg0hVnoQyMVjvRsLflceHwfsL7cuqwHM
ZQg9+Oxe3fK08K57RKcnZz/ovPdpluwQmIelbOMBq4AsJa0HRoB4wMHlPy7p
rFy0+hhHr3hXHkJJiJCKuSgxdFY3AmLPJfaR3blbW419JLSbUivWBoSpWUHE
mjtweGrmi7KeWhEvRSYX9XsgtDquGvfgZszEx/WnnxcEYvwEiaYQiDN77d75
xq0uxwZsPw6dHBzJPMKPN0aA+S98FAVFs8qU/31EU2xbn78bs39PR+mJQo/d
Tzi+fa+e9AjP+XBLwmDooTuNwE1FReaaHJzQvlYSRtYwnKWpwXTslv8X9JNQ
ToUB9eINbUeBY0TfjN/2WKor9Als5bMQ/EWWny6jumrjVMSa+a/5AihvfC8A
hRjLFA6LdIWKl1Fp0q2DLGHErjZgIEKIG+K1DBU9aMNV++avq7qVH+OKtuRO
cLgNvdjWwaawuugR1ggsgafT5gHpyVVxQwkU3opVwvJXnR3U8kQDvaJl8yJm
Rtvu/+jn0CIBEG9RK4SeuliPP2uZs1V9eUJe3Yw5H69EtjQButmZADNyOgeB
51F6PS5gUnSZG7uh0q0/G9rOHKOIokhIW7kVvkVgHRswSDKyfhmxlwU/Y2pW
SmM/74wdE2XNzGkbJS7D42mHslJHdng+DHy5NSsMHZIPyj0RmIahTI9GPAHQ
qh3Xrk9g8S5ExaskOQ37vXb60cg0WDU1qLMFG6wbht6p3zyfh05CD0DlL3JU
+OJxETeHpC0RXC+MOwxRvGZ+pi+BTbJroM4PO4WFAl3ifwSmxeYVlpsyLLTb
HtoEwDmju/GemxLn/r7gKVJJkFk1l/F2mn4WbshKeMcF1XvCF+utyQPw/y5Q
FCftQ25ch/Xpc9uz3IE6FVplkRH6EzKZvmLeemimlQxIdLXHqnTHGf5BjPiY
/rBmD1qak3jrk/wYjztQSCVm9vaASQ9s6woLciv6N8LL7P4BTGRVlmfAvFjV
a4tlG5gz5XFlUf+c5L2vtaAZvIAUP3SGatFMubH4ZQ7DeqeNDPWL+ZLDLMkN
OlzhPlUpJO0CA82AEcF3fYMi/IInHq6CtB7WWfMPtes8jALgYXnsKe0PNZox
NQeKmNpfviCnGJ2rgXw/6h9naiAB4iIpgvyxCeKyCRfcOG9EmZVf4WgCfQqs
qeklpmhV7aqVYCtRDHeMHeJ9X8V6a7UwoZsw4OhpMrvN1KwOaEIj88uDSvB5
e9j5PDaZFuXM8h/gEgZyIh3mkStDuOjpR7qjKjX58xMy+Jzmy7KfCwwApKE3
hvhWltHN58IEwSCmvfOorUCsyPeFAnRFl0GFI2KUF1fdh0cC5I3+wbEjv2PX
HywgejmprdmMPKOIQ6l+/0h00rHjKBCN9Xj75fL7h3TfhT9OusjnkSjtbcQi
Wvvj7wLrTugoSgaXW8T6BUq48qSkKZ//0h8omiwUe/McUtbslBQFqSywxYe7
i9bpDQeiBNrr+g84h7VdEiWuALa7t5iq/WY+nuC/rIZrioH2PUMfJG13WwxJ
JN1wjLz1E5mKkQbvJAMwnFMxmtiwyHojKUgzoCVJGFuPiK5xVJtZH2COTwSG
ocMTN7SfrbWQBMM03wvlVg0MhR7wVNITJIC0eCCxbvKPo0x/qOs93twXf8F8
x++NQrYR5smAFN1GXBSafR+8XjZZCEnEySkjs/aveas0IL7bygIT8SBdNgU2
APc4Eto2/Go0Ltk0di2z47O5ZPOTHRcg0TzUc9Jcs1sayyaQhog/qxviNA2m
5b2c9cN5TKeP13Pk/n8d+pJ7bWrL7AxhOy0auU7XF+rx9TJdw+aXtDJD9zKx
co26AXDttgHtc1Z9XWuL/M0I68c7lT9RWbKjkZNco3BTix8losVoxk1z69fB
s5ABSNzFdZy37FWhG3O1RQ9iAnZbjP0fikzY7L+sqCwSPeiGGOn9JeEci1sh
bsUVmkQBVBSAOSV80JbGWJxpQRbaFghEXxQ/ASVDicuEyDIhjZe7iiVJn9NA
cwG8djndk2s/rwrqaAnvK8djwAEY3zWktCfvD447BBNY0zDpoK67TiNU9zz2
gv/tYrlPtovmbVLfOF7eBhlBs5UFCL2ZIS5YqyDON8/RaGBfQwpmm+Tny2th
x1kP+durh2rfVbwoq9nNtzUY3LUtYHKggYx68mCosDXATRfPq+/oaOwUBzbt
GhwV2ybWNOfY1++M5MU7GExjb5hGAYk47g+z2aL8xOi5VG9PjPn/yL/YKJ96
HOo5H0kuTdXCn4vBabDUAvpnmlNTJTd3l3hIMb/W+iqrurXcenzVcz25Evul
tokTsrcxrD4rgDss1Wn4HAaNAgccuYAou0fizybIOarVdoPmFIc4/hkf7sWD
Z1Dyiw6jtEIWF9jEogl6e65z8NlD/RV7abMlwfiSkC/KqCjIoBorxox4axMM
UAw544VMHDvkQcDVH2rCRwK3JCI6bYFeC5F7R5MDVTeguuzQEiJz+sK8tJP4
vmEFTXSF4jFD45yymrBP7XPb+o6N9CM1E8XFCnnB5OuqW2BZqIgs8TN92Htp
Pko/NWHDL00mY9ny9wmGI5oAjhhgRUwlz6lzL78lOORlF731e+z6lkCW6w6d
2sPmM3jKAfyzdMCtDSaX8/JACYDU3yBTHcwUKiSk98UhH1sgU7BfG7AcjQk4
IUGEMezbUO9IQTp+VPtj8CRYFbox7SqCfrlKNrrGvdW7Aio97d0anlEwLaKV
Q8SG5dvYVDbjHcGE0qJZuVbzSpyjO08Ee/Ljknkg/7REWDO5gWFFjrWVU95a
8nMTnSvifOvFYVcIbTZtcW4s+9qDSqbPJq+Evt2CSHoW453dfG4fsXY+dzYh
6ukYvZ+T5Y5tPQUqEVcxM6Phy/2bHbiM1h74VretMYK/Kr7PdrBMeeI4nfSM
kDDqfs1v+WIgin29SsLmFCdgBE5eZI6K2KdIa4CvggWWaxCvnLBUxFbArfkZ
UgdBhaf5JZQk+zqefvSkrbmE9eonjWoqVxhfzQu6uajXdaOmLEB6LNoUwYyk
+pVhaLyixyOZ3mmFOm2f+9lj82BQP9SxzJNcx9dHOTAWpIVglUPOKKyq8gan
6KwRE37D0Am6ERbC9Fhm0PPbkVwwBaEgzo25KeBxwA3kMmaBeCWCTZQV/8tL
iGwzapURD9ZxfUIs/6jXwqAO8/IM6k/16c4UGTA6D5zFkuViOBWTPORkXcW4
31kz6DhcSpce6LdaLYdqpsHaBY5Ahj0w6maNNyyeU7tdyZ6lnJr8ydcx43rD
vTnhQteDM2MCOrkaS2rPCj5aEGtZushol5vPk4+tJcXfPfGn0Wo9wOBcK1+5
PkA0wyTntAmz0ESvvraV2lYy9exEBmRIR0xCTMnmTVpmQ+phTWM4KFRdnKFu
NS+scdWtSYiQ1Cctt5xcag0vq1DPuIKqR5ezltv+IToZ8JGzNVQSAHpY9dnD
r2JhDAPinkMwIOgj5MYL2Z24ovgPYDZxD0ByOAfJti6YOKGePPWINfTG0Bjw
sZPckihot7rtnFdfbLIFI/p/+VqGpm+yDlDSfSdAKyQ1Fe8/bfsFclLF/37v
B8WzGcntMUH80NxqOU8Oap7Q3mQpVba39wmstEh8wQoaHYm9rqM+2HPweQje
EjG/1DkSS+QD4g7qxSRe2Cu/zQhIJ5osF5o9gXHVjsVNvKMQljFO2ki2QCdU
01cL2OunVdspd70rG70gSt+Q9q4pLVsBhtX/O8tr4WkvswJ1Ncf6FZT8dQJa
BlwEoS9FUc2w1qjyCvJ+KjGJGZmIar4YwKdB/rHnfctXa/w0y729c7uKizfi
3BP3muXxhC33pCYAtWLl2rbgDaCNDdze0kpSwxYV4DYGdOIwaXPXQtYuQtWY
OJdp+MJAbdZhLCqLqMA/kOftuNOjFwU+IoQbaTQY89Y6oeEZZedGGVr9KALc
/RuthcYqFwVA9+mPEFYtJmAw5rLiK2O6SdHHn76NqF0esR5MXrfor+GxW5qr
F+y7P08X2Z22q31yPozgOHLjj+UL4ngSHd042s6cxnJymex1ldsveh8qMGLi
wi7PDG2FmZujrGY3DPiI+cZeY5dLalkhWipEE1Ecf1WvqeFWLC5yH0ZN4vZV
aw3XqffAPijfjMJ7VCQDzVIAffRtRNWqXEygAo0Npw3U1gSuFrr/e0uRiy1r
YXuY+8Og7dAyGI6AlYLyHmvsnxrqrFVJ1tB7VKXG0zz0EqeYRElDac9mBjlm
rW+igt5gPdp8yWNisYP9/8GFLCQzVVhU5eF+295kDrv+i9viQakjj7G1LIoI
YNVg6P7MXF35Vw56n0lGNkPw5Fd3KsFkMHjbBZSZrBhg/znO4G5HCYA3/OkT
Vi5+mOrvNFOeSg2907HmVubcLkBpXKQ8gtfdsytjQl8DpwNXBabiyxlKHkg3
x3OsFH5PrkILg4IlVLWIMrpklLPxspwGGD3E9YQ9j2Xmd5iP0T6OtXz/88c6
mHX4/e2LAdEZyAWcYig8oyDssRdBEKO/YoUbNEGFQJqM8qiH9dQN2CfCSgZz
k5yPgtv1MYtJDY1CvYZ7nwQN1kaBbtZpui2AJgcq1730bsBSBPgHhsuSgCye
YVtrjvR/CD/yvcYDmd4fO2xJArp9LGUkIOI1QrY6xkO9tOJhF1K5ZrtUnNm4
21m2OclF4Zs29MwbqtVHBleB0Bjx3OnOeWct/vxa0W55eByGvUCGEBXpbqK1
57cNfEBvTZ7bAUQTuZUDEXPoLctvsnmqNwvUG9mHcAYrE20nmEzm/QmEm4qt
AUwGifuNbfCxvDIbzHL3WKOT5NbOsszCj7Nslw+vg8nTUeWJRNvjzJdXhNyU
IWoaWVh8nZtPR7koJDljaDe/mQsgosNbH5zlPydNyFiYXsvH49SsUzgsHlJq
hkHHP4bHn+xPWaqcEvaCqWCfVNekIOoRKZCw/v5JhuhrOO74IWwEJRnUeRUj
3uDrCNSBdhhI3dvdd6XykXtbn6p9n645gUrgHfJ+NeCvy3NUvtToMGzQfSgv
Yhmp4EkLjd6qEZy9FK8VoskL4ycWGZvlqlr7hOLiUMT6wv9iTsMmCXzEUs0H
Rj4tHlAfkT+AI2vwjY9xHjbvNB7+JWVXxAV7ldYJzr1se1Gob2Bl0pdNOAxq
EeCMSzi4BEz+ZnUTxowI+ymUzPy+ywbVIlwgTBMpXdGwpJKRruDDfzAQBPWI
3y28NswCN8QHKc7QnrR9Ps40J/TF1JmBHd0maLUfX3of3OLwilqCSVuZzDzf
qs7hmDlzcO/MzeRyNmzXTWfnVu0kCoNc3dY4Z9zduDfTa6p8mhEdKiCiI8h8
kSho+vJDiPkzahjK0W5ijo+KKP8ND1E3/xlw+mWf3eus32ElBxuiqmopajye
rbHsfmL3dla57pvK3qxRiS0c9nDkJvpE9QTT8isTfJjo8EVFd8qL8WWXOvPR
kaT69pJDKiPUeNPit7dIp1cVY4iDQuQnRuyMVR8B4pw9xcDP8XUf93uyiKL7
XzIVKZHkp4oV58SWmt0u7JBgduQJGZrBgqYVlGl08rzAPknq5Z4+zLggHbuF
i1ebFDSRRzyKdhzLjIR4XP3Tr4lMKdwdtXMjih//yxVimc7d4dAfifOxb+xD
UGOughQPf1Kl3ZNoJVLmB4NgnG29cpOUTsIBeYIVssILF3hnkgBD6wSuYxlv
i8R4ez3TnLsXFlfOUIqMpA5O0q8lL40ffoAOUYKuu8CxRb4rFDNK+zuHL5co
lTPcxpL5JCgpirhRQQ6rPwZvEv28hapxyBaBE3Ph72NAmDEa/vsZYo209CFQ
nKpTBtMx0uxq1Z63DePnn52jH4U1u0uPjLw4kTaYDLAHWq3PthcnnMmKcGSt
kar6Tn8EToLcKTqKd3CyYzJHYgPbdsi5tXUx3JkK9sD4QABMSfmTjrGwJYID
pUUJgibBQH903oYZN+vPuVwXG/wKT+tOOgSMsFAIPL68wjtLVkHWa2SlEJ2r
1VaRJvfixsaP+Cj1C2LeMblquE+/BARsqB7k+fLCG43qGr6e8qg7njkplyno
MxR+Ri1vVsGE4gIvFHbgedgbabEFZpeoWgoQxL1m/wBY4YfUsVsiFZOZHHQE
S3IOW6uS9FTt6ootjAdrvVMCvYUKAA45Mfb0lgD+Qc5MoeDRnxyN34uxwnW9
dSGsyEL7S7cdjJszvE9yENCDzyzAau30D8EYOGRhSB14Rv5eT1O2PaB5Kii/
8LRqHO4TdIMjUy81KWftpsdg/eDrQ6TMU3fFIuBcnF39in8fIy3czJTZDKcU
VgcHCj6QCRO5YpjqwhmZLo49ehBdhFGWyYu8M2/zNwUdardSUkuhgjnxQ/KF
pfrPcoatnU2xzuyYET/ERqGiytyu5rG1HGiwCRXUvLWZ6MarL3Zev/1ufWLu
YatrFnwa+4kw9QQRaindGhyoQ8HVuRVbXcDVra805gEwQ5O9yPE+4p2xob20
pSWGHAacK1DrQXgBv9dQJrPjn9Uu2/3vUwgjOqNAhBlIkFclrCVi4J3ZLtzz
+hFRZd3Zq7KBU5ug0L3GgXafNcqejnye8a6X6fbhL+tAOgvbn7rJFgdtA/nd
m6I6b32IH3Deaykbf6AXMRKvGVqt3P5/mh/kfWpA2bNVOcMI7LIbAgNuTlKP
jgunZrdqSjUh0Wg5QNpEspT8G4Hi3ljLRYbeTSKlYPauIQNwHJnH7Hilsa9c
cxzjfZMrr9JZAirOs9S/8rhROR3PejtcNdf22zdvfav7YNfotnQ2IepKTXey
QQBlJPV2iRfN54RSWyhpZkv+hUhSCnZRjDZ0jA02afy1eswV1Xw6aekBzz5b
7Rgr7LgJT/ELTXTVDXijGk2kl+lK7DNrVuKkudpFkgrTY5iiOBaCS2JxSoCp
XKJIxdrQBUbW/s8e33TVEslp2yC5jEQ1Sl5eNSVcsS+gw/US4zbJYQNK/2aI
cvKxPfttc6A5NkEg650vEw9Pt4Pv80UQXwPi852zyEtbKn1biW/HYDN0bzfg
rorxMO2V8ehXtAaWpkdWVTcUr639O3Z2sLb/H7bOPbV/ImGtEMggpJKGRO/J
Svw69XWSllDa/bhnZcBcutjf69+ejGmfWxvK2Ywz4MitKSduoYasQLDNKNoV
TsKeUjpFVQt5GBUtJ8OmTVcWNpprvcJfNRcWnRQpPzXGJeZ2qbDJu4buCTDt
YBR+bbhJwQpEVPucrV8rXYIF/iDniVlrBPMlTXCk47//C0QDyRZrGfzO9rCA
IgybpMmdWrF1k8bdEUdOAkOLy73hhYjKXyOZL1Z5FQP2Hd73+fM8cILEKEkU
5yAcZRSI4tOKpHrmslnw/2t+2CmC8ahILnQq7iPPhvkaCSj7e8JVMKIH5WVi
T3TwUEoJGf6nNFsFjLHOa7ZFfdSXAnjHg+spa6niPhaCPg5aKDmpC9a4te0m
L/yj8vNeN++eg5+XowEj3/HUWp7ZjedGKo82wbm+g/xc3FS1lwYVUbSTK1Iy
cvgTswth+k8DhG5MLPaFTz54nnBJwK7oaMb5W/N2arNUaqMV7eW2xtDD/tMR
JfWi4MUqnt42pOVhqGz4IA+2r3UGDGKkStti/9nYjIjqvDiJjl/OSwRU2H9h
kP2o8j4bvMbI69ohK3dKyZwrsmb4VOEPX/dY5hDwj9KjjwAjxwNLq5RiI1Yl
BEMQFq7QdpMAPcspyT6+lmEiM+8vQkzP4l2vPIJntQTn9M9XPGRBeZNBhDUt
ru6ArkZZzD4U3pZzttzom6cTVq+Dm6K+M/UzW3Kk5TjLMM/EQ/Alz8RvGow6
/4EOIStneEGbJlg2EheHhV/LGSbQTOtwoFi1OmRZldymCz7l9QEPUI3pzVHI
z22O8ksy4zuouGHyncUL61gO0/SNssUDwJIheqL009V9CzWhas6OMoHVY0IJ
TaXA/RmkmMVjnmESAgbEYvoljqpYVAi6qhNfqK1EI+hR/kTOazw11CeNJyGw
OYIumpU8tmfJSsJRtnwxVTI3mpBAJUvt26v/tSvnW+n3jb1boBzo9NOm8r3y
zAvBquQtvJJ32opdn261CQSQdR0jsugIv3g2q+dp8n5m+d+ZOSEn8Cv918kJ
Ae97NM7zs2TMNL71+WbcweMWCMST7PsQW7pUfuZ7xvsp+QIXOEp8k1Wv1MgM
sxOVwcVeHqf1N0+/4WTUhVcvUwZ2+370YEeIz4kf38JelVwYwPoLPHbOlHg9
Gnggy7k2s/eDMlk8LgmGayWzCrYARsAp8pZxz+ozDeFzL/8hvgO49ftVI1Gv
vbgOJqKhnylRnZSVBg77R4SRJR7Au4pmpplJ6R0PdEHJ4enkgzeOHNOjyanR
FOSQmjexhuR+VbaaeQCrugo7i4G/btL6hzS0KWGWVRYl0kXZLnibyVeUtraC
oauf01O6Zw+uY2NZL3lOEaWxzeyYSwfpbqviZRSJpqrsPChIsLJi1z5nKkEk
YfRsjcNSef9sDinNe3quV04RvECqi8F7QzSj4HxV7j+nF/+ZDls7NmEd9pN6
a/Vyj/IDkQxkngF17MaKzt/LyMNwxO2KMN5D0Oco1BNDcQhHUQNDBoeGbrYi
YtKfN0KySlVa62eRva8V0LxhB0L6NctuAfxgAZonPLm/6S7B/1cWTLBxAICT
t58JD8eR+ob5PgO4AqPdBFz79eQ24Sf16xKgjC9kacqHEQ06oolc3pZWjt/+
fRue99iDsEl/ZzfURWGKQmh6xJMhr9p8ThXl5aa83HXZmv15XXEwtEt4+6b7
1SADk8hGQvN3yIP0rxlrsnYvm4vQ5KEOlRWBU/yksxFMtRAyAdQxKl/6n1/v
jkhAG/s8RTkoRcs/IqL6Cxz1GCgIGZSs+Yknz+HYgkQLDA/143PPh7I8K7nK
kuD1HrvxEvw/CNQEYXz+mhxbq+8jN84EYhWuyukBoOIeeBITTSumeirtqXmd
hg8tFTkXFZt984LPQCNI512Ouf8k4QnfJ8LUqOmEHJO24taWZtdIqluTHIFC
E6UxPc1U9yVjP5EyYn6IQCbEMflc+soe1uHB0Cv11HW7CLyZmZ3XoE9FRz6F
ulUfrq29UlBwWI9rxJ6TETr6RJElkhKl0SIF/lrek2Zh74DZVNFcPq5JbloS
hFMcptixVzwGpfVrgpDt6uBt/52wHvfixPtX2DlY2s1gUK5d9IXWA6xNBa3j
7uyjpL+FEy3mWWiH7ieNgMlWkRVO4opw/obi9ASBNa+DmML3twmDuOlyGxoD
L8P91YGplPe4tMGS64uLiSLgZXnxXLAfRMImAXD3/KRakiNPlh8JlRw5u6ip
yynmtgsbZqPMNjlWZReE7B4RnWUsST9vIhydcx5YAFPEjsCWUkzKpQTqZNuh
DhLhq+RI6NJpQVXPR8LyX66MNB78nbc8E5MlKd/kLcxxJ75Dn1rcZMX3k6N1
iNpgwgQIiOv5q1Uh+4uLunEvb47uWqM6tAijzjF34EOvURrfssD/4IppWt9J
7eCAIxj9Z8vVg/F/ODQqgZYbW/CFzuGYiYpLvtWf+Y+BDj7BdTKAUk6V7zIx
ub54gxk2MgvnIT+xiflLwWiOeSTbpcz6rFphCDUhlPl7Qz1hyn3kjfRV3vzO
3kd4ED/B50YXvchFORes0M0SVC8jFQusrlPH78FI4A8i7rf1MKNdsGAR5cSb
0F+M2opIb108ZmUf+/byF47wjBgcjzZUNskH5G/T31cY+lNMSG+IoMD/v5OK
oKeiH0luG6TM2OPuguUgF7Zm9LDFnKzMZLerL3JKNqMpo9u42FRDl2nxNvYF
MqmqZUJWGm3vuAxtGhv3Hy/PabYlZ/vxj2t1rei8EHyg/Sy7LMyUUqyPhQL4
xmakszp+5dLCR2ilZ/ad2+PtBUBSyeaKuM4LKKlxy5koLiODsqKYH+xfyPjU
EW/LRvhO/xIO5gub2bO68DmO3awidFgPvgH104d3ebnFeYc7Erkfw01F/CIn
DOgfLbMBh605tl97smhQwHBCqatBwYYbsV1b1syEwNRJyvGy+0ozWWFrD1Iu
UciAtP3IUvKl01ewYbdOuvWX8okV+hMhjHt8nkYSG5weDTNrBHkysBozCd7k
+GZzAkqAwq9BipjacTtmmUEsBDvdyPrBThe7r+xjl4ZevVqQdmaLw3nquwVv
STxi8p/WXE7+esBAiD9VulOjbpTRekx9d9dbG2XaICkz14c+oEM1u9GgkoT3
vAyjIMVSjSgfP+dPC7lVXAkxRgYJtIjAbX+E0FMkQpAkvAJc6oouWpsTJ+IS
5JUA00DoUTGpR0+yz2yV3nA4s3hS7RjY61RCP8qCB+X58Yzi3abon6b/mufv
EmVOc6zN8fymIO27LNckFhnkKPGnBW/5mhl4iyHhJaZujdBZ20H4tJgHwjyr
I4fqOnWnE6u9V3UWf7TC5sk3r4c7aeFv5zHUukgZ3iOYIAjbltkz2Qg6/aWm
qPDUmAsKx/UPoiaC/ldOhFC2Jysr3Razxl8dDfWlcRkR69AUnbR44vudfDZn
FesZeUhZWSAuMbeYP4ZXxei8hj5o6Q/dJ15H00TXvl/cL6sM/G4Yd630Z/du
1C7ge14H/f6IO9qF0OQBJVI3hlmL/deA9xF0h4BsGaIFDGiBeHZUxVDGj0gb
64mg3z4jk2NGRS3aczvaW7k875tdT4a5Xsr2XH9Ozg4tZOm4DlqSWHzPRTO1
n+vVpoh76Boz4lErLDqNF0Ow6HB6Rpy49D3M78WANxfoRVF5JNNi2YOQQtfG
mHVEcGBgjgXALTli3XEwX/kUEDarGBQpVSGm9cd5FY/eOe4YzadCpDbG9YdB
vT+AFPqnyewfZ8CyM11LhjkpBb2oAqny8lfreqRwO6CQR7sQCr2fWm33uLXk
XQ+EoSI14/8/VrrSrg+xOxBbWT4hzwiOI7YyqeUJElDIlUU+q7QmtfzuSubd
nqE56GQm4o5RU5073rwi4b0M4aALy7MQudQdZnC8lxvicYr1LlSyJC0uhstt
wfwBPdkaAKpjdyNyd/ZMrRg/5GmanP51mFNaP3Dm3vo2Cqfyn4gtk+eO0Z6P
ltgb+Mf+h4NcWtWOFLo4+JE6btXhRsfDcgC55UVn0YznVxIzetNfZmH8Y+ao
9r2d3BNiGKfdHrRPFT4H6Gt0f3WPZjz8ebNDZgAEb7lsc/1muon4u7GpNrG0
ffvLYw92QvfwPWEnupBl7REwJZEkB10GvOCWkL8RljeiqCTZcbXv6/DOd09c
DJojVtMEK1QoHLJAGd8HIKABmMhjbdBPNATK505io0ObLk/1N0wcK3Rg/zgf
qCJnfHBVYO8l2q464F9v2jeLbr4nKejVoddUijTpqB8+6ohUg3nfAigBVYLx
gz/nIhR2Xk9PcHydX/io4qV2jR8pPwYwAlmywM18uMn3taVJ905RNd9qi+GW
VbD3nR5t1ALLl/a7uBb4+T7fh3YCfdWhONrWGuCog1c0cR1Up18ih4ue1C6L
HTn3vTl7pjqNzXAQiS+Ixg9QNtjk5+KFKSMGgaXXBelFF/SwwiZqCwE4DwB2
mI1CjuObCq8bHj7V08UawCY5ZX4cXpBUddAI8VBxSAJYvLwT4LZ861RPI5Gs
tJ6JHkkvPgz1ITpEV1D+LbqQk/vhT82oNfnjxTJeCXSj6ass4qLieAHWPTqj
XsNeZQU7sjUCpvWFjAplxvzpPFzT/pCbkspIjTNl7LNTxCA0NrEbv+VS8lCP
Z567mEIlXf5nsOGLsr8chzTwcF+pgCVRmv0eJEUIfClppiae7ULqQcWb/IUz
HpGE7jRCHMGrXfyPNMTHTGCYrnTLApHuxM4aDktv5XSoarDesIXcRjVnT28b
7BEFsf/e8Ptj8+i4JG8TUKjiMun/fSuk2+aWKZCeQh/+PnhWbIWL0qLXhj1z
Xx0p4N6t6BbnwKlW9N/wmTFU1mJIIUfcCpKVcwcrBYPAeZZ2PxZXSR4DCHS1
2K6mtdvFOIxTZgS5Q/edeSa0vwcUAwc4uIi5WquX8EZG/+z+H3o4pWvK5NG1
Ufvcj2aVV9uZ4h2s5RdiHWVm9DTaouSt0+J6Z8EDo7DOuAj3+E74wQKWThcu
BozwHrdEzZgiI2mM6sAA6KQDMyH3v+/aWvS9z4nZ8tLTIxIiRftqa1bx2nOT
tUq/5Kp9K89ZFGhYkjjM0C0fOYOhtRaGI69o9dI23JFHjDfKxjEwZYEG0/jP
dOUuas19KnQWOaMhYbFePPg/hcO3mILzgbfYdfDA20iGdwk7xsVX+mWQHhtE
BB7l3gQuHbD64/fPCnsxcdaqHePvHlGB9P2rA0zzFD7IH4C1NQSdbD9RWK0d
Er0GcPC4jQBqTYtanLc8Tvc28n6RBvFAaQNrQHPNAfJ++D36jFbc7KQV0YBj
BRGA9HKP015Yo1OiqBA03Exwk5q6QphYAIWTwBDamfSbIfn1XotQbEVzSUCX
B3P7h3QTN/adJ7CweiWBfi79D7vuflyBeQo+9f9vD3KjFAjLjJJm6T4ttREt
WkEBlKgVlfEPOBsT53t72a2XDo5EUdJiE/S2Zesi1PF+AxTDMGMmWJ/V3kIs
01qI00a+1tC35ApN8K+9au5gMpJhb1Dbxkz0obYrJaU3oje0Y4eAzi2Kj3BN
HbV9KM393gk9MfV96HWabAJjHA+mkG0JubW+oCSMN7RPzUswiCkT9Fg9NZ4q
/0+iPj22TOyQ950GnmDx2GAHVTFm2HX7JwduG7VdvzaHGqJgJggoRkNdyeVZ
oSlQsEwe0o5flzuHfhVskOdhSWNOi7qeDUnujIMNaygMOylUBQU2QFI7uwhM
ova+nQZB63BBhHAOzIcQvAaLfYKhV9BC14IDUlNfvRiFTh36eZpHU6PFbqi2
8S+k3gKW2sd2wyx6zgJH+wjPQZtej8L3d6bVF1hjHMqrBiJaFyNrmsoA4Qy9
gGr7V2PQL8yABji8ayo6thFN7SCoNwOUpjbvRWz3GPVSHNJQvykg6OYbFkkw
3CsMuR4KfFuENXFbScx+L8HUB3mz9uUChFYm93zek25Rmf6OL5Ut+8+egbBv
RogAbxjShYh2pcrnDOOmMG9LWZ5iVpFRN/YJpg/LfvKMkA+Ycr3YAu5BbjAg
4cl7mxnKzsTNp79wWiBcAm26aePuHjAFksYovg02srXPQqT2ZSIiwNg+KEOi
z8QDSBj1TNUz7+5TLnC+3bdlpqHjYq0TMEFumK1p1L7C55kUh7Vd0AhzoWuy
nuKAp+M7hEsCpxTE2PJpLevmSDu1msRwZRZCtlM9++m32D1norNU2QDWSZ5u
kHoyKvNIznp7ytMZe2JS3wusVuGHRFLpozbJYlW+eDJhgeeY89WbcDq8xdL7
9ecJf9Sl2sbR0DAna2ESTO8GB7LVYm4g/fSBddhSPENLwzKzwxJ41DXx3F1G
4OjQhVRSwWZ1F2ssykq85YNDcxIUjb2R+/laezsD9/j6/AE+dIFsaHR1AqcW
LIXpjsmnnGnZMofoOlSg7+hFTBdL2JvWlJdh7LiDyNWMNDvot3p1rbHaP40+
knXggcfWuvDstvnf0s7I+D1Y9u9z2WBOgxXMcB70gZPkSrPrvY0HO02uaTtr
D1uSmxaToREgzC0+KVx8DY/+g06bWt5LPljnaI91Z/DAd7gvzK+HdlRZUJ2U
o/QWr7Jr48Js7uE2AdFHzjZ7HDLepBljvcTH/ZtTz76+ZKLA5uyBLVwTGdE3
Rt0SCEXVyIqbwlsnQ4dda6bheaD0mF7f2JH/wO7emZL65xgxRXn73KvY6yRM
pjnjYSqOyd7oVucnx7duXibj9YlPwA4AKZuLISofLGV+fnpu7y0EfVqUo2Q8
ohgkLz2L9u5xiRpe0PTn6fMn+RQD3mP8MydELekUoUOnlUm9oUMYiv+yzwfU
sGOEBtNUEqR5wplydikDtNP0vpJIXDjXQREOY7QLakNiiM4wSmIVntOpVgsl
XKEevL/IfI7F6YT9dA8mPKuAXvh8q3F4Fc9onFyOlRFX0a5RofwCE1XmI6lp
N4xK6+3wXTfNE15563vpmFmG63J8oiurEdBkAlnmX7c36stZdgtA5c0YrVs8
gL/vLg6Rkch1n9ACI8WzQEkdof/5Qdh4FC9o6liUCIpJTBx3wZgOL7acgXoQ
hC13eWDb1hb/U3StkD27fsGwfn1t+4dTfKWcolik5SPWpYG9wuOYcwokVq7m
MRF8kCFBWFQIGNCMWhaNfmxrSOoEbcFFvShRcEWldluDIHx2Meb/F0yBj7NL
5Qy+RFsKQN6wildXTJRGqMDVj39IY0+Ykm1mFwuGLyEy1GkFffCbxhl6Xs0I
D64zpJhgvzhHYmY+Ev6SZpZxX4TOsf8M4WebSpZ32WqNmo5ktSEUTQg+sW7Q
iBlP7GcCC0gugZ1urrmEPyDjjkIQMpjQxdS0CsbygpkkFnZ5IkJlE1ipxs2x
jt+s8tPxhOX2/IBmKMugcSJCBCDKN93QKadHO53VZymZov9JLJBQXVDcRzVl
7VJY+bca6joTpslEAle2w+8zDQGcM0rng9zeRZ1jBMX4N9cZ52PVCJQow75r
saDb9XROTrlWTseRz/sjBANA8s9byzqAaaIf5M7aTMnBsyArLZ6VF4BVLVZ1
F7i4shLUkf3FacLdLfWlCQouXXgjyJr5/atfGxGh27ZmYKfK9BKExM6HZWMO
5x0AvP3AHsVQxd37OdReHsKBKsE8AgN2MTEztKe0qq59K04oYFqSiNT/Nrlp
KUJ8WMJSeUE4b1APkl64sUhz2veDehxo9CJ5pe2cmZ8Yo96AlHapvhfSVIAK
ms/jyYltYMzA4/7FthLLM0LHPKHyvWkAwFXpFZ1W126CH/lsa1ci2J2SdAkO
m5wPc5CBQw2yIJN0RO8YMmmy6DrHKXVdTeL63SBy/dMoXcFe2J9ZsZvQiZb8
x7nT0dgNjupi0dwFe3etGZOuOjlgUB5PcjneMzkgbSZJFucvOp/ZHJiNjMcr
uaY++XV3CwvXwA/boFowqcKrF5XD3cAjFK4sDdMgZ+vai6iwdJXC9JTNyFdS
OeCpxc1YldjNlwCtgfdmDXwo1BAat9Qdxp/LN1/JDBEsxjr4RRUcQz1iqKxS
XUd8dr2opKe9ON/yKWQ+mu61+dEE+FfU/ZCXx+bEesNSQhplWFg5PYFAGP4d
DeNXSJL+FnnHz9nbdHrI6YAeoDbWyIGVBNs5SgFNkFDN3n18nm25AV7Uei2f
s6ksFUqJ3dM4j5/FqI4CN9+pQqGjKi02HAv3UdjrzKgQE5FuU3QGsw6Bu6dY
s1vgTAp0j36JvGR6R1TVk7f1MBFg+TVd2M/RYXkzuWygNwyNk3UpkOnFiYvJ
cWDJK+jNeRvO3c9lzlXEX6rxVm5EDrDNiP2yz8wuER/XFkGMP8PAAZRt/NGu
G3Fwfuu/msNHlElieAOpxI5Lw/vbI8eI+Gpy6Vb1hC4WQQtIjlerltNV5gXa
LlMOvtvvdNMQt+Ddt60B3PlqFK4xBlyYP44oez6OfBWJJQLADB9vJmtOgieb
BSd6IbO1n3gs9tMOFK8Y0hqm9cEub6lPfIWqgTChKaz5qwK4jvP3PkXM9/bd
tRMRwTGKM3FI4tQa8DFnEXKbcqTVHNetQsvWtmwW/p3tqYR2D0JeSBC6PdVd
PTjwqPwu6UuWbIr1mLzkCp4tddR0Qke57fAevwaiz0TsXdtZenCx24GKE/KG
1Q8w//s3r/i/jT9dDyNNvJrE3DqGhxNWTpUMvTJxGjeAXah/98xxr948Ok8N
2VhUP+QB2tl7m6PDnEDIFp0e/slLKBYXygXUf5XJEuhn6wWQq+xwj8WKCNbA
52pOxU3sdpHCG45U7C7h5UtEIKSJaqR6+V2GOfaftKXG59H2YXW3z2oI+KLK
QEVe0Eck9EWZ1D+NGTEzJp2WJOSTfOaYo1fN8aS4FBeVm5QACHUiNdExFeHn
LqeVnY9kfMK0PvIcqjbDyTpRk+A8ebelHilyMrW2Ka8Ne8Our1ish2mvkRqj
zu7CBkWDNR8yNOOPlNPkfT2rug7k0lrOu4+hAQHkPutlJzAy4vlM+3ccpj8p
BTEcDFnCEymYwdsTet5MTfkNa7kJWEKXQp4t3886ojctx6UCuqa2M/P/VzxY
kfsLGC6+9xDY0L3iYJwaiNxKUZ9/no4r+3xzObclXq2V+8+XcTQKvqYWwM08
io7VlS+UqW06WqF1BHyYeVr2O3hRPAllhyhdQDtM0skvvbeSxKyV7BQRKM/M
zc116FKTb5UQDmMayeYN11v0Fw+vj0MuWqKQqZuoBA2xYkjb+tLfkYd2XTUd
lzvFLY8f8GRbHkZimpOuS61MdWnMoroOzc6DjAgFnFgsZVEnRMI9xeaMXFZy
WZTwPoX3REFuVzUrUi6rGF/tnDTGCpMX80eAtWvb55kjuP2dtvMXO7oVDOOL
IoaAePo/gXEUK2ZtQ0xGIyYkhNvHqHFGHLdYLBbdQG28bT/fYJsrCVHF1cbA
9zooAMmNxAmB5OapjD4XYnUVm80l4Vx5UJ2LUGagQw0almE4jANtmlU1DKn1
YY8Fvxy9abQouiW0Q+oRqzt4zruqz+mkOPnaY/CoDwtI/+uHl8EzpbwndCKQ
ZGmazwhehDFdMTKTaFK2ZELAC0hhNxijm7siH2UEsesGiPaLCPX8BuzShFVv
0cExSHsMOxl3EQ8ZFeH6uLM1/iMrrmeg6la+v11HA3zgahdwE81apfu3NeHE
8JJ7H8ShX7Zz9y8KNzBjwChzWXz7ZLdmWPSorlfiV0qTzP77Owq1/Q5MzLRO
YQTBjakrCb4yzUHmk207izh3TzmN+eAhjzl5Lidsm244f3iBBmlENeUZiV3J
meQRP5LGNhrP1XJc9NMFoOh1INha12sx8HQTNOMdTCZAqde/PVRAC0Pgzz1o
a6dLOu7EYCC6ZLqnD25Hr7T9OJ7pyrnJnmM0XZANSoIxHdqB06v6IjO3ciak
0wLu381sjFH9aZYtIjQrPkobHdyh3/UTTLZsO+Qsy4skFwTl4Mo215u9UHYz
FC0koiHdzvs15ixayxIFfrZ/SiuvI7fTuorGjzh1M9nq0sWEfe7Qk+0s02xz
e4s+KKGjODAA1nuzQLL28MGDTW7g62S0N2xYanUjZeXuxWTkVD2NeFFogHYa
EWy1G3QkMfHja8Zh8PVdZzV3HKua9w9kHu/maRru8oJ0FDQLcfD+BuoeHZxT
wo4ncCQF+amZO4wBq8M8b6dOVraJvdCuLiK7nkNPTCLJ326aubCN2k7i27bn
xNFZtve8cAuK4qAA8tTCXtPcMSFtHy2BdSVbJmoCMY+fV6G4f+LwTbACjzZh
kz2jZp6Xfe12vMtOOB9mJgdhGizbcW1i2Yp8eXX4NV5Si3QEq4O5zIlKP6hr
UgbjPIXhpyhe0/TTHptXkTZjUTdbSg5f2HLz0RJekstAudlDtc5SWbrwc11b
wxLH7nzw1DZsArTjX3A26ozCPWmaQfBy7e312mE+EzXLqGiVvNWgOGanJk25
BWRwe+8dGx2pa507pL/QxXx30nyjspGCpQ9/LixsLblB74S2cjvKIHt1xNVN
pV2odM+SfStIYRF4AALruyeXnC8fyOVN7YQM5oYyd+SEhmYcqgQpk30VqAY5
JpbXgXv0F695T0cuBP2TDdNSY0RmK43kPeYaZs5BaaYyWFPDIyBq6gU+e4Kt
1agAxg1WLca+PIAzqhjjnjqEKHRk4c+gk943wd8YcAVeZFpiVFzRJi+KASBB
gFkUIpB/CNgxWqrgAk4paZYVc9wWsl6gOIjNGTKp9CU66SOcUsNpc5i7nzAD
27WqTYzLYHiGqO2OpVz18RoSRp8GI/+c195z18pLMQDdGcwJL9H5F4lOdCEJ
Jt5lNG8isv/KPaK37MvYJRnkwr5hcJRtgSCPK1YMbVek3Fp2x2wsb3W2z+4m
6LKscFSNd6V+ie4GB4b8hTXIL6Ws3GmduOy5lnqe7QPjRPozj7x4KN0qWV1Q
GY/nqJQmC+fJKm6S8ndPc2P5WLEYZnxSHwB8JRY9WE+J2PDu2Pcj51TxeJ1n
wjQjTuTIu5BpiSXwbpAOYU3m3Y0DrWbL0b0TyWZyCNyJU5/VQ3Kycc69QDqJ
E4km4XM/RnXBAmDHT51crPxoFngZdO2ctuXny/8+4mO7uPuNWxvY/urTvK8p
ylRu9Pe4GcjSg8/+mfRLfUwUBlXxNoDvQWZSQxKBmhrIoDbleNo0HPO9chi7
rt+U1jrYjruwIYuE5+i3WWZ6H9QpgKtAwNTTifKRZsDKUWaaS6hSrFq5QwvX
vQQcQurcIhRJyiHwR6CkEenMCUkKHqtWlc1mtoBrH3e2f8PGq4C1Gbwgvc5H
2FqY/Nyg2J9s8RgKr9VZTuNyKeF2aszAFHlA1GzI9D4D5/WWtELLsIdBKVqF
oTVPuIvVFznY/jxyMWq8lJ9JemQxl4fLcgZvzXzmdkrrmiJs/n4fmkibqomz
XUWEPQSm5KS9RGo9zi2jHAcEqtIbWMOcG6VPOQckUYbVOgsy0WRWsGf+1MUr
E0+IVDD+Goipk+zF+nXAJ4ka2pPOFkefcKjED0p27FYPcyPhFQoiBerE1gLL
l2ur/a3HbPIwP0pd6DX8iRbjUw0rqW5d8ejA444qVzcCHzHcAmdEgHRfl16h
Vhsn4ZCMd69dDP5PovhTTW/7UseXCdWJECPgUMWvj4XZT9nrOB8GpPnGura6
4MT0PBmX+ih4/tUaSX1fr4D4Il8ni3kV5YEMfxJdXHwVvKywu71lyjtadhso
4vrcSbfKezjTCuav0riNiiYTKi3P3fTW3TboOzLWx2glpVfpCtRm9crJc0dP
UDkITIU7QHXDLtaDuvKfohELFDqdokI39q/9xbAX6EEqw/8J0CYsSNkEs09g
//Y7DX1H4LIWFM9GWhxHZ5BwqvjuuJLV/hW/ZLxgPosRoMVv41+mMbDGMLcN
yJAMN23NXrdeMy72oRJNZZ7FdozD6aHzPcfJJKPQHupUjvPhVJNix4lBVWbE
ROFPiQgljGITIL6/Ppi2dmJ1vz4zSy0RCNcaU9Qxrd2cp0mPnzrv13FAiAM4
LWjeGOc211ykjRHA0RppB+2PUMuN3Au+F/SB1p84qP1a5GKuNmnuCUdmPn0j
VfgC2+Yhs3gBqfVuDuOqS61Xzya6b0twqOLlZTaVjbVt6jYp5cknaXJA7DWG
9w3Wr9StDuKdOP6IZLLJ5w5DuFLzDpmdo1QGLBQtcHuN83E0Ld6fWRHdXvST
W6dgIabOfmvj2fHGORf/v8Jl6JwuCTqF4jDhaXmsEelL7i+BQRis/gZwcbPj
gU5XylcmRmjmZdoufZlzc6PmSnqb6L1otdKhDCtcKfXpn6BrEssTQBFQvEeb
BETxglHCsMEieXsZ7t6FdQZAkXWydl8Y/6QfNRzrj//W8BqarBKgjGkLnVEI
poDt0fzGTjwCty+0uGxHYp7ZwOZ1G9xbL39+3CqfjbDaiwOmQEWgTlYb9xz+
bWgkpA+diOT851T7qEclmk8k/7oPtUw9HNawoDbfMVT4EGTEi4d/p5Htkm+X
DEv9pJBeJymbwX2uUIcM+xwUcsWzqPQ1b56Z946DGhyUbu5h6uhqNzGJYOng
f3E8RPnwgI5NDGq7gOnekKds1+qfUqmw9B1e083nCBWfTE8RdujPXOouDMB+
pxpBSc1ictzDFlMwV1xVCb/jVlMOHJuatLGO0rVmWVZ0+sIeD2EcVmpA1QAm
UyWG6r3kWWCwHWyHNf23VZQE4lO+OnwO15TzSn9kjhc9yw4ugpw84U/OOM9f
q5BkR8NzabkZ065PacMJLiZrkdbKZNPglmhyC5kMLB2mnHXllAGQUnrDeYxE
ErPc3gnipFNBqOK2wdxecERPDqtLHIbzsCzKT3Kj74CConjEwyuFullnwe6f
f/GVd4jyV1cumyYlw00/PdOvZVtptCzq4F+xDNEQUAE2uby5aoFD74gPVukV
vnZzMu7lp5wNQ84stCXcaOTHMbMFQ2GRTG3ZZrTIZ4gE5pcVnOckeRN7A1c1
NaeFtb8QKZSvqM27yVm23LY+5qTX1LMFWcB1aKwy3Lu6KT7/ipfPdnZB8zCm
Q4hnyVhquKw97+dzbPsy4du65aAk1PWq4ypCOCJ9tfCQUPfMlHXdEcaHB2xh
rEDx5cTIbgSK9oJOtj5T6dl7SHgvfxpHanqLVxgorQqRSiQ0E7tZzEjAXnl3
qDMRv3wUu/E9fvGhoLD/TDFPKZMex2NMMMxg/YuONOferDSL5+UsQbJB3lM4
ngkZ6BMqDw7dZB+wsEm6YBgSnBcbkYE2IUhRlybaagghKLNmBTURPvExdgxC
WQcu6sV0Sgj6jRV+d8ocmZopn0hjvsBnyUhU/YGlW9c+MEXfq+/LvvErqB7z
nKt3DuPLwZnipc8q1zmj0G/y4wDdPsNVtT6b5vhtTUN7T2iZODHZ1bwtxT8F
KJbAInGefQ0+QYcGeJxPVvE7FXO5zlVU6nxA+y1upIXaOxny0FeMxxipY5ak
swtWzfPwRxPH5km4LjLoS1zrtOIqAq5xQChs631I7kswio1HhdG/4N0uyQg6
ZPSaTCnzVFoHtzR9EysHrK1KlRc3wt9WsbbQrwpPK9a81u/8GqEKsV4w2CZ+
TVqntUk1eUE04YlvdwDIAAmlBgHBiR2HmBmTi/EEgoGOW9Z+eEdQrIkLXQt9
m7Va4jw0/JjKuY3XUsFe58zbIyTGtm3am5jnkZLoFER/WV3OBW3ajmBQ1NQ5
nnyzLhUkteqnFIxs56kDb8sbg5rNWpG+pSC7Yfenac6bT3+roHe23tmrMwcS
AbRy4fDnzHUkhP0tkE5cfwa+dvokx5+iWqQy87BA+gHYDKPm/Qr2WYkVOgWk
SMx0XLea6CfmW0jnlLHwGrjMFJsEOccb5yNiguRe0JOlDvjkM/zr2fK0vwEC
hy1m0Io9+yOdH1XbaJSj4K2pJWX4Y5GrzFaTZpASJW2zpNyEgwlKrX++bGDe
yazxDp1Hg4DjQwB04EwZORki8o8TsGbdyk9DBJqlG9oJVmmo/wdOXGHohLo6
t8ZGYBtfQimxDPM8f0BSznd7HY1vJGNJR0lFxWCFvcST13GuMSPfkzrzWKyX
88PMalZHGrqQJ9AKBrquZ4jmWUU893ldK60a761dKewhtCCMZBZwYKjz1ejH
h+ByaeDZGIeM1gynOV7G516SJm6gfB5+3Knt4WwT4TOqGCuK+25kSE+vgddb
EVQyYPTJBiHmRFVpO1H2IyxMd2TaMYgOuW2IO2lu54z20nyevFx3/g3qegsu
6cRSoGlsMtddZG9xnYZb8AyR01xGNmEJhL2XXndjlur1ToFdpxlBuGcgvZ4z
m3n2JCaak+Bv6OBy//xpRwvKQp2VnjC4ZHquO3IPqQj6VTGsQ2xGdQOQji5A
3N0RgrssTQga+V4WlEhY/MN8zprt6e3myMaAOV0WMDnVtpWTyacqK74DGEC6
fPpfCKPBgy6mnOTTwqqfOB4woADgheo90K7wwLihG4qA0NO70mUDFqESNi2L
uAVYsqD5i7secSdV5b/0+pXQWfNiA5MRn1iNv5+6PqgCdMfMvZyppSL3a1SP
nQ5qlMEaRJBwJDf9NDKtJ06/aiXS+kt+WEXjb8qykMudGQKVNsQgiVQrosuH
D3gySZIHoYjtc77jyEc18TJWzTi72tGndYBAiHQNlado8VlpqHPYSxuX6at8
KaPQE6ipLtClz9QPqLXU1B8ULADkXuJlCDHW7+CaKJA1pjGnZL0BFkEkHgIP
bjkIHtxPaUb/xV+9nM1jxCsjLr6TIpc0h/miBVDJ+fLrKz22TA/CCa4fijyH
pJKQdonHKRPLVygTnecjKNcmLKVhccLz8e2XZLbO57BqvXvReQztECF86o/U
Cl88YVybiI1hsCp5UGPfgLtN30buLGxHm50K9YvcRdKl9MZ9B5o/i8M2liPE
wSoKPohYW2ihsbjV8ej0QnftVdKynxEDcnTiM6tAHK3gWGycIjewlhfYn83T
vxF4XEwNufkor2Lvxy7mAvS6T/0NK6OjOyd9l3DVU2mEifCCQNYDKTLxt7bs
wFmcc69/b055T7JGxbHWULh0nWQ3oyChlvaBMcBNAckI6laq+G7DTHIGNNil
X5zbbrEeR8xHbaxbWeW/Fe6IkhYZgcHSdrHsEu21JQT2NQlDyrRpt0yYz4uj
S5DRrBFrkhAlOvRl2lL6uvCeik70n8aljLz4JJAS4KdQ1xl/6KDK4uI7sOHk
h460CZQcc6Ksxas5frZOI2l0J3BikppO1RM2fblwnx+zEcdtrdPFAyMZL1Ho
AXr8OTgBQ4WrwaztbMti97ChdF7EYce9s+5SG/DdnKwjAzNP2uM10LfaAmz5
rHzIV1uMg4cELMTxS/DnFLMfiR6tro974ypzDNTMj2UuCeYPxrKhsofBL8Sg
vW+GMiFJD3p+SsfI1rEDQ6e9wLBXGmQlvEiG44cF5hgDQyE3uFnYgeiv5wo+
c7AUKSBo+cg6+z1XDYN19rrwMndAn7znQStSDaqxbJI429kaA0jpYD+IutC2
vlxwSYFLdHGqYS7cIhdB51L7NmkRdE+fC80gsrSkqJlQdZm/0HhCt1Mi//26
aTtfI+La4WnW5Iflf2BLsB2luapaO6k4Si7A+y/on54uffO/lGcgu30A2JJE
Ihd1sv1POvu1vwFj4YTiFV0HBTrzI7d2WEmsGYXUYGo3dy+LsviMaL4pPHlP
XiTjeYqhCzeFnA/THWAoGbecG+tbMNEnAHVq7Rp6CEmXoCD44vb506THRi8o
/KtGZGZOuDIjOyx/Hh/WwG5FiZBHiTfKOQKyx0FmMNdI2I7UCmnoSPQqa03w
jUDHZm2xApl2Fqh2kLZMivKEWfb1dq3tattU7ELPfYJG8I1TdW3vb5M3kYF9
/uoC+hbIzsydyvbV2I6G0npzfcHllUc7fbNmeyefpckg2woU0RsBRhiOZ1/w
4GVcjHPrgngTA7To0cQHHqd7kbCloemqhwvYv+LHAsUfjazrtaTNz53Ex019
bzogtKAgQcMqh9Y+lMwXVDZ6FwS9RM7fwGu0aDqAbJQDdB/pUOY50c0YUAJj
au+iBxPuE8d1pwhKpFSj2wQe7Y6pKFKxbu5/a6YtNcutnj8X+wceoi4Cvis9
5gw0DyXn1rgL8+YKRCcQRgvr6NQzhpc61RepJRdQJC0H30vcd6gBDaJxGp3j
i0mUE1LRKntO4+FjuFab9ZPJSPMdhTcDVMhEw1neDgt7KV+9OUrTCS1ew45i
DAflx6cuvEr2c6nWlPdqpJJ9Tgq/nef375Ur8COM7LwVV0OxvYPooNhned6U
nfFY6zrV1zpcREVi7H5hAe5SOBqKsy/G5dvMImtEtM3ud/2GR95yhwbfJlH+
2vBU0f/Z1ovdRiN2/qrWm1vkz888v1q1flUOVZ3fuEYebhnyJ8Cyy24rEXLa
JSUJKB7p3apYRbwPnx1RN5V9iBIQd4F9TP0/Iad7XJ9BBODNhiN1kDgcYKgW
4ee6L400LdcHH6hOjzvSQDim9OUfRObUtBpZZdjM+cKqbLJPOfSFFtMBJPax
kNJkY+PGGdSgg/4gJc893/uWf45lCPbeGjsObuS5kPEy8EcmAegwthvJV5EK
d8yb3pbc1dVd29DeZ4aRVcVettgj/xGOTz+yeJ+2QjJWkz5RdH2l8PDpygbo
dJPnwIxhamwj52RIFKHbL1J9tWtRcgoOOuJXFEHximpK81lWY33gvLG/npU5
WKNR2+Ba2g/tU/INrKQzStme7DKx35vsVS3fOMddubCPiJjHxbOtPC64P4BN
plplfTD4+IKU8KGXULMAtv5AHkSkgPCKiY6L4c7rPRA5cevaY877BOYbJu4k
f1MCbsp5wLEoFXGtIZhZExlnHYNJW/7NY+3nO9a3VZlVDkkMVtJluOcwIAJD
n1IPnbhzru3V8rbjG0odqFObr/xtH1xHs7hlatPrPmTXZzkO0KFO50XBEMEr
y8p43QxWZqnPm7OKQUwHTRZYnFJVEaJdV3sKlFSSHWUfM43mmOdP8sITPglB
7MP5d3gm25PkBkzbh96sBghHcxAkQRCLO1wB8aZi1sOov122x6pHhzwb9ZXL
cPj8BLuz71xS6u99KOxCz4H6ESuNK2DkBWhqlzmMFkfrMggyh0LVpucpkfZi
c/wJE/onwYmUw8UQ9w9oN2D9qIqQZUVCfZCCsHCCw/PSS9cIqXbKC741+TtN
holHvMmyGjIXxsD9haVWdiYkindUDx013WkYC4tnFRLP9VqS+hcHtACDIFQ8
MGisRFcYs7rcYJDBbSsSGdr38rgoCIcn35QNSU+R3GGB2cT9Ly0leGh1eryF
2NDnSRyzXTeP6OHkoJy3GIo/MTJ0JD915Vx8BdaJRLUgq7kLRnCpfBH0kUs3
0YpEWuKY/lL+eilXtLs3NLtPzJGWBeK3EGemgCO8Fl9Arkkaw5iKmHfXNY7F
eCEAZZvyRQw9sEbUsqpfCK4JW/cQxpzW+qHveyT5Ify9jETXYugkRvUgzI3R
MDVgAuHtRbPetsB7cnQ3nfofe5SyU+45NoM7aHbrTitDB/wHq+4e3eej8FRb
7QdkfnNJ8A2nvVA7XYd8vaJVFq7UmFVttke7sixgqdUgNscOOnA8C9pGxcAS
ItySMZdwHEPMH4g95GhJYM89s2I7jQi+VyKRiSAsMzX3AuPprpqwEQuu5i+s
JlaQpFDJ91oS+xXgm/cewLWJPIDxn6zevO9SDbltrfYXfuIvyZ4rK7+C9xWW
FHGjhu8N8b9YzNLqR/sbKhp3Pmwz1GEJlBCrEIbzF5P5dif47DuXZxUB+ZOh
iNYygcanqPkQdBl1WRFzhHWe0oYGoTyw/Q3W+JsHXxBk8DPA2XpHwNW/WWh8
BUvwopOhJ9Pp8JsROZzaem6VPMZHFRrc+d7NI8ac/fGcgqQVVHijaIpcSRqB
oyONuPdeH0mHmPbFdh41ylMoXx4YTEc6TjzfUt/IW0OUdrydN/PGdKNq32+t
0H3yFxfCeiBVx613ldd54rfbqZ2aG+fANa1PAOa8QU5Da50JDILT25qEd/+G
VQkHnPCPFhrMx5pQhGyQ3JRnt4HCxpDTEYuj5KWy73PLFG1bNJdlkxvHDzXM
tlFm47bsMOSBO/LMguibZ+/bWCPsJdIePHwRc8Qme9ks0+yu9MB3zoqVZo26
RTzsYWANNGK4zwLH/whSIyiIr7wZg2uYx/AWmeMm3spKPuW753GwIajDv4zg
x2EJfDLFkJ0TYOdrL0iNVYCGtAxDGqiUsnTHg77ybe4YUrmQbYMyJhBYH45v
JaDydoOA3R10bLlMrYjD0/uTFsaV3cgwya243OEVppE1+JqEot35zHJaA1WM
u+v+GrUqCblv50AO3DaSq7k/ghR/S2dASuCi2G9A1AwWU//oLD6qD5FLJgqx
bp+IHDlg7l3vXAsXVZf7a8pMz76AJzdkLe2+T916MMoirxXbDWSWV6g120fn
Ikg0KYPHY/FCSibPVW/W/4LtrXsf+xNGkVyQXDe0wJYRKlrMDr0nhJ9/z3ho
jNpxBltTB3mvj7OLA4vzMk6vqH8U3t93DNsQwyiFGSDLTFNdzc6yQqwlTQTg
d3v46sUDGNinBaXBOGpwtC1UrCm9o02wtY0cI3xyUwKSzXDafRYuiU+0vjgt
dDZPkgUbarzZcHpOmSFDo7FB+ntRen0oYw4wqtgD2+RpMw5rGdiPrV2jnKcH
npp4xnD+7VmNzwtQHjeU3+QDNCgRBCb6Rmh3DKOcbgOTR4YTrpSwc7acfkKY
gF83MPEBK6emopcAAtvyY4xRtVt39aciL1aptAX+SOAacoEDOUqC7NDm0a7B
moPbu9YS8mxMa3TrFwzJKBnOX6i4GthPFX7CLAeYSmfP96GsQk73NRYtwOG1
XPedY1cZkGMPEZD0dNurfBVP5C3JPFbSaQL3QnN36iy+L7GoQLvcdP/F+OFH
QrBKpKTcaAkfM0ywwEbHJsjRX90i9s4r5lhp1j2cNflM5Z1b2+14q26FI3kZ
Gy1peMrs1uNA0U+53+fG4URg2s/FwsNceZlnrDbCJ0NFxPqajw+7cY/G2w0a
FXXCjxhsuSeb01nWiCXKdyMiCpGoDf6rA7YnBJIvxtdMVR9xfCHCEHOnk281
/Yn923sKH0VDql3eWmMCFkzLKAdDMQfyYxYA06Ln81oFTqkgyzuFrB/K3odH
MdyxtJ1IQw03iWuV4TsxmSNVGx55H9LvZPcg+KMWfkCI3QU+TvUnRgzpkC1I
9hhKu09tzBVmezBBRLcpUGS+vpn/3umLUKQMVM7pt+PgRQpMUEsFc8crOBN8
QXw4olF7LHftDnGSYsZnCoOj2d9SMpL/5NiLBpLEhA6RlKqG4YSXEuzbxCnE
yoRNbyCmLssgJTK5f+LNbLYyw3uHqBXeK5Q7HXy1ruF5xOEzjnfMLg/YpUh7
jzsAApLo+V54UpSGQApoAvtQqEBfxBB1tHvZ1p7chOVhDIltgzpT9oyi0PO1
xORx3q9705s+TuROvq0H09oPw/belpNGGl1EJs1FzS8hGWqARvoJGkIbdnbh
Ph1rFRychHAxqUIX8bg7WGY7C1pkhSk6nfOoGphwlpbbuoPOmjykW0DrR4sa
0IaJyy33T8qdC38YvE91TwYUfVCQi/qq2WxKDXDBVfqL/KMM3hReY6NEkM/w
HVK4rcnu6VqL1avghIBbGYVZlG4LqjuMc4CsWlIWgXBwcCGkJ5eUsUhzOM5q
GfTAaBqz9K1KCp1dX6slxMOIAjvwbB9Xi9eR0jcIQ+VhnXK3v150Em4K/3QY
54Cw9t2PJnjjusn7hA4ASDZhu/9/p0SoAg4QNcGgPqcxkkrpGJfFBO3JRcnO
z78MVmEdpIAkb0PLsSxhDZp84VqS77yRDUge1GgobMOI8oDDjVP+fqYtGJ0d
cKkvpmO8s/O1eEWuVtQJdj5wIQJdzdaW/xeZr8QmhRCa6OQtUyWoGKe/0m/W
4VmPkkxsI1tHTu012RwE+cpmCCKZIroO1Ms+2HBTWVQjD0P9eECLemoGpCSJ
j3TImpyvEM1hBCvRDOHl3IIOj6He1Eu77XYQ4GeOOIbJvbsg36gk2D/AyEeh
N+q6qENF/KNj1pSKYfbQbzfcpqSiJOYP9B//CCLUmTKI4VB39yqnTcKvEuBX
Mtun6Ec8uXBhzBmtlbS9+mALeMUAu627Ik0l/AH//zwuWAWeey2C9TIoz4x3
uQpIFs5aZALW2au5XI7zcOHa6UmR+T8izuQjpRmQmvoKWZoLydEFBAHKPxoo
nSCP/Oq2FWJ2gKtOkzz61V3APk/m/CfkP4F4Ln15xBwLH8S83+r4/2l3mQad
ahuxyxhHFYfn2R6S72DV5R2Vv26kmveMliS4AF5Rhi1IBYGw+tE6wpSGssxu
onfmg9KH4wDZArPFhfHgsfhSdMYuG0wyW2Udo7EYZvK6xIwLqvJpyRIQNKeK
487KICSJm1MRQcA4MR1Hh3zWj3jaZd539vLuvdI4exIJc/Y61ZxmjTcOwEsu
Wgj4bY3YdeHP5L7HEiWUFXKXT/X4KYwSQusFPbRPsCwiLYW0pLu5psb0xc7r
kWJt9XC4oWbKruE3tHPUoHggoO/sCRS4x924OL/AibqHQjiDe2XKl7W0sCMU
GhHZeOW9aB86Wd+voAmKcOJki8vhcEGMgrCH2TTjQ1rwwzkE80y2CHiM8Snm
q35kw1//rXsHs2eq1lK11/Yq+j4ib+LEQ8/43Fv7SpRTw8b4e4i484FrhRj2
O5E90kdxS3CG7at9PfJVIbu003ciylH1yNl7iCY0mqkdRiBqqExQGDCEEzAw
mHglUPD/G5LTS8CD2MfIQIGvZCCQmE3U5kgUJ6+69Og09m8NK1S2aLY5Qv5y
0f7/6DaPO922yfLsa12jWSMAu/9ekXLiXMME2Iotuk9akLIpzdA2KXRpNILk
9oY7aAhWsc0dy1JaEl/sW635Jdp9QHc100e+BgOiYclZnZw7TqR6LVcvDcMx
kWM6bimzEiLneTGqquMsRO/j76Aj5Ri1c8WFpUehuNlj2q7VUQ3u1VuFa4OZ
E6u/J6XS5piuRcdy8oYuL0YkPdFSrEfstemOTstM7KXHNLKvF2yk74zoCoyh
7cERbj+MCkzrnGGT4C9QNfOyNgsUTBdUsc7PQWnRKnVPzONcxMrKU7NK2yCT
MB9iVgXLuRB0v5YcdmRXgrNq3J8IeR+e40SBXVL3j5WOhsmtsxQnv9zcs9MJ
hHH681RoshMgVF6fnjjPrTkhS1bjedug7vz8UtpTMhHurviSukamISLO0ZVE
loiYwFSV9o7MlZDebIq2MlhebC51Y4ikUAdFZwKXYmhBVhyDjh+/J7N4gVSa
6wOQV4rXHaj7SATRultOCQ06ReWR6sRUet96PZmymAmeIaC4D4nPpyIRhsZg
qvB/cxRluKlHFeQHlV6oCbkydVieuomMpp5BEIfBNaFahhsmThjM6TOLHdB6
do4WbI0SytcH2q+H+AAYC3h2HSpE8zOZ/Etke5Nt+Ue1hfEJje+quuE3kSJ8
/xTM3gzd/Jen4blN6uZOL5WR9iNAe6T7JSsW4aWuQyDG9jq8RVpk94qwEDp4
imwHxsEZZ7K6xl3/lkIC+fO7qMBKWysxHa7594CqVZ2KjzMz/POj/pf1oEd3
UKibD+fXClbH56YTnwPlxrljaqJ8ufgDla27vBZUdIYyoBq/T1jrCqcSn4Fi
509Et+9XBBgGItcF5T5v7L0W1/8oEgzaKldyX1qFze/bROhuMBoZvO3t7nkD
PBepP4eFuX8Hafc8NdaryNCFvsrozrhqD1MofX+6fipwVlw2grG+JMcD/AKY
Eobdip+DOpbBgZvCr+61kqVGxhHqikaOXLK/IilsI0su5As0CgpuSJvextwy
79xA15LpVRlFHNPzWqWwRWc5boFYNsgPe/MIoFgCd18aKtlSx/JUux2gUN5G
mrRusFz7Ce+DEBpG/CPNatOof2qya5XfWOdgKR3plf9GG59l+od5eNZx6vd4
tk7XP1Root3UMUGE9UjSn0NVbiqMJL7OGa02keTr/Iy2fMkY/+5Tp2lcP+gk
xubFIZXc6dnubN63jjlXYkasGNwRUeKWgixjf2EayfAeNzDf9HiUVBffjPzW
JgPMZaBRBK30L5eWAPl28v70fsjpfqisxds6dKsOtTiVUa9QwRvR3vUM9sRi
TffQDtQuPy70zR0SAac+y/ky+reZchKg6w0lbMbl3mzDXScpyVO/QEOl/V6a
7AsVONGz/DerTt9HQEowEU4Eb2pOe3z06p/321sgfWLbOzHAQM7L6sAbIQ1n
HkozC1qbz6KctUjRiqY1YnOlW3sJriGHh6mEP+io0ygYa/tHGDshK1IjePJ/
5QJtzaudC8Jb3xeCrk2zJ2WF5LpLqv0GNeHvWkpgygElA6kiCzhQwCeco+zG
qV6ygLg/nPRf8s4wsp8ZOox66G7KT8waf1kQkM8QQLaq5rIQbXQzDGI5NjOR
aU5ZCjbYtt12rWhiSkEQMh1V3xYTmTWvWncRx/k3yMnQcyDLfZxbeCsbp7th
LeGQLzz21aPsSOZw4ukxLr6DAPoAWGWwcHLkhwOj53Js3NDONzm/VdnwXNwM
WiEvpZmunpftELEuP6FlyyapC3+UtnU5rxOLCSWxjdl0q0TdQFsdH1KX79bl
jUEM4YWPUdVd/gwbmt4/zOI+aUTqIuiEdD6ua8RNl/VJDB4Le4e0suwcVLpX
oL7oh/Tln2HZhOeaA1tvL+W6iy/3N4FhRVQjOyPw46MipNYS1zRQ+u3fowRb
tGmbSLL7+Rky1i6dI0EkxFAXoFB/BX58rntsh+bXmeiEyePCbPisC8lNOyie
q74t4tgIcHNzOfxCxMcLXSbDH/BHSyjnHhyFo+8vvAl4IrWYsTlknqJH7Wi6
qcYneZ6wqVOs8pON2jN9u57/1jyliDnSECp+Y9ea0ickgZE6dbMKU1FYVI0Z
fXdhdG7H72mjEw4v/LKUDmCEt//drUNpIncljpCJgvDX9LOd38ziRkcOPx+k
Yek0/84cmqOmLlYU8MZNS9wVIvcS3GlG072sp5w/R74R3Pn71mxqr9tnnb5A
V/C8Rj54oI5zBdRR7gSceWdSs/2z21SQPWQ2OBk+IvnFP4HLWJ019cYTbZ4R
R8HGtGVT7x8LRu+4gnllVMSWfixhbxGLRLE0/8S6xgtjKrxrenT8oUyrny6D
78GbRm4H0YDO9ZNYcNKjGJq2m2jC/PcKzb/JJZDm4Tzcsf3CuyOD6dR4t9XZ
R60Kwn1JbngV5N3HnVQsRk55oas/h+s+v/6Pqk8NRkpd4hnsBFcZPc4qUhyL
riK+RFnyXC6pPyVBcCoht1iptm3jP2yjF22KDDyjWpgdBUDLjo757Qjj4IFc
zYicImMK3zH2KtKo1fDk7MiGr8z7PDVpyv3s3aoTHL1J3cZl7TAEVJ8Tpghs
po29OPsvsv8yv2ygeI+fLNpYhpeFCOq3+VDNJ5WW5PPiAyGKq1QLMdRE9pjW
06fkdcvdKkK55hz2KClLe8KFmOT51P1nilzOqa/zjUnABdmCp0MONJmBgOsw
pbBI6//0kw4skTmRaRT6n4wPFJEsLPKq4tXNYYq290UCE9FvRwmsviF8OB8b
dUmg5eb/y2CeYs399+qKW3Z4q5uSfPuAYle7FCpITtMYS08EIEgOnwsG8XvX
+JrAVo1RZTJ0vM7PWpvQyEuwjq1OWwEVKFllyOd2ltg5KY1Vnv4cI9rtv/IY
XhXijbhEdYJAJjupFtCXv0reIWTn5yh2yIutr2HPfNyZEt02DYccbERkWMJN
xeOYYNMyXlkcbpCvSZZtcO3/WAsMArjKH6wXALldnIjINvF6UH+US52DerU4
KPYOQr0gEdi6d1IhTxShlN2f3uLq91xRtDqdsQ9lknsKUx5i1dcjSrvBHvy9
stcLTL7CdzOeZzTdlRqAJpuZKTQzwBk5XbcvvRAEMGOn7EDzqq70+f0UlhSX
ZIpZWy7YS/Sf/AdmHC7nx5sQsh67Vi22mKXKBbT6Yb31UB+fUluxNlc3/1fC
h+qEIX4riu1k/TmatURaLQzW3bDLONUMt9G+HhPKd63JTZtEZcjfFs1uW2mf
3qqBs2mfxaNkuHmjFlPFDksiYwKtP20wy16h5Wjognst3EC+iDKeTpnz0LKc
K9Uzor0z6Y10yQbU+N+hPlf2kZXTp0nBm3A2jENdjiJ1XQPAoWOTfk5B9eyx
W7aemh7KAgTVe+EsQ5WsbGlvtyyUQx+fr0ru1qzYAX18dHkhiULR9iFTFHo8
ajjsrASugcmnCMDe0NSr5x6X1+xiRkU/Cq1/6utzoVueH3FvibduSaLg+dMi
L5IsZ9Hyit78SIK9C1rzV02WwYERt4ehJ5AtOkU9gf/itKLHBQSl99Xee/xc
Yl9Tl/JdkAeNRKvgppabzJxqaWilHs46kCp8Wp9yQm7oYJMX6LaWqhybiN4J
DsIDjHNl6jD1b39l4gBlFsq6T8NweH+euznLM7pe2eCs5vq3DnO673Y4pUml
lLPNdoYe6A20f8TW3fbYFbvMyK0BDlkbFrL+9SClhxbUz/5ldF+kxat4qA3a
R/UT4tvXccXA/00sMIh4pu6diWUT5uDeb9URFqcBpmKkRZan/9r4EGdEnO7s
onh+JiGZEYyYctUeTrLtFBxAQXe9dcGkEQAVvnbXkdJC/fntCuAzHxhYEtB5
nnzvgThMv5CssDNxMouQ8JZaCE5CANxgWXEXeh8J40RNqw3X0dvhNlGxhN7s
Q0+a2mpU+fR7eSWNdyOGKyhavGkjGP04aGRQp/RXzg6RYSJbGi6YW3/R00OH
fQyWQMPQp+YIJS8cKonv9Ciq4fDZfXvt2S8wjfXZfJ1u0xIxmBwbjoRLeb83
oNCfaUoiiiJvi2wnV6xo+i4m0vzG1dTiz4lMbxFwjBsLoslno91JazVwR4z6
dHG3Y/yLfZEl9dfB0BV8XzUll+JumxVeYDjexLK1JKpGC9+S5GSlsXdg8ONu
tGiM3Kw4h3M7j6Tr4nopYCDYxVSwEkpfzknwrRACWX3N+fZvJ+gc3yz+feB4
CxdjbsNEvAJAGTYISANO1zBnczo4XVr4Md/qNqCwSjg2jPWw3oGohNhihjsT
bnKp1kEN1kQn9k4b22GFFo/FbVVwZXEklz//vSFCioliFr1qt14lhj9NI4rv
B+NkY+tITn4hpOvMGJ4L1SrIdjjuwGgLoBVeDAx1bZmj7UzBK+LFJkA3SLU7
9FS7ctkA+suOy8kR+iK58LDmeJVBDLBYTXrCpPB0wEOgwoOVKalvfP+27iUH
MhzS8K4lF6QMEqssSP416d+zUhZMWvIK4nLpy0LCulSvc2VB8UIbsRVEpNEh
e9NxuNrjoAFMlgOlv4H6ROihy8X/5R26ZU5CzkbE+VgCUW3nT4isXL0b4HsB
QY8hqjvs68dJvHh/Z7vP40+mreorLH0JWiRfEMhesPSUySLbOVMrjfUloWlW
7zoQD+Hjs5IFKF/bto0mAp5uX1A7gwiCguGYn967FS4NaGUFN7b7DS+5BEmM
K/uvl1g/cbsxiHP40/rWp3U6Vi8u425CkgyeObMZt5XIxrF8nMdAK88GPDle
kOLW/OEaYXqPBRLKRUYi0Z3bfVfl4RQrPh1D9otcQhr6CjDPit5EdLLABiqH
+gNx1t80dT6wHXKHRM5pdhgVC2v7qRm6nfNZwN/03xnAlph5oua33nqOTj1a
9ODvtQdcZrkbBUVv5K+qd6aG3coDGymIi1jOhVYVttlsosHto2/JloG6aCkJ
ZTbM/T2/XQ/9er1BmJVDrMIy0DZV0/GwtVDpJBi2uu3mH3CLWDquq3vsL0Ok
DxXfOHLX3cZrI9wwK9djK8zMNY86ZUUREq+g8MAoV5sA9WuxR5RZBUWWMMUI
Pw+CkHwTODM01ls7Az0JkjjOwqqKBc1dCvRm5+K+229j0iwVrSz4kYqzVGBt
kh71R4p57atoeFoVrd4Oj/H6vlQtwWXM3F8FdH+3+I08u8HiSmAwS4k+goCK
HbisPJMmVu9aTS40s3L+pid6ckv2GJYsEa+bZ2ec6vTLnW02gtWmSaP2mqju
lJ16hiyzc4CYCdludNtvh1NCa5TzjoFSiahicGTU65IW/tG9Y8W3i4S8b2TT
gPaRqYBmhhdhMHxebN0goVk3cgIs8jtjDJdQxkBGPPTpVxHmrqfA72GyfnJV
a2CfpQd8wy5r9zclzHXftOsLArUa2g1A9XxBM0FzuWLp9XXwexswNt6qhtgP
EfXnyVr45avb6xWKPGlJdt/WzoW2qoI9w9ZASMJnJ9dhBWlDr5i7ik5TCZmS
leV0x5Kvy79lrA0u5az2UK4pk7pKkysksbXC7CX0VLWoPToU/G8sWJ2DRwpJ
Y3kxCVpI9F+kJnv6uQdxxvdbUO+QT4+NdKafNoUddqg9gvr9eIRrRd1FqSi+
YQhiH1I+MWHB7/T2qwF+OOLRaibQYL4u4XyTNd9DdbPmCE38Q3PIa16xMIky
5yxYu4SZSeSWxr6cLRjd4s4Coggl3c0UyE2IY7fZoG0Z6KSLNFi/jRqMhjOX
577cZEN+XJK7f3x5Kpp2VuHeJTEN0aAWzaPI3YZUu266C3O+qd6/et+wAC2r
qjH0CXNTyCakiAS+q75IQtePF5aFlkwYrEioLNNIIGaE8t4einQK8u6DIMg/
ei0CJbW6SGJoutClssTIG/cNCQeCBQLDhfpTjzyvoUvSCtsGWI9ZhYKsOmEn
nBhoKGMky9wef6TWXgE5InRX9To888gBk0ZeFY4XcS08m/k3p8UdVJsx2SS2
NuvwR3Ie0PhbGOCRTXgDCZx7DqlN2+wDxy4oYEP/NQMDNwFNMKxIj8Tasqcn
N98PjGBU0ggqtt14eDOAx0zjItKFYFSwk/R2GztQ9IWzdQqKHdNgXJXGfeT4
RIX8++bELKDqDkVuW9ogRLNqemKits913MMyAkAW1hHPrL73sEWbT+V9Y1NP
4f70NB4inWJ2HElyL7LtpLE/MHPqGDK5VXGq0OAu5zgAWjnTwrmTATOVl5Ma
fxclprtRbA8sXunggXiFRNh4JyvUWEmtEJ1EwQqF3VcfRj3v9Kr1+o6s3X5q
BPo98+7pTx8ZjtaVim9PaugkG/4LINbYVI8BEncVVU1UIZ3xCYD3CixaKCLP
KUo+on2d+wFE3WKiLwmvkqyk4YFer0jdlnWYyvLUeT3aCvlA7pQzf0T/TXFB
+8o6bA2tGPspUtCE3RgSyGpOmXoFwt2GFL8uPraT4psRC1qXDDZ9/a1GZmdS
LLsTcaPahzf70XD83vGoihxs8m4km7xrGnFCoZBZERCDWhA5q5M3sGmSW5Vx
GFeMZnTbDrjlZbgqicYwCQqymvieOoTLHDHJr2dbyqNDDA2dgehjPxFDBe20
h+7mmcUk9covuF78C80/B2oQtnjL+MoPBcIYBsa/drnVh8eDpOrIeLq8vAWQ
VsriRcICWFn87+T0j2nep1OjmHJG5RqiKTG0M72Rg29sNGAk1m33xHlyE0nd
Bp60gDVvxJkvcBGqgbY1qVrSqsCH2vIHYQFwAaFdIedlyuRx/M0UqBziSwgb
s/g0dsrsyvuw0tNpSPqXo2kCaRnFrBdcIVv6pOWMLmBxuQPFalt66Nq82Kca
4QsSFQEbhPT6ruxJAj4kQDuBeMs9nZwbuwSKP+htG66+EOeZ3qMfdOOf+sqf
/L9C34znLZtGwmpD+vC6cK8AETKbknQ8dSN5I0IBI4MGxAZJSUb9BezbBuyd
zuL//6VvJ1I1I9C9B4uio/xvjosOiU2w8n5Z3PK3AKn2UDxlWmpuZPi2eN0g
NTI55WnPrO6i2Ar1kCbbwcpjEeRpSbf3HYalMRNL1lvMle5WnuCiZghoCXSf
CSRcK3sbfoDilP5akYaoZijy45HZvbGYC/snH4jF/92Mfnfm3jTSq50szI7h
HTs5iHU78XsmgfAAuy65QhZhnTKRPi37FZFScq++kvhRv7GmbV3QQn2ttw0t
SmJaQOMehp2qnngUkgvlsNjExl92WhiXHGbFLoVYunsJl8BrHvHfJwvYwj+n
UybqMtW+7OchzcoIR/M+N10rgO0Hubr8pcgCuKkCwHBsSuzXn5yC3Ns6vc/t
3HMFpCYjPms/oDlNsW65XJKFalEAsGo9yy5BXtYmJL+ujTp68mjsW+Mk0bh2
wPtfQttFd8NAbxU7NTTVwsFL/Bh6jxTF9rTPRhX4Bxv/jMHarVYHi/aW8wkY
8bvVmepynDRpoOhbNY3QedDntw7S/ggoEuWNl4wLgGQp5pB/QSQ6PTkx1Try
fr2O5abnjyAXExsTL8c6o24JRB9449aQvP/a1EdJBnDxze5byUqjna6cMPTz
rYVMcHsoOra1H1rrSy/ktEcUTE8/46x6VpJmAG9qfC5eqwTuRXxfuFNYMDEb
6O/0SJze5k4H0OVvY5WSvhHcMOPC0PVhAlNa4izxwhrpjE4f1a7KSsaRjadD
kxKPq+wSzAqf0c/kcs640azz8CxytCFLoh9PdQW4oMmWHEkHYSoFLfW+UnDA
ElqwkYIh+JrfLsLNSyq2fsgUN4wTR+axV1w22AMAJTqddjH8uai+BLmdmlR4
/Gv4W7ykxYNYMZApatg0QxhUbwOOjtrs1dz5wpsfcQSR+C3xajShPf5kAcxe
ZL5FCNULxmf7oAV2I9auZPcPgi6tahh5v8d8SOwNQSxFm2DJ7qtYBQ/rtqfV
VTh9MJ+QNIfSJG5cr+rr4kZezE3axPgH3bsDCPm78pOPfZyMz7KwlNZ60TUF
mhc09aWDcv0IVxT9Bv7O1r0OUpqk+IZ2X6BStB9ls++Y8+8/m3nFkJ0MDFWF
vwQZGLY46El2b3qytK8HeXkn0B460UE6ut2315oJ+LjFj4iBBwnp/b87mOTT
ZbdEdihEKYCt8m1KzfKBJoBo2MwA+UXu5XXsZ+xzBa+Vdz2/B9K10CNrlUme
477yW2GGjknLKm5WVfoZadYpAO2yz06/6Gw7HXjKClpZXG5gc74217WEdVeu
qPcTTRuAo/u5zTmGy67zBoCyl5aG4PrXdXTm907YKOXxFMKulCUJmlNuWPOc
HsEDKSILTGiKkGAISxaYwoUfX0PuNhMpa5991SXWAqm6JM2qE1cFKAwAQa/T
djh74vLjo06lO27uYUDQnKrvo4hOJ2BTypjL967pTbqT6MNN1VqK493lg1ae
GsjykrP5gd2U9w/OnEMjoX3Qkzn4pZrnjD4pEK58fD0i/FoFjemHjK0x7GBH
LdFRAf7ROIbdN+le0Dnui3rnvL99LV2iie+7vD0+lgQVwMBW2khHeXaOuYp1
Gf4O4MiD1tkH2ngInUa5glUoiDvNo1yEzClpOEu0xuAnatCfCMhInka1FEeR
VhtZ7FyjV1D6xyZpUrHX4qSm18H5O0MNuktENoQXa55EAVI1rKJ49NOdtqth
HnnlWW3AKP7ul2xLczPUF0s4ZbqWtWuOO0gcyk+jF/vUs9+e+4XSRACnD/bD
Io33ejy/J0tpyQ27wTnV2BFxrErV4dPCLYz5ku7Zlr02Cx1R5Y3EVloEwXEY
dTe7sJs7CSlwUikKrGV57GlDGmf9RL9lCeZMocSzbkO/vw0+/x9Ut94KIrwP
5ABU2NzdF0/cyoP0FN8qcvr2yEjde1OWt//3cs918KbnX+lAfP58PiqtYNBm
MEnjtdy4mr5TNeNgXEvdq8EvA17cBG4w7HXXP3oEuE03/DD+dpAp7WdEsPdN
P6J8MrAoqCLJwS2bawvsqGSb91MvjK79eeNBj1IuqUseuSJf35aYgR/86A3h
N8sPpayEgUPZJy+BiWOuhZgSVydLLCKqjFnEGkKuCsMVe6hwXXbz1XhLw+rE
fg7d7etdcZZGE1uG2td9jCuN+oqsMQIINzh2hy/9uMmd1x0Po+d8Y4dq+vTM
jpv3+G0FeBeAuvZIrjQPCmdMg4DfSOrKJoxi2+KGe878ndU/QklqhKScVmZH
hzEfNUR9Fgcm5Eg2OckSjh83zvCAA5QpuoJqLXzwUCOzRbEXsPPMMt6wnZEn
iDU1YAlNvjKY6cKWpZ+I0qSW1C5SgrEJTXTwNIN4oAlt/bZPlES4S8JKhlvZ
d50z+oOE0M5h0kxgcOy3ShtPcdHKGoAD0XNIE804jtTDRKmr5d5Erq9wIa//
Cud7STJsuv607DroaJ/l+j0rzPiysgm+OQNzjIn3XSg5p8i58JHbAcrnf7VU
/WlSUUofuGX77YdT9jT5voylPp7pnmVPy08NLpAuFBX45tesF1mtTCjdQnW7
VI1n72FMsp95GVUe8IT/yCwUtFPeKQkvWEHVCgsmsjlbpLoasX5gYdf3TjV9
s/4G0BVpb5AoM7upd3Ios6vm6wZXS20fNiiIrcBUCVcML6M/xSyhRuDD0llF
nk9HoUSbymW9nctLoygsAYqJAHHBCCEoPPsIHxvJj2TcOJFdoJ9LP5XMIJbA
DoKmxKQf2ctBnSN8vGYlkBCD8zR0BQkMSFD01PXaC+f/w8WJ3aMZLB3Ndsun
15RC7LHrE7EQu45AJCBpTGitAAzSjubZQtSU06TGTx0F8LR0x+Nj/7B5c3Kb
ZBpU/RSqx+SDlE1/ooh/jWJgJWLzr+KoUi0dIhhHPJxtGY9trRHMne5wRZnM
5jgcP1baCObu2T3N+0y81Q0FbBOtONJ0JZfJD6qmq+3sCV9AQwydSg3a6bIv
bPAgcocOIzBpQRMmVlwh/gWX6VuhN2sxWy++KSEcmkUcDAro5SI/88RtPXhw
mIbNVXt1Zl3FtI0E6/jVJEmP0LEajBYUDHccey+n3V1kGzqhuFKTV61dG7Gt
mOc+Cb8tuX9sIyh9XwZaRBSodhSAosSdv7GD9dOTCTtiNYYxoDlHerbCjAx2
gDSAIwfQA99QJZ/+8lg94FV1UVdYfpwq6peSBWIK05t8c2RKvhuC8KedLJTF
ek8wncPm+Wsf05KoOf/iSkN7NmE4Ozyv69fcMz+oMec8ATY4XO1dP0EEO/j4
GcszQhj+TTk6Mhx3HraiILS1f14w0DkVtxeHQ2/k0sgik4sDm39LnlCSHUc9
IxbCQXlo0rIv/zPNkmVyPrMIG799hXrcwxfgWOeX0MYFm6ey9FoPZddWe0/M
Xyc6c+r4kzOIoFErZwXaQSUWOzsSdnLC9tjxIqnvpkfUPmKljazb1cgZtKh6
ts5NjEaptt1rkcGTuv2DVJp6MHMAkXhJAds84P29Wx4NiUERd0HeJHO+vkRz
xs591qBAV43ZoHXgaBEDtfPTqW+5yXCQ8xhTw0SKF2uyd37dngbBzGFthzuH
ZwPZQ5UcQYHTMlxNgtaKruMLbL8sehhlwlhDswG1p2qeoE82/XneTiMtyA+a
jpkpuCMHo+NENwLfb8kUxygGtdVPQBcFBccbM80yTVU9/mvugrrD/x3U0yuS
w2jgzqG9cXYyiXxB69Ild5uA0PMUhwWgNzSNeaNhyPTq9UX4XU/Re3p/1PeP
CjOV/yhYpLqlqk4lgQzkhbhyOhOxay/g95Cf+i51BarqdqFGYXyRCkpsQW69
YebQPOGo/oHkJU9AsWUhOvWplLmCQcy20IBhZbjP3rb/jlRmlN140QGSOwU0
p8W/OTK6wb0eJjb4bVuYwX7e951CSjEbarfWlCv6aXm+WFvA4GOFd5MbTCjy
Fg5PnWYJqYlu+9QMi6HoE5J4k5ZepLzUAZvWmgeEUr9nLiMUiSXfAlTVPkdT
RivoQ3a9i2Q0mrHxNHIWZKgjXRr1DT34RZ8KTHi0wWQrs2LY61oWFNJa0ejK
hiDDfHpeuJ3iG/XIlcOjvRIz14HcLOOQiuXmcAuoX9t9Essbcxzak+uTAbsg
tAWuNNCJKhck3usa71BJKgAjWPvpXiQUbkr+XmOUXU+a2ZXCPxrA9GAkeKQ+
PQBUas8aSoRnPiXMypS8IK7bVyl7g84QiLjZmJ2neKhr80K0FHnzcb1YaJYF
D0nUop8TivCnHH7M/CmcbNJfD0FApiStpFxpMg2MuMhkfz+qkUVlLX7TtXuS
Yv8j5nVEcjvKbhYLip+4pUcjeX5dGT1iUt4PrTkfx5KEIAUAn6NVZC2uXia5
RpO+UO15lftfIQ4rQ6FjGQyY6Gv8DcC8SI/bE5s3vQ45rqmXxYHisq72ZdqE
Y+zFyrPspoSQT9JXw0tDR87PgGLtr3LDwvHznQPENaip5V5qagfQZiw1esVs
nirFmrx6eHoaDYhKj1LT9FmTMaayiVHZUJs41WHb3HVjVDZo1RkhlJTruwtO
p9EcVAFnSxstb1In8ZnowHXCcQiAUh8C+BrIAZl1VaGE6Nat5ZugRcGqVg3g
IEQ4qkcz/j1JO0s74nJpPIflSW3Ktrs8fVzYuK5ueOi66gU556hDAY68dRvm
6MZWSaoIpPpcMtWxmIZ+cxKt9DfAQ0ITlTgzEdSoDv3hpK77kpoI9xrc7vFk
9of0V9n3JduyPjHawX43Xm/Ho05N/BOnfVN3CdAfhtgZECMx1uOzX/NOBsNG
OTeHvhnbgfgRZ7NWsyLKzyuJx2RZoOdTxojNPnDsMAPf/f7FeDNujs+7BPzY
j+qs7wqZYuwpyGeSRMhIOGitH/SHuQqIIqeYB1ra178tKdjLwCvq6EuQVtL+
Y/a0aUql+HXOnpm/vDt2l5v+N3rq5dHteYfb1TsYppJ26VH4ANEkymapCDOr
ADW3XBRGw+MfVr2o7bLGO3iihhMnHXfHey00TN0MeOxCDyN/4DYvIHfqJgBE
22/nxsjEeKu6hilo5qAA8N5st3WiPFBbt94Q4Nxm2BxBdzEV0dYWKB2IPUSH
IWrgUhxpGnLKEm7Msotsa5HoeoDyzipz5ob/Zqt/walYsTSymBZnYfy0XMRv
r3kGT178o7IPUsRVo8D2w4UNTZcBREL0X1rMkK0hJH6HZ8NxIoS9Qwe7TFMr
asfR0uSr5th/Ij+otdyiz2lhk4G1K+JbImx3LxqzTAfM6OxWJnV5Y5mT0/sp
Zum9n4ZxVE+kCpjDyvI4AcU2XQk7ghh9O9z/GukhLZfAFaj8xK4NZR202xON
9z/yGT5Pl5Qh6grwGtPfwnnkewI8LMvUOQn1BUHjHsy1kw4oLfWoRi8KAz/z
nBrfxDGNygYYE/n8iwUp10Zic+n4X9vrWYcBHnzrrg+q8Vv73TBOQNjjnJLW
CE/TKtPmq7ZjsNHX3bup+OXsvHyNK9RN5f1g0LswtfNtUPhIoqk55qIWPsuA
1bmdvhpgvgk/Gfx3YacvdYoyCcjXuGQLV2eq48/Qu7HIE2MgJ79sjyc0Asoa
tE8J/TwCzol1as+0Eg9vlEwNm9sWDx/Dsg2sQSeHnvk6sFcHjggqJMjdnWrL
3YNtwvrZL7pmK5zc7//Sy92JpdDf2Zy+9+I/uN2mQCTZXUn1uPe9ULGCaxz2
TONwfP3OmXJvmChLuxOKAjtRWvR+lGfEDefjtnKaGZwBEeceswHrRXZ3rXBa
Vt33cSwclVGGfQY7dmcUr74a909jSjh/noFjmOddEV/+ZFNvK3jBzDWglvWw
V7eMt1ld7A4cY/nV0xU0p0PbPnijKPzjMrRGc/QgdrJ/y36HiUHQ2EIOW/WA
NMgPmohnl26GUT1J9pD+EIyY4DYaybvSxWwhCGVr61FyTGTut2xvrkjK+70E
hGoId1MzFQtUm6rP0SxrQnqkLDTE4t17CxTJbh/9JcWKVyE/v3S1EfDDBtSN
fyE5RGuu3UbWijf4q7q3QWiXTO86L1HewI2wH0WkFbzpuwP131+Ge7iWjBmo
SguYTZGrQ9MYc/OgWClMXLXElTDIAKMhaNZZdwSNBUCmpOvZtLmJ0b13Y0sG
fFYveU+14IDiMCB+D/1ejdaQ0hMvZ7J7yWIqV+eiTzomWHc5OdPpHSUXhVyc
eazua1xibUdhdXKNnT6pweF2sYisi0qik6MFLCtVK5btqUA3TTjLa1ljVmM5
yrEs99CLjk+GpxX9JbPxT8v/AamHjUzDB1msMV6NW3072LqHHUL43/PsbUVj
F1oS2dtk7p1EgRevRo1ma4NTryrpLELyR1eNUpkVhPzRE3f0Vo5Uvj7aPKd/
1iHo0mdobLGte3UC/dfGgR6CqhuZm+RqUIz9Huww1ieHUoke93ePs/Z5XL8a
zNE088/qWXPsM5ck40ldmbKCKSg/9o9Ds5SNP/9V4V6CLdBcbG8lrvz6Zp+b
WT0qxdLwya9ClF/yLPekC3cU3mXoK5BATCivTjJal2vxG53HIz4QI5nE3uXg
yG+Y39GQ1u5WqGrlJpXvley2fhAiiZFjMQOV36ceJQDkvHmJ5kDHiSozeWtu
yW3yrkK3zeTXvN5dYcPgZ8Ahjxny4M59+dcvza0XuJsZ9dUw6snJ5eOLmHGX
KMgo0NNQtE8eUQ6sK45vhmZX4tOjTPCursJM6+B8xUK5Twyoc5aCWrNf6rqX
dtBLPex30FdOwTgGm4oc9JhF6qyefnQCwYlZUICmMDRDOGrWLiA0j3jLpK8s
YgqUb5BFlqGoujUQd/9lofVaiDNvIIg5SfzC55lIIwJ1UXgtlq8ZMoSJPO/o
TFFntLUUVzCVUcgwUbPjcnSAe39QWofpAKdi+XsIpLp5fMCyuL5FM3anfpDi
sXLdoMKBMyAEOJBsxbBM3u2beruebDUufgC9fiRlCzcEg09Dvm8lfj8gcqZl
iEci+Mn7qk5Lu+wn/pBUrIT+I63mynkJd6YSC+S41ANprcZpZSE662/q0+7R
B86/wPVgafS2YZ7PfwIjP681TdgP9oP3cA5RR7XJyz2cGaMK59t/HADAV2To
4cNS3H0LEs7x48+tnfmTh51GVirFp0ujplLffgXxYFJVegx+D65wzAYAeHSW
Q7qMtJMHuefIYA1nFquyPYnG+Z/f3+aAkFxNyZ4S6624CGXbWCbnJDDauEZs
xg2wecG+f7ThseChFp9ELdJOeG4qHQOzaqljBveNtE2YBWWMIwq8LcY3UV9X
OrwCVx10HkJwmovcPDs5GotTjoxrH3flT4CdSacs1qQYiaMaXzAL/ZIcNTOA
77ZQwrIRgjCa4EmfsBvcTOa36XQK4+CFmknQkJrkxRWirgEC/vZ79L2dsjL0
JqG3Cj47AmQRQeC3joiyZeoV1vqKLsK1v/L32IR7W10Q93bHLhFG9Ekq11MA
lzlKBBqbw/X90LDJj7fKZZW12x6uxWCVNCc7Ski3iGPTLNFaCyUgbab5Jzj/
zPwqZX6lbF1V8Mac3FHLB4YyeoaykpMZKfg5eUs+DQQXbkY837AjwNUf8Ijy
i99giSqvxV/y4Ma3qXCzD3cF6kl9yaQPBzXbLw+NjJSOMjQnCBgU+sdzD/2T
MH8LxwrE7V/kNHRd4uB5BkneIh54BQWU+SGAfy7HWnrAmmTqYyZLgr2lAarX
hohSO00CcZdps7xxFoGApQrU+ykMgchy2JXy20JYK9SEBnDd97uChazhVbUt
9xYkUJxc0ZXanHLKKYB3DBCb8bvLWGp2eqHwU9pEWWzaNVDOUF50ikT46gnX
UM8lw+6kXvbqWDoUK1iNIALu8iLEuvW3sNp8gQXu5F7kEChII8WGnLMmip15
4v5Uc9UYN0YumNGGhBkieJwfw458lkeS4Mb6cb7G1bm2yU2ihG5K0PhhDDnp
K4hvPbD9u8SpdLPBq1exynizQ/IbJoFyNT64Dmy0hmsMhTgv7UAad6PbHuis
LBkvE+mwN87o0sJrSI2y1wkhglcqCmYhcPHYgN3uS+k8X5FaBgYz0DmQb2+z
XMnQ78I167+yrN0nYjDzfeblWapoShFjh8X9yTuCi9uKX2TML99C06aja6TC
7FS1tUrFXUz/R7Q0nto443elVEOHxh9WXBWg00gB+GMN04DhElQaDqnqACUX
c6ZylnRlwU429AaE2VFX2dIGv9TGrZZPcNwh4opFwYAwuHLcilCQscw3LPHK
BDFT76xwDFWE+u+YFYIRysOPlJFBbP9FWLh4cFfRCVL8epWSPlmGlzfnz1vT
sY4Z7Kjgr7xvMvsBshWi4UWU0Ucx+4IL5w4nPZgT7XolcCFcge6tkuODV5aG
UTfJHniTjmIWremksQlknWdtEqwwzZ2mqlw4J+uD8rE687nI7JQu+ZJiQLrI
QfD9d8DrfAJyNmVT7ZBj+4RjjCEbSYtGts0746LpNtUA0o2d8rWXqAknR8kw
m11Qb2+C3O/+39wqBp6JX95Z+MzIgmNHwC2X5eSEF29OKRsknsN8jlj/4hIk
z4mKm3R6IGlPkkjfCDF9nop9vnCh0YTBCZnV7x3M1jLYCRRrCOl8agUaXURK
lwgYFDpHgdamWx7B5SpJdL1GrBvql3YArYIpX9ZNW1OFBlRXAbFYyz2uN8LD
6jBXGDkVi4WQ7WxMvvE1VnUg/POxkaIV1k+SlJ9zdcuuvv8UjQvfbwY+evL7
UuZrw3Ko4T4BBA5eDLQBue435Oa/x5r2N1/i4xW7F66qi2u7S6jLu0SW3Ok8
M1/IErQ8YdQ7FW/Nh5Gh3aenrpFi+39/Efmto++WSAoGLw/MMfg8WI4YGPZO
1iuMW1Ifp7utGdXEE82+6FkhP+EbsEiT2VF9Pk9woCyj2DsI4L1QIim5BIRV
5kxTOe80u/MF/p40flOjOrcnMLgq/WcM4vbrCLIPHtp/4EcXd9S6GgUmvkCy
3S5MOviXkHc/FtAGCgc951ocT1Gbys5ivMr6mkMFLUaIqeoRb+9LmXYPKZ83
aSZsCclZx0FLBDwiCCfh0zVkMpoH2OG+9oofQ3G7WNVQn9saEFT/U5YwjH+A
JYJqWOT14HmjczITijNKVWaGUCeI9FdBfq2YJqVO/3Cw9aJWFhBNTO4D7fx2
TrccUYU4LOHAjIwJeLiTuu8iQVmjReklgzoOFe8PJ4qjwvWXcECsfqe1K0jM
F3dMQKuyA3kNWCqxwtkESiWLOOrlQlO3/dCcKqQVQTlfxdc8thieRnrNERe9
vRmumPwLEof/JObfAUKt8WFoX56hEgqJxWJYpkOWL49LgQfPEayLWmYXvjR/
FD2j1Sw1oE0gOLfSeTVgMk3Zvw8FQBttJnQOJxoz1dyBufUBCw2XU86dOBL4
b4cFLc3IP+Wx5Hv1mnnZ3QcCm1MQ49ouaI73G4Q5gC62RGjzBZK11zjKeEF1
MQvxXFW6TFvawSdUAQg/Fo0nin/UNkvKQcYdU8S2z9wojqHz9v1WMcbpSq5o
fDlNbcF3RfSVYCPXSow2/5u0LHZj2Dl7D4pPkDi6D4S04UaosUNPlYPp3Q56
p6dqk4QH0NilcyyYAxYlvp5slCpBPKah7KF4dZUP7HuKy8mbWvBYuX4Y9zJZ
malahYtXMxUtdiRKx3GHx/KdCQtp4oKWBcHT+L+oYV6KmXIDlmEHtt/L3k2C
KGHiupdiZ2SulxxVhHvC5Aa1/jBAQjZVZl0ePc9oxW/7iSPB8R+rzf5sB4C0
7GaCeuYrW4WSxd6i7boNdJjFCk9VdOor4LGFHBDi2oyxRGLgDUbQU0FEnpdE
yN3Qyrv2HdmnwzGizHsbCOA/nrfJ6CY36aeMeraQnlZdDUQnm8eA1sFfXXpF
ZmRXhetQ+A2h+WE8WsOj29NPPYeLUOi7ZQoZsSimmh21hRnR08sMdZ84LlRI
qfCbUpBraqTzYdqPxJrC+s37OB3+SoEqSoBgrqgrLesKY/IxjxGPUbaS8jXw
bBiuxFLiKmg4iVJ04eAJ549E83SNFfV4o18RG15ljT0+Qjj8pW+jBQT73Ti5
HMLsh0Mq8JxJmkhtxKzZ9ylSXzYsj8Lm4YoYEiPPdzxtTxo8RcpP2GsfJjhJ
g0MpqemwP7ywUEgMIwwhOWHSUjmZs7Idj8QbGx1kUhcOlVIH4wPUmcS83b8V
oCw7neHVckJZDvlH10wElb6/0jG+ZFxF/5/dzo4cZ9B7/6fLyBnSgMgIBNfQ
PmcJNt7SR4a1KKkAkRJDOTMBcLm3gjmP3byamxV3Eom0fkZFQGHHW1x1lS5y
dwN0xcUf1DOpql8wO6p0Tuy9sxxkyJfshqg/+u4WjSEtJI/3y3A3/a0zvNl7
B9XtLhqhJvBglNujBhdFxk3H13VfEoCNg9aAs+NsM79RVjlyeuqTTm9Q1qlR
LjJ9l//nZV/w2gNI5tJUUc281yrfcUNbNzXRZJKqUdnlUHDIkEyHUqUD5oIE
kVOnYJGoMfrE0DOY7zSJVMAxRlVJXSMrh/4kYNpfratGO1hPZH/kY/9ZFj9V
0rbgcuUp08xLKRlocnUO51/EsyZpLLJADD8pOg/k355MK68GJyUNeoEqutDU
2sY5Rb05vZ0yixZS3QBW1Skm6nNby0ByJeiT9miGhg12Czr6iV1YDFwrZFEs
lZpPH4IaFlS0AlGusWsYf9MsNsiltKz1jS+82nzflH8R6S8BokPhJbnB3lN9
s59DWqpI1BZKpkRWhc4Hg5siNsRsIH7nI4DiYk0GkLzJc2WcsytgxMbM29s5
D2D+t+1A+1tn0H36TbWCwAaP81SIj4wdAjaIfInvHaurrJEcWAHHwpA/hzHN
IRe/YNoT2IyNRn+uTey2gQwxZ6yQabqtgUQWz8Nq2PtBNq6j5f72VLG2nUv0
ltGjS+dGLxSVsQUypZ7lPG1vqatD/bhGOQeYWEpMn5gTb1puefNFJEkr1ZdO
jGS8mr3SZyvLlkcw9iC9mOSG3JVIs90OXiuXTBqjLMyaJ7LWp31PbHzT9IgB
nhFL3BQwAacyq1ZxZF9K5hascrsH8hVATN45q5jkDuLswUhmnc0une1kdK9N
0Do13pcWB5RXbwNr8aveT9YfKRAb2k7QQU5PjTclmn5zrhnMfyaMF+5rQscK
qA6w511Pd/GuKYth6glsFjrzytBVi/ym2H2D0XXeq8u7iXNnsEigHF7sbXfX
rhMhB+4cPUCpJXy/M6apunsRALMFvWex+ccnes/gMhiPMV3QiVPMwSMbzdSh
c07bIRW6DYfCPu/pwatxzNhLJFMU9Zf7iX6GdzLNIa3iRm0vurJsxr/94ECq
4alOVJ2hw55GqzM4Fh9lvytY+P1HTF59Wy3rLcKNswmaemFAAb2c3nQdYIMC
dfa2GNE3BXL8fJ6tpOWV2oXqhGpaZx8WHOYxQ8lkZztWeziqPuN8iqrGwLht
A2/oOaiP5zQAK7NVFzscgy4WT3OKg8wVNM3E7WMLwKwnHdS4+FRADzMkYz1K
mpWGQPdhi6EKEet9QacKcBH19X6Gh/aFJvikHyI7IvfwWC1tlQ9I/b2SFeWM
PjyRwX2tiuUsajgpHsuRPnc6KGV7Cccxf5n4kkcnWuCwLEWmzvcVwLKl0uuO
L5LFB5wY+Y2XIDPe8RN4Ej7eubEQ2ZFRG1UGwi9fle1U8BcH5wYs60OJ9nsu
z0x7bDlc0PiuDg5SyBhzV1CxJvc8yxSBnNOnzpX0onTiDA00FSH37dAqBdTL
MKEKBJl7UArE3tU0DpR2trpK8lEU2KXFKi3rAE1uzTAUWMR5fLBNqTpobjoW
HS7Mff8k2VIncbbSxB3HyLUrSN/E3P9HS+/ibRbQQJYYcxlxzEVU4JjFXe3L
C8iwUjpryMhqz2vF1vveC9msCBf2IHcPVNvJtvkbI4HbACuxMG+Q7TQN2CVz
TSQQ1jOLIb6vhx/o3Gp2Qi8lbLXmSkSVujFgTQzSuNyw0/LtTpF8bIazrf8w
AB6bOfib6B4ceYvDc3nAPW0ErOPySgXqvzB5LqtSxMG3d25gSep60/vk1MMB
wYlSjI9u3wU4GlBUWUDp8WW+vdPa3wDnTsvqxW4f8T/RfzL98Kv9lh62XCXq
Fz7mnu62rUCCZzRZIePShoaLpYfKI9Wf5P9myrLrtPOSgSOKlPMpVYw/DBzc
M976FIakz/jwwMnwYnE39Ls+c6rHZAr6LglaTEcAL2/4cp5eLX+E3hacduU6
vLkZwqNhvVcuiUK2KcMswRMAshwVIbWpT8Nen6SDntDqPkxjwE7wd1c0Twmu
GC4McGU0UziVK2YHn+LdcL+u7Lly5v3E6F+5Bq6E05UdPWzQO0Kois707zJu
B05ZO9qow+Jb43KRo9e8YVyR012PLEJ2rTYG90gsp85XX8l1za5hCI3IuTcs
kaQql7wCvofqeVO6E+n54Apb1sXRaYaN3xDQoy321bjKBh0W2ynOn2FXRtDr
Q27JMua2JSOgOHl7XdPiYxNNezqGf/WtNNkY8JkRhit6/3r4w6XR6MSJbrCV
iY38v60uLU4fqwthwex1oKTJHZfMHzkyI4uSpezEsaIAF5gWl7jHpC03gWR8
RZmQIKrYVKtJ6YF0SpBQrByfw5PRsyCE04wdMcks3WVbqdYj+0kUweb8TTeK
UP+n6TAjbch2YcI6Fg5ik4d/Y1ZZKRlYetNBZ22cwy15NNvJPNKN6gWK58Hf
PuC/AS1yTsFR29aMFTxtQ0ekqifzSUYTxcWgTNyX5HcGKPwAfoiudbB77AaA
ggUJTpxhd3psimUI4XJGqOd5xriZXF1Yk7FlxCSl+fmOV6blbvhI7K2/zKWH
IDc+HxR7uEsXMMtVEk3Z4RsJp+1e663jL2cx+1UblDWXsNVt1FB7unej0hHR
Q/QwarKPgQnYxsC3koRdMv8W9CS2kxBt0iualo/TmQADmpa5Jq/H4+nNxy0T
Xgvpt5T8AdkP/SQqztCA3bUhHBXrRQvx4zBnc/3XU3TdnVA5CRfiN9bxq1Fo
P7UuADnkoKmZhRdfIjjkmuXWaQAAqVHyMOutnrF3BqEc7+0YAH2TJMiD2/6k
f1xNecgzcm5ZlqBHFIxSZ9vZc+69z3lnNOAT2gQT1KX3Oy/LZ983MYuDbmW8
UIKcBV5pwGcsaeHVsF/gEW/2JwiSfg04wLZG5ywGpZsS2n8BsDNYejR7EW3b
0GMdT5FaNpvg+qQWr+0r3Ztf7Cu3xidbnxXexuh440TzmwCn4CdXqd9LKrD3
1Od+4mBoDkkuxnKfIgJNrs2NxevBzqHF5FLZl6xNQLvOLjY3sO1vBrE81efE
nbw8XMjTnHV0RTtm6G2jOYzsXDukAkYR1m9+C1UlkApddOi3KK5udr14VC3v
BI6SMVGBF7wnkaSscx2xy5b3X8jdNugVb0WuUEn7O78MovY92uuPRQxoOckX
zdpBnINLLBYl8Jy6DNiRlOSTpB1nURKLj7qSpNge0XfbylN22EdO0hAYqhUy
Y6p0SKi40dxllR7bo6G/a/IBhArM1bEOq3RDWtWSXR7EguuE9L6+WSvLtJ9k
82Gs7QZnyrHHsDGiBgJk90RYiF6qzYBzGe9uGhSsLWFmxDDuwZaNTT++WvkB
RP7+rpEY+QFUp8bKfJAQJi+2eDTcsfdxbHLNv2oUlXd/TOhZVbNs0Bprm2hH
67kdlG+SxYhyL1voN+v/tVpABJ83YkLS6UvIQ/fBYQkKt1Pam9T11KhG8Og+
gPFOgY1FtYEnVwmsQhXp+FebhYDsYTAXB2bzsjMXd4B6XJCoQ8jNEs+4O6vn
OpGym6yCKoXN51veQIuLMwg9iMxw2pL6URj2c6+mIHkNsWOixPzP80AO1w6Z
0FmvQjBbupZ1D7BxA16+MWvmv+FKB2x88Nq4QMZJCeYw3hANnvfHsne1qX+C
SiRJmYZMDVPk1tizfuWu7d4YaZgwTwhHe23WCa05dC6UZZzAwKfVQsFEFD3c
Zx7e4dzp+KEqpcWMIRNFiwUuacJJzQxANT9UrnzbCiQRZ4EQFHbYYhNxjwzk
KldCOjjE4rRx+3VR8kBWWxPxg5T6QWiQ68XQiJrr4P735s/ewN6RZDN8BXU2
uI0fgAcxJlhOVcM/59VQ6swg7M3S8ItWS8ee/ZMZnTPpLmQJbBVpdjlwx2JR
tTlgqThIxM0fNzLOkwWEEwws/19aaCK2nXOI74QHbAbksxXU+Z1WuGRxyNAb
+532D8daYjxdJkCcsNcYml3NEYhr2UutDIL1eMn383fCJyPRZCsWuKaDYB5o
IAUswxMd3VH1zdOzKVB8aEJwv2ZGOn2SV4tBxiGS6jixrly8kIf08j3OtdgU
m26gqSAS5r7Ms5RhZ90fuZEqGvvSclxLUXA23gkCEIV/O8k8ao+WI/8MRQMW
Hopdtf2dLg/AvRQgO8Nf3reDlzI0WXBojykr3sLqcrTDEP2NS/+0xCrB4fwA
fie4sSAUP3uE7z91grpyDb+SQssCmL/AuHtOCzd+cOq49wX7O8jGsjNUsCf0
SPZhcR5LTM2Anui2ro6neZoILIcGWRqn/Y4U0coXfvrTgwizyQnabKSncy6N
8oAX4ccUiXpfxLVLe/yjLRFhKPdRCv7rwfaLw5pULn77BtKvsJbU6Kra4ZEb
pKSheE8LExTjC/S97R4oC699qKdJr/M1Plk0ZIfWB5k/5ugeiyLeOwGZkzZT
c57QLgtplQqrFyVVkQal19WYsn2LsSKbL5PB9UHzAaXJmlqEChQ9kenWsTAc
4KJde4ayI5gsWa3gq6s3OU+BnUQceBXIQtr8IH+eonOWXOV8U/i1roRuX3ln
9GHLJ98LAh6+IlZTUk7yXbtHoA5LTrOPfOHobEIZaAuxlf6v/BjPKBQ5W+b5
ye3NGH5f+m7EjXaBSQtHTqNcQYxIXoPQ91FK2TNkcDCMOcAxTEiJB6zPv6eA
gF2Chp53ATak0UACwOrM36CiOskilF2XOHAUaNqFt4vdsGJBgT1jppYif5Kr
VOZbpaafK960Gd8slz2P0KpCvqXrUm5Fzs/DllPgXTzOOjKUID6+k18eOSBx
Oe+ISi9Spm4Ilj6Tkqv5iLa2HT1yTR5r1l6qnHpRhv1S0R1UlnzncGKCvbHk
EXLCavm3kRcOkzPGvOPCv2wH3zAMWUU5c54A5oCiELBTWatePofq6p39RI9/
USqSQezSPtSySRcTQYJBPlPhAKbo68iw5aEjRbX28MokboXUYqw3N0qKvnAh
zjZnU8eD/Fv5ZLHZjTofB/5XxExLzRzbKVw643ZvdYLsSF7uhcnPzbpsHdEk
NZYfLSSBVWBDUcSWAj+W7SgqLszw4y8grVNdbRjMopd4v74RZNTCJszXkkTA
LhRz94GdFWTOuCe1nGG8r0eGwIrLwt6D1xKhScD7XzD6TiU8uFvbJsR6wML+
7q4sW0BVmXARbbt/SEsM3n/5fHZfCv22imzNflLcxUtSECjmPjQpMWoOjpBP
eCQa4vLDRpPsL+XfZ59kVxrxzhR1zIOc6Q2nHwohvluvA80rl13QQ/vxdD08
N9kVH/gZorGCQLlvKqPjiAFaKpih9lXdgtTb6C/kIPAmoRWbnD8BcPU58Laj
4oO+zcNUg0/2qaYECJVHxZ3xKu42manYXpT73IFGfR77+UzXo8SqqREuPJJq
VnW1/kDJ/vR/snrxnbtqwX+p2Bv1VDDeVTe/HpxOlD3vsI2exJvpwYtCXZ2V
/xfnyEtTSwg72fcMW3QCgY3it7gbwL5AK/ntMehj1hXh/YSdN+oSZRKhZdSV
44cw9PF2FWLgOso9H1xzdTE7IgIn/BKd8U6ciPRFYnufHioRF3ZnAziievjS
KJTk8tK0sNtgrUkOgWVG2BB0ZGQpSApGQvOKAE7uezsAnK7uIztygjkkPzcM
kVg/t+pjY8K4c6x1MyDTwRz9XyNN3bq7WIXhTb3yIt5gNHNJtkMXZU0qZtY+
541+XpaERGlxl7pV/z0U9P28vI++1CZZjSuhihA1RV/eX8qUwcs1EWR6UkgV
uuLg0oyefrva1K9CINnbpCuXS1WUM3l+DjbuZTfbvPqHFKxg92yBulZoTzwS
7UWHzngsiMpZyZwSIKc+TRQL/9n7WZfFfggN/xw9hxsPDRF60sK25WYjYbGV
5DcuxDQ3HIqjkDyt59oGooLnD9ks/pRm2iLman+cm4utgl10q1JzOzQvjW1a
zFCxDh4ywQ+1wHFcMzbDG18wJrsijxwL9d7K3UrMGOyEXkMaLxIEjjqIxJl+
VLSQZhFP1RK2eSgIiQ9zvYWhcNlH/8qNyJ8BNPx9j9f5geGVz5jNJ+p+G4AW
LCJ8eV/TkSteNLklXpeYmx5NzurqmpqdXQQk+WDCKgH/S0Yftb8eyqET8PJ5
yE7KGRDEkFKEmuV8ecxRoGaGGrbW7W5MOMuw7YJArRQ+6maaqswCtfhDCx3u
41fvp4JzunxHfftvwSAHtWmR8982IiebePLga2KRek+pndIqYmK+uKjGIqpx
FOMrU59T3iWli/3kthGM+1pjJhD4hd4b+KVaj2JjpFEIuA+W607CNJ/dgQCR
JH7xW2wNbFgbnKMmUG5rV1+wWveww+HI3FcgCe+Tn2uYTjzeLHLRmhydvlcZ
pNOONTyK5lMzH6JAR1NQRNALacEFhFjPqIo5THxxK/pZo4rbGpUhBnMb+tSO
1+mQ4jrQtpKYLE2wLVgyiUH8bE4l3KPLRRkUMxIwm8GrmiOLYEfymKMCiZ+E
LQREEUI159f7SG6tkxnMtvHdDyyPRotOcAQbRPP+oEXGwej50qQWP/xMjBWX
vqy8xDDret4YLqDAJ0u0DbpLHSQ2cFYjMWJKvKvvwrj1T6UMMtEsGMLoG6zE
FSDYA9ooKVGNg/e3ieKx9BAPyQxvvxng7bbQVDiAcMH/7smK519w0f1FBBVV
WlicZoRZM0hfmGF42yBdPu7lcG9vN+8Q38dIiFKm4yS6AdOUzvTghNeE7Ktc
0kYt3KJ5r/LUSrhTcfa5I2wPPnY29ySrq7Gs2SoXDTaa2+t5H6kQ5hE78L9s
T1f/LVtImMdoM6vrq8RifhXmEQ0frvlgEmUfk3UE/8aDRSHmwNfnc6H6sWzd
4ZlCc5SeSpUNvd6inygMjXEhrMmMxUboGPij5YFfKQSA5BjRYidPKUK1osur
CnuxQfN8FD+3IyKNfmg1X/oim8HhmLohDXp+DwMTcbSFP/rabUT/4yfqIc9u
A1aZHeL94JiGGhOHMKLRdnZBYez7rqKssk971teZoTZmXKEfAlrSoJmNQR0G
nG+yrAvPeuEQEhAYlw/JRKORFHydrKMb9TRI6I5mfiy+YTRM2buDpRdkCKmt
4JeWATFyZOc/Ft/DTXWKc2yIr4q6LcSyXDhOSF6lz2dFYxv7w0szwn5p7jeq
RKHL5H4YRE82aaUIlO6Nq/lFWHp45yr7Q6KY9x7mAouCW7TY8NdI/UCqroIp
2WfMXDzeqtdTq5Qrk9n2t8Nb83zZyMFbkQfjsJg5p4muyBoRo80a6NoONBdH
1YSKEWVaIDVdTPTk9XQImHnW4639tPJ1ya4WcSNE9ytRNCmo6eb8IGah04F8
qWzIZIGfD7wS5UaxuzjMVPlHd1epc3MLJA47jsTC65DeGSTLn7R+8QCW2Gcz
uKtBRn+6b9wId8Y/3bz5oobtA2qQet7TSKdTxQFxmCPnX9Gpk1Wxkex6R0qo
yTSFa1A5pyyeJDNOkNVFsSsMJw0Grw9/JYpVS4D84KAAtshkxoAQaxuhR5JV
V55yNKle34GD0A2k/GVTJI0FUVI3Z3RzExoTZljFIdiAEBwdyQFuaWHqfzH3
nH0/1YfwDwgSJrqWYo5jJe3LPfJURGDIW5044PjHyMH4fjosa0Wg2dx0uOPl
qBQsn5p92ObUfkMHldUdZ1QKZVLOuYqRP+aFRbuyH24UXuxJiHfL0F/M6WE/
xH+lqcKjlDJAwwEaejR9ysSMc8JIEZAoSOsW+EIHbqijxDVTv4izaJi4bkp3
WeqkCjUwvNb+dDbRDns2Bw3R2fzS0ZoovXh79g3ct9uDJoy0V8p+yUh0FEWt
iaaYB5Hx3NdE5EJcpP/bX1eXuZd0n+n3nzQT9HgmHVpzf2fPvNNivLPU4cGt
wGk2PE1BYI72rVLb98VkPQ8utR5W67YjdjFKuFFdul4ncPkHIdtZ+NYbGHl9
E0jGOEdYXEL0pE52CJChLu4IQhw5lw69iffR8n97oxGOfjB4mkkB7wG2T6+/
eKhzoHr6wunW84r/c2N1oqWqIskXeG9q68txvi4ojjuBrBL1UGprvinl5VdW
kb88WYa2fFuim8BUh0ZZa3JMSBqesElkwFZtpP2ZVKZnZnKL7fKyV2s/ghbV
ceQl1Y3jxWfR29xzqCkIkWtbatVbGumYxIBOeVhqfQZSHkvetOd+n8vCaQkr
Ea7V4LpYC0r95eAu5Bjygt7nEcP8nTdpruo65xbndGtu3YgUWbKxr6/QQBFk
RxZXuVKGGa24UiYKDqLcmOcPutrdGkU/5Z9a7JwMGHwee/2CT4jSh55ezQE5
5UoKElFs5zRjVQ5GYFblOVLN3cSacAsJyxJ/DjQkMLq/+tWzp+OGGiApo71/
fHgZWak5/bOU9xl0XVcG93KqscM4ECgspfl2DfGJNfgdqR3mxajj/nltsvcy
VKi/dCK9opEJ8n5CXmDQ2EDBngdkmNaSQUbhpaTfR6FNnHXF7XoCdnYzskHc
2sAnK0R5aVt3v+KbvpcvmVLs2K2QILq/SnwIpqJHvuWG7BRIsE172G529PIN
zssl2E7xBOSlQAKGEg0kP2xKieiDosuirnX0M1VwSGkN89fNyYjwyaoG033r
6DSj+LCFRvTLKXk82Che/TW90swua4y+3OkJJE6SUtBavhB1Tog67NfwU5hv
D0i/Ns/o+m6O3vj+lFIZAPEOi8+zVD7GXPwRqpQQlp2HQMFphHsJB3d+4kOa
mVXxtM9iFm3aqonT6M+92AtNZ77XRNEiTI9OL0DTOredZN7jfUN+3ex7wTLq
wHf80GAxQxS2OeAcg2zAJbur8W1ljpF1D+l2CaC4rgn/RFXHrbFTJtFYPUw5
ae7c55wYHfFe8yfE8OaVj7cYEHWghV8pRlYadtXL8846JhHInsN9mDB2dpmf
AAdVRvqWxtDsDxTag7DROp5O4qBWSso1sQ9FTKSp406Bns39tVn5rLbe7Nhg
e8BwMFwfvMCC+b7tgMMOZUPnXRAhmXN1I3FLfPJDMBDOLvmgJEaZle7iao84
ikYMg5TV8PvAZ8JbqsHIxaJa7yVTlDPnm907Y4PPpuxCE0dXyVtMzQHI5zXf
PGr/hL4zaVDh3prl20YlL51cH+1LiVj4TwVIiGEXAqkMUx2gJJmfXRxbzkKz
y5NhieBSuqOP+WpF2h0/THvJQm/IZZ5hateZ9fM+V0BKYgQjIQnRWLNmAxEy
RNIXWhduc5F70Uc2iF7HzCbdI7Eoz+kwaNShGm7FMZrigg0slIsoreTkktao
MYonwdbqK6AtoBPkFzCXt+8GCPW7ZCDX4pbDkZ2N0BVlfU6H461hIIJFzzNP
7UuGBav/go0jeneso+3xDPztLYGy/6z07h6Mp9kAjcjFhjaCXmxTwMKRQL01
DC5fHotQJ6ZKuH34gvUpvZivYdCBS4tVYY7Y42+JMio1LxEzkm+MAKgHS2ub
TAR2ZMJt5NW5n31Tuf9JypbhU4tE28SLlKWZaLnzznph+z9zjrnWe2Z/cjIH
qUpatEIzJBpYvLiaTlwDXiaVUhuUAASDQMwmEaatz4TcE4Gafh0ftO8UL+/c
AuH1rx3QZQn+2JepNIjNSu9T3DM1ws5x47brKpB5d1O4o1ZT33znRwUNY3Gl
DHm2ErVf2roEpAlIndnpNDCJ9vcGnFwxmKzE1VbYZf+d8B/YqmiMs4JTqu/3
CgyWQjqTiMEhcgRfPQ2Mnas1f69uBA34FpmxximlO2O7k9ka4FTIsX+8TXBc
mvxlcrOXgXwY/Ht1bG1IgPq6fZH3QK/fhccTaXK4uM+hG47i98Ss/nMjWUvy
XLTV6GpKpQEoH4QtpWd0IguNAWHm04a6knPCbrSey3Ik2c9NKztN+8PX0oHv
EAIKEx1EhyMdMZ35n2ubvYAiwHHzPBFJDOVqvfogc7dQSAgzkiycoKwbTv+r
ibZtRKqO3ycBLkAo1bBLgMJZ8gtjs/GYUTcf4eW11jKrIyiMwVSMss7HkAHv
RxjCzZVfnAtwURv5Qd4L6yqNjxyTwWGz+5Gnupl9jSb1+ggX5y7EBBL3RGBe
TGpXWmH2vt3IQkqiSg3ZDiT4ZxtAFb0iK9sAxaAqbB0+KIoZH6gd1eueko6s
r9DCFcU35h972z4PzdAiLqKLFa/ZVmjLdJ1QW2pKgl+yx58YzwxpdUNAHO+E
FlVvIt8kzgsBYwuvO4cIR4T4VTsgRUgRBJLsW0sHnS4qkZ69X7JhDFQAGomb
ZB7Bh6fYczf6R+qQvNOIi+y+yccOykXPMMTnFkB7NyjVYA6bCb0UhP0+jPTD
KEtoq0zDF1zVVbMF0QR5XdusBHfq1YlF6ffu9FLymQsIxqBskg2h2A+3l4UV
U5LNHaFkjDnjy3p91DBovgBd5M7M/Mj//KyZH3CrZHMpvIZcCOSzt8xFYGjT
88U1qGRBHaFS442ANtltCGiaTSCVssjAsRiS7M9WefBj4wX3Ae1TqUXTGK+i
XHtpLbHb/UK+maIjYANPviAHSr8IjXzh+wP9vkQZGfhDmZV33tkcFi8LttZL
uvzLBbui7LlWrqs4jpVq9wUqC2JJ8kbqBIzIqEFoNT8/w8POkAhCceBREVxw
fP2HZrrmXD+yiWjptAcaxfLzH/9v3dphRRDgcd/dt4rWc35/pqhhkmh9V1mS
VLlzZakPgoxstd/HlWKff3VIKb5G4wQewiUVck/xU0lfvLyBVVknwBZZt66h
cZZlWFg1FLdOr6PVu0nlHc/yS+UzrLdsZ9Uei/URzWoWQpg3A+pzxuy6t1BE
xN5Y2FDE2Y7Pf8I1pYdO4JnPnLJA580mP+J66VuiPuGQ2hRdO3ozsy48cXLz
6r8EercWo4ynHCyhe8N5h8Sx98EgOw0AThSmOZYSbPuO62yP8gAscgh6oK38
ZFOJ0aPWguCjofVStRLpfVtrB7/gwQgfICcpebi0q7z/2I3oIZZO6rtc92Z/
hnc+75iJPsisPrRr767mnEzm31BBCLv3BS4VQxGR4ajMEoXnt+gwUOej3RsR
pgQjnJgyTvzW7+WHNUhE49/v57srpDjKfVWWhBg4msapfcc6TEE70kCj6Ym3
Yj6K1AyQoeRItQ6uNyra2wQ9rh4NRRPNGur8ok98/a0+Gnsu5TGZREt2mfly
kxT/e38+eWgB8ux6yZckgN3jNRQQ3EdWj2MNPyjHTsxXkLDWsWp33fLYthKe
KrMF795Mgm0mfHESFGtamO+2NHPptnM9hpFuVnn6CKYkwYpfQmhnMd/emiqQ
j5Hs4NB2V9wRQSgEpQA17qC7VpB4lAxXlSJG2nLoFjCh9TcImexgZYXYRpt5
Tci6UN0484x25jTdbiXx6xXlbpHJ8hds2CtEqUAp6pHcr+DcnVUome9UnkCV
Dax02l/9mhi3WGOrQIMR9vpqoil43SDGBB/x/WtAwSj6gLoAzGpac5BX15XB
VGXhKcWHAuUR0irDLlipuvKJnKEGBmndt2ZRXEacJIe0E4UOFj1zcBjgKSsx
p/j3veQOtXJe4FbjD3Ozgmam20TGjBYB5ktvM7jUAqBfQlKV4eaT5jH9yWsR
+q20qkJZMyjuDWXd+a+A98g2oLuINpsVtVaaegaHQhjplAHikRRzPNyGHJzk
OXQzAC7qAf3R6FOLuv2LnlSjRkCjArjmj6KLZb8fftlA7cNUv183Xr8/rvS+
kXXY3MO5S39v6Gjy7LOTkt8gCfnOLZ6iOjc8Qg1TaoNZOQRLtGzbqLHkIj7v
RwmPrqQh7etW05fNEGjLOZhRLOnvbkhmYYH5wnUyX6qjOoxZYp16qP+RYwo9
4EwSy6CunJRl9zmUZCCtm0M6iU8WzQDjicAtaV+nw53hz7FsqoKtxHerhrj9
3jNpQoa1rVI+umVjSiVEJaOsCwdrfI0kIOS2J6aEqpijWAeHLfRG5OnPplU/
7ksAetYorQNTkdf0ge/CXYpvBLDDoaS4cpS+AtbCJSVI1gkbAU84Hfjvbq6T
NLWwrf21VnDCkl8UEe149zShgKVOtXIQ59/wYX94C580qv5pepWWrsFk2mUo
JNfKUdyn+5Zt+ekHDdXCK6arH64U4Mj4+8iCT7+I4XaI9lFnzgKIxgYSGlYl
FFkU50M1QqZZHAyEFiMZI4kUKvFPjAvs8hLbWuwBubhBufReEiPDT1lES7UW
Ddaz6yWu6AljwVh6kFl8zdvl4ZdUjOVngny0RN1lgXTYLGTe19aTwQV4w5sl
C6/H1T/hxHHD7Nqmu0wAZtfXhJUSZqoJMsMS0n0RoJhnS7Px8NStDXLIYh5G
ZmZqpbHbanroohS2lwu5fNdz5b7H5O2Ucf2DoOoZGVYdFiniN+cB1Mg41dxo
g0jHnlpGiCwrzfxUeZ8j5u19An/3ddce+3EkjTYWosrn6erQid6I4o7ydZNI
rWItWVkWGxVC1ddBpN4hDkRaAE1VYQVZDb1/qQu9bvwnGWtdr58+mEVg4VYn
QJxfEkxricyUNljX/s28Q7llt3TI/VKz8+ulAR3if5VnF2dqKHF7jE5QLWZZ
lt3OMG/CtwzVWVFHNm+yua15Qa0/vExLGZ3AG+QwhXXkvjAQhqOeTIiFjaZR
nEN3CwI/fNw2xv3bvAlOoIPcUnZG/ck/4dsSWPqCirkQucpl098cewRt75Jr
m8VrVtqo+9jtzMfE8n5bFb1ilN/zHfIPkpWt6dswT5LprBlhQP+u6i5fjaSw
h3LVWiYrNHqqkWkjxXn24NH62ejQpw/7FmnHcADx2d/7ASUC6SI9Cjj2X2Vo
kZdvq0jD+uDsMat3gdPrqQEGqwg7e3X4dQqsKE0IN96CNEtLFATczFYVGqXx
8xdVmpoFSCg/oKM/kHlKkgw6zfI5K805Pllc/UkPXUBcTvJydhGKhY4lYnxz
3Y29Tbc7B0r+pGDWX+4PhJsH07yA7Y7vfhK3qTMrsL5epbsMO913I0QbpC9Y
ZpXukyGKmjDQeZfRGFTNIJsfBm1U9wG2dsi/ThMFMBt+j8YkEZVIKyTS99up
flCtAtssH8F3mCw0XzDMJa7ATRCNvp/3JJB0MvhKa3SowdA1jUqTvIWiatwx
yV83Go/HY3ci/vJGeoaz1zoLE0RG/52hz5dT1bbZyh8XE9ulGP9FUdG09Nzu
f1P22nDLl/AumMw/Vk0/sd8IKfviE1X55UYLta6C+SPWOlFCl/ZRt4gPXreg
Nc44ZBhAa76OAjKmTSQCzHfBBXU0yaxzJ3WYN79pPWif55LICytzsB53VtTN
Y3RUyEgkfhX0q0l1u5bMNfYcWNVcNAm/usw1P/upDP5/zax+XCmpavRwMLN7
lIJucJreZ+rhxGg6iSXwVlJ9VraZ80HMyioYgjybZxu5Q8qo1ooHDn+vImk6
u6WrSjCGhLOAtKH8mKdBUrgh7aPqUE9b0COZVV7nwhuoxdqmC1fPqF2ToZc8
kEpA3X3TimcCeUiW5Hx5diE91WpCgkY0fNPkNPGs8bJC8kUUcwNaGvheDRUY
8uGBsPquluJqhb7bQWfL2JyRiOACTIzhDDcylhgTMHyr9eIJQOGhpENsA9uj
AcqdVhuIMh0Ebb8E5rPkMspVFCIr6QKize/m1W5BbHYTmIZ1bn2fc5yEJeEH
CvwvDQCrNAT7IRvkFzOLviym3vhyJZRQ6xaHLEXN200Kn5jFVe8XM8KCsgeO
RQfKusvbflKzlg3ONGU+7l/GlZkOcw/yNZ6e6Es4TK7LTjRCvGrnImVlRlvE
0fcsFvReCHt3QGixFjfrAw2IGmZbjpdgqk/Z6gf6O1jS06fdtBKgWMiuqSXy
5csrxJ2M/WSOK8zAgjAsyTgQZfIeoD6pUIcxnjcyiGrvF/zWDqszo5H9g+Ly
ULN2j/RAdYjTvlQF2bFGzYChrkSroYPvwfEWEGgkIDfURjyOC6IAuTlEvw1e
VO2FxEn1JN5EkBr49G7NY/AdkJ0OUbVC0CuQl0C/ZfQ/Hz0rZK75+sID2x8V
j++fb8HMdUpmx6rb21hjD2a6kk26o6HfDBNwpTlvMowALYwUla2MdqWy4Url
Z5L3ypWn+3+OHGMFueZ/QJqRfxgdDC1g8OuhtqX91ULS5vDCgTu1L5pbmNhQ
Wdn92RxW1C0kd0+fBioBXpmTCIeilgsf+QxOFZGC6r78jjdfFhqSowdyXmlt
DZkCgLw+bllK1Z0wGgbFJmoFmuncuzVhG48B2uQaT7hEWCk7Tq1vFsf7i9E1
Ut1TfbRa1ffioH4DPyNkjhzJIITHfsnwlzj0+MPbezU6sPHo7D74B/rIVvGX
nk8/RbVqGNS45p5xmSj9x/gGU77xyZL9yjGKJA9dk1xs2XEvYeWeaWuMAo+0
3ds6P5dr7C3XJQIl/8Mf0MRwmg5hqYXCuNgQZMyCNjzykoYjffpLxqUXbwjH
tTtlSvigbPWrD6XssKIJeZKbLrAE2M+cSAmLqoSm6bMHWvbxOBmX8hHFkNuJ
dRK4BkfxOLBVuJ7Q5Q/vapdgPvLXdJbfuyZPOvW/2gJwP1e2Y+DfSb6Tg5qe
gRgy6D+MFIcMbCFWViNBl2eKNnz9e3wlFUhxzJ+0Y05fHdhUSmRvqkI5wYuN
NakTT/b2WZpxXGZxDhEwtxIkjK60i4MdDY6+dps4vWrdMlIv2cN8GpT33wQC
trUlNVcqHJ1IsnWxAZjm2/vh4Gl9KGmdpUC9mSRGDR4JPHjn5b7WrCOaYzJ7
oejp9/fG+Xw9OQ7JjFw99WNtg8sSTw+ZxzxRe40WVVhd0TSCy/oPt4IPA2qY
Z7nRcP3KkaCyIPDP8LP8bLRpstEcPL12ev4Al110Y3d7glT1Lvgam1dNjnGF
scIYRmDbl89d+klrZYBnj7SVKtK8ZsoVkItcbibyHuksM6uFmtUK7QEjHzJv
gioFDT3WD65nfI/gW0yWpVs5+3G07ArpJ/VJuTvtOZiD8Vm3Nk72bCKJo474
gg/LzDpd+jam1zLnIQ64jGcdvKgMeroTVpDNIsM9Jsj6d2X2q9x99pjlvFzQ
uSuEzNrnOe8fmlD7iUTDK2NTbHHKQwKnHtfJzSublBSmrVl3RdAjKLE6tpy5
/zRriLYly/aoa6jl0/30qWktKaB3RXAgpS3DeIqw2TO0A0AUnN4pVVTV9mc2
2Yzbgtb9cL3QT9/dAefbS2wnfmsoD2jaG9ZC1PZ19LFXdUEpLvFJJAOlG5GN
vEkrzBoRali42fjvnz7lOaNkxGZ0T3lhEjSQkQxfboJZd3EvlehNg2IPk5ZI
ovcwMGzQ5PROBz9G7cdrqP2pt5FRnuyZmo8f85cLpR+E9dDqq9CpBH7B5WrV
x9lpzMDn34J2vF7sieoYdsqncpQK7Zk6MU3dbIJ9minceMieHrrtSz5U8l14
Cjv24eJCZnVdBR9o+4x3eb+bL3z/BdYf8GSbGurQsTAoAer33wLNfI896mh+
aEuYCeHMcWgmNrhbaFM4LSdOk6iTBQ+VjVdLSz6cR0ICLNYaY4VBPNLTe2mB
IUayHAAV/jYDdote7W5SC98f78ggiU4j6/kHLkTC7HZMpJpBB2vD+JV8XKiQ
9QLAOMlAOsJ9N9bIpUYDvutcwtLdrXCezrv1+rpn1WfiDtbzGigKsd0MF35h
axkxIIRIWGk4s8xdKTrGLMo8FvJt348zaAu+KebQRwZadyVV3fKS2fFcU6BB
YXgK1fip6IIreaxt4TCEZzemDgmEIdVm3t1O0AWiwfYnh3ov1FCfNxB+Hs5x
18PeMwlWazaKg+e9mLMuy2B5vzJvu5Abg5uyhQTia6C/yRBbn/ur5QQqTewK
nxzdK1PvEq1xM0PDatyzMECGQlCT4igZYKMvhpsMjXfFhtXiHT0y9BioLG9d
K4nKXm5H2gzyeanRo2VJqPrwdwEwT0btrHSw8cFRjzYnfLi+VqrMPfXlbQJr
4h921gzNX9qyEx1bEyho9ylHyvPMJ7dBHmyqAaazyyc5jDT31g1TIY4dmipx
mBzOh0Pvp8j6v66Pa0N+WDKSvG3qv3FkVFbzs1ZzBnFMDylMU+UVqpKPVkRB
4rCmV4II7zagrrqaygX3AVLkAwF+sW9KAMrWG/SDjy4DWr9DwPlEGX30GpJP
MWjnNihKVBb/dl7ulg+TdYQZ46hTClSnNiXFcV8a9M0ow1c/SKnEb6hLalWy
dZUrL8fg0jxcyfIvc6oBbOOsc/RfZk7FRHW4ZB/x9UrGOxXYJe91VJMytK2u
GHgS5VTIeHz2G+tPHDBJ0Dd9tDXFb3Qwx0IFLPGNS7eS5MCXnlLvfB8rOFAA
eRdrotqndHLkLKRJOwUs/xPv0a1tYNpo/aa8FFO1u0E5kZJEO4BaqpTJbYm/
hgpYr7UF3H5YBHIi92EVzALTUJZ0Sw5V85q9odtgbrInIGX37tltcnz4b1CK
FtRjeRF9Adup6vJCz9GmwhbuJk+jLh+OL8hZV8eG97I4ymlvhqhCltM1Y0Eb
wyd3ANkOfUJuRibW3UkLZGpNfYlfaOetPW9fe/PkJhc3KRoAFcLFobD5O44o
PsgWp64tc4sV3J99D9vZttFhpVnqiAlydpC2vlUHtit5DLbKYyXeXz65qHLD
F4urkcN5gMFVvD8CdpkDWdQUkQOksQ8oYOxapIinVGLL4sofGDQeU1N2fRKT
1SVP/8J8jCdMDbYXXm7ChrQfhEqPxUZC7x50wTlGefAQpSE5DzSmpKNER1NH
9z0RkJtv0ZTGBff/Fxi5B4O17ZPVebL6smT6BCHQVhgvL3vrFubFVHjQ7I5O
QDQVqxuJkqhUhepAgZ58ulWGlVmlTZlA7XWs55zn+WLRKqQlbdzt9JhXbtrF
PzxcwvySKDq+PT89WqPiUOfMmYvE83lHray/CQrv1ogKDguZZ6uXvwEs75Rk
wEZusT8yDuEzv4xB7bLFxBCf2J474Vj6My4MSHjYOxFSIJPS69FLDyRwHDUD
F5JHWDpE025Hgh4cDrh1DmG3qOerKeXxCGb084HBRc7RMbepdRWmOwVwL8Fo
pdAWjiGcBrajpRWySE4UcFedGsRuTGJUx6sGw8VOdy3lhbqy2fGlpc2tKxXN
Vh1tIPEBX1NA39uHEnDh+QPyagkWB4K+3DSBNQ6Lm+OdDZBHq6pinOO0kQ1G
8mBy9FQhQ5rRNKkAHUaitQT/vIU2jpXpOLph26hQNKcECR9ZLaEyMxQrMprT
tue8zFzA5lHn7w61jdLTVSVeccIz5zWxKJcLr3un3QzrcLomXrcyFmCivab/
Aia9pTPy/c6IRELQA3cvPfwy8qteon873+o3jGBcMM9yt80uXXSOEEpGdvnr
bpNCOC+BXlMG3S1o/uvPh0Pt4YqUd4KSRhu6o10xH2BBsXFqK6RA7aUkLzKn
BGMip4vTfPc4vnwsCeVhWnP9S4emQj09CNSg3V9OldiOr+PlwnUJ0gqkdUfm
4my9M9wB0UspuUVpATIlzEXI0C+0p9iqi5RDojIK1Jpl5v/teQN0Q2Nqw3MT
NLQux49hXJgART8RUrj9ddeU359zm8Rgm2w0LVYB7nq+UcDiOzfdLx3xUGoZ
C4IlJUBMW5//CPZH8y8Xyh5axd6/ZsqfiVam1Bq6ErkT0S139eu0r3LqLkgp
hhP64HccWKbNpr709b+6bSzE0QPHYr6jvorPzUyV/dwWr/4kxKh4EK0JIYee
3a8xguIYIFyIWPGpl+CH7V3PXsWydNpXxkPYyZOgMtm/pvFxgsDEmm7OsxVw
Ratl6WCvYZAKb7KoXitextxRnp2gEvKZDlDtf2ySHAIpV1EhORG5soWI+EUm
ABeK9HgKb8JDQmuPQOdvbJG2+eJRMr5YcG5xiRELjBFRKcjJm265utN0EYHS
AONbEVT+HuFiwjLW9RRLavk7Qg68PeZyoihFkRSqaI/HGPe43ixIIdxTGPhq
HLqaLj28XBYrpypBJTHJ4QibL/0jKKCQ6GBOdFFZOjseESONLtc9aLRZxsxl
WlF2296P8Jf95rLnxD6qakHakfHkYqpKO7zuSc429SrvgyZ+y7GNWM8NReOu
wViORYfa4e7ta3lhn7aTKSbEwvoEkeLke7HAxOUDP7Nwq+uxgG0T4RpYlCt4
YRwrz29awrT5j1QT3ywKlcAlXQGV8lN50Jlmthi2LcRzGhar+3WKL7oGDWMF
xIKBGCBpMknfLOtoMMS6tuMJ8UqfTRzFnm70jmi3yCyxxgg4enOEQOv6Kn53
XWaWAz8k3BGs4WrDlZli0ezPcA66Cq/3QNd66QUap60r+ICQesnjXD8P+TV3
yPOrabAaTM2OgjMXHWuIiVCqs6LU/jEhitMSCnQTAtI8GeaTleXJmzZECMXg
QFKd6ydc4jYrGTXpI0ZpYwOsDvxj8cUZJGMY2fBRANa+GNMWXcz27yXWtTJB
VWyljshNGkiURCsSeEFeYKBPZSjtt5RW4ilFiwoyB/nUe5y0bXYX8+/ZtFUD
nqa8hcqP6QR5kbG59TeK1tAAhZcp18z31naRmxCNoqhYkxEa5AntxMusB96h
KiwK3uksjpZdTQ40s1vMSDs36w9yTkqc/8L3sgK+etYlxloh6krxGQFhagr4
nZsVQ19zXGwfRtfklWGxk7aze9nRhRq7C8BegWFwQIPdnoW7sBraHuLrc1sa
wdaKSZyLols85RW1tNNkhhg/3sVXp+F9OQp45zMRfNJxJQAciBJrmfsc2/Hi
4Wm0n8Q5x1kq9m4FdAh0sbYkydAsNDONzoQrCjH0jC0ChP+5LkgZhIUMB1Qd
BBrzm49mosOsPFzNVE7MEgc7ZlSEXASRLIvEbujWfJ9CJGhZcut2Gn1QBXyJ
pbKVF9dAdTmvSuo2XcT+kyLBHijjB+dj2n200EIU+fIlgABYDhQeZEO4d3mW
bam/AXfUI1QWJ0ENyYVHYnuVvfDeYu4TSB0wPs+fehmNFvlMOVg7NXdLPM05
DqgxMAET3ygNeOpmWLFwCdl/lh0NF37hus9KcS2itlSlkAgxxbKxIfrark1C
o4XdRyGu9ajI0VJ4dXp0AvsQ5NToF9HkHqepTBPKWJB7OKrF36SDE6+ck7p3
56SXXHmU78JBwSXmS6wACr5+u5mxznkCwjkFzKV+tsWqbM7lhk4u4YDrv8QZ
L5MxTu3+I3sWp2VkXblpFEX/g/hmhu/EC7GctlQnHM3Nlz6tl3ZGr0ITOurt
MiZuiz2udV70HxkQ0QU9hIlEXuoMumBRZsU6LoMxri+4zbK3k6mlX5gbl737
p12mvLgDRpP9/DuwDmS3P4uXvE/rrrJr5nYJGUp33Ogk8GRgC0dj/91O7frH
/m7fjsQONYp5NWtcxD5DozLIz9txnouMQ0uq3LUmhUzPqf+VGNGOD/MbQ8SQ
NaYqTdCKKXaFGPY8wShAy0Yb0jRNsnVS0O7qgw9nQIVDKle0fDrpyq79NuD3
xxw8Hqecuj8W3L3hK5CwDbSXPVgNID6erwEeLan8/UuQrqA7XAVetBCoFGLB
SPsYsImxvbBgMwxac5m1CYpMXEDuJVO4h7pEHi5B16JQqjQv8qUyutDpxzyG
xAOfqjO5tSHsJazygxDOadtntrV85hBdH31yHsl5F7ioq81yInryNDgdt4XR
5EESmDVijlYHiaBxQo4LvYPAZVNycdPQtNGfCZqBdwH65jC0Ss2YT/5FgO42
L+UTi8RPwXnOBcef7RHyKJ54RL9RJrGtulZEfF0EZpnXLVujlJcVgWYE1RIK
Qj+HBDosoiGlnRu7LAtWdTN34yfagyg1CENm0RT/oO5mHNZ8qfcKvgtskvSK
jT4my50FbtdT7PXdf41KRIspnV+RpKtvoa406xi5fVGkd3CmZh3BZ06hVIta
rGMw4rInUbjumHk+iqB6G3wyJVd7C5JkdX2h37QSzYQQF6kZH+leP5wr/dvV
5IVfCjIMHY20R9a6u3/gs+5wEpUrSE3/eTdhq0tdBCKhzBWIbgov2Bupi1Ou
0kwhO7XK6ccrC8gj3aVIwQvHGlQvLcdFRhdCdJozjw+UV/mg+x6ksWwyJB0c
bIWaLOkFvCMCGSrpmWWz0uidF03O9/MQDpNopZglxEFHUVDSvWuGedid4cnW
Ih4gwvFKjaISf7V8V86g/icIXjOcZ4pMFnmZR8rzcdaatElI7xkgxsoj63P1
/IT5N2/Cp3bFSMdSFYlfIE0jElHzpAWmlBeqrzPtHYhg79qJmyqmnaZgHqfu
riOfbF+8f3s4qrulFQ4W1sai+5ayiWfQCbqysRObu94idkM37J1fEKHB/6aL
xYjYYQndJpV6IUAwdQC2HKZ3KjGFB7oIkRCXkTu2KDleBlcdRLzFYrUpDzf6
PGqWnFdMcS8fg5kzF10fC1cIC//t4UKfvFQendGsT1Afn5b4/Wjyr9XIWORE
6/Ph/7ZkxeHvjLj/VqN8EfhRS/0MmRUBolRQ+GgCBrdBheC9btVtf6xy7J+G
zj5S2DlERZB2/OS6CO8A6JYKcNeq4QqPah8YDsT+kYxF+02NPM4epllAdEIX
2eoecoi3+YfsxjYFH5oT/GDF/lYA10RdCVGuqGv/3GRd5QkxkExQgJ1JZAnr
hPYLY2e0iaLQph4czRDLjJDGrCyk1hNG8nI16oFVn4/boQadpFDBTtVo9OIv
u8CsbH+wm1XCl8bg1cpOOGMBMJkfLx8C5mZmo1Fmb+coT6ydbd2wQ7g2XuJY
EXu1vhG34zSYt+T5U/nZX/gplTbHTWqdlmw3M0pFW19tpUihZTas7ubxeRqP
wW/fCNWK/uti6eIEl/QBm+W+RDDgwhAnSuEte7Pboy1CcqgKVEn+DzRlFq9r
x4JkVFiPNHGeJUczMZkPVQtgGl9N0JtpilEouP6rDtvpASqAxBFHrdXVv4aS
oWltN6ojBOdXzRtbsEmjfkSIi6ECm0bMYjGy7AcVcF/IlGKyoAWKLgkM1PKG
4A23hy24bXB4EZ+wp5ZElZ5t6GpuQxIpP0whMXoy2yGwn2d6b0x5OZqNaR1u
9SDI0cxpkJ/bUvOjNfKc+0JSG66xT8R4Yfg6kYhm/acIkYyDtvuKfbTjhoO8
Vu2rJeAzU8Z0eoJJQBEHmu3HgvrQ06b+JxnjFM6lFcRhSYgtfekVSa4nHLgK
X3RLsV2aFT8rL3VHnXbjE0nCh7xg0EtX5uAFXaklo4Ila+OWlQ/NqECGafPQ
5qACqQcPXi2l0pYrcCTJjaKK0unH7e30Ob0m911NEfYEQeuhBtlB+qb6zDrK
L80T/4LmAPLywzVrlbA6zr4wJbo1KxpbpDRQlPiL4FBFl17TboxDYhDZG/G/
3H8JnwIaF0nD9j4NY8q0aAY2dtgceVy7d5g8EchwDomZPttx8/A8jEEtEI1E
4uMgOKL2hxd7MvDt8BvLBzSU9h5omBuTAy1WuuYt7VUJJMwsWjsb8N+roW5j
Rppvkkdri/Mti8sexITRW6BjYVRnSkPQdr/0nzqsYWinAYMz/fiSqK+SbXaY
83quS3+iESsWSZ+7lcDW0tSbRN1UDFeUMtFqO6jrDlYogzqpFACEpzHjVIRp
rE8FC1LVI2SmHWLJJcKFzY9vNMnbRU8WHRPRcWaGdjvCHS5OX89m8inxM17u
NQFaAk5RMSmpYrJplQMIF8WBmqvdMSqFFoq+wGSKNxgTLyxA4KEQPD0HX5hX
w00JYgmepVQZBmCXDK/0r02PMLVwVp/YvqeusrQbKLJdtiTJ/0R7jey+c+FO
VppXfLHocFX6HydcN8mcfo6omKwVTDr7wM+za7kmtgjdboUjE/cj9qsEpzBA
KdQiamEJBHpfueTA8LTUTlUmOvpWvNqX71MCPl2Bb01geG4CqlLucftzl42G
PrxrE0sqxy/iS6yBGgw/+RDTS+G9hCWEo0eEmyFYKcgZQgvkNFMqb+v5tqU/
Wxq4I4hT/MTd9XuxNubR4RvsRjCVg98SdjIWIlozYCf65XZTA3Z8Ucmt5N6X
dXGH97gHyL98P1BytscFDGCO3qQ13bSaK9biqFVx9kcM7s2gd9k9HcjwFA4w
WnQyoKmiI9qOFjXQLlVhQ1vuY96JofUUNlpQ0yY6gFXpZ9SAn2/olGHUgV+o
zm/JClZzTuNcmueYBzVdYeqRAF8e0cpUaOskPAUiXrtyc50SE+69+a34ZFUy
bVKFxpktwxi/BidP/hiBT488I6DTefGLwX4T+0sech8Q5Ale7oZ7DXrj/pzl
DKvetVZvWjKvjDTbEKEEmWf18ITYDbHbqXdlBnOJ4YqFYO0I8CfyJHPgjA7Y
9e2GOLFN6xbjnUTrXRy6/6RTTqty5le0iYH+9kMfz+XEsnqiLw+7fCCM6MV7
vEMIAK6vdVNOihtHyohrfVFxSVBQyL5RsgTkqpvBCogJEKu49RlX0maXN0bd
6g2zHpwWb69uV+rnejWOwyWZ1Y3Sxt+vYJSpLoTNH7JqCLp9dHd5/fDqWkRy
b/QsjqRoea8nsUezBTfDeyZD+kA4xwQpqYHy09ZDkQozSS4fPwK6Ygy2Litw
v0/gg+SqFbQhmvWNWxAutgQeP8lKy+N233Y1e6gZnOVpQAvXUflrfoylwrfU
1mu3XdlvFtH+uk87xOnaftajcGvefzNqmfsIxPGg6so7fO4l480hZfsaLmFu
V7Qu73pGrGqDxepG36nA1Xq8e0uwcjs2rVvN7LIwz13YW/0Y2oRGMX1t0NJd
htboCywvnKRI2kNzfuDV2YX9203On5ZQi1O30n1HbQY3EGXMyY4uFnwryLfD
KSayuPqwApIc2svNNUnPjthef5EhdLVNptfKQE+Vtzweu/VRSentJKwGEaqW
Kh1bGeFjPIEiMiy27NaNcYUiFgG8lIWBQP/WryeHMCO+8U0n5E4aZTLp+UGV
TerLV85OzzSu8H9MDJ0kv7N64yTGQXAidHGuHbSVWjVIQIJ84l1jran7igce
PWg/bTdNOLjYiPaOeR7rlrBTQjGQh9fYT0UV0Iv9ZkmZDXrOc3LJkzUIc0HA
F/E+2BlrPGQAYn0+xjIjSJEM+6eStHXcDNKNaFg4Q87a9yycfMfzBG8A8Nhc
gl/PcoaGR1b/aFjeKvTJ89ny53Fts+OQlgX67aQPKxzpdoEFgFRddWJ2xnUM
hjXZZ7vihc4PtoKx1hBzEnZl/VAT+vlLm5vGPykuDMlA96BV5fVNBllSB+q3
L5p58WuXTGXyfEPX3idpBgebpAelEE0QBvVwJYUCvJQ/nmtAV6ekR690eTki
klRZLd+mYZ/hFjmciIMRFOkC92DD2axNq5ecWwwE4KtXufLpzIs8sLPI1luC
uOe6BofautRycEIe0w9y7SFj2fXW7Gra1TqpZSYj6YZhu7yVaJ/uP7nk5sTV
x0NJCBO/xbr4mRYMySp6lsQOLu829vtKHWqtT1gt3dYSRbfrs+8Rwng6FBY9
xfIlHIGLPuGYRWrIkh+PxHbHiYT5xxzgOh9KoyHOXP+ujvk+7W9RbavZE/uz
Zy41WzKZipXXSfCqcbNwBWTiA0hVJXxvi1/S5/wNRRKbinPwnCh8ka9QQQD/
jWmB2egd/02AMfvOg5QAAxGl0+8bcUPMKC+F3C1ITKlUYhROsRalip87326e
2pD1m/OyzYlPvwo9Er+ryOaPdSG29zNTRHI1+nGpGqfE83+Vfu9kMNvOZTqp
SHgWDTVz2+ZPxtcWs/p23kQtfw+sgfH20jhXugGiYTuOrM8Qy0uVLkbvRWfB
UW3J71PpTUfCrLmVs2juvxotAAAcYpKuKqG+6/WgJaYTXoFp0xLpLgwxelJd
YqVv10zK4Pp+qZqQgOazM+suInnC/7FD1l1bp6o6KONu33maQTeFo4vcboT6
M45Pngh8HClHLseRa52C16Y0x69ETaVwyFXVNzFnMdfXyCODSbish07yBsxb
UzTI2yU8yp8SUwjU2kQiKv0Mh6CBa75+IqbZ4OToRbZNO2WSiAHDn+7D4Pzs
1Mq8Isp7uMXueUHetbG71nqyrTzudbLQMxHXcqUqlosDE7q+PWSuZwFhNrG0
ETngVQhbsGgNSUbZq5EYXjayjK2m1xBgsjWMXH+DuynEzDvOKIPNezgjVk6q
yr/SiBHQQkctSpo6rDnG1lDV+G/tLupVulmlNnudF+MeadCnvvmaQl6nJwSY
KaXySpexFK7kR3dVfDjmOTz5b+N19x/l1f2aLcsRnYI8AV7gxsd+4oVNBQ0g
0vcrxgzM1W/Sy2Q261Zi7P0u2IOQIwDIWcMbGS9YDKay1LtXdbOVsXJNe/y2
NuOH9RgbAJZ+6kvOZ852jM1v+3PxCWhDIth2WuAShW3BdOIhYcL5Zw3nSuDE
+O9iE83ODzRelok4IJ8NFxlEweNb+0Nt+V7R5uNrbdvYtETnRmlW+eqlddkH
uV4aidWZh2lWolD6iwzIie4d20HqO5I1EfiTJzvbjDdmSRAgUACsON/NKnhc
Vdr5gwgkdYmUCf0kOswZPWJLpzI3CGM6+SeVXELBMISVEHRk2As8wFhv5XKH
io8BZkoBugg2semY+TATkNnV8wTTwXlRjznHc2NMfoPwhJwLyYlDrNOvczw6
r7onRlQOhPLVpvU/+M1nchRZrL9SEEGpHcFRMEhlAQ7SGx42MW/56vbg+oBy
TOKYCJK4QT16i+Zo01GiqJ3zM2YiXU6COyR34KQDJlV12BHvyEv7W/Op0epa
tEIVMXC6vVFHhJO9oaYsKkcfpTcd51RuckgNkKD5YUn61Uc1iluWrO8Cks9P
emrMSq3235c9aANSqjZOKLCo0IVdvgwYhiiW072hZ2PHkL/U7H1rbFXaL9Wn
4gyBncgtZZTWNK6fqhJqtFSKNuA9ZjNXPV+WufuOe3eJws7o+9kTs4FahV86
d4t9uubjKhP2kIa54RcpRDtNfGDWeLNRw+8riHjtc0OV0g2AvRekF39rF82V
dn3q5BhfQoKsmkNTP5OT/Bq/t7/l7BJmcDgyoaTo8sLcYfXxDoO+oKu92rHI
9lIWEsErNyJNbhgLNMrieLQ1GyJYBSSgmZmFLnb7CPFEL6D0cooCnuv/PV5g
wrk2ibz/h4S69nPX4Cpf5cORx34sf2qW9+yxUSNlEEUYeZUOcPf+huYqqjsN
UnxHgG7te0ecfoQxHq7cTChWfolj45bAtxXm5A8XVLms4b/KZqpNxKgpMpF+
tmo0r+loRLHrnRONVHLpJa/uyRG2K0eqCvxCGTk8sDoIei+5RiWnN3pKhtMJ
vHfTNte0zD+2Gs8sruoS9rB/gqbHWEkhctwRBY6zXD2LSZw27urJRUuEbmHz
nP4PtuaKmu1h/YnDithuHdrrj+HqzZz8RImswT7Oi4+qY0ndm4WirDQz30kK
fFKsQAiJLOutHTYaiZR/26ygqhbodc6tp2TMRLLsxlu1d246JvNtNwwRb3Gt
VSv+mH1n3TgTA3SoJNXRgx3L1D4gxn22RD2P6Qpxd32qLzmBmQozB3SGdfTj
Xya+InCGaU7c/JQtIipgtURnHP5FUkrq8yfkbXmx/OmZxiSsvjBAbVeQaGH4
qe3hIlnx6kQgdx4FO+gStsLwwb1KHlBnnrPUNFWI+8MfYJOZNoMo6QEjRX4N
xO/ESBUeosQxIGbo5sgMIsDMiSHXGU0E9dW669ssjT0qIvdrOnyuXHwDRXNe
A1iQ2ywyYogOt/JZ+Nqxai8dbHs2rWsJDXjqrCAUvvcddBZVZHjlU7WIPYyh
3WlHZxuZqKkmBGs5DLtRCCGGISacXcgV4/jlYMahy4/J/RmR58+8Ta5ihpsa
KJH+Fi25t3G+vrEk+QlI0v2sutnPUitbRiwAfg6fnZUJwbqh1W19RBRKlcOF
4gqnkyQE8UOB01OZd2tzsmGly9Qp2KCjTCVY/p9RY5tMDHzSDvKVA1xe4dr9
G3eQYxnPWXBAKt6OFHWeWnuj46LwWygQxvUudegUb1ozUujDl13p3pJZ0FgJ
DAkZy1vZsp1hy3OzzsEtPtcP/5yn4jyVrq8bALnZRKBL2dUYbamytrjtDoog
XTtNDwqdUuGdM07wcaa4+5ewHYL8AfN2c9+OIyiiaDuR0lRwg2z422YBtse9
gb5mksMCGERDueT2lPUI8q/ZleWOsYttjWXbrOZFn2HpHin8fno7tre3r1ii
V9df2AAIF2TEzvHSk+zqp4w2tr/YTc/7Qx3bQIM+iZSh/bAQHoLFwUhb3+Zj
u2P2neN3ATIOzofPbtLJHO3BRX5md0oimrhFM0YrXhJsqSPokKsNueVO3Ft/
/Hswx7XHWHs8G375/nWIVow6sjIyVHBU/RVqUMjtk2g6+zvcep60v0PXQt8G
DXDPh7OAiJ3phx3urv6ILIrTIZKvxNW45kk/j+OhRRs4/TnV4dLxbjbu1hTP
092YXNyJGPet2j4TIgtLzP0zn+S5r/VFGqoARP4eQrPmF+VDc5JwgxNtOBYP
YJZcaW0iVLb0o3r5mA0IRQbs8I87jLVw9dVybhaw2VVbxwsk59LA57gb5CVp
L9/tAdWJMZcZd3koSio7/OdfCKiceuqqXH2VqziRKufHO6DeUehN9TfM6+T+
PYkH2Eg/H4N5o2Lis/qvpFyeHBbeNUJLv9qQvtTplY7Kw4bQtb+G9l24FIh2
utKg3ko7PYCi8MSMaKR2MhETpn1xhSp3E+b0VE4y+9vVWuRL9XE/lLTi6TUg
5vVPZdVwhYJ5ix697Z1zuVpA1oskQh2vSaS0ec04PCLpuriRs3hxhOj/JhlR
fLUMcMwZutMW1jZtX735RrlZ3SECM3fywWZa+osStHbjoqILwuxGrIw0VCq3
Vn1qEIVUHnizVe6gc4PauV6dMFFiNHqNPUSoq+kyMMu+BQ/cRyfPlo+2Srw9
0uN6qzBtpyj3/Xg30X00jI7m+lllj39hasjbp51dJa4cJah9wrBC82KYaNsj
x42rfSe5nIMTMzNyF8H9kreOXH69pr3sOrr6pm5ssVkM5Cx+1MlbZchDfIHS
0KWa3G5HjFh3it6K5BtQ9wN9v6tmaW/ywLl+2Qu8QvyocmxLJzaQ3ZysWMrD
lVVkabXb4NHl2lyJrYlbRQYI55kGxJ4MTwzbW2j6h2Rcd+TB2RBwlcaNMfE+
i0dO2thEqeTDQVkroAA5NKpELUou5gEDwX/qtARxpeIk5sYX9YMYIlCCvJcW
0/8nDHbX5Okqm2/mSZgFTBzckv+HgZWh6GdYHm90wxzO7qYg2HKFy9ycwfUi
q9nlZvWH5sQEid0ZJZ6jiyVkSrbyAKyjwbsntgMdWHop6QikSG5ORyyaptXF
ktByP/42L0RXrBCGuJ4HDLETtIp09ARXc7c7OrYSef3HXxF6dKxSd2n8FfQ5
VdqSSYpSaXjN6svZbH/CXDOP7ZuyQ+Yi0xlDDr+aXipsfqGLgbE3gGAxtzO8
WfxDMs4jdjxaHXCqIdZCNhpvjrrSaVqY5yye7MPMT0hy1yZ2B0afhrgLGws5
Fh5nky9wLnoYMVW4V6FjpmTCapD98ZVfPA9LDhfyS0ZvxXV44hcuQOc02Chv
OCCwIkNMbkG4oUIhdL9KTpPo4nWVFAAmR+r+3Rne/GS2f6FhZDQv4dAp/mkT
TNoxR9s9bQu+Nn+4RKM3kv9pW4NX1NKjpOYIh9UyW2WyO2Pyzi1/V6xCbeCz
Ug0v8J644DWgAOjDFwy2j0nxYovCHOB3nzTKEwcCdZCH5coffKViw8y0Yexi
9DwkHfaCWawRWssB5dFvnQU18KzHCrFoxfW8OoqQCh3W/PJgInn7XjZFUS8M
QoJCX3XDHuRDLOwMtGxSQU0PiMmU3/3KYDKqjjg0TzSUw+WicZX2oTmruVsd
z2imFe1OKJq6go1SBYn5Du1mor1YgY0qM/66gjHGFyZf2TV92AYSFQZlPNAs
jZhSgdzGx6xj0YvBwYPLqOR0q6EDl/MKXY2UMiT6H3zcac0TFrj5LDB8AYn8
smf6KYootBC/j29jigGXwYACr1DEVUP4gjOmD6dzrzQG76d7gLuDjExWyDiQ
EE5NhbOxI8zQBz7mPdTFtLs3zSZTJZPQ3/hBIuUEswPXuDFQNRs6FE293EMJ
CjuWOdaTH0dzziLrs3gVna3n4zhlVuPn/ICMlFw0SfEqrom8mJ/6nFGxD4Cg
RPILPjarfD7yzQ2ynJ7xcvj8sRBaYguKdcSai3PWsaH1jUsrjNj2AH8TOZsQ
aVxEoUUa9bLwyA/tDqqJtYux3NMmfL8lCee+B+Lx5Rvv2cP7+Al8qb8EFvwv
+/hiQbAxPHiMO6bA4v4nZPGcnwV/r4Pqxfqje1oN7W9Md6o8XgoubSACjz9C
0OGMJ5xkYVf0PlYfqmvgR4UhVyx2Gp9QjQxaSnsTHQPH70FdJa4m3qozK8sD
mdiQfVjUqv/3kYPLwWrRrZrsXtdEtIn0b3XC+KgwY4atuup8IcMzRUldoRV+
HD7KfTB0LJ7I+aqGOnCRBjQGiZ19DRiqiuX0HRnsFC+lYlew+7eTUn/jWxor
Z702uhaEJ4dju6UYu+sIvnCbhyhTpcLshvPhVwx9IRBs7Q6rfZqLCQWLfnWB
yVClAcPG+k5o4owqbr4pTt74mfYwRDs8cBRhfKlnEmVKIq2hE9+zrtIWF0J7
eM1bM8337cdNKRakOqNIE9M1DO4KDN/sUCfwt1UP2rkl0Tl4k4Prx2R3y8J3
jIrnOJG8tdtKrtZ/Y8hkoHibUI8QnBxsjIoKQHvCGYr5CcOgTIYR3ImmDjho
iRi7lcUjMVCW5pzjPG0vK4/JtYlXeg79nAtcgqf5M/cYOi84yctqBgfKOyI7
cgrZ3PyEsyR/k50Tt8HVpS8w019pR2eZ6P8NymnI9fGh7BN1Ge5Ue1v5/sMl
Bs36hCsyJb2M2/HvC0UnpSdTCRuYFKGNA/rBKL0uOzS5wPxXUZQzj0lEqUVm
3c3ktJdx/OveE7Ojzlch0GOCL44Ot13M6C5gqCC7iaqa+RxYqjCjYWHHUuyg
OZ0DOMwZwoevElJJmtdEY/010Udvs+MoMNtXIyHhVcUTCxs+ZittDMsuf3nm
FC0KMcpsC59xFZMs0ih7I6+OmJbrk2vwxdWpadTFNcf7om1ckbwNqbKEGdJb
ApgnQla3ObKyYJLU6mQkoKzJKP9XTjY8HrSRW7TkqlNwy30k6q4qiODp30pz
bV/Dgglog/N9tFH3PeULybgmsAkY8pSTk4ASkTFj5fTIREl0z/AzRRw/HHQd
ORqQy7u1P5nGlb2ueyYdEireDpJh/z9deIRXleLMxWRaIAxRFbkrgfYpWxI6
7RgYR14+uptxe9SH43ejldcrz2L1gTe2HTWqccaE+cNTnw5doLKxYXLM6cZ9
yV0nFlhHllOO0o4MMX+iLgvoaR5GtxjmjMJLmYbxd6LKbdPbaK6uVzijJr8D
tvduZr3YJavIwMARKRm2OSchEx6tNjbV+uZxhk3rdhgIA0D4X05uDiApRGBN
XA3XEwCpvx1US71Uik1CU4krm5AzqejUHtojCQ0kYCwmNOVPN7hSyreQm4v4
3MTCApuSNt7bejE/u4WF6DlmsZqL2xYEJHo6qe0JrRkGiqyBnTb7QEzK0ipD
M4fLTNEAfdhkLOhiIstFH2XtMZcqtWIM8vvvubCqkNErlKLQtyx6V3rQ/LDO
i22HklBpFUmOtbkqKj8arwUnmheN/nBA8XWhGyravdjIpz/riQWLrNoDM/1Z
qNDyvlU5P5Vis3ljWBltyDKfV6hqEQPxNu/zWuspYYaD5cF+jzRZoigpuCO+
+8rGq33gxOW0LC3HLmxC47Qq9fJ0adKKuIPBggHory6ad4SRJZcPBpyuZ1ou
y2Kx5R0kcTv33MYw1Poh9ohtwEwhVXG3NjyVOOw6KKglga1+y+2B0ddBk3LK
J2nTr5Qt7jVPqZraWj6my+rbFa9PKqsfVLBZ+yZ7gbK/5mOOI+R9d+CYe03Z
yYhXuuDv2R01pv/4/P92/lZSVNyYbGYeho3ocJ4GqdNIMnNAN3TPRh+tDZC6
5c9U8eE3QvQy0ka4uEpY4WPKg0SDoliV1UV+XBafTgevxOTlh8YfAlE18VSO
vYobf8829QpWKUHgwjOO+qKWtwWh4nuNJWpYyTPqWJHGq60RDHEVrCCXTOgZ
196boR73A4V9wIqQxTI/fv7iquRdgh4jVB9ZO0F6D9f2C6GcWya82S6sRLrA
vqnhDW9gXqWvTCcZKJV5PxW6Y8fWvzuOpBD9mgaUiAS2o1lAoiUW7/Mn/iqK
LAoht05HJAihhRUDYEG6JJZsdP7hpuG7+mzRXb2RlruES3WZvQniworKd3El
tRFnIfxNs2xxMZVDVAeudn1y37R26HW27uQuSN4R1VAEOaRnkkAB3n86v9Zb
npK+KefKM4PTwWsoZC9kVVbYAZ5ZhZcOQel03I7H33gHouRNVyWjvEoGMhwJ
6ucDlG6XMBSci73v3PfHoQgFAeC+SKw5YNClMOyWjliawymSY4BF3Xmd0R97
D8w3MTCO1dXTMdllwnhbqOXAcGsXCtG7GyMZ+uJGYv1H5rcYD3OHND0YN8L2
rkR0VkSMoCvtQQNlCb3A5vFWX0CZlJ9fPL8ZGgKdMbdfKiwpgFUX+zFBCm7c
ZDjL0e8BhgtDAtj029IAqwSfhm4O9nzjaaK6Qv/ioZvEDXkPIk9hiDMYG6kC
nFxsufnAzPDmkfKU9I8BXR2l86aEHb21JsEhtWZuVg4NPXVUC3ZkT3HphYBK
PpyoKRw2QT/usa1yjxyBtndDhxvdkGp+hO5zODtO/m5RKRScY7rFWmAzGnjp
3vzEub84g4GYVcNtqVYNFd6MfaXfDvxx/pfCJE7nPZjWS8kGnSUHLm1tq4CX
KitPJeVWFDoli7qkNTQCuHaAiheSZlc6W0pannznSbld42Rey332PIkDZsya
/QfqG1XXii+z7joQtmCe/LO3CZ+9S7aTnKOXYgy0wYZ0Tk/WU2r+KsbCQ584
NdOEtPnAqBqA8p5mQOEUiH61A5bdivDPGuFGtpIvsXc27z4K6L432WWKiUa+
DjJ/glZ+uDcSORBm9hH73zCiHnRchUOpCKvb0Nwe6M4DqqvObygE9eDgYuuZ
zzs6id8jlZH+jaoAUni3f0JgX0WJBQseEvK59SGeR3hSd2SbBPYPGwBflbXR
UFMKWJ+29UXTAMtVhrX946jn0zvI4k/C0HYIWfzQITCKKtKmHbOZzWlRm9bG
93RnkhlbnX5Y2O5067OHQ4YAFGnKK0tLoZR7jPUsus3WLOJiORXYb8Xqx256
MZYU4R14k/hJvGzCHSB+WVnMXb3U0Iky7Yr+zkCFegD1jOXIcazhkGIcnYRP
0PDtC8UQFP57PTf8GlRAB9YB82ysDhewuuVGTFipQX0ezJeKmdOdCMpzY42V
KkA+Nwk+E/PIlNfjQyOHF3NkYgh9IorIW34skZHuV/Ii77oH8c1xsHlc4Vp6
9V2KyT7SLBROQe3Eid2Ug+1pViQTnlqys24Qdrh4ixpS4r+RmsID14MySJTF
dyhrhVuMNSE941E/uMDpIeL5jVmzNfVlOx3Fl7XOGsHjMSVusQvU57FtnYXk
Zp/qBypd1/F/34KkopYE9AE3zEadMSwqPbuPKK3Ay4gKST1ud3bA58w43l6J
Sowndqt/ipQE9S1r3U7PGFwhgyRnksxHJY3oy928k+xL9LzLRn8fraRuMOFU
kb5DhE19wV8syubbWbO2iKBucaD4C4SQ8q4zBy4vIJTnBcFAfGFv9Cu8xSUs
lFdwivgqWvf7kOHdSnvUC7u52Fe7zxEFOjxP/R9OsyzprLSJAh0Exk1sSyDo
mf+6iF3RA9whyju0d+8NwqrUp8ri3DuRnc3qc86UAXB6tYXVoKGQQAdCws/f
Nk4+kQq+vrNiQkeFez2sacpPcNEzSrguFivz6LlgyYg4sYpWIPYGlrh81xz6
FPeOjb34wdjIHx7I8f3WC1cZzmmJpKywcQCDsnDZJgBL5s/JpkWZXVO9O1O8
Zplibck95K+BjtapeO+yjeoCT7bO6c73lJl4n0sMn8f+ZqDsaZ+piW8c1Ifr
Ywv6wlbqHRPXuUg/NC5ODSJIxZtXZPqmGJ38uK/70cNhSxcL3bxtUCLIlA3s
rBJRP1M9tyDy8fUlPgOAr30Jf3HPbwwJ5GjX8lQSuNXmmfPOUkz4z1z2che5
z8WuDJS71ABlYMm0+7JOpRdVt/bTSlCvy6KXJHdNliA3+67ITClpNCtuHKfQ
3R5O6VZW4OhCpRQ6uvX+M7VSce9f18KCiAe8PFHc8+t1pWGjT7RGinHyXLNf
9DlaCseY0aXDEIwr653as7I3kK/30iZq8/lS//5pHvHbF9Z2gXa2Eg6ztlF1
v64Qa1NgZDDwFcG/o7ckPEOgKnJPEKISSaJQB8dUe/+u/ZqJBoxAs70UBhAc
Gxdgq1kO57zgPu2Kt8W6DlT6ZHQQaLPqtTxcsOH75JX9lIAKlD96TWXMdFJ4
z3CfnwFQ7yp5cIdX8BFN+UOYRoxwhA7Rpo7eXG2L6JW/WPAEu1R8ni0jKr3J
eOJ63FYp6Dsg3rDibq9/9V/JDnNMow/2DUu55a5yMOBFW8oidviXvbW9lFMr
djorpH7AwM3Iy8hIy0qNz2rEoq+kuae/qePxsue3dW2MH6HAm4HF2DNM48OY
XbWr6GQUqetu8+q4n8BqTmCYsCPTAubJFnn8lAcDnU4SFTd03MOeiC3DJuTH
VsssJSE9bTFboKW4+t9K3CnNvGkmR6oRzIqEOM3oCfWHlnw3EFdt4oF/+Q4q
FelyqIw/WuWKRssLaHtRsMoNiOMLVSCqwuKrdo01UzJyeBX1tqY+9y+DrWuM
Qn46B+BpmVnwK58bnfcJmEm7Byq7oT3XcOcvt2UzfVErGaNT0oaJddoo4FgL
NZUU1kVWMl2fRIvT+XIxjBwTAk7kfS/sFArhbf7x35d8CuoUTQiRmLmTKLiV
niHtMAUgKoji1HsCyqY8KMM+qphmFK869rftJuv5/qwZgFI2F1/lx6+ITWsq
Rkh7VQkpUBz7vnzssfWzNM5QL8/4vPQSmyZYJWVKJ610YJdVXSbCwiBSR7cr
QLBGzgdZQFxSr5cGf4HakyIBqtQW3q5w+Q1M+5wjuS5bJ7yOJUTtTFSytJBN
Aisrjipr/ROuqe9EXowJVPsM8yI8rBAOE68483q0nArqsNOM8ku6NHbM0Mk5
JE2lFiUZkScmO+ILpPuErzMPAl1aLBG/UxqR46A8xWMjqA6Wtegq9Ehtbypb
Kjgz7a6d3oztVDwImRGIRERkxsj17BzWP6ievSULxUvSToo9e8eYqm0CpUqT
ZZCGoUkpKEJqvFE+DRUqhRUjXKhKXETCZog7mNQ9Y/mwt+DrGF0GawAjWlip
hWilTl8Uf96uz6yeZtgwe/LDKBU2uZkYKMhIcJy1SoSzKRBHHc1E+b7egqFw
x4TQavdjHjayd7CWuay9uuwjaTeNoJC1jLqZLa3WwtVadeFMLGsXaJosLmHH
a59n190mF1IAePPOFwowZ1jf5BG9sdsrRnt8LLCze/UvisC4kCT9SokAi+3S
KEDZjPP7oUb8n+VpNVeGSy/L4lePToc1z7b8M9qRYHICdXTxFX04iHz9Hej6
aN/hCqLu7JUJVMAGFZ7uV+urP0vlpnBiTBNCN+c1lJw6umf3WNSZvLaAAUxz
99d0HnYKXnkEDvP3R1weLgghigFr95GBE0DmeZ/sKuTZMy0hM/3dvLfiB9HL
OB0Nku1OylIozQAIBA/6r6QI9Lt3NWZ9zdWs0liwN76bM/1jxLYdhe5pFC81
CIdyUGRaBdWCuKpLiClmwFvZvK+beezxiQa0Nnaxg9DW8t5trd+3kNkJwSqT
PGtAPECUYtkSEdATSUeP5sN3lQxjYTfbOMH+7TVvPy8A8vbJwRToTwpWKcaT
/8wUry3061aZm0bsBqh/Sk6iXsEfvWZjd9J+1cYV5Hdm6Brl8ponWa3JnPgQ
xfjWzX49xtrxgeFnXaZGP1r8/NppRuwfL2Hte50Wp6Z8QVjJJw3pcMe1Mp3v
HUlyeW2AR1b5f5m9kX8q+ADgjjOPSyLXQawDvv+mWf3WZ/PMMUY+6O/x3VG3
3Fu3hIwHoZ6lI5WgklZhrbhe/q9NGxLEQjewQ8CQUzlUlGTpsfDbzJwT82Zz
XxbKg2yijCrpA1dhhnb+HLl/YXLLLJIe/pVvlVmd1qFJJVzHjfsfZMpnOBXK
3yAjfy0VmXgKcsQjZ0YQg1S7Fnjoa+eSxn0N5DaOUQSDvfMWkg3+JX25QXLe
8ckARi9aId1ocrlPrL7pngTRX77Hbj3VLl+1li5lQB4L8xMSFy2/ucPFAg//
ivgJ1mpuf2tdPD6vt4x3rupRGKhfCzTWIB6hWv+pvyn+rs1RnDHzoTpEZ4Vt
m0cbr++KekmDoS1B2q9cdCWmiCQaPPuAFhWfgATaGdu+JfgArTsH5yRYSr/l
QdtWHU5Qt1JuCwyHvlq5ejeaexRqcqFQjMnsCp4/CXC3KgSrdJw5NuU8R6t7
ywaSaAMQ342yfvRt8amI9qNNZZK1nGRZRsqPuR2KqsB4IaXbTbVRHkkoRIq5
OH93vQAbj7FLxK91SrmHJ9BW1t50TyXiz7TSTcSs0AYSedfNX73+m59cx5CJ
mhy5ZtxHOqDA6Eyd91naJHSY5sqyquWpKZ2Zb+VRSvCIyxeHEVaYPWHdjRDn
gIg/LXrvrXy8v9R5xlEyYoSr8sEOfrYcZbGkTIIyn0E1ZXqWL55n8FYDyPVA
mhKQCaR+U9XJpF4t7iMh4Kul4T+1RhcUbSiFd4gK6EA532iX9enlserQ9TLy
SLkKQW7FXFioyDyN+j4aF7olJbuLbTCpB979sT0e4FxAc/cYloSjA60vQy4q
ozbVGkhnWY4I6Zr6UOhdNNpOf4jrfDj11u1TRqkEpwUnE6Ys3/TF3LqYVMGj
Zbp5dCLqkJNRPprLgcy+1ijKdrrt2yYF6Okhoz2VqGtXJ6FkdQEq0EkaneXY
782jiXfBG6ELcKAIZ0RXeyIHBWBUF+vwo4cdQetSBZNHsi3lD9f/yAL3a0Su
lma8P+8PIEAguCetuHgBl/Zn7uhw5jgbO0ik7kQMQ4y6H7s9UySuW2oVC32b
MXE/9AOfzBPVC231QWoWn9MYL7JCmh/sTC3umM/jz1FvU7ScOPeMLsS2O3Nd
rYxCoBOLPenXjTZkZO9TuNu5HSQl+aDdR6esFP7NGJZm8ONjWHJcrbKpVxrl
DDw9Ia25EjJ3wABCRPWdh+U80XH7wJ28eabI4I5hOUR8UKQONullRgftDuUY
hdQ8Y0iuTSX47T3ZHubZggwwQ58EFTncQw4K4GAzcRng8Qf+KUwX7Kymq7Gs
rwvnIYmm/ToSi/j0rcZl9JR5vuv9/fjf99J4r/5y9RVOg6sooxf9OFVR+Q78
liMha5CKXNc8tQZPD43b+fXRHwZM5ip1SMKsCGpnOS2v0ePyI014mIwUuSQg
nvchk4vW95FSnTDCJzZAhyYyD10wFsU34oz7LXe6/OAEn9BxURCfCbyDgZr0
4fhbN+HcdyzoQmJQss+XbhJUxQmdw/zqlTOSPCHHgOuvRRhdAXztB1GQG8SJ
MkxV+54babOeYAiWN430ktv1uKL80z6NLeDrBBxdevVJ0AvQIuRYOcFh6NH7
p+kjbQo/0q3J05J2oY21KCvdTzDFKFf7zBM3quQf8+3iPt0BlSjsffDihP80
CzCg+ZCwv90jucRdY+ZOWaOkPNEMq9QLJZQS2oWUbKTdP1XeYLMqD2T3mYnh
u8ZVX9RMMbndhjmkOZ+IrfU4fo9m+pYPLJrRusGFgzx1tlb8NypywPwEcOL9
RsS1e2D8mXoAIWgHsd2wkgbT+U7aTJNZGic4G2+PVH/8v6S4ZC46lKVoOjE0
UtKcEUjXo8MrdfmZzywfQ53Tb7dykQmQhJ6u5JZWCjFvb5y7FFtPkcQAu0LM
BbvbReBgFCtJGUT2gMLFTlCSC12p7XHqqwGB4U8soB3TLHz/6Zguln2VHjdR
g3aSvIDb4xkwUsoZEFyrucB+C+VGalFM8KZbIaEPtlrHmbovJ5hNkCWu43iX
71DXBlMw49w8Q+eE6Ympprj4E/EBHx3mIaYAJDgjDpJi+nU/8GBSOQqP7Xiv
Q8xLrIkMpKMM4Zrh3+b3G/frx6/VyjmikTkgVN4v+KiWZVo4LWC7utMSyybr
DRWXo/nlfdiDIAxTJE3dvYZ25gg7ZjHPQV5tFv4GH32ZIS71NvrQzBD8zYDh
HdfjG5l3P63nX8WbfxHc1NgchLSAsbZnIFayeOShPkEiD7ZQR4kQw0/5EMXp
+Cbol4OQxj6J1l4Ar4lOXTLBm19eECv//i40Q5so8Zt2cA00VhF9NIC96/nn
PTjAG+h6Sp/hfOD+GpmH/ubmtebC+f4lxN3uAzwhqSVj2cq7rViSLKKAZec3
UKis4yxw8SnvwzRAbQc6DraU4ca2JjmZd8W55PJvB67pbF10gXCek84ufA/N
CShi57ifgRMvVwM7d0AnMFYpaJ9w9Ejx0hF416tI6HGNtKxsIvmvGQuzlbR3
Z64MxMxgwthWub3sZSC2mx/kcYrFU4tQGg7Eb7TZSvHBamwXwhFxT4oqvbLT
dQnW7XpSUVF0cqcVowlKWG4BJOhDRiyyxGiyX9GIz9rQX7k9xxq/UeSafWTY
6uCgG7a72k2pTtywzCqcYl8IqY+xD3bNq4b2X0kI7dTy5B87UJBfdZOp7jPM
9gf7Lyo3kEhza6o9X8efygStAaA5zilj9n5PfO177Rt5lzBp9xQWjLkHHBxY
mKLyRLTZlD7y8B3AbLw1iyuZNsKHv/vX66E2fxOfPFyJ94ZF3UH0n+oKggly
PM6ZMoyDC+0HxSzcD7SruTRP89P9vtCRE6hOazPC+EJT3IxRaXJAOS6GsGHw
JaYjwIGJj9QF6wWu+Axc66P1T4tCZEhnKuU2gBagTWM7Upm+Q1HvCJEhjU7T
y1FU4JHrjvFWmpN1PyEtLwhDeLxMQyB3GZrc0QixoHmaRdnO2mEbwqNXfcty
A2cSpF644Oit6g+Ys4OUafT+ttUGZ6zyvwrpKq1QZE+h9Ge2JC074LutnXf8
vgTjjoSBCGJpaTtnXMEReJfebP48IlkB5WBH0Ou9qFZ6p9x6R5EVYUjxnDMG
UJOv3n3oEslNun25QbK1YM3MGeaa0CPaNj6qk36mCF5d9bTLkBb4J1qkorq0
hZvV51CsAUCNWvpqPV39SGI+XRCaCfp/Duo97AYWJ0o60stIszGp9JvMhrV/
ZYwcoeyjKTStVpYnJPiddo0EOSJZf0TWfWo9mPCnR/SjN9uWWeTOblfiT45h
cG7lNIAVqjBdWxcfHyZg+9WAjCsEKMhDe73wwf1YgCBqKEG0QY5HM+uzo7s0
OmdNRTmAZ2HaxgDWEBkFmHQfgX6b2O437Eqihl/aezpJ/S/oMyqbwKPjf7Ab
mFtCvE+EWzvA6QAz1wOtqDlz2PA57dVrxYb0on4Hvi161J4FwvSQLsIrLTO9
2VcJ97irHkXwBIfOwMhBmfWqsnCaAORRaSozOdhudZx/pk7+m5heR9ewM9Yg
gw4Ys7mXM23zJUg3Gmq6F8AzM+xpqgGfp3PLKuA/G1nAQCiY9+JlR8P+4zcl
XSRNQlnTmmsj8Hy3b5UDBXv3nsF6joRrQafPpGFBXzww2ts59gAMuHEtSpXL
jRSI8qaaIe3oN3YB51q/RW3TG0sb2KwDYh5DRKJAD7JsC85phyncnhu9VFoD
YsZsSnz1T56lReGn1lJQGUQRN9SbYO4Sis2GmMNnqq6MZ4z55lNYaXITQgJ3
0OtgL+RWmoSZupnmDenCOQuGpFqUjMCWShbJCtrMy/SE2AmLEqg+vYBkkPD0
WLGwR//kRGdSrKRaDq2l5hEtL8eyA9yp8rPINKD0Q6S52ftWU2jmDxcUO5iZ
7tVWeonkANuDVdZDsVru+YxDl5yFki9VDRTNkrykYSmcbRJ2DTPBI4OqpRR5
fWwR9ar5Hx5E3GqdzjaCYoZHX5nycdscOLxspyj45aeWcaQ5TYhdFXGrhWGw
KtM3wcEfRv2A4o0WHUDgvKBbeK2fW9UCj3qJTaBM4wh8JzZuYhKIUMBptqu7
hlXKEsne8PN5GcKgOc3VQVgQj70GjYmRI6eHQmMntVjsXVbhiAHvMBrD+UmZ
j0Q7SxpMwaxiX7ukk78nXfHjrU8mcl+kdytq0RdJtAK1LTc+uajahjigz1lj
TtJxxP6qWSlMiRwqS+vTgIpDoZ+y5VpfXwNQWO+/nzGV7VKLiP2/76TxtuWL
VPS9XLzs/4LwNPrVYvG6yluxuWZ/xYVpxb6wdESYAdh1VloCPRm7ScqSgrmw
kXTjqSmVsmdevaWgnoz/PCcjgl6eOJpadwR7r+SbFsYkX02FRX1DeC1VJDFC
+4fSY23fK2f2OzGK7GJDAC7CI4EvYNaQb8P0t2Jmd/6C9BsKQ35Fliw0TDsL
okm+4W2TMZFnumz0ozMWzzGpzVeXrt341XB6zI0ATE21cZAchIO09k/EUbhs
sBa0B8t1/qnd508eg3tYEW+xwkHRXbweHaEkTjNcKGFeiHw6ojmS1f1DoE2Q
JF7I21GFQnA6ZgHLa/Q96DydpNkIdGVivZcwhuttezGI1DLQwgSG/mSF1kZj
5IhKiF9ZjijYOFq3kA8+l+Rz2UOlHXVUl3aLvYxk7I/H+l0JRML8A0TpvxEj
B0esYi1hqR+DWfHoyt8o40lzmLERXRQGaD60m7FXlnZqGcZUXiEyLn19VAav
GULFEMAJxcLYgiBylWT5UeS0tDh3ZGbaHCr9ISoKDAouk3fv+oCwCU8CZ1DS
vUUVskSmSc/GTETHhai/P+V20FnqBDdxaG48WsKuy+1XCirVf1a99fhkYcSP
d3Ldi4e3lkW9+f2UdT0sQi7Dm3n6DnMpNug6cUn9wTip2UsGhOFT+jGZmQKm
CwMZwoNY0ryF4EDX00Xd0X0YFcKLNDA/6aZ5Xazx2qikenKhKfyae6932GJw
ukx8lxaBEXpuINJY2c0U17XG+I9RH9EwqU8DtfL+JVWxP4kiO2qLKcPk6JQW
wCLFDG/rmG6LAViVwDz3PWeKuCfdpDzgbOHvTERsWJZTr60Xnt8OM8wyHz6u
2noGQ0QU3D65VYR6UAMXg1g5Hc+oJDBXHG3Nymbn9QEMhdJRA9Ia11y4Pe/A
29JsJGeblAqqiRjfRX75H3Lda/jzlghK16IU35ocKI/AnPUzbFHlSU7nPq9E
u0kpnpTXLDPh5UnBtFK8DQu4qswEXxLWQkLewTbAjjIRgo71sp7Z9xfHKkBB
sq36SwZjQ/DXr/wT2iNL2Clsmpi6x3+4WRZkLYYe9YBUnvu58/ZFVdgwZm6o
nVpH4y4ZlMXo7QznjxsOOFwhBlnhZhruPEnc3/Pn/eln/jsy5Dm1TumgmG4I
rbEQILVkeDNz6x0Y306n0tcoGgoBG7YivLuS6KLJ7UAhKQvT+jEuiXy5EXeH
ZSz93NqcJeLr60Ij9iwSf13jcLggiHgr+VfpFeFTbx35mFdiDyZUaHWHN56Q
TteyPlyZr3ZxHeQHAtnxZ43gGd0JYiQ2Jv+wVn464J3x1IxSPMHRFLTQTEFu
hQNs7da+6yiXke6J2+kG3lDXMJ54dtgK7ftBo3JF9oeTD0NxO+eC67QdadC6
NI/rdW1WNrfJ5yL9VOnI7rQX2qzPj01RR3EltPdsKQFJyftS2790KvmuyCAG
df/BCWhc0ZnDuseqfkrTmZJ4QaGJgxF7FG0W6qyeRNecYKzz6uIA5JJkALAv
unKexZYeWN9CgF1XKKE8ctswAsGZcg9q5gQl3EVcbh17Ru6JoV1kUG5i9qyQ
beltRft/2RnLoImjeGgNwbLNQT50Ykk3GhgZ25vJNffAuOhZ6sI5Lu3hsWN6
cZtbo8Kh8yjZlC76Z3vzOwxoKbuJCErmcymG8wtyzkRnJJnVBOZdbNnxoSjn
mV8u2roPF8X2j0toUYKT6ny7WffEn68qcxPhRoRBNMgupdJ4Jf74GvGnclRx
WM0N8MX/gq3R6NJie2UJCL8+nkIiQ9qDtherEwivRv+VuvV7sYitKNxwYl6z
P0nRg+p51B00SUlm/FHChNWOzYW3ETKluis6w/LICGckfArtFn0gloPud6ci
vvX13yWnHbNMC9bdyN9GW8hgThk8O4B61GesmsKNyW7ij+RJJPsFY+w1nNap
SnrtsC0iR9mXpNKUvwxYMba4LK9dkD3nIS9CzCjE2NNiPOPlGwB/2F/oOoBf
dEswuHujDA6O7P0jnxt2PeQ9cFHJ0XUb9hiqT+UmuWoWYIkiOEs6c3MZf/Hp
FryDzKxZDrcccuFCCdN8u3AtRMsTF8K6dwNXgGS8g98HHDs52YzHwJQN3Nwc
+m0Mg6JVKMFTOToWYoWHp2c/iuF7Jj/zPwarpIZW71yFTgk6ZRnt8QCO4b8P
a0Y3iEsQ0yk5iBzeqUtxybqe5u2rFJ7EjU2DxvIy5UmXxnwouQqFqHeC1EdR
c5CQ+M1WYt7oiECjZnYDQ+vKN9WKKt8bPFa3rs/Ooqap/bE89EDAr8IbENgi
khGs/tQ6zXtK4TjUQC8z3Tsk4ULwtNpLCGTQ+QvzRk56/03o5NX3McgistrX
QYoCVDFApAgoFl+PbmrVo86GXNUjLOSKdh1sRtbpXX1Qwjoa+WM0yEVStFnX
oPss51Z4Lz0MKSRohNJFc+XDo6JKAT+l5A0scWhxe0zwaZiR1yvWpaasmRz6
YlntkmkgMgCS1RTcPqyjqo9EEqq6HFEM1TwUEn3HIHr4MTAMY8mLMmefCkK3
Qg86CRKUPltXF/n96xT7CTie9bvE7ZIGFU4wuUkfHXHJCqcpLNgBK/XSJwlN
hHiTkPckP0qGDjZQO+WFH5qvrmMwTc97fRQVQ0nn8+Qu0ATnmUoQGb2z6opf
OxcIwjT89twUvdaaOeHXdrIjCFYtFUqEt0jMuZIHyKQOviczsQG+iOB3cs3G
qc14nu2ey6z6DHhKvAc4cjLV4OYLDq1ksotA4LAkk+0XP24qADoz1+sYU3+4
zMziqIZvn0+hb4GiJzYeZuM+yN013fAoNG1QgN011cJ27ppDvLvUp8meZs2s
DLq6toZf7AN1mkmH3Pz473roq/NLy9O4Ozup74bdenguMCq6X+ZYduhVXBVe
eDgEAxQFrhNHbyY3WLgdZsK9fSlyL82HBaAeO3fKOumilvJWS8NnP5AGx55W
ve9DEPS/Cyi03QTJHPLh+qyRMHLYhLVOGRexdZ6Mlu//vR2FX4JjRPkP3KP7
hqA9GHaviqzGPe+N/aD7QrYhjsAOPYji3hii7w/sxY5/BPENhEoxSkBnRkHF
I2dAvYayB2aw9IRXyjP5OuyrrVh1MqezQieI+3CVhVQDkrPGBoNZyO34PIov
tq4cP460PXGPUSOoFsJBsQG17aEyg58wOxnfCKXDGO6s4XIdlA5GAjRO/jGl
K7nxhF3LFob6YuBYIYsRGomdZbHi+IcjCUWUKfk2bJGdLjRX3KCvQkAVMKhU
eKmKjyWsPAbWclFzAqxupLL8cJAYEP0c6eKKQ4PpfqOnMh3fxZLmhJ0qrg3E
nQNKjBHLjCvPK5I1T8jmKfYVhQn51TPtiqvzP4wMDGF5euIpI5PIde43rqPC
OukjNhd7JQQb2dznNRDuuvdgmII3JOt6IpZ8MY8ggnm5BT+8blkW4Xhd2+Ys
FMIKM7OSby4K2S14HHBRlTngUdYUBZVo+dCKqfagBMYtyZ+nwl1j5KPeP/UI
A3UOfpMjGz7FWo4jrq/uFKJC78e4aLJr2SzbDutgXuJ5H7RhDV2cZKJ00Cf/
T+nglew/kWkOyB3afZM3XlgPMTqC++UBvJBH7Bb16keGsDmi7+avgYBrPAwS
fypLj6Q1u8cE3gzli8mcm69LP+GI4d0kI43NDWPlHn2NZuCwxldSgSGamh67
gSRVtZITqAKDtbqei3cN23QvMOq9q07BVZpl9ge1MiTn3gQU1wZcVAZAYxEI
8r5/EZ5xLpmKxzVClsVMgpKeb/URn3pQ/winRhtpav/mN9RzqCLAY5g9sOnK
9vALHf0cXvTYnj4amtoiP8wXsHo2Zev+ExoJeLN/3shCAb7rpqO7ROknen3r
XYDNmrDqbOy9p3DXyunFT8v8jKcbsYcIs0EOnRCXgF6oVQ9oRFPoHTeEZxEX
rk5y7rrysrgvqKVsX+/WLfBsI07nWCsDC0cWNO3bCCizpdOijbma9fBp6bBY
LAbPsT+QhTfPpWME0B+l5EwqZJYZRd+1TzNKOFdFm+RSP7XsnS/0izSZzbIh
qP4n0uyDNMdXYV9x0fq/DCygVnhrFgqgZ3t6iGiPtKcbjRVMNai1SPZKjIuo
Pvg3zQCkkfCMXvxj9Jub6aPUVfCrisfQlkuNWKpsKG1/2oBbqYN/v4OfT+Ie
GG77+RWU4Jd0BK20zZFjmjXX2+2v7YaeU+JCdObSHz6gyL22EYQY2Z2dyyjX
ZRF2HJ3UbAjBZkltA5cc6LUYEXPOJ8b2MnXKXIGHwGsAakj/zVnoJQRLPqvM
EAW8RAIS1+I5eydmMLo/HI1KJ0zRO/gJJ+spxMRF3O8Z3LCLaUDgjR4+AHZS
N1WvQ/n7oAloUmqYejWZKtnA2D7PCio2dbpCM80eWth2mREnrmofHSGkVi9o
5t7I6R3KdwAMiceB1OqZDiIpmh44CcGrc2oI4jywIKqAS5M9cR7ySgPCA+ET
l8WSX5hCp5USzNeM0iy53nPkc/I1oZ1XNfCgXK4p1PGp5l4/kYktGy/zNxyr
NDFpFJeZrUDhQeVU1PXO8/9TBGKTsoznH/4HtVyzB2bBDa5JlZDYwMnS+aBM
kn5ZEoBQHYbpOKtPWZelpCVxLAFtY0xm5RyRPikRgxERCVpMPTP/0e4me7tx
cLFqNj8EoEyWtvgSL1g261z9zlJTOkt+3aGm3pc/l7zN/DcQze7BfaZ0Nd5H
dX1tTOIcl/sqPcFhN/V0zoJTBTShoNCgtElanhiUAfcQePThtvijMiP3+2eW
qwhVYv8Ybn4/lnGSbuVQepN88/HHTLoSZJ1eaeKxS8M9hZZjjRMO1NBFr2w3
+DcHT0xkf6sEasm/LyVU92hVKp5HgSQdjr5OzksIGC3KgCcL6eAG5hWLrGqk
iddCzRgcg7BL/rkQwAfscEt8NSbl9pyqy/W4oP32WUgBU0RabU46kuFN/OqU
zzCqWJCsacdpQmSojlrkEgZGxRnzagUZN8vZquiXRKXd0ne24GbqttcvpE3D
0CgaCUCSB2vfKrcQHZ78FI2b6x4ri9YGgK5Q7gtH94E1zkC0ntkP6oQAgfCi
PYbiNh6zimefyI52WC48fQCgOgN/ucl3MbtsNJF2WvgeoXMVq+SfF0pcdmQD
t0lzy1mVIwuHi/bdCe1NCfnmZVQClu+OF9dPxQAsWdpQSQJ0Ze4b/TYawXEU
j0tD2LEzRfRZe8CupCM05AV7uhv28UkU1Q1XCNOMZJd3C+yJbH+8Hw/zvtzb
tXQIvtuiKpG0CdAw0n5ssaeXk73AowXFQW2LSA9PfE/7JCLDuAuTx9y8V3VI
Kn1IzsR1czNSoZZDLpXWGTL0IbhrgsIYgTrFVlDRJ8HBe1JNN0Lfa04SNdx8
FbkATSJeQzsWTZ/NWWNUh0WRgzY3FB0dp+aQAyXnWH2mFB5txD7jVAXMqjiG
/gyActF6RlVCi+cptb39+xveHEG7sfMgMTpI+HA0gZVYWxKj6ZhB9ATYNezk
mOHgoyLIvuP0pEF8SbvDekOarzqzKWkMkCh1FGTYVjTYAoDuJkx36lOObTrv
8g4fGHrm/95BjmN/vZ3bBYSalBnd3a3mexUktz9lrx693jD/9OXXjGcPy0fy
R3HXtbO6v/eh+ngALIR8W2wpK2cc/qd0t2pfUytcMt6cvEuOHsEdR1ARAkd4
ezo/k88QupsiPXxWebpbDREWDTmCyJOD2Li5tYj9j3pQ45i3QVXETcvLR93o
o02TbkHGKKgY4ZwW0K3zUwtqLo1nl1YTvSl4D097bM8kzWbPaOnnp/xwltrI
EpTaGFM7C/lm2/MSwjx729JVmN0l4lvWdx1jgL3O5fblmGHwkHX6saAglZUq
deIzA9i7Kg3qcMGGY4S7jVVMiIGjjo/x8Tl3uDoRpyu1rHQtI5C3QKG6bEyh
bFTUClav9+f0HJKOhkhSrWL4dcvDJ+rrfc08Aa5HEpgNTvBqKe4NVdOhBwWI
6Wf11pUcnisTgBUSfRpk/HskTowon9I2cJV/2ewZKWhRfBCApL3sUHQRhlWe
udPrkvPTKF/NQNdBPYwFUOAUu+W6+m4gLmwRVltCkw3sQtECvsOIvq7nHCzi
KmTzmujfPcMju222E2aalvbmKtbBOKcRs4FYEY5UJcpJ9ihR8CteMwroppsZ
kpE7urnI7e0Z4z2cNEOgUJSzjk7U+e/JTuoUz6X3tAidYgh2Ridu7pUAR1be
wjaj+BKGgSx8QKy//YHVa0WYQleV8LSxQl2D+seJm2aBtQDVa/Sms4ENahuS
TkYfXlKqYVCWX3VXpt2UcuWtKWrYq2zfpTxlM8AgnloQo6hYL5cog1xsHyGU
sGelgJ5J+5CW+m7qvTxQSrAoU32lDaIwTSkNIwFcGwUIooKroYIF5I09ZCG3
amkxnbZ9qDRUmGo3U3g5ARIVMtTdVs4ZmOGZSLW6qI4OC5d27wBB0RWKc7Vd
tGYH/Gpt8gNLBXe8Vfxlu2Tr3hQSfx3zZAajBS/B9WPKAHbSIrENMqfy5l6D
lcYKHUBRDTXsMLlTpQLc9wyOgF24EoyTivx+KUN1Iasw87YwpuUKsud2+DFZ
00o6UEV07jmtZ10BkKE+j4k2yQxde/lLuMLnUVz3E+2ZNkX8ZutLib417NRb
VBNWSnC841EYBvEByrwlEmWskHUfKs7YYLHMXYBduPlWrV2EfyeHCMfhv5eX
BUUK3ybhf9hMM0x2yAAjMgiZAYtrIoY2LVqr7c8AXR4A/+fNTUUQUDMOyM+e
1uJ2f1rp4N6yCpifyNum/esgUf47iX0uQl2nokhzCEymUwAZE5xO7qZL7dLa
yUCZ78vlqiwRau0d22MH/y9CyGYjrZ+iYYCBtrljAkJU++/6LCYGVPZIOunv
pNEfNMXyq3zIURMy6pfT37/lc89pKhUx4g73ZDnVoiPkhxoBP2Tmow8ZaGlg
0BpPcuxpaTq8Xx+XHcBvL6JdiO1gjFTX+DM/XDHFkjbeLony/iS9TpNZg9A2
6BfDYH1zw+1UPuez0llors/5TT49xaXnkgwE1e6J2gofeXal0TBRM2F5Ky/r
iSj2IP8jrzMuGHY4ryWI+SehuHeG+pKg82WvlReF6U1tuUVmgl9JkYbWO476
by4NvfYRbUrhDKtG5FWHLo4bkVUGfhGVLZyopPcMI/2vVBSbmZmwgXYj/AxW
Ib0ArPqsE/hLdTvHnBu1UhNNV6yMEFK6jc4W3JuFibO/4A/14iScrsmoLZ21
GuU213frm3wta6dDn+1qJlez3NNmW+i73fZYPToGngx6uGaQcAPJqyf18Wlf
SWiRcZTcz5LsH++AKR7ReUVZ68ROVtFlL2ndXc+3c8z0nc0uIGuFW8ryifaz
81oISjDw97KjBj44IcJqOtzfdKAgB++ZNt+3yss4q5lm/VgUpuO7k9ZIvdwS
+tYhMGyrUPW/Jrzqt9RAQkmQIZArxOr0wqXYHtgg0ScDMwc4SSW/mUisqbNA
RDDhtvdmxsVvZFSNZ6FDOv3riJjxcLPDdJRmdlUDQnjnv2t/UaZbnGLUux5a
gjRimt2bhijzrcsJH2rqP0Mzokz4mTrEc25nKYABMDXw6yQWClmZCVBEAjtE
KdemV/4WolzpXnJky2vwN2OYiTVopBozqM1CZiMlKk6+aAUhRYBgkNbR16p0
LrgnW0eH7NvDykNBGdtjsTrHckDktC4EVDOXgw/hfhJdoslTEVbMo4qZeJfN
fajQ7p4mTTzf6EJfHFzAEr35ocZpKyyagboZKt2XAQBweLnnnAkj3UykwE86
hKtwFV+DsE/BCR0BxcV53nO4I1xJ3D6vdB6QaS+BgNRH57i0EyfCBF5fWc5Z
7k/tfauVVjY+Ho8vmhSdKR4Z9ghztyWPUo+Bp0bc7Ms35rSNWQ8AB2i9+OpS
gMMw7tnIPv8IlxfVctl2RCL7Hft3eYK+nH04LGfXspExHhAqriUkXSSnOzRj
/GT3QjGo8AttJec5lUFHFT01vi5VR1dspeI/l6xOqik8oJslj/+Cw0RmRof2
1e/kW9+ihcR6A6iD13VwaHlRnEPxKBqpsimo4+aF9qMsSAoUAK9hfgUxJOKV
mQI012hmvur1fabuB8Ti8Wikj9DggAPaHufNKTbSnbfki3fTa5vRjx33uFZB
cWBXPEimZE2DfH5voe6AdDCO/++bpe7ApITBQJTEKa/UNb39DVNjA+VQYSrg
1qYbrT1OCOaWLE0BuHiMKL8Ch0QTQwHp0AjMaSrJTWlnsThnfspbME160E+I
ZsUI8U02lmbD43pJv1pbFJ2Iqvq99i8hq/5K38vbVgLA71h5NgEfVZtw28th
ZeJ9wWuygR6Qkf92CmCo/tKmAqNogwxNoBNRKukn8UWN90D4/OzM2mf6clY5
iYss6jrSbXz92/iRrrUG3CCkT8Xxxhdlh2j1R0wW0HBB0sG+Wih842aBaFq3
LEsVH0WjpS7FlZDgNm5kCvNZtGr1B3ZcIGar4wRo9nAcdwE51Sz4CgV7Rknm
lZhknbWrlax9HuuC7XhKTSlhrI9fFm2mhKMIKqhoZlLAihpRDHYaKThP1Mr2
YgVxc2j07g3Uuv+J+0v9Z9Rfcb0C1VXgq29InDxPw4R9LpdNRFNfVj/QzxFn
2k/WZWE6zFBXNB634VWvaPzjfdXV4CUt1GDIPwimkZGZ92uUzFd9SfkQ3sUB
cnW+Ons3FezHN6oRKzM11eD0hPI94XQQhr4x6D7JUpQjATAj2GRCNvlglreO
8d2YU3lOqQjREoCyGHG+HefQfUVFbUSbSJNg9rzu7j45cXS3EWiyG5n/h4jf
6vaAGRDwTkHxuCgSoymFWqNLdjy+ezPhizCVT4XeUZGXLs1qGB4TFA2HDcAk
SrecGIoCGdi/qtmt2Ggcel92k4SPg7B2CknqkMlNeBTAH55S/l67ljnQdcqg
Mu4OByA1Qt2iopYnHfBxAekFdLM5/Uila/+KzScsLNlZ1OricgjEp+X4gmKQ
hXP5wLV9JVpM6mHgTqsD7IGml0EvsVJF+z+nVJYE3lF7ICz5Yx/vEsWYjCCo
CPsuYQYo1WlJYndAddoYoKk/eZNGtXlFKo/uPty59tovCGIi6zZonu5r0Igj
ygOb68HzmNxnK2AKkh0WEKj38bkKRYPRSXieIaXrr7HnSzzI8cKBwiih8cKC
acK4nmxbgFFWR2sgxBDlVE7XYSnkr3waKPAtSJNHY4CkeODsO8MHwKspQ7uc
KZ12rL+PlZeVb6FHkf75Imz6dulE7F53MB4daDU7gt9IZOiH5PGN7ZV16lwy
wvifeSC1vEMpLCcx0UsE+Gw9Za5gKxP1k6aXd8ixZHc+jo14J+XjYz5Qi6QA
BGOlXIIcCHG8dfMdTWFBDJa3cHWN5cV81v52MURdAqvDKMHF/fBlcyrHqVaY
rMsGpPGULuIWcOf4LP44dxDLVrcXiCu5GjzTsdYec/5OMGTEnkcfo0f/yjNL
B6f6T1dlriZlgopNfmC/ncBIstBXMMcGPkzNo8byK2u6TRk46pAjvHjqB0Wt
gfrRughbK/WB3Amof7+UGQS7JsSmlEuxodEDYSYZbSulGr3JlTIsoZXmzmXH
L4sNi6ALYI8dnCeDjkwR5X5lr4kqgKMIUTP+karIOzioAdUvMvwXHDmx1y1b
Evx9Al76rkhzbcb9dv2TnCJ6KV3UpmWr+GqHhZ79q1xi+PzGgP4sc/X0duHb
+4reIFSSBR56/FSS+rfDnlvFUrRwbqzRUzyCUrZlPEyLui0FXyBpgFNH3IaF
VyolxDROT2aj0d6sbWJ9ImVI38l+nPf6Y7Cn/pBiCY+Rzz+mY3OaGWQoYkAd
NIHwW4jiEkucBM5G40VKI/gPdPIxY62F1mSqVQxWLzexPPAxGYsE9qYCoqvp
NYx4LQdLd7ys90jt7ovRDP7FC/a2VME8G1PLPBgvRwVkxLF+yRdlu694O2Nq
82H7uNURQlaSsqdJGSk/60i/USkixRzbQqyKxVRl+yb9b0YmncIJPCrslsLc
BtH3QjsB6kDNlh44kzmAP+yjTEiVwm0I/cU48R1ChjVczN/OXaA8mogY4Hls
jSkbZj1b/nKg4ge6mk4XNCqhLis6Q6bR2E4Z6tffkAezON8iD9FsGmJ+TXqg
/R2ZtNmeZUTPEnhyernPXbkZ54pd95f4Zyr4Rz5MLH4sfnfj6BSv8YdLmHjA
8CogyEqilKlBWJpWHEyVb32h9k198A+dLzOt486zTH15FbzQ8yqsIjKCS0fi
S9ATVT0OJNHTwwNrVo6t2PBY9BcoWllsbhqSnOFOsQJs4BMm9XKLpy0YGrSn
JyEAaWXYdpAvdqU5E8zU6VsE2VsyjZL//GBr5w5ySw5gBaCqj3KO6BQutW91
CeGE8yjNYVC3kDpi8eh5jIUmUzKTzBilpOCEd0w7Qg2mc1P6gmy5I2A3ke77
0ts4APNdLsa7gmjL6ReESlveiLnfPmB5bZNxqRm/9km3RedqwvlfxKk8EMIO
GHCW0sKmICzfNKxg2fxmvw+Ls0i3gs+qzzf3r18RWgfZz7iYIgoZxO9jPWoT
gic7gWDrqyIRUC4ut42Mefff9iJ1Usx/auXnUjnHuUpTa6IL3UBr/vVNG21V
umyzqG2S8VDr5USIqSBB6U6ZrDQ3Dj4QISdGgxgj+oKhC0UhMvqqNSrbzJzh
Prb/2A6J0kpC3MKvUiQ3EfhLTSgh+GVigPfMr7n69n9Vo5n7M9cb9Yq4O5+7
I9ivU+4mI3gteS2sKd7yAqxz7FrleKUwXJZQ9sSsPkg6F9vj38nUfjBh1ORk
Vjx7Bgd0DseWhNu2aQpQaBI1crX+18UzI2Ogr5dwBU4qX1cuQEy0xe9tv+zc
B5hnDDVtmkZ88n2IsBgTwnk3QEG0pvyXc23VBUfsx2uUj5P4sH9y5A2JDXJe
xzg8tnZCXaEzIB1qki6XXgBdu+Q7ujpq3c/IutNh0dbtMg3m2ZFUlgMuZMam
v+P2cJyREYEseAOMIllskQKxp6w2/dO0tilVHtcK+WF9pYzoiF3cnU6h2IO+
v65mYVsorT3Mtye2HubMOxJ2nuyaV32X4yop3qcoZRZiuBKhq03Af1FDm1s0
hDqnrVWRm+FBKM1WGauGXJJGtXSKcwtQjUthhI65P6SSacJhBQazotxb1mGJ
4CKgCoBN9h/QeqvjCYr8X4SsgpY77ECqKFr9w3F7NgpF0f7eAR7Ef1SrzF7g
8d5BY5121RjMgkrfIJc78cqfncHf/+UGmdgMo3pqbh9c48jJWBdxUVxlhwGi
9kwkDloTwaY/Omo4BxO8P817DFmvrEqdsmb2rNyh5BIZ8Y9BlKyIHvuFGx0A
c9Ea49CFh1VxZSJPGQSumxxeg4AYXBk8b9dw9IQZSUEQVhbmBULAYQzBstHU
H/lHLtbRJjMG3JWZ1b/YVJugElOo7opkB/vwaDjZrdVhhWbzHU1CKoKOyzZq
/Y/v3/lZWB7c3RcqwAfzZUeZRqhueGl6T6jADhVJAeAj3N10JruDI7tqiKft
Odg3IA3ekDWDMNfAlYsFBNi77KiXRtO7Hk0+sXdy7gUzIMOOoSotVNQRfq0z
0k93obkpi1MJvn4SXWm21tH9TizM6ghVD2/BgNgiXd+MTB+k1a3iUOpfxQlT
6L+Ye2F4IucasBzimYIQdUDVom9XaVOHXroiQrcoCHkTbNrx61cZv0yByQXM
EgfTHawT+6pNQHDYgD7G90Nw3ESvTRWzz1SHqgvdxWD8RufZ+3KIFNi8fXsi
QCNfk6jMR0O1zmrg3h7G4p81tdCtWRkeb9HFvzxP8UJjWyPf+ISI59St1w3V
0nKnNM6PJHbRy4nlJtOwZdDIAiyC/BXN3i6jNftLLXeDZvs9MFe+zhG5rm03
n4EAnSpWhVpuke94KYyk/pUQmNw8z80EH4DRx4KalRw/cRnPuZ/xYmdxDxfM
v+YhrKstxB8APy256t+MUXTS1VESHY6y42XfV2qfA89Noaw2RBpNaLfMr9nZ
vAAOjdONje9+wqldMyG6HUP01X7pACGg4vYeZtKPgjCFDNnFcCTwpNHcYR4Z
lQagcR4rNP53yIu0ozx4K7YeiArM0ywMaRdMliI5ZMKrV+4AUSZxx97UJ3sC
3aK7F2fbb9+yidTTpyv+cbLS0OgCqkKi94JxsmStXUNPuhOE5Jp9WoqDxjUL
GZuhWNISYHT2EkwHsrmhTZp6RdTdsS3Dduy8ZBhSyUuKKUcvWGl+ykuBaQBz
TwjBlvzp6eXITmz4Fsan3ejY96WKkceGm84xxAfVnDBB2mqYzRnr9ilH0C+O
Aa38L2fTqzDMrMqIYYIaFrYZnmaiyw3o3tWSVzn3AbH4XufEPsLOAlmzt/Oa
0MqAbd2kAHI22mfnd/nQn6eXVRezROEdxXRTxD+ioFtgCCkkFAsdYld3iwrq
QOWbDHSAeF/57MPvmFryOR2H/yD5rvFApoSBwfEXO/sjEqpcQt1aMNeD3R6F
YTZUTT3CL6sW2GhaXGtTCVvUSzf38ej3K9xRX5ZG0xgPXFbQ8yioOXjDItgN
c5+nWZcHARKiZgWViz2owO/Lj8SHAbcZxFn7JjiV9jalSWV4otsiaGu45Pk5
VZeWNwYH4+1LOTiNHj8jukdfcde6jiegohWm+7g7FP+EHP8pnm6vpI4Th88C
J6CWOqCk+AgsXO4woNhxju0qirF6FlETA9Y7frP04wZF5vcpUzBsXyVVlkmi
jXZPd7lNo7iss6YUN2fHPumoh8Ptt1z+FYaYNedXpghY3jM2o0WKZpe3WWGc
L4l+GTp7RmSob+07WX0ABWuYV5piRMgPJ+qEW1062fQjEpQkcdRSOry+a4P7
GgMGkhnu81nUL9ie9BuRDzS/oipGUYtAHCkCE1kOVn3dZ9fXmMWj3dlslCRR
itTXRhbnNQQybKqfCdYkpJs4+5JJy9GCbYK+0pNMjrkcPcajz4YvWGS/b5sY
G3WENxQpx7wu33Yy85dxBLao0ROHQsaVRbIqJ1sHmQ8AlMQEVP3LZKOKa5qQ
Wzu3LAbkFCZyYHA16N670PxoXIXYFBmZVGgtDhMoUpaB4V+pTBYZcPbzuceM
09HyCrF0ixE4KV1HpasaMtu9S2R9BEKvX8n3KciNS5ZD0RqmUc2hWXqDXgAR
d6KFebhXmgf/bSSDw1oEVZaRV1jYi50VZqwhQGvZxleo/RbXN32x41qVJzi8
Qv5BMk83BAcjljH6SjgnXdcjy35iILqzMl4zQFCzlU8vZB/WUXABzC/B9gdl
S6LB3gxBmUmh6f8MD35cQXVPFleYDDAbR6rqG97eA1mCRaczbgKB8W0dtdbh
w05+HY+KqErMoCOS+dy4KJ3lhXg30reZpfoCrIG/0TnPIVEjNvDAQru30Kso
jWguTAlRoFoY7WmiimfH/XyPNpGPbhJzjwIuJQguT09siZAySW+x6OBUEm1L
jwUlGkb5oGFnA/NBWDtp85uIsi9854j9K3kNjgq4FyT7y5f0vq613bJO9iZU
6cChghIFU8L51ULBIW+ggg8Tj79XoWG0j3li21dz/m7HzlRFB8Ely3Dmb+T+
VDPGZKBfSlVSZrQjkdpevWQYF/MGdy0j6WFW9HvKwfh6ZBhafg21tMqKpBZS
BltOJ8iivbuvYOn3CA+MCilHgHLX5CgtRMy72Rs9ic2ZPt+WKvk9gy/h6FNQ
CfyouXBvzwACgwS///aJc+Mpq1wP7meLyi7ydCmL3L+0PesloJl3KpA0A5xo
TzHd5HCmeb8cmAT0nuvh+CHR2Y1c/nAxUReZMT5uDyKcatNb0msGDWjnFcM4
5GZIJ5zVn7LDTJUm1AnzJmyoBkFrmbvOokxbWdJ1gzqm6Sg+hujiZBf8I017
MibtPqA4ac/UssUULev7o6HIvqUg+7yFR6GAvyOt5382ttIxfhdzXk91B6jT
jmlnKP385hbyxNMKSxuJEbK32AhpUHJF/XXybwu20bcnwocdoSnNV3IjH4TY
SQM/42guQKuBQt6/RqW4/y4xTTyxi8gb5JRTj3diBnpUi//JvllROnrW+zGS
dlM+uUJdEhFATYqQnDO2z7kxbojz1vm58RkbXFnhMSAP+gfx8tBekanvAmGP
npi8swzbarMIT0rEhsq7DJMFrQawHicSMznSM2wHFK4Wz/5mvP+hNGqBXThF
19Qr3U+HWC0q+xi5bx3lmhAw994zwzHvb4D5bJnL6PRPmFQUrBR5uQzenAdE
why0FKyML8HtgqCyBPiA+EnPcX9dJfwcH6IiVlFy14K9hVz3y/2scRKpH5y4
B3IK7ymbcpV5o2N9tgORGr+5BCf7gv7nsdD1oz6pkGb83weWjk0W29OsOcmu
KpdrTTvk7R+9B51WNFot8SuItlGulNbjnJsSRV3ZKarTgz4lNKXXvFTblGgF
PsUawz9r0LagQ6pfBz/qhcB0VmWI1MJKpc6tjTCiunso60/wUUY/EBPKwv0j
zWVej3JeAigP88mh35g9GJpo4ae6vRrtFTHhmTXIHqa1OrGJmzCuko/fc9cg
70dCzg+h8YEMIL8c7jZsGQ4mLDJnrOHoaoqGj8EHrSJYf7PFWL7NgFsLUK3u
hVPbR463E4/jjm+ELEE3zPCUgZwFVt0uLADOpTIarQeiqmAbigZp1aHwBIV9
rZU2glr6uw3fkrHfIB89AK/HHVmsl2OUWHwMZQaZcQbvaeq9aJgU1EzHyTQ0
XaxMBIE32fl6ZwewSY8YYTFIBowSoSPiGeN3WXB7/7LyvygqWsjKoYCMm7SB
kNTanXE0i7BMFU+3Rz+41fDXRUZtOO9UcYkOkMBjiX+Kg5jAXpgBT8vENz6I
uwNpIhZoVAKx/3UChbTnDR5BwjGzl4U1KzZO6pRrMkko2R8yNpOO0oY2P70A
89lTlGZ4gpCOnG4SwUlBBKXcTLCTPg0VFaCwCDFWXz41hZWEyBlsvu78l03X
R7pVKnPD0DgYQudwiQhk+7PKq4ZPgSeyeGIzJqOMHxbwb0PXBOuoD6Ml9io6
9FtPrwPNzVz7fkoap2THIsxrlailUU03pUxafWqm0SA9j7BbJLYi1XPet1Nm
XlNaBIA/bSc7YvGcg/drcYjDheNhUxqjjbUQoSlZFjzHdwWDtD5hlbVSOFem
gnImTL+NoS8KEaXwR47eGqL/rSOlYL/ApoBvF/Q7TDApBY1CAM8T5gHoi/vi
8PeKNQQF1EFxzO6ajIWWrOpwtnLOG9OICW+0Ql7GKUNGsn6rluMAhWotevTT
9KnjmnXaI41u9iHlaQaa2jbpQfVNPMKa7kddIbTfDWsXIC0ppYP+1fttP5fl
TlsFJc6hshc7nAgko2eudRJpN06OCyV0i+sM57pRQr8FESCEBHo0xEL+s4/j
lUAiSwZqQUxl2uKIFXssIkBd8nSKX8h/j7c9WUo4iyUjWRUduRPJXypbV+ZE
AvEVOgXfUS3GvIVl9kQkKGfgeMl6oAUkzlVHsN6vJxjsNLPMdzvvAirfmM4o
fqVmiBhLVNComGnyjaF+n+mHlyg2gChu6kizo5FbD+B8zeQyxJK7YReuVjmH
ct3VUZJqsO+Ea6aj/RQiGcIzwiz4SyJu98XWsl2u8UoiBTDUhuEmfby3AwOv
/hEySkzR6xD4ihrf4FVO/qc+7xohO5uDwLpeUft+0W+bwvYbj5/welCRqjqk
nKT7oMcxIDR+nirSUnYiC9026rzBeZbLqBUT35nY27o3EAwNsoFt1GfU3CeN
uomyjNmFRxuVMFnsXp/9x+cV+Kkbk+JZFY+3EAN5weM21zxjM9S0fPsQh9Xj
Ccibty0K/TJFt47yj5g8XpToq1E1PFKPp0zV1OnkiyGeyrZFWLnxDJbabrYH
tnjcr/d2mqlKjvGRP3Eo1PYoqJKpPL/l4P+bkEtlMmjjeyMz1TQHXsuF4WBb
4zew/qwWIkGpC7IsWpKVNbEHflbUNL5eCN4DenFYUXAvPqtixFTIZnXbnEZ8
luob9gorEtaZnaaETzU/HCi9ekHzBEQUNswcRMwjYeOEIhv6mGxCXbqUELp+
b9SjoJtuh3EdCbJwFWAsyJSI4xrsxHx3sk/WC52y8SfcmLCFPW+217KYLtdd
N/KavgkCiuhD5eIsrYxVhtYKsDUk0p1oEVBC4V83pqEUsysmTuQQjw1H26hm
czaGvY4JmrGupVzANRdlYbwXj7IpG0gi/sdQe9ycOUsOVgTDJXyTmcaCs8/v
TclQaEzw+u9PLd5aFc0bGCnjaCr+w5WZQ3EAnr5awGhgUgAzsoM7P8tSWcUC
/G9dvTY0NayK8gRr3RDzkB9sdU0ZFuffgsDbj9g6Ct1jah6xP1euOisTSfCv
2dyjk56rQtxGPpsk6D20Ss7MGxOqB6YYsOQk71e11aVgswqi46T9su5Jwr0L
0HxF63WwTsZWn0xeT+CMzH+o02czqDIudQ/9xvVKpwwRkKhtlGYdaJrujxUy
+gT3gxp4+18jzFsn/EuKXgXYjl22rRWA1qZ6wtZS59nCnCWnBvsOwueASUK9
xHMLcHZuBNN4+H1DtzN9Dw8hJfD4WCp6qcaXV+edT6Bopn/tZTXDyXA0crUx
xO7PUnxX+elyGHl35jHSxhEub4Xe328a3V4zRpNQW8n9Z0jUgmVlSqxiEmTo
ycf3B8v7lXS7zDqfiiHBu9CQ/kmL0/tf4HgSNvaTWMA/CVgzx20toz9VCJjy
U+BLG2cvL6waWZYO6D9HpnzjAMNkmx+Xmn6ZBYYqtb4UphbTrOlsK73Z3VIS
HcN9IhResBLoikItUrqKSmdZsqKBXxbpE8FKYWRyFHv+Fhhzf3DTHtExbmMT
eHbjleEGyijGJrIP9IzQjOJAGH7M7VNWwKaKLfDcC9klf+HTRaV0In9CFLxo
k6mg5QEG1rB88/VCXYAvdgXq8sgXepOu8k8Q9gmaQLhj9IpCIbHaNUSpafaR
yjISB30X6CvG+N1Y2OKd32IZ90xxONkR73OUriqTSBf/dihXxmyqvL9zYrAP
xsiWoJFVld/B9gGhwIifBqMgK79OLqpXPyoL4JL5MPFZWDtPZoVHPJ/Z6yNW
Nl05AxWbSfR70MLTWoxRK+W611qlYIVRmK5p5U9pnY8wPdJowQM8dSrvPIl9
3EzeQ+N7Kqg/sEwMHoRq0aIVZ66amYTpanSAjuw8LJMSFxojhbbXCFWh2NhE
MvZchlf6EhxGfgxst6fuB6Bi75600Cv8Q+dsxugO+CkN1CwKbo2/VCo4Jt9Y
A6gQY1Xe3hs6tCHnHymmZqY2IP2GX/ZioG0PrMDprFCDjbv2jGbaFE/0z9pC
P24yzf12UpF7SihxMjHeplCzfFQJlRRZqZfh4N7eJAhc4R1w3yUpDhXsrN8g
VSBmcR/N1r8tJqWblWQlHgah+tUP8hELVyRCD9n1iGu5ke1HF9w8JknQ4LSA
F80+t/c0fFDJqOpLUWaBs0vuxA9TrNqyWwF7wdUjh/pqKZnDz3xQZLnNBYbx
UpXliRemkIZ+A3P4B0ot01ATnBpi8IpJSO6LIgviueJ+cLhoECMgcAKJgkEs
fk1tdyyu0c+J7fYRt+tCuy7mp+35S2u6zwoCzG2aOHgUgga++fH9MnXuIJxZ
bGjieWowabdNyA/MGXHVW2u7FIbF6R3f0WrYR+z4zaOOt0Oc+ohFyydsWQc7
dxTOVLKL+n6pC18lkM6Z3NtsnEpk+EH96zU+QSyizCY6Na95BZa6gv7eyOUL
0BaK9MXliAgkgpPX6/+YORJL3ZoBZ1JuHw42prhKTEtf0B/OiEEWeDzqTxbw
VrTfFf5FsRNMR8wKJK7mrjjC4zMWfu5RbOCQyWjwN2DBzvndib8LLgSmlzDI
zICT2pX9qtHqz4eII/urBjlTNY93+XHLsMXXLDttmkjeS1PGRDdn21yB+6/W
jCyZvGYxP5LrTAc7Jc5NNUNUYIATEXdiATajaMGWTBbD/7b6+QuOp0XUZyKQ
9DX1Kk0NXzlrqsLlvyMf2Y5MCgGHV0Ic4zQugoRdvF9elOKKWByNFExsl3hP
AKq6Ujy+TqW/mlH4gO0ttfCSMmB4actLAcR3qTUs8RypmAi1Vv6bPCUjBuQf
UXbyWMD/P4v0LIC9wjzkd3Jp7WMX04E6Rttw8c4L4beg0LxaHa3UTr8ZQmUp
saSPScjv0IskWu3Iey8SUtMvMTqo9C3XcttKQHy6pRrkJMJZhia/cuBhexLq
wOIs4wVRjNUQNUxSkzBR2UOLOsr+EsGXZSuOwuotruVz49wegofIHEu3MXUv
2IYL5CSzvNtVP9jNDClZInUSVhGgHloaGOsxMyy0yua99x9JVi+1hGorqGcj
blQNblysP/+AemHqGS0fE2bHhIDD2OwlRLV9lHERwxAxlDpHVPQqebs6iuPl
ak2R7peAAyP9u5FNU2FaYpxi2LtzynHR3d1lKXJONWHMsfb7/IrYKdmgK16G
WnunShMmoPIYJbVX6iLsxFH4n+DXU7AOTALO7oOIR9oSJ8ZCXd4EbKIZk9c7
DvLsEFXvsk4lknOH1Y+og44VucmnG8ij0AOwIAV3aB+k1/kn0DvVFPIHWrZo
GTWzWloK1p8Kfq4Yw66boz5qYb8D4gey9t8sSjxDgtOqHm5acMewt4NuX8RU
YF/aZ+8+FeBn4ewG0pfcbh2whnK7nx8pHGlvqV6IZrdNWlVWyQRg7+b/svHQ
h3DrDAMZmhf+azdXOrXFGYfUeHwj3zaxe1p2bDtHJ+UDp8hH4xI543kVKLQl
dEMyl2inTgZQP1MO5aOEBRkIlavPoh6E85C3KQVoZggNyhfuEYezHMb9YFNc
t0RTBfULV0REquZpDjXXwuR1B50IiBI+O/fPpM13LXdaaNt0dDrQqAWYp7st
NFv8U3Um9QmDH62DCByHJYKMA6VDKZcSktHm7lnjSKGxtDf9JC2L+eQBHI0f
NsF/xqbrJ+ZcG8v8ovuaMfUqzjD+KRMg7hYyaaskPQHBkwE7rkK+K97Y50+X
rl2JJT4uT9JIpHkQ82xm0vjNs+WriFyV+ijsp1WXsAq/NnbjgOPqqCciHf7Y
ifimTx2Tmt4sBD2JJVB64nADvqOJsio8F/We8lxCU5ZYjdhxvCNfLx5jY4M4
GnNq8fp6LMbDpFtgHjDDWp9/qxB75eSZoTlxJGUCIOc5rt2s86qZ9U5bmSqR
Vkwn6fpB+984RxDYWirejuzqKhPZvJfjpcsq6Ao6o7nMn29CD8NuI5xhJtU+
b6G374rDH1OPxR5I7pfJhrMGgQJTFSkXuLUEqS6bIqjLwqDQUMlYlONVkNOi
z0G2EI+anslSJ0R+2UyGlb4fPyphjpw1rqgVqdFKzaFLp1Op+Kt6r6CY6cK5
t+Z6/5n29kf37Vz1DQR69nc9M8duJqcvzFPbUZpxpKf0nxdRBLYogi5K3CZm
796vX3dZAD5LKP03SE4HEbxjRztA2UucP6kjgI/t3j255AzbwMZ3MGIvmrUt
50cITgIbx6moJeytNGZA6VQILGIZLaYBkAW0mEe1XIwZ20yrQqZeytNuDlWP
ESSFyJsUSUmQcIcil9SmC1YLmx0ItL8qvb46FVs5OdN/57fuXXFvkWxE4bRV
/mrukiRucyERfzygY67FEuvpWyiMsvl988IROg01DplhumAFVbJbX2R9reth
SheXBlOn4E/YctVI8l/x2CKBVwdq5QjW3DBk5Ez9kcA/Eyn/my9Xl1MbBz0q
ww2z2TJt8fBRwGxWv5OD41CPuDcxG3rVUa9jEnMobDY5DxfteGcgB3d+1rKD
fH2m8I3PDAF2vFPt7Y7IDYoKif0yBqhrUiVCZhC2UvgzPJNTmsQ07FTKkzNa
zD2s25unr9CN37e6U7kds2AxLmYygXUGf80/z9/GODbhrFRnrduCWvOAk5m/
RWdKuoyziohFCqcYNiMfeqf1wIq/ZHl7slK4d7sEUh8bUFKZqCJbcniKpD8/
oMVI+0NHGyJ2mhO03mDF6HRhkXn+3QVDSUvcUOb5xO6QDdSeCV6q1MarQv4G
xYYsEOT13nlop7UvkKJTrSqWmEP4kwpxAC70WSFTZQWj79YvegpIW9ch4qSS
ktVJQoXRK84sH81xRjjOx0LK57a4TFCgQVxMxD2rDmS8npJ0ZBrJQb9e9yJ6
q8SglBoblMDprtON02N+CcaZGfohpRPTZ8Jd1vtFX+buwLkNVbA2LPkoMFlN
z3iRewDPO0WMXFIpEPYePqXTqgx8L4hFUf37pBemCGfq83DmpQV+Y1FV5236
gWWXG4fMso+LDbyNBcQy9FsCwKuEe6xH3vhHMwF+jJsa0zrBH4oL6Gqf2hjQ
GE3Fea9DLgi/LYgW6hwnOee2A0sy5a22ai+FJWsZJFNJOJseKnET8pUpJooA
VDuDySd3JkOYtb2fO/MHxhvRcWU/m5luZnMZltEDe5WkP1ZiwEq7EKGsMnpx
9QNORA2Oawxt5Jw7oLwd01f37Nts3si0wuhgHUfdFdf6UG+ZZKYK++Aw1VMs
yBGOmiXgJPxAp+ghLFlXn18LEw03+hpFvRKI8p6VvCjLfff64EYfRE82VRNw
ifm5lLTmncGf5zhkVqzCavYYzlrLXwupXZWNd3ypY3beS/Dz2KEYvd1fNmp8
0FLjTQXXoRwHKl0eDC3bPCEgCK/7oiqT2G9Ybfj8tw6u2tuZ/MaZ/sifMley
azXpyRxF9vjck8H6+DAc9vZ223kuO7DszEpQogJmH2SQ9/M8drPlXykUUOPj
2uS855n1g1A308Q5MvUSA/FUFNoCA6arFfow4pF9YGLOJTAie7+XEyPLwY1M
2Ll3KhG0FkCLRdaDMYav39n8aRpDfFO2HwqPwJecNC2Cc98GN7gHJunj1tul
YXZ10yCcR16Kah1gXi+JmUUp/ct7pvl6oDSoORQ0/VOFZcs1ynyzMlCIdqTg
C/G2NexbzNTg/o+fmxgblhSUwAcwW1jUTqrsqCXbzF3mCylLAToW3K8YNNPe
WpeCRNrLT9r+2gTvCfv9y0k6HNWR1XPoAv0YG69L+C30ZHew9seig6Ed157v
D74Bl6ZhvM7o5SuwfFzXRLlnCkHOsazKP6/GGk1RfE6ouFb51dLBtGd2CN4a
+5EHTa2/DsumtNFFHM8MRxY1R4Bb4f2Ij0N44UQVsAiqXVDuAk4LZcaBjuGF
KfSSkXGgh72wota+1Pcpy6Up8s2s568ujukqUYwYxd+H3NjL7yzsL8tI3u58
WWvuKKmjedJjvmn8p6CIG2z/hlnqJpW+Py3AqxzHoS2tl2CQ9Gv1Ej/Z/QAw
byd57BUh2Lu9aKZZn6IzDCPn7njejlJ57JZHpSvODMRZwCt2Fqtsnk4j9qmb
zcknBkvd7iDxKUi7q9o9HWUldSRMjVM+11kPNCMd13n/pKjQ9yjxEdFezLlC
zPiS7apLSQ+/csvQtkC8a5jGaYT0Q/q4YWd97+4/wwPQW/JAE1aDV/HnmKQ+
cp3G4MSPOROBd27zn42H3sLy75ImuZ2nOW/mfhHlAhj/NDZ+7/sdK+JVptDD
67uDZXnunTaAz5mC34sWB0DXkvYp57stY8naXrcsS+4Diy+Xsr6HdQcQJNtR
lW+C/lboEDuzeywWJmEV5jkAnu2T73Jyys/2pajjZUzgzRMlzxttfD0Qe2Ta
46m38UjGfszcVw0999dtQeQbeCu4lK8IrzLyoYHiDGOyCabJuKyqSv5Q5Wwf
QORKFCHRdjhGJ1r7AvcniyncpabIYVcGQBAoNxYzgmPSEOF5oggxvHf7nKvg
T9rHZddF8n1ZmW+crlhC3rYXOvLCZ6p7Rquh/qhs9a06v0HLJhxpwCWdU/xb
BylwHWJSrykKAoH8h7GmTzOnd/JfJFrtJ+3wX05aE16mQfw+oAn0J9Z9sr5L
LxOK8yu3KEVqjDWcFZXSiESUleMviepCq6dtxAeSSBmoh8YqA1qE8Kpi/+l9
LZBZA7To5qL9hVcJWoxFGXnpotkYYvtUj934vKlNcevxtgddrq+hc3QnTrPb
IshSgFqk/rj6pGJD5xnbJOa+IJB6epoIe4tT5qkNP/BeK8QLmvNhNLRRUV2d
Uf7AcJQOWD4/U7SjDXKN+DK6qeZ58sym+V6NDLPTsnsaiyu7XdFCq95QMjrN
IH0ZN2GWHJ1Qvnu3yrHxSXqcRZbk1+HfnkDja7wo4yIEjVbusGDeVzfPgldG
7Ho8GBIx3Md/vN6KPZqz9c894awsoYcrQDXtkmulrjVSupcoTwuPIa2U40Wm
KOs9OqlH4Xikl8DeySpCTDlpcGT9qV35QbpzoC1vBU7SV1KIgDkcGRQFyJOF
955ofaULNttJDh0clDSjTqczrCWhDkyBDXxergpC/hdiOhj/jESgn8diIuMR
OTVg7DANHbOAjA/XvmYZ/xpMq1z2YPwHyVEyvAWRxMGJbD/KEAm88lqWhub5
5liu6NzykWXZH7R/kEA98N3cjGTC5x4pgyt9ITTybJMCGq+nenJ9ea3Q5OCI
Y6Y0DnwZZwwEKLnCZQTUSl7A6qufSQ3Se1sn+UoNHdJ2MT7GG3dspGWdJMzx
68M8lV0atNIERgGJxsrpvmkaWy9E6KV2czGwJzdmEjFWaKxntyvzJ2lk0K8q
wGOKy4etXNn2ERw2mBwIXkJYqmtVGfFZLZgqSN3ABxO6ge0bnbuCAbVDnG2Q
0MIkjEKS5pfuH3s5D72G+tYkw38sPOKl1/Qo11Ma7OyYmHe5ATfinJyrIW4C
etxcxX0CzK0j7n23JC+FC4JQ4DuWi1PvEUTH+pXs1VubsEec7FQwbIIE54wI
ZQOwBgXpEg2bIA1az8FkzFzhElsJsi4PkRJ9eQbDimbNM+q9gbzH+xhxASBr
ceOO+/pab1/j3yzApOcEJ2BP9ptOzpWGQeQr/EDltHj2uFeWVsZ2gdCJTT+F
Gkjk4X8nnPsbM/V1I0a0acnIVVMXs/xE71y8ys+dv12hAPJRuGVcqwElkrux
jkjgYplhGDr928Sq3TM+U14vDqfODug7BMILHzDMNwV9AuTi+9PWw8LrAy+r
g4pcqhKdHdEPD5Ezpqn0hLHB0o+gWLhUsUZ+MZ4jZHwgChRUnzRkd6UhHQDU
cx3VkcoZhMtqyUwha7x6+o2mBc/x/bazesPYOOBt9kiKNEx/n2e/rcqID5ml
kOwWlr5Y4t5y2aSXeW4isLnJPu93BatvqYpYxbeTtjkQ4n5fmo41DT6Pjxt4
xMclU9fTCFwDI5qMNZ5qdGu2vbmqvRaHWeXHVbebYGwAyG9xXR9gfXfIGKlC
Q3mFRtnMET871SBznDB8p1rCyzxDNgIGwl9hofQBWWDNFbsloxYL6xjSjmDH
Q5dfPRgYzK2L42NQ23mZVbwrCKmq6aM/dLfKjKaq9NfXf7w567XIvvQHbdJK
umj3AVSk72jOxgN44j/OEoiUAUHRRl20ikubxO5BbWqqK/L6uZ4+6AqMY63m
+CrCisxXYyeHh5YU4axqDzsDdGhAG3sJxEreAm/drjmaT0SxDv3CklKsz2Br
hVe/8S04Ev2+WTIPfECsQ0M2pu9SxxmaIuB3lrXOu2N53dP2pH0LIQH0I27m
et3ZwqAcBVadwIoMTRTAQGMYyHfHeMtU6SQb3UMyybAgRe5YjecsZuSLktM3
Ek98ZlnjJMB4mK2EKFX8g8CM2X2Y4TJU7HLLT7KmzHuoNkMRY4g7Q4fdMXxW
Mpdm4XjbJO6lsedF6JNxD+JFXTbF6i8o4FUbqFqzqVCM0R0NLsAb8UKqcAHW
Rx2sg+NWg/t9YWHR/0PoKe9hqG8/75l3TUPHFOalv0My21nDMhK7X8ekDAuW
PegRnt7DbYeqm4dTX736ZAkCj52aytrMT3Ry/tw2EQGzr9cRngDFOM7QpJG9
yNGNecSsyzIa5GBGJoz9Zq3/8BZHvvxP4fjJjdvEK826yUorbfzHn2H/8qIc
F7AUbXFKKXUKJAurlz6m/+YcIoDZ1KhcziI5FICq8Vhcuc3XHGDXVaZFQDij
7dPseW5nYljg7ds7ZZdp4by7Y3IT5b0DQzTxm+/6iFHmql6NIJ+vK/2BIwH4
WGK58DyTMTg99LVx+xI7wTN4Xy9CuYlwuofEspbb+EzrWnAnfKXd0Lrx2MKK
mn2Vn2ae8aZvpAIwjPey+S8yrDVb5nljscxWgl3lw0oOioEXWi7LDwooTXiJ
6eu5soSQ/tPrkfpc5Anvnv9C2fWTurmm+CuRXdfx4bZOWx/w5Oac5dy2MQx7
4Ew4ok5j0i8RAhI9GMPl7vSs7/ytSWrJaZKtr1l4/gbxLWSkjIvkksWAe/vo
AEfjVzMzA3XvcP/4OaKcOWeD4oRTlRwahemS3VG1837BxX9GkmOopC43gR/l
SHWsw8G0iULScuGLMLCVPYzGfXzbHnhWfdKPkPykoxfIfqW6ATENU3Z6FtAt
DhWVzB/pcVfe2QmFj4cLvth5X9u+jV6IvfsaXXjhYjjAGghovnmvsOm5EWbQ
EaA9zkspAKGWx2g0c4Bpz1zNA9UlSQFkt33GI4NWN9WzJ57lovYKCyw35Gp4
H67LoNGuHG7Yg6kIuOmFH4wai6eMZ+Ts299NLKI2hsgrAFjKGH8TD3J9K4/G
qy1JtdgnCuSh/hDALMb2TyaOz+fASwOLFcoQooUKJsa1CtOrPZ0R819UdcL+
HECQLFh7r+e8S/FW66np8D+oYpTG1or17cT9FXOZbWOs9wRUUbQHdWkgNqMv
iS6S3jHQKKT3zGDVsWzVzLt3h2A19qn7LZJnTn30uszcttJjQtDEL2z12NnZ
QNKRoCj8CAQOd+fYEyfFs33jDOy1FzYgUHZIkJoFMPsTe5fcvqkCB6E8KNNg
G+eYvMVuXBKFBmUj+FRApWgIWFp8wh3dqfl3rTsGQo+qiB0JN9Ve/0e6ALyN
Q+1A6+ugWyFOABfkrZMZAJ2LvEdcExlojloa/5EjotLHDgjsYm8s9RYIuWjj
6tzPhWXnOXuk0FSaWekGX9DngR1vloKyau5kzbXb6SofO8NTGW60pNISJqV9
EA9T3CRcondBni+pVK9qfaDT1Chxtu+sXnqAOdSA+6WGqhOSyRJwFXnRta30
2lscVZ/7Zw3Vf1zoS4d7gqEmsX9R4QzVOy2GaBvGKJgigZthYXq9++O0mcpP
hkO/RiwY2raKYpCR6UQ7XMKWWHQjc1n1oUuH2KjcJ/53iBRynkvSfefa+xnO
ypSxwpsY4acUZb7H/u1dSHhrYGeqdGlQddalbpOM8iCuNvfx7L3MSt40XAXE
eMdYIiW5Kq/WsSw6M0vwGSM1Pn0SU3B8YW9Q/NtShZJ2LdlZ/dsU6i7b4S1x
CLPEK4L/YVY2Evftg6k9gLbYPenhIxoeaETVFS94eWJxBxr68vjozZcgi8dr
JfH6ylHxWCu1OPROc8VCy6lRUcEf4l1L2XCPcOS4UBly2Tm7+Whn4dgtcx6/
spys1TZQkmUDlhRKil/GIFI7dbZY2T1OF07S5WtBHf5NDYh9zPx+GdlyAMNh
tanzqhwlzYuTdrUHCgT/b2mxaMqVSGV1Ol63ag/GbrhHcwfPOBnNENgF3Cmt
XAlooPX654NmeU+QxNWZf4ZJD+lRo+RifYVFmd9913mHcgIO9zTl0WoCMWwx
bTY1iwNTd9aLGaHXyrIyvLmpGj+wU6w0yyre4NYfr7OF5IGtaj5V2Ob9YieH
84hq4RD2Ew0QyMe3XVRtJGUIeVqptJFVGkI8c1J0LFyw9Fv8oUvg1hHs/8Q2
y9wDNvM+7LqDNDwtluoXEGgQ8IhZlFYQl0mkWrNOYmlCYGyLVSmEtuQ7wqWx
Mdg475Evp4w/hKg6vWAy5tntZfpRSETJPJeNFshselQddFkwxveW19XCToIb
Mst8ph1K0TgIuBGI53/oaXBssa/HsHLSDQRwwRGCqCYivpCe4TA2Uu3u9fwu
aYLPw5BOgHH5DT2ILkHP22X02oQpQ3kxarAILyRQtSCXVPMfEBH4sv9nZLaw
05dUJAcL/lScezAtWNHSOXsJH33BcYdHHNR1YDlerhS56qLqQMAkuYcI9R2r
mekOpKlP6JQMqT2i+Yl/yZua2jdrNLek6nyHoXn9RP8lRpBGk9PkC4XGI4SW
RquQjmWGIEmJqHfZSP48mR+L53intV0MNUUl8ixi9t4u8Nzl5CCDkvJQfUN2
27t+8jcBemeOXtIbFl9LpRlWgFy6n+11ZBNbjeoYfy4c5BEx/jDj9nPA6qhu
B5O8GoRdrRg4PfvCM+9RXgKicwDIPrQX3YQmY+Yqj7WnIr4FdZDtvn2S+k4V
08TueuNDp/bFoPkjmmGPrh4GjhmVxUVO2erJLczuiHYmy/01QFK93+8t7XhU
FED4jnUdUdFmhS/ybtyub74zPeZ+3xgcW/wTkeOOU3TOLcrwrzb6Sisp3v6j
QtTvvSDM0uptSQrDAIqoZNLSXSYsPMBBSuafGzvj9QOqgqSAEgsCU/3I2DCz
mmKT2pcX5Ec16qxauqhOp3MwMnvTNVPPpzKlay8txgnf/9rqnjL2hoq5bZlR
WUvxJ20J2oinstDQJkzdpHCDdZ4Dn6eUMWof8dBzbqJovxjEHQiOnTCLOc7f
csSpm9s5bVovCkGdZNsFNOLvzMd7hdAM4nwMaN6aSr9hq+ZRdQmxwQnHZUC3
sPIu4BiI4rEEhsGwnZQjjDxOhtrSsGk8GnLZVlFdfhIIcmiT+HuSOIscokwN
58HPlY8IPKZK0Y0luEa2hzisjFXGzUaqWpFuUISKxRhA203IsmU7V3BewAYh
fNK656omF8FbXBTcGf5ZmWlOIgt4kjpQsk99mgDl/tObjTT13IoxzhvoxUSJ
97YzXaHZVfJs6sS7GjecFDoyCv9v63huBv+x6YNqQT14CCGPfFo4Myn+c1xh
Bvl2P0EJDDkEl2lTLdMfVjcCXG13gGTjhbsTV0a6DXvaJYTkRpHgkGjoI1LE
VGRjNyR0q5VdRq/AbS53DROsLJN96gf/Le1jGUk5PusOUtA96CGTDAV51pXO
tFhoOPYuV5OXHa3QldqwwXu8pOvxHRX/BPudg0LbBfqlZCywtYm9XCu73Qxk
OJuq9/FNt9ai35vFXe+rtD4/zxIEfDZykK5IyrEMu53QEtdFa9w1RsH4jXrn
BRDcRMXmnbUGHNI495kBNsCTC2Zr8Kq3hG9V8X2qANqCjOHzoFcJpJoHPTdc
1E2QeqT2ghnJ9JsFuVytIstNdq+CY+BIgABRF5DL6JdfpHxpGplbXVUe0v3K
iHB0evuuN7WbusyWaEjazkB6OHFvjB5J22Q2D8RhKwwdjJLCmQDX4Cfd0VRH
38pUeJYXM2rXhUbrzX0Nx7ryyLUbM0hyQuXLDilImlntz6XVPZ/51S2akoSP
z+RKSxsZFmXfJCso4zRaeprub+xBd5aZ4z3Nd7rIkIfs7Q0yBflVVohNm+Pm
b+TqEuuJxE2D0niHVgIVIFv2lcAwYq3op+gK6PBp/eJwq1ngsDfh/lic3UqI
SiqjVxPy4UyEDvpYPsovF7XrohcT4WLitbrgx8ErcZ30OdsnPgf5HiM3vHjP
3Lwm006lB8UrBmxiE6WfkEDOFW1F5mPiS75sPdYD0tgzIKe5K13l0psQPvgp
UI+78e/kgB9kmfcnw0JOLe3AdrpbYK2wWWn0p5AmBxG/Fc5EiVNMYScjZmf1
h/MTYxE0Ym6I7XomfkjtW0/7IxMNlTTmQF5cDTO1dyE3dJbOU5bwRWIHJGC4
vLOvaQg1QfiQGdr6R3i2nyrff3CBc9dC/UOt5vpjU4j7a3PXwOY+oBsZweUZ
23Hwl1spE3nqJAdt6q3rCwOa8Pk+pDQI9Y+KG9tqQHPKABgt2hXffKN81y0S
m3Db2SwiiEiakZYKHh/1zI7pCRfnwdXUeRxgpHqQ598OlgBOMZ0t9C632qmz
rMIgLzc9ARtuMCDP29ubTdSS0lezTmqU0HtRuQAYDn9mNs+QDg4Bxjq+XKl2
sX2uoIlhmjpuf1xfr8cZzCGo9Wr8OlSJ0JplCeympJwLq/1SIkuG/wI/wUTy
eG/zUNRQkgZD5+RrZdkGKoiEeBiG6E/sAiyGBO2Knvrnl/IEb+nkKZh4w185
5rvLn2zLK34BEoYJf7fiW8BoYYyMcZo6ZZuAiaKDM8PcgERzL4rcYvczMPWW
Eg0Ia2JznQv9FyQ9Jn7wIq5w1AX61jDExSwClwQvd7EkaGzso+DLLd5JfAgu
fPpbdYHzs2hTs1APaAv+4xBL3dnQULkxfvKmEQZUOHZ7iAJiQJ42Bmd51QUF
1+jxIYI0oUApuU3U5m90GZnsxd2aeshYcQTEFCQRifxwSj+jv6iHBrk0/WRA
JP92yWLinZOVnsgyC+DDDoL8xlTRgnG2U1ct+XadR0E+/wApAWqpEpdUXhui
JrLuno3hD/U2EBq0LO6msoRZ4uIoqGiduuM/VrDGW2D2HuzeN8WcKZXWr6/f
pvvQeGYUv7ckFOF1SwIFpDjzia3VCt+DIocSFI7p7/6Nl6yYnzPKGA76QgfR
xGsIeUdve3gu6wk6VlEZvdobE4YOiKk5AmWaxPIAl2feAjwmydLOt2FvQ3TY
mdWBm+/H5KvFnCxl/B5TOa+SJvhpMep7JtffwB+JXAjdgRmXDE4dXui+eiaz
ocyz62/DqRro42bvidAHpfXBOgJkYH0/YFx8/rBdmclRgY8QoDoTSwfTViL6
Pa0ghOiov0FVsuDK0ec2aiL1rizC8A2wc7GcYAtkdImhLn/avg45Jbd3JE/D
FCNSNK2/GT+OVTuAcUGNDGt+o5MXKxxFVCB+TWrwak60aVyFRiNWxnzS+Yl9
PDepOwahXhj32NaxYnXdeOKi0r9DwB0Q5sUh3NQtSIM6UTg9bUuFSuGrctdO
VvNBuATD0vzedCeOgOgV3txm4OFK3EatssiUDPzHAsVbPcKxUfMnkRFPGO/F
r+EURrplhwCUNVkZP8wS+wVxraNw64xBoGVhPVvERy0Wx7W+FmHZBeTLNPVK
2tv1m1/++aUfhQR3ThLP0j3Yv/euvgwMV9Nf5isCpDY/rC+i4PhthgMNUAFm
p0E0y1pA8IRIUldeOGXvr+FaXPKNUQuLLzDbrY39d3PQ7jFJtQ2cpwBdikOr
spntrMSpCovpUKgKpMsC0a1QAgePZ1/3vltFtjONiPMKSAB2Kn2KOcRS/XA3
vOE/btGaWuK7nITf0k/bP8Djm9df6E/XkYZ7Fnyj4zypK0eAeeFaLgFArAwI
GQ5MHCtTlrUqfubxMexYtPUgA3A4uk79y8W1JijITxsg738gjZuGWpcTyIRc
9A68tBdegsXLh7Pxv2bOb2h0txN5I26eUafNhGwLMIQ82TO09Ko13ttBnBCp
HuAE83JHRpuyq8dGzQU2tFyhWQS/Ye0Jsq/lrtj+N5d24rrf/ZtYia5wAv12
Edzkx9ZFH2d5FEw8TwKBAguLJYKavnIEB7XPySmFmvQVIecbrmqFGpRNBGwl
rszzqLxetuRzm64L8AfkS1ubImoddi9H7s+DDfyPn+73PHQxu68qU0BvQ0Hy
DUpKt7e244s3B3Tai2qkmQVVX+sj2tcnHHZ9Z8JbFwoy1evFbat4FUTE8NTK
jqvVuhljR9AS4AK4j8SLbRgCKwXXVBoFJMWqQ/2Nyi8blvJ6mNB/w5S34bwW
Nk3IG/QopSY3YB1agOmrDl+GmptW+O1eVaA3FlqMYQNcyYBUbsVTuA+BvOZW
BNhGKovN8dA4zRcjvFFOfbk8POmvM2XM2Kht4ZR7QYgycHla7rrdxBFq9kHO
qwfhVHKmoE1+ervDsx9b4n7A1zZFmartFwZtev4GmuhnRh10FtRlhIWAOaes
IiTUWP7dQkSurPPZI6MdVMsF7OdyW3e1wyISaYK+P/cLqaSEW/S2w1/Qf29O
HRjLBpry6Z8cEdHFT9vtgyI8+yjA3DrSQndD+KXJ6UbrS/X9P8wxvWNPauOh
FQcWDG6mPK9864HsSJKdmhuaCV7M6I0PUGgdQ5bHDXylzalAbCyNhVENwmVN
ZIxjv89DykTijs7g/ht0WH8wfAvWmsUx2kHZQrWks7H7lxzYhXMfLp3z/h5v
7z2uY53UYwGCah0GmNdov9oLbxHM27qxp0B32DYdpHDRXK9g7JaZVoCQ/lIr
/M6VuBnvm32N2a5DsrNFT/b8WyxUiflTO078ZkwyvsodDg9wiyuotfAUTsJ1
17RSpNpy/h6aHlYMmgQYi3GjE57MrMzXlhmNBmeHePwUJaxtUxentAYLLi2K
hrmA/+fDTrEnnUbnsBLWMDbCHoAtdDmKUeAgqAoWdjv7W1pz23K7tjJeamGm
KHdYUrx92Kdcc8Y5MzNOGFc9DOXWEsQxqrF0AfICfnl9vZfnZXLwD/Fv8MrT
bHHAjz1p4JBOy+QYgH1KZITVK7G2tnyMjPE6wn++ROKs8XedEzQK16muS++C
fb0d7PW13wLu2KadaCJa3FgIBUXh+x7XuMUQs+V4wAPwTxcgYzgh6Un23iXT
f1DSNc/icjjVhFLrnC+UXqkDKhwKUTajC4rj9cHdXgcbzQZPv9oxokrBEyoJ
WXW0HrDYlV8d8d8zGdQdkgdxtvN1WvwdrmX6N+PxsOiiOeEfoZiEC5BC+vqY
JkIhwoo4caKfBMHGTcIUoZmVR/K/YHtbZJFYQZFqupN5e8OzQC2ng2Btqqvr
XJJoq/MjYm+nkQFWC2eZP5MnbIC5I+5irxePyHQWyZBEMaFgjScXeUJVAHGW
AvelR8nPCpvB7wpu0ixcDszJE5RS2mSG8LeCmfOhmhdUg3wlsIY7uBJB3jB1
WYZtVFIb/UoWuzGeGI1YhdhnyfpmfmfErtwydjnHFFghL3J2D6vH9SOeK4Y1
z5/wFkwm6iRpzLvQxwh06CpoOTnnpbCzFA5TZRqKz0HCEdutoaUsVgrK2veA
2Gq7Uski4r5BIJt9wR85fcCWkKmt31BVQZLuSHeaK8nEGwFcMYsNQBgysRZW
nbD5bce0tZ7XiHLTky4ZHMt5TPLhH/5X+5F7kRmrWAsollMx6sqxrBm73Lh5
pKGHM71b3cGHvt8hEMlH6NkI0wZ3Q3DoBsaccfP2U69Od61bqsAo1EJyLtSI
xkK9pnRMv/ptgC1FoAHzEMEdMrr5ezac8wEJ+8pcTOuwq7A03ElejS0KjXiG
1rHVx3FYstW/1t5WbfiqAwwNLJgA8cTqNzm2kd3Gwp5+8D2dvuNT8pqOPoGh
ORiGvENMqZp6KS1j5jtZehBzBkxhXkQ2VZ6PvOVjUCTqdmkgTxhLscWc2aKV
Tm5GG3AhHPTUsb1LFqxx4+9ABg+BrVoqTLBOoIvQmGOAB5esT03qnmPQodqG
0J/BVabRCHhVQD+zf88qRX3tYoWe0PbUUookBaIMXNRspDm/+jXDxNBaz5Ld
lXdeDhLWV4Kei9Uco9EfEdSRTg4VdibBL9+IsK8JBbn1HW8H5ZxUPVDoV7dZ
AM4ImMRsmtGOJW9wi0tC1OSk6zVWsOf/wTkMwr4KM2mR2KgFq21f+clHaLIW
KAAu60gUC4RnQ1dFIJfVxWcZh/g6RYXvKERupMPAm3scq+RPFmMIfr4fCWbh
31gvYih/tXetwgb3K8ZMx0Sn2ADyH1ACK1FHZZ0Iw1w70hUUCTFFJBcxtIbe
edQHKNFCy+HDuYXnlVvyHiFhNf1S/acrtUdn9csZmKQMengziYMRjiflKLOR
2G+1SmK/VbOT9h9tts0Xen+BgbURIGJgu5+vhgyKdZpeurlP9nuXXU9cT+C7
G54qRLSYlFBYGi1PueJwOxAxklJ2MKHd3rLtwPYbgsunxCWLv/XF+ek7rxyP
4oBr9S8VWxs5F0ZkP3mPo9l/O3GXwWbmgFUkeOrK64sCv+HTxy4YeHHS+QpL
GkvzIcrk97512CkvcPLkCaDU/Na1iO3i7XL8skdyQJ7QXa3MwUpIq3RR78AS
ExODKESJvEHNjtz1+zJRBG11D3NH6t6+ImNotlzm0crRjHs2S0sAKn04LcMs
XVF4JSstDFp1YR4siSrs9tsyGoTSao1KvBm7qr2UKuHBe2BTVzM5ymoVKzPd
YyU1Xy6qMkbgz8ZBQKfNRc9jkLJxvJMD9DD+ESZKvA0pLArMyD78kl52jCSY
SVzy38pB+Uxb8N/stw7t0bOTDlq7eWcXEigtuhY7NWZqd4vtpRgCnUezpUWw
zk2DEzWE1/fr/1kMtu1ec6O8Z/iZ8b2pmE/xn0eN5EIICj4cH/4imbY8QaxF
cfMoDgkYPjEtKJ9LLsop6nTQrSIvE6W15+AXkpM7yvYEYZg6O2SQ6oDjRpnz
XLE8XmwipdIDnGiNLX1RTtey7CGS6EmPobKzB7YKfnxcvB4UTqV126LKDtfN
f798M2wcPTrzOx56BlayMZZ3/94xd8ZpmOTstt31h+knu/p74m1hqW3JvKiT
sCaxvhJoCoQ4pUTyE1F2uE+IHkDNB4qqyjNb1uCbwEJPJ0W/YMSBTPceLpH+
/hp02V1tJtrU2/yJt9eBo4kndy1L/Kuzc/8lJuBy/kSz+r3awvGTJgBwxX+o
eUFl2V4pHp9ZgTU6EanNdDAunb1fHtgVW0e5aM0zq5UhMLElnYZP8OwD8U0d
/aeVzpBwJKgMxKOHdWLSBkMPAd/Dabp3NHN+HQlwf77pjhUCFENDZQ5mZGOl
4Ro4igLgfAj0I6FzBZB4/0CL+K0FUcPi1GYEy+VpVzfXnudUYLQVIyV16BKe
VeawDArBzoMkAT9JYHDoUxUTteoRcMB85ATgUnCGmDwCAZPYDrP3hBiXzeXC
cGbQWz6sL1ZNxx2yBTJd/ZO9Ci3iqu+bZ1WN96CK+vXEzBCoi9SCKUDsHKuo
Ug+RqmP6J2BBkmT2wJcFFmpPmdbQJwLZjV59nPupISHu39QKUzP2alzMHKlZ
Z2TJaRzRiHiwAuL9U1JDuCIrqJf2m7qHyr2H7KsFGPI9XUuqRnS2zc6Rf8Uz
1eE3NfPibx94IdQd5UnTNbnyP1AapOJ4OJcdJDdxb19OmuKqUCkxWq+XHEa+
/JjPCv9KcE2yk8YbkdAbbUSS6S+KCPy3YprtVReEGh1LD4kKu3/zfUcLpsxx
vEu2uIixG0wg8AnOyZZMGvKvTepeKmXNXF1xDZ4O/LHpjblHiD3VdAWB9M7H
PeN9bp5zJLsk6jYtglRRxtyGixVew8eQ1811WbsB5Fx1ea4eLtOwDbbU+rkg
3bJzCldtxOe3oJIJapxsBgsCXC4MImPsRaL74yVkLXlqK8LF1RZnIXG2g3sZ
aoa1IaHvCIQ5805igsBPcFFKFO+LGiLci8Iyijp768id1vN/XnZfhzS1tMpJ
RkOH9n1H2ZskLp6wmau9uatRFBQMUE121qhXEU/v0bixN7cqOE44os+6G+nQ
RssKXxubOQ5Ioc6XYUdySlbRU2ji0pq1q38eBuIbOGqe9CCE0wUivA9cl7D9
MRT2sGYtabXKTsAyv6MoHqkq5a6oBvL/eihdeG4KIChKaV9xROJcZifD7x/1
dTU1cnARfxq2wtDWvXH0pEFb3g08ZidNUNXSN9nC5bvoC69XcJvGsJAvRbGz
GSmbGEef/vTvMpzPtG6CG7PSk4oJYe+8wW9uHEH2BOb60YRZHq9qMRVafC9O
wUQQh+/XzkX3qvuncqTiIjDX/VaS9jD8OGLqAtCijDeykomqZyO85yUkR1PW
/euiooPPDyRtkJV7kS3opUjzXjOfKak6XWFuVDNf3gfR6nde0l5Y892keKIp
VQz98Va1lCcZGvnkluqpUQpVvdAl8Pl2h6Ifyj1dxVhhcZEPeFWS61lqlB/U
lSn1OOHc9XzyJcUesR0L400uviVjXs6wBW+/leLvBhm5SJo4hO+skS+W7uji
SAVaBN92t9+l6wR3W1d2v6JbuxED8/ubxTaUgxoXk2xD4ctPRT/RrqYyHGjH
HWjfaTzy1HM9MpvpOJOCvP2UeWWnaGC/kVsFKXt1225y+PZHbocjqjaUNMsp
53fc3uujvx/TIenoET1K5Crt/eobdbFCAKphUBOHK9W1TnOHUfMCgsxqVUvN
8G1toztbKAbzgxUwau7y3+gBAnNLVNjVFSRbTgVbaG2M866HP5//bc2c2U9b
3lx9f4uUTLpp5ydcdtYWK03BmquyilhFud+KPCWfWB7luWK5EcYmOPvlKaPz
uVwAtPky4agmi/N6aLtF+5yr1X6blcoz3BJHrrNWgkc6GPsyMURyPWfHpOQn
i7US/T1TOG9IB2PyxSoeZN3Pp83/zgMcclJFmerMGCboXa56S080+Wd9kk/F
iR2Q+Q7sUQKsJyZXQUwDePaP0kZ0ao7ZFLYdLIqZlhNma2boewvjiw5tL8RW
zP9uxV+aEQLY+k0jFheJp3lknUHmgQ2jU6DOBCu49U84r/JyEsctcPEJOZam
QNian6Zd9FDSCWu4uuUlNA28jyniYvH/eSypCsGoFJg2XCI7jAyJ2wR/tC0w
DHFcmCpLT+oDt1mEQF2CbEyMCech6zHF/Vd8FyBsd1La65hPj7WsLTVsNkEK
JGpy5CI0nUW2fIols6ijd6e3XDDLPKAJ9NTw1w1OYndwzHPA/bI3Omc2ZipD
aGWEZztaZ5zU8Zu2IvXcGabppuP2r+nzMtFrcfFOxEp1r3rn3C+BSr8Em1ae
3vj39o5SKhXAn/p8Tsn6zRF23uEZ+OpDidlPPLZoUI4iURCrU95HKZ2n6UFk
ZDArLuHjk4dZssxCY6ydnREphrdgJlzjtkw3P+1HRvt0mspJr+dD2V01WXng
+Dq+4iWHkhaaBmwDSa5RfTXJuwIoL44MhHtFJ+wSS0adCfELkXClrmikYDXQ
1EyYrP5ZnAKCD3xXY4ND52Kui+qXM4B39KraeueegixPgRvNX5bIplxc6dyR
N0Htioh88zPX6JtIWgJ9wIYf4OGy4IVkJArJnt6QyHCpmzpOdbiFrun/g/Op
twx5FgAIfkGpa+dH0YxA5HJaOWwPqbaZD921E3PsgaRKu9FVseH2qOoD1AQ/
gvVIorOvUj/L9XdqQSV1ykH0Y7d9lvJ4N3j9ZEsFyQ1Wf7PPYGkhp9RBTnsm
jv5+HV4/RvppnQ1+tRciXAAiHUerZ4IJfMYCnCQAI1AUS3ttcGy/ip3AisD0
iESmdwSFf37bKXTfsbrO/SvBw0YTmQQ72AxU4ypLDSa2q2owLnz5K8cIn9fU
TWxScUVmUeloyk9jEiVxd07RCcNl+E/9ewNqxt8PZUH8mr0ImBpXf5aPMw0b
+na+zIyz3JQxx+U+YUXWlwYnMdu2GemD8+ThvlzQuGvilACtBf6r7miv0Vq2
xx54rep9VakExakp3rS5cdVZtslejjdR8eRpmPDbSUOGn9CSmUwvBgEVJs5W
vih86xWXmsElfrydrLfC8dcnfd3ZRvykUUfuUFis407KFzaz8Wg6KqtjcOy2
gDTJsSDjG4QJMx5iCrkBULL2VH9gTr1vsV/euOjKAgZY+bGEf+yjqKZsRDcv
lJhbrj2/+yN3oF5XHzvlD9RNzsgYwnKkifU4UX3x28c6JAGo5aqxBFdmsSdG
feMhjx1WwU6ZvvzkLArVkxMxPiCrsxJLt+LpaVC1v7UoANgptgKH0475ppVK
oi4Pt7gUYRdvNDw338nyDKwnCqoPhY5IxaKASAPxUD0oCgCeIpMSlQiBLM1Z
XKaDf9hv7HfFkVJPCWMIR6kdaz3iWdQU/rAgCzxZ3jwClWt+jbMoe/78j7/e
UDMbSuHdJ+egNrCcFUf87Ck6NBFJNpVvSwIv/v1l1dlw3FBTkTKXz4Qf3+pz
Bzp6zOw9gHgeCoqq1EkvywxEWp9WzDcss7W2JiuBCMuIXnCU3MmdhJxm+WU7
JFMaGlboUT9z+McpXKIgFcojrFVLDKpcrsPzk3HEp1uCUKaMDAUdinupXx91
MifmThlX+R17ei1wpM5y0X5PAxxxnTu4obH3ktJLdQTL1fox66Vvnmc4HTSR
BTQ1eBaOd5gHqs32+D/FxQuRA8pVSSUaDK4QmPCezav8CPF2UmXzez9rB/tH
BxlpoGyyJwJLVXBWp3pfrb7qFRUr3ob9ilC7k3YG9CbRgQALcf3VT07ljbMe
2lKpT+H6QkkmqgaOiyt6SMrxrAxAr65K9m1terGKpIork5YBThPE4OFFRX8E
6JhFv6IbMw0Qiybhr7ETa3YIQWkO5q2m/2hl02/8oIUHs17ai2IEMY100Gjq
OyBFAP3nAnBufBUX4JdxggyAjj5qiGmf3vw1Ki8ShoHLdyZKA/ZMXDtkyx8e
uzuWT9LArBRyrRNmAn5AJMAEQHdgB8IV03rrGHbEwbylPJIezu58kEh5WD9R
mYjrvt8Qry7DfUGaAYvGEnZjrAoAM9paurQPYVjPWw2m6p6NaU/yX7uhBGQh
SGc9PE7+ccDI2nBtjsIWOX7dYZ9gDHRo5ArI+/M6rHewgcgABLOIv5veXm6L
DIpUdP0LYvhKlpAjq6DNpBZ2hj0auXgKr0Gb05TK05U7YSj9x7HUu0G9BRqy
rUtB3/JL42+Io55vzNRjMq1X3dpXoYGYUDtqCASDTYUOLRl+APRAcGEO9NbZ
ReQYVytP4hjnx39lVogfnyLDb8o8ID1B8Q5BjpEJfg2AatvfrwZf5QxlbOWk
zy5VbnEAg9PC+B85514jawz+XZ61HqwVJajVM9vAyVUAyaOow/h23O3XdrFm
ZVLFuKxSifOmLBsaLqsdW6ZA22P0q9CtRNm2mBdt0IMqUy39+3bQUI7ktGl3
AbwTIZbbKuJxyCHxnSnVDTYlPls2qPEpiuAF+JzqkTi9vpYDT7XsDPVDIeH7
W3wI4m5R2bCM8fGbOBWHYCUAjkqualX6LPIBOHNDOC/J3u5xOQVKLsDTYY/z
ZBIx9CgrwU3FMo0ToBpWWyubV+iNtjpiqQ84Q3aHNoCLswwdM32e1i4ZafAz
RF8rxhCFS2/HeUpa08IbcRNv3tUDUvrOEfFQxA/RBVQWYM1qg7O0c92OjKCK
oWBiFM4NCmxeqEhLT/t8cpuvbdrS/liV5AAmhcZkjVFjFKcG25btS7PvbWPd
SYyxXY11R91+1k0jkuob3Qa3jRY+HRdYnYasUf6k/1CZFjoIL73XGfCwEiNT
uGxcuagweSsPeQPKCcBMfRDtuYkrKKcLwxcgEPMx1PvNOBYXGgqhRDOr3ohL
HDzPOthahAgk9naSHJc5p7sujc7i1LnZOMN9jb/IR0NT7jhUtJZE2sBmokaO
jTep12n4sRCkmfwSSO74IdjdDG7q1mC5dutriOpN/l7sZi6LsPYxB027BkaS
CzA9+VB9ycu1BqMu6NaU5U7nYmeb1V0leoOolp5m6KKUK1MIslGlKBVA3fCA
S492F2hdb8x+YzqtxdaUYfKnGhcl4bAR6mhiS2BN2alYhEiiOyTL5ksz4oJx
hTM8b+1bYjuWA1sn4VImGtsn8FNCdRQC8/TPS2Hsy06LxktMRD0IazkxJZDK
dfayhieKBNRbEBLrOudIFYWITlcIOkeF4dfRSfYAeumkfr1a6E/wyqHxUVBo
f0WM3J37UiZpF7iE4U4P96RVflM0zAcEboiFiS17AnW36hINTtUN2vtoLxug
hDmtpRpzsu9rkXx90m/9q+CN+5a+dzxUw6c2a+zCBt+AwblHJ7gG2CuaExfs
MUnjMxZCt9cVaOnNEl2RIoSdFxQcV86ZNYT0tegGIRSoZMw1RE+Vh+UMmtH5
rGNg0OoyBhyaeuDSmAeHKii/TEXs7T4C2uI+o7HUGFvOJDNN0HQIyOoZHYKn
lbIAc4pm7/x5hC+6dNXPG9Syf8UT3Ryw/aKkUwgZb9731v59D4d5oVNFKmZy
Ol76Y6BC9d0ujKZ5iFgweIvjjXhgZye5E1/AL0fQYETV7j9kpZQHv6M1Bnq/
+OnubizgNBrHVYhvdCzg6YGmJr/jnEmmLE3bVV2ne5LRRhYmo84KZ50A26yN
p80YPomO+wgge08fGyU0ZgU2Erx5/leci0EdK8fscH1UAmoC2ZzX2pBI32ym
8EmkyYv8uVvHDUrEMXQLFIdg1dcwSIcEVG7axJD5SyLqmS7HKba+iMtuJWDO
6iw0vSnTooiWezU6FeFXEgAqoEWLvLYO4/D8n1k6mxYA+cyoqTr1W1ejEObB
38cw3bxG540IL4MIrIS/9BdtR8u1KcB5UbQMvg6JII1yi0lYOrQxu+Z4NVQb
mdJUU1B8JejvVlDaLhoGEZTsQbXybr/13dhwLFrFODc5ibp5NNkGZsKL+JTx
1TG23ZKiiuE5JDfmNnGX4gYev9ZMFcjnSlAFqx9Da0uOmTeR8/JecqcFuDnj
G6R/PUYRqGZhysVQnw6ECKK3UJc9gLoFSkkincwwqznXtT0uW6ILCiIA4Gdq
NgAJVQF+fzQmKne5AoyaHlyLB1xjJjJh131rs+9lq68kJrehP0h9uP2V+yep
4VGfniEds/UyghNUWmxiAl9pm06OrmQgZOW2O6kA20dYxSofqiaf9owkTmnq
8MQeTtz8p7XB0nn/OmCWuu4gkDjZtu6P7AoqarpKsFbp1+G3t2jMTcAHSjXu
/pgEV6gclF75ObLgr8T2rW9pyCJSbs/LGfRqJJU9xQvLB5+zXRkC4p5vVNWE
n/5ZuXZ/zVSce9GNau4ZhLyXG70SrHsF5Bi/ezR1DX13BkjzeQzco2yMqLOy
mUaRuEsmNCjUh+yE3k0qq3y5PKfGjRWKrnbXGAInN+NSt6nA/dCicchR3SzO
ol8YJTladXbANUgM/KJ8vLoC5AwMuc9JLGCgAAKZtT7cNb13WHcDh3VosyPC
rLh2tbEIobrY9omUObwCbe1yLI0+brIsU0Wj0OFntHSHAj0bduvP63MO9P3S
YOT1dYYpbRftLnROxsHoc6n3Q+CDrjheu29IAjhxUDCZGFtuOInfSVFpUkS7
owv4dwHUtg/iZWERikV/7ZHbM/QzSvwzqSkyz9PfYHp+B0hqFta1SmlBAtIO
FxIpwhJAAsG7Wffiby0yYrki85/5EygTFA/fj8kmC6+WiJ6xDSGWVwdbsWCW
GBI//dez44lyD5xuwfL2cW+LnT74rsqg7OyreuV48Nu+SPdWdfPz5qVtFBJJ
1q+yW5QOgkU2HNtYwFN80DnGHBGYoQU0HoFGa2Ly3AhXYX8hNpU0trXRbdQy
sGFTaX9IsRrz5VAvIjPtTa5Sw4c4Tckt4w/Kgzir2n+lwT5BOmXxEyo7PznO
9Ixdc9EkTnsBMdxucyc9QxidUkx/Ek+Emt3boYrj/Xh4sghEgCPBbN8SMmhx
rxOKMWk73wsjHveeZErTpITdSqZQfiwD2d7T2777CJaXOF4RgypCTYXuQ3OE
c5z69+LXcNYgx5X7HfggiEd7VlNfENrj8Gfip1j8GzT7sZcm+9eT9t8IT4S2
iJQqk2oz5fwOnDqS2roW/o2lMgq5TGAXkc+2AwHOJbzHC8x+XKDcc65NCQro
5FDWT4+eo/j/LFBVgCKTd6GgbtkfwMH4WC2cA1zhx1G+i+69xlg5APr8OtGp
fx2u6D7N8MwagWqMJpZH9lC0bma1T8c4E07kqRFrTidGOahssvpnPe8AVYPw
YQq7WHVBdcm3U/DSKLlqNA72GerkrKQ6Cp7Vh/ODC2U1wM8RXnx8MTTkGwIS
IFxA2meAlu0uh/oS5WMdDXbBluS/DE2NfvqlKEeb+mkn/sH76WSNpoq/Y00Q
Tfn93t0F/ROPF5d3VNnaFngsklv3WBPu8oZx26YNfjAGg6LoI1zEhlVB4yNV
HkMwtMSVx/e3uOvm7REisIkbXzDk32CG5PrDOf5qFT/dtFISZ6EtNzqyyzRA
PxcQcyNnmHrrQJyfsV/INFOgbU//r4Y0HPnCqHjCE4roF0jo7EZ59/jfJOMK
8NvZMkgGKnvVM9wannx+0u36/JqPGa2WyBZxNz8hu2+ivHQ0ivAtW0WW4+wr
8MnubY8sYc1Hd4mO3prb7rdwgfhyZSjXkv9dOKyvr9Fyemu8Y5WSh07w9Maw
ZNb8nzEcMu5h01Rfmu4Las6sxAtDz1xZ74QuzO/Gvav+kPwhCrLGL6wXIWfE
OA2n7ybumN9ToOWwDPEee4eWpzIQj1UvLFLhkt7FW5MdbXvhQYd7q9ccOkez
WzL/J6iCs92HtHMJ8D2vMHvaovfZr2798FWYMxkHIak4Onp1upmIQN9oa/6k
a7LqvobwNEEae2qtRCEK8pw1FEthVk+2KsvES6H0pa14J1hBlxtUHF1gV3kz
jpJ4lS+zq0eEf7t16IDe6/zweGFOCa/4yzyPHjga53BhodyNvGQUPWi5tqGI
LJGmIV8qnB+Wy54kq6GT2Pi1xIsHC8oxjFwVmSjb3w/uu5baRg4e2yjTWUKd
0Woohx/n41rAUJohEMU3V46lp1kcfKBwAWIl75qrPdP7iteErW0AKtRQNIjk
F8e1RZQiTCo4DRVacsFdWdhEXuH9/VS2CbURI2yqpinB8NfCx14Qmt0pAauc
JV/XZXPun4kNN0Njiz2jRnOaagtfx9wNk36t3hUBkH5qRKIL7Wctx8Fb7JPn
vNbeaYPFpSCANazO0GswoOOtZOvesaCbmraBKMqTttdGf8jiCx2EJy8hkOy+
hWXASKzIurJDjoTRaYP6T1QqQp9Pv5HTD2dlACfNozEGqRX9MJbyorRXuN3Y
gaQGFyOwWhm634r/sDXrZbXqRUPd7/NWx3vX4Eco3iYdq0TxmvlziuFUYw1S
lKa0piD94XGs/KuNGVXbQXqSIZlseFCbsDSp7L5xB8kubmuM+wNPh2uRzr/E
yTBDMPsqCumyHA0UVg21HuPxfqD/TTh2xXx1d1KafwSZObjFhNVeUdsW9pET
JmY2u7LCYTTzZAKpq0bFipOr5T0XUYFjTwHPwJfiZx0X+LwcVx3ufAFJhjdp
cHW6459Zc2D9K3GpZRAjH4OQHwFuHJoEOfjHBGmlvScoMSj45NvWNU1zJQrW
EzMGj5E/eGTlLIaQroV2Zj0Bgl0uT2LaxROvg2Tdlquy2r4+PzbIu5AdS69d
T6RvKWDQ9hCJD1qlQXZ8kZCh84qLakJ3+wwHUYdUDPlZcHdJnJE7565bVJqZ
AupUbKTIQDVsb1YaMcWg0giSDDXtgYvUgJDkJYjDhvCp3Bo3FzbttMSaVqap
XYltTqTRGmWcjZ9+cbZMHEVxvCiyjeU0AtdKhStdYHYJQbrK3C865t/2nmHL
2KN3EsLNpffpVHJQN627E6jbQELoIP6sYmTimTOQFXWGEdOtov7SmTm0fCg/
vIwm0vP48+Db0NkV0oEHoMLKNWys05RkS3FvUNf84OxEKOkFmVBDPcQuPzu7
jZ5eF3J8YuwbVs0DiN+GoB+dCEjjuNozKoJHO2nj0rYpVy3EvOqS5VB80W1l
2TUuG0ys6ml1Hpt3UketsMfgnYhaIu3hoOChBuRRA80MxlV6/V88h7fiZd4g
lWiW1zZhIJbNkh5ZwRpGZ1GtNwoiMxhQwOA3GD58KTU3pR7L9f/9+8oz4SdK
AlVUAnbDtFpZqkOXb1EqvfUs8vV8PwLqfb+kS2KPczLyECWYHazK8eVI7Xwa
Kdxx9MkkBWMQKJJfBm/aNgaCw8/qOtiOtqaJJdco4h4+KUnWunC9ijI5zL+4
GbMKuxyBrxoqGX1rlrluZQbMxDFZwwNmS4x+UsM0r2Pcw6xKJJgRAxk07efy
1hjQEyX2SHkPalZLy2dse4U+YVGO1gYAVWZfKS8wQNNTsDoY1Dp0M3Rzi+kf
SxWoXmUzh7ORhDSPQGXC0YtQNj3YGrjMrDVNWpgvAWA3uQMVBa0dUFoAobRy
4+CN92y22bzdgZLR7QqEeKkBmNsqiVSfq5OFRFewSTuCKwzpbiK3rvNRJsOa
vAepR6JMPouY8ACEnOlsZHShCcpd86yn2udcOxbTlBfkQPUV/aBbhMiWRUqe
bsSSCXILW9vIXfX7eMPtXlmJ/ZG5ZF6TvwB6zCAleWvdNJ1N+dip4vCcroCJ
NBduTNtopMdilmNrGOs856CoInwpBPoZaqLkgUcnWJkzsGrSnGsZ6piY5ALo
TSMS08dASBKTYYTmJFMq8RZETPqcmagOxbWlDwpxZvsANqCq3i/LfcDgdEnK
o5EyNirJ28taXKbFqtHWrQeiubqCpjNSAS6khwWHh54fgWLBadEL+yeQxjpQ
SnMuAsepy55XhUpsMjrsmdl6nohg2WDCB7rrwvE51lYgrVoYhSpkkhaNaMhg
mXKv1s88w9huPaEDmnoE6gPTL9s019cypHM/NBmrYFR07XpjCwKWckxfPNXI
Ib1f6PWXCT3MSlQo4HuH2pIPSCgSOCuclx3nozArXj+7Yhodfyo24N41fjUg
JmH5vf9ta11J5ixOJ5lDxQpNJCKNXQe8BMIosI7iiP4Sw5HPPmneblIWZ7wV
it1prQSSdDrkFGwtpRhycD8AgVVw9eqMN4D4zlrw8D7k+mAdCVhECbhbvB2v
8SGJrlRlkrmUqsRvDSGI1pTh5Y7HvUU0vuY+ubqUg6mJxvvcEXT3zvl26uXE
m++Bhr4IMCWU1uTURPYd3IhIyRTLbxyHcFEp6Mr9pxCdqvCTwvG3E9yuS7zt
GKcQWCFp3uqiYje1kXDehi0fru8kueonBoVVZ16GXtkUKFD2TJBDRUPt0kY9
Nm9BCGbGUYMNGmaDGNz55QvSnbvfMbFlGuvU8lpc7R6RKKQmwz1VPVSzMONl
Dk8I68ADPei5CLsV9SbdsY6vuFn1G7YloRX68Y7pIgSK2BD646IhL7C4/wFt
wHdhYbz7KASiPFmZ+MDqaMWj2zhhsqXKwWBPZFGbubcal6eGGn6ZHFAm9qSt
Q1yNV6glnambtC9toqGE8ObTRPkvCaBIHMWJcRtXLMXPgDb+DTIxsbyuAYWR
+u+wxvZcCetdPIm0gJb+h+i0Rh+FDD0wyYoSg009i95EhOeAkfmtcBU7GnPV
8qLKSFTeQiOigACgTlKCKrrbNspiUySnWKCfdZaczluwD7Q6BtlazKo11dvp
jcYlHQNAdWNoQIFEhEFoQzJNIMajAgnr6lUGdYp+hWOKHcl364mheKeL+EFp
mw9pNziwTJMJ0aNAp9lpHDxBqoZnX+rThERfsqs2f2nOPapZ0E1Rsu2Pua1g
SW/W0YZU/D8qa99DYa/4hnlKPAKxQiz8ZOuJNniE0XMFdTSLV7BQbhadE3Iu
rxknVA3EjeByURNIEoNNkuHIDaAJkBo/SYvT1/XBz/SHI0ZfAXNEvOumLoLA
kJe1d+ZP9OPGgqlA4kU/8XLb5bfaKPlXclBo0ehLqsLF84sKSjp+6170yBhi
YS0OIUbMduV1s1vgHhXBYB98ZxCFaOmrfZu/gxKxlRSywNEwTMGcAAeZIW5f
lLMXPrXLuI6aXmqBC7tVhAvM8YqK2ias4Xe6o2ZvJUoJjCsLgHmKm+JkMDTT
Hjx4bJiYQpfArVHuSrjE1q+7fH4qIZBkYyJ1zsjjnTr31B4KhN1G1lE2zI7q
gBZ/VRcmKQTuyeEGILHJfz6TuEQjtL142L7TypZdNCqpKVz30sapfOYfnNR9
BoMGvkQ7z2niJuvBQklhat31p61AfiLbxk2y1KynDiy4hKreRphpMl8staT+
xxwNW8hMkGIHfAjMUD2LgrsdjADNavkX6E5AzqzgPorxpueAJcl5/+TaYWHY
DyL+n52D4HdcV1LAC5586YDLC+ZMH7+LiYwmO5f++Qf5zi9M//n911VXQraJ
eiqU35wXnUyH9HjL5CzRpnyKatU9kR8KJoo0W0iPodYJDQOF6f3RRvGsXd0+
qGLQwU7A7G4Orw8ErIGwsFhOXGDpj0JyM3VEfKZngNgNV0+qdvzPqDL1az60
8WUlRGYkXVwUmHqyUQKHhNK9uZOae3KOro1p67ux2kgX+mznYTu1Crs5kFiI
LEpGE14q1BKJZREH8+40QSyKoCE7niXk96Ewbnn/15v6+SGIQkYisGHJLKkN
hv5OLAYDHR7SQkvDeNLBAfs9KQaabeQMZyaJeQ9Umm6qxN+2obd45WTDNT7e
GD/PvpWoIEEdXxFWSj5pmTuAQXscJNbAcak2wfJ2ZJKyuOCARjtab0z+MHL0
JARQqdB/nUVKmbBfKQoIJAcsNvytJNVnA9G9oq1VdOb7s0rL+y2zBW6GtYlE
rRFQXbw+OPDbxUyJEl9rTnDTperYipYa3V4f1z2A84En0iGhLIeT2yt2Xer1
Zz9JjvCrdmX3BRrSbKm2jrY9BTReu4LeMdgRZArIl9VWosgl82DQoUfFomY6
iXDcbezE7Qpq++JCPHVZ7kzgvHK1k5fjwU/dov/x2iBc8wCkBZ9dTtjosbh1
DlcgNQQcWrg3M/dRqj1cB20cGA4/0xW/c6DuAyfc2HjKY1vpeqy3L5Sp8GQB
iZ/KNSuuTA8LLdCUKTr8S3tgYtquZ68Z7R82VjBnY27vaXELqkCRTk7pT6T2
C+KJEc0l1LiMyN8G6EKfh99XnUuZ3ShyzMyWJdWEsWPk43K7OsnEQwLfT6JK
ns/3ABFWcuDQBbtPNs9DaFS5gUrGgiuLawnCdMlWt402he9hHc6zqImux+H8
MNukRFPKZJEEh91/rEaFW8yJDV0LY2ptRpIdxH0DiV12OszdWnq0Pa3RTGnS
IJ9hR6ZUejDr8xVT3Td/uLOur5rvK1Rj01+nQKUQ/YHXMXxyFI3bDRC/WRIU
EZcamCIQReVDhAkj6evnFXSL9OXLXo96vN7rgbjUvtg1+hveZSWXoFLVYst1
xgFiM/mzMXvbUvO1yo2/3HgCk16hiGkYo9saF0U+twXVolp6Q2OqhEB+b8VX
+FTdrpbLQwsXyg29kh9n2zJ48RytZ0wYD1hfs/fkYRMPLIGJNH7eTXKWSXj6
SdaCzPWUywrJvIM0J2z78uUDQ1v/ajxoElHJWSN5TOSW8RDW/58c3KXcxYj0
R0rg0okTU+V/omubJ6qRVaX6zqNjbXGic4VUk27476zqL+WUecNUjTbMKopq
/k6qi397fcTDscOlM1kvr2zLBUPMO61/cVKY8zbnPKFoujFGZPxZeYP9aVow
N/6KsAkPEZGT0azDy9VCx0q9oBFsLwyHuwBfSrYQkoTxNza0q3NZVJNnl/ME
+eg++/zZhdXemsy9rgh+uuT5C0n6Mhp/WK+4V9xePc9x+z4pQhe7DmYIHAuC
tOuv3uoK+joZl5dtsxcDA8aCihTnTyvovuBGtA57tOo8ebBD4OzcsCsVib2U
kj7opJOrLaUlW+8oLIcdclfbxKSaeA6qElAcHxgwoxpEFdy79XdpDimA74KX
xDUtDOXODOKFeEwvcH1Gra+0b64UWzKoqqEBruOLYt4M/rwK2MED/OEhfckB
Fkg3TnKi8jSxoWFHZpk5mSXjfCTsnSdEd5jL5To8QfpDnUXAdEL3cpDvrEz2
sHQ4UnnR/Y6Mq8kBH65O5SIBYCxHy3nVEC0neuVFOgnuzUzxYx9JQSwDdc23
rPeEUZ5aO6670fifNI0IjDNag9JSkPDta2Y1u2fiW+25yuHfWc47cV+ZTQ81
UotR5sji5tOUhfIbv+9wtWtg0xQNKeA4E3s+9IOF0nkRFvrW+oRwUxik2PqN
TNEmPOssVaPt8OouoXxlC7fOn7zx+GorLnx5FeLAE2QjbUBumnAL4Pd5vCAj
kTC3N1qn2KtUfd2bx6p1/6JKoi2fyDM2KaND2vJqPJmQ4qxkSf7S27/2T3kM
6F2ANxZIr6mfbShweG2MfX7RS9lq/Pfm3pw6QaxQcUNLM6WOfDnIPFSmYPDo
0x8X1M7x8XgTBrfweqlPqCc6fUYHj14QzWH0wHdnMH51r981t/Rge2oqzaRI
6LzS5kIQu55DwkVVz+RGk6qUD2JXURNT4xfOGN2LWW1AT79kzLj6D/ewK+sU
NNjz61UsMZWBreCE9P2T57vVMMFG/sK0lR6fc6P8hRCep63HZYgmiteaOVRo
egYPk1Se2sEdLlmFgNx7w/mf2Kz5CLMTGUinknG+LvMhUyZ8QEAgsSQimzew
WNbC9tk+nwhdxVyg/NiDdsWs/M0qP/PKNDaUKZo04iFCmRzAB3L7umsGEvMY
EG9x8P0TbffTXaQ0zHe05+KMLkRYq3yUVHr1rjryRkma5iSgVCmsN/HEJXFJ
tnDaE8kbbat328R/Jo+S0NQNQTsKiICO6S5C8k/klomdpr8t1JN+kY4bOeeN
F0xwC4CF/rtbP7yjd7CdAsZMBAvh+pKRtf5HFCot8SiJtNf0PSjGyi0YEsv3
1DT9ZNE+pE1WJ7CJ1g6bLckSp3O4OxqdiK4r6o8kDXVZwVg7KqhS88kKxGwT
eHHIxw47dWAvEcRyvrGD2t+0XpZuzj9kNCiXk75munNyp2upYc7J+W4ItmO7
YOPFwq+v0pi0BlxbM9bS/OqSg/nCxfg0fCq/tn313F1remESdoJJGfvZe/YU
tUYAJgPgZ2QYF0Hiha+ENGAE3I/bFhX/I/gr7dBFNDK+5SPvm8AeCeRjiJSb
yLU7YqhbafnSKsRORGlpii58z5O4JCmd+1LXTtKI6Eb5GxTSScqTD0WlzDNq
/V6qkRBh2b3riTPMfv0TdYIkW26ECoNVbnsfC3RpvxSXhtXM8utgT7IoTIqh
bhSp5RekQ8HIbZpNWnH4vqzaITwLg20Lb3GIb/YPgZ8FJzVX/+brG/F8MB5/
b2PZGzk3PTMtGH30MMpBsWXS0k3nVQTlMrL7FDaV+EuRQweN0P/k/xxp6+yp
HnHUwfoq2KEd43maOuYt8KNIsijA6SHAgDNZm4v2RuBUY38eJtygHT7S2ZWo
4mN7QKpHjrH3ix4LFPPob0o2k7tQfi2s+U/Qu93hHVTk8le1FRTd8d344IO9
vDzFlko3ju8e9Sw9qshRqgRpQcifuT6RSFaCCxspFFDmrv4eLDJJbF2ZFRuS
aR2xTMP+tYwV/btfQ+7rCaIf544udb3mObwxUfj7pBJIgqKebgP3eInaxQNe
RrQSgyLQKTowqKsxRxoXjQFkD8qkhvdeiJ24IHmJc92L4aNCqvx5mSTw4jp3
x5CmHudLVo2e8sgKDsnmA9RBUVxiIzGsCxGH5LUBdusgjnKC9AByyGqyPizS
nrCXFsVFvguoWmUme3qKc/yYg4tUpt5vOYIPIHoqh5n05LWnc4s2krIoXFJw
Gj55UYAgVFbbqGIDX2fN08CamdjVO16ShFVhcE7FlSJrFjA4TG4YaFvNX/T2
0ETqVY3WnRFWscXEcDG5xCkVbUOm3JEJNHmXatbpey7SMBPtzfds0YOq7KxL
/05Kx2sJjYrqxZv6dioPkDrE65IKlBZ+z6lmE+XWk5FUpXqHborHAv9iCTH5
MQd1EMDamHH49/H3zmbtyNkd70t7x5g1T6bHAHbrGcdzzIL+twxy6ImWSJJ7
NM3m+QwuCr+EZpSVI+HTZYN9goHGpW0mUUMjBMOX8C2cGdgA/Zn9UFOieLty
uTz9TaVSEztu3w/z78Vu9AToyTjPSSWD7KnQXo0Cg5Gc2oU7PmWJOVaCHNgj
Tmubm93iuPEAO9zN++ogEw52+xxB8kDUJjpoePnNDc3EXac0WG83D5yegYXa
efEia+PqtKu4AUxp4ew665jMATMRQTLR+9DPBwlI0arXVQZozl8YIzFdpYbi
Ic66LfIr52vUaJ/TeKJDGjvvXcKuT/kYY2Ql30NPWp6qPpueSncvrpS3czhA
B56hSh3ja0c986k7exJfXUzu5QVCuuMe3YkU2ZlIjtv8c87BKOX+TKfb+eEv
YdA0K6qLz2MNobNBQEVwktSpE3aI2Tdm3KGA1WPJ0OZu5MGaiV1PsKmA7SPz
HHO4zjVHOVGVXND0p0j07olNMs6O0LrMTWg6pWyc02zAAmArL6blnG4tj+yJ
2X942nayDR5u3BcbzPaN2yxdV5njD3uD/+tLBsRO34IoqV7ggT+FP91pXjKB
VlloHX1eoI2z2+Z7gSVKLbwmOtSYQkE1tirXJnly1i3bQuy8qqkKfwFQrEeD
NXXeWUlNdX3pa+3OK0LGafPhPJOzkXkXAJ6dk4oKk2UEngJK7Pmb2W1YLVfg
5Sfbg/oq2hMaBnhyZPFWTOB4zd2JDHOn3LZBZdjxwPvZRZu2puKkgJLBnzIC
ytK3Kt6r6P/kKMA5Ds5sDkrqdht59Uo+ltWuswdHAGZ275PcdXk90or20NR+
CrmpKkfBIAhNUpEpwkaxuDTlBlUW7eqFIjxEdVIieuoff79IHSpcDh63qbn+
bhT73BPxlEieCxGOTwPKILeZBDZed8hhR+lQc3m+FRFjMiW1IKhWuBKz/D1h
TiWpC9ZdiDkcpshDpsBd/XCE/uOuK7DNv9Z1+7TDgOjUYMFuahq+MRD0RbnT
+Kh0ssUT6XUXPujwepK7CvsWyyZUowl0yA52f2e/KSR41JqFObuufw9IKQJp
9Y8uIhJyFuIM4fLJ2iftCxzEnVPqK7q4Vlc1qHNxqXW2HdFKIdI2MREDz834
GnY9rdEqFrragHt0SR/ztzuw0HplBoTlyj840g8UErixxZARsbACC422A8Ot
MdSC1vTmaLVGoPRHQStFpOfz69k9gptYfScS3kRdsjBUFm6j66HuKibjBSTp
eMm6xo3RtufJKRaewo2VQixVDC2I2MYtNJA1s237IQlyu5hbq8tironlDNsJ
fLdOL9sLqFbrF+tg6WkyNC9ZFHa12rq1X1XlFHEZ60NeG9APAkg4Xgh8TRu9
j0jzmnAgZlSs1fxKLrf1dEhKxtMehktVbW8GW/z+VeE9HknZ+lj4nqjzfdiL
chOQxrw+Rq0uwAMQub2sKnUvBRNTO++CkaLVHX4Ci+wi67CGF8CmPCEkQCB0
PJodkIkrfI2J4QygXupS8lmgOWUXsDY8smHlY4T8Uy3p2OsJ+Gc04moxEPKu
UfF+BeaCCYvoHZJjot0SZsmga/m5ZzfNbNeMzeg/RtjxSN2Xe1knfCwakbDH
RYoK4E0q/qDzuucHn1yq5AfB2fnOmf+6D7FOI1GFREmK/p+Tkxz+h+jWfI07
kxR9q/2Rn4PUedc9cLNinXitcROzKfijWGSZ36qQ5WfmcuHpjNPYpwHBS9x8
4xh1UYrOQdEvp8wDU5bkJY15XXgPEyQZIEpvllJCLirF7vlLgaev+yzvG0iz
nC2TIdGua6DjRN5a6+RSAyVcLkxIYRcX9BGFnDdVR6oFC0o18YDG7WAUF7u+
QSilwPOXdjnXNNEbhTiTuvKbV4XZ8t2JEywgcEjMZZxzutWtVZAAIw5gEXzu
7ZpRWPWCHyzgY7w9RqJrUqHHK3aKnKfm4yKwZ0ZEWqnbJ6C3HO4u9MZTgT3F
Fels1wsI3h4A2OgyCwvu6nGjExI+RQCAeWevGWg+SXmDrIpKUpwZkay0o+AE
PlrLEhFiFWXDM0UOw80YdPlFAvWkmvoDEsz15NaPyfTb8rxKtFBM8efOL6mj
oaVYB1JsHGPYuI5RgQ1DP0Yh326YADHXHO/p+FWuu/tUjVL5WLT8IHlI/yWZ
6UKiocaOGLGUPcOVdawJ5xx3ErDrzwuO/8i+CA/fMfeWzcvUCXjD1f2g72/d
ba4n9KjTH2Yqz/uqme3PLOOje37p8oSzrqfT49bGTGgvKJRBwAOs61OuJ9Bw
5u/Y9FkcNus1BJ05St+zcxlIiJ9C32MvHmNs5H4HsiSFCMffDqldBpJcAfro
uPEkgeiartUTjKgdKsW2hvZTfUYUTlcf5hal2fn173oH1/QrXPPv7tuKJj1s
1FW2t3f9pGEJks0GkhyDA8bdFnzTdAMmo8sxq5kutqnYxbkTsKsLayDW9/cS
Iao4yPfHxGq+0Nb8neGE1fAS92hUPCvu7FseDm9cm94kDkGi/rPf7QyFJdin
9VY6/d6E0mPIGcgUmkjoOPlJ9Bye3/ReQmsZMLk4tepiFW1h+IMgxYk+oZGj
SC+ylRG8+4SdV5vqnjQiIiYH/Iqj5jnTTwO8/hvyGa4T40AUbM5WDbnmHEGd
MDBHG9X1TMJEKpnO9waygRnZo0KRct6ImEqVBW5LyNR5A9sgbgj/nRELVPrV
OAlJbl3YOMbtEf1S/6erxDS7t2aCjmKkLQ19fQ8+DM3PeI9RWfG04pCwde1q
TZvCOVfWeuOjqJtHIImSi5fsDDSIPX7AedDCuGgt8qVIis8TKys5AM+djrU/
a7OVt5uxHuCh/JKpIEfbIFkxAhfrGFigop673kHjr2eKRR8SuWaSBVpGop9K
85HXsKPgbr/SojictWNFoAFJIJ+952QtB6tM0P0SD6uwXlh30rfxpIqiag1l
XUndK1VK5b99GP5CXcyyQZIAwflQ05CBRC6BuihVTvsQIhdgFj90VIW2iqY9
2bQhgs8rdFLMLMV+U08bbezE6EHO6dc9mAmlIGrK2LpdR00UXhL9zEkbvN53
lsd5DUHF4nvPbcqSKkP6by4Y9tAIQTexkBCr+1ZySUKDE9yXJprP75JKBo8j
p2nxk1RgsrOZllgQ1juFehuOxGRVsN+70hXtRpB/Jfz3vD3qTdzUouFK13ET
2qLoOkiOV/h/uyLlhRSsJd01rE8MbtWnD9ZuS6VaMxu0SpNIf/a+/b0bhJfV
pbosgu1Cu1gAW0QTo3e5uo+Za6T9wLExw36t7i3E8bgF3Rc1wMi90F73j/l/
ZhSa+Ywcohjw0ditU+Gh2V61A9GhvCWEpNHeU+8m9Lvf71elQCoS86MRttAO
JpDR92Zq12FZh1julrVT3+Lp7WwXnpOAPV/4UxJg+pwqaPkwdyydGcrVnq6W
2aVjuSVkmshVxKz77lyczFpLVrMKxXxc8fMMP6x/R6OpfsKp6a472WkwPwpJ
NGFMWHx8zI9WrkLPoc19sTQkUisTAe2/UP/LZkH5OVR9REzGhn6rbWxjSaAX
Z4M3E50qpggIRadBzwS0tDzUp+u7+pN6thYnj8nBXaTo5HsrW2ewqGI6rQH+
QKZ6PVbb6q6TYvXUf2csmA7ITg9WVKeoYJ/EuJEQqPzm66+PsYwmheku1k0h
zB95SYm6Qmd21GPEk8SbkeGE/cNxBZfKtnJgabBhmEQ6nGKpWLu6D/CRKDOB
glGB1KpB+IfB3/ql8V82xW8ZQ5MKuGGlbRhVUIEGR0CSJpsbp9CuIYDuzLJN
yl7/ZOH6eqQ5Rhw8t1ByKniTtCsN30ivpazIO0b4g1xwfqOQB9kZ72wlYJao
W1llsMy40DsoDCqmb1K6TgNipcy/0MJbAtZ1ptmTWl1+/HBCetQCYAp4qHR1
V4IpmQ8Zd9XfbS0wSl6plDoZtkppSc7QCsPOIXKtyJgAZHbNxbbWltOdjxME
uwBOKkjyywSNCJvfKoSwpVatoCppKq4gGjDlwSXbtfl+Wnhbxg4PLGLAJOEL
gbz64wMG+LlF31jZjGegRgWP5Df4B5IExf2+KjXucayeQCqmZECC9m36JjZz
iEzPwBW7qjCL20UgtM8pooH4qw4oY9hGYu/XdkPxepgzgQ5CE+yA6fgfTstJ
G/i0nRvmEmvcQSgpyoZdRL2Q8uLs2Rz84QLEMEsVJb7agp2tu+Q+VSeQRC4t
9COYcdYxZ3qhMR2poKu6AGb+dgfNgfBlOqXEI3S3EBOiCSgfBgjzJgVWEbi0
wjFtAMN2i0Wv08trQ0nl7mV6kdmrlzuilX++dOFW0iAx736H6tOIIyA7V7ob
ch1FzPiPi/8YlCNqPqdeyrr1OUSNbWtC/Phl/MUJHNKMC9G+oHlPM/6WzlqZ
Pn8u38PO5F6I0SVNM39nvDIjlzUhg7nj8mySsKJrlurWHgLlmzlveKz+CEEA
IH976Odcsjzg74wkdpd+dovjoaMBh1ESoT0JrtBPSJVMUMp+moXKmaAe9M7Y
OF8yR3PjkL/c3kNJMO2V2Q9lMMtkihyznwH5Heh17pGCiCZeM1nsXWMlJjRD
nob3aR6yR+IFcd+BgNaU1KVZeWD9bdT7Oz0+BIZAhw+UrY05fiVCNlEh/AOt
zxJ0K5ARCf1rskaV/JwKi0t57U/y7Sm9qNTwP7AAtrf6RJxUz3OMT3K/g9r7
4EFRNH/baKdsb7DJqoDjfWt7K2BBzgWQQ1dp7AUfErmeAaxMaEo4sCKtxECF
q8pfio1GlgzKCTxnv3S/fdHolMoDJZLkN5qZHO2oL34KfjGlVdZBjqIwudh5
Gk7EpfOY1SfHqA38tOmFEHP5JbCRSy8ptTXWxrPNPoKGrYxYRbLhsQKhu4Ra
2/fWjTUXhd0VsniwFmW2JHrGbrk4o9VRDfO4E8nWMw6mhBvsQqxn7rKyScas
gjeWZ2klY9gfavSJxHSfaRYPynTY5QBCWcZsom7d8jkuR7D1ltVt0MmHxFXx
71v9pHnl+vFC5naMKWjVsX40DNtBJ7w9OphLKYbLP7CUx9pktqrr5kiJGqGU
ABxCPwvaEe1Je+UF40xYeIgnkRtDRKpqnS+77iY8voDLP7/v1XT5YjVkLDpg
YnfEHj09VkRDemwoFGeH7bztHjjMbUGjTqlHuIKRlZGOXELuQk6UOIQjIl3A
LixaBAIU7h1C7Yyr7I8F/pcRocOIGARY3v2bOMjK0EbfnTFQI59YLhwjtfvr
AALq+kvIt31ymfiwIFTsn44Lw+cWO4v3wzTDrRCgtWcZ51ti//aNTHLe9iBZ
9R6Z0l3dk9ATYOhmOX8NG6K9SlL4cvBVD1mGNqNIcFVAHcfYTjVRLvaDT0MO
p8ZKnM5NWXJr4xOATU1Hti/mCa2qFs04F3ugxl7GzbG9iqVzff7FU82+SWsj
UtTP1ccB6po7A30Ax9PEmuznMWt33SiztbjgPIkotNztwn1iQgWH8Pou9Mwc
s0m/VkbLe2VI79qyCPmB9UOBEpYgQfxrYDdNKBcckmG9lri8b9Ri7w6zchDO
h25lFJnUAMZJ8zl98FBxbsmyDCtGDZYFzkaefd+stgIlDY0f6sfRR5lnju8x
/4VI7KYXq3HjWt75yzm0Y7wPm5YloXXPYBrb/EwvEr/gby71ALEbV8Uht7/X
7AfmzetllXB2+fz9+hFiXmGDnOQOOeO18ClGXJmJ+GjT7PpAzYAVefHak6do
22forZPzvaJRMyH8uiwkJ9u3dpPuZ6SRW/T+12HAs/KjCts0AvQqW9sSWX1v
9cSG+C0XCAyTlbn+POGdP+m5Qt2HU0HmjmiepE5XZHfaaG4qxQKt9GYMJxin
9Xovzvesyn3OXxHPVs/cp5UhENAX796/es1wX+dBsC+7W/zKBtmZVG9NfHum
7EoM/j+Hm9GV2eafuoSzAY4M9aJPrsLT5OnJaRvN/Dk9icVe3kbPmYa5lRo2
BzZmO4Rvh7BNAYuRK+r+zKwHlnkULPa4A25u1JyG/Z2vWg960w9CfCoOZRto
5ggxEGPhx01BIMOYcOrW+scV+fTjIgb8wds+Wfmxmm3tqWHtD62JccTCoRPz
XkaWs1hnSQc7cT7IBvujq85CbvhPWvDNwA+hQ+7CLe5t+dTImGM7JxPJfdTJ
aDUXZQp+jg0oMiXHkFYnja66lhrbMnNG08YAd9Bu/JvB7eiLOtO9ui19T6me
m9wDz2jbA1PRzxuoUPPGWLH2rds5Va64qQBSNJTS9OdEhrgxzl4o1p7veV/Z
/Oe9suQwfVo44qvaK0fE9P5IjgFAfXcpD1Wd8SiIrdPbYwWU7xQFbOQ8Ptcz
UlTO2R9Az0uGYZwtlu0F7Y6P6MILlXpqWr47X2Z4CM5bgUPYO2X0vND2GdLc
21csnDgxwdXaAkgdBiLA5gEPd2cWVp9kjxrBbulmstVw4OL50H2Rq9KKAoi/
y0L9D3ZgDeTAWnngbA5JGZcpzDz4Y3UbqgyH5mUtylz+79s5do2FCsDQP4mf
8tm219pS2qoIet+fixxquMCtMd4kIf90KeasdGc3Q5bmxaAQWLtL6tYmpbEY
/QJFQjHRNvNRXFmOzuiD6D5Z4BFKQD/jjARX7Qs4MC76jHThfS1O7sRj/H+7
UxdoRqkUEhFqpDnHhMJamqu2IS52+OS8Ymk2R3ImmKvOSY537xohKegKAC09
DEWNISDZIg+Wo/Fw7b8fY2TLChNnfGBDmvfn5/WyYPag9ZojJwF5IhZpVhgO
9As8QN6tONj/KC8wxMiHSWPy33Rt7RmfU0Tf0Fo4nAvaDw1Fu9200Ws28ni2
Xuz5DlIJ8FTOKO+PYXxJUY4uFpMeaGyj8eQIabI86o9xl/iw4U1GhgdYNERy
m5BqqJySgJ+vLqXQzIoYi/HzUHpeOvPx+ZqVUdMPU3qutnFbfq90bnJPpn1/
aA/naYkB92KFadvJ96Tc1vR35Pg9L32o2zaZ5m3KKAjXc9VvLe5V1UUUBwEE
Jl8nG7yddDLacXZe0qZVGwgE/YNfuZ+1aWtp0EieevAUZf8UQkETa+KjU+03
spo6+k8D+iXXl69vjtpVRMmRomdyzU4ADBzHfxvSUwWyQSaxHKdUZFoySZD4
EOGlMLsAXrMrT7ulUlFBiEoCE7QOlz+MpZasEZDhDBZgo01ssv7YMCbBAL61
vC20b/WMzFVzVBTt6NRMNGBrRDEGvFRIayuOi+MvqkvF1axFcq0R02gREyZs
ZzviR4OFVd+OWXKL5kBP0YtmMVzPiGe762Ewj1eb9yzeM1L4ebkDCUPQXu5S
xFhahMSemRZyyGhAlAmmtequAO6mSnyhq3DgS8NT8oknkLKzgEtMrRBpSFTh
0PkDX+LQG3RjCTwPVCVstAo5nxdMAzx2V1nil+3hBnSNepSwK5a5bRKelDeY
dQL72WJV5tXCiq4nHLqHkx0AqMkpEStiXyZccs7g8wixd9n+6a8i/OfSDdPz
wQPHIL80NQn5dzZKVb9z0qBwD1sYcJHXgSu9Lb7YNCGepOIdjmOAu05Do0t0
fPY1Gn+YGrexwl29ITUNqTDY0k6RKgMten8EzYpCY4nxsa0Mdeyt4iO0oyJE
3F6d/7yB1lIHytrjr/RlJuSQzy7e/bm7H80NPTceucIoz+mhsNhvVv2P5eJO
aD36ikBUu1rnQIf2YlGtcIWTf7LyOKXY3nd9NSzF+9zr+U8fZDcxEMdeANrR
CxQQeaALgBHHYRtysJrCL9NoUbcTqvtBzeZWO8/BbkJ/sphh4E3JLSbQwsUO
Gu/I4WLwMExm7QwlPEz3ZoO2L4hz8OkI5xuxtArx7v/gh/ol/F01nmN1+/uz
W+3TZrgUDIaIUnK4MQfmP3g71eqzq9hGj8CxYaiyvKJEqlqDgg1l+NQMzMMx
VNaDTm5md6C3g9rROYX5lc4calwUfVmgX3RH4Nlc8968DecYTDqhU1QE/Jf2
zkIl0EFklV9kobR5h5/8CKY0CyJEgUF7dgx7xI3u9rEMWd6hix11p2Jrzvl7
DNNEAvaZA9C/9KJ5Hwr4AiqDvL6Fp0FlE81RBFTabP8mVvlbdBBiZm3Ok6R1
hA9v71+L3W+i9XC0vtyWtGwBb5VDlyAw3m1c4MPuOmtwZIrmTbIfpTEoHzQu
OnuMw1rcdpGjeDY91U71HRDrDMVPiyCuZwV8v3UQLFz3Cw5t+H/05W0uqRhe
dEfhg5rQwZt5XcyrbA3pce89+0im/DxRwYIDwRUEzEmC9gMnd8x/RaGR7hDp
qJDb3Km9dgVVh9Ks0zkPOMumKSfjiq8AvRJb/XLYj027byA5XAI1eAO1MZr8
dzNwREGjb3qZu/nlBGMwczNSjRKEI1wReiMjAEX0lhMUzv1KdRgUahQXs2OI
B9uX20pnq9ztyKkvLSMt2cA24mCgsyzy+KYeQ353uJN9Xo35AJfq92ao1oY4
HoQZFyhves1gQknHsUspBB5aUO02/wYJsVjf8pe46tNw9GfR2AgaqcsKyWL5
Z1/dHpchlZEzBGl0KJfFEUeEA4jMjMDhUF65B+LgX8VdP9tMZ7Y8+N1yyr/G
d3X/QNVltyjHJOup2YNDVCIWpnJUp02yvYJ1az9b4bqeVTgoB+tZzLulastS
PdLoQQiNAtxK5a3HSFEHIzbCrj7NcU6UYQbYhFuPPflMuP+i5JOP5wbg47rp
wgfXtXjhjIN8zZKY/cDnL7LQv7QlDdOdagEylY2xI2t34rWYTPNPGztoZ2D8
EgYPUXoo196OcO5LgEuAVhXE5ELaKnDInYsn9kvXOmKK9eqc4yzCoIuzBLrY
NdXetAkVR0ZuEQ01KiHIjmdkyYsESqFUoYE7dKpZUGDs+P5/tx0tzwUSSy+j
JeHjVWoJBWxlG1fFhk7PMqOditlvA3RsLrYiJIk3Wmg7NeS/OtnZ6ZghDyfj
iX9/h+jDepeyP5sseVm2V/pbBGvsWk/qK03h+ki0KSRV0WcDN5J7aotu2LfO
ampJH0VWl9w0qCyCCJ6j39DlZyXI2h/1UTTkBQX1QHGyi0zs7r+NrDIdoCLF
oq8WlzsE8P0wg+ExzdTn6EUg4d+116ATStK5cSJFHjwr9eaTr/DONbRu2NGN
v1FDWf7d8pNWyTt1U74phL1WlFqjfWxGI0/VDCdSSVMZaiFfXXW3/3+WZSVD
6KnChN5yA5OLLJl1INFbU2XqQ/EbpdH7C0ot7amoD6pA3j3pHrg/EuV3hNAE
IbP6vvyGHuqbB+wXfhuuTwkl2Aflitmr0ey4GNGtimu57kBjso4epkhPzPDI
Si6mAIGgcTmEQyB4JH/ry3ek5QnR3iRKu2sPhskzJLGvb6SEfNochYTIVNcb
qbY0qLCrEPOkNZVtPChwrM8iNY+LHOoMvn0o1mWQ/OedHp6PXbg2j5B2Bs7I
rF1Kgd8oM1BDXeUZ39xxm2aFnyVXsv6r3eVAO6A06hkrYIvqXES+q4HQgfsa
MUHgQI14ILK0xlLTyy2UDjfkQVEO04/FtTbjTal1YlGRqJVWO3cLgXy1GGzb
62Uic2Hb0wY8SYGTPNhoZcVs9DXth6GCvI4lhQsyAiOaEaksuL+YI4ZwRq1o
UVl8oPxDiiKIL0VOf9fNCMRs0dJ+KlsdmsfC7wfe+SwLcUAxKBjKVF444xJb
ygyoe+i42LRpEDQ4x5U+K80hre6TTmiTOTp0AvzG+uuYIeIldp+/pr62kEXn
slk34tCRjcVS/Mpssl+VHJAfQli+Yd5CsK/oV1zLk2tjRugDRA2tKQKgqpbO
Ra+jLjwgQvkl+ER0fxZsDSY4696KmKXF8g3Fsh9motPvX2VUOW93kJcH0SMT
eM9nhn5RUh/q+FLmOZ6ibDBi6Kd875Obz0sAbLLI/uX9HygWlux67rz2JRJ3
Qn/1oj97gstUZCKt0Vkho+ReTv7/bgLqi406LkK7QA6qhd0ZgwPrOnnA+I99
DpwvBX7aV/sWRUnq6pCxkxRrYApYmUXPXjhCvIX1tMNMOIaZgffLkxjuyWn8
BjE3rzpCWbk1j333gihIX641xfVs+MFGNKO94L25h9Raa/EaGh0t5YRvbjNr
wAuqNheBpChf7ioh+1IIXIg+qEVm0KoL6qBxYRsi7Ewqt9EQnvGlQeLtUyIg
iSrVV0uEnBGxAekz+ro467VFQugGguaCfXyydTtcMT/wgeumKkjyYuDgazig
gF42z2gYnsFqlAlpghwPEazAdc+mDxKhh58ZbU2B8VzKGxjl4+r6l9qOQGm3
n7Xf1fHkst2JZ/OjqgugqgG0wqb19vMhQwcoY2RUhdPBtMdZUPzCsvr4x8DQ
z6a5KV+Sn9qYJM9gQ/5gFa0XjFaM43FkMxv/urGjfVehEB+ES5l4EEogk1JV
RA+CB23yKJnppu9F0ujtu7AuyuvtePESN8KbbaPZecnoJP5uvmoMExcWz1HU
VPD3tx6NNWdyPcstYhzzoCh63y8SOfkNY2ldTvWLD+pnoJ4hF6m+jyzQHBgV
dmlPB2FLArhW74YTl2RSC1JM32+buYWvVbG0Tpr9fbigYI63J5OBjFmYMGaG
VOAXV9ozrmGwGCsRDcByRTDRRiBL1se0rrWN6SKkgImQE6o9Sy4xnEoHUFs3
xNa1oYaLbLmJNRXZao1UAlsmdGFba6Exvk93ZhJ0pmp6kC4CVe3dg3hWYs5Y
zWxkoxYxrGbTzwpPI3m3dfVMqJt/q4S8xUH7QgIVrbTdpYp8sv56ueS1aBOy
38k2jDeV7YW0KTaAyRFO2zotdcMyP1BGtRuQTbSL8CEfzFAIdCFjr/pIb5x9
kCTpAzkYk+4KuLP2fJw5Qz+gC65Up3Yr3FnuYqmzHRG0dKUg8MYYAeN4ajCn
gKSZVkijfixJMGypCVcfmPYuXmT1tUdROExTgKq9YMdCtsHm+PGcGnhWgDh1
qcpkm5pA5qjJGeE98jeh+uBFIT3rZkvePQQwkc4Id3wYk5QtpmKyrBYsMgtl
jaFxLTw2gMqUg8vKryfDHmwIEWX7Gws/lNywwxtPo11zfvrJepPdVlSR6BG9
JP2pqQu+m6a17fBKDmQgm6PStXIN6DDruXCzOOYiDRub7ME0ZzGzr56wkIHZ
On1ziLyrDtL+/3PhbNcKZ9qgrC4CkxqwAq3yGaTxg0oZi/Eb6M7E2o3ET6lx
0NKLX/Ld4tr0JExILaQ0/13smkYdJcDrOPpiMXZgudrsYl7Gg4uVzRQ0858c
GctPcpFvbS4LOCoKBLBPJSETKmx/gIsj62xRHCz1N7awhi2TJJEjW7zCgied
vUiEqEYYo0gy5EMiJj7+6BcUKcNFrzjxKRkyqHk9a4Eebdh4hNtSKnl9OmkE
NCf5bWhHdaomMfJ6VIpSr2xPavs9XIUECrnv//wQNjIHiVlLj6Q3+SZk+ZXv
mXRRrdc5n+yoTsDVyL8HVcI869IQ/nppZlNNy+pYHgFqvRfYp4fMsG8bTOdM
jqBOjeU1QGNzKMZHqV9OzP9yb/mbvuPlbB8j2luY0NCokGm8VmFcJAc+DJTQ
EMjbiCHJ3Krp2oDSkNudhUqoUMCigdYM1AeFMlArmrx9o1CToeZ8gDU33JBq
EfwWphwruhceYBfU20aTPVfjCqTah6HF2IESfwxymZrZbsUdmIqdNQnJiG4h
mgaZY3QBesNhMhaquQHHm+g7R8sQzXB6g0EwCe2Cqkky0fVWUSEpOrOSTqyc
CdL1mT9KICGe3z9Xjmw6TfPiR51H6zYwfDvNfs+fN/qv8BJci5RYLkYHFf+K
85eLad64TlreIGbrGPgk6wT0LqGmUO7reJe3PNkIiUODdDGGuRbvK1GwOOgX
inOwCC2EfYbtmKC+5awJP3MxxSpW8F31zWsEB5vLigC6zPez4hUvPhSuL0up
Y49af6B9sXprWLVbm/9N2F8iTnY5SyD6U0h4hWN329K0SFx3kCuX6VmZKK+j
btfrLAR8q3DbcZZQqEPiibTbuFGYgQCp9tGZQCJTlxSE/qaAsQURnhTqKYi1
cb335RfkdKcwMlf7lo06+PJBWhNmIeDTBeLBTtLv/WAE2gE+5HifZP4kPohS
/xHfw9mG9tHIfDGqzyJLPfAWfxlnYx257oLl5Of65swI3GlhUJ36UsKyhfd1
fcyz9TQ0eev+eO5aoEuBhG3PykjlQlpMWP5L8qucx4GEnttTRYdrK2yeluCz
GZD+TB6IwBTnWCQo96073gCaUZVsISzP55xkSoicUxBLTpOCmPZ2NWziJ75c
G5ko1aARs4+kylza6ZgtiqGP8iTyhoVACaJLPdPqLWw3tedxSas2lQO87HlM
JMzz0AEn/NpBNa3Jrii9fvWn6xKHHx4CYGFQ53jQdF5PolVvUDUlrLOLiuud
F//kj8Y6847eP7vHCvTmzQefw4NXS4aGLdAwuzm9mCSqcm9l2WwlN7lAb9Lh
vX2XntJje/FEDHTtOa3dUZYFqaWHII2iI7570NZ7tycGF4BUMsVOhQr4ix5i
johVVWWQa/K1qpqPJVwDaStiDkJc48RdfZx2YHCzK/yeuuvxEvf50sH5RsSq
f9qRVaXN8IUx9a/mAegDGo5RDQKizJK89o0P6WmYpE9GHyRPXz/xSty0zAUr
gLUnxmPA/+S+A71OVWoXR5E03l+GAAiPl1P4OPGAdAQqLTeEMHwBZpwAgdpP
Gh9q5as5zOp+eRYkLsm3LYVHdwrJVCl49uaDPkqbGCASDs2tDlgGZTFbxVUd
DPJNy2D65+HQNzuR4UQUZz01yfe7Fp5hHboB9S2fL5Gw1i7RpbSv2QjC2wK4
zsq5VCoN8E6mwZgerkTokTNC5epUuwV2HkWTl/14rw41FtjOS/e3hIVXjm4F
cJQPeTptziOwO99CriCs9ofyVTeSVczFZIR6lp4bipxumgrGsb6UGCGdcbFN
91774Bs7mykrP8HnZC0N0Gnf+7YHpqpwiRNRV0INMwkK7f6MEp0iLemZco+E
+nlykh0uPh+ZKUpE8MHWn4/RJsCdFEP1OSNPhIQjVCo7trogTrRj0WTosPSA
/JE+n0k2EOmT4+DfWeCmJygUSX2GxK8RqlydErhFbq4JAzjrK0M0HHxQBaQn
xsYJQVbXwmnCRd7mD6KfplFz2X79ukHvjO4AlhsyTsLFktUIaDi4MpRqcwxo
/w/ptPJySZa+40xp8FIjZZTSR3PwyJDic/yyWMxlpzcTWYQgJZXGCgQXEt7O
LKMOCerk5QfQ/gs7X2Ipwi0+gIKNZGy9/XtPIX8HN4dDu4PvMqIug9Y3evYf
8VNhjqmt7Oc7LzCP5MSPX2tOpFUUu2LF5zlKrgIu61aUE2ocfouPhnBOiLuO
Fv1rLK5Ax+jX297os8wQkxpQDLfXEYNNavBsFo/++tn1/+EI6NJXq68AhWE9
oByrX/YQLAp8r0J5wMOuoUv955Bu5Bm3rb1gBA4fKErjn+QLqzaddtiOI6Ky
C/IdMHQJUMKdIZ4cwNQFacVKPjnRblnAWBT1h4ypIo+C1ZvOXN4twKAxq4cZ
ThQwG8Jy1XHWTuupdoj6vSP6BJYrkBoNh1QrH3TxAPw23m83OKbNAQzQR0M3
4p3359dnpn1Trl3um8t18kArOOkjwJaqYTgKdMwwQ8eR5xhESivBB9oVfKkF
ExhCg2DR+/iOMEaZqy2bjUYdXSUO9OTOpvydrvEyegZScUoNTN/5XF99EVNE
/0pGGlwO0Q18wDqPEwS0zlrbOhhOaKOZyd0DSCLyM3uHkhR06GiOQR5QT4ej
oCAyZb2F7sVtcjzbzFSueozGA7gdZUn1d4j1Z8QBgFnaAJzYM4uOoZCDDzPa
EqhxLnhjsVSTsAEs9LgZhJroamxY4fgQNRmw4xk+E0oUrKKjPtlU4/En+Tf3
JZSud3deL1IoRsgjQLRVt5lYwJzfGWS8ubI11W1hD14WZu7qAA+lx7fZARYV
YqddIcAdeoFYPhrDNzb34/AJESDdLYW943yva6O8iik58V8iGkNKaHulmUb3
J05/oYmsZydlpy+K0OxbEsAKcb6BXi4xzMDVXk4mG7TPsrm0dZYYwQkxhWDe
ZQSIuxds+IEg/8fw6RyN1xGxpBpTrNjJVHO7l6Hh2iqDz+DdrgxuZaeunH5b
mLiKSEMSZZfuYfX1rERS+GB1PVZ8BWfirufxOGn9FbH1vzFi8bVKxApr3MOQ
pF4TjH5JPD1EO1J0NPABJYBc5aA/FWpVG9QeJ3t7DK/TxtS43WxYHYENVRer
0/boYsM2y1NcUZgCvHcxN+dYHAMxa2dLQFnL7+MWYlXs/MXd1I016n8EAu+I
kCRPBjlqv6l8uQy4eTOVXwCyqV8aMD3nncSA9bB7OHRDSOIm1fclkGqYBfj6
qea7lmqfRdMwEZ76KwNMC8c/4xI/7S3yFqY5mRdsUCGttABA0gPiT4+dEXwI
quJC4rSV/s+WC+O7sIzBuLJ085V4SolK0MnwuQyQ1FLEqpEGDr96zYplPOKE
Jcl4KmMoE/pdo/RCvZkloxK/oXw2zT/2J0ympTstB7w0ShFro8oqdeErBTwl
D6Q6uH5hKOdpDiot1Pe/cIsWAJbmLR6Jc4w30NGTG1vAcEyagJka9In7+jH5
Vx5cFMOdg+n6nG2LVV7UUI0cgA4Js8oxGI7DTwQNz1yZ9vTmVcX2Q8OLd66y
o7fgRxgyE5wpR+sbi7FkpbhoRHnv86nAau8fZuJYAHXoJO1E+woRggLEJZtr
sBHPRLQ4bwemfaK1iJeluYcujxxruFOt9lAc9E70wWelaocUGzDGLCc9413y
BOPoD9Eth6ujFUlDQ+642m9cHR4ULQW3YFhLQBTs6JzTIQzapYQBP/JoIPQQ
1RlZkWvksJ8Eoq+iRBiQ7ssgcmiwPRLJgFHIw/v4vCoBIC3ao27lfcKZIitA
C+BZFTni1cDCfGCnZQfh00pCofrYX31/wMea/JtGY+w7xLvADzYWp4g380hf
9/wxygYg/5audjBw7YFabqwNGYBfNyJvOyq67BJszQ/qBxsMiNbc4vgKEZ97
+F4hRNHDEFdVNPUjnVQY6MCvqjrhk+hHrGZKSTy3lBi1uMXUg2v0oeCoNv+D
SX1JrqMw3ozUmWIGC53tQen4CHCggKgeSmFGbgruRXGk94JOrTeWe3wcVhx1
sZQdsj8ZrHgjCKdim1hyexRZsn8tWGnSJK1w7V476z84hb8L5MrD1HRZ17rm
GM/xEg30ZaOu69hWl/C80VZ6GnBELjE4uPVw/hUSHQ/f9aO4Wq9bI5hUP0pa
l/cO9QmTaeyKdcf5ufDoVCsf3NGsq6LN26lyt0kezM/V+CAqgosSv1IYL+wt
Q1OMd7N56yFOXQJM+iwEEU4jvSxrEC/gxTJtA+zY9afs0Hfi7y031ygJf2Bk
JNUjX9xsYW5lODC7i7C9Vkku0vJx3z8JBW+K3oRUGXF+9XzV6CeGvdF4TDoU
ZuzaIuYEHnER2CkqbndqrfMfcJfxkD/vBNyOLL39IbpHrEh9A9aW+S4d4FWW
kf7Do11+oCVWnSWatfhw7p83dyms8NL5G84u872rEahpF23y3w6TnhX6UMSB
nfgH/gJMQAvRXkrw9Z+tDAzZmWH6CN6OeVnWedjZDBq/VUW+11cfKZJF2jML
we5ZyqGNNU/Cdbmnrn4i70px9oHcI4L5LvMZvUX6XpAR4j4tJ7KXNdo9oBcD
4oxIS3AxM6jvx9fNwedJyWzBXZVr+2/OJdR94WzoEp26XIH5WDe590zY2Hx8
uKOOdx6M+cz0PrkRGaECh1Cxn5lJnVGzZNAztS9bMAzvoOc6DnvK1qE6bF0V
WgDkD2V+d4LiP7RH8FS4xlfp3KocgmK5lYtkInXgwN1Bp6Sw7Yoy7wuMAy/P
pQThg359qiiXWjtF0w+3yc7pmKJrrCC9reDoK7kqjJpp9+EqLg2RU8DXADq0
qKg/aU97FJxmzK7wYNUx4JCvYGXXr654oWRtPrVPIdZH8wVcykvmFWAwCUq+
27DYx+8waQhJawFSjmkUreO+OeNhsr0NQfd2wxKE8oHegBUyDIQ8U2/PMpUl
Zu3nlA3tYkXoRDviUzteNXfqS3RT6BWG9xBy3irSWgoJ70kDRfHg4ztO+MNq
+c32KsWQnp3bqlVW9ZjCO0D5NdESzJjc3bo3rknPoxX71TGBFjUJib5hStbm
PpH1YikV/UDnIQRCWt+x88TqGXaVm76gJrdraFXKt9mQTSdd9NFjb/VvVyQI
k09ycGfgM6dhMEyAZ8BbQWMuS1nwjs1DBasERtDA474GJ/NYwFS8tVhNUQOP
R6or9vxnYP3J8BB68xhV8CoH9Ycgy9bavHy97KRWp2LYrlamZi7KRp5ENAGB
pjMiidPSOii7fJcS+dQNpR7UIIiw1zo7437Rnlt1O0/twXWqZ/8RTyHzmIMk
A/s6AJbSlXlM1K7s8CZBLmCabUBYEBknopxWvglyVKDk25OVhOqwC2CT14GQ
2Xcm16OxMtCEy4iVPhdTaghkfgjB7gS189SZ+e3AVVn/ObZyoCKjZYwK4+K4
eAa05Elz5SruhktLJ0CWVc65IzVDvYji1QGduzVfVjczwmyh6aJZXGwflkVm
H1nPekNeTCMlPthCBMrZsBXk2IBM6V8MzlZ/HWz3WFqeeAtKjimze4JcIhyz
V7yCtU71reWan378KZL/LRHeLfM5hHEOsmWYcwWNSrMaQ1sh9eZ3xURVurdH
x1xTyjaxPACIomc0HdMQCL5r+BPAaQgIlnwQqorup5oQOCv8arAostJ8yI0d
eM7/e4VshRTiCCKWa0n5B3ubcj91WS/aHwXDw/BHOfM3g48QQXWC+eCi5NLq
qyVqvF9akAPL9kfRJOF+KtteZeDXruPi2Rp2oN2H8rbayneIawXarjrrZB8r
6aN3iX0+h1wky3CAI3ZPhH7PhS5MNgVUr2zTci/fMCijLUAufjnBJitbod3G
oX3H3tN+WYp52RtgHbkaK3zS2eoTaFNuPdlrfWVT16DrhI9itSIwoeD9MI1+
6rYou6kPfWJxjyRj8PiEaEwih8RlV3BrGeUqHrN85uIueQFDQEM9xf+FyISb
Fr9GqLbRjNUEtEBQe8Y1/BPJbddF4XvwoLXYzxuk9mdwearPlJ0iy0RMornY
oKYumHuvW2vc4SQN3LGIqWHi3wh/jq8bmAhRkRxWDNdPvPSCvKu96dy72dbw
vHtCwcSVKjj1QasOVXHCi5WiAvGfCuEBMPfijcd9n5Crj0lzVW/KwmL51/Or
P4eu3poiX7hOizsHnOgSEk52IeYa2XpfH7PQqKUjapELIXNVyLWKLpAXH2tx
Pnpob5N4dYRRfV7WdhtrPRHP7tlPL11VjUjpjCkODJgxyeJykz2DbvZDMOYs
eaxDojlZ5a15DG/iFMYBjhnCqp77kCwg27Qh+uLENxEP+oS30ipqSKlJHiJL
FIVagE+22kQSKQ5NDhXwGQEKW3LyRN9WHQhCR7i7aA6HZPJVqXMXWeNaiEty
BVLD/Q4O6iIw7Fg26q9ag8tKY8Sb4mdnQh5SW19T8UgmProblnUjZZ6KIcP7
fcIM8mIKJABKHNEaQ4PkfYnAXAMmCI8+Dk/RH+B1f36C/Z4MRDTYdjXOwlht
Ou5OrMO2woqKtUzpZRF2Wm+5OhbC6/EOEfyiNUrrtr3tCkVji9HJf1Jrjqgk
m++CSotUxrhD1fO/nw054bhOjh3I+iR9FW7/B7Araymdjims7QTx+n9FSR0Y
ks6Yhcc7yu3h4cDtSBBpzHWNO/sa/ZX35aTVD6T+YtztgAKqXoGL3T1vLuRF
UFNq5H5lSE02qfbjpdLJKaZU6ZZYTntxhhIa7TK9hnhvNYHqr00hleU2UoWd
FxvljaegxbBu8GnVdlcJWMRHfLJg64gsnuibQFDjy+w3NBG533cWhp1/zAnI
ZGENTVXBqFioLOrnR8WAMl9mDZmKeceViOORj3rbshqS1jpDv8JgS+VHsItV
+hd2g3wMwG8qm0cltXxlw14nkB8SYArqFGaTxEPiXNyoaNE5YoysN1C9RJfu
yARb16QYB3bXwjh+NP8nCcxdHhnCtAaxhF5FX0PQpcujcezM5hAWdMLtEqve
5XqdH6KcLbdELZyL/tFR4dT+G8H1b2RPhmtgJ1Rplq9qbmmvbe5YDu7GAyrO
/XeRsx2j6Wc1GqulbrUQvikP/gCy1M+1S2Dl13xhsfmZMi53byS4MuwMXO3j
SKBplmZij2wfXGB1194HyewqMWQqpxKe74awfbckQhKHsVoXqoTr2pC1Q9mn
cr9Ksk8tiWYJfkFGDlVmZAiXmkFSSul7qV5PyI7wCkSLEejfl4b7HZnnLUTp
P0VV8tkWZB97ndrXQeKuVCghNCyd8H7jOiwwgcpWZn5do16BHwDDD7f5PVZ9
2pNkdJMr25IyWf6Mm6f8vkPCK5cZuDJeyPk59rFAf+4+fiosZ0mYxRXMDTsU
mclmDnq+eS5VU5cyWJumpRK7OE8TkFnho03v1gVVPa26LHFeVHrfDU8oDm+q
MrHobGXz9YPfxwzc0GE8aHAwvHjYH3CSUxcfQ5pmb7v9VktA4zyEyzl5NHfh
SDXa4r1P/kizeNME9THqRmUMaqPwQgzGJC3HkDqxIwjOG+uB+KLYqintTo95
tzi64ofRvuVifDf0uXKQibP7e88syvWxyPh/CE9ylRfvnZwRb1hTG//MqPjJ
vE5YiZOqVvF80e9yaX8eheMFiU97yxdWc0hEFaqGfjG+no/Dp6MshA/Xvaui
ES4mmqi9Wwlm23tylWfJCgwagDcbb8e9Gt6apGMU5w7J3RzlUhcIzLgknxXA
Rsa4WcnxV/BucLjg77cO/5DxborJfwiveENGzh8KxgYXVoeJUtjEiv8Av5TP
/jAz/nuDvX5n2+K1p+lYzVqnbd02xb3MEfb6Yvv5IAaDH0JYHWvOlmOZ/sUf
/sU+wPRfPkMg97NYlYsF1XR5nx98dVIxaUhibzAD93B1nvZaODqMMQHTk49y
P8B8Kneess9+h3ppWg2JVXYrsPAH0uA6PM3uXabcgAA7kUI+XSg4NUjUXEkI
ubDviEMskITGZ+Y9Of1984xw6VtUWUin7T6SRzzDf6QVSpkeMXSjvoVyQypY
eJU4Y6xnjH2gzUrKZuDlPXuNH5l4b17VexsN/Drm3tugfpsgC2X/tTYlpNHz
HRQlFr8J7nLF1e15NXT156tB3u+5SiXqQjcnPCP0URdEFVrh9XHqv0K52Iby
bpZHdapFdm1JsB2uuvvKHHxMX0rpmVSu98A12N3J1Q2ba7fdCklJDI54i8AT
UAMsUOzgbFR4jkEv+heG1yzwIJDcUXjHwaru+PTX5TrRrC1D4azv1R83pEHW
9+pcbv28T3M5k7Bx96NDs+wvmv8q/x64WdLu2HF5oAHwxceCiDpmpUwTEDu0
iuxuXLbMp5AtWHeeI6eATX/xnd0bEXT+jaQzcXQDnyU/j5PvvFd9/6rWZoEe
vtJ8fPh+xcDKT+t3FuiAXa0ajD7fXPoAncEgp5BX2sLwFlw68RH7WYkRQagW
LgOcT1Usl60djzvLZHVhcSOQbRKB1Fw+91ncVP3gciyH2DxsdV4L9jY2XueN
O6ikMyugwIZzSKUM12ZLPqW9j4nlQlXv5bHblNW3juxVCLaZ0m94q36lFyIT
/ir8RTap+6hh+QIH4/gGYa+OwoHF0F38GvkfQMuWopNAOH2igSSJeJC3gS+X
rQvASKasLgc3aroxvqFrNjXSA+yYfChZEc2FaX99wxgkY2ucvpVMkfzwzhjQ
qDt5uAl4NxniEqlhKUG6Lnx3AURkTjJMNvhNhAib4SWrqSIOvmk+8on/S7Uf
IpgdIGrgTTuHeaeyaIMJYmskn5pNoJ3daic5kePM7gtkpDrCTqkWRQChDL9Y
jM33GVGNcujxN7Ah3Ggh1XK+Z9RKux7Qr8mjszMF5SzrLwxyMy0wJxLNpAzZ
u1ObzGLt6BKXAx3QQj6BndNI4+1TAMXSu/5AUcfF28pQ/bSFypfrCr0AHdEl
tDaum19eRO66Qezt1C7w5FyKDez1pJ2TtkLZlT+GXQhbWM954cR0roHw2pxq
kGL+9hdBxx21NnQbudo5kfdtFVdG+uKmFJIRomR1mB4X9/punbQ0LhsEPZvG
jt8UC4kBvI3a6bNRyP1FxyQ7gJ0NCcsoy+Jga7X6D3DEDBS9hPomH062ZEYm
TTOZySoeTM+rMBQYteOYFYxU+r03bGwCv0sc2PE0Eh5skHhdlXbjXAptmwin
e3gL7XMeLTlJ+M3ZFnIf49vGPEHMx0W+2v4hOPUgtMU3r/DH+yfIQX+A43BR
Cv5Mk/KKHOsK0TOZa8qeVezjRW/Y4GQBuTI669vh5EIlxRGKk26aoUIKjqSB
M3Mq8cmuHA1Gob7idQmERABXn6h77XZd/ZKsnw1OhQdCVpcMn06Yzq7jV8E3
uN22Uvfm100wkEsM6U+SaRL+NQsWkpVjHvRl5pIMc5Cod4Pd7ktq4DQx++K6
Db6izCRHGUzVw50F9svNx3EBmju7ak8vRMaxRN0sb9MmSJXaHWF+IWwQ1lux
cB1jBD8OcH6Jt0/Xk1s1DExa2zeNyH5sNrMhCIZhiL9hIf9dDoNkL2PDTe7O
vrng+pVDX+YaQkNCA6Lnk0tEJQJAxXoOpKd6yLLAB0OWYssCzJ4wZcBg/Tcl
HNe3btdEoe4RypFRKOl84mJ858M8SYyLDQnEU7i966YNRl0B5VtvM6unODYZ
vnmyslXmUvGn1R4CXaUGijWtKctTqD2f97VuifL8tK4u+JR77oV3R3kOufdd
RKc25HiBbjfwgb+bSTiKlf3RBP0yRcMFuejccBo2/K8gQiwzlVg8rwrM+AJm
0kJ6CebSE/ByPkX9b26shVf9SyX6ohQb4CVpmNkqsS832mW2EWwmYUuXkkQM
2y64UqAmimffy88K3KcMxCMR/MUmAZn9SVCJJcNSH7dQhA2P8gauCtNMcd9u
PG9CG1v2/HqitYeuo0QAtgSzZhExWVpEI8yeSfKMw3wCmifW61fIxqA7zyBd
EyA0VtcueQKocFBZrb5h6izj8TVb31oulGZGCiobsYSmXl/YotxmChURiDK/
usE3g0dJNV/PGe1j67W3XNGZxBMUU/A3zRLSI3H9SBuYR0weGnM7gI6Y2J/J
TzFqDMfFmmoY+1+PUoLp8EU6fIoqn8+wVY8e/q948euzydWTgJhIUmOKQ0OG
agOeYA/m+JUsO9YJQADzlY8YJp94suda28wAiybwC7iptQRyJcc29mBdjpqS
W1koC1b8yD3arwqHFAN5CjY990OlcfdlCf6PIEK2ff9cUxY8LFwQmsWEJ3fP
ZlwBH9coCRW4S0EullWLb7F6ebtEWu2cQAOXOiXs2IYYzpq53apiYigMMsFb
jhIhzG8SlS6Tfbbakb2ro66/Rv7xQk/G1uUYctU/GFSUG8NwmdmBC2oj7N2z
xXwlzx/DEFqaBXVo6xeeQUIOypeTU3RbecEZHzYAQrQYwLh/XILm7ERGkuPo
QxWanetmtr2JHu6zYS6Kyx/9dcVw/CZ/wFMDawQ9NKMP2/P9J4XVyPgn6kSB
0l36d9GYiy+ViwzCDqQzlKTsraf8yw7usxlj4X25Aw6x2q8QeIktI9X3kHtN
whbrIykjUf0j82QArh6ekat4a7vyODdJMPweqdwcrZbXb7o+Z7sD3y9ZHNzi
1W5p9ZDWAfSQDI7WD+dEMiUBJPRwvS3Jh1CtIctfa8DCWxQ37OHkhUNt/1fA
BKXRDNDe15oLydF6PrPSy/ij7EoZguaJRv1hmNge/YwnnBNSeu80RE3MXmL7
hFNXgZ2TcgDQtjEACGa/p8pQUx0s4AhlIIk0ZsiuJ+ePkli2Vo9/OOjLKgp8
o+WZVOonVTnkH48aHBfZNcrrjokZvzP9PGGSiH0IAkbAyjaktz9Y86gQHiUU
/tigdtd2VAKh3g3IHbqUj7ilzdx4KQWTikm+guFImX2pCHSX/NqT92SVoGGB
BnJ2yQj+hjNCERpLuig3lh7+MsDXJQlrkisaqJ88GWJAubtrY1iN4+DxONJE
53xaQqNRstAhrUTB2+7d0I9h3hePSw83FSpnN+vxD+UGXOXUwFnZrG/cn1Pa
/Ki8mosmbNCHXWMztEUrCmj+6K1AD1ntOxGpAgFu0f03XyDdEH4vkZlV1U/d
DQlKq7IWWGIXwl9bVfoPSmLUCTDmIsXAHgH/XA9nZbHmjWR2OG21JAfLFUDJ
TaZiUOtZETp7HOybQfbttSd1jAi6QwwrbEJ3np/1VrloRcM+K0B9yX7gBXFt
iTMpSRKrlKhLttp0FJDiEqZWi4f399q2qDVjiXk3n9Y+LZ/30eikdKXABMOL
HAu54hO2tS3z8oZk0DEM44AgHoXRDZM7VDISkNn7R98vpGtYjtdgt9mshILf
jLboSmmRFyBMOAMRNRL9TIwwobS/9rAQErrKFoKzwo+HNTzTU30hUifLUXWP
1ElvqWIuV6eJq9TcoPiMK1HpmhLAmOfuX6YUpN8Q+VYn5NSt89w2A+N0Nul3
QB2IVQzRQblkVKHfHB5VFU0dxLrC/etTvfcLrfs0TYk4+guEVbsLeo0/2nTU
gZuY+BmkVIau1Den1XbldbyYzoIQBuBws9VvDzv874fe0iH0Vcv68Ml/7tJN
A+Y/RTsej1lYeZSvLTqALC06oRyCeM7L2jLJHrAr61gYFtshbwwQ1MoORjvz
uhAGIMR4X/8jFGePTBfHGKNqH1WFj74dE+yn+wYVxunizAuWg9PdsH+7yNFn
3Tz9Z7+hu8Xo2SNYp+eUpoBLj1GbWDExfvvBpw1cr9kZ1MvzPB4yS1EfGVOu
uDxfM4GNwr7s3H2Ulq52n4UEvVX8zbJmUXFT51dixwzym5uR6UHCo/yhkC5U
BIkY/p4y7J7bEmkjq0F4wSTMj/OrEXMP8aAq/RVfnlW+dQQqZbibKselj3TT
m9nQVy6xx9dXDM5ql3Jn8MZm50N2BTxia84PMyhUrVVnEU7ZCH6j4I+GfS6x
wwcV7Z30xJoC6kOEAwLeQHAHj0IG+MsNq8f3IOLWu8+qPyWQcoixhFRDrzfh
GDOcCHKOs2W2+2aGjBNruQlybU2bwXv+Cc5SJrKzeVPmARWjQYhJZBD6vyXr
7i/YLdqo27uhAvGBwQJ6UnsJzt85xQ3ScwbGue7Lzh1ztX3K6FSo+nudrHC8
szr3hrv+ugBc1C4yM6ODr5Yg+mJ/lryfbL5V3VMyZ331kGrIJAtJkpFfyJ8l
bAm5SvmRCp04BaeIL7Ytp+3ec3ndMqcT2ri/0eTVy94tiLo0R8ILv85+Ihf2
vchj8HwPbc0ZLZjb8wvaMldL+UUL5uth1JzFRFa3jFFqS2x94VpatBDX7Ylp
32vkcAwwVaxKyRG1pj5SfMY7vEMgd8u8bJbC4nfx1XYdAih7ZQHvPrq5If0z
96IVEX7z0cHw8dbXXxpqcGXaopkYI5p53LZC1l/uFCaF5UP9vyUti0IJ9rEn
kiB3kywfkk+w3iO5ZJ/t6JOuP+vsq/VZC5cfNoui8lJj3UUIRR81SkOGhhKW
/8IpZ0u8J2V3wRaKG01elgRmohWd5mhkLg3nr43Mi9AqxzeIimvHrFpKDApN
dGwEp1BIbJccLvNXFtVNYs1dLjK/y6oZjU+RPrl8K750kYSAdnoTtOzdxTW6
R0OrQaS3FprKWiNcImEmQphXyS+BAHyEIjmqqFC1bzTgRo8WadKsqXiKZIbK
m7L5UIpd06/mFMlHeWnXIIinQFJAvf/k4uPm3FPbGlw/7Myq3mquG0K9QmNk
pmjKycyozJvfnF4yrvvFce2W8LOGeyCPnfYuRka0tsv9BY+k44sSIUvUgL6i
bbDrayfa4zv6NtEfGjdlSz+9oH03itkXNf1k/DXD3zW0iy4CPOatrhndmQ3T
vPoid45v1EYoWBcE3Mspw83C1aVuSzBBaqqYyfGRJv+LGV1xCSCOhcQmtNr3
xTknLVuD1G/zWK2Fsi6Qc3XLMEni8n1g5q2UX9VTHzZhKxzkgTRrytRdT7ON
ZEw8k6iwEKn4FFdW2iH/jmP6t1I/lTEbpw6TJmNUO7BTcXJ5qNPxlGgvkFR0
x/2zeu6mJVuE4Up443WFI19+6+DTL0xmgMMDtavFWO/9cs/96ig5L7o4i2mW
EOxfEFNPvpvq+1HalsvlNVc6qnpnBHTttgZZ90SWaOK0dDaVYU68C3OTATPN
Lrpvqvq+plSU6L+CrLNXc0ToS0gcdKen+/27aE4lbJuuxhKnOlW69J1XTtL/
KXDBZZy5dLmGzJk1BgxJY0jGFSOOcDaX1CRRO6ZaajBqNvEngDxzsRuv/IlY
nGUghzYZPf3/CFFnue/P4D452aix5hxzMWkcQ5WWPqA1ajLGdyjNJNbgcvh/
CRGgNQIRbHVMOM3/egthfrrqAaT+tUdXkzcA4HorW/7yfmXw2VNdc39Zkdab
GepAnN7XZ2Mqq9OfFDGyCu5J3hFUzVyVSZMDBa2zdbDu+QzCObOOhOC2oPPW
YGwBj/kd2CN8RFluluMILn3hFe2wnfMmV3b+OTSTUvFkRQFJMJqma3luoGBD
syynXJMzQScfXmzljzXJHeCkNxFYk89/LQqAU694/IUmvLy7sDiTGeQYvtyu
Ikh4i6lGuMMe6DfgmZJFJRKIK7IYOGYGAMV+kRMLDbBmNrg6OWsXj+eZS1xQ
oszpjksyhscgNkBzrgA5BFpZtGoNpblvxMt4RmsPpZRDufsEsku/jp4j12GM
KQgpS9kvB5gNbvkzWGdikmv/rCnI+HwK+haOdC/WRrow5ItD4lDCPiEutElL
qLK1E9x658xPWPorWZBrnEMT7YdoTa2bIw1bMFerTs60XWZ09GM0zr+bopev
MFu+39+F5LmDisq1zJ2JH83O2EAfZsYyMGrpO031T3GNk9nK8kijhgKyxuK8
fIuWJuv9qAKVD4hr3ypySZ3Ru8xEj0u6dwXFWAaCSxldom7azpgYwzVMjHF4
dPp5aIMf5SimJ0Ah6huRTsiVXs0oP38lHNwaxd8QFWx/7DlZYg8lxUcNR41e
h49JUmgFmMkYIvmsdskEmIgG7VwoA0h0bmBygduuus6fSlGu6V50nw2HksVo
AJy8cBnc/79e/mZkBOKpK2JTjv30hFHq/ftmYGFSbxCnWzvb2Zq5dnXgadeQ
3WSNkqGpwa1t6pVxV676xEg27jtbbfmv+VVeCm8m66Ma6hutf17k6nPcE8jp
dTOBXS/lqT/222tuRoE/DI5kreNGoiW2XceRlLLPrp12i6OhoP93k1+ys5bj
4tPryVmu1EYRitUGrToy2G2qW+mXTgrMELddMScbAJw7f8k5xOZzjBfQwlCM
RKbtOAl/m+xuF/BybwJnW0HSHJB1Auqc+nbdxcj6fr6CZrJsR3gtllr9AG52
uts5h/9eKh9fCzSt99Qqk00dy152zPWyN6KcIyNNgXMsAZjen/ixRM829yMp
sK1Drx+rwEUHenlhWSg0EA+zkvnX32K9s2MtGLkZptTK1SD3nZst+/2G8RPt
DvXkAqE8AAXfoIAbGQw55NXSkIRQVjCACKs71wRA4rj0kjTNiwGx/pDie+QU
6ssHWNA6SAbCKr/SqyNchWbYpNR2QM0Kls0MEFzj5ZtIRuJS6qc7qeyFq9gW
qQ/LW/HotwqbRqt9FSHlp3IZ3L3XurCqikIzNcm5TZiRZ9j7v9jiGhgeWNmE
zx4QYcH69eZ4tMO3SKS3HaCcQzlUVBdR9u5f4b/FQct1yN8wfI0/PMQ0wy7N
JwqWjncHZsTW5K/YLoeCq8p7BfbqmvWHGm3YqZSsVFysYq/VpC8C4InG6WYm
HZmnrTBFr8k9MNS1Ryry+kWwZmugiRLg4jkL3kYWpPLKdcX5WzdWM7YEdePO
r3sSFoRrJAr5ZtwNa4JfQKXOHOBKzMaPSrswXOhjt9iu4Lk1bD5UYUtpEGBX
Ho2Y5W1gdg5nTR6WgXHWLzuYFs+VPc3HmkpRZ0LvcRT8bqMIO9kKZxcQ0bso
7V7p3c1VyZHY5M0WdqHR4k5B0qcFdTPiUrALFFCgH6oe4Q5/c6RnsFx4YqLl
s0Q9RcpqV3GGLxR6FrPbst9ZQ6eJR/PpK3eF7oYL5+b0xOafD0sNPEqvAFtg
17aCqbachfWzu7sWJtDFVvEd8IA3vKvU5xTSIl/SCd0AodZt+y6+E90pezli
sWpJ2gWXmOFUnED5uKAfbmhfsql2mrch3LlT2Db6AlkTiENlhXHqt5WP55n9
o/riGImiqyvkgw8d0btK8SY4neMpnn0tZWZxZN9cT+CFh2ZaAL7LCS9tPQTo
7spVoexLPDDdxh7Xb0BQgwZaDymXSlUB7rqbbfNpgrj/y0NgYpO/HZ86tzE8
HleTwcT7GN/LCf8M2wFbPAA8thKrFH4KeOfXZIJzNN0m2m5GGHqMmm50sgu8
3jCwF+e6GDo+Aa95MkMFsPoCTf9f60xTWKKBzI4Y09qVJGVAadxIrA+1T+pH
croEFh7UnqqHZKmi/0ZFZ4Rr2ZTs67uZrMMsRPPFrKxKDjfrdo3Km6ruROr7
CLhk2ybJit9NHMoPyd3rLObDaFNxcsWpERsNgfpmpYSRGRZO/tyfQ73x34fb
xPK8TUdd41nuILd9nNqP9rbL+W1Y65J3iewzn5UxxUF5XvCJ6MgnTYpFDRdK
Dv0AfPVg49d0oXDN6HnpzdNXpu9LChut+MWpbeqrwYRqW1WcVTVUXGo3DGJq
THd17WgkkhN9lUNbH7VE41nn/Zojce+m8CxH0gIikoCs9kMYKoexPmJqcSZK
EmpcQ5vIuVy1ZDglLFhscoAM/MH8asFmxxsGltxIGys4tW3AKbvXWzQAE52R
XnGLqvUUurrgL4KWbbsfjub+u4Ew0qcEvHF80mZVWzCllkNKnvBgFiBq4trN
WQPlRHvW9uo23v/0WokWDgA5w6lIUmMhz+2k6d5obHlhM6hWIAMbqhFNpx0m
YN/gkpAEe+1ma2pGEgaMdaxe7VM3qZIukXkPRCBF6px5FkSmh77PMg0WIgcm
LxQyIWHaxllyrQacrLIcza+mZO4Qqd0QdwR83SLw+RuTEqJQfwWuKW1olHAV
JJyxtfDLh/dNpVd5JOH0+q+6mJsqfhIVGHs+K/1aPqoAa5wKQ4qja7NKYqtT
wT2QiAgVlz+MaQXqKw3uWhiBQFOtNtvhd/onQ1HmR+hJmr7TuKlhkdsYUNlL
IGlFILcecXrCi0G0iSAk/geNg4JmtndSGNrW9WrR5N8wDdw/HHfdzumJGptZ
GMGAbG1yn2KIQvlLGjmMNJLjtkRp8dXCF7u6b9Ap1hNyJ+AqNDEe6d6CDl5o
yPBcixs89qNXd11v1nCtOKSAIchBxO0vBfolPDr8vLeGitdqUt2dIJlFDVZM
CJRJvSUXWbLM6oSI+sAiavjRwSADYBsv9fe3t7+eNmiOgNDSvqSDeDdN1jCK
twocbpLhAyayfrnJwW7+6Z2imZw7T3owgaajDtKUHjVJ7wIWdyzW6/Qvu9g/
aNuZoLYQgEsxGBXAMWa+4BGAvn3CneNcyucjxByc+IJKL79mWAjcvoGmromg
c6cImI9NPdNchQpXcBZaCiPSwrWbU8lyClGyUCYITieR1nd7pLtpa/AwMo0j
BAXBYVvaLX4Mc48LD8F3U/k92kwX+X+1pS239yY9YT0INgR2YIyf5YW45tp6
TtYNT8H/jlxohtwlcWWgvTRKLrktaXmAbEdoi8YgSytJaxpXOboGnazwE/dP
pdM3tUbTzvo6KrJHCEar61mCoHJzHvcXNiNxm1QyCIHI+WxB9jq0n8vPm6hw
NyckLMSSzhe5U5NYogwShM4mTmZ7B5WEAXgWcTF+YLg1UkqoMRz8XDujEtiu
o8s9RGnXEE56P+tBUfmEOT7bmVArpWuMCbY4pSi9fHFEpVb/liFYRtuQ6EkE
gXvqOPkPBUFznqRwoaA48PfPzNZ7W0E92LGBgAYTgsHTDDE8/pU1yx35+p+3
n7p9aW3UEqptNONAUelm73D69sei9WUW5dBc94c1Y+a8rR0lkYgGOTv1Wvw4
lNYyZFW1N4C7wLOCNjnl/Dcf4P2fd0R9GvqfZNI5PK6pM/Tv5w9dJYJODexd
kfWnY8TPWjin9V4jbMrRRGo7jpD1PBp1PAYtfqhw5s/+/lo1c/qCs+dDtYOU
bTqRbhJoEwodfVm4Rn8R+mgOwsn11611Z9cTOTYSU/CDnDZILlAbZM7yachF
QQymV3OdIGA/w3K1ynpANW71JaikXQcfSiJ5yMYVNsuoB2ojWNkQCNv6ZqWj
XBYub6+fHO5Ef1Lt+tUK7fEpsNmq/Um1z7Ex/1e4pldCbeEAGLfMFd2kxYqx
NwtwVeIVMtTqBAbud3AHB18ScS/vIh6gI1BRkQFR4xy1RHjL3+9gqRkhDDyJ
JKVUJSu/s8eYlx0iF5NRlvbzjN99f7x40dBRbmVfdUSM1xDGIaj/D0XzKMDx
+wAOHhNQBQcZprQ6/TsR0uOHA60rmQLV4zsvqfoS58zR7upiTiUL94NjeJGw
6fIanEsWLFsVAiMpm5JJwT7WKQ3ThQqaH7ZhgLKm15v8H9GidgdWTwo7q+MZ
e10kBCBOwRknGXLNlSEtAco4zFF9HcPAjWnAQkSI9AtJ56DFd7LcWdkhIenR
HF0wMkN3ef6lmbh/yoryYE0euYdoXzW3JGk+bxARJzQMK5DqGxnu1chArSC7
ZWwuuSDgdSN5pRPq5j30MNAlj3Fw3l6kPiOA0NMI7bLZunU1AV/v98xu2q0r
2wYSrEPZStgwAQIJ6SREiJDnX3QrQ6EYkqrBEIBJYIySx+BPlJcB87IDzTia
Z0Q/sOQKF+M4aningwCjOpnlWi3g2xBNsTzgRxrxsJ5rTJvicYzJKkO5l5Gr
pCHYHF9eevHwQFPjQWQHdldhqAZhoqaaZ28GfRU0MSwiWKqOuEmHytgtw7Qf
3s6rRGjsntukTpOVeEBpnLubg3O9l6lr7oL7uB+Am9FJd6Q8jmNACoSMHMQR
5jP5NWfjE/yGqsDc07JuSu66lCEt5DJTUL7g2OMEyAXtePkSQvsDMbvHBPfY
ZUR93PhUGHIEHWPim/1VtY0/2p4tlJ8n6Sz8rw6nsL44eVSpXTybvGD2Nf+T
wDzQoXPgsfQGaEgVXNgTl0C539TjvlTMgqWHlFsNLOwZ9DxSwRUZkmZglIvI
7h4uciOYZveAyouihvZVdfuczX5R6oZb9ZofIseIfgoxnYmjjGGSesRRhTN0
woj9kH38lLmn6j83Etkc5j5v2pUVPdL3F36Hk+4OF1yhoiGdULqCQFVsLj6Q
RecCV1InqomZ5/eTr2JGGeNGcx8rM22Ak9jeEedxCkeae+NuEn3DK5GS0XuY
7RNVfzoZiuvE/Tutg1yvBHUIBJFlnLQQVKxcYv+faL7SKwn9PrbMXbVZ9qrw
GYuAycBgDqCjG5wwAFc+cTjeD8+5Fbq8DzInYvAdmXm2vx1jQQkwUPJBofzD
8SYcyPqMOnncR+rpaRNRGmotWJ0h5ccAzPtBngTL2yxjwH+XDOQ4Cnfm0NUH
nkBS73Op+JkpFC44iY8VeeY1dw3DfYlgb7ov/WAptGudpY7A6yG0uMR9R/Mf
U0kNsL08HBzLExpFCrPZQKOfz15rWo0WzU6xu/KuK5vxzQgFnHRgDKYs5tFP
gTwfc+JAn4W4x5+EmvAASDouTES1yW4f4777hBfWTrwhNRrfcnXUxMUw4BIN
y2jYcOCs2zRi8YTLJe2FeUAsuKUT7ZIxRxbWVsm3tzVYYH6XSCV7hoRL9wPm
bUxX2+ZGO5K5C5t0FA0+ntfO2C0rUiy4A2BC2ul8az9JV0M5I9/ll1zH87vn
11+tnt1Mjwmbij+kY+T1X8wsdpDT6M85nA35VmlyynuHqrPvdLS07hp47V0Y
RbefyDhvkiMM9kOSyCVh+YRqIzUsuH97EIDsk2Ngj8TRrFW31zTIUsXHx73m
n1KEnpxVO0TktmBgoR+ON3/+SO0GJ+LFK1qpB+L88crhxl+8eJ/DJd7DjK+M
xtpY23lYgloWyK32JxvDoy+1YGoLqt5CLjvioytuxUi+kUaCVO1ZkEQU4jRj
eCzlb5WoDJdSwQTBoWNESMdqfEDoRYZFa60QcbIHCFJSWg2vLwW/rf7TbVu0
R81D6RX3UldLCA2Vy1QZBvhzpcIVATMl1pRhPPz1V7HZY+LUb5HoeQ3bpzBQ
sWXEm5txQqGtJerOL3UYE197Ztjwv/HWe5FS3PZPyjupp+lU5gkFseHKH0Vs
PQYnqVsbEndJpPBXu4z08Qvnj12xhTTFWqNK6qI9DyCd1ixM/8RYZ/yvPp4H
2nB7VSO3f9j3xxVHiUEyaCvDc6/BfDs/Igv6e5Bf0TN74eVAZfcGIjtxasS9
Ag1XIqNWDMPORLfXg53VXWuVTxAWoB+PaHvV2xL+RhQuBsGzfYz5kwDOZTfA
Uj4qCB/hm2S0ySa8m5GMURxR1tpD4GavMP5zvk+tXaT5sp5mGyWbcQhAAoBl
6LVbqHxVbJpmSRsnvsFvD7DbctYX7DKXRsbYh+lTLKYvfJsJXEAmrn5caVMC
OjLkHAJQkgDlTuE8PwWl7ATvxOIciLvGBK8LZzSC90Kb68I33zQQDoHX+eFE
dWk7ZRU6DUFfk3r+uu6dShOqgaF/jRAlm/vKN4leXuAeCFg4QqByfrHpNteP
8EwSbW47VxHEMPA8b4bW0VpXT2IGGPjVvopzpOqoU6aBG6V6D+5P8dn6EBky
0Fdc/VdqzHtvK98ScDnGpSs4bxscLpea8lQvKmTQAcHlmea4SJqduHOJ3Ihy
4VhKjnx7A8bfQ8VQDs7kOApXYa/6HONjY603KWhQ+XzpolLtBihCdxcAi88L
oe2isVcuATnYHBB3f129AK53MflSLCJhHrPWyC8DjvY6BzrG2w7ag4EFzXqV
ptJPdGoRZhholRbF9Fpybemz0QFZlfs7mErYAY7rOhwHzHsfmH4B1Yzx/D81
HgZLsPZd4i1irvddRjMYAVh9qOVgmvasOA6b5MAiVZvn15vzCuaSrxigSEGL
1exjEAWw6nxMK9ifvdyFZbKZLf6Wt18HqY00Ylduq/o+iNXmzx7g+udCCcHO
mk3EKaiHpguApaBp1L+lKdVHQaWyhvnpXhTzE83t7xqPakqUIrlmy63iRCEO
A4TDQ3QY2Zhi3s7avmaTzALnCimbdI9q9kKrajdFF+wPsUXOdp5/rrDSEOmI
gR0/j6tiNQd0F3EiMcQ4F4lebkSFlkjRSEk1jVQ6vj8fv1VOWywVmk5aMk9u
AcR30OiEH6Xv/UCqY2PbPCsutc4/kUcees45jVFr6dwTpaKn43GA1wxup5jp
MwZvibg6AVialJQylqJLQt3F2yLCNG/XDrGqoyhg7glXgYOG2qzsHyorBxv9
KdIxgfSE+AWWzu1NCvXbYgUua6HtHXBbbu2rqzOJK+7NZgbWMDERfer6P6fZ
/fNAR7qmPBtqD+yCrfwabeVa5u2fQeLMUcYkxAr2u3wR8ix3wloJsYuZ1dW2
8S6rgmeBj0hL9vhvAFpGrVxF5Ikqlm4jxq0HfJqORck0oKGjI80m5AQhGxtO
180ln3LeJF4lx3Cl6vUyjgqVGOULAzCMLvzRjhzTx+WwydT4u79gfZ9sYLZN
9bxnwCmCmBlMH2MGjQdwcYvaAwAxTvP1jxf4Zjspj8Pz4Js5was29rjhlqZi
6MNBXvY0jt4kopnfK7deuIEaPwAe9MBv5RG1r20caZduNwy5aeUpFrzz4DEp
kIhUmhv9+tH0tDd+gTorCJtbKK9qZfFtaH/2BR8KueC3w07+19uU9JxRo2Jw
gBO8ZL84Di08Juf77xBkMNJqHLfQiiRgAM9laGK6Vx1/ePK795eyy5iFiUHJ
qeCr4hSgKn/JoNZpWuov42932Y7gpqMMxeAo0izdCdZAz3ZE6SnGbo8haYFw
0U0KyEUZJpRbrEdbZrqQ122/0zUUe/J9iiXcd7vjc0tApMZ98Lq8/3dNf/xF
GT0LrlfjVeC86gpyshCgUE0EhUVerX3gQuSLK/PXErn9kHI61fWGhe2KYf2j
c1YSMt/WgMnsDi/kCJFJ6FLkTVmUuyJY+SjIs9rOWEEqU9Pv9HL8h5oc1SZI
7e3oAm3nejQMRye+amvWxXslOHA0MHsvFb3mHuRciLK3873zOJa8lfI7LtTs
1+PfnjD2fX3ih1NnwcVmAH68sMJqbTx07czof6FoJTawBYyGMeEeArIxntWG
jN5R+XoPFkZfIkqn3kf0XwuL8haj+kQw7Q0FinXT4/NmeGwNVpJWY+rc1ZC6
F3H3fnSVEODc0EPSEy3gjPivr1PBxX1H5DS+iCoXusBvY9biIGCmFkLAjTSw
wPryytElZM53/d9oRNJeG153X45l1LMdjc920m4KZrMdQ1tC43zxce9G3kg5
SIPn5F5t3FQ4d/kBCIr9c+mnoerr5PxI7vF4/086a1cK6+pL6dm1TZPGIBHP
yzNDzYJapT+NKk+tY2Fir26mwjwxViwewO++sW0qF3fFiX8SLSJR0l8oYE6M
jCAZS7F1KYxqOZ8x9OtouAPINh0VF0To2mlYBp4IPCG0Kur6M2mhQvFYEByF
fJGpl2JkioChVp4YXUtEnCzMgABJtBXb2HbXyRz57/0R+9OvtbMwEXKzJAP/
ufqnwIb0Yl/lg25BaOsk32UW3JiSfw3cwmK+UyCE6sAEqrC6+fJnLNmlXmkM
/rE5OxrCl7lgePptV/T4CqSq9uwXqHwNlkQf0ht666Fl1nbha+P4tRGAb5te
HmRAKubyjVi8bwtACVGNgT/7F8DLleODEIdPpN6lT7lI3mw6YzCIx25lrLl5
7DT0hd2aEeLes4fR4yyyuVgiZDqbdl6ZuDWPsxDoDJeIKl5YtpgdNFPxXrTA
XNOcfzs7wD3b/Z1bIu5iuFCDKEVFIzH4wY9T3xeH8sFoLpU7Wreolc8PL3KZ
pgo0/hBSdp5lPzoTK23VSeM3zRVm9vi6V4hxZRQ4QQpMnAy9kuPlPlXzLhla
o5tuzPM+msl0c6/qwQMtaA8JSKBOMsMh1IGjCG9vYL8IgwYXDg3R2DrXkptj
bleAAT2bRCyjt/hv04gHl3C4AYGdJKj/3+16mWxl6bFOIYCUrBHsnLb0V1Yo
amOFZoRhwOoCeUSjz+GEXJUz7L8NVFR4/qyj0aiJynY1tmT1IpmNr/CiiY78
kv6dJL5runIOijYyPU0g8lJW2MfhTRJ6FBZoZMy4MZcqsa4TPtQk9cvEBT/x
aYmV0HGij4O649GC8j/cvsjjokofll1LtbOOpYQsmUflc2w+whhDQhx4grxy
UDM63kfFtyJ09dhkQAlnamXVGIkTXAX0um5x7RpHtrNQsG85axdZ5/y+if6z
fdFBUrqcW//ZWxZQCHgOFx7Fi6cuZC7qdANolUodF9O3G0jce4bXWWAWWilz
HEvmrcqu1F4ZuImy3S7xLMa+2tds2IMftwLyzY9jBmnO3LRWb9chv56FlHy9
0ABwEt3D2h04x/6TZp1hBe5rEjcd8fQdF0t/W4xUM4bLFUfQjb4Ypcfwnlep
+nvCdYqTusXunmYL0SOyp/g7gy7byhvLCN8P6DBdxZx2IYTYJiO+e0/zdsGU
BRFGDlxwDqOj0pqrzubWqJwkXVA9xgIywtdnXIS0H2+SmvEKzuvyBm1Ixccj
tgt3gtXoQ+jzhmV6MyGAfwj7c6SRBES/DKJHnJntZvDfHvuwcaSDelqRIVmS
Q6yYid8w64S8DeMKqkUUISStTw574NdCmgEOWaqwMf0KfK724hPrnXyEBC8v
faYSqUYe9b4qN/KB5Lwd9RllP+Rn+C1vuXQsIdTCeuCrJ/Md2w26Bj9Uav5m
OhB6GwspKF0l0m7zP85QaM0sw/fUSniwRCsC/Pfa/i9rGpD6ou1evaiTkU0K
haBHyLRPjYd38P2gaW70+7lqDomr8zD60tLQD3kwyCUixAn/Hik1xbrHBoW7
XJdWKqgAJ3CPnLuodWLpx3xOt0Nr4+7yCwu3fF1ct6gMpa0kS4X3Oy/h6n2V
jv7WReMNylbOmqxW8uRgFsm7FDv4Y5cOgBqg/M+D7UjY3zN40KcOxVjjCVCJ
mcUdmMi/UvEWY+epT65YKqnAMSZKsFouDokJeLlg/ChcNoQI5R/wBp7rTtt7
0nA/q+HjsDtSHnDPPapZw/0EwSRI/MRGjwLnGDpMY2dEH0zpeeLRyMgCm1Yw
ceJ9wxlDf+yvktzUOnkNDvvrq1RK6ga5AfLHEXPkxBImZUTlNIOEXV+UaDuZ
C+6B0s6nGRURpUy6X8lDlWWSBtgxr7CnQt5LDBLpkP50eKqa3Av6Ed1mcQUj
EPX7kqZocRp5LcI3nwGQnPn80GJoeHsTsuX92t6g6PLm3bDIPJ6u7IkhUsR/
Yrb17sYt6wTYI6olHwVuj5I7+blMI2p4MamSnxVYYllZ6IijtgsTNpkdLRYn
cdxVFXnxir/OqWCpPNwa0XXp0BDUiR0GxlAjkj5IOxowFTvtqu+ZapAxnwcW
GLAlWAfmmE/mDMVIHAcH/zDrp79IDlGEEshhau4pxGKPjDL0YBHo/Z47nv2z
iB+CCeN795qGk2vAlHZjk3WXFmbwPW1Db9XPLtTkQdHuBGYUF1V/wiEf+ghC
M0OJ3IO02LleALCFx8HEpgswkEESII280/DFTAwrExI0vEBLAOQmDpyoUZMv
J4IzK4M3hP/FZYU3Yd057rZmNyliWyxLpHznED2mDlOpISMAQNWzk7pZNsPc
aY1b20mp0ViQG3XdgvDDM7rfO4r3aNvy7Df+3+laaoa2C2WAHEzZMRf0TVNz
0sLYYvP99gGazs426HsLaWD+caoxWxmrvhAmg7Fcdx6jq4tQ5ZWTMB/q96ZV
ve/IUiCndGsncHwMyr6EgDDiROZb/0wJFmKO7J7Ih9/KklhSf0kkD4ayxDi6
hA7kTErO8q+0zlTOpb6O8N4J+M5AHCG4A/X2vhKVbbF/xEw+g9TeAnOAcUTQ
AdViVHjpx9xdlhrh64ONFmRX+/onr3gaMEy8bdYeEijl9skUCnh6l2jooVFj
LQt2+/Tq/D0szB6RVHwYndEws+wLzsy8GRjcB5Tr/T+KiaDOXQ8vJm+ZtjJH
6K7t4SvtAMmsAh/bycWBEljpSYx3ce7twEwiqGKJ+01ZeRjqVOcInRCdBSRj
WqilBOsRxTfeLq1/gQMJRCiRGcLduu07zJTAlgD1C44EAWaPv/449RDuVdaX
3wOYmEfyH/XJ8T1BJZ0wM3SgZOCFrQf7dq2smudHp9gcNO4+zS9yaylWmbi0
m1VMbqTEh46iCZ0946K4DXkBRb4jekka5HoohogLGS65n7PNGMiunwMofbJn
FCPoBehbicsb6hUQZml39edxJxNPLaIVWnwPq4rR61/JoWZWfDs2GTAwSTdQ
mTI0kXAsEZc5ClcZJzc8cKWQKMOznPmUYfki4QpTs0yi219uUdNXWdQSOIMQ
ToInJfhSz/nFbsXuhtnngWNA7blOHVzmR+vqI8J7KuQT6C1lbEOin8Zg1pMf
9NNszSdwFrH5mfhYsqRhoaVqgyCczg8PMoFqeN6Cmj0F+Yavi0ZJjjZG7zVZ
q/3BH4jHsv/QA6bbnG62ZJCJFLzWOImvuwQqnx50Dx19yLIGjEN79U+zKnpn
5gDyJDSeQsrVbAGzx0wN+oAQfFzuZkdM0HN+gP1OQ1liJM7TyxWLVvSfo1I+
m8gWDu1IOgRIG2okVMtFAdJ88IH9TzEcRbcs8+5yMyp89wfgY7MabBhntRTO
v5kIv2po9x96uR359LYc+ARjpghUW5TjRia074VL70+b3WS+hWoq6YxrBhgD
KYevweWERWq5ahkE0rDtAO4surKC97FJeygWoEhds6Hsfcme92NGlo6QFJnR
yHG0veM8sbpYM2Dmn4Epz5h7RSlX2NhHdfnhTcwOczlun0kTFOBKqo8coK/R
mGsoUSHe2OMRJqoW7NpEbvUkCBsuxzq19dUnIL47+cgLaUCiCuayLi2/4OAH
ZTXWzov5+U9nuNQHya5j+ly5utSb0xS7vZ8V9b2bazptEJlp5Bd4d4RJB0ba
VNJvY/KRGY+Xq3BuBru3k5DeHSzgx1eAobhEkgTIWRA9r6he7Wl+qJjwKhPt
lzseoF7yctUfbw6eclXnVZVBtp4V3JGw126UdqoPmNy+5faLl8Ib98gSvZ2C
zQaJzQ/TmlhIweVXL3RREMMSeOJeJwKiyULMh3U8kY4qsq5ABRl+7l5MaPhz
n2qJhEbR6hqbSa4a9O8hGSH9EBUgObwgz8gxr/v3NBNQCzxkMs6r7kyPp836
+z105BBu0Y+b4tjh9va4ofzaOA3YU50NR426ZNLaRj+OwPRm+AviBSqmNkpk
FuyV8QQoDs1Ubdlzi6iBThaNOhYphfEid32PhFaPyeM0aSdJG+WysybSwQw1
+wq3DGFk9Y4dTFZpqBVJK6TH9E6SeL7XxkoMJBbD5RZ7mV0txbRNS1u0KMIs
yCLJESflZksJpqlrh8sK4Q8SZhivbS2RsKz98Je8PD+xq6ow2dCjyf2rqo8r
ZB4CCTLCKVnhrziYuM6W2YRLVCfJ0BAtYdQeZh31HrspAaW/Di3ZM+oYhL08
vh0V3tclpTm+GlWe4ICkJNEVs9BHBq+o0s2Ci4uiNHR9KACG9ZKfKHtzUxx1
DTNBidfJ2+r5/nPAvLADM6dnQSbdWAAGC5ybasZUj5GpYOQ0h2xFyTKo19no
0+XA+PoAKI1dpVtQkhDL0zrpaBW318qK3MiJgvz5Expcf+2RBr0RPbd0MjQ0
DiMQqChBk5bKZCKy7m4ZW5cTPZnyylLBIEcyvSP1N4lY+Ht4jFP4CcfLyUb3
OFk6r0vkIviOys4dCY+eNTHtudvhs95zHjZOmVx9O/Ga7wZGWmV4vfJe2rll
VExPWQXQ9f61GTBfSKHAHqcM6adldmm5wZahC9UsPwPWoitXFjZhHFFysaCI
Rc3xVmwacotQqM0BjRm1rH1/bj+GnGSoM0D8OEjJlO3mqBvrertiEL6Rr/Z6
KJdAS4IIHo2T0TUhDW7Vqro7H8w9kYtaWf5kTq+EkRuTNHyYDwxUsp9xVOWj
BM2QH7IakY7uNHzOOon6ffuyKwsv0FALyCOU8r53TYyvUT+GVjJyFXUq/PjP
NKKkSrM5XysitNzDDlhxf9V150s2FYacemwimtCEkkCvmZFrCNuCrbleJ9MJ
c3qp/IoXuWVwWNcHcYn/Grl2xDf69GaNi5JmVTPH3kCy0ZstTVDPgYfFPwSe
bxNKNU2011N/uKlB7re3Cd+WoKlsPLfrTiq9KAkLlHRDOL10McQWJVCX5rOX
RgXt79hV4Zg3srI6VqoAhDrXEeOME4+v6Vd165hEuRArIKtJ6uB0wT/AoRx4
vs8QKl7lNtF+AiWc2TZNijZWGMjwI7Rmf9IcQ/dqjN4459gXOnYaRSTvSB01
vadly1dLj1MYd591dHZE0QS1yZbqnia/4QncY0Rd1xuvdCNcGNIAKT1QJEsD
FQI23tUzu15xzjnMswRlLF6ao6gZUuYNL2thTwlv4sdmnn0Lm/7mRkv1Kfz0
TbUlo61sIRW+01/Gg1quGHVuN5nEgJGgwpIMts+Das4y/jb3MaZn46bJU+qO
FYRdKFJewtxae49u3nJE9BRfekDTxHY+j3KIWlMx/QDzd/xzqPYF2zmY8M26
geFQ/S/flEnIp0DN3fNdaT3pOxdYds9fmcJDGfKw5kXp90XLQXmpJqXQPSmb
B+lWmksuK21kR2nZgvH8uSr076sEjWfuDqp+sfSZr6rYxha8Jop6AKvr0ydK
rLE+0gOKmLDtF+cHftYNJwjLGbM3asOh1pAtEdW3KJ0pwDboJXNfPNjjimZu
nV+k8cC+RdhCMQqlV4XoINFYg63fY0kKA+rujJQzIJU3BUd5sqbENcw502X+
rh4aW+z8w7l/cGR4GM6rt9o8d3V93J4FhRJs/evlbTE7SxsW2zd3odCN16qD
D1mVXjG+xr+vcZeuRPYsATT0eRtdz/9MD0XCHvuOjzPvbGige+pnrenXOVRn
Fo3llaHSXgWnlcQ6fAkqBLAatlXqSgqhMgCBbcTgHQvCVq7TzbyfzJx4Ptij
py016q1CIzA4UuLoee2sr+lkGfeyfFFKud3If7mM/Dr5igSx2Y+ovu78d4yt
QgI6Me1eQtF2VuRNAZfitKQPxszfSLBGpcuf+7dwV4ZUonKOFEb/1iipkOsL
NCjtnXDSuVtfolLn50jU2+OGqLtl6LGrCZ9RMaEkWSeEGDyFtm17uvIDfZD6
J2cHF6AEV60RMFgCkDWdbtSRLJkE9gmLn4GnL+4WS4KVZ+WGE9x82WGi7lCA
/71L/WgClK/NZJ74WSm+gvwEPYkEAam9Jx8LIxwg+Nt1lpSyZQzGcV8xY3A3
5mF+xFbLyHAl2EvCcJJYH+ztpThUWhgBxTNa4+L+ZYmpXy9+wVbH2AbDW6A5
73NfV4yLUJrYDZSBrsqo/TgNJjlU711wS8r4UGkvYrvWBcN2L2ORgm19F4jK
JE4QMT7iloUu6hxscOzYVreo9n4rG7IuEMVGKZvP7CM5zVhVu+lLhZ0g73pd
NGQ5VBcWGMY+rREZA9HATTOuDaQu5fwv679UmOojtzmnPCBKvMUcpN93hEoy
lASuTXpY7oSSWSJrV/RXoZyrT2CR0Wcc4Pm5JkMwN6xORpayymezlsvBF8O6
fcpv6Oup0/HV7sF0zRWZoKKqhzghd1+Ei1UszaPgLA4RcXHZzX60QUEen3C7
uv2SKAa3HZ/FhxlOD67hGUxP/fqkGRX8VKOG+8zSUTTKRDyBi4UAol38aao5
HZFk75c2mjJd9dyL6ckQJTqY19ecuce1VXCxUY8IA4Cx6GvoL9V+YHcqpbsj
BZkCv7ExmUNoYDPTi/ah1CaYrdwwUTUsVkC8mWCMj2feKpuXfBNdgpaXlh4d
fCFZ0OcK0j3kvf7PLtMZWvqVTf3hHZkgkeM9F9g7mxTujPYY3ftaZChsuX+5
UvNO8v7wqin98CRNPmLFaQJBRKQ4prm9leEtS8TdvRvQQW8az/wwrPas2s3I
jxOB1vWFVIcbmfDyBhL72CM9frMOc2lW6KzkugEm2dkTkdMyOZiGuocdLN3n
Dq5IDSz/IbJxpCODk8C3ZW94bamUc7ExwpyiQ5leK0fBzylkRCKCAUkralmh
lMoIb6wGFX85LWZwZq4RUjG/nXILYIeLWJyhi1LkG719iVAR+cM3nXXjwtyU
qv/DKZ4GjDfJlbFZpMmLfF6qchLbLabRBIDNe9F/m9BlrOxoAIBwBn8WVYZa
dfV15Inl8Z5nTWFLPczePZnldBDUoWndBfwA1xHe2+rxktrLKwkZ2/yz9wpx
jFNvrgXP/aoiSXbFsW4AsLBNU9XCeWbN98BlTzIKk6GHEOzy2Mf7N6hW3KK3
8BE2Ou7EZAoGQJoUO3Wx3JNeEP3RKOqKW9OTnTnUTDqUyitSC5crB3C6suCr
E4gsOZnJRLjsOPs79aQR5J0sT+Jx5MEM7pkIbDsRTDiES16qHsRDrj4t3y8z
UTh2TlYtmp/FEj4Rcj/e5n3r5GS5IIotxwqiquDoqXjXXQldOOo04Is+TqO2
toFF2G4k4Orgmus8dYkESj5IfollLShvmgNRLMhXH18x/iKZ1lPjygOSrJyf
ekf3YuEEHSTh7cbKn1VaPKFITOs1uocJs4+m1lzimeTABZyXyg3ASycYXs3E
E1AtNtZ9IgVV/lnV4pfUBMyjhKgs38NVoB2IYJA6iNkGGW4dRCRZm78iI/3D
oElgJHHo59cwPqwtPdGlPsCLOp0wNB/CKNdBFC6k+EepvWrYlrozCfXfUc1l
cftjVcedYCnwdusNDgnhLyguf+SBWuPv0SMo/yM5evrMrQ9X3hqrzopWcAb+
8Ho0Z3GbXe+fG+i4559pThZjrI3TdAYnpBmRD+BdBLO6FgWlZa1AEFr9KH+U
dKNI/KfHJ7rZ0+B2aEWYxDKKK1aDRUCduAu3uu6rJNRJ8wR8qCtvThyJ4ZKr
VTtyhrSbLv7X94Z6I1hm1cXKIopCU15N//mDlvX57RT+J2KhIkikU+ypkT2T
2YukQ1QgTFVUYOqo0xk4qgNp20MgviZS1SHraUI+UarZY3CxOB1v77FP+DNz
mAf2hs3OLMDOuTnBgG779r19oNmlFSr6xI9veWr2HqzSv22WTn+qqodmykf/
qAkvwEc40hEmpNIg7zuzFOfETSYRcjyHrPlQlxkZJXIvdw7mPoQUHdqEWHc7
d0oLcOGMwQ1tncb2N2xC1g/yw9RD3OJRRIZt70etwnmfXrJ1lohuaz9/tTCL
9ZFCBlDxzBlFGv+eJN26c07OifEUEcIyC1gbPM1tRYd/b+5MVs2ZbgqgkMq8
dCTK+NB07fx3IipGBSjQ1BgxUeVdxpRwJgCB8HdBiByxzLq1UOVmsMyloAhs
75Yw3k3b01VqGOlwgonK33kMLtYsDdnHc1CRupqYePWSnGYfRHVOV3kjkiVF
gm0kFg2OvrP/ZgNfa+6GesL3agYw/+4mLiIPMqHlfKWbMRj+7ytLgxzWI87U
H3BWiaElTS/kU8Yf/oOLokaICK6uyoFE6F1JPI82pNPwjWk+bOIXTDqyDgQG
EJHoVTn6Qv73NN121Z3NKB7oqhkb6YsYJpSgzSrtCdar48St0a9H87UyS2UA
71q/UuCMLVLOS4yib4kDa+UPT2tLNoGW6x4Lb8QfoRTvPRLlZNqxv5kPYio+
Oio2DPcHiEIwdtb6238ju5l81OgYVBDwFeoP8+bL1SWs7LFgoaFzjIca/qij
zLdHDeeZdSyOXZ/uvpwzh76uT4YSKw9qgZYuz+zhM8gzd5TQPD17dcWfjx3d
xKUZ+6ylq3nixO4bsQmSVDpacqxOYDQ69dtCeGFCHrQA3JSI+2F8dxKb3W+5
jgp9YudsRq3HSCa9v+Z1M6OtFp7e8u2MkK7OlhKR3RlD9HKvj3GuBeDGNp5L
p7x5u7oHBgcVe1amukRK6KrLEKaxPPSsYiqTD46VKxAqq1Et0PIgj+roOS8G
BGjqyH+sAv/EYriZV8v21a5HDCrRvLcM8CE7linn3iL2ypZh7OvFvLLP1lri
awdic2sYW3ypKzxEdhqX6o6cuqI48o9jwCWxVRJIGeB0JCIxcccTizSAPuqJ
7UR66jCPvppbxNMz+/Q4GSBPj3eAmKitaL0zO4MlGMTbGvgXaaB7kAqq48De
xtzfsugPlNnJPOgtU4M/e9wN8VbVu5wcoJH/HPDkjxSOIRN7vWAE1z8iCF3D
hA3bu7s3mh9AV2OySKy1tIKMX3Lz8j/XFFOVB3RIREhp6ppp5VhaTxKZVmez
d20NzOTPBw7NgUVaAjCzJUVPcTVyQE/b+NtQ5xMRjrWiCIUGve5iuHew5LVG
B0lAuvpvGN2uva83q9hsKxb3KfPgRBeJ1f0RXkmtwALODJdvgK4hTSJOt+YU
wFhwjHeN71msSc43M4qH0g2TBj27IWSt0zqmkpqAT5v+hoJCyaq44gwS02mW
jXGxmlFHA+EhtGBrfW2iiTxudCgEubws1SdrGfYLnDytfYOUQQeoEcPoSaLW
ui7LSnnZweWzm+6PTwuZ0MJoAPfgVrNtMHmKk5BQeIhPQAvJv/iVO4/suNnd
1uiOLx3VL25pAhfzfMib8P4ANiweak0tzPyJmjebK7h3IsiSmAIn8RndHd9x
jI4UX/PXuImH7t00wiCZ/QLVWEhLBQntLc5fyU5C4AXFYcDSYlChgVVQmpGV
IWA+4rmbV9uHF5XRloD/9Bi7QUWAe/BTrfWo5lPeIMdhV/1W0GoSewEjj37A
BdciZNNFDdhHFjK1WK8fXVBZXy+3WoGyvGOoH762t0A5crkBx1iPsuWv5GUa
Aumejb0U3ucOqLUl1CXlOkbqElBH6pYDaqKbb8DeP9ZDhmTRlI9Zkwhu3vSn
mkv1DVeZ+tswYPvGpx8aKAKGzn8DF/qombSlykB/YJWSdpPgv2PVgnC414FU
c9eU355URZ7j171YP37XfyRKpncL6a6UgoKhpoadrS3+oT8wXD0Ypqk3gRN9
NZuOCpjyi36RG7t6GDaAX6xWD4HpCV3UY0o//wfA30wiFrOKSdxXbyUqh0R4
NhKeTNYMnr56HaFWJIvhbUBvLCmSUc41pBSDwBD9azFMqHu4fNgzzh6JNK2C
BSpy6M6SM9cWY/uNe+aShG1/RYm919aQMNLpE1miDs2Q59XLw2fgeJl7plwN
+tyHD2V0hL9KkCYU04a5pUoXzR5FVwFzyYTpLZ/dAsxR3uSpMWRYSBbSKhBm
yC9si1Uf3sQAJZEhosmuE90MDhkFDlKPth1sqtcT3wBGNiokYbGFBsCQidt3
QiufdaglkDAIAaorPAWDhz5e3VCdX9uyrsNls6sqs2zqGjDDPLK2J78pZl5v
0Sfk1UGCLpAAw6YNJ+OhPUURbTRJAOGO5hhUMr9e7QoIPugk9T1U2yEBENn8
rWj8quy2r2PxSd7iunPaJoZBN/RHypygc8L/vBY3ypj/NyyixV7beTvFcRY8
IUthqpPBqHU5p1AFISSvtDBGs8ZPhb3Qlam0rKaAqyDx1AscEW7q7FxleutJ
cAjIoTkgesJXVk6tLbdUIVWVGaGSA1+FuIF1HaUozg89j7kr+o25Z6/e/zgQ
gff9QAXwcvxpAZBlWz//ilMChbw3RYDOpVoa0kmA+uLr+sHpkah/KQ/Ane6Y
gKQ1D3jXhxKdg5l8a/NloalfvhOaHMQsIOKUwCwOeraRGsjIdXvkIMIIssLR
juAeGgsv3/QAP56jzzIt/+yzDSITgsYFZTHyq26JMQ1cUscDBLW1OIp/i3PY
muGssXiCN4pOvWDIR/VjwqretpPVle4PFmW8BZ1teJwQp9Kk+XxUQ1D59R3l
rUr9OEnQXHRpvVCNr8DfO9DJZms68w/OyVlMsAn6mVfQ4p6/jD7iVC0q37Nn
khD9zaqT5o5xp8suKS1PxAshmwQO7Ps+uAejqncEXqi7+NyJiuXZ22XO7qz4
A4ar2MzNhXb5T91zCbBNYKFs030nDXdtQHokMZ1naTmiY/ZfqWIr2zQt7H4L
2F9bKmLJy2lGGtilW1AlCjh3dF7a+kiQILvnxHCbZms+MJwuI+SMpckXLpYD
TJfqaWlA1PI8cqx32bOjBLq7fJyWtTpWSE1ox+fpoWBaTG/m93VSXaB/zhzX
+WFqdV+sBiqE+S7ENamrteVfOEOkj7vkEqNFxag2b3v6SqORFKwFXkzHnk0m
5rKBUHrFlA4MBUQUEI//R+Uku1KskfBSI9k/X8QPZuhtTadxTDii8aTF9Gfx
7QYs8YzARV2a7H184jp43irbjJG9/bMRpg7ki3ISC4nUpaJC1kAhjw0BysaU
5p27oY2bwjDzFVQ+qYCMjAvJWjSEdXY0zPU97lUwzkqYaIrnp6NbZAyPfMbf
IDqWLHJJxIILD3sCQT0iK7AxVMXfIAfHWDjnaq6AxWjOtanU2GOjUXG584Pr
otI16VFm8c6wNL84N7M5XxEWzulmhnoA6vZ+SzeKwwSv3RSZliZBDK3rqq4F
T/foCFO/CSi2WtBVIgmKQlMapCg4uRqvZTYQPTaA/zFV5dAIAgjRk0I1V29p
ru5CAYaErIxax6KYX2ixew4PCIvphJKKdmYw8urkLm7hpLlrW5ycb8ODkxS3
2B3HNITbJzC6xidKvf5aov797U4G21XPllXXnucWzBHq1Tf7L0ZJ+P8pVOXi
2QBuRmuHABGGeRFDB0iQ/HFOEZs6cKtE+Y+2rK5POKWPRWYtEhZqV5GJ6/JX
snNs6dQ68aThEctEK3MKk6MebKDJdAZjvaZGKhrWcJoHU66nYdaWdZ5TTFj5
JWwf+PX6txA0xo8urDBc6gFuDjmN9MWipMqOFjad+0PiZulZHjfRHYetPp9P
UmspfkETxHROd+7+9pCv52zzUnB/jK7LCCsHOc0XbX62Nb4YAT9SJpBSmgrX
kFIlgzsF5UkZz/XSxYi3P4fkTFdhmUj+0vw6hzl1CJpnSXxtEUblq789SKl6
ZNPIDt/cGYRfo1ILOrWJPTrhXCI/1lfxSa2PrVLmvzHogi8t9iPQJlXPDVkX
IiXBdUbPoHPyM8O3yRoQzV/yeDFFTJl1bOcZPzBSXkHLngU6i4No8xIsB0sl
vFfBPNwtQQsWTKXJkwx+gPJe9vHLySZpFjYxFwm0tLC21DXiCIQP8NnuZELb
pKcRn1VgM2P6biKJ7uQizeZgtc6O6WxRl2G21QKlLh2Lo1mv+/Aod7E/b9ZI
GAQQoJ/Xi77zgM1Zwu0drXMywrnPUyCgtYzCwfsCweEJExL6LiJ1H3H6T+jy
TXhTgYRh+fFQgLifZ9dD7bPzMnYT24vUtn35u0h5ftgURmJ8I89WwK/5co+x
IZSGnNcyUwsPeFPF8uNWMmH+mJduCAZKz25YH4f8z+xvmC4T+CILgGtDVh/a
5f1m8egbW3rcYH7VHzGhLhST1w2TY7izhJ7yH7Ci8x9S37RHC0NHL1y0KuiB
2FRpEb1x32fdrgk77xzcl8Ail9f04LuuWNzE09AxEtpmLnhZ1rH+j0wZRca8
J0egyiIMN3PIg0vYwRxnnIISFAf3B4wOb9J+rDAQSZvLPuz+Lctn5JG7fwcH
c9CgqR/9obpxkUvRLomXeeSJycii7k2AHdRIuHLFbiuQqHw7paQvO6ItnHcw
ZGadkhvSk9MnktzHfOO9MbBqIInhYLqpSpgeMsv3iV1tCTNJMvn56gkqL2iS
117U/9T7FGwNO8KLT0df2hdioBtGrSj513uqWnP+IFTSnGLtQUOk4SGyly/m
MZoApWV37AEF4KhSTDB4si7I8M/F2C9IzHj4Sb4FGUr0uCh6uFuQDoqqz5tw
+C1/n/yiy0OWMph1ihtFG0tptFkW1hvtS6qMHgFG4gb8KVx7cVLCwj6v94Q1
uMKwFJ5Dmgj4R8Zr2nK+j7OAwdhOk5aSclLQEAN3d2z75+augYoGScXAARw6
xlCz3+5EPIhb6DCX9YrsFFzvUxyLx9ruNiX1ZzOB6RzZy726YjjtwpSdPsVg
e3Zqc70MZCz+Sd5uWhXVhpM/gxjBxdeb+bMMcJGv5jC/FYatvkeYaDpETEDe
WSEHVXAqFX6P+G+WHWiDuJZH9si2iTvkrmNaaWrdnuA7id5aUTzjKg90FYkG
k1iIiINrHJEBztDvDD+YUPqJhh437kU0pZttAxztav5S/2wAkk7CCk0IVTpp
BMjTyAX41VxwmHmr143g/rhd4nrFxrD11GzUWvaD1IflKZc1NMD1MUTb9jjC
Ja05bgSa6ETbT02EP/BHKcwVedxXFyWkodYIRFHI7LPJdGrqAKDWQ8OghcpB
47+fgA/oKi4rSkqldQMUibmbylqSicEhMQbl2mnWGhVsG39yHSgme3aGo5vp
93NaRroHYQUEwx/Ryq5ucltQclNKQIcOD/mfluWS6v8yGjIdl82W3raPQnqw
G72ivFTG7naB4X6FiYm2snrrA+Aq1dBUJ0zc5BTCo30WpzgLH4I3UxqWrQoh
6+TvKTcaqDqSQXvtF0NPeF/uSXFN2NJQiUmp2jpvSVZSrdxliiRbwV49kEDv
FKOJa2JWMvWAWcr1KGhZmQUGjKbvFf7QbdAvQBJu7onLaN8pca4RDIjD/aio
QP12mxkjP1DRZccxsrCXSdcsgrK4+J4ocG6ltg8FzTle7EazTDQHV+XGOGii
0sujZK+nK/SewQ2tH6/qmZdpcxv7ctCs3ayi1CmFkjOpCpQt9PvzwjVA2DZd
k5BpGw58QJfOnuunFQGK07En/6EPmY9GYLMsaaFHCb/tZ+4klKoGNoVHhnab
3svMVwOkGGHQFtF0pLoJVsdYIZ19EAu7+fBIkFNBJ3BIVuHdVvXwhTudFXkV
77tzmE2Gl/sTsPLV5HD56xvHv0XXWmx2vhID2kUP+wNe7QWsNA/qGnoLMw9i
1YU07vq3jv3e8SLvLbTSgiT2mQwUCBBwFcrTRTUF/g5u/+exPi7/mh0wWQWm
Dwp52nfxgd7XGvy8+FOgAfN5hrYli0znyKOEm68pKQnMwhPFlKRl4khOnXYX
JZGLmxeHvM51ZqmTeB86dx/BJK5kZGj5eGBo0vFX81/8ZGg2JaRyFc/xKUGp
1YZVKV21iLmZHhq28xki39TlNCk2CuYz2vNZssh5BMeD/LDehylprrX9J1lV
DUv6KyzLGBychd/bJ4pqfCW2LG/A34DJO/ImVvKLNBCoutFvAALhHBKm47Qh
Nr6ER/DhhI5Jb2nLFyVoVHvYepHf/aKMUiq/Kgs2yibg+w0hU688cd0tnepq
g8cnQx/UyPzic+24x9ruAQla3mqwXShy4IhlA1kYnvzTExMNHw7NpuHyHhY6
BwVBcDoe6+36gulRAilxsCpTYiLSD61unuWhFL0qRwMlsr2J5FN95IdgEPve
Z/Rskvnw7tXLBIGirBUns9lgolqGOg3gNcHhwO1VoqZq0ZWo1Lbsv1mfmo00
JLlAfuN71zxSY1mRgguQ/jKBcfNZPRq2KngtcCgwtn5q375dVyqnpIpl6ys1
mUJEsyXcGqD+wiyIXP1nKKoYWbcznM5BoP8O+PvOVfzRI2RfxcpEPgGbXpLE
wByEgLwrHLA7KSX2/JcszZVkEFYOoG3k/bFFrwa4ws8xVZYXEMDXJZseTV6S
qED+sNwnaxDNOW45HRL+7DlNrvKD6shaMRUKFSYpjW4dQLObyzvvQpknwNE+
Uz4ZZOIX81HaNvCYBKhSKZhoNZ6B7XzdlV7I2DzVksKBKS6s01fC1IPQ2gyU
hMt7VTILOedsGBzV7Kx0zYVC0lGoerEJYGEe6A2KavuIv8QS5/OVBoFBgDT0
2bF1CN7VVegZLEfN8VWbknxS1uEch5EwvTUaXjVJmUtRGnGKiOXdZM2geoX/
Z6fheLBTR6nZ0XXnZYEIjkQkgeXGL4dDikncHV63n2uI5hSK21Lztp4ZwAMD
ZbkGrDi0dOFpe0gVwIgWtELjvJrehDoAaMIgPyTQ/7g8WQGiMdFixN00kQlh
WmwFYd2b71B8e8NOtoIA5K8wCJZxLrGNnwE/k0pXgKmb6+elnccpzqgxa702
NnSNfguO3dq/XNatK3uRWCUteo5fGbH3BWsO2MsvWr6Xko5KVB2D08ksaYnu
Mf88LxwYKPIdgPL704odOeH/WPgb0pKd5Z8/7JPF+zRsr9I1FCsVVCoRIDW8
yJsGAghtcuGCBF/4/sbV6JqeL3iUGbiGN4laOR23ARnCUCQzF1nOCnwHcWEb
YodhlZFCdPwJK7ell3CsVUEpRU66kCNdAKNQJRYlMpeKMgJDrkwrRWEtfOCh
AR5of6GaP0n28Cm1g9BPsCAdfy8JmCiB3zxO3PiHxzlQcEvTQlw78snrwZJX
12y5BQT6IK1BK1mRfZMTnL+S3VOjRTiVuyQzKsbi8vE3EY/B9bXPfPLkk8Z0
EoUKYqtJHZGXC/m6/D0qO7Eh9rdLqua2qV4nd2GTzznBpDUNkVkiytuVdB6q
ivDkq2Bkx0h83AnUCWHAKJHt6pUHU56YlppDmBzgVigqw+FZp1D5W45jV6rG
RCf9yImPgqWIIjwBA6hOt3D0Xgs3vaAdQKszJs5QfG4zn0+t7+NYWc5pzcjb
O7OJFD5gl3q7ZxbTsi7VyzLhJbvldhypaesoJmaI1sDt103MiH/6h8i52GZG
YunQctQ2ETjHqJ0RQo2/sQbS+FNVCmeM6txFEfz8hFKEQ7Gt1RPzCGSTXxzw
w2UAxYbrAuAwIPLNNb8ofnbpKltKZnEGR32GkfdM3tSTaNDZNoPc7ATqTA9d
Pr0GH5Shso+EQOrp9QYCjd5i01q/7J3c2IEDD0TxRZRKw7KurVCN0Ofgq7Ra
0xNy+XWihD2WLnEjQpfPwNpobRoA2KBSlxoxnCAu/cmyLE2fL7jDqwbJ+qoB
FU3PueSc31aT9TNKg8Dq1Uwp07Ce2mLN679e89NovZ9mIStyvR/jHX7ajUQw
TMTgQO6JTi0DEfJ+dXqVAwomucG/fUP9WZmEMKH5zcuGrZrAxeW1IfcP3Azv
eTRwAd2Sb/SDqvm6D9n9t5L3qg/cNJFuPY3VQBKsENsKd7ylAssvOrR2yYsi
s9Qk3U4qMF23ZlkhDVoaXCwgtY26CMm62HEYfCmSGHQkJ5kWpATV4G3BmlA7
R0lMv86CtyBJKbINTaPTMRGfyNGh0ZBC4MomWa6qHg9l2r44iZKCIvD1Ryny
9KVr6kSSq1M/NmB9Mm8f8uPKZdKu+/Sf6esquq5wmJBgb6r9qNhL13qeAfGD
3ExUvxn/BN9vi/57QgmTzvrEx/3LjNx4vmhuGm6/WrsWRrZN7P4O+T670uM9
BvsvFOARHRDRZTIijQDpxWFfQXkbhi+5tOiwIE3h52+jCWzJ0cq3RhrueMfO
BBBFNMMe162+52ofybOR4SBOGOMqqm1V6UcvfzRoZwgjL5PJU1jXdr0Ephqm
+eWoRP61ibnlTvAHziTAEYbpTp/RYI9l5lmCRQ1h1cSQyG2VL5bX6h57YpHN
dIQr1y7xsb2ucOi0aVlx1nYB2WntPPYB8mXteisoc0P5ktnU0a0SoLgMnmD7
2js9gjNPeG0NXOEMuhnqpD0AW2dlhfsoenikZlTe5DIidAwgvJMDPCrCcOHH
sQ7zjuc2+QtZfLdIWlB6eUxeLv05yCftnwoRrBhRAcxM7jPeUV+w6exQvZgZ
X5hsqrWMIWU/1+79NbypWcdfRorIhElh1jKe5wsk1us45X0SVetFKxfn7pys
Q3G65SKB7b2Z8L6a7I6ri3ia00OTy9nRQyapWVA7ZqdK1V7kiLqvZipnRkmk
XbhoN/sWzWfTyYmnam3b4kQDcPv51S2LJkYuLN5FOSKruKlw842U5iqgWnuu
MvVZPvrUTE1hmlqIx2shZxQcONkodR7TwqdTLmAcqBLtd+JRDS8hdcU2S8Fm
MEw0AOtB6cUZbfzBhKofLxRhhKrq7PBQ5IqBiPWVzUD21druvWCELbN/xpYE
PGnp3ni2+RARQ+SWmzZRE3Mo8b8ws5xKi5r6QvUygPtPTphGYiK9FrUjlW1z
vsRh0eBprGizgTRmtXXSJ+oz6RpSPKZjnCpVFBAMJVXyvcqXYOCUmhu3MHsq
ZaWL/XD8jreyUo6zoufBcBlGztKrrquaFos2tQvaS1FWpocVIoREoTtXFixn
NWzUUDoOfRcKWIkRv0h1ooMrZ9fINFHsQ75aRiFO6rgpStsOV5rHyer6UMtE
BFRa/wvlO3c3yiiWTBep0OzJFizeR1h2M6mzb+neSNsu7H0p03SMfWExEViW
O6Mvx+SyAT/MpggeJVXxHo4QykskPJa+0HZ0qOFsY2qhfXtLyL9gT6fWjMra
zRKhOCkDD2qheYA4uqwOmD2DjoTg3W7GvkE64/ZhCcVNDmYPhUf82JTeH8UG
Z1+WyJz3DlTTdrxL48OqiAxLO36vJMK9YMKfaWyZKrPPOYDQMbo6fBD1X+14
DHskM2ycLC3/0wHvU0uCEbW9LT4zurrJh4rcw/oUOgUhRyRePuw7h0bkbD+O
TOOCpITFlDHm0TOAOz7vKYF/7HiRDW02Q4Q+ZcK/TLs2FaNDnQL909V2BdF+
RnIFDq8AORBohc9W54XH8O3yc5oG6JUeShPxy7sWQkEhj18c4MVxltWSIbyJ
crHMHwTdYUfzK0orCtcjhTU27jC7FwcVgkOWpd9ppFGRGDwQ8pi5neH4EXsC
SdobjTVKN3RTdRLyuj/recqAHHC1eKv8GTl6DEKjZvEeg5mG5xaUcRpBMl2M
9wBR+5dVeOeW0Dxne8rlB4MgwL5BL/PNELCKmy4RGsBtF+jeebtKJDtHx9jv
9gLsmLVh8VZtHEuv49HNYi6nEPh+rtIfjw6dVy6WRqJBnIBauFMihZG8H2hw
Y4gbMQ+5hjO/MsZziOMihPeoR/ZQMaHGyXb5qoZ6k3gLBTemBW6/3iD05Qpf
1kXMT2VfOVYS3m8JiD4CCSWR78J5C1S34dT+POy8bdBD4A47VWbbQztbDwoB
08OCHM2YNDM5VPg1/qMZpak7fiMc195ySj4eHMp8VA1seMbF0dg3NtqUg1u0
nQ+w1KlIHSDwCUNtxrKp8hc55cOUMhBkbEwrBYP/IA940dlUOLhqLkFWMxWD
WVqCS60su+2Xp4Yn3fhNUFSI63bybUvfMRcIcvhaZrPseL7xkMWvomq4UX+r
IHY+l3iGXv7MRA2vyA1P9jFUHoBQg2k1xKZTpvrriBDaj4U+6MmTn7TWtIdb
SoURGgMp+rxTN/uqvGh6vinD/ctejIrPdoFJBn96iPluwzSu1ugUhbI2Fwym
OTUSgJq7uYTWZ2Fs9vIozWLXuZHQmYPSKgqiSZsPVUgkcaShct1QgjnLRrdU
FAGhHfmGkb7tOVFW+V3hrpbHaOdotwP6YISTrHz1dpc4toOF98jY6Y+tTEtg
D98J02NcUkV/REiRwOnhRWTXcW5VcyRNPa8AY0XJO9Fw719BDhlfFwjG72aj
u8rjrcV0JUOwjR3l4tIym9jPGeFb+4ibB0+t64T+2yvZl8sH7HHsDaeGL6dG
kjRGzc2up5XhKzDWlqVYbEgbkcfcIjMlt1kzobMExByWIB6BvKOzCs2I3PYe
cu8o7JY97y1b5Yzzko2H3Cxnye6zdGW5PaIVTicAE0Z3RkO2jvkQDr0FMJLD
v0MBnvZpuQ0Fp3cl/GifScALLIOU0oLz2wuvgXpGjgbP47VTeDCN7h2rHLvN
OqRauaSC/cG4wIvpMUlfXhuG1er7RmTmyFiUyhEFrq+WvT4cFCBx6Ak213hZ
0p5TRkMi0s1hP/UAtaswBqhRGnf7gKWvvpsQkJQ0Y/GFWe2fHAi6NbUqBZ61
dF0P7QqemqFIJgXInF547Ly8II6FVse1GmRc7sKxDqLi4J765V1YtEb8ezsB
aLkr3GbnGTY5o+dcbzGcOKkWpFPunqPJFTXZ7Zt6Eo8hDI1oCqsqTZaG+z69
6aq4AXGR5wvhX02SiP0urwsUlged6Xs2eAre8xtv/YUVS+TyauAphXH96XoG
bf11OF6pVALJj0OQIe5yuR38ij8EGGHBnZrM7cp39OtjASfLOsxqidsshPFf
NMoL6h99Oet1AvgO+xAOV8eRSZxqLmDILqeJPAOBysIlWkTivzyWNZPJOMDA
FsORlcSIOwWDvAXbwpGVGpBPZnaZGtXARYZOcpmTMfHQ2XofkmDk2Br8Lai4
vI1AVeQfJG3ncY5T3BJGKLOOaVsSWcbolP1rGCUv1iESEwrlQf1a8N6PCf43
pSaJg3/0CJAt7V3Ri6wSiGQmHQjePwC0DUY7lHyp1bgcjxO2eruwWy8GwKft
FaxfUw9R27sBMR21UkDbArY8CieNgCcWkuIPQj/zqzNTpDqm1NOLzwBkQgpM
T8xt+lwVtKixxyhkuMafbUknbmypGmqk3Y8dY/SXVh+st6U6aMSpjx+5vNs6
35mVoClN10nDYvXldQ3A9z9OFFEAVQiuA9dg19PZp2XRUKChNBx2mzIHdAzt
GbFFTXC2echLPfcKVAl/oaBaE6dbgZax7cPJH9vs3igcDhAK+J2U80UhRg3H
aTufRfC0JxetncZpOyNL7nJt7CgP1YX9iICgqv2dZ1pDUCunMHjpdBePQQbI
J1JJ7/n5LVDV5zbY0nTzhqaek6qXjwflGBcHaUIwO8tbSyc91CKQbOzVC2vl
6pq3u3vEI7YiJ2p2xU5Jl7oUPmJfJqAilL3Q2UUVoqUuGWF0BqPuE5XH193H
n2uRCOLQ6fJ5oyNUj0h6Y36SmzTEVKK8hDhXSlhW8zPz5TMtDNli2OHBjQLN
KGGb4dikBaOWjXx7tAqF/ApsJ9i1OtwbTM/9B9IkUyddiW1yN4taAm5E1zEX
Y2CTLqWZIRNLlNWG90FiGW1H1PgROwwbHUIUEaThj5Ln+xtF/UBeT9qGwIlR
ddN/GZsHyitlx61+R/NxbmC7dJueme0nfS8z6iSf2BTkLlaWY0Od4uwe3lSV
RmVtPJo1ta8sCHSpoM+8OYU7wrFKvv1S0aJ3nMh6IzUrYmOM9u1orRjK4ej+
qy+VfKCCVv8rqKMehXoyFbyVsDJIJT8+8f1PvvTtYL25ykVEV3Bxocb5MDHB
0nFJiV5MdVYTaZCP7f0AVcEwUi6y3DYMml8Le4EC7XpFvszm15H+x80zI+Cv
NhP11poKTtLxkSlhI0NE/Zj6C07krKTHrd4M0F9llygDCdOKgEPSx8GCOeYw
tzYievb32gO1Akjfmtx0zixFV0CFUn8zNKa1+1LqIVgWwf34r/lCXIMBE4MJ
nshXwALtfZwRujT/nmuRPo7Y5vO6xcnGCk7A7cTLfEZrENSOuyVdQXlg9Aml
yxl5hxwyMPu3kDUeoSvTIW7k5mSPnBEBlmMEFM2R6l51CdBwSjkAp0b2ShCF
+XahwTaBl7omcP2ho+C9ZATN+4K1Tr8BdLnL9Fp6Tyt4LeIn95Ijvo85btF/
y5ns08UnGmFN9JS6J7nsPUQCn2SlRIEFXI7wLkY44DjHis2sfRdUOg+NrctV
9bBQmnZaFV286891DFTGFBOXRcfAk0d/IFRyd3Bsg3EmZecswfhL4IfSNyTs
D6dv6IB/c8PzJDGEazbQxsFXGrp/u5CZSLwQZyMGb7x7HVgPBLj23dA0AcqQ
i9D5ihiXYUuBSHnU5I/Aa28o1Gw2unz8F2AaNy2lEwBz1zmEb0gPIEzQNmLS
f5Tb88It2+EzRsJUiMVVNo4fcn5MkO5j98RfC9q7PvYwgNQO4lxs6MLEUQEb
hOrJB1pEPcymdAYRh7hHIi2iZ+cdhxB4IwH/rtD/aq3ic4wbXbY8UgvP4dYx
ekk8sA1XI7Nx7eyWjjn1wAj+0nNmNEMqv0zFQBLNsPVoK8aLpKRxj/tQl/B/
JCkg9lxmnvneSucAetHJxmZ/e7pGRU4xuWzMYpHBBWibE693syUDmusyWRwe
vOvwFZYygyZV79ARX916L4bvf5/7azQkazwpgafaNKnsG3UEuPZTKi6w6Da/
9B1dNjX6Vug7XlGwlDexv9vo3pjSTM0Klh0LRxaE9rFodQOGxKG5hTvKrGGY
cX2C6lNek3iVPT8JqxFfEQLrMU1v+CzjJAIeYQs0SyAdXYs2TwmbkUjPCSeN
3V+sfLON1aK4XNZ1oA+FXz5u/Yq8wPGsczkXjwLawUi4JaYp8k+cGr3QwF+Q
M2lLtbLTf4rsCt9gWO78f5SS4Qpgdc4PBLKhc5AKAii42/yseu0SpVP0aUKv
CSI1orJzQwHhCLiEKagMqs4kDAMzb7PRDR3R1sGSkk2ylpD8V7oPiI4jIte9
W9u8yrr6kjPUnuRLVUUspa2WsaoRA1biC39OPWHK7KaMNbrlT/xo6F1FE6Ek
5VwVEaz7ERVAdUuO+JlCv9yMAooCIMchSAz7mj+mW8i60ksYusRwXyecy9ll
9vGbK8atAwnGN9Ph0UNHST1q17wrAphgORejPTg1snrtpeBQeZMY2Q/B/8ik
guyNJglobHQGAxCxymTF7M7mPsAg3uAItj05whE86m1qS1bKcQshPjFTaaXE
MmvZSekt9lcdtRQU3iszGeg9M/SkXk10vI3egNMCfBp9/2AK60y0zDDsxn9O
OP/H93QxGXuOMCGz+nx7Bxx2Ow9begGw4XQCt5OtuTdzj6047ZsqgUH+hMLB
wyM4trqaKsz6+c81VpuguvWwrProb63SrOnyTmw/3gP0qjzZc8gz62nNoIyu
zU0Jy7aWHjr6AIoMsrD8jiVKqYjbG4wy9cTv+CNnjct+saazBS3l9UaAyVf/
HSaw6CsY5dRWq7+OOAF9YlkU4ftT+M1OJkRip7DyJqNkoDNhzEy3i8y9rgzO
h6fSjb7ZKXSMOZmSiefKJaXvwdVYBvTvGn/7CKwaQApONq8dBqfv9FN/gOzA
bz3tonY82sVZWigvjWO9DnZyt6E3jjJkoKKcyaL9Fr3cCH8rgmBVCisVKorm
UnjMLtirYBtyctARgq//YslivJW/eCJbQmfTIeqsgbigH9eos1ndYrZbcEXP
zUyDd0J7pEAu9/1IzapAzYxADMKGUIuvUlHYUy/RmwSGxbtcbH3RWrAIEuju
fJvsOPlpzQRtG4Y1X2MBMqIDPlXQWJxWjYNjkwSAEktppy0t3EvP19UekJwn
7PBIDrpj6tvgj5PPpbAQB0lfCmqm2f4v4wZNs/KdfWpCNYusKTjLFmGIfenK
PO+0MlGSCtpJGNpn8fx3NH+HDKk8suIOOucreFPalQMBpdXOZFZOnPuHg/Tl
1MDBszK/PE2NtIkSrEwfe1hfIXvuwHunsoggQne1khdPn72f6qAKHVVQXBtP
kH1pfytHETn9+LjFDiHcShQtDk0AIZ/C4HIrxz/gW9dEmyMz0Hl3Aj4m7huN
H8YCVhvx9qLj/efrpYioY/QtTUuejmP7ja4YIAhfjnnvkubhPx1s6Q6vqpQk
XvKEeTCfRrRbGh2BJGKl/6prCb0Szt0ZTL2u8l5NtWryDsxOFGYgnijUacVW
SN6lQYcMzj8x5c5dfLEOl5DN9wluK9/tkTyQsrztlSNM9bU1Wm0ssDAdiPvc
/86RhN2vr5Uv/DxK9ni0kBN0YsPrROFH77PsHrUl+m1jCGnnSDgkL76MowkN
xrdmP35sAQZaS2XmIEUIGjaoYcXTZ6nhirA/pwqVF/thnb3zfRWPdoVwT9Bo
9Y9+Lc1PjPJWjajkjC+moJNBWXWwR36kc1GLb/WorvYJatdTRkCHQcgoFSU4
SrSjg2ZTV8aY+HtUDLZx2Y3sQoc27WPFot1BzEBJtVJa+jKFwOFd9dyW1Vkx
WuyyJCrBfqyoAI2P1icFsEBIVHqMKWqicqHxSEoI2MyX2pRT1PhBJMvO1OpD
fUN567UQXFkU15SLdl/VhT//1J23vXdNyMlX7uUFut8m2scbB7AoHf9vdHNn
SmDkrM0+dk2kDNwJhNxqyaT2BpBIEaG/PLp+q5rAZ4SR/vhUji2xSeKKPXQJ
EGQht8hyIRPKZ0kHoxPmC9/+XjFlnLMZ3LL8B19swsKv2Mj9NC971BiL8c91
VILU4/HaJiafREiAutiOjzM1IMFYVj0MxHmrWB01OxYwUYnQF8a4BJ2jl46x
3CQLqNVgvIPur9+Pt+3ajTDxJHn9RZtkhVXJ71JwBEM8ouLyuIk8dEtFFMTq
hKpPXQwpaijYbP0STB6jlF7GMOrdh1uGg+6g7l8+RPng/DDv8kpJyLejdnLJ
443aq4Z4jP4MdJ49R9DWe3zHubeJDtmIQAMSMB0hdtygr4CZ/b5ZC76KWcP7
ZE0tIqduEWmkLDNOceg7hOIUaqaDTHNJw7gKolMzTv4cTvyRD9+cc0G7Tb1j
XqZSgdMaBZhYQM2vME7m4VESfUjGcrodWPVPMdP3x8np1Q8RXbPRM0kUUc88
/8Wabx/gF6Lc2+SBxL80nCqFb9GQDqaqxGmMwCjn1MsYgD1W0xrfuic10RqH
eSZu6KqTEs3tUrVGYZd9J66ejK6AnUShK/O5DT4uve6NRZQ9gDbt/ST+LxyT
NpHXw9X4n+Jdhhe+eMjeFTmeEgKJWQVNSV2i3OzGKYqwqYXxfd9c8KC3qSb/
vw5NRWl1qD9h04t9bFJ6+XDNy1sL2R3rwdFGIiNoz9DLziBP/z8S1ZWYbl+v
CR0Hl8553CsgY7b4+HdHC2KBmNhkDmGJSvAECH6gV9YbBewyTKd3CacFsjZn
AoAmC5YcVUisuyBZsqn0+W64/Da00Npk4KdKtOxmcrnQhUFHjLF46rweDGcC
P3jETMMe2Zdj/+8QA/j1VC8TqloAsQqdkNyNF/tOtnGhCFYmN3UJuCXWFXfT
5HuDl5Eu4IgN/+O3Js5tK89vIMD36uC6wVUEk4xUbqG/M98rLxEiTMxcJ6wm
m1rhwvy2qt6hOY7pbiLrpEjR27lHKe1n1uHMv5BNH9wiD/x9MeI+3HkW4xsp
MC1q3NOY4y/DKrTlk0x36Idep7qbSXsyD0y8bJBqKte5HBUdUwsj6hd5uNSu
tjOcXrqnsnfTtgemVWTv/RZbIMdYuRnUGwGZUdZLtEhovnY2V+0Ul9wq5KoN
dxSLQ+6xCFggYrk5ltisvd7SSCJU4oBNOUOjlAuVz+aRy/UUqpq/sR17uFY3
9ZEZ26K7COxusKQfVQ7zTPLaH9FDjGWNL3cssWwOW+jjK9lRu6gWVQVqoE3K
NHxXrjil9o/oTDvZ3G31PR9psDQYpGPajEmET5igcK/FcuzLAcVsyQgASiao
oSsAl5pqSlYxIgP4x8jSgv1WMWwCQoO5hBTtSrF+wyJJNMeuA01n8KvUCCPw
JmdZ+cmNlIyXUR90hyyF5YNJ9xFVUsykncoi+4P3Ev85J35GTxdcgnLIOYaY
nsZ6Pw2hUTBLK32l/e5rgw83gPBp85aL0jVEL9TPgdOk14QMw9jpOD8adqZV
zivEIg1RL3+8kVvB4tNvBHlHukMvY7idiTc6TN0otp1jfmrjy5lfA421o3bm
0x8gZwEnq6KynQlcuY1iO1amK47Oezba9Ls3DSBbJzePxYlkXYebetb20rAA
mGgCIRVmlV6KOiWofXKEf5c1HdQRPuCChhqUIBkNFT989yjxWMYJlsfSFs5G
RiMjzcIqUduVatJXlHhrQWTFjZV390mU8Yakun1KTlMff8BYW/ueISAaB/Dj
sSAYeQD5TaPA3sit6sQJGgxOTcxz5x+R9cjnPivehjg0RfOtggGPmpkVZRyc
OMlyP4ZDNErHXT+aAKcnJBY6OtpXbkJsYlh9OT1gZ1O3nImqHZRZ8I+zDb6H
Vft3UyyVXaWUNRBES541gzv6BerI2pbpwUIQmPx5FJdwAl6OqeZ0oMiMffoo
iwFlEnbwlpDX2BahUAQyCJ3hqCGLfJtMCC4ooou/2b+DUvpqVsbYmtBG+kF2
M+RYnxmh48jGGME+6Is7tTPxZbpzE90OHvJYLj0OBCe25o8F1P5+QQ75fX5r
0pLmuJ2c0a3QwTSVmbT3/W1KwMqJXFLZ+8l1K8+6ycHv44OAnvZJJTE7uDwn
w6xgIUwwZSxZiyVF5pFbqwTywFqgya9o2BoGks4MW462xNbXguQ27XJWTyIB
yuCWVhzWr0rw9Nm7LL7f+CCam/JdbwkBHXltJa9l6pBo6WPm/vq4Y6MRwNPO
tHZKaZk5K+I6SXdLkM3Yl1tJBENH8G+u3bc0A2UWmkTGLdxRUHccWr9urnS6
RhH4Or9IYGAYRfaP+Knb0kfeOUilg+npoRFNt4iHH36kFLb3M+LN9uZaqKs+
8JXmhJRr+424hbHgd4zLA1JIK77h1ccQeDHaNv6PwziJylCqOq8x7RYCj5Nr
OkebpV8fVqNKxmhLPo40ih73mvUGSrC58/YvA1jK8/KSsfBhrij052scw2GT
k2j0at1jgGxHH00nPFV+3ag9bc9xElm6HyX2nDlHwy5shOqdMphA8E6e26Md
dJK8q6ekMrj1RI6bJ6NHOgktdlCpaEIMNlFA/cHhVNCWG7X1JSseNaRkawBH
9242AIOsr6al5DN9yzSg4kHU5obIat1PygLrXN7nWoWAdJHGLAMDQlKAXtVV
TRQ1/P8x9QaKlCrbgHrmRGBbLel+6avVrpuw1A9lR4GKozV5UHr2hcPb6lKM
M0WXXQlNLj1EAJ6aN/tw3qb/fPWDCNXVpZu96sfO1968kL9ZBupwkWJC5tTZ
4Lv68fC4d9LEL37fqQC7hKOMT5G2eY2l2NDRDKeTHWRZknubf7k212QcaJqa
ANO2qGlByjMVLS2+cFSXbfjnzxou2mddkGSb9lI2qhFG7az3pSqcJ4wJfg63
VjEysQebCLTaBZao8I4nmjU/pwh/Su0Xdlpajec2cDnLZCZKBLCEZC4BtDgE
213hfa/GgfsrFXG3k1vFfxyIZRsWsFQgimJ6SrQar13N1VYly5oabT7sf6jz
gyozgQwCQ5lvTJx8DnB8yexPyByRcZh+1L0mlg3Gu5kFMr5YxtBJumhr+KvG
22zt/l/lHVvtPXN67aa//EMQbdpqaEg4Cn2jVpW9hz8ZSKdnL4wfdfBI6zE8
G2HoD7R/D47qAV07k8zG0E4epGhLYqGk5cTnkNWzaWb9nHBx+UilUpEQ3dKP
RJPT5uQJTejLPGixYSvVNT536WvV/JJHm9xD5uyTa/jYHtSkC7KkVPHXuG2m
u0kThKUhbVTziEDQO0uToPEZZ29pnQv9cm0oTYQfqiJ5jIw4dZq837mRNLVQ
lZU3BxIgKi95saohiLHC1q7HIhotbDLxsH9vFPSi5w0H1ndT1bQEmX13NBnZ
eEGXz8+kd+/201e/x+iIBNC6yb76IA12wSkqok3CjRr8vSdgWju/ChCNEhhT
EFSQ5BPwchwFk+Tu/wtle2UgkH2qBcvqDgnChq1laUvm2D7lJtebIQoVgDA9
oexgwWTqp/8ok3hbSVnyjTMvUD6QX5R1dNOqw+YpnrG9ZQ6a/hkK7+wG8Tgs
5dnHT1khi1BohOr0U8ibIu5EGOS49rYJ3woHYd469qozFykshHedPw5FZfP3
4ukBEteWW4LYHd8NdWQoh7egaKpp9ukXLMzm2kqR6drJrkk4LceVkFiWekCM
EI7v6m8ioxNADN6rtQ7JQ56z8uecrsZ8nFw6uJ9QM27Nzpg4s8P36k2AsE79
dtUXMaaQRfaWYf3KEuIHtFAzHiS2WOtvr/Aha0kktmvXW2Ketb7r+i3RbetF
kiCS10uhSf5BrABq4327QkTu18uRCmhpkoMCeJhY5V+5FZImfVb5x3ySdGEg
LKVDDbsKJ3LgqwkxU6pbR1x4s18LNHFMh42EXH4B2oGQ4590Em6DmUVeqmqp
TS1lZ2rnBtX4/oWv6sv9yJrik1YVqgq3oE+W4Hn3kCjRpYtiBD2B8AlQzzCO
IP1/c/2l4eSOrGxTzy9JLAmae05bEFaDy6kDEQ16ETznx3cWCwT833FPAy1L
GlrAglhPZ6FS2phsDAd601s9D0TpDVVPWlWtJ4UrYAZ/wwjLle/4QQ/lBcAc
eHtxaj49si1FwLuqGRs1w2eLdHjZZtw0a7sIFfxYOyQSoCF1o/yFmt81SSYK
aj6hkStdQ8NJon+NcvKjELmS10x2UkhOeocMLxk9Qr4plUh0M/oHPnCiJd75
xQSTHPQ9Wng7lwuCJ0FdcPM7VJqf7t56u+tBz2RTSDQ2FvSQcIl10IuNALRq
ypv1/09sjdTkCr17LWdX5gzBnuODndKzGhmFULMZI506WJlO7LejhaNuGHcY
0Xm2AXhaGkuiOgXZf9pbGlCxUO7THWdr0LRft1xZdWf9fLrID1EDPMQmMLlg
hXcCQenLQaatds4OSzLx0/vxtJsATf8QMU1SasKm8RogBVk7lMlKmoCW7+/s
EnvVCyqIL96g9Mgxzf0Yo+PgFJ+x+cf1Q8IT0mtWYV4Kgw91qYSDWwlRt9Rr
pBOvoz+z4APxBdfwuZe8a5YHyO9J10kJQIAg1W7BAeIr64ikrelrK9ymbsvF
IduOEQYuRWbgp47N/HmL/eWD/jJAwjQUWKjyvH01eRxYTZIzcmFfEOgxe8V6
dzcvDMQoxeBBADNKIKcUY76Vq8Eb0TZsf287d2pkRw0SmggirfGKmt0KMkW4
7wSAarNxJHO48OaFdpUJaZGl7/OORgHgvMek5VJinLo/ek8dqHDzavNykpjA
P9XOv6xfUwvlg/I9VL1jTeY9ICo9mbT3yVW/1u+FtzCOCLah+newJx7TE4zi
i2cXajR/1sXillAewa59/SWh0c153d/PJ8EmANdZ1H0rqhsoXVTwt66GA8I6
hHYmJg+7Ymrrs8ePCqFAitmffnVvBv+q/RGZpnJ45FPwEyOUXOHSkQKNSFH9
RS5x+Nf5o8CN7Q+a8ZdTQ6nqVZwQeb4E7rKEtycfFwTfa8nUKMlNwlKorT1v
ydGggktqG9TDrMjSvNfCR7s48mbnp891Lccvxuc0ALPAbavy48a7XiLpJfSd
Ugc9FtEXl+WtLYfwPlXCmXznJXqJy8QRSXoQ+hl1aXrf3P4SCFLo8U1mTEsB
z+ldmfay0z49m7gB8d0tWgz8Cw04eBl2rL3WzAEw8DfHXQe0SKsLEf5/rN2c
JqrAjQDZO6m1BRVFL+aq42kgaUy1Kj7A09pc4B/lnO/q1zV/L9sNKxnPk22U
dUyJcgbE8pu0GSXr7iV2hX8RI7if4KnTnEDm0zMKyB/thKMH9Xl5B17OkUci
Mma1XqJ3QPp4o0RSLsBs1NLb81fwcVxk12MCChWtEAD4lgurTeo7kljGntZK
typdbeu6c+eZGEASqcsFzThnu60wWoJzUBXb4vGPQSGfIvhBqDM6ngIx/9Fs
JkiF9dRabqHN8Y0AckNi1XKGytIczRyA/mpTnPMCDuEbYjgR6fAP+oB7p2YC
RieAkHVrh5YHY3624L3+FCD/mDBVlhCovFXtxMLmtOykK2Lu0dBzwpNHS97E
aOGhyh0fY6Od8NI8et6Qz5nVeDMyyg8ZWzcyAYl4atJvdkaxtVfAvH2dpKtl
JDwL+LPPGZAXhuGZWHUQmU63YTNsnCTbyUGAfFVG1Bom6K48U1NUnnb57p5K
+C5qyr0K1yrEKy+OWKnYd/A58YUFEXcAJHjaYOETHZivzQNKXoIXEjz2rIjP
rcGfbA5dk8lfc1Z9YM44NGWsRkGbT+aKVjPyvGelKMmlHq1rmVMMDMwHFxJB
mlpgcMKwnIOTk/jg2QMoPqfwNX/NiJ1Xkg/7NsvPvIcrQAk0dVlPaNAjy82O
MEl1In4jZibz24lsWXpADwvKs0wMdalSSfpViAEhKtbY6G2vFXjAO4+HHCmB
mJ7/ozj04R/ppkXu+p+9OYd3/uHWWXEogadeyzqg7sb4ohEinWolYW8t7IyU
xbMvcqI60A4XaIlasd3/KIX13zk1hoxUIMx4e/wWIkXKRqXlfzy48s1DHb2K
1Pwr/b0cIXcWc4qVF4Tsdnvzf4RcNBlKkdfW7gqgEWxb+8BtxFEwA5pUoMSo
z75zO5Fr+bSpqcQErWlZwlOeGizWUc6Lj0SCltQbEZ5vRh3+w9jtto4fFPse
nM/tG6UQINXRnixXuIGZonjv2YQBEHepXUTT/dW/XLX0Y6QnBdULNG3r6dUZ
tofz0LqvG3NGUOfNj5q//7ztbQA00/Dgtf/6HLy8SxQ8VVVIr88ya+oaf0XL
Mg8tCS3XFJZlpjmVy43YlKZFYllFNfc+NoopiDVaZgx5ZLgWV6JYKoYHGfhm
a/nBuEiQwN9JlnaWgNdFzaK/SkG+TM/OQ5DG6laef49EUt69PcWqqJUjiFXa
BlFS5AeUSQNzm4INE14CSkPhoflT4vS9ViTL5PAjRQwL5lLKs1/6LiQ5hjRD
KRz54Uj9MVv4FrOHMtY+hajS+DKqNd3jo+Lf5WWThQGeR0tLgVkjYGC5j383
sgNHijvorktl3o1YfMFNrxtCA2aScfnr+o+meR/n6N5L34l0Spqv5ROXKjhL
JFADDh57PHPx0SmCPK0IrCij1DeuFkBBtwOynfUiZUhOPpyKT8RNnEjMYu9c
ONMdlWfiI78/YraYDdvLH6dYchKoFKH5uMC5zsMo1ZHUPYuaqh21EVc3aCbd
7yi9iWujoLSO4Z7ujNBfl7vJQ+ssWfbSOXYbwAoE/XfinAM96eq0vsSWAjR1
2P77rxlLCGHAXRnfO3lhbYEfW1Vo59jYOeqFJug3yIT9rYQUKWF+QUHUWask
EcVzXCpWwkSKBI439NnqrlQsucnJzMfVNPHPU7RP4zwP2N+PZIco8ANr8+8y
VyfwgsUPTjPsY2RINKw/8nUYa5wjUs6Xwu/icDtJB2mo6UBsqVBCQpqowvj6
vri6/nyuzTqTfURp6J+NuynwcWUUhp2CamgKFODtA6anwQFeo3FLXz29kDPa
mRS/Yzld1kbUsnQzgL4kkm89VybQfosGrqRjzZIS79Ku3qJCvhKurkGdK+Gw
ydf7mGdZRfRWxoyZ3ll2dgmefB7zxSyrwfmHpDQFO60VfB6LMYa4Dj5w4l7N
k2dXz+HCrYDmoLyAfssbhBgzB2JWaPchcQhpBFAS/Pzf1EvQ7RGRSXRsSO6t
HDyFvyydQOoa19gjvB7sVSbw79GauCKLKFrpBGwRnvG5dPvuSh+Emc6a9pKu
wj6OYxDdom1Lsh6GzdDr4QlgLY46Pp2919psRkpAR4Z1tmF8untICn+Mw450
LA61tt9/+ieAeO5sI3f4pkG6hHWoGxcpJ+/m2nPF4dQjxAxhHhUHhup6Jopg
P9Ktzy+CWuCSBUi4YGH+WA6XevALFB1ozDeu8V+KMdFl9SrvyY2gRcCf/+wu
0j1QMS6oUKbKtfKAmy83PUBhZY42wREkryPTpV1JISP807d934Hm9Ll/byFr
q9ffIlygaKBTb5hlk75EzRgFW4QoasnLvXwBLVdBf1l0oJrNFbTyAZfP5QZh
8FIMhgqzeSmSy5YIzTWOs8nBfaEhGqvvJejGUwmTeKUKF7kieEQFW23EXVMT
ClyT5bGC0j9RwQ6Nj+6ETV3rm/wFG6i2N8TTTyIXE8jK9MpmTti5RGzcCCdg
JLRB6QqYZyJ3zi6MSRXvR2MwkxfI9UvV3POqOC5/PxCPxN3i5XWvjyozvpJ8
LrP5SkbcL/6ZkDTKfLS1qTJFkLJxdFM+GdZgp3rXUS6kqlRzZJKb0Gse/64V
cH4n3VvpxWpjNtViGRSvCSl/BsdvHMyGzfr5LD8DpfLbteVI7EE9/mwyIXdd
b+VtByV5iZEKpn2Xs1p3duQsaiB0YWAUQ5GIq4fnEV2XeCvIc60aU5QvDbPY
EpVF8LXe7+DEZztlhFX4Kcs449OgSBnVaw1THbw2aQf7B6vk9E2SiLpDVHMn
l8bnO9DdO94mqlqq2COogpo+Kk3B1BfUapy/17/cvpuSGjb3StPN0cUSSZlV
6jedQgmxPvowpu2IUuLGxvO4YOCoKQcfRz7pqhKCtXHQwifNkaZ34fD6hWZG
cSfGOqfRVV/CN37B9URhORU6qrTXz29QzN6cJ+3Nn1f8G3lKPUxyEtp1umJ+
dIH0pLVLfChfB1NnHnGcPeoR5mZ5pyTngbmz2xruIdGuVmHNJ8UZoMJJE5D+
6fx4E2HvzP2f0HcfchRrBKrkE1cB3jW5sB2j2/ZBzC2IMaWodKRk5lBbbMIH
hJ45IsM6I9BtF79BMW/qVyknVyRwIJwFx8XvW2LzQzH2BWitM0+Cf8EgyejG
09noLOeTh8s/BrdAp4QYBfODMHUpsgvU+xOK/zj/iTnLIfqg2Ayz1xbyMRAr
tD6Tc7FTOJFeXKunDtEmSVb11vV9fAytGrnqWlDHFDR0Vui2jgpuforeMRAw
tbPPUjywcUghUqLhvr0Y6E7sLrKK0xo+i9lGHvUb6oQAhFJ7NFCtmuTyLSMD
rkQ7cgWn8Nx5Pv0mle0AiYYLo2kdpn9hqlUjG5Fd6sGPLd4F2NGcj96tnTqk
rTJXgvKkSJ3VL4qACjxDPpOjn00+0sCsLFDfRmCuu8qxfL37/gUdWs57zhAP
pZdg2AjcA5ZClpDfM6IYHpXn9iJnPmk+cd8UlEnDhULmsbIMxZxcOyRakvDn
lz+XNPfjqvut0OkauObhKYHs5Qx0Xx1T9yGy9qurUsbWshKjVIXdMjwt+mnO
rHrVf+ygufFf3LT4TPMc0mH2nQXKrUGjrZ0EfDt70B+hr0eoYoRbWlsDtqWR
JaQaHWIWzvbUF++GvUHxZvN+fMdG+Ry+A4kKqMBWWCmeKZr4ar7PULiJ8XrN
cXOGVjvbruegNKvNJmlj9XEp89ozQ0KPqi+RypVb26giJ+ju8w3NUHQ9CLDd
FDUXK4aEY88/jhqvsJzxVpBG4Avakzp+HzrrJ01px6NW/OZsebhESJ0I7mQ9
VYo5KIrODYl7VzvJyzhZg6jJ9+H2QzFCGYC6qHbACvKJdc8wIDc+HGrkH/nn
6SJcrs8QzQG3EyXxZx0dbWQC2h7R1IV2EDGXVdBIwZqnaH3WUY/DKDI1lMUp
OUVEVVSoA2Ga6yOkNVYNqN2GRP+J62vQFapn9BtLSMKqAVveR95LHjeflsQy
ad6SUe8h3SO95DCNALcPo7xLrbPezE1PNDRriabj0Y8vxhllV8ucH7vVZ1jR
DGRJPZaBP/NQYYs3ST3OjC5UOWzAfVCuKfCl4lvYs/N5q2nCm25Hk5iVZtP3
n5Et8+aiTWyNgIvDP/6J71++ENwTmx3rxibN+1m2h+vYaPDXfsJcUyDLSIyv
cjIdhoWT6B2YqKQUJYVYd7Y9dWz2O+EgzlPg31+grlMlWkWpyTIoTfuYMbcQ
M8Sc6wpcwvCR0YT9Y1eY6BBdVWOAQSv1M5wy7Qg1kkLZgtX03KtHNt4dLrtS
HuGv/17AVbjLmxl7LyY7HhG/NSZG22FWZ/R1S8d+A7xu3DU77ZAOOYF/TZBU
DPBqpDxXCjvNH4PzffVgIpqEVyAqjZjgTMcLh+G95fORF2uSOXvswgFE5kdP
IsZwMAdcBhBDlN2uCWtl7anW8WYVWdkd/Wfj97HcqMp3Cn/zgmZ5s4WTjLLE
ffD9hwiob0wsK0F/ll1HRfPhkqH3z3VhpSDidusKFNvmSgfq24js6qviWtpV
YwZ7YaNvsyh09853Jq6kdaTNOTrszegXr72rbjqq7rO8LTtSHhjIzmZIuc+x
tfSk26pIETJ5AfQciZvipIpjMDP5DAYo2vg7rcOeP+meSR02Vd1RRKBzgJOn
NM+ycRzPwYNnW9UDcu2MR9wIed1aoiSKHYayNOM2ihhE9J5kIDQAUEmh/T/y
sWGsKfHiDHY7ulTHLGzpLhdsU+WIooB/Ic8Fvg83eK9WX2acDwjZN1jUHJIo
x/JmhxBc/TxIyAW50YvI2GTeqzoVKSmQ7fe5zqijyp8GzvM7sOl+cs2wfESL
oJfNsvGbN+oLM0ElJ5WHvLL5PD08dTglPP+ptv22dAMu+DluwvXaGdM+/lRs
jq2m1gZwoayrqFQE/fM1RumjZOAvzKVt1kaF8Oao9xlcf94y/QYhkGx8yZob
eJcgdBL9F1xPGbKsE3PmIo9WYfTxSDzRKVnS+fz0qAxzq+axKqejYU4SyHDr
9QzddJxvN1oSO/na99LX4T6iAe/PEeA9v7XRiYPlyhZB2qTu5r20UsVdZS18
VzOb0xHG+DTs/eJVD+BcMcFiFlVK5lUAG2Zwygq0ijrOwTgUcOGK955wJqct
0l0LgxeiQUjyp+0UL+YgRAONEbhMjGwhkpIsy5otgnEhFuuXmEyGJSU7iQzz
XSnyveJmhTDV3UbxcULod3McI6tkxYKa1WFxsEdOgsXtp2sVWpdOwhg52iF6
BQsd8xe+i86rMXFFmReH/nwvjFTyCYP+mLPMGCP3HWHpC0QMSLA6ZKCAszTQ
hSHIoCall/WkJ24MQ9Epx5t3wTsneoDd7EC3fYR7IckEzey8TJr6i5obKUYv
2eC4kv3W15unuHh+NtAxwJsqzF6jOuOnY9W+fyl7cPA0Q5efHElpYyA3jqo9
HNqYcFe/MuXlpZJPMMURSbNYwzAS5yPdcz1RkWlwcX4dIVTXem9H3M9otmGa
o3fs6CxlDPWvxqdHsvrG1vvpfoMr3K8uuZX2UWON7VWIdnn0oRsr32t7nmca
MJfKR1Qtm/YjuzmtTn+FW19jyUtOhr5JZeEYC0SeZ4kjqmjXPEGlBSnuWt/C
STkB7lG8z9u6xo5Rxh+e4dtJy723bGvO5inWoY2FtEmGrbk+8n9mm9SR5CkJ
w/xS9wkXqYbvvEPolwnG35JflMKNLONJRR9nI8GQFk4reyw2Esa4ga4scR8j
vB3rlBlDy0XKr1hcqahk/Yq4lRyqZ9rn4t9h4BiuMvI0MUSL+LA+Q1NF9/T9
A5Pt6D2lzxQgWcur7aPkq5fdODZD1ymfwnNEUz2+ta4i7uaJpGc5aAGkqk8F
Mk6joYeEkPybCp2aonAgbfHSurGD3D3rir2V3qgvk5D4S0Rv77nKR37nz+Sy
BPCVL6R0ewamKQoPEC0pMWVT2A26bybhXnbP6LSS7nlNHaZeCcqs/suG2NXo
1+zSr5Cw96vEuWr9VI3HgyG7P0UoQFcC2Z/RBt0nr75GisYSgbpii/Zh3/qf
MdqLJ5+9L0lJP1GpjLMmdSDnTmaXvGPWsvRn340ZSOhmuDuUIkEGQcbeRNfF
k9sCnwqhmu1ZICQTcwqnNOXbncmIvDSjk8TK42nYNBsFRXsGJCqtZpg2qnL7
fka+RrLYewakF5epDmefFjfx2crzmpIxgrvliR5quSDxgTDQ25Dnh93h+3fI
HmJk929dOSs1ickLBJkqZDia0V79n92WVMwEjjOM3G9aSYbiMhnm+golR/zA
gHBsm14qpyYLXNfNGzCvOdmzLS7wpPlWCTV3n5FbRTyDGz4RJIDfPQ7+80IF
GCp6NFIb1pO/CpEoRabTsfNWD9AzZYFi/K1WnldzKoCY59JKpRMgLDyQqQPg
+zqhUQ/vAYE+Ldacl3lwl7RtN5DtqXEi23NRBUQwqVfB//p3EfkUzxZpZa9b
jsx4UEclR3K4BkrsBy3tXTnp8Ivg4yaneuaFgAKOWQ9NSZETrOiiTqX744CP
WlJJ60oSm5EyU/3TyLLXso5vWNO1cdZsmkQ+cO2t9D+m08k39/J1UjUNeeCr
KmpQJQtFiL7x4XoL4D4qBLrypAZAp8nK9ftVNIkXyGmXjOr5U4Z/1t3cBlZX
WOAFDc8aHF2Osi1rQVPZlWeaUzCPURmHf78TU8J71Y0jE+gd/5AV7wKmVkJj
y06LPapSdavHeI/bgJMGdkIosACLc8lI9txHAeB96wF/antvmqwEcmir1mF7
Qznd5hzLVT2On7qtx6RVBNxjkoAAlKMkVTkul3CnzTZ9egxhWcOCgh0jO1WI
7LuPB7pPLi9M8JrYpioYtD9tGIlIZ/OGjv6kgKe3cBy29BzMdC3yAFbdF+rP
FiZeXDzWCwVbL2dtTdjtvmtpTT4+f3YxCYw1xaj2aZSGz6nZteISFy+CJRg7
a+ZBNtxhFv2TeMZWE8OLDMJ4g/HyiGEgmV8QTzmlorydvnJAYyOXhZMKCSgw
937dCDWzIGEPwI6VI0XFQaJ2G+GozRPYGR6Nz79GV34UP/Y2nVWh5sEI8DlZ
9Wtdpg9xOsBfIhEzYp9mgKuXzqRgNTvj+VxLVfHSxZlzmEG4F8YJ8GLfub2V
SCRDbAGmCrw77SprvLU+LP3VPCu8BLCqf1liiDTHY6vxjDzEDPOnAEHwPr+U
aETwdxjDG4orz3qKnBiGSSKtniiOuC4/qQxeHb/2JvWI4/QUy5rhB99O8zdk
4V0z4jt6j00n9kqFpprKodh+yIMMY/zBOxr0a8434vHW5dVXbstO6Akwlb4P
GEleZAolkrMYtHCSiO8FZ9Y3xmkp+BlKMKEbpJJaA1aVJDDvx8/5it0QrVfy
CDtO/H6joaqhoIZRwTDfPEXYhlv93grl8M029T54OIYJNzVK5VSHvUHIj+Y5
VNN3qZqSrBjjD7zqQFIPdL5iwDwvw1GzBp3Krr1XDXokPXVLk05ifOMDU0i5
XtifvmGJP8YXfeNroXI+fhc4ISzcGzEK/CF1GFQWyivO6Lz1L2Nd0o7RzP1u
NDhphHBIXDPoXBaEcmPArkdNZwquNLN48g3Gi6wiUnhHHf1vQ8LpZu11zCn/
U/+jbIBeF4w6jncOAZ1fFzvHUAxY31kOap5BrVqYRKCYhgLqKoD99wfAQM0t
KG0F8a3nnuwNzxZ/ioSraCJGQvNkE28JctaQF+KBDtimfKNQrxlab48W6HQI
RT12qSn1eZqls66241pIgGkn6F6dO4zT0/6OUSmlQOxgAkaXutK7lPWXFjA8
w9m761QzauneYKy/xFseIqWkb3xzSxtIISARRhWVNdWraqdsOpyvR+ai/Twr
M9Q778yewOwE+ZBl/9KDnHwZ20FBm2hVUeg36hqtlaLF9LD9v5YQ9E1MKrDO
+e+Ml/lNrkU1tZniY+tPoVBwBkCHpcBVe2lLMdtZBfYxsHFIqKOIMmtEHvx1
YZFyuwoKttkSAEX5ybIOPD1gj84lQLseJoTjZrITZZp5LY1j3ioJD8KfRCQj
rnymVgOjKa4sdLbBBHAFOEC5+luR2sv21uBxhUKUBnPdY319fOra5usDHpap
WFAFgx+l21FqheCjVZ27+2MkPDU6PipMLyfywkPbrf2MFVNp9w0idaPshqh+
bbUFt6FNnVD81eFg1VroAqc6cDZ0imaq7z4/EtZB4WzdkIhAm7CLhPlS6yYL
ZBTeHRbCF0G4cfKkvLA+mEHYyJ6FAx0FAiLqml1nNQ4H4L4Supq7pd3aKFs5
Jse7ImT16KbJU3IDyk2wDZQITxa+UzeKkIXNU9RJ/l9uoCJHXsHM7ifxc27C
hyDYNM20aQd3FdnI6hIGxwSrPzEICR3CceMEb69ALNUCox/gAA0CYNLrDhm6
Gy3K/FW3p92ko/+xX9hf1RmwrTCCIiXPAnzKTQifu1voOOj4y69T0mJveuTo
GN3dxy7U9Ehi66pX1CUXznJMhu0Cbi79wtj7xyosW1rrnHUIzuIi9AHUb7+A
G1l9kHAujovp9Z9mNSXkpBTS7SXFuDIztlKyZDMtNpupPDvknT8ipBF025M2
Jg60/yAfGJ8GTocL2wNC9r/l+GoRvyO7hcevSlpsjDrGMON2esc4cpYjrICm
Ns9mwlfnAMyapQobY7ZFo5E31haqhdrOGbowHYHwaSkIG7YtDwY3U00QzH0P
T8ybtZ31s7lC0BfFMjZAe0PwW9NEHYwUuhHPOhncKtuKHJtDyCbgndWprzfz
ZTIFKLViAjSE8KWNkCawT4h+o9hrzejzBc/JoHky8EALJWZjL/5mynb9Vs9R
ihMOGrX1jh+r+6f7vqZDC6kTZgYmbHdM18MCbiU0I1ij+Zr6NyY+0Vkz6sfK
d0uKu7cTDn0+HZWM79wGP/dlxUNR5RNcifE6hIS42dzzXI1oaF4i7VELaWLc
F9aSBRt0jBau6TM7VIhu7Ez3Bbr/bv0dKpNQlOEjsuSYOGwMujytz9JU+fRA
tD+t8VqhuA8LIYM+lONo5uqFbe5aRtVO8nNMglRX2AOkvBsITgmtfI1/VK4k
d4NW9ufi+JUBm2Ht4ZDfEe6yfc+J73U8Ukv/P5/WQZKGYo7KBBHClJJyBEUJ
Y765+RszUIxdBTKZA4PFJUft7TjgQQrvrh6YrEDujJmzTx6U9/D0PK9Fedbx
+pVL8QsReyWxM+rFblxbjVC5Q2dklrcBPX0eBN2cOJ2wVmgme2zrr1bymKlS
4hHH7d5kmMLHzmw8NuapbnzO5I0t9GWbZKgKbc3tp5NfKjrajrWZxlXh0wu+
VU1lOkMTCkSsdUO/LF+3mXtkNNmNg3lgkOnR4EIOFAzDOuXzcH7pUkGcYVEE
JZ1QTwQ+cx/4mgbTAb7P9q64bUAEKYBZ7+zxzUg8KY+UR0+Vc0efLK/Xjxg7
9oOJtnPUG3Mqvfx4EZ6KaUi5bvQbOJSvXUg2ljd42P0rSJ/r1pKKw5nM82La
qI1vIaftGNuron0tNDTcZPQVwvbnr4KJmQyACySuFaL+xow/EXFPzhHkqTfP
6aMhkpsZMe4Lp+jOdULbx0rgXhIHuSS5DGJ7mqclSo5wxtALqgtp1bLsmidv
0T0eFj/CxdeV5H5bHVRJJsV00daxg9kDOY4BBG6DvS+VehZEGsfKLEzVrsV8
sgVIYH/Uv6y2aUUNMx80n1SonXBUCUYbOHwyx2XuBbSPl5Um20s/nQFWVoXl
rV2L7ar8m1OARqyg9hssFZ7ISErm61imbUTxsDUHBx2gOJTQsPkxOh8CxQvw
741291Qn2cRHCcy+Xbp3auhFYKqngUAtqF++DDR9UqulCooGy1BDfVRavAE7
E584mNdDzvL8GGUz3n2MubQm/4uiyOW+0YbS8QUWmrVTgI5N+vIMZSICOya2
wHJaK+xFZADBcOBrs3cUykJbv1kkGEnSB+plYlgzwEycmEYEoBdMDllqsnpZ
weNyLFSzYrT2Tr51mo2wztbHuL6SV5lhnVeFOlppaWVlHqLrDcFi85+1Ax3Q
jitlB/vD07C1X/aGmm+D/aDNyasWsEwBNZUOp730GFTnhhryooQebPIXeril
EAyiraaT5WZrppF6+7S4NbxdmqCuStBkYGIFTBepWzfPR1VHx8sRlGgKe6TG
/bJLZy1TsoAWhk1EfxQf/8S6KrJ4dHIKcjZ8dvHTeh/eWHQrHFu/CxbBYzIm
YHAoJzJfAccqFtcHMbCAGQl3PTmSQ1ajR5ekJStmz1fjgcLOVyHp8xAovoOR
HTAnpfQVyFy2mQUtkXmG6fXhQNDr9CjdE5RB9Tr03ctRf2TTuIR9uihyxhbS
MgjqeNVWwcanluj6jWva8VaCcd3bLwFGLGYAuYPPrREe3vNqNlHMiUUzIy4L
s2P8On1KixzYdoHn7skGaBduQEip19WJjFU9v9JYhLOWYmEl4q0tO7ng1Qg6
H4c9qN3mh4HeN+xxOTEKFVtCtYhK8h+EsZmqtpqSYN9SbxSQTBjuLAOKSwYx
mt8uRWw+6N+4IGFwB/McF2NKKfkcUeuKS13jUjFEjQp5hhCJkE4WgLk2upbp
z3YKqGEPN7RtJkNsXUkvjc1w/ZliXs3Dx9lRtEIjaIGtG1yAQODnQtHLW4H0
mVaSyQcplQUr51SBA8+Y6hipI6YsEXOBJg37lm+0tkLVdykY5e8dKwDPg5Kl
+A+JT5OxFu/dPisa1fTSkYXaniELxEE1CykfIQ3qayvQxxFRM3SkdCevzpUF
dXul+FSm0iOPshzwMDhnB+rsOPpGEGbWYKiC+iONJKh6ThYBeOfsVvI0Gdtr
X8E0+MBHGatM3AeCjuuVojohUKx6UQvaURdPuFJiVTRKq+OxnmDVpgsbk4v2
wL9Bbu7eIqvEle9SQ5zfNlU3NCdeoqcyYKw0TzW5tBrVZp3r82f+fBkUz1aq
up5rk9nr7W/6kwo6V4A9lCx4AUO/jwf/Rj+/meoNmn4Xl/CMmETBUlkoZxsk
j7jcJMiJo8/McJ+E8JZfS2FkFuxSOYyptW63qug7MGcWntpowayxlGgVYW6f
PIWdCAHOPIw76p7vW3P9LPNg37xJ7NCePXvZAERiMDgVZdhELECYPpAZGm0u
l01eKHMHQqvdSg909tyjJf+lX2g48GDuUyecJIPRsfz0bFdiwo07/BjZnNsg
l7I7bw6I0PQZFUNpvKPIwJ56st3MoZ7yyYnUj7Q7B0APsCAvczEWyE6SVLaS
6U+vBLZ21jRBqJTYQuwW9mCHZg6p0qTVAgyyoCJxCevarDLf4RNg/2S8ZvTp
YuABcZIG4g6q/fs4O220kcWBzInz8GyFcw/wJKup2BuihCubDbNo9moLlOxj
YzQPKBJpTccmIhZkAsAsyDcJL4JpFNtG8DF4MTg3gBbLZ9b+Jtdje53iig0m
Kpx6rnjqyoIl/6inlNruS9VVtvbiBIy5eQpe6UH7I7ap/Vq8jy8bB2ljuw11
LTW/pAKCEuv0caVVF1tew74oQXtkHx8FVYgWGifAC3WB0BCnEWLrrwzf9QV1
r+hHdNreTuy3TPaI1mpCgVsj4a12218uHLUxUFHbq3sT6k+rMJ4AYQYsqAYx
vjPnY9h0S3WL4e5OkBm9TUh0Ix7BMqkNYfIs+7ImF2co4nW52GSZh5wsHH/d
LM7LTQgyzyT4gY/7d3qfELcXbuvsG4C+H0yXhCMX0NLIDDrHR1SsrrCkqrUF
YWslFIRSp0oxrYNLjDyEfS513IFCZ59wCCSLNrq+VKcaJSYCpQvTkgv6JXyq
YNZqsVx15nl+C+2/FOJq6xzQAxm0lwWa1E3x9bGcDyr8a6+ToaBLRtP/8Arx
hjhkOGp1HOAasNAljmEtVR2qr6DW8bkgkLMfSTx5+MJgwCiciqqAPyMQISk/
LBxID0xEOt4S9E8Azj55bXTKxG/preS8gh0rQtTX6LHE9jyuTlQQLIPMfpEc
UZLuFniWwU2Vhey8JtJIN1KxOFfp+v03G5GBXuL8NFcMrkCI6qN/EGrYRdo/
dv+PHwFDpPFSL5XOTAgzIXCbtyU1wtN5pJS43UX/7HgQ5D9RQVwXftrMaXEx
Wa5gXIhJQvHhgNOi4f+7HqmOAk+WsfFhg0nkTGmC0IiF3XjnI/xTCMjNI4q0
WTt8dC5XZm5sB4w0DKKEYkkg3OPK8c+ZYL2ShXnbNb34OUFziHUTLk9bJfD9
M/YFxvh4M8XH9rmUBxXmOc+PVWDIwrWtLudlxbN9oVyRhYkaF4gCsLGUmH9C
5ytegMbZ9nVAU+5Io8FAIWmy0LPCg7ybQxz1vEABIRi8a1NsV1kvRgKwyVbY
L/xBLru9Yn5KmfUW7RI+3n8b/30PKsSt+oxAyvQ1gv/egSw4gUbDb0lytTIX
cj8CRb/E4J0D55jDJ/xyUCHu2SSx3HyuSkOjm1mcKvJ1plBXdBk/19gkFf6d
6XSTwo3W7UsInrUcSiHukM9fT78nOiRYgTtpRNV8Mq5bI3c28/Q5FqAmohkk
MDUt20E6aCQgnP+lgZA7oNWOkYeW0YoBlwgGSyVEZxmTP3lIaPPNCvw5WwgV
/uqmSJqawrjWNVg1vU9Oze6RCg69O/iYJPihpsCcns82pLGSPLftbSH0Vi1W
QCDe829NekYcmKY0qu1wAANbbW3ybuENencd7I/0QJrJaMneRTyPwydOL0CF
rgfWpq5IbXUH//MjpoxgS9P8r/Lm3UXLKVXrwrIxCIm+Re5J+fKjVEjZBtKt
2h3hraNUtjUCRenKNWtEBT0LNVwQD+F+HG0Az2xj9cpdBgWVyqH6knVL7olQ
qep/l5KUBG4aBomWWDjBgIxDIRPcWol6ju1vH8OgpmGRuOgW5lRADZcR6Q6E
o1FY7cgh6zcrx4mTepZ2Pb+AAexdWo2p3eeuL9syzPbu736TyX5jyAUf63WZ
ZfIq/yvnGfixCCTquMHO9UhA3PSL9oh61BHIZSYa65kk9ACsqf8OAY5SscCX
AX5D+NISKRughNEMxzKN1mFKlEORk+EJl1jnIhewzbEl/E0wtXBdVI7FaDR9
o3UfJ+eB/wId6iFi7aFXePi8Y1d5zYhdXQj+/NNqVZw7q0Vz/pWXuPEn4Tqm
erWPp4Lnt9xZFKExRluu6MTmF5EIGdE0fp7lwjgHsOXDrhgETddWVhA4QAD3
KLUlCP3RqoppldG0R9UiIF0Om4PjkSPf/IV0QBq7Jrd/C9gRxuS7UlPfy1gS
juRoVKrZdtlq45DpjGGKVqD1r6QEyLZ45WuzrOC00T9RxGKKJ+96mBZWgnUr
jiQksya6PWdF0MHWYjAY/gmz+qJ9ChLqiZj8UmthDPgk7J2sbt5OWjCO6jhV
cXJoglZulxp/pBHQ5IdzIXDVuSiRZuSDN0IrzUppgL90Rh6TIJSzD51hiWUR
5w4AZldVt2XRS/YnHiQa2DJEnQZFHNyMhGkbo9OYxIuvjfFu7cdLXuGvDDMz
W3X4bPHz1lEy3yJgFmYnBxp2/MbTdyqOWvRJQR5Vof6Qbwqn8mA5FMHNDasL
vfEJuzGfZyjd62gJM9QFexuMeHPqMsX1l/SY0D7GbpIiUiwuF6W3Km1sQzAo
Iqlz7tLzJmZTImua5PAo5wf2A/+lmAdfmIJOnjFIOinvjjVt+dpOXxg7u+Iz
INIXajl03nWHlooiL+1wFBlTt7bsz1QURun347Vkd5QgbfvhUEVE3t0Cv94v
fTa8NRiI5BC6cBWQGG9ubf3cIQSyN8WfEjh9PLMXWsCfSgfFod35rtI2S08C
1BDb7kCKhYin8PvVqe+pOO1jTHGUbNnn7AsBtJHqPe+GlibNyCjTFLnsBpzB
d0w4nVG90ZJr2bf74+h8i+j5mjiUWVRrrBPqgrNu3v/V0ZFXqEuA7UvbhcLl
YO4n5odevUn9rZvA+rXqyBqJE+uvtokM/Ou5sJvjGqObV+DyMkOCWFNPc7jD
PxvxdEAP/iBRg2ExqdXghK4e5LuJYqkJn0MPoQHIqRSx0hZ28FYalLWwrCxZ
bYDtTm7ivcFzQTSmfuCdg1WyUauX1kJWYdfGBHFIKKWsAdO6giaoOea0+XNf
GbSal7q4rKGd3oC9cjjPW7/7yu7eDnXIbV6ivJjMjE3JjZih49Oib/Li/Dbr
0sCUR+dh/gm2BDzIt/AS0tjnPlmvqSw4cngfsjJEGdj3Yp9sttgLl7o6+cN6
GsESNCbZDSxRqZkF4MH+2nGVP7xAM9X/x/Dl3TqV+jaZjIGZ6v9t1yVNDgMI
hft3uhCxP8Ys/zRCvh1CnymoD54jPBsGleAAjE95CivfkmfRh7ziVF10A63L
bpGCDWo2nwKcOQdQ6royiQKiTD4LYdHaf3yazclaBed22tt6a8Nr8tzGT0w9
9t/VYs+F+MUpy5jszCvw2BTvp5011qvPkevTfCYxV4ZypBBWnq5iuNTCF9/1
DeZ38ThRZD46Z7IaHczipU8fPatys84slR0I9XlT9lcCTthU4kmmSGfeX0Ik
s2BqSMs+dRsMrSE9EEdT+itOYbk1m0Q7UEi7Z6QgLUyASV+FWIuPvtGIcpbj
BihOjCqGLV37E4el+godAKIQI1S3/YSEQ/kD42b7FfckXAuuxkTYhk//K24B
R5+XgkqHkD+YjuO042frtUSpFZAgyTIb5876bRymIqST1rKF19B82b9ZNlf3
VdJ8sDTHrYZgsxL/qt9oHD4Uwclb4k2XUkQhimoKEI/epj+HgTprtTt/aHw1
1DG62hBU2Dl2eblHFBh4NBOAvBpeRrIHP7Td3tJdPOQyJEZIdAXZEwcM8+JJ
T5vs62MMiH9DDbcU0dy8vfi1q43UvIFKTauBKwfJHPtTnMsnwBIkcOeSbJrh
3zfhPfQz4uy1vB9ZZtIyQrupn8EZsialfy2kiXGt3UnTyVuF/rX2O+CzrPjS
jnT5RYuOnetKuNA7K9Ka/LktI+IXEWUQVh16ghfiRV0LOD83zbZ/YGnb+jXv
4Ppr0hiI2CKdaP9C6CiNs1noU1oKeK380UN7+1kWQrAQ0DLl0Q5jacor2d5B
Xu+BpLFsEiVQRIZN9x/TEw5vWGhb0nmtebjtXah+k47tT35c5mYrAhH+HQKa
XzTYNYNdVHQlL/TFKyz+vORprOvvQLxGfQe+oXhfxjvQHFXX8i5Sw3TnYw9D
2fc6kxzLpML9MusocTMXxsuhbpXOoqZXQXsI9i72JhZeEgyyY6zVGpoOLCig
aUxrHotG5tLkOiieokhdePUF7lBy9KmtWjGMgoiFTUXe+4AV6itIcAVxbROH
f6RlQVrARLnwQBes2qQsrZ9ewsX1FZf2iGeVbPBpp9nky4dnPHO61m6BUPwn
cHFFxJGmv6gJ5y7eVXKZInSvuEyLpqGJkgrPqNGPDpHs6O75e1mi+ikSABiA
jo7IWhgan5trsgQxzmvtNlOSMBNV/8TaQtG+qm4IU9m+vP/0xlQmdpHR91YU
HO/sjW/7uykvOq+hDgJPYxrND8rtYEtsHfNoj3oEvj6J0urJN5XC6L9bnbjN
56M4u1d0TR9/4GE0YvxKjZfJWGSUUYzYQnhCX967j+DpnFCe9aEgunrP78lr
4pjm9hZPK+cN2wsJ6UzOvsOORjQFC/9/O8Oj3iMbaJs3O3xb31eDhsnrfgFE
6bWZ2dLQjT7/2y433cZGEP+Trt+5ShPgPoivKAeVLPevA8yw/BznyeA8ymEO
D7RJhXWaVQdlwh2FuTpyxBsRKCja77U6NQCvySrSYD3n5Hvp5wtXHp6GmEtR
Fl8h8Iy2S9zVhKi7dnZThsW5+hu090KW9dHROfdXgyGJg17zpFl/6r4HgEO2
+6Ss8Fe1uXS1YYbsxDnDVPq0SOr7C8hJrGTmtNoACfH8kfvHHJfOR5NXC1sO
qQq8EhGw7fKef4MkAtJUC4X1f2KmVJtNIQkqG8Xah+aCWsWdUQoCJZtKBr4H
VBFebjxp750N0dMQh/XQM8y4aqHxOx0kgLWepK8g61YxV0AX4DhNFp38NIMf
yGXa4Lh7ggHAArNk5z369bG1YQ+rH2QEl4Yedv4GENXwcBsTo942s0ET84+E
ALp/wFlONdL5qCWFrFkxi6RLIXdaIPF1Dt0tz4Wb5wje9D4d4bfDkIGAEqWW
Irzj4uD+iVLvg7erGY/Lt2NL0bqNdglVcAbLbg4QFe1NDhcC6GTaBAaZMbzH
VgDuKuFc4/2VJQiqtoyZVQAOCnrCwFi1CdXoNnXMB2RUcCxzpUAw+AdtuTwm
oQ6nUmD4r31yucsdUcSd3klSreJhodaUNOOz0OR8WQeH4GeFoVNIu8AU5Lvp
Ep+MA+FCY+j5XqM2CW+9q/nPyLQFPujbg5uYnLGWdJZexLPTP1LBadZJXt8e
haZVKdBEica4UKl6iIX/W+IUkW6MZCPIVChVRymuh4IKaeaVUs7hOBac0x6u
aXIN3gmkBHFTp1GAvK12F+UpiGBxU3NZL3wqy08CYT9R6XX8hpLEm4Ck8Aw0
4EiCEK5RwcBGnz+Bf78/P8fASo8wZY+bVHR5Gvq5pFvAb83Ak0QceLLqPF5d
1rjbUCy6SfbV1xApKHTh5FF+sDN5KfkVF/rZR8VnH3B6mPW4tqKQksgTJBRt
L0ZcN36jG5Ah1I4WA9pNpm2XbwdDXu9OrvB2cetfduG9jzgR4hIvnT2PCCQY
Ht5sqWZ+9pXcsqf+7zS2mHosepILRt28e+VmqBozCWdWQV+XTiZdPnJ9OGqr
MHNfeGSo5+biZVIF80dqpSDfuQWnOu/5sPZmLZhrrP3PXppCCp80SSrk4whi
fjVYnf1bkZW6MysVXHf27ag3OTHodmkC5+vpO6lgITz1MeWddAtROFWezh9C
ZKukf7lnQLn9Fk3Fez1xkmF6hQigW7kIDwuRU3o1YrzqQPBvIIN6j2m4wKWp
0+HLUWx1B+W5yzjBZlHpRQgLnGPL2PG3Q5uFps1/2QxaCnW1zsO0SFq00p81
J4za3ftzQ8vAufTSUDDCkBTtzpor/b8UihY2bnoyEt2uonrMZ4VAqs1J749i
iOVj0x7TXhaOoGNK7/bQoMqa26rsXkHejwzSzRYwNtpaBusFfJbabIZsoloA
ePAKolqS+qcd+XMYwyXJ/sjHO6VEmkcOV7jzZph6MrkOM47qosXGpVWkeYnX
ALEcfmqcOytaq0fxJx9xAWVKsBAjrDLhFZd2dvjr1dYIrmZNqV8XJIGWYWc6
Ze7/he4V+h+4+7h/wu/gfVdQiccVmCf7TMjubWFc/tDbfwoRWaYIjUdhu4pb
gkL54vdgfqtQPgGvS3+vNi1ge2JBFQHQ7+G1xWFq293RASN4aQedSRO9r/xR
arOmo7PL6SPKozMjsQeFJvfBibgqCfilH3YGfw2KwkAcZwZY2p/zctkcKCsy
C7tzB8x8GCJbVivtS52I9Vq5X8wFaRxCbQ2RWOQ1e8vluYdpggFxdsaWoGrN
fzXAxvPADlCi49aEoou6RFR3gtsE1zbh2kiLChoeFyerUgsuqSMC9/2kDiyt
kE1WKVEVTjlLjjPfUV5q75lvorROFqlDYMfKAtCYA/nuv509TBtRAKEoCC40
SUzviRAfX9i2ZinC7w75O8e4psiDz2fSXzPllBU75RQ+j+mEh69kSgKd8HYx
2JsO20ZhynE8ITWyU7Ui5oA2fFyHa+O0T1PCr/8R5BhKgssX5NLvk+AszucA
JI3ALWv/ki+YCeosTAYR1c3VCpPf9eM0jAsyl59Cmx6GrWIWXdQsITje+Prr
1mt6RaVkA2yoXu6i7O5p88FyYJNUabbnzm2gPPOcwnEYoqnAdJkluo465NO1
yd+opV+Mjx9U/Kx4SxSCjVd8+Ap+DkzZ30q2N/pzHyUszkP8wXpDGAwORbWf
BcgaK5SKwpyGZp08odw0daP02jJxtZ9n0ex4gff5oF0FsS5HmbSj2lTbMfQV
mSUE4izwoEd74R/BkcPQlD47JaFvcnXWNKRVwEzl2M1H+h1ISvZ+MhX+b4v4
h5TKpHJK13DZ1Ir5TJG8x+Vf3+/OfTowGgeyOTkUJOsWz/alkad1py3OwCJD
rvAK7WygpIZRCNaupUBB7ZShEb5njlblZ4Qmm7NOaBU1mgqM+hBjXhwcPmlZ
k9LklAsOzzc+SjCQeQGJ+Ulz8L1ERHALiiwxND3R+M6PGUBjWF2larP0Nlpm
mVxdedUQsunFA+Uf5yDcLNYzKeOnsBLLwmLDKWrPbDnASpY219G2tqq8E+MT
G1eO8HgdKe5zxrX9eh5x0LjKh+7NuY324PUnIpFsvW6W/JljM2AS/qvVxo5d
KrG/9xlT7lAlVnaMVBFpyZpsi3RMPzBTUvMAhuohBnAXvImS+E6JaEqt6JIB
2QeCKwNVRjdja5MeDz2Dnw8AJK3gVZ98mSeCBBCBXfudhEvyU5opaCPiwBOs
pEjFqUNP7adTI09znUxBetU4R6svq4Xv8yK4A9rDVxmyZ/nSgT7RMycRdfF2
YkEZjBtOurEiDBXhvOrEwU/ZUQx9pgVjU/3zVkI4HTgf2oGURjts5lewZnhF
MgxqHfkNcKb/TRDiBx678zBQXxERX73sKwORMNUOQxQrWczKtcXq84wVi86S
jYUI4n4pa1SEmKqZy62Cwb3+RfP/ANektRsZJkxxqqiRbZirqfIJ7nMj/yh4
uwu2+LglhoMf6MDkMk/XN/VWUkpTWWWOJgoN/OzgQISU0AzqydFjiwkSKX11
kR6T0PcBDXZIu3iJr781/n0p8A0fyEmlglzhZa+C3gQCFXUrW6aFzP7elTZZ
3cmu86n46to24zhNDP3eA0lyqgmwLyZ2PSTIeJyVI0smrkL37nfEliPeygLh
GwgM51SZGJnXCaBju111gj6j4dizxVEHltxTIl8vNkz1ZnSd7vnTQLWyAXm+
3CHyEqdZPkc4ViJ5AYJEPkSaEwkQ+0rrQ0vcLiXX8YCGNz16vbZl1P9bGcEV
nBs8piSBqGfIqlB3sXOZkZrMyNsDmNa8rmbuZQS1DuiZhfF/RnwE7OJb7JD6
9MfxAu+Dcz031quUsbWpLWlL57FRpZj/bIziF1kVZtXk2cuCP3uXvIw210n8
FjhOZMHPQ41yUjkWdM3Yjs4yMDYXRhkZwPg0kLDz+zUIjJ6CdiM4FFndoooY
exCD6Y8qXgHAVDcFwUcUvtDhcEKbHfWnLm5o4uLddXBP839rdZrIUktPXfKC
6lo2foSZUwgWKPt3ngEZqYbql9IPCgwh46uvSv4Y1rm4m7pUnRIFa4s3nVTw
B0f4VyBGjiBcde8ICX/4HIyyWllVFbFLmPx1ge4hqH7K9yx7RYulgOouFxNe
MFQUZt3yb/BU0melHzPO4Btu0b0JEPfINnWd4P2edoejDJXISaNW2g8jtYyy
rWHlku6FS+mp3gl3Y1P4ED6yZ3TZ3Ny63tBrdhpiZxb4V0eG9o5mlm+BVCqJ
kBdrZPfQXsdLw/JsGoKd+YxU6M/LC9L0IOgzd5OF231sl+1QI4sLA0hDiB6U
11sJC1QyvabLlqS3YglIBCHjO/l81guXX8i7mO9cujDMh0d91xG1z3vC9lEj
F/puGmVOX/G3qnQDBOd/18nTg8w65zwHoRIySfPQtcYqjvXk3Fe2TgcK31VR
xZrvgBGHxE4tDu9Iz8zkMemRnrOqlrtXlkS04ddXb2Wmh2LwFmxCQ99SbBqo
IcShMj1U8wobfVkASd5aB/Znh/FqXM8/UdRbyVReABtXAytmT136Nd7wEraI
5xexeLiFA2a2LihuiJPNNAMxkcT4dDrjc+uEMC+EaBwNI2R7Eh/ih8Olmy34
ArnXx3OmoSHp7KdGRSEJz6HLdPQqYIUpPmZ8pfI18tkde2T0IDMhW5BNeHqi
qEBbdLqQDJT/MB/k9D1xRVHEVOofL4HPJVgugQcEqmzPUqQ8N+TO6m+xIcBz
lK3R+6ZNRb0QUu7hgEeAM0JRdxhfDmpaTf3dLoUoy7qj5UOROKUFyMUjAFss
cq+WNHkaWMHHMZ2J0oBOcJt0cCnSdqu6JiwWAziKsMQoNmdyDQqoHs6ux8bP
WiHqqCz43l7/6qYsd91ftTrjuzXFb9C754XG4+0TsRIXGKOiOLP+g3LZgKiu
m8/Um0slZUIVqRu4XJZ6Zq2E3753AjQC9fteq7vaVr2UyRlvHPP1qWR7/Pcx
28L3xxTJoOlkgZks/AB7kNb7BecYFC5tEUXCmz8GmQvjtcH2gHapOUKBSeyN
9Igj/Z3JvW0626IrLswj7BrNgBmBBZbXsCuNsnVbtOCbFNuMntVe9DWAAuGj
mrOAVWm1DouEG74xRYNLyBxmXL/viY1OH/lt6Z12fnDbKPw95/cZOUPF1leo
cxcR1Kg5b6jSM4HubM10k/ahLy/bUhBaQPlfpA82uA7pKxsMQBFmispSp0yD
k1xncpl3QCBx8CmNsMosxnCgp0KACr6/tG9X/2oCJniQqFM3P3kRywNCajhU
GVPcqnpp4xoOQCkfOPbb11m5CPyLRoy/AJMdMRtNeixVt1lggRkL6PjEJzrP
W9LSOD5BAHFYwrigxNCk9t/J+VEyaDsHf+ZyBcBAznXQWhiOJbMot7XbVKHX
ZkLEn8gNofRp22DSdmF/KI+6yFSl+M7+/bp8ySSdPa5wSo/+KLbpIdF10X7+
m/bPnYz496gftyVs0JwDmB4nRxplaFqLmpctXbrxDAOsws4Ps3jNe0Y/d6HD
bJ74hBDHNY7B/vh6+jGvAz5Xrlx4CUKE3jWi+WpKMOpaXUVET3AkFB6OoKb7
gAU/rlMRcxLYZrJ+jJP107pNAaSZYHLal9ypPleOB6yzLzlkOsGQBAR5iNyV
H+uNF7cuQNUY/kaViXPlwqJNSwy58jlixbfwdUaFuIuL0fz/JHL6mJ/HVyDw
TPaa4LuGvk/B8CYf/bJqxZxvwWJRRzeVgPmavuFg/GR/69nErvUBOw+8tRZi
w0qZXfrya9p/tb1oYRy6fx3ztGUBoEPf8ta4VSPbN+ju7tbz7uN9tCbppz4E
PwaclHlQgWC/bnonZXmEjFTawciBkm4acySIceNdJfVvzrxOqxPBP7dzGYdY
KGL9Pnh6zqoOEVjG4qbhlV9cMQGlzi5V4d5Z5kFVXgVamvkaMuKksRThifG7
v6rpOF4B+AjcJawtrKn9Z3n2VLxu3fOlv0lBX9WBaPaMBI7+nuxHeTS55bOP
ryuBUjhjjQGb+hfCHejEJejUd3Z662fyQuQ/7Tv72pjgmHk/v7wO607lL03I
Ql1IG4S2sP9xLzepuzgeA0toWHqJQS4bjOZPYaQmwwzqcKRnNAIWvDnQHxH+
T5EjILZK+mMVUgr/77bG7eslsrCJ1Ok+BQJGdSPkyYhwEZnmDKCS+uUF+dro
12yR9Fyjm4f0HfQjbsyr95auBC1+u8tf9T5Lg6Z3O0E0KgPqhvhbvrKSd2EJ
mFPXB7SlMqGlvEo38afG4Aft3Yf3v+IKRXA0jsmxAL1NmKilfgbTBIBQcqyw
a7+uGdboqrfMhrtDUb0gmGW5vw24ML+4atZ6DBb2RHvl0sy40yhZw3hgyANS
hfSYbQc4NC3gJnY6FQsXdNUSB/dBYAsvzFORrZCioiKglVqaN2LSaKQCDIwh
XFSnMXSICwoZ3dFS+nXUqVF5M34kSzsyEVfoKW361Lm8MDMoLxxrzlRprh/P
s3X5EsCxzGWfm0KqA/oZT+G0RE38t2GxNzH0br3RvocG3D0tVBYJ2LsHBtNF
8J9pcAOaQhyjeM7/WSg9sS0hsprH/9woTOdbLCIhuboraH1dvAfrlSlifkS1
SBnRBqhBG9olmlZtDuKFgBUwyNMFw6S4CIffbf0MV8fBEYiRBq4bpy/T8YD3
dLzo5kqxUchTBawhQtu8Uu9QhbJLxOmjjwSYOU0qgk2AxD5aVPx0yuOx1+r7
8RERu4Zsr3fztHFM0poTBKbPbcAik2oQZvvaCZ4Cu5K6ff3Lo+BxOXh75wNm
4cQ337aSPzW/UTEiMKcQrylcIFt3lXuNVXka6bPbm+YFWjZ71mMuhHx3JUpq
vOg2Mi81CTo80k7RY6UMo5QJ7xIZjybWQgZWV3eUP/rgj5KRQSdGu5nW9Bi2
sNi+4tVdfW+ONN190FeZzhLTEPn4M9lXKxZHQpUaBJgdtTJVl1J8z3/FzDpE
g+SFlaAqOA0m/0rLLJbxySdG2eSw3grNer1Lk5xi661enyDrCSl1ye4Mn2Qp
MPidy/92b8MqdZ7gBmOo3PSrIa3HqwarcC8GreZMCifRT0nNAiAn5JKqM4CL
VD4REk0T5/wLv7mPyLTtDQT6SeuONOAI721HSHLQkMz+CdW73P8VAihZR8ut
5HjohE1XUUjdK8GQ1KtQdVkwoDmd39gTXuCGpsD4Qh6c40Qu9OK4/WTX7Wgz
arO7XktjfBnuNY1ZynjZGC+Aihkr1KaP3lWD9UzN5CgVTfn7uk5zaqEZcrPG
xwf3qbmPozYMg2texOwZu39mSNnYH780xusRo/66/t8ZSX3H7CUpVYgm3RVo
tdwIvEwQ0ZVUd6gbuYFf6AL1JopxcURC/1SCuX1eJdb+NRNPPQB9BoJ+4zsG
BqlEnD/UlfEFZEJiBywhyX7bMEaHprVyU9sQk0v1aIbhxJqtELpmKuYiVkj/
vRIHvFJzOSkVMQlosclYYSoHt8K0yKspVvKScWPZjzoz1sD1UkSYXvS8DOiA
eVL6AdLIutS3+q/pOs4vX2KFXSWPN5i/wFphZT9wamqv6YtNYF2dMeA/AXyk
NbuWsnaUL36P6iLeK1TJjgxKuxs1ErlEd+BUif/GMxcXnFRxg+JfNil/9fYb
MfvJYNo5A6IL6Wua0cJBw+luaO5vo4nATrvfIWh9PtX+MSbBuGIi+t3w8B8x
Yc+WnuvQpnGiQtTBF/Z/f+jHZmB2slZR4Ok1TUzDpYOaIr4PkXd40ZSxTh3i
DvDeCUsW93aq5jpJC2dmFylS39OS6bi5JK11IKRFlGRjKLwuo24AvEnk3mmV
MOpQZAsKeOXr46kpthIhcrKmYBpEAUMUHjSz9SmtVBIZj1ng6zus9RhSFvjz
E3pUZzuL0hUdcFgctTuCLZKtOLyHUCnRcnNuWsgwCeoTyWW2nIi/+UxdH0qd
TyZsems+KAtN4mqQ4wCmfxfvODEBgYk2NjkuSrJ2xj8EkVlGz6TyQqCE2odL
vFS2KvKW2T34l+xMXenXmsx/exS1+P4aS3vM4rzuISxjFC0Lv4BF55Fm+6hl
5TQKIeucT3FmvNnoNCih6BGKTrKvF/DnBYrFwh4ZxFI5uTOWgfzBuqJHC4kT
Ubcd4YkCWR3u3HkBBYZjQiGWo6xmXQDnx8eYHQE9rggQ8igbqidK9KHzfkyU
42fmbPHBhQm4yjOgoxQ4EIYUPKNZME4z2++tGmLZavF/92lGq4D4P9lKpU1r
VU1z/oNOSNsb/3YfcBIdvfCzBd/ouDJkd+qlk/RXAid8RQrj7sz7aAIWjJQZ
vSBqngJz7K8dC9Kc97y3PrOcgD+c4580AzZW0sNOt/dp1HlOWUIMgZN8mf0n
cze0S6d2T2HX/0fTG4z81lYotL9Q6qQqBy6psQkVWABOyZn98w2n3CY8eMEP
nT6d8tVqrrwELRs0dBc5dWMG/bZ9G1PD1d6/gniyTDLuBPvDOI0O19PefopN
60CrObSRAj5FLRyj6gt8kmQe8bammPjsjECEa0RlinJQdZ2XFl6nfVarlTib
Zi6LQiXYSwpuDSKGpYT/P+IsmveBg0rC/tErwcLTLUm5s6INj74gvLqryoP6
HESUbt3TElR6cLZ/gGvCfAU6ksVH9Udv56JSkG4hFR/OgUiqkZ3Frx/tClY2
mRjxcggXv9wHtXVBQVgaDU0+eGeg8PrL/vL4qrpUxYkPLFDa9C86x8VzKB7R
AB9FSVrEIQQbit8J2A8JoaZ9CrBrNpcxAJNQxwYRniGG26Z5q9WxuEepjM4D
7RLh9XmTjpKTCSTSJr7C2ADY9QgSjlhxZVJjCmzZswB+pT2EyuoIO0FieOZD
TGx6Hz1s623E0kDhRLSI7j1QHNOsdC6rVjiqfjDOZTi+g4PMXMUz7+pCY/0/
lWwd1bUfwXhzDGzI2o1Mf7FPB+LnwfyypsnhshZQUutppOjGLMxuiSZ5I7Yb
7inr73ngY9sLuszBiv/MtY4ZxfBIvnrg2VhvsPJ9kjeSzsZTzt1iu58u20tb
lHTEdRByDrSuVnBXNk+qbBj4WcDWSJnBubzlU2iWXkp5qjrRIgrgnvHzMw2A
etzHufv4qAL50cEB3nG7VR5R1Wxd477jf0apXpNASAlhmjcuppUrcw3jDChS
Ap7oWv8s1GqSihFlsRMrvPLwW3PNprZbuHOVTwtLNkr8JffDImZvOpe9JFcr
F6Pk4wXBxf9d+eXKuSRXZqCacgGIuQaZxUNaCVgOoklTAhbEEk74Vnqp1tuB
K4OH/cAA+P2sVeAaLcG1EQ11lxi/5Sw9I+D05ofbUfvpO5C2wcQpMGfJl2/B
Ylsnal68b+nkea9YD4vtYDAbDbrYG3f76FSASazhHgrhcPwz71RsOuTM0HBy
1joy8atikslaI4L8ImquFBtBJCTv0RncZXfhJmRzqCZ8/wG/wIpuVOGgAPOL
RWf+epfOr8INDjUy7eUn5ZT7VY/s/ljwaaKQszOTB0WcpatbNFjNpQpzcUlP
gEWzIWMcjd2EVpPUhu9tTQuyZwFLkdaGM6LnE3YFoM/EpBGTm1KBI0EVcLKw
REl1e3jmm+RIkE3atNaLgu0Shwb4/CJtPDhaeqCm5rxWRmuXZg9qxjKT46fN
IkT+4Tur4bWfub7Ypbf3c9gig38I6Aqo0SsxagyV1KcjnF9FyF+HLrV6PsU5
0jeffwVMOuKYsJcgq/d7xmVgrzKnlLYg7smv5/uwqO0rERhOqj5UOQZELT3K
P9t1TBiXlHja4NF6HJJQH3U2Ud1QkBHEq6kmStrb/zQFIWhOAlFAELv/ikg0
eTiNBH6lbztcFl/q7esyhm1x+4RSeVSAf9AF8j+DU/RvvOB5AUqEbLM4rhcS
NFQ0ZKBJQzofQvlinNswsjdS4wJX1HQUgkB7mk8GeEbEvwRSB2tYtKIwrEVH
wqyZZQuMeWqUjvQtlA1Lvon6B8DbHKOoH4cCVhv09i1cATBifRqV4wBxPVde
I69jfzHh2OhUKnqeaWl3Y4n+HLN4UODQaW+K9AuTtCJXz6ZXQSHDWn4rqgCf
7ELwqbGXFtehWwMTUP+dVrCJQmMkvjoKaoyTp77+8uiOXYlz59Bm4C2hdjeA
+eid3cz1hfMC5oGIrB1HST20Ou3PNQyAe/zifK6fyXr4ppeqYRJvEhFdFD20
pxUaEaqZu6KKtRy9tBAMrfEwQ1YivhwK13vWJzimRnEHdr9ffUTI2So0JOOF
mxFMksiOyMwhkzLAgcsQFDX8DpcXSLw/TuCQNNrRkTtZOI1FQtB0/uVB8jg7
WByL+/H9W1R207xFKzB696eVmqvfftuR08iGgytxiSDKOCf+4tiUCVk0gvin
pfLzUo/LebtuS1RqU7LYH9ijtCss1MUJ5ywB97JhBomoe0PboRUdcj7jMHKH
zS4szILOOX9BwdJD2zET3wrGvpCCmebmi3drM2nRnm/nUBHc5nq3ptpSGHnH
OMwTWe6d6IwaeO7CgVorEFHDuvc0ppq4HkqWhlSbhsF6VFV+TpixJLhY5LEJ
3zAh7WfMs4L9j/5Ssi+hFC7ntEKz2O+GZShWUaR2y9HPMpd3IoMjPEYLbNlK
GijXhNYg5iWbQ2f5vTq8SvpmSp4tgWRxacf75xQKgBFZ4akP4Ck8uSIgVQGE
ykrRpVAoHWVhI6gS+Qr1HEg/ZppbIhfKSMGE8ZcBYVAxw89LACbQX/rXj1P6
8IJTMisSsZ1Aw47vT+5atAhr+QRCsWcDOyilKADWv6MeznPFogXHzOHKn7t9
M21ttG/BGw6rZoOGmJKEcVy3KD0CfOkd/OCdvCtp8ZfxPQ+rYePHb/ynzpBt
iJDR4RsipO5tkCCWT3UgGQ+P0S4m3lf4Ihx8lBemB1tsbd4P4vmb3pMQPNYk
xqjYyCA4JELc1o+SdaZGGI0bq4w92tjdMHGWIY0NLYMyftr++a7ndKzOKycl
WQKLOvC0tsDq7+qwZfSJhi85sCTVqFaFGelpcP8NOp8DeMEi3nPeo190XScS
d23aedo0/wYBndsmGXecu+JgQy4kDPK2xuGne3+JsQCQmDrrjXZ3uHXY0u36
VuO0Dy2nxDwxw334XiYXnWK6n9u3b0LC4a87vpD9Jzdg4VM7iKiZwHhn6l7Y
d93iaBCmOOVm1bb+KkR/s1In3TQWbyGfkdcxaqmR3RpzpOPdngBrBzfodlGw
lToDCp7J5EXyocZY0t2YfFVApKx9ixin8mRPpl4W9KRmfUjTiKahMSCaSDff
B9ZuAxfv3PnrH/+/ydnFSahCgBsgV0yN7IJHwfxN+5CrQuEKqqjkJY5tTxVv
DIG6xJ/MgI2E62vw94p1s8ClA3GxPhdnOUz3y/wZ3ZFtVhjKdRFYyIPm4yHo
xyKncbWFLjJlRJudh//HfZRuQkNtOCfYow64L5z0o6c7feNxyUUW5450XbB4
nuWykcH2IX9AdRm7LdIF94iiok732La8ruzebk3S8vWvytrMknfY+su6VXmW
5HZRZrMQyk5+GWUqkreJsymhJRuXUlxVlx7F3k68LU0fYlUtZ3SM0Umo4CWE
NN6tV0ZqbJye0zHNzXTzVQukUpjuXk5Zf9hTf5CvOFCTLZ6bPuQYXzbzsaQl
bVUm8twq6BSAmXyR1IWFgVwr+Ye+lcUzmhe/MA4tdkMx4bqU4nRDO+MBd4TX
qy8Jc/1kShxI7VKfi1K+SRnDtj7FsyOeIfdjFF2VdV/0tH8iImoi+KnB/gGp
AEh+lhN+URqX0Au3s7LfClBT2S12AQrqtcP3ZZlWgMygXVnce4bWiUuxGmnX
XBSjI0GSr5MNgXxqUsLACxWC9nkSW9WlDzp5452kNFGnkh4qrlh91qmuN7je
1jJF+/cFyFuVvfxIY8YlWVRkxiUOSMtUtZ35K1R9viUJpwEmA5cQOKh6NZ5p
eU2VEl802tQ27RiYO9bGLnKwLTpmhMVR1DLXNp1X5megR/86hFJK6oyiB+aW
5HoPE3NVrt61jTFR0N6mRKZI4yl8ivkhH9opaJF6Oy+NXmDu7yJB7Q98mpDT
/AqmjfXuJtqcoWy55yNiZJqzwFk5SsQ8zuVa0fwuBeFvM68mbWlmaOkgE2YN
iVTfMSNA5e7My+ipvwdSR8z9DUHUitODHQZruYZcJlLdXP7xKOM6GeNZw6mW
1iAyIfmjJTfz5/wCPq97QkVtNR0aZJbaL+utWJvnT9eViTNNOjCKJaYtgg6C
MF+SQ4sdfwDXhy6IXWpE3to4N328oydfZNBgkL/KIVUGOCF1xvN6q1o71Kzd
TX2m0k+CFq3gXesSSoUoRsnEoMsykn3OQGuMgRuel27g4v8RUs7q/AfJwDLr
aQDrzDtGTydfGEkFEEsm2hS+tNVpsSraINUyOpwjz8lDAebKPQ4UDi26WJmi
4rut2yy8hMT1WZkSTfUV8iyJpY15kw5g/dc5upVix1xZKwidFKQqzR3tZ1Ow
PHXL5Tjyq7rwgfaOEAh4jVh6Ll2+VQaHeSCgWbIjseo/2QqbPatz/q9D4PE2
NcJHJ8dFd8IAADemF/2swypIJm605+PEphkwqsbjcWQkJweQ1yonCzNAkREJ
vA06q11626chFXqlnJxGPDVNb1mkNEsZI3O5HgZf8HsAwCynVdJXDGDolPWq
xsTne7HM7NT2/mXg9xLj1pS9mYC2jlzwgZDk/bwZVbPaHRndkBu/qFh4WbhU
uWw9QMEDcoRFNT1lGSJMLYcMlSpgkATxTsS+PmuWOBT2d5BG8Y0ZiybPoCkc
tSOfLzpSE5w8vLR2qlpxuTLlr+G1ghwlvbUUv14lajRQ/9quXVO3oSCBRqwa
M06N+VFNNOIhXVZzRRmHgA4cpDWxxPrXV/FdLZiJA4hLOOjMIpBX4HZH9v+e
MKwrFdXphFyMDx70W0D2bemo222ZJxaEH31FmMAgfg1DQa0jpkRsQtp6HWdH
9uOynjRXEfGWLnjKXTnnVRW6KRJUxqMQMgEwOR9uKEr42/I8SzmeygOF4sTb
trLv2k3RqCOcdklMV93h7pufN1vK8QCDEa2LCFLzrMttvKApmKwnqBmfpNVG
406PnRU2u9tO5zsK7t9+GMJLzjI9rc6yWWZk4bS1toINZNPO29VCpNjtQjcD
qf1/6m1UqH/z1VW1I65/RfN5PWgcUcjYRgWfnt2CtIshGIxUml+GJvPWeNow
UuRk4uFrwHkAjKv/kJ3a6a7lv6YWDZXkVaC0Fxg0iO9YKuggB5XqFtF3kCMF
ReqEpyV6rbuhAR/6rLSXJOOonk1G7BlFipxIqbN85v6uLI8zwi6I31pDwf9m
FEObVBQ8h0UVGtv74qP2bQevUz+Pe2ZyyIYRCu5Pyv7j2RendvaD6RIojVUd
xDre8F4i67QGgptsZcZzNHGWzQoRChxdev0VLZcUN2iqgn3GPEVK5mw1TmrS
Ogp4Ay2DjPrFPemqzGdEXWt/BQh1GR1+twQs7/g8TzIYAyV3rMCtnV6uOEV0
V79GkPvdxNQRET2a5/svqkf1u1EXiqF0rOLBH2i7CTi5MtgCnhI0AnDnXZLm
Ei3XMhry82uQe/JBTWYoQRyqblw4yFn4U9LXgMU3XSdquZs4GzYlc//7M7cu
QXZ0K6a+Dj40YIvvdJihtWFiya3HTMhKmvr27//Sdw17bpKnDADYNQ5D6wG/
RetMdInbpwwuKoM7G/FerJeA7JUw9BrYS1lM2bd5BKe5Pl70DDDK3kQBa/Qg
4eN3NJvdPSn6b8CL6sOGc/iuvMlwrNza4mr1hLEpErAy21lLpxjnMTlXgkW0
tzxmMGrwISyLfsvANaIR4IR5GIyz0i8xwCulbMZKyhQBKVUnoQbt4xVg+1/V
dPt905Q0soz+MeoLA+agWz1ZTiMgn7wGuNeff8v1kHmzeqTj0xP62wA0Pqnz
qPCWAFqo9aaX7dJA5vPaZdq/p5TRP9PqIUpGG7prkwqWLq5z/+uv6ucSn+0L
Alahg4PByp7rLd/85cA83VYgj3IETmHiTZxoa9IBdGauS8aD+ReGeoPC8kfA
xmuGKzHK8ALtD92IHcCQwuk0Oivjk7iMfo+5f6iTYmBdtGhtvxZQaqMDCsG4
vz4r1ruLhvkaRLYKExwPn43QsoQmZunjxM/kw6kinRLcOaYf6dmS9AV4qKf+
Sxjp8Nwc8LgHecVG+Qp4gmKoSdyzAOvgMxytwnw9amv2v6rOGtcbvCySWDoh
QCg77DD7BHpH86yoi6zwgDnmbbkGZqi+h3vp7p9x2k8hl4lKoDnF6jVUD0Bw
xjrXpBZDRcQQetuHZAaZRUVhAMJ6p3m3oMrSKgQIQ0FSt+hx0zAQTHVfqJvt
4lmVjjEbSpKNRFYMTze2K4yBx5+3oX+p90TSUEw9fHRomGFb9QDhzsSX4nbE
N8myll9qMEOWcYOnPA38D0i/Fby/P2iS1V8+ML/dyCIW7cOS8kvsXkX6HNlJ
skH6UKt62R5/oHnREuq0BcPwtOyI12YEVNlZIhs5Uxb0NPhEFYcAjdCLOZPX
fZDJ7DvY8PpHsUN997vjXaEVYW6c6tEP0y1lkKnet9K6hbkPnJLrnEMJvRlf
I+CmtmHxOmffqAgprMSyFXgW1KcbcwYW+dd/BQLCRfwiTMg7cKCdCCZqrU1X
ay5TG0ToldKjiGS4f6Yj3VP7bfz9kTrZPmVN0BazHl28XzsKbKezrrMwfJZX
Z9OCYMlprlLFIFbpfR5I0nwOnA/Oa4EUgG2P5yutdny2xLsChMXUyv9InezA
M9D9aynvlG2bmeElH9D2nkN8e5jVmm7GbsfJ4PEbcUXGzdwwi5tzQ+gERl17
ieTzVe+Kyi/BBscxnT8D2fDEyNIN1o1HIe+34gWfoUwjaxmM2fTd41m9e7ua
UYpPjDPbv6C2RbxfnpIYqCJlLtEpAI3oWw67JHZQXH2DswGe0PFZqdq4RoZs
9GOCUwMh/Nv7b3WUycmillndkEWyyLERv3SrQYC2U4c6AW+OemSMcFCaIQ4p
Md+vstEVloZJz9WZb+LaJglr9ou1sTBb3HBGdvneZDn8HixvzOfhOUvK8mf7
GlghSOpsXRR6DuId8cToA8PtqhgWPbpFP0TvRWmT5pC9zc17mbnp/Ff1ZJKG
nncf+k9qFamfOicbm7oFEBiLK2CXhPCRwHyE5BKvBt0x0uz+kRbiZNRa0LUM
M0T9g1lqGtcVIXa6mCZpy1pY2Y/CALGEy/vwDCsn2/tVJrz9uwEiovYSWRKW
Dw8WPKLinzsxfR0zdtS+/qA/GZm8ljVLq9PFVkkp1loRsn57bkK0Pae5A7x3
bWrjGNerg2NhBRZiDRy/ALDzRWpNA8omeGqDSHDCkM/K5D7eXIG21kKQeh66
PNpfWAiotZUV0rGXG9e+goQjDHRp22B7nc/QHXrCpG4kI6hWYDCOfyqPZ5ew
bbRzcnYFkqJgxQjoIkqAt7FPLbuuAyFyc+xS1xCbWD/8yW1q4PQ2WmjG5wnE
c0Pf4M0RTOyWvy572suOzxzRLGbkD+1npJZH9rCioEhhPa9fMcKnlzlzPDIU
5FN1/lZE31BnF8Hb3JAiY4icXjT8/5GzUIUKpmzmNo2Yysp4AWvCyNgbTvUx
qnb0S+PE5sARoxcYuDQ9UNuKMN9xr6qI+uXs08qS7JLrdtQG/QgKguPIkMTv
BDkPFs0xi6+h7DSF4WT+s9+zYvnuesSzgooixtF38UJq3rvKdzq9FMJ7FsvZ
50y73sd1TgkdSMn4MwuiJ8/FI1qK5DjlmEVecw+W+rdIpD7m20UDBJsMX3AL
Iu4tuhkmqcxQAcLQLK4hPrz02ZOgBQc8L0PQvLREVBOKgXfGUJSB4+itFtC9
qN3gmYMuw6OVOPdtHYokLEymHnDaJsz0Ec7+FK629Xe6ctyVkZ29M/+vyinf
5hHDQ53jZbZFLQNwRIY/9+ZzzRi9cxbPymh9zWOTG5Y+raPMn+VnpxyUfaUx
zSRZn7TZ0PSvKJzjH0eFFr4UDp9mjDAkY6QLornWAQNnpRb1Jcqg7Cng75DL
7Ww6RGnEYHXzp1VFuBlF6NeuT9OuSe5bWHO/mmvlTaj02TY5PCb3V0GZ8T7v
oXH22fImyjVli27MC8kO3F/fEVVIZbaOemU55NZCmLVb96UMIaTbO0pX+EOj
Duo2Yq9pjPx44t+4s4iKqg7rJPf5EgQpDOeIdTpEyuyLuPK8/vVPMo3RWOpS
x74Hc9CnCEezCLZqfvm6LmMpeUWK5H5TMTUuQsvHHi05mN/kR9drCDV9mPSH
lopo+/rKfemrdAMaPzFNDYZUwjZvVMYkEZ1h7q06ken5LK8F7wPy5B0lWif0
NVuVktDkG2YjN5xLTqXLhS90oYrm6rBnwcDufzHGWNG6IYtW2C7xdVWRf8o4
vhM5g5MnbGBKhgWUD5xzFBZWkzfinw66QgWvxVxLI+P31/xyNcGLWzUzrtIp
beHgVM+0HDUk3+BlBfUvSoUdSOgkj1Jn1PQ37zbVHj3T+d5mryaGaA4IT3r+
bbF1JnI5XD6xKuCEO9cBqeeBeC/ww9XCylqLTSQUcSDn692u79lOcrCel8JT
vTVk+ijG2eXvzKEuO2FJD9T5RYOcwMVAGH88mcPARn7Nz/pb7Ilw6fg9Wjdn
7x4nlyzuk5kj35F8Xu0mzl96AhEWGvosAw6AzDAFlT1JTYYI4D5b+Lihj+vX
RkB6SsF8UJ7RzyBitZyK+rSRMUk1UPowKGYmFtQ6EJVW5+fy3jHjtPeQJ37r
2ysv1om36l9rn9bcaZzH44+m5TWqkiAInApO7M6EANPgcyvODLPv3TK+Ah3v
RdHN5nQug5n509I0nUXuewYnYx5tFIosjKrZk+XDPW92zvHg4rYoTQGne1tZ
Q7S84jZhTem73Piz//ZXH/eXTTT/URlqWVzJpYQcFGXPVcj6P65QETTFlDjv
7+7MN9KelA7tSWDZ2zLUo2SWVzlx3fKly+w+F2eR5RQ6ed1j2sDtcaD5Mxi/
eulwT6vt+c+2VkFiRhTZDJhDnZkCyXNYVogeyubksEo1hhXKtt96jVFWnVh6
KwvSyxqqFnNRyHAgQIevNdBYfmdlssON33RUhy20979V0PCqMso9ZfwOhK1F
x5yxRG1RZ/QTOiS9qJfLYxX4uBZv0hqAcSupK2uryfdXdwV2xzH3dOM1hHHT
wHhMmjMnVpH5gl1DpSPE19ESP0vYwrt4H3CD61MyX5cmbhJiL+IdXYiPBaPq
1lu5S/hxGwxmTtKDMKWP8XhFvvIi9HVfzw4eZ+7cMj1A71rH5Ou6dQWh/KP/
jtlNddIknjVIe75lx/8rELd9LmXhBlogy3YjR5wWI2Lbe7RfQjv1TupFOiuE
0NUqxhG6Pi8GV+7mwbEqcXVW587UDhOjDw8mQ2iiNXvYq5Kfc7KWe0lmqFR7
7dTGMZm0Jnyseh8G2vLc7B44z1ZN+psscs4BrbmFDP/wyCrMWXS3Ei1Wg+CR
aCpz9qpE4HTeI5slz3VM3UG4By77q1x4pzk0et/3xr550Q73WLG4F6u/TtVo
RCiZabzfN5eh+h/qIEYTWj6Fb7XsrwHsSt+zAbmdHtpKEgp5CjrDM8Qm9bsy
21ZvbR5bqKAAADYaltPRBCQTrSKBgTqtXF4OSyTPvKIIjk/QBwLv1HJQiGCV
gDM5CbP47KTwb2ueZRmRXL/DjIPfEsOYkHwIEnwvhzTfqk5KWCgxR5cGbNyF
OT2eBSzjh/12Ys3zVZWBMYQ7Pq9Bxq9yRQCnSXt/XopOVxi8gcquIwHcpVEM
BhrqfIt8rQLDxeDeG4KzEepyB+rQ1ieDHn8MRSqjfnubs8zKZOpucPkg/aIn
BCtgOGhLNhtj1YNpH08T8a1COrvSJiEvI8yJovrT1OcflMPn6WqqmorDr5tQ
TPpSdrzkeiT/QELImLIBuyHOGcy53LJZi+aSetI5uAGagkEWtcmck14mbU9o
FO2/tidR9Ssvi2pb9mgSebvLy9OPSFOFp9r6xDJ1ddzIXW0N8+KZREu/5QQ9
dJpPHGY64p7ZieqZixFqt5GlGu/GGznJ6CSHUzyytZo83HwAzKHS/dlcnc52
e6IMdufkID9wffsxtmKgTrOWd6SffSFQmeyz15cqv4K1RKGl8ket5EAbBfUo
/v22GAZsgsii4X0A+vgPzPK3bVUMqSN+2Ji7yodB/7Xutku880HWhC/a3duy
yQv8EdBq7/jDRA19gUVn6sTQEAw2jxzv8y087E5pQFNaDGF3sCcaensrsHVn
XfV7plW55TJnfpb73GJSrcY0eprv39VPuX42EGbkcHZiwK8mfL2ErZd2NYYe
Cq/yEMeTZbA/jLvYkZNBmMkbu1x3kyZZIeIlqXiTP9XlZ6rspDukuROkPSEk
rcYBrdv/czsS69/HrmMbcSoLSGlx7lkmSAMZOvsXMMnw+qlqa784m4Fj62J2
ymYBD6Ng8m3m+cE7rUB+OVOQTiMvCzYxa1MP5jAmQtDr8V+A4nUbJCG1JlUd
TOvLkfvsO+ozhTuvrWQzZ2ribTKdbAkPWRVraspNhr1zc/0EnbCWGYgtVbpR
YP+wtvKKKc1fW2ehgwKD0ZSRUtX5s6SSC/YfkzUdpFY9pQUgN9HelgztuboQ
PewkSmgVLaQ29r31XiEYMCDZMQbC7vWnzSt3balTcExYkvkQcED7TfDGapz3
wRPZqI6wHCQ7025d0IjbJnJhGk389VkZrBnFGqWrgETcmrQVcaFZntiZLn0T
D3UfpJYkTIZVMLzEjUtQdVLNC4G2T3V/iLoD1MvE6lrMfG9FYd3oUVnPiyOn
262Z9Fy7aJSx/yrimCmbROR3s/OkArzUaRDQgnoEqpoE320zlUkxYrpw8JgA
6vcAkXiBYVYnJqgvJrVWF5vE99hTwgtcON9TOaiBf/4GIOyF2SWw+PUBUrDt
Pn6JOPfuzOwichR1iqxa80w8OaYQ12sRqC6ZBvUlwkUMl99XcIxoTYqKdWcH
XqSV4B6gPT+GqqyuU0MH3foYp2QycPneQbnL+qazipzAkN9DFZ5AfLISz8cf
XJwdUqXq+penxlX2bP+mtYDwszBshtVI1Z3X0rW+yI15PZa6gIwwWqDRLfXz
e8RlGiHLeXFtxwp0Vlf5iMwAEXW+EA/xtJwf/Ivdl19uYfHPTnZKv1g5m+O/
iuWrEfZL2VTENN5RlUMUhBiLOpWVb5NZGBxSBAPbqsjKbT320cNkNNycBwfC
yvqP0lnTZ/BvbLvL/3fuBhaY2soy5ZkH9pvS3veJF1oZCk6yoSvX1IN3Yy19
eTloVbDi2lh45RmEJZEeC95SD+TaRmuBjozH7ixW7iRR1hqTCSLnj7TUhfd2
K3zLXGlFlBJtqPC3secGcbZYDkYfWA3if5V9Lxh4Q6FZ6jQnjnJvD5a6nn1W
fUxdI+Xy2iRAidWL/nlMWyec4ZOSdbb/LnCbxhFuzQBIBrG7oxOGBhWJcVFK
DeyUkIvmjcTUgqSEocb6IixCSe4wX4BuY+o7v65hwZ3auteC2TNd3fHJREq+
CRCOgU8878N9p+yjPpwplCLQ9Ny+fe/UtyiWKvpm0EeVjnBBLoynLjeynBoe
IEo+9XefQ+APxkovTRq/lsJgGqDEMkdRVXhduq2AfTygRXva+OgHOYvHxtwM
lsB2zP9FHNJVVbVhdo7j/IHDuZSfO+00hKPs9yC/SA3zMqWi0O1ZsXsdks1f
Rl8JoOgpOK3NGRpFfho+fvyH5CErfwwK8DT1DyfrppSBNi6/jsyXSv+v3M2g
+6jpcNhKxXdfXyYpNUZ88gn4exMaoXc4VUyEPVIY6oaSp3EEyZ4jHjYYoaXn
EfFxoF//Os2mPsbEMfjyqMZXxrNEcfc+OoQmCbpHZb90ocH7npzohq56Ea28
fYyXtCBe1dvdoWn7mgW3ZPgA992f00KT9mkiQMrEbkBBSEfLTCx3Y8wtd96L
yDpp4+SJrvLfHcO+RM9AFdxlQzCgxpJjQ+ZWz6l64m2mmTDtcZAslbkXH1YW
7dVnVlsGxKlxHKrkvYq0Ovvdo7SvU729aFNQ/8PZTYYtY1bdybA4dYdxlUqS
hiEyP663OzTioMTfwQcEqpIKr/Fri20Yzwpcw9rf563gqMGj989dSuaWZ+Y5
GMn/mm5ozAvhdUz8F+Jv9MD8MczssBBb4nJ8FVLV10OT8EAWQ+XyXFexsK44
zvF+aGeCzvKadFPeBDdDMxs4omksKkZZZtxRAO+mf16CfHdL7h9VJd46LDdT
nLmKF+BMNlueAp6Rn8oaUhNmOisG5GmsZWx/ra8W53tp8Vk8riSLNw9ygOPr
oO6AnSL/D2WiYCGo9Q2YhqiJJZjXia3+1H/BbdSU2/nEXDfbA11fH0RxJohO
hIIs+JSpYttTAHQizzBsnFXbUjDx/bsDt0xFJvP3/mrqx9TYwjLhCoQkWzl+
C3D9zJ+JJJG8/RY2Tcb405Nd2PdcQobALcyiGVSXqUaXZii1fRBAorAgzBxO
TniTMJSIMwGdS3bO/pZjnSLLpGZYQ9MDGvZGIoTVth3qT28QR53zdC/OiJM/
7MTqlklzZ/8oA0HGIxyVysmqac1lbqL7azYMyJEGaoq4B5MPluHDf8WudW2A
iBP0228zENyH4GE1Ui6IbJizOyU+Iy19vQwKxYFszkrsGOZUrSjv8BiH6EiG
nsOCxVOy3TcqePNrFGEOdSEALpgRYWgfoRHxa6akzDHn/tQ8FH0mQ/Z38hvt
66vfAhvtqLVWBTe/rWNcHPbPEUyqUp983ga9PgqffNv7YafcGefxIpddNIIx
gsuKoOUvuB0N9G6z9eerMBmvlqaNZp+pSvSg1y9WiBf3BS7z7QTtLs5bHPSZ
h7f+re0paipO/aFt2OISAMy4JyI8kDjRiGRXdbrT4XiZj823il1C4aBm7gLz
SIZn2NZhpFh67He+F6gfCPtgVWWJivF3KP5TyD1WW4w9Uyi4iBdlP1rc1/KN
ZLgu6emEBVAYUfv1WzJimVyHR1sgjgu1DHrb3feaeMYTILOwbHlTSu4yYV8k
ktMnR9GIkGRFANCXs9t0JEAYolXRXf6c9hqxDm9F3ITXqTNhKtbu9pDW5O2T
fJlpr6UvWa8AWWky8CsWKSDyh3N2NBircHF5jvSBzHPIqcp157Dh+pQVcsZl
KY+GFnxb9mQsYDuhtz9iBIeLmfwVTzg5fVircdtDe9FFDjNjUfqE3CcSpsTy
jtx/CzGwC7dNwpTrs8Lgi/gcWC17SNqBx4rBBMYFnVenyXd3I2yu0zD/5o/B
O+j2o/mCoJ/cBhc0kgiVXuOgWBSBmk9hvuecXoaACkvmq5IK1CxfFbtubwxG
tQwXy/cbYauxxwfRSUT85mck9xaoX0Wwi8Dj4FG4VuuLX5E2RjYLHbcLwpIx
96TCbKCVQRKx9bOV7SGbuKB/3eCOx2hz15YXDaNMGMrKBfaMXGgVWkVuCfc6
WQeaXgqdMUFW31HrIHtshPoNjcL/RRsNj/o3BtxDYGeU9gIEQQrtmIuNV868
v1tkC1LTuW8HqffmBIkiUYWdxTdaN2bpVuP1H1jGPt9LKUjhzVFWj+Pg3HOK
R3UjFzPUZZjGtSLv/ioJGcGGrh64n5HtCYTGobb1ptKB40Lf929ZBO35267W
MGXckmV5ZwB/vX/ZWmH+LcPhAB+lWyrNh8Ujb+W/6HKGwGV8k+tm7YdxaXtI
wM245DeygjuEPk5sZGwB4BWMZQtQFWG2gKVSp8v+WZzeDVs7UpKZPVwviFG4
M8+4Rp5lxJVdzHn+ePRoj0MpyED3ejSp80mWATcDMWg633z7mOWQKoiOlV1n
NSunGqRGiPkqsA8B9FJNp60g5GZ+g8+AUgwwCZl7Fr9Pux8O/VpBJaZVDw72
d9R0je7x6aUwsyCDgV8YL6WdQYYaY3h79Q3lhnXvlhGd7YZtqD8pf/Gsq4uq
rR28ImM4ZxDi7YjlcdL1s7vU6BVHFQBXlVdIwyHSMIBnvACAVUcmmiksrak4
fXntUFp5ep3i5mSY9sXiWPG1yOjjCUSiBQoE4wtJTV9Xkx+jYgfLAg/+60I5
uWnBuXByNx62NMb8Hp/qPYyO6+UPVz3V1Is0eTLciS3bPbwkzuaMcLWCoRGg
AEyeqp09YI7J/6KXUVvFeHPfm2nf7GnGlE/C0KyCUVzn6l9jNZROzS+RD+wP
GlfOVTSD2TuMtGwS9/l4h7gYMVGJiIMFqTzLletzVC2sTrG631BBj5RSu6xo
GJqpXFsT5rTOm5014LVhOIoxr7JJro658pBA9PGfwryO63Oz1KsRld6L4Bq0
8i1tSFp5MhtDHeYWS6W1pXk6DIIQdGnirdNJ/kE9KJZW4LYZaj+yKqeuAPgE
vF5/JNGAGsfEL0w3TdIhHb4LKJ2STIGlB/Y3QguvvDhf9snb27FaLQ0hRH+h
OGtWBc41z4pTbHQSndE8r5YwFEh3J9vAi+dy31xbj6sTyx6RkRAHK9+MdzJh
Pnqzff1DJQe5svgQV9GeCl6tRtMap//MpraZB8Kh99IKEqO5FmvCQ+DkNUHf
mVEgm+trp8Ijz9wwdmqEtyLlNawZZD1f5O7m/GuCualzeR6tliLF75stjKJb
j/Isn/K4DS/fpYN5OhC3MZAVmNLYdhyZEzNio70Pvx14LSQKVTZ6O0LVC81D
PSToj6oGqiKR3ASJ6DQ87OW5geGLg9q71JXYK0whJtmzh2tQhrXHB4QmwZns
pHeNJGFbSByibty+WXnrSIDk/cnaazPnmA9XNRTX/1hlcLBYCocMAiIoeY4n
3bS72kBR0cQCVk51oKeEaa8okYFCt06cN8QVz1bfgjyuruzsKKeZ3ab0wMNj
op4nmaibIwVtyGsiPWny6nZw5aUnLtXmbAL4roseuNc8dmwwR5TtEx714QPw
AOm/tNdqEAnOtBf7FaT2/I4jgNPyo8kjCGAWU8b3BZOXam++oofnpuLm5Yq5
EYJ+ck4a0gSoSk7GmdcjBMoHdsqIBssF56ciQQ8DkEEFiqGhIl8m8Fd2kKQE
LU8h6TO0D14cqhsjaNUXxDIX3MR71IPxTgFY1WZFlBgmHwGtlE4eEkfbs7qW
B9hB1XgenVNbeHt2PKZTIuWRwa7rohQkIlemBF0gj5x+S0OUL5eTreiGwafU
pdKwO4+9XWMrh89TW4zgKUL5P1Lqlj/dNZL/lJtWuAMuHdMuXimLYFVY8/Aj
kBIBCoH7KwyONjn6g7kPGUORND1ZMFvHlR/9jnXrdoRg9AKYhhFEkyYVmxeH
xq85bF3LfTrO0gIveVb8NlV+NLvPalvJI+hM2coEdmngJhYJlQXxZgHC22Sg
Lp2QAgE+KJvKL0KD91nMtEmP5k6np7l9HI12xdBayMV9ISAr77Z+B5AI1LY/
gyUqHXvwSn5nQ8PcmbOsZCmLe9v0QTPUkrA7RSv6kdevDOioL6eUWjjvY6Qj
Gm/CFuTz939ktKnzUsVbHAqTlQQSz3yAA6jbJRzO6LXtkhfWABulsaynaJlr
J8A5y/Rp16zdQC2rqVDywqOK+RdL0bgeBZ69ymKivH9ZWd3RhYP7+HAKopVr
WqlrOJB2l9sTI+5S761EOmoOqNjQoYSCM2Op6N0Fx6Idobb2f+h1Mf7CIa1i
SCIgMM4W+S3jQI7z+7qrY7di+PcFNFhE58JWUvHO0OHPsGBlkgvTM15wDSUg
iC9p8941BPz6b3l0kfuaqGWvfglr9GkSVemXkWaZ/+0FSL9Xgp/CeUqXB7OT
R7h2ngzys3g1y/NKo9w95TaMCL1+wdnuHkWqB/N4+bFmGi3RyZzK5KmqVqpN
V+TbWxkzEUBAEXFxsTI1FOfvIa7xVYUklACTfuS3r2XGIbpC04PTXbF1sP3w
74v3HcZXeu4VGnjCWdg4a8nWBlOLM6RqIzJhzA6KYeEVwf0mBtIVr4gtdHK6
HwG/t3B0iyt6TzdiVq7G4CmJlDb7pUzqzHm1WPKKZvfN5hkben78vRvXj/ox
RE4Ta0vVHurbZ6qPFtbw9YSxg+1ncsm5gBaojbAngP3AWqDSNlv8WNv+VsvH
a+CFy9rr+LOPskpf/BqFRBlxn43Y7zmlbemWQ6mmt5vwg4MhZokFuMhCHZNB
1T7T2Zh1nZOJPfr5fiyegb1qovDfABQyUr3j4Yib98zx9GnFYJlUojCum/RY
nZxYvKNe/Hpjh+C9ezh5lwdNmKkaGkuZ8sdC9U3q1NvzI2ZP4KDVmUxPU6pd
fDdpcAt4foqhysIVafsKZT3WzsQxlkQ6smoU06fifrzPT8XuEViA2KNZsKtb
81D5ycSzmhdYxGwNHlbjnDXQrrLoDyXs910h4wqtuGIYlsumvBQE3tuc7zU/
4sdny0QqGZtHplwK/uPry/QIeDMgr44+S8+rtB17UnydW8VPMfBxaE616oev
8ugmjj/cWabmCspGGNnhd0Cxa15/c6aE58BA9sWvSKZT3qewM89ZU55JmOUq
legf1MgNS45Mi/vjxNPac5MoTdZUdDgrXmbNqfFLbg35NH7/ez6PY0oZ4JaN
2nzLRVeL0I6yXCD5d2qkZefQVsaF+DnPmNzOOVI8ku8odOwWG1H5G7zynS33
KFFLd6dya41QAruReeD9yJjnYC6eQK86Ll+1kt6ZnxZIXzQ3pbXli7XoaXDT
6IEPhbS53dGofFEziTYUq5sLEz7gwfnZiXaBYPsTSXqExYaiH7m0tk3/imD5
LOcO0IBtRnLI6CcAfhH1cicOdl3Gx3PiMYjm5PhLw+9px0X3uUa8ACmGa+x+
wUtmGNF0fLm3gGp+t1FH+hVXceGvKXOmswoLZQH0E1/Jg2QYbP1WZ+DUeBeR
NxuZcNK2m7MHIniTsAC6PgkuSpMM0ogtDPwVbVppXoOWLroRSeeSnIFMDWy6
5q3HamopauyviJ6NH0lI4Y5RoUz+wmIXhJ8cFdIxjKsW2R5gkIpNtrCWTL6m
+okNg5xbnvvdnanw/UVjD8uRvkeENga8BAphRku00lpX1DujNsrLkCSnNM2C
zznm3gQG+J0diho1Bpy+1MBo+i98OKZkyIgsr2Doo4vrLkdbJ7cMSzyl4O68
iVamO7TzcSuCmG3uAk1p3D1sApFiZ8P7cw6xUtY4DPPg/Zworxaf4RNm/AGO
pnA+zZajvM9cKCPlmPQXojSfP93nC8PwnEL3MaNimAK/AnXX0+B2lZYvFPzz
ieIVGGh3LQRbHquM5uu0eII774v7yNafkl7o2TbDcvVhRm8Z22Y3SEk6IP4j
ZOftTeDUMsdonYzRfAxXdxr7qAcV+Qm9rst0ANyD+SXGElRAwMu0RzdKxEvg
2J6vHOs96dDzC3D4FG71UUWWKLfMyDcPvglmwYDA681lH1bo9fGOubvTz5UK
pL6/ok5kDsPgNPO9OL5fCE4rHpx7Em8c62qmYh9KzqTKMyLrZ4S4R64P2dBY
YpbeIeEL2v9XeDnC+pDusq58RxEjTgBZn3gFvWJsYLc2sq8xs4TWC3H6sM8i
oUr26Vbsy/OUfMQAHO74tf6xm46oUm33zhG475JM+FbnNX23edAE/13TW3Ha
hWg3r2EtM9Dq9t8ak18tPLBIwWAt41JwX0ABL6M/1RwYxXUHTUWxd706suz4
EYJMDJUNnAPv4f8Fn6o6OVmVFQqilE3tu1XZzAL9Lpmrp08KfyIusNAzmStJ
c4+et+gZGHAhNfdPwViwBGtVBNJcEfyGWE2o1dGD1PcWNuY9+IAXjYVo2+IL
glGeLMP+I/FCLJgvkOF8xph0F+kpXzGqoZ7F8f+0wHIfmwtw59NcmGZF1ZX3
K8kRJZNmVWRpv0eYShMtSWhLC0tJNJ67DV7jyqxW6ifQ1wJaOQzMeu6eqqxM
Xm7Dxmbyn1kHo1wNen1SLNhMleFYWDDyermfIG9Y0xwXQGvXAXe+F5NqodqI
7qrQdLTJSarZ3UQd1fpRr2Vcn4x2I48rYDuFpXJKJ86oqj5hFHg5mWoKRN6n
vbRjXjLQLDNYTajn6RHciQYdNQaeyEu7WVedLqtU0419c3klhbigV14KKGTm
H4lQGuGI72iO1HK4xNnXP/I85R59/+cDBnPMcw6cqOGOckIrmPHGQUyxel2L
q9dQ7T+LG8eZN/XOkCSU10SH2zwnBQtjdCbj+IsuptRdl85levXleuEa/nRX
N8KhvyVi/uIKxu3W620wa6THBG0P3qcXxz1vD+8XVAwScJoQaWlYhdTDhDvD
DqPriL1Uf1L2qfOr/eayCX90P1Cc4Zp9sErgVrfaL41tkm6rCM1a9pE9woyl
m/OfSnymvd9XKma9w7hAPCvJnIy7QdXXkaKl8e8VYBNR9EJyhJPBLh2LTVKq
8lOdaWguebdHf1obCuDntfxXXJwS672IaYBgg1vooET/UH04jpn2Fhav/ex4
7pJTzVZstOCqr0L2/+Mj2xdB+fLUk0IWAuu93v2HuI9foR+a6qwnmgyL/gcd
mZz5hp22A+j5wSDg/s9veJyJNfm9gaa3MJb0cdBQuhsweY/ESfPBx32oSoIc
sDRxT7L5ttEiGLmyouLxAXHMMAc0YCm4kHS5Is3A8zVgVKQ8KeP0cQCxZl2F
K5gSuaT7LXHwmYL+YFPUrqfWqdz9gw7G0m9Jdf/HYPFjLyrlyh8Sq3JvvOfI
GqBXkF7YHl1a3k9OhZZtR7wvdjGq7li9+ohKRhg8TnfqUN+uVjjuGPRdzUtZ
Zr080iG7v4RiYnYy1888n3E50uK7yHqT6n5SaQObaaRzDHMQrEGneco4L5xV
ycS7lcDnXDPemCIdOy/t5SRxOP36ne2xGLpuxWMM0EWsY/k0vlS0Z8tGdzA7
yKqE67TFRO+anRXR/NIsPoVGyCIzvBKw/OAObTv77jGPEccqwcQELgzsSG0y
L03d5yRYB6nX4zZGvIjbKmfQiOxisi53P4q9Wby4kPqjZMv0hcTPM6JzF2k1
U33K2c2nMTY6DD5rMcJVFbUSdp9fl+hBLrfAahb/aQ9RHietLMDq5sEXexuB
aMRiNLExW+yddszt95kL11EOvyw3hri6bNyZkIs9trCuvTbJ0EPF7hbjOtcF
dX2IxJlFWKJ/qJb0YbDWAt3yXxUcf42hT90ZCjR2XEh4MzPtR95+tz1fekJ1
uIzDZLxDAuA2m5hsVn4DWfFL1EV5Wq3EXAkXdbm793f/31xl+FmPCud45w8N
67jDKUECOq6OpQHhBkf4UfCJ3d9ln+ngF47Twe3s39/ncBJy8iZxmTSN7rFp
RITX8NtTLFlfGODMpDg/0/N8IknCP90eXc5HOTJQ+eSznpZt1whfh5c6pajp
h7kWrK4mcOBOSmX8+NHSWHeSRwgGzYQwidE+XxEFY8MrfMrEr5iJ5/BdRy2h
3Q3SzIamyvVKWSjcxcc6E6qkcbgS0T/vT490Tj/7b9lZDabnTDYdnoS5reoI
3j5yIRSCpX41vcazknnn1ip6msZv5bcNFDtjWuHDyDkqZU2sMuuxqprE3x2v
5vJW0qwmbjXOr2j/YMJ5R01dVwZGEKquueQR10JCHXMoR0vS/qpg1GfTR0p0
V9xujSjJjeRMmLZubTcPgSFWme+3Lm641RoQFvyGYnHlUkanWveavbmVddDL
SMA4fbqxIeUUy5QDGrkG2ARY7C3hndYeG9bapKemNuQl1rPHeLM+nurvLJTz
tru57k6tduabDGXfDmm6M7UQcM+82i1fntpIQoeP/zaXcZDChLLRS4Net9qD
qBuRsM5x1W16/jZcLzyUSSIgRz0hxeljYCbZL5DT3YcmBaCKF+13Zeb1FuAA
aau7xfdRIaCBFmmAApSrYkqmhgQrwwNQtQrVi3SFjvFX74kAx+XaFCmsq2ZA
gnTcpBx9xNdIK490xhxayH8cz/xnDPlk/j0A1nODv61sBORzhOQRm4WrDS20
D9rFdsgrSjv1hkMP2nxpgIdjt80GEIgbo5Dxv67Z6vB8FhRgPJDM1984gZkH
1dnSeGRZ5cCRn6/wl7tgNVXGlJxwj89/UVxgJ9dl1MGQAKRSunjUyCeVu9Gp
fQVN0xzU+dfRrbfcMBXC//Uz3qVBPTV5l/0eSHHfXGyvyJhows2AunL2mWlX
QzaPXzNwbd4+ECk/iqjYSaPwbQKI+AWywQrb+UNeLKtaS1xc4u3VhHRwIpKV
aabBTIhvfhXy01DDELs8+kXHgPMP16os/vxRVqjZhgDBGGXT0ixGO+dyzFqM
GZCHWgCwHmnIEN5ySrdQZSRwB3988UIrhgcUInwz/yLWUJGlD8EV9XmwRtrP
MU0RVcVpRviL3LhGb0Yef64a6oa2Atg/59oMKA1wmsVfIYjgDW0BaLQuXki0
pLTkFGANqfhfM/oHl4ayTV65AyIX0Q6IBs+GSCZj+WK7q1nevCUt9cHFA7Kn
M06Eu5VAB4DzkXQag8gYT3Xn9rBQ/MNeX/OmJmkdJs9WsGN84iO0OXjX+Wgv
T5xdtAIpfqhpA8M2Pj9B0Ofr9ky1SXSwWFQzFVehMqI1JCjBqoSXuw04JwvY
qHlhVrb6G+sIPMYf6J1QbSLRv+jU28tYwT/xsZxlDa/kR/zn1fP+KmTY9/0S
NrUiMXPkyTDcN7+tTa4Iv2vHsjzE4ITXPDsVmah8FXvTIgGdqefHrKRo47Dj
RP/vN/RQXFFUw0SmJwPSdOw2DYClubQZ4MpwOR9ThNEUHAIrb43mN0U3g0uh
F1Gd98ARFRZcpNe28TRiPfKpNoD+pV8kamEbOvGTmdwtxIlJ58nMg2viZHbf
T0vn6m31JFraOtuqsV/cTUMeUiBTawatB3sGKy/KZULHIGXmP7ZtiqlJEo1u
qe/JZg4fwtxy/JCkbQ6UHMR0UuCAN7mcx66oehMYU9O/QFzoloOE+gdybPbG
3BJ5KhGtLhsfeM07IYdJJwWpV1XA6xlQgBB9fiwqTVmEvIvXd5H9q9ss9kUV
0BvXPgWsXgaUjXCvotQpNG3feFKMdHilxWl4JZJp0lQJoX7rd6ZaSHQGT3pQ
ql3Jsr3eA7bVayloQXlGC0yGl4j6mzzT/nsiAogb49SD2P2tHzanxGKgLkCp
m8zb7aDwc+OSdcKeyrU/clk10HlDbjUiNYkwIHI4B/EqL7rawRPEeEFadsgz
dPRAqlJ2/5/JX3kbfR0jKm9rf/YCeE5czplUeImZd4DxMROBHsby7uAYnVHZ
v61GhVwCJnbw0O9s0lobrkTYaipaSnD2NsTgYvo+LlKExzNcLc2STow62C4X
jZZQEOZrebiIAY1/tLuvK7ULlCfNQUAELcXRK/gDdnt0mhm7t1tmsGT8K5kq
7V/KOuxGntOC46ulY6HIQxhaLrkj7XKJc3n9XEC5+bJf60F8XusmoEIk6g6X
cVvyRS78m6IaLlP7GMcZkqN81MQLIoBtenB4a3iHhH4oA+Sp7C4Z9XeD4CaW
CJ3aO3BEfBfYsNLLIOI5goXkW7zvOX87R9ZzoSL+XDoKm7wJFyrxuSxHs5sd
nfg6LfCIE2+XFBKrte6TbNouYux2lB1asRImzFHSAE24UklC3iff/BxNKP0Y
rBReoGUgY7Mhkz6HVrmZO31U5de3JPR978vomDuvF0QyS16fhIbxfD+fmg9Z
Ks5Oct4eicg4lHa1/bNhnvP3MVFsER4E0kQx3pBhl40u141W7jvQhE8crRya
kMnCJPPY09E4h4lTKDVnDf1/NRh+woGc03JOM+rmGKli/No72DSja2ZZMl4n
662hMTmGUye3R5i1NNZkRZ3appruoHo33A/ROvhC9iB4zPlWlriupsTRA4BT
/U8Q03ikN5K6UM8WBuA2suR0uqHCtwScra+GisJ95pYDZxtWnrsRQ+eVzeCd
wtmcg5p8qkzbN/lwh27CH/J+JJSTsauEEVQ3v7TI1fLGWPaQTLjP4YOyLfNx
CT3cfXxcamL4joObklM5JmYfze0zMNU5MXc9ET1qnxlvU44WsD46Vfy/UU2p
P73ZKTHK6MCp1RKRKNcU6LQZmtBzwitpbWvc/YY9zDGBcoLCEVCJ/onGqFvH
Adp0BRAWUZCoQBaIqEPvFjB7O2z9ao1hI5pdNdeCtEdI4EAGKIvtLvU6I4NN
23+1CTAo/X3wpohybQ8rq86uHsesye8cFTtfiX0TOHbE2rop6eAvE4tCx3P4
nVMpKXXYfBLrNEhbzmm+pAAA7u3kWwkzE6FfqpnWoYRnof3tf6iENLj7QXnS
rbBVm/pMN//aBkWvu6SztD9kOZnEMihtEm9c5iJ4JFniurn6iqODeeXp1pg3
qCHmiCPipJBKxBgVwrI7kRKOKWYxBeRKbfnZ+j3k66KGMvt72rC9irvTjyH8
Chvlcz9z2Bgv4Rrfu1inKK8rqswfboVgKTpIiUgGJhqYzU5HMlS+xOV5SmpJ
5PnwQtP4MLZRD8inDmVVEvZHl8ooHC8mzMh51/C3oerWSrpE31y7mHWJgD22
2LiYzLqoSc5It7fOLigKDZcv2Ii/DmGF7duCPiKFRE9mHQEPDAhG6gKkl7t/
DdE9At/BsJ12BQmDcNfStiyiMNdeHd2onwRgzi/BXo+g8bhxmIJ+p1ytgG5y
vnYMxbGwqyUyDobJj7oJtirfJ7eAWWKP+PelrLp+58SyIhOlioqheXF2W59d
4X0EZjCSzrSmUvuHki1abQXy63+YG5YFHX9nPc8rin2bZAOjDn6xC3THXTGN
kXFZAMCS52O4NbBGz7LOVnaIHmibCvmOAQM/RA7W3Gvq+Cw2cQkWgMyO02GE
8eVfD7nF7fBf3SXtcfWcqEskyCSaIw25bBi8YicujgfCm07YH2xxanlqAWif
7752Z6Q0q7B+P3j9giipWaQ8TIQaBO771UPEB3FZTvFKAzdQvK8GrLfGg+Bq
lye4cK5U6Rwox/E55bkMiF3wRDGT/O2FW12rOfTwLETJcbfHpDjckb8W9S5K
WFU2vNcgCktdBD7glI+klY9IIBfVssHg9ncpRTyUG+gxI77JJoTaU5K6lVu2
WKegn4LF8WggEXeQS/nQIiFe8Mm7FQt5IMML1hE72/HlAgXo3hYj3QZJTf7d
HOcYfBTIIOYhwiOQGOr78l7OhuFCCAlli4IYYhiGEjN6EHmibzD44JMz7KJj
88UmjsBFJd8ZvcQnp2PUlVPZPiBlFiMC3teAhtkFG3m7CuvD1YOeXdX6L06b
TnSIaK0fT9m8dR8RCKvAQB/069OZh1Z1l8dLlarIT5FLcmY8SiX2f+rlsWoQ
ObSWF+4HP23wy6uOFtLUV/lWGP/jU98VJOKz8jbeNxr8RP2dAG13KzQH9dVy
RyaPWMkj8var0uAG87M0ZDAjEGyiuqpBGvby2X0DNI+yMSQLkNhEqG1gzVuN
eR3VOBH0T0HGErXJSTkYhQB4AML3Fob2bNKf5gsiYtBhzzvipC/ct3AWO+lX
oxKRO6EobGo6ZtYK34BXjzfnw+Ep/8/RSv0y9TPekFv+LbcPPmBYCsLDmHAK
uhHb40E+HQbGm+0SJyk56hyWZsozr8x6put5VdLPjRkDq9lRR1XMgMc8jmmk
PpMiZ8CcBGdtFxu7QvE8svcv4ScclATZKbHSIqd//QU+R+RrQKRGutrm+kRW
6Nx7NQmU221ggDJpLz+oTz3e5Bn+9dDPlEXzvYd4i6tBAPlYGuUNBo91w3Ni
ULiJSu51ryxAX7fDKJUovJspOcWVOmctv9kQqSz3k8lJT7ZOx2P3YCY80bSH
ROOwrxabA4u9d32Sp+ufYIPtMazZevurvabu5eCO34GCnwenLGcGEygHmqdX
bjc9+pJqv8FVzApeU4rTuGx61G62PDE6E5NgywOZEUMhBQurieJueoJ0KX0D
c6MzQ5Tojbg7oXMtK0zunSSYll37wNkfcULtccE5/kG0MgPAmJyUbZCgmmNA
ngeYQxmEAVTloXyb5LKZH9iC5Scy3AaDb80iB8EnTrN3wRNOfT74UCQY9bL0
iTrhkDjfSDsVwSZHxDrYfpnzKaSpaD6pG9ARBn0PT8aPs9tOmR16ZxNuctox
Y8sBmTcuKuCAf2i3PBEvNXu9ho1PdxVq2Xwqi40/omtKhSjVQQ+u7gUl00PP
b/bZQBsqQfa+GZdBgnqBNQ7R9Xx24Y6oiZTrdBE9fOs5AvAiGa4b2y4qRctd
rToKzZhDFaN8TOAMegZ2aSw46gvMIj2EwPRwwymYr4f51uy433D41PMYf75t
i1DSjBPbtssB/Qw0mKinWmbjgsJ5bANlPOMF59w9cAIplSnzQrSvq7PBqaUo
YB8Q1JVxtOLq+JvbiltweA6myO9k02ZgCVmnTLOdJmFNquKXMde940To0t6R
w/ve3qCsIjwij2hEzCTPe26HCsMlMGUhFSVQmsRw5hi8hL6xE4/9jtdrg4yw
6EGUGCgjzUBlcQs4uhZxTIYMMBul1KRIO9VNt0THpLlQiXaFBSNjp2EsTfob
8mSjdEvZjky63/uZSvXwmyn1iEnDGYm+IfksL502GR6dVVHLIfYeaHPCRO4G
nOkWd1aYx5kgWUnHDjCFwovxrXZjTl/2Vk1E+1a3dkSspBTEOfz3iNVTS8cM
bdtWTvGM0zAWQlTwPayuQaos0mYMLzrwjsaHedtm1QT1ZxbkxEdanqVxHIxW
b2f2sN9fCE0NR2DI+43ibigwshdSFhE8JWExx6ptLdUlDpUWqJXZUDIPg72b
AH82T370O3mM5/ivYNabXLSzYbJTAeyT6RzvfwLnDEg1hFacWlZq31a+1KKl
1kXrCxBJ7EjJuC/uaePA4FzxHozpbsRjN6ni6s8xoYndQu1ANH+Gm8vbND79
geGZQAqBm7YD069fT+/EeZIWE3ZZrwl7/7jSUJ2RN60i6odLsXobWBe3b/Uf
5/1ovcN6+WbONuGDoBRZYbQiNVganJ1iu/ELmC6Mi5gsHvLyX4C82iaAlGuT
LelfqJ7coFmtlzxL51mey4QB6/A77wCx5NJd5Euq5sL9U0uQh7Yy3OGTUoDd
X5DNn0m3YGbfE8xOkE6l21P1h5ZIKuaDJu+BsjfUsm+9LtDBFmt03FK2FEz0
IOQL2eoIULgFuhdwaGZD8tO3Y+8WVwC9/o7yXXilySzmvriuJrgYOqhZrzOQ
H/o9wSoxVgcFlHa4eijzjlrcMuRTnJmvVPC2Xs6uuTLUwfja4cankp2VPXJv
5Hd+/qJS/e6IYsMZ4e6siqEdotxamattaJHFJ9QKPd4AtpU/Ihsm/TO+WWwm
mOVHEKWPkjNhgJ+SbwOh68imzw+TDBloVapNXA118/PfX4TonEZPoQ+R7Vil
2NYClqqPQwz5Cjy0HNEhxeDhE9j1mwB63wQfdkJpuGSgkUWBH8sNW2Jvhe55
wBoiN5rk9CfpCdusyQ2uHTE5x3meWGrI06p4LCQQWVVfQxqIen3vVvxpFo61
g/bjwvS9Gyo+KWI/s8AKIlC5uEh+xpqbf+OaKN0uMnSC4Y4VWq3kvqHzAI9+
/As2uUEoUE+bzDoBefviYXEct9dfcVcJ9gYj0dh9s5k1bXGu7T7/JQZdGOZ0
aHL9ue5etrdJTeyIpptAYA3K+0ZhxGM/5Eq0IDqKViQyXffJFicdV62rkmYo
MRQH8TvR4MDWHSYWbXhaupIPo7q/698s6gCw4bQKHvATwe/SNL6nRpxYeEBc
8aB395iJqzSM6Nw5/d59RbS45FU5MuVZb6dEBUPk57yCOEo9NIZtGx87IKKL
Nulav4iBQ1dMCEzjbLxtMtBqzVtIcyoo7nOp96NyNGFPUy1muqSMjJsmIfGF
9eTR9s6u2DTvObQu0D+c2uCiniiF+oD/gHjVJlpakmgrDIAPtLdMGYCX0tU9
HSjFIcXFW5m1qrP9K5yBnbisH/RY4ItVfWmi/nI+RNRr6Bwdfz6thnfxG3NR
pDJiJ4iBsPo7UqB5GglDcxXoMBPesKcpS1czUeCPDtE6k5uoeRl1yseDZAWC
r/VJ2p+F2vdsdMqIOe2T6Y5/UzQxRFpKM8fPETIMuywNpH541+wVnOaYX3yw
nrg9MFUV4qlvD4DEnFTBnfQlpXHspq6PzBTIfSiL9u4trOG+gvRfj6TGuqDL
ON0oO0+TeZfR5ycOnp1LIZqQmgXi5WXCx6kIn1K3F0go4G4WPovqxgfZU3O5
fzVe7bWi61zDbfVB0Twenz3vg7t6HlhIwvqmD4Q0TyhGK8VyjieH251+Ljv/
lpj3pIpOpcw6ZLP64DyeryeC6Ov/JBAFh8al8nmyQXjsX9pUNA6ni3QdLh2l
YHjoZ1F01Wi89stv7APbThza/k0Z+d+b+UVz18+o9/Oa+GtYVntw17mgTNqc
vVa0RTYGPXaLk0eO68gLd2jdk7CahQtXPXbBK5GV8SOLJ0fK7U2S5vN4WKtD
IwaKKr2/Y4Rrs5w8jfBwWclIEhTukKPm5f8dBxoicYnn4BsVtDjYCJsXlg/Y
86cDJ2KTqzsmLIJ31i0KWR7zx1BrP6zkBkfwVeqGgAuedmh0i9ijcdBAKf9x
E71oniwEeKI4FjXw8KfR7jAANtqxSUHmTWzd2prCuOqSc+wIts/vUFxXwJls
cD1qni8sObt5TBsytMNAF0nKTcJqo5gsFxoKx+kGLK0LBFJO1QZjnznSBedt
LDichCCuLXra9dfP5VtZP6pqNOUhSHyYmBMc6FOEJxrpOpI6SFIYJgB6gkJw
IRsZyOdoBAJJWSl6KYSz4tbR9zh5sjtJcXgCaPZCRAbyUZVYcVxP+PxQYvJl
AsZ4qMqCsVz5TaU4V1w4zbeYi7FUm8ZARQhCHIv3Zs51tZ2YDIed00RB0LYX
lN1KH6elfhVTbHEoKgpFXrXqLnld0jlTHiLu7fMgTTXVdXjFxtS3dqt/SEVc
ha6yo57joSF0spOzch6Wd2dFEzFptziHlwnFaRGLNjlXtIz2/xvOGuZ5ck8v
oxkghS9AEv+96cO7RUmm1VaWGomWTJdBATe50kDpUZTVuEwgkOGrwvJpKbWF
OWuNQ06hAuLcRW/LnkfXwxrCOJrpcPVjR7RXgGBCtbtmW+Uj0eyMZ3wL7uPB
sdrDeEC2LG9pID9Ii1HZFBbO8xFTPDbosd1AwmwfvKx5OpQrCmLQOqGlzhov
ah0HSDgdDfVWY4ChFH/iWf1Cj/o/sF901P97jESqOVLFA0H/HA6se1RQWdAZ
6UvjbUlJHQLnrzIRFEPUAx5F6z3+76wNcKSAqksuRrYW8IOA/U0yUNqLVOR2
Px5Fn+SiWjx6PCYzD9xviKHFaU11izhUJ/rm5Oh/dPJ+rJkEYthSCDPamWLF
h47vUrtDiB12rxGc1hrXVMb5EP0FvEUgW1M2sQT3rcHMDhOtYVRIti4rej5Y
cvUnWMlSREZDTz266WokisnubbX2g0QYLBq02XuaCHpd+B4wRuPIqpL2tp11
vMpSNmIYeiyC99FeRz8HVK48zPQOs75x2zAseg6GOHDumKC88sJKSXH5ayrJ
c+K38vYwFH3B18mo1sWnCX3ZtYPwK+mw5MnrI7jrDcABHPfNd9X3KUYHGGUL
/fxZQdeOfL1UYwKPxn0dewmv8ZX9Ygj+1k+NY2FP9Q+x2uyeZyG7E05lc85r
kU0Sb2pAwB5XN8s89lRDWI8PzdiQymFXmfw8Lqg8RNwjW9hSLn1EGw0Qun9I
URyF0/DT3sOD4bqM2eFsU2g3XdSoY5ezI456ALmpho10jtqFRq4xgn2Y6PY3
sYGrMhH/JW+J7GwOQlPARezoyg5ppTvhzzBJILZjunpkBS8dapFADyzYP0qX
u4uskilxtIMUDFjrLJpaUc8PsCo6uj7u5JTmjcnUrJ7xDSna/yfoJ7Ldo2Jm
B3WxBztVmjuQQlI6tw2Vn4IcetDmZOgzd5QJsy1XCeFCcjE55IbEeoocbRmw
6pT59L3pprguj6YZLplGqHBhpps4+JcFVo95om9QoK1EAOzKvP6kqtwV8Ck2
AJ3q+HT9xcRw/xQ+9wSmRwfz0wL1mS8HbxOygMqg+AcM0moPeSYILZiKn3FA
URAkiyDWAs4uS3k54IStvDeQ0cJfypNS/BNlYlVMYH0nnoHtRvbjSd4Z/u1K
4wyjlEDV0I/g5sCBaGMvsSPufLBxtCN6caifaIfSYJXHZBnQJrTcoUWULxOx
Aqe/jsvDPKD7IKePePK40dqGqO41W+taKIDvLhJ5yn9Xrp44EmzxE1xo3qp8
7FVHaJ4VdADX6kvAEI93i5BebgOMSRKG66GzbdUPCcrKYCSd+TQDaqwfVLir
F18ANULwgp93ueS6dxXY5MNFAffv1MxvnohERAau1dHdDK9yn0ZglqRIeI1v
BIt4TcX3/VohBR4lH31LZPPzrhzfu7iIgDxu10k8OIJL304bJ/kp6gUw+sgS
j3686DqjPUNwpm/IsXLa7mIMr8u2uEbaP03EgZAbPw3D/UzRr8CYVKv6gmE+
25yy9Cldd/PyiXKwM8WA0BOw4yFKQ1be9x0szwXdRpTLaPy9a3vyNYH3e0Vk
aDT1IFGTfPSO+u9fOWbNhicqQSivZIG8r/ir5WNbLp3IrRf/Z1gPw2Is4z5u
plbhd4t6zFP84c/CnbfZtQn4ScPVRr4EBzlqyTuk6MeKdWLS2L5HPREZjTHQ
YMLSpyNMi7e89vVtvaz8s8Il3XfKcgwJi3wIljB5gLpOM63fMPM7SqOl19S7
4fLIa/Gv4ol+2HpJszr2JL82VEdS1gH0hVfqs2saNrZK5++j+R7UICombsSf
j5gpuLawJS0mHkkHX/V+WpdDYTJgDTV/JR0CpFK5ZFpjp+x8yvld8Tr8t9pF
6vU1Ki+xLoBQb2/Wx3v2QeN1KTAZazIOulpT4Sy+CTY+VkG1kck0bZJKFNIS
QYrUkdXiwi1sxdCa6WvqQsT5wA+JlaDdV6ky301bvd527DgbJSJYBcpsdCmY
SnG58kl7qDjO4PBdgSlqZUUugWhMrQHHTT59hSIdYs5togqCXnPxOFLhDEQE
pMc4xTDzSd5WtI9gloevkjT2rkZslCBbmjsQD5hhv3kkYzj1ZTVTrqN6hE/0
iIqqXVNONgAGHjWLUaO3zt7tE2sFdOaJv+ESt88e4HY6iOEREqVSOrzTyhK/
epHIIRQmheMMUp+6jGVTW2capjU3nA2/bPA7DaXv22seOvzRxne4LUCIfCmJ
j1n0zjazJlLCLIKvnGX3mYuYLJcoVkuRKWLx8NZ8JPtZtwWB4+cR0ZIWHjnX
HWsGz/nl4H7AKiaAwbU4Q5EoIlqQyXCG2xDGlPPkHix/I8tNEEZPNLrkz4yK
Fd6svuiyYerPY1Mqx+CE6jqr+sWo1X/CR915Ij3zZ87F3JCFAoZSDjTiZ4YX
b2sCyNtPrjqEWNXCLAVa7oHOchlwQkW6dQhrsShWs43UaL6SPKWq4CfkMUI8
Dy7pYvX+m6JISljPDWrBZLMfV9YSN2BL+Uo7mXhIzOkq21u4ozbB42sm64Ii
R9ZDIsDL0heefI1TWmuSp5WoHY5OwC5dR5PGRFaXUOPPuAHKMLEi/vhiHzim
POMr0tR7m0qI3UPXBDBvrVcyTPYd49KM65eagm1KeAwigL3fLnXAGHa6acXr
O5/SgoJ9FSxhBa9yy2yXzkLIYpfTiM/EYjlmwr91wrWr+UapfMi0fwQz5OqM
BBWoCUJyCZcltklsMjc0HAhCPyq5n5kCaltdTiEe9lu4WaioSv+IbARRXH5w
eEnGYFnXPY0XwMtrkBXxwXWaCSBkg11ev2dWkpV6zKNafxIt4P2ICis69fL+
Sj2cmXjEnE2h0Bjef8WkBTjAvulEsvf/u8qml2sBKdZy2GHYa0pc3bMYw9Zk
lBrE4EDTpvOgPMN6B6b9iCs1TyvIqautOT2a2IGiMrEylx0zK7Ep6n7JCfFP
5dbQccQEgIyfEa0OI+hb6bVDtdTZ3A+M6VQ2S3P8EGcJgWRkfsRQs0DtNtTt
SgWzi/G9qD+MARQrcoGfXZgszuiP3lDDgSya16rjPF2W8Yv70B3aO/XUgeMn
gHULmyQ6DqXWE5AfjRbfzTQcXyTh+Enu4z8xON8vnC31qeGSpT7JCZozJ2RD
2U/tjRpQ3K1xkO6muvur1UgRlTYDUV6JxVvX+9yUxMtJbWmZrYXz1XhapD9c
nqxQGpPcCVZ/sQmUgnkPoI7RYuGy5SzUJ143xs1fTqE9V4KSOS2TKWVieBAL
yqKAlydYSvgsOB/FsdTFJxSAujK7fVm+rfIJBQTcZuMWEwrAWEYUVuQRRif3
YUyiv2bLl0AjjPTtg4kz463bvfQzR4VJ6I9QYAdc/peKMkBwz28oiSBf1IBD
/6xKE6UDUwOaQrCrbHZBf9OnpTCqRf9q44fAYRmpGJIsORNkfK0+Lw8vRI+V
MEjHL0L/vRr6WtzzgcZUIifOt7tkGNxb6tJfF7vV/XdBbLyP5QL9M+7+v8lb
Liywnyk9XrvzYmLtZGNuBJLfCOCix4I8LdmVASy9Z+quolzbP7LOb4yVEL7H
YM9WbyEUdhyjPHSD1Wr224v4ZGh7Bec9yTnZG439cyMpq0Aj4hKF7ZgTntE5
bECgDNOxp7STP7V5cxw5bCqXwpkrUQUextQg6gn+CUVCPKPDsHHtNtVyI6/I
d9HaEUEYGg5VY9b7ypiN2ssjgoe78Aqxb4z/w++c6zVHp3xI0Mmy9929+bJ0
dI490ixXnThH9fRiR0lq5AtGrBUNQsYYvqcLEjiWfeVElawPUDhG7s8dMOlN
BSQmGsi70K5PKxTkmuZ5eJpERWKAlknRLnaVWIipfk37u39QLDRxVx8G3Oyz
ywjKYIEXhusIxCJ3Xq9G2C56UDOwkoMwD6i9FknfYPDauL+TnEF+MpbJypcK
1NC/TuUfMqyuzPkegSYaVM/FJsUOz0N0/dftuUE3fOB9c0mlnutcn3aKk+or
D9r6bAOEo7ukQ9UJKXPmghPgy0o8QztOOZsDidrAE8wySh9yv2rJWkswWJY1
WjTSerjTm3VhcN8vEf/VwA0vUEHrw4MxRm9jNUEQWHAjpzu4/zXRR+O0qQgC
dKNF4efFKBjkmx3/QNHfWqwJd/PoY3gqSb3yGJQRmTx/2+X+flA14eMTRXOf
n3zj0QbPSj/z3ixpsRfPsx5mW1wy5q1tQgP4qM51d3clk+3azEUCmYqU+Her
KrNOmQhbZPgJJe+FkYku/8QP4DtI/c3WhPfYaOI95xLznqnE4BgxV/J67lN1
TfvgxiAX/oIGYLZdYSVLMlPUSOUmlYwAGTSPDNocMc5LuGECAIGpfgzJMP+i
ItpfB6ZYciznVnwyfogTAoKnbO0Fl//0sZUDj08rj5nBnobrctCX7CuN1cr2
zwqoIE724r8X9st9y1AE1KosASxWw9OhuNyRsA/R5YnXdP5Fz9EDMlE9sKo6
eXuAgpAJ65xf5rrl2HvbngqIA88tL18LIUaiPqoYX+21jM0lBYj5q/pnB7o0
pGYvJsvPrDdB3GCTcUwdXnHlmA98Eywy/Q6AqK34r4+yGLU+GpbmPtBuo8PO
VBgpxOwv8vkBR5TV2hocvBx7OT3g3MLBFozbjVHo9CJiEjyp4QfKvO1pv2Uj
xphq3/9Z7jbq6nc7Pdi5tq1D/Se1Ukz0Uph7/nxAM0h2wOPIqx09WGJuxxU8
BrWpk0Z7/nb973DO0GP/jwQfPyRDYoSJuF5GEVqtHyTJw6TcfGdCsed6hJhn
3r83MsShWZRWFBHW4LhJ9h6EKbzW9LzpjuPqtUv2CQpMh8o/X5iuvA2lIkzP
51eEQoWypsqEgW1CRH2qC9ZyHURvgSbvSny8S/qexGW2ujQlZgP7kccqMaxL
F8M56WKQ5baburziYepAsrHYOLhL04RjkfjDcPrGMYHs3qhEwD3U1r/zl8L3
2Gz2YikJfX+NoQP37CHGpw4nqkmpqXydB5S6y7/B/nBcuFfVJkoDY+BCPjGj
uKRgRGhzsGRzVJkgdOq5vf5xECpmtOGso49cIiGI7Ujqk54xm7oV1L8koh3O
BcmBQQe27eXHoLrAfDcqi9uRAPbXcWzSxfp/GNdic3Da2PQGNxCQTcbB9LW8
ETCeHkGhrY1EtvkBjth8GtlqH+witgRxUg+QR5Z3Kzfh1+z5DGENydUmg6es
xhGXf7J1xE+Zplec7gTC0ETdWcaKQc8nDzO2y+5APtReu+06u/QOdJseL9fz
vP3jvEk9zl28aIEOkLxGEaZ1WKa+I8FEFF/Eb3KDjd6HKZ/Fs03eXBczol8u
P56TjEQZvckmy86ktPlbhOb6rkVyXIwGRX8gSOi0fX5YnCBweov/P1j7oGCe
ItdYT7SOiE0jFs8pB4Izg58CZdj8k3PyN+IpVi985SFYU4cBiFcGK9um4YjN
xgNxX/VIWIaE8hL0lCG3LWhoRLA4+wYfcmUr3CLoOjPvEE7rroVVXN/ic5Xb
Ju4HBlFmN2oWGpFzNxXBSxa/40Hdk55hmqjcHHI69gOgj8LbycuPwvx7uJD1
hYlXVbFrpX2+0qcrYOUXqiXLCrGV+j5bUu70fOZmAjBW0tpBbWDWeyukTk/7
RfNLCOWWNkxbdRfNaCVbkHvxoDsxHPAn3ng4cR39s/ucL6tZjlq7FFnlLJ8c
n0Btnd0JCd/sUPSgX7q600+LOZMbUP3WMD3JInbIAGLfBrH74ectq7toiexr
5gM5UaCrJXwpYUcGnBBNNHY81dV2ZRZH8xky+MGibxqfS5id2W4U0ffV9RNE
9EtzrJU+LnRNSc9uxwaQ4tQB5M1Eeo9XrU/13xZRTs/HRBcvkAX0AOsJtSKL
7GAWTAwXxCs1Gx8r9TDd/g2DNMM6XLJL/j80PJ930h3mPvckvG+kE+5r8tQw
omODIGR+iPiOtdZBmH2Y3EuMlMlN1WOvw6y/W0Wr/mZHCejV88WdYh/pzQ3k
/d2s3XvovzESYw28Y5WZWW57X0CP37PIUNM4aaGbppXs8PcfIyNmxiW9pdSY
sBYZl1/kryOlDxPSnu0eu4fDv2nV6NrxZkVA8v9gk9OAazOfQcTy77ipqaCK
sHQLuMynKoZA+fzEhffOvYL8JyNBERNfK6SBQUMx6hea/WRhHH/R1JUnUm3T
8k889wRo2HyTjzY+EThAc0pTs6KE6rNKHA2ppBkiTJG2sHaChNpFMti1YT5J
KeOWx8xCax2R5uTQtSDFehUBkmHMsNMAmIGvneH7RL+QZoBy7sCip/QzoPfZ
op8De31arJRT20hDVpbx+VNewzYX0duryppT1tn4Eb01P2aY3cJbVZX22owx
nlOq1kzw2pjZqCJ2C9gHw0D3pHiqEObXQ9Gvh8yl4YBX6WDV5lSA2NjuTB4l
Vof8456S+o5IHzAG5JlHmonOZtRhhH0MKuQIOQgeEwwfYkxauHhDzlRTtMx2
0L5kTVkOqPakJtQmxrLxuPxDUyOpcO4ZgSVyy1a2Up3TeElGrp6Bi32IpAmm
cQg7Qd26fGmNJOS+zAyL7l5emDoWMxdgvznmhRbKUQFKz0l3X/0Ivwrj7d+w
SIG0Qnyj7OJYo9mIot6UpC8PNROUeG6Itmg5o8eTzdS1Gs82pdrZOb7YUEg+
q/3gj31LvG+qYuGibvMRE0paedJaUtedSXduxfL+BpqrZq38lx52qICOTnGX
Si5KVCaf51JtBsxuKgKEd5rhXWPyEb+LBsxL7W/9JbOqTeXCCOqmv56+vccF
nKCSevEFS07W5fDe/IBNkAkdZisP3j/YWb05+TtoRfdpPoDVNukWjo92ACpV
j124XxagMf+omALBQDA58ob8IT1jw2mbr1veb93366CVsRrrq1ZwQuA0x9+Z
u3IZNzvKxqHgrMz21Qs1hX9Q9JmPeyOs/zak8Ju9kXonLhiJnh9WTxfPuk2s
hqi4rofXlgdggMwJ8trCTGB7e2vgRKJT/Pb7ptSqEzmEiaVm9gRIfNTZnRTx
Jx2i7mIGgmYHa9zmnpIun58vRWDEDUQdHnN8sdh8fB5eWebAA8ESia3UpvCu
6DuosNf2UILbScNGZvbHKpJwVgTwiaTSwCwSZIMo15kPP0I6XSmYEm/shUQe
cdRhQZBsWdXlTcwUxr2HKZr7WNDm4nUjaQGwkQJdWRkHJxF0/72j1S/09K++
WtTnoqVexwCZMu7BdTmntXnuAmu94CIj3Rv++DRYRJ4BVxP+sxu8fU715b+m
0ClH7b0TNht6+cRyIVUT2xwEKHgGKgzWC9ci0dkP6LsTJ9N+kCltDUyiDqkh
qp6Z5arNTg8X3kF8mX82vQHOx6/AAih1wkbizsZJy7qjHDAGlhefsmB97RWk
C1lE7iBokpeW4nN4F4G3JVz/LGVH0GTiA+aVl1gM8ukDrT4jBa8h1d/7zV/6
Av1cPt9iVHkL8VHIGCRGu0063R5+TjbntjarbB6t1AI7xkbQR9cZ+X0TKIyi
i7m07S7NFcm7xZjCTmZXohiYJaBruVVilVwbS6/fGkKp4aCOnbnjarEwiBL4
s5Mui8jNpSP04GY5BnpfwHstacRyOKJga4t8Ll+HH4N7TFoOXU3M0EXPus6m
zjAJbv+NB0UVx5VhSqP7MDUIv44fdd0v3JYxWrhECbhLh1q9/xHmoPJ+HOA9
zIgD0AiQJjF4cIGWbocrFP8NJtoC4y5JWHy0FipC7idi8bM/4FbPTv7AxQla
ROHIpwGn7k7+KuLBmn8x+mBdzjg1ACMqb+zOJrAf8aWNbJcMa/dmeL9PI7Yh
V7BRsAPqpgkrKP2l2FdNtr1g95ZVA4G7hRwlY1xNbyDfAOpjVB7nDQ77m7e4
2EGyR2SaySnLcjqjAwg/ANWjJ1dHryZS/Jg70HfVRYtPHLMzo4LzKSOCf6IO
a6CfGKh8wlO9RXzM2hC30s0TPt9uscNeCE//ZwyBbfFjFWDVTe4AXa3mO3v0
O4FKCv5vgiykUQDFeRijWNG+DN/Q0fjqHYNcoQl3h5ZVoZn/vhyVvgsWD5eN
UmLehWfsx5ktUaYvxEM7FFJGFszeYQPHg+2khAu3DoSJmjtwp2jto3RMyrlU
1HmB64ZSMWU1FMDhLasnw7zbOehT8aH4fCVxvYSRsEkLKksDrdhbh6Lv5kfN
Vzsu7b5bKX1EVjg9t60Hl7fev63wQmYMo0yzhJShmUwE+vYwGZ3qucrjydDf
AARjbJoP6T4ItFl9kqOEogh+XXHNDEzWwMTExPJithOkHEKSscPhqz3d4jus
gwfUNmE7eQ2aMqYFSVJ1YC0llnaWdEPEMnPU9SVBHkBsve4H9oa1kfyzOIOO
zGKoqNy0AnJgr4PX5nXH6B8G+L5Tr4w7k2aTX71/m6LawPIUjHgtX5YOE8ym
5dpbCo7oPc8ol6t4ECkyj/QPgC/WvtQ3Z6YDY7PZTte6P7eqghq7gm5o5Qfh
GHNzlv7y4cD9VXmrzrud8Ah3lLAG5FKQHXLskWLqH+EHW8VbIztYxHjKw5PC
HyMCWEm3EdDqvoLRz6Pv+wAfspCCoF34a2K8LhoHQMrVUTj6supXE8cnV2Ps
ynEiOeKcxaaYexTPM5NNxWRtxrUa4hATApIxHB6gu4Qnss4hO+9LjUfupdL7
ChUvrCg6UwAZ9N1cTnVLlUKn2SZtP7Gxwdh9OJeAoTiMcgc+OO3rVnDQuui9
y/oygYfj02dj8Ld6qsGfq55RE3n2Qdp8BnoBMVX+F21pv76D9cb52frZmB6W
DGVyzkrq/Nvb8wbHz1/TA80NyVloQzfJTG8IHPnz5HHIXSVATEW8789GXmYs
eV4HjuwbW1vzJU9qDzsH0atiTdYanPVVVl9o4J66/fnqI9+ZdFlST+p3id01
rf4qr/3JtpOMDz+SRIYG9hpucj+3jLiRUfOYTkFWmu2kF4tGgy2nkcNky8GR
+Ma2S8B+fgUifkmr6ZwPu5QGFlhXA2+Drc4f0iesiGrdNh2hqa3f/YCCAI+K
10jyowKrtNL9nay54FbUx8wMo67Bh2eVlGrrO4xYsNztSN7D+hsjy+f5JaFN
9VFUtVPEpuzmETutIDsc/WBbfbqrK00LO0g8bPf6p5Kx/0bwUfT0+GbDAlyn
9fIIVswGZAyWAzUaPzYvcUZtR4hKVYJ+yjuo/iEgnlPgatSP8Xd1gReCgH3s
6ULfaGwiyWlB4A35OlQNn6WcUYcogT76hb3UdQBrSFOKWMUyRI8OHoaOY30z
MN9xB3CtQJ2+7QpfrBd9O+ql5olPD8b4Pck2zOHMIOYTaDu8Tf0ul/iXyuO9
SMVJXftEtMz48j4BsuD3bjT+38/Ost83jfao2EzQ5ibv/zZdCIYz5XdsbXas
EVeC9NHH8lZ0VskKkNIgxGwrC+v1W8fqihIXlHtWxNuqJnyfFtzzKARV1EZY
I0P7qW8boU9HVKCoH8DECfaUaDeA4iVl1L4UF5Fhu4d+LgfwhFV29Ef2dmgN
HW1Oan4k556Go2t7Jjeb4QINvXDgMm1JIPSIZdLUFpQkA2XHDtmr2WL/hOI0
i8NsE38LiqXvF5M9o8zxTvj+6X8ZbmatfAz4n4WQss29D0/wjf9YqRU/Syll
bsMybJIQlDw+ALGSeaglcGZmwez8hcJFJFrW2v6IaksHQZuYhyTel0SMzhHv
YpFoDfG3RgyuURPf9VwjyLg0MQMSAFKERNfrMwkZVbrDx6YufyMWo8Nb9z/E
aZoMtrSn71hW0U0drFWr1SZHazXZHz4/YohS+LsCM+rJIig2PoggoIE3dRHT
2udfahJna2+axWchIuF2Ueaa/dcM2upN3Lnwx8OWCsH6mkNhueKXcAxNA/ba
Te96d0b77XpjfkNmbogx1Q4M/YNj7oPgxo2QbsXctxYq+hFmL6IOLXkmWz/9
PrW5vEsAg8WgVRia26YF9YhHTF10Srn+N3TUe5ZoU0IbfpeZl8WsReO+eadT
oMxqSD6pejSodmW3B5QK/vgAycckNVuTlrLFhcboqiZzZSkecDLYib+JeL7X
j1qLV4nWTsjGq4VkrO8ByIk3iUZoG0lM+bgMzz3m5TOAKoZM6sZl2iZx86ab
4tKOIC/4Zx6NlLfm+pKQRGTds+VX1HTbjBB3Bd4t8sbrrPeZz/QaB5JnywHL
PQdO5riOnpJPE/dUAzAUbui7kGdPZgk0i6lhUcrN76P/m15f/yesYxL/zgcs
+gqPrUUGcV8xig/aCGnoQl3BY4iLiHx3X/foYjFFZW/4T2Lntrc4MjPImxUV
vhTEH0Mrn3k/8WavlCYbpUy0d4q3kBWEdOWJ+ImmRnqueIYjMGLEqW3wYPWs
6lgmhfwNXs43GjJl093HQ8tQN2FLoZGiOla3poePDJ2y2ehmWvqan/lrIQT+
xRpZc48qEA+axie49u6dLdqCvGPQp5sy45dp/QUq+rxmcDlxBX40bCLJYUvR
KfRyLHqF90vlELDbwRV/Purv9baaKDdL0DDjEhTSz+5lbahFk1wmaZ2x+EnM
aVYRLbMeo3yO6DHupTU85kwCotOAyZixLkwh9T3RDkZp/qMagayn2AA0QfAW
u/ED3+IS+jweN9XucQVvDCp+Px+uP0Jn8ugNb78TrF9mAaBchG+zXrxnePMU
r1xFYpgPfYZPZdFXKNjXXVnI7NENx3JGPq07GEoL2qsiccRFXFQt0YveHlrm
RUENz1zMEDiGqt4yUJQquaFgmLC+0uHuj8jh0iOxqbSldFiu4b1Ubdq8XaZo
V170a2v2ZmxR2ZcWiLxDAVwuSWvwVvWFiSNToxpjaauHrCJDYusd7XW2stli
Yd7tUNVG3J3ITpD/0w0MYJQm7m1fo4UcQ0CvYp3loQIuZ36PlwIFKqU+/Kmm
xvrAY6EubkqQkleiS4g3mz4hNZW25bUojqJlCA7hmrpPWpfSmyXFK+VH5s0U
0R9q8R13H2c6cOZzgRbznrMMQPv9eN87R72x12mOUs3z/aAJui0v8HB2/1e3
eUFWbxh6IPD26cX1qDujEd9bkX/uXXN4tRuIS77ZcQYtbRvbFt0yhNb+C3Jj
zI7YeVz0vvO+pt9AXDRKTEdX7YUcy2HTXESnqkIFWZGg6tocBXkYenN0++mv
W0ah+j+K1xIpoptWrqAqIndYMrFRJYPH/LxzzgmtzkMuLGRu1cp9mnSSqgt5
RrHPMhRa7qP8UGQQDU1HTbwbESwuFX/Mui34TPfn+j5+8FIkKBDCmuuWssbI
py7qA3/maX4hxY7ZCLlCwg6IBi7Nj/gKAVBf6y6Ur1klT59+B6zG6StFxKuX
7mfN8yKQtYD4jeCIvYWoBDbV3/645lqok4fTTqP11C+1/FZPZDJvWoit12RD
XLOGSv/UCWAP9T9RboFFQwWG2bx2+gi0U5kxOhS+Tde15mYTyLPLd9rracvn
O6c5EAZsoydO+AkiHZ08bZKWoI6H9te4ZPal/cCMLRjHRDxLV5ffV3IRU3h2
DfH5u+lBmQdkbDFSfqXpKvtPgdQfOlLDa7+wHfC8Ss2zOxJrACrfDPRml+CE
1BzC3rviE0Gmof/Pmmq5MZOO8K30/8/5qaldqkaTlCm7UYSwlRvQ7qHjzYwE
4ErE2ZX/sAga2luMg95wdjbXof69TeeNY04fMZpUmsVodeWjsDpkSHY97ZNx
rsnfWA9WYe1Ob1t8okPLYt2xgBmcKv0VSCy0OZmGo24nku9/sizCfvMphEZF
7j7gQ8QfyjaQ9FR3Z99dsqEU5Saw5Ql7uJmW7w0szh/130h63hYpOh/dbMrs
ovhYM0lHkq6WqosQXCjWeC1k7jddaJb22Ro5nqsmZVi1k1OI3n8h30FX3rXe
9Jg1TGmfgSIy8ZIehRKX5YsieDtLn38KljUvbR5JnZjDRWci50o9j3ptgtgE
cc8c2RVhqWd1/+bd9IiF3vpLIOka++qPASI4CM2k6CerTVuPiEIdoVD6lrKH
v6qmQdByIVI1OQd/gvsxFuELY/7vmwtBuK8X6xp3q3q8HnSQ6fM91JHXcbYY
EnxfwJ5blLCzLnjDnsbTvKcx3ocxwhsiTh8DSEmZEtxm6qnV7mK2dwDS9iX6
Q3JYU8syYDRq4H3rlVJYr6tReiSIHCVfzrOew4BTuAn9P7FPfTjkHxylYjnw
wfjWL0l7m5BzrGP2naPPZHE7zTqP/aqw0TgmhGi/VnCIpxiSqpkvnbj/npiN
YWOtNwMDJ51kbT400sWi3q1g+jBDj+qtJa+L9D1TXdet3gevj38Ga985wthJ
1h313/dHsGH8VqDhEVi11+xW2q09SygrQ80+GwC4PL2Di5wtSwIFO70zXx2H
5Ho9kcFZoW8/a1oW3tOlgmpmxKI5djZzQu3URGOzKt+MNAJi0gGaU/rejtxP
Yxm3be8El4IeZVGUxSO+3t5QQWBJIJLOTFbGLWxbrHMrsoB01YK9T9G9poDx
esJEnZdkPvsPMV1Lw7F5l6vad6oUlIAV3reROAHdZHCgQc7eISyrgi34aFe0
EYkNwhhMFWYFJb7g3mYpC2GtYrhi5s/BSugczfn9sYTgB4sPnRRDS/Z043U1
mliLUE3fTxu6yeuKgRav/shsrRbn/1UsP9Dj7qU2YuUW4jI7acNZkRTGzqem
3fUaqrRtlaY29HutnCCJjneS1InRvJujN/QPEL1fy9FW5KFAH9yHw5GowwZZ
PkbQ0kzOJ+PAGsBPj2lMKaBdxttK2tiWIhNF02l3ko6E/EVTdmnls0rCvZWn
JTveC3rWOvKMCLQGxGm4XY2wByQ3fn6kSboXo3j3GGtbwF/ZcA/TEnRB4dn7
XzPyPQNaTuIZ38EkliQ0hudNzmUzboyuDjxdoQtT8xFkyufi5AJa2rpQ1Wb8
9D56339juaRvzcj5NHsVgXtSFUQh24gj2kUvELWlaNDK8v1AcDyWkQ/AAIf7
Zl4YuSC2zf2POF98bM7RABI1FsoPRZ82ZZ8YkWm0U1/Z5+89UumB7yPx4uns
lI0U5ajRppbX03iI3Lvwv0paf+lUD7g+euYf2xvU7fU083kG2sMZAPq7cmBO
F32plAZnMA9fVmM/cuTmPQo+Fwu9wdjdHABvkgml7F9bKRAj82jz9sGwbqAz
6TBq7HCfK5IjNI0fgybG8ehtVsdNOghgp8/K3SU9oBV1mRFd/IWi0bdSwl28
EchHbgTD4F7u3Gy5Mf4W2DG6uUMnLnhMk/8zClaNy5QN8XG09D/wS1hWL3cQ
jsynxwDsy3NiGaBRQxWtRIlzgfeVntkYdIaGWrty5KiPw0UwzewHIcnJBmkg
AIsxY9IaIdwRlyQWevK9acjvuH53Z5gGiRFMUqPutIe2CmTo3qU+Rw7+1u1e
NYFl19MslX8uLhzezSwwNFCVXKSc5f/iPW5JfbsbwTmOnOn0rl7CE8HO8i9S
DM5pTUKPIxJVKYD991IiyGM+V/IogkoxgJZNSujK5tFqu+uyFnxApXuSbq2c
5VdyB9HDd0gehnDE9wBE+W2J+w1z1NLI8v68jOcF61GVlSXODnlZrsP7uErE
Zwlweme58OzjeIPipfYD+33YUUrmCPrVHcW/z1QOX/s7MggpYqIjP/R5wC9o
Zgy8uJrV3bkanEoV/oKcrY+dKTzdARpSbH0ScUgBoqXaVWiAVwbNgzB5zpjx
uA3ilYOJ/qNI8jKiiYb2TOt0BgkN5RaYkrai3g12mZWfbgxeyyCppnH90zwf
LLBEod+NR2fp/25jTKu1jVLIzWPyFYAxFzekch+EiOHF0Sn12D2432z5MeYh
Kat3z1SnJJKycd1MPt4l9dfgN9/sD9Sis8wRDZyavds302dFriKjaK3eGnho
BYaxpr1ZdPx6+c90FZvbmu6E+yL7iqA16xdVVHl1Gqjry+J65S0kZMQan3u/
TgBJDobmCJ5J4RsKSINgknZIKsf08URT8t1rR9yqj7WYH+JsbD19HxwWh4mC
iTAF83PqE5aP4enUxCLI9vvpBNG9AS/AJ1BmeIwl3Qn5i8I4YrjK0kc//rVf
m9XESa7za68oGLzRLWV0XVKLp5YfSeR7PzWe4w04Py+g9azzPIPsdPxu2YV4
Mc9jtjZTFYEIrBuSvbshEGiEEerG3Ae7DAFIf/ggs/IvUGvDEwuNqXaUtJRh
R8pEiXmR6NXuKQ30WHKHzLO0CkLcFQQNqQK/t6Uykud6QBCuRO2/V4+zasOI
f43lOj/Yeb8nI/+PaDQxNQOjQD1Y0Dbi51R7jz4j3JUcpfwqTr88LzFL9r2o
p7Ctt6rrN3SkhrwLkM69BDhDPYLyPpHgTZkqFjo7Ew3Zo8wIccZJpGjLaNen
3lhhOila+n4mWh2fui7SOw2v8SwGpbZLDoMj6DbI4lDCfitKy931KvCyRAyg
2LsCjbP6vVV7x8GUQ0OzgfA3h+VA7FazggLtGrosNV+UnEMtW8WYCK4vJiIJ
fWQE3UYLkXN3UYqBnFe7afmZFB8WWevlGYseemqQu+2spIZTrVuRFHgpbEOW
yFIftzJVzPrjlC2nthhEaO2LDONJw2f9tJDKZkjvcYe03viY9Rkuk7NIrlUq
iclvw7Z8In8/fzDjSoNgMMhxrWdbFL0Vr0IbkmhW8s29P7bOZ9TBIWvG12mc
HX+P9wR2PgBxWCf0+E+91tjEavXGoxXEt+1q4iOGHkjpDqhyPzlqVp5etJUR
7dYF6UTuvl597OgzjDI9pOVc3urGBescZWgP12juxrJAZX9XZaAYbd1ME5z/
777tp7oBdURBwvA0tt/GokqNIk/jZCedR0sAPEoH5dKVoAtpPAL6aI9xi8ri
jwCHKvNnYLJ5vlU/EtJkE1jxkh7wmgbwltKKes/1rwiY5E9bu/83COva4Qse
gRQfo2W8HiDmo/fgdhLTPVEomdMNw9EP4IVKMp9uOaYZ4X8MgshhRMvhqBeB
AERQGdG8Ws1ZAnDG0oXgD51btoLtI/WuEaKefX8jozH4uMUlimGJ8ZKJyV9X
imp30HnaqJpxeps0JVD5pjLuLHi//LrX/zPF12l5wFMo+KQnX4Ybe+XGz3h/
OqnzfJOWsyoUyPVIEr19qxjKnTMtUk02DLMqzKY7HMElU8BkppF7VLZgdnhj
PL/LlbcP1v/XudkjZ6hVTGOb73dvCpdAhp04kn35HicJ6eD4ZwZ9TUOiv3uA
iBCP9KqjvFGAaqXf63IJiQnXLfWU7PmD157gbWEr4rwJofdGCLwjxiJguNxc
4X2o8wKD9aObSp+hWX4kA0iNKwv0CEUFBoZQkzd/dHh9C5wOKVpuud4W/OTg
vRgPXjej/5My6IhJzjKDrPV80+HFmD/mn2ccODjxCxtIqGdRj0NKN+kRQ0LG
bsdA6VItbpVCuXTGsPLqZEoLUJ77IUWSYJQ9MijUzzAbtSK8+t7G6iLQyvY8
Orm2s8hn9K9Hi4BAz6V3P1VUmYbYK+Nik+N1N8O0wqWCqHAa9yHnMKDJOb9D
38rOZGATis9faaM7sjxpiMo4O3y3HndCdM4Vui0S5M9gYdd6jEFLXDKgvFAw
M5oyyiz4tmSZDB+a+g7jx8LMmpTv2457Q8nkVkG+krw4riP0cotjuzUDvZrc
JA8LcosIDqmntzc9XgxaOtgdxqPWVr9KifP3vDZ0m1BKF22uBTXRzdSHo+Wp
tQ6ykr8v/6XPzu3HHS7OPVkNZ9mqlqtrBmiFU8ByLiekXCvsqxYT+WA59vpe
crNnbg/Dzh38v29Gb9ewzl1e1c6eOa8w0kvDd4xUdCl26mML3f2Vy1p0qeAi
0I/A/aifN5cQpaGA2d0P3xUBW4/OhjB1pjQ/ZSgVZpPXyU/BlsarfhM9BLw1
IajGGISK9AQADWoFkDT0RzEdsUV5/oZMBaOxyb8YLcRd71HZIZK+ny3XDujy
MPpH7cmC2IW4lG7kqwjirNBKgb0oUsGDFdNZIylRerD8JGbLir6Xvm7Xx3td
vT9n3DF0c3fhQNujN73p4wFzsPwlp478Haw9SJ2Ucv76YTXKM4vPUmMLybg0
DAMlUmJt0vQXGqPaH3BF3Sf6Ty0cvL9YPHixTguYv7hgBwwpo6djKGrs0DMJ
ur35EAc1wiiovD5nyRUgVu8KaMhm6QYfZmWu72RHKZ0cPxXNr8guPSHGMWGk
ueQunYiMMpoM7M9a53OJcxiUktOTt920yj3gs/hpiYa+zTvLLEn+RPfbJXAv
vgvPVTp9Tt0uql/qkFRmfmQVT93x2oBeeetQcaTzlnURpd+qhCw2IPwPsn88
wxQwyGLAL2pEG+qHIlxMZDtnsg4cz5Yf2vuY56FWEjQ0uA09BAQm6N2oDl2p
iR3UQ4r3Q4JryXkpwt0Rsfkgtf0rwx/RdR+9bp8B136s1OmZLnEIScySsiMw
XxYnvmJic3rfYBfpDb/v8re25ugu/z28kmCxe0wpxB+5z2OPjCBsD3WFLFZN
9/vTXpj1Wn94vrSl94bAs0j9b83x8bb+jjedZcF8JPUiJaCwsRIrda/qW4O5
a1T3Cfbl2URv2KYSAuPa/HojP85WOHUFyjv2FIAKpGtdECz5dOv0m/cTnKdB
xCwND+qzuZhyXzNNeuJ1Ppa0KHaDJ0XM43okI+ponhAV+u/swvGx6ErphPz6
d/R4bwM2jRSZIQVEacIht3kFq7zG02Xt135/Nh5F3AFeu1sS8zJLcSQlGNtY
TZK5Q6cHMU+F/6VWAekdDut5eMuiKno6srSZgOwD1Fn4LqwDS++4ubKX2rlP
GwVZ766UY3JNLBmezQNXtlniUDNpqoA8PVWBgWNHJ8PKB8EhldC2neCAJxwy
XifYIIwaLvlMRW/R3leAREjOzOarQ+fJ5kslXGNosCH45MWlydowYYi0HWl7
MIhZ79fS6eLS3e95nUQ1aLL+8kpufxQOIPTtQhJ4iGZnEY0VyirgiZW3lZz+
VjvRITf0mBs3ADXcHEOjQhOAhbakpzq0uWFotRO5+BJ15qwGtZwFD+a02Iqc
MNj9L97+I9gal/HcPfbCsHP1klb/RASeI2MKSBz1aKVmqorChAeY2/8yPmFK
N8wWoLeBCIC0V41lKedD/ljDoVPcEuLgqiKj5JEArq8KGwlOhUxg1WOcHuX2
M/phIYHUVOU8jjVDU6nLipH7nfZab903WmgOBe3sOoHposa/OROgAuRUDGQE
IBGG7IqBhat98oOGDkv8+hh0ArUsJcF6A88kHxlF0dPBvsvkB8JewagN1XwW
wnIkZUrgotssjRT7y53w2C1owabGPPMoLI1E8Od49Z6zqwqMmjbJelXEYRBv
608rBQDVYCXfKDu1k29HQJX4yZFzC+6C7syDqYZlLO2c+pRF09uy2KBbzgO7
DN6v75pH61GJ043FOm/L5hNb0k77b0HrLw/e+u3e+qHkG69YqoI2HLbSxSQr
Q6bmlwxHW7i21xBedool0D87zsT4qqq0lgTagDpJXSWAt3bsP5Fo1nndZLT0
KgiahQ4KPc8qZkcagJ/g6od6tcq16YTC78M8R3FyBf83kVO6pGCSprhcwX50
iTXcKEYQzs85DjNSJtZv5pLJ8qLQ4rHEc0ahlEbG8LxYez4USxg8b0K8DEwY
S6QsJeR2wG29QEBPQKdTTia0G37snLBHM6BL9PK6WNUoXn3Wu/5NIP5ShO9R
2M4LzNv8HxCa72301M6dvtVliw3DCbq4qWW+u2TSumAPxk6b44QyZw9oaCiC
PebXF9nMB2wscc4rNLQxSx0V2oeSCphLZiAd/akiMXcEVem8xyKDpKWpdfO9
9ROVzuIWMVv0i24WMzqOOc+SXGZ9mI/uLTPYz3faermA7+snUP1mJShv68bK
GacpCb9xubaJT+e+EjyPoFkLlh2jyUdnJP4FuSiUA8b8/V7ivotw6cvc8DgO
aXdbZPJWXD/JYQuioogB3UAelBGbvqndMDsIjY1y5VIgCT5pYlkVBkDsjSSD
uTu0p+2sffDK9/Xrr62tUugOw0f0LV0Kg7CIeIDjDMzxEfaqm/nbSH2cPfOH
GH65L4TvVqZFAOphth5OBeHmO0x8oAhO5d546hoQjz+COfLhbSllZQr3SZ7q
LVYXXh0inShmZRdOdnZy7cFszLsUrtb+mRdtokzWHla8aJheBMzsnpBqJORT
wgHYWBuyhux07SGldsLKtc51megmu0B1s1NEjSM7O35Ah4RVHuqYL7PXScy0
dNtuqsa6t7mjrmGDWZVYW7mNvqYrgaBETXhvqRUank7odOCT+R/gBavP6MqT
Eh1TDyfACOVRw5zyVbTBKLs1KBic3tIskKQMV4cgBRrPov4ed3fmpkURGegv
dElZkBUqeUtBg5omv5+w9BDc92CK60luaS1ZhSqziMNeuRbAaHGV7SOuhX3l
nEICLhCA5Vnde4DC98iYN1tcEOjgb8ottrYkqldJhnODwiGiIAK9Oqa9Xzpr
eIPSnR1hpyJglASpcfksqaoaw1/fwmTOQjjKReOIIPXa12/66jOPKFDO1SiJ
4joyF1NtRd4p79K9nYv0LOVOLqNjxZ9SulTuLhThNEL+/1QmPb6QOH3oLd2A
sND2w00ynRdI7B1nvNvLYTsnNO5SnMjLF2hZe1+qPYzIm0TS6AqgMIkaQTqF
W5kR+CtTm90CKaIEqDzPB4eDlLjgb9l1+ABCf1fixkUosycZEkgnSI1DugPh
RAw4s+dekSB6V7jfigW5XQ9/VZ/iL5UNpySHSo05nNDh85IibLi4p2sYUDt/
YjMorZyULz6BI2PkX7Ob+coDs1Gem0DUId4oyNTKarafsa2RVp1xqirh1FPJ
2htOwoJSYqfCYk5KPfCedo6j5K8HM8cKHjrpvz/FfGXD9D+afPwTFzTm2Y2o
h/5Eib5VEECURRpTj4JBc1cUgdbunCSEcAapTxWfPygRNQ4bzNfSlxqUPP+6
QRX6dEcy/fpJ9ktSfJx+bG1VcKdH6ae+GMspgCmvDZc8l73M5sf899+Tezod
lgejLsTBe0zodx9AzDPyy18L4Qbb38zQj0pAlA1TkPn+al1U7lSxQQpzoo/I
eyYTII9Ef+3HlzybGIeTdcNlhQwEPsrWFA/0vJD55vViouVe28J6oEDDgHfX
G//MKYEKMppGS05r+zU25RrC/ydWf54TmCXBIzvuK8eMi8N72c2SjaHFItj+
DVCbczN/wpuP2g+J8UqPM+1Ey8bHuw7jPnASAAgqE5x90TsVFZLyh5MlAc37
6F0MLcxOrLGkLSpQonl2weTwn5V6yvTOfYV2co8NJdg7/voHsDDCLvD7mgrp
xumyya5g+mHrKxkkr+em1Dxva/+zmzosCoeghK9oyTkG9AMDAmnSL13M2b6T
HhmJJ/dJiGv2wrSSL/GpmRse+ukKF8x0K6Ddx+H1aEPEjadAK1lXqTQzbcpY
7ApwtOXzzO8xr+DiENkpdatZYuyTiVk9q5YE4ulwJnUj60/OKppHEXAllk7F
f4xIOwRIaGveb0VQDUcmkAxW1Bl7FhHaLu1anoVllfKvORrKE8iz2yxR4zGB
+A4fK7ZDmIXBdwYVTLB0shtBfJmYtHbHSUaqrhIWKGotjkCtvdKApI+YL6bN
kxvzk6Q00lf2Rhx0ObH9YX2i1XmZuhhAmsaCP8Vis8YmOPBHMLyYKpLD0Iub
pxy44SR4L8jJieNwUvaZTcpxouIt8ygX8RxLAZRne5ZQzFT9B3YjEL9xkdOe
DNREn2N0a3sq26LUyMdq1DYJYPy9NSHCQ3OJ5rY0iNThb1XcYzODlK5rSGOz
FRwwm6vUPqGtRoGbdik1lpf1tDU+FQqNQ1igKZHyTPDcAOt4ttHckEomuQUc
2QUIuBAZoXEVQykOn82in6isIqo1ngZ9xGYzDo1IMvf+Uy1583ucx+iLA76D
TRlHbMMDffgOfZoTedcmAuCosdbGPVviTkNCtHki46facuID0jWaWxvHzk7U
FtbBdOH8FGlfhaPkdS9EkbaHXCXCio0dHY0uK3Ou2pYfMxVMFGbma1gL5kiZ
JvJHak9fSmDzsvY8q6d60C2k/TULKVbjj7Rdd62n3FDTBhIKeVt/QmYaReZ/
dSkAUnAT/fYBWEE+DDY3BzoALCxqTkd74Ng1svJvUMq6DmcatsZmdIUImXuD
v1A5+2oFkZQ7so1DmFhAT047UwkGuiy8zttCi2wpwr38QKRlRE6ieKVmLthB
+4e+JISc6SV9IDj/PMD1HqIB/LgKisGAeTITZl8PFyjD9UJECjxDwPn/QoGK
kM0MOXfYGuOdL3nwugYqVTBakUBChHkeu6XX9ISIRL1ru8vPp15kiLDERkpi
ixVFfnczG+my1HwX/XgGY5pUvh0FRtWABlPcwoWW+greg67eGlbHg3WQ7li0
JIYdLk3gynQ6zh+nKTGdPVJDt3XMZ+DACyX0nnCf7JdWVENHZtIhxLfA92iP
ZreIhyIXJQtH9Wn7Qcyf/yqO7/gwYaLfXY6iPD3b2VCU6jswVsyRKawc5zuA
auqCFRfllZWrhrSnd6pU5tGdAqQ7lBgD5Mfm7ZuFCsoZQkcj976nVzDFT1iG
SAtGxC3wnArH3v7JpIfticyglp/FpCqi9U6w0EHcHLbqgoJpX4MFcC0/jJ3l
32M3TYfZMN+lPYLlA2qdzEuk+fSrGDAh+7Cnj9xqIewPrr3M+nIZmLe5WASd
MPYRdlEgVQuAxGmgauyxoBC+Al6jegXxRODdQcUvBDl6v/LJhU9Sljgf4mMI
V9tOpGvb0FW8xLW439E3xEmjAHlbw9H4ltwp0MCN58Z2duXTxmWK8Zjs2YT1
Ya+LWqj60+n5AzcScYA97fsOcjZ9EMkTrwwdmD2LoW8E7LGJcJp2T6l7vB6/
D5HFSfb4dEEb6kFYsQy3hld2r9N0+T48fmL+GHEb+k3ReY6aK5YHJrDFXNd4
n4HbQ2M9EIuyTfv42eWDGGeqMtVljT5t5r8dkmxlTZ8FHiHUIPo2+6vbs7JO
KDgcSmJ4bTNogw3QvAM9Q61/NjAoXeU7pfrurSnv4XR9eG7I5VARZtb1HHAu
ypIYEAw8AgS/D0wwv6VVhD/rwBYBTVVgB4Z7T3nr9dFUmTejdX7qLgU0BYub
aWBdkex+hkUtvlsn3xyAThi+QdaFMH8b9XVHMDwA5SsRNGwGzRU6MAeofJC5
oaBYLSV6dFGmOfhx8ShNAu3vXkvU6tHOHBYKrTxTE0ZZ5o47OvK7/4XTNsgo
VRDMdQYGFkKYbGi9+LiSQ4DL0kxh7fxonuD6knVQMqUixs0gml1RVkyESkns
ot5P4QdTpTEEW05mHY5BI5GL89dGvFRifIh9IhUv9UnKLHH4ZRduaWJYrIvJ
evUrgQftJMnbZZtMczyxghuVLGVTmK921YeVX3Tg+mw89CtmHMMfWAZVu+8g
0yC5oJAZXl3GGR0J+rPZzR4lYIMuxkHCt4OBAnksBRKkJ/XQiXegcEhOBkum
3XWVcjhhWghq74nHStS2bp01cNY+Yz/kEg/Dvu5nD+YyAiGiSgvxCia1wFgp
53DF496c54xgdPK7wetWyFDw1XdvGu3W+kE323QNLDwwF+i4pQDTjr59jCJb
bw5Pl59Q4O3j9KCMQjlWlRksdHCVOvExm8o7WgVNyrGNG9J5dm/+py/7KIfA
YNCh03l736/eVhbK4Bvo28hkiH8kUwuGppbCLMj1bPCz3no3hPKMdhICD1zh
ZqrB63xoPutGgZxv7SSFlcNH8I4j+hF7AJONirdT6rBsM9XuwGEPpBP1mSem
A80PSasc2gCvcxVMJDbaqrM5yUUy6nVAfx2T7cIeJ2OrGF2iDTRJ8jrc4nNP
7sKbJCJNLQLCyhlWodoJNiv1x00uUWAdvNbhumqSlgqRxGEt704KOzFIOpuh
wKDx4GgQL+fF98ZW+XX8ltZsYJMEPZKs44DcmNNMa/i6rWneqh+STV0nYYMA
r7hhVHNV4XzPyjEqNge/+2EqBb+NQ0DknrAHyLWUrUnxHcYvZCa4sPWK+KnQ
cWACKGR+lGszGB5dGESw/gvQPo2K8SdqZQ8cdoAnF3pQtUVSEwrw4sQcczLx
DRH8DZcWWqGiJTL/0BbX5oC8YWeUSibPLhFwZFQI0Ognw6kyv0ZPWl+Q8kHW
46Ekzesz6Ij9rp9Z0EA8tHlbmAYfKLQ6YumUIvRVqJXXlD9Z37+5ENfq6Ey6
PuCTAgyN5GgMHpkRqP2VhMQJCn9G6tGatEEZGkaqP2tdKvL7lqpKw9ge0D0B
qZq3j4NwUlJLcGK8gClkUWSPwNKRzisocgaOokFChI/0F0ReczAKdtL67bUN
sdshR5E4A9djFGipaWwyFPjF2KVzInbKillSmgJEPMOoBm3yMeETyu/aBXzx
7Xorf9n8AMfCdzNThTSnu1u4m/zK9Dx6lIBz911hiT5tXsKS9w+jFl/QmaaR
KKB70teJwBheajvTJsDgyjfZBBUfs3sSibylwCWIOJfNyBIiUpKgiGx1SRHM
kCUxmr5MQ4dYIYCzX5RrsVumypfOawt+zilVQWn1LS4xXi4J4kF0snaNekTi
lLcR9SDgAWxFhCxojqL0S4m12uFhnfRsK5cVU15LXrIkm+zzzP+wvVhEklnk
axNlQ/Bs/E6UciliQWNMjZxziEN++xBnniIz6q5akJB/WcsLPlzscpVsmMNN
Dznr2nX35vryOiot8d0iKTByhcCUMYgg4EYn5O5m+A98vALiKFUa3N1SRQiS
bze/sw4EDoJqm4JSF4ckGnj35gOZBzvKMsgSfDLKmbnfVs62YCkKEehKTOiJ
SyYKMZfW8mqX7+hhQMUf/3tK6sn6+3NTGOzEy1QsNAvC8b3AJ1W0XYo2dU6i
GimZviJlDs3w4cXyNuQUm5j6NETKHJyUZk6wg8EZzM9cLhGgGp7G3GTiDU4q
6kJEl8ny/NThrelJZ77d1vBITzHTzmBMJ546aocZ4jYd5tZ3h5NWC/bwq7vt
wRoJltwontkKSgUTHhxthSklX32AfQcJ6hCBGTYF5rdWavXnA6gJTDWVgYLG
IvEZj8La3hTNOc9anWkMOGJV2+URPC3xfBBRUGSu+j6fDhM8Pvf4Jyhaj5rj
QeESDItEBs92As13d+sDHnoKtdsJqSmrQ9KTxD8HqHy5x/m+MRruau6hqIkW
B+uGcpueFhOjbWVYAwRTfAqzGnmeQo88z5FlowQpmIPaXjSXLKagvWhUiovh
PVqgIta2g5SKLaMW+RS5o4K7pvl+RuAeZTg0xEYBt8V3QwU2/+Lbk31dmx/t
hVJsNg1IYT0QDwt5tAR5RKyGZy7WJfPx+rMlCpaCdrkgGbJueOhJhRULTI6M
glZr8DcjIi3pKbF/rZR1raQCBDaY5Zl3W5+keB3iBSx20x6dAme6GPdM9cGD
tVpwggxrS+foljRyLZVljwGD90FLVZNohWhLSlnLG2T0ZDkHyrikBFYWUVQG
9mMAy5Wl3XKHL3MaBqWDz9h25Xf6VOeK67S4Z1wVoqUTlyhCHyeC2D69LXNr
/5jiYBLbnDy83fVpiThnCypwLuKUJ3ZPd7wPYbpeHaiINDdCfcRkh3RY74Fr
+xzLEfrdYVLAFgaj2ICFjQZvF2ypYCSGOJwWiGIFTl6+5uGBOiGkZlUKYZjh
yGZcBauALJu0bW2yKZYprnoBgFAATGD8KiQd5Ow7/ur0TH15qN5rq5T8HEU/
+o9FxT+awYxZVXqZ561mKK8ZHps0cFmyGRW3ZpBMnsPM+S/uqaCA7j8hLiKX
WTJHk4fJnzCWYECe1Fdj1/VkGoNCzF/nxBTSfZPtNhkrpPD+WGGRPmgLtWLA
YGhx3c6KeCuvn62w5kGb0SULajJi9f+V+tSm4nWcJ17Txf0Yic9cDOiwsuxs
qJyT5jvxi9uQ4RG1ZdHvFPYeX7Rz1lZFPo26Gc0uBfEMGm6Cmlgy/4npi2sj
FB8pomHABJECaJmb3D/ITiQjt0p2oFUnfYnLVJlY926ba7LORW8rX0ZGFG5s
8Rl377QP/YtQla96/nWIMg+y3UiIy5Pqmtjpe8uSNnyHEyz9o65fwPgFrrDv
s1b0+0OPF6cEUJAMYSRzgQKvR1oO+UTUJ5dYlxB5VjUV94u/LYRWTTpZ0P4/
0eZey23/bZDdiVvkbAOOp18yaQG/+35yKZ3at/BrLt5VFhVi1RGVMcRDNmgA
Ii/GpI7wZ3y/1DjujeRYPcoVKylJCa1c4onw8bWfUM/k81cY2IkFGGVEkujB
y6k5RFQ5xidM+yCxZaI5/w4/O3fNA10/8m95nHVqrKsJumgIbyXHmIEo2VdB
RIie5b7/doFTrpO9HTJkRuETO++BlV+Hl2sPMaujT19aOAFORmO+bbjjqeI1
tEZRbHRebaLdfs2SvEYjroK1Aohr6vz+//1ocH7WOYMdT8nDbRj3cl9pA7K3
9yY2jou//huzoKJHRtDFJ3SxO4Fk47J7OzwgLBRiZI/rBJb09NYawia/cWcu
k75UFDa6zY7wh4s3Px+/DUZX1c3VWOXW0r+kxikmHafsyjtf4gXBRV1E6kQC
DyM4N4GLexNusMzIyxQHZMJFk5I+i80cqYx4ndkYbGCAsWkUVzqw4xk5X4Va
sXImdGQxm+7ZD2JkqGLHw3Z3O+7fUemmuwFbnSCUuWvYaPmH8VSjchVcLMbq
4DLDRI9et1nNvR6nd7sffxz0VO1gBz/gw9G+xyWJiusYVjJpiqhrfGUguUOQ
VQS440135jBR0kVGpMqnvUJQNwcFoTEQRtxGxeTVOyrqtqvWfFETt1xaXyJT
eNdzY22yqPkp5DzWkuOQ6FzFy2W3inp+9WwBlhWeyiD0WfKhqn3q5imBfusV
Kavzx9XATwKzzgozi7EZryTics1pdRt5d2vHXqELtnEp5YBlb0neid4kiVrk
HE2txIn1jrF6HGmMt1RV+qY/1HVL8T23qmy7zXbR194/VcHUE/FRb3xwSp7G
CZL5eKdNy1AVSLIESYn2rM3RLLvJ46LO+4M94ODj8b4A0ZcQLIJKjeZFXtSP
IqIZ3LPATedEFF7WH+3UuWAh3tXBKfiRPbxU70qn0m/GrD7933GqIntzkpIs
ZkGiH3VMzXc8aRa3NVT0Socz6V/7SOZ43s6CFQKOyzxLHHIsUt0vSRfnTlk3
C3BoKH0NRZdTcpVRuSbQeNsFTZCf2/VPNyrb3XwU66ygNZ1QXdnAnkxPcJfW
2Op58o8NVLQ85RwUJX/vveuYm4YmS/k4ZqH8QIevumJjWmJou45Y7N9ddGij
HTcl2lQIo2dvlbEOMNU4epIrdUGrcoqupD04Tqg2jL9+Sh9D8z/mLnyzskNn
gw6twf3Wsa+md9ZYfuCpApkSEM4+N2MD/r3GXnZ0bwnGkXll9q3UNGfRzMq4
elVu1GfwpD2Empvo8/srLLZ0ph9rC5ydww9GR/i6/ol7xaj8Fwcbk5ZSEjxM
gFrZcEYpCkl0kB2VkEmsomLo9Meyo37SEbWwFzsJ4gdMHSmBZ2bsEAhoCFSo
YNEa+4yMtfojCsneENiMVui+LsDVMunWQxIauI9D6CQQTq/uEn52ieTQn2aI
RoHUrL1BM/M6UBx9CcoIG/OXj7YzgnDCregGyVaj/vamXd8yxuIzRsedkTK4
si5p92GN5L2H3tyKhLk2xdQ0CNqr0MpJMhjWbFhU252Q5GdVK9JfHIoQ/mL3
VG2z49tMxUE2Sfejl0tBMick7zklX4++tooGovrVgzuUIO7+ZN4eX8ua6S1w
4UcVKUBA0ArpZD29DihA5+oG82StJaZkeSpQfcKb4tRgwqMIZ6cfxDmeKOuK
GHNMF2BXdo/2TPMUmf5kNwX6RSdgFX4ORRJ7NS3QG5M5iPFc7QX2yxFisJBv
0e8DcUjhu/q92F/PTzsFl7YWubKqb1BpxlyRX1o4Iee5MPLwWGx4jROcK3bH
fPXSHyMmiom0pRE9gX0KNguSgYQ6M4dE5ptah7ZUeDOk4H46n++kvOB8sCjX
II+WtQjz0ABWSlbJuRQUtCYEkIZZaLB5+r+czI6HzhPqNeNuMG/N9tnxFHaX
oT+vc3hPxRD/jOkFzAZtFc3FfdrzS1h45nx/7ij8xFc0cpDZWkPQ3KWmL6bF
dm9bep2RaDpoMrq97AFwePRoYVOWOtG/9xyj+MHw1Ktp1/q63xaSlUlxKfqt
uA5ZngDa0ipYpB7pfsD8rjeoKb/WAWG8xYeuSml/Rpke4q3C+SbP/4dBv75s
vJgiJVFKGkJ/lkMXgQVs7oynOMyQPmWCaZEzRQ90DWRx9HvRwPF92cy+t2Bw
9mhQM3mW8MGM6tZ4Kxbw47TuUdNLpXvTJu3J0fCDcEcPI5BTObCoHz6ffU37
6Wmq5m1BqMA1EJa/pJX5fj3dtwwS+Nmcu91HWUu4xgr1z6mtYy8QFexSt5dn
cxNNu606oNKMEbQxI+ObWxXcDoXbZiyaykZtRSSJujdOTfotcFRqA+u0MsEx
dfPpe3b5xn72IPzZD0Wbwd2mYle96LtoSnToqLF9RQw49pgGwDT56xz4B4fN
+E3xZPK+jBNd0QFsCnU3yHIdQx86fmZ0lrCUIgGx3tPdLbzDCS05hQ0HVu1S
b2OdS/93siSvIIbSw1Z0VVEuZvA2Q9Ofq0F39Ytifz0w52vB4mVEVcq0R4Id
ysm32TlQNRe4iU5aNkGeJYEew8q/iFez31/G9EdZxtlQMsxIRKcedy5pIs6S
hx6oQq3w3TJOFSUs+eqXvtY8cvrMZsYvi8bFHZPsraPmqXZX6erVMPsBbK4O
cV6GObHsw9zgNbRUlXMxUoMVQ/28DibkojBKG6O2OVaaP4WO9RgAW1+8ezDP
HWk5oBdZTLbm7kQfRde6BGkJIULPvJRdnl2uaPtNGKlCAElslrMgkzEl25SS
n/vbVVUnjci+L59KeeoVZBuNz1w3oxS3X1mCSvuV1+QGZZwEKKLJhzOt4fD8
Br0tYCzsRKZ/5svO9YkJx2Ka0NXGGMs1x500rdOEbSgIlR5Azk4NSh5+0O8N
y9Ibq9LvsrAoXatqat5K83t/R0PvtDGhbERE5o3hK6N/zNvaK6Ol/jOVh+Bn
0Hpe8o/MvjjJbNDi90pz1bmdsQt8b5uK/pMe77xz+65UkJowvTFZYg0HwjEV
VRcCW/EGvjQBvhdf0y3sRxxKgc3cp+8lMvTfzVNc+fiqvQx5OPR8fYv2xSr1
jMmzHHWN1Z0AnIPk2xjXY/6TBGatup3xib6AzUanaSbn+iJ8aUSCwGppNQED
Gz7/8DUlD5DbBIgEZpaijDiHX3h/T0Qi4ISvYSPSOrfZXzpzpn8gr5Go6wOp
XZuwOkJfPykVd1Ufo6USQoCr2zrQTi0zYVFC1Hfa0yUzB6uIfpRCZquLJ6Q0
U+reVg1ukuIhSLNb6jE8rJhc0nsg/td4gzOcyhAbcSS1L9ZqLl4aJeNkswN7
rEfWJxeIKy+yiIYpIwd5Oxl5LCZPFZx8+n7chBEqLFMksr6CXOlQ8UPC9ufj
Are+hGCkFbReEY8CCEL6C4XuKPsEuFSRtKBDrhQit4JmhA/lqS2u2HD0AtcR
fN0dOpi+wemiTONa0Y5EeccJS2A//Ru9ox0LIGzB+UQv4tlyekppdqgMUZ8d
809QB4p3WDaAq3UCr94Knco+NDzeUxVfRCD8pFTOtckxBW8y3hssZNTdYaGf
PSKHgND+CUDyApmC554Ta+ByM8RVEVqgIJEAo/Xbz0HyFFbFzD0Cwp0ZFev3
Hp+7VtwGHZbVbymjHk3EjKxkNADGCX6jBl6R7hO0+FpIv/PDReGTEh1o03yE
HNhK4RPfp1EhDp3k3DxSE5LHuFuuzhhI12XvGICbkHMaGObBTYT+pHXqSfvb
3mlHSkHS07vGBDQu2wfSKr//dpG8H4m2rEpz9RwclMAwhDBsAlCQ2CE8BK2d
BB7i/XoMRk0CKBiflFSS4cvwwpoiG1Dp0buVuSS2VXbSFu9+p/EZngC66gOa
1jiu8jjXcVsRKYA/BvR4pS7i4zrFW8KAzhZQg+1eHMWMSlij5oDGdqM26LNe
ThKHF26HQyJtpgOv8GbAL924cE2KTua1XC7iFBSTF6HishckXki9n9Il13QV
veLZ5tI1xlzY0cZQpdIBCg11tHFjlDisuX/1ynwEVvi/aQh2JICuKB53GOkm
lqtbJgpEYs34A/VGWo7+013Q3zrWiwJTJwWJYHyrmh4WiiZotW4P7Bv6dfRG
STKojIjm88ye5Uf3vXunmZMhU7bByws21+o34LwZ4BWLCSbcuGkY0fC6X3DB
mFmN+goWDxJ3bYsyMZ45Bl9Qoa8/ijJ7sVJ+feiTp9K8u3rzFeQE7GmVXFC4
NxaeVkPCFGMHX5IbxmgS12DRXIUQGCYyHI3P7To1uj0YhCZKtXvDTLwhQzi1
XpleUm+Fx3pbPc0fL8YTMdOIJq7Ze3kp3BjpOgYkiefEhZ0Yh64I+/CQhGcU
6UzwDgANQJrPPmzAQz8tSpXh3bJFt/qcsfNVRQLS4yxxI7fzMdm3nBtC26pG
wYrx17tIyEc6HrMqdzvNNPPAs+u0A/qQZk1MDDkCn6FPQSvO6Sc5PeuaHaj5
o/+JMzf2tz55WaLhovYC4g5KvSoeH4hzgipJ9AaYMCKVqVt2ajT007Mq1Cw2
0N252y96waFeFdBLJnJTW3QQ9PIEBGyGzX9caUAT5cowYOw/eircvwDERTRB
7GqzbhyCrgWGwqmSBBTfUOYeY/L0Ix8gpec1bE/nzhDb4i6HlmG38Cu1RZVz
fOKoCB2+hpLyq0jfRAQulVSeRM1552BecOGp97OufGJFsKzPn0mBWPFi9XKW
tNjvVN7CCttu/DdE8RI9eJOPOa6S9X3FA4g+fyqDgqxtfnD8aEUCh5Vh6b4c
LTg6cnSZbgH7KJ5/ae6dP0D5ZK9ktuGfWRbXg4XBoje36soGoZuUTAnmKBtd
VGVBW4HN+MdJDliBdCR5zadqPy1NNSOqolwbIaZ1o74ifQdaJvL/RJPL4/ZP
n50aURoenFuoqz12ex6AEl8zCnFgKyN/lqYoSMl+3Vi5oNUrtRee4EHwxs3S
fKwXGaAUQ0gY26HInPtUuDA1r39uSXF9FB41U4m+6vLmcm1FbWOmvn+zAqhG
dAu12HgpSckTmEzI3bdXjho0q2Hv2l71Ug1EMuorJXJmxxwyzDLYVinCjfc2
nci6kL3Vty2TV2dpLbi3GC03Du7AEuECi68poV7J6MSU0QRxfn5m6pG8tP7M
hb56GvpPYFX1fF/BDNUr5zVgJgm/viitDNGcM84NPIs38tc3JvET5R/FdfSs
JqZnXWxLZNf2Y/qmVVK37V9URvCiZAdggUT6CzfirsLQUf/gRME22nceYmfL
Tu3no6T5v3HMxOcpEs1GvuSJpOHr2ZZ2z9FpI9PAX5SCbwAbRPYBKX7ovhdA
dW39HjQrXykpMc1CCHLRfzdFrWlXlD1InJwTmcFLBJELX+JvAJG6fT4eQXFy
QXqi7NWpCMsP7u4V77K34GaFkVH6Up0G5bisDE9FO6AhF0BtoPjrKT5wBJdP
PMgY/fzLelS08yFYBWJ2wlJZm6IJirUyqT5TuQgwO7PcVooNaZ8gJQ28g0ON
ms/gbsIneC0nHmD3sHlO52zA695NWm1KUUtGsHRa1A3kiyB6h2Q7h9S/IjxZ
k8/5PXDr+Sd0koPzu3KTXi2dNBXLSTGGBzJchewdLK1/5LG8FQ/Lfe3qblCK
lz10BvweZR3KKqRop16zZqVJUQ4BIoRqCrlTj2W2c+NE7B6xYOU+dh1lpN8W
RtkrCuVBJhlRpkCNlaVLThbh7KiG29CI2+P3EEN/gJyNYyH3jIo7UR34SQmV
RUeXALYwRXSA4S1GHsf/HyOKS8iPoOI/T7uueYguiUzQan7XED0EgsnGnW/o
Ut97S1kaMkPqVzpmjO5xdAdzGCPB6++V881FTt3K+5L0JF/HFPB4GLJOxcVs
L7rkLUs7rlEJlfeBzldmZRIULbmG3cSGlGVG9o4bnSi/LLa2mHOzehMHal56
mj0BOxZupXpyLOX+7xnwcPwSIkosSalF4Cr/Ck+Dydpm1MhxMZlGtQKDG9cM
050Pdb1GEkD7xLxny7G//w0KXdahEG9bxZLfjHaT2dNuJmla7N5TyNqgTA8x
HzRu+ANaXjHY1enRqGgKo1sUVuNWLfCKeQIOr+tLvoliPSVos3y91nqSjY9J
B4dINFnvEooWZn3XhkZR3XwnOxpWZ3N6jiKtj+2Ki8zPsozJ6sLAg/Ebw5ao
CbYjTHrAudz9u+vxxyk0+cz3kNPdBpr5KjIg0lCV7FiKU7nYG4huqwVavFCx
bhhrbWeP76uyxDBXQoEDsvOdJJnS21pkIVJNpxsUkek8GoZtVGFChXhMbcvC
ipU3l9EE1OhyWxZOA9dhqCXa5btgqZuTohxqkM6HY2PCWtK2+xpDBNm7dJpM
tNkGak1HLKQVGdsECvoHWJ28LFjFLdMkeeDv7Or0lmP5g07hQB6WyLLwqQ2Y
rIrA/giokKK61F1Tja5zFzdOoFExlodKBhJmTErQ38jnFZW1dUcV/IM3wduD
/u0/3Z0KXs09VfcVrksq7aVfFHaC3R2swTG7p77oPA6KmMaU8Rnu7tuZ7v04
n9fpTKSD00OIawVgjQ2vlTBZIsXtsOgP2ck57p+a7IT+1fuxYgpTITdzcBHi
7MLDzmydvCav7qawTX/lbTiBlcNDVWMAjAfG8juqq26h2+PdToRktRhw/1XS
SsOlXcE7zKpkdLzuij5kXlY3kXa0g+0eKkynZJWRcm55CeUei2e/1nzi976k
EIjpSPjOz7GaniDSHXnBJwJunnkPZls1yzZhcLYNaTjEVNnUEfnGNxSbK88R
KaZW2owVny2tmzof2wEkGSud4kugw/YYnrXNccfJv6KfVAJEi2iazvi18gH/
IuBoG9D7iJD+QyRhZbpSNqJyapaot2rdKnwmLxH2D8uCa/8ql8GHYi8uioMd
2QOQ/qEnok3N/1bj/ljBAuEw0a3cWrOYynljrEAtTeL8FxR6/1OTxZRNpiCu
xaGzJWI0Nul8MiKUCwFvpMR78fJp4DnBFrVXV+oPLYBosbjA9eH7g0bvmUvh
94HXK8MQCQPB7PrzSQaYuBOIveHmqfis5lq7L92iNHlgt+YKrgSkUTUlAEjb
PomIPwFdG0QVYHjSWZqhP/88/Fk7uiauxGjbxFDSgF6lW+GA9idRfq4VUtm3
b1vhOR+pN004pwjV1yjSohD4+K/C3QgHoyH+/89cQlv8kU0obi59/dWCdEmh
vepSUEJdlcd9OYA8BjtuZylieewet1nsJudmGrtXAdP7XM4XqdBUSWjih+No
Nmb7AdP8dvywcxcS+2vbnGVl6krdF4fckxqNH9UcqYI9V1L7neQKmgcEPkQF
a1mmDQ6TS4uoDvkFuDAznqPXYbiQYLTPoZEIjwLr3FG9y+aYpvGBT7wOMOfn
MW9jtkNJbkESmunw3UNRBpV4ebV/p7OX9yRHqH2iO2Q/3J3KpSmOZ1Gx9v1T
YSxdl+Ekv+qiDv8tmNLh4j5l2a+lTwZ3sEBKe6Ri9zDu+SsTY5FulcuBXxuc
HmmK4J5COWQqw4NmeO+3wAtDe+K3RYlnEqbCgYi70S6TmUTFCTSNk8PO+0MA
O9n3CsmJlgAHTYJ7RKE5BxXAEc652YeSbU70t2RpeXqEK8vTeY7mdJdv+tiw
OFdmTDE53wNLSQ7Wpwt42RlNo7LnZG1jNVx/DH5Elb5K5ZLC1h2gVdKrePPy
pR/sr3vhaXnft/SZV79LMTydC1HezmnPdpBOcamaTSjZjOVJOfgvLmgyBu+y
O51eIWDA9yC/5fDhxrgZ+rLeIBVcyQ4ndABb1TpuKbksmBxfHtUbD2SBKJSn
Za8Gj1xcxodH48qjENa8Yaa0x3w5216cXkZSFXKu7FU/n6uPwVv+n6O8FazS
3RBYq4Q0VBsGi9MiiS255Xfk0idrRvNJsnRdsh5KP6YymHBAwFxc5jJj0wUJ
PtF8uAt9+jTw+8a5rNCQXQaxlVo1s9ICj0u8iS+FyEVUrsgGBQChfnmiYGy9
yVFjplOL9lAL8aX2Yj2esEu2LLiGNY6Cl7lHspHtm0/vJnKOJ/0Uq3hcDjbw
bRM4tQJ5swC9jH7f4pqavL19J16T+lXp4zGZdAGhJLN+JKNTHHG13wvSPacL
xGHHtKOZ83XGCQLA71C7oBPYoxvSWolFrFqVh2WJdX8xtspgh4/Bj8ZeV0+k
z1jqujV7XVi3YjW3JJ8N/dVuSNdqQN1VKs/LIZ5+t0aCGVND/jNHCFqmtzj8
iV3sKk68ngJP77gmowVftC44D6I7fKfgMlxNtirxmHmWJnlADPYhy+KKjv+7
YR981L6DVMQZ7744K4VmssPuQSX953Fz0NaCkTwCbVbzSiqwT2yxfP+CR8SY
3Qthm+DMT30+PWemejBAHgSR4gCf2jH2XnJ0+SSYvEHPvnXVAxXFqAiUGcQS
6imqJni6q5652OR6w93M/AIwi4J+4RI63817TgVqZQB9A4/86zwN89O6Eu4C
RUmbaUDTs3jBGGdYRbEwYDQGWdoJXjl/FxmVsmf2J2uDoNHRzuZbtvrZgit+
piX8r91JmG6XzHIrAIDv4XvyZgmPPG9Aq6/beI04RT3htHikltRiVoattcOt
gA1TSkwhkp1G6zwRRxJ9WCHXG2hmrSs64oadqyIr4ERr8MtdzPbTII2q7dXJ
uP1ODHmUoXQq0exA2gEviJkzKQ3ubJPKfYHw8spGaY0VT0vzoeBVBIqaiaHV
aZquavnniIlOrF9jwpdtZeLZp14FM7WKSzzETyvtX8Q8c4zOqdjqNyEUKgIS
RH9Z2w6LZjTE+JqV88413GSKw8zoKdtjiG1jodk7xkonPUPwXx0QG1aoPQzy
IHAgGUnBpjFU/l7b8Gq52G9Lli9vblZ8qYfK0xnxY7ll7sX3Q7WV4PU6HKD0
KuC6k9VEG7mYIChAqaE3OzrVLeQ4yAIlsivaP/vpsoPsSNARD7HlCRsu8sfP
De2tj24PlS9VZlmrEr1/SGXTQ8NRVgQS4TtSE47eElO21Dnp7KsPJTm7W28m
hJG7AdPW1wbThTn2ZA5N7mr6+XXsTDpO+s5d9+PXFiTxEHC5dWY0+0bbU82J
ZSNm4jiJ8rKGZhfCBod+wwtTsu4cpnonhceMG6+VCJULJ6KNfJxxSg1hnhbS
s5O4tmO/ppg27VNLCXVca0ALupDaLEsKryeq4sAKdKV0oc9pXUBsJyFjio/p
rtjdXVuxl3ArCDc3Uongx6nqx37g0DjCsiTYpBYFqtoeOLZyz9qa+Wq+paBn
LwFviKNDYSR1H8qpBVM08RRgz799jZ+0Alq9OosLxSs0XQTqVL0I54oz3fmV
xCcX5a6V1iljkSkrM6L/k8cO5E2/Xg2/bbK13u/DYoAwXp/BR/M3q+Xdo5Fx
7VPbXNj3lPP8EvBxghE0i3iyv0PdERG0MUPoT3yhtxJoLIwWyqsdGr/PG7Ki
HLLfgjdLHfKjIOAcPtfPKE16i9I0u+h6wehqSSfrVRi66ZcJQdzSmrcgjn3O
avtheBL2uRdRiPs94IoXmQq7u0E1A8jrRcCrgs99fdzeTJU9VvFi5K3OGtKc
I+eRG02ueMpZy/BIFzG4uaZMNxEzMZYGIG122oWm5i8JQfRB8QR2zH28P0hD
Y2YHZUVljc2h0njIBxfo+bsTsKbyeR7FDfPU57cudUZuQWeyG4Sb3VK4ScI1
fLT9lFNZlk7cXNIxLOO6E3D0+LcDtHYMqKcTlIDz7UrYUkIyqdeHMZ7ceZ7a
lsCZFkjcwps6c3RNS6SICO+4c3/9rEFDGGb+VsPMy/9eGXT3tDXmksH0hN5j
IP03ERP1pK1Youo5scxUv3/hvx4JDzn9sPqi3tZheGCGNXLEVijawXdoxP4W
eI5Q/mDbRELgvBV2YDD1ZXvHYOy02R0EdNQKP23aFWZvQTmKRzaycdybil/J
j9UlKp8hC41H0F83h/psPqdAVZJ3bbCBbSCHAlJmfkHfWa2miwc8fxh0Wj4q
ZOQusA/jQ6o7RWy730MYKo7dNwN+mCJSDJg4uKxei0kRl0J5kPWXtQzhJEXj
iqwsXuEr6LBN0L8gNyhGVLFPaPZpfnor1o5v7Xexw/ycBbAj2Hw+5bCUqQd8
cUsRCyo+PiSzkQ7h+7W7bNp+A5xTwHAxuEOEp3y5rIdo8Qk3KT+VZLN1bpgq
vtU95Mnyhyq0N88zN3+4UNxDvY0uciqKCUJGP6fkVMTeZRwIX7lQ8op9b4g5
GkikdgjYgo/I3ZjdSVH/8Bbx3Vqc5s2RtjS6+n+LqJ5wpnlxH08T2aMv5Y0x
RSHZRxl01Lk8nrKBLbP4cJYyfaQ3sdeRL2xlnmfwsuGhxrho7iI4E+l2dmS/
WaFpScumEUD6dg/6lOfK9RdAzaNo5ziMSME2PYSFzYiYaCm1D1rDvPADEkwg
3s0cd5TlPQVhgKwoat4yo8iqcWgWEsrBQxjscARAu2JNkJZSXuXb9ANXdr3U
HA/IH/p3S2dItJOhjXPdb/wxQ52fjytOqHhxDte99vzn25tpAYBG9Z78oLEz
nJk3609lmHpo5MXZdwaxboACFkMtbDPnMuqCDKOlosYi08kiHoyFMVNrfF2c
xB77PskJCtXJ86wQA5VlnCOPOpvSZphAv7ax5KaFkT+RQPB2xYX6R5QjpJAK
E9E906a8psjtKIxxOjcHeAXLHJUxfMoqORw3DdPeecq7S6mnHDIF7T4KUx+z
fhR4ny4q3hSY0yxqVfESJo6QR6OpjJGPO0r0BaleDbbwrXzAxkLRjSuDHIzx
vGXbjFHD1gMLLKUx4DNo2er7ajsuFtFT226iD+EdDLuv14mfpmdeo1EQJhy6
5hCB0oapHSku/E5KzYASRtrLYvtXMUdTjOMHxfSfW0gxLNoJpIHdJSurisSP
3EI6TU1hiK39ZWb+wlxahkSWfVVa/sU0ZpGeRAtHN7LKtEIbqP0iaMs1bu/R
HFpBjEp6rtgbvFN5SA/fIGpH++tm/WB+YYUdrZyPqlB+IrXkvJQlmCBr754R
9EcEY10z4uG+PnQDebgojGxIVF+4SYoKq31vzrrwJrBNZqnuqsvyYpscZ5pb
eK2Yu7t0LApMHZJ4dj1mZvBFRTf5xcBSf4EH5MlV+1fQ/Q/NQn9N465j39et
sP4TRZlUWxhHrsGsR+W4EP5QRm8wUEEG2SNralNBQ2TDLAs4nR2OOViGCTjW
jikzUzNFZVzFqtNpYEdPNdvHAwI3nUIYZy2oSGBOXxvrexvD54aJMZahaJ9s
cADrbBIjpqh/6P0f4bUoYurVjuBSrPjFsctB2Y5sL+xN+HKIpO7X24swPehz
C86GT60J82m2+89aYMt7Zgx2ZbjqDWwiWPAXDnOTlcih4CvGkTZXZIMCxrBu
nJ7L+J8o0FV1NTShrbTu+epMUyc14axF+hQATL2EyYWk3r7pCZkxSz6E8sW2
MJwUlvc0St+VBIWb/cFxsgu4oae9uhYH9HeEYP+kmxsRsW6EsqvILzQHUEMT
Mst8jNAGxScdVySeNL3ildwA/Mgn7tqfl0XW/bidzIEeVhH+LGfTGHc4AEYq
KVan4bzqhNnOsiRnNpHtp57txHSHqgAyutwQ4y/xp9zzBl5BNu+cfZ61e6uF
AuF24ntoDLA3a/KzAYyXaLUxxHC9AkxOMBbx3N3yCoDW96+NxU/jp5WGbERt
Gf0v895JLSZ8S6+c8BzZKNr9rPg3OEQEBP3eZ48+qTwhIx+6hwiV7TTvng0L
dCBDG7qOQpvhnNhU2G+Wbh4eXzuw9CJVlFpuxbSPVrpxf8W9FymbnMXqPuzZ
UU4XrBWcGrm3grFK1lNinzpOtRHnwVE1WpEVvu1c5tL2n6UYkQ/x2wwGNieb
zDhZMzs4uGlwB7L5A/j5chRbNsdGYcEVMpljjRGL6MdCEoKxThm1aaBEs2Ti
zJa5UEfclbMeXXCOk9MHzn0xVwbutksOECWya5AtgA8bvmMy+ZuUgWX72L+w
6yAHsURIejLiJp68+u4oUMr7ByxX58/9azIrYAHq+Q8ncNDrEoZB8DcOHSfu
07I/WpV1Cpw3D+mYhCnyhRAzEAk+pOx+rlQ/uMfgtLlXBCJjo5Uqj3VnxvX1
FWDMICifOakU7HMUUbfMGDmyH0ffBMrqksquw4CXPoywzPFAcgRXfVzvWDhB
DXrVeBVFH0TSjcLYtjYJUMLXEWb52PZiO57IKuU/cOowPEOFM2Avcdmw9zgQ
H0zrlhZ22TM0W1WLQUWZ6McsJONTQ8NqHw6SpA5lAOxm5ka9lCOhFMsTGj+C
a5c1BsK9I4Bf0Zm6uqkq8qejdyereSiKYgr06kpr6GJNnGTDdMu5MxFMVKxG
PKSKszgyUH9FqE5q7k+8JL/Ow8HnW8J3q0RISj9F37uy09Cm/kIhbE1KULl7
JJSBaXyJZTft4l6U7ODoZuDhjDensq+I7t0wGzrFLClG4/wo65RqhP/GGpwU
I9z7CIc/WplYKrS2GYm/yHMSBE34SA+hupjMBB9cXsOEOGZCka7DgaroLGlR
+ytnO6Oz/LpyJQB0o9rE9may0EaVudfAJvLDLctsYdT4KcHY4A4+pbhVnGLg
z9o5KhXnyjHbr38Z4JCgvzjC0HjNMpwsePntmftommdUih4Bu7IVYg/QqNri
nR+Oci0dcIqbY2lvv9gI4TKw5PsPen/NkStlyfQ9XIhGnrX5f63pgxLN7ZoN
JhJVvuOM2zF9Y7z8YqDYcyAuc9ERfLGLPzlvtNyMnDCLEo0Pzm6uPx9EH+BO
4jtVPcJBxe3RjKENNV4KZWXeCWSXOHT9qM1krqH4hJMRLttOGmb2ItPKlSEW
jEMChSIT45wDoVr5s6gAGp+vaTMKksnyQRbbf9Y/qogPCnelrR4joevCK0I6
Pnl1/yeonS6nPFg8kcb6P65tZTAbOQ8HnKvS9i+2VrL+NvmByYffJiaeMZRK
vfISnfqLSGRkXm+YVxyMpStotN8ksk3TJD+K0sqhEPjKIdTveyJVrsUaaw9O
wxV/nw0KqUIlNOuR2QfO2Ml3SUZxhsJPh5im4lrxjrH6TKLsAFkaeu07oGcn
DshHdbr4yztmxGmz6rie/OgkkCAigo6JXEL84/ga8T7h7NDoNFlXpbDMIumi
rGh+5d+cam/9kdewZDt1MgzlCNRhnJ61xe8sVdv9Cn83U5A2i+ptlsAYADoN
mjSj/MGRV0SZTWoiAR7+bZ/VbXnvhDqd4VsofO0G1YCGtYdfn/78tvf6bSqE
1gwWs8uqSIkFY2eREDUaVlJAVCGmaslRUaXNXFGehGqLpMS0eh5PPPB4IGop
OfhYYdAeLiktv6m8x6x0nYAOA2MkuRq4rvdaSXYktDKhd/Vu5mdwZMVgvfEk
mrap3ZSq+Z9RPcNyC/2Se+PwfMgI7rJbrxDQGKP3v82155rN+hXHlHOo4FAw
dqyFaZH4ddvRCWBQKIv6i1Ev+YNYBCG8T5Mqi99Dv553BfruZHPP69Wsl9UY
FSpUJXhz44SL7hvSQor5WH4dZpMuVhJShOllhFQv7lCuJl0+AEtcTAko22j9
/o/b0GqloeEj18PPJTpcoqDfntIw4YhH4aACxunxGGycVD04YIoHHFe2bDgp
Yj1+akMaaQ4QT3jM+lP2/i+SAWiM3HWbZjO3LVlyxGx7vnJguLN5w9MsvAxa
ZdNORa7mcfYTHHE26fS+hK6ccC7d0B3+xe9/ukOPvHGkq7mhFmA+WhyvQ6E+
rdVDchfy/QhkT8VoH59mxkahE+cMMH7gUu4M2VN5DrdQX3i3tiKkjpS1f+Gj
6o3HSVhRHnjCsYZH8KDz21BiUAvVjSXpHbmsZI/qoo/qhLI941nPJDG4K5YD
6pQ/QqbiqCgdE6rXXyLglLDD08mZ56P3AZ3sIKRLYZq4K9cHKxw953hdMmXb
mwCj1OZGmmhAOeH8awtFf4wM2jf+wyjOBucp2cWpgLseKaoC+nN7GsiuMNaJ
PJ46JyNc5X44OxemlZYAoMiDV4CqmW91xzFGu/FK5OC7B/KF5z9OLWIFYVmR
PxYoI25IoRPMr1ihdKmF3HyDUOG3jWMwXUOKFQhY1c47SETOk4AKgt2YQ25Q
IzpRQTzth3oaJWqAbLA4Z4s5QVZzEQBkbnoKEDwSy7UFr6TfM0WYsvvjZYVx
J43OHlHQ2e0a50nFu+EqFaGLY7CyNfX9z2RqQu2+Kr0/GSl1yQCu6FrFgj0s
/MbOWmwKYu6fXBXxkTx4hn4+QPDWRuAt0qLq26l8Gf766+NbvsvpELkS7N7l
KlWyN+HOwrNZo8EGGTAeXq2cpVHwPKKvX9ACarJYllVnxsFn7U5Gw718wjSt
qR5fBQvhK8O3uixzheS+5btKccidNx9fM58UyUHDpVkqqFxXrdfNvSB7zUjx
NJzc4+5jkbcDLjm8ro0fUxJ3Vux88Oi1E+RZAs5ZtGQ5kaIuAEkoP9ATaf0a
qhZ0WhRcXWllCWK4ehDw8iJev9bUTEHq3OdwxohYmhb070TJAJGOLchFBj/3
Q0G14xY/c9HHqlOS5IiE2ghHgTwvwTWh2bl2N+qQ2ZyZxHTFLGA+VAoRieu7
Gt1GE2QtZ7H1a1Lx4+yBDa/aY4XXm5tHPKvvbmsdoNkvaSVC9QCnFVx6cX71
6Q28I1DdxikZ21T6vMKj0SYV7P31Et1pzkm6e6KXA/eYrM/O63wvAoZH56jY
aa1KiN6GP4A1EBTi5IkuwDgoq91JgaTTLaZ29Wpf0j/J3k8QGWoNzoBpYTxQ
jmA/fSZ0ev5IqzvZyDjlHAHU9bHEMYFXY6LugX265PWfIph8WRET6Nlyhp8s
2BeDZKrjPGV77dnBxnCIXIAP7lwYPr47rl2cwvW6W6HiW31nWhlkS92/7yyp
8V/gcxTJ8S6QbA8oOo6USC8jzmmq51ppAWZ4ynh8YPnvBLipJSPVFTutiG8e
HSERRkBdTWH8VKEwSDqOt5ThhrxeXtON5aS3IelZ5UxTTHuicqsII+5JsWrs
xHTs6LHioCn/U44beevNkg9YooTRocr2d5VzCuyQjqBpbpj3PDfBEkqYoKzw
SgPaPzUmsRAytG5fPIuE97GCeQXg/hpq6Tdqx7u2edwQMToLxlQGz0yHNMgX
ZUZkhJaovXh0ccnDiTVjcSPUqMAWhcKeN09/o26QBzmrHe9YT4COznHET7Jw
RNojMOudgvwQ7b6EQqh25g/SXUX+2CygqcU8/fpjEsKEbn1+fBsgx7m1WKSv
mkEIYApaRGuUngwor2IYyUS9jVCSeMyEfYmBnJXe3QonRuBAVdtbB6t8hYZt
Wz3YPUuZW0c4Bea089/uGaX6Jfpz1hwtwEbwEd/OvHaQWJNW4VFsrIy2mYAL
FBJLDcK/ClK4sDssZUZSeVjjrwMQ7anSRXC+7dlKy8rclOB0eGr5LBKrsLLu
eFu6hh+66kbIyp1g5BNS0m9pRj9AhHTFvmfpDPqQp/4xuroKe0sGny0gQp+h
2X36DpjOYYKB+oR2rTlRXqSQ2M11bqA+2ZVkieSZuRg8JZDjN9vhJXKbJ9Hi
ZZkJiWvZznGS/El50an8BzZU3AkybSaDbKYtyrgGY6YujYinM4HZiMPEUM3V
WcgSjcHjqGJJpneMgTv2oPZ+tfVGngt4vvDzMwPrxXSa2zHt+H5E7Mqzf1bs
ZA9t+IB4PUmjgS9OeM51XgE+HGzkwF123gH2iQLxtz6TPQfwt3TJ4e8nebDK
p89E0eRKZfqeCpAmuToc2P4fs6O05bEARmsh7Nagx97JHZFXGUodBNqdpe6i
fy5YleLtpE/rV5hAe2ixlneLHcgQYZJJuY0A7Jj5XBuynU/QCsiVsOC4dN5R
y76r3xxh3ViZTe5HMbGrKYAwlMzcYoSQjpSJkWYZaHkzDqSg6nizxLiv+Yc6
pVVbzBNpwhWekTH9sYiHi+81HMCgzquD2676A2N3DvCPulP/TvLJM7h7Ya3p
Vk1QyfYtOIWf7vfBg8LV+QyHH+ftA65Xrl8TETayjgMUkoFoHH6EG7RZWGqy
XOHR/jPqNyetW4OVe/kew1cHwbrW4hQnMHBCx5WwOzmwojI9bb+3vhAh6Ki4
YdCVmK2+0PlQb2tLkV15ySK6B7trmfag5/u/LHABLy4tYSJ+6VhLarFskl3Q
3V2ek4IOW+s9bUrH3DbkgedslJE/EJjluHicsQnTOhp1zBO5Zt3Jqe6QG8sJ
tqbA90uxPeoTMSYud9vTP0atzSMyVeazoTHIVRDdqjnfdGAYIslluWDZIZUa
BkguZImlMz1Nn/61vOZp0XVUAQ5KryEVYDLsJzWtKK5e98vHon8W8rzDj8IT
7fX+6/EwaxwxNnDXOKJhxfV3NeL2vdIIXSveZl6P3riDpiGe/1An9Dh4R4/u
tvM+sZ5YXR3C69AEqfMpu6jtL6E2FDAijCnltg5b7EncdO5fGvzOfRkGu8tl
/Ve9nM07t/i+lnF85mSXM+khL0hBtLbF9ukCh4Z3hbB0zqGZoqdAFtIDj7JJ
LKxdQyvpvVxr46NLvwCrjwcL3d8sEGVOGCOq16i9hlLq72ox766IdIRDQ0Hi
HhRNbVBDxQdP6d53PuFp3sS59XgUHLQEdsE7jefEXHOTI8CkyeJsu2nHbI7+
/sQjHrWV8juMfHHjPToBB7s/COqSMSxek1C5bCGSZIcBztKO8ehlPVGitq+W
puGpGP6u9X4AGtTW0I5sc0puym4ebUlXCFEw9Rh9YS/4IZaGGr7BLTlundHj
khK7rmmDk8NtWN1YhRR6wbUmV/g8cjkW1brJlIaCeI2q9b1uiaFOyCQcU3xo
1baSJsuthGNdPIiZ/0/XrH/DSQgRk8nDYQy1LeccvfimCMWn6PQQu8k0CiUt
v1Alnj1CeIz43BwcttYvqnRlSyT3XM0+oaTN9O+f9/OthMtwopvX0zNHs4g6
1TG7wChBlOHGpNckrLyCWfCZtMXaaHGv89BHz/iMpmZbDSMg4HP5IbnSU15P
BA/9qjwHi/iFN3fG7tTzj1EmNq9uyLEBT2f2rVbGdy92wmzpLHeDb2udnXHf
OYUv3fWG/APIP3HacJ/eefbGfZQEX0lq62wZ3L9BPFBczly1Cogdj6PORwlA
0F4cS7xzkMpd0hVArlFg31AjIsh1pxjsqpQLPaLfIVVZqHX0uUDc2RaHpdeX
EIFc1F1l07mUez+fbtV2r+7Jo5UOVGkz/4w1JHXjmiKGAbQsh5Syz2uuci24
goRnV56kQXQEo2Suhtdsw//qdZSwL9ppsQH5olGsBt37jTxZu2u7AZLgSYqH
dd9TnVSese2S/re04g6wurkg0TQJWaO74E2PHQhgpFcStGrrEf5q6fko0OIa
N79iDzj6Kx5uOHzzYLmXACj79RiP5Nk0QS9ohigdZRST0Oz12XtUXxvk1EQC
08ceLeMf3yws5gTCcz7nVn4V7lBZct9GlmpnXEMIKzoZORMX4IPIOi4GyDq3
w9dNOj7skATEJ2rWdFV9tiKIEFJVRAd/ISJEKZgXH/l5OU4Rzx0sphxsPrgX
o2ho4vmx62kXdek2C5+IlMO4vmqaftiQJ4tVLXQLI+YXNeWBucu+WCuCGEiP
Aa4LCdlF8l0RS9SoXrtEwoBnoBwHSGGBH+I4ZW+RKIJysWvrKTopeb5Mm0Yv
PcGF0RlOyYj3TEjRspXr9Zzkzf6xXolsoCDjTH8JcTEmOCShBQHkGzr+a1jX
KqcOu3KhLZ6Q0yInDR8H+TBdfH5xjwu2zD88XfJCtYaXxEAtz5FPhTjBkS9Y
6gZz+C4FbaC7JDXtS1GF+q2NNmPNRDyJWe7hk7T2d6GLGa/LDA+wdxhXTu8+
I51G9gY7FOC6H+3ElBnCHeomnB5xiIagwhptJEUtPaC0UdY9mro/5vUlgtzD
dUMiNz/xs3nTXHYTIShiJkGJuq4TIuGeLYNIXO+z4/hEvHnPJVVk6sSPCz4t
zQ5CvqgvebSijfp+J6sQeVn7++Hl5M0HRJlGlyBeXVhUcEaF3Tqx5TbDgRzp
+GRW2jTHFcJii+hw386l9BoXCyvut7qDW5NmaVQlR0qPr7ABT75byQZ9DliX
6bVnXNFwMraan1Qktr8YeTDFhN6vS9Kx4Q7inoT8PSEUoELQH4XtBIE45aCr
Bef6i0au1jFNCkl/B+FzJsJUSk2F1QPi26TkukJEZz+gph80ivkcTCYrQTNi
371QCLOG2Jbf0DJ0Y4sR2L9ZhhtTC3RtQmtmpYZaiFD6P3lFXGwmbFYbRk4k
dkyZh0OnQX1Zkv0KE+kP48u16BMl3OA0VdMv5hXyGD2dsXWSM17gltYFrxxq
jRJlW87wQY7ZhpsrC1vn1Y+VeLU3BZXtL4D8l2XBWYVBscHrvwH2TO9uRHwE
g/tgDDImMRT7BJi1ZRTOEQ5/gqZwUOKg5VsOEnHYv2++nc47W6wd4AQwC5Gt
esJw43REp6STm5e7jYtzxOGHq7wN0KQlxS6wmQi4B6u2FbTUuUq+5K9Ql+nL
drnn0vZDozHaiW6+231TX9qFy+9tK6kK5AwYZq2kAANQOKfdi3wXYcXrSnzu
rnH/yzWALZ5aMzA7oJlTtxZASfmpo13m0ub0IRbLX5gK6xcp/QefSqvJpVZt
ckGAs43WSL/wa3Jen9Wf9TcpI2UD86gvEmK1UouFSw4o3oV89OYlNE8ZQ5sw
ZCOuyPiulC+N64l7VulgeZtO95k6m6+NofBqWNlPiYXrTK4auZAp4zfybhht
XzY+3POWPtX3+hJcedvV0T0/qfE+OqhIr1o0xRPsF3uqM35rLHwPurKWfovI
uqAocRcKSYAlhVoqpUdz6BBZp9LWahrIwzrCbaTrqhq3jpSYgeMZTFHa/GGa
FVaDF7reWaudqHUKtJ0ZPx4iJvaN3lhQMiM1wHMgSPOrz9LrXfNPY/EMMPwT
wSIrVXz+TVQgwV+SIzC8LaLKyEKwDk4AOjPrfThhLtLVWleC4bmCuSc5vAqw
BFFXte3xlMBbne0sdyNGJj5tfVjp/6zdqsgJuR9VOYcCocs6c7vwhN8KKYZ1
yNXecaZPqvErQG1364pajW9ZRhyl2zqecqkdwAU6oR9BggunWNTooAECFeLE
bh3ZyazQnyaz/A6lSBok0CgpFDrxtTJ1WQ8sifS0WwTbLABXoho0LeCXMxBA
r6wOU56b7rPRoX7j5rTQSFxiBTBDjuoGn8QGqmRbbCVmVRZDTTEriAdgKEUT
KUhqP82Nl2YhWKUBhkuAsnH5TDvy5HKR5oNb5YR9Jr4oPnB8MJpF9Oj6JNpp
BuCaZ/wrOETJ2wJcQK3xEkFBiExfwngZoRiQYt57Dlqq/I8MKBVM1C6tdodW
U1VURFOq6dReOxcbqoedRMFzKozHbBnhC8JO6ih9AxD06wc0DnObfrVS0kzS
TdcpEMbtdp9sWTSOLwliFgdN1qj0YEpNujCAtgxJGExXmTGabQtFcrNAznxt
oYxM0AFIrv0A013s2EETAlu19oWodH4n5YDxHBX6qB8VsCeAwyhuRn2N7Swi
tKiMOKKlwmUHkb5aDhA8HTZ6PtxvuBzY0bmvkqbf0zABQIB22rUUK0H+uACp
Y9f4dSqSSQ5W/GLmefvWNRm9S0ZdE4b5cGQbBD45oS9jmuZ2bnWhQf9kDCYt
jxkjABBeAcZTSOXZ6KA/MsCrrXvJ4BnQTMVPJIAo6PpQAf/gDAz0CC4vN+55
yQLl/l8Mmi7B2GtF5bRIoW6wsJfHYH34ZQ2S5dlIlMylR8zzfctiSAco+bHC
a4/Y2gunr0mlunSWQyHn6llpv1SFB8QcVLifohmBb/i58/DrvZ1a0Te+VD47
6t1EXEivNLKEkqbNFsNe3MgRtGjnQ7N0W/GidODuzdXfV8eJY8miPeWSsl5b
RBkGcUC3WN0JKZErSpbP1YkIV1XuUXhHvI3RwaudUN1iqELk9jTmvSFXB254
uIeKttiNm2j/J9gOiGciXcgSOwByONuhffMgrAHq4Md0P2wcvt7vXfb0QlJX
loC2KGk9HMWXsaxLmxBPdOZr8eg6R9/PJrDFQsc3JT9lQam4lrY9sXeyh8iV
6lr22MHKvJy5GlSpgfnkq7iwOJ2qV9feudNZUx7O4HQ9D+mKB3XHL/ev9ZiP
LUkfIwY29rY3WxjZX7TT9rKbwq9rz4Y6KqYCGMr87elxwS0RrydTAmrRUIJA
wqGVpfZHCPYQgqWSqWWjQnsyC410OTbJT+H09E/9m0DM/aKJ+qnZ4ByRmPn7
j99NxXsRwlS8U3q4G3rIcDAyTG9QzFCFZEZvJdRD8ZCUCM6wA+BNKAoAcZDy
iB2ADzfhnKkCRMOw/jAmOLsJ9/gsO37NnN2hffYgBQwkTKc64F644WGcYpah
TiIYRvbvU82rX4NSpZd6jNCi/VNnh5JVb2UQtzeew4Y5WsDbZ/ON0ZrDoeyp
H23tj7z80FcrNngdagvisZI3ShbjfzAucRfg7RDjPKNpyfeisATA4OuEGEtf
hAqFpIHSoosXn+K6kP+hRIxOeTbR1lgNTfxFVKwq69QF/Qgdy4qXqgYA6ItX
kuZHSRWeVi2SY8OLS3fOoKMjgLEZkC2EMfiMYKMyYJwVKAVstG6mkvHFSc9Q
dU96tF4/uT6sD0SpRWxXGOR9WLnj5BMJRqabIFDi7XBIx6/Tp9tNNz3VPBn4
pAWQ8Cs1f8/endMHKWq+DG6HhRvVtCV7RLiJxm1TDhKrBtFHkrOBh2I6C/Xq
qBtKXqoXJwxWKlGGEK9fi3r9uAKgm+LrQyAJ88W4oPf/Io98fa0sIhLm+eVb
iVpyoakqQyNFwJEbC9MLH7k1V1zi7JeXI0RaKVeLsNjkwRxcE38SQuswWXeg
aqGV9mrnUhvNwSiOmUapN3JZYs72Fox+4JaelxnScsNY/orBbvtxsPcwlO6g
uejtfD/DxPF9F4TIn8TLfQ8l885rz+SBMqWQ+1CwlCi+EAme2xOMAAHYC8tA
CrQSBCX94GMkPI3CB4I/q/H8XBCGDxkFcOzRb1OtoqV11ksONCkAktqbIOk9
CP4t92OMUV2+FLliUrELIvvN0ZmjFWNyRYkw/7aPRx5+vNKqDd4paCLGWEmj
9zDvdC4dH4GEDIblHgjt02GxGup2vbxyf6WOHwy2OVqRBMC34on9Hn3RNrDT
JO3vW0nlfOr3vWD0PBqDtP+IEWuC2PwCVbaJ8HVwZq3SWpSlPT/IAXXnXTvL
60YWZ3ea1xjHRp/43hYXnyCgZSSWj9I+WVq/jeGTwnsLh7AGp03aYJeQdsUH
vWvUrxMGq/8tqRpbNtYPjg6G0tiyENCQvJVN7Uc3cI1eLRymr+w8xXqUaNK+
2JoCfIETs6ewcY21C3yBaBqDJw4nk552gMN51JLcr7JSd5QjEEiIga685oYm
kFyMQQ8V9mch3h2Li+K9n0/djFFpGNOmheTqgtB2+OmSKe3xU8a79Hr8WMBj
16xw3uqGT36uwAEPgB2wLASrtyJCwzgQbxU5VR1m89RQw4NCglz8c9hW2tmK
l/VpxjJyGoFot3KT92J8JT3ELOgktLaH2xTAPobcmr3K5VtGxYI8JivVDtwf
0y+xLG2VA21GSPuNDlCIkQKvfgfBUjD6nOTswQ5q7QgnNxF78b8iwpjx49qF
zLOpFAZ9nvgeq9OdQu4rwWGgTRIe0enK7/zTEGloyO1tiLPnD5GkwF+139VJ
2kpjoNcpFmVZL1vh5IvVQeQRrMwb3ocFhqU6/rN7NYWGb29JhLB+t0ORRs5k
VNQMRMgAbxmAkElH6hpJYh9k0N+KS9OqTNDkp72fSYo21yifJMi6UCraaEBF
9aJoWEmRpOpYnYcE1KOsTdCOei0nOu7uKaiXt3TKtRciz1+FaqahrANxNv1c
ysBAOZS3l5kAjPimE8Jnm7Ptz8QBYi5nWm/jF3v+3CLDl4oilAfIhezK2jrO
A0/9BgEMvMsTZC+BhUMU6JGQVo6C0iRuOnMEIukMEFjLdhDAv1ND8IV3+nJU
6z5u1OgR2sTBy1RdMiiuxGxrypGG4AXovcD4/0/xJDzcwPdb10JsbJVh18vS
7EGacubJRLi27Lbuu12HQJeIbAmakb1C7uSU2A+34XmzMagg41nPpIrRlZpi
rmqemSa+G5cwJXXSbFyl4N3Eq8SKKhXEiKhOa5LVih5dIq/2QjfERE7nFYzH
nddKYwbsPXLImGBWXxeEM1MepgyAzJpAC5Rm5h7cTdDV589qVesXMTZyU43a
82Q/JSifE4osPVqj03gN3LCe0jyY67l7gM9ZtiQfcdgUTXA8hh8lCAazI45o
SPYusG0+f3h/Scjn7TkkYyk/9bJdWBG+2Bw4l3q6+5NQVEKzv+zJWUG6VVr8
VWNgRnlsfqR6OL+N+fm0A/vSbqljVVPo5/27JxuaU/F3QzJEUXUegb7h0cZ+
ctI+W6/klaIoj66+t3Na3ur75EOFcok4KLXGTtAUVCeC01ew6b5KQKVP/dZu
yyUwE+6YZ23heGHxL3B80yDzNC1L6AZab6BgXNtwSZFQR5WtqFNIQb4P85cv
qE0VdPrzGCX5+NYNoLDpKSY7wQpITupQCrHCez/cQTq3V3nMFG2eCuHWeHqS
wx3sMSWnahXyDEJwyjWJzHwnhY2M8zMOjQiuOVX91TLDa7cQVcnwLCL6mi/d
TzOT1oSQh2tUqI3JsMeHPSx8T+dsSSv9feotWAjqaQ5WbyKAk68KnGHAUapf
JgU2Kl5W0tgFwV0gbnhWxu1q1m3VGxJhw6g3uIuqIeyZQ7YaYk8lYtG4OsC6
7mIa9RHzelY9oxH3ZlKN7K4m8cT6DGqc+m2+Pvxl8bq5Yl9lAY6ezsTeR/pp
SAWpOoawSVLEbAS4FjQxacSMb5+97/jYda4GEdUkXFKtNfpK899KvRoT9I7S
1JeZC+AsUOCoKNzUNLto6hQyUAaWqGL7CI13BQNDFAfwWeLmGK2ffKhzm44j
v4+INGhc1sHTPqz5I7Ss8Do0o7JhHFoVzNIigzr1sX56tdkehw9H/XoQT+z2
jL+zxvWmRrbn1aG8qCnn3KSB2sIkSp6kTnW68ySxKMhiVwzNMLZ3d68lcCGu
gMZoh28lnIoFl4PIHa9Dvu2KTP2C0/bqqCtuatrZrZB/HdepJ0hTAkr7ASuc
dRhmOmUkgB4+AY8BP0zQqoTsPolFXFXo1QApzCqgC4yOIVy6b8zOtwR8Kf63
mitnfFe4ubOgY3G25Rx/XhZjm9GsPvgwDueHUmZgzv+sHrHlEY14wT2HMnXR
2aAlcDiJbenq7d7+KQmml81hexy5M2hbjbSRGJrq2oCEi2+zt3YDZV+dh7CD
xvDJIWuF06jzczdRp/8K2ng0rOKc5F3RAM+i7T9IxbJzU6tD0iqeYan+Uqn0
dSQuLkrJOSPgsgDHRpl1l3Fd61u7scFCt6yS2hoGPal0Bh2yFYh5deshz76m
JsT3VGESm3NaTDFKO+r8ram8ujb5ZVsFayhODtCjKwItQhpeAh2FJeIacAQn
883zpwLAAU+p3yNK5K4fY4557NWUarbZvEWu9TJJWj9yZnz0Ba0WRJzBi0Yc
Wy/rrcOcXzGd19kac1T03NmxEji4LHVgNjb0yZAFe5hESAqvytTwh9WVHr0y
2VT38xCf+o9DHOe6YOSsGGrMg7Db7uZNRIiIVVeOiAOet3WCEoVG1BFp2cEg
6K0CfJoRSuFGdp6DMml2JRjHvuwPh0Assqqurlf9qUnlOFrprONF7k1+PoSs
59mAmyMHgn5OX71ibz0+xVvjTgfPTaekngaivYuc3O66029cBo72dCK1KpDk
1juaWvxn4q29mqv2Cmem5dpJeRul6Temy08yaAhr3N4muLwxZMSboR7Q9/o/
wTEGhSAE8Bc1g9Wn7FcHa1Hju4u9g+zflKmmcNwpRY9gwr78bPoIOXV0ft2C
ifMLd5fFdq2adAlSPh8BUgy+Lsq2xgE55xqHfOJlksQLk9ToQKsBWRGOJfbe
xmm43Lq5SCRQlNRJnqgUrA4Lt/eRAR9efHXudU08U6u2MdBTNXPgNfIXTsm8
eAWlgGoVc9pHXCek4SnruSTQi9AKli1FyfnSkyvqtLpKjuAJ+2z9tpNLAOd9
6FvrSGCeLE+7bCZJ+uAJQ2S3jhkSltDaihMMDKT5DyWdrp/4QSiB38vk6mxu
VrbcI/vazwSUwe9UR5AZ3tUVBZ0yS/ZTGBWsBrh7EGy7VrZhxw6HGAk//lYn
cVuhu1WcNjVj64/RxBONmpPOqwHXUhHoiaWpFsG0GN4V2uw1+jfUTE3MwCFV
4OaCGQMX3RRbdPmdOVUaCdTbp/IWi6OhODfBGeIO38vl/Z02iWVPrgQhO8QJ
eNMtps60hF0zqtEV6gFNqKuE5D4NTpx5/y6CB1sOGhLh34g2XQQXfJ7IFanr
/tlJQHx7GpD4aw2lCF68iTsBeknGfcUGeifNnUyX7wqlHCVCT8Ow+immPIcq
fjktsWE8oXBF8zHEDEivYIuLTLRrWWDNfQ3sh+9Q1veF0NVAsBl1NC/1Totw
nUj6WfwnAgjo5kpED4pcQ/hPFEB3RSNcPJb5gdCpYL4lADSg26BpPuYMNo16
JlbjC3y7RLn75TIuURva46kbGWqqNSX16IOgk6NxiWJtH+zOMb2/yChbDCAN
pbCfBLTLZAwh0LReOSQnsymbB0uf2+NLejgjo/bvYE+jk953oL3gP+vQ2AYY
vBU0biU/IytSSTBQ+ZZoPwT3rnHalGSHhibrIg78VPGdqZZn+6uW3c+SRmn1
c92J9hOeiTYYB6BMjJXPrKhEK+NUDPXhrEzceblhpXo+JMpcmghcZeBt7+Sz
8Kmp+jOBDbiNebgQ97NRg02ac19u0dcoDy5fb1PBnQFCJtAUywcLrl4ApMDS
q6VoR/CR1T75PTC8t/bGLGVCrBkfx4XQFz98eYM2UMMU0jFviTU+W7dkged8
kI5JUTpS1Zl1U3+HbOhxkp4WrFAeMke9pp+f+6RUpvpzR9igMZS+6tClZ4Vo
WSIbG/bM/Cikwb+EC6wFkIjRHVuW/w3vvupXXQ9F6tbkU+mr5fV2bIUmhr/w
wdLwrv4rqPPvxArP99yYqQTP3BjPIuVuyM5DrX1U4BT+40oIOCHfos8SAeHg
nS8J/CubiJR5UOCakwOmb/jCsgpPvAV1a7M2moI2D1X6Ulhsh3Sd6mtmyLyG
VTBjVyCQFElGGQ2IhD3rjPyGNmW4Wz3ddKC5Iynzku4Xt0CWAxlIwBjvPoxf
iHCSP5dsKlhmK4UZzYgViw+s5qyJd0bzPWWWUGBLOxx5Uv7GnjCvOhPRqV63
AIm6oiKm4d3RgNEd7BVRs/IVSwCIzh0QZdYrTOr+oXhTv1g1/xxbeGDdQdn0
FRdvPI6G8aykj1iDciN12OyzfJ2Dc0cVcWZ2kU3Yi8W7VwYIFnhqB8xnnii3
mPttl15hIRbg5Ge4SYDYtsZ/Gb1r0OQvAbsNs3GngbeVEwx9TZPpnU6mUQ/n
uEMu4yiaUvL9ktRxJDV6ShOsYbk17LUX3pWhSc/KankXAKmQ0GBh1R9xDdmr
NiuQVVWj9j3oYQdO0uqoSJm4IYZVrbfg3G8QmJE7M4yg4vercfYOiknb6NKp
niqncXAqcQBDLFTe/4RhxmF2D3u2/1Bj/aoP5BIvEWYoZnvSYJM2i+mqnHLk
Zlz7X5R9E4L76iTsfP3fv9rUt/iWD5+fJ4WyCXbxBYLwEBd+uaozFbrnDp1d
EuoHuBLi5GRgFB6S01JywHXa+VVhmjondauOlsrPgJzQiNEKbzaITmYQyUaZ
kf+W+IDOzch4DwTIZxgwIDETaV6bxrcrdPxtbtq4ts+/OOdqFyzyhI9fwhIC
i2TknECAgRxS9zQPDDzXCs2zGoqxviJ+71Wo5RLCakd1pEr4ol5D6klKSYEQ
2UAhdGYfUbalvgAsV3sdKQzFU4q53JMERGkW/CADWzK+nAjVJEV+9WUwr8Xm
jlmQIMPljXWX84COLEsw4l+dawOLqXjYLiNCreqKMWDsnVcNeVzHdcbBVpZb
xVnXResnGss7F5pmcJXzUj1yUspPEzdBnU/7SN5F6pubBDUeJVAHWjZL7b3b
JazJhKN5ZlLhr1Yhm3Fkkdz8VPykMEpyxok37xGTB6F1rAaF/jIgUB8+J5XD
d9Vuz9kJTQMAOtCK5pIcd2K3hoaO84S+Pm29TCo/7/o2nsIx0vrl1aHZXWTG
Llej/ZePV5qNznkXEVTtmY70D3/9tTbVzmbsLDCHNOFFu66AqmvPOEHONoLs
0W/UJrZxJuwQUWMlzuvBVeuvDVqlYyTt2BGU9Xafoym9zFIkv0VvA0FBgAlh
K9IQRpHaupc2l1+rbdEXa0WYVmyr2LmQ4yyU0URtA+iGrhLo3aZ+nATCAEj6
2nn68GHHyZ4dc9ipqbK1oI3/EMs0BCIJLVnrodRSYLzMP5oN1OQhsD+zocg+
rtdfKhigZY6XgFZu2dsfqvaBv9OWTJYbZLrXA4UXUoiICP4bU/pU6xN2yty9
9Cg7yIx0OOd2GtEtUw2bHkMT8vPsgGjBk3R96SW1fkT+rlgvOStEVaLF3afx
O6a7XKR22Q6gXcTOe/+2SpxK38ppm/JoWjOfMfdlJ2fKAuLqoLJgSiDVGF/+
rLveLTWAQbTdsxebxGpHCOhnFreOCXT+FSm0NWBvLgWoMF4TbdBnHDElE9nd
ExRpPQADPne2xxi/dbVsjyl+D7SWDNHowutbQvd9MBTuB38i2XNNHUzqPwPD
4OvPuZGlBhbs4UreWWZ8AbWYG2qYqNR8lUr20Zby8DUUN+QnPjDXD4I26GCJ
KOBpB+vy3sRMH9mRR8AP1AHKC1tor2tOSdw9LFtz9eP/H/FzsoD3i4Pcyi0t
d7bokOrQZC7MbkIcqpSx2d7AxyUA4oMWP0Ga3xI3KRmajsBpxMJMyboDI0Pn
jXHxcV1Z8toUtCt+OkQWlryk+bRoZyBEgajxy5OkcNqJTChmQNcrpHXOEByG
/uVMyi0pDjrBSKucxoOKXTY4X+fA+zyNadEzOpWHJaEmOI36/x4e+NMSpiXv
K4Hqup3V10laD+uT8SU/uwqp204Q3JWBZy44gYG4uz6h6g+vW++CpRg7ipb3
rpmNj6FiR3sEp7gh6d1g+znh5S02flDoVb7lz5e8z9inoETARGPIu6LiQbAk
c9OdVl9LPIvYieVb1/Z7avP/+/7zGyLkJJdgb+qg9N3E6i+iarBKZPrk3N83
ev+aK9l9FJvhRKgR9ycETkHJKizKr5ZGTyptC9zBmvZsMyiei1jBJoGK7lL+
TwTlEwIEys5+YG0F4RVo9Tl3PzXudke2Gl8rBdeIp2IcNcbNYah+tyEtJYGO
tl/hZryaYNWLhJIZwEXYD1GJE3+ciwDkolyegZdcjSWuF1/H+mE8ChtUKJwZ
0ubgrG2IAUrR3yYZcfKP4IZHfyPm/05xFlB4G06Zz3t6Y3K+jJG+HMSrb2pM
uzOwWuy1zcw2ywTDOZASRjiFfdGHmWuREyf/upWkZhNk44ciYAMFQfXrCbTv
TvsU6K5MRG9m+oufXu/2VVJ6tf27AaAoRtXX3HNoTP22zdVV/Wk+0OdccvaU
9bwQLiHqCfbN2hxX1tt/k0Y/wSjdflfrZtcXXqOAQ8NPkKknwH1wBVGdSFh7
5nEKaNJfsX7/YGoe/c/l8AmD9kWiy/LSxfXQz3h13KTl8C39SWWsZPLrpMzY
TOw509Ljq7OElA3K7I1sjmTCkOzdDqFt9dxXsftHmqPrLCQA6VjEepGiMtjb
zeeOGutjom7s2+ip2K4vwL7XcJ8B1lVZ/gSI0pocDsZK7gURomVEU0rMGkvw
e4MH14cemeN/3iKJQtpAyP0hvYYB6z15LVON5MqVAqtJz2i11B2Cbr3cUr2u
fZ3nMLgae7skFdeTkBO8xjGmYWeEW9E+PXN30HoR/aMXhqdgXwMUuushtq58
17STyT7sUnvMjOiT36oTsqfDY+418fzuGcS6iJ0IASLY5GhVBwP7lUKVLD10
21BwTIucMFeVqmdD6dqL3+Eg8TnewVHNHRPFKFG7pmcI5h7kcqOaDHvMIbNF
Q0KYGkDBMKu5eLdNOgq4BUSjHpiAa/U2W0Se746YzHIrgJo9byHZ7YYSlTcg
ZFPPXkW6cF54vqVHn0WVGSh/7lt/MjBDy6v569lAjodb14LkLiEDlxGwOnnH
VXGNRiG8kNV/Hn6HOXi9JqBTWQAznZPGVLQIpD9BG31lG94iuyQei2rMw/7c
gtjXYVCw17tBkpBLl/XSY4iotYdNsoGAf1RkzWrnByk3D8AhLwwSHiCFaLbx
1FDBNwAIkPB3jw8S8jufeGkqUUIsgaq2bveBWMACogxYPilf0cv3/Hhv8cFx
/BcwBkuPeOtPNjykp5BkYQA5Es5EmbLfE2a+0NDEAomcdeMnBSwoY1kMGLfk
fF0pRB3VXI2OoqVEAg5bp/bN2Eujhv/8FvgUtIcCBjHCunlddnZ+LQDYeTAw
YAky//bRtRpT3Zk5KtQtHet1MgfeYrzfw6I4eDl6P+m9lcRffCh2QzmjiiIw
LlvS1gHd2jRuiwOGhEyisbXVM5H4gR4ptVvDVh5pCi2s8fxNHyh0LS8h5Gz1
w/c2I8k+lJuo0bmHicsYRBLAkiOaQA7LSJyuRSqjc5TNZHp0OxfloWgeOcJ6
fizAmblxUf3X6eejLd3fSUxgxKYGu0j5X45at6tym4zyZ48qBd62uoTLof5e
ZLPqrsUvKb9Lc9qcPQK0mwYEWhR3gqNjueOShu5X9rEQe+yV+FKQrS8XK2uZ
54C33HnxSfhW0OIPchy7oqphAdPPv+0oCwoqVVYD2lSFIeoMvGjC/HTsuZnc
OE3sYxru1BHfkbwiWvg9zrcXOnbcCRVn74xO9UmuSop4BpfHXcRFsHb42zac
hummDwnoQvSxW0xb7W0r2+IFpbX9Fcw7HOK98uB4GcQRsudbqSTE+TLBIfNs
ecBQ63APxIO2xtsi6bDzLh+4Or8nBTnP6p69c74CPs4EIGs2FTkoK5LyCFqB
kDu+cN6rLUG3QhfjCLQLsZwXHewvqNGUS2KMluz2WYwkfgL9ukHy5Oqbb0Dn
u9t4xtREgLixEEF1U5hYjGYm1FwCilDlWnQpmu3vgvCNQABDJGCW0WjbmZFa
IlovqdfUgTjVOJQvF3GgNPT5LfYY/PT8BYANjZmcrtXC07nwH8/uCHT2w2oR
fMf+gUs+bs6dIDn9ZIRkAM+9+Cccg48xsUEcwB/Fpq3YdFgAm8XDv9WQ2wZR
iofpcBMsjlM50jOXBDteREGbY+81sV254e1jQ0nacrAkFd/2ej0pAXVHhF+s
zxN2UDLGXc17D+xqfmVoauWAWgj3fQjbkLm0blqGtzqg1vMfqksKKd4vzLH4
2gw3xr4DOJhbAL+6jDJDaK68RlrP04BrRouTnw7Ktju37GfhKIMYkLPc/N7U
JcHDErkFcCzLZphVOxNP050weNI5yh5wcj03oYWQajzkckDN8DzMzdMGEYJ7
sODD6R2UCGf1otgJmbdLhu0XDCOlu3M1c6yBZIs+TIFDSjftTb9mWd4oVobc
UPG0vjVUZGvqAVwb6e/cWzTn2xqecF4fxux6YF01ZUwEa7oU+2WaxdnReLux
/k3JvQUQxKPtjakAVljogt5mvOEosgjv57yvnbVhGU+hGfHO4DQ08ldESu5n
dmUYMN9R6rS0nuA/E9p6Ru3iCGm+Vdhj0j0JHYfVGXzBe6h7fW6LRk6u+LGQ
YdFtEz8rsLWKtYzyv0E5deGKO7bTzCA73It98v8ANtK+JmxQrU9QdsO0Oiv4
c7KD37AFo5gNJyte9c/XMVmz/kane7dxbtenrRkq+J3ph4U24QqNYlGqB5YA
sYsvghjFCmxyvrLZeBm3Nbdl7NQNFMt+/mjvtxKOxqA31rkEFaEukB8lwUqd
VSxnn/czPNR97Z5GkN2LQ0+3zMlmfP1abpzkYqZQkWdo2MMfC3Tpa+W8HJGy
bKruW14UWOh66BLeLRIdg4uxkvB14Bh/UFlah1+yEQRNAEA+XitLC9v8Ik0M
GHsYa1V8hOSVUZMFEFHmN2wDC0zkmtLIjXXXCOoSXAKtTmPno9XzT5SubwzW
AcwtOWT1uthhZVqZmQabc+pMcj1lzIEkatp64XHQKpohxERdaMMit227krjR
P91pnu60GOgS/C6FicLDRjewB5wBKQdzJzmZOa0pXE3qln9BrEYSrUpmGsfF
N+4/h3/AsMoQ1k8mL1j/fsryl+rl1+VUeTMqHc/nV/7yQ8Wc8hwe8tdQgsRC
W7xxiPrVb+YFC+N49aDlybH2jjVXDJZzb8jPj3zXB7A/Ytd+pq6n793w+mIa
l1VsudStvjKBNNAeDTci49LJbnbAv3R6gFY3QZ+Y+LGCNDkVxAcScncyJ1wF
h6foqZrY/kzThr+e4Z9tuplEUrWmVPaMPt5O6sH8Gha5KHeFwSsQ7VvfpL+x
S5am5Cj17UUS2RcIMjiLEgvfxvdbyrknsx2PUrty6VmCbPXimtzsD0vo4nWM
nFtlFEn+f/ZA7vGqU5fXFiu5YnTIquU5bhiE6xbrIjcJMrQLs7NBY6vXFx93
1h9Z1OGftfrZ+73X8trezR6Rlm2UKWRc8nrjegkFQl+xtttQz71Eg12VxNie
5Tvpb9vbNmuT/0u+HkfPy4Tg21F3rA9sFnGXxr60dLi08ACY6KwHMAWM9Sq5
/8G0RCQnTpnAdmTOPhj7jGHpp3eJy0Ah9BnDRcQ0YBRZuD40e7w6orN4JjuQ
HpbPFZ+1n0J97EuZjDxm4THkLoZVCPijqOauCxtA1sxMu74gSOpJJmAhEv06
RPsncpzhqI7fhCG81xGNNgS3CPtyqb165bzMPjTH15LHLA00RFTIUHd4jiP4
tyr3rogNGy5jJArVA5N5tJa+lC7cRX2XYC4+svq5VNpwkSZPcZFe6lhUDwUD
IKLRUYMojC9ktCBTe07WtOzy8+IyIFCWhH3fA3cw3b+ZkDByRHgOdYbeCVjy
IM9BWk25ontK/bNyYU9DVlKI8V/eRpxQ18Lfas51mBndj6waKxxPqrif1y60
Qp2a9BL8R4QSkzpCXgQAUrI5icraMNh9Pma5mcxNyueHpS4p+trtdnMCsmIW
brS3eulOcdJNnazc/+N1yELEgpM5ZrOvfXZKa9PK8wqRLbDe+maqm8VYPAws
7N5OQI7ah0mqYCIpHUw7IIhQNKXSvVu3ovnRNnaXJyJ1p92q3npizVQQDGrF
uutx9WS/jiQTIuJx7vR6Sb9VyQZ9GYJHVQlurZ3SyKq6VwDITHH31t1tPskd
mdDCIg+ZlXv+2aa5jUKykNS1F82GCOa1RkdgwVpZHcUcgbfDFr0NbZoSJGRN
8l9gd9daqsVjYouLE6oogx+K5s5FyHFnWEc+Xs+AN5jHsAp2PUl/ocGf2XhZ
A/cRF4W1Dhe7m2BuZ0jo9NHPdXzwDmqMNgMODMCYtbZk2TchlXZnsY8Ixr2l
//4q32jvrsWZNVAs3hQFBo2ws2CHeUmRXSNBHOhd81HBN2KL1FJwl8HZv2Uh
tfCT7jy9rNXL4Y+GlId6HyuaTiSUNu4YjymLDw/AQphje36kECgVAn1m3Lfm
4g0At/OoUkN+noQlE4RCXaI7D1qHbq4vr1xbn/LCZIqH+RR+rr7rsMg9Qgr3
x2wkO2V01qkiyLbhtseBU1R3ON0Aci78fyXlXY6URX2EjopxvC9w8zaRYGmo
eAwvCCq84mzO6Q3Umk3YTJz8JuKeHbCf8EUutQhlSSvgkW7fRzFFduFl7jlO
lHbJpztjhSwjD7wHxsEqXoUBgEnXvrZMZ18kjnzejHN0SzWXQxn8Cq1EvEBP
d1Bcs+sDKgfk/7nsaXMoDZJrToCuSdm3p6FEJUgI3UPyzhr7oLu7iNqH+a94
86m/L7zL8bYZ3JyBHwHHqMFwarexuHk6uJNrHIoV7k8uLAhK1EYqAE4QxU8F
CDDt81n5tvUw61DjPBrgxHVb0oxc9lGE5rUQHqlj3fvHc8jxR6OFp58g9Mkz
8en6Vu/alOfZSSLwVRBFmEaDMC625Oar2G0zXg6Mi4oS2y0lPfGLgbbataZ1
UDaS1Fe1oab8set/T/fiC73N12dWioQexd+Ycwm1scay+ZEzi6RzyufJgAlR
4Hc1AJMgtUQhjRDdm2oEz5LVf1MKjsasNLa3yPWhvWqZBPgTJ/OSHhitaMjd
TqScyAWU1JNALt4Nln2+D00CmPrce2MhULv1XaJxF6yp0I3LNNABuBwD7EBZ
n9dtQPZHoSnt1VGFV4m0th4qqbCNnETA6I1GatamIEphiSJ0tEtnPWaaW5kY
gLWNgfCd/eqiT0lzc/aK3cLUKnIioIrTuTkmjtukF8/Yhwx5kAU9eequLtMt
SXOy7ubntKdlAknIi7V3xF6sHnc62jZf5J+ISt6OGMIm5p8A5d61VIwfA7v3
D75nAb9euvE7oaD6G25KcEYfYf/Ax3+Sl7KRytIVZnmxoQpGW23UQ3hjrAUt
azt9051f/Mu5PmMv/MKxjOokHJjeXj+GP7dN1KI1GnpzCodZmW/9Kt4fZxnV
meufoobU89hKXusZUz3i0skLygc4LWg+0fzNQEdxLUtgf6lCtQ3vqi1jDrQH
FApgEfm2YxxWwPWfK+XArhJbSCGFZaeSLPbngGFnt1jdnmPz7G7j11aOMUKW
ZuuVfCrxUm1SkgQFM0COkxrJio0LJgAlL5P7bmWKZoI/iSuz5q2MG1D0FcMb
MgzmxtTT0bijQVqzotaPgtgXcuLw8znljUJYMrj2gMGOreb/526SApSJXi6J
y2Zc5GUAMtSLGdKx2bZWP2eL0nCjHpPSXrdLXz6XHoBSCHqD0tEugeL2WIbL
2no66RynWMuNQwaPYh30agFS6ULJATrq4m8CF28v6l+UciOfc+VaNPx02qCD
eNWmRR59mvz8kv5mphQYvgN0ygFGyGYrqpVrYeYUmR3D2ON/2Yi8AXtVdiG/
obQ5uDWo5cmD7k5wII337Ufxy+lRATyL+pXhmpc7OjqYCBY4IHtxIp561vYP
XWIm2wqMVSB+777gUg5OBlb/VLLe65DJjPOxVg9ypG2UoFO/DxtI51SPC/6T
U5BvQn1YB2HdpuUu21VtM4syUrH/kOj7obZ0V8zGWn9ooQna4H9e49SXwjWC
EITPem+ZTw3Wl5rhrHqMiYX9oVt9V8LQ9Fp5A9UV5e6F7yoOcpw4iWHojy/F
fiXPQ45/uKKugt8RKHNGSxpoX6RDkz0oQDOg6JIK4/L1a817iO6HlD3EPIma
qaKRscg2aGGKOijcOVe8+Z4YjjbpOYp4h0ESqWKLrwj0JqSiMxsKopveyvKW
3L+lCE8gr/om2Zhf12QxPAR+yDddJmrZPth7ut1c32+l9GLoO6L3fJBbK0WP
U13BFLDbdFR1fUP7cQGqByHi2TN1RiRc3/LzlAd8pRax7ch6li4sh8mtgkEC
keAFFa3G7WeJ/FWcfxV6RqpxMtEnGZNUS1HpYKBsk34Q4OUZxJ1iqdjD15Pp
RDLx3sVwghBodFI8Ko16hpdc7f9tE1imO4WGHXWQwK1phJf3BRvutIk7oVHe
iGwoyFxkF21e/QWgHBcHCmtTZwxz+nGo+7dlsPjxjBRYyrddPYkVLsQ4r93y
6GmYISg1DwsmELldxL/jUwKJhRkupQU5AZC+DsQtg0lYvlP9sk35V95nY1d8
e9Gv0JtkpphnDvjS+Zz4CXdrruxNquxc1R5jIut1CXGs4OEUm4lo4E14Rr0x
9EHBFuiSiTxKpHpKfC29Vl3eo7EcrHjb4UaFrlcikVf3gFdc9k/l2cr54qRv
nXTVmHAwqw1qcYeOQ0KD6dJ6zRCu/gcza2y+ftQeRie+e30Bt8qfa2+S4nuQ
whrkXv0MhaENLBfGRETf+yWr0fb2guMgiZ7lY+24rFuf/lwmDZz+scpOFOYU
aHiva6kAGj4zH9nxnJD1pSy0kbkA5bMMv2xztmecBUDw3/Ws7qdb6a5wupVa
6XsA83JPXH331JzyHZw0n5weL9i81eWZtnB4UpjlLLcyhLpHYonvAqEeUiRL
6TK2f7arou48f4vyingjnXS3IFdbd6PRJJwjScu+FwlGtQXK4/srKD1kN60r
F5nG0ga7VSJ32ojAEhZIfM3/92AcPkOGZ5mlWmc+4/w8RQvhOruXzHoXStv9
r3/CgulUNuMNSUcJiKGYXom2oGjzPJfCvMZv0BBrTmBowzG7e1EpKzLJK3VV
G2u+GbLz+JLzLccXFH6mnQ3ovCNzqpyNWvvZdaGKYp9NxWbMTd+izR2v2ZGa
Ka64di4NoRNp+B27duF7MMb+TiH+u09JVtnOgbxB+NRfe5UCX6LKyYDkSGpI
sNDBeoYM2Tjl9EOEcHaKEbXmBN82JbQZLKd4nAnQcUK8dHWtHGcwciWt89IC
8w9SiU0RBARgpQapghY5vqJ0L7rXrAZtkyvCRW2vVKWQuHhy3UUXAsO2rpov
JMtmIg1yG04ZGyrqKYlutDfwDylYjUnQdgG2ptkdV4YcY7u/s6sXHzdpv9AV
HrX1j6cub8z1om0QYT/UZ2TkOlunOETeSv7OUOCSFbOvh/i8oqqu8QmIyHm8
taTK8ItgM+YRcyM0vtzUyVvBrGnyWIiMeYEUQnO/6Y9fF035y1wA1dUl5tkj
COWWWulilYmL+j2B07oU1C1WGcnBCM2RYBR9GhYHEpHRBoFXfRXsVxHQ/1qG
DHA4tnXnOXdnxRTu4O6saBQ3XZkBoDUEw80bVnn3/zgXHCi19Kkrv8ekKOlg
0U868q0+OrGIvIRKVsuwemSgzowo1GGXOyAVSh0H5sVHf5c2LdhA/dsIBkAn
ETzV+b8LschRgsS2deZVObvGW0h+EThkOrl5HfkxJ37MbD0SID6UcIZqQbiO
JWstN2CIek8vRSdFl4K6tHZHVQnWBwshNaoNsf3mg/JKwrOIYuJMEVTri3kf
emufBYcv44VeoV6wG8eETaJ5KLbciS5h/rV85tKgyJbx8I2GYHODtZsP8/Ds
+HcOIZr54Huzygfldl80T+9tsa5oMn5A7AbNYS+CobzIF73VgE0iegrk5N3R
XFE5V7wq8mzHyChwAVg8a2PfXHJOH4prwVazHQL1jneAGcRFDTT7nbUqx/tB
bmNrq/gaHveoSmOq/tVLMbMMFCSZXYF3Zc4wyJBcY6Cn5rolT6NfSLBTRxqo
Ow2tzg1LnAQhdXGfeFHIqzUwEnuU9l41R6r7ahdWzz0XuagYDSqLLY0gDIrr
VUvBJfCNPh0Iuo6k0DKgnfYDhK+J3o8mdUx16BEGMPQ09+bcyOKRYuXYPH3X
dW/fNmn4Scb2StfTUtw1Q9r5pOvpBo0yil4w9iQWAKtGHD4J4lH4h7dbPLZm
EpRPLCZJHeGzgRrbb+rd3Qx1BdHvvWJHV0tMGSP5pigWrgUvph2YMbFvs28H
82wL4kvM5xz+5NzgJkVDcJrK8B5wI1B0du/EQwF2iFZwj685uO20ZxKzKGg1
L5U5I8P7h+wnpvs/vnhwDHTo84U+QBAwgZhcAoE5pklC12BcFzYUmINaUFm8
vXKw6ZqqOLB1xekw9q2I1W2d7Mbo7oAEKeNpdcISpbVdRKVYCwCWwzLKyWZP
9GW9NWOSKsWbiTFiN3v2mwPANtuEywmZfugtWqO1k5lUU47itEZP72RFeAx3
j2t/uRQbmYWOxcnoncM8uUQbBP2eLjLvcxx9g1YlZYSXIlbLfZ76aOkFan30
GBvIdpDu/+5HRHi8vSHdx1AGWYrkPhKAMJFeHbAZFg/AVNnmsud2YJRxU10R
nB8m1zS6BCH6/zskej3BNQuMotJ1A9IptLFJvfQioN9twXM5OS3ekbbGMZ1W
9rqtACDW7db0laXWUNXEBFN8oFbS4NN0KHJY1ji3uDL2JzvLkjKwYWk+8WRM
jsBr9bdDavOeRVu+GPrtbt7qnrcJMwZlnIrzjTG4ezf6IBm+mBQ5l+3XFIWr
kUpxoloe7VQ3wYo8Eae2/z4+lI76hFukMihzGzpqi203QQD0kN8N7Yck7q+4
tYZrkzUYo7b+T2/6kAoTNnznUfRNsmz6SJXWh48tzhfAMgxNWy8f7IPWoygd
T8BhcKtZanstrG+UgZlN75fpwPgOTbGMHBU4QmjEi6rLR5DuhbcZZF6lXoOi
QZrpnTMjV8vMKjPDzAiE/y75S1vVXH4ie54QprcH+TkRzmCPZTTonpfyM2HR
cTxPs95tJjh2IJMYuBTi+S50DLi5h47qGsv1/wAcPu3HMUzOIzem0/EQjEt8
rbr9ihHQ8/dAsdqG8bpRbeUX7t6YPi7NyaoKOsREMXqC0G7CGZG3uK05TjFq
ywBoe4TEs4mf3hjEj3FUWiuGCebL0RaDnlXu4fzDrH4cQ2IDPu0zLT25ppCH
C9TU9hpJNN6fviEw+A1f+F9YYGb1eMxC99uPiu/xKKRMNDokTt2/pLFkGNOb
0CkmW5LR4frw+CHbpq1caoOF4MgoOxxxCNPZdROurAIyitxkF10vFNbZBpAa
vvbVGPAvj7fUntyUZvzSWEqSUpbY9/A0bHcYBhSdrkS1QCK2k/5KJ07pnmVM
qp4Ec9n3vcrzukm+idP3mMC2sZA8cGJ99VzvVmGfiEdgKMrvBRmWj89mX1nv
1la8n1T+CB85Ot8PTC7vmIY21tPvYQl5EMaK5NKFhjykL1Xeq38YO7/Zeu9C
KiqSH+J/mE8q1/EIg+qQ0I+9w036ROzGVEVPP4DLYYABqxSSQqqMzncdDEbf
t+FxJLd7MS5hXetISLmuWenmppcSEiVykKIgtC35cqQsAusa+zL5grakgFHG
sEEmwVoFst/FJx0+dcQIT6Js6jyHzyz55N7U9RgSCn9fDs4TpQjDSj/jr5Qz
mVa2MW/M4RlT/yPU7FwF/wXvtEYGaeqIwnM840v/3YBhd9wpQna4Wl2tRfBU
9R6fPuLwr/3jwmfUfN3/ZeugjWZkrqwbv7qoVqdxoZ3/4n1+mx2jINi+HvMp
y21AyKZ2qySblxMFm+cGq017RdxrEQ70vPCfZskKRPy8Xc0YaWF0LXMjtKk9
4fisFQhHtRhLxZzSrN1fq7NclRDGtCP6y1yGb+xM3Ys3zcE5G4a2DQb9oEAV
dM9mLp+3mE0MkowlKCkJYbKyIjHMBIYnQPgQK/RzMNc6SpLmXF4o8hm2j6k0
rMdk1teLNGSLsvzfT+glDohuhmadI4WX878bpDA7UyYFwmoc5fr04c82NXGq
YgJZ1iGOPeCG0zIlFx8naglt8K0NEJ7jDt5yeZbZGmeLoNd/L+ehr5VKbQaD
XKZXO2URxm8H45dJN/XVH9ih3TcGcqB7OccztC7LaMJJGPjNgZPhysR7Aa1k
4LCDdVmYP4Y0pVQSvRl/MIchAudNn8W+h7Cq4HklkuuqBtpGOFggZrtz4HvK
2LwAqaOCcBUDtagsL4a6foVGg8XTSrbp+8qnH7Nzkk2MLRkat6W3089DauMX
4FGRAzrpV/qxjjpBtKPma+DxBQIICc7vHKYm249ctpiDPxgdrrxBzzFrJ1Kd
YM82qJ4zJPuhar2cXW6xeHVYDhIpRV5G6ke7CTofe3yR7EhxVGfzC4Qv86uQ
ppoo34EZ0GzpSApxyLUEEDssjAzkGjwPQrGPy3GjnjtKhPyg89OQLlHplpy7
6qtPuP2iqkc8FXvGkKZIFrKtw1wWnQIB82a9Ju2/rnplFSgCYnhJQFOZ6vPY
SofrTvf7H69zXse+TT9wcMReQpPebw9kmkd15MeHalnxZ633CItI+OvNzpLK
4S9vJD+qPLPr0qvBOfGZ2iYZuNiHAgyPkwQAVPjVnSv1k8dRstGJbtPKOLKQ
68Er2I2DVRI4LCoEFWIjWlSkSFmSZ1eojKHknXQPAu5jjbCDbA9ul6OhHuTK
bLGskJkaCAl0DGVwx6zjq424mXRXj9488cGW/GJRksjN/oumAPIuCm6rIrkw
brT1pnu3CUFkaW0sHxL6AX6/Wvlax1g07V+L7oxZGTaIDNsw4HUkgeHyrQhk
yC8Eczl0eAKjp9kVZco+18ttyJgqYISsg6220n6I9e6xYe47UVmjqAEsfNXA
fLvT2R3pSkTKPNfY7FV7nI24N6E4x4/hFNs+bV8Stolo7xgDx2v+I+Fh8/a+
LEmnYj4VM3BifecDH8rO176qRPNt5vCxCcjWJUSNKj+QAEoKGwxb2PSgYeil
ZwmQl6+Y+BLSaMwfXlFGc3rS/xFAVArS01peKyM5pmg+tbSLl9ZXidDjR/4Z
7ygH66omTK6O/qgmdmDGhkQGweEPvXuOHaFFDfaW76LH/YXKyFckGQ5iBe+p
s6bA1QYBBqt7qoW0maLe7uqoGT2qu3dVrUQu2uoK/5Nv4x1NwoDddzdIOfDH
gWOID7f9tny2tfFP/E+svYKTeQ/5M/w7AB+kHPbjpeNaKPM/NPkK1Z2NknK9
+X0nuRYbDaBeiviVKHkLEXA/roTiYX+whJXWsm8a15E3ff2aI2h57MxgTFXf
ve96YYy0EDitlPLV59+p0ZNTVf4jE/1QqSwWhHKw6letlYvVUbdTYEt7W4F4
pq/qO5GHkyL/ZUQLGS0VCH9InqTOUJ2udH3efnueR7/R8pVGHpK9UaYWYVbz
8kQ95/U3JDv9DPeJPuk9y0QiVvpDpXkAVBQj4ZAMITpUm/t8nfLxO90swnD2
srk8ceVXmea0PZas1j4vqYjhNV3EjegC+kHyjMS5Y6THLYToVhi7IlLeVda0
jZi9lU+8Ct66Np2z22KSGGKl8bPWJIU3PsTK8pwAz7GBHCfB/5HWD6CBKDvg
tsrzUDvAI214ZO9yIUO9hX3B5PmuKOo1ZkY3hx5vTM1tMAHW7fs243WCSvVP
9CZlMSpHP6Ggw1qv8BgN5ikV8I+Lcxh7rYKDWrV9VNafrUM78I8jE0NRYIJX
7K/03LYQNCafV/g/WqSKLzcz44CtB5J1SEj1NJo9ZN3FiCYEqhBn5NLhe9ox
AzG9DqgTdOAJluGBI0FxIl8gq8lBz057eJNOEv8DIHWDA4p0KC2V7t0wDvYR
LYKFtfj4gyr+w1wsQbPl6JN+HQr/m4/XBxvuTCEWIQjpq+UTaqpPJX67Gm7N
LDipJRvYgnKFo1xrGZnHxIycVhMyzTfflYa6nzVL54z3HEEankDrJBOQlTpI
BqVJTVRpVXcLV/k1qOtU+YK7p2bD7tbaTsUOAUOV+nRaoFqak0eOiQkaQZhH
2d4xm5sS8v0CXgkdliq5uOSnHXVkIjgmpfw/LdPrvxS2zWPp94qWQzeiIiKb
7CNKitIKkd4Ix3W38hLSUk6V4/WQxfciduQsuEgMioTDk3do5/Lw92gXi0D+
B9jf2Vy1r244x42sUe/dXP8w7NCeRrn6zYVTCr1oWvwNSVFGNQqdHaoc+wSp
z5Wm0ZTDntdCnetdqqwhxIkO9/5OibbWZleAZzc+q0nJGC5jXxOw5S6sJF7H
0oo4PYxMHn+GCKe6vYwU2RdCSoG2WwvMdgQAedSmNKm2aSQBG5Mf2+2jxlfm
QmSLfnXAa2oXjuxq+Aj+/es+tbLOQx2Bxg8qVwz1o0babYA1PTj8VwQ+4iA/
4q0OYHa+mJISmZ5eXlSkSS6vxFwFXOXEDgC7Lhok7JGLI02ZoxUGYzZ9Xa43
rMvST+AIUimKbvSVVYKjVRGtKdUnuPux7skWkCWTc95Rl0UsLljDpGQ0BycI
PyKR7aa4oJKwoHC7DDPTmciGbBac4InO+9xkJf5J/br0f+2KEimu42ISffSu
hxWqzec7/XE/vzn+GREC8M1aJ/E5t9NeBvKbZLcmH6O1gLCGPOBuNS0z9F6Y
f4bfA0VjqvrPYk9/Wag842jnp017B/E5nnNlG+xfFRW5jrv1UE8SXtw8HXuT
T64JBxsy5arfLAZElM0WOxwsbalHNo5wnyzK6zlS+Me2fD4NbnW7Lqeh0Qpc
8z6jetN+/cDrX2sgNvfDKI94ZEi0vI5c/Gh4YFI+eW7VLAd/aVilkD5JGpou
KeHanRcs4pjvlQbmd2g6wRWCDNFsxsURn5iFTtpveroFp2ZiRr5iTm96alZd
UzDPW/4TJCXx9/nvZqAgRwgX2lExEG4DNXzk+SOQKHB6Hphpft39dOkPFae2
ULWRlc+N7T88DMqS5rDEXBTFYKk/LjS9LPLiK/4Ejz0Hw2U6DKZfNHmlFFfq
0TmkaOWsNBq34nlcjOGXgUEz9rJpBuyfR6j5/4MxgEX3jdJpim1ecbl6lP5C
/sNf3HnE9EXFwN8IpGlIeOjKEGEwZiZESrp9AfCtS6H9HgI1kLjmA7eOKxef
yopqzVhs46ELgG/1vWLc1KfBMI+B2YYe/4iYB0PoPrbdltYXaxfn0O2Z+EH9
AzF0CqYW7Vr42v7pisWIznn6U/wh90F+yTQlZF1+I6lMAYqwhzc3W7yk5slg
AazJA8hUdH8uQEBJ52Lk96TVmB+ARzGsHkPdDjE7d31BouNQ4pK1ViowpvWh
BgYdE5GyIynjKbypM08GNakbIpv2lV43wTagWarrYfo2Qt7pHLgdybqpDr5/
GNQjAOkDeD5fuWaZQObYaQwdfDhjdr8ZxyFGotn3vcHbDi7GCUD/ypGy1ffQ
IFlgTvTgddRpo46jmE6pMhZUp4thRgj8PlMHfAOAsYhZrKcTzn/AIVpgSD7n
ry/FzHY09E8NNdSJGoRt0ltc2nTMQ+9B9sHcOto0AhdAku235DD6SRBgq14x
for//ThW8GQ2UGiUg9VpZ/h2ypFEmuVQ3gDP1KXBNmn0VThkCzeVxBrjnHIu
BJQxCYDUM0QmoFFLHj2ybsvIgLEaVXepjCtzFLQ+ReLR3m/xQlTTX5k94Kka
kNQmV4bBmbVqNoCn65ZBDqQ7Jx4ctnCdHE0vDCsAix+bOk6r03Iph/uTvSj/
XJgRggSRdb/6nfGZqeo1hWyTvmsku81Zgnqp2IkATVkUwTv5ZJ2ZfgDB8zBk
3TPy5ubjOPbxBE3441EqpB99n1ZdYpHrOJ/Gy8EpvcWqCFTVxIqLBEvCql9x
7SGBSjP7YC/Pv3Dr4ioYgt8pEYnaWnfCq9WA/NKO5Ackfsny8bZ0YjSedf4e
VNQj/7Rh1SZBFpONb5l1dHzn6jY9HrXjYpRewyPKuDrgmbMjVrm+f/NE68Zy
EGG7hBtggGBZ7+mekStv90WlrXnJ/GQVW5QzZSJEiYF7+/OBKbIJ/EFIj5Be
SO0yDUlScPOivT9knaMQV1RzUlurES/ZHYVhis9yr9xa+mm3UdoFAb6bOL42
nxhZvRI85xkxDl7fyUVBs3SyRW9aDbuhxlpe+enRj0Z4ouvU4cYjyUninFjq
tQfN5V5G9SxX5ELgVPI+CP7ugBKHJp/ZU7Qkq9YWxpjHFiJqnNugQQ35fihK
Aa1F9qNS5YAH6mW3uGPllj1HGvl2ypTm19v+YVuZ7Wxr2k6GIAVg32OV1UJw
7KBzQDOQxTDrrk76D1qOV+6vJZ5qTtx20TYRo2w49stwxEYM0Y0pAFAigAry
UVP8CrsgjbSVtMY8A/l6AhNnqg59A5SU0ZTJWSTk10t56AteEYJR4eCDnXT1
vjEDJnrpZbUtn5gebJ+ClQTDm9QTpup5T948dxeM5DMYShArwKBElnFcqWeH
H0IJ60zSesWDDfGWGUFYspliCj7nSSK4eDOSoo9RIbUYr7Pbjv2kbI0/P6k3
lQcZvnjJTBKDiH2ITDjACCtS7D9jHwnDt77yi8QkfETGCfPgq5D3WpvsvusC
TFE9nskQyEXBM/vKI2z1VekoRg8CQJ+nrZTeCsNLi65eDKUerG48Etqwg/Za
dKNXif+YRgFnBu1qoMRi3sCdaF5GhjXsuaXs3CACBSXvuP+Ih1/ZXENcC+j9
QKaI77hSQPXoMwV4U2nZqd0auI2N5faXQ+8CD8f4wZvUkWJpkUTLDGU1D0c/
KL7DMCCEtoVe9AKarMGeZGFsrLU72jAYTQUx9hFeDlLlLN1djUlXycQw11CF
Ukjc3XO2U4Rmc1etQlYquDGaxijx2Lc32Yzn81xIkPBL6w/AgNoPP3OxB8hp
AjVPiqcj5H9c6uo+J8+mPQkjRVxGAZDyIfAVE/I51tjNF8mKnqcqghuBA2Cn
/sgK2fliAnwOWyepYF8HDdHu7dxWfidczdUzntWyOGFZr5Iul8vSpzKcIB93
jWyHhb1td0yA2UoZ02eLiVVBJzBjOCqfIh9CBzfkgpZeJlXdCRBIsUP2TBVP
F8wKOlMmMzN+3ENUWh2hqPxLVPQOO9n1ZDMIfZqharFfJOzT52GMLU4pQ1rG
21P1rvO8ffO3OJRPjVT1whe/euAbP+uxILnWnG6CpdcFkO42apAJSu1k87xc
SLpvIN7XIEFtEPdjzfPzOnpjYC4JR/EhrGubdOpd4fNSUfB9vv50AOmoxS6Q
A8t1lppsCIw3YnNyUMeLMFw7E1WKX3GLD/qhjiUSpVkefrecS7rsXJavs9Ih
CKFq08JoFRC95mu52JsMQ6Cw6UfD7S0DRdiMAtsvRezJ6O6EHaGjpcMGr2JC
RR/xSl6+mKeQnASdSdPiRaCH6Bib2HZBbviHn7zsR56DPwrPOB8niS6gX0E8
PHfgzeKREJNNUerEwnWnaVWfPr8pKIcJKrlSc1tLU4deKrlbOyxR5C1nq3TI
VqZfuU6J2RUVZxoATdDP14WEkQG/nEWSxZmN+eHT1RJJaH6d0z11kjcWiLFV
eBh/JsNWMU6NYXKQXH0rKCwPNdT7J9aOP6BOsWn9dRCIJ7EH5Ajyq7Ga9cjl
OmthVVk6XaN0AKYh/EhJwGOtd1r0AYspoBypPsJwE67rpGu2eoogVFnqWNGj
xODFZ1vraJoSJwTAmZIgjVdIrQddUQgTwlYOCi54ONhspFAD0aye5GRmXjz6
NN070HEMuDr4CxogZU8838WLLbcIgbmyTY85MOZmzWejMpoNKT+N/5nxGB8L
sTN1BLJdUXMKmOLRjvj/jasxHKAzhLwOyW/JiWCfqfCKTrAOK/F8Eax1xZNR
ZOUnOrF4EhRnQ8X3kA/9kbGr5boc7MYSykI4zfMLeZuL9vQnjCmaCzM1iHJ7
a+DKNgD6v7KjZ/Z39u1LKYPEoFXYeB+smgMp7y2m7jcnvIUC8romk7H7kr3p
SWL6sURRDXGyA6Rrz0KaYBFn3my7J0+yg857usofnSCu9uJuWyPgyWJ7yhS/
gOcM1rYJt/qoJ629+lT6xHZI3KiT90Fl+jG55WjlDUiymDhZ8bD75VcGvpaU
KT2xavqgTySbYcpqz9aO/rnhzTQwq6YJ60xq3ScMQvOTOxSJCSKh0A6r7fjm
qpeEXbfB5HyKulPA/aHuA4IC+P03DCJTXhzkRi084cbfbZpVEq6Lg4v23a1n
DzMUsfYWsEr9JcZbQd+6MCmgQ41+L9TI93j15Aj+cwSsAFsono1HjDJsYaqW
kVaZopacsZYbHflh0PYYiIggwl3Afpxh8EJUHQ34Pn99kYiy5TDV5Ky1KIZb
vfD4vKbw+LpfDJ4wez69+dFGffvLiwRK5GozbQJle+UfkwmV8UBZV4kZMTbS
iKTLRi8qTSL0jvJueMUCB4CPMIR9WfcSJSA7x5aYocMajSma6USLkgNffXux
j8S9O5XVpmPo8qUSV3uyqyAzEIaAAzxUWhwDgr9/4/IW2azvB7X79vqX8LBH
J+QAHJbfm3vD6PxsZrDA1h3W26UbZfUrK4sY3xmVGoxQmWmxqZHQL+dooNFi
G+Osui7zYikHuXgrhmtD5xQ3FteiCX0Jm39+CvgNQbwNMOnNXJpEn7ANNedI
e9b4rdh+fuO2nbVwHUaw5t6J/SK13E+EfCY3xKC1g1VAysvUVk/lWCMgyfd6
WXdxMJAWlbC57MWJ2bepBzaDaGJfT6qkU2QjIALvs3qu5s8Kq+jqemguw3w7
8RB9/KMMuu4u2jpB81aYDwzo6vwTmSTFd+W2kZCUumU6OM6q7NjSsNmDzbS1
SEUcMSyieEYU+jfi08p9folj6TZA1b4Pf5wsHS9kacpGqrzr2/Da0JUfFscf
K0Yuy82t51pTPsWNbZeKm7qmeiUgNeTHux9Y1juRYD+4iiYgD17nhQuR5PrA
n3XWNG1EjGWgfLcKRj69k3q8hpfALszh1909nUiyeujlx4monnJL1i3jlL9x
d48Z7mAs6icof2RagmijJpNvgYv2I9o/n9odoL1cfpIQlMJPc5x2rfqpBZyF
j/4U8WIgaFTmz5MY/oWKdBJ7w2+m5FMT1Uy/MAZN2C4XbDT/g7cBHW6FBrnk
rPjXojRDzgFWrnVqZr/Asr0xqXY7yBMn/SbjDNiDfh+LfJzza5Vl/olbgPh+
qomjnUDhReZbw/hwthZra5uZ7rTff0HFute+Z91fKIcz6M7LVgovt5+kXPzD
TxRkXj1ZoLRO851UYPUKpLmJAklQ7FeTdRZxpDb+w2FVeT/I5wdpIjiJzgtB
PWxNz8bu77xnho54JwrJjqafX7d++keW1JxsO0a1PRFaRm6VP+AUHJ+S9s3j
M61tlnmGuAbTeyb6H17jWlI1VEOUqrkKt/dQ1RH8VlVt8sDhuxmirL8c+4IT
SbuQH7qRGNe5w74WeAE3TZBUmK+8ETm9WKOBaSFNyy2L7G550tjKX3PJtmfl
MBVUcPrB2EEeOeWALbzsiUojHNwn63WZSewOBUByT8SteTWC+vKdsWHIygtQ
06Vh1jZaEgZsMWxROiCxMLhlF/x1+bywf/LkSHb6uKKClha0oOJ4MdiuwaVg
zqGb18vNFubAbnJHlO9z/nAtao3KH7V946cqoPXtvyEEfm0QAGp72jQjU9zk
UnE6Q4YhXULCgExlMPYlg41X8PUKjVHcgvVCVDNGEgd2p3L0zuMssqjYXdvs
798kbQ+UCQ2Uz7VF8DHRRcv5Lj2fjLs04LHNru7IQLf0O6LYxbMZcLqDet6w
dgf0M98ifvdAgb6LDZPHwkYTK7/11Cuu+U4AzcXJmNBlo1AuSFWj3Ezr5aRm
BwCoONC7nnmGy6NEWz4SYzH0xKiXwwz5MMjNIHxTPyzN6V0WOZCGcwAEdoOL
KrP2EyUgRI81mk+iEgDP+LdsKv8W4TUHxVDubjZJtjp9zi5WzTVx4Lwi7bN8
A4tejL+Ds1oC9k2eUczqwvTmyIY7B2iiUngpixkuCvBHg8QapCxB1Yaqp2qi
qV71yT65OxRv7zjexRVMY7iW7WRPYxNwm6Kqb45xayr1SeNoTyk2rDLprMzK
do8ibMwhcQjW/hTRI6RJ/luTfUqnWWeS2Z6Ui/ZmnWafwaArMn9wFFRHmnlt
7OOeLunW25G5SANOoGWLZgcT2fxACnMq0S8rYn/W7u0izWQevZNrkclOlw8B
faSw+HWwG40zWcxJJ9supk1RCPGgUmhwwAmdJvWvDb9F63PKDgDeByyjbjkd
genHYPCLsqG9z9L682MeDnjd2cc70nKXAvMQxXHkoJV+OqCpPKnPz87WDlxJ
cCYjJlx2IF/NLb7AOX/xEbb/1EXXU/gjvwsyKNfdd44SsonP+nh37VAyxfwx
PmMRZPkhXFWIhef7UYOVuKZtLbpA4tnWeUd5kSkmEJy72/2o1W98aHfToYQ4
TcamtqPAWaDDBqOFZuwVLT+muMvaEI8pYTTJGOZOJL+v1KPEmtMWtHi3rvM5
MgIX1RDMYDcMTyj1ZMUE2voPa0f8GFI/aBYt9SQPSHM3ySMaxmC8k4dblSFg
Lub/qU6cG9V1IHp9mtMVMlG9KdsXh1xQtos2FHbeoNn3coUdCqC3vWbJWL0G
jkQenEib+l0UKapbpI5N0LTYCwR/Vb9fr6hdGAQ2MV3QVIpbFzamiFVjhqmg
vQJEYBWVErnSC9yJTAdVLEnBLKxBjsJUqSIH3kmw10XtVx0C2/Dv83mBz64l
k3/iLMNed27EetQIz8L6lOkcr3nuHWtqMciZGKrDpUXZEvSs2nII6JJN4j0n
peEQAi7nILeYMzy2gPB4HgsjVqfQz4SacztM5VxNQ9fzAHRzUB2FRkTW45+/
uLoX+oXPcs+pEB4Gf5LgNAXb/3VJCmXOX2/4o85MyMgr7HAhju6kJJXpMolO
vBbK43fJBnVM1gUHdGHYFxRzyIKL9Rf5DIRkZeCF2RUuex7sVNutWMPe5w7V
7+W4BJgZuvSbz/s77AG+KDHcyF6lehOLJkjMcQQ21zOlaDvB0q0vKpX3xB5c
qnBElM0FioVkZxwod685iCviYSHsC8Iukt13NT0O2pLGLxQylkfY43BBElNP
TMHpM8Nkwu4As6IU0X9iUfoIicBCv/P342Z2sIMERloKR4hxSGfuQoJHdjXT
rl0bfgiM97X5OqNsg8LOEWendf2mk6RMIr1rzd0mIrH6KTmqFvt3Fu+9wZdx
QKfDZryaPHC0AnL5BKoJ3wcXKVC2ZzYvvq4c9QM6rnXCkPvHmMrGpRJElw4o
GF/HK0dEpcvqX+WZ9EgDi6oVscyKMh+IqinFneqvJFZXLhwSUPF+hcba+mKZ
abF7yXYKlxOqUteB6EFwHtGgjhaVnDl9H9RGQoznsJgTzdV/2DKoU1FBdnX/
P+62mvMhGaacM0JNIePHZAtkK3rP+tAQJPf4AjqH29GvmsunyFuNbFixOiLZ
eNnzHCUiPuwKwq3sVJpRz1kxIbNA/aYuEUIbjjZ8zZoMMpJTp58/kq0YQKLu
FG2O/9SIDc5yUAN30ibPAxsvRTCrQQFKtpxj+XW+nRRmouwZPop6klNa0bnR
ZeOEJok7ljMsPdlHNT/bCOTSltjLswcVOQq3E00CR6jdOdyuJwSKbqUZhHpm
IbDoB1Mr+sl45sAhYXGMbF2rR+px1pYVEYxJx2JmMCJ1N46GvkQQxZ6ktQjI
aaeknBsob2rF96XRk7efxeEESj8R2DUkZT7CPVqUrZUargtXlBTbyp6EFIEk
GuSTFBtvciUjU9PXqjYof4KgMZef3RhUpQtgbqwz5ETifQ+JqdniQEUX4q6D
EN2/5ZxJd966FxVOOnfe8i8Z4yiPkQmdcARhdb2pIHkn8WXzO0Zx4kv2doCT
GzrrOZMXvSdfxk3T/Zc72LfkwsHedsMIz6I4E1cu3hyZn3jj/O5JLYE35l5p
ozGN26cJZGbk+2z3wymn+hc+Ou2aoTE17eGFnX+OYsdR8DYtfiy5T0ywVjIR
bQsKDh6T7H3FVtRXsWgNlBh6F5vJO+hMneV18HLxlNkr0ZkbyAXozIQej1Ze
S7bx5Rlv//mhfTVGpCFD0i9ZFByaohQuWBEyIXq+9qgZFajyrBLgt7j8httN
oIc+LIVxgRYODYiRoe5O17sQwzif/JoiLuUj7IKZaatJUrqYxzKWzkrQDFxe
4/E88P+v65JYkx49AI4lLjkY2L/pFxLpsCZGvjy/D+PWCrF0IXO5K9IyaPlV
SEYZjqdYwE7r93BDMqWVpFlKye9N0Nm27zb+msyzSQquq2rrVqxsFFaf6AGC
+NK/TzWHZqkJtgsFZJfUdzfGGBa2E0IIk7bNg/YkwdryirEFHKBaPiNAHacW
7Kl/qmf3CnGHT3mGNHHlGeehMM2oGZrQNBPWysJ9F7c83BUI2+xpcwhqxwJH
QiGEsY0RDFMk35wCPbksCh8WBgTReEKR5fhgZLVkrPD9LZG10lxpUSqzIuY4
3xxDVWBNwVe9irBSLr2pi7b6ORGmzV+Mr+LEYjMz4jsLZH4hCmpUqIx++oC8
vM3CCNe5Anqybg3nePsFhXQhTnss9jEs+6TGdn6eXP11FdxPrI8KBGovEQ0D
DsdqrblYVzgxztvzn/aX+Ao9FGed5wmbbhnqNAq8E+B+k8BeHxGAUhbxmFaH
jhCAND9XcL9hL/dCViZPPxtFwOjY7yo/m9C/zwXmlQZL36HSvf38itgaymXF
MtwY+mamAuGKa+lk8z8HJWQgXwEfF1Wqjza6/HBoJ4AQEsdlWwDyVjkxjf0I
yB22u5yNF4E3bOXjIRWyj+Pv1gmA2LKc+o8FbaHLjWL4eNKD4f8F8/hGexK9
PJMV/Lr5ojMuBor0wlNOX/qOhw2/y1o6wWvsWchLVLrVRIX56Ztuyd0UQ2LL
FX35pDHg1EWOOjmgcUbEi3FcWVxxBg68ljtQ3Xt7SYmanKo0QT+AUW4NL71B
nEV25wxIrh0ELlsLJb9kNNSgORrh88d/OYltnJhn+ut1MHoqqWKzlUKnP+sC
naGJDzAK14vs9Y4NiuHLIEUuLh0/OUS1ykfYDDwkq1xygeBQt5Y36O5ua8Ga
5uqNHo1yZhE7QPyZ9bjJKtrEVT2RyugcXrgPMR1CCF7CFietplP2eTq9RZd9
IXPyZ46YaspJ1k5j7UskZDJdPUBeOpvRnBK+2z5GBfGZ5DJpdMoGOjDMIyju
GUKjj0VkXJudwiSFRiOvfD3z8M351Eo1Lb4cmRgw9XkxKBf593t3fygTGRVt
7eFoaCDubS4UMkSISPsKjltNUFLktj4CH0Shm1YKIQ+4qpHfFAdOiPR1GOO8
WxzKAdQDCxR4yLO0kivSby1PkSTjztyfcuoufc+46N3v/bwBjHt135s2Dw+X
2B/m4jLVZtR6ErWSlOyt/L1hUxNmFcI9S4A0PzPXIxVEMSL7BxzqsVO5iuCq
a0294Soats1slbfU4AFMbRz0e2wRtSRTQ83aJsqLHqUvSGKlbWO4hmI2calS
6U7ydK0lKu6vV7iV1J55VljFKjsmxcZgj2JK9f4fWk4QLNCTnimO5uak9OZT
r1o2s73swwmurOdhcIoYpNljjNnkIaOB1iok56HY8HkUDLMg4IS68aJHxVxW
KUbP4wcIIv29YMnD1X6Mu8h9I/keIQCiNJA/vjHnGlOkCMAWnBug9Pei/6JA
MGAdvqx96/72X9HoJY97Kf7Mk1gspvNgTXj8Xw28qAJW2DtiPaIdSKQXgpxF
niU1KL3PejtU0y6WpYEpXKK0IwwWt3dHESuQeVoPlERzuVC80Ue5AWVRjM38
+ugpMg4ZIn3g1M7YxUhVnj5xrrkSy/zgUrkfPeDQFIezRqdTvJ8zz+q3++uj
+AqdgZoV+dXV17JuJfAKryoR6kTe6OvPaVxEMxUyzjicaBkPt4cYlOI0SCZ5
0/p6IfH7v9xik6dxZsDAyaKyPeruWrd5eSCXTLblObhLr+Jq6IbJnxcqie1A
vXlZ1QgKphO4nitsQrxCfDc4ARjPzKA3VbBpUyDANp5/Kma6ta06I68Vbokn
nGVlH92Izu2s+8EqSksCWGSWJz9BabECIP0xc5UhLyRoaOGCJlhzmmBZ1z18
dswqmAZUFp+wd0EdnGFGabdRxPzgyfKXWeV7dEcS+AqpCcBvaHoOk9VZfpuZ
wz9+1gjWjnUmoZzjCj0KNNY7gMVOhHmlVOPM7YGi+PyC2GZN5y2tMRNJTJgN
QoDxpMXgozMu2MDjOrj+vSxolABtpKB3UIUS3HsUIJDEhkEAIr43Z1oXzi47
Xhqx62VMbVnQ1Z8usaZXFtJUBZROi6BibryMkOOCWA5TFaySbMthj9Fs9Xm+
rJ39DGyeaMgMN4yC8+aY6tfa2AtRyfd2bhC/aXvh2+5H8hmS73Vb9/EhQO2V
/JBRblp2y3WyWta/OlTdqosduMtJ2BF958+CaD1o+mAw28xH6DiovMko2ZCJ
c/Bka5IlzxY28YG53RAvZvAi4QRHHzOVpqR0D/xp6xccEnQsMYXr1VXqzXNJ
n9FKiLek6MQyzpI8eVZ0X2NhHbIrx87gUlnFSlXLW9X0oZ0ogHxivzVq763f
kAxaI75WTQPHOzi59poike0fUCi9/lpIfx2pGD328gj33iFkY7WrR9B4qT0X
02mlfzDaY9WRGo2fLotQ5d9l/tZ0HOU+2HAbdvB3hqPx5OzwXcD2P2cBA53G
pJGBo9u/y/4pZYDBgp7mdRpgFijgkbCJzzprR3y8xEKlDil4y1fUzLkHrik5
uyHlXKkMEivDNEV/1jl0T59sD8p9ExfhoWASd1xUJuAo0IU1QeJ/Gq/UgPvx
8WpUzQOYn9LRYOLiN0GtHtkipUejPBwpioF2XAj0ybSYYbDfU+ox1n8aVJMd
ocppxRVKIRciZAIMALt8M9s8LW/cwFhjhqUspEUr/DyKPDxf2guB0R0xM/SO
R8gr/Or2CQfcwooMjz89j1AHtn3C94XlnsIf6Ojq2h2pSMOOs1dHbZuWg7v/
VWOhAQpuTdrZAH9EQjx40dY+uw1vKKI7jhNhAnt6y5OT4CpPMyZPOW99bw5H
NUaVpMEHVS/7Ah73ebDGf30NA6HcY8hETEULcYnOrBDJHDmGAG/jKL/fzcWE
RbfPImQj/E/ljE83CXtTyBAYiaKL81XgPxzrHkZwflCVszMOq9h4cZaERr3G
3ilwLIDLlEf01k6d6NUKiayPRNb6P1/UKmZBZCEfMqDx6VAOL7tnuicFpQZa
Nq6JOxwCwS9yelH2Dqd0AL+jpbf+frdW95uJJ6it0gB5Yw0gT8L83d8UL/d+
QilQOvYqpCNFXxHW1ttgP+CPjAar+vQFP07Wgh3XQnqt76/szGBi5y7P1NBW
Hb97xkziJCV2y+qkoCzVBuaCdd3V1zPT8MaV8O+R5OpXwVkL05c3+5oIhLo7
5idA4VI3S4+XX53fBxf9jdSh8vZUkx6JlVj0527ItozLX5BvUBZNRM2bazxI
vZjd16/dAT/b8P6KkHBqp3wvOP+pl9I633BMVcrUQ24PfBNPRxAJxVBrPK1V
V9q1zODn9tnt7BVFQxhoiV0pYFWcLWUP1ngFZ0mW4M1T6XwtKDTZqZ0hQYW0
lNktNKxkz6YYDqarErd8tAXPxwhtVGMOckCX004vScPQj66AvSTBlROvI5Ti
iv6XCyIo2j/uOffjA1kHlI5bLOex2dgQ2xd3vvtfy/1Kz2e3mYxLcqfmNjsS
IfOm+w2Eh9B+NmF0V07VtLSwET702p7FVuhmKlrhtBnAgy52eIz7XxENzR7y
Hle201SGgg6EdF5NrnjGYgT5lvrSp8xSTkCMsP/QDf5E5VCRbtvkN1qVfWKx
PjKyRl7bPJBGQnzmAVnVyt2EdEk5dbt2Ht5NCwkxj+BQYh30yqn50uPay7+y
6ZPoTQIlXLDgdzCFYOaPtF33/QzjebJSF3/q2tC/SqamvuPhyxHBbguMrE98
4wI0DpU56JL9UpeG5c2+kSy2xZ1D6/f/PsKCuv0s/axKomEc5AdRbLnqxa/0
dNRSj0aKBu+qCDi1tGpOaoq7goAy3S5ymPMt3dAy/lPDY8aIbeIFwJp3rj0h
jyEC8p9LWdaGLIpR0iv0KHTYdi3Tv0ZDp++FlWPKVC3OBStONaMZpripQYdh
XZskVGUUWjjPUUa3UBqJLlPzgosl5VXnnp6JOo357NP/o4rUHEEVoiY3yoP3
PTa48BE3TUvMSsKvjZbYeWKc+CSz74NOuk8QGG1jM2u7nLlzevFR+jtsWEi6
C+CNdoalJu5CEkqToeKqyPrSwQXrdg3ZmqmFw/aV7mSDSDOdZhF2q63xnXsP
jTbPQkcHvy9O8A1CA5jjRiG7Fi4Z4RZMjESCdaqHgr4BfUGFYUUW8UmWVJ2w
+h/hNR6hmqZKgXNDQaMItPXRRKUmqhywa4AyU7nhStVHpUY8AgACrAzR8x3E
Fa2H17HQF8MdUhtAkwyzKLh1BjQt8dW1QdCQmNLsd1PtZubQ8nWX8VmUz6qu
mbnVZSXNAG0ph3OHgyP/zSSWkhwYvUZN7HT6RN/3k7kYkwam8Ci4ojwotMX+
8p+fI6EY5weT8OoRgJzASj0joVYHJuN8HZ+aGDjIqpZEgwxb6XdhMAKIq1dg
Sqv2MhL0jpNCzO4FCylU0Vu1ZGEXw1ODtLpWUMELnQ/izABQXy1wF3W7O9T5
ATlF27kq67oIDlQuXdz82Wtsi+tkvs3M9AAOeYxMJeaN8HBSgWMMd+OLqqBR
yi0d8/AkJmQWBq0SsUxpUHIsLL7J0xGjOFQCfJqd3Xq6OI7VKizpzKCRJyXf
S7FuudJycbGK54JhElU/oWutT89gArzhJmscidOVo0IW8TqixJJ/o3NKez9I
+wQGopGTBoPNzGlEOC9t5caSffF2wmYDucBK2frBfYLgWo1LAmCc/Dd/OBah
C9pzuEfjXmNf4ySC+JMsNrOzeoWqqDfln9x3Jezh/eKvQ9bpgyvUP+UCK+Zj
48F75U9KwnBnPtL15VXkuUVH4vrCASUXkEchT3sIYf4BmIWTd3AStYgrN8lp
kCJy1JIIrWN8RA+wBp3Ik3SsfTgnvpXSGDiLQO3+8jBfx+M3xUoWZBhIfILZ
jIEIsSKPMk4sbr8qWWEQuTIfCUSPLgAyk4KnxJjWUndcyTQOVHs5kuXsVX/z
mPPp1csfuXVo4QOaWlEI/kqDjzN5rlvqu5c1oVW3oYPtJUOQcSILTbdLeAum
Y5VSIVD3NqZOyq6cqEEmK2ofuu1zSaNiGAIF1myfJw8EV1lCXxAzBOuQ+EgA
yMSSkLKMlshJLEahQ4/7NKzF+6Q7GqISsFK0TZy8PpFh666yGM+QM3ChjnVy
Q501fR5fLBbQmm2Xu0gp3Sn3BWgoH+nqSNTrHZrT8hU5nCN580zDnlFVafHX
o1AFM8TJwGE4Djfjpq8OeEmuiWFnVTc6qBikzfQWXsFICowVIv2S5b0BT9p8
gQZBOe8DHRs70OmVvlFpNGqe4fnBf/2Pkq88kDkRqqGC2eGyc8MzbrR+V6S4
o2UpLMbN4K4hT2V5hrQxjtnQDc4y6E1QUVlb/oXMssJexTj2SPW44vY0xUgn
tdP4EehpqNqA6NjIKrqdaRG17e7G8Ac0dNWOHaqp/hO7dHgDm1c22xxnFJ6J
Fnrme+vzn8dclnC6z4XdDV8MDBxnx3YLVVFlSOsHvfdwr5pDqmuK0BuzJ5c3
TPxSoPhJ2khJi1cdqOybZ15qlg4O0bZjyaIU3z2fnf3umGa0UopJpDfosBTU
/8XBlHJbLdUYSKKlGPqV3oUThi9kzRVNO3vT6jU9vqXdg5Fw45jSxr2SYF4B
m28hhp88t6slf6vwxZhRbpMe8MNSi1BW1VtXlruswvOG/P3im5XDl6fK/crI
PZ8MsLyPrfZkViTUpIvUbhCnnoTtXmUXjpfuF7TkRlOtol2Gx6p+1roaTsl/
zTHCP2o47JU0mcjD2sMx9ru87mTuqjwzaCwQgcYNX/tyCnQwO32z4Ft5X5wh
1cj7n+EjIdvhFYsYcV3PvoQXK6IRyX4ELzwso73G/+Z3/aoX+q1WOpB6aJ7s
ezVnxmVbMZC3VSd+qMacWLwf9/T/sSSqGb+4L269OWc/+7WNuR0hArAOLnq3
K2Cz0lg6LLeA2UCtefcsCvtAfs7IsgxCFxPrHRAUw4OVjcsjwcmx9ztWxGf5
xFoCpem67W44nfD+mE0MeBwJ8gVKebk22v0MbDwpNczlti9zTiMd2B82dqyk
ZDI80ws3YUoTyw7VFw6a5vqw2C2A5GCegsAVJqZPtDDGchFJ/iI9i5gmEl8H
2wFtUQyPhqzAD5LzEHpC8z0obecogsd4x28JBo7DTaB3yX2948pXdm4qQIFf
qRRJcaJisjcb/90oUg6CVBl1f/7VoNqVSSLCJ2giZgywd5qHo29ptM22qgMc
i8tPqcye7TdoCmdQ61WyapmCPF/GqSJZr/Q1GZbLH2k/RywX6VBUFCRUiC8O
RzdzlQk0/FmAkbFpUT9DbZ1o4vitObuCSzxA2vdZDzPgthNK9u+DvSZPpZBz
6LXiViwFcnqAOKU4YdZJ66Qegx2oZW9QR13PQEJvMV+C7P7vAZ6ThMnlX/05
lmHjejcV8uGO2M/Tu8vWZmSvHtZudvD6dX+G9FYmfAVw2+6J7JccW15SWkDd
e8lPuXBPSAqYkaQxrc2eFYc0DZgpnZwptCPUR2GEg0OeVST8JpSLvPjCY5RQ
7qMVwu+nWCBzsNhurST2o7z7Gl0czhD+AptPt0PU5AJ6fycBDfpcN5I3zlL8
lTKNUJyJuzdmoCOo+u/q3dejx4TWwifFya/uqIpUhFJH1QD+6dYvhaJE9wb0
EA++qI/6tS3GUHLkxo4EZw0o62CbcwIZlzZYw3y3retOnb2zuqgcUwczQ85B
maOMcmcYg9WP9DHP5wRW45IoJT8q8pXWkN7XidSyfJ3CEPGd4Iw8ZzOrvZ2W
4mAq6RD1rSuULEXV4avr8gwea5R9+fw1+vlhu2Yo10d8qMzsSxUeuNzlP9n+
U1JmjXeRTu46WwvRhl0K2lCTempFaUxV2GTxF8dJJ/WQ9MyJNqGMlbabzahj
0Km89QxgeKFtWifkk4VOCoHW8JZoZtYkH3ub9WAcLPbHYRKp5OL+Cm1HS/qK
zOBzgKzNUafb8GiT4KBfVfjex4G15Sl39FaGPBWgPkxU2z81/n584IF+FO7u
wY5cjDn2HILUw2a8yDYS6Ev40so6GefM9LVfLBISAASMqRaetPv8AQJN+rqS
dRT+g4znhH1RYUZTBnXPHU6bNh9Bnf6Lj82lYacuwccBrE7iS/bacX7MiSnj
b9Zv7C3E32moeEsmBaOh1lySGkGYP6Dh+BcDskva3Fi7yOWZZuEd5MTXr5dA
AEkqMerHDkUgd3P7goLWbm2k4tEMeouEAFaS+USXCEL58sGn4fBztD82DFqi
JvvuOHxt8tzKUVRUuD825pxTzaU5BIpYTXKY/5Ay44bMrC2gPeFN7HZdHQGS
dHI2IdbUqpMa3lPAva8fMqyFQWdObGggLyqghARJo5E2F2EwT8gwS7nY+ADN
Ugjb0oca2Zw0Tqd3+SNw9mkLGzYK7yAmbeM84x622srcT2IieC3a5vemZoQe
GLuTKGds5oHNQcSSFv5qJSjGkLGDwYm5CC34I4fyAH+90/+zhEVCbzKZ72U9
meCztaY4glznRUwp/yahQQvuTV7nzvWFUbtPPtrLXToL6ohiKk/UIFBLBGwe
+7EQ0IsHVsjRm9RnL0yDL7wz150FWdWsJr49DGqmq9zK8/H93SqdShzpnNcc
aBYK+Rhcl7usTreOnE5ZddSxjKdXTdHHSTq0wEu8YFSH9Qpep8fHxAilI+ic
Ytbcs8upoi/dUq+X/UB1xsj1Jc/vt0x9S+QsZtVAi1Kes94lnobDdLqp1kE/
DIRv7nmOkNjrDNrf0eGw4/KbqkvL4TO7q1byx1ZG6wmFUUPm4Vo08vbUuhQB
8Ei/IqKKoxx2XiQlQxeAs4H7S8OP4JFBmtDc15QjvUararThtLLsLxgZNyi+
xiB506j0dYfTDNBjHzSplrb6EtIspHgn4tvJnn4TkWpLSAW1ej/6DnNdKO1X
FvcqNFd4+6s4A8Uu3HSvALCkYhad+apeUmnoQeGkj/BKCjYIkIO66+4UkdyY
nqAbivTOg9bZL9/rAaXIv6SASGG119bGhNSc0kE6Txfr+UOM755dc8DxjPsb
Ew1+GR/w+wn4fXV5LJtrbjgAB418BD357PRCo5FjKqAB+ZlGqubqlhASSi9e
UGwMwj7uGoXS8EbKhtUdCux5gPDaXYxDLzXOQwApcS4o+BKiAB2dfEkEwNc/
cKbSEXWPUZ1hPOl3gb5BJIKmqk1S86vT5cQ5LHlBUs8uPAJFq/zKwz060m2e
Ku/OesNnWDbf2ChV4fDiJ8lqJEH1GXvdOOUbU/ktGSKI5YuEd9lNx/nEHjVF
KwS5PpZQzs+31e91FieeoCE9RrnIpgPMuJ8FLSFTdDyBp95DPMd1X48I/qYd
9yqFpgRz2hIGd4AS/H95gVMOheJ3gEObEh6VOGqOI9G52EghMO+THeYr5Tk4
nfXdw2ayKKSb0sOyFz0s4TjSs1t1WxpXc7XdEBoZUMtZkcxxDkwXTX5snDba
kNzFFwtNiV0liqyYyTsCFg8xjYxfg7jddQdhwhQUQH0rj+nEz8J5hwRRV9mG
fbcVvvMnmtJvLVZcMLkTnFSFo0G2mwgX7A4mQM1FQKZf9Fyfjq1AgtH9biri
QEz+p0/WYfTaFBPK7XLTmUlQCZi73Zn3V3Xb4IfAb2aTc7ABk8q9okxAFeqE
+dP0Ddu6Wt5P9LKjrgQPXX25XCEwPoXExVkQ/cayjKFAlovgDeKAYoSfg8R3
6vE2apAoVLm+Ei0/a34JYKyLUW7+t/vVdgpxTNNrYw7m/YfXban3iviswjTM
CXLo475EiT4BIKSRxxAMMTtoPLipudBYqMddzkwcFDPTjfwXzudKDxh0pnsB
1YZkQGkDuPih3SWeumn9jlwksKWCidFAxBcrybOu//++7pwenEu1MOQSO9Rf
LS8i9wRHxkQlILrCsxZ91PG5+X8XUl6IlDrIvUTyziPaBfNd2YKfdta1NBgY
WIh/8kWDtYHZ+0sIB1/o2qKPVakmX3MB9ryJp6ZQyfLP7vD3h+/EJ7BZmEMY
63o2AoJHnhlrjlf4QLcXLwBPqe0iLmJI8OSyVNqW9N2qQQjCzYpr349lWtLY
sSiXTPUmzV5bcrnkxcPNh2q+4l90dLWrs6XB7grRDudPPOGvTVyVxyl57Ivt
dES6lvwfFjGJw8blkYUqCvp1afa2QWzhp48Kuf+lq47ZM0oM0qm3sERBfv+e
+NG1RpCCidorsY9xp61yzPuIvNn+fDvmY63kWlgJWP9T8d6pRMhW/P92TzV5
NB4KVA38fZgkykdvWl0Xq7hSW806af2OiE7eVS6c8AYskQabCfAT0FTRErjf
faCrsxTZAqDRdQssfvsJiwVKvNBUT5vA251WveOKPs6QVbNbcag+QAAlAiQ/
ngjWnq3lGRszI0NWGrgUugZn5Px8cz29b2KzWTkiWMgbUtixUs1uuUyh3xOe
/zKszg5d59tEUVuhnnlR2y1ppJocxciAM4/ECjGY9gzOYhTOe2jAIW+gWDpz
Ew5DJOO6cS1T6S2mx0rxcK1Q0KDZDnmLBXWEOGFkWMWrJayIxJ6xrxdmiHFi
qkEZLaGXq7/UdsxZsHNeaKYbdAdSF6Rx3G9TPm8QGvKK3B6vODFhOKPRVk6+
CoSviZxu1a/H5DtcAEkKMaHlcvrSUpMq5itblT0Z0EE0tOzFuG9Z1qaWlv/b
ioikv6QnMZcCTMuTUwGYcCBkmDEoeA5U7cEQgCjezA+OlMGaAHfvbGOxNxbi
4Wd+Pb9AmKna9yPeV8BhFrjcO4xht7xP+NMQhc+XPaUDSIaJEbiBr/jAlZd5
w+BtHdwPFzYRpN6yfos/9zoWZQCfei3JDguvVr0Zdg1TI7KjyBWLaUZF/qZm
rYQCfh8bci4t1WliQF7QJXHwmtZ4AP1ctNkdMb9zVqM4/QoRoVdBkFEXtusw
FzLG6VaQTYFTyNvUClJx7uFUaY+pyMnqw8UpsWosnbZLug9WRHaA2oGxyVhY
mQRdNJXPd6r9Xxs7NUXZ2VESMwXpzhmIRFtJkiSkCvEpccb1tmBMFXvRLtht
NZNuffGqHEJobyiLtIyWx4ZmDxcBwJ4Q5Sbe02/xD1BPohqYMQJvTJENKTd7
0wuL3/oJA7JcQRKnLcnJ+KOejpHiZ2GvTnjJ8W3fmtQ24mBRnAgM4Yj/PK8A
UpQ9rOtufYdruE5VGFy/ymqqtMJtxDRzxr3JxVnZWkfxRkTqIs7/lSSG13Nw
ZWfUN+GeNlIgpddMSmuEWru5GJwfo9KXEHp4e2iuSEQzpnSAQaLAtUP7xKS8
+p0lTswLgXKEJ+edjAPQ7gvTZzf3YsKfqM8ZadntkChlyeEnWe8jjYMTVBkp
cJG8sKtV9oTW+lBKw0csWDSPgFxr0Gxdt8TH9YDzQOBzKue6uyIvo1U6Vo5K
9cGNbbd5KiGeIraP68X75NRKulDN6BQmfWf78byzJk7eUnQsBMD0izumSZb5
Twgle0WDHhiC5fB78C4DTSDoFjkLL8uxo+T8GlAoPGa3bPy9aYPK8SK7Mtbi
Q/tdcjQMeTYat5i/szmqF6xw0YdMx6s/914jcYeQ8/wkN+DWvy79cxTv5soU
U0lP6Y3U6tz4w2/Qi4q/hssyfcZQX69ESWCZCsFBw8Igl9NQe+u/3Ns+S2c7
HR2LBONLKjiafLqQT3b6BaKmikCmb/FDx6RH0sWhJIos2BC9m/GSst8cxyj9
YlgZmNsduBntIdySZDkhmOXSgchlDgSjIBA5SfisYAsBktkY4VazLJnEV8x4
V1EH/xo/ljaIFtui/Xy2cVvKsl6ykJfB+ArOp4WNgFLBKRrD8+mZQnimvX2E
nNKSj44dTUqZuiLqIVbQe4TxokwhSYrNXZ2UxDai8zaSMmJ8o+Wj3JMrMQeR
apaUDp9F+0rXlzcQioYFZSZWZkJ0oedByStKse2wt8GB/asBsBivcoLlsWzK
BCnjJ/rb6BINltUV6MSoLO8XWHrkaVxxYj51gE9pmU8EWn9GTtzqL+cBkHBC
bpIIPd85G8yHSf51x1BmH0gLsJZ5Bn5WEzbiYLlK0AHg23e+6Ha28+rN5R3O
0t29LAaR07A6LuxMDCL/6OL9EXmsdWdbGZbA2FoNNrz+tShdRxIONiurJddC
QIDJIBIpqcqmEGJC0NvZl9DL2MdY5/8fw2QclsxooBFt7gEjxxUL9ghW4oyu
pOgLogvyKeoOPplM/+t/zailne4rA6QbtvrsC6s1bGS903etgPwcXU7Ap8T+
+U6F7m1YhDVNHO+/80F91Tv9srQMxv/ogrDzgA+8AKq7rBjYwbPe1ee1t0s2
KgCt+rUXPodkfG+vz7bDH8BjZTBcWhBjIWzz1Yg3eEWW3KGvzn6RjoIGgkmT
XYBKKjyAjrXX3rf5bsuJ63FwMUgJydXVmGO1G+xKFcmyir9XWJux6dhZ6E1E
IEYo5m9W5bljI8DcyeppRNwvTDRVE+i494iqiQfr84lnp3sbmw1rWTMpe3j9
c0Ih5JL6dUVLP/mcClOqk9CYsm8EtUyqVWutM0TdpKY1hyoCKCEH1nJxtzTX
pdQdFycFNOWwiv0UYdlESIih79e/rnEja5SOPxiUHSaQFT375HoWTznoIL0t
ZSaNsU3YjYQ+uRPtL1+WmvYnSMaxgSVVdHFHmHrXKTMK8pCS/ukB8nnb64T0
tzHKoWRaDvuONJAFpfIP5XJ9ckgx/UqO2/usvwlzJxeaw/HuZnzvpgmiYXGF
7orRgWQJ26cAPbRVjig4Q5Got6YrO33HO7h9FbuXB7x8OX1otA4ANKkhiHTC
7U2hrVBADDl8boD2SzmS2jNIS3mgR400aE4mXFCGPEw+HJ6tQmVv7kTaOOjg
6rmE3fQiSWOpnXBo3raOFtxyx3vxwL4tN3kMy8a9DIiQ34LaNHYBy3uiM4TO
j3vl2lb0xJQsObUhqk5OMGCJzPlt/z/Tnb4DepuSzvES2AD/N3DWJRkZ1tsa
CIAmkOaTJWvM2nfW9JvXMa5+6xghVVLmvQuTThCNtGCH68VZd13MxgaNbcHM
INaKgMWjxHWjOMFkUk/+3zBj3GQ93C6NNgW7yXqNveT2tES/BlhlPhgou2gr
L3gJZvBm20QPDiCqc72cDkDIETgFySNuL4Z4YpTG/dybqOJvr9oqx1i1YQyl
l4c+IoxRVlqmqkazzJjTPcvfnGyNsyeL6uOxye1UCdfMPO9szLyIxZcqU4/w
fE71MoVm0F2mJKe1rmgL7fdi8uR8RecpIBuWee6Y8emXnwTL0imnMH2ZDA65
mUv33m656CYw9qTdc9zUzWVMekgsj7Cf84wvd2sOnhNZ9p9WEp13aumTUAvZ
IAELng3WfJv0+fhnbPB3/OZ6xzP0KgKbCRojhQFR+bsakm6G7txBWUAuD9M/
xzF1og1oKhOBA0aU7imNSgS7+yYcjNDOnCWrNrfgIBFPceD7Acn5DVYP4xyj
ck4lo9JY8xjtqyyo+pBMIz6rrJidkdeYiKF+vsqG2YzbL5BeglX+nxPJ5DFH
+OMJPDvzuwSR8d89ZV7tW2iGcps3wLwuZN5B8E7rcbBXFyicz+saeXtL9sE1
wbCmwdi2NncAzZ6k4y1h5pbzsjfs6MRStzn0EovUW7BGtHkydqz3o80ZdA8z
h1Oa2eG5Y7IIQ0a9lx1AKjtcP5LBu0kGwl4X50CEremZBRep1kIM3uJfObTc
9/A5E6FcWoEnS6DUqCkUd91kVJE7KWRE46xSZWmq4BqD8+8bJYM2naINPJae
CCx32eO0CsslD8uP+eWNcL74bv/jg3qK2molp5APzVbxDpjXX8K/YDrV5FV1
agq+Uv1avam3zjPOYJpNZO5hN68EzsDCuZoH3WhISsBrsw4r8dXzqsVGxagp
2s/8Qgg5vkwKGlluK0rV+uWjnDOF2YfJDzjwjUkBTfsbFOnr8JJK15to6Wyb
QrQEBXKVYT7bSm8OyuRihd6ekVYRX5NgPm1xQGYS7egY1aS7/sY/ZCHVOCuj
1GDO1QpEPsQmsju99Wt3SdpX8L02AitAxcA3eylDCibGD0Q6PJUD9Vttny9D
A4PFLJEiWEZzq92r51KCVzfYWzABgkmytg94fUKhP9VPmgXNgrVu59lhCr2G
ZUhi2CNQIUxrnvwB03FcgIhGLmPWu7v/F2g1VFUqrzRVu2rSEBTKuq7XfHvZ
HYHzJBrgal2dZqEhXqOUQM+jYSHTLpbYJW0AbAQ9/lfeSLb/NvvhuXvlXset
+dp6V8RXWUt4j14wS1HTls/vCXwE3UrFhEEXaiGjRHG+mBtjrJDcYCp8cDTA
Lo9DkKgr/9YaCOXz4nNqaxHdLBN6gtIfNPP99AOyO1ql8oT84ejyzetqL5HQ
7+HED3lir9vd0PzD+wYjoqg9CNDfvyZEwRdPv9oUnI9GkGtd7Cky8lURfpAJ
RmGXku1BuO0pFY8LVDZ1NV8zOvXM5C0J37Fof1Gua1FRWAKK6PPWS4z7/Q7P
MfJi7nk2slbNL197EbcmRNRb3vTJzqDvBAIXU86dHSs4hqN6UupL42uRARWY
wlxvn3WLSqLAm+jcKYooK6maAJ8utC5GQ4N/ZhTf4vKPfqnZB6Hp9eHlfOC7
A5GBljhaRp5+N/K0r6hUZ2xeCG2SMXzDwPrwLUl5YaIj7fnr9TF2lCsjh08D
iBksEYbXNDdMcNi84hwFA2a+Xsyzw8oPBvRaRuJwjRUyHyNRGmn58F/sGZbN
u69c47iEFslaX+OET5bAvRy7DIs/cHp3uBOMPl6akuzvIJ34Wg22MFPK9jZ4
LWBrc7xbhX9QhWH8dVA3WmxbJEpFA3ZrCBROdLL1m1DQmURmYY39Ovhxi0xR
zGVGCX70QqBhhSA5pu/Ynk36LB7gAaZywrsmtT3UVe2DGSfyx75p/7nVv6hb
wNjYxERjaDkCaViavqZwX2OIKCizQd6kXev1UHmHhHnj0WrnFGQ8wFzA1i3u
jCa773jNxE+zNRD9YTnVe25EQCwL+l6pFYdrTMnuWBpEA400782Ly2rU54Ih
Wp4XtzC0JwHsOITtO8wqPOTGI0ErakNJp1jSghhHsOPWGe6vXnlEym/srsK+
sF0/DueM5R5JyhhKq4PJNjwtip99KA3lqUAGQdkZC2E7mE1LuLriNUAq6GS2
Ajs+ru24+4qrVpfrcIOs+z0pcM8LWoQwb+6JT7TFGiKHXBUNIvQij+lyEQT0
cN2CzBqEf0j4veUhIfASlXqwErNOxqtnTeY9k54am+ibR/Cl8AceGzQyTf5y
JDT4h2DTVkNOiyOa9aonhGiUkGsNPvBrtm9nz6ixSshd+QLjKYr/s15wnFCx
QbzThQ8qA0MfCujSerDqUjsVj15hEk0gbLVoQDDop40WvY0EK6tCEa20hmnL
aAEgub2nCtoxWp6JAxuzjObd6QaeW62Fdb2u3jYsQhz0K1DQChngFRU+fJk5
6/F/Dt9yd8BSsR9YhAVQCaO1/wydByhmHvRDEuv3ke1wGWtt+LbevasLcK9q
1WrjIJ9vfjHJXnZozq+IcH1I4nh90lCkLYYT1p/07XHnKs2Zeh7820Z1tnNa
HzWT4MUmIiQd0lYgyxQTGOxZIUtOhpYZbURut9+l8mqFslXjaWcOtIWgvnlj
pfBwhvrQ6dRbyE1FTeaFHp5tdFMIIaH/3LFoffxaE3BD7UErleo/2Xr6zMEu
WbHpSvjDx1l+MWnMkUzzB4WlzsAkOD5WuPZyYYqc7kT3678mp4fqw+l1coYp
7q3K+0mpR6liQOZ+BJauOlU1jAzA2w5MFJbb+6s5xGSs3q0qPiBZ7tc/0iDs
kduTJXhqpVx2AEiorRT89HRYlSMjlRIKNZt91GOPm/imXOBOyjLx6Pg888z+
6aP4YAxwcQQzinRse/Yew8dpbiEOpJMcrI/LG8BKfMM+GpA9ZaOb64du0Pn6
LDmX3Pr2zhcRYwci2fiESwBQU9/8pnomZSAN5et+Q+Ff99ZxmuBL16qSCtkQ
bYnqgb8eq0zFC06OnlOmRRHfbxElIfjwUR16E9zF/ZMYEp16CA+UrpXe577p
G1sKeyzfJFeRxz6CmBAlRUAAHGO76k9nFlp8KSeqJOLBxOE8ldfa8UWdj0dM
8QQny7imihATQX1Yo8ur9eTBHyRRXO3DRvdKrl2AXq/tWeteRqhmBnFCfmt6
VMWycqilS84D0664fKiMGTDT+aK7/so11gHD+fDrLbd2XJAx8/fnv9I/FslX
i83IlNPsYlSh72B75dGySkMgWBbR95OAi1JfMexFrOAfn8d3xOU7BZs6Zya2
SAaxG65sdGKSY4w9OUmzUQ1owk6Yj4tzgOnO0BLknnmSVoaAjkNf8uIzThyY
ITo4w5cQw+NaxNc4E1tHVAjLwKf2o6Edc/Yql7s+YcYevfRpT9LuJXf6hB6q
TKNTUl2R6uCNX1lqz4dmIcWTRTt2Y78M0JeY+UUARIE23o6lFOrwPWejG3bh
VSk/iPcPLGWv7swFKIygHsoPq5DuakB8S5hYSzRK0XnW28D8g+k1000zp9lr
cSeT4k8fqoO7t74fFfzVEnPobaZJksfc7+2q7urem7fU7QIu4R7Zun3ufZDk
NsNFiA51uhJPJZYkrlsCeSZ0B4oYCjABcEKx72KRFbnTv6wusqysvTwxNsny
35FWZVlOj6PhmhpAnBevgWSfybc2jfCgDz9ulfaEgcc/yuWwNC63qqOBKwq3
oo8EmNulrXWb8Ba8wi0cJb9UU2445stZy4ZUZmeiMLf6NAzs7FmQ/MgycGiD
bInwx3xf/KK2J6aRUSxKQmxyA4l1FeiCiVOl0qQCspBgPpKGNqm20rKprQaH
sa51/+h1ZQ81b7jfvzoHn32QcvfYywSILyBFL3r8fSuhtkd1kpHvEsHVhw40
QfHTZQFO0OxPVBfD5PBUKVZKu8txrrYByYppEktsQOZDx5zultUI+O/qVOR9
g6ISOdJE1vJ+Jk3NhRZMNTNGBWCqJNq7/OfgIFQQ/W4b7KyRyCKTkhrHWB+o
FZc5GL8Ivgia8CpOzIXzJNuy9jkn2mWJdP7YeMZ9L1DX718/df6fQ20Dkw60
iSjtSN+NyQfK4IRziJ4Mh3UKEz7Nbn/+ptZK9t1J91wKzbFH/hmhAKS2d0rq
28wJT6tz+5hzfKi9IeoFPsX5kmVAl5kfqqO/RQxPpeGMlj4NZPJ1EL27zMMu
oxuCd26Sf9kxq4qLuaubACXgdYrxk0vK4NzRTLXEvkubPmXmBkRqEhs4zbdo
mfB55pK347FH0KTc6CIQP9tGmbaMVhqXYoPAFu6KL8wpi0k9XOueuM1UT093
CdYJVtPzMldmlG/wATH5BE6Qd00P7v/WTAGAIUZzZgIYgNgHSdp+4BM+8FG+
JrdV4a7coO8Ao97XAgfLilOFG1y8JBcM1VG9vNAzHcFYLW+juoZ72C8MwcKb
Hz2G1zbCGSZjwwr+lynx0RfSjDq1JXe9UbA2jx2BRU/jkOIz2eTYC6ZQTBI0
b/0wNRN2m+O9Wi+5YOLiVk+ok5PxUTqyLeNn1OzJ6FBcOPuvnokn1zwCFHPQ
u6123WYjc54V0Kt0XaHY9PTY+eztOawHfbxYmw28jH+/be22KydR8aWOuFis
Cfh/Kloy2zIf5x1wEDCMYil+DqoyaQkXd9uq8ihkEpY/+dSlvApUKxfvwcfJ
eiNJHwDncG4AI9E79fOpKRQU1wEn0Pmn+2YcwCldfhPq4WJhd4JRqimOKQ8k
bHiyF0bsXxdn0BJlpbdujeOLjIKuJzgu0CDz394IVR5+/SwlKqPX2WEUDYcm
6F80yG50SdBNXW2WvQ/emQzrVkRJ8aQ2f53VyaRQKwMhupGpedJC/B9E2hiZ
mC0yoY+ds66S5QQkoi9V5Zq2TH6AX4Kt8B2PfdfEdSXKa17iGmC26icpkuFL
I3HNkl+N5g1y2GJWa/hxou3ukzAtiwhjQKwO8T4gvu27iOVV5Gha1N/rjkH1
H/NzN2LByGAwOcgH9UMjN3Oa3gbms4u/hX2x0KuJ1wpAqVpBzHn0c1y4gKBG
EaCSJmC5HH1BNgSQQxtf8iX8OexPVgh3USXbN0u4W4kkyuhdkiJ0Uy35BceR
kw+x7CG/lRItkrmSkdDT3Lk/gtI0USX+avoWJmnVCPd+2/Ssak3FqzAYf6o7
ke1B2cJ9uu6jZRFZsWvM/c/5ffJ9Mv/UbOukutKTWYK5ZOon7HT3sGZ2O9O4
6maoHU01/ZwxOj1TuA26M6AF0OzMrzTJ5j5iMrgAyqiyBVvczIpTq4OsOst8
g60A/SashSphZunsk8C/oaf2iVTLNCuvV9Rdf/2y3u2hAOeDtExk3zQ3cWkM
LbyXiWZ4yEEaYRdC68Te/sRvlgeHOhKL5oD9Gt39wI0R5QEQg92+B5v86aP8
9YjK3DO+azsPhYmT5nc3+HNsgLRHIQK1JG06aRNaZHZAHz/xbIgfP2XHXTtH
OJDFKBvD3yRN4wcNUtWAVgk8O3K934Jjv96IghWNsPBTBvqbcjowc+RIWg4y
9/J6zJEO61Zj81jNCSsaIKsNj7Yrx6CSmJPXeOeP7FZvrlxieIWGFvkvK4yu
os6o5KwUiDeVDwu4EUYHGfMnhCQtEiVlFaf7pu4MIQ5DCOUeXSZwE0BJanB6
qCpK+DRJqGhGWNruaDwyTO3lWXfINlFBl5VOUq3ETb7cYfqWaIM8QIFQpxFi
DbTaBe18sAaXU9IGzvyVlU8hwno+zbOriUGTuacCyJFuqg6C1wOGIKWdZYrD
jiJa1B4TKUlvNsruaKpKicwbYMY//2boRH8va9Ou8EkBOME/q0bI0U0OENpm
RmP4ErIxEKmruCPtziAhjzPxeYfuWiTPG2UfWuXSnqR2voe467FC0KGHiylF
aovXz0/skKGjkVqi2Gt+CbzsX5yBDvGBS8tNbeGJ3Bo7g3zkGwdH8r4/iZyG
zARX21ugDElzhJ1E6AkgSHl8ueNOpROT9+KekKF+5VZiz6HCfW/H/5e6UWKb
qy2Gc2mBU/O/EPNKbKa6V/Pd7lqbLd2b1GeGSY0kfNjldEjRervVaCUYdmc4
nuJ9mQ0+fIVbm4GUGf22Hm69r1KxXSFVophmif5zsFMDAM1ZGePiZewP9ee2
/StUoN2Z/gde8G5cGtOmSviNRBrnJjR5Pk64NQECQk5A7/UEEqnjabPCAvPE
LX2TYesMC80lZ6LVnzKkPknU+qG1b7d88s3EMIoFRPAYCJHSXhe9HWmfnjCb
NayNRCKAhwmVD23hhd1x/ZKtCbVR6Sqfh3Pqv4IsQOpn9tOzAIXHyI7a4Qn0
mIhupcpLmrG8D6Gwc3zytcUwjkFuS0ttKeg0Z6O/8x1FfDIcCd11PJoZuF9D
SIY8nRtw0gQz2MlvWg5gegGFzqn63mYolnKwhuRHVLHtOQi0PDMHTHkjAapN
nEe4zPuViOPbLYQ+2mnnNrCNnlwXSRMF1lMR9Al+VyubrM6LxTTxgm1zKMrl
g/EjlLeokZ/I2lQ8tCGK17ARauF7+XtTHjWGa3bZ2ZzKmnLsjzqjwaW35DRd
mo8lb38NaXsLkSR4Iomay4+60XuZco7PrOMHIF10fay43CEdSRlnBtFC2R85
6awC2qfNQk5zqvVSdEVZ1l+SzrKHX3FbMy8q7HbkUvl10qcwHECM2/taSIvd
X6Zj2ybJotNj025LGhwkT7Men5KjiZ+/JnTassk5P8+3Rt51rnZE02zzdXMm
m99Qt/dCSysTeZ5gLuvBOLAupjVb6/b5MlULTsmr3q3Ps+De2Y2CEESCjCnw
/mA1IWzZrgOd7DzFbp2NfHB/4Rw7Zqs/hCkks+0qPXqeeu6A7g/wSmdUQaWH
5c3s7+liRG8dM5qgRiym1acgl7RUYtBrtsArb5qL7JdsBsm1RNxT8rdtGkTB
golcpZL08LGGmzx2Ob0awPdMtYi4gHhP92+pJ+2SYzTYxFhTdKuTLDWixqNf
Jdv3lSZ+PXB1ah09TPhcjzx1llW41KvuPxd2fq74oj6qNLBHffq3OKm2uHce
L4ycFZbgZ9/abh5zXpeOmSUiyYOCT6BRoaIOefi7iaIC2tMKJNWiYgQMPFsr
HnryJSdKnyWsUFngUCRAHWaqLan+KLZg/CQ7Jb51VpfKr5BXSNOdekdOgZ80
gUMLdcAOMzRe3isFJTycR+/KyhTsfMdvwIbVBFNtZ6ZRl+ug7gdVC2lsqtHP
LB+fY6mPsV4Wtk/vd9xTylKq85z6VOZFvPr47nFnMkaB8xya5p7FrhUCRhQ4
UQM5UjMfRqVYVaEyz9xetk3hRP3YLCZeDGBU9WAlGBGkvCFTjKR8j8sF/Qub
E8sp7Eao52+EWFMLnrlfk2jl6EOeOnLKdgX+JVXl9fobA9ZlKvUTJ1ijXrrp
LN2t9qgqXxY10kSoXO1rnZAWt8FrOu+2e1RURYMnW309+N8pAKDUrNX+JTuT
JBGIcXCxu0RAQhOXXbvuHYyG2UxrujJ7gfMIBE21bJEAK5QLMSLVi3pLnMTO
NI3H6+hZHx1NnhJkg34mgz6sZVV4Anq44ruCmW9gVSYxr0Vs6vfdv2g0ULgB
PDuWJ0Pe/nPOgB8VKASkCNgMWsfQC1UM42jivxeaTON2u+ZybYHPG3xs4C9k
bV7H0uyJX65RFfZo/hSr9zxwqt0JHPF9LYg2WM79V+tPYU4hNL/rpYGb6IcC
7ocm/Vnk1pBVDZCgXO+fdqAmcfKqeXNHRHwz5cXlh7MpbkJPZaP/ZeH+dMtb
+npydtrL7zTSuVYjCoOw0gKwHI6SlAA+Yt56HqKQdy66ORuLwZWRR5WOh64M
mJ4WzdEF0SojIXBlOAHSlonnFzmje0VSJ2yLmTTTsfXanakoPK243yhxcorw
o2O/QEOBxZKeNmzh+aiYV/D4PGzg93iv9Tto4pq8J62hVAxE60PahbWHiG4n
rgTAFWeVyfdD/MxQLxAz4EpIIsKJccfbmsN8sCEzyZ98ZXDH4sTL+pDeCXvN
ZNpK2shq6dXPLLOnnpH8wCUEoYrBmWMgOaOwTfMxsrmIPE4r4cGWnUTA9uw9
S8cLJtLB58NZ3l2Hk7OFfPl9lu4p4t9DJMCP9/ewQfRBkFiqe5Dlwv8NiodR
+nHZtQRKG12WO4lM0Ay6zkADxy3KZ7gV4SOOGQuTh983qlej2M+eTggnGuMW
M0bz4jflric1xB1tAN02mdWfbfxx3SB2ZzmsVt/YS9EQ4qMuhzlVdVSjT+Ob
OXiPzL1Krot2pk6W5O7nFCZewJTvE9mirmwQ4ewvI6ATHbda7P1AycCNKPse
qUyDmkLT/dDkX33P7Qkj/Cyu2RzM3kgE51PiAK/fcKfSV5d5BTJsdVSMFRR0
3SG+tBtbHsgyvbtE7yyoDkCsqzs5GUxH0MDSB5G8RxFFJtpZCIQkATqh3K8S
8QNJqrBqr5U6Ug1P45Vt2hs3je3wDskQe9cC/jZM8FE8S/5P5hkdDvaewgvl
LgFi1zxzDEZ6ZTUIyKfzPG7qIQQ6UuVp+JfmBJYAa9VlADsCNNAF/YA2AGxD
To3+vZnILWG/I2ZQLp45Kh1whqo0PSXPOEbj5P/BeAagz/NyrLCiR6iqFCsg
0wzxDvmOqLTJwvH7DEh3rnJYdd2wTt4jr7AQ6v9t2AZGJVeqebJnYJEbwPvV
oua/DsmXsbhBSUpY2UTZo+9x0qRA9PKgTlm+Lg7IScgVkmR5Nud7LS3oJyJ7
vNukR87gssyveoPaIFOJKInN2FGYDYTpReM8SLMlLMlmn34d04Yc8ifwd5eM
U5nxv4IiRs02OREJq5gqQEHGDH2a14EAMOflU5+QiWB3kFqwG9WWyzczlzIz
lylrH42JuQnZWzW4hfv+ivWySPPqsNtbQlKqSwInJvyqkqRGJyR6DFTVY3yw
p8AqaCoZQA7vix3Yf6X6L0S0wTFuEmciVrsjDGlRyZz3v7Y8H8oPp4OU6PAE
1zqPCBpb/CCe8HbU3YtLj3Y4SPqcH+W6FiH37hW2Mg7XgiQjHCOlhwfZNqhP
csSn4u0vtMJJ3LwGkpFimjFtrI7gr+N8opbMVrJCUMFwClCBon8umJG2LXqM
HcfdIBSV9AO/ILyeMccHahVxgS+NgVWKXiIFkel0rGR4tFCQFnBd73TIukis
Vt/QqPVSpq06MTbNm6SRaQWUxEBM0pR0z/pV0ymdaM9jelATYnVQzrCTHGPi
xsRur2KSQiSqVHSDh7nHAOF/xO03rMTKbcy0wzLiNUh2Ooobk9pbWmOm1KOD
p2pWli3xdIwWG1Cw/9A1UOoOGe/UYIWRhFO6WIfNDOoue+A6uoNEuCjyhfgt
kryqn6gn5qRcbUCy9RM93ublH+J0gD2XdK3HHD0EIlOMMmuBy9HdtQEPfqHK
DEOm0so0S2S5IoGjOnz1M1hNBci6BO4nIfxebBE5Olss1+IHtNAawANiTmap
s+ojqUv02A1sNWvy4gxZogt7+pXT/k/vgy/YiPQtQHp0bMFvsKfV7AiUNQWW
JBiTOvEnc8LfTSX69e5f73CpS41S/ijJ3anLRScVGr4wIsaAee54ldVALweW
J117wPEOuE8T0CdyrqsgL8QlablFiJu8zDSGYC+lHIZwFIEk3Rnf2nZs8HTw
BeVYrkwnPRr9WQdt5DcaNvNNG4v416ySFFRNsJwg2uekexRDGMb9vqtXidDB
3XaGukHqMjEdh7KpLewHWSQtQqFucGYnk/0A9M1CId4yiKy47QxHSWKIH9xV
TeAWd+FV4BL5kQve+fi/IzbOUApywIWbJ9b8q4xYMS3EztN33BQLXZo3ct7e
xsrLuZDvSwr2vNb/iytYWEMt41fteNTW9FXv7p01BJrjcwEdNxfRmHF6B/c3
5syRC4AIfv4m4d6HUU556o7sfyhlDKat1QWPdigl3WUmByEOV/DKXtHbxrje
8LVUD/OFYz9OULCTy7UA/xc8zXIMC7jk2f4SD/KDX8EPi0LUYmeUwbpW2Nev
5ONInIHnSGDm+W0/LkhdyiAerTuoPbtde8sU08/LBUO2y1BWQMKRlMJ0ivBS
nPU/wx8umzBIN4toaBGxSbndqFiK2ndtIQrj6hQWJ4C1WDYPQQIrhnr2SoE0
/Oap3UodbPQfdr/XQnpm3sA/QMZdn7BL6+1Ojx9XFOzsrsznagndJSBR7rjE
WvUyb2Cv9uo7bjmtITKwU8npLC7djXvQXNF37ZsVosRN+CRJ+w7osn1U45ho
UoDiklo02eF6tn3OtfU3Lhy6ASRzOPril813CjMoSC2h086Qd3x5zwgY6zkG
GNsbyjgiNoPoEPGaZQql+M/A6aYh0q6YvkJn6dRBJTVG5cuaAvkv45cHEsOj
0UgeIJ4HGFv2JjpdBPHURwgjIi+mHlCU1YeI9VdoWvktH1A5gfsBHBqy80ow
Qg9huftQvmqq3r6lPE3HCMKUsVy8UPB32XWbvr5hfP4eNeiZeiunLvGqsGnS
wj8U7W8A4DU7wEus66Kj2keeE+DuZJUnaIciOLpbJowguL6h9SmAoXn2Wn9y
K41raiWQzK4RLKrIBu5ATMWK82UAeVxeNvyrfSTC4UCu1qiiZVM4GJQBh/I5
b6XrO8AHY3JQVAF63RL6wvcnxFUsjfmucNVcDLl7trxkDObDHGwwx2BtqMSK
lpd4p/N5N52sKfuEQuQWpbFoYaRgWo8DMOMPASZ7iH2VDHhXsoDeYB7qiqPw
dYX4JFPODZxRmLQ7GGK0kPkha35Oii1DQr+ZPrx8dws1bFsoJh35jN/BSGAe
Qhsn7EnQgdEurgRP3GgQ+GYSXprgB0Hi3KQ4JWibGGqP6bYoOMtiCxs28iUw
nG2iyqYurjqdRVQs8jiolnk9fS//mAr9ys0onBQDWKLxeHVwyTDo9AyXV8XN
lK6B+l3XocjDEDrn9ii5rtfC52T+z7NP9tbqH05kqSU529a/krbnlDvwd9I9
y7W0MQmSFXTM5dbn85Cu/s5tLdNOVZA+m1gx9H7m7fmyq1tZuv7op2y6nq1u
VFBbiBMZrZUf+SDm4CerEL1IbZAlIutCN0fSgMqcdw90Ro7iDFKC+z29+h51
v51bvB8ZfqReFgtIIUrBggYjDJrYp6YdXqH9OQvnFVFtUbHBezztVv6sJHPg
MCPw3+0kVxXJHzj3SKc/Ub9EFeFmxQ5xybWsPYGE9ZXxO350IJy6M9rGoFfd
W0JT98XpHmmK1tTk4rxyZvX7Sq0eOlNKsTvXqK+bJyAHN+PyLshFEeHkgYbW
uKxhNR27Qpu3L+Yprk6aTDiX+p4FKoVskGMlGp0UiWeDRLNn4mnNTVk5cZm7
Y1tDN6D5+HUxNu5fMXW2LBKfWlpEMk8TMbRWTCObfvJi1IOzhtgrXB7mVTS6
BmMoNTRa1tjjOaIabO1qY+2e1R3XOdeCBVVXOecnTIIKFrtT8x8sd3WejK8E
naxXD7V4DrsjpqLOsFN7Lk4OtvVRFfnX0Z3RsE2eAZizfEnKrJTJ6GGhR6pi
7lhSf2ktk50qSFRsMlh3bPOIue4xprU0IwLzEa3h2BQ1yD+YdKoUwOsgVVjT
4SAhNhTYDfrDvDO6DboMjz6B28p7H/lT8i1MFg9v+/auiayJV8bJWooNcz+q
RkPMb5JmPkpG6IfZVZuS44odi6mgJchAnl9KbffYVsinHevHz+mYlh6TBIyo
Sxpjb2G/IjM5FshF768+8+ulmDPMSLH2Ijm7NAw47ulwBXcCDxaum5wXbWKX
TwjkbwYlEi/6sxlTl03vK5/V8eSakeiMU1AP7aSN0s5WOr3k8XngYnBDStzn
iQfzQPQD4t87WUpSNksTybYFz+L2og7iSE63+hzI2Ac1xlb0YXNmTpYYo4kM
X1hIHOZOYvX6bxCG8S11lpZ4GnKc+60ZsaZW1dfTO897RCxGwNbcX5zpT3dQ
5wvYuYy3tLJijOIKwig6E8Ro3KEmdK5SStRhggEI+1lXhjnQNbdSd2TOsjNZ
LFmy0ksqwzLXVy3V692Ib1yYzb1n814YkKWme6XMUtd8y4ItVWWz36XdHY0n
y2T4Ay8jD8+VnhrHE1XlLdz9jz3HKdHVjd/1EJEBwrSXhvS7Ll6pvvvmBaQt
op1I4psSYfhlFEWZbQbm4n9mp9O4P+l4DOCTmzoSob6KqHTW6QhiYLD46kLw
krinjudvKBFrHDiu3Ankh0hgl+iNU+4MWjWUcVF7HCE3xE1e4VPY3TtV2hE5
7bcQ5jLqQe6Z9xEcBLjRSRGVJxwCR31OJlHg5yGo+6M+/mPmR627mJ98c+RK
6IG9IP6tQb3ktEttMicWWqTBrFM0XW0C5uQB5m6jKoDkMH408CrVcU05Ue2e
7EcachaOt8fVVhQUwEwQDhN24ERRtehhv/fAu6UOwzy73AH/pVmHNTtjn/nl
Kq2SkTLgHN6p3TDCVhlnN9fGynBP0PE0j0CXmMZk3oz2SmrbXv4IPvBThjw/
fzZklyAUMKXnPlxsRjSQWrVsNptdki83GfXuYuuax4dUwTgtd6eN2mBwl/fm
LywuvY0l5XKGGAK1nWtz88GsV2OZDf1Yygk6F+0jF40q2cPzaLtK50aH7F5b
9tSQ/VSQ+QA4MxNd7mSyU9UtykdNWw7o3SgXCbnMHb80P0SWnj6LkhEbhk62
Af7WUqHcf0Czt6ww1b66M7EzzCJQMuCKS9dectvgR+jKrAcvixnl6pAvNQCu
RNP0QpUpaSG4QblBMHEb1oXmUYE/MXZT5GHWURPMtwSupPfL5J8D0JFv/iI7
rmPb2gigQwP6+j3ih8YUOrHBrmbOkgISz27N+Z6wNQGtsjHTwr/wVRAMZu4U
t4Ke596PXGPCQEL9o2S1JdhtS3Q2AWXSa+MA/ztv8UmjCIipr5bYbNsrAZ3b
DkJIA489OVVS9SlfVkrS3TJ+GHf0nNy2nNlk4FGuFrA1k7INYgzYitdXvhgg
qOkg+PyK47vzjhqxayEPTeraQSJqLzkelu8QNtpClbC7HdptBK6rf875jVBY
+1AUdtkP3kOpMYSfZuady8EhtVDzdVwF2GoLiowSDzQqn/CHo2BFmWBokWQz
yq9/LJPlxWMn1Ix/VRUrYHRu8DF46Qxe4ipXAzlVWowgjEUOe3Giopps1G6g
+e320u9cFzn3+Hhf60D1wc2s29hT/ykcx18nwR/BM40rUz2R8NunSYG5Zm3y
UrQ9IQjeZzG9G65TJ+uifc7mou0qYTJPVZWNm2Qq0fTeohSjzijm2GxkjqdN
gIxC3iCgbtoLc24btdNYF76u/Hw2c8bAHT8B1Nxm7XBozhI4CoKJi/abJutb
ej+/ty50KGRkfSnA+TpZY/kdYVScFJuwH5OndrP3FllERWItHMFl8k+lUaL+
IEk7z4ynRcB1q3aJBDWDuYSV16kdC1b9ALpupsnXxYeqEW17OplMCrx2lOOX
j/xYFdoHAkzU52UaUAuW585FWHnMmMp156soTMdcFd1FzwNjSEcAtL7FogEo
zWOeH7Clgg/5TJulpG049B27GkW7B5+CN3NPqv8ef7dCTbaDu11xSM0g+Mwf
UU1534hwEdvrH5EYJ1SmThTBI/+zdvtTj7pyfgkE9ix8G1VxAHW8pvs3I3hb
xnndHLEHVXaV+18zWYjIQx5UoXyw/q4oAYzUnbug1POx7ch67Q627+WUzGFF
tQVQct3hUNicFf6vhGnaaNlll2NuDqWgpR9SezBu5j7DePXbbVoiCJQKOhkp
4hRvdtNB/D8xjSeyzp6TSPbzn2H7A20TIMZTZJnBR5bKylmu0em+BhZF3yTR
IWubLajoS1J+uui/9/JHTniFXlfWxLaTZ0o8pOegomGoMVvDsm5XJ6KbSCqp
T/sIMABg61v5P5I6L7MrPo3Qz0PEkFa/UiRCNyop+JnK5lViizjXGgfTOERX
fYJc1lte3qo8Xh8O4QVoQ8pShPxv+/Ua2QD/M49hY4N6t5hUuPSee+ONwLdS
QglmMgHHkWJRsxaKTE0PmNjwRW5fskn0MI1H7W5Mp8WxSsz4tCz/Dl71ge/w
NFbnkMLKK8fwBGghK6pTpjLD0CnPKrUJsNGFhisOHopWIz2F0X0Xi3xiJ7sN
4faPErHkBRnJhmfDkrY5WZ9F/hzFuVZsUtd0KrjlWITPf017M/3vQo/VLbP8
LVIBOeJTuMzX7C2lbYnlje5LXS36tWlngk6EoGt3QgNwdh+JVzVs9RsBdAKr
oUHEFNxixi8y6lWTpJEfzWNigykuIBcUG95RjQdBqMEIp1jkkYJhxCfgJkHz
oavqciJf6WvPE5b77UTOzZ8dfSu3mJKaqS9+TjRPC8D69h6MH7uma3f250uT
XetcXdhpfZ7vYt7lbZrrhfg7IeAxO07bnr608PWhRuDA8/Q1pd+t8cHtFkrI
6uh9vvoblJxo3WczPJXH91PQ0YvOk8hrv9y4n6Kn+o3I8K9l89DYym//jzzl
m1DicSchXdPD+ZqhUzfnpV84mSJz5b8gXbUQzNAk1bXeO+/zaRu8FHJD4eGq
Oq75U8B5J6CffcUIXr8sn6SvjRU9GX3BY0fMEg58F2GBu/WJvfdVSYVXFJZV
/mhJLlYaBpsDweBADrbYoqtNUiudgd6vGtOMFUXWWaikSj/Rv7Uc8ubPFD+w
9QVXDGzqgiHHXZtJP2H5/Cjzz6F5OlT43Qoz6BdChwj3kpUNLO6O8bAzaZft
TM+axM8Va06mGeAqwEsxpB0IkFzzm59YHeMWPr3FKUKtK2xvcfBe4Ix1cHCn
4o6k7T5+T1+66ZC2bSFYlFlGNKv5ntmHuJsc4CLXmfP7UvuBr0FunMqoFd2D
9oHEeblHuo4CjEPmuG0GvpcyoT4DS5v3uLcy99G2bEYU1VCSA1jgFnDf8IRh
56S/MaAjtyj5olMzW60pXLp/1+oTpYhxiY8eDQUAbSCei4WQLZM0CroFsG3e
HM3HmQrtrzEDhZaMbhJMYFqrGonjMmU+FN/i6XR57x+PmFczvTG5f/cJCPvP
3yYhG08IlaQoEcLnwNKgpXDLtd+51PGRSrNqmPmP//COxU1joydUTIdJH7HU
0hiiZl/nVL1RB6AM4qX5G/J4Qvi9ocUbBStwV6KDgxhpYoBlyFoV6DMMMQJz
mYZy+xy+k3ukhKhsTnnAXxf6h/dBMPD1QcQVirERqHgoGu/9ztD8wKOhDdo8
xm9fDaNhHdmCrAEz4AvNcnm+nbRPnsVmaO4jeN7HusPIPCZFRY0Y1qDEsZhP
jyvonGhWdxJPZQ9CKGdAjwGW86vwOn3u2Q3jxbO3458PiKMTTk/6GXNQo9r/
1dHd7KviPCWKymO7NhziEhEo9TJIhAoo2XbwoOsbogG52OxxUxSmIFHHIHTa
oXf2l+RyjbDMQcmIadTgO0LWUqr++8Wtlo1SJMUsTOyV2JYkzx9L9bF3opuO
YQMrcyrTQBCBsj8F8ylQ6vyR/SW3Qz2vvCx8Hwx9U/nrcyh4A5vRDFEcBxNr
0qjd98nNzgs7M3t5nmPnxSMb8dF/bXuS4zMYkfZXpYD4cJO7G5eZ5gSPh4n4
4mN4EZw9J1vbmWrCUULpmeL/vXAUUhvcT5c4EeebyARMtA25DtwoYaIGgsAo
3QKby3AVxsOGRYMAtNmHV0NMLjAha75iajrXwL6C9QkPz+1XVN2Splv4vCPd
dMDZu4uHmqAvsVct/zwHQYIVh4JgxgLwJlEs8z7SMzgZB9PX0ZWdk4jddOzV
pZ9e6WfUWFgb4ep2YtoijzETzSdrPOvqsYrRp12NOURYF9Pp4JQUJTrCVgun
sVu0OpeQSlFV7liqiXXsyKv2MR08azdqxfpLYhmpQkRj9KhkhX2hoAiLeV+q
zqQGFGyjz5wzgZLaH4p9n9pATPmY3QJOCoxtUJGKl8iH5QBN5JwK7eZ/3XxY
/a0TB0JBYrQ64ZW47BOOrB+4kg9lj1lqFwS88zrX8dSSIK6qG3PT/aExHBni
XSl8U7TBxFCBhVr6xwFOwZtTbvFQAANOM+9xmxAoskiJ1ygF4KglwaZP9g4t
a+5p8vpdi43jxSv6FgNryg5UcaCM6IM4nyhoc+uS9FoEWltTmSDKQDUttd3m
9nw16B3uvvJcxkVs0OhUr6znK6lfUtHDow4LnBPuPqW9Q4LLBGCYqJjANCIY
M51Sa91POUulXEoNXcrM2ogElQW0//EygyjoMKWiUEHjBJ1BqCpMa8lIlqU1
hx1S1qpfARGQQjaWbJDgPn7B9kkQyZr7iT1DcvnN9k79MZO0/CznYbFBqjV2
nKgWDwUVZVW8tqtvcU3n3NHJESZxsNfQHO9larmxk5AXlUxNb/6zb1dCDq7a
JtpehRXy9DIFDr5KfV2eu4yUEE/Nwh9C/NRqd/biyHCdB2I6eZjQBc5voSev
3uqlHG98GxUSzjj1wnnb39+HSDSUs7bKRVrNKLXaeqFDebW1jelcN4XFW9M/
9QYkg9ktkmUmVT4iQ3ZmlRT0t9TrcDF2+k7hzw0bepdEAfmS6pSI98Pwchy/
zmAtf3+aE70E5Sz7wDPVAGLUb5dJScerLHsKvCy+4v31OErpTMkdr/PILK7N
KzGx9VDBbATjRl8CDQUFQs+UVyAumN1m9d8wz2ykNPu7pToFGHWbC3WQzZIx
b4aAxMVETi7eT6MAX5NtLswhCwBmgxb2FQ9oY66MydPPrgdkWZH4QFZ2SSVr
MUeIxlKqRfSIMYX9Gbo58KuIAwdcQBEOI38kVLswV49mvuM73kJw2OCK3FEx
DVNvZN4dtmsLUi3NWrpV4cYMIpi7TOj9kzYAVHNljkWfTaPhFMEMrKtHqv2L
JVH8rgKvBUbzgZQGGhO93zsZketxOiGicP2tXRh8GvVk6GAMm2VzF48+JjIb
oK/b9AqniiaTPqW6dRRC/GRKq+xy02riJQa+X07V48q159GtQQxx0WzXPKnX
4381WjsSEa8x1ogyrS32vU91tdBcXf7alX7t8rmu6FAgYGKbV8qunuPLUD53
WUlc3364patI/nXZc7AXbJsnRAsw5Z1czRMnZvfPBiM2cNnilni7KGLNK9go
vSzA7+XHOq/VCHyRvKOSHszjuFahwa5M02ZSk6Yr3ROzFtVNWL/TqzCY/n8U
GdnEHmviqhexhxQ7URvQLB6RjfOOXcuom6yytiVxAU4xpX7MS/0fm2yv4R8Q
4My0j0IyY3Oei+7IU16x1no/LDBD3gWHcoPl/yLzoH8KQUJgPtxTTM5hcUgm
rop6xyAsJcv0tcTAoMLZphYb/hRilgfdy5Mdrx/jURkOOhRThWw2LSeCSa+M
N2wSkJu1oVRPd34fPEWmezqvY/m+kWvcnyn2321VImWH52/aBV1sGkCmcuQm
5vIZK5/uE+OoLZo7n6zo7KwD8QwbnK94IcUur70aXbY1iZvwOagKy4jIlxXX
MLV7DB0+zZHksW+7rnxAfTyWAdbZ8XyPIJRCWEb4dqt1mVATlkIY4dytAVhB
Iw1SRHp5atTG8dlQPqFtUOeCEFTDukEPV8TSvJBfuZC1KXdLVECisnWrd33e
3QfGQg6vAAMEnVuWWZqY3p7+XgaKT2bV7cLg3OL3BjO2AU6439PSI/4Ck+gS
hcIyLgmrKWOmboGubwg/t5ofFp4NUEcXwyUGhJNhUxh3U5ZCN9qtsjtBDxhr
vHVUOjTL4vFz/xBsbZp4yT5Hpni3oWyRv/U3Nq/CZszRu8W/PC14zfoM5lBS
tyw38MyfKhWKJJ+zxWUrn/BkSQut5X4rdTaBf3ny9kVNPqGWknSrq1+NB152
EQVtplGY2XrvvEqgtsGJf3lO9MBoKB6H/EiseiQvwbF0pP1D7G7ICWDrznK0
DUkuwTz+FB4jGl4lhHwbbmktcwHbEptsnotpfXFKQu4EuerCZpQb6uVOZlGw
onX29vb9/GVbEdDax5iN7JkjvRFaP5HDS494UJp7M3N0PbbihHP7PW9x/B2q
MbXzTxVwgtQf0fQgNxB+PGN0Qkm1HUGF3hRpoku/gx8Hupzm1at6BnO4sf/J
h8NAvzismsUe17J1zhZcwarkJvTD1lLRDa/E0hTaidmFgi1jjDjTGmdvKHQR
hSiEIF/+myzi6u6dCvMs4JsXC4sWtJX8l4P5tTJAPU8Y+euUO6LbCBIuwjPM
XoCpIISV7Q2R/JiwpTUHNeIRqoqUAr6fcKGLQGTfHNDAxjxvMBeJ9kPcdkDw
1OpwmfWBuVlhPlsoC5q2eMXmFLw5nxgbcWyRAIfHvWlu08gZge0P0ZtbQ1IX
d1ETs/I27nz3Oxu8lrfRAtO1U2zBvcfrvH9lowzu1Iix+CYCh7UJBZXUWn3a
MlJ7FGADqNLcWim8aO/o2GwAz+MDOWRAcpusW2Id5URdmKZ6A9retaysoCfF
6e4aZkn1tWYl5snnk2AF231l9u8EWt1l/SvVRcKhu3uXVXAJ6LQ8iLK31tV+
MFuN2GMflVchk6XtjuE+NGMTYeK65Ip2UaGPbOo5V31Xnn9n89k/z0ow7QoO
k4vjPB4jMIRyxX9GJaDMb+nT8igtq9uXdR7ocz0tQoxy8xjv8Rqj9DYCczPS
swFpAhqYSPiSVmhS58RJOzHCSUL5tXfq3LujZR3NQIDN+fSEK+sYBzdUEMpU
b/P4A+gNMO1eKqk5Lxk8VkXqpOhs2FMD/jN/axl0UxNvtOq4/aNIHQpKfPN9
KDkaAnxhKz3JNlxro4S3+pCL1WsCt41uSK6YgHklv1qFlswcf01PL/ateT3Q
DvgRrgoQ4LsKd9swfUlG9ntLS5dVwtkPxprvQ5Rdn2PmLe+Jnt9drh5uCdpk
Mf1qyX0lXOijAkz7dzJoen4mbrrZZTUXID/Ur0Ynl1MrcDKmMQnwOuKc+xuS
1BwhhPWBc1n4rNfZU6JtJD+ao/oLPza+rSEgP2nTy5H66ClEhZlhbfJgi30b
LvLWGwHni8QTuayD6tBA5fkM3eBr66kfOxL3tVDbbuUFRMMOKo7VO1uTb8jE
aw4evGCL7pHOW5rBKCPIAtxzfJcHlaqWZ0mYIz6jM9kb2GEgXytVFaUiqxAk
tTYLVtoyeDNKsFNjrYiFiJR9C2jyL1AC4OIbGuBCH3VHREjM7ikBYWJrL2xx
lP/2A1QqTi2Ov/enD+ApRlUNBk4fyNvhbBpN1y5ArKEM0FL0d91NQnbDtFa3
Uu/hWFLH/ruusyNOdj5ON+rcVRWkJfpCk+1KY6LRdOYueOd0YKrDhJS2wGll
KKCdz5KNk8OOeU2Bf2fC/ceZ9RisYWol5EHNL1xInQkYc+eUEC2yifD4sMze
9zcYKMbZTvpj9jjfXF/8rMCDLmAdD4udCiO0HI+R6pf/nA1KNXS/v5jSq2tw
xRRPBZxU2klM1ycaT0LXapvoaKWNqBZAx24FwAignjdJQbt4N3nHqeDa3ZQ+
fcIIxuebiibOgLwvtxIt2k5lPcE7Kf3cOBHxs4oRr2At6JIfKj9co6Mohfqi
nPfFWnbSRTZgKOJHY+QKmN9BkFOtO6J+OJANYNWIasLqD6sDHh2WOkIiKGAr
7DZ5rYiDvoRl14z8y9EEHlRZr3WUkw7HWH04VX/jVfLmy4cONMQDdedI/VBD
pIYXqLLRTnYecp3HxUtc5NmasvkBn4V0KnXxoOcqPSLabT1LC/+kBrOwaAHB
lMDkqGCoA5A3IZK+bz3Gbhz+3wY98FRzo8ikc75v5OHmbvXKPSV1DiOxoeuw
uKiH3Jb5gkJf4BnsNbuZcADqy4qIt5gc5zMPIV5kLIC8c9IjXrmcS4uw/zUB
aJI/5NE1lBSO2xxllu9Gt13KYAO0eonpycrTygshXni3+7RpxM5cBYolx0bg
mrEI0kqmBZ7qRf1BoqtZENJkXzYNOXd7gaxk9zJPy6YvRtxFq49UNpKS7oCz
5WvOQX7waUk++v4pFYTJXHa7i06uY82pJ4A0GiV5zVotROAxrGgHlUBJeu6E
cuz8m4kXVST6THKUTTqnOUrr8SFOb5mQTWUK3LEhX87XglN3lE+dWPDqu4KV
frh6yl0DntzhLeasn5jcXNKYRhX6E4L8e8YAWaKYOj4IVSAr01v4Drs+rm5+
G09+clBAdmR7Hs5eSr9tERu6rAsk/DdaJebxDC8tS8BPhU1FuwpyKpGmWazj
DlR2I9PXv8DdD46tMQnrIU49woj1WYJHXDOaIYa/32EMCzDtYGkb945nf24T
GoviSp4pOfFZtvszjKFzhfHrEm9qWtfTpqMaKav4Vh4MX184vLctsORlyQlt
nSMfqTczp8zJ3bJ/9Uno+6A1qcPPzsIvrcV7iHPNe8POr2ZDG7IB23f3oj0d
MdWz+3At21MoFeg2CkUJNnjXlAqiksNx2LZ2TtwuclYb3RL5ugLFLGw2eEEd
AZ394eTn9iO8QDaa3DzMwj0LOQ9Q0J7GSjvj4pgKFpgoQiHCXlIbVN4w5Ah+
qxWKqp7kU0iqvCHfdg/llcCcTX+NGELF9sqVEv+dFZSgWGMNtLaS+ECLr0dO
q835S/j/crWQ/zTVUfOJfwZin1uYQFe40V89EnNrirwklQVNsf9nG/IUrvud
CbQ89OnTL9JOz9qiP1Jhmu3amaizQSnO9xLZXY+kwe3MuoPEdVALCwMOEdRU
hHdjN52Ceb93HJ2PzBUtDyh9yAdMyy2Ytc67g+QvCsI0f76uUlhTZbXOPbvY
aNXV9ZFwrwoai+jx4uYnEqA/0GWc50WsmDV2UjYQrVc4F4yZsOLNqXEA011Y
NjmFI4kwftO3zdQfE3y29HS6JEUICsMjzfbLRMXHHjvKUSUWSC1+amcaOgT4
b2pGYZtP7CMImNDN/l9E0E4d1n/ze0pJ0/2ASRR1J0ZIxvJm0rw/tzcARQU7
RL3BUXExwcbfR/o0B2oyRWGJPFkDgv8Vz92bBlKTKEw78LA+lEvzgdEhXnGj
YBG3A2oyCAqLGaUtJZJxHQ9l5XR9roGIsVm2VUKJY3/aHMCMDop6zZl4rhGk
S7pmCeR0Vjzh5zloLLsVSnBMabWaY6D+s5v/60Vq9uluk7Dp0kD8DuyGW7ud
IHC3//l0tGc04WvZKKDOvt+yMVO6O/5BOB9HEyTEPFujG9HenK1LeAwyKbaf
WR0hZp9r10dhSFgpAvsorBmqwhNaNR+CkfIDdDqMOnRHQlxUUaajnabtB9sW
W8ISAEzD+N+6MtnvLJvy6CGPlz0Ws4Gx9sLNsMpQV5v9Y76TwvCIOZ3jarLa
zuWJXKuOyqipn2BtiyOuUh97kVg54un0Ud3DA8uA3WDzrty4wKYoAap69gCm
bImHnin1QOVHbnyYnVpTBKvxnlk7U4+HR9b/+xaFb/npgzsUp4+pAqp0slhz
oZ6YBLlXuNffpI2lWT9ZsC1gx2sEr8xAehB4zqqnDdCCequ7tkGCqmue0cRz
pvJbPqMMz5QG7ihZaZbTehKlit3cYXYmWpmRhyz6GYtBFvGTDJWmy4k42kRO
xetrIOoOrod2JhKYSpYE/n93974ui/jJ+0tqaw4p59ti3GV7H7sAN3h4GCru
mF7hPvJ819WnOmXNJ+AsbIkvdYOi67bZEYFDxVTv12X+gJokU3wgPveK4ETu
zWQZo6c1aCiC43BQDLEMtJSlYE9a/uQPTb9vI99w2qQb38fBg7NV0g+/iBw5
L/Is83UuGisvZzsfdh8BWUIFSudIonN1ppYpCPMyCGCJSEmXDGmGQefnJaqx
OSJjsiscv/ozhEST1Vm4j84RX6BqWJn4ABJN3o5GoXJ7Yx8TDvWzXu9fXMQw
j7ZK6By8jf2Cp6MzWPOWtiIPH1J33yOHppVsIWwhr4s/BD4Xcj0FMXAxKkuF
adCafd39RScSE62M0jynmi9xiqQOeRRONFzY+HSiYYwge9zxcjY4j77YjQFR
N4jMg4OIedq9yZGMvUToSCRe6VxP2Ane16wJ9e8ultb3aif8Wx9rvB2vO4on
heXKzRR3OpE7XfXEdOEz+Jhu33tVLKVtHAUSBPrkkj5b5bdREEcgzT4Ev4CM
g58OUDmKUbz/F/lUfG3KOIORqGhGX6jIAT+POtdRxf12Gwx3srspmnK7Pl2+
CPlw+FTJ7IJe0UppAgcdpyM1FYbXnssrg5TyF/3cMB4mzgjYFaxZ4BjSlh4t
LCjl/6hoNbuqfPgwRrexgcDwClDsF/DkDFSskyKYFHcMiWQJeuj+ajctRHbr
iI8gAfWdJEBsBvg2HOkBbPKvvb8iClGKJC3O4A5ojajyvE9BVfc7CoENPBjo
jHTXuX8TePLkDwXk0kqj6cSrFvOOG2RvOjttGSsnzwvST4iD+dTToa+w9+0g
Sq8xSVBgPhKeysLrWRg0nzk2j2aayXBFvEogo6RvTq5aNY0ZOuSz+Nd6PdhL
JBPoGVuNyNMT71IQ2tX/426SwOQNgFlnPpSzkwCEXeGKTfdigEq8CudVluFx
6TJvkL45epgAMZjBzA9q4a+Z18n/9pWp/CrTVjdr9Z9NY9sNDKv9aPD8IyOi
5VXvyRbyHnTuGTdU07ZeKnxjk/LyLwmLzKwhtoeqxJnVTnvzUlirkoTE8PZO
vlFKHXBCLwGd6P7GQ6CaRoK4Q/3ioVLu3n8rl2JwFXudc4Prf0jrCjy/vuXM
bNhe+XsHdwmAv79r2DzZKlrVelKkHIZpkmAbMCTyf5HeRgtTD/tRMbfBmbF2
sDtL+9/Jfbfv5nukKeuGeVW1cZKIogVoKqx1dACDsfJXq7GYqMt0ZevMtWV2
Z9pAV8bJTWSq3K+FZXtbkYLqEd3M17v/G1lFSjTxeDOxDQyi5+k2spXUZPeI
n+p4+08cMSdGJGJqQOTzbOK7ZwmoY3UDoLnBXkTD0aGj4U3clFUFQKuXshC6
xuxlD4AEcZgB6LjUjuUFHc/XlN4hk+MdPMAiZbK7FZcceJq5c49T/pQxz4FL
fc9ZAD+ndAB0H7m70mTnjJqSMIgUs7sqbBbSnFLeAUVfDrQYL70v2BMskvAT
DKEhe6rmsJ6QyHQoCSDPshJnSC08uISzKGvUZNrPxj0ukQC6iyeB1SD5jTM1
OkhvECG3qTU6NmfZGZtpRwDKjrWFTXzniSrDidDatltQ7Oe1J8G7Djh4uw33
Z3HvJLp2okLLs3mNNAwZGOEGW+Nu87BMViyzip2jL6XUqA/ij2C8QjOjDASd
NHKWutACNdHO6UdWoHwEZsTDIU5/VeyNf6wAQHgsnrFKsCLrhoFKKrYQNuzH
u4PVPFwCxMhskziJLuCVfEqUxWyZeNSCs2jNxYwe6aC0KkbGrsBEru+DzXKg
UwPFC9QM7Mq84N4WeDMo6WgeoQHAEoFyHSrMP6TVFNDQmkS19r31GAYWM9M3
dWtTXo7Ta33VYTFAYGprQnWyPonu/JhiPvDdODu52k/zB11OYbNo4RY+fNpF
QqMn1SU35P8yaKBsjs62xQXE5SSu6+zrBTGO8ZRH4VqY9i0l4wJPFOQRsukU
ZlkHaDrI5mRWwri2/uHoCTlsClwTt43Y5pXiiPi2eo8QoyL/egiPVGv+lwNp
YK8pifKQSSTfiMrkYNWLPy8MC6CkYacBLZYGEuMcfjQ+jqYRbMOnC/o4xKUw
zESUtuTf9mU2nUfuD8X7YaUmgW13wlzB4S7CvxjWFiiEwlXDthPUQPtcD86b
5XNFit98XxPwneDe45UMdw78dwt/ILtyGEUnubnCVFrDfur7kpIUZvW/xRJf
CW5BNcvSHDfiRKOlRLaXkI100uOhtrLLKmmRUiauh6ENIho8ebolN1RFwDEd
vzjH8mZprzZLF/lcZpzOadtNVs+cDwxDwxj3am4xqmmF9m/8oMH9heqGtPf1
zl/EeE6Or1dHX8YT+YCIjvp3bt4eBek/Ndj+MevYeIjI+P4hYX56RfEYKGWs
qYA/wG9ZI/12h9sU7PD5eUpfTzRTcqPu60cK6cftjxjNj3mA2bGMAXg3ESzV
/dZM8Zc4kJfbtN/GOryLHHiqsPfL4p8eQ8G2KvjEFqxYbYMFTK7w+OjeEMmK
vuVoPz5gLekBKismdU/ZHqSPMUQ39lLhAJMJ+GKt+5qXrnJ8xG2j4l9R5/PD
apAjI3Ff26uERSlJ/3P7QGHk3cXqwrwlmzgGRp8z5BvY6BdfaMfPvj3r7vu1
MEwWklRZ5Zz8t0cKLKVrlOPcRDfO58JFr1BzWQzr5Lxt1Y+kJPFhbhJ+ApaJ
+nKVesh4cCZjlrHKF9ZWVIowDiNfnNDsGOO4eDFXHhWi5uhLheqT8Z1guW/8
tJtKfqoOre+f3Fwvs7kmA3/xznEBgxg2QTQOAd7pi0k5HFNTRiIul1RMi258
6EGRHDkVnSTbZc7tcXZNu02SkPTPo5wGQu5V6QcgaDqwmO/rJRblgOWIgPYw
iweBjy9ZOOHQ/T3VndcL6Uxe95FSuXkTlYREdZRON9uuEU+G3tkRNXWuKzud
+lZNivs+cEHIC22Mg6rga2qX3bsPDD0530avKME63HS0lvi5od2GpIBrD0p4
1D5uhhydKJZWgtW+vxIQjU+2Z+SweUfcjHhUcE4571Ptn7LRrvXvTkx1d8M9
SIVlvQxEeLPXSaLFEaMS5Hz+HjW4UPenFZWkegMrhZ1dELnu9J4cXdpKfU85
LrHztMZUbtDNreEMvDk6iS16YIjdhf4CEvMcO4/AOTIxpiZju47OOkSLLTQD
+lTqTGdi5Cc6d71aTFQnFBd78c6NthirFlutdNHApysldKtVtM6gwGFBpP6+
aFeDloeuHuo83OWB6FPtbS7pTye8kZxtJxx9AHxf4pOTjDpYf/TQ8pWxsNNG
W44MTW7kHOCVYEHT77CrErNWgWlNlMUO1Gbv6oXMHgtw1gPZ4VklEuMk50PD
1Y4UGRv7DicJhZYxrqJHeUIDY2iMfCCeJRNZK1uLo6ZRIpFTpGL2SQmZsuhi
1rTMLCbzWJ/zUCRs++Sh+NkUBwxxOWNbbkByYEqFqVjoEjMBgujuJGy5VUKw
n2fZtA5wGTKGvYYei6GEPT7TiU/+MPLYEosA+v0pfW3g2ZlC5Xmu6VKwKtbX
WavDFxwwifJPNEjfwht2zZkVMqnJAh1vUxezNWLkAxoZUz9aN3erwoWrQxWR
MnDLEo5lPNvfzdXXBhbyT9S2JTLiecCsGRBGpMUGsbQd44pkIcbnCS+GlTT6
OWm4Cy9GzdQV88VQQIwYeodVQatNIwPC6j6qhn7m0bgYSAHsSmRfxj4NGx3H
FMPG/8bPNDGTGM0L/6caSXaT+EyG/fHhzVCru6L0CsdqZz0QpC6c0onQTN84
JcSTSiRLg7+HARShTkeJPyh7093xHrL7isqIHmLhfYx0O+3BVfYtL+2DMPoB
HT4AUw4tCl4DrGl0rBL1/lTtVntzDY2OJfXZxnCvz3HsFiZgYKl1e844RkDc
HUUMc/ghMDw7PaJoi55T1FJ1DGGSYTKbv9z36kbM+BsfuKg3B1b++4LjwG7g
g9zeldhutomavYhbPpdtxKiptybyWZVkZ8FbvfJx+NmI3DK3RW44/yxTBXaK
P37argb46SUAcbMnO1oBG/Ltc0FODrToI+J0OgLkaNkYc3/GmGeRKm5vE0Zr
akgoZ3GaMH8DHJ9C0f0ZV0lsUh/EKB7F1ZvRbnhA8ZpbTLQ9SYzlD0ixhnao
dOiZEDm+4awCEy2BBb6WjvLAhtD2VXU+RqvXKbdaOBxI+n/dTVMhT4os764j
avwDEfMifUtas9et0WYS15LAK/uXEooCv+4jlJtRaKel5C9y8fkH+pCGHCKF
Cx2A3eme6GFrYR1IJYwTPe1SOS/vCcVJ2PlWvFisbnZNwh9SjWa/tgPm/caK
i/h4i0Z3txhAURj+plA9GhjmocIqEZ66vjlSkqtLLI3msYC3qR+8lTk8hAQc
XJm6Krvv0gNHN7zB6wH5ZPaNiCXCh3nPAjzS50jqby3nj8OAifvLC1rvTh8k
VKwVyGfiRjYe7tYZ6IiqEdn5HDJZxa1LEXKAVAnx23Y4nWpHXSBf/rfEg7d5
u9GlCzBiFD4LkBsY8qddJPabV9/JANvcjjeRdD0bke19NjUOsjJC7hNvfjfY
62mw17QojIBJH4eqpiwKVp6La/tHpIfw4u31QWiZG95bRgAyGp35bnT3xUap
I4F573qaRyL6U9VkAS23nv9WINqS5AUx/2RqIqzmYQx4PGZTcmsOFj9hDyBr
ScLdbI53OVYzHK3ZsVzFc+qDHfpwozEyweA6JRZ53GMTXfuEF6m4SbxylIJ7
a135U78xoNyO/XG+3RnHqO99FUbD5iwAHHwiV4bpCYBN1U3Z7XCGRZQUSmnJ
gxe16LRMNy8fPKLzi5y0H5ZnOfId5WuxB6QQhRtzYrqoh3L2E0PWW+0J1+Cd
uMQoFEMLB5oMWiGDm5HePHZp8fhXLfEwmBqLc6OBwQ3RFWha27BWdLxTk4PF
DoTpfNkHz78UOosyVbTnxrVdWFMIyL/d3tBHWAdhcbrIHM7yIg0p9zPQfN9m
izRmK9MRFNHIVw59HzJB93FExEuBuuxk4gd67Zz+bGeenSGQzx3Kx0RhRbXM
QT2CHsD4AW6l0fGxl8Hae82nCPT70wUaE0LhJjBTgBNQUKkcPipGmCECk518
W6WpeUMXXIC1SVxi9evPa6D2JALk/Wfp1/Lcw6bMJbz6i4+HhH/AE+GpNVXq
QqBDAIMSC8W7/K1tCvP7ErXQ67AcgApf/UC3ay+NEy0Y7QTUTCpik9NY/R7H
CGWjMvNVFogXWlSivmF6jaZ1ps01czYHE+nL53YVn0FXO02gEgcGIWZld/gr
5Y2OeiHZfiJRaAe7ony5SgaK1EsxNwZqnMSBGbwni1ZeQRIsuMEUGnpx4zdP
IqH5BPjePnHViwGhgGThYo1VxgF7m1eNdamZrQovI1F6oIIQUydEuB5sKQXn
knTrsHx+f8EgXaesNHbRCjaj+tQsm9RfthxvrBc50GmX7Vixn2VTBM3L0oHB
PUjG8AHn3JiJGLfThwThgyzetKUH6TITJv/J6mxahbTqc6gyFg0ov6ddzfup
iQdSjZENBMAcTh/PYeJys8SRmQEwSnNmEn59KHnx44GYBApgoU+pJ83650BW
pwkfxAOO4rA6OAQ5rdKSGkgIgHpw06n0QVP9UZJs8NSOdy1U7Uqrkxo8VK18
CA7sMEm3rzYZjj1/TlPh6KNrfmiHg17rYyMPgfN//agY9ZQH22fX90ZTkcdz
J9qyQODVddfVfb55OOtsWKtP7U5/VXijFCFOXzp6gMo4jGzBXOJwPXqFPv0t
e6ZzjLtT6Ra+AH0EseRoNC27kzvcANLncH6WSqsbNUilGQ6ZnxsMpRz12z0y
wtZ2d2rhwjOoUPwMaoAuYxtMYkbM0qpwlYbARllgEaJ/baCqfW/bpBr6/azu
adaRIPwHKvMGJYemMml1u2czEDYE+7SWQDvPozGXeOdlVvwsfd+L5RKM9FOe
39t4Zg+P0a2cKCS3RzogbxLmpY4dr0pL+q+sd4qhNIgL6OxkzRP1rrFcXTlV
4QSwiLN6RrR9149H2TdrTdzEWP3eBGuFj0KvccF7jhODaE3ioyI0w4Cztks7
IHEy1zUkCia+GLsS/otDmm/LSgBJ+eFc3CDVKUqZMhZM2GOuJnt9mUwSuG+X
ZneelGG70ZRiqesR2ufxyR6VjTO54MdW6L/H3cmvzCFlCe2PO+81lDihwzDu
nQjq9+gThzae6v4ppg8fuWfoPXdpjBoXh63gD0TWnNn1pFaBdtz4T6ZOozA/
DdAo65aGlVRow8qQS6qFFXl80Xn00rRcJvJgYcyAmAveXFATgK+7/UL2a03x
1oJv5GN7dx1E288O51zKhZ2TvlExNMggeeY5qRyb3vrkuaRCEe6uGk7B7V8U
DY3xrVOxtxr5Y5kJ5D2HQGuwtQoyfm8SsobifY85W+S5I1QVS0/5OoDwKD8E
krEQEUZYaXKe9tpBYZ5WI7z+8XXmX2W+T5kV2KNcOo4F0WD8nyaBIOBfqAGc
g/BPP8l9RuHJMaeuUugD24zAToXIYOtFAaorUL7B/uXEqf7SMWE5ioxiUl/x
+hFoKmSy2W4qt339noEoCfDZpjbAhG/D8Vphrv+T4RQtHRRp+YZZo+VDbw3s
8gqX5LxZH8n30CFFsXuZ9mJQ3oDjahjfKn453/GeOwt7kE9eFO/MMe4UqfMJ
U0lazl4PTyPLqijjpS4LVL+MAO/dMSFVSOJHa7j7SKtYuVcxkIlDV4/ZAC0n
eHCsKTPX+yQQ9l453f6uPs7G7gVGdCuYDGUxdLVkwA3c/onW+xOxNCGNIxeR
BSnClnWwahFrM7YEo/DYa9IdORj5SWXzVeFCU0aF03sg19TuJ8BKsAUvfvyc
kRLxSU5rwa6aiIikNCepxWMsG5cgRH1xa7qXZQjDW8dA3iszHouLwHOm3ymq
YUG7AMlCTXgJgCz8n39VfTTCLk4cW4vDPVJ/GPkFAmnzUR9W20gKHHVuYYkD
UpSCnc/xyFrHrEh4v0rUC4sQiFu7jUvTtJ3hwJWu0Al47LW6rNuhFMM0MO/D
CX3YB4Tv0K9CjIi0aO6F4jXnF7y6S/6yBe1IECwIZGNcuSfxKpI0c6mm3PYG
dtJjsFuxi4EwwrSMJCSRDSwHvPEKHOOeJFE1o31YTjzT6aZQ3RWlpN40n5hi
bnK4NlD+0aVTQ8jd/E1iqQmEbkRAJEETVvCm4UCih5AmZPrKY+IMD78oOG2Y
5bPRoMm+FiYrPRfRs7cv7AQ/Nji/ACPpODQ62gYwkWKkD+Y0AIp3DRfjDL4u
WW6hNYc1MJIgLM0x0kQSwj+n/sQVZCeji8lS7o9LId42TMgnNPuiewhkYBSq
URkfWqBZjfAvsa2+xxdtwX3k1rgDC/MWVaobOCBQ7olAc4EKCyw/09U5wVKL
MS8rt1g8qYJEnMsy8zxrcDeyOkWvFjlGedTgoKdWtmicLV2RdXYctPXv/npp
FRJOz6mVL4jH7rtiAzJOCqooSCUOwpbG6x7yacJtGBjzJWDtLP+siJJlSvEt
rxGFJpt5RBhrNNeekYciqSXCIN/83ycSAHONjxSATmXNcLeSRWGaXUur8p8T
S8K64VsLDPY9MREAC+/9kXrdPy/sbEhEyiyHsE3S35dC/gAd/bbgwyTtpu/m
ggpkzJMS+2XzqcgGYw9sxth91t/Fyps6DQuvj6pFNStqmhlDDj97zCGCb8xB
Lapgm4f9+/ZYwoPNAq+6N0mQ1q3r1au+wC4Ht8PSHIII1ZWKK/rDk9Npvtss
+Snc8IbrFO4Rs5qkUL9SgXXI7h1Gr3jMbSaNL10Vr1+uiqMHGU33+8nS3+xq
HaRsDgHRPERI5fdLtGhq5m6XWAlzDUgTjoeB+USUiY1bYCzsjwvc6p190uri
BBeJrMH/47fToiVCoJxzYeTmFOFD4eYAQe2eS45Ws/JI2hTpt0I6XTbTMZGA
OUDsM635hfJLxqt11hNWP6Q9F5P+Np6XKAeIbjlYuKadbJ1EEzLUszISEraX
Vh23u6gj4fJSYwNHbXDjJjFLUlgoQZ7vnSvge8Id/no1oA99qa9XHu/cQsqI
/CMm5RVTRv2vF+1BcAjsYOH1S5S1nAfMG/a6DvnwVzEQy1I++rCqzeVjVW4e
FtWuSRrJoQWTTZ7zpLzbEMSkKr65PWQ6lvcTm6N3vW+jblxkKGzyGO4sauHJ
mr6ehiuugLKR8+pIvzxuyCHYu18Nz8G0F744cnCcU64QadMMZ3+O+h7lhAaO
s3bmB/GJDhISYr7w1Zc/7zP9dI54Mb9HtWYy1UAUCqGCzq9YDNNDSPrt/uhK
AVPRmvn3ndIM54cThpBNoX/q6srUA50Tcr2XLdJv3AEhJ81BxH42hSksrY/P
pnxk7U5UWbreRKWvHC6Q+xjQdbFcJIKWTzguOx4icGsrhUDxoda/GQqi0IWF
39ab+aUV2usAipTVGQtsUFZBu15OKVA4ANGdHuQM+uZKZaLSze5737lXBcYT
Eb0xsBD0One+6FyTrONzxo8O6+uj+j3DqtQxUr7xEIWfQAG+AhwjmhdOmY5u
D0f59o8K0/2Ek6wBsQJGNiiSFVu2EvuLb1seMub5blSkyabv3K9vEVEt+ctk
2K6Rf6KLgPiU2cSpOvSYic7K4pIedmltR1rWlGhn91QmypnZGcdTCTFvL7SL
RLV0WB/22Z4cozHR2ev2tFbfxNOiNZt9JUZ3P7aw+oyFG/mKU8cwGA2WNhth
anF06HjZt0KdCDIFkkaV6mGEc3zW2CgoZvf6vQnR42s2xkNkm2Y8+IRoT51x
hCQxSskZ53E2uWJ5zy/BN8fY2T4fzSklHdxr6GgbosfiwdUJUqhIha+mYmle
OHNiBSelWcWAJ+zoKUHD2b0YZ0eLPWnO4zHecpyMkDXWFCZQmLiGDHtBn4N1
GdMSUWI3At9Rk0TqIzB4JCxziiKa2vXjsGRJyX+sK3bw2OzepMNz05yXxiIP
4qYfB+9OHu+HCZlgoJrowo3QXwKwVm0WvMXSBi+6Nhd9pdfe96frA+P4qfW7
7y58OkHll+E/pZl4wSCE3/u3F9tgF/42gMg1UQxULfekCuxnNDmpYAdYgblg
mWWfWOXYqHAFr1EVNYEmRZuD8C/Q3bAN894c9UJ0jyFepm8cCEkl7Cejxdlk
4/mN+e/TxxuXKcfwLklsOSttXqxZeHYrhcWFOCJ0wGgEPscbD1s7ZRax3DSM
sWSndyUUty095DeLzjlyWi0RAazdCCTWUkxAlxBK3wyr+d0d6jA31zMYcV3V
w7Z9AVkVpHcQWrIcwQEN8tawb5iYRraue4wj3aIiyf6quSrBcNLKZKfT4obr
e3A5Pu1QJojRR17E+IDY4JG6ZP641s2cjXoPV3JHozXHV6/UCSBkqotjiqIr
YRsFI/qt5qU/iNSMHv/5JzkbQEfUkSyIXhQbqCENOHKrsR9HmdUW4UGMLMZg
oAHW2UHnpeie8i66wd+GaEUHH5/APuD9+i3gaUgVrQA+olIckUImUTGFGkeI
nLKcuEJ6bn3H4XlkQRWHKkDqS/fNTrMSWUvCEseM8n9l1xdgRil57VnoqlAG
o+A7Wq/56UwGm/hy/IEP7vz6r/LOLYdzuKZFNWTZv9JOppOWBsddOcA+X1ag
p8MCMm5jqlJB3Oo5WxfXt89hWPUILyPQarwapH7bAiOSIYghD/HtqXJe9dAX
7uGdGbVYT8zhwYF8QambJf10DdKbNyN9Vi1LFhGFsTaNQz93uLnZ6vrlpL98
fejPmIsiO3HOJO98a3W3jYMznTVBt/rE8pw/373ef4cPw8EfGTt1Z9xY+70n
H3E96PSDG+annrE67k505GX+rVxF2yBmSnfSiqQhx5BqPYyylmbyfHP7fZK6
r/Q5F34rN/OEjDDkkDxUzQP9R/moYsuHE4fwsrKWszF5plZoPTJyKCkb5dre
xGWsFuIil1wL38jgaDLVycrc++e6yrt2R/ZJOEzAozsfkAL8mcQqfTXWGB2x
/+wsAO36n9Py74mny6hv++Fb5GHzo2ENdy2ZTQ5h2AxvSoN0k7jXCpM64qEg
yos4Gd8dhKdcntDwYABCcYUVzepgzVrz2uc7mt5Vxz0qxlIzE8y/RqejeMce
z5pDrP38yNKHcAag4jQLNvZYbEemPUhBx26gwcEHKbFTTSzgfABbWI9IlDrW
SWb3NFqQ2fKSxCb80x2rlO8fqx/IKPJw2SWUxz+mCJvO2s21QAh1aje4oQ9F
G6Dv5L6loOGcS4Mb6DKqcFjWKN5XS87Fbnm7hhjRIQXtck94w8hvbq7t2FDn
e1BlePUPvk/CXRfHmDIf+GCmn3/ZruDqiQtWpZpa1sNgIVDFAWjG6z0LYDtt
UxqhkgXrimNhpDnAl5jXlITpYig0Xmmn553i5R4EyNVIcI8HO0gjIa5B22/d
1LXN1/9vmOPRvYC7sVsojoA1lb7E6L92NecTq5Jr3gk2gqIYPgMDybFVI/iy
kJsq10r+cmDGwwoilyUvcweON6wjCdeOs2t1DvaBZkw6pXDqejue/fv+DUVI
Kqfie5ggLyZyf84aUthxAyfgiwCIVMVYAmhULOgKrFDbXykVx8SOfBS/m+3U
Yn0S+0beioxtyJ+sorFC1eo87T3bZXP9exXlY3Yvj8Ign6x+viNCDFbwVqu7
YbTUB7ETaO/FsJfqmEGrjOM+g1tx1BPpIS83k/O+VOdoosfcq17QqcKRXZJO
GMMVDBGrhy4owP2IQC4GwZtAmsrFlZnTPD3FFX/NKX6oGBDr8wXCaHZwZN6p
GObMdYSpi8qsU9TuGWm4+zgZ5jW4g8mcy0tczylss01hCkRd3dQ3NjrOTvtk
odmsXZvezG5u/6UWtNtT0qGNX5YwpfSzc362MJxd9TnfAWOmpKuyinI4vUoS
qm8Poi31c3Z4A1VIq0m1HhzzC+p/G+0h7mTctkHXZcsOYCRUT1gxIdZKEe3X
iHTGXewiRGIHcgQRyOPH7YqG6+kRBvLOakrT2HkQjUABi9gVpnzjTeZHDnwo
9djmNyNivj9a5kniImYwuC1nvcc/9F53b6wwWnaepNZHjQYvu6DwgoVji4TE
mdzezCSFLxuSG5jg0sJT6Nke8+g+BP0UeEhxzQPrDecioe45V/fE+3rwO2V/
5fWLjQFm1lFiiwrp5CfPKsPjox34bijrhBCZ3xtZBlVimNdm3XkSSzjjJHj+
ZdaqHnCGKVNik3XCs4uEARVkxge2CzVQzlNa/MOfiI7kSh0eXSEIMWvG0cT1
rduixVIriP40HTsG/8285tCypy4xTMd8Ht8zulu/+QE88H7lQA4mHGuZ3PPp
cQx/i/bBal0un2ZOI1tE93lPXfLEvtynflP0zZNpqOIyRHPZSjFBx1pjByO8
X1EOJ/1XTnkseD4N9CQqe6HH3guH8IBHXaLISdWqIjWmtSiuU7EFYzqHMo5V
bl3d8jgHEEgtu8Ma75wPwKVGGVYfOtVrpyE0tgdtPSWdQJgfyJ8q9umGP8zo
+bBDOyzYHd8pCPOIsuaBZZc8H6XLj7lEPRFfv1/v7K/kiH5phoGR8GXMbv/s
WyrUgVUX+gPyZSW1zascqaEsy9iRvvBlza2hNfoFr7VLE2+z0a1yiJBxLbJb
UlDGhwh8yQ3FJ6qrFwMzCbtk7G8puCgWD1FDgwif1nUZf3DTKIi2xT9TeqdZ
y0d07Ns1z+akIG5fALubJx/GCLGxRULS6UPC0BgUc41lQ5Bdb8Vlwsmnd7Qi
FuLhzQTxPGqdPyCBD5yDzFxRyQe/5zTa8G8r8FK0GDdKq+eQ9+8uEMYweIK/
gf0zdJuaTtHubn2eGWLN8GhzUVejuLN8ainXIpyj8Usvww9WBi8MK1nWBiaZ
6eT9XYsztfHWgqVB/tTh0YBQpYheRdhl+3k3KkPFqh5y38NzQuhiOF/mzjDM
RIil5IFyvJDIECwDR4h38x0D9AFCeh0cR4nXcy+D0+TmwiQbg5B9dusaIbNj
A0qREU1+2UL6924Bb3HCXlSbNolvNjXHbxhn3gsiw4subDGb3FoMFn6ZYvV7
z5engH4/VcIOPZegYVk10f84bZty3JTIQSy8MXxQa3FHAihH6S48oqUwsNGZ
JfdpiXV8HKY+CHparwxCaSXEa47RpKrByHWb33dNacV/xBAnZEs41SBDbrEV
EQ7BDirMUxiMUGtEyt23hx2h0L04jjnpRSvec7cuRREZPQrbk+4bvh7vxYUk
+R2Z2cOiwlkhJTVkFLwr4wYW45oZduB7nQ8rmlG0qKrgW7IH/VNwnBHYEz+0
gilnAkhPuY1ajisBTWXdDA3FCVtahLaLrbHN0BzCq3phNh0YYca7J1wCo9AO
Q6Lot2CXBKJvUD/BykXGD9KYcgNxS9O0DYuWkAtOwYd3lDsC7Q6T1A1TtsoE
xUYB+pMYfuPtpocmQovjR7Q7WtpWTOjqhPxFC9/mbAoBO7PLvIPq8k8XU4aT
jameFrrGYv5+UcPsyp2A4I1/agajpYO9RYosjI9PmpbNUNndEEp3qdZKR94M
ExPVcDJbdy1KFpf/WKQUpbSmhNllNoaqi/B45C0nz3LVDUVHxnBZ/ooWok2L
8+r/CkLwPkrkWiM/bZq2sD1QNb1bNfCKZMQc8UOGqRElrLwX+XyJq8343ISI
lxpKu1Q7E3i24S/iJnDz9GrXSixaAHvqJcLsSE+1ew3sEqnUTJdbTvmTTKOs
WqOGoECUeIjFjIHHI8yJ9rJ6qIePiO5pg2a3wbKqjJ25zjC8MM1xzzx4KFC7
3dbF7bhCgTN/F08pJpVTUbslALrGdIXRGuAbf31WN2nUFx4/oa6cMfGIIk1y
eAuWj5/TbLF/LvwgMySB1mYug7UgyXKwVeFUbsMg0w3h7m62IzQjLOk4NIpF
JtufO21b6DHeFP8UkzqPnWxhV7lI2MvHx3RrHxDO0Rd6wVehWpTeOMi0qsCz
b9ToUvB0kO7CCIN+IXQvTWQHVrh6gOksK9ykRFuG3k00QGo2S01USfUUg2+x
rUKZyDhEDeDXUrDf3TV5RXJXpdVDxsGtmm3OIpv0sZY3zBPUHRUnEZZcXQUh
mUmcG/HE88KYtPjXEPBi3A/XYFHep5pUHlVy6qt0xNntcRR8aB3bBIRHHZ0X
wK/NVjDfntN/qCIYYoFpYl90AyjEOl0mitZ9zpBdp8ag0gRPUM1lrcBInDMF
Lgjq9TaHOKfQEMEY4lyhnB0CUWbym08cp5oNVhXmQIkrQ+xZLZ6BNJIN4Y6F
EukvcnoIrR8aWdm25XXz9nXj6/ma7VPkTSD7WT/hMqndZ71HdiO+yHDv7YwF
Ib8LxSPwgqYA+cUzqNJeIlnkBIR3pz/JcCoxfxvf9GpedzqaT9WCmGY3DDHJ
jeuZsreTssnmQBRqZv6f8rVdY380gMdA+WwDBBqBytIENE2iFXwzicw3MdFE
aA8WooyGxhJWRuWnvxx1d/1rhr9dUL+89wyO5UnjDE5X51K0qdb0lhqyPuAN
KqNB3Ij0UPPR+SI2+bEpn51g1H8IO+y3tz0G453cBqXsTY3GFVRyZ5KoP71p
Bnu4aOrjVszIXvY7MwEbwp41o9eVtbuX/SMqi2V2b6ZdhIHC1uQ5IuaByO0S
LsJ9eO+UXJjfJW9PBrj1tOxCYNSSUuBPf3bToR1RKbQQd6nfcc+5vm6qqGWV
4qIVdcZVAw9z+I/XpZaUX6f2xXEvBi0/ifCwKOX9UhHU7Y9l2toA8W+Su3IR
NbU+XlIaFNz5GqaSeujo9oYdUwwxUObXTDV7VZJ9nSZHqFMApF7XjwcCUm5f
gMw/CI0vLfEf620rIdXtDRmgbl7GlMudqU5Sck9OjEOlKaw97AKWMrqTZCel
m4vQhf6aZ3qkGd6YnZLAB3e54nKclwzgYfjMsRjdcQPxPf4c0yKqASVQZ0tn
fIjOxLpDwh6IXbGQLINGYQ96JFAI1mxTduCEmnjVnrw4OYxBEZ19xp4zot1S
m0Mn5ecx5xqddvcyKxpmriO29jCIhwOWdGF4Q/sdaucrulPYf4rxCUQvBC+K
EYT5UpormuCnFKr0EoPCL5kGHlFG1tqX1Jj5Z21NpPhsg5UpYiP/qHUAeqhb
U/EU6FQOwWa5XOarnLKrPV5V8t2NzXrb8K0bI+JUMMfuMUIATDG3XWZutORB
sZdQpF88rtvqNOBXN4uk15sJbQV5chEJTHtfxJfU/QXkNST7O2spDuxqU+NI
zVy4/XjKtiK8W21ckQ7E2m2pMrUnlY/0TA4Vcz8yxK/tYZL4FG6ru3TZ+iRb
vQrfwlSXO+yUBes6dycSNevw10ko3g9thMeBAzCja3372odFEug+wmZkvJbm
lUfHmoxawFyyNfDt4+wNiRXkwzEcWoHOFROW8q2F312RTxKoMvM18PiujSkw
w0zbPkAP+z/ObvUCTR+pCFLx+gfSeAuBd6UpS7eDFr8dzxQth+h59X/OPfhW
Gc2wLxTYQfGv+/t3GbMBUbYITBjXMJXlcmcFp1vaTWvSOZtAKJLQylBj4Xxc
caX+VI5aTFNqWKJrNFGTh3FJNxuRUzJJ3pMPK1HJkYpNQZCu5UdiBDBP9I+v
4ewejQyIBzwx8pOaDF79pGTE3H0R2j6eoMJn2QiPFR+9+PT0Xod4DHYGykcB
tFhgVxheoHwMwNQm1aRkdCyDdut/T5d6yiAmz37EqrzbfTON1ufvW2w4lmnw
wY50c3YkgEW9y65QiXr+65/fKukdZZQrVB2VRKpD7s3M7WPXqJa4Evi1SVha
yBY4xp69iq9rIWHSx6gmRnx0jzSdsl38LG+Q4h9Yv3QiA9Q7NhpDN2BLgACS
2Ol88QaB+82SHANohc4Ws7PnELTR+qkCW4upN0Szw/t2ZVre2nXn89fbwv9f
aRPwiZqb0p6Z+0UxlRMLVBnv5TEVaxsy58CHK9JBTFbDzrIoat6GA7ZDMZ/f
dSt6pD8OaLvkaP3tfbZvIiH8Al15lgVyuqxdeqz/9r6xLn6rV30oZj9CKv1s
iRm8aLyepLHy+t16kcn/rgj8fWTdIt8oqet78KxJXsMWSBwScmu//SZFpHQJ
OAhyggh3aTYFl5Xkqdy1wLdYpuYMl6iP8yWxkMO1VwKetjIE4Z+O4EAarlny
DKb64sF2QURoM9/JT4VGKljj1B7v++AEjZfMWqBTt0lwGQE9WcYxl5afLGYy
RIcG2mje23VBGBJKNChss5gaueLmKMVZWA+xh/f4msgI3CKS+ph03CTY1/DD
9o3TOlOSprmnqLJTFqizmyU/Y5RpDGT5AWAUIuqKwFaQ2336A9wt0aMwcrj4
0mf0QEFzWvxEM+AzCvgweppVg2Wehddo97uqnqwwUFBG+Yhh/Pl/WBqyhRmk
1pMbYXBdOQUm/wakaDYWI/UcYMR+wjdOx0kzJhx3Kxd5W25cWrvoJMKMZXUX
ydSjee2oH1wkHhbpP/FYpHFl+U9JhZmBtsbQg32skH9DfUdMDRgNzj8UWXCw
++szLskK15Mn9bUPh5Gd0z6j13Pzd6vR4dQXQqOsvRlTGfKaxxY96aKy5m6J
g1aY0Kqgf8HKVLsVdsqczVXqsdT6dz2ZuNddQvlK3hDH/zgVbXDMbwIKOlz3
67xU+1k5VhtVo0s2qbQZUYOnTtHCn52mq6lo70xSjPuNenNnGOakCCq+6hTU
95VjvkoZ0zvtgEbLsOqK5UKEV40+Q+wSEKEdbq17wAuC0wAvbgchW4Q7957c
hC9IEokUtqScyzGXb5keRgWaHEz1mDPTQimCQ5XVSW8sOXuwFT5uubGXySMx
K3Tp0fZR3fkwH1aO1OXA39N43Gfke4KZP+EfZ4sZYV1TbAFbGd0Xgh9j99Fv
W0kvjMUqA/NET17H8wLdf7zc9hVBdx0XOyu0KR40y3ljEXGKXd8PPuyXq7MA
OCklwXFagZ8e+sASyMj4Ztr4lDbaZLHT7//tyLtrV/6ZbP5YQkUQB5Esh5/N
ykze18Duiae56tId1vM3uY/yxKLU79DhFScnDYsoLVQUZ7THN/t6PkRfBcEY
FiVAbrDs5R7R09VIMwdMj21/D7fmqdKoTMX3DryK90sqsEnfUA23oxwwMAn2
1gHoR1r6g9bBRFaTwnwYFDHlPq3CQSLXip37InjJFub1DAQNxqEU/2USUh0e
TPZdVkOHyBpb+V1nYp/EYZeQMaQJKeYRILKAa601u1vBIrKmhTsNC+R+kphU
UyKSRj8AAjHdOWnkHYQ6Nbqr1eOuprGTGwUxvOutmMov8zaR8E5LPPsYcX7p
wBDG2WtDeH03BdRdKcpXg8E9Za3IHfINYMAbWfJiPA2hGCBrCCEgq3tsA+p4
lGzvIbBa5NYDjUyTg/iQMWDPSF7g6jiyRqAVQ0K/ON/S6dsaO6taJ94kTFHs
fbmw2/BiQDFtHlV01SoM7epRL45qn0pawO5ifEzUr9lnB6Dbwd2Q5VODKvEq
uExeDoom7gr+JCYoUzvIk31+ugj/r2Uan00l+l8zvLw5Rmy0RWwltiQ2YbjM
n+kbVSdUeUtKz/MdWErlXtUC6POrAss7tLnR/t0j9UuvaASGr+d48YesHNI2
XEqC6G9ySr7BAe9foW3wj9J2LFX2iUK+Z3nB2JjNRgzH5UpCr3fBMGHPa5a/
v5JbBsNOVb2LamOuzQhpwZFXmt9MImd//OV5g+l6v01wvRM85ZMpUv942rNM
5wchHCOYdpE4bgtoXAdZibb438QoWs7TWicHf6BtqGVtx0EhZW9RhIDISXbr
rsVKxjghrJliIkPk1n3ONmO6yhLaeJ+pUSIkNaQLmUiwIceqUSLxAOAiagnQ
G4QByknPpuiSBK7VSJpfEhw7miX0LDDKpReoE1n4v8vziCkPmgQaiLZg+BSR
Y7utaTqH2EpLBgQHgcryi6BflPSJ39cXou48o1qqoaHCcxKK/ZfqIAulG+tA
X1jpLfZAvKjYjTf2uC6MzUlSYLuUxqeNF3HThu5zUns6vlNVEW8N4njmcyqo
LFx/G0ozd0thB26RGahhuTyXTsVXvx/dtgXrd6nMFrOpKOcrv4QzjH4R9GpO
cyUy9AxSOqjsx/z1wCJ6EzXn2jAi/Jit1fQtAQTqNlXHlPTUALn3wPpbQiMP
jyI2quWwDV5qY/IdtN+h5NTKbc3/hGVQO5lG5RjeG5ckBgKC6he9rwWLZDp3
iU6WQTcsE5ZggD4J2ZoLtCCjvhEHOx4EqfhuzvTkJKgRJiPM8gJMvCzhCtrn
ToSL+lumTz4Z6ry3KkIN5kUGlNrFzJt+uJTnrFm6vOX7izalM09oLO1zdCiS
OJIUeAfZZTfOU1WS/oE1q+OmyG2eaK/mbN/IAJyJ57slxsE/x6Et+Hs+d1OH
PgfIM1GD46ZpMjNKKQ1FK3oHD/QQC4dTgKRISPMAKJc6xfkoFCkgM+Qxwh83
bZLlQOcsqkowDEf2UIt2UK/C87Dhs3mkpErLF8TtB67cXLpQpgn3VCmSD513
u1xW6HRs+rKdf1lqEJUEc0aDiRdJp3sFN4kcgWQ0r/rbpHdMXo8PeobW+moF
abY+x0f3+mCNeTGZRHnFeYS+qRXK539tQtA/utAP5qEnDxodrdYhMYlxAB2r
O0tUCLaSV37Y1+hJaADGCCrf94csfWYZPtGjS1j/ByF7qlnTohmJy+YvJdiM
oedZFkDx75dHDPUnOaMeyvE07/rJd+Y/kjQ+aLczB0QJtbH+QyIdirAUbV/V
Oa5WeBUy9WJIf2jKskwlAlzX9/pFPj9zOENAwk7BFyxCSJgQXqJ97TI1nFN6
YLlBotglN47zLj8ikmArmQE1HruqSLvt+M4F+usuW6fT3Nr/wjDU0vfZrRgs
GTr2pYEADBl/BDqDVj8EAEOuqVxKNIJAVAutqMDp37+icaRKzxJ6iFlmUOSe
belWMj5CJr/+MuMGd2tuNGvWVF3VpTgRvdLkdTYzyvI9T6E+MyWJIW6jZAAc
41solEEHxBG3mlwZGZhrjRUjnNSJQE+q4bHYdAHNrzN9BnMoCMSTiovGVlDW
mj1l6YISW8nS3Rt5EhmkNqwNhhUXVYPCPiqccEKgooYTYpVpLC+yjFggz9+i
zLj7yQVvTUqICWlMtp0Spbg2BLNCNr8oVU18x61Gi7QTUhALdULmAhOTtYUO
JyUK6bB3nzrTXjwWtP5oPRRo/LbszOgXJRD3hJgCMI5ohURq4p+rY5zvk6h1
/a7/rr6+khbw1Xh2ffbK5TrysGWP2a2OlIJg3KHBgWIFvqAMv9KEdDl9g+4J
S+eRk4Y65Ibg/WetD5N5QL3TRvlxEbBpJjpwlev0aPheN36AkhrF/aHoMzQ7
X3pi0bXO1C+7zAfsXXtMSQ/WW1WWd4QIGe4kyNTvUSGowTUZed3+t1QoYR2M
TYsTwsWi2LBY4hjiMyO9RodtNHvv558bomliYXL9zmZrABCFmKRRZRB3dP2U
5D1YqBD5URdbxUfHD49h+Axt8TIv186+Ak2j7CV4/kEOMvYm/ePfMreFj0XT
0PVD1opuaTGWenor70+BKQce5vxBLij1gHkV0hjsdrWyzWxQo56uzOb3G0LC
B/N4lJSdoFBr+6oiI9fyZmF9AwTo2Iw09Y4LY3MBYGoPefQ70PhDnY8UXpsm
8EdJ01MythGGusT1z7ejiBMzZTOj8qGrOQ1YEnqBVi6M5MAtakLTSlZ0umw7
AjPB3oW+5mVFjBFuzVb1ZlnFzaSF6DZwTDPvnE/9YgCgSqTVcTe1pPt/qhgo
gkYQn9T/uARxSWoZMkRUcz0GfS1TXwWTFWaByP8xJD5w9+Xoo+nHr8eM9Tjp
UF637Wf/x9twmVvjtXuIECtvyiPO9Z3p5Q0oni7huMAfhh5DZKKaJoNS+PMc
tCxkH6sHnoJShSep6Cb7cgdDU9/lVK3A9Qh5zFB8qd6MN1w9u87mAgzw0oUc
3pU1jPGRatiJ1l3BxqPqwTgNHYU4fzGqZTE0JJGiZOYiGpE6x2Y/Jxwb5/h3
XH589TNZ9yIDzdHFU7uEhB6lQgjqNkTv5GjKEUbGDsUxho2vKZKm8tWKMn+v
DO3FcG8m/xXAkhuRSVpcOe8DDBr++K6D8JOs/A4EdenDPCBUXk7XgFWLlSJo
ZY68qcdESc0dHYBE/WjBrms2dee5VMsFuXedWJqX7Ow6lIfatQF+Az7EUZFs
687VKKZ9TIp4OSR0vnuSsLVXtHE7irCi2mcM9LS6jKUuV36ktIzyglnKq07R
MzqgTGkAtFT1Rby5tjJL9eU1VcZa5TpdP82YiG+j0Eucpzaoq37OPRSnSeOm
CuTyrBhfhodpiGxL1Q361Y9q6OLXFi1XOpXvRAuh54zzMWfT/LwjEytdYEv7
jr6jMqSbZdbFhVcp7jK3NsACTne/YhN+i8E1FGQVPeUtKZmxXcZqC4D5tH7b
aeSwa8IwPmoULQgqLsGxbdw0AbAW6NFuP65gRbVqYsqtG+cWBWhceSezaEhn
PZcrAN+qr0+y65pf6hUvLqNw0ucpciX26vFAHvKTGpUhn81DH9oL6aO1fL4k
abW/flUZrfcnwNGfrVAKkhyrWv//3zBvT1GdI29rHtDzs1cMNgoDnEWSpQDj
KWDA0xGTMfZP2SwQ1exytdUSZQPBhltDUm9s4YmMr4GvhgRYvdEoWtuXl2cW
cQIkFIUFyGQwO5lzOSP4ov4pJI9Pq3rNnJyzGPQWR2/wbGiSlagYBYzO8ipp
2VctL5GGS5lo8NR+gGI3PKyB4S/9xHcgZ/Cv0SIccv2YygnBqTTYbvKx+38s
QaMbchIfHCoqUkruuYiovr01deScwHwAhC06DbwJSzavBiXggH/MSQKpWZwp
IhTjBMvP93deBwV17dx4Ptf24+Jegr3VHb/qu8xHgQQENOPIaL318QZMYDYh
SbXoD4V8I+POSqkXAh6kjTI9nTjW3USnj4MhgS1bL+aDhO0txiCxw3dErOtQ
2I/90gjc5EZvqu66mEg7PhvgggtYkXED+RMQKk2OLr48lw38rNuVG7xqaY4J
EpUODZZJ4dGA0Cwv49MJYoqCYMMcpM86DRhf2UJjcEt0a1/yTF0WrUvWvR5W
dKluCEhDuDZti/VyDduQuiZNNGeICANItxrlatLQAO6+sQIvh0TwnijZlH0X
gwqhjQN03e3tsaRM7gApHGjWVvXwxwScW0eyhGMtBBLnXkCB6g6yyjWlXds+
Ji3ND5YF/yO//UukcymkWwfd3va3o5JSOX2nALpUvNk8MwOKPz5+LmumAvRr
Yc+xAZyEYO6U7dKhmJDEQ5aR/TU77Swtrrb/Gb3PYrken+TNSGxdaBEeTP2d
hsnUIs/jrtR29HKFiGS0yfAoy1skWbt1E3/Qe9QBO0LEwZl8X0trqwaMZzxF
5HuYvTFkNHtIKf5leHzgePNKVN/lts4eEowC5cxD/IfYXijuiSBGv6yDOv9J
ZZWmUH9n9di/lQ2ckR0UuyyQUGp6GplyivesOzis3iDYgd5nYJDmZEp3zpYA
rThJ7bhQ+FHSM9X2dwDJrSex7sdfIJ9zE5qxYRSe9fqH7yI+eJ2qSAvExSCA
GZZvWbUaIX3B2pqSD5aI1KEi04rkj9W1fipaZA5Imo00qh3FC8e4slT6vX7u
0Iym0hFY7VC8Sa0r9AWZqYsqX00d8woYEKwuIY9el5r8pMS90VqaYHfGTS0V
qHM3JIIFwjsv6CXeJnOyJtZn99xtHnbZRd6Hc0zSs4SrETWkpt7cKwWCe/On
a8MiXL8tke36pTMBHd0dDdYUNTBbm3g8Xddy+IHIwOAKsNPzVadpMIOaqIbN
1XsMBdmRxQg3a2tyEt/rWunnQnj7GFwQU2yNcgqsUdyA6SHml5zyJM1hY5PO
sfxN8tYqF1YZoXXQoTuGi6TK9+EUBcjKpxGytadizlZhkyxOGNgLtf7XMi6s
majJ1gAW8qPMV/wy2/50g0GW42F2vbuvW0fnnQX00FLRzG150fabkbGAf7E6
kt9scrb5qWRbHxcxZEaoqrk2SBjzBfKph8jjw2lfrgauxv7W/JR+lXkhAkew
0tjUYcuD21Kg8vYv/UFXh31ced3otw0M4h62seYbB75pY5QTX3FBrOIwadER
gjHJQCcOCo9g4Sca+4oZvuJEbnA3ERUduyC/s+n82Ei76VmsJeePAlSVNNBQ
/tk0/PhurbWT7SbWHmNa8ScGZ97pMoPHnnzgTaWd+sfwHb6CXJn46JPJrfIl
5rxP8iYtV452BAHqWW2OXk8dlnpo4F9pRCWyRUVoMjbSJs0pGwhmMxh5Hqsc
8+hBfcG+P58rug44Bgo0E73nw5SI4k+QFCmTHfzPw48xZbGWtwoC1Kn8Cqgc
0n3b4e1sqH7mAUZf4StCNgFKJVD/NBIENMESHqvyDJpRAZA6x3KZxxs9zYkr
rQ09RL1s8oocSiiNUSjKCL/NwFPW1t+ulMfyKZT9/o/1oNsL0ejJ937OTyP6
54h5R0rCGle/wPxLdm7vnieZKC5PwNxWSyiu6M9Y55K35oC4LGtQ5nL0TgLO
ZHBXzu5erlRHKkzTYlw5pCPG2YqVqtalf/btC9i5xrxRPOviO//QYFn0Wu6R
KjFgmgjTnea4Eq0I7bgKcmGHaQ32vuJRmMXH7MiSkD5twMcYJRdx7qOOgukT
4sWcMvwv6TldKbW3Lm7LB8wauVa58iJjSNzzS4Mebdq3mdU7l8JkJ+p7tJC/
JHG7w761Uk9TdKChqILjRrQztIvyUqr9fM3pnkzlqroiRcXtQvmU7Y4Izs0b
x94ua2mM048tdkK9uwETw7DqSbbuUmmnVbgnc/MmRJdv8wo5q5oqJaZ/xt5F
FMVaSpaeZvFDe6kF+RakU78bnLcnGmHRBFDiYsKP8NapcVc1omOK6mLjK5e6
QGia3a6yvo4CylV006/ZcjeWctiOXNLHFR9QKxybW8k+TqY82YSme1GbIsNK
10lkXT4sgM1cyPTIO/zZ2hI17Mh7G2fMvHe9+mc5VWqVjxjpApaGnp6jwRRm
rghCm5mzC+85ywlMaT3g05G4eMe8gLLCfy2U2v4uKkr5zxnf1xVg1Gw/kcfl
vqY6cPWx2qfsGFnu9EfxyWA6Ir+VsmGbMWeR+qVwnbKHRdHjWKk/elfWScLy
DypLePM/of3IyYna0APmTvLsSM3p6s0Qcq7z10p3PnEACVrZMVANtD9REPXQ
cVuBPj0IGR0mjFn59I19qPvQTMlDnFMe8R8OSYUC9heP/C/mtCIpDZiBIGrU
PnuBGwfbda2m5+UJTxplWYtXjKSU0sOLqSlUkGGUmLhQSyUpXocEXg56djSn
4r/R5ae22EhYraMUPactjDPtkwCyNGNV/r5HMt5RUcZEHEahlZbgDw4ieXlr
ikTdASZayxAGrRZfA02+wPRSpnUEJ1FFzoERAetb7pqE7F2i+HEG7bWIOPn3
QHcAUIIw6pO5zS/eXR1sgCwytavdpkbRb6sSruUTEGYoNop5elS3qVg4HSXC
AJNfw9JMu40Q93kYkfVTZf+i/s7PQPA+yMIqEd5CP1Nq/xu2jJqz9adIN0Yy
JyMnGQkMjB7tcocDEmc0Uzh8nc9Mal4RJUe44aw17VEGFOW2e3XtmJCARwC6
5YfMTxSbCGqP6Bur7yp0IG3fJpVBs1WRJPzSi0BxRMRWHCyvYyVHEh6lbPn2
YKDoX76FhMNDLwOOkP18S3Brcf5s3NU/WZqKI1uFyB2DaMXBBZrmsvrnnPPD
u5NL0TQy6v8bUEaEeJ4CMLuVihkiPE9j/yu01V8AB4SEy9B6NMX0wPThI3i7
LNX52s92pCUIcuoJv5gf+W1BIB0UCg/ywm6vc3zNW9lgD5JFKpsTpW5BF/nc
cKa+lmkRL5qxfKgUNqLHJkdTGf8CTtWwfJWQrwfHf2Rrr5mDNJsSU1VS4Lu6
Z4cfJn9wgwhg2B4lHPtZUQlAL3CNtbvPnJ0Azi4FZnt1OVESoDek/+UlmbyN
3PwMoTjtx5PfI+b5Twg9NaE+FgZpG9MZ0MPjdjPl/UrmA9ef1rIxc+43C6af
dChlLtnTUuBFsYFscHohe8Ew7nfYPVhcGRIDs1Wvaoj0qAgeWjMLJF8V1TT1
m6wyoVnZGuMiZ+xwoGlAiJkf9AoAzYYeRckOa4Zo2YDQSLFxFaQ3OCjgtWpU
MgWe4ifDHognYEJP6pREYCGhv8ukdnEWi9l0Io5+6gh+5BHcePgZzfUOeGOn
6jdSPX5N7vBgxFT8HNrMCurHLgIM9c6zyQYhSKKOaF8NEN+0qJC3P2/5H2kC
RfRjNWUpa5J5BWTEr5XVBp2vxe7Rci0olPEGjZIlQ0mMtz+FKAcquZv5mOia
OADU26qXn1zVUrfZZUnEW9nccbfc0c3ehMm9DiUOyD/7fuyF/xlqltSY+wwy
R2gz9QNoRhnxmsJFvwasI/Yulgkm30HotGzKBG9JV2UUmZJWRPCSRWnBtOZG
eNx5tBsbELXKaHbUrsUPIEc5qow4dd+KesF6ktMHR04Ek4rv3Et1SSLS6SgM
yG1gBGHlFPqr5G27/nV7IniO0BH8Tu1kgzF2Dh7i2R5VcFUvEiPGWaacDxbt
99hm8G/hlWWCINlgV1lSMJ3qmqu+4Mh3hQ8hH9z3pqv6XvRWJrdO9xgbX2RI
oAbEmiyfA+sGcwDHmgjeUhEmVIZGAH2UYH/lcfkuaV/xMXUl5Nae6bYK+Yte
21S23gj+6GYSy2WcYYzp1IpMmDqmXbUJyDQd7XMzBTXjV58wG6GbiezEDRcb
7slIy4sNlZoY7KAitQ4YHz9vcLr2BMDTb6dFiyeChVz2aa1uikyjKOZqHnR7
qHPC4BzXcPRS3IrlntsuhbBq3FxC9uHWFtDQOVnqb05F8UyK3L0/VfCyBE3K
eDPMbgg3LRO98r5mC7hZaPj+1zWF4nq851DYNaCM6oTgmWE98EQzyObTAro4
J05YeZWS2tYhpa7ORRemnmOjjMTll6wG0LZiNwo1dmJ2Bvne7ZySMLMIkVCr
SmpCLnYo28BboE74/3MBTOGhv5Rg82ht8fb+xW3J+4DypXeXHonVkNBrtzBe
apPm8Gnv1bE8EFhnuzq7nyAYVTKv8O2zgAcb0GhAywPkZbFyIDQ13BnxAELs
/aWCDWYMY+cUHbnUis4dLNx64hpj3iSbMN+EyUv3SZDtwR0UjvJ/bc0+Gse+
WERQMw6bwO60uQLzDU1ySgBEyAaSvsjMVCje3kZj75e8HXjt2PRBvwxoJHLD
8JkLTWIO3AqltQ9r993ZFeT90W6vE/HrPCbA5zjLyZxBLRFLp34iZqNPVi4g
qED/JRnCCCOoUOU5SKm9vIdNxfuhHkqcQSpV6dPo+VprkAiVCGSUbvYMNdMZ
nTjuNDbejLKtlAVokpbh2uRr4AMMxjGrgDIq2LfbCGhLgxzs4C6Gdy+neqpR
pNlJYVIdLPiQTMy6OZDix9n2SBKr+NGfNyBDXnr6JvcxRa71U3MBpITDHt3K
kt/yGeY+jZSC7f9ys/lYhsCsJL5wPyxDcr4oar2aXtZQvy8qkZDalkHaek7D
k9a5uoTH3LsEPHNck7ps5r7O4ON0ngVpKgBGjJ9Z7saLL0UN12l5NrJL9Wbi
tUDfbGzi3yIrfzBvPwthqiEQBsOYUwgUKkW5zF22MGvAIdQEJeh/X+4wGPYM
67kNt83wN7BUOixQlWwjf8pYv2oN8x+y+BlQiJFgN95XTlGuG+pfC36y41tf
KzAT9avO8goqv0AVzYuMqmsjaSHGm40gIDdHuYMT/lJJEFA+/VzN5EAfavUe
ULCCpfzxwgBp66fc9eoPCypsmk8f3p6tmp4bNKfZat3TSyvXYPr8b6+mJe+n
W07v9iMeO1U/lRj5cNC3LjfeRL37WA5OkZUCpjM2ZH5pcFTpMeXBEnFxUDsx
6Sr5abqEcJDUKj7lRLV4grhOeJpyUwArSvbUnucUM8gu61sIpVD9ysCzTy28
v/+8kcctpRnOL8NudvJFeauFHOewU/kPcn3bPapd448/xX3UPW0GJ31oCEZ4
JQ4n+HesfhzYLvEPS1B/d7U2ELQ/man0tK4dBtmBd4pU9MFjCMFqJ00aa3aY
BYWv3WG5DSDWjNTQFliS4jsv8upgy5Efl12T26jFLwi78kWwkiSfhimCppMX
dB/U+0jhiU574JnW42Zq0jOvqZIg9aYFqc8JvMLsioS766hdWfuWB2lMXBPv
e3zyFOGzTui3WBGxhi1jBRUaQuZfljoUWmP8EoWisg0BUxVJdokM4MxqihlB
XJRT3ZYPi+pscfesYunwGnsQpfu9cFlcPDRu6cXB2Ddvc2qecpe0I6QpMiPH
vUZQcoayBqsWz2miUikCwmuf6ljh6UcEw9aPYt9NghkZ4p0nyQkVikYcTPba
7avwM8SgNfWQaXCGsNvy0NpTH5DRFg54yAXU3AWqcpuFbixtt0HxhCEzeWLL
qUNM3t0i4JoSYDCGCmzTJFyA82Otw2C1HBrM52nPuZjL1tSNPd547hT8rs4z
gilWgN2oy9icML5d9xr401h5SmDrvYDPbpckQDIuzo87jbFy4/s+JL+5Vbk1
2jDmEGzM0rI+u83JbSCeWlHl/9wAXvNCtn/o1mygkRGByhWzi0FXePx58+4b
lu1NL+7jv7sCbr21ThgmtNyC5bmgCLg79l0/rNOxQ9dX+DuLZ90U0NWtGth0
aSEu7mz3ATYo3F2/m+2Ck6yWHAhkgGunPJYlSq5fzuTZEaTughpFgrQUooii
4vPzoPiowlUUTisK/IpIenX1x7zAW/XgdImNPIDTn7t0msDFcAALs9n3YBBL
hpUeFpw9E6Lh4vsU7o5meNHSC2vYIYiv9kwfCI6rJuoNM8U7CJJw+If3SXyU
8OmBpaNJR/CXl5aMyVLnbrDkoZIBns6BAyvfp6CRjtlBZRu9gLpmBkHc9GmD
eYv8SK0zibuzzt6EvDkUqyHG9wZju/iFP8eN6vsCMK89dc9LtP1/crrrskmA
pd59BgUP9MIdF15mtBzPBcOfpoKIRX4veI6RjIV820iEnnmrhxnOmR3a3gdO
LvfAmElJtoAuBw7xxj1eSWknC1VfrBtcUBndfyvVf/aKNYRZjLZo9bJup/qp
cezuE2QaUGVVuTp/GXJsp9H3JeZA9ofrxFmlc4RCtFwGoEKv3MWgvY63Qg3+
KpoPS/XoQ8fV6o4wVVxR+q7K6pCK39n+ITPQIT0m2zkMC1+AzKJDJQNvp+Tz
N/UktstZPcwNwjrUSDRa4xX8OoAeb82KMvx6F7W5AgRCjBuQ9IOmFyQeGQVk
IQQ2RHVtxqL/NXTOhoz7hle1edJTT6LR0HIFOVyZUTjbOKtY4XTh5fVIoAsf
+ZDSB1sSz7V8MxDq/uYKSoqs+nWs1Yr83OXWdOG1cjGbExVQdRigFcVLECUk
NagiV2SE72SsXzbsB4X0AKw7i9lc6f1yNVCBr6xNwCis5RMfpBBdSulG+YQo
ZpuYZC8W+TgrV9SWeqGQgWUSk6MiVbXQckl08U5qQ/hxqalb0D7GRinrLBpw
pWpT4lv+4y37ydiBkfr+NWJqAONklbzm30lvCKRWEdIBIG81BNxwr8teWT2D
AMCk2/TVEO7gLNmeSNXjB9H9jrjFXTa0WsaeQTrT9He89Uxa4/BJZRHssv21
wg/BHN9dvLlQ3RKewtpYy/BKhzvfZ/TYK/H1geFWPfZn4QorGiJ1bJt3QAUR
GqR0j1YfIZaQqzeYCRFq18OZtby2U2IC6vDs0GB5HnESEpU6zVbScaxjzaPR
1xcz9lp0qE2eiQD4eM28BXPoR2FMHl/gnQg6EHmQlJV+mxrLa32DSjEZ89q5
hkjlctp2X1o7pY7tXEBgpgOYe1MugzMhmlV4fLXqUHt6fUQv51+5/L103gCS
Fb91W0XplmF+zyV1r6qoALNqexqlFhIUhp4vYwgCbF48+ITSkiludZKmmhWy
zmm2jNpRDoB+0stPTTFIj/BHNFNg84BMQJ5PfxWx1OI7cEC4vuIzDZjXbN96
GRomU2NxwH2jnz5km3s/MKWfOXwIOG48dEzQEATOQ+UqnnIeH5M7pGdKGnsI
02qumRRwtZcWhz21rsLjEjxOyK42RU+AdYSMVGIKcecsWVww7o6uqmzormaL
p0ec80uTKERCYdZeB1srlYAafwrZfqXbGPBLa46lRdJV1+px8M7XlwP+uMgY
QM3B0nDKaa7M2MLj+FsbyBpTgb623tsRWx0jpPQ9z1gu6jf9cGU3KvszHgRb
UCWEuQY+EyexAySDeVHSn8ou+RgVyOtlqA5SLMqWdCvWlZIITd+F9byvTRg1
NenNPTuBAk88h1fDY6vVMY0OWW6tzSlgkrzlBP48IoWe/KXaAfN2Am8iJQ5b
Hpn4d74VCBCsaQL+xrkSBZOq9Ebu0iXbxBMBzrsAkFUXClZHgiafqB0IzrRV
xSKI3Fzsu9R/JaPfQ74IeWzg33OV3u4ESyxx3pfxixT9hjPAU9V03cYXCog6
mUaV7GXmVWyx0K4+915dR99hMGcDWMATqNFf19cPEtWoDuNbR0flmVNamNSv
oNdpUIoRdS6UtODNMlxfoSBqYOomhLpJigtqkw55FNAwcyvig44qGYBGuIbo
eGksS+0pj7vldD2RyfozKNpP/+SM7vZVgVH7ItUCUsMM+QxHKnWJPBfDTrVt
zmh6vSbjWUrrhPghgFXXWsOmvia7sT/oY8mFrbaxhGxPVuSweInRhSU8uPSG
J6rRnlzgoagvs80CfL7TD6cuU8KSS9j1vX5Ud6FTjaZJTbPB7NqQ441lfWA/
IoxrmSrNmDfOu+1TC59Ygpfq6M8DxQnnnY5s3UG8Mct6oylOFxUVW23p1UQk
59pCXqulAQpJbV+uGE5ILjgNKycrOcKW3RLBDgVOg9FUo8wVosS1sHrZnGZQ
MVAhRG7WO4h++R9mF0faEcVH5gcWL1hfk3Ohm1YkBH5A8tnvQnpGlMTDxirY
krL1crtuTcfJc+1okT7Ds4i27FWA7sJRtQdxxS1rERpdVT0CWoWKjNtIwtfg
TV+3hdns3gSxKyNk4Oc6T/vFXS1z32ySEueJBMpb28w/42mlwugBgPEHskCG
+tH45XjT1qdEXhVZfO8+kkE1DwUlhsYgV/0xJT+PWt6awWc+LZDN3n/cVlB0
OXY00Fdhi+Bhax5g6I2VlJCjpt89MNJuu0Pc15udSRScMkf6DpaDJ3DgCbGe
4OhP0GDFyy2j1m5sKnwl9BHnlNpc6ZbzCy5mCJln849jXPnH4CqfdCwuV2MM
/QE07zrTKZ2UHERTpWmt/JQqew6zDLyMJJN8I6X7hkFRy2yFb08Aa45PrG36
sLKidJznaubYi2fkct55et9Y1iBzwY92XHCE1LHACayWHL7Vyl4kQpNuWvjJ
n2pv75FDdY84r6uztgQwHPU9GZT61uXBX6F2qIVIeURcsLevd3elFTXxl2dP
BIc9h02yuyuikunNEIp3rvhEtwUUzFW/nd05f5S2qmt/J42pOUDrVJJ6kdwe
KvP/vauzfGogEiimNIICt5lcllJxJCS9k2injagkWSzKROEEXgxaw1f+XNw9
IOt1LZW5EiHQlClnp3ww2HznUvCD0r5yJi0IkQ1pqwBitK7q3TiPzHXxoPdU
p3xHy+nbVXKzJEFYwOOQk5kP2DLN+MYCFdZ0w54usFTgaUTuU24W4evZTEZi
IqGsDcDd/qeMeXBwSRGqIK1Pvn0K2w5ORSsWaYh7Y6c1nPlMj+yKxgReZyMq
YqRjH2oIp/BHJdcj3za0bxurdlQEPxqBHagRgdxT+168d1cZYAzK/WSz9gmK
SBqMK6vVGoINg0Yausgkb4g7u6rswcZvQxDp18yWXyOIIxRvBjf+nhkExwMB
BbX5KjHDh6t5MmYw4V4UOD1M6jtiN4p3EIQnytsWim2ZWVehmFPtOS/3pmTa
7EbGaLzrgRBP7jQWE+aZTpHjaeS96Nnhdlrvb3MAkpSZ27HdLy6TvBOSF2+k
tLPN8P3d3CgvlySXDGjOjGV7DDlWJY9rbMcb75mXOt/gHLXT56KTtPh2B6P2
QIv/8/9LngpzcPOQ3sUebfOHyWr4773Joo98nWxi+9ZN8OqrWpDfQFEem4ch
0jol6jyS+gMznzsqd+bz0xcTXjwUnEkEOkfM416rzVF9ye0n8NykPz6Og7iP
jR+ieQsbZ12d+Gv3tz1CEXPkG6mJxp4KSQQIz6tTHOr1U7y3JxIpbxZa5EKe
QToxKIVtxm/K8knwSmoxUkY+Kxm+vqK1GvyEyA6BsgkCc/9zHmco3klUxj15
oBL1arD6CQC8qQv4501TUKPE3ZIXFH9d+n0NWqVj4LxMCZ+qqisy+zBI5U3z
Wf3QbKnyTfIVXv+/dJxSeaMTZkeaQja44xxbElzL6UYUGp5k/NBO/qZXhYJF
AQQfUNNBoOW12e4t70NWUSYk6mINoeTGBwBVRPUHU6W1CdoVd8s84yNsWNMD
XydhFuEDcndftdofOuzRZgW3VVH1yFIIgAxgZu3CucoWsordfEYmRFQY6dRK
0HTScluD60i6t1UO9r0RVuFDhJKYt7fWfmx45qytmVFruQWpLFtm+6WQMMP+
K7TePf8mTxnvsdhNPqMa2sTn4/SMrISBXHEKm0Zx9EIxFhr5d8+0NAVJBJ+8
5e//Vz3vXUh5+ZAumRkZcxq1OWvLdPryVFKgCcQ5vztWSznNTPOsT/iAbFM7
7+4neIZpt6IHb8LetdPrPJvsrZNnqdlMd7dAyWTjzAMQ0ZzczDKsn1NiW5y+
fTvVuOjt1FmcHP2jIkdWREQyMvt0NKhb2haPWc4a1XPUH/0j4Y1SF+CoP2Qw
zkUpiDnAcIGUQ/6gnqwZqf+irPWU0js264Z0jf+sYde3wD9CIYx4+PXnn9SL
XCGU3JHskgEjnRjSHTYSBgZHcoRd0ftCHJqVssQkT67+rEtShpTNKhT8ST5i
BnIU7nQ6KJ8EvUkeJXuMgRFRjCQx54dVKNeU+1XySsm6mrbfk5l+bYYtMKGH
mTvbvzBXcvmfb/4BNTTrjYkKKprKC492iEHbCtdoLJnyREwaw3KQfZp28Lkw
ybUrCjI8yB9fwPwI0XDkOsVescmc6JgXYAd2wJzWVcvLcqKfqs78Ew+GArhW
faHDl81C8nfDEjO0Tf2bqgSYWk/VBy+9rZKW1ES7ffysYvHGSZW+LazPlMSM
N+nvi9T402wV49YHrgi9xum5pjznIAPhnYfA+F901Dq7MVzAibIar71XF826
JTFZCxzzOPaxuO/XK31g+xpdKqWEthvHH1P7INA5Jv8oQQ74cJQJIPK095kR
3ptO0xLd/aglLx3sp0oTGGFhmycqUVSkt15dc3zGRCcyhdTgeEbpSifABTgN
9tRWHLo3AjRlHDOJlyhbJEVHP0vCfOESyh/+Fzq1EH1O2ONl4WR2XZtKgYHd
AVIXy4gHlTMYweUxEDyAh5XtNOxWpByG1+rcLzm4SuGbHdz7vsz7RYpmzS16
uVzb6pXwpvofBd1UlKtqdTAU119H1/b7mXU66Y8sMMwl6/ZfgTKVZwHk6xlG
qPB9cxdx0VQs1JcHYlfmghbAd33mwH2mUH7/Afgu0ABAaH1+DEjV4MMQjoRI
o5bsdCgevv3twXOxLHJQAvSruFSWJMJMJFgeVAnDcpsmpbaTbS8KcUS96Bdp
3R3Jl4NGLFcMlcSYOapsT4zBG2AmRYE/jhtT9uqxn2hSIzcXY10NkANLFQdJ
sR2dbLIBPOkr71GGgGpEeiz9ZMT1E2EVqKAOrppfKCeYMIqCyZzPMdmwzZo1
FCChpTjGz8FfNN5ICS+72IeXq/MLZgT+Ukbdy/xPYSgGswh3RO/1CeYKHGaS
vQYH5xA20JN4CBNI99DjnuYe/IpM6yY/dhF5xP7egjEG6VWPGZfm4oFN2wM8
NEpf4YWFKKHysX9YuXBv6MLNDHsrEliJ2i2cnZVig1aoUmgcVC6ZsUlg+Ia9
f72BZN75HKg7u/kq0LcYER7lxxlwY064L95v9PDB2H2TD25N3gwGfJ2laJ3r
Z6u8ojvZvC/9QNDfYudlD3WuwaPycHxEXaYw8o6HuYd049D0rCKnoNtkjh8U
kpTGPSjys7WduwAy/ULL8LniBCOFd3wixS5u96kyalTG2/ULN4VUBow/jtiy
3y9gNcw7yWVpTJN1QWfy0H6X9DAe8O9XhHYG68R+CW4HkFvUBFKBsYatmvBH
PDDVhSJc8HL+X1RIaCICyYY9fYQqA6LL/48pU8mvw1SAN5caokmruC+DsjeH
I/rdHel6p40evSukHrSudj0mSwVOpJgX3czF5B0jf/w9g03AgpzaVXMXgooq
6mn8tTxYKw1Wj0VoyJAmzcbYW5o5jo7QU7oV2qMLbev6L0QhRTSmw25RvF/V
BgHQZLLHwDYmyk4IbIs25UAGMuGdjnIn+CzPSj+gVF8Ljlkx9pZRTSe4Ma+e
POMwF+aVSEiJmCjaRMC06drQ8rYENO99kOMOGcapQ3KNKRLBLL0GThNg1gw8
B9D+j2K3rpWhAGZ6iQjfXizL48+RGTIehCfNp0AJJlvXqjZqbJz4V0AOFGJa
77EsK5w5sfU4sJyMAJfdy2+PIUkgIESAI7jg1JYJQb+8B83xyDB713kQahyU
pCvzVcvxPdOI/3RAby3ew/bBeSwrmvVe33AfVPK8I8gzGyTMT0sAL+4g7mLE
U21dBB/X7ArbeVlQyxojyu7xy6HcQrceufLEL28BTcMZwVs/GYzClPvAfh1U
ajhVLHw1PZUbbVSghEoM/JJ40XaOR1u08z4TC0SwdtKznq0yVyVDqQTpdVH0
PJtREmxsKWyRSZQhfe5GZb7Hr130u2JlIUqBbwTp949gHtRQ5LIIr/imFrkq
fEUQsDzP19w3cryluidK0LZKUYcce3Wi+UFahC6/32CKz/WAJGy4YJ8GWEhH
b6cW39VSqsyP8O7fJaBUKQM2QYJybXksYgx2w1+nXP+4Jvuuq6tOy/AfL1I7
20Fud9dcZ6IRpQX+e1lrCKI6bAsy6YL55aYkhbKpCePMajxt+69LuET7if9/
7N/SyCBInl730sSGKUYiguXwzeWfdtlCX++rejcWiCwth7LQfAYN8E3Sd9CV
rNyx03l9NlRKOhiIB2xtUBv8SodwJKUWevWz2jyvCzW04O2uypgYm8qR0gIU
guiEDoCJ75ABNliYZODcjdaMRONnVbqOOq5WZ57SA0wN2cjJeM/Rzf6RU/T9
u/AuExt7blyEvvpiANESbgWamRQXbVZBc4OBNUAIKTIlGTo1TK722PMTpqe0
VP8sSf+1mMIb8wNbcSsbKFZ4XlrbQQRmuVOo7a318KfuSArxhFgMGlgzZu5k
Msp4a6xd3HdCdBMYSE5OLWRScDvFqL9WYnKp4EEyCa5I8Mct4w7zIInF8oc7
OjMqK+wDNq0GZ9SnzL/A535loLuwc0NIBi/IbE3iSMbGRqFpj2YQp/MUP3iT
utbjj0JhRi7+IMyNgZkiXfS58eFvG8K4aPoV78vrIoFJ2elS9SsMWdvDDlfG
m2IF4ddLF7VJo5JxVOEkCS41/l2lltmfThX5/7wjOh3VIzny2/vThcp4ZozS
dBqHHpJDQTedD6YBMS0S5FAHu/dQsMSDN9nGXMNL9MTXByFwRGjtnkRhYM2i
ra+VJg/cH0krXkkmZ1naacOjq3cXhlUkud2Tf8Vhm/Sk2A5JtNAbWTQQKT+N
97VdTQNkcSQNTrIWqFaiyd9cjoXTBM/bVTo+5422mi3xjGytmFgvg7ofyTAo
gCgih8n9RO2tIiE7ED0rpCjvdBND6pYJ/YIuB5nevh37ZmaLhz9tyk3gAik/
JMGELjY7BPrKaXwoXoK4nI7/n9nueQlQc5suMzy4hZPQ9amuQR6tWfZiZPVC
A+GWs+q3FQIlmop+FuPlHOt0yPZg2mo6NR2ujGzw/T4KthGL/P/KQ9tZ1piv
9srjtstLzRyVcfb254A363V/+EnN8QoaiINQcVQOVgm9n2orjFYoIlHKhovb
b8VLTPfGOPJgb0cTHYAh05+KP3zlAx9eyYuNoM4Dj/zwdlB5iAyZJaFZ4Ps4
EMPk8GbY2Mfemq5J1Ce7NBIFp2PLF8qL2RpfB1jR2UAeVlzeshPWMMeyZcsJ
FVPUZrdbsQODJmyBanChMu72ugTJ4LlcmmkZlD0kPuqtsbvj/zUuPjBA+5Rw
mNEF4zizAgjf+TNxw+FL5q4yplgw1g839N15BKX2bz7laEXpdXorhdkVEHDr
68dcQrXKzNyCdPdqFhjyreu+qMNqUME9FZ3vwJkQneV0ndU6BnMzc4hJV5Ny
d2l8b979rUp9qQnmZJCvfXa/0o4/hrBofKzRhbw5dgpAVQsK8vF/NRtqc14j
9qruau3/JRNVn9ciRyXP8v8IiLj4QrLSdRasc+k5qu4dSRulVFZ46pRfkPI6
u8NLrAF0tqsBoo/j88iuzKQ29e1M3jnuxn3/uJSAT6nnN7CAuNGF1D6rqazV
ngDn0AQk16h6VLCe+o5xl+eOz0lrL5J1BPs2CDueknj9GuyFYnjOAJgnBiIf
+H3+AYDr1vLmzZhD7hb+0LFDmhiYDPzeh0mbqmWUhRt5z3kGWJwJnYqkUINr
GdkzykrPIoSoxpZPm/GNFQ50WJt5iEKGuJ3RoBSNYQrdznaejJ+U9c5pXwBV
pZ9UidlyeE+eAXNPHhYFDIDgxvsw8dEu7jBwhBpge3aJ6IdECV6wDsFKY54N
qZzvzINB6Ifsf/ADzua+VonQDp2SMuKAqwX53YDK3JWhV2SVnLPAqIjcfwu8
23fTrqvbmyKUpcWHeFG42Nu7nMAbP5YzviuFIaelJndtkWxTQXtFH+SNsgHT
rSG0r8s9rfdhjiWMO7/3T72RdprT1cu8GM53L7GT+Hog0sZ631hfrNHHorJn
LqpxVz4gC9TunbjvN7Iv1VOTKkXxYgfseKkHIzhf2SxtvUzR9ca05+PINGlZ
91MsHVNXU20DDz/qJHw07e1zw0GtWLMGxpS/EaPtzd2dB+79UEU9KbmLcFXW
fFDz9ehgctSRXNWsTvmbwSP5MjJJ7cXHCgmoxLeOPDdX8hvyAaLE5FS/1taK
oSGpEwKFT2dNgMdhgJKqOQEyABBxoV2fBy/6XZFtggwj1BFLst8KWng3navg
ChQgcGtSOqYrchieDXHRNiLO9+crvjLpHhxtvucLxHzpc5Jwc1cfOD0NrwtA
uj6vagIxQjS/TVDoYZ55UlH5KUYD+bq/WSaVkTT9pZpx1/Ryr7xuYY7ZfM8n
Q96dybAezRqqSoIQ6aBHBooeaTqDMhK9eD+EsvzkFmIMmu6M29DAZfmfxtUz
Fo8l1734aJxCdi0KQVXRfRW1Oj3mDIpDesQsPJmWsfnHvdH3AmjYFRolxZns
V6AErA5Da+1CLnS9NZSJVUG5niAbE0hk1QLylUFdWj0egCXNemyTLx8+lcbM
cWkrkpju2Y0fFJmzCFgjz+duRhRM+A25wkP/XJvXCKarQbZxyiz3S6zrHT7T
2g2f2mhoE5Tz84zfC35xYT8n1aU5x1vT7Dfa8e4DMjtdFsUSrq64pd9yJbv0
9ISYQHlAKV+0s/wZ5duXXOE9rsGZewufjs8aULGSJ1yrM/5QUjLL+3soZjqf
Fvl7p2dShwIfEdAoiRidYXFMMk+wVC1uD7TV8QiT5b2XzaEyLdKQDayYuF6N
d8LbD5Hjl5mL5FRCus2cb402ybSir/eIBmGx8SO9aGS/bdL1BCsrutVdwnYg
q/tMlCgoiF0hWTzlcAIT2+3v/UcgWXWOdjneVJbT+TkRc97EBTB+9k8Ydk79
ZwH11KdpwDbKP/w5ZKjqMCs36TPzK0X0qWiSWMJ3azw7WU2oeMBWnJ+99Uz0
8gKgc9gFgDpKCqzKZYRFum6YVH7ht1DLdK2fj9HHhaLZEWcZe4OtQKCBdK5m
z/pVkyLrLMYBH53drDrSnkbUDtU5xlaptY8xbn9fqUxbS70pW4QiGQz8xTIH
P952RaFOEz6/34XELQVoZisaoLCPf/HfFisuD9lVtloYp1jlSSG6ksw/GwNk
nZTUMUDBsvUYz86GyyX+wYIwNombCEWYdDbKndZE6m2ZNGV//jD4/TSgbMDv
tPGDgQrkyYRDXXy5V5lfM6JDN+RYii/Hm26FFCtLzJVoLiLBLKT6fljy0ttX
HrKpIyTGxiGXqTEvplN+ZPdFYNXBz9RmU76Eeju0lRunlZ1ZCENFsgEmAJmy
ZezVGytyDB7tMB3bpSsli+LXUz9WfIRooBY5X3sxmhlqYDE2tVMWhpq3ZB7z
BMyLlfs19GlkgH7ppI0IK04ILbM5vbEyhvbWMxb7QhZjXVsFC7BN4u0Vk34d
eRA3W7z+S1KCcXLF4sU3o1/sdZ31+FaLStTy43+UJU33Dx1NQ4ENUfHT+9or
YBE4VGmwMROEEI6BXAxT/Jh6OLGXOAMeOb61qP4C/pivM+g3quQJkfjsU/Jl
q2LOwBH2sNgh4GMvUQ0dg4vFWNm0fX/Fv1EtNi8nCUPc+quusDgrrC29ccWU
fvTeMemSFjxDNpcf7DXwkTSgUdz2KSkHI03LvmENMkaQ0LbW+bFh9mPlIg5t
uOZx9jHmPfoL39HEgr95d6OvPdZKQYiZ+OtJB1jc2HnGnZ1ziSdNavtAoYau
zCb2FvJSAp14RZ5BXzjHXDkDYhy25WxL8yGQSG0Wtnry88/i97Ew5XISJEYX
mmlYALnA29oolun6Jf0dD5coGgKA0lfoDonJekv0s/iJMNp7TOFSk12Opp2n
2DMB6Z+3lIpwxAot22ft3254e0uLN81n6BM560L4cvG6iTaweFXHBzJgWblX
1+ZJ+xfKsZzH3YC1qzKU6Jf00ZRnn7Gjoc9IYyqQyPvcj7xiVSl+qbFr0W+Y
hxBBnHSl26K1zYdiOvbOVsug6R8O2QwaKlVIwlk4wLo1hhqBHhn6K45fS1ui
mmxmIo05tqGjlXtLOSR5o/JCrhCQ2zq3vFQOcvV6zZTrPPwJcXb3i1LRiF+F
9/mJb4raprRG6Ps56wZBMFzl2xAs/Om1QJIGJvhw+dkv5HVzp+JmiDoi2l0M
vskja40eWkKSr2ynts8nv4GSbq06OQcS2uClEHGC0sdHDxymgiwQEIwRTso2
rq/7tC0cv3sh4wLaVagZaNAVWq8PnGtOWV3n+9L+dnMgOr1MO4rLjIWL5G7B
n04U8hZmIrj/UKt1QzHiNbg3cr5Cgw2j8VM7hZPcXxkaK8wYj+2jeThCCWtM
TcPEHcpD+Im0A6mBRlpFPzMjKUNJIvJd2/SOXyGu5nnGb98DSXhOKf9e1BIL
QF0FcEUwHvkxWx9iWCVU873DNfRW0KbNdxCDsGOTMU98OwX88UkSxcPoqPKI
DUcPCSsD18zad3FyLy27ApAM88/r230XiPTAAW2pdrozAmvd5nJY3HNxw/L+
vjuUftLdWGv46cwYrQ+GttnBmOV/OWt8EKTs75vRfp1Bv+52eYSuNjRMt2qL
twXb/vrpLB579FDizGrnOGsqkKZ66uf4v3c+S9bXkIZzt6POtp1/JSdyLIzy
2Obj1DiFZSNITBXXdcn1CPD0sIjx5n3QSBVkQ4r3ceOst2Hi7/s/Dz1oc2rI
wsYtowjim5Z0/CBzlrQpnALDgUzqiPp7Q4CoiP7OlCyCRZzqa18VKvgXvlvF
LHXfmym9eyZ3qqVLPDK4/69Aki4e50n4D/XO0P+pSvljRh0Xd/cLZUEIqIqB
WTPqzlO1/ioLHMtuxUJITl4B36pJi2icc/BHGhWYmA9s2lMKcksoHvFGn5f/
oAOtgY6J7wyGLYfFltqZwaBqtxHzw5EVXRy30ZSB2+V3XxeUQ1naWl27N1Ol
GXGHlbU30M/YAhK4/qsLAtTfFXonSaQpxOi57EhccUgUBLlaur1V6Uk2mh/C
cqGq6+6OSkIhGJzQQ5+3uk5sDDxianfOUlN4XdkulYagH07CYiKfjxJaDcy2
NeNBNyPc3sdmnFmnttlNDVGg3k6+jX08K3vPKbgv0DzYyYCZRkjiWvh0Nxlu
33YhM/tBlMEMyNbEAzJnQebgsbfBgQ2zXGkoxGAfc51zt/L9XSvd612uB2Jr
Zu+aLo0xno76vfe702CSVFxOICUHZd96ZUf8OwQtgiCrlwJUUVm6lyDnQdBw
cRiT+5pPtHZmx9bTTSIxR9RshgstRzp5CEitrjfYzyqzXKPmcPY6Rs0ACvCV
9LKGhkVYy5oHACD7AtMl3vsHKy8zwJEhtPHud2WuSNs9LIpTKeS8mSCXZqfm
Y7zm6ZwkrbFq9fpzcCOr4amof/kb088qOdoIymQyne8ZLH4lDNY1g/X27DWW
M73EA6Zm1MSf1iU9kY0fOyrRqapWavoAVIvIk047rO2KFHks9z4vTKyjvNGV
BFG0HLc50qXn9dnn0DVULCfPnl7ojx2STQwDAO/qlllwwfjw7wVZEBAk0XUn
7szesxeTbmJXY12zTIJyvl7+1pMYBSJEUrWnuXy/EhMobFMbup0r8AJinzk+
0NDlBg2nKMEud4BnzJOxYMvli4ioA+hKTwFHs+X7A2oBTEehF7V8gUh8mGPv
3D1t0tE3yimUc14GXMrI3J1Rfb4AS8j4thzR9mHMB/NNlstFHSluADt7zPSk
CDas5O7hb7RqL9vpAVxOSAwmjaG/MY3SNpUMDtuPCywwf7LdmnDkod+prKLG
8GZLvVInHfVEBCbmOYNpesclwaSHZXGpUAfJlnsAc4TOndMRtKwx4KPCQyw3
+oLTO0LpmNiP5qRhojuGNtsbthHI3PUWb0w3pi5s2/X2XPJMBWcNLzlNDuWY
qX2S0kFKYZqiY6mx3UIl2GeNJ0iikxSgP1oTL9rIsseF5eB4SA8oqRImuf/T
DboMZGBPeqDoL/ANbVpFvjL7V5CDjyGJiIHR3K0apo0h0Q2IjDYsY7oit/lv
sWuMo2WEfilA7PTIEX0tX9ajYojFjKJkR87riXBPQgcd0jWYftMtnG8JzFQu
OR3bILWGV+dwL2jSyEbFTganHPIOE2yizSZGVAv8oh+bgMuzhV6t7If090dI
CypglrfjEuy8TOYtaj3CmDlavPFZLiLCzY7cVu7qSIbk8N8mySXNpAGiM8Lx
pt1lC5n53e652FovD4p8JDUD50GVhDDSJMRS841i4uEgxkfkjAB3HQR9ejNt
vdgm+0is2qj4FoHP3mMgvViBk2lLDZ3UQX0EBcLL/ezIJnGQswrqFSON+2u6
COn+qO4joYmH0KRFCYlYQrpYzHDBIII5iCB1CPog/hy6hG1w1/maBM7Ff+1Q
WgMtjnulB9/XM9WH5Kbrpo99T1tXiMDagcD6zleb6hbdc+YkAj+YwFAhCAFJ
qftXNDgnYGwwpV4CzVn9kId4Z5Nib0R33g4vH6DMKz0XFI6uJDMIhLc7PhpQ
22TF6/b3ikVzlnMNBu2sgW9GhQmnmhJqHshgnBH8edqNyyEG0Hvn/qawj5nv
+Bl5rX30TUs0HociJw7TvplzoQcHbaA16MlR6cOT2gqBroSB2VtNpubs7c05
tbMied6zC4xkG/ApMtgiGg11dCY9qW1+kSW83xFh8fROY//69rCq5Wza451q
yQmrrHrSpbft/o1zlpnYaSNA2mKXVHfsdSb0coAmN0h7g1/VpmesN1319lsy
rR2XBxIQumrRJlzQcZNwcJCoTu3ZB6vMeGF3xPO15NvGYQTUyuegpODoVOik
qgUdBsBHaVXfl5DAEj0cLTVkeBm4p7N3F4rSrTIQmuiRUl8XmoEkkrD8coXB
R6ARM113ndJUNXDKKaobUaHZp8bckf1K3nPQMuVOlLkXHM7a8Hby6EvQzXrV
eui3GK2Ko52OjNY5Hd+mlMIeZ96ptpwLt1gRbYmX2KcpuPjd1PPeE4h8wGRk
bDsAzqFQP4YHhoHw/L4rCHTE8maWlNsxmEFB35hXXY35fer6PZVN9wrsboIF
qmmuf1hnCaK9Jqe7M7/KOx+a19AnO6wa/o2IcTCfQBIo5knOpF7EEzB7K6kz
N+CUi9HmB5xjdxwiUWs6pT9//7oUKMrV1z1jY9yCK+1fhimVBFNrvSH7iyBJ
/3eVoLKly8osb393cUxQeq3n5FywzgDWH1Yjm1m08NFsnI8XcrG2S0hGTCba
0rALN5449X+U4IIbQmLVWYEmOOw0+4RRfeqavUBbRY7Ad//8BIUm31rWLHjH
7IHyiJtz2jJyuWG+7Zbeo0V8b0wfxYSKEDVZrpUH4lW9RsDjFSiPrP7vZvp+
L8DNiFkb+MPRBm/m/qeMAeh6hkpTuTh/j2+B3FXJqXWHq41G7zvO7Hc5JXnV
piL8Xc9M5DLoh5nv6pJeWaSaYNesDWbTMx4FwnsQ3Pw8uj5VMk1EBoNJj6wP
cZtOMHjFB/9q38hdOqjyIOEEd/M4Tg1Xm0HjNax23L7o+eeksBjFc+n7aRCK
TL0ndOGwITdVHJiny+TGj8ttPlgZQCiWJiyTLnfqlX1BTkmcG3Uf2J+c55pE
p6eOH/Y5o7iGocL66Yyocxog05XOSF6iken73Ge0gBB2RP71LUlmsDAuBsBJ
IdvefVVczxehpP9QiEgWb6DNqDmV8+LjesJcB3RjKwz1eIXVfV+0KL4oatxp
xEXaDHxUiTAob5SQ1tWP7Nl7wVTdBDxhau5eAncOBqV5uHI/Aw7U/wO987O4
eQOSSGQybQGSBuefqjQrI13OovGz4IN6p12Fdbu6R7VAcn2g6vWg1PSm+vQY
1LMavhHoWKTlhUWs5ViQxaNBXzWECQ2f8UUUaRENjHrtlRW0kipJnRs/4sVT
z0qcPLlhyCZuBvFgsPnbd86o9GarZ2bdnoZfFCDnHfHPFA84oO92FHGujCk/
yo98rKnhX/U1Nu1OyQGLklMS42xW1h0aKSmoOCm3gS+l3RDb+iV3b7W7MIXE
AtYPVLX9FpRyJA7N8q4004Bc4F0heMO3o+GIkp6SanVMwVGwZIHvLMEwUqIc
qBOdsT6dkiEhcG+g3oJ17XyiL58sk0zhPgenWkONZjsffrkVjvKA2KvKfStM
90PzjFNDFKtQBunRVZ57UPjZFWVxO2QH1kBQoN77GbEvBF91jGDZSdv+Iq9O
uEgHsdPES0HUVlpn+JHti8Bm2A6uaYo80BU7Y6WE+8TjLzNLlZQwlQiQcFX4
301IrnXe2YW1eZffNnFhP0EahSgGrH0p19B8hkZP67bCwgaBebinC4EiXEcz
xyhS+TByrcikk6vZ/xvnz5BiKu0ViOsd88r7hoquB4x1XAAzpsxmsjSdufGd
8vYCzumN1bTQ1RtvOK73T+tL+gQ3pWySTZK2ZeseUxvPpmxhXQKq+FZpxj9M
u1tg0Rh8V8pxJid67xbMbkoOmnEYKxhQWkBM8mPFKkHBTUUDgiBSB7s5YaJX
u1Dg615z67w0obvqvk9azJz4twgjWttRqnCNkiRM+k1EMSKMyx/48PtfIZrN
kr+14eTyhRtE66+FmcCyUxuvysWP4F0but7makMgNGNgTmoTm+wMLFYjkEOh
54E+D5WYEEML5eo+OiKvzfEef6GC+aeqVxuT98kpIlJ2TzK26+BpdsbHeN7/
vUCrnF9pxqhKrrK5xsPhqOFyJxAjvTngokvht/UFc7l92Br2PmnvL9oJe/nZ
eTGQBXmi7F2BnwCA+GGHg01KHh0Vo1oQo7CXLxolXF6BkJLfoLHaRzJPGdmN
ngBMZ9CApM4LcwGtiF5OihK6lRP/pZnR1+xB1wZCmycTBmA/kPQGmYZuO9fv
JCdGDhR3bpykj7mKY24AjHa52kmSw2o/I8QwAFfnG8FBSWcLSozsFPxRBv2v
Ym4q2dn5fS4OBzdM42TXB19ZPKMsjXKz1VtZCnzkBNeat0EYgYzFkpiFjZPo
TGPuOtGUYn0kMoqr4CJP6X+kKRwLJZuDMU0ERnpZDpUQx15Y6+piOJMdNaIL
dISu9OCFsF+65a6a43OsNzmei1C2wntZIQxrtcDnjFLre8skDER7B4SC6u7z
wrkVl0soZpcpCAvaIfo+asqXxcMsczTJa5IE5SSlfC21YAiBFpCacuMllHJ5
u4ROtIbB+4g/JNNtkyOEFtAoheH9OMpDQII0eSuVh4depBYVLOZbdZzj9WvG
s5jx9OnC0uXtt6bJFaINQ3gKNABGA1Yu7OPo78AsJMu5zkV7aAUtta920osg
sIo8I63rvuV6d91yQa3siuqNglYLkpTTNFKgguuFh9gRwSaZgMVckF5m0F1R
iFFf9oZ2a6o4n1a8M3D3XEYpcnEIXWhSSyGv37Qz7mM7NRLBdvoH1CxhoyLc
n3+fwU4wGIyGz/Z3iSS1B9ftOHr+uiykTUDd+aadshQU3RxXWEyQZLwc2rqg
0IsmdQ+ROOzk1qsHud+6+tVdd1lGTQ1tfNm90oaLz7db1ESmmLhEEnxPmLr5
sAtI5T050ZD94eIwhRHep88LvRDJMxUY2xc/cPsFoARwnxzdTSo5fdEdmrY7
2KkkWGF6UC+dzvSrEUpUH5S7n1SLvzeP2qWzJ6UH31VTq3K2p2zTREcOLZgW
3A+LBDzxQfzUr+F7lXEtVayxHXn+w86KfJMZQjOx4D7dn9IHRp0GN8P7gdd1
7Keag/bJakswSAbUX5OSIGvsB3YBhRW7imftGgxOC7aWwqvFO6ZvB5fDc6gl
7NZTpCRnhYTZfW0SgwETycwMkWAEfXT1A68YNw/0pZslIMSmLJUPXtYN9AxH
3kGsl3jNNgeX2tqIH+BWDnUNnuNJbV8TCtgQROA0dI6xENws74byAgP3AYuS
oOKVXNEOKrkrIW0NPrMGporCbcJ8zxq72oMX0/RDeTD3Pfik7zMKe1vo7QHR
ON3S4CJnEZPbkYp20NL4Hc+7dkvYLlsOn2/1ZD4ldakEUhL2WpjkpWsE1x0N
1OPf6umQsA5VjXtDxoVqVM0DjfUYisZP5mOtPeE+6/GSrDjSxCrg9Q7DODP1
yufzvpk0PsirvEcv6BcGn19+o4SDL6YlsIpBr3qOSTDGxAUOrhFevSWh9281
sP2tixPfF6j+KW3Bu2PAHoKzQyg02ckTlf4N7PwiJ3Mm/g4RPTbsAlH+Ti5u
jM4WY1ejDwiEcjZEVn/4lnqYlB1MG60GU1WTT+iA30LHwhIbvGxiriSooiBu
zPUshxvGoJQgpZZZkLWgCchZoiLTcrgLfy8JnjjzwPCnNiC4l9vLjP9NLtWC
SVqc98r8OrWgNnB5xsdQNkGAX+MKmrOR2L7wOaL0djty3aomKy54l9WZtspS
ZuoeA9nERCxakyFXDzVYs9ri3zdw8ekv148tl2pjJ+4KGo7GMHVRaG1YeY++
IGI/eBa+4SAoffk72Xq3Oo1U+vnmMTfIj67BuzfNfOyDkuEwkxyNXJPhwspN
wOAOJIhxrOjtc0Kx8DWwPy2xZwvjALRcUihJNG4lex9CV1UfUjoBqPEYcJV0
hwbx2I61IsujzstWr/LQRodoUAKemEB6TkV+/9t0GLVG3814xu2lFQCB945G
BmyLcZJW9lJiAJPFuM6rQC6VQ0MmCCe9C1szNQKTN/V9HtsqtdZWKK4cb5Al
siJTbM+jDLgPaP2UCqiSZxjPkpYVSszJlS8rVrQBPdWV4Lq8rF+pTHZ7DXqH
RjQc7YbMQzr+3k6Srl+oIT6sZodKCUJvnrHwfKtbUeKu/kZiRlELXum7nDX2
y3vxjXyYYV1f342nkeNBMr/4iQFRaWVt8EWvZCwQKy9qRdOuxToqou9JXOjO
PKt1k7p1mk6hHnrKcqRsj0UqqGgXAaaXOLbYp301AcX9PWjzjLSGnJuRf6mt
BoyzBGBn71quDylVQ6zKysh8orMe/KJDEJbDs7fn+fhmx3shrsFhAjK683lN
Y79VkQycXOguf6PH73C9JjnQPSv8c+lypf65w40kI9F4BNd5JzsE42gSXNb/
oPz64avzpmqsSS4eAPdeYB5B0NL/cpC5CQ1LoaQQmaodLtxRUCDW8SI7ZDhU
FPcVgOe5KdLXNhGxxv9fQdSMommBDe2rtISisv8aFdV1HxuKLP5PwAmo+8En
Uw3ee0yeDY2n1ilfM/1qgxhb3g1af263XFJqHZXgcL3xYD2KAsFKeYhUKgE3
A59RyeZvcbx4WrseYRQxE06FRkMtXPI6+tdrpB+da8DqUA9b8zzreRs7RJvd
jR4ixELC5KBWWdbLL7QZSZS1b7mENkfDjwndPKKBVndy8IkNhbdaSIYgV/B6
xhXSJRprSPR75WTII4ZJp0Erf+Bkg7NCPpUeTpjsHLtUfZWqSYzdPG4N4wVL
XpGCIDmji34rpmqq0sRF6Ywxv7qgvzseXlF0pk4K0GwzXKjKC3/yAIg0t9VA
9v32Ggzw2kSPtyEdKB8+NNmpzqCVB39kFVKWyplUMzBlO/9weDIgatlhx6nq
CBVypr7MevmbXI34ylUk5Y80OSljEAUsQPCUP5kvYUm6GawYaMEMiJGU0fJy
NtyvHmxi+qs2jK2+FZPh4AZfNMrM5pJ6PYEkOT4C2A98LVyHMD6rRBu88gTG
62RngbuKoQNxCnJvSlsLVZEP8XZCt1ehUOY13ydTF7JUOPGh9wc0PmXYhpFb
pwpuBpTxJder0YzROyJArr66LH6y73IuZvL+UbfuGM9Ga0QLB+Qx6DvHo9q8
685Hh4kAe+alOC3Kwk1tZE5grjW2msG31OtrRBYov3JKWIFqTds/za8ECtIS
FPdFleSUGHtQMXL3O94ho3UwUhQiBEBepw144h6MVTEhSvjUgR3ZIkC3J2/t
RD9sGtGQV/DWXvbFUhqwE4zXHtEXnhJMk5ndaVQP4HAzFAwy6af8pwnCfAq5
sLIKnt6vHrxB4I0X8BoQffdwlb9hq0m0GyWcQcmOEE7TzrV7jtpcGOVTpBvk
IfUhlBvYoM6oKG1cvpSZ4fbbJy9rPShrgJGhuk9vpMg+gxsOpA3Ops6d8kcj
jofYBNLevpIdACWifsHTNmwXMVB8nQgngYUeGzCSGY5VDGqUTaBojs1vLuEH
0hAFScOH5bEOXsdXg02J5WGF2eD0MWPu2vXJBiOoqGzJca4Kr+4dWD0w5Stf
tNo0dXcA/gmng7dAXC+pM/AB/ShXCdNzZdK61s6Afu4L5sek4c/9BL/Z4uLD
anpUikqglz0WSX75Rwc+Ok68ijeUd4NHd+1S5awRHYmlGSiHuYAlKFnEjdHP
MyRzdxa6cxFCfE0+uoHx3+ccLI8N/CqFV13FYWC29rDv7U1ze8kxtjRuKzYx
/rn9tHTtWPPhF9RHr4Mr1aeoop8Z4RuUti6f86WWnXcjKaf6TsptfJMU6Bs2
U/kCjQgrzmI7uifPmTyu7YwnHosWQkLDgd05gqGSNwbGBrb74hIA17STsfo8
K9a5kN+1o0wTK5qIk90uD8WTFWeJFUD1cKXdEWSXpnfrHw1F63MaXUB6EVPY
7eBAJfb0Rh08eIYnsdD9suajKVh5/iTwRbwWKv/FzDiW0VAckT4VCWLhjUVd
WUGDBd2SMYEDHpAzrLDV3wZRsf01E9z6Y9MQTmoArIJ3dYGPOaaI+Ib7uiI3
GeTOToXRJ4y2TzRuD70d9sTVvf1BNO9C3JKUmwtfSt4dC5mqZ8FN8CYrvGWB
y6Yt7UPV1v+K1iiOHqIVf1gHpahxE+EIoS1W5wEXkHxWPcF8DoYtAf9PJDIk
rS+Qu0kZCzCugGItvXHq6ArKeP9HzmNxDZ6dQSMCnUY+ngIceLqUFfTz1xTe
1fJFg5RLty9g6mwWdS9cE/BIZ+em96EpOvB9k5s/6qYBllA6qxK10Y0j0C/q
JGHJoo59z3XKlu/ogeWuubrTNe84iplOgFq5mbv46TMxhNGZzn57XExDMcsF
CV102Am/Jn2FRMqttGYjLTrwBfaHvwNmQ9IgXjrz5TA1jhRplY8hV7cCnGrv
1hggjmtNupsrQhYCVK56/549S8K9p3az6HhVGmKdy7DXpe2zH3uSdd+jrgAH
vL9y1DovNDwYM3mvtDT+DCHqFcTmJgYOXT9DjNA40JyxOIbc/k8grlJ/rYII
/l51LCMrZ+VBSTzY8TuLOeAy9aDx0YOlnYcrkryU1sz1KPnZ8DKnc9WlFWzt
oL2gPug0lnD9zNJkikNhxU6+39b14dPSicr79PmXSurQ07VDfW1PwHPrny0c
2h6EM7RZ6Gl+kpC1ALxsm6hgQXM2eJA7bGTCmLbXuRB4QzzwWf00KaFyCPpN
OiWp1SfX4M6RIOpZRzFFgJm18oQYnmfXFG7yvH4cK08L2fWoAnjYCjDHh4g6
YIxjXg0z3nAUtb4oK5rh6I8rtVdCahHmmoqDE7EbU3DOMG3+xXEd1Y3MG9G6
7tX2ytVVFGC3V35LMyLePBHseIe/zzn8BESjIi4Luglx10rdrvgYDRSKfzEl
ef15x8qaqopiPjNVu1dvwC1XUHQQjneAhSNPx1HHWFVjqpS9boRbOyObCYoh
vilio6a+TLCz9dLR/zcye5bWFrN1V0yvwdFuNHSUPR9A+EG77xittzM8VRA+
mDLRjZnhqELo2eyK/h5/tt0ZN66UczdeJSiPQUgsJlF6ResyEiEosWS2oEtD
BRUuvxdLeyPNq8UTZTdteEz3h1/gXzXQymCaE+4MWPH71P4JCzbdbrqZ4Iig
FetxsFOwTFxGbDqKPhUSb3tyx4cUdn6v8L/rEc/R/M+62gFqAfY46iHWm2Kn
afi4AghPznqZM48jqUq5uNa+jIFpFdgWgsb3bn+82RxReWfNPyXYi00zyR9y
aadSSSuEZ80WOASGw0xoG7oLFX2dQPa2YndsGjxL2FkCqt43ZVDPmtFVNorm
vW20VD/47gSqQEeWHR1JFBYfJpalfolD6is8lhERctUD80lLSriJnEOx090H
WcG76wmAAkkYhUJuBh5otlj5fXmhNbVWjHuzEGjuxofvzPoarkw5H1iYXJxi
6qQv7fdGERc8bCDWUu+vi+C8mlZexmVwfFj54mCcDUuEd9/Vf0BfqmVz9+wc
SgpSIWRA3Bm/Gr3+Vgy/wg73pQuvS+uG16RlH7XV5crRmvL/kgiXh1nLPj4y
ar23sYBSDqmqAbeCoHtbNArecygdaWkDVEFL9eqdRRYbidyebE9FEB4at/Qp
CNQY50LrGUXvZ9inEo/hDkLnSt1y2ebsdcwCy2ES6vC6g86iugA/XhWk4Ie3
hn4s1zypfwOtk6+zYiBkaEQTJL1ujzRhpm74E7vpLNjgvGc1K5z6cGNWPW7q
bW+/01MpP2kLg5wcqUD3OJzEpVZKJnlbOg0IwSPW3Mv2LKgw+ml3fOcQGF10
XPTsQmjJAHbA3xg01lwnqV3G6xxphF7ufwb7ql3FO2TOAMIOM7RBNB0MbP8x
EPd9M0KGVTU/CCbbGfOjA4tSMbIchFaz2DTFFeLioL0y/PuWTNeVZ+FpA52A
BLJH1wBxfM+uG19X0h79CCAJLtIGDOdjVpx2lqHPAtF0G9TcbpYY3EyF3BU9
+MmMkk6USYVDL1ZYpYAUKQ/0/T3KzkVTisCxMsJeaYvy15y+zKmUlJNczuep
AgS0bMZDoo/5wdocNrX4jHjpyeSDQywt3A/f05GYLrnDfzBo8AQgLNCp7rzk
8x3q4oyw42bI5q2qRrez6KsWjmUjz8AC5UDEtSdoRLOF7Dp3fvY5bWrWANnB
AkD1xk+VdaqSNE+pIimEcK4IAIPd/klhJDYXyqusEs0I6L/86gkYBzAp5WPP
SyYKuLZTzJZVzvXlDkv/pSikfTtob2GGdh7bQNLUKPzJV3fDi0SbP7odSsEl
YhFcgzT1BWCPfW8JyvpAhl7kupi1LPcyQXUOKANyIhCtp+Ao8u9VuEw/mWNE
JZja4zw1kbNxzTJVjI07bAs/zW6bgVC1kJ6E8ubXU9POG0J8JHkuZlq/KYHX
ySq4AZLj1zYIWu5kK9Vlxz7Q/ZhalLi2NTFu+Lmqd/UWl81jrmWDpo/TRvrO
qySYX7WiNkmvRCx4+JfFH60EPeOxHDpGKh0W9med71b0CgU531hUBTan3ZHC
7I4pO02y34uw0vQMEIXBa0XU2NPAQ10zIWY1b9Lua48DLebqCEIDp3nInpcA
KLGh+XiRLokeGD8Wj6jCR1a/0ajRWQkd+U4V4nicTBZsRVIOLQ+J4b6Og8oN
nSXuFpGkYefDASESasOIl3zQtB10ximJRSp8LYhvdsLb0tntz/Ef90QVML+a
90XtMUiX3DZIE1UjNqXcn7lCPgxjgOYUWmSJG15WfMZC38n4YelY15o0dtT/
8hgh35OZn6mbPg+zcgErfPe2DQ3xLSP+1CeGaybn+N63sR84CZuGp2w6csc+
aDTju6xq/op5M5ndje2A4q79piQD24jhrmbbNqDx/OltXTRKrPSzltKR7jkH
O05dSu8ynzWQgW+z9mj6T0j9MC7lqwdVAy/j9Zpy+419lPB195jXStbEkL6v
bwvOnewNt+CiveI/kiKzCFyI4SYidpJi7eFsC9FMVoAkQcKFq8Cn1d6ggdd/
yF4auEKfjf4YogeP/F/Nl3Rz0LmwxkA78mNc9V2CSbNU1UpQRTh9CfAscK+o
/nQMWQ0FBQC2j/+YxYanpBQYxrL80eJgH0w1nvRG5sSt0a4xMz/T7S1ETNBB
BcNwujfw9XmeGc37sI01fCncVPG+ZKL+S26ybA7JrltEf8ilX81hQoIGL3qJ
r/wvjC3rzDiL4zNGgfNu1KwwzMnEnMRwRG2Ejp0+HxJ+se4g1ZTG49DVyejV
9IgRWcdzCxoUIartzNiv0NxQepyek17s2OQiPNxyhKmx61zMm0XJUmYNNKtH
SDuMVmqdb7F5g+xZSPPuXi92Bcis+k0bdfrKi2l2qkM2wrJCFTxfL8pY2/YD
pfd9Nnc1EElLghZ2rbHM9pX2lShnwWQmN/JhmVhbor6WV4a/2OlAHmvd9wSR
gCtKJewdZY0xYL96V/E+EGqTuA2BBI0qU2ce9OzOy2IYksY9v6Eciv5HafrX
ofJE/Ygo+kNJmS6czja0/KfB+8OKnk62WE+n/lLZ317/ypwhOmmT44z5VB4M
URCgQS6bqs/Y9cdwFbOsggwMFEGucILCump6aX2ExEbo3RrBDwutx9YPAGCM
0iSCAgiqUwZdHKdTT5gK3T6iPSbMPQCI9kAdRJzAGrxlig+sg5BpSWY9dPa6
cG54TsHiCDSJAxH6hJmrQROERx8fxm7BlJHXsdlM1AXJsHvv4uRE6oe+ScNx
ubbnnOvne+OB3o9yd1qK8AP8JymKefmrUNIlEy8o5zsVpwbe7o/T/iWiKRur
QRjYArvaPLLEaQIFtrWWCspqBBeQmRo51a3b9qrkzL2jJTwJixSn2vVjRW3j
23emtAPVNWralwLxvIqns/Oaqw0DV5oX64CX+Sguot2FeHEqtmSHLFG6p+I2
ZT2COnycFZEfkcEAYxkqhEgmn0OQIRoqniYsQcCh5vHiQA/9UsF1pEqdaitr
geKJaCbzYkBFr/QfvzTn6Z4cvO/WjOMsdUcNTceZqmpYFlghLqR9EqFu0rzp
wN/VbxDxLGQ72UimdI+f5+4ZJmr/vQlduzwK1mcq2JhnWamHUC8y9X0qc0wn
tCxToAXg9lbSb7PlwHN8Jj9FCC6zFwpbOIw7xsTBrVzbKMhsyosHOhwgVNLt
ODf6qPkPfcg5B75hlfFSU/Lba7AFuyp/4IqeYbn9hjjr5xKE+EOokJNCKTi/
WlcrYbXiWB1rvnpaSkR6Iil2Wvkr4Hv67ntbEtvL4FDRfdpyLHscvy5bKIJ4
jfw06egU02aZR6c06hfRpzrOykUetTh2U3nGXz6O0hLyvCGSWMps/AgWmUoI
T6MqcaXfl9CnmosS1dsaDKTOeTFm456j3HjSyOhNOAaW4XH0FN/ABAupZSuJ
joj71uYNw1zBglTmz/1ls7jytTwNb+eo1S54IA66wZ1J7vQtrEZ8xQIvnt+H
X53XmMJU2ZaD9PD6O6bYiayFcFURj5ivFIq6KCn+FCn+foGmHIKHJXq5ZsaA
tGiBNkZ5vL9ee/iC5YVKdl7Pi8vZwFfnmu1g1+oZOyscpM9fq87v+L0YFovb
BOnWdXzmuWk36ZSEgcAf7IPiLhtg3MmFL7WT0GH08u3CISmSypxxU19q026j
fWWih+wPJLKO9GzPmBJf5R6yQhLMeAeAVH9yKKAQSL066RNtrPsRusyRr9Tb
T3tHfKTOo5Wxnhw1yVxsgYeqySgTj58B52vn7M9svD3e6cp238GT1HCSoLbA
N18WkGjw0vILabvwBzhrXlYLBx96Dh4qNEOqiK2iaOMI2TX/+DsQBtVH8+er
D/Rrh/Crv+kZBweE8/SzSxA05k+JzI2E8QlSt1SMfs5PmxRs+OHPKpSpYdbF
VNxEq1y2f54EWjBs0eWNs2iRMmtP+mOpdSZKuKbPOyoGuCXvUX+TcHPB1xMs
RX+N4wVLJwCBsPOQAbV80xIXT1pBU6DtxzwSRz+WnAIs6sH8tWN+bFzPISGd
Hi6LP5Le2a0x+hIN91yCn7fHJ2fJxZKhDtB/s9w+Pwopx7/f4UyZmhWTGh8I
tOe5lF35KE+Kqm43KVx9Vd8khATugljR/XPHZ2ErDnHdxL1iwE2nbd75xmq6
KRq3CP80ihJOmMpt9EWQqJHySpROS1cTY2Ld821OmO5YKzoTuTgfJ+3NBQCh
T6OfrCHDMJZmkLI7oIRRzmOvk0snU8NhM1Ah5KOqR1z4Jh3MXlrG+xmIE4kA
PszoXxBMej723v7HZTvghfcERjod4gODOS+vHblQSQIa2WH0z36HynwoDUNP
RKb+aT7ExEBSJb0Du6aEN8qvVVlVJ2OgsbuKuskMU9FOm6QqE/a7FgGBwxLn
IipVHOhZjrXkRd7xQ77SD3tkidAezVAbK5UsPQL5svSujzqfbot2UWFPoEYe
MRBEYPWo6PUfGITXgwSOJEYJ9E4+wREH+sfChpXeCVPBN6/4K+8jLt5KiwjV
+ibpsqlDHMq//u9dYEcV0n38Cyi5uJF3ECh299fvAMdd3zj1G6k4y1VjZTdC
tcPO3Yd3/DvA4EsnLYJqKH44hkpwNATJ5ZQWfKuqhmmmksxu9TxKT1s+0QfB
7GkDEKeDm/OkIiIvQpTXVmzdOonlX8eTtidWAK20XBosBmS4hYIInTSFCigW
WLUYeNqejuJFKHdN5GiRc39efdQYzO6ewEZYy5nZZEjr3OSnXSNP5ijLJ5jL
gY+FkvGrEzv1FVoTQ9Q10Tau4KF5h1bp1SA+yfHLrgD8f0cGnklZqUdQ4x9M
d4z+nAu2wHowUYEmquCx76dLBtPcMa1LK9Yj3qZzDAGNBOSveP2IxdmPIGs2
OxxjRNk8JZxVa/YyVgt9GwmWzP5k8RtHU934TJpShn5eK1HXdi9EBchg1Cpp
kv1j0+VP+h0FVnbmjteV98mRj0mYOjGtHZ5tYunD6/SSZTQfzUZYL0asaeus
gWsNPQjWLOcUAcXbXNrTpjx3o4lDyVyRW5UqBRu2iI8Ezmpow5Id3xawmS8g
Gg+RdzuBj62ezzN2q6D1UKtXe4pHsZVWas1SrEVDvab1SsCsKFF8Wr5Ma/IY
V20PYv8uJtJu04I/02/fs1nEDfsP2po2kQZKwbGGIqYvp9uAGX+e/KN01cD3
d4+0twF4P5VDbrEJWK6dKPJZYg14BHDzDMIKsw6QbihJlyi0tdwFTXnGTJ7V
91lAwHptebb3c3Dw4EnQGmxYdOjIfiq6V0TQfNGmfwT7SWLloaqmZL3ps5IR
eMgobnOJccVvnA5DuHDLxCEF2w+K6UVBJj4YLAlztQzqvbBcdm8HlLm6zHp5
kh8gS2vNhGJ8Hi9xHPI45KbmZoMICjPnYiXKnvgUxBEXqXNiDd/9lGxYLRig
Q9ev+8egbw2YGXlZmwba65sZGMJ/MUAlYUPPNYE/nhhNdwmZkJhYBVqAAAhV
nw1NHyB4K0M282R2UJvV8lpLTX4mwr6avFkdHFY3uf56a4Ej/QJusWDS5pfp
qa1brgTe05NY/tTDxzudHP4CBHVSgOOcvxZPjZkNs6ChxZW14QuFbwej+qQZ
ikoh7nXZDltHvJaa2OTD5R3s0umVhC0qHxV3302Ckv5y9ri2Je066FjJ9/e1
HYWMiyq5EEoHSxajxTPqKxsnmygZke1HvIW4bi/vfi6k6nstZQ2twlj1T/aM
Joc30ylcxF/xoa9/+NwoeuMa76XxeIlf1Gl+uOTfImsqDNCXLKEruxBr9fWd
L8NemC8gJNIPAy7pskdVr4pqi8p93vUn92SNEM1COhC6iA83GV/+n2JfFewR
oHVIOItTBW41rmrKELMYgQaW8XwvowqeINBD43USmxMbPwh2mYvRiUTs8znx
YHjlYAx3sNBHvv0eD/JvQyvONfmqIsV9tGC3yqITa+MgAf5Uc0FcfX9cZAmQ
Z+xyyf0mPXa3xHFV+iZ8xR2KODvlLJ7V2PLVzXD887WfLRa9rihJUgxhj3/y
j51Emvyy9UdGVygVd4UNtSUoevHJsTEZX0sv9A4vWBnP2VhzfGVKZWozrYl9
sG7AN8hQY7g5lY/xf17w9yqgpYxMbTWKdEwTkCYtH1koj1ecXw0y5PWlHePW
bgSz7D6tMNbRMPDW43tSdipkR7TAikXMbci9N5BRAZ28RhhSADrZMjLc0rNY
bU5n6S8e3Sy8Xwo/9WXttat1kD+dalI6q7s+KOhm20i95Er6n4TZRwOk13t8
qN1/678zsY0ees6tCiXiQUj/N43zOtCB7OxKgWVo25NQmJu2tmka6IYhDyjD
kv44efLJJ3V+2t4a/jaDSBgkTeb/89RdcXLLxE1zXeXkyuSuMhVCz+cDlYmj
CBQOy4UStqUnAuHsIRfmG6djVSEAS7wMpgXoTZWfXbSsptpDzykY4iOIpiiF
i1kGv6eojMsKfXD4Lhklqu2Iqe1nl/tChRZx8k2/apS0ymEUxZQ1yCS8r7E4
V/QtqVPluAdW9q7qtLCwnPe2L/z1xwjdlbOGe9/TDqbp83oqAzuWCnMiJANO
Hax3FVd12vL0U5vaA+hgwTMHshWfq/3xSgZsoxpj5TjYDB5sn1nuY41zmlbl
DhFkBi7yIrkynJlqsiiS6RnbbVTTbM5/4NL8kTuQfo5PuBN+MQWpEYfyhrNb
A/WrjnmcXhjhABfpQJntbVzjiRmp26bTeyoGDbGIv2ThdP7p5y3kFPnFZWNk
JdKe3QsDB0wfwZpOWjfenh890dkpFo9SyyebdCZf3iZ2cXU2Yx79HWyAXb59
i7zD6tY0t7lyW4LIaoipnS/vudFF1CfdmWSat6Bw8ZuerCbM3gtIc5FrkI04
o8B120DioWMGV41HhOjrFwx++GxN3+ajFAAG81Z39TsiHq/LflgVO3Uu7lyD
bj8B/SWRwJF6U4AGkdmSvSIibAh5nrStZIkNz3GiRCk6fKps161zu1mEEEU/
lgum7+HW4/4wnYygHxZYGlDvQtdeKRkEnryU12ub6QaWGNqqxIR7F0DPO5Gk
SoqIdbxCFi4dLkIKRg/6Ul7Jl9czdnIcs33haFhGX4TS1gtXtYj5lCIwQiem
rKcQSWidI3m4CBFjli+4aj3qglD9b3Y7NT6B4NiWiCHelTzTTXOIRfpCHdxT
En9Sdl1Dds9NCh05DljnQUo7g6Sd1f0szcWakIeZlIxkmYGRWWITKUoOp0C7
3znsKaifsgMA9rytcOgt0UPATKWDW9QcJ2ELJlPgRbQWDK6XwTvvDrRemypd
/uOUg9xdGCfn+GkNBWi60hqrv4XOopvHu6XnTYW01+8CfR9UlWjdVz0veXt4
PvfUgf1J+vSirSDuhRexDGp8uPuBolhQuaK21vKTDESZGCv8Msn3dYzHiqmv
IKogBi8kFC/r+DattZBxY2MEHpq/3lr4N7tpTtlJKuDa7dOUANymBaLor6tZ
lIvio6Kp8L2u63SXHMmRd67OtVwO5bVwj/QfrUOcqA7bijj/NIMHTd/onwUu
IsBgA9PkdpCZa16ppzktPeYV8jWNX3Yapd1fqhm7AA4aQrZ39OwMH9ORbMIC
IBPIbNytgHpXviqFr3xUofgtvdDPSgcKSIUuykTpHvfyC6mUURR8W8VmACqo
2Nh5lCuyVYfVgLxl3A/+KbbxEYdJqeSh7WVtznvw7lB9BPdn29BPVbd436lb
rm8FmJ0/o/fHUfWaB7Gv0M0X2c0wWFZet1kEK2XVb3WNsXHEidXI7afy+nQn
usAJky9VcEafDbPF2nZE/XhrsIOKLg4c/g2ec0/3/u0h1cA1Y0ZVQ85lqPgS
ZpB+WPRFj7AcYULeI8KJtSmWYYtzccbKuPRhinKI1R8TS9TQoMnes0gbr6OE
zjJQodfAcOTv//PfKO8OQt842COjrhsAZyTDwBuhF6zFM96uilJiKRzPY1BF
BjLJT6efKCEyymAh7os3UWAOU1uNVqSlFRn0zHcm3rqkmkkp+qeaXnIzYe90
QYI4j6MulnEp2v3Al7pBHfMEYmMCcxrGggnS9TvTlraf0uLTYFrIpTX3g7BX
KlmKxx5QbjBqoqU+IT0G+Xe5d1eZCSxZ4fwIzEpLVbEDCwRdBnOQjNt6B0Bv
Y5GyzpZ8pk1THi71ORUnmH8RaOKIoDdfQwiv4K1gPZnyqZ4j9bEueXHEWb9q
GL+n6mJOHtZBADUdGwmqBY2VJp0FPSiEUT77KS6+CHLjydTrq9BNqzqTazT/
8LNk314H4NEzPkwxDAICuu5fOB4Jf3X/bxkY1dZcQGto5T7/Q4xaTMIsyztZ
ghq5ixSVDqtbDFsCvYRdZEnj0RVrXoXJh0IKP9Qw2N5Pgi2EizUXFeQQelRT
yydkbFQaaWcP+/fEOReP765aUr8N+xNuVZzVlAJvZGnopIs+y5+p5x5njQAs
IouGs9DeyTlh7ARmJX0/hvNarrvPIR+xVZjcZ73MomWNUELeCE4A38dZH8R3
v1SmvCQiA4eHjsXny2Ywq6kROBcnB0bf1b/xeXTlQE0+gzNleje6FGmDmPQU
GZkXyHEpm8CkUeRooj0WT4QCEzLbclSVs+WQae4NrVstr4lJDjSf64bxMUc8
FIs82Xk5zR64l83n4Bv//HR3LLygsMPmJiOItRHeLMsMv1gfPFbQQ7h9jETN
H9L/OZ7hKorTfhFqUh9KJbkLAZOrdEdhRKzqIVXeaIK1WICYmaN5DYmq9Gmx
dsruGydhvl/yAmUVUHmXrHDmI4jAndKTjTH/qnl/XFrqyrqSgk7QcQQ/+azt
oeg5JXGsoYiutf8ohzeIHnRhFU/r2CIqIdXz2D20ySt9t7CEqeOWSPbesxzJ
tGojvFAIE88IHj3k0Ss3sBSLcK+rrCwIpWQvxAEYYmAoFiwSMNGWh8ShL7T1
dIfPxUv5QA4SPegUJT97hUcOIAZ1zFvky3Hzr1Qke8w3cIY9sxjczsfsoZlz
5H9QO4vyCZ+OJygfxMCvP8NdQOqFT6LeQT/2XrB3yd9a1EGZVgHSM+DUwjbt
I0it3SN9R+W/OHxxf48fckdau9Sm1J/dSPGVjOvVcEKrgU0EPj7W5StK7Efk
DT9GeAtSp0mbTD7H87uFRyQkkOSmNCDgMv3ECDjuZr6m/ig9WYRXL3vczytD
CV+5ZjzI8loh0LTwUpAe2xSz8aSS5Xj+Y4FVHz3QIZEribtkgBrhCewuQ6r/
6Wb73TDggDFOGaswuJoZvQAPnQNkeM+X0hlGEpShnf1BK1Wje5v6BT2i/tl/
08EjRKGPNf0xj288JBWdSJj5ZaNLbDQ20ROU1rBd6QefhntYUk2RLhlui+q3
V2eJkS8G/V4u3SQL+kJ5TySqeONxXwO3SrBz1hXvzHHPaxztBuG3gXiowzhz
8I7agmdpwPtV/mJlAz4t5VPEczwKCeI6bpQgdfJ9K/wld2d1iMX+F+NC+yMN
ZX7d2Pq46TyPKpfHgDWUTP9WccAj+yRW96Y6gBvgLcr3n3mKwLr6KNbRK9b/
ta+yaBFhscd1kKPdbJ1D+mKESbc5eGVuHs1/uF37F9Sdk8xiy8ltf0Q7mzF8
MS2Es5BicIH95fk798RAW9tXoHK/eVPFVTdYIWjHenNFbu4AUdVivU7g3WoB
SXF5DsNlqaqJWvCbv//RgIQ1BWTMWMXEZq1D3nBK1GMElesWSqCphQ6/IVfA
QF4x/oqHslKmbvDE0gDiFxjSbteYG4/Ef/QVlN0Q47qHmRaC49jJGD0vX5Za
FZk6D54It5IpFVuivUHQOnRURzAR4ILeBm8Eobvm52GJDG/Y4CiLQZA+hjtd
Xb9/16/IGHFV+A3U5nBJZHKHw8/rZuWQxA47+vPEgKVOFSR8x9diZiJIWzmB
q0RqZniF+1/XsTSe8lqLNdSFmEtXbFHWFSfhR7BwVoaDsDaHhuOOL/M81dr/
JZ0FgxEVBVkf4LmvNVk7GZt+ZgCt3zRAr/IotnN5PKj2fKYpsygPi0L5ZeoO
8UDOYKoIqSq79r54vptUlPDZnxNYRjj69ZFG7+c/JN5JA51m4Vyukf+ARNpp
zNYZs+tBKROSIIm8roa6XlqF1kIaiL3j26aZoEahH+0lzxnX+Rp1VBDQqAOF
iVKtnpronvAH5RXD6ZQ3KcoZz+0VjxbYoAwOC2w44/FEpn6+jYF2QRz2NX7E
3DbFf8eizP2KGulp5QToe2PRCGhSicchu0XV3XbcKeSbl8DFk3IfQTJg3Cqw
wtGdTMK2OghLdtGdJrG5qB0nDs9i/bgjrTvuQ6dvWRA7vHlWIihsUkTPyPbm
zi3zclhRtkwhAHFKu+l4SDXNnpBQCrmGUN5aJLkNdbAEEHaj5eCvOoz1P9lf
ZEfw9gSKjQj9iCkDfY5Rfw3tEvNb6LgWtgQ44Pipy6MNIxWT2QbhN5NF9u5U
JoCzxZATGO89mVX5dhIOJQ6bHKIP+dwVL/GMh9WMwGtHoufRKaX/FFOFj38X
ncYGg31N5JWJlRRwkX+DNPQg49D5RCInYBBGYgSQ1SWSTfQo+0Cr797n2zWW
bUNS7zZEEObqRHRv2TwHynJfLsOJXnENo4A5g2KDZv4j6Ike+6eSViIi50ja
MV3RVm9oOCZ56wrWrC3X03J5ctP3ZxxvFxJgW65i+7N4gOAv8Nc6VJV7LiDJ
CkdUFyd3CdDn8FOyg/mCSgJugGEy0bjxNKuJqyGqlyjuqJDfewQsA/HbBXfB
YPT6V66zjyBciQ7OWRRTwsmrzSYRHAEZsDai24Kt/+jVXE4R75p2nv4MiX26
xZCqZxr+gkhWuS9l5EhIAjmsdofJBE1M1SVlbKr9I6bZHSxaLxS5SZMCrocy
NMukaNln4qqF7RYMqV5t+VRVpwj315itINTmpv4IML6JJaXkqa8c3zr2f6k8
+qH0jX7PQE5fCYoRJjPQb7/UW9Dy5n1DsEJu/D9RauWGI7yPjdEcSO4zftzX
h5KTN8FWeguuBJJkEBFo6XkgqBhawkJSETDYZa4Y2pBtISJ01kutUPEz4w4a
99MSSJCk/D41WpnGvh+s0LDR000igYHYGtVOZLoESJ9v1Vj/Ag3c4BcWzXnJ
hTXKCJpksEU6U+c2cqYbH9pvjtyVhqXqJLNnSxp7i+nxkDdANO9fy81+AnG6
wyfO7qGMfnr2tbSejaSL/5FrK/3wK6hL/QZM+a0mK45eu8+xxQIn6HPla/tt
ElTSOTMfPVFu9jOsL2f7oQPpK+7kknk3brPrVWKLOK/J0LttZ4OBNHhkDNgF
ZrWh1cNdHQpcUnZtyBdI9RaKK9B9HbO3mgRNq+Kevf4uSVmlJGurk1iPIycn
44CAyo3PUd74uPH2xAyY+w4cGc5jmytFBhBw3dbKeLm5GiIEYhHq1JvUTWI2
qZC54vgZpb9kMChmMDidGa/GWXMHjv2mmbgXbpIBSspPQ5k8zLhRsPXI6zNU
AtNphLS1uU/ZtyvKRpbXFcboZdPUiKW0QeA3BAt21BQBxzQ/wGm4wMpmX1Ew
rJlA1f+t5ONoEavYcnNLAtmoJD9kRQsri6cvNc2K0/ScZQwLdAiLI4w0XkwR
dk4YYiObeTg+lg2D9vo3Z3z+Qqw3mSs9LqQI1s7J5eDMlD1h7vXS/98x3lSO
X+hq/5TKQKBVlyExIsPQgVvAAw1QtsqXl7dJTzPer9e5AZPUYBtFFc4jtyWw
0jMUe23q2tfkD5unTJkET/hQIsgqnxbJncLrpot/Xmzf2jJMWtWksS9MoAs4
umt4MrwpmfudvBpJNV7BDdtEBq6qeVGzN+yBNhEQ8JWU4PDYYUMDiZrFjH8P
Ihmrs3rNA4Zo2w1/k9mdRaQdlYQUiMDKhZvVQaVjdeYVCdz1gMCXWgP3DX9u
BJ9cXhb0fMrin7YZmdFqxfKB8fBfypJQbie8R6Kojwo55bnsdMPI1kmSe3HG
50FMoukzmvs/j8WiNjWtPV2qpaS5Rk4m2/gFPDO3zebyKGkS4ECPXz7OtOh+
Gg/07jB1HEir4Bcp5cF40mgD4fW/IIl4SjcHXNolIYy3H96ZGLvQkNdw1XQ4
JF8NoG3Wn0yXJ7zdoQOKxc0ERqMOZTMbBHWY16im4kG9MnlzggF/EyWbH8nP
A0IsiQfOVysYaaiqGI1IDxpMETp3wNLDDPK4wlMF37DI8Iw3zZ1Ijg6Zn9tl
lG618pFgX3hcKPLUFnI3J1TrGfXZ3KUoVWM7asKzXane3xCBYsKJVCnMYjid
LKXvRrmnwK+7kPrq5904uA89ehr7DCPyP9nRs0HuWQVxIf3tJDWN7sHPTzPS
VdTJXa1JQWBXmjE8kocso5BBgWyQ9j/tx8Qs4sxHR0dBivTjUcwWDBzXgSJE
Xlgw8bM3Oa8aIFesg0SEvugzy4kGyojRtzYSvnzyXFmML6wqA76labBvX2rR
gjTLg1gnZZRLlZoHMcgWNVqvKz/i++VK9iSv8JG7eF1wrEO8AQzuHig+rJdX
W/buPpxlRhZtrC2eQxfuBoaTFGA+QxaIVeONQ/kL9InfQio2xzaIXMMSCP1B
RVJ8PPyCzOpaoxexnYUD5xHv0vxslOhRfkbmtzhCaBUkBFz7eSw0d9OcMQrd
vu5a36/fVVs001KuUwRp4/1Wr9wRo2UzCwtZzy911uEsmAsSp/WECb2EdZ5I
a8gGeyICKdDFleEVd6dmCmxiTdSyqZaFpVvanIUaShRp3pPhHzYVUEGU6T3b
hbMCjmtm8Rl24p2OMTsDl44JozL3Ii6BRFzMJOlPQNRqGmMm0+U/uP4rUp1s
ZOQ+x79CP6bPXOG9DrjdnZfYNyk1VAQjZ3sVcJsb+vuX5Nt2hKV8qznjrm6O
WJsPqT/0YWEIu98P11UmlIb2tZOaJK0BWaP46kgv3xWsR9ANOp8MIlFsSTCm
wK6ekdfLI53QMRjEHFh4kEnl28tlfbMMKINjWGLY8uvidFdOAJSiIp9ErS7K
hAkXBAbdiacjLm6lUQbS0sh9gM8i9TgHivoxKx1StXeNV9jFOomM5EZAxKa+
5hTQOLkH7J1Tf9BIPvnQUPEkLSfIxObR3ZI6tk35+LYvzAduhLzuKX+/j4Rm
kOohNmcKAdQjNsyuuAcm9bDdfTEiY3biA4X4M7ilDAiO8T0/YaHL4tNB6fJD
iAR9wLa2acTTPeSt8cFJYFFnPY+8JtdRSO6mDLC1cPBn5vG5Go0/ZscL5ts1
dOghBRaUn9mgZRZUtdNC+r3ISVyIjYJyOsYaf4eO77D1PxwREoMMP/4MMAt7
cAOJlJ8DrWwEW92xTxdJajt4Eoub6vmWuNnFpVTJ/bquG6t37LazSqRJqJ7X
9eMtw2S+V85iEwLP4t9EsIUE6eNnr4gtJFdl0Oz+MtPr5ZOoCFw6+DD3OplS
kbfCpJGLjj2PsuNLA7/McvPt23OrLDoxt1qK+87BXkIhmuNgT6jD8eo3sxRw
+FdTLovpaZbKY0TWMHOlIwy0YffwxytEEE6mkertD8WQATFsAYfk55LRnUli
zXXUDpoGVr52NBui3MlnDG4Ss49b4k7fN3ZCzXVWo+UxaD1lKT9WNfMfc+cg
gMSkjWHuLCW2feNFyZi+5P1dXpr8IDvCosxFK/D3FiDO2etY1kVsRk52R4kh
4zzLvvb+S0ELd7m4R8LXIW5I+ktXh62KQW6+4ZieoJPa36tCh7ppnCgu9iJo
kr1ZaWkzPG9AYU+xpA9+k7lgZ+/om892gftKVHgKBzrw5FPGfTvHkz1s2qMW
ibyW7yMTAlsgil3D/lxXS4JhmTJ9BMyfigr2PZn6swKN13iyVmlpSTMk1NPo
osZa8E0T3ZHLjTd9l8/Esp+PbDLqblg486rupgqoL7eigUQ6ErtsMnqcPMhc
S0JoWid/cT1sAeAQmhuIYDdCe+mdtgEwcDqtsUhIZT+NbUb9eo9czHcA1in5
ZPbgGClytdcT6EZexfWz7hAVLiJyIqZbGSI1yoPzHYLZCf3k/XyHiTV4UEb0
9J5l289RM5dXt29d3I0+yHG36RK6294p78iSLnUFLhfxUb2AU8Hncy218BD5
wCj7whRQVmwFOwIENRF8892eopTczIPIEfYqufO243KrhB9FSYAVVaNgdw3p
Ati4D6E9mpDAoLtRCRr3bmFcbhdMLvtA8qXetmwMo4uhs2kJY+iBLJlgzqAz
RwgCat9dQMKLDCFLspmkfSz9rB8mqceJA8T09i7x0mMneV3Z5rI46F4Hzg5D
KCLnFQCuda2RkAWSnuFzmw30iq6IFRTFMp4oHyHZBiabKrPRqsKVGRAyH56N
sdTSEosWV+QV+iQQF0Ho/J3vJS9+FtWwiLlLusmF4F066xVnBrXPigKKIouZ
Z2HenzfxqcHDrPxS8AoYOXIa15wCi1Q4arVRHJ3TExGCWnH73TvaoiNBYAi2
0pZDD+h2fMvyAhm6rM4ZlqHyVx0AtIuCsFxrBXJk7XazAb2/uwOYpEKCVxlb
WwQ3aONlbCzHRXhVLPVaccbL9rOyN+3Y9R2BLss40k7RzSUw8xR1HPuFNx7W
QfSSAQocdD1mbwyzgCNskGxRmQPYoKayGFpij0E3sKzqaNJ52v8S0mWtB7xH
B+4q/GYKETfrorrWqI77y9FNb08+eJjobbNTD9j0CagYNFtx/pXfTP1Oofo/
9O1KoNXacNvhDXhiZuOVfk3MRQwsFHCeAMzRg5AUX6SvgKQv2D6vqvhN95DA
0uKfw9lBWNlCrTOeoebAI13Hdl5XxIzecMOyQlGFaB/MNoTdfqN3024c/n6Y
cXiREiIMJ5kOdHG8oRtuk+3b0rHYIvXT0Omk14jzKaBiDh1ft4zcL2UC/5H6
Yw7XceknR9a6msh37yAP5Xfw/KEUmrI1jeOlMPsolrB/hyVR4S1BqTPdSIr7
7TSpL2waL46Fj/V08XVYiM98gsDHLh+Y3DFSLZDmzIKjjWPIv1KrcmRz/pbA
gvnjolMV/5Iv2NGyB8G6AU08yKSFfJVyEmkvCfOqYoW0b4W3TltmRRZXLQD2
a7YVpOzthXm0TDlQ+khAodnn/gsIbUZEpTY83IKGmg9kh+MP4DSdtMtaPImN
z0/6BTJFPayunTsgtr2iyt/bDEAlGrQeeaFwM3V/zvs3QfdN4f9SVahB9+k5
lPzpZHO5K0Nk0RehjsRH9BtPpcWoaA3POiGOeFTtrzZ/dYUV2IemaO2txIiO
Y1Vdspob3GbqlnX7TGXte8h6OA81mp/6nq5rl/V1SzUpGYpGnmm1/gr31St/
cmhnSO3lNOeCyYIMA5ZPdHBC2dEYaVija3usUtrEB6r25xg/ZbAu9ASkpe/y
H7tyFzPxQqFwSgXQoaMj75scqohOHBdy+QJ8j2KdZe1eTycQ8V7oYsx/j43W
B9WkEl1sB6NoTQSO3NziHB7/ZtBnUnuSJlcQhl5hSMiYFi7UhQdJ79gmWcJq
zF0kOKdY+YylzxJR4IdN3oFtOWZI1vpRjHyj9Cn80y08KI9kiW7EaSuu764y
/b/w3TeLBDX2j8vZSWPYyfaBkhUSLMa6lRakb7xd8KtVmLdiJpK9ZeaTep+L
PP8Zo4vUmEnqOrWj5VyqCwoTw2uNLCLIuMJtWALGd9Z7kHCS3p/Mz6ATzb29
9hy4BUXJeNki4lnlAHhkT8tWtG4xxW6ONZWsPMbWyBibKoczrKAmPDyvBLdp
Izz5Hd+Vm98yfZ/ttynw9/guTFALUfvYZIVP+VYwLbQYqsHAfo4Sr0QV9Ze8
TJIVIPHPazIeoWhYT/9laUFNZCxkdDvW66YnH3E0vbbzxFgp0dnhV+zt6Qgr
a+WyFax2fUdotNYaqTUriGIJ0lO176Bpb+/qhzuZemUaI/JJi1LI2pRDA+3G
LvCprZdMlOaYmkA0aWzK6XZpeg4qoRonnuueoxLei/wDcYiexM3MzGoUNjvl
ARr8fr/ArYEuiOg/Po1lw8cuWRjdH2Zzt75LCTM0IvCIBlFqz0jVY44cia0Z
CJP4wFWYYJYZsu9/Qqw1iQcj9rAYdHiAHPv9ZlLMOq/g7FVSKZSTx0P+0T5J
ZMszO0qnKU+u+8Wrou8YEG3aXSmz/Z9/e0ligAM3j2IxGFwPDaFecTofG92V
p4LcLBAYdot8N/fPE6LevWVfQW/Cu5oj5qnGYXynde1wRtzhHYnyN4mrPkwD
gj1NzLS+N6v2oU3Jb7nCWmiJL4noRLk50YPC0CrBWOBE3oEtKlgxKtlei8Au
c8fQ9ST5Q/OOwvr+R/aPbaTucgkKwKNmIRREAUrpqQa0qp3C5S+mMyD6jxA4
b44MMUVJ4e1iTB9278bcON9dRgPNu4kzO5BjeyjND4aAKav4E0M0qH0br5fA
GyP6OoePMCYMcul3mr/r2uq52JPRrumrQzySJid7I2MQCmj6iG1DF+K/nS2o
X2wvg6/dbOJu/pJ7gZNffflhG3kD31cMjRlrktqwCCqYCCWn1tN6HWhE8aUD
wEvjd/AtueyiV5EmC7qWnXzVweMLJru1IDrHnqCUI+JXuVTCDqmKL7yksXEz
G8JDUJhUtqI73CyXBtehLt2OTlvDngWZR0VCy0elRMqYUVZSwmcMSUZdq+NQ
t/XXdFe6cHW1sIPzxxCyI94N4vUonhJFPtIoFn9JfeQn9fAFulD6ujd/oy7S
UnZ+8D4D6qo7Pzr6qCa+H3jAywUwOzR2HWwfSmXCU1hCUcGed5EsPgIF8IBD
cOuiMGT2xuRbH6B2hi0ge4BReLNqLPbfQYsMkZQdPoUrlN7mH20dOG0Ic7XM
csVhNLlA/brbBVIJVRWSziQFfjm6bPy3k4RV3JVhieT6hoSmROaIGpi/3jKV
v6Ire2/SOOpsBVGti+/qyhPqest1HTxpwNL3KxH6OfTlgfimh4SUy/kbV7sa
Tm8wf3vi3kljso79dMxiqk/OouubrSPqbWD9sdtC1vBfIKCErcxr3cjq1Tdi
aVnBR5umwZCV11UtuCw1/+fJJ5LVxxQKgHxV6qtvupH+1TxuRlVxENeIY6ml
+BQvDO1Zt5yQuqbtHRHSDJ0t89/e4F55cbH+qGH4DpdF1mh3sZWErcat+/I2
XHV4X4bsGYo8zMwOGPTHZRM0gHB64ckHNGR2FwFh0UXXH3haVMy3o1Px3/Ka
+CkuAsXpSer8jmMuQLZsrgL5WTncia/Hh1Mx0yggh6rAqkgg7imtzwXY4AAR
iDovURcIHe2X7Xau5ABDxJ4YxNLMnE1uwkBGO8MHGDzkCZx5PZ/dXGMxqO3j
KJ17gXxP5XmeA4vKrUrayTr9Rfi3ZicTDb4INOV9IeYGXsN0Tx6YMymIj8wB
VQRaY/Gcd9GuqfKGHdQgah5IJvv/rSM2X0zIVu0A7O7avFjZ+lm76AFqZ09z
Vd69SdWtUHI4dt8WGIJixut2r2LvX823z+9ebL4QjnQi5cZMbJk1TvxklVzL
mBZqyTPsu6Z+K+aMA4OKEsNwWiJYySt2w+w/ee3LhlwcGPrkoJluLSL6nHEr
38UcYJapcv7dsUUcSzoU3DEM8PMsEJEe6/B5auMoFg1GH9Zc06e3fnxolGGB
VEs19preVW6AobyfTnwrCu6xpjTFnUN0lRp6OFmM1A2g7Q5o9JNlAAS9XJZU
j42Aw1D8rI8RcwB2hmmF2oJWOpZbsV4E6JQ4G58VTmeTkVkeuXHT2Tbyi0KS
vHi6SfpWPTGlCbHrhZQECpWDozJGTfdxD/Zwj59OyjqWpD0ab0pq7CB1sLE/
xpg9nscvasDNmLle3BS1r5XcQ0Q5i76Cc4UG9hw5E8baKYG1XKJV+rOYHCrj
E866rlNLr5n6G8eMOWFM7twZKtACzyp7H7HzPq55f3VV4+oPEPhke+r46EEe
7f6EsjE/4Y9Soe87/uv5y8rT3fCrH54/CGqaalcnbEOMrjxrzeJG0osWzhy4
6TN5O/urYCPIpZKoNkilmQ6GHzeSOH1r+L1YobLFK13wToKGPfopZC30cnjj
z0Imz+fwu2+Eld/52ttbJQ1E85xLwq+Ogu7RhZMbsdf54T9ktw/Lvcn7Le9q
qsfoinCcp+S0CiHv95uAAfln0hj56kujmuMHPrJWORqsza8ykAt1ujsJLnP5
dIquSGxUQT+/nqqLeF8QhFpBsdAsv58YPX7c+qtUn5Q90AlNHRzlJtEek9sA
Jmw2ddJxhfQL27V4vavd/7PnPRZb4ixUtm7oiQIrBp+7fbsEsD5/SBOJ46Rt
MFElaEklvsipRzquUqaWyQpgFJUKwrtD8Fgcl8+oKL+PZ0YUD83kB5QTKGCY
1lZUOkQZHPkEL6R5JRTIsNLgniZCfPjTNP5+RhfJlc8JKKtJIH7lkZ/MoXan
Lqd89J3TB1lw7f05TZsmOKkU6XHaTnznVpfu9fsGcprEPS2+K5B+I9cmnyxf
hhHELnyBXIo3a2ErHNCLbL/RjM59aU+saxheRiZMOPW4v/dFDryuedlNYupc
bUTAlAyC3RBtM1t++VIcWJAVHL1zyaxSUwxvNKvGBffDAApMPR2cc9myuzX9
M/GVfy09FXzHS6BrUOfzXtrKd9RRgzy+Wgt9G9p+azNMD9Z0EcD2cJBCwIOh
FpLM2VEoZbKBlxqRT8A5Eht/i1Lpsg2wzahX66OorclEZjnXwgqevZ2n2Lpx
5T4UL7YDUdBvnQzw6RHREklsvvSnadE/rKKcuC1XLbtQqIP9/ATJ4QJxlLlz
BC4rkwWJ/DqBVgILDuWvxQh38V+TjYylMBJg1I4x5TA6Z7s3XDLZZY6Uy3D2
S9X35UUK+4AJskQM/A81T6XHvtEfld9lbVJGmxvHty7yt8c2Za/JP2zPu/9d
kqkQLoTwe0CaZebQ/1aCQc3dptQ5LEByTaU1mWetpIXgwoovA8Iv8PJ7i1xf
EYTMvkT8DlsygZ1ktIO5uOp2Hzb5/FzCpnKWH+J9gnUM98FhSLArVNkSF2Y4
fFQvJIqlTwR/7tLQKB4ne1Q4JeSyq0fIxLvIQbt3u+psJI18ZRnCsjRLO7Od
wkvDdT+hlG0IeMf2PUIVDvIJ4GSOXsjo+Cio9Za+cx0mb6Aj0ooM9s6d0w1M
137Mf3SpH/olKyjQDJshPkd0q2Gjg7GdmCYPi2cDMjxRAdXTe9wQXl82AR1Q
3t345QBQmF3Uoi67AT7iyMDJqW3MJ5RMM9lMqGIxUf+fb0S8/MIslAgVGdMo
DlaATPoLhWSocMmKsCBwFQSzFHje/se60kKaxEC1qfXHvCFXk0OanT5Ac7ng
wjTdb6N9HlXL5rLbwINnuU9OpyUApoIXmY2ze7vfbJsbU3qtyD4UUIFmt0Fa
uxE+4WEQYXv5QzH6spJ5VX65pnWkk6KcxaHEflequhfTA07AKxT0wOLSBqxA
rFhLgtHNwzs3FoQ0eF8yRY3Wi4jgzy3WNgVGlmPLO2uMUrs9aFV6CfZcK5p0
akLgSbNg+tJi0dUNWjWaejyaFEfSPhUGQlp5Dex4m+Odoxz4riGdF04GANRm
ukI+80Mij4CsvpAIlkTGLNwFuTYA2zZg3Gs8tGInUeKRhmNUFCeHuaOmDSLI
AWCHO1p8U6Y+KuYoU/iIpZqvBxsaOsl3t5IMwTJy6tvbglrV8WmuYtLxYzPg
Z/j2wymMAR8x4Y+TTB5gEXAxv4E3+8qmiD4QZ56+LWeXm237cCTrwrSl8L4A
I6GpVIJJRxxezLDjtopVBtnd22qEMCmtt9EoOFn3x5jp3p2fqqEuJ1xLHHmQ
AYTBcqf+Now4nAiWH4SlZF2Xpgu+HAbmAGlXxnuiLaqoHplRLcoQ/RjEyz8a
lSyfNrNifQBiXW5Cn1uS8zrLAh0yDCvXAV3IGu1RnqIrS2K/zza+pZ7bVza8
hj/hIzhO9Ub1qETrr3crKrcX7jlBha8RLHw3Rezmk6rj2o+gUB17HpzikzdM
dKPO4u0AJFs4CQ0x54Tgh3xdt7UC+9EJpjmMUFGVpL00K1sHLbnCYplK5YyJ
pWSlvY+3iRmkrkuUGJfkSUxTCIdiT5bbjtrhoitkOowr4XGg78ZcPkYEvkEs
VvbSMBMVZlKce4HX5INJ8rvBEuz/yS5487CEMv8HdDXTmGVytZyF2bGi0LaX
shwvLT+6oGTKj7fupH/T9tiZxLZK2kQnWTqkfSUACtaQq2KWBC4zwkuMvvC1
Kee2UgN3v0CHLQUpBJRROgbSSaYEPjN4we70bdkoDuCgOltas94RW9WM+1f2
PxsJdctOp8WaGqNUsTYmYWj7yB8g2jslJ/e4Ss7q8m/O+0sHQ3y0DxSv/OQT
rAuaQz/buA/uw5ahJ0nrwAiOTSM0oxUuHVUST1bJLp4SrUA4Q8ASf7iFh6I6
Og/vxxy+W1Cmpg4lX2WSLe82YSXBlhknDX5S4SeN1kfqHeOyBzSg0rjT6w9R
eQ7YawCJnbe1KSyQ3UvB/5s4dOri2nEx0F5NrorIBv100TQhQ6ow4h0Yjjpn
Gwaxzyu1O988y4JXO/M9uIbAZQa5CLk5CIZdjj7klIgHGovd8K7hR9PfqZcF
noruyTtdFj88sxjQF99KbvH964Bhto+TzzTjl/XDdrQq2FOSofOqu2M4yesL
nl4T4znSAXGXo2HO9xKQWLMRZOeEILSP0BPMCtYzxZO8nMfwA9oSUxlh/dF2
EE/qYa3hVB4SEwfNjWi6bueX8uxm4EvMYDprLU7gez9WG1wXaLwzELTy618S
LSnc8e9iyUoDdbJQsu3pXvF4C47mvMRHtPc+0kYYRo0wLc2jv2sgWRXFkKbv
reSEYCBe3XfWR9A0hexTB2X8wy+ua+R07MIgz555k28PyxeqgaHLy/y0vug3
61QxmzLbpfaQODv5AAddvm60bikXzDtEFZZ+S6WKACVG1ct/90jx/6HUolKU
n6fNaZf8kXbaRkYoko3E7xVEF0UbviC9xAlsDXxyugf1a6et10mmX/lKvwQb
xzWOx7SDOg8Qnq8VKkxMVNpsgkXYeIPZ2hiT/JSpu2mJT570SHrnBX58YIHg
6J01l38Evz0gxe9hG6xOsV4AK2W5U/McAV6ifzhN42DUquFnNr2eC4cJS0Ov
wL5wbMONX+TA8fl9o3kjiZNL8EiqVcn6foj7YW+FzTxsvd8+e0cvoBcCe5J6
mwklwn6OOk31i78gCM5q/A8m6IMylhoelUSx8D4JBRJ/iThAc3521FOQs+I+
A1RRStbjuoofjFzeV928nk/1lxXhzR+LfuSsgIk7fQo+qKhIqiKC4SldjKoB
n0bKByTV+1UwDPDFsBVp1/PdXmzAEHG7q2iuFh02NX2Cxi8rRfRs7DD6WCN3
FJ9t8UcsCDW/2cNsEWu5K/0edFZmnBe16yh4bE2b7ne+t3EW/lyaHGq0ALVm
StZMUramHj3dDnVL2rYR4e4L3W9Cd21bGhrrvLKHRtlrixbKioTNKjfwc8cJ
4faokxrI5e+YUEthIDENazDjwo6XoJbmSmgafgRcYof6N7ol9tNtVCAyZQPB
6i1RCRWbxMpxeTt5oRXwQ9G7WaqY9+zNfwhCR3q4/HuNChz0/14a2SLSW7T/
J1z0Hq/kBpswONdeHmj/FvCuqRIs+0MOL3qH/6xNADLNsM17c6HhpkFgXKG+
POHKJLDhvPc+1146UsrTtXw9R3wV76Va2NpK5024DwR5hOIM4QeChq5VNBbH
vV8t7pUFqUDT40+epFshIMgLG8FP2nj6WvXgdjTtmtE6IbOV6ODM4luq3Dup
+1DB33UxVYaTd6ooteH+HGmYNZEXl4MxOaJcZa5JEleznMkYp/HuqO3PnPdH
22CY99OjxA7v+fWhl0ULtC4pT9CfraPb9j3WLv1qkKtEBL5YzUeU8et6ArK8
9OfV9t9IhKd6syWZFTUzsnm414PjwNZIWHF/B7ON8Ce6BZlWRt7hfuBtlqaJ
jUKPVQVWutQbyvAEjHSZFiNi4vGoaWzebIlCKR4Q67hgiMgixEAZcRpKc7oI
MY9nlYQyJoCnRngM/9ax3gXd98YU6MR7bmHe+OEax5cCkRE2W9k4Ukwuf653
C+QD+E6fCGKiYrxJQkpuy7ZiPRzT8ugq6qMZyEq1AZD7fGNxANory7WpZWFS
Q62pHNmMrmkJVIsPAlsvH93+4DvlBq3RPuifNtBZjh5ZGWD7sF5fb+ZFHwgr
nTTOeJCDuLPckvKZrUqh2x2/JcyLIJUqm70YVWGeGotdD2A7rO0UtnaNLhlM
o9furl/VlTnOAlpHYI+WLgLzulEKfNXdkZhaCUiolPsGDS2KSTVTd6vS5mAC
At7EDJROXPuxVzk5v050h3eW7QoIBgmLzcvSdcudSRy8K32WU/LGzoMRgJXa
X1XWwr2Lv/xD3wid7dOtKMNaxUUjmze6SM6HxLtzj9BwB4kaU0XJlsK3Vqyh
SOko6km8SmhsUMcARceGrjMMY/etJArh7cgUrvlYhLDQCTQfTXxbNEoS6tMB
IiR5rgXlHGxXMN9hNHXJcl09yXqiEB8AMmpToKDpK5I18/iUmV1sqX4gM76F
IaUwxQKG1Y8GG1UH23iFZ0ZooUqL/fs/ei83RqhBRH0QJaN7Nn9mAv6Avjmi
dsa2mk7PgfIH/8QmsEy/M9lALCrvYaMXw4BNztwWNTZ0C3prg+xpbLC3dVDj
qqnxten26vspHAaW3uTzRR2o8F3Fj+8Hw57kvFdwyepMhbHRLmnKyt7BFEkb
SsCdKE2qRDDEjLUFNsJI5Pp2EsVecFebm6TZmRfsJercewU3eZhvgIMVeY+M
UYWlsEs3hydwKc9tVDOx3FtSsQru9KTTfByHpIRU+6xl6uWKNQpN4cz4NbRV
HQdO2hwk2hLHFey1XOyxbZ6/L4+Kg36XdLx6Hka4rbuVlAcxiLL79TQo+Vbl
28nu7agtlut0Pt3yWXrExxuBkQqShUSDWyQKY99Rg/1F9sOGXdH/mH/zXrHk
1x41RytLiBTeuD9ocFcVwywqdM4B0pJhtotLWwiWQQBL9CEIqUHlRLG3C0Gu
WX438hHkLCU+oKF26jjgb7jFe3NuOLw04jqZmkMimmAPvEDl3u7ozzJgzAwj
a+HnHm/xR1jeutoecAQIEk0N1/09tK/dRxqYWKvQ6HoqsnmaSxyMSKO4ARzP
uPSLtrhMvX9nVHzzGhAMgHoUY7dANdvy+qHOWsalPoRq2DoDzTM07SmmX6RZ
yPIQiab1myXO4gSEchWmfAC7EOavtLlZwFJgpPK6arVmNuuDwrkywc/ylNVz
mhJVKPDcpanB6pySPVBy1e2uREbq9JCq11jFj3dTOcdaUdtnUg99LXRWCNu3
pnHGCBWSCmOgmX4ABRDj6qkTit7caW3kCL+jCiy1CAdmGPFwpjeVqBl9zN5I
lbYyz9hx1dvq0wwajjSJeWoKI3MUTMmPYE8vI7FgT3oeGIllBBW61T2OoAM2
kKpHducmsZdIX4CVtomw2r6dmfCtsYuAmabbDoHMp0GCUB4Qk9LP4UQ7bkUB
mm8Hc6AqCDTRxafC/bg3JYW21iOVdS3YWHxgCOQOlGrCmhCco1QiWMTYVoT/
HsIJtYzqU3bGMgvc779twMAEfFb2h+JIg7kJbS6rWdRhUX5U/hFuY/FNKIkv
LEDks7Vyt3pnWuwnVqLy9AwT8KtERynSRSQR0RZ8aKAWEtvXar3ORy+v+Jjv
ENxa2m3grgesmBWHjhIB6Q2OJVbCJ8bs5OiHDWDCLFwlB83WbHJ0p0KEYZOq
/0LsCyVPXZTVVZrU/i7nBP91vwtXdVjJjL8M+p3adKewVt9Tsa1wlUjBolJB
fImSXcUHrkxkLQwbS+HfTHkHOgn3UzZLe01jdcLv3DlK58la6braPcvIDCOa
ISNUoPOz4qIQMmrzERxaAbZ2P0QbZqujG/pnpcl78W7v6kA+moFG81M+ZKjP
Es4chUdn0ZuVrCUyoeSR3h52tuLc1Fw3N55TT7IF/RqCk5K4fp0eCado0XM6
eASG8xFE+ajQRZD8kPtkgGXBwP4Xnpp08k59XYLXep9y8EfROoVX8X36UUjj
FZbhUOmvFOR/CsYCywuxXIlyYdKuBR3w8d1xS5gz6mTbBHxOWJw0NckF5aO/
HBEm9ZvvQCnMEak9twZGSJs4La0avxbDxZuzjOPSNZ/Ive7EfzA70AMYQJgj
nA1GzHawSXREm8JIClFFsjmLB7LMW5bY9Mh6ISs6oGcn1LGu5GmPcaAHN2T0
IVqq4v/CwOkdtdoxJTsNWFayjO7p7Fww7AELOcndYEIctGsIXgUczooBxYBT
PD2EVDl8kJlretGsW5BGjOEHTs1gm6fF4/tWVj7Kcy+vKEl/ZFEEK2ZnTVyU
HgU8trs23sbAHaHu8PsMdKBDQ3nbmPmKCh2ezwI4lMVjXm21jygLes/dSZBj
WqV5hT3ORL96ya6OUr69WhUTxynBNQdd/Qrt1tUzq4q/OYgRze7gx9YaWLGL
I3VxJq7AMdUOl11F5XMnIeQ7SHfwzi3vK68clYsMuzhrP/kFqnaqCtYpd3G/
aZXV4d3ucxbJigk7DTLjaI4cBTxIz806iezSlMIR3El5Uu7+nCjSGwjoXDiw
rVD7qPMsWMcEOiVuaZ452VdPZFdkbAy3k4rhuRmnWW05JtrvrsDHauetUdaB
HSq5qsRYTmeWNTwbaKbvpDsMQuUVU2lAXDyHgJFkUQli9LLRfUgZyZY9cHDB
pZWzPjV8cwFSFOJIWxMXTI7dXCfw2IDwLzAug24a8kDrSWm0+sxnLN6C6WU2
kjysC84stGfWmGsWvlxNeArh4y3uXNCec1LMRyUj8yBgDukigZLRD7Sn7+TX
tUvxh7MX/Wa+UpliVQTCQROPl4kUtPakuzPegtQVc9qy2M2euiAFzJSeoFJB
3n5cHuKi02drZIKkjj56E7/ekp9mjD9Owzg+efehYzzhaS2fr0WvGWY8HdLB
dc/hgRnNsMr53Hk2wS0oJcJS7B1DHwcBIWPJ7x/LqA+iOYUegtwMu9/qSMgH
hydFLgf31m0+AI4LKBXd/GAMMOvm3pfbioLlIRd3saObeUyFujzgfQUCdoI2
cSaMvN9tb1gYyWNFrFzGMe5iaWCeecVIQE62WmxjxHG7KjZ7haYU0vQM95Sw
Ol2r8SqkrrKzdRMaAzRPehCd9YX/0lFtgYt1cmWzbRgonKQZyKA6974ats0L
EphoR8jxTjdsxwCx1PwXOoNovzU+Vpy0fqvA0WqBlx8L7VTOWBkoGBPc0IxT
k1kA0q0ZbqE9xgGngEQCxTvEJGOoeUB9tVbwne3Ly0G5zD4OmjvTOcrHD4gW
unZLee5fQmmQkB9z8vJhuNKaOy282uv91VEUk2FcXHaNc9BrKoEGlB8+u0cE
J651FDLwFtSTdO/MezLurATP8WHyixM64LPU7N0rX8zc+Tw/6tQMA1iFB19r
MOd7onSB67MamzrKFfl69Hi/x7WKKg1FPCAHjMUz+BrUNBW1eabRaoDa+lZ/
6EFUDBqv9eXRUcFrGQZvih6ReCv6MiJNTAzhP2+inQrGkqxKP822SwRLkJYW
s/2AqfgEmDs9YFkuQ6QoPNAV4MMs11su5vKhKo6rVTlCF+swejTOZNfG2jSc
tACjPBoXd1Z6SzKIC49J/2XXuMEQGYfGx094973lWEfFtg+4ECcXhARjteMb
9DCRr7CeRbOvuaiV8jlGIEtag3OXiIfWQHxyFuV97rD8ODc2LUPUEcmYRhLK
FyA7WmlByD+CNyv4SbNG7+w/e5uwtaDSpHXAoxIKfpNFMz+tgmYbJDzRhCxy
1m7v72Mb8LZ2Rr3q1iGHzF6b8m0h0ZPn95ZA8GYAjVOdu4+qbS2KZAWvjP/H
lHte/u4+WZMD+pzsIHAOrofin2f9Uv5Fc2JiyI6GJ9JeL4dWujmMvg9PbkWD
yXP1HWDNhfaQ0NTSpXDe0ewhBMlmH6sUohYSnJT+DIXu63ERjEkRDIV+V3Uh
Sv8jmFgQM72PH4fky0+kQYdG1ufbECLI9wNn2v37d3dHWqNEnoJzpG/nZVel
miv9aiwHkiBD6gIW2Ay7rECVsJEwUhzfRf4TAq3E7KWC+zokO5vgPxmfYA4S
hR/uhfdpf81+kH0KXP2dEiNXd+gpjbD6bfp3XvjPYeuDdAVjRvi/gPcfPRNt
OprOWR6HHaoMxFVeClDZi6zLhs+q0bx815mepOcz3DmeI97uPS4JSmf9NBso
E5hQlXP3yWeVOtzl6YPez+zM8ahmwi+4trzjIZtW1RDPWr2U1SmMpk5oCmA+
lJXnRiLieROpWE6ZxNT0xlDuY68ohY0Br1OxZIdizQAmVSbqzZO+A2b92g55
xBWK8zfn0qrov5sxE8ag1XPRgrK4XZ5OXLiKn7sxUXXgRcFYRCSPA/+3b90R
MM1wpxvmTvRhSmplJ1pHiPxlW4xtLzt6HyiMGdVti3NsPsnFtRjArA/2G0t4
gIouRCWRy7hrVI6HyG8EVjtUVUlFUiVoOL9vpHQ/HWvXBmYmONp8pLezaaWN
FBiuXNtxpiubyOdoDWdr7KwsdUzFu6745VJpAhzfTVaD+/YEUVH4L6qFpcpj
EoWLnM8VUbNvqpAc3HfGBHTEk+N7OSDPePsaGofydvXqC7G7Yl41heXwuClj
HNPz0G4JE2WrvOkCISeaQimhNbl/5KfM7+9ijbavQZZ0PvW8M/YwK2RqNnb+
mwmocj5tDdj/F89TQT4TtuGeG2tIb3NuF6GYZ9KJnf/NKncICXH3LsrNwEa2
eYlStOrBprbjhYX1Y8QNSZFATifSp26R8N5/tqEIoXoYnLa/P5uk4d+I0bTh
YAs6xjuxiFksD9pNw7tOCeJd5qfhJCzh6WCYzzJ0B406MlcuAKMQhKexqFW+
fLEcgYBnQksF2eNei8lAfUaUOL+vEgCldOUfqvI7ITIEBwz9aAseim4IyD/2
agmr7VQcd95osLUhLymUO9Fzvy2rEPc3RTmr/dXoD2MiWzqHeYU2+THy7HN8
Tz56tmf35VQroLzxJDtxWeQUDo8IAzOdgTT6r4LvgHoO0AqR39mKLGhUlv4Y
Uz5vORoq9Klx510UukHGBmmeLSbxEjLqvLYNF9WgZK+GR0KAz0fqVzUp6OPa
aX4u07oPTo0vBdiHgEu83LSGH6T3vu10VfpHsAkyR2o+w/fxiPsMreCqi5UF
2hKiNx4Liqxmy3RP9h9DQvb9yNT0y3e3BonCnX1XavwZayq+GZcS2bKPFs9k
25ulRvVVGy3c1LAXYbZ4CuKxgclz6MkykrYMjeRlun71W6SFQ5ltGHQT7Iou
jggcg9qnUH8kzAyWBfc/mK0yQdZqMZfkyCOm2xMWmWxs78Mtg5X7BzXn/3TW
K8fd/lSU/jDcesfvwTRnUzE8iWNTczdpfC5ejnNgbwrJsMFR0nygXEcUuFmG
jCEWx2fh4nxEYLIVseFl3G6534FVDswv1C7eR8BZQz+nfPP02hIK6jtUphmn
gyWM+N/5QVguNDTUu7lRt007qDjsFEFnTAQFO/GBD9IBqoREJaLGrzBrP2so
jroVYeeIVQt/cMdIHiwmn7j+e6jKZkgyInkb36n1YnX/rPAIh/+VoncPGa5l
/AJNxwBCo6pRmSDxZWkJ6nc39e9yI0TWVoL7O7dRfOL5qvMsqbMUMP7OEgge
VXBnwN8ekTdEpwDNDg7QgS1Ze/PtyX7JoxrOGvkqKJuNYU/4DTaEJ//47fla
u1g14ReDqx89nOTyJUnzd2o8PbWOL61S3DoZpTA9oYQzW7LWsC1wUFx62RKd
E3z5KtMyq67L+5VuAOrxJ2r4PmoXKO4lObzlFjU4/lxQucxPvwmZ2bBTjuIL
ebZjjRU+8tgM+C70JR3rRzX+Zmc+z+RHOcXQW1oWL31wHNQYWj5adHrIjZI3
tFuluM1fEKDVuM/9B3V0dvJED+tiG8hK3TSocoF+6vzMbZir3DJbQhf0dNXR
O1/6eP8166e04m0IYezIHFzfHzD/b+FEAh3XNZoK3M8VLgTeOh8qfSlt/BtH
Wdor8G3Mvx6iq1QZyn8woK7MYkgYjBmhqxA2L49Z4LTbbrFB4miBXb9a2zF+
tD2hm9eJTrq1YFQ6iMJseYIlm9MeLIgAX/GlYlTmG3QVwEPqNhaEtXo/zygr
6q3BNvgRxtHePWE/nQWLPqJhEFVVNpyMQmYv5OeItRcmz2zPgN/STlTwwZX/
AQybV5+C4Zx28YRGXce/lEgtoQGVpbqwBlyXIw1Gh3mt6np4eXoarxn3COLg
wjrtlrasaPfjxJamSiNdLn1pTH6aPIzZYKzHWxjFiBpGK7+vQ5vXv4SB6oHB
JMH4ILb1KVnoK2rb/95lswS/VBF4XQ1RTSlKS2FDeY/A9tvXZaVO/dF1/tN9
/9qgcZOfAWvRtz9+VaRqleILBZ20XY6pR25i7gWntv0janitOLBENzrqPhny
vkRaDedJzSgcWvzS0OV7o7PGEa1Ozwpkhqc0RY+VsWjFRogroQKmKGp6nFUA
0s4utIzuZ6nogeZQrcqwQbcxV2DmcWiI+J8CteRcQMkL88r7LaEGXqng1BSn
x6aMTlPSEShKk6k0nAceNIwk7JHHH1YknSG04mCMMGmOIYmYZ4xOjsJM4R1/
IeG07iLa0T89mLj7+32GbGcIL1cn8909Us/QhUQDur77qdleWRrqyIu1r5R5
0ft4eBXcrjUTSKIVymGwtQMoZJwmv7CU/U3Jo0Rn3+6v9AwCdLbBj4lGmh1r
juBNVavaNbl1/saGb76mROt8gUHspRLMsOK6zjL6TV2OgT1rU7nizK5JpcKV
txPsOS5SLvK39M8MrPYwfpl9g4BiUjacUhm0n1ceUjkUW/MG8tHWK3uwM+NR
QPwAZ3J4In+BGhqX1IuZ/AN+rg+MCaBX6Vs4inbn28XCwhIoheKXYswyohjq
ku0DdivUFdXph4SZqUGUY+UmAjy/LAnLpf8/grx6KgN919k+Qii8hMfBoVVt
gDOnlC53j6BMUqxoQ3aqlilN8jRQpMtUpPm2OtwA+m52AWrFeVbxOqFXWdVn
MReMJZetWz9VFTeLWUZxjP8iY5Q4T+rDR9wwoHXct2B4vl54K13WoM7dXvCy
WAGZu+HV2junfaakbdtF8JrEp5OXcQIjUnR++s81pqxPwfIk1yoVad3W3eQ4
6OlRmLWj6WLowFsI5qduTKGMhj8EQoIhQGgwbVbHtkdPrTjOB0jzWvehC5b9
F8VVQ80RihiG70pCwOgFxrCNXGQiDsBG1pS2oeBMN2srku2NJgoKtD1PkEIx
Sz3EqEha8WI0NSZxeUqEk60hI37oqWpqFUhKAAuysKAvhh8gb+pwZ7Zf8eNy
vI9rrZpDQlfGK7O2rfq0eTlFphc5uCqxYVgA3lkYeum0/Q0e0G1vbpz9O1or
xX6T17qN32saT3EANHGQHEqe5Qto3l9GmMK5F5t1FM9Jsbw61Of7CquAqfeT
qxlwa5D9Jhr3zwCXAFg+W1mpN9iZG6AA8YKTxa7Mu6E+/SbfV7ISsJf72kXO
7vk2AemCw/4Y1xajyGmy5KKk7foLVXtCgkIoc4gHxZkX48iJpHjB3wEV7BcW
bI3FGvXKGwD7Gq0/M0Bqz7mvCuomgSPXkhNEaZoe5Y0WpzrO69Y4bAGO/Afx
LnNzJi7nHAM2TnwqYRScvdhF62ux5UUmd+ruXjnafyd53ObkL3PwPGp7LzQF
3/HbZ0lPNeCLq3whec4Ixj9O0ttshLriNPnzoELYtMxqQbcDEYKnP/vd1aw0
4iSnR+LlyriXSlm9AvLYTvcoTQFwQASzjEj2FFu1/e/P2aRqq43X43FIJZPb
DqwaL2Rel+Ekx+v6YiZgTBrkIdJBQua62o98cX4OIKyA+UF27/FhOt4EBJbc
wp8peBxcWjleS2SBgHBe8eZFfDkdOlD9XT5/jc4ZStewUBRKBEqrmz92jWVm
q+ZF5CMbUj6yCyedyKDjNPjBRwrxlhh7v6PgtO6oAfe5MwZtyV5VDKsSHajo
cpetq4BgXPkR/0z+GTgf0AAbJcl7OHyPVGs6TiI7L+c1nbNE/A8xRRtvtidr
F/HXdZQxwqzZE+35Dm1MAIWoO1bWjnFcPRpN032B71DshknRCY+v8rVVgubo
1wvH7B5OOmCjemab4D5l70yf6fm4I48gYerupKvxZ9xiJpbOYbiECXJQ00f2
VUr4zjVRgW9+NSpqqhYIYAfOMiLVkJIw+e+PTnaE6+zWLRTYQrFq7QnoDxXz
xbOzwk22b29fOR1mSm9AY/cdveu1m1nbS0fyZPz8FBYfBYEOJPy93rXymXM6
6wT5q+e8P98hsiVLdGr7cYcGIJzz2gd50h6i6bT2Azj/WO8zzzMXU7UVZ1oQ
wSjr8UvNplV/dRN2dvFWSlaAUHKqI6SnEfRyQGPkESM4dPZf0eam7ivR/C4p
/Jx8Gvz6Ma8ihiXGbmiu5DI+1DP24ZRzxwBKo5M00WmzFTP1kHhiRO4dlgHJ
Jy5MTRgZRonzdspALOMQmMB+ofL5R66vlmkHI2ZwnNCdWX5KrPaOsLUjIR7n
F0USeRTQLS7ed9T1H0MMy8FU1QosJiJxif1QjfOAh+SjHQ6fmuajuxuladsk
2QXeMukHR80Pvy1CiHHzdUryzRS74hNE77X9WfU9IypBH26/+JDMglmh3mcE
R45iSG3uhu38ZUK35nrBflzPHifDS8KFxdRUP7eREatNL/DtKNlD9uQkk3GV
afYrDBOOA+BjLv+IuFV6Rgd9JHTdUmVeSfgGf2XN9GljwsbufPMu3lQ4DKLV
xCcIVyCi8XdQW6/WjnVT7ELGP1Y5Xsnohrz45t+HHbTc7nDBPCy5ZO77uBP4
u6hraTmQlVRn1RyR/08XKzzUt40+sy53+Nao2ZpLFcUrCUEg8D5gJ+Bnj5C9
/lMHUhY7Md5ISvckM2p0ytPiN/tlrPH/sQh/67MFVH+PEXqWdqAXVyh/nJT9
wlplFJBuhSjMcgPdlvBkIXiBvAONYdJG7AcekpZQKi9nyTu1T16EcHORWUtr
2AZetdRJTcl3WcN5aoHFn4F3o0hfVE33EfUEiBqMADMYeBI0mTLhIvzBW6/s
EQezEerkinz/m6045JJMTtXQoa5/e2jADDXKC+Z3SO6eVyc9PPITP9WWbkis
pEwukft5C6DEP+7dSA7W4tgTAPiw4KvQXtx+YQS7rN887iul/O6O8y7VKdgb
BrdOQJgG52kVZ/gGU1ChB9d28B0XOhWGdt2ruBVJ7ka23uo0ypeInYqrPCFt
oVSrUePXgLseu9oJTBTEcjGKeFFIfS8LQpITjVnCXOWXOM2/ajRlpNSzbVka
jdEbGIbiaONuNnXe3+Bw8th12vriCkOFJEu+ih5o+0hjdlcuylqqx2O4TAHP
cRnFf9SggrP+EYvbm28gRS9CuJ9c61rCllb9CeK/FX0jTqzY4LZjvUNCccff
YLQAgngPCDBiDwati8EDjoOxr4bAQqwBBlhHyx8o8CFjYq9IIIjlXDLA5YrS
YBd99dQ6ox33w5xW7jVVFjcxza7OjVPE1xjorgBhN4z0If2Y7Kgp1IJ3vMEJ
imOJEDl3hejxdrJ1FO8MHgrExPOUv7EqTyezufeFNECfyUjpQnLIkvuakXqG
VZ7+f2hNaVXUH8vV6Rv+c1+zl/NgyE5MWisenVfvzvZGdvtn0cQROxDWceVZ
uwkLo4LzjpPSsEcDj7QXE9lxQN/UgFBMGyCQItSL/I73dtODwmP5il4xs/d4
WePWGfcGr0d2GO0J4Iiuge31y963Cm/EGEPg5UGI6csG+jBytgocvw/tDNVb
/azSdvPQT5ZHLqr9h0xL2w1vSWQzlhMcwVpT5eIwGJLX8tLUFCc+hbQlxR16
DzGiMsjL+jBpr8mi1YuIxmc+NO13H0izGDvMzbpDgeEnZ02xgy5dnpvFZOpW
RBO2bGls4Lf9SB6aE8yOpDKImlA1AZPvaE1op/Dtg/sIk/M+Lq+mhG/oSs/t
Iaeag/0+vJZYzpKqEhI9ft55F9Js3iB6ktLz0sZ1ZfbjZoc8C/TniA7nKtwn
Yu6BJKhVOFo3V4fw/swCiFEdzBc3jw9UWQAYLB1rK1LSXELPm2s/1RvkWyKd
F7aEKTmXDNFEz/Mo6wK6iytZBYrBgNQOcL98/QZHqtGjonsIVNYe7T1Ptqys
n6D+pBhCh9f819n+WigO1b2s3rXt/Iv5OynMC29wImuwFj5ubp0ROzYMNtBi
RPxtB/L5CIqMcYpiqYQ3JArx24QYlxnLUEemb8cPmCCfnuocwR1dBY1almpr
Ho1VnxXdF/B762c7yFyMmo39d299rjm5ksiTC30CYkmO1o8NMPg2l0oX1Zzn
QqXla+4/5GUvTlVcKhUgc72UCViPhLjSsnGf1ggiSvKZz83T9dCC0sIvM0KM
rMwL/VwvIbOlaKHJfdlku8kBgqDl74Ul+vCUG45AugwWAKPkANFcFtT2hIQx
GGqSoX8eN34AD+z+bPfyeQNjGHEleGQJzl/6kfej7M3RIRwICRt4U3lOdB2K
iS27BHbTI6baYFsOVu688SGEaX2FKjUqJVi+Yc1H1IA0vBXds8hTbvNYHkk1
4fAD6khmH55VUhlsaZUpiiQcr+lm0XcQK2EiqGKiuJxUHkCNmhUYmWvAwFYy
Yj1J1Ya12aiPrJXaPuOJtsrdf0IFKhoi11lXuxdUebbXzznR3omQylkxbgPF
VhO6wgC2k52X7jVO/1Ka71MWHeUaEFibALwQa6XxMtptTo1aCW+FZgYlQ51U
+65ErhFHHbUjD8xMW989iJo2bvMoMwi0qOAWPHu3GSTutYHyHg9jhjdX7f85
yPI6ndVb89jhrBE9ZNYBRIetWC9BH5wnDJ22bfrjsL03JPj2xnV7xjizVf1H
1Kg9I9dpKEAGWeLK/y7RPdy9wYgNgFp5k5yKiM0O/AjwXLesOagKSbRTzu4h
RgbNsQWEgmsrAZSeUG+vZIdvx4TgRR+DYP51W6bmzT/pkcKPgpJLl69dFm9y
RoPCml5pP2ooj3SeRfN5hoVIeqH0CoF2cDkFqYMtAXZZ+/llh9ishgxiR5bX
lmJF/7CT0A1MsQ3ppaUraszaXtRdFWCrDsRXun2gNRkssOpO0+Jp63sbjBqZ
Cc1mq+evU+eNOTcmZKdQ9wHGWeBFs8yN7hu1WXYfuuzS/DrhEyQwhS3MopHM
LaelB0T77eStPS+EzxJ9w0whgMvkk5qyAp9dMoYHar4a/NCwsUOmZYBzTQ6L
S8GJOMtwp6CbCiwYlcoopa7/esrnZr46sW1YvzyivLg0JIO1h8x1SFYb9eev
X7+94u+oJrjfAVOt+/veAFiFl/W4JPN1twdT6+yBnV/QX/hFKmVG2pqih+r9
qt0QmjVyOHuN1llTyKxKb1tO5hRg9lCwoLGUMuZGHzEDoLbfdTJC8yxVSFtm
7OhoJpMJl5o0TqB7mUPNpVsH2ZqiTiD4hgkIGrwl3+BfLXOtgMGvnhEqMs7a
HQgUVrrn1Ks5h0YWpT64KK+oqdZH7w8Dyl2x9NXETUOE/1TJGj7Nrwb7BYgS
H/D6vRbjamB0zel/Ce1LXY9ItAJBSFpU5P6+Unrz7yqOhVzNGqCRu4M3gl5f
KYOp6u+j83Fa4bMRIkHjBakdFHIHS9oEax3NxQU41f5FKZ6MeExXKnviqiaJ
XlAj5ULJf3vxvZjpFP0ZwudPHbECvx54QISJM0a6BK8JJ9tRukmQesTDumnx
meIONioEAxcsCbcnitaDZokoPnOqo6JUhKFcWwI7zbovtcewfY2hq4ohGLSF
vTKzX0Qo3k6cUPkDadz7dGCChs+LqoTIcuoINH9VyD4cWvJFCSHx+F6x0BTD
Wf6UYrs8HkNn6zImTaI1Mmca569xdi0xZhSWyDMHQPy1r/C8qMYQBQB9pvJU
DPne0agfnaDjaAkt2i7ZfWek/RWJ+uLOINAX509vn8dMoE7TcP6WYoEdcuhy
DltlSLlqhclaJxpyqaDCGw80c4iSJVKRLL+Kdc/cf+HeJPImVPq0M9hHxZIE
JwY15zgACGMLYf0aiy6BRXm0qDALNLAotHXq6c+HW9/SUbCTkDiSOJhJHgIu
j2UbqFdpuYIpFkdHQgOh3Db8ouB/C4P+aTGp+z6dNOfJ4OcwXCTTIBcLB5dW
RApCU6psOht1cICdc9SAO5m9hh+Ww6xD0nqjrLCPL73ZJh42rBAC7+cXOLA8
Yl7BMi2oL2qFfZ/PYXxMHCrqJYkMhQnREZzNlxN1dD41awSwUPqR5VCSQieS
cNT6r2l61NpubrkRajn8tPUa5wEvyEJf8pTcy83QapDYWEIqvOhCYKfwnHvk
MJXKudvgX/aT7dKepAb0g+taDdgHAVYpIrN2mD32aTaPi81qVDnmI478wo41
VKrUEfUx0e879CS6Xe2fLhhxWZBZWT31L8dAN8fBymSXykC0An2cKJE/s1lK
iWpEe+ON6Rxlc3TC4T9zxOKs7Z5VDv24RlTs1+ek5JhRKHBRajU12+kNk7hZ
OlM6RAnJK638LGJdE8lHZp0WCO0SI4+L5wcvDgFL3UbeipwhutyusXziFg0O
cdwUy4Xd0WRFojks+8ea9z/f4KoEN9JVkUcgypHnAowwM8nIyr19BSVgmRc4
33aW8UQKQM+XAnoxvTxsN6AHqp+IJTJKv4w1t3oA1rvWHPn0yh4i5WU1CfAj
wzMnM2z9ph8FdGukbUUKT8ks+QVHRvYtyokuPZVmiwRARLd9ue0AoqXDzmJO
mMQVfW14ldR6s+1eNhd32ydqJnCUN2XZ22rYbPyw3WHALU59bAeK6J4pH23g
6N56Qh3uxnavED1BO+A8w5LdD9WyRKCqKq9NFmhbdvdS7nMySMxwxv+6R3KL
HtkNYmN1Aw1Bc/KLzC7Z7ouNhPw+GVa3dqATNPAiDhTRGY3peMdkCwhEPT4z
qTSP+NdH1fFh01BN/5WPzvfbG+puNYTo841QskM0YrvJ0KUrW9AXw6JEHNq/
baHrs8xHgMne4CKZ9CKAGThhiqvlpcLXgKx+e+hzkwRkk7IZ5nADH7GOptlQ
Jy4/VK05kcK7qQW+nJ6UjzjOjSQVLqIiOikiqPzH2jeK5FQ6f7e4EfbJdB3e
0qdP0DuNfxztR3BW4IYDfEr+BweJrsi06KuhcFfaBHHPuExFP7NGc/ixIVSt
k2CWnSPN70IDkW4lcMPTE9aWbcyP2p66zVkn60/EoO9zNEGvjndy9lNed0MU
cAN0TPqv9UP/QToIrwOXleWlG3SJ2wLdzukX++ZHA7oFbjKM8+4qiYeY4qrP
J6wdV5c8emM2tPMSQibGQIXsK2vKh3e9m6uSdiDATBQkjBBdSE14qRvX4Qoe
yGRNNjTONE3mob4va2Nra3YsTry3OfQ0cIb08fuvyyo/EoSm/nEdl6GfUa/l
m+R9VdtUQB6XV1ql6SGXIiSfrbxjM1KOd654KtRF8k6ZYsJjQJINZFJQJspK
RsIX4ZEnKOvgviWKmoRAm5f7mGW9wBSnhwewghI1R2gSRjUPxtdr72Bc38v4
4kDHGeSxNf5YyeplwM4WfochOQrvd0FbDbtheD+wn8KLJt4TjWHV6toudAYh
xEG2fMxsuaTDLMd1D+PyAoRw/ByJY5aoSgtj8rivk4Q2AkYdIoJgv5n6txAZ
euynYtyDkA2lKVic5gOjs4ULtHV9lRgvYWjmOgwMq+BSnA/JezEABe6OZJs2
vKTco+FlKmHn/pwD/kl4R5dLqeNDOT5d2iyOej9FCJ/eoJD4ygcSmCCdQhma
MyeDYBYgMbgNKz9o+J93CHs++3VpyBlpvIi9VYbEoMCK2SRwyZlxb15li4Zf
8vgaxVVtDg/kn1rwTG7ELye/oqsjCsopqVnmB997FhJspPTjmLE662/riHX1
pTU7w83iI5yfqq3oeMYkGlcA4HBK/PXjMvNE/iPsuAyVdj6cTfOLzxHte2cv
NV2YH4N43rNkr2boq2XVmQ0rACihjPAmS//XCsODKgTgmPm80DKx56RuWu7m
xIDprnWWizx5HGiAPcyHZZMwtVO1uygOcbA5G+4WNZ3KWZA21bi/+cs5lVm8
3Qu8nsjE1S2Mi/uxRTpEPHtovmWGgREyEni8Nb5z8OnGmOrtAxhKf33kjKNZ
XXBvdEY4tdEWxc/tF6sCQ2OzEU5D9byvfZsFu0Bxr/mYZlLdwxUWBu2xz3Lt
EbB+KEdSNL2iJh6xNs4ipqNz2nWR78hI6yidxMNE8ZsyB0sMosNlu2ByKQMt
JawiE/UcP3m3mwU979gDIxf18PN4TGovqFlfjrBaNEaDe44sjHfA6KtrdBbo
Tk2vHV5JveaOsOoe4AHnFXbyqj0fkrpZ98MZVWiIA/0B3yCQTTULyrDvsTn4
kfiSffez/bjRigovgbOQTGsKSRD2FxhOx597KhTQPe3DPIVDw8iGzzF+Fn7P
e7pJhqJf+/fWdny187wsOtlmkcWOyAFX4BFrlETrKc6btfsugAYfM0YIuCwF
877RYGn2JRuDIUO60UI3b03s59ajHafHv2DJHdtn2D3OJlnC5s4M6+F/meXI
7iZsanZatFlMb5Lza7CwK5xdngDiJirL+QmET7MHodszyEMN3kE2+Xv9fmpz
4PUGUMu7fSzXCzSBkPDQOZMGpOu6x2cfuqW2TuhRTuPmy6u6e8gHjoX46qSd
nsGYqVHobaQuwKEHHQE9sx3laMSdBINuCeIsNIXfxFMtwH4WlKDT9VrDcU57
O9eIU8cfqCJxs1nfE7EonVF+pJChMO5Q0DSLV75yyGp3jpmIprlXLIsiHOOa
SFZaWrPfTSJOGILG/bS/Q9+oEcGz570ymCmmoR2lx+1l0VC3zhda71ZKSrC0
1nHDHmykllKvugnDsWykAWaA4wTqmfp1a1BJL68MnpzOyb+lXRPj8ZoVN+yH
E/WtWvsr0CTy2zoy+Pybyt57XyVWzrvzjg5PauKcRGxpFzR8C7R/PhZjfwnG
aWXc0HwrkygcFVWShT8KIW/X2eugeeFtLVwZvJo+PU/dTObQHRYGPA6IPlb3
NyGe0BO/Npuv75xh6UmDFKWpzXmXjeoJaDgTiufqe5cZKV6IzYborhzOPI9X
9UTCy5znM5dFZt+EPArFw0T6C3uoIcVpjsaUM8eDb2Vb35wFZR6Mmf1nKwnQ
DzjB0FdObs5FTlp7rcdsX2iia5Lzwe+iVG3GWgtSa/SrlNb6J7jD2nocqIcQ
p6qdac34PHKdYlp8ieGBI9Qd4X3rOikuyDvmYpqEyI8SW+kcJDCbCNjdr9zQ
1X7eBl5FvOSZrOCRAGNSaqYrXC6gZZLdmNPESVLy63xmDseEFn8ISm6G/1iF
VPsC4OsgFb2/i8lWtTiuzTRf6/Gb5aQQUYpTPIC7PDBjojtkl61jDozF/yS1
bmLowrfihZYRGaKORusXKb3JUbll0M8W61uQcyCU9Z4XCld1m5gOQWmDW8Au
s9LqRaqnLM7JC7Osjyl/QtVdHyWnaWX1JmamRwhkmXrln0NPOpS0oQG1evSA
kuC8wV3Q1zoNgK5VRxilyd5muIKge5wljlm8Vt+71Xk48ONmPhiAG9ZCgDo8
XH4wiUaSlEGAMySogsjStj5rwnUuxabWSrMs2J/4EpTlGX88jnR/b9lbzr60
00Bskc8XncQpGX4VsXJVehC+CwwC9BN2InfbzCEbfivvyV7oW9Y7hRrTvPIs
MplGj80YfVyokzoI87KGvG5KaXOSEqeEdvXtWmYHbpVIjBWjBaEDc0sA4rHa
u+0NxsyOtxZHh+P6ykYpzKnGTUC8XxCx2le3CLSb+R+DFQoWrrg1kpMQhl7e
5HBtexgJ7VSMg5nPqytYOTgQMJhQOuatNX+LnpPFaE0aSUrPftJgGe/vrYBP
Q/bMHQps+NHqLJleTTvYatwSwS7TacvnJ1wUCBGD6RwXwQs8y0mqtaoloBa5
bybborx+w9Ndb+gnlul3lF0SOt5WZmRNCm8aqoMvA1trBK13xJxyEvelIkXA
9mBi+EMMk3dLnE8Yep+diaOmOer4wjhQTcWuexNWUikCyk4C/o/w8Rr+jr04
sfVuocRHCqREtNXwiH5crW5K2VDvzMdqkOpaSp19gs7B+0zOzAATdwTfepFq
q3SSXBpFaw00QE9falcA2pI5hSQQyfWPsPkH76SnzBJiqK7Fbc6OSROHANRn
7IExSE0FZKk1A9gZRg6pxTW8kdGwPkid9er5MxVd1XQjWICoPIdVivEwhc6K
hMKmibcY2Js1LlRbARbBdyNrM6mFUyMIFOeri7j/8GuvLL/Tew4HKdFkItdY
wGlzhgGoEk7WrxrIDinQt17axOxI+dVMP5kvnThTvCJ39rREFa/DOralVQcB
L6Qz1oDKY87pzQx49tffm/FqlwmBj/ucMkEbF441hcEdV9KasxMngpx8b5N3
IiObqAzTKPLAHsfys5I1APzYp1G6SRbFFdP/FvjXM6vrhD790Mmr7nIwOQGO
zOtwSpxgp033ndGDX7+Z8CkxWFOf/34gbxgF7Z5XeFWdbHxM46xhvmcK4Qq/
XBsgYq+83x3mLKT1PFhyQ//k6MW9YfMdWFCH0zBhbpBaZ/ioJ5T9qtJ1YxZN
cZ6lX7YLs6JUJWfkmUNzQU2H2+X1ZWNLhPzV4UJQxDxEbvJbDF0DXLxMrT5I
Phqv3uTL6k9cEnW7MZL2gEGdCo7/SwK9iV5xdL9b46I8tB2dgjBLLyjNL3BN
C8t0uHyGbA9gzkU3uxdwZlFRKzszAvwG/i+srhjh0qTmUoaVhvtGkglHbIvR
NrNpPTPw0Pxai8OJ4LotGVA0+miHeq6peEOaHM/ccjfs9UN+URDigpvR5YK/
NU6hTCElzH7paE34tXfqUHw5aqD3ut02ywKNu/5kxxPN7FQiGCA9iEnGRuCv
c0ZwXfSK7n9RAMYt6e08vWJ5emBCdZiB5ZNxFn9FzDqMMQkouRfXXUFzQp24
x7mvAp7Z3e/Qvcuf1756f3tepzDy+IRdHz1AujrUjsC76oTbxYeMeINOAeWR
AiIV7TlY/WrqSGtDTij42cBF4f997ezCCGmotWjDgQqeCuTk6kuwtCH4rU+Y
YIFlUAQyF1laNIb8ke7gCkRul48IIa3hYgOJnWf0l3iC89zKUkDOt6mIzgNk
GxzUC1jALbgOzgoLk+Jr9M8otUKsHY/fIsf7FcJvnsoBbZ+WtyeGiU+0VG5f
fPH3xLDg+RE0F+7/yv4nC59vhbJ/8xuRVyOd/43HqGbye61Aa71H79tHpGaw
TgXh6T3gFj91DNXPb6UUHLEsD9eRrLcUcmhHY+xvL4ll9pnmAcekrwAAo2TR
+Ataw61r5rVl2JMP1iFXyZQ9R+8Zev4mPIwma7n0m8TPCyRAKbHCMCnm4Ix6
Go9c6TPAitxi1fwscPD+dmZVJZgW3ky4MvoKg7tSDlUud9K6JVPYxIWMypyo
J5Q+qK3cW6hG+qewD8hNDGWYUpC/2sZ3wrRkCSrljQ6kGzx7c953TkoRTm18
J+3OkQyErSvbW7SVNpoiFkyVbFwDZT5XoqRhbE7FZ5idEYDgPOWlqw0bueme
h3TZ+GeEU3uckoChW294MAVtpWe/oclPq8E+1EJD3p4MNRQwPuwYyNwUjoJS
OBsnDaCvyT7v66RFLo/Oor5YhyAEf5jey+lKAB7+gR0pw0Li68yAeLxaYNeI
ZRkhTFvXIs+2wu1J4KJVmR+rH8vICNQymVDKPmwdnsZM8P6X5T1JFn5dn/IM
YVr8Yse7ZeCB4D1yPbezM6mzV2yNPDJBtJ1petL+IqndRGJfobwfAmxIp6/4
vbO+k8rHgw8TcTo+PUzcaevBekKi8UGMsfFB3lRMowpAl8zz/sQ+B8oPgpou
MkO4DvKDF/mK+SWB3Ik7OWhhgrileXf0VfB0HVCtO7QYlskPybEjkWpiM91T
Tz94rFls+zXwqm1Wy9DQ0F6wVUWpqYPy0wmPjQC5oWtxpiu+VqbicROfuXIg
W7IcYb59yRnp9hpKrafhB8uLmQW6u32uhfymvAghQ5VSUK6VtfF4nUpXA44c
Oj1fxuUqlq7ENOXY1Vx342GMskULIpin1CBjnJg8EYyrbwVtJ270YD7uZzl2
YwWtqYTdOvISx2E1zTSLsCXfzSwYs1NI6H99vU7Y4XosLmXaWF84noeBGh+D
b9cG+sS6oDuYj9i2hfwWMW4d75oWaub1hjYglVyt4BOpi8wmwhE4c+OPAcb+
ZqhzDIDcYQj9Xe4iPL2MrEurc3L12vANBQBIKQBaAwxayrisOp3xIacDwEKE
sqb7ouiFOnX3Z+/pNhPuuAYeRYgjfOKbMK/9AxRpjYWMg3kXREt0ZWJ3Z9eo
8fmnjOwSWxbl5ua3XuqzYoBNzWGvD/SYuP2BysofGUYy4GO1aEXvH42ZWaBy
rnFStpVEBp+G1I688pWMebEUOiJNPdYyI34KcnVeJUrExeiP9s/S31ASNXlR
dCroXc0xuv2IgHHPrXAPnPfNhhuQWGbQACDCuxNWHGiUn7O7ytc68LGomCvP
1DRNrTZNa715//qj3/rgx2VdzJKkGz1uozy3YucxZGUbOVMiikbtytVlvksL
I2TXzwk4dSlN06Pc2P58smuUpxS+fTqJiSbVNY0dP9g0xFv5Qti19y0fOkQa
yhU+3K7WQOVWZjmxGqsKXaiNMjvWSKlp1U7BgfW9D2QcSPTKJBhGYp9lHK12
tyyt8FAO3b7AIu/7n5k0SUOf5ZCHZDVPuv8FpQUtMRjUIXh2Us+qdS1qtWi1
STypb8jeVnvUQvwIxW78dhyFHBZXVjt0Cn4BJxmex6k+H42h/dUL2fnULSN5
jtXCeJMsAmRFKW0znLu9rDl/cseJTPcVpQPrvC13BTPfyGmf79CyIPfOA3KF
wi21bHNQqveUp/bZ02q+2qfrz0jygl8Do/syc60Engac4cceBNNrm+l9Xi9t
2JCU9C7g1ne7veWWdGY24neN6/2m08Y2kmCFOTBJQ7SParcZn1x0rJjomzdv
t3UMYJhjhxpRyakQdzveiWfdjhnChyBnyTQ89ubdD3uLtwd/5bEYU+LKI/kl
8XwBGfeivfgMS9nnsB+uH+rAw8NFismZ3b0PLoSeaI+bX+XXbtXiBOXdrIKM
ua3/p47oF0hNBm4wZMOlzAlOkuhtBRoMS7DBD/YZQn9XORzvy169vAjJ8/DT
MKHkdf1vyFwa5LcHn5PWLwmJMswtAjF0kD4OFF4A6JOiimyHVzr3YWxIGRg+
FoDX9e0Vs9kpfwEtnwCYmyodbWMcrvl662oc4/fEhxCAzylxZO1U+oglMBK3
Eh329h4lz1hNFi3ohBBqaM9OGlO4Jy8CeMi3wLeE0Oc1oGhcRjs70l8XG/bh
Zn5/4ZWyOG5jVaNnIsBNxV2o93WcIAcwlhuNkXOR12m3v18mN1jmf9RsYkrp
NSC9QxADbQ5YL1ddxhkOehjFQszr/XDrOXsldaXHyuSpKFFemVrDKe0VaKSQ
HVIjl39AO7XVtNFbJhKoX0hZXjos/NaB6ViDErzqP3cq2Gw4QhlMWSvMPcrn
PlDFl2g7qQRKqHzzsTpMv6/Rl/PyaXMXxn0Y9qiM6HogFPL3P0V9vNGe1pIg
93Bj+/dqXEZ3gIIt3rJkT7PnE1SImOydwrtqZuvNrvlEPpg1fJmphAex3gG1
tCyhpTFZ2kEp7HF51STbVujTKJax6v9Lq//mOce5HUBBoY4/MRJBWVFgqXef
KL3I9/GU15AvZNCxY6EWbFEdolOnS5U1h2+5H3I3NXHNvDhD1Y5KQo6hRM9l
oUlqvVIsVWxsVP6UnkgvF9Pi119KpqOnovg3STeYQJny29+97sRtwOv3jSHw
0gdqcFksaBfvRNQb20dGXWqmPMTyrSthu5YCYqeFXk+wUIaE2FrOmiFRnG/e
3B0L0ShrQzWL6rPRTZ2e6/gWVJfedkY4Ew1wGzJd4LNGXDdZE8TWG+gFKqnO
ICYkLu3dYbF5ulyiX+MEz++M0H0lKE4jhupjfTdbSsYGZ1yxP1dn+LAygP9n
Tk8pcHpZ8CEVMFWp6lYMTcsNEu/A84if46MVASpijScCmYf6lNdi58loP2Ny
vxIRYcIxjHKjCAuiktIUMzL6kSkrXWnvQLboNsYiqjyx8ie7ldbLEVKztaKU
bxkTJKAHheHn+Ll4lK3xoSiCUwevhcLHcs37jYIOA+05KQPODoe6ic5NzmoS
EKlAgxqIudDFQXLlXV25AEH1u3fVq7YuVQpSSTJBdbGblNg5t0eWdw6b3cP7
a6aOswaTPHjeF3GtijKqPHPbgsvsIDAENhwIYvkGKoRFqx6t0YbmGWyjNQLX
1DJaWMZx2P9YrU/KY4cu4T47H3e3KAEP5PKxkd0q6fE23uki91Sp7HT2ROqG
2VE/jPzqXt1/u/F+bGBibeEYc+eVYTyT6V7lWKFn1NltXelv7UMdOn59khuk
z9ozOasOh8m0Ene/9JGxRw1mmGFZ138dS+P2/jhLuhqO4/WJ1zLom0B+QDvY
sXCC50RGro3GtaSUtYKBK3hE7yuyLg68pyN+mIcxQNv8NvuNijHba/6k195U
IrMhgQ2Rpi3knf1yffIqbcT8P9N8+BpDBNViYlC51hr5smpdiAoezQQFZJui
APWy0V4YZiyXY7qcqVsQ7njA5G82suophySFRkTVkPNfUr7IyLhWBUvnor1o
6C2hmxbzKtMY86W7qm8nu5l+UT0TNS4e+F2DoV7aTvwDv87cu5imn5ByW5c/
pJyXOAq4+hd7if9vzZaQItpt/LnzXRoOlP0yCAvbAU78s0dzGorR9DR8Hf8p
lvVjVuUSvcEKK1Y5Z3FvxZ3Z6QjXobciyaSMaRww9YtvAoXb0YkjEBEOXfK+
b7pUTk402irvpZvmQD2jlcSW5PNQNadmSEIiRtOTq/ddtN41ItwOzNHwPkn3
3SgL4edCD8YVdlUhVJ7jw/ehdQltBvqUurLWcikHfGz2kYmBYQNk4N43WQ7s
30KmYb5UP3hPnKs37jCxxHXXBgdtK+2JV1DRbt4nt5szGemxS61BD7klV94a
pWMNvA/m06rZ8f6CmJ/tNQI0bI+9ChIjIaV7XYSJIduXywL4ZZXwBI5Xfq1X
M8JqjWxFgeoLkejVRPRxJI3KEDVKr6JGeBo+4dztto9iiUszDTIxZ9qj5sZk
w8hrZYzX++gyekZTBNIlt+DogmcdVvK33OVSTnSghQnpLilFur/0Whu65owK
6VYv3CTRKdKjK98hmm99kerYmToV9QFW3X5K95iOQSEVBAxgz9y/OfRSzWHT
L+Z21MU5NT9feYwfcAikvi7z8yYvLd5X8xkXx8EY1Ag5TnpeoU5dh7SgIrUV
TFddtgxh6xcXcjAHIdILb8zCVPbEm6s0oawMbOfP3/KkE5BaFZoxIJYqu4DZ
+87Qliw94mMMWsTG+wq9rjy2vvsQ68VvTm9P5gFLvt34cDz637Y9I/vyt49M
FjVJuLNFyrjzwf0nU4LKZ+L+Zcv53OWx4uUPNStWT/G0i/wo9HFNlv+k43PM
bNZlvFyWmWmVttyiui71CVZ+kWb0h0hrJ6Xosjgioj2SnoIh0+N0qJ1/nuCc
4IQM2bR8vH00/q21MVPmG4eBZXVvEaCxt9tcSrU7dfEA3MSDPZ4EmPciC6zY
C+L+CJBJaRavEosPFlzYrCmZnI1Bsj/746VStapeKDGKyuyAE0aK41c6UlUM
dTemuLRIDvH8SzbwFPAmPPLVjqbWF4OOJSsa55c1jsZ+UXgvZEvQABDlUdu6
2p8TfEjf5dOV9QTolVUD03t8uP1Y4+XHt5GIxhmFFu5BTbO4dG7dJPIuSSuC
4aSofIr3CGn07AzJ3ZmjkCkF3bhUEHkWvjrF9eUDW/EM3TmbC9diMx4FLh9D
isTHP7yJJp3zMWLwz2zigky/Bjx1BKUXUXsllK2DVcq3QAPKfDK0QM39O1Uz
zri/vioa1LQjrjT8Uuqilw+oI80lvLB3uBRqRbhMMKVHKaYbltGZjyMKulUx
YvFPFtcuoMbDlmYomK4Y7cPxnvq6leFmHFPb3wD+gtc0L4GnWcM8uVPiuaug
agtxG0eFwSUxdm43XMqpUobPW6hKiLAWYCRr2u9sg0SbbkUW5/ZZwjwVmdX3
3+iVZVUrGeVYWW/e1r/2a4kYCUGHmztjUVeNItaCnJijBnfsDPVb27nPR7AP
6w/ZgE5MknwmFObHrzo1DOMCn5SS0UgdUHmQfR0iUyiJpeG/PRHVNwiuBmuw
ElPgWGxm/fm8/X7J8PCrm2rxAw7WIXMzASCXSL7mv/PhhoyrSlCeYhRAQngU
XMnkxcyKZUC+m4Pw9bwOyL+8qdGf7KrpnLYOamdqaS+x1/7FBO7z8IAugIDz
3h3QoVuRUeIyeD21iNmmvIF/aFigmUnAI36qIbYICXh+84b18MWxZsuzJxwp
UKLCLsZpiQskZEK8e2AxHR/4seQ0QU7P84yYYwYmmUGmNZJI6eW5t5KiY7Md
kiNHLhA1whY2oUDFICt9nqhHnbvpJ1dhq/nuNXXIgBfIAml/r/xItgXOmstZ
O0Vqq1NvSMbjZwyXVKo9b0HtGYsG/1giWf3mpHrIxUVA9WxEpRaXdxwozswE
DojHIRH4gOY0d0gsTk0IiBuJJkPFtvUc2EZ35pM7ev/di6hOqSShHpGIk4TL
nHXpfRsp3vZ2C7glhmd0I9cWc8UrRbKZGvhmUO7aKIMIprP3zE1NUQyD9Oxe
GHvXrWCsdaZHewVmbFn97y3XFCAMJw7eiEpfLTHgauq+vHqdat+/zaUAYqn0
vIEVJuq4S+cZfCvtK9nTNcAdjT9CSsPvyer+PCqLnWGWPVQvvios2v6gux4+
brNpdpPV1bu3cKsChcj1pO3Q/PbCnKhrCwiLcig1WfWaAuXGw4d790MnJGVl
kFyxt+6yyo7feK4YwryFYebEQUphPlslPLedq75iDX8GIP4K2zO6lWHL9YzY
vUF4EbdY/USeCy9/j5TIUYcLVIS8AZGCTc9yyVS2M2BjhizyHZN4vlkZLzXG
Io0NF0jz4K/9w4pdJX/YTDluZHMzZcaE01o7UjELNVr2jJwE0u/x0n1/9ASk
1MdQA9RZNYOuuGSQr9LFOmdJ2R8WoSRA1WQA5DfALKDQ7P5GsbYQggC919xv
MH7WX5bYXfietsIDva+Mt2nxCJeyMmMDdKWd8UKtoAU4vKrwWXO2x026dK3d
mHr/xKk6Lae/Jv5XVH3afO5xalob6S/mBQwnshybbNs7isYNhKpDwVx9PDar
AR2kKEIn8XGTOno4ng82paSCt3M5QizXjEuXIuy5dAfx+Dde0Pa+ecV3KWHP
A31S/3E4cVFWmbRBWJiP/Ic1AKCKnaw+rpt6+G7FQ+RqeJglR4l5mIingx/J
ZC6n5MVe+lmXKYCGNRZ6BwHeKSs8glmv4eqTm+BiXUrey9+6nlOG1tLlvE4R
HKISlJodVsSGHgr2xPpGJYbu4hEY6QhBceN8eg0oaH5DVV0p5+gKDptCGN9L
QKnB9hlOz19WIXyiY+rtNHvrPLPJwuKTKa2q0WLWkjgusM73nZtJtEyUmS9y
UjEWsqj+thkUkTuAxQzAp5rSBI9yfTFVSyr5/WFaO7HEkWASioxZCMlZXTBh
JqW2XVjN4Rs5nTM7/J7Gh8DxY5tRv8/dFkess0sBVSYSV9eUat9WfaZTYMkN
vrhKBc2sSPLW5rgNfA3gE7pspX7yWylhcmq2uDB2FXQ6GJQLN+4aCR/ZTjJ8
8/5k/u/Ygr32gv+BsMexErJKfNzB0ekE+RAAFYniSj9haGCir8g/gYByw1Dt
KddvT/sFW6MCIwbxY5l5cUs8a1hj9V5swqdI9AcPi1AOR4IuxtizhF0Hftzb
fpNlYUr1j0ahT1tPUzlgHSjWqyfArSDe1ql+ODW/KpJoWDiWk8zUOrwjwsq/
dOeSWhumO9KY+cY+CWpzNQOP1a3Go1HrkIzcc9AtXZe3mOVoSFgvjT16Ulny
2buLpS1ujuYSUYxUQHoLEx1GGAS2Tgn5CNaZLSqRJ26dzBUJY3OSV0MrcCVJ
YpbHX+yGRkmg3gKuqGoNeqgLwMm0LEXhx6rRkEKkDnW6A82Jr0UgSkGI/w9M
KOG0d8w8GGieio/K9MeKxup2pds+n8uHb4VZJ0OMO+F/owwpdDieuMTwuf8J
wbzzAo0NtHuqiyTN33id/W5BnxQat5PbO/Zh5I7kNpGYkyjk45y7HGRq9N0j
kOBV3MIbTaUlPbbBql5GkxIDyRM+UDPqDpswV8HyBr/B3QcMQcrL0Nm0JzsE
6aeEdYJqGMnYquePhoVi6iz+lF9k2H08+e8vLuw70o10ffU7SFUdvvRoHwE1
kI4lNm17SfSN4odxcQtcOgj71MWF08DTvEyw0rKQYcM34eitcpVaU+RG2cTr
3SuA6+ZZxFPZ+h0dXqU2Ut5JYZzV/YqKxDr43cZD9fEfTU/zvEGT0Ott5pGU
OSZI6d6J+sa22G+2roy4e2etIzwRrgkqdLL81MAIT09zMnuIpuUwKrc/ahIo
vNkVSneFMrl0iQupNgT4RuyJRQgaEx3xESNuWSCdCK+V87caZNKsne4pOIkp
1HWAfbxc1xU4g6y5+CXqnmabYUxdmG+9tqZAyLm02aLeZnnns8h6721n2X9+
O7deCALihVKnd8mND3MAPFN2LIez5vyc/ZI45ZDitKZ9Spk7BdlNabOV4YOV
/lww5AtZKmN3Csxn0o9JtxosH8Df/uaBJm1lA2AE0ZTzPuogMTl7+FXIgiRZ
jvjDdU1c7+dxgi0p61DLBvH2QiNOLUiGvpbXb5nqQUrXQijLan/65YUXVSgf
w73wRhJko48lGDXEdr/5gbrC692l6P+0IyA3EG33CSvvzcDsY4GKSeWI+R/y
u0uaTJcyptw1Qr5+CC1oVCorvVZIsMpBuxLSyF0AwWzXA4HXwMpsgsflsrVO
mmwq/U89btpAE+mUY2g+B15BqAUpDbMl+UNnvtHksvVryGtp71PF65YWEFUB
4rbXdzB/n/Bo9RaYonk8UxlV76hdzQwLUHZh27Cq/TEtYhtsSLtFiBnC7i7M
tyfOmy2if68kT2GRNAWUVUCaTkeNPOth8KDOfx+Ztl4J7NUCo7Y9vMZh5/ml
MnJ89VDlnFNzR/845YI0AFUnhqcCSOK7JtxjJ4QAHjPqvhHD3wFGyaAqAEXY
T2zonQZnnGYBBTVByxd7C7fQ6oR4uxOAr2KLuQX+n1KOMFHLKtmDp4m+Z/ZO
HW6kssPOaofiGrr0w5PUVrLTvNFB4gFO6h/CD7ZLgR7zNt+rUHP2RTyuEDyu
p3q+39nM46WBdYXVvOz93hKg7wk7aB9HNNN8OcTStC3FcNsGDijUPMyEjpqt
AUoy2GsW3jFZDmGMfVrFGM6AFT5JmNWOFUoWVvc8SBrInI84jh5mz+rJBwet
mX2pyWRHuti8APwwLYugj9iTZoC2hPZERVW6/LcMOk5sYe9ymbHGgPGCoOJx
oX50ZM+wZlqhpFtmj/vNWU9oS0I826EMFWBOojbr4DCXZlRxbB8UutumW+JV
D2SJwid9cKJlB8WimRYx9yrOkasPseXyxGFdxNXNa6gLRhRZH1URZetxNkVe
xzpHC4gRIvqoXIjruwJDRTakhdsvMmc86SR8h5M3S4R2sP3I3Hu4h0a4BIn3
dTV12CeZCrjy4L7AyYmdUTi4HGysVB7L2GG4VImRHwd5OmCiL8f7kLLSsBpn
z7B1J2UtEy3sY1oDCFOpFrNaxHChNKw6vahKfi3JKZtv8mi2Dvk0qWtLwtPc
zuw5F1RapuAakrkWSFiGEgHDPJIUcDUk9jk1oB7JI8ELPSzw1WmMWI2HsDRh
lt/qav1NVHzm5TiqWRdkE1HUO0Ql8CtH1RDuMQwR8BSm/cu0F6sjeQiQ8MmP
GV1xFXR65pkDNf6ZRjfnGSg7jdhfjwNTLTT4rx81+JtEyS1JAyk7kBNIdC6w
rKuxzu1EczKnHzpNelUhQsxJcfAek54oIFM8Gx9Ju0FZkRixkPm2oRQ3Ui31
8lGkI21jJdEDWayQ06djKxb0Q7k+S8cHFvHZy2TTXuBY5qp+4zrIflni7H/B
gbP6h6qHauCwBYDUnqWiMzBR0w+Txc0I+zYqh0wKUSrd93XSxUvr9bxNXC03
qcXY7htbPnbe2zfnH9AbcG1sDrS4xhUetcd/Ob6QIRsy4bzBj6TbTbl1lj6o
IRcyQAs8aHKPhfBMWrBRogYzz0mcPzB9JRpjrDQIJEeCr/SmZmpNV2lj0EO5
/t4LDi4Hy27hMtVnpT1o0KRAnvwRZzJgGpgbsaHTubNWjxMpjHNaCVPpx2nS
Ubf4byfgKxf7U8ccstd+/lAd5cv1/x3nzmSvhgir2Jd9qEi4fQl+yLNjI25s
He4AlhU7ja50KxNGtekCMkcc+AJOQ8YKzIoloXasib3SAVDzzN/xMposl5CS
ytxBzuxR8BjrZioPJRHfS7rys0Sd+VRWmOOpatGAweipLxalc1aobc667ZLl
wtb0QxgcTqKXpCo9lsYOUW498iPyYiH5g3ZaD0WDVlDs6LUKT2CaUBPP7QKP
4ob8SdSn6CDX/uAgyMNTM9AzIlRRHa9i9KE17tHBO53pi4MubtDzraO42q/1
42+R8KqAUjshaoehD9ujP2ttBaFAtEn5GUr8l5oBQgXJQBB0ZtomQ1Bpl85j
Jk708wcWZaMkKuuGZpu6AHg2aKqGxvDR6r1eRuWJg9CvlcDdkpm5JiyiD5mi
190lg+LZDHam6/wQ0JchiiK7JxRP0h548yOjwGA/ujOO2g7nWl9YO3dkS7ur
4DEV5ZE480KtOXNs6OJwY5mqE2L+uta+XqHw9vx0iq6Z6TImrzykRPqxuKWy
Ao9zr+o5e2GeaIxN3blMSDt5l9COJetW6t8uENaWpK7/J4o7cECa0uaZSCCK
jUqselHUISgMVkqUJkaCXQpRE9ErFzPubpwdctuRTiCqZT06nmhBwdUbjhKM
eOE0p5Tw0KlNm8ze0T8b+k4x+W5a3N6KxEjSPLot9FfB0Y874C16K3w7gqI4
QhEzR42J5JknleJbZtXgMMQ44mDTwJnOoW6Pm/ZwFk+X6cY075+s923K3ocd
hH1Iq9Dtt6TN4JlmRCuf6UGPHACNWznp3abYuSRR00bjIsEWxPxMx/Y6byYe
tPXnXhyIOWW0Fb5kY6ikyiFjHTOCbZVn8eB1l78OKc/obmhzB9KISnzOzCYs
aRZq5WVhuOk1KgzoKSSQaksV8e2c7TQ5MaEsC66w7PC4BJCopG6PxkFmWpoU
gQsVzvFmFSx4NlL1z+2dKOok7EqGsiQepjQhoH4GQTXjUhPjNCTqL6FtiVFa
xecNcncMipTXpM5pInZp0l7MInWBVUJ5h3Zyjdjh2gI6G+5I7RDSi22JRVmD
0vejqjTrHUfmiCNjF5RnLxVJoPrUc4YorzRaiNBiKxAFdVc8PYk0UYEIKMhx
8HaGeoyyf+9Tc2Y2MAdmeeB3CR0haHxY2vEABuEkh9qDJKmkjwWZhTNS94TB
es2+SjRx+xeS7kKryNPyneqBnaKWLNIFAnImzQ0muITRl473M6rmlxmmVDQY
yNSVXErHeCwpX2BeglwPj8U2tKjUvvk9jc0dfVzAcvfWObaMK4ATwJnoa7EB
tve1z0bXQiTT+Y+C21CYkYwL83ibyll1AF+jq0xbdiqUtpQxj0isgbhEHpNF
k+5K8Mwn6XUe7lsAIDJdulGP2e8iXrAag9gz10W4ZTwa/PoUPjvvuu0gAV5F
tt0ENa4t6SWsGH3iCWvAyh/dE4445cdQHrDyV5JZHNiWLEnLUWMBVWogPwHL
SMd46S+V5vwCJMGFUzU/VPOPG6phcwidJCWuG/aSMniake/9A1n9dJJdGwdA
bhQUH4WpznCJAO2g2P3TLJ+Jh6dQGnHvSq1Z5qKNCDLFjwBv7Ozj5LlPpTzH
rLmeD7XzL8vQtx/GzQeKJQqy7uCFaXrl79xjBZWYwSydf6ZaG/ZwjUQVgxik
PNgEv06v/tE0Wsoxf0gXcf36+UVqTUq+eNijgM4m35aysX0Wz17y8QEdr/00
qf825GzoIvv6x1gGUNYNwEfEIqMSYk/8dzHKZHrsp6U5F4i0z8E0OE8bKRQ5
Vuqde/g2pOySOIDyr9MzTNyq5UaWJTsrQIEoHf8HKPrqurbrsv1Q3AfQcZMZ
g63XbAs3zWKZwXsA7vMvJbMIeM8AVECzlWYa8qJbN88j2XKX33lf22h0z8k6
9FihVQOsXS4nSts3PVF9xeneUQR7cAzMi2NEsqs2kYjlrNtAwHMLaDQMWDWC
B1KqLDfiyWy6nAXdKrq6Ij7lCDPVstSqeka+UPowoG5VuRxi3FpISgzOkCAT
fRDWEAo12tzN8nkXppmS1pmMg9o4AhVHmWxqBAa7swfIAk3t6z4LuAbpEISc
VtQhBDcTii2wXWpmreQZGrCmlPhqBbUsgkfod788wlVEE+GatJ/udvAOZqfW
tS96UcOo9Pf3X3UGfHj5Ro6Bw0WKp5D+luvvcEs8hTaRLeN7W4VEBuxVoLAZ
pqQIZv0tL2n5e3zeXL0MrDqY4j7ODl+vGd573pc3oF78aaJtnEQRXtEISIW7
1t9x+eyaWpf77su0BQVGYr/NCwxKeC8mwmtIQX9GyNyeTHBRwBppiYMLt/+7
M0SZSebPUFjv4btMtNpBmoRJxtqCn89lob/vDZ1Kfg0sR1SdX/zCyADlq9hG
c3MOL2gQe9basoDtw/nsiaT2yT/1vBPEY53poYCq4+ALRnEzpg6P3OAO7r7k
osPChnoS4b+LoXdZyrFYxIBZ9LAoWqmdZ81IPirYWgBsPtEfMULXuWHPCm3y
U2EG0Zd6BzDAM8iV5Wugoi7pD1/havDrHRJuiovagd2NRJw/hXkYDhSe4yea
m+RyLnB6ubcTC2lzhX7CvCZKF4B2oYfHANj65+iJth4mf5rb8uUuzB6ajBow
e6E1nE0hPuQnAwza6KxyOyY+kn6b9VkDwTw+8eXZnUUJoYtHRTUIWGORJhtx
eKiHA3PkS6eFxgAiG5UsVikvM7k1ERYPFTrZ9B08JDGuFc3TlaG+0JXTAjZI
l+U/DwVGF4WiNKCqX8IVGx5PdfBhS7pc3wIHZufjqCKcQ1zqfynFrdQFF9EC
XoUWtCCyPX3hgNt6DGcBPuGOH/YArAb/VCcwMZywfRRWghKaA0felROFs5wM
ciwxvcUfQ/Cxjj5RVdFPk9wlPNI54DxyBJ5b5PPx8fwrzHB8Qby03/TRg3hI
+JIbIMZEBuYUVQ8kdSSvwQgP/KAhuSFUgLiNhUE9bYrZiLx0ReIRKGWS1jnr
nMTj+uAiuQraKBe1oRBMSANbOzLF+s8LG0ZPsrXQ9YpFblQdKxz+9qotE2/V
mTunY8BZg5WcKvn/JdUpst7m1IhmK3oQqgfVaUwNG1ZFjAYcO09/EqFCFkgI
J0WWny2LcAv0mXMG38YlDYHtSxOYDuPGD9W0YxvLBQNQdVu6p6o+CEAHtgqE
W98vPPzbX0uOa42kEbH0LQjEJETLQ/64p/6GIKUkzMpuF9ZQlzq7H/D4zcqB
rYJxIVeYzDXsm9lnkajb6EQHDTPHO7s0g4r5HjFdt0C0zu0kwiAv9wdd5BGA
Lui5zgzdaqrKJNhKEDZ8X0AVNodG7uFFK34TZTHmwODdEBQc3OGjHuoABvMY
aViIqxgwkOrBYG/c1uyKH8zNGk8ISgLiQoqY1ALGJoKUTyUjQrIJpddQRYdt
8yJcYtRfhtfnNAWix4qUPi+1/7QdSOcr+xRFvV5sPa43khln79z9IVPO1oBE
43SfLB8a/EeMhptbz5tB/6iRE4ObFF6yysBFFSrW0j0Ri1HCZFJKS7O/2MLP
Nepmwin/XhPYmDDB2zm7z5+f89UAnpD+jlajd20q+HnFN5c1ckyH9RY5FPz1
pEyxp3qqTe/vjaWojZWUjcp+ebb/q+oMTW4XOdlW76/Lbo9LgLlv7ZQLOCLc
GpYhKgV1o6sW+VhMOibJ98aZhMjhghfeJC+K3D6t3nGstRi5XItYDdtDbeVJ
/2CgjvGVT4OD54cuef8i9D6nkybVEGH9BLazEXFrjeL21piGuLj83JTSGfP1
mcDYgHzvE59XIhYEJMIQwhDe+RZaMZPv12EOzAuAR4fKHomIuEa0BpASjSSY
mznBk46GY5v4EvnRMBk+j+j1kHCvus+R3qxdAIRVkBepEVzXZ6TWxK96zNZs
hvyf4aL461KKPbZsfBbBNdl4z0EC155StilEQBgrzxfa6hEu7Mq6YxEwBDH1
2NaqvEmzr0gZTwC/8k5ty4Aiu1mUr5XPtrgYvqj+CSUCiFPkNXXgDFpi2yiY
pfw3SM902TD/u6fiCofrFucgiHQ3PF4AexUvhfqLg2dB5WUChm97CvJnvbHI
Q0AO1iPWXqVlcVHFeUGUP9mnxTcptCfP2vHueHV+ZDznXy1r1NTGpzR3ZCbV
p7EhIPvdAFKnKDlNoprol+G03Mb9WTpkJaU1vOUA3HQBqWUoIA7QCBvHN8AD
4tlhCtiWUqp2OoVB2EolShNgMUyt38a64kbIjjYRJQLknCYiridfkY5rn86r
iHrG+CkDP5hee3ybaNIfssLmrTdGq3IcQ796zzEopVad2wZ9Yhl9GHXt+px6
aVIM6fNANrhgh2s61Guvu+a/UAHoccQK5MaVp4UIprv3d1TbJfRgtj4SFpdt
f99s2w+sDXichguYCkw+rwMOlJnobupM3mM49AyJIbqfhCEZ0VPlB93pIsBj
XopZzqFF+C6+WKkcht+EEWXZHT3KkC7Fqcf9YnPuLcjrmRYcV24vnCREo6tV
3z9ubImJ9U2NeWMraV/hj8e4GPlpLRKUxIgDYxE6WfPRG3RgQDTK3n34mvSV
wmscua9bMpy1ywYE830+NLLKVenRKz7zUPy6c4I1aVVeBlmenKnJSKxNu3Q6
ZqKNlNi6Qr4eyooT1dLvfuxfCl3O2kAba9G/rmZ+G0Gk3TjzlDjhzGN67P9l
u7QBHUvaezEcy4I0qUj1LgwjCPcFS019MafS8i4SIyeJibTBP1CSxCVy44u1
KGhb7tIzrDEuAYJYOMFhuKN/p5VGJh9uevKaSvy1XOreetWtUAYW32OO+I+d
zLJHV5VaeSgQMXfr8KYol4RHw81H8Sd/CRIJ7bOvGw9iuJd6ek+IMDlcq6Zm
K+f/fmF77KvegdHhEohzyL5aiKk9UdAfs/hmG9lp1ya7PjW/CnDvbRY6RBAX
a55EHhffKpPaG1Al62WdC0ZsphyvLjhRZpVfupn21Bbipvx09QQPZ87yZ1KL
FUvjbOswzC+/Zp8GwxHsocav/tSYFkmlv6ppXuQ8eOPzJ2YGdAxCQSQyQUVU
ccgYNfbK346IcwuW/fSKIIBpUTFHY1zrWp9bILwVlg/5QFd1MepCG+ziUaJ5
Xp439lz+o1D2q6WXAWMk1sb9YzDde3tWX+JN1Lsm5EEtXcyX+WPU/NVkqn4u
A6vPwtJcyR/qVXd/YEwNyNV4yqWkR3p3R1ey6ruaglt4fVqQ7C59klAkZjXp
45jW/FWjkmWfMRyyxVNmYA8nAOmsyAMJ+1hw3NlcLvRkwx0eRT7Q7eTgtzmT
QpoJ7OcTJbCICWfToAEEBr/oyOPmFlOawUSrxo1xkBEVfQZYEHkREBXYVi0K
+owv43YdwBIbOqUGjWsmB5PaaVhCq2UeURrqKqMKhTUCV8mJIJeqPjxQeUUI
gMds4Lgw5M/d6Qd/vKsvSiO+5bh2WvIvlJq8oaTdNqWBZ1JRrvbzbXXxDaIY
LhRctYxx5AYf9kr+uJkG1nzJUfVOoo8sVkPOeeLKkDFN7RGBDRNQ1TFAQ98X
gRXUculegtRBkgDrtqbm89cDW0PXK9cSb5fsELlkI67c1uUCf94lOZZG7ncL
LZeqxm1CVNOkO6iJSjaJdFKXqlW0QfYs63jB26QVoom2StpxYMPhgzWOb7fX
sMnjBp7W0xtgoUYK28VeiW3GfFwePNixTGJzb0l58KtLKpYlvVUvlOZgflbq
dUkro8yOwZtqF3+MKt5Fub5R2UF408AaotpXIwdyMybe1DY+n0djSpr4Ckpw
jsaYZ2EZxX+ya4DGKEBwPo7NaLVyveyxwpR0aGVtt0DbKnDNSlNMp1QL5i0a
XVokNI0s5f2a6OY/gitb4iIwWZIcBbuBdDMaYLiqUQlZNmqr4Ffl/LkVEanb
2yx+pA65jzqiO+1W9LJDUuE9058rmSk0H+xgXpkBJcIHAY/ydXgDNPOXj79S
sDzx29+PnLev9We1H4vGInFNias+0wjlmqRUdP5Avn0FJPjLT+xcTu0XRqTc
oTi6XqszUxbMkMtcxD3yt9RFPYlI27ucMAv1hUIsIGiXvV7ifbPscHe3Whm4
ugPOvP/2qCkTsdEfHpcjpFffP11vp6KOZo4ORtbH2sF70YbWbHkFYkEFHO37
i65qX68VmXatyBmgQhqQDGI321UMoUGNVNax3J16PyZ5IhdM7IrrjhFf73sn
pSxxA9qWMi/nhgPOmRgGZw2eXDnkcXnBsFk3a5HBZGgl+T7CraXbtExmfyQe
e5uIX/uPuemm9XcKrNn7kl3JH7OtlYT/vw3tdw1dPhhneNoBQz+kTvFdFveS
lTTLriOcYoRBDCQwA9HAUJ6cRsIeWKwvNXVJ6/+pC5/tOHnWGClOXNoCFElY
ORojkdZp4hZOhzP0s2RZN5Hl9GqV7BYeEvaL+KqxrR/YNd+TZFCuwsX1z4LC
6+2SAroV74v5L2N0uilkCuXQnHhFLTa7MW/O/TOpmtX+07Du4l9wBF7nSNPI
Olo9XIPeMpuVNQxVIt99/W7Q8736bv95nPXny/+aeTJRScbpyhUyNSEdHOPS
QHreM6ysK7PZGbx3PqxrCTEhTx1yQg02dtNDxC0AFNiZNPT6AvhKTDT/ODwj
PDEFJJovXtP+SdvdCUWBqmhau1yMBGCTONlq2PcStk35FBTdH//d3Acvd1GI
nNj35JQ+kdrmyzGtBfBNeEg1Ife3eiip3DjZ+RZmqg3U3LBZN0HL0fL/CA3y
tthfh+T19cO22ZJpQtGCJGpi7IDrNw/0kl7UjIzopEDgA+8AH6aDusgbRgWo
eq31CI+dPYvKFLjV9BjhlV6Qfhh0rSo+Nb4Rt3ITzBz/pdBQGWW+DRhNdG+/
9S7l5Rk3C/G6obLyIMEgIl7w/UEiocyoiVSe5lPl1MpCOw4rbYKxvIGrsrt9
xpEOJe4rqKscPZQNdu1xMJqH5ORY3Thhl/D0LVygfjuoLf/+NbTqadQWYBW7
dwFn0uCqTqhIzpIhooGRiuQfxVl8HPO/Z4xYUuupCMFKbUhM4880PghDhXn/
c8VZ09c6NsyrvOzjxYsJD/6sehIg6ox2teoBRZbxfYDSJLMsHfzqmASFpPka
jsfbMI0NMXrQ3pUUzqaKarrD7hs78XjuMb4Q9eAjk0WztUvjN4XLk2YSSI1X
CcrGKyXpYjyHmg6iUx6qfjNNmXYlkcA1I316ZrmHrbAvS+YLyHeml/sTHDVp
xqK4/ri+btkeCxE8+zVx+m2kzBx1YbhavXq8X7FgZjhs9iBe9E9CFFE3XsE8
TiyGdUUG5qcAkMS4lMtG4ILrR79HD1AwFQCi0DmAIlwDsvNE13ObQOZef3QX
vBEsW2W3B0VLHCjfgdOZEu+Em78UpCTB7sUYsuXgX74woUr2zZVWzTUw/dPr
PYyBZcXZxkqEeEcBSjLGhNCcg4SokjgiX4DBZMXaMmLfACzezccVI8dtsSqh
s9ce8Xch6nf7HRP6d+Qm3LA8LuWzeEHEHzTHiht7RhE59oN8tTZ2lTaIpCvo
r3PZROPZc2yyjyCNsuKB9sth4B+C0nyxc/W2gofAyHtnh0u9fy9uWl6FoL9S
VlkkP/l2hM6OMTAwYbGkwsS9xtDnz+G+/BAN4z1StGM/d4ipWFLA0ET0nP48
pk3vYXIe3CGvMCECyStWyyEwDh5SuspZfU5sxeQihPg6iJCmV9FIFZypdwf+
lJIW4wa1vYzMiiLt+CxQyYxlhV8MqTYtis9PX4WrCxZpRPZHqVW3bYJugOx2
hk5xu/gQNm3YTbVhIQqCvhQgIhOJDRswpN1whZQdL8wgUROVvd2Sr+nEqgqs
0ZarF6cwPO4y6YAnc3i6tzT8VlKtHQ1omnzfpqoBRLdBgBZxAzrzNqRGapuy
tiehex3uhvFeakz7rpCZWsENYtlZ6/uPe/ePGIaCposUTTHGyB7QDwBsfL0s
DLLaFGRH3HW1LkhV1V5HdlE5P2stDFc9deZh2kQAWfRaTjDJK3kJpvzfYNLn
5XBZM6pp3mI58ZLDh0PoAFjfMfnSnh7mMQFgXqHXqh2/DOsuC8mxwI4gV9dd
2m/0iUTDEEREMuqx49AAaNkxQ+XDFqNDJ6vsbtP0yEpy8hE8d8DRhKH7oaVl
3oRVdkxGuy7mVlQlulGjQl0/GUVsHfhbhN7Fu2upoHwxYRv9IQxLEEe8MR9U
blnr3XuQPRWCEHiXSYgzrQEut8lSNGs36nAaVfi2OhhBFsIqrV+0d3LlAqpI
CDf3AREkogtq6qI/n20PNTgMTmRhKUEPPfo8w4WJIzEk6WGmqPX24mRjJZ28
opZSpQPHaD0foRMXIPsmY89iQaghIcB9YgvLQV7LTFz/3zx016x56KVisF3z
GD9mKuViuGC48iIEkjwLAyDrEt9w/BlsqEBSa9Es2jFUQ9yp54iD0sW1vzRv
axqYVmwPFTHjJrZkP6jcSNybCy3bvGJ9HwXH4Oix4YuwA/DV58PUOdMiPm27
nkGkalQ8stCX1vLGPsz7FGfcMtZzvBchc1eu5E8o8Xq3+eQg9arzxeADS+Gr
PVyn9DBhQiCtF+eVJ9oegOZnlBb0ydF8SEAC87khbB4r9slMDJ7IGMiSLWTM
12PLc9TPhLV8XSlJBKpuVwFN+jKwLdur2WWApuz7CCYOqSlJ3AoQdHDimuni
QZkSjTijM7NgJhoWqALhisiEP+i7JqG0tEbLGUTPjHyihLzNgDDf7ImJdI0u
XlksqIAMlUxNsQFjilDyMwEPWe9iGJe0r+zIzKvFXVlQ3A44JNqS/vg7hFd9
k05UZLSmvbJy7BxBYPS12yIbiUewb5RRu3EomlZiGQYojVE7+aindS+juGFe
crvemwxpeuDQYXYdiIdkoCm72oH95h4ebImjkNB0qACt/L5e/hDqeJ8F8sqd
UvlEwGJDuSPnD1UlgW2zW/8vnu1b6JpiQnK5iTN4H7iaRGzk0KMpjdE4WCbL
qHMmetBP3/WtyQf3BrGC3pdM50AZZTG+mIaPxzbnbAJNeaYrHfYNUjrQl7nN
QMg2U1Rst5J86AbVtM3y/etreHaImkU3y8qGReayWRDf/tIO7LuoDojdH6sf
gn1whGx37IyIToMAqatAxirMDY3gRwfgTdymaPNFthRYyMCRgt7iq2P4hNDa
WNplRjQtk9iwMmuo+55X7mJ6i9DjSabK7LtuWAC85mp5qtafWHGAN8Nfnv/x
mDVUobmPazOiBs1bdW3HNVbT+6KvfuXnZCOg9z5gOqu1p1KoBO/c75xyl5LK
xvghB+Mo5MEtwc+bq7IBFFegyaqZ3iW4N3ZhdsXQRg3O52I9aXZKfvB77yhy
KEcL9Jz+mwpKCeiz1r31eSLwZMlBMT8Zkm02abk79V7U96M6q3TnrqvxCmZC
Gy0erMm69F0EWsXXqAXLXR+egSJc9D1XaaLrN1tvWNDEZY79ALk/5+6uuU+k
uLvHJY8LFWsPO5qpxRNzX0jv4pA26L50n77qIYWyEgfC0T4ueMPQAnacDB9Z
mkLqlQwfw3o2aNUwhWRhajXZ7vRtL+j1Ul8gCLViGxLrT0JsWhcmJM2QyFo4
M/4JReLuAA65TmKXthYYhhHwl9gUyrPiVjKXwy/ebUwhx3vvo4GTFPmBXtwL
Sxez+BDobi1ro6ZkWf0UhMT1TFMXqJ1VKw4kFS3WNPGXq4uEqBynN9Y8WPPi
pkHkrwTJWLXbAEv6jJ/0v2nPJMvGaORC4i1c4yRo6m5NjwRScrdpCiDGHUaP
B/TwsFPGuBhydzknLDvakJwYUGncZTWUvrUQicH+vVMvUoSt1d5/xmCDG/rt
pE40QiWpyyqUXDU5TumZ37JtVq/zzT90PX8CxIU3yYiYBsUYqxtdmPbX35n1
7EwjU69OY2WpB9tTi+8/LKtYfWa6aVBJRMGSXnbVZYhftgyoN0iKTkAy4bSa
GN1Wdu+k73vlf91Wcyj/Qoprn9x0cq3oqzon5LrKSGilYrbrewT+2ZQIa9XZ
U8O3IRyGG+ub690M63DB/14Pq+raj3stcR3DrhAXBgAOPnH5pUeuEmffxpfu
MrvsHD9gOIqHKir9s8OzBhdXRgLxTATMAJeNe0WuvKVN4+vNrGmLriyX9v5f
npUQ9I8Nqj058OKmkHeE0Ec7oig/vm4VZhXtuQYE9OGNlk493ogSfj1llDZR
BMp5tHoX2UfbYc9nqQp8hfJul5qaGRQ7O8Damf3TEX+W5dyq+lkEV6La4hkn
MZi+DZTcces1LBE1xoUCqs2pbkBeLcTi1SLWMC6igaGelyqEC8ud8ZOU2Rni
7B1t9zy/hkPjOboVhykO9XRXgsR+SDkx0n4iEAcEWJVmVHp+PxZr7nyv9zj5
FxfugcPnfEiip4gsddr7PRTjIKwkLxGIm+5Wq90ffeS3rFq8PFM7WzZcyVQh
tPP0ZEVyUycTfWjQQxYXvZBKUaqipMXN4qJk/z9ygkEeOotLvCpnJVg0c1Ai
jat2o1DdfKcv0e3I3HaRMFWfJPnMDCfpYSAPTZ54vS6tPz3V38qzXcJE1fGF
6pQz6dBADA3lFzlLKs9ykAn1dNA8yC2N0DSCLeDeLaSBMpB/bcMK+jelQaia
Q3vczqtvzeXqBDECegPMq1pUmA+RoWoe9i1HlWbiBALo42jMjtGJLW6RxnRj
RMRz9rP/dXE3yVPWc2GqRkOCqG1eWDiiuEzR8OzgLFUwc/mo8Qc+kLqaCWmO
E9QmSfxrnBBr+Kkvh/0vQRn9t3vQTGfsvhiVP1btRnPDr90w+P2HaAKY3Kbk
zggmaZA2DbWGzAA+lxUWmI/5mQS6FRJQyTXzwQM6M7jefvqI8Jwh+p6sWdtM
KTysjIq5lPWlKilXjwGS2WgidzlQgqbzl4t8zDdxX3axkWYP3+ULKHHPifV5
M01ocrXfi9NOCx52q5wPfsoCCFPxFTTTXkhu139hO1dL7OtpB5ND5Qu1ElMM
7y40dCZ1G6WKqc1XoCPpB1YFvNgQuumQXhVw+RNWqznym+UmbEXVYP317zLe
gxj6gxt/vUn3quuNjvDjwNyVfmnGwHuk8WkJa4mgCjrHoLCebz4SNohSIQeD
6KKpgFqDLmfnSfPUBTACgZzd0UpDyCmsbSZ7QtgOrvt6fYlq/haTz5ANaon4
JnKwI8XpjLaUOhL5hvCaIh0pVXbJ0m22Wpfphms42gxhPeOnUU/FvENWgMWh
qnx+3LE2yivG+MXzLY4Z2PQD2VOUQSm31QVUWezQz/I/nGRUoxV5s5jLpgLr
9mYeUhf5GB2mEcDxibwmPKgvsmiKmIGX0hWdhZgMZzAQXPbGArQXScm9AOY8
TyloVC65sH+YFndk91/vC0Dd9KVx8xlqWOKc34PWIvLFWdcTcHbzi98SHYMn
djCuLYkak7qZLC8FLuaqPmV9pkpri5ZF2x8cjtYCCGG6ej/Rj6u47a0ctTYS
kQbBJ1rBjeSUk1r6/ha44AH47nfoFeFcYAWoLC+jgFhHxjY+48+OQGyjD/J9
2L9OuiZ3hNke1oVWzqgqojesJvcsOSaMAwhwhR7LqszMrR2rNGu3G0ySXil3
8uPNqyc4FeGQg8XF2DzaWpw1E09Wnxs6NPbPVn7L0FSvd1mINOyDa/X9SMeb
0JHFl053fY+NEbywu18NIkfBtmQWOBUZnXq5KA82g0FLEv0TUECWc205den9
Oqt0zE0fnkltEEqFBE0IopRvNYvo8cX+F+P81jGloJBECSy9tCqzUiK8kKdy
6wusUvI5lr+eWkQ1ME0GqC4+Ai6V6cS7K74qRiwcpS7ceUjlldu+oaqUeTno
yXsk4rtQPYssenbWNURF4WQK2wkZJ6L1Wr48N0WJm4OpNGQSQ7rhMJvOhW2M
Md0i4L91kytowerzTCgV1MoVvFnSRcNIeD14rYqQkweXQiGliODSNTWujcsx
dO4E6P/mi+fQzbZUsmP8H9/O++SLWSQSCjoJWtKalGF/OdW/7xBMv8kElZW+
hGFzRPg6IcOJZuTFCPjNfabLqwNwszDDLjbEBumYcuvD+et3bMXjN6zAY4zg
fzRuhnuQ90FzpLtZHsng9VQSWZWYJ6oKEm/wpUgF4PN+g95vgyt7ZuLjMGzV
t3gYB7Re93hoh/xgHUNRA4apxy0/TAavuwuD0PKz/et6/+sNcNACSyZj3qYp
YhKJ3o46F/MN3pco2OAfTlnJsj1IB7CEH1MTEFXwoKFwJ0gV6yS5Ew4TCe79
weiaSv9YR0gnTPZZhQ+JWM+WPn32YETkEJBazbZDZGaZk2L+kCJZcZP8UVvT
MfxT6/gyyEkbhA7nqauY/tiZHlw38LMhUEXHBbTzI7IbcR5mz0nIdWLtTYGu
T/Kc+aJ4DUlIgYkrm/uGz48T1neX7gF5EFpxF2V0a3fgpI9bLjJWLWdiNQmw
Yi0wVKSayCxCd/uFBYft68QjB5dkirKfKoC4P5FtK8KYNOswTz42A4+SRGtV
swwgh63oXPQyxhk6yfGHtzXag782D3XATzRca+HcsyApTodXXhKcQcmTcTKl
QvpKssjjviTvUO6Bot7LHT/bampHJa/PoboziI0/osWEJcvoWhT7l+ihiojl
jf19HIJKDUmM1kUJ2nM5IMOjGD5RNs9DbTDFgHU1O+NX4jPSH2/JDuUsL+QF
8rLAjqtn6/eybOLmcZjIZ3Ah+42hcbmfH/Y6ao9LS7fmHF7q9kvkzqmLbpXY
+gHv0F525czRbuSgVcROvjUzV88WDS8b/+NN3b3l9ysO//YrBSPPU+MX01SM
O+UECbm+bF5fXj08Xkl6QYnVpJSXZHuAHfimNKcH7jDUtdBSTFA9rY15Mv4I
TF8Gbot+mv+9R1HJct8C93uTKrwoTci1HyrqQ5d9uwPzZTwv0D4bWNSnPWyu
aBfoQVAAzi219enIJJL7qUyVTKugVy9nLa/urcO63S9abUPS1PiogTDc2bTU
YfNKR4TUFTm5tZYffiOkFvXGfQowoaI5UgnpoTWWYqmLluJuRFJc9omXXXel
oFZkWOEahYrrialFFc8PhfGfpsgSm9JojopZxUcC+Ych9HinAHMyhfEdUP0/
kNpIa+imQTDL8MOGpGoPnJ5W+ITmrITU8WHaqWydNFZz1X6XkEj4+WSZouVQ
RpYkhcwEoJC2aRchq3uDHyRr4eeBuevA8Wh/4BNmedbtw4EYSHjioCyZZghn
L6a3jBTH5BoSFr2mbY4PUK0NzR5I6K3WcRyu6HyU5gDtwIkvwNYic01RLOKn
3++NTRKsfteJLnZE4gGS87uZR9rce+A8Qj1fYm2icN/YF4K3jtFqW0Js3JqO
w5LY1k70MEirL5KU5O87D0h90OURYzkq41SZptC6rUrENUJrGdZBHoQrszQ6
V9+a0GFzM43+3DwVH7i0H3KxytA2wldb6pG9mj/7S8a8pfRNXrMmVuRmdusY
LGHiQshX62sQdQz12nQhzB9o8SB1QMoEKcgMSTTYdOVnTiVU78dowbhynlKT
d1Fiskw8G9H/NDHj3/mS/89Pdy5hk+jYYGNNiuTYnLSBGtZo1GcJHaFe7/Bj
TL5FSQ6CM3xnQQEqiaYEuTkt1+mhlm047eiNyUBpZ4RrGfj5mkaTN/uGyVWs
DZBYZlcgL+LjJzprUq8iyAtytchJc2iIEqtRudO3raONleYHQMYHIwbxKTPz
EZeZHd9YCP2PMvtgxOlrftmPjh42J4nHZtvBPEAGXKEC091pryzU1e9kVZ+3
uZc31lm09DmX1dXdHnSscxeajAGKbtDqsb3SXLsItd7L9v8Q9KztNHuW25Y5
WQacc+YJ1Ff4VgHlcV6BWXLdQLlKBh8GBW/6aRtWeiK5gDykZ/atuhXf1FlN
WTNpGO78rUDfl8V7+HeU/P7QHhmOYEiyKRfihZG2ks1DSVmIo9rsf0MpZ0cV
+cPYeQugHN7gOa4L5RxTJsvjuTCPFuN0vnGVJDQZk2iYwBH+Q19u7E6gDAtd
UgUGjh8keuXKN3B/92LFb7c2l2Nev6hjXwQYxyywtFEXNYfSUvYB6+PT5Gdd
SyMr6+hG79kSGU+2SrQDWrOsjfRyL26YoXeqFomSojBzpuIPcNZnOvrU7JTb
A8jIHQ23TK30mD0+rEH1CSX1iD9WQjboqAVnJIZ1joRKtsMS7/bQ53tRq+1S
S0x6B2l9rr/PYw5PP3+aa9nIXEj7YW8KU2+Vr+HXtTc+kcMp3mhuJkgJvgS0
86rC/RaVeKUfk3Ne0leA5rYURDs+6GnDh+vmYBZLrcIVVmlq8t5Dsa3KQZeR
yr5++C4DYErqGvuAmVvdNRhQ9RGZzRA6SEwnjwC1cGlrd9zPqyMxXAQV0gbA
QtN4UblibKqma4cwch3MEdzCMIBb/2LCsem0AKGGsUH/7SJW0jbtsCIGpjwN
Oh2mIVS+kMWO0SBq9K2y1q7djDnLdfbeYZkm4lKa9qVieFrGpcHIPSoHT3Gb
d0WNsESBycIUjJwEWp/s7sxq49mMeK6szLv4YBAQDUG+tfhvE/6KfHOHdbCX
yrj4kEtCUcU+iIfnljZy77fa3XTHjjkpqG+oZG0WBm4emN/j/5NVboNr6oRo
2XYGUrhTVMCsNzlrvkif2GQk9grBbwOqg50FDdchzkkVCTTBbfbQ3p1pLwqL
SxEbtAnw8jJAzroubLLylSYpryVJ35W8+i6T0O4MLTIC7XTmLQIYDQ694wyN
eWpESttAflatWiPpP4x2umqXL6jIusQ4GJftH4S7r1rCJd7N8bcIv6NSfGb5
K7ZjJkQ+e6Da2yxXwe370LjOIMCKE0yB/P5dcD3FKZkPkkVKqKhFI65+Eg5s
NSW5rDcQW4E9ABqYcOO4MpjW8+s6TL2i+p+0niaB4H+T3/RXSjr4xRBNObZw
nr26bb75qLb2VR7mMmy5kQTkz2+SxoML1m7sS0z9dqsy12Lc6YURJifTdGOH
qzMBEClLdQ29wXHVhkExCM2tUH6Ba5GpXGQeGVvAyK3AcJYMKBy6KGdb65ZT
5EgaeTMQUS+LmsJ4+eswsSpc7AsVuelR44mndmQ+2VevMQbDELCoNvWrB7sU
j97Oa5DjIv+DD/K8MB+JTGclGyaW175keOMJ/tqXvlgPOvDJ7dhIokzaFBde
N6fqIcHjnL+VtU/oJlmIjo1TtT6qK/PpnQnmCUafeZ4TrWqt7kx+A8GpjLdG
e/ro6ConGR/faVhMI6ugbEv4NXi/U2PL5GoBG1XUmJGMgKFCeuN70Zq2bpi/
qj+3Fs1Yrphj3YsXtU8DG4XZnDasglh+H3rTm9NYgA4NfnGrX71fDrXXknvm
GdzPfH7KVWEqCgyPLtraJ5HvWKCCSpOM6AasWOwTJx19mytZnpgN8OpkWg0M
/MzQQu7nbN7z0coZtz3JUJUbzcisnq1FWmyHeM0OS1GNyDf8p2c63LBvn3gg
TQNV3nzQ+qKMOe/kQW/nzdGnoEkbHin4wRAn8nkGxyEdjeqXYwXVWWVo2omQ
Eatbk8GuhMXZgOZy6OamsQNeqY+irouMZAEjh2rv2KNxomqu99MN7aF40w06
euAS8tgxCQikddwXkjC4Wv9HgwKdkER15OiX23LKzMXs27tQwgFrhZ9lNxTG
98GeWr5KPHd7f1NU+sZs0MK0G9l4+/RAKwZT/q+cvVZjW2urm7eFyVaAUkng
C+SDq/7XCB/Ltdsw9KhsK8vs9pkzh3suKRMcxIVbfaQ7yHyYe2j8B5V5cY6o
NAo2VgBOMYhRvxtZlu4qC5rd0V+pT6nNIA77mfHlzfsWw9CH540KtMOZzSJN
qtz6yxrwHximQf+udRs5HFHqxPRAUDlZ5tQ9d+iFdJP3Jh1uhK3PwES8ErYD
RHvtWqhVcR8Ouyh11hyyR/bp/5qR3auX5GNGFoYxs1rcIm7W8+C4leUHXfPo
St5SQD5qaF4KCADrUTnM2T2HkhLq6xz47VmGDnC+ONdrg5ayNK9mLHhYU4Pi
ZKaTgnfyrG2gsb6qma7qs/kspEAeo7480OW9UMs847oj2jXRH0lxL9CBM4Gz
dnnNXEP/ybR7KuGRoktFMYc6y1e3YhrmwQNakhzHGF5W13xEdaldt/oxPzRu
SoZ6jsZsnnKhcqOdKc6u3hm7/tnMI9RSSkEJLECNy2UNE0BjdSKCLysGETYw
h7E3JqZU1OxPooVR8ODZjMMPShvn0tW5rZ+a/0Qed4jY6hLAgCiJ30EHxRJY
n1QuuD76mlsq2W7yvx69L+oI3rc8KU6fK28EbWnyvdbh3qnDA9eTs7ntE8VW
xCW/hzlkUP1hokDKdFw6Bdt2n+EVKYE5be2sRRRDf0oJnrsL0E/IfrI1IN+Z
7T6kAWqZjhH/2TOA5LVZOQPF5SjhmGKc2UFdMhT61inwkSoVkhCrixg6mgDb
Ql/q9LRYDMcR/WpMY3b0k/ERaVcY6naxqzjHD/CXyW4AGhUWuz3ns5pUQOKs
R+cjeO8EzAy6rerjXJZihFjTbD3wp9OC3DL3DI4GGQRMn4M29kB8mlwMv3GW
Jd9ZgnyEgmh+OBR4zh0BHg1n7q4FLKu3opc9WXcky9LHagIvElo+NoJMZMW4
qZQjwJm+8Jrg4QwmHPHNiDNhIX7+RVRs5k7nU+QJRqX5OL8O9eYHMFnLYURo
YPcFYaO9L8FmKU9CTD09sBOHE/sqzZXGw0/yAOb9ItHC2FWRkE8dqggSxZP0
UK6wWVWr61hfK4KKUs4j6YeCGS3TGFU8H+ZOovsbpUhuhXYWjUbQukf0h3nQ
ojAvAdU/fWb6kyAcWJbcjXffztXkUJbx6kEzCfjFIM6L3rqhpFNAyVF8XPYr
ski4/xVZVjhHYuLLNz5oxY3pH30vcodExceAIq4g6KUoKXf1WQdnYNrOdLEg
XXNYsvWabZUDq8Tzo59xFHUrs5rg51c9H3mRmGCBTjL9Bd5dDFfqpUIq07U1
qgZH77sOYzutPcgWWp9oUkqk0MvIuX0EM0NACxh9kGHWS8KROz5idUAQRY3K
hi/IQBC+FoOUqxl0ssCOmTm46rJoQrWMrWklZJDQh9JZ0RXDA6TcZFqAasFP
qKAn+1j/OqzrexWvsP8EHdOdsa+8klicE6BVHQmJ5BSEUQOYBeRKSD1eJ2Ks
LGZOeBofBpmpaCzc63vBfLrkG+pvjEWSPFrtkGe1pMMhQjWBeJlYx4YOh2jy
ZDWRcQXSlibfNKZsFD9OqGgKUFtpYi6fci5Hfc7UWmNNup+rjI+4MsBOfCHI
f8JiRL7VTZKvOKq6OpLmCKzpTRREqBOXjI2BdN+haKdvlAaa2R/wr1OY9LyQ
cxNVjaeSke7SUWlndBPzonUKxk+0RdIkFSMq7l6pRurGRNC2+Y0wT0JEgL8C
H+GAPa9GCwT4H9tZ/DeXaIscDpx57AtqpsTGxZ9Rr7QkKtXKMQgcjgBkCC6S
BWU8RYwlDK20+UvDJaCNnd0TIVQj/Cuhz5jOGEkB8WTi6hNpb8xjp1xbDXsM
wumlB0hMlBzvobMaw+Yei8dnl2HxA25C8jkewCHV5ais22syQn3B6v3kauKp
zsZJlcnNkYagNVE+aahV3nb5qPfwiXznRkBphGmIUE92qfofXflcSgzY665u
NY9jZkVdmix/SXOOafwUJnnNoYgN+B5ajU7yUo5T8DcyLsZFhQStFg3rnfkW
ky6UepnZ0m6b/MEiNKIUFltYXQrTVyIQ1QPl3L835bI1ii46Izy7LuDcOrYk
EXxIHp/BMSZ5QyYpM/09TUAmuUnAkSlImsDfAwtHYBRPeUVv2T3cFjPmklDI
m6ftOMGHWlTOaI+A0YlkkLnVRXXsWi8DE6BRCHyJa+ZP0WRMYUzFzPXjWE51
t7XQj3UGP+qEYFF6BKrvXuktpxkCHd48z6ChvKTPnDqpTKFfKQyB2vxaR6j9
Cjr++OjfzjvwXNQxzBTpIu9HS/4N82MmkJD4pRMfk7rfWOsgG32ZiRa9dpNB
+An+5WbTMRPSbte4UjG1VOMWnsw3c2z9vKnNn2J/0lJlHgFC5YnuCJGfrKvE
GiStPNVTnPVAaj8iwFIQgf3LADeh1iGJ8M6i5z9kD4m0NyXHQXVlr22VTHus
RU2Q+oIRyRQedG65vRyW/ywLdY2ZEZTjIWgf+QQ2ItnL7LvYlNAwGcO4UHDb
pEUysNUxMTqoxIOHr7yKhYdsOiuKSvH1+pNKrSIq/2mZzMyrC4lPX/56wgfV
tCkFnmSysKncyhn/+N3D86KDmB/ZRcvuQHWqHq+2UKZfQEm2R7cX1RXGKhuA
xb7ZmTNlvqDzMY6meLHxW6+IvZbwT8ie3rycdaO5fr6a8yWsdLi+gU7FpFAh
nZbBxgDRIAfZkcTTELuY7WEET2sEtcWRoOIq4a24XhvWQW2t4TF+kNXTB3xP
VtZbpmLYNItRHQ2s1IWmMwttzG8hqRbhv7LyWP2BAwyYrrjmQd66o/WSHXO8
O7rhVv3qOKQpxtWSS1svsx84pT1ceOngckb9BKsnszaYCdom/sr6Y+ehaHrD
V1FILzFq8Mw+XN/l3xJ3cBr3S5OpcCDOawTDwAkpecP7iYnCYZFmTOEtMrIn
szd+bNxfPh0HIO8q99+Lnx3zhjFOfz9cIMUZ6ytUvTbdVbRvveCvEWHqNozk
DRst8CDChpZEft5Tsi8jFpi5KiHO3451YI1qnU4tOlOdJNWrg/UbNctRzJn+
vWoJbmW3hF7csFpHPQv6xewsrRliyAbXq9XM/cfCQYvDIgISy7qJmjk9imV3
SxNwcCPc4USQhziHSH/WuXjvF2GEb4vEpcsGlc8ogBF4DGnlMiglcHGr1aYk
IoJ+EG2Ew99pRRZ0WPgn/i/5d68l3SjhbBXcxfRmaXfjE1EpJwVXrcVipkeU
miPRBaG3QeY4Fh/y63NYVA7P5PQeX0LzHuJNJYVZKe3S1GFpq5wmbUkccp/k
4PqxsbcDs4Ab6EK4nqUT0kyz5pAFxn+7tKJZ6PiMNm9FCfhg47Ry1sUeOcas
Qor2D/MC1+W3Z8hdjBKMrHD6BxfnEfL4wdQZUSdojIdzIF54bmJZ8ew7JzIR
M4RzvCCwHODgx3XYYG+hTa45mtcP2aOyGgRj9T1uqjxWTtePGp5cVY97mKT7
Wp8cadsjscxIG2oIk0VocSqQJuyJ4Mgf0YDZ9W/cyk/fWar9rdP/jsHzr9OR
U7qIz1jR+DkuePD9y4XPrfG6dvEt2tmy9DZ7JaD+9/6gD0lb4BUCytD8pVmq
6+HRXq8kEylEQAY1CpdjZvVJ/SQuG8VLpP9EIJsLnq1svV/1uDnlDG1jn1qI
7Pxyijx3Qn/yNPLDAv/gfAzUMjdOuBYqT3f9L3hUw+GLDXocyeHLLR63Q8kV
GPXlWRfBTY5LIOVLZYdEiLg52YOnVvZRCHQf6z1z1GXAvcdCsY+42aR1oKY5
6qwDgmpzPEoY4cocrOT4YoWFn/ubbr5Em4kPWZlJs1Qw1Ya6ZOAxuk8biSWd
U3U8/iwCVhs3sSXBIC9qmLtiLfWTPcqRq2xECfdds65ct9NvkNQrNDvkJDIE
x/mp7ucsxo/XOP1JvJXY14v/BXQPFQAgypw4sCwAMHKgB0HrQU/Y8vSdFm7l
VXzwpemlT1Fqy6Z7b8RGfnD1RUYG7x7EUsZsWwGDU737dBvn1PTNoQ0EwsVu
vB9OAK+W1Wwm4+wNlwKGjrXTdygyabElJY4ntcYmCW7x8LEKlgx/bhX51RMg
Rh0xgaruhth16PdwdEgXpxJFVHIyiO9KeBn/6gHIbj4Jlg/rxF5sM46a9IMI
GOjQlXytKTCmMoC3Jmjoz2zERCVOXItcGdwukM2rwtp2WJQzbr80zA6L/aeg
r5LOh1gJNDrE5RLiXX2n9iwqgFBGsnjwrv0AOlpwe5bSh8dHlEgie/e+HqJ9
RwUxvtrKbuIWOnXWnZ08xTDo1j6SYj1ikR2fmKRYrrbGLUPmNiNfRhJkUaZq
ZK1lWpLumwWH6i0eaL2iSVOeokNjJLak5xBj7Y29tCLZvXWoeFKQ/94/fH/2
ufGcrsYRRSqs/tfdmr5u+vyma74CmVS/JsoQL/cakrd+gHmNlWklTUicPFZ8
l3cvEXTx175bAsFhi9dJxbKdc7L285425rganuI7//UlalTfkL3EMFLYBR7L
blcBlrltNmv690fugRXkkBGmGm5Dwcujf39KAWPQ/BH9T+srdeDmeCsofQ3Z
F6AoREzYn1xaNVqyegpto/qyJrUllvU4bRPgq3kx8GP21E4+ZU7iJamE2BX/
mu6pwgYFkT15khBiFajUQzcsHsiRjoAdFurIM7MRolCWqfPoZDUUkDw37L1C
zaUIaECAs94PVpMX9nvRq4xZv3cK8MIFpUQy5L8xJtR3FMEd0ieE3/rTPIS5
KOOCq6DIBn9CRxTUqdL8RFVxcqCWDwMghuMvsxngLWrDyJq4Cf9k5oOXlIdL
90H/pOnTZD0RJ9ryQZN3mnx97GgpyjDKzZS9Baz2NGlNukW+gg8dUXm/a3F+
LZFquwV6INU3ebppZI6LkL3vg6CkjrlAxF3yNA4FgNqUfBDBrYAQLyuv6zfv
l84sY58M4/EJiB/YZlh8kga3m+UnNbxhoLX82fFJokAuSbDB+ts7FlJqFJde
11Ru9nVJeZ8IZ/7IO2D0wAdEvve1ik/+O7EOWtw2abwRC1O6FP7NGEfmYZMS
nNt5WjQ57lEXlW5PzbMST/84RNU/Q4EDjBvIFBQXrCju6PiPXYmMU1N+c2lS
FEVoz3sWg4eglgEQb+KPQj8EuDmdo78gdhv+flW+ViSjlX6EERvtQrdgl8qB
GebUmJHG3Z6qgmKCC9jljIi+N+3UYuIE/TzYHwVyR2DyhDcmLnlxPY9qgmmK
8NMaa9vgGgW1f6rL/jVY0WXmVAsWqEEJFXgvuXo9sSYtSlt5Ea6L6zpr9Igx
RKL0dbe2FxhYyVwb/BKlEJuXPbpO/7shydg/Na1MQiqsRhvc8GrxfF8Fm2bd
iD2sP2Hwedp1ebyVgUATwqCvVPRO5v8bAm++vU97PKWobKl/tEDdJlpHrovE
gz7CBztEa/kpJwdcYvvpSNYfYv2A68Hcm8YYon6mBy2+ZpvgU9j+Jk9CBT2i
jQF5SS39JhdEeZQtYIlyFQXzo0A69FFB0VVPFDTin+9oIP5YlgSMDCPjiJ8W
5ak+RON8nInGt5X0v4RzsMJw3IJplrIoLvuOmy2pMCroUVmfYUuEmMfJ+N/2
AG/0zzjRhQQtGfdelyR5yomwrkvzfGQzoe28s+ka7PPF8ASN2x2ffzfIktxV
RZHQbhq7wPX2fvlMlb1jnrtTov41fgd2tC+RNx212NtBSkN3Q54w0Om9mBNZ
OnHNdlYLqRotqC9+NvXMWMl87PxTb7NcPM4vWdv9x0lMCn+3CzkCriPS4snc
WV0RRqH0IqYw4Tm1pwz3o7eWVcqVWTGCZZVAsReZGG7eU/+p/BELK/uGB7Og
+c55L9JB7NCceBzHNb2aiJEE1p5tBv3CFTZj9tA3h0Qa3/cKbYdX8X0ulucD
+UOFvfKnH58jK1hntBtvAniYn4VNIfopPm0aijI08KIVFqRbuT8jI+YsqtFd
H8vOl/6IU9sukTAgjZhJBG3YqNetOi1au2X4xukcuVBPVfGtNCtkvvZpQiKL
kkn2Jztt69Z8eBFhWREQ2jPG6xbmonYp4rNL+3acwsARsZuvcE7sbtlERiCE
XqmTTJ42jC6kdHVwI/71C0uC8YnqoIPqIDV+BsCzaZR4uk7b19lfbf7kPM80
onGs6KVJD09P5A7UNz2H4wRiTYoxTZe/D7l8ZLV1BWuaHHgAIP5DcoUBHnAh
CCbVoFvRPMg2hNM2kzd+rxJJHU4P5rImtZp7h7LV0xPYG81lp4TQAwQeGhd8
IIBFcUW4YM/9I6dYkq86waYf80CC6MrGTbqr3xHQr2fECMjuQFsravz3MIEy
39exuisXHcBvwPDkYTPuwHDlLP/L4JfRy8De9aI6fy2RsICkx81qeyasBNae
keLoMfmUjfd1D2R0hcfhtjYT9CZObT0AAnl4ezP1duHw7imOPRXXoZY6Gbtq
ooSw+QaVzOBX/Yw6FrXPXVOjUL8uTP2zQSP8saUqeMGazCQIP6yXO/f8s/Fo
Az30M6aaY6cMxtO3pDot7Tr3Qer23O+KnIJN3fSLks4wkavrD6Gm+z5sB/e3
x7qhH2OuVLJSPftYKhuuwnesL7GvdMFWab//GkQM09na3GcvkQTWrP3r7zLP
xsBT7wRpzLAMs2Ug25UKX2yfyCU5hXmDXeNy3L46GnfPG1sa9EsXz2+8dS4I
ddzOo/8nRXpve9S3ozoMhSlZb/TkEoJrls8rXWogUHdTZY3Bv6ElFbPm8Y5A
0/kIqCtJhFoTkd8l8xtNAnTQD5bKZ2Mc4HysOhRkjxYepn6/YZQ83kFrDwW+
vk7C9Uw/YDezgOJHTYieYPEg7jv9ISYH725o2zWFce/fVm/ATPxtnaUOkL95
xfM9uhRQDOIvcsT6G0JmeBkdl5lt26JxxynD2F+FnEJ8KtnaOwGU+j9fiu6U
UspxqR1g2vuinVyb8IxWA5UzRX7acxP3QRZjnKcyBLM8N9AD/KRmbmyXuBFn
6KfqMI+dXkTEyT/YeJJWpPdPzXTlqjt2BSW5jm/R+tjdpwRZcmNhFHWaxmUh
gaVnl4KiN/+wQau1RF7ZDgTO4nEaMQTXG8Ixuzxz04bj8ykMyLpu7QBI6ax3
R8JNzm9ibSrBnyjT0MyRLy5ULz9Zu2PWiCM0ESzls6He5MeYYPhFDG7tuO8d
iZM2skUCgQIuhNVCQPg5kO5mPQY5INOUka565SEIbWmC2dKFsiGM2JJjyNBG
8lj/Xs6dBHEMXrfW3cDAqQK5isLjbVBoCE8+gIjMXUD7/HnNiaC83EU2s+wW
oLmp1wdyFtbIfUG4lBeaZYeP1WsDxKZGVDsxInxSTJLedE5gDMnDtaxxoph1
9zByY3Xz9QQo3rf1dMja/5WNU+HYsR3vLDuVZtVcD58yaGjNNyGbAzhIg9ju
9vblGibsMZ1PLmlrPoLMCUCrewgbBo0JHPl3osUd2OuGeTylhTeqyUQ1WMy4
+bdhDjR/0gjO5oC6/sgRDshJf+JqqDJV6Ohzhe4S0X5dEnrXsdD6D2hjlIXN
k1bEXAobGtrmdJybcZlQGTSx7q9z5PNG6Z2b+ebU7n0NMFU4p01auLvh/cCM
LkCuDVZWmTrb8035acaSEnCNRvk/YDIir56dxnp/cdX0Xq1ppzKRxonnx4e8
bjm8HFLwxNihUUip4gL+JklHmeil173pHoDaCJ8L+ZI6rGAvDE182DNngT27
v1dRd9KkvB6q+lBC4hvk53Up3JCrvzckpzhc5iSGQPm7W+48k4wZXOqb5RNE
mRIuPN2G0ZzCa82iqFEDafFDujoCaYJTPYWM9ze9S9MQFUsPJYyl9zy/ck1v
4YXCdk16d9ouwnu7HvQzCXjwUwQM4808CZhDl5F0GeqvFgw3D+/f/5Nv4FXJ
0n0FMebqnHN+Cio/2mUXfHV+V8Kl4urkl3MB5/SKYw7ZNNiPNWe/yvYFxKGo
XVvPt+zs2Rc60e8BAcWzikOrN2eo5U3+TwcfxY+x2NnR7rTKf4/OIbrT1VjL
yIx6vjyD2A3wKHA2/5wZe8+DgUaTYJy3Ux4t6fmP44kqFxjwxWp4EM2TBNY3
2Al+lsMqdvblygqGLp0jCR7voqUhM4Xyz/oI4924PK2bT1Mslagy5glPgQK7
kcgMTUOlv3+OaMat1OiOSCLv2/a1kJIgSjGUr79EfsfEloVhcxrbLfGP+erq
4d6TsMaUGsDorTawDlpocfuxnlxSr/sfBnONn2gjsnjtN2h/Q8mHoNPeSRyT
fvB3U0f8yPUstz8QhPmeJwY97SSc2Llpr3x5VjmmrycBkVXkdjJbo5GL0kZr
SAmTJ6jmM1sboO/JK8Z7wojibO9NPBGh7jBX9KOVrcYUOZyBMvR3e8tX56GL
689Xr+IuY8OwSylWZ7aRxvOnr4wCYnWMR72iVJacI6/BO8DVF13aa4iCJZpn
dO9nYuCuqz3D8G1CH4tcrSU/DaaCRMjjlElBPX8jzVYgW7LO9M+Xq97JDANO
QT7Y3R2KwrPWAuoM0CyGadXPJFLGuILtd7kshCIwR74ckhmoSrySg4ROv5b7
GHBBqP/iBqTzYYl3MI5gy4kiuvVH/1dxM8BLJm6Bgt5tCGdeRgvc2gkO601q
M6zboLxNnAlliN6M89pgvn8MAiyk0GjLKRtUrZPO73ceOS40bdWaKLExTNh5
xXVpHlCpcU2Gt2SiWcK98Pgf91Dfdz0XaKgV+0B/yllEjLQp2HrSY1AtOWxT
tUgyNXRKYMU4LGkhw7akDGJV4TX0/KMeqT2ZlvRO2CdaBtNkVW+44QU3L4ha
bXO1Xf5FUVhoH4UTNz/pUda0TPkeVohEVRTl5hh/du/kT2AhuR5TzvwXXzRH
w16UCzC2klR8EkP0wunDNA+Ifd+y+Ta38bX0TBAmXp+h/9rm/lJDYAilftW4
Xp+EaAe7JF35H1ZNq1+3vtvl69JrP9AsImAQHsfN3kP7K58Gk97DRRrWChmE
3N+/fDiUTC+bLTaRT/jVb2FdNsi/v2CsqEiEo8XOqA41nyBvgh1MgWufn/gr
Df28X9URrYohMzU8xHjuYyO5m5Hazw2dksdimw03BVE2mRsLU7VpkdGgVr7S
/YpJ0k9E7T5M9OwFrKz8+0WYBE+KNAY4JAR40O9WCILbeI/uH+OJhHofXTn1
LaUXYJlUF3S2kAAjT+g2DL9nQCq9lhCYPishfNWszOyrqYMtcQdwwYqMi4Ya
eQ0FjVFF0N+RMNAapnohWkSFDQuHrw+nNSeLqTAvknkVZ4VrbKve5c1FfcCK
KOrXLa9PR5ZJ1eVbmqg2jpKQvVMFC4zfiaQAimMVJFKV46URYnlXy41RF6xB
g8sjMBaDiL9E43J5tf7DVKTJ1IhQVl2jEfdyY8g6BwQ1Lm4Uwf91HkwYrz/V
Q1Bb7WgUEstWJsMTdxEdIbciS2sr/euSE2fJL5pypKF/NxZq+VxQGHqkwHWU
iUxDoQ4g7wLvRa4FYKpjhfSoQhSoQtXgvxSu1c/qoAr1aZHcbY95WBbrpi/z
mUKUV+P9oWcoIWKcwA0fX3b9XehDUFGWQVbQ2X9kiTMJxW/HzG2BI4EeZeEx
TCKJZUHZjbPoUomm4XEuHFS514/y5r+kEaigo9k6zYrR/4LElReTr+PJeUhA
saygQ7xRKIjIgFR6oauAH7ahJZxcCvPUwMPaBhi7wbOCqQrDNTdkcl8xbk0R
G0p2fFUthAQJPa/fv/Q+cXAnoMBpQ/ZV04cfDr1QQEJYOaL7Edc8Mg7d/3xn
fAIe5hFOBr3goA4DGYLqKvYjRNJQ1xCzDBFutf6HDM3/D74Z7rn72YTsc+It
WAn7TZS3vyaN+q6Nz5rPA0C4mrCNGpyLuPU4JQFqiArOd9OMJT0vWApRTLrH
b7t0ZvPZ5ObVhZXTi4Z+LI87RXigaePy2bKi5lJP/ckpDnneCd1ByW8xYX/6
xeovgLCkph3vWF9o4t354pXmnocKdoaC+cSonno89a8G6ATsGOF0WBURLSvD
wuP9DqBb1eHWc7N/FACzWvBE+X2aURGEE3Oo4Rswi29U+Oxrvl12WpP1nH0q
6SZLV8MoyUiYehoEcp7x9VPxfX39tjeb5cG4Q0zcokk+qkAabqVNxJu5VH2r
+gUMRFcyiq6fA4JN43hT8E8CoKM0LCo+IsOAsdvmxD6uewm3WT5gU54Dqma1
YFwgMK/iK23qHMyyckq1Z5QzXq9loQVTD+QdfsFTSOVihIwuQZ5t+3AWFTDZ
W3xHmUwW8nNKK8hMUl6cXvjgOB+WCX5ZBkDgfLWc722JBlz/5pyCNIUJq0QZ
hf/ye+gV7tCGSTGQqezfdc7e+1O1oSBFeLAfS+pdhI6wWlFFAwUI/Q0Pyc4o
hoCRlVBy405B43Qlp86hSlyxfFV2jl8DVTPM9pvUpYGgKBXieoq5WO+sYgQt
JYbiIZ1e7BhWIZ31mSZ1IDw5N3wE8JLUDPogubFZByPFsMUwJDm8QfhOaBXl
0/3rMeTWK08wKJdurrp3c3W+6m7IdVF0IOF5bJH+zFcPGhOj1tjhGtqiQXFt
XV6FWDshUwsm17jIFWn1HRWTN4Crz8rThztlS12rIXbXUvZ/TpqEae9GZysF
RNtO5pz+7m++DlIrj0pd1DB4d6uWWS6uHwvbjs7T54uhny7vv2su1nO8rZin
5vKtKnYc50u6BcvfDkaPdHueu9Lw55wEs15192rSA9V1BZJzX2fn9iJk6KFn
P/gxQTNKRRMeWYJvjQEFf20lYtF4uc6yZJAizSimczT2LST8qFj5z/eUCClk
6iSJ6lsQUGcCk3seLpEKsEALdxjfPnBBWTyZ6ZAeQaMiywsHQEW/eN/oe3BM
6tM0W83ldYDAa8tdI10y7BdLAKR4XbTYTeLs1vZA6YOLfcXw6AcWylkZjZLl
MKEBEPzWSN/wAbGW8o0thf3erWM6b83hsZW5NqdBNds7prV4PrV8BB+EX+aT
Uq5q0XE4uDLkc7IBGulHgPJOxdiqlVeY28FrErrs+IZ7LdXwWwMZP6L5Jtpb
On3Cze1ST/B1cNmExUqMe0erd/S5KNlXq0yhWnNKbz3RgZfcNHV3UWRHvwZT
e38pM1p/BVVtgp2m/rs36NsEYQHWlfDEBadpEHI/98h0c8G+tAaur068nCV+
mWRo0IeZ2U0WIMJ4bx/QF0X+zarvkHBNmuuiyWefLJRZ6I7KcO/wh5dPFYic
pbfikwUR5fHJkvy8+wWwP/hKIOCQCuBZZAqY7bcNWHxnebOG9DqQwSAJsvsV
TUOIEqNtiB8XDNe27LM7D5PlkU/dkh8IP2iMG12B6ODjJoIw9J24GEaGVoPg
coWlirE7rH9xDUYjh0anzxcDuGkWTnEa5ingy27obxcf5FH2yIR+L2JKS0cH
OzJkiQtmIK8YLlgcQqeeycDvr8TT84dsWna0BN7gIlxXm91V4iFXQFopFXmN
G9/6G8a0na/2xE7/6uebF80kxaEAcwvxWa9ddXdz+KSuAd8adS1Ku6i4IWxz
tpKbs5s7q7e76GPAyxpYGccSYPwhlFOKjYRIY8mJYjNofMGzgM5CkfiMfj5V
zMSkSeOXcpHdQ8hk08quz8Og1tvXMQGUxabERnj1GmwMn6ut2uI3d8KzgSuW
55+hsjs+uV72aOxpBVKtrR+1ouQbcKvrvZwX5QboRfZf+8zWSLFEVr9L+xuA
t6uBURdAyxsOsfO2i+H4joQ8715EL1jlP2iIwd85MbDlFsyQl3G/tp3MAkTc
5+FF7pDcoxGhCt+n5jbf00QLwzBlTgPQRl8L+zqlN7DcLsi07ojg/MM2FoJr
4eFgBIO2lFe8UgdxUpE3mo+lOKEjZpgnqWosUxkvB0sKVAH0E+huc9PUumRd
hLjdaBXit9QGwLiu1boGpb2xB7484EY+jaOoYgN7A1Weof3gIb7wUvpzTs5R
P5FBkD/2aw3I788MBPKma1gwliRHl7CjgBsa2NUIBnyHDNfi/JF2UUcFaNem
hZdxfhMavR4zw518WCG9aN1vf0jcrE4BuUlu44F6PoLoWXGBTzKHojic4lNw
COZ/3i+VEaX6++x43MlpAH6645w91zmXIUuk9Y/Nelm/2SI/+7l0sRTe5rbi
tVeMWSztW1Gb+65OBS0QyheHsZEaLt37Yj8vNCiyVKwdUao1ab3ZJqo/XV/Z
46k0WvJmvcWmuRGPThMdVlfZUHC6ZiMpdw36DIv52B50yU5H28IbbAtRCTNZ
M15D1Arpf3+IJZ1Wze76M17lBfQUWmSX2BSovGVFVtHsRsDqdAFBxeuK9TCc
5Wl4nreW6QOUmxH5iY763uPHsexsg1ePC1FqT6UZ7GKlwHSQB4hEBkakRKse
E4PoAH5wTmm12GU8Vvfwn/V+eHXGmo9duo3D/IuQaSZ7PwyH1ltsX02dMsd8
K7RXQtuEUFPIwl8/L3tvtG81uBbyBRx26tjICI0TKS3J4Q8sHvsvQEOyOTmS
h1ZvIzmobzjpYS64eCjYieNxLasDbOclBsPSI44gZRrITzib46l6Foy/WxxY
8kfffoKSeMpTHA2IgFEzY2sGYUZEVUJdKUIfJdREnxtIIG3p/VY5vNyVEhOP
014nI7lWD9BK7sWqWVYTv4EChChyQwgDYDChlVetN7lEh8i7QQ6oR2VR2New
7X8L1uSYNbjX374ZIHNUNmfUBzXwiQI23GNzlDiyPzi9MKLktQBQwjI1air3
+X5P1jDwLUBBUYuJCVhAOyFdyZVbTuuJcq4yQNbWSK2AN7tULrr+orzuRy0g
b30msJYHWzbfvuCQ4XDhgONokh6H9z/s9U+WDdsoVn7joNF3v/Th8zrS0M9V
b+u/OPAkg5Pqlj9R4oXYdQ6yKyQMk3ZuFs7/0ZitnslAcsL+vq7qVX7LuM3T
9mpmqGCzd+/ngtRD1+8NO5/eorhcsAjnWgzfohz1jileTq3bZaNiY5VvPBGF
9Ps49Cg8zSHQnaSzOxcDFCXKT2tsmugyP20lFxP08YcXad3A3ZogvR75jqBf
U3C+FpP3c11DUCkoQd8dP/sw8/BWigMBoZFxjQjo9qCWu5DYc+zic22wMX3K
g+1+82o21uAeHS0T/UpLZvvT+HNWfLjfMIMjfOz7LdzujjAE8sBOVy6MLG6C
H99DbMRAXqTTcvRFIZG0jDqZIkeWe7L6SwuLU+woMGBXdb1VFkkw8Ggr9kG3
mVI5SL8Bbw0J7X5qxgBms/XLUuyygisUNB/UmegzF/b6bTjOY0FMdgAfhwTr
li22ClTwTFTUej5/yd+Mv5sEQ95Sfz/s9v9p4hXsulDm+oUS52JGMLe7BKZy
ANGVH+ZZ7pr3pTaTnep1fzXMjja1RRycv+B5stJT+zOdlOIvdzi+mwa1utIk
VfQue7RlV31xvVnCRuDYcog5ku4K3B+m3E1eYiBdU2cu6l6BqVD7V1k2qUDn
/+cfuh9q9EPChI0kk6NYarBvEHYj28223cOlkhmfvJJmam5mMJJLCKY5xPt9
KWg3Cr4gMOaRQUZJn8ASgT/vA4gwKpnPlHmqDEzKjVjQRoANDCGqPX+qlWYi
Me5ja2VJgcHMtmKW2pC+1lKkOd+dcj5Z6RPCDhBWBDAOkB4GSYCx3oAKSRIP
yZwmwbn/897wRPuaplqbc8g26ZokPUkwUrZZU0Obb3FpSiZnUWkBh/23Uc7a
f/AnXijqXTpzb18kiud2FUenYiuvn5AkEBve+Zcxp2/EFJpFFjMkndPlEHXe
tgG4S7WuYlsuUu347yUR9BD8EP+luZGcs9/9kRAGgSCRDrZQxTAVEhvl3A5H
bUv4B5Wwodm47Mf2Bnwf0P1MDkpfSjsI6K5KuYrwvVdZr0Hw9XKJKDjFmeYm
ZRGGPVeRGcYnocGcvAiOTPvtk1bWgvNTWQOeMz7i7Y6NRbgH7YYWlGXh73Ap
lMAnCExzqbVcOcii3lxq7/HDOFs/TB2yqBpNo/5xJ3pRWQOJuBbVzN/C2Apa
kTgJ3kxiOL6oZU2Y5zHP7artMky7Vy/gGu+ug0u5yrkk+8Y6cvOUvtbXejfG
DRcQcNWA2IDjEU+lg1gfv7Y9Hfv1NONitGIuiLMBYUFzWaZXx3DcHrUV0+sl
UtYc4Lb3BGtBaA187oUCPSZwMjixhPZEH7GwJAyvDbeKnsoqu1df8WyY1JVC
LzUfc9yEmEIbC/treJwGOihqEA6pD6wpQ7hjjDNSB3dudxsYLFxtJMpo/hdR
UwJwf0tuf8E6U8ZKVjzrFtvvOUZjeo7hcZaamtWCxJxZInbMyApWvdabWTE4
yOwnoaLWg3Ot7f3LbYsZVSa5BG51OziBeNbAun5WKJ31h5DF64OQAkheMMhe
5Sy2i5bO6hNry0K/3mddv6QWlP8tkGgnJjHeOuu32MgIQMy48WCtFYpAxdwH
ea+6shkXxkv/4hWFWKkA8Jhu+m1GHycVbxux5Vheu/L3QivlBkhhUCQm5R7A
n4FHFwlHcdGOpB9S0OgO+psDvstUHmGlaHCM39i+PXDn1DJ59R2uywXmdfkc
Jud/Fm5CnicHsb+Cay0CO0q+QZLfIMzMdre/PNEHcb1okRttv0wIFkAUXn15
VpHG6nW8ixJTCmXX7iKifObprWu8S/gY6+P8qsWQDpZm7fhePRpcM0yhos1y
FNa9Fvbm+g8v9B7kMuxO+5Yx+I6PRmRu20zm7gJCBeHzvAHRdLIeMjlV+Iqb
902Cau3qdvPnkc5sUOFQ2HE8nV1Kz26S0g9k3EQ+B7V9DF6B8id58ySMK7Y5
HflzgQhHgGRZMOOcabdoelSNODAAsXEoaaY9wuvioQSReYVpagCOyDEgAaog
oeNi4b4oP33ay3iqPA1wwbE2wPY5exs4EzQ98A8B+5A0oiTqxqzvTqtU+rwG
3JLP8QJNOZfwuA1F2iAO/An3rfgYVYCqJpcn9hcGJStdRMZecClqC2OSFZoN
a+w7dzx5gYQ389E6GiK0srGx14z2x1wSPC162XxQMIH5Gj5vqQsAeXF+rshH
2TMNmobuYiJmlaEkVaBByzuS/7nkoAkL9C/SWXVWBu7F2aaMrF2mAi+xnhqL
L++0YfeDlWpxcnkM911q4F43qUvEWKLVZjdsYHzePt7bImoGVMH7e9E+GlN1
QuBYAhwVs5Tcllav+41OwvNpxBAhgc2C3xvKYis1uUd17TgcoH5hIbFO+tq/
gO9m9RGyoiZEYWOXlBTpQWF4TKbTTY8vg6wv7jxUP5DBWTCBXNz8cwZzRBdX
Nt0p9WUWVSJEmlWBmHll+wwy5mbLtYw16eduLNaAgW9yrsXScU2zvc/Q8j+4
YXH94XTHB0mc+kqHhDA/vouSFriwtMoBIvXPr7pz3vgVpfe/Q+CaE5GoV7VZ
JegA/PH0aJfmKr/8X+jGStUAEE5ty7p0uYNvM5RCxcgd8ZBCx7iYiu8g88PC
8moL1fRo6HdfP8ysC37udwenkpOwb6VkmO+RxopDtPYx18nRaomTBGj4om9w
jAsw4S6OfDJ/+vIoMfVYoi7uFnkG/WcojMF/qr3yb87tMOUfoNGMIbwaxN9k
jVUes5QV6Q4/AxqLCFn30FRjjal7oKDilE/vcL5M0bUhUfwX34ghhkkib6ez
zSScgNBUMADBIu+CB2KRy0YKjgaV+08sMeMklCH9zoFyAg3WLmsAej8uRHTH
mOTi8T57P5KjdH9qYBlej1KdPIfzGQqu3TU8V6evfqF/rxMQ979QRVdO59i8
vNm7M0yicWosMPrB94Y0Pq9e1NGcEnQFrQ2TJk8m50xUSOTgAYmFPcqX73Zg
aUgoLzWPfIScredqcS5v42qs6lXl0k9Nwos/vZNPFs/XcchnVku205W3ZwlJ
4NNSHQOt9zjWnztNUUPzf2tM1n432b2pSUJmJw7ob9j+vYclHhaM3C5AeoQG
y5SPpt05BjJfLQx+KqwoyZJGH4/mahsELk4U1x8VFYVWJiDf5aTAUFJBLHE7
Q32MQbyC0jNHLUd71z+rEhcnPsehTmyxe1I853ohHpxS/TpwUc01XV3hXYe4
H1aPfCkDjSVg1N1YfIHQ3+3IZawST5mWSCmr5ZK5Qhe8YSoVLOErXFW1HoJH
+qE7BW/oL6GV+BDO9ADH0qf/1rNDqu20NZerf3fTREBQ458W3LguNYtmiNZT
H1cnZ8liKrTQHPBNBYLnZWQYjGNNJof92BvVIsULGE6KrsY6bKXzwsgm/l/r
rRkUmsWAQliltFEZ2qMUWoj/NWVch0uwkuL0w0VysqdG6GaTmGR4GUBQgkQI
V/JacoT6fTXEaFnYByIgEpfyQxW8uj2Tiid6r2i2R7lPJOelkcP8eYXnd4m1
zRfuGnH8V4w2X+IMWx08MAhmlruTTmglrpiqatI6xvfGrQespO5KhhET6BZo
/M/mwdLCwA9SDUKyjpM8dA/IV03eLyWXKuqZDvFrEkGMkg+UqEqT41OP/dxF
Yy+SKAgyyQ+5Dwdb/OVyvErg3HXr0sRzM32QEZRFXCZHVioU0Z2WNu5Iq719
+W7qvUASlz4+dWb8KK6w4UwHlIuaJSuDVPbVNeDJn/tmnl6x0xcBbPx2n+3f
vIFo7HC9Xf8RF0eYQlh8r5ojmeERtWiTJY4i/U4N/T3DiGT9N3kntbptwEFJ
v51Nvkt7+LGP0jLXZ7i7pYScy/EqLwzqyGkGFMv3VSAIg3LbomFG4W+OABpq
+q9hsgH8YbEeoJ7YNbCu6/apHLYAVdMbDZZI9RnQ/bRUo1qH1HlQRbYty4yH
BI+UeeQyJgpWxkPKbln5qhJHjID27KfZF1uI5Wzbxaok8ch+Q12LcZgSdxSC
NKMwcV+thgCkZ59Qzv9YJ9HRhZmYWoPbx6/jS9VlNlzcsLEdvA6niYonF9d4
tQ5zdqBE37hsc7o1aTxumVjJ7UjJdpN4orxEB+PlSzqoR59+rUYF/RTB0yk3
Y6QxAFGBQgToDNQgaCJs3XM2lq3kcbgvNmH8CkLtHiKYlpJ8CNII+EunpD5D
upes19dg45HCYnjfjMztjqN5PpTJmB4bMStyQmmJRIp9KTAHGfSxTxx5nayD
GOPfU+dBHlNaWNAz+RBB3Yvslhlq0HStcCBoYo1tfS0rujL1O2CKj2+EiHSE
Zq7iJi7YWegdrA6kZxkze2kiN6keBSyRlavKzeW0Yx039SiDpkyY/OOcqaRM
mhdrx/vWctLjl/5iy9NdivqR/GrjvJ7nbrx0KyMVE6l8UKn3R981JTx5jbcj
e1/uMlhyC0Ao7IbeSnieoYo1U9MVw1oeppX9dKQgMrVpWYqD45fpg7Q+DWNT
mUzsEyn7UnbIRKofe0cCX2/cv8I36Z+/xbR53jQAX5OrYN8u/TyLpu6JGuoP
MwiUYCjPIwwh+X05YSZB4V57etktQEkGB+PtvDUPWAfyZ9pBaKy2/uXlHVj6
cCNnJx568SJ9yR1Z/8E0FlFvHaANbXGIcO7CGH8ke6Sk9YIcx0EDef9QO0fQ
vWUF4vHhrOlgCJ9X1piiPG27Ryw+WBJ/KoGU9HkVT7daoYOiW/9TTFTEVIki
8fP3VqFgB0s66SUXAW5b6zCiyXho60mc1DXP8l5Vk4BAvwjKY/3KiH7olrd9
N8e8GvUQ6oQizKGEw1r/BPzJGPg0gML7Yom5E/ST3NjFwhXB6chdRiAdRPAG
H6RKgxX5CQDGDa1jCHjLYj2fdiBF48heaCkLiLyIxDpQfaXZVQch6IGV9Jn3
ckHjismatBZsYwf6BeV+Vb7gjsgsY8rKQcHRczTGna41C+HV+BCcTE4he2AV
ud4H+AI+BFHhSgTe4PZ34Uwgms/1lezw6Zvs162ve28CzfznJjS0XNQgSq/q
hvCYXY2lPwEp0U/Cnqk0MBbQtc/5cEhk6LXvoub9keaMMWLhN833GJN3e7MD
yewRGu+dcZjmDXyZl7+yvfpacvatTi9MA78iIuPeAqpSWGnzszl09ADvw31+
qMHtEOTdMcpTf7sdyoQMFpmaqMCNNtnAppwS5yhMdEiC+jPLVjrY2bW5ETEm
qFg2UCr5kJAzBHy566e/z5ZH474d7SbaroCzlihyJB4RxEpJA5AAuSuSkL1f
7Qqq1TxXXOOkuLt5CpyrvMffQ+ZkgZDN7U/J9PbLk6kDw3nbhwsqJLLcfhra
VX0OsHQizXHwE6rb9BP652R8RZHr844y0HvMwvcyPZ6MQpgdj5F8wMdRfTQe
dx4o6Hmrk5pjyDQgo6rxzNP1ZGbeOC7qL1dK+44ay8ZCEPZ8vUyzJ9/Gd6Do
bJX7PDjS7NsZwEcZLzA8ERW/lDKO5YtZelTYph1l3Y/TLOQ7AIC0JoDIak0w
Y2ZDakZSi133ZKBvsok8UTi6tyraausfOMikzXjkXe4+zcL9dSnhIGc/QSR4
YABMgQuL35U52q+RisDMjZ6APH1rMrpPQ99Ms9j+IO2t/WXkk3I5YbE0Na6I
xzANOaC4P9GpsRmsFtITJfiAuAxNfKu01gOmbUm3lZCzDUm548tbXpHLAwLM
06wiW2RSkaSDU0xdzF1bY+SXYLEXLZI/Rv4Br1c/XR7RkrtqWg/qa8Fqz8XT
7rjt1xgP3u3JcTk8iS7Evv9PvmzoYxCTxuFty41y8lThzv+Ato4eAZsXiCcN
zTSuNUnktPqz6kWQOr67cOmH2LKwBUlA4QD1MxtsNf10BLMOILY3IuZTL3wC
BPmaD9euqVbEvigWETt7ATIhYeclphAwzKNUjJy+3Yo0damw1YKBNZ+rwsnz
B65Rqc2Fm8sAqE+EInzzpHGJp6HtitDXHWBK54iWlhF69unS7DOkjH29VgDG
ahVdSZ76bsD7zQAI9PUQgBsYkHPju94KvBiHKA9pQJ/AXm0KMW/9BR8xPbDv
Q4ozOS5gJfuyHo/TEtwSQNx/v5EKuq+nwb8VrrQKy+p76pJqjMDVC0IK0snd
yjnVQlepGweJcIKJKV20WftyP9K/68/05lCUfSxWgI3BHIPo0OLhhO+16CgA
Z0YxnxtP8DVE7fiCL4KuJ1iEE6KOscN+BNDqlGEoz3ubMM4T8VqiChSBGCL2
e5ZBG2uvHfonjARAk1dXYMJNmnLr5r0XpDGeUfBPEvujK7ptSTc/wSX2xBK5
rUKEE0AZlPuGSPNn4UfFgxuc+yRC+AtJON7ZxDmss4z73k68FNtVvN4yAnpQ
LkqICoHPAX/EsPw5ezGEfDrD/ptzJJmX2UCf76xgUvdWudjrQFAIVui84ERL
2MSXXOM4MnggUGofctGbEhmOuYsbIL4EAMbrMuVNAuaIe8yegOcbsSXPW7Cr
yJ3Ejoh0t+CNZOv9vMWOJIfG2FAwdiivMvwxnSRG9JXyyO9OFC3WokMK3/jO
NQhYKCmtc5O1uVqHYeAFuaaaUK5BImyDtMc7igyNmD2fjyWK1iMw/KuisBXn
x3cQjhXZGTR8C2DFJGsLnsWbAQqBTwwm7ylO5VYTcYnXoXsGQGE7Xgqcv9Ug
r6f4Y4VTMMnnXUktpRHlt5hrZ7EQuU3Sn0lh/1U6jsfeMrggnubawJGZxHrS
wuOWh6PIcQm42o+2YC0fPHLnrC1VzZ9ltELlNAr2Rqhn55wETxrjz1JxF798
2H7c6lbuRTkA9UglD0pFuovNoxyGeyQAnw9sa0SuBWajGTIz1bCkQN3o3oZ3
Q2rnH4ifuHYQhWxox4+OrDYHd/00y7wJn67vWqq5rGgZs34n8+Q4I1SMUzBF
uasOqUq5F15h/qwed0/kGdefi8CCFfO27/PVz+gPAsyDtZLMJnYWKKrlgxmC
yZtmLb+FaaDeYANNZb7RfQg+jBUENSVFcRZ2rSEkcUHgNFnZYKoyWKG0X14c
FayYzj2Z8TPOS9mkn8LGS7uI0dusy8ilEa2MKqbwWlpBNOLEHl9V7QfmFrp4
ACCuLBbsbqejsOmKr77W6TBlIYOQgeWSMAyBQ2sXDdKV1Nh0PuUOJHnGgrDZ
XDKfG0LTx7ZcsSGh682jqL5hf7QE5ErBkIQEqWG3nGBkXCyODmr1WYMXlxgY
9MPanDcjql+Xwr49/oekAHw3HOTEg53zhjt8u1HwqxPCzSbWw0Kc8eN3Fn47
7gIdIygehENbGF3fcZp36vmnvqgat4nCp9Pip+VWOrek1WO14x9kk3Xknt1I
blUHKJyT5XsPc9VF4VQ9lps50jL9zt4hUdtjOq8XrrGhBPDMkmiwsaPd6zkd
MevqtV92sCNokCgvTkjan3KUaIwwOLxOGIO6Z4aOHXRgDlQnK9wJukadwItp
aA+1qKEnS387M5iWCZq5bhWsIycfeU5Fz6iFnCFry1ZLgliEClAo4oA0V0M+
fz3QI7lwMPXdPDYdrm1I/FTtO4nMCsu5SXe9BcMSQZ9RCgF4s5F8Py+CQg1h
vTXYLRi2bAJAyr9DGjwEeZnZgr1Who3xoBlstdFCVRpv1xipqOVTiJJXihIR
qJBRNsC97B/mx9aH28o2UiAvYC9dCGp6vzUekGLNLX8j1hWWSchlARr69eOK
EvE24TNyFHWCe24wkO9YqXcnuiWkl2DdFV+Ev4rFjJVcHM5fx6kH+1ao4hxy
l1lDTxohaS3ImpyPTCZBugaTRAaTmGXPrbfV5THUR7LKMTF4DS5rULhV5PLX
nGERSAol1LZav0pnhc9vwlu0AVhSr6Y26Se5fX38EHqi+cJyMwg7WoNUwTHY
B7Q613UcYrJVryJPfkqygCcMny4RpGyxjyQUuyohaeGRyGr1G1Y4AtH++rXH
4R3FdxHC5W4SZ1p/dOlg9lrY7RhgW+j7PQTXlVh/1wj+mD/HaVnTzNb6f+TP
FPjpIQaD8tnh/TiM+Go0wNUk4zhmb3vx1eFn9AfUffS7ERyQ1SGugNSzKWd8
Nk3FQcpTWrv+eyfWOQUHQhbnSp6Lic4N6SHZUisVzE/Bc3lYzA/g63jdsSkr
AYauB5utTvp2rdlSsnszoTKAU5urK+OD+1Hlf692gT8vt1rKHd4QM4Rjkfzh
P3Cg8SMoMzDfRRbpgX3SJQ093SVUJ47pecgremtkO56sqHuxINKP9H2BVmUo
PJdUqNmsLLc64980g4vpIv5fmWWYblm/e2RrB53DacRQ7uvunB7QrXEGVZP0
heiW56WGeiLMTQN4U2ViA0SntzTm6yk7TS1n60BNMgBtM2/u9AnjCw/0MYsr
3nQ+INSm4ykjJyZgavi3pXshC0xm+/7paJldtVfnITHAfhNF3iLeiC9QXUAt
9wxXA/As2866vch+xNtjnTy9NBBrbP/kWttmPIgqRd46hFP2K30W7PUt5sRl
2lLOzOA4Yj3JU5mH5kbXAtTkg0vXtdkniacjeZ24MN1tlFU2mCSLD/A024oD
LuaHYdzn44eXPx20+LNBv/b2/iT6HCshwR7tN07nv4bOv8XgApLHicCS7+jI
EhyMsb5/RW2qX66xbb59V7mQZMccsS3X7oGDzljkexeen0k+8PwgqKCBpyPo
Wex0GS5S6htQ75SRcO31e+AKP3rkTuVi6Tqe2+VpnWv0dwh4PTT3bYx64Sw1
JesrVyhYc4MfW4DYRTWlO1QY5Jz14vngQ3j6P9EFnPWCKYABE+CENZEdfJ9P
MJMD4BDTr+fAMoztE5AFgcZ0Dmqz2xVwSBiwPFPRuVfQE4pG2GVm4MDYKhKt
A/6a0ZGUtcnv3yazNHVKqKTGePp4RQY4/inrbxMnuKDwwlTYl3G7/rnE3T94
OJsF/nkEB6/w6lssJkqgM2eBAtYchx2kOP/z7yj9gxNsfqJB9mVVRjSsE2vG
vV81TTRbm1dIhdbXgd5pcqq8Ko81IfX6x4ML1BMLguEtMmIcopW9wmeWemDa
KlJk8Gcsg/LfqrGGRfSPBJcdstjKnMY46Rt8NtMXK/xtFESFW5uoiK02jmBA
3qDgPAkIlW+Az4tovx65Lcdcq3xuXs+3nqyebjHzMBY0HwgUm2wFCsco0/Ga
iGwUH6GfPRxVBp9z1MZ5kE5NmPGUiUvV70Te/lbuvQ9zHcOD8uHgF9UhbMdf
e1TqvpABYpccB6UWkQK8Oh9+Bhz8qi+43wO9WW+bai7/LkmkS1Vfc179fR8c
Zew6bWsSl5lfzKqqSV61yfwpHIPwOjLRIrV9nh3OI3qDsLPgVVfEUEjjjP3e
N73gwLHa6/P12UUrjGCfAU+k0K0sCh+wSqxleWardopmIEiKok/Lyoqc7hMP
8Wt6jTIbwzPCuCVx4yYOxSBwlBuWY5mKegs3iLcIyrnQw0F5zbB7ycOuCy8i
4P3Psb6Wu/pVS8kQ4b4O3Ced4lIGkWpo2BAt8DkmYUBSVtJZvv7xXvoN+ivx
QlHdPAKF3ZEOG3rPfCDxWcrPt692Li0VgXhXxcHwP0wjCfhpYUkZkBkX8xYv
zQJydkiRqZiw4G7UOS50ZEd/WuyKfRFmiT5xaimAuDrSYNOEKjSEchjd4yR9
CZ3Ma7ep2DOIB1KlrCDn1y2scqXxSTJc06Vr9LAcnDgNGjiORT3cfq9d3B8s
Yi2x/wOsTymi3HTW8wJqQEiy7+oAEyCeJmiuPhcOsN8atpVf7WR0ASZ/jZpY
e3KaKixWLm0Gk/jp1pfbYAKWLia58F925pxQp24BC+vwmIiv6auwljDldewS
papyD9APUbYWEE6ii14PqUS4s6MmrszJX1dsb7WXaSKsgTvflxJUMuQEuuoU
xND07m8/hlDrGnyK/g9Hn1VeN5KNV+Z9xSmIxqz5Lj4/HyOqTxza0drOQXLR
Hnmbt74NvNaeoyxGeoRfaTYsuQMsJK2mGj7orOzr8aYlU2DlugHw6eyTa9xA
EotTrIq5bWRVSxvwGpzZFcOZbcg7mr0GyIIJgUnz4hC1znF0NWI1p+n4OhGo
bOyVx+5HVe6AaT5mB3hx/bLs3edFJ7gol/vEMuORcUFa6NPwZm65VKmBGOrV
HtsJQAmSYwiSRfL+ZAoblXhapy87H2HxufjJENp+kht8YHBb4X9vc1iq2x7R
itMHp4lVTJMWr8QNVF26ZC58r72jqQ1rIUgYCiRHUWzCGs4ptdhWWzGMN8sH
BEOP+jVTBQljxpIS9kmXGUX0kLv+DeJ0M1yP3FerX7vCp/tvewm4fSl7K5je
UEP7aXL5ngxj4pD3uaZmFyqRUxm00m91SDfRF8BAKZbbOtrzNeXy9f6aF1qV
V/NxeU5YTvuESEjS+dLSp3mOUCzFqclJqC7HaG5uWgAErd/q0zXrFces1mD8
TN255l/2SjW6CNDqVNWDmXUKU6uhKYlm3OF9yHxAKDUDoj5TotLPqyQaqPnM
o/uWy6JM8Xu9C/kkPVRfuJL0tdLMjJ5wKHOE0j387Za6PNoCAvFNv+tUBknq
jVfGifCYPG8fvXp/rJS/k+RLL8SsPvR1ZQcVH+1ohPeeL+N6sPgcNCBf/V/Z
vHLU6EVRlBwd5+JVlHa/halKik6ZfmZz3rN7hAxdN67nmthjVSwNVBD5bvVN
9h8Wi5mM6GaBg2MA/5WXIZyMQsraj1fDFMAzh143yMtvLtK3WMWjtjyn0r/M
KqoZAerBu/Ne/tfxq53i62u27wBkElR2SqbbS1a9I5WKgRWto08Hz1DWefq/
EhGlwuXz3tfiyUJ7mrDQbwn6taTzDyh4abLuzHbw3MB8/UjwRzSC9VSJz6EC
c6seAv3lMfwNE3wDOLVhWAUJr1Ft+nT6T2a5d8lN+qX3KS3BaWp3il48ch89
1E8suYigjJoiLDoUMyP+kD0mv8QY7fbVWuOVBjgLlJ0MXnkxmplBSIFmYuXZ
ENndVgzrHpvj2hQv+1/b5RDpRrmM7C1grGHDErxd4e+ICmyqOGCaHrYLJmov
zFRabvlZZwdU1bL/9fAzZWmzSOxMy0U5EfjO8nRId5DBAzkB+XDng/MHzqtA
IwVTdUU3yMRAmB252Vw8cc/evDVwMNLjcwFsQt8/J9CISE1QfmEDxBhkVKXf
uq2ijtCPORdeFHHFe+tEjASQkA/1tKN3PlkQgBxRcA+Z36z+HD4QfqxY9sxu
in4dHg/O1kbMaNhAW8HbDexMbkFh7o8nB7UGUU/wVajRPiG9lmF4Ksb0uhUo
rjFPcJ4SVgMrwoGfhTeP8X72WqnJAJlfhNzhqvcPBzgfWVOMRC+8DG+ogCTm
Mv+TKevlJDHEjFKzVAj0gQkrPvpyy5I0X8JhaKWuEGMt5SDE7w4D+apb13Z4
7c83mSXxvG8pk2McQ48vmn1w7DvuJ3ECB7VYw0uMsvjOQ4SOPFx+ONxbV8qm
vRER7cdkqFt5G/y/gIovuWuaWDWuj8uKIQ7AbOcQjbhCVG8HNA165PqF+Rf6
g4kqxS/eYuuWsnnkUkXrhKs6Hb9niLSr429B7hTfT9IeEzr/pRm0L4SeI+61
GSafYsP1hdvXvuPHqMWOqB8Oi4hWNze5vFlmkn/HymybovVzge8vP/Wd1Cqf
up3mFEvX6pwiyhfXPOWnHt9W1WkwAmgKousLvqk2L1nlgYzlAQuAqQMD4TTf
/8m1h6qNcdrfOEReqdwVTqMT2YmwAr8zwBv+vp4Q5g6vURgCzHKyxmgKKw8z
9hC1f+vMNJKHAO7QHvRNKIHHreVyqsrYf5lEpmoqgjSxEInOaVcbh5w3Vn37
jaXWDVkoiYnw7Bx1lb77swVLn8v/HFJhgznie6SdxlQYXAa98fcvehDCy8PQ
0T6rYi4pGJy7nE/hfn5X0avYn5tTxlRd2+gosyh3g67sDQAsOfz/Gh4rIxPd
TX9sz78FEZRcYhecytR2qwrMW9kqmWWQdy77GpZP7RnHjMbLUdwMrPS1U+em
mVfpx2PU3Pzm9mF2nQxsSV/RG+CYxn5fahc5/ExNiT7sR89KXxg0M8RCR2jL
JzqdasoTkh5j1oVBnWEbDQxozvF8AxdggaL+DdkXrjBncth2necg9qKgTPRs
kKeQkGWwSvWyG/Yi5pdFDIA1Lz3Eh3WKTDSLaGK4UqIJOOgvPQvF+7Ybd2kY
Oxk77y/nDhvFhnMDfUlADfjHs95X/fNoBQH0gsMLu6kUF90fTtjzDPI/9Kz4
uYHMy1ITEJ3HRCbpyV36mMDDILcNH5Ju7jZ6fyRgjphOkMurswZgTRosKg2u
IVMEmmMOAjMuzJGoVcZY3VV1NsoTpKSWYTajvxLDBccg2kKKOi6Dw/ihQ8hb
5qSNLYBmtfJoq1AwQ40QPSk4UocQHe8Jw2NRk5eBy6/pCHPqc+jcaOQAdpUA
qpTOYgZPWomMv+2yuPBnOdPj5LPBayCFgFiU4i29xWXav9Y+nHZu2gTPPPTk
vPhESVJ9dc7Pj2lW1KhDrB2HG5gcDFfAKUo3Rpo8+p5IWbDaFkMyIBQ7/sIh
Jta6M8j/4R/ftOGZ3bZ6WKMTzNXgweD3OBGgaT/vqaPqN/0IqLh2Wy9vmoLe
KaVZs2pbxrwtK7Vatqe9taPNfuzpcvaGbMFXb5Atm3N8SgkszaJSKcploHA4
XMjUKzMh7XLWLmddJDngCUWkxZLkZNlWm7FnoahIo73EkkKI272HTwgeIlz6
ve/z8b39qB4xcu3jNRty/qvwHxfiqJK/Bii2KwPctPTHLs1J8ij8HdOhA8L4
lj9tz5XWwA6H3kQO5jqeWyhvyMzRPsUfap3opN7QqqTuzCiidFncJ0wJHIAU
In4FDSBDhhNpfI3BP7zs7fDwpsef8ATg64jx8/lbnqj5OG2OL3iPMwzCSsyX
m231lNQFzaY/TL106Xpa7/5GWF9We9sGPnoCHdIwsXhFapHRZ3eNzHgJeJUv
Rw1fcLmlpMCzlezDfQM8sRaRrTSGqYc71kPGgrWzajSOCUjEhPzGFMf1qTbD
IFUFdhqRmpg1MeH1xzckxK5u8Fr+4T1a1LfgmkPW4C28nEUNxzSHISyqw8SK
2m6fe8RGsDHouv0wFMZcYYTLZy0Uxu7I1AdN3+e1zf1SFImoWL09Y3Ojs2pX
wMyNNgirqgEC+MAbRRqq7+tOMtep1m5S49gcnGjFI6SGExvqcRzhcHPQArIe
FhbzQ0gQ1/Qtpin4iCWcMe/yJjKJWWeA0jzbEar3gFSQGKSVlGGxYL4s2hby
HU/BUakx+Kq3CKWYVJv1fiN1Jc+NvXJKb+DR11Ip6CqS9WeAjWvINuDDsBEL
U1QCHaX/jIzwCRPqDhPBej0Y9xm2SAPcHcflcBdbfR9a3JL6HM75YZnchu+n
pQxaLftOvRAE8bV+QNl1j+sTFpIUeU4KQk9iB+TPXVgqcabTg4QZlPahq4b0
09lvTeVJwwitpL+NsZsg3Xh+Txg9pB4Hf+I7pfIx5aUhPo9m+O8W1sS+8HDs
WoizjupOcr5HaRpYL5puc8L/vyCZGpqpRu/XGfhJqKY3l7X9fy3xoaRuywnt
MUJ1G1mhifKQiT1ZqRlbnIRMsx4NLiI0VqAolv2Ulwioh0SvLjxksUkoi9Fv
68v5l2UW6BIT/qrWWjYyie85IRChOF8OYGR4Wr90l8JtnnzsTwC/KHXNxhil
7iK0TEJY7R325uIw5vkKGtSx6J/2cj8U097sdc74YNaXIwZUUR/pB31f6+iE
OBDIpDUpvXNPfchyKjV3S54jWTlGYKdkRF81AbMeNwShtUW1C9g00j2e+6R9
5CAM1/JhPpEXPqAS/OQzDeQ8gyd6yIMewJ48lS+zE0VSOgzzBWW87TXXexy4
3tW6ViYHLDu8nkdlw/6vAVOfoPEoDsTelvRovBBhEXeILGq20u907jlu4Syq
Fpr1aChUDVy4ismFSiOq4CGZnLPe++3lW4lqFU6b1NvA9POGXgJaXsNAOhFB
ciubE+0JimTQ+lzfaUmZ5W8QqBVo5Qq7OGs4tZd8JLSaPOI5NKALCtYGukPi
i/fp8O6gEkAdd7ZiC4q5SfoQRlD3XisCwWg8GNDVX9bkXzd/vxsxqAHujlG0
+U5N/Qg1UBDG+Ns8Q+8aCpB8a/tKRCVXR6W2aeMujyYJ3iIcJhmmaHcXSP3y
FhDAiDSwgvqIb5zKcOVn9ZHdTmVIBLe1Dw0Bi7+lSFsDUbdZdIq+Z2oqrqGS
qETmcFi5q2600sj7GJbbPmUsIGxnkY8q6GGC5azEpCK9ABX20SG2oDMtrtCE
AyoelifgwkhkxoQ/H/jKgGgwdcmdaJNuJp+mGadovDnmUMT4mGaw/fjgo+PR
2sNc4qrPgL3d5KVxLcQTdi0yJ7+mWZSCoGAEadN7FlR657NUcBiMacg2kOlx
nP4YBTJ4Ubi1S1lZCgKHBv7TN5t9jtR4TOFu7tG0sqE/2vFfbiBFhxEeLX2U
LV1psgnA+HszIBr6zBffFJRpx1hdImOWnt3cwT8YLNcgObPnJISCsy1AqvI8
m3IS2iu5FhRS0LpzPG9yqXq+h5wJE6wG4Q99jNixQ4sUcpEzImDeT51OfSOQ
HVubkMBmKtxpcNaaaR6mpmVpFyLds9GPfxISORzFee63y6erQouWNp1LJ48D
ay9ML6qCj0MemvWdhfkuGoGOXoKLevmhYiDlp6yWatitkPGXKMMRg19NBrZz
AjFOAC9E4jwISkK4L4o6lCpMnMVFrOKSZQ5UArFhc7VEF7uDDXG/N5pPZamY
zTJrl4sGPxEr2szHiua8da0ns+GDBx6bAdg5uK9BQri+BxB4h7VckbwTfABC
I+trf+Oydc5foGmj9jDh5jucMSS3F7QqvM085W3/oTx5SWbIhclbw/ZeV05x
PA0iPQN75/z8aHy8yoWkD/BwV2WDWFI3qpo+iqkvO18mhBh2I3QyiMC7C1Pm
+aU0Pv5TnlcvJ0UIZDLzeRvSS0VOT7LI3Hqhvdr04EfVZp9okpRfnAPeVR0H
bgNWohcfAiuW5neKJK44MDTmc+TvAPkBQ9C3hinbq3wQj03g1ctprzjqQxI5
cmTgQq6vjxoA9eud2wkY1yajlI3ncdzkqLd1o0qhkFmCV/R+ZSrEHQIi3D8z
h39tQtgPIZvl4wiHDvIxdGuTQFrlgEf/DeP/WAu6AOi3PwdlD0zkOgsqf+X7
zvvWbrUPt8LuLhDyB0zWdlgIrHvAWCO5+EIDiBLMbkMG4Q9u2Vq36R2F5MYi
cLmwyytS9omWefbkcUlKohsesuz9XSMNLHmnDfXD2sYm8nfEeNL7KWyM2ycG
2uy0L01pvyriii7P4C5ODPUGro/Ave1tYGRM8A5FOyq+wonl+cU+ctCzpATF
S/1bTVzpxj8ROB/8DcErLC3dj8SYlbbIeOaTgzeaChXD9r97P8O1myi9edcZ
HeFNXlMteaG0yDG1iInTVxxQED5P4zTFejmaM4hDdcuz08+cooAYIpKNRxj/
Nz59rmoReCNRRJv01c6QmD2sX/uW64H0kswHgais0D8EZ8i87rXHHbybWr7j
NRmNQG7eofB/mA81vdjMLEzfLfGrwQJSg2/wCJKO/V0GHLXBb3ML+rJJPIqJ
goI0ZjuzKCTsm0XPM8rmO+vMeKEFstOg9iqm0ICMJOMp6qSbT2xAvlI/n5zU
Slg78KQ1WF1BpmXfIvFYXsO66y6u59edcsLqkrJ9NXJAA+SvzTt5XvbsmviV
JKv7A95ffOOmsSHyZNtNsA88C4JvHMmjUWX603xqBin5r0JDePLlr3HarvUi
CA1ZKptyIgTzxAk9FlNdcoFhjIyqQUfhU4QarCB9T1Ks+j4fHmfEwkj8/blE
D5VpAZe0mxtGBtg87DP6nxMNVRtcGj2ciJH/OQV6R1yE1uLnTN+oOm4Q9HGI
4jFiT8ijgsVEnlm9Ie1jAKJZqTGJR1SeG/cFpvsmo7dBJntYKwb1mEH2zc27
ySZeFJqyyzSRsPUTsurdhv9zsGQO0awElqWqZcYDty0UxgSziUjvFg5uJuIG
n4kCtrJYys5z1w7cWM58284qD27Nrr/1KdhM48SLc+JwWG2DdmAi45nDUR19
mSoA6dA2Ih1oBbTK4qQeHoJql5RXAN6iBMZZ+bvnKBGChdTVajKILVLQq2W8
omwhfg9LIz0NlcC0ji9flLsnR6nYq1Ky+nHfAq/vAwz+cEXcyuv77FwKCjIv
m4AZCCVGwW90JCKCqP0kBfvgVjbQn0mAw54cbzPvKmmo1eYdsv+gQqHyTJZk
NRsGJs/ThJ3ZUF2+xp1AeiLwoxOclla9H6p0Ce5ckDnN/n3Hzv7zWMGjFR/T
B2GEfaeFqhvwiP1BrdQuMOBpcQzyNSJ1AmohSbk/ax0M8Xser+FmBRuYhgiW
H5+L0RtgJuSq4J/AHv0U+aUtcagAhZbIKB/ZaC7XVrc43EoThagtj6KF+gpV
Wq5jHan32/TiVBui7JmNCqj31kCKsvcfwcNcyQgp+REzf5PHArMdcH1VF4VH
EYd8aY7G4AC6OZ/FeOp5Da0MVru1hcCIz4EBxDOzMZwkhn2QP21N9O/ht/FQ
y/YAkNriIsehHa8vMfob8SWYMoX5IjTZWoqMzQH+BcL/NGxNwXCrUmxFh5jZ
rayhjSenNrHhnKu4VfUiZr6ccafPi64OcI3XMs40LHllG0hMEZv283xiMpoz
1dkjcGiqoslAYZBZDI3UyW/Tu1H+q50Lt7/7HUrKlqRZ5gicBaG2cdGgbucB
SMN1dI7xjxmDhRb5B4cuqqB60CHxf7GmG7VhBjo8hS0a7u0jw1RStTtEGpih
nQZXLdxgDSt6FDtKEF2uTGLqgaDcwNfjoxy13IEAFyiw/4OMJnhyFRdEhX7I
ctNBXED1ckQXOdebHetuLE+yw/Zrjc9sFGeztwmQxu0h1gqY2YSXhdROBPEu
VSFkJWS4DkJKbNUSs3dZWM0UuyUK7FD8Mkn0GQ5WVcyianqbR4hqpzci+8dw
EpJNRh1i8RBaubq/omy/yAPJhzkZpPCeuPrQBV7wPfhziP4+tzF1+vaRh9h3
LNbKcwWxgQSx7MZNnSXIApe2siDr0/PzV7bGSWdfDHtCgT0/I1RgUVtQJz7B
FDfFQ41ChKu708W5fQPDH11/bWQ0sF58OlnHWOwNQGE62KkPCZKJZ2LGYU4u
RU/Dnm71rX8ah/O9ajwPeyxXds4zimIh+1erqQx1aNxjGlIgyu7lZk67BRF8
pnf+mJrHHtqnOVXh6opt/WUlbJ0GYKPS6pxP/FlDPy2EBzi0WBHV+Thytdyo
8SrLzei1Q35FDXSn49YbwrUqodBDomcEfTFg5m/KMydfLjSm/Jsr227DX1Of
lpc+fAUDg23Psr0oxe6lQ4wfLzIz4BJ4oYku9+Art6t45muwzws8G5KzBrr4
3i5R2kTW2v8NbKPa+Jz4XhZc67T0CIzCd+c13YXWOQCEZeWfVeRlBZAXLsfl
c80CFkcH2GWGE7/2Zl9X/tDqrA6oIybEiOhv+ahORvdKLW1jRRN4DS1BnN/C
nW4XCr37AF13CAIITkUP4GKydMPqyjKzRW+NvSdbMNWY0pYqMPEorMAVMIvs
vSj+eq4yKtDQU33OggoPl8X3QBkYEFNx0crsXU0gYHdMeMdk36enn1iThzMJ
N3X3Z5sxPQhVgCA9hGAWGGusQYpXJQAJIMGjv1YpEswhnU5c2ZyL17yf5ca1
sqXQ7ya3DG+VXPhOyn2PXAEOOoPAJfqWM1XXGLfqb2WTmAXBnRQ+h9Q5f8P4
E7b1obD3IpvN7iPVWhKKEPNpmv01VA+tgzs/8qz208vtI2AxEvgo+EoVJxPo
a6T8ZyE4s9CnUAuRQGwnVACwZVt6tRuO5AIV005ieUv3dipbaGx0lTNKWBBU
wEibdFSxXE8Z5gvdKU4o/az2rPoVsg9rDoTTefzQSYiQlEtzZ/ODbg0B7h0M
pAGPFGp4EojCQuK8yZrXnCu+YmK/uELY7Q5ao+AA2iwK/EbAZdp72jaUypWM
+lGq8tBwlEhGY8fUZa+2SJribQvFIbDfuF9WPeNhrtim1imI4jUYaTa6/ryK
Ps2i5F9kZuyu6xdcyuICs2Lq8yIkhqpaFa1axdUgh1YeyHYNDqzZ7kCRNJOn
kfs9OPAUyNNX/ndR1Je0zx998DjKXeSan5JWXpLPS2CQrO+tEsWXiuZh4O3S
dzHPq1DyJbLfZyPt4605VEWZTTkrHgg4nDuT7coohnZ6N+02ZDH1PwbDebp4
q/MshlaFBZ+IXta6kz6aAFZR8ocfVWTrZl0et3cZ0OIOhqRa74lrrzDT2dGE
7eaTP4v45QLIKjbadxbGeNrgWZ7TbPMklRHxY5t4vCGPa74042lO2ymtIIEZ
rvLKBMT9wtYwA/QsRiQ9JcM4ctTPCnlgnUVbrjgapDYpK6/r9WS6Y5scCHor
3kiKM9Utf0PLQhTuh8b/+P6LxoGCmu74IDScyzRVNsxflPhKYvPYs20X2MN4
uLJ4v4JpwV6B01vsHrx5qJA+apApp0s8i8NKguPD99oanLwedZTP3bwMsgQ3
50NSiRTkJi4GrS82s7QXbfg5oRSuYzWuaYHoOhvkBoVj5oOKPEFx1DjybYlG
nKwxX5vcSwpYNoaRMgFkaQuW88CTLPYXyIOG3F0UCrPGAt6MYxwH1n9ADGt0
qUTzFA2jIetny4w1FbL2SEd6NXDpQdYLCsgMspBvisWDSWHfQa2lYSVBkqXc
kA7tV9WsHgRsg5yZ1sKjrfPb8QNzRl5eukTHmRT7hFLEqmD87BzHtyRuaMFx
TOvZmnOVUb2xwA2U71aM+eyyLB2gmnRgBQt5UgyTxls33u7JKrhZ4pmyrIev
v1k/XvAnQXU2KWv3lTjWi0vfrml/GydiXXBIT4/Qk5cNQWymqCca5MY/YgGx
sRk870G1IYbQR1kj4XXaRjCXHAxgdogU7xh8ex3dC6alauBNx0lF5d8b79Rz
SAupcnEo4oEaLU4/eeOy/b5wbRgza1//7AVY3Q3uPRI9PYtDGyF3gy9vrvEx
77fJdZJyV+WG/DT1y8RSMj5RcU1dfKk1jJIw6Vtr95poi7QJlGaIdQdMNsG7
fPOMHAnOv82CmnVCTRM+05avrIwfqVFRAIHdvLRU1lPmjgfkWwZa0YdC/Dd8
t7ID0hiCzyv6+ocH0JrHBnDgr3mNmil48yE5Pm7OJCdoXcSVUnOx7zqJTN48
WFQa38SO6nFnqs4pTo82O8Go961u7UhPxVcwbgk3Ghc6p252ZS9YdGooZ5FA
gzksl0r10+G9SP0KTSn5Dov9W/QgOfCL7fVktvd9Mv2hB8G6v534WO98x2Qb
81jIOUyb8kMcwrb4JYK1HybNULW1LeajIV8rM2WCA7SD2lBJBf95uwhjthJt
Ke8hlUYgoI5XBbHx2tegNfHm2vv+vKA16M+FIjhPQcBklXi6Z/Eq00UEGX0H
hmuVZJvxcJ8FarXMzy5Tl/iyECiuGnUGKojcS7A1PkWb1/CRr9m7JTaRE7eN
mql7Q+HFHKtOUn01DvGOembjODOp8mlKBuM6gwvhgE4+DAd5TKexXGLhgE+d
QBfGVF4iUCGds4EXJgXccXiHqQzfEi6nJk2j9rjD6OSdx/D3rFLUnbHGas3o
vfD8QFsBzabkz/MfSn56VPmoybFIRuWZtRh75DcfUtF4iq+RAf74WRWuZOLH
YIT59ibBe4vs6EuCxiZmAo2AnnBesEEaMk96sKTesuxWh/ER+o7LZL109qQ/
SgMr/wX11S8ogGCdQf0ADw2OW1HQrpqH/t0CzGR+ldCIp6rB/5vdo2pKz4RC
/FEg9i7fuhTNfpIJtOsEeTjYhhxnD5dAPkzE4V7Qn1trk5n5WEjhzRvVCFuB
Hrhv0aVPOiS/BmYW7SpsM3p/7+JMfq+B/AaNQ0zDiKAYIT3pXd94ry4S4wHS
QO4cU5811i+P9hqINluUcnmpRZ/3GenUuIgdGn/r1wFfJlUuy8Oun8s+3GLX
FnOSAnrBuo6dTJQPA8JMK9ha4/j6hue6fagU1HAUwk7lRy3Yma3x17Mgucn+
dtK6TKaP63yrFQPX2AWk6+VU/8K/Bdqwb+CHjQhqVBbEigtw5pHD13GFWSAB
4CRzEV7KcZSYz2XzHyZUBOOr4EfCpoODTt1ijueELtT3mgVQlZ0hv913xIr+
T9BiDIVQwoB+f6YzWaz92eqBDsCSFhJwjjmm9mnZYHLQd3v1eu0ftOQOdIhE
aJZHTBwuhoUMdrUKrhf0OiA76evO1FsO9Ir1mLlpRdoNXOMLqwBU+8FITb4v
hlZcxwwPqUreaBGchDOjDg3PLbTPTPB9Y40t+u13AmnilSIQKJZZkSKVgWfK
OGAVN8gnH6njP6gnEampBeLEc77o4doPcJF1mo3fpLkmNW101INEAufkvTvi
2VYEhplEP70HKNJh1pCPV5Lkodb5S4JueYSiPRuYaSXDHCVbXkSogZU99oV5
nhqvs6ANGsxuZJ0stmZ9Q0nSQDGx/lkoMW/6L+LZydVUXph0SaQnUaBrXQG/
57/oClAMti9iDF/4I2Cr9+PlKqoLZ1A3p3PIi7Nez0U6p94U28W9TZuTcM8C
sSXx+BBsxJUOBcnKnweia1AvGSbVNUBlAe8b9Z7WlHXXPqy3O/I9ejUThKZg
yn6WvtypeuKDrZQAjq6fM3DDODiMsTTBlUKCcT5YUm7nzWQ1DbjVt2rhe/rk
HZffvbOyEWNYqe3IxyV4hU6nnCXaf+K8C0K3R0kA3iQCVp/QGpdScp4n9rYi
FHJ26bF/70hw7FBQoPMMLCXNaIfjfFRT3HIBaPZec/ZPzWxKF3FDqdHG97iz
klDz6bhIWa8StJgkFrRqcdDy1DjMZvKlVSNvHPbZ/M8QHnKy9AIhG/AA5vce
VXgtQ5c6iXakSJINgYkb8sNTG8gwsAv7BdEI39E+o1QZ+LOiED3zNaaAXIqq
4tgtdWYPglBLeA28i5YQFLOd8WRwVtJzWgsen16M3eEqnaSCPk0eLQTYWWXX
PMj7+v0cZXVF5A/8qkiseeO01uOEepCSN1DI5f2F+5MwnKK0cRoPV8I9asXl
sHahfB2JvnjpOcYuDc3q5q9/fQ7qFsITOpNZ5pk1wKINvkFL65a7uVIpVS+s
Ml3T9u0sDZZJp1RMnx1RXS2V33a//VM8eiNNx4dwDomN5V7bl2+S+raRl1fI
lxKDvifn1ZlZj48vikmTGmBtmqey3qGQYlYazi/Jv9HtSMafyvK/xdnGAYqQ
LO8Rmst6Opsf1XVAZgTsh0YrnEp6whoLE3HoTeXKckYjsiI0FhKG78jvyY8o
hUu4vkBQYne17zuTlo65fI7w5eiZ4It8XNaTbNuox60auLaFuE6lRBnKXqy9
IOiZpeCwK75xNTsjXzr/fMA6GihfaenOLtFTu5Ot7u4Kcq8DRFGaBMj0XXLO
YDA/hFxeWPaOQXo0hUWmrQFLeJM4DKGR5whEkhPVHRtsq5wifJEjiwmThXSQ
X65FZLGx2cLSwxsW8niB7n3/8uCaWMcxF/FdQFlB+uYFrCZ8iLDjiIm/jpB9
yY/3rqktu0iOtiFFWRbcwScwM/WDyV6ZFhLhdm+9OalDdsCAecvYA/2//gpw
lzYwo6StqY3tmI3OGV18eU9x4K6LQJYByzQwd0mHdUgdJN2oFXlf+j4cexyL
fsNsnZ//eu1mFPIVTIFmbexqGiHuRVBiiA4NlUoYFudve8zXPssO2Oiw4BBQ
q4fKwTPFy3Vn1DfT81FEY9Y/H2WkG9FbO9NgzrjueUaVRss34QGtO2brgwDI
LkWPT9waA+h8Km+IpZMqQAMm5VpbZq8vDqcsp4ADMIBAO4C0KV4mZ5qmC1+g
Qncop0VoB0A07ujn4XlDICU4LKLKZjhynti824lA4d5rCSAlwuz/VW2j9pfu
ub2/2BUqNO1pVoKor/rgKVS6Y0HQH31Pkn4wff2ZqB4ORdZyTWLX7FGcPsce
6GMGJwR6UKTXEVZF6utsBLxWZaz7FOyT5mu1WYGCDPSjO8uWgMJwSNyF5FOF
I4qmCDc40G6xwwb6VB9LOB0XXN2vwqrpVT9RXRIRjdmP8dRGb5EpH6ke/Qrc
i6S7pSNAKsQW/ucR2mE4xOsfsHRARoFRu/pkFmF1gMHDRfZ+DnL3FsZqTbs9
HpkNUs4uwEaHr1wlGdByNLNRhr1kRU86xJrHjhUyRoAbw7gZ0qHl9Pv9lU0u
bJwgjZvEn7WE6UkE5A8bKgMLUpiajXjZhKMzZ/5+SG1ct8AKTikT9K4XSFVT
NK9YxsyVJ7gWeWkGL1jaOfIe+JZlZovEir1feeeELRzpw39G8R/a23eGKZpX
+ue015Phad4na5jNqGyKPSyhtTTSMavAxQ3XAHkRO/7Pe7Q/cZ4c75QmPIvy
7lWY5ao42lV1GjguveNzaKTjiKBzE8YdtGUbY3RtToDQMT81UvMF1dlKbMjZ
CfDug0nNR923I0HNoo6jy6SphcLUnmCF2VtJ0I65s7UN1KCOWxG2ZTniXc0e
dMMqHcE2rA9RtD1yzLveau9yDd4ytqPn9imey/SBfrgPvcQkzyC0uvNbq3rl
CtPfQ3U8S3x/RLr9GLGlPIKRcYHmSAlHkqwKiR83v88nHVK4Ezs43jJ2WEXx
ArlL9zamxbTgnTuWF82OIqKOxHbHVFT570uC8WN0BIIvPGf8PP6moHL8bJsS
KQrwPbBlK8lnkRoGaB33b1gVPsPAINmW6hvf9oaVUxo72VBPdwT1O+Je03fr
mSa2ajIYeydNwdIApLXgoYGKo+Lw0tNP29EZ1KMPR7XQRUvkhKCk1KChWZKW
Dw6bczyHRTfpEn0MK6oRtV9RQH0eKuymcstiefIvHlGGXjJ6dmEzn+LOAWV1
cLKZZJoDu9KxBdbnjGPCe2ah2sEftNmIqyCt3Qhp/x1+s2QkhQD8TDkIYt/h
uJj7k5AxeNslfVZtU45ds2n3wfvsPpqNoEW3YWyx/z0jVjpZtxM2/+pXrrXw
J55jwNNaFPayLvHPhSwGoI5/41H4gpsDAukfHFJ8fZu8kR3NwC+XpvJstDbL
G6FXYMu94E1IyFVO/DAHtGeDdGPKL5w/+9YVIt6IbEeoV0YBzhjoYh0NSQGi
wWVD0Z3QEK7p+VkDlinV6AcsCgpyBG4LGms4wH/3fxttqy3tbZhtqMlevCOs
dK1vpxODXwETqf1nu03swP23r+wn8RuVJC7Xz+JhqV2mM6Uhd7cf6VBsbcEU
xT35eCUETTBqIhiz3ZDxTeVbAa7cBuwEftx0P232lH2rIKm0maz4+ctV75H5
r3oAPAoqAHx8jmuyN4mU4/ETv1b6Yx6paZHiwHA3+F8IoXqi/CvH0TROpXpJ
afTncmD+JXGZBA4oUo4j/JCToUYHXD6tjjvMEHsaTa+IGUfCaoMMZs6AdatB
jVppCqyw7nNyIZ8ETRYxKo6gUf6wr25KA57uK8oJG9EbatehdvljB6kfSEjI
j6q9eGk7rCjUnt8ERd95jcifOJmvfD/C7majKPgYKyIuKlKrhJZb7C0tx5xj
xJnsv9lEHxzyrR/yXLvI0C+j7bvxl9WmjFotJ3QFVmJAh0QPToPLCfkQI8L+
YM7P8oA+eVHaUMIBusDlwRemtSTC/p1gt0f7AK5pYhtX/0V1NePHTW1By3P4
sEi4jZv+2Gq6jxrAi2eyg9TWg9a33r/8Xe3QBRby2PlEMPFa/BT5+Qex91S4
2IhaHPZfyCg+lUcT4HvDBGiWgAUigRN2UmHqPVEkfNRrOdydDOLz4dvm2gaR
0oyiWgIwj0OFIwzv0iV9u1wkIBJkozdwAiHcKNE0fMml5pSmQBl49nLzR/lu
xLH1Jb3/4nkpaOg7aSmXYFAqpfTa781d1FSyd9kYixvME0ipLuB2TjxVuyHP
syod3Prz6OGlLjlIrZW5/iGZlod+a86m/zX5sTj9rdDfi3f4qQpm60JGNjOs
t0YUNkec38Y433jYcBB9WA5gSeuuuGjf7a62XcDkSRyt47wXL5Cknqpi6UUL
BuRe6RjTLbP1OwAvJo/Kr5MfbC1phFVHZ42rr9rqjIGBFuNB1rYS/mG3ngOt
I7noc6x0KkzWWGABms1PWnPacO0gvw2TDx+GiPZ/kODiKcBOmZH6I2Vn/sbr
PSA0IvrJHtmYZ7FT8dBYKdMm2c0d6WCPSIOkY6IIpn4HGAvQuMveWN7aIXSq
3sr3Aw7bjInRISt3myNyvclVBDb80ttbFw1q/Np2GBj4iVEt0PTuyVqyBP9E
wRi/qv0aop5GBVXkUeqHWOBrsRfziSyHWCL7rgTdMJc1vPm32ntM7iXAJoTP
SPn7abcPF8g3YJqIObEjCRPfbY1fSfutg7njb2oT7phGabbKSGdZ/0330Uhi
eq7g7zLSCZsOb35CZi1PssuzBe4iWRMnrj8Mn+JrMxnCon+HzhT27hJgtZae
7PTdY7Tfm80MyU+NCxvc4WRNdDgLWECtjsC9BHObV8+nnRQk6ZxpDy9CAhER
87pYGsViXHQ0kckAnMal56Vj2iE+hTo4V1UijDm9QBqaAesXMh7GfjVlTOiF
t0EmLD1Jtc34esxLsUG+eJLMvmLu5T9KZeujvzoOyE1a88jUXvYaOA7k0n7D
r1xqYzzpmDyoK+MiCW0AeAD1jiJFrv79Q8zs0fRoQAZM1l+3KTtVEigVke6l
O/NgAWoHCH8TEuAg8SP4d1k22m3d5rZI9q9ZqnYajKbaYKqN6DjGI6biJIjS
vXBH5Njcmf/nbDliT3QwPpfI4HFCRxnqFyDU33l+litGqWS39+fI81Xa+Zrn
WXu9wQGMxG4KmVe6cEkf1poibdR4mfLkvn8gLlpG8ZiiAdGwRdccjbsjNoz9
AsY/mIgzzbMpVAFPPf+DNuNZwVPqQPHRJFbfZmfchECEnO6u59uHyWlIHAGi
0DN7UdfNN8Rd1VYgZ177n13/x2XVKndg88O1BuNYx+Yols6WXZW67V+JCiFJ
NSKGnllhXNN0i8eFq/4pC4pgmCrO7rVqm3oOzowOWOrwVtUVM6wKMX235zNk
hcdvLhVfJ0U2BGmYyiI2VpsFG9hWI+FvCSnnkDhzZFHYSjxEOrKyJsb8evPl
aTpDjC4YNuIl9qKLIa/RLbVzWaKg5pd7P06m94ImGD8XqTF+k61nGesZKMwM
g3RhqvS4scYXUD7Ixgyw/WSuDsRtUwmmSLAHMwdl7k+q7wWlk7Y+gcSE1OpF
KzMb2HbRM+kMbtAhJiwZuTiCsU3pA29EN2VsEnAL5NHAV6S1a/tKEYl+VQ5E
/gtJjJDHQMXQBwIlCHS3KXh3CsEVWAHwmTI3GDLdMEMY34xUOlhiayYc8mxB
68kZBOhemVZBFJr/3S7ickMha1GMxrFaxhTITUUnDMKe4FoDVi3c40ThFrGf
zGCnksJ5voMdktlKftuTaoIvjAVF1c4rR29S6OfKtT+oWGwWQdUfx5VtSrq/
ehAh6Cs3wj+DTS/hq0Ow8TLSlZzJ/h5yGnDhcLqjsZfYbU+GAwTdRLx1kkZo
pYtQfhn9EbwMCdmHhavkthy+flwWustCAX2a8MIB9cvyttIOeVKg18IildFx
h0LEgx/KTLHG0Cvs/co37EKP6w9iknYQTl3egeKDZWWhd+/I5VfZ+WeZ0vS/
LWwkoNWWn1oRBo/6dMQkjyu6x5dULcSzQxszLWX9nliOQJROjeFkx1Tsg0yx
Bsqquhh3FaX2yP6Qc4tjB+WzAH86pSfxxr02grxtJnIZiA0tKMLOGR0Q0YNj
N9zMmjWBYs448Aaocsgo5toXgDp8S6Q493BMFI49QsnX8a08/xaZ33EN+lBa
wRDfh7GNBbed/4k4tv8akFBAYtBryoSP1n5Qdi3C2tflcs1fOjEpv/yxM9If
+Nu67XeTnGggT7/Da9nm3fBhhmxxe7C1UKOM2L9Jww8ZBmSTvXJJWSqoZ6p7
ippD9nYpaL6gYmgDrgQNoVIICMa+693tNg3Ij74tOIlJx/3J5VmKJJisBaET
loB1VhY7PRSyc/CwMWbygcWeJ80pkA2J2OF6lL1xgep+fuFAFnKJ6R+UP0ft
aX8TwyflTjivkF2n1UaJ4yY8WkYllCCxYeQ3so+Eh63mJd6/URl4IKeelA2t
kv69UhdCJd76+C+5ubPcHZN3wMn3JQWOgXdqIu1+5dZsTK1j3/9x++j7S8yU
nmabT14PY7TsRo9bdS8NeexZ2jZF0KPbr1vDODuon0tpen3hNRH+aW844Fcc
mv/YYbQ5yq4vyrwMCLpomE1w9SMKPBdm12w65k5UNtCQX+9+HWe/fVxAaPSv
PINwNm4O5Krj8vrRgIMTKrPPIEQA7X+GsjlWYqo47CNi083H+6D6ZYUf7Jxt
JyYSDZar4lrD9oVds1QayRGESdfTFKVYXgfHxw+ojcTunD7Wq/xGinwaeBS4
c/p9YkfY5m2gq5hAWwPF5UuFFKD+gLAWlk77aXipcPljddfYkrxo5pR6koA+
Z/EAIpHsbdNQK7r7RnoBWPIvdz8bLU5+WXolF3fAlvsR2hPE0P6LX/Q446jE
dpIIQvfNQLcbV0vlCE8baPd5PYRhPZMtqxHprTyy8UsGVvkNpSx/hNZCGdHw
IaLczBr2veZcagNkxYe4Ntyq/jG/KdVbrnhl41MFQykmvGYnRKh4Xbv+yw/P
mPqyyzAlly+edmz3iQFh7n0lhUm0Z8KJgCPxGWNlFspdmWR3a6Qkp4scO44l
WK7PFG7csk0W/3Xf7nceQSy2uWtMTxEAjGen/Esrgd1YtJ5WL6WstOaXWJYe
YbltTtdjfY4ais1KSq7YYErWQpd4TolyQDC+SrE6XxfpSUPOi+863CKr40qF
rMSzeWBBVLDMqk/d+OQE7u3VX8QKCnajkkFK+AYKqNYrU1GUr2J2nW/K0E5P
4YjYtTeVxdRvbgfMVvRI4NnLQioWY9Q9M/53C3mravqmlm/YbUCsGn2LoMy7
P+gbIyltkQJh0bzOykRXv604Ny1rqx6k/y4BPu8XLAuTuq9rrH5JeYhfOZUa
NNZPwnuoeFnex/dV3NZD4Oc2SZdh0cQD4vSaoSiHtgii0/Ul/pnaLDKWNowu
4OmQVMuRO4mJy0FV/Gfoaybqn4BJKuDuSAk5ziXAofDkacYQQ5lIld6ROWDF
plMspyPcNwop5wZD1n9klccemOGwsS9ZdOR6O/Jgdtzg4Afh35Co8LQ0zY2y
kKnH3GPHTRVUaNKZlVPi10UoGIhHBf8yalmVrBwwR14Vwp0qxdl7XfdllPSZ
M+iK07IC/CHfb/mvkC/Q6v/9of9cGr2Rgfq/FwgXpuGAfOWu8HDai40XbKAr
hfwPiAohxQMWlKU1Drwjcr4Yp4BR9ov06gZhzKz1cPBYdwoOPciVaiE5YT5H
EOXMpFlTJE/TXmRGUdOh6X4Yy1BXqGjcyONAvWnMbzSTg9tVA5q1k0c55Qqq
WWm9YDj2CRktbf1QEvcCQZD+4tB0ohi6KaAoukECySUedwk3gHuIEoG8L82v
k0pjLGv2Mqj5lJZ2SRiCKjfWW/kgTfQMzpvFo6A9YSXhSfpt7HQLVhkKonLu
HuiITNifkHAsLBre88yNHIbe/yXd3qgef5J0NtQlvSebZkpWD4tCZxpZ/sMw
FKlBAtURPqmRCfan7fNKSAXKXl++ORY5b87MEigjtThhXyE5TGtoAVtHJUVu
rZ/qt2aDk6veMkEXXPaKjLiYB6114B4AeR9Ms+Y0iVzWkZS4CY6PSKKdfcWi
+6oQ6Kq8qr7rSasUY8n9CDevpUjoKTj5KGxJZ0moKZZ/0yTZwVkVv4aHpynn
+a6vELERGC1Gj43ulxJ9WIxNoUZixw/BwedpcsF0CeaGYLA+1rb5evel4ACQ
LbUFkkk9vDc9/XKUhnCgaeli1sRcFT8DTurNiGYDaSOE0T3Lt0/hh1WPvDQO
WEq9wT/4F9voKtAyIE+z2NjhOOMcC5bYTwDfewXh2ctVqH/OHcn1S7x16sUN
IVPJRY6c1CNBF/sPmzidizHFhbToZD4CMERXdmuSWST+3F5G4Ocf0rHZxf+Q
j2wzyvYQdUBV9iliWRWVUy+U9XS2XUrzGT7j1U063GbkRpZwIS7QI0RBtC0a
9lzN1jmc97Pll/y0R1MyEXgakIVFayokS2MJ/jlmuqx72ViKgAPV1ID6Kgb1
sl137bVD2gLZz804VGgh45jdNfiMlJ5121gp8MysCPCc2GxDw0bPPGp7tkKd
PywKmQSvHogq9g6Ly+Vsv+xBfINxoCdRhNUDP8eVSTqxr70m0nQ6+QltcEjM
/gHR3od3g7Zn/+xCyh2wBsLYJBjb0Snkbk0sALJwbXqyMKE9gX3B6MoRH1xy
gkyuC7DVXgBItME4M+uQl1hVlxktKMBEl9wEg8GT6AtTny0kMqhCJzJJ1lui
sC8TEOf1wqMWx9M4KbA6zaag8DsbomceUi/3pxo9jpTaj2RO0dK81PFxadcU
a0mU0TC6stuixVPmNemnX6VIHBDw9MkDnqfUIjXlO8e/vvVsOa0fAYGBMKh8
+KMNwWAgaENweyAz1UNNk5Rcd77Br6WGS7uWH4OGl61sD2fingadG+XtWCgH
bf/ui9lj2Z3m0OZFgDA7M4ryfYVIOS4Fc2vZgCliIDlXufPxmIB/rIKdrKHr
cKRDDV9AikhPXEjUtzM2J1YVo4Fq35dzL67UMD5Oc6cC3BvQMuwDG8LYAlbo
gxquMKJYTsVdlJ9UZg/RFhmMLpapwiTpftjZtDfvD3wLNF/IZbgnH9yxc7LL
OD8+RVCvVna0Mw9co+Z/TySt2xfIozgm61p+JDrgGeqZoXqthKq6dkoc1BUT
/tCD7MelqCdSGGYw1cdm0QUP3e9sy3O3aKahAxEnN6cszdpz6ktx+TBqzfeP
nGT0xM8mxl653gJ/7UCBS9Rebrwatq02aSIDeeDaDpB2fHuDey8H/nmwtnP7
ApYgq7eZ4Q8+LqEA/ZdwNHkmJDo26efGRO9Nh/nhkqFqQ7YL0UTqci8CcV7u
2Qo3fGuUKANxhH3esm22a9+2ReSzbY+YlLirCyCt6pfFnPbt5USt1RMlT9zl
v7BMPmMYaDvTi/k154M+IQYEieBFgICh5eRdKUuJKwdBwS3arRF0BZWW5ajr
ejN5SBC6iFy2CQY0BQ6IYVKF4pHlYCnCrsG+Qw6s+qw1ZBfOvHFha1bacF0e
yxcJzCuTUcg+jq6k2MdzMdJvYfLpYJvSl7LPP/ZCj8kiOlrfzjvfHPb/SUTN
RZLeNjXV3N/i4tQpJdF4SW2N6mS24RxYIjJMfGy5lwxSIbD9/xfeuBUqg9sT
XHQFD/1yl28a89alqiGJ7tV44L+NkwkEaBhkzufrSsxHFYJMG0i2JaizaImD
e3Ijk5fElM6tUasiahC/jc0eeJ9rwj3UIJ2q1Lym+3lhkSiJDKdbTwv3jA76
9BXx5CeqyUZIOedGCB854JiwLibvmvlevDIxtOp+hXmAzZc14Dsc5zOTe/6j
I2Y4h9w6Ljbd/S3eUODjjaehVi/bWhSh0AyN3Sdi2ZdNcwmrhInjiLEgA3cL
Sgb3ZIG2BcspuGUDKqtUWFqHbfnAnsFYZgDaUcg6XZBaRAjLSf42lFQy5vl+
FcaTxpjeUKuSS7OFL0iWGDERhxTpILj7ajtjqzJtCzpyY6mYSadzlxc5JaHk
4VnN59X1eYZ/nQk3FJbstjKrKTQjGngWmq5KshDYWcUNDGbIPnKejUeYNgDa
FIAiEidfmezkJ58u0jiBa2c8SKmn/SEs6ibGigmKNbI5+43SUiVH7mAERECW
lxQ7hRJut6sM6wgySunsqhmf6AcnYgocKiK/UOj8lCvS9tqxPgitn5j5eeIW
L4AXSVW8p3X/P01DsaNrkMLVSKNGw3zjCn82iKNbxXRoTPAhPs886PehheBC
W3HHDgNNRbCufWjq+ON5dJCrZWRHJ0korG84cZ7k5glfxzTqhSNyq0hcALMr
eV4u+fHtQKsnuF1fGG/n955dgGQqoP39hzhtSdx3OulVnw45j0dXOCg7dKsa
OsnM35RkNYQ9/t1gSszjgBIWFtgnEFFMm19pTVYUiXjiibu0eQ6eNujhOpRQ
KABWHka1hH2nys13J8RHwL4/NX26XE4eOaBrT/r8De55LIKiVE9LptVAUkeJ
TWxg1ULWp/M/+jK9E/JPq9IavgnZo3PSwVRAiZ7DRtp/TgGye1yIR9NYI8Nv
wvxuSzdAw6wmV7LSu5S8fHKqjFUbZLqhU/LstncjMPhpyDQRdP5ofxK0zv6k
111xYekoejYTCDY3NI07wXs+ecat/E/Gcn0SM4t84XNkiu1eP8CUlAHAgJHW
gRttpzWCYH81zOzTyl0X5nUAt5EDjmMWhbo5pPFDeza9ptVwTsfKQQn6sjrV
WXkKy/9+KryLI713vtIc5y9cU6935Kq1bBnyoCcLgiO2kji1G6AujmFQenXw
NzWe+2RLHtiEQ31ydKnFJRxLeTK3WGpwXD4vFswT/aGzOuoQnW5uMwotqFPE
WNVvVotqil6CHxiPWrdyxG6bH6/C58yl3jV1CbN3WHBCuslKGqGpmAsYlWF8
s/q60khPtfmOYI6TyZyJylOOJ4jsN/U/+rb+kFk8HYjDtToIguXRXWCA8kT8
SJggAb9VlpF7mjJcWuHc3wGYy1bCLBMxp/rUCugRroEQLiUnNAZZgSLwbjnp
7W254gyM0e+BrTteUPB04tgVoa0bwkXn9YRCXX08HF7YMbFhRkXwdovOiabv
s7fpjTliGfCaVNqlBSvLjzJ5LwFTwuBdNDA0oPn3NAkWf6l0yHrh9IFHUXK3
xCZNOm2rl2vCd6svwePpwdc/spXzP8MvJpEHpACi4RGKL8j9tHFwcFXGUNe/
SAPbhRHc7OrA+g6zWJZVfInxde2c9CphLS+lPfWmpe0zQVT9kT/1t9dPXbeq
NQyXz+DGNbMUxbwdZLgLD2OKjvSLN0jRTXyn4LX8X82AgsPifEtEHvJZhQ+6
0943L6bnbouNJ1oBvcDMQNuuc2MsaoXn0UZHj9kv5eybUC/mh/8hJo87KwUS
7Yk/IoVlLvWpCCrdIsMHnnaHDahmuBO4R86TPrWRejOUuvce9vqHDBgsN/pO
+h8iVW7UXEdQKkn22YiheV+YQ/ve46n0IJaTVFL4B4ujyZz2kI9j2Pvfbhy/
yrcmrpvHL5Qf0sz0EQ4LQgUNZunVE0tzjzOwfdPzGAH+Ra2eaPKddppywL76
Lpnu8gIBM6b0yjW4M0J5pvWU5Y2+OOiBQZ1LkDYQKdPM6LA3lhJd5Zkc90Fp
OElysIkAL9inNM94/gJAnXh6ZNeSzxXpShm4mS+IBL/eNB1MBYKU080EUYWf
pEIoG2GcQa/sJ0MAn//WKOGk2nejKv8evp/OpT1fR2j1JkxsEPUvch2z8z/x
VWr/3eOYrQUkIzhsMHKZHDprUSP1RyVsdxs8aTDFFsC3XM/H0Kn2b6OkTi0v
Qsk1SXue3tvEBlCBe4lt4NMfDYKdzqD1WkrQTOBPSajkrmHHi4aUfeUfZN0x
/XTCaBY+fgzPOR7ctM0o6kOhXFNjRKmR/MEgaIgx3zVgJ1Qy/ER/FzfZtWE6
oLKCnYxd44wW/e80RN/sH7U7/bpA1FkOQ7xKL0/q1FjAXJoTvWfcbrhTQWXt
dv5R+bsfng7p4sNMk11DhvraEv0ed454Z1v8tHAtxuELLsoicaTDOqnkIZeY
iydIqpotbguxQxg+0cz+UBhUKaNQZTt6AMOXz2ixb+UoLUv8BaIaNyP2uH1M
kQZOSxRSvS/7UTdsDdm1LkcV48CUEjf2PNlvg8mqEZ/o8wcBX/eT1vD4mRZd
3f4GLhtvungJOHv0RJBBINaqU46N5CVC1Vw0T9uyuqKozOIJR4+8/sXSiLND
ihwqopvpNFMO+xGsL6UEDZIOWYpNs68JSR8hvrwxdYMaEVk8tcCF77jgF25P
mcdPdksHn2+SWumIOIqcT6Onz6JsbDU7JymSc9FvxMvwi2sIz3csBXnGE/YN
54W7IqsNKBbQiX9SLMA8nDptageiflzi5jdp7hMnXN7T30WgCshPeeJdUmaV
cL6KQ26X1R8t6Sc6PPzl4TkbgYdO3Jscjgt/Xd26NDfirmBfjdfa1scY5Jim
kuP5fcMB44p3PnHv6Nh21tbELwxzeI/MNk0E4SmoNmyktO4a3iGyj/Sh/saI
2cpPbdrUDyBzdmf30RVJ79lSkdIHi0UU/blDQAWqUhypWXi+465x/i+5dHnR
R6vXuJff3PlC8UwcMfT48ejlzDPb+29eL/fvd5bMr4R7ZPsA11/aV7rmoKYs
2lFWArwqPDuw7kY/uoj73IiYrkxlED25RYSzZaXRe/F3N6aVovh/oUcI8/cM
yDxL09E2/Pz9aeAZca3yrS+FrdZwoxsd/PfqvzdBD1yTi0nagQ0cvxsaoUvV
O4ziSA7dyo1+yM5ZOhoBnVU5HcoBFGm0F5eKGtI9Y9kCl5TTlqUZYAdqMxi6
fdKr4oWIjwUHfyf3Qmx3pVDlIhvJ9zjoV4VWNku5c125tVa0NuDc+gCchIt0
ehU6diKEKx7OxSlXnmZ+HNSb2nlahiY2WUAARy94Y7I5EdCRWQjVFQUf81JA
tnE4AW5pwCuRkBQ0PIa7hvZOup1vqH9NbUF5skj+QFc3E2wzKaCzLnqEQA2l
zYJ2VH26n1QzY1lUTzX77db3QKL8nofz5QYyPYMA/OoT82ioZa4g7y7RTPsB
uKNRj7SBECUe4hk9ASifkhxlriBdWNd0PYGqAEPkAlUCcTnZNxdJDpS6gFHm
6g2XA0gruwYEpCfpXlZrwieVGL/neKXlUG6KkcOLtos2Zi7+sY5BdvrSJ+rA
CRfghoVBjMFWHZfmp5aua8Xvvh2n9qXJMBIzfUsrUvR2JhCEfjq7SvPKd6XQ
FKeCzkfIR506tXn6Cg9ZYLEgVsqSnYOUnqAUsIIxX0TEz0P8iTfc6x2AYm20
Nm5FUiFC3ZdCU3Knlc/Gi00GcsbJEUKm9XgKFEK34P0bbOL1s8CpzMyM/tl3
Cr4EWKO0C5AWjd0XuOFmaZp2CCHmZjJKpMgD3UKbsO06tS/u0ztY6CUlCTH1
UO0kkZvPPy85HOMVlCItSds5/kzFnDnkZ7eaUZ0aW4Bv2xUUui8G+NvUfelV
9iWzM9FqfzmjSuL5jilumiJFyKl6jz5qRnhx4PTtP5HvglIqErjw+rLzexCk
fn+N1gcJwcSgQwraZlnBmEYDPDh0kMwE+REFNgK+Vs3Cnjhgzhy+4SRd5Xg5
LkGW8JC4vZ9la6Bb5Xf96SMtsY/PWxI7OhG2PClsf/G7qBLxCgJ1pKAoI9pc
be3AsDvCbJvObCYkogSL5NFZSkP/QixvEZpMjopk0RUS2mQl9KjqyzJCGaJz
g4yV3T/0SUrWYbMg9TfPnquTzSROa/aP9dWEJKjja1Ht9uflv9h+7UnRARui
4XBcDl9MgNGL8z7ksFPROSS05+OSO6IfUfRU0aR+THxyASNT1ksOh9wqWizY
vqLMykXgh5kfQQ4ArGisu6fHzsdEwKVIeihtTryuikV6JY89sacFfcXGQBTA
VCQnpHzeS2/aSsCRY06qdjRX6I0UbRGbAYYlkE10bVpvVPbbbiKikqq4sBJ6
pOKH28b5BPXlAJemaRtApi6OCM7VKu5c4MNDQl8UDRnyTOKyBuuIfl69WGWS
sWVITF+YyEKwhTinzcFpmax2wiOnKZEf+OY2xkElwqJ7YuK0K8KjSY6DvRh7
Wqea9MlVoRV++wMxjCvMNzTtaFbNgACdjH6SkoipMj4HCiOuenF8gGFn/SLA
zJKJYGFe/bPZbHwJYrHtJosVqcRHS5fsm2Vk+XcfUiNZRB5+NRwJUV2J+WQg
TXICTtBg9aDi9MwoT2hEIo+fj6/eSdABwimive1d5IMzswPeOI2/Gso3J7RD
5j1lL99hKM5f+n0aRXaYBqvtQVuyN4aMwLpw6qI2iz9yIOW5XOrk0QnZasrt
4w7CyNzBM5+m6kIZ30jt5wMYiMEPB/rsLblyM9g+ln6Lja2XcotYr7mGq3yh
EwaY0lfutoGi7OW1MP8ncbYCzsjHJyHY4GgglM8R691yF+Drdk0HoJ83Dg8k
1CCO9mgEP83L0FHycHreCZe5qoo+OTs+5Z3uzSkIJXGmxkgQiXCkWovCga8V
x9Av12MHSO7lCl7aKywAEe+ZfI/P2zMC1NuqBaCq3zVTqMNXtJMK6ud7WbLb
n3KkNDNE8cFYucGOatBJmYuDGNZ87nmbmQz0Hnxm5Wc4XUqg/Qo6sX4cWlwd
lGlz6ZYj65mZN/Cfg4hiPqQwP8vpUk127Ucht+Yy0Ij9LzGKQAcwLAgGlU1h
eDZ/dhiOlFQc8oenOaOE2k0G1PARYSVmfAULMXo6l0kvnCuStrOUD6p64atb
lYalFjTFnKy1OuY6eDftL50fxOaamz1uW3PvvVcX8Dm+R1My+gqxBWaztwDw
e77u9bL997+eciIpFnI/9M0HHo5glNPVqdpOpIx1LnwfMSIAEKHmbyTBKHJq
H5e4pWvXzD6V26BBYxHbBs5rpUbjiybIeVmtejIa8ioMbz/8Bb2zMDMUmiHV
rpcIpmelQcJ2f7yb9Lbd5UNCWivBmY5bab+P0l7azjN96CWIDPMC+VAU+YEq
KMmoGuz8DHIS8wio1s0Izr9HmWeysCXBYtHDqOxdxHE6aYvj7w2GcvKeslr2
WiXNvu31FAw2O04XJ7dEJsknFsbrek9DfwxiPY67sPRNGJZtzl1hD5Qc5aWl
sIWmOe8dLXY6laj9nHpnmSEQ/huuZml2gYjhzEYI+/3Ltbr405Cl83yyRxVS
0EWaXAJ700rybnG/kIXeIUs/St612H0+JnH2XKbe/lFs3hPqN0R1C4u0tPP/
b8nFxJbMySlTJeSP+hJYTGOmbFYTWxmgM8eAdrXBS+8ROdTI20ldeP8KEav1
d40YssAXVO2tpwX9i+GD+QwuP4Bc4etms+VlLspqwRuZ0FfLqN6j3a0+2/Vf
vMGXz5owqzOChnefCe7+rok328/SC7gaRl16Dxng55F10PtSnZbxaKXx5Vad
X8aNqqTQ1pN0U9IKqimqmIp1J5ZJNd9kJvEQU9WkOKXKgIBfOFBCfpTwxlqo
gPJdEaLMy06dHITzoWkVlsYlcOjb0mGm4fH8ypX8w56FST/VoEcNYFEtCX9x
b0JxpmUBos40CtZSvOYhzz4vCv+JhqYV9HrKs9CRDD1V8bqr7MyBogw5nE+O
V+424Cja+yAU7Yl1RXfEzKbkc2Z8bkY4zbKpp2TN88WxuDcnjdWB/EWsasGO
Ln2ai9TuVl5tEavtG4262TjceYQlwe18jx8bO/E97kFwVLvZPDC6JwsmREhq
X3CtsiIoJixKaVi78eImi/rqREgIHgTxWUwouKhYlj439QgZ1hilve1et+dg
Rf49pKgl1RNZbSWmcvETtt9b7WleQcY4Stk6XK4z4JwDp07WhLdL2YttXNws
O0Jg0kZpE86OZ6gd9X5yhTcATaatIuynbCfA05RGs8Jyi8iH0mSMOExGzQAY
SER9RpM/MiaCxKRSVWC8voN8ITj0K9bfyLoCqswVRnRZ+UpQ4YUTFNIIj8Oz
5gcQpCoW0x9bV6WWQn6r4jECdg+eKe/8veBftzrRmYVO6uStOOUvsTiQ5c6i
NXDu3wL/J/LzU1EbteSsphfL4af63azAjKf0njfRrE7TC6vxXUiGLZKa9n1d
ZaO5kIbtKsnBdqwPzje+fibz1IcmV7ZY/isLhSUHGbJddesnkOJrhpydLM7q
9xmluU4efFzkxHrrMJ8qsjpUX3TYey7kSk97Oln+D4UObtvsUXtGHa5E1/To
lOnP1IsfYstglTlH1KbvXceVxd3G86bgpI7DtOof96i1I+SE8HLN+p67n0AS
erjLwq5KkTXI5gPBEy7CDteAyDCxbFSBnXCRbLpEpxqKLG31KhuMpLl1EcZs
gRhkGM4P5z6pWmzOHqq/22BQ5lsCnKlF6fUIDd2hQzfQQMF2HPAwZ86qJc6c
ddh14MN0z6P+6AfG7oBLbVP5yxkjAkc7EVVeLl0f+mnrOthWDO9dv9SRGE6R
CTTl6SfFHKeULZA+wzkrGFTzXF+PsRCYEi0p5EvnGGPVcwcmyjKVfd7aIruC
VBzSNhp7O9OZW+3m1F2tzQoKNozUwUeIlBa9EQvFG6zrejswzKCdwIvunrX0
8msS/Q8idoulDV62ieqcZNlIeHMf1h9oLxfd+2zo7UjKD0hDmaZX/ve+7cBD
XcXRjAfFY8OuWTj6eVXA/tJiwvQLz6LWMHOYMVuYUZcXlWKEVYXDeeEqznwQ
8sv76J2q5SXc5wMVbL6o3Mo8u8F4g6IqT4assFFGHZpDWie76zWhTNIDxG1G
ytaN1+ypZsRp88zoPeGBIqyqsswxjzV16qxi7qzOQoWmObdAYovckzHiIVj4
y80gcGuEk2U7VVm+EK9JaSolF50IrZX9LhswWOJ/qUrkR8r44V/tp8/zPSHb
SE6sNQMFknXeMvmdLBjwu/m40ouAoFpmXmxb6AJPWQ62AcZzlNbvOo6cBMNu
iILAOc9iQnqrjdNKsFk8t2QPm5C2FtcnSgFw1Qrqv1o6ccdTd+hufSkOK6c3
vV3nbCoD8kansYL80yAN+IGsiwNGo1I+5rIAN0ENS4seanlG9+SAncB9w4Kr
OtyvfKKIdN+shuNzww+HFCDPBrgTBdmXnlMVFiKSXO982SZUD9XFPD8Wv2ip
7niRur6D4bTqZC6ynwQtqGfaDEiTPmUGdWuNWo0Htvwy+My4iwYcVRp0b8MT
jmN5ThA6SsJiHI25BHP5OkK/qTuyByj19LdhgjW5G3q22MWWDEpIK4ywNd6n
twDsNyLDCAj70mxZ6QiRfKa6vvntz1LIpdWmPV7k9J8RyQjyecHewr83pQVC
XVyG2jSQ+autjRHOqkOse+EV0m60IJmMCZqjBQpby8epYeDlZejiIwwZ5h85
yKf3pMTe2NW0QetvkMoHx4lSppDfehIN9mLNPaCavogLTRZE13N7g6oyu4yP
rrL55J1e3KCZFlzea/M6zsPiQJ1fSBtEOGItyRWDGDx6w+EZE3bxFlxwNhzc
FvyvM1HRKoZyJDdDg3DZD2aswZ2zBvXv5JcGyxnKvq+LT04TJT5JfsESBz6e
Wgyr9ZrtDocjI6JHtL2V2MORZ2reMVYflDDGnti8yj41aktBvDcKx3uEr4OG
34IACR2zJTnaClMs+d0vXUJpuW4wCQk2U2h7LTsCNT7p5sjhAJSOHzN5mH6L
pTc0ZLD66NyBJKHfONDASLbwz7dimAOb7yGYtpReSVBJe2c0y/Y9FH07lkiW
33A8UP0879DqUCED0NeyjMs1gOZ9jTpmlbXGUog3vma29pvkaIWfIPcYtwxH
VHSEO8i4TjqDeB8H9Tt6lmDvad2Rw16ucr7WMAZRfEWEHqOlTTWP0dkqDcaX
XPoys/npL9r2pTfd14zkgsZ0OeoeNbStAiCDU/zmiaevmWhUE938uIGadlPe
dNGWutJhWebUqBu3niY60d+ie4Lv/LBvBdSDGeQKDYPDv4C77priPyMl3inU
FwAoTivEKSZ0DaaSKFVcivp/wjiSyh2fc+m9NhhcNCUGcKKd3bVTDKRRQKRp
ytvK/34622xj933kn7xsUMWTG4UZz02lbaALSnbgC+oRp6oBR98oHkclWI/K
dUQ+BGRXNdPG7MOxb9rNhbpvy2bgV60Qti4lUrF63hJsQS+e1uuyly/RbYvk
3FeZByd2TVBs1JOs8bwScYp3cnn97vyxH1B5RqEtZSPl2BsW+MvNykzJDU4Y
Kww5uJ1LxujhOUk4bArtv5uAh7sOJX+D/HZE9+3djqDJvE+I5UBiCL6POVnc
4d0Q78KKuZBbkEabQw9By57+sAYeiMZ79qU5dQnGWfaTaoOD4KUZPGxAcS8F
/DVluJAjlVckwWip/SmXQ5ixqJug9mO6iLRMcV4EHKxCER7iL7JOu3+megyv
WRcl+zqeUFbLbjakqjV5+CKlQXFXlUbpHNA8GqDp9dTdZc+S6dP0iIToHFyH
K8PbXVBKMmrHp4IZYW7xpkmxbaPwwWlBunII5zWUBL3blzWUcodGhkuW8Qcp
2ikOD2OLXvfj7XKljujB7nWy0Xp+sih/cYYlolz+zSJ9VsVtxXTnjtungvLX
kQQehtxSDaaVv3fGaInqiQ0IvkLrAP+wxsQ3aI4+rrvP27pD8vaxbf1u4+DY
GLeg7oYLP9jF5H64jUC0UsGdsfExTNd44q5wYmDcgN50JdeLJm/KIL9lGMWb
32HBh3qBIs2aFH0+9wdRkbXhx6ZsJaGq0GTppGmKi6dM3000WoOCxTmV3SKB
ErjVFV4WrlFXltf3uvqKeiiLNr+PYE2QQV6xUvrROtKG2yZM+hq4iFUfeYXW
Itl3s45CoDCgVN88LPXWR1xa6Ct8WkTS2zWg1NrotpPwEa8f0u3ivYb83Hwl
mZh4j1nNdoZbJkN4J6bQWVUoi7ZMLjv7BDMtrWfpUREfBMeO2qU2X8tgtV8l
q9UXDVqIkSKwG6n50FDB9Yg6BhlHwy9exIL7k9NjKjAYn/IYrP9Cphe6vSm+
bdsGTZLPqppzURSJZ9VxmtGG8cllZ1L6yijRqyJY+de5bSAbRvtSaZK5qd3P
qit52+efkFDjPMlWqlH4+1+s9gQrPKlZtsVR2cVrZIfR2ui8jrqNjcAfgliY
YCjrvPd4li1Tk+rSm0OR1p20M3ZVz+VkQBZ7GWvwp2Kd0IiG9MZ7fwnewRAR
2uqDhHO92SnnhtuujvLyc1sheHI8jmwLobvpbfPXW289UO4Rk6ak4e9ZL8Hn
ymd6vkj/UG6+x5WJk0J9aYmTQNlfkTWgk88EJhvTPdhpaGwmGakI8fskam3c
s6FUfdTKqANLWWHh4zMcVXxdnK/54jgAnhP0CPOgaZHMd2I186fikvkeU8m6
NSqDHyZbAQQIQpQj60VAiCHX63fTvBUmBGm8Ub+wtjjkYKTpHAleWA5IrKzC
R2AYNGPn3DsNtoW3eWBHA6d/hInBK8Zo7fcXtzKJqi31u0LCpPkfVnCkp0I2
Ih7n5LojyF32YLkKXnd6BEo72d/16kgE/4rHhhV5n2LAq11U4rU6Ton60lnx
SQ3s89FQTwwzA4WUYH3vkn+RGB3wWKNsq9spe5NptTM6/Kj06xhHwggmrbZC
H99xBMNygXEoPkEbW0Jt8zw8VKOWlfkVEnVYqTXIjZkP6YjupfrSa3cF0ttV
bhHdkNtPGW7/BmyA9tm9CdxW0Js4Rg5rG8UcaI2p1gbGHexo3MaOjduHsbmv
UtuYoIGoCEe+njOYtSQ5+uTYsx0/qHYxJbdCFxSXMEWum6BMCofPXn4sVaOl
7N0M/4aMNMTFlGoWYRyvrO3wnbEy7pz/xZxRGnQyurW3k7A5TcTJgUxQrcMB
e+q699P4HFXVRExqwnpILwr7Np6/cdMUcQrGzFGgXfeuXa7gyALoflcLz1sN
Ibnr2RwCdfDiA7rp1EcyYnbTQsANcExIBEFig5GkfQpmEpZuqfkMJ/lyIAPD
YmY8Kv6iDo2Zs4Rp3iHyeXyHO4LyW4lUF8M70PlLtO1j1AZimIdhClcdS3tF
VBArd2EyIMbrpjpvlK9qyRhdFD0UvpCh5zI3AisDoDz8/bnsbh7qaSDs9TFF
a3TKu3yLdWvv6OKCukqIlUxQlsSUSo5apnFlFzeevTAI6ZPL2GhulelCBEcJ
+apH++X4rcDMyD0HAOujuN47O4akcf7IL53zsID/7hqk4cRPcI8YvPG0c0fD
CszjmczKXSIZxDabt7JYY89sjtnw28Cb3YMR4PAOHPzEyvok6Ly8RFvW9XeR
fV7Di8XOWpAMAmbBestf9hqcgMwXXjYkQdFqN4lE9r0BGQRrxxmxXlwN07kF
FwpuDYn9ZARE4iPr8Qfl/CMSxrxrAfLgvafUwMS9BQsZEP14rjF0teZv9xZO
dD5pz0XP+GY3qLWnN5PKNM6L+OBqA8Ivcfmub7lM2ygepqHoYRte6gT9IuHn
47SZPKczK4klzHYwUV/bw3zQ4D7KyVqH7Vfj4V0Nod4DC4iO5IGeSFBoPxfd
RXKaOit2iHB5wCICvyDY7OQNGOzy8jIsUWzCFgiq1FzI25KjGqjXjz7w61H7
XzT/SfHaNtfiaRsu1x5Qo8VWb37LLya4eEeebloA4IUiQILPvZb5DOFIUZpw
eMGG5EWMpPvKrwJcMahzVM/1h0lyPQtCSw2ByUF55mDbun+SqpeCYT4HKmHA
9aWEiLuz2birfg1TCVtfkXTIEr7+w2ntxwWGnphaSiZ7h4Iucq0RvXC5KUd4
OVcFG0dfWGJa5WujtDlagepwrkNOSKj36bRLPIYTx0amw8JicmbtnyTZuuRA
kUJvbn26VnDjDX8SmBS0oqnXC9U7GZbPpkgdJjP3QJhhzmss5FeR7+aneQX5
mAOKVmMjVwYrshe0DP2bvfh3Rt4X1qt7wOb715RT4NQvZVY0dVp4PwDl666h
ckNR9uuB7Q8MNm9m2GYxu9dHuNEZGYdP7vUvD6LoFtLBSEHZIjWCCJdZPWzy
OeIToS+FX3AywomSKnQWxt/MNl4G8CpdVvBVArSOQo58k/QEh1LsUt2Hoiha
bHSXOS8xW5PG3B+oj1quBDdd48yGZ/42SP+Jv7awIku7r0iNj1LmFV4avIx/
yQMtVCSSTigvwF/2R7ZAi6DrlD+upRGJ0Ha/Z0cppoao56VE7M/JTc/vBFNF
RAwzAYRxKJt3nR4ohcrrfKCfIRBKyCzyC3muYZFOwDLOBHSCA7aH6A9V77L0
RaE09+rELVy+XwKZBVrgx6QnKxZC8vYQtnhAXfmDaDz3zi6CKY93FU0PIrWb
TG7jFgBjKqbetdxlkhkEkVCGXhecLMD2OG9l5ZHGRMtcz3G5ixIRr0s3x5rG
gxS0sV0WpKGzReArTi8tZYRAobkrN7bk5ujFPm01BcxSUIrq6vfabylzhWLC
m52RnRfhaQFSwjEliDyhbTIrLs1VTl6JvIytckXa/hpEkulQ7mgeoqCAiRZ6
UYu/wilUl9mKUtKd/axcr/fGGs9KE50gq3vfEM+WBSqFcahMHgf13J8Ktary
E8hA4eSWUmRRTpS8zvzMAoSN18lukKTFP6l3TfqI/KNjHFMjMcK0vMGOVJSh
a8tcC0KtM3zQ5iqXbqq9VubJe2JwU5a9drFwhduBxGH0/XIQmRo0L66eggBZ
0VVpvNxDJqYJnFftnnILFY8qqZMWTJ4RUPNDfaBAFgYTrJ9fV+FeTwLqKTub
zFDD/gj/WuDPnv+JnKp3Ob0lrDtmqrnlSNhx6HYBjjXqellNbqiWHxHca8Ql
gRBDOJBtEqZSIxZJXMszOt7jx8cNFj0jYhmgyrHog3ZKiMiVYRaZ0u57zSU4
CDti3LpyowKdnQLXeF3+7f+57/Bkq2wSNPyKjyGVQ3uvPVdNOlzqXLaTUA/h
ppumj+PrVIeouDUPWNWodTZIx+GDwEyKu1CgTUY26oCc3AwcFFkPP83dMLCD
UMA3/NmfIDTjgKmHfcsE6v9pLLgGM9Yu9ssCysDP5lWqUPyQfZjRW81pEzK0
3JyoqAg6LcqGT2+zmPz48CmzCr40B+LQNlR/wghbl/KNOQNpnwrh9O8bbUXa
fqAoGR6H+wVHPVtCs3Yp9SHEK3f2g+EuH/NmxIjrfjYItv9CeX9isxpXprfx
devroI9IqIQbQ1bSM1zUJZtV1IIs8E8UHOE3SEO36cAwbk9w2L4FT3rst5xt
aFUAUoR+6tcV6BV2rS4cHAflQxDQjQYYmBLDZmTv5iM9WbQdxnf8vPJwVY+S
dz5ZqGjQuNWOfPJQ+ISCqLwGcpkFW/4x0E8ngUsa+YoAcO8khE7vRgWvC7hP
Ndc3/p3YWFdLm3xJitcS79zub5vCs+7EF3OUocsxC1GZ8lbXRzRqqgZXKbjy
ZYRRY4hUNhthwMFYkmL9DYONmEwftpPVgq67s7WQ/JcsAxwhmh8thvYAuGoX
34fcgNre7lZmt9pbUrD8ybRJCTXRUaKf0JT6eq0oFdLf36Vh75S3y7mhJn0x
PAj+RziFbAxoo9nTkhrU0VW9o61wO5YKPAb3ecH0tjo3EuCJHZmU1HBnFq8b
14CYOTxuHDxfgSx9m2XhZCHN1EFPVMmFO6jVfRr+kInMeh3oHrBfzwYx2+dn
a50aSdOwwdyDTSxI6KckObY4sFJa4kPe+IaIUP1gzz8XS6oyzpI4V/vKZyH9
FUMbuZzAwk/FC6mqghei/OjZDdLOX8acLSAcLdzrJvqCNxYZcKXp1BicFwuB
2PF2pW0OWNUTKQ6M/5BED9/jI/BN0KfG4OPy61fAfXUwmsAeRPpOj1J7u4Pm
znbQnTsA14+N1e3yub2PksB2UTc+ezP9MSTE+xObahLM2UkXISI3pR1Lr88r
ErPVwKK3s2JNj3IZRi9tCHIMrSrK7dr30Dth6Nb0xAu6v47hm814YifxDaxA
e2l4F6Ff0pnPjX+NOPwyB8rT9jkZTjyDaNWH0PxJVcK7bUnW/NXAIps13jAP
inhyME9Dc9xebrqT4CdOavA8q+D4SrCDOeHiyvQqv4d1OEbVX52oUoE5kTJc
QlQ5JuAMUIBfZAUhekgAXn2OZMvWFDUZ4rUEj9f/yPMxyZIFCVvdrHQdRoMV
3nJmEt5AQhUezp6dvN9/j6FrFqvGhDw7PX2pK1pnTJPXLHzwe6FAPQzJ2cSQ
aj1J52AH2U2STdITZYQP/6V0HVFpvlhBqATGvMhH7HDy6UeFJ3FhAoWaj7IK
fidWaWKn1QCOZqCl2UUbp66ayCHvNwXxTMwSJbcQr2fkR2tEoA952JPosky6
0fqVYPbLaHSiyVIOgjthyT1fuW9BMqP7AIpTKKWpa2ld8dSGSwXrchqC6WbQ
ZK/z1ZaZ4LczBWtSSvu/54Rk8RKEdtMqEkGTGyngGgmgT8YykzCx0UjdfzQq
o8u0hgKx7UOtgZIH200JaDk7avrFESSq11Y5FUYuKQoTgkCTJFJRnR/2nMZu
jRCmibO9zIuEWSjS59T9P4gQ24v1IylecO7eX9JuoKNs3YQm+2RtT/eodJQR
aVcZFl1g2IorbLfYb7Bi/roCL8LiWa7ZZ6jY6PXxcjLGyaSBGm1Gl0+ZC8bK
hUXPTkTO4wKzeYQBIMTSOvcUTv/yTkNEM0xBPs26gHZGtxsDZouI9MTh/evJ
12sIzXUhuEsw6TNJjB31O+7gca+2IOakQ4A9rSxjkmoCA9QXiuZbchrACug4
LAgjg9cKXMpKHqO6Morsge+ys0iZR+j1p5wHCGr+PzKC38rJZmsByUdtmAQ9
5RPBOvGoQA5KAJrfl0+S3F2h5kl2FdROk7e2HF1XXRXMs6pgEco4DQwJmQI0
Gae5IF11fTfyID2P+SqkOJ4CNaPwJHPsfJ/FfJASgBVggToIf6Por7+CkggD
+furU1vVDI0JA9SUGOra/sAY101tw+zrbwIELxdph/j1khwuGD70xE5TB911
Br3zH+f/ebqztNuzBYnPY9P7oV8zvi9T5aA84FIXTSf2C8i1GjdcjEJSCZlP
A6UvxJm6D3ekcVzW0CoIGiGw15tvqg0NoPHvLWhjmjAiJPLQGrkGKGdFt1bQ
CVN3x+AF5l3/ctnlAWCzUKnKjB2Y6JV4gBSlPt5m5se20SKPjDmp36B6nYg1
XGtD5kK0ePr/oXv77pS6dSDP3e2C+YbDtco/r5bd7GjgWKPCVTqdgQqQoySI
P3wyMeEGDq9CmKIwgFIXteMp9A0vWOUy81I9y4nNHXv4LVH+6BGZWeDfMoIk
RDmnyYkQDkpMhw/HikMP0wstls1fY9HSwShjPzXiLLAYmrcD92yPileEFv8p
OD8n+v3VU1Ap1wyQ0OmEaq84GjQSO2T8Xk8vfycVBnLJd+8mAIJmpw5YLcPz
S0j2VRd7BHTIYcGAr4Jca8t/JxHtijo+tVFJCLTMsLelzVOkorykIZcgnLPc
3ks7K97UkFTm/XfKVj6GxdZZKGAMaWkTbbweeWf3BWrqf4Dj4cEUrhIB3dGk
RR9GyeMg/mcpNtmDjMSgXlkqWAYpVbyFI4pMMP2r+G9z9DMi5Ta6XP0qlkco
cQSHiKPjM/guKvZbKsysE2emqf25mmnnm/62dWM87aZVfHW+SBpKdUfy8pIc
mrswkohy3LsyZADiiUotqlBxyxBV3/FXlTsL5O5D71VXfLREkrcDVFk4O9UW
c4RBmD9MVeG2++j6760XBsUL/oKyfr38/98sSaqFwLbUKW9V3JLsJbl7sofU
m48fxQPbRaCuCrmWYH5D+tuuejn9BHFhYWof5gLKCm4q40EWuZIRFHDR7z6Q
rsMjuoJ45mYk8m5LXKLd+wEdoJt8+uwpovNaZ+i3pW4y9WTYM5ppdpgH//Wv
JN5da0pEL+hFuEPQ70uDnQsiqFpTyLasJfPQcwfff2miD+i0/IohSPcQvv6H
MiyyitZm10iTBj6RpypKzB19xbcZOeIsOdBD8jIxalTFdMml1TDBk0RiLTNr
Tl0dO9roOav4HJXdc7ZNi+zDtOlNYcc1yCsWC70T8KsM1ZNMvg+oAw6S/ii+
9YdVUJ0DfemEE8v4dEg6oV3pF0Cia932mjGKoqolLyDTiYV0Ng0RPttNpzP7
DAbUR2qU4IZP0nstEUbLSWpgWbfKmLwLnasAICSIa+qPiJ29H/j+rrbFQrhK
xLOIozEm9OdMXmu6GrJ3EDCzyORRdRTtjd7hOqgFSkiS/OqIAmd7wLfP3S/h
8EnoBxSVd4wIBlfidCtlvva7MEzkJxkDvEok2PaOLuJqFL5Gt4A1mdUuAtmw
NzSCSYuXpTJDyZaqSntLd890eQAghEs+TKbMnBNF0H2u8rzfJM7VsNBtKm2Q
wwFx9eaBdgHSbGbaUOHxLTRj24uyEyGlq3sHI3164vXfwB+T4lUuepp5ajWQ
JdqEb1n1p/uR2Tj+eYiiiY9aJhpyjBkcNVzuTH4dB4QoyFY4CsPG9Nefcxpk
qx/lOdTHgFDH9fYPchYT9GtWRQVon2soP1mVcud5CBzl/Z5s7hZM9UUloSy5
C8S5+GgZS8UYt5yEa+iaYisZ3wIBVN/IZ513kS3xUJL6t9G1XfiDPrho1ZqN
q3ZBTHO55Y2ZLfOSXIsxcmWCC2V8yhitNdn+BFDGORIPbdVPbHb97SNJmrCp
xaC+Sx4h4S0Yj1L6DJayPAkxIc1lkPeyg01gfLQDdrcQcKz5jBEZiWYuUhIV
87qlxVf6ltleK5wf2BgGv83upQ8YFSBNPz49/L+wDEb+RYi7E1KKBHin2r/k
piGEE2/Z1dSZWria+TY3AvESWWq1KGyO2KDG7jeHy58BxJ6y7xOs07c14s1S
Xk7j1+/tWbA3NdkJoC8KNG2xIGqKhBA3Oqepk6kcYHnWWunknI4yuZPOSqXS
7TkL103/XitgDr+4seYE2R3yYzrvJYeKP8E+Ex+op4TpceH0C94MfrIW/qhE
Oh7NXTONJsqZhNj7sG5exUAJ4FtT77iP7x6A/TulTQ81UX8NNw2PhXCvi+w3
UH5HV1Z39q/qP3GoU2cdRgWrvYtpiaAQr3jBwVanD6e9OvdMjcxHPTV8hxD8
91dSpEbbqY7dS6FWf94e/A2UzlKY/JkAJdRqaGhTEDrQIfNf/uoh/JFCXFV2
3gHIsjqrfyxoCXHYdsjRdFdtU/WUyqNMJA3T93C7FGyIOENUtWZ89YgrjIqd
XEvsGHgXyoBIuvzLnZ1nigUjhYquqZi63zxH73rAQzCDl/AApqPEB2hU+B3/
lkbbRaPZFB030uirFaMqXWboxv4k6/fP6YjBWyYn8XT9DwAc4vS4x6qS1bBP
fqav1Goenk/vBFsjuY+gaIhzy3rdyczGw00rVp2E5fWAEocgpDMU3tNIWANQ
uHGjExKWIYRJcPa+jj8+1szliRB3zusMJ3zK4uG/OmioMCcFra31zzXehhRx
Lc6uvWLJXsjxaJXK9uRzBhipgIm2M2gl0G8E+Zey9YfvS5J+kA/frS9xTDDa
3Q2t1xr9ngA5zGNFMPK4yX0219uT5dQgifHkEatiDkYiy7r3XFkrtWxvANL5
G5Tow+VfXs+AHxIVXfk4ClOgOpWBatjn67O9hbh2cFcZ8ukI0uvQh+aGGoUw
nYlwqXfdWQBmDL2sATxSiO0Q13uttUKjGeKPQZXOfptda4S0XGA8LlyGV4g0
gC2ZOBlsbI1Q0c0KUHatKMPixr3O9ApWlEl/C8S9CbrFcvQ5ZJH73gVYWrYi
MVnO5Z47vE5oqbUxSGh2+RuiCfY6xpFvV3GAlbFwnaIN1LN2wrLdv23aP4+n
KaLz9fNN2CeCLOvHFxtoNDoQszqmRQ4VFuoHN4Gpt0iUxLCAKDgAA8jGREJT
qtwB5In3z0InG/YkrI1hOPFZ3jtR7skXwky2PYSjynbyY+J2Rs9tye1XMvUR
W7uVuPeGM+MGvsABNTUGG2vezzF2o8XN95xm7mqx2O0XZw5PW+Q1JAdD1QRS
xHAWrwJhvwrUOr57vzmDqv79x3tjRaNLftJWGQb8B+5/08ax4uc7RLpC9hwP
EADrJi+KAoHpoIPvo6pFSR5JJ9H6PbvBNQI5Yo5cg+6omLHWJRrurrlXTsOG
gsUfXYZKkanPJVFVTyB9KtEMTbXEX0o7MdnAxgHh2AyqcJ4T5clgTC7Qq5Cw
j1MC6xSFYsJ3Hyh3iNut3j/qVpCRSeu0azXk4kZPbdxIXoc+szoC13xRcLM0
/IjvHNk6QUIgnkPDxFhYTd2vqWkFCNGqRq7bkOWtEtyx824JFR0TUTnuZ/gD
bbkcja32s2lrwe5E92ydCFSCUtoh4Nb4MR1wXF+0MjrKG97GbNtg1B2d2ptY
UPjNvyz3kIOBDQhl/icbWF2KWoOomZI9imXmMiTMuw+dohudRWoDoBTyshso
Dutx8/l4YatJMYDWEBBUDSEbYV//hKZduKIzooGEyeGQEtEF5l6NzFkHed8E
wCtS4Oi3Y458FYbjkMsRXplP1r91WIyvGZDiy7/Bhe2WPy5UKP8xpYwAWjts
5yGrcId2O1Wsp4L26GYV+dRtG3QhfC52nJxBlY+GPnsN6EwSs3kMB/yDrmvU
35/L3UfwcdsTGrwhEBGp+RqP97wDDhfdSng8k3HwHR5Tr5sy8pZ3gRCTghGk
d57lSI/7mpgyGXGUC3qp0KksfWyGBar6+y/1byBQ9UbEBb6KB82LD8k9Csv5
rZ+96OH86D42BsMfGDevBJ0b9Rc7mHa3EhwrLVjSFz2pay5jDtNQORY7BjWq
XGYDvZldr69ltEBhEg28ncbObC7ZazxjkreauVxTatlQS9q9Q105g26FiCW7
99yO0YF7FpAyzI497UAFKTJO5V1lG4SbezxBuvCvulSTjGAGjTJ5+iqHfqVk
uwDy24GubaistYirByu8TnggLhGHKN/yL19wLus/0j9idixlSFIh1Eqwgio4
nMmiSWkYIxDIPUM+hDwAMgK895BBnzzH9BNrL0z3E3hZF4Rq8rLAtx5bTEd8
MAvHnDEkPG9C0rajOFqm1psup1tERix1hkDyDFSdV3rDrPK534uzivXaw5Y5
Qbc/E9Xt1MO+X5kcPYExN91howW0l2UAMMKTt1sbAJCaLYeCbuMJTgA5i/Ri
pmizKKKJWepeJtWFEQZOSQRbYaCyupcBN4UucYTEqXhH0gbuVd8e0VweMUFE
BTxhIepFI0DlluPmi+B5dZkEicMeGBWZGrN259f0pMWOiUieKnwZJaEm0m3e
Br+nfgE+qjCaRefLIfuF8xZZz7kUQTfwM+sxiVFVRvnOXFuJ+1H2uFVNMCMT
cAix8Mp0JrGnWzr498gAGy8XGoMmau8dkPG/5Y/QKy4x9aqWd7meplEW8dwu
Tz/JbWnf/a1bWH2n9o3HIgvm6ALS4dJV/XixnoQm0+QqIMN6HuEz9uyQzI4d
TT1GRVEdrwaPKIzYjYJOf+eo/Q27OEx8U5M49N39Za9RRnPcopZjxBBusniZ
OL0i03uMjdtPdxUwNcBh1utcl3GcSYOHOgow/tOUWfjnrDi5XtQOhDjhGh4P
h0hq4/oc4aN20VWB5DbH+NvdoaSX1eAMv431zxrgldkBWRkzAwyck9SOpc12
QiYPdKTlaDFRzAZQ7POFMKXuqo1PibTHaGVbrcfKQ+lhObIucfV9dKFWrFjj
bRxDZdGNLfTUCoTYipA1SPZmmtMJdyg3FDOP7keljs/vgvW7Desn38u3RUL4
/BkFEmVO9p4HEdjFJFH7dwysb0nV92iphubUR2gW7TPKgrOCLElsL5gz/C3u
BCaWspTxKgTRtJkiE6JRNXvToMnLgE9IPsCKP+1gA5sCLuUVUz5ElEseE8KO
iPElLUf34otDg/el4j2Xw1VtHcSA5vWeWj3PH7JTuEWfh0S0IC51eTdAP9JB
kVKcR2pLB5/LBvXfiGy71xDxIrZmt/J9Lpjut74eviSnfLNSzUbIGjObByEd
9hpvaWMNYm4x0WoFISgZQhc4gkklJuTDuOwYyuB4DsFDUSnAIhN0/d8dZf3S
LiEpS4slbUVKZiEESmqGi3uovQck/jmM4DN7Lox3NwnTrxxWBBth7V12KQjf
oZjPXdWaaTn0Yyl52xOhjpbixkWIZJCoENaNObNCKqJcLez3A1eXLK+xdZpF
hNMxMY/6zo634JLfoU73tQO6H3Iw2fy9kKAo5g5RH3BHO8WRnRj2Md0g4u1C
+RhFavYp/cUfkg4uYD3S10wAkT0gGnEYZk07lKFAmBq6bS0wimv5zvhkRZ5T
HoYHUdWlLsRYZGKsJu2VbPeZpFQko/pZQ8GVm3SM2NThhH6ClWNfStKKnAjl
lWXfeSbrWfmzjM1PLstq5mdPPmzA/ZITgXb8eCEdfZ8CPX6uqpknSJnMZZfY
fslZ2pyuUan9A639bjp5Snj80UX/QTwhaY+TL3rd0GGLuYb1LFwN/6iK1d8k
Yu6/g0md9u5KP7ffNMFUtuKxO5O4JrN04T/NxCMpOeZUoujx71ECzDqAANFJ
r+HAqkx5rWTvqiA1vy3/2ePZYubZxypv31b6D2TKPiCegvZ7Id4uO2Nmi/Cd
q+TAnD5UO0U+UPUxBorjI+Mv02/OqS+skix2A486uL7Ui0qP2/mjigMwyyeA
x3EPFh6tpD8yQ5RHRhOlrcfJVDLAs5V48sYuf9f0WyXdU5GVAOKBQwOBCom7
NixyfOvGEEDtYXkXnv/MQ+dHLsxQk6W/qVQv0JlXRERO7QL2VxOL65JeJrmV
PJxZ++X5iXRkxNp7JLTELucEQypWB209x4IzL9429F/WGgO5bUF1NuzUWRjK
3A97mWs4/hr2dCvOJTvNX262C6yVkRvoYu4yphSksTqOx5wOJQYFH2HlBwIW
4M9r7nK3MCpJpo6nnoGPVXDvazmZYkHO99aOJLZmxF4gseIr5up9hKhYKlkm
eRCk0LiMhAEH6LlvklujMWoO/+0pmkyZo9YcXd1XTEGOalwetX+ieu2WW7wb
iTv/DMLAcXjkK+/4KgpuotsqTBuHCKDaU/p5LSQiWzRoy/1bgEjp2D+D5Fj0
mNhIigyTXPSQgzmV3Bp3XXXtCDsc1dx+0lETosM8/Wcfqxeu2JyI7nTAab35
8zReYtHjVXqNhSOQ6mIpCte9/oTaZtq6+FEDQFqMjTPYxK7WibL5Ey0++EmC
vKzrXAh6T2SrQGKeqSJZW4a70OYl5R9bt9Y9aRs6iXJfVfkaFJ+GfRM2LxgO
Ul9INipFhbBYxxl9dAoq10eL77zCMh5+6OliD+uZICqZXQMvZ3qtiOz84ysh
nN8c9t8Ia8CCCKmulul5oXCQdcU4ihys+uNtVYEmAwt7zA0pWlVhrDF1EQ1z
NFTVok+Wjr/cKPQXbVhHZlPQiAbSBedmWJ4XYA77rhilLAk5lLryf97ttjiJ
KI/XT9j0KWMuhDxe/gWdQxT74MfQpvfIxK85BNQ8+RTjLnRdKMljHCFU19zb
9oLCwr4zfenKyPYxLCxpB4tcVyUlhBnhSFxqYhvd+BNpndvE6VArHj6/0bsp
r0r7lvUxrMIxLAmxsfYVg5TC0ZFS0xU4G6yuVkKXptZTPY5oYOYRO16EnKQy
zGEi4i/p8kyV5+M7ewzYIGdF4KdPRZ4Lc9Ilu2OkAYQu4slpUMLM+IVIcXhv
VSfirB/z9pEH12TktF2zAFPpISr+d2Pa6w0RiviOvSN6ByDEhCWx97AGrLLK
6VUV9fwLwqbVubzMxro9jMJry913Fh63mqm3jAAX48D/SGt8G9YVPn1ezMJe
RB55Pl8WnbDaoA806Je7XyXCjnOzoIToPiuhtR4HmikAsUeaKFfkAGfvL/o9
ImFNvE6NBYNcoJC/OYr/cBZbtG+q6Xj9iUB/Bi7CHb0z0SxO9+XfV4YFwHee
9AwoscYGgG+n2oKsID6gBCFz/c1l5i9bwEIF/W+BPRjiEb2D895wh/9oXj1t
CqLQeBdhEqUa68Yq4AEeh/2nRvpgdW1t58jDqFlJEzb2sY90Bb/Cf5iex6y9
CLMZjc0oFkbBECXAEA3khNjHcgAxnHDVom8JtqFAtgVpAoIDNEAJthWcERfd
3zfO9RsiS55G3lhcXsyfJbUbX22YVFx7u6i+WVccSPk9bgeP/db2vz0LQXfi
dnI57dcD5PzuQEFiazniUyVInpWnHHtBhe4dujArjf2pyGRS/H2Lc6VTHMRM
S6OEIMHn0jPe1pURlp6Xmmv0PTzf3GCW4FmENi9VugT9PWF9bRmGM6/mOvTu
K4zWsa7T097KOdwKhE+NUv25Ur1R+65an6thhgB/3CLmbC+eljEeWcvtg3EW
PfYxNnprGWNzRn326wEKZyS0QnIbnKJ9Z0UA4T+vdtPsexZERvhD7Ml8xmIL
FXAzW8lql3vhi47Gsimh/X68+zorXomqpA51Aw98FBh4J2iHes4gsDH8ZSJk
Ftn3XMcHQrRYgSyIeTkT0ROtnZVI60wQuCURgIavZwFbBr+9eHP9SNjKOX6c
KbEaWxV9iE7W7WeMfC32Udf12Pm3S5qCR6WSzLN53WyBWlZPfR0YIBkTfXpw
vuN7EG/0sJWtBzgwSV1W/vfDxiHiAR8ydc5WoSpA0Wo1A3HiwJwyf4QrY2jB
P4/sBb2lgmUqMKZZFl+dTYMXjivjLsePKEw6jrGIY1zdT3l0z8bXFojvfMpV
JCaFLmS3WhtS59GJYoiBGBYDzkDudAopg7kCj8dz6IJwhkLBeOy/UxVDb9ep
au68A2GGobEjXgTTjd7QiGKkIcseJwvQOAqAdTOLVskchDUcH1h9GHv6fodz
qf4Yfg/5d59ex8C6sLeATS++6S+X6DvgB+211twaT7la1g8CNELeYtv4zYTQ
Z8YeRss93cKhgXAX33aAQgaeecd9Z0NUyfvCEnaDTF8xqMtStNFBsu0EoEPQ
B8ez0XL5oYnwp4+9rkd8mhADLSdOGD6XgVAYX1Rq5jUlPA6ZPXx6nAwK8MC0
96SQ8uTuWda3ub8fbT3NHfU/vT3bBrZYYYM9hi6lPzCk11elsZcvHFGnXuOC
a0ADkuqViTAgPX1Wqtqlau3hGEs7cbjyCzIlGKU0cKmu+4wMCBvE9dSvJ0rk
a0A/6lKH+vZrWhc48zjN3tXEb+En1NSeiPX5OkqEN1PydmC/Zg7OizvMthgp
gfa9/UVZAxIZtA2hvOtmUKwvqh+0DnwafmHgxnvGgJzD5RPklZziVT/cYTWQ
kUBkYL805dVdlA6NAeTf1HeHYf4TzHAFD1jsqnp6pAlTcy4AYEFQJ3ehtBnU
O4ZvG44dXOwBpcVrQVcqGHPSDL74ZyFSUugq2sU4EKUNx46q6yjwc4zyUn9n
ZMvyRf2Pyn/k0LFfhfItUC/zKbMUt+1PzuDe1PDUJ2ozqELkwXguzdUbij92
QlH1l/T2q/nGKICrr+iHJ9wFtOkGCrxgn60V5cPNIzO/cekUng8U5StR2r8s
nazDUXF6N4vWpayVowFmmrJtYAIjdWaYPG4MwiPRAEYWR4GTKcnbMueNFuS7
kVdZyEHR4PgHPBL3c4yyX++ghpDEeT8hQ6rKHMfyKxUR/8QUPllfEDDb7XgP
zgKQjTtr2Vn9MeitV62TdjifYO9j38pSnZ+Mdrt+yrwllUMXZQe7l/jWYCw3
4hqmK1DAvoFwVNHpcs76PDYY6X01NYCPGi1PnccFrOr5B0cXkxMeVb193H/P
lvJNn+zDe4o0A5hwJvovjZiKJv5mExXqYZKlqbm5cIsOIHKgylIAELkx60CV
Iv9wffqKxGsNcEKhWiQR7t0p2Nx3VYlkynDNLy3wsQYb4Dq3Orm19XOj+Nun
kX04FjippDFMvtVReogXJBt6YRFipyzo8FKr7/jyKXrL1eDYclzn8k925H4N
y8r0desMuj38ig==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "221cqLfSQtZLwpVKjUxAj0azxWo9qWyTHel1yyBq9riDaTa7pjyEaEdGOLLz3wcrK5rHulca0g1g9Zlx/VJp3su79bVOdFJFOSZrof0/9wf6C4nAWrw+2PgJSzMMKpaFLO6gpDFruW5083aTh1M+Q5KnW16yLzHWGhpxtWHi5x5kzslfPRMwe4HyZUYh8/FwJanr1Um2jvkSaUjUKvojtHUTdbUpkWg93bqHvMIamskBoXE1RlpmKi8f6aB+KKYZdQe62GuBvsq0hKAGvoshzq0uY+oYQi+HFtXa+Iw+HrTGnVkTJZzU8VjmBPZM1JgsJLzj9o7GiAlzXrUkgASFWlfLR5ulJmDqumvyGu5QSmaBdbyitBSoaTFTYp5OIrRcCDNxoTkGHkF3KZ+gHbkWBylMiYk8+nUkCUpsF8aZBipEcrG5v1EZmcdweg4px0ypf50S3cENF4Gc3GXS+8ukJybTyDhe7Z6Z+uI2FmwcucnGui9pvUSvfENocoxztVt64anypiqDJL0CT6GWDPhXxrGtOZYIXMTAs5/Vk6IKwvjKirr6qNdUz/Xv5rSdu1NQn5/9qvjF3+Bl9SytXcpuaGfdHCUcD7pvYn+7zhenbIhjUGhzeF7Bb1LwtfHKRLEGmdEsUAmfzq8SZoFm6qYtBh4alNbmkDZCT4RdCo+XMbWDDkqOncHJdkHJijS9X5IzJbhdrhCPuyP7UiIa4fJX+I9IN+Jje4mKw3lvFCA2BktI8lacqjX921fLEuX7ZEfPDijxxParSjrvdm1/VI45htM9Qnxd0aEQV+xXaoOVoaFOcnOuwa7njSYzJ73yymaJUlfpbWplklBlfBtN3+4OJAQjRYZc7HsE+glE2u8WE9HFeA1bs5bTfx75Q+qV+i8szUIbFnLWCJi30gOZyW0Vt5ZUHFhbzT8BCCawzY6y6iCBXeI6naLmZHTWeBQ8b47xX352oqiAtUj29DdfjxVsZqYcxk9TQV9Y7e7rr8fy79Ol7klHSso0KY6VwxueHXsH"
`endif