// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qDk9fCNVPRJK7SyAsmMRZ1PaofKq5845kZ3uAsAFvYZoYJ5DsfwB2+i/HPgx
uYsjl1KKdigwnqAy7C5e3C6DP7p3c763+O7PJcMjS+H1h4lTRhlT1qIaZwB2
JvSK+lfLQ5YNtXVK6/kb8YYXR0Yh7oqOrkmtVpFONwVJ4wte9emoddjRS07t
u23UJ9cImrNBnNWAxDdmaWb8/l8fJf4l2LdJ7Tj6/WyPkTpwvvktUEAu5uxK
FXTXIPnVTEhlEJbCsudnZYbqRq6O6u+k5F0ZEYuVC+zhDbtCQ8++B6JbLt4z
lOLe9yYEaqEtaBIHtuZsp1JmmqazApnMzGI9gz1Tcw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JZbKkjgjj3JNvJvrfijY35t64ut7QR3X3l6pGI3hUVy53rD53gvAZKSveOvv
Bsw54bEAyv6rTe+FLuKXNAI7T66Kv4LlAPy8gIW0QZLWFdScYzDCnz0Asknm
DakeopGNUD/vRuM+ko5LWoD7mXO7IDZ79/FaZx8xHoa6DCgZL8+leVarh9lK
EGIu/H6rEYIog4z8YEgn0j79rwjYTu9IncS1Hvgx+aoiquhJWQtUNH0bIMHE
j/1+KWoc0pMOsmNdtEVnL8FRi19qoT+krhXeE6zehOgLnLxDzahoX0cMFSeo
c/ECZOKw53E1hhtDCttgc6uI7PvPh8SGdW2OP8GRqw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Puu71iwg9E4jDH+hnStOfMPIRaC3HDwJeaLB6jy+aEB0nr1KG7NPUhOlWbrv
riGN6ywkfJBuVvX7F0zS1oWlIpRoG6dIf3jCC7HnxUhHS5nFgzYooJImLJU+
y/RiEYpg1EuKTAWZdiS98MtPu2HB+Q2eJglNfES3qNhHHoHO2jUvYFWOOeQG
NrVgrqGxJyDHi6buE9kif94tVU4hUpHduWhoBIZb8eNGGiaDsTFVQaH7CxGs
/kCAwbAQKzxM2AZUSqIpf5rAiRb9JQjLpLtNChBToiWeOh7tBViAYVs8mQIf
OgzdJ0rlpP87SNPDtozn1MCTrGHB1d3VFaDumgVpBA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pPb11kNiy4tWbV9vcn6hj+qWF3khlBwMty/S4qp8r2mZw4k0318TKuI0z2XF
QksXmQ77q3Ra+WuPtRVeTQ7q5q3eC3ONf2gpvnevwbhA4lm0CxLXP9FTcP5r
Yq/2eAzNAjuCpIl71kLbCBrhhA8n/K4vf8XKWUyrNwUOhwV/5C9WkHoDwd8L
dCec/KeYSRKoxaRBlkX7CWT+PSTeqxVDf+Bujy3Y4+JVUQj++OT58QWYS1sD
001N7HN2oOLG/l9aJY/IcHAj909y4GEV0/hWmX0HpaNdAeiHWQ35S5q7BVb0
U35hQhzd8qRH0iOncZMXBqog9zcJqxPOpIyn1YAlrQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
q8bb1hXbZthf3xvXZdYqeEushCwc4H8Cft4vsaY+EUK3C5Iy7lpgYZgzsVK0
nNK23oDPZUiKO8u0P6CaCbKZlYjLCZ8nW+ZMxxvcXMXm6WQoAzKc7ehQFkwS
Nhpc5b0N13saM2C2Bsvc7H+TkHBsgSf2qlCGpK4NMA4WHL0Sw/E=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
xcjhtJl1jKBufXdX4trCl2dDTYR42tm1g3rN9b0Rs+OCqTfuRy0bzfGZO5Lk
UUtaLQOrfa0vgju43rSX1+TJIQ4m4EgjeSyrO9BiaVLH5DEycL2V+8ZxGDAa
kKI72Z5RNtWjLAnfgq7dgL5VIvn7EBahrIrqou9EHslIS7JpzIDV48LEnxXt
GB4+p8CIVsMnVzhoFqujEllDzSbjPx32Q48yapkyoZmmY7/kF2L7aPBbzB2k
qwvPt+kth4jqiNgL2xZHFgrPmBqCqlrjpbg1jMh4U315GoQLUToeQ/WiGxJH
sjcevEq16MiSIXeeCfpEy90g1QVb7ifpXB1qw9y/Kw2/QqV1b2Se5d/fw6hB
3NdWIzXzRBE0jbr9KgbzCtzZewOePRPZXxmGZ4eF19usy9xoxE8i8M4ksxqM
YVSCMsPgUNxW/9AW/6msQU2OsAGVeP/jh40c4GM3uXuJ9Ty8K3gxNOZNhNJz
NQvMIKsHsMHq5ZAv6bVw5Lg3dmCFXqsM


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SPUVi6SHi0AaSsdB80SzwmXFduRvP8TKsZV55nWa7bLU6DhtTkYzZwV9H2MT
DnuCANjWl3IypnXbOUGbp7sxlhZOFXZAcX4J7M2OvTMfUBQPgoxzT1zrkev5
gLroAm7BfyQC5KFKoeEdIpVg8pHH+X4Dg1DYULuw++OYSGkJ3Uk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jVQYdC7P/7nwDUO0lAXIjvVgiM2UgdiIgCi+mRcEWStw4BezmyE32Fa41AjM
qfxL4OVnCTdkpMpFdZthHh72d7JDlpnsPsK4zhoHUVa6npRiXCh2sW6/Hbjy
eslqVirds8CKFEINCT2YQaeh8MOkmP//6exKhg9mOoxLot1ePZU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7184)
`pragma protect data_block
JkfztkRWwR5jB+YezGSQflgaBIgjVlmRqqLKdCKdjwmN/5TE97EuvdZPl++v
hHIn3zKzynTKRUkPrevpn3n0jh52Dza3JuVzlvZK4ACkGrZc10m9aVtjXZcA
vVE4A62cQnGjW2dlvt5OGEked6ofopRosSv2DY8zJBCaleQ7OYNvvRS5e/zy
qQsxbgzcPr7jeHeqMXupQSznvzE0KoCX2kpaCs+j0G/jkDX9TlD4XEAnlGaD
QIMoVqTlt911YQZkvnn1fZ+xC/ZnsP7kt1o2+RRPdf6V9VWf0k69yk6w1NaD
guyFjwpzXBsQdGeMaroZY3cjZPXmAsULHK7+gza83qGxJcyfXV7NpcKD7ylA
QzpgH5fiSXomNfRcnCU8R0bu99dWmh078w4IAzRY8uVTB/g3G+uJLW77RNmb
1Sl/QzAV5l9LULTlm7td1oRtc0pvUl0uJ7B8y5P46Jxw5aEQ8TBIXGi5aLZ8
XMUPYd3UTWQ6CKPi7nkBQqCktlplTKOtkrq9EMGNTBIlRL63b2qZX88TRT/s
73b5YrXdJTlXQn8oxyKvKhg6AdGKDftDk2eST4hzksoUm1Em+THjubD6Ipue
g/tiDhNtrkGzBe2bDW+l+vGsNGC8NrwhdEetk/Kok/ljUGRcwxgHiCZP1gfn
vXKnoFBKOWNlTwsFK35wVcARYzOjPtg4qkfSQLDbJmc0LcVy9ITZiuL3K47D
VFe8ueYoEHV5Z571/myVMWOTBjAGUmCXvMDp5FFSPooXyMIj8KhPo5X54f0R
nDNxnbynsmILjYpvx62TLPsX3v2DOA8zBBU88TQ2oXJUhCIAqHlKLFlwhEiA
HxhSIWqxpnLVpFTCVaM4WcGWUC3A/lwIPuGEK3PWOVjMR09w5pXOm86Bdi6K
QXiPlYKHSTynRhc74gWoEfs/2MzSD12qgPLvIX0aD6HUXDT1WVrCZZ02XXTQ
jrLRGt+Rvo+CTooTXNEV+hVKMWhOCMQHMjfZvGrcuwAalrVeLve7InpFlLp7
KQrWFfBB/hBQBryLsyHt3SsbdOhqsZiiWkHoSK1z5bDa1pjmTRpS3K4gZPCP
kof00QcH1gyw1jv5eJyHsHYPygXJo6hSoLo5cAzFMWXCRLrr/me03MoFAqPJ
c8nFQSSrF82LU2FMwHEp0V+A73kcXcTPWSFQK+K0sSd5YOM/wIvM/9ESKaIq
Z1ynkle0Kx5B7WT1ROei0SLK00cFIHYcgKrKLkHRm0+j5rMtY+nCP5aao0oB
Jaf5URHSo+p0r6CRHvnC68a/poBOAaWS29bjkceM3AQqMHiRGZTMJGOYSSYJ
0q5hrIQHYOPWUJiTrrK4RKnt/aLB1tgF0xpi7PYbolc3PieRbZ3Z6InLUJnM
tgcAoFZs+KnfEVpX1RaX3AzLYSLbIlg4emY3FpnhSDKW4Oz/5lVWCSaRO09m
Hrz6jNnwb/rQrB4K16aqE4Bb1BqgzQT2YDTvxOa4cNmFk0UvAWvnaMwaIYtl
gEfvNu82wv+y3FyMZVu79xCmNCcw1zQ1wGUnWnqJMSatWGdFWDZRUcK+9oGd
Cgy6Og3AP9RqSN8Tyusm0A8BKJqw5uo+UJsTcPUm/9w03yd6Cvaz+rDUlZbd
5XqoLSqUkpU5YMNfuA5tWFxxsOErvhSmEpWGiJwif+cNkM1MIzYNpemETOlP
xoql9XXSZlRYzBcaLBeEUO4sVSMWKSjJ7O3M8c5KhbAMjQmmODUwrctEKwtu
Dzd7zQEmebG4LUkbQ0wTOQzIwpg9Htfy1/rKidWXwPmssh3Zt8E56BcPLc2C
lwh3aepWI2GQj38nWO1tmfq0E9UEdNkbur6zmg1hdaOo6wjqNY6hzUFLH5gD
/t1W2F60b+I1mcmAokJ+dNf+kmQjXHAmJ4Zs5XBaCT8p6APgrOrWaf/9Wlmd
rozI/sxpJetrre5ibIfusitTGJBJyX/JsgnQzdThXx3ajia1TZiZLhq4/Ntd
PoId48sUANJWE1CJu/YhigRDML/w92CFGSqYXeGdzAtWQnaQ7a/spw0gPnIB
d0HYci8z7hd31qrGnuKZkHpjcypk/DGCK1paH/b53qLuYlwHY6EsOnvV8LOZ
wNMSQbku2H0JtGL1fEbvScv2TAVArhuSKtFKsqHDyHIZmcByFEbZJAMhhrGC
vuiAnX+ws94KxYVoWJf2XbS2cobc/+beVm679eYmu4j0SteOSIAI7ns1S7bS
7bzCQDSDC6NRFNoWPU1GrUo3kz38CBNjvAof/pxtb+2WLbzpP+bx0brDKbLf
1cn60LTfQ+F+w8UPyYw5wgcsWdMjGTTPN6pKtVyuVmpOWjvVI5cXwDSJn3b7
q8E6KWL1mCoBNe07sBsdwdiE2qj8JyffGLfwf5Ve6c+sKHnwvAhmB3hXGo5T
tj9p7MLZ/VwjQaFFnZadMOamDDw0w+eEPeuwyfIJKGkanhS4RAB58JpSg4aB
wS1HpJUf+c6eeAxDNqcPuR5jugs0TPBcEqBNGdG8nyMnSsJCeBEj1s2XvVmx
7n9T0aE9z79FzoeLrOrymt3qOZaIlUwIsJHcdJNYld42Md3/5ew6p7ZZ+T5U
AvvdNAQup+P8qlUw/7u/ftZVdYlmweH7jHR/CYmVR/7VDb+lyICV9UYlOngg
7pOdc/aP2fxVQePVEo4XXQ+w7xZNaQlHXNfLhPn+bEJH0Em3q3Cl1R5/ClQz
MRhykxyUgD6YqZOrGx9Z9UoSJ19lmhc+CdJK4ovaVrEea95Nj2Qhu0aa00VY
AKOl/KgVmIzx2kCD92PGa8YEWdFGPbl3ely16W6HiJ5/lB4DEhWdK2StLZip
PMZwwnwdXKX9RLFlQ6d63hOaMcimoCIgHHxYyqJuJIGwea1ESSxYL3Td92vH
Vzfeu646oxE91j75kEKOyZMRuB8/dXlMHCL152cn8rLrw93DSv5elDkiJbkg
2903xqPSndlL4b+ReA38D//AvYTJnKISlVUHn2Zw1hsdXOHFh9Y38ugRIxaR
CNz0zijZCDqqQm2vvxvLxE8RpKpJ6yDbztn2XM0xEbXN0Z0XWoT8uPm86aLv
eCm4zLkDbh1XumOLWoubPPfA6yeUmYls/xg3J/wxAQMhvB3EK2ZLlZbMcsT/
JWoqkjK3/Ug64zeJsnOrx5F2Kmw9FfLeecOEcqF76phKQgoVlBoYsz59kXoz
xWBn95blZ0gI83wL792IJYZknPTl9Ng0yhbzxHc7c/snt11X9M7s7JIfTfrE
tvjCMAKY3KuOm47NWxqld06hCz1UdzM1g438S01i3E6NezgB7YJzGEVJtwha
bck0JfRAWG4/wuennjrO8uw/9sGfoqYJwrDIIxGq1NA8mk5pHqwU+LfYtK+O
2SLloo7ns1Bul3+hmK9edc43clhANTSXj3DVlFxD9KLkd2L5W64MjjJu3Zhh
qOsNJCbJnSRlvy09VptlAJpXgox4mNeM9fleKFMB0Z2hAx2IGyCKNQG/THNq
GJLMxg+OxI6ibAg4vugvcWk1nFk8dU0nzIVsq3bxlAk/YPDqB0tPsxmgvUNh
ZqqLMHl7qmYBxVtBul1M19QeSsZVvmUbTVI+cX5p1nDOGpy28B+ntzwGF4G4
14Krj2A8RGT2Jpy3NjS0LZetJY2jZWj8zIbkiEogxsYg29tVgY0GiaIm8IeU
97aj5BJrh4XghXk6DSzsw1yE/X8vpHnLZiP+LD0+pdNsIlOYTQ6q4cqN93q2
WEHHoZ+2UdroSZEkEnUGkcHPoxNmCI9tHKCB5DCFqN1jK2ZWiVpNq+wNZZB1
I7mEdSwj8mAFz3qogYQUJK9wiDFOep9SGzELaJR4P5budNCluBprOMvwysLK
Ya04uJYKi24jJzSg6iMajN/TPwzp07ONdcPg9e+VQ2NMBpQAwqhLwFJFyH6N
Bwx4drzNxA6Qflf3rxAWEN3yaJHaAuSXR7lFpxgnrvXomFuIWO+PvcqY5RR0
z85RTYKfIDxexOC7N3KNTMIDOJhsosInx8jZUbGa/7DNtKmYppvpD9Ln/S4I
RWe3UShhkBASave8btSSPpsYwOt9LwSrxm2y70oC0L+m0lIlkgHH35J1C5sC
kNlhB4tg74Be3RyDh66AMF9/cim1N+c9o9yREZr94MUEXSn8IXCheb32BOa2
Cuql6lmaZMR/TbNv+1SZDZYQcpEXPqeQMwGaPEwopnr6jABH9G8KpkrLYZy2
YE11tSbJ06IDWnv29IkKdoHJfj34h8hJDmgf5VMWAQUqJdKM8xdAnwP9uJHC
nKOkOWZzgV/39L3WeijI2dVXHZcDL37sxMx4XwSFOPtC87dpJGptteLorfJ4
yzmFeD1xaRXtP5/TeVSYJSOQwFZWw29NoJga6mQ0fTFuIqzp6CghQ0P6+NGX
8cdi+5AFCxJQDSAJP++jWc9woDIR18PDhoAXqnTupProgZavSauf4HtfEuMO
5RREgfw+i7PwzG0mQ1xTIF5SZ9+ABtRv6achjFwKW7F4SSOlEj5p48To9NLE
1R6lNh8Y0vI2K2cm9FS8RRuTvtzwKLbjD8fllDjqNFZoNDhO9i36yztLkjPw
+4DaxQbuEp0BsYDoLdmOoVqB8OCaLh3VzJPLRnnAo+KvhtgMBirsAqWpkJZT
mAOtzl1FOu0prMXLs7AxRCKlJNimIFoAZWt+Dvy0uD0UFqIrPAXtFG83cXYi
DreD0gHmbfnTriWg9YRWoHzIp0wH1kj9kNZ09QPwBu07uQQ7Zs+DcWE8QVc3
0IxszpjT94nZGQm6kt9J8pqkeL01GKFK985XBNdFu57lETXvubtM7yg0OxRs
CBKzIaYL6EmxLKxXpW5GN6mYXaUMeeyp6FFSFgAsKRWKWB4Or63z64WVT94v
TpnpoyPdxXFn/FxDYGKRVUUCwo0ZhmNCeYC7+RSmCKk7vihHHZFsuoBc2lVC
pCOoLq8nn00sc3gl/k6RL1xqrugyqmOqJ2b4BHNZfp4X1WAWm/aWBYtqflA9
nQyFwMf2B8WSi27sv21pdwbKQa6YuRkc7KZybauDuTzN2Okv9lnXiB3wpW8T
GIYir9N+qN2WF9DcJqOjr16BhcHNLsgE6tQuxJHtujA27y49LUdAw6X2nQjI
KS0s9/DCheU4HFQTyqqOK2gaYCdd2pJefueZBXp46V47xS+53V4q7q5hdYRB
8+6hrbQTAEBX8J67FP+AhZNOcHuZ+l2LBje56hC5hQP1S3Dvmc0EPeLzuyIg
jh8kk4bgDBcn+SYZcYU5TH8qknILhGKru+pQ6w/x43E74ev8+GWXrgHLGUBK
iiq4I6UUc1x9VyY2DjF/WM0lKkhnlr2OOOzhqUzeAJpuMBYgERWendjfdiaD
00MoCHRL2rYQQg5xwJDMwOu2FmTFGLZGsDb+IRf6ATLeSY4JJlVtY3CGltaf
U7RHMLN6m6No2WvfSXzdK87s2+8dFN/AeAkZCJ55zz1atkX4Zf7uFU0MqJP6
n4Q0l/c6sf9l+NY6InfejoTIZLAQ60DMsEYQqIuLKmgt2QnTDBke/pDMPbsV
bSQpoqf5naEWIy5yS/NSIyVIl0n4E72oX1zouTXaaPNucmccTC8vQNhQ49/R
OJSDqWW5tmwcGsjq0Op7JKTYXkvFB0YqUdgRcFg4dhZWuyJsZUcjxZhWNkW1
kcV/zdiXvzBBZmDahb9czGukYEq/6BF6prr+OunAO4YGcxrJP2XKHF4hmpOF
+ykpDh7VAkzRrGD0tmQvkYyX63pJYl1Rr/fwi4ja/U7z3Ymk+j5A6MTaXGQ5
Y/3qdnUwth2hSpr4WLNn5I1+cAENwj/mInY40Nmj60KlRVDiG37Kug54dQTz
/YfI9Oqa/cRRc+wmFgtLmba6aFFaFogvoUSdNNJhDxhGkT5kPybwXnkFQULc
UYb77TFCHytpEgaTun/fhDU3s8GuvNiUb49NnhEbbniDCryUjMrAo081BHN7
5YjXYEmaksCBPin1vSZ2KYiQa0yeo/DcMh3pFwKXYzeEkZ4FEu4rfJmfQE8g
kx1sg4s8n5bGBfs7k4mXw8xae+S0XhBlID5kHnT9R2r/HcrpQD6v95K/Wn0F
OZM0c3m9cHozA9rscuMczyrXCsriuoRPdCcK1Buf+6bucVxg3bq0qw35sCx0
+ZlefHhZ7+q4pPVpG5TQGIYUuyKv/ZU0nT6bxHx4yl3kYn2g09t7DrgoSUFa
AzwXcvOsIpXGaALe9WNUnrFf8iBKAZBLARA4yQMEXomiYzOTSDyws/4tfITy
yjWTfe97Hj5EYo+SDXkVu2Ou18+m/ty+ShMhtyu709ngXJfY4eQOQIahVjrq
SSl3m9W8ryz7WDDPyJTjvb9ZTpnb/8kWL1cO4GWc9RWIcOk0dnaU+2L6H+vA
7OplsRyZJKA1LeK1DTB0CRpcCXuUf2SBSOZxO/YxX9pPJVpth+D/IcAF6OAY
aLdeNxsSFjFx7NFFLe70hyxavricxzRntN6zo+N2A6OJL4ECcts2ITvWxvSv
jbAXOXmIdNurR0FLYpeJhFoZRDd2EY5AGBfF/ReEiCOYJBHqnGcYF9lG1Q/X
5xkHr0cwCsaz9zMx1rm09aU5F6VZmdUCFTOHGuttxJG6DFcU+Wwnl9Cfr68h
pdqL8OGWoygfhNjd+GVQ7YA9J+NBzxFXihGSA8z18GT6ewRA4dsrgYgcjMQn
J1vngq7oLNeX+G+zKjJF8o+U5XxyJNeAnQqVjGY9Xbo8lcJa8xF+GsFaoXoL
Kby3/uG6/oTfPkTq9tGOjcEl/N5x6RfNSmkNUjLIRvF8vAYBeH/Vhea6ooM3
/dCRSqIki4k22KJQD9jhQ/siWe3TXaxPKEMpkVs2V6qwOrFU66JbF6R2XANB
rLQOzRCROfK1Nn0ruRZztEyD2LoXLBlahwUe6K7SWzYiS7xojxUvVmPKRtFC
GaxVeuRrUDLKns9rzHxo9fNzFpR3m2f6Oqp1FkMtVen92z7osVpJuDZmgeXa
58C6cmJkb9kjuuZo7bZBmQQvjOFUNGknkRsCtgFf5g0vEaNMe+QvKmAswGUp
sJaq6kJWIKgTT1chZfkTVmXI8vfQFzFBCz0GXEMjceBVf8+7SLikI4L1DFqH
BOxWHgxBV/GhoswlLsb7Jr0Wo1Z13ncxElrVkIQEp+Y1se5XQzTFLCBWwBy1
sp/Eg4JN+tyUwaF4M6pNAYBZTV7I7lgrOv5LShxwd3JLWZLBAizElmqpjYne
XH1e0V5F+MMjHiSFlPi0yWKGlPbQsLpiwQ1vrhxkZTL/ktf1xgyFMqD8XR8M
FBah8NT+H7SEr+EEmPs951ftu2J8cTRZc8dyoHEO7wDF4p0vtUz/8xxhIJE9
Vr0ZH/yD7cPP3AYepfc2ku+PPSQ3hUez+ZPVqZaNdriE8DljNxYece0IQY4H
1l8x+pboK4bGHc3sV8Et+ycFvXAHQaD4KSv2gZ1ECfXOsSRDl13rrJ31iVyf
1HZb6zpKS+EZhNmm0HN5FgkP9gZ7t8mODymMclYDjls6F0qQ4S9Yyo8P+ZeJ
Mr9WLoc4r/7Mrym+tCy5QgKyKS+2pHb+c5uzRVrMIKk+xkqg0WINNSH1enQI
PU2gVyTIbBQcHrvacsPj/ACcUmHc2FXIH8HAJxDWQJYNnbjz2qONHaktli48
fK20x/FLHreSdhOIG2k0wEEPS38aIwMOw57d7ZNAnNZLFk+0zQrrRCEHaNWj
VxyPD+04q/i6t0vMvXjNfOZH8DBTccD2Vf7ToteeGtWg/K55DSW+Ad+V95rN
DZXSl55a1LKEgwcQjWD+AeJbkEzbjMNF8AaLxUED39Av7zLkTxosOnZt8oEW
QNeF/Nux0LW2Q0qG4uJKyKWUEElvicrXHDyyEAyrYhr+5w9Biba2k0YdYMI7
hn1Deek8z4E9ADfIwsxBc7biayPeyu0hYSu9El0Ng5/EhoDg0y8jYaWmxb7y
vlXXQFHykwji8DUkY6GbgWgoNl3Zk0Cx9p0tTW7iVQ/5eDsLF8QDLXOwP2Yp
AAzMvwm8ZCrYxYTGhIep/4ylPHQtY5UCMVxgMuy5095Ol9EBMZl/KAAKySYH
mu9wS5ykgvhBU+jr8P4m1GjhERj+UMqFmrqU4W9hkKBgqiWUzh0J5hi0VOh8
pCPVvOuV6RFc+1p1hMj+wFHE2zecNhjJKrciE1trJY5SkOOB4lvXNkxV5cAk
grnKJmfh2t5phCsjEk/weaDZOeD2+5gtx3ETjiS/mOrCKgSH2nj2vipSLUAG
z6vXZgEdHNZdl+adEMVeawa9ExVj2qss1JbrX4rdN5Bu5EvstcGtWiEgaZeH
ewyo5CC/jRyfARTqGP0XpqnTvxXMFtqL/gNZICx2Htcj9/FAsICSkCUensJx
T5+y6kByUcYk/toTTr4tO8W5DYeaZYbmygDjbz8avcX7oajL//Phj2Ur69mQ
LVU4Zlpv0PQo5S4fPAA/q132szS+KZbA579q2e1S7Ygxvutxio/rLv4YzBzW
bsQf1dWOmfC8VvfTPDb5dHqeYaESofnjETv4F4xBCMEvmcSf7YvF5LviBb9P
VH2kYb2tfLzW7TN2dst7nHB5aL707tw95LwlR+dE94A+Fj9AV18ZLNTn/eL9
yiZFkMlsuhLwnbgzby+pRHzQbX5ostKOAIGS6KCnATLvuh8ssPQryYT1Img1
S+nLrCv3gkgyTCnh26RtXZ7Ft3A47FcKMmxAyYIMHLbw/zall5MwnNX1mhix
ibnItxIwRC7K0ahYQImmkjJilzqO4i4Td/1Udib8d3Nebzxvpi6FOuO+sDJ3
131uZvX7PT8IGI37GWdXCwFBpjvsBEUHtvGeGV7Xz7gWK5WWjHr3o50OPxbR
BTIl0mSX4JqCl6/eB8B8VgzweQ45k+XDBYy5axkL4gLgX8Ht8rUjzq1Gc1os
lmKfgT1UhApUjO7cpv8YG4CQcOfKO35P+674zPGKeMcbq981UqdSOWW5V7Tg
QVjgGIvDKo4CGjerGqAt9TA2Qak1DUM0C+/bX7LwpX/7s+69cbJxdSOmMMy/
NzcFuTiXBlBi88xyHVQUICUt10pLTpbwkNLbQxxnBSVNRwiVjvE/U7GLwndu
S532zyRhgfKUuVWYkc5kgcWj9ujREQEbcmS/OiltYScYvh8x2WDmLI1q/Zqh
/W3a+ZYxCOCzsenrmV16vHshRJsFFCJXM/8EIVYKuB7AsJVsAHds0knkNH93
Kb9BbGzMJsWktSsxjYQtd5GhV3qEtfDiDChTSdCr9Jh+3eQTr74v6dCyg4i0
h23T2Wx3j5IBhtd93Ue1dwBQGId52evrIoPF9+wSONKss5KppGSRUv+qH695
WWZuVRmGp2qQw+v9pzwzGFe4yR4vfcazr/6IdS8ANELgoDtUkUM3yAOxG42J
HRVSPpzqgqUMKW3/FVxGfCwUYU9TOn2s6v2ZeCsRNnOw4Nk0e38qoHiBREax
t5uzuO120dBBDjJmHNVAH29ss5G9ga+S2IgL491VIw4D9gek2aKsKJlN5gpB
e/oLsFu6bvIcIcZrwlJZ+4+oNEvK8wYGCnMf9g5G43FPVYc3V4flb4rM8YrR
MHrhhBkKrIh9dbRVzCDvzqsa2uKtBgvVfguCgHg=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpegZBL4/wSSI7PGGebvPn6OnUco9/lcGLQUmKPWhuobugiKuRGRXVVtAUlAkvADIEOXYt22u002sOq01I9F2YMPFT0x8t91g8qwC8xmfCuwPj5BFj+w8SNBn0gngekmOF4X8jDmCje4rx1MZ9KgyRBLSxprCF6xIv5j5SNElehqnyfpcTEQPuRGpFCtIJpl8XEbV0hch9hSmMA9xpQzwHWIHuu9FOC2TZC2xY2Grc4/c0QUtqdQoM8qJsxmDkC3fNW0lX3K17cYZI6a5h0t92Iaa0nPB6omh0LS//n7un0UFGZuoP66NNbdWdvVdOwOFSKpxT584dfvGv8SQPWI0HVzZT+wlUcXEeqtQpRgyykrTB2pQ64EfZEfKdq0hgxO+mD7sVA8kL160dHj3NuQ1VFbmy73knCKUdy1Hv1Zq1pPBhqTJFYVCycrG1EzaOVx/WJNP9KcU4LgW07RlOkwFQUNhPN9UcvDN2/iYtqFDD/b89GgkMcbUKBcjWAFXluD4Lte+8SqNWtob1bUy4sopPEn7ajaTGmZ41tUNWgdrBP7Y69QSQN/X6RCb9BdMoxiLTCyD9Er1kuJrFp0ZV2zsPfGVyZDtF8SkgX7I02Jbv4hCF6MpB8G6EGNCmef9LKDG4GIrwKLkojOFiqpV/x7DloZCwCAUIPLRPrdyeN+VU/4hN+/ABOgfUj74jcbMRSf0/fySBPN5XhQLl2TyTGrDDCVUClAJKspj7NkWqHaM6URjX9xq4gU8h99Mr2OHG3QbExgxKaPZ0XRWdLJkehIO5FN7"
`endif