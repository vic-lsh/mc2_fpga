// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZkuMSisQSwrK5vVnPCpNNonpsijdjYg5QcGkbn47xnHGhcmpTTADwSszSo1N
PiZzPUTRUkZMzKDrcAbpa5NxB33xXCIHOT40479yxqJOyIdmrrYNjgMEb8fz
4tYMEk2aHbpM8hcKvinVvMf6I7fyZtQWph1tWjsxPF2dcO+DUPcU8002qkTR
Y49K8GG6In2bbIP3QCk93zeiEYmzrDiccYTVlJlu9NH3IW12Uz5EXIf4N+as
UQe1G/YJS5Q/JoDwCqmUmSEmsYPWBYTsQ0JaJel9OcEq2gp7z2/NAC7cYrz7
95PC333lw9EdRBOEVml7Hr/6UyEyzgi6xPRaASgWnQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
E2smnmSiL0VT2LtZgOh4q4s+QngxOWCCcOns8/GWLkF7RVWtQun059Ql3XZp
PEsq75gyHUAndLi9ExyI094Zqer6mrvidmONy4cXtqqwtewX1L2wAjUr6DOM
5PKq1q5YMC8sxxU0uAL+UWbqa0KY4QF2zgZal4JOHCnEnpKpnakrvyAJIndA
OWQxeN+0cDRdps/Pk7Jlr0MM/4I1QYg0ia5I3x7WvZs2/SjiWqMPRqSDHgl2
QEP+4OKMqEmTVnBirX08l5Tf8I4SrM1CrY3jlKqljSoTKpzPXeX4t3YrFYhj
7gFFuaiUDk1omcQAUdEpP3/LRxBFQJXlWpJJrXJCGQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
sVRMjI0DJ6dkMEKCGxkNF6/p4fEGFI56PP1D/QQTNnWvRMpGx1EFCPn17F0K
h0XDSI3Sd2Kim38aWgaSdYRheMBp9ln3b4IHFROVG4I/td+IHnBqbgiZmY+p
LYy3Dg2U3RoLRDUThHRHS+nl5BzvARV3bhxNfKR0oTlWt7HY2PpB67o6ILCV
qnIu+8/o88lpFgYuJVOMzCz6OpGKvp6AS6ZOQB+QLeihcP/4rN8i14pceROK
zZcwiHDhaco9U/dvXNZ++UXNwuB9a+iRSbc3/e4aAJkc1F/vrkZRSj27GyNw
2N/dAUTcv0VdkfAn4tp/mOGv6sWoBndODPjdSAo2fQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cVsQrXW6Qi3JgkYrt8l0i2x+n3gvUO4ViD8mEKtLigWw4jGVFmwr88yiF6mQ
FbQyfxJ4z9NinmP9p0ergptljzki9K9AkjAzINUxDc6+Rmpiip5OWgfYfwkK
7SQ9Ha/kgjgypSRj24GvWUzs0qPZAd2DQsmlyCQ/jumkTkLHEpvJyx8ojJ69
DqNeN/sB4rn5kBgFW2S++AqF6YQaialSCnjkNfEzS3TNIxczvuY553ZqfPuV
iUBS1R/4D2fH7R4WlxjdG5Lz1VSnIseNPIkYgLAqF5QMN3i4fpqYvtHo+sNv
/+fdqJVvz5Aw7n//v7em5ChevjRCbvJEeJ7+DFIUxA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
h4Kywy+Z8ljLFMe+48wggBOOBwBY1QJ3RXgj+TXkqu6IPnonOvgi0c+cl2l6
x+WraTfCmvV6GpZp9ZIrqmbktvXb648k1qpdglWGMFpXi5bUfmzcD86wG06W
HGdl8e8OJ/vjA6FWxC0xW3sOHxwQvXdy1aJ0N3MZcCg6MXheh5w=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
qofJxN223idTHk5Eb4cH2VrM3TL1OrWoOE3Bee+AREdOinPxBUXp7vh2IQPP
NXb9UmPWMMCSdVtqF30gxHXnjrajaWgzrL9Iqy+eTXZ+BNokyT0Xiy+R0j9v
QPsrOI6PMPCZTQUeO7CP9vwUKrgmaGLF1L7WWzPslfruJsmA39cWu6mXEgHf
r9UhZsFTfMrPCJZGWUzCMQrGdtxgD4Dxs6bBpsTPqgoC6knMVp+Wc5MTYCMX
+waztNgAMDiVj4QPqFP7S5L1tTiD0PC1FVlsMJB0JZ7/odUKjh6mt6Ve6qDw
r86bIzRGFTlVgReEZkSHbaS/d/61zk1NhfEm2pQuX6xueW6gDCSK+kfOyxFA
RWiITt7EjoxpKk50a6jiKo+EOu3G3aU8O5cbDL/9Hk/Awp1jP4E3DNYo8Tv8
zl+jQ1aomC4J4wH7N0ZSRR5v9GpVSEbEd5Gm4yWfscGzQo4lg2Q8XgCmSVwd
ef5Lu08JmEVc611tufFFHs8ciBWkQ3HW


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tbYC/SXpByk06LPj6BHSi+xS28f+vCjB7l8N+Xcu63/2IzUabuxnsr0tJ6Xz
ERAh5iCcxB+BkwQo/gLETHulOX+Ggg/xBaWAoCMiQD7pXna3KEOeTobvlh/G
oJRABMFWAYDpAZpD6Ca1aRA/WGONDTilrC08844BD7uckGxIEhI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FXjPYnAKLSJZNLxyvjHYE1/H4hJjn9ya1fnW/lqhPuqL3cVnU6+q+8kpwj2W
aEixStDwE3U9TtdZQn7/e7wjHBIlMVxD88NMMgaSaqCVIy7ZGNsmfGVaTxVB
clqm+M3FrBNk4KlyjAYMMd9wVt+sGJl9LAGZ3x+FEAfIN5aR7iM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 18432)
`pragma protect data_block
kRuipdTzCVr9ENrvEdhR0YhemxgYI9BhX1qE54O5NoEuYPf1Ydw37QR9H5lm
VsPVt97CHO+ULyU7QGUXFNxen570n6VpxtwgN8WuaouZUqj0kVjANf2UAMvI
p803MqjgD7RqwKBqQCBsI2b+qWbg65YBt4/d21hbUhIqwLXKL2sDZP05osZL
fKg2TBZTeI6eyWQV+B0nUs4tTozq6k/tbRWD0J97TM+GUu43ldz5rY7I7cTa
dfcbnikCh+kiiehfxb1hGGfzUBx6jPHqnoudU7KAvoXLDXhzMXmreVDgyfPZ
krk/IH+OBR6VRgl5OHPDmnrywiIxF1emIgGRBf8BXgly5DKeTQe+xUrogYj4
msbiZOFDaoZwj0JSSXqXEJHy0PfT4Q8FrJYnuj5FFrS/2rR8zMX9VzMkUk2F
uGjEHLzo/Xph14xqQkK+kRjhrb5hIZ1uiazYiqTxshQzj37AO2xqgJ+E8H5P
5lSdcMgKPrZ10kLQBqbZEP7ug8+OEMXyghKxgIGMqMZw8qVEMKhYEsD9leZn
g4mpNAzwmFLgMHPYbe1AAfigKElqsNMs0U/rDQZVUnCfJp2DLVqmfkNCSdq1
blEhNY43am+zTU3riH+ASWIGz21vvDPB4TeeNP552ctPN1ciEl8uiwL2LNbX
/cHK+wToQDJNKU2PKsKqh50TRjuaBtTzH8CHxrq2wYj3wJGiQxn4LuvmAHVv
uplNNxYuVahJN6ItfKX0vIM9fatH4l+oTeX/opBmqzixGrvBIq5hPJT/6Swn
zqraEwV83/Rn2aBchMfmGJfzkjBxFaVpMzqHQ/pzW2B1wCQD05x2VlBFj3lh
pqDxXtt/wzs2lvfmRHAoSDWD2tJ87eM4j9E8sM+8+B+E97IR6f+34KZaUrWp
LSDK2sarTMvGBbP9rStJrgm1Y+MVpqg4kVUedrfs1TeGcWHENKcG50vogi37
8+JVZ3q1IwfeyperRDTt6OCaiO74L1kiJ5vUzV0XgORp+SFdMBEwTED90ihR
7ZgfIhW7c1ZoiuTlzWHMrPDGDW957PwrvDkls4Lpe9SOC0LbIw7wU9SlBBtB
OL1FtGKhX0t0T76wyGslN/YixY1//8+GZSMctUVHyVW0gn0aQeIBogwb0UdV
eE99owbcFD8HVK5jFj/oXNUw1ZiizIc88WkPwEID2UD0jDWSih2swQZaWDS4
UcaQqchLULjWNv+YTWgUd0d/CxmtRP/WFHJNzzufcV3KHs98NVvdAhoe2LC4
LMOgLm2eQR3BeUmnzboOoAcn/t/iTPCTxzY6/7loFJE26KejkoAGHXmhBUkn
op8Ng/3j6rhYpEkri7WAr9NXBQeo8DCAOaHoDQDwc2BXksemZEHaVOzJCm5Q
LK6j2xrPF+vkzZfyZzOqm5NMbB0gEySx41KPw98RPyKjJgiVmseCuuLjFdo/
rxLbGL408+crGKq2gyftRlnsAvw3hjDZmKyAmfpa5UCGIveAucamvnbUJVbA
IKVtDGzZBC+nMATuxhHwGtB15nESwLeBCtcpeRTjOoevtF7GGAtz8rKraCCV
617q7oWpkvfe9YoRUqC1bxCb3V6WYvfnLV4QcjIrxRbkV3Nq7E+dC8cKwCve
Pufyahaa2f+Z5YeIBUSjCHl2I/4o4b5em7oSI6JrE6EXPTUJkNwDZBJTx8vH
ggOdDzymm6H6tPVPbOkx81bsRjXs3Ue1cB+4m+zIOuT4ZCNbYvmHHBHGtoav
OEdkh2eOkXNriGtzeyIFsLnZd/pVbRKcHLvBVWQdfDIsP2+x8PduQposVuco
qQcGie6QUC/si7rqHWfdIZUPpULTKgSQgfOSHeI5VTQguKX1q+TFNy588dHJ
6HZLrmbWVrDGQpvX5IbDHX2ok/Jl18BOfT7kX/HU8lwlOBPL6YGPJ8gQK/zg
EIQOmGvkNdGb0eHcqA3UoyI6RYBmDnWWCAXR/zW5D0XxdqEdugNjGjtVTv30
aA+0Iq/Fi0whQ8qThWlpH/bqc8pxOK/QmKP1W1Q+KNGCtnBydxK9Bly99wvP
0xvj8dJjh9eaf9uicDzdQsBeiKA37IIBkqOca4PFq5xNvwSuRYW+1g4fgFZR
R5JtgWWj0R4wjOy0Svs5xRZ9itaslcj6wSlMNUHjVnQ9ByDvzKT7B0yYdQ5M
fxiNuyA90fYOa1FTZQQuPM5tjuFFeusLwPNPuSpeRWQuZZecMk7njCePMKs2
dn7nhHeMrTjb0QbYYYKrB0b8SV3ad38UE3WCjKCexmDHR1uPFM2hYrQZ37s+
l0u9knWvmXXpUpyktvhuJdRQddQ/GEi+Eb0WE/E5SQ6lxxYMK4EpLsGP3GBt
jgwTUcL+dV5Xm2BxsobS2/jJMk9EHbZdXWLxq3G60Ms9Efed7s9CHyuu0E/X
IHC6LjfrTWSFDrF1SdIRgwcbiqnMnbUKAlEF/iX1cFNSnkoAXFUu52jXbVWH
yOQ9VBJMoO6/1VDC+JJ/g0zI5HBUG5MAaAkrsil/HIJGfJ0GnDwrHlOGVEXG
y4UT1EVwfzLpSHE4wN/3tju8DomXSpNfexcQhCnKvHxnY5ClxbFRyPHpBdIM
cf2Q4flUhXENO007bWY5usbo/ZhL4dxInYptWfrxC37pspXsqSIXhJANOneT
xZ5MWF0sjpT4c+rYxGNDfPUAElGqd1hOzMHIRXzccIoID5AwFP/WNR5Wud96
m45JeuLDmA6NIaM69AFKbVopjZ+Nf8bwTu91tLgRHNYQm+z7iiuJGkEoLs6o
NUrlPiqtd8TPwMdN8BfKxa1wCZdLVVZDFH7leOnQDGM/DvcEV3tVYkLOwfKc
3/ro4ouRAxtU7s/MmSZyJZ4bDT7+IGG0oxTuInbwoDelbZzgGEqboLt1qD/H
ORCSMj9Ogl5SuRNS6lyZ/5Id+V0RKKPqfhp/OLkHrTrzXwPzPFiF9aG9zCY6
HAVQNQiRkULz4BEJ4KuEJF9REhcBGA/Hn6O8v4tT/5HDp9qgfummmtITAyxB
uXfITQbyaPMnk0v7qAk/W3G2ej3CguiW1OaE5tfaRpUaZzudiGT+XWar1XyZ
ClW5W+PIRLDUvDi3QmlDNd3p9KSqzksKPA2rVIvdxeGQCQtDU5lDZQLkG7Ia
GMx1VC58sBItDw257h1MRuLTQZ8Ivh4ariUbTXZef7EX2YPHAsxFVAB/3FID
QN9IynMV5ULHczeHPn2YB+v27dbfDflWaMrJ3W0PtOfGCN4fsU1a8hRPj/Ph
0/q+SE8+/+W9+PdlUhyhUKsjgyk3e5MhQSg/ZGJDfNUSjd5WqKguceyQ7tdz
vc20M6h+bYE68MuuU7xaJLkl6BYZQmn5MREmkFHF/TQkoSVxKGqe552+SSUI
7xffHCILKF0ONxM6TO7jv0ZzZv65WtUVQl1ZrssBz5ffWdudePM1qnDo8qlr
t8aa/P3XNHgnJ7uetbXwg7EBJr7htc+bGaCFQaM3tg+ghKWfakK3p5qHGaoc
ozXhwbvOCQk7nW3I40n2utSDgU8sRshee7B1dId/nNP6qOI8qJjSsuXb2w6F
kp7zGf8u6UElST9eNWzIQNlOEgw0hCULiv+Eho7AduWgfv9CLYrZE1zszoZ/
rg1zKoIlSm1ZI+ocrFiRBHDymBVcj64xcd5prHWALV1dJ4g+vu0MD0JwTPLQ
NDrK7RVQY22Z1ozE0u29+bR+OaHe7Gdu4+I7rsI+sTj+67NvA/fXie/YNa8E
J7K8uyOkpO5IHj/yIMqflXJA0PRIfvcfXE++NjtOZLBgXvfBcLdEcVNtuO1W
ex4x45+YAjS7yDnVUAPDAkKa+TpbWZNvEmfGy+Y7Zz3bhY1lVDQi34prdGOl
GMAiBh2fYybEmhbxQ1P//iFka3Yl2RYdrpta8UEUEehsbISdKO58x7jEzsvb
226wkKG9cRj4rAo21SUzsg+HvHgBwl5x4P1kBrEywkTRrJigUhXqRGUwR/zc
r8A8JYJcyEl/teEusZq3teoRnqkKkDGYWS8kQifmwfgrS5WpSrkVV6f21wIl
+iZRO3mDuKkcR3/NZTSbtYfkicaR3F19zw8rQj30zdeQ6501BRVle6WRuXI+
zRFElUUklqmiaALXmCN3ZUjJpqNaUPRKfeaFI8L6rvaf0avYqNm5XoGqhz7I
Vzy1No5MZvQsxSXwTeLlNFWPxI8thTMPTq8Cq36Rrlh9Vu1tI53/a4C9t2B2
1bi9Rj220kWIGYwCgfp0xOsZfrYMXsyL2IGcfGut7acPUn1ON3AZrxYYzT32
pv++SBDBFHbH+kvPdGEsqHHRCNQxlhH+spu1LnI8CnszhNQUrEOLBCQO9N3n
vaToHWua5E9XkF+1/QwMoDjWzsVTbGH7sYK8PpPVW2/W3GvOmY2uFMLyMITh
9j0xjsmmU+6CioPG05+IYoiVqZwttoarkzuN7sdkLQEmamdhlQMzE6xgd+n/
JiGGm7BNZefdgbL1BuwWJ79X3WnHjR+llpf9+OKJTlFiAx/RjXK1Ev1gjPyn
RJQPS4uJs0f49ZXAOAjKxeo3AfEek3bMVCWRTbV5P56KICix+lbj/vPVvN5v
ZEnKpy6QPTYyB9uWPuct21dlOUXCGljBFzXIu91xQUnWF+wrqVgKkRjyaUCA
Ap9Sy6UMtXWYd6b48pq7vlpGfRZxdzbS324uQcgI8GzKYdmsTcyo9sffaQ78
2563dvO/V8cDFBfn7Hk/v/SGkUjwvRDUb7qnS97td84IDXs+mxu3ZzS5RJDL
2XZeMs14dSchnO9X6pAOAgDZV/u9h9YETGMpnOndDDYxaJ5Ado07WhXbiBq8
5BYfyBvDGaTn65hXPolPKy0xrkKSvPdwL7f4ftGpNZEMuih758Cna3RFzRWe
shbDf9IQuseB3ZXPb1m3KB0BHmTawviFA66/TL6SzwJ/ogdDa7AIWbczaCrM
2KPiLJ1AF0yKSidj5Yk5wTXjvp1lBBwUaqaY8pxE1/Xb8s+/c2z0dvHkopAJ
bSZctSkaczZxRb8dGQ/i2WZDGEzD5LI8r5Uh5txir2T5BYkJNfB68w41YHm3
Sv5J0ZrZbswFuHtiJ/2A2G4xcREXNev2qQPeNvYFYZWf9ZCyU656AZnxy1Ax
fgaqwwQIVOD1tjBxfBZiaC+tT+KdQtchD0RBevx8lJ02lfXV3+EEAxUbcT0B
E1vBR1F2uvnLIQxl11Y+CoFFEHSsiTR8k/G6OoahjAwJCiEX5vaFPIo7fCwk
+JGx/M549mK6UT60glwjAvEs623X9/6OWnzk1CDwvqSGAFqT167j9okFx0VK
20ESZEYputQgMu39EgeTmFAWCo57enSpaaQye3ToJRO7SSY6YbLWbj3kJZl8
TxhpjHs82J6L9f7TgO5eX7v9tCdRpGAkFTb+h2O4Lnp9ZJX+n3Q53ZkJoaD2
ZBERJAscZw3Xt04kAsua/qHOBm2kSnQKELP4GKDKjMr1TSt8TX30xG8B0DED
a1x30tftztQwe6RHg0GqOvszDJMjeL6a6wyocc8/2iKMyxtpeCwDS0Vdrdih
qcs5ew453Wxl3+TZ+xVyBFGQipBUpyL5o/dDWPVG+lddOuLT25ppSPu26Hkj
AzIbmDlcKAQOP8lrCw9bcxbmdj86MfoX/JStTfTyrCydnHbdC59a04y75Kr3
O8oDerUd0Igo/yAdmeJCQOexndDAQMtSctfcof+PU1h8r1rJjNE/OhddHBaE
UplMEovj0SNv99+ks6D5NycQwYzbNyeP7jsQFv9QJlyLvv+J5jQW/iOLHT6E
xuuwBJ76+QgAu+NMOKBvmVmosEwpHDhYM3BTtXSL6ndtGe16pxGHJKyrgcgL
Y5IhA77eH8WA91R5yKC4+PqFJ0JFsSlwMutOFYPRcJv1mSBBFPz9KHhjGjUR
yuNNWxYDHDRrePEWdp7nCeIiOwa125RhSu0Vf2w+F9D01zSMxQs5HRZAzeNr
jARZ4UHBSTAH+vFknuMaERks1qXU493vHYaH10GULOiG0ieQxTeXuewUYmEM
IhtjkZ4dRKy8T64g3O4F0p+ZmysfVLambQXwOw722ghzyWlFljqk5zG8LDZf
EKIQLXxMlw0FbJnT+lNbOKrs8Y2cQgMAcq3z5eu4GyPNIf7BT4bxP/XHNvLF
D0vRNvA6VKhwAsFLPEUKHKps6YemmKVifcpEh0CwECV5og6xyrNKJu/sEbg/
45TGTZ1YuxmXtarqtTGkg+oA7a3Z+Q7IEAenI34fE1sqCfiXKRcwFU1A9Z2w
O6eW747yVYHzTN0/czva70LmPZA5C2U7uWZym8twdV3RX8GGkvQej1ZJvnqm
/DumWo5wheVVKvN0sSSFnkUAf6DpDxqH8PGhvytMyv2oZp4IirqGWOoOXQD3
Rb58ixPfkLO4tbT6ycI57SKNKsAboJx2d5ebLKUzEP2/WpYLmkptnlFlWvVU
evNqFdLGXaWf0jCHtemUXOZQhjj7ou+n1789UCt9zvEkeCWDdD6bEwSb/oxD
1DhA67PxGhZEwkM/7Y8aaUSvAYDBfpbdlkVL1CH7lnlSaz/qoxpB2PZXwrKv
mjCodytDDJWQNZNGgl3SPeaH5i8rf7b3eku8PwOl+y3tCoqX7utaJyyP6hQX
mEePkE0U9EdW7r5pdCQAroN3hy6OXVf+au749fblbp+oIpG4+TJ43iNcco7J
x6RU9d5uVxrzOp5lMsit4d98wuhqf13vvr7hyFNds7WGhPdFYzV3GK4oJXP2
ZWVdvicHBZ46nhEOM1p9Eqd8WX9Vdb1v6ceQ30FRgiyPdR8LQgv7lhLDHgBO
8r5pEQU1LrbGG/zPz2z3aBGo8RskJ/pwGafOLCD06fiBWHEOfCj0F0mwiIPB
W7vo108vubAi7Jk0FMHWlQDOsE2FwflMFYkEpHNsmE9KMA/QozvBLECdEzJd
30a7dagaMYf6lvVnrStHrgOBcdY0L/Kimr7cN7YIDvmGmOuFovCqswypdYvY
RNBe9Hp28YgYMLs5RdLRihPMP7eZzq7DA6FZdgaWOlU3NkTM3wgok8HsM2HH
WjO95iDmNZPKlrf+38FfjoN+V1HBwAPsn2u8OmDD9IIRxohl/6Cyb1lf0YjY
kEi0PdG2bVH1xxtYCI4aba3pfuV9cxQim2svRBLMVtB06whyBep77F0P1Fnf
akHwdiWshcONMnhUI0HEwYCYH1w4/TbEUptZV3f3ATQgpeZUar7pP5wdGdTz
1lH2DvApcuUOYVSfrBvcrUW3PHKM0e1QdhfGTu9x3ucqlQgcId5/mn9SXvU7
k3B35011/WXP+YrWnwdY6hoE8bVFaydV0t0dIPIQsQyhhR4J3YMinRJNiQ9j
Tyt24nC98CyFk0V76UcsGI/5bhZCuPZ9PxNRZSl4aOaJvBSKW2v/lpdrrpsi
tFKTx5d3+GVqagGcBsOdrv4l/DjHHiiYEd3K4/NT94O1BZbu5pfPD6SAE8Sx
uzDx4YB4gICh9Rik3cSZVSKbSRHy50KBPFa7Eic/ES9qjOSL3upiZpAkD3Uu
SvdFTjmdoSyStuXFuJlUKKezSgIP1NjV9zXH1XB8p3KFGlZVs8/evu01Gqbu
NXZ+aIWYPBSQj227uf/SJUnzIphhuIE+O2x0RKMXT7ngRwnM9dUDq8Lzy+rF
qBGkho1BCytjXkaKU8J6exkJuIZ7RMdOCt5US3zBMC4HPvri0Uto1L08TKWV
nzkLte5AQ+J8creFcgYWhGzHUl+3/7qHTBOQ7Zox+GqsF5+yQUWuFiEUmSa9
IE6gV4deSnOQC6qY3AWEM2BHt4Gx1zXXzvc9bgSIukhFmexhZZ8slZIueVCc
0/ZApg1MVeargaJUZLYeDP4i38KhBhcz0w4+NpBBbJQvvPLbXNV6n3l9PZbO
0QZ6kD3gzFVR1UGcsTgK6OdyrKtEc0ZiAqi5U6ulqBy8UlSyyUzaCUibiRuC
fuTEePXrmA9K208WRo855BsjCo5/wFfc3jKCiBIdN4zLPvA7ShR4IKZfB57f
O7guxuBIC54CYbsx6LzD76TENo5JgHDEPtSadtwidpcyr9k0mU5Yh+aU1JeT
SVMVUb5wtpNI2LGKlosuhvSaw4KJY+rTmxG37qa9eDSgkiSYHZ9FfN5bQkk4
ugMlSMmwuGUZ3mAk8/jUMIcmszoldhGrdzpm/XKGH1e7NPshNYd5sPvScNA1
FQuq1+oCKZ0i2rwDu4Upwu6I9cAZehvCA7DWHvUNqTcKkKVGHBn+WaxS7sew
gb++knsItjEpjeoixXTywNHIXQw7UGTdK8HyffK259ezAkbJSrB/5Dp1UBdn
bpWbeSdAGBumLDMXXKqF3lizdFWNH/tsD6zkDmlliH2EHOvfKk3uJV8G2fma
yEYu5qPTvOQHa58G2iJPz5TwlPGRr3ssVxKBgLG9LxGQIdxZoFGlqPh2JZg5
XbhSTayx+mfAJ8pUZ4jvcrwkyBbIcC6aNlvjbreKh+1+fWDnE4wZqyMp6Ogm
py85+5AT/JJORDrJRznIlyFL6SJu/SpedVUIj/kOf75ZKF30n7w+JK2S2y1C
jjnbV+mElc4gtSwaxCQV/OecROOzGnNwet7gppMZRxIgE39e2ZHFKXNefmRs
w/tMl+fdMNNebC8YWDHH5YcjGiX3u4Ab++XGexE7q+oSVAM+szhb/TRainDL
L3Cv7LjZGDrOEbj79xJpKqiQIoi83EduXezC4BweFeJRgehLOFNOAuQkhb4O
3gLuNAQszl/SpMGI9Zr/ywF8qed3zP6c6cKJDTo6Kjl3fL+pTvqCD10TUN4a
2VJUJ45xrHlqOL0BbFjDkgtOkH86h7QwE8UH8XNg/wNaVy9iRd8zMhPjJEY1
7pR4F2yKaECeJ2QtVp0gt64lY+4tY1Fqc/Pj6WhcfESf9SuJo9HWfh/W5T8a
5E/mck73hGZJiw8CeX0rbMkZiRy/dpq/mu0ZJuyhFfz92Lpf5+4X43QEdf9M
fIos7BK6Q79M5/e8yBgJ16h8Rx6WpKeKgzaB6jdz7V+JYMYsJQKToXBy9JDN
7DMMaqr4hGK1+aj9POxrw59sRpNjD46A1hxJaMhH/URUyt/+gufrTyN3c6Eu
8XG/oMiLpVY7x+XbZgS+vgUe2gIHJbw5ayr+GEov2ZnBVI6cP0qug99ExDSu
wU3cCM7Fo/iVO3A5y+bg+Ky23mPoQIZYAdfDpi1x6LVHKX2K8YahhVqFH1Qc
Dm9yUeIZomPWefPhv5jIC7k/++puWsE6bwNbyj6TzaiOdbEWuGBlLxlYvNnh
qrhQZxOB1XBTH5xJ5d1RHv3TJy1GisfI2uPuW9HmM3ma8kxiYnWCzO77Elpv
bMwQdYwaPyoQf4jx0OyG4vQU4PmmxU4hWXmNR8AWcSPVm2flGgXfF1SJ8Rs7
6lQZ685JD6bwHglldIQ1208kNwm7OF4hzL1T2sfL7Ul24eUlzxbQMFoUz2xD
1T0k5luRoHXsy711hFLnz8mWfrzMPbDr4JV5Nr/Aw08dUX9W59tHylqfwKth
aXis3kO2dGMiiVhHbLA5Iq15L2viWeews0ellhFO1OwM8nf9JNQDxSOa1ypD
mdMUO1tH5L/EzQGLYdfC3xF6wVitENxb01Ii202koRT5xX4L0aCPfxWTIV4e
C9yxpOKwhR2SLp20En2zzDV2cN/Ccxv2lJ7EDa+adeS6bK4e/59XKtxjXSz9
Fcoml8oTnsTt0QLBjtBLQDOgd/EBEmSOt2yn1Z1pAOufOyfvnlzHsFghAEE7
Hqpg4HJUzBSJ9xKEdzUA9wq5WDmqtGnfogr2l04svKZ2mj0NNwsLHnAVRCX4
vD/V+TrLXFnI2zRipgd0sjZkwxNEDZf0nAg7eaiK9cJLdx5YGiRY9KWaAiLG
TxkKAsXI+Wd0j5oMEghmHskLtRDtxpVH+TjhiSvLUodwOHx65UIUkQBm8pzX
mYKcQ4ls44F5kIahd+yQQo0RebojHHCDyrO0FN4+bJLZ66XiCZGZo3UvGMGE
OjZMrwNDa0fh+XdhMe9kpcf/RJqbtT9Z5M/mkYY4XiUVrwetlj9u+PNYcQQ0
HtJ7r3xaiY7vdUc14CbbtCvap5pbQWmYBEWvWcN4eyMk9Sng9ioJaant2tWN
J8rUv06yjtcjwmHKek++Lrca9iR511LnCKAzc3Y4Npe0Ea23mFPqPdBhDofi
Z/WliUhP2PgxrjUwjr48+9ATkRGib1437y85L84wZHIBnqgbkozUlcSJEBBk
5z6DtX5GAYjkxxV7Id0Z45w4NwJZRp2qXv3kHsiItaTicv2qlFCMtWEET89W
4MC8PueoF4NfVgJXroJpeHMImuopAjoyxrXQasu4eqnM5lVvMwGJvInkWHzE
aMcoBsi8qmU83rrWLKFEWo4MdHRf2vZLsfgFNbpiPT0p6OAuBxUsNrvmTcvw
hXUUBGodrtsfkGSksJ5RsevNBRBKeVd+1btPCOV8A9mazlb5fWgNIfwd/wRt
fVVYPUKMH0IyW3nRIG0du0nfMBzWIkdZZQ/9FbWZnsDCsMTiPmN2Nd+O2rV8
X4FOp74WRCfBo2vBUFodMXb68QYb2QU0mAkQkHRuyQj2/V14Srr6A9BhWjbM
NY5L2KarweNjbeQ1EHs993Jg8CLMLXXOpgjp5IqvJwEaQLvo2uIKVctXaBDC
8atZPohHu0fH1kMnGXqbRYTkq5RnQggN1dUxEHI2YX6k3xa3CRS95JWiiYDZ
hJ+b9RaXLU12KlKdo3VY4QLiSjnGGs6AsdZKnECfamJzqN81i8pMo/9ayMp0
H1xUWuJkaCjrSsxUjs8BuxhQtj3eMy5iVm6vTnyAhVjxMrKh0glC/iX+h26X
K8kAGOyN72ZZwo+q1qTn1cyeWerspYaVs6Ms+r0hQIPfRw8ovrFKi1/NlC2v
6hNZ4wiSYLhBA7opIY32l4VeacLgpcOZ/Xf6wD9aGTT4MuXF3rJWCFka5CtL
ApufOulCuUz/X659Gn5kIwIE7+jFkHxVa8Tqu+qDiMWFOUXcaWltJDcm2dTy
lZUC+k8pbV8O0TDaDBR7jNJ7KO6i3IaQeiptlC3K4oakjncDig8pWMyeY1j2
xs700Wr15JBPD6FHt5u9zpzOItDQ/yMVlJnbsmFyItmFd1ItqceWv2Zld70A
B/iV1tOhSUzzomq8HL2bECPlPeOFK+Wn3Zercs7tfm3dt6joomWiuwRJab6l
lE8XE1WLt1PUyLJvcJCexvCYfYDJSAlHbciK6Lt3guY2sHkjKXqHODIbwqwY
ljBLchyBj2KZk9y82mH4AuftL8IhOa+aemxSykUNsvvZxfmFaMGjX2nmJi5N
vOAFrzEcpQBYLIMK65ViPGBhd9cuUN9tB5zWdKb1/1mKl+QJ3buTr2iJEwA0
OhgVXhlBlBbjJtOYiyEnlrcZoxDYpezkaqKd2vjT9Td8eTfQkuuwlATXp3wR
s26DtdZj1pUcTxZ9IBeYT56TeeCIEvAaG2VcgBH+Gc+VuvBp8WiCv6btMudU
x9VFf0MBeZYa6unIwHxLu78hHC+evv2+suhpeYPSqdNezv0ZFg0VkhbMsc3l
IT6/z1hihngAHgCHCcoQfwkaIF5TvKKVc60FM3smanp7X9g2BVE+3WoeiA//
Piba+ColjY+jSUEy9cENxINJZ0EsZeJAbb9adCnTQ9sF+udeLJXvJsszIDbS
ILZtgh7WlgW1dC7vbB3Dc/uJ54V/aIWh/CH60R11EOe/aTObY/l0b3CzIbLO
T/kvADqC4DnGQbDZn5+Ggs792gxFa6oGMn7xJ+O+1aH6wu0oTmRyD4VtL5+D
zE/EYhzomiPYoZ9cB9R1qFii82dzDmBZDxgsSa2pzcFAmKFLnhvCPP1Zt+Mm
odj8jpFIRw5sURfdzosFsqr2D1TtkYpqpY977a4pyQxhFfY14NDHVy29veo4
t6YlGVQBvOfALyuXAy52R+ZRJRCcpcfwRwRItCoXndLMPlaXzZngoFxwzVzF
pnco7CIrcIdN/QdJDylxFoSd+j1K7rtrWgt3TVdAm9Br20YsvJPlNpz7JTH6
LZsAsy0os6Z8w3TLNTOb0UvqH+liXw6XQoL3/IfaMoK+J3ymnmKxR2gf3Jzc
vgKFYKcPa+uTk87KaEmmR1tLVGapD+0Yxj/bPOFDXgQDbTfjKC2Ro6ENX9T+
Jpm91B7Taep+WoszSavotZaxhiMThZEAUH0xrj9d2VHD+IwCdRm9zyS4I53O
tZyz0cJyoehCLZokSUPyeMx4jGDmmjyXwQ5UvtdB598k8Yhi6ctqq43OsO0w
GsRS/ycSMzUqVPlfInKvyJ+G6/kZqnveIz10AXsxJNApUUqBmcUH96u2U0KP
nk87jGrqYIwG6H4iO4+TUpHNTb3Wid28Srbl2IzdQp3ZXvCgIHZRNucJ7neP
sWEMhAvVtwia36kF0ZrLXeKMw9pLhkPOVn8ScAT2RmbSyHyQkIe+6WRyHJcH
iUg6ER2o3cYx+GD8SFlUTe3gd14Be5CGJvmmmG1MdHIDEi2TUQMJJ9SHtYhW
dtqeqArDrUwHRWZOgHuNOWXqeLm3CCgzSaA14n6XOy2mHcUMDp+ANwwELE8j
UsXvKIhCTJ6prNP64p/PCRVmSaywHklqtQSEXGIKqIs/XRuN0gGNxAZpXv2c
I7h+Bcl+7L9BLGlIukgUdKgZQ/6W23/YHxMDuo/zV99kKLWY3yXDw/naMqcP
q+5ezwrR7w5Enr+f9lFbXXFlciQFlGxfmg7PiqjehvcfeAOJv+ywICl8dVMY
eAlABmRysB9AqQDAVn5A5+A+VqZ/BRB+tpxYJptqVte0ObOf8FxXAY+2lK/z
E5+WT8QFkUK5dPxyH2TGT3RQ3nIKIKWVCjq70yyxqVgVIGOoiVDwoh/FL//v
as/ezzxVfYgxVedbMccuHeA0Jj7AML/4Lh5PpbbWlXrRqxQWGsl3CpYlIBa/
60IY0q+5yCkRhMSq/zuH80BIwjZRAAKsNY2lltC7fbXeMHg1aWkCVbK43yzm
5te7Qfgo44k//vIqzwl3s4HmR4VSq0l7NirlSvlO7YC31ea4ykamjqemEKDZ
KSuIY/mK8y9SaK1iF4va5SDbBnmvhzNAarCXzkT1Y2+GBzxvvUwTzYkv2ILn
PZSPZjURP74bqCDjWeD4OTRaB0erh6vPoyAJW3Zc/cTAAbo6IGk7LSiaU35O
4OLB+DouzliKQxTe6D90v2lx2fZvzp0tRokxbb+c2ujxa82plJIGdg8hRl+m
j/W6O7vQ6BDEfwFO3/3tCxYDMp3wRsgDF8TmydfyyCpoT064IrXSmqzo29OC
455HtF0Aiq/lu3WS/nml3SYi4tqSZMP2DQ+yBLM41O1qUdsINATqZ6byqWED
ubheu2GATTZnV5lqV0oQTHdipn+sa/19hX5zJazINY76ggjFyO4FGo2DYM4k
iwZgcfDAD6bfbAptZIy+cxbc+HdfTj7d2UIbRVL/UzzTbvxkEMW27ti6A6SN
nuYm3HdBhcTDaGJWvAcTANLrVIHMIJ1NNXyUZpuiHiSRDCztgPob6iBLH0YG
vWOd984XagpaTZycrv8lxt/IWjWNPgzLTO0zWSsb9LjpJM9LjjRwvSLiDJUj
knMwtjK4tGCWM51r+Go5k+0fTJLcYxynaMPM6VBMZ+A0UxMgGI9BN1hOW8Vp
QGS29+p1+vHzif7d2OpZxa60TQQJcCyBNKzeS5J/kenH1QswaQyAnWBd3FOD
R6qldLLGGbpkYTnejgaBorIYLQUyE6n6uV3bCHltNU/JPJaO9cqZ5vuH10KZ
AaZxsDVK858mIkvMCakE7atzuDTMukLnzYx9iPWUvibJfiHU79CmlIWCKDa0
GUVaramPHffuRV2CEOyJffgsBKruTV+rCHdXpR514ZdpM0c981cirmVqh5Bd
o7R5swV7KdimQV1QI0+XoKfOPjbiJewEyQJ1NxEqsvp/UDRSupHc7LLE9JRr
AQHEHCCqSnToZ92lrYHQxoQVXdmijet0Nuxk+TW2zS+X+GK4bEVahVkbH5XR
u2bfi8LXrSFzxkZClaHmIRJyklzTMOwFHZGz2vw3q/mZvYdQb6bPs/gGiQLx
Di46UYjgCr1oPMxrnwHRSGT58kfGLcR1KRmQ+wxCHuZZSuLwwvIeyCoOyeBX
rpx+7CfCb9RrNRvsRUsN/0pIwZsPbFKYBjCctv+zFuMWgi1ZyZpEqqVmtXTK
HmNCNN1JY8CKMI1NfEadoh1JK1ZiKEPEwTLjLKodGI3n9/41NMEuhL/5H2s4
rnLOj9se8+bWq/ioVgPbjEFT/D+fwgPp2eUf2giOgmUTA5TtmLs7yA0HCgkh
TU8/5i6PmOGYppT70p4/ofIDKRVFjsAFTbNCY2R5Rgg7IaUX03V3w2EnW5CO
XWwRsVlcJyJt5MY94mqAFsUnh1KbBeohnHQylBNBuPfVl8KwO2vaWgp+mhcJ
rAUgM/zyxn8kBX0iYtIHtGzqNvNPB5Z8/GzZl8AZxCFJNbay9f+rk5Vk8CRE
tv2LL4tE3jT2XgoiAtaqr2GnyyF7zJhsRaKB92HpzhJPfLZb/FzyG60mJPf8
ge/6Iwi/6/GeEOUpnIBmSTyC8YNQFyfsAJJ5VBLWb/z9jlIzvj+kOc2uh5Zi
VHF+GRRhItEepO/8jxkZXnx4rNw3c0ac3iWpXelzhMHVr6rc3cT45HYzrl8t
C0R7iMX6SGT/DJXCMCqZGrfHNIfvhE+6gcYeh/XEbS+Y8JBHhERmo6skiQvG
3PeYkXW9nb1mMj4fjICfJY/ZO1alMbfdxI/BJJ1/8QfTLjQEMrhJpXSa98pV
4xiYqf1dnLzUojFBwRt3V24wHYAFlI6i3l+04/uzNpG+qaRFD7XfAGOCA7vF
vVyN7Q7OVINqoEZQyQ3iH+vF+F/sc/tx7nzVvYDfJHtSSTDGt19pvZGGeyAc
T85o/DZzgOS2OuDk5KSZCMo3VpL6oeFauDxfT/Jg2OMSdKZmu5kgPZOcWxZ6
R/ATxn/wWNim1qmtZxpOnn0/B1oxcuQx8x582r4PbrH37XUNAF2dCkO4lz+Q
kPYzKPx/P4Ii7PjhhYNZo0FDHazrA5RAMHEFbPog0tr+CHaLtcUJBaBv8muf
JOSN6tiVig+pJYv4Jomhg/tRpokX5fMWv76wnwF8ckkF+/18z3gbILko/81Q
7Jg0JaQM5Dc2bGOvaa0FbuE3MZAL2jcxh8yOP6mxaxIG0g11dRW/21oc57G2
8wyAIS1CRz1QtMTDdx8VcgU5m7Sw2VWCGWVl5WCF+AB2vwxZ57UNzLKyIDrZ
N8RrzF4YqQOI+MnO+amRjijZw5NDwi+kbzVpZW5gFzRJF0q4z8k1D4gSxpdT
d4KWx4k16glZODvRFcsiUo3qeJF3iGaKtVNykhZ9R1czXA7NzZVElZ+Fvg8F
6rOSuMiN9qWIHY4At5cVK8j9Hnbo492brQ5Q76v7t456guFoqBo2FANgVpyV
8MMX9DghXrn+8x2PWa5mlYRAxdHXbytgiFfbaal5Yuh/HkVbjsprIsXLxFZa
LqfXbLZkQRh72xzVlo0ddfhEwxXI15Y1ojzhkVM7GKH1IGe3l6DVVgi3SFbQ
psYreL6Tjom/LJCYawCHxD9ZM3NLNjMkRyynIZQyN9+Vb/xYiIzWmdzrnPk7
HfSaUkn3JYAY/x6tKpYeCzGkXZhBTJZkBntdCF50WDedFhILoY5SenT8sztt
zjJwdClSkSbTmIJErh1iWOyLU3eWGBb/srWItPSp2+/OF7B8kaJlqWQS8FWX
AoDufbPpcCevslrtez766JRhed9iZYdRa37l3aq1AMDF5oRlYoA6+cCfjL0i
xYgs8AiUcl9qDRohYIwOsDiCYTzZhpeHupqcR+PcthkaBSFJE4XUPyk+qntX
SnyszIV9N2znxZSisQf/MQRCrPxSl8aSLKz9ajO+68J1eL8g8DsHBnAuKdBo
gLX3C0u36q06ib5x4jBAJ5DSflsDmJDbDrJ3jMCa5ALiwtJskbQCLOoh3ykm
ssXWi3ndtTlx4HC11KsScuckfQ5nDqoN2SeBxKVx3QrTRoCDk3vA19tqwhse
vW4TQCzDetaGhNH/SOuLJ0riP0WiKrq9bfrtZBfhDgX25rcg/I+VU/40c0Ob
aJ57hbiAuRyJfsvZ01YAtoyy5ynaNVIzj5W60fzl4po8xIXkcX3p/7fPoqEW
SMpS8Jfb4TNh8ZDoQ6oOEgcJ/wgU4mgd4+ZREcRULnaF9LemWGVlLuspq9uo
Xp8d/YZzcTqq+2jJhrM/NYHwfXLn11R2u0XcNwXw2RBrSJFKxHz3trPkmxH8
Sa7XZ1RV2N/Pl7PHrn4/Irb1BH9iz1tCbwuLpx1GIOnaU8R0JIHjw6gOmXk2
k7KTHQfo8iJRgqP3mZqUU3muRlXW2OnS4jPGqp7Oek6XBDrJlit7cEqKg2xR
ptH0Zjf5j9l3azAFXZBGL0QND0SAKKQU0DGqVVTdEpXccY9IxH0NjK/qAKUN
PLHM0+493UUF6KnJwrk50JN27PyWhGPhF2P4di8w8teoVa/REsEhWfRAsW0G
9GEQM37iIspz9004OYSPxXr0tCt4Wxmtx5EXIzhVuxENzTbsXh63mdcDOFFH
ZwfljATcz0ni1p1CK1qvUhfKjk+qB47DN1aVL5EDt72Mz/IoNBkM7O73QZ4I
j/ZvpeGAqImnbPl+x1il+LOqiTmDD2Z4euTqa8ba0q//bApDWlem7NVtRDo4
6c63gl0pwCuOwUxj6+u9dfEffMvIqpjGkX+ObP/D/0JYcKPrH9XQ+g4vbh5w
o8mJ0+XOBk08XINIZLLkZ/uaYqXHt5HiPKAh6o6rpgLbWLk5tpGlzoOzBjAd
oeZNsh0ihDtuGcqY5KCjsWTnWXH1MkTazJY4GkHp4zMjjzJbl+YPexIRtrgK
4FLdIinAwZiy2LHkqLqvl/fd5Rxda7RQ14EGOvP7aYcRFTq3aqR0uB6yxAhO
wrxqsJVHm+wAVmds/445T9FUQPV9SvtkmaeLNB/VwbZOApDXFH7uL0sPcXMv
zE6NXuyhtqu8an+CaSEf5GH2loG/YLjjY2+kXNNhnLYgbfoU9Dnplk2C0fh7
opmjGri1nPINhdaSpdu81jCJZNNowKauEhrIxc6PDCI+3FW5nGy+WvVtB3iu
3Z35gvE3M0lHYLxVnUAaJyJTniAKuXAH9rSJZpzmMSMef1X6yx5pZIXSfGuS
osXXmNOva4poYkQJPurouLCwuJygiZfBQtHb9NyYAQuZ3T2VIZGcYYcXZEj8
WdaB3uZayXYAPwBJdIIkuvfdM5etLc+aU+jwnvt4HxBYXIfbNp0FgtaCG0HY
aBneXj0xoQpjiZeQj7woqWicE1kdlpCzxzMKlLo0P2yec968DmpfQ81SxA2n
u0veFRSx+Ijp0LuO+SCfwCJ5n8i3Kt2ekt+BrNXCL+QgZ2kgP9I5rUl01TlR
1kQWaeOs7NYmxdlekh9/Xbzvu/tDMOjw9uQLEuZRdyJk5zubnxw0z7qT4T5o
vXod1pjajnOJrTrzdodCGUghlos/OWOmTHvrsYHbg3M7XK8yRutW9gRZK33D
rbUhO4/OfPHqWVk77rYln2JNdy6rLfdmmsBrP9wi2S0ylcWdl9mP5GDPUIML
/9P+VPn/P+40XuRnV7Y6IwwHllEanhc2luZamY6oBpkYesfebRLY3Eokvg8F
8/4RHgW+5uclVkQKoyPINorhGGwVUi6rk4/hgoPWVDcn90ySDzyxnsrfVY+3
wKjWprLzHfwNTDVfeJpoUyn+aVz2Bs45qIVsFLDcrWSxnVSe0EWHIvUNQknn
XpDUMtGYbREWhnKHsKn4aZVY1tmKjy9vvUbdLWmmX0BblvaeMGFXTU1q7yzy
1c0g2xI5svsyeipxQ5UWGKDYUtWA7zRnclv5b2RDOdbEylCdNn6XVkNlzsyz
n5oTf9Kb1URoTjT5CaoGaEsBnX4glexKdF27OwkakpHYrSVYQddI0fzyvKP3
qf+54NaGaZ/KKOT7gAXkRuexyrxFGzzO9cKRbSjszu4eRJVOqcFVN6/kqnEa
4Nk+Eg89mVR3L47mr0xbINPobZXjd0JkyhvMscp1zMOc4/03yn1dIVdIKRPv
J2Ru5lP+RmNTZ1yWbcgHp3Y0X2oXY97TKnwy37Hy6IF/yUjvKjnRjOGvafiq
FEi3Dcj7w7z+MBobTaoTM9BmSJ6KJIhWC/daXM39JV2JySbfOpIj49D13L/K
TnVj6cz0BmjfWX1yaIkUxBaMczg75wSVszSptgM2Q6X5jtM3IQWOe4hFu+Hj
/sgBwJQr1rUTtF2wzU2QxJzvHbUlNtb+SZFffqRxFracdDl8hLFBHns6RXCf
/b1imz9SrhZOOUkFuko7sZArM0ohyXbTXm1kP/sOdanmATapT+5GsIjtbGPp
KpujBJH3HQLUl+hOteHnHJRXoZA5eYuo4M3rY2k5YZ1ypVVtAHr+oDYuoxSg
UyJBmw9snzHYsFFgaq4oDEInXjDbaooVgsRns1xpHCoctf+tGQICMzXXKa2C
yz7oIb0ZIqY/Ua4wtJIyn1SfI8tCaFltZUce5JX71ZQzx8nPF+OTwdkoAEf3
tWhxNKbqj/EXiuC6kWH7AfKP7jiJ/DEUuua0BfWm+wCAcqPfVnffHdy1bZR7
MISXNriAu/l6vrv2oxCb1L+ocFVJaoA3x+GMOs/gP12KmHD82XNhLg9ZPQX5
jqe2E71ARNTJDbCGlv8teqlTLUlpXzGcUeJBFtNuuyeag6MMFH79mwim/w94
iAko9ptwve8nGS0NLCOawrfT34EqzQzKRcspx3IMFiUxruMOisviFNk9EwOw
j9x7Pgs0eIh4l/gFkbz+6ebPCYzSWBGlMNk2YB9dfj6o40avb8m0Hponw56H
Wr2Yehl1Qw2mVpNnl1iREnGjszwVi3wkgvSWvRxMdWw0mWPkT0jzuECu9cS5
OERt7yzZYqFIBl7LkVweewDUAlVQ/RDCdlwdc2af1E/WUVb7qQ2ypzqscYIh
tg1xX0/Kcq6zk3URNulGQzJxIGW6rtLb4bn1cqhB5TSYduCAAALpWmM4y05p
WI7r57yOt1SZJzAiTjT8ltD1EVBEIk12PCcZKxwRbrH+zyyYRcyHqDUvpbca
lGMEWjNpjA5GVsMpqlwrKJjmGA3wmJKaExnR8oLb9AnTCWz63/RscjRvKQXT
kGXET+XQ94LlvmS0s6HmN0MdMA9XtIj5L7XnEsWO6F/yln89/IWK+aGvQzJz
Xcebh5Two/Mu/jSfWV4mCDEBkZqxF1Sf2eE+zwqgfgV3R+TedhdJ1r4f8AJW
Y42RA6yx60qyJMaH87VDAd1XJivDkzZ2V3JzixRpp4b5XtxyIdRqyBEWqA1J
zEc2hDgk7C/fL4bf3YGRHHetjqnV6YiAwgFnjZ0ymTjwOF8jiOFyuLGe88vB
SQPwC2HlTw83Yk66STp7iTqAHn1otbW7z5v03Tx42ZD9eWIXfT91qgGS14CQ
mc0rQvyyjOr2w1kUCJ19GQ0yjzvgkWbS2DyvAwoXVrzToO40PcdVxPlpk22s
uYfG2HHcn3pIWPbYjXx3etTfmpJL9skPt0qA8+jS0BRwHiFxtW/b5HjrxAph
hTyhsi7jlvjzvNMGFZYNg70MfJOGMR3cgfw7wCTRq+srcajM8pFeiTZuMF0x
yNViyQIy5pkZLuENTxlIL4W2LwFWiX3iOPRTgqsQc+riWxJKpyp9Muk2EhuY
72pKuHXTWNNv17tRFbtoiaXhO6Z1scsVgmdHXJos2ULgpR9qBcWqYWWWrSmC
0cO53JBiFwlSWmfr6B+rrlqe+TiH9iMgC0lWfV+7w/7ycZ1Naoi6C7euZFa4
I8DU3R7BEz3xfaO8a5v8nlM+9mUvAHviYQIoGsj7EFqUlWcVSel6I38kaLYI
3e/5B5H9muOglm+oCp60BHMENZvpYZ30bhxWWoTLdRGT4BOOOlDfgmfsytlP
l7xNvQCRv+2mQlgWtxuds5IDla9QiD0AGa7R8igt4A1Rax35M8viwHXjT11O
O1tF8wLqppS68B+Eel4Dp4JYUgoVHUYLsL4/CTZahhIp8HEf41ijuxp1ND30
DhE0gUwj4sV5zkvYdkjTyQvkp4yxy5Cwoqj2YPDUVA43ZNfp6iOEJ30FRjlV
kJwMlMuq95ndfMKBrjDUIIrKAHbh+iDQ1qiwIma8CPviGoOTEPCp4M2up39l
bvbSkDj0VvF6rwEBBBM6Swqmq/BYuosjxVJs4OZthf7CdFJ/gfDoyPAgeqep
ib427moE9s6O/S+3rJA51RvejTR9IeNhIetErPpQSB2NHI/7iHtSiHq73/DJ
Grw1YOMtzTEsjoiNIr6Iv2elF7LYnEp3MOq5SyX6H7E1ZAQYEq9kvAP1npGe
qau7d958Bkq/qqACWymq5hId+4M3tbJt6a/9v6xIolYN97AWazeV3uY+i84V
URMZ1Trogc940XJqt3w5d8GQEo1daeRNccqWA6/gsn01IiE9WT+v2zfqWSSD
PYTgPKwE1box1nqeQHeGbEkR9/dYBBnpRQqvg7Z7KiDV2bXWspBo9bSnwM3f
bGYVhoqA6g+ytCqoiL92CYAIWKWe4KNtBj5JSDNatNzqYo9/Yy4xCghtoWw4
juWVmzlew7+anSJs/2a4ODvr+KW5JPH46XWXNrjOhE0nLVauNBGueqTQi/37
8Zju04AODgxlG6RTmFCwqjqenw0GTUHjpj+O+ni4QGYnDRrSEghPU1dFtfLJ
dd3ChA2wGSvp9row2I1vfYeJ3TYw05OpH1Lf+HLRhU052qke1FOmns5oyaRy
HKVrT/YfiRLMCKP59lJI/zvWKllr14UCcZ73SggHNLCYJVTKmUbDx09Jcqln
4HcB2rxRkfoe79VE6YcQKYF1lOCCFBMRA2cMH5ehoobKQtGXt5muk9XzBCEe
bCBn7rE00/5dz73+9NTHVOXx/3V/tndbJULYwNMGb5hI+jxuKoVmCOX1xUsa
3/rYeU2u176I7TDxQmedEILJN5BJwCz8yEbzm/GGs5xc9Eu3RNQES7W1cTlr
i3eFY2Su7LSnzoVQwnS2lxAK/zz+pJ8EX6O+b1yaOL0WVMzdHji96S3oG3Fx
zp76WtCjjGCIzg3b42/dovi1Rspvo1NgfJmdN86wjXRArQQTwxx9UBRqu+mi
EyqdUt71nQZi+YVV/EOICUvdXFLlxphYXCJ6ya7EjXLJUrYnB7p7s/gSXqrs
MCLEXoNpEVvE910VJTD5RX1a9JQlxsAn5ATxKUrmziWHqj3q591ZTvDnH0hp
DO/lX4LLhvAKhs8K6q1n0KlaLF9+INOxtnFFAazUCK4LtqYuDxdRoszp9YvX
OoQHCyFNxLeQgBDQ8a6TeuMNKCkTqyhMr36rWpNznrqK3eAfhBbULd1bMhLc
5DFIsedosNzybcRMhZRc0J+0qDzKx+iKk4ngxD0Fpg49uHlUORvabQLqhSPL
Rkq8rya9SDlSMJ5CGz5ryu1Wf5l6i/veoachvNzB0pxYN8lRqH0EnNiwtjRI
FTW4/QEY8T+6Qj0UziZpF7pxHFJlJg598pnU6cWsoXh+QraLWUdq78e1L9hP
a7Oql73dZzQmVUhXI+RH11rZi47SXrFN2Zk6ENbhghkk7Ac5UiHaXfJxYHNr
onOpVMqE37cZ+kmBtRlnqGGLIsREmwMCBTG89o2t5hxrbNqmDP1bYXPygqMl
tqlvMNdpgvx9ft69t0bqsXVpToJ4wOCl1UT2KIB3sbNqlRVfrxhStCDoznkk
HpVhyGeIyktYD0YF11d8ZVhyWUQj8zEQ1tm4OdkCt5/3VE0sN57TSxZX0zAz
tHcgyzU9uHHiWwVc2oeHzlHKWN6Y6WRNPc8GggEqsCN6SQkDuF8c5XgdhgLp
xxDs5c5EznyWh9wYla1+3uKhP6gkjEC8SF9tqwr7bAIWS1xekOLBqN/EbnYo
QC2/dOLAZ/YQOsJMu+gz0+4/CCtiKnMjnCdd14Pvh7WLgXqwL+EYJz05AONT
2zJ4E4pZyHe2HvLKnaUqlWQ2dg+lGRUJeBWA7ZzoRWEpOwuKv2HWh2rhK9cG
5pqejjDdEtCbJPN6yWPfxK+/xisRHAb5/9dE9gKgkm3wJhBdfRyv+rc+fDp/
FBm93HvmF/40FFMBlDuw8uIX8OrU5o5lD55a4PH4z7N/fvvf1IujXMqbxtwh
5sl53baa90RcrvyeNgczYHpqXPzyRFSXL/2HLD70bZl/hcWokHcGfz7B2cz/
Su63rjMmcTn3saBWRsKmCouE06+Ju3p8D2IZyf7OqqBQrMHGUWaWVffVfcXn
/5YfjHO5gBPJ6LnN4exIgRVuEj8BjhBInoeinMaxy5cDz24hkH98OfK8wklK
OHGvDK20QI2voTp7lkPuS5l7azN5CPrGsW6OjqsVfhqZb8GVhP3K4VvBnsvI
WJI/pmzEsx3HASfyq7fSs5t6Gfu4aF2sdoO5X9jdgxic8fRhQKnV1FGZuaU1
6qZDRoPHsdtNuFcFUJuUCGblQhrwkku7UinpPpp54/NPucUsIrS09k2scNMg
ayKIlOzJRxDk9rJFDRcRM2wbfcUKjGSiVAhMZl998EqtgFmguhOrLoH/Ns2B
FreiNJ0SPe//9deEaA23SffnnQH7e0DDy/DKTK3K8G3s5QPmYdtWkCnWPdQ3
MRTR9ymkZ9xAqVtHyTh4m6NBpiljEdKwv/XNiMH39K8Sq3fcjI/slZjZazCi
ERb0wqwU8fiXTP77lYJP9s4e7e/obZkYEcj4zVnIYVPCsbCPYI4YobwOeQKx
r1JLl42TTJqV2DMO/5xhQ3y8O32S9U+o3hdoXubZbwHe6l9H/j9V5mMinXvV
GgCJOLSta53ZWRQVhMEJGMJvZ1YmKjpEEV9YnEul+yga8dTZWqTOCULvTkYR
O5kBEaSUs8RuXvTiW1MJ6fJ+Idj7hlFs/3lLuXXmh+/vrqRT/4rc+HuY21/M
ue2CTtfNF9jCy4o2hIPWY5ehjfvFvOKbRkjhqmOHcxz0hwZbK2PziL9af5cM
Oub0aTDSn1skSFBHpZA/b7Pu99X2lRFrNEsoEB4G30asGQAROsU3/gLiJah5
s1cmpBDR+ggm66jyg2vAuD3+gMD6FPC/Pkw8VaS+n92EVFyH0jSH2fz6k1tI
HqsmDVYxwBpkTfeVPShERxiSFNtd49IfUudZjowHoloanIFDepXh9Qh55e76
lVcmrPgBwcHn8KX0A/jwoT06aPScDAU17SpEKPqmZQ6+MGh/qw0xP5tHO4Jr
TVAS5+50Hgy3bCp3XTYznDUSYaWbOTyXGe7yTkwApdBZHD1GHeJNdrJscSYF
U8HXrClGQSivi8Kk8IzZ63jRlpILYuZApgIy++tGJl0V+wzT3dHJJ9bDg3Th
RRoGhTpo3RELoDf2AYg0z2DuBCiET4ke8Vk4g7aHDzJX3IAgso3TU+HSXU2L
wUkJfHBV53mra58OvDteZ7GjLBq3lV5gWG1kY3aXBODhfCIas9gZViTGnJvn
AoBbY7uVB0Dk8UE/5uaJWe/YaKqsDccV6xl/9p9yQmUwVnx2zX4sjQ94m/mf
BtMcMrETzhMRmWONVyXgzdTKwvD6wVBSGPMc+PiLJ8RS44va6vumMbmRjsYA
F2KUdUuSNE4//neNhxZc3FTkMCXua72iQS7JY2lREHY1R+9ouds6nHyauQct
Cy2Q6BkuqfbWOy4fMgJFgQG7OQl6xQCvIIhiGJy/dZ1djkbHTlY5ckjwUQnY
QkcETxjErBbcGLDJes/TAvHZ7xVZFWMDww+bywDV7zmUvQDVW9RbTAW0wwZM
UXOqLFrHv2NWq8wZBN2ikd6mBAZNAYjOIBF7U8l2FsUJurpzh64Vi9kkcoVv
kPQQxWcBkQA9d+8K9CMmiyFN5ql3kXPEmpLaG2ywBT3KAw/IPtT2DiWJc1Xv
mhSmLKXibrQtdad+l3wRz5QGh8rR+inxqOaEJ5vVUALxO6niGG0rc/Q0//8E
PbDwsL2IO0nVU6M+U67Ei9x75y00NH/WCh/MiFLwcdz8T3D+iR0UR6SA+DKC
uP4lBr9GzPkwPMHmVJKwUzvzmNLBgtIsBHdY3Z6qXscrngK4+ZlGUHSx561t
XbSaTLlXMfMAbtkdHOaK5g8PfEvkEWmo1ckhquZ35asVmXau7lnpo2LK2yBu
JfQgjZanPHQdumvFk9OhqNi9jrwFdv0htWAdO0k5zClJVvXe0wPhaaQMGXgp
0A/x4iGytn1b6WUPyuimJHmeJyvYfqZPI1tMErDLCM9zrB8v/0+ZTDHjjF5O
+VGiP6u4glr1RuNscbt9mjj7DIFP2hI4dFMBAYv4SP6UMmi/U2SuVVhLtHuF
c02xZuRze7WbK5iYB8zK0e39ehx4I/TJh0MeMmddOcB3TbX91zOM3mSud0Xa
ltdOqTOxjpO4ygXN3IVnW7OKhpDwlD//lzBFDZi4udB0xIL9bRE27heceVfl
2ndsPLGzTjewNVUeLg168DKw6QvqV2oJJjinkcMf3yTjnIrDX6p3b83jXATD
LnXk6aqM+0mzm3mF2EsjxIdJiCf/GwgMh7R4uKYBac0b+em0GIsvmY7kfRAq
0vRWbAhtDfF2Ch+k0F9BeDAGKKd6BhuJZcdI

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1JkOZ6oxskGfwquvaBBGfd6xzGxUNfA8T4HyCEOQPKKCWljvkCkmcXo2Cz4hiXy9RtNA1QzSDgcXX0H0+GlDjkFr2LAz4dCy5d/KPo2HIkffjpC7AEKi0Xnf/cFRNHSf3lRm4j490XpYH10g+XTeyvsMgeS7+uHHDG4y/i0MFYivh8OJVnA6Hs9dkGrJw51zOcRoF/3E01ws0DQBw3B92vusUivsXEvRWE+Em4XjfVUj9ZXpTcsbw0PN3LOK4PxUalm6t2YV6QRJEtbXvgyb2mR1617XQcUjgz4XIgCTJ9HF9KglvDqO+smlQzMxsZrjnLmJmSDKHYw/C+gdnk57H3MJnJdzSDCtOR9eRl+cE19nrsHY0Fo5OEbTKNappbiYO+VRful3RNql8JpaKXonPaG00xS8BwU8rCPqKQfaJA0C3HVsdzYq+dOBout16nIWVcLO3auU7cFO05bV3AIU9UORp293r0+joGcT6ictKgJYFUA9jxI5aZJx+xDmop4pwqhCDcaSqULR1XJrpeuXBXY0Fze+B1hkXU38W349heqwlD6o+HBtdKUK2+k962eD9I44SFrotti/6uDdCVIWWX1GygsMmAfNObhGXuLlG9yD8FNYyA9kQ/x+/lva10Zh+6cn+doaDSlSh+sVL2fxIXl+QfO/ZiNE7concPEOP0jlSG7Q/SjE3aB/yhVG8VdQDfcqv5pLnzd3QaqhkqT7YJr3JfnJIfYm+XX0MZSsVdntHv37Hsp1M2WqtZ7VcCxM74rCp9PkyhHLwK1wlozEzyD"
`endif