// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fJzVYbjQ2WIDc9WZWJIMijZ9exLKNPLAhB67uEJY8zEpaqtra/MGBl+GJsOa
P4z8ABbEBI8QamG/Ni/M5mRFv0GUksTloezA46gOWb7pTKYZHFKiD7CfT/O1
2Qnwu6jPKZv13mdq3ZgsNcNX8NAjY2F3ErBZFpNNObIsRFmpvLHAl5Rqhd57
nYTdrvSWDnA7H3Ki3oZfxkVB+3/EVYRfTBObOPCF5yDqjdkVPuGBxDFWZT5c
6BC+bffBTKPSEv/MWF35i8wRMkESJSzOpMLscNWunS5nZ+txlo/BbHThXZDd
3Ud7o0mjmu7pL+Cywnyq0YXQpEt0DDSmuMBv5GNCmA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OmmaGUxqrwUBoF5TPCXgyeNjsYx0dI4LlV1EcuGWm1jSEyUgUk3iayoiMHRr
+AzKKGnH0hBMs1JCp+8TLvVPPj5D9CLuQL2Vt1ljQTJdl2D7zgiv4tGnbyGe
da7z3+Gb5RqDH5wogROOH9qmi1sj1EVxV2EvJbTrlUsY3QPUfWvlXY5xKlwW
HR4xjL5rry1HxL/ipCO2twt9JNHGT6vTXTBzzYELpuJ7G+2v9f3Q9BmNOcC4
LGVx8fw5FFOmuy/uTfTZmeVxH39XH12BQZ8xTJrwjwJwco/gPkTrsKTGb+ge
GorYi+EA0tytzqdHmm7+gqBa9Vsj/JKgOu56sOn34Q==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
D5btDernB4U8D56ySVTQTQmTod9ZhONLsT0UNedQL8+pxJVM146OMsYJ4g4B
c+Eo3doOFQ53IFht0QAY4H9lPYHe2fE9fpmVqLhoX7IKmqEPoZ60D2AWJrs2
73amCCYfHurplLHfD9OugNd2V8DdaDIaGgUyirQZOKtbquo1QgGfE8jY9rH6
0qBK7mu9trC24x8TRdj6vKgdQkIUY8ybAkPXSrQLWkebzRHsRmslLegLJk7t
S6D0uw/d0tnK0bVMCdgghi6W5KYinAk2ro/TgkMwwvXTCHPMIF8kqpQR8UvX
YFZ4FR3B+wq+rTXnV7PwmxSQAl8/NR5k8OV5e6XZVg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
coGGD4EILuGVlMiEF74coYzCzeFSSc0aPdfRKuV3/FIwLGvKTniPJ0kpfIun
JcsxaeEtpJOEEv4iz5RQbnDRK1Z3WgF6sHT9L7CPgL2PBFa1wHXl6PthIPtC
Jacpp+HwRNm7VamZQB+Bi+1CB1E951gWHCx6H21kBIFx7PCsLt7bIC3aOq17
rHxNMfZGBtDdqmTXca/qkaFIP84cWzjuPfSvtPu+8C07xxvZ2w5IbijRBu2q
Eh1KSs6yqbtlw7dSjjjVTtbDvSg2P3eplWM2Oig1QkFR1+YHlZZgCDygiVe7
RM67L4lVYDqy2B8BOj8mD1mG7j3yIBMXM0V7+WFsXg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BEOSV0XFQtlNfpX4cN1wEVjLxnMxCDcruZmdjjXi3BpTC36ucvfaSMV5Btaj
0zvsFlBvGKdjD2FIVRWhoqz/RFiDfJ2pRAdG0/ahsyAWkO2d5bV2236L1KWG
2WQiInfE69wd9SQnKUCxIePaJoezidOh9EncXd/M1Y6b4I3IpZ0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
hLx/T3UW6IyywKyYtJs7w3CwLbMziu5mjEGd4LRaga+ACZb3zsMjoTvQNPts
NRXI+4BtU047rloXHXHJm4rcL1EIZYtIDMdjHQKHjWvwwo6bXK4VnKgmYa0P
Ylp+6lUdlJv1B22dIzG9iq+YB3KldXSgua7CQFVG6CJLDBFG6LURZj+EZeQ+
jyuIurhRw/7+19WyDD8tXRbo68t66C4duLOqBupdj8fkXKWHTYcPIB6lyVQG
A5ids8bVftWlXazsQ+6iQK5O6B4zVCOYY6SbbAobxYAcyx4z5WPazSdh5gQW
QyoFdC8Hk8bACofptN8rr4j2SjqRDkC/wPEc+xNy0XBIeLTDsgvOu5X44qsB
nNieZNnUeFPKIZwzVnZqtCOsTo6tmfsxhziooz+OSiJhxYvkvpY//14YGdFY
X/T6B6hYGPSmTmN1l7xfEV4GGABlrI2BymUvlU5DFmp7ZSonJOyhtbmNEmQs
tOQg70jQjHAA2CxkAgevuehbAVbKSuUE


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ij1elRgsy4bU25/SQ1dyXGyBZ4rN25FpsdSKrtk/jaL2vIBxPbtFweiRBOpv
ixO0JLVJO4l43oRiMTf5kgGQJqocYu8il9FrKrE9AmZe60ygJ10P18NuSlv8
14bP0VUMDZCVchFdtb6/AL1rkSlb2vkWGonNxsy0kizDVXarxZc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
r81w9ShPsBqKHHrd+FozBjZK/+rW7gYQ8nmpOO6nNgmlOJFW5KsxQBteDdpZ
irkO+HVHptNnznAZeWdUt+McyrbfYXNGq5S6WxwCfTKenPYPhHn9THOVDuHP
mhHq1IA7fQptM4qHYPfSpkCANdAYRdhA0ApK0zzrjjnagkp3I78=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 666304)
`pragma protect data_block
0Fe8fL5Ib8X/7e0sj6juClWmw62fobRhRL33ZXoOlFB3pBurIKg5F9SeBsEl
eDOWsxurIwpBiaTawN5YAQ5YehxVIfIZyGUzf69GobIKtEwdXcMNpDW3NvIw
4Wbf4kwgeZba7exSXbvVHK8ewouUwemm4j5RLie8oT3pOMkyPVnzx8Xp1EC4
e3EHfjcbD1IXpCulHw0IxzGGl8I6mvGxTdKxoTwbrNLYel8k1dIvKSteZj2B
9lKni1eZN0ax55Cq+kLI1MkSzYuLfLQPuseg5Zbu7bMMhJ2xY3BpeKE6b0/I
abetyOP7zpP6ROs09HYWjcP5czl3/ne0i0NbTXXme1vA3LgK5HQUfglLQrwX
3kdhZOn9JAAuhKA4HC0eWbOwjiqhtYpDRBZbrYp+l39SjLlxCKSweMxnPZvo
m/lgGGfQMUKaAkzjqmQbihS2wny2xvBfWx0mTpdsin4mKwJ6VHYoEihhdxkE
9Bda9e3HPBz10X8L+odEDJNpdX4RNerVspMmTdrxzZ2+olPxbaIghfjt9gZX
o9ZlBTF9NyktGCLu2OfL8OPw4fFPQPMlFX1LDALZ2Hjxp5i1B8vFCs7Lb9rk
4sjr0/kd4pHGaSa13IzW4GygLuaDwCozYqhIyWroG+PIKhsv+c1uhwyp3DBl
vMkuwQwtv75QjLpGMIK/q8uqtxjwxbdw7SBjbusVOoM2E6zMR0pJXnDsmv5g
3jkUyWtP9bqfW/sx8M0QmTT3xmX/bHPqZIqaQGAnLe7u52HkOOeP2g/z4ZFC
RxfthDOCY94cYDO5j3yUdzNYE7zfenYl3815lriMnu2z5qZ6Pc+zPF66/Bw0
wlwIASf5VM8E5ioMdWsCIuySSEBSq/gF+lQs0Q2r1g+biaHRTWwPoqXltADE
fiRaTl4W+qFIPSRO+ZeSzJnldqf2mw9owBwVm8YRkC8rl6c52Rir9jSBJ9RD
7CWs/8Awzr6bJCTlm6W6FhxRSY28g1U8BgrFNHef+GrT2cjj+QnATrCJ1PFg
LTIn3GuF7CtL5En6vWFe4FCRj8vHSrOAO3WC9pF4La5ncSwkov0B0DIO97B3
yjSjak105BmuSHCqMyYNlK/gw8xTRdh/56Y7XPyKzXrUXh8CQagggVUxQqVv
0z1pyLH/cjaEXltAfJRgpwyzhDFwiI5GTLEWmt7LFvNgcTdJuecI+AZO+cwO
rN88bv5S9CxPnl0iskO4PK/ww4KzZBgJHaGGK2Xf9mbyjNs1KPNtd9xKEoRp
Wss36Tos8SNY/vh3zHjydylHHwFLzzYAMcNgO8oD/uuN14A/KCb1HAhJzULj
DUya7cq6iFsLUCHmlHcTMEKaE75sl8zJmLGY4UrDSMeN7TOo84y3rHZeYi5d
eLN/FKM45D0r3PgaiR1it1i45JkO+ONLJZzsqSqQJdjkF7JY33VAtLRMwZI6
yFTS3eDlnRnPvFiT5YyM59tC6hrVxBFO+5bpMUJf9J5DRGKHweCKuVzx2ZN4
K0bwiHEHtvLCE5nbU3Q85NOIxNWmDvFa3PvqWKoF9kQQy/yE3CyEgBzmLDWZ
tyf4vo7bgWiWYaC0YXmpN6Lm2aYYGzvEPn589tKmmwNB8+QDpSPL/qVzmXXV
GjLUnM7bzxkKNOovYneNHoP74HxVr8CgYzUy7u8+ZtEb14FiQuqf+MHEEIEM
vioPjPhVt1Jlp/vnLzSv7z3e8LTrenCENKLO68jA618Fbs1yM40QH1Ehj/ea
Nb6gmbuVORNStvSRU5HfBfH7jENW570BTmAA1MGTrcempSUvRKAwHGJVocZg
SRbIiGhaUT0oZWtNqwE2rO5U2eKBqk5XKS5kf9qgkVE/wboKMEai5xAHGRzG
w8h3UuVyXOnOHySC8dEIe5aXqXkCWei1YztQahKKHVF1o58Ls01dTGki9oGm
M96VYYsl/CvZPrx7Qm/HDIrUGhWTKTkJp7lB01rlqec9BLZPG5x1Tt6uX5qM
85XiZoDMgHeFGuBTY3muHugGRw4pRvbT8A8N8OUPQAStfgiOcngPQtfiLuuI
2sYtMzDlZ7OvhST/wmoJWOgtdUuorLm+2fJE2w6Lz9wVcHe+fpEc/QG3qkhe
cMK8dBRgKhC16WUygnXHclInihpbYsPl27aEVP5UkvUYE/baCSiDc0jDFQZd
e46d5yVNqIkRYcW8+5aJDE4LXc55Eay52g5dt+FCbQqbd9ttxrmFVQsFNYAc
ehoGi4eQpjirOexsRthEP429fvKRC5Xzr5T4d2nb3lUKViMdoEgvfVQFBqtw
/OwmK2pMTfykDDiWbqZ7jDr+EhfPq1E1aWbmZfEzpvQ0LWX7Fz3IsgB9or13
MCVfSQfHez217X24FRaHuPVNMRqRkcciBLr2uiMbWpSZWiN2bCLmjwYnE64C
5uOaArRBKEiuzZqQ3bpDrjdnWDl8XW4avwV5W3PTWn38oHWMmS63bkTi96gY
ODuNnOCQYn+twXVqN7pEJQTJW+0S4cHVlG4s7alyEH6JOkfZNsGVt2WB2N5j
7nWQ8AWcRFNhcUbdUO3Y1mJbn2ZA5zJIXj9Py8FLkKThPW7gnnBm6kAocOBL
LYYT6OxHsEOnwjNocfzJQ/wBBwEhJ6UcsneopOvMKcAzxO+PEEGmCQE0uWAt
ejtef2VbjC86JtfGhs9da5GcCJR+BnOiIcovEpRq7hyDHt2GgutRZ6MfqCEQ
yYXBMJ4tRvKLNYQZwMEAAR6VokH8I8WXefJRSnZ0ffOW3lC+CTeTGp6NEIMM
h4qxMNTJ6Ow3XHkky74F7E8NkmjBn6ukWfWuvPt/pEK0Za+BI6yfqcI9+SJb
j5ku+FBtXr4JV/qNT4SabDyeUrDGbc3grtZLOvcQBcsIn19GL2VAxXcVlm2o
Dp8d+X7GEmIcxUxfZBb9Z6MV9hXbXQABYkRHUpo1yqStofhrV5QwuxiuoUqM
0bHDPD1JXrqrjWBhQVW+ulIriNpVEtzW4me1TGMr2Qk4JDQMu0F7arHe4Rqd
hZj1HkZkUjWjpbVPZ40SQEkVwjHMglydTQBjRtrvfxCHy34L9hLLKaXAshza
+p5QQb8CjUc3MQYE9KOHyoutZ3b/pGLz8N7B/vZZUQi18Pi/DCqAyC3eA9os
Qg2jBj5J0CWDRT3XX9Q3VWjI41oWvSmICEvIxB64A+3m/JRrYvCmTXfBdkbF
Eng86E+mC/sb2fvmRpULWCnoIZHbsUPfth/lCWLE1Q5dlA811Y70WQkdbnWw
kgMA08i4b0hYSNulT34xTbT6nCh+3EhX4WL7OTP+vuz9rOHFTB473TLq/2F6
rkYfWlHcNWXiyMj+rKOjcS7B8nJhKXv93zTDylp1orcbTCmua7p0C6CiZML0
TekFr1wWH7uzY+eM9SUI7bz10xDGVIbAlcPC0tqqjec3TZTm1HvkgqsuoK9p
V7o/x1XdSUTQBSzGhxfEBdw23Z0flVT00KDww7ZMIFIH9/0mXUgQlsC5qq5a
PtM/nzl2nVJldVZsQKpzxcz7eNyuXToIo28T6scpakqU3n64acCmg0DT4muX
vQheM9s13G8tvbF+DAViAC6DNWDKCg50FuUXeVbk9Mg8Cqe6bbN/r/iBi30F
1nA1s54umS92EJU7eVwDIO1GDPfDk2SQZWT2qCEUEjQa0Z1C1rcgZNNah/Tk
zqhGxXozA2ED93fsnhgx3eWAdi2YhtRWyH/KY37YMQUF7WXKtKlij50WMesV
+XkgLmaFW2utgzLexIgGDyuURjpXHl6lLU111NuS7PAGs5H4ql+I+V6MSDTe
ag2gaoRVTo/SBWAEkP1hSniCB7ITw9fterWf6apnxIzFYDk2wC35T4fa2J3k
KYrcYc9BUkTdyaoQ+oT5J3xLVegykpPsDviBL+igGJq5uwTIMvPCSxR4HurR
hJPgd2+hJey22ZLQh+7P31rwDbY90rEvHf+fgTD2QLWoOgy/7Nhwm55XjI4n
2gLyYrnS0fviEqgTf+qUm2h2QPwAvXGDQVSZhOiQpSrUubg19w55FDRbt/IS
CRDOsFcOmaEyiF5GNjysyqh0zg+vXOfemOZcuALuDhGs765ThrBvnUSr3xPl
sFwV7kjE/g/BBjS3htqykagirbJmjj4gwITTX1om/aUkyHC2e2IfFHngW+WQ
wvih0/p3cKkGSZODT/4KsoTGFJNeD0FffjY94Mam+N9NdeN51xmZIMILgZfd
f9xBSIrNi/JjoX+TuN8upK2ElzddIZzAUrzN7kr4EB49pLSETHRC+KhGe9SH
TNq3qCR+CNosoR3upKgm4FzBBk22X19Y0eLtbOFmANX+4/D45ENyfLbdL1R0
tPp6gQbZgNjgDBZiv8ooYrz0LyV6FcHYrBlEl8MF3mD9FsgmZfARuvfKEH4/
1o5TNvLZCNTEleds6jTCJxd2GMksIW3ed82bIiBjQhoX/uOOCf54bTTyRduz
RdQQbid0U2px3U/j54300xcSC2xCD+hak1Duo5X+MNbwpvnyXBiRQ0UbhFxH
EqD7HhKGzfOiJ8APNT65qbpx1Ctfvlkq2370rJhSRPNcGG6q84pNKUuW51ab
4GdRz5Odkcstxo//mRlJJayg7i8q1RFkaidPg5CtImfqsf6aDAVCTUg2KjHo
DiFf/EWIGDvCuPDzmY17XJ8mRm7q646yeEcquXv9XhR1sex9P8R6odurhpk9
JfrPzMdc8QhcQ6vUrKSvXMdSbyrLDOnHGjcJrkcUqYriL3ZROOPEIEVrakKr
SuCwoOu7c5RJN9A1fjJyKoyUoX+wfmoWip4N9muTM9pv0KqNDbYo0rbGUKMU
fpZcPvlvpYKaotl9cbvhe1hHHuRk+ztKqc+YYeRfv7X6V/EDrLkEJaMrGiGu
Fzmltbuq4Y6FWfuxlg3zqqGgOSX58esvgKK7eKbWlejEioTSoc8NWs/CpN8E
8QYk06ZH9IEmSFXReC8wxAIpAhJJJN30bVy5Cn2Gl90+oBxwxmM+K4pii/qv
e7qQPksOH4KAbwE+I+tbBitiiJOP/QY8lbfPXJrdDFFxc+7vp7SH6wwOZSko
zy98v4M+dfJ+sMoLzN5K75HNdfGjCwXz9x4VdqD1YDLf8as25zHdH0ufKjkx
e7J9YI43kYuhDtcrqMF27QMLv6qtdse4lm5Tk3FDG1hL21T4QSfmRJmQ9ZAY
YMOzxuWU/PA4dexGNHnvbPqn6QfMv+hSPb5PxVtXWUZjGbOR19d6zKnaS+4o
JON6crUTihQbfIayJ3kQihKE7VHe6/NoTfsgSHvnq8H7WZRH0aT1AP7PtrnA
08C+qrLj1kOffzzQzyp5B8iWtlOO3+/ZtFCf4hYNYr/eAFihv2/Z8v64H8Ww
XznqRb40R+OEGiCUyIpMX9pT8nVmCLBcTtX7n4rIqcrTzuaxX0XBhRVRZgYm
QbIZpfLWGnRy01tIdgtUXuzu54zmgXZZulAq8E66Y9bxL4oLBPaDjFyrYihC
2c5zwJg/ZNwLe2iWyXIafjnqAd1C6noUvqKbTO5VARxYzNlo9fCd0tc8cakq
qNBQFI0Zo9wrf7nRtovZo82UEifKQwovG2A/PPhsuPjzrJKqnVC3a+eP5LQ4
QRT/TvpJ/ZQtKK6dOPM/aG6aPJ4w2s8xMjZkNtkuIcdOrwUMCb+MAWA0ueD7
sK27YG4wc4GkeiX9xDQvnZ2f/QvJcvjbIJj3ZFEfsC0yhDJVywXIfmbpulX7
vixVP89tmtCv2HETS2i1PEVjaqqGcpVJnRpiMpss7z4EfXwjQA6nW/wKFfFs
Q8IJSF/t8q/QrHDCAtxC6o3nOLH9uqTKfa2vfxwy4n4f1+rm1kSEtb3/+DTA
GYs6B2Eby/YSLtBZh/o4Hxbzn85p6hm0Z3kZ9jT2h5+J+z9A8clDPEPkWT2X
HuODixzuCHtqlYOLStXOUjXNtxGMZQmOa0dC7abmJshUY0hg701o2pIPh2pX
a+Ew6H+dIEkFjz6GUi0lWr7d4FHCYNi4BoO35MnXDykIVcVZlmcZyXb44YJH
U4k4/d7EUWZKs4piq3o9C6IMkQoKOMR1rSkKOMTjfwQvXEkAzNk6YgIJVjZs
gRa+AKFKJWIGZIgsTDyeTPVDknJxW9qAoahxZ9YvV66rWpnHI9o9OYIHRuJ/
GGNFbmiw1y2YNtxRR8qGaah9OMoEGLC1/CUnNOrwjtAe1LmCHIcXdS0DS8Xk
7YimVr+rQuLLt8/WQ8xSh9Cdq9HNp8qUPdD9HerOGsTz3Ib52C8BrY9R/bzg
4igKihMHBdabIqmqEoe216tFIGnE4TB5hNYPjHPPfoLWnPWvppIIpoHDBa7l
7Wu6PkiuZTSTwrJoMPskwVMu7TRAB8RhnBISKfQkmybG0a0HUBwYmpOkHi10
ZeN+rZHjb9afx1E5QhgCQTfoVenLGDmEl0Z0TiXrzTvtmr/L9TdtOFA+jP5z
awRGg78skbak2sbT0MveQr1x2JK029DTJRD1UfyKBfvf+/lWajiwbl/eWqXA
uQrY0ZllNxxtKJM+IDzB4ylR0gGEHhIiXLE4S4kB3hmaNhxxaC/nyOqQBHI3
qCV6F5vCHn5abr3/2cvfSvxVSujSm8uNKb9YsRi9+Apa4Zjw5r+G9CKJa1Q5
V96rsXpbim/VIg6sIY/AnZHkmOLYPM8DAUA2PJRoPLut+ZIrLcyqmV8fGfpn
UiAVV10wkytR5lZErMl5BOD32CEPdAXgR8xY5SIkyedd/KsWSx7Fshko/rap
iIP7N7pD+RvKWHftVUA6S2tJA+D85OnfQO7yzzEGtcc6enUs/Cfk9in+6Tev
ZogKE9bm2xPhlCvKwcd+0JT3V4GaGKWZJ+jxm26A88AdU58bTXy1/YjLMjxR
GTc1wOep6mLfmdTEcauD06B6nnjxZUfF66RjjDH0eHyNM4mZaL/LwIDqNbqo
+oQJFiPb8sdwjU4zkQ92yJh7WgqnxsvjfHYAMUIcE8VDQ3B8/03eLiiMUQnH
1hgLEatjPZ0APWM7MnVo4QLvRQmf/yXe7qZJFv+T1NDurab6tH5kuCU01Z28
B++mo/CzvjYqNkX018A0OtqXHAAlik/KC83v+NUQzgERa/a55Ug5r7pcu2B/
47LrKRQIB60NNRW0L6+jW9W9JSKNWUszZ+sZtyNWpSSGY3HmbJ6GKhNfagUC
PUY6UK6SSCQQT8nW+rs+54gRPjLu7v0yxXZo3nbCydP0gmqzmPar1mHetD/a
dyIVQ7lvCYVF6v8hrWyE61ln0bL9saaeBWSo7/8eGQXcW9KSxQO7xH4mAYKz
LgPcAyTY0aCFTd3sj0gJflnf7JItjFhHiYut7Q1Gm01lq1q7j5fDZYfyvAbx
4WJJZzBjl5K2+NiyHTmzyD1WO46X2R6gFQlxrtQq7HJvxp23/cjjCHvmkI0C
VV1OoJGpN0Pk8hTX8PoTkJr0S8HU8uV6mc1hie6tlP44SSOOxUCSGdwkuIic
UeQqV9KHrjtdj9SuMxdFqpy8JiqZSwTU7v48y80bD3XShF5lyYhXeGJzFsWD
i1i/pAyAQC/qUUXZm02rypxSwely6Rp3Np2IkRCKtw6CCbzx8LjvjiMI9OTp
UxtIDy2pGIs4QneOgOkXx+kuwXTC19p4VM7KjuK7liRFxoWQPLAtzBLXYbde
1s6HrGPy5B2HbDaiUcdfUnjGzcHGO/1mvePjaze9S3gaYz3dNe78NKJ5myKL
f6hx7SqgvGu7plHmLsZGcuieY2m/JQ0zpoupSGovbgD4KTCjcusuJz8vJJTD
rMzvBkFBdvi6wxDj7CLiDYXYh6D1MdZBv7muKlHYu2F+NFjMEJvNbFmNUA/c
zlRIVR3Yt2RhBXibGhmv64o/JggZo4YLYg8u/X4NfDMuWDwfbkprIlTiD9Dp
vkOfrX4vRgn3WtwoLaXxiyvBcYXVnvOy9aNFlg5ULk4zWKjTyMB22yduJHTR
jm4g8tCsWRyLHk56mCin9FbvXts+0st0vJIAL2oUrYz5Fkz8SOq3WHYJW1yV
T+quYXrSaJjge2dcD+9/ojUi/YE8qU9Xwk/Eca8SWj20D6N0rICtHOFkus11
9KfSEXAAtJH3aAW30f044zZPT+WS8ZqMBaQGQT6O4C1hF9JSOgdhHsSzFRIg
ebqn5mZruGjyzlPFWkYnekdXF0e8Fcdo/IOuHRE+IqFUzmJNpi8MSHpTHwws
iBorJwYTn24/g8LUPVsLihrY+BCC8LaIBJziDCVGJRS0WYbGWVjmsMLUjXV8
G15AtmkA07A4YXeBUlmDy0HNVEY0ssa911lWoQjTjI3gtycHm1H2T0HKQMg/
kt7KXnSGG0JFd7NTYa3ZxwApvEaeTs636hsoxlya8eS88AUnwTOVQ9gwS9Cg
P/8dHnnDW6/YLn9tZEWNcq+GK5lc54Hx+hhzLbiw/23fLtTykNj/pNxm0Jxb
x4waE2SZRYGLh+AQ1l8AywoaNqAKkXMh7gVDDqvCY9p2pZyEdYlKDBN/EcBq
w9xkJP37++ts6XU/CBW6zXCo1cyZr6/hYg/D6LYG2c0p0eBZHPGccY/FQToJ
I4LRo+7jK5LJGtW9qunWfUMhAS+AQVz2LxQqkNCFqj0lk/vWiK5db/aGH/iR
YSvpJeS6KLRM5+HgzZ9cOibv8WjwwGBWQjt47kHClQHPXjVjyrvml1yAmf9w
4TnRmo+bLF7j3cHCj4X/qrnJC8HrbR9E1deDziGS3439tgCSLUD0Mk8JPWhS
DMt1QIrEMpFoqFx1Gps6xtFSLpBAcxVZP+/XteWRfshNqFyBzg4/XHsckImG
cMZ2Z1joEimxzLOeLsiWbcfxM2YBDHGodIfdNskLnsNbLjRTQ52kdwEY3nOJ
PlEK2qFkGVqmzcuAUXN14u8dQPkM750Bw6bLYsX1y5lOjX2LM74kCzAQa3bT
bRrQZxj4DFhK0cGEre+x3z3ztiO6JDXted04bpBQDi4JeZlsJxH8Qu/of93Y
Iqmp2Vc/lKawfg89uFeWJWCi5qR6namwf+GWGpH5C/kwBNhaJVyTDWOlsDnj
kBv/9YbHVpKuLfSErkMGd2fJi0GeHsO2mEu7jUxsUCACjln/uqonJX0UOi83
8Or3I28hFm9m3sDaL0RQuRH7drm3lcbXTCXWNsovtt+O1HlVkbnz+gcWv/nk
DPHYInmmwFo2eXlwm3pU1LO8Wbcx8phN7Rpd4+QJsu+dA+nD4ThhDO18DmeS
82cWdnNLH7nM6x6Sw23cmIa9LqShgGR4kaK0D7Nrbp+uA0Ip8bO/hYddtw44
rn8UivjBYsh2f34hUdljH/GsLEy/WP0cSzeJ9X2LQb1PRlPGGbsx7wpDElsK
v5c5YFLahJpT4QX1OQuKV//l3R3I8rpSRrInOY/HMwgkt39CvGp4gs/y2SL3
8ydI87hJG/D2dbDUVkmdxTmEsxADOuGHGl4ivtXkeqL3Ke7oX9om3+sKQww1
6QIvBqpS9coCKOUHGnj7uEla5w5qthvBSDFjWQBhrZLuduIEj6pO4o00FOdc
x5SWhnmDreBIYhOnI10VQcnUl+gfOslmJotgoLes9xE7qQ/auTbGByHXl92W
+6vNh5mFjo2S5jBYaoGqF3U/2LXarXFYBUykIeaGMIC87RVsnhowYqJYUrqU
BtqE00ghIqLJwLfL1uovqhBHgzuhTNhN8QO44tWpXD9jJgvnk1dgG+rOdEgD
TQlXuvnosFoo14kGqR2ytu7Ha1X6VHFuZKc4aYpNsXursRRax0uCPJmlrG29
lt3Ndiybv1YV79TddBsVLsivbxV7ucIwT329YEH8J6Bz05MKFb3N4rPP0Fid
3j3cQN3F16xt1yTZUjRzYMyMowEIiC4qOWd1IYD5veTngzeNJRdhiBHNkzkq
HLLeZ/hDtJHllesxMG+eK0DVLnJV3uyu4RVJ+4S4xMZNOx7cZxw544gFkEm4
tUF+zLgUxJaFeTyncPfOtCEGGC68DM3ZHnRJRoFMt8n08P2nBL0/KsRxG0lx
tkkQQZxrCOkwxqruy9cZKn9g96alYmMZDC+QA4tPOJb45vWFN96gRCDnKdKr
Reji08dj9IgQ4uPOLQA/EqIItcis2cFJG/YbD5Mzd3ouEWNKhQ6RJVPK1gwZ
ihTkEs6FW5jGYZJoRQ89191mOjz9zTMzZSVRadgMY0CAZ4tinWOYVWYeuLTU
7fCh7L78bVUDjUvIZSaGvvYRVo6SGMZgXPIAWXFGWoUvkH3eYWKka1O0jTby
l1ac4kqm/ACm3G+yr/pc29J8HkQ1+4hf9/52BpIMrZwZtrCRkGTPrbNpsE9P
umUwcYgVAU8/RW9wWYv1+7ffkN6x4dAQlN9Pmjksc7iIAMA9Qw0kH2BN2kYy
VjSDe+nLIW1Bvs7yJyxTTy5UMvgKXpPAvyulhMkGRKp4gfh6l9HHtbvOlHIz
bolNbavjOqj5AgJGE+BsctAJelrULvvFdGY+/4DWeS5mPxGPk9FH9bVmcpp6
VxcnUsw4zIchAgJ2nPCJ6s15KfvFohn4UDW1aPWyGlAMZE2VwSqNNjKULNKc
kOJYGrUlMlL0Dqu1c36tO3xZFIbT3HV3Hww7SDcg8+PYx5RemhyQHAACcTY5
LLvJPMH9wFbnQtSM2+IwVb04/vI8pk3sE6bBHGiw5xfmM3wIB1j+nIZgRGpJ
ybTLbV+XgCLBkwQ4hmfyFXvg08O6BalXXslqQ/9oIiL/4oydwl/KcRQj2t3X
mRZt+E5dNxsC2hjwocAa6l1XPNkEeaN+Vepe9p111meALAKGBOiUDMnfl1pL
V3rnw+jJ4WKh+LUbS8ChOjF+WZzce2CV6R6P2/HTnl4RJRLcvxef2iKqH7E+
yW9lu9nFPVq4/AHY7StMDaTIbWJb/CxDaxfA0ykgoPBv325vlZ2AvvOQWOyX
xp9FM6IFUq9I8T46dco/fGriR8avxF/1p17sCnkvCXGCKk7Df0muRrcyZV1R
6lGfKur+j+KQqyzvNgqCDtEIkRmSU0hu/zIy7LsYjh31C3gd3U/bhyql3sbo
z6ooMRnUAHnfn5LUt7cn/DRnMpKtT5HmSr8FeAjcfmGmKaQagUhumdlHw0Ke
+lmD7l0A1iZPimq1fXlojqMksKANjCgt1f1bQLjPgSNVuyE9WTLmK5PVJpU6
5QmDoLym45DtIMHXUG+FGAyoUVrNJr9JIZ/KAHeNiHcNN72+nzc+sGL2opja
rLIimIWpUAnmvZWflq864O7tUpGlvr79JAPSJrgKwuHVuEc8yWjyBWIoSl3o
YbK8eq89M7ABGwCw0FWnW1LuhRGg79maICCENzSHldb+RJeeVLkQvGWbR/yj
M42LBmZ0EHV+HfGJVxBzLFaJbxuacs4e+1ZW+xb7ZobIq91aonCJvTA4f3Rq
q/dmjv9NflFs/AKP1OKeo3I1AJvBfPWGylCLmg7/5oddvKQtgPhtzzEh12c7
DexsaxXSmxhvaiBqHuvE0q6iJED58HLHR65/khSAmHQeT26V7KykDGsKf98G
E0Fm7vCDRD2nRjuQycK3IqtYzYMCQC7drG4/QcUqwD9aV/1akB/HDhtfz38z
Gb6BbEDkppsvDDCOnhJ2214I2NcwbLkJ+jJx51UgmRyx/I0jUu1ZPQO15R5U
dJmA9qQfpcia+5DXTz8S7p2otrHyiPD4NnHDkynrJKzDP8B2MoyqBpZVk8w9
N92x0431Ql9xbeMwELLu040QMuDbZZlhDJ8QqQm/ctLMCCxQdOu8WltKTZUV
MxkG7/jMda1EnjZI6v0xuRYgmke5YBCmV3qx+6M4yTTwKWRq0Sc8/eSpCsNX
GwhXAlmZVvwJjUSXfDsuzNoRqYCLjvI6hr6Xd1U2u+BuUrqcYYmvVTae5l6Q
tW6p1naFLZ9Xs8F4TBf2lkqR4FeJZd57w9ESr3HfJ+ChRp5Xon5ZtdObNpW3
aKvND3vrtSQBlVrmtiAbC9LWMuDtfKjJIbRgJLAwj/0B5iaOXuuuF1S9FBay
kKXtN8NX3XonsReenl1nJ+rTCfu8SYXAtZnOowG6QWhCPTSZuRSsUARYNFpy
iG3KPERoFQhXUGyfBPi6tBZknS2D1R9qrWLkR0fxALUBwbta5RKbQh1ETbHS
VQgzC7353haN+kj2ULyrQ5KF1A+mrnut4zGX2oCJzBqXn0wxLoFGBIOL87pd
6I5sQgHtcBlBBdMDLeoD7q4cC5vD6mpelHpogpjI5rB4kRbgAKNta9Q5vnYy
yxS31kLCHik3QteY86BchNYf77FlGZYCjhLDaCMWL++VsmbPeeIT4ZXQT2Er
VD0KixVe59PV/NTiY6+9xApThCKigmirUdeLXw/3J6T6BYFQajQgPhEjIF/d
cqd964cqt7S9Gt3YwzDVNqtnT8o8JRNABzjExMDsopCiiHemQxUr1bw9TYz1
rLriSxs0DnM61fio7DcqNXIPJgfprnuGR1xbLdqoRD+mOFoLBk1cwg3druCU
1dtuG5JzIAx2lQx+FwexC324ttCwLeaszNC8UKMee+7KthxME4vB7IiUzDz0
r7KrkcyEbmnl9XUuVoFyzXsaZ1nVvaM1knGV2dwbooGhdX2A3d6f/wuahNSQ
M75RMtdVQU7QafsN0DNNWnBL8d9GWG222IHdVWV0FMvE1AliwfYEG4RF3AIX
QvO4SvXPWSS7w+2OgNpaLBrHYt10W2bW/JRLg6Iwo97d15ZB7UvCAiuv3X7Y
4PmJnqQIgtOmy4A0+hsWJooLItfTtoxiSjzmzLbgTaNAxq7nNFkqR3W/nTJP
9rC+y24jE2EN0j1sizKOgDiriLF4QsUAmszO7Bx5CVrfUODfIthFvd7jtE0A
//+jPUF/8s1gMGrT+jNTIpRUEJfgnouIHmcZHevuHnaUTEVqjN5A6+2b73jb
qP0wEmxTMwbSqo64NA9D2XR1bSanP6kW7g6jVriyUjiW8rAbqHatyBbwHZY0
6cYUB+BDScT0Xf+DNV1LmXcn5Quy5mcJv6yLD+mV80qxDrMR17pZwk17LNyC
mRivHLpqHKYUBWbLjkToZZXDUq/xRoSYrlIDedpZ26tS3fcOx63t9iaDnQ8d
jTwMo6Ef1vu8vnFqt7HoKWyp+OurSjfiz1o1G1Shro8oWxIEw1I+tP4Vr9w2
Ik3p58uuDRJKfdCBdG8H9R45qm9SKOYbIF/CiQk/S5HIqeKCt+2anZw1aQaK
aOh5fw6Fh4z6ZYJcjONntvPFRdKUQr9m1FISGNmyKe9Xtv9A9p+IW/hphiPS
5sYUwLrmJB3J9bcSnyASi5LX6smKFVMQi/mDM6Cb9sBmYOmldyzL1vVTWbQN
txS/C+EaImvHEK6eAuIoRfqXqwn7sh86Np/VaJPz8ZCGwqxUshBhelDqbxJy
63I3toQs6XLZ90NuPtyi+HL9LzWvTLGwF59dM9St6wxYsNQUYLqiISrV9uTK
JwiXX1Nms1S/pHKrj2oNjhHR+NhZdQG5zu8K1cOb6DHC+PVcRC4/4UiHsNml
Y0p3I0jQ/0uLa5P514KgUzLobIhfkBIh7Tz/ljCp9tAw9N8X0Z3GOlnz0hvf
pdu4FVamDqse9gPjgHhK8/ZtEtfUcS9bjB3FTdhjUmK3pPIM9rahGaLXlK31
SNDcsOtaGpPPlrYD8X2nGt+UsIePzw4hR/Yc6VSEv4HSBVraNzPwXuu7lE/7
8TUysSvFPMJPVKRqnKkpfAYq3iuHWuzhaxmn8cfzLMgFq0VmYRkD+Jjp/rgP
UIdChFVlHk/N0Qlk7dz7HUGuYWFLByxcxcpKEy/M1pB+DWZyiVfkzcFIUILi
uC201FJDo3Xf0kHDPFFoiTk970teo9Beq1ZoqMaizVuEmFXt+2/UMc0M7N5w
S+WYIWoDKUGQwkNu7x2E5fhnhMYFesOajB3cLkoeK3F0LwFJAIhjEExnGVfq
hp6mbYfz8EaknRFDQb4/cvxSEidVQbRT9tNTUzId/4kzymc0YZdSWq8yO4Fl
f+Zz3GCF/yahwBhk2NoqUOgjSMXu7wbD7xsemEA8EL0rxorfkn+zmn1j8kTu
ywxH6GuW2SJR53qmzQQvobXmBPDaBDFVn/SEYOKsHVSdeRpTh+1hgxTW4yHq
SXr48z6wbgQGftzh4BDIHfp1oIUWf0vXchtOQ1aBaoyyso5vTHlzMWb2yTL5
u3Y7tZheXGb3DTsTuGi39AUvgNuJckgqTC6VBJrbUuuzu2IwHc4Ex5gtVyMj
NhC8C7eejva+PmIZVAoeOxkbej0WK2Tk8dt5ljRMv/i/fN+9MJ8TtveoVN4N
LPlRdbaz5R8CqVEF2RkbktOFEAfacmGKuf2qzwLq/nFi8T1oJbbVPoINyaaa
BFQxhd3H9m88n+PxUSCeCtWlRzflSeUANzVNBTVftPMc1iR0U52P8iwNbKpW
NrtqESxlFHPNxKngjE/ja4fV+0hnRrevq/pCyrbyqLwOXm/wwCxQnNg7Sr01
5xqML7gNEYGw4BTQuJit3AepjpZOSxMOPKSpOQvRN4uDtxgDpuwD3aH90M9m
IJ33IF11F1iv47uI3epF0OASL7j5cVl8j888IpH+DtJCJuY2JYViguBkt0Yc
whjT3Zlj5mK4+EiHZP1vQv6+f03OUgnw1/ZLabRFqrGowZEvbVRYFYU1rqTe
t/5pgJifzD6rXBEtf3AdJJMa5XiwI3vcQoJ2TkkRycX+sj3raXg/qBjkJBtT
NYIfqhMpGzxaJjD4/LtTkJAy5TX1EafpPncRJS1nYDX52ejkD1Pnd+hiRsnm
1Kxu+dYQCymdOkWnXmTQVWbsb11M82PnOUZJ8B6o7BlkyhhX6DO0Xpu2Mj3/
ufTG0Xg6WxhH1kyjON+WxC6ktm0sUmN3MxWHkpZVoOxhSskOflD98VF3eJz/
A3fj8M1Gtww3qBDeEMykxaLD89gCZaMJt9tO5h86aNwzVYJJJyqmnGODTP/T
lxza3a+bwdBfW9ObWjEpycMIRuh5GUc6ZAQMhTtJWGvuFkDJxSqcl6AdCwpJ
2HmnFuVRgIUvFCSsHdFRSLLVTLJBt9PcAYIIYumwPsOWhDTaCGZCnBtZ693+
yrq19o+t37sY5J9hWvhUhJyFfJR+IOBFv83uHIhqEgMgqewYmNvHP/N45yzL
YDQYnt9TVpf+vkHQmwp0c6zTYXmcGnbfsE8fEVXbYhDY1h8KxcUrjVq9iS+X
cSiDIUaYmQP7N6pje7mNsQHumE5qEaQnjIauO/LvsnQqBsO0ZN+ZYr9tHlec
28df7QaOQS3hu+UXW+Ypr7QnEfHbQNma/jX+Lz1TKQtNCZOI9nh+a6rifftn
wwFoyw93YsNWgAPS8T3di+Fj5XdlIkZNtRNQbzg6g5thUj7P7edhnGAAG2AD
KgECElo1LpJ1j5SH1Qw/Hk1P3SS99Fj6cwfTfXXys934aGxljpmx7CSNF/GA
9Xicame/LaiUuv632j7FksQEzzDH9vLbXfYlyFzDX5dHmzP7b0nWjkNyvxtE
UB/l9FXN6PbBYwnFFmxBGxlI5JX6gPxNe576Xy4ClTJkYE2wP63j8jAq3Whz
EQkFldsanOUNptfBDnngZMrQG+7Y0btUOUZyV0HJlKYEPZ6lwqvXO+THAUf1
fVv+uIEfMwHRD5ENidynM1SNELbY9M/CMpY2pRD0wrG0XqxqsQ+wE0a/ZzvU
MvPc719LQREKiyLDALDHM4K7E2L1gk08oggfsR0ybAM5Ts6B/dHo6pR4wXvo
DrciUzzVX9vVoIGrYnDpLIBRcF7h5gkjyy4x/E1GX3fW71fnAFVe59fONf4G
ymFqpsh/aZwVRavHLlAqbWC8rtpk35LBya+BRptnWKi13gXvH+siLCiQyG6X
7d9LzrtM9pLVTBirGslsmN2zzmXBlQKRdb6EYPXjZAJDWm+WDjoDlQmjW5Kv
9i7MH2qwHg5qnIoTba1AihvLSdBFtwrV9ssS02BrpQ8GZ7MuIheUyVSDSXPi
MfVRn1GJqkqI/5KdIcdkqjMVLVh5Oj4AAq9RsO9t1pUMZLbjfI/52T3uJ6NN
CAd2NnWpHr9YM5jhsCupC5wObxBKNR6xwcdJ2cQES6BpgzHAhCcGArlft19F
//ifb6iZnWuQYtP9OW5zO25+dnx1DbS2diWokrRTkHS20/e+uov5lLK1SYs+
GIVJ8d5cGHNpqcuFRpV2qU6yFoz+Rb4pWAbCim91wG8JnlkT3pr5ZrCe4yN+
BU76GcHJSAMAjGOdPZLExc/WsJj+B9NAs9I13qsxmHLyAeYh8EA4dvTUfsWS
W1xUV3099FMS83Vwgi5BW+V22ZdRPpeee3Qxk9s2Mm2clX88Yr+jtPhhzcsq
AxYCf4THfLLgxoJ/aXUwdq3A75U7DHsAzYddyLPQOxBvjxilwbANKpki0gY3
eLFJMtN0ZRDnnQlMFzeBURXUuj7049jOu0Mzcy0CgnvCNm3zPML8Oenya/Kz
ywIwXwNylqz20s5biL3EEYC3rbhjBYU0FJSLNIolOM0VWDwNrdC2sNamxTna
3dp1fPVYRRZJYxPOmPnVr3LL1DSDjfWQ16omi+tJdh6JN079Gq8lrZ7WcgE9
BYKm7GXRPePRddinqfcWBw750OVXq9r4qZ77Hp6ihV9vXQfH/UmMSmyGUaAN
8R7gfaMueUeKYDqtECINqkbUT65oEnlvfNK2kdUyOOudfZMh1C2AXXQn0+2u
vNvKuA3YdjyGLpNwiW6KeIqTj/Kc/zzSm2JlLqWHSKsM5iHAiruKW/nBPDQH
TBr59Nd6jfpcJffuglCGTq7b/vVU5pHdfV7vwu4UK3TJIR3p1AnGbtN/vZGk
znyrl8/rC7eLlUVy5Kt0n5/HUfw12q9ExZTJlU3fOyWZSEpS/jQbyJnkTRHq
H9tFLpB/NqWHDF0qfdm6YmG/XgWh8PUVfRS7cRjInBw8nUkDHGDpPTUo8Sx/
FmNd9QjnsnejwOSuUK9bGFv2B6bOCdKfxdL3F2hqSlIdEkFEvQfi4RSUNOuS
vvOKu1HydnXylujDNkiB+aQdESoCENB/a2Pe2hhusi4cCFw9d1er/XTty5Gs
PeoT4PagOu5g0Da4kcITwnvjnGuwknjuWIBBL0vJXveR+UPI/1RhqA9zmxTq
w9uA2r0vFO/RjD38q1+y9CzgWHmKELBt/U7KTSurTmW7irZI9Lo7QyltOpKY
vUUCXyLiuGp2HvPG5Pvt9t36qnk9IAcfKqlTq7owe5KhhGC2v+PdPI5lMVsp
PQDXZiBGaHXY9wnkJy0//a2e//hx4w73CdX4WJDRXecLoZB8Gbb6Qwus2i3L
iQoW6ZlQO9kpUGlrrdB0uM7S5rge5/Pzp+XIejk3hi2smWGopddkXxApzJJv
yR7Ho8uzPxEMs2JpWpTCap3J+/bF5NVsW6254gB4AaQQcJnHBD8Lx2Je6qo6
H1iZLdensR/osZFMMUqOAYKbpGbMClTHzhhC5xzIxafr7YFeQfGI+3NeiuPQ
dH4LDBIoOyP/UKYIT6DMh0gVHpZpO0vCPvUKm22LQpGXw0bL6wWAP0TG3vyP
F66u3aAqt7BM5q0yBheh0ero86PQ5QhHl5JL3AadM5uRzMJODPAyDcuxhF+A
easkthb/lsnPgNFQ0+LkgfbNjiIwgiLcGVHIle9AhJI48FenuwWXBmKeNXud
tbmv+rIa6ji6BQtHiSgddyYgvmc54rBUEoPWDnVX3xxubFrNAJMX+o2WSLH8
PcWKpahrw2c9ez+aPzf0tI3v7ZDUFv7SZ1WNVrtHxhZpzPO/+j5VnXwPUr/H
zUKP7REIwn4t4zD5axwSYMCX+08MErYxxa3ZSWArzqln5Caey5IsyqfFsiPJ
4nfE6gliOPkXiTHORq6xjTRJl0F1lOBB8Y9+yeSwBb7DG14eGxyTZhc9+ddH
0c1MW/WxdDL3DIy0xkgvst+ACjive2luweH3v30qaLYdiQybEHC2agtWhYmB
cdGW57lvuNBVnJfhqhgOsCIidCEO7L0hxcBYvekeTttcCt1Vva4wiSfKdEpW
G72NkHDvR5f4g0MR/yuaLcXb8ue2RZlkEfo7dskE9czN670Ovjfn31HK1I4H
xvry6I8fDgJSccfS4wiQ3E80fNpXNk3lRRPJ1/fjfzpltR6ut6AxqW6xPdfx
gld00S/JNQlg1q12XI9INhek5dOftVb6fOhoAQ/LSRXoMPyNuZbL5BKmNZ7C
GOAI7T1py2JpFHsOUUUBo/S31MvjIR0CKOkhB5Oq1T2uF62kLyBpv3DFRUfy
7O8IHk53Ctbv+gl4DTu2TfihT5U7QLbd3wUk4qz1fs17wkVZxm/1pP4l0G9A
xMKk6I9Sa8Y9MOECyvv9lHvz+4l1T/Yev90n4BDUaz2MTtYGW1GCB2hM41VZ
St31YMMqx/Me3eqbqmu9LmNLB+rTPtoj/nfoFrEo9BX3AscPM9DZ4/uQCYwj
RsLdV01fwuJ6JCJ0VMsAoi5I+j7gRoSgV4F1HwyevgIMiHafio3xOejBbLSD
l8CbyKDLm0/Fmp9QIAPKzjMUJd4YgfftAF6ICAFetxYavl7p9hbLsMwOVoa1
G7tLOTxsIxhhPvWquMv1jrIttjczQCZhueBRTqt0QbPRQDGMwUVmosQUrb/I
qr/5AOFvKJ5361UYmAZFGMDtPAMsZiVJ2FNZCGFDG/3JmNzQBEz+8RTyOAAh
mq8y/2NGygOka7L93xtkURHhoqegDOfeJOUdXm90+lsDl3fDgjRwj9uY/ylF
pX3jV2f3eUsbZwmSbbluD1ybFRFLQTbZWjcsgmqcBcNbpo1CB+hYyz7e5mvI
92O2OUOerXYI6HuQTjRRnRVAtrBbTNMfV3ie/3WfDMqvyK+CDknNvoMclF1h
TiaFhaIv2xiQDC4UvZ7px+w1rIR+a9jI6iOTXfJqRTLevXbq4AN6y6PF+2bq
6fwVAv93fdUvFqRAYHrA7Utr6g+Y9l1pGcPRX4aIv0Z+J83gjDsVMCv0oNao
Rq0SVdSM3DwnAu22kB2+YxkM1l5yzCjtGnoQMZR3io1QXu/OmR7K3zMXM2U0
e2eLqaEsv3UKdd3xkb66ITVYe5JopcfGZ9QHXQbwDddf+KexpejIOI5gDK6K
bqjJf0OPwe+MpFTcIwlSMIDZv58B7hfcLPC2jNYDXmeVWiqMkUn9btIb67hW
KJCXZsYxcLWr9LI7UBkxBGrE+QC0QnxmCBoimk/3MkNViQ8eYqpSAsO2fn2c
lXxg+R399ZpcqnZijVsmMgwJasZCjCiOkFXLCiTdvYp1tuS9ctCP8gIOHChP
II315llfUEJxVuoDs9lVlvd22tPeuTuHHCRie+mEeqbNLFd7IHUPRCV+49gq
SzWxpskTvwQlPDb5o5YbUqHE+WzFnAM/axsHIm6EZCZzhT7V7ZL/OTFX49RW
92UiefsJ7uSH5uyZgK423/XEJ16WYkpCIMCyVo6SWyaRqZjjXS5Cx+1sV2ni
d2QmAemq1h4gcqFXRmzSL7HHEN3mCvPZN94W/INe2jU9Dz/pHckT/nA+sZ6I
Dej/SK3fOyOzsIYBBymkj46cbpwLj/uNZEcyl17zNwPptF4hORq91lMg7rOG
32DVInKrhu6H78Z0EL8vHjub8nX1/hcp81Cea9mQ+HmUT0cUXUSDiVsSiLSk
tpa1DRJ8wzH5+K/Q7TtOnV+0+hJmAd0pv7CnCdDWlL562UkvVt+JUfEz4SHN
g32H3HVCJVlY7OQqKJW7LwL8WuYJn0ydyAXnfJlWCRH76tkJlnejg5+u8scV
GYsomnrYHYd0cH6zJtyguxCqVTDCEBmtfpHCTSj0xmfx1RiBMFaiEjbWW7W6
CCS4FYSoepzug8SIxskiKIe9JiGDk7GFYbRqWbNDmph5QTsRe1WQT17VyQfY
iOzuDk/6VBUSDOODLmLQj2NhazLPOcV9tnBmWPnFBmY15qSQupvZSxOdfkR9
w47sCWM/bSEoe/gFyV6TcAoJXCZ0xkvoYHW05HIix1ZNo0+kHJ8LFYwfy/bZ
NU/kT/CYQUDplURxH2JWF4541zTdgwcAU2C+TSOhIfPZ8OoFF4JBCTtIcBPx
T5/qoMh2blAFzXaOUoea5MwqAGFXta1/JNr+8w2vAXBRszaQXaMixfcbW0Md
cowbgPLEuWyEpHrbzObtcnDrT3aPMmF4xtyEdy2Hoxe+oEMImAtvKRbNroHq
tE0zBHqFQvOPW9QGZvpt+Ybj+60A/QsBYXwO/sdDAH6DZXXvh38iBG4Qlrss
uopKBHwohTRRl12vTq05hixghhP/A2jnJed3BzVsySLvj4mYZV+PycQ+XAOm
HzpuG9E/JfzY5Upp7/tyu+1Aauakp5bQSxs4Tjr7mUMRNA3WyUy/mmUG77Yn
IDUez5cmwZ/GrW+Ku4Xiy4rnSh5rJmr8gzhigCL52Sksg/EBsZtswZhh5kbC
MZnnY9ZBTVEjkT9SWWn/NdJUUZ4nVrLgDkf6EXlvgSKEogpNQT0aZrbJG0y6
g9wnLMNU0/Tf+eXIvmO6Ys3FJxKityGy6Jz44DHxTfvaWVShwmM26wyKBe+E
qcicNk0p/6Zk16Y8UcDwK947BemxQ77cRjVbA4XKUvGJ/WZQFgWH1I3JuHNQ
RwjP+qbv4iek2TP3rlMaZcDwtCecaCz4uLR8UbrG5mUfM9x0lsUE9Qa3yH+P
237S0LUJFnpUHVJ33nlRuRCseUKQM06khCtLwQNWWS6n5ApKxhDJ6UwRNpkD
iXgHGzNlv46hxT1QdOb1SSLtwAO0RQJ5RyPXJMDZJ4hFNOBsrXtZxwYR+aSn
JUw5ptplto+qQli/RJMyrxFmKPftJIo63x464winkJXsGvInOSOrlenHQAct
+2BVxP+e3FXbQblMj/w9Shonk4kx4OuOdCPAI/xyz3W69Pg4JnJDBC8jZsMn
I8IWWZZ33lwZbCyh45Zzv3GFhfvw06EDufljpff3qLqu9QvWxghPjh9yuERS
m7mVQTFMJKVjUw17Gh02g5Mpg15ewMlsgw1hGeDrhdlBg8Vr+5KYNgct8RmO
AFm+wKzwQXf+bV4Ona+VYxIANteiQ87vjM2M5roujsSCpEgH/fkm2Fec0Gr/
4JMVDsjRTI4tn7T5boAT3fK5neAKZOMMPkK41L825hq9ElBDvqypbRCp6+Vk
3rmIZGg1aGLoUFPoQIMbe99qhB5eifByDpuo3UDuI2r2jqIBM4n/hQvT52uQ
w5QsvoJlutR06nb1O2MyVdtr/iTj++q9c/sVrsxJH1dJFMlSSnKAxKu0jdt+
ouJaNH1syLDpPMLAwjjBheU9brkC2Jk9qjeg13Wv4XjvYFdS+L/P3QUuopzR
T4xp2pgJTIa6jpuy1ak7YXrzwwF5SZcWM9+sSo8MzWDA9WHW8dW6nld7nCiv
JLGWU9PC6hYo7OBSfAo0ub7v2CZoS1s7M7c4+f7Jge5e031zJbxbiFhjJ/dJ
+52PDeJGlhsjZtS1iZvtjnUFFzlDXOdi09st6Gydvj9KuXnn2Wp5ihl/iHeq
6WMMySRQhVuK/2BkIM/nBW6ZNyXKIQ4eoQ/jUHsQuKzzay6IGnYGr7ydmuF/
3Q9JGyMASvNVdAkDqfe9SOkApKpxCdyfc13brNER+uVtk1CFf3qb0dcGWo3X
QSAkSDkLMwnLD/yPmzOCNEfwGTKHQOSoLyiW26wfKYp79ESPvoMzNeaybGIY
RLJ83uTIoOHh5HzEoQPxq8TpNnFVk956dwIgDDMPBoI2LNeNXxie4nQ84kTI
i8UA38qd94k6JNyr13Mg4uZkrK2zzlKoxgd974aizTLG8rURdAQ4CR0QBJ32
j7+MNMmgnQoyzUtIVa2GIoaab5MYWndQqFh5DdOO72cgLjWZSHdI6aWvNlhn
mzQU1APbGLFkEzswbllnZqL3zSZudR6Dh9ta2Qdmyws5ELKHx+UXh60Ilyr3
I1ipPQKHqRilDSalQ3t3YWk7j3bmfnuymrg2EvK166URig6JNOJPDcfqDpaT
D/ly4KOPvTcwGYxl4v6eDblP6S35+9DsohmDR/TOOOYwToT9umB6jEmy8n7e
dOBL1517GYRzjm4Gf4GuUuePV6VEEsw1CDmtExL8o78+F15gMgq6opGpw2gV
XS6p+QPrXpI/sSXIal7mpgHm90XLDd/XhvVqcikxmqXDTDyAlZYSp9A0uj+K
C3hPo695tyHf5NzVsoNVhc4nEP6aZbfHuPLV0sGsq6l7R5v/TOUrN95bMlOS
QsjJ3R4fApG0Ouk+Vw+d39DibauAeG6Jpr41xEMq4oiYfiFLjfLkBDyMEZQM
A/YgvB6Nx70dQSYSkydLP6m4ZOVIWEoRYVNac7TxjV87QvSf3syhRu2dn7gr
UflOYidxN07jh9b7eSx+TMzzHeSpfmpy3kLNujhzsZM6iLlfyspxBeqLfahW
92jp4zpsKlPo85P4Ve/nZfwJ17uU7UgflLHgYs17H4SoipdJlxoyEgcv3XLy
+TF2ADFmgNFWxtkIdcpoSo3giyKKIznzCA48CT+0N/L9arNv8dy115B8FEDn
j2aii+NoqQTJZH4yLPc9qnWpArmKpAtIAI0Vey3GV91XDhuWSFpeThIWLqlQ
Kn6tFzQUx+JO3OksIFiEwPC/7At3qdV24+uZLs8gt2rwPnLxLJX2K5OF6Ep5
rHDqsMqhT29oc0umt5cj/eZWmc9WT1TGxaUDv6IKVeUeojK4jEJFDoPEks48
ynBICfeq/UsawY41cShrlxhhsmd1FQWp2sePRL9X+t2l+krLWMJ5523JEmmG
wphlZ31eZ86+Q/bHGIS+WEeZdO3+hXWAumpAhIlcVzMWoIuWSSjPMvHb2j/P
grWZ4CfKOllFqkKaay2z25hUNFX5JnRUuS320KEXIiy1zvEai1AlIsRJ6oNy
nHW5fdC0B7ShEywjg3VPLjxYG4hoE6uo+z76EfTG7DMfSYMtYgvtyKtvDYTM
LknbBSylitOfay9m537LX9Qp7hFh452qnOn1ybTvMXpuvxVZLVUWM3qonxxY
hK59jJsXdkcPsPM/qMLbG4O19U3cEgjh/YMUIFokl6Ci/TCfl652UvsH5uhB
s10+k1izwoxdP1NBAgYFBgNebMw1s1KXdxXicJnumcu0m8uBWCIiAFxniMLn
XRA9BDk72pjEpQaTqHIzhJDV1OeZMhfy67+CMdRiK3txIfR9QAU+Cr/PKT3z
K1ULZ/uixgkZ2UQ+OAVAgt5ZCnoxyYowaFN78zra+blKGHRjZjIfggUuS46a
Xr3RUHatsPSmEJ+f7uLKFCWnudmZUAORCJKecAAHBHg4aRyNc5h9gItC+/mD
HrZ9zUg8fcHNflJfBhxx5KMSL+Q/qLfLGMs3OwX/nstoeDUIB4gIHD19IGfo
SlBumUYou+AMxMwvmbmS2Iv0EWFI+kEXN5zq/ubIutrN3s81b0bFEuHTmyyx
XXwrtVYur/U6NydVZVnw+G900nz1/8hZ9eTeWTXsxUBeWHHrtu/TKdJ1dt5U
/AT3HV2qmUXNNqQmgCYgpoLS5hvez8sxdveuenlCYVxGVIDIrbrsnEQEFQ4Y
8YoFu8B4txQgBuyiD5D4lPliSpOVskkJTsHLfRdbF51blKDLxy36ES74gSPv
oPM0OQBaauHEhZmG3U5SwSZXexK8TzCEg3N3/6cczem/bsTPIZEJNujktx9u
FxNY68o8WnypAbgMI1bdBB0jXkg888I3oMIDS9uJpvOnntW9xCbxhAXqtkyQ
lLWQ5D19VCoesbznqUrUYQ9cWKpuqL+zB0a6C5T4J5XCHmIkzmGvpnokpw6r
2njhx5FmMZ67L+4MOWcpDr33wklAiwPnPU9hHF3eQYRlcN2DDeo1zAcUxTss
qbsbCbCVnNPQfsZJ4uCWcgaaO7UEzm5qFpdEB0rgH6amdcsGvTmEanYISQ7n
aVg5a+SPitjyUDjnD0sONQQ3a8I+vfAs/toUE+chJfjUUT87nLqggxwr1sMK
iP2zwDgFzhNrDsjPVYHPF0QUxwJViAtYeELODmQmJAJU79WHAzYCcd8Cvkz7
hAzpWMxmXhIKvWlo6/YK63vrKcm+VI1CrrWSAQdGXIZzNvLhH70Sft3Mr6Z/
gHrsJwmNfJaVGsbgXs5/A8kz48Lrk2gamN4/2JqWE8AXAZ2ESIA9egZWuIc/
FjjdnOwf+3BSZD0uVuSUVpDpUqKyeOI/lMMttD///Bq0tCEg5dwcefvRcSUI
ZKWQ2vskKK5YNvu3hPIzJG/38/7p5hzwt9Q+5p7F3WI/c8qm72iLISMvD5/u
WYvWwfuyGET5qzK5SAuFcJbdeoe3mH+X+gzy3qFg5YuHd/ULF/NevwmuxAAq
aoLH3Yz9GbMksyOx/FHlcey8F++FR24ERoLtOJ6MMLjvhGgohDPus48IqXbX
cf2LseX7P4G1qjzHYFZ8Q+gNuv0/pOLn0BIY1+nQg2y1tlSHsTE4K9N6ZElO
YOj70sduaSsSe0rNhm0xvLKCP3gDuz4hip3s9q+Qd/KdTrHubmnDDCEqQcP2
zUWT7TezUvFhFItzO4yqC8z4/vbF2Eb8QeK2uAo7wzl3l6MVMCGlorOu2SQG
PqFNo4q7AJxPiVAEAhxaTufVi0P5BCN92ulRS+gNiSfRBCknB6LOormFFVNB
OF7byBsL/svt/txasQMgcnorciAnbYnrzq4reNjm/ZEZ6+tGCNCsZmg/GrTW
4YxAvl/rXXEWT99Ct/ru+r9xDes98cksqOpmBpzbJ1Tv9DW0jAiPnEznKvLA
4zsZ/+K5+/0o/6XAhDUxcP0LhiZ6iFCNqeO08hOaMaQ2voX2qvz8083fdBJQ
ujqlLJjrhj6RGDWb1MbXjYjUi5qmDnhhWopNBUsSwegg1lN8knIhVZVnoyNK
WpOWbsGMK3tsiStQOaaZiiiHCiQJv0arRmXEIuo9lhhs4bqe9NM1cPVBVH6Y
yfkedKYFRGHWXA+Giuur7QLFOSntFOsxti99ue9cFc1LqG0bzyU3DtDRheGK
WoyJa+mAoSLnDTCyjBdmBjyXsBolCYtRYpyv/xxvYqmMDaTr+qGHSY+Oo6gL
8UHEC29N0Aao5UIzRlTB73K5IkoKOuPz6G/NjMjrXN5RPgAKDO3wNvysOqHo
SD+NQfnU/FInv+BWsUbglwsN+2QqqF6YpYnyVRh3d5l9Ilodo7RzoS1C7egi
F3SDKHNakHoSOhirQQb9I2qEMWt1+wHZurcY75XgfsqwFvaSEGrKlY86XkUK
e6zrUXKSBJ+QakBdqIZ//hkDU/FywrY4lvtdHzK6AF9oJoDOme3rFx9AGoDA
pM0Z34WSTUB1+Wbz9cmK3JmS6TftF3W5wFvR97nRtdnH/G3SOZ4J+DogsZMw
bHctj2s8k7qB+abkOQ5ETKn5MFCpNPkEOr4wlqxPMZKytyJeZFX94PTy5m9i
P7XDcsRxJ8SDuwD/w+uo5u9Ma0tjiEkmYGi9VQslgA6rjDn77PsBUPoj18jn
WFTKNGyRUGGepnordw+mqSORjvsk6TSZQC0LdKw2RxgoV1gYqZMP30uzZ2bk
RPa8Ii+xDftM+YJGJGECYThIR1lrlumjkFFSTzHsF8qY+ccF+iC1Ctj1mDht
8+xaBH4DfNeN++N8WPNh9Yc09Pem78rj6DXLsGkckKABSdq1xAD4g9X8E/c+
IkfDkhij8TpBY1gBrhtV54OyY8SHK/+193ZcqZTp9GAKwn0UUXOuqTrUbwv3
tLoBbCLGyqN/t8Ut+sEGFSlhGm/qtHlrK1ILn5mP9vWjv3qPWgRRr8KcUz16
WQZdoiZkTBl9IBX6DGDaSPaK4S8J30mK2VyTGBAi/0qSQ6YCvFfisAX4jaXa
9LfjoBfIqkOf/Z1k2L0gDRc8wLgDeBNMEuYxVdA7pO/J2ETU6uUQYSEeYd4p
HJ1LP3qZKAmALIU947nghfk3JlwIaaSTFsEg/VoV1HoZVKQL477nbqV/P7fH
CguoI5eq6QwxW98UbGywXw/wb3LQp2mpWfh3IvV4D83dTolOYPhNx5wbfEwj
CB62JArpxYWhDBVbgqa3EL1h84CR7ICOG9WzSthkCuRZU1lIS5BEuPKHDoy8
39aOlp/kHOOAvdj1UCJb1fcHiJMmwCeaBNuSedwyTggc+rwC1coCTmM6t27r
7GMopQXYVMUW+y7H0U4ljOjt8mDytSru2Bc5OqG6CYXDn5fCe9spcT1BhS+L
lA0s034FDuxEMlSza6KBD61WCF1bexGDVgTOgS1A0jVNnYHk64TEUFppGaKD
Rzt83SL+lGnCXtJRsShuNU3Jv7GHJ4EdsJ2bFnpoAkoIPTq96gJR1Id9isyK
bINWNLEdsgIjpzynX8hh/3ZMLscFmXxq0tEvTZqJXD4ngXrBUI46xobvGUSn
oOBdjxjZsf7iMDB0E/IL0zL1gk8PLve43iS+jX/OcE368DerifauxgLXUcjy
MfNpgBcETxLP1C2XEPi3/9+srds9/b86vKJwVRJt8WFsyjMuOMvhUd1R5/de
SJ0uWJyXGb/kNsTnXACu05o0/2exl61xHM/BxU5iSacO6A8m98X0muuyG51N
3obgkfIj0fXLolxaDVYnY2ZEAIOIMUxZRJ9nXP/9f1CzZKO1E074oHN+dLGm
0FPSNW9JBz81MaotVozHDhTI7a+RcjOTobFnOa/CjUzWyL0QCp4v6j4FpcDV
pfkmcdVV8a5/HJvO+ApeB/7/lbyFUD6PbwUBv4CLeQTKuSBwCxefEOjZU0RC
LqstokZ5FZVibS6CoSSOVF4iKZbp6xYDh+aJjzQ/oRKt+DTbLcW8uiA/LBME
/w50EjQeJEbzXWW7+L0WWD+pU2qpqCEspqY4wyceOM4tCI3nWUnn67u97ayo
bq1zXxEH2YJibngIB+OhJ17cejs/F9gEztxp0V4py1cnaufrJNs3V9PW4vNX
G1srpPHDPlatDh2bAu6m4WKUK0NMyteBSZ2UJSLjOEyWGtraaHqEAiHCPTT/
5UHMI3A8rALHdWBNthyul6mN7mNh8nr5Moxex/98Ll5dNdgnXNqF9GWeU/iN
OpaUOTIRThusZHXrfanduUNkxf0YG03UrkFw3ITo+j00ZLxvKWXx45SuEBjy
/uiXTZ3PhpwBKeisBFXBf3ZFqhlcyb1E1IbMhSOmOW9UmaXps/yVAd7MO9Gp
LEtSU6puAheu3uxu4zKo5nkC3qt88epAmlA+ENSyfUJxVpwgOj59EAoLHHzp
wVaa00EhYy/oIVYIOR8D3ZnDEib058ZzublubE9hvgVi3933LZunmKS3YHiv
17B8hUhOQo5QWg8UXNaj1XsrnzHQ1SeMegv0G1gdTMplLABId7px1TmrrSA1
xZa/hjJrBtPnuFuyZzobs6Tk8u23yiam6ze6K4iMDQqQ8+MLNziFXGCXjcpP
JJtxpCU2m4IkQ2FNaIgDrNBwiviwXqEIItpFod9GU+JViqP8vAsHsrYwFt+L
ZmLcxa5QycUqI7+vkqkqEUjYj8dobuyMRPAhOWQzYMyzsrSxiLGj0HcHN0AO
AWiQU8+02UjBzMe60hBX1vL+qdRfjqbHN9kZqTiivJH35uW8cvz6/+ec7HCw
HqFzNe9M3ihEC4JpTs1hoteV1SoR0I2WQ+iuI7OdjqPyIj5T9untwZJ63bd5
bwlzGuLhb0znXxsVuBcT0JHWazLo/oixgORMRUeeSnXzH/UK1R3ctH8r0WzV
56fR8hAuXwkKVlzFRi+x7gl0TlXI+L79Fynu+wdPauQUpOCGnya0hkM+d33i
/E9eSCbpRB2vUyTiEbp2/WUKQXBOj2st3hljFIwobvGY+3XqxiGgk9jQghCw
HBus/Xtdrcz18IiK6qIqDvNUFr5/Y4rGi+vF0Yp6+sPfj49eVWKdZO525Nge
+v3XudqM+het6hJDYxwMZnHGKKtiXGnx9m1euaDWQclfYjxulSwgz+lYgTki
gl0I9lTpUYlSgB/SIgSVgaJOhSIYkBtXs0zo2rTo0EAj2kD7+SjRrtW6grdb
8HuLqQyzBV9wfMND6ROrerm6wuPHIang7Ds1OnTI43ywoChC/ZOYkFAJegat
Kso2h0g6P2uA+UPWbC032Zhh2MTPcG1sD20A8u+js/JPIZUNYWCt7Yv0uHWT
kUvQNQcCZ7xVpwX7bmqb3T4glNN5YchYL25XEVAfJMyxA9VelVwAwf2AzQ/T
sCvHzVGU8/+k+xWI2g5HJ8ivmPGMH9yPmcTklfSiOCVYCrBsIPn233AoUzSN
HRKuZrJq2GZLBl5aiU2eJ5fx7GPMhDckb4Zl3t7TQ8F1HkIXqrzRU6X7HryU
yb958n+vhEANNltbkju29atgfjM0hxvBebqQvyFBazeaKxRI7TBT3EVQ6nWx
bDZNAiH+PrTrr00E14Y9O600P8bYpl/1JoNA0ncFrvftXwe/V1pFqyy9kwyz
xnbCwkD04hAujPni+5JIvghWfiju6qqgvq1/JBzBAX6aoI9smdgfI2iG0e7q
dghmvAp71uKyQiaDZTJ/OIYEa8IWe91ddqF62x61Hn9+VSLPwHMlNBXvXIDc
Y9eSYgPK3ZE2lHVptFSeNUDVh180NQke1S97SMm364xlqAzoEgMXawNvw1HJ
CETyRKP4gX4Mt09SoROW1GtmgLY/eb8/mAQA9vnaIZVoaOTCBswpLRWiVPSa
es/+GeJ0mBuUXRxX1Qc4BQKXS3eQeG0mrPwwTZCXWrw/w/VJzqWCAM3K7L+Q
2VYuRrIA+tGvwlAdkyupsPHz8m53TbzFDLrnJy9dptyGIrkaQi1tCqVEEyw4
528vP2cpQo9pwNdaxgBEj0SscByoqyYw4I0x9yovFTVEuGGz1vDbWk/lOEZi
FSCk/w9RunRK4AFRq1OY0PRiPwz+WhfS2PNaKxM422a7Fyt6kXz11jtGeHAp
lvqR7jspyRLh+7wImsBXFVf7sLcyLMeBsgnzpW/7YcM+jnmZvlWyydfjy91P
DkzWoVi8oSEC9RaIRdElF4NNMwz+J/gZZYGVbIXJlgCAIjhrLQtIh8Owl7/r
xKPayM3wSzeYNJaInIemsO3eCgopdLxghGCBkPut6ENExfREcWtdXLQD8G7e
r7uWUax4zWBYZyzeg1oR05twlH1++eGi4iv3+8deR1tVIVCTye2aaLU0tLPT
TbBhxb0A0VP6eaNn+f/piWYautY2t6t+xvbObEr8BcMd1R2ewrSe/JFJjjIj
fmznasopOzl2N68o12TDer5BVrkRu0vmV85x3y9eWkKCmKhUxiF1SzlhxlD7
GTqITWl6Sk1YiEOzgiJweDWG08Wuh31EFcdsZ+nXU0nd/mTYAEliPzKTBB1M
yPxk/7Z72G9ZOt/9bO5PUA2V+je3G5Il5BG41v0WZP9NagZS7ZrMdSzdhpTS
1Oy1gAnJZWBsG3qxLCE3R7LsYYu17kEhqMZWaT+Osvdut7uUMVjQq64sScFN
LtbEVA0z6DJvEi5T2M7j2WrTFs7Okn59wKA8ncXi4IPXh7m5tcx6Zj4faEmF
K9IGS/Zuq4IGWd7AZt+LEEp0VeVvqwn9+PX9yJz3aCTZsHyy9MnLE5BGJhvW
wG3t1b7VhvOYlcId2yGQfBUbKt+a3i+K5Gj4NmbrJTm50DAXx4mdMrtm6BoS
ehpZ1L25Kh9EvD8fgNuPyNCkiUrHPp1YSjbKOTkqyHYZ6hqJLNbxsHbPLcYM
TURQEnKVNsaBZIhIPUa+5v/cTlSV72x+SflwijkC+6OzYDBnOmprAeP4i58q
VeXk5v8lLogsztMuzLqm2a6SZ/I6p0q1fzzVcBK2FwzlTpFw3AMUmk5LA4uU
u4gsca4fXixk7+xdn5rARrg8iVdndhek0FTNAzsnR49mcw/fouuJX2Ms1rnD
JVIkeC4suoRQm3Pkje4HKK/h3BAdEVIAOd4abdgQldjiRzGJpvkJ3X1ZDg7I
ABYxvx1ivZHMNPctqDAUIt9tyl31QFJx0jKkFK4nGgXBirX+DJ2fdlOkG0gJ
pebiRTsf9qqiSPYl1yAsj/HRocY/UYF+QUwIT6Y0Gv0elHpxZ0v9TFLLpySY
89v1qNfFiNC35H7z3rGQsH2d1UJxATj3CXC7c5yaveDCfoC7B0ht4rLJS6R9
hhj4bh0nwViqPi/03nDHuBf2AhJAf03PcDTyj3g5YaC+FsqcHbFp+RFvos/Y
nPKMiL7/r1wW0CMRL7SZImcj9FJVs4qGlRZZ4Ci/2syz7Vvcusdg2Vznb6ii
ykiUY0ej8SX3r5g0eHjQgYutI2BmL4URVBoZLighHDKSWda6PbpTKKsG1Lo2
Kk17+sMUq6C79TtHhsVeCRAckrdxv6yW/Gk++ktXB5+pabqhxvS5kwG4nRyi
L8BTBrluJFHjMDfBPX9h6l6vKSsi1MSIXPa0uAfCT5mutu9fPX3ECRTZ+E/K
VsWr60PXCDHV4YSD+/3bcq8Vir5LoHShSgxhRNgqsjklNmnRFsBw9C8/iAW6
hxATcTdzQeXIi0FfaX4Xa027Ybx2CuA+zGc5YS1cs6McsNAEUTKPEjoEznSd
DwR59n8TguyAnSXGpQIAMKGZxFvbq/caSbtGKoatAGsZYITucpHt9SkqjpJl
OsYXk9k/u+BJJIm2PdcP50aXu2/zOzNtYfT4fDCG1J7Ch66uLmPhDnAzczjI
UZTyObFX6Tyx+Vcjl+j2GLPVMGafiPXnw4vtEmtp/sJlV6GrfPCNOMWS4rh4
d3y1UMYux0Ji9GUORNKq0H5rjxAKA6zTovBY4LPqgOoDT01sLPWDbWyu5N0+
p+ZbikqJLwXPTkltyfqnnANG98CPNVyGqeSJrv7w+yg5sT8P9l4sOvcsOEeR
CN7L378AoRptDIquhi/cd7hT0u+zhpOchUfdqJHdM65UpY9WEZ6Q0/QokhjH
ZESAGipuYnkk1PsrCMT7RvMaKT9RoscpxEpepm+anCxOgcr20ezHOvC0rjV1
bNNlBlAlmFKQIBORvHOmXm2SR+9MG2r23i+iuaY7N0UmL0TvjfgJ8g68psbu
r298DSKFku8dqcggBgdml/jcPib3cPkl6p4Y/Bh8b3x/lvkpXwP6plA3/bnC
m0sWb+nUK5kxbm91nJlSaH6cBiH4zzuQiLrrcbciFMi9TKbDSIRfEDRXHUAs
B4/llpfLTlion2A7havsNopJwxL8Y/2TWUcTY6Uhk5yrLZfJaqTv7qjSyc7j
z1q3WZvtveHSQY7+up/Bh0HgGDMh10ZXj1TLn+c7EmZ8grfga+IgvyclFehB
+WdSWRbYuw4QrEtyEUVv5hRRQ1SKxOa15PSrFhbYBOjpUq/IudihE/QHN3Ab
l/bHoH28h4g04iC6njAa5hF/g5cQl16NJqR3LPScCggRlVtwnPXeaF2eshON
k55CBiaa21d3yjRCE/ePa9tqqaeUhofk/bvJRzYv5K6ddGIiklKiJeo4+Sv9
L29m+2z+YXGr1tANI25VhH9DylWvxGHa7SJGeDGQdpgW/RbDAIIHgo5ZqpNU
D+ZDK4I1kpl4mJIqazxQNkGji7ODicw5OWrVydtcxNGZZ+5j+Z1mOp0hSpwU
ffeLCMBzL3MYOKi3v4SEXdrLKWDT3T7Et6iiNnwb7/zNfjyX3g7z8q9Y9P6A
w30hrh+6epoLlIma+d/lzoExJ3uWE91EDWnr2WGyWjClGLq7XYq4M4a9HRXp
rNWXveDvrmYJpe4US4GKjbGMPg3RauyVk3WikTaoRLRJ8oWxFoWfPhrpzS2B
H6PKKI0/c1zhzXm3o6eTec8MxitNI0e/UKCA90Pfmbs86LIxfmZcZZ7cvJ1D
gYTbZPeOSaXZWU3XTvRzuHr6Mz03uopGdyrH/uySUuPpvmBojBZ//qGOCr9O
9sWpi3VXTPiXcVbUeWrh0ynx0OnnsrwmvLHKuupZGoUwT87tlR6T37PB2pRx
pWTWXqBXbh7GnErrq7pIvvYRFeoxJGPxU1+Ras5Ot0mfjY811jpfa+ll2EXl
FsG+tYK6+XdAiwa9gbRL911CYgyVIKlwQmkHuNyopK7OGUgtfgMvoILKF9ME
Bdacw8kNOo96J9CLxm96LH8euxErjqm7A/yVEAC6XdQ/JqJp7LbphD/SB+7y
/3iCG3GPdmo4rP8i6EWIFsMSxUAShZ6aR8e4f2CVckIgO38QCdoYJZ69B6HT
ONZfnO7cAZ9WHK2gdCFwxhqu8iIajQ8RUCmK2rQ7iNWjPAGUtTB1mP3j4aSk
NgRaes8/MXn9Q3/V3tomiR7/J//8gUyUeaUX3V0BK6NPaXtW5dU1NA1MDNhA
cX5xY2jDlijquVurA3dnhsj86rBoxWrbfnmedoYXNiz4Or18V5AGmazWZT0h
ty5Ch4iNR5XUpc64kBknzHDz+dAiNltRGzwnWqg0s5ofupuxUcuMZWNXYoPS
Y7n27Nuy25dCxyD/4fE5xoY5UAPdE1CM+yQ44MxQ4OVkIK9RPOeO+RO5INZC
Qiq4+e3QEKL0sd5SWUowSD7RRZhGlTfKrtqtUtLsxTlVNiyazu9uOsKCI/dP
gT59Tv6cGOz7UJGlnZNYfqnjjXmWAXAwZPANSPSgX/j3rxD2Oz/SV9SrVg0m
6gLAiTtJewb6iICP5E/nMaVlxDxTLO9jRCQyyGJC87CKykUqugrhSz2E27C5
lXePu0qje3FUK/Y3k0zr7hpi/gRbMoyUvl4TChkNd34fevMkyArSuoZQE06R
L66IPcqcn1GOE+gPCevFWPqgmlgUZVAyDrBfz4kBMWlxcdTaiTsfdQDg5Vrd
pQac21d4nBiUO1E0yWXXPTTEJHv719pBRlvVmfw3Qo2P+mESf6m6xjZt0k7E
pJ6kUWjqzz7TTm1Nxb6kqojtjICv309hWGrMuwhgk92zrPZlzDo9rypDezfg
m56pybL9xA8iSpJY87duIsC0DvMbo7pYBRFbSKX5yzfN7mmHxfHq/V/CVfqU
+tmDxP9mU8mOMG3OqYgZaTTdY2FnhSNj/ZLjSR9DQL5VZMZe20hUp0GQWDuE
izayOey68R9I8q8fNTlG47NHB02YHOhkU/3BhowYKdsxJXpV2QztXQTSH1SW
FI3rVuEwmKZAxRb7xWbbdWLQ0BHJoPLcrNa0CEQHySdj0pN0l0APLahjkqjW
ziY8nKcdDIboukKPiIi/DhdAOLJqR6ElkzzudkF0WV9X6ME4izkBpgHOxCXm
pPoaJFzBS0lKBdydTvfIOC01KwaLOShN+PHj/ipqklqJyoS33h96fqqWtDqE
tCcFIFpDPPjvC9ChkqC1mPMsvOMXwVj1MyNeVDb6g7PkEKWjO+smHZYL2UbV
1ovm37nR8g5tcJnWTvae4pYMpwBPnltHwNRyki2TN7jDnsUzTYssZziyFGyu
FVkbYl5VPeC+nfqxVYXLTdg0rb+mvDR5SMSv6XcxDYyQ0JfQJe2pPU2UwBSD
zxD6s/eRtrYpQipqlcHJXLAkeKBBqqZXVn8BejhhAASIDm9Z0tNT8pbdPRZj
qY2Yd6l42TX4VKcgJMmDg5tXh7qietam0kIfuyMPxoGi1g4SP1V/hQWbZlRh
BFY4MVzWLQ/PH7PaSGCXPBsqp66wdxTZw+1l3G33Ue3nYrcJqj5uh7l0UIfC
9R+a3AznNhou+e5ti1MZ6vyIlAJqbLcgnoNhdgmIrdlN2GtHn0skSxk3eFhK
MW9hTGh2+LtC5MUy6cKEg9BdDiqQQj6NBEoG7u+YH2+ohdQ3ZxRmDKOkeVk6
BsIKHsD2XjKAkzVIvpy8M6NnpxIJTiSPC8ch9nHeECWjJJBB/HIU0hXY5c/S
j1zeHbqSUV2mbUVK4cQkGrbZibP9UuI1wV3JdbJZONpFTbI4Eoi5LEwjrJXy
Etp1QfmozVZPyKSPV3JljaCaZwq7tEW/zinic47Xjdv+iCVVAlt0iQ8wOaZ5
2qWGSSH9VyJ/5d0JYf/FtDz2cLm3MvasJ2+3EnEx0jIiQVwcLgyk+XiEtlMi
+rmJajgh+Xqb4Zbo3RHKbCvxTfBq2QwJXInHD91OfXYWKzbrMKnugseTNtMj
gdoGaSojkcUxudyk3OwC8erNtM0HTv7uhtjlIE6YjKkbM28qnvEziueVisoT
dcZHMY2m/sy1ahRSMkCz3bU/3u1tIM+FU8sV8NtaR4zdIsGLJNLHyoIDEA2F
VEfqVpOFyKc5xOEq39ljDOWm1okDDESKV5JKEtVhmyjkkPeBV+MuW7FvNaNg
tpVW8/kkIZHr36imc+Q0PfJZn3wIDt0QkZr2cko+sIoTflKbWubnK6O59jjj
iSSaJhxcEp8EFP6Wa5hESR/uw5EHnTfby5D2aSq3XUAU12vC2+kuwF6FelXU
cl9tFIHfyurzhIVfh0m3256qYLcziDKxyJp9ecMEk+uORez6j1mLZragLeec
sVzXXbrnnvbqivEOCFxylMfToOg3yA8IzBH6kTY9cPq2UTPVUYXEoajDFaBc
S4vL6rgyTq7jld0gC56G63AsDM5mgI+p+M3vlvCVUXZtbByEiBFDjSgzInVR
Y9Fk0Mqjr6TNvcinVzRuTvBkxsCAPlGEqS/8MHYlKT5PdxphQGvmOoQ3KUoa
kb9dWRO9fGhIpptsk4wilcTZNeF79V5YNfcSJAc4ickouSKSa2X6om5aGnwo
E7fLsrIJJOW8EEPrxHt26DG1niK8gJOtRO1HSZS291+NqVl8GEHvSLSXvBpu
9HDH4p4MITOzTizydingbyLjeUInsF1wLw/HGmzS0Esio4AY2B5AM3ysF8iY
RQz9KRU3thRGBaX6g0puWR2BPXw58I/UMdmPbVUGzXWDSbcvO7QeZMx3Huvc
niWDsQgK8xiRfggbx066i7+qmXvNB0SlWUOdsJpxkkyer6xecWWVuLbusIoo
tMdFU9OQNbNnYlV7RCHqsXW3IXdDXfY4kXq+So88wN+AbEMqXZcQ1uV0IoxR
hUdcYIxg4547pD/9NIAOvMjimh4DzkRqPr0xgE5D7z4kytLiZEaf5tWAZPL1
ESuYRrLB+79ArgS0qx2Oz6If1Prxi+3Hqjmam9NJaBMK48gyiqPnRMyCsatt
VB73YfJ5qBWBJRkooY5zJ8RpgFAke6/xNoaBpX4QrG1FyluCAg7/T7dgYLA/
KWNFkfhPMeou0Enb/58JVntdHn4x46mTjOQkNQMjkFFa1uoQ2sgzs2oDZpJA
VtWJIki1lLX2hayV0+V9Co/ujz2bjEVECeCr3/MQj3+LKIWgkCjGxiZe/QQ5
12UR2Jf684b3DILnGha34TpTXmd5u5+sLgGxDGG7ljhlFb5K+72W/GdebOQq
G/nPrnow0daLOs1wBrOsfKVeAF7ks7/iVz4cV5BL6EVFbEQSgFgN8QAW0qaO
NMBJxT4NKLVUgixXFF10tXqTenZ4K/y5aC22+01NAbNTNSzMwjloC2t4IQt2
kRQq8qc47GYdXHXib68O4U5GdaU6LPUz3rh+dCGTYjm07pyXn3daWTo9+kGN
cTdCUM/W/m2WT76U+mpllOb1L+bqM6RwC7N7mF77u3dr0Y+99Q05tJMmFWL7
uopVvkEGAmbwYT3OUI6Ms8lLvqyN9laZL6EzgDsq+tcfBCi+KlrSUEMgiwnS
aBaySbiPnqhGNjho2PIkyFMITnlVUNmAydFCR3hQrzQGBrHecsCONlf6DZkJ
FozyyHGMiyjlyn429VFFe02vGYGTBIxr7yanXTAv+iIiuKj/rgEkwocg1nQF
xxgA6ioeYrqAkczvkQkgIXT+Yq6aKDk3+YRjabkwGbbob/xPR0gHTqrRf5A8
TzFXPF2KwSTVZ+3ykhv9jkSU5NnBCZ1gs/11Nb2ZwdFLP9zezPkVbQ5S+pF6
I9I+LJXewegWwZuisbMKj8GrxORpAzDtnAHrJ4bElWm2gaCpkKW2NJdDCbi/
k4nEwJ/0UnMEtCzGzhRA0kLKqv+Q0BvI/CuzayRU9nwthattlrEI5n70lDt3
H3q7SlS8n/VBpK07DxSqv0sD7Wo6XKgYkJLypEEj6KnQIklqzeLwuokwcrpq
dlcsiG8IwQFNOo4p8vqUntjRJEFmt5DKYXWkNN+enuja2ZGrDK816LdV8FrB
So8kP1k6Uix/3k4Gfm8BtOVVuLmy7Mr3QOPXYlcC2OCT0VUTnMp/K7ee2l4G
xgNpmBKrTA7Sqx1t8n5xruKAatGb1BQgnOHDAyOPbrvbWQ+0OQLjczAuj34R
Hi1HX+toBmLRshZbIc9YiiyGgvE0BOM7LCOe5vfzMZm1E2HFJulSK41CGgF3
BISG1Hj45z/4kBe34oAIItGoQfPoBO4i2P31Telw61PeVN6nKOivkpbyedN+
TKhGxNCraw6g7TIe/GhO8ZW27/cfO6q1RTbTWExXHUh3tIABG4IQqOlx8MXA
gFXMshtgd7ojalS3nneAf9EHuu3CYP4UbTkBli9dPRqWnx8irb2bQom7a6Jv
TSHpn7IGXqm8Us3JpJdmHUqmI39H9s2rK5nEJiCNp/EkN9hXmQtvgS+/lgrg
f3QYdCV3hJOTfv9Jun1l9aNGOG8/LIYMF7qVK4aJ3ahUDKYw6iTHzqBXgaT9
CDYX1+YzHIA/Rufh40Ymi91q3lbjVU04dFByRNeWaUvfC1JfBxRnNeIFiITs
lq/CFcaZpN1cQaiOus5gQ2y9RxS4gfMMDMgQcA12perfeyMD0rgv/doaeGrZ
MfuSerubIe0Ck0PrcGD/KWcaZXWKxBMjzRudloXsdQyW9WR/N4B0RqAcIcrf
EmmZxgdUQ0uKF4b8FpaNUmbZdWiu1WXjOZw2wChcywLGhmZHhUPeMFJNS2nD
DQNMkGnqoBWUwOoazMNNCLdhB5t+/R2O7EVU1fget8MPxdZc57BxYLKL7oU9
gpLpfxFH/ZCd68p2ov9WmgTR4qBMx3XruiOdtgDOH3s4QTHaLsy1mtb+6a8T
9RrzdXt/CCe/k1nF+wZzNHZ/bU327h+YQkzcyeFThnC5+3YrCkVQxNKPLZlK
7zYglwARYs4qynENLgCFus+RAIIhP9wmF/DOABcysPHDjE03mdBQ7JjxPFb9
ilLXUJWKtR31AUS8YA3JNo2J02fsFFFldxGFQpH5TbVqPi1JvUblLhvN55Ds
6xhkscA5Oj9FxPjZcRzz2bPGPkVaLxsxMcs0tjIxX1hIUZXGvMscsh0XDv7m
89rrAoFQoSia+mYiSywEZLCSStFAl1Rn1zzaPHurh6y7loyifugItfd/gM8c
ESk0YORC9btyBA8gBktp+s/X7b/anEdTfM4GL+M1JUHl8JVDxRBAR/bGNqz2
Y0VinhepyQwxKE1y91UpfKRrv2CkpdCDdvY30wRzFwne5TP+Mw6nnjQBtvqQ
+k6nO8ukxtgFDvNpURbhT/6v/n/zP3PuGfShU7RRNg6vbkYQCUHL4juP+sY9
eL42yR9iLBxRo5PKyGlNdiLUGNCIttBZiJpNBI5ovhxUdR7M63L8RIuWJiMN
z33HRtrZhbjEP1vghgWJ/T6zZyKrJ2pdguHPMJwnawuczFOrmXT8D9NjDfrg
eQVvvx+ZKYvbjTBStNYhjqWgL+5FoRMiZfG7xgb3lnhphHXmigs1WGOEaby9
CbXFS4Ny8otb/J4fxmWxHPuMyl1vbvSY07I67JKNS3AEwIooShHUZEwGggNx
rNR5IPb8Tkt/shqEs0XbdbOpOCQIBrR55uUcH/bzSN5ydVyiW7vL5yXAcTS6
FUCzzVCweiJf5tp9k9wZA3yXtmqw+kes5Bk/hjnXl4KkhESD2Nak+4lcOAAl
M7txBQVrsHSuCUCt/a46YuYm9l+tOc0c6YA06YjhzenjonBcvYVcrCl+7j8i
/SkyIWSmlC7o0gvxLeN9EeuhkCyDhoGGOrUVTa4Vx5mBxd0xB00IeLoPXDXU
S3LMSmenTj/9R4xO1Vs403+azTDzG1rQ4lEylzeKJEXUD0k6mbpZ6MepO7JY
bcLgzwt8CCIcYZXfNdLhgzfSSqJqPp2GlQ0t0c3KwjqKHYtJ7QAOuzHEv0Os
D+q7sxJ0InH/49M1uBxsW8nsVs1sNzjXaKyUG7dZJjpgKdkldxEFiu0D+QgG
+gFP8vO+SFRZ35yZ2CR91cIrq2/uxo86zUEEZ3yTeSPvryxiLAAvJEW5Nq0f
ryghxVLOOY3ykY0JnPNzMV0eBisROTEiwIENCT3YLRwQZh7enpqvb6+hXUyF
X/XdPcbeZkDS9x0nrxfIdr0JVrJiosuYXNFIw8BKLn+13zweuR4rruJ+mIXr
C+4WKvOX0ZP9s0pXMSVmQu3Eq/F6xDeaMsoO5BhP3gE2SgcQ78Y8rGfZh7PT
jemJpcjFdQTZ8stJw/LCBEa2qcHvycdDr+6Wnr4Z/iKDaZpD6IEih4RUfrvB
iNVpQ7Ze8kFXcPNoRPhlCNtoGJMt1KmideNOjgsr98T/l4YOa/Lg04I/BqeR
ZWBQnFbKivelat3wA7Ww2woFvuPFasCXcXvIypZgqX/3OQ93hGT7eOibbEas
0E+oCa6UREFLpM5X3CJ+51o+pUUggTzqrs8fDlvkrdsiX/FJJib2S3PGd1m1
frmctuSmRhtKN0uFusYRsiWsvRQC3yzDD05Tqn+cL0T3sgnFHBNdsWaE9lg4
mMsBeP7G6hLzN4PFFtGf1jlQbRn88jwjHFcXyMHX2Vhm6t+J5qpPSghjXZDe
0UJcxp9BbRRoCvNPQ/zuTOh1SjQsqvdhCg/YG+39AzLcI/XnY5AgmZzj1I1/
2eQ5uGjbKhe3hrenpbTE/5WVuUHHD3ETbublgXTA10LFvGwFinf/YBB5EqyS
bbtHWI5HNVoRZyMcFOfnEyDs6itvWkamHx8oBNbWw/56P8D2O1LPryZPybg8
iNOrLmK4brjpCwCzYigJN9lIECMua2fR5PZLj3w6IXci+iE+YIZvkub9evR+
2UNAi/60iVTphw/wih2vM4I4VLK1Fm7MBMuYuyC+Bb+Y/DcbUstatRfnfW7B
NN557EnXAyNFJcOqfmRvrz0mOPxggMTj41SDV+wEQ8zc8ba3kPtT8SaGi8Mz
XOLYC9AoD12n05lUJMyoilKBpXOBu/nTyyy1X/rsat+7SW06W8uuxbFeHRB6
epp1z8P+zB4CIhdxcT2lgmmk6RdJ3h+vUOWLa98J+ZQAyTCtaqDqZRke+SYe
rg5JMqQKpBw67tsNpC4lv9KTm53VqoIYydiZk1gK7JSI3Wce55jbmbAtAJwn
ptRqmdV4PsnE5pPqXNOEmeSPnzXS9aGbqOgW5n3VJ5kg5quxJ17YiGCgfAuh
KTp3TlaMeWcF4tU/aGUxCzpNQGKhrByUORoEURijoSwboIBajJf8a/QfGtEG
gSGwsCnHx1yrYV+0XZAsibdq5EHS6A5emSVoZ/WVDcWAHasMyxtDBMUqkqa7
a2Ek7fj5XQ2G0Ec/l/mZCg+d2FxgLlxkUmvDDJJle433HTpRFHbGbn+r4l7T
wm6TyNppDHjMWI0OCSS6YjZyRHYpI10V145EeZt8jl8X8MhbX4xpGHFY3kWC
Y/0KWtR+ZlSN+X2sHveIx7dPNTF6XcXNboKbbo9hEKIlWf1g4FPhPBkTKp0d
OhfkO00UDftwm6hwZknFE/+yG0fYSnf79pmavWgzDJzKF2ge/uwfpgnE9bUf
aTYOjJL82HWlNtIxJFIQuSx27qjI7/Gw7ZohU64NWMIdlhWqLnB5qIAndGO0
xLBLRW78ckjbX9p6euZGSX4jeJkF7X6heuCEXNpGgHXf/n6RGO9qZrnST6mD
+Oe8JH9uuyr6+cCmX7b1jV1TiZm1cQlTDWzj8FjX0vYaxKmxao8bawNIifdw
hOBXSFrjXYsgXzSrprDTnrI1778uBHnGNd7WPvsAzL3Q+lbwlP9qXwAyLG9X
OqsyhIw5KBtE1+gJ7ytm59MXZ5RV0yHQc1aQnOziOAh6uQy4xaceBMjkjEBP
Eo+cb/qGSlw0TIsIepdow2Z/Gcwhm2W1DAt7MNAUD5y6rmcHovwjA2eoFh1z
ZYwrNyS4Po4wOQ52JgVc26DOlVsQU6HGHOsnYsMuOSg3Z8ZtngXxIUh2bx7b
qxWI8f/QfHgEtaOneblMkfT40ZGv6azYNzy/K0U77ebFbf7Lx/JKi/VW9FjW
Ep3Y6bClSuoteqoYPMt4GGngudGlTUjayURrLKFKCTPJepDziwL3s8nk+0LW
UqC0NP87N6d7O/yWG0ebKJZR572PvL7pOeFN/jXLzlL8WTcg2Gdq2Mfo7vmo
2NARDOrAtStIeX3E+pd2BFTLqVuFR35S31DvZMGLWLN0tBkDHIdQMUEi32Mb
Kv9PxL7uI1pemnp2mmJKeo6CYn4FkgWtQCG6q8qkgylmcdaORzYYlRm7u+Cm
1WIVVlR3T9x8lVLNUo3epaUjG3lZt1+SZdZalJUgB8fL95jhVlRAaVpmROuM
tnx+fKYO8aIg3juMfQuN8ckMRwAW/yJLH/I55g7R0inoXV5tFAketOrYPBit
j7Pnm1kA6ba/+cO++Yyu/HyR9T8za2m0HPGyPAwDcjfIdZ7bpIc3yf8NjoOW
crM6tWcgEpFDJNP9uzD4AVQZnZC4hyDo1Qrztxpy/eT/TDy/WVlu4ndwXrW0
5I/2Ti3Iby3UM0neXfXFOf8iZGSbyv5YU3KJIQocxmH1MWw2pxaoYryCI9kF
MFuPQ2s9ZTzu8hI6D4tjzqCmfVJ89rpD4xavFTBaLahYzRSU8P0m73BosORX
65wNlkqOHa1o0yQ/PoNabafU18QJmTOde1aDKOVIvo+viK2c8VHxqNGpXOer
m/3ecbzeHM55OXvW5jxW3INHMn75rmSXN6kpUBnSGiGnwfsUCCBOeVcnJvph
9hMMHciPKSNMjMfkGpJrqsna131DhI7iHIhlsdq4i1ULK5xcdJg0UAIxE1zu
0PHJHqqzI9L0XdnUIqkaEd+p6YUB7xS+77kwFZcdqcFdL1ck+doCsbYNexFx
fx31f015LbGqowJpHFfTTdNqwSaPbk8+6dTcAv7ukdmZBFfkCwyn95e+zpDP
JVKao3w7IsK124xSxz8r73+CqXbUNoyIgCjCfm/puIVex1fav+tZgTK/fz6W
QfKD4Pojy2LZjGx6pZaiFEokFsjrkXvadXL0TayK987ma3VzEEUrkX1JW9o1
Gnxtrn08/fpJ/xlnWgGTWBdKFwMsZYFcc3WhZ9+klgEBdDpKgAoDqsSpw0xt
OsiLgVQ/qYMPNWyBXsaKt7jBNusSg0J/ObW/pLn3yo1MVvjYNAfcqoyQJ+78
1zaU0rw/lTKk8j0bFF+X9glYgStI2tV1NuT84RsSFDYsxhbnXpkdlM8MZQq6
XSvX0GDtSDhbU4M0B6z7d4h4iRghnPUC0P5LTpEIEAw6SuBGyKdvaOsFpEYF
SDgWhGbPdADwd5y94z0sHvoZDKuN5X5k8BTcpgxiSdzsmvWVuL7OzlYa5IS7
Fn2tz3oxPen1yA/p8IBUbRG0SyNNR1l4WSey94ngPWn1KMfEfCS1G33Vj/uJ
4g9BulNUoVCl1caG8Le670IEfQhVZ9GK+ZGJvXlN2mPf92mMkUN/y2qllcAi
2DYATuRplGcdFCaYGyxYBRgyTGRZ7kdlOzIdzpP6izkz4VuJmGM+RI1+qERf
UfTbC/XdI8QM2fMBeyRYFsH2Q0yYmSlnBZWeNul4j3pNF4gEnS+Ec0Yei6vM
R11l+ULMO3Y8cbFjoHElc9qkMhA3MqL+bdOe6wNbswPSBudUIMRRJnpdS0Do
D+RytQ8YC5wFSZ1Pcnc9RXF7rXZMCLNQN4cUduC3GwkjABoV2A0wfA9hPQjN
sEifXDvzXWOHyoSg0h1oXVzlNcWxR25XsOe1RYb9GIel6BWyQDlsFDUNtqTj
7QOkBon+KwoZPDVLIs3Dry4Pbsiudsm8i+lzPwkancF+2FxqePoCberaIIDw
bI89Ww52zFeBndFWec9dmyn1hku9iRlc+wbAuMXxpB/ZYM5EkHG3K93F0Bco
YUglql24haMfIr+iwQWOzV1/zBkbheVAzDxAzvqYSaN18lP7qBu8tGcIzoSH
QZlmhoTefjjNYh6sV78t0+9fJzeMpRGnTphkK/UVhnmA/jQlzv7W+eG/IyqW
EaVtYgVoAMpH4sVuaF3f1TFz6aP8Ua2LwWGW2mYNle+faLXoP5COVX6LikOT
jAsg8jouLi+fS/Ds2uNO9ERDgYRoCEJWBYKbqE7mizQip0Vgo4+tmEuhjx8Q
6U7+Ra8+sZjbzEhMRNuS76XDVIBo7jwYOBuhk5Eui3NCxHnoja0feOR4un37
lsxrl5/QPIxT94xYE0cmCO7nYaeC557rXyZqkzWrHv261eF0E+907/G/vexL
QQT+p7mW7PhSFqxC1k6Pv/G8D5+dCQGBlOz4nT6Tx2Ju0QaasqdiGT+hEgVb
e24UlqSP2KIbAMRgxemlhsc+yyN0XKz8f9EAXonn44Gk5b5ja1Qmj4glJtOB
BGvzgYQZFAMuubW/1Hlibz+3Tx7jZ542c32M/pdqrKwnJZ7y7i1/NeIf8I9c
BsZL6avDh5bBA2HsVxsKpR0kpLXt4r2thBZXLGozFC7qSbFbmUQJ2ralnHNc
wzTQxnu4U+F54mIZx6sU2NTXRnaahWKKxYaqzD8DOxCbBiaeUqQF8mVOv2s3
/zHWFj65cwidva+ZPP/vhFcTqRtD0DJQaBs6hJKs4ySwxrgdjvav3v7I7wZX
8c6zdJF0qalXbf1KGaiZ/8oSGPn0ZycBLnWLceFKYjUH6r0agCYTSwz3HHrt
MWjfei4hyYNZm1h2E0UjGOD7OKty8y2qE6Mj86moQzirrSbaqwJpb4dz4LyU
5Y/qCUlw/ubia5tTLYydB8KLOcSEO2VK1THy0oyBK1VOreUpS+DQ/kH2jQYP
qCU3OdAHCr0CUlVBOJVhwhRJwa6fW9FDbOO/Amwubi4AbA9TMFdxvkMFBbLL
RqBdB3KrI0es+DTnCu7xf3/hbx6frhcPs2fvPsTPv+MDlyLvK5dYl8SmbKvR
YwGZr27CgBibhLf+767SeyvbyZQCqd4B0UaucJA1JLBTLOOzMhpRos1CUXsp
QDe8X4f2SdChmSyCpyPABSq5DWnyCMWT58GlQydUs/DEN/w6bzPhQh6fU6EF
ieZ50ABrIwup8KxWfGkcXKJyvufYdR3n5HHiuzpz0oKK39wJZ0ZL1g8ZkXRh
PJxGmnDIxfSJfFHj6WwaUr0wT+O76FFCIk1IzWUFV2fE4cQjW2DGSO/zOm1R
y1EblciCWFQzKfbpqSiJytWGtT1ka6J0+O8xKiiFA/0kdGm0OcMskTRR2eHz
JbeWd4m5y0dREFOC8TZ0dXN/1BYf+0+KoP5rSr6Ndyz25sFHIEAgJjvX+CUn
QHloT2ihDSEdY0SHbx2ronBoO3jdAuhKwLwDvrN5NrfQYtJO5s6DqFnxWyR7
5bF9UGPe5EpwW9jlIl9GOT86quB5VSzeDkVUy3DQQfz8DdiEotIK6wnp3Zxe
7RdKmims7KYx5E/COM0O5u4gk6Dya0Sy7DREcDI4F/p7SvyMy/ZwRMQYRjW+
52x2hv34N6zVEdFqsQ468mbCKkajZLImBft2XIjjBUdRZOrqzc5J0Oki15wN
L7u7yVtCcuw/8GMIi01fm0RUMaoyuCo/ekzuP3CyOWJZcfoGVYq0g0p1FiDU
EL00ZyidnxHHaY/9YuOX+VTqqmhr9rqZaLgQkddZvZXRKF4CrvmS3jHDdx25
FnAe1T1wfTpD413nq0cYoFtfG0EqBDRFShZ8HDPO1b+v7RctQiBadJxhhaFH
uO0qMYe0vcTreDJHMKNRv8bprZR7fbYyjJpHzudk2r6+WGcgO97cHfAgRjRh
zpaab7Lecs51AE+/behQwFC7+7y4hRyPyQdaV1mn0nr7tobrVF7jqYMgQbMd
cR40nr9Syg7A3eA9yTyUBFVdBTUt2RBBPbWYIUeRx36HSfsITr+sCEruJXf2
n194JJ/3HwA0jtmTrx986Uo8ST8gjnyxg00mUKJ8WlcTL9kglGi4SvCi8iw6
/h6BENi+uktMP3MVBsJ329Xx1933QFnodquXwpw1pa77RAC3pgZn8R3majzd
an+jqbObonB8//NCqTtGyLbb9A6PMQoa6fekM62QIp/7Fy9CU4sQl/zkY0yp
VQSosiMW6aNtU4lOydBMqPzIix/7k8jNdsVFlFmWI8m5fonGuAokTdUK9Mw3
raCSHS4PaLlFmk3wHP7yYYvLdw0is8D79Zz8EjIAMYmJRABwqFvAuGfxsbBl
O9M+QIVczCXZ52t+ziNzThYPxNR/Bo73OFLhPdGLYJQ5ApVUvJAOQdgLwNZ/
5DDxJp0hPm+rQFe5Wv7/1P8qJuac11zTrE2x4Y2Qcyfx3H+Rk8lssU5Rw9K7
U+lDnfHEcRvZY0DMueIyWynfKFxgrUo6MSB19TF5LFb8qqkB3nCNyNqlBjLt
KCfi/Bc8msMHTX0DwZJrP2WAAymt/JqJzju8B6PZxzU+4hI189a0s8XD2V6h
GL/t7q1u7e4Ny5gXA4AOgRvDngwQyuXyLuBwur5XqxAYBd/jEIq+OmKA2dXr
qyhUGEyckGvleYIBuocx9hycSPNqxpuVhDmM7SgNpKztTqRfw/CjueKJ2Son
SQCtLgR9ZMLj6G9H2YkQxw7y4/IkwvR5HJwhcykZX1EKvnJbXVF5sMefAFbq
kS9uhm+wumcnodjBPeYimVnXPPnkDtXM3u5ERdIKlEisHQT78njoCiga9Qgc
5u1MuBq0eNCtJZZdFfiK8pM9IKfi9iDM/WEd7BfN6TE6TGSHz7IjucxY122M
g8K5be9gz14/dt/PEdTq0vaCOS51rB3RcxxNnp+e/GTFTkWshjZxNaHD+77u
dz/Y70VrYnlMQJcV0Jjzn+V2jG+E45TQJ+BH0EXYZ9y2ju82J5HjHF97YnQr
5n0czh31u+0MByRFP4V7smfw9AYz9/hosLM5t9pbUuauOju4R13CPbmu/YtZ
tKvHK4wNFeiT/rsNDsWatYe17SHOIYFwj6sjuUT4qQIz+jwZLcjpAQsel0TM
6u9R1pwfyeS5DwTEipiMITaXACy+yZumsUMAv4OH5oOepYVwT57I+JE/R/Xm
l4PTUYiAkNk2TEwMd02nq+NDJ3XmdJihzo27vgIC+Zf2tH52f0kF7sxxk2Ra
Nf5wVe1gDr42IKYGh0x4KDZpwfahxF937Kun1EysaVzT0v3783dxXolxT/iw
HkOqV8gBvhBcS344HHuJRO589ja9ijqwcsWi1WiOihdTgAeEV+kT5Qsm3D/3
peJo8tMDE81Q0StB8unsC/cLsEk6XDuC1r9IuKpNuw7nHQKt3n6V8dQnwh5Z
HKM0RTvSdvVzzHh4P4iqENIjpeOvk5WhMgO629sDO36KpJzL5cGwEUqsPGss
eLnNbpNGIu8rf+ZcLVdNtRQdSyp0lcEDQnR09weizoOnOV8nb5qObOzNvgz7
acorQoeXCHnAD39CYQDZUajQTTeYsvXyoSTJvYhj20jdAP0JWCZMDpgGwJVz
cmyXnzg4hXWY2v9GhSTBitMNpRe2oTaK4VgBY4bJs64RB04SKN9A4olwuvLC
dc20UdQwDW78ECmaFf93/zVQY1TfIueQB3zVzb4GJ7b/nms+1sGUXdIazjq7
k4OO+HKOuTVJQbluIoyzO1XZMajRpPPN4mtlwggXxsgZQpWO6WOjls6nT9if
dlJwiybLUcnQ7ZZp1HaIOiFLHhpveRcby/bnNKgM6KKDoyMJ6jVimhLibRHV
qyGOvR1PGdItymG567zxmZcpTTJpT6gq0j/FjYOErPnwLRvcyL9XOVjWttvf
mxvE9ZkTXlXxoyxpbAj0smMxPuH3GBhwpWE2Xn60vJdQzJHhN2rXmHdqYjZm
uKtnmUIvn+mvYkRba+B8qcTLcJANguS9/SG6rz+zrFONQ/1BjQp79ZzekO98
xJpBK6qs/aRVLrNq2uxW3i0KiawPWfyJCeqbbWzPRR9rPAtLW3HR/gsdzMWu
LUHslxukX8UGbbrGcR89k2RoZzU0kqE7dFtDakOhe0ZzDwK5QYk3nB9/GpWG
N2edLSYHkZ/VzP8Lh58cveW9RHM1nFC+0sgbCOdiKucrOVl90xmCb+eYc3ds
2imRbs9PeVRfvw9/pfRLYRMoEPxl4uC+vRG2Us8LW3FFhheiIo1j65aqYPYE
2apAHxoXD6KDZFmpDjY+mCmuaVsQSUqRBT5mGFO5pYStFOb7OXKkLalijmGx
jfPU24qdnnRP5i/4I01kn87f8finag5vFcXX7Ro8FRysi3vfwJSRZi7pOI4E
Dy4a5gYZyFb4E+53Co9E/Rg38+QAqDVxGbyden0K6zVtOtKl1Kth6k11kp1K
z+ccSe2BqF1gpzfmbySG1ziMG378RzKGWfpMigO4XzT6MWjGcQXVKlbxlU85
yreCMDl6NIfpjZuJG4NxvEl6jzF85XBwBdRRJ9HPxUM4F8LlK2qKLUjdGSn5
pEznL75rNvIAyBu/O98dckWte+dqrKHc+PplUQzpzhNN+W9o0DAc9+AMmMkH
EReEM5Vjx2jK925GklIFL1XT0ZGXEYl0zWBH/mi4WCZZnDlka52qb4NF4CFc
DLaS/MyWMsN7vuaBV8FOiWQnvOkjFK52XXjjIcaVCCMwfDA2SHa6ALXEJmJJ
XyqLFIMJw7H7IE9WooY+9uToyv2ucNMb9G87KhYcoF1MEKr0lIf3c4KqKfBx
CnfP0/8YYCVUVFdtXM4gTYm+q4mgio3YsWCIi+wRJZSOZkfg0byPm4intBxM
M9WCAiRtUCIre6oZEPr6NEGbSWEcgUEQczRvRpWeGWOXhSC8akWF++d/xL5J
0kM8x7RXmfKQa4wYaL1pk1PiXdyxf/FmLDF9G68oumckTI/dEodCTA0lnn3q
LSYmrzdU1Jmek8RZgM6YN0XcoiffY8hyLzuRSrtE/9EwiOk/EX8V8culbpMs
rdgxlxnBaRWbojFsHlbnxRIuQ9kBPoBV+2EHhxhnwq5TMAvJ3eYBOHW8caKk
jZNY7c25r1Z9wx07PxaoZVdwgkOCw8gb+YOQ6I/sR16xejbuzMDsL81LOBkN
5kcljhLfmkoey71AUxT0kuLLbJ9deZuIl8piyI5ca0xnfK1d7c+f0R2MZ3Ad
0Hr6uSh5jsZLYYEADEJhp6PQ6X3RpT7qugbrFwRYBeBHd2vFd/IZaaYHM8L+
qorfLC8yg3ksdnJsno+rHJyG7qX1625UX7tYUi7Q3AqZMw8VX0XAnMiXiEtH
P/e8mAtLatyfZCxuDfUHxb74xzY+kKIaAzwFKliUH21oISE3JLGW78U3dlKs
wYpMpytHX2TTtzEMfvsWR7CfaONU4jEerNlfadU3kuL5K7UqwBexu0LDXhrH
3QwUaFg6jIfmzUG/8dfEyO25Ydci9mBHVnc+t0pxteJfan7VKxAsbB7lsUzc
9RsTyS+RDl0FPbuAf7Ib0VOBEkwP7evqI5CcokEyJZgA+w3E1HSWgNBLxYzT
qC6ps/v6IhTBQAG1hWDM9n6fgmDYLIHSKMYuGYpqHryq2FRbOqim7OPcjM3A
aKx+DgEUn+NF0iG2QqWbsFmLuznaUZb/Hk8FrbOLZz19tAhK2fLsjjhHeVcY
/IEGrDdD7Z0wKJvRn2G44/Su4vU2toTBAXKtxGYf86AXhap2trb09XUYQOvr
6q0n5KSN8SoPFyMGhAwPT6LOoe6s9WL4QAhuki7mL8bBm0fFODIzLzVK9s6o
a8najUstAsXqfJkOnYe03Ez7pPlEXrGOTc2fOS6DJFKPO39KHXgrNWr+h++F
mt4WgKkCgjbWzviWbxIoIY38c5CuAVLrRFgMwIA7L+/byatZcGAAQPYD1xnn
uDN4uSfikEzF8lZu9D7LGpgR0iC7J4dkV0M4vC7QnbnPshgK4QEW5AFcKBns
XGfoVVp3n3A/bqYFt28Rwddq/WgRUBoILNlB7j5QxhewPD6XtD+3Cx1HXL+c
weDfaPVbE+cRgBNyV5ym3pBtW02m4tOCBarLVTKi7oiRp/tpm5aF2gRrP9EF
WOrPNdi9DDEdRZx+Ue0+i8TBjF7tWRpCGt8Cb2zowZuFieB7TvsugHCWp57Y
QiRaMynmsaTZbSkMhhMQ5I8dsyizy+Ev8lKsDrOAH5jgNVKKRM6v8tvrbR/I
U78/BQhjV59T9v6ju3LfK93NiOQw9UEVjqcEvo5UNHqguf0YesbN0HroPbu0
pWHC8tpoVAHFgO8SNmDVTnUkYHs9TKI4jOyUflYeYxIcWg5A1CXUMTtzt4r+
K/GpxKCyF6owpTKVL79yvUIQbWxllX6WOToOpDKsRUutl8avBiLZi95wFEza
3qgCECfuSsAegOp0FFtGPG38Yq2riddea6KZe8samZdNRRaF18PzXE+0TSDn
YqDaVjajxQ3Omia8BSWqTc0+CifBFckiFbZw4rqCWHfakJSQepl6MKecKeQ2
Qo10wRC52f2RRGUTIt4ohqbibZiO/xbmq3iqiQh2RgS/Lujxxpqn2hqSKOg+
ZlS5zab6fn5SRS+TjfXyyXETG+aB7Kzrtj/QrjwaFYVC6PUf5T2BBF+skwnA
NGBlAcXvUiqiyGXiKWLck9ypq10YLzGo7aqLgXw4VICv5FQjwVn2vkdt/qVV
1KcYlJymxLLPcY69ZmNCABZM7HtDuoVx1yyBEYa27rQdhdBOWwS/Id52LM1V
CnZzbV+Bj0ion6yM8/SCbK29zgw1Sg8xA2cceR9EPw0O2v+5BJ2j5Y6s1VCu
mE9T8OOv/gYhPqg9EMlLL0+yrMCCNYZlrvqw60ggKaL67CUconVKPVS1mxuI
3Znj3WNC7yxut9gdy31b5ZyO10xSqmbUxmGzcqI4K14bPKHw+PFyYlaMRpsi
aNFLn6ooxc7hjRYeXYuSBtAB7CSxNtwncM0uKFL6sjrhDtYF9Wz3iM5Tl5NP
Q2z8PSb9+hTY0WVraeWZ/+/BoOgYLrPS3Y2UR0Jk/2WMMnYlPT2Lk3XO5hOf
KXCVuDkf1F/L4fTZqwCcWbkHw6xhAjv++cklZ5BFmwMCFOoIm4tInUl0kH/Z
oG5PLe+bqDHsF7XCnAc8AtW7EXwQ9TIgrk56EpfwjYHrWtMgLCXbR9gNk80q
achtZ+XwQ8j6aZZ8vFsSRLEApqUkmdSz5hS77aLzyJrhHNV1PbhGuAz4vdOY
wj+lcJsgLrTj1SS1GuO8przcBIAo9bnu8s42IPhLHTFN247bJeA3126Rt5F5
/mHWO5OMMH+Te5YlE/701Swrp83vTbJ4InK3ifQ2kQpI8qs9nBk6mOvYoMm9
s/gDiokj3pFwBRsBnGVTLjQ7YcPHAJcY/wkLH+4pVM9x+iH3/cfRhCyAGCZR
R38pRxNR121kpfUYCyJK5pNB5PKQLotJvtrJMub7Rhm2UyoNLvQHjJvPGUtx
tVRI55ht2aM0j3/uT1rLE2ZpIw3TGylZ8l6uHJ7DUljWDJ3d9OZbzkcTSzr/
qrU1vZ2uXMBZ/r3p0+3wI7IfNNHlObvQe8UFtOsPhhAadGO06HClVSPB25ww
FS463U6Ze3JMQzQ5wyySqU3orinr0YC8JqmaN6HoQFgekqx8TBHpqASeJQTC
h3Qrr2sUfIhr4eWw3c1dzRq1/v+KRqoB5XqtbdRPfhctIBhC+ZHoPCNGTKNd
YhG2OgAbU//nc44WhDt8iWbt6p/3wfzHMrNjN0dhGYfMWJ9MviQ1ZgHk2J/3
rEx9xrtfAd+sB6ATFxdOpzHQK/prLQ4dc0pUydTY6Kx7ZJ5H8POfjG47mlzk
BrHQTjy0xuaZhMmRzxKzSOlF311FKlBu9mKmA56NZtb8D2SgLa69UmxQo4/H
E2iw7BvxH88mbdf8NTuKbERim0RDGxr7hWO4B4tRwZm/+VgVajL9pflL0W+j
KMPyF6rwBnYOZJCvCmPb1w0swz5QJmX2HRFaDuyKuAIvABoaYHFGyuEnW/Hu
Zy7/EctrztNdwjkdskiS6NyNmk3QizHCp39HxU3Z+sTMowMxXZ3SK5fduBMX
VkEBVwo5E8I9nhNQV/qVJ30n1Kd3Oz6GPF57rjaCKhkFCrjXHHvDt9M0qsZk
qVcPhKYMFFcfJm5et/uvhQaNJk/YLpFNwiXLgDpfJuzvUNwzJMEm4qozc/Lj
aYDsspUU6IGf54RwPTulF8Mx1JNN9PIIrhxsNpyJQLB4gPHnUnVa2x3zPr3z
fvM6KQwD+XTyejib/ugoQFhXQwLFlbDR5TNZCO8feehCAq4K7LJx2YTjScmd
XLGWvm1nPAtfPsO/ZFYLa6oKG7qrbHc0EJSZGZA6VnH91IqYbTQxXoX9oJ20
Qo/Uldg5+P5kVJKlvcAyQJRO2PbEJDGH8OzSLJaClKSi+IL+HkTvabCiu+hq
f8wcS6tdPOmBnIbeD7bH1+Ut0UC2Vtod1QdOWBN0eacdIqBXMZT+vH8lOZV1
G8dy8WS+Kcuv67FcMUKLAi6wyhaba3TQatSBKu/fTQFh1MOH3JGnbz/d5JAb
KJCzqZGGcegou+YiX1iNQQZUeqH9pdWhqAYG7AtyI6wP6IqtHhq4F/+F5/+0
NbFBC8wNFV5CkfSEgfO1rbW0eQGlSKrsa7vwBXzaJxgBBEb6HOlvNYBXiXaw
8i9tviTByvzjNTH8Yx9S6YkJ859L4igBWMJsZj7ue1Aio7lxQrwr3JWCOl4a
DH/wqbuW6B5u3tzG8ImcBKvnqZ83UrbfE9KgRF+q6t6J1ULtfDg5ZXjaSiUI
ER1AgSOSpb41qpbr1xAAulpfxeZFvhCFZjPOQYBaUYTY3yPlQO7XDJUtLhPi
V057lCs/PmXAgfkKhBE8SDzWjh86tpV2IJlKo3qdzB5Gk5YC3rNKVP43pv2P
8Yeyjs7M+dvOFvgcbR72bV7Nj0mUW8A8SHOMny5nkJna5TEq9xWooreuQcD0
9IRsHL2ObydJHsYDzXhu2dfdNjnGOAWzdXKpjU0A1piGjYMLn7tcRfwh30eG
ugAP153FhhDl5OKggx9S7DgcFzyw9tgah/v2ukVDPgdz0+g+GLKBisRQYgpd
vS5T6F98gST8vYvYeyudtMStPsG6ZGLwFfWYHRPr1kkwxjwTCFD90IbkdYea
DGTBVCdwfsviGFHMk3hQl117To2oyRuNMAcLh8S5KksRpy7r3lHklfU4R3Pa
uJVReFFflfAT7ehgkfA9SSLxbZOuRCcq7jEro/kcmAjU22BajLwH1hk4CjU0
yOU2/r8DeIEXoMad1jpT4id0cL07uoE3DxnPVIrTiPLFeynOsucGl2rUBgpn
SggI28FWtSIQ5psZAsejDGHlCJTuPqzrd3aEAKLjzmqk2i7TtcmTjG9SUAiS
YqNniDtm2u2lWXhjKcfMVSPKKjahOulvIYlPulEkFmjs+c/GaoAKtyhh+90L
t7El/lX6tGbKieRH9Q3/6cwRUII6DEdBrfYtOKZcWp8+BDykEn9G9MFBtazJ
n2gODjXvNFx2nz2kKUgUjMuiSn2Vs1NqlJoVFQBSODNXzP0Ah6RG9Nh3Rz7s
XdOpXrouSZoWbGqEefIAFtvQet8T7sl1Yl2+Zji0DufiGUFT+qkvcxC/3V27
I3p/TzXEe4eoITwTYF7LkVmUFqMnPDvIrIzExp8/5E9kF8Z0xxUfyqrKHkjd
eGRkEBmDoDkXsC67ngPu7YJIq6hnFZLBJaCxKBZDh52YxbbKVj7HlCUsfIQk
uhkSH8+voxKtQMWNdLoMLPWq8VbZsfbA2TCqUuS3sQwIYnnLr5bSrwOH/1aJ
/9ic7P0PaWNfPwLS1UbCsYt+HUkDZ9hd5UWuytZZJhWG8058r5pnk8bTSnbW
KSmOBab9omNSE0U3ewiU0MCDFkqTzX1/KX23dqbvWXRBcImVxh9RUUh/21zg
TGWWsNpNNNPB3gWmY8ZFE8giYvyU0o92cY4Xoe7rFoVQ9uL083gpS1RMVrGG
jr8vaVfx8VjVONBTWqybfldnT6pYIjXI37TDkWAByK65wW493FAHeF5sh27s
IKYFrxjRPLm+//jdix2OLT5j3B47MzIFZCY53w1YN1Ko9o0nQt0wovq95jW4
Q6MNcFyQPjr7QJilzYk3ceZffl9rPyt6pNXW/NiQigYsILqUwGiskvx2DUL6
+Dv2Ll4mS61vrQQ7YJX2FOIPAYrUHBY8HhzOf4tisCs93Kw1QLnGg57kqEkW
Cl/JnMD1GNDbokAwY8vPN3ujnx3KqeLT1z4/ZszbskNC+REGh3n7snb6OFmD
X/QuyCGSp2adkCPq2I7Tlue7Z1nAm+0/LndZREiLMKCdWNx8/or0EvsQQX/a
9sCFVDGX1BjCxQijwZ6BtQU1Q2/zYD0W0bgHumE1AeB1V7iHQAuQ8BM0bul6
nf6eOISFhUT4X9pNaFjfZRGW3RYrbX30SdOScwi1EIbkgql0wt36u7RuRsq+
hj3Iz16UpOJMgL5Rh+oQvzdzjJTaYgf1LeNPYV5qGzWKfhc9xM+W6jqMgAbc
DnB5b45ZV+4yAAPKE0BL7wVIAsBGV06dwgcasArVHK9ZRb50RKwPv9ibXR1L
7Zo/FY/0BkqhSTiNu0vI1Ke36T8FujdEgom/86oi7P2bLQ2KyKdmJRxxE//n
1+rNdFpfRTmMTJiPUNpnRjlIEiW0fb0uauXaaQ8pd1yyG/mzPWFJIYvhXMDU
yu4q1OOK+fdUgt/rI8S54iM4xDdCO6C+MeKzv3I0zdPISBs24skK0esJDQ3c
l2YtyyyQyhWQIGK5RoCkuqPHim9CFeJHOYYKsGaM4BzLx+05XMzfy+OWVoP7
hA80elmdbjmGAYbwto1UChoLuiP9cHtz082/rgI4j/Qulg8y8ULCqWYRYTgX
OCiaSIEqOStMZQFG3v0yeU80+rwUx+8K1+FG+CNpL8h/2VmP4IdjZ9vLjeWr
0n5wEIL4DRnJIvC0Mnrnw9VX5uRVs3TrKFZTK569Cm8/K2/uNi5yNSvBMck/
rYV8TWr/2NNjpNYx2/gG1sqD/2E52IWJIvn/fzXuurYlISEP+ckLZxOCuO3G
M3ho9uGjOWQJBOsiuDtGEzK1YVBytGzgPLxIs4Ek6TuRfI1FS6/U24Ys21RI
dXSxsZISs7YzDBemZGm91hW8ZNWpa9Fihgu+X4o3IYUIg9ZnBJJPPzygtKIZ
QK1xgtZqyGcrS8ekKblBuXWb9icQoQNWGZ65UYHWJK4+xLmRADB5GzI57tRh
BmLDIYkjLQLxihOUF+pohTKCTEwtdW0gvkj2Ccjg2paO2w/ka9crAXV8fY+C
ed8RsMkEdlB43foVEEAeEkit+tpd/jFPJopE/5OlD2yFbBcUAnP0VchPQIcg
HiPYfI/2ZiC3EbZvlLAH58ZENK4mhL0YUGOP4VHP3MbsWbHhrWloBSIUDL+X
808y3pq4h6M4vRl134pbieGplMI8/OE6phgSXQKQ/TPBrAihMhxndzwgso5Y
Vv50t5aX5byUuVrhSuI0dV2PVgJkShvtgwk6rFnjL3WhSwoCfVxLQ/O6jE4t
ihdt1eGp1xbw3Z+hjLRx0FJi7SChlZINEKoTKYzT2n8VUG17UdY4lldv2bAM
vgmUxjgLPa8ar7iggIyRw+yzmt868uqezcxizVdu++jLt7HZ7kl//2pChRhO
BuDNjw/wbo3XaU2Sy3vZS4+kb4E+ViPAosSCXjNsnI+nXjQIAJeYcJCaZl4w
DZZaeWhTLaB7naX3iSuKoxvMg/exvlYmygCxWHie5CwRUNUbutecxei0eWGG
4QYc4MbOoSeSbc+wk35hNk77S7zdA13YOnfZ4PHYyyRtMcqUoRQy7C8FI4jv
XGkbQz+Shtmvtib8vDwLPGY+syJ4UINlo/sjgt6Hz34hbIXEgn2X3FE8uC2g
5bMpXs7Ab+ILtoEZ41QRM0QMCif3eoW0GYqWon7Pyn8BBvIUpjM6c7qYI8l5
yFrGid/CdKqUY3NG38jxTmAvWzBKKdIXSdn0erBFy6Nol5tA3CLOScwnSZqj
S3vrQYkYfeVipJJBUuEQReyRCNNcnrzWW9487PWCFA4ajkCdn1QrvsFWo3GK
BGyoftFcwt44G2hx7LcyMdQr0lQ/NlpHpnYEycWaMRteyM8K8F9vaawvHUT8
imgfPwoNunhyIlNyo3X0s+NhRaBS7X/eZOvASSchHcq/eWU3Bc1ftaOjfF7H
SqPKHXpRBn0xhtsVEzncMZLBoUNA3Zt6BmSpcmJtLwivmIdolozLqH+M7i8u
WrBbrrSMDMU/ZBTeb85WDgwZlu4h2PI+57geN4jKtMHeJz33TzOmQEn7KevX
I7/OIU7mhortyYozeWM/aWcSyZaRjes49Nr8tihxUcRM+VVZKLtpjrg9xmi2
Snj/pBNEAYv1+MKACkdq1q4lX886UgYQTrmwU1Hl8GLYFpqjbof56Zy4OMlP
g1h4e2UnPGd9R9xXwquTUryIys0yxhzHQwC9b/iaqoxt3iEmhWg73kzREoiz
KiAaRFUI9TAfqJtAsOq/3DAnBTZC9zH7Eusf9Ls/131YD9nZOwYzeCHsmNej
LnR2MjjQu45jokjXwvtcrb9KUva7FQg6ZBl5T1q/ozZCtPJYJFaIP3oheudw
tJQWhbUWdn29Odb0yebfTiKvlD9fOZ8Lqmp9sfwaic8JmKknsoXiP2Q06c4d
poJytlzMXMwWole1qjI7+ZqrtZF6N8tvN3YpOVKxVRLOz50BsGBYt7DtzSqR
rL1Ne1plgPeb6sWWJTngreIAvFAWIaCV1+dfYHm0C0X7dOTMws9DuPvoVTGW
+FNyK+hF0GsY8bTcb1I3rM1k9Cxykp3ixANYUj/mx8y6YGc2xgaVLKML8MNh
JgI/eVwTTo6ILpIgh0zgJ2pQIeuBm2vauk1JtKo97iklbF1g2UWDufycNo4f
sB6qqXiXH+kU0bh2F0T2J265aSaXXqor3tTKbROnR0msqrwRK+BVY52RMFLL
KtZrzsU55XDmlkvjU6rFT2kALoKDVrmOrRcOzaL81aWDiTQ6GMIMV03TsPI5
ft1S+bhZX68kGPXOuYf1Jes7yvK2g66THU1txEHilHqySySrsZNPq/n8NWA8
d0UwMGGu3XqSwkancPpd2CCJuiTMT7gnTD+4XQCEahiPJ0N1vi5h4hrVw5V6
Bc+Y2j1L8j9QIHv95WDnciTbg5Td10FlvvdEGn0W1+LeODDWfBoZrzqaTf5c
P9CIS5wd9ylwufdqtgEWDPmO8Paa8R/2weVm/BpoL6e9mErcweAv//H7x40k
/RUfYoBeGIP0LvgUrjkxcgp0zqARJ6WkT/3CNz7b6n+13sbQZZhSMMj138uK
qIYiKU0o+IHrIJfStIWw70DgQvc/iDNPdStF0q7wNRVtV/hE7ahtfADvf13h
V+6VTGn6C3gZFSIxLKnh6j7GtsQG+/c5oxohnHd8zXh83FF8a190EzAmGIoh
P1BNUJS8zsQAod5BSwQluVKWLDsYop/ut7MmYCAyO4DiGY0CSS+YFNQujhYD
1gasvLHZUUi+mZAHEPvxvpIwzY857bBzLRupC90P8L3Pi8zc+vhp5xSmEHP0
2tW4pp4xh/HUBQx3ZhwZKUd+T1O2b+/VtwZCRc1chmWd95HyUigE1qlwWDzY
/U7yEL8v8yoj8eprJfwiC0MEWuROitLRlvVKMwnG/xxfIcU15eo9XAbyp/zM
zrEHyPeUz+xiR+4K25/9f117jc5zsGRjQpeC0HCIYy3srIMhA51NJCkrskW7
4yzPUqnEKm46f+T8pFoo15O6i0rMNHZZNvRgPWpA7BTAL5cg/pXMtvvBLazV
0wequHZj3J/+nT8MHKRjaVMZnNWgcKDvYwfox52TcCAp9n7D9leqIStfOSuN
pSz7k3/a2p1/cfa1zTgYDYndVIVX3qjHF6BSvUKHVyxod6Ch4ACwyxBLqCOv
Ptf3KNt0BywxRdGQNkBLy8j4OT9IPBk0E3UlLFxaO7D6OCpwkizagrDjrs9f
exReCGp4LFwb4qK2HL94w8/kNHp65XjZz+KIMFK/8Y20w7lTzVJR7fRB3r8c
74jX7h+RoZLBn6yJCOmsYzUtJQdnCF1pQY61yg70qlnSskYhftpJ7EnsAw31
XNhPA52O7TMOTkdtd5k2vvWHSBhj06cGJIuRvoBJz1iiTTH44bswxIaF5udU
AZYcGOYybo843jgNZW3GySs8BkmGfnC+lHkqVpfGiGcbZm0IDHB/Jz91C25G
q5XzT+5Jn4Ct4Zy+b/Q398B+FHuF2rp1tUj9DQ1M3OOcLbj2b1d9Nm3eRuex
/G37Shy0MO6R7cjGGnQ92+19BW7bco0Hju4oC7VsHkkHyIUIhUt/+wSeocKr
ITfrE76AISMFF2CTFlt4ug4tS7MgdGWJS0gSDz7Wg14dR/9VTXcShiEAba4S
c02t9CuwDLzQu8kLYmpwuoEeXIN9MY2uJKr+Na9AAi6Q8GGLyahV/pg+n/cs
T1Xqn4JoNrHlRanCMZc/Cdr4UR7Rt/pl7fSMHpc+ox+Lx3YjJavaxMxEZH+3
Z6j7tCGH3+OA3wjtLTu7XJSNpvH3OE7dVquD5DYiHKMkBPzvEpajKWF/92Az
XcfmILLCMe6OaR5MSPqbPFl7ai06HnfDTq3g7BzFleP5ClOmURZkTWs8QM7K
i4NQts6VyaQPtxVs41TTihaYND+PP5odOmLqpw6agb7MkFiI1fL0lxNI3Mgj
NpYA8YC4M66St4R7yHmcCQFUJcRWn0jCcXFXPwjluaZPtFvbhLNblidjG65Y
jQyqL/qdn1yjdfh+Hz21BsG4+hNNF4tmR9HLDzaiLFUamvgmJvUkBMyVQ6AZ
4QIoDIHiZqV0hjYjwG0ggGkGmiV6HOtHiRW7JIB+s8x0bG5zxuWAZh6GBSEn
kvlYC9tMHwclht9E0a1iS+NLt00NIHpJdJ3GlPTRQ0gWL5zpQscDkcUsabHF
ZB83HRCpEc0wonHF5LKyugSx8YoBYKRr02rUAdHJe1nwsC88Gp0QlNcwmSLm
sS39JkrDD7s7LWwB1seFXz512K5Sj2yaDE0bbv/TyaBhqIZn4xmCYgv3SogJ
Js0OS7zYEjRGK0S1fw6EV8ZBocJUJ75hO9H3EjvV5dbPCvcWGl4XWzMzysPu
RUnIJ7M8iCXZ889CaSsc9T/90y7JjarrjNUImwl3XIbAtEZsUBo6h4EwIQhY
+yGoUQliobo+v/o69NEq/qKrdWap2J7y3TUxiT37DMRgGfaTVPN6muXpy0+1
CBvlnKGl9jXz4GicAbFwWN/xHVpHSAKsCYkrefj193WPzSRl+FFABQ5CMKKY
FwdY+MkSJkpTgfnwDehDTDWLBu237KtUJ295WOY18z/tDVc49ZQj3O/Dax45
lnfEKKOXb2GeB5wkrhBOEzn8H0RgtF7lWBkPwPzjk61BPRf4DJIdJZhJIzHc
x4q+Ae8MoUqiDFZRUdU6S/4o93lcSv7c6zx7LQ7z9AHJJlvkA0y2OzyH85zj
AVMnz/abuIjELYSSI5UfZBh1vPcb+TVFCn306xaAyDrPmmqmKaxgu+pytfNo
E88FvU+TQI7XBcytdoCWbMilspLOd0RL2Z1lmbmuTvF68yccj5UCC7RMzKAz
aG/cevRZN3riGAoYUhhf/gt6ti2633Y2AyGR/huIGjIANPy2cBkBnkYqOMdL
LDdkm/F7XE2ci5JsCF4d7DtdmuNZdFZwbkkliXuvu9M8SmyAWxOOhQK62GsG
QjP2R1TQn0T5LNMXdWnnBwAwrdJvoxitWOU6yURyAje6yt1KKkH34HZyUVd9
DWMTdKGEIwPcFOmui0jF1taPFJrKQdjwNKSsFtWjyDl7E4R22kNPhcZWsv9n
k0xApih5bw2NYQ7SpChkKXYu3Y6EM+bVn0A9bwUYq1/edDTD3e+8WZNUnXNc
ZAlBFhRYJO50qtGTPEWeXjjlIxq5KQ3oOVyjr5fNdknT3ttkjoaDPjxH6ygx
1VdJBg8JECSDGps4pxeBa42f1eeNb/tg5co3cdAxADIJP7bpBJUZM4JKNcGo
/35wvQI1ZETmSEfYDlR5lJUSm+w/EjWR1IA6VDCTG+Lsu9vCuF2G+9jzO9Gc
NiPGDwSFUapo6IGbbH1HJBBZxT2Px7yZyMzib2HpJvBKp/WxXtwwF6/yKZ16
F4WquC3kWrdITG/TBqxJcNuHu7cyExDTaylkdalhsdGJeUNWJ9LjjVyISFPO
gMXzEE8UXoVwbSn2SWWNPJGoDAJwkaLiEV8crM3ChABN1XOrnIPi6fjKx58L
On8w0n/6uVeBz7ng4AVHwzY2EnSQ2j7Fip7nxcScAJ23F/9Sdmr9qTrLfgpT
JsET1SP7Snrf9jUfxGnnHsEmC4JcYsjm0RSN4c9ScOy4kaDoYa4rvl4Bsler
/870FTGfNO1tEEz4uXcgN8SrbAmBrraFdzj6LMJfHpbJo7l9Rv/m2D5QynBx
dmno7QxYI8BmdJr491Sr4WtYyBZnxGjua6T6z4xVbsyoPbhmqKs5gw9Gd9K1
Vz2G9rSaC++X3eNR2KMn8oDXtFMR7Ay4aZktenTUwBlO7hFOC0PGPCefcN1V
LKZ1ULP8LgR7I2DrZxjn07MBawYz/PeVO/E+maDc+W9+kUrfS4nCOxVXwoqQ
AVOX8YZvjVMNbcdcx4EUsUK8Tkr2vnVZERxNAK5Xh0x6UnduZ5ip4AziU8uM
JgNF3JRowsggpbLYPM4QoCHyP8I1uYUl/tHx8K6+IYDT+jCmBL3GiQ8Tf81c
WSNFZuWHOFVNoGMChrIfmUPXtg/H7GGo57odAtBX09a4fHVxlpB1FMrvAdL7
se+HBUvMJrLHHA1lUFQ+xOcOGHwnxk3pxJi0koCy8nc0nH7441ojLxgfAOTs
Tljw2FgwfeRHLmOvoI+LtakgxaUjIeK+EKjgn1oq04jwa/wA0Z+WWZhHDKPl
EcRRM0rDDlv+MRBnj8ZwpGcZFd30Www6uJNGVs9mHrM5o7KyDaRJdcG6mHwu
1c7KBLKHe/yGJve2UTlXNBJBmuMgNI215mBs17or13gcHDK/643KHYOtJaTE
5/OsSDyvwQ3BoOHHZ1+JZATG5HiTD+cL9H57OS5iEJUwyD2u2bO9RXCjyYeA
2+v9eVmfs0NWPo8sNIoa2FvbYw8zqdN4uop784Ci+mOy2sWhCmoIndtHOPTt
F3GDIXieME+LYLPAc4N0Lr5i+wLSff6oIyIKDys8Xt3uV51LCjg9wGX4pTyz
bVUCd1C+2rRXcGnCZqtCAhzjkTWGmZqGFNjDatBytZ5wGlZZ7ILE01BHJeZY
JxNPKipMKRe+7n/QHgG5LAHNgZg58ut75guV2yIOPaO//o6Pbqa41wyqUoM6
GEXrifhuf985V7QGjB+WdJHOxvbOxXx/cv8q3+QkiNF8XnTWBSlO8VD9FsjI
EXqPPmlHBAJhQ549ovM3H1hvMuVHEmo0jppLZNrCDtNsz/Djt3HEG5RmDM7H
RBxVGnayG1i5xYZ5v4OY5iS+P6ff1oy2KWbtx39l2VeMy8yl++mr/UdnndCr
MXY1TuMqyFRrbJQ2kKe4aBW6KNjY2ssZIlmgqI7EaMRo/BN13Y2SZvzuSp5z
rnSqR2fUJl36tNB1ySvL/EPvThstpfsCfA55zlSJSxywnvGYvr5UyArjPpi9
FGe5wuC6K+LhphMfygAHsb68A/vrjcQTcP68oZtZ2/Mi/4ypIRb75yYDmnou
q4Zj8CgrR1opPXHEDLzApCcM+qFRvujzIbdrsr2BcIskjVNnF2LVF4mQMvx/
NimUgQg6S/AwufC17yEs99KcP4XabiuBYd7qBjDEx5/ZhgSaH8l52nC33zcx
J3s1nh4CrumBFS97q2o0tRLSeXU16h4HFpaS1mAPax0DmtYZSEBawyOg2fVD
Idvzb0kXG6Z5W9I4HatS+WvNQFh97wIcnz/VUcf5B6jdB010BUC2hFZIhFS+
WEVFkxJtmUrXD/XXqFRkblwAniCyP7AQ/Yii1Ct9pijeUVH7tNOphMrhaXV0
4IPI+F93AgfmoJ9V+NK/zDqM6Lzcs/M9CkJgcwjvj2STyXEhFD3EodCVlOcy
HjxPIEyQalpQqAYxOBu3BqTS19YlUjRkUTZ/xmJE8qgqMzPbz9qHyrZowmSP
ghHw9cXhMoSEaRyZH5JYqFZM6nEFnsQYQFL4i7LnRPj+TEK8KvY1z9kyKq0T
8bYTBTUdm1dp5IZooymH25u2esEzVelE3KpQd48OsSM5o9O3YZvBG/5NIM+i
DX9ldSja+yNm/TSg3PtYfrsXb/zdXuyFJzpVIAJDXTzF4Rx4WbIZFyvK4w4S
oh6oZI7sUW+Md2MsUp6wePB1WKFOMQX9HSPtLAMfoZd3Zy5dv6u+rh81/edK
6pxBJPY45OpYnOppHabivs6Kao0WRDtdpB6i4i0YS4p0fn1mzppl7e32urK+
yl4WuWUPeXVZ7f4t6QuTh3qxQ9pxBsnNNn/vdkEP6JWlaOEJbueLHL4H88Mt
DohJWch6zCUbt7ZThjKxgoozdl+YiOm6OQtyct2UEwuwcvlid3hAO69NCtD/
vWLCuAc6i/UHLU35jXeXpj5p1za0pn7zaHqf7IWcp14IT8DJz/O4SZYf34ND
zNkcRsCll9r9lNYOEOi2Z6NpRIHfgFVaYNe3Rz82esVbJSZOeTscG390Fl/M
duS+VMq4mdKzNMnPFTWg0fsT8L4JbXOybkrUY4hWpbBXxAwDr1l/2WEzFEUj
/A84OZPSNeN/+lmOc8L2mf2XTeg25Mhfa/m1mSOWjD+niGiIaxNNRVkaWcOJ
LP4Jd6SMwjmkJwwVWkJC2bmgAvKv/iJ/fAafOga7V7Arymipn/VO1NkkrgxG
ExvHhMPhLVBUUZH1uKA+E3Tju9gwcXhuuJcaKb9VSB7Y8mz6TmqpPp/S7Rq0
2RzPhXZuQY0kEhfkAD/6P2/2LVLHaPQw6T9FiQ39qlM6LW7JxC8MkVhhgrux
As+8wHDxoTCNaKvWJ508rJy4a35k/Xqyp0J8fY5o5ocpvvGLdA0DahKP/10i
SVeSasz8wPyPP4JXt47TZpUIyQOhaO9RhI+jgX0PyY7D/hLaqr6xEX4CxPWz
tb1CN/Aj8JiAL7Vu9kw4W73dF4iCBLEDwq34ljdV0Os4+jnCL1pz23x+IcKV
4lCPG2dIHWpl6uaYbQEH7Ixp3JOOGu6FyKun1SOZf2ompalucVlFmBZyGDl5
/cyHgUPQ/LU+HNCvESfw/yxsyRxmEA5qNnEsj3+rd7jJz5vm5iGtSBgIfV1b
+MhD8UA0MzBSHLplvEKhM5cTYe8OOnj0KtcLryBQyB4VuSNMzBZCHZhUtjDf
fNdvUxx8pxPlzGdmhXIi/DYkvHQ3y0qCDf5cjAKqXQEFAVT2pveck35hCX3T
JKXH+IXYeOp0LZ+42OuPIrFnbv5gFEW+quMisoI8o/Mtsab3X6ajszqa4QO7
ld8M/dMQu9G3+kz1XqagS+PHrf9fnzn2YSWZ4fLLRaaTlAqXp6IR5LTDfQ4j
0uh8vrd1CJ27HKQ7/5OSsHMHITpKru5skvtBv82RHzWKi5xFVVk3OBq6y9js
prBmrreCRVHw+HeBY9yGxLWK8zt1FMQXcsX5XD5yp1Ze+OZ3GH637M4FxkIT
HRg+20xpIsAh4T5Mu26HQDy9cHV+TVrUPzxZzYqJyBAtAvi5o04WuFWTJQdZ
Gcq46FlKWtZhIlkgAnkWkzPkgbrlDH8bDPvvbrZRuQZKs35Ri5rpQCBeZ5fj
PIBXDLtvhvdP9kzoCcP6vt29KjoCsdfNA5f8GTQDO6ZomJ2j179/eXbvS3V0
7NitO79GtGBxKyp1pbw+fey+whgJIPxTCfml5qy4Qstzvo+OwvZNyejCKHMS
nfSjWF5domDH819OtK68YCgO+tbwtr1NDqznnQRhez8PfPQo6+CwHY6rLbWw
cJDmLosD7H2vczQmquYIdYLJRAzPAy+Dkov8bqV1RfVjIIZURn6nn2595jUu
+KDOevO382b3uLGvBR/YQzKCkNjLEEd5/dSGmA8rnho45dEFFS5LqFhO7Glj
wLXH/NZ0hX9Kj3e250KQJabTJIBnqJTGSynqEpophTE4YVQQ2oJWxbnE0aie
6vqydaQ5cxqbsXokYTkDLiPupZnHTpIsCG1G7X/9Ob4C6zqzLXIEB9y1Ri9I
onKizks6eupX8VZ/rubIhxgyFONDPYerWLW2i2yeddsd5eNvNSUE5HOpGK7z
LSArZNJY0jMsclkDlvYQUyJeNA01fcOaXMGc0PAnGj0zPq/Zp9gvbQ5tckJ+
6BuI8jaRE5+kEt5ZBrcm8QSBN9Ktp76UWLlNH9ARIEOX21tlCZHnR5AR/Us8
+UQ2iqwBk/Y3wuTJwoCxGBOpDT/4QUo2hERUJb+3U8nLM4SYPl4cqGI8YTdS
Q82WAL7hDUDR77YVu6jLTkZRc1+OcWljTXa56CazerBKWhQzj1hkxs7Oltra
sP7/KHk7I1UZpCLewvZuilf39aELNJ4OF2OaI+tKdVdi4n8blpNX4HN1BJnS
zidhDFBXo0Q5ggvIGhDlTDhSceNObIJYMbogPBrRL8PQGO1BFLdCf3Xev+69
23XSB1awlDiORgQBh/XgyKDq6USStDHllSq4/bNOguKeYYrzdFxVEPxlyJSI
vhOQjUm0oSaADu9yEg/r7DMHPWE2EckyO/8UqRr20Ly4R9k90xxvdFSHQ3eE
XOrkpLizisMLEDnJ61Nck0R3U+q3VXnvDfymgYBUzpOn+B7s39Q4llWHqD24
0y3KtzRbuVoA6nrdj9Li/qf3eZv5Ixgux+V3KlyLw+klBj5KgzV1k+MyEPHj
KyGJJRwlYe5zyrGv5H81Y5pDaHAwYwd9/xPVZBNASN7JHhchq+9kbtC5/a88
+KW6XdXHjKfU7Ua4eKorntTG52gFM7+mrhvQ0ReMbXaBKhnIDc8/eN7yCWdM
QSq6mbLDihVOLF6ivRXemhaeItZyt6RJC5jtks6uniISEBt3avb8Nhb+7ABW
7/EdG4F95g2+TtHw79e335abfH76CzSNrXWKuWdHtVbSm6Bpa6uzgwBmCRlU
3K7rx+vS17Bm4lnNdY8wgTCIXbdLM85fSXke4yUdpCleWet0dV4wtSlA/FeT
0SUeE4+K8n6inwRJ+RiAtbQh1oOFsUiY1wz/yaX2Kqgxw08dRHc7x8cUTav8
ECkrJ4Bbibtcb5hJX2EsZXQn9KCxN7cYmtA+VO1Z0P8AuvbEyCx70T8D3GP6
CI8Gt0qOB4fElj4ZF0JCcIG6MkGDQ5jSssKYDnME4W8r6YSkmIn+VExXwiJl
UmjX7m+RuCO1oWWc/EICIGtk6zCXWHFa7mlmorZD3YHSgGWwmFKmpqwzc0Tl
/4+g2EeRkoE64YIokezWIJI6uICYEuhW3K/518u5Sieeeef5XmVWTD4KWLDU
0QI87ndQdTMeWwEm8L2t1Lz36B57riQ+sJnxfSvMDS59SIZGcfZw5tFkMPkR
RgKUVmvvhgs94UpgMtn4t+etzqsyWDaSMaSeaGgJroWQb3sqAdUMlH4hXC5s
zmcN3QeL0o9h+ZrIb6wBQkd/2Vo0azr8rheVJHsYwxVYOlqgwZGPbyeIOvDy
/prwEyNsbr815eKPoZtpy5G/h3Q/piVK/OqUw25fHql/UBOupRAGc48NDOQI
fOOfA5BlG4PImPw/Xrqt8zLHGqYFCsrNN4QeJ/3xiBbdIG/Eoo5j04ScoZqD
UFv+Hr0ZoHbOUg0s+hdttHic806xDnRJO2OyKr0kOqeOdTec/LVaioX4PfLb
3538RH6c5LrhD/3EX6idOrCZjHl/LObJgnB7a8wvOVUr5lyFxkDEgTVHMVwX
5ul/er6V871lJqrqT4tIxfTqp73wk5nuIVIwJL12lb+hIl4w8DkViyxcs+9V
6bFq0PGr4dOS7f4LEoJk4wlfQQnI637+bYI/Rhd5j1+DA4BavfypDeOeQnKu
u+MMuzqnI9jI/4fuRozN6cwFB7VmoFY+sNn7xH8XVWmvc4lIhQDUpp2wLlbV
9Io7rVDCdqosi8FiEoC5zmXolwtzBFTxYyMVLqn9btOZ3x/MPKU+K0y0JfA9
gS4qiSBc9ryJnuNQK4SSTyKYJBsD/lG1HxoYbbHxMn80H1eM54enfGcR1Lma
ahn/EtrpLOlyomZCLbDQUSQnlNl598Zu7x87zqRIpn4dUFv1+cgAM1w1qHrC
pizBP6EK5G36Iwol5DvYjK82fZs+lfHQfnq0zeGd318GfQi0JxpXhRhidkCF
vrwMrS6tqLUSHXMCAb64Z4vZLopQXvHjnE/yib0z/i+70fURWcMvfGxpLStw
0DpY2aGA/55uyRENlAFTFb/Ogtr0W4yflg2YuiIp+q6SYwmXIShTtHy+N5Kk
YVNHBfGciBBE4+ojxIerKv3huQIkKBPRhV0B/RCG0CwRr6ViMhtAUg2cDXNu
ybqCmsYEZHnOITSZoPnoIaBhzlVdMXrEex297eFpuurN0R2eaXzDcb6zJrxD
pCxBJmLxeOJL6DALr8j0QDRQ+1eLzppiUQkr1G5E/46EAbi3mS37iXbh7npu
ta/NnsohasuxKEfuWubKzH9i1K0yS2U9u21Id8AiAWNCBwBomQ9RWXWpsAnO
DgKlNWQYJfvzVXcBQp/dpJO48GwwVAYyc5foD5zDvxkG+tdYFQ8IH6ad1ZGI
Z3QN863oFLPhaKtmRjXPE7v63JK3GFrobyn5/UOnLwdjnuuMrFA8CzhngrsS
S27gmnzOUZr5hhLseFtBJr5OGanTYRPBEKTk4YFUhu/K9f+kVzT+7DW8c4IO
WFqeVfAXo/vxAWP620cuI8sxlYuo2K5GKSL2pR5FSjeFWM9ukw0XpVu1DzwL
YlnWwODveOpEjVOSnWUxI0TDhNmJ8S2edhYqHrvsTbAecnGfewPrefsJaJql
zbbIR0MEh0Bhk0VOetvLTG9af+Yv3fVOjafjz800p4vi7Xwhpmb7DzqQuKmj
pO2y1C/tyPNk2NZ9ZeZfOizYrTGe6T3+deTQvgP8iZs+x9xOcola6+P9i7FD
zhBe7HLLRXgQOExn87Ho89msi6crw3SH07Z+fstFm0cIlgP0cg3vtHTdp2BN
ZS780KkZ4L4vJsA7i6SyB4KC1XO6LnoyP9xyK+bj+f5VSi9DJMZGhrMft5ni
EDELFKBVg1Che/dPcELxk3pT93RIEt4f6Hp5niz0G0FwBzKju30ySEqD0E9t
I2geksb14RPZ6pbNREpb3aLZj8YUiqbvYUwlikuIj6NOpCqFMzZX14YYiUN5
ewpeYJzHAHbq+99vOkDpCYfyL1AjtrZaI1WLQ/4PcThOFiUpLOKDMguA+LGe
E8TBf7ZA51nDmAeOnDiKNfEwVms0/jDaBZA2/bGTZabF1nXSBII+dKQNVM05
DASmnBpKTXJs9Hn7/8zQK1mnR/CmBdVr3U585fUtjEXzSETn7fXrZPDY52Iy
7H2FHeF2cjjFSHpNR7Dx9sygC4Zbl6I2ncZaD+Zkozn10LQfWZNkE+jSUBZd
wYnDgTi93IhrkCd4ANQoV3uyI4bEfGQebQZAUsuRbFTTjqL6W0rKsnlxqINn
PHmJ6n9LsiEMFMjy+YN6pprYw70Oz6aRq10S4xLoq18BvjCntyKgG+t0EeLc
oppOmKw9SBcsjACF2Uun8VeyCvmMKKV45XncUweOlqvR616H7IBZt2ffdXOj
Vo5IBCHIwOj7dUQaMj8P09fBqHP8UwVUpeuYBxisw02eKTVb6T9mhSSJlppC
+/PpLmaZAh5eAzkGyaYsb1qaG71MaM/yOW3EcBxpd26MM1EWbQiaQgsR8jo/
0Z4bataMCWfvAZqFcfxCZ3Mv9WYMEKcloQ66tcneCf4I0s8ayJ7Lzt8Lkp+v
FugHvvFsmTYZla6RjmXhOkFbGIoyOJcHUMpawX4uf7mQc+HMD9WOKjykySBB
eXqPJq4AQG9NyY/JsT+28qEXkuPJRPjGGND4RZjstt4b2GqsiTDlbslLkGjJ
KLuy3e6xCmRqtpfLF1uXcq+CEMLW0G4LmWwRj7JatphoGcluXpzAhidkZnmo
FpUmHBEf7w79LL7OIu706kzhLV9nuJhntG0xSJRGmd0sFS5+fGUIIo7NTijJ
BCSlYxqDR4J/biezqlZsIx5FSn+5mQSDz56uQFkANHgXtnqFJT1Z//Yh1FY2
JcEHB53lv4LfTbubxtgPCedzKXR4zLZ5mGf5GZnpmkPZxEflz9eLmPPWju8B
qX1XhvQDtY9zseFYbNntgV/el019tJnpX8cpSAqV/ataIrZkAijsePsTIRhM
cfkz+9narZaWIT2vbIhzkwpPZZwJQhym1t7BqStt2BHZXL+JbJ0OObvGpiNN
1ZRU/Tb4SPQVcAZk+L1nVLX19kB30zGEl1RcKvdQEmRUMuoqm+fOlNnWDuKi
Y8a6dSE1II1XSHLJC1y4qxb0zd/u3GeY5nKBfGLwcnkpCZr2hixqD+OsgciV
x61ZNmV1mVe5bUuZy+DoeoLENnRiV6Hbbuwh7q5K9AI6RNTDxMZgJgpKugCA
YCyUJatTY6yp7QPrYOiG3XlSJq9z8SezE/mNBGrVT6K9ywLXRj4bXvn0PmdM
VYiip1bptMLfKAIqc/qV5AVzsetLmX55mO4fR6IGh+DwI8apIsoEyzUa8zuM
cK66PmD4YVemOs2lnRcm+Rhm8JtgGK/Q02DUlsEBDETwxhSs+qDiDeYcBjkS
emQmO0eWc06Jz7t3d4Mui+DtF78NSswR5bRVoNrclyeiBsJwzvZa/Kzvscsi
jVVHB6gazEIP6Rac+52Q3V5FzrFcH37xmjNm0sydmoOJlk4vY1GvXSXGKqa1
1ybE74sATXWosVUuXtuXG+QtqYNjzPTjLq9UNJtS8kiusdZHUwtQOjcIWGVC
LWluItVbrOz/kkz8GI68SI/qf2Dy21j6SVY+URmlpxvbPpYUe5JBEVtyNE+1
ZZmn1E1aSZsm4ksAgNaCk7kXl1Kwk+qJ6nC7047ifxfEu7UAeAwENMVU3MAd
qGd0M1OP7MZ4MxjuO00k0IVbKKtyMYlH35chqSlYQwkyNLB7Ku1poc2BX0ZL
MNbVw/rbaYNZbh12+yiGA84uOeZd0A9x4qC6Poe69zvDIH7D/+0Dtx+snbDx
1sQSqtL7f0Faj2PvyGSOX2rNNeKbjt0fhSu01bQKT5dlMJRIHJ+oPveuNiKq
Bd6JeMlX9H88pB3Kzmz5T/S3mnJAjxbemivM18/IZA8RRfo1++9fqmLClLYB
0Aj+eF9LViQ42b98wTJhTq3tAs55BPIYxmL5SbrxedV/O56GHvXLVUA70HiW
7sUX+OWK8XbybrejWwi/duKJhUr6dmUWgz36KjVSlxn+unDLhRxO2on4l6UU
z/SGZIxAEP+aA62905RCe37fGCI42kdy2csjpg8MddX1bAHvtkRA+u0Apc/l
yZRyelDE2OGLsPNJt+Ph3ZkTi9Puoyg178MPWGk5V5+14Gi2p3TJhIWwsmmq
3jT2go6BHsNSlPTVu7I4+0oq+RtzQrFodyMYiU3uA/SNxjLlu7i1Cx3omB1n
I4utj93El3nvt6nRDUb8vxw6M2fqbFOIQTfNXW8xJ+yJl2rK5IbP4o/Z+vbZ
m7skK2Ggyt/80M36aU0jIivdzGHKXWnf+UBRf4W0sWqEBn9w0axiLh8FlgH3
/Mb9veD0JU9GuHr4Iom3NDnyL5cbeeFpA1z+nyKHYxQOcWRIJ/M8tJHgpT7a
K0pTckk/K+KRWR119qne+rUGpjydZvipqEXfY5ZpfAK7YyV2FK45j76ylOtf
8oU40gmrYuJIOYWuGUemlQ0hN0YyOMAe1z3JZRLZEWYDb3JqkcK9HVZ4hjDX
Qy+Qv1eXsyUTuuPG3DrTV2LFSy+ZArjeG1zJrigwsbrUhk0oUSqX37U7X9ft
hmMuUf6OTXjP1+yO4MJcOa/vRuOsaY5uqfeqdpCsj4YdzXKOCrcm+wlNFAlK
fGhLg3GkAmBfFxaekApAAAiLoimdU7V8JnwuTeI8i1yZpVpD1N9KDOABqK+9
z9mnkl+hK+FxskjSFy19sWWRgw6oippWDCu9Q18zEp878emfsGmOx5/ky4bO
rPQpHjXcwFrtWNwkK0+QkiyQTIcGOzCo9NaHhOkHpAwuwKNbWJeb2P9W7ECy
MTlhbmLPV0IVX1RoRu6yZkOt5Enl+MXcO3tjuS50MqGc3zd9HswZSyth21Tk
oqyIwds9fv3M404bW6nrfoiBO6YrxjXyBg5+l2eHpvly+SZuSVtiQPKIU6h3
r9gm2ZGgkYmDAUyX28eZid8owXbrz5JEZuKVy8g0d93oViHCg8r+mJ1RAb8T
/T+VPW3dTp7TY7J/sASowUfd/Tw22h0NULBtD4kgzmSZRwIXxq7YM5KK6q3x
Jfdm1uAUsl89XXe4eXIKXtZi5feZ9a1BszL76bipU88vyOWQKWHQMl5ddLGK
oAk1VXu6GE9MYBLXIo1J6ZpGkasHi2dBJHD648b7Fcz3QuDSbkymrgXEsTtO
VE5QXMPysfXx6ukT/KUuCgHykShicB6TQZKy/0bWt4FDoEfTTJ7nBT4yVSYo
UELOdqskl/lVuDLiWxY2IMa0Hrs6ZAjZAs9v/hFZRwRDvturgKbbRsoAyTOu
Hl/F+mlE6cNfgSpNDVmvgSgesXQeM84njodSdYX3uHcHvL3Zbutrb4I6qX2z
cFa4ATEKt74Yo4kt1kfC0lWpvwtz8gWk6gVTcV1h28SanbYphtV8Q+Nciv5L
mVwTRzsHqA5KqaIzkZ3yLLoq6JKvXXxjYmRDlOLSyCUwEV8mjnCqsdPnA9t4
mH61BRI1N0RPtHDkqRn0LoKQhbYlgDbvMvXuV6GzSJ7sUHh2S5jcoke89nbW
OkNLfMPomZw5aRGZfAqeW/qv6F+DmETAqi0T7R6JHLe+abp9q2nNtxO/l7Bc
DSZPuq7HKS3isd088L3TXNaKPmg0IKUHavhmRH52GMPEybXskWcOM4d6rKHD
J6Cvuag7Ao4M7e+IjxtbX/Rbfs//VSfI4NnvxdSyciAmIK0Tj/7WjpKjdRen
zhCEE+5VbpGV2VQe6/82JOu9QqGKYJtf/kWInmN+HjChFqb6czt7AJHiDOsr
SLeAAzbiXibtC41R9YytDwKVYUA96qaAr3WVs6HhuZjQupLoRNMjo908iAQW
T9d1kDsq/S1/TY9Y8+3Nh4pKx+VkVNj2kAME466Hiv6juiMIyoxIPM51CCbA
zk0vK3AgRkvXV3WAw2j9HwICoY77XJhpO7NvRM+m+oUThk2YcB94qe2upCPA
OIHLMkNSxUYPy2NfzP018oZ/p/TYzSVLu7ksNCig/0P6x6sCOoa/s49g0Qvx
MDIPQ+lBg1GkR0f5MZvkQ4SaL4eP7dR/4998QxKf99TA/ZEzQvYAHoYFvVRV
bw3ysX7hfScbTRKYlWsBhgMXGRjW11LqPLof5cRnM6sVizqYAYRbnYiP13sY
DqtlTxSJILDy4rRJjIkejAjZWrA0cdFGzByOEDx6DqVqjB1ebWuNsbxdSZ5y
HszLjOBWW6/o2poR0cjIKGJtc639uL086NBjCWiB7hcrjpAal2pjTUoQuIR0
6a/TCQ2XOZzYjZBazhQ+magOaphyI/rFwZF8kfqV1IaKGStu4VTWkZy5+dkT
bdx0T/BQJTqXLBqfdfzx265f7G8MezhKzktRwSfHv71CkqZ0AoQ0ABajlr5Y
cTMhxYwz25hpLoeMkNw8D488tkM1BnViOO8foPVa9UQHigFAwlhbSc/NAYvn
W7gMxD5+fQAxne4qJTjTTXEffZslyAO6X8aZrU8lJVdV1YaPG6KLYkWmgnYp
YP8Pk44aLO7Ii4/623mhgsJ90Bai3B+9mIa+fSavGsxe7fHNqcZ/haDMlIbX
Ls9rZjUNke4US9ymdHJHOaBZd6h5OWVeL2S2RwtbkzqaC7lhd8B/BOaC4Xno
rNgEJNPVPcAUVGus/Ir6dYRtQx00FNkrLR7NPHeM3EzM4W5whPQpGR7wz1vm
QpUEuhMMFPqYZB+gS989kCaHAo5R7IivCxkkD0316+/+/OfBRlhbKsnn8i8A
2M5+Ng4yE4uSi8QCC12Udkq1aRU9x6zUpSPhPQI/t7YKeMowKsqncd7l8UMU
5/KDd1SD8eZxqNk/HvGMpfIAvQixy6RPqnHXvvUkYYmJc35SC7acmNxcwgH4
kIpW3YunQZqBdTUjrEw1rXMcBhu8wGGnnTBT4jRK6eNSu9BX6IL88z7WYAZC
6ItUlzYH31mhpAUCPJu0Pi6XM04olL1h47MGltQtRtC0JDZNXWuBXJo9e5H4
WslxNF7UZsVoRLX6Kc2vUKdhL3DAqIumtjX+/gc6Ci2Eb4hlYPGQAZzxqBaW
jtUKBS53XvKqekB3od7SS8ETn65/X5EHq9lHGDcsT7NrpjgBX8BQR9VGFoTd
RO4A7+0fNKDgunGlzCoMLAq5dtAcEmawmlqWV89sMOGFTwHHSs9dFtW0DfH8
0c54ojAQMvRr8BPdhepE6wONClAYCXhHCR5MIv1bdssmpFtUfCzVq/DdbqrG
q8+5QqFsvXsteoAFzthRmZniOZAYBds8qFi+DH2Ag+a8Zqfgs6LP3UD0mHnF
Job0gnD6ce65+8dfbCy0+OBqQLmRVwR3EY4mIuYIBnPc8lnF9z8xA1ebNYb9
w6CccKFJgmhMSzdrwQKv2AW+/k1qgbYLZIi8Hh3vzmDE9erMxKibn+8vnVmK
o5To/7rc86LCSUaWTsgoiNW6PnBi2Nbu0rZlNMH55ga6IPMOMU4j1660KcSY
jqUQ2UJsu2fsYHz8kViBSn0xwEsg2Kp+sucTsnUzgmiM9HBLxT14NOcHK0Wu
rceCP8vY3fVW/gpH0VPVnKLkVXKgafRZlw3QZp//Jsy8lGuyjKUvFdyg5C2O
wd1oGawvKnwYRYJXrLsZepo8KfilYXm09zSvSCScP770ikoSWs0p1Hcr37Gc
QT1lwU1QMSmzBhj0XK5gsmmlejH2+UPuMc17CsmizDBzvLgQZxf7lIpOdmRR
8bhZopkFlBproLoNsFByGPzxF8EnRGe5ep/yCaen2kWKSzgR7UovxhmxUQrr
XtyZbXJ9oXvZP6BnwD+Nj4ceGMpP3N4lEcTyTlq+Mv1LRGPZRrLUPZiuBx8s
6t7XRnFNbvQNS8PqgLQSvxpRqNyDIWq/pprtgFFusMabeK/6n0AUn+dzyaYa
VJLfGdkQW4TPwitF4Vd5w87JAXaA7f+TR8Z6gqTJvwx4lN1KU+DFV9RVPGIr
J5pMgDmc6kjmGQPDuk9bP6mnEqfX59CGL+wMMAPYyG6DgxHKTv4pEhNfQ6Bo
OdTUHOba3dkglp4hrKvvrGI3KqPQoDdCNZeXaN06VoElXGdxmhfB4rcV65CJ
sghTXQd82eVjtvAfUrZsGRoHq3JoudFiTnopi9tMhGiNVK5dAlcRNaxe3MP6
b3TazseEePLJn3TM4D+j5IxqpJlzPz+iavSbIXYgIttrrDsaogV63MkHbNfH
hP3QyDLytnRUqixqlge6R6IfSWUVdGz6tMr1iGlD61Wz91hyVdNhFIBQAWAD
N8CfPEtqObMlj+m8+24NJ1Xmxy30hHU7vafW/WNAar4qZTxtMcV0MP2qJ2KO
+fiV1Srti+g3NPmgiYR8llZKH/Ed5ornn0wnaA+8hQIurCIFwgmspzqXe0Nr
p77rHGJqsEolJwTPRcHXzZc4hDyPdbI23ifRY/UQ7Qw3x7XRc7CCMNKAEDPk
kHkPAgUj50W0MwpdYQ4EZGJw6iMcq/YIWDjsrjIQeEJYcbvCp9xJQJpJGnKg
8Q/S6kS58ZJlLBsDHHEv1mxa6CQmp0o+UgMG+CQFujYSWcuk8cH/OObYItoc
+o3W5S+muopYnqdZF4i/7tyBrd8dWVaBxfUZPmDwt4eJXoivRq2HdP7PqKQ+
8QBknU0TklNO/gCZ/Uji39v3Xrrnf/3Ljlx/gVLSXZ0ejzCQzadEJ/KCEby5
4MLKumaTPrA0lebyJcHkM427sko2jvcqxFhjJTakwOlV0zWj9XuFZwJsgjTI
0SV8O3USd1qoisvJeI6JOVwrkbE4HyHofLmGevUrDgX6Ux/GGkRfrpIc5FRp
NgVYebkUfJg7+7PfBnG+Ai74QTYYj+ZwmCMxIlQwUkkGQt+sHpr3qJgo8eDl
qqQLH1H5SMEi3mcr5fEEBVpofjUB6Q9Dk90VNbiFzp9fuwFlUvvTlOY74PTt
cb5gLB+kHxeLVxrxAUGVlglVR6Rq5lpYhjI0LtOZP0Hyf9pI2Dsm5PJiA6un
Q1Xn8lKLDxdCaUc2Vhs6hcDcTFien0avJo93FK2D9JHCSZXz1/boLJYmPSJi
BKi/SwkEtf7Bo7p8riRn9EPynigNsyTwEer3kZuAjkPMfEML6CoAi25meiDR
7RAhRAacaGLtFZqSRQwrQM+OWS63Uad+ZzTrJVc7Tvo6IbIlV2U7lfGaYHpY
oUiB+yd1SOoBkC1PN4rNCOn++9tFbxVAAh8b641iZaOKgm//SAfo2hC/0ZVC
sn/JnDrDLEf14H5maQRiaVb4RnpOtYkvvs6WURh+2nCYvVdLOismoRGH3CqD
9Du+TDKZ2OACUASmPZDp4NTbmxJ2PYGUKAx1A4LZsmsIAckD6uo7xuZXBUH5
acefhegw1VQwujnbtf/qTz4+pIkn5k/oRO4Rywww2YmLORyli6AVwy6zBmwj
O1U4C3N0M3bKwPJKrqOz0yPalHbz357xN3JsYZdi35TmTP6QLyEh/c/4OSLs
MhAMvp3q9zQ3n/858r9nDjqTfb9nfCWw+2/xihrWFg9Mc7Qe360amSLFwiil
A5g7qaMuU2L+jJ7vhpvWOVEv75CUnG9CJ+j9MkXSud0SeqoA8m2QMyeutsoW
M4tuYY8I28sjZ0/UazRb18oabDqX5T11Dxlshnl2kXZJZtm1ABIxBq2TcRH/
HLMwWq7auvMHde513nK0r6BZ5vftttyetUVV09lVW1yLzPCjCCoFL6CZ/pKz
PrIoBETWovWSLlz45GUT6OeVTLrZlEu5C82jlBYcGZ0jj62Omz8b0qNlZZk3
MMJOtiBzBYtO7kKict7HLdBa/0zt1Btp2OCeUaB5oyVb20ciHmDnMDsxOAIk
TH3B3OF4sqJKV36tcO/FP4K5351UJLemEXI4tzsEgrpDOCetoNKpzkO9h8Bp
jwWeKhBzCLEzy3bF2pwjufNJC86gA9u5BZq2/ql2J/c/g2B6WzF117WHMBrE
Blfl/9mUo2OD4Ha5OUhg6nzx18bINKKevIDBTexlF47yFLcivCRAUT3cv1zo
73PUwdrCcDIQo4hlyWrX9EMbhmzdr3YnAq91012ty0FxFy2QGNDgCMD7mLlz
y3g3bGV23IFvceYAo06Er1K5b1JdnXTmB+9JvD+i6q1b7b5S06d//kH5fVTg
Pff9wbAJyYflJp1iVNAkdgHJRyd2NZmCcl8QQvsiOFtt4fDstk9OBjQbKDPk
5BqsHMz0cr39GDS4gkvQJp/pRIgsclzj3L5rAfo9FW7OtO4jbePFehsxDESu
hNtW3P5Pw543CPuGqqA7+0zlKBXZ3GrIprhe1A/jjNACvr9CjKsXizQTn5WK
WsKrFquF5RUr6F0rFQ1nY4YVvxEAR/jeEWclLh3v3bC0UUe3fElTHr5Hiomp
/khnuLmwvdAgv3rWzQ9qMeX9+PW0jzZ2/9wE2lsMs7KGmvAxdr7eF9gJexqw
G4WEY4/b+H7lGAbF2BKwsn818VbaHjs/hI8BCWeN+/8LligxeJ9M7A9vkT8+
EVykBIUXELw0SGUXl421xpGczQlL9hxoMCts1ZINpdJa0PjgPIAtuQjEX7n7
9GyTD/8pDKj6cROykAB+siJxSfAVGBDxUcxcI+MGY8J6+0D6rAUR8DVhJSwM
w/cnM33og6jhuJPPTiW0CP6DIwrY4PUEdDDWKaaho1n/8RiiV0jh6YS9cY9S
FCrwbpVOZMPuDKtOAG0ct9MNMp0rFtpVhf4pqB6QBZiWPY5IlRj79ddu0hRK
fNQx9YIZkCYYqyWTxuSwlqzdLoi6wgrx+2fZNLre+5FKXUl0vMTgXhChbcCp
0FzQ2KUahKobk8W7AYielmOPxL2MY7eUqu2qOfEoKeq5JbX3cugIEn0QlpRg
tXdjasGatQj3KS2Dp80nmXES6Ed13cOPo995SO6leqnQadS11q1iVBH/9qlK
nPIWFXUFL/dvQJZILtJYMwFhmHbsilJZa1Uumdd+BNusL5zkcHZiOvFKucmm
k67AeNHD/zHtVPiC+FwxK7gqhOmRQSDK78g61FCwc7JoNPLgjmLsBGt+kp5U
I5ASgRDO9mkK/5ZL00OYt/lC+Xf2BKFhHTU7pU91TnSizSNiWTrLAVtlEcvN
iJWCwDcTbOECzG5Vm4gJgwvaTEsxQq1a0uox5bOl1goFKNfreHrGPjp4kfh3
JlpKm2/OfwSptatg7aU8YQZxD+DHALFR8YODC3HjC6XuKJJwuv+OVhvjLSPZ
QECPSZmCzJC9F0nXi2mPGqFjHcdpOQfzI3qJEOmHlkjS8qvPhy1hYCPfFRYo
q8BXtIp4MGQSfq5vRdv/nVELJytToOCfbWch6m1ZkR6mDKcu4+e4Tu+8Xa15
Qlmkl7CcH3sN5HVQSco7F1V8gLwnyCG4fos60aUMSwMVA6rSnQX935DMoILW
XaVLuz2sPhPZnwcfs8z3DpFRWnFO8f3PvJnPLH5/1tCDXrjOjP/XiXqx/2su
8hC71sAB1SPyvg1GfGobOV1FqMX98Ly0OY3Z1Qme2blxWlg34sDuYChWMDAi
o4IaAk9KMZnxVbAPCWbbSzWWZfC9/TZJRx55Mix8pImFBi1chF9Z6RFewDaz
Rmxhv0d/HhgrvMrsQP7EgzZrUW/72mC6c07HyKZBsxBc4qTWRN5B1797sAuP
1Xglu6//dUztCirxa4t1F8tjTBkgOKAjjQqr308iomoPDcmfSTn6Ze653sAV
Kmrz5xa+w/ooqKUsxL1P5zSoNvyI32XNi2tFsGHVHjJagTwJI8Ymch5EYY4h
CXBwaghO2TJlF+xzQpWCkrKlWpttoiQC7thQQyKUb5EYWv42UCYrPfzhG3WR
MH5w5ClE6lX4rX42LS+QUqhGdckJW5pGgKHoRAbYdWsWME5HQIsae2EpOcWI
FBeMjJ7aFCOfRSoOlgQSlC+KfdX4lQowp/bWjKYUZE4wwg7RZnXX6wnvdQxQ
p5u8Wu5SLzemNOyComk4QALr6uNGzeRqZTX2xv/QxQEdLs2BHsDo8HGXrKVY
B6ZnpR6RWfHVyDAeojUJBz9PTlcq9E1dtyoZdV/prwXqHcNg4hIP6QNrCfC3
pkggRWPAU7Zqh/3YjtUsW5+1ylogZSghQi4BjO0Qd6AOZBBYrqa5lcaRYjg+
vmg2K4UwdYjXIaZdGuSieIQPVwVIjTyzl8HnLKb2BUUWIbG4I1JtiUaRMW6J
4JHcEfxFa0S0eKNTbIsS0nYFat5NIosj0opUeyC8lffqqTYs+iIxe77boyiJ
UGcvp7k6/Z3PZrpcNJkPowsEG35IgQjACiyS+aPUQ02pRpL14DkfRR+SHvpF
DXzTr6De30c4PLpIPVdepegyidPCfrXCmQBXGe1wz8sGe6NOGhEdXfrWf4a5
cg6mc69ZewnK50J7VuHV3SosrHg08DmuYxz1NfpE3MHrxV27wlHDjIHgksL8
Owez2hCtG8//VsLwGvbisFT1V380pSWxW42MyjNVAkr5aLJ7DBqnJgXSfG5p
4p4vNPV795I93SliQPLU9suAgW2N4HFb6U+dqVIPHtigGM5997CNJFjASF9j
Q1Ni0X1Zt9zCII2gL4ut6X5CinxZ/bqJd5BUQyt/UCOSoGISNf5b49i7C5z9
18OiAvYmb8F8vWgYLCssgLbRSf6oEXRm4AOKB2OGS9QSEXip4N0xH2ffqRft
AKyJBgXWVD1PwVsnM3zsltpM4EvnX9axUNu3JhRgVep+H6Buo4XkYEU84NJy
LsLblxKH7NSsOSwV6zifzEiNOuZmqC7Nysm+A3cIz3uo4hOk9p+ayxw6vcMH
0Rr0tZ5BIvcaNyrcDzGjhgHdLeYSgtWe3u1a1LSRlPt+noYj4SFNsrKTLoS1
hXQsCLDo3gszzkTtEtQKj5JyvRfxubsGDb6oFXf99owhtHaJYoJU7RhBwOlQ
L4sxtCXF6EiC+wUIsgh1OGgaosKxkcZlpxv4ZooV39bbjFYFsERF9RJBqGW8
cLA7ZpR5fJf1kBbgIAgkL9Go2cdc7WWeLIW61wAM6tA7x9iyGB79Fj1goEYL
C51AmgLA7IrMqqlsIMhioDD8EQejuBrEMKqUUHQ54Rs70d7XPSQI1Ze0Jiq2
Vy5NBEwYjqBmrkue5sgp7WjLiqNkcB77I2XHWAIa2+zdRHyCoZVrwxtsXX0E
K1r3DYWhDS8b7+Ayi57MALN5piDynuMPbCN17B62BBqdAPQc2qzuqURvUwHm
/5gMkBFTug8r1SuF67PwyLI6tRO/rr6efKbX2B2LCOUYSgFSJkx7rj6r+Jaj
RWDpX4oAmRtOPO64dE7kEnDySIaHjxqMgvqrZK3N3zcxYWUdKiH4cVYUC99y
j04/NXvO54usTnZlKNeQy+xFtMXor984GK+55+QUfjdIYEO2TxrnYAcHVxIe
LA93Zmqlyw6DtZiu+7sYHIzq4LjMQYJ59ZmhTorbph6/tXkYL6fsxa/Hp5ve
nRSQnepBOB7/YZND5Rnc0MVnNZa4y1TJu7lKDXP6LzzQeqyEjICiW06rfIOO
lFOcgjXhppAMfvAJQMmf+EvJ+xxiKnfO6xAtvYz0RfQJdl/LfWtvCCqxnxJg
iIiWma6lkNHa5+1oftMMwpBZ4okjKOqKMntLwqm5joeGAW8ZtmbjS9syC6Ao
BpQFlJAaavyhZlzeBdnVuVeSxJGG5TYddJp7nUj1exGd0YIdRzwI+BLfAJmL
VUt4aXT8xPuuQCH2LL2Eajr3kXFrhxohc0u1k3+lbo7r7NLpRSpY8BxgygEr
1IWea0Wimiy6TE4ZS5mgysqc/yMAD8T9pH6neyfzCfb04SccWMqWb1Bs3e3q
jCn5tm5RTAuBj6FkiuHzJb/MOS8MgMTu8+jgtvMxad2pUdARjxT9qMJKSBMG
0EJd5ensrw2W9Zd2QHwVpFeMia+FRKldoLAR3fXc7rcM114LVjS0Od53vqzK
RYKIUMVVS68tG8noUwUkFjTC8tTGf5lsS5HZPqXUs4MywqIp+cxOGxVGYdvN
AAa0JqU7wiX5OX+DleUNxDG3jLJNVENjUqYBuR23JV9Z07OlpdtZ8cDypm2w
fN7P4pojY288hYbYzFXy7PzEWcZ7fArPDTdcpYyqZV1ddhKyPJfM8qyXdu5B
291/h/NQN+6SKELM9TOjlMGFBqheQq0tANAnJmeIkGNjyxA75UBKnduSgyhK
Ufy+nYvoBViGDrVmhQIVsWaWgcxipM54Wvb64csy1uhswEPSW0fMxVaBJ74C
tVcztRinU1s5+2QCK3na2jkGSqB2+PIZdyAmdaIv+gqSDhMWrScymbFF4Vp5
p/m2LJA9VKnUuPWBBaXJ2/5faGbycZiUW43JxxrYWprG+0kVI75b6u4z+CyC
npJNDjTupcI/Kcwx/VORb1WSQmoCl9qrnsFO5Xz2fGkNr+55E8TsqHPzXVIX
ERUWZtj1bcogiazX6GjXlLxCzQLim+0zql5xiA0X9JNlJomPJZpk1xi9gqvb
uoZQ+n17tRLuUYId2srgM8mN0jYwl5CoVpxbKslRlfSdrKmv8AhWr3FmFJiX
mMWQjksvotiPb+GHXN09n/5srb6DXT3FXksmWjZF2DuDnPuzGkrEFw5Ae8AS
RHHF8NXc56rAG0ccg/ydSAoXC4PnRNtIVoGuE7eyXUwZk4bPZNKF5KfVSs4z
3DxHPeX9WqzrnFSLQNBVlNzQksJOxGiTkThW2JmbxHixhNMYl10K9u8DVlgl
IJcY2F73MSMKj+wGd/cth+Z/DOnha2f3Wb0VIAm4Acw75kMkR60fRz6ZGLge
nGy2WOM2ffkLl0J8NJcc7PxZG6FWHZJsnce44IuRR7IhgDyDuX736B0CxDD7
YPy6B8dTw5zOPERhQePfK85FqxRt/oKMI3iSupGBnlIj0ON7Z1Rlvm7o2W6V
1jZTnIs/lsPHRHHPDOiamsHylsGia823YAZBkCB9Dk76CSHOkIGFBihtCyC9
VVV6oF6UuI7Tm8bwYuDMU5h+gx8WYCpXwXRtXGbP7xh9Y1rdOngVGmxbngUJ
AvmiEKVkfFcLgshD0fHqGGWVz8isVbSvBz7D0XyGVCz5S/JfMjo/N8Ocu0hW
Q337mre61HgqzB9ZOnw24qgRmmso5gN/13imnexUrGvu12Apq4N2BjWwnWPg
LmlZnppX3ph44cVjZE1dlGt98QQoIb288H63Bec6Nxq+rNn6RhRpf5RCfRIy
joOTJCR6lDnSAC74UvmBYUArihiirSF6EZ6OfXalYeVcP/0ZVcgdkjR/do3K
W7Wd1ejFHcAmrvY5qsUtlvlrNjJLyD/qqWmNv0oAkive7b6P87NahjSg8ofZ
07m2XmPoAI9b1PqQs6oIy32v/bF2FAtoYSJtryFt2HPZhXmKoVksECO4Cry4
09BqLP/JbhNLdIREBOKO8BNZ6jDNd32gfo8U3PDSLxzD6Gj7/xty0vGCCEvA
i6suwr8LQ3RQ9vOKFOo2/msYodeBl510ZzlGIVuWE5kbOGkXrvnYO41638WN
O9ZqLWd55GsI8WFuAVvyFIOelLJcnlaQBGH5hN1Hay3Dz4ycVMLjtcwmB7y0
lx4QgWzHz/w6tBB6dty0J0uE8IqKlMlpwfAfa1l1xNUoWl/ZRphgbBYRXz65
9mFxU/gvENzXFEC0H1LJ0AC7PrvuTtOjsTqhyn6bjWc9k6A/TvtnvhDniaxb
fqRBMjE1ntRJO6QHnhNLDCBiKvTkNtwAoU917A0Nh3TryLpvkhbNlgCfpr59
KJkuwqhtv5dAiBK3tUBZbG8u9t5lSAVY5HnqyiDEyFm3mo48Ewo8Nm/EHD1R
brf5YklgP/NdpLJQGTUXxkqx04SI0DvRXa6/wMo5DFd+jppZADwD4HP+hwsB
xIV8Iol5V11lG9QwWnGLGVZC5ZCIxNEbV+cHwg2Ss+nnqK9Dx+ubq/zXa255
3sgwhAGKQSZiGe9yBGIHTDTUDnV5wwkOv21mXBsyX1WUfPesdbhag5UsvDY+
t2tPfJ/2kVAK07fWMEXpPM051BKB8KSuCYl1Au/d5EAP7vtBV/i2YEzpIp57
NIC0+O/UDrd7umWQR1RjRrX8W/cN4T/4HfQl4zpbJHjDG4ZkqudN8sbsUpXr
a4rAv52ao3MKtVsw8SWmCDDjhSKQv2QOZWnvNP2AGODWruWpGV6Nk8BXIaFS
NnB7ZTwfdQlBkf0aVTeXANRzlvBFUs0l8dvLhcbVubdyyHIeUr8RrbyvTcU8
9nVvGyzQg8IStU0KR9u0PufpKwHzW0NjSTP0UKbwq/l+q1daFWUkS0jUFFyv
6ZisqIL4DsDAcUClPHGFVcUVDOZfJlz1gRRfFWZzOwT9GMfhoMs2mC+dPxfL
dIrdvTjuw+5kJw+9RC1ylwpz2XT2WleGGrcyoXwJXTWMcdglTGW7ZJBk/nIl
yVCGRuHM/Nc+TYPV1vtcchK7NsuIP/08nzhsVGNwBwvmDYPsbMuU0Qz5rsvH
nOnRvMGRnFpe6tsvrJPAyWHIJwkJVuenkFOTU2RgmoCUu1Nz2L1ZT+BwhDyn
EBwxBotynxnpwvRMRaqv1iLMRefULoE6aKXLpssxKpXOLXynQIFW73ZKc3GX
bBU4BWneg3RkSLW5juNekPG/B8X7bsTCog+IUMRIr6LgeA4ef4oLSvtMxr5x
bWAtK5ZPpTF+mLSsehmYfjKhSBNQ2Cg05sYwP1hODhsbqTQvHqiFYYA6ZM3o
j2vKFGZ3Yt4nNaGQEF+BmMsrxuC1LAcTqIuSuc1QcYPQjI8sfsfo9rheBQkD
ufug4anq/ZKjkPAYztvmd46Na0Hl4vH2LXKWxZkQAOW55+Qm1BlZlX/4o/JX
TnZO4/yMGBObIO9914KkOdVstK9sDvWszarIwq2vvF4wvsRlXXws1bi3gBvR
CsHxE/UB35INTOyZsR/Dfzd9Sf7k0RqiDyY6ZMl/QSbMWdQijPk9K1mdmszF
V4mxhF2OF7lMhI7k9a8O1cb0Df0zqS6htPg5hqgVKNAd2VhXZbfbfsFL8Psw
+QM/7SzLvVbsfNYKGxhFrddPWsBnXFT3fLfgWBO8lqjnhKHgD5uMTmRGH3lX
SRqNWlT6y3YN/Kf1Wf+1C8oduiPotTHquWSXpGLGdett3ZALj7xI7kbSNkp3
q4TBFv7+3mjuZHWH1n37MTcsoB+/1exBR4sTxIwKdhoT578TB8hs6Bkas9Qj
BZlKIn90hm02fClap0l8ekp6uXZcN9IwcjtmS17PSBp7+HwLRFXuyYdtynhB
XtlSEbLPravCPWm6IN3sCpO7wFpnXZI/QuOFnr6fzaDBiYHrsDcE88QXC2dj
EkH+7vP0z1se3GLwSna5XHj6HoWD0/FU9l2I/m/LKFWDSvXAa7MdJO/1H1Tx
3sHgQSqhHtllN5UkjX9NsOeA7Od4/OmYHvRMJ7NDrRtizyUh6MKHlTWzRBla
LRH7VAGvHiH78oP8XrRGpFWgQlEiFA7bD9PVjap3dyuzoU5A7vx9NP2Qc3Yr
gj1kB6vqQepEGXTmbZzbUT45YlJ6ulcuuKb54bRLQTnbG1190KWrmhaPc0Y4
tfJ9P6IeHw5vMT/Uhe+XU82EBSzQGTJeZdqxl6knkqpV7E/O8GaaOfLKt6GF
eSrQ7HNdBZMGxKpk28mVXsgV+LMljnKeFMuMjHDAGFqvIJThvJZe1F/gwCqZ
RS2lpXoQvWQgRS9RWx1lwcA0QOge9iMGyOTgu9jk4rACPqCGyH3A3RbYLaQH
4vs8Mafnw5vYynOG5Xk9BAVDx0RtpXhQ8AIEaVwzzCYJRXnuTylfhig+QNTy
0OaGMQhokfqZHjrrhxaiHxgWKEoAS+a/uX7cWeGY9JHZigSTYkp/6LiuMIPH
/MX4mguzGCjZdj7SY+E0HiDwF/Quv2yVvOyyzfgJtGTZtzbTKVEQteuYJXuA
whyh/r1QqhLlOAFAy/IJ6fuDEJBexda0MFL7qnpuE8MNHKaUathXacwGg7b0
oAeIwMGTalHuEPNhhbx301VCIBYcbWwAn//UtBWSoG6n1daRWcbZozVHsPHh
Zh/+KTvEJn4U5TGiK0A6z8jYgXQQLVRZA6V6uTEMuOM2fCCNJGtYftzjPT0W
UGLSFV/7fdynmcV9oXo66eGZIYMzP/AUj8f6BP5y9lcYrVVnuN/j2g1/JWTj
6DqQ/y3y8JGpfD0SW4fPnI4v0LVXlVyxY9OA/P2jFAwNH+4puR1Xn3mXqdf3
9nZAMFBweNdJbmf5nN8VIwlQD/uhwWBzeMC6Xhv2hISsyq4R28DfXIg7k+K9
O/nVfI4EwPsBNjPVl3Sy/C5ZI26XWrBRibgNND+igTyrO9Rjd25PEpDzkgoy
SusNqjMotcewbXUVtek7QKf//s0wYVsyUoSz4DIcIvN5N5Hen5Y6OQjlPGGC
2vjTrgHnLlmyEIbPfw1faok9H7ZLib0ztzE82DBZZ3UV4qbOkwAJJP44DZ5D
0gSgDiY0tSXyDY9aWvXuO2hVQJ9qlTMJABiCAVNgYe+Zuu1KCQ8z7jV+fFyZ
czG29n5jXGrYjxAuWx9d8M2VEoVA2NSS0IZ9erGzHRc5+SmRPdeXv6Qqig43
hCLuL2soHlFCeEBPw2unv9Mr632d/c5ui1YOHcrtZUFkK6wFyHL5NQY0Sr2N
Meo9+2gqXcq7xW6ed2Iq4URG11cSXXOCYDJqY1Vr+CaeaU9euBAPBPlbGEBt
PdfZ0sJn4tN1wc6qjte26RvWJy0PqKdnjlmyofE9dPyId9Bf8c4ZFCaS5Pat
VTFrogeNH+YexuNsnMq7qLoLsSq0BDDOxfPFljUEnjEtfVRL6Ix/8/ihUjVO
jbsqnToOg2jajCAh1JZdWRHZfTsKVjyUxAVavF/SOkKc1w+3yOtntb6EdH8n
HNNDKchWNx+D7M3rcpiqhrBIdmGCBKlMIDQoljIxGOZKQCJkc56XXbKg3RP4
XFnjKswJ4DAsobXEFrJXOt7ujtetLKi8gwB6/EGcHxTUZVtXqauZ75G0MNZy
BA/Ae7/ayBikNjIFFrLurG6Ax51gVZUDFsQfJobS7CGQfapFrZlRHiFywQCq
g6TvAamua240slcA9gS2uZy9wGKakNpyKsYUyBfTHlnkNgw+Fp25MoQoUtSi
L/2umfNbiTCY0HVZvicU4rkk/9IWTLiObnDOEQCVd1jgMUm7K0iWLcTtYEnF
9C01eZ0aarKvBpAVmBL0MLx7uZy9pMSrVPWUzU7I9gSAa1LJ1mUM5U7t96fj
Ot7sFxBiT5aS39yX3EiJRl/GRgrmAZ5Ifm/2+rTecddivUBxRJpI91tsbB/5
yTC14sdsbK9ZwXS1jyuwfsPTmpsikLsOeaiCUbe280Zf7jbkZXtb6RZkmg8F
X9U/wm213KdKXoX2U3387JW9f61T5g2FhsHxXUBpEUCconNnPkF35xv7yiZ3
bmodKPab0aNyMv1vmCwsHxoEHaCI4p9heJ4mgxwhR2atvfjJDbBb3vpDIZVc
rGwAwIKe9Oma1p4tX0XRAxb1pCwL95yjXfaqCCr0n/AGUg2HFGxT6332GXxo
TfsruS1HA7EBfYn3wAbISJtKbxV+HU9WTpNkowRb48BmndcgUwlnrvgmFkCR
n68+0TRPxiyAQjnb4JkuqEfpcKi9ATjhV3rRgSTO5DhMgAy4ZJUC/loxi/Rf
4rwEPWaxTzWvP3i0aF0SkBikwmLkwCgYYn/a49An3AmzcUAjoulM1P4mVrS9
QFPB1cQbzB18fennM98cMB0BISOH3xQTHHgwNTwUzEXADeK523nNzV5/68yG
4n/ZRekiRpPHiF4f6wJ/0fxfIoU1qE8v8igvYN5jCFYfCRoCJsrdmkPOc3f+
nCCx853PtbNX9Hg0b3TeQ9a3YCrXipok8XHmDd0ez1SdHr2rZl5/2yW85xiJ
RDZWpjiVJJaOD3Z3QkZPNZuyqkPjT8BZKiGZFUwd8NilyOXkqPV8+pEFYxRC
D8/sj1E9LuYwOqLOeqnhmzWbvVqrCmbK4BSg2t2DLMNnB1NHnWtkS9iD139O
aEB4UZOUhuoCay0nmUUT0uEfjwmBbqaWdUgY1y+foOpL10Y+oYpd7s+xWJgj
KUBv+11TPLQO4sFregJoCcEpGJ3GglKd4ott1158cI8L6JztHGmKmRS+zEvN
rkLla9wzSmJRPOjMwo/nI4Jd5oBMll+DUwy1tAYemSUoGqtC+Ofa3R4maSxL
bbFYuo0GzPwz759Qn1LQRaJ/revzk6EKpEZ6GTTorjvbZ0GHYcyOAM1AZKQF
pjs+d/EiRZVWffyk0sLlMDI/cRBnEzi7aiux7gUUCh7SiT8OSw1FkEYlE7TT
XH3mj3bUQDgwbs0i0r1BRnHzxVuo4wjSPzPF4G1AHkAi/wXgEIHr6feDmJEx
sWFCVsllsNJy5TV4rPmAx+6zDFmexFKDs1GPHICgUBkMgUDFvETR+zBWe2Jn
6vJKAKp69bDRJoequJ5GtEiUIjtKX0uvTy17USnN9OgZK5uHCBxuEorzYG57
hGuezGOvLpe9gB/Tw1+McrlW6OXUoEYnfxN4pWAgwqCTP1G/7KRA9tCrid2s
Ovp3tZaTErsRJz/zIpJVqEwP7J685+Ezbeejh/Ihf5AjmpqyKm5onnsVqjOG
ZLre0t6bQD5DHrxi467eehQDs9cj0xrzUf9uIjVFAH2N0Bb5r5cYATA2Y7zx
O9D7n01B4wcGLQlZ1dABIY2hrzMqjj23Zs4RnWuF7l5tgWX8amt5Vz2Jji4h
5kDBdGfJbI4FCui39Ltma46eUTkBrwP6sggNaud4vj0Tt7D1wUFjOT4O9rLX
goWTBf+lR2tkVOjUeZYyOtz3JIBvGVOBZXXH9qtez5wXo5yGoh/hON7YU9g7
df3nOjN28SuPb11e0ZYmobP6CETUgPLmvcJCN2wSOYZZMTFZ7oZXQVXfc70a
ehp7OsFON3vkMmtQAMuzLTFmVMdrtDSCoDvtacMz8K4q8WBRaDvuKh/tRenp
DFHDl+xiQ1MVteXMVpZD82Yw7Tb7TzX67O4sek21Sc9HaqvFwWSai2rHdG2r
Lk/KhhVW63Nb6NMywy5sVemwC7sPr3M1GGLx/wGT2bq2J/JTlnPhlVUtyhQ+
5zgMOHuUeDQamrIsgsP8FwWtZEeNQd6GKY68iaIbpwDvjsm8T25EP4y1q3r+
gCKjxxTUgkOZagHmf5DNY1BlbJg39sN3/qb8jIGiil0Xj2Z+rZaFIuiLh9eC
uTa3fngOxBLdVHUicRo/bAO/yxLFbrYFC9ev3tlmVGA4KCxDzLTIlzPzBkqX
ns14Op3qt+c07shwNB1MPOpaR9rAi1Bu3ZlfXT1Bml/6dHaduYg1HGjQGa2A
H+L1pSpOhbI+I/as86omEu2/U6FTRxHzOdHoSqtURtK7EbC7CJddUt6URxr4
yTiV4WizAThZGMBm8AZHschDrTD8QOgLxqVwQ/LY5YyZ6hhEeuewVD7PHGav
WvmU8mm8db9ju/idvLYLN+7JXGFRzT/Hwxmiz5tuKFv6zmwV7Q7fuRXsEvdw
tEQPLadeTWk2me04BXPS8jeGrtm6rZbvhp7A+KHlnq0SroFAP01XWgMwI/Tu
sonex17NMNfYcFFzSOS26TGPjEKYsiAPYHaVv0Dmq9ejod80EYTwkiwbfKh2
HA/0C57IfB7VQw0xlbjvZ1DXXtwAKZ3S4lQ7eUnjEys+tXv63pFT5XETzmou
Z19Kc/uK+z9NFM8I3kbMyh1isfl797EqzvoZ+dN6tF2r3jU7n1REvpgpmWpc
Jg0EsGrVNQdD7NNgn1uw1WvrrMbmDyjFKoi0bpFOrFmd8p3/BRu9e2vRDAc1
dV5Wr3A6OMPceEo2pUVkFNIOHa3z/Vr7QxapnPl1HDLbza5IshdKk9Xvr7TX
EahQQwhY9jd0+WHiBRsrTPGhyNiHjTioKh2x0N6iwjp0cVlSilyCftd8hULy
aAwR3nM/5sbUjm6d+D+B1GdmR0BQkgmCwr5EDjhs1Go5bfWoihHMh0mbBljO
LSCHoAqiHhCgflyZLFzkn9ueuGgwrGz9vYFZMNc1iAW9loGPwYIh9g6saL5d
CODznLQjH8B0C6cH8f08SidYNzD6/JhFKb/mI3xs+t1E+2NjKLrUJGBT6u/t
JLTZPHimpE/WyojZK3WZCSEjNF01Rlu6OvujmhdSCnW3J54qcABTaVD/ad+m
3ZD6NM7G2wgI8IswmGqHSDbVK3hkG5FwMyp8H82hW4Ib8pqKaY7qiiNHdPyl
t9D0VUxpCyYHdj7cgAWXKpNiw5AvkNiFoRO/gL5s2X/ZCvhmIBdwLjQZzAba
GYNxe+s8ETACgyHb78xeBv+ZwoxUK0QjQXAz9JI9550XwFxbt5O9V0HghKzt
6xh4deXzQKLeYtBnE9ICDK5944rQs0UGatNIoB/O5LtqhWbM6uQVrEmBy+VU
SqTCHldks7U7FZgfSPA3qFxgYPo268EUEFdlMpLITy8NHukwCuwASLD8qjf+
RN8Y5Brszdt6TgFJccDuW+aeosZtpfrNmRXmIYEUyAQJ7E+bOuAovS2CHcPZ
ifM02vFsJjVjUYNileaQG/Q5BUgk9+MW7pUF6RWAIvr52FDAJVULy1aUSzZW
UEKD0OVm/c2zKYfaBXQSS1asVDk6HDNSSSx19f/hDKexCgBLBqQ0otj9h3Yk
ZyX6QEuyscpk3Z/6WKSwFwT2sStz5cgOtCpwVaW7QL6aHZYXNZGS/3Cde/x0
sPyQ1K3H7kjK/X4BmZdjXZGhMzpDOJCBdO6ICk5ZAWYxoRnvs9YsTt35zcfw
pylpDAZdTNVJQW8TrmAOtq/hDYxMC4b9kGGxa26FFiR51yCJjY1VkYQOjzLD
mWFtvdEVlrz/94MoioTblu4+haYwTkerzth37qXX2nkR7mQ+2kx3Wg74xjbr
SKjmLUQ9OzUEUqQ1BOqkA7NFhUB7Vc2PGdxu+tN33lZJzaOPHiaAwir9OZKJ
ONqAD+u3QzdE8bUnS5qd5oCMMgddky4qbZ1Yz3ASraCrV2idj2VQfSyrKRgj
/dZPN89kBpnKxT1XCZekwe4woQqnLux0EExmCC+yWdkHyjb4RqwLiM9dBv/0
txptmBRMM+5PNIEvUHPtS7Qy/Oo0aAx+pU2YAWtIQNc3Ab9Dy0F8teMq2UHb
GLnBGCbpIwewxXA/9I3LiydXZwQpW2pQVRPkyjYxN/hbQ22uTkpNsuByILGM
KHAw9AAksOGX5euPxCjSlUJ2H1B5hv5BvSnNScHvthbQtev2SaP4azmUncym
sctx1xV/OuywVG13QSlQnM0SgCh1HiXo/lA84RAWGJoGfF1BSBWTZD27Raun
heTQPuAWx+HZZUpwMWLQgmSYCt7Ahk8LIMrnlRb/8+UP+zufdtfvc134Gvkv
50t/kuov53thH+myHDnPo7hiYJvZxw91NuZukONJPDD45NSTnBxJMXa89Q9P
OqNOcbl/Rw1UkDfBQeSwBlTlK9Rj2Fkyi5G+mvaViP23OlnR2KMdBUdeRNzy
iyPVhrtAQ/YHNyODTKRJOs/wQ0ypWdExlSZN/UFZduQmu6H22b2a5CnOpesc
rrus2G6W3TXPh6az6q/SqLHr1HAlPmeOoo983SAWADOxR26gg8mP1W+Q7nZU
o3w3cNMT860SM44n+0o1K5tGAis4FbAzItk+/EWr6I8EPNKXdRM9K9k95vlV
fp7iVB031Lpd/IQAw5uxrrwqaTJe+SfM8BmKBgoE/ev5pG0c2nKpJO9xG4g1
u2mnLd5sfgXmMesecWxjvf+F3xpQFaTi/3ey1rFeQnINBf3N7xq2tKE7JfT5
qYDUive1VV+EsoXv3PHrzlcB4u0pLyPHxE2tqaW+wr0PqZZ7KV3GkPnlKaKi
vZHn1Pv3Qso9ev16/Lll0uN6eDMRhXankM8/lR7en4xO/GKOqDhIMGKi/zxl
sOP2FjbFCN/xdWi5seMGH9bnaHKu1yQfIARVS0rYKkuLJB437wHMsEEF48b2
cdZdG0IDM4V7JA2HpG5TxyPEVke6qi/2zj0A5vK8idTlKRkcLVhZehIeymmV
fUH4nKo9i7Ar75CO+eEyycV4A18a7dO6A7eC7Gb7Vf0pezyVn4zheKLs2izd
Tpjq+7+F1juYD59zOi9343CVERERdavzDECUGpI2Ia/QNHxf2m/fYzk9FjLz
zLDP2LbU55RVf95yhigmlhBiQNfzd477ouruJfDb8OamyYy64IzqnCZQ2Vqm
4ZkindUX6N0frRZnwa8EQdaoSuRD2iWVeF8OuXhePNZLB2ErS1MN9FGv1hDL
frOHLzUMTcXuW6ZaxGAccfW27UsgTykj/EMpBfE3+QRcD2YG8yQOD8GBQ/M1
fxVfazW6pZ6AcO9LAmo08v9PudiAW8hltvJurdjrhrtPTMcc6TovbxGgh5x2
Y+ese2a/L1qF9IJnzsc91smBvZWkw2qPxrs/Nez1rqh/L+d18IS8L5xXn364
ktQjif0Ilf5uYCpYL2MyXMmpiZ6+/tS3nhJIZ5x9q88fPxb8KfINR5rVNGAa
IqNB9Y5uWKyD1kMpJ0yA2EEcKj0MAV+5VsNQY5jAQga7A8jHstNFFuYCk0kL
hzcn0AsJaan9uS18aKdqQr796GIHnwvl7jamOZ15fgw/hBlN3lLdRvK1DSUc
sDe3V7XWoqaRlLNhZfay3JPPQ2Z3FEZT38ky7CRKPLJioa8iynqVJhpm8H4s
KKyUVAMWvglkRvJfmm+Shp4xtdVbWvcX4sTOdOQ4QPwZie3AHpnCd0RWr02k
befE8Kr7PlUlKqGOqCI7swbn5h/wy/GdRnh/JsA/akAK9848WF5/v8hcHaqu
WVMOvdeCy+Lp3AeJ7f3iKALCL8NeJk/MAke6UAK4PmbHOlfiodz5M6Sl45lc
7XWNYevwc0styOg+LVuLR4GJ/ihzcznCPrNwUzzficKLx2B1gp0bZHqYosXp
2Bd5lSveLUj+4tRmnpIx9gwlMjdVB3S6zKpZYULPWEHQSKKhUy4q8jfghotM
4JMu2e5JbnUhYpSZ8JThxLYD5AlRUuMY07MjHidfUZRES9wf4Il/VMZCtfVs
B3JguwfiDATydYtijm9mg45tOxJCznW/m8yd7z59MYzQVg7gEpjw1fM9elu7
JrCTaoRzn7ZW386yn8kKF5NawBZUOsluHK9c9QdYLrNjAt0RIMXfV1srQsqT
LPPaaE0fo/7gnF1QIY4hWLSbxx0z3C/56ak4+HQ5YE4gsK9HhrXlCryRd8hb
VWI12y8QxIRbfH7yOnF2uTQHQ5L15EhmyARbnPILP24o6QLNRUGmJrDfP8CY
z+jNzkNfAydS3tElDH2WchcgmmhTox5Az1mVzqLcM+cOTU17AyN2o3koStS1
27bZU6d+gpu3bo7cOdUP14ldSBLs8hMmFSa2FJbiOa2qpFgkbIroo/+Az2OQ
S+LcWmdgUq75ZXxOoSKpSUdEIE/mkAUe/acSG5l7w0artzs5PUgj8ssaZ+bv
K0XbKsYZviUdtZWOI9M/iR6mAh7OiJCSLDP4GWE7naDR27GoZD/aRISnScwM
LHdo78aMkZ70UQ93+V+v/wPWX3j75wnHoc3Cf8bY+CfPHfLZ7yjXyT2CjGkY
iac17yFnXyYRRrPDvl2fn30mLO+hNJDFiMnweolUhNoW0AQ+f/CZQOOE2sJf
m2FttdGke4cmaym0zSv2Mw3ibJQZBtlnYs1bwJ/qbgDxHZstx9H4TiKifM5s
NdRTGfxh+twNJSqXFAXP+tbilheDPFra/PQ1fct8RFvrMrn3RBtVLgQ1GIuU
E2EQU3bR1ap96bobJ51SNh4q0dr76C1vjyGOChK2pPlCW0B8ISpNBoETjhOX
E+sziI/lIUC9pLJrTBsG+HGA/l3MNLButS4FPkjXbOSNSAEpsQAVR4DJX3oo
nMn9dtwW37nmTIcC7WF0dvOI3rJzpmdxHwl06BD+jhLkLw8qlaSXxV0MgUgR
kdzUwdDCKs3/izwPxtTI43p4D3tdHyOsDzgLoKUnRli+V4OzC8rO742vwdkD
CzP5SNU2u+WrwOXK6QhVV6Og+A9Lo+qvBogMZ8xY/I4vLsBNpVe/DPquFBd4
7kUYxzze7Fj5GRA0S4uPCj0IDDRc/dLcbAMBSZ4n9H+dFd04MFXGJ+CNprMg
mjNuzqMdWIa1OnTyLqRovsvX2JU4ig+2nOX1hSvxT7J3jVVYU1DkC0HMANsT
F8xCCEifaj8b+19t3Wn6vbKyWpMkIN2Pw5ns4lGbliyzbHrtEndjs9itHgwM
0j2WZrz/wjVmHJZAEkPw+u7yDO3Mzlgl0ggHXrBLKuQn5fhT6U09+zr1YKw9
dsj6a9HBfS1sEYFkWPonwkgc48xbujxDiMoUqBG+ud1LGVCSVrsxYuFlnlb9
b2mRuI9Z2tzyhZ15Byme6/J7vyLSQ0jFQUbc2bHvJJEqW/w/b90/RsrYcjsv
D7zKiUlvcPFULI1xmRPEVU10xkmGEowqaC0qDE+3521oItzwS3H/eD3cQh51
yRwAPUMo/Q1i2fMSmk8zUacZTRPXocwqDJb9bG3S6J5+8CR/skwsBukd2G9+
W5u1jF9c3KR2aVnazQ3GUUurytmAAaeA/LLruWt6aGx2kAnZ7/kgPS4vj6LW
0cclTzhHhjNbGEkhDmyh52QmjqA6uNAsIy0/dR6yre1490OsmAat+ZmmP6lj
6P0rIqAuQTHCk9j1uOhYacUyq51J5SV8VaxWfoIqlq5AjoH4lkQdyNQfO12f
bzJr/P6kfvDg7v97xF+lSmvnOsj/6C+swc/o1EiA2vSXlnBceEfkS9njjmpw
lMCu3aIj4cHbPlMH12qadtrYbF5fwolJndxw1iOsQ+ZIo9fQdFP751LASIan
LH137vWj5G+rQRunwj9NHtz85I2+I1Kb4u3c3ltWZ9sMoWDmnOsryXbWpnCO
bz9yug3Znfm1lEQIOWnd0LUn7VuzM4Cdj1fp0S9cMnfVkHR6od3QaVdcnG/L
Eu3Dw52ShXdc/jGXBTVQHIKtqAup3+7dZBzAVi01wna2JS5GqhrYPFIuYYVZ
88cfKtRoxAHSMlip6+HVgU70MgrzXuXe/Xnvrrr30VHnkqJxNUH4a5aJpy+e
pQjfy4gw1+ktIi+f4vkSGylANa19YLCIvfXL6tW5j8ikuPz9SR8AGsTUnb+5
zP3rjZSFwo7Q0c+pRLGdADFryA5hAEMMDnXbnFAaXLW7QD2GnAtoAx9zBhBr
hYSIcKU+hbtoCAk4uzB44V6cSVNf2cRJcTLEfJ5YmxucGF+8kqr46vRKa8kC
4RnJhdy9HNBAY3GrnUmnUpZ7aX5PBzLemvChmVLqVOME+KsxnM6ucwB/hXzW
1lgyNkwfXHkNKN1rOpNhRyC8E+JZrARmu3gnF3FgxMW0naS+wJqe1qdP+9Sg
iat5QVuUc3D1news8/auGSL0VwXGYoQRb/hhTM3GjNPYQniSYKufDdbi4Ra3
uzivxK8xsVlZbwwVpJ9ZzybwubM+jNzCJLJAL65f1iPqkuhGABOhjqNpghdA
Mus3bavPlzUZx4LtkFEadpdd8AjaA2dVL9R1dgz5Sp+kKRQfQeeJzXutT/lw
VjbQ3JsRu3XkKhgn1T+lUhJcwOO/1BBAWX4thsd7631vu775GI2rM/chuiBh
9FuLKMoWxg00ujIOWoLRCBEq8epx8RoS6Dqh1VQZoA+Qy1KmQgY0/IK39pni
QKvtDkb6V2fGgpK6qo71LHX8i5lKhZsmnZJtTl7vo6jAoCjOOGDJOBFiYawL
K0O1HpK3rnw6/9ZH17J8dIBCRXneZzVDMhs3o8gWU8YJX8yYnKe6xJ6Q0xXY
ZhnfiCcfFgwKjHK3LiOZ40QrZsYUzdna9WPS+QR/UkNI+k5zg1oRxoJU2N+H
NMfFBlxU5eF3gvpsH8PFOTdcio4Fc/IBKbDlc8+t74GGnlviIhTN1+C4oOFn
/hvz5TvHmyktMRW5hORH9vodXBN4dYZNKNkl1b/ZDHxSPujpQ2Ec/52HJmsk
5KoOw468ZvzFGbc6MJfNq3+YrxKuMznFPuOUVEIIV3JSiQdTzX+t04sSaVeT
FzKYCb98hjYQ4A2S1jTcIACeOy2HscGVCoznw9qzKcNsCZ3Zt9xkjcecehVZ
O8kutMJQ7E56yO1SF9v27zW0OMqXmhiVCsQed2io7g6Zaj9pI6yA7hsfr9N0
J++XYmoXDoZD1zd5ViFlK475ngHjYivA+gXUBo6ddtZ4mDO+IjW51DcDesDW
A5KyFD9q5VGqtGNsXxBOpL9nh7s7zV3mYKYmUimlne4Xs71kEYFl7eDIxwjE
/4fW6FRRnpgjLY0QgGqI7SeNLHBiSHu8bvugywNrdNagUPE0lViPigvbIuPS
9fN7+068ilqoOHifjPx5AnzxykiiWEt3AWVbRhuLaPnJwXvdXP17TMHI6SUW
QLS+yckEXm2ppuJkC9TR9aR59Ny/YwJhoVMI6J4AlMvdDOIToUg2d90JJq5b
5ni9HScARGn7rT89jk8DPzu7j5B8TOUpf2ZkIGm9GnB/SF0gXSCRieL51nXa
ETl3tFEI7FZquDFoQMLXZRQFt7Mrhife7AQ1lca8iaq2iqSJjZtOEQ4Y67kI
Hz1q6eZxvIsvrCv8+KUTpoKUCY7dGRsfBSzFy1o1pbE8GRsz1/fh6gVpef4x
/of3H77kUFzS1cdPq8Wf3sWCGTODCqldb08q/qa0nT+yHWPnnAngXmDaLkBY
jZO8PDXBVwaY4n31EgKSwe9bqZ+rx8yTAEzLOmc6JO+WAoKolGUkQvtVLyCM
uWeC80LrlmOB/80FQqjhgPJvcx+virNxcajaVPTAok+kyU0nuuITNHkno4jL
vfo6fPO2ph7i/8UJSx4kbpgiDWUQa9tbNNz1UkR5cb6EMZK5E5DPUmIU1aLJ
T6fCgb7ye5JfnifbK10vZYnpWkp+HKEyq7tV9gDBxwkyWVarVEIuhvMsUbZ3
3ROUHRzV5SipXyk96lNHBC6F0EkSG6DxyHKw2WxluVs8IlZkLt7V1Zax38uj
o5CWdhjMD4N3osLHXzNaTdjK1WQkA3Jdyv7nokq528dcU+t6HSWbCRiRMEAR
8VgQWqNHvW5XYxwlEaqGpalLdvsX7/H5EVAIxh5uadJSEmgaWPh5Y2ZFT2Et
Q7mq4jSEGlhmce5/UBE2k4jtWKivVmG8XOni/0iOTc3flyhLz+qkD3ryIZ8r
7uJCasQMBHLrz2AMVGIMfEb4grHpkFpCiw4hhAu0cq3WSpb7Z6uXPj7Pxfxi
tyAJoDFRAJlLMut03V8wDPC5DJzpLpfSRF8zZhF574APWRzwndUUJqeb0X2P
bYGUSJJWde4/KnyMFLAfAjUbjh1BwkqDHjVyYZRUxc0Ji6DvtrxmLJVES65K
4MdfdtiH51IeBBQ/UD34XD+/SW22lav5o3UZ6OTzzXhz+b3Pt4NyiTEJlpbb
LPJhCG4c/Tb/pknSSI4wH3p7dFG1YMvlsbfk8A8sdEcprxDQc8LlphSbHT2F
XcRFgUn9ssYeEGgPNKcfhqfv5sO/Fs1MMeHe2JdkcVIotnWgPLvtMHgFX89T
dlM9XS7tKbx/U9M5zc7UgkXiFvbGhq64WxGLWLzihBVzVqzagApspguRls9m
XeMa/f8A72Rare7DZFFXssnmzxJwGTdpBpzWBIZwO1+nL/h3UaM7ZeUGkb55
e51RMsfCfuZsKCiw1B0ugg5DNNXdiUETsXHe93ew01iEGEsLlolomavg83x5
Wx1O2hDpMrbXeH424GrwA/q1BcRuz8BFTRndzwm/G+bib7QyIb/nSY5iym61
sIBqcuIIQKqiQvDg6fo24zQHZ+Z1jyweDz1f0pvSiPx1MnZwawrcR2iUWCmF
5/vrC6gV8f88okhXsqoOzLvz2HXQRO6sr88kGDpXzA5FiPZslNBnxx/OXeEI
1tBIP3Fvw5WbdtfNr4VUOIanRdXSKu9fwDmxXg1vS9vrRT2pRbB0mfqQo5l9
SPJAQk+sSWgyXckEO0Vy1Ss1prGSbwsjh3em3ffczjWNwbwPyywyAtuIh/jk
nrQeJVMRRbWVYEBPZyuDGNiltW0729oaii0+ZfCwv21YOlteCQmlc7HvAjXq
L1tofJCmE/tt4G9IKOPA4Df66GQFPiBe/RI4W9SrJIQKQFAvzU05mh0EgZuT
lFPEx4zpk06vl7o0gEnDzTrWz+he3eMtZTUMMjzOD3TVNff8CZgsM1cg4XBP
UKZw2K/jBWrLVylGvNLCIqtWYrKOIagYCz8awE1bH5e+pPh5ONMa1OHvJa+G
5YxWxF5TavEG7aBQEzI5W4RoFkd9LNBFsoqIbO+qFfuHKzspQwOoL33NqzEp
Vuq6kNtpSiy8s5c02aS5mjKSduoHyILke5LS9IOGj0WPUGJ+Vtv9tn84InnT
fK+IgKHJ0CM/+ypc2x4KswZ7MJJAwfIzwnt55gUMt6RY+rTUZgcC2sOVhQtf
xTapennW1bBEZ9b+K8rP0KhlTXj2T6xZgBo1PXTLyiVCGg/GO9rrTthN3hD9
cnPEAYaGUJajxd10Eir1Jk2e0ev+3drs02+fkPujPUajTiy8b6a/cKqp6CQp
5gnJx4zxPojVCtH2LPuwCImyfz13jp+FZp5vV3HFW7209+TRND02cPs4OwNO
cKImdYdCTkw3d0xtvm0sdJthZATmro4Zvz3orwhPf4S0XWoM3aVqRBg6LrHm
IAqXKoa4DGSUWMJyfqkrxkzhL2S8kqeNb3Ffw5pnqZdax3H7agd2NfO96si1
3MNbzWlj/JRbV7IW5+/tfncrsUt4M1LEjK2EsRh1w4VdEuvFat/fES1l/QVH
2+M7BWXIEyGdwNN/iN6f/My7sSno1Y+m4Ho5/gy9nZStX+b7R+TcyUA2MWiW
U5MUEp3b9nZnmjXe79UHbrUwwhAbuze85udRsteRx4VX9+IVyJWd4I0O1QYk
y3WM/zE+KhTolJsXzCGsbhrXC9P2PneRPsUMsEOp0vzvRWuQQ+kWQPvzx/WT
SUf7WE60unvU9QHtEVUf+xzf39Hq5JvgfDLpPwqMVmIhv1fivQiSG35DI5aB
vN8ti5xh/GGysHNb7RAJHe/ie+vSnVYVXG6wJPIVQECumheTKWOAKFNOaB3e
1OGLvKyKyDkbCkh34rTmtT84afNBO1HVSQHc5lNc4Jam8PoQ/0ygclFZemWE
HEaYIFtrJJR/GXjPQ8hFRrM0wowbAufAK2ooOX30W85SvWpTeGJC2e4SSB1R
h0D8mBzUAO0nNIDwYLv9TdTeBazaSGi1dMoHLTz3Ww0JSakDIPyrv2p7ljIw
YwzsUcfRjWYDNcJnphAL6QcDvq4QcS80r3Dv8H4uaZafhpiKSPjJBt5Ar0pi
XQ9vgvIkMYS4ej0GoNlV+lmXoUSSG0z5mjjh8scQELmpjwXJrFyIkX9b/SiY
oxmkUnIzzo/35hMeJmx3c448wSfXw/4Oq5dQVZF+3sKxWSJn/AaX+hs+sQta
C4+a7dN2OM06J6t9+p4zTHdxb3607viELh5D0hn9hQ4DZgu1onBBz9a6v5Nf
BNzeP7tYXn9LjZcCP14e6gofKFbld6BdfubSbhB8fc9y8L9F+JYGTSANv7R+
HXRyhxwniyYw5nyaVe1GOA1t1tEMTUjRAKvt9NSeen7GFjHoTvXxomjp4wNj
qEfxxvdkllPv4mLWkRKAZ0ksTKvApumdYQVU2tnAyYIdpd8u6+CgDNBbA/zx
TjuQh8+MZfRzzMqyVbMpBbjVqATkHxKrnqr81hksU/urWYCXP/JVGc8p2yhh
jgx3oep1k7clNWFkUx3GpYp5+VX2F74upshMktZbluisJJ6ZVWFeG6zYNwgz
rDkqKsuiXVSpQf9AjQUOa9O1/gup7TRvz9oZNqasbqqD12++VSJpt1ni/yCc
M3lk6Wcl00iRdkUa44KKur0ikd3cuzkBYWCRTfKWqN83Yj7UOv/F6zfyfDzq
HsFprqebkIVDvUG/eA0SFVHE6xEY37UFZlebwBWcpEajGxYFcJGucQjMAPnu
D4cUYIBTxNomPQOzP23fvKcaF2OU0sKcZeEYUpxSguctPrid7p/fLe9cwijf
sgaENCF2R5+7YZ1OalRlHF1O+Jse+Of3CgBr9WXKUZgH9D/uZbVJ/rAkFSUs
G0wAEPz+SoAnJlwP5cgBfzmxd77Pex1idyGRgRfyShqbjp3RyHqLE55x9rq/
61xtngTSW2wFmrwvqEgRYkob445D7qZH31h2Ar8NDGcTNgESupb31XKwZDZC
Ylxcw0rdkCpPR64oF12ThKo9qk0HdFuBkW6zv4sKfbBdusqJTGzWMTduyMVD
nEh0wXuB20AfHgRBjkA4OXaZupNl8UlO6tsQJYvTtM7srzqVVQmfi+eDGt3g
KGpWIQmxDjVnB03aKMsDiHQ7u1jOJiLHeMl/XCmIgkO+5Oarn9PZLh59YwVv
YqcRgI4FFVum3TbMONK17sOD/RppOKg3FgIGEuU125GVrdFAPe07r1ai6/cm
ijcfYdOg1gF1CnEUveE8wV4YVbe37/4NgkMeZzEIMaBfyIANKW6GQSfWugS7
toqz+dUCSBImMARYIwnPvqmKU4YXmvoeEGVsan2n1F2dhbHsKeGq8hGojC1c
4tCuhqcsopJNC2C0wBK/E5hNZH7n4WC129zthOEWfErKzV3OcB8jkP+A9g8c
xU9fn+kBQ6Un6rEW/L+Eygzd8JE2jm6F0ndoJjz2KpvJj9SGfiW70DTXwNrs
ewJNXrHmYm+cB+h0x1Dn6zVpnQQ8cpVJ9MMVPDIF6Xno7dpjYoT/l19inMM5
iCC1ySCNHmQnDaiCKAWEX5n43WeCjwVun+aYLv7CJpLYH7twoFeLzplHq1BG
1jfFiIyieWdN7Zwab+NUe7yPxdmCcwBZhwdUlV/ao6CE58NqKCFz3B6m/4YW
VnJbo9szjTZXClljXtTqRRFZY6aOb/8XshujDmAh0qaMPAMmhKGIonnTnlgU
WHgtwzswbqvo4MJzO0MvugPC7tcWR9eA8TU+oP/VNTPBU9YMXhdxi+pPoEBH
sOK6HFt4Xvv7YLLnosc8sHBQ8UJtgXzuC3R5kySeq3+dVYfeRh5HjoZ79s6o
M4SnrBWJ08vUfk/IDeU41A8KTUnXkjwexz4ZL+tLD4SajAaaSwrHp1atduOS
xdnNt58lhDx9HdyXWTkoQl8C53au+77RdmUk8ma4XAeFLiQ6GV4FTVpMhG6W
AP+lrTH47i3/rU0pDF/zhjvuxbrTrY4B3V6TWU6fnY4RH2qf44LQaCeQztL8
Unf3o6CaTx2mwHxRk4byGOuIlyMYWm9uWi683Q9JXdrkdKFcyq2mSGkcN5FL
93jO0bM9LgIqfo7stcsriKqiZZO3PpUPLlTssYXkbt4pk/F3hCqXzGNIcZjY
drrrVniGf0B7dITBZnQ5vDYdhtv3Vk6utYdI28EUBlnAa8obEgr5uNvaOT0u
k0wh2HTe6qF45EOshUxbAnIoBi4jW5dx8/qq+aI0GYwS1VLISEmSVxh8mnHf
X6ZeLwRVLKB6HDIjMYTIvNnjnXT5JnRxvoVtJDOypDfQ4i0Xly97vc32BvP9
HCTLhKQZyLGy11kdcR0165xlnUYNbvKY3rO4L1E0K9c1wwbztKTQZ845mSJF
d1m/PrqoxAGqAWZHZkAZ2gGJa6Zi8JVyx+IHV6AlnIo4xDn4jcCSxzN2KaV6
sesyOhz1C6/4GugsmU8SbyUNETqUGAh9zoh7zfDdGiQ+YCJZVXFxu8wG606u
uFmnaju4N2/bduyXurzfjzxiD5F4bFxq4K7+GQzPdpmSRjSLePf5KhQWQiqV
2XK1LXcqZKm8bQ/Pq0gQBT1o1oUyQMNoNwly/qt/U3P4F/5aFkSxBnVnQA3F
XTyRfe0dea3wFOs4c9ti1FIORBpysGM3S+08qUGra0Fk+zgT8eFxM0RA7YXP
lVx79qzKYGzW2oKiUT7LTl4YBXv+8838GPGw9qkitYcaGhjIIUFIlXYJcvAj
QRRU1jA6Vc5biWH+ds7ThA1y41lL8+mBLNRl9A3GH46QZn2B0pLtcv1/gtKQ
IT4TwvJNqn6KueJhoJl2iy/hOBkL94pOu1AfUhme2JK5FQbQlhrBvqae8wSN
3NiXzfVtYfiZ6wwxDdbzyRJ2v/BcVTPnqbCk7Ub+7xh1f2RDp7p2A3TL5/F8
KkO7AfPqgAObsPw+Ddfe7255LI7iH2XU3+NaisFQ1bJ+mz4giwuBx2yGWA6A
mRe1lLHA5gitdXRXsXRjeyeJZWn5Gugmt6GOuFWn0a803LHTTSZh5xWH6zOz
UVxUGnODFfB8LodteJgKb1GakeNiA5jYZRuQAE4HOj/eT+VOd6nZL/LqSZHS
JTSEfmp2/vVbUkJp65uNIcHe+nwsHk5FL4Sgtcx+WKL/G7NRqBQhDiA6OVHn
xoavdW1TWGY4BCU1Hq7i9yObjn09pKDfFeRdBodfiHbda22q41OSqxabmBNg
R8i9D8op+Fu1C+mtOFBcsOGAHmY9ymsDCR7OBLrmP144Y2scQOoH4ClYXrdz
qypKFcenvHZBfQsAj6yPgmNRjsMPiQWTmcKE7EcPxx8Xx6506Gf07RlkM/NB
5SU4JwwP1WKJv1JcR6NynEvqrTLRhb4doK3b7pSx+QoBnHdzpvS2soenttng
FBN9fo7zuZ+YDDbj8LPHKmL8q86JmHh7HcyNhBpYWq8RaKj/cRx3VMebKBYv
YuZvQCXPNDwsrP3+Iaogh4ct0J+0ngIzJBtzKb9Hnd1lhZnkq3e7SOnAMP4M
1b7Lub2qfoeLOQej2OG/p0WCjHKmQPd6EL90hf7vk4DqEFzC3aok3LRHO/ac
1H7AhpW/zFZ9NxoMTR+bIB+YbWrS47S8wSraBVt9i8pnrysUTYmn2gUBo8rl
y8Ot7ZmKYzafsjCLXNn3bTJECQ0AXr4WkNHbNONJimuJyA8+n2kScNawZquQ
NmDkB/rhbvPe2LYhDwMkDOoHUZ7U6xOkfRsCvxEm/g82avlAm/WPw7WazOmN
c/+iKBcMfd/x+vuR+AZu2mlk3uSX5czC1UwxMc+f4lSKMCEFII9YKe037ffy
IppXeLW7PRZ2gML9UNvAAp9/qnrRZaQ2bogEUQdf0z1a6tT68hqVPL9NSWXO
Ema3+DLZFuC47+C/7QSWJwnQ6lA1jdHebSK4TQNYt7DEj/EaYwF4afQLxsZ+
WHKPKsc00AWXZmA+0d5nLj5uHwhx6waJyNprjAYE/Ot7eCmTh0Gru5lBQzyG
rHXZgbjRJVOMSHQzBAd8XWHhC8mVielAovDP+l7eRVEt7qo1+CPv+suVtUrS
/XaAL28y2CTZoTRQOfUUj0QzQeXfDsw/DtCfj+NHSXvEQp1BmbIkOa0zrp3l
pYl4/wId4P9KPHcLKL/l49/gJDqR+otkCGKFl8+P4+TaPfNHyLpTkJW8GHd0
vbdoicaynedqDgNa9nbQW1vW97W7ddzYvF5WAv3Bj13/xz2eqUZjG29Wo6wV
CMUCYlCc4qVqg8BrgfSzu+UN+orNkaBneJ2upjWlRxyjffUK5s22EZZ5Hdp1
/cb/tddy5KhCB7f2C1p3crhH47vRvlKL3kjC1n94X2MY+BjOPz5coJTqnTAr
SOM1NKuUxHAvSclm2C+JjJirU2I1twkIf4b672DygjSJSRQzTsxBwO6iBf7Z
KHCenfPbTl953j12dvvMWAD4JkOp7mqMC1xnVW/uxJF8kRxbIIRHXDKAwApZ
hbo+VoQWMXzVors2Uz3G6en93hT86AJObkpCt7SqCZkPRMKcz91IL3QOn4Em
VQV38+aqj9QE69Mj8a75k2Rd6fonIiuvDFdtet+T87Fd+fJkugfnZQ4dcklQ
ha591YoD+2rHpGnmcbTVOsANdSS0alT8CCdfmE+xb7XNUsak8TugbaPPQ1lG
TI5RXUrzHYEL2DNoz/+Bn427r8Da11xaBbc97dfciibNc0qc12v6tR3DUFC/
Wgqy5v8CDnMioeN8gMxwLzvHN5VOVRFKudRaYdDpodReupBiHsmQAtk/hJet
UzNJY3VJVXgaG2nPnemWoi/XZ1sF3QPXQ5IPG/KrHtP9lt2S972WRYys1WrN
n+vNhjltyLXdjivWCv2T5a5LCyVaXd5A+r18qRP5cPzVJcjj+U9x2w6YPwg0
gRWv1+7y1yvx3eVhcM52fzYtjAUL1wY+m2elFAvNCvDbbAyLslt4V5leFWGF
T6ob99Epdl4/TVFQKWOQP2jnxWlBmI7q0PLz7kx3c6ybQB+3E12bu0UQcnKt
Kk7SKINtOhk6dZeG62OmHlLt8ulAGCCc+SarLsJL1w+RKLOrK/oFEOILcxLB
8Qghuefvl/ZZ3Imak3INnLhNzqf/6APEiqqtAWFWwKt5Twisho309Ylj2+an
nvQfhpHiir3bd/4TowUWDZAHSqY+s+5Q6Gb/3SA9LFt+hsfN7ROCzMWIfImA
7cNyX+uAl+UH+nsYzdlw/nnwWQRyTpV4n38vSZHQn5gomCJCULm/ACeOuXVs
VO1XdRerZ1w5FQqCRnEj04FqLg+daxpn/qsh1/KCP1z8ZLRIXaKxk5nkAB4i
1xVXPe7EbaP/wByMkS3ENh8I4W7PkE2AjRwpwO4sE7Pc6zT1VqK/TVAY3AzH
qvwbW+TotUwzzZrJhCT4irWVyJzyaj7mYdLWikL578p6zEYLj04+P/bP5XnE
1O/AAmpSkrnwBujVhrzxP0rUHoE0iJW5b/L2tf4u5/KyvDw/fsjMiY3tv5Ij
b361CPw8cBcR/JXWCuXxpSJzyX4i0SAsKHeIHQUAyqZBG9FmmRaV/dNODRSF
R/wOMvr4LBX1retIEow58XH0xNr2Y6SXW7B6sUJ9btbWkqGr31qLqaFXfZyb
AEXvQgO4Kw8EgD8OmQlLup5gzSzgelsPa0m5WfBJqYvfcZntcTLhA/VVeqYW
Mz5H1xaNMRLCSzQ3AFUQLhHFEcSlOH8euiYlGxS4gMK7Wo0Adv88XQHbIV4k
gA/3wPmGecp/VhM+lWQil28K4/FsahXWXAm9SQGXiE0Y99ETS5dS1tF3oyOw
Rs6T8fBlOPdmV+PvMMrjIakxml8Lz5MMHusaEYZoDfR8dQI29uMnP+CM6ndE
NvcO1bHJyQ9ckznbJ5/Nl31L3f5jiinTV4QkRDmqgUy+gVs6GaNHsnMgePmX
WVBzTX0xoit6sZEC49jzy56e6VlV8FjJ19OvLK8EpF1/z+OEFJ/XsGqXkA2o
UVJnYPNqBfEjiYjCD6tsPpKuqTCllxUzSruaIIIcp5/d48WPzz/zIUDesWGu
9iMAGM4K+GL1pKWZsRD9bCIXSnVRo2Y6vF7OubIdJ6l5uFFSg7ZLMCeSkRF2
55fTCCqr8cUJPckNkkmVEna/5MPjxRwL7y/MhLoNxbAvlxLklxOC5Sfw6pyn
TnCiXUXSCuFMV0yZwiL558VNdaN+tZD7CRRsVVY3toEehslha6mhRWlmgi4n
h+RtZjX6HxTD8EWB6q2gVaWeMCq+oEMDIyr1G5oaRTqDWMlNQE17s5Ml1MbI
FHPwKR5rgb7LP3lfNpyC1rVZnnpx+lndx2k8zQKNAsSG3Bq6RHyuPXw5s6Dp
ULv4Y6bKkMknm+YeA2rAiS0YjlLfpdenwXF/yaq4uAq7TdF7e46ZpDLyT9ae
pW8n0e5iwDd0VhSeUqGbdfLOuGTUiHy+3fnrrmyzV1cZnBvX2ViE0ISLZ9Vc
qXd3WDZBRah4wLZF/JKuwlin6TBSxiIPHutdAyvznno7fKcUdp6Dz/vdDAwG
YJdOKvczbWc/t3oXU4EJA5D4WWeHnjazbOe0BuNnQqan7KJRd0WpG4g4DlgM
BRBka9XyrR0tDlppGTSLY8rBvSXO6C7GcODMscGikOhjMEoYmlWyMHq4UM6T
YLf+j7ldDuwVagtHmtC72YK5haRFwH9BN8yEijPQ6OPB7oS+3tbk/P19ne78
vPLUdQPQJmFKxbeJ+1GPmp3wEzXFO1/7lRdPJU51mqrUZwcH6Kyf0Zd3bWNN
Jv9o33U5CwmpaSxjABwco6f75oE9SkvhD9yjlb7P1wXOEB2X33rncCkTBjZR
aaiCpblYgsrdnstbgsUpSysqbzlcsamJCK0zEPUpHrgeVlWKZw8FBe6DPDc6
LG899q+serC1ESiwTUG0YmBjcGMVPRICGzCj2ueijkf4t6LwoykBiXpESTzT
gjxQDkzXIbAeaSbz6fZtxF6YSZohJ8FAsJLCEk0XTPe07r41sCiO82SNyNbW
hM36wsBBhw4BJVqGoj+YzOWFlBMkBuQAH2QP499OPBEK3DKlddiEFZOA990/
80RpMjLBx9MzaT3j06Q8hfrVQVHNceyVHQkssusAnHm4zzSPSHBExNXH5/xh
pB2GTKVmFD3SpHrst5DSiVwbD2JlsRsZRoZmw6KCcQyLCLZCbOoQ/1AiQaVT
t0mlj9GhX0/smOgtv8GVbrKzH8C1D9az6xv/eqWTCrZltzeafeDAFsVUHySW
XHWhUQn2pQQwvUL8d9dXyLt5hE74e9iwL4NHNHYWj6NhRiPnYS0EqOleYgKX
qrCY3rjjOOWQJsjNQ/enWqkyqFnVrpjJ/OdGPxCwU+4ZHKkX24f5bSqzk3SM
sq4h05agZjxcXsTOYIPyKFb15GDd628WU7+VIUyCZDLAF6gIwP8N0GBSIPo/
NvfW1nU3QXFG0dIICCThl6Spx7Rl83Ki0CPPvdgfsmd354hQdO3c032lREpI
UrFOzu39IFDVYdoJhHp3UsqlVrXmJkHvePPg8OCVeMmDCaySpmBb8CzDHVs/
shnDqebtO6p4f06wuZbN67Lj2SChN0umAoKOCCNVKCpJmDJjcE8wahm9qu1O
4XPplf3A3pzC7LFNGghQ6BQ7J4tBvY1jK1edlGVRbVJTog4fSCN2Vk46nW99
PC6aSxtharWiCfsx8qwLfYmIV6jNU4SK8uLMV/evIhhBQi/WZ0T6ccbCKlIE
KeYfm2LPqWGf01TLKu+bx4IWjNyCd8y/it2Ysy+uT1RT6ICWj08cf6KqL9cz
dNJXI+Ci0an+pM5TGo6S9dfUkuw15GC+41IfPTRYIphYeF1tp2+dDCsHtgOk
XaPjiJrUCT5RL2DEywDGWulyos87QgM+HeuocguEhR4Rp4cS+5axvpnRlWxc
z8qoWWE+SRR3y693HCHxco5aU/mxzx90DMkE3g1QlSQZk4AJ7NxpLuMOo4tB
mTGBKGA4Ccvs+cXnitanyihuOFY1CVd30fYJ6YknkAUkkhk2YGpWROn8E+PE
1q1SucCPIVOHFkE01lgdyEezyrDIqSlMOnWKkdAKj49ZJoduFs9rVAHmJUUy
69S7/psl0X2Jqe4S++aIHMCuye7snvc3MIGZ5YB7ple2Vok+lVzppFAIrmCp
7LlvwS5en6jDnxfapB4V41wORRPfdq/YoUrSEYmKBoXJzcV92fwykG82dgB5
c/5Zerw9ERLBI7yHS2ue/Xq+xR7fMUEpdgnQf28Voa8qPD9ukA/uFYX3BAji
tvHa+QWCEHl7vJ1wx+lHenN/syNAkIEMRW7NYXwoW5UgG4Bja16DPgKV8vIu
/iybWJ1mLg9PRNh7XQ/bwDod9oNNa3Nt7niK66DVZV/QfCct1p5UHd0E5l1O
nkBCQx2OmHZu3K/k07k1bAubMecSQXmggY0ZoU54VtmbVdjeAuGZ/G8WvRFr
m/2qCH+/URRvHCwmKaLLoGKIk4nbkf22IKaMnU75SVtq1nUaRyAeqJd6yyEu
potqdjTekxWt+ud3+4BRa/IHIdf7uKwycjUtEIowk+asp3aukIe1408c3d1I
3oa/YFiaM9SgxXhcHOBbf2PMx+nozrWYmZEu1xH7RNkwMpTXYBX5ZdRLRGF4
YG0m1zFfRjr8t6VpDVmf+fNIRNmKEXdOWb4Amj73+j8Cu+mF31fiJHVn6CbG
IuyDjXVGMuD5rb1Yrc3+t6OWeCkhVGkvnXml1eqVlJvBXicE5oLln5Y3e31j
sLK7aEkIBAG4orlrd1eAV2yyOcG0TCh+WERWhefhZaiI16boZFi+JEZsTWG7
lkDZriHFNsBMVDaqcFFTGh/6e4pbxgOVpnFcztu81G0Qe39keFk7ILmd/lar
FjNUTcVvRu/MsGcYD4NgDaGko0cqEH/NCLwX8lsLGyCV0IaXbp5KahBPnJw8
fZm5o3yIKnb0TuNNOkmJRcfDx+DFqf6SxoODOZQkqcO1ZBhuZ3c2Z6QTPbgz
QCdlNmD5r0I1JTk8AvBam6g6cBn2M3ooN/DbK0zCSS7FpkcX2YxLBa3dWjaU
Wu+rdCwrALy6cvT8nYNsKyVQ/bBmTYir7lf9YL/abpqz+B6m5ezNgMQ/7UI8
1cgOJXmdwsYqaJ0R1gzK7GOgxH8jUw+CmgmPxNcd4fA5xWUW/WirdZ7Wx2Md
NrMFW5Zlspx9SiXRSYrpiQao0o6QGAwD4Vn9F5eQBSDtd+1mDyA7U6lSlKgG
cTQ0r6b6tOp43y1QKlSIBuk2MHW7y3A0eAbI83WJc+hTgzT0bZ4xpYMiq+5+
WXDuyZeXa+Lo7lEWb3bwiXuYq9Dka6oJ5Z38WIQgojelNUaoqSzuzLZsuagK
nNjTJccXY6r1QBy0I/FgpMB6GGljaTK4XH0sfIIzk9JqkTTEgS6pl9bD6f5+
93dFdAaqPxEFu6u6o9xZGh5ZJf0xB4p2xcy83bOri/kQUNw8u9h6xlWNdghY
U+05G+eb6j1aRvYFiZuBrICGSv3RKjJ5x8JfqSP/11mQ9i2Of9RXHYI6Ogw8
blNnEKYfnktpgu4nquo7UtVSHEKKlG0+Py90Heiz56ugUJE8K9DWgOMOf00F
FYswbtP91zXpYTUhVtupW1AwTPaoXxTJV6C2F55zg4x7iFDui4r4N4edVN33
/H/ThJd6oB9y9TGne3+dfeSw9NrGcTngLrtdp9E1RdQkBC+OdZfFygaX4xlg
vH2+Ma1bSUForBoJmSF6Av4MOTSVH8YrBbdCY8qCXxsIywYlWZv727qHToqp
6m8rBNSsgWOIYzbzFO1+/KH7CC32iPm8HG9AOkFMVb9j+Pc/S6b3JNnYSz2V
t2+gUum9uHyrkstgr8gQdO7mKEAlQm3RabtZkhZeveYiuHn4RMiILJuln+EL
0Q4NgyTCWmjDEpvl21I5HQN1/04Xa7KEI/qDuRmLkbcwBDgYbhiPr7hj+Qmi
JnVpYAJI+EnTzSPRer0BtUDAWGheaUSZmJ1WsLoVh2swE99BIxo7H6yMgu6e
1XpXGy2Mr3gDY/nsunBUuyprN4xPw+m9UMNoYA9IVltAstc6g58ulCzMrIGL
ceDMu+sBMOyQlzGi1eoGjUsT5u0Eake99sJvQFywDgAFYT4y9eNoncPkb9ak
aH75IO7Ay53iY9T3KRm1M+En0bSLCKU0Hz7I4f1z0grVICjIN8ETBwQmuRTr
YlhQZFB3xDLeZKV8n3M23PJnpeLIfj8wuhMcnIL1mtA8XQX9hzjZXDOqR74Q
xv8F5fMj4T+eFIGbsw5MPo6mE1SV9SJoNFb+k02LVYjJXjPZCdPQZw8LKqtd
U4f0TEWbjILZfsJZwJ0HJ+hJFKR1WPIDEPOUP1umLdh3qbmeXjC+HZtb6RJb
B8RLdgppdy3dTSxrp3/Y7KQCNjCzKLGM5QVIX8JP0Cj2bTp/8o1+WSf/blRb
BwqGcWitEHE9tindphcnm8i0ryFfYUSQfxm+adAeO379+1BIjwwRu1S6U+R2
lZaPSZjSn1kPTg6N0BxBOw4CwFJgjA/JR3sZSMX3QP53tjpZe31BSPd8+FfX
1E+pt0uB0vOY/m/VqbzKfmXjM553lL2zVZlN4GUj0ANlVKMQuAHk69+HkX9i
CxgxOQbc+X7Fb3zsvBv0XB9T6BlA8rH47TM/MHn9qtfmKsX/AzN4dFAZYrqc
8vViUmBIe5TuvOtNaAu0LjLI4Z6GcaQgO4tluwhpNG9AVMDuNAaNfr5Dm4XY
ntIrzWYiGcEXvJl54aLvsRb8zcduMTk8UU75b16w3BFBHd78nelIbW9op/Mg
lGAU/PhqhH5X3OlCPd4yJKf/jelInCLXDvuD1Eovf9MRf1iCe+O1Jf8hbsup
8uqJdf5FI6Y6EMFdTgJ/Kg+iiofSmZyTn+ld3A5592TQfc1AVid2U3Yngnhb
fciQsE3LheKieNl64HBVEjs4w2cONrEIXlseBhuGW3IVs/WDLqCnPvw1T8Pl
G4SASZZe/OnkpvpmRxWUvt5F6wcNwN/HgDcpfImAchvuAQYpvFIOSzbX2txk
JvZtJXPK59/gQw478TYKcuvhbuYFiKm77Gl/v6ezZeZPYIc2x0BSu2K/Xt3s
9RuUE9IwmjEm3jYI4DVyiveeCu2HOL90KoiOjw1AOznLQrb0sn8LhlGK9BDC
r1MAdbYblo7Em5wuR0UQYGUJX3dMhUo9kIgUFxNvkSv/WYg+BXNCcdXvlzCx
8VlLE+TQfkPVyhkhWUyFtiYCnN6LZy/hqYyjhFDJw47UZbzONF/w9yzkpiFt
o3zmfnt8e5pcqmaH57VbpJ/f7yVvmjE7Qr1I7ZrHcDSPXXcPldtPJ+wUkJVw
Wls6bAxbVA9u1+AgNm4impLjDONgEN95VsEr6JwGlmobibmZcdSItXToFKZz
YO2XU0LeRijaqt/oS7Bm/Alov3SyzYSJX3Mx+n57vuw1ZsJpH+5hyPSUfxAF
S3OPRu8NMJHgomgPku4jBAv8LpJZ0zEszvuFQ3R7Y4OW+OZmc2VLZhFjEJHK
X71DNYNujhtOT0ugRPlmc+TmO4267oRM2gdC7UjmCSJil29X03Mv05fzqPbs
HeKKISBbhyqcr0ERNnWQeExEyr3ttvfdw6/ahpgl7SVgxQ2OvWCGNufko0/R
1uDHlM/jyHhjcfHU8vFs5mU+OEbOUVtSxOga6ONl2NMa00d+FeBPeNmU9eds
VLJNnhnTfP7i1uYgjZ9G2EKe0w1/ugztU3ozT8nZyHX+KPbfm0eOV0epLZIW
cBHFyzRrFwHaR3EQgjKKh0qCCq5YizT6Bv8rXTZEW4X08nJU+6n1Y6D2hZ0R
FaV8G8eHv3ysbyqj1vC0CZYt5pcZzkYKRTNBPKWJmbAMy1N0jcS8ZmD/3lsx
E7Xkz2IbUOQ2tVPZcRNxy6gdnoUJE+XZYQtxkzAdlLER37f4ocYOQM/9L/4G
iY6Ge8u2BZSnDwfAH4grAc8PH7nWWZRktP/IU7ifvaX0AUlY3WrL09Qw/wBC
RrvNtMZhCgc92m+1Z5hKEk7jylaHCASKiROnFobnZsCxxEScPzfZY94Mmyxr
/7IYLQ+EFP6s4f3nn9q2Fw0XrnAwE0Ahehw5YW9lP49ncWoxe5AelYvTBpsw
0he7h2v17qHuH/VfgRScVxnSCiLSq4y49ZAur4HSZh9+jKT/TjhCI7lWmoIw
PIBcooDXOzgD102PRTddn5w02JdA1ccpy5FPFwKl6tqCp37302U+TA3uQgfZ
wmaeZmo2e8edvayDj7zynwDqVczi6KIdv5wdHbINfhRTK5XH8FPFRCaEK6R3
o6LT+U3joKW5vRGoCaCOYigd4UzCO4FxHRHG3bkYMFe/B/12YI8J83bMuSaS
RWmVNPoPbLkp+ekcjgHAmxWo0sNmDZCvMSFARi5kAC89m/HMb8mfpPdOq0XN
Nw9/ioZbuDzXT6b1Uy1LSvEcbYUq8YMAr9XJF7gRRrOfPWs2jV/j9h2M0lCE
EUTOX4YNiMCNh0Ta5fYob/VKunGhE7Q+jhvmomobO9BZyIUcUm2PXZSYYUkn
s/QXNlLOmVv8MJjxtaiC21hq7TzhWv3694J/YbihgSWPQY8vmwlwjuDsUpLG
tSyfKXRaaNKxz+PevrqbwLq6HkB486kLneXodoge/MsA7wIL2rllyxZn1lDz
UKadlAk7W/8PcfqNqBpSys1ntkilMB4D4VnIaHXLxo76UXIZ9mSsLz5FqWcP
FRjD106kKj6Qz5IoAloc6XDdy6ve7hoIWtB8pp4Ns5sFq02dLSvNlFVOav1X
L1e8s1Oc9zw9QYODo0rFrdVb34GTlsEZuR4bTZMg8JeVhWESOkjXy5NNmK0u
YeY7dtRyMa1tWm88xJQ7rjQlWjdFtYQMG2ihWEpH6/gdNwjPOUGDUfo9xGnW
gOr/tsaIud9NlWEfHDfuHX0kWdIzJ29ZiHZXXaP9fq43Y80K1BnuX1PIt2wC
azd+27ajCo2Sr7o6VCWGQGwQAqynyPYE5bIvbmLmMmWZZ3KGzSAmV6pl4Zl1
8qoe5HGP4GeHEfQ0lAEheYu8cKGVpx/vfnWqYJVoFYjzFGIooae0sT8ZzZoe
IJNawLm2urbH+TnOxfLbYr3H9i1m1bvI3Kd9p0Xk4ag76NXWEmF5/qAspa1y
jtDu+QN9DfgvqZH6ko7AViLYJl52RD1d25GUZ9yVk6eLETixZy0Y719BrwAN
+5NGlJlQD6z4geQljmBNmH4jJquTRXgbEK2Wsap3sUrI3lWNz7q+AC90BmqA
ryK/Na6bVjurA0UKyjPYhHjVnpqrV1WJeaZPZ/krHMtFkcZQ5i3fWDuQ0pQe
TPDmQ0+ODUyJW10O92Vdew3oVkJrGuEDwPJGPggEgTIsPfklhrQepE4x8b6q
VYFaUWWsufjD4BWYmRfK/q7pENmdW1z3UcRCb7sUdiirbOnU3QS+WOcoiZa1
qKfAUUM7U+3oTEgrWF+qsMDH8HdqtHGr4Qbqv1RoJ0R85mPRbc97LPhzVIoA
G3eRFSy6kL9QP5PQ0pfnbKngWLxdOPo3P33FwGadD3ibJ80yGKfAkg8ZTtYx
dQVFxGlWT6wqBcLhzM5+7TJ7tpkalARZv+WS78jpkczYZ/bpMMXxZlmHRu08
pePKGGRPhrstwmgyHXXrAzuFmj5gBJC2caYTBmlmc+cx1bUBuY+9RenEM9HK
SXgaxuqSNu5MQWBy7gSvkTgVbeziOHqwLnkwwXBKOTp+mRYbc++6LEYhZbIb
py2MeZhSnEIb2iY1JVFzV/jPvxJ+SlloQyBvWUFFZf8IY3To8ALQDg6Xr/Be
/0WN9xl8qG9z5qKI9Dvp/sYYtKl5jXYYTir77V+67Nz/G2ayLd9vlRXhsBHQ
W/RQpCpppYJbgOkj8rmR18rFvbIuC3MUKF/YHteZ5SOjzzmSRGp+YjxvhIFR
H6ZIMAbceitgXV/unKolfWcSoVk+0ZkbSFWpjPi2qlYJyYQFl1rp5SzO9efc
qS86cAN5SurW5k535gKTNLupAG0l2omnTUROgmy4j1efFQi/ibrjxhzlV8f2
YjW5jFKVGGVrDw5G1M7lZdPUj52x6GXQJ5pFtaGzpsQtMn1lZtnAAUr4vAH4
Q/+qAGcUmXamtmUCzK9PkCGCDJtH/JmSwaMo4LNyWoz1YEvjNyUDe9qKIgGB
iWu1zjRzXjpvWYTEr96ofJi27FovdR4cP03Mb4LmdrVlwnmHO6xHOkEtptq8
NIFjf0Q4HD+zOilb/PMRPRI9bVoRXT+/jvfRlMC0fCtyy4vNQPgtsbBCybx4
u5DSTvEHmUJeit14OPLEnWGe5zTx7c9X46cwnza3Y88jnugAisOhjtmIOUVz
X3+iFzwi3ZR+/JdBxJ+QfWlSoTZzwJ6SlGYwOme036nff2wgKj9vVrUrd2tT
XYfEAZC3w7VBQ+qCOK5EURvLRsv8HlEr+vqvxle2ROhJg0AymfGtPe2qbVaX
+naQqKe6+1kNkk5jEoRFdwc7K2bY6GVsP3Ia/kaBjfgWUWBWjHwnXjLGJHCH
Qm01RyO+EnlD9/ebEwtPtjV7In8PMfbFFNwFozbmgqKfTTyZME0z6WFbS2rH
cOGn54c2YkNuBe+fnP5tpYLBDrRksUOTxf6t+cygW0sW+Fo3P+qOcrQR9k8G
DWO79+fR4U+UFqP4mQGqMAj8kpnJuEFs9uni7DWluuXYLpLPYBWqA9JvtAF/
32DfpbeFWgxdqD32I/xmCoxTp4sXWhq2dM7lAD77Jsy/+DrOkPVXB0VS+jRm
bOpSRXlCPDWhNxhC5eNCdZsJPg29c2f9xg0VxuzBQ5FCjb+jfumGoFF8z+Gk
HNTnaLNXPxmRQAkZFsJ7GJekB9KTsvv9TWvvsxWNF1Lc/MSx/Tr+Qs+iEmwF
zJwpzunmyQ24ho7+V0RdIW+qFwDp4XA4fuyEcqYaq89pNLcPwVtZLBoy1Gpy
eeSl64gboeHidJ03UU6qx9f5gAS1CjgWFPbI7m2CBDOGVQxMe2lR4Nk4xn/a
8+SNK363XaKo2vocR7Iu2cgTO06qPnBRBFq7DIejzlZrC3e4YFs6SFSYmv8y
vGP6WrBjxPmnKyJJA4hDVjumrGTBXAavhYxuZgGMd/Fw3xpvti1/MxZ8johZ
CMtIgn+2X/hUmwdcNtyDIOUlKX7Y/YDJ7a74uE5JITOXnN337Qa1OwshWheM
2xU4rjcHRGnBZD/2UOMMwV9QOuqgrH3+e74NJlOq4ZwylDJj5St507bL6XIB
cD9+W83kiKIwkFVAN4Ijxuq0qWoecAUP0wYbTHfbSv0gxQPtoP1gA05kTr0n
4LFEiFQWvIyG85drSTdL+j6Je6bbbXdqOxJuu4gwpOJSxq8fZkMOqJNlpV4z
6u5MDBN6tgnSF+MBvyfTNVffUkBtkyDhfUL+abuD6YX5kUeY0dUWkb68r2Xd
U9ya7c9R0WyZKOF0OIHSunY8Unb0Uf2tf41eK6VqTLUd5y6MWjAYQARYr4oc
7jLMZu32NUzmvH22cJfw2EHAFwm+dtEXhReem0uE9M4jtsS2nNvvHfeyBRym
KNnsTST42qj6K4RP2rA/hg6FggwI08gCu1ANlbvDi5gPC+SRAC8i6MyKpkbS
GJ0bqZQgPdpAokhJDfc+rpZakqhPTGbEPbUDUhtYwjZmKnteMSaSA/UqzHaJ
IkDSFvnapuAoZcLsl9jkHnPPEaK4AWlV8xb+GHDixPiYhbEorqXLpQ+i3oA2
bczWxH1cdQw5dcvKmDHcWWC73hLfT18UN8Z39Yly085mbyzKSijTeFeiKfLO
G8BPv5T3cQphsqf9gux4+swwUqMXyw3WobFAHji4K3LrDol8e41NxcNvE/rh
IDl38hePLaLLjtZCyWp5TzvssbSZulDjNQpVOq8clVI0uMeylgxQbCwXpIeJ
gopeGY8lVB5txIwPUaJhkJHHv7p/ahWGAYDsi6bqNuWPcE5ILBf8YCyQNIAj
V4Z4kjQjKYT3/KwSTBwXu3P/frFclMAWqgG2Krb1Jnrux0j/eeXigpxXR+6F
CVapw2ntL5qtp2Q/svUyMiZRkwBwK05Nq7MDbuEMSARTkzL5TvcbrNDPiEVP
q7xT/3h4qfn+uFklfigxVKGadm1e8lNX5uOAJ0YBsj26bJrs2lRwP0LVp8gd
dqlUECa+UEQa8e8wJSawR0xT5h6/VKGMrenRGtnv4hmaNZ1V4fBUW7vLZvuW
iXjIZJPj9m/+NVuOl1TvMADpeg+ZNqC9hIn4ROz6DLkewp6v6ZusJX2nRxrZ
M6T/poeAh+MHmgI0Ca31eA/nk8KHhzrpTHxUVcLwNXdUCJBM7NbRw2zgKI2Y
eA6GX8+J6X21/ivVo6ZuWuA/EmFvPFl/ewTuDlxMoJkP+XmAmZh1wYylUZBq
tth6B04XGy5tnaaxb+ydSMcjiQtmVwMMT6xFHTbaLR1D1lvorlLB/iN6moah
Sq42g2e/OGEeHCp58SupPRG1gLgle/UEv30vLYBiuoVm0tMm18Z9DyTpu9k2
WQobmVP/FMLbi95nv7s5xGi/KTIFxkNnVwQ06gi2MPth2qwACguJNyW8aWUh
IuTcU1FWy7SWzZ0tTAlQiN8wn2Tc0qQjhcmywi9agVHGye16/XtWt1cAizsr
ONTepm4N/vstUNg4BvuNs6XJVeSfUOcdZmsdV4UrnoQCB3JvwOKXT+M0Mv4B
fZ6Jsal+jIUm32XoCJrh/3qid8c9sJc8TXBNnm5m+tnfOFJ7FDhnbKiiKScS
KrwlBpWP38tNEjCcoB9Qs5AFNfH5xI7+t9g4hZkgD6+mJre1ULO3cQVBOZcV
drq1A970KXZaQDzdIRJ92ikL/sw5qbVIgjfjni32CU2a0inD01nyr5iN/whk
egxG0sqx2tn1fobhO0nJwCR1Kf/4qGKWpa5Y5zj+G4y7zzWJd9CQTtK58138
N08AUHrYA62/H9c+oTF3xqlS6wnrMMFExPE5T9u0KWzAGKHNGSXqKFvxPeAk
zJLCzKYt8g/9pFUzvsSJeNCgntH4aulBWSWX+QQOOttVHUxN3ZFBD67aYPqa
uaAFhV1yqFLi67c+tKyzsYZNmt6qrsEHgJOHj+HKZ8QpMqFr3KxE8Bd3V0x9
14z2/hcQikfcY3esI8yqskUzBO37jRN7Xvj7kp0POfnthbuJRHGcC0cN8V/u
kS2u/8yew2sJfpRCOI7dygTR0p3V9LwSZN70CuRppQR152dMXI+/8G8FdaAA
ij0pYuNT81T1l4sw1x3Y4jaGyRLQspg3yc2RhXbPZEL0HwUmZMhDd3zjMFwC
bV+xXyeJ4FgFlMtFBL8F1Uw7EbsHH/o4W6Kf8dFpieDuDrb018FaCqTx+FME
KcaqhlaLCbFe25Jurvr51hbEq0khnzFsAlP9dW0dj3O4KioloL7W0MML5fHR
9G77PokBIvPFxHgrjsGuOxHhzl6ZyQI/XiZwvlVjp+GLoyjXKAUJI1Xq7z4g
EajD4IcA+0CBGoVoPL/7H8Sh2MyTrCE1oUlZLsFMtRddtGOFEN/P8CMBUTvz
foExP7Mqz68o3zg9mrYkGLEHzAWBBt4sUCeKH7QVevXAnH8fK54QRhDteJ3d
JLKRyomiQkrC8x17tUOLI876BvNpVIJAqnmXIE61E+BAHagtyRMNrLstV55F
388cS7EkVdAYydYcz03LS03JFSqsK1n5/x8NlBuKw7h0xtLgxg/7v2CnWBtk
Ycsd19aks57r2YQoCTOknQ8dMSHNk2pwlR24fjxQKpG4yHbMgP7PKOGLKKde
pTGJSEAhRUt77wtaMPsXcAREbPEGFd3G0GOg6kiDBoy82A3nIaLxzJaoaX/H
9Pc3dgwitxXsahuNoghj/nrH3InLa2QRC/ZV+PWjvzTeaw4+7kQQl+myJu69
dl3rWnkxot2VfBdRmBIJzlV+izpnJ391TlLEAihG9uhlcA8Xvk1FyIrVY8Fo
wtLP6lwuXBUWAHRidun+l8Z+3U4IF07mjdoLgke4CL0QvZ2rE0ROF/5UVAC9
gnpV8IdZiaxxKe2wI4WTsnUCQ2HHQtQ1yws1GBCtYzCIG4H3FwphuI5fUCpR
K8rrK2ycQNmR5si6xdQs6mzHuqRELWQBjIz4lNVOlsAGJlCaRgmuVCn8Nr4I
M5xpn5VOgXz7I5mSqcl2dXPqioak2igQ68t+e2H3JnBt+guqy6MPDqQcC77+
WPQzXz6K9OUSlbr/CCzQrTAaCsVBFDGsMwtSedROKEKvPwmApk6UD0kQnFJH
XghTPEJujBB3jO3qDA6hFdNXlYzstByiX+gs34WXkExOXt9sBEbtW/VHDl35
46W9iHQcZzmrr4WdZLJ6W2aKe6p89NVJxkKY2MeMphGNbgemvGZCIOwPQiyp
NuTtW7arRXRPvJfcF8PWmOU4BF0JRemwil2vxodmPcwu3jfXS0SIOz/yXB4Y
PqOWosUH3iL1zeTsy3y1hT/V4atgL+PGXUD34B0TeL3ZRg8dbGkZlCHxbw0r
EvFAMTgndjgAOVbM2/y9t9zUUc5XDuc/gbiTxv++kUdhdeMnKDySJCW1rGAJ
tX4yf19Tw1R1xOzxVrMxYxPMThufdB6rjKB8dQk19gebz12+vjSfzMcUPWNe
ZXABGlgyNp5Tyd5CZl5V9+GlOXNIxY3DxHLPsKyJCoqLvqcsksxgRZUMETJc
Cq1lhJHQHb+Qg4rNkoiICE6HgGjx1DywqLBh6OSdAb/uzgVceZizvKrOzWhr
eW25JoIe6kxmVeArn6uIEHpGbd+fGuV3SvnoDZo0gjZ6juLi6vMj6BC4wfM3
pEQHMFXOwmaf5dBeSWuPa5HdTWYZRhzidha6zJ8Cc3jX9VLcYqSxVbGuc8Sl
zMnDb5OOuUnqC5PVYdHQBwgF6DbdBNR4BEwy+pHOn+TfwqIA9c4ACqxjmMpV
7YWNZ4CRYmGuqupj7j+n+MVsaWdGg9JwLHNeHQWCRTx90ymMOhq3iycGAwlg
l6I28cieQ4/v7oGNBlAumNUDuhDM4UzSk1XpQ4uhEHvXSqnn4sw4FXyJLfCE
bTbXhKkmFOj0D583FumQutIzXUiViRpQrQmBdeUsmAyoVXBZRCuol+GgalZK
4VLxS8G60ZTGiFquMFmEGRYjjcR13EMV4llh6UWZHmSwPDTBHDQyMkG3G/Kb
EkWPSOpPGT3yf7CtrcRrQuRYr0XeDR/N84RH3+ioJk4uB/w6HGXsay/J4yMk
To/nyPvNc5Dusai9KuBs7gZZhIMVrtKJHODLYxh+/WVfSjPyw78qOZH7b7Eq
lwkbODv+flh4wi/qLfpo5D/+i3nascGuqjfmLmWfK6lGJ0fjlTsb71fOcgE1
+DbumXdYLlubo1UXmqZQo+NkBX/oTNwtLGkyP+35YjZ8bE2N2K0LWQ+7Vstf
fgWQdDV+8Vn160n9bKEew0rqvYG5yerAN3qbWinqAdqrSkF/+/5WjdM5nZ6a
ZgkUuKt5hSjCpvVLYm04JsCJ01eumypGhyj2y+aV6EjJkh8TRT4WPFneIxeN
lTJHlAt9NoQNeN5tgHRXoCWPuwedWMDHyYThy/tSoePOFrUs7Wn1gD62vYjH
jXJu4MPePPwywFN0XuA3Njvu4R46r/a/C7KgA+2f4QGRkn6iOvF3oTkTfXiS
GpJTNyL09JsIKB1xwJ5EsRbvbOzWAOHlsoQrvgfQV9FICDY5znPR7njWITqY
9hpDX9AyNCEM9nQrbGAVJ5kt8kfZh0UmDOjzNJFSpBuZI0I2Ix0oCRx9OJ0S
i33ZLRT4LCfNCgvvik6b2JuUgXU806iniaXRHv0nNHPFEVn3ceMo/94AyyG9
8g/dW2POFXFd/vCJUG7+pF9j2OUqoZ6JHz2jtGNs8WSPH9H9HmGfxNZk4vkO
q+1SmRlciU0LhA+4ME+5+U2/z3YyHKYMswhy9pXYxftNW8y9mOnp/ihLb4Hy
hl6RlPDQzh4OkWkc8NKzBSsBSfFOzQqSOU1zj1HX0aD6YxflOzj5OBgO+/ga
jObUrGj/3RJBPPaj9O1wC47pTjA82RV6Ka9Kx2txaE9GQjGaFUet2GmwxPDc
//6Mr6Xpkw2kMlDsIKA4sZVvfudQVk5aU9kxAwhs34P7as1vtgv5HPduvlOK
vb32shgn4u/tjnmzvSd3lmFBdtMMArGITxYc+PKM4F4/99/rPCRWs0rgY1lc
f5c/brJTtW9wO2+nB4Tfv7sA0MqTrKaTRj+ii/hWkHLRDFJMPTWui9nCwewc
VBsSrdOrMG58OqXt7CeHhTVXtadNxlDlWhQehH5t0Jmh7gh9kVmSey4P5aqS
nSL0FRFO0h3k045W3e1gVfZpLe2UargGoahfxEl3w7fmhlnzxhvKvNu2Ynwc
/1x6TaY8E3FGXgdyRaBoHBm+lCe8pqOUdE31VoxIBWvb1+F0PzfYibaJHccE
3uywj6y15KcZ/HMTiwm5Nlra6Wr+mzNuX2KaBVEy6JVR78+L+z0dk0ex1K1a
giTtYWmz3uVzTxHJ4Cv7vDKT+xsfMptIsivGeF7zx116m3gJ4358bMYJPEqD
DsOmNZdBirrsFFmla4oFGL75e7zoyAUJyXxHsGH/OU2mH3GA/YrUUNE+9i97
kchoZETGQvBNS7wGAhX4R12uiZkTsYRVSL9Efx5CMPe/Hodpehr6Zgm9bmpC
CFgZ3Q1OAIf28kmHL7oDl8XPN4UIPM9tiojLnV4wtEAHCUVwHkrt9sqsNg/8
lBcx2UNFeKXo2CHTy0yIxJAfLbyGmMSBK6tKLMFlCzGyJZ4quVNAtf9Wamgd
vNljiPnimTAQFvmU9Xgmg0jkRxDkJxbWEL+8wxC/f8/9VqDzaho29qVF80SE
0YvwZVPyQAHIwjyMD4W6MqoTcuEAVjaH7Suwml94RWihiTVYB7e7iOg6fVgD
UN90ex4DuKHN3PL4juOO6pOtD4tNvNctpuNkqV/F+aSjC/mdhoJkCWcMLVVw
Ohj4WPfZp3UhkED3sHK3qHO6xQqcuUverkKtpPf/H8d8IlVNCEZuHj5Uh4Dc
nEkqq3OJ0HTTWzpUyhkSZVspYY3OEwmoskeaMh0j4JJuJ7l4nBIrSaGN48W1
Cqa8erffhXDMYkZM/oAC9w6WvG1JVGETskedeahePGFbF82TvGjvhMFETHZr
8jW8FC9EY7xtGNnHNl2WMkA07r6OYoed6vIsfd/4QUYGWcJulrYwwXFmXKrG
9CSHt8IEyaExfaA86LWoi8+dmuNHdBNXPw0iy/ssjgg0LEybrdJHa1VWAobT
lYQSPX06Ht6G/gxeJD4s8pg85xJykNqqAMZT4/EuR/y0GhX19cKglO6ay4cv
hq8oFwL8aP7m+maR2ZjcTfgzr8garUPdjeOrkxu3JCL79rFlRlZvFo5vHDvf
83qdPi6jFbDf6EeUzMiho/+TV8bDU4sdnxLjWovhgxuye5vBumqb2ousA3WA
+nZsBTYQCxXDB1UsUxb/rmGFraSLSF67Qj6sQMF7aDF6ojZYyV0W7hx2yWLq
IrVVU1cmaFB4O2pOWH5o6erMsIdwyXDyargB4XlsfWUoTPWCoRTA2eOxFAwh
wiFrWfAcVq/ti+K9LtteSllcM8HF8T6XbT7XKRrywWTkQBO+7Niq9zkga/e7
wYZz6Sc8MF+65zXqJ6ba5SY4DFnzAvgiCuH4fORkWlu5bdK6Y87lUYTwglNG
Ci6OB2b0Iel4UtQiCfx2+qkCkV4x1bB76P8p4og85+4S1sSTyA3z1X54N11J
X1HMD5RKIRwf7JCP67NyV6LXJKndO5S95ZTcOnz32JUqzrWnM0Th205l72Bp
lP5OCogfdfDi6lAatSrr7Tv3aQfnI3jZPRKsm/qDvRxS7KzXd3UcevVxeJq9
TpSNTx8xlMcbhRlQOSmnUVyPpguKa+1kobiCoVJsx9OuF7rzOvmOZ6QXgE34
hZCKlCkJr+/GR6up1yt+Tx1gYUdrSAHEWFwQb5F9e5m5WHpOQ3KSbRp5ip3z
c069JjX5AP2OpNKu4TEoRx8wyNP9lEpqEA86g8DTEQbOI2UIXNgYZ5m2o4MZ
mnMmqEJX5y68SIGRtUVdQRvNz4jCmYs/EXfFNSA0MEY0Zar7HFcPm35bKcbg
LYM1GohONwhdQNEd3jWx7xn6u35D/2ikfFXjlj7dpz1j76zf+5gNOk6hZh5+
dbnp2efOlnvq02qcssKw4icw7IXGylzbWQMmmtWDg4jkba3sFNDN80G68Aa2
Q23PpXnyz+CnbzT3pigNqIpHmL3sWX8BiNNoSopTk4N/vxokO96Jh1XJq3zl
PqCf1CnRLpiUM7QVagGc2qY0F9VJTZlNCbxd6POJxlmZHIvNSexTaFztDCca
PBG8SvTAi/FmxchwsAB3fLjQuWz9Jmqvh5ty3b20E7zO/V6xzjSGltPb4Btp
epFb8e39uVpWIPO7laSM0BzpJP6+9HMCXKj5pbgCa+TfpfmMm/xEcKS0jIxO
FMSZ1mr0hldT9qhYKF6FOkOh92p1TYP7RpquaATy9djcthAemS9boabrZ0gn
aVp5L8G//zVzTfqcIoJHwYN1/Cms5Ffa0cBa54MjwwMT2IKhRl2XEj1JqCuH
3OnIhplJgDehMWHz0Fu2CAa9BIcwjERQ6k6XeWXvoPqtjO3x/+pNUCobBP6P
FLic2UIn+FrNGPw9ZS+IFLWCQOGTd563W8pC2HkqUiPP8hOxHbjH/UjC3rqY
ZNxMj9+0LXpoWE/bC5Hk6bV71iXRqvQChxHW840/1XMP7eUWKPw2hqiAUih5
Pfs5WIPkxSH3HB6z08Wn9+VpGsqlq0KnRcFjv66bNBOyuhyRJWFiR9pR65nX
tI4YRMGicBYcyRC6DUEK8OPfQ1Wa+Zvw5lXfK4OvDcyhWGLka2IvwpZ3al90
u+yeVBrhS/cqh5tbbWcXnwBzLWiOrUaKN/66HhSuEpoPg8anfkeM9PC/t1ob
YaLLYQUZbHhI7iMGYaQEdOZAFYLtU2pnhRtqRDylR7fLXBDT2F8cDAVS0Kqu
b+OdomIEOsmnZMO0lkbXKq17I9D+DHf1+3ASwu9sWC7iewEoM8PYnCs2122v
9BLFaBG2rMx8Ix5XFnJcztRGzfF3L81ItBO/TZLqBSfhFE+rwC1NTWuBJ5A9
UCaU+z+sZkJP5tQpL5WMEgZp4JJpH3w+VpFcMxpE3pr6Kc6HyAgj+2vrNCDY
a3eB/WN0acWccKPgGm6jKR377KaYvf4FP3rxxXQS/mdzwOXSS4YYNFsmI+7+
i5q03wda+lx7gnJxZEuMYubF73fsAVY31fV1qqhIqk6Gt/r4r7tp1nRipzyA
Y4fqVwS7c3dG1l4mZsX57GYMEWVC3kYXW+Lt2ohmKVvyybivq/iCt5MEEJDq
mQ1T7GMlfjgaD7ROMQv7bEraCWozrEAcw00ceTE1X6eM5JlmbePj8T37zBdr
jXDsuc70EnDMjnRUs2phYpzIFkaubC95ulU/Syw5V3tkwFF/GZd2RB2OEpVE
23nFhBtN5hLR+gX7BpA4mppTal1bmGZpbvYz4vhKNR/kz+gVM/TsxK7lP494
agBOoAefo5S15zqtOETisTOaYj5cN0z/FHm9n+zUNvP6nW/dxwoWuxSS3rRo
3Gmf4rSdgdVpLRhw3hIbyhDkhtFrqpB64WD2ADCIpmGSSAxLR7A1XhMyI4rv
EwjxC3+QHykYE6BrPmDe3/wxiyX8IZwMUSaABPh7o29mvr9v37zSkSt1z/8b
ZBW4Xf9eOKOEBFNstCDb7Q2tfb/X/z7RpcHLwe1l9epXlYvqVD0mzCFcCYf6
AGLZmz5K13tMh2PpM/LSvF4zsgsNXRj0ptmRFOG/Y6HMsyJ0HZESY+quXVkq
f/+qASPSvtgP7DOKSYVjwj0PHSl83uXpCTAiR1koh/RLLt5f1R7Q9CV3dXmN
uJWF+xq+7It58r17QSUnm3t+XPp9bh8ZfSxxAj8E5SxE8AR6KHlGWJhhFUk4
/RqyK6n2uqg5zi8VHCZyZG3kaawFXjqF8Pw2Q6s1XbbXKfjEae37hK2soZhw
XIOhMxAV0fYnr+Dk/M9c7v8czoYwF/Xq8OHak0FiUE/r1lhacpQ1Ri3hL0+w
UoEmZMAYXIDuy0nU1OBHgT2ybLov9Io+AQvEmlznEhXPuCz1E9KueU1a1pa1
6vo4kxx52paIKwykDgzi7yMfSsGvFGL5CaPJ6HN1fxxOOFs49Gkjx3IBH0Vi
7V5q5OcKQNORY89yis0cpHDusuTHg5+4UKEDqDMx+KAUTFKV4dBkIFo+xRyZ
i+zCLcirTg4GVyhpHKGfs+WjxcuvK1BFUUwV+D9Zqswo0viDaNQfBCBFIPCi
v432NdU5RoHMRbWRnC3aAF2NPN23/jo7ruSzSEXO2D1FJ0v0L72y7HFB9rdb
oPjlk6bYhthDUR4EM1Vq4a7WkjNd2eux+6H5FTTHw1lJXEhkQQ6YUugX1kI4
7MEJqMCcj1Y86wuaNnf7Y1APqI0j/NEj54Vm9/cXQH22oOXIDuPiC6YaXEiI
39DZZxvkxJMq3pFIkNqjiX8l/mhltsTeSJCErEYbU7aHkuyf5Obj13mHmqB7
VjEYOCwfxXsllUBhIqCtDVEEv4tGzD2M7fVAD+r0uSE3uxGc6jveKGDdeeq8
EAT32cVWboRLAqfGjKj+OoxtmjxQZUZJO2KR0gjHKjNnpTkgSBdl/QNzcTA5
1rqXa9ij7E1M9F8yUABXA/kXrwZLTd9+aqTsH273wmxoMTJ0bSXzcP0jUanK
f0BND4n9boT4XT15Bl0P8393EdcnbVwS8/pnGhKFskisjJjD3IfmumEPHqPT
c4GqgXNWsh8IYCL10C9yAtbUDjMnvmeL2D7kZZfG/U4uvZyPx8k1mNJfepGu
9tgNzebNcFmrikMz6Tu0GlMsGlrGGSVaGK0886Icqd//LoF78egwyiMH+7e2
19m8vE3OqmhZV0TDUEATBOYeE7MdQKKy08rz36wHFUths/4hXr2vKltV6jQx
XY4kjaFeijgUcSKBAV7z7zBXmNuSaGEXcRsy8m2x04o2MHqdFzSHHPPJUEjb
ilJDExNiTXqMwfFVWmCERWIdn/N8rbm5a9nOsICjsUu1H/x4TVFFDSjzMQks
SDT4ILIvFiGAggPWT/jfhwXQ7Le1KT4IYCxiMwpXFjKGCoUV5lNbcAcnDE9i
8Xw6C3G9iG0Jp+TrlTumUfMX8JyzM4N24CXPhH2YrEqInzvo02bXzF60B4Zy
+U4/jyR6jBY/oNKLJnm29BzE5PCvcXTEbMpA82XTDuz3HXB9S1x6NATlpwg5
cqXHlVEDHNiXAdJGeTWGiVLAgZbApt9uTD1J8Xs0AoFoeii4TR21klbNeZXk
pLBhGn+WamwOfpvkcRABW1ZEgIXzgunov/Mp2ZEPzCtEdxJq12mJDX+XSjN1
6HlaqYoDdNT8uHbmhynbBlR0LIvh6rjfPwxARhLYHnmWnkRJZzuTjP2bIvnL
Ce/ZS//kzhtlEDddQPS/Lo4ShWu0zCMOnIKw1LVkun7zBx7EB4LQ6aXMKvrh
z2wjI2z6PuP1MdCn0bYQWX7ju1xDMBxkyFU0idC5gu0/ZzlbLcPqfCPcvTL6
5s9SuRNBg7zuTj/r7ZF3hGuMHOkRhhABB+hUI/11EjGq4mKY86g6/FuL+4pV
onGw3NQWWb6je+d/mv+5q65zgI+7zoWpnnHOBLrKVnpOQu/uAvELFtY9VXF+
eYDvIMBMCKtYdPtTAzKmeDMDOjQUvlY/PsGw2p85LLm7u6Hp094d/IMg9Wms
HAtX9+TDKjdM7Lcb1I2s3lWnKWPGJG8ULgdnbUsaFvhN+iN71DYH6i9hoo/P
yaaWAhHJDrBs8gcAXRLkE3o/dsMtHQXO/vLLgIEwOHdR0J7NohMUQ+8GAQ9f
ypd+r5g+sKpqSX/qyPuerPP0QWb3IERZOMvA0gjfGAgSBvHULHvMTStapkgN
gFrse9dLzcqhwUIJaxIZEUiUUF2Y2pJVe2XKM8seaXnxwehxeT2ms1zs/u5n
1mccoYna7v6SuFHJPhSYZAZGkn5gRicj5GVYy3wnoEdheu8i+PwhlZl3m/pR
vGOXCBhQtBSLD48RfudI5YMCF+N2nk64n5L9MuvUBCdVhS0XOKg8z1JYNL0B
Bb8YpREouNHGqZYoKcvnb9xBpDhmvR2DsQNAnlZCOpj56+msKpF0ipKnIs5H
wgCKmzoPzXKdnsLVWiGq4O304XfFvtZWnSt5PXifbc8BHhrMqEvQ/H7CMrJw
kyf5GvHBB5egxjuAGkNzpXQnHakHFkfXm3rzZuSjdcjmKq8+gZ4urcemwZWJ
2M18QHUJN5YN/yL12oJ/ORy5h0ZfjHBPfIKkYxJswatd9g8ofwyD09NHjRLQ
EUg089x+WiU6NTzFAp92JUeXJkWLiQhmQgfPll5QDbQIOMINhG9pYnNSAOnn
6oqrkhGaIi4/S8lQc3xgZBKhNFjJnAFYv13hy266Ye9m6t3JUVrSeoWgS8ua
pH3s8Gndp21LN9A4pZrKZegRMiodG9SjcxQwz2OmHIvHAtXr7wb/ib7PtBur
KSsV5dr+IklCiJbTTEr/m2fJCCefbJqYwvlrGtJDBgfV5LBhQEufKTM4R2h/
vkROeNDFTVDejyM4AoJAN/AoKy44A6k5OhdXi9GDlkViA1IxvgNctGtnd9ac
cDeEnNKEO/tnYHooPtMu4ny0ZLZMIW/0rqk7sU/bUeQ1rNkXRVxESUhN3oLi
hke6wOjf12BHyhEAN11HEMT4cWUcIf6t8eLNq3zVkusin1fZRwSYfIpXyZfW
iY8fukN37QM+j4khDCR9365Ujo5pIzzZX39qdSf1uC0EMHNDYrahroNNba+0
L6cLOgEZe3uSAIL/aTCoRQltGCxx36pNPpyp9ZcXKr0FRm0dIJ5OiRdSMdLV
vzVWMzXpNQuYgRO1UNNk7+Luin+JZWLdRnU+8IXU8OFqvKWPEodPF/2WwkYD
rFXXP3Oi38zNE/s0DzukyVIkG7mjzfPIYM3FVfcQrtULJZw/hmutF/nqjaFN
dAjLbXSfxX8C6sstcznfvcI9iQc6sFJc2dPV2FYP4XTZDr/nDYIZ4GTqG0OU
E3o/MMg16UU9yrEuOVcS0BQjgOoJ6rBNE/sKVfnSYFgpFuARfDmNN96TMYsr
I78uOdH7aY6NT5BieA3yVKiiP400SYUkt6rzgsdJ2qIx+h+OuSathWwK3XoC
DjY//wWpDr/UHRV7jJjMbaSC4S7o431+ahAMX3i2ES/kQTmzFPtsWQhgb5kk
HQOeMagWGdFABP7cde2mg307haS9qojUhn+PFh9NFDfZ/Gg9iNYqS6yji/FY
5BT4q4tfeX2Ih467Xu3TpkCTE2H44ocy2GNqTESVN+IYouUGNFu3+3MVfkE7
Zy1UyzyoRRlptnQjY8SUAhRcT6/Ws5GRmixCenGvnZNr1wx4RtMwb/xlJJCw
PNP09dacoQF4IhFGaqjTqMrlNyHFae84TBT7yHmExuYmsXJwvcTLbRiLpKEh
Si3EQNfXnJ7Ix7u9aSRdjdrhkGu5CQcfPUPnClgXT6XtVKn3GuVE+BQ0zedI
/KazxtfDFNtbScs1iaqhH/b4onz137eEMPMN8EdIinp4xJjvf2wOWE67DG1m
AYLuo1hg3PiKNxv+3CK3w6U1B/B74lfbSwW5+571b/bfsqtcvjSq9i0pzl0R
yrkU9f6ZkPqXiWWeQ93PtdKcjlV5BPdC3l4ZWrCgmAVKxSLhTJ9yzG/XFEB/
MZCjT7v/3i+9Uu8YYKdXgg6UgTz4P7QuvPwKQreIYgvynmIWLD0223dQJz4e
f8MUDjHiRcX6wXsN7oN2pZTtORRlPbrVZYcOUtup22ImF9RgxRVp94UUEC6x
r7KKZ7cijXcy7ZPrttQ1kncDG3mPQsZ0MGNMJdvTrKL2JYN2zuLi0Itu1hAa
7MTcqU2LQqmHKBhP9sbP5LuHu9VilBAhzxloPPBLMTUSIxVgEV/QSwZRFisR
6ynca8ZcJOnFYgmcW9fAlPLjjgbvIGemvPrALAlKNwK/ItaPaFdiaOUhymx9
LjKzA41frvzZR5L7aDAenEcojJU8giosrd/q1kNJTZF1qMGxiDxex6PLBNmf
xfXRCnzzEyl5x+TsptvrtTfSKCWLMy0BG+BVU8WjrGBgvV5E4tNsCRgL+zTw
iIGgjmRvw4R/SEHWZfO6mEbsnZuc+OrgoVw6oCQErMI6ipvIrN6sUAIiQdwh
ZQ94+2Ayajsp1+HM8SotV9YNaa8+vz0ryhi2JYBjURIazTRVY0w9/DK/qQm6
rRUQqcvGnnBpKCUW/o3rk9PYqz26bRuXLDWdWGCgBrnKXUn2h1Ou4R28j9kG
cCyJdc0XLQGqdqmQH16RgaoroU+Vprb/9VCxhipZYteCq+5/aI6R2uC3k0mv
kwnbHUqSk+2UVuZa8tiSuycVp4MU9j3f6CfOZ7ul3nxAzoqawyUKEpGVj/yO
hMHQzDoQ9pEo8BvD2pM86a1sQN/HuCHAFcBi9SSUD0JKbuiK1mEoEZxtURM+
Fb7sKws7rehar5BA66LkuLCZpJRuWWFyiefQuVQILlixY2FeemY2WM04KIB1
+rI7AVFuFW27qnGoS248egQi/sGJAsAn9x9sht9U0NcamAVcGoLdGRkFW0OJ
ZkkbDEX5t9IomRaVob88ugGNgilxENwhZpUTAOpXi9+gioWEjbgt8SSnz7di
jzLzBmXSVQKaTvbmETKFpfMsOBElKYioHWM9bpwxM7ECM2cbze1I2P7QdYu5
l3z+/S5VN0bwFJ86atwcS/x2ZizEeNdnZcjN6CuXczPQCM5s6RF1EymJ/CR7
zOFyQ9Ok2eHEBE/4Y9hmc/TthIsUOhzCE2OBX0piJyKJtyaD+/ZRet7qcquY
HTFJYcqQjad5APJNY8ZBBK8bd70LtrY1ImrLgCvYVTeXnXTO5mb3+QFaGD3s
PICzHt4imsKQVNHdhYTBZhppb0U9im7NopkASniBGuRaGw/TV8ItuQYeM8ri
yeydD3SMVA+ulWg1putPKbVByQPbX0mZNHC91PU53dpSG2peQBzof5SGSamI
Si12y7kpIA5RJBNU9UQIUEdreFtF7ovrcu3uJEh1+Il6hlEU0XJ4gi/P+KK6
IMWAIDrAIo5Gyblh04ypbt77vQsaw41AWQpvfgO+ui8EAuyiPj8sxzpz91gp
IVdQRTkF3oq0MXI3XUaFgI5DpnZVKe2ajzqZvYtH4V8aG9l0JxQwKGRaTVXO
6GqyCSzWAS05PJj8RKkd5JHQRRLWf7KugA1bbmua96jPRbkbhngSG0x6aRsT
MNEGQ2vzS72sFKp6wm8kNDZsipoL3LDftD8lT/qB1WMnYMijnr9wFm1+nzxo
n7sZQBJWX55tNV4xaDfJ1xzmuC+kWaF+BTgcawkmUkqh2XrWaIKXxBRqACH1
Sjj3vKHaUCM/k6i0boUzWZ+57NC8QwaihH/hIsNyPx/UbC2zahKAhXS3bW7r
HWsPqEEXMd7bb1bvntik734DeLx2ecz74Ij8BF2JjFgxlYatjO3JsjQYqTVF
2FrXBr06AFbO1G0gmRaOE7urb01S9ek3/+BwC4thrTpHPbfS2bSZZzkSc8l+
kMiOcvpqflBcyVojmqzoHmI4FTNOZ0GM026rMHWA7Ejt6qvLlhbV30fCKBYx
kDQ6Gc+pL6G2e/MTeoWBpycp2FVi6Vl5NcoIZgdYWWtcRbkf/8CWT63+sL+b
jXhy/J26mpaivAgPxAt/es6fCUjuK5OZOWlByUqCYw38LbDyS3E7pHo4r0iA
bV+yqZ49tU4sTifBeu+W7jGLrqy3HhQrTfmOHpF4DbCW6XzIbXvZDG9GmSH9
jozxP+bcW2J78ts8UT+VO8ER5LUjQ2LZuq4ifLgHGhct1GBs57DzsGeOmwXo
PdznwBqXSAQMhlHZQen2mw9Y4qF50XePNGfqpLFk43RW/M0Lzxm5tBIBW8qf
UA/Jy6zDs5x4YY8rb0RCwVg54+pqgvzBUyRLWwKFS5m+16e+7jdZbDQMIYUP
7jJAv5wEglYVHtzCTyQ76cq5xhZFWjV2MjV+7h9w1c+afQIF9wRXh1HKUQVo
0NdLQcQBQKk5Y+kmbekahjGvUcQ+e1Lqka7AosqyhBn6sBwgj2Y9F0x8o11n
D7ll2AJzhHK1aguEKH1e+szIWfQZ7eoocqe0yAh/6+T1kYwd6FE4z2hGHT+W
p1lMONS+KyFWT4OB/3/jOXBZkqHZ9YONXAGfHw3BcFDdKOYmPRV8jL6dPJlH
JyoKd/0it3CGALdofxTSQq2qoy8v1+Wnh7IRnYEBg/WYXWl09CUb+GzYppF/
w5CVslsz7/j32VofBH/zPBCGGQXW5FpQOvB291VvYIO7PhYBwPX+WtNywVcF
FkwPJ4sdjYiGuThttu2hZqSc/Ibooulu3LszagKFdnzeJlwalZQ5rRVFoD8V
Kon9dkKCpgYD7/O1L23+4gzpgLvtTs9Zh4iUdoi2Bhn+UWReX2W1E1LF4795
jRFsWXh8c+ZJABaMV22hLhPHOOY9MiU3Ack9Ep/INdda5z+m3oKAPxBObyzD
Zsrj5IWwyNnhmkM15I8Z1fN6c+kFnEQ5yTDUFL22fyQWIfn1vGVow+/7kJUk
8DcKwiaOtSJHwf5KIr12ihwbswXe3KDMLKexCyNOjQKtS+D2iSBN8BxdMlhs
D2wU6qJyMuDjO91MM49B22gF1pJn/KFGRSk6hh0XakufZLCbqQVDEhkp6mRC
Tmc2cS0vg/RhgESesHcOoKkesXUszIdQB+aKHsTCYKsxVnOdslADxKjYShDO
/UivFx1w4TIR47eIMY2vRHwjwqlZuQsA8FXn3xXtugDFfGuDdxbCu3W/iY04
fTBBoKPu2V0FXY9EmXOVLR+EFISDRIdTAMEwufFoVMq0BD2p5/b/Wmin6I8f
LMVLep/3qh1tYhr4N//yfk0gJBG4KjEGDQYRq4X2g3aDGuwH1vgHS8otqPqZ
0Ck4dIbLiyo8vN1UlnXU5SS8aiH/sPEpHsWAIP8naon2TyZDTYO3XpHWJ8vd
nS/15+NZEJDut/iuQCQI5cThEyfGeozjUeRC95D5K7klxaxa6whagHhhwpWJ
FUvmJ01TbCKIO9ArjNs+mE8aK/z7ztEj69/S/JwG3Kj2qHfcO5lHFZK32m/c
SQBB14nEhY1MM+DSokX3MxrjNtZVvYqs6c3JTBjwJczAFBJVWDFyBYO1YUp3
JAtwH+jn2g4pNtDegFaFryarBBQaiwN6zD+cjqDLiJeE+BKecAd+angpV+Bh
balIOay4sjuWelt/DOno5kmx6T1w57XCE0Qz19mlbm2zsPJTqJtmou6rEmmD
dzy3wXs3geUo6Lfg/1Vwfbfybl//x+cmq9rsr+lMqXWWtY0PuyjUJ4eTHc91
NPi3U6SujfBVfrqBrQPZ1Ggou46RmpHuUQd3EbI9mGpeRFGok42WG68WPurk
W9xQ6Ik070mHdTHljTcF7utmJNIfZh3wF8Cp81/2I4JnwXon3sqR83jSGg3/
hWhbfNlq29HxzgvPlQg0iEzlW/0d0O+ngeDQrP4z7Lf9ccwFK1ebKUwOwZnx
iIVyLHOus4vQe45f6cKYgqxaptrCr1sRrsykPwrspibd5b5fq2BEOm0CAMLl
juiLIJXI5BARvVLYJj5Z3oHf6rggYzKl3ONlZEFNCLbHhrfx1KK8XW7RNp9H
c6eGyymDwOe917g4Zcxi6e/4gchfsnn4QtK764NS18xRsGb5N8ztNpPwUI7x
SADDXl/uezxyx3d1HcdQPVbxd7EQ+Un8fIr5JFLV+b13/hzdmHEeaQjoeCMb
5VOetaHsFIlew0r6JBTfkN9JU1CPjOPgmmqI6spU8R0br7W5RmqjRFLWcVAN
bcDhM+S9QE4vXLrtl5Yt1IZ79oIXcgAD0SI5tT5xmvjhi46UP4U4Szblsym5
NxTgqpPTojTiUZdwfR9ssgp9KRLl08+v1Iv+1eGKbJjLNGiDJkkBiao1L6u5
UtSpoTQrtclvdkTUeghgKHx8v/zTo8FCWh356lHC/SNx4kFpooTqSZlGaJzA
8xgZH7+6b2NEVn60NgX/K+zbgaCqL4SaEpvoZnGk9mj8AsBJ8GtmRKpN4AH2
KzPLSzsLXexD9CdXMroXfgOJK8nSmVk9UhroqbssD79LIePEEFNuYkrT+d2r
7e0WDf/CAg4vO+QtL8/FKltrqDixyeMsCRXZgRls3mk6G+dKyndbyRb1omjO
HDF/SSPiDSDhg5r8Bd4M+IALJsRgd/oSMWA6ZsTFKYr7So2DjmjV+bGC8GZY
xtSIUZTfErtNVbuLJxZEPZn37tM+7UXSw0ocUCYUQHTKwSVKl9O0DpHNdLJ2
1KmqVsEVCVz1QJZxIE4eL/Zg6+YF3G5glSe20Logkxj5fjZjMsk0e+W3qJI9
3y4ribtQkXmLD4SUyGYozDAGkhrFI/Rb5yyBX18WMuHbQBSbQCOwzdynPjuK
TingttedhDt9oiWtHlapCZyo0GaOYJusKx92XxA+FEcxkzRniRphWbyn6KO7
0Sc0DVH9VsQpNwom9DSaHlsn2+vSwJBQXbjmOL3Q4NcYg6DoW2TtlY+1gXlm
sgSGqvfc2zyZ6anvIOJzjuuoYjshpSSjjwZG4sk7ZNBQkeSuZiOoVgx49Z50
nJuaSLiorQxSHSZFBVCaX+aKfAX/58qit02UVZE4ZwkoWraEZtxI5K73OHnl
b4OldTbeKOwqu5it2VoDgdOczRI7aAGNoqq4mVbnFOWOOH16gOCBot+S/bZd
W//Sbz6lLktQzj8tCYEcDdHgsPEuYXan/GzMUbdAz6sdSI1fadDFWp0BY5JJ
i58RpzdICSkm87bywojAEr/wu/V3hIWdphHBfUCz5F5A4bXc6XGtzmRXvYd1
mJlkgeWOTKw/d6oZDl0gzUO4wPWWa3QKKdswzv4wGYpZpKOPjDs2UYs1iaNH
Yjg9pVW6FbtJ50qoaqHnzXYnmkdzTiYooug4Vjw5sFmM0wher05U65YVmFvq
a0vXvc3UW/LX5MOa9P0ZJFAJ7Pbvxckwm+NikMXFBx00hEd6j4XAWxW1u8yg
M5u275CB56zF2EzG+nnn8mUnfxA8q3iPdIjE0TjLRQerRZkf+45Ff+pob+G0
ygDzLa/r4chAlp0Kmw2Jl1VuvS4VrobQoMafEPj4lXKEEcQ9ceh/MytgzMSD
KZl/wLK35mu8fpz2vN+A8XTGlSLktujzCCKrUf8juBSCreZx/2GLR4+oNdQl
ffD3TBXcAstf1j6afIEsRcZvQiJ5at88fpnlUEbsTjLQoWe7jPRUm6z6Ooq2
FNB5WqtpPz/XTSdBa8l6XpsC3XZiAYIRDiex95HgFYwcYvbNj5Gg5UwAq4iX
QBBYEAZkSx7tpSPaFO7MaP8NMqsYvc6Xt0ZrNQF4uRvEgXzkMin4xeCREJOF
6fc2HGoAqiTVMnbXRVPMp4n5UqgSkfWllMfLhjxngGWZPczrUuryR0opdk71
k9suVJ5Pr0zrk3gzWLWLscsV3dauSP11pHx+Gdri8aL7YiUdz/EkpkCSdfpc
C2Q42Da+7dE/JjcFhRcY75e8s9C77L21F4JKCnwG4SfMrfm07VabtMqtXsdO
5UyiyPSArWZ5BxMjhGerwLX1xHSSNTZu26WW+m+5doOSB5inaJIpFTRJFEZU
M3S/zpJrT71FmbO4xM0dvrW/FmrHShnbE16Eyk9rosjPJrS1p+an398lBjiC
InTGVPMNlWRUVX+1k4A4sGAfcHT9LpHgNhkkizoD1v7TPUwgVdzZSJPTt0iL
7LvvXMobluYMQL1cgbZRPT49ux414S/P5megK7kJdpVZU1qX+biNATtHWx3V
E/WIGLNrI4ZPNNS3PI8SuLbsM6S8btV1QTlgLf16QDzfjYBmZxFPIsyoyOw4
DyLl/3e9m1UONvb8vcDHrn+As8u4aAC89GfRY2K+0pPDg5jU5ttSKF3QSvLC
8Rs97w4hhMaSjTPh0fi+CLYzSYa32uUi13RvBS2pGwZiMkRk+NHmZm9Zjr6R
yJvjtXd0/dU0MojKCamKBzRuhWvedCVPFwtvE+8ohem+hWXy9CglQWc+DnVs
zQhJxBK2rVWITTZEWIG5it2O2FKUmmffVVAiUrgXopnz2mR1GfQu/1xpIy8V
9G14HssMw2jeAn7GAs/FvOhSb2YVWyD/lwiv2OUuUapuokuRxZaMjHrIO7Ws
D47fC0BGmKvbenZez4l+P+QdZkT81c/sCxXPcWET8V01I1qRs11scoZqVCV8
WGqXcxtBFQ2cz011dmBQqB9dSuLTINhbFWm76yOAtt36y6IIIA1UTfdN+QGa
igA4SBjjBAh/z9KBBVVBnO+0xdw7buWqlAP8aZsi4BkF+pUXJK0b0WsHeUAg
IngtQ+aXP0oCIvqg2oG4d7SBs1u/MuCzoBKaUWLBUs6j2HaIyGrEeSpLuiQi
eUx8vieL5gAmR8c8vCcsz0OF33qYCSID1/96PWxP4hA9BeOgpk00hDL2evWv
pKGV5DWPuMHvW/gsFwiD4urSmr2Ij/5DC5C7UV9kosQ7u4qGVs2fRV1RLJpl
usKOWPv8T9PtwkB35hwSI4aaJd0kSwFo5c46Gjm1RVXEkSCAJIus88Wilb6A
/UHTpCwVOhNk9T0lrHg9IIqcZPOUkN1b3rTStiBeZditbP+GmFFiTUNclpcs
pg/2T7m8lN1NyesM6iN6i29ZUA3jH+MV8/JkLxQLkvc4JI35f/IalDqPdJzO
CEyhuAI6d5ZOMwQGOYNWHSG/ExnuHyxXmmyZ/NlTEdQSewzOjHrfD8VBhFgo
Nj4cYL9PGqJpOjnfgM0N3ytV4nij99QV6oWIv8/jRt8vm/RtRw8DFiWWevy+
ErWvVF6yHE6nSO9nn3AYzpZfrXjSyCfv78EKzPcZ0xbFgGvInd+uDoRY7Kym
V3Cq4qqXdLVFmSaY2KLPUFzdlPrlghOeZGVusdri5l0HRqdbw2py0P9VqKCx
/C/Wlz7GrMvg1nSNh35r3cXBolqt16zb6Tt1SBKotjmojrdj3QfyBa1Zswxg
Mu4jrmquZxspdq9AzbYn6K5wd3vMYJeGVMMO8yWHsofk3apVIAU2GwygSnIJ
whzPjOpfAtbco5tXi3qQsibDWVjvjtgFek6oYnHKc7/WvpHBytaHsVbQjXRQ
1Rdr9Mnb0ogPXHQa0v6lLJAgRGptsYONarBPUwDwJFWRWLDHBcucSwMug2F2
5a0UVN61UdInaLqQcLdzsPw3eneSsxsIwDDiMlFtOwWTjgsmtpD9RnOx7fhb
3hlKWdgTb1tZMfBi+uIk3DnUuL7y7T057U1GmcOqUT7YkSVm4OIyG3sinnIA
8qp/9jG4trxKbaKkUszGRTrdNAUiMctwQbM57KBPucZJS2XtSQr2QG8SCPJG
D9lYA9yYAq8eB0239wxL3rf50SoOr0hBRHehnmzYPkAljBLJy7c8EBlsWz5v
avtXpwHX55lPPajWTex4eiHilvSizKydX+J9FtasvyhFPfYp2dr22i/rKfTB
u4XBgD7sKGSTEKx4h+wJ+7oYI/FysHr3zTSZNDDspEakfQbStfydr31aBnLZ
BkyE2qPQ4kJLt7bJ212Q6rKmgE41zrVSHvwZifqH4tvwpimYEwggUixJ9P/u
k4hv9ccRBtWX49HCPE0B2GkBcZKhZ4WyzO9vy7/uG8FI/9XrbKqhzaOkXuys
RRKsK7ZcQk3rdP0NzZ1hBbXRMLMPh/ZCfueNtUBU9abocrxwONt8aUgxHz0W
YSSW7o+HL8m+lNT3it/Cx7pP3HDPxBwZHFUbz4KmjIYXIF8hVgTHr2rcbb7J
YDTFi/YT3giHsO7WVCVLtm1acb87WRzIdU38n63cymA/3gIk3zxdXrtmmzvJ
5/3SGVS25ZDlUNC0eEUG+RGlKHIWKDNaZE/M9QA5EeYRUrZR+ac6hOabpg3c
0SJg8r8E3Wd62me03UISRigdC4TUBV3Y/3+JEdV0bVi4hgx/OHFogSBasArr
Q+FHV9pKOBHL+0LN7GuhtaYyta0WWcZDhnE08t76dWlbUtSCd3kEAewdvT1o
ov9OHcJI1657xTuJoztxsq256U81DUHyiihA70JdCpZFe5J04Bw6A43+ohTS
KoRbQ9CSjSZ4pQn7bYuXfkCueAwR72AjYbCoO7sUnGfSs7BwN1qj7fZlj3BJ
ZvBok7O6waYI1Idu+Q3eH778Uhcm3xvt9oxPEt1Y2qHXn8Lvfn1XAHL5jQ/c
LU0bIXDU31dx2B5p1jUcc4KDezwMtnbYXS3W4o1wxsCKH2E8ghHdK/SZNfDf
GacwZO+NgxoOnCSDY17rY+z21Gs8vP851QlZXentnRbEPiLT7czlu4dc4CjF
GI5lTNWvxlsFEIX0C6X52dw6XMEw8QKX1Owg7mCzwsORBvjN38VdlGc7vWwb
5iDldWFzn33ZI7JxokdknSmmLmwtr7PqSVbFVxgJE+iwy+yBDMTGT+J8hOzP
95kSKEWZc4vnDwN4iPMtYbE9xfk8IDCwLLHDFlEa62/T8V7cZpl26T2Q/NJJ
vHkIu+HsarIStVwO0b0T64d+MYVS4qNy0UfRIp4bVTGmCl1O5lw6JYl+xtuQ
iOYQu2AXNDQBt9uXYaHeQyXeN1LSrh+E81WDfzu/lB1Qbf76G9AttKFDM4LC
qCBoYhRq3VF1jHLJ8skSD/hS8UTfR4zKXbnbG11ljUw+LZZAozzEhidnyTEy
+NpLdE6qwE1WnPe2ROaw19i50LjsCqY9S+z0uVfR6k7vN4FwzBehMZBO2jfK
tA7vlJbGEzUhk2UAa83+jGm9EjSn8UhrE9kVeMU3zWQJZUWlsc0mWQhhoeUv
3zy2QfNSO4Mdu0d1FUOJ1mMSXjE0Sb6qzgZz8SkfLVIt1yAA8B8MCjwfXmyz
JSw8Yguv439GPhTDcEh5+KpkemG+X9Xfm5WMNt9PTJevtH0kqnPEAHJ/2UFW
KlNzZA5TgvS/KmPnbU+JyBLEjQ5qZzitlPQxaLrvNWBaKgXXjkxAhYgZiAAg
9g8rQkPgwneNlCbwZbSaWY+njNucIYdVvQYzHk+u3jrQE4wGaW2CD6Vyz/RD
UaaSQVLeWhUlP2q1jcZzMTkMkNugxNswAwZKJwu6TxNarerJpE/RD9PXpFnG
4phNqxDY0czY5izQJz+M331Epmt7rcy7ux0EJeBo822k6QPmwQNMRdvtQqEm
SKDdfJ0KH1b2L0DiZa/meVLCsiTrUlHYUXAZl5SeeieJ2xDH1hb5egNvubDa
5Y4/k9pe9Otz6PipXk3HNop4kxs6GZefaJAPk9hcKHhHoCzKmJ1DkXWRs6Ac
8iezUdNN0Zi7az+y2929WTKzBlt/SnkHwbIF7q0EVz3GKjfnJne4gkkSpUnF
2c8kNFsicNM4y7mukVXugztM9v5Zn3fD2VudOtegQFSZ4t32HA91oaQZTG/i
uJs8BhjAqpExaC6RPXnU2bhWexrDE6u8MJmwCybgxFzEdxTGtmYmtKyEaxRm
aIadW9kbFMnwaaGAXleasUWF7ICdxSkCvH6ZZjYZNVoBEsL2r5II+VJlKPrZ
JG3ai/BwS9QA6xobOtFESul9rlnoqT0WKUTi2nVvRGcppt8TtH1W/KEwQ03I
8hnLkF2gfheFB2Q6Z9IHgH602o46H8v0Pt46ZnkQKTgUuiCVD2gNX/D4+HoM
3W5DhliemiVPfmy1ORTVtvqsMckvsQd3yOWvM3C+t2Df1LDSDhS4DscVUIzI
aEZIOVb1boxf0O+LPH/PG/OMGiJhVcFjFOV/DfNX/6i/ed5LKE5cgpf8gH+u
p7oiaxOrAAztGg9baRMgCiLh2qqtY/FnVirQjkIPS7SxatCHRPv6SMikhj2A
Hmv16GCaJIjqWUpJ8gzwt6VT87UDJNYMZUHrdqoXwVIEffxmWKNqULBO74VI
N2BNJGATY3whFnZ1+nALoc+4gHLXJB5sIVVer4WJQNKIg1hZ+eq6NIMlGgB1
B13wp0+TrK77zt62vX6StMJJgR+MlZqfa5zzYZHnrFZEWFBobfj/Utz3shJp
JZFSMxkEu0uQ4K3nKQgGVNCtmLe347ygqyyGu+OPus9BDar5toeF5HEkSpYo
hE1yK3ib4/LboWrvdp9z+HF+nuFphf3ZP7jn00SGUa+o5lFO0olOKkf5qtrm
v+M63RdMpDtRIsVBXI437icVheo3OOdw0hBPAVW7eTaXceR9Y/64qRw6bxdE
Zf2uJ4EUojsosZgnY3g8l9+ih0SdhWyw+dRF08gjt4y2lmlMKLBDUmuwUwGT
CDcaaKvk67UeO57vfHW1XXsVhp2cYwnQTkOg/IsYiFrLJIlSIjO4iDd+7/eh
RbZQYIzoCT+OXAQLq48W4MeOMcyi+LGHl9sdGzdUwGovh+FQU3GgWNBlvtI3
UAuNdIKnjN7hneMTIcqDxxXn4uYQ9WCDhwgg2nvlPkGlCszAfgcZQZHOh5vR
V341Io43x7KUEEcYnEQOTdjdjD/jJpAj/OqJC2avJb3mVlSGjU9O41GC2wOx
Wyl9VCdvTl22YerwhUIxADitfu1r8hXJUbaUQ8InQLyFEXVbmDZASLywd1ws
XfKOfBe5UIUFeyvjTxE0CtMCGpL9oJj0phzXjvVZo7lN5cXIljZ0Naq6D+mg
8O/MnSOsThQpP7F0CXj8snrgZgnB4+Bn6HzIWuEWENGRaGv/gX1dlIwN1/gj
m3f6DnauKpqw3fYMfNj3Ugy63uOAQPZ8kCEUsti7/Fj/7iDLeedeLlkSbCXw
dJt4fx2f9mVbbYYKmMDw0OoYsfgj9b8XlSIS5Wq4m49WAOpjpbhRkrdVmMTg
e9jwYGi6+nrwczySyF4jo/tr5txFy86Vp/SrI/EL2SAKA3QhkwYLSyYfOVS7
QdUOsb/be4E271hwuzL9HTKoW/Bxpp7+Ka6TuAlqdIOG9uETUf8ezSmYj4Ix
obn/hV2UvMjm46CXTdfAKzPrRNx2SF3GADgOf3AVBjCibxI5EbftiHbfAosn
m8lJCuK/r3h7WGH/k+tBTcyE6knLu/J5JLgAgt2L3/mtLvWgPhfjZqX89YxK
NIG/52QPtf6CdRTp8O+4Pw/E+jPmHLVjNCfO0lzP2sNXXzJ0EIFlbhp6vhe9
HMd4Hx2ntBedv0V36ut6NHqgQMniYR1ewtR4Hv5LkqlnGt1LJsAAOzIMp9Nq
DSz3cUoRb3fR4+UQq63uZUFsXVBv+ptJHcmR1u+lsDwpFQ6Vj0nKhVG2Sr/G
knQOyUqUYwFScDcCPbuGlWNbPZCl/Xrks4GLUMwrD4MueFKXcFN8Qoz9b0Xi
A2JuQKwzUsLlxvZEhMXQOMn4ymMqVg1LmeRWUHOWyhwcu6lTPgNRGZusOe7y
APdUYjAe/asSDOXEpr06ejEQ+/6su/WvbEkL0s8cf8alOsGqEiL1tD+1SqdF
2Yehr1nnpqIK767jayWNmdfCrmV9O5sDVA6cIPjR4Z8xMcHjc6q8aVC1vKwQ
LnsBVQWpzGPKs/gIZ6wpQfrC1wPEaqNvltPrpwnZ1hR0zMwpUWlXLviycagI
hap0dSMwp1YXlIN70d0ywEMxhsaLIElDTK3RWt2frKPN+7t7bGXH5Q8UxSnc
Tj1Y0TfX49Hb1cJMq1ZyqnS2j9aNbiEqZxLZDPPcBCoh7sFIfZH9q1Np43UA
eowe8BqLjTAfMGbAzDDAsxUO2dKHUQxG22kHDsSajMlJ2ahVXN029Fpu6KDQ
kIoccS5QJ+v83a3e+KM90c6Da5yEDjtnKifmrCbxqdGHo4+4PzkBrCa+UxvV
RVok0Oh8eqNq3JZsQyK/9S/o01ilwvLtCWNKd+BWHPPUCFFmHaILlw6c8KWv
tc6mYrwdOCv4wprvxQT905KKfIio9JnrZOBqGJKVagS28CvPpIO/YUwTYXOc
QSZXDeKLEhDOJ6kmIAS74mVuLOQ614o//aQqWupoeAbaC7JjbvhymK1REamL
P/MO4amg3usyA+FPE7kIa2gY3w7dgMtZ2KqQLyZlrMus50ayHmoO3fEHb95U
d+ZrFHxQI5nmY5n6Dlp0zYJolbJkp/xvq+wDY2xePVTYNYvYLwNyeQlXzX5e
Bfy6lLEcbJVUtHVPgN6h5TsuHTGtxUI3TPb2bXd+D4/Q5eveGIUfvXwqqPiY
XO9rlcr5hUzI+gvTqVsN8kZnkC4e92ji+LvC9DmigvcUrjOKxnVFxEwsqxhj
BVEAQfNJsHClVIISnB5ZsOQ2ug04xqf31/RD9xI0PQIQgzyM9D5t3/bUGQFt
i6zf8lkgX06M0NfPijoIkv5yxrR6JcSmGvhvBsgyH97ZFRBIGlCdyqOSzbxH
tBsi0+kJffBAkWuwbJUmswTQE8wPNvpCl7q1TBEPWfkH4cYKUWvuh/klDN9g
7vqzxMfAMvFdns+BVd9RT2En/A8croVJaQxaB5cm0WR3wI0Gdg2oKNAwdPDF
34eSfi837SAHrp7ro0zPcK+JCpOzRQZuyhqymMYc475vLJDZ2sRJn+nWPpf4
0N0CXLuqg8ADyLrp9VjMzM+V3SpJx0vF+LnKFGBsGBEW5ALZtF6+6vHj45gV
2IRhy6Jy+ZF2LU6pY+p1trgygoE9RYeqX/H7G6JrKKabAGLko7Hw3l6dOhcy
JHAHYsWntxQ3Wyt8hcwTlyRecfbFi4HZY41Xc6FelYrcdE6iQUAC1ZXtn6eO
D7ahqjWIqZ5mnNSaz1a5wvgFw7MWRGiDupoXlAvof2iTN0k5hKcQhWBjdQDM
JZWpwPSvkrvZr0kIKi4QnddrB6zJzFSbKKc8GhIO8N6ttV2UiFHl6EHpGaQd
tDdh3R54T+XbW7rClndRnUCZwxqfFTTa/uaxHYe/u0ouUUgZcxbKvYQqUeuB
rDp8klK0PyknPfwxybmozhuJfpBoUcdNWp+dEWffXUz+WbFVc2bDPArEw03Y
sbZaIA31qQLorbikMkkoc6Tkoa4OruePQCaOiJxujdzI3HxL89MDMApgb4W+
vYz0Ij7/XoWdtun9YXESoPtC7i2bT1b9d50jr5AFNzn9vUnKYtoevIrgA6uX
A5lJmwgByJ+KRqWNhlMT7B0WRXWe65r8vFvHeU+x/OWRYd/u58l5tC0tKtWe
SGKqrOvNLr7882vcM6Ryx/xJYsjm45ebVB5NtS+yn8touVtDbYAY39aBMnKZ
eAcCb/FkDPK37mA6O9BAtUCmbFKW+mYgdCAVGAHBzXkvU6MgBJq7Kb2Ha34x
wJw8R/HXuM7hn1I8Cscv25OC4qPinXSfiRO9+q7efl2xdwDtNr707VSwo1OT
jMGRKxTPaaBy1RxRGewoTfXbs2xmeW2ZxRRn/jgqwZUDBClLMdYqcIqxZmBP
c6iA/ihXF0y4Xtq5kYD/WjJtECocXGOa3OTbSbN2GZFBO0yR86zEHFab17K/
EoWfMRui0Inuxjrk8hcyeee9z/OFxlgWQPM5eWqBeAV5C1GixT+dfzu7kZ4K
LcwXj/uUFF8ewP+gp4+ykoKJI1iPZh/igePPQnwZ82EUb+1mRAcpIJSq9/iT
SNxPCw0Jp4COUnBnfSxIy1YJ1jflYBHZ2k1LZ5qazP+lteMEJHcajxdYbxi/
UeQSvKnS1gWpI2W7Fuk2abrHIxZvuKl6LonizLjGBzZHZJs+ii44KJosrBwz
doiF9eLYVnlp4KpQEZfBy6QlhXT9eAhzPaT/rjHI7vkVc965blqsuLibmr2P
WHLxcVlFSrklOXWvAjTdZAfwAJ8yUyYgdptNv9bCpSRS494MUmwReLEhXXm6
sC4yOOkV+CgXOakLlbL+dU93ffnH5n0dsBU75XxcP1VurJZpWA2Nw3HqiToi
tQvQzehng28Svq6/6JZTG8BJ5/PJ9Q4SoEiIvrTjustyGCAzl94+zo9sIS65
O0Hu8DGuo9B2/WyCV24i3j2fv87hTfbgL4ZH+uNrjegSvTDbkW6zTgPqJ0kI
UO4IIYKLzW4W2xTBGtlxRQnNX3WLBrjJJIWjbgXbujEjBcmLikN7iqM2KNVW
3QGuyXRS19mWv48TvTWfNOdfnUb/gqT1Z60PFHrk7L4o9VuGFKIHtgXv5/AA
6qoUQICMISoPdoINy5c+HGufhCmbCUxTO8kWRU8kaMdDIFw5QOFays/n8wHr
uNY8YtiYAmHjaGWagtwvCY8xn/wCH3HmKp3iQ902dqvkkOSw4wC4MYLKyG0t
3fcJWIvuWjb98ljz6ig2gB3iqU82SWWezKXgph5K0TFrBGwA6QV/tWlsHBPJ
o5KIyOdupGggUW5ShOzKAPgovD7H+MB6RxnDcou0nphmwJbqRBbx236yz7XN
9X8q33Y6akpBbjFHekJC5+wY9AupB/aEq7G23F5KG/OHylkyIDpWNg1T3Ln4
5oaAr1M9j1dQcjP/nXEE+ypu3DaKSf1aVXnmNVx8afb6X6ilmM8AZmp+Vc2c
SFBd1RyAkyj0EGAWY74zUOktSWZxGLn4mBzQyZA8rSDQJis4OhlgPrIfE2Rb
z2Up555eZdMunKlqRIEmxBt1VDS3iJaoWt8GdQoeFsOfJWuUtVZ0Y9UAmnxe
78EtC+3q8iO7lY151qj1jscWB04OQ41pZMuNUqoTplnJHr8MtDPayKBnwfz/
lYMO/hNhFEiwZbyltoWs0PWc5h2k0z+VZQfQ7plqBeKmEmy+OsNCXTXNbxA+
FkEZqpyCXv7mHRQZYzAQEBJmmXD6zwBoKIMENOlwmaa7fHYH9C5gnjS/KBoR
gxk83bEFWYmvOzt34b+U3vM9+lq8WnKrTGBTqZ38lQde132tNqwz6TrA27mj
blbHFjvbuEgsxMc0ix6M5JFrmwa6gRWZ0IFHDHQnIEagdNgGwFCd6T9Kz7J7
e7QS9tIK0TL2KmU6CKQwttpszxJZKTjRYZrPIcL5iBA3RiddxIx8ypp5vaww
+WUluJ7HfF05m7SLLQ05Ov9qZK/8bhYjDEeI22Ieoxb66yJ+6+m5gMApadfJ
8pdCuBeTBN5p58JjZDh6TNv9HkiP2WUlGJEy2urAraeC3G233RxIxWueSmAn
4wopnZKb7C2HmQC8GhqB2A3DXlg/tk5/B0QkPSuekuTVs1EoUnHAa8vuSpDp
oOpRQoIjClnrXIKe4Bg5tmHCP0fH+pBZDo/sbNTQwXhKOjkIoIT8xoVF/fVT
/dJ1aT8UVp8cRCzQphJW90jDcEhls9flKNAYBl2FKl9/VqS9f7toAUbsiDul
/dAeY3Unlerw0TaWCN6e3SzyjZeXkT0fTv4Lh5MlCR5uybFpshoMCjXhxPdh
ggGTuo0YYNScXMg78mu8PEv9fRckS/A/eBufdUjm1DkabcJ8K+Y+oOzAraz2
gRfGY15k3iRvSeuXrxZUbNdCuIeTBbEFazQ9jVgIrbrbWshfcC69bMc3XVUP
8u9uIub5ut1X7Jy3FG14mEMYXsE7eiQ7iPK0n6pHNu5+7d57GDHHkTagJ9YJ
4h5IO8HhxWBPKSqm9gVXGZd9+XqPVgV+fXfmDqplGL9i0jvS6qzB2buXXX98
BoT8umNZIyooBdarg7JiW553FndRGjHOVUE2tgtJT7Hg3F9yRb3t+nkpY9mA
VJWVsNwijzvPmn+sOA4qBn0H1nZWyu8/5/jmxAmGt33sePyVImCiTyEPzcsh
AvCaoKtm3OAQZMx6d0k52i81+9tuVnjwEP0y/zPBStbFF+Fzt9oZhRT2Bvbg
tJoDnCzXzbQDXz/d1+nwVfhg1PkmtV5h33QPtN1FiT1c2rsQdLTdXSllxMMK
IGMidnNYRVjI464xpPMM/Uonyb6zbk14VAxymgDyJuSv3xvXwLO5ki8kTOyq
5cnox44LS6A3DtRx9y11bICzQy25t6/R1C+nZi5sWUM+GdibgTQEFvHFyyCf
Q71goWxKfR+5pIsO7LDFEznOc6iRZMbSB5alLIlIIdo+lGJiIGCICY4H51c+
e4LCaaTUFItxo2tKN1UyA1Bx1z6gDyF8fqEo6Y3CJay5pMI9jnAcFW524oVN
ouOv5KHD/ZEjHuQYbO2k836q6Uod+aV4hi+h9gDw0fq7GD1wLlc7MkIpkjSf
uy1IwR2pmCd058vkmtFbWe+Ay55PbfDu8SXD78No+WXIwlzomT4p/F6CAlDs
VxTFf2rQcjYIi/6qbjU2XPdyAgHzLQSUz0TZaKIYp4CZAV0yJBJQ4r3Tpyac
tzH/JQgngy9nOxukQAeE+QWFEikpeIlyx8KgHxfwF8edCDAGi/9I55bJUWWa
FD2QIslR6VssgLuael5pQyPPI/T759LUIOoiyIuG1fV884N8P2VutuvBO960
Wd0duCseATeNImI6GfYKynwFHXaUTji3I6MJlhxOghZ3omxVUxd8CMr/p1AY
6srBiHMxGya90BStq3TEIw04d0hrHlSb8jq6MEmYOUPAaecXsNfNSv8LWzSQ
OCtMMozcTiW+MirLjf4/EAzCRR6Kg1STLE3r+AAkZYFFq6RWs85APSwqrrdC
hWOvDXHx3cfTmhfYRdTL42AoHKPsfaTYkEmjybS3o/RvWY6lypBT4KKUUsf0
7blc4BTVFMP0BdhkB3jhrZtf+rKuoUUa9ro1xlOcOiFaAuJjtD0mRSxdPcfn
wwGBKq5PTfa0Wlu6JhFo+RBbqjSwcVLahiBCyPGDZtpS7Da1nNAChpvCb+Ja
NZV+Jv8XTM4mr63smQyPZ187wLwG1oG54liQ/va/v5PCsH2SPTyzX7+YAnOX
61t/Kv++HmcIA3rySbnIIMHio1D6Bp1OrE2uqqt8vrAMj3Z1tm6XC3ySSqki
l6vxrhpcD3a7fuOqDP2Ca3c2745mCTG4sAEp92CEGMAlYthbhsIzsXQPnY6o
J7SMuOVUib60o8la+RVDXJoJm+Epr3b928TqnzCYtNoG346rAOJove8M391T
pXtdYVNBpT9PLn2oH2CXUj8lPzOyIBFSE+Da4TDps0Udhrk8EjZ6PGbjspqa
eDkglV/8y6E9flnSP/jl1fbt0XFBDcQ+Xx3+IgRMWeNuGv5xQZMLIrXSk55p
cw2M3+XunK8OYH0sNKw9cRmX+zcvcVTHXWvYn0DOwvvEXzHIW29uAKWwXldF
VHkL6GKaeu7b9KO0VfpFLit4OYak+TzJ7fXFljaSs76mdn90mecCV1cK/A82
Lg6HdVi9z4l0hYQocOtfqa3azkjDWtU+QHaW2CVAKZuN9W2POFfcqMFjkRcY
L0/tFcBsPGE/mXaC3UhPiyZZ4EE0sNf1IsibX0BVJs7mpnmPKXSjukrN8n09
g9fU11AdVTv11pahsBXmkd3J5c5rhGP2ZXWgV5ms7aJwaC//WVChLmQExSqU
JAEeFuH7TLFql9ngMGQcc4N0KElgEvxlOnMZXZbwNxP+6PM8NCMRkTHTBiw5
QYxtQAk1fYQ2gigcCdw7mmFUtY09yjxYs1LKMxaKwnxF0jtxmZTJj4/LkfP6
qSI66A3OcQox9031yhxkpVovbtlki+mPd+Bj2L9sz/DZBZ/C3Vqt74bs3zk6
wQrdk9pBdcCB1XEkOX/JAL9YR85mKSpV6mTpiy9r8+35TwMJOZs8IMGqLYdd
nDQ9QvuBn/YWVBXAOCLWTElqrXpN7bHWLRhzzr9O0579Bk63/eUntG/JsU9P
vZadSpejgN7jCkzrKjr2ok6WMHrDZwUkdhbyAIjXX8vk5rLEvWT7MVHyH52f
VCi/hPoN5khstKrlRn8M01QCcvZka76vNO9RS16Px2481m2HTPnQz6Hp0Ivh
re+HlC1N5DxKIkacSqhXZrhtnjI0UZbWK22r4yVcQcWs5RfDVVjI4IIhyigq
aFakQbGDKBTxDr5icqIXBHoIF1TUNWjAlHFSF5xsK2HT+RLiz60m7jVc/lYi
aFnXbBhDdIq1s3aSLtCmrE13WVFZvKKj48thXh38OFwpvXWQdFljmphb/bk4
62+atLbr1ReQbb4Kk0YeVkudh0U5qIfiJNfOcmDzN6QDW//DboKyYFCP66ou
lmSJQe54O2UnET3JKhHF/CEhMTFJTc+L1QZ87yZM+uVny0Z4qruEORKGAxvt
vaGD7/uEdmyzSOx+set72yao/vzeNlrvxjIMKGAa2si2dFzllCsbOK2/CO4e
ZQhY9ZETr6r8ZGGlsf9dOBPnni8dsyJUfbDQAmxqXby+atI+qru+eWq0mi4M
9Mqrpk3aUnaUiWg5mqlssz5nsrQnPDEQ71MoErQTdu7h8ZjO+pXjATfdlmzN
LHHv/rFq1BIDVPcFgtWjmT7DIe+fkWmz3EHcbk02VtA2tgbn8SrPxGUicos3
DyXrQIe48M+jXzQHLV+Su9WHQIlm7nEe4NJ0Gt3rbO3df3SiTxYnduO6z+50
/XXlcgUZnvNfvpSSDSZK2y4eaAJ4NAK7mt5EoWzH6y9uFmQRsBbmyy90FlFY
ZRtd8USVRX+b10FxVFt6qaRFB3GaF6iUYuQ4daFUQ25TnCG13CO23ATUT6Rf
W4WUOPLZAiJ5/L0dxeooLULeVUNLOi12D+oWfur+s5MndnOkXSYkJhoZcWp6
+6eCURRWI7RZ8FNqvfVqzyHBDEcUO2tmphWBMMP5kE4lU3Lr96MXHwoh2JBE
0LlY/yIBWgwrTXN/pyc1CPQvmOGvJtzPYPEc1xBFLP0okOJ1dHuvCQFcJUzG
1hUlQ6XqK4FdoYeP2itIEQRZIk7XTt/Eo6fPc1T8OK8DcCo3T2BXuBoCdkMt
nAuIbB94vFoFB7uAAGIC4iaJKq5VUJPGnnDli1qTLAoNSnuN8HDmvy7oX4uL
X/GV1mg0ekQ6vBmTjcl0yPgkTiTG34iqPlEjFwTj3fuLl4jLJOVB7Ge7fPJD
wOSNDgNT3FqJZJ2ioQKwRSUGlVzMcAr735dBg+0IiZ6zh/C7569JtzHUSFyM
2+vL5xlNRoD6H5nCX4t8TcdTKQ7UZNZv6JNj2jELsnj1skuTj+03/RfjM24w
ig64xZBZmyyEqAs2tS+bJRo4hklcYaIhUpa4esjeZNPHyFaeBcOlfVowham8
2SxpKWuc6Dyj44KA91wg8y2U7PVOq0gK6ouPDBnvS4/YyDW/8jQxycVJ/761
ZDxCmruwYVXON/aANDkM2s77d3491FzR4gycVJNT9v9Jg4bJ/2TjNDJ7PjiM
Jyw0jdYO2hdbrGpLooIt+InX1ZxCsD8zFygp+euEPPA8s7V0uFSjNFiQi+nm
lO7C9DDY61+Bs4NrBd/Jx7IDzEER9pvrfsJdmDWJ9DEIy4jBaqgtuz3ue458
Z/K6+rfV3nuwjd1/n41rjD4i2uO7hpffVUFXZpKCR3FmtC6ICLiIG8gmoUFf
GKO9xPi8XDVtqvJlIRGOwCyBHfPRc0Lzwi7KKRyvkPFZN8N8KFDbK2vE719/
5gun/qPVWX8IJyc1dL6ExcDeoD76FUydADgRMO9nMQ4ImTM+JPX2rWXnnVbp
53Y4dWpOuKPXrkbNxXo7o5rEgBvpz6yhr+qB9pqWXUrlENsaz24AVeCvF+9y
9yG0VpphkKkjLDkyrRvV5pV/r9t3b860Ofu2JuhUy/w7YTeeqma2Q9DfHVUr
rHmjqpScaTEnvjSNXSYv43RpAd7cFZ0V6+ftIOt7ZCYOtGPfzlt22tH6jlx/
utsBTM0RflPbCXgKWumrRYVK4Qs+HjCOQWAOuccin5ox0TqY7okHZAN3Czje
COKPbY3wzfzELVJ9cEPNlePHe2AyCtM4qz+PkQeX8Wx/sDWeOwFHOSrf8Rum
MHY1u/6CI8tnkrJYz0vxJE5F0M6UBgX4vUKt24pM43tL7//mPpa0pmJ+w4Av
kbsAUgNMrJLlqDj+wDyxo1NUywFb7dns9wN0YNPOmtyvuvxyVZcvBvXAiFcO
/tQWttsGOg2lZJ+ot3owpk7+GmsTw7P6KFMyGbH65lm42C1zqzmngbVsr6TC
eZREJ9+RxrnspbYuTtNJRr2UYrYOi8U4MsrBa4VZpAiy7dHxgbGNTSpMdak5
K7nF/Qw5cG6qVeRCSkIzKZnvaOIeTQGrobZQYwRDxGIciMH6WaLpSwthWjLq
vjgq14nqb2y2RwGsp8oQbWCHVG+MuskobnIWouyZiONvOIfl2/2KK5eUaAcm
yfldv46H7Yy5uxNN9mR+CmLb10vtR1IVCszFmylZRAIYGSsEHkMrFOhkHL2B
mxv7XOh6LoTVs8HEGnWF04zeInmpJKweueF24++K6CAGkQpF63VHpwY4yf8d
C9anh88wS9d729kNZui2wtkwlFBt4cBEG7aZ0KZWffE6pIGAkz5mUcocl8rH
6Si2WAPEUCksrQLkjwJoug6EZwXVa5KAiy+MsIp9cBLka5X5T1S8i9/3yXlr
qafiNeczt7biPKyNDRh70aTrQd9jDgwkw4lWskYP/bWzVA43anC/elmyi8Rq
MPU4H3OiG28V7sO0HpHcRHMLt+9TtzHMWFnH4PsV4qbJZ7+iy1RvaZzjmKzQ
Q5ok1rnWtX36Fx32hTSmE2Qkav9XFLlXYVkAxc5b9A31e2ws1rfDuZZS2ZL0
KfC92z448rVfDjhsTQ2kJ//nOjjI37CLUSBvA3wdLssD67J1yKamkH0xIxpu
9WjQP6oaWwA3JoK9xrzM5Ua/s0GWv74jPdFpnttZYRqQ7iaUeM5KJ1nOPXUy
KCvkW/dImISWDw0jKauJoMIqfKTlWqaNt+iFnpkilmIyq0WXgs7pX1DZD8Vr
Oz5zQochuvFO6N6SuR9dVSzxBj1tMiseXs2irWNZ9sHwBTCBzU3wKtU1nFYT
hGuGIzG1rxiawNbKqTsvTxvtD3SkDkxIDCq4+NfWheT1Zw2eCo5fmwny4QuT
twi9dlmyP6J3E0dk6riAPZY/y3LUAVYtg4Vc6ZPrNW9v4bqW6sXGYz61eZp0
/NvKByjfT3LExMab6PdpdjjRprggmoc7RPiFzWxb5ZcuwBnghsPx8Fatud7A
ZLq/PAxKUm//revdEToQx0KjHXjd21/e+W60V4S8bRWznBwIrPgvPRAyNQXN
fyd/LherHRraBCY2YthK3ikymrf2VZPh53e9TGWUoeHRH9gEZb8Xl9uJNEkG
/xYjR9tsn7bLT4ntg/g0N3OgBHvgbmYa6Y/OiCyw2Vkk1fqcEF36AHilmY0/
1wFEi62IfG6Uwx5mXkChWgMfX0hpRpAIve2USZGJ0tdE782CaU8B6B6r5+Ta
5feb/jRjW+HxZDE2lL9Vq6BjJxVpM8w0zSX+z8+LIsdelEmLxzW/rz+qFWjS
3oVqtc73mGzBUKEX4HaiYRBESE6HeOwUL3ymiFj3Us60xEO6NvsR19O3AtzY
CEfn1PbVvma4b5JMGoHgp527bgtLPVIl+CuPidHjQ7+VPWENnfvUFUwwVcjQ
dVwnIg8k+jtPbkSdEABdtXh00IB8vl/LHkYohemgC4k9FruWI3b4KusXFbFw
ixcYMqUp9Gf59ZY8B1B6ydAkJh0EyjffwDJikrW2zj0Z/n+ZzcwAzjUR4edI
fqO5cohJ7N+ASHlu/f2dvtqHEqvcyfUQiED1oKiunK4TUlJJMqAU+9XsxIq7
/wc65tc6pAV8GwwWOO6jzhqBkQVNynqnZFiJmE7BsgZGGbLKjffsKKxTbk3p
ucFkx5ysL36C1OVsKsGRaODHBWOqq4mzdZsPa9fiLQL1lujCyWVyQdApEjIX
ONHxLmUbf68WCRmvLPq38z70kuCLDZobvlF/vms5dPXfnKmRBmuyJbjtlxQk
qqcM10D+5aPOg2b5CLRGRSK/gUwjwv4KR27O6scDGKWZqMv3UY0LFcqGVJor
+XSHo/+EWU8UaFf+zxgQscdVSOcqX3MFDxi4YgqXwHonm7pfUfdMCLt/GkI7
rIprgQM39bi+X/WRTZkWScjDjDxE1VEeSeibfPM5rnTKaqSttSYxDPObc1EV
62rqusE4M+wqAjvgOTHL5bUJdjA65oEF652wiApw7d905LcXiJAYAroUNf++
K5Ugzm0ahuAfzozNv6wJ2i+gkfWNEBLv++xwJGbsPRXdBAv8wSgPPbnDAfbf
1HmgTRStreP+VwPVdV4onSA2Jf6WGA7RUNX2aoGVqpgDG7fa663xk2AyTSuI
5PWW4SkdTd7B06tW+T+n5Xg2/DXPTBKgz8R9/Bgvg+Tb50EkvPCms0qhiaAA
h9MMbhlWArf0poluFFqE8j+AukSvVcRq6VW11U0jdLAjWvBxVrC7KpW/R0gq
CzHquENTozcyA+sd07K/6D8gfK9sFRH5chP1Wy7HbRVXcoI8KMUfdmkpAB1B
YKr1azzSjbert7HZ+c9bcOYzuBsS+UDD9/iWwspNAc0DTM7EDk6+hs8rxy2T
fSRN7oYPrCXinDmM1TcwMA634zOgdf5BiV0QdBAdbgJLDiLQO3nOsJ50n29U
46DDYSDsy7B8XSOgtnxRq42Z9hfb7h1uPXHN6AqRfQ5ByLyh6Tr3JolBTqBl
afDH7hdgjqWiXOaePrLyX5VNPa3JrG715GrhVLLorq/hnxTfe25IVRFMRJot
Zg3KsTZtsNxRWtBJ4LAH9UmfAMbf05oWELTEVLwuhHzDYsl85BQTCqdoHIVi
i9iMpVdfeJKEwS0l08DfK+j01QylrOYn5qhh/8GWyTczAvffcu/cFq5Hczgi
tWKHjEgxN7TYmw1Lbn2E3IEjdYhWYsdEAbj+MEcYhYV/SDn5xgPbTMS9nWqj
UJ3dAk9Nydh7ZWe956n3/bbky5p5I0GYlrD9f0ojr45t0TmGwea+Qdc2brHq
BRas5OVvg0Gh4MVKekDbZOrVq7E8H/BbrmpqhU/5GncqNDhyylPaWbEAu5Lt
qOCWsKH2jbuqs0ofXt4Q6w6s285XoXYIVg5YSZQV7m74xRIza3Uto47UaUBL
GuzhgmUqG6nkKwuqN6wRRlJyQW1n2/GQGIUsY8s6MiZRNpkByRfSwP6F887/
IZ+y2NsI97uzD3wtnGwumZoCw/I5TLBCkBjX/FOz/GCJc9Svh8bYQCwWUE+/
VSgs+wiy0UKN0N0FnnBafH8EGshSiavKN23OcWQKngGwYpx67aotgr9ttv5D
H5hNxR8QWuhoXXxSBrZQ3m8f8Y747Hvi02D4OO5vutW+ScAlgy5GckcBZQ6L
iiA20SaeLu6CmF4k7A6iwipW4GBpNucY3/pq5PxZCEwysx4FgJMm3zZfyfIB
OV6tWLDqhwgqIObsUldtTSyWao6vXHJlhElJO4v61gG+tGxFTl3Kvo+GAF53
dxvoLeV1dWyM4qWQoL0ZQPa8t/iCa4XywtVcdveD7drQChiGrZ33mq4zoF14
TPaImnCnxr/QVBOttq7fg3Y15xAYtSk2MhDUhpy8E6WIA6v2m/ym54+eifOR
TCRL9apnx5evhonc/XbF7jO0EGQHYTZmvKHCIMHWaX7is/OnI/IhFpoiqcQv
166r2QkeJS2kx0s3Ot7sc4CNbC6LriFjXMXFXlfmkXTWiNaopDbxViNbzgMt
zBSioMPWx1CbLpUTcx2VVvpnMzYSjGjtsAZqUvGWevC/HLJsZO3ckHQFuVdc
5eb/5Bo6+6aPAy1RPmsS4szw1AUifhe74oqteFD4xB6bXVzsh0Bto4tNcmj0
oBekB6xTJYFnyF7kw/u+SPJNWN1IGYIyJujh59+Vz4OXInwrqNBwmn2jox1D
d/Bm+WuOQxDEwjcXP/25B/LUxarC9lFywOqwVRif7AoVcITxL5tzfBbnQkpo
HonPlYeEgUmxplpwQ9EQebzLW+7fzmEzlska4juJTEBD5vtYCZZ1Mcr2ibFl
BB0OlvW60VWBAsEsjqPJIU1HHlQhpdWtzNYjF0WP0BCPum3kMN0uG/VDpB9E
pLT1LWtMBKumW9B6RxziRfgP+amQbAvwtjbZudctOrIHA3xigTF2R3Hz7LcH
tBT3/0BG4RbYmxzFFxCUXM8WdvVPd4igbRZK06iZzB3JSJS25UAZ88FU6g3o
ZD+YlXKQBHgILB+FL8ybKqy9sxKlmQvjcdVL2d+8zChxEd5Qk23tRklpATTH
lYj6L9brV5A5PiXEaGE0wJ3QOOyW/Bs5bsjF5uuv4eSvvDAbALVMpTPpbBuE
yIQnT4yJJL4lO2ZqNEjvWIKEAo0dgE2VIWSiQ8pV3+h4vXzfvZenhzcIMAyw
JfeF8aFbg6aC9cu4wHE+TJDPZRcH5hMU9ATYyCZHoc9lMR/KX2HXpyH/t0sF
Petw9ZG4dojF8LrTwtLOKImphkmsvMNWURE/FkRmPcqmeZ645UI3KhzA8JBE
E08vQWbEW8x/6MPIUo2OjbkZktvPjYcUl8Py0RWBXKsyyoVX19FkEly9Vbbk
nW/sR2/cPaW03fZoxvOaRxRNnNlbDdfDEm7tBv0o7yCxch4M2lpLSxuDMPc8
73mim9YlmTdyGajB2IIHyMR6vj16ucw8jdLof0fPSGjcI/8IyFwgqqyuB3BG
/08IeksgiqtG3g4rP5pYsKsKrloWO39DBa5cwYFUoDYMnbdouJCWD+9PC6AD
n1GY/JS636584DbhWpbM6pwhZnqqSnC3qaOc1Axz/yD3pmrftrexyVKlDx1U
r4Bl1nJQGWwrpgSzmE14TWtnXjiwdP6I+EZWIKZ4foQ6idgSLB5lSzTZhvz7
xGXnUfJ1uUoOzIyIvfDrn0zHzMwUYy96+qDEoi6WJtsTUpQ/dDE+pSCc5YYF
VHWvG0DTgIpvNZvcgMz7XPBV7g+dpAb7SIOCddezHpEuAHo2NwIVttBkKTbk
V8hEA1EsQGRGndWdWEMXO2VQJaHw3s2B2PYIBCUCtPp+2eG8dnOLqUHFlv5K
4KezbibutWTSuz8QJqLn0KPXcZN5SnanNeoe8oHUVeLq7hbGTchRVkHe61wt
krgcHxtKqXefrBSUP/gJkHe0T9NiNJ+3duR3fVRMIY3cDdjtAbC3displzRr
ndyAA4LVtySY721bOaKoe+2G8EhKRnE3NKTushsjKCm2Ctde0O0jJ60DMP+w
xtstpycDpdwkwv3M8z+qBk9sJfmN5TuM4Z/VRitjsswA3kLJAjqxlF7HkzB5
cFY9N4PUInKWlH80kfrVoJgJhjXEfI0xaf9pgOnBvPqngQkCfjC0tP8d8c/z
6hnco4otnEUHZ7g6GqgvhrFgueq8gkBBF9GZdyfb78cyliIolKmxffyZ0JYN
Ap6ucj1CMvJ1K6Co2oL8LPHu4/a1s6Vs4kaUwA9CDfSVEJB0Z+KsQnINZjSw
6jtu/gtd7ii1Z3iDNajIfC2t3nXxBYFIF7dqFNUfZuMaFgont509LFBxBTib
l1Lc30C1qv0Bde31XrNWlpw41Rsemia4acpl7dZxKRj7EnIGbqEjJ410IZ8C
z7KCEtXrjbJ22mccI7vs3q8Lm15sbBtzo3pVWbrfWNtxlWbhXGrSpkY3N0ph
n3nA7WFR8JCekoHFytcD7GMYbaIgJP4UJNpimrFj/lguc2OtNrlYg+hiS+G6
WEjiRvVNsx+0xqzCHabqf/KD5WcBLjl7K+hWaEuKnYnsu5eJm0bxujzIkP5J
QwAlctDe/M7xDF4LMLBQ2feg3DfLSU2YjB1QeBI2LCUNhxIKK8X+WzQVCI2A
EsbLvLWWjGXVFwAf6FO+xelqw24EpEVDtVGVzo6p9LrkUcwaxzWDRjkZ39li
PZ1emxpSSvTR1eQslnSOswDm5LLSKWVGYkyullele7mW+1KTkxgRwLyyghPZ
dIIwivmpGyfnsRYTBHP/I3YnbKipJtNAD8ghPj8zNrKb2JPqVJWbfa2thCW+
xNY+0Z+cHiOC/sn/aMKRKaQQ43rK9vqT1a4TtefuZQ2xyFj9QukhAz7v9CKV
KnBUbvqwX96p569HtxviKRtkelNGy5gBZOM7m7OFPSkTurSFhvOpagwqntHT
3OMyi+VHUiGh2PkiU7zKOzsoUeZDI3GN+OlLj/BGUgmCxDcZLiJ9XCb2xnHa
EA43N9ENUAwFWDl7lxqZ3VUWFDlG8VF6h4J631l4bVHgkKXOyf9zr1hlymWU
ebuAJM9HIRK0P/C4eQSZlIno92ouOaXa8C6UV62AqWDXwx/3aIKxllp38LV4
S2ROGmuC9cwAS07XEXaQFJB9c1bzAvcRz4h1yK6ltOUYP2f+zLK0q8vAeqcT
Qw3629rhFxEut8yAyQWy8+clHJk3LsyVxrRaYwv8rZ4jY/940SsiGY7Zv26p
ZztuWAfJUswUu4gd5bihvLEHTpMAmr9u2mNuhvJ+T0Dhv2OXYbYPkdzscEnR
DeLkPzW55eLR8SoHN52R2fMKGG2XJ2X9JAmR4NEumXzki5RJlpFR6Vsdgusb
ErDrRmmGu9Q3lxJJCZQXng5QkXQ2K/XX21vN4U3TQnCTA8NO157d2u4TMrRX
3kiJAHmCYYZXXeIYdOP5KXvqwALXKXGOk3hQESgXVn0I2/Aak2S2KBgembpk
RRLbUv7DlbdKvOCDuNxN717JKSP25Xb0gAhFwz0mm7eLDE1ajnw1B9Es3e81
VeqvGBgDPLf+OZbAlzCNXlV5NrQfixHC/78IpWg6gBj/phphUMtCL2T+p8a1
Q+k5YtheftktocLcq23l7lc9Fd10rxOQwqsr0qQ8CtapwjGBqfD+T+611mr4
/ZUhK3IguFtlLe7e5rVfcPMGpUtw37yA5wPcbAmZtx8KBe+z9tHTc7+XzHl7
eZvIeULbJRBWZ3xvOYs0Bnnd3y365rk8mwBX4Ak7mRfbiLufkuHXU+qAsQ0Q
lcoHcruQ6so5FirTsTpvh26MQJ8JLxoewdJy4JDKFu5qEC83TafZ2IrWVHEy
m/o4ofnAHPIvjAi9Yji+ZXnr4fXKUp4lxe/G8KxIOXDa82hzl81FdDoodtlR
WZdlE+P+unnuJXpcG7ECb6/tDPaou6nV4Dowy7HcMMP3mzt7J7a7aFhiilB9
dLrBFnQon+ELFl2agsHqudnDlsiBugECgeGyYVlKqeXyvqMSK1BNHB87IRRP
44hWbnVGUD3UJeERX+ouG1mucCg6GPt7Q0GGJugdbOBAyhBbrFMC4Leq1f9x
Hqixhy/2Wvt8jhX/2EiVyCKYtYczlfZHpzcVrpN+kK8odUUNE9oDMP0ydu2D
QNlOQQOeHN9wyYcDBQ1/7a+VzJfXO+cN3cDllfnzrUPxsddeFwQD4gPE0dyJ
z6MnMikso1j0sfprKyrqHDc+OPDK2p2IjWuwX+XEdwQex/F0aeGU5UP7ZuFm
P7UYPo+lIAslS1xK8qGDXpWFRPluEfeTkL4U7uCEqbo3fuGMihqOf+nEX86X
9GwjfF3U9kuxSrw6bG3oT80ofODnObHJzkAQm5Tie/dMAOQE8gAxkOXUMCnT
Iei3DZelNMLMT45draFSOZYeAERYtK0z4MbLts9b6+b+5PHWLVJ67p/TW0jM
C0Qd5uqwM+b5jTkyWPFPt1hKpFrqagjEnfSPIieCrkW4EuDFfraeMgDYdfsL
X7353oH2kPvWobnuBV2Qx2KppuBbS7qPpewViojCtodG6/xP+skaBrm2VCyR
5aofHORrVldKKYX2RsZQwMBdg4mEmgJ9mJc6KExHwNXxAaVyYsd/GlUCwQQa
02Gh0iL+kgoikby8rMhvc5Cogq+mrTP90WczKte80+7V7SadvK8RejXmkrAo
I6N9wD8kEY+eItLH5FFUPIHH9H+y+NWhz/UNu9VNmerFnrMmg7fWD+uXnnpN
KByj3e+AabHvKNdN67lSO+0z5Myt+A9/yjxx6NK9GmgI4EQACwLNS6F9tbqo
Fnmf8Qq0xTz5gNujPiVSxzvBj/9A3NCpqqNpmTGg3stUrx5Rf5ak+e8ysvTN
b6LKD3DYCoDtDU3oF5aTEa/hr2GTy/TJgAtMUKUbC+LVvRyPuUKV7TLFHLQ5
RMJ1m2UjakeUmUXKTaT5+RMolvK4gG/Ab2zYoyYPzC+6ugT4fo4nDlFAscRF
uURDmUw/21QsabCAWsAD3kCAhM4EPCto7+w3cVSS9GWbmLeCxIMT0TppIug9
9O+7opiwbqBAHh8U4yf8oMmt215Eiya3hI/DrG7b2uU+A1xx45xIWs2WYwDm
ZhEa1Cb3Aq/YwWxGmv3ULMDaFWihuwQDKsqdLUnEv767GPBlt/P7ocov6j+L
h6hXjhuo9omAKD7YrZCTIJKsuTkTu6E+LL0afpNy2cLxZbtnHC42uyNtHijz
L8G+KULjl/ag9QwwGk09LwrFCaNIc73f/GlAqh2Z6oReWYpPiozoNsHIha6G
/2QKIsFxj3pXHO4zNRPIkbDzUYNRv55tp6HR/S7X455Z65UXdZwxXJ0mMRwt
+4gyLUB7qBzS2LWp+jbQv/5fJQTv8mfp4cTbLf/oUWiyBgP5rwYeE0ikMqjp
KniEFBrW3kONbWc1Pw91dvn+UZtYocJwTh1w9BylrVXgGoNDC5haZvhlzDqM
A2+c9iWU4Fm2b5vrsC0gyMLvfEFr+HQX685+/4mavgfpP1mgPPZ0dXboTTTb
iPgUlyJYZjXrAdeH0o6sxgqgV26p1J2kqjFVmtWS+a8Dkwtc7JcE3VTw+kqg
+9uAkg7VvZbYVwTxGzGGAdO/CvBETAupKJWmBM4TruvAFbnlAdkHjAKn2z0E
NVDZsFzYH4H+YhHuz3/1E6SDgUfCdY45iy8WpGzn/E4XsclUyf/96Ayp18KJ
eWrmXI8N/pgn/CprnAesjJFzuadR7qG2NC1BczY5Zb8j/JDLBupC3KLmVGJn
t/BQFrocAk7hvX5IAdEiRyaQ4s3csv19hjAf2sly8Ka8/Vh+CUzwZyMcifdx
hVE8katJgmfqh6oa0OVyZixgSxskZARPJ3WrVHZG7HeXQid/23xzQIzM17v+
Nm3M6ayd7DJfc+56Nzs7NIMoOLMZPEmJlRKJggrOPNAY8AKPHJQHCjDlCFOn
gwfqWzsltHxYa7LsmMc29zR8/PvJ+jkq1laWXVA7S1p1jOwLlGyXzV2dl2oM
2LIjH9/Vs65jxAmVeBx76VDhqUqrnjwhnT61O/6t4p9TG/7ENMULoOEKjHBV
LtIdnxYKThocS84YuV7hy26FqUX3SwFdouPJJvRVA1ncsGh2BZ+VDiYG4Sdg
RKICNYJ3eMm4aRZnQEEbjavgUtdgI4x1Ps3+wqZNwtSDAy4rU0eLZ86cHWBp
dSfhtX80sm1hgBN6rUxwbJJ7BuadhtH7/XwOF6oOwrf+J7BH9R/U4MNmPzGi
pGTyiABvNJb3/ZTQfgCHhnw7ut9RKNORb2xAmzGCpSzR/YqA0HJLJeD3PLOY
1zE2oY5BC2imTSG7MYV1fzvKT/Z0cdQ4YUroutKB2eJF/9kloccIWvLt3ipR
CePbibUjSz450R6V7NqY1/bUdnvscHw1aO6dEjY/4xFTWYTn+T64wxvkV0KQ
xS17sn8EJIfibp8cVBlsYrsLu+aHaEHrc/4koIjEEY6IxrMaPyZlHSqJOc4Y
eMHTntD/bd5WAqDcxuwl7T15jaUCujzetFhFbmE0W3wS/rJ9WMsDeNvp26iK
ZRp/o/+dqAKW2DU0cowAFbVlL1HCOQDomf5M9Oi9t7xbA7XutBl+HwwWYal6
zEbsHQ2EqGsxaV5qjl3Dt/PjKETWwSy39am02lQ3ofHWr48UuEhoad2B0DBG
Q94JhIN/BYINN0WHeCU2kLtdFW4C3+a+N+3UJWjtmE9hJqOX5YubLX71tgJP
1UTCE9e/3Hqe3WW4JFKKFVb/PC9Yh6qnV549BF7glZB1iw/13xA2yUVP/cVE
4T89iywytkpnUcuYJsUJ4YWQlfywnILf1PQgYg7fi937H3Ahq/0ftp47V3kU
xOIZrit6J6V0Sr9BhxQ3984GG2W4mEDdC2voOrj272qO/2bJEgm7DgIv3jjS
BWSvthDyEnE6oNf7SRlwRdYdrHfx0fFeyIkWR/ylFlwn7lOlq7unTz7wb+7w
kD7Gyr5yXtqcVhlpPae/hAj+5TDTzW+z27Q/Npjm7NBGhEtPg01wQOb+Pc+Y
JVdjmpb25/tN3kEz72ePPXgh5MAa5h7ztRh5BtlUJgTiTsE5VWk6qWbqTj8p
0SbfZxHjxt5iuFjueZKLt2N1CSot63NPzEnPf5f1EfjOJdXKG9ZRnCNQcjJt
1tqVnIbVgLKdrfVVb0fT/360zZeGzjSHklHALmUSTh3TaX1LsewF9/PhmzLC
nNCbsl04+PAzt7vwYpe83VazI/FpOHZBiFVCgKU8klXdiarKJe8AWIfjOjTY
nxG1QmFUxuOD5KBVLqNtNSDrQrwAQcQlKCASIipcS746D9/z8F/ou6DOyEX5
0cEy0qPe6VfuGME1mmUBfpEFTvbLJquvREoTd7qPPL8T6kdWVdJ2BuxwX+Ns
3gleQ3OvLY4Mxq9O60OHxXSSheG6LHNsOdKUjEsOQIAMTqJn8v1U9QipQ58v
SFT5UCQV0l7UU+/HRAqeHIID9S6Jq3ZGJK1+HpdeGJITM/uxSMzpMUAMhswg
rIH/Uquxa0s2zTAbGFR3zBH7WuYkR2JxtmSF+boqAzs5Mns1R75pGMzqranV
fhQ+gGF1g6F4u+duvBkQr/6huHJzq2W8+ZG53HoL8NLBVNxsqWw3NgJdJ0DX
HRWlkNa3aapVCM/l8WmWtC4kJtaqWjY838MrsHty/ALIDuGe4EsS9j+5fsuB
+HcMAfoSylTy/6l1THZY3u5ewdrU8kN70cipilgnkg+RfrRbwVuKt+5xwL2n
mt7tP9JUpmy5jIyy6U59roGEd3gPmlgJkqooct1yVEd3Jhl0x+Y2mTMYeaVd
iCxIEgIoMxc1TPp2whqsUX1K3hCU+o+yJv8n/GAetL05aUeUvPalDalfx63L
oqJ4BuTpYYd2nV09IKNUEjK2CD8DVClyHcA7KFHZSKUmZnghrYGn1aR5c//R
SMwZ7kjye0ipc7ZIIhW3AW5E6kHbhCTC7uY+bxOGv1yx3bbzmKSUO9P46ADR
BUnw+x5lT0Q6cWewivUtVIbIaIFL+VsRMFL/6yIGvHmQCT7JURW6GTJVFptt
M2wIJE9Ay4zf2YonQdGSfZzBHl1dMKNeE3CtcPLjM65GQsYpB/kIte+GErFe
q8bZhLSz/P/4tfmr/FgFh0WwoBU8xqEPgsfxStssw8gCC3urzxcGZHbj9qYq
pSGGtNvMjIpXlxFbuI5e6TZ8Ru8utpmyl6HjoaK6FcVtpI7hZicm3MVFU6fD
p7e3SQ73BtdwRs7o6kQ/YSDPb+gGMTrKbrGyB8XSMup0M6iLbGbSwwv9cNaa
FGO5AXAOCyN/ovqIrlLJzix+gOsegu2I55683+ydy9j0ucfRtIoNh7L+KmZ6
oQy7V5RFIOBhyHigTq4+GiKH67ic2VAh/MDRNYJ3BcKLYkd1iz31qXL33PKM
O8boWol3XvVdQ688o9aAAuef60vUegvhZg0V3L+parW1ZlwplFcUzaNJJDnH
AGBv9VjfoUB3qinTH2LvTrptxZY5zioAroOtlGHWaPbzawcLWNqnc+kqSWYv
mdLOYHiPiyEDGLsSORPVcwHAioJipMMSA5Q/qV0GYZ5u2L7Yr1HFLjF7NbSe
wQh/AIZm+auT8Q+W2Jf2nq2TFRli1EoP7g7JCbznw0u/F5S+mvPQNYOB9vXn
6nEWwYe4RyyYMXivO6FSi3tYeIaTehQwq3ad/n+R4Bvz/L799kcVmcJ/1lGs
N6Syi6vnKyoSYBtizfigUV3wKrQdAfIoNJbBV4lHWA7kdbjbZv2c+cJizXM9
xWf3mrmePEUc/aK/ULDznG64J2MB2xyryxDSzCBAz/a3PqQ02zsgqe/ErTre
5IbtwwdSf3ty4ZrFskiVprczOwEShgb/CThSgZ1AmprYYfX1LfQJW0qMQaVk
ViNn5ou3GVHIQ4cMHxa4GyEtDZc4h4Zg/dWew0P45Zm+VLK1iDO7nQCp76MW
zjIXw2pwr1cAtUrf7aR+gPV3Dd9zW9qbi9XGgnDWxHpdZN+WMu5taOzRxpTM
CZe+Z/JXOXpiaytdIuVN5chWpkzcD/Z1ZHx9Bf3ppUseR8vSKmAAbSsAMHmV
ZZK33ZdW2CNpmTS+YDQzf5NPwWfGeKK4yWS6dkUR4A6WPA/1MiZmjjXj5jTG
9vzj9eW5JpgsQjLi7o1U58hrioWDS/NY7cOwFhC47hDU/JnHEP0J5H3+Eiqf
8ELR7UHxyh08ISbJA6/469Lq8vibevSfTuR1UXl/sfKJIaeACN2rF9VZhnr1
dcvK41GlcZLl/sOUmGcVihuOsueN/A2PleB4Te3arYISBdqeHPPEjL01NTcg
FlPsvbduzO3dM63Av9JPeVsvIH1yUEiTsxm4bz66xmG1ExBiAuOsRm1KAimy
Zq1kylbd8tfTOq9WGzzYqVEoiX+yHnmNq6w+J7rDfIOzdJLbtXMlTcd0/OAA
g78B5O20zx5QyN9wwntjlDVqQojdRSqXX34ELAB/rg1a8EeZXfMqqi0rVO2E
gYiqB/Xc2tgM0wsgTilRUFzFEz1gqfFRYkBH9szIaqtcyjWTFZMLPVCt6jYB
C99Z7gPEhjdIoIkjJZeiWSeI5ukLxKuHa7JuWqGN6jWSKNTyVneNqM92boR5
Uh0fUi2JQTK2NBPQuNLaP4x1PuXukxelpAfLb6Vk+LjMYctXuCj51W6lrucN
bOSqlaV7oVA2nZromgCn+64DvqcyDix7CItqA3RXEQ0oF+Gwgf1QO4ptanO+
rQjuurq96diHC9Dmx95j/AiToo36M63hHmnPiSmdpAr5ADRyyp4iIhlwBU1B
WwTXgL796xSt2mHJVzHQsBfc6WE06L+lOtm7Bzts3bZy39Ly+bqL4RO9t+UD
xUzjsR9zCJ8gZVS/c2xC6+tMRBMsSLkyQ4a4lUL4ivU9kQT3RZp32n9bvzrU
OeZnwVNopVnkznThh5ljSWDXUS3wf3WJTOlwKot3dW7GKxBV6r3Me5vJSFv1
JWUs4pb/eBiCeW75hVzcFSqvbM1/deuOBG5/WHMyG87SCZ/XcxCTsy56SxzS
8LnADqqftbX2h2uLXd4RH9QNYlZ+aiR3TFBoERDYXCOzuJlJmqml3/KxQzXN
TD1HjlMPG08K4m5NzqF++POZi3KmtfpRWQcHAnLnngGKDn2NuUFEnNUZscfG
3ucCSbW7+zviIclWp5EyOKpbIMlAfuXYkbkJKhhXwGYSqEFgNZm2Yl4hU5LP
98rbC70j0QURwu2gB9/Md8yDXPiKXbFWLdtgMBlnpCBXtre5bF5lYotNw6Rq
R3A5uoh3jmSiofjKOSfCoE2+K7obYBHGJOYzx9x7ss89/zA4AyqkcMB60tEH
kjEY9S2n2RhqChEV7UF9losUbeBgK+CT6sP9mIzYMqyIjkeXQdKSaoQ1FG4m
ScHWxeHGpXZDu5OFOtySd9KypfIDjelCcI2HVe3sMZXHMjxcy8LQbTETj6c3
dRrdWkXGdwWOIsEp+vDHFS7axCO5SvoqZPanY1qrZA9Yn69sUZh1SusZJJla
t3uZs1TLc//S/yMKnd6t6VOEtCpWvOlXEyHQg2BjIKsrbQ8XG15M56lgiXJ1
qwn5vrgYkJOWsGhg0hac9Rysn+EqemMEs0JmAJAhNJe8NoTNugaujOb1v0aN
MbKNIE8seM2Vlvz7AgcumUtXCyVMjhvJ4Ducv88vxQo2SRl6qw2ZnTTNSAPg
7P548vEIrc2ZmYhytIEwkw33QmsE8+dolFxtiqA4NgkgI4RilpKBeasBIsLK
CZSxecrXuofKlHMT+Xc4Z4drWPlyvD50KYmW+oFrW/8htcNflnSjiLVYfipf
WksAUx5VL7oQRNFoLHD7Sx0o4ZD8i6OtgZ4Al43wWNCkdQTomdsngOpufSOz
iPxwvLpcff+g0Sq86iOyOHqtI89GYXtdSRWhy8/WsyaNxT7nPxUp2E3h5waq
24jMpQx9kwasWdYO9Vbjx/8Z5W2S6w9URc0VRL4CQIpi4zyRL+LRCY2w56Je
vAhGNyf6G04i93ynxUb3Ov4rMSk3gUJTOozRWDHkrslT64RrXAe9wloc9Imb
LPXuFPbZFEWDOZgN/fTDFSmycVfYIzrAbcD2+Nq5EZ6R7Y8aFQEAZ26BcOdp
FPqcaxTx6fX/gR3AhUrwebIvZprXTLK/J0EK9XjlOlDSAav1GighHKhNIduD
lb5B2H9gq6DM+QyLGlUhC0U4omKPA8gp5xHeTXkbx9VE2dNMLj8V/KnbIAeK
9SNOkaZxLRUVnuJLkyKls/TkFE1Vgg7P8loap8xgI6IQD5QWvXLgwTQp2Q1e
kcqSlrzoTKTRRr+HHkqZ+09xjc9PaF5jUdpA4y7KfmKpe6yg9BU3qMLfuedA
9AGV7rUKtDblni3zkJ4q9oy92TrkzUdziIKzGggI+a+PshLeED5LJ1N3+N4G
mbiB+JxWoyYVGMbIlUG3QkeyQddBl3wJUKMXPTEBaJoau6crBZ6bIVzwvJkn
6UEQ5P0yDxsP6skPSAEXR5kl7IQK99FWogHACLH4d0qftraLpuDhxjmy8b2h
npBLBz7/5Xp57t0mr8FgfJd8et/Q7DEY4fdPWLreMz931ZmqPa5tXlhX411w
TEl39NoUUNx90TiXsmayOl8om7eM1CrqYE8WJXunvPNzjzhrrxdY0s0VcRQJ
7H0MHs1jCfqLSoaPSMnWj0s1tj+l3Ew33ZUJZFALdMHK3WRGfNbB54ZfH0MB
9GmrrFtMQu8hFFckdlIk2l4OikiaQLOv582GA5ecdBlwq1HyfIxc2h20vxbO
NPCuM125BUcDm4ryu7pw/9xDdd/16TNjTXMLq5Ns0nO07YmeZL073e/pj0LY
b/It1Gw3MayNu2RitWK291xnOHak2xFOvfWzzjotRYEVldYs6TCjo5iR8ge6
VYAtfUrUZq2DfAkick1L1hbSby6uql/CkUc19+Cbdc4CNq2TysA9eo+s9yu/
OxFuKPbla3DKDO5XL5WSk1NF9E6Wfs3rDvbaowdwWELY5E91vB8hhBNDSWUy
8Y5sNwtuv/Kg9O/BdonPBEhSOsfKV/c5PrXC13DpeR0DY/ymlOQMEzV/34sI
5CAyRFahtpZVncXzqLhjdEZz/CD1Bi+LwmK/4RFOTB5Wqmb/0TCUdA8FAgjo
ecfjHi5hoo0WTa9WbLW9d+ryBGjljDE2j3QpWqBVVquuw6Wt5Ce7cOPyp34R
Pgrg0KaSCYD860mOAL/Z/6BYeUFVOYsSNX+Om4eeQdAKNzPGZ3SI6iWGobme
7NAE2Gb3Jvjb8VNLkGpUhQ4WZBXCWdQX6n5H6cu8pMOpPsGV+W1px3AaUB5F
NSKRt1XHkYL2hCmwaDUaFtIh7lBpOmkPPmY906zEdh/Eq/mUa01noflJhYB2
kpvuRgzCV4gN0wGhVe/+eO/ATDnjVM5ogTIcCMAS7by3Boi3wNxnCJN7kGIT
VomN/OjPPEl2ggR1Z/IXHbTH1p8bvBnpgwJdhYqpML/RKipGuZNjbEc23VdZ
2mLSPQXu/V9al0SS/u3mc7q51fBHD292zeV9SBXniSojdwtNaFv5+tRO5Fc/
HXoNQPF7ObKrxXKPVHVt9bKtm+QQIOn5oyGpwY0BB1+YIl1It0m+ULMPwgo5
Ln2tgjW6J6gkwZz7sBnuykP6DG9j03SHSidkg8ruTSZxvSSEnye/Ovf8NSYB
3qFqHK27W9mbZiMxnVSUtwtsRs/cTVhH+hccG5drLNUuGufpOu3apGfpRmLw
gjBFHQH8HP6hGszbDj0/bKC8d+cgSK33gjaFO08defeCFOmwix04opSGOioe
vA8fbxaq5V+iXYNWP+oVSoRJkh75HeLxOKRZsOZeZy/YST8wSxzfLMXfJhST
6ZCVmSqI/fnsQ3LlDM6lB9sjDQ/EXELfDGWrponE458gQ19u5GPJ05rDY9Ws
l6+sfSjye/klhSzhE7uYMvBTKjU/1gpjSYodxqo0Mcz9g2IaEd21y0yDJnRj
QblRcFpXBq5XqBX6FkDFRmcBOs1GctIL4MU0DJaUHYcoFdVKJPomeafrIg+T
QvotzIa9F9hO/dAkh2eK6/s8793KkVJaj8aNIP1smedaaNdnYZ/IHjuYOSDd
VE5HxBAlysr70pZM8cY+SsWtSZ9sA6XjRrSePd0Uy+9tgukvLrQpPv0Eo+hb
EG4kFx4vrHVu2XVAGBjqmuCHt8QqJiIKwgN6qY84QAT556lvJp/F45/HfIv6
lR60xa5V5RyocXHU9fFDCf/MmHSY1Ueo+zBNrFg3eS3UXyXDxprHrDdCLpNx
2bZhW5c7PJv6Gv60gooW5Nigu2DGvGmclxbnMFdBntyf9zVvNIv/9GhdwL4Y
psHahX91SbPWbAALpsYM24yrqzb1oexMRQGPU2QIUKShzm2XhfaD6QISfmzH
rabqFpPkL7dxhbbuMPKky0XNCYxvsSgkk04odvf/3lCMgjCoovOd1QbZFWRj
/zKEZX6C2/ku4bE+WZjHZ/gTNoY1sHycfcWuFvCJTHucemKoJmYgSdZK+WRO
hHHckzGmVBrcM6rt7Mn4TBQ+L4k74+i2TsaX4ehy8C6NITfu88umesl0O/b9
rp/1yDHfGxdLGoVlRJ57nntkrRMwIsQtaWEOsqNepfwm8DD7tX187pGEZqqI
mkd+2WJ4a1liTrcZTQZLEGAOOgii7xLs69ABTCmpMM0SLpR1LKns/bUdnPh6
QrYJFL081lMKAx23WRgwCJzD7jYH0AJ8uQ0Ag+m9TPwd0TVJpiQlfChqf+Kd
L2o0YyR9lsDpu+JonNJ505AQp6kUrttIdrq8giPnWMT1ISp+9eKdGS/WkeHz
bP/KwRnf0Vd577Y9vMe18bppQcENMTtg5oAgifvbb1U2lKm5Iw10OB9Hzlg9
H7oDrVw948H/z3fQy5/2/tynubA7dEp6h30Ad4God2knaBZlKOOCyI+FPqGJ
h1vWayIWml9VS40TdjP/btnCQwCvNTSeBrcVl16mdAXJc9F0CZWj6xZgWjE7
a+yEoMHZ9BYpqv0c+6eL7jXT4MqUyAlWzS3a6XXe5dvFwjO4G1iW/ZW/QGoy
ia9exRNmivaq6q2/y3KB/CahRxFWDVSC8Nr1sFk1I+o+DjWI/kbe2Rce1acH
7LG7bq+s2YwLPbjpD6XBMWJBOtkW3Lna80ILRWWxZ/vuqWkEJDkW8+qDSOHV
Yfpfx5X0Nx6p3RKOti2WDu1/0K4URVtY0pvaDCIR6LjvS/Ts0usRnEOEPL3k
8/+wgX7nGckY4YDKZDUHfJceb1japAYRqK1WPmaRF3tuJ/imNprc1frgfGXa
M2KesVmmKHIVEEJ8ulBC8kmiXODjKDB2VUUrjfzAWUMZ1/8YTQRAtaNW2dRS
sBML7+44gTdzWDgi5/C5kL3PEzn5NTOU/S941JZ8jiS5fIc3iM/i75HoyPgg
HI3bIkXcToHX68tog9D82JHBAX0lJg5tfd7bgemWs9nva1ZpKq3uT0YkNc+G
zftw7wOCu+iNWmWNwNu0SndGT13au46U5OBA6u4oTWHfpGYkezlM4tW/5695
g2MmidvdvJghh3GXQR5unsDVEWn6dTX+XciAEQzBqsb8BrnLTYUajnKwNeQK
xSGVNBmbRG+l84UUc6fzA+8uTPKQK32VKf4mraiPrbKRviNyE3Gbi8rlT7IY
UldpwaGbEnrdMhm2EndB8TD0STbDpzXjyDKocNEARmd/Sbg1AyvGHDOUOXIP
YZgN0fJyJio1pE3FUgJTXtJZsJqIwnixgq4U0UNNgE8E67R2eaDgamhC8S6e
d+Oo4Q7bVF37BxJmIoaKmLz6MnXnwda1fZmEzOk0xRBDOE6Yn3YauE7PRLiq
teGRvUpQrsUqpePcLrKcHzPtvWOSnKgEKZ0KWv95JUhOKONmAr2dH+4DAzDw
XpGznOYxcFVEv2NSueI7VbT2GmmWPyNV46FjQOwxHKW9RkbLUF9LERcBK7T2
RfDoSWYY3fc+oV8HCviODpISrd3J5JJc5Krs5AoOeYcDCPr365INrqZjswMX
mGbbp+3swE8PNMBRzcpkoqhkAywan9I12iD+cXsakG8/Q+AUyUTaEFlBqGyb
Uw/iHX5zvKfzMFh8WSJ2qJioM1C3eTTXFqXCVqEm0CdYxTKtYnIaThWoqhAa
rROHul2zKkMBPWoGF8vsGIyVKdJqmnqqozyJFOErlpcmx3NvXM4sXMJ+E+SZ
Fb0vb1DP6LXMB7EFSwp4uBoPv8wt76lhmz54HqQSUqKHm2MHWlRPMJk4hxvB
8pCJpT4nn/IhQep0JQuD3uPCo05eSnZnvqGxvjG8Xp6wX9BpWH3WpR3n4eVc
lJ/C0SGJxQiPOLznRR/wOK8nmRWOLkMDiHnhsjuPrg6vBIMWJ/n6k+OooJSg
3G+XG95U248sciUHh1E9+135sc/WCSAwRDGwnOQiHhPVa2q9b2H/OIWBiduz
w0b1jVVG5h0gayntGtzkEgmd74lzuHOxdKeqBpzB5Iwi7K2DO88YstKCXWKc
8pXEicbv5o5L07ddWkHmn/0A43FOZ64OSlSDUAvClXT7l5eh9hm0IbUyykA7
8IswhaeDK/vu5RxMtkLAnXgAQ+VD1+8uApO0+CN96ikEoZ2Aho/vUa79DmH8
cs0Hi1wLyQ6OKixvKifnIXFRvN8LwrEvQf/zhAhCtAkMSRAAqTv6xdn97JCT
S3ct3RfTPoHjk96PJc07CKmT+rzMgsq7P8DU6E2MvzonN844gliVZdU1+fIr
4May9pQ8R6wQpeMdvzQQ7KOqDlHCse3QN1t3Bbw7sxy9DMglH1jzXpCsFN7M
q3GRDh2Smehg2D07gS+Fm3W/v4VRY7UmHHIpom2xUrmrkQuIiEhCbqbnS5m9
+trxdWxaGT43CG/d1l3tsGvPi+D5BFNxCS/sj+LEDZV/IzJNtLusVKJxISbG
NxivLVPj8MdQarlZPXuRJae7vs7n7O1NOqTENEj0jOVA5QeqDeHka6Ek9/YY
u3/RFppb2zKJmcNJ6F91J9WSEJafWgv7mBAK8k4ETQqZekSx89pLPib2eq5t
ybSu2MN5QcZ7JYxrGcKyorGuFPXeZSQsN7Yz1gMyB+zOQQX/3e/X8HULk0bo
OEN8EGE2KHNW65WpoT9ZElUaaI9EO5jZx7wxvCP71SjW2I/szVr8cQ/Q8Wi1
3iJv+Yl0po7Gba7aVkLgi63ygP4Eb/PGTCMR8qaRp8c9nmPUBjp4pJblmrCX
FTu697Xr+6gBnCXDsqjb/TcVoljwUlwMWfMSUCpKPjGRatmPMyDG5L8K+Uo+
0a7ihxBt8PgfjxgSZotAidVFwoIgZc+XMEfc0iq04Fa+mV0lq/Ha4/2ZtVhE
jZ8eYmv18Zdw9m3REIE7eM9q7dN5BkEXUfhUaB9jJZcwe0hiqXxfBBYl+8Mk
o9adLBtcAc+w/NBBAz0el6KZb8mIk+nUR1QPK3Q2valcwWX10/KABjKt8y+N
8nbWsLmnLTNg3m5Ua0Ny6sHzD2VYIFVu9fnvFeRbnySfYfm+44wuQ4oXDU84
KMkkhckQbqKidCc8JlSiiBoFAFhW4aqdLnfvP6H0nDK/rRNYF1bLi0/jtLwU
WEawm8dcmSNW5tNTfzDH9tWBZpH+droaMVSKG2sceiZb83ZspVS5R1opsHqK
Akkcxcf7uWVZTyE+RTk6qEGmomaWNzsN/QZCz47xDPVCPgpHSV5dLfTC8b1d
BFp5i4HzVTW5DokiDQyqG9PSZ9Pslpvt9bWtk5S8CxproKKXOMwIW8JbAYZd
aNyi/+2/DKi0gCkowN97/LCF7MoUSxzHj3fW0bZDeOIUUKfa8ljUVk2hUfnN
WFv//I3dw+SW8wFCmCsO8OLzZPvQE66GUrZvKfyMZolzU8ys4D44kGSeKy5Z
VLHm/P8A4PUpxC6OmTiM/6SbhWA2ZgKrzuVuOKG5sTbQY/Gi4jiuVYaJuyk6
yZzuxmxER22IEMpnvTg4QFNrLQp5nKU2CcnOa2y59iO7OyGx27DSONq12n1e
3f1JOTVgKZ+Z8bYZ7P2uzx4W/C3PvQ4H0+HFpGEoys+6+mWZLOX5Z0bF9iMf
xK8psW2+eKcy6zZ2TppELcjjvh9AeStld1LCg2P8lEppNdNFYFFACA2DO/Op
Fb9dGu2MMdSkuzdHCIgRSc6FpdHu1ScZRywuCi3dPOKwCdsqPmKaaQMGeXW7
PadI6XIrzxzeB90GtSARDN1cnmloxG0gUqAPdddhBdm3YZLHfI8z87P+eyit
W4OMYXj4ULuimqs3Bfl+oM3rDpVl3ePIGWQHgS7svPjRZVlxaTt+134GGsRS
qDKpb1agIduH2hvUr1Wnic6vnGp2xMX3E+bg/RQJlkW4/i+PFEY66b2AmGc8
6K3FWPtiO+5+d8OLgd2xvn0GtHPFTyJgXoLKtu09Kbs9APyylwDIi6WouqLT
jv0d0dXUJgKIW7/P77oJ4tLu8YdaIrcqxD6U6J4RQsiKycCFfPUOhjKi3T5i
x4KbyKn9L9kKh8WCckKUFPgsmJaccXLCaMAeaOMa1e18lPeT6Lo+ouVtsB8p
vqe7BsXmfhqyaA9HrszQFaF1/gs2I+52E+1xaX8je9gBr4pDRt3mhethu4Xq
8KGKF/c+PZwHCPrnG5gRT4Al+t9hNxwCizt0e+SpTb/61wYcpyQpTOAsoS8g
8KVBmOLq/JRzKzBqXz8qfvkoNwXI2Jo0giMMR+4g6amzIWOPN6CD5RD12cZQ
iju9eZ6F58TpALC0pVye7eZgUHGuqNeyMrtEQt//J4d3LeqiUUrJUy5HgKRj
eNbRUjzTNDXMu4YZX7hystLmtjV6USNZGVCv+rp0jfhL9F4zBHTm5H36SoAV
qIat1U8g0PPxDacuajReKYy4FU3dKCMCrDksuP4QgKcU7fNCDVcxBlVkWsZ4
FyCajoH7NHkU/5NRvdw/eTyJ9xYyOtsqpS/UO/V6t4nKp7Z2AgP1ZT8JWC9d
UyeUkSRk+ywf6BCuL7n32zo4NJxUraTEJyKAjk+oNrOBhvG8WdsZjyfF19Hn
BatrkDTFa4qxEauD5ftawbJ1aXM4yXfF7uajqfxmfllSjzF+G01wqnd0mUG/
G++2FTX0jqhRoqfyB+01FGtReAVkaXffFYd0OzvB5HUHhxdOFj7EKJCzwIcs
NfpLEUOHCNhNchReVb+CLJy42MzMRdkd3VSooUB0Y7imb1mwj6b5rk+dt5av
8hgmaPSR/lKX1rl7zSYJ7mM1IQ4/CDOeOfUMfeUWAmRCn3wJLTiEf4NEoKEj
8YEwuUDOnwvoPeaZvkdYbCCt0Ew5uFsV0MWNSqLCAJORrM9dwE2kLUtsu1NK
jUa+He6BWXYfM8q5n5KRtKX7Xn0dcdj6d0Zev63bYFlWx/Lm698kT8AMj+dZ
xaRnvD7r6iHOzJWIJC/NP/7WdzwH9kJwRqVuau4t2OBq3CBqznzgjvd+vSFD
NX0pC4bS1fKO9VMT65MnTfiNGkj5vQxO/OWhD1MWAP+hzOzez7YJrGbnx3GA
f5C84tIC1r7f8yyKk/ULLMNfe5rCk0wNEi78iw5rDE5wUO73EG4RjmmwUXTB
g/pTFMlyh6WsfsG21m6fhrOr2j5b3PMcU7fSwiou3ygqP18X85eSV+RoxVVL
U75uncW6KemBjfwsdo8rtnIRX59u72NpxM2PvRidoQjt4ZZX7WYd5fbKPsjr
eBXGG3fuVgMbMBeDjtycOKZ2uYLfKRKT6sH2h2mvlWZaUF0n6iQB4gY7b9Tz
AV19AFoDpnmfvn8j6Lns0uT8hTuNcOqNwyrQYhkeuE2dnEp69znnGW6Fi+ws
ogBSZp1MHMjpF3P3utG7fE9yvlELkbEkcqRUSQyUW69qd/VpOGR+6xYI45HK
6CZE3kRtyXRevCmHQ9UB5iDDy+LNLprm0cg1BShxGEvi+cm0NSI61r5cxuOz
zxVdqwh59Xqm08cKCWwULxsDMi4zEn8vcNTDkEjppq9dXpYSFUDeJl7TzOvd
0IipdJ5BWR0mn/pglJgW3wKJKzVLx9BlAc0XkxF6wFhE3+aq4/EyWZ/bv9zB
u4CruNnud2neO53RqAdtNMyDMwqXQXj1arLyINGSvl2Yhc9SsqKdO0OF3SdC
tL9+cDdUPeSjEI5PDnGOkrYCiylPh9ds0jd09fcFGIuX/MS7sE8MYgJi+2Vx
Q7YR7HzXDqKMLMoEeoTc7/D0vQepr8afcZAYimVDpisu2n8BYiP51Z7ZquIZ
IofokCiOZ8G0b4+g5n9Gz52M83D0LaQcjJd2kh0wbeykI65tDelnA2OrrRcp
6LmLTwrRFn51MKII2iSfRhQ5j3x20YOUnmAiNO0rSG9UxNyORdc1MNkIy9aM
Zdfx7H5UrwDrC1oRMsnsihtMt62kZojDIGR0Zm1MY88bcXNHAVHUK58hfwc8
0LWQTxm9XkJ5+0CFA6FrSFyTNRWWcCI8OL5hitazSa9ceai2OsyHUbPJGDqr
DEnx6a5L2+KiEcvy8P2tIuynzNeOu0F3GORyRG8BYxjBk+ikdnKvff9wFCcx
k1KSMJauumiHx3MeSSqgKAsScMVpILZt8lHWt6tFanDWj5qhfHxjnxndSsVg
bwLWpCTFz2XlSh0OiNcWHK26ornRprRPF+SJm8W/vNUM5Acw5enMjm/n4Dk8
aetjk7YbA1dh5LMpJW2P9gBvH2dkAc6MOY2jpFQPbmn+0oGc2dwM2/5GW06M
y/iIQbN2HSQ5Bv+RAZ7Wi3ixCxgEWeBQ31cay8ozmZauu0f+alfa8LlfMNHz
fpuWC9iIjk+6IXsdqyc9e26KSJgEB2XjHvfBfiIkTL243mPvQuGIY0GrsNQa
d2p9cRBvBz/b5/wFx9pkN4+4GkP+wryL26onrZWPA5XtpSePSzv+bcMklpMJ
8e/cRgw5bUw71Rhq27xRXiB0tWu/HNordDLWqp6A6W1tYfwJVJpFcAWa5D+p
zgFhMLSrFJIckE/Kc20uUo0VOjR1/phexpqHXBAYGPGGxbcB/XKv/HudBBIP
sz+lyRM3zhRfcfOdgTRz1coJFlnXWvXTJ1aMClMWSMNCir1NOXcler8jcwuY
o2Sqy7apK7HFN1CYYMerJwMb5FOIDsEETBUna5uCqDzinVJMo8lR1/UheNI5
4wI3Mra62SDmsmeeg+bZSkR2nZy9Edte9pCvSrJ/KLAYUmxP4JHl3/8itRV4
lpQao+4/P6ce8MlL3zEn34+h9WcCLQe0mvhbJZJEdOuDNlxMr8fmWhyLE2rU
p4lx2tZDA4oqOLDC73k+lKD1tWsXCavawjtqOm3tDRQ8AEOfQhxTKLq5a/+3
n3DRcfIz7toiulLn2vKeqlDg3VlkX21DSiYvLxGkPOvIXizAsxdZU6B3gRwI
IwiX95IyDZxZSRHnhJAgsVxjraz6biK0eIIrvnPz8nRCc4T7c3L/7PB5HCgs
GiZ4aOT07Q2hsdcYNczJaoDvUuE6JRn8GTpaIb0l8cTe2uxufPZYvOL32ARY
n4JBp54p7QEKL6846Sc5klsGD8R0gcmPMsoN6ECwqz5NTLSf4Opb4S+QQCLy
vUrEEw4X3AJ+hF5NUK5prw9y8vMTwOFFgAwphfc/+9LU0LoCvqr64bwPLOgO
8NtsnWcDnkDRZvfjUgySAmDgjWPjWgWqkxUGbN1QK/eaAuNI+NG1kYMdQEmb
mHjSBmSAAhkE3WpCWEYcInp/AGZQ0S5O6g9JuBiSCe962wq0QSmpKMoZUSDB
qbnpAawus1/Tf7x9E11DpYIA2U3pV4setBCJnwjzSuLZdtTy+9JbE3Oq2c5r
UPFsamdA2q06jTLnaVebUo/2vLFz86w3EOejNaRe1MTJyBL2AQ4EjJz/+eYr
ZyoSC8kKU2NSK/kY1RpY3oilpWWgJW0vV91oMUk8FEp18BIhusTHwfgAqO9S
EUuoQGmjIpUoKv5auWAxIHFtuHk8bzSpRvrAgJ6XBJIMEwSCs8PWmUYe9bQ5
BRv9Kg11l/BiWOZjRrj9EqA/9ta2L++b7Gx+MQpclMjRVMF2BpfPJ3d9ZYIW
CwzgchZfqI/aB/pOfWDXv0zMj1usnn3MsIFOIv5bFnEuKIyGnFgrOWlzk3YZ
dT8WCapxl1sNNSu5QTxsD1oATUR8DggjsW+Mszwrrs9W4ucn3CIgsma3vKkx
Jfp2IJ5XAyXEJlEdVHC4CmSLVihx5d9pOigENDa/bkNyDLsJ4NDJ9j5gX4HA
Hoewvlojidgx+vnK1Ljs5aEH4+m3v1VWpUvhnDhHSExxa9UAjwtPLJmq8uj5
MLqQ++vNYRPlkZeFIVSnmlyM9ekfGk1gUyt3ydpv+3ABYdSCZnwaBCjCLnyH
thUUFqA5QJpaPCkb8e5TKdyeYS7YyI7Ybq1gIuFbECerohvftRpENVlxla9C
lJBnEPxuACxnP4QRtf6jQ4kGEsYdAoLi5tOfG0VdQwUoYClrEXykOgAmYH8g
9cvwXw6Y2AWZc3/C+lzHPNBFuX0D0We+CvOHA1dsGr3r1gr0K8naRl3LmA/3
Hn9wbyy/R8mH2Tz8wzDZXRuokTbARY2i5Hgtk1jTZIg+i7fllVmwFJjeyLzQ
W1ClmVlI4F0IbGz4CTyfO1FLHktJo3POy7AMhLPvMe+9CsVT7WLMKq21oZwN
wVsuOoY3P4OeyfvMyYRqJxmEIOzRfbYzBDzUSWaRvQbSRosi8SOtio4h2Bht
TcbzQqG93PHHHuFtx8cyoWwsuk4tqG+TR6rvaK8M+0J0tbiQuvyeZ074pbyG
ckwv99gesn0avvAUwBetwgOs9OfTijOo+wuMoz4sYzdPzbK4AaphE7651gc6
7hPiHwk18SttfslrYiHCBbzJzwIwJBbEzqxN80NsZkbaNxZ5TzT87ehkQehT
75HO1EOgioS0UcFUO3nfvwK8quYTqXisOpNaTiCoYeVv9QceNS2D7Ubkt4nc
3aWjPV/B4K2uvrthPmMaRpXBrttKtUQjJMfo3iGXActqtURrFvXvfbRlI2jk
79fMIbVD2FDKDuwSf9nqWAHbgkESEJa7IHD+qaihYOvmQwlt6WOa50BtuJrs
EjcROiS+9wRfeJuJUU5G9GnpnjXYLe75TsKF5RRZOdWz3bJ5h2ELsX7bPyqq
vTP3QSiOEggRySp5r0H9HqReGIfgfFHppnipXMj/AhDXUOQeuyGiYejwyWQA
QNNVMg+Q0YxeIGcqE0b9p4dEzJuDNO8y7e1QlJoOC+QduyLG8xhIEtejRja5
hmHPyFZlHwaPUcuhkaM34q5XAVdRLPmzBvmiAEa41EcLp79H7jCGFdBUGdfW
oo090MV9HrQZXP5gYboS+qUd9hml735/r5PdfZZzLB7lQLvpm7UL/bxMVGLm
1h+BxJwaNTEjF2etlsFIGKF4wfDg2cx7DZorOjdAtnnzd/dCxx3bioMv3QNu
TqcMBzCwHUSC55As0aDIrVUuDw+CH+/mWsXpR4Kjq+ptiTgrusnAk5UaDbb4
r6175BvssBblxK+rMir4RgAIP5o2dnP/GR5BW8caLwPYZ775TrcFdetPnzhl
OYSpXd+/QDX8mIkCvhRXMXxm1m6ZxCnjb2LK61IntwfEVycDYSkeNOIvWxei
yWyk1EtfYHp+JeHp3ClyXwQJ0ghq+UOaLsbOVJvvKBgmqLf8YYdGzKOVe8sl
1+Yoj2rjUohnOWmZoGJ2FYdLHb4FfV359oqV5QpsGdJRffPkRIbWo9K6CZ89
ekF1454QJh4lvMjb7qMv+qIjG7jR3Cke3Y43wUrTsaccrsPv3vzT5TpA5QAU
BQOfNq5iO1B24/9GqRIbZ3T1Bi1cuvLRTez/uV2VRqS5TXu7cber3OO6VKUO
b2QRjj1Ag11QDezDU2OkXSk2nMsfWaYSSn9K+1Z7rfAbBz7atNWu+VdWlIfZ
ubQbTemc49pLNNd69DTiDKJgsb2abNOEPTN3oyVAu1NsaDV56reX8QztWO+z
VMeVYnVO7QV5Z5KVLpfXERU7UElYDeWt0RcYkhU5/5q22I4jWmtT7vbYEXKE
E3EmpNfRhOYFL90NVayJfbjJW8NQEYhfhzJuANIFTAAI8HZOMd2ISVOOFp4n
gAFnfDnVuu1PbjUJXp/NJqg3iTmZFnRUEyQDUpjbKhzSnDatX5FxTrUnPiP/
KoejuTASkfx3sq5e0cu2lgYejjlVHakUlIg8smjn86pUEZP35iJuYurt8ds9
IOAO4Bz/3KdRFUo9khfiajhzBSPvHAmy8aR1FQ5e6zEDDrM4ygIBsGisorpL
SIY9jAXUOVSyfSwNJ5Wh6wLNdpzZGxL7nzYeMHyipd8Pr1UQKJ85k0fOwCr9
tbkOY9mWyVhXFeH3mgFVctXC+y4A3nWBWEQUHl3zI54nIolADUMlU2NsuvRE
xG33qSLrAtzwFeMMMAfwK8uJV2HEZTju+jqThVJa4HiKhF4YCIIFi6q4sKPn
PTiebI8rLWI7ktYrfFJ0xJiQP7WypnIEg0zXfZhvnhY4vL4ijgfd/yniZLIf
nU4iXQpHmMaTXSQY8BF1hB9NMkvySD8l8b8NvpUHM3zILhlHaO0I4MQz4ivF
kJMgVR0+h/2kkQznDh/vubHeYijJB/z0yTiify6vj5mxEcQP1QAJaeEgyTgy
meL0Wc6zDBoH82Yk8lch2bbQSeKdgGHCMz4JSu1Ds9+vGEEEK19yD9A1qvw6
ZrJ5XT7IyibBLADHp+keX9YxQ0ExKn8dtNRY/0e5/L3+J9Lw1RzsJWNxK+rf
3+mph3ij/BNeG2YkaYpHbnGrAs4+vSHlt1+iScZX1oQ8qVvVstXC9WfbZDUP
h9ml5D2u0LsRUleG6u0ksRuwl89DybYViDEiFXzv+rS653xODwGlE53SO7vp
EBNUaS/OAc/d8UT5L6r5Rr4IZ/PC+adctUMZsIEI0Qrc1DXDtOgwPMyBEhOV
xhnsYsm0Q6C1tSpgYXEkN27T7vwpoqA1UaQ63USZvuuIR+lEjeCSu2vqslet
rSGVw+zIKzWYLBQ7xuA4XElBmm2y17bWRxQw2+HWsxaTMBI9TgVGzTeOGnun
lx6gJrOWlfMedVKdV8dWohb9by33/+1wPdu31DlZoiQedvqrNbnMzYWyoeJd
fcvByPRcZjphNGcfEbARtQO1Uc1JY+c2Ym/yxlPGrdfPK1zLUbgo0prLYcKr
5xXtzqI8KkowuUpcS/S3oZJDvYuRNKsJKWnhvfUwJr1Q9IErqE2xxAeBalg2
fJxuuG9Sf8Bn6GyvCtjJxYHgwt5j5CoZcvZLU2D4fkpy9GWyJ8TSvsOopuf+
JHQ+bdS6jRE3CaiAK2AVPGsUq8NsHcfcZf4ocA1WCc2J5FOzVwoFklYIzJ/I
+cR8L7Y0hjuJlZGrqFwSFyEd4OICbS2gpdG+tyNhyIUH0XoqfJOf60vnSggO
cZojHNk9+bdYI6pmShY1GMsAeO65mg/LD8uAGS7GrLNLuIxxdq8W5gAaZaR9
FKkQLOeXDHWrFi1sIJywr/qYUFQ0htByX0QtnVofQh5J64RlpAa/0PW/iQDP
Qe0SjWkhUQiaaAfCMCXVZDgLacp5H7dUv9oP9KwalkFK+CgIjrx3/Nkv6yjD
ElBpvAEfOZnY59ZRi1r3EN3phyqY/qHn0tNqmwcVWs8JKFRwn985BZLD6Jhw
uQ+ddF8mv0LaOWkelLE2B5vcHa4D7gfQyN3U8oLDHQzB4JYPS+l5tYonRr12
BNltX1UFTMJlACM0V5MgwyvWQ1AaoEy42vKsEWVOTe9jK1OcS8QAqV6jpSep
ztVwJFCqx24qMAyUMSjZj668nBwbqEa+r8Wmz2pZ3Sx96vd/beOTxREbNAc7
d/dJgAbbpqxb2e0S1cg+gYdURnoL4ASxv3GsenJIWjZGcfPAzycD++7Gh0zc
jDtPZq/RkHY07QLTXIuwGp23NJv6mg4A+RCuan36v9dKBhDS5QxUJHE3Z/aC
XA0a3edMPbDFOJ+D3r1oMmmqA3UMYjrmq/jMWsAZgAgT7SvW4bWnmVb9ulb2
KQtIsaIIBOcpQDH4eaUaxGpgfCIUV+ye3gEZ5ApR8+PiR3z7Sm/Zu2PTXtoI
yb7YB8XvPRi8oP8Cldau4Gys+myUMujt1kk+ZWf6KfGTvMB6U35HMFXjnlIm
hkMwo+lhNXl4SwPn5f91LpSMigVqw5mmdeR6fNsHwoQ0GQ/gU42K1draIro9
fDVvv8guN1zUs7/mD597UcvKDf7SgFirsxDM6FvbmTMQnGg9AnSvqFWKDwls
tGxl+YMgP/4XDHrO9aZkH5E/CJGwmfoEegGuxkE44hHUJhjh7zaVoMHbrBDz
c3byxvk1NY3cZZDvqMxM5Yy1NFQwgPS7eW0fj7wJBY3qvn7uawbTRPzXz4Dp
qt1GaaNXsDdz/UXYwaWHXX5t6s6g9oZ0NC4sBvC4qneGrgzgSWDCkG6t851C
pAS2nWPTpqMuUvxCqYH8hhKQglyyn08fGoi4vzPQQboj1m5l618NDSLp6ryi
hCvwB93rdkcqrfSMZKKpWDazszkODKuOIMF8bwmmrby0bAQoEa1/J2tkq6mE
o6Il+Jk2Ocm6jOzGe3WrQ5eZFR6Mtp9Hd15lICWH7GpKDZXvhgqNtfJ9QWX+
4zXEwSJVIBQraaZ//DXcnFE9wcHUE2EkT62wos6/02QqcTEnAZVSWQe67nwy
+Xq66c6ivF6qn4ZXseNuZ/MdlZNdDh1ji2CXqEITG1KROhg3V2baq6eLNUij
uYrfFU49Nxpb4L0hrzsmFIfSuB4StfGFisDa9y1Cf43k4GCA9oRT0IjvomZv
nH75k1dqhh0qrHDCHq0NxRKPX8dN9T5xvDb2W9/ZseIlYNO7Q6Hj7Y0Lb0ec
gy0FRjK4Zs93NooV5cIiHLic2ccQixOV/CBAEg0pJ+W7rUZO7JeKC4fK7OEf
zt/06DVRe7Aiuvy2zvo1bnX3++7E0cubLBfZEtjTViAPGqZFGIC3svfggGHD
UMFcEhBxItFqYyvSCmHzXP2AotDCSbTqRgbMOTxG5w7wEceXk2QklkhN9aeT
Gg/zDPnfuclJeOc0UEqt432+vEg3cnU91mxR/i+ZjVeLfRBn4z/x8KGzBJZV
KF5+857BE6skFBYF1STHu4eqzOCBGEi5bciFV974iogzfYqIOHBYuRgZYQKV
BbG6JDdU/oMCaXmVZaHx80iUBlNhfxy7tMXGqD7kywjyqRyMxIeRuoTRQhdR
l8NeEm2P5BY3vSNi2TZadT03RM7MDHi2XSFJLOzJB38WkuWEQXS+/V04CJ7r
Z4mr5Gtj/14tq0nd4gsUNBOZ3/A5KMgR9+g0NSKKm7gZsmP+MzfQPC70oiN/
TUE8krEh49DsRC/uG6tE5/dzIV9KpxkpPUun6LVRLIlR0CBFQlKB6gk8RZeY
B3Yj2s3WGzuaf1Sf/jBVn7d/GEENKOiZmfoTCceDSZsNV9m6by+K87v5LJCu
3fZF5/EiIbk1wMBDTrX0AB0ilO0/zmGiocYFfwSgZ3a3pL92dXGjjjNYyTGw
+EQ3l4tL8Q0yoee52MSHp27gL6WcnDbGZPkzM2DYYm02yj/5Rz+KoOShtTsQ
NA7cpqZLPVPIXz43k07YQ6oA2sR/Ax4CoKJJ2PHLuFb05QKNoRiWRjljXRWm
5I3ZJJVeC3HPiruZo6Q8d8tOhq9xGoueu1AszuQbAkUXjRpc+6FYR/dpHaJK
OUlgihiDFj9Re2yMdvhZQqvIt9AmOsJtQcm79cPBpxNOe4d3T3NkaXyPleqO
MxCDoEOA+z3UhzQfyjO7yKxWXbuVuwHN4HNzFfgcB+ddJd3gjCKG/2f7+swK
0SiHotIy0nTyqTJFxaSyREYWN2jFd69OJ1OPr/pvTUuEHnp/+ClMaIcqIWrh
LVoTAQG1G6hyqeynkIzF2G9VHnN6/jTL3KilqSe1+D5VjN2MgJt0LPhW8+Nm
sL1MJPx2EDFaToIlU2/aDk7pH+GCXBTH73YRPkSI7Yq88sn8VBrrqhXCr8nD
yDlxzmxPOun/b/cp+QjRRWaRKppvbY7Bsm6o1ho9lPLCnQdHUemVl/XbEoGH
T7E/8V4VjdMlOO2pf+AOMyVY1HV3sLMovsTxTTuA3YUrg2qJKK+RagZcLpVb
TeN9nFdVuFQCEK3Ts9uv6cWHaBXs6rx8An3Q4cawZr4WDQ5GByfDEcLX2qb5
54ZAeu65TiJgS0UUlK/JRtU/+MAWYAkC6F0/ym1a0+n3qsHi82Tk0OJiBhu3
/H6N4DCkwJKhbqvONHoMTjm43cwGiuA6ITCRLw8dXFusuj0R0cgEXaeSOzto
XP3mITF9s8P+a8lzlnAzrLqlewPVIfez5NJJo/+NnTb2i98SqoJI1QNkJB7v
3Nw7GluWoIrnIgL2WfG/NDasgKRngksO9m4kVkQAPt5pGkPsgJaLJbju3Y7S
LptFfbET5Ud9bLC/ERoduyr1e7KPHRP9qVJckHLu5XHUB3J6PTN2NqM3IsxO
wsZPOquJgjxsHEuu/eT1oBWchBw7mZytSkMuC0B0ZIW4CymjSAHK+KYupL2S
w9lWIPLzFUIUPH0Ucmozb/IFO6aN/7eZNwWWr1uHIVHi8txSGx2bazZSMn9a
SNXZNmcPSjzcCJ2/IH26yZ8qBWsEAASZFn1ocOS5Pons3TiZjgD6Z2XOtEIU
E/efOL1pzI8eWTx2CR0Z0pSnh5B96r+sbM0JKnuCuplFfj3whuHVqW12g1g1
Xr+FQlq5cgSygAYzz2i5Oc1DPeSXwSoJjTn8veBC2aT9gVHf/YU1LEic2548
q3ft/1oOmVIdFhxoeNPTEgdSAbqQGzvya338dE7xCcPGzZP6q1QRleQT720q
rLNOhVyUNX2RqqczOyZgURuhSogJHv07lkJJOn8EIRzkG72RaT7NimWBPgTn
ExJWAA8m1PMR80ZjMIqyrAcSaEgBQHGLRz0iWlCPaYP/BC5MLlK9bihBLK4x
e47G/1LbIrD/5G/ealzd6GA+7S31uCPwfBCU3qEhheApmq2ewPcTwq87lMWc
6ypBGzWYt0KT7bYR4U57aOqmRkQ46LKs2iZfmIv+DD8IWKTE+8V+gxFrCTZ+
qKsAEZ9AlBsbgrpg7YOdfedkOnlnGZQ/kyAmRt4GTf0a7hnaEPhzVr15QuCx
IU1MLkMX1YkWtqtV9mRVWhtR+5pZ8kLulqRwvaajpuasSzfUfrTwabBr1+kt
rEUjwTN9+1BjMZwxn/iG5OS9NN9LhjfC3CO8FQmCPaoK27yLCbeETy3e1bJV
NvK4YD/IiuC7AXl+8cruztTXjDCAXibQ/hJ3FX5IS4hekPE5amsE/AsqZ/AT
4igRzaBO5ukMewOHFOg75DV/DZX3xQzxEh0YuX4SkmXoe/NTefVJJCQB4sB6
/t8A9uKCaH0QtP1P5zeUHXky30of5Ufbwo5+W5zpo7n6QgXltqghxd1kQ5MC
UPS6b/vwyknQV3Zjxy55rxJ8Ec4RHJjHvwLVVVwQ8u8dGslUnHF9+ZY4C5O5
3iJeZ7tAFv4oD/YjuFxz03kAevrhZLbGUc9BnaeNjIwg3dfuBI40g+3ksoJy
hMniZBkrtvB0MB2LuXW+vehNKEVw4b7SN4rzCThLoqr1WIkHmtZ2E5WQU70r
cvZqd4dzThSeiOXhW/KZkP2wb5jGR6EstTsXsaVyoWj+9lbg9WwqrtrBUzvc
y+GZO7lU05v4fqVbB9qN92Iz23ylPw62cd5d+P2K7kG4ZpUkMkofl3YUfaeH
NWdmYsJBhHqJYkGoomRfW/P38PZj/LeDqTIQZhRmF8c00JJj2ZbZpHcPH50S
YAKbQBOUgitZYnp7/Ah+nlgPmfKbRSs5Wrs6S63bIIEICbfMNQgUhim+sE26
2Wos0lNG/7Qv9JqaZs/0LTJjzcHCtukT9qYeSTvjSK+pcB8I0A85tX29Paje
CEhlLIeIgVIJ4RiRMJLMwblmvGdm6qL1kz5cRdAQT/nm12X5IwtYL7CqrvKI
oWtX5zIrjxE7VTYY9fmWC1F3nDmZ+UG9uNZq/jalt5u+6H8pJa8Y93hKEkMn
RMg1g/hH/K9jkY5iZ+vi/B38TNjaFyUUMYI7jeYC0LxbbTmNksfNC2bME3xV
3L89lw2RiLD12Zz2r1mD/rL5YJeNKvmGML2HrQ5yaX2abx6ovP79a0EmYSLy
DjGGSnY07VC8cBgDblYoWmrCxEBN5ZfDmNImedMkw04topCJWloIWMInbG86
nTI88cUI6Er94cT+e/G+BiL2G7O4J5kpw8f3Or1eFg9LT/F5/r+X/3141FML
feuhLDmKYEIhsVZXd67pyCpEe2ad10bDPzCLz50CjD/usJmKMJylwYieevs2
0YzD3bT7iVUUpz3fmxR6U5LjrQq9bLLIaQcgkoHJZlPZ88NvWEpwxeimuVKh
8HXuPjsKXdcZWjDrLHOgwK8cqkUSXnUuqqrcVmwS4cV1Tcz2UmXBKZ2GhuFv
uFUIENY0+WrAnMsqmYf8VTV91iq73ZQGU0ocUuNioM1kZLq4vzvAcwOcUA2W
r13PU3n3TncHFFIoilnd0LtCAkyVyhUXf6/r0oz9hOHtHOsxJDtH/BstTuBk
qlxnKabtfp9OIWzZBre4dT0B6kSt/OnVSqcJv1OhQsVaCroyORSVbp9Mj9y+
oZLutqPNCwt2gqI749mxM+fBslR3CQTFSp/LAYYmBJ/FqmyoGU/VN+Yjqx9I
yfhWnM63oPXOuje7XoZ9QflOV47hDp8kI/A8YsmZgiFmib9P5ZsRBRSHsEuQ
uBXQKxDBQO6jIlcqvgewXH+fRI1XMD/enf2NBYOTaxDiTApGHusXNBel94iO
LynXs/Yxxlg4t6SHghHeJUzkbxn24M0XFMV0dRaORlNsJQKo7ReQs9rm36N7
04eaMqURXEfBa+pr3+T4UQsF73TIPCQnU9QOfWUl/s0V0EYsQLBPj9KqQ/Jr
6MieMNdkMANuFMyzzPTuv7gB9um9IJSIzwIKbbntMoUSMVGe240TTeq1YRF6
7T1L2I9H2pEuzcBqUW7aUoCICDOdd/gT0U434POhty0ELpCiOLcZWCpYpJK/
+gA7voZhjTMWhOhy2XGT0FqvWSJG+RVKjX7mFNesphgqNo9B+hCLX3HzBLV7
6P0hlAu/jz9dT+Sjmh1mqJylLKre6SKRFldFI8YicSC8gv3I2bO1C4WkCGyJ
UZ8S9IgwyaU+1pbevY3g7df8olcOjZo3fYqkB0owqlqmfo7jxzxevCTV1grE
Ug5LzdmwO+sIA6U0Af+EGnc1AvuWb+olX66JkUHgUQstcrP4GrVzbgWqa0Pi
ccqP/1BsH4HRs6tzEr2rj3owG2FAHhFoZvmA7YeB1yCy9j7ee22LlW4AUbV5
vd/LuTVU5WvEW70EZajFCPSqGaDsgx2CZN0KiA+US5S/oGLwDG8olctmabu6
vzUW+AWFXXFZt+TjW7HhOMA7h6SnvL3CydCr037Uz7YFQQ6yRMykv624V5vn
GXEphJ9C3gvDGT4+MDraoiP6iYRphPkHfX+b1h4ZVaBsBR6+FsQQ+GdGyKmA
JnqUCsKpGBE88NJ9m4xbCcm6CO/fRBNEV8kStDBBP48M9P5VCNNeHuZTDHTP
l0zjRI1TiGmIY01qU9TEcS49tRP+RzP2ZI30aL83OqSqp9CniVkPt0zAwBcp
68dRT+uPFXzUwfo8Y2UDaAPuSknk/veioCvlxLV+MO3nFeBpSvcu6SyYqkL3
iu/WgZSrWudELZasf0ODHb3Zaed+YhMKzAgTM1sREq9kqPye/aRdQBb5RTwD
OxbJqITxzdLn0s55kJ1qlNeSmelSlYwnJzvdFNG4c5jJyG5WPvH3bHoMZv2V
qB4bPWcBueuU7+aSQ+guwjAA2rQnpq9sFVURGHxwGI6cVisxqDN6gmtfZVdI
vco7udtH5xPEbE0034lgAR543zFCrJBeqq7ijL2PEKrbtGRIlefU8nxRJR4o
zmyB50UAPE4Ixe1Hj2GNiUjQr8kd+Ltt9SQdvkPL/Kt67dK6O4iyquIshrmp
tSq4QO959NsM4P/9JbheKnPTuJ65DWLkmkoLj4uLY7PTP8AXksa6JeJLkbGC
+s6WRH9Jd/03Qu8X9WfZHk5IwehEnvcJnoJR/+5nP2UtAYGTbOMsAejFZ7tM
bciJCyjNKksqpY4NVw84O7KsdTCRIpuIBu7KaDWfxeWlvZejTlV5A+N1feLd
OF/GlyTI78xZETRm7D4KnRaL+QLMjkxUwy27J5p3xEL30GgCFhdjhPmsmKrf
voEMRDCSPbXd6M9ObDxQ8coTZymxB7pHOd6Ds5pOhV3AmYgzXBTlGwOyB+wq
VL5Xl1rzvIwZjlfDyWO0SOL9eVEDv8wEUlPYNV8LIWxfmj5yRgU4PBJK13bl
/bp/OTBEvwku3OZCSrOJ5BBp8F2hatSCZ5wSumr24oL61fO6nZ9UzhpONT3J
aEBK+N6tDiQv7c9gzkG+EQZeDIRYlVgqyee6kZdK8mzT1mR0KEAx1tzVE/WW
sJCIB3K4qNZhhLThXebhJNcUhZn+Gj+fw6wYIS4bDjB+TBCrkFwmMK2J8Emo
IHeUgVPxIb80vWavG4iTLBhQcYz4TOofDcu3ipSxd9cnpkHBW8fq5dI6pprX
wWVn4tHX+L7MmQWrpdt63S6IRLAGk41G3wdRN0TrGVtpLUgY24FGGXGWt7VW
v/FZU0jisS8QQeVW+625nrRWxLJX4jcb+fv4RE5Gk4+t/Eh9MSQl2Qi4uYsw
TxLMlu1NBUKY3yibLpwGKI1xop3TKuZzJitbOUlnHzh7KMXoJjCd+TYCc7O7
rXWisHtDDpPoqhaiDhGaG96y5SVsKHd8J8SMwj6YIJTKeYhQmrIPcob57UNA
8CUXDe2lR9+8lmyfta+P3/PVOcqNlRewQ8ZBFn+YjNl6vfizxOXteS0omZCt
+e3jV0piFhfNzjSs1u57Dr32Ijt/4N0JwjJSTqLrUmkPQ1ygvCa5/d6TEzi7
2PageCAFSbaVGK5/RAIci11+6vEY2hKlNbS6Z4mXxYnyeXd7xqR3z6ObEZGf
CPluwIuWwYYtQenZafDGIfi2TL+zzcwojyMXElYn/c3x2glubju0X8FzoIiC
P+joYVa4SdmzoGLVUdoYWeeb+GZt+bWCAXrD+Zw8I8lHPis0NOacvjvPn1hc
wv+1gW+Pvyqc8B9/6q0BioGKBtVoyuNNPcvTBngs742vmltGJTW0j/ebtHr2
cQk/djI+HybpF2Ka7EPqg2lYXS/glFzIBqErwJGHvflyMBYYjfTE1fU5JluS
7kSGP8IqNt56iDWLkcm4MxI1JSBINC3np2GhnuHG2XK4/VRvRGi5Zv+yo5BP
zrGKNFzONwQwOsFB8obEG7nUEmgZHCJeACTK7eW+R8p1aMhGAFNhiLduPfxe
5jzBjiz38c3ketxDI3iEpwwYRtTxd2Z5x2JMN0FJqoIaAGketS9Ybkh3aRhe
feH65mWFVwBd+CwJjL2dBzucW01iZTRbvQZQcaC0l3BVn5gSaP8Lnd2UwGhI
1iU9Z4MWDXvHs9s5oLyX/vMJEf+HU/tlDj7g+p12NRkVM41NrNC5B6OssUW7
5uCLW4KkNQCCbR1dXqxn2sNzhZfUAOOmOz2xOZz9e7OMYLqN1EySun/zCzMd
TXp6E9fToYrTEgeiyWHOYP+uoU+6DWX2vh2JZfLCT4XP58t9QKsPJIPwjEg7
Ll9Y0kbi3xQqkD5h8ZacUkZewbFdgW0jvMl/6JxcDJsSIFBVbl6xHSp4TIoS
dKwxmNelK6jAQ25wXsK58Dd+jhaMsiZ4hnU7W+fo+pTQ+K5sFEz7g7GChZVA
RJ9XoRlErdehekI8TRpnfEAreUUurTUemYZMEpQVXOYxQnGj1xyVzqDikK9N
2LIKnOLByG6IbkZp2e0mMJxmoce1lP/SZmn/LQ0t9ONbk5U4Q3vYT8zQtaA3
tIhVT+rj4KrcwM5ajkiTdwRyeL+eZl3IBwUKLQ4i7PcGpgQ4sUBM2FLsjO0C
HgAfqDqk3iBOvyB3ovz2HBW0Q9hIMqreC62lZOD88ztkcwsJ1hbK7+zLmnZm
dAuemdiYu7OLe/WPLTAP/TEEiQ+FhtXy32UwOKLRhqZGo7/JoiECViuqt2Pk
wY4CaAjoLeeacmNxNF/t+QBPb/NjBt21/GE+JJuqzGscxfIW3O1JfjKJYVl9
L7NUa1jXMLuSDOHxM0USnEIe3G+Er1TT8HdUQ/aU0Rw2eXbiYg396TYusxM/
0dn7nVUS+tHsrVOot980tX8eHPKmxQPhmqy5vLq4PM9Xn7QF0aEX2bwJ8Hxr
m6DTuX2wBSMH54BFOYnRG1tvTLxRXBevWbP6Q/BLqe5qj9gyGwh7ClaR86r7
nGOXLDR3qkhfTq2nKOwSPwEoMfVqH/HLIqd+tKIy21ojyTBy/4+C8hjsbF0y
05QdE6UsFuHgL/7Gp3doggAgf6KjLYqlyxO7IyB0uyfEIHv1Yo0YFwH4oxAE
sJM9zNb67+cAmO9RLh9Rpv4GafvhZj9v4tKyUJjTG60XtycEdur5VSu54fx5
16n1gwqfLaA1liKHsDn7uIeAfHup8oO1adiLb5uhww0LUARNKrVE43imkwQP
WGdEKHJ22D/EVaJlKKh+TF3FNjFL3Iq2qUxGdQ4N/4M1sweiu809PuSg3MX0
bXP4vpPYHhYYwMYJZVmbZnc+CjSd99tgW+l+l3I+VDJ7DCl1gBigT+op0V/6
WHUwgO0wwsMRYRrKtQHFeIocqcg5fLi6JOyoe/YRLnvLLmEhUcvoZsAFGhu8
iqhSgLmxPy0lkc1jMndFkAAFNO/0yHH/egfsC02GlfDcoJL5L8GTpD5i9c3u
OmOgeBMdlGKB0YvBa6A2TxiAfVNufoy/waLm1Yo9SZeZYaiXX62QlbJMzFFE
W7tb3N+SD4/nFn67DZzLPQFn6cCX9Zm4K1lfb91Oz9A9kMr/w0/OqlY3bE7R
IYw1++AYzKe7ytLmGAgE+br1bjwwa8W77a7tDABNhnhfCW31G1AbWskgdFtk
FieQ8h5di7c4pjJ+NSiCpk1bTA9gvbffvGohIMLJ+nUKh+nMNGZJMyeeEjNL
RwUnDTb8ETc9WIw2RT1xvzWPlTTqiaMWQpgMSo44FA2jDnRqKFzNYthSUaaD
5TLpW+y+T2Oybj+W8LihxDWr9IIvURhxb6rLMuV4yUL17CZ4BngPyRZ8tYug
5/zbspG3OIn6bkjsvSF9gwZfaK4fQ/gSQwjDb22cyZ0Nsm/qpDFuoZr9Boom
97Xo/VklkiYhoha6qDmVU2VhQIR2/dKQrvAThr+qct6EiEnda84nT6lw0iZk
IKIZ60YZ31ayAbzPRLOBu0bZzx9E/OoJCVoziPxfu6VpzhlE2X4WUvSvgnee
0CrOvAq9P7tEka5AFGQvi/bqga3jR2US+10OSAgMiGQz3fzcpjE2nMbQDmm8
lbEMHAUvXyrSZmMKqT4Jqgemybqf/60iJzcQ0y6uvohcsbULo7oEBF052CL1
J/9oexb+3NCtlKjJ5c/PdRDo/r0s7KqXyGTTJ/YCIHfciPuU3KK6PJG0urp4
/IYkTw5W5V0d6xD9HDqMXw+06gDyJ/EMKg4G0abZignWty8F+qVVGBsQTC2O
UXWPV19CWJ/G51HKY8grB1g7/XDNZRusJe6KnLI10TAFI7TAlOnqnad16vKI
DkGnSCHVr8wOgDI8xx7nvILtIOrU0zN5KLqawwVy+j1y36KPLDDDXaqx98CH
47hvNH6KHuaaU6k7EbEpVZmkHfyEXmItdeANSuiDl7i9ETpetT5wydJ7rjyK
JJDxTuCy0hfOY5SuOjlTJGRFNSCdqmiuWOsmgb43Vs018txe7LRA0wuKq1lu
82Gph2dcqh428RKIj41+/jPsAolnTsj9CuPczu8GK0HzJclOQL1zwZ3eO2Q+
zeSn91Roj6a5/KYqs3xT3PCJeDcjMZiYh2+MY4q75Pk7F+5E+k7z6ys/HwdO
8EjIhKp7WG9nEHjSSaNfPj1B8LcuHbH9y69zAA0qYi4ydrmT/Mn58FdOP1EN
dHIZfDWjy5Rw9xlRw+cluTe/TP6G/x7euVe2Co0RERzd8c3hvn0lbDuzKKJL
TjCpstMJQeld4cNze+jWFXrtfK0KfAqT7Vzi6izJ61DsLPsdnTKo31a+DtTA
ywaDzJ21ZIacFPkxl0oBSb7IukTbxIeeuB07cEZyCD01Jzx0Fal57BEmKg4R
f+Kao/lyzzcPavu04vEiZ3GB0c7iybJFK33F4HUT2g6YStbL+BDpbAOZGIdq
i2mEqHvv7Hf/nZ2W8HKvFK1nOlAJEpLgZEqvt+Nw/PFtC9VLI0Jskejlhp46
ZBXEBmjnGk7hE8LF+7Maocl4hVv2EIRmq/T/RL12vPOR0RF5J5m3sMgNrxj+
zXmdUiq+kJDAm1hP/AMekXVPqiDND9cRT/GDCwbAgKP6kJsvYD47u6u+cdvC
42BG+Cy3mT9gnNMZgVnc/RwYqHVxHotsgP7LB7U/xCIFNlq3q7c1CuG0NPfw
vu0VBN1FpViK3fDBqXDwQfgKfxT8fpJY0/5+6mQkWzktKzhn5tBO1LwS3MXZ
1trCUI49Jyuy56/1TEaNEvPa9nJJOYOq+JMjZrKz+vzFHBP7PPjRuYntytAw
k2CdPKbL6QRh/sXi+Ftan1NUnpDd4auW1QMJGc9y6Qmc2i+SfTGAyhH2Dg5F
QRlpP9KpIsgBsRCzJQeN0YU+H9wnpYsAa1bCUiyXlX1rZd3/IVAnwc77KxmN
cdCz8HzN4WkuBNaqOCUurjF9VPmj3yY+YRGczk4qRT2A8phzStDjIrILPIeN
TQZINURS4AURzRtA2trtPEEBefLeKpkJIlxYb3lsmkKKfSZAJHXn2seja1b+
zxwT1OO3AkA2g/3jksrM10dE3e+Ut0Fu2tkELTCuWplbcG4IKGP/G/oVUCE0
85AnC/7Ji2XwNQqmvqBxmrljXthONbWB5Pik3gP2DAuMZVGdkiCI+3AGfin1
mZqyEXrwHvV0YmohuXPise1QOZE5pdIkOi41m3Voa3POzMw53hTO/gy+MKYJ
syv7iKmFp7UOaSGVVtCB14V1V++dD3N3S/cnxWGSL9FELiAGTc2VlFBsCKoI
5nql3DNx5tI/ucSZf0F0cAGD/lIDjhpceBhcVgrVQk8Z08FpSarGISPRf58s
Az5qpILl7t98nOT5q0aOA0ErSGtchJ4LB9nVWHo410fkFqb8KP7LE8zK6Nq9
ok/PiYCKbGcZtoDY38hdEcf1BGGbbJxqFE6noESgv8VvmkVjq1eC4YhEEk2L
gz2NqjH9Vi4Fy3FqHnA3GGbFbnGB4vElzMk15WvxO/M3Y0vASopLtS2g/WaS
a/7Yv1vIKR1xRR9OrMoBk9nV8+YJELuSeT1ETU/XhVi47wtfHlY1BF/Q9a7g
5M5ZRVyKVG/H0gnWdbARugOcYRlF+d4LeBF7iaRYwoMHN+Q6HqxkDcrTCmzp
FZV+x1T+DrPww9PP9w25sK/O3G8VW4rofIIPo8BvL+Equ9DFScfjTJSBRUlu
xEjlSB70K6C9lbS4W9xLyvqu2zKjX8sgTGKrva3amDDF35a/L8Smahjocwee
EAhoq66pk7FGyRsSjGLrUN9CVdx7UULLWrJFTHNf2ywnHEvuM3eRRicIbx0Z
irgL+um29v6YGmTPu3si7xLdb1eZbMTRpMLD7zUUgc1EvdPT4s63sFCeBKoO
ZKnLj0spAExvFQQL5ACvuMStxAK91PcvBOGWzzo3c51YPAbWDKcXREmg2gPF
jiMOptXAzBlEUIkIQJYaWCoZgG33D5v2ci2y9ag4U/CtukhFbaoaTL03ibWr
PItIJbel3w3wJEeTk30rW7Ohi2jH/fhlx73yqEOQhN65SX7yhU2AcDOf5keS
41wkx4SQ/jSET09CEEwAEAo77UYh19UbZp/D9TxQUkZSHQqoxBzJxwdGDUGd
mSMXTgY8orSfrO2s+EI1rvh2w6h9FvJgsiFVxhB4UcS2d+VA/uVzxLTwpnds
SAu7CsUsHnGmWdBQL2OZAesjbewWHog+G/XfCaQypiA+6A9YGeRbsJULqWQh
Idgz5LS7gapaLZqupBeOos+mnRf2WbEVEY1Er0enOBSxuDiVwqP625Pwis45
fZqCWhQTJ7B9tu/9V2F3OrGfNNSPSvBvcBzt975bBl9QmcwZSqeuwDuWuvFp
qNCb8BhvXfib+IjADIGn081Hvbc6IMD7v8bFXXZNfLEeeG44j7/q1Utr3lrJ
aIvnWPurpkYwcTUsDqGGbxqhc6Oo0yZlZ9sA7HQGnXSEhvXNhdgppD32clkY
ni2kRsrq31sdKhZ2iS/epOxA+jf1EQVCHLzrCCCR2XsmLsySD7z2+lir4C7j
arZm7T0ETPc5HnqfdqYTsYPUQ8+8ITXqEBXSP6D6KNHKFkOjh1I7HHyceJLx
OhaszET0u/P17lossNG7kSCyycvpjbF24A7hHUDRo6SuvKk4DtXcFXOSlsqk
XaSDup6bPdzZMiJK7IX9Ksa+/v5U4jdLPCcd9JXsnlLpfyhelLJfYyfZcMpB
DMDoFuHtWq0dVtnrCCfMwvjaWTunUbRObrZiukdCxZNa17v9cmRsjsewQo7Y
EWhPUf/8YRTd1L1TIJ0BnreyOeTeWru2sR/BvjKAa8H43dXKRcwoZhdzxuIz
fa13/rb8T7D2/b3u8IdS7dXKxbEmxMa7e9NBZz5ws9NGiLSafUaD99HJHIZx
iZXjcQDb2wiTk/uVKzZDYW7t9XmApKHpNxn+sd8SV5/QMcsnX8evF7xoD0wC
oSq8gu1QBHPRZBFc2G79FxW2gFDscwYJRUzRh8HFG2MjsyKBW5k+PONwDZoH
+/FzvcmPUJ/IptOheWzcOeGa8iViFM2t9D6DuMBMpJ+cnU/U4R2QmFsAkKnY
/2z8cSgMCNNvHs0IJpfz1uRDLBekTM5L/TngwzRuraPs0zMYKKDuABivyktW
Vdfj/2PDoRdGD1ww+yvHykbKQf0EwmZhzodc5hk2EF1/5XM3iH7ngfLmlYkd
w5iZfZACcfqCNd2UlCNcJbuStFzEb4qI0lrKMGmltkxAqwHhhkt5x896ecYJ
tr5O7HXQfkgdIc6korKBAO6RIFQj8Bp/aJBCWSJ9ZWzIlWpJSppGzjHMB5Zs
TivRRmEp6I44s3DMVs4t4X2i2Eg49M7TbFLx4JNXM86Rvgtl444qhHmfbMMl
+KzjmccbyGqe3mf1UI6iaZFs/TQ+AgdK0A44GQpurJembu+/2lTR0Q+yoXWo
KkwFcl09Mxpnkxn4p7yrBPECHy0ZLlcB9HhzTtvM8QAZ1+fFwkPcAzLmSVU+
b6cC+g2puq50sETzvMejJgbnNQ+j28t1DGS6juY3zJ1qQ8/ODFG3lIHtWDlS
fWM6I/w0s3vu3v2myjimxJ6jYxjJEd87lqyluF06fEJqo7Mwx08m7uhssfq0
ZQzN2/gssikQ/oHxvCmADjVJk2swoDe0r+OaLbGPb7wcG4fyp6nv8tKdACws
vcF6Y8LIADoaqAFqqF7q9wpMnBtF77qEeuE+1h+E78VEpjoKU2p4M/efZ6DU
oBBMxUdwfdZFsLv+Dv0LWK9yR4mfVxx2wzKAmL3y+vEmkFgmNw0JV4EPyJlC
7uuUYbAp8z3Gk9B7feNwp7SMqcol3xOL3tedvW/swJ9M4asmqO/HDfVfPUor
7r0TQtD1j+4QFNyPyxxMzlNMeX0uJeiuy9uJAS3MnlY+ANJXLBqj2NA7y8dw
nfVkG+07NJ1AD9GKz9IwfBAdTjD780TKfA7VASW9yPub9h/+eg71bqKcyZmZ
XhLiu7jdyBzbB2eDPOFOXsBmqxP5aXElZ9oclM2ftqxKWJxuaakd6kROc35i
Ev144ySliWfmuf+ijzqL4tnc4rV3I7VJNcvvTr+QpMYS5M6patduf+pshR0u
042wOaL4Ty0i7FnIsxG27uOfMn3X1IbIzRkNU9uNlozoJ6VCnzDBkQI1wHP5
xylkYF8gqMCOngcNs8V5MQDH6dyclt27Xr7qcxXtA5fwNlFNCtEPwA1iQLB2
alf0VEoWfLHv64VDLGJMYXxidSwaeqNtB9Yhcpe72nE/CY1h5zREiOO4nbcR
NMOwG8ZVgCZsiK85HhUH6KcUjALBVC/RJc8vRbOIYfeaADUIc9Jp3TrehxB9
//HQfBf+wxIA+9PZLkbIjPmzB4Bp0r3ojdALIf8VL80uJtpic50U/SoIahUv
NpASCH0rSkxu+kp5yZ6ML7rfOP0oSVHjBULqaIpTy5POeI4uUWoEt6G+Vw1k
zrdjYxLJKhSQUuI0cWdMHqsuzftojwoYmvnXgsQvEw9j6NijCvxhYiuXVJ6l
gPeTSDmSsR6ZGO8Lk9dukK39Q3xhLXixHA//gZaZtxPc9OXk8gxtpqwa1YOw
vM9iOvorgYxrC/0bKBBz+TwPq7vnSqvtLrmm0sE21a64NXh46Xto6LSV0nPt
I+AWxr34jmzaqV9Zv3hyMQ2rtKbKNbHZsXmjDV2x/TSrO10vNTeOkuJUe0lW
5yeaCELQdjJ4lBc2G/TBZ4zo7VuhAhfWymNegJZ3Ew8LZ0fkyNh4roYZat+N
+TfB5A4PsJQUtqqrhy4DaZvQ9s2HTlk0j1Mrow6xgmIuy/Tj9nbIAvDLxYtg
H6mtVHNl49TA5CIf7uFdlqIj/hQxvpBVwidPhwxrYAaAKQXlF0T4AqMBNfaX
Bel7DB9YEd7oiZVJPZ+vCGVITAMC7huBlltaSroBp+qc+EBfl4e4SBP3R9wR
AF736/5fxH1K90kOH+e+upoc6LyIfsBN2XZx49t8BLhszfhX/3PiOefNtYr6
YKlEzTuaSMGdVbeCMS4gJIm3jR41Im+kxjXUyWK0QC/4cIRLEZhqb6ib/7ho
xK0JJ+aknhLxlx0k3oE41A6/h2YKuCT39XRx1ZD/qOPie29aIiu4D/uhsHvi
9ZGfZyZwZ0UHoq4eBCIV5DBrXbySTa98lIp6xxs1CB8PEDNSGDygZvz41IqW
Jb6evFYqhsMiyGEl8Gn417BKcDsj3qRdhXILtTyBp/Ih/Y3xK78Jg6GZpQYV
e+nRdQnFndsCFB6eaxXqozfHDfqm9HVw3HDkZvoaP5V/JWpTJWtaYOFQpXhq
hrc18MX4hTnvp4xTiQm3PgFaR0VBgOOczn8iXYQqOALBEywYd6AvIaK3z50I
Lk7Aovj75qG7ESNwIVPeHxjzlYREi9MntthLnrr2QDqnyLOdqIiX4jRzExYC
k2Oc64rgohc668aThvVy3Gs3PmyagPC1YPB02TkLqQJLvGt3vTmRWZrNj6j4
48nn+CjI0DbLs4VZPb59uGzWyS7/xh/4OjL7tp9mPPEHbvo+nxXRuX3GjxUw
auDs9ee7ZpjY1mhQWpF95ld6uUlPRcX3gdptts3vB/79udRvGncmBPA7Jf54
TOs+eF5LW5wMAaQkrea5LCZlaLCMEH7NQTpOn2cbknLBMOKQw2BIDtZbhlzc
HTikDwZZtABYUp0sEr38mknZ7DbwF1xZB9+sGfDwX78v3PbpCsbm62umK8pY
EUip18fprCVmssLSRqEd7svzkh57YpJ088AZrGIUtattlsWnkam+AM79cY5G
rOPFjfUlvD46zeCRy8HoSjSDa+b38eaRw3ZjCcT6XQoVT9aJI6TAtrezxczx
OmHdvGG5mAjuKKoDwpVcT8YsboSMJcfHL1s6QsgCCpRLyz+jCtQCI4NsiIHL
fFWKGA36VDfp1+//caA5DpJkuN4oFAHmTmqDU/hoJSH9fhWYIpyM45geeNlp
3XGiTQfm3GlkwYQ6wHQxoHgHlJ9RwiccLv8qL4ODM5bmYlvQZDRKTOiozfpF
664vFhgMNsewv8f3h5VMJXkzDkeakl6En3WVct+hdCpDOppXt5IamV83PV/g
Vdg4+bU+H2eu5lkAMimf0AzrwFfkcu455ZiUAVyrpO8gmqKJgEiY06SwvnQm
/V5gnpYJeYIIpdt3CjqT0PTpkZNDfsh2X66zg8RP9sFzd+q8l5ELlJwONkQi
f8Pyi1u5mWOw5VxTOc5nluiq7REF+aYVVdQhy5Jfdj1g94vgmtkfSXg1IiIX
XzAqIEbmCWKvIYZTRHoxZIV2wEOv9mT+bV7WYWEU48pNQOKZTcB0knvtLXdT
qp/q4mugjsxcdxLeVGOF/IhyRtpALHB/EmAtegqWS4Q9CuyhCrJrDNnGXU31
BnhxFjWPEVavmJsgLKyWBLy4ECPOSa76NCujRHHoHuKxcp5FtVclRSuQf5Sl
BN3D+cDxprkh5+GUXQtBJPdmDfNkuLsRYHyChJxUm/8j5cO3i1oMgBUYE2/o
CD7qikdP59pxVXo3cFGQRpDMQ1qtQUcxYOxmNYq5EuJSQWjQVZgps2Xk/Hsg
XLhZtiAmKpFzD2buRnjXfj4PhuF6yRaZXZrK/MQHs2hAJ8Oo5uuRFZa4WlXC
SmGD6htZmk3XyUOULroypegk9yh57jhqCClJyugjEZZtMGb67zOkflzVRUcP
x93lYnBvcF/3vs7jjdsEiqyISkLRoUbfnXA4Uszo4qEZkyfrkuLEJ1YIRYiS
FfC8uOdORr5ynYAwvsnhlhD2qf0za9jFVpz7PiOcaJfvtLu6NHHXvtBUiUBJ
NbyCRkmNBQNbwc44PVOf5MSkVkID1W8fQ7X/rJhKLp6MID8NbmOKEc5xMy/o
A/sRDm5rR6mvIVgBP5KMAoyAsB+SuabkmMydebVXQZWppBWs24U4YjoCSmaX
cW+acyq88MpxmqKUfmiVTqpBzZkBzJl2C6D8FPp5uR65quFTcFmGpv8AaT9H
w724LgxFIu3V7k0kYS7vRZ6njYev4MGnhTR2VCtZRigKOeAV+sXjfWLshDy7
G/M7xgyC7Rlegw4+XQBIfeh9iAdEoMepwmTLRPrwaYgPoeAEZdvazPBJtadl
J7VEnd+qbPftIRzRxxcDt/A6otdpBnjW4JebDTstAIL9ffWzCvO2C+bxAtxq
6hEdQJIWtCPhAOT+IE+pE20KP/ep12nGiUKjJ9qOZ/wAEsryoLMkDhjqs01b
c5IomLePnvh0xem/UDlBfQef6T6gkOO5oVhvx1EWYM3+QbP54G6Vn5hmy4ij
5uR2NeStaeWReHT/Xk1NK08nl9Wmc9nOxr1mWCUKLiaDucGEiHSihgTCNcfm
NDXBTLA8eOV6IsRyZNtiADxpZ4TJuEChkHl7dPHcMCALU56k7iGjGU/kjfR/
fu/htuxr4Y1jPoAF+UlR6WnlEoPh0BclrMxzahznHRk1UYBW6gTvY5poGgpA
Cds1pkM92Uzwjdsak/Wc+K8yL8C+I8wv0XwtyHmkgZWWH7zjizdmSzSGh/aj
YbVu3CvUDhkaQK+KeHdAkH9JtkFuHiu2G/aZuPFZIqaYx0euxv2uBRXjBuuy
wCvAI9WpA1Yo2Plw0IGhH7PLu9IbcvvN0vzYzTKh47OxSTs88JiAEUFmIUf9
9SMmR6UWqHvqgEwvBgUrMayvLXN4wSk3Sk0y/KKD7ii17my9lFCVy2u5mUrL
jpRX6sopf6bszc3zZQ/YC5OblxniNu6U3Nv+BzFlJJwAy5tQEEZJIs0L2GcF
lMtk4KQfCut4Qhx4LoueBzdRDJmNFRjPq3YF8TvbQs43QzxeKDJkpOWhNDmf
BRPNmsSIwFKHa5shyhSQaTMBWPrA7yweQeBnXxgDoDYLKVxrfb6X8S7BtI4b
zMiFtRGU9bB7H6OFW6g7nsZgDC2DM3yzk5HIbMbZwM/sWFKv06wabGdclLZy
00HK8TrQRgMmbQy2S0LIL9bqHl7J/W5cgff6kHX2ot7enjd1XJdl4J5d3wMX
/MRXq2biW3sKFYx6SkcwwYl1B8Gzi5B+ENZQ72GczWvs82x79XcSJ005Cvys
OOaY19TLWCQtvmfSNjYqe42HcSUvqSTF3WbI2y1VZ0rq6SeGRCHY9scL4fTY
6Tc/Jy2sbUXweDk9WHAR7sfI79QM46LoR64qLfBNdgaWWQDw9IiHe+2xac7L
DNrUBmSveDUVbZCesyjy1Uudvd/otYKzcyCxzM9jhRxgHZGZk5eJUB2oJ8/y
raSCfj1UE/r6hAxglwMdM39erN72iE6Ua9zGHnYuRahKmFmVteZlrdeiV3av
M1xdv1Cfhugr0Ude4J82ugeR3xxHkJcV/sAaSGROdppHaEiIJJtfu4soVV61
zGjFxEnEWOf2Fiwr9UPdRPmPM28LW87VPRiiwSjGn9MnoV6yCwlHpVRMzTfr
kUB6zqYIRN+G5RsAnky1y2yRaJ16TroMwxCVtyOKiNqU3MUKxqpPTlAf2PvP
JdycqMGn7r8nlsW/9pGeaoCnI31nNcVoAKrWaevECO0FygA5QdCkoqXYFLt4
mOUex9z+wvM5dEYqKKEd9kaL14jykzjWFDp2mgxEosPFaMda38hTIr8Q5IS1
Va9E1rPLLRY7TIPC+RN4lKTjn3niQ/XEEtNy3Sjmh6yxuoDV0ZiPaaK/wKQE
HGXsLTOs8cbY+CVkkBdwnYHiA2aq0AHF1xzN+aQc8Mm723rU/2pX4EsDPq31
9RAp8FzV4CkSkA0MqJo+WvOdBWsb+GDR8yTZgvP60eEYh034jWXjAs57bdMF
a6i7opvL2y6S5XU4gcLA9vXNluT64bYOIdtJajhkH2CjWw8OTy1K82Jk41V+
EOA6H28lcSFVFxpgZg6hs3CDjin/9bam2ZqaCliaRkqmD3VjY795wAx0rFu0
Ms8tZIKnwyN6CvfXS1zu/8NyFkFAqnx1WhIx8TJkAIgYcLdtIyCTTvD3Yjyp
8ySA9eRFPPKebyrx03+08YDHOZSaXZDH31eQfmbqntYlBfwnJGxupPBBGN6T
cwJXT6AElqk2NCT19ll6Y0DNRIPXmHL2OYTSJX+SOr75bQOu3PGwtcz3T2UF
fbdW+vAv1J8Yh6w+1CMb2H/i1EBWa2U0NeJlCkNpNvVTIpRrbeA+VYGHakFB
FcCyW7GopU29vY46wV74I6qx+yVNU7i+LQeODGKwA0GYXaDhfyg/WPXICr3a
jXG4FkiC0Pdbg3+0SxGNIV8WVcLi+BNK1di80Yw9+wH9cT/wgffM2AAjeZd6
khvznEiZZkmia7AE3remrl7saBQFRVkyNAVUSIDWHVsSF5syq+uk0fmEm8R0
GxVNB+7bJnfiraLhJFJ8yYOEHdovTJzpWyVVMmGDYFjvA4ZIcqO9wwWD4OmT
2tWARFOhvsHJhn7/9XvdXY0O1J8pLZCBlaBhpj5ZaDfkUcyy+dkDyzVEIMV5
yTF/IksfcH3HPsatSxiEhZOJxx8iG99LgI5eRfM9mM83Ry6Hdw0B60gNxrgE
GRvM/z0Dzr1YB6xxJ36A6U5S7VcffCEptxnJSMiR7A4q2rOlWxYUj0dyztHv
+4AJkJ6KXLnFtCvYXTwOgZG7u2Z8NU5jTcUbgPDaYZHahpF4JANcBBQVzHsy
g5l+pG4D6h91gmNrl0GzLypz11u0zpWyrRZn8TO8odhF2WB4/4hqIZU6miOt
RsqYt27Jyi24xdBKIKDmDq8/iqg2nN7uhnWnCeqqiOR4ZFBNh4vlV9nhrioQ
Em/O/X/uFZdH9lb7ljvGObtHC95mt0XQvYztqfDcwcMPfs7/6gzUUCu2n9F8
iS8CcLjVeUl2z1nYfn3R9zlZxXqWyXkKqDYaFi1jj/uuVA3kSyZsGaDHeChe
SorSNrj8oEDus8myUhQZzwdhYM7LNidPGdUQPzmATPaApTHouRWZcfxm8kMe
tI46VQSrLnjbeIqHJANZP3ZnHDJvf1stKs20RuIPTRR4hC4tyOg0nryQt3aB
+7cLEZ//lNjtHc2/RQ/Wi2v4uabva8xup7kgzs6VWdUSJSvfof5ZS0ZnILzF
JusUWZqYw3hw1UFH1/zdDqAxsRQpQ9A0Fo3PE3K773QgRiYOryXIlwC4w4Pr
0HhxbefXB6lOyVFssqSVXZcPhErhRLdAHyJJXwfl822qSfg1Vn2pTi4AGMcR
YiYHlUgWMT8A7+d4NEtrsJ80ecNPmaAxaNiPT/oSqMCkhwreKsTrMKI89saz
WHrgfIbVAYxQzP/SZCCvKb+yv7lNV6Abr5HB9nWYFfa0kRD2bvwso1lI5pqS
bQVp3cEVz2nazjGrkXu+HVdgcFSWuMaalmkmu0c8xRcmYCdGSFC6k/O5/wpK
ST6mMhPGCvh/zSKaEvnrs45X1KruHNfFf4F7mFFTSC2afGm2MtROJ1bjjehY
njFWBE8CMxAnnwmUJBqddngmGvm6FgdHI52DexzUMCgUvc2jIHc5RzqRm6w2
8VcBEAWA6v53KSgjq2UYkhN8DeYdQm61cSITQs/yM/bCSYAWlN16Wpz3jIQd
szClKQ2H8VyyiMXAMXTUFVPwXK5Z9Rz+o4zH7RVcI7cnqnIfyrbjwxYv5IST
MCbtaSlznTGZoPn+caNK0wXGcTbHUucrsRepyzW34EfbIVjVRkfvsQGUNeWJ
ccVAv8CwLFaPOqSjBXxYeuewtDMKR/wDdD87c1jv7YFuBC49m5MIP6v8YrwV
rJj5CJLBAFwpLz9PlsJab4lnM+RG+ky81FA8p+rsHMXsHKdpqCkj5oGxqxwf
gtSMaNu2HSmA51BTR+Ugc+65uJK7jQrc5iTcqqZkGspCH1c5MGUyExGpAFxN
FRgchmgAmd8BKwk2qj4kr+TZWGMw2kPcq+tXqjTqKHQCv/6fnLGTaxcqBvvm
qIzSB8C+SLXmSp2xpcIIzucEairbdIuw7SYloRdo2850maCGcwY7grCwI4u/
MJg5uyzxLZi9Ztw9HILTQJgGk7AvYxh4DJkZzsgqstWS7qkmwZZLgbqiGEPk
+owVuFdTbQ/n+lImlxGYzgKVrcrZTxHs4XJGtayQaOy0nxYJ2jx771fI3VTG
4dODzWmwzkJGKsnCvVq+FAuKNpPcZSNKZs7HNsMvTYstkCbJ21Dp+OvuoZMH
4EHlwrkS2zeAPMVdTf6cyHMItcKUPIS2dZvVF0xXztRiDpKoGogEiTcatJH4
lyy6cE0TkwJJtHVe0jKSnNiSpDFmA2SLd261/zx7dDvqDfnuEFCGY3e+YT8H
CsX1WPcCFeqLP6a/briEa1gjkpqtG1Ddgu0boufXGFlvsRGS/AXry8nvyKm+
HDcqbAaVNqg39Cc/r2CLdtXVv+I0HCQW+4Hpz4iaE2c0Bc69wf0FBjZ7FxG4
CQwVbY/3Wr/fhavqR7syg+r+LTMDp+48Gse7zxjXVmfc0vMoajFI9jBeBynp
O0GJ53FWP/tFSD2mmO/i7HAfegPt1WQ5YFKpr2yjNyqyGKfbRsTaPaYSPFPy
DQJH2ECsQnQkqJEdfIOo15KO3EjQ+2GoDqlWqfiVksN5u9e/8qP537HxGV8n
WiuaoFMaj73vHSAXPiLHQnJZ9iwWGtDpg+169fRXwFDeNHairE7nRibbrlA3
Y1yjnl4LoSydRcURj6LhDOyhFZlqCOxR06cgqjBcNG7IqTqn5Pq/55Yt23Lh
JL7v1POrKcSBwmxXP+rtCY0vzHmdiZ8C8YYrk0ifMmiqBZ4nKuJhaiK4lmJd
iQ1omsmC6rB+on2nfPFXIvB4VPrCYHrQhWhmfHbanCLHthklUzKJU7NCTn1q
2h9ktrb7WmAU3sGvlasCNI3acJjcmvb/1St1T0K5nLurv1a54iYaGbs1LSeT
vjqFwjIP8EwOnvgIduy/ScdCUIxSXqyiNBLNuNCNgwUvDUkOmL/Zdf1U0ozD
3N3TF2/hJDHC1vxbFtQKdBWugLYSGAJxIJUsxUlr7/6ukTgEaIpnuOJrWkgE
6x5ZK5YS/MyAoVTMn+lNLvkqFX+qYyOT9QHUDcqruthE4+hlwAaSTF3DCAGD
jc+7FLyTpZ3hN+8IOGsnV2j7Bue0QzzyqZpCa64I/sMkfyrdjmZYiB0yGIUP
9RvSXcSUHi/ttiVf8ROo5gAKArI/Ci1rdVq/SFA8sxNLG3FbFtROu9AkzjBv
+zDD55nBYmzfqJGX7ZCAx8OXOZd37dOdV00iGm86Au4QCrwC8BHx9XN9aF3W
H/tee/JI8TIxEQE6iU1EoTcqbQh+WVM5lW+/u9HjwEJ8nUX4fT2tLY6MVP17
LJ/11TzJnbM9/S9PV7kPYFS2VInPLnyAWBQlt8N51bJHa+OnLZj+vhsXNpT2
VW0gIOOH84LRHy3A6yga3zoy8UfEcIYM8TgR/dvMhvjhmRiTIr6Phlp3WlPT
A49mQYrkD7EN5b0ExuQOvRSE8+zJiQ+eKqmjSFBnMD7aSXtpkD5QfzfR31FM
c8enQAYOK8KQK/H+l8+6HohKNzcLqwOENPPuI8Yj2bSJKQAVSvUQ7rfO9D1k
Eiap1Bk4pwBadApTAChg5i/h/2mpV/g/aY/LC6ijgvZIOmx5tj6UtTTV3VWM
d1wdT4/Jo4bmQx0909WGui3i+922iW23/uuRwIZYs6UxYPQD56+rX4vTSvQI
1Hk0LKDJr1PcurX3qpcpoVJ6nZFQgxBrppEou68XO0PQ3/bLIS+fDTJnxAFP
wKPykLokcHlDCdHeiayPfdgKWGNCMR3ennHsah6nMAUVZkj3Q/ZU6aMywRZ4
yQO6toaazROEbyI5MntW/vqHflI64qESX8COuFr1iEY7Z2RZLwLlxZQwVghX
Mjzg2WuqGjdj9BPqNm5mKUSmgfk/LHln663Tk8lyv66GrrEhPvXBdqk6nl2B
jk2dsnXSH1GEhhyOLAsmkzVAuzPAbO6yH0FbCA7ZfLT70GZyZqLllahJ1i8H
MHxFMmsenzYg2xA8buJ39XKz/I7zCk7ueeNQfPRf16g6z4Ig19APy1S6pP2/
9Xislc/YXemYH6Brp328MZd2JlwJwWktq00CAMhelVkQ7GrQRkgSqpWKnlgN
9fwcTpl8SqW88bwKGJDgwlwB6U0KkcLuhQnk3AFAxvZhkyKJJ4BtRH7kf0Zc
YKEpwOxYA6ZAX7y17Q8v3zpCuLyqOPwZbE20S5r6IkJVACiq45NzsldB2HMm
o7UbY6uWQ6RMSMrGETOjZCODq3/XxJPV1AVK2k0++nH97ke3n3HPWqNzGfmO
1+CoQhWGDFgx4rWSMQDzQ1HF8yKcDHr9g/pZZIkWrrwe6gkGLBUj1yy1x1cQ
xXVj1JTXRdZAumBhffkzufhIsqZxJs8XRtjBknuEveKVju6j9n4aAh6XrpTV
b0b0Xvkvf+sWQwAvaC2YX4i01uQhRj76qM0gJ6HJQHUsMDDW+EwR/A0MEz90
in0o/Sf2JXq2pCvDmiafEuvqXBYlFLzZxKObszTPQeSGDlHOAb59Owl3KNVH
dDS+KCupunSbRUR7SBTdP3Vry5fiFjjSW0yM5l2lqYqinxbGyXgPKBMtMyLn
ltLOZUXeL/YxlWEuJLk3b+YLnGit1VAOX2pczVMt4QO083I6nLhcF4H39Uu+
/fpu6O3unpIf4ORFBmNqDZvx4qasJ0F7AXavi2AqjlLj4/TWduB0dz2zK+jo
12vZIha7wXZs+BiLb70DvK9jhef9l/MzubC0mcLokHjgxv+nC7QFcLY6QGaI
Tncj8QQ0Rd+5b2/JN2UKPla7/oQwhsKV8mBeaSZk8fnSgaLVjKPGcRqzXHju
77WB3+VLhE3nrQoMiRIyjWworu5PqeqA8to8vTI6w1gdrRFI/ykKbIugNWfO
sbCThi9NfpkUzzpGqZ5MhpVqirInPjmV2D0fxIfo/g2GzGvGXMYU8k8zh1M5
Agd48vtqDC08uzuwh6J0MbpmbgGL+VbPTabr9JRWIsC09Gl+NO7jtKIZh6wv
/H1sp0D7lp3DhAeZaMtV/rftCh2bXHQl/3Q5ylUzdx56e48PxDAFvGu+7mMq
aRhE0ssajK4BFTtqPL4KxLOB6qziIHWpNOuD/aG3zLBBs6nlcBmtAX1KKCaf
CxelWPwITpGaSnEpjRLVsoe/Fax8y/uRUWHpTXkneOaQsZLYZjn3bokbpD1T
a3bLN5wZN7d9BjdVW4csS35xV5qi3Ufs4ApF/cUDfXa0yxIBnUucvWuBzNz1
DLHBIvpH/ivEIz5umEyvTjIC0JBWGRAeQQbEwhlAm5NTV9FkpA6McrqgCGk+
akKkOm31WnRUt5TiL0uZkg6oTcMNj6npaemQlQwFC0HhcfnOf2bFrx1+evoS
9Mfy4++YOAsn7H//GZtLjok9rPJrFHYP3TppdPU6ac9vND6oJc1p0BCxamZ9
sgh9MZv+spb2jBqZU2YTCDOAjCbUGnvWVc2S620aba5rOpWKwUeRlNYVGE6l
oZvIaMLH0KcyQhGJwCK6TuKXGTEOD6EijCaqi6ozgw+nqWq/gtCD3wCDC+rU
UJo7cCl9MrfU9HiM/DhMlm2LoR2kOlbVlLbWmm/oec+4kWZcwgfzo/Dr/C3Y
rXAWZhWx8CpDKXyb/2YTJlQ92DtxiTqSQaqm5Nz2hMYXkJ9CjOYgrEb/k7aD
HyvLM10lW0YcmVEG7nSFN/cd4WeaO5zZv8x6siJSwZIEXkK4pUPlw+3PQ9Ot
OYgB6LgAbQVYp6NJtO5svvGc0gnPNiRGm/erqnMDS8mzgFroglq89TOtO5ry
JLE84hPTLDawRuglPaXcxrCP01DnzdhIY4OwYUXQKi3Wm+CC1vKdvCnmaDgB
k60AjHtW7q1mSEt0pw1FOxI4rS05wGnDiQh2LvHwFZJK13Q2c6THLzZ/otFA
7TCk6HH1a7YJe0TOKTZ7403y0QIljmZRns4Q4f02Ze9Lc+RQtA4eaDEBcSfn
x/fmsJpH29WJZxdTKJTOi8S505K53x+c55QVmtKaOs9v+Ajvb5Ckx/DE61Sl
jZf8mtvvP0G4sgBM+LwE80H7SoXybsDz9ud9ACOP+bszidce2DS89RispREo
TJ8C7xbHgvK2QeAQZKee1DyDsCjlgCizO+ASnq9zMMaNDlHu0AliLYHApUL+
qVLb98MaQhyUXlY4p3TFYENnnJ3DQysYXKLN9mUyAIHKytVHayTqlmn8nmPN
O4xaLs17IetFVO+fRtTehksV5dSfMmfvyossX4RRwc19vZ+b3eS2+1ZBPqHz
AWg71/2gurXAVDBopjTcDtSj9RSPemfht25qpw3sAJwUj3q35QRG5UENWVnc
gpVqQrZP47rXyBY1s0EPN5uRD1Kf1ALi/UIFkOtWFw2Q1PzK+Sy25brax0yy
/PJcoIwockvToZnWpUDX+3brywqFR0S5Le8fF3a5LvI0V3Qu6wMus0E1m2QD
k71g4sA1NwlZpoakXZ9gio6kQOtViUnnvew/EKLTqKqPVOzpjYVCdkfBy7gn
nCM+bFbO9fdFlwhYL6bguVy0axFeogBDqCny0OWv9hpK55vcBPR6qUZBexVk
IxGtg5LNoG3hqo5asjxu4uj8UHMisi4HumDYRPbXVpjn3OmLrcb9qPsw8qce
8KbsN6J4k/Z9jpgjqLDO3QoySEEbIb3PcP9v5cTLK9nOQmZ8lF9zBYerqVFC
Km3X0KtlAZGKBPjkKkK6ZnJ75JZXLTMEfihvQAYzNmZTnMhtQDQsLdmAnGNL
xccMGbJ0ge/QR01dOEEsuh4Opyzg5j97ghhgeT37YGcyyh4Lqunf2wIPZ1ya
nr+6L/rCpFROjOgRWWX7uOHDyfQdx20Rwvn5+X9VsDPHcKDoO/M/TQlzcHMP
MbwHRtCYcdvZgXin7Z0Cy/r6gpU6rjWZYj91zkBc1VaeLnICDwu4b1AJZTqV
+KAqMpjWlQaZaKQIw+TQIE7oKtBOM5bxC0Yub0iarwGiLdQ9OAeK2fTFhMvp
XqCUv52hasAKwj/s/yctJujaU0AC/uKJE4WU3NPqyfF8Lt83CnoM+RZD3w/M
wveCFxndSvcsXAfdA6tTZIwqUaDsfJCTQLVySq9t6/dwyQBbYLClAW3W6w8B
2p9KfuzncDhG1PR71V3hrRKIBLEAy80e3pSMvrStkKpncQcFEcQn8kEeWIdk
crEsx5m4TCm4QerKIb9IZ+coXmzc2jyntvQo1bD5HhbHAAnD/MUFQIlLRMOu
5M6TYdJMF3ICVimZLZJvbe7drZy5pCHmtTe+WbGjI50FY++P0Ffnfys4SJev
AgPnYaZgGlYZZkXb6RyO9OMGjPZoYKV/LvbZhrD5sOt7dSGPIv+hvI6/yXwx
Rh2qA/ucXWVWy0Pa+vtfS6m2nJ8fQNzr3Akc6MXrzDvsWgDTBudcv8xx8Y71
6OhCI80DXkVJMdud9ZX6boK+Eoe6Agzg+dFBzNewP6ycMK/mIYPmBLvWTTqk
Pepg6c60Jubt7lTvIIpPgCaMqpuYbO+HoKYWNBEUOHxNSUzvi4BbNrO+dR8Z
Pf55nhBdBOz1kZJBKZjqsFQcrbL2rH10Qk+ws3PsZASZ1+NZA0vVlAKRP+dB
DubfO8ZMjlbkX5i3g62ReSccXdi0Ax/hHZhGFX1niAzj1VLtJwOcp0nhx1EM
javFn7fXmwH/tKdh2zNf4hSYtcNmE4Q2w7bMSFKWouWCib17LUmo3ADzeYzM
PA3ZnyxbAadZuI/FtHIQlTuMwbN6yGh50az+yHg+p9upUl0Lh3aV+QMUWGOG
4Bv/JPU4s3wA4fHa7AjWKxVakzrbTRRx5c+Jiz6cCclx917d2cc2DtEG2h18
r5miVwu3lW8uJJdb0Po2hTeP9qk5LcO0K2V9jCh3YuxIA2y9tKNSO3PkNJdO
Vzo9LhHnsR6e9TMO3+vEi2B9dCfLFg3E80fmd9zlG8cDjzC4Js4auBMaxwrk
EMvoDLvJ3SjboELyPxpvLrE00ukOTcpDEun+698Eb6YG/gy221+KJAj+LmqV
jQ0+fHQ+HOqU9FYtCGeuR30A6JUvFCeh66cAII9U0obYAvD0m2yPU4ANPp1U
P+EQ+B2bqv+kL/QJFB8QB3gynNHHZO2E+TfYFv1Mik+moIN3oV9UiW6H6m7S
a8HZEkqEPhU6W8WKTu1lDjgWJpLG7kz32B4w8CUvjtoDP8htoXT+PwGKkCt6
GylsYPaBM6In8WdORYklBlNW4/rwF56r+mWSG1+LGfTQ44KAh3eXZJlXAS/g
A+Pnx7dxeZhbO29oMxKZM5TT8u3WtaF1ZKlzg5NuQbYy5P03FoJktSIvXyFe
CRIYOH5imCboDBJ2aY/zE5r19eF/ChWRWPFox4cCmB+ZCETVRUzIR0HT8Sdf
4n0/d7yycmNIlIcrf2XiI4xq5nd/r+aJi6rWQR865QryPJUbRtGh0xAq0hh9
tCioKPkGiz5NV9nrQhbRWY4P3PaiqQ61q1oMi9hzm/l6O5yWeaBLbJbdoF8q
de8g9pvnoJkaWaWMuLZaajClxL2HXm41KoIyh2rXhM1lrCxReyvzIGmxrPQS
SMD3OHBUMjr6lfk5ilXlE38el/5zxcLZaNZbhjSRguRHvDxXXcQQY04Y6cxw
usUCup6sPodNBX7Fq/0H4lgLFMwnTto/iPnaDFzYxiQIC/A98pbm9GOEzXUF
6Fq95JGhbDxHvvoRfxK49l6jgSpTzpniI/c0j4KVCHnAHZoZlD9Qw6Rex2tb
44CObMdf95koiouTmEQ96QcZRV9SRBUcYIbntvztodr9szLl8WM6ZYyE44ru
GCFVhDcboKuRqwgjWF4eddz3Nd1kRN+3IA6FkA5+Y0z64vwIQ8jIk2LGHjEK
BgNql2N05S7BImtq3YupsZYVixayS0tiW27//Ofk/Lv55woY2lvZ8pTNDH+c
eOS3qbYmCpSuNMK0V/vpPUF2FOruLZebAXA8OYahrkW4QM8C6MTT7B08/00e
Ryb9O5FXZNQ4ttbffvT175HyaRboo6qJm/V+LYcv0+O79SzPs4j7ogRTNF7e
AHQUvMfz1KIn7LhGHQfF7TRZmnZPqYF41iDbTIL5LCXGLQ2NRIT3Mc2YfiPl
1ozZGS0boZPh+POex+IB19/mWZTNvuNC3/ryXP5Z71FnYXL0NPDsWaER0ioT
RH+/A1eOyfkZti0rvXnarhFBVEIoCf/f9DYXzZmCC6FABk22NtDo3cgg2fmp
vjY1jbzedGJDbXYiAraGn9Ra3b+sTlze3S1ru5STfuv1U9fdB/jzFpIoiGRJ
5V+5sU0vtWIiHFm+yrBwrJ1zKSdaoVjxBjQYWr+ARQLTcdD05Pg2MPf7ohwb
ayAa4D9IYoqTENFIneYQv4hCZIm0ihKdrEf27vZd+DR9JM9aYDKtZjzTQ7Od
MeY+8PwFhmmW8dZNje9NcpLvn5x3KTaZUsN5J6maOMqUe/u4b/26Lc5iisfU
zzQceLEJsAwz91nt9l68HKUJG0H1+RsA1KfRf6dM/Jg1G0oysNbbFceBXJEP
SyVsF1aDehJGD17OuN3K1Zy30kcoOPLQ81nIheFdK5VbfrAZumCaVI5nGpZA
s7dRDl/RmpjxSftQJlZYcjD5Fmb84rtfr1vdro1flE9+oYE8RGM/4LESOlfq
gDnQKVi7THIrXzmOI+LE5NozQfTqMB40NnaUBfOfxEChfhLyzO6cmu61uLpN
q03V/KiEq7sLSTb5mjkpXY0BSxVG0ctdHvkGEAChbPi/3C8o/iVQSxidSFtH
RXy+uzfjNFyyrfcy7xGBNSl1Wyr1+vShPyvn4no+0l4EEEePUKLzPZ//9Ffl
3wFov7eOk7wCk3UkV/6nDUjnRql8hk7quE5tzMlzW99aHdnvjujIOZI8ao/i
D+CdHmzd+Az+FVtCkIjb5eVgZw01UGbdC8qt/fC0yPqwIOCpruQ7Patj6UTN
qu9d14rc+PLzocmqHpKrteyCBLbrU5EMMdUiiqBSSb1fUtCR0KKbiwb0FPmd
9GzWraXMVz1j8DBD7SV2bvjTWsWTmGgAcZRJnku/rXSIWuKzhx8yI0UydO/+
cnE6KFh39tcBuM4oAhc6flBl6lz3ArdHcg9I1ueImtdzKRaeLMDOhoNc0esg
ZhhFxNGOjC51vTKvN7KiwoAcAOcvcNK3I8XuoWZDzYZtd89lZ89xTsrRF9fj
a8UuMSRFKh5YGHzBDTTO3MK2vJR6LeVZYHQ/BukigFDPMRdyE7y5jDqEZD8C
rD2rNLEipX6ySC8rTVpVJOKkMfAyQiF/BelcThVXJJaoivSWZooBv3mcYDes
/4TcugfJ8Ni8OzvP/OKA5FJGVxJRCiDec2bt74ndmyPC+s9mvcpbi3+x5EvX
jC5/DkE43Bj1kB0hV6XV9R5/OobIGIIHLfmhBvwCGZ/LDpjENSErR5JpuvM2
ATfZDuSyDlm+fEtvZ1f6s5xlon/insODXPdgyrwdhVnwj39zBlHq8CWTo7yK
2WN2nbFjK8/Thiq3WaHTjY3mL4NNq/9MaI/89AoVUgxgyeqoWhjVq8NLontW
lMyIZo05IZY6JCAAN3tU14QztlZjbkRMxDKVnHRXbvDzEmLLCdXW6duu4flJ
pSMLLQqwQhsVz9f0pDKvoq0JfmTZ/yYxoRvhIvvmVpVXbz7yMnqhvv5X17Xa
oTt4XBY6lKhefgcGU23QyjQEENeln2CLAkjG0Qs57vqwXxlQS8m9SyXy+YTs
u+kFNwm7r3VOo4Qj8nNrShHcZWLzLIo/2Xjap0ENggym1BwOtVPMdXPo/BY9
xRRHPGtlXUyy3SDlYmEpZvzKRhxHvEHyFvzMxaaZq/twb23h13AMKuiUnia4
j5HTQD3+yf/j2Ahi8l7c3CgkZuabdWpFXkYhI2IXYUa5haB2+MW1sYJV245g
Yyk/sqb/dWbBrczcYWqmklwiC5h/nj5BIgo8QjoOWv9uCgNuth4lG9Q+/bSS
d9driyXiPzi2r2Y+IYcE5AbaXF68NnyOwDPRqoENddDaIGiNtPcd8w/IouvL
4m+eJ7t+DEiP7+A4FA4WdU1w3qsN7bgUcE6D41R4PEYi8IeKpS6IlM5rANBb
yso8aE7inWqJEiwt28qbAhLsmy/BRmqJhzhiyeYduvF3HkVkevVMSXi2MifB
zVYymFp+YF4sdEkZqj9iSU2oGspT/IXqNdcd+fiu2gYMnBZPSx5N5Hj70fkv
KeqdeGSuMG/0KE1CXvpYZUslPn0n5Snti5LXuQ1oVsAJ1hMAD6XzHIKwUoJz
mJdHZCT802xkihG/reMmDzh5VAPN+H0fiTIGhyjKfqbG81eydRJ2TWD0E3yG
2LB320J+y2MDHWdqWZu/QmtRUjzBcV6iZ+NBGq3JWmsvwZshcJVt97GLVWiC
ts5gzvSzsw0r2wIvnY+7s3SnwigCbiLwLfZLHrO8LhwNqnjA6OXoc6oYlwF5
Yp1kcyd6KsjoM7QajzmCUolzk16f6M6n+jrVMMnRP/xreXnAsUjUR1mMIVr1
egVA3C0fqnRI+PXdx1hbSUezpCBeJ9nfnmtfzKQEG/yX9Kw1ufL+YFuU0ibK
iTsLmkBvB45gsJRkfZz2G7L2SXrCmNtLDGbkaEFD6bLhoN82leb/dFNcC+zO
x2GUaTzTfBZ6UJuDAWuUAr8o0xEIxwG8H6oAvvpUQvMGF5ksW3iRg4zdQFA2
rcWqvTJpWa5x2rQNMj4sHO6yTk9U3B73P7BuW0Dw0JwccRSXIpODXVz+RJnQ
YxY8CYz9B5o09R5h09108+ss6rO9Op0IGamAC4BSIr9s2aFn5+kTZ9u1fw6C
3l2yW9VHVwsTX/8D8LtPuP9oTG/BnltxZoYYLXlqXU3Omqh39+RMFAESxiEg
SyLgJnQZ4l0riX7RRk2MhKv2CYULdJJ8+4c1bAR4HyVTNB/zP3Kir2sNA+YA
rbGgJJkqgWhVLlW83FZghAP48MzVIerX23qwTNHGaubrgg51btpFzJZeoQK0
MLcdRimRC0vd3WALp+50n26365l8PT/3w4exxV1s7jDMVnROdkgfR30p/vXR
xSOczaMm2FFbDNf24Xp7A1aV7pP7Q71pEkq2GdVyi7HfDnqH3KYzTVpsOmwr
zGphIVh0Elp1BUHivhEsBAJyzgVeypWRC5p1j3x7AKWo7XC0AVYWBZP/9nZ1
vsj1im96BNPy1CIUxGQkghwmPgP4E8uj8P7VycC4OJ6Is2KaxhI8W6aV+sMh
E2Ji3j6DW9zNkPBhyAZU+h+lTxzeSK09wW/yxY/15zbHiibhxjZCgPnTfTgX
MMlyxP4TLW3tGCEdmHJIVslsvhEWbAYM5inWbhdt12PjKcxTsfrSyzTf/rC5
cT1yULi0caKw3Ryr5PL7WZPvhoL8MWacpHJDAPhU+abLr5GUEQE+bcWDC47S
DbRUeqROXA/8iORX+L0fxvCeMqRlPO2/qYZQsw6TZ7yYxsbboSDhIi1pBN5t
BtP70SfEk/c/uQV3bgZx1CLuAZ4SPAZ7q1D6mTjMmtgBS7g3FGsP/DqeuX2Q
GCs5gZq/ZAY9Mm9pj1JUAjwYEHpX6MAyRUgjYtgkglD3Y1nxn5hGLJDhJoy9
wgEZh5aPvPEPWlEkeW+TBihdS3Gawzc4pHR1SGQkwnwguT0A6Z1ZWxOMPisH
bF3vGWaae69RjjH8Z0MlMrp04KVfMncOkqtmQQZhCbW2Ur4ge/o6koXdWo+N
/CxfbK9jUs+8na2nPTPOe+wftfvkTgKnOMSw0NaiJxRDycrfl/v93QQMpf9B
by9u8Nh3MC8J3qqQiB6HrMBSxgIhqZDt/AbFY65/pzfsW4U12mFDzmAoKBl1
ufBHW2LDefd4rXLwopn9iU5L4dCBQxHa910c1BgKcd6aRiz1pQH5lDR61AXB
oNxm1MaD0BD4JW8ZzL5A54eg4HykFnbND3kbFc27/7xj/AiBfqIloqUA4U2h
eodAbNAzgxK6/WFavFYoRLPbTKnygmlWwg8LuY7vaN3F5q6EZr2Umk0/6h/X
Z2/xXSijaBSBvNtd0cFt3ihR4wv/51nYh6eqH/YIPTCEfkAGWT6DzWKyfopC
n/x3ugtOr3DEAC8agmq+FE8qz9jhzbz4fnYIj5/tI9X07ohu3o1fdCTmNk+8
H4J063Bt1W4yYVc1BDHKNVN3rxxsX3u3n6aT0sJBkAi7zNKlDx87HK3FP+Uv
adIEhb235FyxK8v2u/ejY7cfi3f7ZVIf5ETkcoPk+kUVE4xq67RsbbNUfIdY
J+BhN5bxp9ha7FNi4n4PkPsayInnUxegAl2at9f7eJFxVPi9D/vlDE1ce/Ms
Vm6spigYIlYnPB2Yr+QU5jweF/VkgFJ/w/Z8xyqoW2WYU0sm/F+/BZxPek4/
CszkjG1OtKpwMpJ+pJMIWQGcc9dxOpxFVxTUA9qcHFKNFAtMCFWQvG6ls/pq
bc5O7+OatNWZVLZO1yURYomODFNocy4WxKx2mQmDZSjtiz8gYEn+G3RCCuhX
DMj6jmztZfW4J7lyCOw9qhfg1rYIbQkrQKdtXYFWoIci0JfQPqyYyTScpnOz
8FAghy7aTylEfy2xqowjTgcJPc/7Uu4i+CTy77kQ+MzV4euLQdnspISYejQr
2t+8xkbhQ8Lwxij2Yq6GrZ7ZH7YeDo71oP2MwypIjbIiGS+pOvoS3OMybE1/
qGfKiezGtAyPJI96cUg5+m94pxIzybmNYQA/xiXGykAGafn7RnxYriVVBWxZ
OwnFKoEV26u1soHQRuQWHSX/pP990zQ70jBhcJRWeEZsSQIeAAGOWcM2GIde
TTr7orf4/GZ4WzgkCrplbRombsR7e9ir6RYLlnzF3H+Ma9ePtojN15JJlLHL
0XYtqE9etb2P1E1dwcVtWZBDSasCw7QmeFuW/hLdGfLj23AE3dnkA4O0uHGD
O3TENvnnC1MhKCD6uRGqDWZpG/gCxG8t/lHPaC8J4/9YYTOefk11/xERsrq9
0JAPY0+5ASDW+JiFjoXQJb+N5r/dZ0O4C3vOw1+TFsHB10ajIT+HNAX+V6/Y
HNTRQPtlWoWPDoBELcEn9hD+k1oxafzjwovvszasZH98lLy6Z1h6FQBWp8HS
bgqWxp9IHnd9T8xRKcGm8c8WZ8M0BCCZxpz9sc0AuYEGQ38dW6WJ3oL1bYpq
fnupI9ckoaPBVfdm0yw57O7qY/qSWXCzOqpqWEbOxf7fBdmX8YBXEgW1iQG6
w0M1qIMvN5gxiz/lSDs0QnpEklQh+pxvohRcMiwSHkX3vLnkpDgfJtw62AbW
jMS5laIAyjyPLByC2kr5P9PDKWD4AVRQFUscMnSRIktHQis4euGvu2nl4mtn
OjnMkg/Rs+bV8ZUahkDAOAbKwp6jeUSos7sbSJdtQ2Fmv9vvFhrOypTDJ5Tn
9/p9K1H8slYqJr4qu7Qqehs/NEit4tVEiJuyeMpvwniHxkNlNrguWDVQzAbE
wrKx09TQlPW9T72jcfGuC2OyvkXUKqdHkt9amLI8wkn3yJNpc+BqYG2dasH2
MzaDWWX8U5Og3asb7+noWF+L3nkCSBrw4CnxjoN8YU1OXMcE3vFpWmhlpLkR
sTRVi8dTISflELBl9mxm2WfB3eYdfVsWy8tXhABy/AUM02LXepdsqxSp8qDi
yWCs3puPwwkovmfkuOGxWB+C/qmKsVfHMUQvbS3N9MNB6BZ5B0ybfuKGNc7Q
oWkapvx0REV9RvPZ1aLgeLYsAvRK8qZf/1k1Ky7IMSNvYImTIky6m4NEPExL
aekwcZnAVRBo1OfeD/bkUbo1tFrLdI+Zx8lREH8rI6NrJnI92kKGx/lwGnDE
AuChGzwlWwx1SwwbgAov+HVj3Y3yHK5utKNPmJgk+Kz4kiPEsZl36PeITctT
PnpqGr6IRFdNXLShxZBzaH0hM71WXo2moqRAYS/V57iFDjq/9QfGgISldb5x
Q5mnt0YgxLs0ZaK9gCSoPb8UPBcr3kwP34ZnJSgAkdYGgxL5XV/l6ZtNr8XC
uNECNxilh2R/i1ckQKiq2xNwZHgw3zjU/osfQlwjSpHUJhR+h1ish8Xilxt2
5iyfYCU5bqmXmNiBOI2zpIi2Qcxosr82PGY21XDpOGuwjSe6kPgSyt02CVtf
Gza6XS8UIcrcn2IVC6tiWXcjtu/V5eqzc1tX582kf+fx4sNI3V0HHqxAW5YM
V18yd/g/E7ryCHlxt2kIPIWfvM1GrIpwGIlyYUrDucBlC717szdHUadMlYou
+qvbAzmogyXTBvblmreR2uafMDHQ8ypr2EcuRQzaGemhNv1T9alvdK3Nfr2z
6tKnnOfVLZnCMSE2Tavow4tKnfCL8doR5/HyrFocnXelcivm0UWLGAekPlsU
moc417/S58Mt5Konjy9A0KIGdDQVe4X6W+qWiMObqoLRRroJe6Ts6LJXmssy
Fha/ENJ02FVasPdXG452ePwcdVJjltoZtceRqVOi36pTwdBo1R927ceAnUQH
0u06i2Vj8JC63VuHPPfhJNSX9htOVZ+WhCQDCsyTQavLN+bVnEEaLUSXVIXJ
MMe+zVGkGIgQIS8kh170U3rRcC8XefMyoLFfSW1JxI3eygCM5hGeTa/sjHRb
jndn1o4HlEd0osZXB0Y+QPeW+9VvPoqxtyaLYExaK3Vqdz9j7iYh3IebshWV
hYwAhbi3ZX7XHPGXJJCzn/w+G72OI82bbOawe8ui2tEZ6pw+GDQzkshdqIMV
0KgS58ZL5wHywZcVFeogMI7GkMMv5OxaJMdD673bNNkxBWbS0qVPt2MZpUWw
4JZNztoRZikM0hltw17dle2RQW53hFX3ec/+wn3P4kvV4LkH6VFusYN6BEAu
T53Bbze2e8AqlvhSfVSd0Jo9gVHW7PP+YiFYiMuZhfdMF0IDMu4EwRfWo4Rv
DXyMosWw1N6W9cWYxlFzsjQXiWTZTYsk2dXsdn2Le4VjStopV1RB6XrfCxnq
f838pu54IKLmrRCg0EcqJpKvcAwDXniAw1D3QSxbj7zdiMC8wfZ3oHMGjajF
2FOYh54xom3TrkeQPAHn8mn2LAah0MrVtPuEFLqsA7oKBLa8RCJiiV4FYcz1
i2VUchRO6pGtENvLoa2DCgQjb26lutWQuVRPDxI8F9/Ry71iYVnbbqhwBBnP
rpFKg+UxDOiTur0lbnPrlo0f87KM/uZCknc8L9TIqMPGc7VvGXgNMNe7mp6B
NQREMXdwr1oqxdkSVZYNGNCe2rBo9N8h4ZRi2gkQ4vSBLSSnv22oQ5im0Mq/
WS4yLZKbxZWA1REbZeJrqY6mJJuK5G1YB3k2FftjLa+ey8hLVvuH6XXzPsMf
C7ixfGUtB1IYCJywKtuBZA2deAOb74AgckWvmIASlcs9THQitAUqdSF+z9qU
nEfEuXeL3IbIO+pUEeNdXfw3oBfwuNzWrpiv6OGvGjLq1EaTbC5WdMbNS3Q3
bt+psYfng4N0SFXUK4d9HwEHnYdNQc68qEdkPv9CTQLScH4Y8zlRemrJgBX3
Ctt5sNEhfbCoNQSP2jTDY9eCnuF113SaSw+ONM0MrAuu/1EIQ+dd3iOfnKwk
lCj1TquUAMqWlvk76jGzrHjQzwrB3BUtyNHI5UuC6bK+ZhiHzg6uo7eAoSV4
1mRMOHk8IrL6EWoAupmy5taFFhGctcKfaFYg/cW9Yw89XLEV3/RbKEHYy0rT
hCpAhHy9Ts/WrMlBfJ7w9AOTr+4qBMEZlzlJGXmYVrAwrFu/jWTMGtxmgV5N
0UvoQBEPaC+hbq6F5g3vL1q7S06AhM1riedBqWbVbtvySZ7lbjX3TYBeoRy/
oLj11ZYEBV0UN9kpWxJR2m7zK7ZD9Wdcpd+J4XCi/83IJLCQoyClOI3dudgZ
4g9HsSp3bAAcEtkmHJZvWnEPcPBZ0ycPsXl7A5nemzCBwGSSitIplAVYlhA0
m8EXaWne/bdvhASsIaHe2ptEeMaia+LuIo/twWcr+leXaGBoiQhR/CuadtTz
QuUVMw8v+Es5oUcMbRsuEtnaz2JhCEwP3VFhAOWMcXFzXn8JTmnDkyyRZiMH
ucb6dpCTvFwGdX28BGWuiP3IZop2mwuxwFS6oYMx3mSjSpR6ipExNogzo4fA
s9JUbTTqtFIFi5vl9qD9Zf32eL4htPlJPxK7CDXzaK89ERVhSqgOd0W2F11w
iwvlTZoC2LNxAoUfh/2hx+nwrfRyFyGpeTroiYCXP2o8qbxELubidLjI6/A1
OeOlvE6mCSa83Oz1MYm/CjedrHGRw28Qe8DNcpeUY98Nmj33FsZCg8z5YwcX
TwqcIcYIIQAzlULqLb6piNJEj+NE89HtSEmAIVElN7ZcbhjVJcm9m83tGKHP
eLL9x5lemb31LDHQGUNdbzHFfE8OET+9FRfVn9t+h2s2Jt09jYU9M3NtlUdp
4XCeHDTWO3AJTiFDGEhDlB8IclkDyUSslIstk3+Q9YCnot0CgcaE2Yd6H0g/
4bUEsLn4J0Hfx7AY0hm6T9wPDRHvphJhdSVc3SLGcnqQHz+bvu4MFCe6/lOn
QcRRgQ4wueIqUob6R148UMZIiu0W8lE9CQgwQGWhTJqvjzMetm+GxfgUSDlZ
3LaWwbKTrtwcVWmWbmtjgDDZf1eOPvWDYCEyFv9GoTe3vfNCogUXEK3hAxsX
Ls6lOuZgmpdTJXc/DBWtucYnU9QR6tYYzbCnfHFU52h9qJHd6x3m0DbDkimZ
Y4q+vcITMezN3YoSm73OG7ImoA31HR3JapI1ahTFrlNYw+xD9TZLrCVaLUeg
mWRgBcNryWZJKcitkWxexJvIphnis4/ZWja7ZLBi/fyBOfZETKCu49A/KOBV
TBkEkyYZbqEjfCW0qTZSvtBzh86w1YCypuFd++pk+Svpt6b/jq0Spojij+O4
lsqB8xY6RzXfyMY59VaHw94fcxYzovuLi9HC6tsOxKM3ZROJF83YIPdxYPJs
kfblWQHuTuWrsPP5WWB8jXm+WXSIC1SxJW3Y386k0KxdCaKkKPa5OeDFvOOO
vwOWUqfBIgYRqGCUcWQIMQwKCgjaP/zsBQabkeMJil2FML+/Y8C6lJanyho/
sF9VZmZOxlGUekxmfz/msPBue+ahAB+T4+VjHeyxDPkx1DDSyZ3nzvv/uFgm
OdfnpI5gnB2pVIHP4Yo0BfMB/D6zqNvO2rOfdjwDdSl4KdB+/HYTSjh4ujUE
tRwvilD7cfz6/9sJxR7u/il7IvsKBZ44LS6Mi2cMOBMKbKnjn2AORi1JngxG
8f6e70qobKChfXmM7+hZ2MBP07ZA6io5xg+Ovj2lVSWc9M0nP/7Gmi8ErALE
V168uuBI36R0VPQZy4qcBTfWUCW3RU8ggW9XOZJOBcxe58gb1CIpQ+PtNipP
9amAiW24XvRQOWRmly3Vlq1qfVELDm7RY5dY0ddQbLSp1dCo3YpBi+G+EBXw
BkkDINgsjcsnXXV5qxCzat/A70gDCjmX7fKQNqxpXGOE40FRaZR1AQ7ywPD9
GlDPPkQVqIz8oAzMxmhLdwxcjMxlXm4Aqa9uTUXTdYzXtfdm8ZwbIw8e0zj7
lC7jpauvDYsfuHNzCKXo/vLqSFeeI7SBAteps7cULbt9CMEs5NxWnesChKy0
jBGwoUqbnOpwp5TlnHc/9dN0lnZRpD2Gtnnq19sFNjoXCfPmDJUVsN4is3d2
2NdDM3MIsn/OJqPVenny/zitpXdXOZM+2wZk12nZ6jcbtNjKDyMTy3Ee8aMW
aJCLmKlI3gl5sAgMWkkkvksOp6E6d/VkdUQ4avFI5o/5SUBIeG7UcZLhNe18
HK2/sA2XfDwpHQK4OGxlw2iUR6qROlqlABwdhNosCBzVrnch3gRfdirMkh/t
vOCE3uQCCtqJ0fcJUoEd5LW7BipI0d3YvIPbEPoVR6GKV3/Z58T9RQMk2qC4
ivsDT8oG0WsHqUwJjBVQSlvq9+3FC0uYFutIW/7rMZVAG5BNtSQelClzb2yZ
DzInjNTDQpXkbrdOd+Mdm7v6+909LEzq+86lmuICUOXfj/jyW9afRep41y2j
p1G/DsOa0krHgn8pd4SW1OU3c1sl/2i6sUsRmz9dlACYYuxXrCd830bx/BPB
hMTQNCC/JcMVzFZlH4nItPavDE9FlfQzHrcIqsNzjRpOsuc78x8QyNDx/Ee3
kKghOP5vNxkM5rcm6Un1LzC4G3LMTsMMElwuE7Hx3W/b8Xg+xumSCr9a29Lh
8bh+F3KPBYvjbCsJd1jiZlRnwz9y47c1KtZb/oO5OCjAOLNMtoJif0fM4p6/
LLXFtPRSOdzkp0kgI7FVag97ANkcrDJNzB8TT8cx12ns4/nDhnUAUihb6YDE
MXtoxRLujljnAR+WE9B396TXYZzytDMdJsiFPxQmprqN7bsOxFNA3969How7
Rx2VaT/q2bCbwOxsxYkRUWFE2I2MxLCyvGCR0vBvpOPUzxTuix7GNsE6qE9q
yCDYt+p17D1epcf7N1H+Fgs0EUByzdoGS1ggA+xjxMEFhcL8m/G3z1FbALv5
6WpVM/rDMk1Qv44fteKaGdLMK7xOTo3UeY3cFiFVJq/EW/ArzaaEFMXRMbfd
QbOtSFkiaLcNhPPnuYIva9d9qduByPNpdqWgz7yJub0t0u5FzyDja0pxJyiC
dxn08/83TGKNhDfaEvNfmhLWaXjW9ZP+kZttGcX8HuZM9ZFzTpXOKWPvRyIV
VAf6mRr05OaaBeLXXiEMyCBifJOauTtECa87Qck8UE2lJOhUqUSevQNLKblg
O9pxczkpMiK59fnUNyeHaVynv523tmuVjQw0n+Chus12/+8Ax5Du5mk1DDtQ
SkZmRkB0CtpA45Nqw8U6bU4nzdXzqTOP63obaLUnm+NwPf5ucJSZ803c57Ql
FmWRBi8d9r3A17LoFjxDd6C51OGMJiyNVO0xuFPi7zimtXocVzjwZHXC1QmY
VNP3ei3Eg1iImGpgbZ5aDUcq0giis9U69ScXHMd3fXrV0FgTJ7tsWISsVEbl
sq5ZHYZkSkG2oUOpF3TiLUeTRaSmmLaQZ/Q1zBP70kE3YCn7X52eUynZ/A0H
mhI+Wg2+rBjxWluK6XPYSSvClQle93BKQ1ovZsc3eqmutqxFsQr25e2o/pS0
l/3xtjQofanQy1qNqgdO9JE4hro6/oH/uRrO8J6Ozwi+bfmPajHOKC6dxbtm
jLgZMr1X0s0vlveHKxZ5vZhuqpg4A7qL3wFNxugEJvK6//yka/IfA/kpLPTO
bO8CckNglh2/cE3gmrnOimDspSiU/emfJ8923mlVzI3y7kTrhPE4u06Zfd0M
6rqDgOnMNT7jEmrwg/AdDOOMSEueldJEqhHyPW4OCIAs7qQAck3rsJESMNkE
iELARfOTX4gHtz5QdGisKA+URgoqwHxkOpjysZSjiHTBLQsDqCtoN4s7QZAU
22o+O3D9GbZdwfRD6a46KPQ/JDzA+PPLhvF02a+arZvYZ3Wp8lQCk8OPoqoP
nEgsa/HDw9Dz6wrBIFL8YUO0MZdF5aBx4vwtoyAxt3U2WNFIByLWJHQMcMre
wxgROJc2glgwkLYsgg/HM2pM7dEpqv4Ibx2lifGu2Ogxw0UXQTnJXao0sjUC
o56TVB/G3n92D3ZXmzI7Ggz1w74KLJqZ/zYVHM4JnMm+dXy+xk+WJtRs14UC
2+sIqnwZQB5UaKAeJNVe38KZ8AJMk8mvu5UtnirwphwhYpq9gT9P6NnVwGbd
gjTWFYcnWo4o5HFH6+dh2637lZdwgNd80G+i1jB2BBvg9MZN5BaIKljLIUD7
sWZHSbHqop7HT/QN0ZOPM3DyQ5TSc8zdC0kT53jojmbn3T9VpiKpoIEVuQqI
XfG7k9iNG2t1qrc3n1FxRFx/HfhWOidrwWXHJGI6ND/8Q3giJzbljGaGvgLW
sRO2WBjukibmPqMJrHQQaMsIpdop0O4rL8ycnOS5n9Q71rk6+suJfYSKU9Bj
dinUbE9XNe5uPnqkoaIGclOF3Z5fNUAoCHNahIn9kiisEf0ct08U22OvAb8Y
VAbgAbjWa05kE7LYWzxhnTtc+4aaefKcw0GtFxDlht4FnX1pQCq2F1E3THl/
DuyeabtAq4b8qsNu7jFPo8lreCfUA1ExBg/fHRDK7L5hhx5cACiATz8Yb0uU
JJBNll8jpFVRpWWIJoPlx23dg5rZOPlht3RUUSAKnWHe0HW54CLZBN2JPDn+
Q5gSm1aWgOdqFnktaVPMJR9x0jhvntUw5Vu5iT7iPoAaJxamJ+5vAeaUESgf
4iwy93UrwogFi0VJzw/9szCTqkQ02eeLh/23cf0xJgNk9AqtQw1GzbitGWS0
3UQsylCzEFRTD3XpOtxsX1KRFaEJCD7pxgnthYk7iN7Zmz64vagyM7Rwjw9B
zA9d7jSzL4ZVlSt+uXJpizwQzXQh46v9RnQ5QnDqxrphQkYjXSxApg9PrI2J
hMvwRaki4/+es2Gs3irYlkeZoLhoD0r8qndZIkvbOLa/G0kIKSgj0t5aiZfa
GqZFl8snYMwRs9jzOkxssdm+5GDT2g3JPi61v/2ei1YYnXyi3DYafo3OOlPY
WrotxNXeP6FLJ5KLDnW21BlZRbILoIxuYukZX0sK1aYUSlyOHg+rxJUFiK/R
HKlaGVJvi3RQ0pyPKN19N8ge8axhKTGQ5uT6egtCzJJq5y64Vt3e0nLpV+Iy
i0YpXY1iY4pDCD30Zof3uAayspOkSbEX9/VrtifWCIYTb2j0KU3JXNTtrrIv
p1PSVGalMLbMffV0JxYTY+xF3cHIojVkX/2+DWovpKBtHkMF40oHrQNdeVql
FC/iQwygarPGTSE2tiz8t0mcx078iJZTQ3MgmMviIZkNucUNR6LgCYuSSluS
+RnnYEgzqQTO4QTDNuoglFJC/VG8jOCzx4gL4oGs0+fpuzyJYjQStFHV/dlp
WddZA3nAmPfBk2TEQ8RG4jZqRyBjao5sYIqm5TBciCU93BUjCTJIAVpC9mTX
5sxQaigwuwRAT3gkoq4uOfyz/ckJ0v/E1Kiq/57+jxh68xPIJoTeIl/NK5d+
0pR0h2V9cKOxmZfg4v6js148OWSQNO1mrl56bNGpFqeFFdJ6zxemjS+hfy0P
2kkHA7yW+B8BqC1BX6tEASC7PXOzgiokqQjyW2FHiWtBIqp3Oj399/4I6lk0
s6vKTqYNOFRC+t8DKx5QXRm5CxcFTuoBtPvg4LrYuS21vKFBFRiAyq7ItDEd
qk74pDVzDtQuHFSuPS3lIXabIIifFa4qEZrVa7gMJwkGOLu5AsdbQWNFORno
8VXt+Y7N4segPJRxQR/JSGLxg6HmowGuaAtAywIZrsuHtfvM+pK1vUBmKcMQ
B0yq7vSxzeJyv7zbpgFM4epO56R1AfwwnXjYpi02d4wqabWvVqwv4wY/CCzN
kvLHY2CHjimW0B82oWFe4IXNiC7RcB/8KJwXOIzlXGHzTaQDdNHuCOPZHY6B
sx47WJeNNAouvdL5bpp0m3wzbaTm5jxhhhpRN/FxGniNJCrOMnrMoM1bjcyx
SC//rfByuzOFT6RApmIRh+Gjwpn3eR1rI/yMhloh8h3UvtTo6o9sD07F72Wj
D2g9xQwqvUuh5Px9KOG4yufLwjInqCY7ltB3UeVNB5xexMcJx0Gv8hOtRab1
ZyyF2r8lH2f8glx9ln1LdXYS0P0ykmtphxU843QnLhb4UTFgm5h3MmHBFajG
mujeLAbJmf8gG1woGu0WhemKmjGeLPSSBcd8YhXWbPo3L3Q+2DUS1deNHdJW
Z0o5Y2DveYLccKIDz3pagr7hUVqzPhK4exydyxFt6Rx8UMjy3kOJsRj1EyA/
LIoUKoYnCZPTcd0yygRZzkW94tC/1Em1RtXMfvbqMCY87JbotcR1IuKEr/lU
KAtiaLm/WRNWkHiWDAZ3I3exsgUvHcLaj6wqH4GiQ+pBYuCnmSgtIm46Bfyp
bGwt9UHn9UEYZ4rpiPebTxtIKEB0geM6szUSBoGEujm6r/1dyaxTxGiprT4J
e6276BzlZ0NAgH6Dz9MrBJWCgb3/J4q6eZxHztmigNnmD9g4tOUkVMxoFXym
5JO9i2RlSdG7u8TMjYI8UPiFbnpezReP8YEbio62SE+L5w5AM1PvEAlp7Wdb
fP1RHavbR2DwJ6TcQIAAcCeUjT51NhN2QQBCiWKEQjh1wWq7HRSC8l+wOZzs
r7lzVZj3FZNv0ZXzKEaDPLv/kkhZZZWIlNKbCMi0mNSmd0z++6Ogw8/xefJj
6w5EEM5nqq06NOqJgVXkjZ4KYPTmbDKUNulw+37CKL6o6CMZOReM4/6Ics9h
xCWFcAxJZ42q77r+Gg9s97Ufnq3zmc+vOvpdXp34GN2MGXZL0xfFgb5j9zZb
ZYaijAOsVoE5f7qXKLwqNUzgsq4F6d0H1wJdQUcdvNeBeM/IG1POAn3JhV1j
PfGVRrnBPjf5Pb0+SgVG9/nKmErAYp0SoObX9zOJ3fNWp/fnkoMDA2joTmC4
AqoiqJ5fZGzBnOLpf6QjAW3OSm8Yu/pTLxUM60FVQuItSkkuR6DpUS0TBJEE
cPLeYn/fX+5imPA6OQ1zuG+43Y4aRE1DLwhv+FQ6l104+GRgwGdHELgdhY9P
Mkvu/ZfDKazS+e9x/N6y5s6BgidPSNewrxGZLG0uDZexHN/sFex7q1dz0JG9
+KwPzeftiGT0JaxJhpObh+17AsE6tLRCa1qzLA6CqP84CqDfOyWKgEsQdYKD
W3KDL8mccw1AmcjY1Va0dkHKkMohB3erw/9DKKHVNNSN8b54HZhVyEsbPxNw
OwiVVQe2O00EqKwmMhWeCNfPLzFHe5F57kaELmRfzIeGyejeVOmgn8/yR1f1
wCKt8G+asPTssnwlp6cX/K+PNRUAlOHRPmWnw+L9tsNfc40y1qR/vYvE66PU
G4lZvUQMg3JpuvirvL01dZw51yKBPjtEzBAHAa7paSuvI/ZDsHjAdYrC3LLY
KVNQZA3KyG8AdDVOx3+Q4Rv59JnQk0ZrijlsoYEbx0I2QkL/MHTiJIP07uh0
ej0tbM5HHdNKvRa0tPl1hhNNqLgrpwxOWQgwLqaQmcd4m7Z0co34iBo7NowW
P2mHH7a/MAOAWcv6S/f3JsA/FZhwSfK3SpGhH6eh/qvd9y7lH/nEBjSntI98
iCSyyG5StvAadkZDTiNeeKHgq9JFshfJ0Vov0opJwf+3jlA8JiSC6D78b1aX
bvn/EU38EMVMyNZsHfYAcxu2RuB8nsN8mVVEegGONyK/DoPurL9TitpSv8sm
olWfSf6YM+WXS7q08iOINSKjcU1/eAn5QvnMQC+pjpoZd9Co9AFvtZOPzkTW
0T57j0yhd4wTAtEC4tsNMXScoDBhd5mQZXB2xfaP0RlabQJyH3BAHJZ84o1v
L5TfPXT4R9HhbHb/vuCDMwGQOmnY8k6VkcLDSkTAyF1lJezvOdIEhjPK2f2W
MYh5ckE/yivFU9cwYzpTivbuMVFR+6CtiUnFvYEPWRiuYezZU2XWInsjey/h
Azzm1E/NNndhHjZtz/PBCHYvH+oWAxOSSscl3tdPwaYaJjDU3zXM2MRu1q5S
KUn02LnyEqay6UzdL1dAyz3Gi3cmfoazGyZ+cjdOze/XqktzC6CkSsomIsQ0
KOPj7SxB8S5FbOgWCOu1G5ofchmXcKPDDTdIlJIAJH9/lbrc3eNRl9R9JDkc
ReMfYrMTcJYkd/1L2Q8MEt+yXUc3un0JYWOAX4i4wILnpIGlCT0rDMKbLNHZ
HlP8xQyUr0QpIL63f+K/H2zVYcxLufL4Z4yow+5lbwcz5selHBytQ7JFNLEU
yhie0zWUIocVuiXq7CYCfQxqLJa8wWw1zLXJrivu9v4GIAIBmGqCCDqaEz2d
vodKv0n95ogZVB2pQifEWMtfgPxYPVQhcBRZml1oYO9+kN+oM1EiDpVx3Zdi
ldYH+zLd+ajItfKFhZeX82LPc1IQBVYzFMmofk4nf7BdpIsS+Dnsj1JQzDLa
BFSfA2t7vesdPhUowLy5oyMGXdCsiAXmti3Mk1g32BuSTXvOmiWB3MbOy65o
8s2vJkyxTteZw3DyVvyyBdAGwMMut/N3LQC5GUiW6srDZXEl6qNbn7edebLJ
C9DRuPoCgyCXNS/Z+k1a4CMg7ZqRQ9LJxC6D8fytKYnxwXeVym+yNIGtIV4Q
RI6m6Gqro2fYpOG7n4Xalo/q+JREARi/Gqn8SD6L69RxbP90YHH9Vsm8eHz3
uTA6+L4IajNAFxmGnZt5p3N0lBaeK6qai0nyNQF/zkZeeXJPyZdfKuZxWb8Q
//4ZdbIt2V3bawsukD12hCz0czy08WHhIGg5v6dKF9ZKJctcOY7Vfw+NMc0l
2Aygg6SexEP2wwnbhyUCLJnqJIQpLqUHJCa3ThXda7huYrZki6EmmCVn7BQ/
IhCyGl1KfeDEwzqNeGDzpK9zC5EwFWn/t5dbCzuIws2hunIaVq2KHZnX+j2U
U9kpaEXauNp3JmN2I2COSfTqzmh3R/tdKk7ztX3Xqwbtbwj0C7jU9VKKupQj
MYGieEuTXgIUfZFj7X5lVlJXWhSwYpMM2FyGONCGMG8jH5GjZVQJPL3Ccp2d
DViBAqiaCuLgIeDt+MzCxU/4SwpMB2L+jRIHVKOW9+1Ex+PMrgl3qBcLlFFn
I9EaFVBJC/ot2ybNScAr8xiR9N3oEcKM9eGpVRpQUtO+H+s4ECyggFizW33P
rc1m3HinGPuWcGuRKsnrPuhVjqPDgMccSd6NDrPipiN51VGnALTpROfdcdr5
dA8Ch2DTqSzwKXFiEmRaYwcYLJRt+t0kov0TjlYOgoV9kqyXjzwiNXJvskN2
7+ELRlU1U3hGfQ7rx2KvMGwXq6tH/WFUOIdftHXfZS/OXJG2IOBwGRou0PSo
+dHBOjY3ufEL+X7GBEi8yugp3qQMQce/Vjlz5tWaJ4pWB53JuiSQFCHaKefg
SzTaXwiEAOYyksa76NIDVoiKIBQ/10FBDgnz9dtls+J7+3EgLiuUY9/7c/Lo
3rir6QbnsCNOhvU5Iaphov4x6ymN7mIQYP6/5SJqcNaLVsxJJ7qI7s+BDjzv
ACpqny4J4CGxptvupcAOHM3N8eB4xFMYdJAipJDtqwj3NXodxH+xCjE1JScv
8+fAKee+thmmXOIIzqZe82lX92dsTdcRQJWux24fVOuOOJcr+04/FhuetCAn
KbCTvVWaSZ6BrtlhlXwj2I2slOQSDaCrnhJlYlNYifE5H9iArFFDu+RX6ms2
HnOh/UP2aZV5G8MWHkSLU2kiwWoUmd2/4BL2U47sAiPYCry/w+wJJXaMR8/l
IDD+oXgb6cnBrvKe6f7MiKbr1w2h9FlvWABtOj8byPpadJ816AmzytcNngjU
hlycmvsEkhiMUJTdwqLpg5gF2lxbL44WDe0Nuw8i2iGNXx9A66/lTWPW47rs
XLjCqwibgnNGzjak0p1ANvcryu9AH6HIJg5MpA4PW3E1Av7YM5TpSdarlt0T
9y/yvc/kLsnDSlWFo9xKo11FEWReAWrDB+VT4iJnS53TJAcy4149Ph7v31dn
Mp3dYJzArYPEL5YsB0okcnusboSc3Niym4YLomE1X9Dtn+yzj4m2phwbnFp1
mwqj+USKxgd8tNqgleLrnVTkNS4dKSYlhkZdpSxN7yaN6lBj1qINoqqlEVrA
9fFwlEbDuqL4kFse9Zh5XI4LcsVtItvbUpTYNSaseY2WfAOCIMG6G4AIHwuR
p2k5ko1KcwVRtpyf0tTo+quTLYyGaNJA1QvJeJTyKUVWkRuC1mCy/hdl20Y6
ylx6fkaVMXMVg1HFeN6HfJ3GjzoRJSAyRCDS4Etec9eaOg6MVKzU3CPgi1gd
NcUVWLFzGC15wNwebS3yWHrgkyNtPPZfgFMtX27TjG4ZIE0uDmwKUEG2Yepo
oMDHOUSDcXMv7jWAloOyGAq6+4UOObVw1GVoH15rNcPLuftcOmFtX8PsZxua
ev5v2S2WpvvXaV814CS4KVyhkVEULO4c8grweAwEow8o2EWDuDCWHAQojMM+
juNb91FuSh2Ujzt7J+JHULqtKGp369J3nWYS+ZJLfRS/b9WLPOTbLXXshASR
meIOlTXF2DvWJXAgIGYmAiWZ2DHk0jjptx6a3xcEvR9p675WwIT0NZabhQ8A
NaKbqSrz4MFNW/hWVU/iORNOSA/VYuTtuBzX9DH6Ht54uQHw9JMF4RRvyFvy
b1Opyrw74nYfwkVULssLTszwcNM/ZjKXW/Q0T+Qvmci7MmA5/NJ51lNmDNAq
VJFtO81eHs96/4/jpNQ6ozHtu0CI2V5m2UM0pXyTdy6bsK3BQMT7dmYyWJPD
Oit98HdNVSwz45UfWTo5upIgt+PYgz/FrYwbMuwjXAS63yfquj7kMAMd+O1Q
vmGJs7HLEJWN9BHEycgUqZqKDglVE/VIe7Aw8K0LZRMNLciSV2HJ+5zRvFAl
hLfOXzTQn2Lox0uNETUHC+kyhw2sRKjms5UMZ2NvbQCANQGM/UarsTSk1V66
KfhvESwWCxtfcWL3c2Db/F53QjgEV+pBJWfdaZERWinIwfqJTGj+kNPAHAws
Fmpaol4sXE0ucnmqxssRLWgWZoq5APUPnDmJqMut5EtrCHpKVOR1uQEBBLEJ
QS9lpAgh/mxtc1SFje5U+oPeF1gO2YAu6UI4M0whwUCNzEj0Sm6YVVI7iztd
VFtStheNUJHhfT44SfHVdES9DVNk9rtshGBLDnqJBTVqvNG3qEs4dzvHMywR
/LUbgBw3EFh0Mi68tLu++EZpbmj1LZwbAgYtwKhXAA28zJvyOLxgF/WLoamW
oVL6EE3W+NtLog/RT1V3GpLPgkU/n5JlF8Uqt780Ik4QtfJIY7eXk/47YqSs
9+0lVc6D54M8M8XntPMK8SfqaVrIBaCNwMZRir+aamYiXy2yMGxK3DHghdM+
LC+5F3FNmsx4O9WMq2rEETsKK/847cLcHCwEQw0EuDsyRmLCu3aP7xbyg6ev
YCzqmQRwZW/dGoEE6PvBKSXg8XIw66RTkzijeBShuZr+YnOES1fRHZZVF4Au
/9yAPoMzdsPU5/THsbe4rWua7XD9Hmvkf9Gr5+fdMDOT7M1FqufbqalXSIAZ
lZNwEUCtDqT9Tq1zoNSsvPqkuxnQZgNhr4T2xop766dqgYZqC+k4OhjpeG89
4rcLXcT7uTs/wMCvRp7a6ZNMdC271ettey2ft6M+iDAfjYA8R2rLHUVL1NUq
uYqpaqCEqElnPbKDt4hiae1DAbvSUAGSRVXWT6+zkQPlIy1jecZioVUNABfO
yg+cxrhGXfaF3FT3xy+XYIAu037IoyI2/wQ2+5zSlrgIyBxxgl/T/P3xLFqp
ixc8ar4yttI/uZwqsLLgMcmfLfXvYzL22gHGxWl84OFjq5dcCyRlnIM7Vz6Q
cop06MhNc7Srrr7dXi8e4iijUjaq4u1RQ/PrbE2FBu3zcOyqM4yGElwj6ONc
NSql+HELCHcwno2PHAbeSL6fEvKHgKzO94oIpXztCrjIigIkHCpbSVsFrI/0
HtwNrLFfN5xRQqbtpKOa6PfG8xnnWXMJFvjtRSnvCGLtNX4NGcJKEkAt3GD8
hFHEbCOAbImeJy0JqXvnqmVw6eWu5Tu6gn0Q3wSNaOChG6IjR89lnRhDcfCc
sVJZ1hq9Sywq72ipmhjJ2c1099pfBn4iey4ZyxE8sgNRGDe4dewyZYIZ+6iV
NzBjgNqcBNlRhvSE26DjccQldkXuf/ZwOmvurtKOuKs1MwD8yK0izkPLjZ4O
pyTjSEQFnCIPSii2G+f7qLsnquQoj0SBNTlzP6XEt18OlGkpeKjFejzeuOVu
3wcIxAwQ/Co484nki5nfXbFpaXgOGNBI4hr3J/7yJb9t71squSY9zIpzfERN
EcPOhBod98oqtf/w4W/f+NPPVeuVpXRiX2sR3uSdYBXBkSNnu7fuKSEyEZkD
YVwHqiOrmDTb6DsRBjrcja9xmjAeKDKCb0ekDUD6BXSMtTwlDikmVVtgMrRq
3xUHIQYdFkTXSAl1H0KkJ9vtNqsGzIVJ1QsqBRU+RM122oBOTlzdZ7PqCsUA
yaVxyqPsIOROuIDC+YJkwawKYFbuTI5cJacQAt8nsOOC/ARYnHZDd9WPGVHp
W7es/3/KL4qHarvGiEaUO3ybdJc47Gt+8XEhoxtKQnJqSNcAiRK8y0sfu7gJ
DFidftHAbKihkhm/dX/0H05YzIyHWLgN6pgmU6cKvJkQMzXwohXjuUedv88g
KAxIg2rGkRe4vwVK51AlzvJA4+QozvWEmNEpdObuoO5Jn+K1vMUub5CbODAq
zeshgWGSjzG8Ui849/T1efKEjK3M8RegqByyhXrZ8mnFHKKmX4pA5B4e5Bdb
WiJZfVu+OUqMUj74OPAcaJb9sjKZH3dP/fI4yXUKDu3vDwYOkvWL8/sjl+Ss
n0zyC/yr//3NK/okZYeTdSV8EZkppdnan4VnfbuXfqWG8bLmIXCm8JwCteXI
s/kuoGbV8iKP72kS1HDa3NRmaUaH02qSveXfVe+z4WbuNCX0FpmAX3HV1hIb
OxRMXQkGpBr/1UOb4qI+9Q4hPhQrGvvnkYSZkKp8mJOy2cf/aKHWoyxACIil
ynJUJSP4uYCalxwBrWymj0LQm1uEEmc+iztpGdo1sAttcYxMF9YTOcL4mZGs
AQN84Q8ZwgwiFgV3qkrcA8sfCj2wvQPIpb3Ob1BtqRAUfe1zTvFDnwSosqBT
W+paIcPHB7uAAK0WrC0iPa9VOP3Ewk3WFX8X0T2+fliN8hl9yu/V4ppyrJ7n
AISmh4SschI6uTNAyXKVs1+jBAxzyFK9y0M4Rn36CerpJ84ovlJikxSvZ3j1
Mie3gsc7/JLUfLlsldvY7cNzIj1ZEOGuM3fwhg+mbnIO2qobqM7Pg3jCG/FN
B3BNhr7ZxQO8mPmpZOC8brGRkPvO5DJbUDpVpN6QxYUlSLOGKNKP7g/lA6zq
aff21CbRx1JmgkBCaqzIlTXuINAaYJmivc0Ju1/jXqICU6LI0k7ZH9rRj85c
xvZpNwZ5sBCFB7ETXxbIeY++CcCe3uQ2Hx7LCLXclshf2t8GSBdq/8i75BvS
LFqOjgDt6nh+gDbD4mtr9tc1zRlJHMXw66ewEsXayzNZyw7DIO+1HUz/4oGT
JbFXKOJ0axftZ4/dx9N7/wNbofU1aEw3x2AgmEa9JYEwYEWoDrSfa5CaFsQZ
jkmFJRUJmAJOuuNQqPA3c3SO4Np8Ylj7X1MpSsa5LbwKJXa+Y9sNa3mxEdHO
FD0I4+BYA2jL8gu6v75tym2SyH1F47rKiGM+yTjR8iUd8XOWqnvHBuhWQbPu
CZK1EWdrCdi78PCnVy3jCOltgkM9XwqLV0CIfWgueJKnvR0xILn/Jj4HlQGo
HKLArQaQpNlGpM/HiRDBYsMLzqQ3C5T4Zciylndgr/qNSn7xSRrIuFT3GGtz
RG/wiaXHSEXlXT/ycjr0P9lrN2hhOtCyqQwAMUIAlTpTqQkSKuM6XGirWRmw
yRZn9GVGjJfdmAnaKAy63D5EZvwYxE2VCRRXUG+cinII92i2c/vvO2BEdGa+
VKzDRTBSNWQ2Igvr45U8WjbZ9d/jquozei0pwmgo4IAk/+FfPjSdZ/Otle4h
zfGtTwYm6QcZI/LXhG7F7pO3rFl7mbVc4LUpFSPfatG7OqOxWdlVjRg9YYN2
9V1WTxMN/iyrSLRe+9dRp0zxT9CFNrsZ+N8QUc7PItFR9ys74MzablC8mgD+
1TKs88q7arboC3Tp4kbl80tjrszak+/juLMWcO7OUDwT3Agm41p1Mv77jEyz
yFX3+EBs06OQNrOZcMQmw5Q9kgiaeKaKTAJN7D0TF6g4o51QeQMbqne+NZuD
H/AQcr9Jz4oTaN9DFyUFLtf0qyJfVAyMLcLTE2REZHMsXAmJ8nQcbMtOwZDj
WEyLN1LISQQ/PfPKRKkp4vVbUWhOgS81GPOFK3MEiGNpA5nzVu9c+Uoq5LrI
9ddAn9LSca75l3okbyXkD/Vx5FK16AdMZCtI/ZUBeYHK+jEq1okwW34ww0yQ
WbVMD9mtWr0w5tZ1rLsSSQoZyW0Gvp66DuaRKYrFMC0FG04wDg2UPNaT6+gL
x9hcY3sMCegr+vV3jGq5A2W6iHLmHPMjeBATe78M/HMhIjiY6GvdxGJNCg6O
LdgFQYKX2z5kwP1pxlGXLdnLSRmQ+6si1rGgvC6Rp9GmfVvsGd1P3LIhgvNz
v5eKcyzIG1YYAw5qANaNXO2SVbJDh9U7f1/e/P4lrTrWwtKdkWFBxyRj28Bd
+2cyhwLsv5DsW60hVeyIIPRxZHt/dysvbtbuZKDe/ZkKiak6CZlJS5xcIOQI
hciHqYu5FWal03xmJaA9zSgjuKFxhJU0POPcdf1kdZzo24oxakClp4HLj7r6
ytivM1B/fVlGqMSBV+L+3Ni/nafQN4y2OtnuP7faE46IbRlmyN2rllUCUNav
ysddnO1asR1Eqh/vBww5vB27J585eskNpNlc31vJ0ag6gNiBeMSCN90TrDXz
BSD/UzmKRE4m5Ga1WrmxbqLlUBHajL7omwJs+LAl/BIBFr8R2Rw6KJ5o8jF6
GM4oTIe7E8tACkWkAVYvu5j8sP1gwNMU9xXigDtE+wsAhTyPyC0AOd1l7qtU
PwGy86AxAYJflz9/PNOr9b/CGrFBkmNKf9fW9Vc/TrNXFwMddr4ZBc31XC64
iDiNYgzOJiINdTnHJg3WsFj9z/T/OM530xT8kyIiThM1dF2MzAtp1XAgscP5
itWwVU7mrJFwLICJCDW3iLILDA9n/nioiocZSRwLbiJkiOs6fFzaOh0UNXYG
oeUbsp6KXf96+GfXHYj6mItCN4hJ2EweEZzBxTTDzGv6ueDQQgaSvAhn5aN9
3MLyhQEi57Syqfu1U1lx9bVwbYDyYFU4GYKzr/kIZXcVitBkyYnPMb7WBgoC
wmnyFMbOJyf7wwlm4e8jVaEBAGWZvbZYtHAB6x2pyFX7AvgzQoY0CAio/QMC
nZLcQ05M4KnWZgUOM2mwlpJu0ws8CK1knnlghyfmXZPCAyO2g8KRrBtHtJuX
anA7zWOshlb31LC0AA7s75eqz73GXP3v2srRcNs3v89XdI17Kw05VYNTofrQ
9WkWg/3ebKCclLYYTTZ0OY3IdBSoSIyLphArv5HGOm3I528VbbrM89S4n7KN
/7qJYuEc3v+ZfaAKy/rnI1bNusvayBN83zT3AUZNTmxB0xtBor4O/OFi4sBR
U+jWaE1SPl4boji93p+AWfjO2fUsN1jem5+zK7gJpynCZ8W2giISPuwX8603
nWGVccSE8QgWJ0eGbrfGDU+9glAG91jH9YG28QxHxT9pAruCdri6cNgYhGx5
HxflakLyTyTmZE1Ublvvt0HTHYvqO/c6JC1U+SkPw3lgn8bWF3BJCVyPw4VO
legSX8+pD31OBdNgVIXsjHool1C8sQEGqT/NfP5mnLNtjY6NTDiAaeL3Hark
EkvXD7ZyO1BK17iTCHHG6JTizsbTaXs8OLnOFk4gJceoQCX+aaxLoCNg8hEu
qRA3uRCvliUExu8NEBUDZQ1A5/sxC2XUKIUsT/P2t82/XMQBvm2sL9RFcZhQ
HKmdGiTGGk1NhKTaa/xH50F6D/bAhQ94hDRSXT4gOlHYKdaJNe0qEsmqwMEi
gpIb7fAuyxZLaWX10ypdw12/2YwSD5jRytJnmzBMBnqq+4hMBL2aTT+Y+wnP
USo1IbIYpgWP1+7OZT1+n0+fFx+Bpocxga+fPL512JY2bA03RSLZ8a5Nz/Sv
2bok+Iac5apUD+FVRz7RdommwQ1kEEI4ijOHzs/UlBrzaVTXPWq4OvV7NaCQ
gCTrTEh5K2HgoFoPJpoUmLBj4Af6yDiFrAoq/9bSk6qsVX/e+IMkUGLbBZN5
eHizKPwADoLrWXGPioMgXRERbmo8yGlMmTfzH6C91oyEijA0Dno40n949+6W
8MLUlrty+88OsyxGKqd34c0Zm81DalccX5Aftl4SFT9itkaiXdsO1mT+KoHD
ZjZ8XgeW5hU3WnNDZfEwLIV9RkqQD0ScwtBY6frbQv8VU4O2vB+OWbmK7fNH
cH02fb/JlETa16E9DMi4hgpO8tDGanaFfgL7yQqzUqd4xQ6jPGlegBKvwLM/
1BzfR6KQdWPXemEiAnZlIqP1deO5H+aOmriyTIQjk4ckj57rq5QMc47LEy0O
yj8epPBCta6ZMlZbOroQI6xjUPmQwagUsUV2xa4DYBF/ylAZ7aLK5z1midTm
BjFjhhM/deiyNT0EeUgCLHah+gLEbq0v2kq6gNalMCqf0ztLFQYXGzQP792P
nEkcAvydbyEFhM2E6cGLU8ScPxv6RtwCSO7U6VR1Sg0ta+QGXmhm3N7VJ1I5
+oA0S5OoE9zx7rPDt5kaz3XCpciehQBlpqSjfdkZMDs8W+gEKLn+4/X4hbIL
JI4v7ikWb5E28bp+/ZMh8h3tCHnhiuxCid41sXQtzTS9gpEKPV0tkOjEsZUu
Z71CwNxRGZeIduWEF7EdYu5QFKKrrih9LudmPrQ5qA2MHfTqW7/GecrorDWg
MTGFtB/NeFsiP5rWOY/tSFvu+XV9i70sUgtkCsXrKzLsDSQZt1G1upMy4Czl
B8SYHqYtOOCErNY5RmVDU989cJLkQUInNDkr4/MI7vrk0SOZgqf/Q2oABVgR
Z2JM6AquHokgUTXoG8hnYLO2gIuKRe89RMEJizX0x7FjYrhENJXH+n+/2t/o
WeVzgN8RM2GRFUlqAucgL5YNeWZLglIk9jVICJzVVVhFJb8NZ6EDQwfspoVy
08BMaewQauWpeauPyKVT3E4U+xtfPaRg8Nwv7k38eLNS/pPjxb2FQQZHxUt+
A4+3nV/04U27Gzoq25UXyIfZoMWcxEaLc3j+g9/uT3PPXY+EzI5xTRVMYOMb
ZKsEEC93HqFxlFTgu8u66IazuSsTbUrI4RK7Pe4o3blGdkr0Qk1mwDkvqhO3
Jh+Zygod2nzpmgJe62MRK4RS9WglAehK+V4iUssmDgpYXvpPeXNEBUHPiPN1
IbIohQ/eNd+iERKK7C27kB75ykpTL8HakNPd750oM9Tuiw9yiqQhf3IpoKF9
ufDgf4/X0kkWRZz49S1xtwpKHNx8ZHPf1/luUVikOZq+lnJUBiblKMgq22P6
RqMRW5LcoLcZxZe/lOaUHOImZKSx/aEHqaWef1yLVq4hv1nbka0ATy4+qbO2
WY+FEl26BkTHjsP0wa34S2t1fw7lSVyNoS/bXaBIragT1hVtvCvN27Y2aKPm
gG6Iw5dSh0zB2gZukAAUo1+FIDC1wpd1ecDoGnThK5aAVAIDLq2vZ5Fi97c8
g0VZeKyeEKYiB61hvZyg9GS6jly379dPNTwYQnfJZhTTLhqBpO3tJW78dflv
8g9nJF3KQ1ocaS6Moq6KwLK5kQZHenXNRoCAHNlrxShiWUqrMOk5ApxG+aM1
NsEFcyactiifCYbTwdg5QDlZsZV0tvzKQMF2x+Gt2rndJ44m6QhnINLyGR5+
40gDRGoY5q3iu3EIjKEhsYkNlIaa/ZVwsccWiKI0Zz4nd01zO4JaiOU4UtlO
n4nmAPFsplGpvJrJh5YMXp5siedZhsErQ/PFUYhVxZ1F7IhAMIxB2VaztWoi
NZcnHxlo1wpgOu/BCI7+mh2/pjEwe+ehJ5GLWaBKWB+OGYsekLCmtlBto17E
nnrsbrb64JCYn7zyxSjlklDXskGOb8sM853eUdlG0vGpyF8moL9lpJDO1xJP
FsX/pAvm45jW5y6zC4QYcSWav2jLDzrEaqVvMIZQDX+yVX+TrLIrT/hqQQ7f
sVd2emcHYOttTd2qTdOYnvhcT5YvPD6/vtyHzEuiCnq9Y1JXivYmTuptrQal
h6YDo5AcCco3cnk5/1TOyh1F/abIwloVE79hLbZI3VMm0JhlBLzjI1rHOLHM
ywly2vuho/DKNLpsf+orbYQpxdzxJ7UmH7qxX3tO07w5Z+4ua4o7NPznFG8D
4prlPNNKRAHV5deHfTpOJKAIuwlyV6JtyZ541cXnyLSOCv1xl5iY+N/3qP+0
pszYVpvbECnKwntUA5v3HcY1n+9/Mq7l/5ZmN2XwsohXPRNQZ9SPEddwPs9R
b9TvBjldMvKafAzlObhv/zYgjzNaHRMYOhjDZwgKzsQ1XC8SDdi1FwGZat0e
uhxHzkDrcne89zjcHKcwJsnUH98XGaM5a+uGIWiatdohN+QYLCCzAKmPfYa0
+K+pVhjXdZA1IGDXd3RF8jRD17hGYy/5NzXDseMnvpy4UezE9u0caLhcUWIO
lZTVBD6DHCYUeZ9sNqz2aLutjlnJBdwnC7ATohZsTV+7BD+FWuZ1u4vgdk+M
J7W7mNOWdBbXFgISQCWhWrio3xuGycAN9aoTqLdCysBN8+6ZwTSSxPxBe4aE
+Flw/1Pg+IL6Zgw2uc8fGN6yucPIwpw5j+MzyQ+J/lEFRk/66n1ZSpoLdvBO
nb8zSgfaonLyZVm51c0qzdoWquvP2nW61nZnw3yh3hpRMiR0Zd1FSlZruEmV
lS+5KqqSA9BtQ/JNPCFDTHkJI7snSqYmx0AGyngJGzjrqPYR5/KAqfX7WGvI
TTozBfE+TZYpNOBQij/NnNiyh/lxfHI+zDRiXnzTQhVh9QeE4qh8kroGT9w7
usqG5n7yFOnI4VBcpbg86cv4uwrNBOLJpzOA7TDuIwkIZj1uJeaGNVeKOsc4
rtBnFNaxbSIM4GiP+v80z/FtyF0Tl5oLdIEv9dCTbbRngx9lPq76d3fAoks5
Amn16wgrfNMlXCMgEySPafvHDa38+ZX9RjIQPRilWslz8VzN8Zi4p7fYwZG4
kZAKaw19bY3XaYOoTv2RXyQzXterhBkmunUct7i3nqZrQ2dOjSU8xIJ88S3k
tu4EEOD5dTBgYH6w74iTuUy0TFfQSwcBWCco+h7kZdG/Ti6jUgfu6pu6tftb
X9/FvUiEaqCOUVeh1ZmiISz9+2MBX7J3uct8rMYYF4lVEk2FvqJcIrFJRSvO
udTOjzh+iE1KP1RT9UaXJDK6TBLopvprT8gy+CqRBZ4qoeoT5KlnyeeLqL4X
oKOnPruK7rfODciGNsmhJvbAydlu9fVueC74vGYk0J5DkvimGrYtf8Mvjdf0
l0mqFvYgKthfIMmRyB7ivo9tmJCtZXHSdTCxYRy8lv1t1GrG/xpFuGYH9bNZ
5MH1p3zuWQx+6PfrzGmfiLPxmcL4GODmyfosv/vlL5FGzGoaYKKbergi9bjA
l13ksYYKns+vltwrCqvOWdLUzVkSRVCQb1sEjiBWRq1cXvlOpPTZgyiTdBLA
fbixlkSq5ETgvJXs6wEK3tlY+hlp4siLPsoGmpqRaxDtJBig/bt3B5mzMhOg
eYZZNiHfDqMVuWxEO2iVVbRkgNLdUHdzd94w2IN00oFXdYJb8oIqS8h5CEhO
MMpc8OlWBk/XKOChq8QgvQ2upkNAp92aXAMem8qKgR7NX1Kf1TlmxI1bP8hR
W1C/PGm7Jw4KHdjagxXif3KeuQsfIeUXe7T6WUJOzgJBzSSGXMj9tfLkVqf+
bpf4dN6aLPf7/1su1SJPzXB+unYMHiUYU++akO2ibQbUQfcuMnyUxcd8dOG4
XOrDYIaUeHwUj5AMZOSkGQsAg7bBaK4AOS7qCbhNicLPQtVs7VucpaYgJRvT
V7n4W7x3k4yXTr4MPKfHXD/OCoZbd8/zYw8V+uodk6K6kuU5zkDv7HvZz5gK
qyQg7W1sY9p98Xlu3e/DnyVhxXbX+uOou86C5zywQkl16j0x1ZNgw9BrLnCD
zTje9u/bDwIXW4a0f2TOjdKRBlzRyG/7b+IxdyGzRovBb7UMZBVtaUh2OAne
WWLJpNVPB3oKe4Y8daVzHIXsG1QT/8oM+5w0lRt3SboAMxs6hFkXoorQg1Nd
+IQKWdHKyBMtOQXX0COwE0SVUGMDWCQU5THMnR7nyo4AP2bsyflxRohBMmcN
XtEOmUIDKXOQJjxxqgNZOrvjzDSkQmZiqFbPtxtzw2Cg53l0htxTqqt77Ugp
FTGio7PHyetB6SbNlErQfb6Wvlh1OsaKtwLUW340Lrx6nsLfjGpXOuRZ1qiZ
lqX1n9u9YOKo1B66WceG3n5lAe5Utp2UVFz3cCNl7yHZ6rLvqVUR+C6FpHRJ
V0Iho+qFW/NndS8begIPX0Aa6KDHr6h8cM3m3Kwyy3M7bufDxSunaBwTzHiF
ksOT6hIcN1Sw3tJRtFQ61LAW8mG3Q/twyyDkDEgdnPNTKG51FeQbxBPXkqx9
MTfsLe+B2MwRrDy7SbifM0PaupA3t8ql1s+vxZZhC7YQwnYskkMKxsxqP5TX
MBtcdAoYVAikS4cRe7nSueMACwkklGqNqo1wHHhU7uDvUtW3csnsACyM1PWU
Z8OdNkX9iUrE0AnVSgwQZqWR3AOhiCLFc2AcFuhTY62fF/74tyKAvN6N8W2q
OlPExSx46WQqEcVsr1qE6r3bm0bXARVCIFe84wuyltCssOu1WXsHuwUaq1Ut
+xAu7b3JLAbRj1pzNSdiw1/uPBS7JLqtM3FeP3BIwnBJ22eXVeyIum4Vc7l6
lV04zeiGNd1gyFJ7UDhFHZRj1Qc8maDR8exFEgEBhfoMbZqoVRFJ0IxPyHpS
Rqx/06FAw2DgPamV+SnNtulQngM2Grb0Xcjew/+h7k4tVu3uMf9oGA5dNTnk
VOG5H5tk+JsmwKWM+7gL26BET6BUXEuH95Ndajq9Hx6JyoAXRwT3Gyc1Jojo
a+zviiIajsQSmNdM8gnm8LfewfCzyQNyytZYV+lP6nWClsYPG6nVMyE/Vum8
P9c5kZNGg3Mm3gZ3/1a/J/aQ9wPU2ZHKrVMs44Lm/G7Pn7GgOqRaTjaw6H+p
qrU4X/N9z/wmG24zYazC2rszwNjsznk/HWDR6HoXCsRMV2WUmo09F0CQWcJQ
q4GNiL1POgAmu+gr1JrgrX0faAZLnLZWp7PIg1jJv2XqO7LnOix7YgDg2pIO
K0EwKWmg3p1TXp3sbXS8fUGCTXd2cTlLspTM7mltz0PS6QznDVx2DF41awOB
xeCSqt3jqkGVDJzAYD66IRivnA/qmDRcWvY3BcKi7F73ks5U1Q/dGIehPVlq
13c9rjKRkcmg9dbFL0XWkjco9yE1tu93+wp5PEjT0HsztweCb4/xrs2yE9Ia
dC3JeIb+F0iTNsg+JDJydFyo6Po97vokC7LRRSO0ZmVAu8qT2gVLbZzWuATx
lG3BvHP3fKYoKISqyV8loKbZ8CZR2aKFM9v1Ybf1ZSCVWG6gqLRkHC5xK6vh
1VzOq79R4e072i05qYFDnjy2YH3lvEEJVA3lix1zPOPP1nJ31qRTvRRlFENh
rSMq6oZS5+3wT4qRiPhmO4/KSGzseqH9iUuNItzWj/A5sJutDnC2eynZNKrb
bHrxKMUbNgbFvpknhtUcJnFiPnaP2IqF0KjWDLXau+TITwY0zABWGnAPPu3C
oZpeCSfZg1KrTjTZysUVb93zTwhQRAqv/FZiS54qsSZq6cfe6xjkq4KW1D6I
zHmgA3NmQ8qem9LFi0K37rE/YnUBvd/jjVQEYPvcDx7awQ1R1C0PcCT28B/w
CVdoziBXgpJcgSD038aHqgq24/C8W/YRhE2HUIgedpQzD8YQhGoN3pyZMEze
cdZCHHgff4yCIjZ0Y5rfcZyEKyEyWdeXfbO6jeO25+xmh2VYwMD+xOPLXxrQ
ZwmCPwp20hphegrvtefD1EEWqV0q8DlGexjO4ZydqYOTf/pQGDSyofrKfTCx
xqPdpeVCf8T13tEwFLNSkdqLzapWUSGLjGCVP5SRCQopgVRImiOrSmV9nRVk
ejdLK4vCqBhjNbGETEh1ndarg92bdaPXC7HhHOb0UffHecvnNFgofYg3C0l9
yHxOxJyurznUhELyB765RSL5bI1eANkJEE2Q68lLgy105JnUgPqZYkTtRTx1
YN8WB/F4QtDw3N6SIRSBDbmBBb5upGCTBdVa6hfH7OHl82j2hsa8dT3RaWLU
XPa7c8XSUVH4FYmjo+jPG8pdmd5ES7b1qFp6wwu0S15Z5IE2DGGB01J/8J3p
DPJefB0VI3mYf1bl84eyJ1Z9D3qUYG+jH/uTZKImKCOQqmOtMRM8J/o56DAt
eSJPlE+CbTLo0x0UXbitOqePhPfvBWTrjg/KoKQXpLAAvk1tJzf+EwGN3X0B
DepcEvr/sJUtVNY7Wy0KP44jht09c86OGufWhzDi4EeeNyiZEaIgxltyDgjJ
+3GC2RdjyNTlB2LxvnH1Vg7U8GMl9luKHEHgkWef6FHdV+/QN4BBhiTYs+R0
Me+pTOS64KuveHkNuyscYE+sxJDYnX+JIn8WeYfA45jYfYpSDJ8aD3qOt6Wx
S4fXHZUNng5B947tc09cKkNgSS59khjPJm9eFwFl2guDoGYKz26Yf/y6EXWx
KJCrAaWvuXPj2hG+qgXz+AUs2ZCV4OF4PgL0/KXgjV/I5ZEdGdBKq+HDOkfX
2504lomCKclE9MQcXbXk6AdDuvMmeD3iG0K+bg9kZibX3e6yYJykPJPFwNOs
VjEFPXDS0T0rj11nT9+czwrnJ2vMR+vJuZzoXrfgZscl08J6ByZpei+PMdlS
nkOxnCT3ORsxzXrXwfWmac939tzXsy6MXpoxLmZEGFVwD0Mhl3JKQcR66JJS
s4fi2HDwy1ED33tsimiti1i2QMIHRZT71IbKoOrhJZNq+clJcgvkJ9f4O3Pq
IRlEakD5PqIJkVu9lUPHHce23gYCW1d+8lenE/WV2LLBjHiJ5F150PZBTO8E
VgnpV/KBhhOQKWxbXHbQR2JbQxRyldrIEfVymcCJmiziVHU/MyXQhhTMjE02
omegUzMRa20GZg6+lHvRHh/lCwD3O3/q/TiGWTVpWMfnVJfn2VE0xwoZOM5y
Ipf72EXoxuZSkCP8+YCHA5oeHU3QFeDtFXqGW9YHbb7OowIxeM3tUy0+o4Xp
CowDo5W3ffKGZb41XZMVJLyB8LxVgFrQbZeQT6MJI9GwxOlMdG1NUJ2pwsOy
M3CZFlAyK7s36jWZgVx6pON1fXenuF7io1knFzpmo0suBWN2pUqU8kNBkX1q
TZF0kJW9RLEOWLSbWjQRU40TcrZBNAmM7fi2OVrrwu8JAQjcrdRcU5X/8N80
azSHtRG/znPwF0MZ/L+FaDz4zxWl/zFUMnw5YC7ODeW8uN0m+i9upzfLYn/G
uYeIlaacU4e9a0ELQaKEzMe9+YWvB5BvsXKqR5LiS9DBsT1aAguYua0s+f0j
7642atZhOLr4LTUzuxd3gNPemJlwk6aEKzq/gficMyMhJaVolYLqcSgSPb/N
RQ60vNZejIXFWYVQocu6wdOaeCN8DrCRin4vUP8++/JuXShi7OsCpkRS60S+
22VghXapjTffzX7rk9xrpx4i3wJ6+wCuecBuvZlA/aPdv4eKoZkvBRmlucgw
IcaaZBfebK0BEt3RtHK/zQCaWfeP4WDua1YGZ8fBDPD4ncnEuvWTvSHSZ5US
gzP9sgZ/HiTJSEh8mwx/7gsCno8TIJzisRb4KxdPd5HLlERn6Om998L0iTzv
oRiHRHCEI7yam4N2FYC+RMYOfJN33Ug0Oxw9LEk7Y8Fd9qPXxCjxFXw1Uknv
pNXpD7CML7/0X2liOwpzK2GnxmWUFVCzxjXR3Lb3WOSmUbFPz2Q8oB8AWjLL
Kai0uX3uWfivmkytfOO1UPRF7bO9sSVLDA9AKgwNToVxeynPg8Rm0Q8CLRr1
79DIHgKTZ56j54ySGJwM24XaGg4FYzjhSpQEKvxjA3x/CmFUH1lH49q3IUF1
UWid9VjsB+1A4YKjPBuBN+wVtqaKUetHDyM0TJsa0X4k21go41b4WODy0j3I
7ONy67mwMW8QzsoUT5eECKxKzJKgAs3cWyKUj6D0gsATsO11TXuRFdaBhYVF
N8mfBLmIZiN4x5DrUAaXfF4KldXp6Y3XiQPmf99Dz75P++Dr79XBlOKY0dfY
B2I8rtctLLjv4kQZqJB1A0IngwTwFMk5YxP/PPCIdBSgvYTo1mHKWVQKjtT4
0Gc9efOIrXrBQHXvWO+/ChvKmtR56iBLsGGHhsP2krmR2nLJh3y+AjnwJVKu
IQzWaym3CKlhN938hkVgdh42lV4gLI6aovZdMRn1XiOn1VpHMwREbPOuj1ct
MqHjgRY9HYU2oCTLx6MOJZ2AkoGixnWllzxUR/CqcxB2vGsd5tabyPhvAEta
MFJuRpP0da3M3M4yQptmLT/qGQiAFFGipJ8Yo3f+RKsFNqlSXaSxj1otFIvC
HzcY/scdsUIlek6ur35yIeU/PSDZiN7rfulr+z36+lIWwEDYmYp8L3C3MGjr
kTYbijq7fuJMdYp7IQT1RE+7hECKjr5+ZqihoH40gA/FTyOrKHsGcaGmvEnC
SJjBSdfHdl83AjHa0gyqzifWWPK2jS1cvdCq/gkkPmAvcK/92KMcCXGOVPJN
ZeLFrMN72yCRDynY6WsHsYMLZi/v1nwjze5UZE40BNYEzEQwhruDQIl2fLuG
7WGLoO1YelMJug4PLnI1Ihjq+Zcvua03hJa8hsCFuykzQDMWg/GVwLlbP7XN
yv4GkfGRNcE9eqzXZBW3EtbttH3lz6obR0dJXWi3yaVLOqWa8dBndjMKD5r3
n1NHK6dvd5hDCUzQ3/siekRcoG/Y08OBpz/bUTlfZ6R5KHNwfiD6mMrOfk5J
K6TlduXUN0Y2aoq+/7SWnrN7H2+aOONp3JwrKMqLtcV4XLYGIKP2LHfiX2wy
ohq92TfoyU+oSESD6vqmqLoS1h3nrT3BgJwObJ7rEYoMnzvIur4ipmo8ZslG
DVgo3XOCmz3gH6BHsTnMT/OsyQp38iGteaFsNrkjhZyuT+CEcpd6i4xYJ1Rn
dZbadvcb8wFuW7nZoK/HC+dSOy9NB1+t7+FlGaB8FzRK3sK9a+9DRE0OhOvs
gKPNcCZQ8zxEO8YIvbqBHOWP2jmZOLTN9dKoupPjCqvgxllv3F2sYVHbl9HC
/uxcHJiQiEYROX7gkl3YrVkmnC79VxLEuOaSP0YyYamQidisD7quwT8YopP8
3NEauG2RovQQVDMQ0q/QQu8UdT8L7ZiafVbc3ABMXRSFKUWD4wzI3XhoNefe
FOlc9IOtkut9aDfp+dWxQF5+Ux//V/C21fOahKnqNr4W+Ju6YTq7llmJDHmB
ivt1KXB+GKFVT2yITV1ThwsL6Sl72WX7kKs6jMXV7JRysKFQ2/1erIomuaao
YMZ3dSR0KJaEEO7hw1mDix63lCnurWf4t4WU4TDWrRRHulxAE2vy0WvrnYm7
AjunWSUSibVtl2OLV9JYQgp4mgMx99JTHQ9vsJ0EWLPr0z6/5jdStxpP+Pgb
94Dg03lAUt0MgOgRm8zn51Sk+GH7oKmSiLHguR/tIyh8l2bdsM6SdbFsn2yd
LXNqRZrwleAeGm53h+h/Q4oGd5V3RhLqLCH0q3kyEP/6yhnOfyv0nSOaOaBx
Ng52bufiizfUfy1UFDR32vzkb2+0tZrFCm/UYI/uQBoA6/zNOkY4eAEYJitH
gJGftv+GLjfLvB6CWio6dlDu+IdqbcQYaJ9nwA5gecFGQ+gL91WBscqock6D
/rGjlTlGjps3aLzi+IPszgF5VX9tCBP6w4xO5/1Mj2sNk6FGZQb2fctNJrbI
ZINzlRcIi1diOXQtRwgwAsmm5iqV+bTIUz9cTNHGIxJ/3V6wFGkCLc7LBgYZ
2WGarJjHg+YvHWUD/QArNVxOO24h4spl4Wt5B7wc2CjyNSIdGwYJDjPnXmxt
Q92eNfLCC6v5optK3mOYlfAi0BJYDYAoGKwBfhd+VEATzP054aBnWlph7a/x
ZwQ3Jmlw9qitsiWiPhcmtKvp6peixWCjCHZQc6Et7pzxVa8q2rb/bDUM3C0k
QvUctD7u7xPWlrUlN6763GFbRa/iSrj0n9HmyXGI9LctWYmQy0um1NekauNR
W2/nEQW0izNvEFpXsOJUWBngSkhTAzK79sRgTu1wHEeQRsSZuBYuQHMADtee
RHlTQ5z+q03JQhr54vAJbk2YAFCERlOlaA6iGhYAvJtwO5PDTSy1eRV0kY3l
FjVnmtcgggvewMSsK5qsx9jpQCrvpn/9OWFUT0shr5X5EUW9ToFMuVB5xoBT
rtTBbPl18Q0Rob0V7vXk7pAA+oXhRr1NmJ2ZgZenUdu4wsQdmfjAyMELOACv
VHsGYb7DwojDo2YwMzNhqYnXgMrAVKSsGtpJ9RuX3vd491RWUeYMLny0ssYi
Xqv6BT42CQkIasc6wKPWtUsXsC6p9/nSXxsHm1zHGuFFoBeUhvW9+zMlj34M
flJ7lsS7UkwZCaDEFdqN3v6C33gBMmLTxhMFiz1w5Y1j6CzkYNK0Av+4K0Lr
x0sjwvxq7ZPY956z8HVpEEHaqeUrgZjakwvwZtB+VJJ07eYBsG1l/OTwC5o+
lgA/mlCuVCJcsdxOFTx97mkc1kB4Wq8hokiS8ZKc8kgTpOKXEbp7+Ev2Cc+n
3j9S3HJNsc0rW87RbgrW/gSXFR5PzzfqKGLl4SLy8uaAFq1VekVcotZCBfyr
VuXJDa52MpOJtR/I2BXpi+k2n/5R5CKcinIKtJI+zwhYs9H7S1w0RUl/uTnV
2XdY4ivenq6TCbfpDg8AlUWD5kAx5U3Mbh/m2uxOn6AlQ1HCNnYzVR9FnToz
bLVLBTOsZkFUXssLnuXP6n6AZKesEGgDko4wvzVTZTfvhcr/IRoGiE7mhUp9
x4gvPYPK0b1hP+h77quS5sZLlwmQsbb6UMNzIPnx6RLYc7AeLd0HU7SHTyAn
++fYG50WKGgBod1xY+3l/rdD06DtxPMQROivFCf6OGhzLRKkTXEaCssG4Y6d
mzp+KwzRnlzsVD624zLpn0BHslf5S9mItkYw2JwYZpQ6VeCJL7mlyvpPDYlo
o1iLPxRdpUGsi8Sn8atE9c3ERmzB47VKuPy4s7lt/cmO1tFTZa8c2yAfeCka
g8WSEMkmUNHXTECTLL9rCKzv7cVWLkzhNCAF1tYFJ7X0ooZ3HUUAKdy8RAA9
qpydjw0Re7k/MHo+NL41t6kohKaIXbyKGcpzyy8dxfxiFJFpA55MJnnPf3qK
AehrJScAEeZCJlM5PkmwJp8LsrlNUG/ICGRPDnxe+0v+Tv0R6FYuwMpvldXJ
oJgr/xD41l7ytdlj5Oz/rE/BCM4LSUxl+OBBTopUrjdEoGa/qXOG8n3r0UjZ
SSg1OCHepqLMqU3RFjD9H7NerhqKw9nOrAfIXv1FaRvDgLE6oaeYAfjvOvei
+9dHoynnAdGLjlaf3pbviGhWsAW79FqVf7NelbM1dZdDt4+gGHAG4ikZ8mm1
7/UmFzcleiyMsu75OmR/DbdCZwJhQB8kt/tcULpsGQGa+o2cNHu7d9O+rAT6
ftEPMn1DO5R7KEuirU4FBcnq96hqlOblmM/k+aR6HyLBUjvXhEtXVxz3hF2N
41nV7laXH5igyOGflBTviQMR55UALkqT6iCkNeLUrTFJ5vxFSXN+WEEN8uHD
g6oLZu6Ies4o/6WZz/PFHPJHT4YWifHUqh+fxSiZdjlifWMUINOlHFr/kJ0N
YUm8q0dGfhWwwb2+dWo8Ctg7wSe16bC0/Xi59dj2Eq+zaprSCunUmguhAnpz
El0ESlfz71bG3GFMLpmBnQhN4mejKVvHsdEi7fJyHtZ73tW4HN+pjkfIfGST
98QniwXrS4QW6eomJK7uor6HkaKGz09B8158RQKq0oMHDCfZkmDQvbyRq2mN
6PDjdLW68LF0O6xJA7MGVX0yqjyhnODGzZNF84gnssNeqU64ZdFDkz/+6qzF
MEN7ND8+soB3Hd2kyLbA0dLpEl6kGHuBOWujlExuLSrDJF+828w9jUCZDHh7
UUf1zfBaa1R9Lj9O3o5MBG+AH5cnIQL0px9/C43Q7iPXvJnwCKgoY/ZN94BH
1CRQbAq4Ww10ntmYNDsKTcTMarGgg7sqN3GqnosNE8FySE4CNtVPbMdl1ks6
q3zVmJ7itC2mMtwXjm+qiO2iSllaIVu46V7K3pXqlUl0DHT7o+ToHKqI7eNo
0SMqtF+HXFV0m5k/uFmpusnMuAsGtut3MdPJNzIfkSyf6c9utq9Dsj7C5Jwr
veeBX8tzJxauktg8kot27vE3vIxJrZX2VG/99gZGHVtZxLAg6b6ZJSuIYPVk
leDDsYqgKiQQojS8kdupGlkwW82sKuJVj3RAViJBoKp9j2FicsnHp6DHkG9n
GAUF0/I+QS55d1ozeFIA1yzx9mxjaDzCpkEJpcEEpz4qdqz3YsEm8SbhZX7c
RqF7x2BWnsAVvn+qXw6aHOToP621rOek+681oYG9Jb8Rci3sjk2M1bJCd8Kz
I4HXBqMC47Ot1YLZONzh1ImyJjXadPnfnzCyFcyyV+xkWPaxDmkOdkYi20Vg
1VyWnw7CniKvqunBihFJ84GLCBulrmBeAdcO6WD8n3CaldZfFrntmKwdJExE
e0x1z9uYmIsm1C4N6CDAh5RaCCodPevxVviSWYgEbai3DX1oji6MUycYlX5G
X+v+/r3P9xCqVdl3GEv8QAwO4Hj8c30rvtAcHCxbVsLY7qZ5yOxn8WvQym0k
zUytWhJQ9feyKQjBLgC0BFi7d+72Hud7rADndz6iallRMBq9CARYR5dWqoRa
M0/sCZb9NPRjgDk5kIH78xpcOEghoX+5RLykc5B3wSjtdJWNlw9CMlbVIadh
RECMA1L2TjW7xZ1TQtnnU5LxcqvPYfoJzkQLPVwiDS9JFTgwFNtfwjqhL0Hf
c5PW4llF+Ov5VhqVrXSV6WMpm++W35wy5pMZ136Igiw8bkDX5RM+TCZDvjRm
tZ7kZ8oNAd8tsfAy5t1WieXsvn6MOVYCc3lOrfQN6lnDUaMZ+bgyHgkbbpic
6W6+gDsRJm8oX4r2UcfN5raw00pH8x0QS4PFNEoKcxPEcGG/k/1vnqHLgMRc
zJPGqzxYt58oNCQ1BKYgqXbsBbhVLLT7Y9nsDICtNArGetV8yZlrCm9EvTgd
sZ1PcaWtG8Cm6UitqgCqvLT+MtBVetYAtn+iV+pB0Kfshd035FbnrR62ZhjB
f4chaHcesl1Vpj7JxoJvH5jE7IAs0D69ypkxUD+S6bK26vi1OJGWsWSewn3j
Mllh4SFTGNQSwmmeOT6cyufOBHNfQY+E8SSqAG1waM2IjSqffmUk9clgWUaE
6F4MomTWYTwGdR6qurops+trOu1SM5v4uOWOQhXGqiweOUWdAcxr9q++Qsnw
wp2Awrn8Iolb/ssjEo5jNT91/b/Ezz1PC4yy68Fjz5w49o8fzx7abEAgR5pS
pgAecJ+zW34xhS5BPhhE+fcaXERPqzdRZsP7Gn+d+/HCw13qQgTvHHrsAtgD
E8tQJFVI7Bba5cB9oCSp/spXznOXhDhT1eT+RvTHZlR3sV/9qs8R2snzoOOA
LN/paUpINs1493ku/LlWOMNCoeofJAUd2kruvE8oQwJdb1MBFLXluqYRnQP0
aWL/Nd4WsJ6Y0BiHswoL4jUyofDLQ+DppDjPLz03PiaQg9EB2592HWi9bmNW
CQQnVV+hKh1jJNSOzwvk3eBop6aH+pzx7Td2v6uPgnR0yjfqoQRzlFKoCvwf
XX06ETwHc77S/FxeF7DXHy5gNQtbUiXF8WBZiqsCZHlijpANfC1PwO2sq5Ts
Lh90qCP1E3LQxoi1/Zkjmb5I0RqzZy/16cn137qCLUMWv8Dzcv8WL+ExaMEk
rFWo8v6QrsOUCs58lVbruyISdSTXkLr5h2jQgnHcdHcsky2/bz0mjgYMLiKk
ex8EwxagJ0QNn5i4tDy1w8hpwjavuAZHAc0yl9noxEKvKkXRARVF/vXvwonz
69zEG637v4zOzxCzsFFzHvEZ8xk2QiyqasDGhfMwhGpPO+7U1YpAT9yzKv9V
JLL2mBSaTipT9M9fMkTtFJRDoZAKmAc2Forg/ZgQiY0Jh8BqEzIYoYy//1Ii
iFyymcGVKEfbxqLV4yQQp7jPNCyL/QDpB38Eeq0dyVYs0KpceXDL8epdMxY6
oNtuWj4qMgFyfYkdRToEi9MJsV9OUnE/IWvGHqrtG5ZqwkOIb3tpeWXcMP3t
cLX0w6ZMRprEfDsHVbIoC2OTCwFmeyP0O8O0oNVyo+mqoTBmCSQgQOs60+tz
xzjnMPBgOmhrSyW+wdVs4rXIHJXyMD8qvyXDw2AcK2/dIk8vd/XWyIe8VU99
3bfihe+Ezj/4e161I5hDZtog+ZCO+T8Y4SheussdzqVJ+Y55fpkP/tPg62aO
7sGJPfL/hZG0WNLH/HNqttFVNhm+RXlovbOIxhTch2lQeZ6b/bNjsmmzbXpt
5QtbPy0YaZiWaAWKj/7/3+HWOBBKoJylRSbuHtD/BemAPFu/ORU+uLNcl3qD
S2jmlk8IxCi9IDzhZGooRpV2eYvRe7UlINQRz3D3QoA/fXKUEj+hCJmdy5zm
YwwjszNcwlm3yZ7ogh+r7uw3SCSn/Mf4Z5+viq9j67gajB1PdNQclcMTuXF5
JI++bON8exuapqkMP3nyzX6HJcZT6NTsiyicu8nk8kxsvEUF9jBOr+svu2c0
rMRaAL3yF9O9f9cM7iX+9HODF3JGTBTSH40FFJzF9q4XDsMGzt05rKbLAS/y
eZfZzDEEvf39uBzc+ZYDqbVhK/HtF5BKUIkPSEk7au0K+TqkW8AXv1P2AViR
L1sox7iBgXSmar8NIoFz7OgMu+nxF7nvqNJcHcjqDFKGz+4tGKJJwB2rSzL7
BgYsXe54VKMxbkM3Al93aYAyPbr/mM/5GlbB3JpNBcuazO4t4gtxg//iAWw5
pvUymvzQentsxB8EiX/32KXw70axzPopd/cBapn4Vx5WbDm0rYYGQOk/8WFa
u/rCL9tX0t2frUy+9G6hFPLkym6z+kSkt3hHc6u0Nfzp0D5wLHWWT2h/zqvT
mVcXp0a042Rg87FkzDE4PyK9wKPUNvHB1Yp6vUZSbUxeTNQY4p+eVwklUs3p
6jK+62IJwfeykkZ1cVoosYuSjlbgFAno4Chg1EBprqzGX5A/a1SQ70kPepwD
+reheXy9sOhbeVqdfoOnteLEB9Fu5qWejjUDVGP54pj+U5DTVgVQ7DZuYJ3p
uwR2QC8GY4o95rrQtZnaauS4jtA63q7qKS9kKyExdHzehWoZ4z4W5f7U04Mw
QR5R8UVb2Ih9I0egqMRXPF9oRc9JtohYLeorMaRXk40wXgR6l8KcuS/Tj2KZ
31Yy+oYaqwd+XxJ4TiQx7kbVEBjb3vRoJAx+u4ChFpAOKh/beQrho1sFOXJH
uYJsAeUvWekYyHQ5q1toD4TufxNqneEa3iFhSLSkrrIKmrew7PY97VMYsAnD
vUGPYe0kBafYrJIkOI2/17qgOqgF26yMkJ5SBEhN+dN0gEVKKpvR4iiwf5na
TDWGMCDdCO7E2zHb3kIoN3CPa6wY9l3padzhOiv+ZeaPOt04JfOLnM9w9799
2IHGTV+bN+rV9VTQUSmSpSeLpcnoARdC1EVhasIjOi5ZeaXG6IurhEv04aEF
qMVzCH50fnbxKLGxpkQJhySDHLXVFdyLxvWyXtdTTLPPvT3QxjoQjaPWxqyZ
bx9vR0iFKF11uLQSKtbKCjbXD/ah+8k2yD4+QBTLrZelI5mHjB99n63NJCGK
2XHCvEQVAP7LKmCjiebRvMfsWxwPlTHOv8ZWbRhxI0j1mYtFwObujE7J8G2V
jW4oDo8i7VfjmhAovw5z4wIKdTNrZa+S7vfEraabb3Yx5njgtBMi5Pc5Wjsz
O3nFBRbWRPnllsYy4KdSYKg4CwkUL6Ebw5uf+3MPnmuy1+YC7nQ0VJszIDKL
oQMtmYUHbfIDvBs0CbhDnmjewxAhWz1tk+tzn4NMxA5TBQMwC9D300w9+pwH
HVZ6WO46x+ZyDl9kBUjkRvt5pz0S64O2lzjcx2QOpGQoExSFPYTmBr70fW9V
dwp5lm7zr/HhxWxFys6eElCXH7sgHoD3hF4hoXZzd+wmNu0VJ+7AL8NeBrWB
MZ7rWk0LGgY8SHh+eLmKRE1MGtHvtE17kHSJjlwHss6ZXYl8+893vGH8Uowt
s6dW2/ket3dEUQY1yrJdzUATYyInjnIG/LKsufpApFF7XXpjuwTeuy2jHZvj
zEUdbwdYTOuRKpYpwa0orVcWPmd6y0vdyQvl0MADfdTaaNQlk7ydqF689Moi
0jY201UJQ/e1MHgUlEj7bpBFdAcveVFxXXfUO4O0G0Zk+pXf/VVYBJenC+A3
2CfKFvwJgDAjY4xuZNUCF2db0k/4VWqZU4eJd+KxqyrS0LfbzQjA0gDjXpkh
NvhsZ47CeEvdGxlr17ZUL4kHInDGPN8YVAEhg8ccO0cYCP616Pn7n/Krb+uT
v5gzOo10nUusLHW15oIrDjBMmp/3HUy1/9T2d8Oqr6UCtyK0mMFAfOHPQT9d
3QBaIdn9K7saBayWUczFlWEnOSuM6NpESDCtcciu6Luji18dwMjryCOqir3O
yz5Z2VvjjVIUZWtEF9BH3YR0JjsciIF8yyiAvTCFgOFDbziplhqyekRc1vo3
GO6w4UpUKPMT+ulS3MBgWfExRpGTSWiYh28yEip/kMKzCpP3sbZJ+Vadr6vu
9E0KcFNTsJN+2sObshMYnvIaBnF6IZ/rZMqpig4a0KLVCbdjRpXAe4iIrCuU
spc1NxQ0n8N64dlYudkbqqC4TxwS0I9nNNFAtjE2gRxyDT9OHKQMIUEJaOJJ
2ImmQvd8z1DnlPZrafSew0btDdQFbcyU+HgButbtlBnuqiXVsepyOrP8VUbO
s9nrCl3I74tii2UNs8bIBnbS27vAHlv/OtMwA+RQ5F/45eOjv5zXZosI0Nb9
pOM2PuHGkplZnlqd2yZ9wsE1ei21a5lS5+4A1yzvvKjWgQVGLiicLRe9fMDi
5CmakovBO5r0U+XGlbEftxzUIocEi8qUGKmrJ/cw5GsOUTzwhF2MW0s4oDBC
Hjmq3ssF+7H+Jb3kUI4BMf/g2maILdUhdzpipERVouM/KEUiXbO7h3c+MrI7
ejzdw935SIxAF/l86+l2GSj8j24XNXkdYEw+qsJt0SmqzU/Wb+nSvy7bX2Ww
yWd8MRr9Wye1CyF057znX90W+IXHVR1grAqBbybLRYmNCiXeJrKv1Ek57U+g
4KDmvWF8fsu3VHRPlLsMZAnVNdszKU3Yf2ROUthRvei38tinvq+0Sc3of05z
9Od/VaTPIMV3n7UVf8Ixi7O9fKglxn0+lJGmw/14ahudmujVbPhmAoBShPiQ
qdBfnvmCr/1abBhVO+PyaWn1HK6eOZ6DwqGAZts2rXcSv4Cl42KKGGpsiUZL
KvGvrlS+iVOPkGzM+oWfbXMuqeYth5k+GRRrVkg/RxkHcXGdELPC369SkAe0
2AMGZgQda1WACy06vr9F3C/xDf4/TsXzu2QcUovRzN/ps/kzoUouFF+IqUoE
w98NbtnszduoxEN4rXfASVUzG4V70QmqRsW6K2gxZ7E1Nz+wtMZThTn3HjaC
RIl0BnQrlDmhWtCLxMhrrgCWLVLcgF8QIGAUiFKG8DHoKcqJewlCNFl6SBZ3
EiqhU8VUX6r0zf8tpixcFnbrZRk+kwCg5G1xERpG0TkiYWA7F9ftmFdWrHr/
FPzK63JuOZ4dQEzssSouDWd6ERFWFP1OQW0mzbYRp0aB2awy7pjrGmiZ5R8e
Vm0ise0ZmqEaksmntKDBEbQfeG+SATHOPQ3/WlY/hgRkPnH/5SX1HbnZhGOS
BG2/DckIkHDAXdYflGHiGc6Q/E+QoZcig4tIA8UDLho1YLga6lQw4Lr/b0BP
T4eJDSxD7Fzy8CfqKtZNUuzw6NmB1AgGba+Y6opOznTPe00gILkP5ZpfOeCn
w2SW4EzU+txP9omuj0BFBVoaZcFAYqve9EvU7aIh4qnI7fX+0ZwEJEI3t1XO
c+gY+NenR0apv3vUawlUvfZPG9CuwgCVBtwUifWB2dj3p1eIKCuy6UvxUy7i
UJvO1RHRJQ324ZXHxWgfpYTj35dvmOfjx4VaT1+lzeZz63sVT7h9kfTbhQYB
kipo5G/fDfUlDU9mnIMpZLxlrLy7woeMZuLo4pLBWhcMlH2orUbdVuuTx+g6
+aIbm5gYuAccK3ck5/20gz77MkxMxlNXbryA7+BHfrYNKtyONGgVRkDgRVKC
mbB+amvd/5MxfTGiCz67pCoBG/+WIES8huyPLborqoa3LsQZMLu8f6jRijYe
5Igc2r4bwGqhf1FBnHD60CgALZrUt7Sj/n/QfkMyZDZr/M4CbBFdtoCdJ6+l
opFktPfGLuTSkEJTXzK1Ifxt0zPuenH5FmSRqcPFPZ/kVpeZZZy1NDMMhUo4
T8WyHLjCOU3z+rT7yvJeifGJ2EnbbMrIjlv90t9L/AbriMntSnVoJib959yj
edcnlFeVAYoMzGzrV0zTemAmLKACeAfwnFpUMjn4K6BllwrJ1GnvtZZWw9eb
vInL8QKJBu5Tdqw6IOply4yeKvyFMHEdaCslVaaWBqdxLdxK/hJarofR57OA
Ng63f9VDl/tMZue103IWxbhFJOw+9sGV55xemtQfAG5IRNLR+kVNRLsBLXYo
iQ9ooJrfwlZ9eKBXDp/smAfiWdMvTuaRgE8ADw1/or3r8opkTW6pQ+lvNpok
f2OoB4wkYbyVr7AsnWTJcxmmyLGi5Yq6PhhF2y0lzyFgIqgMysL/AuJNBQaX
ADqw1Qxv7Wse4xth+Yn6rivvIc0ap8uG4RlnaWFi6VRM94KGVCE4AeryLG4w
tpv736lHtIQXjn7rVn/7a+hNc19fVz7D83R1z9HA2O9YrtMgbVfSqL/EjB4A
ng3DCuCPN8l3QipW6SxlxeD1RRGFa0eWQKGaFKHdGoI/xuyEvMG2diNWqC3B
Ls10zEkr/WRDWHxeuUAFEdNMHlbca5QUy5SZ2Cr5p/TsrxK/L+MdrX7p8CNS
4uZK8z8qdYVT8/5OkQMFlNFIXhE0luL4HlU6NjDxkRvupuNl+rOGbJrTc8oU
6MawXxaWnO50udazJ2n3pd9kfCOl+M/MCR66G7aPLQKBx8/n9ZJshi6oCmLE
BoXZo0Q41hFJjV/wv8P1bWb5+NjTfhaXVg+ihhZVNZaNk8pW4THMHLs9F/py
9xKGn0X92rOrpW9xLIaRi8ATVVSkZDedTemkYHTEz/975aNhoziPiYGsvG8x
JYPoPr9K6TaqaYxHCoTVCqy2iW6L584P71zv/aC/CVzP1qhRPn2FwqFP9m6b
CFfsGNVFRt2OGx6ZupFlqAcYx9TGlBIyKsAbJ3Z1iMVCBaHgDTaR6pSlyZT+
PuUbysgn2O0ClxLQ578ZcynqZxXd0UPi8iy8U25FOa8q1ItLKlvXpgshiHtT
4aTXzHpxTMyK5Ke7RloQ/7UsHDlgOyw3AAXQiZ6s2ej43vKRQrgrzsWBcugF
z22Ht96ZQVyuZDve2GEFbrHz5Qozd6thmJ/nf3QyBEqPziIiYlHEui6xep1/
vybt2FfDvMAHM4dEcLLq5ePQa0GmNaVoh6F8QiyNBPzqMBMT/gJ/wCrcvGPw
54JzeqKxfK2UXZm0E5NmvVgM2YFrSF0UUN+sb+hmirNW2HqiUYUd0aN3JkMU
hRirIhmFUOGWaVCgKBBrITR8FRGWPwChRh5sxXk8OFRi4h6IkpJRP2ftm7v0
nuT5LxmPBogLRHR6xCpFB5CIdOe3sra5aUdNU1rt0DimzfhkyTWYjcwtpk/e
hH2d0yqpDXKSsbfkerl9bEFh+XrcGs2mFjjBsU4VMkhv8heGvISVgjuaPODa
yIaWlriKBPOcPsZJlMC8WjyNjqk7tzTRLDFbhglwFRm3xEYGsboTbYCyBDZW
/bfGnfaf2LZGb0FaHPkAysofZZN0C5PT1tEyBC2RxSZhTbr2Cc2D4U84f2u7
O/BAdVywXaYI/2h5cSRQZ9AQ/o27QAeU/bXs2AsyfimCWqbksRAj8j/22Dpi
0pnwFqcQfZaVIhmobtoUT14C5TbRcdmZdd+w52YmgSXv/SaeCSZTYOodiou8
8ER+X6dK7JvqPnKqGFbUZkiAu2dyx3AZIm3srJC7OWIhCwCI1yqUcw3uul/s
1Gv04ubfxdIruiEUJkYtgDJGCZr9/7OzsfvbEyhBRPx2JAbAI+Hk8fkglX4O
Vx5/DXZ8kCmIEy3KgTTVRqpjjNO4auSC17vS3wT2nWMS1Mwe/FaVkrT3f4br
t/Y+29ELUdNiO8GDH9FVNqj9oTLBdMFCcXnjHp5Pp1Gur7LKAA5f/fAF22Pv
mv8uus7fHuKLBzw9HTh5lOeUcI1/nhJMcCBO9atHELITb7IJPA8y21tiub04
YUNdJ3OwfcXtAQaLbLEvFnXTrx6ClDB8tWnSix4KP5jD/fMrl3veCqoOSXjb
sezRt3THoNWZoWNiJBNlyQ12FMiGS3d62izOKvuPZZaD2lrztSzAB/clh88m
S3bFQu3g9ONHmRmioYxmUuYxCNTISYSfxsljgQiYAD5Se4ISGIhhs0o/Tm8H
dbaWocADyrYTO6zkPLrn6jUNHoK+CwGTT2R6YNUM/PAF6NkDCG9U5ylPulUt
XTXF5dJ033WPXeU21XPkSagew09iiLhm3Z50GVQeoVEprNjQU1qM/U2yxsVz
MnDtWRQs8wFr+P4I/zda6sffh3GV0GsZkF2fCIESTP1ER7turtelE0REsOYS
3F/E1Kr1nBJUQ1U775XcluDfgkCGUfXaFR0/L1aYgSPTblv2xgYd9nLui7ft
9hm3Tp9Y6rcthCkQgCJuh7iWDbxomFOwiT1IXoeifNw3XwpvuLlmyVzdnWVB
p9co3I8BAsz9jbME3uSLuhywYB4gJiPA69g8dHqkjMp1QBT2AtM/N8/QaSbV
5Agr3YB/z1uIRe3D26wvDXwFFaXf9+8HXA7kX/ZC6Y0KFHfLP1AViQoUht+s
9klKMP3+rqnYBMoCXIYYSDkS08ViOKblN7+SeFQMB95grkcBtmcAC0tldJ5X
H1H/xpAy/aI1/FXWXQhPS6+rmVUX8pEV9uo8bi8yTQvyyMuh1fNO9G0IEb6/
kap99JAg9+l+5tLF0gp/ueJnKIklzI27YmnYDKAASMPtQll44QPmPFvvt6di
LoKN+4yRLepqyk/x5S63S7RHWboc3H86zctEqJSKNvoKGDQ7Dxr88lRyfCZo
Omlvf3cdaiCe72/gi2RuyTIqBMxP3qLrrdjb8oxrh1BbknngQVxttnMU6iZG
RJVAsxe/rOBc5eVo6tahY3+mZkruCVv2cRicp3xn4M9wF5fAnOFB0k085s2b
6IpZd0gA+cR+LobgOmag0OmBplVDa1P4fyW0hDPh1UjB2YGd+PJMbuoUYLbt
qMJFGInL5ThUjCYtloi6eW466xZIDtNiOrRmC3hMrAph+duNUTNRH+76X/6f
VZTFcXe6XlmxWiWJz4PQYCLTb2en3m0qfDez/MRZqZf8T+ycLjA3aOXb/m6I
erKDx9TN5fnnBE6RToWBAnLOJu8lvaC2Gu1YckpKgasPp/u4YooKAjtRBbjh
5/5cT9ZbosTKWWHL83MixxU1ZYCREhI/NMjKg7ypcqsaK1v6KpPh0T10wyMp
E3tBd8ULGbb4/Z3Pd1fyh2gTGu0ofS9jooIdrzzj2NzWvtFmRkabRYRGe5y1
Q8jex0nc5HKXtKeY/OWYzRTNPZ7XrzMAtWPBl1nFttd+zBVPYs2y5xQMT+kk
mos6wsKQY6+Lar7iHG9v534xPHuylYwMdGXAjCauhE8pDLZCa5PR7/z1fowG
AHIJnyiYTHXKkOBjmwnXenty0IHm4KxCAwKC5EkeAOzX/NqZ+akHcJc0hTwy
3hnMrJmwXSvPshbV6Am8SjLUrFmmUBzLi4O+Wv9gO8YzNipDBKagbs68Mx8L
ycXfh3i3nlP0oqvy1BMzY1xrrCF4ARzixtVUe4YAoVmqkyTzSFhGhItoBuLh
LCmVIQpFqLhkFU2s7WPFUq+qamGmaQbwyvVAUKmycyI5y+reg1ZsYq/inckO
f+Sj1Wm4UL//quFK54BfTOeW6UGOJ2P4stA7nawQ4xfWd3tgn7ZE8zPkUokv
1y9j6U81DMsj0wJWYN/mWz8HSIw1fbJoWpWtMKAZxI6mDQ745bYMyYCYTQmf
W87SsKr+CMnF5ctqV//g1Xt8+KjJpEN+wIaPSMs6bcZv2w48VsSRhVbbRxSn
2W8xfVbBoi2lzTlj2z5EVRCILqDnLJNN4HJTKIell+U6oCLxvl9NEgiv3NlA
wVDNMPU32X/V1+UFz1sdpRweSdpSby6iNFkyiX8dYctENVISdMMqRv2TWqc8
0JAzSsmM3R2IVQzPJSYlbA4YhP9bNQleHT7DFOtk2NBLXeiKXJ8XV/CAXfFk
eL7KDofxnuEi0RORKYHZ6GykgmjcEvkqN5wnoF4sRW6nPRzuXncsaXP/aCA4
LiHPiArGPwoQRbp5SAjAO+mvQYJIwrhrUOzCB1QPn7W56rZWk3Hxe8GPq0JI
ss4U6tW3d96homodVz4a4sAnUys13xW5ncgY0m4LGBFn9o0+t86YVLl8d4xU
sHcWtzwvFmn6TnDRgIaMsQdWygrLL0UVTv+NSlkOgHwuMYYmL8V9PF2mZVQs
uIzto2GFc8jELqO2es9rIVslpoEG5820JblEt80vmAidWzf/Jiq2F6YSi71m
VDhDIBsCCiT7zRtWdZS6HBmQt/J5XUHpbTSmqQUeoEOTORpdxrwLwGKMvjox
0UJdXBLG41QewHlLNBZxgA8bRFsjJoK3tuzHgY2IGtsMkMZk83CxL2nEulbX
CaD3EQnQTV3GTz/6h9USfsvJQ2mMdKROLqG5O+pBlsHSWA2iqZYndHrxM3gJ
TAHJyy+Qv2EbnAVeBQ8au3dntr++iqcy4+B1GWZYcVooDQ+IqTewaCTZxp0Y
FWNS6p9AoYR5VYAqA2CjeCQRUzCKcHMZCdDIC7/qK6dL3rSKImLAT19fVume
MwYy8Zu9u35HxskDqK+iE+QI3UYh6tDrBgHKBeNAYMCO7XcYbfNKlyW0GRJ0
r4X6H6v+AtxzG9s9yym9Qj8Fm80em+8FB2FzWpKDkFT0d33XgGsbjup1vFQs
Uh8mGQRyWCrpAWAEhFabpCDPHGvO1FC/EKRWItyWOYnNQh+8SxcDAT/MZM9l
gkzJQAFdhNc0QTVqa1q4iDyYpRc1S+rZrZm6L+T/UGb93xVfFynlb02odrn3
GYYHIldFFx1sGmm/GcAwS2Di9NRO4zRf3Si9UMhPuG6A0+nY17j91jJXXdGD
S3No+H/yfOFS2Buz3ImTYw51uZbTkVX8dwAxNoxw36ngpUNIHzqGpu0IfkLo
vREwr0g2J7+t0O531T9zUeKv3gLopdiAZXRlEZyD5rfSA14IB4QV8L8pIcMv
GoA1ldkNyjoQf41vx8eMPBbG+vyOhvwgLTnMEhmmGAsjiHrj2wQ+sfY/SoOM
M+rH2ZUE6+k2VgGzNXkroBj2kVe0kf2iZX5hhriOm/krWrOefe4h8rngpWZC
1nRP9t/VudcpvwLZCiitnkaCnBegD65NycjI3jmUPFjvvy2gyPts7dVc9UHo
kQfrXzBaOo67Xqy6d15ZXyYwSCniQfUkwWs8KBxBB9VwYg+3rZK7sQvimTz+
DKJCqHdcPiFEmWi69nRoYesoBqqGbsTWflGnAcqPxaZUnX7hcK8jdRhhUCGC
LBOiCbGc1fkVeQWJrT5g9pjRlwOUKMROo9jCg7DHuQjPcluOXyH8g2UJrSAB
/7dA5hfyTbxyX0BATPRPv+d/lbVfeIAUq3vCy5+r/SOqWxFXsF8vxOkfALT8
bkj3S6xo3RjJJdpbZLqZ2ZBed9HqjBXltF9okH7iW3sZK7FZCOmqSZfe7gVI
vBe7iuOrJK0S+U6LlDzHEcsRsf0YgvmcJkFGHzag60HFk5Tma78QOk85Gc2/
VVSgjK8kGPk/0F3x7x07Wa+d5FFv4NdnhNGJ0is1Nn3E4WXM09Zhbq3Iah0P
LLa9SXnfLQnaXfj8hU16MK5xhRtNcs5DZHBe+zP4FgMs1ebjNUcJq9G7W7FY
iH9F9F7TThttfJm/I6dvtwVFoL24RNNF9uZk0j8C3XTN4SWspomlEcrbxBL8
zgbbEpXlwKl6bjkdMbJ38fif3+fFnReEpnEG+2D6YnMO+VzWgbotHhHyHjT8
k3QuhOSlWimiojobv74PPETSuzdWogaUI6YnE62jnZDghMLe+ysXovDD8MOI
u3Yk6mw82dT9eK/ncfBfTvDpc0UnyQTZNxXxz/hVi14KPKykVUMTCy2uQDsv
neintm7P1uyBhdc+aebJx6uBdi6hAs43d0+pJ4BJo7Bwgoo9Sofg91HyFZ4S
IhorDF2P/+1uqp1Bph7/eRbzr+KY7/pCXB6kvY5DTmnxUToeyLNEXk/6CgeB
jaHHCnmADBZ4OX+ovL8+RSbZDASKg3/Qvd/KPaYkAiVlpkcNCYe+uSQdI31X
uhz6/GXe8gRgwway2EkIEMSLGiKdfeYR6P0Dg76FjJl2HwHBfje7U/QFj/ja
0chBmq9rMzrPNfZ1Sv8Zq6tAN+sjOOdmOrpB5MjLaM6cvNh0gO2q67BiyLky
0nWyghtG8KF3KAqHfknZC7G1YP1ztn96bZe+jmjE8x/6vLj8DYxh6SpmiK4q
/LAJyQB5o6oOAypC6TeNB0YYb14+6VP1aURR98GZstJ/hjI52JIFRxGs4amP
JYZWyc9Z3olf/1gVhpt+7mmZ8b3abq6N06loUxqPskBPk362ukJPvEjpXla4
zoamp+X+L4isdyv+8yP2gEMIQ+RiturkH0yzUKUTp7R7vNz+4FprhpnPsPgK
fZ3aVW/yyrWT3jZWq1bzSorYHUOY0zNnr7JDie6JR/S9rSssqMSYTn+hyr9h
48UpkImLhianIOHEz+oSE2EdNeuDvpgHpZc4zCxasCkP58ixuS+ie8vbztVC
bMgC8NpRsrBDVLBu84Bnl0EF71clGNOihjk7PKoG1vmwvyy6LEMq3qEcnuc3
VFwHJ8HMzT7sDMzmSi2RpANRzgbXa88Hw68cXAh4EdCb09fXwjdhaqM77lKW
0hySCQ6CrgQkaoXnlcyVEdDYrdbdyayx8Tv2bpQbmmXvH+TdsFTVMS54KT76
YB1Gsl6Y/F1nZ+hJ2bcfgtLabZDIU7uskt+vF/zgDPSQ00/4ghxU64JVieXD
xGbpDieM0Cz86TNbREIlKsqojrr91wrOl9FyE60D0yJHDnPBj84rYUz1Ddus
va6SkD8S2eAP27X+eeWIFoi5Dx2JcCXbpioTNf1sf2CPLOc3ZThkS2iSkAXN
IAwTUJOfa0lmAi8ggDhY2zYoMEBX17eZuEwZvmAv0W0QRz162G7ZPGfbXTDk
jfsIe+RvsqlJll2jc1/qJNuQ4Q69DNRFlhIO/La8AQlVEVIt6wMlLlSZiGCn
9/I80dYkl69oKyqFdWa2W3Pcn+TTrFM3DZzs5Zb2OUZB/rptjqdRuSLlFUjy
11nhJ2BzRbDqZxvMg7si0p0TLw1dE1prjKuJROaczZ9u4jXqvigjyxgalTCE
8Uxt6mxb8QfyZgbB8JR7NHSEM4/F62F4eTU1eI0Jbytk26jnKv7lNSeQ48jb
bpjI69uHLRlfLFvvxPd6C7hbfUSreE0V7zbYIONZkvT4ivJNOJ/H5kS3NJ1U
ZodkOYjlfv1lihSlWgsR9adydo25KfaqdZguNqj/jwwaEMoESqR7jEPctj9U
5cvyQpMKSxt9bdw4qCeHQ5IXhIFHh0AmK6MypO/Av3M1pZeiuoP5Gted+PHN
IHpToI7gH9YmQ8keBmw8IQ37E1qaqgXoS5ZHWOrkoNVJepfknDa8v7buBoz7
Q25GxuCVz6eYJy076z6CLA6xUYnrGvDBWe5AmdZFrsfn5qbU45jZH3nAqfez
k2ozqzHcmNuDMSVF9j5W0UbLbVd2iXNJKOZUrSmVo+flW2t30VJgY/HwDtzg
WHD/Mt0QEtdRaY3DHdS8HOml9AuABOf4XRZW2nP8YN6Y+w68gDOoI2IXbrgL
d1Ga5Vm8DHC8No/og/uP/DGtdS73bruTx5Rn7pRhEx2pB4ddBC0rBKKZSkqq
4a5cAPsTRCRXB/hb3QxihuaYzmKrGD2AvH1DCDVpm5L1hfSq/5RCOodeo29P
WxiANXkheC6xvGYQDBBroeM51mfnA1a6kQSZifeWcmv1BlhhbnPpj2iQkH1O
AtoUPMsdDruLka+iHT/VK5S1NsDC7YOzqIm2VkbT+H8VPLxvXdyOK98+EOwX
dew3qXURUBGSlCy+DkdKd1fpeoulaIlR6fBpmB1IH4GKhv6qluUOt6Pep1tM
dAiz2b3++9f28bz+wKIYnmGw3LBHt3s3q24Mlq/aKaFHD8/rDlwewH2TyO/C
2P8MHHZfZMSzv5GIfL+CYOA02uvTxBikSUp+096jji5WjJV0tbLYxFJDZRSv
FyhK6nPjy31Lu8igswOP9SpxuUUGLSsWc+azqkwr98QCo8prXgbfFyM2otHc
aKMvaOUnZKI8jO5c4e2oEjwtPv2I4QxbZKArbdnnKJkMqdDswC1JsmtcAql3
UUl0XRdpKFR6XM98odnrQM2mOOUS+w6r+fSUTozDm+yjuN7RG0PpQ2BJ0p0+
jVSDsJLhXTIBsD2MwbuC6FxT/U1tRJgmkC7M3eI+Tcto8+pwj2wDNsmk1xt+
wusyYetRpqpVlE8nTzlbEFWnCP0eCK5UxbFN6EUUvlIhYHtoFBoWvR16SSw0
DQNXqfZkmYzFrvaXKnMZEQPyULOjvC1yRnkR4KhOCJUNGR8EABFNWxzRL70L
uvnEuSTDjhM/Y195zn3HwfR3yR18hz9Nif2lUqXCnwmWK6fJhjogF/tjANPb
042TFVFiF5SdLBXqZeJQMDWMWU1AOgrr7oGc/Ncyl4nrqaQ7QLonTR9/1AzY
Dz6Q+1RfZxv6xsSj0eRq3vPW3FtSCefaLP9g7hvGlYGzNgfm1nBnHJzbKFU4
HayBWNBLXzO18ANcNmFlHEJh8jatOPHMSpDcNvFXDd81qlAHjy9PnN060WGr
AosrELEtFFLpmF9SQb81s8EIa1pP0ndjAi+Z/77RtsKqf0dI/tSKJdcyAtRg
bDznLeEOWAzsWBU2ggt6XEbhS5DU57CtqJlhkJf34SdsSNRlvxEdrhPVXfVZ
Exb27gzKzk+H+dwKitImgs93sGlxuXwnfHn6USRTo54hbZVCHS3xNxmxlrjd
kD6Wj4pHkIDpgoP6gJnkU4QJhAoXyWncYBQLnH93/AdqqjpviVEyNh5O8oES
8KOxpvN40ZXkykmXeTtytycKJNLuaUjRqIxqlMnbOEXyUo0g47bQuUiK9hdP
DJekoAKMbywUQUDsv6u/PIHitO7sm6v+xNsH/HFFYFwcNQYOX6jsGaLxtFrC
OXuxAIvkAhbe06dBIFob4BqqM8vaA5ibt1WNnLiX/WvVAZgDIU/gOJW5O39d
/SV35f+n4Xr9IbHbk0OHaEq2q4G3akQ0eZfARDHoCscu5qP5j+H5ws2z72xZ
u3znS2KFv/yZAxll12owWWxTx9r4MoBR1HI/I1w2C2ZK7+VFAOJlB/ToFM/l
UWZ3qExapNwyh8lWBcv02RZbFZol3GMNr7tr26IAo2VV7Pqwgr2BEsH9/cLb
6rfKDkkTXcw9Sn4UE1OjO6HMAJoxfiHZr7B+DHS18IgVUNxW15pjR7AbNIdW
a/D+JSunRX0PQmgV39wRSaSZoETXVb78MS4RoLJVpoQqYUUnzNMY6PdB3sL6
bXE/f7jmlJXJesXPXrf3rfy+blwlvmDs94KE5BOEq9S364HDBv9OZmx0UnrX
MclH5SJw5tZTbXXZ2UTaS+rucnxJ6/kAYPD2rPgFuYdOyZlU0A9CInG23fjH
v39ygaKuJGskbancQXrVV23nb0AUbPnhY0Csg83RLHygICcdYm6kb50Mh0Rm
YZTtuIpHbkJeni394AJcHdzyea5u0EcSdWV47rsWnXITi5K6oLREu+RKbAL5
rMnVlCBMnPQIEstVo7z9BgadIR3qkdiiQxGnnkF3V8GW45QRKzPP+TxckYI1
BG9bQew+aydZF93V024fo1o8PtlzpSjMAIZY7Quk8HQG4bYqQWIyFWeCVMkq
S36cGYzxJYVDPMeINALFSSEk541oc7z8zc+jOgb76kMBqiTohn40rLZN7XqV
MGEsO4RVUShsUb8xgGwUela9QUAcbwr/DI28AB3VriGQ6UHWkZU3r6bZwE7Z
1AQtiaVwxAQhzHy7iVwHh1eMEO2cHGhgpIQLAvxd4QyW1rkrYFSj/yUqzFAL
o9Aif2pAee3TQXHy0oaoHH743+Hd7QjmAU9eI9mAZmLFQdYFPHQN+Pxc2If8
fENZYFYaaJBFtwzQdYefaInzBIW9RvP8OjcTRXpyKhwKpY8bPfYHMSuuuDMc
DJBn8CG/V0ERm3PshzjDCEbgmt78AijowpUR3dOMPj29W8CW9upjqGtF0mZg
fyy/ZD5DaMQf7IdOZtcl8/tPYK3WEHfIX0cAlFDr6mRZhiltaKkg22Z3KcV1
wWCKqd+0np1C9HprHtQLWbR9fJFpZeWXx9FjjZI64GNWP4vMl7tt8dTcBrR0
mmFwQbdJTsi1oJzyBX4Whr9YM+mN6vvcfdSd+IAAVYTOE93gFQOJcYTFuDe9
KGKHbGd49FIb2xUyr3u8ggFtoV11+6JalZIbQhmgyThw275W8S2aM0FIGfpE
fr0d5PlS/qc4XQdvJmjLiMCuXxp42G58mOs+Zo084D8u7uq0fsr/mN8NJTtU
5lu/k7LzUmhiVEmb6UDnqS3U3E5rX3QKCr95Ynm2KRX+vWKSH1N0df1p1BBE
7cHKDD9Te4VrPdxjjVX1yN3evd86NOSZBy+8Y3AdFCWCmmxoakB2nOKy/FUX
eQNJRx7B3ksxMWVaGqd7LRpGvyhgioE4DN8l/CwOl3ijy6GJesWwBdDQ0Lnh
FWBG+k7VzzeQhG1ENoNutd/TdDuEGz16HRccxpKnq4ukIeKXYAmAsCvX2pre
o5T2zDMCgtaHNCN7UQfv3jM3u8qXeNKZQ/gD/2+x1LotD9OEH6DYbXeoopfi
gePlF7VaAoKSRSADWiALety16EAJzwSbnLyiAN260vfDlR1+C9vZFmwIu6xF
Zsllcm9pZ26P0TrXuXzaQeKtkfGTw0e4890jvQ9p3pmkbXETC2zr0bt/uATT
XI8/OMWBcZTBar8B+Sej38V1POScSz5GIAr675u1ymT/M8BhkNtxVK3zz/Sm
vgzpgkp8Ww/uST68Q52zMnkUqdcP9a2OW5n0Gpqvl/mElxZOTKteJwTNzMQm
uJXN46i9eIauQY9HVStl0h/Y9lxOJs6bV2rQqqehOHnFoX6gU7+E9BDJYUyI
Vi0h5FQDYMMltlsd6YzrVlSiHtZZZltwYn2nggIl/ZUCv0xf1UUDcOG5qonA
pUggl/UJDNsuxEzwxNk+tS3zKNo1Y5dX9akKls/DHo9IuO125ZEc/j5kxM48
CUJXb3Teg5BcbBpUAztb/8Ohu6tBC4jvwz27BWCvfLoa3BpgGmkgxGbFNezf
EOprnjchj1054o0ig+yNanfwFIeJ35S8la3jaf1yXhjEXJ14RwJNqAEXtfrP
r2WQiji1aTLXr6tGaoZUXNh02oh5o7y9tKBNR3xrHsPpJcACAuszpwtY/OPl
Iq97IGtq5w5pRU0pb3cpa2djPwX/xEWupxaiLOtghyhRPYSRjbKCT90KDeQg
SVuGA79GN9ETjr9A8p0ES9RZ86Bxm2RBRRgiPyIaNM3m06VuavlPaMgLizqE
YIEbExj63SfewCGcJpc97U+NIOSxgds5ZqbZUYqt34HgOcQfSOVWpeDSEFLD
USqthmOh1mU0RIi1CE6jI5v8NUUrU9klsg0ijEpVa66rLcfyiuZFhBwX4F4i
l3TJAN1Gs33Vn5c9Uv3WeZitpUvdaJaCY2wc1LXD1tKFGCHkqIRXk8tcL66E
P9jhGHO5cZ2hjyFOqXdpRJt8kERUJ1ZwgVBAFaTddteTOAkiAuoq+mlZjFts
0qJS1FLthJRtgqa3IPmUySgdVXnW4Yl/1zR1iFWHBXGjxH59eV3PH5C1hyIV
rMUoTyMPqO8IvL+d2tCy/hkAMA2pYT9ein5ol/51XJYsbrD21rGYq0Ihf6RT
6tryxJFc8hTHwrbLqUDfCF/5uLF3cr9GvLTMeaL6KNsY8FCa7T6KTjr+bM9K
CTD0rDxQuCQMsZ2LB59hgh/u2ukkfqCgmW65SUnKaU7/o4ByXdjJ0Q1Vu2tw
WliBgrB+5MzJgJHHTLjjQAgWkasiSCqbLj8z2gCZbEYzoVv1VYIHNFcJdAIn
qDohwva23AfrZzLd495n7UdG4rbEHEDv5fQVpnTP5BTzKCL0Lh1l1rH/RaN4
nX2ANRsxsfobbEuZGkR9QPrXPWJxHuJ7BAEFJ7F9pTUK3fBDTScuk9zte6iT
kJKrqLFe1Rgypqkn3L7+lW7oVmCwRLz3ImR9noxT8U0mDpky3riVKyYn4WVm
1c0h8L82LOd9oXFS4pIKBwKVF2JtTCq9Nrjz8Y2EEVWzcRgQYHEYKz9WaUTf
Fcv/pWzTrlRdKlmjpYQywPhFp+QPXeEk0aRX0bnbdSfK7qns1CSjlTr92RtK
cKz7+VQSHRICwpGsqQbItC7Bau6r7XtCMkG5pLGSBowV3qV0wkIkmMD9sDAU
rwYet/kJUjGL5MxlI5tnAA2DIH37zdIEdPvp8oo6ihErT5pvFu95rsu1rUS6
pekNR/GJhhrrwsyn+BiDeZBfRlaGPxqiaTzNlHYWZWoGL2frX4YiFpBNK9kx
8/ttc78KGJQyEyNtmFPKMgKJ5VD1QNPnt9tFEt9gMPh+TeL/ubjIGMDsTM6v
kPkaa24C6X3PWj0NLXtQ9sEwj724aLHsGW+Ef0x4yGQlc3CicCyWHWDsjjX2
vw6B7xHmXnKKRSBCwkg5UdPJ8Z2YpLO4Qxbm3tWya0eQx3LYAdpu96mtp6GW
VpGc3Xn8hdLUIO+eeRWsY56e8T1vqSHKT1kJIkeTbjoGnJ75Bi8EuT4CTDVv
jV4s4T5ePJyV9dpKwUl9L7iGe6w05e7M0ES0sHSHFugj57jSibO5AWAhhYCG
j0nzSDiAezN56h6GoCkcAPJ4ZHxY6F620TaH8SOloZMh4KG3sIIIK2ILpSXu
NRO0lbkT/FmWU8j3ftN1SjWtNywcPY7STAWmRLTiKNrwS2ahDtGl8Zjma2Pj
Bvubp4DBSMce7VdQmVTyMOHflPqgmI8Jh2bGqloWjdQTcGKj0TLVCy4RRKua
wusMd49hGWeSsU/5gqvsGO3E36gslPMwi2in3ReBPwYxzCqzNjHC6oIgSsi5
glVAKo+9sTAezDewS9ypwGu9VvpwhWK7TJnUefjgCV5y9hRelR8qmWcm1uT2
lFLQXKDHvAb/bgkI40Nm8YVttfyHTUWB2z9Z+9dOIA4PEwWzFgxrODN7WxuW
Qkl+1DOtYY6X18C5Os2kQMcn+Zv2FvH5IeujbV8spxlrMAJObIWuDaHKj7us
CDOAiyUU1XVGhiiNqcO80vPUB1/r2HoKNKXwJApjTSQf4aeejtW1ypxW/D6a
hlKhJSf7xy19o3wIJlC4izem+7gTdfUASWKFQf23Qw15qvpZEveyZmPcxYiY
cQlQMPrzz8qdJXyK/JsbgedWt6iUZx191vcigx8d7SjmpK08573r0MK4fgLS
G9TBPZTh7qfkr/fV1AwLzxREyszyB67Xx2xoNxcdh859qjzc9HqzSfOkrZet
y0sP2qNxudcEjKC4RvonG/yvKA+yQTW3puILadQCDVa5U72QilBPQflE2SPq
DmHE4dSMoWPRA7+iWpd9OfV18pkhxwY38rFLl7gohQsym3g+usOlZtag930C
NYDnZRMC0RVl0JzBtNmaLhuEOsYYMXunzGNRqQ9SekLNpI8FP3H6AtEOaYpG
dFJXQbWfQBL448GvP3/mprFN4NjEiR/8MwgpAFvmWUKfLIAXGKIUPVkkwpVZ
3QRn7Da/rAnPSG1deM5csqEe6Hi4p4zOmujhcNUv8a5lQ2f6CrcHhIYKxheG
vXZaxrj5xgts7WmkotdMrW3Ook70XNhloeTps6iTVNVZuCszFaIHZtabsMKg
5oQFW9rK51y1RECIsBqH3XABaJE3u1EMRL5tBbEI0FPEAycrjYTPVHZSw/JT
54szdogQp1m8U69qv8dq2ShglAEXUgGioZc77G1GTvdMRpkyESocCSYxm+90
HQySBj3SC8Q3aKtCYqLzhnN/n92STc1pYoa9Z/G/Zn5YbVhagKLthcV1Wcyf
r3s585G3k6oVQFPYJjRUxvZKAoAzlqJ3/4cNmKEvlznWM4i7KXcgXzW3DolH
04ynp8aiooKV4OD86saGmDKQ0y6JmQHLp4J3GohBbYOnT5zDsURLFyJjpD9N
knOX/Lhlq3MjKYq94nGOkdMSsruB1m3Esc0ptuxENVq7PFpMSpRom4vzEkX9
0Da+cPmqgjgPhz/7X4GqAb98B1kiLeocaM54LefB09+KF5nSAk/S0HZxeXSU
+vSctyEpm09KTesiFZptTfGpe3ZskS9nuwi2FZKJ8xLVuRCQqLTV0ZKvLnqD
AgtSN396sffQ/GZHyeDrBxS7yrsa6H/mGpaomYOolqp++ynSbUPTdkhk07Y0
og08sZk8Igf4XxqaJX2OoWMizfLIZeHqWjPiKjZu4+JdUF85RDCER7sjTwG+
d72lfuteFBgaI12exH1Q3VES7wr+YSfHPA/3KDFw6Y/xlAOT2x4OHDZJbA+J
xmZFS4kyC5zeHtCpEuAw/GYFM6Yq1fht0Gtehbbjqg9Vo43VtUesTLzXVLZn
V3u9SMoSU3TjffuTWgC0SL7RB22Lcj/hb75KVeR475VmUy8cdbd0FTQb9LQJ
AiYvIzw9OMrObTMCuRw4xsemTnMUc6i+pPzuamK8f1sUbOp8iMbdO/c9VdoY
wZNcB8UJfWIBU5lykqIpurbLvigfLca9M8HgBx9oCrMIVvNcXfIqB1HdgHWW
sfKANaqSbVTDxqbeHqXBkAEQNDc75sFZrp9tfsdbiY4f4vniVono8xnDTY4v
Rr2efub/t4HnO66tOKUnpoQdMagdTVWEy62iu6jh0sLPQ3xrP2ArbZb+bLCl
mJ2s/vHqJdonG0Oau0BFh1NWZsNgjnfSmv/GewyWupQxT6/4yT52HuV6SKfW
NbZ/yACyhbx+vrFwqJlmUPXgw+K9cs4xr8xYWh/DAn5CvZn61mZn6AyAKdiT
SaoGncShxgDSxdE3H8Mpi5bZO7MzsR+8m6mHQfe+nKjXAt/+h24xERPVbSuN
lNqci5mdLKmxBpNvYBJfbk6NIKa04BVURC+KhgMbyPq7IWCQaqjCfiK0S1Zb
Y+1qdhzwiZg/e/T0oBw1hPQHFU0jki0KmTpHVoUOPJH8h9O5HrpMKzqbfwQ2
kP3RcmVyuQfiZfNU7kljJ6ks4ka49fPjqJVvjznuL4cFmgsGZgGpeAaIz7Pi
7XZKtASWeIvA+6DIUlpeBjplw+SPufNwi/9OUrXTPcIAkN67Nizgb3Rhjwg0
gltbynA0K/7RJLLZZt64r9xrosqcC975x8+iBkMp8VSsOBnia9VPkHS+LGP4
0rijkp5RF2ijzZAIS2GCgqEyz4YMN+FEtMhr37qT3ctXhF2n5y9a3SwwMk9l
pu8U52/2r4+AlKiYwjvZ0jESZ+AL0eDAs+aiTfDdL2UdeoWqmD7zjRW92SCt
758FELTz84xd86lZTamWXMe/RnYTxzAczgF/m0ejPKTPr2d67Hi52C+06oyH
Q7+hx4Bu3XeaS3J+s7oaOQYDJlTYwOTsNQ63mtlTUhOnImeiuVegXtaHQ09q
5HKm//7gDc3O6EeftQoN1nEGUZpWquPdB685GgTQH2gmgixh9mlE2vyeHhGK
8RjbSbDGqRMafGYik3ID3mpq7mKXG0Db/2HTccXJCjt1hDFAMHNxQd4+DfBl
O5zYMB6eUcjL17yvpd0MKd1GKTexXU1cvC/JQ+tavQ+jRM1Kecu2sFHsiUA9
BO3m7r8YLOjPVfdmV94r0GsHoiXQUVMABI5C6c6FAfybK33sCf7atCmB1hQd
j5Yp2VQnyAEJGM6UFJOLqs33/74r/AMg0+9ojZvQ/HWnm1yxY5BjFWJCLYrp
KnGho9YM7R7bB6WAVN57NW/1bbcT65AGoCvXv1FiKDT7yIA5JMvziv0w20Xg
6OdjBhXAN3+/6lYMP7AevmLF4yTNcwazIRAeLLOidA6CvVqhQGzuCzud9msA
0Z3KBtN6V3zg02Lr4G4RQjdDQ+4cAGX6gQgoaTYNtof5rvEO9lv24X29Ndl1
6GmQj9ifV0DCHooripelXSgMGczQrbWyIyWa+VpEa//9R74SZjLQra7mZau9
jMj4qEhAGMFbbeR8EqPqrNfbV7ovhyDeVLFqMsw7QtQ97rpskzKejvtYN7Ie
Xi62c7RoeuA/mVdkn6XGAHkxUtmKWl7WidylfewbddHWEmbT1w0Kq65P1mBR
Ioy46lqyXxr5WQHTGkEbpXzqBAYKXdO6bjE3Rwb5n1BBBLyC6/jNxq4+HwSd
NAK38SDznxEN0rLVF9liqOnSu/rI1aQ+LxR5oJqoctvirNmbKQXRRIJGLtL9
4vqtuajHDbH7zwYlhLbC67QOMQZA9Y2HZbHQtzJ7Zy5Bks4PY9sGcs2ld5WJ
z/LIzku7sXSu4LDuoKfDJlEepNq5ld4SDebKNLfmqkr4cHUI+E+Yl3MtJxDS
XoU2Sybw8UqSN0LPqnVDeAl/fyQFbq/8Dh+JqCJtRoKOAhCT0u//jG1ip1Fb
4JSDaNljjijbXyH+ZoszT0JSHqCJniOkPyufHmyO+veqEHHzXDB1f/VFcPEd
OG9dVzA+4iMAdm2zgzvV9TFHbSnMKpbWwLefVTqYLVy19Sk0P+gvKoGeEGMe
DmN59Oc3zOjbTxkzwge46alMcWvsPOz/HutvobP7fHq9TL5N5f+HMEp82iCG
FK2dT49iY4Yawd/vf9CB00VmDx6tEflHPaeEQu4UIjkdFwWozp2voiFePGv6
UobeH8V3fCNMhU64SJ0YWHrAb8Pl8sLPAZDfug+wrHhiE4CeTj8fqVCfzQbI
EhWi+PmryqNS/GXmyCNAiBuyCYyPNjj6O5vOyuq/2htTAYXr6NeX5HZFTkLW
tHCTTijPTgB62dHf45DtAkP7T2vY2WjD1huj3CFka/4tdokDnvJnktEKkY8i
WWtUSys2FSoe6LC2S1OY3jlKNkPI8Uudw9Sjq6BqYdNI6vQgTCW2EHjdrY8i
BqGW47aP0KNhy3bVqKcf2WckzfsdUGBbO67xO+I+nh78Ue1Es6+W2UI+lLxr
Ds4Mmiv/k+EvOnvLrL7AwVaNWEhTXZJN3ZOBbTYZFMBko4EuMd/2QY33IN1z
cttVsZLQ7oOfmAOKxOgr5xY9LDbP0hhwgSu4hievuvwPcPtYhShDGoOfhW88
YPiTBYzHbejG070KRYedLth+dakeSF6TjV71koR0GdrlxukOVS2PhFFzKsWU
IWAIjHjDiqOuzsSqLb6I4pr/TfDEGMn5n3kipLdiUnDvkiCX7f85XYfZnBWu
m/KtRn3q1esd9agnALNZn6akjQDRpFbc1x1UdhEfGOSlxNMcP8krQZHTV5oV
Ts0mTGP3jlH5REp83qpZ7+flm85J+w1cxyx7KSGh3EgMcdQe7vVNLbVPMzwq
fNpOQwIArodGdYjqkqCjeHWHs7VzyNtVXbTinU+zLv9TnqxUCYxmLdJWVHi/
V96AyBoSRbN6JTaEKhOFJJuCGaAZ5pOGCX2BKX6wS2CKlZBwXDMQvk4l4EUw
Z6jBHCBVqJ6GChyA1C4vC2hRjdE6v/Cu3cqJHZ9LbtiLLolfbfHwt5sAnvZL
PMTKU+Jdef/UKiVG0e9Wga+ISGJlRByM2zilc0lQODV8xdgi1IhaWkdPthX0
YY2H8J6mZhO7pP56pQiFZG7r/l68UNUJF2LUbs0jo0vT2iQD+C2snIvmjZOm
IVViNhzkQUIeZN4FUK3n7zte2q1nTjshFqM+9Xb+4V4TAEST+FZSMX8TODas
Tc1RbtnRVf40CDA7SQGADQkz80U917zc21ZNE87snmAPQrV1+OWAk+aszRqA
BR3/6GczXix3tdY7moUcmRZOSQHPIReCxbWeiutDh+5pDuJ8+29rk6Yb19NJ
rrbP/YfyG7+xrHvrnPTyvlqN5ampFUI+yt7DRaUAksAk5GJBstpuEnos3DgY
RPcv+P8I2FOoL8x1eKZ5+QLI7XLXX0P4vvqef+mFMEm00oKqHE3JPyGBTUTV
EOXU69xRnyQEjUihZMT1l0nntxdfF/XgjlTf9lnVAf6+sPwSuzJ35qJeA2L5
7aXZ+PDP9Ux6xocPhRYhVL5MB99m3Lga4bfr7ULCOec/SUoKqS9k654/a20t
6yZMg3+beuiCwesLmK99ln7bTPbgJcwlkldKS9tdn+HaaKoCINZ6/KHnfjWn
/hCdN4qbDjHu6+hrKEZxlILNIyXLPm8GXW2XGqOkfBzqRHQFvzckLV958hei
PhFMXf1ZkrSkvHnWl8ILQZX5Jr/V25cgMV3AJrjiuUA9WaqbGS04+kmSyJSx
iFjKWW0QXZBKzi7K8JJQFX751X6NFeWEKv+MTKS+6DphyvYU/TDDO+lXIUlc
h16LlH5om8eIvEysMUYrm7zY9WML7qVqBjsKxD+SDjkTMS9bU/wWrPfN0kKy
uxu4ZfQn/2uBNFUEw7fL6U9T2gMRnEgV3UC7lAe+ApnmC9ZHRm/X+JRuzgoO
OUHr7ywTHTdUH7Vhzbgx6Lj7PqtN9kS4PeEBT897mdaHOhmOUMekEIuWnDBR
bHne4vYOQqges5lfpeB0+6+l2vlxsSOy5BxrGALLz9r8K4vyaFsEsFyL/FNw
YSs2c+O1eeJdyqP85WdNksLn6IhErz6jmcoskRCTv0201+fjh7XQ3YR0vmJQ
jEef6CP7Ej1ttmd/OsGzKYyEYB0EmMztLv4lAXokaXg3TH/BE9Wty9iB/yEm
H9N7fwbOsS4/nWuAB/JLgS77nqHkDEHCCAjcKmMHRNNypp+sBYRM1euatI/V
/Gd8pWa3TpByXcs93MppY+DdiSFHuKWtkV5ipEaVjXGhzBaj4/8J2/TtfXUT
FmPfxm7zyAMli3Bzsu3vPvUWPooPiaYttckzyS0vKrxp29Apvcp8rrJGEv/8
0iStp667HAI1GVcSCyeDCxahKZabOUdPcgeCLytJ45f134a5wjWRxdd3v3cp
RsrKBS7/jWHTzV9N0o1oDF337/KPpwtffHB21k7KiyX/YFKVz81FfSkCFtnU
WXJJG7tTLZNA2yjNt64NLYEbN7Ep3DwfKtpwdCPBLPzehK9Jfui9oXC6EsbW
LUWTZyPH3mfWQT/8YiXnNTg+jiGJB4tyHM2L3M21DQJ67wGLCJ2GBWeHN85v
c3SgYe39RILwl3//+cAYv2a+T6A4igH/l/PvZ3PyuGphdCFlATOrPDXNmAss
pDHMHj6L4/KKq1UuYVnA86+pRcEcqUJzkiaFq843vfPkD4WdR//r2G+4SfEy
QPdnbqnDwfIdiiP0sstGSiZ89cRZbItbnej4S9ALoRwnpehElnRPGeBayzPR
KquhYakLBceBWy+yW9gGs/T1nBXB3tpAoLimFfjlR6lqAC8fGc0ldclX3rso
X8LIGilb6JuoN9kYBYPAX7yjJRgzehTUmo3c/QABHepabx2tkWOn+9jzOiJW
YJ3mww0HFuC9nO6zzxbOpSCK1O2edA3MZjtzx2AnO042Ya2wH3O+I1xnpmgA
1oe8Pimeusf/K+39h6z5+a5NzAxWqbI1fI59OONfSFUZBQ7mnYJWPey4bprY
y16StgeQKcN+gI8VdSpbasZfaoqkWi+CwCWRSnuw//onVkKdW1dCepBI/Hws
okSjFAA2iJ8GxvDiDc7EmzkWDYrH/LMekIEI1aFTOQe2yAYqmIpmMyH3kV3v
LFR5Kh5wXm8luX+bswCfWvbts7vZeNt+A9OdFkeMFiLIth389HGgBUYlQRNl
e+QfjDsuiz2hA+6ylVhfQJtMs5jkUaOVFxxrU4o9nXiVw8XYW87CltTtKr5x
VI3I2RfdKzfDa5ZnvNY3mqoeKnAhjgT6Fs7V+VcrnKDqp/e+o0ZuIjyh4gyX
PqOaVV5RRx36lRfiolxUFe6joQZPYzwj+9lKSGcTIjpmmaYMxpp+wKghpNYm
0koKQTSOGC+oJn2PR0cyEuy/ddnjZLXk1IUoqTS2KEfKVjdSV3rHR5cGvimA
ZoCCwccoL5/VtnLxjWW7MAF6LGdagClSUJsaVAkhXyDulIwvSwg2p4NAcg1E
qy2cuNwX2hLPwn/cCPQ2ih5LBb5yQZcmPgsdTSVj+2CJ6JTi+psT2ZOZUw3Q
60KUuDhde1caq8JLDL9fq/ityvJ+kqkSMbOfk+4xIENiZ34qp2XtU99j+Wqe
6FDGCqj4wvXJ5OXrNpRCLjKRw7wTcYtXsN4SQGMC1ANunSnsWg9zHH90UVil
3kqEvU0s5Dfh0H+LepuAsnsU9pEZqxAxJGJ0zUIyecdmjWXuUlk+PhRkT1GH
Ls1yCpnHF38LuSQn0IV6+Mj9/OEMyjjjYGURuC9LC6CGnPBqOfWwSNETZO5M
dOgl3mVeoBR84GR6sX5oMAfFPUrkgCjTRhEssQ7Jv0mct60OGxwI+Vzb7tSJ
LWeHhFLB9N5f/PlgzY+pm2Q1S9FyKxrUwUE2D28YpYUpwvOfIYDn2/jEjJLd
jOObYscOUVSZVKySMcbCGD9sRlj32wsaRJz4uKP9n7j3X8/L5lIt1tgcRbcR
BBP9gbgbCqaa3E6lwmLtX1voQxF38qBcP7/abiEgsB17Ud790RU2jlKm3QxK
6up8EA6U41rxaVpdigdKiqjPYJ4qHQ6HU9EZtU0DDzcGmwQ1YojdLLyzYLOC
eRnrY30lf/aXIHlGs2OiFSihMCitTpt12VRz47m8XyhJlPx0/Zkn5ZtBgoQp
ssOuwmASbCUXs81SkM8FclDDd/8dX2ysxYzjpmLlojfz2kN0XPwLgCXh3COP
WIlobndCaQoBXGDPvbYgWe01h5X4OygQ55egTZrXBFpLLOtSGNW/GLzviqeB
61WcP/baeaqLaDflTvKrv/p9UkatkXN+nsjxmiUZsWlr023TlX06Bixe22JX
bwpIcN2+l6R/+eS+wsCKx9Zb7SgLBRwIaFEM0QqS7bJt+YLqP1RC4F3w5MBW
Z6DFrw/ZAzZWeXN6KGDpNfXXFSD+sVeX36yWLNzLNx8E/UZx8lYQlE9ryKUx
KbxAbvvOgq5ypJFBkiDOhknxAAaGUFaJdENK/m8ATZxXmcKo92wCqJj5xSdh
kBs70K1msikwdYDZGyKO3S8XkTdEzHxR9kK1fgkPhd7LOzwVZq0XfNWj5hZ/
VrkMGcTHcXWcfjGQxwW8SdJfXW3ONyxypk8s1kMTMG8N8uPFtL6DRJBRtPNs
WHNxLhFrjL8rYFjYrjzFLy70GtraP1rydeSe2AovmdeYu7+xQx1EsfBMPrUz
MbP/aSIhEAYOkVmioGNOnaW0CHx2eWjlqYm467SGsXQJmJiK/0YU+36JX0Aa
sHpdyov8AGUrSZN+KW6xk26eFRBz5UGJC9FkDuH5KnqX6P6YYuK21kI/mH/0
9UeWSkq4HnHKEN1H9X1zFOdngBd7zBZWhnmWOuPJePzhM0TsuKZyTMgmVBcK
ghFNuVZ/khHlcduqfh078vBZUfEeqTTOu2Ke+7usWi5aVpcy1SUwZk7EapNk
jljuGFT04qFvvQ/P8tQ1CVruAx/kps3kMRo3nREm/JA7iy8j/Wjpx5ouZXMf
4qN22oSJ4PdB8I42yHTFzPDrasvfGtJOXwKXIGbdY+Y19zZSFiFVqaA+D281
o+msbdME29v0xqbopw2o6LC+0xirnvL1dYnGbt7OtmuhO+Uy2gB2XPVYeKg4
U97aAiOl78HuTyI4ZjxLGsxCJiXvOS1Lx6ctDbLW1MS2DU+JaIEh7UxpiXvg
NCwnhxUbyhOj2I1ffTiUeBfCHJ07Bweo1oOWSYO12aEcescB7cNSMPiVhqlp
nybCfH+AjG/slzd+rVva69X8gglx+wgfUruRpMLkNa1Nl6WAOzTJD7GUqbZg
//YXWnS6RrEZMqdtiCZ/GxSeI82eSAwkLrxIroS+odLxVpRtfDwJ95lxbKDW
99z89iHTYT83UWvRAoa06HDDQ8HlVwNlqUdoXMcMvbp3dr3fzlfz8fsQoKMJ
hbNHtjMfHye/1MZDb2HpqjZKPOwt6WywL0x9u8RQBELVmpQRb+zvJgRQjSdY
xXqClYZojgOH6xUX5t/ehfjX0ZPy1q/TiP9PBNom5e1cLZiz7umt6SifPtLm
NcHtxHFKtDW/ZGcaN7op8Lqqid5LVLYgnU4NFKV9pGL+9nTqHi2VUgN/iILk
9CKpj8n46XiOmucxVw2O8aKMHwHox1nW0YiH4qBIfKd3pLRapzMsalKFHGx2
q/QeyMxueuOw6+oo8KRLV8b+SZxmqE2+9xI7Z8B2xR45iT9k+HTI1xIbgbHE
eFc5vkJBSlcLF9qST51WkWTKWvfo0w87tzEN68WtvJO5csdPtDjegxwfSnVO
hdnzRLemdLpjSju4fJhWP/NQ+qL4u5J0pOIrLZwPEBbeB44GJNLlzK3VAqVw
W9UX8rhSsYnrKwIIzsRTJ5pMU8FsW4QEfuBwkiQYYtBL0I4KlMdKTesiFU3j
mbNDPnofT0PMn2u4PJX7eDrPWSxPWWm5UgwZWnf9VmFZD3PZDxDL5j6q6Mvi
bO+v+FeypJa3/DlSdg6m6+1v0GnGyJ5xBMkbScUa8K6kabuc/VDtXkvWMLsj
YrGWCxb8xfIKjtznVtzma1lxUrAetAjXKnG5+KHwtl6zxg5xCCfxdFMcTMvC
4Tazo02irKyn5By5TtCgmwZYsaDotxV5GCR7rhhliuMafuO7mSnkOrZqm43C
bM8y4XJkAbSQ5fRk7dOp9w5H60ZPhhXw8JSUEWkNM9XzmNJ98Fh44YkIdLv0
4Owdd62NrW6aETF2MKjGpTWTls9whhV0jFi/5JnNSVGAflPESTFG4DYpGDmy
ZHaooB4beAyuWw6JlnpjCulk+wNCABIl96NdGPgpxqXL/kjzDwJyme67buJ2
B5hc3m+jg0c29Dm/R0KBRbUnLQ3T7IyEY5D9biYkx+Csc6Sh6fLw2QtQ0xMy
hwECkpy9aKi960G7vreRR0yzckwjH9tDaANOFPOVz+WyvLi04oXFsX/ZOLa1
2qgUItp3pB5AD1NMnbf4tJy3/PS84p5h8QQ4g7SKSQzHzVVdSyOiQMhSWvUQ
61/nhppJRMyRuHj2Ri7A3SnUrDFpJ3LuOkJ/b4oIQVBiQCFz1mtnbBGxrPdu
QjjatQmlyOzgmmHLxfBY7/VDbDJBRUd8dBRF7ulPSy7FjgI8mZuUBErEFWBT
hmywVTbN5sHh/gIQExaGhMc4NA3OJqCKCsnJjvkjyL0wQ0c8ORf80wqSPzCo
l16nRQ6e6E7tSrWgp0KiOu0E98PT+EQTnggRSjxkNpaAeIU8WjP53DiPDVsD
LcCASfPw7PO6DZXSlzm9JpucIjh32+4S7eRlDIY6H09RxUmTRv/9k+rowEik
vaEVR6mqTjkMCYo8TdvyVuehPjULSAMYjYYqYjqf+K55vPPiQPuhGr4JhxyD
GnA2OzgIQkjrk1do2QYgcf0IVs9zTaAjRMXd3h3SDLo7Bf7bBZwKcD+tbB36
OGKMDRzUNU8cyEMLVBe31hbez4VubRHK2dFqtrmLLE3izcWqequqvjX1Zjft
heucZPnULfemTeWEK4Pz3zXgbdFX6vnZwd9aROjNZRAMW4gK0/kv/D9YIbrT
31hxty/GFl1eND9FUcwDWle8ROPrylS/ye4d33cHy2l3JCUktYuvN37MTZll
6ehxCrBFkVZ/nIe2TOguBKGv8PM9hJMr0rUaLJYpAwK3XuTBTSoc2Z6++EYT
s1E1jMD6mx6iWrbEsaATfYe0j+T5nuDc9ZlN01lU/pA7if33/3K84JKETue9
Sd5AOY9HRqsvISH/JV+VCXs8+99XUFZidxhqssThCZ/oIY0KtF0NTLOJaTjL
/WwOti2vVH1OST+N5IcMjJW5IQZU0XjjUW8ey+4J09Qn0pvot4mcDRJQ2Owb
SlpiBGrBhe/gvosBdwVwumVG3mpJb3cRMdU35uTqyOmgCpqOD5mRh1ChHxxQ
+G/Cu47tsSFXs1IEyFsaL4MDLZNm085rpXdtQ+nkEQ2zovg1dmL9PPNY9RJj
+Ef8L6ywkK60OpUn5EXWMP9y3/Jsf7n7qFhcbYNTJIt4k/pZu9M/ai9Zx90z
qNmyfsJnQl4QZ7QJH2jpxuTeEIc0cxdbHahzUQdmddZXAV6S216HoFfS5cUY
GxzW3yAdy2P8NlO9XaLtLGtDFl2N3b3i3rV9Xzb0TZipzQR70DM12+C9wk/W
g2W+prGWKi6N9oNChTwOTMpa215bYBgHNR9k38HY9Za4ddEozmYDNtxEj3Hj
fam8bIw0/jUGBZaTkVaWm8e3qcw160a8kMVk/T36lFr5cMNnonUNDkiw0V3S
aeA0DN28kV4QmSChndn+mk/qPVR+KDXsd4SuNLjsfm2YaRiGGdOr7qwKRt7x
tGrnzmX/Iecl4/FMEvpol7+KiWnxTYCVAXz0pX/xl+6EaFkJEOlIBYbRGKOX
zX+pDDFGW8zvsznsgfAgda+Fpo9aws/sy5XKIrT2Eq89vcXwmVASuc4FdJBd
Q+rOR8iwMjnhyNydX2vKcaNtt0d8hKE5W4+LNnnyjrdF7EKs1GakwxiWHOkE
odE8BD9T4NZD4Vpn/ktxb3JdcGCcg9UOYnrmIxNEog54M5GMh+ACO2pdNMzJ
LIGotsU8coyIBd8upOzWPtVobe2HnOEDibFoGTObDfIHxWcXUtqqPODCViLc
+ATVqVfXOtij1TixvYPs0jm8R/2elitEIVf2UjdR7NcWU+V1widhvRhx258a
w569KHhgyy8UtnXX+F2VCnaTVNGpKupc+JhMAEJFWHxZGs/3fsIRJ5mha1X2
MJ8sGM3sh2Ueo30aBpLBbq9F0dDQ3uHXA+AteMoAD9hHin2PmejwbVSGysm4
YphlDgUw78vqzL7SWB7TSK/GHwyp8xnpg1Oa7tuYCRi4LYpSeK6FD7NjfC5d
fYVqKXEPDc4eg2gYCGRye5zy5zWRrr8JwM9pLqhZJjsirnq0VlvLO6GTvq4p
ItJi7k1/Xn3YsaWAqYjdIlUBG+e2NzQZk6DmGeRaNzeDpSHZHWoqeOhiZGQm
ahhCiSQW3LCTPPel0615ttvOa+QxuT3Vh2RXbbrviaQIfUVPxzZmWHt+pjK4
gEuPM+KSVaho2P7db0VKqz+/zeTY1o3EilWNcudqBBbybw9BpTKtzKvX1EYP
MjVIbnZPgBNYxi+YYcTQU6RK4nJA1yKXOvUywGjT9UsjyXVQdXTgyHPxDk4t
Pt6CFOFkGZe973TNkoln/TOIKOM57LBTE3bzroaAtb/CjHhldAQkaqSR3n3l
kOPwd7hb4wHMxef1d0mihksg1IsuB91sRUzuPomajFcH3yPNqI7EknFL4H4A
6nueyvuyXszV7gnHIZvfMsQsfafVCMVYS6b2c/vb06yzlzbtAupl49gkrn9w
lDaAVMYJNh6l/flskxPSUGZ41QfWBeD5/Zpm1GEIQJBy7QZHubrJF0MtDysA
7pELT77KptYZ4LcavPH/0ss7cxULOU8mNE2OqnIKWNhq6sdG059y2m98zgmK
ONf0oT/7dTxJ7THbeQpCCLnnYAME2Zq/zgizH3trodJIRnrwjzLcNZEExwfT
pc62nsK8NUHuMl4/iJ23z90KfOsw0nBAxRupOAnM6GEefioF9Xt/bYpMIL8e
uZvfoZMCGwk9RGwAA1+kIUmznn99unJPt9SE6nqiQEOxRXjYaaAXbieH7yno
ufsff/Buhym+mBkYmzpkJRaaJCpce4kmaaw7Uawc9GMYFXYDpFOJjq4zk88C
KSCm+5P3XJtt6XEMQWBjM6d+NNCZsQO1pjyJ8zP5jZnhIZHuS3trmKf0XPDp
Yg40qG5hIX7VB5TJnz/lI/sNejSB5ozpkVzYE+zKgRZEp9+dJu7xhcSsUIJa
vhPfs7WJ4kpLiZnQtcjlnSQeS5vw74b4LoTfXZqnZ2jEz3MGCROX1WmRiYJz
FfcDOj/IhxuqTrKkasNC/UMnXsQ8orHS42DPsIMocN6Y1pXE+YW5DZFLWsO9
RweHhVAHnH4EhJY5xsGbfjQmZoRwqkUIO7HiN1vaD0GoybLh21BJhRN5K9WK
4hsogaHA5wmXMfOahqye4vUOvHERru0k21YF/90OUN7Nn7bkVRFEdAy5Qauf
0prDC0R0DNGrZNsVFwlpK1a2MVPNugpKLY6qDNhrIOpQOeo04n6w4W7wpfHc
ysKKOMk86jLyIyyvWI/mMxJxI5ZYtBBoi4JgMT1+Z2w0IlR9Rb64i0Tncxhv
KPxnH36ba3VVd3BjHZiN4MvNimlB8oP0PzVr4YytbFVOCDfl1rFXaZDRWrN9
u8aL1LejQHuVdr9y/+najUCySKQvWQBflMnRw410egJKtuUMFPqIeR/2McYC
fbyUq+3fFYXJWjhPMViFfXwncXm/k5Yeq4cb9s0oJxo7TSEhr+zglNjfNrnq
PivOSQ4kXfUkv/Vgwu42/MnQrixwOxGastfEHcakGQnvNE4e+eDofL3W206a
FGaxJ3FHqoSCD6nNEwG/6X3Tog1UtLa08Zz6Rg/Wq5EGlRAUdqRN55B3hPZy
CePA3xBXyjbtyHSbUWerzLCBcb6hX+wcFT5vaXlSaxadWwnCUCBnAQWAcbZw
fQMnykjLNNP0zdTPFfggRfdRZQnW0P1MVZ0UJUxPOv4cXPYAq30dJwnBZSja
5qy5jjgKDFLy2AfY14NDL8BtYyC6dAT82l2J3h73JKNcDWjw1L6EVUGz4G0F
i3WiyLqwTGUrjfvzdcpV7QhtP4VTboMjld1sJfN8zdDxGtHhs0faZwqfGrAJ
ea3qA+WdVWUlKgRG2edPRSgDfeDS+0NN21zjkOiBqTQbYqGLYSWkfD4L356y
sPUKU/8qI94XtFFU7gdIit66lw4B7r4am1N2vXiv14BoooekIAlA3n3q0oNI
0Lds0/bIQpwLHJnwz1bJrk+SMH+1NKDV1buSQosPXWtg7xQtoTPKCr/BfbtV
45QqWuKk1wDdgBAEXg7EJyns/i3vPROErNltWbhdcWRUBVQl+InDKI/1RZOe
5QSa72Ur/o6a+4me6Ug6cMhs7Zv6VY2p/XWihHpAaJDdKUfptgo/JEe786+K
SzS/lu6BParsZyzpidbQ4a9NWmSPahp1H2dPsWnWf+0/Whe5LCTscdFur508
kW9CG02M4pQRGkaojjrmxh2ugaaaGNr65WGmKIT+Gs2SXlkZtxQpQhX9veYk
vQPPHxJBXKnoDZc54UonRojuYAzAH7AAcBY+4KSYr1Fk9CqTdnFBCeZ+d5N6
6HQ77TGD0nVqBdtrNPCL3XSObNbW/mVlMRbkKiCSYgY5ush+7yhcVkNtJd25
XfoHTsKuioaVoVbXxxqlKLGz/JJZhAAJVu/xv8LwFnDZRp+zVbPg9CRFFNP7
wxSRT87sp3lmEOAZgmINGrMT/LMVO9PQZ53bF3/UZD/Eyy8eBq+hUmo1VSAb
3VIjM8fVJ1s2pu9bOiDoX+KZrw6xDgDAIKc+cf80kptZBySB7+1gOv+5/56T
Ijt6ik3hfalMU9s4uA1HwWU1UKnI+eg1jj6aqvMdLoNEkeC8Q5cQZIP9T3SD
TeNIU7kwBda1SE8s2zu5P3Ll1xQR0z3WwVjgmYoe7mgaOFMpvBC2FBlcIpiR
4SolhX8k09IlDC5brJP0zQg4DKlz2Xt22yyw9uteZRCog+7BsSECF14FTjOb
OIQ7g7TcbDCCKoe1q9/SHE4Paphg86PmKkDrz3zYsUDZiikn1hGKYzCvFE04
cyzspWoVFCmIfLBnKK+oKZ0liExdbmrBZkqVcql1IR912TeJt607qa9tC06f
thHj5v4qafqWTNZO2gbzyQJcn20VUS76+CzniXCd3B2vtRRZD0NO/mLlF/P3
8bgQnCNKh0vo9/UkJiwsEnXVTqpXpUcuhaOEHMT0uSYCFtlGLL4cDNXPkz8/
cCPGYvEX/UpcoOdb6eYZE5Fce4QvCF5q7Db5VmJRPvLj6Izl4elnYX8Tho3+
FrZ6Q7KFQxEJf3IdBkX/LrVamHXp2U6EGDKk5c6YdM+um0J87qSQ3oIvGbEj
ciCL4LphhkD2x6yjS1dCdwmRjPatg/kqn0U6b2NQN8i+JuDO/OaaxcXBdz91
/HwHI0sl6olHTZMoOhDw1gSxgPy85gifwZf0prgK39Lz64nuLXvQLaO9F5BD
5jPcpOmkHx6/ZzYPNUI3pMflCLd7yD2tj19wVWF3LDB33TxxZqmO97NRR8HV
JCNeP+Zkw4eT9XPOgnVC0ipiIsfPHfEZ7zacqOljcL1qCE2EM4bCd+U6GoV6
NVm8qaydgsuuN3LxmFbuJqnzF2U+AVQ32Qt7GlV8HfHGp5duF4xaoBnAbb/B
jjQyzS6MInq2nJNp6ztyi/v709W86Du4KK3zuMmUzdwdWjCxYxTUlxniS2gE
dxAVKwt3HCJJlLkvGBte2BzmaUeomXIClQoYGQ4biy3MpDrbCifr8gE1j7Nx
IA8GbMApytEr9BZok7AR2dMUFaTw2Nrvuvw8W8f4tecscHRW74sC62w+V5t7
fPc2dIo+IwVxihHNxweSn/EZhlqYW9yeeLrHJTpdDPlQh0+K1Py9hTCvFJkI
i67zGBxJgzBH9LxqVGk8IhD1fJMIlhMqE6XXAg2k86FwD7Ccs8sGigALv4iQ
Kpi4zL83YLxV9kxZXj1EV1go+nge5EGK95aSTxQ79sPQTPohcSoXjQ3EDL9u
bvo+3Mvwm9ws7jUB8VXY/YZY3wKZOkIUBXEnnj5ASxp4ztLhk82tCsdt4u1y
PZSXxeyciKUf4tfZlMg7v37KWoWnqnhiNE43zk8CIwDO4Bg3VjHTfrj89rqw
s4/Z8vgQjgjFYPPtZKdntWDxwaRvB22QEcb5eL9KrBmdEod5sGJ0JXy2O4Ib
eRHj8PE3XsQ0EATP1i6jGYlh8RnuH4fEQCfen2xzXLtayUUIzNnUJzSxYWAU
4vyJMdU83ooSEBxSoi1HMPdug79cZOuDMd8aj92p4QFAjeV8Bwv1F7aGK6QG
sH7BTRtPTk/1hBKuBuU7djHbc+mnFpYm9UfX5DP9sI61ldSzZTR5ukn+qJ5A
AeAt3VdOHk7DQ/UU4I6vLV5x8TROVXAqu+1QGYFdXX1DUWauZKTCEcN3lCOm
wdV46qEDNLHhzSzM226QwH2hNVsI/C0DccxKsOeznG6t5fV7HOoPUYQL/bfG
z9GUNG3NRu25zjbBEXEHfUzEOW4t4ioewMZSiSi0dRDtElhL4obyuAXI5ue+
o4H8VFvh8ccCHSpAnG8h8A2x5O8OLP/aygca+RyI4SB88omuVCmUkoiEkNhJ
tJDyum7M/AGqrsbhceAfcRQKdS3cvogssx9N3IWOyPOZSvZZU5KgZHRFd0gq
trdGrfvW5LXaeKevg86Bu2rCrWt0w5Y2xzLoMgBcp8HEXuLYYn8Yl8R0sui3
7QbS9gP/EkV8VqL4h0nrzVB9haxz0PzeKp5qSUY61xpV1JWMYIRQC84a454Q
j9MgZ/R9s96ioUP3VEr6n5kZVKgV1pELywkedbntuglXZu4boIHDr79g+ktG
1+VsOqomsMH3Nd4uaPoubE6uBs30Qoijhy/Y1w4xm/Z7TgafCIpInOc8Z2TL
PteNNbWPWU74I6JzhoqnrTv2JS81muCMqTp42vKBG2z3LDtRL8VVkm7fBhez
g0JvauytrnkjT6sfI2X847Kua1Xuc7UKhxx7/0RSNJtrCSfW7B6iBrwYkbPo
b3pl3ZC8wpAHCjnoKtsewvyr3fE0kKardO4Y2FHTyXYyoSydNlOgGBlIcQ1G
geatLMul7noJkJzk7hGiME8gfbhW2l+VX1HrI0+aqRHNDvUe+xWVgJsNUQw/
A+gAhuKzAMSvGtd9VOyV6qD7UD380nTyGxV/d9DbPU013CW+Q8Ll6lGvcAUp
Wn03KQRhcpw1BY38+6J6UIphNSYsMHLf9ojfK5P9lNQrLwJ6D4Ukr6iJiASW
5JwMsnBzM8lC319USTQkb16iPCCqfJFkHoMZ6Nhpa5zLeoBk9PGuqgisQEPb
CDxyf1V3yhDcrIFm07lkUw7Zy+w4WK3oI+r0U/Ee23eZRA+L9HX8kZnlUVAa
4wGt928+dKPW1D9pV8ffan4E/HefSjNhF7yDn84e/yCUFg8ImkXiKW6Mx6Jg
xphwYc4iN3d8tbWXga0g84/UYzjUiIecRjo1JLBKAiijcPdnMRIRf8MK+4Fb
lTHAogcX/bStCzjMdaj2/smEEKEj2kWguGyva3odnjHyo8WHgmysy1iUup0+
93RwCktDCTb+vSpSym1CcDHbi2/j32hCpL5Cfoud7WCPYBxf2hx9Kw3Xbfiq
81h6LCNH4mP5e4rgkZ+FXBIXeozTYJSzOXFIg07m6tAM0kH1waHU82uXZSna
LF3H0pEyTmiQV2zwUobePXHGi+Mt6LLAIIAhCxrYEdRq3obQNUAoeZF/Y8ZA
LUcyEk1xuOvtQEI16GtjJxA1vAuR7YVejiMGPq3zaxVE5LXOAvHqwctRZb0e
Q7fKb1JPv/SVrJ23P3UrLNiBDMhIIfFPnxcL+l+8N/Nbdb85sv4pkbCfSrWx
Shz+kE+am1vQ1IHvk4EANrIqiCIF0B6RRsigeYVPFYoe+YZP5w/oq6ekS8kX
X/6+ZlfsVBcCoa2mUXAaRgGBc4Xy6xVurTFIlxq3KhMWTt7heHjqyLoO+3Q+
01szSnECPT/m7zvUkrTKxEqLy0ldf1t1qDc4OSMeRydECjDtLOKW77WAvGNg
+fXqnkl0R9C/0pRP2wEksauOiy7wpiEQSm6NA9sOE6uzI9ntV5bzxjE5+1rz
Y9f+T/KHzk5UQghos8hdEj/N/+YkR8L5ecz1RJ3F0jMpeU79RgXwWh6OK77u
YovbOM5BEUXQXVWfUjW53YZcLAeDqQ9T3xeE2yV3qyi20iEAhwthi5FACz1O
nWEqi6edyYwJ4aWafopylmka+va3Jki1fzE38Fe9XK9w2jp+dC9pw8A7U6F8
0d5jIsQIExLo+biwsPbG/AUlprlYyKOjyGRrIK3iCT1ck83FWxFVPqJEmses
hgZgQnTR3WF/4Bsbv1pijvTYFUJK6HCJJcnKnNnsJ9XImn8agiC1dMlLuBpX
u6C7oubU4mf1XmYx/AR8Gwbj5vnh9jla3JUiRCM+S4dvJGxvc7Gha8MRmXEC
+lyJf6cJ7VIbJflURpdrZ5o7TM8c58IQ1QJiB//zJolAYFVXpX771b2yaboe
XPCW3US6q9Kh1AFU6U/KcVvXyzk/Gp3cWhb1M6XjflBjo5qx1BRVKCNSeZg2
Qm7G8nUgSqo+hii0Jgkdg0rcBW38is7Sy6MNRk5f7FsHVi1Q8nqzaE+igy/J
5j95AqifK50Mi06fQg57+e7tBRDR+vh98Lp5Fgd4o7GBSkuHomsEQqvVLZ06
OAUshaQJ5/Hc9eZFsmWUpjUbSeII1SXqZcEhKWKF4CAusCN4yLvQv8iwcwfP
kH0GhDStZ+3Q/cSIdhnK6/pLYB9rtmYRD5qbGytKa3N3oa1ko9ZPUZgnyE9h
Uh7VVX7x/0muVVRRUprb9y/3tR7S7CMk7DpCAlVt3LfDPavlEdhSfl4tj9HJ
UnKcahV2NHmuxAPGwkCRvjkKdXNzHRUCXGSHOc9RmRa5MWMM3TXM4EcVIJtG
dqyGl6CEZLmLMCx9qVo+XWQ8MtVxil2DR421mBNEHfgeabIgIMcW2nZMOvsH
0enVuWcSP2ie50Sf4U5IpKULM9AubAI+FlHxECKac4Gi3eT7tR9G0crGTUWz
UzJXJrwC1nF72uoCWMesKOYtAo586/zp2i93FYxWX1O3mdjVdW4SOpodoeH0
AcdcwC6ezKVn7M6/N93sU+Ti24T6M1hzi1/Zv5uGZ3aLVDn56pMlhI5Odqg7
lLVV9dQJWd8xp9abxyKGUNmfF1rWBXoUVrQnsSGR+LKCvQDcB4f6N8luX6RA
FYExAXM8rTOQlEZn+5Yz2/upLpumwPHPLdaYw/aZabQ8I+/URBAy+qP8S9JL
u7ASgwO8cNdgEoU8MJDEyuNUAx6hcUco67HqZ46QpQkpyX0nlQDWe1wR7s5x
3R7rT9Ka0Aqm2WGsVyptFCjki4+fjg8s8vm8jOOeo2Zn1QM2YLeNtik+W2Dp
QlAXlW8RKIC1I8hF9uFxtnIYUWiZetiRQJ8yS50tUx+jrsmgRPqfOWhgexm+
qZVcZCAS43/0FTmMgnyjFKgMjsg9iSTALxn3BSDZw3qpj7Abt2aKBv6lSlVP
uSYxVeUz84tXdlZpTr1StLLudn3QDssWxzAsVNYKig5KtC40apbl6Lq7l6zU
kgJPtfXPC0s4/IIEwrLtfMrpBn4rAsrQ5ghJOBD2udUm+LBiQ3hW2mTHktXc
M0y+nT4KffmBAyUS0LDBXtwdyxkKkBeVRTVDZemgl9UNFVc44BwOSdRetZZF
QQVpy3hiQg6Q+OoE4XI9xEqqMJ00SsNYfMc2WpMlPrGVDJfJLpuV7XemSm7g
BdmlaqK+VzeWBI3Hx2aB8FUWLMYMgT8yEgHUNACnTZ3Fqaz5Ay9+0dLJy2jI
l0lCRopbCb2uqPAxHql5QVAS6dL6xfiugk1rywsDOy14Us+SLko0LvBryTDP
8t/qPyoCfWLyQqfoTnvvC5JQC0rsQ7LMgw1YXqTFY5gsKYcBTo3wv7ygrlc3
Up6T1aeWetYZswdsViwfani5uXUAXs7wQG9+Lddm8PJW/DeFVJnAhd3YUgOU
r5Axl6+AGmc+0fEtqLf3xfX5WJiLsoqY0Ldghm4Mw/XEkevZneWXkbzeP3pf
hexeH1sE59KJAe0bBuW0FE3qPaQlHUDHNlZSHHX7OWhzyevIyrKfaTWlxkUj
iWna5jSVwz0uZeMo6eEhAQOeu31BQGPhBcAbaT5sUF0pCxDJPHjEvY6Ki00B
dG7PimHSl8idO8aV8x4WSMMJRhRfNMnrLEkyS7eJ9DgF8mjr5hZdWnjIaQtS
CbAa7THAdFVp/Kvsef5e+Eq7UyGFVIh7yQKIT7MMpTzYcko6xmi7VOPUyKGo
qKgxznTKWtD5c9hEqqQiqc1ORdZpufVJ3Z8KKB9q8OYpI5d70dO5MX7F+6Sl
SkW06AhBD4hRbg5AxVyosoOdol11r38BSML/P/1MbqS2vioWzPMAQ/DmBoBb
hsof3UJp1KAFellzPRFMSN5GPiT5KKCr/EIVfM2bC+KfBsJF8QcNOEdb1GUx
UrVCw/D3+E00ZWgRTD8J61FZEcxSaHswC9AcZ0TciKhAG3bQ8WxUCjp37ipT
zsEnQdxnGSq8S4Tvdt9FiFmOiJLzcWsBY7717mN1ts+MgpkfkkuCLNOd2k8z
KQq1OOYZ9eplIv/KDfilCpsJT0an9tOvuqQ9A/ce8vO9YUBrnX2bEVt0E9tr
bG5WCHBRkNZZG7ze9pgpyGMDjHu0Domwuclg0IgjMGXDpSVTHEeyN3/32UAT
+ORdis8lF64zFCNc6v4f7A5qZEfgnAPFFLCvzZWy1Hc02PMI77oBgyOibhmr
wDoMFJdDliNE7m6uztTK8COzmwtxdeiev9aJkuY6MtJTA+yHga/ip2mf7PIf
SZr08PlOUQFZ4j5P4cbCx2M1202S53PB1O1luqgadTuP6j8qbLGcsAMB5fRl
2cVfK9XcKaiVSytqXZXm+6r/MD+B03RI7c3p8Ok784R/SbyrkxraaeqqlEc8
Gtpzhoev3hLYN6stsLA6oDVnML4/YeJcqYqByeO6+Cm29j0rDNhUKYjJLiiE
AYMixqCFgi88GZ8tp7fKT5J5j7CoP3H+0ujXriR+ZaMON3jLKk9/rMC9JtiQ
JKcZkaeeRuiGnDRFk2MFM18PDFSJcmAhXFlfTGtgpTgEEHyORgOcE7K8OVH0
AIdcyedlduCsA8lwlGnDHGFJ/HzQP1yYYa+OSEyxVTHdRHRtFOnpgTXI2Nva
wcNd+K0r0ccU9Aol+k8+MelM1CIvCuK1RYQEBkNonSLEvbI5DwyN7Z2q1M29
fmHe3CEqlwtdXmOXjXmCXrOBmu7DKM/s80Xd1eS8xeAaZW85m4hKJd/SKJUE
2B8PDQ+fQw8I6SFXBN7C31JfBuW1iCr/nFxOi2mf9qmPzJH8e/KXvLSSatAb
LXB585wfokotknL2DKBKb9vBm6T+AFZZiZSikJ/ypWLR5I4mXZvhO+ISl8cp
bfGHUtELcNDHbanil+pCWvMOReBlqS3id7gxGdQOs26Pr0n1Hy79QO2U+7PG
TCxDnmFHdvGl1X3/GFA9U7b9nY1iNxIKDieb5D7tJYw/7WvovrHui8fOGiMO
pUaGV0V/AKylEq90ZYvpKzZ7zhCPZp9Wp0Yja3VSScXwrfaATApcjLCNBdg8
Ys+VToNdS+M+ELH62I9XplCZoryx8AETZ2ZPOl5icDtPOp3G4Rsjtsiilyf2
RPozTRTJrvIVjMfiX5vVJTdhMp26brcHCxbaH4hx60DeR3VDGqwvwMcv+Ic3
rzeXJWkL3RwPIWTiCK3prTtrQghKCN8dklhWq9cpK0ldkgCSgpgHH9mmnrtv
Sx+hbqAHMvlJ6JR1T5LQ9o37xb6ULEV+k/LOqthf4AxJz9m5oA+1MrXvaVs6
C+yqE59sNnfLECJSTIO2uYVZP0iw+/FdXVdx0pi3I3+V5MHStY7zhZEpxZFx
HI66pamaLFqoZjLNyfpMmK5NFoT2MTD9K8LkiVFxb+jjHjxj/l8GSVvYWpmT
2GYBmVCqOvWEzH6OZGChleIXKX92ztssxxBbyUlEFLMlnPht1ujB9xXoZzd1
OorxL9865hrjN6qct72uIRVU8gaLx8Aj9UW2o4nh5qHwZanUOsetCh4EAn1I
AVl/uJ5zhRREfoTg11ssvJZxZcMxhuriTov7RfYiGy1KpITbptYa7WH+iGZf
6Am9Bx272fyjbsSZTPGDPruzuFbuS5IZt7n4J1XVtDHfHiSiwdCh/7KpR0i+
Ym2sBKcJS9w97UHllHJ9sGsw/wiWON8CFQZmxK18wl0/mDoM7QgZxq2/BW1B
BJFMPQrQb9bz1Cb1CGgjRpCbOW+HHxsXJUm0+NuEkQbIrJeQjWgYvBlSh4+F
aMJimRrRGMaNNmP9r2YvBA5jYhFc8sq9CLZfGelPAEXdbM3MTtac07fojXa5
xUasBei1Mb1T4uTWwT/Bk+uaY+RRe1M67vFVdpas8y7++Rqsu0/qjF8djRgX
3Co4PzGC9k7CSm+2E/HDFKze//Tps34ggxIK05sEyqZi+SpoEWF/S5McGXsP
HbD1DwKvgUCHo+/ERFjPAYI4R9RioBOGmlDpEOdCwHSNBDMmKnGp4pxBkW0p
NKLh5b4bIs8OC8Vl5RYvLgymqrOeU4j2WYToNFgZRyAL2HgmaUUjg5w0h+Pl
miw7KiV5h/InlTT8nmi/+TbsRVBUD8LERGEK8pVhtVmS0Uxk48WDKJ3kCQ+4
eIKvLdvCGpwsk8BgjOyIQnOa0nKRmLvmM0IX/ILZ0rPPiNxr7knAvQ4Z5hN2
urQBAEJtXH+IetoQBHrRNo66MXBMQ+Wb9ACl2X7whKP4pkPxsN1KaLfN+oB6
VEppCSUcVhVg9jBt/TWg4z8XV6zn7W9/FnSSVEAkwVooqtEvacId2WEHnkVe
6fVXBQ/F0G8zXVtsgb+iasQCKzXSI3cWibHwxOZEKbo4m6Hzir7rMNKjXLfb
cFwTmcdvE/Dwc0XK2SsUIuK5ZEhlNhYhs22tVweY1PpyAIFFmLThMowgNECB
xjPBcNlc+ptXZa8G1tvZtNSHRKCzChsq6v+oCHMotWBjoCzZ9QsUe46ZXPDC
tVsBBWebw6D4Jezq58POqAVIFLayAV+VB/pw7lJY06atdcy13bl9/a36Xama
zKPdglQja4qOhttHPdwiZHbVcUbDMzrlsLBemeLgU5pAAtC1bNaDREyWxNvl
YYBj968+T9LiGJ5MJoCB4esoMyQmr5G7cGhSrWsXBIcIUPUpkjINoGWtzO5D
PQ07qdbZ62FiyY+19BAzMThigOZ1MXPCHq1wD0R2r7fkxLyymAiO9Y3VmM4q
VN83uKHX9D/xkSH7Hug+0fzxgRkKUCuP3AYOLss/Z3xYAyTkkbo2ULGKCj49
OtuKAmQXQ+h6b1Fj+z+nI7CFou7cOGL6YAgX6uB7O8HJVaPaFr2HoyokVlIe
jdHPCwO89QB5ebV+rVRyOKZ3tx09v1BkEXsALCaIc3eivVHh0Tci+c7xtk7O
1nKguK4JsabntKxBjP+N6jDsl9fOlf7626x1iWveibrn/ZlvcK45kLFmDRK7
qGxsN1vTKvfHZFRsEVh3qmldAPoaOolmqmaB6XaeyfEHtm/IdONR2OpeIhda
fnLee/KXSYxam1zpQA3+7hczl7ZdJgPM+QsBSziEvbus6vx5eimZvAeVos8M
PvVEChGpkpKCaZH+zwYJy4b052qNMLCSbo68aiwq7huyjz9uhf+Dc+LjHGnb
WM2fpflQhC/7zY5b/wxQqi4pbs4FPDWMKLj+d2SPihyuRBDehAyIUHwHh17s
3NPnlwf0FTxdSNp2gD3U/5PT/qJ1FwkyT1EYAPawhA+XOrUyj9uZW3l40czh
OCGWetdmJ4AbSJb9hSqm7CS5EHH9dsnR4/SymSUwQ9p3MWRQY+1D9CkG75Gu
CNr226DkxtCizktHS6bCDkM9YUrerIjK73h147dwm9XioKAGLL7wKqvHh24k
Gx7CgRjYM3j1C1V8lKLRcXFhgmCDxNJe2Q21pc9Jiy1YmGz4liFWgpp2bsln
bHYVW5E31MHPDbWWlhtUPhsL609h5vRqUIca8h7aqziuEdm/AQOCSCBXJkDQ
3IMtideeeOUnq9J+4nRnZIUjj7LNblbwPtufA5N8+Oya5FSrt9fApOc1y2uY
0fHNSh++Do8KwUmqiJoyYH95cHlrA+kSyTyzN/XWidNO5IhV4BDnkQ7h1TTl
jcoP/pN3JxL5uzqUdztbWB9uHOxEeFTD1TLqSy2wawfxdOoWR7rh7/eYGezv
tXdoUwyE9iAjBXsw3Hw+IgkPJvUQllLvsHn9hjEUpDwM263mqM+IUAGjw/zj
27G6aj6YT239KgFzCv7Wz31HTRyqf/eAmF+pT/pbXGaRCLj+Ie2pNsHl9Uzj
Lli2IYlneJzCdRcJlCE5JO2ThTdrgnRj9gx5IgnMTPha+YSPJsqnIqFT7SXB
vPPCH+zNS4o+eR+GQF+5nYRdBxtu8x/7vMxT6cWdnrLa4wL5OaVvYzHV6G4z
WtnZjBPHq06u++OJkdFTP0ssgDFp4XrUXi9cY+BSkKfi3zZv8mJ4wrCKgYxL
/o6tLuHma8LOHLyJWJ1JnxnKL2Ig5ggoWvaEWN3jp9lzLLtaHRSx9yR308Ts
DdhGmYsMW1NtPpr5+00kHqY52+WlZSXUJsY1bgA0G48SVmUJ0cWTgwMmDKtp
7YdU2dofZfqka+g7COSD0gUseAjQR/H0jueSUeZSFEXQR//2PgtB7CKiYSTs
QbkBHjlMxJiET9FtSbVnL6iOoiZhWdQ6kc152mvlWUv942Z5GYTwbWuks3Yj
DSga/eWJ6HJxsFsL+zMKlqbRYxIIX5bMxuRKTcBj69Hdbk0czRLJ5L2xh4la
vo9Yjrook4UiuGLIf89Kq/A1297HTKZMkeo/fr2HcYW2pXjcVKj7+m7W6TY3
GLPnG7j551otbKFDmI2EhWIyE9MQrPv+ciHBMwtr4gocKams38tc0FU7zc9H
x4xEJ1TYgY82N1IxiAQgSXCjzYDXSI654u4Ysszvt0qTKq++bfBY/ZRy6/ys
kFmYxIxqamfTsDcqgtavU1gJEun/34OG1+msn1JYDZmRRbWKI/8go5IUBmhv
2m5VF+3tCN5XVAd/t1QQ7Ls6cfKSrXK9ms/akwWvc5EaSMaDqgBo/TPHt9MG
kHtVhNZcEm2QPrjnojYXs0/wCJdw6/IX7TXlv/1vh8NjHD7RLybVJ1h95kXA
dNW+KEp76IFIJKFUXXgyzRIEsMumzPcLeQi5zViXZcZqY3Yhr86SFXcGrFIt
uOYtGFjPvXVUUfzfG9rlR0YS+tpQCM17McktGTBsF9fndLJX9cJP/xuOQbik
+K4ooxffAM3cLQsGnkfXIvRxx1NdELKP+22ULzFrV+jb1zRpIit4E9gFxYq5
hYGzSuFfe9cRc1ZHCLI4DiGkBk4ynKDUJCIEPYUe0zuALn5JvM8oxaRoAHz9
I9FRCsuSBGSAufktA3iGkYkuopqpw9p+wF6P9Wt60bG2ivqPb0kwC5EjfmbR
GWD/iICdyDlpztJ86w7lfh7TBn5BR5pGFbFLA53XMZWsMq+vNHxGrOXEOchJ
A50LCyiJKBVWt27hc8sETyOXhRxWDwDuiLIlH0xmGUvFGPG+RAjlKpIDm6t1
emd8gzBeD0Hcu9jx3/7FIsqoX+uvJ29zfzxP0q8WX/y4Y/rYzwczt6jzDl2L
4Q8IPen/p7MEyj8CPaC3Oa/r352O8ZlSgOXDkT/e3YdPy9LY49nmIw1Y90KL
j7vOEyG5uZMOb0PLyoWPRnvA2cAcjVOtErLYHNX7Mh+24QYp3sgJk2tvCo3q
MmqPGwEu/NtzXnB6tTP37IiqMl9I/638S+Ap4yUIEqzkj/yBT4MJkytzxWDN
zZaMxJbTJCIcp/RIAt/DwgsUKPsgwAP9/I5zkPdQE0PQogwnZERN1OkwlXjC
TyGByeKniGdb6DVtLXWMo2bxl7xKQR1H4qkC74EAsivyyBMxNb7RWkQrlPCd
XJTdKg6UoCp1iiYXZQjAn2zE0VwUgWAkQ2LxtuiHT97NOY6EEHdOqTvHU22r
F21TvgfBIOSAhcTVzOnNDiAB+zGX5/NmGaoXVV7U9cALhopxXpKdieGlrAYW
D/fdNQ/LdiDS87Dgc7lYsnM+5xwelqQNwUurSr+vaMISZl70zBb0XVsIY+Vj
oDEbLa6f6/Hla9bhix4QLgb1qeG3+wqmJVN59i8cb5jWu+j8BVS+KKKULILC
E1lCu5WaJdU5/+2XuEho6rDJ0T5tVRXCo6JAqMYvDLPc1J7SJoz63C7vpQiV
umFok2f5pv4K69hRJZQX/1frobxkCPKGqnfxMimGqkBwMkZyGpTzIMtWUE05
XbkQyYI7G7DEUM2jbT/BXtFFn/MgY8cAH8bnfP1enFAEB2pPA+UL/eD4z3ME
P/W0074ldfHZypV/m1F/f3gvRb2SixZNLTi73Qhfl/zOWYMdySEmM7A+hIzW
DtB9DOAhX1Rc4EgIgGUqmWELKFot0Ln7en0BaoMXNZmjk3g1Nj8u10i3VByR
ARuaQlHJCD8XF03KRsVwM1vgzXVs02PRg6h+O8NmvuOcdAD40fF4Pli27KMt
FjIyNts2dFsNwjeTytJ2c9igVyRKg9CoOz3yRuYNrXri0rxKFU1aEMzsnc1Q
IXInfhfRGRG5bNGSglVM8eayEptv5jROSKWbIwwscrBAqLE3+vhWjt0XFgwl
WbIjbaDkfrZNYwENe4UQRq40i5EurNRF07sRhw5vveCc70/g6/0T31RHcxVx
tJVBhbneqt++Hy1FUiDJcgUveAmRzpOmnupzlIt/sYyYlEcIvsQ4KYHJPGy4
vpFEBWXu4rUcN51y6Xym9amFuZqXdF08Iid7rdDulIL9nN0s0ngcU6WL0AQ3
HqL4hFzvShPhlfJ118XPVsZLXA0rbfGtndJRDB1NY24a5vlWwzmiTY+qwClD
JWqS4TIwxCn2U/RJV0kRLf62DfLBB+CbD0Et5kdMhfXDSzI8jvxVyIWw2kBj
OwmaQp2beokvB+XpQBv+e6Ep/uVS6FxOkgwOO/gEyqycHA2k5+l2iXd8BBYw
X/NAOGapillp4/adtv10uYY3rURaQp/MAcpKjxSH3Y4VspnCpOxb23HW3AHq
/uwbao//cYlwSzfEda2kaiKd3CPbn10OgB5PGxYcY15hoZaAoOhW2vFFdR4s
PjVS7cOfljVYgylhKTYErr4dsKOmThrp0n0IndQvftibiVfsHfn8pu/bdetI
89Ni4Joso73PQkYbQ2BzOuMWrt5ypmI3hYbcaAuDLLiGpvQk2uMClWkv7S45
whCD1SGVP4h2pqp/s5BrNiKF6L1HwHpSOTBonCipDb2sj7AmwCmRQt5/ZyXi
P/yIte4LGQS6tl9fYKk0FWo2XPIRux2CW+k7PqGetk4mXlHpAmiyK3tiRNuK
ecrO8LuBVwGI6O+cMUe+JgOugpI/GHcLXTUgBNQepRps70s235tb5TOnxNZZ
8IWkiyQ3gmbUL8+CPAtBg8Cz6dJebgPnJf0czjCL/lDRcDoCwfSk4OTnvsLm
uyyKJ+C3XXZRuRY905jx7T4k3r5L333zipo5yVtr95RBw2PmRYoeT1PF4doa
OWPU9QhEA3lPJUQdc9DD1DBhPhXNkil2IRWmC9/MANkIG1ime9XOpMILlDik
FkA3vMsHJgwuOTFyqn1pUWGmM/UuOgCm1dw5PtMQHDPzb4f31PONUTcAd32N
+RS09zwuC0daNnI/wFmikhMxM6wIKW8tG+V1SOP/+P6sjMij631G88JFsPAa
tE5xlTfjqkbPTRY6R/VHTQCbD5kXKHXowtG/40HUV+pELGAgoIXbhgb+TPZ2
SfNZIkLX+NVSti5zFXknyMroA7tXmet+X1s42HZZefY6A8Cbv9iGo67+nyaW
eAdA4BplXoVMePyUkAtzxSZYvQOuoiGW5ENkYBS6PwKR3s7PoH7DYtzjhUIJ
rqo20r6PkyKXW4m2pxGwi4tHB9QfiKhS3PFhFNHtKvoSzcBwyNs8v0FFPuiw
Nxpj9DRCg2UkxiGHfyxoXWPBlPIFvwnHcmwxkaKFzPjU4ivXR6vBjO0EXm5q
7Ap4H8tvJQumTe4GTS4i4N+KJOk+A1NeZnhLzB22rVKvHwgmsO54uCAa4NRM
rOP+rfGL6/n4AjtFuVQqK6IPYZbx3kktaeHJOdxJo/E3/SO9dOUtYRsoQMmQ
TDL4SoXljLaa91TCaCSGqwiKiZOQUJYNuCwwrBZBnwHwZvnXihFhRGvR+21c
Y/OSpw368YxAOdmC6d2EBh/QzcskJSa9yVEwcKgwhWZyuYGbVyKkN9tgNF38
lhvs/pvhgd91uBlCbTISzpOPp9FuifoFAW6heljDuySpNVRYmfgtC4t8ZiA1
cofSQ529+8M/KMBnSjVmNNdfWU7j96vYySElxvMPX3+7Je6HffVjsM2FRKcG
KOZ0VZ5M2pNFzF0vMYSaLhVqBOa7yo2YEIM0IO6SWeGHnhDY+9ELAZ/Xda85
58NaLY2XI/7JLu0QwUuBpQP4B4pKdTAUyCvjSBEIVTefZWwVdw8uxw3YyVkz
7SaW29cYhbXnRpW7ue32chED3KlihXOBGpacLTVI2X8Vm+my4W9C81vUEFN4
WPZb+qWjxYWNRKbtlSzuXv/ZrrggOl6FGL3RdjukPzxHPcpLtY3UHrKTn2XB
j6mYJQH4ULMRksXvZ3Yc0t7xtTexVF50OSv+ZIfbsK/aEWh1YEAsGB/Iqelm
sEPEo+IorDkfWTHZiuE9VVRccONPSpDyF8Rn7RG5TEC9FhQJnOu+lh86dSDf
PRmxuUFvr5/rxgrlrR0X7YbK3/ZRykCCRven0szPJbxYWlwUhN+nCzPabN4d
bt0lyhxueydbGyQ8uql2CFAvVS2M1l04Kh4aLR26ANixK7B3sJ4Qfd2a+hdN
eQIaDD0L5NBIQNX5eInnC38eDXQTVQAmBThxah/u9UbEqvYVd2k+k8PKKq8O
1zJOG2B3S0Rww/bgOj+gV+FuN3WJcQX3G419N6lXUK4VDT22Iu/Uji9TbqE7
1k6JEC/JAvvmJAH+wF4N+Gj3mwAfkU9dwtVPIQ+Ulv039DWKXvNteSYpDrvV
Br8HttxrmTdOanNLWK72Y6VkBwO9ijni13ccebBU5icdUkld84iVkM6k3gcn
fjRpX1dYgl5quH69B0oeQhcC8pneGTCC0M/hW6cQvoMl6cg3ZpKRBaKAy2ci
RM8P/4PcAhUXcSLXjH6IaGwY4hnMMTQ0bulV7DytWYDYjPfzUZ+2gf/NBF/z
L4tGGpqu0K38M13NMGhJkL/HEYI9ZaWVYryOaxVMsghnQILXJc9ENQStQkh6
dP3Tlz0IGVflomk+3NyE1pi4m9vpK/Mwst8NDtSgWvhUyiqkZach5/CeI+4Q
1tyL79Zh+1YiPr0Hr5WHisCK/OJDM69kdOI1QnVi4bvvGKjFuql1EzCeqr8K
bpqdCr3vE2Kw/AKx0iTO4gH91hb9Rr7cH+w5TTDTe92PwKtIXwZTkhuaahfe
kIPLH+4riu6/Ow6JRY3J00x1i495HR/MdkRrjZrNEk062s7fXUnk7n0fkiwq
BoKYc5Iz8VYCOzmUQET8zCtv5BVx9hi9JsSzEQ8w1Kaq6m9gL4nIVyZ+rnPA
DfFknAy5De8S/o5CcZzAMPN5YfgRiHrp9bJJeFucpwIxSxFUZZQSGWrTiUHP
uQ3nyIl1Q/kdyxDRGV+S3GGIrcuT8I4M1dKddURJoIFaJBUsb/VNtnYARedN
GwKfh4Ru72y48ZliwNnRVtkVngeGV517at8Y7l6UEX/FCo7kR8fdvzdwv+og
x87WTQrlW9x89y/Qhb27yhS1kr3GRq5qK9JyP5bKFLHMAjU7MauX1eyI/clT
1Nch1Axn40G9fh8l3eYoXHVC7Esz4TRZJ+ZflFoePpZThBO6UkqKcu0/Y63h
bCeAp7RvshifzWEhYWQrP+y59YWSO+TBQxRI3CcS8HBsGEEpImaXSClcFNpz
CrE4tnzZ7mDN0qSMoCCn5exOhsblsL/uI+Rpoyh0Drp/hRMjigDGyQYc+lB4
zwOMT6tg93XYZYhjRD40eWoAgD1fLc0h3R6lZLmzqBzOzByq1hEVSN+uEczg
5QfgiNqP+XjlrWfMjGIfex0wvjWDWQswBlowDmrEEm6mXHRFl88EQCdEIMR6
kNen22PnzsS3KMn6ODto1kzGPQqaU56s4AAOy59dvlHCz3UmjZ1NDf53UyXS
DipI3jdmFU2UcH7ckpV1yDub2Rcb/7bJuYSZ8maLPN/WGEUmCKCmL8mfCdl5
J1KfH/5qDxGJrcGWaC8iy33pvxBL7CMIn/UV5MxCkA9kKU9w5573lxeumTX6
bhuOZiXXKJXVZraCBwfttoX0qebI2oThtsVg6aqekJLIciB5kKpf0zfE06cM
OsSJb/4J3hZpRik/fj9P2r8E9Dk19JUWxB+vdu1OM8W92q6lXk5OWmeek1Zz
3bzP6oWFQMVgpDIe+zf3R/M46ZV3H94t415WEdX4FVLZfK59Z1LBIqLE2uzb
M+wTVc+Y6if3nsNnbGDHkta+ga6qI9sFd7Pryz8OLSUur5bAvIMin/Zxqf1V
SdMrJZAySIxo0YG/pcbJgJnOggQA0OthCdLNKd2bIEp8ABsY5CAUjzen7LqF
HH2/8U0B+cfI6YRv0BnjQ4+fNbrWao+US3H5xI7VkN7+2qOSKrYSbHFpYWQ2
zaoQZ4Jh1umD1ElLpNMgcxPMo2wuEhU9K706ot+vFvm/ipVBJQxgjodbBRe6
B9c/kvZOCm6BQNWmthbmcHFeqFQ/oUBis0BmykDxL9Kjnp5KqCCJUmgrjRss
IXQrHK3DtHeTuYqcML+aa2yJrrqZsXrNdHpZmzFdD9PAh6sH5eeeRyxmp7dl
PoFddLJUx4kAm/iZSnaW8di3Z1wfnyA8DwSLy7Y2aWAZJwwIBIVG10iGSKFC
AHa/ucFTnnFQ4lRqbAkILh+kMlthn4VoZ+/fiH+olpiLpBjtXSUS8gmh8hUl
svOoWYKsroFQHrDVWO2URyDjHNxnx0ZeiQI/m/a2F//Bhdi3CCG1rpQFKTVT
hBykPvLVU4Bj06PQWDkqQiy8g7MoTwYvYtNI9Th4JoU711FVOd8RQP8XTZSE
S2xUWL1WgnVkTmFlprSXu9EC4DzMCU8ag1/YHwVTYwH/q6FzYenatPoizIOi
CdFobZqWi8O1G0WFmgcfA10g/Lqha5DUrdflh+lqXaiw/TFsOv57QCQEasUs
Klbv4oGhSGVmXV8ZRRXykcFME7Esd+qQgIyT1Y9Z1DZcNJcRyGlO0SB8EBqt
tqORkRoR747PczPUd/eFBynDGmdf1mth1dgDjWrgt4oo1xxaqbiyBjsr0DZh
NGPJe4bpY9KhMrU29/mcrqgb2Im8pSI3l6qB2Tj1qGE14+WDxKAV2VmHH3UJ
4viN+GkXbF8l+sv5I95+YMX1/sgs7ndEnPi3926wAj1TMJEE79TrHt0WwYBL
KHtYB8z569rhRSg0cvTqjlBsd5BQ/SWsAjWMajuTK56tZELNbdjZk8Zt8BII
lEwWlmlXFNlfKosvX9DGKWeVgHhQsgkf5f1zavg2Xp+1qvQ9SvhY52DfqZ7u
1f6xhLE+DLcF9rfXH6LXrThUCgM4y8tb5s/Jb8G9XWHTbA+TEE1OhAQgu5KT
movCNlbnuDBVtkCyCXeUD7LKnLYFqVgZDBa1wFsrow2FOyXREc+oWIy4hgem
josE6MpB1ZuFBbDZNR1mhtbWooxTnckvWfL7FkiIJKi8jEXbd54OH8UrlYjc
2LheYU7oWmH05vlUqQCVPZdbGuBY0M1mg9ffqmoC527NcCk4MIAdllwWqrLr
HaI74/zAwOlANz4XXF+ecfU9nQCL3rwiyh5Dx/IeBk/0BaU6VDYGRwx2Vld4
WNbev/3ag83F/btvTr2wtxj9ARtjL9HsrGXvhinafyn05S/S/+8jfK+emEMJ
oWTmrPm2dygIhk9SlQHsRBFQLlJGjO6aqd+h2IRhJbSvhL9za64q/ha4Kq8F
7sdqdEwWExj1oYnF+qTHoFcFyeUn0OPoe94Eh9hZ8iqiifpEX1q/rDxY+wr0
pALcH0JbJQW2I1DgoCLsKeMBDownEjNwunLJQrTn9c4KgJi/27Zo0X/CDsDa
PEjparK8aDFoWqIZ+ACseOl+GHII3zoP6fodaj2od3MAwZk0Vu7KYAS3pz4B
MGfcDHoTMfrJT5BM7KKNUaejD8HDtTyevE+hINAareaecD9DcdOUF8hUPQkd
zDapck/vppEFWCyYjynElYrH7eZ8ZAAWPx3QZwcs7kKdCq5bbBUII+vV56mV
Wj77X0zrZknIR0EI5N3XFkFwO+6vjFS5ROaiJbooSQyAWE+r9KkRgmiZUSnX
ipxsAapCYz66TI7vPUUjaOKsWHpm3cpIm/m4G+NVLG76heyU3+6MJfCVClGk
BDCAEm1UJIHJ4edhPv0IztfqBS/Q2Ymy7m/NiZBH7mmsKsjwXUfrLtskF7S8
DM7Km0RaF8Qd2NF5ykAT5BDU7uNDnN/qsq+uTLOwSv5C5X0OnQ/cYfXSRUM3
naLi3lTh7hF3DpPVyuZNCq0VC/rHihcuEaUYljL8pPv774FTPBciDrNhXBTY
vVOuw2dnWsUFnB29ilASZaCq6/v+qovlk1k992X9OTf1bYwz/qik+d7JHegF
RJ2fB4OlQFpKh7dt0dSJyh0l09jAw5q2Jfh0Lk8xJIkoTXId/7fREX2Ao4k/
TnXW8ZAe5YFFHJb+UWoIMa6ao+GYPPTImNdi9/IIE50kbnWPAM5DqWmuzYZq
k8c9mGRTSOAe6IlECmXdDMANVxrArcFOcO3o+QAfIeQ28MDNuKm6nR3q9ieB
NMP+y+wzHO9w8l915dJMyL4GHLOgb7F4u7KJCMtULey1KxPpT18Cg6QWGPYN
Bg4Yn9eGDZZIM0ow9RzWWBZpzr6xUisGDuyk6kiN7sNtHbl2LlDQIiWNBGBQ
sdkvjL10PQyKE5XAl6DlAcTUTFeIVyShQccBJ3sWV/nhNszxKqtuV515toXO
34bbWOjuSjLjQ36MZJEkW2VoUltBWx6/x0u3meLciP4LeLeqFF+5d5TUB9IJ
okJ8LugQXFfS2mNejB87ggjQoTSxSqwqFXEfZUibKZVfqSqfmUzO1uySmljl
43HnO5Zr8ZZroDw6wXnkQwqcBCi/DPJKp98wpjDDWl5gQPpn4JPGqF9afAxu
QPQkVlMl//4r/JKY/YqiUTy0YwpmTIDE3Qa0U1j3dJhoo9jsX4ibZJv62CCM
igZJgNJUdBFzuh3cuJa3R/IszkxfvwgkQgchCQPzlPqrPn+iuTb91o8ovm3I
l9DbqfDx+GtsFZy2rjUHe5YJm//o6Tg8HnxaKmKdRYNmxdb5R5HUCdbuoFy0
EAcokK1GUmye2fVwyImpbWqmCi1jypfaxTHQxVe166eEcdEBOqTqYrqE0VAJ
FpRRJToKJTCR6ib5RKkkN1nTKS5YpzrKXRdz6sJTWHRfkvG6a3AFsfywpDPD
0iEJOvWa4ePh3hrU9VZSTC6xX341oH8S+Ephel2zJhqkBmKZldiF/0qMFwat
NA79p3tFA/u3l+z290c9NpI9WZCW9C5p4G3qV0OvNYpUOASyBuG9KfcD8pht
/TxS1NQJdiJNgtZp6pNFIi7PvwBHq02KogbwK41nWoxbxxk6cg9fbWIBapkY
WyIh7o33eAve0r7s1VHAGwNkU0WkFSouHK0delN7lZiUjr7cZYlGUcDTplIa
yQg8k+2zxEi+0I1WGLKllKr7Igw8J9ZTPLspFB/wleDRqhho4KCmFn0GWLsc
ETbdyQv1S65KOWS+w+XdeX6Lljx75B4U7uXpv8cBj9V3FE4OA8u9H+NCHxiV
/asqdJiMWIyoPJKy5/CJOc2feZ9S/mqC83CCIYv6MpeLCdPkBQNSkM+3W30b
FIRKK3vWvwpbT2RqBSgt4QYe3t7rF0++wTqEfL5qgcydELPpcloCBmbqrxHu
IJ06BhEolecF3cM3AEqbKiVpcwmhmBtc8tJxmpFZRu8H7Umx0qKDdbGmX6bG
cAzJBNwlxd9SxjVZnGvvHJkWR9YoJrZ2VxSbk8/TVSE4btdcv0nRIeePEWpE
LwMMd82G/k8/ENNLRZI7f2C5MX3dROyouAqQDRPs650/BcQQ3UgiYboNBJH/
n0s8o/0vyL4OSx93vtl6/0XNQ9sIU/OJD5FoGHpNJbRu211XYTVRLrRDAd/8
ddg1qcBxL2L+gc559PItOPbIXjB2lFjSjASPQ8WCDgsf5VIJnwJ3fSn2jKCa
H5S1gxV63GI5Uljkk59TX8H1zcVOUL6xPEUzkf8BD0MpMru1SwAXtTQaQFfo
t/8CyJC9rAwIWjnKgle0n2S4IJeZzOWyrjhwyGEdzw+ch1ffJvHHn5Pa7rOJ
pu8U9LaoZYxP/SAK1nqhOqhaSXikESrzfNXH1iZOgrliXfcUoh+46f/GHdhv
ci2DTk/UBNDUwKWhEgTN5zdoJkOcW2JwOaremAQMytiXBxjv8xyLdx3hmYTA
Ewkk5SgRuSSS430a3Kg0HhHk02pXUkNApY9TEcAzm+XkgZ8mvLn1l4o43F8z
UoHT2+j1aJ6s7AlYEfh+jRqA1EdcVgCTlCCbYjVYz1DD62oUIK+yTA74adjv
yhafueOyi9/HU4S0YokNAT4CmLIS68/dL2JA3RXRvwVorc5QIXLjFfrLx1bv
O2z5gCIcdDMKQWbUwjseNhCtenH45RmIS5ceO/S2YSjAD0Jby9S+B8bUDJit
iP6E9cOiCZfLOM3aZPuDECqPWJzg9fb/VcyHtWlOhu2fwvFlmPlUpHT1jLrV
dstOdVSBXib542LPti9gJaOlcqPVNuuJ6CzUQTsAwMv57wvxtInm8/KxEkxr
VdRaoYJISs1eUelEy7O+OPtFA3G6TZke03Urkafe4a/XTeYAiZlfTHtwJE+V
+vVdp3yjQxttroJ1XU+8y9bjICk18uwad387p5HNMrpIUVwp/p8bJ/NmWcnU
x5GhS8ndC3GCgn9IerKOos8yOb0jVe2fYgH4NP3Ii7kJGNMwm5QZ1kCxvfdP
hI0mx6Pr0D9hRt+1z5ickJav4V0uu4wi/thkbWH7qeI9BOQEQbxvX2TiFvmx
sOwZI+6Zdny3+c+4lwvPpfCbJBkzfUD1nhEqraG57AetCD2oPFvf7eTPlUtC
jJ1XbfMFjqqxyHpoRQ9f2TKo0F6SYf/6x8PHzXYKNOfmDs3pJevpmRUMmEjk
DlOXCIMCrjbXdtf4hRdF9yzA6v7Y9zkH8P5uWjb/mxlxv+RJ4hJ1uZDqrxIx
kNBaJQdX2AdEe+ydZ1XC9H9MYfIL77K9EHFU9sjG0KYb1P//OUQn9fNcAd7I
PlPFq3O4f4tdPK4EpgNj0fkSldGR1BLftnT/PeoZPk4v68gW88eNAkP1ijLD
TD/PjAl+vo+03eKCbzdUW8pLzCRP4pla39D88PClbMYMAaxZeY0zKXRIULym
2aTfszP/glSW14y+yBvcXmJUm9a4mrPCefJ37rPDyEfvZ1jg4N4TpAH7cGUU
M3zOKugzrdYezFfaVV39DXauc6037lONjlU85dEfgwJbMira24aTROOA9l/W
AT/lI5V9T44dIVGkfF5o+Pb/ha/5Odx3Ccrbq3zf0Jbbq6EUPA+TxnPKTxy5
GAm/7lqj7eEzqhQJXaMJ7RZ+MdeoHf3fBFLpUf5XqMNl0ArLsi25ovhv6HSN
lQHwpzakrruOuGDIz69Wev8Kjarq0iXtsAj9NqP4LdH2fuLwqBHEkK/2MRqI
lEW+FDVQTFk/qiojZNj/4Be0BOMoHx/NIzjH0jP4RJYbUyl9nbW0TkFbOCYB
zfjxheLzE4gFVkR1iwY6CmMmTtc+xo/aYJu/J/Ejbn7VxbO0JyCja4Vv/eOF
dRBACmHppgD9Z01e+6HWHEJGz5sOaNdpmkMjnBprPczc3hcZcZbCVFPBeI4b
cGgVdJEzvM/r2FHQsVt3rd1KPwbtzxub3YqCRcYzCyXHY2J2wUrTfRRAMxqt
smNT9toMQGOAiAwoIiYvIXt0qowMl6GbFF9e4rS4S0nw3ea8BvBabj2jJE7i
z5jvGz38a9PnXXNGAsRLsRY5nJmzilLut2smYyIqb8XUYDjRr93PjqdkpsvV
LrexAkbffD8RSnaNZWouNml2iFvULqC5B+gdnKcu8WKZ0AlbQWiUCapk9Zol
tosQphj2i25QM4h+m6JCd3zNpGQcUxpfCkLvqcw2SfGaIpI5W5pmg8nHG9WL
Fnb7nR5S+Bf2Nj8J3O21bGji8xkvQTcWBYRsSLViofH4cN5xGQP7QnOUYJgB
Tac7RKr3Pxz87kYqssg7CJaqSzM1iGgICXLODogstAAVpFpNqEI4sEK/DeYA
gSfGD4hX9+g1QGbEY/TLbrRf0zQSQkSh0PicUp0j3bSo4UJ9/xlfBzXI1f2G
p7oqcLsGC0nLqzBr8MV/YYDsThpXarMhctL0EXY66cxsMpnaCLNuj6oachH6
SvNwnEIfWdui5sw9vzM6RWE4k8wE4hN7sW7xaQOVoVdGHnnJnxOJ4c4aX15S
l7afCbZKrhwQJztrCw860+rtcpAzQ8NaP3bs7QPXsx90of6HQy28oN6JDUDh
mRejzCSQR6y6FCmvFNkZ81r425hKuUDu15GVVhobAbMs182hQBQRk8eM4nFP
mCoOgDC1k5ukM1WS7OfhD6RBV1zWfveajQcImxO1kylFQaT4tTMCMN+b8k7I
HVt6BWJ624QRnqygL5sepX3y5TCUPx5RdSnW4VYfRL8pmjfHLjIf3zNyVEX7
UfCc8SesNh31Iv8Yp+WZP9VjHYTpbr+OnPGVbTmRYdqXBq2/hgQ6fK73HCYA
mWBWs1+D0mbqpF5Bycub/VL+Acr5AAm6WkbIQuucYDbvZ/z11rNpL32T3X8l
LywizhJMTKdSuH1vLf3UF0tdsIz1EQ3+U+pRQVjohJuOjMC2mLlwtQ5r3W60
RCcZzODImRf16L9KV6pGt+g8LJingghGjawSk7uIB8+edlqocE7ljfeTRa/7
1bW39V1ftG4EgWifNE/C/epbt+e3B7KAvvterrTlcyOEtk7R2Gk4kH+/DHuX
hRjf/lyUpIA5LavMW0FvU7ruBmVHnpRj5w9mRJYTVbjYu7vm2cozimivz1GN
XHwh1+T8yFyH4GNSAvxtYe2h+xPOZSovdxyZqCvR2+XYIuJfZV16Qhotuq2B
VVm1IMpZUeISqzBtHW3fX2prkjYNnuX3kDRUBaUA5kD6+jn2+0Es0/hDXf9t
RTRkfdMj7OXzxohPItVDGJO6KB66WObC1wCRbSoN5JZzWdzJNZdXWEtM6hW0
ETkYrg2OV8yo5S4z7MFjD3NXIn2vqOe1va4uuR8KH0vuiHXapTJo7QqvSL1o
OH7pruOKT9KhGrtjtr7omJp4GgFNazmK1HnltfWLZVEu74iVZq8zGCBvh2WH
QOzgs9znc45UPDbBYR/kpdJyhEjCA6MESReKAOP98lbxdBBtow5G4a+HktcX
zNQrW55swIF11qnsrOMqLrp9Q05DJLaeQz3r41buTlHbbZygH2nyxnzuIgbb
YSAQ1D1gsC7aGurd9Ezcsu3kO8ArDz6Hj2ixBsN8QQHPmKjhZJwbbT1UC7C7
aB+jRSg9HlgKR7LPZF0JS1QMcurUWq+RFg+oMgBq9En1LVjcOZiHSCE0dfsQ
YxhD0d5qhfSueNt+UAlDwF5TcwjNmffXx98M91kkF08WQb7dzrIw7O3urCdJ
vYyhhZY9KBmbLnoq0U0M64z5UVuqZiJ1295efEjybx2rKtnBiR91qeglbP4/
2igUM0Y6tD27ju4D3uzotqnSv9+60Gx40YqHhSpdC/POlfjmS0hfpeBVUQ7A
93GH3k5xaL3AKY6ms9TxyXm6f4IpYxVs1zSPGLohoBECol9P9J8gtaIbeYF4
nOXIyUyhAUBfTioBPxJyHOsLJYO1SnxYD3EW8js3w7dGkqXGKN12lKuNX8g9
/HADfaCDV5nnkYW9DKh2s4wZwJVwQOpHiwLWg0X0w2Ro01+B023a3nz87jVw
T3JIphetSq/gXplxyV0F6CY3/Mxgvdu7SW77vnXNjqOoVzzHPvgKaBKr1RvJ
x6aHMuN6wLYsTURFXqe1Z23hABUWqKU1JYSRexXLZV7fEnAeBtJ+pwBc4XKM
vRbNPn88AG6mkY5hdtJjuc6nXe++kMIpYQPEMGMfaY1GopgCXcYmitqu51CG
IDMLAcskVvysoKMcSL8XN0Xqul0O6I72jorZdsPtwxax5u1nfWMO95NuGrAG
Zt2VAm+ZrrcGtIoRKRcIaYr59QseGL1nlRuCskMuSMYm3nV28caziggPtfS2
acDOy4CRDUN/0lO4VTUs8j8S1HbQIDrjgYznp/l9GyUu6Xlr4kEcXLiVa1WZ
gpLVmjhsqoLdZE+a7pePaV1XwPQWfAGWMpVnZsoEPjqmMfC247UFSsyFlzp2
5/GgHM5hTKu4+LB7GsOJOcF7RU/RiBeZo7SNrXLT2bb5lPZ3MmbHt00lhZzA
Z1h4phn24CjJz1hvdG5r6676qlQfXziMbE2GF+vzfkTuPZGMDeE+lJ8KwZqr
aCNdZew0C2EGM/sHGKjglEByzelqRK+q7MM6GEVYMguwPxotgKxwB5ueGEHD
tgQTNWYqhAOfJRDl7BgcuHSfAHOdKHig/lCX9jKdEdSDEReHLbAY1wm1wsSk
uCeLgzm1Hqd3SD4qHUAiGHNcMvPLKgptvtdXo/xGU2B0tqgs1+Zr/kItv8Cd
Jc6RR5V3p8ghF3PCW99np5PS+K1D/lRZqv6X00QskjUaxipGoVbDUpL4aRsX
6znWQVr7cI6PmCNyGu2/26yb6AV4Ju2LQ6HvOaiBdoEatFYswadFkJjba8vq
p/5cwTYUciA7IFeKyxqaO2eHu7BM2/tYXsAFk2k67mjdtT0OAB7Au3/GeX6k
JoPmfyk439f8y7fk7GvRCKEvJudqxaTfWKxOEuA0Zjkuq8GBqjTM7lJmD/zm
1Zj7RJrF8g+uMzMCEyIV/7GtuuhVr0ptcH2/NlW4itxWZ1ZRtRWroMROU52m
HkJPxpMJpeyWcIR190QhEeyygD3bRMsC7VDSNaC4/NdCw88fjHRDllqJ0mWs
H+YiTSte1lzUt5iExIL5oBZHDQjSasUuCFA0fzIYbPLN6hZfNDtvguCTkIwl
C0LTSB/WN9oXTzG6As2Czc5ckQnSL4QMXEbD8svn1pp/bXDrVIHFE7q9CpZ4
gDVPpMS0QdUHfkQNiGwCapLsgjAAj1OHy35LAMgXqr4ix/NTu90+/LqaKrFj
A2IVl2URCfIMW7fDg0GcBk7J3e4H7dhgwj8xA1nw8GrpRGXqRxyJRoG589Ue
ndpq2H/Yoam+xEsopADluw74ugAB67a4LMnochexyEuoJenFOAnrU2SvlBTz
16c+2VcVpAz9pzpg/40EWF0UKmRZqSF6EsAWBCMqUA0KK9AZtSkGZoaIs6DB
mzPB6OasZueAQneaUk1mALAVj+AAVcGLkvq8LQI3UGSGawGPS7/P+PRp+O3b
NIFUc8+llIMS3YtWUMbvhGX1VdXUczKOxkp0nkaX/npvz8rYBjLntVf/FfDp
M/ChBRPEWN75pN90SEyP25hnJl9qxEIzkcN13IrfyqlBnQrdlf7gq9sB8Nu4
MsxwTQK8AGtpEgQahTySqjQ0fvuzjIQboFmnmRM9IMVqSK2kQk3PBN5ikY6l
4zDawRNyjriWv9Zhpnbe75Ud7epgu2kPJ046hFW4hIIFnnhqhIeVEzfm688a
B+d585WSGsU8A4l/hhZVi8c+pgDZV9lqm/1jxPMkepWN0Jm0iNEiSi/othDy
DLCZVyEBJpkQIasJL95GjeBQQUttkMaijYyiUTMm+oA5fCSDEdICOWZTN3h3
NIX986vvfryZyroKkDgll4rXyHlyf6XoDLuUBXJ/Ri4DZ43Q4OOoIlrbzEMj
k0sCqDBquIkmg2kVJXrCXy+nJFrckuiiArDndUVyLQ80gXocQpj+dK6RBvep
4Kg4n24VycWLGyY5FuLPqCqw2mKWAmtmBBbwlHuAc9cebImga9NZywlSl3d8
xsdwp45rTk7yNKKIT3HKHr7sE4haFKKKEOsnljjJGurEgM+WW9gjDunLYNPp
084Cf6I/wrUhdl2shDJU12+DPrAfDlauaGIXJ8hMSAil2n+sW86kDhqtxoYq
rBLk8WWH+vsek9mqwlN7AHMuAoudvvf6krZuAlhJs8m+dMT66oGBjg5KDy/p
bQFJPwPjdK5Nzmzek/4txhge/+xPyJZb+Pk6t7f45w4nAOv6NbHOb/KDveno
lbsouYU4Vlsp0JRz7DyDCVXPI8D0FRH9HxYADmhlcCTh81G4m+h0wkPMDoAz
73+w1wLehm8wpf0N3WeV41sxigJPKTV8t8Krz8assoveYCJrxjpc1VaijVgu
8+9BddXLlfMc1o2a+XEfp282SYrph+JbF5xjdK5rbQkdAEzL+HoBGD/HUb7u
v9unJt0qhcQwQ7gnZFZFUS/a8UElhYtDgwnYeeF4GvcLasPE/PMfRMLAYrWn
r2fh9qrkBaE8YQWiH9xhsSKI+RpwzUr2fgaZBxw3Zexta2Iv4+yTqhXChYn/
td0kAjCPoyPVVVQnyfcwacJe8Z46CQnjj3K+jTkTaS+eVQocWgmahemJzM1u
ZP2+A1fPnnKzhs+MJDbAIcnW5rzuWT9AIo2ZqWZotwJ01ZqSzsK7N7OQs+99
9m93kcWR17ocCmNYPK63rsWMwWa0j4M6Zf/KfrUuEILAruM4Lh7jisli6xVG
XGip/n5EjhK2F3ekrL176QKR9GB3M6ddZme4x7XqsLEcTm2E2w3Bf6CyyHFK
CtkG0k5g2s5qnM+XEGhy2VPLk/qAtPI3C6prS7kD4zZRjTjlTKKuXi5pJ0Dk
GUNoFSjxZPv/NyWQ6v6asvFaSvw6YMd1ABDngzGIKFcnhmLgqNTCWe5xO4VN
2MOV8tKuP28aKOMmfJ3C1gDbpin8e5XLw787W05guTkJbB0CrLrzS0f1H/45
sYUSbSpPoE5bBqLh+k6hOqCXlPBec94V+8LXeixwlnpmr2Rg1cf8N3a1T7Gt
mcTZo8DRt41lt9afQZk+GLTLD9THE4sLaf0C879bLAe1m27ckPq3HOoMCLlG
En3x1qP0ss/JRzegPfhmAkDrnga0ZAM0CyxrcLNZ9gzfOkEazrzB70uySTFj
zkCnkoMls0kAb+LZ6x6+hQxNGmqP6P4AuuFsL0sRurIt4LRs9owZ5CowZSYT
md3GJ0i5mrgz31bdiB6Qm24UKkRasXTvlAVn2UCb7Y9OlI7wHZDzMzAsfttr
Cdf9WvtbaAn9r/plDm4u39rEW4oMzseiozYO/yR+h9Gj+t2D7/No6HOmd/ks
s0Dade6hUR8nLgBUZHDo3UGVyexJLC/bik3CJ23+ZU72v2QDfoVDaaeyk/Gc
LOFwvrdaaNLXn82QynAKPL1aVRaWKyhydrupS8itqSybxScd2kiiqwomTTTC
zxQjchZiY/rz5o22XgFAM92wrP8TRW3fVDdNZRq00tfCU1IPXlZqi4BnMlBz
FAwFLPDJAuFO74kB40xcmgkpnywTryiR02Mf63U9AHgd1gQx0D6A3ZCPJiYP
n4hvUm2LnoB9UWH9U53DzQLC184vPXO/eGpX30TbrjkWCRmefvsV49CEhach
L2lVqCI5mr58mLW8M7Xw0ClD4N7Dl4p68L8eFM7dLX8i+0OFAPAkWE4jzD3P
fnBt5MH9LQKvyiNHDJ8fgR8oDmaAtalxuLWyeoR8ioooGpiYiOxfyOKRIH5z
Jk6fW39DLJ/LoZllhrwfyEBteQQ8vxRyZNjd/L2IIMoe9ptP1l4B13R3oIz0
2/zhv/3FqjbAkZAQ50eItfEMuAD9IJDGiHPR8wfU72KEsRR2FRB8YNqWJBhq
/Nt3/5RWpKYJdGM/P4QUCq/jODwT3rIi4mgcRmMtD/dElkPo+5AiyViIYGEY
ydHOw9obWXtzKGkg4ZWzTRoI+p9Lyi+bv0g9IC4aXtpLcC5vsQeAOTyq2WyN
XOywlVl4WIZSY1lkYHqVaDaZmROJK+gzwm/ef+b9jvATWnJb8+YBZqh6hdx9
TC6WtGCIAuarPrha+hZ0ZZn7G1XBhxE9fpeQW6EZNIVSlyfEfjbhDJJv0hNV
pRIxBBuo5OF9dcCn4R7LBNndKVaQDd+uzfvoDCdstpHZiDiHFz1lmxRrOGmq
VcZwrTtmeOoIjapHrFFb2FgIil7EPtWJCb0FB4wvzHMrGWcsl/YANTDl6lQc
YNKXdv9Eq3L/s+nozBuaTBK+AfTC6TEUEcxdAFqZL2jvoyNqGzxtwwUj1lkW
4Y8lBtTV0ETr8PkG83LFuhg1fKTsIz1O0i8eh8fhMJa7w4bMtcRy7yLE/1p9
kHVTwTNXw14680FIDYdUdvf5H8Cq7S8dQSvVaiBw30NQa8n7KUdrS7a3f9RA
KVMXBPEOxiyjpzh/1dmW0HLxe62wwCnhcAWncQQiclnXI++JrG15nJSLkXhF
qzvVwksh7WYJk6gJYlgtTaXRdQFCM/5MBvCzcC3m1tJOBmmsx80tFoOzkNgN
mrIg78rFAU6B05wshOJoOOZkayZKOHT3YDAvFH4AUng8F0TZHd+mCk/H0OBC
eB8LsmlAxf/F4n+X4faAGFAsKemmkU0otCF/7O2xZN8pTwhPx/RdUcYF9y7o
KU73G45PWxKayZ4ScoPWYcF8eemA4XLaKF7ONSBoH0cAkLvJlU32Fti5DfbA
RjH08tZzdhG6bfnqSUToSs90XXBSPMdD0c9afPIR+MZuoQtMmKDMDhyALup6
RKhSisks/IKmY35ULZWVW3uzTY5EnegxnT7ytDnVwX5FgZ2D59CzrVU5zx+8
kD5m9Q3X9NzNYhzSgdEWv4cXPG+B/tZE0Sjca0KOh45GWD1HXIxHO29V+DRh
SdsnvsxbqE8Yyrssd7ah0OC4Fb+r73e89L8PvG55DgesNRvHFk+rQfFF4sHC
luQse8PULWVh5YfkzvmBZtQbIfzuOfkQWTQqtBhMgMUGtLladCybqYPEzJiw
dY2EBo29YIjJ3pyhQNtjTsv7RzTJfez6kMj7HOGMfEdlZ3UEjVUirlVaz4ky
6nYm/8nPMmHxxVvAhpBvJhVkvNPqf0TtCKuBtf/JxkxC4QOHky1OQO+IImsw
fsyZds/Sp629bFrW+bS2YmdSGtXrDD6kwQ2IS1RWqgu2Gzf2+f1TiJTAQM+T
zv961EzSb8vEssIHS/xBVpmeq36IfmdFFwk0NnhfRrqAQUTq37Oc2lZ5QOmY
JpVDI3NoCiAJ2Vtra8R4FbeEXjR+cGEql6tpkH/kg5feoKeOrxkPITccIV7T
rpouZYfdk8zlzoVUoV63rEpxOmKRjzTKdEr3WJzt8qsQBFA5TeT9pLMk7ltL
aH4+vYR5mzMJr4iNieqQF2wnkClbIOHgFyt3rQxB5jXq8zau2Jb9jiAzrz6s
MHfd4/ZRVxPacLC/NbZqS3WoK+JiSoNR6VLqXNv+jS3hE32pZJvs82tFgP3p
+IeTzvjzh4Wnzdn6ysAXVmGtIGwiPRhDeEEkkEeByt5yJK2d2ubbqcC3WcWL
UgpjE1toMmXcxMbLj7RNKjsCenWzFAWEUfeiPIeKyiJbhrRDx0+JIu4L9m35
M9i0KcOMH3qU2jHzdvifmD6EIaNE0x7FdyXZQFTqICoYLRKPlfQ6pS2Y5lOE
Jns7Ud834WrtFXT2WDJXRzGBJ/nmk4MwdOUeB4GF0+tNhDga6hkWiTYwHUjV
nia6g2HV9qSg5biknuOIh+S0lbc4J5T9CSks2MGj7EhmjJKOO+myTd4MgzVp
34hvd47RHRoCsOf/grFGyurS+M5IkJUXHSD1MDBsfPVqIOsLIo/Zw2cwtQxX
Wx5YayqZ2EFbkrN8SuBNGAi2y+uZpJgVecT7XPdbxRaBLxr+CsE6lzpYBnE1
omzpjzXJdk0hRhe1INV4rE9VD7WVT9nCR9OBMYbzgMdSCGSXuPDa+RDpbYmz
SCwLeYFlF+YgeIasHhEX4uBTxbTVXcNC0sKClEVvQlZhGBp8TmXrSshZ2n9J
Yj5x2oB9uepbdjL17ddM9Pv9Yp672gYuQZEqqFd8YSy58glZIh40IP/EqI7D
t9LxfARO/TJziv4GXiuYSxRapt7BGAZ6tcRrs4mtzjr8uJPIQtnOtxEdEbQJ
GGCJRYPj0xV3n8r9B1rPfhO6txLxAEdJBSANH64wkwF1zRf1DxkcoiwLJ2ko
/OIZAvRS9F2PDi2HhpU4bgtbzAMoPDp27O71d/693ZX6MVwYYtSspguUyd5n
6kY15hwrrZDeTJJsee08jYtyQPTvLxJGgOpmQDX3jPTW0XWV3342fWMLNSVy
O74d4EBWKPtZxYUKjqYEEr73i3vv3rfIlB+jQl/W0jnW6R9vH8hrEXrdKNFw
rzwIlvEfcMYb1+hbUyQEUsoggSvQ6q5aziUwidYBw9tVS6bIaAouU2/Pd2FT
8zyshZg9LzRey3Z40IFx2GGUv4ZHeSLE4SEQPdh+stiSe87D9MjSlICAv2hT
wk+W/A9RhWVJ6/QLeFJhLmoEL7yQ3CpMpjHad/3dqjSy6RQv7xf1cv4O+zi5
jljHUm7opsrC8PBxnoh+ZaOXsrZd7N2zPovwpQWJdrJ3svddw5bkAtkb1i4a
Oc5FS0MtVeiycA/a/L6Q4BFvCzniN+Fw0IScVuaKVJIYuVgtZJHYh95OAX0k
luBebd3+VubIagDvslBv/R2f2ADeE3AJpLY4G7O5lwaOP6P6z4/r0EJvpnUi
ShDNYwXkqSoC02IXJ/SsNz6uwK213A440I9RoGPMIX+WTjuaI2s2ze27oBhg
gZres7F8Lvs1oW4Y2rqnvqtGphdGKsct6T1diUujhyrECO/7fQNJ+l/Z7g6d
IiwCUCRRI3wpRULwpPwrDeHgu2R8H87AucxVmNdXAzWDUQs8HK+ib0tFs4wE
WnEFkRZ8BuC/AjudgQOU2LFh8xe8BVOKi0WNq6NUqvqpVnFAMdeScttqx+Y5
wR8SsiZQI+OyALGow2h4+6yeHJuYtFdlbaAf4ZJlea0i8XIDnOQ/Y6yByLA6
ysH5cn9xet6J5L3sbnhOtGsbWCPAQCs40FSmkrYJvOGv1P+v5IjmFWS4Zygw
yVc+uSi5FXfJ/8P14bJyT39QHtrjdNhSYYXEqaVUOqhk2AnXkpbDfISUvCXv
SgKiTwpj60G5fEm2GCi3VohyeJg0LVg4bIhPWiiXapsMd+oKjYzEWmJ8FZzR
VlkD5Ld5uAZhFLKwGv9WwFb00F8SxBRzmT9s6AFLnqKAK3+14U63Kbh6TRgf
mUmciz1XYVTF3Sr6IBTwqMbGFgVYwpwQebiFzNlory4F9JI6Y3ujfqmBvTUq
l6n+/GGPqs0g39ROuLuY+0MkEejIt/DNRO1dedtwYHPfjcXQBSBHIG0xMHLS
HlIpl9Myc4ekN9Z3f46TBjDzsd0nUCb71cWOpUKna7Ar/SWoM858t2JCSdMp
5l0BeFl/aiJBfxZlf7rs7wmanzgqv2vC151ia+RZKMi1pQzLT3x+Xqv8r0Lh
lnyqE13ODq/CHEVPta5n2HPLhOGBRLhFKt7323kAZAQIowqFnzXEyFtIL8JE
T/XApEWEURj7q1W/oXUjYjJPyLM8hGN8HElCrCqJrIPh0IuwVtQpC/IcM3JO
Oz2j9zb+qVRF+HSz/m/EX0YhinYCdrn4o+kOwRM9qFtGE7XiKlrKn4bbqpcL
24+m3D8yF/52WywiRJacFIpwdlzEcTW6zM/wkbhpRMMoionWBZ3CiI6/6J13
wxQ5R+eVlCw3Y93V6KHpaUbA5Gw8F5gVDSz57UJEf1sZtBEaljR2IK6v5HXe
DBUTJA0P354xbT78E1gGox1JSi+JS0u6dBHJwQfYhbPqPDWWMwgrunJsO7mQ
gl43Q+q4GIttqQsFJdyY4QU4z33Qo6Ommi4Dyjm2eYKm5oV1qD6LIONOkQcd
4FswS6S5EH8b7rFAWaFL07S65QrY+yEEwvYGxe6Jv+/tZN9M+LrkXXtf6K4k
U/rucEwBB7wVyZNeP5oXTk1/Eziu0fZLFdE44bfsNH3lh/d1GRsDGavXMmCL
FDN3l8WvNdPACKsWfnVxuKxzzSG66MqlLh4eLi23hYYbdjx7Kxe9U4kH12As
GHyO5owEPtoxSaYKu8SzG803/yw8HopYoxz+BK7FOjqku2z0H/hlhnz/EYZg
T+GHy8CH5ah9dR7EW6fDgzLOQEjg0BV9PsGbN75PBzXt0zG8aeAG10oIyhda
mgeSRGvtSQTO4Z9VgjRKTPRjumQVxp35rGVGuHCikt4kf5CrUftn3DJMpyVb
xsHyOfZFVm0rBi8G3KEQnS99qfOo6mFMq/iOe+Pa1RV2VvUd0NynQ1wT0X74
MvVwusEzbPWsiFyqZ0q3IgGxaNKigHsZ2PA+UsFFVPGOtv77i93hyAre5+ht
G1bL5VDfJ1DgH/6xv8NBSiDKOkhaMF3tjs3Tj4xpgcBowrVpYpxdM7260wo7
hxA4Gl62d6EuKRE+EU+qHD1YrYDnyrJQxLMoRFxeaNB4OFkXcypu4Mx46v3s
4RO7l/vfmNTxIi6qCIcdZNIGVFWXlrpROnNUwLgv+fovW5AryiHCSmKY3Lbp
NUmEnPsTakR3pTQtTg5qBg1pelsyPIGVUrr665ECINMzJexUFsves3U5dx7o
sKI61pLA9k0btvLYH2NOozI5OXRy6c9p7o5x0xWTciXnYr9/rctH6Wn/jPcM
GOZjUL4sQWkPAjBBCwFqAPo3ECV6cKTg33ljtFFG4xMD2iGjxkbQsrNJ2DMK
5GyxklPzAS/r/Ph/AXLylGr1HaK9BwzevbLwI2Qf1ieX54bmCCM63/tBdJf1
PK2Ns6VoatMeUj2+zcpqsPL1NfeaxYOvVMU7KgPyK8ouwx9l2dY9varmGmAO
5Ni0xtU9hvzxFIHXStlolCfCSN4gQ2a/tX7Hs1zdMi8eMQfz5oSMlev0Ekxy
ehUO2moLnZgUu06XY0PtTNUnAVaRCHzJSZP2uJ/z2MJjoAiH/eumEQjqngP0
1HVxSuwjZ6u2L3lbBXfVB0mt0PnuzzzB3t40aoZ1hwWZvpjfLM+eqKEc6DLv
18EhtXPj+omgZseRLQ1v0EBvo30HBFdG5pv9wZweg5hTB7fg240uKGwk4Rld
ZdAfAotsj8OMP2xHrywDnVoswl3CyEi1rN92WUT6oF58eP/vMFZKvcUD4scB
OkgMEDyc8hCZfIOmq05mf1siFVb/j6uUfUbn+OTnRIW4PMFmh62I7k3Fzi2w
xpSeChaBQy1S8cypPPer1Cl/v2GLRpF+qqnaoI6GZeoj2krHw9GyONjm78i3
PjayFoK3Ehsf9U0UW4woO0hyX7oNORPByQ6MaGVoQNOOAc59G64CN9enUyFK
5HSKIwgQGG+K67nis7F1ffv+isBmwNruqOpasRuYcaFxAw8zHruQwkhrvIuS
IfcTzGL6LZbkHBVE0uga+vuHf4AxIcJDtFngDjTlNW41sbvEgyu+O+yt3osV
JrwNp6KulzAUzj3CwI1g0aGAoeIDJnfpdtuxzMGH204bVvRbPKrmPdxokHou
OckYZb1RpcGI2ehura2Sghk8QFHBGjgO4Dtr75VSKPZkVURbtJzBzWJCWUdY
yNjKMolEUlL/7kjtQZ8DtLRMbxsMYw8E8qiqd2RbAo7N0V5mKmYifm6Z8Ctp
glIB7Zswg1zef7lY+CC4dCC7H7SBqeNBi5dEIhfhYq4kqU0TFV7YDtYBbcZn
m7bASfs7w89hDwcikPMR4AYgdsqIJXU4Gi28vhmcCXoyCYEtpdou5lKeDMRx
X9XftWqQZhvgyNS1LAdY/OO8dAIpQTQ3CFbqablatYTgT7Fc7j4pFvbbYy38
fZKO8HWMdjGli85bW5UMm7KPsJAcWA31XX//SZW1flq4DlS/Ugv18FNJLTHS
mAVmOxc8nDPTGlDuIXJUb/k5iUkpSewOZNFUmPDYppgXCPTR68nH4Soz9Kvv
VAKX7ogYRVl7Z6O5W4Q70y1teut9luldO+j9BWojSNmlwXQFCaRAZSJoqjh9
Qlvdlhc1XhVz3+vpCFe8ggrOOVagLZVziyxGcv3DbRfjFvQB2bT5qAX83LiM
GsG1hqU+pkqowRo29hCcYs8eEQvC82B6r1tfJdi2SgHn2ahXX9nih+tEo0Jy
GZ7s7oG57WIyoFEBX2K1BUCT/QNLulgO8E+g94bWyLaM43gFIHWYH4zahAul
duVbNm1v9pg4xgZmtlIPSS/V3BGmwtv4wYfpid/ePXugMOUbY3lzhBmh3Ao1
NtjqPALdFm8UaMocO4ZNrjF1eyaWgivkksslmAxWBnCU2sB6j2i42kCgXc//
gQqAN2X7ng5fquYRG4eSKRYWNePX4AW58qpHUhIimHWoIAdnZANKDETRvcaE
35kD9NdhtyI9ql0e68XKwxwDwB9KXfmNERwURIXMzIHX2z9hDq/o9ZWsdpiv
mV2sPH5h9UGK2sJHlq8owqHsq+n162Pk7UXfbr/W/KhbNeM+N3rVlxO9fmpq
qKNHxNsJnhGYRtDTRtAkHrGr7qGL/20mpbUOyqVwwCzKqnbb0lH7WbgwIoWA
F8C5znU8AP6kNWGSY2NRNZEcURcnKqrZpHlsgEiWH7tJ8FiyUhzUuuPYTErI
dJ1CUZzXEhyIRnHWts5rrRbPLb2ioQiFTwIFeDgXaJ2JhVzquIlivnhS1CvI
IZZXi11Kcr0rNLpRIh4SVABYEwfErO8ITMFojb9Wj3EEILPORazxv48dthT6
L4IH2iloR1oixrM/IQx7uImtKzSoxToJZCLOlystGTWF4CtSmlKpZ+qq5L74
YxwtN5o+3gN+wW7syGFEcY5QFUl/Ga+e7lVVrPtXjHeZcaV6qQrtKB/PcZjB
1QgRcR8zw2jsjcJACAZlA/JvbPTGJ69IeN4DzAObB6QUiU/isldZgPlnBpvi
lEbU2geHx8GgHNWyqInz6D8ngsvgaaCSdiWHBXSi28f/tY1NFuUEzyPRbE7w
22PgvIGXmtFhfpsJ4jcJXHnN7NBlHxfLv2cqazvWh3B76HbJmdEU3wjcbx2y
B20HfQe+BSDz4aJWmuTf6xK/Esn1Jxoem04DypPmjxbt7va8JJF2L3UM4Xw8
UURLAIeuHLJ7zowX/8XEtF/IOV16yeNSkm1EKWLdoXVZRPhiujOvwV52Quj7
IdUpK4PgdKmrPHxZ6MuSrN9SK5Fl7xfzSbMOBsmKsZOlizRhb9/qPGBxAntO
g3wgtl4mkrX8X/VcR+wBcWzZ1ItjPCbf/sxcfqGHjCv/KCs84ihjJFqgWuCh
qEAG7+APeVGtgtxTQNigakiDEHLSuxI9nv4n33ITxKswLtpqutneTe+B9o8+
+lT0M6eaD6XhKm36E5cMn9apL3ugH7LPXD4YMth3BIGs94DgD4SJSAk8GLe+
TkMOxDE5swCm5fI+gM+RvqFZbAuwzLy7GK40yXm8FGWXu9d1i3E743XhDVxR
xPD8IO1zzSQz4bb7WHstNY+Zu+/wU9OtY0OKh/yjEcd4uIV1s06/vjP6pSxb
zgAndSzUW7LnZH56vE45RaWSYrbHWJDR8LG5c/0kYfW5bDJBF34Kh0CatHX1
7SWHW0htszxwe8VW/GaG7XyD2aWQYX5ssL/sbXiSAzi825Hh+ToOwdk72ePg
jWQPtXvmoQ9po704FhpecaJo6RDxA02QCyY0lCcJRgkLFChoqLDb2zrkHMmX
qJjzOP8Q+6XU7ozrFzTZ7gHcdqwGCwFtnpkltATp4BFw3tqRLAHKhr8NvQTA
LllX0enFrMvTNxFpe/mkkYZPiBEbgUcAUCg1hbkKo8NZLp2r50VlBLRfYlFe
8jrwHr+s4DIpx3ghPTWcBKpVQqWzz862465d3cjd66RclL4AuT3EDKRPhdZz
0eFjw41lXQTfygXgeiqtI2t7rVFSf+7XI9g+2hfaFIklL8KQSdBewb+LzqCH
mWsleb7cQmPuujdiEhDT3t3+WPXrOoOhyXknzX0nLQ9rAyzNcQjlozOa5xQD
5FLayQFTCIGWjdwR9jYCy/lylYu71NP8i9fJtOxJ2/AHAThR33aKqg87G69b
El2ypDbEA7EOL4cUjhTtZNY0hN1+ptyOVhJNuL93cW0lUg9URuE8RaPVaze9
XI0lCwN96kbbE7Rh+buuOWpEgLuWS4CBxh6uZVKiLWp8QcHVbKymfXmkce/L
RmpUwFRN785hXXzu4L5SAb9TJ440/Wff14RMqVAJStikSLQry0Xd0z0FFBxI
EXyK01mdX2n3O3TqpFlIPSO7wu8jPHWPmlCaGCLXCxFMwVGK/4xoIIxdutgS
3dENyogdGrazR20f2qWQRkTJzUikfGlNr56zQOk1cgOHW64TVNilxU5LyLj5
jH+i0DMdriujNw4dFG64Oc8ZJMgsnrvw1c2qx7NrYxlFK5+18/5PCW+Yxpi+
fKCWdOYFXGxrOQqmPk+yLFki0G9lppcZy6LWrmSjdlxuPl++FjO/YIpJ0EBH
BEfkpMW3ttt9Z10IMn9cG83nunPrVseBAONx3G6a6tJuFJHq0PfALSaX9Dm7
oAn849qfrKVPMfEoHTMkBYOQE1qw7nQZWGoVrdVMQj/DPCqErvfLHaNDcYiu
j6n3iEN8UeZshSpzvOvMkvw/SRJ4i6Fk4FJRvTOi8IDyvjNCsmDD/BdfGhNR
2pTikd09O6x3dc/Kjhwt9S6gvfOGUslkHzX1lIniRl2NzbxnNvAogyNJZfbP
F4K1/qA9b9D4NtL+AVBD4dQDDlhBOTV9X+hJoreh8QoOyckKK+J4zfigUqhR
sI0PEw63zexLc41tWPLMbWoiJQQlzuXInM4f/5llNhQAxnnRGmodZ30j1NMl
FMBxHpxiwyp6YwFjX1FFLsQVQQr6y2w6SO0bV0+p4JeZhGp3IoyPRkIyyKWS
h0oAZ1bbw0qE2Pl4brz5kYWLj1KNU0+4+cWMZUpEzk9x2XkANcqUNDmbdHL1
VU3zuq9KAghTGap+mWCKpVgiXN6PoB+x5twLLfUDxSbBsQe+Ti/c1QexZKuY
BN2R0ayDCEcy5Kq3rNnMl0l26iKEh7Ampbe0qCECjuCCwnQiqwyRjO/nkuEs
4cgygYa/lC6mvF1x7X06nauDdev6ajx6jSAtMQW1CR7qsrVTq/M0YKfeq5K9
l/4t1IyhItLD1pE0mNj0EFiKHZRyMPeg5t7qPqQbbwuqjLI+/K7ihOp0XWhX
33ed0U24Wf2jS5MnjpCi8oEhgnI8dmvs0w6suQkkaMEeuIF+il1isqqc7eRu
dGuDJhBszoYmP3yTuW6sloapezlFbZCPp4TWxc/LQoaDkqT+l6urtXoJs9en
SPl+oHUEw5tEf1/yQIgvNuZcyzpOlK0Euab0dSFNNMrj5q58Oeufkdns5L9U
PMgf3KtY+CI3aJqrLBpy8FSv53l/ZnUMKf/qjYgHx1RqWHQTE6YROFrZzK6I
37+Nr6S/Qb4ZlmP0rT3pB6mJmtW2wUy8y9ER/yk2L9BlyBDvwhlOyYNqwlYW
7lIElhhHvpPzn7PZ59w0oxHUk5AvahF3x+67dF+WVll/t9dR2QcKObO+s52o
J1wbx0Y+MLBL9A2m68Tm8UjFtCHYVAK0QPEczp/oEqhzpR0qnHb1JIK2NAVZ
hsKcRG7eyk4BiDHZDxuUnq7rOVQdjFLpV5GdxwSV2zKfwDhdOnEsYgZs6Qt3
lPDBvmh240X/RlshYhR5ZZVG3LhOYI3usucUBs9q2tfgMlLl+CT0DWFzHB0V
jvm5n6oUrl3c+vbQfJYSgG03ACdj4UF5ZKqwBi5Cz5lrj4m42t5BiuFZapo9
f4Ww9jZNx+OwENn6xe27NQkhCnaZhG7CMEatbAzreqUtMCXWyS34F3uxPU45
3IQQRhZ/tX0K1Bg64IhWvEWgII7Efu8kkCdCP4HjH9THae8Iun4ntjG+yDW8
RadiPwVCs6PyGHsWpv4TFxiXV5GLnuOxinnVA1wXxH5KIQ1fQ78PdvciO0GT
lgf9R4wO+ktw1pbz+DOYD12YD/+wM3GM6HZe8EmIrxc+4Dz0wy1csqXb8fkR
+IHB4HxuRLGiVTmMgqpP0DjTb17z/vWJnFrM6o0vY/QzsXX12tlukbVEsjx8
Ar0HZZB6YPqMFAFyva5CEP74APd/2exG+eaqyHWRFP/JQ05jfjfNhdEtWYTd
Tdbzybd1bi7KbC0o3ZmIWZx8yfsz/9FuUGw9uwtSKZMuO9xCBRfcGbaLnv6j
AUc40hfNba5z3PNEv56HjQyqWlO+XAVkZdsb5Cd6IEbMZ26MFOn6dKia1a1W
e2QdUBwtDjqFt49XBKvcvO4Ip3dhvAJv5SJAAoi5Lu/yoQ8qY2Eclq6AYu1N
LOpkxxuXCam29DRHVJEIcA9j+it7EeBWTc3TCpoUQ3yGVpxiEwjELyTsZ5HY
7weZBTp2Gg80P0jWF4kGsvR+3u5C8cUIkrYlmiE9d+M3njLzRVqe6awvDrrB
pRcqroZ2Vs87qaI6zGCVSa3frOWyVaHtQcFRdfGYBANwBWD6hGjqdm+J4BHq
SU1yFPxH63c2q0tCq5ZJmhlNjnyOCzjQlgvjsrgckQW6biJ2te52IVun5/Iu
bTl4xa4hpfbwZc4ll3/02u/QR+sB3jcWYOSppyR1mXxeSI3auxWFKGw5MmkN
UnoOlcEgNzfFsDHUMZjRgNlaJvmwomWlP111nzLew5d7YQg+WyqoQItWVSVr
tVr58RAGC9S8Vr601fmmCTf2kI7a12lUnRoYIgjfKTxJbmu648h1b4os2iE3
Z5fIx1TE8vQVxCjFUdoWsCvph0iCd9X62g5PNP/j4C5zDI4ZRcjSnl0UBkhp
p78mbRh0XGYJy7g6mmzKSoWuxFEdrrCnsfxUXQpkKEOaiUFB4NTPlJOKtIXy
ehtGC/2icljT+JExT4eLYBn+/5pLLEcx4Pss/0rzod5RHewjbb21cVmqdPoD
HKGOJaw8cra+BfnZ6vXR65fviG5cL0EFGjyVVJfI4M/OF7Qiu1roI6yYwGM+
bkyNVJHRy+Asicp6BrYv8gJJWcGffhQni7FPizxM7sBsFzM6kWOTihlNnIY+
VnVWpaQ4qqpcpHygexZ26Fu45ff+a/2kU8+Zv/jd9pW/5fFMps9fCRAkwAbb
5I8Pl9MMOCU4U6T1RfulycWVoeniD3lD18s5pwidVrHA0SL0vhxzY+v5IUYe
3EPn36dTTkuaf0UMMsc7/fQhljyJMlR2lh5cALiZ2zYyG6Iz4t/ffRWYAh45
ToVP26ZuTvPOOtMjHgpVGnMqBfadCcCf28ca+/Krn3Davm13gKBFxHkjiSmX
FlPQOOG32yudgQWvAEGvfywPAOvQtOSa9ZImVSr5DVm1SsC8PWw4EPr6Pzw4
Uzecbqs/h0UJYejMfZ8D70B/1wKV7WKCv2UWvNJbU1K+J/2L70r1/PNr82t5
/ZwMrU1QaOoWjyIkEum2THqoKTuvVU3qQR+smXz37haB0xLMRjE6y38KJYwJ
YbEhx83ua27xfeDBQjhaA9piyjqKUwEG5CDl3QYJaiHI7QhXLdMoLrmKa1Kf
BhuhngLJ7HgIdbuphje9mnzcEGVKeNXVm2AQvoL8x3QcntoZonJkFWTH7WU3
adhynIjh+wV1qHVA693xwW1CQbg/wBE4xWPoNyweNcBQdIJ6ISi8JmWL+lSC
aiY/l6BRhciIrZN9Dr2XFx7nIE0ZiElPLMHzKzSfMafifIvT/0S9uNQuoqFI
jWB0TUMS2KNgDjmlGCQMiHD0XTGzGl5F5oxgM0rRFFqTDedCwHXn1V+AFSY2
HpJ5kg3fjMmF64UYkLVYLensE5+MsH7Pinj8edaQ8ZflvFXlkCXrM3BBdUbV
d6GcQ3GuaSSjwdvZ+pU9Oi2GnRpL6lXypFZs5nZfvwG0DHbROkiqG78d/U4F
Ml66esBZ4kTcvS/WK2he2QpCTURu3D1CW9A4r7IApGjucb/R91wUQuX/dK3k
FpARig9b4rdsyJqUK1Ow3m2TXiqnMTCbb9AFdkVhUV3F/sVBL/jPbao9Yf/x
Y7UemHr8PGDWITwus0iSgZa/Y48TPwvgU+dSxP1NMt38YGlAyrrUuGmf5MjD
5XomTqmuVgRLFjqwk2+YBi3xFs8OsOjXYSLN5cLJPQofgauEv9jHG+yVphSe
hX/r+M5aQvkbHoTNsbJsYljA8+fR9d0Dwk8JCqMc/B1l/Uuvpx0zLS7Rvkee
S/1ZTrgI+Rvqow8vFJK8QlppkocyQIFjekRwmkIgsvzOj8DVm0uA7me/JT/C
4pGY+Xyd1D9CmCW0NWIMtwQbBqcze6HVo2HoZdVuv6Zw3lWATugSWrKStjxR
zLm9wT0VVRUsor79RXzf2bf8H79ntfSWoLCv5Zt6Y703OxqLN7+wFkAYt139
5ZlXLFznWq+HIYS8PxWxt/21iwfVwr+LV9BCG0Sb2fFL1kWQxMYp/5BF2mBO
pjmUgL+SSMuj30gAeOJie8s7LXSzlqLxszmEOG6H/v8eikVdByuu7iX3m7aH
BA0gZ7LNeA3lSsF1RP9JRVmG7kKv58rihWr7fOB4de3H3sje9iNNzvzp0GMx
L9Y5fre+lNPPrW4duhQtZIBW6ubmm4IuBVGplZWZ2FumtjOI8su6nCDgg87d
HDIPpTBVSR0nN6Y+muUSiw2CJYL0/D/+cpdZ/KtwkVI2hpDVmRJjGIyzSE0O
rFMgnRSCOfQJnZDKCCDYZNhUYHSleL5GAJSOzkQS01noiZgD+GOhTNn0K7JA
jzQmNr0hB2yHRG7RstaEyY7DjMz8YrwMyaKY225Ufm8uvNeCK27KCGMZx73T
C3rP0Gkr1cLK4ubT+GVU64FdtFvk42F4mlApXTZPxKqcDCTnXr411G1ZlhoM
Ncr8KCU9kEZoW52e9xALqJVCuHXDBi5XZUYLDDoOMebnmrRuqVPcGRhmxTcK
tnjiQh8LDnYmC5tWk02V8DyeAYSDwIy/NOX+4mCV+jzyefTLxZcVcivTCSPx
ph7GdZyM6Kh+8zDf3j5eYAIjRbtOJqkxLlbYBsohbHbA88tX7XQpkUU8jl9W
dE6IBMynVLH/IQVoskSoYR+C3uleBPcptqDOv6xPaGy9cflnPHCslRTJRinu
rxH4iuNhNOq5+Kil54yIIX+qyA+oDU5mYpFGZiRvaph18BgL+hmO3EYR0YDI
eXpQw5236zQOKKCNyJCOH+wgr5+GKFoGXkNA6063JTG8QhUBjbnJAmVCA5Qo
4kbleBal3UMqs9Bo6fA20IM4Lsv3HZGOS0I7bmO6iHYtoXCTpEGExPOcdyaf
dIjnCYegWUBbc/fKzTJKiruHBG5hQceAdrt4rPd+pXIa5hSyK/osKaMsGxdW
c2yIcE0SycrsaUSpiIUktLrpg9YwcVwOdhkERsyp5bTkGLAngG0l9jfmhwb/
a+H/LlXkAb71x/N9OfJq27RvRDCNqDVODDuAJNixSMsBndB/BwbzRW+QOkRm
yu7loR7+h9/T5kmrGOmNvOkoLN1cIBBWR5C47e9/3NOP8pPs5+xieAdTOk56
A8+zSsk2rwfLs0BMIY/4EYzaG6z/kbAq/fILwvgdC//+2beuolDVTKlVDcvm
XaaXC8ApCb/9RlLtp2haFTQYW7o6/Hdfy8BARNtdIKxwgfYLhtZWemWUig8O
6nybO9a867ba6yloKXxcZVUucCAVwvy65ILgJB2lI4YK77fn9CLgMohNKg70
i0OPcYQLRx7mhv38omoGC9wURcwIiadG7Lj0vgDWm3XGtxHR46UtYOLE2rDK
zkwao7rjH7GNyLWJJQbEZbF2ZU9I4v/cp6G/vRLEjriiE9t86jQJxmKR5AdA
nIdmggb5VDkdwOjZwlr7k70czMdVseqfUzmNtqpPxQWglR5g+7e4OF8GEB8Z
f+XPmlL1n3l8PGp3x0Dm8Nvotg7dO8c69Ssjra6AAnHNHFsh3VFcUmmUZJ41
2e+pVp4k1z8EPqBl/VOGwF3zZHU1fMQbbRyStGq06PFQ7iz4q7F8IHfuic48
VmyG/UFDxAmq2VXpd7gVQENPVVA/omh+NnZ97i7x1oKT8BZf07JzwLollgRi
SC59IG45ChBLlNN7/OW8AoSAzwcpgYl939hgbfKgQUdBQm/DAXF75baAyIjh
y5yBfv5wg7X0s+EUdutht8GXhs6IYDu050a8RtE4/lWg6JvyfAG99f/gBRte
XgNi9xT8Z7wTBDpF7yplUipgJXbPhl5052cvGkEqqLBvsDP0jskAJzTFo/4y
GmjzuJ2/4abbdIg4ZBEEkH7gcbr+67f1ng6OqC1LGc7/5zxVI+uqh2ZA2wGx
GGHT/sUN3XejwzwHpmaKI5XmldP3VjhWSQpG9Mki0VVYprWp0CORkIAcp3F1
VPegOCZi+pmhgysfmORG9ouwYlFPig6/vzNSmWMubtGWGSzj2vQeQIWm5bo7
eqBxE1FygOqe/AwwZVRH754mdUoRDzIBnQyUZXa3sytVhXBzdEUvs669oW+Z
R4xeY1cnPoci/03cM5J9p6JOQKXRo0vlJUoDg5m966NpgcKbUrcDAKzxS/9/
DdeCCVM9/FjhqquAcGXuZCc9210jtNHlp9Fn5v2cIfgZc/xoh2VWOLsKszA1
t94vcE9+mKFSM23Qbx6x4ddseJYRf5plJe30zxQLdAanHTAzHiv2Xi73cC4Y
EORFw2xUvbZQtq1sNU2jjOty4EOdLEI58DXZ6nist8Q/oFx7+XP9yMchj184
ijpY3fBCaH35i4+xZZCLsLLPuUA4Al+DFVvgqBPULbFb89MZInSg0OtCsWim
nom0pMBxHqssPrPvvWUKH1WXUzsQkd+Tm9lGTFv91xvrLT25ybeIkWXi2B/c
Crx2vF/QpIVsoLofu3yx/UkzlG+TgjnnF9vGWkWix3dSq2dmKvK+1Np3y2lE
Xs7kYrh5UA+AfcVQHNtKnr5x4fCH523N7IT9VsluCKUMn24gzerjjbbdzjWh
jh8C9IOmk4mN09+01t3dzd03dzh4Vw6VFdnvihAtKXns/qQTnDGloQJzmMoZ
8PWKhLpMT0/3UT8w2cAlaGSejM0YzIbAvJ0E3zOLhvpFq0N0NfBcxHGP66BQ
EAs4Iw0tRw4VEjhPHEYxYJCFWUC4KZLUVjBCPvOlPtuvoNdKsRi+8reRaOWs
B0+STpYE94PoI7vKsyxjSoRujEfu38Ce+B8/SJ080rWnCgYRK4msRpGKZIWP
I1btOKC8U4oKXSZK+2cLsViOH+BJZiDFegxD90bLkWvIdsdA8yy3DROdFrey
yIws8grQrc4cfWr52xSG9x9pWJTYCsJTGIJMhsj8x7JD+8i0PY7A0lD7Js4a
pzH3HUFohlMr3KlgD6cE+dXiQNM4l3ZkpcKuNi5ys9m4ia6ZwkLL02I6W1nK
DiRI842gjcDMQohzqoNfr1bxpS0TM2iuKx2+jJlX42bsBHeeJIUfJXjC2K53
7rQdewq1w3S3EgevRCGgqUv8D642Cq/JcuU1EA/qyGFioBViWYL1EDyNQ8Tb
jWi5pZWWeDkXcqZ6ALCuAoEgJx67UvRqxqs79MhkG5XZdJZhGI7ojrDvtgHP
p53mH80XexkdqoulmbLIlMhi+fyxJyBT/byRKUl36lN2SaYDLgWmBhD6efqj
pLB/Xis/YrJNatVE1+jWFiBjP3/+Hm3j4556Je4UIpKL5+x5Ukb9Zq+xKK5P
7XYsFUDRBAbxM5f4O3ArpAiU7MKT3tWNnLN9SWhKIUKBWO5P+QK/edtr8owK
fbzpMnKoaviCUiHGZptBCqCTjeWqY12XZEccCB/sIC+/x7eKFGA8i145bHJI
3tCYYks4Ni/QwofvPqbHBenseMFu84zMayAPnnJza8cRQQqf2K3BtPsN7FoL
q1K2aU2xyY9VMcwLkMwd/9i7Tl/vBBTju32YLWYbmfpsUzXLxH9zmCmLP5Sd
DLA51VqwX9XRwHgRDlXgb8uSRxCZR811DxFnXz+h+GORpxF4pOp6jj2mtw7D
z6/jSRnA8Ujg3OJw95KEkWTDqF9o25yzQe6mXCjw8rg6HX/APSCOxtwTZ1KR
2B/RGeoFgge+uaG/mmevcOGOU1mhSGukTtwhPIKXP1syhqeOoai0mbvUPSez
46IGFUfj9QhE5kiYq5cHYaEvXQtE8JnuLcavODJahhRX2srQE2mu5fNRa6bO
2T4VTdNi1/eEuHSi5GDgMlC37S6gDoC1neEN+lw8T88sXdvgpedxfUNHTSoh
3ZjfOcca+TZ4I+Gw7/+0tQfLtcUkxTcLCbBiLSv0/HxSwUOgzxsiOpdE2hqA
gnsB9ymvy6UnG3oQueg1ZhqHwandihNL8j23XcsPJUWVQvqX+rcPq4ViQvbW
YErr9k3ZgKI/IPZKoVVGdIq8vZu8Wvtzed+NEZdeBzwd91E3mo5fcSdU2nqD
QZ9jaGuhSI+yR6D4ZUX7phQeHI1YSQgEbO3t1VLq8krSUJysJ94CPheAOBVT
f61FCSEbLw8r63OJVHEkeMVtagXWemAu5+SrH876McVZGhPHdM1pgmrpYuGP
R9Hjcw2tRByhhPJ25SaeDcMV8rP6IQRlBS5QnPs1NO6y0zoG11QW2dBg3SHq
+oTK7DcXPevRZtyR8y70+YIjezH5vbJQY8E4Fofg6yaeGIAS1uHbdynKthb4
uferU/MTVa4lyMehUMvhtD+EHyzIj4Ym1s8S/tfuR93wf+k0vZw6TMMhrAHR
MylcEfKgtuf47X+rOm9alhVJcYNjEJzOI5INe4gHf6MrmRfBpQV0afsLXNNf
bqpW85yo/VlP4e0BeCupX30oENuKLGR8CKmNyzTUpRL5X0iutI2ty0f+JXJ4
9e3YVzfGnn9sx/YPZIA/zHh4j0WByuDK5izWb6O814ifFNYVJj18RJqwcY0s
oOL1mHVMRgIFmQJ5wEOZi7xDWez0/tZbbohNjraOgi2QWXnYHnIcALOrmFKe
7XgsYWgINLDGN87j7gbUyg8wYOBrBJblGw7//4m1apY13E3AdKv1aq7s5mMt
QET0/S0A7P/HcNVS2aqje+fgx3+0vzERN+NVdapKADbOscyh0MujkkB7sIQN
je1ycpGiJ52alaaAMlSU0y3m2CU+3YugKlz0wEJvUAodACxO/y2vq41v3Fg9
M/hckElPUnB6+v0A5cani4Lc2POUSJ9pGd9SAsnlxct+wAAel8ahuAhuvv8y
q4PULeqEEf/X8Bk9IzyPlT6Ug99oblvCi2zC3l8E3ReKOZ2lcyrWQ1pnR9OT
Z+diq5vf4daWEVLnUqrPj4wZyFUiFLG69MCk/X4sz4Yt1QAIc3+wU0wIb5bk
iT5B+UtZ2xCO7GUu9bKIZCNlzGCiBm94c/tDsAMwIuvTT1o5zWsGFPMQRfeZ
Hd08AXOi1PSSyLqO+KJ5dPK8FGzy8YGrxz+wlKv56mgEQ0O1Jam4Ty4P9Ok0
wFRVYFuWN2XzmgI5hLN4GK226ybGIRY1NjwqeBm6CK92nUrwWIP5FLX+dDbS
RDFLV5lEFuODVXwUMNiLIrz9Kq6oDM+SBPmrkkbUc7Gt3tz3xa2EMeKYayWA
EMeIWbKXpMy/b8iOgajKH7XOEdb6EFAd8u8YwATO4NgsDh58J1/d9COW2bPH
Ut/Lugef6/J+/Cjpj8HDsCKRZoml7+kemqSgfnn9uU6xfg0YH1M6t2veytym
DDd1EYyV2m4AoERHkwHBWmqI8oOWmC+DoWOYJwheDnDjpqvWdTfqUdkTZwhU
vv+QGnhJV8kC6971v4FabPWh17JAXdh+MadgRAwbv5KZLHlxocn/WgrI6XZa
ctCDNkBwNkNaRe0+sbxFJI0pO2/nyyuuIh7BOi2Rh3Wy2SlOhcpK2RVjIoMY
5euYwWLSKiwJJg/Ofl6KoqsKgSKy5DEfdwhB+fSFdFEcQ4MdZ/hQy5iPHqcV
mWdImH5wOLtglqDS4i+2G6a+vyv4WUOtcG1df/kla4pT+16p4CCdCwFxTeCG
ZPuMYp9oME/1BWv3kJS58ocxQ9IFYN67wF/0CyYm+mMAGUtOrFfrXl4bjM1H
+2BaWjGDwagSbTooT9rJg/osKjVqiXB9xf3t9YFE5GSJIKb/GwJAJET8cerT
inaQPBNh99gAfT74TobhjjSm/mqMJAnAH7a/tduArd4bTD06g1fytBdYJUHm
eTbb70RJOS1xdhSFO586Cl1rw2vQcs9EgSg3uln8+KW4ww3z/vz/lZ5ew9aD
0wd1rXppC/6KR8wMooN0EduR+LCGK6mZnfyoYJcT0ls517fMUffglH1LEopF
kcUG92hfdgfeVmJ7zty++sPiGSeP612xyoyWYZ0RsHj2MqdMBkYdgTbPXBgD
6VmkWp+fNzgQbkpXX8dfTZhueqDVGQfKKTQWTHuyzqzuiuALKtIxEs0ZxUmt
2k+7AdLnecR9/8q9N23gKeYzFHsUAALRvSQ0GN8yCPjMQo1K8HBVIQECvF6V
lrIYD2Nx3w8y8pFwc2Nld7MKwfg6NUd2ni5p0AmIfZnNTc/PRMJxhFMsjQTl
Q6cDMkXyTnqzdX9bLPsWc5tcM3d8Zdgl/GTDAp+NW6wP2++ZgGD78UAjEC5e
ucBYk/gU2ZloqTOqeORVEs4LWe4RLBG2ox84UMSvkkYB8Pssg5ZrRU93daml
AjhFPtPCKrgZE5jOlFlXQRyeNrX1q9huD0cJp/QWQgzD4wmllUXLrVfefBBa
Xonh09IwrKm6Wx7nddlsRcDQ+/hi4xoFiT/6S+gub/kRKxXzaqApCCWnxKVp
/bQjmaL1oAaJeESieQV0zybcFhGd3/mNX0nflnO3+/qIJDrw3Mvd83OqZFpV
2K/PeuCxcpWy98bZm5Z30gSU3257otqdoKkB9df59wkTB6jRFGXd4MjW0LPy
VTyucmGXCEL9eKA4b/7ShOx3ErKHyVajMbm5HMTyVA86iBApDcz9BwLTUFYp
tZhXK/bi0cidDlWk9Gii1rJkn9SjQVjWUtzT0UYMbddjUluvK4zOsNsiQ7An
eMTdS1BwT/ApltQSTpqP0vGVjKuHWPwWjDdr4dYcpKsLHdG+TvqzpJv+G3CW
8+Roq9MZ8XarzeY0e8ldB9i6NfmCvo4vlS/P1iRDXWwwtEfY0GEIvP0LydbX
Bu580JqoQeiYj5DllUU0oUndOBu2cGrRve/lyiP2plEPY2bZJ3A0MaGjSsh0
Xa3zrVDNxXrmMBDRU7VFwZsNJD7MKQG5v6+j/d8xcHGjL62ASmQeJNJDarlH
aYSdR9ApggjfjIQCN8VnELMS4K4Op0LL7VRq/pHyGj/WlRx6wpfgxUCoMK6W
EdPsCUgB7m4dYv3iRe8nzPXh6i6ZQoKjRlRW4+dLbBzq/cxxGwOYVwEosp90
Knwxp0ma6xXYt14zy1OGOLDL+yNPKyEbNrExSYSMEJQEgqNTfLqcBSXLRr66
iueIKlT8c+VO1pIVXH/KCXp85kVurOj5qWBrmgjN+yqIvuWYlwx1wrqo0/6l
amqGQc7jK5sItM6/GHcen2QYQMTF79KCgvu7urue1lqceKTGxxz1Zq5Xbjrj
8Yjin0QWPvfJnch8SJVaYimL+FCCRmAd0zR15FDFPjiRClfs/XZCpx3VeTQj
dfY8OABhSYHTb+lrPRzjEDDXtKvDOpUWJyNcBVyt5S2vWBPmVo49FkeNPVFz
NIfMfuS/OE+LMvx1wK+79mfmkYYY/QTOWKCnCfERs6EFgezetj7bwVktLMmX
DSiYfpu5saQSxBdqwwkkbVq9/No1Qks7m9Z+JKoJ4Rl1cHpwHzW7mdHxmuLg
nqpbUBFwNTM8FqCs54TTtjWk0xbU9C7ofEUDNHIzXnKHyx1S4UQK4F+DZ1kV
Giuz0eIAgbujkkjlHykdUSEXmBC/taAqrKztCAL3B8FAa7GIiLPjntry1n1s
QM7H+dTVUU0T5XU8DJPPJrfvx6uGWlHtYD55MJXM2mKf9ae9PKo+ziHTdwO4
7kBg2ar2EP2Wmf/ghxW2wqPBv3oEiwkTj4jb6hWxwJQkt/HARCuKXS2wZKhV
4EbIUa167zPuFQFfcZ17CGbKJdm9Nf5j0keNudE/kK59d5k4igymx7gwiEHe
6nNSkFXNFxlLd95pOZt8vUyyS9kcSGOMeIt3vMKFgsYVFSFxTnL/5f13OcHr
umi3qhNTojuH/AzrieBiwpDDFzyM2D+GX58PRWVDeGQMfaTnF8U5AxN16TDC
XoniC1GLZZ8BJNOERf6OmHPJnOzvz/CJruH1FYL3q8lKgSRLU+hLrzGAp0U6
O6E3EpwBQDv5LscW2iN44Qas91U0MGFg6cXF2dmJ/1uueojBMhLqEcvPaAz3
v34OoJcCbKUFzfafww66OpHWr7EJawxguJMMWw3RPUL1b1q2Bfw1k7ZivO6s
mxETlg3xhAQIbI4FmVw9mvJvDJuuKPEsNC9wY/h//Uv3aHdvMBHXcB+YKCAh
aQzKWwpint9o3GPq3gjrfeJJC9Yc5rT5GT4eaJDpaegYl+o/5rvO0J5m/jb5
xq/Uf8YKtNITueEyFz1rxK5Ug+hx2El5DnELt1IF9DFn/Bs29XX96Q9EqlY8
5eg7aq2NGIVd2+kWjlQf/7Ubmpw7hsMiQ34XV5QRk7tK2o1ViWJumkLt0Bwb
iVJWikJKZgNj7Zocq+AyaxUWhU8RQNapnbtuPcaH4KbBMgaoSxn2oD+oDghK
GRlR/jT2hPkf5x5pUNULlod3nSmqKvTD8W3CVvjegFv+A7CrhvjXZPAXP3kx
uSyrSxFZd5O7g+8ksz7pd4W0s7tPwMPwcKkiZKp2JwNfSTnxDSw7yMjRoHUO
dQNck0ewAyUV52liERt274tFMHUStr+qtj374WwHD3B96d1vx7UrV71+g7nc
rxPQlVOtlsoZ5Z+V3Cyhw/gMW7xiNakwjUu9Njo2hnySs8aGAFqQLFLavjqg
4stL+VTXJpGoOqrMw7ZkIyqGRSlTsIFZkV+/ApI/rIcZSx9hAZijBpVbKnUS
d3Egj3eEAsA+HOX5fkPL4msTjK3zx2iXJ8YZjl+7iZy/cenUe0/VuGOoMwNB
+b7qZ3M/2J87amxTO+0DJrAoBrI8+tt2hnA8VyYddUVRhWaie6QPWH3ZP5Gj
bYdq/s92tXAJGKoMtswKkrNBPaEbhvArTB8GYok8XxW3HGy1lCQlqNq9qhjB
cB0HTVZGQgu+ckukE69W9W9KxlXTEp26Q6y9Gm8PDyHBdM9whFzp6jQ5OYT1
vr2lKMxxZuz0qOwuIW/QdAzD9fYHLq5hvt/XaOTeXRWjFXqn0U+5z3M+PgfN
O4qSKEioRsYxEerDC/P+ErmqmhU9iZTuJRmrbbwHmbdlh1k3LYm1Ymf9V2zt
TolYUilhSoj3LfkS63XKWVd/slEA/wl4zKhsSjQUybu3KC1uwdjoQjeExg6y
+SuZ4iMBy+NuQzVNLbjX1hhcqqc77/hDoKmOaWrI18ejSGdL4AY9fPngJ1Ge
GghEUY8vGQ584DxvAcG44EmuQsRdZtPLEITMgpOTKnNlsRW5GKEFLJ0wlm59
Y5ZUDXDAuPYMDMEiM4VVYx9VWvZNqBoyN0yYtlhgG/o/ps55XY+SQETHVonO
v9w1w3QZlDzzP7puhiuST1N2QXLjZJX4WeyGOhXesrvHk2wsRjCTmPJKpnXU
3cE683SrW9BfVxbwTwUCxlXE2Vte8JH3+toZRhqv/b126B+CnYffzD+tkXl4
t+BJ6qPEbM1v1yOHHqEnWrP21HhH3V857ngL3KmjXX2NUoxKvU9/wGvYM0gW
8x+ajN1HhsatqsG6ycLgnn5RQxPkhcsoGANlqZSAigPAJAVhzgA5tgBE2KG7
w0Jl7fN3erHfNViwR/2cwxRaz4zrMyFR8KBWMMTny7umPMmW+oRfK1rBtjBv
W97QHeBbgqHM+dv4PXkC1ciqliwydGAoiZknw0bPEGRugxrBRnyr+FOeMtZ+
+GslejbynxOL9x7YuOE9RM7xcNhHwtINr1aAoEN3s0xDbrFZa3nsRoETQ9f7
Q/xgmXI5wwTodopITVjgnNrWVkHYQUFYfvuJgiH2AveC55+xP04EusKQpE15
gYnk00YWIsW1uLZLK5CDXu9M+K8KdpimZ1now0d2hNXteLXddd7tLcIjtPVd
ierrk3mOZFScC9AdjHY4bDnjaCFCPYEBMP/XF6qtaILNJR+CUKUGcWAv02qI
WYKlmKjDY/VLEIw7ke7Ayikcle/KXh6tnR+oxdS1ofY0fzuNuW8Ksp10mvQM
otBuxi/RyqsOa0rOmyv06ODbwjBZj5bnhQd34WubeTMNmDvnz4XvGjCOoNJI
yVrW80H6YbYashLtnSPVd+YkrheNeGvWoiUzx+wQtnpV5XjH9ozpay9RipYf
tjmahcEHOf2u9JQZbaepYKBv6sNRCW2LoKYScQthkTM9FuzkEFAP/s2I5a7X
3LowAFM0L2/Htxslc/79TBCzP/cPZn8k0PK1tAzyCxJWZFrm4HPdELTevp3V
37rgtmh5NO5T1ejykEr6ibZTyDNc1rpVKBalcO4xLSCZjrNeJ2V+hJ8A7Z2e
DOc2V7ONiJ09rxatIxKIljX4j9VV8zSLkl06VsSerHOdUVKhN7jedsGIPN/u
G0pwUFjHJPSK2okSU12smUoVtMmtwd0RKe/c6IdWXgLcMcI0op7bni7Eeyj3
q/OKrzwRyfddb39w/CU/qpsQY8Tjrb9WVd8KTGcpKxdRSGetlwh4QgXpAomz
daR/kxXA0DCFySL/bWaQu7/HnoZAl/BGrGUCeK5iUnZAeeF4WLWcq3QASWti
G0t/VWpk1QxuxaEFRTQLwr9xqjw1sPHsCzQRu14Tush4J8CORDU3momXD3CN
Y12veYpqFOi8M+P38gYiaWrOsoTB92VvkIdmDXyd34WlsCKcsVWaNqf2wNmS
AnqCTkOe8L4cptDlQbmF93qA6o3CjPvCMeMjK3OlfAoPmT33Rjw4tC9Oge/b
jAjLdDQEJDexMMDLbXhLaPlQPuqqguV3//crjALJ4gnaPCDaE23qiIqnfEdB
Cqb8k3Vkpo57pPR/n7PyKYwxTrpJqy0IsDblvKQU8yl4xfbxwuuLS46QAfLK
4rocta6cZkbNFetxo5gED/uaoYZdK/p5xjjTehlL2XVCNv58uBfbfPmy0c2+
+ZkvhFgDWVpQNv0UjwHI+ttih2PmpIK1uwXU7lEa2Aa52+qZo+Qf93ouz9sX
eLglPOqXoQZpnR9wh0AcwFnuHaIfM8hGCaCCFlvhN0XzUR47WGbNyuxsqf5s
PXUmFXMsIF7aefl+RpqBD9d4J8P58gHByzeLwzVgS2CgO7SiFYEr9lcr3jUR
+1I8vUSUP71apDDOEFRxQ4kC+3c9dKkyf16IMoSk0IpjOimDdRvxG02D27Yp
HE2AE9q1DqQkrJv95xtLO6oj3Qj3y4Q5RVaJ+bZJjXFNYVLunv3ngPcJrb98
Q3YTFoA9JmVcbnsJRv8L7AtRFzwLDaY7LDD+ZMpgofTDhiVq6kb6zsv/4lXi
8q5mKnXdzIZuO0zxULFsIHypfYqKnenqcE+eYoOIzec6GezLCyS6NtD2/30m
Ccml5nPfNjRrOt0dxDB9Kx0r2QsfE8cgdJmqUBYSs7u5wM0iNVNPcOgnKkDf
4SN4Br51Aw/m/JCaMmfC2WLNTzmymLD8HjUpB+sTwkiUsfVeL1ysQzI4wq6q
BWFjCv2MivFpuQSDLY8pKSGMuVa9bXfcqO6BQ+85BxeITHDkjBX9R6RjrNLS
vwRGyANPWJWfTlhqMVFbWIhjQI1QtNfYs5LvY3wpk4iD1/l6Hay7ordcABzJ
hRZsVVoA/x6Ypk8lOkExjuoY1DyPfAwJtV9arUQSbrZ6dt/F+WfszBaDe0Yv
WQsCYjOdKQRCd43yvo6ohCNqajdGpl1y1T3zaskWFBpTQpkOLVmgr9l6GeVr
wuHwwhHEH7ZsAPCIzTfu6benX0AB9pLI1qm41r9YkCr9GlWOCev9RhcUco/H
OaCFjlRMtacYXRZTMx0I5NLOJ269RODKzVnYaQyHkUM64phqDYS3LXSQwi8X
LO8xAs8yiCB/1zWh8WNCGHnzu8sr1vWH7y1d5K4Z2Go6xUCkzKUW2AJ7GI5x
j3PZ9aJHoN2gzksLTJPu6tZsd+Y2k7Sw7dJrpybh6tYZPlOAEeC56VIwLXLH
tg8dLmF9JTLLG+Cs33eNGG7Aa7LobUvWKi0i9lGynz7eD5zoAnklUpM0Xejp
oRi89vJU3U7GAX/mQHrYCLY9Df1IL3zRT3Hh3mvMJfdszjHEVwHntbBV14La
BEIu/sgZST+brI8GM8ivbBvLTIrtR77v0kheMT2FUP4PfNKg8GegLJ0w435d
wzRUJtzNOhmhrAxbwvbWN4Crw+6SI901QX69zPmcvXKfDkPNRCuKIZNkvJ9T
d3E9b4dDEAk1an3e836Q1sxSO6iAblECT9+xiXOUjsqXe+YSeLTf7bdpKWxW
3KL1TWClFXsBLFEgsQ7XgBywOqMGeOTJD0vxdIY0jfYardK/7KOVe6rJZDkL
BNQfPUuHKHfVXeThkw6Y+y1bYb6qg9LOxoOaJHCh4vOYHjf1A99K4+Mi4AgO
AM9F8dHzbDvzgRgIgZVrNqH1X+daG8sfsKRgVSxf8iapUiRbX3JjYGYzDcaU
9dAlJBs7YMmt8HjkQP13f6wMYWZvpUJnyHcHf8Fqfm6ABGcH45V9jrMy2f3d
5xQuAdom+j2jGzWvXDSwyCRtepyI+zSYJBg2R0fhIiclOJmSaypsI9qE/0QA
ulNVBN+sz7lJ9JFhBplFpacTdRVCfeiC7DZtW420LVo4tJsR54LnZxxsX49n
jyrHIwZooa/JCybmVww0UqKrrGGRUj+dgW3Pyqvos3u9BQClmAF0G1yg1uuF
Fjc27uhh5GpjP8HFMJzAeCaP2mA9oC0EUWqsDGWFtFwvm8eI9x6XnPfY5YL2
mNgQuQiHTO/k9mHAsC1DqY7NkhnuVkVeUHiSSTNNrUd13SIYIiYPjTqwpw0b
1V7dPI7ycOuLldqxHqTGOgw+GZMeFaZGrkQBqTpzJVt8AX+SuSZUV7SAa7E9
z67/VDQFavC6aWynbYfkBBUbET1yTkm5Fz5cfAHhM0j10EvCcWKZXl0Lgd8N
jha9bUwO+5rcw5d0Xe+BXg3FalljikfjxBmoZfrpJwcal8rOj/oUlpsAvJtQ
ESQfqEbxwY8FmJJJBqwHqzXvaSPDogzJo5knVhyBjEoe3Garr+qtIFxNyHSM
8Dt9WrhUyxU8sQgccxlaAl0nmDTBi9f1bhgzI0WxEBLE8kJpPzhJOTzeHYUf
otkOsBPUmV2vaj3wxie93N3N+GEcmKQWgzYYV2qC6CiKo/RGyA8RxZwW9pp5
8ZIUulBrleLmfUVzgMYmRQVvBl05QC83Ba5nFrAg+J0tx1sB8OBD1yC4Ebdp
UF5n62d3VB7Lq2MztpLkC2rDIW81H37P2B3OHrfgc4H5ZiHeIUyLdwMC4rLI
vJg3MDiAZirEx2nyisfJ13opQphVrQEzMogDXdY0VY/mHQ0bkIo6fd7yeMnH
1fS05HAB75C4stCEv0NRcp4BYOKA1yRAAFg5edm4zk1uyv6B3RkLx2wwzTg+
NOEuAiGOklidK8QorntQxWhqc8ed7tV7aUY7EDhBne6oNorsJ1BDiQWP056s
vNQctFnJCDTJrxG3c+wprG4HwaYcvOZWdfBiGNgMvVeHJjTNUW6rp9M9elqb
vpYBwue3IqLCBsM483IGMT0QDOdHdZSRFi4XYxiB1bcKwQDgpE27Yvor3SbA
VTcYlUUT9Plm4C2RcdNbm73hOejhh7n/fiIVyWOxYvT1SAgGNsiLv/Dqi1Tp
Fq+EamOyg32ZGGlSPXcYwl5BVNia2UedDRDkK18aezcxU9gwz1jQJTCJfbmh
eQvpiapOgDhCLzhyVC0bqcx554SD9N/ebpov7/jtAK4hXQgxBXChDWINHq13
otrVUMDPdyAr4QVtMUdk4zxHOPXkSruSQGL3oYPL34nX22nesCB3Q7eEFzd4
lBD+Vu6ZWGu0/ONblyXgqY/iL0m+kmUeMnJ5Boi4LXZmTw8ZC5OTokD/pH/9
pUqVwrqFFQI06G5WzBP0tYMY0EGo2AAtTWBQ3IFX2+mLLfttrOx78I8mFIS/
PACBspenWludBizTCMcnpBBWelLrVxnXG3bCyhIUfD5QZ9rA2tiO+VQ3hUro
l/uZxBvsbLvMNICbWLPvwG/woZVDuHJYoUPX/A5coBA6wiNw7mjnXqvl+h1b
W5ZDknmMiAAgZQKSQCX4fTMxiSlm6oDWTCpLxbFMvAQo1hXxoSPerM3hNKGi
idC/DE/zJlUUY66kLQE4SjXSYMSbnkKxjcjbnukvAP4O36CT/7mwL+FXiHxw
jc8B1NpMy2mKTLSUOxSsFJtV/9oItf/S8gdPciwtRpMv+u+XKUF2C12PO5xf
duFHSJJPUtrTIgPRTCOGLD5h3Y/tvsGa07GePt1PLiWh8O8JKr6fqNfP9UIh
kUHd5JcByiEaDo91GOEM0QQC4baRuWATd99WTzqURvJblXpPfcLcSSli7ekN
6Nc9k9aHt1UdqxC3XCnaweG3dX+7qn2eksNLlhSq9PU9zqk5Hg5CT261B7ap
mI+2mONoKFq0MufcrfZwj7UQJxM69QLDBlZmgsyI8XgH/D3k77Wi6NfQAzF8
tsVr6lqDDT4AExrxPeLMS5xNCmhP6A/pAIMwyZJGvUeDMgnxkfLaBjCHBGeP
5NZL5ZkDwts/FUJ1lIe0zT8MBhaFlCwpuFBwwyqmN+l4MZULSAF65wzh55we
NCh0zopVH95e+iF5KQyHG30MXYU8zIH4ZBNRH48Zb+BQtfMG8cUBI9gNzenl
DZVTwmn9OQWP/N6dsCmkfCifgdZghSr/wXHBKasTyRfmzSTTEsQRHzrcdPAV
xUa+Y7ddi8xRj7z5FKm30AZLpRf83+Vh143Kmnd8DdLHqzPp2iokcL4I3uCQ
Zj83iVORb53zuD8X9c8bChd6+qfevhQHiV2L+swhw8PBu6DVf6qgc2PzD5lz
pGd+rh+Ph5v0mQEqYiV3NUeRkLNDHsWeI1mw/qoyeb4+KRbGuHIH1cuIt6gJ
DrFoCP/fjv5wpdLbjlyLKST20JN91Rrb6osC4Kz0sCg3Abgr+E/Qp4Za313w
bnq7yumoQf3a3U/o4/h/0iy+lJrXxABEiaRPf4X5tC7p6kekXoniAxYDroRc
npczi+NdH/D67d3vyBIv+N3+f96T4oAfkMb7mp/6i5zX8bQG9o4m+BngvEt8
OKwMt1caJBLdZWDr7fberoNyyQnAKj+PhaP47QHLkxqeqO0P8a21llrRrtPP
WcsF6EpjMYozhC9x3jpjDMb4JXiBDdCPFCtvLRVlVBs0OL7a8Ky9JGXLL8jB
uz8xnMszaF0El2hwZe0LVNZxUKJGgrlC3KlnhozL/1zhuZBCCCNzl61M3IOZ
Qu5RqEWQFFXuNQqnSmT6zM61QjAWGOCHRDJmBc+xXW7IW44Svnq2UxoPei32
Zlq+U9Uyl+geoQTHFHOnFKBxJkK3XaANH/xJ7yd2m30PDD8n/KqDKb6aXzY5
jrygTb3J8xUZ5Y71dco8GcQdpkBDgvhxLncNfZzuFFFg6NHxlhfVqNCcHhui
+o1cLyYFHeWyxfZ/5Kb5xdUNkpiHBQ2pM8ES5cQbA4xTzGa7T9s8ufGQCT66
eOmUmBhGYwYbHLVYiDk7fsowUeQdhfvmX1JT3mlkm+8HFK0VvdnYLH/JQFhY
SfDfdnUw2Ky2T1y1u5gYYO0oa7B90nVZIsDfJ16P/NEigg+JEabP1s/7xjHv
+2GQ2xSgHRCY4jmyV+CjwbyOdLUnuG8bcjJoksJf+YAakPa6/UBMeY/RAish
xiNIl/gMsjlhpEQrQ4jIMkdmORP5woUt5YhKjlJkjEbXKHcWZu4lupKnl4h8
wi62DUwHUvrBjABNmMg5ePJFgifAwtE8D1m5Re2qN/G59tjH05L/Jdijs1p2
Rv7wtKMUY8Xmpz9UFSUAcBxeLyvNnl/dOttzxiSvTZngjIti9fVQIpqHytKu
aIEmUYzh5p8RT6N6gjpRpG1DMkqGEP9oZ9SIQRI6YizQUke2fV3yGg4NPiei
PxI6rZuBciSlR4fKVztYMfCyIHkfuM71njN9KLyIl+OGpkT/ggxfBzy3adPQ
aSIpWv4rh0UBpey9+F+Oph+mzwRbSIQW9nPKBucBTZiD36GqqLZW+BeVz45z
kSDnozScQKZk2BNeMjOq/SNClGYTsJJSslUAut7LK/rv2BQfDR51vfMWNVcE
ls0gpMDftzeqqM23di27yZAiF1lr/09CMigMJPbLh16FK2xfENiqW0ZqjXN7
GehC2bCatHQ+mrRVGlbJcd1JP39ewPm5AimazvfgPkZt5zan2ozaOaI86Sp1
6L+XUHkmnhV1jM3KSRWqr/eXNfLdq07BI4AIWpbSc35vrxJX0V+JlvgXr/fw
bs51j+bZuRdB4uft/sTGPX6Vp3HDI7QEVJGKe/JYix9CVOKvZ9eFloBKnZKn
b4EixqBylN/O72uYlo8loQIlqssoPQucdFhT41zYbLab2Ff2s8FhN6QJSsrp
hf6cm11U8Bgt9qU+h4Ty2ZhBXKLxpAKZsqjok4MwLNgAQSU7PXUBBx0y61DM
7qW9bDKdXOGP1Ycmo/U1G9U8ZtaZ3TG+xzhiielQ3nkZigkk7VsKJ+6VJUp5
k21pyVsF9WG0M2AC/cUpaND588DZyvQ8soWlUJJHpaBf9I+HNS7BZNkPvncb
JZq6epl0dvts6ikHc1u26JbY8D27bSnsq9EXw80etGHZjNj/x8IXUA7NcKR0
JQsiKj3SmJE5RTq9lrPBOWD6zqmqFV4OHRT8BllH1XvRqUaU+VP8ngZ/3GWu
4BykedKQXdxaLLedEofghG2w3NgDojDX/h5yHphFH3eg3c13C7QmEDcVs6Ga
CVk811BixkoS8x94/GlAaZhNw/m0yJ+oVXakZMQ0jecVo3DIpr29qIE7Km4B
+q7LWqFi9gFjONNAVY74GKlnGHxiStxvEpCzKLUvQ2Evb6WB7OmY+Im8cRxV
9xtoK/Tv7BIXMzinF3CYD06w9+OSveJaGsX+j7YBcEa2CIwkvWKLheQ06Vup
qoZe/4fo6uPaUpS3i/M2WJDSLsUx2QcCncVmhinspuz0NDvXrD9c3dmbOyID
ifYbQEJiLlxXoCThBIftGU+zk5mJBjWk2W/mWzapuHx80PoqqmhiNqmWe/y7
JI2NNTmMVCj8DZFrIQO6lAoVPc00Itnszbz0z0njsHXzGtd1NLA31gTaqUSs
K+6Q5fUmG5yaYKtOb0v6okzBBHknsWS6IwjTzXjvCfv7jPkENn5o8dCyFpMg
ThcmTNgTXLiXuk9UM901kYr2rkpn7h5WiNNV0KbazXXixUFW2YVyd3iOeRue
yTS9Cd4iBWI53rgvoVF0Agh0yIj5Icta+C4EKm+ZnQ9hLz4YXLsfWJ3jjjWi
vYOsvxlxGbLbSwltJddXglgx2m/YCTmx+gKDW4JkyjehfxUP1M70Ig128+vV
8XLJVxHDlYaHWxNTEhEJS1znYT5p45SRq0lAOL8CnCwcaKT5sDgYt29eKbAZ
aXDZKbL54PotU3wnZJbcVAtznkRw0bLQEQfi8o2FOBFjjCjgB6xSClqziahW
I7UrzGRxqDhzi60+MnuxLK9Q4CwAPbeujsNs2D/dEXAEGT3Nw4oH54VjdtHB
dVYZomAmpQIH9GoTLvi5D4a/0yBmyfJuHjF2omQgmAT5gH3pcAztl6t4a7JH
yx7AzIu+sCwc2YqbOgAuJRsrUOHfFI1fwkh7/iw5Ry2GA8adp1AYqadfVLL6
toeJir+I2gOek89PPd4cY+pEyBc195Cm8hTRkDK2U63LsXIDc+sqtB9jurLD
+XtiTCBzjxfCyybQ1b7h/b8+5ixONt8Q2t+jr2f5d8lCe5D9GFzDJ8N1yru3
c4rPbnop+SjjBCVkGYpiMsTURF1j5rfRWFd8RXWnlNgC3vAG2H2aA+NOIpHC
5nQK5zggivwvaEM6XIjGo/kFQa+ZqdMraPta3J6lOUAp9zpOpMdRx+duML7k
WYA/DiNep2nbLrpVO24vx/DAaXNl5JhGEwzdszFZYrAdhVDURf2g8UQ1wgQD
bPHEZuhzKUeveEBoZbapwucH8Vq7Yzd5fV8wdSV3lC4QTBSP+qJeG/RNA8pP
UpufKxcE01sqC89yVPd+37isbRAnG+amsed/Zl/g+NlGhKLOB55FgCoAHLOt
f157SZq0b6G8v3hKr7kZBHZSJcMgBRWwwoMXSQjhB5niEQ4xYSF1sOadl7bj
n7lx9Gl0R0Q2cXAzNPyGPGxrcdu0AhPWj5IHdoAFsiFic/XTBoMqyi1bEaZN
BAbY+QtZ797og6PNVaITH8GSSYynywAduuKCxQRZ9LA0ibUDTOPm/EDvhiUV
Oed4YVjO8cN1eIr+/d9emwDvYXEm0PakZ2c9pfOPFRMGx1q2MLxexRVJtMqO
ULoDyJ3DHNC6fB6iAgm5nyqOMX1mIgyFF1GPcpfad9md1+xjVruJCzb+VF/h
UIkKUxocKAXkSJprosjIo6Dl0AjGUrH0gFo5dgifnMWgbVg3wOkZn6h+kL46
wjIXuNPs1nnF6VHDur4iLpdguo6UaWsku2qAtDzInm90r4SHoeyjrMzGUl+P
YG5O3naEQrvqMJGHuTqUC7KizKTQv5CfMSkH69xk9yyI8jPHOW7Y1zfyE8tJ
IpOhVJEKM6gnwwGxYb7g4ym5nsorFrXBfKypqpQecN1N8hwZ/8SEEwNFOQEL
XHBcUSHNxl0N7T1mxfXogb5FAOKraPTjueVi7xp7GeFPrR1Rm0jB9PMifnhb
xIqai0bheYDlZmH62HXzFqfjC1M4HXdbS7Wor8MENidlNLsCC2jQKrxcIptw
2L/HKesVwUZa0KonySpX/8dFcy9rNzWx16DBlBbtoEIvjKPcM1kM6P3u3cHA
ixFOsWdVgGNwBqnEqGi7F199wuvvdHOTdm5I5qhZQuyXU/WQPwfVKO2mvcuz
tTJ+OXZygn4OkSuHsc0/2N+2akJmaBqByZY1LDAHeeZb3n2/vgbd3JooBekS
sYr8j7R/CkSkZyVJfdeNwAny96mczsr3diB+uXu9cBxv2j0foUTXxz/tCn3O
ONdWENcNDE9y1tlenBS6jM7smkMlb9zuSSA/Z06pD/svxxWPnE+T8gaXPP5s
fB8zI0QgL4Zq4c9OJjevqNJeARizvCFuXMj9MPQvbyQ+DYI3qviviOoEDdxt
Tke8tel6kiHa0s4b5KbECH+XDWiV2/OVN/G7UC2JK2nS5+DRkDNC5VLbgXKQ
rBy4k9gLbUV/qXOhiS+ovLQcsLOkSTdTYQUUrSHI9eAmpifqa4qNy3qelblZ
lgvFlShO1fLhcT/diVPb34entd4mBFaDIDVyPAhNS9qtkGCNZ9nq1XbrhVSS
t1807XKrBs7h/cyu5Dmu0dWbXVFXxgMc/LT5rDpDdOGHBTMUG76Nd1myYh3M
Q5xxPCuvn9HLJwS2y2B/30GALgfea/y4Ewbr4w39rJN0NnyDzl+EP7WyVBuK
VHQ57Bi13aFNG8qhmep3h4p56EL4YxsIvztHrH0yljQMIKneQLCm6vu70iXv
cGSR95K6TrvyBh+phD4egxin/Hb8mqoq8u4UPTA244tpHKljGYA+xoyQmXJq
JFEXvgWQsaY7SRQA+LjRpazoYPGfCMQmdHk9E8mvZsWrd60BUIoOf2dlfB42
EbtFPNHuT5Wh/KtVdi+1pEbO7tJE4Y9CGS7S435oQARJsqA89QZlW4ZJ+J05
eTw2ktHFy+qtuse9AauFP0sUlfiWcGXyX4nnAzgPydp5qT4b1p0zEzE2p04R
tKUNgXRfsqrMoS0P7M0NC66y+wJiftdQFQl3l8Er8PEB/4UrFhkzFBKjE1m4
k3KmkIB8m1PELLO8JRkzwwzv0x8ARyidS2nm+R/cRCTiVzJUNNvU6rPMwFAj
ZtY2y3HTAy2NxF1v6rSSJUywQvS5XwIHIqkHxNO8oqVD4k6drrpUgDsi96IN
/ESohCcdurcAzyF6+J78xf0gdguj01qRFhgWwwGuCaFuLVbT6+XjB99/nC5B
1uDRfJ2VZy48Hmkm5D1VFp69YsDnlQm3hYJsGS/yogIw4ceWn3GUrPPEBXxU
F1P2X4/hL9Mhz/TPBrmyWDvEQeeNHHaXad8xg7cdaxCf9dKXVOOXj4noIRsz
OyJ1To1mzs5Bc3sa1Kb2tDDbrZY9YId+h9L78U9mLgRXrTuytYhjvUoEgIzD
LV+NfME0pSHZY1PLmOru3BO0xehgN4t/+Y7wJ+kSCl/Msmb6+LuVGcwQ/7kM
CBqJ4Ch/K9c98B0TkEX2wVkDLoD8VECN0mTl2Put+6kWl1/w5DCU58Tx/rIA
g2rhhHussJBV+tk2PN8V2O3XGrxQHLUePJn+P/YPRfbZ2mI29l171hinQb68
FkuGmSyKAMU7W2JTS1waslgOm9OT04biAUfWeso+ZIM/ywIr6FkgRJG7A+cn
fwBWY+OD5rvOQJ7YP8uErVSquk+9tFcl1pX7oaZP/dnwgajLhgM74Tq3Sc6o
nSEXrVd3Rdq1Dv08S5GgvGqtaahINBt1MT1JdQ7RqgBfInXf5NlBPc5+8zAO
qKjlYxeN5RVEtYmjAf3lKhjX9m6LYWbhkCGYGpg50E0D4Kjjrvamxveadivv
Vlog59Z3p2BA2j0OCoTSHL8pmFqnK+9B9Dz942UqIObsn51ONKpBlmeLda9F
6NopgCjgnJ7qCRFrnTC2le+5stErG6bpyuFfAF4jljumSO4QbUkytC+LM/YG
SZ/Ebr97oLgZ3EV6K80UDMnW4Xdi5pDmU+FICgLRsgajrQaN6Uv/lxS8kdcH
3CddxEV3sDHbwoW+qdhrZSSB3hvCfSd3tXyrCphuaAuPctBpTAlw7ORXc2z9
RnnTPjZ7ivgaQNWxEHCcgPH2jN2inC7etWFE/gdfzcdzBevzr+4Rw7xaVAJo
I+UDfBn5OB1sMInk9DqSAZbeSKACDNXW2dNcpR1OF3usSwTet7FZTmSo3Zg7
CETNCyuvaoWfI4je3MXSwQ976bMRWwyKFr/BSU+XBgp8JHvoPBEZ7LmDheuX
qY/feNyy2pGtbe6ULRf95/G5P+1JE1XQmnAQUosheIjc95iDSn4/YkZywv2m
hMFNqDVDevKxxQagqhxQ0GX2E/Cmxio26AdJv65SkLDoi0u714BPOEqE/z22
LR+AjmjXgoz951R1uKnt4fItBFDnmii8DW96smEjU6pnojzaNVbGCyJLi0KF
UTtUAjNZNjggT019/3FVust6bL+rUzuflKhYcWIIk6a7e6SCwxPZVmSKyX6b
hnb/bn9qy0GavpRBaoEH9qSpBPr5p5T86v3hGenIUGj71+D/J6gaHi5l9cqZ
cGF/tDTS2M6Hgfc8K4FFfdM4AVuLBxQJLzBQSUpAM+oQBw55i7qpJWGZE1qG
FDMpbbBS6o4vV+Oveg8vXlbJlX1yLl3LBJb3Nr4Ost/8Y4QJaJlr2DhiMjgp
xXrXjtkyMQ7FGKyq06AC4Mgb1ZWQCUTgdDiKorQ6KmElinXSuKlXyu/Sn5GR
z/ZBD2yHdXoC+gVBkIlWh86G2d8FRo4H7oRf3qbc4yF/A+b1pgaI5UdpMu6e
MRV7bxK1cqNO/bJKLu+zzQd3fGCE+mBQf3yLQ+B29rO5d9XBMucITRL+KS+r
tVULxDo5G/b5zLitNO0rKUt0Sc8IycjtEiNonKmbwlY6Y7SSp9QK0WFhH8GM
0lD08AG3frQi/MOcTHIX66mKgR2t+gygK2djhMpe1n2zb5NiiWNspq64vmPv
BPFS3yqecWAd4eNbQ3W0ThQjmXnx6hUVtENrIdZryU7J0FT0Wi5BMYJ9eeav
3Wr+zoAjrzgVG2O7P/V661y2jri4V6Y1rNDijGV+hI5Z2Dy4bNDnskHCQypU
VSs8UB626mi+cxXRNgLTl5t+st94MCXTaXh1kQ07CszikFwzVM6ROtmPz+7y
zu0vdmWWDyRQc/yJj5595hyed/jDU/aaFEhQzpv1miEaoogGXBYthLyNtV0F
vPvcSum+PH8HjLymfczlxnBWRmXYszYlT1+L8l78ZzXCFPmwEjgfkw0Xbd/C
Q/CiuCMnoZRr6qH/c8L0OM3OpWakaW+pxMKGhdqOrXXAFczN63yKChgU5Yyo
kqGMjNedq0YPMbX2DM+BjaSBkCqUrdFpRaEOB53VjwAoZdJzTcOvBG/xkCz+
eKB7SPNPbFpyxuurSsSwWHm2Smnqzb5aqHcOZ4fJYfSDeB4xz3PizYRoMY9x
Y+F7voIKNq4dVp/49jdAMvsvzlZ4vz3z4NEVwhDwjvgJRIlyIFfVbQAJuIwk
D7oJuxZ8lmUl8v6XRwOwOJMM2IZIibsAjlU+CVOEnP3kMtTNOrlJaVDBiSjP
Ocq03MA06zSuqhF6MsTjHuCl0WWoDWwsAX7u5lBDgbhMiJjDkprLw4TpktYs
NQMTmBzLoM+6YCrJoFUeMcaD/9mwgtMzdFufcZAAjLZc9Ghm0BOYwC+klKxT
0UYNbSWZAjlnxMAaLOblYvTj471mRAGyOLJBbVX7zf+8WAQ6SBnSrCibaVqP
JwLA+VcdORFA6mu1SoGx9DrX/SlMDcVgfdwMujq9rBBPMgY7PNLWiX3LWKvC
clC59Kn/e6mVn5hWU/5d3WbP45GVvDDH2zt+nb/II1671QAK1nOxi2FMNrkv
MAruQBvRIzDaunailp7rdeAPx7AX3QP+B0nPlQWMwX4/L5FtfZb1YR8h0ah1
eq3YzgIOHQ/2ddqVc19zh7Swl62gDXUW7q/0C7pmaz6kfntGCx+TJrdXYa5r
e1GHr15fCiqR3F5BrqDKPIWmUcdQSik1KSo8jXmovbssom47vx+bZ14kH5ul
HILW2Q/s6ERw+Fw6VHJdIkV4riAOZfUVkLRSGh7WPDDf7tCTnv+WI+sw3+zY
g3MioEDtFb/tZ7jlqzWtW3+wnhbMHuLWEoblrTwNgkB4IhUST7Xmar+JBESq
/FnTCzmv4qDkdY/uNxuwV+UBG0eqbIkJlzeoarNOMFXWPliXZJAVHp5WlvxC
70h1e4ZZRlAcPeq5yyC1RA5KThuQ4JZ6HGqtwqaXUxe+duBLa/0WrAcb1lyN
W7916q1SET+/fxJU+TisktNyECMThiRfzakSFV8bGrukj/OoxVE8R53m0kMc
X9q8FIzbE5VH0AyGhTTT52j7oTvR3PgnMFZFh13z3N/RDxV4PxhKLo4uDRy1
LQR7nAnPk5xk1fkYH1/GRynA1yhk3wBZeDj7Z+VzgRrw5yVIUcMYFuDKnbxx
tHViUTe23Xk2gUT8ej0OvcIo28ZunGaGV6UNueDcO1YKkd1bQ46Sf0ACFdFP
Q+Md39REozVboJIKMCVmqq+v19YTUMuUUK4rHyeesZUDkI9hP1BQmI6Ct7TD
CB47Uo+/UAjNamG/4n+rkJVInw5YPl4rdD2i3FtLvxROWSWUklOQcsxdXtMC
EezHHi/zpkupbZiZiBkGupKqAFEpY/TnE5hEZXoI5dyU4DCtlIDgPUpYmGt8
SttndLQC1Ia3JeJww4L7FyY+1D/HJ+6vrbJbVo4N+tdVdH6K645gDidFX6LY
Ou9tegh6gthA7F+ljMkOemAgWWgvj3fYoLkIivXwbvU/E1hqfDCTLIeT5aHo
WtT5TbbLiVKc/Hy8tjASLykVWG8oUGT6BJWWQ2ZkxOWP25z0lF8R3EoXnGeP
jZnnANHfnKPaRB1GFkWFfvMnD+FYgPFMbCCKufRWJBjvgF9NhKjczSb+Ma8N
Z6+JGhEp+2DPCyKg49wfke9CjTfaJvkuOjCN5oQAmZB0EINkpLpEgmjsWp1L
MWHv23wEIwUGHtn4odQUDeiEM6j6rS6w9OJaO4s4BbJtmKu5eF3fuAKuc5BH
Y3UCcWZkfbEl8Etb+3fjhl91EGuk3jdqz/WfVXGekKvewWkDEyEu923WCS8+
mmXBUWGgP7NIrdhtaLBr0wZaBR+ALBNA8SdjtqoG58dS85sxPyY3qwhQyXfK
QM1eTxVrlLoVOhQWd1StiMd63WgswmrtaR7rTPAyonVOXdEjyDUybC+FN6Ff
L6be0DeWcFS+zKOROFuaOMf86eVlNWFB1NiU8EjxwJig9kIPrQpQMACqeR0i
SvTNHazO5h6uWzpq96IoxSUGdQmkDSnf4OgcUFRXZt5l1PIMfITV25EUQJOU
xdE0pR++mH9ivbbrk5zpJQWHr0BGiHLuipZnzQsJJj4Y9VfwUatTgQCnc8dD
zB7DUCvxXmfn5BlQ53zJxc8/xOrNqpQjdx0ay3GAHmf9UGI6zJ+2PHgkRYAh
mHV3kl3iCU1zIu8qL4aCKPS+pBV6xpNDbH9/jqMvKJg9scZEDTV8O8DIS3oA
3VvMpYeFiVBApHR+Mt2UZZvsFyWDwIshnwIr4uz9wQJgEi4zPbAmjiDv63TL
4KLAWa3MopPKza/B212f7e5U+8KY+m+MPvakw1S3QfqoL7hJkbs1TfGIgAfX
q9LV6AgyJYSrpiG2hqwXradNaIpc3cByXBQK/71Jl9GyR6bHgwLcwJjxZcSY
qnmXxJiBu/LSzGLmOqAzsirIOzlK7Ux45OP4wZVxvRzuAX9NVYLsZ0snBIh5
RFPnF/4PQpE3DgoU4zrD33vQDD4KncClTV/7kxlgNBq3ToPz6xAr4+SrUwTG
bElDKAjZ2BvdAylqwmuz/XYKGIJ09l3AX8kSNiT1cBc3AsfxaarJrY2JqD8n
a9sDn9ZlFC5vgG51nVcp03MEcYaXA0zcH5O3vWNgCS2EzazYl9v2v4U9xG+2
PIzmIWuzYTztGErmJ4y9Qgq/iMl0AipPZ+Ax7ZtUESrRtAs1Tam47lMlKTXz
36Cs3Z4TMnulpN6jBJ7NdATEjRXC88J92JuB9nE4hxvm7CaEZ4tmersHye3s
uhB1DcxHYsRANTBM8JbW8/uZyoPpFnL6t7X3bfqM/KfZQJS1TRpTFAQnp7io
/gm1iHjdzlGzMQdoIc5cYfzcUPyTaj6xNlvySVEVNb7fRviSK6LWy7Zh1TfP
a2b3BIpN0eDuhm4w9baOqv2i6ZAgStSEdgxNI7iOn8I7RtNcBsxTBJSJgss6
/toKq4RpPYleYn+D8XMcGxm0YdZPJOqOLRMQIBaKU02bB7HoGSAx441Y7SaN
VhA12gjxIFR7pSgAoJICTbfdwa2b7IcddHx10Iu/MpQjs3dVSePBMlit6tSM
lqJ00kf/Ut381Tw1Iia2ALmakZKlU4AjtOUGJl+CKWCr8WLTNJucy91xKWN2
r0FCJ3SU1E3KxwROafSx+6ywUIJg7WrX5RuV89qkcmPPwJoaeM4UxsOenjO+
EwjhIjp7JwJ8jjIqn1FYFlKToyCUij0uo+bocEM7lJ28sq4j4p5OUQlQUCQT
+o2a3Xhod8lMSuNe+sFpfnvjmohzj8IJlA/ZG9LrUxy70FuhXnlCbcNeHU+T
UWOHT1yZkptZnG9SLf6/96gYoT5cnejk1SLtXwH/IB1OSYtqFooyfRjvRaQ1
+wqp7f9T/DKz3A71CQPEjKMrbawSXsvZARJ63USqBpBWosslz6HU9Ztc2aQv
3XTzy+VMy9O64B1KUAZc0UbgRxF8jlNb2nxNHJUlK7mHiXbll/EAj2EAbwlp
yafFquXpqKW9VQPmWI/EGkOyRJVImtDtovdLOgF05+ptLzZfrlNlk7imVKtR
v20jYb04IPhZTJvTomUsmfNcw8JBeKiazW5ZesDv6I9BONytXtnU9+l4DwCT
RtbGh+gMVtiGFOkDGJ149DkQ1zzRnnds9+Vyk5PE5wVDgM7mLUZhpIqfLqHS
6gGI8miLK2syVx8kMhmMPmfdmz/aS76CjWQdV4F0NOwfvBad+Z/2cabSMiYc
XqarMWCkrAAmeCb1RUnXtkj503/glsOWlQmtrN/S3YZ9lr5/LQn9fCHUQnTo
5XxU84umXal2PyiONXmBZTSMb9jxhjguKpzquB76iyAakoCweNsaRK0Zj17C
C9MaVYQ+5nCzQ5BrDUM7xoXmVPqLze4LJE8ClHxtU/jhm2Y45gP0Griik1ae
1JfhPlKWohoIlXAj+Gnvkpq4sFKLiFelOKE7VsUplIfuxkzFSnJul3pCAia1
3ACn1VY7rRUnR979+GwECVgrINsuBOwJq6t983Px7ddSAjZzIWQ82xEv8JXh
0j4pngWUYCqChwnmV5QQGTpkXzLJ34oFbiHK5dZkpYgA+qvSeSf/s2ws7WXI
wrxdAMrWD616IsxX1oYMCbNCUGkIwvrF1SoblbcjeExUlbuClfHYelzMIN2R
lBvSQOW7uSBByVBSzkpoYlM0faABR6vYnWOL2GFkbOAkEQz56nRSEKvVcCIe
I56IB1fgiYBeyeFZCu/7GJNkJ9epxY9XMZDmEtxisf0HrkQf7lJrrgdLb3gO
x496bd/mjfRh5ew5kHlnjJ1yokoxxmX0OG8Y0bjfBS6Mfz2WMII0AykvSUHe
pFwwWZpQMpsKxS0ro2AIsxgk/spPmOpEWQIbUQnt7gzoLmzeTF1mSqGfNaUz
x2smM/MFKnfq3py5fpan0iAy4UCapLy7tFyH4/PBX8to7g/dLVSc0M+28IQZ
HptuLR2t9AcXzP7luNWIW8M6kxlW+FaVO8cFshVHIuZuoVkOp7XRI5Vrsg5R
1iXyWuEF2RU0Joiz3fkfa1dBb1Uw6rHDi//+JNO3RrU/tJ6/DnKjaPLO6y9d
FqqRaYFsSdfD4tnePjwSM72JT2ZR7fJn8wVdJZmdE0usG+DZC5QP3dADOZpS
+sZ80gp2G1DReTcczfD+KLHwpE1r1C+RQ8qS/Dk253r3eVXjzC3wLL+cGHVr
aJXjiGzepVWqrWZO7vr9Hu3Jei/eT8oCALDYlzM3g+q6C8v/FnhvSrRBvwFo
WLomSQzG0DWunRR3Z0Fald1CkQqQpau1BW3UNnOJIq4zSU7KPFKbs9Z63s+S
PQHYYu7NNDmgrn0IiQFvJHp3Fnee8UqSWWBxEkqe1lJ7XUI+kQzs1IHW8B2E
ILg9nq17e1QMPI+17VtC5oquJDv7mxdDzMNeKCDeCb7CAb2bZfMVpwML8E6I
lvChI6gRNGB+5c7ry5PwqlQkaPhVjDKalMOuusHt/moLnvTsl6Zxza608rgI
OVOx4gmRaSuT7gwHPZArQhZNsebygFvBrtShdJoOoZqiIsrMS7RU2McPUSKq
eh7rMhhvwMi4o1Oa7TFyNDICf0IkPN4ICcly4qX4q48dDJXu3GA8H3TEpqb6
7tho43uX2oCft8/Vm0Dnq6mChngrAIcwviHg1PF6nQ7RnT0ZR5czwgfQwAQU
KmTMg2Hy65xSRR8lNfL3YmEdtVUS3WCbvfI43QkRbb2+h1i8SoETAlrIAvNk
z71zMDOgsr3d79nvwKKB9Pj3vAjz9Oye8e34WOoSdLT9S/VLh2Z8N8Zm4GLk
w4T2/Dp2N0LGI3LB+FsVYXwAqZDXTRh7iOgzbZJ79aBIq1tUlAottmxtCwgA
ivX60pPuoak6mzPoRbX3keMhQwUO6X5ByZD9qrAIZztc7IQyx5wcCLOD95YK
AQXvwxrATNOyclg0F8FjKUd9D7Cc4QA/DzG2zEp+YS6drND/fr9svJOLtmKo
Rx6/wjI8eQgd0v2zbidXJccAi/VWvXC6+pwmDlXjuowxvscqwI7ucSgquMqr
B/6AJJOl7FSjxrAK5l/CqNlE3neE7h1xfqcAxw9VZaXmPpJLExAxB+rHcCkD
iAhTyMasVpyeLvMrH9aNowRw0DB15+5wiDrQULm8+HxURGpiFNKvFC2B9Cih
Lmtm2U/9AHw4rG+zAwddVVCmBbUfZe3dB4OFQnodDsWWL4aV5cCTvsggKS2e
p9RikxqgWm4yeJbdmvco7xlhLRXS7fEx514Lq/rMAgFa55zhZO9nFCjZtYJE
sq/ZMICydAMLgzLi6HAVYlZsVSPUnCCyKTB5eNLBPbS9IgmnZ/Wuqd6ArI8M
x6V3NzQmjTl+t6XjUhktBvhEEW2uuCemf7ga3tbGrF0hFtlCK3ReQsPbDTqn
p5qvah62423wUH9tYA3M0LQWR43bGtETnQMRu70CXidj08Nc2uzf9GQvx5NA
XTbHOY1guCHD6sGqWUWHUICMjGKdt2eBovSo6i9GWyShNNwCE42+prmAEnMZ
OuTaOdTJuyCHVCdKb4IV7gIzDoiEx9547n6MJZ96C3Ocb+4ZSTIDx6ZNMjFv
Jsl4XyFG1d8ynQcmoKkCbDSUcjBE7jO5uEtg5uh1eO+sDCEhCvZ3zuOEqzD7
oBd+vnPDrfRgsLuLkIhG21LriBurESl7J3S5Vh7jw4SOPRiq+g29Vd43Gg/o
pXp+Yt9ZSUKQBPDwiZ9TtM+iVM2kIFWytUD0bG/TYm99D45+SUFWSXkTV6oQ
IELL20XmPMQxz+HOoFZ1GZIR6f61LTbACYXhmcfluoRrI6MpJcyuNxClkDJ5
lc6fugXIt6Av8Lr0AN8yGpLEY8ev7vMnmsiVZPN+VbhpnGRR1nqlvdTlouM7
T3k729vdET5Uv9XvZjS9rMsF1CxpMmzJrh5IvXFaIOr1BTPI7tKr6boWMzNm
wVxAgkxWYJQeqwgOH1tb9WtpwMGRtWtRcMA5SzT2ZCka5IrFIiQYFW2m8QOO
L4GDOT/FQ3m3HQcZHnxihTL5volD+n9YJ9EL1DcQKMjXHixuyM6DtH5kl+/E
i1ryXY6r8qysFmbV8i1qcP9YXAdeOhZoiB+497//VIA3DqfnEqC3gtsf/Mxf
4kmYMrU+iNE8Wx6IAKyzL0ouweAULRIhicLC3ovyHyphrfwAQq5KedkbP+mG
tdJ1Lgf5N/pY7M7jdyv6OA2eOvy9MbYM1hrFUV7HDWOUZjXWSEcLgLzsCCE9
YOZ4kVUnK9zvvMVB1cBg62hwrp3+/cNTyEtZHppDK8rUUyOyJsQbH30fvjLf
ux6UzwcJzGJn2GkvV0WkLbK51+mQ8kgb4U4aTJhM4iPAfE84VZhpzZPjdRxp
hBk2zYRP+IPPIfT2tda98SnczJZJCNFoXAv1ZU6y25fHkum6iUPvxdb78mZ1
peTxfH2nMfnMggx7ZLdeMuJEMSxJfnLxfp7g8v5X08M2M1rnIkpz50qIsmDN
ggHxjMjusNwTLqeeMAY+buesw2C3z8jF6dTWgtZZXakUjXVh0mElK5T8PrIz
ubrtQBnTkAqzng3uq6s1LqJJu96jdkXIr2WSFpOXUlklHksp0kKHqzDo5xUB
w634FM/aWmJFEhNGDBr1QaAo8lHkyVi2uvRCIUjootus733EJQ4pJkW72uxM
gFc9hJI9GIMXoAVICIW9Dg3B6cX+UkJ/OhdBCyMwYAdyo02Qr/MoD7XKGcwn
ALTB6Jufi9jGOLAnmTAVrt3Z7ohapVM8XezHs2hOtT3l1tAUavxxp0DszdPo
TPBdcj3K0eR9yCqB8gqdgKsRVZpGNTx7HlNs/WTm5V6shRoUJrYZVDSehVUR
MV6QvCBIruAmDHhPpGfanqNxw+lidy7mi+Z/z1NPv2h3F4+qy2CycJM/+mgi
uBsLE3g4386G/d7esQvxC3XS1/9jUemDpHvOr1T5u2bMuyI2/I0rNEmTkYel
s4pTTRA35dgvMvPtHc+Wm8gt1ANaLhiwmi6q0pH8VgTy9HqZgNrG4DPNMNok
nmBFhPgRE3cpTOJxtH94Sk/0qJZpugbNFM+/XnGK7rYWGmcoA3/REPwcjeuw
Ng7ksNyVbqoXnod2uO6UAhqUHEO0Nwh+seQWOzRwTDOv7+gstNGkzrmC3Ct0
8xJzQd060DZWqRu9f2diQCNF1LoktF7eOhBL0/1CQ3G0PfNUbWfUvk88+EVb
731ByhgmqHJBGjbtFncV7o2PtJvfGCQgcUVLISx25p4V4ShnLNSIlOlBeJ7k
8M/eIyVQma+B8cIXSqxiB5ZauxjHJzK4qxY7hFbmOR1B6w/C3zKELyEMS3FR
TNE8IsL2W3DnOWvUvbkKXbuVv9fp4Hfhvubhu3X6zIO5nvjPTjT7AGqnMmh3
XvoNlSTzaXDce1Dn6OikY4gbNWlQah/TeT3TY6faV15U2fD3+ex/LjkJwh7j
9cZ1wQLZBKb8YHMm3pr89oI3qBn4Z7GQznvLy9lCkiIUKaGC7O+A6+2vMIdr
Yf0otzkR60IsX33OWWRFSPDnVHAKeV/GLXBWLNB8Tfk85264yKgjdhPZWzL8
tNDoRWfieTXS8UBxKxdC4ePPky8MUydLX8Xt5DchamjhvgPSsLA9mGjEKZBt
AjQFjlI0WpCWCQO75qJxVx8uAc9Ajs+HYkdqy3C2DesdB11G0JfTlPj2jfVD
aLJ77Jd4SmaFBOR+XaVRy9urZovWKHXOyJ3gXx957/qH5zRNiXpOTcu3iTbf
edl4IVIFGpRv2e+ZAZIYGsP792QlTF2iMyKEVik7oZvysKay/VXQERTH61FX
7lKoVLXwKP1FJLM++aBCJdL5y7taB/mJvs1sNiAk4IJy5p71I5JKj8wRybv5
jSI3Pnn/c5jl9bKB3n1yjsSflwW4Dmzrmp+rV5P/opLZ8KC7N0laXINHiRTN
leKazKVEhFdyLIfI6cyYuAo3zPvrtE9wk+WmHuM8UNSQLp3aLIFewVBPjj9J
qu0mdbZvU+HXljQH1ROCtiF5oyRJtydVtYapnRppE5haZo4MucTSJ6grmqGl
FI1vkjTqh5v/mMCnHfP2FnzMLqyKVQ3hnoxk2Dce/Ozgy4o5WA7s17MAg/H9
NKW55VEVCFkQFGvfyOMZI++lgQzC+ijPBbcP6pI7eG/uAVvIGlU3gO8yBxY6
EbI3qRPfm4MuYjIfF9CnujSaq7EFpXaMrdvqjQDq+ZhefBDN6ySpR2gO5loG
4vR2x/pgyeZkLktnrbVz/Q2JG3g9ucapTTIme9APxva1VaLVUNuQbkW8MRLM
ipiEOGSFBr1vNRdXoSWABmMs4BqxmsU9WUaoukEVVkVLmNF/XV687G5qVyDN
176lFPHon8v1PBlvuRKLEogAbp+VBHy2ytSef//5Vo9eiLV11qaTbUsYB6aL
zn7tE48tLRk0agE+nwWjg+cIMJ5VHNCsLvk9lQ6gifXpnbpt+8+iPP49eU76
kBEihtf4x/hDa/m7sCayohxv9SOw43GnAkKCydkNvuWCcrIEnQRoHBhoKvFS
boJ3ApEMRf4iU7khsVU1Y+dFL2mafsjnhUCA8QuyEhHyUpXdhXIlfc4SjDdf
gPskcT3fKpGJERQw4QymcBRHRBUvR7FtXcFxl0Ms97AQZZ9yStkkr/PbGJuc
99nn8PAE1EGM5wRXJ7ZIj/qv95Mc3KvfAAkmgdDBmgPB+jjqUnbQjTZk/Wx9
o9XHnibja+No00thTVvH2yTBc+ragtNYljaQByiZwXo0KDvA95kna2RMJLaj
219Oel6vJKJyLt7D7C3Q9Q721svl7PtphiNwCghYW2ua65fSBPlyqTKw3Aec
/VpTO/GhUrrjpEBebtpkAtCEyJNJ+vcNbJYicwXMLQ2l8q74ZEI3Krn96xWZ
D1r3FLmyApZkopUBLUnXAM4zp3EFcDePpg5K2HkO1whffL99JfGYLIsrRqUl
VOLHr+rV+QcQCbPVu4Lz2jjLDhI89MJF8CwYM74ZjMeSHFiQYVyKLzTS4WqL
IgwVH1+MZwn16i288riUse64h4Witw4YE2sjDKUSS1T4pzP7AWkm4cToJ8x0
IneIcilm3NYXicXsz051LCChi12CXLaD5f9AaZnewH0IZOyhLAFIQg4UjbC0
AzhY9CwTOZbwtJmsPhaztfiJtIsX1Fo7wV4ogVfz3h69Wsx4t0eeX48T7JFX
+DtJspUGvP1ETLkvYfkTI3vQEguGo25wuJB8deYOCKurD+hEUYVtPXpMOGbv
54rOU2Dc55FCrIGaAD3TnFLdEzIp81iC2dxKp0kZLqHQK3R12PGYcXlA8EAK
RP6B43ydUff0107wqF6WBmkq82Bc/32xn++SRaL/6biXqny/b4YEy5b96VQv
j4MTpIpudfD0SqgqqnYWl8OIVdNk3f7HKcvPPgJm4EVlp1YqZCkUWAXLsnc7
ZvRVSXufRB1d2S6Oa2QXeuIs1v7X0gYXNdbn1YWbCAYKhqKtxHdqL4PZSCqq
WIX/G7dkLm7LtW84HNBJAYvcY+ZP2595eRmfJ2YtZbWQx3Q7H92yP77spxA5
11AN3LDZsU/m5Kmhe2WkgJuDfYvglLTZTIySr4fJ9fndLhI0mHKio5JOLAAK
NPNdojPl528+SzSxOVZtfHiw4Zmr+XGhTKEQBaNQsgmFE8gUuBF+d+IaezN/
GkE6bKLWkiUJ3hhzC+5SKGiC3glNIMVVYR3Gy5+FRXKYLeooh6/5h8fX8X24
KMAPIQnd8dfB+TG0+udNwi9YaOTp/dWHQx4Y6REWTu/2R3ozO+shbyugAzLM
6CrbXTES4B/sjTGS4FC3VMgs7eDaJW+Eg/E2F/VeKKRbG5gzKfeBw/HVgCeo
qQQorO5X0OlQarm07hpVxBvWU+k/tMm7HOZ/IMX45c7XfHIgno7g7luzXp2t
fo5hAu57UXdl5C9qaxIpNGjR0ge9dU4AyFqUX1rT+iFjuLnVr50aCRHGVL9u
gUR7aK2NDMd2Du95iW/W9klndqeGoTP3R/LmQQ10QMArM/4VUygJJ+WBvF27
sMdcq7inM0H/XVCKWqKWqvW4FERBTESvSvulwsjfUKms5wyL0Jt69PqdTZQh
0obma0ZmEGqM1hNAcfI3S8f5O8YuVn4boRI9Wx9ihBR2u68sDo+ysbJHX+vs
GOgjKHPeNUYbmnRF4EHePt2EP54Qk6ZpOazgnGzPHlZWux6cnzvo6H6dTVE6
pL1DPIIrSP0UbVrlwlE7ihHQhJRpi0T1N5iYpX+A2IBYgygLObWZjxK+WcGR
pa0bvpLszzey4tKWg8Z5mWjI9yAqzSZp+v/mhI6pxA7x53WhINHWtyHdfb5Q
rlIAd4CJK4+1KDz4nT0kpw5iOmm42NXeg233bXqa0zwCCBo3fNtnrOX878ct
y8ACcyShj5GMexyywN41VbdcRx/uCgin/kV8M7RpHhVGpE6KK5vwveojjcEX
AYv8P4gUDoGj8EaH/EBb7HEvaNQyOXl8ZehoV2as/JHp6mspUMPGqYB2dmyT
tkcMHh4zOEEAhviyLjPm8gK8a+u85DIAjnuvXgk4mFQKGQK0528k1txrY6Pg
6aWI+fG6ahTXqFl0PYcFBhyI3l7JT7WOi9LcrP4De45DjNz7mzPRUvBVZevZ
Bk3/cQWKDMLXKEFkJSYOmZTkU4Ww17m+5bnLYfjISQ/iuWQn2kxRZCfoXqKF
x1bSKpq3kGedCu1X3aMbobCtOi0kG/U7NiVPI+5E557dPXuTCJCEw91u7W40
XlmxBkhHOMhKeBEXTki88S1zoKdl9Dm+2xTaytGyx62H0HhjGb1MBm0U3dxZ
qT0MPRvKETtAtnAn8R8GkhNsWBsL7Mbi3es3DPjjjUxlsOfS43mz+RjhCLrX
tVD7qzstMgNvdQLfp5Q6yoM8HB/H7BEKLp3KcUhzzjBdY9aPDY3OlHYofiWw
Nu9dKZC3zNgyCNODiWU55ATFvyoLOQomzj6Ff+q0/1hdzOn9/jmePobR/xNX
zcKgiE4xCxHpLBbHc58aH9P82TiP7ePGpXjLjhu+E/YEUNTLE86oCBMrAvdd
AsgSihHjPR4IIvr/KfkPxfFL4Oc54pVC4EE+pJVu+tfVdfR4g0lobiMJvXx3
Yko+MQ8Vwq0UNYflu/BJavgv8NEy5UiMEQGoGSkPmI/9RkUGvFkc7lbnCvw/
IS1wUyn5xWwU6xE6iCOOJtbLVLdkkf6EDXpEzIlXoFA/I4f2YFtL4CqCQjKi
yQPWo2P46j3HpejZXZB5CZi2jDE1VS1QLjvCXLsXl5bZ4Jxpj5ikPeQUyWvV
uSBM3K5TTwVf7dw2UOcERPNT8TqhLJbYeEfGxNlonBhYxFSUP+aYmiK/1mNY
hauqbPOTpAYl/gAW82FJ3IJ2l03qV66IGP1cS50m3ieIMCdRWl0hwZo5GEgZ
ttt1e1KG6CY8aPdBE4lXE1edoU64qfb4lUh54bGvYYZSraM4G5NoWilB7lLr
LFzTKgRkFap4ZJ7HUaWhST4oEXpYjnn2TdvcbeEiXmMpRCgvryi/7ValbgJc
Abj25WSn2klHcjm7r0t1kK1AfPuBN/8+8XRUBwPOQqUkqHrKtV07f77mv1Ld
J0zhYeD8kVeHyvEafUj21u3nn0Y1c3flRNr0wZzF+MuOR5QTF5Bay7i3ecyp
FakLe6fqVfeMgxNCbMhmMuwNqWKO9W37alifjZeo0wnr3mu2qUa9L/zvi3X+
5iTNmwv7DA5QqoElURsjS/nK05BU+yfmOp1PcniAwzQh7S4nVdZ9gAUv6yp+
0ZrFrOAoh/2P4f4XuwY/9kL9HMUfIE4Du306PrFNn0+B7BXCGO3eRLApzKik
mY7m5c+RtaZ44P0lkUG2zDWK1qtLBL8ZTRFceXB8/sBK8iSJuqtY89hQtGw0
G9Lenkf0bMrKcFxY6JW24m0Zl0MgejtZ4pBZRaYZGhS4kbOEQIZKbnh2C/5M
C6FhcqAuzjuyhM2vzzIoNl08MKVjEWNzqq2JSYMSrZwCZAyyEMeVV05Bp+NC
kZ+RXU03bZb+NBkl5l0sLj4WAO94JyNQfS18ZBw0bhPoAesbE0/Bbah1fjyY
zrHVEIDQfL2ZaLxMRW0E6TRkH+bEcHD+TY+YBbk9APrkrcN0m6fqBZAaze3D
Q1A/TA/3Zz9CyxVeACcDOe6c1WMOeMLRCf93d0PE/xbieXPI3eRSI+P4UAnw
t2CZT/NJ9DdT8NC9GJCSwXy3Lcal23wkhMKQsJwL2KIIGUAuqVO7c4+RzNYQ
30XZGpmDicPNQRAj3hVkBfIu22BIChY+qV6YA0ZbMCybywH70qqi8Whfdbmh
iGUht477sJmwh0hxgsMTF48X1nnRDKvlhLY3/uMLfndtcjVbW44hG79KEyV3
29h0xgWYZqlyofgpaxWbEFbDY2OEcP+jsF2ajc+zXhJp3Gqsrer2Pc02DQaO
FFTpEVObGXyuC9hEr2hguS5aK7qwknA+peMKEbGnj+47mSbv8d4nH+SvpRKL
eGOq7NygDbc8BFfcNeRQ17eufWRWBJz2ObW6J5iHOelHVZktUDodc73jPR2C
jI0H//TNbogXMlrFeAyb9aPC74IymdA7FosX2j6JrsRadlxBihHhxJUeq7d9
3buG+yxne4bbVKSvZgexxOc4O+YHtEpphoO2m5jdWz3RFsdWPtfbFdBzD/lY
uiyloFkfs8bYhBzDswDfLHP36ZP7MnI1IUvbMdlL3QIBTGvoZDf9/qnu8oLN
B3YmVpkmdvie5ny2AfW8hX2/OUL+C2q1blpFltLOphLJK8HMhSUG5vM01/5H
4tK8MtEdYkSUEBUMwH4HeU9S/+Xd8VMJ4wn1u34OcGfYbLiYawRPFaJx7PtI
3zvzueWYpvCxInBa66OsUAshgcyINTDKelejO1cnqmIuV7amxtZEvKciXs0D
KnnpmJbIdpTkZKDGNnbbEH0p4PDmv3q/5CU5v6oTyVMZAKNyK454aKaGoSEF
U0Psine4AK7n/oIqYb1ky1qf/iMBksIgPNkXv22NpMlCybaXmJd5+lyaEbeM
OID58Zs82kPplBV8b322aLz/ZlBXpyPUsqtaa8CACCL9etYLC4D3RELFBIGp
tStUvQF0LyECcU6JHgVdwNVIm0MjwsIFCObQi6KrXzI0Izph2SLlPpO+8DB5
KHv1Poh1hT4scNmIApyeH6lUHMZOs7DoSpQxWVVxmD15rYg6696JtpH3CF+e
AXgslCXkoMPLc4JveGZL9fIR1Gmhw4HGvXGEP+GzogcxDum1E39gQY1+STOR
/Wm4kTckP39QGPbzSozh1sFJ893REaQZRiqrLyynx969qPoIXR37gkRrKA8A
QOSgwisodQwQ8nXtzOyD4DG/j20g1gArZpoA1NAREn7e/1f625afuBX4LBjc
29irN9d+qnvrEnDKlOUy4PQolpY5etzRtTdYtAIMwR+ZdQzlRpV1w+9JO6cZ
QdXy2KbZEU/lCEr9DbNJJ08ktbJtH+gl48EpwJY/mNh62ygMmhLVYklP6sUb
pPloZPRiQcUDAe4FbRtHkhYx++HpGoQE9Os2rQrHrCwwHXEryirBKxkIBWJx
Jwda45/wqAub8/VYxSHDJcyyKb4tYPAZnmQX8xV58bMsArbyiiltA5OqDzpA
3noi2jzOu1i9LOeS7Vm2bDkKgRl4alzMw1KolYcAz1ctJMFcb6f2T9gwaoRJ
DNZaObk6hXiXyMU/K7jIzUUAc6neRQPqBdHEWPV2GdZ4h7emEIdsS5+yGwrv
RZh1BLs1GkSmy99drehdAttPEcGYRYdBOj1+Kl70QB58TNI+brlpfD1dHOYc
BW29pyftgjYw0Y6cHFJjntfoA5Cjr0661h4WPBPithFZOBtqHttL4ih8YLE9
fBNsmV2lJ58MDyKVaW/PKE7+qCDCdcLlenSdN791/z138vm+i4V06FPPF8Z8
HdyxayCwbksikR0yqjdk/X4MH2WE1pGarOe0McIFgJMcghcaMmjjv/a8NukR
hviKX6dlrrIas2sLS7UCpT5S7QASzY1A6aLgFR+YEMUhTbUZcFHUKBgY9uWD
S5CzNc40XPlAHO19SAuK7OS194T3PlawvGL3r/xEm2neSafOrExBVSdM2dvt
6v1VJ1jKg+2qQ58kHdYmq6wZV2mIdO9DcZcC2/adXwdjC28nGAp9fqFtAo/j
e5ClXh1G8+yFvDbI4pbvBKIbKh0HUIM9VJnNYPeCYNBMiQhI4MiB9+9dsGpI
zPtZfocFngWuHt0fX/vFxiTU7WREmP02CyCSfn6cm32Nfm1odltUTu6K48zy
ppFx2SsIZ42qwx+H0peNg43nEBr5ANskEVk9nqoe4qoXWYG0zIhWORyWbfUK
0ksk4c9InHoDWBXMIbwKfOBSdk+NOXX4b13pPnagryrO7uGoYpxP4tfnMGcA
FXqErKFUpQaFjyffHuJnMcktL2zBp2VnKlTvgai9f2wlaxOXkW/BN9NUI05n
cEbgW+5mUjbIqw4IkYUst/OTfESru5ioA8RtpEwp2JwGn8/CrVkIzGEgnb4D
aEnx3ulk1MyFWd+FeaxDAfIm0Vyqajwf5D/TVRvriV587f8Uzhkf74uCR2qL
sUbur6TIIwzwZQqNhE0QGaifoBb4DqJ2nG70E3gQ+cRsVyf7lbmRGbJwSU4Z
hBmqHGEbTUDxUrGUon8+ElzjXCPj9l3fsjwd2bpERF8mq85MVBII1RXaIv36
9LvZrh0zhdIYyIpGebDT3AbU4O3MIxWcR2VOuZSt47gIgpBCS6GceBjLbHra
VZ0rruJvwpN0DxO+eCUpw9v4PJKZItgaL6a+CWaEBIpBSL+LUCyArecEaAHz
ZY9gdfvjVrzJaSD76sGtstuRAX294CMuk6DPiL6PCmm2XTTDY9zoYmXTYYgU
l2civOcRgmKhU6bx9rfyq+i7EC77s2MIDw/C/Jq6lLr1p46qNAZaRjlY0X64
ZDbF5uEU5EBjxScaWcgb0BmdB2lsVlWlM0v9vUYLwLj15vEy5usBC+MFwgU+
CHNFJDYx1Lf4DSStob0VGfEBKvUyKDBdoCQF7fA7ZtPBjFI0TXjhFuVQyOeF
TkWpEB8sCJNqpECB4jliCop2/Ml4wWUEuUqKK64pgHzxi18Ga/74yn1Kkaey
37gyD0XBuCwPNotNLxwrEPP1BKzVrJ5Y3JCaG5qAM/icFWh61FUVoCqlw2BS
AdW6S2S4k+wGuxfwGNgH+KA21xqYNYejkzJ8XhOxtFmBOpehFMZgQ9GX2HUy
nG0t06fQGdFRSiot+HFaxA5o+UZYF2iIf/YhHO1sf/zMe3+jS4OdU3ioOtcX
JP5vdxW+Tah3vaN47Q/BNwIVtyxncVNhJksmshQTDll9iPTv0pinqLuYjLny
Pv7PQq22712+IuiWxHWe93rZSQ3esr7+uVY+pXyNR4XHpyY9r4Md6Cwa/rRt
QxcjyLk3j9qEzCLRBQElSUctayXZ5FTLfBOnL8gKST9WZet4ynmX0cOkPKRq
xn9/no6tjpCl8Xwz2gylWQy1ckZUg47Vuv4B+ZmHoPoxgsyRne595t1irRa7
XjJzDv+fqL7oatUXPb/hyY7+ib+T+JWXWC3+8LwDAC2xSlbd5Ap59whO5fv8
5IeS1uOCd3c2nadqY5QXdtHCXY+7ONehd7JEjpF1IM954MBpH0jQy/CZplXl
IYPq9kmeEcYKHaDUOYzbQy4OXv078WqDr/VxbVT2J7BWo2MEghrDCA1Hp964
9H6y9HBX0HPU4JIVVL2/ue+CmgySA/HWqs2AlGsK4uctVouwdM7YGBPsaxQ8
7UZrVTeWx5eBMyuOWWLgCqqbQCe6aZelznNq//CuEqgK9RT8g7B0tTnk1Klo
1SSFvJokeoXZ18dbbkZfU2WRdgofl4s0XJG0q8iINE6UZ+N5Wk56mD/gvN9Q
QDOMYx6jaiRjUcT9ROpNdSGh+6Y/f2e+vK5bkx2IT3U6sAx7ZAaTvHeQ1avO
ld2ggNZcRpAsovnbviY1NnxpBhiK/99xzu2aMRqvXbtV0ZwewTxoaFJfkiFo
couyZHaopI6qjb1TuI1l1RgP6T/55zsjzjKDCRc0M2Ag9Z0bWTjM7uyPMcax
LsfXGMZQYeTEFFqQgHQkqN1aZWMZgfO3bPyjQJCt+/ynPGjrZZzAsJ+F8bvo
qbZR3hqdWqbsmDYXtjRLNSMdV5ASGx7ggXKDU+cKs/6YbbYLw/xeZlLnbz+c
ZPjTZBXOCykLs9tSZLwvF8duCifnhgNz3q4tFsYtdWrUCwmwwq+IRL3Susji
xWsE79H0o+bvhHC/xtzsKTi+Gt8wGViyHPqngqewYddd30maOXQ4sfwEFunC
b2XyYkzPAH5F1NDUqMsuGoZj2tEmDCspYnHvD408CQf2xV3GKvyDcukdfSeP
AlTgnqTwzGotIPVid4dN2+BnFZ/yeV4+WmsbkMOp8TvUzh/qFiE5PVXHqPkB
XEeJLJ8Aes6D7GuKyolArQnn8beQ0xemoxsigYzl195rtYEvpHf24iSZC+GM
tcubs2BA+2qq/cDwuG/qNmR8Paq/NnLVpZ977QfCWYOthoggPIc+z5PLqaoH
KAK0HHkdomHF23o205pqeFf6HpzdbR9cQDWToDB4nHpebHrtoNeTCAkBFZAY
YtH4Mtgnm2LHSNMr0kCepcxEFkxsNuo6TUBc4F/6olkC8MU3TVD3ZAjGFGSw
eXbSiOmMfpDok+N5xWeNh1q+Mzzpcql/Eb/aWQEAa4VrRAhRpdlx+66wqzwO
kPIhm7ZdUV7esogs5yAWnBizxAAdZWoK6gKkHlmd0Phk6qs7wxAXVasOX+Md
i1dv0oToMLUvCsOYKVhVekSfkv8uT7BYJK3GBMkA3voEFhOXRjsCxeGSM1/Z
BUvoo2ojCJISu1EBX+U810KmdMAR0/ovaPYGkw+/0qooTajChgr3xOhPaggo
T1e0RUQAuehyRJYuKZR3C6Ritn7E2AGST7mGeTIQo7Hfg2Gqhvdst8tFG3Wi
N/5lSLHXjdqhbzjpngtUSK4sC+47mx6j/Yidt1dwBPCJI9bDhUF4b8ohd4uh
CDd84uzOyDdGkOTLejkQ/tbWfQahda/M4LaHrtueJCsflT19KV7fVTLr3B8e
s3Qhij2W49lta5x6tnZUnfJno2/IJXHydD/ZTwBu0ZcZ395h77VgYOxC1RBq
nA8hADgjgZjB+qnkXpQEKTACd+LcK3TdVUOrq4UGoNyE1uj9WOKw1bO35qSy
nQLUjpBB83SQZCHvAD2Xw+Xp7r/lrasagB4muKr6pNbOLT1HGvxFnqMfTeGU
V8ztbMrnAyUlY3gQMNXF4Y4M4nD2zpNPkkcHDKtzeHYdqfp7tVyag7eoGqGM
X22wQZrgCeqRMtflFxKzMBKKadJkeqdsPkK+rkM3/O7GVVMA1W+U3gPYlUFE
LW7MDvho+C5rdJV0aCx429YhA3WEV2fDDD7LHQR/goo2k8hy0pAlDpb6Gkjv
dHjZ8avdlWWbF13e+PPL3Lff6UbWteb00LR0PpdMI0+Li9/qHJvngDbQiLqp
WlGQqK5pe/qkL6BQVFsPKzoJm8clFUTZMBn9y6mZGH3lvfbDlNatGgyJiBjd
Jiwq/lLKp7bQQmsUU5xopNd+K880/vvC7AodlBL1X1i4j68Tt/hGamw7pZ0D
fXzxLUYxzWHVakzHzuQf19eAoLWmNL2cV2XuXCfje0Mg0tz0dZGl8oCRAidz
2k9x+Kh0eT5TOpyTnIyOdsfqJbtyobhhvCEn+YPal2SfGmHh583qFxIRB8vM
0T6xz2PFcr3WGCvQjGZqXdN9tACd/gnZmt4mKCRqtcRWuz1GvSt8dvRe0xOL
AQQ/g+KmqZWN6CbCPcojntZbkMkSxfvRuFmLfKIumMaJXL7zIjPK02rDf3n2
d35U+mUJbB60Q21+ESD0H2cGAAjMvZOPZ/j0/p5OfVKWIQEQJQ4nvH3EtZkf
iDpaId1ZhpVKl2Og5lYZ87zHRZy4aCy/51MBroBHMde6qz40SQYfXxi8r31M
xTdHDUKJZU9sDnQrjZgeztJGL5l5C1iG+go6HKbisoOy+++aiGDJWFMYZdQg
73TjlzjJ5UqlboVctDIdVPvitYaLiK7SuXIMb3/I4NTWE2gQvy74QS9gsRm9
y8n+MQGZPGbzSkPqVzJggHXDaMO3pnEyfWvX24yGYjXWALU4Ouwll8nmUj/R
uBTjbFZXlM1eajd3mo7jfIx6/uFIf4dEOHVBeOqMCpILUQR+6NMGAV5rdT2c
NWlBC7dc9Vt9ZxD5TaS2M+LGOQk+s6xkyKL15k/BUJhMZmsrjtOpigTe2dxI
ARGjG+wtJzh+Xac5dHsukaLt+njoVOWLqf/5fBVz/lJmJFv7Y+v9pZYKIrGH
JLBX8mhXxnnsg8WHMP1Msa8p8bzWr2d8R+yZ6svHbhZW6IBhEPbnn0I6XiXk
R4i75AGAFfdB3lfKVmW2b8PPQcHjLu3ZbyhJ3WXHVTc0+faaCdfoW4+uOGK4
3rwYTRXgCzpR0tINbllDrZZhCjR2iycSQddeEKdPBAhv9c+y3ISSExqw1/ov
rzOZCFxZ0za9JK1Ur2ivQTXCqK/iRBqjrHyi1lsNtqWNDDea6R5Qto5448oE
bOFJ1Ed9dehoeH7GOg+Xuy5Y5Jt8N5BU/6/Kihc8dCuYUtfC1KhbORMb91uy
HmmIyLSL4GDPJZkh1KUZ7xTSmMpX3gNGninm/tmS+WY6aT02VkQDJJi2CPQs
YMd/nAPe8RAzMEtYB89aS/qWPP3/+yBQ3eOBTvDGe4207+7P40CHuPE7t/4e
c3I5RtGQ4F6YDRDibfFahuy4e+4LhqQPwxdXpayg5wNWAwpsb1zktf7w+xx7
Jvkt+KIhYZTZTg5lLumjJLjX+ks2B4cbvFr1Xv+9n/ruIrkJ9lRdQNocQUnc
ZV9+Yp5UH41gzC28FEfEiwKu+kWKxQ2q2RxnvCB+S95CKTVcfBevCRtgIXU3
miz2O6sddri5y6+2sllq1bsRfAqogCXBvC3oSN6K/oZlJ57Z3Hzv/Ia+m8hC
ctasMIoReuwjzeTy727kzlzA0BPZTmD5j4Bkg6JgfeWgGUyDiTVZHOmpw2jN
mYgGsmUnC5AT2jmEnirvRSdoSrxGLWFxs0iZ+n4a2FyFLVqxXwpOeb0VdMr6
urQC+y9Cn+Bdv4xk5M3cJDuEBvSbZtKu9F+ni5ewDfhhObx4E1+7QApCjq4M
X/6nY0IMt35y5burpCgDCUFg2pDRaggL0OcRRDZUer2GImoRk8JB9OmK68ZU
N3YPrhBfaMHl2hE5AYZyZOPUOesS+VYt3kiq45dvoFhVKC9Ufsf01oM3/pwi
px7dmKouKS8JpD2RBMuZJhmYDIZokBeQ7t3gwaDms7VgelQkN9BWSghi5LrS
9XJs4iX6r7y09HS28GzVfxi8JjAt95LiYR5hdyu4ZN8yi2XJF7bQZlMcfsEu
SZ2FYZB40eKgIvRZoPq0+ui+9JtAdJcLnjj1PG7wlloj6C0pMsjEiV1T3GiG
X9DJI6b+fIen/jRSY2QJHz2fRocJ0i9G+TFJSdLzrUupQrMUM80xLE4JCk5i
Jxgdlo1vWhOR9R0R7WupEJNzU0TVp2/qjsKNl42QyARGkvRjw5oRkpQQTlrg
1ALdZDP3OY6lpJUzS6hmjDWXLKhUy0hMlpxqztAwvhThuBYn7xnxoiVmiRnb
fFErFtjzDr32BG9uYRAloqxPnRlygOzPIS+Wpz8ekFpLieseTDyyJKc/7ayR
MSyel/pVeDIJLdd/cEmfph0RdZkFplFw8GzqOcCzSgpYxxVQSEaTSBnM/USQ
RnKGeST9X0Np1dsmD4KpMeDB9HLcXKLqp+odqhE6XubXbESqX8imqZyW4nJ1
82RemiP7+ZQI2zrhjgEV1dYVfByNytSvnoaoxqcmEa98LxRLxxdFFklNUGzl
W/yaaPw7JDDfvZUgGHg0OWETfJIOVb5i2GxDRgcAXIeNYgABBW/7T6aAtKCS
KmVCKL4+mUZE01THDuH77QQvdBvx5jDEUVoBOfl9niaVpAW4C/BS4i982VbI
f3QMF4H2PL/8ouuPy1pHra19MYIQpxauJb348x8xNJoDR3w+3g53aB0K810O
Ua8YIgzKEtfSlT6Wka7SV7t7PnhC6stl94T9WdxaKYuMsx92J+SKVEhF6xpX
4eObX+ZvOHzlYZJ+g1n17b9qe49+vwz3jpiVnO1+IwfaKvfe6SVGESKeAxQD
PAsUI+Hcg0URoq3OOKMNRkpgc+gPD3Cj/SwmwDqUkan+CaCQOsRYHiGwfCpu
YvSCC6udD9uuko2AWaiXewgFjrG5ptUVaHvlqOjyQi/NAbLgAUt3fPkS+E6g
JxEIUPSZsinMSnVJwrjZn05ljxl7+CrOQBNvIoLo8ZP1WmCwLeO/qJ6CCRqz
V0FjXdvF3hNpz28s2T/kriBpq9JgV2zAqCN9/F/t4eH3YtzVla0PrnXkS0FI
OSPqVT1yrnFo8dUun6v8EBxkj11M4wJAEsg2q6DJNMuSQI3MUu0TleLBDrOK
RbGrfwGZWW9ZOmbDNjSa2n8Pz8MlVyl6gl2HO5Wdu96OnrkuasB9WnpAMoZ9
3uVHLRIVEtXgAX+MbkPc22ArQQF02HD6Nl7qmCW7dHRoRss2Uyt4Y9vjqzOz
WD0w3gtqHpqjQA+qRmbU1RYNOyk/hu8fXC8HVjNKdW0VazlzEBu0mXVx5MnT
uZsOSnCMqYKGW4GcQpGxNdt8jntP4iHmtmgM+LxF7oMoFoDJq/9Q4q6LqUzB
bOXVoMS6V0Syiw07aewdqDhuFi5OmboxIW8gsXEBK37h9ug/XVWULTsuny4y
pWbbGX/4I9Ua/PyMCoLTbk5RbLM2iiJDYUDr7Cw0tRPeu8DmhP2HhfR7fDPQ
xfY/iv8zcNHl6GeKCRXkpjz8rNJ3sNZhwfW0pfKP74AtxZdTo/zIs7NunB6L
REDs//hTpD4TUhdSvblfkyNp2JZETrwrPHnyYd+jWlzLZIZyiTpCiZ0zUIQ2
OT/BBoiifckIp3uHZd7B9UP4OthYVRkcYa0dGHtvnIBzGk74YpBce7jVzCyb
K9rykDSV/IhlmHIdBO62HcKLwN8l2TDiRLxJSuHQscseg8DMjQUIgKftmQt3
+1tTpnLGvVyEbJwOIwxt2uJSaWRTmWnXoWI608bcLPq70lmN05sfjlFIwbdA
dnSKwoX8NeYXxhI5ON1RmAd3+Pw7Zb252klVHK2hiOFnVBE1xkaaZQAxQuUJ
VJI7fS2leFGRpJR33edbLI6PzapEUtVBqeygTqhnDj7qr/JKmQIQ2Divc9HX
6BqzMxbL5mmFeHjaeW0qguk7kZbw+cMik2DC7JWZ5W0YRzbwXUe2QV33l6cO
4FckO2/q+P9u2qjSbVKahflODDGz17JGqiTX2iwdTV3Nc5f0VKlfDK82ufUC
BNFX4SQZJkxn+EvMvzXSCDK7duS18PXDCS54IAHHFEpUkg61thTNKNxzbmDG
uxlQsXDGHeLLHAnj0x7eauAmfNPQaRlbFn1QlcX9PtUoq/FR3/P6AotthbBx
IxWrBBvZu1uh1ehu8s5rgPsF+YaW2OmsDvaJT7uJuK+MW5YXJKJUNtNWb/xK
WRztNpOaZw8zUyan1N4wF71q4Pke0LBxnMmGvm8tuP4ziTLWi4tLtsfky8u9
ViGKO629gUpxUBavQ/X9wK6oL/pZVUROevTOkTCtGwlnOfK6CJKn0TnPFzof
L+bEq0aU76immXfZA0ZwiypOBSy/ek8tU72xaS3JgkHibvmDb9qXdpbb76zd
XrFU4v5lwCW4Bff7OCL/M+C7zZCfQBP23qntTDLAXbO7oxfVNp1Nsw5Klnl4
8ALdHVm+IfP+dKCn2KDYzDKw4iwcjEKPQYGKs6e7SJ5KC2c9HTqTmVZE53YZ
8Lhp6dHcBZnROJ9LemqVj3o8jNwSRgCV+E9a853C8czXWTZ5w500xp7Ql3UB
D+cho/IrvpM3f21dGBUYjqintnZ3+QiNLuoPfVWwvBikWg2xkZdBzrQFtd3a
HHxT38tlS5SAaYPVTByf6Y7aux22om2ZKdHk/g1W/Q8dzUlu528gcedNxcQy
TRl4to4bglhw5F7OBvN4lPlwfw1iJNYuNIJ3WJr2rEsCAyOiMy4JpikxTGC5
8ui2q0P0SHYupDwymaAUkQcQ4rxDIhLchjOnyc3suPZkhmmpclntu7H3e/54
P/RCfbwrzzF/sYILTibS2/7zy93sA3jaeQK/VRb86pHghg8XcYo4svAQFILX
gHuGAECnLkeHSvFOxQEmIkB34aXMuiJIfpsfvt9FbNBsQTGnnZ3ezYs0VgQT
8bJPtUggHQZfToifxpmrcI37ozmndek8h2y4Adx2ANTQr679+YbPDXlD4zwz
I5/MIpCUbt700tWtVCsPua3G7cfhD/czTEZM7OwcP/I/feSMt1V/rqx7S2Jx
F5hf0g0XH52Q9iMxnlqANAFikOdsgutsWyVa4IIphaH/enSCmkKWs7RUzaF1
83QkteCert+6y8InAsi15rk6SSJdDd/HXpwbpESuXWSKMdg2yEU5pRNyBzw/
X0h9RdYBHlU8h4W1ooJ10SPE71RZlJc8fMxBUCaMaokt7JAJadJ50KFWmzz9
rdFPeYSL4etpNGtK9V6RfkTR1Jh9YkKR/YqnSdEcUumBsee1PIUcNZoQ5GfP
qX2OF8GNl+2yyOgTcD3q4h7Id65GQWI0M958gpwNhXvdN4P/FXr7LALxKVIU
nlerPuazmQtZvcUxcBGsaJVrgev8VAgwGUARS0Ydy5s4BzqxrqCNsgSk+699
ZZV/P0b5X4cTrDF/f1KLvZM1MlNqd73fq+0os+Iid4mGI0ZLH/DY4P/Hr7df
VyeDIvGqpD27XA+3elKZtZUR5dKioLfxDyMx//FX+huT+ZmUKhqcF0UOPVMz
c96QeNOVXPW0+SnjwMP4SrYSoKnI5fqost/UcVGpO9JwgQw8FL4TY4QYYefY
VxeYL0l3NlVY1TX3jXSwY20BPflkRiw97FnDFFGIIy/fxMu+vmMzjGDjvmNw
pAjEFHM3o2Q+DOJtmp2ZKzIAvEX9Lu1s4EQyFSFWpXeHF6nmQjQ9QAi0/MZW
JPe7FQUW7jnVAbOictOPvJ4ED+l60q/04CwOQDdS7K+YZ43YbwMY5mdsWKI/
2a0Tg2yPeUOHn9gd4Dtki1Q1PN4fGa289mFlswJWBiF/4cPF7oHaONgksWdg
hkNMJzQNclkacqtsYuJUNt+hPJg5MiMOFBRE52d70HW24ja+6H+O+ezRuQ2U
GxZU8EQop//9YCt+XJsOP+2B9KevNkjHeyPbnFWrVYCvFp3X+bc57+f+mpaG
STVGMUVpaX+9/tqi46baknthAhuddhSV2sxmGv3wJeJtqkQ7vJ8Kwxn9paCl
x/7NZi+e6RrkTzwTu1/yfHEz/7ZFvQR6TKeh9s8jXClusH/wZC5DFSkGq9Ok
cHv7yAosldViVU3PqbYh31vYS5yHOe3lw2d/buDTKzfJ2lpk6MNzRJhPlRfk
EiNxf5EpSVJBhog/DjoWTYx7G0ggzMrbZaol73UtrWoJ8guTLwdCPdTYZqvL
bh4TU0n48Paa+akEG4UgE7At3uaI6QkA4bIj5kRgnEoIJEHhK0HTjv0kpBlN
LFCdVbtQvsZYArTFLJqoWcCylZzYqeWWoatzI4jfeWsVoavy+kfSVNc4dEIA
m7lE9To2aplkIKGy3Dk3KGry6r9kLj1MF9mcWcKXzLvGLUOG6zoyaJX2yhvb
I8Ny7CNgomHAdjpnWYe/SGvxtyF+HMwfEPyPDutDLW6f8bG0ld6svczyN668
QZ5JLkXChbRXG1w/JFmH/kjKiYpN0mMHhaIWN3wa7RveH8X+CamGS6r4wNFP
wR8Na/uUJ4yH8YUsbq8fEk2TD8MKZrBiWTL1ut56G1SoUqlMfUZYuNh5M/Zh
j6TT0osckVBN77nz26AOIeb1irDfq5MPjbxGWJPONm+NW5hIBvkHzID4IAs+
dzBB1lhgvp5Ck7pIVuysDgt6KhDFYTcqqtUpRPI0g2EC3tQB2bKLlZqlWHQK
0VqMZsRWdXiIe5SYdaKvSdTBpEabjaLZqu36veEhvMYXqugx3jSPvPN6A2O4
VgAKNURvv0gl12mzY8hBJBRxnvS976XCFKaUGpmil5+5WWKA3zUQm8/wAtLa
UhLJuuGVTA4L0s96tf7K62HzB2HY6oqwfBvRnCKp2NRCL4XIZZHBWhkQ4Xff
JU+J8/HubE/PQqCKSbZVJf+vATeWDIbJAT2+jERw3GJsSkLDoYBIT3mkk5YD
FLb+TmlDkaHZhrvjOnA9ECdLIf+o+AXwVwpmozlOyKDMvlSon7mUgehuULrw
6KqCYe686j/6gwgNtcdxMeNAl4gSCGkK5+QaFA24l+8/vbR+COjrZ/176DQF
NxW/pt2KscHGsI6xtmxmVfR6n3jasaWHy5ZkYo0l2pd8hPyKpyU8o0pzvIGS
p0nn1J4UbnfuntD1mWsFY5/pi/HgyLR3gAMvcC3JhCWbzFpRjbh4qsh7UL+U
kySUAzMi5PVyJfCBB7gU9PKVMDxGuJWe6ttl/uqQ64dkV22i/ZBcLfAV7A7U
eKhNMMIvTLHZpvEgGVU61j82aJXSAvH4SaGrJlQS87ctDaE4pZqTn5ov9k1x
APsCCOdf5Rhg4wGsOBYZrDOf2fPYcYFzBM+/J/A5uV5ujzyNsRCSp0Te7c5w
/A+2fmJ7NkCoQPJOoyrnvVdVkV0ZSJTBju/pi8U/3x7aU+X/B1jAqZKiwjsW
hIrvC3wjYgFC8GBEbXNblKZxbI1keYOx6MJUzB2drPePBK4dFQB340+4cfMI
tUEm8a94I0YF0FlUtt+OQpkPQ6/n2Z0sOx0B3kfPXVJtQ41UCZ8u2ozaiG1+
b4vGBgEtMT2noW7AGIJa/wUOGO2I/D11rLIuxoeXmDbv6uVtGiB/joPwzQ02
wTeyZy3duQycjvv5eFgN2n8QgNoIwp8YIIF8dHd7R5SV5sqjI2VUnVuJLKUo
qFRR8iWVevj6XxJDEHH4Xeb8SXk5aYVL37UdaRT40o9yR0dxUO4kDyI5ijmy
mJdSvu/hvtfYyaz4sgsRQscqIoFhNdeBWEweRbjen2MJ0XuR6To3s7Ntd1WN
x1ZIptgXriTKd1zgvMkEeObbl/ILH7CHZIDWO7ZQpC9Wha2Zo2Psz+/z5d81
R2MgEYHq25ZqWaw9FbJTDYZXFzaKTautJdaKQmpUqDJSC43XUwZqPLzcxePQ
+SYsMiwKE6VS2ZhMrV+pKRraSvpcbjcUCUMxWXa4bcbgXay6enJiTPXS2h1D
+TSndlir+C/bDLuySSudF/zQWB/uaLlrx9vjg7rKCjtnMxcTlY1ofU7n2v2M
TRVD0tWNJwP1RiM7Ygt1JVFLHi9Ry3EaSuVaB/mio0Iikd96Wfxz7aYXpgq2
L1ozeBciLXVjwURFvK6W4SAGBTMkKwIo2UG8c4P4cvNujk/NRmxmzpt7YSFM
VrhqB3If1ufUZ2vinEInchkOC6MaAfxgfm/yNEe0bjI6AvmHC12xpWGg3NOG
adwqYIVAPsH31alYmTG8h2JmpTHrpkwhLBzAUdO22157uVeQk7W7i08NAFIo
GNSAG5MsEF/qSvOeQW2RedqBf4pO9LuX0+T5h4lwTHsKYCuZKFCuSHbyzmNg
IMC/PuVTXfEOp0HUqO/sWbKf6vQJB9DIuBi3AoYoTInaxARu4fG/HYPMARRD
c1t24bju+xrZRXHXBdiUOODJJn/yD6V9+OWNaIlftp725gSefWTm14u7lUTV
paJtOWrC4c7AOr7ORulKOWqFi4gXnrrQqhkLhoCBkK+nDFKHOuw+B5+7t3tD
gJZwegvxQf7Tj99YhQ78Ibw+dZW0lY/ZF1dlN5Zlkj3dNVo61N8pLSWQw5Qy
sLPEjC/hiIBn/c3+fvgFGuzbeVPe3yvpvvEwqOqeprZ2QoFGF8lA4jbBZ1VA
LKUF+BURbD3lPEnavHQhONj+pFJyGXjxRLNIhwBcSz8I1WVUBPgj7R1K9OYJ
/kU8bPGaZFAQPOlN8nvG/ll4zSxU7WqPFVViYOTla1PjUjgh/sXbR1GzykZB
qspt7XM3P2HO0L+rHUahUNuYjPOzw5DLDVE1AqU202baoQLL7An+hq0+bfgR
sDrSI1K9TES7RGLTuWtN3ejnNWzS4rgLCOESvNWiheK8oqobF9SCo061OWHa
rxciD6tpIpbLaDanTS82rcvlhBLFnUwoLfTd6MtJIRPXZfYhvcfXl2Rcd/Pf
H+xI5L+uAot8TFqJp2bxbTQ2IImbwxETibpraLSY6rf6Zg07cw/9oG4gb6DL
D4MqoQHRyHhqKayY/Pac/7PMgnmwXGyHbk0SACnVpIlQa1aZqZaI1a+t+ARf
2uHW52bmPjNl1Sq1PGMTM5lnEeJFDjmRzq1Qw7XvLxXuxy0wIzQ1SoltvZNm
EM0iZQRfSig3j5EcKlCq0zoTp5xRJa3pdzqb6EJQ6quQ9h15aXjf8nMnrFtK
o12Y9WrfbOd0LVGqUOLPocvxFZ7Z0fdkAXZTzM8Zc9WOr8oe5E6B8yAefYSp
SD+CQVp+1ERNCSuapQOlXtd4uCLZQR3FSqSr+8fdysAxkOIUKGR8uxehRxD9
BlFfckS8u1/aLsu/Cyzkj4sGnchB/mkfLvaNDxw8+tRzcuZRO/DG5RySLPly
iQawgXQHyCyC6zj+gPHT3EZ13LKInWVSrsc9YJOjj7BENyHMEFBHkB6+m0Jq
UC4Kj1UKYgTf8ZAEZYo/At0baZpanSdCXupQ3IkBmEooxB7orK4+ZNoFcsKm
egRtF0CXkbdA07LaaBolB2wtKl5/RgYGtbMOFq3Yxx1zsbyki2u4xK1Uq+9W
vvY1H3ljDwNmCri+fDxDQIZWiwlKa393CGvX7vfb9HjZemjaidqHqNYBbiod
l8/RcXWdbUkidolHPTNwYBkLdLWiWIAIQ0vReZvTFYM/YXXoiXQvlJZ+7SFf
wbzG8elKiAXKoLSw+V0h8fUhk7xdmgTBkFK823nKtFZlkBOZAtyXViOgtwF+
YNyJVv67wF/0dE3N1oMOig5imFsaDCKhKBEbukpu9Z7srHmsDvRp5cQPil+w
26jG4hzcqqIZeuThEeiirD5LrHzLNV42u3Rb5d7m64aJMZGEvpFhzfSNGCz5
3JA3gDlWxS1uvbqsyB73+hzdTaUX7F+UaAbZdmUGRCh9O7yLLFH7oIAcumW+
kGWTa4euch/f8DF5jbRfv4RJbkRFCTdLHMRViiiT3ZDVbUy/og20W42L1vgr
0ByPVq59eKlL6O5QAumjeZPdIVObEExoEZEI/i8tUq3N5eRMEoNqhPoyDxtt
xeLiR1TdxIMryv7uabxIZWCWWxQxpQTJmnRt5njCtVBqMFnx0TofXYGRAqF0
fpxzIHe2PHoDzuQEaCHKH/jTq1+7pkRuToXn878GMlP5OSL94N4nkvKfA4ez
xmRU7vPni33BkPJHY2ISIDHjwHdp5LWOad+3Qo8StxPuMD7rfKus9LHlXlEt
Guu+tNVJFHlUSi7A7YY9cUnpputBTY9xkeqsjuaS7HxsSaioPfGBq8WDEInR
9hUavsjatFPDUF5M9Rgpk8iJgk/3wY62lARTO5Fu4qs7bm9SNcjy2SM2PZzO
TLMLwR8oNRKW4qs5ZY1E5pOPfZNciVsAdc4A4HU74mL8WS/c5H2z+UqY/gaq
kWnnMGa0w2+erK/kfO952IMiiDL6f61wHt89mcha8q+FIKxGJidAjjGAtGwh
04sjjQYHWfYIyx+rKFg+YUK2jlMIaEpQP4Gqxuehhk6ETGmpxMKqkMN4hgzC
X6LCbLWBqwKtZD4jI4cgVTYPGu3QbstSRgYF6JoEFueFTRusOLXAUmyCYZcS
qG1/GqZzW0GiDXHfxbxwEQEtoZQW+t2Ahy6RyuYi78EV81H1i3gT3bTRjgOG
2IpRWKeSs7kVeDLNSFSnYYAoJRWjjtjx5ZbePmqi5LcwpF8ptwigQzogvJml
kNjR2yfsa2H8PLG+9VbjWXBrKXb4m7eq9xWF1B9UosD/VGsJxcwQOjEm30+M
LlPOKY/hGai277MJsD22CA5nvXfdsOpSKaYkGuj4D9lVu2+srxIoSHKDoLfA
aHH4YGsMcvVznMwwpLcPBiwt1sGEDj39f1nqaSUZ47Jxtj52J3Z9b9nHjO4b
bNFX3tVZf03cbbprtYMLHC4btaF3koz9JU1hwcdBhW7/RwgWiwdCJRnsO2rY
kkAn4y+s1pdHGIwtyW3Yq0OzxV2grXO+Gmg4XIdbYHSUF6eqsr3qV6NrEgJ1
AlwbyYkIRu8ndx3UGHVcwwGBoAWqMu8S3BMmid+zeryDD+0ag+OmxXY5TfVV
g4DasMGLDwkhmWj7gDA5r4cMTJ835rDY5ftPACapg8z4OmUPD9Nhwa33G825
bbcfB8HQfRP/+a+A81Ws8nFmgp0nAZlvGJy2FU3zNvh0c/xciXKczgRXIG7L
TOnQKTQI8+/haopXkQsNWz/Y3T8CGwERkFxUlgYxUFmNa25IQKklgW+QC3Ap
YnVQGjteRUFt6xoxxuZqWqAE2IjeXYa4KZ0BXz1aHZEYZHD2OnxERFgNoP+j
9G1WQbSAvXKqSSUihFd9M8QRa0jvZdlMAVwiJ6czbmCnNbzxl+Dnf8id9Qhz
QISQCngU1sazkZP2xRpsIfFLR7GNA6eNzQ2F2KjnYCN5ilGuIKsh1AKV0ey+
ouzP4R9mlHkxy0q0YqRct/ml73+F6YDE/gcmy7YwucmAlFyA/wfHzEm/6SaM
vHMgwUGxcx+8f5/2EDSjRjFsaFbggX/qepDfznrSF5RnG6pV62Lwvs2cDk9k
KOr8mrHs1Rjex/z1P7w4h77I10n2kjW9Mg93WXeR2/QuGD8ulyEBkBHpNSUb
eiRXgl3tjN8oMqUtSIFWN1Mlyl0modBZ90Jo4XbTo4hz65nbSOKM/tUg7F6O
0aWC1q9k3vb7AfhLRdh84Zc9YDaGQvLBHNgpwqL8aReFliPgx0qb2+RYp1Aw
6jFVk6cQzzbQiBA7HquVhns1jxghzZpMrrkg4tlW6laCw65HaEKu6R1rDZbR
Qwo2xbIzAx8gyujdHF6oz7mcTnL7kxGfq44F/MlBDAq3CEvA5AUK+SsfOxIW
w/PKoQzaYVkB4h8ptZO0zAjB+BLkrjVBxAAZeFWSd6NwWFnuc6cbr61LYL+2
kYqb45abN6WvtITaJ1LjNM/vZWRmxg2rUvSXTz3XUPxTn/LlzAAViQZNP9nP
yMKgYPjp6jHfKKozQabnCS3pRsKtVZi/LjsYmEnQwuQvXlBKZ/++0Tc7Nbnp
suy6HQi9RoGIn+5Rv8WCuYLVVB2Gn1DrMiK1ZeMwgCHwqD7llrq0hK9eNJHj
1zDYan7DYjtbkQDbQcKguCTgBuoKKH3Wd0nRTZB5M2gPAp2U//yAOKICaMbI
eXvxdUdeSH46kHmUyJzCjtx8/30KgWX18BnkJk30Le7y8T9v7Pgk0mixQqii
Uzh/9kUvBb8PvhNxULKjUpUqNPxXsOvrDpTynzCzOTSlliWsXmsS42Gfwtc9
Pi8cV/tsnuzPQ6djG6r77BL7bLetmATI8hBICa8kHoiB409hv1ZJLnO8hQS0
pWL1pv1TbhtD400zIJq93MDpOP8vNd4y3AlJNFIRyKLamAmS9BHx1hRpTEBX
RwZ+BEo29Gko/sJHSAkojbWawblgZbt9QAUoTDUd4Dh6R2jKK92Fy+A6O0W6
wgs7Cpv5L1HqSGKCAi2Q1rMvbshwjxxMz7eWUR5o0SDy93rpwf0HgnB/6Wom
K3m/K/+M533iZ1fKhrYU9Q2LYX0UQXsTqYPHH522Ganh3H/gqst5BEc7RQT3
/T+L5HcYsqNNwNGP2Um/0MJFzhUVTYJmigrasKGZhsZbVwnIgZLqDIbpeqHG
h7qlWyPO9NBTUrEJA5pE8m/ukmy/hx/6ghpoQekOF9C+hvx2Z5JmC0TWHwfk
4OwqqwnCmbRskyYVwlf7Y/bBvbxc+BowY5zowqffA1/SSs0WR/ttWFbqA/DP
NARKYBK3seo1tBENgD8p193y89kdLBolW9uTzhitsmBNRyTfu4v3lq1UP7y4
1iODQc1NAprTeA+mHGqsoCgPl/GqBb3am8bI3bCYT2JytYInoe4ai5gsOpVg
qm+SY82HNPHi1K6pJp7UYAiB8/VmWlrGuaLhdAwp1jcx47/qw1Aieb8Rnpw5
jR5Vlhz+OkPlzP8kLJEdS8BH15nlxiinhS0rGinzrmn+Fzz2CT1zgJobwiin
efun8TpTedfsW3ttCmK3juvpBqvkQLekK8gf+zfyh4gu3EW8N5i/QTLID7Ur
G9wmkp3URhbVhprZWVHCxzVVGIwUYU3Y0c5j06cMUMZvnD8PERzxpRF4lZBO
pOHa+dS5MB2s8qLG8dXfuMU7QOEp9PklsF4tfVTB5VtHGHCdqanAtxUysP/6
2baBXkwAybZt0nuwtk6CvWonVtLqNVgAM4RhDV56xLCoC1knk7R0/9YLs/0J
PrX6XgcM8otmLJyp8Rh3CZ0i7KtWGJvCagccoK3+2KDTq1ci1ajlBS8LojE8
IGac7jR4smwxYQF6wceVBm+krLWI899dYJ0y4pmC4/yh+L5S6SXFQ2vQpDph
cjWjAm43ST0CvKlirPxYcgSGPYMhg3wn6oK9nPS/PqcGiHBHf/1+fHPWyiHu
lNdopCoiiZzGyQwL6MU7Hl5MrDI6jLJRwYsAHlnduar7nqM0q+hBq9R43R7Y
+2aWo+84rmI4wCd4PWmb8mLSMzI8KJDQWWoM8JtKbWIuxAI99SE0VOqMRZcr
pUBYBNtQMYkqfZMUZtUL7x8m+Kuu4H6oSZ80HFd5j82zBAXZyitrr2O7vPNM
YCrgXgXugfmBJapCY3sBD0HlpQrZSl61BKoMuXJ9AlphhOvMPD9dylqdjf4y
KFG1fuO6FD3Luyor+UIjiFukLiXl3Tw25or6sFUYK+X8xAYoTVdVFdV00qQS
waYj4O6MMsvfCcdxCS88zH/Qzs1eRCpX9TZ50bD2khrRAlLd2Ai8hed0shpy
oyarauCYZmualcCpi9omSBDtcFNE3s+0h1ulUVsSL4jQwFsPegezY7bTx7oS
iBnj3CO5TJiVIj91CJWk0/GrjvpFjRJjA256CNXZsGtxH5mQHPaQyVbJxB0J
hSZEgXVj0lxJ/90rxNss0ETHM8cQfj+JNHigv9UGvM41ne9uErF9cdJCWhAx
5Zw/gQ6bz45lTG2Jjbz2IGFmtdboW+040nkjKQI8thESIF8pG9ByF3CoRibF
5DaSY8wbg53kLZ+g61GsIbCheRR3ttoOLRHjWGW3WLdLElCqGBJQVUUNTQ9l
c97199MJ2J544/220HUXExYDKSAeuAgAVxha2qyIyizgDBpB0KmFfkb3YZtP
pFC1tX/oypOCcrXdr6x2OPnryge4cu/SktaP3UqN9fPzwgFuk84PH981Bo4D
kCKRiYvPIdeR1gi9yO6ilvBnvnG5/1/xZIVq0+64VVVKCoYf2aTlcjUqyYB7
VJmmPIoLS14ehkM/b6ChxrGBszl66U6YumWFFS6rp2zlJmQriJhhIzYQ7ZHN
XGo7k7jGEoH71vHRtWvHpR9fsKqKOnmUEfbk5xiDIxqa9UQmzhGE/ckDR5oT
zhq3yQLXjJyuYiZWM18eWB9qgI/Z6NMdklLZ3rm79cuDY5So+cLicsiXqiil
TgVnQ9YpxH9ta+XsJ6JSG9fX2NwiewQOYIYauPuqBc/bjUyrNVHvkHuU8w4G
SmXElGiaY4v3o+RRPygHli91cfHIPVeN2WvpF3kREjhXcnA7+hAvWjGQWXcY
ghGgH6EZFtiVisYddUvqura6RNv4nD2Gmw2iJSo+NjuHU/2fQIfJ4F8cEjBO
6UZeDzaoLobReOqW+17mlJsSi6yP/UxP0jDsTrBrY6WCDa3crFv+/QFfTASk
mO3+CKfXD5LSttHOFQuIpT8Dx5zLdEhBohumTVFw3qQOPp7FCKL1IizL93w4
7xgzZ5zRFFOV2nP9/oy0sSYeiXLLYp8cz6r6Cqjd/U4Dp2q3uMprQBZPYJhL
exeEg9D/RWEfzT48S0Ur6VzuiRDQoJMn0F/YgZzfURQ2o+70sxTj+/6JbBN0
nIqmuBrE3Wm4SkloUzXRiQR+oqMk1ni7M1gIGRIW95OPuCCt7hwFTbLMaYBY
4R3LPxuqe2yEikNA5KpwKQuj/y4cLfjKRSQBBbBOyPRfXvloVTFSEukKgpoT
zmq/UuJ+5LO1Sb+/KI3Jnh2WF83PbsE8RijrTwDX2xWZnSKUyxtnf2phX2Px
0RmIKbj9Gfin2AWC8FYRHHGBviqffvOwfSvjBFPj6Tsd/SCavhBFvW6dAkB1
DmYCvIBKUDdOO4mFrZg0SChNn52ypXK7j7GKv4TvX4hksSmYImbrJPgdCxsY
JoOmjUsvIc0B9HbZsomMah9L/kH1tsHBjLuM0nQUlWFkBBXYcg2cFBw3YSWR
KvopjoMUozmVxHCRuv3v3bhATbJzQaX2y67RXU8gKSp0puz0fyb4LIr3hXuw
oKr9QbPxGdaSlxOoOZrgDx3eU+EzkCJfzR8DLAoV+uJNeNvtIqHzQ72Rbuy7
dkc94gMue6LkddcecuEaatbY/YlQs0AsHUQPPFoepQ24e0j+kINRAFLFfSX9
EoazA2X+DUJb2fF1n7VOg1DUUT74K8SaXI/H/kjPwiBGxrFbH3PwuHSJ6alN
Fsz+lIAooN4/iUt4DTr+hSj1z19ZnRva99ZgubbSeZQHkw4RUXKyuUzeO6sv
mpt1cYqRFaRwABUA7C+HjF1He+UkRHIRg/cLvivcjMZsusJL+JIpFSnCPHfx
qkpQW/XntrxJD8lcoj5oSV16CdpMlagoKO3NG5jXEXTaXA5tmQf4em1N0Fdq
fWXvRks5dnHM2+HcZYHuwiSrUFpiIemM4sF5v3DsI8NxAyDuClU8nJJ8NUdY
csf9GVkNUc+tcFzWlsWBGAnlElbh6BHLyRoePi/WVT6nRwTd5nhAoH/vBLT4
eYtGnkD+w2v0mHcmty6t+ssgrDZga7d5lYBVKPaFqRPzzNDXR9h5mYY++TAo
OZAyrc6ehS84VkrxJnz2h1FyiA32+ukqBHfFL8sIkPKzmQlgRQ/wkuG380NS
Dx50HK0j1ddGyiAueOewBKsNh17EMlAjjKEzDrSvmsL6YPMxxH2tDM9o9QmY
oJnZNxuTu1irJ/e3vYQfE+VcuTN3+FpsPey4aBz5tvk21AP6g5yfKIqmL3Xs
4EIQ4c56EdCQlCwQLEbylZuXdEs8Tzir9ofAT3abGI8MSKLOjPcbGhU+V/Li
DsNIBRAdtcsfGYGUKcfvJ+jpYJBScGCho8fazF4Eovf3hJHNxYQBEIqidIOn
ySXeHjJeDD1wmqnMbXFU+wuB/Dk4a8HM1+2nojy72mpyIDLPzqhELb36Uy6v
iSXZg/rkCKrIQQcxbgmq36fV8StvnLvJ8AU3aQkM6hMwZQ5/8yc8sTfn+kYz
fODfGCMfq4OEXkqjvhZtSkU5jLz30UcE7RZhy+NrmqzUlBq20f9gtO1x9TYC
xO7bwOuu8Qp15opftT8PNG8QQq0fGEIkJ41UjpkScK7Go42xvHLWuzH2XKUR
gvBYplPIBWpulhL3eKakvEGaOH6YrddTWxq580jp/kVJ1mv1rmrM45AwrCVw
q36qknD6Bc5o+AXQs54uNmA6tn97ZO4oArRaRr/XE3tCAXBYWb+ogF7pvuce
0qb6VqZZMz+n0lF1d20qQ8TYZBKoNVWXBve2jCQd8aMQ9vs+Aff4wuUgw4Qd
PRr7puCgV1pGPudOb8X4VO6NSEGwTQ0XWbN0S0j3rWZyHYUYNqgb7Zlt9pco
Ur2OAKAepFrfv8izA01NKASYTRS8EtWs0rl9P48Fc/XXGsloGNMlSe10DLcY
Wq4J+U0BMxtxlIDFVNHAaXE0DJS0i/3k7i1fbzbQWtm37U5UBic7/v+kdG92
1xouQBEx6ZTb27AnKUrPjaYXnyxmgRyMs8QCOB9kh5ldpsavt5cjOL3iD1kv
ZYpeXvIWAY87LdosNA9uVA39wms+ITWnG/PPH7Wq8oFAEaf/T6HAiAjOrsbC
iMpeeQAVu0x/jt+kslZVTmxbeY8Uw4+lJqUjgeg4hGE3ByjvhVvuH8KdNaC3
zo0aqKjlVWTl1Wd5O2edNFAFoxv/WKhwPIsxJaGwUbFvSH+aMiBoEfaA8dDJ
pfM2SJTCscR0FbubAx7O9zt0cx2BZSktSP6vd3ShtDZNtOccPb7GkyFxrRjL
wT+w1FZiEDKN0DgQuoA1DBdXLr1JKqql/3vfumbQ1ScoR/PjPX6ilEuu+oIL
ZlOwY+epYfVZaPVBrK4gy3b1vsmQU4hibAlghwNbh05dkSaUR4qmuB5VkMeL
lDtcodsNd5RxPKdETm39KGOuGZRpzxEm2XJtDYnr++q3KDJ0xSR9/2FiV8Ex
BhWa6UBfvD9xpBt573QAKVoy9HQZKZRYl+fHIeDK/wxPRRwgtzo7Ay9bTacD
Kt8bEvAoU9paZIECezh32nf7v75/+w9hBcr6Oa2C9psGvUMkmJrN4TUOX3Fh
vneBGbGUCROeG2qGmo/y8NaLu8L+9ujAuHOnf8WPI1w5lg0hgcDkIop8c3RO
soXEH2CMjfIaDM5RTtbFmK/aY5ZpespDrEHc3UDWRWeNXPaae1QAn0y+bOTh
jEuG4GmC4kQOsC6AtQNeXZDlnUdJnZ+u3uAEOQH8sgH4Ne1CNhZM2p8gwyi4
YsQCevMPawr3IwkCGnpZlXZye+Wx4lSCeHTE8dZa+obJC8KLZhGSwDOn0d8/
4wGw0E2wK16p5o2RGjbsCbwpll0TGb22VexxPgDNyQddDyCKqDiX5KIRwotw
/fyWhGQbLlW0uAv+YRawsjhJvsowveZQEKSnoT6PrCt2lvqH+BS1FjAPHRNy
7so85MaUCQaJyyVTLzLVhAPAjkDQ8O7ji9AZS9lKq/5nxAayXPtQ2UsiG7Zv
lHVlyOKo/9EfNKSrRGHYTkEU2cO83ZlHqhjhrZ0jw9wWYGNL+1bDmVsP3k9j
jcA3IR3MLZC5RwDLv8ciWXjRaUc9EN3G5R2UnJTNj9NRPi9q7bd/sp9S+AlK
DpwxttfNGrL5CSnESo6lQGdpJixgj9dGmzBfww6l9wu5gTTP4jaAc71Ngp+w
F3R2BySJJuvj5uw5kf0SVv0OpM+WJ/I42yvhWW8zaUeosgnLc0Dyi2jS/XHs
FfMh4aPH4qW3u3ABq9uFgsTyJGvAA0GRzU9rrTjoNG25icok9nIUg7bf9lC/
GreXByRJ2Pxpjvi193XNxG9aywmyolKOnM3g6LycXv9hJiQjjcGRVxqGj7Ve
0Sx2xJ+uyqm6iHXa+MTeVPK2U9OiqO7HsFpPCVEC+W1nYBvkKDdnQeoJo1or
K4X3jyZimnU3jjZqL7DV12O87IzD6Byq1vhMEo9RsB6QgM1rdys1kUsCfs39
IfuBJlp1U12BokzLZaN2fX0fsMwdBvQS+XNINVjxq1zHZ8W5E+BE0mPcPWgu
aFUMbjq80nXqMT11t3ciChfYJedQWpf2HOtutDIC454rDnn6ASfN0HhBA5WK
KMRjOhu45JKqunzIzrOCmfIwsdL3+TNuy0uDKRdarXLr5265p4GbcxxSLtQG
GqtCJ357qDuDcRRMbH/lVURpbkWIOhSkK1AGk5mah6tsywMgYwkbflr02mg7
P4RgVV0aG3Rze03CyAqj0ea2Q+MXIVEi/gKa3kYdGK+SpaKNHCI5LpPfrabL
HSu3JIn0FFZdIPw8aV3d3nCQ+VGT3+2nbBelhr+FaVcrbBZFjr/e7mMHQpuc
BdS+yGSc+s97avNO4TQO+t6zMNichgGI2XB95CMlXHI8BIvSKVwDWdu7UfEi
N4PRhO6/XIoiiCn8aug845QEYECB22KBUayKEGaOVyRswELtNlo6sDRYLdRb
bqTmG8tHmjzgxGQEi00+U1lMMos8RUlf61a5LyxCEsvQOa35dR98zuRvoiyO
UlPDjZlDSl+yeO41fS52LHVf1HmzcIsGZioWNYM4PPXnKyorBnueEDOde7Bm
4EubGW8rqhGZZSWkYMob15uP6dP6jOllf92PGGfDZ3T2jjZyLW3fjaaXk49/
zvctMVTZps5sNIYVxqpJPzJFQ5kLbtO52mJE7MzMP4dAl6345wcf+RmNrgsf
UQoVuuJZKJDuS6+gaZY5WbtEO+a0IVECPuaMZLiei1Pkj6Is+5yzjZcjXYbt
xXjl8VGRT72Nr2gj0/GcIwc5R8aLN/dhUybpMaCQM+/cXKYgzroAhL8r1C6X
w2Y1njZVu8K9kB4IDkblLA6ANBK1Wyu2Te8Rb31veZXcMCrK2h/IcT1oUraZ
xymEArV7i8+l8nj1cPfK9PJbZJrmaUHpJjv7a40Dgj+8Z+S9s3CmRn5hcTDh
8MZzmJ4i0jMai9YqGHIWQQofHwPtkDTpT2OltMH7G3CA2pVifz3BZDvCAsV2
MnG32zHuKiY5yxPd0wnnf85mvZgpwM4Mim21qbWUA61pryuEW6IVmfArtNyW
zVVVnRpuU0BQ2aR0J+QgmDqRCZPOjYEZAiVylgElUJLXuQoQTzso9Mk6Bwla
H0O7DBjHkkEdkxjfaymSehutNgO0sQANsaXxZdsyfFlYGjHmQa8E+wpfR9Fk
IdP/JsrSITk2IrJlU7Ty62frsrrC+4gkAB0AS77n+mtCqQ+ObhoUxPRIM1dg
LrI9dA2HHLgIstk3Kc3KrpzAu5VWyAFSKothlJd6HxUUV3cP2T4qi1lldTvy
eIBDMITk/SbwCYQtlMAaf7S7wEQ9DOr5MtDRSx4dfq+i3B4M+NW1B8SKH/Wn
zpdYVuxYhyUZTVCocsmPCvKrbJcHjfrtNNtWDM9tmYu7nGzkLAgipqOvwG9/
5PRPlPpGXheg7t5liyNyhJmv/+u0erW5JOZqj5ZEszUgz2QrjOah+MLGhoIs
5pAJRmXg5JWT1jK5MX0iZshTdwQp+vRQgg5BxJFHbFVtXT7wsjTZXHcnxkEY
TBsNjqI0s2DzlIIyrVUL0owBRGTxSGJ7yNHwX99etdl+gr7GfTMDUt1jxeIo
FBjR0latuAgIL1eAciN6CzgQIyBPlNvHIkTo61B56YUtc7S/Q9eJsopgtlAu
Zh/j7W9lZc1ngi1wpMHsOhEuhzb60SU491Xi9ZihtO86ONusqRO5Zu0jQtMV
w0Xr+ySJtXOz2aL+/tXH6nT0fORIbc3W+jNciFKLJC5MQtPR2KKxDjrejK2J
mUpcCdN9SwjT6SxS4caSkDcAd6DuoZQRjtE85FERHagSfm7f9CLf7yQn5rWY
4YQP3AbvtDG4adLBf8Ee7+u+BggOOWH9RtApkL6vTWxgoP5UJe1ClE8wrMqr
2QA5bMuUCieAVUW/jV61MyUCMDXBKIMEkq1z7C8Ud58ADQ4lyxCyMPj2M+my
LqdLY7/ffTpi3UQhZXXAyNyxwwnPz5m4oVRKVXA+97r/i5yIWoU5IianjoRF
3/fjQ0if7zsv7pk+hkOfwxoruV+UC0meSwVFXhUB9iTUA3dTds7ay4DR5KuD
ZzpBFzsssM6xXsYLQ1G7JIXbnp4niRP8mczrwkPSRWrWj92JUiG7mLSn0x5Y
6c934IPFEPl0WzWbeziHcStiNMxzooyHiyHCNKn7cbVXNaR/fnc+XtmFAQ3c
kKfy76srFYFjaUIr27U0WTgmzixcXDM//qaSB/GVq0z3NP6fImXvMup6vluh
X1MZydEcd7Xtmd2qcBiGnthDLOGRYYzhlqVym9q7r0GAlemPquDoCOgDYuv4
HIYUy0/g1AzaCht4txuzOjnj1U7J2p3e5Ew6e5+gzChT+yvaqylrJIreRaHd
/LTW0vIBuSsQZ+78wgWs764DaOovxGJVXbXZ4ZjWR3sBAbDtuhNyzh0tVWP4
cBxIB6/oDFfr1eLqJXyZSFWf89r4azpYXycBL5ViWJv4agzt/goPMU1tQXuS
oZrxdxzYsXYmglvYgiaJYCBPYiR4qoDLAXEYXyLp4Fe3cIRlqOvIzzkPCCFx
aKZ0VkLmUQZ23qUJvKHP1Y4yi/cgxd7G1uk61dAs8Pizk26WaZqRsVR51yDC
CewPLzQp5bdPL2906Lp269PUaQLvP7mjX9x+Cvj3RY5ukmsyZ4qSx1lfdDYY
Wbo5zyKL7v65noVqo/J9hPu7GdSHgwPR/Yhmz7fnOxC7W1F4HRLB+41iwTuq
t+OBUaafmadm9aCVhhtSpl/EC+KpYIx0FNAuz7lHJZBQBdbueAAWyeW2Bspa
0E09qtqK27+G2Y0QnyKqPyPdP+LwjI05mJVhbkSTNLJucfVy4JwAaiOkhWjr
km8UVvt5oeVHDuwEUp7bnN3tz2i7Bjq0XK0t6HdVRp1F6mSdJR+beaYMYq1w
sDNjtAPMJkKi+4BLScx1zyhr3orv5oRrJ5WRftwuqifggHrRpdKLt3gVHeVg
y3aSGMDKEaw57Z6zpgYxvGnnl8ZwQC6zxpeX+WvUAApN8uL53eogxUO9cpXw
i3aSaDoYuUEqVult3qF5CT9Mw0gEPv6XC9sHlGriGXvoftXy1+yCClV+OT6A
s9wEVSagIyK/bNdQ5mfkCKfCK7Bv/fB9P4xcYYakNZeDreRcSJXef9COGmUH
GRAHBGPnDMzXrY4uW7OHTWUX8zNHI6kgwRvkuq63SOzlX8/V8M7PTu5/7eWf
1WGS1UqoppnPZedPwZT4g1o6jcwd78/XtCEQEIFhqjgEvXfXIbRp7AwPeEyT
/mcOLmhBJwm8Vj7I/qlgEdTPPF8PjLNMLLBKP9kJqAI+/MYh/vr8VZlsrlQY
g8Yh4/GYCcBkkNL1uEELUMg+K4/TC5JctTSEfVIM1Pg917Cw+6grcS6AEf88
cA9f7frvgljBd30dII1xufhrH09MV4CfBz2at6Bda24g8ETiDzpIKzJStE5R
38EzEsKULcSNZxDYbNZFrALATmepjKX/BpHFZ6wZxNH7aCU/LrPXlUEIXkhr
iqF2Dy5/mLg0XZiexzVcOXZtxPRXXJn4UG9BzMWbSUWhFlg5/DOIhUvPLqRv
L6LD+Cl8WfTYDYnRzlhyF3wIoKGiBrII2n4qnbrg5s+yl+h4kcb34BHk43Vd
GC/f48s6HBy1klQqZ+fchUN2fC3Y/DgN2CB+8qaSAyrAOfQqk3Ov6vyN+oYS
dg6cWirNhyVBF43K/D2hOZQ2Pl4GNn7HSLh96WPuOY0O43XnSPzO9IksQ8aT
3pEyLNRzDNGolln6Dx09ecvy+7H0Ll07EUiyVosPN7p8NACUwY9WACN+qZKp
AIjdcjsLZ6hssUwDbnkznNi4dKS3JsxJ8UUkmulC8WEIpglBE+4SLNXUCTXi
zwnrhCvp1xj0nSTHf2a7arwd+WD+ZaGY1XtOWDP36EcrqxFFiNhGGAMFyaam
XEPebf7mYyXVuycgquZUGBRcoyW4T00lRehB2j5Geg5YNwFhYcI0WrkYeh7V
Z0XRfM5Fx6/yjdMJ0rrxiOf03Fose+XhUQ8F4Jeb+tIEHMYpXdyo6F/1XGMR
aJIE9a3qYXfSikMGVKoTq6uUAs+01dmTJxEfiund6USpaTqZy8vVcb8fBp1M
ZQxRVelxa7tq61CpldwlwsJpXgY+DbwzPpr5XAoLjhTqTWOwbQI/7aUig1qt
ycGe75nnmBmrmYljxDgxzU+Htbn8wjl8SMeJmq+xSvhsdT2MaNSU51LnIOfz
OV/LRmqFG4C1aRigUwXXsxhYHR1Y1GX15zhRoXsBB2VMecJzYE+Mb9VUEWno
eKE6x3dpeM56LRywgq8bmzRGwfMsi1/59FSYnbNw/xhZxKLaOnZOePIyxjbv
fLjBki7Te36rcOjIkEpCf6GzeXaneH4fS9RAClHi4ydl5qOXVBurdkXa9UEz
digDNi7umA8QhSeHnspuE1M4zzc/NInQ+gkX/J0Iv2MlNUyC86DYNGoPCFgA
aS7bLZaQwR9nfQEjvA3D1d6FFSqtEe/xCJjFo5opUVXFYn2NYzPVGj9SQIOt
HdwmZkTFB7tiDzio7+mKssaxZnybJkDdEfSnuaY7JifS+Or7IK6suP28gZ7K
AxMK29/9jmI1OWa9iKviAhGrgU4VgXuz/EyIaEfmjqna/SrhnUZhbYnUO/Az
GwRn07gTZ+8DV24f3cEht0PP9b3N39dTFqrgJbBjnoKuSoEfEAN1T+N+ORjb
eoriELuqVHa/7IaevbQrNzDMfxBCRxoCSc2aLZb2PgJSDd5kURHiiGooSi+I
7p3slmw7C9pgpHafq4V2e+0z6qHxl32fVPzCyZiGhwkhLkw++4u0e8pEek7B
7F8NZAyqKJT1l+yIpwVFEYqT9zkC2FsLcHD4CwU4kgckkuI9sq+7TjAIV9r9
z+hTsjea3htoOG1B3WsplLCDLeWmNykB9xaoEJAxZwulWXFmltSQXNUQjRFj
BPTu4QVFnfvhf8omjX34k7twT4sXbrI2IEsteE7jlxa8LBXuHkssgATgSuUx
wG6oovJqQz5dYMftGUOaLotDR94eR/lS8HZg5+Z2HGxN0w135qGmkk9FKRRP
ackIbyze5a2/lmxT1bPAY9heoViaGFYd4RSDnBGV4ylus93AsKNm7SQO3gwR
TI4bO4aqFmm0LLgqPjObco/iKvmdotvKsV2uPS9uG6G+n3BZVyvDQUdpXLQR
5iUhmBukGqbyH6VdRqCHSuFR9R47jVCUxTKiujD4+VTkTQt134tcn/H6V0RX
teeGHwGLIXs1NFU7Rkc6nV7Q+4ZFgaGEwr+sGE0xYnZ2bkjJwGddKkUWK1U2
4WWAiIkIl6qHnmvi+UDnzPsRWnXJLmztWnumTnewTKjARZ1TsKOmTJh/qSfY
NziaXz95V+Pn9kuJIzupA9jZiTs1Rdjo5gUWmubST9xRmg0p38RwKJnZ4dRy
V9qWZPu6EwU+ox7NRb1ewb8fJOs3VbCFWaHBvhm7HJTyq4sxb81XUJ9lRqfh
Qym+rvvCrKd7sbrqiiVyacyH8TEX/WxBCDuvykMT2Y1fI6TY1t4RXCBIwLVk
UXGAgcokbo4pWcW/PjAjE2j6lMcx9irmq3yJzXLbO68/ZoQFTB3bDjMuVzL+
wviVavAUhA5x/TYZClbdZuSjyS9YXk19EVvSBMaEHLHlVJKgT+3jTPxc1Z9+
YwrPTHad1LV9roaj+zdeYIqmM9xwTfW+UEEhzxceAH1jw6+edIsl7TczKiZX
GKXsqekanjjXtxzJcm1hHbZZwqQhYuYrglt8sVVFQE+VGX2w+Y4adv2tq88u
G1o/PSdkCq3w1hzevpoT2Zim5ivDIx/yvZnDYGSmTfiX/ikrsvgnuuQAezKT
5ZrMtFBG1ezmAzDv/a3jurMV+3UC1gkYorCSZ9t412KOGhQd0pbNdMu8spzb
uIMFZ98lf82LQs437P2Fs/F24kyOcHD/xsKeQxl6HCMK0kgN7Q4evqaKswu2
3iEf82VYfBzNwKX/9jXIG+TytsnyfqJbfhx+bB2+Z1tGH+f7kdgcSSIRgrdT
zMob8X18MLmTzDTwxYCGRBUkwwZI0lnLrcrNHLpSXb3D6LWbQLUHym49QjMh
JpxKOA5JE3hDrH0Fc8Hd82pYIbG05JuuB7xt56aDXxASeCc6SG3fkDnl/rbg
tEdUV413oEasFTtaK/cFiuWcIWckyt7U+bhesnphq+hMxhs/Y3GqqrTwApll
VDbmu/rzOsWsH1hD8XLxHDcCXATwaG7kC3Xo7zvmF0eU3zU/XjaWy0/52JUA
lgFBCuzLVFc8AoLFH4N16h0A/IBQneTlSuDdc2F/keQe3QP6FnZqa0LWQv1T
pzON1Dp0zfT1tx78sJE5sP9Gnp3BI+h1fWBDV+iMn1nVVXYgu2KdUrGbvyl0
b4URsPX3wzehOhygyGQkXsuITzS0F64md8ns8UaaAfWOt9Pspvl8TJO6Y1Ba
NrKChPc30q288thamM5LoUl5JmLWlR2GaL1sh8fCGGNtWJfW6vphzIFTTMz2
F1wJSh0qtjh49kY/pHVw2WpKRtZ0XUvKtr1p1bhSuWjCYJDxm+8VYHy8D1Sm
xV4vf1dKCQUv61RnUzREvRLGU9A9mhFLyYZa6+I2WPRyQFoGClyIFirKsac9
DLjETpPfXkmpYhv4+UrMtm+A0kXYlklHRtBNavdLJNYZIxbDaSDZ82FuJ+RJ
Kzr3fyvcb+fLz1MnIdNHebDpY4Amj6bhLB88KaJOkM2W377uSdfNw/cs6DGV
b7tARs8gmjTGFk/LuELQL3GHmh1Sv8lDJMeNGcFbQTr/fJbe9MW6VIYgp93n
QYKhSJ5vZElfjYc7Nle2NKn/OIKy6BQGQ9uviQfjTCKwTi+OCO19nhQCiHsX
FPTd2FduShcUNcZLAmoxSogst24lWbOGmHNESD9Zy6kpcWX38ngzAqiW24Tr
YF+pURRGVgl/gWmh+uLaW3PUUpOVxiB6dRcvYa1BLychq3Jt4DVfI3FzL8UD
DOoli/N9I9mAr99ZTUZ5C/UXl+IlXXlkpg3Hm1LZjHZPNoTeAzCMAnfmgJD6
sl3GOOmsvikzP5lwYoPT10twtvuXtZviiq7H1Kymnj8oURWpze9YHS886bX/
h81OOVWbCEuF3JH00DWsKLXEc7VYcosBFB7/9OTDBOsiJ+QJTZQ48LXqT2Ct
zjm0Wwei7v9yUeW95PhJqrSPtkBTQDfKKV6ceO5vrrdFh0Uqgpxw71AHMZ5S
i06D6knMb97pc3GvbCC/Tx9yvUASPb/RCiB2BA4g5tzg3v2Om89RLGyVETg5
Cg6+fCesOuWGJ8Wus4YkuI90mdk13AqVrBXnz1L85zFHANi+djSL/Frg/e7s
nMc7mZeVK5LgGlNFhL7QLdcuiw6fT6jBXGtcUG+44TU35pH/VmMcMc2/eXes
Iaik8vPUjE4+vra7AybdlQVuaB6qjn9EN/rn1Fq6RtWC9C8IHcEEzpcoTnYb
Bq9agDDT6SU+IkASX2J0Pgm2i9MMqBq82pZFTtKTAXjdXAOF16vMlyCpafFK
e/kjOZxR4zbywXgAya6oD0YrJdVyPG6mzFxYsT7ojYAQDa+RiHLi+3NIsZsV
DEwtRAKrea9Q7i6wzQTkOM8+8QoWl3gf3vNbM46BZV+LW1B3Uw8y7nhm3AFA
IKdgNao/vewWSm+uuglPPIT4Dc/kCYluFRC4i6yiYgNDcf9sBkWnUSoWSnEZ
ZCyq33fjOF2aZF5X95GIIlkTlD/OEsHk5rPFgrKjqZTkyTj2YvthTN2Ozw1O
JUg6ftmqSrd+WeOGkWwKz1DpUviEE/lOGWl4a3g4cD3k8EAixl2NkSh2R6Wr
ZlsQgXuZaVbJk55pk4nSuWsrRGeCnprL3t13fLgwPUSxp39ZycW5xczZe6/6
xpq6JeJfKG8ZghQ/1XsxBW4rfDgmD7UX/F7ksTvGp2YUNgNL7ZTdwlPRHM8g
TkBMOzWI++pxJsM+LSEItHWafzOM0p+04oC5bwW8khNGeYuGlRRc23EUuDfJ
nqgLZIYmcbIKGt6G+a+Tm1R+f6kGdc43W2sEB5eMUJVFqH2ET9dElCKoVUsy
LSWqNFjpD0/yNd6fYfkf/+KhCg3HMH27clm1MIGqoHuaqnvoaTfgu/afSQIZ
E3tpu08uwNiOGAmaoS0WMCsuqqBipKMTJZkwmgwtXep9q+NN9WXfg3X1V/Uy
x3aLzshamD8cjgMlV4Pb73kJ7bWH8ls/7DW9gct3BhG3g69jIacxku1QwAyR
zHb3sWH8uYsvoDEMCD0kyjjksnkY9mM9SfSqS1ME+6DjqVGUfbFz+9FlJw3I
q55eo9TkYcWB3AihL8AEcBzl7GwbRzNXagaOVAw0J1SobnxA58JHZl7B98pI
ISnRT4Yd8g7ZDXFNyLNBmn4SxbEl4F82QZlCJmqr64rf3gyL8BVuc3yny3Gs
NmDkQPuBhaQBNmBaPionph/j93TvfC3WdW+ypqBRCw2ad7qmu1Yqh08edg7g
YU6nhVJ4JaUwIg2FKOOKLONDfy+tIaC0/bmwx5PL25gz8HE6s9xTCZ0gqPv8
YjUJMaqc71n+2NErqeTjc4xESFgIydf7n0O6UQ/M8A3YK5310PzU63MU/UMj
xsnLp7tK/lb6fLKBW93VhzphETsZhLA2Q4LAJiQiJfB/hIWJSRpc9u1v1ini
fP6dFuGVhgWCdgKPSQawAXmlBmgGXbJGON1ZMrOk44vokEY2uU78UEQ+mjql
pJRwiOM6z7MibL6K5ix+GstQmQO0UKqdFi3x5XhQ3CFBZx3rouQQ4PbhUNHy
iFfDYFIdDSgijqu6+oeN5s90+h/h1fRqiIrDvF6R2uwdC5BGJpq+jyihIKKC
EyY8/+2F1I5RrGkRy2bNFY8GSQOyk9v0kwp1CeimbKm8mlMG6K3BeiVG3CkP
DnHnq4YuqdkiB5Cq13ZJjcCn7zq95tCaT5vJ317nv3DU4xhh8SYUOoNpXcvm
ALY9sqRFy8CcevihS7HLcXQFYw06PxVdqM49l/s6Mhxx6oxjY8BpTbGHBkof
8dWRT47BqQOUqBG5cJEXj7mRuTEDlG73woj6yVhAKNNlhoyIOqUm2okS9oBO
PFsD0bHn+dA+jw+CuD3wbBkkTr4RZUUWyiCpqxFw5YDzGAGou9IXdGPXAFwc
+QCZw37qcx30k8+DyBl4qRbVSDKUJoXA2S6Ww0wDbmnanAhsD+Vn/5d+R4fP
ylt6tjfJwG+890gyjzTYH3AYDolxvwd2g4ffd3IUj0qh9ljpcLcaHwRsJMpE
/0jKwJ3Dq/M7CzggghzIJAnsC5hlDBRxWH1or/LCyfqG15ccpSWEsQyZHnXd
JofHXJ+vAjtMNbMDko8mq8LsrlDImxW22gJwXmXW4e7ch4G3w61wXIFRODjE
OiWd547usmtpBACAqx+RUzhkzbZXekBZKm+bUxdX08JqoA2el1ROEWgmiagt
mgatH1/9d4UCybNCYWyAoNcNQ5bY+uLTWfyGSFzd5+P6vmZbMwa+YCJo2Akq
yPJZn2J6/plqib4zOfhRR/bWgSR30JKnTaShovFn+5Scmh8IaUW8q0yC4+cJ
PLlCm54O37cHWSun9FnLyv0ajoJyaOpRBRrCdFOSBho5dJCceFvSRtbX4gkx
RhUHOKNZ3/zORpL8Y5+irjYqOnZxUaANSUqy+n43dfFTL1c7K958xWWWaCzD
fFznX4dZwXwxQbgyTTjncudXr3hLY1n8RTQKVzWujDyg8Se4mSNymhBmbHnD
gs1Gq3X0zAE8P/wQKIT9nrXLh+vOKQHD9rMgqS20KipWcAAez+KQM7laiJlf
2XaUqSozdARVEoK0yybRTTcP6aUp1jLXKpbN0/+EzjET2/t1bMWpM4/JTlfU
fnvs3Rg7w7y7K8qXaaIofNc5gW/hS8E6YUm/xIGMGXxPWfA0xd7aw6ib7/ob
TRGnPXiOaR2znCBkooB+RXuEOjh88Z5qV1pxm4hy8ImnSUeXxlskTZaWeZ9J
JJ5iw+5CNkYu7kI5bo7GQ4pVorJtNVHnJtVJ9yqEYfi7njHjXFUQeIM3uR9O
VKbP/ET4cmjd3r17T2X0gIqZb09sskg/ZwdrgRpnrMs5c5wm9dScwoykZIWr
W/jNRf84mcPes5rUkgjcQD0OkyO5+NLbDpSaNx/PZkb0b/3nmClJWDdc5xJ9
ERsnzCG7qpSGg8IT0vui+9nJlUtc8tvF60uHGOHksW28i5p6a902eNZT9Zdg
bPcuYYtnc9R+FrD8n5Y0zji2xShBfFXKa3i79YcYvKxA0Rn+/xa8XV5D5wYX
cg1JEY3ZY3qWseOvGfzEQCn+JvTTbBxz/wdnbpvQUdo9cYQ+bbW8YbuIbZOm
Y0bpQYypim/112BWhk+0y23+/fKdgAA979noVRGp4X35OCBLY6CsJ5CEFlph
1mt3ll3DuzYHFu0w7hNUu79jyAHUW3d+G6Bm3g0omQ6ktEVTyHVHmdXIdAAk
NzW/qrRtH0/iU9poRgzUzHuoDbF9WkFQIPYL48xyVse4tGmcAUAalsF5tgHa
kaYza8GS0AcCO9KwXkOwmG0veaZ9pshsNeIGaygVEQVb8mupl+XfeI7L+vrn
DgSs+l5TZrdX2ek38XnLirRhGxTb+ZL8JweQnyXtCvQv6/UEQmK2cAJA2lFV
I/DLnwTRtBj9i3oa9gA6+Aom+j79ZgeaGViaR22KoUkCXS03nFK1OO4e3YVV
4Azxa1x89OncvUZiKZphfC3WXj4zeEgzOz/39JQ3c9hi/c2Xfacm0fX6PcWn
MjQ1Jh8G8F8JE95FXZYoJ8f11mmI04bQS9LSXVuagioDhbfHP5XJqtUMr62m
ZGSmlQogWghCS8MXWCXhROSjzqd/Wp34QtBrn5Hlm5vvWPowapF5h+4l/0VF
ghjU9KkvFLyGDZGlRCYfHY+E6kmbvpP9+VkKzk0idE+xNq6W7eizzUjvjpsQ
/a5AIn9YZD6QngHzMIEU0mrMIasA2pjrYKGY0bLu+4+sFtvju3w4+oGdBXNE
+27e8kMJiBShSQNVa6UDCDbxttlLhtI8wv/mlGvqmeizhJ42UoPCnWSp3JD2
tv7jXZ+25e6B2aDZDSj3lgMqF+J7UWZ1ti3UTdes5+dVz+lVUz/mMiTo2mvZ
395fRIUr0UUN5dHVg3MtSjUwVBmTevIDPilWNReEbRgHl0cOPynmokeIiluW
et823eZWwhG8/WjDZ6njaoGzkVy8ssWsnTtELHNocfWXqFjkqovH72bo5Bak
oOC72ypS/aDOBYuVDaLkPbbr5/ZV9MFPoEt/AdxHBiOzzJvQvr9IERNurSYQ
UPvaj43pb96IRSUNIueWzyUaRyckrS2wz4jJi37OO/E4Ygz8P5wJDICKMPit
okrFvSnXvhh5Q6tWIBARBSW7vFn67qpsjDN4FWXZytnn87QRrc3BdIyhiZ9+
16mW+FZ1/mqNZHoVJskQwpvVtYWfxKoSRWqHxiQV0SUhCwHugHVk88i5Ha7P
rkDcxSM+K0jFqaOqi3nD+47KzmukpEg4QqG8rkXDLsYbkhKOJ7z9M+pT7+N8
+PS4C5aOxEZv0F+XMLtUugvFiPOGjSyqy6sCaR1FLMfZcvFLJLUUyPUV2hB+
jytOhTf2We91uwB9RmQ39v0dleY+ChbXKgSVUma3MtE4WGnXdGjIeWF4fVXv
4D85tTn7G1tlmAke3WbPGUk9YXpKK2uwjqBIQu3fcyV0PCKSK3Ezi9RTApgr
iyi9YNkLyWYzcUwIZIjfIXPapAsyYxX2RelLVMdGp369jXESRiqEUEJoNbrR
KdrZfkfWXsIjTPg1MrDFIezjDKDTq3jDEHJI0X0OLqZfhHjQCVHwOMa5Ojtf
zSWRRurqJQmfBbhME4FHPE6ls7P6Nzmx+76u7muxd12TCriGGFtVl9nlFrOS
n0jpaSkcY9BOsaSwvHn5nDpsho3v6UUozh1AYoF0jpTV38db6JZWy2bu9eLU
TBVt4ZLvBsiKd1xK5bpd06BNK9TsuBKXeW2PtqAF44oZhjwFyYol3Asi2dqh
SSlH1jGN520ml1VNAq5x9uE1BjWVFXsHqN2lz126iR9Ad1hLULzihdeCtr2l
/VflMNdLiJqDSPoCxbULLQi2IyJFwDHHfmlYpdysd1m12QJhjNSZ6O69+obq
131wttBIknjIs2svjfQVYKBNfdkToG/o5Rl6lviW3PeIGvnfbroymJtE3xKq
ktLkuJlzJV0hp/KZAaI0KqZDHoDnX9dpS8H0T5JL6brzmOXBT8uG6j1y7Sfi
QTUl/sjRQ5pYxJknX+euLXPREImeB3uQK/khcImcdvJZCseHVDX3RM3igU4j
uWCQxDC9tIol8X1oSv3uJxqPrSVBdCDI6gKuHjUaIxxNO2BkxUJUVxaor7uI
E81z4UNYyZRh8CdNOVeCjPRmsIKq11F44GpSznoPkEBbGxLAwYUvMFROJddW
JteLUnVJWfNos3QBix1mKigQ39x4FCvQzoGQJFMkvzYlnDGmOiOE/Norc0dO
ICnMItgh6PFJ3CtUmkwAj3f6YfZ47vu4oVvvElPmWJva581nHDnrkG0R5ato
gVmmadeBJpRlgWy6/kBneGv5Jn0HMrpi2KmwTfyhsTqmpMERZb3JjU6pBOJU
FUCkbZri2PAgfu0vuLguzQdlNAL8R/2xd9eYbTFejbqAe2j3C0mWNn2Ddd/U
WyL6q+KO6l1CghIMeDssynUybBWQnRt23ZnnLRrS+bBeTMNbczOK6ijqaYuk
q/KZS50QCZgKVVjGHIfc/eotZlmmsIxixKJ+7STy+Coi9F9xxO9z0FtQAYuN
FoPN2FQv7xQ+naBDRfs+3RFoFyfcio8+/+Ht/ke06U1bKIQTFVCXYBTfFtAv
CALL7W94RzsceQjcoct6cVxns1iIzpGB+Vcia2xKTI42medygKShFHOFUlGz
709Uf3rSjNxSpzrPmhBP+ACnrNQYHTiMn+vd+P5Hari/ViVlPrhvXEbA7hyz
Tt8AwwMmGnRyB5qAJw9tFGT/9jCzNDTU4OPwo4XW46QJBIXtCV/Ule0nX4pA
lWqejAiF0c7Ewjmty7e+O0M4q0Zg90CdTjGW22W8L4CoeTAzj50ro6PwjUCG
jizLUrhC7T+DVpjJXZEw9vxOWkuYRHwvMFlXVYYBxDVO/ZIoKZUa3N7HBXdS
6XcAyVYmJTR02FPVqjOy4mYDAUCF4pay6o0rZft/LqJi3fj0DaDLGP6YGURY
XRmkuAOYUOKbelH5lrl2nNmYv6Wxk7fYGdRBfLkssGjU7CcAyefhLvfo+4AE
PjBjEgnWf8T0tKwd4/Q+gQlr23ZaoxiZqxvc9QUd4jMUmXUEmUQRXqbClJnm
cxZwrd4qMojMGaoj9kDdS1n5ZPMC0feCsylRoZZcxO6sNQD/HnjNy2LR6pPc
cPEEYymYflLwo22waBrsc/BOt5DoV1owO0UoCMOxdBLp6VPmw/3Qd/sS8c2K
3PO2scYPASe1pndi9KLDtlNOcTp4cOOFTU/gfgB433qAaEuuTPN+IM6pbDhV
VPi541sgkTDJkBqQsJo6oqrecg3Pzf/O9cwCDNHx87GuZO7ePnLfgw7wUTRP
kyDsXXT3bh2BoP913XNxcauW+8IOJd4NBWHSZfYmzkVEYompboCRFsrvqFTp
J/eP2LYz4mbjZgLUFlIcy/JiQ0tpCFpQHC8ucLYljGuazsvV/CZsrVEnYb8d
k0jzvcitNIIaCZMkV55LbY92VOagGaQ6p+NLdthDB6G+pk/JYSzbJwDUpnun
NIjfvmRxiZ5thP7CoSNIGfg4j7BIb6af02TaGfK4DMWAoT00wzMktC/oJNWK
6/A6nGRF9rdKR1cV2MfhnluEeVo2c8hhj52NAXkF4pXnzXv6WJ2EeZt2gJZC
HyKI8SSWnTy1ybG3aCcE6k8ZJ/nE9sRB/4gETS1AZ5pv24lTrA1ANMIQw2b7
wcHp0aeapgfVgHOJySE/rmJ1BZ1yg9nRa2isB9F588bNoXfei5OUzTQ3sVls
p5EU1mYBr1xMzIX0RJ84/T1y/oImteaPAxNtbFNOcGAiOGGW43SecNvmB3ng
fQhgXPq/2+SNo1mYyi2qN/VnNwdbXeyfd/2BQT2DlTrXRi42iaTBjSQS2WNH
K1iDcJg7vlf+Xo1LPWp0vqQGthuwEDuUGPhzr5Fyys7Bx+ilq+LxWKn3ikRt
/3mxtOgLioS/ZddjGEkx53bnoAgHCjCkRIU7qI29kanjoDtQsLe9I1yE4GJm
uqlf9v7LoS1OVKpmfqyK7D25R9z1E50xdQRetgqyPDQwWIlEVZ2pC2OmQBUS
kXk11+6qhNoGJkGsi02pAEflSo4kC+76OPQ9xfxGWy/T9r5wZaEYfSramUH+
WuKfNA9IBIg4HMN2hCZJrF6jPvSmO2QOx9Ya/ykcoozsVp4t+9pg0/RboLoc
LReQrpISUH39+LQnQd1dTJhyp+bRYUJXFfRxnIwnCewe1mtwYfwWX2eR3Onl
1oJLQw2iwlGjRPqsCN1ENkwnQWxwiR/rkB6nvqx56l7+cIPj6i9hki4jVYXb
klouaM2cgfklpHyFMF2iubTAzOR0HiBPEzGqdGcooYqRCfMKsvNqSpfi553+
8W5thG71PycMkamqg1tki6jd76nmxEwJtEwXgyJs6oQCmS39bcvJL2LluWjj
+mUNxxhBkKbSZs6lH2hlYmc8OJa9KN2X4JYd6V7AFOZYdUzVTPgnOQNMgAlC
vi6qGSYTholA9EtJL39yoX3prgoR1uJHsvJec7tPp3Ko5JxdvUS3Pn5PIAtC
lB+AD5bvRFHeuBKEE6X+JuFzJZ4uZrC+pArv2+xognjMQ6Kkifp+rUm4uFC1
rLzx6lIywPRwCr2DNz+UCScPAd5xGXpgWwMGb40fhlGOfGL1P+HiQo35WS+B
hP0Mbig08Gvqfmc1WlNSp+2ppYLMFLxIAqxo/uR/95ZbnjsEBjlW9oubx9db
/pJ5fNcc0CD/fXV58D6eAAWD0EAQBCe/XCZiNUrtZaRXi2KfvqauSKvrIFhh
FhrdnkXlv896181RTjQOYyf41bxJU3vtoX7XbtfQwYnIAh+1ObmEtvyfKiej
GILIKiSpZk60PNmAkpl1jUyaciBItk4gH3JVmb8Lug0fdMy5rlKq/SnozVoJ
SlA5SHBtb53MaQ5ekDl2FhXKPJ9ME8k7PQw8E8mHgQJkDs6D3A/pGwreAlji
LRbuwmp6IjjN25btunJlIqHaJJ9BHjj6e3UJbtaT+YCVRn56jHQx/EqyPqNV
3ZBEFhGYByAE15MIohzopSepHC0VAHuq+HH7kBafhK1FAhzfJkDcogkNv2tC
pByRI+iQ0iBfTsa7TP4vOkkT7J81VSr3l/9szjfXWm1BgrH8IR/IR19HIVTL
5NwcQGHAmkuF4hwhEZtWc0dIhMnOJEJkePyiBW252qEN3FyhB/MXC9kTpPjC
rX/KnPWzyL4hiVb4Uzq1DUHQ8SqwW+niun85imilRTZ21x5touNis0ItbQ66
ZMZoCjirHssOKwF8MKls3Ba7nUG6l36OcCUZQ/pvKnSDop7Y6iGAEuqvAV5i
2dDUfibyfVdju18C8+H4/BMxculTDplMMMLHVD3MWUMYA39QF6W0F7ty6PEh
xmAlX3unvweaMje+3Xw3C7co5THt/Ut4aOCM93LT141DdASps+CDlUIKoWrs
rXoobO2OU5dI1xI81M35rQCpMF7i+Ht/08IvxhohYb8ejW2ZLWat1Xj67Dy5
dc9LBkBFDIb9kEtSA7lALOICtLl/d1B8IDFWCU0BmsZEB+oLnhkEAOx8zVXc
ZkqkTYa3HaPy8w21gd7BGzDQ9WpWyGrtdWgM0bAe2vQUYR3TywuTy4fGB8x3
YNMiPx01kQCxPgnLCuLp44JzwrlC81i8zgvCk0uLSb18/D2fOjXnn6RCFG3O
UofZIKArFU+YcCHg6AbqGMdu/X0K5SmlKKvY+Sp4ZRRQmT6lqZnLhWBmGKlE
bWPUrngcAmVFGp7rgtHRjN3HS9ZC4IgrzqRF2ziJEpp3S0+pSKgaVWt0oTde
85kDqtlyWzU2qDtXnXUtdk6Tn+O6cKBhnBPtB4qC+XNl90WC0mVQW/TbPE2e
5diVudGSyCSZcXwo+S1OdbiDakg31z6jS03NdpPahItx3u0fI2kgsPhrVHhf
xnQ5Qn09bQ1yrqquuHkeVDvtO6UutHMTzJY5ir3c+jsavEbLioQ9ikltQscP
oBjJiqwPYHdhiLWQ9wbNpsj447fCavxRAEu/ko94SxZ2UtB9qpjTedr17sA6
dP1gNDF6vXQKmFF6vggyFlvIP/+krruv96uIWQh7bFmDNJ1f0H+cETtsVY1h
PdWwBtbsvpasVuwxqOqA4sTW0YWTkhnOjlu+6JqTR4hW2CYa4heQ8R9rl9wQ
P31/fE0YmTs7p9o3sxv+hXlS1JYoyO9usQjk2aIyBCsDyVXYKkfGiayiT/ma
szTKog6FPfqdPYvyNwr3ReRH5QUkwf4lWQqMYmuAV9+yOWEj4hT6yS6zbGJ2
jO8QDoEDawJlbvkx/JEqqkl5EV6JcH8Holn9JCnL/olK2rxeqNFjSRgWbhy6
2lq3UCdaz4rj4OrrfBq7lPFI59zsyabLzUQBTB6KerLNit6PhoQNP2qj58NI
V8ReTorYbTehILhZHkc+1gLkk2mqROIHlJrRPXybisWucwMoFdRhO86j3PI+
6o3QhefbGOiiPekx2AxrLy7y/39Qr5ThHSvtEad3ocZNPj/BvhUIlErlnNyC
nOQAhXIhPDM+0ZPjQG5MjAD6ZuD4IVxY0/lro9dmKFJEFJIx4KmbXoG8Pxja
QGOyZ+0z6RB5Gk9QU2RwNUmjQOJ1JRVl1tW8FD193b+JBi+vU9dj33Ccnjnb
pKAL6Cq1aawTCn+q7lkAgaUEVnFJIxbjyeYLNokxrvE9XSNA/gvfTQNpWczY
uKBipSnQwQLTkjN54Dy7dWrz7+qMmIsNx7JNNj8SeB8Z2I28OLh3wMG2Rp/O
vic2r6A2xVnfW7pCgsVWMAg0OCxyVocer89QvDjlFQWiT+Kr7D60+GYaDIu3
IfJiOKd/SvxJfaZZPmAmr1RpVshiaXnQeuQqWPuVKvg8wIbUW65rO2aRk9lX
j2ShM4qW4v9RMlbw8S8GAB7kvxwTCjtQKEiStVHHsTlp28kauADmr1FC5a4e
PB2vnSIu03fg0FeTii9M/3Hj47qp+zKDd9iUT5SdzlI+9N/eIV5EI69JKMeL
WymD2nq4dIm9g7+ySayiBh6WlW91bWD+rGDkyQ8nhhpKGdwoN2l6czivrttY
l42TsPE/Trvxof3591XzBgSYU64zqhibc7G3SJgu/aD8jresi/iQVSPdXLaQ
AXxF2zNvMcD8dZNooogUiHIsl/GetCJHc7UG6duA0ZcCV9XYkKONOURyVqJD
5iekAFE/QbN1qbjWWKE3heYTQn63MB8mqJVYKcd0OD8nQu3TgbUR7/ycUdnf
gkcDN0kxA//iWRQReCSsfiBjEwyVEpNiodvDMMohrceNOrby4OulhhoQo9D4
1l4WRXteb2GdPxAB2NvKlL/K/dB6iacTn4CjcsQwMSR7TXyDDK8EATOsjwer
LvOWX5r8Fb35xFo+g7zlwnCNW+0F5njoyLD4qMzyazY+h14KuNaMkf5uXEBo
8DcfKb7eZ3iTL5CjIby/I0ttkcZdJVToNGmYDt/DnTDLCX1h9cFMJQ4cBVUN
EMKqExF3O/MF/PQXNlDFjTwzX03uQEPESQVyBvJ7Zcizn2wy/C23/ZOX/66l
s/PXsSVAFl2gg3vLhwpobZfmEojftO20cMG8rum+38vPcibVw3ovuThc2OW9
4cV0xVQoFInjP3jowmfRjF4ch0gCXhlV/lZ/BxV0QiePfKvJERA3cS6a2/vx
ldiDimCBJ0fUmpxVL2BbnX0/zrMjTNg28HnSxxlGEJO0JIN/i8RZZzeOkk8d
pkXtsOOz+CHbYK5PMUCQe89BNBu74/kiXpEKHAh1TTjgTCWBOg0nt1LJMwCl
NL4pt9Lg4kzSLSW4iWWcu2tKgraUDDSolpjIn7aC3gNXF063RSaNPNWqgTMR
nA7Cq+IWzUthKfgmMtJwgwaQi00wQw56KM3G641kZ1x+AE05snLIl9D6nt8s
GhjlRCUhipN5p5mQWHMQgMWrTnndLhHy5rybMTqMDSk0xZpMIKNVJTZwmhnc
ll1re626phzsnvb738I9wJDyOiIxRo3vMxUjNvCgi3ZzIm5YqBc8izaBOCmm
8cwCrg8IAaHNF/vrMy5Y66iyh3H0xgKTH5MUfBbGHe2fdg5ShR8TvotBZgx+
faYw7jA1c58xHwFmUJJ89GIErCdvQ8SJ08YlLY85xvjy0Zs5hk573J/ywkFP
YN5nvLqNYCDUQ0Gu+HuU8/0eWhVzCnAuNP6YReQAxx+1tW4/tWRhAHGyhOLw
a1IU7qMc2pYmCrXggt/nZfhTmnLPgRjK+0nudnEr0xRmgtH/nlMzKMU3Zj7R
55pt323T4MrkzXoCI5fu3QHx+rBKT0v59CKYU/O/BIDqIg1Eaa1zn7mgmaQe
oRO7nPW68xU+eJM6LXQoGEcNOryr5cuVj+iAU2eM3xdnw0PYdijFnN427/tr
Heo2sglmIkxRGefv/eeKgqn3P6VlfBVZS8MWbHEXiyWmE5MQipp0BVtv9izM
aEF0KoedNjphf98xm7HQnupEZLnOpnYtTHByrEDENDoeTurREW8B0TgtOJwR
u28pElJlBTkzV6tH3H1bz9jxt4ukNYuvnTIH4Y8W/bb6wVvGBTBJIkiT+Qa3
Cr5sp7o6PQrOIJi00c4T6G4TLZo8GLCT8UEXhlXfswsxTMSi2fZlGuEI3Lm1
BSvImpM1cg3OksECEhUCKkgtYfau6jFhIV+946eBjC9QPILABP0LD9xLNBNx
2znw4c7FtV+ub2mlf+sTm/X2xwEMnyZRdsxskVrXhD0yxpijKhzaHcfcDgRr
YGAh0zaW7ROW6A6oiUg8Y925C3yNcvbkCpgatHTtzxqjNa4+jM3yhhHiSBW/
dqnWr1l06e0yLN0o/98arshIhZrBXirUmjSLmUSdfARtYEbjb3bsHwiZJMr9
/YTQ5mtPMEyx43tW+ePrwo/lWymzxse0sdsJbNuER2TM7YR8cbvQCz21IC9z
gVXW0MTxDYzT2Igca/CxjVnLkJjdQN/wykSt5Sj3P0GZVZIuxAkcrfgLZWvg
Ao1ydVMVn3UCMd5zokvS3OwcY5VD3MESwcL1w8yMVxfsCs4NopEUVZrPlmAM
TKBqtJwDOFQuwi6bRah7Bd0YvOIJaczN8zw37NWIj/Wq1rpQ/ZQyM3XMswyU
7RKE1Gpq82b6Xa3FpQ5US7MlrSS8dsG4NrLQ7EM05m5sPDe5W6K3vcGMG8Jq
zVIYZzGY11bifa4aU+JtXmnGZgWtDnWr6lTIbhr7k2wFQOutnaFsOh0ur9/g
i7KRgy6MSKV9YAf1J+Yenfg0MY4Et6SSegMKmK63NvH7DXuicCEr+AkIGRXk
f5giUSKHNlGYWhznWXotxPTpvhiDT2fIz7ZX2qeAWEsU6gnURsNqLQHDPQE5
Oxpb04j8MSUIgz0VnxkmD2A4Hs2nRYfqdzhsZ6y1Z9XmG+3PjNH8HbyHkjNg
DJR0l+L/Aw7K0I0xtMsYE6Z92a09YDVCd1wDRCXwlxoReEa7HYm+uGNP0oS7
Xu/50ds5ThBhwB5JH+Z73JaWk2g0IlWCMVLkDpt5Har9c7qHOWA1AQ7gCWps
QfxEb6aSUOgFUmjFsL5aymwSBLC3jKf9tnKmjSQgw9SYnssjRHQ76oyUXZ4t
Owo33/rT0d/4tNspafdf+OLybJk7uYAsTi5dQFEzEC/KVJivk/azrLreAm00
qt0QgOoolHfPZ6FPC41Id+U0jYfP3fuygA6OFtZzG2Yl+TlIMXJIs22ehxy6
dhTChSgXdoVvhNAI5iPTy0lMv06+eDav433tSOrrsSUY6Btjb9cdTBjQiAa7
lWZ4esOSvI/wmYhP6eq+zqx3MpKYQtM7szqKW7xEq+QMn4Z5DbeMEXr7vKd3
+xB+Z2AUOkhH09VSfS2XR4oFQ92dpJJ8irl/CLHPZkVpSW0ahyjazv66CgUV
gc9xAgy5YeDH4dCjzaDIORB7fYmOlU3/pLHC/2IiUFreCPNZW44i3sAuSXNQ
OsTmgAnjOIJjWDkm1OpZYbuNiqJDKawuuEU9cgrRPIJ014eWfpNPKwCnnyaA
LhVq9p1eC/w6lZEzHZ3SMrfU+aFavY8+Fkmjf24nKNPPATRW8L+KdwypnI62
CLy+RLO+JqbTdy47XAMwAIvj2wLTs1uJp0hm84rfNH9D9NCYHvelmHcvnD5z
Qf44ZsiJ31mDxfqpBeaFwPyIoUNBDE1LECXeXnaWVPDsuNCEuzVUYZdZ1AI2
41LKSrhOER8sX2wgCuJ9hpw65JXVBKZM+NuYdBbSrVpEDkvVjT89orTIq8gN
tlqocic5mN2mPvSEA6jZKEhKepDsueClT/20FN8MDcl2Q0QhrErwFcQzQqMS
yCtUVouawqBCnw4s991oH9OS6fdkbArhXfMQ7rOk2BYX1B18Om/YbDMZ2TNt
t/eZMWn+nuedyA8qM0V3wuhFRWWRTqJk1OdjXpAyjdW9rgv/npD6xfU5J8as
icggTVkxBtdnkPf4H3PKAikRv7l/FxDK+0YNlNkHuu72bxy/vknru7e2K+1N
Mz9fv9J3gRnCuCnOto6lxEeRWMUArTKrKiVbSreadovWh62iO2HKP64q2sBC
yhmPmayRVlqJ347URjDyxr04xR8BIGpyB7bmiY4EGaXWoPRpk9iIDQsRkYWF
EW/IkMSd1EhvtQEjXbGKyYIINPbI0oMj3fdb4Qr0UvkjPEPpSGlZTzeLbMOz
/N7s8vdEL8mbtBHxoaNPtmCCs2jzKlnoaghjN+3orFQKH8J+VF50QjVxk42Z
yRjUfaBXbxtK8FnudHyro3mJ/LciK3NyKbuVJdgqN8b9V7xfetx6dFLZyY26
vvc03nHmWCFbrSesqYEqsqKgvHzBJvV8wK2b0WZVmik9rperHW9C0VOBBB0e
+Ap7UHbhr36JXkRC0mZAE2lD6CVipGwklVexDJE7GNzrnatGNdkmOv/CiW7Y
o8kVn2AYfjbriPrOQqXEf6B9qdEIYYxOThgBRKY+o4eUsqVOpwXc9P57vtNH
CUiqAb+JmjodGQtPKlpUhZouDWK8D8bs+MVAhoiuDFsEbz9dnhyQeYEV3Eg2
9LOD4cYjSqvGcsMBEx0q5muJl5BigN6VLeXtI4rhLw9DjV/b6v8Rt/+qZml4
h86emH+iaCxEwjt6X18u/nhENO588D+XKHpQBEbKOgKwY7LftmLe1iozMRC1
1dLUikAuw82l+nULb7lfjrGrHrdi6kvuSwIWqN1pjUwoLIXgE5PR990P2V9v
jQzqLLMMKYyD4CILSinATEKRDN9ah5WAOWWiRI4epX1UFvvSGlWIHt/PTr2z
NW5iwQduKSfkEGr0qDnJor+PbBsp08qG36NsASCebV/RA1EWZR0o5snRDSwj
PcHKGE4+NlHZ7ZrUE1Sdxim+UQB3tphj4L1vpPAx+rICHEoMDS8fMbQI4lfS
iuG0ssujDRbTjD91eMv7/8w+OE/8Hhikox6lKWVCnwOM+JWzxTgPK8DsE0jJ
wxbF3gdRf49d4cuUUxzkoOj85XswhPI9GIKfMBkMlKRmmhG4ODPCacbsMmVE
8FoRnpV8duhwc2jIbUq7sOxuIezxo8MgsWae0wsJyFsB1Rar8rcN49oZhCol
etaitp2cZXGTPJR2GwjIKpA7cHdQhO1BeU2/CWMOb9b6GGdCSyq4XE+qK9Sb
J/0IJwZuzSesjFCqpn0wYNFIEpWljaYSSGhSdls6ex0k2jKYG6M109v8kWwT
vnBDiimZeCSOux7YhOPs4gfPBRVv8r6ibZ+DIzcgLnabhPl1JuAfGw9l1Q66
0MMS8078+Xk8Rtf+P0/G0nD0AkdRtOE2jcn/iT08WiBjUQkXGZdY/qO6ouet
f8YJjrRE7SuDCuNjiiaefFs5/9yIfAKSwCwSXC+roxNpbX8/x58FOwKJ350j
JGHz46vAyqIOHCBSX37x3QLnj596pBnZk0Y9WKWO7GyD65j8CgYv+RmbNYe2
y4btHEYzTO4YzQkMEvz76bBYM4eQgQGWCSnuTIA04uSn/qhzOa6IlQB+fj6V
NiLYVV4oqyNueos5MHnSgh7UxlkHPToYnesJJHGMRqGDZ0GDZZ3yDUZHYMf4
1wiWWziqe/Qpmwo+X5K/m8xkTMutyNCiAwyEWthHDAuCd4eXdWzrLkaC5Iig
CZPQHMWO0b5Fegt2AOqLmUeyzYtAmcJLkRCumUoHBQkt9ymnrKCYdThrK3db
NUfoDyLsfwbdlJVH/AyYBK36xOiSalaZHiGHF0sAIHWAPBv2wdYAK94IVs5B
JhY9ZT6B5GToDUGbFRd7L8M9AZXBydr3nvNwN0DyN1x48RSYPdjrjqTTIzl4
Fx2PgXlzrzAlXcHW7HriNj3nxLP/XyCCcxjJHGf+aYa0icG0xoZlVePQ0qLq
86fUu+An1UWR+p2v7VQlH4zZQZUIPR1ve0BR0JA6xgasw1aK2gM5E0/AcDSg
xeyBWBdde4CDHOrxlhG7KSdF43xm9T7Fooc3z8wpapx/tjbk9GOA+I7s8nD6
FSr/qZcMhBiWX2rnqgiDRwtr1QdnqDKNh2aPGHMDCI0N4HgdRvxSKH/6RM6c
BuIpzOlaV+pbz344dODMnXLY64T3SiGhyDSSH990YkrlYIhY/nFyKWmRmfYh
okxPaJtohapY7L2etln1zgmAeg9yGTrb2K86rZXn36y8LkfbCdwDBCvQhhWb
1DJYd21hSHMjEbsnnVJrTvGGpOzksYrdRgLgeXsgI8jHoTZq/0DS6KSx/hgq
Xq3X5qIoH2hK7IIg9Y00XpiD5tZkWKJ0Mu1wquKdEmLzi8k/1WkPobDLQ4iQ
rxY+c3ktcN4jAXyvxHiTNuZ3byxtT80hbYtvaEiU9kPaHzeaD9JqKpwKtkmD
y5uOHqsnI9DPsnaZCCngdHGRAH2r1PnCbdPFaIKqyRx7yuAJ+qNmsmRdSxCX
dD3l3lP4n9AAxE1B6EZGxB5a+8sTnAqPFWv1Oqjo0ehfyzdlWlDVDibjW4N7
qZEW4zx5o4UkrVfp4DShFnHXgr+OQbOqbqP6eFwFmxVexLITgNQ6rma/6ZJr
bTegSHI2mx6Kh26A4kTvcJGi+tyILnB56CtM5zZsezN9nvQ63ii2xU/kv2x3
0GM3T579G5UBEpaE5iCh8Dvfle0RjYiYAIUNrDg8AvOuGcXga1c56z8Js0pI
DHZWLiPdYCGxvie6k1lMN3aTrTb3n31X/Q2bly5oREiOEwR6Mj2Wai/C1MTO
EIQpHh6QWuKXdZc9SSIUIuEjJ0m7cujnrxaHZSmgOYqlb3DlQs20NRqRCRGG
R7k223+AtK6j7fTj6473LWUvJ/fUxB672ExGqIQNyEgJOr9iW0ilR0lxXoRI
Gl4LEBuYyH99DBmJNGhIhIEWJQatTr1I1LSbLonkg7ep59EZfslBKdvyXyFw
Xsl8TwJRKQjZVPeUFOf9/00ODa5WOn2FyX5CCT/XDDAdoNCBtNPtx1fgdJCD
JJksXoAUollwlSwcnvS2MhtOkm8Ludlq1aQ2ZXNV07R3kj7ip+eiAuWyQ8z+
v7pPKh+bYp5ov+AREz1ZhvmaZloadfvtTUMW8mJLbyH6+BElROn9xZFxRZvh
CRFN+HRJHk23EQov60N8tRXojwaHnDOcEcyMecPNItcEQPFm8AIkgiJrIi+e
InHHK5sDtLncVcKukL7GqqCmuwbJKGnhBFC7TnrAzKfrod9rSGgy/DuEdT40
J4uMdP12Sw1MIdiRxVZUGoMq8MUCr96hcnFQudmyPHaKSx/wMPgx2YNzqXgr
2Dp56DvGHMaz0sWs+yTC6Gs8ULtSLoDFhNIi2n37mLiIUZW1z6IC1cHabXgE
su3ZifYW+ce6Vw8HssqEyE1xuWZtZ7vOdTNOMOAIpUXMY9RequmNGU9xggDr
VUQmrJPZBe/wOx/7c3uRndLv0KOW7/TBjSnKnMrR0rmu8GDvnKjhd2CZE0Qh
rk1oH1IrifEq7YcnR4119IP6JtphfZX3OVV1yzByMKRm3fAfWiuc4fv1dWLQ
MXlPdzloz8yxaf2/lbB6DwRERU9APFkYMLj77MaqEe+ahvNR1pkVjhNAhhMI
2wC1XfXVlf0iO6eBzkYSqCLE0K6lJ9+RPCFUMp7z+sxkEmVdnil6EFb7p33S
4FEMWzT1ZfuRztIubnqTY6vJ6a7Zx/aZoOJTCv/y8XrnB+1zxoPPLH6fKvu1
yupOEsuid6+I0BEMI6Ec9D8u7aJgL3r4vs3lcHfyUtNkf72P5dEDBJEcy5Ki
lBeEM6bdrPCQtuibMRzDMhS73UbSVNANoJCpZ2HnW5woJu2Eq+M7BIE+g191
FaAHd6igVxRlq/HsB9JBXPojhzThN6aWdGDl0g/2upTaBciGUWAgEBWrPHI1
mISKF9uhtyl5oR8xB0SyUposxEiOTTLsy4ePbI5CqDTtvjjXu5pc4GRI2zKQ
uhj4uMWPPTMbrMtnyPNKqSThnRwg4/OJEa0dRoWCk9uAN5t+OAxLVZyq0C36
O+Z9JojHJH7OurTm6XBpt0ska12zcjFJLbFflt4pLFB9vr9F7q5NI4J1YBeo
9WhXYap7ks5EOgBbMzPlkY44cIwL24eRvX8a9kPAqiQZtd1gpJ3z71+KSnIY
P3EhTRnMcLSzmpowVIYTFqxAAj0mW6Aup9by0jRbuFzEnma6RqmF9Ozng0VC
axd3ukwolIFpJAkUPnZ9b1nwqVniDiITDwthJCGualji7LVwn8xgkMNWEmnb
GzcUSplMVyDe/vA3OXin/4ydocq3wVbJpP995KWNXd5Eh6FFXJSOFuT0XzTE
WnfQLjU8civyorwqKRwl677yL9ViRdW6e0SRtXVBGRxdmj8BdnCRwjBoVqg3
KDW6XFb9+/gyP5NfbfOBgTuLmjaDHs/SFklq/vB9eMcaZD/eI0j+weqKEtu0
P/V9kPNQwxeM4yI50kYwKihNaX6DxqRKabh+Edz647WF61g/j6Dux8vQRgcW
6MF+NZTdgxmYjr7nJIN6PYDiC7UTzCPE2Q9uSMCh6pIiHJ/UL52mNE7QsLmT
Bwqu7aUITMDmhOv/sQBGPJrIr6MK9PF0YUWSEZiR9QRrfR1oCa2g0k+bAYZL
h4vZXHcyBQBZVQkxqDh7lUa0UXYZiH1zyNk+Ln+BKzg9sAq6HYpEj0eQVO4k
DfmDMyHeGzqQjVxDfM8691toVZh1HEDqvWhCEYA8OOwWmF1osAqD+UAK8FA7
0z8lsKMGx08nYbHlJLhdXv9aAISCfxICjdTatwfTE25Xuz/IKqvfTXZsD0l+
9E0odS+546r2YzvqqiNbH9nSRkHF1M8uImDjdG4iB8MerrNeil718o3KE+/2
E2NW3/9ZsnoLGN1BIqZ3B3jB6wLamskgpVtCCH5fMqW+m3uMDfcrvvM6j8Rn
baHWvDptXrVbW+MnSDE+WAKRjAdcPWV8C5Em52nQQJ7G/kZWvPYUdGuarYMm
ivmrmdoGh6nFoJ2kV+ubo+5F1/GmZrKBc/0nLA5sI78YeySAnoAnn05n0XuA
YtXXBy2vxiPzBQshZgwyIAcm5Vn4jvvd65rmKkrrTZM9bIqJw+3r37zE5995
weSUAdYorLcDjVhOLEn76M/GnZ7+FasOPuYXB7fC7jOQub20gZkqbljut7sb
wrHhLVTdqoyWl32C25CgHQBVHY4ozi9IfdtdhxH8jSxs2KqoZQLJO0Y5gIeR
0XAqfGAPImPBKRlXmGjHeZKGrau2Rz4WWAvtDMdI+Oj71eXCrTq1/F+EUV9x
oX4cpowPNrll0S9kcNDmKmfAV9Z7xbfOkmZcMuK7siDRF5M0Km+RIo6TQKE5
/w/9YFz7uIOlUNHzBAXMO7Gqp2ezDZw5JDrzr+eZycpliNcwIWqTn3Ps6z0U
CBC3IjwCQnJk/hbeYvpS0V1ukxrnfqbmiQ8wvb9zViJUWmqRFgZFzNTWo1oE
bPr9ZgXS17HMeBxDe1BYpwySuyqHcGCdapVa/8C2h+1LCcQCydXoFbyIoU0m
jHY6YXDZybUgz7Q/sDUcPN/9rfA/Xt6Tu4PgqctQEGDdCdtX6x1uNtfRGGqI
X5F+Jy/rObwLP/0nvsWSvmdSafSO6cJUTdxQyFfB+O3Jdl3DLhneDn29rN6O
Jh/0ugO1QLOwaZXHNVApSecw7UaNJTe41Ev/43bGjwILXRXBUd3uCuiL3yxA
yNbna+UCHaSHZhm6m2Ug1DW0r8ul3FuBohnqUwP3v0TU68zWo6SbP6HgE9xf
2OcR2BPWwS57TV+isJJ+HspgF8ZYgATZvqQ0tP/O0AH+noynSNk0d5Eege+n
HLvoJ9yHegU19rBXQpdB429vu5HUOr8F/FwOVd0uarKJTvsimMmFeuxLT57F
/3SxUVZBaIAgmh58Tj/TDHAjtukb27tXSSOH8itwRr4G9XbXj5yMbbloGb/9
u0QKQnRvBVAeLVfYC+UF1luPjeKUhGoTpmiRm/iKM5Zh7nNDo90+EmHf8UQK
8A7UX2jTtJze4Ix7e3eaEDUV60lMVl5qDfiS1b45/rNg6dX8kNVVO/Mhqxyi
h10Iz4YIRYdwI55inAXsLfmwD/Z6rKjxN0OeZOMaEBIIjwNPtR/TfIa2ZGh8
0gNph/lb+ky8Rx6IWZS8rICuBaskC+mTYiQgRqCCM6Ge43sSQiRQ7gwLSZcY
/figTBK/IbMlvy3nzbZBl5wa4LYHuM5+nMO3S/Lz+NoeoX4frSJ6gcxanMrq
9qgqENL+JQMlr+bM7yI9PbcysPIuHJ9jd0JS1aqTEvclOY9Xsmei9EI68vKP
Y1j1QxFN2hBymKcqIuH0B5qf7Jnqo8dT6T/VuNlDl4zMdAtzDyk6YUGWv11L
LUkYqRB7/Rm2Ay5Hxb/PXBUK6yLIS5UtrAyXjyWX6x/VeWdt+ZQNowBFyuB/
F2KDhtMmhG9TQnjJyzuBAParFV2ePmbqK30bkiWfjvzS0TNEsdJWYUyB72l0
2WDNf/5Hc0bDw7iibHgMqJ2hzMNh0GGf95ZP/0JqBo5VQaCSYOZQMtXdawft
F7VO5Ao+ifPUOEN/8HHE/0XpKdbv6HCGd5yMDF7pFa5zL53OuFF/H+sSHPzA
Lhe1s6PI0DnQ5cYRVR+NZbRlHq9cY/1ntASXKzYx6h336h/2n71hSCQBf8UA
jYUPZY/45L8RX/a7wYEYwpiqLHg9hxLchYWklSbY8GJ19jGkKcy6B0uNXVom
8k8ecU+kcuKoM6xXn/rcbfV9FbK2ikxnuxqRsAn3yXKuXvbj02X51H5OxluJ
wVmb8C2cpY0Q66rPyxtUeHXQ5Fuy5HB5hBL4Cwd8HcAei23Np3La/3Xy4lY0
LUn92ZYCbQlm5z112VlbGaY4E3HOnRwl0+DhFMPRyMoozOwxIJk77OO3piYS
8n3oLR0hbSTs+ApJFTL9wUVJPSuHGrB0R8fIqxV14QrKa9gc+Pnk2eiOd09S
+PO3huU4T8QWt4T5uYUl6Wd3TOQAIsaoE7cveQofbrUCxoWAKUZz9RuCoObr
iSnbl5bhbfsSJ7RV9RTrC5F/6JtpN/vtvoRkmzy8Abeoj9Pqh/IetMN6V7du
jPUJjXKX6p52f/edX0KLbtTH+Zi9jAIUPQQNDBcJcTPCaBtL3vEMMXa8p6im
5HcLHZsMtYAHMq1QSL9sfecjLMQKtWjzn5TdxdjLjLGVsujIR9BPvamJ4C4R
iYNGKBIh9yA+6KiulC9JTggzdZX/dethNyyWwCncIn0xMlRKm5PODY48+6sX
ZGfyESd6MIT+gIRVwzR4LqNMrPQhmyWijMoltqBGZtejLnq9gMSOb60RRLj1
C4wK5KnN4eNgZDOwaOl9uQ0eamGNR41ju+xTvWL84Oi+emxXsG5XjZ5UgABi
bQUbyCupiq0goBbEOYWJwJstHghvmSV8/GN7EN345w5IvNkcmE0da4Si6hS5
+984nkYofjQUnVCqtMCGTXOaN+NZGS/2fes7a5mVx30GODj5bd2mnlToNekU
DOIlL7FmJTmene9E5ocY6NoNkFpaAU0hCGHfjy/G0SaGbv/9JxAXKaOMJL0E
AIkSrLIIp21qZGqk3W/l5WgmSdGcM07PutoT7y48Zh7JycJKWQpRlJrEtn9+
zT5xDIg2eBXuC+xv6gAUQbSefXQh2ZVOJqMCPDMg7KE2rqsKAGPJvz7W4tdY
qpc4+VvGv2wiuxz4Bz4N0gDjbtjDd67+ti2RGvacWU0ua18NanwwTsn+kYux
6v6BMRJ4j4nLyBn0t2suv//vHRbhbO/xxXxsK0K0zTXREifRMlkKhC1hwqSn
5sHium+VqNzZoxA86tz7F6+ocYyEat0LYNwqGA5QK4vSnzC6TcxLKZ/A7hWR
7h4rWNfPwVwdo6EW8QbJCs8IEn3LZ/yquABiLIMku79mPASkcp8ecHNBkabp
zstDZtcwWjD1ufR1xr41yDtjidc+SZJYxv6t7HNPnib9NyirGdZPeLfKTNmP
jkCsW1ya6rknF3TyC04vD6mTGt1J2s9oysZrMEOezoH6ZP7MICIP+8DVBl6W
zzvco8M1Sd2DBT/FmhYGx8z8YUd+ivbXZRXD89yhuUVFD91Xfrs43+l1lvmr
SdLy/d6/c3qSScxpg/1QTuRAHk2jQmpllA2qWfpCcVJUUrzfduvL5gJXvODB
Y69PCrqwPP4s42wGUV5tXkpXi6tQL4hV+gKxcOwgymLSfcZP7MQ5yHHvuzDM
I4jk/BPiDfQRZ19+qBZ11S4rChun5XHEdBYwSuvxCnwY0me/WT28rqg2Mg9/
7zGMfpIq5QF5n5/dTTMLDpWMKnQrZ6KwfpFR58NXEo5CtuwtoJnBtnzdYT8J
uy2FXnG5oWVyFYf/VfwBAD232OyQ5lQgWur5TojPORWTRSyl2hqu4Tgukbtn
nGj5C5K6QFy4QjQX65ETSlh0vcSVSlZMIlXtyDXmdNv3Hc/wWvurWWKENw1Z
M7C3cr4onFlWqekzwfBwCBJGQFQgwjgw+PKyQfoexAQYQEzEtntPHiutnKjY
ytjneBADsMyq5l8Yxt7WoIzvfDkS/4IqxT7cL4siWlCcWBPB8zx7+LjUXFgn
BtAVaREGZgslhHNJTxgB3zGwQ1y5hen/8RhksBWYxo7eA2XejUriWYmFv6Tm
0dmQopqQqeynZW5CC9b0GjayNdcHPEobJzGJq5XEo1Tfa307mqUj26lj+Nxc
ofvQg5HksfwpvZiWykNaqAjS4W55stsVqkehw3jX3VJhWomQsoVveapzdt9o
++7/J2aL9lzSjS15x+BhDWyQxghyiYx2AFXL9Ub2J+uS9uyi/xqswNHajXfh
XO43H0DZ4QvDkv2fddkFsW06EOXef8QX9NypF5c3/O3rzUJJ+Icd0bk1dRDd
lvaM0jsjO2fBhFYnMlEf6Kc9HUyMbd6RxnFgRLH4osmp9NrGuyHAa3Vsj34r
UsXTgBco4IYh/lq2J+r0BExClxtgwVYaEoLLd2suMSTh2NbzeOC39YXkZFYa
GFWlNYzeOdD5USMF+b1Iya7gthRfK6SktyYr4Gn9ruyWqqfHkgnx0edlCsl7
rcxdHK13UZdnj94tBThCIeIn3vM9KeO69/fqfIZk1OoxcQr9jJzzevFPpgWP
ST9ixNnwxxTP7DOFcqaIh/qwL2JTrfH59oclfesvf+zC9PN9cNQR9zGMiDY8
2gqBAXB0fuQszqhXszu5tbOH11b5NVRQ6Of+PIupjV02D8WmiEJiU2e6KUpB
vi7fpfDcaD5mXEGMHpGXTCWIuPnZp8U2ZFLSNSVjCFJeTvsLQEJNQiLWi2cn
zPo6OLrwC5Km1jp6IOIJblnu5mA7YPzSRG72a2HajExnrAnHw8czD+ApXz0h
XqNbRq/ShRWsYv8uWsCUfgJ8la0ciJvywQyvih/UY9l+Khl9uz19mkR1jFw1
FY8zKYdA3w3Kz9t/MQV6BhQVXk8UyW/Nq6+pQ5CmsHXOen0HOqMgs5fzPxGu
O6cHOlwCqE7f3WdeLUvmb5F5IUL4MoQHCLh6U4OZ132x/ujpGaK/VXU+3RXj
MaG2TXzo/4pme+zMF6n72g/Xw0SVbZ1X2LhlxvhmZblwAYce3qup/Cfri1Nh
U6Ru+3IiowuSGJOUTAogNeTyHtlAPrQzyuUMDZB7l+rDzSFXFiF8OYl4Xdes
EOU63Z1jXpHJXp6+kJ3ANfCX135lyC+0N3cIOxmmRRyeaRSxq6zTQRVT6HRF
Rdq2B7by2CgodIgA8bTHWgFxnbOMDV41lAQcQHxmNmdUv4pZyu6m/+7VJ4ce
yAM3Tfflfljn6+r0aI3ADFa6DVnWOjEIKoMYHyiyKfhuHcrHiXdvfmOS3Jf6
+xFfmIjedOgBgbeRnDdSGb0RIwMIfC5U5wpnnUKcFzPf5vil0C5cm5CWCcEO
3pzZw7iws6ENnE0pMAEqvT8AJgczVZOKIfPDNZuK1nOgJv0Z42SafYwpFIR/
YSdNGgJ1wJxW0pCUohMZWtjGiZxq9d4FnGJz1zYZgvDUq+OstznAeen4k/3n
UXVEaZd9o4w6X/NE+4Gv0Ptj+vwt6uWaceKYf6vB5lL/5m71KLKQ0X581I4x
q/EkhLRH3yK7uvGvrR2B84J7SzsLlkbLzYZrXqWMaC1FggHrlIBEooBxzHTZ
+aVcERs4weJ0hOqdE8OW1BjWRKXAr7d/Hkm7RmUePdcdDy1Qwtze5jr6YR+B
leBDRKsv7sGHHnTqUIzM+i1iHsvmHIOS+65VZ1Dl75yNULuhT6EyuhcBcscD
ZEBDaba0pK/KUFNPjzy+TmpJtSgfLTmHD/WETl62p/jF7aEqWBkkAhTOklz2
fr3bnTTRuUjyDcAVlaa20MJ0Vt4kHCKxMW40o1wBSpdxoEdeKxxrquaQzO+y
1nLCCaXs9v7iGC0CkZy9gRYJruiDaSP3yD9UT0d1YJ9QUT/6P6jbg7bJhusk
vihotateFrNuvnriC2sw+PtRAzoORiTA7VREyGVTKo3eTq42gzxtGgyrkXKE
ewSNo+IAwdSU3JDc1g7pAwIhQT4C4X/iZkn8s2hBcD457HBdc40veexJVr/B
YRgTVnhqaorH9RW9MwsxCA3+fN2Hcin1A6pl24tPVbP0ka/MtRNvhy4lL4BS
0L43xJq1v5kUwEk3e3Mn+Yz17E6Hu9VI294pp5roLVKJwYuz/YZw3kdRzDc4
ZmcJX9JUmNcEmhZahRVHm5kf9gWXIudiV4E0TfdPPXRzuFL6TESLt8hi5ayI
funut+vdS9oxDEDU90lJctyph+ncnerXGfXf9r8kilkoB4RJDFdbpIChf5f0
sYShVJVR4McsXAc6sMsRmCNzSLA1dslmAtDG6wD6cJlQNSqDnup6NPrbQg3m
0hhmnAG6jQWU8IxHDOyuRXQ8iFxivm+vv+YMwwhb9w6iCv/rjMf3UmPjF5hk
t2wSwcaS4YnBMBNB8WJ/47yAO8Sp3Q2iTwDrfMrhp5DP0If7eXZFU4t0fw+s
pT1o/D4p3C9RfJsvuZ3g2Ot0390tsEETx7IxL0mqh29u+C4Whijv9t7Eb03+
609WJw5o7OWma/YHBkJ7Tg0W5KnO2rfUUX7DlJe49OVCxsNMoOSexLEaZCA9
9KZf7ttdeRntE3imekq+BF78OtWXYWuzhiGvsdGobQEcn6lTkCssdfsKYp2O
ZlzMI5kdyOLkO1KO8+GSW2WBwzSHsdWqZHPpzwtOprLwF3gLbZx5q95fP0OL
SSDvV4IDO3J+2K05KSCsz4Z72dVwTU4e82ThqgVI/cqDiAPMyDTXGILB2P/j
fJKiefjU2lZ7cE1cra41BQS09wrHP8PBtBtnC3EqWiLaPxyc2ykjYeiBZYx4
Eoi/w71keDOAPSyxUvaU7jndRfQNmrlpP4MgS616j6ZKz6UOMNU5jq/vIJgM
fcIv2U5js5rg3rCf3I7AS18ft6baIO28MxiRS+UjwlSrdaJwXiunw8xKjtAa
ZuUY0TBkgcQjZ8MKm6OGEGclE2tF4Azp2+FU4gj845l0zGlawdImC7Vw195a
jdCqfEyHF0SPaqDzyBHzSB4bn/43P6y2+kEur3iXjIelr8VhKlfx/OYQw0D9
xYdpA1Ta5nbHBMFR4P6sGGAZASCwQf3w6BeYDYX8UU/K+W5Vl3wIz1LTrqee
h1/Y3FEz9ROsIPUIyYaWI6chxXuQS3OGY3ZEH6R1LbmfIdrPavjZSFUV/KQN
Hp+f3A5XJZRT3WMfE6Sck3K8lIYfzivWBkTpj//ewf80yOwSIxnuU9ZWII/9
dRWK+yvLmtZBdf1U/Y+DjP7slldu94sQg+F1gB6gOKjyZPABAowOtLmSeegb
QrDHPDxmsX+IhS+q5UCg99d1ZVnIDiXX2A5/LoV5r43PC68sF9UkHWZFAZW3
JVolzDZvVo9thVJBC+U1ZEfSy43TbSYvjH0G2YzupRvmMsznLzCZjwX8Hbsg
DEyT7cHtLENlA97FEiiKPRJm4fm7pbOV6hdhJQ2et6DAPf+uA9Sqxr6CO0b3
RHxAqxBgrXKTiGWDbBkiZjpU0/1jBoXrSSck+YccL+2yy4HvhzoLuXS+MEt0
0UAxaTzaBBm7+WntXTachPDeaXoAnx4CPC6eqYNOkkwdXnwny2trh9bi89cE
e0BMJmRjJYn18J+ZTPWbjEGSRuWTijPi1c7Q6kxm2vjVBoWGmij+Zes3hW0f
rLNqM/015EjH7vQXcryW3HPr93bwSCoLjxqpcFQtDgO0B+7rnfWMlLRvdVIl
bEXMxyNugE9YKwrbJg1scNgYiOgF9xCij315rgKko1RmpCUxnNgACgc5bM/f
3C2aCAgeXNH9TMJS9WPrTj6c2R75rnNR5ZltgIesuMsHreXz0mtmxogzpqTk
TFzJg2thwM02QgORtAHORQwRq0IYpGsDlKbgJusLaohXMRgVBdInMQ5EyN2l
TqVPmgUoSoO4Tc7peNJRvQ1r+XvSuu2dzf0SSmNbmM+VM71gmdNTyXc19b+j
/zpRXZHBbqxgd5wM/bp6pp6rFpUddTyEFQ2bB52b5AsEE2g/ZYmn3IYaYX4w
6RrMTWjOYzHq8Gxk9AiAMeZup5WaOe7lF2uOCP1RTF0hkusX+wpCPvy/LdaZ
/s7EFP0LMnCap8gD2bdTbFruZUtrZ6uBCSD253KS5AnY7BORk9HYndguMnTQ
UIkmKSPKJb1NSigJsx0AsUUNKtlhxbsAxQMiaSd4Nh+p8Kd0+xlyGSVIBxJf
ZYOVVIeX95J0YfLzDTPJJeQedCwHhQtpo4DlTQDYAy4Est+d11pDrt4FUM1k
G8o5OrU5R4u0Iu0FqSOzzsKQDO6uqE80fj3KP1TL6etcGNSG19nPj/S4wi+R
OTG/No7xoRaMZTOx6YubCH4ben7cxVouVDE0vzKot31V5ig2r8mlr91tfMxX
AIJhRgSxRdOncG6Mxhdz6Qp5DouJ5v8oefmj0Y8Co0RZh4fO6aK/Gr7+BhUU
2PUtQKJEomT9tHcy0aw2T7UCwjdIFfMwZQtT7r1Kgc5fERqMpRj4JmsK+ZJz
MoKm79Utly4cBSedYJ//udDLipgjEIdfCJKyHBlxnpVlCLSAVIjsAqnJ4DFO
uh03PkSSRW2HbRYJcOiUpwSltQC+4J0vbhYfyBvlxcFassHH5GAGWMlgNl55
0vTxPnQ2w/gB5nRx2AcYcUC1H5GCPpMfgz4SGHKkXDW8l/4/Vj5SmCchg045
0q4pxldYk+LqcNoZDmafkjlRORJDg4txO16t1jZEOqRS8t+vHxmYEtU/7nke
/Nyhqs13MSuizAj6o1VgN1pfVaTFV1Qn63OTFgY6wklCuUFLGOPKvXCopINp
pMacYzoo8cTuCWUYchJpvIWJbZzwo+NKS6Qc2MoMIdmgdcxRHrG/gmZedMUo
kNbS1ebJORwIBhY1Ir8tNiwRF2dagi3w8LAdqsmqS91JGUgkImxWMAlH4HRQ
7QIc2qXGr82LixPTbNthyCAvMLqfCIb8tn+HRmDlW0ZJ51jbIp2CXR91JjxK
YgWQHLz4bmdt88uG/KpWKhlsb5siJEZIatbOsA9d/ShzgcTgJc+r5Gk3hgg4
D4hz6DwuPEXc/iKAyYU707klKovPcwaJD4Ep1zMvLCQUrdMyyfcSWrz+kvN0
wuqUWGA5HdVETtM9fLDCKG6PUHWSI6YXoLQT64pBp0bOrU16VfUOuVk/n8Sb
2QxbK2g5a8ugrfBLH1vQ1ErERkuLnuXa3N71BhpWeZlyYPbkEULwllBXQFcv
qYkwz3RDe12YvdIqTJPe2SNVfaG18cbGGHUhpGOIHmgKC4WQ+VoFncPj1yVB
X+lLG4whfPF9wMtCEV4c9H1EZlyZLOGmi71Fl2C9GwBNY+JLKiowwFOIlMsn
rzYshZqscfXgMjDeHY/EgViVukSftvKqGPZ2kyGdXJa64pF2xInT5bkNSp1s
WTUAezbnisFDtZw9MadYiGoR69uvx8u5e73j6EoNCIXfrtyTx3IzGacEjwpp
Hh1fac+oeIuZAXH20vERKAEZEL1xgJkr1/fg0OED0z8cVxz4BfLg1pm+1dTJ
8bWUmhNLevgwOB4y3r+VXIOV6TldZC6iJSNOY1iFcHL5y694YhZ1aBpajUP9
xQ8XUli146hhcsfybRpyJnCk+tWhsUU/ngmHvW+2k6Nri5w32aBI28nqTixD
G7Q0raZaocI2p2zo+Pw3uj5YH0m95KRsFsBQblsciRKsb9MZPPqTcpNy3dN6
2rDit+li7nqcUhTY0v3C86QPRHlhCN+mu1thQyjFCwBJifFGt99OIfoS1wKM
iKXIAu8LmyMQHTJE0BMbwZ+bY0bAaJ1YfWatHUQd4tL9Z/iC8irV2R99YrUD
hzwZT9WV0vaul9Wj78pWmzfPA9BbbStyJklfUCY5C9WI0nYkypnAbds1DLNr
EBn4AlTm2QLxzVmU2CzHJqltnzS/66otzaTos78uhPKVcmz8sTJciBAR9/3D
GBKUHPzPaFlV8YNM7Tq03+5bbCbnPMXNaC/9wh0eCNo+IAUUNfnk90sRSVlQ
Uj+tCJahU0sm3nm3WJLt5WWGKNiV6UhtjGf9w35QzNPG4NYsmkvCbgF15X9+
0TOFdgN4YUfznJh7Vi8mCOM/g77U0toGT1i337nQEuF/uKK51lNdcz1IDApf
0cc6aiXBvIh3xg0pU+k+F8wF2z5QYz+UCvRbfP9HRzEPyNK6NPNSov7pNg5f
aLyE7fXh3FJE4P7uA9FKIr0/TnPDW9/VRidw2H0SLX9dUajCXy4nM2ALU16I
xC3U/fREu4ta3XtqAbpjFVsf/jMwKa+ANNPKzRVZ2fcs7SW51SqCTZZ7OLHX
tDGmeZUvHHyOwZyVjEmbewUsrwJqnyase20giXBIByayh5LJn/GgHAyHA9+L
q/6el04OZFYMBsr8tDVqenmNvuybokRfCS/UyUb0kAD4ZldYxoLpVocYujZ7
n9FqMmV73PQOnJm+sSk6ElHFUsEZnHJ2Q6yXdvoMit1HHzqwjszqhFUkDtC2
WVGbGLZAAJZlVZjaVfbFVMdCndZmYFO76tRZkbCv6bG/XRILYinmic9DR5Qc
2gqMYcv+tgEpoMjaLdDK7lwRlVadxHZnEgkZPVtVgisZo2ric5ipJiNX9vip
7Ez5q74hJ+pjlBqQVBDP6MkmRjY3weHk7hwy9vFAPGrHsjU8uQe4/HLwZpln
2MOmaqcjEj6xyXQbLJFkoxDXFd3KVVo3oYXEM7HOkfPAoSxrbSnPycqgxZdY
T4P4raUR6nGFdTi9AJilTbb2k5T41cwaxTa24kvpI38Jmz+vs8T8ef+ocBT0
t/Hxvk4RE1yWJ5wyUT+aOaqKsSGV5C9SXaXrXhP2xxPLyBUTPDO+UH54DOVy
dp22ZI0ox/FhiteEe/w+zjWT1kHC3cAQXC22NelbRE+kD+hF3JRrMD6Vye3n
Yws2JLKsfZYUbRMAOFmmOgru/GNB8jaZGdodOcgU4XhrIQmlFUUoOx5bLgTk
1pW0QtKCKpYpgMt00j1RCM/YhzlvF5C2qkLAYmkJ79gist3FRqdgY7yZebtt
nvYT8YH3B9Q9+6SibKzZlu/uUm78XP/6txrH5mJB9kOa9mQkkdPuIWDddooW
Ay8WhpkSrOX7GgWpvlhCifsQJQyJrYYEX09TVJ3/T0Ro2HkfmfBdlwIKmpyH
WR3yR3TyFAoTsCz16kZUeSr67BfLPgxdKjDTMWC1hljwjwnDRmdoatEs2hpz
NZ0+mAzDg2s1FzPqW3hrNZ/UZnEg6ilOxgxErH+F/xueUNzmXNl+q5iDvVqy
xh8fsuDFBZ5ENNVEAALRdmW0aZiTMCJTxjlRUUHE+MraV1APnIR7sLJB6JH2
mxZ0gOMMPOfBJD/sDQYJ0PdENyhX4EuNMa6MGr87nGJCA8xkebzYekjA/P5u
95Qo6W98q5aRvC3W+0Vgt5Le6VLjk/Vt03KKH6uEqix1COE3LVttxVSujzQg
wlF9MXsvbKHx3mdgYQdOZvVhPpJ04mrACvr4mivnbDZi1T9CsnXwWyrLl4k/
seQooza1Co9diP7SCAFYIJ1HS+tDzoiucng32pvEO7+mm7ei0HBqjeKyoCFc
pASjz+JgJ09RQBbwO38TTQYIwhGQbougBaOmgdtzWfyJOf3wpKQOfPAL/xRH
MEwKLgwmDHygZwryqdnMxo6FFcrqSWczurm202NiVvhXemgLGjm3iOhdmHBh
WIIBXLVFQ4fHZzC4uCREpsZVhk70rMGwDl7Y4uPT6SIqObmsZKy6KACDWn6d
pSBum3uIA2WLZvfZJRPUChxDY+zwdrfQZRxdUcYEG+yNlre67cBGfUPdFDP8
zuEGruiEMlTjquAyf5zg0JlqSKquy0ocDze92bsU+wjlahqKQEW77Py9dGBE
KzMvdiOupyeCd8dBa6TQLcl+L1Od8lTb6AkCNzbPOedHZn3YA/ZFhioZhg0m
kuZrwrldsFsJ5PVaXKr9891Y+dWBTD7sYzkx3NyMEjg8YyJpG2/9s01vs5Fz
043mQjxQokQjTnS83YUkm7GHOdxJ4ibUpZBHDGZMJVRebxL7mnuf9Ac18DUx
83quJ7PqPVrWdDkvdoELYbHdghz5X8Oj6wiaxqsCVvCAIR3NLOiygGeQpYkD
EkB4Ac50Ty8JJzD24Boh6Nffu0lRVIpBLRPhsBicmvJdokCWQMa9r8k2XoY7
TrjX2jbpnQYMDuarMYl+x/gTzz7u2ODiKy8uSTqsHdFtTU/YxGXoW03ZNm2u
2HPBxK9XIBDgHxSEhOAJGSD0F/8psa/JIbqCgwrOm1VXuzyLZcWOrWCrGthe
XFUMQK+aUaCZorrP+n6VjSY+dxKWJEKbZLDXu6Qd8925iD9dHkQ7W0gc6HxI
70Biw0DkgnGoP+P45oRQRZJXNya7HKp7nf/C1YYOMd/1X8bdIeBerPp0yYcP
+FMzWegYUUIN3AClod9cOL9Hw/cZ9erC4pkam94xS6RY3k5AOtTTShzrgavI
G1V+v9iGHBwbrWB8vd2pRBVzamRh1p522xZZe/3uKZ9HfIhXdSoOiJ32exr9
Re1COPE016RHZ2B+LGniQILkVGeiYIRQi+OMM1VOobvCPYfA8ZiHCUjTmx33
Sky0OKcmvYbw/G0N9AmGKZc2sZxmWVibbeeZM5pVB6xA1vGiwSx29SOk/P4s
ig0NBGJhXJfOxH1msWeWmETvJY1gMeE0P8jghmDya4b1YqWxReNmGgC5Y/3/
JfHKWG0DH8wriWuC8IirKrFZrZubl/V6JcEGu6IKzLZcOh75RGQR4MFUOg0a
9321Q27F9YdPAxQI0hZZJj42wRTL/ceR7Yl4HhtHHVLIzLmID98+wCs8fW7F
TPkp1ETKnJl5EGe9odt90F23NQiRcUoE/BG5qo2FgZX5cyj6baNhA5a3F5oa
PEfwD2b9KKJxtxBmwy3zTKd16YdQfxI7+ZeiRYknzrcqTwmhvOtblEEjCK7g
u/foleqfkTty7riwKVJdbGJ9qmv4UfkqtnkmQLgbwO7Z46NkvXlbw3yfzN5C
Sfwh82azpwFIeszv0PoUbeVvGDs1Ol7Yt6IB6WDuzO5nlPutrF85f5lC3+y8
YCjL5PKZwGaCwFnz8imE8IaTw4RcGMKM7oh7KqwH5rndVJlUNnloCq+zmgpl
n0SuK3JARD8Rxs0BLlguN1rozTo2UiU+hcapuM7gfh5xqXQvP9F32zg0VYU0
chShLT02pbrTfLENoaxtk9uZtJb+abg6FP5jj/jQ2HPTYKgt+kv8fDaZFTNT
Y5d39jaGh2sNLRE03tl+75kjP/2YRofwUEU+weih5Hf0vyW2S2n7oV6lRoAs
haJ3qzNtI4RyDJUDPu/nZPhfCit7Q3X2NHOk6K/NZ3UaJTOxgxt8wYdm0B67
cQpOqpwkqs/sgMxZ60pg7Z3BXcWevd/N0+wihLxuz/9eMqRGeXluh3hHShis
7Xtx6ooDNP+Pmx6dSk7m+JSlngbmomimJVXvJwdV5EgzZZRWroA+AH41AUAK
nkHZW9pcClcDR7+bfsU00265pdVFrE/lGnBHLXe5JCvBswEZrQ1oi57+/Yqk
wY983yEYord0R8sVKTJ07LQQw9fba5BZBjcogkceUyEkrqHWha6xCQhovIit
cV9af7rH6EXfkaAIxQ7tgcP7K2qwaDGEcZXuK39VnXo259TFCkTPsEyBw2ca
7fiJd4wEa3nWdDDBI2vDF3vJneJtX86HutIzcwUhEsA9OKsa79ai5mQlruIL
bvcKyKAdBGAjaDOehKuGtoVhry9o1yl4wlf9iaLTSr0TF7f9dgyfVyQdlnYs
mXcZObqg4h2ihP7ffIzlA4uisa8t2FiuXbaKsdS+SULFmk2zKYqypgD+Hpns
mSeFThuIMx8NqKl2oobcYhLkHaF8U1FLPyNAMh9FNdpgZ8671+t4LritPlij
lzC5XztR5XBa1CvAYWIekFt4iT+0wRJb7Kp7np3QRSxj2rhIO6KvyQ9GMPVX
oKDHZbUCR5dtV/d5AYp3AQZfz9CHANoJd9yVWqMBOrKMZxYKhvoOE6znH0yV
r12yKwggmCIADRZA4LXmE3WvxxWLZRs8GFPcRHjp0sfetowXH+q8MQge1oV3
jawi3bPAzuS7ElFyEY2M99jA40Z6AztW9+Y3o9THDtAR4uOyMt+i7AwiHNkS
0RwZrx8S547ZaJ/xRG4ea/vghdxzRL1EqSAoSfavTnEuK0dJi5J0e3zadp9d
Oys46X6P9PpgyWNNIe368OUSwqJucsKlLDj6to7gkYsOqp+wi714UHETs6hM
pOZarqkwOAOl2vlS6KA+swWcJO5810CQ3D+wSRskh3W/FAjbOdg8sg1uv5K8
OeIlaGYQ53cuYRuntnIVr694Q0tZo8jQvkK7XFZfPaOK+BOP/o5lxqB/8FQt
qRQAhCteSae11HCIOU7/Ek+BaJ/WWqlmecB5T6q9K3T1cupLs1IdkVPbSFE7
S68afa+uX0ijx3kNsnumsOKkvkBY0+OSUHcWMVeUz5y7EKSt2octT2HZTRvF
PXrdR/CJ1zpveh9FKHL1scSAy7dbXHpYHw9JlWbXjzKsxefuAizJmJG7F6nr
YeWXwpFXioK6UkN9ujROzHBjs35kT70OCJWVAL2/zk3cTOmPOfzKjLShgzJX
L/3Y5qDRc+40xCwp5/t04XzOvzYGZKT6vBnD5ssG1ypK32fP5EdeusD3E0MR
ogIB+tlgPe0I8pRKoXJFGzxdkRqpb9OS0TsxcmFpOwOaOAJA+MxOritKecVC
AfBjI/f8p2htvbxbplBYMzSXf65c7O2OSIFAqZMy3uSm4Df/Na+E9fS4y1+P
8a4/jq7Cak553xE3gkMFH8iPWIUEzKudfYkt2eWpauiZYurGVLZHBQCssSA+
hFMtTTga1KArDia9euI0MPspBqRO7G3KhhMeNdkQN74wKW8UZLKz2xkg8F1V
dk2szkGeVtJWtyZtYH22AUxvrLnQyP9fRfT7FTCC1svy3MuYf/Rh0v9i4oOR
p6TZbgxFROfUsoiO9gQFDLQJdLWwKhqiRTh15Goz9VKWmB88k1KDquZIBxK2
/WDVVY6BFH9PAFKilOL4NqvlVdcC1FvGcuEEEo7qBXxcH4edDnRuozWIGHaY
6pKuS/0C5BlyUEVUEdpeJ3CSIj9R+M+5HBEWtXTg4A6O0ROhON3UwNS9bQzj
Ez8p6PG8uow9WgtNmpCmi8IbfACZ+UIiR7HY64n/p6n90w1gZhU3sHEYO/fS
ddxfAJUXKoTFJE5N8/0XasK6UyMEnZ23uTDXT4rJP4B0KuxAAjRkaDqI6Xfv
b1G1CW1Bp4y+Rnvh4dEooovWYiYFmYVX47ddysLEvs05ghullyUDVaKJVLbq
+Zm9q/ZphLQtwiEnw9FzMQP+bEqLoC3V2/+cX2PJ7BISkV9C/63aobrl2YrR
4d/wUWDohVdwJCOgJYqI+6d42UWreGnMzj/bu3LNJOaXNt6iUTdw0tuOghNg
9+UWdhB042RDHimPbb95eRZkqD5lTVtZHhIUwLjgKgqP7PmWbTkRQR5c1orX
DQ60uUS2D6kgwt4IA/f+jmOtFGHro/WyKP7IvvNQZGyVVUCkKxqv+C5q6/mB
UXPaWRTe03m+X1r9i53EmLrIO3HyyjLGWStGHRYunCbaTZOpda7hVZKNLNwq
l4eqzZeYcK0KS2dveADRDolUU6MyGRB4GzFjM0vzIJxRvwHp+KU9V0+fwQaN
3ZZsYdldkLCEcjPRdjATjj7GaYmDrKjt/3DNJVDe8YlO/BpHTDD3mAAzODM9
Z1Zd0dMNGNdnp6J8nrzHo8VOQI8NQzCLWKxefecbfOsaLTmvZfaqo03669l5
RAoF0jL/PGvsnqMOnFC8XtXkfhMHdlNL7YYO3wF1dizorIp4qzYY/EMNb2D4
w68FSHgxV17TtLL2HFJDIXjWFkWk/51bmaOgF6mCkgAYzpteni88hHe1CVON
z64doJCJ30D/92rx6jPsMMIPIZ7vEyEzuxdZ1LbMWydCOGixOgVToQ/MMxfO
EcO/d6OXFS0YqMWfW8W1efPbr5VhJal7fTFGWN0bZ2s1EZfHB0/vVoKTeLLA
eY2fQEnGrpZ20K3pU7bvRalMfwJs5r5qFvVOFJpbpKs+S33/rqwAmzrfFLxs
1H1iM565b0B2CLcs04Q4OjGYiv8hjE3UF8Ww+MtgI4sDOvkoixs1NSUMGDHo
PBuFLiHUcHKmPDrtMzF7xX//mZ5oUaQtKwqWlsLDv5qMjbSeLGVXqAv7UJ8S
c6V8GYgbAzXlMquavlRQte/CTQz2tAWMKqDezkBO9YCHJGV7cImnDTlXFYrl
U2i3UBHRafvcA/D2Zj0H3mniAO1KnMYxwjVaBoFP5J2vTpsMUqmCK0P5vKUs
aSLfPQDTtevvnyWq9BAOPXVwjDVrXmYZkTQ9j3rzR2KLbLzeirUfL2dnwvAO
GnXlYhkBuJc/gTCgC/+VKBs/pEsYVWjAjpMuxMUNaqBEzj5GtxBcv1Ye9Do2
QzgWT4+FjY0Y0MQ+dFxFwCB74ZFANV/N8Fu/N/NZFrzT+APX60Ntdxgpix8+
k1ENXriWxn3Ez1yp/RvFmeuvN9N8ZR5znVJpipGrqM0eg8T+0ZyNUWNNwWAb
r42LeLb1tdLdllaLBbxlB2w6/bZa+ofhx9LEWxySmeS0A4QTFraXDNOelNFJ
hauPvgqltJJzvsgfizbFzSO6yCmtNxbBG1PJSQzlUnq8QPVzQBdcvolAoRx4
t8DKhh1wjh1jYvUdEuKeXW+92aeORMUw42WhwZsJcOeaIIY99RNGU08WXXPO
1Q9J7c1os1qHDfFLcOQpEXJ1/Pn9AN2MLKWRerSpzoa5qD5Mq83O0kgC8MI+
4evLdEx6niHy5r0WOA3k6oUFbfqDNCZO/0PYtDdWa56wTYfxendyK+QcrKjw
Y5lFdyuNf/m96Mn1BW+hgMI/ufYJHN76VRQPJTKc8Uq1j5T1jcmq6dyeFdu3
46AiTOOLP0lP/HIE5b30bmlU3nCjjcOVUyXwanez2hFEkz7fc0sGCGqO/SUc
FU9Sz3CnRlkpR++K/xBqzJJT92Sz5i90n2JR8iDijA957L0PGtZaQv8agJat
eG1J+mW7R9yhBi7MzmdceUxxaoYWXEcdleYnjbRwWPYc9+Acfyw4kmIxDjCd
9qUqXXSF2Ado9wFvzf9Xqbo7Wnm4FmG3rQSrPO3TaTXNgMw6+uTmxNZcEdNb
VHKmkEkidDvHDdB73qUSXOnGPeD9U5NMktL3y6llQRnfULfnG0FtmYbu9jzy
iru/o4wbam8KtBTgKyzZ34athdUkdPwJ2h7mXpzg4M7hYoeUtPHDLp9wFZjr
8Pz5IdFvYaq+S1B6KMcf8U8JZ4ysMFiCdWqnCc0qu72lr59fIF7BPYBzFxUG
Yd2rQsPWWzWjvp+cK0XnykhyJep0GGtil7iW7lRz3Uzl1Z4spU3/Yugn7C8Q
559jPeIQ05Sfh3SI9FdE2qtoIW63EOhBIjfyuShQqGB/ECX0+Sd3lpjhRmab
6xpoCnsFygdWfLYaOgv5XQC+8NJ0Oszqod0LBn8Z+VCYM71PRQQMq+tLNHQd
q8WqjYowiwufHIdb3zZH62Cs9XOgN799zH4hk6RDZLjWI1iIK/yap5veStNP
Fwq4jGI0VTEK3FWqoau8H8RE6Gvgg1xabHQ/+5G+9TUSWkslkYSM0O0fLp+F
Ct+ryCDMQoPikehwCt/tM7GdOG9JGGBk35WMofDpL0OuofnLxCiVeZZQ0b5W
yhO7lA06SK7qVGhxfSkA1Cqq1b6XmVE/kgGyaAnU6ysx11z/tVtazeE2Nah9
r1nkmEM/qNs5IDlxDYn+J3fWRnZ8Un3K4cIuSBKjujicr4zZtKirnCzeOVp+
D6aBvNM+mvfjvIlqcX1MYnhRr109lWH1ieKnLrU52nOzDWoVeTdVRoCKJkMB
AiaAunVBb2ynCLb9GjKZ2Qsgqbj8ofca2O4pdOHMPE6WbstVVR8vtvvi9Cab
5ASfN95sTiYvrLS21q02Y1/L82kbLytDKqGgHbYvqpa1+OuNJ/+KJ9YvXxpq
2hRqU2BFhfK7gHEMmcWctZgi69FDhf8HJyB2sx9iG9uAVkZqZMet/yeZIgTW
WR/SeWP1hAPfijLwJOcEcBkkc0k0/yqLG3MDXY5NcmRYkP/fjqjkH2tQsdHK
TL/8yQ3qw19zahGn6RG1xm8w+heXqxKEAJe8VPysjnx98j85wgTOiJVI+2qC
7GUOydjk9uRdcn4cZpns+hTifknEzcup28R3EdGrYwZwaVhndkF77tvzDyEo
Kntu4lmeQxtfjFAVt47rOrV2UanCv9Hu0bBka7vkhXE95KodE4Rw8kCndU95
u2pxdaLN6MXRyzKvNfdvAfVFE8iUQm4aYvxsCzP4LhYTUHbJvq2QW6oJAM7p
UA8cuy+hv0YgvjbyY4PahtLqS4w/mAWjlthZ+NIm8wJu/FE0ki5ISkyODKjo
UuMvc661ML/2Sgpdu/i8K0DfzCMFLnQV/asLHxXpscG1DmjcFkvFhOESsmJN
GrXO2E/AwFV7gbyMfIK7xYiMEN1V35em/57qekJ2vs0XNKyqNq27v2f9BGqW
XStA+wINvSWCuWX2TVjsMAlXzQpeeHe5+4W12+tRCa7V5rcZTcFH7MsC07UK
pqkSojnXJ6zBvRRtT6+kRnSoVHgtkLjlVfIDr5PqjxzOKUkV7ASY7kJ6Bd05
WhhGUZqiYbBSkEneiEQZP4wlJMILJTNjKlz+H80seYY5UI/yim97po+HSmpi
BoLlDiZW8yxdpxTjCC0r4oK4gIZgl88lOJ0ZNzbBFXUhy3ZrOAJAvlpGCa8P
yZVLmCo7Bp7qOe2n7hN3aFFjgN1783p12Zs8nFEyMa+wQfw/z35vLzaqAZQE
mnMg3rYDc+Lq1aV9Hw0rlzaNHVEC6Vx8N4GMtnPdLmvQReT0/HlmKsh47N4q
Pa0RRiq97mNMJBPhRrZAwU6L2wPoPV02aHWJXE4lZVo2hnCfPjf51ZdQ+kgS
5eDfk6cVVDoJCopYbhcvjXj4W/p8aR0L8vjbnunVJpxffqQVISg3foXUPbga
d/5uVPqICDqTvLkK8BYIU/luwHioO5rYaaTWKvFFrLurf7iqwR6CVcw+Xxcy
HEE/d02DnFT4sFYx+4mGN8xq+cIX0wy8bVhL3fm1gVcGADAy9zpAhhMOCnPP
BbBDUEZV1I/+byOdrTZR7bOtBrGCN9rwydkct+t2+rB9T3b1knuBbDuEH7Ep
75a67F11SL7LMApai9CgNXRwfNig3zD/DkC5K98NDd3j62azATNwZhg/4HIp
grYpUemKCJjWAYq8x1LCPcMPRPqNglEjPeK98fg+KgwnTNH2AUV39Ty3EKJK
iFQInwyHN3KkCL3mwlsXGVILbo/CpwCXlCgkcuD55NrWzWtX0vN7tnyNas9Z
RwaQ9oqdQHi6+8q7ieb6xqDyxgSycdlWZUXvOaEM4N3cNpAlrMEUi/lDDyad
APqLBlaqYkwyvSpGC8o6WLqE+J1u/lMa+h4mc4ntJd5jiYMzpALVsbMWCBbL
GxpaArGoXy6+qSG7S9tu15GQKymlOn1uryBKrYcud0xfSJTvkfAfzBvHHjob
W+D4yfXRdOqkDsNyaFgveoG7wuak3wBsZ7MyzFcjhontvLe7jLfKY+K2Lmgw
UPkp031Exnxl9+uTlUUp5ZpST5fNlPd5xxOx9lpBDkCLhGZtTvuVkC9TwkL0
3cnIRfxU8S2696H9A+8v7XY7HznyjmUjlM/VtlvHP0Mv1s/+pxtl0CtWEysD
oI0SWKHbqxy+2Mef+C94vd6tMDHHg90okXODSAlfL+BnU8vuJg/AnbnC5BiK
qh5KiMWJ2UrA0meQjiAn685zXdcpxQHHAzU5f7jS66PpVpp9xaYlkXFtNMI6
qxmv6p+nrc4XWQcdTWqKScptq4ch0gm/RdedEAAO1qkjtUaN0ZH61nzV3YgF
oKgrQYhzl3mX12tTMo+pXxNojfn+0Jnjp0QfFo4GocPf5WE3044NJ27q2xnr
M3szehhDAhNFElcfu7QCcwiDmMMWo9Ob2vmB/Gzr9ih/kIL7LjpJ3uDo8b8l
Oe+P9wbcMerT2u8bCKRO7Bf6Xr82GUMB3ZtyygxN5r4mbuyrenw4puEwIUj6
/FlejcUdDSNCba2nJdAKEVe7qUwj+eyIFMgH0p/ybBG5SAwLDQUq+/A/ZgNX
zQfLkvqDcfILkxBWSbQiImeCNhJ/UQTFzUc+kZ5xshIOipeoe3v6B9D9w2HT
kfrHeKW8/Ul7Ik9aZp+Aj1zoXwMVI2QmqerZTPwnv5iFisJ+3vqAdp6WJ8pe
h2FYhiIX9G1FGfZZLnoLacJI2MPqL7di3TM69eeubh/YbBZXl/EWuGCl2iUR
mJFnCGbFJRWjCHpG9V7RD03JlKXeNyVDCOjLeWxiS+5hrrFeSii7zrozK4os
f3n23bK2nfDuuUJ9yHmjg64167mtwdpDXnZsGXO2HRoSP2DCQ40+SdUCcNF8
Gs3xE0czKiWJHlGT1y3idJgHPK9b6aeRVq27YjzhFeVaU59DrKnLXYAH35Zw
rHntShnBWdb+/4WcCG2vWBLnPn8VGyNpyIioVj6wSMOTLQRW3mBewx6liLCo
E+NPRCBqCqwVw+aZwkW9iueDPXQzZIwGJTVK9oK8UA/FGZwUmPjOoEePkJOI
Jb2GhZAHUIW/7qtRxDvbvR+UOHJ8UFvXvM5mp6W3hBsH1pzQUpbwnI5CI7Ug
5XAk9CEEkfSUpjLUuwZGS5XRZUROIGrvZYbwiAtX4/GL2xFYJZZE6fsELj3Y
c6KNlAkZWNlznLd/5Fuh04p+0hj+2aeXOfjNn4wbCGEDfi8XG1/nYGcBzee1
I4pgwzgZP8CK7/AWK0ZRHOz58r9usISpCezyoOk00NXhwqFwVz2Up1JGIIf8
aQYutVIK2GLikKPWVEJ0XSR7b0fKBf6HXfLmhRzFRQTdw/qu0y+rgxyZSZ3x
kCAlXMdQ2+EBkXy9uFoSzrYTJWYPwnN0vFCDe3BX1ymFOaooBBIBlFiXQMd0
Pkez9oVUhh6P3Vx5CcPoh/0AqW6afSzOcPLUgvL9STrNINMt5O6fZxjbMAOQ
kQPKz3vKBqAtxBahn8fVUGSlzPI+SyFZVMqonRE1G1zu2wO7mySFo0u/W6+7
U1m4Dc2mCbTI1XGYO2K2ngV5qXwz1flUopFAPIuzcrLp7Msyu1xcF1EZDtW0
ybXkdKTzmymfcTcFLhYygD4BBQWTUK7BsvNY+0MaShM6lntkGwxNgSdPwzDW
35pY8NjJTR3K5Cx2c4oFGA7g/gCkSNuzSw8W63V9PZEJlp/xQlBpIt1z5BqD
tQfr+rEXGj5l39wx9SFDSbNIRjBTwAwh7Og4xgNNY27DM882BxFaVOvkL5d7
Ie4twd1htVYp8wE05f9S74ItWdilEeN72ld7FYlaS/RZ2RgHOoQ7vRREQJMm
9lgAwo93zL3uHxgA9UO0tNOTkmBmYu7IAfuAmgzmFW76lyakLcVv3/gHn4Vx
M+spKc/kb9BWONrdcoBbd6+MTrudwFMYAddIuodcp/rn19cYMbASYTbe225i
dmc7DKcuOrSb1U8lf8rhpMCL0BIWO9lkfC8xFN6Ub1J/m+jxSc+Uh5E821Qv
37xW6I/nHBNCxKKaDOxpD6uJ5OMrT0QwebwN3kkGfjLtHM9JnCTvLLKQnHmx
KCJp7DPAarcy36TfTT07kWxpF0w2YOStQQegRjn+FZbC20CBcZBEfW78yXL3
dZomdsmUwIMIYwiIzGp18FXtGZYd3ozOXYO9vETECbhkfGhZ8EIhNQrmTEkt
GJjS23dKdW267mmMLcGqy5FvjGuxEXG5/9kzs5U08ACFYu6GEZQXzkK+XPFf
hYdq3HlqAw34ad1X81SEkAdPta7L9ftMfml6WZTK2ms226Hqr57Mavjq3IwM
QRbWSb4E57fGohgapRA0skjZPJNCO2i+nyMYM98LY5RNAkDdY/XRAZFs6BI7
9Bge5Mgi/zmEVP+5mlc1/5a3QHxMadItm+CUtFkHpjTIukm/PJUKt8JmZg4t
H/W5QQIFemgxIcabOIpecgpggv7CziKWMHnp+ibrqBCsxEPTHaVthNN3F7LJ
6oQmN/yl7EUIgaHvRVRPdJMQhGUrgRFOJGMD1B/+dsenJky1yKowW0aqdBn4
koTGDvt8ThY8jPokpE9gTK9Oa3ilramiBmSCxFh+0cNBdTB0is2MTDyCwmcY
0QcOHaUsck4OQy7XfwiPmDFT1uuALY3nw4tfSOYlM0VRImI5itJaFaxYuZ0k
UP8/j4WA8ax/GBTgiEtoMo06Hsr/ZFKVAQ8ka40uPjHccXKsMVJStWR+CmRe
BnCXgbpJRWRlmiKWfjKRKFvxWJgaPKscuGjKZgVOYQ47c5SmSvvjZrcc6XUm
X38Q5pQY88N5LDq4Djwxm/QgoDUxwhhER2ujmF1ySRK9Su95Yw+FicE4oVC4
erkU+Gf/u9Q02oEYxSzY1oLj0ErW2p7L4mZKLdJVDf7rnJaVaExkxOwfEOaX
5FqLvFZEtHgHF7CnGrooV3prBZ5jUNNsmX56Mpe/urxbkvnqlIrjocc7S0AJ
Yz7hwz3o+2ObTVHrEdX8NYd9I1mkJWduWtBj4Fv/bt8Mb+r4s72+Ub2Bh3EK
FmsaHnUnVkZjQA0t9tMbvjYuB+ffWrZcewd4tL439Nj9a9LMtzvrKHJxwpuu
Gs3JcZxnFNbrFXt++sM20ZHytY6FfALZ5pISW4lQQVS8KOKqliK1Zvg2y3SM
yIZzp79XfzUuH1bJ9YT6tCiIGwoxB+Slr3/ztEcqsJ+LdZWvAG8nGtOkQcRF
3A/Ic1w0YQwvoTUUh2aJLcaLgFi8HD4NXx9EsAm7wyRqLNCWPEp95U0gwYVQ
zSCVJ/TutDnBRO+/HyIWF2emYDNBzS2Nf5tpCFyDywcjee6/XGd9h39VOn4+
TnRBDH26V2i6HD8uXjVBNPrk2mm9Ur4CHlfVPsoOF2Xsb8VsFUlMz0SfMMHA
3Ij/PAjCZJmk5LXcSlPfmUMGaoNvLf8esBQb2vWB5QVCAh3NBSOVDpXiqMBz
bIIi2kVMHWm68ciBaQLz7dAsdaq3xdplnuPlddC/cBtJV12+4zpRtvqoJDFx
pbgBZkjMvU7GL7XYmMRlY/VPd6LZYzHtWYtN+MZducRX5sF4Q9R4K9O0TLdq
MMt1H/VElkJzRGh0+hyqerzk1gG0MCKu9ZUNNuTfd8fMss9PkxkkA/ZwFi8M
dNpLkcNxfJRT+LvJOBFiXlH3J/i/92CZslQ5OtIS8MvtEUT5l/on/z9yECs7
tN9Btg6cfZX4hCNd/+h5vTa2KIQbpm4P+CTURIhlm4TkSwhrPDuQ+XuxQTlT
NYKr9CAFx0Dd9AOD4bdV931HhxkQU7+v1krj/J8hTugfFYIB583L5Hste65e
wcK2vVDZAaVHUlF93H6aMYxK3geS/uYSLfSkibrWHWojE81QleYM6BQEhqrd
n7aj+btYyB8nvXq05nFtkjbraI5jJWcouGiQzmozGJazpJInwLjgKB5L/R+C
6sivqma6n2biHMlGXIlAOqQduiQK8DEgC2HcDkJzcszqhBqqZWkf6FVB6juH
bDNzWrCNQYY3/25deDJnSeIfVnwoqBkxF6WyaiXs5WegaGC+rHT8nJzsFazv
Rd1c9jiKO8Be1+C4yoAqrYGq+QfRYXXi23kQjo8AAPVrR58aH4gIQHVl1ALC
tKf08KdQBFi6Fdq4xzbD4Kd1AOqPcTRvE9ntLo2LPbSa3hKcbhigpVBOXGQr
WWWNvDK38xJW8GYmKjzQwcf78NOLYE9QrgbJkun6/6yC/wREB613rlKTvWMJ
e8xf+e8eIhIb3+81VC6sJbE2jKjf3fWeBkdTBQB/lIRbFkVWCpqnt132BIxb
V53LpPl38Z4SLjD44eM2I9XR3whkHGL2nQYe/bOAv7xdoCHJTa0/OZa1hukt
ed3lFK9OlMQbIhAH/0x1EpqgVZ9L13b5i7RuXTJtalvb4aDp93VNWntD+WrD
G/yQN9GAwqfKaoeV9o+OhLIa3OOM+cShsfeKaEkZr2NXdIFIXjUn68NhVnE2
BMszU9PXU39mH7ZnV92eKguVaHU3ZYwYp6ikkddIQ/IIfyyuFYKSFV456/b2
JtsCKGkIFO4ONLe3mU93PMgurJIfP3635bkUsamUUlpeVad/+cytNlkXr4E5
SgO6sv3xFngQ23a/cZJaGTFMbqZsJ9E6L5Xmvs9p8dRvhMVlLvq+Z6NSxtyj
UQDg67zdNY6LJgG22bUD47MrUDNf7P03lnOBCGeeon4PAMbcSsMmRK7a4q3i
hj+uKzCvLATTbwQi19OHCzM1hTVxv7l7nxUpLc/oJowM2WJk7p4IXdgxNR+Y
Lmyu9+nglOZ2dAkJAWdEzZwY0D2T5oWT1K4PzgCsm7PaVQuIa3uo8bGsFpVb
7cBL+A0zdhGKWROgXxf5gL3imZOMtUMZu2HYL6YphhVDHvlNkPxTMIxQgL/U
isOx/nMVT5zMcsRc3Z97ybcB+JQ4UPE1+ue5hOEMdzkHE05+LJBXETt/Yi0L
Tx4JbEUeeFOLoXtyqjzuEqVfh6Xdf0SRsdhA8G0X3XKoe+wMZWpgleekzaHR
ym5fSop0EJJ3uiIkldrTmpE6SORyn62jsQ2CNZg4S0SrvggBFSN1/fXJMoVB
klwfEp1SYxt3b+44VCZcL2D3dZhLxDrrrNvnBpCcsl1Gnw85NvyOO8dqjsOb
E1xdD8QzpBjunwViUoz2U1Y1UCO1mqHQoRhgYLqn5emdYQan9SfTgtl+jVBc
Gui3iAMBpxUiz3rOZxhPki5wuuct3HHETkGaEBJ0K4uTCGh3mu8/XAozSG3y
WjKM4LEk1GAKv0OOZSIkmtNa2xLprGJ0CDz7JFKM/3iQWFAu3/5WxcN6+d33
8HJWNBPu00AbiucP9OJuv60pDpR0LnsZBcjGzxyRbRdMZuN3QwIWnRsKr7nq
F94gnO+H28JqpQ1G1tPQecLp8GbZei1Jsc4ReWeWeKIRWWhXP7O8/fnj4FZ9
g1vDKV1apKehGkVAIDOIi41fJ7C+6D1fr1+6I6EQ0Ku2gFFhKlKn9iB7At8E
7Zn2XmfNxg5439m2iSg7gyrIUMCGI/j+wbKq3bXHosfHjIUbZvbETjhE7VOf
2ZwFkeIuiXVUDChfTBMbXOzNlOHzkphGyG8/pK005q/r8vcFpGh0BY8PW5/s
pusFkuf0hJ9fNXrk/acm7OMmJSYDCazXGxXfxgjVpzvBIHOuN/1c58HAxJEQ
E7p80RX7AAT5CS/wJppr5+DvKOUIJ9ukMT8NmZWHz6eiWvvr0F63/EBlrr7F
mmuz4KZEFhmnGyIOOgmVi16PfAA46JAE0Osjt9NvOu8edmwujsjq6cjhEuUy
arFYSA7DlKIN3t0LNASkR16Aqvwc9qmV8dJqR9Uor+lF8s8TWBd+mPSFhZ/K
6Flu14j0JvYwal1DK0amhcqx3iRSsDQoaqm1KdIsH+ikxvJsjEZ5T7hThpYd
AElmUpIiT3KnfzQIkO8f7ZrKS88GoH2CY0qVhqo7ZlnV1Hx5ks18Qr2R7LWa
GUoO0+rXPWI3V+0XqnQnbo8eSc7RFCpOLqdWoZ3CU+8IhISXjaajpJ1NOZkK
9TUw/Mu/q6oETT7k3cJaq4zEpKjlAX3SZQYfR3z0NFhJeelwRdEz9b/aOPH3
KWUXGsYVukJ1ZHxpA+dPn4f0Fhq/6cIDjrbIC3qI5zpCoZgb6tF7sYwjYoNx
k5l4ljudwvPBGN6DmK6fVfaqA3qCCjNX9VXG9opfOS02DOT75xNRKGGr95sU
oPePBoXWmCgTuYZwBnyyedJgQCNjjzXBlgnxbHJJtxbfrd8q0bvFAPnjpB73
t2ms18OmqB8p2vxfMuxRiDa9X+2llut7l2Vbh7oZX2mb3gGO29BnshQEoMA9
vkMlQuEicNl6QnIpM8OHu/QUUrk2xaCverKABxjV2y8YX3xlXCvH4onmHm2V
W5YSgmx1+JnO80pznDaMnW3pQDnZFnYKkiICmJ1SyAXGyHCMz7Xa3jSRgN6k
kLynwCuujUm0CHvqzwoYocz+UhSgeskHDdfKLEtj6SG9XYyQ8GPoNHUmcTCl
2c5DcEgR7iWNR+MlrmKJ0N/830JJZnhhbvDq1HTDTXK0wu9tsjKTucC6p9qh
q15BUe1JjWRwFptGApxhnNancm+JhMpJE3NpSjs7bQrb8fX9HehmwXwggG7f
06x8SkMM7Xt60n5m4pndeiq60tHAwrsPqJNokV5nwnrstPjoRKqOUZVcFclJ
a0FxhYJ1G8fqWmSyPq0DUS9syfwjg0KB+2X8cqVHigm/wyvW8JyufNNoqasf
HP11o6G2eCW1Dpg9ZTFL+Cz1djFgn/kOOEmF87LidRIAsDxemwQM7VTkbR66
BmOUPScKG14W0rdWHspbSGYiRxGyyEsRe0JZXTCEHR7XKwQqYrw9ikI0wtV/
HK/uVd02hF1NHRgx4tB5GBKNQ1Q8z/ncqt4Od9A4Rg07HsOhXIjoCHS/gYGG
ufYpEUcyPpR4D1AXPUwU6agE6UyMqraoOvHhBTv4Z2HKbIjem958bjMYdHFd
WS6do4c7hXDtI5Qla6fJHcPAiAx8sULGchhSzElJAMlF4Umo8a8/K4Tzh0+2
P9tMk1WUOYYTmmZfdwlCpH/G2FHyWmlpDqVLlRljBfRxvQvSQjHdCH+gst4g
6YSowaBxPr9WKtMG24pb3HLrUHf6P5mymmSViPicXVsU42ElPhNA83zVU5Tv
wRUO8QCX6ssuEdSESMkmC372l9iQ9iUpoBToalVpwFLSitx/r/IEcyWrAXYP
hEmciJo2kccA2MXeSqCoD/fkiExHr4girhPxEjfFK2kjvMaAEfgRmC8vsOad
U2bSS8Se6vGJNGfq6IjitwJ5ox4TUjAyn1Q9Lmqo+DDuNOxWI4IK+cZlle5x
fJvLSyf9e/Jtrl2mhyma8JyWKpv5KYy7ffQ/ephDJ0w/sxguFsW6n2Som3Zo
iEDCokcQ6deyFWL4++k2IT7GIVA8xcucisQ6aXzVe74BDnk/jRqqkT5h7sZ7
Mpw6NalyAMf3IeawB8P+QU/VGPrwd2afIq684SoHupB0fN3xsG7DjWFySjtZ
l4ygzNm2yndmRZ78cI3Gr9lzqU6tj/7d5WamCXiwdkn/2NhHN7oDD5oqR5X7
4DIGhGAXavT2ZoQkDzUs5IlG3Ba4Hv5d4UYii4NoPQ2OJzJG3LurVw8gHZIY
ZRz8ZrWSAPAUG9CCQwMog0wZTragWScbYNGtJkbqF1HRuRWfOJKODIyORFJ0
PfD6PR0V7h6UsMSt3GMCiHwe04N7HdRw+5odn5sJ8UalLnhNLLDeLSWDRvYs
l+0sMiVgyCMOq2uGUXxD5RHSLX+4FDbESx/VYRto7CUAhWCoeHGpeVkYFa/S
uOl8kUlbMp4pmsXzieWnBo6NcrZulj+zlxNfeDm2H/GtGhXXpImIsLoMG/yM
6koqHCSfgNRvkUPh1AYV3x7WyOhBuLWS5NOzwrcwEYnkaqBx6CbLg1b0uyJw
B0R3sfajz+wBE6iGbQocFOwuOBqionIl1rans+G5OsKlSlffNjgwPptnweG9
KSLyIBcXdsllkP0KigWxj3dDwK5eh3FFpt63vSeqCLO1UvCxWzj8ImSJMHjV
JPlmHsm0Pw1i24DbJkqSoKnCkPNp9T2YF66RHF/QFRpjUKtVDFEuE9rE3dmq
aGkup5NNzz8YmPBVs2hYVIUFdisk35o9sf3c2ii7LySw5OwuPx36tRnJUX0X
93W2GndJUrgjoHTxC5YlFGNARj1zu1LBoNkwrFUDE83LxjyzJkx0vBEMhH9v
SF94eaHrZFlxTf/Ktp71yDy6m//If8HNUOUEJ7HNZ3YheLa24vbClSeylCSz
11v3wr8fguzxaCOgW9VZjRc4q7wmdwgmU4KP8ySUV4sdZwomgPqcC2hGQhVF
VEJmzXS9i9rZe7rFZD+6b0ZF//TM1+RRsEfy7X6FSItnxiKGfTTYaUcMeD29
n1GYAIzQArTGpWjzgqbPkbMFhi1iuv80dfC9blkV7rGUDuKyF6emMbJjPZvY
dWBwuYx5v8tKa3XtyNFngXViZXxO/g5HSZUfWZIADhkFWUUa+7Kb/DUx5XTf
+2YE4YYAPedAMJxEzoaNfKngAiyncoyC2aGlyvbwOGvvJMhdDd63TeTOSGli
lU6r7GXXUaDiOc62EUU74ViwRrhXgVLube8Gu6YiRF1Cb/CHRmafNdOydCvd
Kx0hoZEsCW/BTEjWjy6gwxGKZTDeb7TmTcYl3tlelcUC4qtAENNawvpTlc+k
Is13K/LMOof/xOgPX3uJh9UcBkT7/xF83d+sqgBVcxcZ/Vj+yBQ116uGwqlW
ROLZ36ELoV7cUT9P6K+RoRzNHZSyh6fNDZ43lFwowAlLlMiEZUpZDoQ/AAH8
wOwcZzojDzMPmYiIyNzTLiwlj+i2/t+P+RDiQG0HaytLnQgkhS/VNkBzOlsL
bHcEKqxQYO06bcmh7ggnKE7KWkzUwjtZetxIJ2Ci4hMP3JgHbVO9PqM6F9LO
zqG7pgC1NMhxRIb7zJd710tR58ekLAm+vxwJjsoiDN59oZh5NYPGL0EZTF3U
BxcvJnf/X9GlEKEgsU1PtrzatEe2OZY64PP1PFSYe56DxyGYN7N5YsaenSmo
tfUz9FAHpOLPj+83KLIc5sHh4eb+5J+SDKj4XfX/gVgkoDf/tiizJQYfvA/i
utT4bZPul4Q8VF3B3SxHZ+ihrwmCUVTK13dsxHI/C1MOZvlVH56/gmKmarKM
Btk7PEet/YHGdkIx/3l51LeIT0OmR0IXj+tUS+C/EFmu7L7TLfd/s/8j98qo
apitj3UjAQzAWj85IMqRsZbqCk+bIdjHrMJ+EjNLFEycgJm5P0qbPl6ukxHF
WUBpHT6Q36yDlYPscAeT3hLcVMiQOErwPL/BIidIUdVsfQ/NUY+FoX8SDfij
/49P2CBDGtzZjLC3teH18lsn/oziqsjSuGIKUf2LjijhOmqj5zggiPBQJmys
bzq5PtFGv7glhfzMsLapHN++k48Y5VAtjE/OTRvxB3T5Xbqe99PSOQy9DEMJ
RmSOkgrGYur/Tr6TI8+j6gT4ZLLT7r8gbU//yUfBhdrJfykiDUgsBA6xapYD
6eTClskN0TS0BZwQPUVjhDtwS8wfVoxRnHBMC11N9YskiuBbbMS9m+mgxW4X
Fd5A5IAPSMWdpQ7R2Yj+vJqu5rLoIR9gnh8f5s8hoCLHAph2Que8yrovH719
tn1MeeVDokAi0GyDpr2OzYzpw+ETgUUioHEJtyr1zX6kU++Ib3Fo3s3xccrS
4S6+5Z+xOX95iyXI4J+WCdXSw4zjq7KU+IwpWqIAGhI8SWcZl7YHDKP/EgdH
H/dvQ1c33n/jv9DeKwRQMsNQnmcV2dIJcCwhJG/nGyOtkb/10UWocV9Qa3v7
zK3hu2nAbei1yLPJdb+lwzUqeQtSdQzaD+DSK/82MZeYAVqO/Qw5Dtcc/KU9
3SoYaK7ZcqlBTCJbQx4/Rlk8f+FJwn2AJBO9OSLxd4P1Mu7Fbbx09Dy5tfFZ
RoawEKjobUhkaMt8TInvwtxXDS8+2ZmIoL7iX8AEKbMcczej4yUqJeI9FLEu
3i+IKflR/JGtUDC4G5ULhdusne+QZy6KLL4ewiRugmlt2TSpPFFvpgPk7dJg
dfb5wF1UgfjpkovHtLO1wKCCqBK3acRHvSs8qNMNmEuoL+NVvpQzhqoyedoW
iTyL56rrXHY0BzHmJ+9utmKbIoRaI69PbH2yVe9SQ1FArI1CFu0OIHwr93sz
Iz3JGj1e71OQZ4i5Kt1ZLtCbAXJgWZJm4ZHIWwLufRDFbskM6Im4j2MZ5nVh
vPW53lSLODouHZMx8ZpcgkeBPfBCgPIgesdgKcmVQ8CL5vrh/CvSqbU5LYNh
AcM5zRcR1YmHJU84mHzttqyrDqlNl96/uLKOiMNqqpd5dsJGV68KDWNDUz4b
nrkwYLweCwDhDMeA3/mrLZoX1zJHCY+L3WHC6nbvuWMbPGLG7bFJOUugJJ/S
xW5+FWLEdSOuYYwj0gEENT23IUZDmgjv9y7bFPGXOMt9dxutjyYw/45dUKLP
QSmuDCNmDSqwZvnx7wglatVUX7V664h0P4gkgs0ugqN5FEHoYjug0Jbmkjmv
GWeUlNb6VvHjyaO2DdV+M9BVHfp+DEbNs6XhLVZJ4pS0JZ1/Mq/5Y1SFSCVu
yaxuSe0dj6ey55NHmJ7Lrkr2Ll5sUxeB0Ja8pem+wkYRKN0peoa5eiw63ChV
m2grcCcOrNu3LQn9CehGGXyO//ePN6Yb14hc4l5ZcT2wwCzRkFZyRO17zEBF
pvxEieV0BI034wVgqkk8wgKHDUiM3WaB2/eSddJ9rm9URC5ZbxRv+5Ethvxo
YnTNu7Lvp+J8Y7SbVKhfGn4lWDfPhf+af2s+53zOgJegNZuzy3AeC6IT+XnG
62uH+gS1yyN1qzY46scOlPdnyuA6X7ABOdTXZ19qdRqBMjoJ0BTvGxFi3Uk+
utRJN96QcmtVsTXibq4B8MeCOBv2pV8Ss2n0xxocidb1negzV3u/XFOGzASF
JEzJUfehBnCVSeCNjXS0i4gNjvCuima5oG01RcN4FsKdV5L768jlTC2dM8Ke
9lfEgBE59caCPPHSsdsvYco8yCd3UshX3ocudQU/FUgn4/OAExaBagWlDfuo
3FyXqf2g324TGBUdbQeufm2hDUWb0FwuB/TdtpweDGv2eg8BMTY85u3pGJeF
kzQEqjdqjYxwYLziQGy3jx1xHQ8NbGb/jqn0TTD8UILvRYLNxKyfIPI9anX2
jTZC0mEVISm69TVfn8uQjg3MKPiGa/YaR2gmYMV5hp0u/yPN6yRwjvmtRLpa
IoFXcEuJ3bJ8nxdIo2J6FWj2kwXO9i7XOcwmbVYgavJzz8AId5lIW8gfXII6
llP8yZO3UhXiV2c/kJyZh1D27NDKSVnoYjasQV4/zmeo/R0X0SR+4KOLjgCk
syWH9rlM3jXr7JGpPFzEdHSMpCeZQDLbVfG8TXsqiQLFpQr8xYaxH3MSM0gN
y1LK5NFIuDzmi9wn0dzRnlnE+SbwX1VfvaYiVPx4kORDnwJnKqFcG9v3m8Qc
VUSIDOq03somn3w2kktmWyCHe9qEaUt0pGwiULrVvv7sdaNKffDO5TAXaO4e
IQEXXf8a+qoeA1UB21WhYF0q7As05VYmaAH8cnimg43e7GbF7IVccx2339hQ
H6PnCkqzjLN8I1UKjsDeFJDo4rueiPgtImL4MgdN/6lh11iPddPHzTKXBs+f
O76GqKskR2JzekoP+MUmCgl8aUFuGmNfLk20tBANsYIPCzZnd9xcMsd5qZ80
3wp5za/jd1t/GEpF3JMHi75bNYJnQHPrsyapohVBUbP3Nx2sdxQsRPu92l/i
mUKRvfeCgT4Qzd3Gm5z6LBHimFd2LdA5NyyYkp1pM1udFxV4bxGeDIpZT8Td
z/Kq77Se6BAZjjjSlewqr0j8rHkLujBdMpDXj90FL7XHZU9mdVaX0GqgLUtA
xB8+hRub4N4EyKHGohNAHNulHA5LwpyWn4yV9+abcBdt4TSGpIbR1YtExMiU
NA1DfsmA4MbT7sZFWzf/hCcvUghA0p2p2KuIL4O9eQB0NtKEOKj4Q+BekGos
mm5O2Lu8qm8gspz81b4E490frrmJUQlT8C25N1x6pxkX5a1c6wGN3PdF1iZY
v17FBi5mo1AF3PSjbZYYhYWdXkCQTFSHrVvDtLxlZMosSTTPkDA0PjOefSm8
wtJe7DuMx4yd0FaCdH0zEZfGO3OijoTvxs2Oz3sO8TpbYo10nRasAtp3AWBc
n0QKiE5MDU2fxeilkrBsVnd2ayD+/n+vsl6v980ar3kMx+jTmrQdD8TK45lP
j3T6MBla09uANRrTvvJ1yXsLHsK0jU66wRt4TdJCXpgaWWnJRuKeqnHUxkKa
IdrV3kGXFBQ89JC8UYRH4/78aLUwcSdKJTsvNdBS5XxIgdtw7RtW87Uc29oL
PEZxGgEGi6CrxQGN4ZGekb6TVXSQEBFMfzHBjhGCpT5wpg449MO6jLDP3Na3
rvC9M4gpg/fzJ5/HxjEoG68tEDcxN7WIBa8LnJMlxKHUrFkUHZbdSALm+bKp
DC0uIbPqD7nhMjkwlXlTvjX6FLsL9ZfqcB4WcAzug2ehY7Xy1/r+qatVo+/F
OM1GGcaoNNnvyrwQ2cJtImvoETesif07ph2vFZ4ujQP3U1OQNcGfGdXtncQo
OxpXun2jXprrNllGqSicXVf2b8RO5uiBszb6kVToJWp2z6umKnMfOF+FwY2W
uzjAwcbP6IW/d1rBEPIZKCuLksVvHY1cSK9UIgz62h7PFacYyuKQv4EZdQvc
jkatxs4h8asipnYzx7PboDczgga0jd/qyVzKFQNpvpu1VIRKDsTVxpQstrks
w5OVXg7bcrS05oCHjSavzvTkmgTDJJmwjmXpkgABBS5ZH/4DviGrQ81VBOUL
8F3nYGbWkW9EUx+EaPvpUZbgMgTiljbwNj0Xgowqp9GH/lfC0cSgxSYfrOoy
ZH+CbpbFBjuEIrC898n9iR2ufus/arFAvMqy44k0IQmYHqS/EUEiS4xSQpwj
uie7k6XwaCUtCLNnHrvX7VU6DHFW3qw8Q/BapA5fCbMwe3d/Q85KrQwZhLEq
dI7AZe+rXnDEb/QambDmJDTmZnaOWTy6XBxPx4dRDTRdmyJYdQ56QoVyfywb
Zr50HeNvquARL5t3cJq7RHk9OVdgIk9wOUKhDNgvgmctqK6d3DNJFNQLmnY7
0zrTb/Sd4gfySFVyulpGi9CNgyO42xrfYw0H2YpWJBsphPL41sIqyKcEt4o/
sXe9NdJpAxparg+psGXfpGomdM2F860djFaRO8gF8advzX7FYKi5hLYd25xz
bVXXOms7ifmgMy2DAld6iV1XZtY1BNB3gJ/S22VTcXmmrCz/0VtxqeI3FMH8
i+HkXf3y7C1bG73zP+C18Oglg4rcmfDtiR6xTYNqUMxrC2Zzx0VqNrwjAV4d
H/Ss0WxRdA3D/D/ZJB7fun/1wd0LpVmgKR1vapj1bTCIihMn6huAlz9p7ex7
Pwyr9s3oybYXewFws6+jHhSSd7P4yDIBwQuDWK3blBb302j+KYpwUbKUZjls
QZQRY3sr5aJysd0LjjfqfMDsL4p9ujoA5dKWq6H1r1g8ooTqUOtPSHV79hSM
M1uIFNLzE198KRvnqJJCluKLUbe2cdlsWfJWr5eLbduSGfRpCFP10qBZnH06
71ppV77YjcLX+kDMPpV/30LUY/XePqgErfHsrHWr2PUPIEfcObyY7A7ZVa2F
7EtWNzrf2rHLXviIqj8Od8GdFbqMbkVcKcNhuViuZw46Exae/VQGnPRaY7gE
XbEr9Koibnsk4P+lg16sOii+tj+kzK9MNsNCkVBeM5Mr9ctueRrP2MjLxjaD
PvflcM0PaWTsxqRlHInM5ZzCRe4FLPeIbJ4+Q6dDqvDSTU4xq3/QbyeXl+Uo
T8uvYxTc+F40baXChGgtX0wGjwOKv+jAtE4J5NOMpMBvJMN0LR5iKOgVM/W/
lPtSr2HGV6/ARVHnPz3egB/b9lBcek34zE41IAPT66ODLN2RwfgwKcuoIPbQ
5TRb0vzzzHFnD55wOX0oWxVvHlfm95NkwKpmlwNDI0FYTdSJBIKVTCP9+IJh
SWWhJ7kJFl+k2dr9zw3xxseR9Y6UKMK9qGAqQo2X38ym/ctgoCf9UHqAcrTO
RkX4ox3qLcRWKJldy3NZp3OqW9bz+qb8TTPbAYGkv+0ey1Gu17NexLVk66zv
Jg2XgyZa6AbD8Qvj1rtqK+IpVxqEqXpeoIVMX0QBcMxUo3TjMdLslq1TyBGq
edC18OOue8nilnNmWZykjoh3i+6+f+HdpxbMvuQPVDReN+uipe+7yXQtew3Q
L3PkMdPwsPDXnnBGicvosyyKdvxPPyQvZabEoTk68h8c0w1mjOg6cEv6izYM
COYAOAxNkjwL7YTtIkAbXdrVOOZNcKRRpg8iF0yGVdRriLXixDBLBHBStu6z
2xF9imoHlyAxUS/ydQdWYG7LRqKhMXz+6ZIH+FqR3iM+XY4c7tqJznFmJwrB
tQ3g1dnGSQpB6qlvJNlNBARlqYqW2rjUVZnyVDOvNkbYLtR50VPt/OsVrd70
Xe+9qktt2fZ8maN0hvdUpP0lutZN2vwq40N9zeU4xA4TSdKeQlbcUUUzEAVM
fC9vfq9NNUEWaLaIE3neRfpFNc6vUgn8x/1LqNWq0Al63JrCP+mP7RTkJnDI
ZEXaaLUKzynRDXoBAUCWlrtMCmMX86o+1sPqfWJo5NsM9sk+ig4U8OTnbPqk
m+Ef+M3NFPsRHjxLeQxzLz0RcEmf+m/TrBn16kAFK9Qjue87ZT0kjw8DKKro
m0y4NBj7Ca1GZTz3/iFlCjCznOlByuU+U6lMqyh+K1hpMIBWkXT7XuHxYVQ/
EXXIuQYnoIWsEf8PdITp9F/OQDnZyMdfoGdbVvuPdbiZNSR1N1/wvR4A21dF
5X6OE1EJoKctDQeTlxedL3LqkF4IiGBNECqamsfdvnt6c7MDX/MWn+H4Qgxo
KoD+Mia+5dplYGS/0fHn9G+6lgXA7BMUhHDZpPUaqd9NhUt2IZ8GeGvmLm1k
X3b9F9pdlHu/BTkp+5K6GZ2SNhyZrZ6K4ZEfzQjM9Oa6GVTGoQRExtxBoCJi
dmar09NBp/pE7CknXsgMUEHtFxKUjN6qnyUTdB1n20WQmbS+62TbUaZa5Gyb
DhSeil9mRIyjK66C5OIbuyd+c6md+Tu0WIpDcOo2udDdTtGZP82hNA/2x56C
oXBWtcU+On7xkVYfbusCIHlo91YslT2R3WX6ne8p1A8BoTJApXQxqRi9TSn1
F5sVf81Ia//Q1X1Wo1BGS7AexEQdxIYq7Gkk088gg8tvvmvrdG4hRQziP5RV
cAJeIloHxVg7XYWA74isJvxJEKa+ud+ZqHqBe+buz0MFJqYubxEvj0miGbzp
BSq3GLk69jJM1HOuRZGu2bilXGGjTfN/L4kNh9zTIoUzCjAODB5hm4iLDmPp
7joN8yZgXAWQfUAXvtyu8vm2z0BAqRSdgygxBeg4ZgwbyDxEqKZi7LC1mnbW
6ITa/CO2zTy/HcFLWIo+MUcYevvNzrrEdhYeY+x8DjeMPVdaVo34VmVGBVb5
U7f7Ik9EXHtU+Fq97cY2ALWrEGrbJ+aafrtAoYuwULLL3CEQktVsbCnTuse2
PEIgojeZ/HfxH3mDEJSNxRfGAG+dyGMcr/cntKEkFSXLir0z7Gv7iXr3/62l
OJ/btDx+NZ7Roy6tjr9yWhM/iyEL3phh5j7AM3hCn6tHpRtHnk+2oGUF9DyR
pfUL6r42vBFI3VkRJBN7RVfzaFaWQi3wCHI7aK21oiqi3VHCfgtbHsXmZnvL
EuWekZ3itgKbGDZ0vF2mV+thrg0knNXIqlCxfv0PkHwdCknAaLraHDPAmz6o
rCgGJ+pvrgrZeMr0rRfs4Aje/KcOTwMVOMb3V/TuYiHkgI6D200oiuVS8or5
5Cql+0PATOrhN8CrH44KMGx6K1l5ZhfaYmX1hjBY25QvjpOJDPlDdTLWDDEi
i22fkkooZFBp4de5qeXEnuj3a6fOKgScx6XVfVFfGqvj+2qPtomKnVsb6Ddy
aXWgprYU5yWLFnMpX7tdnuFmF174tA9BjLVFxbcUFACek7JVzO1aAQMAePHc
TBmKmSjmllwks9FqpX/ZSqDCaY/ZfXP+++YL6p4R0u7m+0LpagxirWAGKbZ9
sKkXKUI+mtDFpiG0DaBqphtBvutx+0vI4tVlZ16XiJNkNPKTYlHZbm+LFLDq
oFJ3VhpCn1i/raXaDmohAoCQOTx7ljbMd00j3LMxYDPc12uc3u1NVTuEBqcE
P6cVmZdOGGEo/5mjcRc7qPwA976D1wbyNWWuY1+mC3e0N83uNhoZACgIkgDI
kMKKGuzDNZfWsE9MsTKp+y2cMqs0MI0BGf1wLc/C8f4bGrUuNhP814YYmK1O
54234+Ut+pRHfTimyZ2wxZM6rz/cBhjs+QdZpdBNP7l0pnYJcX7D2KG6YyUi
j/2X08iePh8n6/kjF/Pc7IMJyO+URANcMEriVIv5m2yggrN6Lj8NmWKRp1Mz
EqYstOcJCTeB4i1CyxHdqJYLzxge1aJQipH7LgsT6E/icrOg5jfnOexdVSEd
FkzjPbhH+k59thl7s+cSxp7sbSxLm3vHRNmun5Rd9FTAIPMG8tOwkE++Ljtn
grrDBvrWgdmfepsXgifQKCBCz1MluRIftTfD2df6kTWYWhyWlyklxlATeXjv
1yV8oZNxs1gH5Io/FgvgOZri44RG89in+EeqOomLiC11z7B26ZwyMerM6+50
CEGIvtAQK2SLWFpqZ1yuy7gN2Nbm5vYABeyAojwF5Hskf30ZqhtWo/K0cDcU
GT1xVGydHnE7VIvzvLA8fu7AAlvtikJjIE80JosnSewC4kQzQTJ3Oq759wG8
BIzYWD/YPdfFqiMQH5o9+EEKk+yIN7TiqgHPnm8hcD4pjPVsw1/81DZemhuO
ALzd00SLpssZsvdgeIkgHeEG8TWEPN45gRPmbhXB8yQBeLbpuflkPwcjtfYS
d2UNShb73HveVq6pUk3prBbz+KJvcyTkNqKcYnckITPSurOdaGHQFD7WM/v1
h3vGGzniuUx8n76eATCYBj9nhBnsn90Ppx0T1v48YzBjzl/dk2/0Cqpb6AZb
35ZCO/iie1mRP3YAau0rHhuih26QKkyJ1IpRLIEyXkC7iS+UdtJr6bxlMeS2
bOe+VR4VVF1PCGbinE57qZvGU/1cvsR+eH9U56q9Zb3n8WNcnJAEsnhArC/v
i7PqiE1AABXZfUtiuscgZ9UzFpmn3C9Z5PtBUN9MKbHuwBumFkhFC7ahRy60
lIxF8TDjuiGQnoZ1uX+p//CpgPBupEtLzmwxbq4G6fXiNJaLs1W7loIaJWBu
od0kXk4npXxRlxiM3+mrexNtyWZkXFE6XpX0SO1UMnDQiPJLK681zcOVguaJ
8k3nx+HrpM1vA+lMEWd/zUGEC2fdkvDDACALi3d9v/ShNvQKP3vBS8FXVqk7
FSSHXiYL+Q0ANgHDD6pCTT6k5rUMOTwERbaQ6leHSIJ9SAEa38FJpdmVO47h
icxs5prt3BZAGVEgvgVE6OgSbEO8UfvEJkLHUALO87OgWHGCAHlghmoS/r0L
Mnr+VM8bFimGRzIp7CDsFsuHBdBXfoOiakLURNnjkXYc6QdBvrd2m+DcEs0A
M54mRPx5ni05V6qlTSQnLAvXCoxPP6Hs4Ww9NhSLZbdY92h/dxbGYvuE3V6v
YXFiz70XiLhw7vmzLFvb9CNdNqSw02avss1pERBW2geDqMC5alMt+Nc7PT/O
dFTJv/AUVG0TAjM7f7UEiNRRefWHogtQgte/bgbBm6Zi4lphp4BsR4xEaoqV
dOA0ZBI4FD4VydDcM9rAgVtQK0HhRdd7j5BW65mWlsmIMM46qknFgZzqYN5r
S92Ck3ypn2Xc6C0A5AYU2QuaK+DGp/MPFdGY+tGw9soBmgJpLmcWUvbw2jNA
bvhoer/WS5EWxDhBbD80ogEf46ews9gh/UpbcLzAvdJHTgWpKYL18TctXcAw
/Fq/ASskMFqcPF7Q2SG4h5L2bBZq+Q/yMiwbIs13kEwJaSxtBu84tktd9YBs
G9pHoOu3ymWqTOnK013e7a2qTKKQK8S0PDFQKkZ4rCmIu72CrD5st5nrxQoS
+VBixJ3XsTI574Aq+HdeP5Gz21GCh/5BnoCoF2W4Q4HMZ03bcRA8awmKChpJ
8ncCkgWUzfAa+FxdJwVeTfTbF1DlWjrr7riVYZ+KgG+D8Is1gxkRflonDnF5
YetSWGeJdA0kJh5pK0vDGdxkbjdMbG4fE7JSaUbvrO2JWoS7Y+WpFYPuNQME
Qf0+In8Bq0YAKGcANUBM7gPYsc/amwJ1iEfdxcXtNmO2Vsl6x8dHBxIdWLhR
KQsH6fjKbRBEze9eAnqTJ2sgsjm8j3kTZEXRMHRuYy94gDv8E2ckVa0Vpvt9
2iCNae/muUM1LsI6KeQGEG7r8uDSpqNe0tE5+bQ5SQ8AMUOICl4SC5ID8KL1
0grG6DSxO3FNnfw5+6SiZFl0mzAKFMj5PvZUKwcKk7WY0dLvQAf+kQdKX+CV
SaKFJIWawC7n7A6dwU5jAsNUMsYD/64GJD+dyazRf1FcNQY9jB7Ki5DW4zNy
1+Gb6REl31a+3VyyTD72PKd67DduMKPc67YyninUow9xfbDYQ3nxD7ZYknC3
Q7ALBt0+5VcZgfBLIKD2vH4ie5gvrwukMQmcj/MmPqBfsgGVj4LCzXOR1g3i
1tQy/NgOvGUvJcB+6tUVzvDCLxNmu+EZZCLVxvJGoJwJsuJS45Uw7KhlSy37
7xfhgD1JDgHAsgsWNGxvR57vOdVWxw1rfgbq1ZEyUMl1eJhQEIbGXLCfqHTw
WRWO1b9BpFxCvgQ7NEVQjKp5IXTLxB30/H0UVqljZLMbxgOZZbYZ8AmkdAb7
NvCbKIL6Z0vjA/4pUjDDVSTHpzcXhKfDGNFDwKjbXh9Qd/BdoXoWgD7e3BsE
YsrQAoNrhIAjHJVeGYT8pwl2Yw3x2erl2Ekr6Y+JV6W689hNOR5ykRCheghi
BvfqS1e7qc6WtATSHKnLj/CHWxzGTvZE1dR5Du8lU2ZTpdxx6mjeNGt2xl+r
3/kaQl/P7Ped7c9EXAsHrwDF4a/TzL3JnyDNfbyPOD7ynVyJamX9dVx6C28V
/maCOamLmRYnULoTjWKDjsnpMBHmrUscjoP+y64eWLZHDIm7yAjLoF3lH0a8
o8NciwgpmiWBLDzkw/1KriORRrbg5NpYrXRhC2N7ExivORoeUwMHLgLxH6G8
CJxX5DS5vPzdldnR5SbvQYmu9NKD3WHpMG1lTT6pqc4aDeTuu7yd48BtjJ0D
VaehZEIZifceIGIZjbxfyo63mLRQFbkwE3MO15wZgNbazfIN8dDbVh2vlckP
E0RTifHssCuFi1UTFHwqLwFoIC0U7d265M4exRk72QERKbUzp9sMwFzuW7hV
kdt1e5wEHVYEqijHKlvvEOdhUYMivVU/7G7PIo0j8j5Wbjj4d9oSQoVPFxqb
UQkRwYOekOaOX9kQJmaWvnFWkmHspmorbZtc9l1lJOQQ+Abbucato7qTB5NK
a+Cdj/P0Dapjfut1BaU1o0gHAWIz0KhntYqq9KqAtvvHebOaL7zIXOzXuWhk
CjLCHCN61y34AyRkiyV3UoN07xcUyFvnTpo+mptJI7Wjr72HCwLbeHNsb5K9
ow8p7IKXLJUPQuR8A5gE4cgCBW5TK6bD2zQZdKKA8KRPqLEH082sGuOUBSC5
8tXOMu0vkPyDfeA8cmY3uoB3VNhFRCIBnCCghshrGAfXu+DwvUJ3paQIK5C1
IbyxOGBArOeaZQRugUVZqo2Zxumn7dLNfyLwPSXPl+cC04RBGC8r+Fkp/xsi
t9SBgDWgvzR6Qsg8QmQhOYwCudZcHUsb3Kz3cuC6G8r7+h377MsEyfIHni+d
kaETeHbwIBbgEi/x4OEa+q5SoYK1hBynXDxwE8oTUirs7yveuijG8q5Qr5fp
pJL9ndBrOv9uAQ/+pbOzdoOj25Ys/N/c17Vtbq8Ey/F8M3O2HrdurGaWnNt5
19i7UDrTgUOiBzBumJO6uQy2tK2TeYxfotVUpHCpUK26W/q58q5yoQ+f8l8e
J9/2G/40a0M8cU/9fsAERwpwlWumVr8fgdkXYhmd9bwOrhOq/DMEddA5OlxD
jCRw5i+NzJFpoijXRlj2IxxsTpYgPOoU11kCHfeMyVPElkTX1/wUwNCGyGaG
k/ybW36RX9s/9tFbRrHu++fDHv8mFFQdobl5vfYOBK/zbe2LSvixHfkqUDNs
O8ZS7Q9VN6VNHPFgl7qr+2F0N0pS/6mE9yZvJGDcRxzXYoX/SxvLIIah4D7X
3jmu+ij87FBrgU6X2fxl0ejNwYPewAUa/2+xTjP319KQ+Ak5cQhUv0KQk3G5
8dTNbdEOrwPG4cLI2yOZsF/aYXkjXQRGum3u3bphVF6EwiaZfKGqvuZHM8fC
FxweKC6eyiKm2takCXL5ZlrHKDxpgOmp3uhdsqZx+ob3lTx2YE8k4O5WRgXL
ajWbFfWu+h+/a6tjP0rKTBPQJOQI/kBp9OP3oQOF21oXLVg8ItRwGfVk9caK
ar2CtBB8l655KGq52dAdmOigEixzzpijXed1wt3oQDi/Urh1fkMJK/qEOeey
SpwKF7J3j6lSaanJELo22dIeS4EffgjaHbc9Y/bJuw2OdkRh2U8HasZfmpEF
0X+tAFQi/k+mob5vG8FlZPby8X0z1KJ15RO4BoGH7dP1f1T4jKx9qvyWP/ZB
OWa/oM28+sqNBZ2aoRjiCvMOqmdWTZ19TNDYWeeCL7BLJ9zfaw+w9PjzOF/W
wUbcOOxE1fj50K0euBeNSIiys2T/pWnXRtlrbr1DX814XhOlD4T5XSaMo8KU
GjeVtkl1WZ0zxMDv3UBn18n3IUQ1C5N48R1hVpxSpP5ijpt3ALUGGon3WWe6
bjJGNnMJNYVooJEik8nq+PVThVvdyIIRpbVvIfO6tYHElZxW3614mqV/CeCg
i7TX5KPhPbnXyXOVf9HMH3sMbxcdX5B0gkQ8ZUHQYoymvQbrYiocIQl8nVbU
ooqZKxztfAJBVX41Sf0T7hK9URaFibpxD/KCN1y61OIA7l8V88jQKzGqE7Kl
b5nsyGdPCb2V9qea1eM0ezhQv4s9D9a3oubtvmje7Wux/RQ6K5zVdPten9ax
atPVIHzFwM3hRfYUCJLAZwzpLfeJF9w9fiR+o00V5M7PQbDyw8fpwGauvvKP
y5oaEuaE44ykLzzDhNvDG2WuFfwJxRmMRshYhTMI0XIR666WWh+gLqTLHIMC
5x7+hAbkCok0iQ8sNBLrAKuyGTWAnVnvAyVhg3WgIS7xshy2Y8/r7AASVcUz
E5qWp5f1IexZA4Xx2UWebsU9RC0VdNsl7QvQhz/yyM8thdAXadHvowdtml0l
i7FPVpvaE31byS6xVh4VPFGemmzXcB97S8PtASX9One/pAXIUUu23MrHdS41
GUbnX0iiOajK0KCiZdJL1syznBZSNhU/+MP8YhKTHL12pSGIYcfecLMxpecG
eiWTsOnS9ET/kFbw12Ncw0NVby4GmDb4PwoeP/+FnhLCWxhi2ds4UYmAhMPm
Z11jT84qjGUC8wuaU4iEhT6Sx8/OTY5Rv0FtqoUnRoP2QSj1KcHTfsssOHHN
vYCpPxQldwrZH+9B1c5Vth69CRjYu39KNz/tpJ6hZQwwzNKXQ9zifiJwtHve
IkaDwFZrOmcTpwBO1y66wF7Mcr3xHthClp4ZGXezetz8YqVsDKRYM8eMxEic
TfbGicv2o24cF2IiUJIwIos6u5eMOgSGnDC6Xh6us24VHTaUtD98qFQWQNrg
LJhbMZXPp6rxQFs2tyI+EISaxSAEb/OJKFlnykgNuBhu5C/iK8FeabI/xTNE
ip6v2U6XyDmONsf4lahJIiJe4Fxc/epSz+jIFXR48639/Li17d/wE3zYw3BP
19II18Rb/19UBfieV1OykQJwG8mOUSQbcKfJqLWzbjTjMP19r6XF91t/z87i
d0ivsMypBeZ9ChIVJnKgJvKwQfkAztzTQbzk5PfoRfxbdLjSi/wttVvBkBJU
2WVBZmyGeUVYyPf1XMrv/2hC/D4y02Xy8DT0XE6tc84MeLacH162BJR3Jx4K
IN100d5mndNlElf5Hom42Y5Ai+cQQ9mYJE2dtMiXTQKI1b76n8vcRUmJiOEP
avc9omi46GLLKIjaLjiivwLvAIiT8ZauuCT4bGrFaDFFbcn3Sh36GFqYWuif
kF2Lw4G0y457R+ofRAxLUS/scnYCL3V1UUbm5A9FXX3orp1sWCRsIWKKgT1U
TIN18L1HRRJkDqU4DzwM4UEOP8f1sBAWeJGgYGhtE9yGfLA0JMxNXKyySKjy
8aSROCmqQAxt4VKAhVLzoBG26613yHVti/16ODlI7JiRqkks7252QdtSJ6sl
9Rd+jY1SoW4v/yWtXXQdwaTxB0VW+YCwIKRJgTgUD/VOYfpZKFQsQc+47HEG
jLAWrAtzDFI00Q1xrMct30fZHhdfLUnCMXu5IJ7h+33a4wvdRTwkBFmEf6UI
TBEIWKSRfVe/yLcfUBSrsBf/0pHb1mlgfCyNx/V+iFn3DFoqMSTkwQTRO3zD
FIKdh5ytVLqA2p1tcQD5ObFR6/jC2HoB8CYpS6WxCCyGri/gnIgOqpHx/peh
4v1jBTRiWm2UnG4tW74k/byckqov/MYkuR6C5MchZlHfQ4aRmAz1jcgUyQZa
eJoAjhlahvk1BzusthRg8WDNghOKmOe4IpK7Shl/LjqecV17KljqTTg3lYcV
RddI2s5w5JT+z2u2doYbo2bkRbeK35qFWqi/7B6fMhqjOdm5FOHqAq4PeZWV
pd4jC7MpfwyYTYuV2I/yZSAi0bI6v3xylA6QhNz9SPj/7lUI30p+nTNqHkHr
diZYn1R9rO1VrRo0rnXG31MXHkm2xb8Qg1cR3zPTHzg8NtuOQA7OyEaUXfGo
TMKqasSkfsBgAb3yreEPjx2L60c+gUSsr6vFaFkCTD1wg+hh+TywZSuPw38P
xZQc/me71G0PrYXXBdoADVw4Qi1QziSaWljbaUHV+3GYyriF2UszWUDAo4UZ
8Q6HLjOpI+oOcZYS5DnMiL7d02jDVA2DeGDvR0Z1vIdVtrtEBrDW8hIrnpOc
vITunQR4F8DB6li/XgvnPIkszY4QxgcjMyTqR1A8eAsccctSV7/zG1nK3dYQ
h/O21Z7ZUI9rEsGXmZT1r3YTANRsrglsRUsPGcHtRG2QGmdrUYcXi1NPKJDj
sgFBzBJ42er6BTJGg15/cCllZClCqPjpsQt2RQhYHUmqwLdE9rhCbF7tqL0m
3xrxac5XLhBfQwystTmywd1HmLzGl2yTeWzc2z5aZdpffWbSV284sNUoOYXm
kpqtP9K9566Hy/8+kwRM/iq56z1pBtdQmTCCwzZ4G2hCT/B7OD8U4rCQGwCk
kuUu0X/oT0JjL2Ux8SwoCbtTEnB4pko8jodWsgxnoN9osLZ9WXDPLYtbK/V0
5hy+3Uz2B8Fqv93KamCh47XkA+Oyo66wtfj4PJLlXsGxV4Ze/LgoKVXDwC68
p7rCFlDa2Tjyi/ZfQheUabyT5ry74lLEeG2KTQRjN9BH8LiHxb7jpVaCVguJ
OS7TxyephgnFSrbiP2x2hgvYjuP3kXUXLXIJZzbDl8p/untMWAFj3vUpOD1I
Nq3dOD8PlOn59VOCdWFpJ4WbHMHW+UjX9oO2toSmCmEfSGyu8Elxc0nNudVx
G/lIBCyxN9cfJ3HsO3nHp8LfGjuPsxVwf7DVGVR2kkxHTrVw/75D5teHnNQf
51XG0ZZaqR5rSmUvuGpY53/u5fRG6DjPGzemNJacBlDmGo0Zb90GRlSelXPS
+cAHA9HN3iJREDIihDPb/5EgQoa3IVEjese5IJDPjFP63OtABp3XJKQ66M0G
aQ35/7lHFviybrIxI9fZUYliKn3ZXRLFJGWn3lRjoU51h20o0r2SMS4N3NUC
7r4rmzTxdQisGusMfmbtF7AgbBvYg66oR37GyB9tpYZYntdzxnD3gsyxLIyS
NxYqRc+kh+xG23rf4BHTx68r1awmSnY74jqhqWfEpc7yuwjiYJuoS20S0mdm
7HVrFfu/0jP58awONmq0Vr9z4ONX9WusHKFW2ee3Fsm/jVxT4ikj5u0Tf3OD
yycRFT+mke7oyb6sfPXfRvSgecN2r61HKXtpeKwX2WVDimMn6ZmulM2TWhbx
PO2ijaY9fkaH64mz0Kz50mGPHvFrKtAHppq7pX4C2oW6tqeLf9km4qdW7U9I
f7yJZdAiBVk866Xi75jRatpsJASxOdM+MF5pVCFNLuImhlArv7KEegrTa3pD
sE+teO0EPiE+YMKZF3nt7Y737TiUaIpaqNZownuDZdTJvtfW/AwPbEGZNDmG
jKcfcedTx0H2R0EF/RfCNEk0hxXIPUn5BSeeKK4CTV/XCOydNT5v83rqZG7h
QNO2+hKqjUVDsdwzhYoT4d7KNLxClc9pVf/k9+c0X2NYbKictdOev9skO0Zy
2x/CLqAWy1s2DY6B2Fb8ydhwVi2wokwDxsa6dQSWgLOscrT1+Ng/BBbvCJaA
c4irZBbsyov5S/q7/QtiVMdMLpqyNumpYAte5oKU06hdcgRj8STS/Eb79y8Z
E/ImykEdlfz2Q7hIHyQPsuaBYGc7giFMG96bUQa42pqmCs4gd347cbyV+Tkt
wGmHB/8D23+lzUtTSmMRLrOERXLaPy13LwgVhUhib1FRom1hgg/OFLsC6MYl
VIGlXc2v72hzS3eRdmKZeyeQx7PML3/2koCrncvTsp57tt7G0uzurhUBAyTE
B31rDYh4VFkKPzP3OLqJsOhtBkadG++eL+T/x78fBWW+vcrKaVHDn+8Qh8eL
LRorxyiYyyjOA//PgK5YytemxKq843S4Q8JkwB9urbJXEOQGceR0kXkJyNOg
eLq6IsMuUPyDBgR/yl5XBd2pQ0qs2EJsboRrcqDiuAqBFXLsXwQJNgyxho+w
u0gAsa03bl21TIgoPKZxFy28N4U6QMQFjuozsz7TDCUzUvTUkFFTF/M8gmMb
nACVH5IoiSSuqmQ8pU9aXJ+wAdE5mClLgMN4VVSopyyTRcTG6MzTPq10g5A4
ALyuAlH4U9ko3Meys6BRYoNZQH0HI3BK5hdTCIrbW01GeXBu3R93NPdUVFYb
0lgGZrjjLDDNpNKA9QTv0/BScJ4eqVbRB7rpZegugJA4RM5SuTSC3n/0dTcZ
PwIX8M7xfwfuAT3P4a3SVeapKMkwwAe3KCc/AGdmbUCk5Vw2SNp6wRHNcfjC
aBOez8ifobMthP0T4bNVQyFK7Ex//2JAV4vch/a701CpYz2MV/sqzt5cUvOq
RLl3iTWCS0Xbnasd7KhvkXcpB7CpUjyReNHSsF2x0rS9xh/ZiAAtyYfP98qR
0SFFxgXZAa/c/o3RfhcgCJ3YDzKQl6/haXC8AoDSaMBYH8FthtD8Iyeo8u84
AFRtjF2PQ1PTWMS5YnY7nMMbYCzv0VXENCkavkGATXWGG97iP0o90sz6GOi+
sjYhD5vETBioZ03M6kBccs9V9KGztwF53eupOeAnmuWxXXTvc/wZCuA1pc/+
ODM2WrBibtb8QMdjFGWtjney7jidaUzYYO3/xfJoC19DVCNvVQwNGsz1Qap+
OwMHqBrgBiyjJLOwJSeS+JSPPKow+KgvKm2W94IGIpKjr+Hv5NlDIjc3YrNs
tFP/eAx9/DOG/LxE/ZwwPvnbaN7uvp/14cqLsi5kAIfgaKSq69Bycne0/hOX
flVBA81AIeGUoFx5ZUSqBG/99vfxtWBBx4BkYRsbpJO3n1lVuyH0Jpg23QkM
+1ucMyV4q7b6xY9TeUFekczul1cSVwj80054saU//Yxxwdk8lm22GWXgwWoB
O8HtlpbIqm79zVfJGTbskW19vTgKZq8x9x9haMAauHakzK4KxuxA9rZelZ1t
Te5oEAhpn452UCtggdSkpAuJxlSBfOjvIsZ3g+2K10/9GIxH+irSgAw2sozb
Us2Gey2eSC9a/r5XmojuJV+Z5Jc0l1hnHGI881H1RiaYRNfnX6g+30Z9j2XF
pTHu4GoWXObR1sOXZzmNSYBGLryUA7/H5meYF2H86OFCIKKUtw9Co3nBAs2C
Y0o6MKhrcPEtRwaGHtxeWaDvLtZ4fnvOsFmgZnEC6Wp1IxwU9fTI6L4RDyj5
BYVkQ6Fjc/3Dn0HOOorjLTJMCyIj6t2PM727+kqA7jWZCiPKA9t94vFCxn/R
//X3uQioy3Igi2cdFbD9gKZ8oE5r9llvJifOyIzpGI2GLOqn/FRmsfJyA2ZD
spPboJQ5n61osmqotZON9f9eB4GwetrZo5oSEqNkrNO4iwaFN7aOsMYAIaAE
WaG+L3khje8aYPqGJY00sbbU0NkEae30U3IV7kyHzTJE5kL+rK6KAq/BEQmK
rThsbCapoGhVX0IBVJFJnMIuV6QxKKAKPDznh7qoN0nwTPx0eUWFNiufN5TF
iXsq6jvwZSl5Yi452j9z+oSYk7o4vf4eplpXASERC38GE0JA+3tJVtDTCF/F
lnS7LyxzdTmUijWQtDwQnhw2zp6D2bte8nbX1HgaXf2j9LUsno0BJcqDEaBh
XCKzIkAY2tqBLXQ38rTMnWcWt0+qYo7n8MSm8Sy+Foa3idsBCXjjcHJTGupZ
rf/DpSalq5DrDgy+hO4ryeTWjMNxTfGtNrAeYObTZhC0rhqJAptLLf4Obv3C
jC+Mo10oxBm+BkXbExjOdzj8QiFQ8Dlei0g6x3nDINVscKxc7/fRBTNfpLLA
lw5UaBCgNwBlK1RwNeKyLUl1m4HEusCyBwZXYt7XaN1PD6o99c0vU+UJWZuC
tAdAOmyQn7Ygctjrd4rZ39M+paDl45hbJDu4sxXka2UmHdsNrbqivYVtlwJ0
ye1S4X3uA9IBdhPKrK6bsp8HJJc4hxUmJcqooC03a11b71/MoLRH0sycLW02
P24Mz3yh5gdfVOXwT8u4Meqt5gONgs5l1pCfSBS6WcluWL+Ak9ExLoI0luNM
PN2zmhZ1fhTC5UAwbuXoN6PNpyYCuKvOTLCZB4B9wFnMDi610QXG4unJz+fW
6+kM8V+j7fonIUgkSrCXPX86xGTZNXyr/ijeAU2KTp33Bdffd8xqnZUVfdnJ
DPpVwX2vyqnP8MtCft9SAwZIMULQGSeQSTKc/LNOJwi9mUc2LlbRdnBOvwXr
oVpE1gd0Gqx+0H1HI7gz6H5i/wgH9JyQ3Kcwx0VMcfCearUTbVu2+7eIsga0
pu1p919ccFmUCOWi6LCUQuM/dqJUkrrF8Ej2TEikGdzLmHi4L9Ss34kQUyFA
nL8yFJKG2aJJZcsTL35mPe7SqRZNXzMRErlM+8mXPyJk+viEEaZpZLvwJTWt
9FJkB+VcCW3oypxhZtPfjzGohwnaOOicJLW+FyXRkPjkPhHmgFDYGBCrjLsv
PHgT/hD9W9588IxhDAChmoDGeOketfiDJCVvl2lsln+bgikXPuIzozn154FT
WIICS+kjDq5VRJFRKewmk9LDBGWESLH3PZIbuANjbcyAJaz/sWrBhyP3BerP
+vatoh4emRYYYfmRgn8FC5sNeog/NGQbPwByZZc5uOjyZuwyaNRQdrF1NLZU
JsL6Za7VxL7qzRhJzIXUTaHd/tJmABSxQmdbBX/vyXyGVO78vlCuAGM7bGmM
2XC70Xy6+fu0SFONH91aIK/j8gjzDKMPNF5HYHxQ9ac41hLWP+DuJblTdGYr
G+CJ8y8D16CibiwbgqcZTUee0Blcz+YR0j0yHRo6I69a0LNKEN28pdNu2ezZ
0VejzcJDKkDEKVcYijFJxTgVv7+oNgOjoOLp5WvA1qvsib2wvkQQQ7YozEiC
t5KBRaj9xspqFrG8NX/r2cjOolA+q1AlXNmb2uC+LaoONMBzpsGOGCpVPJCu
YLnP8fFX5CX9rB3GYa4kW/ZAssx1AfDpBRR3wfMkV7wWsyo0FHnbzKNMLAII
kbgDzrIpRpNzvwXREEVgFE0mZdkYEXbGfqsC5LA105GNVumhH1eF8/LQkZJs
VBzxSw1G7w8ct+faZPPN22hjR5BXaHs7Cvsn2YZEoib1L2LTFjtME/aFYNpR
93ouTZzHSXZNR1Tfsc62o6XZ6ucrgSj/MeSSoSGmufIDzq3MenaHx3MG5GOC
zLtUX3MwGLQh4RLO+QchDtstw0mhTexmivRsSze1hpwuL+fw3IZspXfTMKES
Cu5qSkAbn5wnRaJYVONp/F46mEealhpZ84WlbDOepl9MyNTQqWalTGPefA12
L/S7lKIQPTmWP3MRsGZOlVPFIGcWizWm6yYxhJ+O2U/Ghk3u06e5QIOYmjaQ
E57/fCXG5lGJHrFnfVjLQ+o5QSgcj1GDUNlTUzOPGGJfzFalO3WZGWzVwjW3
yVNRhxe/fGEl6WnQ87K68KJ3ktZOH/JtSj8DyvilKYvfuOfbG3zUNbZ803Pg
FSEmStHQDOMJZAc1QyxrNDk8Xl0JLVQnSrqqrVks8iXCfS6unhrCptVrngUe
ZUNR4ttlIAM+yh8JAlBLoffZmrYIdbkRV9ej8A7U7c67Tw7rYV7k7BmwjJer
xr9XoYtzqYeLJLLnggpWe5Ok6sQRmu29jZvBMMVV8qbn8TC076bfOXwcpSff
DlTziiM0GL6erPq5+cYr5hDTcGA93sBO8IarCz+k/fmKZSV40/v9Kz1x5UuN
mHwGpLpdPurw2FcxJ/cH2RUhWzk5ydbZuQTVRyIU+xLSZb0zxw9vnLJXEayE
Iezs6UIawAhBaiaNTf1ediA8kuHrQs664OZRC/ZkpSPMyMmJ2koegWVgt3cL
5c/wM/xuISkItQNbf7uqzavUCObayXickjoSY1FizTq3l/BEruIdDzU8fV0A
A1G1dxoGnnOtrwNxTJTkTmsWb7mhFAFuXC6vDjVZ+pd07HRq8jlpj649eHvp
2yKyRC3BWRB/a/Du7yPan6jIWzfFQ36RtvF9Dtvw+iJBYWNpAKn5Y+uvCyEj
y+zEFFqLrYM4xEo87UJdiIlu91x7rHY1ikVwGS6yCxqtsa0ghoA8hmD3xCR+
OS1UdPQhCqGJ4re05+9/Jc2JbeDleFyF6Bry14dkAst2YptDKUa4MAJd470T
wMfsc3p+2kweHJQIPnhMRbRf+N1VbVa8pUxRmhhOKgFAib3p1n207jZW6rb+
9yIaGkIMp/Kpk4Z06QMby5JiONhT3+ZwG9wBtFD2XQCeWD1vYWsDxreLON6I
IZhU/2EdKW6sFa6AcdDbe1e/cuRb7oDt576tx+lbh6V+5ZpGQHkb2Rd+71JI
L8DlcNZgV8CW2KQqrcWlFlXFwRM0z8i77N7NNgFnzto80WY7iEoukSfihtw7
bXej5DJUPnIZppr5vzdbJdNA39WLnXxDUINJCXaL5Rifp4qXRjYf0S00ix79
4TAXp1nuaI5j+Q92d+EuTXj7vIDQcFzspL1YtJ8tSj5/teaCR6n9ntOwckKb
GEAKx0OmNSQoTfIRnDEDiwTox2v4QAdP29L1A4dt+LpIc8g92Q7dogjuJ+64
Z6pQI0jDYGJiATAmNOPlV8rWI34CMZ9cLz+dgh9e8vyaavuf70U6JSuM0niM
x7muM2DI7JIxO00/q+9PpSUf1pTT+qmqw6+pre5I04wv9OZkh/2xemeY5VzO
jiIwpaE16Gb1cEqP4ermf0GoRxBul9XMLv76x3wfucW3II4svp1GM4M1UEap
5heFP/Wyd1UDLl1SNLfvzqxPJhzvD1gyrT2dKrat6xLMbtBSMyQqrEkJorfv
6TfO/n+5P2B1VysOzj99ML2UudpQHb+djfj5vQSSMsjKHP8C4QunuJqQNx+I
SoKt8Zod8vFVJfAIC1LbliIyYXmBymVYLKO2Y8/VmMS3H8pTq7tYzuJCIgpX
nJpkrTpcoPNzeU/7fi2JebVCSYYUjj1bMI6Cpaina2v3aiYTDtiIqVQyzw5D
c6UBGskRTqijI6GL+XQjLsPJO7hih6ccQ9j44NLsZh6OVmO5oUrNJGKb5NhR
UjeQrRI6UWg5RldR2It/MXwegYsvYUzWY4OBPzeZ/nXOoXt/B0Me8ulRlNrg
7TquoAjFN5WTN4w3FxDm0x7DnIiUJbIWs3TqGz/MOPpXUXhlyThXSle5oBD6
XQJhpI3794GElDzuwD/RRUqwtvElpsOGvzt+peKTrZxhpUxFqisVQ8jxi0zT
tXp8YzLfsv6jPcAbwoEC/835zMbWoTbk3f7sv5Grlkewn/P2SJ32+AXREx6i
eLR9rPH4f8GSal+urIQhIvbFoIwTlM7Fnv2P/50sYVPa2iVxNGqND0ztRL4E
KVXbA/7En8W21DVTuzZ3Hk/cSWzZMXeXtub1hHhB18wUE6oa1FElLUZ3fGnR
PhQ3PxAZNqXb1eaWitYZH8JmtTN4/muG0M0d7yK4E5shHdE2K1kld5MoY412
DkkYwelfuqMWIDzXxQ4egFl6nEogJZZmeDp+sW3lVW/GWG6+LiIhT30k/nQO
2LQ23jNem6s0CKXo8fEFt4fN4r2JztjzqhYL9uQpNZX2c9C4lksFNamHPfHT
TA2W4c2vZE7YCCsVKv9rOqz5IZO6NuGebbB1P0R/XQRxlq3rX/vGVuUzOGPo
vvdbrRubQPn7hl5osfTtPqrsU21M7KDmenWJ8nFXmG/FC8inMY0hLCKt46tW
KNLNnx2QMRVvkLiRfPzOdme8D0RAkGx9sgVwFKWPqDdBhYsMAFWQ+OWR52jF
0K2p8tIptrZh/tFlvJ/efHMB6AsC5FFv5MjqBdPUQQwdz4GXTByCfcVB9eoN
cYh5Jl8v4vjbJAtN+tFw6U1TQmdSVgwGcoBMQsdG+TOMSoYYW/Bkrg8eFdJx
MeI0x7WOPQrq4/SnxA1DD0fl582uT/2Mn5bHz7hlLOyeHZsXXw7NkyO8CoQF
rkiPQ1aPjAru1IZnJVQXHPLs4iYDUwzSfRDPoLIwTc21G7KkO5f0O9zOu7Ns
UeC8toLUIjH/+rJvEB1EbKYICkchF/0twtlpdnkemTYqoHvod8c7Q83HIR7B
RsaG775RUfQDUYXKCHrgIh53PCowCOf4ICYi+ivLFEtJ33C36YT1s5qLaqxe
FIEDx+4HDV802bto4wCRi9MseSh22uDGVKA28rYVMlZzbdHRngx1aeFIytZ8
87Brg4Cqhfo/O+BZjTAj+3jUPT3nlHGxUlUzIeXP3BZH2qmc3pG7Uu3PG4gW
/BVOUTxOMSvwjiX0ahVhpeLOUPz5RlniQE3V2PVwIxtYj9HEoS8y4P7Tmbtg
ZooJ/iJ+0cys5P+fGCZu748xRZ+eIm1W9Mn6s0bgO7GnUtQAmHBD964D9TMz
AzPMC4z9vUCdZGuZMdszu0Grmc9ipfLNfPdC4M0nDbxGlpRCpsDYNy5biZbL
cWJHzejLiVi/48+Igow/L9Qly7hQu5Kznu4jMOwcrij6983GD4kGyyaxMMaM
63kgxdeUzvYcgRY7Fpfp7E5W6aGmGqbuIMUvEwpY3S9PHF6Z/K3nYMdMUjsl
/UmBNPnmxhPL+VODQ31jmu40B8VY4fyLZSZaBP9+wA/ON29DqyxLuBqS7L5K
pwy0t0OoFvOzL0VmgGNpn9a4RsxRalXnaA/1mbkHDrC/v7obV0d/yDVQPAF7
B6vRxWoCZQUbf6H9Gc5Q5gBljui8rXxWKc/IdFERHboHrr7G9718aG3dS0bu
yGQNP+r2hrXUXk2wh2S0dApBeLfHGFCHd+0Y14BigUKznvxZFbVlTJiD6ahL
3tDm4oLIhX9LFAlqtI3VpxkwQULF7J+XcsFQr8mjlKP3e0SJGSgUmcWydjb+
nayAXc7kWBL7ANdWmFb70+BAhJvG3aRq4F6IvSB2mNkvsUYbtg9t/iCT3W24
W2s3IzTgyIayBuvybDDFd4omaSNnTWLg6hvDDDuSblwtiTH5UM9Tf+lzoRRW
zvRrc2hdUsMiFAZTEsX5abAMcQnxr8NliaoyB0nkRRAliVmO0+tmuzwDZ6tu
zMcZ4Xv5MHljGDaGDtVbleer7/uIvzgkspGyWMqg8/JEBmCxso7k+G4cK4t7
ScpqP00QAL+SIE338gt3eKXLK+ugQR6i06lhgt8i9bVprVNCYXmbuRx6jII3
iLkh19G4ySXGD0yVJXNer6eA9aAqt6kpN0lbzW7ieb6DqrckgXek+iXkjaCh
8uGOHABYMUR8FkjFWZk9U8+Y7VxljuntTF35zlsEw8HlqHk/Ggp+xJd7bkv2
X0Ww+AjOMvTznKOJCAi+kNyEopY0S5SetqdIqcduihaFgYZAl0o5lRuKbusf
xufkgvzY7Uc8krhOXCGXX4mtYGcM7pEpiaaRonYi5vhbBb1Cj67wIUEYC2NC
FcgUu2WwlH1wQ2REGb98bliQP/q3riNDxqgacoA1pycgVis4sVrv5fDlQNVh
u9RtVaWEfuB8DhLtdUJ6Bs677njeUQlIcfH6y6akhuC5zm75+sSJ9bStgP1v
g5nPKaRY5+U96qRBg97SX3BCARxsStvIZIzKlZiPfo+yz4GaE6by9Q0pkc0Y
gH7q9aPglnhwJisYJaYNYznLt6FgBRVjkAHzG7uM/mpfOmEvzONarATECn9n
Z8lYTdn/btD/6YiuIm33EqFWSKz/Q/OXQGJPoEeW5VjS6NO9NnWneRu6k9RC
qQBDBfA2qI9ly6aikTKQCtBa5zfRmTYft7xQgXUF/nDLqTUpwtBk4TAwhsfL
bkQKN53C1PW4d7ZPceGTfZUOgiOHTNJz1+wpHlxOOyvmIylwUwi6B/jjQtWw
HmW0JxSm5DaHNM3sL4hbtvbHNnsZYpmO0jpx71y0djut/ERdgPs2pz7yyFM6
HbJxsGTEalKges7oRMc8bgySTdvKBe52f+rkLODs4cQBnqr9FL5+gEfBttcN
FLW9D/MruVOrRP8DM2krhGVfZRCWtb2VgC7QRJh0CemcrRF06IMTtkj6v1Wj
Yr1ZFPpiHRtL3MM72j98KBGi0mcjoy5iWvMvlvLJhStdlaXKzxs5pyUwB3bZ
omB7Tl2h6EK3w4x0I1819PfV2RIdimIGbXvzsRwhkaPXs2/XfdGDIJNbKtQ6
cWzND4JolkoOnp/m6lqQtypC3le+v9g/3sYAJ5JLl3nIuIkJKrc//ICQweR1
8I89k9ExdZeL2ogj7xxsVoNIOSpJuKmBajfp/pvtERCNc6OomNzT9bLPxcYZ
QhgH1543k8ecH2ONMygyvzbEi/yc9CeqgDKOjQdTaayG6k2vWdXhBM7DVQ9+
oSvYDZQwBq/GJUxvWueHk45iWt+UmwcTlZ4zsngUIiQ8khfJirjzqv3hI/re
iGxVIIOi1N39PLU3ozUXddjZAJFJj75mPiJruyEjzRK6DKLSPnMrtcBBRCWP
DgGNMa8gryZHCl/IekVNQ38jldmftusGmUQDC3mdRij6tPdwDTPQR8wH4h2n
T5ASea9y7oTsGYZwO9XzNbUegSl5DRobRPbJieTyl/736/7vFB7I4n5/ur6C
2BniASGHS4Ob7+6DXidXlDzxQzG6DK7mzQvwjLsOXK/MTmTwzqEuQqNKR2xB
skASESnnLBoPvd7BnnfUvgdzNDPw2cjPOq54/fArH29Dk+2nOgjKGhrtJkhq
Hd1283tQ5rNBNr57xFajyduxbDtMcMZPJ6maMV6zAOG9cIr6cy30upqH8HtN
fnMlAhJDdzZ/2izT3zsxCWlRTjHVH5150hAbzgcMVwK8x2oOsx5ZEqh7+AYg
pOhxFPJHzHEdlZPUEyf2hkAud0uo9XpIgm6lf5uF0MGZsYPzwySjJe2gltxs
IRpFsqLC53gdkImmbT0EpmqysuY5IneCCjgK5E3rs/0wzysR4YiBejIja2We
HRvSZjlW9QKEcbBYJOZXp2nydm8Po7nzSS+/9Pma0W8Xrbp2w0ePuj5/j/Tn
9fO5HBfJoC81eyNl9N8P1fmHuNxYrIrHV97epmBU0yZRtcVIVHbB2Wq0cMTJ
JjaQkLjnwkjodwRp2VVaQkyR7CFabnRrRKwtbGzJ/F0HAs50dP+k0HOJWCGs
aDx8IBI4zFESW3DCRuuR5FRj4lcdPoKNcurt8tDgdVJMTMbfh94rlXgDV3e/
hb3Nc/Awc2VSiqfatv6PzuYIjHGguJVYFB/Me7DU1gfqezMnDX8jqWOQGqLA
fdUxKjNtg5vRyfqnXyZv2o/TvpDq8x8eviMLLj99sUs4La/PSvXSnMgQF99G
H4HnPTdnFVUIsou7d26dY6ynFOM/S4OQ82Px3LIx9qu8HKL+PK6X7i1OgiZu
LnWsyX913iV9NOSXjhXfTLANADfljmoCJNzI6tW2klCW0/sjtFuF4uwgszvA
AL73kYOGoLk5NQDBSQ5NwaO84TwrVIyIc6wCEo06xhYIcwXVBjVV3bDfN8v6
C+odZgOyrPk2J+i708fka4Z/dT1kcHooOWWHji0PHlqSCFbZgmMs6czKwan1
Dse+0MElZwSDGfmQ3KXT+PM140uNvZNWhzHTK+MNRe0nykqqRE+oVA8zIhnM
T0heElUd4cvEDXIWRbu0IC5epvwbXRIdSBdEoW6ZBNtqvviTd+Wi7pf3BBKE
oXKT7VA+mnNwXe+oLN1pOXsyzWDjHB0LtX2/jzMVMINpHTH5hsdO157xpnBr
ApudVBZ+eZhO80YU/LXgXVIJd9VMV1iIt+kdpXGZPrykxFnY1E5o/aH5FelM
W/q44e1sXKbXTNJKnPdp0dCuULEjmOSwXfGoWzAvGJ0/hDAfGqHaUg1kZbSg
88YxPX4MB2nCIUxrrE8dj1CPkMAxtsmPAZNwXauhoKfAOeyxhUErIhgdqM/U
6blAWGqx5kje27TSm0x0prAsOr6yKTstsf0bbXW652MfKgk4mMVMu9osaM++
TXvruexg9eM1fhONFWK1b49exLbkwnaJajtpjA+DsLRy8NaalrVaFz/kFriE
d7e/PjpySgPhxWxtutCn6ByTI3SgA8svo8HgYR0fb8KwHQlVRClRA2MvSNWB
zuD/2z4ie+C9CmHdHjmASEGXFdzi7FqFkVozkLrkO6jyM8EfmDzm5sGrpdtA
8lk3hY+OMKU1cN4gvbRK31Fa/FNgTlT2vi25vWQoMGfgyD73A+BuM/w582mq
1XYmFXnTTHz3sY5qo88Tb8jm62hqhwb79Lhi0HNsW0jePVIxtFs2XfNSjHz+
5xS8pGro9A9i7P/nq+IxZ1HfqWZDb8oNUwsMd9Jdj7k7j9HY0u52uvcKX+Vn
inbXhVdSvC3s98ksrFb8EVY4M6gc0SUvY8B+BbmbBd4icHFXLR6gpUUupIoW
WUU3Dsc+zc3fQXUxKuj/MhyxTaLMpUujIEpbx3GJbgXzv9SU+n4lter9YuCL
RcBeTe5VBUV9w0ZHrWKrF62MsNVaZ1t1ylFLRfnZEugPxwKqIZvB2n7rTfwh
7vmMYbyb3n78UmHJa/QfzrgRhoSCrsYUx+X1TuXs3prpvqSKgniJDRACGvSE
rXEffeipoTZtWqRrwucWWMntplzdFDkvcBDyWKyN/vbAQX2obCn+Km6XLGzC
1N86lF4UyaPEfEGzBvkDtTKa896SkH027L+LzK/xRtFkEFiopBn9TXYkxB6w
7KUkYzIciDdnQWQqUZ1DovcqDyKwufBfw2z1OjJgPHR2JXedqp4UNBCsJn7J
z6iDZ7CbWHCarsuCzSYblT4014XgjJgsRH7thkgIkARAaa7t1BK/imNJoylV
lWswG/79Ea0tS3Lki+9U9OBNvmE5xPfFr8JDLZCxdpZolBRqaTbF2a2FMs2v
SWOOTIZ0kMw7AMqzrbuM7ccO1PSwG6hhAiAL4ZS85qs1ihk3qtQkDXd+smX3
8aXc5FwE2SKTHOn1c7DAZDDCnL+hJX2SyItLjVz9o4VV/m/EmtE2jkRMlLyS
QljsykCnA1xsPTZM4Dobm4Q0Kn9lmbHUL8QHmrH0VFowlPXuuHVZkSQkIzRW
ddIPCuT4e0gG81N8aWANGY6PZz7ymI1v6hXYOOYeekaGV0wPs/GnN9qYhTwL
i/8BV/+ISqHlq0qV4VCJSbniHdLx0yVUqkvEq7Veesz+VOgdT6VDyzLp7auH
uOEyXdVVrX6wGbYLx2EiwQEBfQPl0iQ7Zcr0br3FfhsbBdboMzC40zgQXEgQ
0I4lZudRs17cG5g/me2j8HLi0oOO8ciyoBW2tMSqEc+hCuPFYW0RgVCuF8CP
KqkHj7QvDpBJlYz4oWZM5s/K2fsjDrCNMvX2jAeuayHQHHY3JUC+k3UJcM67
AG+LYL0I/TTjX7Wl1yM5IRkNUuHtrMkcvdGSZBEzc9tVtVnWzYHxywbrHVnp
8KRliCmcK7pNyt0e/oX0cpAlvNElxEQkR71xXv7qOBrAQ50uSLU2Lzeqa7Oj
1SPPuShJcQY8qButFG4VL5f89DaPccdnzrERcSgXckIITDhlWN/VzNuM/J6f
M2gTf4u90fZYXJoIBWRHPdzjH81SQintxP/B3szIoRum6oIOtuUJI+Nw5gIC
Y0GKL5zGPksr0xMUl8zySxZO7avpCoFBFk/nomI1w3bJ4gH5IwK0M82nBZOz
yOU+yoYQndzb/RV7lDYYQu1mxf3hCfUDEaBjn8OVpaEq16QAnKt2l06apCSm
BT90QggQiehtjhWXedKrpPjwI9d5xPvx4QmOmdeLA+fkscnEJaJ1GS+bcgBX
bFrxMDEzd+RO4YBDygtpq7KPcpR92sS7zxHCr7Hz6HtDVjSimJhvq8yudWmy
gS3MDQ75nbKiqa1/JSrH9px18iAUKEDE+Ur9Qf19xyHlDO9TBR3YzY11KfJn
Pu2z6aYC9weNxIXArItelywCy4IBb8xXo6D3XQ/CYxhEemfiRlFp42NqwbYH
HUaLnOLMCyA+zmAghN23vKGDsEHJ/6co+nA4Glbj08IOOdCLXwnfPjdJ1jla
968kIQ//fFwl9UGHBs4WLmf7g01RxKbsUp4P9AfRFpEoG70J5SE8yK7CylxD
ab/80LTi99UkDuBaGjlk4eWfSoL4pwue0Q1SiaDPwI5G27DI3O44vP4NUTND
mOVJ5WQ5P1ZjSsqL16wneWj0jTpqku+lPpbYKnj2QeoTA+fxg8Z1sHeG3VkK
Bl89mVh6JAZND/mOspziPes72nIUYM92OihR+U5nsl2zTYNhqagPfboDVEl0
76Ts2lTa/5cNWvzLPAcoxVHXOX94yhSDvSLvU6wAyhZ9JWUY0L3mVE4Al4XR
M3QiqK6TL+vNiOJ1Mr5rkIwywJ6M0NOUsZ1stEWf9A7JSnWSDuyws28Jm3Wy
CY4ml7O8Ca+pOjBj5bydAjyHhZDiDP1sCTfBHws9w2Lr+WE2YykD/5WZTSTa
drTLnqkoTzmchgRI2IbzcaUX50xfMOt+eQ9D18T7otKU924dkSv6jnY3BhKr
jjxBo8kZD2w7eiAD9usrNaZf93YmP7L6lWqB4/DbV3Pw6aIymTDu5ZjoxwlE
y+ERxknwAbar8EooNk8B7ZHgwWAMLsDrX5SvWOV6vAqEU5mm9KuyF4PE6YZC
9VdLHy7zjcRlb4hV5ejZrDFuhYLfrHCp55wX0gu9udMXWBsTXVhqIwgG+djW
/6slpRnQ3KJhv+4A5dVCyrGMHYjEOV95DMUVSATPJuG+bPH3x3STHdHa4sGJ
1IrRqcpymQUQQXdRspkIxlResD6+EwxAthNDfo1FGufqACjbhNnBhj+y6cEp
ZV84XcOLZIRdHl7B1Bk8MuRCljSOC5Tn4KNbyjQuacfFS1xh7gVEBsF+dLqe
HI8DTx+fsQuuKWq05Y3iGCIueeTU/5g/Nk96zdVoo6kLxUOAMhZfmQjucXSm
9rGzlnPqHZJU/76o3YS58wVTlXj6j/8ViVMksx2mvl5yjMgjKcCKsse6LgKB
lVrsMqGtBs71xng20WzYZFV19+/ohpyMgU/hMpbiolBA6JsXxYoLdACTRvpk
R+IT3ij0kGE3Pn1HYIUsFG+Rb/AOPKMSV4Sg+fIlVIhx9VKWq1lKVPXd2ZTo
nxigiswsQ1kWil9gZJ1u4MDeP2EHrnNsw5J/P0q62Ov+9B7pzRnua5qybD07
xjhuwsEYw3fr+YfygKEDQq00lwmxrUwCwlt1BdUiI0PTPojlrnkTkiRyhTSZ
h3/5cf3uhZeE32HbZLSris08luFcT8b8Jk7Gn8vFYemA9VkGgkGU8aod2ys0
hHnCStWnXbLx5aGkp7xp47Eb07DvY29r5H5qy6TnHpV0ojBvUPwqccNwYXPp
8orukfpPCwJFaxuaQq9xhumhKUifNnzDxbDthUqZJ8TEMVA9IaXMmzsiVFuU
op43x+8L23vd9eHt7OVFJkGOj6pcGPXLDMqH0GWhcqamgNbMLbkdE8OIjwKe
+C2uD3r/pGwXXWg3+VMrUpQ6X10kpfmdaeMwi/jY/eniJa+cf1JSE72dGD0f
tc9hWAuZJmVEgupg95dTIesqlOyOvuCocQRmIJDJlm1RHwtLR5CS/hr5geHy
uOQS/T8tH6zmKHsVA8Vhh98yau+CZBFSBueU7XofTcwkVXNBl4SUDrP91nw3
5xtOTabVcfwyIrYJzT7kli813M0G1Wyyx9MkT7u4PCJKHbWuA9ZxDllv/UD1
xQXC2/4uPkcR7BB01OLecne0WQxu42jO6XRDmKiz9BEXfuvlhPu+p5oblCWH
WzOcQUZoS/yOXFvuPTynwp2l6aKeNL8JieWTW5rFZgChL4YeqExRFtjZaA30
Nae31Tio6dZNKB30B8xDvaMTA9CvytUaXYWIq3f0j00rHliDnZA4Vgr3vcvW
JWykM/MN4BxKLhgsirGNeyazs/T2W9CtvLlO+5MZnxW3uanikz59eiJdl8bJ
VbVA4keLUVeN0m3N8SiYFws30OoZyxPwrUHvoCOs4x6ss2690sjPk+n/DQ0u
b/U6nqWSeuBny3oaNyV1Pz7fST5BsD89mhz/yKfB7/so942PYatxXK6fcSn7
35UeRgQwsL48lQaZIpXlyeckac9tfNU9ZH7m1xPmuMBcohNVU1f2hC8lJYAs
NMIt44B3q2ixFumX826axIMAQURsKvZCJlBtzkHiictrqS2wo+mgJnvYNwrm
VAqF00ZZoIFyY2VRHB9ughFcKwWeTh72wVXUAvz4G0UfUwnEQD/8J1lMsxyG
XsKZAAZlSjbqZ3b5HNn4o0VgFUJRi6Ayn8atJWeCMfiiEBaf4j3SuqVo0AS1
KAuinr3lQbc8OqhRdF93Ou5nX1cwFLwoS1NIYKdPZkUztL6DTpO2mSivyXiu
9j0gXIBY8s221rvgBxkynE4drRfHQczrRpDX7NvZSey3wkjvzpSHE8pjdSRh
IoLNX9qwdLVaf6mXKCuU5w7YMcDk4IOa6XEO/1BEMRDeVr/YcNYGa9WYvu0T
fNbwu7AIkZDU/0i8BXNzQCDnuXOROSn0fx86fDHEQpx7kkZ+wWI0NzUXRB7B
UcXX9lyvK46dwaDh9OEC/e8A/HFwWH4iyH82gyeH2qava+YVcDO4390UQp7q
XydMatmjx7u0FyGOvUxy3r4cI9U/AVmPvmByyhXmlw/iwAAXMpvv/sCkrvZ3
5eSiMdl7LujwNevS6FZh1bASPak7KAnmeI2lwv7qlDRTzEXWvzlaJiv2txHy
vfEkcr8ZWcR0wxz9eYYzzDa9x3mxmInbdxUqDt/DZvA2FidEk6GJ+jzF+AdY
Be+luMKuMYDjWQWIBmzMXjiOMYO0f6TOuudCS9rWLLc2nijZ8N6os7U5t9MD
Styjz8aHHkW7NgEMMxScmOEGKhrRt+I0dFLFIWyI0QJkBZeywMCoTwyilDxt
SttK4Uf9JeYbDRJMrLKZ8u3LVtbzEZ2Puc+axT9D7X2mmNGdOo0nyrsPQn9G
2GY+1B0Dy76zSIaRGQONedSXRDPMXoqn5MkMzSkio+bccq2ciEj9IvKimBXu
LrJD5z0dG4Bli3xa2D7R4Mv8fCgkmW2yW4xIcnGk/DW477yoKIHmCgbC0998
H22299doUlRwLU54jiYb93QgHFWDLocnL8/vhoNh2leYpXCNRwBnlgwdiyk0
34OFVro/gs/7s+DNZkhfLgv/6SyMeETh1bvEJA6CWB36pMiMLe+5C20QbgtE
ZaaoNhsgjXPG1RFgDmDzleFKhCQ9xjuQIdwQhMcCiLtCdNITC9W/Cq0mV6+v
9NFxwC4kpaxJqLZfa23PH8lBveFohDH3m3q9ep1b1gQLbXhc5ve3vor/ANqq
msJioRJPfZmL939vvUq3J9QiRoLFIRZNKVXyvAYuIhh3gnACh6w05NgsPhcY
eAUJJ6xB5Z3iJc4Bbo0uhd0EALl4BcJwMmWNcGkYDr8wFO0Spv2knXGkWFpf
DMAerIVFK9nhyTUsidGE49vB3t0gN3C3F7fhJmUDj1bBsyQoSORbymbcgi/x
+GAe3dDy1eiyNK3kqjJYYb3VjVTvIx5RBblrkJgP+XTiYnCWxFLaqlbeo5TM
xQPC3zgZckxIi23BOlCRF+DNpSRRIZVNQPRaA5wO9Cbqpnep/ew7+mCIDcOD
s7MiQ7AuVzoRXZNb9zeZTatf2zvPWCvMr9rTaRzzw3xN/zbnnIO01XW0nXJw
uAad4BkwRrvV6iSbiOmUb9x739YUwa0xQ8TiYYu4d7RUgVOgwxcQ+aobmujZ
CML7xTl8mbGXUXivbIEuE0uKCJkSnr3MNefshaWRhZcx+XvbTYlgPVdPDwQf
OgMT4GTPWWvzPfjH6H2jOiIWwRWOTxJdVMzIdGy940uFClAHmM9GubXy/+L7
sN1CLrtyGXhowva8ZKulDiB6yPTqvx+jYlCxFmMVlwtvtVnc7p3ksiuTOc9Y
VxPQqYGQdoHzQno6YvQFhFIeHljcSGuxN0M4gz2OWCDiTvKEamAQZ6prtNiG
TpXYIvD6ZtvVH05AV+SuyoYxhNgllWCP5SfUTASVUrSErzsAuf+NH2nhpQk9
/2T+LwRDbxk4mFNxxEPZ0LFOZhvRa2lRBo/f2ZF24kUZnxHsr0bKLDsN1aKO
xFpbxAuoaiHrR/3JQNT8ncFaLo4Zw7cvd5PY9WPGeGZFjmdaKGEl9ySQ1/KD
TQ0fE0Pg8diOK6GHcWeTXEggGEeYORYZaUHo5Ewy64KGo55nYP1Id+TqYNd0
kBtkozwsqw6r1F7rQnkhsqCpCZkLYo/ufq6Ft9eJcl4sErA+xajs98P7Em/J
l1VFq3BCw79tNBxUX2p14obtJz0rZi90/H/wJfaMmts7th8FbIy3VU0mh6BV
nI1A0weH5c29k6DN6/Yod4H6B+Ieibsi8AAgATtxjT32jXddNg8eCXEsgoVM
eW269WfF5yB8yDmeNmzXk3dweRXfB1SedLnnc4HTBAe+Vg0uR7lkofQVs/QG
llFQYkWZ7DHt9ccqKjYAy/gIcueRMsUbw9CqSDVaPwrypq0RKJdYvIN336dq
Y3wSjdS9KOEvcIWCvtkOHOysRgW5yxDuEtey4fTuYoc3TBf7jcIDaasgJ0Xr
v28hw7OgwllIBBT715ELabweVlgGFiMdlTSndH3yXfpavUcdUVWP/oHwOWmC
vmJG8OEu3bp56ep9YCAkV+JX7G08BSfB4n4tuonBmC1vOqasrwBMfoqA8zGH
TgJA15reGUxQucoSaG1l8IiW5gWN1Wn6CN1J1c8v1WR/1QepnXUM7SwiYqFi
oPbeFLxW+gjYyynjAENRLUfzLXl8Dh/Ti68JApHE229+erj/oHVOwOECOUAt
s7i2KRvCrDwjNF97BBHxQVR2Jwt3WCcW/Tvuor3WKcb/HrMUH6ksSOsM2dXm
w2HmLPDBsvzDxogSFggnjoUeQyOTZa2qSb+6lfAp2R4QJI4wcOvuiI5rngRD
Mus1tLEZGnoDPlwf3n5uB3u3lbpCfYBVseUgaGO5XzPGSz0uAEsi/71Nd5z4
pAmUlpw1Tg/sv3/6A7XXFrs/6E8EZWnruxaBjaUJ4POWdjecHGQbgwIAPl74
NKU4PpNdtm80DlubsWoSpBpaQ4Qtwo1N6OagGC1vdiu6C/me4aSkqtxVNzg0
NUwOzCnIi5IVD+kUhsju8lVcWI32rwpwODA9jvjR8aXA/e7zQYquRLKxHOK5
Px9CpqAFj5Yim51ruz7rt3+pKausY/3agsEOW5ga71hXgCBf+SUMpOXzHFIe
+5HXBRpa9d5K+Ff454YGYshCIYyybrIP6iW1N2QgTMELZaXExLTWoh5l5Qad
tkuKsvO98GGw4raNp/8dEMxTl2vgGse30ds10HFYHZZNrU6FSi54kJynsLNV
8HkBAITqatRBPpF3W7byY1oTEk71La25YCCVibQdsvA1ab0GpXuvJ/2ALs/F
9hH7KXuTBdcvVeY7LitcUOLDZi1FRm7c42wNAvMDGSoxRHhr3szej3+rj8HM
6ytT1SM3stwXT6/O6xxEOY2o9IOPEmCYD0s8fAaFXFZql/6hjmqAQBsyEqPo
zQGF9ZVOfohFfaaX52JAOc6yzjL3ya0zUudMHsIyPc0f9W3MT8ttFHXUfjTU
7S36Seeck3MzMJsumqjXVpz6sik9l3W2+Swkp7Vyt8mQkgEzfvIh5mOcI/Kk
TNdNpNpNCYEFJnnYpSrjkZEeVnZ9nYY3Rmd43rjLrI+PzPNrWqcl/N7CVs6+
kS6CCG/n3P95QrjplysiGLyg21CuKhj4BuyTTFc5uz3Vq4mN8wqJtpc+1zGp
eskyp1Fvvnp0wnw0m8XwpMOv362dJ9Im/cupZLaMFGiHNfgC9Y9c8dt/5Ron
mkG/ouG9ZPeop3V8lT1WAJzJgEU3+cDfYZvxLbpSnJcrRHVJfhAqomJSvGce
C+Q+YZ0qIrlq2yJvFFozUEXt0UK5Q9UYnCX+EyBP5xGNvIKusb9lUlRwXtpO
tRVt7p0rjMqf5ZAF5vl13nv96Yn3GKAIbTD9TKrqntTBvEm+uNO7y7BuMrEY
Ggceoi/GWpbjudNipkaLVlZd1dzQ6rDb/dkJHcKe2SEeJ1v/RvPvxlyvPcel
a0u/JE5qmcCjMRzks0nay6+935ipOHhoMG/9IeX+nf2Yi0HciZKB2zVBGfYN
2mcq7/th1rdQU83u3Ti9Dwu+qujVm085r7OqSve9/4ddWxMHW35ucLu94AeX
OqZtcmiwhxaW4qJm/ZbImiUgmt6sGxa+1dI0uyPIN7A5/jSPin/tn8WkWfuR
0QAu5AbZyzxyAbgvf3kXROp07f/DI1s2VqThIWHAKwch9wcqRCE1IzFQip/D
n6ZiY5u7RFYHo4mDHT50zYpyBotU7IFkz6zfWlIBp3x1cybZul+LoVbMXbWq
DY4kE2r7bDOF+4i23mE7Fe3cT6UEegR7YBF7HOPiU81Lkgxzq0TouszmYLV+
NXPCXBTr6Eg3anOl8K5onWpZKI2fmlfcjCmSFtVWESxw8KP/VeOEln08mmyg
SSNZkBYGk6oOceziKLKq51XbIMx41pxlTYgXlPgDPE6EE3GSBZ/v6a3oEGnV
XcLD7g41NAOewsBKmekT7sJ9D1eXn/Q7C/zfVT8UoD8nOg2DTKYwhHqUdxw2
MTjNvyAprlMLkK4LUUMF2YQf6yCvDOAZLSr8Q7kNa/VkiWW+DLkGe62/PxIZ
tHbVmZUYhvG/bL6z73IXcg3TdaNUzVvU4LcZHgD3ASa1M+SITrh7buiq0zq2
B+3VbXcs2HRJXmOUvwOg2aDSbbt78wmHOh9wAcBnXd7ZGRKZV8cnbEeGJfcM
KUp7OPr53aUxQA6aOlvSvm45TIS1bF97IB+HyBycqlvdMM0IRGFqFJps2Ca9
pLhqg0AApWhl+F9dzvRjS5Rc4PVsQckCh5WlVQLsm2RWcopXR7ZxzPtJYchM
NONIUJw+OjZ/5sLQx45EfxcPKgbVxhOVLDHqzklBMJvM5tDTY2EaGIn4NdPs
xJEDFn97bJfrAE7rO3Zs/5wS9TuMiSSQyavfz8L8H8WUoGXYV96AvIHclRNR
UH9eqjUEOISofqXnAYycYGXJz22p9RJWWA9aCtEfU10x6M9qCfwQyj422IOQ
53K0oNZOTppHNgy/wuDUmJkc4mP+Bu/rKxzQW2e7X6+fk1lsdku5MJQppcT4
00GYnV72gB4M+a5oC1mct/i5YnQFTocq8oEmWgJUDkbD8yJuayCuc21SZ8Ye
fydVISIA1Wy/wRKpiiAwgM6FH9JTDCMbp69f4fouZx53+PBT49ntp+PeJVg7
GWq66XIec+jEm9NN4nE5GW/RYS3ycPhw4GraPUQXCgQPX2yYBiYH0cVomx2x
QLuHvgJDYEbyC2uB+1EvT7xNLo01anDPXwG4VDABp2bySzN4E7+u5Bgir4ni
nnYrbK1LxTI5FrrJCVGZekvFN5Fzd869SayYi0Sy2GPulXCrIpuGylA/yFOK
b6nl/ZQEKn/AYba2U5ZuQKS5FIWGHkEpXJybzK1PBJRYfdZPL7bvusac43ml
OUrK3j5nOirX1/rq13TeKOsdVpU923aS4XnJivy8YPI4QOJQLBEYY67ctZlJ
kizZ3bDcrmJ3ER+9fdJV5YEqoHNC4/I6YeZDclyQgzIZNClVUFWNJw82Bu35
D8rt700aNhhVvrn3AYO/2QxRYnpe29t/IMZExbB8yupkFnhL348Gj2iBMJHT
STSmT4+QM9pBzptRus3JAS5rEOAxZS4nj0usmwiL16q3by42whbBta8VBSh3
mRJU9btT/X3KR1bg5Y2CbMI3H4uin+6zP5pN/KPUf//xujVMKpaPW0Vfvp1e
eZ9t3N08xDW2Qvx1KgqqbeOAfMNy/1C62aJiClUwCl6Be8zW/kRDTK5g4/8P
DM3AeESkdpCcttVwR+nteY7uhwIKXwGm7ZZ2SiKh35A/q5grvNm+Eu9tRfxM
siXUFxb5MXJEdjW7uWvJZqOB3PKC3W9+mVGQ8rvLvBNFMUUEZC1JwknbiXvG
7FmWX8Grxc9GjmcP9Hz3t5LSclof1aXgkBymhcxkCh04C8qdyN52i5vqbtEn
QIfzotqOn54zQCQC39+24n1EBEXcGgzfTMk4Tc6h2l9pOwTcZseUbmenFVGZ
8/hIphEDpTmsQc8Hu4HyxBbr+3wMGUEjIadqj97wSnfiYl3oHl/Yzho8xAGb
kBSsh61/Huqp7W1kv2ikqaxVADTTXBNkNJ9lG6eR6EVHCK5DcJj81mQB3/MN
LnK4zxPx/eKECo4RPrC+cdJcWyostaXIVvkYabbztb5W3o0hNmOFkGjvnYSY
DVOAb/t/NXYcu7i7OWVTOeRTXZywErxFSS3rXA5XmDcQLagXvN669pmlMchX
RAve6My3GLy4Og0/cgFqu3YL0tEy7tihhp51fOJK2tlTgN4vdGQl7NQ4iZ5g
Iqn+N8U85At88Iyt6gyH1PvEl3uoyi+BgAPqLXGbubH/2OyjPZLwoEUcyBil
QSPpTQzvEIkwHKbBhz0Xb9MUD879FtyVfg3TjH+Kk1OKgqxR1RfaTIB6yYHX
jvkUfCLcAzA5YJb5elhrxTCMpe6fv7B+xd2vjeNf9BPhcuzogkXunAmoEBzi
+i86PPmv3PgeoP7UXcEuWhGLbTt6yx/UJVPuotmqr3hQ9YIhUMYFSiCoydbY
it7Q1L7QA756BRV8RBYUscArFYLRyb8ZsnvM9q6eidrl2y/LpzF3rsIQfuUb
c7dm2VO4u00yxKUtvQ579SasuAcS2Xq+UkGsPH8Bl33I++3Qrs2gCJyN1tNa
P6UHlF6Yv0D4x8XZ5BbyUYD7RpTt8uKJG/SbioexED66veaaHynM3vQOYMu6
YkrzuW4EVHl+UrEaSVoKGxmN92jSnMTdTeQxzXnrDQHbql9J2FLUGGprYPEP
Gp0/NCyJrgb6uRQ3EHKS/reqdkqITL0EYq468fTIlu5WRg5vyQL9VVPwZHri
Ol9rjRsjB5RmZtxoZ4iou8HaYGynBfvJqj3nrWNJfT2gMmN0Kcgfy3rrwFAG
appQzQap3a1o5up8ANDi5benAXBFxGXTFY5NAyjeRop9SY5E92W/nC96etul
Q0s8lhWLtUlJ44uds2nHKKm7D54XGuobls7Us8PAL6WA8nR73ZMdHLOVG0Ny
Yh6QyfTCs59t+N0ZqR6dExkP0K+kJS8Fimcw0yb2UurJeMSQJnvHGPerfSNE
OKKyPjXSe+9WUWaT6Nr+ArZt/vrYfeEE1x7cyC16x97ZnILIkc2wy4OHRzhr
PNfUaMOv3kiv/yKrKU15aH62mD43rN17wzj0pSL4663Im1IceUSLMEJjbZFo
hSDu448w73aCmoYJ9g9GYHFgSZZDzfuTJGOBvvtgx47T1rHHp+FixrTzD6x5
eaeXtjrblFZA/N9VcKP1R8fQpIfp1ADmg/VFmHQlBnVq0kHr/tDepTYiEm8U
0ZcLJ5A1uOeqrl1t5zZEbCbVXkbaUWHXci1xPitCJtYnUcnXzhWrgPGvq590
Li+VvYjFtRvPi8eRrwxzrz5Qd+2hIMuyMHibB0rVU5kybCppRB5fXW5SK8/C
pc0YZpSpbA/xDpIJOOpfpcIQG9nIqyMKUFe9Br+x/UeM3J8RPnP54Ef21M9H
wnjrOF1VWJvFvodrwSyCF6w2tPvYa+fBbY7RpvmUzzSrn62TVUfyYIX4ZO3J
kXJmwvkZpnsV9CwBuQcdpPV/e/4nFz/pIDJGUq4Xc41XsB7tH46LpU1A7Uju
4HgrIPhdIE9PDJ71TXVR7JfnSBrzo1k8tBRJDAnv1M3MsYfSgELTWz9tfE58
7INQBXgpKc8Lfh0TOYjcJUtRuhFz7nCEtpMRZ1fFDdTfj2rjbYS/gesRTYrr
9OxwtsaD/pa4VbyfqfTImxuu6DR/G6JOzX5o+40eFEnE+HFIozwvmWk7Rw0U
/Ws6e7En1ySrLkC6oepQ1kWUsFzu3Zs4E26mPhlbI4cm6ud1b8hsqWtEGafK
g4QVtqCtfWrH4hWmLIG4PUgjlRVoLwbu634726hjn+p4wdToK+GVVGruoA2l
Vbo6dAkIHkVfyeJuVfLksf1gck7x3r7rTffP3OjEMiOC6qud/WnqTgyNtjAO
yKDBKu1IrQ1Ps75TH93dDoEhoyMj7zQwOP0crSR+Q1WP6mYJG6xirrpWqQO1
91wMlVrrVYSpXuzzdh7JCwWfuTgMka0wIYA+Op+8qyvnP9oWTNee8QVpzw/P
uhj98TmRR3CEpqQ65D+9C7IfJst+R7cIpTNmkOwbc4CsEQ7iZRnTz8XfIUd+
0VU8Yu9DcLbaX1k/XWGa1d0kahwJk5I5x5RwjdjFFvmPER3vBLpHNOtHm0Tf
GKSO1TlLmp14SkaTLTJrufie701LuEQ5wKz1SXZaTJmf8rJatjU5zJBTu4k9
pBEqSErLd132UboZ2wSpIGIYOmDt22bJm4hC4K9o06nPbGE8GLuONbs+SdHB
inujcndyJ0G95UmPwcgj6QtECDeLTkh94UuXmdaFYukEl3DnvGWB5fsgJ1S5
iZfmMgqPkkJFPpGIHbVfcNVj9OZrNgnZ0SDcZ8TOX4J+3MUO81L2DI8y+BSw
/91uTI+ee8jpbzRQPeYUgI/knroRoeDtxfqgVHv+GHP2s0Wj2J0EmCHyztP8
10sVWcBwYDId5iJW2+L047wGvBOHiHgqn7QugFQ0Lw1eHvgpJ6NMAnwp2egs
5wJtZlNKI5dQpVfpU6PFC1uRxToXayZU7DLOi8LdYqSSM8RyNT/mGIoZwfKY
8NMEwRp/m/OPsV6Al8fVEgmyVptC+bH9iLHGgANk2dhYbI6IwfspMoThq8Kj
4H7wn7w8Nu8PZuRg+vJZvGp2Bs+UxWRUs/RDy4cYm76cccBXcmr4pXXhFzLh
rSL939JdR90ewHIi+jHLzjOHIrMApsb7yULOfMt1oKQuRkSRteeI/38J/HDC
4gY7YU7I5dVmvz4aTSmJ8df2aAESq4Qx/p5JviHh1fA9bFZO/4sIc1JmK46J
F5wyAENFG/bkiN2qKRGk156KehZ83m0rFgg5A0KZw+e3JcChJfRNKDPEXMdZ
iC8jquGe6ouZdH94WExr5Hi9ViPb3CM3KjRy80iLmgcGxz0EfQwcX7S1zqAB
CADZ++PCqJfdImIFM7qOYGFOvPLyRSiIdAoEm48Mh4l4YojoHiSxAydpDdOR
7j2ads/BelKuqL6KgCc8uqRNxXQ/82gJsKjggZMYlxcuwnwRGUvCPhXU/qq6
lXmW2SaVK/DQRIh0qui9wVODZDiYTfYxl7lmER3twtg+qLM1A7p1oQjEUlkc
LLNfZVH2z51h8I5gAHpoCtuLbhCCzfHfVrj8rQcwXHZQgdCuYe+MBZq0KRjT
LoW3feGxjr/LyIbwyoXmURg0ggYQmGkOtH1RPZpEXpK0SmRrIaqWL1jnlNNR
X+Wodv61mXi4Y+dK4oA+rhaWn/Eb0tcNu3GU/UYVOA7NDJKBmSLPLc0Gf5eN
2uIoGXu52LyhF4+mvtNDjgaU5+b79a/47kDAeJPujLRRV9IyyEO/5Nv7JwGz
wUFRTPmEgdvJQVla7by+JqINZZhutseyOsbHAenIkPMlif3zetptr43vjbpp
qqombLvzLHIAnyy7h3mIh/fCJyXxgojN64tKuJmhrkQiWyvQjliJfJmK/DaL
Mzbqqa3J6CNtFa7wGUsxScqbtY2SnPUeyLVYpdCd8y/VjfW401MSMVhIeqdJ
IRL47wk2AeLuNBysmePfmK3Kjb74UavHcK1VtqY3LaEtjjtElE2/mNMPqtP3
dIO1oF2sgLb8I3ATIdr8ZviNAW8CeeF0bw8UiJVacy7w+wx+gwTZN4aIUSgx
AsvIqsbW9mCVMbK5dNZRslzt1c/nmMIMUIeXkpkis8aSkKQMo4Gya6CnyJpT
maFvc1PYNz1FlvphMT3tUObb8GQG5rMjDktVxVAqg6YsxbiuZb0vabxdLnzl
MDJViczooV356v7UCL46I22JhvKkn7HFtzmxeUzin2SPdD0S5A4cvSX8EnW1
nx1qkJEaEL4mbb0f0v20/rtspHzV1SVOWc2G+vJJLW5KN/9bYn1axn966FkT
fpCs65JsmeOvsUbeOBragtJq/inOADdO+ttDS1Gsz8CfTSypxTGzpY+sxIkt
jkQYPS3y0rEUPB5q7HZ8ZPfR0PurFTj3bP/BrxiarFyHf0m+Yk6pSJrpMvZ5
zdicEeBttAhOsReROSTTCIm5X10hN6T9/AF6lYCpCh7aJef3+/1AvemVtupJ
ircHIA6f4IGICi8GXdwNm/RCEN/EDYSri0DkIUkCu3rxscBqvWTaM4U53ota
WImrLU86X61toV/88wfdyUsl/2JGFTE0Lot3nYFs+/KZfLOu1jjovJhKzTuM
wppXMgx5+spVu9pC2FVE6AFIflIBvotWUs0mN1Xw2698rKUfWj50gcBZoJJU
ryGRuP4J54f0ynX6/RVZil7vslW2vVmIXLUAtxsinnLypc1OFZ6gV0KdCpGh
cw0kcKiI8hZzvK0Zjrx/IfUTRBIUeHPRdLDbp/ARzkxNcYjGgGlSGDDLCrZw
XFdyUo9SKMev4/bT6mX17Uqo31t7JmTQd6UV+P8IgbOQGxNC8mrN/oNR8ZCB
7X89fXhGAMUPtdbSPl0STNNCIJdsP0Bw7VmVY8Re+4Glaftpg6rG3kjk0NgT
fshdSbHwhgBYA4UO31l7nWLQwFuZY7r5UwACkFtohjkuLXKDQ/YTJk2+DcR9
2ObipgBW6PDfMJalSwVHSY3HvYV6EmDD1QAdDviuTLZ4xCKvuSsZ1p+buzFh
2j6NrQ2SVAWORR8FZ4ZJ+/gkVz6uWyU2sowqaJXI1+4gU28xRg/du6iyZEhw
YjjHfnqi91V4YD+3HTNPCe0PAj3AoO4CWtZGSa9H3DJv3uMIgsGY6XuivnS1
yyVQJQFSH9ehNIc+i6crIfbMuaxMIcCEs3i1efugunYKQKLF/382/HMIdAEO
+IjZBuX4yWecwsdH0HE4ZWHJ1SOREwY1JCce2tF44fQUhgqqQ+7WcdFXlWGf
rlW7cxxdRzJ66ybAMx6RLANL5gscfg1pz4GIIk8eKldbE9iEDCKG8hQqm0Qi
ovnJd6cBr33ioyRdenDj+Z2I24YSJ/n3g2dfv+b5nxaVqSnEdHufULV32aS6
We0CK9fFVprDvG18zKYIGg7qQxHTgDxUYje25DJvV39MCY1oPVvHAJPthIAs
/UFlNOs3pzC77GAh0Koiw5HKDsp0k7WpOUZ8SS9eDU+cs7ogjtTlRJSeqhd5
daCnniFRaa+beSS6x5d0Uf4+f9+hYxDHWkYInds2whlxR/JrgNwaxH6FSkOo
X8CzJ+LdMy94cnPSaZxhDxDvrF69vfC3Gq4Dkc+EWfLJ4QzO22M3HVm0ZG6G
SWuAZ0/Tkp3kp6TD12yCnxjBh7CXYyCeQDDr434sNICy8wYn+ul4ZpNDVl+s
2JY7jc4pAVxK+i8GdhiacS4RZKm+SasNhjqrDMntq4owobl/xtxTHVUT/pfd
Y7H/nSRyl1gj8ZN7E1m4pV3A/Ehr3e8+H6MMVLzu6aaG3JLS3jpzlsyWkuL0
/aNeI9y+Jtx/w8Ur9ytO0kP3m+kBDf+wxfE1dmRk/Wle8mFz7fnarkwZLs3e
Dp/Y7LA/eY0t7/lr3flTXINM/sHLYSUcQhjxTyLhLOSHQaZ1qyprfe7dDusK
uEdgu3ftrcTI6h93LXKmpkxBGsDs8yD/IBpXEGGhKwm9LYmRaC9znofV9mpE
lpeISGwtmfMGPt+kPZMVuDXnkDylAerud8HGaXffQCUVUtHG1IskkYwcmayJ
1wjMoi97SzELdmJx7sGUqxfpsJx0OvkKm7IrbmzSz5cMJsdi5GarPxYegjub
J/h7iIhbXmiBCj4NxK5I71jHBrdGsNva/KoB90kBIVQUK6qBAVV3Asz1hj0c
IGWq8qXn7AefayJh9d4DyWmqYqUh7c/705MMGf1BguhfhKMjqvOAIdw8jZvh
aPK5f299Q3sVlKpXHsoef5jV2kMn5sSuEi7+snAj3PthFgASOwE8bR6xeiKY
tG1scmYJIma512ON0xpMZ+qUCRqX4JbZG05qwHMFAgIFt+y2qgXrdu63PBac
NII0PIIIyECdqWxvaoPQeBKuWn3gek9CpHlG7wIYeJjhyaaiAPRHrbEe9+aQ
itJnoNTYB1WvgmhvqC9dXzMFMonV79EFBnoDEdnuQhTEMURkqd2iLf4427qG
HvLn8FJLPqrjB1ltrEsJiREvXnB5LEsK2Al+r6ikxO1S22peF9y1mm8qWHFr
NwkLIxEHs0TsLm2mOjHEixdQjEqD0OmhA2McVSxJ6NnLMdWpKo39wNk105Ud
s/RRuYPK8mJgTA+mQTpe/gWRlCvWCw2jfNcQzB1cS97ndLT23+0u/XGTwPTr
GmjJbA3EgUYN8kVmzhcNWpF5U9RphSes2lHVdxDYf/LuNV508xvxExhTueOq
eDlBeO2JKs3jP3Rca/CkBXrOCol/3yNwOwqP4MGe6e1N/IXEsFscVHhtaSqO
xMXPkBWB9gvC+XqV59dXAgM30lKnLVeAP0bUhlA5qGW8VHU2EgsTejaYn6Go
OQEJQOk8nnqy8K+hrPgnXn82ep6vp5UjpehccZoIg+LQ6IID4nyqjakubDCf
BWcnbsTsFY9qrdfUlJyAJ+9o+lvUwGuYkhD4uWKdoLQRKhTYC84nV0A5myOc
gXQ+CZa3dc671Te1PTP0vbBsSUzKQYTQfYXEPIJabx2VlG3of9FsoM1nF5Vh
AOHWyDtsihxIGHrqJeCSxuRg9M3KJIMQRApAvIsOwNjvf/q47pT8Gw8RkGW5
bTstwhfVpnDJ7Mj4Trbt6VOoDEgT0thXPE8n7L7Ux2NyE/OmjEigFoFzuyNH
czMsHsPZdSj5Q+QXRfjP+vDV5bgdwfygh/rl0WC1lxzHbA4jbVJA78b+tOyw
wk/2qnSYPQRq3/kEnl4MZWURz3DqYdeTqSXK0hwUV1pjiwOCnfoF49uayrgw
y+GLRDoGzrSvy4ZOdX15eZ6agcJo1BSV6inIWnMTE4WviyUeF6HUMjhiVlvL
nXJK378pXvaObCJgz/A0mefZENbzxGiiEbCnuE5e5qEcT4WTaPgGzkvNl23k
9K2QoU7K9Y3EZ0WYgqdUur99hZr9ebrcAIRtU0DMSQH+Vlpms0HIbxe/0j/e
gFtapbguLwlkS0NTMsR7UpAc9Kg5tSnok8RbEnFL4IXTia+1Nzxls5nFuYUw
04BUWB6LI11nkNFVTdimImn/wdz3w044H5R2iYjd4KMaO+sNcv8i8I1KudHy
3v1P5OpjAngJB6IvYJnrjrCfc8v9Rqxyi8qLibOLYojKnyRzVC6yMFfkCZVl
Gj37CYXDgxDMJnb8rWR8eZ8wmUDMPczY/YHpgtgH9CwoZAjSSNvsHQC8crIw
MWoSPA5L8c41BBUbOnnxGVnLDLH0iy8vAKVbDlEwVuxG42ip8xZHgzzkBvu3
tNmRWDoxY26Lym1WZqfcBv+gGF+BjSb/q2E+4gzzENqJ0fuqyXMSifxE/8fQ
SNL7rDLMW0A0myeyDN9ftRvdqHBlvGidU+uVTI5m2DW02vrVMWQ2SJehoHNb
RbS3CU0WLeOUfez4s/KZqH1zM/Tuy5w9YIGXLm1Yz7ikQDV3zipG9F/NoqUC
stLD+Ttp74zjA9/pDfppMPaHYrzIZeDbHQg7cvJGVs+/u2ZrFl4H1zgjA6aZ
z2jRKAKKAw231EVMubvRrZXdNy6fjMMadX9J18HxTNbRxaaWr8PYdY9fphVU
BQPuG6v4Ycw1cWkXJLAm35jftt3tmvmFfgnqlCUDcyn3gCN6V0Up04UPQl1t
jxc9p0FW4owLqaeOIPmG1eNGu6HzCV8v1Qf65dEzN4/0Jv+hqBdqbNJ3VVQk
6pQzutU+EjwYKQLFXLCsaJYmIWbztpbAk2QJCnQTKK7WB/94BZiqa6+3ubW2
MBLDrS+Z2sgok5KoXy++sjmi0gbUEOEY5jKFyK+syMo0t/RymXj0PQdJ0sui
uuaNPA1sW8m10Cmraq8mmWJEgKcq2SMQV33F4PW2DXLd6FV81arUtR1cxu13
bv7X2IgNo8ZDFtAry4hxhvM2DHlusTrC/Dg/3f8gmCTj3UO7ST506tCNvaIX
NXHNUN92xln1L2pWMPZjB/9mLmhjfDgv+rcr1ilYmpvwdbj/3R0G5nlZj7Wc
S0qUyPza6DnIZ23/4TowYLDfyIGpaN8vmWnPLVPNF7NFATdQSY6/Ff1MF0Gi
qEQ9jsVxo3zsEzC3f7GIT43sKNeyat/Q1NXi68SzujB+mFLqRcrVQ05ZkytS
5qKlu1nJp/xbwuyY8hplCjBdt3hq8IDZJGTX9y3WdE4BfPGOllme45GjkN2V
ubNYDcRbQlEU4rG6+6a3LTMTDBPAN5zOT2ZHAgJEMlqduSUocAJXLxfCAsqj
UzhgvtL1iczpSE0MgfX74VI63y4PAJnnCIIQfFyJJeWMhosYXG43kT45OIJK
h3QXyK5+CnJBT1dcR6ML4fuhp6h/IdeJyrBswDVpLJXLU4XCP5Yk/n/X4YQg
GBtyv0MlBBppjDAiCeHYWawi0owe4HsQKfRvmgzqMUi2U4BIcSe/crDg+qiM
T9P2P02TAK4pmmCYkxZl6QLjhZDO+a0eB/3a3m44gzz+2DFk1MgHepP9E4sm
b0LyiXFmPLWGY1hyNcEOlGgnaFZGM5HKh+VaGh4TszKHVJfzzLo4xSFeV8Nh
FPzxBAMb93KJ0qiIy4tKENXY45owkO7k4DxjEAFGDXzyF8gnEHyGq6h/jfYl
Ly4GmljAdVXO3eL2AAikrPhpbDLRCL/P1t7FwRK6o9iriWXDnb9XVdecjK/J
v6jUkmiZJQSVBL4h4xyfgCUwz2qZwt1eOzSznuHjMt0vaGlXCGwSbkdu5EpQ
uOpf2RBCv7uO7hGViHLYUuN4v8RK5d7Wo5ITZuQq6JRGEI2V9TuU6Ts/juzB
QJ07fl3rENQoJb05bQ/n2DIa9NTaCAOsy94Y2CKLdTKzlI6CuqRVv3X9KJuN
Z8p1w04Vm3v+s6LtDpuwTC26tQjIOZHHfgL4XmhWFQKCrwY3OjbbAQ7QAa6v
Y42S4udZ/Vh+QMt41hQN/k5SuxKPDqAmUUF2IX3bdOk++11H9lHBIsjCxu95
Q7gtqpl6VXFFF05Mr0RmWIxuZxEhVGEvvMqlI/2C3QO+O7497Rwi7nLAa4Yt
rfeKJmthGITaAYcEACOfq7W7jd2GgCu9XOvxKkjywGoeWbccSlZWquZEcAoQ
k9vYAz8jJYixaeRsmL2TpfR1SAUqONfQ/ODO+qoWZgXDkW+fzNtmEgZ3sLpD
Qr5TNodfvqDj9QGq6ehksjr2mRRd8sy7ibXz3qQ4FbYG2pF1xKo/MT40mcQC
BUm3U/UuM9MLvtVcT0jiLH/HtC2GYEjq0Ub4tN0/8sX7571guBepUie7NrS6
fFECPVoeRIFbYUaE1x30tm/wyhGcZuQ1h/rFUkcsRDB5AE/AXu+7tiT20FeD
BiLsggoCLHCE9TAlqMmcDyLbZC27/NgGXvw7OFpjjApj+bjcCNDaO6stiZxM
e0NluBjL4sDkglh2V5Aepyo6APQFl8BgdJByVGb8kvUSSsACsyNRTfnrcDie
4eyXdfOAzfebIWJ3X092JdZc0z6lmmwyPLeTd8Du/BjG69UzD2waXXg/Qmdw
eRs4KUQcAhAhVuNBNXi6kzRcpYcTEIuOuzDzTv38HFIAbk3hn7/4ymk0RAqe
Izgzi83XPLJULizukTPVqtJ02AduRQNMeyfMUSnF34cG9uXxqhVpCBbdZ16G
XNqPnJFBPJxOcvIscZ37oqoqHCjyaWcLoPPjyaET8ZK0UjJ60/4QHrA/bgdZ
yECuya6fA51/oWDa7U3uS5Qo2Kh6NngImvDW6spLUjkrwcr5em/ZzlbxJUCm
9N0Af4r9Q7vbrh0XVE8g+Kk762sizNy7DHInxi44aS9qLrThQigMAA9vYoG4
nKOoII36j+9R1q7q9KffXxISLGPxrzwmYLJ3353ay5BG3sMKZfcI3Qjmj65u
h5a/xfxFUD1KIu3630TNktdzBAMYqxwXS26+M688Cn7andNBg806YMWnaVsE
cFZvYeR9SL66BH8lLZiB3dxYfxYIvtbphxfNhgr76eW7lqZQT0ne+eklu2LV
QD3tuLQzO3OJ8iUFdePYP2DKCFlxX20epBiQEgvaVmJTD3Cl7WFgrC9TNzQx
kIru78Ir/Jm4tSsmCVOIupI/GT3DDGNYrgpSY70ECB3bKy5+P1DFjQdwsksl
ZdQYA9eAxXqbbj0fUq++lt6WCIS3DVURvjZb/6mChiLpgHfiEoqCB/XlFTj0
WIZUfZ8E7+zQrhGJVzNFnZOs3tP66Pnf0rwnC8OmF3DtaWGs50t6eXXV8FZ5
w1S5AIKy8RecHSjlpzD9cQEYIZX6YkJzucc00o6WjcNmdzNhoKAGKaZFSlKE
M7VgV62/1moejcDLsx4h4QcMYjLP3eaWvTfqpG0CzZz4y7o+MUamjz/jUzk5
qIXl30svIYeH1JChczmLn//QDWUxWs0IjWQxoMehAAzHJAy5n9g3KLDmOSYB
AKmX4kRowZaA4eKR5yWyoKPD7ntKAQKz1qioLFLBQYJ27dG0DrYtZFZsbVxU
MgUSPo04Ju03gfZgsWwF/2Wb9mE8GcC3Sj2jf+IeGd69rvk0wW+DFkIkAtFG
SAN9hceCUzyhHF72P/pJtd/SogL70k9TCr3jLfE5/pDTbM0TQXzbOdymaL84
ez5VHETpSBPFDukE/ZCIVPXyq3lAclxzg346P4qM3fzYq7mVhy8xyVF/vUtr
n8+ivd5PPXleasPspC0gbzPAQNPY70/u/D7MLaQHHFCnUL2o9QCSV5YZtPcA
aGUOoaTifRded+CaadMBTbOeB1fHAkXhGu//sA4Z2kfM70MzoWb8ynjKmFzx
QhyvVQAR+GTx5Zi3pGEFYn3DS36qAgSi9jeK8qUPO+fF7XUfDDW72CsSY5mj
2tgk5KwnuMXvlyKFEdpHlFiB0uZyutzAG7cFHzPNzFKXs36F7AIIjf+ecjut
N2zKuZIKsPkiWhJ0Iyqz0UjGsfX+2AzhueS3+bSsxum6mNay8LpC2szx4XmQ
EvYJDg4BYG5Nxog+LMznSy6tUvm1DhsSUIHeSDpPY06MuDJDC92XgLJ1RFc6
SYO9XLlH4S7Fud1IVY1e1N7Da4ISIpVQLBT89Gs6L1WwBEmZSEr+x0Fkbdr0
W2sO7Vd+FA1YVq4MprQ1afzbwFGFotQUvfAsEL0nonhK5anZwg8imatveIzY
pWBMZX3PsbusOe4Eb5PGnDywfLE7dVd//sXqTallL3C6biX7rSxuAopDjk80
iw8bWt9zxMA3rENIm6PvurZo82WhCqQAfd+ToBbzK4UKK/RqMKxug2DTZR4y
Gth6lGGL0ESv3+BC7jR8fBd1qR1fm8I2ZfFLqjo7IylYKPRaRnpUreT9BpZ2
j34m0biGedtJwIPYmbzkbs1D5p7mVcPD5iRLn1IpdMeF0bwcA22wnMq9GfNh
+80rKKsOb3aAuch99B1CUVYwi0J0ji9odfU3XgsGH+PaUhV2vAHI0MOMIaM3
JSDqXsp/4CDqn1ItkdKJzS7zCuNCzaPOxeWn4+4wVaoT82UXkUDFcR5tCKTv
s/nAKOswl8ZnIA78MD94Hr4cgZtwD3CJLpoeYA+u45Mb3ffmW8dVeYAC+Gj5
uB/2SpRiFmN3h2YvFvBkhEBHeOnrLw5zeJpXosmolnwOIeHoQ+yjaJ9OZdBR
ovUFll+l9H9vc05QXX3/nz08Oq+U/Klf9Qc1RNaaRjcoB0/iizssyakBEikU
a7WpJuX3gQ+fXQuCSL+WCDk+hwSueGk120Mit6ZYY9eFb30VPKfmm2zl3N1N
ch6ovRXEa77MNi/1GQyJ2eloF7sXgfUTswEZbYXr1UtaS3Vt+G1uF3EWMUbs
dWsFH7mIK1PrECMcLJ0gQoNKa9EUIYUJJtq0Tn3CXxSs1pBPs27SsEz0j/0b
oj2JPJR/QpKbPc7tEx9jSVkqwZy9SqzAYP00jmRqRwSAJ7HBSCaRl3h1uxwH
9rVABQVT1Z48aPQzdnNVqpV90kxIAdx1nImyTJWM06Lhixu3drGS0IpwHxBh
2USi3dbptEacVrA1T/VNy5hrK6yoyBCn82tbrQ6UyKNUQdEfr77oG2sgcOFL
coepfkGhztAzqBnSgscy5waJ5CuaIYJZ5Hd4AYNIi8S+ejGrQpj22DDVC9MU
kvQHAqyCQTZ4ya76JKbioX9G+dIlDxnRy6wY2fdDFYTNM+Tn0PYC0t/KkS40
xOnvczZ4olpOxThj3Qh+pcAkW4lpankCdHSMBpUEAt0M+z0vDDfgvrHxLA3t
lGoPokVhRaTKRThTALxBOPkCUGPBhR8DdTx0f02gukwAcfDiJpa+QTdpieqX
hT+Sb1fM/2qtpOflX9Kdhmz9pDFITcm0jEWdi6ke3rJ6tN6tPOh+upSCTqCJ
UeCe4BMdddVUm7Bc2hGnalIPzIt9oUoZLMxRstIQWGvX+93/Jb8ush9DqcLF
bkCcM++ld0VYg30Sf5DRA/5wjoaQFyc+Qy9fN6AGjkrU6v08BZPdzcMM7C7F
bzzZFmt2TVAoSUi7U3RQQIl+NqkTJRi1ULasPk6YZhOyI1cEjNafA8MhfiRA
i6Z8SX/NPTjCvExnC16L0zpyM/AaE9GQzGOeZmkOBRiPHgxxjYrRcB80Jufi
0Cq7e8EXo7GUSbIZtq51unTnzsQxx3vQZfII+zCaUKy76/CXPMSiuGaRtBmT
pS5xttZ9Jmb0HYbtiJVjwmqXfYYp0izSutQM00DO/ofreg5F9M1G+zEOjQ8V
Lb6ddnrEd8FluyptRnYd1oUsJIcU6hwFSLN4Xwmy5Iibsuc8H8eznzaykKPp
0IrThLgaCTjnuM6/2WChfkQbFtdEI4wUDwSTuhcoi1NEz6ZggIjBHkEhhAtW
1seB3ES8PaNaC/NO9MK74m36Lur2Y9Oc3kQ7VXLwY6qNmIEuwXP6eZTRO8/F
p1OBx+3Io/dxRzEqK7310s/d4LC/Y6XZAL7HJy81wdvbm87jWqb4MV/jmtsp
xG86m5+Ok7YGL2F6xIVnQRDXZD62fgxAggLpmcLTBG4N0wsx+Ib4QUrxec6z
E7MNzqiGvE17I2F2FBdmVgYwH0wkGxwYh3DgvDyDH5xecbMoa1UJX6De0A+X
WRDd/AU8MxOQH+NHRCGz8irSEXRgsOsZ+fyddOuJRmQoBrecLead5IKiJWIP
ejvIse8T5RgDZAHGSyXFJHdC5A700h58YINAMro9QuLvciWcashuxatoFWbE
3YGD2Dma2UoLXvOATfrCLUF2kQ75aWrdE6zbQAEFMJqKk5CTOvq0par8HOph
WV7berJosLLyrgNFeTp9LYyOPGsTCLSryUXtvas5T3LUaWdfP+IOAn1EQ9jh
UlZuJA/Es0snIVdodphCytH+/tcp/JTHjm6QM125hDi29hKwHSIB4bnaf9qZ
eBPBvEnQ8FI4vyQLPBpFGpSdibfX/BJPrIl/844NhB2800gtxA2uLaXK5K3h
PH1eu0F4IEqtsjB6HBgh1+5jGkCA0ZDWSgElDCn4zXpu1koNr6ajz2nMxZjj
AomMiPDEBiiYOfEj15MJoGiVbTqPespcd6JahPItb9KDUQZKZmPbyukDOGtm
l5NTQYRwaNBK64BiBJU3t/wFTXfLYbYMaJENsnOWuY7pS3wbY2Z2WBzk8R8j
QgrnhVyegYktGIiA/wvQptYGwyshs3BU8PBCln1HjOnCv7aft3rlIAdKz+nU
mGIOqSg8hUhCQ5/UWthExnVgZLK3JvFOXneK6OWU2K4Qv8njbTAQMKZY30lq
udDnX8OH5Sv6AmGAXG+RT2xJl1OomjxspiGPBNIAcuFGrlVDS6NI1gksDcd3
fpC6h+BvqhoOhzJR5tTQdDOzh/ZXxlNEhu3QwVU6iZvdslrspf2WGD6c6w+T
RqihfEKnG+/83JYRHqTNahUYEgKnUtOlS9pNfGmuzeV89RpC+6O75tnOcAfX
sjqg34KcM3OoNag7K+ZyhPjfJ5SLtIp4X6Qp9x1EBDYW9Xm6AxmKKW9MmHkH
pAx96whLu4YDu1pwc4XmcEzZxM4PEVQadGRXiKfJMCQc+0UfoHrz/o5gafZ8
mJCPW7TlhWXXnB8wG0Rg45cKbaDr2TbdEg8ZcmZ7ENP5WCkFt1MDYg6DsMAf
LUKwn0X/1oqWFz5Wi4IEZTgyWP8hW998e/wMeuG6+9O/mcOQ4w9353rOWKZp
cDQ7MYI/FrEdMcIEcIs0b9Iq/X/MPqd4KJDGGnIxOaiztUkpi41q+Bswk28D
1NpNIYTegTiz1Q3R0A/i36FKE6jkJGHoqi4zNvOaEX61OeSV4WAFVTtLHpcO
rrTlQRdbkG7pIVXz4ho5zNnxoHwW7NwbIClPH9vR+yWuk/grxLFsDIsBoOdN
RxbUsbwgSIJHB0/IlrMTuz/tCb10GKfxcGVUoBlN25HaqVUAgBP/rGBjkjR0
xLuh4l3AFk6PW7DnNZqOlPdLHctLreXfOwY4gCubZw20xUE/3lwxTlAcZ7Fm
LA5Cp/PFGu0VcPC8t7zxL2iIJDdw/evt8/h6uvAWgm9D+8nvipVHdhm5rLJk
QxnZrgoh/bK35kxTWcWSXrEvkY6YdDUsPiprMrEkFYQ1Ry/5aHDb5IHsyKP1
7R0XyduAvUgIPq4clgRMU28X/VaNpxjbRD/NDdlAmtw+KV8tIzSQE6NhoB0A
igLTcl6x7lFp6mThbLhNjlgxp4PTERDjyG5C1AkV06epF2s2YqnTPYOssQBP
saylx50LiobaCLT6/LiVYZdjwt1HeRTakqx0ltKJ1cMqQ0ZhNKcwy/wJiz+D
txiCNlo3kfxuLKHBakx2v+qEeKH9dae9BRY0sShxtsjDRahmLiox2uqLQ/Xh
J7/HHkJOCwmH3Og/Gew5dzMfi8r1m/3oRWGJEOJ0+uATF5ubHeCmibcBOR9w
yivl7e1ljRmGUar778I+xNK9Ser5CwqvKEwJYrXgs/uI6PUcmxpOepFhZInA
P64PWUMLhBJWLEVwbWg1vOoULXe5AEc/yveFcj5c5kKMpRcB6bHTIyHgfMpN
cgzeIexhy4M/9EjinD6AnGJXa+wpTYfmMgTxUR5W12GHHoydCGNf015BZduX
FTwglq9Zv3JP2gaGbDMUi5GAjkCiN+wXgpWKph7ElvwxqW0RbB4uK2WncgxA
GvcL4UAu0K7ImJtm4ZrRT0xxkugGlrkP3Gxxk7/7i/QoCGgOFdmhFV3sSYip
oslDQLqHfNc3k/OP61wAcC++QtjJfOrzAtZqvqxH3w5NfasHmBX32qLjtjsB
fovsMyXDRc8GEsSzm2WMER362WwxTpvIuJxSmDa8x6bNpptF7Ltyh1clVlEj
9hneyaxKeUTjqup9IZqpx+15cJhSKUGetjvX66dHP01unUFqJ4TlGIelakeI
d3OUmftSrCsCqCHo0jBpUV2dkFBEMtak2wenN9kk4CjzRIiG9qyRCCsBPFws
GLpNrb5KFW7nHsjYlBv+83PKck3o3w8aic2Pvk2LxbMzxQTO4wHp3MCFbGWI
9QoiU2wOpIb0ma8/Q3/82xnwfAdCHdqokx8wc/9cW+1mkGoOsIq2XxBUbs21
5CrxWbAkivcxd4EjmHs7Z1un8sEC0gbAAiZbzJA2uqX0eNwPP04DS5lQTwkq
fGxfrgZmEhVts46+OUt97+5g4kLWmSRDe7bmkFciw8Z685uEJV9I6R+oqk2S
1gFAMZHaN6NWPGLdC6rBTOncrx2Cb2x9MHacTurmn6pvPfCe39cVlPkK/2xs
KNI7WhHzhJOC7SbO/FWNoIkUq5bbWvL+0SSRXabUYCjfAH9M3zaTL3RXXIpA
AzbcEF+Xy9TzwvkwLqcPCXtZ7ooFkNSr2ZfDF2rqvZwoIAJkqPNGag2+RR63
1pJD73JzN7esYNNpQdEXN/FgiHtpuoMnQGj+SuxlE4BoVJiNyj9o+g/bf3Wz
hLgyRNXN9x3x3abvSCLyHwTm3Kk6Hhcs3L87gmeyBKSsstcDqO8fRDtvn1jW
uXClzZ2BSXczY/GQf1wUQy45+o8EtfCnV8t/rP5NCeZ/hcJL7tLGN1azHLy4
vROmetjsWdErzKbba631KaNIs8Dbt64IkU2Zr19pMKTjtaKWr/odtai9CH8v
D2AOTnMGJPSZcg9RcSXQHQ1KeVb0FrpDw/lR32zuLAWi4+lG7d6ZUWkOmOmj
ZuUK6yKJcgKbhKywNOeTxeIPCEZjr4Kvc8zn9Tl+OQUveVg8nsTY4GARuk51
0JM6VxnWyWp+4T/nP/1UPq6Z7GrTsnRTp1PfmOYkPE00OFXFypAYKOOLqkuE
k66xG6CgZfAbeqajaeLmqOZklQh4WgL2IO0kdolom3a4jnAHJICO9IAIQGBt
aJX/A6ucYTia0TMIw+z6PUm+gV/m3K/sA5B+k8xxCiYaAaqcQG8BU5pWNqit
6I68pKEsb6krtWf1n3BmhQXp+LtCez5vUg51wNcQzQ6FtKv8jOXihqlJ+h29
0Rzu6QC6I1W7IBOg6GjA4x3tU5gM7CRqaylbfLtHWZEiRPMAdOEJG62KiunI
qdVjT2rrCwPzw69DLZUDqaj8n7Fw96VV8hlAO4rEwdB0jjEQ+4sjQJcbmFOV
l+2N8BkqE0X4rbHiM+Eqiuj3kC9lnzdAIQM/lcqcrJbxB7V3D95n8dzy5PKD
TowyYAO7F0sIOBDoCKRpKTOebmVRHc0inCrMTRAjtszWzj6LDGRZIm+N+4oX
SBax0ypZpj1PXu1W3lQVbg1UTjaeVwAugWeF5aTBLOlKZ+GZ63L1z039q0Xy
5R+LmsFr2SmKiw/IOK/nY6tSuQthi4gCYTctPk2YAyQ2PuS5IVk9y5JoCPqO
K7TTxcoYpFshl+YEkTWDxs7cAfFLCzbAHInpFND0M1TZ9KmgWntOw3nfRqhH
w+23VN3k4VZXypsHCGYDzXmW19Z0VCUW+I6+biEuCmOjV7ne7nQN+64tKI5z
RgKQ1MEv3FrwTC0RbTg323AnA8UayU6tRpyBiYkkZZNMXUQv8NHbZHBEvjrK
NBZY/DK47Ttb02U4rPAJHlcUHk9THhAtyQyqE7uit/pOTDNIjuGKtK5WMPsr
1uQ6vYmjirpy7/m9SmpcoEmEMb89oOfeBdSrPN7yReZoIWmmzjASukvfXmZk
SmiUb97FFjm25LEpKg+NbO+UGR2hkcKVyRo1qPgFf6X1TMamy+Kc9fI1s7t0
7ra0kC4J+gTzyIell9Zyrq2hZgv4BPI2KpUq5SCC82l1k64w6BEeQglk6eyx
SxtaqNfsbiIEmntVtPqCHUyGe0RK5CSgX5MFfwExJg1fgnNa4f+JOcdiPDPw
QnhXCEFDcx0SUXcihNjSezk7TiDsC1Vpw+svLS4hjZq3y4vBmHTj3ZFtM62I
CNz7yJFyTdpuwTnQGZbNknJ4oklHTEbc1biKirTre9uhr8/Pq3fWHJoMKidE
UM988gLBYso0HbNp54KyNqOqyEyMQC82Bj8oEWlAvDvqQNymMCtYAF6HSgoZ
UF0bJ2LX/9+b5HdBrnwFYDhAGYVvqRkOmifkiNb4AW0AyyFsJreC3xuBjHnU
tZwsEG+K7STgeTcBxMlq6LRKY4TqU+U3pg9A0xHdcI3KqaVaSfT7RFs77zes
hBM59LX8OEcWG9pWKYJ4P9IDXjViIIXca1DepgF7zQ0Dsw7qOEI1Di0X5UEp
brzisxnt1tTTnyGrNehPH7WW5+cvAVNTYuhjwEo0kufHlD329dIV8CiPJ9I1
qw/QtpAnj7WF+6f4cqJcxNNMS5nDRWb3+nqimmGFG0LBOkHBR0uiMlOhLIZh
mFYCz/lnHmwkMllxxTlGStLrplYiTQPQxr3ddj9YnUhw67lvQFrS/f+CKTsV
3az9ou2ySBa4O4MxKr4elE052U9Y2qs5j6SD/EV4GWr9w3+4AMc14aqa0Jvx
m4TxfUC+VjTvZ9AdM5U492lqDPe+v+R2jMWWS1Tk1UHa8/GcmrGmNL1ykoe5
Q7ANk8+jXnpg3bLplVXgYtVtYVkTxYDEoLetbuiBLR0Hh30pGICViu1v8SJi
C1mDpAYA4HdNXoRuZVJoMB65+rlCySK25GP4qQG5TK5fWmvp2pHTR7mzDEDj
NRDJDOcJ0H+QnvSf+uqT2eG2HVOJTlstRENZ9HEj8m3oVA/qoKiGHjJDnmOK
fhoRbCOXaVS10RjA3FL3ZhdGVpMSRVrhc2KPeKlPNOmoWH13tUZVwU1A1yDj
JeOp2pz/w7ewAiV7H4ywxMZKlsRvSt+mgUPP9r0TXm+u0z2WxeZec6gXRkLt
l67yeCT97NcH2UqA7EScCmc8OAVRfHbmUPo4VJMdPyLXH1eNTK5l5DjdRnV7
xw2I5nVi3xXzgCGJhLHAXrwO/YtPT9ylGbnJNNfDRufIeDEdNvKztHCDl6/t
Bu1+a2msFwSgwDrn16n1Dvdx7dEzRq1IGh5A8YLIm4SsEAdQkncvYGK2TtM2
MJvFeK5h5xsaUWViBfcLJuucFOwjIe54ZLKgRQTFSTGiHTzxHIxpXCNDoMDn
AIncQGHfkmBTw37l5ZkzTRupawnXWR/rsQ4XHrLN2j4SF8TRWfLB7H+67vaC
ZW/UHDUDecWU30cGZxzrV80UicWs6/yG9TLoJe+ZKLtK6IyKTMK88hCwHkUQ
/4+byo/U1Q45cdW+BB5xejUvPvmRFOwxP3dukFAF6BnO2Kd4vQkT/gZxKhbk
JN6uOyktaff+wz2wJAQB97NuxCTuFWGIfqEWA+bRBN/X7kaBj6JStsMSaWTD
QslQOnY4DnVXazAhTVUW9lvCzhfkjXDvbTzqqyu8aEfN/OkpbZMSCM70fPYc
Cj8xWuVxGz/ztaVbOGPk3SXLuSXvBgASxzleKYpU8XEj/vqjjHFbPGFGAZNZ
BNuFyyDjGwUwLQSMKdfJl6D86Eh4qUDafP+zLWOEfE0hpTgYYUi0yyyDGKYt
UxuWV0MqBALx9lr8dXdL4/gzK8127bZkiRdwwFgBTaKvKvNZgNvf6inCY0c1
o7A2eNnXGOd5prWSYtWcYO9hfIDpN+jy4Nwe9gNsgA4PsKMhBLdSAfhPEb0N
tUpkCXZoDIF8Yi6hIr9X46UyFobMJbzOCO6Y0ydvtB3aiH4UoYd/lvaGrzU9
Hz5EI6OLK4vMQdCMIDblWMD1XHX0gMrIQhuCJ0TdpH0A3zsv618B/uG5GBgx
QbPLUfe2WguPNNF6eGjIUVpnaA18dppoYO9U18AGetzINEJlt4I6WV73B1Ol
beF+0UwHdU/w+TmQ7OYhhAeJtjhOOGpwhBDWWol1y5MFjT8DrnWqUINqPMrF
hNEWqQHc5KeGaNK2DzhQotZiqVGujtEU0wccVMq01R56Tz9lEAtUDsS3Ox1e
KDj/coY9R0a35dLlzNCpT0jlIjb3V645vE9sVR5U8jHUCZSYUQC+Uksy1l6T
It1znQLfXZGUSkPPv+dbtxr11kVAY8k6pBR9+LzxzWcrwGYfFTMlNsGkAGar
m8INb9XI0oOosDtY37XYTJ+lTYGn9gqtH5YfkmE25MYyyp71y2oy/wCw+H5M
0n1A7m2b9NfYev47ZUrXEMdBG1g2Q+QgKi/IrxrGUqIW/+Ay7qpFweW1sLPV
iVTjxSSoSqyIUDliKHLyVq8lgiKu2xqAiTOmEQlUZYsCYXIGIofD56JawybM
J4vMcEFcXvLq4lqRkJAzvZ1N4AK+Ac0j4PVPEWKM/B981ICH8ekgFcdo++Uz
e4tbIOl4jVhi90PBoH9xb5x+sDG2/VbJQcpUdiwRRJwZlqPRLwIKSLfDeKKp
0oBTBa5frGHu1JAPgeT6wmYKHynRNbnavRWXLdmif9xU4hrvMgkIbxUv46Kn
7Q/VquKSOw6OSuhxnrK60YYFz7Wji8FvzKja7ORXMhiXEsC9nq/vhNvFxiEy
rSeIwCE/PB0NXTe9PoiOXwTTp8pJ0JNDNophOr2wUYHWd/8F216hqbFZH6bh
m7tQIOg4GyKnMrw5YXcqr8EFdCT3UulFZG4xbLgjIRwA6F9VKTchPRLp6DBS
h92I0SVaC+k00key0mRE4z3bcwG62DYU/IKtcaXOHU4f35XTRGFIIMNxejbc
wYMd7XMFxETcq+oz4TbFzp+8LUKjVJMZrjNX4Aa88fjRhl1Ej1cDsFzCaeyd
IR+l2hN6RfTEoBmSARAv0fco8TVTmVmxIDmxpWpqCgbLvnLo/i9kidlND915
N2w4RpYVx15AS/fo9/ti8hBESPeJ2sKUoTcuIVyBf6JDlQ8o4YNJUsq4Epn9
XuZ20YMzDeO1HNnRGd79Ozmt8dvUWkd8BYfPHdLllk3JmerVLO/LWD1XNqU/
YagV+uhnEznFWrCKst06HFqYct8EPrpJnJri7f1/KND53/Dom4kHOjbVD4xy
CMxHH5Y21SxkjRaBOyoQyXNzSzwwRD8Y/TJf/Hz2Jl6N1enXpXcO/JTKTf9d
lReyj7L9jm8EaHMcpytJX3N52zUzimIxAf0CBYWZpsDqEuAJ+21M91xRICrK
oB3qb954CpXG/qUelelN2UF45rJPrdeqN9h1rCladnvRKcdmnSQMRhJjJMHf
6eRe66IaafVeejmWc3+q+0Oqd3LVumpod6XqJHCaVNt2boDojX4KlXhPgSOk
v4IUcdOgh98NkBKbf/B2biG76CXPmwQN9X6i5yYnL3U4J2wdGIHQ1FlknM59
Ur/C0JU5N0EwE7xSOYqXGF4slMYjCIoGcw52PvKoRkb7IVTpOX7+qEayTk/p
jlffGtmDY2OXpGMywn6W/etF0o65tZ5EczwVQSVFsriI5b3K7Jez4wd0/SUz
qwT4nAsKXG3E0VnONF/sSi7H/gLQUFc6l+t74ZGQeQ3sf/p7aY4spqt6J8Zl
etRVL6T1HSdOAi55qRCxt7MigvRJ/Zngjk9Aogp767hW13P7CUx+LxlV1wXS
aJBjXWu9ygUvmXytZQG4RgODKfk9TV5nhIXDUR3bhgGC2avmTr5ggTJqULIT
f5KLyE/uRW3zIZ4REHTg0JkPRzw4Qe7wqG9trQq57k/m5bIYQIhJtCwsL5vt
P7dzssK5q61zu0rKucG/rN5Gc5BX5LgZN8y01oLcRDcntSAi+3IDief9tvSW
n8Woqp4leYtoZNuTHJxLV8t4lfdw5kSbe8E8UrW5zq6xr3eJGgewvdVJCovS
t0dNH+vmL5GXw8gNo0BvFyMcV33P1UX+tMWzGSbNR92iOBa73kjTMIn41sL5
08oRXBpmJChimDUlz3eTYHRPVfcFUSJYeo5HfZ3zp+sSSJ7uMjp6BOYxZC5K
ATiZXSg25O8vc62lQVopQChRC0NCjX/pbTG9cskNc889ecT8Zt599VcGJI5s
lHAU54eiHf8aakZNNCfo3Jk/URS7L+COji4LsgJmtzBK5lcEAYwXTC0oV3+G
+4hLifMB3mTi2Q9CkJmfFzOqPRmifnJEpJvnb62j5fe5Vrpe+WXHJhbwR3Dm
myhlVPaagcwLWq1HQKoBIbMlXGHdIfA2jmRZ9USswBNtMnBxfXpEDIMhN683
ufrXHpD7FTa1NxMwewHcZ831yq6wHyMPpH0MJfAiCUHi0sr4UKKR0vlINsGf
5EmWJpm6E9ZUcPm/8qYANvVctWuhlxnOCZ23DUTh8zM95GxZAn6UPCplAFGC
0/CPrtvJfuZgsXYaSXhxoOnW7mZ/wncY/g8fxV1iL/TZ8u1S2pyPRstsmcuW
ZGWyAJiccyh5ECK8KDl/UXtIkCNV0i7MdwC91CpzCkpqpCoeXT4Dq/gYpAOe
18Htam4OSoMewaqrIvugCxOVdxg/r7fNdo37W2TJ/CPLPjn/5L7Pdu+YLhf4
g+LTqdIbQlKMSIu6h+hWC+8RnYQALvBLKjwRB6WaLc7eG6uIZ38hbZh/cOeG
oxRm7Cb/0tGUr1w0cIVLM8JjTx/TJKFWRxqLrVbV+FT0Y9y9ykNj+vDVJX0F
aautRv19DqSE2OEEky8192OCHfTDTm0/AIacLp7d3dT4gSyOeUfNzlgekAla
C1fkf1P7P9QTaD3UsgGMLNVPh7L4hLey2zJYR8TH5zMPyRPWrTTUs/IV0Kwu
Yr6LeByiy4NBvK42Lo/cSgCAJGhw4LaZZBUXAAGiLlHElKlBPJrJyqtqIunx
5140g55wL3X5ouwCZcuVnkGE7Ri1xzK25+qEl/pty6w8uLltmug2YaZ5s63C
oXIP+S86rKdQNXgYeY6XN2pCHerW5uFiQx+NzqYuEFlHM5D8BavaRdH5lMny
AsOPdmwxUUBrd6mO7EraxOzBwnG019JUZN02nV5XzZEonRQbYrqoG2tS1KYr
+C1bfrrb50ty54X8+OGF9NPciTeI+1IrZcqWiJ6yQH1QBCBgrejERqm2TvO3
OoMziZnByL6IKqNj6VrG5f+tgQ/Dl4XXcRjPczJBQSQINoM1PoeDnkTWdeW5
GnihNrYPmm/KKABYIci6JSYZcVSMgFUUO4472razO1opVRLJ5uOyoSTbl1/H
9Viu84KqSLDOFmUph75lzgHO3Ucsbkx12ylhhvoztrn3078IBLByjP2Tnu4k
4bBm2Nja6FO2TwM+3omK7wFOIlQ1qcyLn50lqta7Av0FtPdKs9UX4dC11NFz
n3wcZA+blyNIpyk2jYyO6uy6Pp1VA+9x90lQmhXcwWCD5Q/c9BuQ0VrdK1r6
PRrivHaLXzBVb6ZvVIKFxGjbo48dcz14WYkva8c7MFCTyhEMxD63PIJJ6O1f
hNTfi51Mwf1trjPNqhkk52igeaYOiByo6an/qlcnh7x+Zl0BllHPqJEPsWF6
MLt6R4aM6wUGHqDN2NEKWATww+1Ij+Btx76hULNWaJOWR+ONhYQp0yPf6V5b
tX+SzSf3vWGVm7b8gB3Afsi6DtUiAfQmJFF1bobx096u9VzHf4bYNfB2w/oj
HZhCm2bIGs2jLleqVPqKruCZEnOnJWucgr/vnPgsDBe/4glh392tbpPetcJ7
x48xB/UBNTtyim5toUiAjMXVaB4lqfSj0D8VwuJkAh9uQ19R/LT+JL88pM/X
Zy7qpX+fLy00GA5u+0tHFrFvQuPq3BlNHzjmku7AYHiI57SDwQJwHN3zfiO2
5ebaRzdTJn+RLv17ggzc4pFP+VvnsN2zimB733CelyaMpWag+Rs4yo6gtf17
eo98kYF2pyq5MV32AQ368C2Qh+xLIKPX2JOM7ID7jDj7Wa3MgDQLHoNqjupH
6GPJpa1QuGL0Bf5Mh4F7kvFL2zrCRz8tTcDvybnVWrCH52qK8M3DOdeNMnGq
sW/WgrXFstZXAzHzzNQ8/DexDCy9aOFl8PCRUq2iVhhAzDlk2mmjQYuZgZC1
XDWKXUyolQsRdMavfZmJ1V95eNB055QVfD7YHQGhJbP8Dr6Hm8mXijf+ssc+
A7kiIQQSV5hP6S3+F+gOiAP5PuwqBKSxkTRu1PmD2dcI83hO4DhZSK2yluzQ
U+OXZnol/sLJKKpmb2wrBDA2hWLM/CHfjU3t7K8VxRJ389TqaVdzrf2BbqzO
aIQVBvXnTYcrx1HIkKH3chJPACvL/xWpds2bA7UuuRpw3N1NDD1ea8pC91ZM
ZtthUZxT+cCAHEFClffvlj8BEscc3ApMR+djtCvM6kiZcTHUqTbQQlVOzUe/
yN+uJta0gU4lJwn/ML1V8vwKe6b+z/UwOtwk+HTmE59u5xHDhRBLvXMqEOQy
oRe0siVCBKtwn1DspArAfMeJLfUdzGt5amYBTBR9+H/Tqizikjtsr2B2u7dy
Fl4iUeK0CHIV4oX4viDorAyYsJK9egTQYem247roT51QQRD2rM/bHM09IcCG
bBrv0SNFiNBdqDJayOiXL4WzxyILei1wiNQU3EuAx/q/XnyaxLvwO05VqFjo
8QTsdU8Tpf/xLi7fZKPvg6O+iOrNWNgeHVpBeTL1b2JtNP4Mj/GLl5v+yjnV
CoK3B2MP2D4qLlt6G6qF/2ykG0Z2hqdB8NE0UKaRSS7z0ZYf5UAi30idAHBR
cSgaX28RYxDLuldNDtX4ebXM1EhLHC2ibU42Q0Gg0USdNG2DL1/zA4lA/Eur
szKT6gMW2GPe0V9ormEAcWLYUBabw6HHXULRvDRJImAnFJ/RPEay0BNpU/qo
HLKjdAYQKQmL+UKU80Ybn//XZwcKagnfS3YGm5KgLLlzpl2XZP+Gq/Kgp5sv
Rhu7dHd+UxHZtUgdGQXzoHeWrwqNR3vTz0Z9HMi21lqHlnD/eTOtx5VN5ipd
SLP+Tq5nwcEoiGrIDAzZfx3/jEXvCrGcSGH2UBUxVGuhd5MDWfMZOuf9eo+6
4RVFaAbrIWlqYkd/Ph+pG3bjSWH5rcdDSwQDXVfwLezlzYZGJoTLVjttBoJ2
9lfCRoO7fMkJ8HY+6RYIAsnNBLHfnFIdZl5FVO/Gt5lzJMoeduS+ibsTQ1TF
+KvJigcs6NBPcIBI+VchDwfbW8EeGEQwLinLUFuFe40e0Pp+4JBQhGHWocFa
BPps51Xv9RYLqaA5TSjzgUJoz/WVmQNzKIdoiMUHRfdxAIxk1jh63bu8eU4Z
+gni1WkDzgWfKMVL3PO4m/iCodJy0BUW6M5YhsipFZidpBzRBYGIn2UiBB8c
ZKFEEeD1AeDGQkJ596W7EI2mvaEGLCR/nrleOs7AELL47FG/Ksz/AhGaT0Zj
QdlxYcvkR6l6QBdUMjPa6VcLWEgpNi3hriJkJBZkjLM1SPkdPpccG10/oKDi
d146DhAhV8m1YKUQS4Kf1Cwz0ydEvCCQvk/kq8CBhzvCBAXr+cIJfgfukpeD
k3Mn1uPkQjZuH6M1YZ2LKR8SlhWlUJng4GEIDApIu5RAxFPIcjOtqNcvkYgH
Zr+5wLtQW9Y/8Mbd9YwJtXsJcclfdy1oKog6bMQnZRjg3E/S8fgemAxbLmr0
0sEJTuNMhfj0JOOd3A/AWsfPce8XWx49ElkzJpzws0mZfbKTSSKTbF/LfghI
pDLkFqvQFQ/APiTtsxngSwyq+6eWqPZFfXVN727B5v1nHoI6LtyhA+OiD75z
7zcyzo1MfZCj8kCpeOUSUYKr+JN5GG2yhiK+pYZFr9PKk0bXsRsVprVEFu4R
HOABtqfrvZ9z1QjCv/RF6lKnbyj4EB1WUA34/2IRHz1vU+yAbaEUN1ohejEp
ApDW2Q5bSQEuXpxty0sG9ndKSH3pJAH+rPqdZsRmN8OuNWRT7YYSD2uqY856
kOAvrW8LbNelhOlzcmrNwDe0k7hZEpUNgA7686TPxHLx6aRQ8CIRXcDQdIhS
vu2mdcOL0G1XdbtKfXowKLBE+i7nHKocEOE51Z97Wuo3/V0RNImlL7H0RNQI
7Y+lTN6VzL339fBZWJn5N4vjJrk1M+LbtXNyW2XwcBEWuh1hb8sWFiPqyOXt
gp9Qq2IHTHNi0tq1hS1llWy6+ZzxfKtwgJujo7vFTZfpXJQA/k94s2Eswysl
1TfyLDYymKIP33cTMpnvkiY7Zo/FcyPtp+GJWQfoiMihEeZmpttK6yTD1ylB
L7EctjvaUWqqGxN8D2H9/7GJSUzQl99g2OjPo3tf9ozxEcyINOGoRk0DUiUa
I2id9+g41fcwWHp2RwL3+GJ93zqNLxg7nPQqRov/LJMG+fGhUpmoGOuRC5wk
5xGJ+c1EgI9JXd0tUz5y2UpbEk7QDcJj3rzKQxT0iosB1NSJ6pmfkbXOQORr
j5RzLEQ8XH//EDAW5oTyJ+MezmQMvyscvWuaWYM3144wbkUxG0R+nEe6YIf9
w9l9U6ekmRJvb1uj4tqvv4/6mvRNMNqA3xq/ygn9sA4q8WekjVQxqthgNEJ2
bDOQzpqA6UBesBr/pojBDaXwN5MZViRBfwMj9XroPx0fvurkey7uqLjkk4Zp
dkc4aON7tNJrp0izohumvHeCBJXicbyqPvWe4H9kvu6lclckWryl+e6yA4ms
LYPFzFBkPQ7VSp6l5CinqDfDoGo+bnU1xecJh6ZVguXYyGQ/QKWXcuaWnUzM
4fHOlVyzFZskTfIVECcmqjez5WRz7r2fpufj7EhFO4PtPJXuwJsytg1Ml7mi
0Wjo2RkRtjFZlG18X+wJJnMpVJdyAf8qH0BoGE6qJlPBbR12nXULVQtPncXu
zsaT3WoiXoHsPg8KHc+1Vw2OH4JcwUm6EcnPG+MbxZo7iGsaNzMC06vmCd00
bC3m0tSEn19UUWrsyTSi+8xutOoz6JWptZTQ0m1VCj5fab0sgqhIVz9c6F7q
TE0rjsOtlr82DdEIb7WnpVKZNfYDKat5rlTTrOBBGrzLt+WgjZw4/sO98VMp
S2mwPQjViNCallySsljXsUldxovlGbAODSPBGv1+zekepphLlibK5a+HpbzP
bAeL5xIY+yc4l8TR44P1VCK23BFjVfG+/ZP6m6gje9Fvjek/b0S8cfB6e89T
Ig11mQiu3SjDv616+PkRijxAdcyJUvoQYa6kafajBDnv9wbKs7r/Q2wwOb2Q
ouwFQMVbA1QeXvLhRPtbgMxfxbCpak09NR816JNPtN/U8KSdPN14F+5JIN3s
8o5RsgaobHrA6ho+zMUZP67lp1FSa+eyZBS1N3bqlswyOyHuwaHCsqPiuf1M
X9WnT98twvqtdV7yWoXXqK+RZB5dtW8tXa+gpnqqVTjzoDBCeGkw1ALGY7FQ
X0M+qMxiY1Wl9DOZZeap1IlEVhTwUE+pKJDc7tO/942W0KwQM89dWCJL/9NF
Ccf+frrX+58V6IIerJ6UG5A6U7cycRwOjOJt0FJysHkNh1U58eDjfdV7eY4n
8B3lkwZmoCR3UzJuA1gBeIUz0tqAZKxpeHteJm4VOp4wZaLxaiaNcfeYEkiE
mP/M+TeKZ+7kMvtF3odQTry77EuHXooTnYd1esmZowWogIpCwS0M8ivh6BFf
knr9/WYTk3tThbTIjF0Mpdzm0yPgEUQxfKP4V6gRmtxSvj1cmkSW4iurf8Sb
0o3wRhLr5BiMavWZjKKCxS7iuR5dMPJcsG/Qr3XVlZTr2ka4BaxG+a4e76zM
/o8nz71exKMtqRXIVr/I5GS17Kn6OatiPS+pRxdunHx1YAoj2CzPE+s3/NRb
lXCskXeeUY2+puqwwO9YX/m1CX1+20y+c6hJ1M+kHaRbBC72Rg4+3qroDO/s
3VbIkQSCG2F5yQF88I/v00jEZ6Bqk1thgDN/TdeBAdOcjcNkfvY3UX7RXkP/
RE5TCnniwa9rOodCGK1wzgCrxol83O7jOKqkhKeyHZrdkpsKMtiDt83MNwUs
6SL/iytsJqEAqkDA7Pulc07QPsR9FeCagW2E8D44bxExmmAjlRzzKjCU+8q7
4N6VbyiWP0n7AgsM92e7s9PjA7aLrxVHUt4pPnJuaukhDy9q8Uhciql+GtcF
YFHcMMEjm14Sr1dnYk/qa3qp49YrhY/liRmMIX+pgXAZeSb/74RUnGMVt+5a
/YRzn6TUoZE+oXLaEc+q7Zrs4RJFXm+SHxHnntg0KkeTj/ec3lEGXoYGjGT4
G4ZlKTQ3tJZPXUAKxUCVkt4bF4YfrbPVwj6Tq2m4u3CPbdU2IjZKEsJFuYC/
6Sc1MMMxu/nuzvOsK3OEezP6QqocHG2MIHKJIYsf03O3mUP2RVpoiOVh6X5T
nxEsi882I4fRAxrT8PfWk8P5w1yPNDNk0v1w3kl1D8mTvTpjr92yfthEhJ9m
4ntUk756PPkqDdgG0RF3ntfSDNGD3t0C6b3nZE5BxDKCA/3KOqM5Qv14M8PF
6xtQBhNVzQ2qjvnmR0cSTsq+aGcPy5Js5SBSch3JC7ozfAB8a1OU4IuFFaaI
TDCnMT/tRThY2dY8gXPY6gJJWFxC9jTt1vjId2lJkl8UkHNaa1Ow1pHdGlwe
s2uD2P9TdARG4PmaCCe/A083DYQVFfbR8cngWf/0vcD4B3g7Y5YKCzESmxcu
S9+q/7/JQDcZXeUIBoxDCzOMJ3+Z0ussWD3qNRtVuk9QbHTINAX+Bq2sgVSW
nn4IdeX15l+ICGBUlFi5MwXbCd2emK5M47FYMqquRh30cYDbbLf15ilJ0v6Q
KxsriRMmnroUVvBoUqBcFyIP9noEUG83hT82LXNp4rykymWGs6iCzQsC24oe
+D3559+BTNqxbxmFKBkfZ2vwb8PKf2WXP57lw6Q4i9JaVVdN+EUPW4y4PKw7
L1VAkS0l6ZQu/C/R9SxqNSXtnN2ExaanPhfiFfMWR5+/XFDznVEdYZdMxH0f
DZRkS4rszlz4zI9mHuHr8Shuhh67rYsgY5lZX6DhZRpZEjpUD5b/RZauOfwW
T75nZIdvOVos89+jqXjkWjRi/WWkIN8fyfu0qXLC2S5ZTHAC+I685AEc3GAF
/YxVpAMcAPxVl0nfQAf/nxyXOISS63rZBy6sNof8vhZywhv8HWG5ukHV/oQL
0MV1i/isWPF0hdxEcok2SbPBh+79ybyrsaW+p3aTCRZvJ6rXZL73Zi1vZ/Q6
jBRRM6LBiDTqgJ9eE+zbyJwzYpUGSZ+slbU6JrXlPoamc3Gw9JcMpPZOnVQz
bK0iwQJROFYqMGoqbJphSJlgNmqPytksu9T7UAOYp6O9LSCVpu5SeL/hFtbg
KuSRGm+8XUCczCAYVnEPdi0/sniMsE0hrdY5ABA0gIKHOmk1El2IyxqwiPzp
8DfGVZ48CT17QuUPQY0065I+X5WzqxnXxVVjr/nsNBjkK1puiWf9Se2JncDi
oi3BHnsyjGA3SmmgbaNxkWk6GxxSTqPi5OlQ8mXjMsw7QAr8aHkYmaeEobuw
3GXzfNaeYEW7FsE66DRMW2xmI70bH9uBUg4V8AinJlFX54AP9jY86RULGieP
+T2i2f/ys0nb1R4g3JcKCOmFUb+ThuP/ndnQzmTVcioZmTtWDca1yXhfMVc6
780GT/M9LCTZwnWLsiSsBZIjqcmhGmTpaMehrDP6BOKtWss60XGYWEtsNt9g
G+iD08pAS4tfGt6FFc76lSJOrn+Dt1rrh2plSvvLXz9XrT07ePe8A+06N5w1
VoAnm6paT0CLpiz19dLhRFBeBgGX9QQdWhlqMnvAzlpSmCOn7Kc5NLaRj9IZ
BXFdZASufafJbzgrCEd403xmwUQvy8LX+rU+R92vClPxp3BdL/J84RytarVS
LQWnGXlrpcgqgmaWzw0wV5x5PYRIUfq9WxnpB7ke7YBfyPNj2pAA4Ee48luY
XcRLQCTXTFmvpfmjv24zrRIlshLQSQyH6NV7On2wdcTnK2+Cs4mqgx5ZFRHO
nCalAlzhELCIU0jRumTY9ZiEVB1iT1roBikTQixddJitwMW/VRln/KksScQd
DLvIRHqDFjwCIDTY4DUrCCRxmVIr8nLMYtElzLofW3uvrP9ycq8aL8Z9mh7+
mb0LV7WPUpW7Zdy3f/Jhu3CD/6O81mcTOJRa56ZGmTWoGxo6rSgbeGuLjRuD
zXUqVc6aITHTt7dn++fexjczYmIGs7RmxTQvk+GNHcLJUvGZmDkIySP7X4QA
BZVyZ+moOKYT79jXJy0oDI0vtaJ8gFnlatuRNWAAQXoVdOUPOCBIPCjbJULI
dZw8nfZ7i3rYBYxvaX7zUy9LHdIO2UCANtVxqYgF7ZEaQMr/s5+TcX6aOO/F
75EiWwYjTNeauEYkSbvx2NcSWIZNf0oTyhj+/wRi+uf0GP++yQJDBOthJrgb
wezCbPr1hXYXJ/fVPnwo9Wl5NX9ngS3h6QcTZRdVATnxts2AD2VoLy7rgsD4
sw/WJ85CczQ36JQtBlp3wl/9DU19VRUrKS+MtWAaJy+u5TGuic9VLPBA5KbL
q3FaJkk+kr3KyBLG/0gvRJUM2VSkfPCdh1xaypUtmoMZg6BpuxhPIrwsWdKV
FKtdgS86PVJZeOqy5SfRfHyhIUTVId5Sq9Pb7Is9YeWmcuZfJ0zgPnZQaNxa
73xpSkRnEqfwnNRJrkFI7xmF01Brcyj8nvmFyb+KHR6XGLTd4DdthN8eDT1T
u5srl7/p87bNUUddnIbXwVlIZUaqYikJ/bJPAiuuIP/i9oVmdRKlEcDW2Nkb
gCDERgsh+vlAywA1T0E3GQFRpejrIMS/02K9/gR/aR6aFNmWJt2m1u5s7gdi
mTppKvjcdIqszVL/OyWa/r2GJ/XBffJip2x8JanWobG8i7iWoSWhSCEFpOiK
2Zl+fCw+Sh11bHhI2CcdcgnG1yEYBT0I5zNeT9Vrh8c4lwQclXDId6+JZYD5
9/dS1FzI0cFKGeVMCSS5yREXpcmm0sV5JhyXM8iFpdyEc4bn5t/ftYI61mus
ZMcQwvr0WBeRZUh3E04+sP90b9lHXXQdCswAU4A4IAE5uoD3mQ3BHyfZLKEs
MLw6TUZBjPLbVrJaLqeVcIJ3EqGgUoukIws52g8hzgaq+I6rTLZtKSEhBroO
KjT4udMrbLyy8JO1L3+ZOZS8/UXAoYlT681/MDPEuNoU5OA4hwR5S9Qty67j
NPs7lSkdwl+rAHJpx+Xr6/RYbJ58fCLmSsGVyQh8YYz/e2yUvAvkzUpouMup
SNRhmOhYRsVbr2MMQ9ZJ1pOQMxrpq00kmIf1G3XQC1E+SFrdYqJkrS7qDuUB
28fxFrGRw+Ik+kL1KW7E/g5lPr4whLfmrDB3rSrlo1x/2aJP3+4OSkvTTyBp
H1ZGBMyhXgFmq1Y85vr8c3jR+CIezqnGB/TiZ0OTTbpOdZ0WCw805zQwCIW8
c7hJk6iG726pWMalJPDtxp4u02Qp41+f0qxURh+HfZm0mAQrj/NMrp2h+Z/Q
enMH9znnjy1Drjhm/M8CrCyv5ESdzcmdgN5mK35LC6aVPE2V7OQRH0RCZJUU
9ElciC2Y6VVTfSKNO4e4R5cXgSvlHWf0KctU8+l7+SSqcr4dUK77cmO3L7hv
o7ISZgY/7Yf8y+NSzi9rw/tlqa85bVEI/pW2rtcIwfthfheautkSpgdnn0G7
Shgk9TZUOP0IukhHj1n5jv3ycLjyaFuogB50Dc47iJIM5RSzZzkDsHLzSb2D
dQKsAzDuUDeRqJObn/x2HsGAqDbWgIG9WTF3cosHiJVzJD/r9AOlWr5Df/H1
Yl1LP/TY/uuyDtzwMraC4sk/RWLqr/+UI04tVHYfkGb6PJ0DL6igmQI1OgsU
Jc0EkqXQForY9Ckz5x3Lq1qSXVHSiSGbtU5myS+cgIKVME3Gr/FyZmPFUnZD
GxiHLtQ97tzkJOpu0yo9cTpRtAIkNYjz0vn1ajwLuO6DeVcHXjYEpGwT+Tu6
OoCjV+AGfeJZ4nzTsFThdX+WmQCd3hlWzlT8vRwq3d0HwVcRUKy3EBVie/kt
1ya/Fx6Nr/fTAXoZk8OcVpt4+4+isdFf6+AZTK77LNclJw/iqDhs/TRcd3ZZ
Apk4/gZmv429tf73udD5iv9cpTGH7nfaXO8E+GyD7bYF1Q9hOMH7HY/dghEV
vFRYzQm0rOTUNICNNUGDr0m977WWoJT3zX5O9tcHKgzGjL6/x2RzBwSFHzDi
jeJlEwFV6ss1aUMewLSTkQGNrRBvP827/MQUrwbGaA+Jy6XqFUDVLQzg/t4X
ezn1dovfT9FL3kukJUo90c/PnApxDRBZITWD0HZ+BGxeJ98uFXOK/5SW5rEJ
pLjzLcrofeAhj0gBRNE8rkxHtOLN2NZFRQUZR2paDzlQO0DnqZtSmofjtu1E
FIzwTiJiJLQP7rmvyVdIRSHZtA13+IyMactbT/5w7G7NUoBiDtvne3BneleX
56gxI6i1s2QW2deg1fLsGd0VLCVNxXp2rG9tJVbvmmvXV3AXgySHWVUGLeZD
aIpMhrANe9j82EtwpDW89Sbom/r9je2XfWFYYk3yXzTCaaJx3rWfYOHp0ISR
9GI4WWHan7n9wojOFnu0RG0/n5l+N0AtsjucJ0//hKuZyxNs1ofyrrgJOF4Y
1GLURXsAt0XL4lhVs3dQ6kSokKNG/jZO0h6fGF7BNuWAiiR/M2FghzcsDaNO
bTcRaKcJL4A8m0u/v3xc2VpObFL8u5nFpyo8GS92lURAQOZrvCxV1mBYh0I5
pB08xKLeG/Wo+r+TMosye5WHoQKYcZqkynCyJu0vOjq4OKa3jMHCEcounqfN
uKxRLmKLskigMKvTtN+2iB6NGzdmQ0uLO+6DrY0X/iyNT4g6PWyENoya7v3/
3z7c417vGOmIvCcfc/662kPsHLcnFV5OO4rKd8WMfm1PpMrxAk/3zadFTS3z
HOizsXRMKHzgH+t6asUunQbHMbtNV2i7dcHB9ydHH2TV3NB87dcdEj5FogvI
pMELTzgMeSPjS2ReeIs91cf84Zy9TmLVzb8tIaEWOfJoljAMG6etfJslGfpP
BF6ecdOBKLlVdaf1L/GNiGAwlYsk4ICC5/sNzbYUym8LU9ZFT5kNDPnHug2w
E6+rs9z2W7TNLXomSqZMCd9KmCai/BVmDIGbPXR6n6AajNdgCdsWKpw3OAkH
uoD8hs8SObVpQbzBDjkQGNNR4N/HzfIv8yCOHLaFNuHTwi82AmKXN7okXEwI
GWLC+tLR+UNRQOauqZASjDxdTBCjZHL/aPS3wcffRM7pF7+9N6BxD1j0y920
9+tc6QBCC5YlTQpXh3lmOJmqmHD+pWX4R34EdRkCtZiQGjbaHjZ9XxiClsig
/oXr4ZumCpc8eue2wruDtCIfS5J6BHr3PVQsh08nn/j4vajpI7g+docEcCr7
7kAzvG9IaTmezlkn/mAvSrfhsXoVIghNIdDYyZWvtTeptk4h3v+54bTc2Org
6hTlxJpv0UvxtkU+o4B22dmr/xJghpNAYfunKh/7Q0OZbTovMLRsiFTeamit
KJmB/XoHc6zUT01WclmF+3c66F1l64p4UZ2Fjf+f5j5+1l9pncbWC+J7Wz6+
l5zXjcOnDbcmicBk8j3ZmrcWIhgaavLTHEBp/p1lkDaPT1Rjs9aeFZ+TTJMC
cJSaim8x0sgkN3ir9DCOUeuFimHJQ1jxKd0L21BIs64udDe4CdVtW+yb6Qwp
vO50+ytuW3ioChSC8saPJgLjE1bG33DGzAjUKnR+zFdS7sOwrGe7pwvWHI7y
cmT8WQYne/5GXg7M7LdoHwemEqw0k45fOJ0eGdaxQXXPmOyGeY4ac8iDdwjv
CXM1zBH98nB6xlT135xFwbC6kbaIWX2FwBsFz6t2FEHkhVJ1sTejqsPeK57Q
X+BrIPhU6ZKL2dA7/1eiFBZMf2TU6SPQSiEzqtDL4B7FseaPGGnga3h1apU8
xQ5iNX/qSoY6EJ0S7BkBHFawDvAnj536KGkSdBFi7RLFRxwNte87l4D7vB6g
AUcHC82sps/pg5dcdRoEr9zd+uXjR0c4eI2i/zPFRQikIzKma/Bhhp3cXqHO
RajIRQ39ykxQrNekvQsIcen1QY/Kk455NyjPq7Xl5i1oGq2ccTlaRRaxRrtU
o4maiG+iUcKNL2ZRutXe/sDfdXib7WL0oM56TDkY5rQeDzZcy+9LnOLo1OcI
6P3+MufLAl9faqJ6mY/xnQ401ZcyWAuVdLsjWWLV0hKzEoruiVtm9bG+8nWe
1jvdMHCa/lEeMJSSCHkBg0YVwqTVsIy+Z/0y0dLKekeZbrd4hNPMEuqT7vL1
zY2XCnm3OjD5Ef3viCOV9UMIENKaSr8IsalQCVpgJN37AdfNr6NcrOp56djn
mPFDWobL0/47F1w7vMtO7RQ02j6+Vwq21lCyK0hTqOiyXZFWpIWS4hb+nhEc
rMiVKAVeAdGpYNmye+pPkDRhI4t8TZ8A6CAdKew33OogxUEJaKQ3XGjDv50X
6TSp+bUzfJUodp+WbpAYLPFu+6p7NPKvTWa+n8gnIqDxJ1eQHRNctcI4s2g2
+KCleYexUSBGIY8tz4xaypWUAHGJ7FBWJyu7AMlO+qbypJ2L9/KbyKMwj9zL
y4GY47XDlPiGVIglmDt5pshulzfHB8xkPa2AoWpj94FkEE3Qsj4G8+OMGqAn
wdBBeFVZVDugmjQ+kVD3o0a0DiGEs/WtHS9E1JWjQ1PSqkLT+uUJDDW8RytT
iG3m7sWdkB4l3NWyRA7/LCy156HHrDNmRZdXlFmA/4wO9RHchswi4qENBtdv
evya0NrLSKNfn3dsb0Tdec6gWoql7jAtUy8cFUqoYXsnG2BT6Gkm2AGNJ2TS
7vuWnjj1xFBwszCAYF/qRDFJSVuuwALsM1DYBShhbo5JtrHRTLCaCpETqPY6
PfMQQa6SdNHn6TYRiaM+R/qtKYoC6XHElkc3RDzM8HhGiG3goBt6kdk96+2J
CWkQKd4K/RmQRZqK/Czosjr60ckIy/Ex82uKnbvVTNSrUoAAM8trvD5ZLB33
1tKtaaAMRXMORyOVqjoTT34b43WniBdHc4lwF1D9H1JxoGK1RSWcZEWye2wi
pFHEmJGBz7WRF4Kqu3IcaoBkyi+cOpF+MefTN4o7J1i15zybVAg2FJB/q/Vv
b0jv+DgvrZcKlmKu6tc7s0VH4I90CncAxpGL4A5LWhOB1xdiJF6EZFut6Blm
dxCrLmCWX8GPpG7a7rE9l30q1CCR0DJRc6vZL1Hc6HnxZ2pV+v6FPeTZHuwh
iuM2qvCVrMUvSrPa0l7d6pbP6WPoKzNuzInqqlXHb0Nd9ir4IukSQ4KDngKp
35fMaa8YPVQ28P2eld6j/B5XneURwxKAXzOYMUDlyd4v+Lf/EsR68/ri5ZDO
a9T2bEqbn5IP5UjRyTCV44DOtEKuXb/fZ/5SlnbP3l/w/tdTctlRFKsSOleL
fkV1KxBguFCqdDwae654YJpRTwU5nWYUmMBs0ZSDHY3jAWLkuVF/rq8JXu3o
eBTb8h6WxGlACPjbv/fOqHmRV7wgwdpcJ8qjS0eICoU9XgdL9xztS2jdiiPQ
WnUlsOJ4At64Dj8jrw02ZQ8ya9UyAsV2CqLnq7+4nTiPK8MBIYL7Txbxakh3
lRaokhQ9J9LYUbyjYM2TAC28/tN+474jR9p5tcEXRWBy7fb+of4TlfMjahqQ
bkY0Ej/qQD9jpEz3yg8XvLUyDWDTYTSjGEIZqHwm2EaHhPVqebnn1GU9ROSl
n0Gvk2ym3IfnKxTCGwhNV2vRNicxVssdorHhXqb+iUvYQ8z6VjFgLIpcHMBr
t7cyqiCU+/RfwlcHrvxYO/9oYIPV+JDThg9hh1eM2kXfSMUu5CeAOGoKR2QL
24quZtRXFAn0JdePYqdzrvayDZNX4rfHvc11C15XSKyufWeeJoUPrt+z5dW5
Px7Tt5SN1exQ3g9YrMoGvt1Uy9kHJRGksYxzERAqz1YAc4TtzZ0yc2UecmhV
xCRrk0xPm3FpOVZeo5nzsHAH++Ea2Ro90ZmHfKnveKozC9E1Z7heOT+yPB/N
hbov+e82lEyECF/tPy2FChN41X5gK052n7r53LpOqWRBJRfxMPdfW+T6u/45
XZU7n7VfmADLSP9x++zkJ/9BXfkoOen5wv8BGH2bAI7lOdBKn5wK9UXIjh0I
qdeKD9hIwockkAF8d8a5wuQWji8oXSerP1hD/H/8uXKswQea0dzeBZNJ02oH
YSx1qrU+CGScCHI/wkC41SoEYcAJqQ3P3QrEaqs/gwlLXVk6Fe3siEa1L3jx
NHoEdccQCXA6XLjW99a0uaNZuRF+/fnP0WGlWIDzHTfdSi1YXvOqZ9mDOxXE
aHDogFPyQscTjBj9E+wkhLNpWZrqvFTQOyMoShHSIfWPSn8RPCoIOonWUmgK
X96M3LgUXh2edSsVzwyJoTXczXMIMeDIIDSsJckOxJ/mv0kklgB5A1fys59c
bMSaglerTAOEBYdkAGU7AABtbyi4pq3Thfi5hUfWDKcAfwjN5hRmvolZYPbY
gxw2ysctViLliymSG+hALEvJjk0rcLNJMhpIPuDqxqvvlXMkwEBS2cFcD79H
DzZNKU9CiV0WM8idvWx+SHxZWwBATfwR5lLW55v37+63dDkqbmCkbDd/SACS
zIXbYpcWxFm7XBm0gXn65MaP6lx1pwDxJo8lfyUuRRTEhC9z/+T2x8xBtzZN
fisJ6OVR0p22GuwJd1cswXdS/A4eWXwYcmvduSpqEMZrO+g/59HGuHuRiT1l
Zc0Mot1of3jKGiV9/nK9J7TgzdogDdVePGrzr3CxBMjxXBGKlktTTwH1XNLc
XtVgQuUBKOVBDLLmEiH3aCXxq4Bn+6p8DgbrmOkvid+8Mzxra+4VA7/baWAU
+tNDnJa7Z6JjXl8rbqnl2GKAHw7mZY9RQ7F60oMT9/Fa9cd7MnaXEm8KSFUx
LgWUF2sdRZJ4iFxqGhkGL53GyyMA/FoekEa0XQnOyZg3gHoWyB3kJdOG4h5c
qQr/8dfazKkTTDWzsaFFmV79t3CuE+fNevDIuSKiG7h7J2P5H5HVssPWcYgM
K7dKOwMlllqW7tQBXMs6Kvra/cYOawtAkt93iwBN4TK9fJRBl5N0wcAQuqv+
cwLXNOYX0IQNMzndj/zJ0Bzu+noIZcd/otKF2zJ5o6xFwQqhyXMZoH5xlVLR
eu3+w6U4+19mxaEHqykLL4bEr9K0xijE83MSJOVQNmv5SHhITpWRC6be4Ngp
BMEcdFmEsLCuM8YZ5UMuC8uvVEPWoG3X/66kBc/uzUZ+0dH/WQq9IH1hrPNY
w0KVWpx2u38W3gXiJe0S+Sox6q0j3Cr7F94WRRNrqf2/t9F+FgJKOzxXgQCo
ooIQRJ8+/E10x/MeDgSdpS8uOLyDWNUebDsIT0PkY5PdWkmzIgSNAWT3MvQO
46eH55o9gmSsKtAVNCQRmSEpNKYkjRj/MYLlPiYc+krOpU3r+3/Rj8jHGpFN
xJUA2gxWsSATpoukOllWjfwIJs1pRhWUiBACQ25EjQsqsx4sXg0juJctVEDc
9aPPqosu+v+pZ4JZhpJvz1zkluC18327l8ncCmRgE1RqhAUtSaGirdNfwKJa
SSAn4QGEeQluu/Kw9cLo39zv07HHmb8QeUD8KP5+wGdb7DI5mlNE4DSxUglO
fG6azYYsesuHNsGy1Z8pcPYRme4CjQExtdex7zUi+VVSJ9Wyuggc3ThiHo5F
EDXNR0Elm3JolKdRNJbGl4AyRsqKdWhswrg0mOlRP6Q34vV33SsMY3moC5on
rMSm9PRSn4Ijje49ZMx+Gn2xjn4Y9J4rsCWRJebboaNldJiwwoaaY4CqW8JG
lSlkIQ5kpKtxUxbbLfBOUollOBgQPY8YkqNNSllgPrLPdLIaZDlgkIUfsQY3
Ky5OW3SD3q8pFGsWqTNSrya1XDzloUeyDp7obj3dL9vDPYnqhcbY1ucbD1QL
iPgkQudStFu+LYamp6TdzJH5Qanqar81DVimjHutKjTb+60aY+hMJZpfrh3j
8EB9So2a4+5sFy45D3QCAXMz05wfiUGWblMLeYacD0dZCmN8jwB+p0keLCMB
YGITVrNMjz8MiRnzhQPPfeRtabITom1kEnao4R9Wp1A7avw8aPb4SzTymaQi
ExqMRdkGXFuEBW3i/5LYz5THnCWUvw1LqMxCmdmW9ZxJHkImlVMiOG6R2MPb
iWXtZ+ZPpEkr9bOVrMmkU09cR67IgHc2kERFl+h+Bgph7grvxPLr8jhnVmwr
/qDm8HCb/mNSm0ezsTU4TXC/hCmGnjt2E1cj5DTGL5yiaYgp6qBKjZL1rKsc
h70QQ+3cJ095psUlXB492TMowmH2DK8+VPd9uI+EU1Yfc8Ed39zW8p1F7gPd
OQBdbyPQBc2VUBr6e6ajCawL49lnwIxv+DsufhqFzQoc5dm5RBElRe6NMDf6
FAsz3CkO/V/2gFkD5/HA12owkEqSIG/5G5aYut0L0g6/0hPMXo0uiEfp9eEk
llJlXfFsC7c2Cw6zUCvbgxH9ZGwRayXGqJ6AFMcNyOaVpPPjIiRuzcC8pQ/N
9fr74QDCX8u96Hz+XltWvNYPzJyLN9ev8KC49FbGRJvLLK9DuGXAa1MV8O7L
KSJ5OQux6UrkLQUXMqlKMtSPVh4IepFTeE5D3BuIAHkIKPN/C3M9qW3isai7
9QBCVT8Ox+O/ot40RaE/Nwii8/Or7FoyLlIki1gPguAS6O7HvbIOhqLgstsJ
SfpPEfW25J5GaQG4Pne2uSAML1z3BRDKzy3/gkvQ0OuzzXG5FTH/aWkr1+m6
UuU4l224s13XJh8gpxlCJTduUvdcXMsI5fZOALzAW2oXzMMIzh73vIZI5B42
8j4Uw436in5R7YcOrsrf2LJofNYt0Q6VHlcuqb3FL2qrRAiGVz1y5JZgH5uN
lqc+x7w/2m7/6s1bnjFK+F0QOneqsr+u2al+X1gUDX2P8HYo+cAWnq0iXs3K
J1LGLptSoXFEUEy1ZTd4gIkYX4zxiywpMxLtWFgQfHpIluYcp/BhLkPV/hy/
WUyXeXrr/kFajP/iXl+PY3PcwQPgJWujqaj9RVvRkA/z1jGn9FBwiWFXTaLm
vLO6HBVriXhmzq3tIS3qo/vryPMl6pabHE3yAJheJtMc55PfPPJL3W726k53
Aw+Td4hw1iqTzcCybBTensHcZIX9uq++qXEBhS+3Fqk5hRWIaAxlgit0ZCQS
9GVj0DCC2ELXEFde7N3BlWlPc9cRPfjQDyHqeGLx9Vj4VaBjemd3qlA0GTzA
pV4Qch+EKMprzXsPcJy8p2menJ5/LifVL1osACnlkchlFbJu6che9quEwcO3
aRGXQYPO0zpqoEpdBIc/dxYQUWn7TRJQOiSH4M4CEEyZyxKkunnsaxWobz9H
dHXrlNjHOJeEj1bt3YWozbivO8mUQBaRk5VeqRtKinUc/GaBgMOAcHPww+Bi
wX4a2MZUNA8V30RIl75b+Cuqs3j1Djcc8oAg+O4S5ZXUh43FA0f5JgLGrCI5
Ci34xohDs6HW3ne9o75O0cD58rS80OGs2aq17PM+nl8rSmKxevsFLCAM/XaS
ee2dlv0lI7JFlla9xvQn0/brd+xj3Htq+vUeYXUVu8ESxBox9RWA7XN+hTEz
F8XKcvIoy+VZfyhlGfuLTTVy9mNzHmNAl+leShMXT9qi5b0u1calKlrv7AJz
CFyvltP2rffNIadd1ScCa+RlsIYJ095vvpLo4OtIDtnN1eckUYF4y8UyjixU
2HRIrsFoRJew6Db+tUvf8vDwHqfdzh4k18ysD1mpa5/YpGguKo0ymCI4BCtA
yRPtOEFT4H70sn8OTq8DhfVkfQVIK1W4RpduVdvTpO/wDxJv4LgQgiza9D/x
LSE1Jmr6hyVtKkJR7lDbuwQW9Zd0Q0PewgOB/QJXR9PSwAMq0lUpwqaEhCK0
FxtcmU8oamKHVGg/anSGzPVnD78Un5iuYq7rsuq4o3Reff8lh3APfnNUvdoQ
MiCj2XRGACgA46XJQqQRERVwYJjbPpWzIy75CitKVKSPpIdsRaxXApRM86IM
l4zfSrqnPemjko4fYigMduw5sTdLWfLQs3l3//atcKvkxyMwvZuQPX6xzucp
7BlOKqJT3IPbUDPiW9mahmmutaYOOar1jeevRdm+zoLngHWYgRBKZc1wVesp
aSERkeo6uckIhi8OyGr+hDiU7vd98OAt1dY4of2ramiF7g7imCfl4ClWwwPA
XGWINbfEmYvHfErKdmiScxVWRxV6vahk6NddKjREQaeQjd8dWuNflo4NOXyL
oVfCfovsqOotxkYEI+VqL5zi6bo23fum3PNyqmWEpIOtzWXMfcxdHg1sunCn
B+f7J2SEz3LbNAeXJ4sPfW6SjHKxBSFV7gnqlI3wCFJmOrY0u32RdaW2pIuE
D+rnbWoch2bzrO2r+QdY2GURKoNyYMFTLXrqUTz2yeHNlmYSCw8oQyQcSaYt
rKZmL4DIK3xfgzE/fpgLGTrEPn660I4b4LqJJ0jDXaXAtkbHtPez0hl1n3oy
wdOn2Vf40PDgWHq9qX49NTTrToag/PslLenmP9flXKmtUC1+1j9U+sGAxK8Q
0X+Nq7D4/wwgTQZnI5+xbebAjRmTlFGfg23NfiSq88F/ZjI8zaSzRp1JHNGf
rE8movvLv+RRxL8bD1PZ+0mBfosU0aUI9FD4eKMhKWzDxrzSdhyvyoW1fJu7
aM8IJ3cVjqHF4/3mVd2mPiGJ4HSEL2qdTZehWF0vaR/hcwAZPKFcqJNzeBzq
f689hcnL1x61qeIee/bjCBtC8sHQVXCXgucx5oUBYeBRqsWIjly2ABjOucvD
nE0wJgDAtQUp199ic5KhQzx/P81uYOVJYsfL1scX4pINBTjjBTB723EdGyxD
7OwadYLwtiykOjZmkWc96GdMN0C42/ucSzAbsxzQ7qfd5j2JmjSqBsk7Crqy
OtjqEhRhpsNA3FG8qpRUT6Cs0A3GWstVOcRohI1bjikbHtgefpQRP8HHDHQh
sDhMO+dXttt64521SeeH6n9Zycuj6UkDlk5IzFSpHRS7x0XDTZkVC057Xf0g
1ghk+yaKq8TwYlYhYNza2KL5hdKt+HQng5k2puy3cFGatU/jIz38ASP4IlI+
bCL7xSiUjMQcEfyUkg27omLaXN4SQGKjj8595BvdIFx6Nmm55bgwH/kIVqHe
R+2rB3whdK8YkFb/fI4WI558In/9B00/+5y7B+RJELwN5gmkrUaikKWKe5LP
EKkqGJRZWwizCpWv0FLoVlUiUI38j1JojeP2TSbsZ9dfeeq78qPMfMXQedWy
N5ejXuKb/vIbNLV7tZSMBZpimDHf4Rn5E+Y06R2OkjvcGeNcTZllvQ51spF9
8eeWq5isSyeiUe4SIghq2bUkLYd+3/kY2fqCF4dPA9KaPHd4zXNwDKGIWtnl
V/wQVTmMxwwxnHSUs7rRA40/h+fjm6elm9wyxDnjvKi0pknqezngnu8qmopT
smQLrcoyVX3CM6e5VLLZdwhAEWZyuNEdeopCyZ0fQhtCrA3Yb+ayGLd65eOw
phhmYZs3yxg3Scg+W7GMdYiK1MqFSRhUwBbZ6otalnVlhAg9BZwG/unlKpmx
AKt8j33q9ELH45PYHuLDQrA45hybtnO4f7R9trSz9X+yNYMc3cATt+Yzt4rb
8b7X5B3M1rgUqWiM8E62KZCLK/Hxp4iuW2OhZIP0JV9bsIyqFItaZYwSR3sN
eplPzROHFJcHqXcFN4JHcFF61T3r6rT+od5a/gSy4He93L5frHg5BkcMw3Ox
1ARh5/2woq0C3kPZoRgd298QSDiZvNkU540i7S+GNPABt/Y/hOzT2PJZW2Ss
4cdjzTYSfBQg/Nky32nRRpuB5Qa39dX1d+qfeeu97GpjHcMXgQ4EsNS/839J
Q+TuTQdTV4SHU48Sg2hfn0Cy+GQZDNcm7pIzJ3pNhUpR9KykuWQqGCtkaua5
i9d0d2iEtpzaR8uKGQwmAfGyuFks5xDFb7JfHMJeuEqGlDQe8xSg3BvHOAXZ
ynX8TSo3mzWJ4Jvwxx37+cbDARN+Rv5MlsScqsrz4I85IBTfdh1UEsmCBKVc
B+rWp/+EZzlhcuiWBgG/FfHpJljEHpSeTkAGZ6JrpFLt9jqs8XE5QK4uZLo3
ARWuOm4r3f0i4DsXZd6TphJOzyWba2jqRU8QVLbkmfZ5+Jx4/Y15P0dp3irP
uVo3t8aB4mfRnhy8GVRG6K2R+WHPRqHgpJ9i0aqTG61034r9iadvKr/PAEwg
ZYCcHLIMGwqNThEYq20kBZAblzcNtCE68g0CoNe9oML03pOH969/k6jURCST
JerMBOlkR/YnmNXBwMvXxxfaa521dJVNYgd9EQA8eXAun4CFWhwT6LmNXte0
/5AyCMraug63wJO9Qx4obgDtr3orZfHcbVcJnFhPXs93dx8xt3J8gXiV/wxI
kB5HLjgdlwnb0Mh2MMFxVQ1XML0MnR6g8e+01zAEKfY67+gx/aT8P1tBY9LQ
u+QmAx6x2vIBr9Sn0RmZ/ifI35zArMIF3SB8svnjzFewDn0aSh6Prf4wVfNN
BHxNVMoR2rD5jHQP6GmXx8uSL/Ge6JWbd+A9LQGwlfaVEs7xL9k/EYrBsH6n
XLFvysR3IM9HebJifIzCNG2zGF8lM5JoXlv71kK9D8P037GrIlkaVd12YEDe
a6PIGqPJZvvERZThz+t8TApRNBmni/722LGNKklto2KeDqaKbmy3FVJR/yPP
sj3cb56h4ls/Iee5KT4caPbVCokTKyYEJPwBFev2iqW9ZDg9sJEC5hGqlqZP
UszHpFm1wiFTR2VAe+gUdsGwSwigsfLKIa9d7clLyizERwd5TVhuaSaSHSHM
UMLkk0QVzKPyLH+rwg/6LCmCVEGq1lZunzE3i1umUQ9AxgSG/NBOxv9cQvjH
yRYCrElLCrYUwG4TP1aSW7sDP15lqQr02FRACCRkw8OnS3OjoX+9g7Dqi1ZI
wsehgw0uu1qUh7Bg+WnDVBFYaCA+T3ZJ/X9phUFZnMvCw61CVNEWvPv5Zme5
iSUSsZKE1q8fFDjb+fTMiAsOIq9pe4o5T1C+wcL1716PleyU5ZJpeT7tKkFC
mGIoO7kLPf8wv1z3J9Pr+HDZWrqw/3g8hBLMySyKGK8iWewN9LBL5xMNDMLQ
ZA/xgg5hkhwKFFYk8REHpPAG9yTCDw/UJ+ihATzWxh4jYCVX2YKyyxPy2y7V
eDvO0ZUwu4HDSQ8HHv+DqZK3195ax2G7rQoXsUepg9e1E46KMWdV/XeLf7rm
DDb9Hxdaq5nMN1tSDlzgw0KMk0OGSTbF3Gak3gWrT1e4trSHNgiesrAO/7WX
5E9aELQ8SE0D1p/zWKohGXxK0lgoC16Zt6tR5sKfyE/jnNzCdLMF4mfdufTs
rp8tv4XYmEEa8DdcYr5C3CmzbzcYVAJYbcBdMD4CGCapzqArz85Km9w31wu7
vK1WWVuCVVq82EMdg5VE9u3n7wg9L0Q692vXNaNQIJGAyapszb33wnGTX0/G
BciH+HwDoK/Q1pLd4NoEVXSmZUXjO18++chHw5ex0wnoIh7Uq5m52CwpvduD
pc+nig9DjnqkXGkbS4wTBOmo4pY7f7Z+HJvsruBcJ2ERPES37Lnv2bcQHP7r
xUMvtwgOkdCwsq+IbifSA06f3r+VQ3jQfCXt6SzIfoPdxfw4ObT/oS2lfuKh
y5MX+q3iFQaoAN4SHOsDtIyum7Ge7Bp7gZvbQlIZGZhgca/xqspTv3fayirQ
dZxQnbqzRNHXqjcNK4kFJuLDdkijkIcnam5xEVHWMZoPDQVZPuGSHr8ObvyW
8yJC/bQyc+ji0hGWlUQUWbQZhAnascTyOGEjdzjqnl0lDo5bVuPr89zRun3D
BMroShggA0ln5hhhx+g9ubSLEDFY9uQlFzXrO+5c1UqsFsDf+ZT9yI8ngc3K
kHNnDRVQPiU7HiBbf3bJWxGxU5/KwbL9/Rd5wUXK3KPlY02plbEgmpdCCILP
lLLiQBv+gjVpGGhsvQy8/FnRsgQ6yaBkbvJHNDlizy+ReJkTZzlUhvSrhjCJ
5J8cB7fDYTn6piHe4IKLKnBlHDjxhw1otIFgj6IwQVEquQKhqOkniaUc1+0F
Gm9aO/G0pRc58wH7SR+ww6PslduEh5Nzdk8XGMjdyLe413iPwFCAp/aoIqz4
N2z1DThsJM7hyHi6A0vJkPMKnuHqlSMO7EXlTFFj49wwHSZN6P56O73wh80m
hq8xY99WdonyzUYsUBmIVAGXbJsW31V7yrEDrwhc5ByetfzfiRLuRtmhRoH0
1/KIVVLQx9f/bgszYWNjyL+nrNxrP14SSocNqc0mcIuaoRrU2aFWEhWcGExF
zFpH7joDgBmYD2EUzUmxQhZ+gQu2htcj47Rq8lo3SAnyAaSfJFv5/O1AQW0h
NBugY+8XIwdMpuUV7t6Bhp6TtibAitbDVkUfJsMaIf+o+ksiKiym1Q6XOMVZ
0rgHwSB9QgIBjZr9Jqu7hyrdIMKpjby3P2mXQMUvStcAvRnvRrqRdhn5qMJ3
4wtLe6NzcN1prXnOWlIqgHAsG6APpep8wGP+S3lCko9TXTLGuLZ2ZvOy9vNe
9iwgn/gvPqHId3YEsZsIvks+h9OpcsBYleI5tzNjwxV6Wihxf3owKBvVWrZY
A+eAkVBPnjgOUBR99yC5g7tPuazEGsHjRfnckgb3MwAu1uJwNYKnTW2gIR7x
ke8twzZ2+XrTBnik7pfMUfs0XypCiYmssLy1SMUGrR//jSy7yA0trajCD8eh
2HGP9aXYTuIuF33bNnkE4KyYRha/MkPtepuj9o4jxVV6NDcWvgSNBXTfZ3xh
D2MNltDtDaxeUV/i+j34YVfwqW/MQpIZthm7V7+eQ7EhdCpqIl8HN7sRU0ne
8zJ0sFd6qUGxUl6OGyBU9hWJ/Yn0DQxwITBWUcQbRYu+Qwi/kdcwrcRO4piD
XG7/bxbgUZ/mtASn8iwjIKwSUkaHDFTfyeqNOJmh0m+tuTr2zNG5gn2baWU2
hYxMog7hXsk2Ya/9MJDjA9XOmdvcPOXb5q/aSy9fSD7jUFoTzvx+lJNh3r/H
IQsZ799a46u759UX9N29fy2uHoAqxSJBM6ZPBefyks8KYstKpJz9MEmrf6RC
JSTDWmHyACBGt3OJwon1icagxD7PH4q+751lREHvhm3xrYIbMIZdsmOeeujD
5RLO/i93M50vflW33iaI/1tIPQUY2uy038Ln3gQwol9+Lp/HtA2pacMSjJ3+
Yz/F1bsduUw42E6DkrCvVa65xoHjZ5EhBGOerwH+Mwz3hKhUsaD75QtYCQtn
z48oWN5mt5mmT2VIVTrrlxljVxqIdaI2O1j/XZCTLGBuDhhWh9dQYd55gx24
hqKe1AVzo8jlcgETI0/bh/YFKz7vcFmhhI1H3qsK/pO9xlpiF+E9TzhJi1TN
ffEqLf2c6UH4C3+7hnZKWsb92xNG5MOVzKR3sdrnGzg1vbaKF1oIBaVkGnBT
wPbd/FgpNw4mOUCSGF9sWsHtZy7e/hyWl5bSSirdC+1qjr+qcnY7VeNbbzY7
S7ePrsllIWMVpzTGFdcZHs4Jtb7+7hiQ9hvqljz+18HVXgTTpX8ZfOwEso/4
Og2b8npETmVi79GJto9sE0H4NO3MXeIw40VG9kzUQqHEj8i2Gq5L+zddrO3l
mlch9hY0Yy4aPvkwdByCrXNcQtoDFrEGYHjONDF8WU2lXz2PKwQzFHZrOCX/
7ENzjGQBS8OALRmfnem/1YifJodtw97o7QaQKBGlocndqwx+IlMCmulB0YJ7
tOpHB8Ijhr/P3Oonwyqr5q8UZy0QXrZx51AxqMymze+Jwg936nN6HOBN61Z9
IP2uSu8T6g7FrVe7GGXGv92QGngtVSyzwqS63AaDGuCsR5xNxneACw23Nikj
wXAjW//dLKbJ+qJdjw8XbjJVrbBl4ApwRkwPOiSPKCY15hjJVhPIyOpFtnHs
ilJQvBCxpYj6RuhPxbC47zCkk6fwzBpEi1dIiGbODRTIsn1fztO52rVxVxhl
aSyK+y+8t+zKFKNsz5oAd8wZZpcbl34zMgsEwv0ZlHBvW+n/85vCArd57B5Y
zQMFZDzLJYitq54eoRh4biG7DmbaXHvDk1ZdNWpRg+ewvVqMoHbUHdMEBKs6
xv65ewmhDBWK7H7eax8rWzWpGJoufvy+gEuv4PWKLIj/p7G0UdTruYivJyww
l8qUk0nCX9igJW73vV1JoxfnLkEMrP/7uq/haeL8WR+ofpVhXopq7APY7Ffp
8uZDicg9Ti7LN3Oqapxa0UCczWw4gZLcw/na4lMPic4ADOMq+nCwI4Uru5st
zDjzifd927O8zO6aO2x/ei/sWdQEhOjuavp9C6UIJmNGpOSfECbjZJYzBCQZ
W2CJB1YIfQWIhdAp1nIGJCnYcWzC2uWeVY21vNJz9xFmPJPYv88SBVxvagI6
Cy9PQ1rgby3Hdtd6+tx9KC9tzagi7F7VuSAMbcA9Pj4aJWhBzHQ3boP3KsM4
ObNirmiDtNUnNxQdoItfC/Iuf9vZOtu8LxHiMetq04Cuu+8oVsSADkbRl43C
CjbHjo/+9SY9fDo3OV2GIdaa8G4lRX+WLObWkRyWPm38CJgKIfeyIMWKvscy
WalhZlTvrGRZyJq5NV5f6DRVz8OB0Esww7u8NOzTfjevspPR8wUzSjfIxinb
GCHOJ/jXoQ57AoPKkYC2KduQ4bf2lLSa6uwU6IAe3d0YnfzVivYu837stxjd
VKreGs+X4eveNwGxsnk66a0mYVR+8Ja1FBKtYFZ3EPRkcHx2lAofd2gHSseO
rHjXONONAJLX1ECWc0jnJTWqgoycJ5ZS71HHNDiz64N+k0pA4LOD/y2WUN7f
851daG4yM4nxsrC7y1o9YUqg8LtyK4zyBhhx8kPOjXJIYW3v1zjJvOO+BVkM
zMvXbH9hQ6MNEWK+Al3CkZyb//0NUA3PDqtkOkurflAu/YIYzL6FMaZTXelD
ykqXCLODRE8YOEJl+R5zAuyqG/2sjUDrvMUbQBz4MpnWyyeijNL2ZUvedqtN
cUFpIHwd+5tBknNsjR7LguDZucFCDpoOR9hmoHynJuHqcrEuviTbLbzvCTxu
IkniAhzmepGyCby1gpXzYUNqcZ4fFOiYAdb2k6PIfzyk0K4NNTypjeSjpd9j
Xek2nGxqjBqzGFU43g3LTE9aXjfYDv7Hblc4RjmGZPR9T8yns8bVhuMtBFrT
OupI+Zq52rLrphNPxdRPuoEbpPQ8hhycGZP4Nnuw026xBPxkxcF2Vd0RkEN4
G2YOcfi4R2/7e3B/9KxDq8t0I5Q4pik9KYGLIx8kKOdcMwtwXYyt7n+0weXP
VyqBnCrD2R/M1QWMbbGIEcr9Yu2RsG3C2F0eO48dEz5x0i8oVxZmeS3XEUj2
TXG6xu7oe+3vDL+QqLvBZtnrG2G+65PlxXMoWEyMt77cUfmcubC6B1qQY1PH
TI9kHjV3bYa1r+caj5FbLdCGOtJX4YUDUUTTo+Cekd66fPGqzw8qNxg09tRI
QvbOtBOmMt2RSs0idjlS1XWYJno3QU0Bxy7ckH14ch45d1OwVg8Qk37hXD4q
iIuY3UfvE53RXWYAbSN3mkmSZUBwBhd/oK+oR9EztnNljlHTj/pcxfXqztV/
TXD50YbUyj2PqWWuzcgjEP6wIdw4ywx8Bt77ScHTVoHta+OPJf7X1Er5SqwW
xjaW1jLFIzYe6MOUq+er4JN19fF0AUzbyzBUwc4ntSxoyT6HnPStSzgeAf0J
kN5DNsSpT1T+V+dMO7anN6u4nyusztvFavOqvGuVFroBFV8ec3KDh6QHdPWJ
qdEzUeoMjXBSAEtm9v7KL67CHosJZEOmR4qhfgXREV1JtQyYMdp2ChIgI9FT
GCLU9ZIE17fJWFqTQ2lnnGtJfRqFtMbvvFpLpMlnoM4TFKYMNohUPcJ3SO6x
8FdTG7MQylUmljM1jBHJEnSgo9APwNv6xxoMVEfvnqTiXHkmqrC7gUAkXUUW
IELQAzll0qU1h+TDdJKaSLJQjTtYTRkMnRlZdiAU5yePHzxcCO7mf8n9nwKC
6mOm32ozFCihrBVHYKx9w5AsW/FdnHqNawW4ZCAtEvWiqZjBWEndm2Yl8PH+
hXT3MbcA7gY7MxB2CXLPlIv/VZK4UeuW9p653ii/LQyj+qJ2z8sUZHU5K4J4
rQrKPeTgYFElM5dluiTXksXGIbsWzLWytMz5ApHgoJlL0qIKO8tnPjqmjj4E
HMK+Bcis3ruDH20veekN70yk4xKhssMghvNDIBL7/2RVnc/uZPmYikUvw8oR
rfibz47dPzj67W6Q7swEJpW1DfoCYUG79bUfYGNchzN7ai9w3uyS+0znEDEb
/hN+wsr3zx0o3ltOuI4RaHj+15PX2ruvli3yOyVb+wcdEXY6OUGdM89U2Acg
eRTI7f9COWmVWTpLzHAzfulhlFlWTy3d0F8iaNONfq7LUMHhQirM0Mimx6Pl
kPwjmiFTE0xWn4aNbLpMP/q66qUxbBTXTm/QTyhQ/0YKn3wy4l8ZsFQcEW1V
w5CEUQZAxf444i6GCjDx69LnF4fscfmHEBBLELlvvVRb8ppsoVTmhH+mg760
2RTXat0lgLfKODu5s+gpZJ2gPbGrQaxgaQ+BmMXEWB2qiuzslpTj3ZJnXlGM
7OurOhyYe3YQiJFVennp3BqvADsOfefaZ27BjEqvoBntk8aF3U1DL4Mo8ZEe
03s06qqt7KKqUcoOU+NJ/zLefrVnf3lhnSyE1rO1KTl1QwNKB+pBGHAo3bQx
HBWy+AY/d15SSs3ikzwyRA1Ez4woMjF5a8obyMg2MUJKT92cPPd2NpuP/SFe
oPK1rNErtSXFQmizAMRgazI6n8o8Zi/hL8KmfR7tF7gC+SR4P/MeV0FPdUFw
dHrj8gZDc1OvjWrzF7U0sF7q4lt9oIrm1NLAl2+0NHn8TLXODDiI5BSzqrmg
DVS4pid0GRn4HOTtj/pYLgDl4mEY/90fC2GuoXPYPNMBnj9+Sqn9WfBTj4ls
bYbxk4nzPOBIsNiKz3iNhxyJ7F2kaC1SBfAQ+XR8GwYgWe8YDlJGMW5Wmg5j
pUMPH2Ebbd33RqTUqDxtZqCe0tujfL4nuVT+5Zh2Xa77wmOj/0wL56wl4SLX
YYDo1Ktl5zflcc6BdmIm+ZNrv99p791+sM0db0kyrqZFFLOK4tbRo2TBM42I
aYvSNFZXvphmq5ayds48Mxry0YP8/0dp0faYr2BeLUI3mvFDtsAYS2qH6nku
bseZpSLnnwMoqG26ZiYFYiM3ehRYZp0yCotETbCXjElAu+3dCY7duqw9ziQZ
1MQTWrLB8wD/M9jEv28jPVPITD/ZlS2Ki8KklYCQUaBXvTJm8poaibaaEn4L
SbhfTv3fAHV3s0vK8+i2h9ItVvw5bH235WzzE2X3ceKtKv5XDjjC4Sm+AgN4
4jzlDLPc5nXDi2z1Nc55wsGVqL0K0d7clvTkow0lRQoqMS/LR6SasESBSrvu
44lOxFjn0iXRWjYLdQrL/NZ97P14eDkcqIRz4NDalAu1Sm+7pN1Qa9xidOxW
yeWiOSPhybQvkyRPENoKRueKaJUQ0yuOmXUwIU8ilYyB4fDy52v0zBEIRcK7
o7t/Lru0Aziujfwf7MHKNJiIVnY5qdnHWujnoerAkKY3Z4h3eAL1wT5QWKh4
Tq5rkpfwlKiOwZrmClw5zNPN8NYUPf/aFxCWTmg/Yttw7XupNwKrvc9jeexT
0razFLFfys+ua8zUCZuE3ojTptEqqh0oftucO+O0h1Mg7vXAVQGgKK9PzVtv
KCYCZMYE2RS1jZbgMUspG0ocxizrN/ArVUPPKEE+PCS7twJKhSJ2cWT8Gs+F
RDz+S4Pj9yGqq4wxavQH+H43rgPdWbTcHkwV7RQHk+sKXV333N0hCQpROxRT
42bQ2tLuTDSgxGnm1Zxnc7l0w0NQDfbRo7lrHxfq9obCNr7+qEPdSRZM0avw
GUeUMZBNvthfaZs2IDhJ3wNUBe2RyqVMqiQmrPGlmhX5TQxD30q60jp3qDx9
Ad3i+KZzZ2BWRgwvrZbkkr5hC0wVcA16V7OUKJhLo713WKinjPv9dTahThb+
3RwBhJBOsobaZEo3er6ycVsxv6RxZnNZp3T/XynIQ48AJl46kyGP9wq2sp/+
nZIfUWLi8j9fyQV8vLvmVJvbghR17d/8LyheC5xNnAFnr6hIRdRXSImOPA25
fBFMogeBI3glEAFZAGB4KPkxU5y2gb9D1+gAED7EjBDhHg0RG02hvLYmZn2X
3yMeCRpVWUL1HZ8L9YFSW6HSchrjr6NW4bd4K2zfumdwcVahVNJgIGaeZekq
ah7vaENTgVIkdnCfSdtSFeiwWeXF1SMEwoaKLA4EYbnKK9uWqDK78Z5agLS1
COzphXUKxF1SZH7Am7tGjuTBTBaDLBx8EXgYKo9NpVO8X6pUVsLjEagfncGP
onIPt4+fguOYXs8utPCVWh0qqQS9OSeqqpA8aRcYM9RL1xC6VHbqZBLni2KJ
fqyo1Lez+TZCAoJDCqT3WPVf6lSjLIss3bIWQMdUvCzjPELKq6+U40vpWF5R
/fBusMTKZ8Ijq0tQDfl+tE3hoVFQOSNLMcOsfpAQrj05ZpQZ/jzGoqTyg1yx
/Z6haynqCJUzNdOrfBHGwHvXBzMT5V+dy8kklxf5QVz6zh1d2VDV1mfZ+5Xz
vrsA5s+CuH6nlV91ZQNjXg/xL2TrKg3Ox5ZM+HNlyUr/ACZjfTnsf2qlqohz
MmZGtAH3gp2YVqcIexNprK3JeqPBLrqK4Kx72aTo8JmTrIgDlATl2H7K9Ycg
qgZgHUOPYaAzdvTLyqidPBUyS3op5MW3luiaMRkbe6ZqxXUQcTh2UInKByX2
NyIDRt1Qmik0KJtADb+L8jW1esAW7m1Y18ziOkiFEaRscEyF6sy80KgqDjAA
Ep6Zub2b4kD8zVdTuf/yUwJxTZzjOdvlXxtw5sze36G+vCmHWAt0Lc3Yt6ik
oagF1ILrum/S6xvuo14Xud00o/AtXMgTAOcrxzy062Bqb800sHTJHqFBfsUl
csKxTzb7PhglTW1ZtICKrdUcsVeRaI3BthNsIpm/b7zImaIKR75grwh8zxkp
Xwz6YV5NIUbcJnwKbMCmFZUs5FEnNywbbAIvoATZ41El/venPz1IURph1DIE
revNbh5/K2rAu5MKfEeAWaaDQezHJLlYA4CYx5/dVr+iDrTbhpGK/+uR00+W
iAGREHYPxplrsUt9+gGxMc/a+DMKuefc07ny/kKXk5SshgwE/+UpVpkcP1GK
GvJ8A7fuySN7NWN77rLsgmfX4T/1a3el6p8JZestrMlJ0qbockDfkVvCgpa+
nalihJrt56jn7XpYHD7cuIZFAji0bEIRkUWDVYwRzBuVeFAq0x48zd9eDJOC
o4ujTFt8WxKP5jQ9PzJi4EYe9P42b/D1NmP+cNBb8UDT3X5wt+y9YwJhGpWf
Z4vBQ77OtC+u7Tu/u0lw4hSrRHS+cSE8lkzFcSPxD2IcQrN6SLqy7IpJJB60
WP2+ezE93QACSYXvmjQX8YX2MtJqZIIBPsulioox7Gfh2pDoBbwzio0FSxj0
Vh9ZCY6d1NiUSts38yiZ+7gsESlZd5GHNxumTyL0fu+RlzqJD6tlZdGGrbIw
VdZhmX9fh7OZisOrdx4QlEgSCUAuk8DE0S9fXxpSpBPLqzo8UTHKXfvOtRoC
9bJ9s7RGJr51kE3JTNC8qCA5kDvMZsygHwpNqvqiek6TER2feXRfmIIxIopb
2O/8gCG279Zf1PeVSuiMhwK/H6/a0PBrY8paGSK3Jqs3Emj2/thHcTI3/YW9
TeW6CbQ2Hv9L7vlOA5qf7YHGHGrLLFVr9TXeA9a613froM3WYqIKmTZhhrNN
KO6cJ5HnL10BMcNeoeGMUTwoQYmkvr5eFPlqeCHNC+HXbaeOxfbyMB7PtYVl
6KTZpQ3ljSluMTxfcPtRR4TVQE2L3qdaTguRTEd8N2M7yNF6Ktb8LBMMq5gs
GBLYXAF14XjSMYpBlmmZFPilmSnIeZN/rC4scHdYxcHIS9JAeqkfVj4EWMB+
MUPUtkywD+QJQwL6ZysHKpvbA2IREGm+P2+0zSHmug34iQoYnmSY8gfOrd0L
FjUwATkUyUtbufe5PQSRz7tNHUbbgdDFZDAQsoh9RfRQe4e/ofBlgBxCueu7
TgApse6PbgDdtCprdjsXCKTfQ887zse2bTSoZIuT+VqDKEDQsnmJraANLNIG
/CZBY493GuhEbKelqhvhOfmsw9ULEgBSXT+3W9gZLRUxfpL+t8EHrUOw43eJ
dXfnqPg7aZFW7HORtgN3bXKr/Yxy59925iTSPxVz4Yv00S1VsKey+F7qjdhO
PK4vspgBBf3pFgi0BcclE2i51b4fDRCm9L3Rf6XiTZ9Ik2C3CVMfhcTjqvGG
AewU19B/ujg37U3XSP4kCiUoPWyeiP7SpTI6REi7awESJzsqV3RAHWTXhrwU
Rm6pNNuyuzYSGn5q2u6qHdWB81U/Fq8HzMAeewzqW508JeJRJP23nXBjd5Iz
Gj4porJXLzoCm7VgCvOntXL2LUPJTaGPaytM5y9Ehb+fTcX1V0NYBkIr9FF+
5NZaZjrH3ImJ2WhHhrO0QpjWH1a7eoDZWmsZoQLk6lSTC8dJ/9XJzz2jQEyq
5HIx8IUtaqGQU8hQkr7XS56c0VwWg+UX5oxA9Vi+/t2FjPK8ZOKDJ+6PV72v
DVnfwp5Wp4vbPqKL+sR/JoqP6DvUjK10FCHMsW4oh2Ox0hDXfg1RKlBquNSr
Rf0vordbZRyLhNXt7Z+MZXk2cJ0w7xWQPFzVvstreaRck3eslut4L9pGoLUu
gsyPNzeCaHuQwiX/s2TQgCJCUtz4PEZ2NqF6bqszsl9Ym2Sm41z5CEnxE6Yy
qhz50lGktevTv4I/ChlrEMHTPxKBDcb+79n2xrdCvK2wCJ7YQVnzYH55isOl
C0swmMwzPG3D/nInUsrFpmfYRd6dRD9LMJ7v3FoPdVWBib0psvFmad9reOCd
9jf9MMb04TImRJes0q1WbvmBardNQB6HGwcTrZk+aJPhpzL9zN20QxYAAgBu
vgE18Zx9dDcbB4VMO/s9wSU2zYPkez9a6O8GBbAbjQAkny1Bqpskdd4PWOyZ
wpWr8hby2PpQpx3sGfzFPJKGhfzIgcoXgXKMC4tHD9xNKZdEyxaFktQxC5wM
dPOExqFZHtFfZ5N8XLEWXeT7RpBhwiDpUtUWqEqppFJ99ZisLev5jZkeC4t0
w3ZPZWldGGkgRVfvlSPyht8Oa4nRoShK4gbyD4M13p7FFjjzFAYDZF+lgBl0
YeLuRbQa1XFFKoOQyXw/tXLXozE9Uy0Ildxvd11sKxsWEkWUKbX3TF6rXHO3
gPu4tiJBuktD/KBsvmF/eojADQfzj+DvLSO4NKI4WPG/5ln374bIcjE8GStU
s5KCg+68cXIfGUdBAc/a/jl8kLvQg9szI8YmOHQsrUS2aIb1/D+B0DGKZ2Rb
3CqIYbx7+KU0Sx9jF91ll4ZzQqz9+x4v+/Rs8chI8PcLf0j8vgRDxQjVS1E2
CsKoJPVsArDCodfpaFy7LpY1t9bsIQp5lzSV9hm0MLeri38RTdu/iYcV9JRk
ABnbAHKuiVLBy8OPLqomoDwusO8fOaQOLYOLXr50orY9py/PeIZQXpwtiQtk
iPj9p9QrNzlIibZH+tpazdovlnXQmkE7us/Aa5YdaEs9gjsdXIXnBQSdd8qQ
h/02Zvn0ldx8tY5i4EwYgy6PlUpgPyW9klgZOCfy8UqaCNH2If6JtjOgEaJ7
d73reAJlHxP+TwUySgFIaHDxjA0MQ//2NlkvlfxK3PwKqecQUfIiN3Fc/Sdd
fzPmlQcCwX/Ow/5O1KDqY4siHnoyP2ta6Ujh0vT+J7Uh0fMZfS9e0/wwC6sq
0R51zH4WLxc/0Ii8bsoqO+I514L9Q5jUreCl4U/KeFQSOfvRvkbhnjrYqqjs
6SZ9yOQn+Ff3K6Vrjfqu65tX3/88G3LUrScUIks7yFy7tdoVRUX8lELpRC3h
sybkdZ7x7OWpAmgkacmP3qkt1qi1evBigLluxPiKHyLCktj6wCSVxsVKOuBT
3NUKT4vbneyJL+osWE4ATkgW5LKxIygxGDGmKRNBy7Fejnc91/H4zM3jQCHE
Ve5HGhuasgmTgPDgDn0Nt18glIX463Sg8LkIgy57leBzpjPCpCPufVuvdglB
IahmAjUpjw3Vz9CF5b2wD5OH5MD7OHoGd+YhrxyC4YEF8SKrfH3nkg2NWC0T
o9LeGus7XlRGHjjCR4xmibNh6R9fwpW/rEyF2TH3P5vUc+cDiaabgLEs5QBn
WQ1vArQ3Wsnlmp/FyuLTvK65KM6V1I4KmeRK46x9cgJkBvegv1yE7jjozRUZ
lvVefOu6Mz0oNevKsrZwfYl1ki5L+mY55+Mba3Ag6VLOh6A5/vKFXAYO2llj
i522oRbUB/WfjbEfjoV/XwHXDH1KoXHdSZOvEfRMxyGEJbJ3F7K+Gndax8h1
xZADYuAqNf7bi3017GtzIR78T9ea38FRF+aV9ZpLCkpmupMBhl9nGNnoD32z
TYAl7/uf1WosC2EPUI6KL7no67HR8bY4rC2g/UYea6Dz7n5kwQTY6u9iNYyq
AfypTs4xmlsX244iIRmd+dCn+tIJcztmiqqNH7UiB/qzuO7ekHewDh0frv7p
IQtl7+nHEbG+pbnAqeD7IrAFBrxYUR4FaQgZjvXIeEL1+BCLWW4LjnYgFI6i
wlpDHbDJSHhc3E/vpgKc77rHY2hQ5QYFORAUAYVbBvps+eBry0/BbTjs/pup
PTEl/knOf6R5Vuwl7BFRl5EacsvHQumu/QsnFoaa8uw4nZgCbcBvsR4bpDr3
R260+YVsxbO689rpk7OMg8F6VwBZWUqJ+GBAJt1Ash2Hvj22HErrM7XKK4N8
9tmESDXgQrojiIfkD3HVBng2QbgTRzFdnxg6fk0u9tINFnq9v3kNW7MBPGu8
5je4IBawRP44Fgif8ftSgu1eVSB1s5P+b7q4sf44zECHtWSiZozY5Hizxp5/
+SA8wiEeXwObgmq9P9itHwoVW3/F9Z9lrNMfkRQDIW2qvWw8FJdskSMw20/2
FEWZ+MEPbfnokfvbZZCuHmR42cekYa3xQKpBW5L0CDHZHbnxDR9glLHGIuxT
9s1Nv64rE9mOR5q9TosIOF++D2kgNaCGuJPUvNIspUDftNyGr97ZXPTWZA/V
XDOpO2rL5v2vdofcy3kx2pFGguWsOcOazXa6plu3rG2dY+i7/4AOfhI+dRRK
Zw+2D6Emi9Z7l6l4UNaa7e9ETP+BH0ai6wKs6UfGZuUmZCBqvznEk+Acm6xN
pzQLF3EnkY3OKBnNqLT4iq/u9jaTYCCXY9viUoSt5kRj5RG0xWgo1tTWPW1W
WK4lGY3GL7HdmEYsPCQfsDNKl6GZukdhWAmjFA8Gy89VNmlsiNXBTbJzxgDK
AKapmqX0q2pwKDAwTH6BTd2NjETfL9j9k6nhYy32h+uRCNl/K5BZvTLEbvJy
9+m731nJdELzd9D6iz7TFsyENXr3iXcAUV1rc+yq6DZIE2VwbCmJPuGqt8SA
X4O48b2y45d/Hkr/HND9mfdSwG9hymf3mW6ua1sXzlk/EpMwWD3eRmkkshQp
raIPvjSEkD8m4oTDb7m7a2rdeengOF6qsw8JLcUvrTUFgMULlnEjBnPLohiZ
ohFctBsEo0Dmb1hA0m2gDLNpxSKMCPndG5ijP/9H9jbXU45XoBCtoMfbpyGe
InY1UGrcZRvR1BnJwf4OEvO0n1IbNR7Ex6so3Ct60E6e3ZqkuzvXcOIevmxq
400GSjALXCZdEKWqfAZBUzOvWro5tabil38vP+XN6R4asYIxhd5OqRAvj0if
Fzb1lr9eoI05QFAYD4uR92ybvXgn7WS7c3oY12Nu3zIxFAPU/In0f1NEDa0W
vqnaIMZq/j8xfkCF3rEfYO8276hW2Hg7a5GH0/OpUs6whmk4S8N+jMsxt64h
ivdtYdd7F8RkddKDnn1ZozVfqNlNw4C6vOrfDzXO9IJcNozkysHgKqR1JfKu
AOe3alNnsplQ20LdHBN/RIUHIDcJqvATV+ot+H3Nk/wBFVoKrPNA6Lh54jIC
xwiOyiwhLIkkhkzl7XXh0bm2zqrtX4Lchw2ohXT/DCqpUk8qcUJySlTw35Ze
PvgvqCYByfcwaHRKx1eeP4ufDatYY7cOyyLtnqIGys+Qj4mEhWVhSd2Ln09x
ZtCF3hTnwpmdjqrxiuEC54gL6sQkMK1qWoXR9fb3y7PAlFQ0AssCxUvQ+2f+
DWa+nFZO4qkiA/8bJU1rwxn1gXRBLRTFFwBAhnSJrYV7P2poT0Vcp5jsIpj6
9b567tAL2Ajv86HpwXM3+6n/7O6iHL5LfpTpFv/s9bREXYsIFBwIR2XMpPpv
c2vC69TnzCDc6YOVH0MLP8CES4gdYm7RhqwMWSzrsMv/xWvW0+WcxKHLB1nY
Ot+w3RxIbc/JixLnrHBZIQ9XL8MH3oz5LRcCQmQOeZPcjylBciwq7QW6HLhn
xE1fcy1Mhyo4GRS/hoSeOB1Nf3Bx/m0IFOYHzTpTYNZRXq7LLfr6ivwVa9Rr
xiLnRPRmGj3YnaqFSDTdHKhdsWS6oe6ke8OkcZpfjXaRh7gXo+GT3kgh4GRG
BdWNJvrTJFKXi02jt7IVeRBjWaemb5HGorVZqx3IY1sgw+8yd4ow1cJDzYue
olFWEpGt5BpNYg+pcvlqhmioCffZPPvSHlfNfn8+aq0n4YVQiMSZXWfeH2Sk
PEo8MiEBCzj3Bukgmsad9+d+p2SZ6L+GVyFQU6USaoPlZiOOxitcoEM09B8D
uROIFSScrx4YhgjDKlomONJYUHUt1Z6kgD1zhdl/G5RSf8LF7KYngYlOwkr1
fSEE0yJTlkLU+ZqGFF91kHbWt5JE4h/W9SmG134ttkavvYM44HlJ8swgZi7R
guXF0aF2UTkjno7YeY806Qorc1Ininkpmg0wXeiH2kEwZb4hRW3uVODT0qIR
PWVYT4li9lsK0PXEVLCPiRgT1h4JNWT6NLiNZhIm1tor1grb6P4GDW0V83gW
QOkKCnsUMyuHrrsO2v64I5enEIb4O1nY+nemTo7TJslz6zNIEVn4YR2eWFBt
XO4rc5F2exwXH3U7jlrJaFPCpovYvacSCHKXHxtyyEipRL2IYCeB8qSABRCF
AfNGhKfJKtor3gZ/LY9t7NrCD2mmcioYrbr6UCk+ONmM6cBJcaBELBvycYAS
hMbu4CNrcMw0LW6uHpBnGvo6+5NzXWdYArrfimQ8xd5qVO8XM60rrEdlEM1K
0DFqutQDPiO31WQU55ADiO9A1lwIfL/+U9Cu7yn27UEhn6h0Q9VyhoJHt/a2
k3oUPxX3H1iZshapPej77mOzd4ub7137rjC2McxKfkMR55OkQwEfBSy+Kcw/
wz4DBRPQqBeclM5I/mlJXIRS/D6P9EozCq/Vb1IUfAROMMkNBPDpZDO7fLdG
bZ3fwynwtvxrdhLg33s5MSVr3Ue+0pbptbVRrtOedo8Y3N/DmoPqZSGKPySM
HjXX0Xyt0+FKIG/syK57uHq/decGnvS1AmFuhfQghBtxfwjWKutsvjESY65G
KoE4D/YcxgirUQdRh1wSH9HbSiAX+Kr/IeNsl7275gb8TsBTmdUmXYnfbALL
WZZRdJuIYWi1fmwpT6H9JY3xDbJSvjrUEEx/q6s+GbddXAZ686bgP5mTG+5/
TgKrvhMpUsaGcKIeB6KgBL30HebnIDYV9r5ClvdR980e3rpFWGTOxX9vOJW5
qPLX9XPnxQ2brS4l+gQfNmwgVwRCWHUomUhfo0WozneXyTYC8jaA1mJBdbaB
RGD2C2JoW+106KHdAkwjDIS4du8yYbCKJ/jviHQumhZ6G39ZSpLNxqiYR9b0
LuAa8c2NTzXMvKiTth2+FFxftmaWC6AOLU0Cm59QCi03bLaTYMRlXMhD9+S0
khgg+BTggtFa1E+NFkISaI1DiZ4IlD0E0nVvKqPD7d4bXxffpPYw1hm1aZh6
LyjUHJvlrMxrkAVJJ3sa4tWNA7WxSP9ggL65keJNXIPK2OGZqUVZKqfMipL1
7aBKpuroJg2ZOQboMt9MkPsq79tXpvHbbrUA5hwP8b+AOGCmZd3T4zt/M3UE
drGOht2CJ5NbZDQ/wAvvzmJfKCkzuiyAeeNmIfm+myfoGwg2Rmxk+nMHRUc9
SodC+l92Zq9Vx2Jbq/5aQnIQexVZgESHPupFEOo2hlthoBr3CLrhQ4B7EyLu
sDicCPb6IqyGK+Vm8s7fBdP6nb0TcfYXgYFhCOngTlnRH1gHodubvqrlOKI9
RuThSPx3ZHxwmUK0E7xOsMrruAP8Igzcu/GGpRnEpKoxHb+JP22SGaaYpknD
uic7LPVU+ApK0xG28rM9uA7HnZw2lG3zi0HWY73RCXOa8eS8cjzuX+F5SWar
VBJ3seV4ynPuT3JmG9nbsB4a4bODjCcElx+rmSDML8qCav0ATAC4gF5Xpbyv
/UfpGsCZuDa49BFDIYJuKCrs5Ik/TgzQFPVJpCIIBCiE+ZHjqzlsjNvK4eB6
KogcmcsE8MSfRC/CYUFG81La6Mry/SUoGrVQQb19DtTTfnuuZXRd6u6qzWjf
ne73EakX3GIlFjDdQJMIy3RSG+0FZnA1Kt2o9FzFExXcqg6i4pLCRHFw/PSR
9xcYtiF4/jRr+fzM/Mx8upEWT+5dUPRHATbqvjWcjHjT9mBDi2X9MhC31N4l
zFarw/ay1rOkBbEr8bgNYlut66mN6RIQeAAsbCfJtYyUTQz8Dry1k/33aGAf
Q7hh/kM4uVRZuDYjbJd+z50x18yyOHpfFYtoIwKNPJs3+tiKbaxe7gBcibkf
fE5ZzEtUe0Wedz2ZU88YpAmL4bafze9u67a0fFJvJcBwvhsB53bNmfMeb+ie
6dAGr+Ro9xgdNalXcGFGmh3raCzBKHZlELj4oad4QLoJ7rJWiWTD3uYQZsI/
pNskk3g9XVUpzHQPY2e/X5DfgqmuRks3dxPFT12TKiiFJwEDR/hFpSEZ008Z
8THeWqNQNTVrN31bZwAs47dcfMVT8X8X1ypJ8StCu3mA0KRzl2FnUCVI/A7M
TjR8/ZD5JzrsvQqDZnOPTlqVl5sOyCd4ABD+gxklFV13PPuyQ5I7Kd68uQ/6
kch7gzygrhCqNhCZrhHX7Cl/nNpEQlOumnGVvKpbnuj0as5heEBVQq2s+W+k
5GHqOqY/7DDRODlCI1d7lPh9xP1GCTVodJxD+MtlMT5s0mxRnCn7wwk4K60H
RhkHq9PO8Yz71g+7MEbcAPTGyheawVvSZ7Pr1CQ7sA3HYovCaqZuFX0KiiZ6
6h3FsWgBLgEj9Mm4PrYLbGKLzGJCLv/gJw10+NE1K5b3gSFaiqXWheUVlGkH
BYb+qHks9KTy3eaCjqJMwvVk6X83emzdvGk4ttmzcLFZqThokNU3lgtHe2BN
LjPZ5aPn4EID10v973JKW2qhHOffpydQPZouRXXxIxPlHujnXcFTk404Z3PD
+h8kr7/SgbjhS/qHweIyMInOEb6EhyyCeWRsjiskC19u6uWTmC4vsRi3LPRl
04bjVXfWIY/IZMY7rCiYmCCTpjy2495fkZ7im1Wj5/CZYpfjaUQmrrEs+WqV
f49Sy8LghPXmDRFKEnllN7IpzWuaSYaThJirLz+7xnX1ApicPqdiC+6OOlj5
8TxEPcSTQFkk8eDEl44yDHPMnwA36n/SbWMZQhAqaGPRPDzR0UDKjqUYAMJa
vtXn0nyFbGCOxCmheNjusre2huIy4Lb2H4qRFLYL7DLxIk85Bhzck0nnack4
Zc/rXVY+X1h6B5HDQG1OA0wcGQmAs8MXWTcE5AiFmSgGFJkoaKm0f41T8TNH
Qk68bOZoPdptSYJWVYFH0UaeY4fpxhPnyIfnXQ378NKVpzI2YH28T618vMa9
qQ+Ua3hGecn2M+ZSopCA3CFa7ZYaPTEMsSOUhZULcnd/RDuJ3GVEPFgSsJ5z
257DsSuYWMdvV2tGp/MM7bOYIMnRSX7s53uE1140wbkJLYTmJrf3xObFeDhd
df/Fa9zPASXWuG2O8YmobIvFhSI8TzUeM85AbmjQ9A5LwjHxjdrlVwTCjlfw
QoqRAcIp1DZMUX3Mfphtulw0KW2lkNZEOBjD9EM4pyABM0K49WxTDci0zTEz
cdoGlC0lENpT+pcfm8xP5SwrSIdvUA3XL5cnEC882Pi9CEaI/HdCioIoPm0k
G7PnyOzGTLGsum2ZnSvblxij7qpMYuek09W9+qbcm/GlW63Szq7Kc2DgUWQk
oqAFegLww9Jw9RXSXP58F27X+bvJr67uJdcUSeot/bAtdNi7gEpWC2LYQGJD
km5vi53mz28DC9QZ9HYuFnNBqDCOtAwEznN1TcsfKOQPdY0uN91P6Qnqahuk
rOuBVWTcnIbxZasjf21ny3mGG1sJ2p0qcuZbf7n0G2+Q40oxFGXCZQgqFVuI
rACKN+r+ssKXO4MkjYVl8GmrOizuVVSlHGVNup7tqldxFpPc30vr/ZJnmtdW
OaYw//hBD1jnqqgV0SodSm2UIFbg4eyiKnj0PRuZ6dIT/guzo/ClpYeHXAD3
aF+CpCZNI3E/tSOJ9eEOvyyt5b4PwyWSsSr8K9OXDMOj8RSH+BaMrWF8tUIh
6iCru54NGTF68ptWpy7rfmUH0Z/COpJsAOWhQjtrpvOuyRf6beDjVjgy6f6q
dr8kM3rr8aMM3CMagDh/0uwr6uR6y6o+isH+ag3Sa6UcSwXczxSY1ZwXCJa9
vD+egC7e+9lowNoM+2pb2UoNWFkU4iAvu9ArXAwGQFs/jS9PKB0caiQ8366g
qMV1ZuUEIp3tv1B5e9pJboTfRI/vHOlyCsAfduHuRjLDDiBmP2TLxDX7Y1oI
0RdYG8mMoML2gFCqtfeJV9s4hqmHA+oM+Gw1mRp1/CLSCTDB/51kXPrbMFwA
VgHvdWDqo9Q2GYcBgxQAu82bi8hdIRdPX0G3Rf9nBiJSAaVQJsXLEwN6ZFyy
l8ZVtXkl7dv9pcuiB1Z6kR7ye7SMNwShKG9VLNvBtJFRsQxqBUTvzMvJGcPt
DkSV8+NQb+Z9aRh/eSxcojly9xG3yCyGV5GLQs2943cBUKBxO+2MRbDvolIk
mXWkm++pBm+f25yjwi2UjbWu9Xf1uij6lIaRiAQcm41g5BUE9ncGhNNaJi93
e0/DOUrfrHCzqqvLv/ebBV+f9Fi+w9B1waV8Wbu9x9xnnx0CR2iOBT3eXN8X
OVvQLYNstFmUQ3apM7V3Xuizu5wZE5xGOyNoOanLxiKhFnP8abYGCNrTRKqO
m4YsGCErIsNKQeMbX9nbmMIrSvMy0hcx4v0r0KpHs4GGjM2NrOQ8S0xLQ04x
8ttGr+rR/J2o4+t9FKprraxzgrl02ofbkIP/NjdyLgG00P7SVEkhgLe5LdiW
6sh6Y73kZkREhLwUskyzU7ok13DPVvcHaKey16uJcx671y0dv1ITFgYcad47
vs7u1C3szfN4XKvC4agLu/KeKI9kujK33HGKfmuDG9ks5uRAvulcUu0Y+nhZ
TRbmm7NmLnY9LRgTuJvvADB5vawmWT6mLZAk6h3KORvF31GxqEqfOQmKd6eR
syoKxm3BaveGYkUXlsQFmKif4coL35pS9d/OwBTpePUWk9fgH1WuKbpfYHZc
ZJvqEaV7WZxIWCJYD+uGmiac4FaEWpY8+jdoQZG/3VRZx2nO5weYh2yJessp
OAJk1l+lN6dqP7sQ0QmCLnqEDQHM2/TO3/I+Cv1i8lef9hkShhC23kV1/R7z
M/S5g+fnoBiSz+D0b4BLJ+SWcvVA+8kbSXiYBpQhSMAJT5OidM2cbHjL1+pM
fcZwWoAJfxF+0jVteQBtLOPVureJNmL0snIAFQPRFkeCBwrgK/wp6e8HhWiR
GUL0BR82kY8RFHu6z6dXP/D+NPmurEYn4Gzfsj1FC8+5843tLpgXhKQyIsOd
2rYlvUM5zw3HwXXmsQhwvv3VHnBzlXIBxJh6Qla1idjtFbD6Naf3BrgmfrEG
DgOVienvsSmhKScwXgoTxV304ZmwJCoF1EmidrqVIoAIyen9EJw6Vc1b+qkA
bzTJMt5UEgPPJOM4ynpwQI5p5B2lhTJbfzxATs6F0aIiOiBlosAJttFb4KC+
XyqHp2LZGc1wP/OuxKH6tg0XMetzbYEvTfrpcaY4Ew74Xvban4K9mlEWjqr8
oqHnzVpx5JQ+Z5cGgZ0ui+D/Jtq720pSlOuYYNJ8UoeWo8Z1iJC6U7w3xbwg
8b3jxtQHZuv9Wm/xd1G2esAerN1Gyrx9aMZRnM8nO9xgSkQCt/R+vrOGRlDW
JrV7OMAu+oTfJT79y5ALqv+FFblFCmAySqDmuOtOg2BHCUTdL4oOBkdYyFSl
85S5olChndvMM1FhrwcV7cvy29jvDWrTBbEvghK6P+DFt7YI/DKkgIqkRLun
ORGEJnNHfHAo8pFNGnFyYa7z+RJ0EiyK1lPz5E4w9gybjDi5k1hbojuyNEuJ
1Zc0Jpa1h8qStTPjcnslkMCEKvapDZwxkjmsa5bQy3uceq70hlbyIgNzCP6X
SEe82tNdMNNgBHjSGYRJEX5UsrV79AjBY+44/PlFz+/rkbpzhpZybDDikzKT
8IE+3YQXBWbVthv29ImfqZ4lbfixrDuEyL37U9H8XbIqz/TirshrgXjUVkhK
JFdvb/V7RdTyVkhFAzGA80bOmtYDLmuysgNh+UMH4TKJqTQKf7Y0YDKrwru7
BdQ4Nt6cJf+Lcxoz3BxFPfiZ39OsdlyA0YXqMM36I4RASptccgpWqf6YSB4h
aGf2Fq83jmRwMUcCKOJ1sA0uqhNiyDSULiluQxz/ZNd9++M4WDDhKl/1Rlx4
d57v1/yzYhRg5mpNSBEE8QSixeXBHFeNYvqu7EQTTFv+Bsb9Wl3hU/aW+GSL
lhiuxn5q6EzaJmyBiCyNxYpu6hpue2ZsXKVFqz48q3D7J8DY66rKQmSHmSju
KeKejULWRSCmIyv2a9abPKU5s0mpKvxBvGNmJesnml+pNpTEWEPyaKo3YinB
7lcB/DbvQxZdahEmuJUuDvm1vob6iZcbfl6SxSU2vxaMCrEkgLUXlUQe1/36
l4iDppfY0T4Ia3QNlRXJAczVgpRufzz7Nut0j9mJxoZtuyazwRyfddjpVx20
yWYvW5VYd2qCSv9SiQcejz7uQbhFvdkdg22ha76Yy1hiv4xvfL8EpDTgGZpo
7Gk/sQQyuBdoqbq74BbW5bympkTZF6vhJj97b+6dD1P+Qc2pycR9dM+PI01O
BEtIjvqc/Q7bGQ4O1tZ4YmYHoSuDO7O0zmIEZoOxF4cu3kHFKa1JjzQm0gbo
fEegPM7CzRw0mRBih302G8bwXsME2g+eZjCQhvT27VV8CWXEFHbuUHuTXOQY
uOpmZHzeZZgfdmMCPrtbtpY1+Ncx0UEADDY2+vsrmMQMWImBQ77wBQYva22x
YvR1t56YnVUA46vfN61SZqKRk4t9npnggx/ovNOdsFR+IjjfNNZnFrQn8xxv
+61+UDWR1lW9JWwYeRkl24/JfKEdCM+V1WvfRGziYh/d/ozopBpOET3CnSjy
pvL5XWfDpNI13Azc8hZqES2zWYA0HiTTCmueQAGQlCM1akFGq+K/6110O4XY
h8Zf3Vb4HnHiF5xWqxn1xqRcFfb89p63hD2HD+/gklK1VPDN8HatjxPAUFHJ
2Gmyx80RNcLNi8N2sCmPiVq8aRnYgqDQ2umyegOcAq9ZONsCgxFMpoleVhSF
z/lNfMczN4Z3wvfjruKes1nsOZTe9zy/cDdZXofmI0m2zovpyN9xmLU0TJYT
bevAC+Mo4q7iC52tcFlTKmtZM3PtEIZd82/3I84c8t+N+1DuNfSXmJ7OD3Gv
Psud8q9lH1IGrhIspuuHNQex+57L9O8casGP5Q4BKlkTo/9x9xsSzY4oodRm
/1pVCXQ+g1i2f0TT5heZbCE5tSvPle8TE9L4UlJuGqLZgAiaJa6RrixPovZR
sgThTwTmEGTtfkGhAhdYXZe8vQPIzbmjm2R1bFTzAEMwIaX/vMsCycJmpTIG
Ft4eV1X1W8pTsN2elYtBCDF+2mgbjQWYOdlI7fhCcuSuk5w7kDSTj6vGYYKr
QDJl//LhB4mSZutJmS0Ted9Vl5GFlnyAwSF6Qy+dhySV+goR8cM1OzBELpm8
9vGdMnC6lQRg4tL+ld9r5HAbB9AbouIzfojj2E+cefu/LxljfrvDVlioWaaI
hsa2e4iWg2KlrQCK6ZNoQcwpEfaYf1XappQgrTNqi1+QuFYaiizTqtUTeBI4
j356codp1WT4kPqo5QAFT5wOmAF6sgpLz0l5QS0lS90YcIxhBC+0qf3wnl4Q
/t4mwAn4Jyqu1/TThMuFkYww+wE7Loj8k2Qut8KvbPGobGL9IT0vs2gZfjAp
z2UNVFxfc3BnlzPok3krtKwK9IIfIi2hO1dmwg7b4pmc8HP5NQmb77hC2hrD
UEq9EvONyP4YvyA7V0A9B8N+lnpG2EfsHa7Iui+TYDiUDcwzhggCf72WneSi
VPoahe+RebHU2PoKY3yc7k/gYTWMxNNq71WIqFGCn/3tkSjiKmlw7yKI2mlM
hPJH2K20YU+5bpcMaxcXPE+irVvYScfO89zvQQBkv4ooL24SEGIvtngquNLD
6K7D7HzS69jDdNhf7cgBYUvCB+88F4i89YqwCnG1JQVi8YK5hwwS+DKUAdfU
gz9jKKZrAmTx4pzFYw29nqRAazae+V9/3Wv5jnH6bJYfC9f/q0UA5lbS66i6
MAUh4U4iil//2sOvnzJm0aUL5vHLAy/msyqXbkd1Xf4lZwu2d+5gIYhDmFPu
YPILi6DzU69uGYd6evg+5QmmjjtxTve9GBlw1Y4Mklk9tTfG4rBU8QCIzmiX
HRdupKiv2R9Ma+eLmZMN6nSoJa3lXoZPkjqkPpkhpJCg5F/LbGwDBVbuNxsf
p7vCx+gvxh7LWz3Jhp1TsPoEXiGVM/DWEhi2nMJWOEi8F64uIOPW1T6zQlFy
3nyfPXPsscopYF2C476h4iXj4vsrcCfnuM/H6NlkgE/c8dXb6euA+RroCc7u
U86yV6bN/3e7HUqio3o3okUYnkYG06E5+jptOXvGgjlkpB+PpOysFoaUnhom
jbYuNWYp8kBgCkVjU6fIc5zDof7O5/o3y31i6DULVQ2PAsjS7qhE+FsmO61Y
u5IQi42YYPgAlsOlDTFPnV8JK2V7I2EcauIGOqmVA9idxB1uED40AhWOlskC
WF7tPOW8HJWY6ItA/ZGKKg0E4YS/zHGCGLpOUeX6yRJpkvtNHyqFoMHysoAo
tXVSCiuDYN+DncAYCAoq3heae2O6wOhiK6cJng8chSaFt695/IO9uqXdnBIW
MA80Jq3+zBfCM0Cy9XUF7+VFKMRoFOYp/45Sv9O3M0qMcCAdSP1NdfAyptXt
Mjmw5Pr2TpWVruFHQI1Jd5Be4ZsV7d5T0S+fGzAQlZ7P0gltenSnZomlJEsC
Kna67B7ljeykCDShBHukizz5RlrybBYGDoihw48oNgeMqN48jwsbmt/nSAlY
bf0rrR6NJhWs0F3XRVPXmOfZiA54ONUxK0JQV6eX3p4n+Oi6Tn4ksiRxYdVX
/PQd2MrObkjvLXVKpnzWIXKyLQjWeYVuo3LXQMqRE/GTTZtnOaE/qBB/Pci5
E8Va9Uv+L+CduO11rmHS0alNPliJXkYionFeFvbV4LjtmMArbupxa1ZgPw0I
KgLqe0Buont/3WlhXzo60W8XoDYwHC7H6H8m67vS+QvX3yiwcbeQbz/yvygW
O2und8kgYnBguk2erTW3jQp46N0phaYiJ5cR31OECxyApb0DZiv0oiDegTKj
GVZf2mh97Quj7Wc/abHnJacwYH3fA5i3abnTOTr2xG7Yw5G8phLc2OvL6lSb
Dgrj1I4b7zhybkDpv8thI2ZdyhYWL4qdCXiuB6Yo6x3eIQzt2dADibDbZQSv
D9roZOR7lRX18n1ErIiMLppCVm76KFe3/ZtnUhgqOQIyCb4em9Nx1Z5W+VL9
Fih/5chQo2MUiXe1LQV72YDAoS1yCwl+mkl70f4btZqpoHzj1IDA3+j7HmPa
im9HQ6UnSrZCF7ix4OblgFROUngtj0spoqzNkiZhia0/zU3jjnrl5/Qre3Wn
6yS/V+FbfLgERhlJBRU1BMYaOuYyjfl3gSdlepqNglg2WAO+FfgESCGnhVim
a5ueO6Ph1xsaz/RWn7XfbZJGMKsZUlufsjkulcOPYK5MSvxLlnxA90mxz+Og
HHyd7WknFCSQxm21iCgiE+PO0cu0dyuyPfcemCdKsnOzFoD9OLLSjHRZnUBN
dy64CPtU6Xy5BmA+p7mRy1uL7I40WVvdHxYdK6zOY8ug4bWZfeeY8/AnxBAP
I70JW9WnvnCkfeXmCm2MgI4C8OErO3dOFVcc0WkHQBrw1NCAcT6dTXe5cLE8
h2gal/65c/G4V4Hw4s9rstbfBAM3PpAB0gqzQ3NSWT1TR21t/fbpCfcN5Bx9
1QrDCGif3FMI0/MolUgBS5jhTTXyWRyge63BYwyxusFq7+m51dWlp1xyjKrf
MNHBnPGAX7vA80Rr++2QOmsYlKtTnQbGaCbCTmZrcrJJtz1cjaINB4bUfceU
22Rr0yp+0FNEm/H1/EVJ4fGLARqPHK4uGnULwbbMFSmG31xOZipyUiFZYom7
u5sZ+iI8AGNp2QBrvCCUxFoeGMjKFRZcGR2jdek7afXLvMFOMN+FcTJdkYEu
xijFMIzAHDoScggWM0y6+agC1/HXXUv6qNC3mF2yWQ948GAgtLDfq3xjrdkc
82BNyXfsdw6a9nBrWNdSLtlHEZUT8rekpI33x+7yJbQzg8qB+dSmwOTvZD8y
YYxCcO38oLqu1kciZoAh1LJW2VAGEGEcUKa6sSYFY1aS1rwlioTzBqu+IfK5
pWsLN9/aT3QGJdX33mbnFpvCzxTKBGYVyXOBDizm2HmLQw10ooPFqSp5R4oZ
faR/2AbSwzKkVe1nC+MRKGyhSdhzDmEMegEj8zWFaIijUJMrXdkytYjnUn4E
aEIAzBWlnQPuK2C4/aP3QynUwz+96e6lHTb8jYbJPLSk5ZlAs7SeoF+Gmwpy
krohcA337o2axKbTAsiVswhvIq86M+KzZSEerMlohhOisoz2Q9KFivnihzaP
kf3Rn/pFAuLcxNlDQ75sX9YPG/t9Y1jsNUNWk7HVg55hu1i2GDjNvlQu4FXv
N7HBcYDiWTPi8HhfpNnyUsMbQV3ND1ruscmRSj9Qvctz9nrljvRGFEnq02QJ
hmF0NFCv8J8Iv7nkrb6UEBuKxYW9/dVRd1FlvpPexKuiHuUoyjsGfz3xu2oL
r3+0Hu5aydFgY/UQqWfsKQ8hHl+ZlqBcHak7Y2sbpIKRvChXKoGuDi8Tmu9D
Cej2oCQf7sSQseVKhmSO8TEJVZgrxtzOMk/o4LTD3tbpPYl/PLuwyBDL+WO6
SDOORZzd91rkaAGm8hRSu1s2z65Cke2D5yF3g8s0DjkkVtFvu51f9exLX59p
JqYYUPWvxBPq4D2ZUvdJf6Wpei+yDoB9ZMr4r/Q2mpEpxbjW0klR3wpagS6F
OMxWUu4S4sj2QEWJdYYCGMfYlIg83UVfgKF8H+NuEPb3axOvMKD08YHUN1gj
49yl3Mh91i2Fr65QWeP5W1SPut0ThwgCw2dK5zTAOQTUU6hHHaXVo/gNcrEK
BN6GdPyIAwSFIF19F+MKXJ3W3myrEAw13d7kY+ORGBOxQz+SA7WTuKe6wUWr
KHqpNYhmRUh60uoIv6wGmQv9zS2zk8FoaFnPtn9+Z3SQg2B8XDjJzwAL7fYm
WVfLk8f5X/DIaGqlOQKAaKEfb4n39CVwqyI+E5j+NtG2+iiJF+Gb7bj+Zeiz
enZyre1N+o2C1d65Gjwbj3XYE80HyjL6mnxuHDTM8h0aLR9WB7HkEY3zMY5f
6axXg8nUdsjHMmmJUt3EoTID3D6JB27pelQi56k8lXFQx5XoEMW8VOeevuCY
6PtV0FxzeguiiEEe/G0ecSPt1yfo3wKGmoNmQZuJnVyenX/VktDUymG2ongt
TylCJCe54iJWS5kXbcBn1YiY4uenGN4yuGAnG+zPHJ7rShj+jVGOibl/LGM8
L6Z2EZwIiu5ayaQ7f0pgdI0UEzd9/af+6jW3+d+g9Hfbsrtd5WsIoUHDneSy
vJY9qtIEwndTa7tXv4cCfVfWhtarCXNeJVqs5DO7kiDaTPe72mtDyZEtj7YZ
UqZps+4xt3FsHNicVhEaJxnN+97Hh6uGHGvhpvKaCAsxRVimFO33mK2WCsWi
SjjqSMCEu1Y3rsOEwpyryIBeB5Nd+0oyb9/2GKdEbbOd3sUpHVAN5b5QM6YG
uEdNyavf0OWulxfdG8vm4ZxVw37afD+6TfRX4G8NlR7YVFZTOBrDbEHKFNyJ
P38VP+1LeVwk3QZHTtXJBQUqpY+8Fn9oZTE1JOmDMk9bn8vuKW4D0SRiL3hQ
6cKDz6iJCEFn+zkZ8iJ+VDKiO3wbQWahkkJDZuRrUDW/XBR2LfY/3oQ04iLC
zr3WtS5vg/M4xCMBOelIPTQw38vOGL3e/sM5BFhIsj01+QE8x3HseE57p8Ud
O+HhpcI42VJAjJ6lPfK7kUlvCo+vuN104Yuy3/S7h2Uw8735z0LmSeHh2SZ+
vQ1E5g7oeg2utcaP07MQjBPKapsYXyrkvQNcqFY8YCrccVtx+ecHYVzTdNw1
eEkEGpyjdaXDGzA+g4LAijFQEyAeX91INqaPDsWjOY/1OeNMddqTtykUmxK5
ieWSi4Cmsxe0jBEVikSqSBA7R9RVGhyW665NCB3E8hMkRwRV41A2rCWOwJz1
MCogzGPTDLSui2ZVRMuot1ftdHHcdcSO5n+gWrxPoO6HzePSvw7iH08FEmeZ
VzswPo0Jb/Xc612tqT7VcRhdQ8DZd0YC44wOpNKhnD1lZM72907O4RDCpCWB
ONCMT0awfxs2havc4Ug5l2drJKNev2J1/dxnK5B6dv+VufAWPG3zAD0NPiVz
WylOycqdOGmyVWY+huzpx2F18THZFAnhAnQlvEl8CKZJyAdeSJ1VUCBS7NRu
lp+Tt4I5U6KvHZtqTfwZPJYr7XRXT7rzA6HKfHeAI2DcIhOKDTaarpJpsMy2
n1jXz1SSX6GGhqlwOpGRHS7gvdfLOgRYqrUGF82JW+RtrSWsEMvIgiucFgjF
7Q7YeHzZWVqQ4qUWy5dQBqK3hUtpMmlGF5vIernxQw9lisGzz6nXBCpLkpQD
xoFGJ2YWxpadL4u3At/10aiBGQIvFrL5q8CdKV8FBWeLLEqFzVPyyfQKHwJU
1BgKCPFYKbnPOZEJJ7DD3OAiICk9e6/SdwkV2R7zdOom+5U6b/vqlQ4kbM31
+YsALu88DttlfIXGhxbeUqOyEvSE7CZp2VXXIfL/D0c3y1Y7yd6cSc+w4fFQ
PMrSVTkxMg1JLcXDUL1pw0clDAakhulVILzF1OtNTzAugWkiZxCX6A+b7uaq
fPPyW0hPCMRiuGRHI+NwsBrjBQIKcCeA6ReU5tMvhesFjOdHjrus5OLu4Ytm
WvPSX9hPGSvt7ARXKuiCuwl3Xe/z7tPZACyXYronr/xg86m5+/fplRlKwx1G
FtzkB33v2Q0+i1B1IL1QouRrb3NwlJGz8TcABoVtvEBU/9zDaU5RrjLvIt0H
+t5o1QoJSKP3IuZVKPg7go4aJlUd5kIVJm9UV7bpHHswBch+bTNiy9VI6x4b
SFiPbqndjIxgFijonuJ/dwxEkyIj7s2DX/slRRNktR1klybRNC4crqDtJYau
tlYIp0INMZZeKVWfkrZF6Z9HtH63sVRj/TfI9QmOJjfjK/0vd96Hu6/R8CZ7
du3ma8rMd+EoKhUpy7BvzaAALFkEVzLdFElGQM4THoZ/J6J1hEJ1a8B7WIaN
uP7VswU9uh1Wkxw5pamEbPv2miXMkMSzwhr71PYXUkW1t7hWuuDWESbfeEtT
R+XLyyMJ/W4LGXcJBkat+1Nr6gj7NuUuM7JH6Dnypd16ebVSSKdtZEk6NOqQ
gEYp6+lOtfznAzc9ak1JMymK2AvkaxWkLohA+1W7Afyyo7VUV4tFeE+4zLD7
V2jn5+0a6SFxgtWfisVn0epqyk46cOr+V5ctEsgutfM1tULAJsJEOpQZ5LOS
JOhLkqBWVCISMClxyACigGXwQDf3B5iNkTsLLPgGRVL9KgFGrH+hCdJ4Blcj
OnDK4aArnkWVcpaCg7pYuJvbeAEoQHLxRcJNM1p+oGEx9ncbA7fs9JgNi6/I
MwmQaoj0Y5tNfXJ7TwbclwfV0qhPB7FJ496wm4WTbBeyxSZ6Y3DszGAL905Z
KKZKKdhMYKLCL2CjsRf2zW0Bsxe8wiEY0PE17Y8yrfMrUQulkn7mFkFcbfox
xnw5ogmAJkG9BMvmUv2FCJ2s84UDCnhQvfth19U/ae4B1xhsIs7+Vgt9HQFf
uXqFFEN7IomzHOU+uspsNflZU22Y6Go120q53imeHDsFCrY4FFoGkK88HHXw
O8s6I/AEiEENlNpZMfYJmN2ZI4QO+QmiXsWSnxK9AYXzZmPyo8m7kW+aM3qH
/dGAqylX+/YsR6FOXsCYIips8KkAJwDvN4lc7bpuNewyPKnK1dbaMM2TREFQ
KArTAAeoSBdCKaAR1Jaes+1NLSg2NT0R1BSb+qQNnp4GIe9TRA6uvFGhbenT
2+9aG7WThSyQbgL9qRfIpv6bsPrYeH1BlKOg8h+fKTcm5w618FSFKEzzLdQo
9wZyLh1lq3yvhyr/R5egRjYdEPKnmt5Uiv//w4XkhDfIEGJE8f2y+oeikQHb
VlM/gMOzFeSonmBXwqK1Z0eT0HBnBVmwumPCfk0/S4bC8gT76o8SPNys6gPK
NwcYg+021WWNvrwhypF3ZQlGm6X1bhcLn1o65WQ/j8bmyYk7xOrgc1Z9A9ha
OcAt+uSQMgrNUXLSss/QSUVVkLFWQ4D8CNbT0xls006gYEkXzeymxIrR/+kT
c+Nk/L+7h6kMGvHhhNzmV3vm7L/UaUUa1A5YVyplGoG6ptuoOtEtqiIrCQ+Y
52/QwSFIb/RWLCABtt9Bohs0PlpTDMbJcGs/S4QizdsiQqvV1jc9Wa8ZjT6H
i4OXliW8MyIIBSxijQvF4J6s2l01ctfHhWZu9lDwDWJe2qTv5fk6T/eJo7t+
nQwM60ldEpHn+LIQh2bLUfWZAgpYeUXXXZUOY/nHnY33egBhoAwAJ1MenAJw
6rMP3NdHyad6WoRpPNPzBZ3UbXsWsGfSXzhs0+l0T7ttkPfay7JMkTsF26XW
u5EYBmTeKng73t0aAY7TjDK4REG+9Tv58Og2TkV1Vf66QHfYqDrOXIsFs/cc
7CjgM9L65NJLiXS6C5OAFudKhE326G2uOJBwbPQcaUyXfuVMBRv7UeDmpgAn
g7t2/ax9ormicctMJozgWsS005wpR+P68vOgpWq13aw6z+qEuRnhmTLdxaeF
O9RyZfSwpAMgG8Gz+h8tRAEBYPBJ1j1bCs9ATCBEwPgrmUat6zH/ciNEST9O
bM/uOrA9QImGWn0ep12AKS0dDQOywB5+iGGcpX15LWJBNtHmxuSYP377+x5j
lNU1AIf7ML/Yh2KPmeZtRDswjvcMaLvvnSA11Xi8mOY5fkcjGhapg1EPpUfv
hr+fYPLc3gDsiO/E7IO0mqO2zsNjcubotlA/BbPuGRidsKpuPA/K1UlKfQrB
lerjKNuMLJ18aUxb1aNadmRCVUacp6y5YqMvHe6SRLLWNWM6Q94R/mRSoSJy
YDO928m0hy0ePpkOox80xvv6tqCnvHqiQH2LpTwablO4hMiiItRHTuN5C0M5
i8/U13xV2f/jOmPcz8WOBo9SKlrO4OzLkFFE+iXhoteKPUG7ClZwSfBtwy7v
ymiirNTs8KSSb+k2zR/O1Gc6tDlQ7wXnO0VaxQ9eVgwOib7/UFtr2XgCtUP6
J98ra4P/SOcUjDcHSqIzGZXpMDLsfZ3TeplK+m2yAiwc1lQMiKjyIjmtBsg/
pzT/c7rTc1CREpdv+rdxZTrlSPc/Iq5SIYIApd1QI/kyCuritn6LaGUYV2Ax
L/jJq+umTZKgn3svH5OMRiChtGJJThAzPFFGZjBzSnoM4awcOAAffGehWbjP
3ogRHMBGQKQ4Ze3Hv94PLobaK/rjSFe82WMMYqkQaNboNcJ5pJFZo3KFxX1X
QdiFTEBlCxqcwUYN/lqgw36NjgWc7F/wSf0LpGJz0JYjLQRSqEmvnZvR2bq6
8AGwKTV+RN1FlNyhSnwofcYm7nP48iYwKeGk2y6rJwNtdkmlL3/hjUI3lQta
VL1dgxqdRfatrUmEPhdtoonMzrC3sdQSBtEN/M7mCrtAbV1yG/g3438Ugfq4
7naZpk/0+vnkTseCGBfOC1wl5q91MWVaUOVGSUL9wMrm3Y6q2F/lcrF5XUoO
yItrc61eu3+4FVwf3IQirJ2tYh61ybswu8DUzCepspKkrL20v4+qw7l+iDcK
gdhMPkCVxL5Oo9OmNDhFn1w2RLUkVvDxwNepI6ix8Z30JCStDQfgi1N1qsMt
dlODTi5X31ca23gQtyHB42hHScQvU+6p/L0tq+B+yjKsDzYaQ+cNnc8gOQLI
ZoVjwBg8RHzVQXCteVx6XWYsCXPaR7TnL/3z4Zq71S2s0dX6NHJNcR9Nu6a0
RoPp4aEjUIBlp1w5F3HvWXyvPov0N19AxVo6r8Sco9JV29obv50An9m/6+XU
B01M08Re7T765AZMsnAVqDq1YZvS3BV1GoAn6vElfWKD9TN/dWyPHVF1PMXm
HNMn0orGfuNqaxc5pgpmjw6u21pIodpJkHx/jnJXGIDYNQyQVrMqYf/RyjgY
rtxcWggg6jSW07RmMB0YqezqknOOQNP9HSfZaCRw6M3X3d6sMwycur5ywl7X
50OyY5GOYJgqGr+IZ/6qWzH3TXvnGEUIRixmrLyTtpKpfXsxro3mEQmPxBlg
WuGNjQF2JLy2T0x81i1HWzdm5TLG6FCtTyeLwdc6uC/Ps39b68rBPKieBVu2
zGmNYj2i74On5D27BzPYG8l6oMwRbsWdc+iPKnimfEiIKkvsMEO8hsNn5Nmy
SzLGIvUwt/fExUbn2kH8CLgs28sLh7bk/uQXsZ7K3ggluAP5q/RFxhG8d1jY
3Xpmijzjgs/Vrh2kEo0pgOW659IOZjVVrTnbiMwI13rZcZxbl9OhlZ5TIM60
TxBuOhEV0F2H0uKVN8BTkzs/+QHDt/6ekSkD+XLkGZprzJQAbfjkyjxK0uTr
FPRtceLL6K4E9MMbBYN7UHxTze9Y9I4xPZ1jslgKT2QMkuKjt3VkeVrjYS7m
Fp67fComPOgSjcn7WL3WNURQUlmlH3vfZ8+oE2Zw2CBLDW05DbSIXM/An9LJ
IDAkWVfLECa2/MQJAmB0axdY1jsk18KDsbtMACmOsg3/P8R08hi8hm3VBu7/
7Pl3ObbQ1YuypEN1m3Q7sh8GmoLBVSPH3G6hPYuxMTMsl8AWjsrmEt/EHvlJ
uc/Af7zWqf+zqVskpA3Yymrfz+dff0tNSzbJL2r7t/+YFXuhTgHpskEClmhm
ABbnT8dglIQGFt0Tl1ahZ1rxIF9aawQampoC8CFBRk8nAS/iNUSVSPdbzQ6L
yn9NKDTjQCkJ8BtHOpS9uYqLYj8YxW81g5R06tDYyJfJ9wrRl7T/Py/MIZEa
d+8dREOBIQKhzWcUV8PCG4Lko5T0Hi4srUNVsUkooZziVIzj6km63f8m7x2z
l2+jxb6nVqHcN/iaDfyQB+WKlCv0Cx5itxS+TEMdDKGB++iSZYs5/ywjoOVt
s8Yp5jw74SAlm+D5cgB5DKH5bkotoss/J23EyHvm+8Be3MmLhWYgtHvlVsKh
LAvrTst3rXM4cOmExqdSXyhCSLFjKLSyWuD9Hxoe6kNh+YX7pN69fiHa4eQF
Dg2yrqSvwLOZLyXYj5PhVipes5eVvpUNkeuCLGLcS+dnSLNyugJk4ft2VAia
0Qhqahq036qWX7V7PXcprFb8pMciMFBs88aukIiTdbRmdlGUEtth1VVOkCR4
Mpw6pOyNfn7T9lnHnRef4ecykO53e1zraF5+XtJYnsPlapZ4EQfQVHvDhEfM
fFpReE3Bg7KCMhueKAv08M1WOOolnIFp4qWxQz/o88LDhlIUlGSKLiPlQshq
j2bcLd9Goop+SehZB7b9P2jX1k1hKXXl++n0Hw+tCt+CrW52ijNxmCQj9Fk/
LXQYbvZNrSHZINjgMnph+sMDdkqMbwQHhncGQ7n2SdFTw8zpdHqrZAv1U2sV
aOr6vhvVrPVQ1jwOgmip+ypB435Aymrka1+4zAPdejdcmBDjB5tybd42uRf4
hcIF+Xze2UrYOSHJbZFANQVck+MiRITdYOV3Wrw4Zk0cZOT1SW1fWznRFstX
ys9PtGQZPT6Xiv8z97dzK8PUhkTwGQK1d7ZZbiAkJH4kBq/SFVM+X8tCRVAk
BDum+Y0MIEdsAKiWYs0ZAH+vcJsaV6Gumg+GY5o90H3TvYpuXE6zXr8FQ+1f
WgkbAz6pAZJURjwCADXtmSzng54cfxNLbXWS1zyZlkDd4kpeNYYkFKYfF7EW
YWBGeazK9qSqGG/HwlQQZYpIRILsVNVJndIPcuHF/pjNIq0OGZXcJ3/72ef2
0BhwXBH3mIgGz+5FJbMvtz/Shn0khUW+Xz0gZv37ciyUd4h8PtaPHnRwedXg
bzCO/XSnhupVlb8dJlV4Zfi7JoBQXpiingmr4MFadUp7KAVkLafiXSJEYGm8
Fgh+i/vTPJmf/eKrf3ArblD6zqCDE+bfqvhEgPW5M74mYdhH9EFRGp7Bpx/P
MlAbDj1OMIon2WDBZPZexlQSbL9KXTbHm2N8jNMF3ETGf/u6Wn7maFYVinzi
7E+jK2vy/Jt6vbkXF2IIKA861SVRsh6xA5FeWYTl2ClmZMhSnAXHmhg+IyTc
iuKjO33V4wEW60nRvkWfy8rsZ7b337sSYsVctAsywjqj2rogUV6z63W63+IO
+stV/z94aO2E7kCyDD0v6+pqd0WKEtlcXrFMfG/FzT/dheYuUdpYonlsl9qE
b+xFewb05FTU1TRuQlB9W/uMM4FB7SmTskiCxg3D/8FxOp1SVvf77brteh7o
Di6+fhA7hhttAih0HaRrlPdI5jlz0hHnUaoqNwT4Jquzm/+CVI2OmsC2GOXx
Na/CQz3sTHDJSXCMDXqGUlhYNuiTWGVAKnb36YPTH8Yz1Letv+u7FXB51P3K
Sz1Wm+Jhdd21KL3A24m2wH1v2dBGQIGIwL9iUFUtjxRAfXBQ2djFqpFIIlnj
Qq0v76p9x3YJ+V+Jfo1nR/5DMk+BfvhagE70vBjt+IT4Q/58SAaqI74qmrRp
okFIF+2ACZ7qUrfTdE1UY2bv+7BolgZNrmhcY3WDt4oLxCUgPFi90ouCKfWJ
L5zieo1s8zH373SxcQQnqL0GJS1OULH3MJklNrjaQ3LXJPZOhm1H9YsHYPPI
Sw9qy2OsETIno9QiYz+hwAVE6F7jmkI4S7BRLh/hvscNmRso8dy9Kq3sRQfo
X5HZqY1fiJRcIdBUxAJriXDC/kYb5w091sH66V5AHo4oX5XuX5m3S8uEoBJ1
RfljI9T8rDP+LndVH7saoN37nd0rGaIPa9z0ignErHAT/liwUQydZvNC+v4Z
XIPwro/WjirLJSmNvmDIN1boe/xLh32YqnV8RdsAA4QCoV2HfSRskwODcOMk
bPBtDABG2i1kRR02sGSvRi05tf8lrRIFuX1K8SN0LYEWWBG6/gJN4lsFB8BK
Lts82Lc8GjAhn966ulVB4TdPsPFQKpmq/MlrFpmq1sj33Bp0hC6SWi/4HNY1
uasN6hzJLHAMogqB+j6aT05SRb5lUZYnkMvWsC1hrPSn1h4cE8h1cvAxXl3B
3fWeB4w5gcBopSgibizb950VEfVnwvZjHPthNO8Nh/k6FwKwSMZrWDVlbron
alKnBc4CV/zDvqCPHtixNBmUDnLNH4EFpl1FYcGIrT7T6SQu7XeYNkr/8SDk
4OUs5UskGS3B6u+wT+aGwhSwLOJ/0unn8O/vSyfoQ6w71eQKMuoKBmaOTVpQ
FZ+jErcgsg9NjDLsg31v1FYTg1icKRD+JIdYzxbz807wmtzD0Id1YY1cBERH
jtIWhO0UDoR3F9O8SbmSF09njSQsMmVj8fZ5HRvs+arZLPrgPzpVhIzMBA3q
oZwtQ+5zo8fGI7DQ2KnHPsB4Nd0EZhDrr6RqngLm/hBNSTDjUBIQISSxJ/VC
a7bCk5V8RNtIPMoI7bW8u0wocFrNvF4JgAP7zfTQslj8w6MnvkQZ82p+9e4C
tEX6E8C2nHug4k4DlCTk+JMHBmWKEsA2eC3ddmJ9opbTwEA03HHfwyML06tZ
QvFCr3HWLijL7AjWZ4489BG62Qyb3GRl8SHzLEU70KT5eHde4LGXHlNASlrR
pDBGwZfK34ptbWG/1DM9rnVWk1BJlcjX0JahhAqQ0GIozmrmnMUxKD9pnu/R
2b7UyRGsAaEMdCOTelxh8CxhxQzJOvVX0eWZK8d877ULN0K4jEN06hL97KMy
adSHr2M4D6MCcWW+ZbdwQw/1I5+u1SNgz69P+A1mqmuXHkg5xMAURIiZT4Jm
1TXMBumANFItqE1U6H9oiovQVr1YZ/1r0b7Pf4q8kmIrU0wtgRgJiCgsz+Uh
WB/6puYSXxZsBxK22m6deKZsKJ9Z15vLRZ6QKytFBh9EkXpaZfmuGMjfoVCY
HBIO1+/VGSTo1U16GS/FhaVoBM2TfqQ//JmRN/DvKd3uCp3i4gp/Tq2X88nt
QTrj2SVR7KREvkXldh2LuaTZZBzZhGZIf+kSAIavS1gQe8EQbKpy/5OpvvKd
gySAq8AWg2UXsXFmrl68dTgzCnPJmlsUkE1F2NnWNWU01oa4N+OEY5D5b5ny
uj9K0OQzNzMfBh3vFDvWbhbexagmZEZTbNEDta+pfPYmUGzhJ3KBfHqSu6NL
wK9ebAtDoNXmUULPyNQmuEdck5Cqfvfwev1njZRvQlMDyeeV+hn8/1gcGrAx
FJiNdpLa4E/+LVyJZ9oMwNoVYVjkQ9oqSZptjd+5vjw/+WG6VybF6p3vKSAt
tq4vvA1VUyIsouUuItx/xcGNHMf6FzDTSMtgChWUoho+giGyuZ6ofoxgqO1r
zz/T9xq10v5WwCDuJLZap48+7D6CvkUF6cGfA2nJ+4H62+C9g8Wc1yXaH1Lw
Ywe6qbfxBZ0m9N7qgb42FQ6zrtbDnZGsu6VB9K6zmc/+tefBSWL0GzrwCsqm
ovzpBQGmWBBfcuH22wPeUYi8L1LLJO387oNuwgf09qEgblvph8WMkPjNkbYr
FEU1K9O9hpCdgj10YvWQO8DtUvOr1x/SDmZhic/IFWN0a6yOFdciscwZebkB
DF4iIWsERIzEG6KEQE1ZKwtebEzzTXJVHcoG6oUTEqlIA0DEd8d+FcCBRgve
f2IdHSbStpXITRR+P+Z9YYbxvbmzFXhbWxSusCGUz8lk/onM7Yslgaw9Oybx
t3MELdqD7K7Cov0jq+9hpbQhrERgoUzajHVMf4Ye2/F1qyqZC1arCgcYx5bv
c/VPEVpL2tUMubvP0s8StgYhPjN5dUTuP1VemNY8ZbwLMba+Be1alkpj1aTW
4qefu66BTDqBC7b5WHRx7RsRe5mBQ6laOk7GysKax1GiSFi6AjwSGUi2kdvp
kq8+FGq8zCE8Sak/m8BXQiDHg6N+lCzyMDcGKIX5YkKXlKXV5Ccp/cqNIaGt
xh29c9FAr1KhyM2aXTVaStkPKnKlS2UENohu2o7qlhSHZYoI39Adv30FSck8
shyG0ertu0IiHEXGWTQHMtJewG4SPiO4Zxfwh/vnGTvuFsREKJyxFEsFPw4S
sasAqj3k28rpiroRAqVeYK3qfTW0tJHNoPw2ZVvfJ1LBpI4fel+eAimVWtZv
AQbMdbCN+JPZ974ktLJSFEPvChDLVEac15Xkn2Dhs4aAeBPFzqeXljVDzV7w
MM6S03Wwh44tDcI/H0BDieB9ILLBp5OtLgW4i/mG0W/nb2WifsNPtPQqiEkQ
I8ntcaGgq8vYV70f1WtrskVgMfHYuQKF+lfSodila8TLCTHMyhlovx6f/+OE
MxfoRZc2O06mRo/W6H2F8lqiUntre/gFFh95ewexRC9Rtnqv2dwIZOWqKlyu
MTLvgq1vXKj+KzGRyWpUtYOzpbpNrVkqI4cmQ62yzsgemyF6akGAfgfvFuJz
BH4iFV+EeCAPjyGHMwscmNpCzG9/XEjWYsHKXJS1RD2CEtCNDxjOJQslItDs
npmyYrQ6Jk22y5gAVvK3A9yTyUMUohb7JhNUqOFczin0192OC3t+SqqQrm3+
SgYKNhw/IYyyl2qKInX4aXmcjHZ5z7Z5KCYtrKUm6umdS0P/zdz+tEOesejN
EPMEDJfDYyKCp3Qm8tzUHOJPURzSKtNvlQols5nC+IZ94HtC+WYJ3nwHEu1w
Zg5T6VE1fQhUHNapPJdY11OHC9iwN2+7kDvPbanP6LZpWLGQBryJwofx8Ddq
D2IeskjMTE73r6P95c+hVfz2c8M9oGnJbNQq31hf8537T9V3YMN6dEFBWWMH
O+ga38ZeIGrePX92z4N62DNqq/mpIG5vQzAbnZoZM6y5sTjvbSwFifLHrOsL
arU663krPsFhu4fGTcqrayoRbu4SYcR2tENNgGCX6fhn7y7EtKSVyXZtpUa0
+An+zXVeJFheWwwGBZKIDCcJ3zmGadaCVu8jqCzCNrLWOg91YeQgOpzG7OyM
dnpASo4+Uph1u1m0TD1KXqzGwWviFvN44PfyDiGTS/Cly2T0O0aG6IZGGEiJ
oj1mQuWqdVG1p/TR9NKS5Mz4/ge7EFOyiP/IMFE2X03jcmpci2ac88kgROPI
AspcM8mnR8pRRj6hX3kFKQl01QEGa6eaEL0Pdd5S3DZRzmXIxQw5fMEy7v8Z
6pqpOLY9GH0jFdgz/1aOoq5YuqGispoK7NevkUXOpRcw5DPzvmA74WxibBdf
4oZafYpi32ZkcsThcfhbBy6DDSFY0wkijGk/fbnz9PN64Leiae9xR0CNbPen
gkUA7qFAFXnPPvqeSRNo662CG0aGEsp03cRoycnVKltnei18nJk0uCNQYbMk
WYrzhI472j5wIiBqFRnv7u/rbPCWSP9f/2M939N3ylyfXZbxeXM/Bq5mqti7
m5EoUAoei6qGfIb2PkBBmJJArGvHUXtT3tQmPYVu+jTqOSgMMuhHzW76+/Bp
z9p9+3StCg8NyU8MtKmtDObjouEZSW2Il0RWKB0MHfPfeuUO/bUyjnJKlc9c
iShYo85NbO5KEzvzZDjcVrrEdR6kP140d8YY3eiHZ+3HZC49cSiUswyoPbYD
Mr7Kfh49+34GhZ1E3dReGsSznIo/VkWSxJSY0x0t5pkkYLNQTWWvGFblSqgN
eI5MzkLuoNnn4Yiv0JqVe+d8XiIe0a5EEW2taWLfj8I8NbEBGiuCvom8Cftt
YOUx08tmbB9fxlVEnze6orXoOJWXpyqJI0LY6nw7nOR+JFXQapIjFSUglJ4p
Iu9JwFvRcjpm8y9qD1ZHvlLSzckn5dHDC0v/ZsMLeZBgUBELptl75NSgJPu6
XNiPe3W/u4nmWNtGYYXW+AVJm/vHApy1OmrZeAcLQS7aWqRvQBttHJoBwol3
3OR/+S8h4MtzSxBtqaxyK9yqCP9NPjR7NTxQ/m3NOqJQb5dunvZwEuUDACXK
dUTw2j6coZsPTdCROw0AT24sv7LgBKETbnZ8QexjC+8rZlePD9bPaEJKjjrV
ujgpz1kQFKPKdn0W8c7LNBLc4CtXqTTJJOQcJzTmZaeE8SkE+fT+tMgqAn+M
ZbsIZM0PYqQp/vnwbtgeFppo/gm47/rcv7if9AyqUGNccgHmt9SzPYbnGNXx
sYYMJygMqUOlC0qB3uFlsxi46r2Gp697jSlzeaMKM4dPt8lHKLoVGmODP9fI
ZrD5Ko3shuG6AY2b8sktK8NZu4GYrcbzBTES3WNxv7P3/UGKQYQhegdXi8CA
+yEOU4Xyo77ZcnlPRTS/zyUAsWJ4RIs8+qYshdNpnPXSgWYJ7mH5TA6P8U8/
85LGZlnti3+4GuBXrXNFBKaZZJrtTfnzOgtIW9srYJrgBBLp2Uns6R48Le6q
KvpcWwD9Y1xbXmFel0TrtMfBotTgXD0CsbKsXpEW69AP55x0FXBxQnND6pVh
Qy/q9yGZSMBzA+jnFiMxI/JcbVJg1Qqpg+P6stZjho3o4LXiv9rGBYyyfG2h
GVFP2FvxHpblH3Y+671NEXbzP4HUH5X7eiEdDnML8NbunU7bA2U8/qSG7Gwd
VJNZqutDisUZTl2dxuU9A6zqxfWDkkfTWU+gQZsjbkWmKDs+dstSPiM/O/rt
QMo/zU4L39+B+DwfaTYSI3DukBYxvIcDvgyr/rQ3YxA30XXonQ9UJqUk29R4
sgADqRyCPqx9oj4/qVeC5PTdIbK9GQ4mccveglSi6kIiXAzeCEJHduKEOFL3
Ue/sUMWitNfiDAAP/Ac9ZgQ+1cLhiOjQ38avf+8R4m16T3MoX3Xu4q4Htm+C
11Cf+o8wdY3G6hVjI1qBppRGnRwqYxCvyWdqWbCL5377uZPtk1/tORbY3j0/
Z0lBZsTr34IoJ76Vflx4jKE5ySQ80q8n5h7v/mXpguAI3/D5f6B8ocaH6PLk
e3IxhwNmeIiqYGSKJ2X/RvqvyqNMxaF2kr2bT+ThJ4wvUW7XrnQCUFAhaFbU
cv5WFrSYNfWbuq53VWpgBqR7lveSCLuh3/ytqPhOhfdC9eljU3rY29aOkEFL
TVEDdv648tQ9PAdv0cdxB4k/0RT4vdXozdolZmz8/q9bGW0GEl3hLYaZGMxQ
o0yVELGIKmGqlzgcKdoCA4u6zPrf3IZNs6ZeL46HxHHTJAD96yATc/iOHqfq
v/SVyY2s47vHz5nNoO6g6iQczZ090dPnz1SMwwFZZ5RDy+D8hYSy/9vkFLbs
a7BnurnLJQjYBGe7JzqF/lZ2JKfUuwvqTbXBpDwW2k5ZK7Zh5QyQAGZUQqom
naTMeUTFRKez/cn1vG9FIbrXto3RSQPx+20R2RgKBNCiBM4C1AZlN3QZOUQB
U451oRg/D+W9L4z4e6GYYEFKcrDVBixYylpGl2YlueBlp8yXMgYRGUoNsEvE
088XgUT4Oo7axLWazxbBZJbT1tWAVUnmyI/u8xzEOuKXZfNQt/6LQOW+BJ2t
wcnXI1nXIevKc4kx/F0Q41L41sOQet0j9XzACWOpsPhXFAL5P1j1oHLgeJkx
wCQneaPUGCCMXIvCAoLsKJ7tecNezXUe1inGmgYP5ZTp6du9MYTiHCfK3tYs
/dg1MKUB1miAHjWd16VE3clgVuqYctz9DbFGGNBJ6dK/ciA0818t2NjOr6ih
+SHNkdId46ty+mGJaJGmtaajizEkpWUl5bjgyE+rxMuMfiE03nTyoifCLo1O
Rq+hsv9sSM1o9GaLCNTZW8FxkEa9Sfk1mUldc0XkTxK3jyY3V58bMqiiD3n1
x7BQE+YbZpEbWOA22fQ92Prrr7xBe78bzGXf68sjxCYvkOylmNbpJWXNEuM4
dD2Inm+nN3T7uUQi6Mru8KVw9S1DVcy5VEI/mDFVQbZdOdHQcVy+0qJAXHBV
/LqgO4F+FERE5M3EoamiaYeI7qCp5wPxJf2NUYNmOB2VMXEbuVc5Cxc7ue7Z
GScTUnNiirQuwVIELH7Ztqa4mlto8EsTF90neuxJQgfhNgEZPGWQSxKKguSi
a+O4hKxR3MYvRZng7oEYKfGtlxqRA/+WdG/j7nVnKkliSC0ByFAIIjw2caDe
m+LpG/yb/SPtHg2sHg6TojTviMnVONgLA8DqF5vtq5Y2RdmR3qp9xX8YahuC
9P4EgQtIu6DPilXefEuFMDM2DQYeP5Scc5Aqq3L7owPmEjEQ5pxbeHpRgget
lp1YBOfkuF0dgToj9/F7oBN1bjolRoT4LQirMtofmX/5Iy0Reb7QFHHNLSKq
aSaiZQdBO/hMRoBu0FYcrtuP2W/7/uEjJT1xbk49Juo9goe8MTI2kHZwuSO+
sFTIFfAb1EcEMZL+K8H3flgXwn2LwEOlKu/mYR4u/U8Av16ktKADKaVW6Hgi
HL106W2sbcZmd15vamsEWX67BEQuaL94D1cPHNLEB7kvJAIQs0AeoVzRKT/8
kokaf1AayklhNHlC2Ieogv3R2IZktrSzCGj7kJqkHMBQ2NWk5J8aU/PCmmVX
RuI2IqX5SHaQWtA9hOdtB3FciAJupLQaNiTQ5vOd/4Uy/b5rSqiLAJwSeTJG
OMiaQUGsNGwAxexZagl6fRNmheXDST0w2rmoT4yvgLgd+UkXhYrtfTswyNTv
I9WbEOXUoWret9A1v2VUMd/EXVBt2LGy9NYQJZmZnnJbsM5dLgK1tQNO8A5y
H6bSsJzckO7m1dQS6bUM1rOstLvQxU42iBVV1HFoZ3O0qFYst4Gs2m+G+xWE
RtcnerbyeTB+b7GdnSLBpOuN58a+ts6pu5Lw9ySNIqP4rEtziL8VgV6EIB/Z
iwX9tpy8FKJWKQR3Dma/zPhi54Db0qv3NJNcgLFM008ICkYVfQcmkCPshWCu
NE4l5X1iB1QqXZ65pZ8jeNfhlte2D4VSfvdXGsnhEZCoCXW+cIpdZlUMFNN4
AfDwS5XN4AipVg0XELaQ1rlJ1GUPnNZ91Jd2NIIzmUrOqmXRXyUZAc7oyfsl
W4dFxS6e1xti9PEvKPTrCfqz3ENxJbDMOi85ufag2d5mjhd2UA4wYKcAyoHy
7geu9Qua2aeBI8Jh2lks7kKgeWiEVDup8A84CksnU36VoRsBRJvacrTf687X
a/+RKzc/SalD61UYRC3xtog+qqSViEHZI3JRSwskaj13IrVS/9ViD5K45LZc
vduKI2CRoHcyZ7UOFuHUfsL/w4PZPq8q9HZDIlhxC4811h7N6dXM/DQ7U6In
k6DZQWPa49pgPjsN9geXQyviyoS2JM6c0qXfSZJKUw0XPu7vhkdrojOkC4dj
TKe+jV2XuvQKZB8lR6fF7dRzjmOXFo3O6kdeRraXtoFGvmlSOIaeCid8vfjt
1KVTFL1b2hg9b4tuT/ny2NMWYo7vdTyACjY+Ks631hxCfMjPV8XymYpsVqhr
cMm5lqLqFSM+2Cr+RjvSx0CzloSEmfX3J7HOrogd1KBVuaS5NnvY19Amx4I/
TJOJfazraFHjG89My1eU+v29anGe94MR5FWHeTb7rvoh9xnJHDe0XcclC5X4
+u+5+7QfDKSXcm/OWa0nbdhP5G0aPX1EbHB9WAD6KPIOA92fYs/7aGQfaSSf
ivRUlXayM99MMgYByXx/D4bfMPHZU6EirGcQdYaCsuxEUUxTCUTJC/69noyf
ReN383T7+5U0PclfknsJAhvGNrZNX6OhX3kpxz45oXKDXH/aP3DPoxheHJNI
O3mpvQygtLFYeCf8fSvqOOkfPjix2qs8pU8dweXBzFL2XLnk5Gn+OakZWgGW
W9GHvzKQXilkgVtl7GuiBicg+Jd8IrdS8VFCDHthPQgaUa/mxdwkTCvfJo9J
P1USEjTmtu0AX5JMzbsTE+weZwaQAkbB1zo0fH9gyZPxeWCqyaIT1luTCVof
eWtOstiPARiFvWjgyHLXkre4T27TVY/gVEYAX8km4d055sY26G3a8zfMTSgg
gK+ok8fSYnUwGuQlvPF3Q7QQPcTRxzDiVahiF7qT7hlagCYf14rKNgTJaG6/
jRCXJ76cerX+HE69kV+LbRodMP6EsOuUKvJbGSKFX8ssmHyHIrCTfNFOErLH
jQ5nUDMNqQCJrXd9myOTJ4AQaY9ICs+S0mbsJGJbFd9CB+mMxuWea/jTkfZA
EEcVEVbmRH+7LJ0j7JAwqkkFYcpcZUCCJoagJkgMacXqYaIRHcxNHm+CggJ6
nnNxSlQ3pag4fDbZqUizN04eWNL1dJk1m57Lplkh8TdWalR4PrFTvQA0nNdR
pFYsS3vjby6KehRCAuZXlQN+dkF1V0iMzRhTxd0n2oBmEvJ6mqyTS0mfIG+D
47jVc2+EUx/L7mr2osDu7Q/x2krsznEmP5Xf79/i1v6Z9qYvIBRPztB5xLbY
1ztmx1fnIuUhi4V5r0iMdUauES0HS5tWvVn5Ner9ExQ/Wt1MdQdXg/ogyJFs
DAag/1k2SHK1t6JJaElgaqAheNg84Akr24JjpcEXIxeatwCvbTzoTaqsTsq5
SoMy5BtLmUSDsHzRAfkFZ+AMcbLRbcZVWd9CHZpDHvNdbE04iT8CwPlfD41X
zPtUSgm6fHAPT5jZLNPvEpyq9wTngsOZB8cUfBTKCTCTkjxhIPDFKUu0TtyO
QaYxAyg0gD0pAk8d1V9tsQ2CjeOJmEQe+L3q51RxPt2UysvwH0A+DHWWhbRd
kI7P0SScQRI+iz6c2xLvw+qsyjQOY7Qf2Dkqx0HiQFuyTz81kfbTIGUQQcKm
WmrJFJTsTWFC68W5ZPVj2iYw4MJ/f/2BCIZe2nkTfYr8xjI2hr+9n1fUNNh8
En3tlmNM1YVomHwXiGif6B3gKMry3I+Vzk5dfn4clTjVicRdm6xXSNtWEfL6
ll0qvuisHWNb2AjCsVB97A8yz6qdK8yduWopzn1jVYFAMtBEiCRPda2eB5RE
W9c7MuOLKdLJp8rtrnGhVsSZaSFEwDpsWruKW9oo2HFJJwyao/gUOQDCHsst
ogPjhYJcmjNk/4dfoAVTrMBp/71/my4Ky3DwddekM4Ol9zfd1YSj/YNch1VW
3Yafl//d6WPX0dIHFjXJeC0ItkGmtJSSE9cDtyyqVXeCY8n93HdRsDB9OAil
QD1l9rhwsjFJ2Ds/1ekMej1Y8ZcaJPYL6596gp0Lz6ImujQeLvZKqoa0H76e
YeMigP6DHV1TM7rG6Bt8ASsDtBuiLbq1r5Rdtjko11Nf31ZrAXiPdPOG1Wjh
1n+5AM4cjXx7j7FawMYGJD1pLqSrGR+qO3KcHOtZ/hJplWyJJAkRC1WutUG4
21ph/inxtzPwsWFwGHiQ4jNTkKTuELoHkht2Xw1O02QlmH4JLRrKYUo0u7x3
8QPFoI1qqMfLUf8zNdpKWmLkPOk4bg7gtRhKzye9U4gdNtKimVGgOynVUs9+
EOW53QnpVYBCU/X0fdpl1MQndQY58pdAgyp4LaFe6bVgHhH0UvFV1XcOM4Cl
zIIzJnFUWrt1JY3UkRPEiom4am1/yRd9B3OELXz7LqyvzmNPE3rjAW6EFLP0
/hyg6/c35U7oCHH14UDh4SFldz4QoMFGfALm0w//hfWbJPlAaxqZGrAAxs3B
eqk81MQMs9tfWTzR19nKHHv5flK8e2oRh/9nisyeSRJkQRK+64Wiw28vXE5D
OuAbzd6nSsv6hIz20xe/BbeLkGOSenLZwGgPxxDpda4qboWgb194PW9C4ntl
dbxtc6q6hExwy533zmqyvd2RIAJPMzj+ILCYvOQhB2yHpkiknbquQdJGcuM9
Kg0W5y9O2nj3lcPizf00jjq+gLDySb8JhVp7lClYAalvzz8e+2TvmSmy3mm4
dQgWoU09MpwbW+1HtK2ZitubweN1ORgLD/AWuKYsBVGK1u0QLppfpPYzFeLb
Qbz+lCFGHLCwGJlYV43bRxlRb5OBk1lZviP6LPZB5NYeo3JcLgwOchZf39Jk
J7Hp6d2p5LMvPsOvd7OkkxPSx2IPvPSxvbvBy0WjQkmKqaYUdLpGgKevnNL/
OpTvKMp9zN8T/LHapfGXY84C8Hc+0MEF2iV6h+K+OMV2ptVbYtSwmwIWMxDf
bHGuv4in5UNaiII9tO95RijKPzf/QapIRoZxF7eOYRQFqEmWcMt5F46/5BdM
zidif5ORaehSMLzOvFRmlQpcnhixWpC9bK44rsJ7/PLwYdU7QYQDOuJdh957
E90HnWGoex2eez0cJza5QcKBTD7Rsfy15lFZCOw6VL7JCCuP+4nWhSHGEH9L
RaXbG3BitHRCyXmQbvehHGm+66dk6WhoBFTjyIZlZzpfZqDKXGO7cZBNDmcZ
FUo+Cv38KMcBVaPo7mV5k+xD7lF6ZyBb19qOtjQacL4G3v/IULrEam18Ukhl
geazWUK3+7zopNNedab8tf0u5urQIlydtWVITFwTEZdsLl/JDDPvAWp5Ie+Z
IqmVOoIIf1pzTcoN8/w3xASY33zNe88HMUzYZkXAm9LTQ4miyWyep1BgSqzI
8BZRPb9jFub+eNkz2C90sUK8td5P2kPJogIPB+gLkD27TTsh5UxBrPxaBKV6
T51ibXHDS0XmgvUSR6TmUGfqR3jRQmHDrNB4LtxODrdgmv1oSC9jczqggbXy
k6HkkhC5NvBtzQWttRBE26PBVzR6ogEw416QfKXxmgPs6b66qPYxrUgzelnQ
V9eifHBtCbksqaGbE2lPpfOeGM5Fe60xqLvfs11f1Y5Dap8XxlBhfSaBsxmO
qrVswU1K613Xid+dcMmXNfHOE+351X3/PdyxP5+/EtnHBKEuuKtVC8/R/6vM
lOLwRu1mgHZGf0xl/zVmdI8lV/1M07v9WDJgby5cQp4r6nEmDfuo5YrVVnce
9j51ySDzxYC4ZfeTQza3i5s9gMZuOayyl1anuqaqAjinzactuuCtSXKByefI
vKCriHfy/ILRh5EeztKd8z+gbRybU9oTuJQSpXc3N4XVu2Rq7zK0JJHK3OCQ
4Lq1ll9JNWSan7NbTvBamXXiQHllM8IxAH4sQQ51JIVAbDeR7afo4mpp0b22
7MkZPpFyK5GHjE3plfhSiCDvJUY2/CXeDsFWYdo6q+zL1ScJZ0z0CuJkZ1dX
RzDtbkZAGusnconKBLfoyQR9hI6qoJ7ycvgcUssVJhKAWlylsfcq5qHb+Cbk
xBsvPbDrrAnm7xWapTNYWDeJACeCuInmpIaHBu7h3BHLJWkCKmqINq4xa9f6
NoiJmv7QpayVEll9dJMFa44cVmnas9epY6bMm2oSHiTPF2eEZicXDYzBhfru
NM+tdkYw5OPrCrsf6eN6ETY3wjjR1BQHA/1wPJfRXlzj9SEhkxOjJsLdpBnX
y5NKZqj7EofRezogbCKbg5/4ZNWheSsaW79unKacqL6ZSEJDbwzyb7nn2K4D
jLyNMNEQUQKxDULe+ICA0JAx7o++brFzaU/S7T5e+2eMUjK6VhULoETlhO49
+a976o6NJNigRS4y0MjwSCCmQ2cgytiOXA/VUdCuCr4tMywMThCOhA3cf+bf
wWmv/9XBth4ZXCmesH6+ALmZbDQUUQxWhSjZxWvc+c1jGwbWXhH9bw7sTwwq
hzq7uzm4+b9i2fWLhDlZvMXYuE9gLH/D1pEr5henk7F1p6tHBIDDNNb2eVWr
yxlDZLjg5PEIeyrYptA/MFLWGtYtEmrfYH36PU+E7remUcnVe+XM4SHyqlTi
g8TQlnjpQYBzgIpMRIT5pX0DIqNPw54jtP8YxdtNVwRk4hLLJpVu94KWjbx5
7qX/lNU6fay7kGzf5mqo/JInC2X2OrMPJOYypbNgbg3l64MTe5ee+inAJcGy
FMu18YuCdXwkgJ/XVgYEbJAMTuTj90kafQteNPYOF3aY249trWuHqIk69926
lAu8til0+LeX8jh0T8KaLZ8Jn61R9rrwjHXJQszOXJ0Z3VbeFkKTf6fKIMd5
Jz1CyEvL7/Q9HXPbhVuIjd0MlnJSOh0iKalXyFG/S0qXnj6T/2FxTB4BCe6k
0cwUq7uG21RTbZGpbaMsyNPILLN/u9ox6av8wFHmWpd6nwrXm3g8wJeQ4JPj
g/zuO1uvir/vEWul4MsT5mT3VNkk30PbFRzDxa1hP3SS+MnZqoY1tnCt+sZ9
Abnz2X+dIfRmDlr+YySeF0r4ZDW3qDsSoSZeXmtq5D0offYjbk12iAJJmfj+
WSeEn/eu6yIZQP1mGy/w6rqQ0LGKH/SLIWoynAoHhiUU+MvULvE97M4B9T1G
50gh/oKi2Ekpv3cIQZNB4yGv0/o7LDc+eqyjDueZnQwbm+3EjkDELZnU5zyk
ksMm+g/JgFzppyI8GvdG37EsKzKCpNaPlim3cC+w0CZ/POBwaAIZ1BMVT1O/
GbHHRjU2M58HNIuRcWjr9EaGECKttKM3UyEnVpiDB9lRz98+zXDC6Mehn4He
A9zvY+ecz9GJCo7Tnf5V4Gt0d/SgAV2nSN/IscFszf4xBsggyC9fhG1G7AMo
URNE8VReomLp4etY5fuQbnv46EmMBII5P2LLtQDzpVVjA1xtHmrXUQ5PjS2C
bnVnXN1b5yd66M9Is7r4lyXD5oQoIsLB74SIoZcqHqQY6RusbpOZVDI3FmTr
5mFLrY870RLCj5lqBQYl4P1kdDc+CnxDfQOM77Khreo6yW0kknkDprtRLi6M
dXcijgzam6JyY40qRww02n3GWHsN2HrxQnR4H8gBFYFGkyl745/rTBQm8cEB
ozFB0LMY1Vu7yGo0cfsfYHUBcBv3Y80VzvXzAG7Dern4PCa43qBzcy5IhRZ+
gUHURHE251I7ZdpWS2dPdIReb7oufIQhCA1s3IscVHLCEECJOFn5GisYnJpY
DMYDm4f6Ty+b0TLj4QQVV6gaJn29MyxmBxr9Y1VFDQjy+0iXPqyyxoB2qngk
lgkLU+A32TfhuYlgOj2pFmh3jmxksBneeORthWc151vEIEdPlAFKWip5iqpu
FIq+/kWqkb7r2LSc1cqL+KbCWxLlZhkOIlkuMfi71BD2LxgoGYeR35usfoVP
pImnRvcIAdyvuiXXfqLkPu/FG/mXAjI3RDmSnwMFxYAIa+sbv/sXx2CYy/FK
q5wHOPsaWr+m5SLih2KQphLBBj+ZYyzYoQhst0zp19l7NeZff1O6Bp8OTAty
qWBODNNLVZ4CdHrF4L6PRB93JHshrpdUObK09PCjsjIe8zmSDddW8IcnYIRI
lI/sxgKCFao1WqyENPyNnkDyWWJAWA72Bfsy//otq2XGtrEsrV0QeZgzCT7e
a/1kAOjG6EvIm3mJMgFrT/zPJxUSk7sRbpwEQwsHFHbVAhEgtJ83Hbw1VMmF
FhJQw5d6qt/oDZYvM7LIEHquPTd8wJO2Eyml4n5F8wbsV9vbbd7c+VGkyWhJ
HZ9dxjqzV/BzxdW3ROncvPgsVZH5bDQ1Euh9CnBrYPoediVfWrcdrIFo1zpS
nHJ/VLTdxy61+ATKnvq0+GiM/W6Rrn1qIrCijg4Lj9xhqPE8WK2X/nI9mvwB
yTTLGIwuCFodVwZH5BEEVNkejMRmNarVdqYVBbUUsZwGEStsVTM0m10+0nd6
ge2GI1UwFL4abiobDqxPMmGddm9Yl7odU9YeXTHxwSTCFdkZzAnLeZoKVn1/
LbYPEeqfSa/3ez/DJzoy9lLy6N1aEivnpmgBHDqtYCjdhPFVZnAt+9/2NbKH
1Jk7sGz2w/Ccn95GL5VXkGucf3r+AWMW+xQ8pKar1ui2++DPsMcZpCS1tTtR
tT15kmGkq171gfqnHQu6dlYqzGiJWqKAZ7m2if5cWAGnaau1BKZ0cUGzw1yy
dq3J1woKnr6qu3u3A1kCMnM8y7ihUBRp8jmaH4/T0DxuRJ/aGsD9gqfkjgiQ
BOZS45ch1GjrRYEG1naiKriR1LviTWtA+jaySfHGa1Z8wXzhKXM13zd+FKuM
cRrRrTXzQLzidx4/xXOGaR0yiWAWaTb1NmA54OnG5n3QObYclCTQoExVzY6A
Hjgl2a6yt8ehLRqSckaR377NFW7F4o8UOeQnv/lJd8vobevfsl/P+GevoqhN
IeWpPNod6Hb0iLVP1KSEDsfI0HzYQjCIRbf/2fu0ZZLQAMTIOxG6aade2xUG
anX3KtfNPkO6bavfz7qo9FPNNyMZzNM55tEceb/vkvMBuYeTs5X06hBKch7+
xGTPF9+QDbEnsgM1u22jo18baMuBAWBUKgQLrJXpxfk2FQOuScMKEDX6bgGE
XuCwlel1bPKIFHdpfsDkGWCKrMrmMPt50YrPvCB8c9zyJdxSd5wkHR4vyb/q
PmhYBesG5ZLpRINLCSfRT60yo68zAk+mvMjvr1iyWB+xyiYdiGjXUjKWjdKD
Ur/dr96dPFNbfyHTJd9I16ebHF69wpEATFrEKok9EX2m8HvraZnaTBBV8fin
admEZgWs/b16CAq0fzMeujDmPXyB90MlnXQvo2vFcnSF0CHnL/8ZWPXQHpI5
Q2OB7PPeNolQsxHXiqN4AqNOT+L/Xp/3maG+7FyUd+fniZB+2AWeVB0PyvD1
Fnb9GjRxzx5/DRkScnm5LYU0V8d10J4qewBaaL4DNmvV2Dq/W/ygfWiUgmwP
fYLtKnwVsgRTSWa0YKIidH4PpCIfKwtZIELWkckh9hZEQEUZ+1EY8bhwya1I
Xl/+QfOhLkk2DxaexFVgmeJGj3Xfso4GUQ7D3W8PNWsKtW1zTVwfMM0VrlnZ
nQKKk96b9lxL/yDu3j0cqe+yR7XgZ1UoiLk3On/32KSOYSICZyMbK+4NfD7M
5YXd1acaZZKp5RCkx3g5S5Tk6l9Jk/l8//vmx60H/KmfWcfiwEdCSAUQ1acb
bEAmByZEn/xpj1i5Du7qfAzm7JwW4x/zS7F4xdg+5aJA4CM7LvflPGPPMNle
OBfC08fcP0687m+QcAnXUN4Zb9dEaZdMf+dDv+6Ip/ZFLhOeXWYsHm3UkE4p
hfv9xKZAc1sa3768ia3JYAtBOJ0ssJRE+Tl9ntZrJ02WfAucS+9w6yraEhMT
5PrNTdc+dUPsFChCOJNHj/GL/ARQDugbE74TvssU4HZ518icVcLt917WgOnp
rFTnbYW489SzIwZ6JviQIj2G6kYb1O5J3Xe9J7eLUmSBDOogWaK9rg/IJirU
eNaq3SZyHLtC7bQM6pGbFjIsP9Dhxpuhi+Q7XL0eKDSx4MEB2xXtUrHRtFn5
jn8CzyXme5vNKk29+C2tWCKcfBBIATpVW63w5I+YVeK458ycrYG20mu0H3pH
EtFxMRD7sMNh6enyTeR2HJaFf3+qXwxb41hZi99h18KqM1KHUlv3NQC8mkV/
zpO3wOzCejQyhptlhuT9B+3eNAHN4KbpPBYIwmOqH6V0SpDcbCdnrG2brbNc
hDiGuRtlJrpdViwDzjv0mYoNENnllPzOvRJ3/LXZrDFg5PLHGsCIf2n4TvF0
bNpd/PRFQ4ThNdpolzZnqTAFIvFpPIAunoGKYFmlLeefF30mpTRkQ1PRRBHC
oZmt3gbxwJllcN1/WMwJbENiLqtpkBakhPlkDPYvGeGIi417cQGxEI10RFI4
UtpwtldN/PLR/ZoDsPgHQ1uZvbNVQIwEIXwLQKZY6XTe7+Jk/cE+fzVq5HjI
cq95UF+ePPEpPPZCasQJRevUyc5etba/oPqk2TSSTrbLFk2UYr1waQM+hcwo
wzEk7ZBYIPwJEibR8f2kQsBDQZKUytgunMB8MuBhs6Mw0wtdxKbXAUMl2DDc
K74Tq2emP2kdKfo6+laQehWLy13EbhiwClVUcY3gMdgkx+pidS2yItwDkuIr
OIGhkkBKrl68bCBd7OACgokFumwhoF2qxo6j7fpvdgjK16yq/FP7S79rm1YS
M4Pm30IEOEEUf3xrVUZAIIicD9YPP5PzWe1R7sHCt8knd4xnkC7JBDOyvnDm
TDOJuI5UNG95yOk73ap9XF/M20K2hWGyu0oh9bE86WmzOJHMLrcx8XnNoq22
o1GGB7jgfBrj9W9GnHz6LvwUiw+vkCUzTVFA36LWHL+Z9aBa2K7oprAXQZDB
6AhhdqvTjPhhH/fFrMdE+FqAKBxnw60DYO2nmb/SlgsJDmJl6mMcwCUetoAT
n57QTwH0nc7FeDKM3D2lN5gR2E7kCoAIXU6p3Zvz7HQFPkc6H/sb7WyG+7V0
WccgGCZsERBsyTumjpNzLWwuHHMQk97PUEwz0sa5vBWb0dtkF1OTLWWCmk0t
NfKN8i/txFh4re6BEcWf1yLF9WKbTaZ8p37rmCL9YX+Xo1Uu7AS0V2Fy8vrN
xUX3bHwZVpzWPnRQ6XTB8pv0wxClcGcpdeKmHw9K459N77xtuDFY2/8NmOU0
dp516G/HTDXlfQU+hICrdtQZk4+1Id0VSQsj/dSBwxGCA9QauKGj8sq7pCVp
LWGmDTuOTeBBOG8Hxp/dzyHS5aF8RNeVerPEAT8t/DoNnSoj70GopxjaoKxi
Ys7w58hULydBwMFxFkWatAzL+ZXTX3eo/tf4GW4Mn1YGmxArCPs4hMJd1h32
zUymYEqdinR+br2kpbdLIy9dWhR2aGdK8kswhWsAjQSQtjDBo8LvdjeHg+0e
z9rBldYrOLFbhl6qaTq7O3fCBXSu9WuQTHc1KC6vuY+5uKFGYIxorJGNWlag
aIcmsPmksP+RrF1z0eN2Tzi+S51EMk6kZVsFAnF8mO1JoZUwh8C7I7DbhCYp
DxCfthwChEcXiEi2jW64OfqNcDEHKB+apML0YnHhBSc0Y4AAUdq1R/FBF4JT
+S9EODPMgzeCliosMztzyRYcTqvSFs/NtGctBCk8S0ErA7/NrZ14FU5wo7fH
KGELHsfMRapUw3jtkFdR5BqntBWrJ6QNZJauVDugeP+trCkShUElUHvXG01N
cshgx6B4E9FZLYyidnT4To1n/eUn2mr65ZM4Ws4PK7sWRLJtrRhD3vQgj3rk
wgZ/CY2rwA9jCKhbooo/725cU9Afyg0YWdNCYi/9tDFsIYh459B3gsMTZ8tz
gtyADydCyxSOcJQaczg1F8R0AEAZ7u6gBfkDWZVhku+1WvEnKQFiEIs+yYiQ
bMAr2iD/StpgJqopHz6voZud6C0i2LO2iz6KJS0Lc0n52cb97EvWhoVPjFWD
+Z67LO62cHyqM/DKZlD2GswajdClRATFL7actLNTvrkvlJOPMe558nRyny/x
DKhas6YIfnAl+ZRr8NiZA/Ecc+2yeeM4kOOmxJtp2PlkHx8lMwx8HBdEId2e
UkcuWYQqh7oMjKcdTqBmJLQIGfKlcTbhzzhNUy3ecxOHH+pfmLpt2ndCJfcL
LA09KeDlt1usWSHyiePBXcE6rWsVC1nJdZ+CSmdCB53SoB/1mrF2WVzZZrIY
KL/K3aC7SuNpQI1eUhTuIsmJwZYxefA8b2aunE6aiVqNmTLIZYR2ojyHIgHy
sJZ7XaU9JKMxcogC8O1xW5eEYc8mAU8lk2T3cHFNsop1CShpLx5ZXYTytdPg
T1uGycQ6v3Ilha+KKIyjSx9q6gjlyHAzoUpXaavJIOyPegoHCR7YDeHYsrtc
SiQpMUfWPYykihG9aSiRWrTBWnK2meE5wrObI61v7K1CWHOvshc82kNhYlB6
g+187OGKQwW5fMijjrRNgCFA1jnh3WNdF+DkZlRzhlxsnrefoTTKG3Ykff3M
Ovn+fwYysu4St7iC3yHAVdlkIFNg5R5tIMN+Ic+GmisfX54/9PpojBor4SDd
WYpsAcBfeJ3KzNRo9e+z4PtY1u5J3Vns70Qi2CSIvMExT3WLRojyEKt4cy2v
5rErsPyWQO2q6eMTVbBPTYdPani1xAmFV1ezkQ1NVgRA78yPQmofGPcLlXqE
p6MVF5xVYguo2WL06/SLJL+EtjU8nqXPxWO+ZAamEkWvDRZwI4JGTaoojSXo
ybO/MCuuS2JcMcHxxaRtV3z+u4WPYqcmquJNQ1F8kfmNg98/4JZqlDANSauj
R0RAefvHZmbw/b/YZwvqKFTTjexr0PIrDbdZGdSpNSkSGSr52g9VShrjUsPf
n/VdHWhXZvV7vdVxWToepOXOdWaa5pIfzrQwJTHTYKtHiCY517SmmPKMloKD
EEYob9ofY2bw9T5nntcCoCV8fdmxnac/1VGvQIfDRu5cb7LMMIkQ/Umg9yE9
uiZ4XFbl/ZkKwOwmYhHZV2aIyde66MtUU/91/pq0QORxKqtSw7hR/kEwGOcC
OXvsMVYC9o5ZvEot7eAfYSepcV5T2dId0FWx5fnZnTUiWqDzfl2v2rg5lYcr
3NoL4k2zVMPCdSUwBQqmWPbY0VNq9tD7emBHasdohwrnJXLJ1BS4S33Yhfu4
XVFry/a9eP+75RnS8wIshM/ia+zVzAXx/cPd/aAjpH/as+h1QH+WPgc497mk
C3oD+9CGDNzlBa++D8Fokmk6m7TqkLVY1pVYvA1C9IK15ey5m+BWxru6N3CO
7SFiQl3YWc+Pa768FE5zIuzBwbYLiAQOP0S4016y83wjTuLOv6Zdi3vPeY6v
QFywIG4hImI0Ia2uciM0pR2ciHHg1UBzVTernIRuiBUtUtzEbmi/ZNPQ3BYN
AaHiMute+iwnJlpaXnsr2Yyg/kKqZXTFN/2bdY93sFKLt8lZGw/QKvnOAn8a
QB6CBOhc3GKvgXj1YTyv7vDQJlYQjh7HnAmWm1+2lSjvldMCE5p/kV6/S/Yj
GtH09P/5aCEkdXmhfO664Ovo09URdf4AIwNO/fKBmVT/osRTIpSYRgrvYAo7
BenqA/aqmHJCk4fcaXMVxXPe/W9GmVmzHeFsqcTxeNZqF69s1o45y8pAybYz
6n5CXI6iJRdLzF9S63o7/B7cYDtLnocLnhqX+WN+Rg8qJKW6RmqdiE4wSaKF
XLMEbHytNeFzwJRJPHqvOf840LEqetq46xs6cRqa4ZS/5VJRNd9VF9d46d8Q
m6L9/HqfwbOH9Xf4OwOadEmTD/tKOjzuwAf0sgauyztLEy67QLOpiyTUm/x4
yYILvNbbHsoPSTeZggaXdzbjAAkr2QbUJ6k1BMocFGGnhJa9oglyNLraQxDk
t11jOysNmUPunISQpjfEEhvYjGgWu9wl4FObIfgTHHYco2w5Iwtks/ZAuf9Z
a3AYejLMyjTnOzcH9VGqwKRhyM3TbaFCdpTjUj+lSq1/yceUcDogS+qOlsrG
IfiSdEaWmiszDy/lYqajlc34F8DKOLw6lsE8yHELprG7PVj5UqUUcHS9m5P2
SAOh7lYGE033bmPFTQE1+NS+XJEcg4QwpMVXa4CCYBHP6x6A8u2c/VkLyF9v
JX1qr9eHNgY0mQEdfmU46KdxCjsSg9u75efpWaVQZeYKB8kqnP5/S0RrJX9y
Shr0UAQpi2kYgP49jRKkK25kauXJEOZVyJqfkav1RCXWyfnR44PFJt5RL+f3
pYZV2/0iPd7klDVrqMWspkotBoN5VFPJEliKcP67oAFSBc70HV2XcYJSFWc6
z8m+vnQfGceYKubzZi4VBO3LN0vNNxOa6ckYTGevJbXWTyoyrYp+AKc8VyeA
WpYOYapWhyLnXshWEK8DbJJoyhtG60X1AL2l2qJdXK4zaytlfTt+LV9mBG34
MwtSr5uOwjtgeo3d/4rhNQc0kK+iIah8qYz0+nDLTuDd+7Zy30bM/h64Rmwp
wUkUEVOMU92sPEskzQ0G6PTugfR/1ALqbxo7fITwAzrebzonEc+Ex4/dZnkT
rBR93X6UvjsHzT1G6lx1IJGDxld0m9U9hENKI8HcGTcBQ/NtxrYWKU3Cd7gw
jGwlQk1AjvMxKLPWCXdVnICiYcwM8KztPyY/nSjjWqUaKFqsxgE4t+zI//VD
KXlanQLFzZhy23IjPaHM1M0oDdjpvMnEVukT9eqqjDf+2jUh7C5323K16vui
IFXfSaV+yT32oxJ4cpDJrkIxeC3oQqAqYrmmSpCybLfkp/M5DpxJlR1A8lws
7TOjUt8RHciJ6bkWUYcF9+lYDyKBj5bz21Rrh/Y58lCcClkp3f+36ZH3iLws
hk49FaDhsqnCI8zDTihEmGPXEqcGxhgL4w6594QPvpE+vP8J+raDfBZRkJ5T
5tT5ixRKgHYpjzUh1cQc5D36BlRe8ChEZUiSM0n/fqVg6TXtsf4CGw0WzPEN
Kwvv9vI8y9ET/k8hE00J90KBylQmsq1zGw6cs1/GRbSU8NT2YZvEKKiGorSQ
396wgZfHQKzv2/HL42l7G3ziOlOcYl9ACMzSa5PP4XCvlNGe4v4tc7uL+ZV1
Ka16YpD5MTzH+Fz6u9G12PzZiLkIHRIq9ee/vBTtZmLjFhMAW/nNzH73pJH3
PTPlE89GxLwGXV33iwell9WUPNEwA7CLk97SIhLwUDSCMHU96SjDLPOM+zBf
r5RCdRiOAqqi7HZvrOZBGiuHd6X+XLAY/gzdLXsLftN1PNB/n9dERvN634Pc
GEyNRNfT9Nv9dVJBjvplGTxk9nQf41tupqVur2r7U8vp6Iq5WyAVKu7q+mfq
+eKv6EFNVb1HEBAZ51hkLZXctjzJ2xgC0t2obiNgDK9NcO2W215NUbfRScx6
aDmFk83Ey1FhM4k8fzPY7AzG4wCxadGOSPr8X6TKLisYiFqzBTPXQz4eoMyE
uXy783FXxXGiRXx4k5VlfEz5XsXYv5aaP6/GauztPxhmz2Ik2szkzJNWGysM
8DwLB2pYiZYzuQ6KQGB6e0y9Rq6k0CeaE2MltjPzR9keRaf0X2QYJwiScZ1a
mKN46n1tDuul3zATQPHCfJwxjeO/fOIaHfAm3JtvvcmJOAMvgRUUNZ8V+Z31
gICEsd16UC2qeWgKj6qB1bgXgIgfdjT5uMZEz+Bia/hZ7azy0CTUDYvC1dSJ
T1vPfuhriqG2EkvR5Mc02bj9ooKh8QLV8mIXbns5Jvj7+Kpam2j3SXpFXwX/
oyuxkoHrM5k92lv+0CnCwJu0mprvvpLeocx0zPXM+VoCdsaGBQhSXFX5CLNH
L0cHtt7W3on9DolQDX2ufk+eybktDq2/owg5SpxbPcXL4YsMbU/KTxgc+dTc
0kznbieTPZ9sRE0NRCI2XN0RXipgHGKcJ5PR2/Ki1xZhhzb4NLpFhth5fIwj
VPS6lXxoYm5xu8T2VzW7SiJW8lJTIUb0e7ccPqGvgtuKx8jmMaRCK28Yismn
S6AfMXn32BxElXKzg/TMg/75SEKc6jI8YgTyG86dAxgXwb48aAF79aI4jo7Y
FgF9Wr49gCik213KiwtKiKqT7K3Zdfe1jrlF+kwxdb09lADiFOpYY/UcHmTF
ZzEMODkf+ymYAYq/wMqP5fucWH0Jwoa53TBO2BN55yZQbKLkoEMrEoutk4/a
uafiwgFTBj71EbeJfU7ZjsWclR1uhgReHR6S6FyPHiGQWnR9VbhTJUVm0B5I
4+Gpfomqbd18tZEuoScS//K2uMPc1Aw0gCMCdHTV6FFoaJtO6NBV7EytWCLY
1AYBVGHyo6AiEHNG9O84dfDExijXKdvJnzUfskFWiwAR0zOVgZDtJQU6GFm/
hTnPVrmRIKIQRc9aGOSuE9Wm5MY6FuXjZT6NjbrOuKOF0QZbIainA9p/ItBD
I0SrWHJmaz8EK5Gr2N1HH+ApWZZk/jNRfJXX3tjotcX89unQIfhQ4vNxr+j4
QZnf8X1R0q3HpDwIZpqAiZgT2JMzJrhPXjpLmEbp9x2XrEuUHhp54LmekcVQ
cBiOZeyPQp/96HnvFKPejvOg4DukHvnbHCL/JJ2GcEgpEeUODly7jnoCjksp
HeF6/zqW7mGQOJ0EWU9xM1Y2VtR4318nt4akUkjva3ZEjhiqZsuzP2wWJ70j
lx2/ghFHRDho37PKRiT0rHXOpLLcItFFQsZMSv1D46Hi4o6/rA2amFv+bfUG
BSgO8Fuy5vCaQZj6pmXeJfgkhYpHDmfn9XhEt2XquNo6cBt3K1BddgnK2+F3
Kt7zkdfJns15/48G+n9EcDaAqXPsjnBHioyvxfx00c+v3AbySkhlOKHQ57IZ
kq06ZxDiskjQJsqwmZQC+qFbPZnPwOAZJD29ojjgamOSaZfhY58pajf//Av/
jlBNLSKq6aYWLlNqUhMjC4Ryhqcmbd82sk7F6e03x21nHMViuJQOm7tXQ2zA
UHwrnHX6D/ch8VSsaWea3EQArNlvRPSCy+QgZUAcN9ka4jh6CgnQ+ZfxdPgQ
wEpkORscNJb8XV0Wcd0QhgZxNwAYAWKNwwzoNKRcIhWnc3O4snFpsyo31j31
krGymdjPcrUk8PRHQLVFL7nZtwilaIyKKNyVp7xcskXllhxThKVZewhLkjMx
4VkPNNOivIk2Q9/F/QlYdGMMamD2hBiI/NhfbLCTC41hTQOxS3khbULhpwt3
i8I4dcdlK4nhiE4jvcI8E5l6na9zhMhjEV0dqYrSC/s40ICJ+9PlsFaLsEMu
e6f/0SGVmrB4b9mi9GN3Nq9eTFVjVJ2nqfis91mc7OpYcgv/ga9FmB9vrb5V
paJ/NxkysCFrvICryGKxGIHD+OTT0BkTeyw7NmP2etZL4jVqb9F15mgSC/Sz
TCHZ4Jy5wn8uhjWquVM+/x1ltwj6DNosMz/Ydc8y3BPlY+D3gdvu9aWlShRu
6x3mte+0Nz4e6RoDtBZaa117AHKIQph3eyMnW0nRuLpI5SUDWBUb1Ahn+Hsd
flSnnpx0o33d7d7SbNsCSmA76DbqwOusHvF4zz8e4FE34HjJ2IPqLuHPztlK
n/d/b0TtdfQxy1OxcnEj0FVPqP4uiDfpifWYJq1hmKnazY+E2/0XNRpYHSYJ
w91G7NdwjdLqMNvOXeNp8T2aQ54W9T02juvu/lhDFAvAOYHGgmub0xITQ2W4
pAsn+vwanPA2vnpV6GTDxyC4reVubWBmE9LXA1hOZGe52JCmgVX+i4LU/d4y
Q0dFA/Q8DcngshCviim56uYVzA7+VdtF8tGqUEeh0fpstGwS/hw7Ce21O0/i
9ASBS8+P90ap0+FbfjEZsnE9KVd+LfESvOEofaaGUjU42NBwxA0yp0viod2e
1oIhXve8n6tKNPF23UHnyl3wut6cjiDs6P3wlabvQPoxdS3IxZEurY3MtP9H
+Ldwn8wN65sZF7H+mHYsHiRwcTg5bb0AHi+Xzf4Y2sp3DQM03Z2dlrnLXT+S
Jmm1jd1LLE8Rp/GneVzdgISIG0FchlzrAfHuwxGKu69rT2xx0xgT+Jocbq7o
vehTIrkwjTgoBjtHROtkrazzDxWQOeAcYMiWeUB1nDvea8iz97mXkEaUZGlb
cYYx50aXze+aDj5GbhaBUouxrw/n8SvZG8iCTm8gfLzLnP4cqUN9ZbF8tVaV
Ghs1BsD39NV2qzmMa5hR/dmEdJVZZFvVfgDSr4dsjjNkPqao9F+7wzfTr7w8
Kf2AfITOGwkUmlaW6oHBrWw40V2AheJoOjMpSMfKeYZKgEt/3wqbtdAHF9JN
NKQ65Y7UM+q9zK4idCJiF1SzL/ybqV2gnB0KPWEUCB7R2mqt8YyPV3084Uth
+A8lRF/vJgvhm3ZTEbtyKKWRRxMEeJgd04MpKbNtZKZPjSkyniI8V/mdOiLK
gHRBv5DEaufLl/FvU5zlVmm4GxkI/JL44yRt4RUP9w4XiOVGPxffEuwmy0m9
pSbOsjYoVC49ofwMKiFxnqhZxX4lU+gX7u/KmrvTHUPqsIhu8tGj9su3wumg
t/c6+TKkwKtevXhgfbE27WBubLAKErCV/xk3SiWvx2GyI/GKAdk/8dwdtEI9
Yx0yjvxsqsN09NhwnVae2WtJ5wy3edlxPvUMsJ4CKOZwATmb7MCJGYi7S3Fr
XUnB4TXXXyFQ8FAJAuY4pbxOKqLytsrCKVcvCSmIyuvyw9UZjzxFvHnN8lTf
gkeB7bcwfXkwcT0rY2CzfiCDsKPWCvbAjO4KUt+5D9VsCstHxtRm+VSfiyFG
TQH4SyCIVBObm1vP2pSJSaMme6Q7Mbjt16CvKPRCNUwBiFZbAxmNzUF+pkLz
fhLihW9x0k2Pg09BXqYiohlX5xA8YPkKXJluDy6hL5T9cogBnv9GKxO5fxJM
BIFvwm1j5haz3Zl1IqHFKjGt0npYSmMwR1ZvMZhy8XqOIx4GA+8W6RrZ09kV
UrA0O2FRAVg5AkYDAlaje8GIpa5uXGq7i5fSefHylX6m3+p2fBgqRf+C/mGS
yvxE6WVzbQ7n6MMdue6xW4FU3QiJE7x/ojZks6fobq1cKH3gZLkNC4TAy+L8
NzQimtSOwvQVzC/sByBFAI2jfofR322OdL85iL9GUbOCiJ4G5YMf6HI7ZMn1
Ezy0z9N6IZjbY2IvshpzFMR58VnvrEk2svc7bpAEiRtrnREexUrm/1w8tmnG
W18yrRpZY/1swckZ9dVYcASj2Z2vVXdzETrrxZ0XuXGRQnINitMFki5I1oXl
l2jaSuFhzsTiRi7QV+QVpyWSNsRizDOT5kewvSDP/6SFYcUxLw7414qI0NwO
4z2mfwnTmIip0dC1imDafVuKPwl78dyn2xRXXKGqMBct6w2OwdQOXN2da6Wv
Csn+XmmuKgHiLusByyCR1IDqewm+KAeRKrLCJFXhBzAxmf7DEWpbXWsttfl+
5MN/+SvgGZIIGd+61DrEXZNpalCHe+vdXUnvXHd+KUzY3YTYSJj1uBBn1B53
ttx9VsyhrUmFcM3jCVNs/zVkB+WSPDfhPKpMFuGH9LT6QR+rjgpKADl9L6zb
LWDKiFxWSJBDGwLlykG4f+lGz8J1gCAr1MN1XozzmrCaV9kYvH9r5rHCMLMw
K2u4QZUdK/FKuoeUny930vNIQly6qeh4jZuYcStgAqlP+dp1FWH6jYtQQ1Ng
nAI53yqnd3izTKGNfj0PdwdIa3KLP+Wb1UA8LSWTJBmSgouTwtM6zgFoWcDN
RB+YTV3Q4haTR+p60enYHAnOD9G7ZXY1v+mS7PIMrYiJstIm/KFdjREbl9M0
8FUIhs/+8Nt+K1vOlISq2jZVQclWmEfs/IWqgAVDc7kCxlpyBBOHawUNwJiU
ejhEPhh7O8lyRilPZvxiIpMO44m1l+bOBj22MYn1asSpP45VtzZsd5lBkUef
SRLRUivb/tQ6teUpBR2Ia8wFUoKWdSjDYatit1sbnPdCchu2dFlFOThTS2uE
3XoiAB01t4U3OA7DLCYmZEtfCJgE7jaGIPy8wDoXzp17gutYvIApOYtEq3aQ
Ne8nXnT2TeFkhY5D5k+KWJOn9F5ZjJ1mp5rFfjI2OOE/pPqOUGquX7/8oaJy
cvzWqvTC3DaEF9sEOSnC3pVEPC4nAQm6toqgSOrVM388KZaDOyITgKmgkWTD
V7I4TcgkCl6wxPM9kDekSPsfSMAs1DRhQMF7M9K2mwh0szyTrwlj2bomwrnR
NEvf2WW+zi5Sy7pJh+4IgV5p/LLXdR4Ai/zk1yCdPyNa6kmz1rXTnLsaZK2N
tPKbkqn28AVLkQZ14yQ/zodql8WWYl2IH5vP6iLT08H/zzvZv+sU8xtIj0Vu
2iMko7R2njleXFXs45SgTpVRKJtFNbPHuyhKesXyKFGK1yk1SmxGiFlU6fTn
HKywo5KQTuuMWluW4U8YE6LmKkWL++yEQGoFe8COliSSRm6LwymDH/z7ilJx
GIafbbbAxOEMzbAXQwgd/QeBhMdKh74GmymBolR2BY6ZeLwFZCiYdbcq2MsX
gI+HV63ivKT7YAx+ywrkvqBl1T5U5vGSo8RcVMGB/sgx6ZTs54TnSeb+gY6a
PyigWKV3tlHDAJQr5URFmAOyKaKsLPFPU3dnsoPvKG8grfHb+3jT2EkikdhO
7QLVt6GH1tOy8rxG4b7jD3K/Zkj0dsCp8gXEZ1wohYnlyKrwJ66Pemp5GY0f
nHDkZRi7y3R/c5HL3tJRxXvCSg0Ulff47eTmFdGEWM2qkkbD9OLvcALjJsLp
YQiS5qf4FsZyv1fO6h3x43JiRmGHA0yXqz4zruGfvHC/BKLFBicpi6axlB9q
uXZpmJYVzLQqsqi0NJ7HomOdlhsqLcexEOWkm+aDjPpH+bcZyFwY81vOeLjf
Jsni6cgGiBwBtnXxRGUszEFHGL+6Oq3lyLs6NAMhZrrxSSpqjKokxJ/ecFMp
g/Ei0n8BqI0sd/Bwd4We61sYjCZ0TvIrkuqMdEhPjKV5Gp1qoSCwyuBC70//
lm2j5VTYeXpII7hX+19qDF4jPmKPa8cfbe7YCIx32OauDUHIADdgOwR1EPSZ
NFJg3YNian/IcnUt3TAL4RoDLi0UdWI+RxmW99v37sYCGomDSdtaE5tMtdsq
Cdt468SS0dP7AM+gaf4RUAsTVnV0bbQtDskKDhxk2X+V1gNpK7aatDafgnJH
g8wYengDdGZzhOaNZnPkbvKt120vvWmm5hhiQTL7RF/7SWfEReFOPqJKSjwy
qY6C80UxYlPKCfb3GRebM/Am1PJXYnh9mBnG0vc826iOA7kcnBLaQOvT/P94
g7XkxpEmFPBun1agdX84HL9t7ZS/E2hUFUXS6hm5DfgmjrfkztnOFOCE94ME
oNKI77myiPyggcxik/bmy1NtzPSVEvQICrYXdifBuqssVwHIuLE3lhkGEa1n
1E/hN1ZgZD0m6SSpxVqL+kwngcBHGW3zU109qMKS4+ibzZHWfH4fAueAYxLi
lALv3LWy/mneEzrsirsaVK0/c9RmX/CDp8++LJxYLAZXZU9fCUqNSCX2Nxsk
ghx9mnSvn6TCGMbgllxyige+Xn9AZBjNnIhJ91BXjbcYsl+wAV2SNiCitJm3
ntOnIN5vdk/5M12iZmNgCZgudAFgbyBlHq5FbnURo0tUx1Ct0MLVZXakymwp
m0cxFJlQ4IOUVX8Vl9+1FDu45it4W5lst+CSzsWp1oZDv06QyrqZr42O/CNS
2l1kK2K4uEBeu43C9ZTG0DM8OIRGWJySW9149/HFeH9Ijr7+YAOtxOLP08aZ
8D1JMRWRGqYQQ00Jia/kH5iPCqyrJsqvPK4IQlHnpGCDNxTsAjPX24bJxnAK
vIo4XMjU4UxbnBnMcK5yEFBLwvhGOseF6/nYhFztluQZSy4kbEzU61XiN5OM
HLthlr2sH06ZssR30KwCj22ogBP8M4nP78uJYdKWBlcjRg3dpCtcjj3mH2HU
816sqaZsEXvQut8Wc6S4fl3nVAsOnNVvhWkvgGieNRRebtLmPQ5MhSc7lkpm
tNzyDZaCSxta0ErwHK7eOooh9xWRyUTAF8DE42adVzP/fqOEHxn8qXPgNvGm
yx4gylGMzDRJ6EV7iDRr+wly3Saj8PvxP6LWmEvlFGZgUHA7i1zeopv3kcY3
85FdmAaTeiaQ2mBCsKiB/1c/OloBg7axknbpvYOi+USuaaAJQborgIbGEZmG
Zapvk3wV1tPb8xDFGrO/ZsxP5bvnmFGo01reYalYuii09dvtEZ+Thb+U8pzh
p3GRD/tXhTgB7qAbpp1g49sWR6Entr2BJw6w8j/3tJpXaUBVfmMnkMnf7mdB
ld16rLFzZYYUJdUQ+AEbZd+BAaVEEt+8YBm0E66zRZ2zBZ27LlL69rv/5elx
JBbtTg74o8Y6yf8kUCf7AO3O9aiztWznodblJvl5KVUs9F8rehwnNp3RZsx5
638YKXeET4LjBwo0IR3zJ8S7DL4D7+MgRaXz1vXa/1W/4HWLN8rw17aP8UPD
Q2VttS7+to8i/kEUQCiWchcRLFqIOWPM5lcFYZY2HO/6qHVnaz8wxSYDuzXm
n6RPr4WqEZM+A460iuymLwPffqpioRl9tEoThmntkupAHS/kum3qt23ZeyuB
0KWTHzRwgLm5RlWMGOReTue9mo1B1JC9VmpRbJ+sQ6OlI+LdNlvW9Ku6UOAH
sclldODkajObljUIkgsOvu2qUXe3Zax+JzH/Ib4GxOQe4R1H7Lgam93H7UK5
8+wmXPGCdzWbbU+hQgY39sbAau1wyTOQ03vVkByEKN/0P6qQNLFOtSRjolnw
wTmjam6RsKi++NvBeJ94uTqwDAJVYtPW+EmHMt9u3WRKOxQ9ie7llek/vEU3
DcRFhMkBBE2zxRoJTOX+8d7d+U42y68UdcrscwKZK1EMtErKh/ptN3AKDNOj
ZQu9Q2s3bdy3+dyPChjebarWMwtenLy2kOV5HdzGJTotpIwBDYlwqjHPPpQf
BTqdIFBg439uCYEAVNeEO2AJhZjMutuso1gkdAQ0QJrd4d3Nsu3ws5BYy2R9
CdWYnlvVSJ8Se2VAvjqIG+elUK7Fko+ShZUjsmrhKAyxmszqdxZzv7Nx7KIG
XKEEr/B0LElP2iZ/HYzSTU2Q9GOBHRiIDKVUWAcrtm3IItQPTQYZana1l0Yc
Wn+qAT3xg1qd6pMkdvu+Wu+VUyzY2U9F58ALL8S0Jw0Hd4sObT7v7yBFIgkf
81QWzcFOgzqqXI6N0x5ZU6inyia8O+biC5DDnW9WoXoA1zfQDsjGeIRekpji
pHdWdALWO2RXiEcB+UkqSdUfh/IZJpIN1Rrp58OA29HyL+LuBbLUct9S2+w4
uzs+WWRU/jFEy753698xREMfQGFDjThJCRQOqcC6WINHLLKRS80tkIiYeKTv
r2xFv5RlPujbuTJDMf9EUUDgYQKRNJC2Z1kCKCRF2tCwOiOwYBlCEeSkMuKa
uJe3xGa0gx9WWCQW98rfSn1X6PubeD50diAT3dKSfk0WQMAaojlHKcAUkBhC
MYMXodpoYoIPE8a+c+2SymHV7FQbWf1JUF9tpb6M185pIRQQAGU8HeS5ZUnN
SUgDTkrNvSS2seWtKdENhLGyN2DzmQA70oqdGYGDQ4++5N/UDc48th3jVWYa
VWuauG0VOG9CZw5fUdoqPcDEF36wL08SniiF9WOQcvesqGBBE2zUMrXdWZWo
F3MDPu7yXgMUTdTfFTAj8ocXpyCSbnilEthMEI7/i7CUbQ4jNbW1DfgEfhPJ
hoOkMTizplxbpZoeKxcUY0WpGhfxbXdJLXW4sSSS4XY0dkXXgGZyatPDz401
h0jF1YiPM4k9PfJfkesjyFSkK/UuygDllMVoYewQ9X2yPdligQb4zmYHcn3i
0rQToEX+USraPopdS5ZvSlrnG3Zggma+FECWLU5FBm8HrxsCOwOK1ec4epWZ
FcGDi9vgUggD7TmxfViGcAngDsjQriajk6pAJmdDYfZSIZ8ZzbzIISfLlV3w
5Tt8pvFdh8V6zCgNCukeqEjvYIoqj+5BzUf4toovpvpfYUVYAyNWyJdCR2cA
4eGUs6+ABCXlqn1ec3T0MAqmPc5jq3abNid30GkMvvc37eCjKop9oCu5HWFk
BKfIrNuE9XvDbJVLj89U9hZMV21yf9BbRrjgx9NlI7fHrFJljEZi2swcAxV8
UDdR3xf1CwkIMV+OUdBsDYaElMBDz86BUoToYxdv6hgnPJ8PyAC/rgkV3XPk
P7U58ey7IpGmk3TK1Mpx8KIK5mqL9xgvFCDoHLj3AThn1zftWUtzpEC59x/r
93srmXyFmw1yY5jhnx2g+hT2tuzQBQb5VzkXwMaRPFukXw/iwpTwl7FuY2aw
JwGB6KbqxU1Qi9eSd5PaCvU3NObXnW1ikTvePrFtlfdeQkj1m8+ekD1dOqSZ
vZlXngb1QigyFFClbmTT65gtus4EmijOCK9w1U/AUIcES6IngkDeGJ1vzTw6
WJgUeEMzxDAKycGRQozfWB1M9qnqP1Yw3/wWUK/57231/ThUOqhAhpYKaAWr
ATD4d5mg4O+rAHctcCdS2fbG0cVEN68a7cz/qp4/A77PzM+tEZRQtxVBrPPK
JN/ia9+h+0EwzHbdXORTmHxjO0JC2UJpt22HuirdQUj3ZfN+tv6gbmfJFRoX
YlV6B9yP+Mn90crB75R8PUuOTpJ6P6/jO7hmRi0IVnEsZZnxSY3Q/o1lzQGc
GHp09SMQ8l4xSVLRP0cw3GkDpJbJlpNP2U5iLL7alHyB2UdBnHIsuHJQCbkB
muiVswuXR+NAFuJcISvVy9PZLm4udNHszE5/hOfQGGtFP2KspyHc3kGB/z6y
w+0fg1HgiUw84ra8XVae2aP4CxdMwoczq69fROQCCdjOoxPvZstMd6Rg98VE
Ok4/nwLkQx8KrWDPSP8Vwe+7EukRWiyGsTPJJqs/uTfGJtGvarlxGi193ZBt
H4yalY+aL9SODusUwjpEdZxLGrld0y7FbsMKp4UEy/G5kNpN1NsaY17n5Pdi
jNzxelJtSRAShoYoMS7/RBhNVUxVpc56WJL91FiQuyULqKpQP0whnIq90xKm
ryS5gZlKPpsdDENJnirbyf9FOTsB3VQAUfcNIxd60GhgmA7/ahSDzsuFJLL1
Jmtbt+8HNSAhdptfs3zVfzBuIS10IeeVlU+/WGm4+cO5VxQNPp3Y8NrxKME/
DVK6KzOyZ2eogsGDWaOAnzW+MJZaOK7BX6W1CTNQVSpb4TWhTXCvNmns7f/I
hYVFsAz3KG8Mm6XVvr4PH8CFhXMepPvccZ4MhZfc04qhAWq+QpqjkL+Z+8mE
tcvWoRZYPMTwlQDX3D04IrjzXXcGxZFTy1J+6Aw7mBpAVLLlOOuaCiLFOuRq
7WATkZW7RLZ+k8s3zFa6wyuCqgnDWaCRRKtd0mQZPGIj9W6kAMEAX8p/6Bqt
HvhcVprYcCnI0zKr7TLurRNUCg8TcjQquY1hkPwM9Pwo6fRR/4D9FNkJUE8Q
4wOx0panqlkRpaCOfk31CiXBnTXASBnxAEMtyAyyV1YXpkX1Q00+F2LnJcXB
sONEi7fQeHKYM7CTQat2C2ghSxVj50QchfMJ5LsTEYWeVOu9YsZu/T0VF8zr
7QPBC38dqP9SBwtPld4EKgHXveSpsBiH+b2J2Zxze2U3NaVO7Ypgwcv/ofYf
3lfeYkXXDXIX70GqPxPxPfhxrX3jDQHzY8VdvKYLn3V1mVbNIUrlf0XJjqic
AWL04qZrzJIH4Rpu+7kmHLQnKjrHKI4ycfxqyz9WPE0xHnuGc+QTasvJ2MfC
68ZYkL6Udk6CHX8TazJ2n16Htg1wC0XGO1mGXHw+hUlrjXywip6pevqCecMQ
ADbXdwhR/iGv6Q23+yp9R77H7AAz8seXQx4wfuB4XDTIVYPXYe/4bquVrjnC
Plh9xB1AIRBWQmezYsWuodHrRsD9RZXmL/qfugbVMPCido01zF6DyMRih0tZ
q1/sjE6jZQkKGDP3DgyCJHW0OzTEKu3Co8hptpuMkwF/npaDvewE1vpehbER
SB+gXcehuXdvGMjNtkoKG2Gw0ml7oC7wSGQoeHdJ4IuaCYVMAsEhmsY4OjSP
vemTAdWn972R+zDyxjYR1PZbuqxEJTQ2imrnHG7vMWspp/hISzubEplCdkk2
4QX2TbvP1J0XlJmOf+qF0h0LfnsapPpaZBw3CuOUSw4xlSc3xpTtXQpBc9hI
tlRsrC8/07fK4sbIgGQXl/zIZkp5XJc0iQXdngv3S7ebpZTm5k3K05+fxmWB
ojd0eQncV85AHnMIhMvZCgyrzXAgKmYYTI3ynMppUPll6ksSA6Mg+hChgFRF
c3HThxVrfiiHrp8M0rxaWxH1g/Q8jfVJ96z6j+DCRd3fYsFhhPqUBjOler6J
Q1D/zGTIcCCgokaekR/eA8qXsieUWT5qtByuG+bteUOs+sWS1PssWY+MC8ov
K0jnYuZanZ8MqvWyQesKTJ7atAul6qX/wVX9kbd5t6VvrqPSkPe35T3NjhuK
8Q8YnBLDrrRVSMYGxEzAUztzN1YxD2WbF0hUnZWw3grIWw33TghmLRCnCX/x
1dvEp/gpmn7prLHHRxtMM6vO3aT/qxNgWFluDB7BP384hp3rI6qtx1L7lQ7A
H5C3B9L3fThDmPSMiJR0WZwY6YIlDVSr62YiaX+VM5dPgjqsDNEEDgA04YCz
VlUcmKbRMnq9JlJvJqBuJECvhdFU8bbX/Iy2J5W336wBfxkK/hJVadKkMQ+t
0w9fw9Sq5vZJxDXGb/AAPjGtBdZGUE1JlYpCbJApZ8dzYufzEDmVmMF5Tdb9
epqscyVeBoOQsjpMtQNAcAYFXAMiRQKL0nbR7hH11VVq7+n5nE34akwh2H9R
S6T3pMCtS6YLCd29PVZpHThFfMXFUBsrTr6RhUxW58hjpnLeG+9Mj7ViVSBV
lZrYqcqNvorjmuiKCnRZfehzXgZKYKdrzc6fK+AVxrejddWSd4da4lVf884o
UdfeD9zIYwuqoFYwuTE9geSHZJBfrn4XPjxiAHbpe4p8qf0koVx3Mo7V+DN7
p0aLwVbRO4HbmIJETobTnJsliDuY9vLQk+LuaeCh1seuYpW3SrEeMd0A9oKJ
8t7r5iX4DYPfvRugqu1pfjcFkfWBtDIUfrWZXfFp8OFbS8wrFRovnEmNoFur
5tDz7tjLM7R9gfGdJCbri6sHYwrlJ1H/vegjRaBqw2mDvmtCHGrZMrbowV0R
boRWdZ9NAFW4a/ttwO+1a9rH7+EXlbTZr5PWGNc0+b55MxvLoCfUH3267/J9
5if4zcAgb9EzLXttwlrgZGWvSOt1XK5NsCpIjI47kGIzDNo2j8euBNfYk6Q2
PxZ+vCNrdnOAeUnHRFrPE6gcPpQND4s2EbTjP51qRngbnSKTyrzxZ19Y9YgJ
CWTmoi+rhA8JkDTWdmReUEd2wCQT7scLIFLdfL2PfBx6gZ86Ec91+n9Zr4nb
CPVXA2lGrRta4MfZykq3tuioHR9lddnPh9n40uSFQVuPt038J0I5mrcSq55k
K4l9evLxtEIK0kJUp0I824oohJcboeXD9ErJZFXJrdZ7fAxTWw8zVsMH0XrF
8VqMKiI16tVw6M/woHpRjvS5rARaNmMcD+ocf8OwiNXG1OUnQduqDdtXgmyK
DzJqyWAUs88oQSELYAxM6YZgFMPcK79tmGv+PL8EZBVGZb6B+uehWF9RNFgA
7esUN1FmmWGmU8jgP5J62Ujmr/V+uPrtOsG6uWw4aNsWpLgiGKdND2GQqozl
KhhON4W74yfhbTLQfhtSExGZk/A14S9uUgJwu8ge4ctLoKe8RX9kymkxIrSU
1QVzAhKAYA2Xw79AdjDSUbymzCAMiZ6xSXO8FmW7JvCto6NWyn14HoOslYfI
WdrqkQf7uJHYd6LUbRy9yddEU5NitA85n7vBwqDDi16mg4Nx0fpemZsg4vSQ
76PtMXcnxWzMczOg2t9L3uXc3cWW7BNYEvFsCaShNl/fIYbKy1DvyJwM7xl+
mMdTIcaBANSO9NAM6Chaui15sHOizyR7f77k6urMyDnlZKl2jW+zL9sBJTOG
r3tFv0LHetUbLl7r0NpklxiKaSAr9ZvrirHErx9brWjt7KfzuXCT/V0hFQ1N
KiC8YDvBOKrQGOdJfpV/uOfkV3gvntRnzAcyqR4Crx9NWk/aeKMe0mNbEmpj
Q9qSb20MnzxZ1g2IM4aZVibfVDNEkVFBZEg3cGSPM5TP9L9BG+x+GhJpYjpe
ZT21J3mHHBhgLkcpHSH6AE5OHxuMPfmUH+yxlrXtTrHvXhvkHrACquBlXBeZ
vfSxX3Qj9SgYemm3h1/6N6HrWpK4P/ySBLypQqM1FcsgaqzU4NVkgAurN8KK
wxrimGXkpcVLGq59apThAt0syzr+0Vylm5+eR13+JBBjk3jHWRAq5yY6spmN
LNxFlKC6/bXHx8wmxEYgmhORgfMeZQLcMB7pa/W+sqcMpUAUUFf4dEvboXpy
Bnyh5wpPTQrQM1PXUEkWWW6tLEtf9wHGZfLIsVd4T2swcWAZjpqaSNqw2dbc
XNktPHcy2mjG2Ipy+Q7nVvy58BWIVIs95s2bcTOfBlWU6S5in72DMouht9Mf
23+aoQBED6/ZZIr9amOu/QF2QYze7QvNWCOd3FF/eitmscst63wel9dslYD1
DOqsHOkHdaYFhPgkPK/ZH17uZb6tj48GS7R7xTEsSXDFFiUrPu6Z36oK0kEV
639tKKPwo/JnBQkTHu4tsDsb0uoYO4u/f1nnydhRMnzI6tkuT4BovuOTnzMO
wlTvZIXwOiebUrMI19r9teqpnLmbP/WqPjcEQLAAcR2oUWgBl5HaPgzj2jNa
Y3J9pBPj8FcwYMLxsg4+0z+yb90YcnKBbZyXc/mt1Jz9/4Ry/KBXBzKlafwq
wWwg4MCB+eKsWdp5dHPYEKdpv7LNZ+y9JsuViCI/olwWkPbRlelYDseU4g5l
RPUef42tFPFxHZewuhdIb5j+AQOjo12r2aVSf3l9KUFfZCEZ7GCkODMWwaiE
nT8F7xRR+0Ec0z13bouh4PITwTkR0mamV0mg++B0Mm2mKhF2MxksRB74g4Mz
/kXOxZKqYYdi0TRHyx4kHR6tcYC3hSeWReGwdzY8UueegUBwmCtJ8Z61Pw+0
FpQp0fbKRZOHWlyyr672ltUhbebVHWy/FovtDgGLpYYaY6vL3GhMgQkaQuGG
boIR6v6J0lHJwZQxokzOb2+0q6aY1vzYNlZLjuC84qEU7LHaV6B11y2Xflnu
t7Dek31bFsE7Fuo1bqIQsRjZVXhP2SNtyoM82C/53T3BLKll+zusGQThmUBN
fyvuVYNk52w4Dm771HwW6jW8niBfsH5CWTpHHL0D4+rZJJKWOv7/ODH984W/
2a0ij2zCC8uq0BLdwyrsvmmRLgsogzZMxeIZBB60aLmOmroDkrSD/hOpLS0a
qMrfRwTb3vn/yuhBtorZdqF4ycfv85lUoif5nCvQkSbiOMTeiAVYo9TToRRo
h6U44elOmsswpouZv8dUKKVt8cBTXZg+7wH6s+Fyv0tA3GKInElP26Hojl/F
aaDggYYTxj2mySOBrC81JFw6vc1m8zMZ8wjrd0rpMzFuEmUnKt3kQ85DKfHU
E47h7AXB3PtpnnZjjiIjS5ytN2N9+FXNluY5nVARihc3EBFj/8JVDl0qaCi9
WzsTIJVkSshvbj4PFdxZXUTz60J/ccTKTQ4XGV1Nw2Q0bCsJdSgIrzBnleyR
hPNOEXaM/TT0piRtsX29Wa55CqHzjdSepm/fvn3Bfah+Rpa91rRugfwTy58M
r/Z9Zme3XrQ2v7ygK3LlDhfqvuAEau6n8cVpJmkyCqyoMW/QbR4l3KFjWAIk
3EebWMISqjbTifdUGnEGhDJPmsZp0llYhPvLTkVZBefNm57ZMBEYCcYrXwDE
EhBIrC7hhnxXMQjP2jZXWYtEiMMWvof0zuFbjUzjYdWTgP8ADw2k/LKdF5CL
dWfnMbhvV99oOIMOakTvwqdlmzneL5iQP4AxEeRoKhTjfms8W6FJEDb/8iSf
TPXYcGJ7y0hisWb+TqDtF+YpBQhZ9C+ceM1Be1Igi699DqhPGeZS6w77Ma6J
WPhrvc3p8d+4s20Vfm+JeA/wKMddEtrjEKzVwOkwpSLP3CQ2k1kyEC9oNPAZ
+Mqoz5tO01lYg3ZWGNRqR6p2962loRqC3gtWZykdE9Kf7u9w64UmlEcQVM6W
xUSa8HgDYloQqX70moe8oMBTgRao8tlDlPEW59hmwQbS6dVDEmssgOrDxgdm
fIP1pU6FX1FLE6MBuceWlUsXoJm6JqtocENThl0vjnChX0Iq4ghz68tWGE4p
lz0nr7gXKfPpPSYEmhK0elpgrKDyDpY0j5gzcXDZouAYLlpBL6+T1Mw3pa+G
GIEhYtIT5bEuq6s0+ezXIsn6D6BnzjjYNLuNb85YMrCFyuglkp8FGc7jkvFU
SRd2krd1iGI8r3D+vlA7yDpH8wuGTBD4ctz1TA7UQ32jkUBcoetFAlKs6PHX
c1HZXofgjXjVZet5H5YYpGGf4YSTJZUW1Lyo4WU1aInCeZI+Nv7JHR+FkoDx
5gX61DGq8n/C8CNzspwqvw4Jo7v+x8xV4i77AJgcjYIW2Aji2WJxvYEwEPF6
JEK9b+wYDrVQCxyNRgB4Yq4Ntko8Ds7CfEgLenj7eoB2LUosTsnEW2ySfNEr
id3uC0GuaI56h+1Ba93wbcv7IrCRCeV58yAv1X/MGYNaLdHtrNymhDspBHIl
ZbSbA688wFI4vjU3FQO33Mruo37yYwUbzSPJkb5fVFARo8vOYNYBUYyO+ido
J9m9PEpzP10BR7Vq2fzuOxr4Ctxo6YGInx2OIa40tiknLV8IramUwHEOYM2Q
HFE6XXRKqxt5Vzu51uR0k2PizhgMoaFOROOZN8669Xa04smh8apHwUo7nGms
BdL550A6C0Sk+jnflrYWhuodbHS2tzpBIT+UjVIls/1FFqtuL0kykdPF93WQ
rbrCsCCR5LUxHF2QxZjcb1lHxkByzYZLL4i1zM5x0LhHOYeqwOJ4oCMrnS0e
Z9iFgq28G03W+/OB/cN0zCDctrBjkz/auadiNLm302xd1jZ1aXvv/mjer1XP
qp7xt7mdteBC+NPw9ZJ/W37y7XE/XXRAuxxDGXcdUYzdOU5qrkrKs+rhrio7
XgsBtvTYtqHrC6Abj4S1HwX0MZnk6vI/PzLl9Hw0eHpXYNmmNxSTOBTVP+/5
bLJOdSrMmeHfxKr+SmJvsRr4d2xyRml3jPt4m8SOYvwOsRwwfB3aoIbtoUNx
2awEyuwJ4gG9jFo3xetaXZekp1gnb3BkKH0AutO4izCYoZFxjjnn4JYOFsC9
xtpGCrJWeMRXUkllmYw01c1h1d39YmRbCi4KDp/TbIN3yAHWJU6N6E15e3bH
D/z2+E/CbWb1+/mXLxjoFj3MYaIvLsUIrzAmsdJsISES1MzOSjgjXVhpvtXM
jpabfcdFUAlnmIn8o46F4WGCtHGhLGHC3o/Cj30OxZj2EW6Kpya1kDg6HYz6
n0UcjMiP+/iqB1PDTXOytHaFOt5HgOJLTFBCNPC6StDLJ4nvuN2wJWIyFY0T
S+YQNIa+7vy0B5bi4RWNR+Ny4AJhdotJBEgQxiigQjXBZMIafH/CrMwAiYtm
1XosZeygG5b+l/RS6+aXvw3PSRIYXSprBSEEudAeQSRlIomShxPl8uZ4+4rz
L3ucaIGYlW1TpSTvHOiCd6d4pUBZ2C94biB+cgog4wj5/K1RsSU8VKrTrg1L
px9QkelAgCfXYDOkXZlJGia1nCjHYoZIyQxsXj4uB4vQBy19dCDY0FcgAlvT
DHm+UInli7x5sZeu9rUrrNrb5CfEzd1B8y1kvwmV1LM5p/zae4hBk1XDMh1M
1rRENWcX5G7sZRNgSxT/dJ3K7wyIxDaphhtjzlmhT0JKH/+0eFIluXkn6GOE
sPpHl/WHLbo8hxh6QPbCXcXSPiBBmWouX5TBCVfn3caYcjO6gEiUL5ZGygD4
bVxV4pARnbehqAsP4oipdSRqY9jiqr2nTUiEDNN2tAZdtOmR30vjfF1jbq2C
jm6Bk+yyIQkr9AStrJ7LYqV0Iscy3bsupER/WdAN2mYeZElAXFlNlMNoB2JZ
z7OGDkLZF44YXPkGKpLKj0kd00w7ICPvnpv5xKreFEyTl4HxVtyRsmoS8wT8
NnXlbGP2HIAMUSIJfvag4qk9tvRvkdLHHHMYR7FHQod3pyGcY2bk8cCETskU
5OeNquMY9yLbdWkCAoKyKSMb8mOTZRblT1FeqIBYbA43+dPhJUbQQr+Ci/oM
SR9w6fj2CsFvHeISVkMgWAI+RRNwibmg/yRbmEwTzl5yda++RUGTGBxu/sBH
9OHb7TI9blVcZqUpCIP8+MXid7eXKpw94+jCR0X+RPoLkCVE92xyFMfoV4lY
suu7IiiTXLeCiBnCkzn9iL6Plx5vuzYloqjBc0OxXwOVlxOaDNz1OMO05Opu
jmx+5oakAc56UQVwKG11YBN0JK6jJC3PbXhX9GuoVMVFk9yo0oHE4f7H22V1
0dXt6xZMWGK2C2DByyABhP8S7Cu7LohBUNd0S4GDGoDgBEvQUgpwAx7n0mOn
AMx8nVCgS/K7R72YTqv/wXIlfm0pY6BpTDn19+0EEsNUcNEmIwqaPmHv7hXo
nAzd2qXcvU79bozE8bdyF5NyjXPAHg0ExHw5utOIxBVAeYIsh2CnvbtBo1gt
KJDXZQoiariQsvALllxD6l2mRo1sOmLVa1V4t0QSPbvs1qxpe3UNeVSZkV4W
tpKvWDE5Fzkk59XnsllTSTNmdeaz87a6i7l/irsS5atSoMzV6xO2vh/hETCe
27Sg8CL6Uqxh/67MXoscUWEGjHCTCV5rUP+PnEKarHeCBrerJDaUbIFuRxkL
ohvSRcg7b2J84OUFXmJjXnUDdXex4dgICdfLp/5GagioVMd4bkKpAvpZtqJn
JT/SCBJCySpPAAWpowiJg8rWIIdVfMrQQ4dcgZoQOJRDYTKKW7Axoxd4AeZf
DLxBH9KYftGnq7TFGewty+45RSIYaoo2hmo6aTNbVhzVzrD5A6cBXHk5ud4a
BdcdxDDP7RlM4cl17AW/T4VWTQoBVN8jeapR2bZCZAzXfWceiVw95z9ZoprB
2/dB9yQQPDzYrWtRkhnoZC4KijDSsUa7eKeQmWZa7/SX2Nf1MJVbVkRJj4bJ
MVqKN4+sw1FemuTqXZiK//uCsMEdQKer8vtYZRd50yxWjra0pr7DHp/1ShTH
sIR9KDEOgPI/D71nakOtsxzpLkbPbzc/5xIauSbf/nBATuhl7w4TzD0hdbQi
3hCzGasAg3xqwe3e95HySteOtRBEhyiJSOXA8uOMUaneOddcuSHY2kIp8Xe3
gLDVq8nT5lkoC85hhSyOn1VJKqrUToO/6yuJdOxBXCDpAjb69+dBVx4WQLR0
KCbtG6oZfvskfKaYXminbFnNtEW5eK9g6WxO+a92toVwm/Kj7HhbPGAumT5J
fQTa1gnIRsbws1Y5n0TgPEJncJdNU4Giqa/Z/EawWCUJLltDRoz/dPo6hGsZ
ARWdmqjW2JeW+K+y39ggipuSNepr3wrtZTYPJ/Ii7SJT21fzUBUk6UWWIwOy
OLRVK9MNa1r7ZIBPqf5mCQ8SB85DqfkOmZsApxYJDDnTWXuC1EbQ21TSMR2O
wymci4WB/7migh2D2GvdUGa9RrCWW5Xy4OqPxUn+tfpWHSMD1IXTFg0ybZzi
E/mW9CLSRNofoW9pqMQMWVEk4N576HcgEdMpxbKfLXZDiLuQFNU/MmR/uFKB
bV14LPyoYbC1ynq6dEjEjG/YL3lCHrxUGhgrjJpo8JPJgvzRr/QR2oLRHu+S
A9asfA/ocv9X/3nCtzMxuG+saQ0do1OL5fNeKqCqrHcSCdOriQc3QUTg1Wml
7iQPtW+uYLG2JFdYIGgveaF7RYT/QCY4duuxhPvkJ8sj8ao2DtZrnHPAgVmz
rtBR/wqbFQYXNeCL68OY1AAUHU85rjWUfXLbFaWAbcZlnhN2uJYKflZ1/ff9
k2oAxXj2ymKilMDOQktMLIlHK9tuxW3I36WF1/yur29TcGtGY8+kOY1/zSHl
Lo0cPoLR9cUCnYXNEhOPdiz56j2KUBWre6lqXvxJKa2horfB8Kw3rTrdWaK1
VfJR+xA9qxARlDMK09QoYduyYGEsaiHlRC6ZwXh8+bAGCCPZnoNy6sf+qaTG
FRTfRNMHQm31Gz4G1aWdG0l1YINOvWcvuykMF4M65caCYANe4j8DGpD3UpGP
ZtbixahTAI7mAHSQhBRMS7DcYwPmvcaVr12BIWXpMnHvQ6iXPyThu8Pu8C42
Ds5IZmXCho/PEP5wh7sN/4zZxo36i9vAq5Frl3/E5TSbYbaPJtWwR886k5Ni
L6Nf2/b00QsZPef/UJ9cR2RKYa5VYrwkFHO01zuXb/HOH1XfsUblTASYbrvg
shkGzHaTcJywQZkMMbbOS6n2r5CUpxOkdJbS5aVnvIXz1HLQTS5Czco/7YLD
VCn3T5eXQNcemCu/+uSTZrPUcJjmKoJONNOiAgsvkiDHBgulMF3sp75LeDtf
qUDiEYVDae3WUxsHliOFTlc3vK+CJtEqf++hCD2kir2NzpnMHHg7Jj/H4JAQ
JeZQsz8sKWOrVzoc9KvsGok1cD6lCNrJl67Y4mmIXsuzlfrKJCQ1jwVVrsxd
GTydasLNUL0372JCLxmVhB5rxlnZh6J42Ub9nzXcjrkD3v6zCDsvvXOi8OdC
IuVegyiuwkAPfUVI/BjwYmsHwr33XL5j/x0RBVMqQhf2TO5hnZfzRqhrlm4q
yV9j4LGDcRH2ObVoo8WcgcAKNaDf9+BsagsZNoiVa+52YWHG4nLMSYNpWjop
p3ctnkHOHY5Scgj/xNxqYdFYh2dNCTpNB/Q+ehTKRNjylubn/MU6ei1iN3f/
qWSEGrBq6ByuI4NPMq5LiN2wsPfYfG/7iS8Ylv+CcNt0tTJgV6tL1QO1iEBJ
UysjtJ8olxdW1Ut1ruZv2aBKI1Jg0tKnmKh1UsuX6liPNhXRSsj2snjDip6h
i49OoZrBN3YafhtlWNXsNw7/AQDMXDDpP3sZPvjDCpRs8obSJ9Sy1jJjZgwb
FtXj3aYW4uUvdyQbjjN6OhVObg1CrNbmtqEppaYGJ68U4ZOenmQgnp/GdS0m
LDh1GInMJC1U7JHgE7KRgA/KbZidcNW+UGI9qczK5pvl5eXuvp+OjbJFxaGA
b027nmWfpGSbgoJFvFHzI4SLHjfstaiEuxafqA1vQPAcBEpiAnU9y6l0TPcT
ggAn3FvLMRR51My3tsD51Xt/LDxHqC3TYn+kzUTyWS+2rayt8wZxbID50hvk
hOuTAl6sjuflefTYqHuBA8JKT4Se57QOgr4r3IoEK3ysWuOIHplgNBaJBirs
/wyc2QOhATpGYQ70BTjiOxOh9dOT34IiyeOxoEl8UGxjnp9xDVPi2TOFdjjM
aRn0j8HoOQULzz8WNOMnc+lYzR1m2pPYozhFaeSTPmfhBRAJugqTYZX5Tt/e
aNM2q0ovyOOdRexwgNicRhm8ekUKhl14WA42CF3jhDb5utyjAKjyemPKyXiE
+qSPevMwk1F3tCiOHRyQ293+EPWCx9B+b3rnvRwliKYSArQCk+9IGF7cO53c
8QiyGPsBIt14CvE0rseA/wGcVW3SajY7ut2TUBlLI4EVjCSYaY5s2ZrPxNm7
fi7QQpyn4xBI2Yg7WkLAMTcEuafBYMLvTWKQffI9cQkctlJ0C3vnvlUmJBiO
5hyRPl/w4Ue040tvJJEurHLmVs/lBr4Hh7Hn3aTBC4zsodrwSkTXj8oV4LUj
cRehRiRtizKajQ3TGSuzfljCXLkmtHTKGyRATQkdO5/InP//WvdBGDWPJqMF
b2wFV325ufEQR7Mn5MFdvdynAEPGyQdZ6OxMQW1q6Ht7FThSDaEAvFztJ3KZ
PgNfHKLaZD9HaVbhOqyLqM55GsivA5fYPCxroewz2kkje75rsBT0LtaA3ljv
1soxEK6FnIJNI0DvTXP57XHcf8IMuj82qngyA8N4axxq7hzv+A8sqH5qy8B+
c08jRjLzUF4gFi1XMPuRxelY1ezWvnZ7y7KTlJrRIqJZ40gtTaq9icnWRize
rAdDaLMI2EI6FRAh7HdPac3UnVR0+d5cAmuic7jkhZ3V0JSd1u5nOqvso5SU
ItOy8FVSktbftapBArVvpj7+p9Wd4HjgvwP3318SslgE8rF392j9x6CquX83
mWbIOm3ZMA2LPXDk0tHeMHEpI7ZiQPyCXeZDCh7E/eY4KhuZFUCbl7isaXfd
sSgMvR3XbahJ4VqsflJik9c5aQgEsCYNeZY/elLLEbnnLzsrKVT+UWfWDceN
o3JWfpebJoH4y4TnXG8Ct3YzfAfgZ1Ca8YLo/dX7R17Km+46R1Rd0XirT92Z
eLgf5azTc7dWfvgok9r2RKwGo1nXzwiKs3lZ6kxnypUtUqoQLtYmer7+nThQ
OPmLNaavG/57exT2JycWDd3PStyP5ZxRiz5jZWnuikaUIlwUE7VxE3qKtbOR
Ec+V3pDQ5rMV24y/ORusO5JaZmS5LlrCLQ8WDalRPTM9UEYJ28gRW+n6YK2w
y2XeLnGRuT8wfVzcXa3pE1B1DWdTyrpJm4QWsPjy2nEL87+783NlAXeib+09
heP0+fvQaDhiSJwRC4QMVnmlOPbQrn9jN4iB2eW+ReBwpTY3ScL/e/17mQQ9
BC8mlsPbXHdbqecHuUnhyJ6z+r9S08TL41epPOMEgPKtTH9AH3RnFj3kcBDu
rweB2NGd5bnktK1kY7UqTqbKNfbXKHqepDcmqDeIVXHf38Fbaefb6eN43Gvz
ikQ/EmKS7Xqr+s+Gw9ja8Gx/l9YN0wfgsrquMG+6ymPXc7PI7XJ/S6vvtjdm
8h12pe/4Rfsi44Ij435EJHEnql7X0R+HuXMLakTWVmrMXf/EnnSqVhYQOdU/
YuXJEl7mahz8R9OVgKrhActRPQoS9sanhoCZ0e+F6Cqfjxf7NTMPTiARFwj7
WA3OYIcY+wkD53Dg2E81lDBwkXRY+djuMDZlH9QRDn4DY8vmqJ0JHqtpvURq
BBxnTQ2jPcNfkaNMQkfmk4pGsrl2n3KxsD5JnYmhWGTfdcXO7vxeKNCNuO/k
2NO00yoEPFaWENy0QABkKjk4DuC+YV75rXvVEVKL4kXTEzn7KeJgszvpZmH0
OqQndsorPWpykehrvY3k53+Ujq8Z22+E0F+LgtqffR0Zmdxx3KHiOuCDQFbL
qWgO70TVcl7/garuDQHPZfUXAgM1nAlJv0i3qfxj9tyqWIL2f1jXRTaRquV7
NEqwdFex5/Zr+pvUNE+lWwhDOArrhzn1z/OTsqjjs1LoD2d2UWVAgKsEB233
yy0EwgDGCDvMqvEZ05is5yvuurljxu/Pq4USwcH5c//+AdLw9mvH5jpoKv5C
H8PqkK7LjjIpza2vkCb5x19/v2ArbXzWND4Af+62AmTku482437Z9QElP7Yg
6W+e09HI5oYQrrKp6sKCDryQaQfbmx+RKV4awmajw5IKwaeBl9jK4grxQlXk
kVeIth0fthqOnPALj9YzjkwRufAZJly4A2dABnrV65e2CqHyGHP//liRfze1
jxub87lJpzrnzy0T1SNRVOiy8C5Ft/mMc59Taif6PjCIs7HhtexOh7CZNswv
ZfQlFkDk0p/x0JiCHmyWSQ9EATerTesHrSHiSmS4TG3FbvRnlOZ85HpcSyv6
C3IdtoiZgTHckU7soUN8Nu00UfIGPQpY9ExvGD+Asvms01YjPS8mV36mXNtp
6LGbGexh/en/2zC/cEKgvD/cOpad98Sj6W2SNOoBFHaf/f5O5ZTp+4OGFlH/
enNOAli4fJ+7fDUEWrAh+IQdS1VigweugNI6YK66/K5jsgDUkXz1NLHkYsEG
PMd5Rr1ix/Hw3gWaWIVlOb2QQBUtqMbpYvOi/zTSEDgiyRtNt62QBmOceXVD
elM9t9kzKmzuBZDAjhe26woDYuiicg4Zo10V/OEhJB7CJ3MJSSaHl8FJqfJM
/XtLrW3K8ZW6gsJEP4Q2hDyfcT7F2PPe5BWZs2sGOBuNjvarZxQnxCIjlCcZ
o4LB0H1zm7XR7+9UCREHGO4+8U3WAyf1XDThipIUHeNV1koM/FXHgd32P1TZ
rJxCJd4dD3ZCupPJ2MugWjcri7sn7e+uy5Si0OM9XEN+xbv6KiiO1J29dLOM
OMPTmlE6UhK9zjtuppa/VoNWNTTUjsYKQLcP5VlqDMT+lG4SK6uGr6cNrm2+
DN1dDUlW3DdDEOWBvE3z3WLjiYB+ZYymcPSD5VGm+d44w/l0ZODXuuW37RVY
Pf7AykeY/ZfXL3/eYYjdXnuMopi+jV1k5+VLAVYwCw1/y5wMI/fQLYEQqc73
ePDdwnrRoasQrXG2w942aP7F3RsVzaZmrY8Gp71PZOdCUN6yH5fnCc1Bf34U
/o7EFWVwKZpxH6PYoC9rAy3RwP68v11Hqo6M5Pi4004dDkGwySKDeb+ts5Rk
vgLYenZ2eoco+em+5ilpbxTNuSW68DcIO44hiXO2S/EdmjOAbI804fE2o180
h3MKogxr6FbGmbe/Y5c2umks5NkKjcrKBk4/VtIi1JWgq2Jof+4Fga4KH5jv
eYHjO39LCWFC8fm6VMvaPThgMx0cPvckG2kHMGsbFTMV81ABcuoaQ7nBz8+s
CY1g7kCGGfi7R5arNJL1RNzwmNPkMwwT7UeZ7gWsMSo9/9WdkzvoM+ZMKWTe
e/1V3EOjdz8YGmQHQB1npC0db7RtjyBAB58j2FAln/LwltF0WfgyqVi99Qc7
c0veM/79wiKU+7aigNbpQkRdlVUG9Mwm5YduT0bJKAxqrbHOLJaVFidPOOrM
SjHxcEsM+jCqR1+5IswjIdmss+pSEOU7x1OV3eKzQjL43DBZeEYMlzJbrMLr
rsUizMSs1a/MHwS6GXBng7vXnQNcdwD55D+62SGj1frhXj5sz7aDQTH40JFk
euNfPo85Nb47yzlyFk8sVkvyxEaik3PZkoTtIp/7C2dXiBECGiBwSv4dG8K9
qt058TLCxrMNFOCLMmPd3P3A45s3w6khKYdcNebsrISmfuAM8fJVamzBO6aW
QvqakCycDSuPjsAih0FDpdOuIYW5EfFP+LBw+3RAGUA3Osw+hIxx1FZl/cds
1rRkpHqpgTPWzKzqJsnWN+L43Ft0QDxcToKNpIbEliYYBDRW/KhXgG/ov4U2
j5gmmA+rZOFV1ui3fXxoQ9DneJqaobEXDyEGUGITCDFpG6RrRB8mXPmQP42a
KDh9VUsRGn+mQBVFlWD+ZcY4G68Z613qQtOEe8rtPTTKwCrafAMoPp25kQN9
5gCD3s5oRraNz63fW5tciiVMhIidQsa5jmV+1Twd9SEnfN3H7khVJY1dydat
E1hdmvSXvXBK3mLPFpHLZptWs7heqLWFJ9EljpsGLu2yeHeARaSsH3BKTWkV
b+CaDO0tZnaT40cOFb/miPyxElpfin1deXOJ8jjDdjQeIsVpWWMoNfBSuTlT
rOayVkmTg5d5PgIx9XblvjY8wQuloV7zpISUUlBqC6414lotHktoMIVDPZVk
H/Yh03cHWS3WmiBdIGfSojzFSYqty3Ly9QuUe/9eg16majtuUL59lOM382uO
6+XgLrfSrJ5cRhWeiX6HzpYdn+o8FdWe6HEM7lw71ORjltBWWYqyCN52sddh
LVcNE7+YTI+9WDUi2XDwsm9YPkm2V+e+06I4d0W2fHZQ0r6U4u+jI2RWlAkj
K1r6uHJfyyl5QuIFxA0+AXYvbsMIj8SbfAuQSdGOh9ZP4a6aBHlwDtQeZKGp
N7Yz+1se2yRrPD+FzKDj0smjdFkZCdZaLegfx2Dg6nAexfq00KBoWhvVnKrN
qBjM0HUj8M1u7wyMUSkWXrcBNcXhh9jog6v0qfcIYCaHPG1VLDxUZH2EYXnI
wUEOLKPs8W+AnntWD/4T9Jl+1AZIx1ClEUUdJqYMUAFDm7syfAIGMhKu3nZs
ubl7NBYUFu3ywXQrMHzp9fUGFCYyTEn34P3QQwH/VuToA3n6H6VIhEtzYb6j
2fRhcF1+B8k7x8e/nsOwVGXmfXxiotFRylrNkD8IrpLT1oqSuGgz5FQY900+
nlhAeOQweyymGQ05m0FS8sVFWadR0GNg2GIwGV9PfNOjDu3xrRCOyx1B+Pge
cQI/oDWtK2Vtg9paqVFInSZ0uizI+hPMvwTI4fHZWU3Gedb102TxZ/U/IVGL
OT3zRHNWF/Z07n9LZf25GueIu0oIQP7JYRBPxLS/yLg76nTltBHXberLxpU4
XuBOSNXsiUk6w5pGdYQ1FBgedKJc9D9/3nQQFV6g7RzPMJ7g0nysehTFqEqd
VQccQnsNBnZThuZ5GFxy5XfIP9M5zm8t5gjAEMblSWinNlWVX/IGL67KhnKz
ZQA1uJa9Q/GP9tlkMorB/+DToWFp4D0JEWsY/WQUkusFYFJYH9nERHFNQLfA
/hDGZMPiZGEodgRYpEfKzEJX9NPNhs7Qt0sx3HCJ3usNTd7fudgcS15+qaMo
fAI7uYg/Hds2/bTuLgZGaL/mH5QhwdPa+0v29u8N0Ae2gdrnSiezqhBCDM5Q
kxlz7T9X91INwDOqfXN8FBXIVca8846VQnLW8rmhc853PBd+IJMB2LHPJ6z2
XooLTyEiYx5RUJJ+umbCOpxaVIxIOAyvfZuBXA9jwtEZi5QmTCvgzhz6qGOl
WTtwaAqlnRtGmv6el5ZUIl32q7dyRo+MN02m8crjvosY2E+hhzg5w7sH7Bud
oWgcW9BksOq7f9iYqY8JWZNFKqHMl8qhp6TwPKgYIr/4LFMe/3z+XdIE7sxW
rnDvwOI8vEBwofVTcRs3WwTytj5KgdX4XNMp8jUgAvFjcqx7o6DzPU0urmAT
f8KrtgrrEB2mVsS0Sm5D0Jt+6/qX500JF/VrdY1Mc+t4P2GJ1SmvEdG7JYrC
csH0EObkJr48MqZZr6bcVfH6IiDBNB2wB1nCyE5saJqEVYw966oALYv2iKS+
ZIc8nIZKy5J/nAcRudPlMr3de1Dn+0Ey04CF0R29uyOzE8MgKPwis60jDYqh
W4VuIcjAm9op8i/tNuPsm7sHPU2Kxa7u2cjdTXaEEDdurH7lbxDsDfd5bxbZ
ar1AVakOcccdPqsVIR76OeCI7L83i4QJ0bdp9ZlIv9+uMuzlQwS7bA4Qjj7s
Ke9R+J3hM766bYBxxO1dwrFB9BEz4Xl5WhtmE9v2H9hz0BeYwXwrsXQu7SBS
76FNsFvvr4TZdahwMZq9JLhq0I7oCog4A56JcpX+ghbGuO/gUJjzCODDNdUo
DhVI64ip0GEgdzNIDkAmDx46GQCJTurrETJx3Mb/6xKNj2GRnyaMdTMaWV7v
rpxZjWDW5zv8jY3C9eZ7D252bbtzocMiuIh6RpOGhPwHSmPK4CWoqJ9Ty3rH
Ekc8paQAKvlAAmJVh64Qzr/zOC5vLttH/OZ5JwcKdgDFZJ8O/liJeYJ/AkTi
kDf8Z9x6BnMNU95JynHmNcIJWraFjzNJh05gESyu70zVryZ6dJnTYLiAXVoa
pSQfD8+wDkjS0VG65D2RAdSES/PrfKl44p698hDprsfilFt5x0Ts5PK/F44P
fqaXQ29CEhEAlFd62FssPFwAkkPPPvYDO44Xrbg65YBucJxxSA2mIqFifLuR
1sM50BJkQOPhkw3KvtL7crJ9vJM1pFHS+VDjIJhVcPfP+VydRS2hSE8aWMDh
Icjqc/aOGSyAwWwdhO9UfZ+TCmu+kdPNODVIPKMkDD38s/YrQVJGzQQIhijz
eXjmgfg0QWARAgwshwIRZrI1uD8WgiYkQVM35JE/TzohRds49T9fz2GYjPsb
TZ+nirbiOmaqbmfgLbgsU8KOfWjIHuYHSB0UdK0BGhKh5BGAVBsKs+epOqqB
499WD7ZzWUpcTl5q90170FOgvjk2cRDKPj0Bb8ab+DRHEPuIyj2Crk/szbab
2F/A2NTIaDJ9ofWc9/toaugDyllmsnEW0L13w/aiG4uoBjHsvGI/Wlw9kOPV
VrsVzNUZnNnkOeUK48w8c7giqO41rhkRhfEmUp+ZdRkdRGfAYlUPR9ooPnfv
eI8ISec31JI8LQ9Nv16deP8evZFAJnKasZgTaEzTI2qOgyak0Xw8cm3tyqYU
keJplloOkPRNwHPQQX1rtJlJ/TLiFa5mOHtmWnICwAjI0uVSdxCDhevLQxRX
dhAHY8UYDvO4pmOCJIT+USIcuqNMr6resJKuutvHN+kuLf+30mo0M+DBEHf7
iQRnAm3RR4zMUiLVv5/W3FoRNvOfgjJUJt/UecN/W+nRvARIGOEO1pe5gX7l
lkGt1yMbWrJBIFg0ZVTIBDDRwYbbrfKsR8iV3DH4pEsMLb5yR7MxglkWIYz8
DTcc+3C3gdEznZdQEo3GfLJ9zq7xmTle1LtX0bjQJ2DtJDKuHEcnks9OdFok
Tei1O+ZZOmXq+w/iZla+tZ54yMxP9/uAh1u1ZRxl1+wZxMo1WT+F/M+gZ5Qi
gdugQrpaigyGIl812a7K9AHS1osGCbbNs+10SvdHqoYikZtirFF2To0mweWR
XgxG8Fe52UoJ4jYegGZLx4i9iEq+F2w6fdDOITEIRX7yRxH0vhJQ3zk+hmtr
UA78NiXFI1IaDjUymLXgr7E8NupIi+0OaZRDB3fr7dxPKWK9wKysjgO+JqyV
xzfY4X3nbPX1M5Qv65uMneHC1DMpDbsnf9gtTfJX6tez3FRTU+oMLWWDA1T0
sXfHP7/y3R5Mo200NYM3U9xrr/J/bNImeohsozcBOm+H1Xbp/tSWVOHqOmuJ
sD6NZOjEuynLkfbI1RMDRn5CzlGj8S/2CeHH9a0m4YwOmS4hJdHOmzrM5xC0
BptmSiVm7PF690Q2xZ1OPB+Stl8z1N80Zet6GTR9pajvB5qn21da+X2X/WbE
Xri2nb1AP7aA7ORg2Hkm5OdEXpDCDqd0qfjzHWBsF/ln5lUyKY040Zj/bXJ1
MMgQ2vsLsHN/MWaGB8UWLsTCG5D8q5UlVHYsq23OkbGqVqfoE9diubrUXfEM
Gmnask9wR/UADxkeaGwx+Yh00uIG6jv2/jhRLA3gWF7DN1kxjtqwwVA8ratb
+D0TjuAlPo3DGO/ph98ZNSJyVxmowvtbUlrEP6wY1CLFMCOWoDebkKv9lJdK
G1jOM9Bl7aIsudWku7zIeFtelXSMq5Z5smBuJOOsE9Nf7c/ZVSp0oiUox5gx
2baow8Ff8Jexcc24mq6XmSthzPSFCscogt9T9h+T2XR36TBdEh2SFXUMpEsH
oITlMdhWFxSPqpDv76wFEiLOCPBaM1MVttwYaq/fxXbg1uo21X/0YcnyekuM
JW9uHr7r//RYRDHH5Tv0EGuYG/+AFnI6SHzy7xzQ3ofRoXUSNFjLoP6JE0uI
S9Ln+8R4Xo6Uh0Fob/DjLbEzqYwsdNPVLvQaZR+f4MvUAGJtzPkoPRxwWRcZ
FaDZvHT0GSgDqJXmYEjFfjkpvFSfEXh0v5pBlZADcx+3YXsQvmXIwRWJl+I3
dvmlqoY+R/ebTyxeUbepE8HWncJUBQXP32Z60RFs5qsroG0UzUbhMM/8zQEE
rYyaIlRs4JPjVW1aSwEDxsisUOMXpDIL03BO9SBkMWugQhUAJPqyNf+n9gOp
cIJfSF0l4a4mJLeBYEStDb8/B5bAn9X6hkpXq9hqnZAxmDy3tXpE7/2wzB7g
6boRqZJHB8gkKJBG8A7L2bj5YXCl3vvipoxiCFXhvz/7m179zuuTW9l5I9pl
vpJoQ2Tp4kDuFME6qPUNwPvzdYvjHLvS/mdemEWdxacQWsw4H3CdMMPecadE
ay0GnckyQ0ZNrypNrtBn7btb8W0SUVEcV/auE6Q7UvuL/c9kf3dYEzScZ/6g
TzUsPLHJuy9WhgXIdpmZKiz0t3UmHe8n9QrN5NliQYgp6qyh4Hwb89MpQ0y0
Gu7k66qA22wEHq6bR5FQFIWwOaBZHCiTJY9+TIFJx4wF8WtRUodMW/hs/sP4
nnGXFZ4r1Jx6tvk+Bc3AB0IdPn2mfiPU8snll03HSG8YCC2JY0f6OGdkreA4
G8zV7LHyXWaGSKH4iiWSylL+QSVl5ddNsrYqWM8sb2ZB+Z8XTurLEtys8oV5
OlLUdquBYVrbfN5Z8ICgqgXYQvNVZeTsMISZREsweAXZs77W89L0FuASoEEI
uu9w5ywq+WBB6yK66aiYH5tJ+IFF4HwPrk6ZuTB5SSZAe5+noM+KbQHQZ3Kc
48dA5HrRbkSkUqY+RxZJUyfNnoJ0vbkntxih1imdUZsvSUs6vb+WYI/uu/cp
6awhpo6w5LkxFdEzLu5IiDopHw3ZMm4Gx4dd74kwBWKKR/P8SpJ+VeTDPM6V
748qJ+FbJ3ipL8hV0M+oHgn8/u1bLePzHmFjzZ5Y3dEj4PtWexFaGTrDCGaM
VYkLyokKLpQxRVaFYSAEO+DCgthXIbsNFuHjt1SCmLHvv+12X4DGjmy05haa
X0GOwjo9UWcH5WoXmh0CG5kOhO2dKQw+Jn4fLs5tw5uv0KAfbv9wADII80Fd
T9YwTZCsMnqR8sTbd52NLPaodDxsZNJhZ5TrmcH7tMy94r7nzk/Nu9WjIYLd
We+vkDoaXWSFpL+grXYjrb4j86eI+gYosew8cGVWSOCsyrHJC7fi8CYVtQ1U
N5iUdaI/yqORLuB/KMQSTdUA1ia2tPwplgo/66GfaO9ZajQRPkFILioAcH9W
uXmDvIlA3LHYqubhtD14P84JAnPjz1nUGOnoVoo56M+uegeus9gQaQKUebPB
8i22DrJWvpEbuj0hz430Zb91c5xBNmEeEM77lyYX1IptFMiwnCzauXrwuAfn
QaeSig+wCOwEJanqlnY9GbVS7bZ4oPadZAMRXCh0pcynGso4TrAaTG9siWQb
O/DMia7ODKsXXMZDOGmrfOeTliCwYjfQnllNz0PpojvuLfyjotjjso2N0cJl
7ZuaRut3nfH6O7uasssKGOknXX52DAiloasuQgcpc25hUnMuECDdsgxNbFEx
2JhNOaS44F+NLtc85P6Fg0nao5m6Rbkx+LQdzOfmngOhoc51HjVfVBww63lH
D21d66UB/uqkfkOu+lF4IzDi4wToK9eHTWIQcR1Fgdrk2s3BX9cX90fsZtja
G/RewxrLbsBE+TDkDWq1qAg8wlzbOsXrytMyTeRvWt19LpBJJaJSfi9jkReJ
gnbdd4GDpSRD4Q00Yr1mDVtFzfLE1pqCoMI3pT2q/DlQHOIDLfSM7MYsTzOH
08EXSDYSifax27DAvFUBkhQtWgFNXdE7+rFRE2lmilqv3vAXazRJFnuK4BbS
FQjIYQVWGdME9RgXFjxAozMjuK8Ox3xtbj1QuVauZcQ1pC4lwLDPGX4agVfD
4tFK+u+uNwyuIA7tOUaJDA+nd9LF+nGi0FdLco0yW385rednyvY2unJRm/3o
Q/3Gd8OTY9CJVmu4KEbeYiGJPaadF+UD6elRIUn2loTvvH+3vnBGSO15i3/8
D+xBzBMHdNWou64M/G2DLTJBn8Zg9WdeRtFDI0UiCoQdqtyYVJWQnAp5sp1g
Vo4PIbS0MHQ1KijhxKlt3h7y6noBKF71O0d4gSHq46I9ZivYecfDMDFJ7IXm
H6A7PlPPiUTiYPXGaZ6J9mwcGqz8Kz1ayyeNJNqqrQjbKNkmhtLLg5La//sZ
W88qkiZyagurMEzjRg9XyOx9NfPdE2+joe6iTqrDcr9y5k6hbCRiQpkg1YBC
c7q2nXe/6ZHZzCeD41ofLkOHJRQGpTqUM3J8Jr4lW4FnE3LhHgqYnpIQmoO/
kM6CS7CwxvvE568IXKZpM+faMztfcmBu9XhsHMg2q/uz+RMZD1tR9Lvm0j3q
log5K0DakkEsGo6TE1WMVewWDSdHasDTsycSUD89zBIDwvT8g5q1jfeUEz2w
OGwoijLx+jfs3vgoVKzjJ2aB0nOYPYAxpmecCNvhpsDSSw9RbfdR/MDJp0WX
03aMFOWkFocAlZy85Ur4H+rSZ0OCC/r6WmwgLBQc5XlZ7nmFimKo6GLRumAJ
RD56hmjG9d+Sp8RHGqO7NU8gmIkd/bQt3lliahO0Ls2YWUl2CCwQQos+ebiW
cwbbASCXRvv1DmF2iZAFqxTNmGytKtcFnmn8xQPQT+tKLpauMhY3eg7DCQJC
uq7q0zsLztf7gA5OAV4l3cPMjBb6ULpjIrt1RdLoBOzFD6qMuHxBmSu8jlgl
c4cV5pr3spMQ3/aJXKdFmYvvh8KDS8/Jil/EnbIEMiZsYtLrOypWN10Vb9kd
yVY27ZIglN6+WQ/BVDwo6K1V4l89U8+sHZLBEJc9khokn+isrON5ImCPiuqK
0SdV5J1gG8vwAs96PqF8d8AmI1b9FEr2datk2pXxGcOtBG7PfB2YhpR7R97z
i1p69/9Jjrg0Qq15NRjQvh1sC1gUZlBDaJgN5DHYZTBszip9cgWic3K94B7h
4WJWCtcsPvSDOGmEGA+7wFmkXUAKfZ02RIppyEY/mZ8n8gONP5iORoZzPMBM
GCVHxE43soiKRnlaDtgqxuGwk+hPMzCL9mcjKSxGeDJykt0/q6jcQEWG4Hhm
qEsDQ6ak2rKycYc5iQ9OvriVh1eLC99LFVDed0pMPv9FMTJPZkWG6yAKk5kY
XiIcFHyYZWbOhr+bf4ep+fagTlvrYuhlnCESYkZ1vNVnovrWqr5BO5EnflAU
8a0ZjXBOrKDHz6YkgTQvbvXogfP823DJaYV6oKapLf00oUnmNC1C9DUx2Cuu
1NiFWFcfslbeGWXkf8vJKTkF8YPo954Bc3ZELSNc/PFpfR8w44gCjwxhsyGH
ot0vyZmZVxM172ClDxiY8vZuDFhCsS4KzPDfTwxWRtXt4pO1nyHgJ7BtakDa
jwzNNSgumNq2KlSb7Ms7rs1ihdXqxXAniOa0l3vKvrYl7zpydhiFhX7ixS/x
bvlm2pwI3xJxKnAF+R0P/iMsOCQ2J3jbCXGM8aaNvCwljOkmvqQdcGoOI9Ns
Bu2T9zXtO1uy7AgbiG53fyPnS7ej35elDnwjSFT3ROCZ9U2LZB82Nady6dB3
vj51U2D2Rdc2gv3VaP37HuuuTL/lOvz+0O5fBSGrXoKywmfWOwNFJz1ZCtYY
nDnBZiDSOj/j2qVNVT1OcRSFVwMq7EWM33aKmT9sjxG5s4OzfdGAbU92Oq26
v1As9vHXAD/7zePor16W719NVvryQcdrPoRtqtC3kR63rjpWvXgg1LQKDIDH
aBgcj8o9TcsEdvsmglehGvMXQi7GwiJ9+gSIJKWe9U2oB2ZypJj6LKW/p0fi
wA+Z9jvyNItpISaqPo2cyMImQqh4Ka1yNdGM0s3z4aIjRT0r8aQQMyNv+uYe
kyu+xj8ga4/3dRPytXpY9a0Hy1LEezN7KFCtMdViJkXYEPyH4fYu9+zeSegi
bHnMt7k8TCzbYXx3u6GBV15zw8dhvDsvIDmLlBqkz3y0qFsyyJROuxCeJUz8
rl0pzKNMa3eC4CA8CyCzyyzbzIKISDc+HnsDpAywMdWRxzBMIkY/KNt34wEp
bWa+qS8V5JPEqkCZ6iqdaW2bHoX/XJDrEgec+s6uRVCymmcCwhd1t8udcZ2x
vk1cFt5tSy5qPVGJna7RDbVyAzTDPM3SMmKzj8TQHUJoOco2iRZJ2loh2A4W
yWEHfxZoaCOdVYDtu5JSfx9pc5ZkD5QZcTwDhCrBA5sZA/oHE2Aa8BJExUwU
h5RGT3VF+0PgJb6Poyk3U8H71kFpoRbdM6fMuaaGyDq6KafMdzwp8rpV2yK+
YNW0eOU5Ynnqy96DgGb6N4y7lq5DnEZfZ7kpc6PJ+RAwyP/Q1GFV20vEWT4t
zmhssgbmDEyBXUnD405rmR7mFuvKqUXd+pIsyiiqRdaYnMWKt8EKBVOLcyJY
oRK1KZpWhZGKVPOUo8uqPLw/3n2xaNsFZS5bx7rcBNPFsCCqblMvdSA0/mQm
lW6379WwPOjmHoxtgVqfeqKOprXjcMuObiZRvH/jATAcZ3j6X6tduPXjuzIu
SfK/78Ary2Lf8mZ+LILQu96/JJ5XuGShpAuHDr478UfFpNjFWSJH88tUQ2xJ
H8cOR2xE8L6gu4zIMr8ov6lZL+7xuc9LCkq4FiyLuX/yYBxJOuVMQmgRqSkQ
wngCS6Bhw3qN/xvGAB01KORqsbW+L01LkFSdM9/5SyaoBwbRjXzA3zCNUKZv
TflN8A42Gu7qNsTWoc62jFAQEFDGnCmJG4v0QuX1Nib3SqpGi7b2g0f1le8d
5MpDKrVkpObzY8rVSJMtNheeBumhcGu3vhW0Ni5HdXDioZtNIvHop2iQ17dX
IUciya935cJYwhYWq7vQcZ2C2GHBMBFKwgPCz6VgaQOq4bRt9Nb9KAdv1Wks
tsKVXB0Ux4MCOkAWEYNGptJu4GQMANeROTD829tG7o0tAXQVl9rB5z1nSqRM
+X2FpZGQGQfMX20Oy4sLar/SwOMQQ9dLXbNAIYZV04Y6v3KFoXJNKT9A3X7H
KSSoffo0Rtwgbq8/aHpa0/9z1gDHLhto1IlUXZGOQS+X+CRBxH9At5h8UY5/
/haGYqiWQjXjD21Jw6yEA3TvHd9qAo1b0dDDMoVQk/s+zeIHWB6dDLOG+rOy
EB8fwvrrAMhjvgw4hC9kGbRDOgfT38iAiRUmWGPK3rPqX60pJepP4vSsIRs/
pkIwJ60U7EJsYjYBzpNDOOHN/Tu+jNva/vM5x7DzZkBgre9SZI8QSofa/KyC
6PGc1W56eLV3N9GbWgOoO4ZphqImSsZCYfRq259F0/IQZsE6CagB1xa10ZNZ
XpWg7WYKTZLdmNYKsK7FsANcLxlCFztPpWvc3K/839dFLrAyQw5tzSohwmYQ
672U+aAgmmgxh910DjcCiTjGncmnc48XXfABKB+XHIV8kHsKYDJxIR4zEaqu
oyAzheXYkB/ImInBlLJLQwZMZugurXeVVxDDf7Auozptts14vuYCEG0Ectrx
ukUdYv3/gv7Ar+v0HCRmTnUbP8tGMALpK3EUi/2YK/LT0FCPFJBqSzWIHDAa
pFUQv6NHqMtEa/lEHz8Yf4pi2izvqU34m/rAulxTDz9A6Dp2Y1E11kP8jSWP
shql1eAkuafbyH9xxbST6UDFZgfgD0MJwU+1jRa/45eXklUk5MfsknCMnJQN
tivGsSHSCpnWzEFLs0ihYSdZY8mS7j2L+2Wf29OFhCsclHutNNfH3bPyKTm6
hPOSp4iPAzkIZUPSRX5H8OXHxGGPfr/JEk4mWNRO6De8Xgw0zUt0SUL5d0bJ
/amX8Ql0bxcYf5uCDLrVAfb62L0vVJdp/ZKngZis2jB+HYqy6w2AHPkpVtHw
Zih/MK2xlKHP+RyaaNLd0+DTVNlN6ymbyjTD5VfOFG6SxZRedV/NjwHR/utU
BahuE/qgBlJfOfPoQzcl7LorF+rBjB8MKU7Cwg+2guPRNQWj2o6EQ//2m8XZ
hRljOKkZjJ4YgsOw6F0eOP5yb/o7XAQF8G/jLBIhyL1zJRjeXBuT3AGDfDPo
e6+7Zd2gCqH2Qvu5/SM3UQNHKHNIoeToY748dhXNCzPO32D1cnyN2COt8+VL
RM0K1VzPUF95rCTNAfngq/5F4bgqYmSHsQdirVTOMGjmRKhwbQfpF4CqKA0D
LsAKn4w1gKLpXT6PH4HoaAagC+g/eZwpBGSNxmb8pZlxOawrBu7POeMiNcVY
sZQV/BCBwlcfA1Z/f1VqdtkP3lNX+8oqJzCGcEBTO+sQik0DRaTAT6V18E3H
5/eo2AHxNaE1dkjwNhm8e1Ie8c1lRAx9Zf0DWGaUPyEBRrIQGeQTeMecLJjr
Er0+VuorufjG/2DUNKMOLwuUeV+cfKAOMVcQibcWE4gv4OCWe1oBYi0AswR+
8WuC07k+v2lZfrlFdVc8xQWJhcHBQQxtWQ4gM2EGfS3XcEtPuZM5RyCkDBb9
7tzHIotmr2aB1CCwu4pnwES6wIp5GB/9FAVFWsCJL/KHZNVvs3p/334pJQnE
KsumKVFpZIEnku2hrlK2tXOb21q++rD2i2JOJf3MVv2wqmPQUHWskTUYZuPH
hSL4Uioolzte+W2pZMdsKVspe6/Vb6I2c2SmUiPB7e5flNS8lI3IHOERfWWw
oUkcVTWXlCTvJuaLqpDn0EAiC11bTzF+1QEnjWdLsW+GUtd7wr9ePgKE9dwD
E5apogLD6q38L5y5y7PKnjj/gBoOZTV/sUV8ugIm1PsekiZOI0orYLInbva0
yjxmkxcsg5WS2RnnlPOPQjMXNEGp0UqVoluS0mTPyPvUYZ/Wy+sRG3om+KsS
WjR0x+RwWaWeOmYAfJxQkOxwY/ci66aIb8RKIkHyqNhyrge2NrUy9SG1gm7L
DoIQxfMcN+Qg/qboY6r7vMReGYmO4d/0ADNTLYkRoNtgstXupdmX9VSlN+9r
cmY3FN3Q9A8Tpop7kip25sNTWeV4/5l4ydlgrgTDTAFaCGSwUnbl/2GX2Gnu
46YeXAlUjoHkQ5vAdt744a7atZ0f3LkuM5R0Y8eDkX0iijGYwbWnaVfYWkmw
OelwqXvv6oi+tCv24WhwxdHLApADLnTPSGwlylv6HnyZQpYjR+fH3+C0WAyO
0Smfzb4n/+HQ1amXS0m+60PRfbi8wWH669zujUyAuSlGPB5iwwyhf61QTPEl
MzvlrDelXjnoIKQm1L99Xlq0TjFGknmX5llmb6RQCV8NiWSn1e5KQDuAiNT6
az2c6U+zjkZqH6/5EiC1UwrzwyEPk0XRCWjrtKZ0TYe3RmQl2x/TOG5yLH1f
nDqOiey3OoEnNosQCdU5mX5kE6SroZ0QfJK0U40VpW2qNLe8CNqQycWIO079
lXtn8Hm5kLhEgqgR91JSJnLM1If4lHXwVmYXiw4OvW4UTayW/0ttYdWfQWSr
mYvQ7HEptIu7Hdoj+qXJzdDsbhvMqSlU99A64Try1xNP0OKnUYk1/P0Jq+O3
puk+LFMXyVkToypl9WisM19YjxBEYmPj3PswIy30JM3v+NJwN+vIc1EN7cGS
r+JvtlGpQYmCwlo32fSt3+uP8sRCCP8naqoi6AM5gGBng4mDNs7TA4Mp13Co
8zdcMmdjuzyfkFP1mi34lzYTzOla+CGqh58U6WXaEzI/A8tYwmW1M7YNAHaW
aXmMJMLB5XHjeEAH/6721N2o1gAwHkUgZ3CoDJG20ObJdGxkAQGbKcHymMMB
XdcbOhQuBz1PVgMW4NwVsVdVIeFZJATOZJc/zrwCqNbC2o8nGmBfYFYRSs8q
KlYN+xUV8bNr2AoCK5N1DC2dDXDcR3gdG26ZPCWECN5W3jaKU1sGMfO5F4nP
UKZEi5YDIWJI/tII5xMFZcjPWZTNPNvtBQvm64FT6tpDoqz/9Oy3SXqt69cK
laowjEjzRv4zJUhqln5NYRRLau/3xiVRXmTtp76xKAcwAdZ1ARrkMWeELLgj
9vge7sY7TMR/ycFK7tZvjQX9xZVVoBfCoCNAogH1KTakdny+A26KchRsDM1d
PrfbKlKBB8GX9sXJyYAhBC2wH5kD4tbr3snMQjJGnyLe7Ul7XpRsX2x2CGWC
HDpPfNeXwLtyFqADFOTr6FWU0nIIIaYuMwbfTLCNWlRlRlAhia9PF9i4abht
wg6t8gJtqD1ozWFDxoX9wr7MXF2D4LD194YXICuMAhPVvE5cwySOf84hG6re
mE1CvSoCFa4qmktErVYe85it0+sw9Oib/L5L7HYs+HOGDrFEfLASQ314nWv6
ydQcwjowA4YFg19HkDyQjwlVe+1J4WDoKl3p/DMeJpSUhfJcs+vYCMitR2Xd
mElK8zXK4ENSS9QYaK8Y5cGn3bgyFR14bCma0W+1lTy8E4fvt/Ipmy2GjPXs
REs3ovnpb+MGhiNrBU4P6ZLNOkC20R1hVL7GoCDy1ksMHVpczZSKhqujCJ+9
XNf6F4z9j7tzlvDNm0ER15CX+IXgxVkfjusGbx7xs61S7iO6xYK5Wv/1G66z
n5EEfQQbtUxeMVq+Ks5OSM+YZtrmwXr56L7INSdFrCvbF1x+Xy5YR9hGv25v
E4cY1uTgosOsANxoPEhiLNqxyQgXbF2gG87zJG0qVjhgIDUogeHPND2MOlJ9
sQhrR3XnxZtppIynI6Z0LfowBbi7+7c4KwWZwlzK4VnONG4YSr7CcklNcR0l
bmg94uTpnRgRj43xImaI8gu4h3Kdg6ZL1F1HkCMiv2Q7BRv5soBaVmrbCDxo
TOFk0b3oogYtWtJE9zMsy3tpN9cqHefL57k6hYG0DILhC+AqcF3KVp6b/EvT
gtOOY5EKsGXCckD7yHgN3h4gt5iPrRWbV/VhKgN9OzJvwaxLtgsR4hpm2Tbr
zt+tP8/ABqCU6xT59dAuWFaXZ/zE5KaMEj4lDZ4kfO0eT4j8hvrMn35ztqyC
2UgBZnrsKNwC53Q3MqQiixDDWEAP89Gqk7yywfcjmoioyH07ulmhGwVeZEWz
qLYV4tC/tun0GrTTQn1U0FkQ4N1Q4UV9sD05t8WK6p6qfzZ0i3ls7QR5qFPl
l/dfE/obyWZInNXqIQ6rJNQk6QXlUclU28yBT2tLy3xVXa5vZCB9XK6MRphT
SHc57i1s10tDmf303j5+etLs7Sa0PdX6AZpWDQJiLXt56fX3wM6ZWHCubD2J
ZGG5Cg8OtSekokhYF26zdkhcPxODoStxN8GhUWslOxZp2h3DjxD5txTeMMOQ
GQzR2qsQk52rFvopwF8aq/NZyRV4Coau/KcGXWE6FFgCrzAS0JSFFGN7AhYe
AeUT6QCzRobZvIlUSFBnSCCJTHtB3ka38LWgw3a0orSJwnKEowxrE6DV4pi2
NjnouBZMAkhr7/G3ezCtKGuTcNleMayJ4XaRIwRp3CekvFG1De5jte7Eoayl
6tHvhIz2vfrFWUAs1XDhrG4DRysVrjK2QTxYgpdM/RQZ9PMURxeB73k68ZwE
8sGfh6D6cWqrRm/TwsKc6pQOBZ9YPknM0ohpKdWoRb69nfm4l7TCKGVSF/TN
FpFMfvQe4foNI02XErsqCYziRVwECSC98ajJiMSglw/JJ1jYyAXwGUc7TC/K
bnGXABVphnW7/LzzWtSRRiXYHW9a6Co78Kf4lcPSbqK1HPOCrvoZVguTmR8S
YfaJ2B7Tr5ilGSuE87n8OPf4ICj82Duef10+WtENWrbbnI9Kcq9XZOsJLabZ
jjIJA1nmgWusVYs9f7Fcu7j3/ZRQ4JPZibOokPuo9z1jAz1ycTf2BXJc68yT
cZQ0Z6g+ALh5khCz5mL3IPJGPLQlp7wAJezFMPWGkqxMchy9ujZuGi6bMJMs
sXeI9Xc2iywOPAVo1+kwLcAq5FdKbdQIIEx3zRAei1MdZpv3PvPpHZi1Rf6f
Cm65YtLNoc8SQkhqSpTpdBfeMLJEBRrrQatM3D0tom39DbVMVhW/9QdtQTT2
9Be2zBhULDZ0D40CIkwoM5aeqFd+YADwx4HKaN4nO2KrdD1TzCdDCxFrZrz0
wqHal9dcIkBIEB/RnXOikBRIEAu6iOrn6ruRkCIydxPaisov4pcjfC+Kyg1s
KB2s6ZyzfDWf3CYZWjUsFCOlc98nTxHCL+HMs9M7IPyDHuA2XzUa+qfX/xGX
H5XCpdH1Xt+rL5yYhqIUi5ERT/iOM/RS3QYHRpdBAbxPRKXtl+joCdcXofU/
R6SspXzhkRi4vvMLUl+H888rX7J0UgsU+KqL8KEajxEpWfwVrFCU0D3lRVIA
AyXXSnrnDvzETBK7MU/mMgYFlH55uC8fqGv3xOlOb7zw/nLuqKRuJAp6GsCT
pQ0HBIjRzX416ptuc5FzIKSdyL6P2o4W38l2AqYVroT2LrmGzYZ8DcwnL2wK
0PQ7FEA12K8XeSzF/Ul0tHvou6Z8BTPubK3FLMfR8Wym9WcNZ4eC7j1kH6zo
qaC6ygMt5zN8oiVICC2DeEMr5iAdnXOVfV0TSPwjLyyC59BPxA40ctoFgAIl
LLiQAz6DBSNolomwr7wCfIT/3vSD9Xzq6VkZh/oMoDYXC9vOEibwFxd1XAy6
w6tKyozw+6kxanuSwwL2g4keaXhTHohsIXHd1FiB6qG13amkV7BApFeL7pIF
bhq3aXMJ0xjR8vqysVIXlw5IhlXeKVXTskNmlKwN9Ti5GjOHXjTUPqkP68np
STwDO7wjVfFPbBBT5qJ10FiduhGWcYrvc/29wMBjeoy/VEjLrur2l6L1vJQn
ZYzK3r2kI/xBMPSt32xn478lh0B2l+bCSbvudJlI0fKdN6c1y5/wJRSbVo3U
b2YBDNmM8ilNtgS7hVo0VVAn90vPYjHP+2dh2reNwqaB9PTIdoZBrOKyoPZq
CEMNCDb7t4Fsc0zAX1ZBh1BBvs8OQxmTRFxRHeShNf+9PLi/ETLC19GaHaa/
aHxIGHtZjJzFG2U6trLJeCQFLE8Y3mqiucIShznFuZrMPUsDgDK/qPXyKKCY
qtCZGaxbuD4Bk5tWI8QnVyuI0gqeSgGntk2O5Th0ooeNQMpCKcdVbOh/DfSq
NfkqbJSWHCKioD7cXtR/UTbhDTiViKa7wxsCOC8jd9dnwJCY3ayBNQholGqP
xGTMHAD4Mb+ZR9JCo+wTbJpB3j0nvJUuLhioiumlcwFujxVCQzWX0DOXpra5
ciqKjO3eM+q39CYUmvaSpo2PxWXCytpeb1mggobxdANwGhZbzrbBAI4THWDc
a7A+Y6XP+ylF8tn7kmg54deFMLMWjIx/EgiQVrV3e9d/8MKHwJ+qB1h/D+Ht
Uti+YDwCi7nBYhMQvsoWfHLd7mbsQ4ovQF3cxSF0bv1XEfM/FIRyQ0IRpoUo
M1j/r8XIOmPr+A6Cn1lRnSuLRKZLdq62aKTtowuP4TUqRQemdswHwxSeUOLf
hnNAOLPujpi8IOHAc7I7Hn93VEmEQ9pKZVJ47R4QloIYgeJMIo7ooV/8kZ7P
kLGpwOMrpSmVgSW3pjcUPrJBycBH24IxKfaStyd9AFye6Ldi7nUmgW5nPP7y
lC8qFNjmF56nkX4jPVRCfW2W6YYL1SZYCp3fdWUE6oBlcLyV0TzQP7NOaRmo
t4vHNfka+itoJjIW8jfvtjSCsvaT3tsEJ4blhjCcRzSayNuZKKUx5yFMumQD
T699YBL7KfTIWwUFdLc10ulk0ipn63bBfoL4PhdbmHEDfw4mA/gf2u4ll8ZI
Has77VdP7brlzrFTbyUlJVQiyNOHuCD7Ht+Lyih21bf0uCk0e4Zi1lP2q+d3
Hqmgv/cbwP9sepNwFHMahn89uWpj0ZVb9vNs/YRTLSGAM12o0OBW5EKvwP2G
3idcimtgKq7NAqD3Mln9zg+EgcZm6D5mmGC+HjoSz23HAimh8YWRfQgbjpoL
9EJFXWPfro8hOIJOaVkMkAYa9KekhjDP6rutr/zYgH6Iq+paVCewpL1hIYbt
tye0Ge/ASpSsDkXkCdzUKgcbOg1dfAKqefiIN5O1nbCZGb+WH4LOw1REfXPZ
EnlgYtLYA7/YjH2XK2qSaqJtqPHuqf3kpY0NPwF9/tCoS0T3jbh5yYDL8mr+
7APF8e8rdMOuNKubYDZAWU3SLVvNQ6CKGg/uSYjGRHff2AsayOD2+VKa8iAz
Pk+BYbTaCuJqcZg4Gmv5L9SpJ7j0yZ2c6wl6mgqopJvewa4aXVW2GSC8xdaq
DcH9QJZk7HJjbTtlx6DXoKEcQXC/3UJxJno4lj0iZusvyTUVTTipWMiUvpSQ
X98xySYQ4251B9cZIh9TxlZIabslQFOUB+tFVzvOuv3uI9dasfrJEuzPlJlr
Etr/iim8z54uiyn0YSkpogg0cMLys1tLNI9y87mUn6no5f9835J1y7FUEDe0
FZ60XBJpDlRZAJKhjgGKdJjrVhqQk9Jpaf7ilFarp9Q/JF+NvHavc+BHpznT
JOh96zDjFgEStehr2DY1qHl8mD7dejG3QI552KR9mFjzEpw6JTecRDtVeCR6
jZHBRppz26GmLt2uZNzU6raiRnmnpXwR/KQ6On8w+nOryFTgXCid6Q9EE6yn
1v8SPqUAnN+6ayt8tHLMHksqinHvE7e3GANIaRlMQmjCQERpu7ST3Nxvvv+Z
7jN6GjL1FaoLtmmW9mhZWyTWFS05H6OxRGyYA/xtjB3dQjDpr2AUx3Ln4q1a
5kZz0L82bUaUnLrYOg5+5Tduo9N2eeJt6jJ2eWLGJ0kO3wPauc5gD9l/Eef4
QfNZanfbRzxH0eBAou5l9X+ea8uGsVkceygGekUSpmNY+Y4ZBjQOD0PGFNJC
6ZZYicXU4WuJmItF2WC6ktDn2KvyjoWdvf0in3hFxTSKfLfRk2UmtxFbYoXL
A0snsFKYzh96u4MCNfyaYqmY1It3rHZmEejFxP2rSFSfNuybADJIhbZUSSmH
2ijGoI6RrZc0Dk72Mh1yQ2TUeKL0l40cWxGRTVNox4M7mUnYEzLxBAeaDeAG
OO9CzUgnA1zmfCaVsxNvSinUkUHQA0sgy35cyKKMkgJ3vyVeUzToa6wEYxkf
njhptuc2AsHN/6XdY/y5jAnzBfZIzl4Acf43OVScfiUipP2MKU31IUEOPNFz
icJFlSJcaQ4IoYwjRtqAJ6rM8CkuGf70S39nsgOj1raydedVCjaL12u0qQ7N
kS/zyVxvFlCzNSH+cJAKnSGXVvKsa81vTk/WFqJFjBkXpbRtbbz26YUHe6fw
Ervs1dkQWTy3gIfB3ORIIbjDQnrdZDgCmN+Gav77mtdJ5EN0QfUIg50oUyod
1cmTpy6L8UuOm7lZ1JPBENq8iPNL57cQrLg89elXgy7WqtHLzIxxoogajdjF
Ys/AbVlNmRWzChO9qAug6hj6TurTfJZVGiMHV08XRj27qAZoCRa3svoJ9YM5
mkMSeydt3Uf41WSgacHKZxPC6HYt5aMrqO72uAq9gKWOdnrtopEM9UlyZA8P
d31h59ciX1a/du12U8Uh9E8Ry1AUN3Xl/NKZQf0vd5bkpTsXZkFezBg6R1pw
onPEneA2+FFtOIqC+xZe/QqrCifxQi/Q0nFEZd7zSc1fvKEYotEIPTzGz6td
+sOLePgtBXb/G8Mm1s9xsgVAx7o753PX5H6pSU8UtPGcbE/M5DG/7V+kND64
17AXIb/JG+/gdfEoQftWZwCNH2dzW1dXh6irD8jzV3XSq8ElBUDPOGQws0A+
KnAcTOGsyYhxEIsyaQsV+cXMjrhVsIxJ4BbcD2ng5na3GVZ1XNt8o/PBu+LE
gmVx4y1vdqJV+f5QCoAjpzQjOjvfA/v9Ufk+ablyy6AJ0Wrzlr4QkrrBJorr
Ylft2Mx+aw6ah/lOynAK13LaHjTdJCJ42sKEiwVINK2UmRwVlInZELKqPIYr
bZTOU48ika4cyIcoP12uLACWMTHrbtnRfWOxx1u+6uypcG+y9anA328IwOVJ
yt26Q/nYcq9zUCG7YR9K97DW3+LFGj+UifHhTC1wzsTEiQg3rkUmp4cOEEL6
cwWv0Lr5G3EH1roleaXUKuI3gv3hJAg9hDwXUUcyNIjAELr5kZXec+TKvP7l
IOZ00UPe/c74+tAk6sXe7ArkR6sFVH+dOOqZk87/uwH62nBf4EHyEX0LjgIa
1tH2VzR5KeBLruz45L3rdoHjPea0mg7jm7LPU9GlIRCCC2pZ/804t4UxwgFE
JMoYMidjdMP/Ok/wAAGd50kZFFFow61z0sKiqIeoUaA/BpycyqSyIIg0gZxj
fn+VCfqCTJjhAa3PjclGT7icnT1xHQWnmZGICs2OnHgekZuqifvgDO8F+srK
FydwYX0fOfUKn+k5oWL+6h+avkyhJJp9wWBmKdHN/kyrk5zBGhQ5OxZwePIc
2ML2ktU8i9xssFnhmorkUcHAiSR7lrm49plMdQkhFAF+LDBQfWjPKxirrxoP
vHDguuk59Uemn4g+aSVNTD8AdWF/0WdK6VC5SZwsdr1YPoOERytUuxXZ/CYA
9xEdFl8gQV/E9VBiTBzZ2LdtycrQdbihBWjcog8vnoWQsjL2hHsvW1ILIoh0
JYsjV/VC1HjK6EBqwjxP5l3/vUuszrMbQIvDHL0lJ1qFhSu/J/qaqj3b4UY3
T7RL8wu7sIZ2o+BLvvPSEwUJbN5394ioviOAif5v4DY/TINahMpgfMCElhB2
QK9QHT/beKs+3sOBa6NnacWpGDMw4oE1mpD09HyxZ+v6dvbXBRSkuFR4beR1
sLj9V7VbysvkIcNMvM5OY3igg5I6hdnxebAfSMVeIJbdL3fXHxCMKWC9DI2Z
d3RWVe2jYk8COFxYeJvEPtpILixUmTXijRCLgtigCDf1PxBXNtWOlrO5DSv0
sMwdIX72xhz1VWGUAYpml230xKimi7Tn7liDBRqTtRtZgjQq3iHWImgttR9N
W50Tua30Fz7If6Km8Y0JKYxPxzisbkXfS1i055CrYe31aPsSNHBDhkTVLOfm
YWZEhty1ErLNelcAk+HWE+SSX4uROLEIStKweGnG/7eEg2vdaRR8YPAxWSng
7HsIlWr/10Y9yGu5/2hMU5qnYk2xx+kESq7C8YxQMktN32ZQrZ/jPKu8N8Kl
rOrMuxdgHfIcLNXYWLH500+RYmimJJ6K520rge/+zrm2x3E1dFbFNoG/cYqy
Fy1LMygJ5SRb82cL32JEOCJAWBT6Bb1r4HLgm7yhG/ouEFqhogSuOsh4rpyh
dAUQzlqNnalhqsQFOr+F38mZGFRO9cqKIw7q1cAT8XgMZ0WR+0Bl0uWjVYf3
vjLtwtSPcUrR+mVNONh/Czb6+3ecEKdGDQ28JH2GQP2TTZs5HY8SLUE9M8/Q
zZG89HDwTR7Vm4+nOr5p+CkRhxSGJYXbedcV+RTHb3xYfeb9ZNWWABog5QXg
Sm99IWNyZ9y3bbAgOtD5SZwH6Yh2Zq/nUjflH19/51Brkkz4DGWwX9J/jVPU
rl0NEbpw4mOq1wNEbgHjnuKAPzBtfgKArQBZYS3drHALigxmPzD2BeLBb4GW
OGheXdnvWQsKNx8h3Ij6m+IJ0Hi+kzRtf3U8seOVwZxp2tPUgPYFhe8ldBze
a4gh/CicoCwZnfV2rlCy5vtfoYPxIp+hq/3uVDGT1+wmRK59w0DR5/2HNINB
Wq78Ab+9UY3vGucc2BSDZ+1NwfUWY3RNEnBS2QgJW4/VA/U7L3DV1L7idPxt
/YsJ19IH86V8NORIPcgdiSjfg7q6ngaYw12w2XhQvhQt836SQfsHRAyssbEY
f+Qx8DIQ2AJd+2Q0h/z47YZ4TCyh1L7UF9/g4d67+CizepQLLB4St8eMCsNR
MQMyLkUUxGBT7q+GBpSTgLMRlhaGFAtHazCkSZKEYy2fhr/MvrRzzUtjmryR
1G4brlXoAAUn1L1mh7SnwbFI/WITOvb4+M1QSzWmSeZIVZVOphHxR0CMFbp8
68Fm/8t0792Ff+Na/i7E9TGoS6RMJndf3JKuW/UmV/r8sjd7eK88qyuSR9gL
NmUwBv+xXvfggH2NPVX+QzSCadq2dL/Ky0SLLw1KinO39HQKBV2u2YsZlTmr
zOoQkViluX2bGUKRh2PUqBsGolK3lL4JUVlSkSj8ACpDSSRyYg1wBOmfzr+H
CKWWvybLlpT8kuF4NvcYom7W3vbGVDqJMQAbZPpZ0A7dC3jVLfsKM5bDlCg3
As0PcQovq73+RBSfCwr6IUfRf6U4J+Hw2l1aQD3sFe7fS6LQrpSBKL0mwNtd
0gHlaeeU1WQ7W80gNgS73mcK25SEjB/lomOsMhbCo8NZbbs7yuAzn/1g6H/Y
uA5ZwHg1eLxchTxx84cPbJrGl973Np69QuRZBBLtLdqLd1VzzbYyRLIk3fH5
xygMk6b3Vb6+Pi30PAgV9mgrajC6d8hxnfeIcLS4oFrso56Z+M8rBpztsm+N
R/vfeuaJUVulv+gfhsBNIXNIcccr8byRQCgAf0YNgUbuTR2aOMZJla++yPRy
n8C8c+fukKocfomWRg8Df+9AUauT1YR3Ik+9IDucAf19QmfyBDoKa9iyoN/p
IHNkTekirC0Hqa1bzXqTf3/dBit5F68+zUnn2qh6Y9PaI4u4F4ZUxON/X19x
FmZIInEeEY6Gk2KDx7ELDqIByYvXZzsdZau/QlKI9oWHMhGm49M86TFTmFgq
Wsdppw2MhgQnMbT3py56i4+ThgAc7P7dV81tNXcwixAGWzWIZpvvo2bLEdbr
cXv27Ooif8cXDsSNVGZmoFX7f9YQpPCr6/mOSjcXqW3pRJVHpI/J5Rm6sW7N
t2W+c2U2NsKWzIvrlN49zIIAz835+R+iWyf6zVmS8PBHR4RV/TgXHKrv3wpo
tAmDMx9fjlC5f8bxRsZKIDNknUycwCNcZ9i19CIb1PIdD+yMfCMtW+CbMSpB
6IeQUVYADlUr5Q6J/ObIrkF/Yd/D49UtDyrYkOxEZ2k735mgaEloxnwiFC1b
r5RPwz5mI5kp7lBAWntn7pDCJWEp7NAg8rCIegg4Q+6Dyee3skKdlB0vsdC6
Zlx/D96oOWzZgU0lgYYEdwutY0SPDydTw//8r0eLZY+GBMzdUtZr7veBrA3g
ADWk+XL+f6bVx5bOGR8kJ1eNdKjaJYGU2paWiSn2YrYLlyzrVTw5JhtzY+yU
Ftej3zxzBSlk+tWG9xUHTlnfLwYT/2u1F+t+VjQnFPoZ89eGnPZ4+a0EqPbe
laWcnwn15dLAiyV4dwGvBjvvFGfrbhhqd2prh1mh4y1dhHXoERcpCLtHFzO1
oEvyQw0LWEGpC9MN92dj/kBa7LZPqF5/O0wjXkkyq5s5gPl15gnb1G6S2S51
LXn9DbvdykLmOIRqYp1cYPaij41Fxq8QD3a/qBqK3iXg9kBYmBopcoQmY4vN
IfANwtfwwchgszDB/e6SGHynkHqBV4HD1Q8MxyUGBSw5J6FQCZbS/rJ/cTBO
3syCX0pD60O4mICcfsXCT7uY7z1rZIOqM51t2dZh1jeCAdLMC8v9PPrZrU2w
y1z3jhXuUnH1HbjCrd+QuAeKB6kysYGHomQ43MYSxbhYF51mt5cMYRVb86N0
4043sNZMFRmmsKfJR4bGSXcyIUGlY6l7C0y1/F5oDzIHakx63GdBvUXyZGGN
wf813D7LyjgeGWdLObhgfzUAWFhhuE2z9HHjmlQn+uLkXxOE3vhFjv81ZMTq
BFRhw7vNy9Um/QyG/DSWKoTj9N5Id7R9T/Lxl1yFCwwkwXPjWixa4/G6PcmW
5h9HyVD+Hp1KSCy+p7tK7p2tIqdXQ5t8Ore6pmkjmLkGN0p1xd40n8GP21Ot
aOKxoeOmtbqCpmx4kGzbk3zRN01lGShGBy6hjjBpCPS4zPelnbgJSTU0d3mE
wL5LBQTIpNOL2rPe0gvVGnOlBkSDI1h4WKVdjVV4CM8GMdFxubxweT76fWxI
y66vE5fViH1/s03NuBd/ZnXwGk0jmVg34X6uIo40WLUgm1v/0VqA1Qe4up1m
vHpB8qvBdvEO8mK+jTqukTPmzziWVHJktJ6+K7DSMuclUg7WgrOBhI5i/p6K
EcWtes9qCReMS5fgvU9g7fYOsliRK8wGqRL0hrUu2vNwqUQTaCGpe+kR0YCr
7d66ER2pcQdsE4lnI+DuOiI1kJvUyFGBRBSF/sn4HbqG7+FCbkwicZqHIWAR
z5JnDQtrpgOmRmUKMx3AuJloITMgmlXNw7EbOZRJegSPPktUUbkkaEl23ahD
yItfkMNzInYLju4KWNAnPlkeK0blpVTdyN12aBbpw08Huat72t7VoS0ii5My
xP8h6xhScCZwVP0Lb9kGTimA99xySjGqydsfauJUZXrkzenEUJ5Va8fy/M9R
U1Dq8dSw72JMB3O6HxIf+uXbLwrhnlIFeOG3YuS4aUquVdsZGUIc6Ek/AU7A
sStWIY4tQzFcrNxAao9CBQL0HDeS3AWdpNLNl1i299gxPaxERlI35+eQ9Nq0
piFVm09P7ShrnEAiZFbj9SwB4qWZCyZhF/EoOa6EP5xc2VAbJm5p3If00jVB
mP9SuhTY+xpp2owGbHzskVSf5HQdFgD7L/E5Nyt9Hs6CbPexyXLuT0KSP5Yt
rSqYY9WIywlG7bjrXk6uJUYXEv5KYwAXlOsotuhsDXXTKP3CLK7w0G/Epeqn
gFz5ZpAOrHSFnBKr6/zryhnObcdNU5RP1oZpht2ihcO4uhSPKk5EjUH5lhep
5y3hKQQ4K/nQCzqCQR6YPguQ29Y5KKreq/KnmipZhlLOBUTJN3EdWZNTRSHF
t8J5JlkzW7CDOwaHhu1nelB8UHc3tx1G86AkMipjvmEHvpK/nmRKYin3CXDd
6kma/hNXY1/PwIJe9FKbOPajhwxPruI3p9BOpM8QtAytWdTwojx2cBzQlPTt
05apNcsmmqVEU/lod4zWNOkOHO4XoPWJ09TFCJAcSUJ2QLxuPLgQSwMKga0Z
ZhTdzUOJydBQ61lg1s/2PnOzl2rLSaSBbSkkOQ1HptCjcgU67G9XZlC7d1Q5
n0L7jl5KWwB46qZt8ItfvyW7GulbMdDBhFsZ/JvJV0/m9EVIdKKEGc+jLQc8
rX+mGz2aebjmgqiNVGddlhw124xLzJkZeQV1trprZiQvvkdgQpdpDm1owXvh
icFra6h8laYpz0g/9In4ONHMADyWI9cbz4w/UmNKzWdmLK1lZACUYpdaNqse
qtTAjFX09X0VURJm9+3l1vuOuegIyLQl8QDUmOR9qf1vN95/MCGPL409ulrd
BvgF5c9Q7Yi3l2kK8MWQvDDq56Ei0RQoFZ1mYTr+jzOLQgIdg03uhmsdBqgx
Di4dGfDx/AQtEpnNW/kxVeCnCdxsQRyYLTR4zZugr01+Gq9p77CbAa43Mbrj
b0L2DKKXGR+c+pm91AxBXCEo/3ZrRnY9TtU3klGvtOpcXXltyjwaB3DLcFab
UJCvTwVNbpaSyMzlC1ViDe1vu0a5r7ltIvmH+KS0HaQV4NFfodK3Hj2WsGK6
9Sq+QGgMPWXDxbPeG+pGrv4QVmE8BhwI4HXOX+KCS6vTAJW9iTTL0mCPX/14
U0Kadm6EgdyyJeTxK3EFCloOefvy4upHAIpPxtjELiL/+FUTAreUns6t2UWW
2jHBoe7Pg6a53kDm/K0PfMswB4aEOKl0zui97nDKTWzfI1ya7z5GweLi3IWn
zT1RLQD9zLNEiqhiK9Gi2CUXhHpjWahDKDJSpnFnW2uZ1xywwlqk+Dutd01C
2cmjd38eUSPQ/40hKdQ3/A4cEcF16iX4Lf0W0DM7D/65MKoqIYDvfYIMqnuE
jc2F/ZLt4Iu4CuWRIZriIjVDOKG4FdxEPjhRT0DIS38iTb+huwIn0/ZRrZL/
n1Q/qPiFsooEOYeCDHrkT+9MA+dmuyTwo78JoJEBNlT2XKiog6TNwUbLscYh
pYXGn62x+mIwgsoDJksCawvCnSjN7hNW0IKXRmERm+Z7kNjSzzU/G2HT1tfI
ZVa5YOP86yP+6YayoYhq+C9WOsgGYBa7eAvUra6imEt8hN+vrY03hsKBvx8K
/wIpv8y8Ly88UgrvGbti1vMYHC4nv1nzxlZyE4ZOXO0bFtZefWuA8ccEVSuf
ANFncPV1FhuFGN62AwpOo3IW8kcXg9ja02ZNUNKQGhC3XcE/42+AjeAd+bGH
FYrg2Xfe9phiBRedyRbNkrIKXd/g8SDhBkD+AMstjZZ/OJRH24HWkwlEj09e
lDvXNRoy7PF6qHyIrKWqf2IegZtwIa5xYhrGVvsr48HS8GiDwB/2UOZm/1E+
C/yCLX2Il/+C7baeXSVaZF09Q/d/vQHUbkPIut2f2cfORK6j6wH5vf2tXmuz
Cq6fsp+4cMdhkleCE1eZKirmNWSIcgeD/XL5/l9aP4d8atVBlhUd2YzZw5dj
wjmB3sxnxr6bIxgYH4KrIWUx2OgnvcbNkAD4hWvCT/UOTDJt2VYRchAq6sWC
7jKX2VYJagbmvOs+DdKtdxwv/fOWhAvBw1co8DyHNS04JtRQO7Yuk6YgG5yX
jSZkUeQFiLCI+Ztw7lR5yY2Ixv3yyBKwQzmMBTsjuWBmX4g+KJLkUaXq4aiw
8lHeD76e5SvfLM3rlqBqkqVOzRUFzb26HTIfIaq4dILGH+H4mzU/x4FGWhc9
fYpi4bZpqU7sFwXEjaYzMa5FwVxsUM9QgjYkawER9INzFAtYds4e28x09lE/
OMPN/GrBrJbqFjFQiNcAMXCTbot8MECr+nGCBgPY+15h+G4FFVXgeEpMy/0a
RT6pjup+ohnJTOERCPk/L9K4VeY/YMZjGAZM7kyaU9/x1f0BRLyqKNqd0hbT
KZ9+DXGZ/Xxbi3ckmaH7T95jwhJzwsGVuhwXZ+KIEeCDQpy4vzkx08Omppjm
r37zw2AojviVc9p8LgK0o0vSNAC/ZpCT0vPG3FWM+I71luIYeUf4+IfoJC2F
rcv6rFRe/SgrZvVvV3a7hWNwhtF37q0FgO5od++Uzy/gZ0kdqpXwGDTcgo4t
uKXtZniNkpQ6nLhL3dvkxSXYcC/XEkMabVDmBXJa0SaFj3Zf3MgSsvYnU8Jb
2x0XELlQOCkh+6p4HUU1XnksYRdhTY1Tl6UVzDeKFrooqEKdh4wfiVNYV6/g
x5jfGz5L772YndRYopERhA8XEM+lZkdX+dpl/QcYB264aFofFQxDaqavzZcU
2l+a2zQj5dAindc62T9O8zwBbimGeDsUJ75V6ipYZ39BTWCLtA1FIh0luUpZ
WzR+gsknuQgDKN5gc1ZNkU87esnsZZlWE6uymww9VYzaxDRW81Lfu8JtDRC4
MlBRT5TR73td80pwKu/q76EEKZHaOJ3A3PyRpg0ZSoP91OXk5vgZLKsi+/ir
53fr+53plyDz0fhsaBeia4UMjgtwsmzrfyN5NVs3FBYznAvaKoI8+9HJ/HhL
f7jKLmpV3h638oTl0qvqFjk7dixIyl4/nKMvSQiGPwKo4Kbd1jNvNlUWujba
JF6o9/Oo9pZeANUBULD0ph5EVAz6iOrSSo1MNw92javJrNYydSmxRdAqciWa
77nt1NZ2VJPkpOPbEW3UdWEVq8YJAKVkq1qI009JKkL0fPmbKoTbhnXmKAtu
R0B6hai8SVaw27GeoN/EGwNxcrT5JMi68L1dibIyqMoR5x5sxgvRbbWssvdu
rn4w3Cydd/nxIXFDAriw/PSj34vQ3eqJPXR7afcngigsVDv8tPK9/kNSA7Ri
QVjHlWsYM1/nomp7477JvrllujyLNt7webmDPMlj+jvv5IFDbKB/TPJyB34v
b8xdKgyZQi8kwD0tc9/F60d0LCwoLBiqKkrClpF0zrJiEpGcHjwUvizbh8z3
yS4712BV3X+qJehBLnMXfNAqIuY9rOw7t0EhdRXzAJjWWhSJ8eSpeEki1AH3
tHCOY30V/GI4ugTC05b8mlrl40KfEUOkSI5WcmsNoBWMqUu2VbFUJ1I5vrBp
QZvd6eypbqWQRSS1X++I8yLkhbr8qmv2qx/IXKUKe4hz4VU7UzrIqfwY+rQK
mZRt40MWi7CpAfGyUx/F/G4A8ehwALToBckeKuOxY0Zj4yfibqKRqLIru86U
9jC5OrtNrRRFzdWVpYOnI4uOpnlNA7T6n1ikH1w3hezItIxAgDeWbvpwaBg6
aqs0YGhNDVyZU3RHZxGdugm4Qs6WrOdUoBHmOci2IzfuR0xwMf2+LFTS5AKx
V8DPqlAm4sacLMaa1QWk3dezpkch5Qpx07eBxD1fcW0/iJ716MtPIpNqFNVw
A7swoNFFxIjJdzLrAxBVJYMUci9nX6ZVAoijKZTFNXb00E1JbqUT/3Udbq/s
6mDJDtn4r44ikpUCJ3PSSIfdIawpcmNojQfZT9SE+GSCsbWMq2Jad7voE9v5
zwIYZt6zAko7J5w2gxBqq2IyZo9GADNrOQHr2ZNDb8votP1jl3ORvdTcL0by
0WA+ZUEgBetkj2Rc+rj8RAdQy0QGO4kdNsgp67HTArpowsWQ2jAUTlqlpHCL
eUjKLLwIZRzqHw5MrIQ6MAZeZxj1KTuMmB+YeoxAJzIxt+g1ubGQTfFZ2Ka5
8G1+osiGyPiYBV5F+F8LtKJbKh81JDXwMxarivtn9G/KH7b+yyet2SGbRCWL
aTRJP/3dvVNCnndAPl9/QSSOBg4Yho50WIao8oyLufwdnF4kw5NpJ1VJ5ZhG
LxtvwVCwqOTDQSZqSIcJRFMl6jfmiCO3W928G5nVlCBcpMx9n3nWF/7G84fb
4VeEANEYL/0VgPDD55WiJwJZcTmi2nr4jGuPyFpEGsoBvC8gS2IcN0XVQfVK
a7lVRr0tx9k1zQYt3/2L0StUaRqdW2LjwuM5lzZVanuFko4dcY68X/9zBb4l
DCmXnU7GVy/SSmyaAGwsutFCb5S6omhEnOSAwiTl3qYL1y1i+oFgOYp6FyvW
Pg2XDYa5eqSC7+Uk8k8w2T7pksUj6zaXshdU4OUTZlGEGjdsijxWXII6iUg6
NO086I3kU/s3Us1WV/OGRlhl3nzu5nl+l48CsUmjB7ndhJJAbnGqd7vFLhls
pGTRAYOnzu9I2qtY8u+9OBotBygAyhrw8yqS7k+dfwOO7Zh4PX1cS+StteJl
JgoN76vTSeyHqLrCvdtKy9GCu6/574IoWI5RhDhuAXH+l2EHxRmqtKnBlNUF
CFyTkRTWVHewJBDELX5elK4AKOIiIN+f92ptu/WNylVMopGHH0wkkaEs09Dh
qGeVbOD6lgUZBDtY2NarTgaYugmgEXeETvFBVR6r8m4dtlMdbAadBc6YairU
oJ6bgB/NsCZYGDVuc1gjo9op+H050p3ONcp5cHqTVVo0sh2lBgz64IdMQWbg
ttf42yY/Ln6CsdqK+6nsVwbpbbdTkhHwA7hr7HZftKjBiuNDjJuk8z+0DA10
ZWTAXW3XSktZx42ghVIF9o7X+MiwJvdiUcmBszbwtCZv+H30r3UvS7EWIKDl
jcsDyAd+YEthhSNEPEMpxK7KcgA0eVu1df8fdYWrmE1QXH3W63L4ik8gwupc
M8QasAijXjQx9TECra7TLcAUiEaR+BCT2/oXbOGBoO1kR3s94YbAUPXg+ukW
c35TURgCKQGWZ5v+RQjNKM8fkNLHJ4f3EFyzl6HSjYBXXjV3sPlADA5jUxh5
3SlB6z/pEXpkyetIbJWk4vKxp1mSVgWuPS9fAifuv/hxaeooGoDub4VoANAL
eFJRijIbiLhTK13phtvDmcJ4pfICS8wlIqZuXsPyiMBQrryKhcPvwxHZFhcR
uye3HyFIkykbqwHA52BGkD9qYE6UJpHkdE9YDYd//dcmp36aMSZY2RQ2QwPj
+viIL0wIuj1uUEzNt4OH3MxkNoaEINhgbBigaeBQKjl4HpMpuAIpgVxmZUyF
qYTF3KoIR5m1VFYTz8GPixxpp8oAbIWsaPIiTcuyUpyWywreUT9LnLThuQyS
15H1YqCFZ7NZvHzFreC+54qviaVbd5NXkJbd/GwWXyIBHieSyDnb95CGfsL3
66nEHw0cbGjWUDg37apEch2gu+FYv0FTTJiw2pCpcZZTF4KG+2X3cPGS/TaI
lW5c3NWXfr4jY8oOmD/1uY8zAsmEDPA9SsgMCXzfVldaDj56QVTTXZnx9mzJ
uqjhNveey2tSD0wLIkTLSk4rzT6k4qZIfLR+OehhEGt5z0IPT+7vcHH26H6J
/iZSUQwoKrlvMRStEvMOYH3DfLRgk8AyDdx1H1kRM7Q0HOHMDITxEdPevgYV
o7JRdxoVpoDtYZ3ATOkIA0yGgmcqlDRG7hgPe2bITf5spmbxzzg1zqXY/ld3
/k+62WBypptRoMcBZKIMWC5Utdnmw76upaUE5RuqqXfct/GVJVzU9I9MpAVm
tDlhsF8NlYu1Jnitc0YAYeewPveTD5by4CiUPFdDGwUC1U/rnU4dmNIyF12L
/XFzP6BCbjvrRbGHb3br0paY/7AgUwWdGgd8dqhlIabdhsXaEIHWJ22yeYUT
YE8m5gnjIXHXV5ZguHEhEDbsmSIy4t4dAUJFlru7Xu9foRmvsVEPp6ZeQ+Ya
Kakk8AQEzJBpCPCKrUb2I1FNEHMOrXR6h5z/59dSon1z1tuh0m6NqVP8d8C2
URbOt0Mm6NARHtIH2wmXL0gvKHCXNz+cCXsL727rMB/mB/2lvEqz+2egYabJ
fIkDQ5+Ib9Pk1QRtGt2GAzr6axqB6+qIizryo0lmY/4vkxYhV5Mi0Wb5Pfgp
fE24+Mk3yeDx6fI72bJwhKh6F9TJyQ5saNybZ5VYJrh1cnkKONvJH6Dt00V4
KhpEXNfCDruwZ9GxD+9VOVPRRXtlpdlArLZL4kUoe0LKQ0N4pCQ9hsjd2/um
/f/zX1bjggM3FtT2dUvs2o7a/irk22N6E8Cb+S9Rd1bchHnK6dUQTKV0QCgS
WZtdwwz1tw1dnso9Hi4lDweLnx4n9a5t1qfu6ClUqb/reU7szRF7Voy/iBjO
qy1rRwP3n2jG0RP73y9btW2xV3ACqDYJuzgSSZeB9CAvYCIu5GDtUvp46N/K
sEC5OH52qsVIvC+a0X+YCHIaIZnsbx0qiBq8ElaAddEIECHJ2RSIKwSp+6rL
sQky5sdpq9FFvMO+keX7QsNK7srAgLROnVPDDGYRzKHEQ2tz0tDy+AsNKiRO
+KvR3tiZFu7GfZ2ZdnE5IgrJq1wW1oo1Kw2mzpF2sCQL7PlLSuky91n/yNtR
5HAwHhwmCZBGdWN3Mjw4xTJU/nq7IyJlLsTrVhVza0i+GnzmX1T+0D+GYzis
eLlPy+z/XqfGsdVrSpW+zEUIP1757BLKWg64XDevz8Ri2xZPKbdgra4E6QIX
hGM/gwnwRwbJzdCWmjRJ0u5JgrKuO3dxqDv5AheHyxnzROXh+eLbuq6Cfaqf
SOokLJG8aospMF/fkHenOnec7D0anG1Idsc9gxlm+V16fP1daSR86VC/2Rcp
PaEMqQvsN0SDmBgnB3be9Gl0cDzeFo8xe93gNQO7GXhdffoOaHbEjoM5ozar
O3ncTLs4vEl49NhtJXvMIM4XFiAxft6FVucKpPP5gWGGgoH6XpXJCWyczvDZ
6QwZ7EEnH6pRUp8nf2Z3aG/xMM78Cgqo+AZqMbqlEuETWx2xIm/KW8PzISXc
KIZbAOtwH5pdPYei7NMqiT9MGVcbcPPcTuLdLeuXKjsfuF4hz8O51aEnu0zW
7oxZvXmW4aEuIr1Suw5a5Wn+j9HUWzew1UcIATEIljmnKfVOm2AmnJEUfTG3
aXmVuBgkSfygOwxF3K2mA1snfVXyTtBNqyqKk56tOjOKqasyEM+iHLr+WT12
0FlSvMglRWB9NWjHlkO5J5GFYee5Jb2vjn1FWiwkQWYx41xvHUjMCs6WU5lT
+pHve+t2GvtNDUYc4+Ldnl51+8d4JSRfUCQE7HXZKd752P7CN+t/rmYdihuh
FBIS/vjkW6fiWbKhv1c51KEMxhtwGNC78siNPy/Mhd6evw4N9HNUSYp5JjUY
wOWpe9iLT2npcbxhcKoe0w0WkcwGUZ++jRfGnPfdmGNZ8+kPtBKfMJDtgxra
usEHe9HFGQzV2N9nljOHW9JDFdTq3PahDsivq7CkAbzunmG8o5w7ucZAmC+W
YpFOFxhmy1i1BcCmhOHCkwb50SdK158MCGHHyi/ZRY4JTboakXoMtJKNil71
UAVfcLRJBc7isesNXXVP4LP8/S8El5XskxGIdaEk3KCnsKpCXcpEaNWr4dl/
HPJMZ8/Q9SgTaBU3A+sR6qffVe/t3OJ0ESRH08yYpVW2tHPAjPSqmL04FXFN
cNF3LKJqVjJ0nSS5qZWskFq3/56Cf3BC3t3lq0Rk1S0SyqOjkXol619x0Jyf
WLNfDVHXmPoSWx/WxcG7FG7QCMWTFmai29IBNBfpejw9RZVXt8c12uYWIPyq
cQv0xrk5B8jOfuFMAVRjMh7a8P1pzdIeCVR8/3f6FObZbH7Yw0ImuUkWNVh4
5osoc2Eqmca+Ahx3YeYToyAYXipis03bMhioMQDYhe6n1I6ZJufnPa9lfusE
4wNM0+Yatj7OS5m5NbTMkh+xIQ29SQ7eX/lj8HUuxhIFrG6TX8JniC8dUUZS
iooP4quwvngYtc1I3IJMLy1VkI6UN4/ToTb2E6BlIZawVSYyLVaMA1t8Swbu
YydbVIHX19OVwAujMh5wcs7z96JXncvY2gn+nStb1SOvoaFOpzlQJx3pN31C
521HD08h96lIkjStcl+vSHotBS6sm8mGoyj89LOjez6UfWKhiyeO9Iv5Km3P
zyFa/f1cfgoDa8+B1CY8ZtIzEDGwMPpgyFW5+cCrvA25cffTyRvEf9hXyQi/
ngruHQK5PWKoTg5zQMzSOVSlAi4y3hq3x88Ndx25BLcrZazHKNVuReWA6T3h
kdkfOnuZ+v2AoThrMGpsz6nxDNG6qyqXoQ5SBIfDJDJHb0bUQFkBR4Rlm9Rk
jhEHtvlxBgOOHfkuiUZziy3L2OOfhYyv0gyl0J/CW4Ao3TMQBqmQYGV+LzlY
Xrue9V6FLPLeIqdID600kaSMuPWyvo1VTN9zXmB4IONRvYzT7LUVCNAiKVq1
CU6tjY31y9FkVBIiRre4rv4Pl8gbeUdYAUtLiMxxVq/lSi1Gp/4UhCwjRIWL
a63RSBkqJ9Yj4nDI3Ej9F8sVS2hA+zEJ1GqJPy3PK/pRrFyKZ8BRg83fLMBE
7fSr6CSQD+W2h2dRA0Qnir2tIrlO4MetXVEyb0ynG8WdrEGm3RBeaW5jbcFW
1BTZGWg6NAYD2rZgszOQ8jJgPQScEPlkAp16LK6si4ERclAA59UnK/WjpF0/
4oRkWMbD5haAiiYvY3+2zc7ZN+AcqIx0tFmxepm7lZnucfazsS1U1rfpWj5y
9IxaekVGL4m7RoTrrohxaiCJk4nDtzVT2c8xMAYCevi+w4dzwM3hWToJvKxl
IqbmvVuCd8neVdQhlrNoTDzVamVqTGJZZSNusgcrWkju1iicnfvI+YgI05am
cwjNs6ca5sdVnQV4m1/cAWNK11lsOiO6G4LJZ28rRqmiXPAdAtNvut6tHUFZ
nBKLlHjloBnsfapRFR8Lq6jtqdNlHX4jJrDzhfTr0zTs4bL6b7ZYPPpXNDeE
W3GCBGBoAEOi+B5OMTAG/JK9d+n1p0/KEgpLr4EjZSe+HO0sVWDcglEAUZiN
ro3zn06+IvEnR1tnfRCBqiEnrqQuJ/oMxqdE34MWYtuP7xYhsl4+6zFLq4bW
WhIMiw93FxBU9uYUL0UP5fKu1PvtwjvywobYIN9ewzKBZtc6zVmtvjDZ0DyG
oYyMffrxzIbCIr2IEzlPqATCVf538O4xIclkTZJDjg7Sd8vvHgatKWZp3dzJ
Hv1ffudx3dHrJ7Plkh/Xz8Ug3ej2IKL8x675FJIN1xSuQJqReLfTn/2gDtQp
Cm5fvl+coQ4n7AKLXHl85mv6uiOpVkbql3D4PubIzt8wqoH+meS+B4edHOTn
MQDJwY4r56ELq+PXJ1EL13KnSI2botipd+Shrmxl5mup1oZ03cTYUc40dXvL
6VB3JcMJkSnkogRkvHzxHMEJO0giKsscn/EhRNeM3gafG+G1Ola+YN1CE4+H
MNUBQeIjeNF+4R9n/MKxXCpkW8UNeKCw1oPxwxQtRwrVVHxBo9mRk8axz/Tx
MarPlRHcwOc6/Ht+0gUrhJwr3TWhwAIB4bEMb6X3KCIIK5I5P0wjTh+W4mAh
k4AiIpqC8JRocwGY8INtFfo80hQry9cJlLb1fwgrV2Jz8kabu6CKBR5zmPd4
/bKUTWylSwNDDaYS0kgXbeVD8liJnXZGM5i5PLmSmVfMQLnNYreZ5BYPsSCU
Dk8wv9Cd9ACxTjx2oEUgrW2/6OwLruGYNfavFk15Ikh4+S8stlwQmqh7xLTz
hyPq3mMMBjzh6GQTwWuQ2l3exwrwEy7jcxATWkHBxBJHEXvKmhVwk0AuJ5PX
Guvy/YoK/yT7QNRiS3vVXLPe0uMBEL+SoDMAm1jWlfGoLwYNbhxVeO6ZkDk9
6p6R0YwQQQ+phtBndwXQ4eZyJTN7g3C5EcJNS8kHIQE/hvJaiUOpUikzCo3m
8jGyt+BL7K/YnNn1dkCuTwnpvp5yqXri3/1Z3VKG6USZ8rl30JOJhGXv8oTA
jiskFA705BtGv0D6uGQG9Eg/uzjwDEKmXXBDJOHCNKbqAKxol+4ynk6D8JFB
7dnakoRDkRE6H2WzqVyFHN+wbGiWKULL6snYzZQdR4ecnVamfKGFSSm1Z+Pf
LCtGOUOXf+fNrupP8RyVZQE366gPRUnaCCvUmlhvbyVSgNKPeaS8T9NgZ5Gh
49z59IvryxL/DwAvA8+kuFTZye5UdUO8dSYqeEUvBka0SOrRr2rIuZGa+n0r
6NndbMubqZZPbPkAxr8IjkgikTXx+ivfqX/Xxe7yj8TjEaWTT9ZEwQ/VttHB
zJruK4jLrtfNLbV4HDKMD520DXfDt/o6hs/1bOPmS4B3Uq1zwgJy6VVycvEt
etegMTHL13obUgGdqfYz3kDMRfWJKi3TuWw47cIWVTe1KTAWuQ7UyhBjn5/I
AZgiESznkdNnazW5eMnZ6MvRlSNY1rwWhv3x7wQUxo+6QoIGN0S3tSBDiLJr
G1DuAfcdPOZpwK5yE6C+BaW6wY/uooGfojNs3fZXInQFsJa8ItenlFV2nD5U
IYOlcJQdPpB3OuWBB8soRLGZjOVq55MDk2ZSn/g25/C6b1UokhW3VkVUi4p0
SI562AufzdH7mAFW2iMHoPcWLLPZlOvoR+Zkb68EJtAoe/dnPFmbXaaZB/qQ
A7rUhRH4CpigA8jChHkNaiBf4ImbbJVM0HE94Sgptrj2iRn/ADtyC69aaV96
dXq2MhW9WSZpjKb69VV6yX8bOpLd3poYxSzHNEsOa6QfMVY2uBv8rFO5KYIa
h/C0l4AfviCC4txsOzIRfScH56Mz6Q6KeefgbU5q4LhOk2OY61VxxMXY8zFm
SHm5N3fJreTWFUgflNmjokVCboskGzohX1jgN0jE6eJAbw+odtJf+g3wMLou
Eo0Ar2kkwQAHAzl5h02pvXKjFhTlXXFDINZWZ+tCi8vmjIRUrDy7pWsaH6DD
eVQOmPdtBZBa+RqM/u1HDSGHKv0kaPEMfyFtDO0R9gRgX1xzDVy98IXWEmsP
jBrhoAL1AWFDRqpbn49WtSBl+E/d8m4Jk8KF8H2D3xMAtCSixH5f8wtDHn0g
v1NaWoFMlxTAL0dlXxZm9JQyivTXTXMkHPQuy3sww9ELLEs1s2Sfybch5WY8
Lt75g8N3FKURWyEDBzNYbkD1v5YUvlNlayyG3vNbY6yQNJd2I12C4pioc9//
YGMB8RoKi/b0U0BbP/1Lmg/XSQ87jQSouif9co027jr5iWPVeXrxAiJTd5Yb
cguVDw4FzOp/L1wNUDnk+fW8iz1VbwdXmHFAHOnp/s/J9AWqnfdBtmVUqTh4
WutiHtrMqaRbUJ3cLC9s8uq6US46fj6jIkd7i03i/QCxBzLTqBclkeikbX6H
KhJ1E7Hi2ol7WQjQ+vM00gLAI7SwcLnOPg3LLQqEPF4/gMDatQgwJYZ5Pi0U
Zz+NMu/JC9X4bEIZTh1qwpXuqKzKVQxcr247t6Yy7/SMppwuDxFimDEiHqNK
GP+ecI3IOule66X2CYBwsVPnRG5SY9vJk6i5cQZ/SdE0KtIEoml/uEx4GDVJ
NjNszRz13Ox12G1LAgWeqemiSjyk3gM1VmNSOpMDe+lCPIAz4n5qwXFJ8wgo
SXKF3CjKPvmxcE4uRQ3hHm8+boK0BCwXpmI3XBwMGpq1vHPuqpWwW++5foQY
5d+z1LYpaJce1WIvg3qLaP30MpeFhDGovz+aMrhtXf6on+RCefY7bsv1hdM2
cvoGPlyPrwKCerAzoZV//oolm48K/A6vLueAXHg5sPq4U+A1+vuQEhL5zvPa
N7KKZGQVWQGTdYobpqWNTMq3Fb2Zy7xX7j9wVyveuqfhW0dc2w+8hmJa4mpg
TJUCFn9yqWGdX1CxUwyJ85lqGHEHXokH4nvakJ+3LZ80J23gEgF/HpZgR8AA
x68LhJra6FivMvL0iiOlnijVPPSm9HqK/1b8yBTKqNElJvBSnHR3WcDNf4Z6
YLK3Bn/JWWTQyUjBNuYrBXF6peN93uOP3VC8RO0M2Hre2OoqJuiKMb6WHr7H
tH6bVMTsRqiekb9hO4OZuyYfp7fh0wEwjA/HpjGUps1yzvzxeuopVisyAWTS
BIe2bJQWowkPCn3FymOEZO0cMW1np4XGjspdCeFXWKzsPYajpE3mizvZ7etO
RocCUXwZUlU4Ix9fIf/uPfvokkRrtVlrJoTUu2cerOVmnpmmD+kHo/9KacPU
r2k34mwZPGP1FeLA8+WaOM/6Eu7uhF/WQmSnv51t8jnPWFno5gPQNppvurws
8MkRl4d8NbC2fZgiSTnsspeSNpFIC4Bb4M5H8ugVlWRriIqYC2HDR8dq/9k6
Jp9eJtXIQzf49UXqyXNQLaGdzD6Zl7fcY94Mk8PFESDnbw3FrsejQA5p5hgB
QAwf8cR2q9PS5U1jJyrcrWTg8tL0LMailZFyCWFV6kE098wFK6uhFYb7Qw+Q
a8LZWXEWgAtG/6UvbzJBo881mpCF/VGSAT7UzmhU3ToqA2aY36VtHpb9BAef
agMWVIv8iDAmbFjysxtbmReGbgTxtt6pYP0NdNDlvDU9RpyhyPkaylfCfb6W
uyC/nttilcGHiV3gGw1njxTS90EwxDF+WYJdhe8TzLcA2ZjT/iazFiXD3G6I
CZJI3L0ywwcGi4b3tVApXpZOsPXYbF/5GLRuszMzz3AZVqflkI5QeGdqKGgV
T8YPIem0+JT+9OhnGgWWuNKkMxB0zoq2Q7aVoCtIUfjEVkdO+3QY9gZnuiYN
G96SXD5qm71h0ZgMlmU2f0Lk4dQ4fgGeWDu2VDK1Rs6D057NrIetUvyNnyHy
oJxNUto/UvvH8pzp8xUNzY0qM/np7AIEf029LqmLqm0BcbItiYTipKoHeBBx
ET4atSXzGADV2lGsn6NiVK4QvlUoXLgEjPeBqdlgJcUh90ny2CotO9lPNtsQ
Rb/lcmdTVcveJWg6cSfY7QOqJzbFam95f1janprlbgoBcXocf2Y4bFh2euym
rp1jRqczD9+5W09B9XHCWYMUUeKgu6o0aPTs0SNF9IEOR9FQ9DTwQ8ozCCMM
KLtV8afveJ4DSUjT7ug/6oXPoEqpS2/vVT6Po4GNhqLz4M3UQFldESWUpYr7
6dYEb3D2XZsYAL72hqNF58qn3bb2/Aa2rfTRTowlPE9ubUGJGx3y5dc4UAOR
SstdFoZ8cU+/LprReMcAeef3SLLly49aYsYFRNa/oNPLSf2jXqrSw9sVENbW
kuyttHWneqiJ8ve3TY+xnbEAcd2xoS+Puf8f5dEtw7yg+Gg1Nd9aEIqKX/bq
R6JJAeSgz6TmotkbNe9IBEEbfPdJZcRninERr6PBel6MTD0YhQQjnEZE+uEC
KWSNRhspYWFrRtU2EnupVhPzF4G8NKzqSIi16oElf8UPxb0u39u05HkPCy1e
wzWKTnVbsYg+MBBSyxfLD77KUa4fLFWFfXbk66Jjk6OqewU3Xu6AGnClvhRB
ITeNTpQGRAwRE1m9CbP2yKYBOtc/jM0rCz9ohocttGGRjuewyf+CYI5Gt+ZP
hLK/S+B4nd3R/Yqp0Yau/jnW3SkWme8cTJo4g5xfQTU+5UT5orb7XrXCv7gu
swdco4wfXtVLa/JxnmPEsak4ducnpC9o/iAvtrPUqJE7J5Bpxixt4uM9pxzW
ulmrJivWjXahNhy4JLlwmEibAODeT7rasPMRQYtJDJlHjKqEJDdASLXaGRPw
osuWBm7RgK3/2zS8XzmGvMrLLwxniv6mYR0fuyF9pynSZDAsSsU68KIhuADs
ttYZSceOyUX8/bGlIBUXjmYriIh2tC3AUc8jbVeDUnJgvPTwcGv2Vp+Lsyyx
6v+jUqZptjxzdtYehGPsISgh5T2W84z0h0mZolmgEXMKrI7QkzWrAos1GlDt
ibwblqi2B7Kz47uJT90z97HCQWa2lotv5sjPNkfqnwfOfz43TjRnASaVDOTX
01A0Z7q6UT1ewnePty5iwl7Ocy3XQ0kapM9vjNF6sGtDNTBSqjI/t+m5ZHYC
yuzdNus1u/yK3axlguLFm8f6y7Bn1olR5fxx6c/ZxxP8CLjwTk4a6MyErTB9
iPwrtgUG96dtFF+lubxv7/BvWiUDEUmEovjX22WigPF/vEYxZLlFBRyzOWpr
rwdiDSxMGt+Og8OuBbYvh5J2t9s1eScaoKTyotgI7GviUYzE2nNXo06iBzhP
Rwu/FNo/4xLtbTCSRpWMRxc8kFIdypiJoqoyerzK9Y1WY4skhaBfrWkUlEt8
0Nr11XRVaJo/RdN8CJfEtcVm+q9BSZU7vKDmdrWtRNcsAC2U4M++U7HJIC8P
TYODwtleiVYoTx/2MtT4vYM3WApgbx0L+sc6OlWY6rjcJwVqTyPTeHBCC5vu
xCuBzMEVYncFbCE3D7crAz7f6AxqQrR9sH3pWJBxjwf61/nNKzpchI5bS5wn
fQCWLwgXoi3zk+70vQuzxNH88STKf+np3cTvMDiboVe5uCCOexGdqN0ZdO2R
Vsc4b9M8NL5dfHUQGo0c3Nbhguxof8+OvJrq+KG9YEUm29DR0oXTo0X0wjeg
jlX0YPOIs0E069GuTgrZDiuxU11PMHVgH0oSPLU6FBJ63RbC45BDQRtR8qru
qCvsFzdaz+csaqxZppnnoP0zYCEo0P0OVEjodISXv9OsNPg2zqmVpsA+mPUv
OzV5JHbh0ABjJJ/pnzEIaNkVX7UFEBijeuZp9GZjBcr20K9anNKhZfp5X/oM
YkzBIJ0ady/RsE9mDO6SBVMTdLQq8X1pddh8bujNO+jZ+7m63cShYdrRqFTP
fP8wzkiM0bhGbJGWLT1WjM/xIbVZcL9DuPC7kYUbBJX8vrTkocl7ln/FYmJ4
V4nyJD0D5nXjb+rbMxg1SIU0IM+aDxz93Xhu1NJtR4kAf1J8jYBDIsdwfB75
npj6dlrTugqClvBWTR//L7nA66eZVbFWdno5uV/j/Cr8mZTA/N+/YYmv22GS
SUeS5+Pao0AONgIYO5faz8/Um+s1wvmmECk4A6COl0VANeCc1GbPqn+OpITm
Du2dblZZodmPQwdVRxWvCCXUQ/hlo4fF6TVeJT7G2X3w3QbY3T788KaJpCoU
aeWmC5FaSR9HdSJWBcpARkcy6mP2BsrIjcfW2zRzmdRAYKnmox4gZ6uZ1b7H
tkjo5IFesvUGmp5Sx47KkH9+y7E0NSUyjFFx/Dl3uRLD6EpGcE9dxaE2Iaev
nbEyY+qXK/hRDKQIQnBz6IDhTsacaTsoYGF/UO4Pq3lz3WI2qGlHbqABqUmg
YL0ZhFO8VobgbNQ/CT7dyf7AaNSMZ4tmy6lLNR2isZZsIWsNVwdEUvT7cwT3
mpk+5AaF3qucQ3Tg5bO2y2UxJitfHGgTla/KDPvO9fjMljEZJ7dJkE7kmg5r
FUxFbhQqclGi3UqNgVUTYuIMg2ayekYAgdbCzeZUUNiseNsC8Njsb9AOUOfo
A/dIB6+kS0RZG9LmLdleJNFc94VnGnnht4uEc3eG+ELd6pp0andcd1a09+9i
7OTDB0XqhQAabvEDkL7wOcM/GL1igeeXX5KpydkX/K+rtKa8zRR9H49deSxb
gGcLMNpFhVYmJcVS0Ovem4m+guxK/AQzI67axZvZs5KLqSVVhkOrr7veNDfO
4Wa1agusBWMWqiydqWbcRhevXcV9Pm9YPpKQR5q3dFc9DWZUVZeFUUNjQNrk
igUVsu2ofquc3Rfgmk5km0PIsFATWtmJOS2VXpcbGZta4Hwgw6vmqaH3OaAV
eECCXpgFTXMpWcHPf69BBIkR7zCHAgTVSEAgSNjMt3p3sPkwfAPMnYgNJc5l
DmW3QVbwjp625gx30mqd3vPYshBvT+9OD9FVFiFV1KcJPS+S28coWR+R3LUo
nVSRa2X5pCY6ZSn9d7tAcZSP2KKc28ZBWce0OqCr0O3TPUmo6W5WEiyD6KIo
G+MFc5LhkS4A4jGTa8ChouHLh+mHc+5/VmBM62rOlKrLxS6BaX1eAB+/CTpk
xr2M6Pv2phjOLPGR22nc6bfI5XLX22hFp8ECnVpmhxoNY23eMtJMsG6YuLig
Nq7EbOMwzYoFsIm20Cx4l6ofApWM8o6rB2+jhA8U+g5oeDwYU24Ocs/FTdqK
FUetAfLIBfqEq9nBJ6JB9nUXiUdJ+ECCmgte7uVWZj9zvfNdZzqPf/FsUmaT
n6P6+2p/0peCArvkastF3Oaw7T/OtxQWVNepe1zEzlNocZIsHl4afNqh15K9
2b9gp/BG43aWHcAXxL3bstCW5wBTkH/Toeb/hQjPjNAKdlCv3T9WVewPPLaY
+6wHD17lDI4jX5TfKLrsc9141B0zEufZL2Ek7FTadrG5USId032i4aTJlrAH
UmT+DIf4z8xzQ28bm5vDnWVNki3SfZ/ntf5CntQ/qF4mUdZ1UBxiD4T3EvNF
6C3l8Sc5bdbYAkYjnQ0a8iu/tiBJqbPKQ+uf0PRLQv8geUaRcu6tiTvGIxyB
CgHAGXO2aWzn/4GBhIhbvBg70BzQXpzojUVHid3tYsKFLZDlCFWC7yFkfDvc
TuZ/nWT4MLLi0oXFfcqrzo6k8mjrX3LcSb5Fc4/WMIXLczT/LKSMViZp1YLD
OwRwneBlL4c92yvicqWAME1heNR5Ot8ZmuIXnK0oc8v8D0UMOFBJ2BqSzMar
d6cOkTwKpCokO3Uh6YD7VeLIIyZIbjZypl7Ys3Jo53QqBmt2d4K7iicRhbaQ
E5Bv1gU9nxRfqsX/6Pttee2AGHE2PQOPPChZjeaDYI+eCWHftxpWmwC8DmAW
UwP+li7BiWhPntHIS6uHZXh9b9wao/Ox9pQwGELze8gNQ+38VH/isxEEgYgT
WlR44gV5FYq7YA5USvbPtOjlxulJEyS+2yjf9nm0Y2e9O/peDdJ29fqGq/Rd
R6rslbOgHuAtXyK6KuBs48TcYPcr5lfgo9lhzPlIktgQLHx5EZq5CSsVqw1A
B1hKa7GHd6u/lt4kZGHXHxVIqGbEQDSwJd3VI10NSXDesytb7HyijkXdo3vo
9XY9HlypPu+d2p4hH7Jj3fdRJtKxWzaFJ6zj4gAK6YHnRa8FEB5AnsXOoxXn
RC5WuO8SYuBspLG1B55eLAGS8kFFw55fsAK/yezAlGbI1EeYhLn4gCUAZahs
Aqx7HyuuhYxeXBOCU4YlcIkeYPaj0IQuerUTk7G+0dD0TbYQS3aistBGNFV9
Aws0IpTr26sNCNvsyeNlmCOJzKFT/7tIbXThQ3+Ldxx+PhAT01GvUw3uxPjO
4eE6K/WLC4tZ7OIj9jYHzXKVPjAPNj+RTF+CeA7mCDZWka8Df4kumvMJJhQm
c8CbxkzVdwrIdOua3IMbhIeGGFbitoKVQ49T9dU3BAI6Ld65u0ScQgMXuGEH
N8GF5khJN6mEZ0fmxigUtBJdcFXaO6f/RScrbbaoDbY8uhmRDdWrhSUk1lmp
LFgaUxX37Mmb4SjfXQtA0d8C4b/I2va1pXGOgcNph2gLLCs7I+DtlVRlkIGF
QJp2myC+G4AW3aIzJBu0pi7/iPGKTQYF5vT759IDDfqRkgAXOAFs5+0Q9aMl
shEF0bTK7qonAgAfKbNqQzJL6xRaMr9KJ2cYS6Dt1P38Q043BpVIU80Ow7ev
wlzYu1ZUaA3WpkKlffZ47Dq7X33ZSjEnibm7sEBbqv7NbQQFuS+uViSqXwuT
0BhahpECAOiXg0bmQrRAFyzrbwY3B9NU7+kGEYf5ExKpJVLB8BUWqV2MG6D8
eT3DW/EQd+LR62yuFWn9FuON0Jf7wMp545fhgniXSzwBbU/dciByqNkN+XiL
nCtYmiFAsMVSjM2tlO6j+mPTkjouLqvDmYaUtXfefxuQB3Bxrnw7NO9oWI7U
s4PdBYRv9Az3uj6ycC21jythLLO/j2VsbfSLCRNqDMt3DbccLQrJJegaODp8
C/uiZ7FcMvUv3cjoo9uFc3XSIb/Ti841tf0SX4kVxPUzkUJY3oXifuWGhR8p
6bpbowd+wbNtuCsVlHT4icmuBwkF6Wzg60MWVHBAVmWa3xvh6zcNmOJm1zDW
s7bTln6fSsEJcTALaqqx8KVL/xvYaBLN6oT4A/1RIY0rOHcTVpIAtI5/UFOL
iW7PEA/B2RYjyyDcEDxR1dvwHng+Y8HpwFAVDuzLJlWiqYRiXSIn0T6av9cW
97L21xL0Ttlo87HnUVrsEGTX+N/rmhTCY9mL2ew5tvCDnHSvlnBc07HaTtfJ
gT2HbmFAxfEXiG4EMQ/ofbx17Y5jc+nLF+hJOxzPTyhUCJZTHOXsSqn5jyQ/
kuZqsN1702O0VEYBcRV2LNf0o1gUNRh4ONObebck8Wk8quUOJAN35MrDqIyX
MZPaSKppFxz+cHzPObhoHeKvoWb72BiIilK1lphEyIjGwYe5JJGr5GLximzP
34UlOIlFjzqSOcJwygJO/KWCNyRS//DNF1URKcO74V5BC6BE0ly/PXPzev8b
cKZ0mn/11KeoWBchS7++bYVSGyTwis8gwOE6LphBebdK+kS2RVDzs0ut8x1r
p1SwLfsGcFdDkvOi0g3M+Us8ehUySHeeBrocD4PJquHoFuCMy3JKucMjA4ZQ
qvpnGhR3PLcxAdToLzc+H3XuT3GG1oKZxR2YV/qW1WALAisw9ykqhhwO4cIx
kP0YR6cSdoFPvuObZD2hP5nTNHgsJWOER8v8055wbLAybDx6H/XbMV5lITKv
E1RJ1xVLCuAfKFmYOOvMebxsltQIN52A8F9lGA04zPJGiGNajgxosUwiWrNh
QMpPq+WSPhO+9MJcPHgci8NBBcKHAejuix7kdKP6RQq5pF7tbnp3f1aa5+Ox
LPofckhlaXxUvUF3+oMgmXD8aZGloBh/NugedB584gIxodLMgpTNvTFnUHpI
nVZpEnz4OinKH8vhzu3Tr0TYuQMDAjgcg1LCXOeXbY/vTt71Vr6tjOur79EM
lYkas/QdMS3xe5JtvXjWOPJ7wnbLqspUgeSEwdwRp8Cl2jy5PKWZ77cXW2Gk
ANszT9JQTlRWBMdKeEA4H85bLiDaw9o2VDMMNghHsTyyRuCELqOOsMGsQ16L
uSjjUf7+VhsTf8T/VhUGNyCCEUZFsDWsbzfCz40ysRWOCWyMpu37+M8hAal5
9UtJ/LB1ckp3mMnjqqz5udvRM5KPS2M2MUCLca5QFOTvBPU1yJm6vY7gDEue
s5hbr4u8zeChlzrGTYPy6l5uG79rH4CwXIp/ftU4LjDZgY9JdvwNZke01/WO
nzTitPQTGrXA8DvoYMYoHHcItPiH6N9bYi4x92WGBn0VyeWewwgX4swKOG2T
NPtr5PCiRmN4V+TyGrg3ZUTgzHKB+NQqoof/qrE/EQKynsD3hSA1t6I6LwGA
2+Zp/mkhzuJBuWu68hlGgOwRq66YeKHGtJW1FgiDt9VuzFPQqH90iadgX0QJ
c2eSgTl6Qaa8Wg5cCAT7gj+uT4u+s/wPKDL8dtpl/VMaYMsvFnAQe+U4jc9A
aFdETjyAUQNfc62PA2YYq3OlkDe6HGHJp2RMjHXuynpjAZjjyBU+ChfWFCEO
FwX1wDJQ2ZmPm58dyKltJUCQKjeiPl2kZssdfKpyPMMvoVshUraIGzD4h8Vc
KnOC50JEYREksv9CCvfns8G+pCxjvelow4PdcY6ipBUTjSVRx0ju6BWOzS74
gx++u7PYHQjzbdb2MgJO16Vl63EXCr2hp/xpyvZ/niuWMg2W3u+ReDeJoUGi
cQXw9xvjOFkr4C8/KerJ81CVD68DhNoJF/rK39OijS7FmCMeFyslXOVLQ6ZM
11IILS//G+UIkRdD81xEJe97aM8xBwI0/zhZKlNBfXSHXHLKWMBWUwehoSYt
/nQHA7qkNlx+RBv7lJJn/zS7MffJTRMnxSoNTZy2w2khgq2lwQbPI4dmstks
3NBrADRZFgkGG8ItQYDLh+4/9R+aDYHeK7VmiuopuRzcs9uoh7MK7F4RcQ14
MEZUSATi+Zuc1+6i6PcXzMAVPPSgMCJbQJIC8x9mpXNxBx1tPsBRy7WLee1A
fGPr2CCxkor4ceB9nGeWQ+qETjKg0bo8O6+CvZULs7OMeMaQ0L5bzBl3jEzZ
pMVD1ohMVMjWaC4YaebFVhZ8F6/OGW9lOP6J1nC+kDP+llg4cCC+p8V3Dz5C
USlOWQuEM9jmfXx5zbv1mYGfmuKSVbkDmYUCPCpNWwkznC6keH7xf/UEJp0c
th1WIpKjtePCRImGej2T6rVZ2+38V2n2uHFDBzx0t2labIdtcYUf9tGGqmnb
Dkf8d73djQb2O+gwla9VcQqn/PgGYEJ271Cx7/xRWNEb/GxxZf0LRw6254Hc
XNYpBdsktyCOxkhxKJrDZe29OvPsKFztEkumbaEAtYoDvSC34fmR4Te76Yvz
82KLE0PlSrlAmq5sZ9iJYaFT7Yzth+bIBKRkAkckwf+w55BZ/GzulFmCYjJE
eZWm2IkPxzMk+rigjfEvUGiT/j5hssq+2gcKTLxoVAibICJk1uc+vfOmABFs
W+LMRryQriS4DBiDt5hVPKvL3b2PGulQ0hOpVV1DOUgCt53ukVDB4zj88K2/
mAPzsQ3k9nzQ0SWxUjbtZ1VP34h9b0DxQovBSkYYqKYWO0tU8aMV8auw7J3n
QbqXMkDpwpmEU4VHSP1N7i4AAFVL9BKangjj6tVBm24zo07y9oKP2sW/jEvK
K+1by/YFjNnS1vb6wJIo4zxwimlyUrv14246YWJcgjAOs1kctE11Dd1XrQlS
cPUAzilsTPkkC1/YV/MFud1SoXIfZkanTESyE74hT8S9oi7VdIYAYknWfGhm
KCUBmGhfsbwqjRyCTvZMFAL22cVvJQ897JjNAytq9MYaeDnicHVJVdYJalHV
IYQWLR9K8dzyv6qPeN0pq9ss5CgC1rku2z0vWX8AOR5LHJywZbTfZagcABsI
NH796i+cN7dXDu/bMCA8K2llvJZjNtt8TG3h5W8uspxUMqx4hJorUuWNxe+6
J3xXVMYhYYXhVeTQq3JgdEwUEq9QhD9LcK00V7MxsLCa5fzmbc/v10JQLROO
GvwBjaxcIgVq8cwqRIe0kGS3O9lUK6vq1J36AP6UHdUPCFrtqlOU5Edj/pCV
FXgIiuGdVCS6nlyBakO5mUk/fh0kx4XTMb4gWPPbQsWWtE4kWfg2bEpx3BXe
pNXucBtaqXW+lthEqwhR0KYr8PoBdmx8yLO8gZKJaOhpAWDa8VUGwfbHyLkC
wS4igazYpGgKROrYohd+dCrd0lfbWAe/kEUR+d++gjfeqSVQoOkJfyQFZBh1
vvJgIcetn5ecmAs6zVFW3Nx1Lra1TQh212s93C8U2vdJS5orjITmENwqoBxH
3eYldPV2JgKYKj/Ilv2eHE3wX8C5MCkyaOrxZzT7NtXHLgI+ztv47D9kcFe2
ME6GCQW6J0HONnpMyWNulPUEW+D04aNj7p1dX66OvRDxH5csPm59703JIpsP
fu8xpLqHgn1id0WgUyn42ALPsQWt/d7Wfx38lf0Rma+8zGOKDPcaCVsSHukQ
5vtPnXtonEGNMDAQ14ulIcw1z/IDt4qqTDFeiKqBgI1pcIA/VtUqmOGftag3
sU55ZA4hf1x5/3h+kdXXHMr6ZTNzlzS9JNL8OA/GWB0reTzi2mi249cvX4cV
/6pz3xVKsZ9xNbPyVCU9ubIw6S7L4GNKLF2vPS4Pv52kepcnX+pCuNBVTFh/
N5wmRSssy8061rSvUwiNP4i80oMILnzW0iMTvphaktq8OirmosoRPX0l6Tt6
HPMIDbel2tHkUvTDGd4Y380Hdt65522n9mpoNv9Z47nvVSFCdtbv8jJoG5O5
+TOcJvVrVk+7nYcS4VilDQqEPpjT4qLage/gwAPa3MIdWPo+gchcIhUVQ40M
LvbgyVHrvu3Eo8ntIKN5AjyM9wyuZvlSs99MxAq6e4TllbkAh/5wtciB0M/2
TfE6k3v5rdt9SU5yzTuOznr37Eqp+/o+ie36mN8WJ7TG6ery3aLTl/EZH09l
EGqR94UK0YgW8GPz17VHhagMIk+jDXdDIuCyPZtMFQoeRitfhLoJ/tRiYaWH
Q4BStrQYd/SgPYJsWBiyjVrH3QI7WepOr2buxdFuGrJYyGWEnNaEWxtK/zGn
BKdDf5W1lyHq4npAdPTcWWf97BHIpTe/+cmTBLJSOZz50AAM7ltKxZwHqP8v
FWyWDkZvW9dOBNF0hteqi5FIcILrbVuEbiI4R2EX/yvMWB77Qn5qmAxP0Xsv
nUFXHU+5z0xuh+BDdiy0Fy32OqeiLpdaGM5Dnma+xIGWPf7bpW+vMolwHKMu
/pDM0MQh/YLpGvr4KW4jbiYpdrutOB9/Roo9PcyBCrOBgudgYI3CviOHBtjs
3NuftyGoxFBcZYVCaqimfUepxjiA6P3eQ3vOvh+8CKaVih7uC1GhSFSjsps9
vSOFQRoJZs4dgWqNzQg+cnQszR2jEmkcknnSIpod5bD8aBOO57D/gCrQFH66
jm96vjxAV2ZOmK9bAgcMXOBwsXM92sfUT1Wv4D74PuO8WdOjtZbF1kl6zmCM
6HXCAzdZcfkQ3A7aw12wJfb/piQcl43jduG6nl/9cqsN/XmJtWoRh7/pex04
l6PS9mPX4wJpDAUQ66a2RrWSo1CH7LAMm/dU1qiShHIquyj63skdVvUu0XB3
O3LU1meXd3av5DIRxpl8Kh6wWxCzjAmzAmARX9mJEmZS8dzK+pZ3jDTAqiSQ
FBo/cFHA+xd8yTEc2UuFs14totj++I5RnIo/HHuEKhOKRjX+tMJ8pH8bpgkY
E9M7r9RXeBAgBIoCUxMIqAPN18a5hkUjAXcW4g6WwPtdd242rUCgM3IKKyGs
zxwNGSf3RMLKwxLEA4zvDbQ/od145Wzii+rsDkdR9QabegfRxpvdwmB3sG1H
VoBKWEWfEthW1OnD/lSaBNyAtl2V32enYWPKxNfcVXi94hh1HagyhAj1BcCM
9m/YSK3Y/mJW0Zzv3nL7FPOSoVD6WGgLgl1gzVBE9cKB43S600ztxCib4TMi
X7+m6hWUUOBwM7TW1PK2Y/28SCQCs1kqKkIqzt8uFd4eNZoUka4ZOJOVv84H
Stk0Z7GrHunq0MFMZ7yO0LAPccgcRR6RhPd3Mo6JC2fy4kuQxi/n0No1zzff
MK4GmUD4FkD067wx41firjrEwAsgZaBU4F9loUoqsPyzc7GjnfHOpmKMXhg1
X/LTm8ja2F9B+hFUIzTzwAz4Q56HMmef8sd6GdTjDV8g1lt9ho4xAay/+Fn7
9o9jO1zrfvR6FngkkvNfItGarBb2A7fYn84WyUmTlo8KxRVzox3+XsMkrTOD
ym80MtTjlOn22Z9jQC72Tj0QnhWrkY57vs9J0xE9ruBXiZ1UNasePAEONUQz
cmw1p0OZns5rNICR6AGGvNttCxfoXUl/oS6XHBrsuKpUp/xas3fMFweun1Rw
zXvPS9AvLVhivHMhUBDdqCDAuB6lpGZe10xoTxXLhHdXBtMwmsinaFYxgDs/
msEWs+NtOWEDa0M8t6Bd3lckWzmGan6kS1e5knJfL/mvhOLjrbYD9nGy/E7E
Bn+KyRnmY7hpGOt4qN3579RXY6P468nV4SZJl4IuoXnAbklkN6ur0sS6IZMe
4JUt5HixMVN8PHh8SCt8YkrmiY5eK99b2LitpiWro7DKwZAv9fqdf1nMPVFy
3WXpKhiCxiJSixpGha9VRdKpBXu0vBS6bUMJ19wPYzCc+1My+nnWPFqR5qLR
32GC13M7DzTVXFGDuQIQuoETP/MSVqxPpGCDjA+/9c6JWODN09BgmTaUtBSj
wv7uRzBwlLWIKM1AJ8D8KPyZscz9B492siViylwn6oyTZBk9grUtenarCL3R
lk/kdUD0ugRRhpWCle2v0td9rchwMFkATSIkNRFwzQu38nTbIhB/7xIYW8ES
xN6UNh0tV5LGi+f/66J3TKvJweDMBvtGSPPvfr2uO4kOoUBeWzUcWzDchEKl
cxl9dMYU2xCkol8P6kx5Uzq3K9UaqIot7ml/NdMPYUmM/Hd5dQzUzZS01fi3
ooYF6ftAOhGtdZXZSRFERZHNiAB6TTJu7x+WunLfI+GNFoPdSM1+94TbiP76
2g8H+ezOHEFAfcsnufPM8vUSDUN825ceEWwTQGwYEmhKNLNCOwWa7RBIQmjh
rJga+wYQe5ZAHZ3FD2wFN8jofMKzpJpw8SeFvChTFovrDeKuYY0hR5BTB5Ko
M90snNBh9mnXx9mJ+ANGv2ZxI6DlFW+SVOWFQ7JXVt8iWWa2ldz+ROVt82sK
BfuQq9KTKSHvTtAGnC5DEImrADF/hQ7rJsfNTG+MrUm4bTu5RSRVY/Mj9ZQ0
zXmQRHb3aj6zLmzIOmKZiV3eS9V7fl8FYm4Vyy0rGyutGBbH8/8v6y6WUwd2
Yb8MABB2ybDPfZZOK6DDyeXeXWd/jxsjGPrpPb8CP8k8BnjMx4ZwT7K+9Teq
JgyBiPKKE136IKOlDQiaTHOa6SWZny263/SS97aUqVyKwxyuVBUGMTVlELAX
5Icv01bhipIU7WYnLuL4NpxhCq8uUmdsSKHSh8xR/fcv2pLPfqT/2hzf/3Au
cEM9O5pcVlY3bGCYNnwe4kQ0rRzzRJuQL52bLsjYNmx1GHw7JWeRZrUEr8Lk
3CjCXTn+odTR1xk7uxej5ovXiHtt92mMZQ7LWkv2Mvrl7prLbn1SuTUlk8iJ
TKQOe2Bt6WMCgwkaIyGnL/jjIUjLw1ehizvX/OHkK2mmUt4DKdCXYfX4lA1V
+Qcq1GIA+zk3xsSIf1ihLdyyf2RbYYuhODBCWIvv+DK7oTAEDRAG84DuYOL9
USHTUqPo6oS0z7BXvXYnMJYiQG+4oTZ72P/HGPd50ScWyshr4iHu7U/2lXgS
0LFIb3HcyBF+U26xB+C0DRyp8aXkoRtMsd5AQVKhnlGSTqMS5imjI9LTcN0n
gJkH4qEpY+HLn51gna0J0jZPVdBYHfaghHcYm9G73xLB+AKdw5WMMEIWqcw9
y/X9TzNNwdOgPTZG70jrRBRjsXHRyl3AUGFBRu9QvQ6DVxsvmu1Km2rWQDML
nP+QIOBrkya3la5IBdSDGWVWi9ZGXe4zOTwRO2VCd5QFG3zakVUHqUOVeLK6
5XV1ys5H8QVll9zMSF9jJzeYPSPQ75rqcvZPVAIYpc77qOcVYjCSE8XuIO1S
o2h5fS1+Eb6Op3ZNXP3yk48HyJxxR7U1Tyi59Nzl9K4cFOcz1RCkf3b49ZLW
kVsc3aeFc5HvZfclfZprLbYsNO0wuD9lxeAm6Z5Mna4uBm+F+ofNLhVgtqg6
CntivgGD3zfQahOq9uJ6CNswSz4wPgyi3BPQ2I+3FFPoJIKozNPNBLW8ieZp
ePwYjo/ZzqilLBn1f1+ETZFGihPfJ8sD9XCcNp8JUCSClnN28pAum14riRzH
CsFe23C6CgLxF0iEtR/bzsg0jp3/L6AIpKUN2VpJKbhzMLQSGKhYVPGjlDWs
h5DQCv4oA3KR706JiLonHwy1GYFx8LeTxoIF7WdF74V2HjKCQq+el6lK4Y9U
e3hWGX9hXJ2wktRx8OLfsN2xGnJvwhYS1MLsO8Fz1Lk7wfAhQ8zCXdtzfUdo
qF91qaXPY734rh7C1p4DVJ3MDPN/rxEAnpT2bGJ9+yexWQUqxsvy+yPWc8R6
F7Tx9ILEZy6UWcGX1IV2rT/S0gGfHNAzrzSpICg/MPk2cozaXvujn6qneXib
V0ZVjfGwkC9EuP1uexNjkg4Cm/fHEXG/GZtFg7UwL7Ss29zHzraKSCQfv6gx
upUCMo/fz1b2O5S3QhQfO1zxrmI6/IaId22vCjQ5asBoU+8+D6BGnosCXF2o
oHMW8mAX2N4iGVjcwmBnJc8/uO1dgNtpWi//sTdaPHeJ5EJfPPgkRw1U1cMq
XU7u+n0yYjFudPPJz0Roux9AsUlNfeE2415YEsNifH+4rilJ4szKjrDiF+O3
DiudxVRk75TwYhKu38AXXSzhnAq7ZAg/tIdlSxsHZjGGddxv2x4fSQdfndeq
42YRea+QRJ3gE6vaQvKTwrHWceH5QvkJM3aUzsZmF554N4fz5aROzWy9fT0r
tXKrli2B4yscLghTAbka6MxhQuVaVf/rPlcC8d9/wW5JvPSeFzLLUp5qpcaF
JwukAoV4yecggGxcfY6AUZ3ukzWURHJ29EHnAsTOveaj5MokVRtbT2+mf6lY
Cr66a31Y2TTEIqNJpZeh6udubHtX8jMtyVI0Srbzs4q+ZOs0YJ8l0iU1mPj7
R6ChCSbIbTMeBMcS+aU9MdcQ4anzV2kTq/9fDNGD1Qd6l1JLIdrEOiiRYnax
pm7ivEboAwe5J0rcQfwbeDm6MN5OmqWZnRZ4GJOP0mbPJ96FC5K6L0HvsTlQ
ZYuiMVZWssmM/+HG0zwhhKIyANwlVaaXbXPQbpxkh6XZoaq5pGNnxrnpJNrd
sE/2d3OmG7rXzKPawz24QN4rGZ8sPDtU2EnIJt4HDSHLzSLo705vovssNVjQ
Q52cVK6gGT6UM+Q16ZQ77UBRiKNe76cwZHnOrFSv0wEEnSrSsX8JI1gPPy2q
Y94oB27CCG3CftJcB6Z494dTzKXQ4HlFpyhEhYQv8mCVro7enyeBRbtIn2LD
zrzdOyVftMzT87GdeH8HPKSQdo1rXcHN4LROvZEn8qCwoeck56/4luDAJynb
inV35g2JdZ3bh21NkIhKQEVs3xxc6H6K/letjbGNU5Am4Kd9nSJoouKxynkO
Df3zGvJuuc2LqEUCFGxuSPWimWQvSs6+Zeh6tfYKSW7U7MMnCG6raUcUim7y
CLBeHX/it3xOSbeYoBQdZfHmFhknUKew/RrsAKJ/fWddDQgN0JO97iWgVSCY
kZAtd0j8YSnfio9HGl/ZUL8EGF3QmpdjvZrsekRevM4QNkK/JmlD9R/5hfVs
Vf3yNUTOuYII0e0hi1NxB/aZ9FoPgEAgdPLYP9nNNvgVyJXhuh95wPQWOHvK
1S8zWUBf4tM3oo8Dk/mneivNsJRaFYpt3h98fxLAEsGgaFo442n71o/629qe
yc36a6BK5JlGwm96aVTAd2bWG+4X98tC6o5DvbAOorn1GNQbcDxUZgJX6ORf
/naYgJLW+oga8CsZ860Y+VrIWg2IGHmIaH57mYCYFiqUGENZDaSpv+ipHmyk
L5JnHoA/+3x/BPGuxcK7/nh5q0WDXqdoA/UDnbWcDavN67Z0fBHimVY9Ksr9
La4AhMrHczp8OaBOKPQaKYA9Nx3wzJoGVGVwS4Rrw8n0a2pBW1sr7OcxQIWQ
E0BvXiI+L8TVykmsysL3OtUFwJS7NnrdRafppqr9a99mDkxsXR6GCEJ2JJpS
T0JjusYLYghNoeyoYzt9RQ90vmczSjv7ZJ7zJMzSSw5f236p59L8YIqBInnW
do8uxsuHls/qOwZbnbtIFNZZNIGyUbeUtLtAAwV/6x1kzYxfqcsuzSaz9ZIY
WAFgw4kg2/Ri7X9GPyLktcoDHns8gSY0Cw1HQXwzZ+IlB+5WQsOA36x7Q3qG
lcjO7ElPFUAXqzBeCc0rVUgmFdVHFRzkuaBVUs3IKxW2lgh2p2s7+SM9zp1W
NnJl/cCssAtV6KEeSkkiNtjDyrIftPNT13Iw1KuwMh2Go/7txRj7sXBLd9sx
SRPNcBJ+LilK7mkfVqtyg4PqDfKA5ogJkKLQmcnpU1JxoCXPsdE0HR4lQxeZ
GZf0Tps7zhW6FDdfvlMhZojwQEfgdYzL/muAX+f90xrIBHXrzYXy8kyLatut
JfTOiVLmFbq89OfwRprDNnHPMTdolvEsJqAM5kWvkDanW6n4LYPpNcnPOtsC
KYccraeu8td6V3V0JbJKwiyAyraPtsyO5k3HqQ3WzRDsx5zWafXhWpoXYG91
+/afqQ8lR8THn3fu9HxJ0oepJGjTEWNM8wk9RnkascCe7IVNM3iFLgW/9Mj9
Cm4DeivN86Ro88lCR5PGVcocOBXGlsvl4oiTUdWWWhYe9x/1MeXf5/v4cGpO
VOCo3heIrdiLMsEDPCEg/JGLozAd8lGpqt5Brm3SaMGEZ2HEE4XPYf7H/MIC
1hBDX/NiEJ/FOUEy+R4A5pJ0UR4QZ/KL259qc+nDdSBNhZKu36PDTLjjjEHF
Y46Lj7EgmGL7HTF8T5tXZe3fhfnWJ551hn2SWVt8I83AqoyM8aS1EnRQf4PF
ytb8Q1SMDPjKBSkYUwc7/fgIPvmf7CXPkVV3KkWTeGmSqt0/7xSlstfMEZAs
kr5jyIxC8WmWAwdKddRczmsSQwh7u8ZXGaB0Fv87oV9mHwm2Edl0fuAECX+H
a8yndXB0jy+I4DYBBkpba7C4oOVOyfbZNLh+oPoCQyTGoHh7H+SGz1f6sKtN
DLcl/hPghmp2rpHJcRFmmFswuSAmrnUYEZ1LzeuE9XzV/jD91hCYRVR76yk/
ik9mwmQS4xp2Ali7x95KkbvXJO3jyRNSNOLBZVJLOi6pSjI/q6pf0+4KiWjh
XfO/PlxjcFz+g3x3BtD0hRNG/QAxc18HCPwq9oo1gXOxX/k2BMiWX2jfYYWe
YWw6S8elkm4J2NbEejfWz1K+lHki3gd75Jmm7upagLeynYuZUkFol3l5MQGy
nHJQXbjl8FN7+MkjTOB+9Snb9HP3oodISoY6oMS8/ERKKog0/tybN0atBvij
mhm7d3HzfHdzgQR9CBTVpZbH1/S20jcxG15XByCNLrly1s/RhdeBYY3q9PV+
vlMPj/jLfcZZsvbpVb/Qf4sd3DiBf5v0d1ASuvVODWkuPXMAhp7olmShckJ9
sYDAFJFnfvUTlEfZfRobyO5f3HEMUQ05jJtYSqJHvhWl2YkmJUXpl03DECuI
pfwtqVDoNofh2UB5Vem7FKI+K8QG58dkFnFF2RKp/y735UEVqm8HBXfmozg/
RBs0uGv1AV9TeZh4/E8xVTJSox9fspNk3azywEmBP8b65w9GlDNpXsw/Zj8N
hijHNVk1gNgXN65lsoURfmHJKavPQdvdVnDW5sQI3dmMZiIcWF8bOPzA+wde
tq3jnf5vmyNHRnFbg7GoaUi5fP5LyU83X8jKABiZrFUdpEWG0iESS8taYE6U
3SVaxcDkTQMZpWWDa2nRC6Nr2ivzWRepvAdLu8+e4TQ8nIZWD8bRduG9WW4f
FClFanaiVAnPHq9F459bzK//+G/DYSORiNcbYo5jnBf/otcHmJZ4Z75OBFel
XSYOBuL+AZ8hJQ+D5FDuamwT2D+1twViDcRu8gOwvzvybq/lQ10/zByL5HUu
OaL2dL/Ut3ekc/8yTu5bobR4cwk9RnhPJqJ7KNkSkzXsnNTDKouTCAyBD/Sk
wqHsjTCDxW2i7CBdc0qCIxtGjKeQAwSjXG+EhuFQAnmCdC0ApL9ApmBoLlgJ
jpmQA1kP1Dy1yz6ZMyBfsP7QHxYb/4TzqEfWi2AQDUfCpY/gXgGL17ThDXVc
cwPfqdt/+zLyJGffi9Qn5/c3ulOwov5IpKPm8+QEaIeM8RS/Xffn4cfu9wNo
74gp6o02qq0ooIlUZTfkwTAtnPo9emdruDG51hR6BQq5ujrOFiCN4o7BZFgC
ZbUY+U7dYiEqgKkB2E2G1ezhMTddh37wg1L1KcVzQF3P8cSoiYmwFxlaCdo/
4z2qRYX7uhDkaV2/YxoT8kKksK1a2uSBRgk7/3EKkxtQrlRfbxUE7DJAU8UR
G+Ft9vpFCJzMfzFj/rndylSX2csZiwSUmQFMFCn2jbEQcgWqpRqyNTxMcnWB
Q5/7KErk7V3PPK37jbQV+vuj7VGzBwjQvXj0Aji0POAoYycxF6j7WZN3kb8T
D0FX/2E5fvsSuU3qXCFUmZXKbjC9MpcFCvOzEXGuowELrOhBT7TFpph3iD9N
2yELV9LXK3cPbmC1yFgOPxXk79FDDkRxJsIkBfufMgkDb+6V8MT1J5T4XXj3
Lm44BLL/+29ETCVdR+rFfZ5486bJNebUO5LCYlKaZ/KDpJRzODZf0RO4L4Dl
XhXZCfyHMa9ezM1mk9tlbzdIMXpAnmpoHIUbfJNyUH8bTwG0ZmnCYKc6ZdML
IbABZxtYrxon1ky8NWRCos+9qkayvd4loaQhIiuXgPROttty9tjXo2KWTjpg
6vipOTRDKz2h7Umf3rb2EkiIfSuCKmqJIfLavs9s0FGYYjomEUIXfuSah7KO
qY/YP5zTdn/NNwZJRtg9YzpLrRYj2MraVRWMdtaSEwxxdW80jdp3R/mCmqHD
J2EwwzJuyJ8r8qwLkw4IyGP/6fNEw16v00bY9NrGKJgUObsW1ZmLX9FYkfrK
eOtXngOZo0jP7wMO6iEOyeId5d+cRBNPXTI20EmnsdqgrjVpko5kwWDXz4QZ
vW5PXej5tROic4Ora/Msr1ezmiRa7IP+3pg/qCY7MHrPZVmnd3H8q10SrLzI
3XHcUnfSJGF7rcPbpHqwUt+LTqVdoMSeRKnb3v70cQLM0INesJlgKRNhDD25
/pezyr30SSUAReWlzg/dYbwvAaOoYRWVEoxndv8yJh3LB8Morv7pGDYy6T/W
8IqiLOzJ0UPrNNMq9ThxnVLTVXNg5zVX5yDo6F0NHDlA9gZqZ/y1R9i7rOoD
wEOWnjC4aubnZJv23fVyTRkMUrMaHMrVeD3jOn/egeVXJgBs4RfJC23yUC15
ksVqIu6qJVNf9GDxEybd7ZkOvuyG6Hdc/gQ1Z2WWmVRBKaCFSrEnQK4Fwf7T
Jb14UEgIJcb0jKqjvud+6Z9BVkbgECjs3XKw9hCapuCOMQlblRYAEUNigalD
rseyi+U5ziGbykkWOi2tWf/lHAZ3d4kv2n/TqqapSWAxd+qfxCCwUudU7Wot
e0W985cP5ghP922DvB1hjoIxhlzPHJA9k341aoZ1LXnm7joHiSY+ImsND3r7
UNWurrjSdmFicDNncZbG5RwtV3LjzcA/4xgUr6se3n7bxKTr232qrapAwyFO
redkgP5v/XrhynJBUdrwF2tv9Brtr1bodMvQdHJlc9lieAiCwpHhTVnwxHIh
xqZrePdNUO+WWUsWi+nrYvzkwFY6VNDwk/ypMblcoXKqHx2XiCm+2QSYtmgN
PQVqpXAOiyr3ZksHdM1BA7lYU+AyTETyHpgsULJUiHloJ1J5v9XspBcADDh3
mwxqCZhKt+kKchbpJn6kW6Ye7/ccTV9Bi7303CrQYJodvlfxq8hsMm1cFr4k
LnwVlRitJE4qWF6AG+w9bUBO3pwXgL1lzd8FFBQpKSyk0aOZ5hvwbnZaaRBG
l/VVkApATK4oHA/DQoOMsAHdpPxk8PpdVXTQVghapyvLvoC4wcq7EmH+r3E4
Dy7hKZ4Olc79ktRVA6Ff6BV/zUgjP3RRN+FPbf0/TLm8tDrR7u0QkqRcUqMG
20bcH7a6Mpzh91Jk+9A7vpZi6sNh2UbAs001TgYfzouQmpeErVMwD5LOftjo
Wne7sKkacXBW0ykNzRk2O2Eo9ARmgGLxKyzsEf9264BVOfmeoZfb2PStBUCA
JhgbBICCRoQ6u+IJRtsnQ21VftYBuUt/FvjhmYYpP10BlqzCh/i9bwKZ2ZDZ
ZWUOvta1KIBaDcbpG82hQ3nvLLYBb0lQ7oxdC0tIYSvuz2OToLgNLNcXKqCj
v7Ul4bDogSipaaHJTd6BJHqCieleKu2JspmHCs5RWEnJRAaFbP/rorulG+KN
hl9ZRN23r4CVujb5RsOKL1pE6//ZnJ/GjIQB9UODvZ1vuBkHWEHCvrquNhoE
2Qc1fQZmGcMSJpom3sgvkM7UFjzIxUB9H9Rgsi4GPPtGqlWMgvST7cIjobCU
lR14Ms6qVa3dDAOD98ty7H+xoSDXLDDVvsmmdvRnLWDDQgXdSpKqAWQ8Qq/7
iVYathQ4zXaXZC3fDzhyPbtkVcQYw0In08aHQUHDZKxhEpdH3oRrKlYD2/CP
9KMIB0P5hpBqfi1feJSHGvUGDTo5FuASlATGqC/GbU39NX5Irr2uvbV1Tgro
RIV7XlnVPrk5Erex3fcXsGaKifqk1m7Rd1ispH3SKP/VyVhVl2uqN5ef2izN
mBO9UUdCgOq7pCzwmZzNPOPosjaFuI4EUs+cRmJBa5H3DSvp1ts3iAnINwKT
h+rrSicvY/66JI+Z0QXn+6vIHofGlJsrUMFV1X2t/Yuw10Y9KPYzyGceyTFL
0fUDBxGMs8nXWgg0AhZmdk12IDemA0Cm81regy1t01LwED5joGMWupZ8uz5a
4KrB6Ehhe3trgyUe4SRIanSEyUOhD98jrwflJ9IPeiDRos1UKSi8fgdEuJdy
N06XyZZ4JYheWkh738a7YKsHIIl9mdOeAY3lct4dAmV1ojdg7i92NaWdOtce
LDQO7uHL0sKk/ML6OIGyLNVHN/e3V5HDfFcZwE2JxaP9dXRKlV1KOITR7/Ra
9MR2QRJ4m3vP9nRwCjS2i9I3FaHNsiqrKymch28MxIj7+JZkWPF9hRxauw24
4PSdsR6jsv1/lnDY85ICVp4JnJBkScZ6GPFp96YX3HKiRUG6BnSVI9IKfY9W
qJUXnVqsApVGvsiqKNmmM8NdNG65YLn/x/7IVmovKWWM9ehdnyzHJVw2J4dV
pf5Utqp/oFJc5XisW0TZ7R+7ASm9NNLjSleUr5lZeCgHxnhVeBNGZT8OUuhY
wsSs5DxidKSbMVJPQadZuS+qN754FNvitBlVE/Nr112Qwi1D8Xws4ztYuZ9/
0bnD1jZ+sRzz29t1r0J7KnYkKrymW1+DpoV7rG7S+1IVJRLXlmiP7s3WfeBx
xzgMfslL7pMigi/V6nCbRw1uXKo/Uhqfs8NRAErUf47YFeHpdXbzRmZCh7//
9NQogmDdsN64ChT00BWrPgh4taqt+fpZMiZoqSwvXfnWF1E/gaoioUqlgtkV
0bH1IumCzfndruMUF/Sx8Q8Y3ZHyTWPWphBhVaPnizdbxRfkhP5VJkoCdEMX
QjxatXzuCEbkOZ5emuo6yq8NzKs1OztBvZ7jS/rIjGjbnoTi5vR7bnnzPpIk
GHbgoFKUT/dJaoMK7vvpIDIyLxcARtfHXYRS2QYBBQPD6IDzmN0gZ9Vag2C8
4TFJDgaGn0OW6M8flayMb8nAGG+U83ni27g1k12M55fpnUOGr4HNRIDTg5U0
nVJolP4sYjWh1QQQYyoS8T6b2GY1Es8Mzkvk5aayeGgpGuUrDCsqVq/9WAja
Xxs3AHVIDyhf72agPppCHd4nWiipOqdtuH/asITp8UNeEGgckUjfU7FhWjaB
3tp0kbXpBUqo0XJ0qdMsi/m8xn/YGLH1bYV8A3/orAs/ZbyW6HMdJfy4XG3l
V5HZRKglqq7GmhqckVW6hPbrKtgx4Giz5BGMCKm1LVUeCIRkzgp+qA5kGst6
PaC6/Pl6RuyPymDMlBp6sXyX23CbMrRbggv3M2G7bb8XxCLjKSLqXg7Ui9oK
77G/JLC0AJLwH4Qn16Ts0oghQ+xVFuPwNbXZ0vOOt8JXLQcAPZt3CM+Vp2Jp
uTzF6D9ovMx9kZagqEu/JIjxTGr8M3y1ketWMppB1u8EfHHXrs6dpgmBoC17
OEk7RBqlbHWv8jeXYsF6/OoW1GpPfh9m1UjMjkBaUxKce61YE9TH7LeySIew
FhW4DxP7vi4n0g+HLyfVdzzUPD/gWnc9HI57WeOCMwGoEuFNCHMswbt2jAOg
WV80JsskItVCNV/peVLoLVIAaBpox3K5Wpo84l5+OFcUg8qeCXVF6r5uJH7k
0vFH86vXcbjq6fuHnHuQ3Yk6V/9oFzQVtCMnWUL9lOoM0yFm7QNOgN4LNSIM
G6V77ouPFi3tvhuadDmwKaFZGRIk5+niINAzMUs4fV+4iVXFgi3ICnzUwOSc
cLXdtElvBqEnw51EqLQwB9VrWQfKCrEvbvb7E5il+CW7QM4RtrkunHJnILLU
eEEd2HvNlHVMiS+daS/Dp7rQWud0n3XWmHqertdQT3q0iojUHB74GsQLzcMz
un8FmSsBjeSkMYy6bVcRn7LUuXS73TPAA8LOta4Mr9vFoe0u5R3GvPPlbw5h
saiB+cdvycAZV0JiSz9wCWFX3JUure2VBSL7p2z0vNaiUYZGi95ifd8wjGCy
Cc+9CerQ4EZQsAXLyl3k/q4Q0dkQ86TUx9aBTUreAPXeMD8duBC/ZYFXK6Hi
XiV/zBgTu//5pqWy9xsVxSp+m7a5ow41i99pCYM/FWWLW1lJZoltJI8+6zB8
6x6GoBOvwsDJx8BnvsDb+3M8WyjCrm1Sd8EzWvVQBU/2JS2kGlcham/yCXjx
E03XMLwOnnicvobUSw309lFx/Qxrxc4FCgSrlZn8riwDIqcCLkSSPZ9FHd1X
6CRpBWPXodKX/2gUokx8/N0V5w0PQjh8aR8DqamLtktA/KQpL4vxydCB3MJl
jQZFNYpKCFA9pdRnpFdg4SSSwdWW4yyWN9qw1AyP8jY5FrV+a6rDI7Kg17Bc
FIEeuAGNgyE/nPGYAvfetEHEJY7fUEU8I9aW40ihzuYKcw5acePejfT8tWqc
ZqF7F9GlkodR7MnzBkRuB+ifFtM/arrogrAVsYqXCmAfL7MbZrPlTT6zh6Am
Z1nUJQqfy2VIDlQkQHhK5v9PTohZnJvSanFd7XC7Saww/6akqO5N305xz49x
QMOV5faCBg25NGFsW/vde8/y+I53sZzlO8jzgm0OBLS6RM7i/LltAb2ylUu+
BRaQUiuzvTQqM2Q9cR2HryL4cfGhelVI8gWBwq1SQbQZE0w+R3s1XWzfjl4X
mRPTZDTeroM8G1mjH7rO/d2Tiz8hRcHuxo+d9fR1B4WtaIcPrOM/UJdpdVvr
W5vpERFdBWl+vT8/x2h6EOLJkJhyuYnr/z7A80AJr8paNslvpqSTQeKJRq8R
m3tbeABSNOG04S5E44tTN28EUBzyx3mp6nlaJLm9fecL6k7U2feEGuAPuLUM
/ivwtWaOK6hppRISGN4Ox6rrM/dfCLDoB40GHybmH0G3oPNn/TQ3MLu7ce8M
080OtsQ4uZFrJnkKBARuQR3Rd52pUvlM+L8gLTRtr1PpDDBYN7aa81KUjTc1
2vl1V6SVrJaue4LXZgha9iGo9oWIn08ja6mJSyPuHwBypfZBnggG5lXIyqcD
hUQvBto96ZxGlvkxlgmvJ30DuCOzZRkMgd0spuPCU3G6+ghaYgLIqnUBVU3t
HqPBt6Gh409jo/iQdN3IgEVq4fBUs7k6o1QmWGJlN/rSYSH6TE3EeHyjMjRN
FskKV1fEkBj5Z5NUvyWwhOqmfcoSHyszxjr2zyvLczuQIBxh7AXJaEq/976w
JrYhUYr4lz0+ramfRvco8tdoRBc7VfxJAVV6vdDMRwMPz+jHM2cCUme6apCF
iU7NUzGPt6N/71YC1LatjaDBaiOfLQ/AUOZD2hxl0MpuXKYxajtrsIsikHTv
BhCMTnd27W6Phv//yv7B2nXnAiJ5D5S8SyeSIEzdR995Vdbjl2rvWK3ftqps
1UrEXfFXRAG6CxssH82R6pWKLneQjBg0reLthstGWPa9/tMRaZoNzn9/U84H
tUqrv36dJjigKXEijyBb1bMImhM+iVXCNrxYvZKEj539fpWnu8gnkPvXP2ln
HeZVt9VTr7aKuNX/G9RDd/GjL0N0gN1mKjhAOZmu7rvEQuV8sOHryZO2tWhl
BxRsQ0k8BJitHmSg+faUSTmnASxZW+GzCt9WYk6rPMd+4A1By5iqZJizymTI
xUYx16uwIavgWpHeDSksY16+GS4o9Jq0B+eLEfEAQ9Q9Jny6dDETuQfwgRbq
oA+Gp+2vC9ptl0ncBLnAzIXdhvSrjy2S9UoifsHVdrbAs/Ux0f7zYtdornGC
4Xj5VKhxegjLsVjO8e3ecJ59jNfMXHp1osE8qSWIhfEv3ry1cKy2/msXr087
xWvUefwqu2/Li6jewbAYVr0LDlqAPxT8pvIFvoCVarfPYMnC+kYMC2LE3SR0
ywE2T/is5lwdLdhAqTPVpr3vwSsttgd6LODgGyyPl854idOjVCbMRIVQfGuU
vvq7b9RCKJUZW49xTx/zNces5H7twxDnB8ev2xb6t2BbjrwF5YrZsE68DqE4
zw3fXqiU5zpN7lKPJ+Kc+58TaDIFefLhEGmI+TdzWG0YoCXvUhz+5JRUbP7F
D40dyVJRx4cFXj0Mp/HvwS5emEjICLCvoDL/O6Q4idDuulMZ3+rFUkVWAZeM
uJ+r2v0f+PeW7S2sz2kPYMwwi/Pr11kwXLNVkzplB+HM9AacCWHzpqvsr1ZL
zkLWTh9l3VWxZjQQila2axonVWvV0h75fVCTMBulz0NGc6pxcMIKKC22iYYl
zOLOBovuS1o46qPeIdWI/fdbbb2T7+GY5ZZoXRV24BcWP1BfEE5lX7z8C37B
toiU21E4phU7ep1I9iw6TTZV04kKR2jq83Uw0aLloX31/S66mnZ67fNHpUT1
3C7OwCNxkzerjDWjYBt4u7L1aVOFJzlcTlQC3gMvntBOWH/glb0wlpP9oaPO
ArCZjC/cTulXVZET9EMbSK8UlyMWUyeBK47MSgFG52BPUZ4V9EWWT9KKuHfM
pERROJ4CVRC49lKnKpATUEuouW7p9kZBgi++kaPa27GxvbpSYvEE3wlXgeie
3sw43ALuIlb6W+CFbVgkiXGVvp0Jooqj8R7FYPISfF+Y7mYtwlJYvER1HELt
t50pxoEXeSZrMdcvjoirQ7WF65f7HTMCXUtcWyIgMhyxLYyWy7KomSCGRzMr
uSyL8YpI2ByfpnxbyRoKKxtFiXAweHkC0LCkF8hPGTwuAF6DCyxLEuv+Tnji
KXnpxPi+TiamwYyI7Ic4YYYzz90iNLW2CpY/2chPeatDz2JzQWJAcIKyfovc
qHlBVWVyaYtC7mpO3apAv44VHKYnvbFwpA/+gZ1/eBAjy+lAMVd0RoTHxybe
sFqXCuJR2gztt2IeLM3zjbHoL5hgYyODxrZ1me7+3rQUvu3ElEMBvh5Hk11w
HZYHlLFW4Abd44/ZZgax7n3CaPxuOCa7fCFrLemln3RkdJk77JvycQNi5ypW
TT0iqGJP8NyVrIMmHdc30k0GdP0IcT9GZbfAvpMBlqhGB9Lg759EVL0W422r
oFDPyE17QOaDeK18y2eXvr+km/xW/cEUye2qm32P2VZ2PsMsUik5n9mqZAmc
FUJAbLOIPAtntnLkr9yjuxmyq82XcfVbR4DffisxbWA0Ob4Ccj3t7CSaa6BI
JCk+nX0YudCxLLsgSK3EUcgvnnZq3TOoSJouSbncy3FPqr0fvksu95fiePv4
BMOb3CHpgrW5uI41QjzPYZvhiDp+IpnAewORuwrtvJ+iml8P86JaEf8TCDXh
i55RrjG1rqHFfpCUd0/W3lcs+JKyp5SiRm47l//cUhFjEE/51IbefhejjyUU
tIhKzo65Vt9XArT0wOLmySnn9D3v6VHfaqr9QcHWpv0IBsUKJSiL1B3goTMa
drxEhPI5IC48O0pmSElnJXfABbDX68O5hgdfrrBzoy+t02EZS/ifgRMQ+7eq
tE31XL3OqVAggkDe2iKD4STaimZcQ6XlZ5vpYYHvxTTpo0UFY7DpFuvs87+G
lJpjXiuYnlOGa+Z6jZJkyR/dMd4oOcsnrtfOWiN3wX2hMA+90AgCICgFPzd2
fhFqQ0f7bSsCuKX2EweBFYOXKHLpb4DegUh8WLgAHcUQITdxWkRnx7wuge0O
tV320hwJBfrnjcR/s/3rB6HyZGw/VSWIcVfmpeB+o/vk2yqWaUcXXBcQuAm5
u/7yVGseeFlamTJ6Zn4NIZwuEp7AbuJSFNWWl+us5GVgTw7o9VNybPcJbbSu
dxpIIAzRYpwujVPeIeIkTNITt0DfU0v/1VV7O9siAbmoZqTeVSjy9N3eERr2
tjUyfldqbfDqdkkJXwI2CYRGgiuezKkLcsTE2YXp2xRlVgWQkAf/rZAh0JEg
ZqyXIJtzH8ddNzpr3G8izZkRTl4sl+uM18EvsY3dSJkYM5L3mSwxZjkCl/xB
E1pOKsLGcvontWDxHP2Roie1uoSg6Qg+5QUsXVVURI1UG/kQg37SrhB2P23N
Vk2RsJQ5sgSVth2gJGwdXWyJqaSGA6ROpOXS7hAvt5eu6sRCyjev9MZmoRwY
KriHjhEddGBm7PpGfbo7A6EVVgGNeL1fW8TliiuaUc5/16aTPDMgfMH1kbF2
ZAD8ll5vUuGc/+HBAWuL/qvwOUGu1ZJItFxw7tpE5Xa6ewECn0jmF5EiCWkO
pDUCjxl/3zxFk5nd4nzwMSsb3OI1viORlg4/3yAEpSaNN1Pim550zYUBL9qn
6LKD23GnJQzVw5YZkY4AyE4686dxmFLDwkIbFhdj+mpU0kS8Zckw22B5XKgM
hr7M/ts9ClCHgOvf9rFWRFAp1xwJqdgbyrrJoKtXCF/p36d8Be4TuNAq6C49
JoQpagQK4+agqPE4Wv08jyTF9QYXibYkjrs9YMB8ZLoOAnq1KMv9H+VTariM
u19FzRck5BPYv1yfdp/8xHA/FQvjI1Jx4Raidc8JOW53D2jK4oFgHgp1+ibD
Xoydtio+X994kQ+AkoR5RT03uAk8TJ4tE8HIpnFcwqXjM6uciiGc3sHrgxEC
0d4eH9NZiRKy76Iv4+13uWSEsMUejR1uycQnTe0I1nU28mkKsaDe/0Aa5XdH
nG3/xlgChxJysZgSvhSXZg+AfefuR/WHoYg/tul7ZjHR58d9gtJNNNOrtX+0
zX7lwbesttVXCKwRj08TFOugBAk9OXJyBgwgSv+iumVO7GUlvkDWBn95UbRz
nQj0gvNQeTWZFt+02ihlJIiMtLap+9pAjWAyBjYXqao20Eh6cL2rq78ZGGGS
JCGwY5LkAHRjLDhIGPDlnsFFdl121DWcCv+ahO476EReZ3/SgmLS3eqtSkEF
GXa7hiBiTbK2pMuPXQ6siVj+6mZ6NXf9A2dL9UgBGH2OdZxzaz2eeHDnkFGn
56Tx3tM+MayNUQWKDAMAzkbFJlscFgX9sFb+I10Z/Ax0WdThSmaBpAaFH9K9
nlikfjqd62aK+5Fl7bo1OMXEc579Obi2Fcgz4eYEw4ioVkP3rixpeLrU5jMw
s4iJMyhyezw2hIlY8NJW7U9WZDsTn0DnFAQmcaUFH8/qUWGlbRd9lVZOJkAP
VJmfm5L42kMOs8maD3YuRgmBzArGXLQdTyoHdttWMtOGm2SU8RcAyv9HBVZD
AuM+k3G8oHa3FXqSD4yxfBTWpDQdJrcdl4ULmo5u1CyvpNxnd1O2HLiJdIa4
s8HVtU3cqAx6l0aeJ883QwEXXIQRIwTi6CxBIB0SUGtihO3bHlqgGVDwSSbv
lKcYnFYuf3gKHDu+qK9+EbYl9A6h97VzunlJUn9lTH7FaKiahpWktZwawpqH
NVda665NJ3nF4bqGXPhhXZ0Gf02tnHVfkrZdK0spwi8qd99+XO4nDkt0KE3+
u9eePGFm4Cq+YmMW1xt0tveXeZ1NIaxIV+uRSd/RQc8OlglH1EiwOSYQ4cFb
Ocguzbq+wBI8yXw2+PQI/3lrY6d5cG9IkxIuw7P/OjvSeK8enXsWCFs9MF7B
yzdIytl1BLr2xDC5p+iTKUlfzc6ciTJIcrCHo4zteFBolXSj6uZ26rg2AWtg
YVYzgh8Lb9KftooXG1t5XuEL5nEGA5FC9ibyXsivyOM19V8oK6yChQvm6V3W
T8GE/GSF17NGNmHwbRsBHpuHzDJB5fJ0qBll1S9Jm1APZzCN0gtSz7jQlFvt
syhx2dqq1EnFP4Bi3UgcSh1ZTePoLocYgjuuPfIgHcddIAnsv7J62AKu2tnz
Sx7kZbZWrCF6TOctUhzlUFAzpoJIqrmxiswtrshENjEnk2KBYTmDKcXWV90b
tzEIF629YFye2M8c+9kwThctXW8gOEI3DOc2nR41UTuEnH0CVxoKaEmgR5RL
uhWcEE8/cYijUOqc5Dk7k0lDjVGkCJvpccuTLOLG6lazBzcko5aoFZmQo+et
EEwA4umu9d3R10P4Phdnh/oR7yl9yJcVcaiUzN21Kq9iYG/pnRqqWKAGkwNX
esHOzCtYD9p1+IQrw7g3ezX5B0QROfT4hlkjOPCzYk5Mflr9rBCvNofoo7Nf
GqgxUVDmujtkONsUJ0F/pAh/G8YK9/dw2JNcmYYuvnjfgM00rPOpabR5vNey
8s5VJeMMnSC48lEZ8IwvuWvrNXvppieR0jM7+BQZxN5jWAwuEUDVsZsQQL06
yX4h6bhirZvQ+KcJBcwbmgoQOoRpCp5ZTQdpnJ3juokbfyk+45H/uvSdLugl
8TAuKemq3dgke+6zXAvDz9pStEhuQQfPSh6202A5/iffXL5gPzzZWaata7e7
GUXdLGbvitReiJsWKkQ0mj729zDBANjOTuOMfK4jNhNKPyRVwJ+qa+8Jozq3
L5n63WwSR1BF8tlPS5fGjl1Bm73oBTFee3nwFSW6YIUz+JzLE0Xz3oselzx9
9trYXa3m1g6wFbE/H5dGk2DDtGAp845vZhGcvFj7dBtNxX/RVmkI6mz9No1t
QENGV/H0gcTDwoFdB1FV0W/gEv1C6WGLLeSKGRmxwPN4TPQXVRX2pdSui0ym
iYNz40NL2wXmLbuE7jQ8e9IhpXnn70hv8nz+tsFMrGh3BUWu15FayU1HJs8/
BZIWX92uqQGzCv/Ryi6PTjsbWxdgyVLIjtIVjORJ2Zic0lUWSQi0XdjdBERV
VIZw/33XI1xUbkj8+O4teLstNNGHai3Tr8j+YFj3ESfiLjXH8miOnrqVgXhU
rkmvGzu4ykVQVyU4lNKuF6uxGLoW7HXtTAScvZjQzJwVJSpENscEhyoLi+LN
1Tm89O2T3tLOfoubjQGTLVPFAbfVqeCOBIZKgZqFBwLDGGFkmsaYg8tgy/On
5h4hbkS/xQXimPL1FCgouosUbITgV91rcUPiqut92QSmJnt03Cv8DxaHTpZ0
WFs0VSiJXmiOI0zejhzDhZNQyKf4jPXZolrapyaQvuhxjQ+JMynvM3eYJiy6
yrvFIFH+suLpad5KyG45+ouyJZI0Ei2Mw8V7DpDeMfUIaj9nXeJ+rgpkYCuA
bTiGLQDiJIisNNj4k1smKw/dRIYluBm/Se71Du8Y274QHAcG2+sHfllJ7Tpm
Esw9AWJPRjLNlpzo6W9b6fnHyPYFLH4B/8u/hFSh1DTmS0z0NV1olY1eiyWc
LF2mhFHBl8E45dj75XkbMHU6hSSR6ZCJPVm/egNs8+wnhTU0vHp1u+ufyb7l
G5PJoQXrHl5IQtd82+cZJRSS98MkoDaV00gHiTEM4HSz61Gcm2cmgPqJ9A2i
y8Y6PqnRE4nQ6S3UU6DWP/1/lf0Q77pUNbv762hjenv24RdffjyBHRM7k/hZ
WhxCNJttXNZ/fgeqm2z44GuAeNVjUK5UaQ7GfRowbod+Yb0iy4Zk6ewByBYX
CTX/xSxqbxcVMpIRvMDSRqjhQPfHAHD4RN/Dfc68muEfsjzSjBKwNyXpOwY1
Wp7beODZpzltObL2aE3Ts2KldsIUDPZQM3fr5DyJ3vigQvgaL1UXENEs4bsT
YpWEoHWPICvnkdycQLBG2E8oKkeLFR/7WlFu3AW82zOqwPCZipipR4uryZ5j
VubiL2yH3ue/DhjIOESZSplZn8J3NQZAGl0MSKFMOMwpGSZ+qPJBlm/idw1c
xt5bJRfolcOVYQ8fUNbnjFpoiQyLnVHGgHNYdAkZ+W8uLuvA/cfioTJ9l0Hy
rwuV91JhtCqGtMx8dEEFnzx27JusjGiZ6QyfBTaSkJW1sYwEt4yCZCinQkO0
HqIX0VJiD3PJ9mNyCW0uvzGHlec1GkuMjlER0aPpddm1ktlrfyMMgLyIwfQB
4WoGMTqbez/FkkbiPb7l3HWvfmBYTYnMqSDHEOyNvN/WSEmzzso5adORpHKd
ZlP7m6ANxtKduzxLW8B652edQdGFA0QTcj26HVZ3c84p+rMBkn2fYyCI9oAH
3JsTSX5A28biB/wbtHlfeXj/bQPyFZ1rVF0pDTaluG4GY3LuzwjL0b0QPD4+
QPVuAd4+baENTrVsj5mB0gHJ6/w35uJi4JX1SDHWA1pAucqlRyHEbRRIz4JQ
qALTZeXLF4eFPYNU7uKzWHeeS5hzx0NxEChfk98gxiKtOfDN3VVWCiHEgrGX
J7qSxnVdLPSQFooNkL00Je07cGIO/+HfexD3id/Rcm27VtuqhDxjVULuJkvO
OHRsCA7H+NdHhiWQDbsPtAoDbvd+fzz7Fewn14M9Ymu1HG6iIqFzryqlt7PU
fo97FwUfZNuLm5d1Xac5xv8/JXTwR41jY8DPRaM0+MAe0GFNMI/mKk0F3IVq
bUpWWfplHR36jrlESuwuKkdXFXJCK2in5I5xW5HWHxWGvxPInPR/D1Qyfzh4
Qng8z6/p2gJzY35i/7BWDMq6LNgECI0zwLyTACGVR+1INM2qWDFHkL+fHMR9
ovybkFXxG8Bw9B2ARD/qndMroJU1C8tAG5Rs/uGTgvAHWjHUYLrZcHywI+1x
eQoL9bsT3F3at/wMRR2TGkL4z7a5HinfhI8Q3MSMwfMl7THPqaB/axrmW78q
CmVIhtSxjQFRVwtUsLctZe+YdF2a8qRqgDpHXMDLO7u87TYuyy5YTfUgLGfh
daaR1yCRuApjJytr3YjQroLdH15QsNWlea26nggHv65T87c3HAUKhqGHoEpz
iw2d03O9PHiMVIp7f45uUbQtL5azihZSLo6JEOaQDqLA43aKxpXfL5d0VikC
HQNrpRQNdI1/Ncijaq9ZKmzTpoKEpf/DttNhcLqV3S1avJD4iHYiJVUql4Ys
AKrUmr0R7LZ19pITzfdNHbF4vSTSMZ58tpX/xdZ3XJz0PBUSl5lQNrRYGMcc
Fkf0UkdsJfpj03nl3AWhX1ZIpO+wjbhdt7M/4QwtDFv4UWwTb6Lh/r1HWenQ
D1XizCj4PUxpA7UmD5X+OSmPs6p0VfKQynC7hPqLzPfPxmwwMtGAcGzHH4Yk
E6dGFoUnY8hhn9FhjnvPUQJSA/FgsiByETGwjViiCfISG8x83Y4Y/6O77EyL
7HkGYKv6DuQQpqq9TeRSS7GoEBD9YXK60r/cmb/HpThzRSzSXcbX9ss2A7Cp
OWE6ARu/cshO0uwar/wG9FMBDW9+TWX3eh1oV2Xz+yLYMRh8Gj+2MpFBq9q9
V0s5X80lByixf2dflDUL5KqkQWq/uv6quh2F022tA60EQBFeik06avumk7+N
WtadJfQY4CkpoOLqRnT9/DyFgzoOc/PQ+cUbkZcGCxMPBVpl+NXBl4vS99s/
krDKBAqcFgnlx5KYW3BjnGmjYRYll8nnRVtgqTszwf+/gY1tDwTW8IomBI9V
5U3QmRisBx9U5zlxArIZkyab+KufYVoFqjhVU3Kw5rJE7TcjnkJqLzF2242X
8LKLEBA8mXrHAek5l6F1KV/cWQpdn3vDg/D+p4QLnhiYoK+QJSDDVYjUFCIT
0f31URvmC1iw7256E35T0GtjGLYlhK4Uxzohi+4bEDXhtPhTiT8TMC0RgSmC
r5LN5cmCbjAyzIUVzvc0cwexYns01C0pwqlHMueRU8F0O1PfC2pGIyWIVyh3
Ms9ZymuX6S4zkUTGp0PQEoTG2Pau+LcNXjCEiD+Zwijb919STNU3Te7CW/fD
53lTLNhGtL9y+SRDhXrWblz9zWPRNu1O71NFUz37vsf41LPzfU0LpqaBXdKX
28XXCk8Vx6VxYM7xBZ1tp8dkmiaBZy8h1q7Trh/hLGZ/eFH3z1J1ZdhPh67r
7F15TV4bPKUWFOqBy3JVKysnwLQvTaFtklKh6vdgBlID7mcdIPlWgsL+Xzw9
hHQ+HkuYY+ASGt3xomkH0Exo3LrZS2z+0vNGW3qnkBKwwcdHwyrmNO66OGeH
qpwU7sPCiFoHaCW7FoMc/p18g8O8YnnFNcoNqmSdFA+U2+HhSiGd/NHMSnAb
zbTAqFUn+ldK+Bw2FOpw97djoYCHuAUlP5bLUC3z8MyJNExJ5OMhWUhethxT
YnsHu5a5lQ7ExKxF7dDZsBP9DqeRg8W+3XwhHnWWzTIsmE7b4w+42n8RXGcw
HX/s/gPsvHhEM88xqnEkxfoE/T7ZnuvXAHcOL0FlhU2QWp++RDyq5txbg5MY
WH2y6RpbZtDZrupShqnzyuE77Efo/FuDPAsjn40F8XOa40YtwTyxb3PiMz2s
ubGVbFopltXTYFo2ij9tH2pQLBn9e/WaUebVtflBlkh0lt8YsCPTdrnEeG1D
WbRIjL/tMHenXE+mRLg266UX5iuYU+y0eWmc3T/LYHbMn3RAvNiZcD+QEB6a
/QLVXJou3N36Aa/mrGCyNAkuLXM+Io0U2TlRoEFpJp0f9BUKo/K5LJsdQ9RK
QYdi22rpM8uAwCRb5Kdh4W3pjpw9og0P1qPe0YHdVkFO75DONZEmEjG3I5+2
t+3xBsRgDp4i4/xte3EVe31F+wPGQ2bj5TiGIrnUD/VmUJZjzHOhMJSvGRx3
Ny1gBvqUpFqCvVvdKMaC4J1RHHPJpYV+mUsjd3R2/RybIWdi54d4ksU01eRp
bbP9Cz6sEtUZCKn89DgLV1Fu6saazX3+xYdZY2jCXi6CUxQVm6hBacl4KmVy
v/PGM4dCJendfrtePCpz7HC/QPtqRTt8e0N3mfmTzooYf0ODSlLnLFcoYmTl
Wf/xGdS5Kp1KFKA3EuQ7R3sMBJMdECQ49jpDtNIBTr+ErJeE94sTKuAOWo6i
CQa8ncpsEl2cKE7HN9rOBGKSQgK6GgXj892iyeMy0W5B6AhygcvTHObkRQdK
3KwXlqAW2jrfISnROJ6L1ClL4k/Wc0ZC2oRASGfi03NXMdwNFMhJImR7RVwV
BVFNTbLZ3DDQmMnPjRDoLB+1ZjLfGdac4bss8Yb8SbYr80BVyNNfYbyFgulk
zLB64NxRO4JqEirEVHfYIKPN2Am8TfDdj3m0P1OZCYkxhx9BxM61PR70a59t
S5XV1SknQzorEwbQq8w2SLzRtdMWQalCuy0xkj/XWZLWwltlrkv0JXT44zZl
YpSTsE+3e6F5x41fGWyzOG2lZOltC97QanyKZadbFjlZ7lNf3fKwdzAMvXXJ
HzVS+x57+GbbfuFhTUP7s71u5Z+RH3mA2eHC3yrOyHjGF8L7KhSSEgPzG3Cx
6trRnJj/BfQSLMCzqBFtXqe+tvRLL3G3EKc9kXyoju05KNkG6pO+UkjhcBkk
r/xPSLbzGdxPfzwG7ebwN327Ee5tTMA1/Ent5kr5leZZOIoVYI/X+IlSQyVy
0fs9Ei1+mOzeMRM+6B5zWU5GJnq1X2xg9SeJWKZIBy7NbbYThRRCmX51oauy
jlP10cibczCM7YbcehiVkO8eaZdcIEObex8tl/0TMs9ZLDiyNPmylAgm6s/k
exR51qxCwOkQ7uSZwinOj6Bw9JZZu6z1MviNk6C8c5e5zilrns3YLYV4TRCq
scRxB33Sv8QJSAi5FKmFq65aWor6oH/prEHf6MmRhhI3+XDz/ZKB3UuG9hMi
keuck0zpgeBfDbntALiX7cbQgS3OEe/EhVEIXkLjWe0KWQZ9ypZlVlxecsGu
zAoU1y07e5j57g0bdARCneDh0cpFeySxCvyBFXfAK5NPe93jbAhpSpJcPntP
gBsRGwY3b3g5N8cQSyK5jgEPzYSYnDI9MDOn1T3IGfF607zgn7DQAoRaT/iE
HpdIbk8Bn5AiQ3ntPE2LYCRGbkSSP4kBP8yFHT23YVgTtfoCuTdYvwK6I+sZ
pb3fdR4zbVkGJLTDqLL/kujEoWL+Ok9zdwO6d3Ml8W9AShZWUKMwqMlSEw2C
lcoov/j8iB8ISPCzutmf+wchqX4piufS3mNbiEzSSyZ5tdxca0IdNBfZN5Vf
OosU87ksaj9gT4OQccS86MS/8447XqFKeJ2hALl2jQ7W/c3AkrkuQXDzuWrf
j6Kx8D8T6Vu/UWILmKZGX8AYUebGKlZAVqPEmhBzl+V95d1S4cSWIWaqfsnN
D2CBBbbpdl5OAkhmHNuqpD7brHSflU8DZWJNy795oEnc9r/mxDBGzkF6c2Mk
dpzwqc5WEs/GqOSi3nUtB1ziQYbjQ24PzVpr0j72U04dtU3GyCS4hrGiDE1Y
mXmMt4YopqI1aYo4+D8R+kZCsonxHJ+Sc9sg4v89ajqtGACd5lQ0JEFBWpMY
asu53jtyDwJzm3bfZmrUIuM8Xm6sOo2vFd0MQpjEY/beVNOMgJCY2xqPH10r
nfbALVnPKrlP6wnYGwPrs1iImjaaA03hfFFbCkqZnMKF09XVt4A+PZX+h+iY
6cbUcFvRfhYRH6vDSnorlGb3+AS9NSMASx2YDn2U87jmFvJ8S6DgTxQcKXgj
uPwfXKw4gUrAklwg8pS52Y5+g8YCKjCwWftDfAx0elm2C02ovN512dwPM5Ru
8448s3iaZWcheeXvxEKQDl1K6HCGc89mQbkbiGV4+gWonMun2/PLSs56keRP
HMMZsBQLtAFrfzT46KpnFGOdie/0peMOkoRRh7T7C8t8MboOrWoTbig8TKn8
oync4HMo0N60e+QKOqZTmOtpdwmGzl32fAvzMshOYmHSpLE5wgz3Anws4sfX
tKlj+NWovAs9UK55XvY7Z+XB55EO1fcDHvjOHR0b6oKuSdH6IhTeeaywZ1vA
5OJ1BrBiZEB4kX19F6OuJUZfdHCnNvoVIS8M7IqMGmxEU1i9sgIW6/i1GNQP
7UHOZp5pybK58igOVmjvoVg3dRQPEm5MiLpjocRyceLJBnnI0MdlhnZDU5N0
VxghvJ7fONvfEm1l3gQZsD0PuHMI2LV0xCMz1/zoOv0S7G6KM8B93rQRW6f1
L3DNjZGsFtpDD5ND+A79qLtJ7BvRTn0oznNvVaP87ouBqdE82CNiuZ4VQP4y
fKEayFFyPRiXuQ+NvnG0cy1V+KcTjIL7Cp/SctpYq47JPrEk96CN2ZIH0O7e
xdHd7DCCaHZukr218em/Rrqcv5AeGBfwd+H4QJDiIDodswCUea8KpYW1OcXi
oTAMJn4dr0FbKNLz44Q0jXHoKlD51KXiKdKmP78/9/aCfUUHrcXoIElK5tAa
Fy16q5BKaNpK5UUzCgZ3eUdnES0AGnRI3um/HytcZANqYcE+++jwrSgvpQ74
afWns07MFoWtrCXZB2PXMH3VjjznbmsnVOFT6Xzysq34YVZRObjr+bc92a4w
ytBEEwl1ohbJu2/OsGqBC5TTBCk8iBr/8CT8O3Yz4BxWoAovd8Mt8OEDGKlg
QXgL2NuIxYud78HberzblV7Mltj6py3iBEcxG5bFMo7NiXK8II5nmwXwLnK9
FSd9Akc27cO6TG4l+d/YOTqdQq77DEIU2xIcZ5xy8BOXItTHNHUzjxpbfnBe
zWiWwD0Tx2mymVWnXLqBnUpYSrxE+iLBMpOeZlscvxvMXdw3+42FzEi/WTbq
hlJna8rqftAHgIqN/e42J3EHmz+MJpdH1QxS3AGz7PE6ULgglE//ZdRiYl5E
zCUgCN2gjJTB+nS8QuHT5mwug4JKinC8+gOYWa4S8X0t8U/ARpMxLCAeGqp8
15Idk7lAjfzCu9dE1noJ8EPKfoVzyd/wfqUQms/Es3+GSrGPXdiSHQVSxlbl
vOY/WtZrQgUXPunfRMCPspz6BUANeMXsxX86OWNPbNqsfVy6Gr4bzUzGIr+g
VmVmYq9pcB0IxkRR48uj7v2j5KfiD1jHV1YPoYZ5FESR8BoRbP5Bkl8VTxGl
0/MxRRT7HalWT7mGU9cD1Ic+/TH0UT5X9oeHKdKSe3e1mVYv7KrcuvI0cfke
Fv1tqHI+sWyX14YVY/v4Kqr+tVcTLe2Bqukgo92FgRZTjyht8J7LxXbEGUdS
nqv4IbjNAFuP3vcYu+Sp2eC+1rgdu4czvIJ2Pn/Ddt6KUsJq/JgGxb9AfaOp
WLqOuHqhzD8iuL4sDE5yA4kMWZzx95NfbrfdbR+XAlTiuSdT6GRnnLM1oDqO
S9BbGqpuwZtYiyWO5tQOxmlwE6wMTgrNhK+hMWernOmCQsw2ynaVsnTj7pkv
Vqu8FilymTZSwhMR8X2dHFLddtNaPC4f1jSQP79bYoriUjzTtS/BYqZjo2A8
nP4P5KNzI4XGmj1lG0N7wuIcuTTrGM2iWEmFz6G5/Dv59f8vx7yiAeiQ5XFk
jsaGtp+VHLYpf+MXG94T3p29gbspwJ481u8MVluG+ojorItKG1oBDRUYmtac
y1QvlOvpG7odJaqSPDPQGsQV9ICxA0dno4+hqMxmf7m3lMwZNgTifE6gxi3w
RKIeftP2wrbR38Dcur5dBChLD8gzHKzVTKubZd8Y4Qh3Gj2tX1AlfCHt1TAF
tU0JRiONZxVV2IdvSSrcBTaY5VxxQxEhWKgE0/MOGXsEcVgX3T4BNCofSXNw
xpmTEoo2L9RMvaDBNEw+iozkaKlEwYbDSm5/x8yDxFPgBDvWKR05xbgMIy1h
gC6XqiI0gGQ7mZe/0svaZc+Ttoi2dw1to9EqDoD+60ViaWBLPXLC908W8+ZF
jqluZY1cmYzZrPDouxRMM7i9zrwYSALmOdiMNRjKisRXDU2CSPt15VWTvKzm
oCY45zJEYyhej6BsaEOEzXLbu1QKLqAw58ptDXmIWsSSZ1YwGjR8EzoYOtAs
EioXl4gWbMJcZvukBXRENa/WD7COoFHFlnAlQ2JX5cDYQzSR61GtNbqPOhRl
fIFcmiqWhnREMdhjRqRosTIuoF2Ri2679nT+mGcPrNJxFRSRhCGsx15+3HlM
+IpERA4/uYL2C24MlU4RSrhWDxcB1vJgg6dUuNa2vupoldrLJUz+mrp498Tf
jFtRADO0XOTljWbt8wOuPy7IMjSJXfPRNgAjQHfkUw2vSl5yaSJWcE15rtlq
f7eQh9igvknPP7ChwOeigXfvjZg46T19NZeIzlBGwgG+qIk3ITs4aFIB4rki
cWImMr9ugCp4r919iGPqHHcU2kojWeIjXyoLsEhYkJvcrlSYmHRO/UlhO6K2
ChW5F1+54mfjb8C8wQ3t0fRpmEzunrWM1VPngTLYLJzLKwOJI4LD+nkL/Zzy
21fclpgd+U/UANMsGqJLh0qZRDeQHnLAQlLUnnH5J6lmqtNPInwrabfTbF39
PlvSn3AiR+7Elj8zwjqW5evgJnLThZPgMFJ5xLNbk6UuxW1S2FZuWXaLJzMy
+Wf8bkcqCT0XGhzNe9l1QArGU0Zphd9TT6+BH7lmY2XmcygsovqAhYBM7zCv
JHAiKUw3SAFTWj9X36flaTDSrwWkZL/CXHfFIrgqGp76zb4+zEFxCG3IyH2J
wudLS9ecYRTgnhKunF6OIDwzs9WEBDbwxiezGrE/EIYKY+vK5fEpCR1UyEdC
JRbv9Tmc8qTyqtYtQp/fqgFxeJ8Ol2/Lfcw0ZzJW/iZYg8fNZmErkdrLRqIb
95dUNr8JjXwe1oaGmG7jc89m2+TBBy4Ardx8VBrrieO24tBVD30OmBbgu+gL
SjuKWLQlryGTuLBgUPYjGSJ++JwJ4Qqj8re1WEzt8vUumjxlqkxVpMUzC7DY
QZnGpppJvPDVd3cJN0wRE0JFCxFFSud4Q990RLUvlWWhUZY5lNvLD2Df0I3q
K9vOajYr0N7hJtEhq0JScHCh1OXgCV9IscEUHpylfLq0ZSJAqO/nzfbuW0Eq
onq5oAvbwiLwtj0n/WFVnrpgtnYf8lgIWqrIpVe/bIehWAqzmRR5sCEOCrSb
piKLa1aGC+LDNp0tyR10bZQRy+jQWowADZJPj8nf8KsHvuEX+3yvNdcTFNA+
Y3erlPc3lCHfIiItHNZCw+M0er9cgIy7XeFuTyFcYO/y87d7cb8LX8vgYb75
0SX7PO9Aik9j9I7K/8P9YEh5MuzoekMM7fHl4zCI+6uGXW2VoyJpebDwmNe1
yD8SV5bDz+VWQKYYhKPqQhNqWUspO3ib8hASZIm765JcrZvs4iwVQVJOHsjq
5qX1FflQOYxYidGzvRue9qIQWbBAIEkRduC0N07PI1906abKz1V05Hm8MrDB
LrqyKICBwsD21lrgg5BEnOvDvtqewMZaKADFgd0PjWTur/nSsxmuJ6IaZ+h1
fuMSFWEjpP+hzHTgMnt4htAdCCVTyKcg8ZrnRyrYQGDumOxLdjR51dj3gvWs
b4C4S1vBUN34CJ43ia2Ci0Sh8oJmUt/My246kaMO/aG+pwFgXD4UCzg9rsh1
tp+eTtcVprBzDXw0ybLwXzxiQb78a7mO8qDIxJBjgadNo9QEdByiOEh1Hqcd
to/lsrjWnDQT/pUshEPrRKUNOZjeMaizzsBadg8HGe1M4O2l0ggVB5oklbTJ
UyOmeI3Qxq+fre8i/2YR7gLNIofG13vHqY6d3iy7FezfsLvAFbVMDGhDALQ1
YHCnTFqqp7HVuX08dS2+ytAg7DRV20REnLBaY9uqwSA5wa/QaJ0q/eDoJDnd
0DqVZ5BuScpBzSeawvuCoq1slM6GUc3VKZed9H+upmWr6vOqea7N75cwcSbW
mK7bpReRN4jcrUcAE6m/zJgyLrKbD2LcnnvS8RSEM1+rHDnfL1dexeCorj0s
hW+zES5K+jcLrog3uZ4XLiLu8fteHrjdy+OMqvfdnpucm2H2FPkgqJFNKofG
yS73LyRwHrN9sT9ICBDmL+HZHKshl62ddMC/UZfFgt/WLS7BWAucqYtNw4bB
5b7w3Q+8LBpIY4v/3dq8u53I1h57z4T3yFwtXGxVsP0E+jEVY/Qr/FDVUQLE
Zn1kBUzmqHcGrJkze11fOreoeey8zZoo8X1Zk/nVfOLpieMiejPAa8Q0DTLn
0C7jBteMe+NdFyfBKu82J4tCHCrC8AHDtv8juAABifbHMW6UHX0HKLgAjfAp
l3f68QVrI544QldQ83QOSCDzQckfWY9pgHWKzgWceibdBWlIQeEhmF6wKIhu
QUIvARu8ns9n+g5qCgZf/Vg+lnjnXllgwpivGTMj50613YbOBfE6PeANgQbH
3DqJiBf6ImJXdsBK8N7czvyyKDwUb1AM1aHdEp8xEGNpNaUPHypDd5lMWPwy
hvBuoFY8aWzrC7xkAbrItqjZs/JPBeNVeDBGZ4lo0Bo6Td5ey829voGJBTHR
dU2E7CmXiseqHESg9vK9BXAlac8q4t/UhZun7ITpgsWJAD+AfX8LGuMb+Cr8
bqH9Eim18RptQZZ3ZyiH+VR+QB5XRvpC66xfNAbIQz0vW+kPKUOMCHuULrVc
Yw2iI1y3rfQ1KEagy8ctIlq4uFqlxInX5zYo7yrgq5uiExsYBtKpI1Ssn/uQ
yHwizy6T/4scH6dX1nkTj4NY+6DEJwQTlnY7v5ZhQoDELfiJ55OJBiQujBMD
s69qT8718Gk226BUFPkJpzCr/zthV27j89XqmtnPZ/Oi5YGua1wT1W95YIek
NRy7XMDi/VwbkI8CogXAfX6IIOd0BbY4GcETKaGH4dkVb4IzqLLS3xLldaHA
l32em/yFnUgrfClNQzNTc06z6lZeaxqlNj1UTKhMG2s6yq9Cc/4VLJjTIy6b
mBg41iBd6AhE3MURFoB7VTjQjPgUU8Zx6MIzF2dUYbw+LgNxQI3ClK3vxPlW
LHQp/W0DRENccUesLXkVfonP0BactpICGilRQECTr9bEsSQCfXt27/9E+m0H
jmk0wt49nD4dfOHUj6katRnEvWjlpsCUrVzhx+TA5dEvVxqe2nqYYfWfIKjx
aWn8kFWDVDc9VYFqNqaJWGhACRERIIqIsx+DvxT/xN5pJ7s7LzXmZOEW5abq
VBQukuKVnlksC5s5zmNPGaxc5POnCti+Udi2j2iYLoZX+lR94/K2qv+mqaJJ
W6Clm7onKuD7b807RMppoYglmLUNo1aXl/6MY/A3GUhqOIps3nhSGhjT8Ui3
ZGrM1AhemuqUdYZIRn5ThZrwOx/sxOQC4q4YSv75jiGqbIEYl9ZFnoVxLyOc
VfWnZdYNiLh5LfsyMmBXugh/Kc7FeoFakLSno+eIVW9LfYrhsyrRMwiRxCrR
2YCHztRBIVBDj2AQDvIiemMtAoRqEdU5g9+pfYIaeCSvpByYc5F38hcO2X70
HyGt3pGRDWc61YICymOr1h57tCzZe9l0f2zStC8Nj7Lh/7hfqF4qzUO3klIk
QYuid+dZa1q5M04qb+GO9WaGsSWLDQ7HrAReGpQG7amg5TJ1za4Jf7WqmqWf
EEomxQS0Lrb5puJbcfPUB5DDov+ttZ9FaBSUYj+aqaVw8w9CmXFsi2Nu2I9u
Dg9VCdAIeK1od49bInFpnodWN0i1MIfQPuutAlqggrhc0H+PhvadLr92w5Py
whZNUP5pj1oc3kvzUfCewINeb3gTAPEeWdXXnE80eUb49gakQi5jEnyV746j
ImB3k4NbtRBjg9/55toSvupzB5Z1DXLNb5POu96/it2c9EtcyIPiDxRfLtvZ
8jtHXa9NEMoPgsXz9w7rIe5811OHKdrqDXSX9Hqc7JIrKeEvYv0RrQqgPuzn
zesaZdtpQDLo6DEeBq/kePOLJtaniHmt8swnWIRXT6OHEpbP7D4y1ljHjEE4
REYNBr33HjhwSKhzXzG4IublQdkxehWxLQpn6Ldjsi2z2pz2qRJsj5HqTsSp
VQRhlvA4ad2eJehFBHl09TAo/YD8CIQR1VHHNpLrBFwLB6149KCBm0nRaALp
jvelKYscG09RN9cqegT+64GGyQXfoIu+5Pw8vgPXr2ZcrbzWpuEwpy1LZ0nz
gEM2iIydtSXEPirRHlu15ylVXuaDwGFulUh86cZauUkWJMIkFgZfEHs+bmxN
jgmKzZ3cXivZqx0UPo+OSZmZEA3E8cVqMu+R14ceRbEa64/wNZyurkaJWUGL
c9fKviMp/cNP8lw5u8axN9nMTW4bzQpPYFJcc9es5xMQeRLJ+/0JHJxU2tb2
fleJcLLTbF3darnYK0e9sfSmZckl4xO5QBgA0ckASY3yhUTfaZ77hjL7V62U
jkujOZ2SriDgxK0yxC2A0o56UOEgPGwGZU910ZAadvJKoDyG7k7/sUpbrGrV
NaDFXmXuRO3e7gzj2glTtpg7JvGqe6gSaT96vx4FqREGaHDZtnm28LjKqgyp
pO6nfU65nKhtKJdUmJ8huOJbRggWgLtTFKlFu1xgfIQhY8mlyk3iv9/pvZwg
zKRhTNuTxvWTszFfOJcjZWQGmeCbUfOzQR1vP3emj7yYmvTSQ4gWMhANzHII
mY1vR+SHoIaWcki+docvTsY61OuFylggYh0Iwsn/bPTHNCKuqJPhm5BwAQi8
L6bcMUPrBC/bVdTvZyROddEFKa/CSk4loz/3kk7VknAmbNMSJwgr1dkPSXNR
dH6LfZPwW4KIMvDNnIDgoKEmatVw/mAEaWy93x0CG1GaPlep0R8QR2J9cQcG
0cbWxOE1ZM/Cup4U/C4eTha1d825+k/wMu/Opy9hIlYcs6YgtmRBWFshiozi
kj9QbIR0e3sNdl4r0utTTcowkD4kv79Qy7O/mcSLHkyYB74v1ZugRKqYU4O3
qW4EMbU+8OH2sbJsiP8pZD6bEIM7p0xCj5lNhbZJRY4eF23PIZ3yyn02euEI
7sABf4WinrtD+W7dJTGDEQA+2I5NXrVoSM+4mb7jMZLyyKncnqfUh0VSSCEB
erD/Fy7P2sAuwxrMIBlfAnHZaDWHq6m6QH1WhPsEjxcTAwbydMvrLGjU08rw
H2cO7c/llffO+VP8uqrKCqqovmayplABD2SJj4H5josKXCt7theTM85CDIHu
0Cfkvr8oloFoeIKYrsumjDOiuFpYGiJKxZi9FwwQFd7wL54aDS6MIz8ERlZi
eKbcKdyqaQJDmHRwBvDLS5F5FXxdx0cpZ7O4ADNvnVK7+H8ZNNc2QYMbDFH/
zI1agk4poHmPnjnQHCz0hygIyOVkv3BhwGzbyiB+1NvKI1yW2vinz8A8lZSA
WalMqw29DXLfQ4qhqq7co73V2+laaviW8j01HZNUwqr9gcszClJuaU6xTuCu
B3nWscx/hVSsgvDBBztHrmBWkskNPel9V+BCm7KyBL4lcMGz3jHFQXgFoOfJ
e1cPPZ3q3mzObIsDRc6kidhJx+Egj+ZsBssQ0pmm7pyPTGuuu2vYtNleXGWQ
pFcud1jOFTcR3W9zWBwoXn0IaFTQVPN97ibQ5E40yOnNv9u8aKbWApOJbGOh
PJ/5H6xDGbzBXMiapr8kUeXubRwCN0IqEzLv6U2Po2ujLjZxzkUFTHBjt1+u
7Ho/seAIDmvLT5EwABwEDx/0Q1VNOGBQqMhqc9+rmjZZqEVg4NEb7xb3M8qs
x5twlg1LHWNsDPrFqEB+MT/lZRS9fgsGzFjAwknUmYjE0dUK4wUcTZR3rhIZ
47ihm+VXLpPlf4g9/pKs3iUnNrKTCrLtcmtp6zqphv22BbN8o16/Yook5z7Z
hmTcKwBCKYMp86XWxmAu2NhgzOuDMk/Wgb2K/Y7h0L8MwLQvXRO0a2UwQ76y
SFBGsckKjhcGgfMHY8zdA9SIC2b+nbSPt1TI90Z45BM0AxP1zcKI5RDrLIF1
HlYTEBh0ssIu6B2hk4MrlmVBDLWCoXMmrqPlu6fKqoWjPww5NA3W2XujV3Xr
cHXCtjGLWr7efSxqfadKtG/e+veMVAp5DEoI60CT9gFcasVOQWesgzujMWpZ
rjizTOgydJV7HmmuTCraaEx5FaclApurOaq2i/MHXqk4tRxjdLG+b+SfzGvN
DNYyO+4qXYKRh74o/c2GBQnRPZEpN/4tZfrokvsi9u9+Nj2wDJCSK7ZJG6Le
GTEZh9H8DoAL9JM2FBSYNrCzvAqZzp9PTNhjqvBR+f4dPFR0SXSSXrA4x1sb
epuxpfIYnv0PxZ8UdvSBrZLwbDDi4Wu7sJy6Br3UHRljSnfM1lL8RSwEpw/S
8XPTI4FZer/R5KwY736Vt5bNshIODE2RSh6/Ci2nyDUrQJL2h5idzCTgcCLc
1SqZzlX6QGS5eU+Mvg0S7+uKx+rDe8u7NEts/Ixd1uvyalF/b5PBMrR0ELvV
KoWMIX0yEQpzMix/TFUdwE1chwS8pxlXpzPpMIdakiDTy7OnCEIIXs6kGJlT
uQ38wfcB8qotAI0InoQGGX5KgjftlyLR6Ekrd+uhMNfT/UM71e4nFzrcy+v4
1DNPYF2aYoEDrogA53BYQ0s/+jRMmIm0v35+35mR4J6uZ7uCdXBLOvCIypsC
efajqjCaR0pB/RdykO2W4gQizIkTXtwA9Uy4CPsSMB5Nxh3lkRkJbbsW5WZm
svK89rIP7ovAk3/saa4sKbYNqdnosa9eDGw8HoK4g9FDimAjfyKJG4lllFat
GATykEJbdfromAhG00JmsfTL/AKbDIDfsJ2jRXnCti4f81t7RdTAZb/ebKYh
5CRE1OZq3y3vusvy0WBHV/V/OQv50bbU9gwcSpXXA4+o31eVAiMxswb7tNFY
KcE8IGLyVOHMHTAUnUtE8NDTnzRv/nwFNB72RSSMUYcSyZI3xGOVuV+AuM9n
ApgHdGr95OkTQUQUed8J9oXRvCU955OWbnzS9OL2r50cf0CoCKdKTntCh4HL
Gr0+BZSmV4sVWcbLvg6usZLf2W/UxF2Z6GHkn9Wi/HMV9i3u5iWmQm6gvuyw
p2W8QBHwCZwuUT2FxqDWP/s9Hkj9/TCm/+iGdcixnPKvM3keYFPOKEt2Kjff
fufK56Usr6RfeUy5KJQrUf7xlPJxnjPmmOJ4gfJSXASRnveZnHFk3GjcxrWb
B/7vjRRbyPIMCfcyj8gDes3Qg8McaNEZMDAGttexWGFJ5tsW/MS6zhf8RBgR
OeNVZyVA18ipcIsTZlZ9lnkk1/9RSpob7ZXlDpvEDKT30LyHsIXyjxUWdxJw
PeNRCbZJFo1VqAZk0fn5IEraAckcVn+JJkvZtO5Y6mF3jz81iWlmlgA//l3S
Tb+iMqnHLdHWJloHg0rnjzijare89PGeG0YO65KAhs1xbYkTAQaWHUfoM+95
7RhgurPuRZth61Hd+y90TfdfB3NIT2N9CxZDMTlGAPtHVnbjbWtdZfuYUh9J
f3yPvdpGCl+fKmbkvJMdnkI2GN4ufW2SUE22cqgW18bNDrcZGIco8WogJJtU
OwH9WtknQNVos72VneEZ1lQY05pp1JC+qKxLLfa6xOUdCveE58xWP9ad8Boa
IqfwVhIu4I/wCqXM4Lu72AbAuGgmos0s3rmnLPt5cOhjylEPcuKOAWFWO1yA
HB3/pEWdXXhDxa73XCucAZXdrKw3pZ71/s5BJQRCATgVQ2K2Wbie2IuMvVaO
ghuiQ0KTJsGz40dc+t7cGBPOeJBqq2I2eql6KCA9NUjEV271oSpz/p1EIzhH
3uWrmEqbVW/pcJTmeFHZFaRh0V+uBUt/kDPQMd9luBoi6saIxsO0v84KKtBo
3qExI0F95r/foCtuRZt+4LTmeRV7Ctgw4LTvvK5ga4Pkwhaqt6LsK3EUY43e
je6Xsj+REg9Iba9vej2NX9D5XkvyLQ/yZhgQIFIgVnI8xBygLhdNEhqOQfvh
JNwpE4+3j4sH59N/CK+hxyxJOCKCxh6WzJyiRXFuWOTojpEUnkkFt3ZfpUxp
9UEqp7e2SmUsLPb+ecMwGWAm9yilFZOZv5u4V5xVhlmbPGCY+uccQlMGg/OW
SfLIbV1FIlxktwrHv3jmlfNA1e6QHFfTubymFnqjvgRyiYtdoKogw/M3CM03
QfmY7AWUFjMneQCKDCUZi2xM5K+GFg+4OcQ1Hy5fGFVvZVJ56vxtVaJCTYv9
XurLURpsWuh8phtRron/Wh09Q63LV6kWh8QeH9PyKZk0DGlq6ol3Uz5E4DHZ
Gd7rpaVmlGiB6Jr7sm91N/EvULenXG94/TlVfq5zn2HyRUg0aMmUhBurU7GC
bdK/RDN8hqFTPUDhTIWXEpkYdCZtd6ou4Zeq8Pq0C115a/SYDqX9GISI1JK0
ZjUYFwLzSmyv4M7DjsCxL+gS3n4EDGTzziDsWjVBwa5fvLx4iXnnKaUWcfy4
KpN0c5yjOhELhpmk0RZoQVixY95LJon7KD9fgMO6ohKtfPqr5RG0AvVva1w5
DDMoR56U8FrQWPpkYyFLO+7g6oYqFIMpiFSFCHZo/SDSBXZP9+ukcAmvSFY4
Q1/bA7SjlPHanEucyohWDUq+2MpsfiausZ7KEjZvC3pBcuCVy4WeS3xqAgC0
fGjOexbL8vjkTP3n4XaMq3x928tgwUfTGGRqWA7jgMSxBI3GstwTZihrV6iH
hrhDHnQu5ldEkeHvOYrY/bGYjBgC1CgPLaBeAudsetmnjd9V4c0Pxi6ElgPS
3lUJE+HJ8DwEy9ZV3oKUFZWW9cyg4GTOCqeQUVsiy4okOxE9bxSv7Lr/FYHD
ZF9JQ3IJUMuoDEUMT26klEQyigEfq9RzHqyp9fkmB8r+Bf6z0Lztci9LOVpc
M4GLMrbWZOa1PcH2GuocRe/+cWUHD9bdgKbCpxi/ud7Kb6cXWdtDEXJjA+uE
07PikVwo8jLNpUUlYugYrHSnqjZZ1CRVeXb9SxOgEPjLZ0BYaGnIWVBNkuLg
nq8FdI3RA9G0okj2cg7Vdksy3L0R/TuuxMo/hg6tGcWdOGsAdw/BiIgk8SjM
a9N4KBwN+RbJCoc2cOH+TSYKSV9n4YM6Ux/+NvulYQSgOELauer9ZNWW1ziD
O5ZWY6LwKmexRjbI4ubAFabFCG9Nj+zRbiBYwEeQc+Bf0DGjoBWct4bnfQ1K
2z7Nnz8wleMG5WM85XDyxYfYmc0pmdEjY3uwI38qJeWut9367h4bmgOAF1Gl
N06W+CwMTY7g8IcjypLb5u3LwpCeInnOL8dHCLnM4v4c+nXEzrWuC8oWHmh5
w8ez/C/rgjpz0Mht2I89WQvIuVBF/KQEmX4vf7/zpfqL4kX6nuR2fojr4/gf
lrUkWU1XLQO+asYAONihilz9GUFD+R88Pdt2pNC2gnVflT4X+F7dtKhxjW5+
qwvqrIoXVNInoAjjtv1hoYvJSi31iSh0LlC1pJnB3of0P9huJZ9GgmUJCGJo
pAQCSbKy8MvvKQteoypb6GjksK/9egfNsP5/M8OiiBQPK7ck1sdrj/64Ov89
5dS09wfzYVJPVzU1ITxJdm+vWsMbPrGGrT2SZNBJr6xxN4FOYyIwIXAd69+L
ABPaRqLZ9gokLTeOYLvJzVQl2+AUvRq8FdCryoCu8ScSIm7xt48ishYFqBCB
Eu7U4usmSh3wMFEkTP2cuoF608FXXIIMJrNnGTAcgM75cEvb+YHjGGZVGe6k
AkL6nnoZ1ySO+fH3I8+KH080MYaRZ2STbS6pLSBTNMGPTp1PI9FSPWDanf4u
h4HbiJEXcL5mju/wkRlYooFx+y0ypNHwRWXDXAA17vw3/Q+gzrqw+nPIU3GW
SS4fLEyec0f2kyObM8Y4eJdkiTxGNUEdVpkdTy0Bbt8H+Ai9wimzqU6TYMtw
24Fufzr7UH/q5nUvxPYI7tuLpAf5ApZk0Qqod5xmfwM7qL5z+JCBLGehXgzJ
ruco9dU3cFLvJlwI0NZP7j/zL6ttNfcHa9alYSwzzPNBE+rTGEDa9gj95aw5
c9vPqpkMzf1nCZ6qbVG9uIxYNW09DVzZ4Bk04F4z8cNOPhAYr6ZfoPEey8RB
RM+5wrb/Ja2DEr6Fjo2GJgc/wPyHHHfpKkmgmuO4oKvl4V4tzn/C1D0jfL+L
bJEAVe269YU1Dia3SJf/YDPAuTTncFwO+mm1iFVaACrAUallsK2RE2ab2ZvT
jwacsrfd5TlQUGg0vK1mSugd3GO0FTH8q5BmpcVTBYeplitpIRze5RCD5Xe4
3SrNw2TkQyeNHHi36Uo0I09IbDl26dQlhy4UNnQ8wJuKnyUL3FElV0zDeSIo
QEhVHxBMq5e8YcUW+x+OYWrtvjn0fHLm48jlv1acOVk+5646h0HMch8mahjP
tFMNsIjXEtQpEfgR3+UMdzziL5EWVxmPZYXz11OCLR244Y6gV17Vd/A53msJ
UXsKttMnCxOQ/7zF97qPeE9jVz6hVo3wfBXOONdlFQphKN0lQcjUyGEwGbHd
hW1bHzsL4S/Z8djLGQfzzwK18B3i/b6CCaxXc6YDy+cC/HAeMeTJA7ORhax1
tzszLqXuVgWVrj63W8wl0AHhYPtXuQjWN/KH7VJl4C+zLgTcXoP9qf0lKya9
O+bihsphfP08PNi9wkqEHbwPdauTIw23Y3b9qnb+Hxcs16dJdeZFr4IFPZZh
5o8ihknlSzc69u0+/2EthSdaxQnZQdGm2By6m+yGnBBaJefALFW9m0jVg9th
3lgI93t0/kdsHbN1dZJkjwHyXxH3yPC8xTgJAzOuobueOTC03rkUZcIV5w/a
M8yecvCPKuLRE6xbmTAX6XZ3TZrKr8N5rbXDG0x0LxqIfvl65wM0tkuM2B6L
UwY1eAOUjnhylOEKOEp4Y5z1Ge+YTLJbiGOBI92Jqa8j6sVNMJ7/atW4vGiG
U2AaqA1HzUALwHCi+hmoauoU7yFCt4aqbOMoN3HlneT9xaXp9jJVPRv7Km9u
d66vw4wtu+eqS4PC2VoBFBFWtzaVwvk2ge7+5/PwWLT8TnifKlscuBG122i6
lV4aDfiIorGqNBq88BeI7QCEH5B2XXNSKszdsZLRwsLk2z1xtietbAM9V6h3
Cozs70NSiBP7Kc9iboaCOK0jXDI5iAyc1HAMSnit07wDufLy2H3bjEYp/gWy
vtp4dXz9CqTptFekxH51XmGyhRU2QEz+vB0iITOGWMUa0UJ2BxbgZeWG7eMF
UuMXT+wwb3ZbqxGk5fg7FKh3fnNxMozXtYNDR1SqZXOpbr1x5XjvMQWO0FjS
8PmbOhSHRulvGec40p5gPIElQ7LdeEyQitm0Ecf+JFoe8vuX6jjOJUuUlPmv
9+ChYSQ6H+8XibJpi4lCTiMU/RfdG8WB10QglYCpxGaF5IIigQ0oRkzjZsNC
CXUn+6KWlq90EjyaB8hGWudiAyKf6r1PBWd8t/3U/7T4WE0esplEMw47ar+e
IwZdhWFwH9rzVh4rkmeFf2Ch6MqagZRxiGeyCSMDuswpy+35JKG5L7px43FC
SBNhYT2fsXwdH6S8jZgo+Qav42f6ml58G0Ujl2If8wK/V2hBEYMbbEPgFq8n
jcHiaXack6iwH5+hpGakNlAJ8GqBanFCaSrzC8T2sUqVLUmlWeh5b5Pt64xN
D7mYnCCUoraF9n+UzS9JemD4nSQDYgv2sjtnV2VMMvD1PwCAnPz037pDvxB3
4jcqRkl2BY/T6FxQDiWXfU4STHicFGUN/GrhVLA65kFn/vFwecYgX0ftVq4h
WC0CunFn4n0XQlWM4USvAQyJ0+sQuHc6jZCt40Ge7+awsL3VlopwkbEKSvAH
o87ROfv5OLfOJd2GAR5QN9LVRh32nLV3kkYVd0TJ/MzwrGDkNAY4cAwjbMM1
sn5rkDyGD52H+CNQ0W+/OdF6CUh0+QV17qYhvqOe9NG/9U2IDxxlRg7KtRVc
pFi3rlp4cUuRsbnaKjp6O1S3AIPPwZUWHm0gK2duU3BVpGc4DLHej8hqmjhB
5WwvNO2sC9jKWtmKYfkdX4O6loPhBUkavHB4UO31sv4F2nS32KVrcdoGzIwx
VvFCWTi/OHm51HOom7dBnaTfE/W6p9n+aatrBXFJzUEzbywXQd7uZgIYXpzX
lvcRnYoAQUy1h+1M5g56hCmUIdpwt07biIskfQhScv5VwNuMJJPcd/Mu+388
MuYRN/rJE7cU1OQmJrRXO9gGuDSLOXewDg+yPcxJKFL/W5QEmaz02cWaG3sO
fHDwJQlXP+hrEa+zK0gNhKKfnRdtY/pl2TmapeMVQlPsow+tHMmzHCWquN3V
p77WYc/5S7UKDuLHWZooQwvyJUNTWwzoQrFEoTZ0Qa+lwcKT+5o1rM57/vgW
DhTFrhr93pEWvrPXkfAJYGOYVjvfVCrZuSXh5cr93IORWRSyuQtRilDMM6CA
QL/aX1HK0O6kCIthB2iRsAHvBBA9i5DjKQSlEqoxpSWJuCE78O535Sjuw+nh
CBk1swHIBAtVeo1v4J5QZz4Gf6sX5EGlvM7O1iztIfPJI5x5HKIzPt+o11Pm
S2doINn9VVRqLAkKry38gdmZGDbPBLXakjXap6JJPcPK1RkaqN9rnD5PK526
h/RwspOGKMsFwkY3IU5TurMDVdACDEt+mZkMC7nbnTjQ9xqJ4721bKp9755E
n6njGAjRXRmIlb/K2ylhG8UVn3PmO0OHbhvlies2VNpFacfyjMqLHCsDhr8T
GR4d8r7br2kE+piDxiSYPtjsFtkmYuc3ttKey4/e85XhDLxC3so9c9FihnxK
R81hQSd2C+XPnpF3zBQTw0RmaII6Rwp1M+kNxVBjrn6g5S2lP3fXQLmDO4Ui
IN3Nhsu0Q+nId0TSL4gC+ytRszRiC2DwU4WLFrcDeL8OD15+Q19AT8Qz/tdq
ZGYAtHEp7YOdrkZWN7MGauUZt5SSzbcnCkhImSc2upUSqlxsg1sOkHvpA7Ye
n/CAtBfpGzf5J4AUJIMubE2IORbJXTuQaT8N2nfokdob1/NhrHy7Eqeqoe2v
fV4/sbklbwu/pxzlQrA1CNydEWm39c3w86YYLhnbMSyeAKB9FxqAJwiPN1Td
WeE5yAew/AyNdMyEVnJPy1BP1PfuBM0OxGqot3v0ddhojqh/T0hucfhf08D/
O5RanREzfwcOdfhJonmwNXAZMyX0ukTw2bUs6ovO/ICSPP/lGvHJxN08sWuS
fmfwIBVLolmve6P90zu20TTrUasgA8ljPcNNltqnEdhMcMerRbq3CRlyMI+C
eFB6jjReMzD3+9cyRD15NgUxD+B1eMClztr995SuKKNhdWEZKNk1DMZk/yli
81iWoAhkCoEzxfIKPem3w3aKGnHoXzxZOJpWsqLcAUdBQQLc+0HUpr7M6wgQ
JomUjF1XflskJdZRLyLouJ4eYeELNXteGvNFeTvclN4VORpDRbOmef0RlRk1
WN3+6+M9xDPc2r28/oIgUtT+7Fm5d4cPN6jMfwLhq2nPysHZJFizWRjTIyo7
awUA3k7x5U1e0zYFleKiSkMUqssnSb/yKljLUDb7i09uqaTVbLPNnosQKx23
9ehibDhY6gS8F9JfY7dpFkiy/3Bif0VoK3FhUsnHJ+jBsfCUTvqz8tdj7/vc
44zuVr2vCvWR7SAkmjYhGLV5HZQUuVb1W/CEvBNdRJbtqu8d36G1AlPRbfdK
AO34y/Bi5dJr9cb8rAQ8ETFijLdU5LPh14fzDFGKDOh66qPqVH72WtJA99Tq
oXI7OgEQwEEUgSa9A20oKa8bf1xJmf5HppS2RVSSIFLUpOchelNpireyAkDn
DknBpLZ6ZrE7O4LmxYqa5SBkwoTMZX3c/1Ba8hTGLrzGovWZJ2ULscsxv7Ju
Z+Zrerxdbw/wPrg04Qu67YybFPkyQlySaSMJKHW3PgaqwLQybcfvdePTbMpt
IMODFzq/vP+dLE+87J7wemV/C+sEx7uwKDSqxcHHy1YxKhod1xc+NjbosR2b
E7zExvjWkMqzwkbyDuPmDqF5xrKnBj6Cd+KEow7Mh/s8GW3ftHy6J7Q+de9y
AiOkuAzaC8NBeDLlCwKqvWOgvaRAYL0RE5IwrAXqu1KXJzzmV0BSc9TWQzaM
B6EMzI6bya0JKC4N8yUqYsVWhNOyzBY9+8cXu0cWS1crBZ+RQ3naznAwhu+2
KuqdqZe8diH72RYIEoRYdxljtiEQLOvb9plwb9RXuxDVvPGmxJ/TIyi020Tl
zY7e/eQP8boz+MvkQwO46CkQNKExE8Fu7H/ooBH3l660Nq2DIDNc58qUXqdf
P43uiIVNJ4d+3PDCRj7U0NnHhE4CwXOH7f0pVChtqm3ronRR+GcnIpmMuWdn
XSnA93Euz9WJRCI2qIAw/w8BJUW6sIPS0jis+2YWu3adbpQU6J4nhdB/uu06
SPYcqGfWV8uEZEorne5wOLXNwhyFctCgzZ76CKneLiuyZDkcf9CVX1F+4o8C
AVvbRYylhG9QmjlfR77pvz6JOyD38/354DjZNoSBqCHgRXtZMDwQxpiaKqHe
4QfdhLWTIZ7GvAWctHzrwxvchckBCr0C0xT6zw1TsOtBhD8HUBzAPYgkZTbU
74xHavQ/L3zjDSl9/LYCHQT/b1m96oEf/nRps/Jq4RUUMafF+iw0RHqrcy+6
2zGzYHrXKIVwLBcLv2N+VoRH9314pqwcQ6SFiJuvygFdogjeFvAWg2zbbjLJ
1AoQ1lBS5P1NdEquT3EPlMjb9Q6UYETjPW2OtbzJZCln6U0Nc5lBlFsUxpDw
TwWcMFCFOAFi++MDPOnoRTRS8CWOmrTS/SP7ugcdP7mcrLqh5iyhm/uNkUVg
fRsHtycZpr3SriKRnFZMTGPLKB8a6A/QymAOwMmolIgc+UZIujz6zq1if2op
Y+M05pWunKVCCJcSTYBxI7pIPTpCzN0ARcEgJBU0dqWbZNFIT9ZQ3hJ5ZmaI
hXzG5hBt15T6zxVNOw/IoBvkRqnkCF/wgQueKcBxFa3y4+MrSP+rO7ZpSdu8
dnLasiDz/3qhw6PBMNuAjxkcwEqFhdFq40+HX58jfYl2Wp6ySKwy4d2TG8cu
7s82yN0w6hl7Yx+A7a+ay6cbjaGErAh565iZeCrCPg6xxljLIwoXVy9Ox+sn
3MBugOpvGmW6ilbyPZd24J+gILaac1dDauaCJIicUmasF+JiTK2cf5YHaivJ
ewWVu+DuHJW0StI9wwsTj6rRMMDaufCW3RIyjfDbWd7/cky2+5Fip46hllCf
OEKMX3dtm6x3p+2CM2lDuVTPPxcIgsxgEEYGu3GOop6GSBsCnO6bSacahrcG
ujuRDcRs4LE+csJDlyhv0hBLdAAeULr1EE07r4tB4yXRWAEFRxuHDF+hJUz+
8YwkxEgeLEE5lM3ryxTNURaHTuKGg2d+R8mtXRix8TV2C9xDqsreNWvQD0/u
GJca8c6B/+2UBZf4TnvQZOWS/IT5yb67N0laIbEemRtP8VUlnwGVkfemmnTp
lHoWqgpImc9z1gTvTglRJ5w5IjWdR03cJlymSdJa3XiyozbyEpjY5CIrc+/l
mS/n5pZKhK9fr3xv1Zz8W0MLv4hhw1mVN6ggiUzVsrRNC9iQICjg7/Nhafi5
whISD/k1yYA14b1N+Jy0NIPLLBclntZZvbiCshLeNDQ6oqHIVZWwwAjLlCy0
AR7Ue4xLHehbhVB9SIdn/ZRM4hlkEHkoucmtPAb9dtg+nMW6rutxw9fQIBak
+3tO4M7PLJxs7IiItlZoZHuNUqlEjMuy8uT0VuT6ZYv8q3Jm5jocvm0Lia52
xjTW4tia2tXNy3zBr4M131FOmQUjfULiIJFVhWkNwv5vHW5DsBF22zaeqaZW
RmCo6VGsC2vUJUDKIS9QmxAG4NpSZ53L3VOGpZFep/2t/z0uXPEGEyrI+dXx
H+pMcjaWl2xXE551s1n9stk+Xiez1+BNelDTNcUzmydbpOV0hel93pbcPSvp
rKr5pZYonhE9E4+PU+49KQLDSWY9F5cUa3rotBoautq794dI8xZppMQ0+z58
MMQga84oJmxTAG3G78lj2aNyzTU/Gp8/ncacb6k3V7QbIompPN6swoP8RI44
Kh0v0oO7JbjqY1DCW0NpBGj6rUmgrRHrOodylN+wdvSNdnufhT4nytpJbSgN
Cpw5nSK9B/doQRxwdwDXkATts6iOIAZ6UVUPnN5oC8aJIgRq6brTh++1+C7T
OX9P4D5N7tkqVI9YoD9gve+8VFnFC/EPqFQ5I4dV05Rziafi3PD8kDY3mLuV
WfKvhi2Oi8HzUHH42926WfyeGoKzmvrLPoUmv10L5yr3/eb0rz3XriE0Axh6
pK4q2Lxmvc8HQDEj9QMxNGW8/FgnOmbkRcJeQ7RdYeIWl94DNlYSf5R1xCzu
bAaAYcxq4AXwV8eevrUpqJCyW99YFe3H+unYYQ69R82VqN61xh1yZXgYvI4I
kgMrZH1zAlbcJ08LOQ25oGka/9Oyl086oTaIF4CF1kMl/QRUmbqCrIJfuvq8
zhekhSsfajtyp0hcj+bj3/vpf6hydp5In9TjWwR9NwYA3o1WVfZYdgGhLeES
iUKkcGTq1REPAMTrd8xKHf61dMH3/6j6tzzuPX1tg2ML36AAxbBpp29bzPbg
KHULZznlqGOwal4QK+c8pbcjMuhBXzopssWp2a22k+DQDqHlm8ns4h2BGNAv
E/r1aOw8LLrGeW5vOEIva3BZKEyhlU21NL02jL+LM2D1w2WFaVeLrow16GwR
xwvwbdezRtQ/VTJegndPemhyXeWfLeePBDVRyQffI62qJNRXPqmNghUYz0h4
AdZ0v9O2e8CmS/+rrg0LIsJMsXTuSiWqZDQm0qc3zcmdimVV0bkFIYr/x1Le
m9sYtRDHxoVjb2pB0bhq+a9ihPagrvsfiKTbRc+Dy6DCztk5Qc66L4cj78VH
uCNL7sxZOi0JhpTDJW4tY5dzNFZmix8uaS4Dw9ORjLHRXdQULcPXak+cW7ev
tIlNdCgkDTxX94iK0KYsb6VfgXIld2C0yknnev3ojWig6xQ+khQ7wpreAISi
H0peadZ8asLo3x5hUWRRY5LpjRHkfn+vszeehd14da+sgSgJKtGZKdIKmmcf
4VGi1KkLkqZ0X/cFfvM7I/HyZqAILp3HDZVdSnR8cqZd4xSe7fGPg4IIEExA
kBOBs4wt2OMHMHed3TTvUz30nDQ4q1FQjXDXSrlY6mocfR3g/15edU6e6S9S
bM9QiHw7i1vpfjGXWmmd/zmU36M6byUqr4oxr4Jsq4HiEIC3DHObRlzpsoTu
x+xDMmeAcpfAi6oN/WM96zYMbCNJgDHZxoA0uPGNgewgqjD08zsPuOgr8vPQ
vI76jtb2zlObwvGt/FaClFP1gt46mP2iF0GD6euN8xF+rrSZSaPx3K3WXAdE
6DxdEPv02I6N5z4DQKuVcl8uMKtIs9VR3obXbMlVBtA1iv0eUpPU9DOkGw9M
myW2iiKiyGMsTmhH4LimwXDN0QXa0Sx81zGq9RO2IC5vLuhoFr2bKZX3s+/b
vyAQk4dy1gFqZ1k3OVMl3zyK4ilevUQIBmJ7UgCm/eT2XgElU7F3j/gEgJNw
VD4yasTE0+xUN3nSfH4EFV9pNknJHX0EIt09RY7Y2jjapRHyYFANoo/6CptK
3yfYH2WY6iKyP1SRG9m2rBMKwVSMz59c0fBlsIlcc/kTJdIs5mizdEnk+CE5
XJmIV52lPMhicnDXudpHOFZGkd4p0afPpppaEN11GaoxpHHQQCasxMHSCNL4
ytwmZ9srrd098spkMV7f0LzNuQ4mSLaYkuXFziXiuo2K3zPqLql/8SZ2nqyU
cZ/48XdaELDB7i2/TKB4ZhgM67ZRHBdq2SmWmT4kTaiDDyZG79Fd1+F5guPc
dNElpu+GcadsJ7Muzh/1rOAvRpLsKBbM8fnFZjsx1FRWwKOBjOA7D+8+hRIJ
y063S99d1OgNPKEIZuy5Jg6aEzaUkmGKQvL3JyUdL4anB6qPrTs7KQvbGP/j
a77KkGaBIHc11Ql+4Kff4tABcudWCpiU6YXt2k61rFDMFFCJJgMVva4sZo2M
npWSODp+SEoT1uaFgB7dIGOMTO5paluvSw2HQTpt33SWLIMnIv9asV+qv9yx
EM4hhu5/sagiwz/ywcvrAu9GFz5GoYsx58eb+ae/yVdRfe9gSjWyGMePoZR2
9RzV2kgHZMgREaOAO/aWThPcGsNWzH2VZaQTcTwcu3P8zAFiozBuPkcM/wBO
od86Z5QcpK+W4zkeqaOWDJlbyBmDhifC2v68RhfmMTnd1o+Mi4Y9uEZxuzgw
cYBK/BEoyBPGAjPsQ5+JL3gn7RTd/DiJmev6Ii9VMqZLgyKMXlZGKbQ5jwj0
Koqfoo7RQUDg8lYKbyuD3rBXmx8rGKXgct9VOo7jQGydZ5olcd3jBfdgdgdW
+uAvcwgS7WKwGS70r+REpl23rKNS1BM/XSmUC6rfILxu266/kr3GfiHPKRfL
kEifiCV24Q6QXOjY0ictuNJlbEOqZjdvnxYeFs1gf3uCVQ4rmZfhB0gdMVAh
To09a/SKqV1e2a1LUna7+W3mRpFe3plEkfNoTIMf+ExutCOMTJz1TnlF0vfz
QnNAqHEtoUFNtPt0/Ps/HAJC1wr4wKG2jGSesm4DIGLIbm/GC90ka0vhHp9z
B5agDTj8qtQ7eQW8noj6zxVddbS2eGM/9w/gbd053HVfiemC8c5x6rpcoyzD
P/IfDcRJWx5X97H7lxftYePQ5qWX8mfPFZFKkmZ43XjeVQrUPD89Ikhe5aGz
Vlj6+hYRp9v8z173y9gJjq7fKSX+FgRbQErOkbGoxWQaLtA2ocULEARdKoyL
Kv+h49Go3Q1tAV4mgOW1Sr/U+rq0WsskmKGRPLjztxUFAPpD3vO4g4c5UBWN
bCV0xayPb5NqfjiLIxhuGc8aWfek8zejTMeDX8PjxFZcHnPm9W/Vczd+F+VE
6UMfu2dIg9yr06XhfjBVIYlt0KFBy+KCI5dX+1ukPsDINfJSCzdsvAuZlv0G
v7jsBB3YsL/z/AEukmtVW2o1ayhdyL17xpju1IzC2qzxUb+QA/zqNoPj3sBR
3xpGcoXINcWeBMF0KAnGUNSWhuJmGc74HgKDEwyv5QDF0XPLnZDDOSaJvb8G
2AF4lxR38thuCOJUtFrSESMAE+1HjCI8dxc/0QMzeoWHQFiGpHK13DpXu0kE
co+79VTNx5uKK8W8A2JVOpudejsMeR7j0xMBixdgdc3It7OUFLnNgvMJzPtD
yiiTocWXD5SjO0I4Fh+9eN49ljCs5DVmWBLY/AnvKrrqZsQ9L4xMwl3/THbt
IdBhfknyQmfzL8oId9mq46+4sv+NDsDbWHAZz9UINf1adz63YA9C054NN3Ud
ZP/XgOZrQNTbGyiwsyhnMQa8YESK38hYTc1CnwG473ut66dg63io1mM/Lr6V
vN6dzi65UK+F3SaCX6rEAmzwINfCo8ROTsJr0jocK+chJc8XUScsqknAvQzz
h/AwpBtTUgNyq1Jf2oHcYW/5vHmSC1FOuzG5vm1eoD78u//MkMJAbVEIcjEj
bbMcRD4GPHz6Dj5/s/dvyjqjPbg0+RXO26yrDDqIIbS8mVBTXLzWw9UnS4nv
iEDt38xT2wBASBFyexb1Vebyg9WhS3vdOGdhTve0S1q80aT5CXLlDJSye/lR
uJaNkvRzbh8MXr0KVrSH2ScN35xbVhuHMB+ZuFFtLdcMhoanlp4vQc/UPpRC
kntCQbOeJUWKQYymMwaRaGm9eQaUhiTMJ9CVC1Cprjmvg3xUT3ii9TffTR3o
mFYYqcQTs72srA/oWrfOWHUX7dImcRKojXCI+njGxUauJdzqzITL68Hx4AoF
C6S9TadMVolqsnor3EIfXg1sZrXTiKZYs2c03lPg/pEmibeQu4VdvLPkt/Fn
z3ufriYnm4g9K7RS4MVMRl6DkbZ/ZDawu+cpYn0/fMVN7pLdEBVYTFU0BiTq
OsNEyAGSynjtZgrlEMqZPVt8fbXGA9PlcX4xOnrRYrmv7DVGsfV5xNMC99x4
II+lSYpQqBcBgAOqLmL1lMmHnLtNJQVq0SaFO/zLts9DtPhazj82mFAeoxhN
hdO3xLNrhzniJGgMaYKcUON0pJ/fKlkxm9JMRmpWTj4wjzhy5+q+zUGF43H1
NasfX9gACEn1reZ/s8lcf7KhjrVyyLXYXK6o2UzuENzxWdwVfZkhmPOANJj/
yYI1cQJ2sJu5hDeXVvzuDuRUMP+frPDAsaPaB2mlsEV8Yp2aGavsqryhV2iI
5Gz5Psw+1+T+Vp22uGkq7gswL1WbRB/MniBCIclNgHIE7BmWVRXuMCp/k1xd
AkfylgCnxTpP1MdI+R6XDGVIfWJZxwhjySdsArGOOwemsKQRP5jQS39FlP9C
XmmZlJkQgzG51gDIxBGMakTIo+H+MVrepBjHeND2JS7QHVbf4yUMPZa2/cRo
svhM3vfQKg5NhVxWpzphs4Eeeyp6C3TvcJ21rL6XGOPSKBXnEcFEwSZVj+yK
0O+u2ICzEoAMiC1uqb23B1gyTrE5S6O7ONzxIY702/27bgWsDictvn2//sj6
oQO2vcywXD0UZWtWz9wnNUF8Va+qjM6cVgJRhwGR7yWzoCPnJL4pZtKIDxk9
hvHi35+tnp+KRFKjBmpMBvWgW/GZmaCk+xb7h+NRS/Kco9+LXoYpX18oOgrQ
71EnK1SB6SrTe3bpwCNiE1nDGU+9/U9GCG/jrea5/Ka9qj8ImpVwMAFWzBWU
6xRfyXA3f15eTS/L3JI+Hidu61X6fIU12TQZcN/hMWBQNa8yS6Da6Hhaqa4n
J0YP+G60+Krsfg6dZBj9AZom1Zf8VZRPpoKhecekN/rQXLrE43xEuV7iAFnt
W6kHit64eLZNTkvjiLw7dGGafyNrl01ii/KTKTSyPm34qfLyU6U6mG1f/pfR
xHqHrr//6SvlIO8+b8qdCo0HfTzrXMSGPQ8qD8rM2+pHUUe34uUzRvxHaaya
qL/iXgFh0SKZzq/qRH7FoHbc8/lyygx6H7ekroFjununb+3Jrp5ZI5H5/7wG
fQrjeMYeQTC2K8NF5SCaSWT/f0GOkgyhLnskQQaQDBj///yd8VWuAXNL4wkv
4M1yEPkpdWXwzNiGypOMXuzb66fdmVnu2smQFnkA4ZSQ1VJOT8LlV7Uyd2i6
T1lSxY+9eOEMv874zREFjQeVNxCfYwKPuOIgNRbkF/oUKLJTq2NuheoZdQJW
OnOyey/e2SlLjM/lCPozp2PN5y/UpLbURykLAxB7kuikI4hX7xLcVV4jSe5q
fqa29jga2yED3fiwGUv6y57aRpmX14HdiyN0bDRaYt5xlUY/h7tKdspwC7oY
/luvOPviXmpVOnOrHizHlf9k2zNenLrIyfhkyAjbfWNYQ26Sj1+NbyfuME2c
xOI6EhdF/TENn0okPaQRJ9nriq7Q2uCpuec1xIPNgwvDS8X1PKjuZoSeZzv+
aUuv3C7dE28AkCs6ZLmAe6/3p1tOHq94l/ZstU66LegD3dSqRRMzy1RPRtA0
5j7iVGQ/mRKnE0FJzV5Kc0gDVdxJ98U2IJ66UmCpNmpWbLYoUweF4jH4NmI5
FnZrJLeyPA3iEzn/VW6Pfwp3W9TL8BppCFE8t7o/TmUKe0oCw7gCOCsYMQye
8+tuAySTlZzxznBCcWugJdNsfq3as6VOQ4kCp6qo2CnM1m7ztRMSRHhrC5/A
eHDeRT436r0koyI4mx4yvt9Khmb7eS8QToYQHDmGehuhBxuPso+uAGG9LAfD
4HIfrk0Vls50A0y7xJfHRccH+WHVbLIjXVAqftZrvgCIGpfGaNEsE+5795c/
H+NnzyFxX9G1vZxqQwYwo0rFbT+e2+67dmkaet6e+CWrKWRwNGZQkSI85BXs
RAy1ZMuKVyla+s3Ab2KltcD82KwAEdCzVpN9cqzgDkzY/jjWaj+hK5s9kzRY
GTOqWeZuoIUAAzrKnfepJVtSyC0Y8cOMnUUCPwKrJ9fFnI1uAKfzaT3i1sT4
CsVqfX4BFpP/tWDR8yWzJXSpD3+YMJQ0wPj0e4qSfFj+M8xYa0pcBLecZre+
7MBoGPv1Qgyz3tok5uPeikMN8zj9QC1Cqwgnk1NtmL6TFMJtwK0abhZ5kIDQ
X2snndXC1QxlxZRIO6UQm7+PIHoD8dyt2z6EnFk6fUYVTFqrUwrVU5kOZgjf
HmYzXOXe43imJwb+nP5EISayW3eVx54qhOtoDYU/0MtXmZe5oedvczEmYJCA
p50Vuw4Vg5FATlLyKSYuWbJRhWSFtOoUmAfiOOYSGUNeTvqfUjF0IKBVnIya
meObwLKBw7ZVUMeWbSyyDF+JNyGNw38NNIza+156fxzqB63RWFjkfPIlZroG
eeWYgqrcnTcSjl49EFIPEh/0ZFd2IEOX5c3G09fmhzr0n4G3A/RZgxAtMYOV
G2866t5unayCfS492mxULSkG2v9Gskg+YrQw7rKiC5bHBA9pZVdo9PZF1KIm
seXs6+s03Us7nkvrJCcui6fYkQP45rlCWMA0XwbNjUWpbk0P5OssgfUg0fDu
0FHaHtleNOhs/2dQLGtjcnla4p7wvX4wkZnaYTKjol0soqs5paw6NWo19g3U
naE4Y1kV6nC3BwWee8FJ8QjOA6c1OOTs9EJ5U0HDi8g7V1RABav7i9fmf2y+
Bcf+boSbzAtkU+YNntuA6Pjhj4GEqFaZ/4uegmdjVcprfPKF9XHA1YGS4BdV
Ts6tcviD7CtIzO+vczV1Im1Rgf6U1gKSI5NbSz35Ifb/TY0ziG0F4Z5W/LRd
hXRp7YOgSXOTs/SNg2hrqaHTjNoWYhNBiejtz0S52RvleYN6LFjjXlb0kZ4Y
9kEz8/neo8BAZZoNElpSBggEsIL3QaoTB5pMpcp/M/ptV2uAfnkIyDpC+lZs
FNccOreR1DTLp6dnQ0ukGxQCc1mkOZTxJjos2/gmWooONG/fuVcQsPXTmDBu
ETDQlubkzBg/w1GWa4FTqSknMDfW0OljvrTpmfNnENefTwARQ6oV/keKoEIW
3yTs0CL7FEDId2PdcOev75WyYBj2ZJ8vhLnwWZEOAMnMRpXYiODb/Bf29BdG
9/NIS16V9J93k2aGFzJnFYlYZghp0x5lzlk8fG94kuqL8tjXFuSVSbZ/hDJp
u5bHqlQinsfdHa28NTKSpFFvbZTcB2CNAsIlCfGywQQCohsbRxxQUcRg2WqD
5NNzujy3YarVmxFzAbr1DqZ9gUKe0Y6uOrOmxnznOrAq3qww46vxF/gtI+2D
J/CUa/32EGfQP68cAFHrO16qOOBbl7QRBQ+PQOSfNdiHHm+XdGzziIFXKVFZ
50v1vuf0C9SioL9RMfbofsHCvmyUo60SEZOPZmSCxQPrhKC8uKxsawTBiQdK
jr8TP+CnW9XDGjKYm8ZbNxPuWz+BS3TbcoCnPNzyAQmgW4KHZYcmad4CIzKE
cnkzrORS6akrKosp1JgDCbIeH9CAkVIYq855RY9+jbrJbUKyIuFexl+7yFrx
0NP8Q5DB+9hxiW1bv03xi3Oyc7JHMzPt7N6w2X52YSH17geOZb9A2MLNG46q
6mBQjUYgMLdmj2I/UDa+YDmQN6bDQf8/uVIJvwLh4qqJLBxkVkFImfucfBOb
4y/ktObmWKQwMnpdb635oU2+tFxee9qiEEzHP9Nl2fQzwgIth3UzDaVQXExC
BOJBIXohMdoOrWk8Yy07apLqe6LOUZr/M/LjUJwspnygAn1x4e3ZlL98YDkv
7FATYDDk7Bzfh3SbqgJar12saV0Cduz2xq0k/Yj/OyqMO1CDUCJM1JGpay4L
/kGQUKBqmfnTLSCRxA7PE6YIKezrUs0xx/t2NRuSKQm4F5eyMUO6iWpkF8yl
DbfJ5DDjcvk+/RvzgbXrj12J7QhSRfB0foHoKy4xY5JdroZhNRHeJW9e464B
7ZWCtrzh47FH9vGvCTtiOfeKEyVDeDzcbiznemAiA5Vhd51T95A+aiw0Y52x
KIg9RChSaVjEONKOpb5hwF+W1r752qV4tlGSQzQL613NA98G/BFYJDEAktDv
ZdyUCXPrIuGoSWENPcV2llNVr+nMh8YXZY6v53u8M7uXmkeR3j4IYnmJCLuh
srlOn6P29/MAN+08zXnEQl/5mlQ5I0kbeFjnNFf84celWJj/Bzw+eoVrJH20
s6t4zTIkhxFAx+HC5/GRXaA/4whDYj2vcvt5BwKjYxDWSakqQTLY99A+ta5S
XTakJitLtKrD03XygHfHKN4gzDZGP35Me1oU14pOQal/gf37lrl4GB+ju9kT
iY35T67yTQWPDoKo1lXAsBKrQSeMfw96SeRrZbL7Ix9HaE0ctc6ToS4w4knj
fB09GccPQ82U5JuOXAIx5btaXgCldyZL+9OXFgMfM/4kRtXyKhxrNYoqQUVw
/0xnEmQuZHRWeDyJDAR3j90PBW/GDWPXS5VSbY9jZazV8i28sohs/LwlCuCr
5KxCAEaJdhyqq87ge6kk4ZsOwTJ/0CBGHYUrEctiFxBVR4TYVIt1yHv524rm
3xvCypsPIcXuiAbd35eP5kSlSM2hkWGAr+cAVq6dyBDYr91dnMnH1LpDstI8
zU85JlBj3Mh+oKdPDYKIDWdhW6g4KsMTjDK7ROAZ7a6NcBljYuObFLvEEl3o
m7q1UbHLYo63Qcv1JWHLMzdvpSNWS3ZtJWWVihMup7OhjKpDC5PE2MzBnwMd
c4MkgxulBaYX8NO2Ir+ibQvgMm0zVM0BzVennnm7ftS1n3rru87O8E055v19
R3h5GM6WIxq/RqQ1IrzgvCv/7LP2AkkFQmSP5l07IHLQGCWkqJgW4gBtDpPQ
TvTi1DmhtgXDAbOAVbgq8Ef1xOxeYVMkBAcmhstARjYh7Dlr1IGNn7n6ulRL
2gdP5/la1P3oUELvqOqCaES7g8qlJbJ9FMqemeNGDS9R97yRJr3mure38RWO
NnBWR8eU5w6x6RZiR9Z3SkT1rU7Ck8wu/pL75ORyQsdCPnHFyj2rcqEEWrPk
zMfxu5aVbl/pHrX1iLluWU5c8InoOG6+Nu9u4AK7K0+MXKuve7VXTDAyiGwc
2ZmIrm+NLxGHPasfSYXdFvIC+lFYfbj8RtJ+khJT06FkC0jNqyTsfOzhSKQ2
e7FAFFcppR9JdC7pVRf54r42gy+z9BjF6cdEHq/wtfYHQL1XmPkRO5r/m8tV
6R2Q5ZVfC/qZXnQCn57TTQpil471wbNMT5ZwX6B4zXCrt0jBv47RZYinWBvE
d7L3r1v1WPUrZS+wIRFz+2cF4uL9hqmi78k6ebcm0QVaCNXnGIV7pqXG3vq8
WtTPBg6H7CByt8KOAYKJ2hyk8H+iU/xUeAb/fnOu6VgVn1loueZS1XZhp5wT
DIqVPGpzGji3PvVyII/zIjYAZT/k/QGq+lIlH+ksVuPq9gg2k80MmxeICYfo
QEl2MQBXY9KLepSscjEnHRKOdSo3w7e6dB497l9e4/jyV3d5SjOJot4TmnJT
/k3489epr+E+PeQaOJ9NomEUy5P3FMibO4aRNgkhmBD5AVsKjoeivlaW3Gxs
UUu8Q7nvjB4V9zm60ZVD3/ltNtqY/1NBBMTu0ZUSaJSw0aF1QuEqR0CLqJFK
4S30UFYSPjZR9lyTn++NYLEOgznBCr2Qljo9CKLiLgnqi9t0WmKmMG2hGyR8
tdU3Ydy8xPlPtS9dY0RYXBLkWl6y/ssZ7LqFF8o0FNITwlSLSwlT57+6rFn2
ANEmbkaMkhnUBvkw7/yO08sbNR+9b2YNC9CgvMkuGWT5NDnN4HzEgfpOcS/0
AMU8YI6KonMwIA/er+GzLIjUn7JbzCvg48imTTwt7eeIWowz7wF2CNzUFH3t
oPDbDhz4kvmVL8Y18iQMPEtiKdB902coNe0sfIyxwuIM2zyI6X5CHrjcx2Kq
7nDpntvY5LLiAdE6e7Oce1Sbci+FL3okc/ZFTmdv+/lu96SFN7Tii0uHeX12
R2iTf3pcAvRY951n99FZyRIyzelyML0AJLk/qPzS8bYS/w891zGwhIiij6Mq
JhDG8w9u+olw/12qLulHT8fVkjszEV9t3FvZZH9FcaONShQK/cC2hG8EwzZ+
Q4agJFuPTntfGkcljQFXGnuwWRRhu6etf8S2LCyo8fZ9Kg0rXFa8B8Ny1SzO
8utlnBAFmX42X95y2MJYghO1bcyNkrf+55drNQXB/HdpI4Or/t85Ezgv8GnY
eOT1KGRxqCN/8zS9KivPwCXVXYWR5beL/eTtkAtPS9nV6j2nBSXB78ixUXgn
BoYRQ6fJedYrPtwReen5mQqnLXhtpj8kx+TFP/DWYwJ69xt57oqdAtm3DJx3
WyFFZc/T9UHlnZVkyEWX6odoEudue66j3FFFZ4MSAxJStOCrxXCweVgNGfZz
WPE6r28PD3n0VGCy3xvAYf4Dzk0LU3zUETdXp85i3eddtx3TtHI8KXuAzaa9
eIo3w1+4iLpKERWrL4vj9JYTjF9PUSQ+wieq2fHBL0GywzSrwYigoSKJ1izd
XI+4PKnMp7wKWx7c7TlXYnq9yK4N4rQ6tpr7FcHHgj6wDBP4Hq84zI8NOdEc
ctWjNr9308FTWzN6nNHlAqIkMCwQfH5PkHbuHfXvTBnEs6R26ELmZ3GJuKhA
un2iEx60+RQcKZ8rtsPaRr9xA/AAr936hwNaLmg0AhZVihzPfa9MIiUOjGe1
lZ/cobVU1v4sSM3k8tCNCVosFhezHVyZXHRA3GMnUjXzVNA19nf2GMgb8VFY
ovgnqyEkFwU8TASsfAhJ2hFV0OUFiO3fZkflW9Xv7YclKIEvwn1+ZzeA1Tla
xuUCbG/9Mkji37BpZ2Hn8ziju4RW6kQon2qiwP0aw5XJtEMlCWhByniO6wQp
bm9++C5SR79F2PjxazaCeGXUb+DyaKIRafyT6kWgGYBbuu1Heacw4/sI6a99
8+qDGGWL4vMEukLcTFDxRWc0vj/jlLOMzGaJse+sp3pIEbvnTHIvEEcG4Dzf
KEi+2TeMPWv1eJ39B0hm91Dkmg6fRMDafTh37MkxHVBg63BhaXw6BgKt0y8M
xXN2AJ8V7lSOkwGNQCVC6nayl5crSEcU6VO9J/a5XhLbTxu9HFx+Z19EZEaC
uCSuyABi+piM3+WT4mfe5j/ZeVo4k1bo02Sqt9G6PlGjRF7xjV0+Xqkzh50D
vG3PGlhyquvkYUr6RjtuX/yuVFITi9EgkAYHgu9OoFzyGBxkXSs4X4iiHA7E
9SECtj7enyzvbwtgYW/qKbNi+dHiSDyrzJOBiXAkV4zEiUf0R3VVVaMgF/0j
83VIRf0SP4uBT+3mv16+27ZDL2zhqMsIij2y70TVvbGy1UPa3Rh7ho2aYAbD
c1ocC5ysIeGaByR/nQVAxWR1ckjgDFhn4uLfhTOh1kgpd5OKrPBpWVEFS3E2
XgYy3jmEP96pW9lctGj0FepzZq5SNvMS67JKeAzcTAQac21VaFXqBmwm7gGM
yuP5+LGhOoDoRsx/RoYGpNUeuAWNfG655p+td53ADCRXmLwR+wulC9TaBzY0
jQOi4CSjhrzw3gDPeacga/eEKja+XlTgkbpKgMmc1KfCGV2BQPLhbCg4+w8V
EK8Fj3zsHcp+bUuB0y4s8HLP34mNKxGZ5qqIQwVSSeJAq06MnnzjN7kvfiZ8
eoxiaip+wbM8J4Y1oScaR3Rf6wSJsdO31bB54MToQSxWq7zFipaRJl3kUI3j
SxVYP0L09XFPD+TkDukRpULOkArHucknUCaSyMmERAJZaOkn3lznlD04xrVi
bPJLDUFZZZ3/8zkbIwuv4fSuQvXqQq3RTmraU/UJXD2lzoweDU1dOHwV+wC0
x4MEe4hcpE3YJkgttAXR9m8jPom07Sxw3HVwrXiW8YNuirFFBn8DrfA9y0HH
7Faob75Tv4ejE5G8WmV9fAf56A0L+TE+YQvewYf1dVlin/HcP3YAE9bXU8i1
J40h20EDWMaOPoEEoE801CaRSRHmF8wQQxcRMgz6/KblxCWmbAWlxmDWeE3I
q4lX51nHmnoNMZ3aaR/m+qOwIKpxXtXwEi2RjK3XFtQrQ4vhZrrJ8rK7Dvle
8UZ9nw167gntDETGORa4+dXOF3qeJ8RnCT7efL9nOzhh+eaSQsx1e0alzlL2
QyPIg0csE/wNsPdQgDrVaX04GHTQA8YR31FXZeOiZSgOX9LSg13X6Bt4kY3m
2A64UoRZOxVDzKhVHXDPX3+iZhS+54hbn909G9Qvf8jBz72NV+Yzg1MQJ9dJ
DbALz1ZVDKXiv++2YudWF82OYJbWCLrZSAf5dQ3mCJ9IeZ+/3AhXP99G7coL
4lD5q3UMCRRuMdc7x+BjCS/gHZm4vNIirolPtFYc8PooBFtNSsINRqMQWqgk
RHt7UC47/DLyWoaHIzmfEEbCcPNRZcinaLoLiPqevOQbOQjvKQ3F2RuKNxd7
/zYnVvY+sK1IdiWKba4Km5rAJpKBZlS7l5R0OYk5T3gvlPmrTPJifvkIoacC
VMvrvApZuIUo1Pz4g8sLX3OOSb7fk5JaKhXJoQx3z7g8ewRXeK9EDqi0lkN0
rGudz5MhwYLW+34F90NEwgp4wQALWyGeAd9Cyg+SoemQhFG5m9H62pjonl4x
FIgKpIchT3iJ5FcCzkNVLTP75hd5+4shUqsUrC50TMi+93qEMQ7cLz70AXCx
L8PcbD7SSgTsS4HcRKK920oZdxgPv5IeZiBZ2ihN/RZTtYZGuBIrwVA9POQl
wYja73bit5dy8PZvcR7FGwitlFJB6lUu/PeFCoXvjNkkO2j9cc3z/vRp3MZ7
vIb3FmlDOAlCYVK3tL0L6DkOCRAyGGMeLs5am92pTDLUjXA/q4LiCq30t6Ei
j6ae51o5esUxIxyO/pHyF45vNZ8ZP80YetBzBFnoab5nDFL9QAfL7EwaPAms
otLdpz/dw1pKgz/kF+Q0kqR55nPyWtlKrChOYr9dQTcyMDIwolllVY2/rmTz
YhXU3z34fbB1hiZve3II78BIVmBKpKZlX94rOYgG0fdU6VDTg9suangZLeW9
ImfHLiCqu/BvLcAwcJmFJFr+qZO4GfiR7ef4/Gx5VfJpiUfidLZld3eZEKBI
mpABofQ3RfHrJviQgCY994Bby4nbiRhN7kZuR2vRrKrXXTK/FGhcIsw3t6FW
qDfrhTHFDSO6SsI8EUFD3VTonJRo6yZsx4BohU6iyHECftjoAW0iTUrhSo2x
yOX2Zvpfb3NhcEYzGJEpqvSkU0uAWdFOvWqvZ2SX6emyTLSEZI5mzNSguxdZ
jJKIJppugP0vjJ4ZzJzjGZSoTyatzhIw/NbL6RMN8PiaxlD2wGaSwaZi0sFh
4NXOQetpg1BuEvxc2oMjG7miIzfB5S6b/NV/HjaY3Jmfc9FpVdVbii6t7wWJ
D9EeX91huRYNlZLjWIoO6krioePq30EYRKT2NLTnS2IwlkAA5Zaqdl1bd4hj
mMc8SwCLx0enGCLR/6qM1p7KTN3mOiOo94Cw5+YpX5jjmULCe27XzNhA3mn/
1gsBFj9eoHD8nZ4hE1U04sxZXBnosmOAHUgpqi10JoQxkXFpSCv9Ep/MDbA+
GtnX0fDZp+cFWOX0iij8DfznPiQC3hzQe01f8zE/xOZecYCWgfC4o9ivgsBX
jUcsA6DPnUw2AMTU3IpZkIWJJfYa6t6hxQrasgHpTUoRnxHgJMiGHsRTF1an
PC4kRaWhSFwZQj1ZEVCr2nNnvOhMMEtWi0d9MNaSGitZv3ztVUwrcXFFT4b/
7oXOpmAG4TmGWLLxxE+JNiCFu1RvIqvo5DJadkQHDgoX7Q3zzCC2qMygGx0M
cFWzS7TtoG255IRCsbdNuxQdvxBI1nL+V4eFZ/sLm4ifBtq50sq909M4sLWd
IgM4ttstCOW8uthUylnDfeXjbK2D1gZ2qZ5MlGieAfDpckpkytrrcMXB9xh4
zMlww+ILwK70B1PPACUKwvSJhG/665ngTZbIupVAAgFAk0ckpGr7rnSyCErY
0/IRRpvcUbr/LkslQYKDOreVtZvT9GWfWsLiQCeHY23sLREe03RJHf5Lf6NX
mWpQKbe9ab2R9vbxZWHRG7Bu0f6LAmUdvkFMWkW0wJbngvi5peA0a2izu6JR
K2ipXv/mUJ8rPo2ruT0cjBK49iOpb5lzzNV2RkSqsyvrflF6ks9/+tGYBaZw
gJyPuOx+lFObq0uRSKkkqIy5258eaBaYMHvVwTKuch2zFR8Nl/FaKeIxSR8r
tTFwb0M6eYsN5BEMvoGt+2Lm48KOxPCAnEeRzrZoW6cjmDPFCQmzyVQPVd8e
/SijI5A/65EDkAqWg7JElS6hgxvgFvK+md4g9yaAr0guZV4kCFODjxyaeXS2
bfkDajb19svPEHC9EC6Z1BfCjL6Fwe/liJIrlVVO9Stoq1+pim5X/x26WIws
vkwDZqess8jdZFz+p0LhCzXhSAQw9mznzMPgiYloI+ECW+IYsvGrHItJEvxI
U6uTgxjvfoeaO5/dNaSnMUw18xssptGeb3MkeY9AcNqcTxe8WGyllSEK6N1R
aekm5ja0ePlYWNeYU4olzSui84vSehzgFGidAEcLxswQ8CTaNnbyBqz1Xm5o
AkiPNMKHFkxRrFYXE9CATg4kTlkovk5DBPgYZ6jDsy1TXU5maNzkOmSUEFey
U6o0fFfzpTLpEVfolP8/KTR5ibQGiNgcPhq2CD1uP2IPsU1xszg3OtPo/Pb+
Ksp42QpSa7n5Q2phavmAH3hGPrp0Htru5pBL5iauBimpgjMBelD3FGpAZfN1
WgiYWVlZBXceVUKInNgytXOgDuHFCmGUeyITucWk3BoqudB85JfBmbGK09Cj
SYCP5jeJCkABMSYIA9eeouxI1q8QwIWRa/wbMhZTe2F4ITI0WM7CKnEYS0J1
x/BWADrDKVM6XoNVlc5W/0RxQOm8+bpAPljC6sIuFhQIhtp00vX3OzHV/iJM
lhsqUcUF+V7J7OumlDTTBqD9SXgKZU4AeIg/TuqZ4njyTa+VrggSD2ZtXGBY
uz8zONc/cdzMchow9qDIC4nwRenivbJfQdSb6b2I+EYaXs7TtE/5rzNRxPeJ
/yIvFtemOtEK3newjxulp5WplvpMdSP2NxRm9abpfAAddjU9vkrootYqH6vV
CrDKwIlLRlu9M5+uryRYoVd5Z/eip8PtGWCO1o4tmBST/6t0q39+iSSAZX75
t2dYpIWhZJhMn7hQZG3rE8B+Q9vjNrPjex6Q0QxxZH/V1bnW1pqQjChEyc20
eNA1YQPnw1lPk6Opm4pNgCaJy6f6ITyvIazqeotPHJSRUTkAuON0aY3D7D7W
j4dVt6KRaqFuJ4KHCnhnEz8oJK2HxGLSHY630nzG2DZuR0oYTU+YwWQyBGyp
BFddIgLV9ZugUczTtGVUQLq4xx9IAF2YUiaYcw7Zl8DdceRKQgPZQJIYCfCr
6OsWkOTculXDkKy3/jthk5RNAX9LKUam1liyx3yygtMPOoBHM4f6wRfOz58K
XEuOdnpOIQPvBmAe0l3lSbxLhvCINXAnlkfA0GjayPJODakpjw1ug9nI3Qik
fMus3uiHWbZC+KvEyGhvwxSHf14ak0MTGEBovGdBAKz/lg0OQnZQdVsujlha
LbmElMHRurcCW1GUdUJm9+tWZSlO6suQbr9w4d5iYNvoi1mVkT4Msp3Nuvcz
XHWICFqfyHZrn4ow2bz/Z2K0WdRTQ9dEmqpCu1BnwmCoBos6xKg3ECeiPjXC
5G8cQRpSSaYo7xMKWiT+qWVKexKI8JRuzEAW50/SglvO8Uw3emnxS+jijSsX
M6MeiJqQxU6oFA8X9sufPQnpfcJ7ku96F1aVKPpVAxLhnpz727M3zloAoPUf
dwv/v7gSJlv/I37vHUi1m8969f9h2KQzck1lhbOPWREzVy0d601nnb5SrBTk
qhlRRiI7rdMQAueRmvBMJe225a2M3KzSbH18308Fc1oE0fSRPe4+l0Hx2wIg
WNmk8e5tvI43ImA+yteTAwLMe4BEpRd1OHGAePc4gKDe0xWEKGz8ZjpFBDPn
bQ4eXB5aeqEXHCnWpv9I94vUQ2+rHjXB/EGoHJpcffY4tPtrHK+6OyaeCc4U
pRRxrRNt5s7nk4z6xt6nyV9m8LmPwQ3phR9SqDpuYz8ItQR2+b7UsOUZmItL
5lVGce8v+R5lGSe6vIXjQ8r5RrMmj8int3e949ixU/x6ulh3gkGOxlWmD7me
SCUGfiBDkJwdpAsgdGwKitC1SGDrRPpjXXmp3HL9idEgkiuu3+yOw73e0IiH
j1+LA6J8t7mYjGXLd0iCBHRmeyzHOAUqEHCUQBY9rSnf1/nFCx1y3KDaV1lQ
u8/u2NGsRnEwnOxkv9A/d3C0eLjalwNwdSWG5uYb/khpasbIrbTlebXnGK0O
pV8j83QvLBm3WVnXijFmyQkJHIS1sv3mqJJ01aqOb9+hwKGNkbrENT3FdxeD
nkCCNBiAaFMJXfkFdYN6aMnIkHWJVMGJHXZJ/I3Bh+s9XVLsGhhEiFOLL3QB
pWxJml+QQtH/Di+VrwdZTn7pgDxzK9KrZKkqqwzJpe2bmTEdfpjSWZiqSsoE
aMRCOU6H80HhtCus3Slb/3/Cfvubs8DFsdZB5cfPN/Cqarc57kl6ayI5Erdk
ICZO+f0jXMHGMWv6y0zBgTpcDRSUVc3dMzx1Ka7b1xc2M1Krj/ZUMkcCePnj
vRsla8CnELAqlE+9eBhv8/FRd5OjGTkAhLsGmwxoKkJFBqSQCuBFfcrDVp6W
rWnIi+o32SISpQySepZzDZgyCZTBj4M0fCLS79b/R9jkejobV2U6CUOfZwDZ
UaSYgZ9m4iOaAMdXHyOP7s7Gwo53Pg8d/Q4Zf4z4CVhYWC2cugO1iFUGp6Ig
hsI/1VReLYfy79OK8YM73YrMLzh3KiBh9aIayu2pgXxmhJNz9s+suGf+OKqK
HY1vtlLNziBMsGbpVIf9n2VBX0tgVPIdmjnPLVPRzP1FxG0Qszk+2Spk+ADf
iU0SaK4FWAg07XhCG7LKiYMj/MyV72BxuiKSOLTWf1K/WMRO4I6VUH44CuzW
qrnpTPgf+lRsq6wEEB6QmJGHjUC8ayrqNuqvgGPGtACF2MkkwaggGdXtYKK1
EaOk6Ty03YB/Nirb1aO+L9UMHVjINN8h5co7Jy/SG2k1mzMP9Snq/NgWdctl
0UWTBmxH0BopTA4HtQNp4lkrX1ctHN8yw+Eemr4pbERkvbi7dB8a7lYdDudS
Xb9PvEKxiBTkoAQcZTU2KuYmRZVutT1O1JGr5BtzVWCH3YmtlP4RyABfxEAr
U+MazO5Qn1WCtIjhzIOztwcyIT1bv6b/1HIofEqJfurIvKNMDAztXns0/rg8
gFjjx5PyJslKk6crvHXG0y0sSCepODoL2wrbt0aSXAOIJk/VeW/Un7S8znbh
ZZyIEy/pOEVjbewOnZuFjW/8ypm8I614Jwupl9aqLdJLHX08kq6+UQokWm6z
Gkx6TD3PfO9qknz8FuB7be8vt1S6k8pFVHovHgCJnhGcYyxmGSLRgHNY3G0k
NVzjojNxNaLr9FyZNZKDi5px5tQqn7OGpAquBvSBQykyfwnM6grsMqrQ5n+c
/uWLOqRe6xT607PTx24ca2q6POSoP7meOIEI3enEsoogTYLlbA3VLAfvd3VX
vDjyNGBYXQjGSAPZWIZtCbHss0I9Q4aHde2IsJboC8yTcp87W4ruVT2dyyNN
9SLRATE3dK7LRBOu6clx3y8H77Ov0rSOAeQnICj4V1oJHf6sPnzWjiHzsbA0
NJkdBvE/+8X78kFvd04Qo2b0w/UqB5EZKJG5URixRBmug4ggwrQTs5w8pKSK
iqBWz6zDMGjClgPYYNr9eQOFw8rIZPLswKeYAJjYhPIw/YhL4VkItaOVczzK
kC+/9A7RAJwSE9FSQdQPfQuQQBVpuU88URzhp/zqMCs875xDOU7aCgA7ieC7
UqUNz+1ckcsmdd77EjsRqatZAc5+g5aJIpS2xRGFw7tDBD5+1PMBXU0sYRux
73pAubx8O0wll3nruqKUXbnIRXXGf48fHoBsXlXMw4wyfp4QMQA7bmkdKjKN
nNwpGdCxPa+rNNdU9suXGFkP5yi1ix5tFH3e/ah1IfH7CiPHhnFzKyHgxIAk
A9fM9IZx1BCTYwJe8cbtZnwUwOzCnzFyurhJsPoe4RuUjW5OwULie9bx9oZu
aey7wh+h7CTyMQxBJakVj8oPt+hszhzg6vOmjnzHuI9o7ikCpZMMLLYTVI8G
DA2V9G6ma5FePMn+VfoBAcD91Rmj1ozRCZMDpzVXjGifkRjFqp5+g4vccu2Y
QTagqyoa1zvIvdruJHUOHKyCzp1F+OmuSZqcutyKq3xnAPqhGF91vABehbn/
dMY3mbBWDr7HBWV9qjsPUf+tGDEvpqWBFQY7QDlcBkBryolUf69SQgvQX53Z
ONcirPz9RrXXog9ufGQoNmk56QyLpnzIvsRHg1qCMS5s4nie73D4uAkaMydu
rcRykaGmwye2ncdQI9HThy+ZrWBAEGemRPrMiLUULzUFp41xSwloaWyqQB6x
oCzAda4WA44BCj8orr+rHiBpnoPcL0m33e14hGJDD7k+0N15a1YfGVhOOFZe
UKEnkTHRhhWJZsieLLxT+lWIKeK2Eg07tROtbdz6b0XZ8dZ2ZwY1WrseHJVa
22vph/TPhyoBXJZr3kKQtgxv3UkQ4iWChrjOOhKTu9L8ntMmmjf2LV00M1w7
E6OfCtdy94GybqnVn8jHdx/VrznoOkwNdQX6+NQtp/nBaQ1XOGcdM4l9cKnV
K/eWT8uQGTPvWPZkFjEURoxaATmisYqX2GUZVwP22FiNtYhvPyLS0Xx6I7Qx
A3hyeZXBd8xJWTXyfHgwCVrP2l6g0ukNxcxm/uePHeB/1a5Tz2q2iIv8ii91
uTqQDZ4lCHqDuDVtwCED+ffMC5TVeasCZUEs5N9fAqjVnPOkCRgunJSwoPhc
WYOGAbdAwq8BrcJQacgKoBmAJwA5AutsaiGo0Ued6YyYU+qQyBEx2klruA/0
45z3+g//T7ipc85rZsG850imqche6DolOk76qWNUhmw9Nj8jsw0/urUUUz5p
7pVC/59VPZ7YnVGk/E2iML7PrZ/Y6gudcEPhY79GhX4hXQJYCmRW0VzxJKiO
RSKewP+N7B/NCIw52gSx+MwuiilkJP5lqVGTFUQzliaDoWL5ruqT0ZYCbLhC
awM01SVglJaCRs/Bl1QwtfrYUwTdCoA83Y4RUtp0YZ+OAeU8RroTDLc6A1DZ
dmB8IuMICdutfRaiBlwJS39yoJv/E0E+8n9QQCCGjNJVxOCbMOKB11iHUL/G
vqFcX+nEYpWwELQ7zzwAR70pp47zJIm6yrxnNafwPK6v5Rcn4JMYlXsIAicu
Rv4T9PoGAH6G1muR1JP3nLHjNiMKElzEB98JKvYEnYHuRuRf61eOE9eWO9Gz
9gapjK0tZf0tJTXEVr281EOcs7jXalxquZOLkxC8lO8/t3XyiF1eDhQesJxp
JymWnRU5kXYSzUWLYYJeMi3rYQ4J2XcqQzISwBJe6NwRPbKaTYyVcpQrlTZb
gxDzdovCuSOFzNFT1I/ZE8hBPW4GWb7CTatyTGoYWqBZyHpTlCD02rBHCP3s
8wo3vOWHKzmHp612WTkKMDP2I/IVjYxrP6+kLaIB4PUsvajNZHBwEXceVKgn
s4a3hwOVxkq+IqgUT+SXU0OwIctbDFDTUB2hPYDx12xjO6c0a+DUL15aZWTF
fHE5oZCyjsq3AmjKjPR1N93KQcsOHWLfoADa28Zu4SBsxfh5rmxPUOwpOAYK
hUDvmMB1W85JtgfcZlWhxwVl44iOxU0YVzDLB6vzcQt001xwLLUcWlOvbM1u
wEAvvPDpe2l1vM1zFsRUUFUqXJ4WzXul82YJm5BcynYyC6CYv0vLPJ2rYu3z
HcZiZBO9KSYkeMlw9RVB8bVXF7VLG9c0p1vTdJ+NF6QqXFS6T2tKKK6/quTj
r4W3a6gDOBdA8G7lVu6oluH1Srn128woXfun5MZI7jUl1p+rzY/z+TDvQJUf
KaFqMfw6fd6RrgE2nIOkJLBu0rNDISuzNBI//o/1cRXvhVIwEJfhiM4E6dI9
CShn81Xy+WXs6C+QL+qTM20rUqXhK8AGkCIh04wXd/O4GZ+JR7+5I56oPgh6
QxImS0lu1jByl4JLveaH3jJ1cic97vJgyKKpn+/SQcLQX57xg++5vUF9T+6A
9KemUL05esqVm83xygS3tP57v0JpZwZqlo7GNGGANBdVm8LchzgAMwhI+6N3
nKwJBkZ2kKSFcGc+KKXxN6hcLeczd0Nym8Cv8g1WTRnhYlG7cryj7vJNH5Ea
Tzi0vR0IUHfA0shy+5vjhhspZT+I67fpId/v5H88jHm0BHP2dKwGgL53c22A
ZHiDZw6U8OQwpKUi6Llu1eC22s8e4v/Y4TFgX/8XjlZQvHOdJXOlyoP8by3K
0cEKaGDMViQ+PoahfeNzKt1ZGFPrI0XmMkqzr84aqpNnpq90EpgI8tVvGfUu
xLV98+LCoWKNrrfEdvnpgE9jGr5raxPKCYvpzstru1Hd/r8vApemzQwGHXTk
55tbWI9hcI6od+tOD1r+j/C9wK9ePxD+4uZYY4Tfsjzbl9pcDLSPHujI+Ndv
ZJjY9qwl7aQKxoRYwxyxtuSeejjVr6kmY+2XN4aQvWxPMT+l2KyiedzkzfKU
RXq7eZAmoqaa2xTMP+qly5LlAcYgSFBvPfZGPTJZo89aUATrz0VTSwD91chw
C/z6E/6n+wVZXvmoqAxiJ3PvsCLhIb8eWgAZtG5cLs/z0dMyh0AAH8m9GGsj
5uhsBAGyiAqvofeX5kfDMU3q3ZiJi/rLEVzCU0GAMhizLLCOzCn2ATwA2ndo
oUsW09f8mShLS84I5A4G4mGqk9zhRWII7119LbC3Ea8QGnngoHtBfRRdcuzF
1g4HsB0JrxYUdJMsbDAMQqgBCxLZGdGMyOiC8wJhosyFMeXImupQliNxl/Yd
uIjrgkVmEPJRPYnWPMf3RWC0kicv+CkocpDrXVz0Pt0mY0JEDffG2WxcDOph
TSXV8ylOMegYGvoGsbdZe3DeF8s4cWjwwadeWVOuSVFy532dJVsh3mxeXM/g
YVL9WouubdbzWE+2Fn0PD2dPB4K5hTpE+EoF1w4xTPp/OVck4uvX1fhn8oFF
FacdGjSKKDY+DrlzHxAOOLm/0P/shqY6sLIo3Ai/n8s0a8mm2kEPKPAH9vj/
yL2n6R+IrabD5MmuDVgPJeRF405xQvNq6EjpKDGuO6QPofpc+EFHdVdfmW+v
rXgo8Bd+thWDH8mJbIUJRWe4jigOlS3aR1wqQjMP7ufeAbEZSq7VjWpETend
84aO4cbA0ix3ppDs1VOYgaCt0G68wNwL0+ZXzM2qGoqPoBN37H2fxUTZqjps
V5RvkelZ2ABBqw9EYEHb2yIXtEXkhNaobNWsMcZveVS51Q91sw2K2mWTivhd
vgr/5rLzBirD6C3lX21dUGpm25ovqtsefJFHo6BicEhZhSKbE0zeieIsKoda
C9jEJ+ayonW9UkgZf6PMxWk99bt6a7XH9oJi3eQEg3+afOBhzj36vwlczjAo
Ju2ZPwrnAgE829NZH8Ce/x2jchul1j3Tx8nXh1nb2Ht2xpZjVuIoqDwbcG2h
VwGND/4JNFoxLJRjEB92iRuNeI5ZWcgKyHYWUNUJsmZNSRLkBN+RiwNP0DjG
Fzu1b1Gkq7EybNB4QEWaCyNOFRW/1pDhkz+nXTl5PGfjVH6mPRrmHx+kQ47E
WytI53m8NrjeE6Mc6P3SjNiLTqVKcj7TgIbR3hntBYjhdJnYUorOd4p2nyuZ
vfiZgLsZTjLZPFjMdMJDAyFcZLvnmHnyQMSaTm8vL0qlEpONFQIeBahwvube
Dy5SFo2Txhbma5c5oGZcRqkzfYqLbjUrSsoLpE/2xytUNQa2BEzyfqrWJtj3
r33mXX1UoOZnPHyvrKEHYE/kY1a16efkkUvv9TdRau1zrYE+FI5vruai3CkD
QXSlU4RWAtoDErs9/7kHqhPBVDryyuP8ppWzFjQ1YX1za6yOtjErK4V1xkCv
BGzIF8rbENYKDZTg0ienZHnaocNhReK7oFn93qCD1dIT0CpSgThJq4kIFWqK
47r+cWqTuxN2d/WevJI7anBOjtiMIAnbqjzED8IdY5EE7cSIQY1Hxd1+H2IW
3bqhD5EtUQGaSuXOS3KAgrI8AZ9QWjZfpWhOm/ARbc8Mqk1Aw3vWSavnAg2m
sVyfaxNU42YQCSLacIiCGWLCfWYztvmAZ7lLA27kprJtA0LfTz3qqYEzX8Th
5eF33PsA3lZ9AgMVqoWyeGfHtgp3BVdve+qaDGHHfc9jLj3Gb8odRs3nL13i
ZFZkNBnGeTevTNBxZr+novwaSdx8QbA+w7bgSvWOYaFu/qXfvBPu7UETGN2f
v9WC6sikBQjZLnyN9gWjqgrMIhPz3KI6o7mj4qRT75kUt90GoVP4bQVZm9SI
tSNVKzIZWDKDSGL2+U1hD+XHok7VWnmSLPkClVnxKo7NExV7airH/cbUMdBa
gyTpYo5J3D5MhCKEYOK+csf92VrfI9J77KUjmThc03xlGw6//eumtW5updFp
qKcVMMjvXDNDBnENTrPv7ekkr/wdP/TUiw3r0BiJP7qWvkLqRLsrQFZtysoZ
Gpw2zv6xx0aMjBsKWlGvEITMDg9cEuswyNpdalOAeBpRbEdyUQrKrERvtuBv
R64nt/UpspuJ1n8iJgd4FYA3YXgX4ddloUJZ67niRs2Ah6FyDgqu41e8RDIU
NJEVk7Cpa0uSTqspMiVta2L1X2MJ61bU3WEARwHaT7PvjSaDdLrrZsR62tL8
MCWIvtnRFfAJBzFfZ+8NnaBvJrfLrxPG7PNOMkrsDkSE7KVu0aKViJvJFJJq
OaY5/NZq9Rhp5KdQXm9cal6kcSbl6klBijHqsdyOCjLfpS7SHZbS57AYnZ1R
5rpvIXq59EMI9AQA/YYOd7ZFNRfhUjmR9Ibu/r9CS32eo+qAYyj3jhDtHBEt
sYU0b9BSBVIChJovj0auoMj99kLe9krcWA45dagV16beQDyOjMwqQNj6th4p
vDlTK7fLc6QwomDLLVsbqN3pVnXMRMikcKYCsgleR1aq7QjLeRjCeP7SRnC3
xpyTLgaYxDUo/pgAlrhpf28sWvNUDXF7DN7x2tc8tDVlU1Zg313hhThLLmay
zsOwleT+WfiYuTGTeUI9AvpcmzJmPEMtYYIpuEqvoeVfu4/GYJs4nBL1pIyv
7tO4NQg0r92qRTetGA6b63XCt17BkdqE1nUqzSF0hrsKzLJtvay+aJ8M3B0X
wjEyEJZZ5CtWhfRGeIC12vAUbKlJrm20pmyn0grL+aTbPlCngVlLtk9I0ewt
47uB9IeABAdEd/3JFTDZndQc796NO99xRrQYLbtN0f2SUND+zelDyAsPOc0i
1HtOEl8IW4RFwMcC8hNlMWUT6rx8XTm/K/kFd2aTKWIA+fsuAP8lx6+GnCfF
6t/XjZa6opQZrvSskJzFhQwUweZU/qlQAFJjl0ZdvdyYoBOrQ1GSiJNUKTNw
VdikLPUSEWALUSJoYXdvssGMHDfO1nHEhHYc1Q8rNocwjp2jQDlMXUhWQP8a
rT+y5jua0jIeXhl1ckkaDCEru+1m1tLJUVq8aaBflemiQszITB8yw2wl8OOS
YO/m7r8aDTfkUqW9steWtEphHoy55Sqc2H+41qe0V6MSyU4DSmBL66LhUsOK
qEsEDXexsa9nIn6OSQgdYW+4Yt6TZmx2SVsDADEP3aMTK9AdQlhIWk/lyciU
8R/oqUwvv5LIq23dXYeKVAbEEhQo8zCDxZCkgHpcHFcXOS3+FZFT10KzYfgc
ZIIJ0OyM0yr4M/C/MznigltiWMUndBtzEeRI/qRbpD7/ONOe1uYyfBlPWUe+
XQJxqpJd80OfqMF50EwspWDZhKPGxStcbhjjchHeDgz68FF3CD3ozVp64e5V
9H63C2iEc9XE61j6EdCrcwEwl2jc9YVQgac6gDZ/fU68Zk/GgW5CnDuV+MSF
Tk2WnXSAnrcFTfIs6iDYOZHUpRaRhBX9DTw5wMcDodl+TvgeJHvE6tNKP46+
IIrHVjyt8Edrj8rsWGoREz3DKfRU4FQSp2Df/hfaVxdVd5QbFPXNks0rnGsp
7Ni7FxVGooC/hQHgbDZgHElJ2X5fGdiqbWtt4soHdM6OSk/3ed/FB1gsvZ7K
fsViaBwN6qUKvTkpXKeqeBEgIOVxMzlPBQrPVmZcgfLg8R4nFra1qscfaEaU
2vGjbo3Z1xNZWGFym6btrsAtB+sGhUEtedsJV1N8eMtfPpHfgzliIFYpnB++
Zvq43bmx+HPzyLNn2R6tohyJWkynBw2NVLTbA08nAU84b+Z4mbawfik1A65r
59oY0Al4Y3X1QJaNbnk9dPAsEKsRgFnOEMraFYHiv7PqH3OOQYl6sq0cNyPf
T3WLrPKSBH3DReYWnR1iyBlcS/53FYM2ilDnNbTCaKVS4q1RmTVZzK1aebXD
fwjSM+aqYK6QtSFcoqJypLYauoOrkRQrBLDYH6mQ1cEDmb/QYH4vn9HxcuhF
wsw1jauWvFWGcocqxbEhLNxtkG+a2bog+fxQ9gojeEZsr37wusx3Uy3sI6JG
+ig7x9pJavq+Py8n7xLhLXh4ZTWlcGCbqenIrr2/9T3Vsjy2WhGaGrjoHLTk
/toitKt6q4TlJNVvxtwsxUhijok1ZX6o9KuS/m7d1ziFjUqmTs9VMkTE/tFh
k6kw08ERGT4+oTExjz9zgKo8VVKo2a2eGPE7VgH/k+0511lplp2q31fj4eWI
h3SLLsZVIsOOQDePWgu4HA1GgJJH0a9q6JWgjtnnBdEFul96bfRArkuDrkWO
WloLdObKuCSyImuXj4i7TS3fa6oj9CIIbt0+TFbvKBIWlFfVcWmFqc7vynAr
hZ3teQpazL4aSAHBEy+r6QLCWSo6zKoY9O5TmVrMkl07IKIxEGATbGg4wzRM
YoI0tNOHX4nWCX/oOO5EpG0xyemgSGUFcRA8iBMTszp7jdDwE9cLRgEEZemh
Y4h0hj55emBtYeKP31DPs1ibAx8EvSH4IrLAUbiUBcPwZF+GvXwv+lItnwFg
v3kB3K99IBu/0UDYBzZJQb+JeZ5Oqrkpu0+8YWKaFZPtN8CyHL3DSSyw8rLI
HqtRWjQ+P6990ag/hktKSYLDmUXhp4Aa3tqAufeW6dwb9G5pdreCj7e+W7e0
qd+Elk4XGvGSALz5bL2xzVxoY+kAm3SUYkhKjJmc5v3zVo/rwiRxfj11JX6T
BNy5hvKaxRzqTA7VLifh9NiRfMj6dotWKQ+E6hdEifcSYI0NI1Gr5uTE0hhP
f0IWdZOs6opNw9wuEeXVtvTgzB/5L0Xo07nszuCfwfggV07ks+fLtzOU6vLv
OcSlfplKC/jioQk6pFRpsJmRTT4QCHE86di3IwmleFrnmssdjvkvL8Fg9R5D
Sx6M7cZAn8rD55S4a/z8HKWoMi79aRzG/bolmUjIl81IAdis/VCHmxAmsU0a
KKA22K/W/Lv2LkwWQ43mEYUtk6L1DcMwYIOkHEhZPy4PnDiyPZVufmeZxO13
ZT11SDr5xL9PLocEU+BIBMdE8e/Ck+tsIIzN5tiYUeg8o/leIdlQfAPxmO2k
EMYzdaqMV57p55LwUGYAVnZIdpBu1KFpAmUOnmBoDkz0oLaLWwaeaV+X06bR
6/3PO9k44GuzW9CZ/uTfFFL/DVnauIoPVMyqSIKxQYflZDBEPPZUBJndNkTz
kapFou0aPnhzIUEOL/YW3GFz3yCibD9+qoto8RNM56PjfPLCYh8mDXtcBQN9
wgozeYUgb198ISR+A0R3VRlmo9g0lF7SkqjKIXwUItx9kJ18Nx3Y0uoSrwkG
wrT9og0nSxm00FRYedzMS2b3wYvbrd0bMl3RQcqtiJvKyuCCnKKuDorEscv8
zQS1ZgOU05aBL0bRgSr8rxCCKW1sz23b/VxsVDoosXTJ4sWBgbhqXVs5cW3T
tFr9N9Vghwd6ltDVlGRFxfmD5Yr2DB7QSAnJvfpay7wpXi8LkR7F7KD9C0JE
+ha5vYbkWu/YU1PY/RzAS5jPTKxryYAI4CRBdp13iwd++83H3V16YI9Alk6O
IzVZgDajpirnCqKp+hX6KMZtTyWb6gN0u3JXxrTtwlTHfL5V8kUa1HLYzISY
wWuWtf/WgZglIMqbkc6/3/QAaIYFAqBJ1OS07/rPBzpO6MxhI2MrTIB5IS91
2YIfkLkLy7mDSKnYzLE2h1nh+icN2zZAHY2Eby+o49KqFCK1cOSS/GrtgS/4
VdukV4U4RXPCaaJyQDvcSYoNSVOp9lafokcgObIN+c4QVQoWpWko3Ya+k07+
/rwbD/TqkFiqg1wXOOYxjMGlIDmgQsfjEIYq2zpNWace/9n3H0TG8tJ2Brw9
r+79IOQZD9sO1NCUjDMqX0G7S37Kss+uXgLc+mob9CxG3qxF+Semz9POQlW+
NZkJCmyfpM54oKgV9+KJJcLtT1T9W+Ja0RpO6KTJ1aj18W34CAL7gyWtu4qv
+a/haLGG/UJqTsMyBBDI96U83fDBQjlWFZIFAObTZxJcWcEWYK2KScpcwG3+
m3bGI7RRdjz1QGf8XdK7irb72zmPK78LerZ/CqzXUcPQBNtNz/9cUv+8yjkV
Nt/OkAIhe6ccN7POdYgfCfbd7wJnMes4p/8WFiI6V55NGlnYrZXSWx3eEL79
vogO6kTAgAGHohEuivyS87p1EJXDd397E/5n18e5osaYEteWFNcsxMLa6bgN
nDo7/BSzxCFGNmxtaJTkQqPdxhdb95af66gPcAAWAIh1gRdQqDdqqiBu4Q9k
6M7rv0RW+/xNgthGmtXlwcw4rgiiLmVY5nc00QyHG7spiv6Jp4PqyhYpkc/s
ilVSZevl9A0FUw+nHTBnJKSsIW4153hArj6VbZXR/AdXmVbz7+/K/GW4Yofs
+3vtrctrT9SyOg6BsYk+ynC4p5LF9p+6wmlnI+Cdf8weOHdjYoK6giRI4kwx
F8WlljiWqmdi/uOK7pplCVz9hAiQo0K8uKq7vuEcMtOUDLwohSlETcf4THjT
3X/Pfyzl5dGiRl9b+1Gc+Mva3c8w9mwZJWE2lV6p6IJ/clrX87Gd2yLxHfhE
S1L9FlVX/PG1n3CQPEDZuKm8Q2+HZLcIJnYLZhcdRNQczDf3pnMz/cJEU2y5
Yny7XkgbLxctMyij1ki9AjGqG2VZFJlCAphCtkLdqIDk7M6SinuWOZmDoM0e
CYWWZlQi2rErQuc/ocS7k9Uwvua2otMakSd5IzDyJXpyghqtEtCGlr5F2WO8
oSZpjqnPRYU9yNrBGZWK8YQQR2mQtoDFyWSvgObcXMo00AhI14Zl4CgOG0jv
LnKrHP1D1xWsLNAIyOzqCyI5lr462zJTJdIBadGmiEmhhpnAJrURbWfCPqYf
w/rT6LlrA20ut9hcX51m1wMWNyZY+GdtQH/ET0ZQBYD7JTkLTfo93fQJIzgg
Ql6j3cYgT3Q+QRTGH8sy7we9k3RjnuWx9g2Mma0yFUBYEACaj1P/k0f2WAxn
Jr31LKQNwtu7n7+vN7LGcc3SIgPaaVOtbLIvB2eW0VxvehwC31HrLog16xs2
myTIjHcNlxQH5P+Tpz+B8lEn/2wy+lrzeEyLhF4X4/09Ogc15BUSlkW06EbQ
Ux+x4k2QXGAAvpdVUNvVOwHZDL8yhGksRMqJOoos9O+YhW/FN+uyZtilB6QR
6vCkzmyE0tpVK69bCTtQl0+8HaAB0RfVhd9fatlS8RCGHFI17AW/72Q4KNfW
QmG9vOtm7tETH/obDRoDSeBKbf/SzA3TpNG01o4lQcHVjwLJq6sXBhBor9wR
ibXOAw/LbCGwDRpe7rrtz73RA23JCdTH7mkPawVmi94xWdK3JXwHAjC8ZTOs
2nEo/lK9kXml2s4iK7KI2hPfRfIKvZ/hnZdOB33kRn/8c98chYNGaD1P61fr
GdB1P5FL717p9FIgBB0k3azPIWIaFi9brm25aJfLljE0dHiYIkPmEgEMhb3J
TL2bKY7dP0nH4Ol4WohfVZssqJqePf1+UnROzR9HxDlmObZIBBPrtV7StKZU
ChgVs6et+ZuBNG+P8rT0svm1wctD9CxGseDHL5EsWcjHJtStfI8g8DkcO3FV
iYKYv4aCLv9dce59e/MOTWDNZst9cx4t/vj1TuZvMTrbKKmy0Ep5gI2OvUM8
fzWT4pR3iwRWXQboVMydW9MFWvAbKxWSA9/UWXDLGx+8TQteTqqGYxOeAwUi
TSxTLnxbfCPgxqK2geSOBoimGzbCO7Ji7e5l81DjDJUdsYBi7F8vK3gBa1BO
SSCx/ZoOUlyaw1DoBD+OEsehMqnHeUChgA+jzClUnQiO2b3FSLwHa9lQpc2m
vVD+1QrqCJiic0W6UBza6h/FF1iooGeCgVJT9/CyVtwpLgkrOCCpy2u8Ai08
+LrEAVVX8+eIILo3rIghrdh55UgXpcLa2yoDgy/+cHT982HwDhGf3ttB8EkD
qXdhrPZw/4GeZ+4F19AggeGhwro2aVLreWvcFnup9nMVGGO6Cndghtg/3eK9
N3VoD2fwTBqZbMQrYR1F8WG/QINc5hgDBw2r+psRxbRH1gxJQa+seHSqFc10
33E7H97IhP6JafLMIbzLxqG5kjwNfcIAMjJ3JE+wK61NElixYB430SKilpes
jclW/MCdPluY3ktNg2yuzvkbThFbPYjlhwK9UNWrMhl47EYJ2p48IGJlPu6h
+PLAP4X7NWLmw965aY4jcJe2oKfKVpvZOy7zLGvbZ0frnh6E7LV0gOIjt/n4
L1Hu9B+oli41PC+CdRrrFWlVHX/KcpZooK9avr/leVt/dyPpxaywdtBy8qx/
5+i5UEKbIJoPINSsxIBKCYO9koidUkLsqSuqStoVd4nPM1DYen0ZNUd55kxa
1VNHyzMWRtm0YnzlKrWD9NnrMsTPnJdfKQMMD1KLJQDakinGYSvrJfA9ibPP
oZ/VKVidFJ7bgNHT6aTkLuBxQ/Z9ufvlsJzYRgYiMZBrVwQ1ShufkX1BsqLv
Iane4Uk6OLG3PMoz0YqLr2mIfP3/FEMyupiRsFZKdV+IrMS4r+JoUL9bXkXW
kOm/Wbng8FCEY4JZlRv2BvHRvKNMq46kdfmQG+dite8uWVLhMbDHNz0cGJuc
msTSFTnbt30ZjGfbEFprNIKtDO6pPOtLLmfBvwSgOvr6LgmATUouZxNEvFkt
ulWyAJfoT3cM/wK1qEL6mvxQ67j5sL18FgWjvXO+A2ZZ48LWWox22fOcXKoY
FiIyIR/7wJCg1qGVVic/JARSqJv0/BXf9EPS0RW+pmUR8eD0mClAdim/mSfO
TxnqJ/PV6iMtbaTwGnLxkijHk817CZEIPFQWeTwFAUJgaHMxOVUI6o0lLHsF
jtKoEsI+I8sDRYfciIDb4kGR/d8KizBS9J2zS0eNlwu6rwN/K0SVISa9BRm4
RdIp92L86HdOzDOesWFo0gJOMMLCJsudHxZKT9iCucXWs14rOOmm7WRzLXWp
HZnf+/QsXa3RUn2c+SJ62JjRBkbPJ76f9xtWe2UOZnRP8uoELrmDL4/76iWm
jQgryRBBv66nEFcG6JoHnpVeCc1stC6LBwUSFOBYYq20griR/Dal3z1orObU
8sPxox8UOwO/z2sZvQFMS6FjfyEtVaZiw0qNv1bS4x1cv/LWCe1CN15Vl2N1
XkNy1kqzxUWHN/eM0qyGysHL/x30r40r17cGH3LImGvkdQNtWEue459hY83L
hfQzPQf1c1gY+NKqEUOOQDb14p/mVyZqJ9Lxx42tBIVacwblbXvyC3wa9v/e
fp4TFCfhv6cjeHSNvRL9yptEAhQA49hbfsv+zVOeiom1OxM9wrJn1D4w32Y/
KG0Kxdmbrk2wwhzqxwauj24+5zm4F5a52bzLLttBGmgTRH38Pdk6mSjTb6Ib
FaiTaYWJKzhixKTmjC/oyTLs3qhcLMnDENcf5dF8OYRLlerhq7XZDaF+PwvJ
zVa4oN2cwk1dFDggQ8Bh9YPT/Mr70MUFfBzl5/0oZuXYAXaz7ZfMwDghkSIf
y2X8Vb8YBLZ1IVz3b09A4o5Cmb+2pwUV6Uul7dfqC2lLTkYRK0zvn7w2wXHo
UfHvuKZLU0IYqd1xVH/lEKIkDoVVVGM9dtHj83QCq2SAyHHoKWEmILyJRQ1g
keWwEk5f3xp8Ve489dJ9VaU3kt/BcSo1LO4/JoZNAZ3KLpvrLJcdxrjlaumm
lrJ++XPQ3ov7/WdKmjiFq4MYs+zWQLz6lGFwmrMuC3WnE8CmOblSHBjIby9t
TrUo9AqDlUFa8BiOQmcXT9bjF4Y6rfT9CB+mAVbMbGLYvw975JmjPvZWzjer
UqLnu35y4tTujYHxVU0rY98XTmqqdedUT5qzwQ66zJWFSnd4bTzrZLnC0drx
4U0Ut/Cvli0x2/QvvCQCH5P0xRC9uZqQFQF2QNRbQ26j89yLc+u2Ews0BPcx
ERaxZkrMjgyR4RqPN3O8ggp0dqYSe6WZBXRaEm2zLEzhsOUe024lY/8S6wZ3
csMAadsO/zEafghVNH+oT/MwA8EkcANevBzlRvLCAtfaVffr90vDZK0LO0nd
io4UfqiQ0SHHa3+NPFZ1TWW+eMK80rI2NvmApvcwZxvXCWWMH6yr2Qq6kxWA
MupVYXMn/WnUdk6+ERrRzFDT9Z0+C6H74PEXhWjryc9ZVQzIENe3DdYjtgYo
Vsb6T/CAYzhrgtN02MOuSc5cYL8gS3qWP6rIvo4ioLBmLfZrUnYNohsZQUsl
gfv6nK1pp/ty+TrgMkzfQrgbZYFZURLqCbPOzCysqSPJ9QOVbmMfO6Vhr3ls
zMDZZknhJAxaWtJU+zwovZK8Bry5WMHhOQoFhyufl8lpHZuNHIE9VycX0kC4
kgaAIrBmw0qS/5IiUX6hUNkzYnmCwokuVRtbOvFdTYISx7x/UHsbuuhagLvC
+mt/Zt5c6T+D0LIritzfSBgl/7f4gd7IVee1e00qJt3M0HXBY/ceOA4dt1kI
Dm5sTDFuXD8snBop6En5Y65QCzeiU6xVyBMwMjpolEI9nJ78WQiRQioMPGc0
bUF+WE+VTu+IRQHtUIe32rKFqoMua0aoqd5Gfi2Fiugcyqh9d5HQryIl921c
M93k684BuvdFBN3hU1i9eE22t4TEldnFhwjyR6WXi5rLUnikV4dQ0s9S58MZ
6HRDnNTIwQGjSOs7TaSGA9XswpgFIZG8+94MQAxAdLXavTmm+1yO1a5zBY3n
eKPI1jHv3IrIzHlgNm027zkJ64nd+UCPfelVhE+NVWdeM0nM4S8/eQJ4WoRj
0LABlIDzWK2aFUG4PSTltfOb888DXFbXAJmmEQ0Bs/k+b88/+hNqW4HaOqt/
nE+XiSxHHqwqSWCTD/OzPofiF+9/GUtKwJJDBWxkLvlEZjeFD609G7FUb0we
ucQMcve1Z8MVlcKhkYTHCOYQggvk9iXMxjSJ1YNXQF8vf4IXTY73XLclhu9r
l81pvKbY0sFeCtRBExO5BbDAUqF+a0z0DOK8nwoPGwPKPoQbCUabBhs0JHZD
fMuGIXxjKYdobk+StR+Fy0kFTzcY+6q3Smf8IpSCr6dYrH4PB3wfkuBUNQ9w
A+de7+4LTuGQGbDk64ygCksv8veSiL5FgJgrn/92wrGWR3NI9wCz1PNLCW95
ev3elJRM0M+vOTHA2BpXLFC46H5M06z/xoGEmvvgmHFra/ePzdI1Bwp+6e/Y
cp4EygMA1yU4u2XydTHRLFYbUwZgcB1/j0W3Hw5ySIe27sOb9pYXEwk1H6AJ
tGxRdTTA9CHjQJ8IkDw5HLUqxaQL+5gD2YN4YsmhxbXcqNWH6STm/MniH0wm
pTDJ1Ot1UpMdNj+XV3I5QtEeHduvESIFUSwi82ISZYabbxEY9Y66U5bE929k
sQTfgOLZgjm6ALR5GIJPdHIQ5Rk+y3M2xd6SM6niqfP3ElFej0aD/IFzQJ7w
bA5Q2gkEPdPKrGg/fPpBUBrXH0LnQOfWRJsteutCYL7CMYyqCuz6nFPHUZjB
RMRTplbB9vXj1GlOz91YFCWQzpI4ANQxgNURlNA6VxMIX+NamLD2YlDAoXd5
3IOeDEIMCU2Bf+TL1xV9WrZ5PybEuGOTqBnriECm1Hc26kq5bioZ9qaGrtU1
9bDshm1zh2e+KaZfxNZBs10KrUICQ/43eKIbhDnBQBAOpo16vzstfM61uvNm
ey11TKl7ErctsIiDpQugzPIpl92qBDOZMbuJgRwtzzu8J5SKn+3VK8665Bbx
XsjjAW2EhCPFBGtDG7uNkYY5hj5w5TM9HZYi0ji4mZTAHmLLpBz/bdIl8Hal
hG6IAXLNcVbyFVTd4QM3Y+BRsXIJb+ea2G55fW2Y9h8Gc1v2El1L7kH4aMrK
QzzlS/MLsLR9lLSsQEgx0P/Gbx8DJ1BUq8DEKHLRZmn2j2BLG8afC+wML4Qh
7p8ZojnPS0X0Opb2Y9oip+SvGNPN92ov/QSpcZ6mAxDxscz8upcbPPPesziV
U6E2qsy8hbbhQUdHpKmwwtV2+GPwqDDXeaEDRhIXMdkNfb2kn/x3cpu3+UfM
gV9TD6OfViGCihe28Hq5dZKodUxzvx4PNtSL235sKHxsXg+/W7BG36CStZKW
ljOijxVT9D34VYMB7MpAwIDj6MJicglmp6t3jW9qvtynxBW+VHjXxpjGY/LT
uZtWgi4P4FF/Mt0hXHsBVWcQjCNBEesAYhLw4P/x+BlbgciH92YbdPJtVyon
HSY5S8X5m6WK/Rz2ZadLFpF7yKU5LK9+LVLs4aml4IROhXnmrbTe9Wr1P15f
KuICVKayNn+fd3IIp/rbO6EzjqXtU37UhMCWbWSZ4dq1xt5Y/PuXjMIi9QWs
IQgBR/sYEJedl+2MD2NAYIVxFd3KuGVQ4aK1/gaTngPGUowc/fliFZybkXPu
rXVWTqms+Awg4P9JWrddCnklkk6mbdSeit+UDPFGJRqziTQ9VMKnyZyY/n96
Ka++u6Ba1ZHocYxPtAuT1eMvNFpbbiz2QjVn96o4b0PZvEjKn5PlF5F1MzXE
v4aSRPCeW/I3FcT9wJ06snnE6Hv3sIEOKDKAzuKqQk/CluijS8JnyLqgWQHP
br5Nl5b99CyhF4mzyWZOybdmcnetC6Km+9epBlx16PZBHi6ayTvOEM3aV61q
zVROSi1TsSXTqjZIy3HD6fk0y4FmZdH/wmUdfRZnEoMl1zABfdgAVigu4dNG
zx4SsjkPv01gV5eV6ol5Up9+XZBKymKPJbavKNKjS4FApFVwSIycfDaeBFcb
e/GaYV3JNRKr0XMDYpY3V47TxkIXFYrfZHuzPHhb4LEfxr3nkziou/B4NwTI
RCbgVc2orevOAPjFr+w4KKKKXf4OQyXKQJMequfvbAVddudfVxjlED2rjeXw
wVM1nBe+TI2dI4Ptj69MYq+gFcIoGJMrdcR1dc53E/HEwGdMWMEA+pHV3pUW
DFJUybWkZUOcj8ro34azaFYfATN/ZQBfX+OZgqA9U0O2KxYilYRjsaSkyvRj
cfLSR78+ZYpLXD8RlAD/EGM9e/gDJh6jgV1GrvpboWG2mUjySc/D0hnk9A3V
e9PVF/APmquH/2X9B/Z9EBtgkz+fDX8ELS+iIL+F+SIQA0eHmhQVal6DwObN
4H8FTUItGUymREKjPVn19vKbtOaIb8/mGmcaWhCAlMb5sT8b/6DtGDzrCPNU
aYQ6oKIDJWmoDXZ/b/IfZQhysJwG3HITBLazcb2wuzNB8p0C/1k3mmK0TKeI
JslN/Hf9ZH959tLaEFHEH7KS2JwOwot3r6hspe6aO8PZgpJQmPoX74fiY9hN
KaallG6Rh7b7s71gIfI0j7QmF/SDQqph4icQkYnPIiiT0JOP4D2kn3adIb7A
eXwI91YINTwu8eKr8Hn10zHEdmvmVG83wbBvAXj4+L8TvZIg7lF0/HSJgYte
2mUobUjlG0ceGMRHO1rIn5dwpxSWUJvz+7VRIilzh1bS7s8gNYWu3hrCBixs
w2v/Yv/gSj4vzCqHI1CtNG4LEhN3bQ9XZ8dyv3qj3rzaEPqu7KqtMRuKjuG0
/+CIgcCt9C+Fvvx5A7j3J/S8RX/brZe/llXhJVQL5vXlkmapMt9Asve4svHk
MNzowLCFBpnAhQYTmShKx9j1PgSxDru0G1rVmpY/GRnwSyoPnurjUAFhQuRb
KWQ/3+8Vfh/kgWm86lo94BQx2g010y6o7HGWSXWNabekKB4m62fUDNxQlag7
vrrFSsnJly7tgVFJktRCg+kaw2D7qT3cIf3eLyii2sotdknybM5xYj/YGCF7
TdKYOz60IojjSAdPDMmYr+NzhYClYj6tJrY06+MxT40USJOz0XC5omaspQmU
nbctr4P3gi5POUIUMb0BtpYQlAZhVdG6rB6GGb40mHTu9BeBirDKm3NJwVKn
OnZNu7f4JR944xlQ8B9H2dBzjx7GLR3t5fCDPtFPRwdHDtRBKlOi6o5t5yPS
sh78utIHblxGEDp9jTy6TOymYFAt54FdZcRzTWDujvpiPSNfm6Onyeu0mo31
etxp9wYYjbmd50+h1axP0h7aVjSWA2+BmF7sNgsAPRurCvc9aMLe0Php2vBN
d6EEjd8AklKHsx58TMqhEv0ThJGjwONF2sp6RHcfGvWJh0UowjxJhLXhI9pr
aV3BzK2HWALCEqxqMNpmtNwS9PdkMfyzf4m0VJ0loLF96+oPjXhIjT7hk4yu
hvU4YEfHqRLJX5Wrxp8UCdNCQxoZQqID7wjVdIqYl7EnKASaDrl9uPLWfwBs
s33Um7oa3tqXHmJbm19tXGADqzrM0314npY7/rfYK/Khv950O8rfgWtbdYE+
pWgYxW/nc7SiFax8OL0PZ1mO2XZegZyrjZssSkE1kO5pftE86OLPrKTnlEYe
cil9LDk/SXYfBU3a9EWKrfi2uedZk5XUvaH6kZj/VqBBgRAvB9M1dsw+9Mc6
x/MZ0lHnHHqhdutgY5ggnZI9bohJuTO5UlqxdC9RedVvIj7mOux/TFUoxDCJ
y9I8Pxqt+eu0r1uUnjlufCyR434V7F/6DyPgEH9ZVu6XRYYn7803Kl3xbNQ9
YggcmIpRGWFtvC2Vk5O2XEZNTiyoTU8eeIJspqAh/YhAvTbBz2nVFlVgGfil
ax8uv8DQYivEYrefDMpZg4tyq/PWtFsOlOWisvR8Hr8lR0PIsJg6tLCdlnyp
uEaie3sxFssci2Wxje7jQayhUHmEqPzoK26XlMs+wimvG9cytkRgbTbs+rtw
bJ7STA+i46QHG5M8TiH7udtujbWjBWeFQhdQQJWt5NRn6FrUb4qx7URVj0uL
Xmf/CipHTV+rSZ0j0Fg7Y3YYpa5HAe/XzwZuCnafUj7wz1A2ej9KltwdMClI
e5SlPm4GQ2wdONG7YMNcCNag8yz/WMogTq6SNQyWGKAOOm0rFJUtTU4HJO0A
eTvBp7FzCFYqDe8Zoa85Da0yOJRIZ1+ioerZjBldL1DjYnOtDcoKChcuYwAs
0uv3o+vctmJwrfeR6u8U5UHrLU/jov0Pu3kLZkFjVy3pHt7MCgydTy62QZxT
2Hf+aVo349TsC+PT0RmPyOJSFvB7axciC2Hojz20mQOOSrAvu3z30AaDvjJm
ollMTu8LI02aDiglcvR1xLYPIPBoWS5iPHcLr8CQWOHaJks92HgDtxZYhjm7
JBucY9ev9s9x0/dfB9x03DSjDLHt3B1HyQXKIkyCJFRN5lXZPLsJ4Js4EhrW
NzZLUCi2VNj+2rHn2S0oG3Q90alejMm6LBAaoZUhCDNABPH4HMS9qtiWSeCX
yWugYUnOLnxiVvcG8Z0+SBOK34CHUZaAP+lSxkEwixPnOxB9mWU522BNOQUi
wXbRbdyI+a83/Zx2BmXgsni/7UC5hPOEWM7J79y3dC0PuNFb6LojN2PbrZKk
poFBlwGuvBDwTabB44j4P11Qu1fA9MskVGb0gesbRqLO/EZZC0Sy2YslFCLg
ilDGqnQOsq/ckCVoRGP3FoVSNTknEX2ghqopVzbYloq1yyDKEjhxrkUcmHGB
K//EzCRoJ2bomnT3PwMniuEqO+BIyR214cZ6rce9ZqtDjT7CX9Hg3QzI7lvB
h8pqHzNIXR5X8XR3a+nlMH4z1Q0xA7KZhgXSAvw0gNnAXtxHM7SdA2VrGoi3
TKWntR3lKYEVyopcg68uoOoFlQUniE3fEot83ulzV2MFXW4S1kUViUU9uhCg
wl1+jeIiYMzsrhkjU1UJuoYsRhZwi6XBFuV0VN4UqW2SGg61BkuaPWiXvJ62
a47yxysq+s2Kyqw2CoAHeXAUovszbP4+7wJiVJI4Z9/vUvS/oj1GFj4bQ6i/
qWRBaJTdk8Yxyh5ILdGNo6jqx2szZwjK4H9PGnEpnmpFZwricL3+Ge3kwNSc
aL62gReexv8hA+HvNcMJw0tkP4G2RSjh3303j8LqMq8tXAtPI2U95e7WgzSA
qG4N4Ew8kJmgG+8pA88b091d205N+X1+2N8zItpnXMIBzdyA0/xrSOcoEiIM
m9+IgyVmufH0KT532q2hJX9mBa40hs+wrwD4zb26o4Yqa86n+01pD6unO1gZ
ORdrkDE614SGozUJMTasCJ0w2EW0v9UzqlE50vyyERphC4C++3tXp2icKLP+
4ehVDi102mJDv9+MZc7cTxAMMox0hT6sEhrHm6ir2XfgnmjhmU/sZV3+NP6V
GAjTkxqw/eEmmCb3Q1+Ll8zYp+RyZjEaKs/MAGx6h3Z+BXH7vk4BawJHFFU/
K1l5KDUjWqWu8mkKFuiLHojvVJJrXqE+cC6b9C8bagcy0/CGCKymfJZOrXKN
fnTxPTnXEpr3yztRJGBEaj78VQgbVoKWbPRoMKiNe9UXMH/IM4qABsXUPJsI
js2Oq5wtz5i4R1CH7XIrZLkNM6T9jEocpLiX8XJttL2LHiaPcS2ngtlKUACC
JJoNDMtRgdk5BtsXYHrCxZrTbFPOJgHfJtlNcs9chHb1uCGg8qd7zdyAEqrA
8i/YM4WMPEY5HMUXI2FBSlLqLg0dbpQM0p8yA/FQ2L1SLVOVJQ6tSf7Z+bMl
NGO6O9kS7dufPNJorg8mhepZdpQ3RQgzvfuJp6SORK15RslDpTnzKWPUwdCJ
LlW63ZvgJHd8TSBEGZkQxVlEBg63u7oEgsoHmuB4AMtdOeEMwweDM9Cf3S1P
d9R7/p4Z4fNYNewKbqogIDpTtfTUdFxNVBwxcw4uwagAJLn8+ZffsJiuiQhP
q44LF0bYjrOWHblxR1BK7gt4mbAne4D9TTwkKTyYAHUvvnv7JCIMK2q0SUG9
9Z+vIo6ZdFpWhtmQnQW50yoHizgSgizxhe67eAM/VEbxFVWY+Sdlgs8xb9vI
uA3wCMoxtRhMC7fh+gbtFftjeCn9AfaUOoR/fAWI6FKO3CnG2IskE1kzuU5X
LMFHt0aQg4c9CsYaTQJgsatrQKKgSw30T/cEm3AmYWA/yXTlat/h8GfjIVHH
UZV/yDxplPK8WbPhV10Bp2EKAthzXwqNwY18A/jfJMQ84ssuDxpphUqdfLzO
X0+TTVW57Ro4BipTA0rqQHkc3vBbn8K7VjKw/H+PCI9VjmKb6GwgxA+CcXJi
6DUpKWE3fcCz40zCD9cR+j3kOPyAJg9v1E39M9n/+SFH3ZmRiyWC///lyU5q
Bs5VCmqdxFpgx6Yr7rhTOlyAs0tESpvxLjNiRT/imD2RARYpblv2r81mBuY+
7blwzl/npvrir96sIw7U7upyfG1J2TRggT32GoWX/9CcSlehoQ02k3G8LtAL
GthWr6arGI0+uP5Uf8clUe/zJueZIAq36+IH0NLZuLoMZ6iij5hCuZuiySbe
R7h3TCwTd3RNCUphkv18I+3CWv+MODKxR7My4WRjNO2kF6wbZEBfKZw4Hz5L
eaXIrYtCmgvY89ir13vpvUojmphW5M6l5Sm3ctSbOgmUhltDElt0Q4PkDSBF
3P1tlVfk+92EfnMstvcc4OiAgW40pKGy719nQfoaLE+rMf8kUEszalTH/6d9
pQpNP5O1lf+iFck5f9Nmkf89NWvMHi6+wucT5JdftBYC5VXMDARyaPCzYnqR
FVBu/dYuEmZ1fTDMNjjOA1la1lX9Lm74PWDEGQHeHoX5sts57jzmp396uJ2R
e8Dt8t+pDQ1ZFFZyfOB22BtkZjBs3kshawnShwEYdErlBy0zCJ7hO6hS2XX1
/I5xDKFSReeZlhxHRzH8pm+nMI00UAGMpubwFp7u9Y7boITFtHa47gD4gC0t
zonjyXdTbC4GZ0mx991X+q3B8UQ5c8H4E9S03F48r6O0EzUoj/RqM9mI9Nie
EyKjEEnrB9O4Cwo0CR8i1BMGqkF0NJa0T8x34mhKJsuKK/iQrUovCBNjltZU
Ynd7HFHtyzrgIK1QPoRw6/OfXLh6frdUEctwyksmRNHnMAs/oJQJWA2LDXCT
7aZmgZJI2swh0pMNgl44lbTeO3apWqTnD9683QhniBR8rX0VTaJh7EPMPmSj
oXJVSSlpuoPbFa/4t+ygAaAxkL6C2I13JATmSnL/KPLyJw/meqvlPyJJ2OXh
AJV9Yp4DLyI3ZPI8mCRNrWviOrVefG6PVe/8OnA2vtg3zq9Z3fBpT6Ra58QT
tJVLwymhQY/yyjm5h7ToG8eu/SPa1xQgCJxlqwF0Sjjpdj6KvE0TSbnI2oqT
8W8kV4/75PlQi51cRDjOpA3ym1CUMm+8Cpv5BeBA2V0Y8tZ2gmraG/VIsYXE
YRfYU80ctw7m93J78rEAU3TpWs+rGJeO81JLJYq3jQhxWs9p5XAjE56KeioI
RQhIIJUP+B61muU3NCXdI8DczeTCjs86xOY6Xa9suQNyGw6x4aip1lnNAGyz
7EY6nHaQ+aR1TqkdH+5AY+vCM6plw6dQrvHU6RGh2LQZkQsCcxaq8nah24OY
NjK7lRlPAT2wJfM3zMvCLtAUS35tSq2PQYqoXZ4BaJC0Z4He8RGArkSkWTW3
QbUO6InZfHvzygS+U7uHyehOPXjcAm4CPbHZZOM6zU4k1dP3renV5wCh8fmK
l1BLZ0oNLySW4bgVS0az6bVcnJaQ6eolcVgLjM8pHOI0F5c+qg/ZS+ky6i5n
TtnlmnUATHRPflNAQij96UEukjCgkObfH7ewmWCl5a59XCt+lEtyHGOj9pnO
/eSlIPE9Ov3huqkS9hOAFMWx6EBvMsXFGBGOmjw9TChzAx4Y+FCtBzPx24wj
nZCdL38bjD0My8v3TUfD1B80bG4vJsMWR1CvC3g8usM8Z6fbcNAG+5lHjAFG
CxTMlo+6iNk7Oml932JTMWVfuW8pdvmhM0vSrduh8x/dEjxWT3+zkaqWoFVx
IoEFfEBZEB+H648luwNbYyfiOG7eWPbCDZ0fjSrck3zZO86i25RaDKc9NlfG
0fVh4XEuY3ybiRzBZFMeBTK1zofMnPl8wPrCVpEPYuSirCd4xUnYhma+JJYY
uLP6JDjvdRNqEpbkjMy9UbEO77M3EIFnTJYhcuM4uaEzSAXJpCdI/TZ05nMG
UVraNdM+BPLHUxWXh8kdYZa3x3C8fdyyd0PcUQRxQof731uCDCEqQL/bC9V2
WcZxPqObOfLMC7mz5v1RdkJVMi+8v2IfgtFRz2IdZspOyL0vpDM5whPmfv59
FVJIMk4AOXtJc3NM0RG+jj5csVFmBULvFXu8J+S+yG5O8vBQpdOD+dZ9EOMo
r01JzA2XzywFVLXOogiMU1Mk0po40fcp9oWRN9pmxRynREjVxQPT+HmKJFi/
JPXM9kezUG0efesGQZmSErwmXmCLVep0zfwxlUg9A01GDkgSPEVZH/kUWAAD
PjcT81uVWd6vUP46LBX0qaxlLAVEJDcnW3jdETygmYSQVkBqztnV2VYT+0sX
E82zxNVwfmaqMJ/QMkIgHCUyJ76S73qgLN7tJqRyE1BeCiQyPIBvgqdelHdg
kzYJsGMJU5sdFOxagSiqEn+i9nE4jPJAJEXCAHWG3Yxyu/y3iYEhE0vLK1Ns
kS4kAzzgWDsieV0ABkI35o1nzIyPMgTXdYquVIj00+UbBdhmfgxR4XyFLPsG
IF0+s0AeC+YnKesTGDX/UHezX2RGPu9bRiiJMqqt3H3VMWnAaS0FgqgWm6W9
3QX4Bbsv8yQOGzFNRtK/JVyjecF1pfwdHG3Stm9cQntnQbz9LN/Xro44p0sc
KZWP4heR5T3NFzPVLUEph++oXE1BV5VOsqZeCp7nN0zbG66D8eehzwHRx6Ue
TfBRAxx5fNBaV10WgPPBp1illJYDXvWzOSW5vsaon9jyTO00fexN2HhKiTjc
z24+MSn6qq7Gm3j8GiA7MThOeyWyATYWbEgtj5ZC+K3z2uwJuVCtoPQ813mZ
z7bY3MpLbFG7GMJp2NIvII2wtEna92HsO97GOWdaj6qx1tRBXdK9fx1iU3IZ
tQRy0yG7B7xCHIx8ChsNp5kSGGla3JiaR++SruubwPsh4RWv1jR+EECYhBKM
aPlEZ7N4rNavNr/aK/Q83TGMxklio9+bMiTIz2NyWhY9Jn9C23+jWjlrcG9j
udK3aPu37VIUZ4/xNfn1DkBrurydWL58an4O1bKzbbHv4WWiKc1dSrADHj6x
fTvS7syItwSkES3N2bSJnjWBJ7is3uhxKpsGo7OwYxuDR/Q+skmL2FmTHzTa
zpSfICw3gteuuqAc+bCR7mWHXKrrUy1voObed3KAU0k8kOdmi07VAyKjiFlK
JBV4p+FaDLktrBxMyUZi9hr81f+Np9rlL3sU0geQvzVDvHPYK2VbI+2dtJHz
AFFDhxe3pUoESEQv/Lzmh30Z9w11glWlQymkNuNFtv8TKSllqLOS/1GPHwfa
iwwTLNb3ji4Il86n6YWplrtBW28buoSRb4quCIL1hrI+zVl1BXIKwah7oDkR
2L1ylAYQbSUlcHlVPYxTT3vaGMGrGI423ykvyKyyjMgkm8FjXfIE4SmnRzMQ
QjJ/HJETdBa8ednm4HAaDiU9i54zn57nvBx/PPmhhzUuZYTLLOdbaqWX07c1
BS4/8bdVT0w6xKW+dXgRMxkfuzw4sMwhmbioLPbo5BqfkBJQAT2IYRZygk2p
r28ExRnT9fcaAJl+hjbik917Q+M1g9UWpzf45eSVzM01hW58IS6c9wXxXSPa
8ai32L3WD8W3MCiaQyD9lH7mfUxAkDSiW+SEqdqajUkygNw36jWzsLix8G0J
srRoXwQJ30Da8ohM3vlWHqSNqzy7FMk3lAfTQv2J0G2XTOqsiBzMbYyzcDen
ECLguRnVl9pWwsUPQe0VDG7sVDeOsaajj08ZaT5mj9+eZ3z0u++GtsJEt7NL
czXalEmvmJYt1dSLlUZmVvNygtKaga83V+p9nahz2OHY54QEkHX/0sSTV+uB
I2stouVXsTrh+R1gM7phKZPoDLCRkW0pAUv1zQrVqolLZ1dm3L/ZZkYSMzg6
MSWSGR4fPOk+CgDILLxf0K7Hz52IEVJfCJhgWzZNMSyaAd320vm6/7ef6VvP
w9sZc0JDk9mR9hAYerfclM64hggdVo6hwcupsBXKH3EoiM9HpJAogIGJ9UJY
K/ywA099k2KfHBFPpSjX1ycY7cb2nqphyIbVxbKjUFu4NC+3GFXrNUTWvKuQ
z3RVT1WItwkGv93+Y4+78qd4lSa4CpJkmQ1FA0KclITl5Wde45XktkiPKlgi
Fw0yI6lYBDrJ0DhHBw5QCUKb4cD+PfKHa/QrC2dgn+N7T2FRU9JLncPI3Dbs
U/oHQf4//ZNNXW4pB70CFBJjLJM7FQygZIPJtb3DwFAjhPU2z/ur+ZzGI3I7
bt1Qu6yzQbJ7G4LMHtBStfV6fqEQynpDwRUy2HbX7iEquiVvkqxetzEBd/Pj
HRQJ+EKwE08dQsQ6pqt5OKr6zTuXsa21qZFUmNQBeijUNjxWwKq0UWOCOng8
zSKraaOtiupWfNfH04khvP0gAe2mzsxX6UGRnDCSAX/TtgZPoFIYXU3fCiPB
rYq5utcyayAsMriptTuL+oZBo0zZS0M5UibR31vw+9VkrkXLDnnN/xaB0S49
LLveUSQD/mcWlie3Wn5fTCBha2DyPP7U1zZmgvqmv61EWdF30c5OC8dX5fvt
Hp6sNYKm7HTFvWXf+IMWnBQmwRKQtrF2gR1Gp+/14Xt4zIpcebCkjBJEUHq8
FAxvHniESZ1IqZRDmYIYX4yxdHxu19oin/GYH3mob2cf+4Ie8HPydQUKp2XX
UuqwcyS+Q1Qdd6OXxSR+Ok5IExSBLCNMzQwb1sDy/4O4eUopXcuqP+n98gVb
31BxdKf9NFsn9VXBPm/MTUa4mFxfAGknOzu8c71OVeWKKDliGtvTOXchRPbd
ssmKEpyAaiEMowdB3RTZ/GbFgDprfdgWvc7ZQlQdTkRoU3iibSw3gmcuTIFK
roV1+U9MSR5jiz4uc73MV0ime+AzcSqfb1/YIgwZg/6pAgoA+Y+ChpiIev9K
X0ZOYvLOPC+Djx45dA+t0XjLD7J8tXzxBdCwLaj/VVPoQ9hL3eSrQ0+92SPJ
921ZrfRvH7Axv+I3foYrnG5s0ceBota6EF98VHij/tXOQfNUIUJOXiaiOD3X
bzW6wE/dFCYX4mwZQqtbqtsFlhL6MGJmaY9DCZBDrwXJXujlaYXDS2XhqHil
1t0vP2raoJKjy00s8ggf9G6+LPqvs0NLDCyvJ/Hj4t9BV1oOyDhdbvEhK5lC
6rvdS5ro3P1VVzJr8uMmsvNdw4W17H4Ge3/k0fJmlId6xyxW1+yILaGugNaB
x3EbkeetM8Sa6+T2ySmT4T3vOIGChUTj/1i981z8yQl9Sdgi8vV/vrI7LnVo
VMHZ5DW9iqAo7it+7BAG6awEJke9T4LZFyweUenx2rnHORpfSglCDbsEfzmk
vZhOhcRaMu3dg6UJIeFrO/MGhMnZjN2L9JhZKUAM9geLMlYsSI8/nFZDPCKJ
iZWuO5jniD4WOts0O5PIZEd0llZSmd8g1PZpDSqNzanQpvcuc0wZniqcny1q
vi+45CzYatSLYRlwXewpXaDgE+WnuWKtls2V6d3u2DSayYuNprp5LX+97L/p
vQQxRhG6KvAoEnRVcLyDmT0adguBXaO82Bea5DfSqQv59dwoxblOgu9hN1uw
/a/hPWLm7hJl4u2/kTXv6iaY1/GLALdQj37alUaVQZpW3dHaII1+ghkum+0l
d0Gob9hdqjdwhb86i9wA6OehQ0J9/ywD+KV9kWBfmyedHFz+8IyNotCmlhuS
7V0Mmt0WQsn4s8ljC5tgWFKkoVySUTyXwO9BlfKT2k3xFHp4Y6asMC96aO8S
oBPNfEwH9QfEc39u2M8RaYt2TKmi8+r+XH+V+XH5q09MQzSe3gFG0pvEzXKQ
LhwXkor6Z1b74Ty1axbNzvl13piXRJukPGkNmgb6jHXJGpjkQYdErvtsVEgv
coDxUVYy7JebPPjZGgso78PSTQYE3pWvFhV91wa/bzhfk/YI0/dYPOXMjtR+
8y95Fcccwx02uc1WaaFDadAQoHZPzh1mFruELsICvkwT0oXzai7ZNuvH2KF9
WiApzG4tFmjFCmEumxmrCCZIc98ebbH8EP8Oi/PKvRJMtEYNgIjw5jsh5JgN
4kFPZDRxnPGufYkrFLn8MNwxJTuR/BeZlIPe5GewFIQ2PBIJnuUWUnaYwPEo
OdPaz/TotiIyDsTdSPO6UT2rjYqAYHMVCcOzuIf2CLKeH6OQ0C2gXXV3mbjH
M93v3iGyBccylbsDe3CKIKtXXhU5HGkgf4o0P4L10h9IClkthnFdV5R2Tc8x
2wY40XyrwBqUL5XGoP8eaSKG+GGVhHG9IKdHdzLBGA4J6m+qOSjq192cx6a2
jYGjYLVt7JHzeJM22hCLijYRvVbEkWbnsjRQ1hs7OdywR8QaPSkyi0dUYuVs
WSd5M25WKM5uaPMQNZRZL1JrX2ouC/n0nQYPJijDMc9D1uB62QJZpwYYJwOF
Jw6ECHKThncMpApXgLFKLTJdso5mgqdqMctODjVmBk2rKqoadyJXHtCQTy/T
r9IO1V2foO00Fcegs+oi9A7zkp3OYihWN9BP1Wi1nVENRe+bdT2GY/sZabvZ
O30eOVjXmErXIikkjMozYgg/zUNcRll5cPBNNwyz6xx0DfhlssVoVuV0SrE4
7Sl02o9rE8pQWh+uZ7G8CUKyJIKYCmv7ME7ORorPXyN8kMF4aQOViVYXWx5p
XLId7DcvxlX3LkbTgEXEVO0gcQxzzgvY9sADDTVTTZSxMMHlS9qQY1aKJ0Vj
OnbrEbCsZiku/u7Dk6AVYwVsKZguLHK9Z8Y8+R1PYd95/mpHMwFEh3x105C7
A4SA8g3fpvlO1n36ueVMhuQPlqgVeeOtav3ZoezOYo+o9bAuoEBzI89FSsaa
dq4fyBZhP3UzhpryWvVtHzxBfN4hZGmDH13afa3z0VdjGUtEnsBOmUeLBRCL
GZVKsqAyUdHDR5JhDzJFvogptJyFTsMgfqRwhbSFrSNohBXVLCHPLIvLf4IX
n3+EZL4jgAQaX5s6OsTZkuf+/MqeDKnn8L5FEwPNDoCAalXSOhxrZu12UYKb
xInfbdLw2wtW9KjYSJ+ymK3TGjnl7UmAFodBdFyDpKEB6w2xnLKfq7w6O9n3
tKpbVG6U0iC76cvI7Qvmvh2goVp0wlLLc2cE8CGsM2qMoWKHp16T7LCTSSNF
1IFT/Hx9HZkCMSPD6HB5dUSq+4JKnvtvArGHKVtwXsq5Bsv+wFQYH5oXSsqr
bUEypjFGl5IbpIAOVtS8SKgnIVP4URAD+v5CgXiVj68kIbEDrj0piTOG8Nyv
B9ir6lVZ8nBdjhDjox87FegQSh3HNCURSJL4xOuoThY7CGLyngxMqFcb1zuq
Z83iwaYgZK66sjzarqQ5/fB/5p+kUvhe9yBDbOw8kQ9xlxMQqzUh0sE+VsG+
t6qCD1uOXqpZgLziqGLhUvvoJiRV+ruOmCevBYbBbxF2+B9ZiTY7IASkE9Nu
dezLYF8jp5kWsXK3WWakFS3MpG+wHE86IAPx+kbWJpndjAZoIN23pzFP8ADO
fdlx3KyBxH5a8WS5JvOPQEwJzj5ugiM3NQ/I9WIr5TM/JTFP8ftCwPnq86B4
SHYM2za23FCphZ8CIBaBRjrAObrix1/Xf8qe2LNRXRrGUBgsaxH1AmiFTydV
Mek3d5YG34XBmhhZIJFH5U7t82OyUbPKsW8A8ThWJdrO72+amFDRpRlElSrt
yXOzZ0hgR2n9Rvsy1/pZUhtEQYaVQ+HVAmRTs67tc2m1BeUEjcgNCj9jjR6A
Lpm1mUxJvizFaNq2kSBTrEYhawaWSCNn0FguZ3odQcRbTyv4/043y7uTM8pM
Jx5PdY6uzl3+LWl4wwgqoN4RCUjX2/NwSgx8r5HI5HYZJNuNCjttGlVGvFEm
Wozac8PkvHBOvSX39Rp53ALRhrePUTqnB2BKygh4pt5Odf1K60WbHNIFenX1
ceQJO0AnzGG7X4MetPDW/ahqkgHBNk+2hhbYrqM5bPKmNy3AlN2dfmqPPt8p
FHUwWLBQK/8HavGb2e1r1XNvb9cA3j/P3rfeFyldm2GZrixfOM0X812a61xc
4Pkx9RMorBzvhJ5XvQtPizq2rNwyLzcjZnVMBtsv3f27t4iPX/SZ04DDuFu4
/nVed5ff5XRKvzWjBfYSMcFbQkhzYEk0JPtmAPHhQ4vu7q+XHyUuf7v9xnnC
JWech4TiIvP5LuwKx+r5ppPtiJXg4zJ72WQ0UAG6vndmSu4G5XBsAaYAAtWc
w04wIShqzh0Y2vDSkIZ+ARVGoVgrQPb0JBSHdZBlzLCsnX697LmedZhaZeW7
RTGyd+RSUpkkqs5++KNcoHLsMBPJRHmEFR9pyKqvskgGX7BwC76fgip0z9mn
3z53zlorIIw80k1J+x5HZ1HW3sj3+ve95IS6EoIO5qAKBmsTKW1xEQOlQJfD
vbxT/eP/uYkuFQMKgicCEN3tKZCDHEcftZVaUcLOjTEcYYaXJ5zGvf20KKSt
WVIkvhHa4B703dbTWt/fdZMPAnQ2SOfP3Jm+xnHKPNJkxO9sUbyDt2cDMvsL
6h5EESm6/oxJy9nv08FHramEIDawt01Jr8+30EgxEf/Z7OH9AEfoZYkRQyZa
bCCb5aI3ru0+s9QRrZPOvXPahaP3jzHQ2i5eWMAHhYLi35EnR6RP1XM6Na+d
y7Trr32fouQIiyp1+nygGsXb+2ZbmaZ3MU+Rf5WKZQDHtOh7LZ8Di7eEWmMZ
eP/wZv6P5oGjBeEW5kEF/d+uw4EcC6SF3W4tfwqj8vf7rgDYOl2UvJNp6iXf
SdiuyzWht7MA6w36RCUsMx2bilMEcFg51R9XPirkbbh+kl+MoaoXUYMWMOLI
Nos/uyUytW70GFErCChWyljfkE9azgu462RtCQgoVsyG0r6Ym2z0GjXRMDEn
WSSfKUNbfmPfUcTOEwDid7ubVqKMJ3KVRgBGZbbHlR56vO7yw5+0O2KZveXX
8c5eTAG+dX1/WAQ0WHh9tK0v3kiMuVFHPX0sC6dNLWdP9b4tdxdFDKEGiJ5r
r9a3QvbNa4qtqrkDLtDKmoPzOZIBxXtFWrCkmWCoe7PXekqJqVsosSKnmFrb
+c1MEfXagS9lAvXG3sNI9McmaNTV1P4hsoyvFDglDb0FFBmXCHfURrg/7GTf
pZOrlgl0oloXdQbqc2BmvgF/Si4Xfta1S4aQFmLu6QipntJDTiIi1Q4RZv8Z
jMc/gCeYUarpVnbze6NfxXMBggUJFld4DWrHZIGx3iKOeYk1bjnhJao6E7ol
DsqFGy+yhoz+nYvhD11NvcuNrLs0/B2th/EBfX4F0E+5bS4mRfGcIGdiRoV+
zQYhxtTsCrFMjBIxV7osyg5iT3VH/4WbArEoZyHviip1Ys/s6omf3Z36n8MH
GMg/OoKsHhTouDqCCTZtm+9aak1v3L6FiTCNCvNlQRwHzFFOonl/87v3bX77
YMhaJOtU0MPzrjiByGZrmb4dXWaN3LL0xjUdIx5j8nMLyrLYf2COIRnZhvxP
QnL/7AYerOv0q0OICcM2GFlVCjEmCJYxr/IfxhlnX/Ci59kygfEMs3RiqyqC
/bT+edrt4eHdO7plcjpyo2RwPVlDEtf+H7CymYgxe8YFlDP1X5xIcDA0CKwm
28UDRdOpA1QKMFCIZaFoELN+u3FjNuNAy4QzcDIOyfai+8di63l7rEfVLnT+
bfetXXyUUJ4MQHI+R38t8eCKvFpSmYNK4OdKiz0YHF2/9/QRcGzzZ5fAI+SN
/hCo9dKoIFcOwR3cXGvBsYrQgXdEvIidXGFMz9p5v5QiJTJ8AsO1EJgIdH7X
KzP/RMGKt89hzN9rN74CFl/HEsM85r5gSKaWN2MqwMguvGcyVlrYt0vsZgmq
EtxrbW6WRqfusQzJ4tsB3ZEn/u2XYgiatymXO+Etfpuyd843eoNSEfkVaHyy
lYAACXpwCQ/XXwK8y5j4pjNSu0y1i38aSnbxiBWrwss2GjrWv+6qXEE/QPox
m5wKRzlTmskNZONkwU9REt2Ov2BxjNr2/pYABTi/iFLNPkBaGgMCLPaQ167e
P+UI0bG7RrPL1Lj4ZTRUIg5axp5HLiOZsq7hBDUEhaIK9UGRpIqa27Rfuk6E
K1fOFENqjnQHlukig8i9Nrw1FXf3cLPTA+tt6JS7I4ft4gYumobefvaYz/AZ
c2m1NnL21eHNQF8k10cIVbg7iL16IwZZ+1MPTD2MRTaRKglDZMjkuA77bAF0
47/TyYVdRGp3qn3V1TJ5NJtvfs6YaD0tvx6r4ey67cZyrUCBcSLm0sbOGT3g
R8ZIhQd+4tCZro8wiQrEZfUVP3y9WjtPlrn2PpdgajQRMUDnvqby2jO3OWLz
NODleOmqloVsKQPkQHa71wHupQDZmy3sE0171mI7YHrLc1hy/W6078lzhJMQ
kUHwUtf3/KGSAs2aRZLwilkMvjrO3H7Gayi0V81bUQF8ej9D0jvgH/24lgeU
9dru7Jai9qhIPaAfRb09kYOgGVCrGULF7Lv4qF9alufoFkvcY1J5YwmIpn7B
upXRSyFjb0r2w38ueNlwOP34cjegFDN9qgpvR8Ae+tQOC58Gf2wiLYGJ98TJ
3BQen7Pd+gCeBG8SDyDzM9lgfbnam8uKWu7bm2buNpo578x5ELitOJq0O4u0
4ekC6wgLk3HkSXzy2Jiu8TQFrXc6LxkQ09SKTr3tEPrvlBjeEkfAEQS91qvv
S69h20QhJaqw4l8JyBxpj4L5TtOsq3fdzwHXuMcV66Rqx/EZiZkR/Xk0o5PZ
/sv2n0Lq/EwnzERo4jzzXGMitWWXnv9QOrgNTkXHI318IuOV17ALSkqVQ3vH
2xusYixjvpUCBY4THTKNGri6reWg6+gGUupZF0J9YnL1W+vEPW0JEUBoIQx5
bQtluxUpm/gRSpU6LsRBOcqa8txJLaGr9rC1BT0y/06nYL6BNdincTy20OCu
tdosbdpRyssVCohFDUX0UViN48R03S0aez3I+aCsdAh7xhiBetpcGktrcLA4
dDKccxOG9H+yUUGBzMeiTlBWjRnpEZQf6C1d6awtDNpSD5vxevwQcBm4XQvJ
Z+TXX6B7zRQrYcWYSP3mGA4BHR9UwwII5mX3cRb+cylooSjqHPh1Ef1MmZcw
N2ss+wrmyEQYr/fcr5VgSV7ec6UO9TlE9bMveBCib4Cnmvgs2JbIA90G+MIi
DOvF0gfHZUdzfc5EGTr5oeALZ8gf6AbckNqxeDvsUQkQc0JG+h5T6uDR11TF
n5aOdV9T6TJ6K+pUMU372HEqOCsr4nL8f+jHVAOsfGs52REuyDHIwKXhiFjs
81PC8PYC8BKGRXIMW6fYthOfiDnfuqiDTtyYWNy/0n0YY10Cira3AKTch5mV
3cmd1tt9ZzVH7z8l+hM64v40BkZGJ8h4YXQqFbIRxA4Vg0wRHE+Apvecbz76
SGtd8I2Cnky3tjIPcu0QtLG/oADGlFiFf9fGyCFmDnAIBcZ1AnHTV1acv61x
Cka2BxDmMBwy3klJ+SrsRHu2V0TNAGd2y8E/4noxYfgVzLObBXyRJsZoLasn
SQODxwMVlCEY1RlPr0Dz3n5r6Fwah0TCdv+hh0jpNDmwf25fGv6dz6/OwveG
RWQn8X6ycgszWR7eIgcabdun6LsvbmCC16s9am2CeTLVu3juMcPmZABWTU/t
CKIZtslDMtc1K849hL36SrGg7eSup3jDL3cycfZnQRtnUCO/lQYX6fbE1ap4
xq4fZC9thU0L6Zb2g40JXWgm6nZIYsHT04ewHA05RupB5bvKwqFZqP1XXbgh
QEULBApC2gnGxtYhkoFnwtk6JqvOJfJ/2wGccnkOkuUKpcHiiFLGoyDEwUlD
3u9mqhEnUcI72MHLVk6djQlix7uGh7JjD4oU0pWL1iVkVNDCSeA1+I2tQQch
4T71QNYkHkLayqJgOD9e+xre+okYFU+PWUQoLk3B2t/2RWxU6lzvS6iGeeNY
No3Az/udoSXi/N5wN1Oetthwh0FPpGPKDUErr6j3b6KytpwCPRQcCpXAvqLs
czQEQzGItGkfeHd4xrvjoKQe6c/S3eQkH3p1UnXMYbExbq+Tviz6qMUK7ux+
8gAD6dBKKCpgWnZGyrdkoWl0ZqHmiMw+TD5/58NRzw83Lm75BbxDz2mw5Syt
/ZSlvTC+klASZ8NAJTwsR2jeF6wz4EMHxmkI3OBlmfInvgXloW0otPyPKDfR
TKgCVy/EF/UchljI1H3roZIdUEW2uB4erGPc+CJcv7U05wTdCrgv0A6CqT00
tSQ7jq4giDyvMT1o9lhKYurs8v/OcD72r3JGBD47jOJRIpp3+Zl0MomX1ugt
RHAfU15UDZ+KM02j3M83q+S+LUD9cgKrNAu95pIaFvS/ILHpC4326zGMjGKN
0UUqmZ79arusvuAQC8frUaQ5+bL+nttxhP558toiZHs8fq9K5N5Bp1h+t8sM
bhJUt5Rtiwtffflswfuz0vjVibPwyU9DQp0R8l337XWP7FSySyGfJIvxdBjd
GydZyDs25futFBbLDto3SjYzziyhFMGCjfsiIXxzdgxIWNFfBb6WM2Z7hFVn
nsGarvcw2HktQsF9AiqpBggeKDX5D1MQoaFefLsmArp/qdTbefT3rzQ6awwP
8iOqWO+ZoZErJF3GptPYHLdF9GTAdWu1W5fzaykyMroAoLvGUMVhnVpV2jBG
8k7AUetWEeCOarT/+S868CtJ6r2oMo61L41D1c09W/WF0fcqwhTMKh2P9+0T
MiWObIgSfpBLCH3iaHkNKag3Pl3o8hYu7mm/XJf4AOtj5Q0sda0+qv0pTAxe
TB8QlAe2QPQi3xorqUqCNAsDBe2N59IiVfElio4be0TFX5pYfQlTc4TmUvqP
PEW2w2NvzoJR+w5UiBZK5OgzhX3ynGpXAwd9ZP1/afh4lSl8IS1cxEJMtiks
NtPgBnn9gYVpYQd2J4MyqOpccHu8Ij9oLtoAr5CrmJm7hqoVM+dZCowHFOao
kJCWI+knieOz2iP25YIO4HmBZT9JwPvdcGp5nAWes3JCFVoKvo9Y7RLOLVMS
7hp7p5brSjuhCnONfdizm73Fe5PCbKKUTO5DMi3QVIyIhx3wzo2WjdRbSSwc
Q5QIUdgQMqwvJILUTXZhbjgf3sMoVEMle2KyrgioyH52xN7FFwmArom1l6ZW
HjHy7dVLvFZ5a1N3kHOFcvlXGLbv7teC3u509EcRzKjnbw6b0USY3p2lyA+L
MIlKxNXQY7iZjB9j3rA61pjlUYFEV/7EzN2snrriHSESbaY7OW7N/6XNApGL
qOk0BvSgyW5BPdKCrOIUF8t6FPoNio3vGX4c5U2oIR+00Tg8KgwDSPqLjiUy
EO3MNTrfBtWvXk7Kz4OteXyAKvG3EWQvkMtWV64eOFUDyDDqtUQl6Y9an84D
RTg39w7aYSKnYvBm0XwjuA4W6+WHmSHCcpA9rCc13eGhB+RlrDS0yd2x2f10
aNX7/2cTZG3nvSmb3pdiySb0TR4mRXMfowXsJHuSiDfpacY4cs9WJ4jQteXn
DKTfh7q6iEtpKPKwqrKwWIuV9HjeRZgmgzn/pEjVTg2aBpZDQd253ml/cqvV
SqtxdsrDzXRNkHtREsmvBl0EvRTMEpADw7X3zSsxZqnqXuar5Rxob+CL8USj
TLYIR20oY2pn0InimTKrPY5tsxPFEKT9Il3yeytex9SDgT6ZnJzjFooLdmX0
4Da+zYIAVEwhWJ0Ws5PGEcJqq6FpnrFsgYGgR6GVlp/auXBg4n6U/IUXDn6R
HOAHUTCRnnAnrRLujng/h02CYJw3QMMOjj+hwoURKre13ZBnpKo7nj/HH3lg
tthTSSyH60E0ICjLvtS+pUDR2concHtQHVdV+PqCtDOh8SMzWhVRJLN0F6Rb
Istkd1CLA0MDkCGkjwF0mslHEbeJTGRB+Q9Qfp/oyhC33028tOZuitASEU/C
q3NVdShNbAK3uylEM4zO3t1EGlSDaAdwIihJIbZIcDrFmH857yL1+705hYWb
X8DwTB0CjfJdSWfHL2rXQ/+YkEXpu57avd2YlVVGXBP/ipU7fC6ZQNBBL20s
BYLenna/wnkdHlxLJxenvlbawPEIo2ztkKGwMoCpgK4nopD2qa0a3dhANJWh
5TZexiX93u+pTPchIrJp2+HUe9qwGxUlhy7RwswCFynv0lOoCsMGSEStB4eo
d+9gxmD256k7oCbQJfzVUBF/yIqx1kwxQ8O26uQo4lhxm0A84N47XkUz0Alh
xjosDzq0bjNUzg/zHGNv689nkJ8nXOXUE+Zh7ctht1ce4iCzoecA6F8W+ek9
O4c3CldGH9jkBR2NxzqHqmPUEMFpo30oeQmpgQRViMU/suwmKo0SBjpPB8cD
7KMG7X55flej/F8j4q3JDdZki+R97QmFgUyqb+TrmYEYPMUgSkXKFRUICgKG
NUJKiQE/rDrSVt3JM4NY+JAMFQLXrgt6bQ9q/vy6NGHDIBE+9DHidBizMU+h
kBF0pIacgxKfyS2ywrdOsAam2LyIXKudNOkCK2f1CE3ic/mnplU1q7pW/QWQ
8nznLPhLfaj3I91rRkmK1yrzy2l1p3J4hwYWWX0I7hnBHnFq6zAAjANyxlqc
w/w/HegvtHNDE2I3qO7cL9BPioWKCRzxgEXnFwau2KK+u57BiLpyXQbF3mKl
Ga6BB3R39Ys4PXTpcwoSTVKyHHLupbQyKLHK++LLosi1F49/RKieeq5tq6F+
W1DghWqTcw6ji0z1tzNc+BvOdcJL9w0YERDO1mlqqe6ECcR50VMd9ezDOoB3
bUUv8K1pB9tUP0jjec0czEZfhoX0uj6mbWzCm+Mc6dYkh5FTKn4utv3SsX65
oxrHfzqteDHCqaWdTlZA63neIumRLlmCPHO4D+D+pFVrklLymu4qNhjMIAeh
0NplxZMSG3nbiojaVzV+n4x6AXo5mKBpsicsHfSk4JMgjO4xOT7baJnO1gW9
CPSTYc23lqkDSk0Oz/8YflG8wOcbHzIMNZ6Ix2hvgWNcYwOUpTQbT26Gu6dE
D/470B0FraYpsN8GajdUPL3vohQKgW1BHXoOHU9oVdg4E9xxgSf31TLjLDE5
mPKLSYZhspl207x+yd8xtwsXc4aMPHagv5HQbw1lZXw1OlgDN6PZdOU69q6t
25mzRyzpChupP7f3gmq7OZOhnhIcmgaTHJ1RuYFiRNjlRR/ZbiP70eC6ruW1
ETvhCF0ez/pNHtskK2e7iEg1yHDe/B3MjzRJKcjoIL/Oacb2akNwMoDBVg9E
6f0VhNov6ILPEXjwnZTORIQdvJR0EgZwiq1zApC5z+PLtkM8YWz2+bHkTjlu
RSTYYhfdprUuJRXtbDr0nHyjIrXTuLiF9ib6Pd70UkwYxXnlnaLgBktcLgfV
24xtpdVp0t0WI64WtUokwJTSVvJ4KYEx9PVjyzrWmSdPsfbeEq73DlhabzgG
+3WU4644V0glrPzz7gDYnUN5ggVMwrsqv2Nux3vWVxUeUYmrEpyJGGCm+D1u
bt/RtZBpDnNym3mbMPfRTGe70EWFiPc9vluiH2X4lNMnet55y5Mk290iaoVP
Kh07PVmeLNQoE7YhnbC+2lWHBlDpIitt37Hb0CZf+OJW/l45ucmR44M9PhZ6
0xZBaRaGx8UoiVwhgMz/uwQdrLCtZMoWgHvVUBMcqne1O/gmh2YI5KSa42z8
laPNUpqtDv5GMBB26Amwa5b8vBzImueZqL9n0mbXt7LsY8ZjxRVVPQnI3rqm
IN2MqjLekcbXUbzfEAiRRlUdjUd9kj2T3kxDzwDXEslr5wWnXauwjPjVmtkf
r/xxGQid5QNcz/fZRQqEshvPy3IZen6v2+2rdSPxk1Tv+LRMLqT13Gw18q8S
tEP9gwz4lBQket2Zhxa6uJtlDIQhi/4EqslBJVYSS13e3nID9gFyIhH+J9Uw
Y82E5hJjtWd0UAwfS1rNBinpDi3Tr1wNY2hAftOXjwQgP5vKXSKksBXx+nLY
FjeVZeSGeamuGiebLwUwXwKmGiffjQ6GYRJ4CVQWv7o8OMijcx7TyYbdASWa
br15VRtZxD7kqibP+t9O2yd43yfx2l5IoIJq8QDp0RyFjoz+kWin4ySJfZxN
eu/FnXyamPqiy5jxgdxUGbHo5eTxJA3kH6XLF/C8uYNhcMVN9d648+tsxiuD
7rDDyIt3nHHUBtFjOGxtfw8l53on2zYRLB7/7Fk+Ck4PGdZxEoN9jVVUcEQi
Sk5T4uifK5fMvKqTqNJPIwnl/gSlRUMW11fDOmet2mxuVVuTa+K7mZ0qY1cf
wKAFKel/G7SjEEENJBcDQhB3W4fHJ1RY7AAdz/41PVbfoiRmAsy/Xn1Wp/39
KXJeNia8JljWQhKd92vFI9XBiohpAT+XOLA1nc5FmHUWprdHOSVvMZ548xbZ
Wr8zKqlISeTo1wgMWlhEj+UbWWBBEaSOui7AJ07BaQvmfntjf24D1sx2NMA/
eikXp6JRfF3WTEHJdn9ZYTuDMj7xHkofpZ7QJzZD9d6vNaoLMwD0CL7qztvu
cX9A/XFnx7c6JAWJc9mqcscBlrOTw7bn35zFZKee729Wa5lCVYZJTo/3LNow
N8J+NgwM9uvNVpfz2FhUZOJE6qVyD23fPoQ9KWMc/pirWCmdmjdHDC90jSGD
zggIUU45flKd105k6C3Ub8IXLuihxhmJKi/wYqL8UIuRhaR0e3mjFl43Y4U6
pAreCZDZuHSU5V9ah9KWp9lm2pknX8sCg0FR92RpA1cC4m56hbxNXPw3QHiu
mB7Rcxxg52VDCvBzDSfoy0CirGm2OrTtmrROU6vtwgrxLEpVZm6uaqoLfUcZ
tKdyP/BOIJlpd6L6FZnhiZEyymTIGWAZAcKpIgwa6s36SOIWrZ+r0pXnlZgy
4WAdJqeN9sZd2Sh3/FMuTKjTs20GKhZEBJhFYPNaMT1eh8bURaCwlddu9lNJ
eaPGOFEyDmHUCN8mSMVHlH32GVa6scQ6FHN0zj9ukjr3REVqtrfJVkRtTapt
AwBBfiHCQk/VztYi2RuuxoNvfVuS9t5Y3NoZhArZqpbfUSN1i7l2V6H5YboH
mmUV/w3kuiZkIHGZg5hvVhf1SCQQbtAFG1ahUqza+UkyITWvweUqdG3Ji0RI
WHtKiKrBwkrnQSXqabr/0zC74ZF1uLVDZM40CmkwTMamay1x+PQ1UNuXtgmJ
Q9lck7j3O8eLtLviFFhtntWdHPOWeepiAw0J1CIMuvwC3AdHwOtND5VYldXp
YelJc85Mi05u5cWyqFp/z5JrF0aof4anWrVJ/khWPyE9iVJROAueL00XONqp
/fRqxXXAnFHrvvDFNnANNDR/4qnctOwXWyr6CgeUcVEDJfcftwlWPpAVlvdG
aJJxfKUyRksePSK/cn85Aa+ed5bUl1SPOsdgxKYAPttDzhK9UUIcaYM3gGzN
qX0Swc1dMYThe78gLf5ss+KTeCtDpSecB1e/oW9LLY54EX16p37SthQ9t4dJ
i9xqsQngw8vijo77kJFpJPwWd6IKE1UwXjcC2gOWEvSs+k+VRD+tAd2qrHBU
Uax9YU0Fgo5Uf+5Qeju8DyeMP9W/2V73bvTTpPQmYHOiwg0C3qQSDo2VHIoS
gbelH7t1A7Xmfb8/o+1+C/rrzVV7p0SUmPfFt0aFHMVKYVUOiJkKJnxXrCxE
Bc+KtZXKXPSQG3/uhYrspMdpUNFndeq0lHYTDwP1hbZjX93u77RDD2jo1xid
s7RNZXlACokqgPTJg6oahyCGGAb9HisPiEp+rD31LxcOMqbFu4q3y/12Imll
v0E9SVHUOQ0eWlLdeOyk8P3V0h7GK51hMRjQvNfMq/6hO3qfJ+ALopsaqn42
igi0e3J3V30IbpxiTtCU8mav/w15A5drhYFgZl+YkyCO1fAY8zVGgFLf1yVU
OR+XxjIG4TUoHPWc6B7ZOXRIXvWCJ0RH+8jgygVsNeBxWt7HcPIYyJI9VycN
iOPi3YbMcg0vFjsTTWakuaCYAi7TGZk9q6OM23/sHDpDCSgWpgyOaPNXHVvh
qXK6AIzCChmhRlG7PdIjR8LiW/OWYvI3OJvF1jjueoKnOaQSlVvRAkIbNEBK
fIZv7/BMy88Oek4pZ5yggX7DilsZLUubHCb4XUBHwgTBEXhUqORXH2BpT031
rVDHqnEc6y8Y5TsU7McssXLbpcX52VAaejA9zhf9l80PB7andyFHeJ7b05ir
x3QKEyBLWJBRMmBs47BMP01+KJTNwiGDZz+d5TFZOMEP9WyaPvAMngMHzlfw
elFyaAzUGUhOG1cvyoKkzinNPgcAPmcFjyhPID+ul7h9bHY1G0DBw5zfHaRj
VcBt2N2pjtXAJRonwGQRMklIoxKYGwSxTUI79cDmzyGaatdkzwL9267UgiKt
TF1/Z9+NwfZ4U9ndOO6TqTPG2OQPKuqQ6V+8/4uCX1Dziyhm0XfTeUQMQ35f
PnEdLuCkWKfFLokwxuez8IkZdcuMnwKDYlEciYingc3Nihkm1PnpqdhXGdxX
CLVJoIv2gP9csPlwN/B4u/a8QvVTzJ8H2CghhwNAt88yVo4UQY3Bz+S+ETyz
pb5Ys5jGu3G1b4n+4wR79MQDCjzc09NeQ/imib71Lb7z+r1mJ8c5m54YZlrQ
OBuX/y0K9fD4JP0vjcq0TEXYHEmekXreUZ+G8upBjnSqza4Qu3RHFPvtB4DF
UF/PNkIt7XSVGB6a4TtsnqcyLHbVO+0JgQvhG3LHF+B7nH8Ptuc1lzQ589Th
eLaWgEl+oXtQG3K316WaTlOEUmb96/w5evfyp3s0eI1et+A0iJmLxd7Gz7lH
ZxkmHOl5rkGc4PlhOihK3GK9ZKy0D8UfvpnskOBnbIsxHHPz2hIOZdi4vx5/
eqjpc9TccZjARDmCiEHDbL73sFNkyYwgBV8GNDAHofnfmEL0ZrDqdzKyZhLe
5AI6LIg6z5hrWIc6JVcaYlsqYNvBLT4vydVgQWq3VqN5iqNTqkS5ZzdKYbXu
B5U8C4mlSiPA6EvQCy5yNdYeGVrML8YnKPVLVH4Ni3hEY7kp/0eDQTz9W/Qf
zPEkkV8+V1nTpFXHUt5zXN6wIiMdNtyNQ53XjEx9RFAcVmXsQMbPg+LOuAdf
qhdmDwGLsZPkGPAIOswFn5nJU+gkTgh7Z7gi7xyrmqf5KGpjK7fnnMbzIfMH
xRH49ltdM4KmiNAIYzBZXBcnAQOuvr5Bt4XwxsECmBKGd4KNE58JT8sOvmyl
rtXV6Y8EAy9bAMFdZSfT68z7fwiEhVac0YWMpyH7F8bwuYZcoHrWVHjED/fE
IQ7lX+zN3NGM9D4Qkqife7J0x+E30KfH4iLM2hv0vtOPxyioMYpLtOQlWIg5
ijCFDa87Oh5o6dbISC8MhyK30uq1OgaeuQuQEFJDldi5DRejm7VI2P6qPxBx
fnh2VUuLqmo/gmD+aP4UscGRC/j+J+aTE82+shRx8CsQ4gDkiNJBOj3rcriS
UcbIp7CYAWMf+D0htT6u1CBG0wZcRTjhzH6dZx0ILZ9jvoHlWVj66SWo/I5/
afmKV7NxUmiMIWCL9zoqzNfd1UmE00iDv1dYabMDYq6IWFxVDnud/zX0GaGi
8x+hukqQn0HnPUfB2g+lV512EdDfG7z8bAx1OF7iBlhAdfUjwh+NGobHrK9Y
rqKpNmjJh6scTqw5G1oXu7C3wlKgxy1Dv0fawNkkXYfs0pze518ltApPulLy
a8Vx8ZACNEIgEru7HP4WRWXt1rPHmfCl0aEFR59gYSFacKIVXBEmEoebhEqe
YiRbKfgk4TdO1ZwbvzwKDXN6q67sb4I1dnUorVcykuVHZENgeDGTZc2B8NgB
3pxIIEyBIao4Y1+TWxdIGXxwR/Q4B0kTxTgZG0LeXCG7JBY8jz/xChfEpXxF
sAAAglbjTfeoNZHOK/LSLEjsS7oFrT7vWsxHpIuOUdNPGmRObI7AxHK4lWi/
L5rWnvmd7TraLFWoMOJfVAHRwO9Z5xUShMfUS+o6IqZI6AKhVWEO49Onsq8x
4mDkPHX6KZnsCnwnLru5SV0TDAnf54z8GjEEPicUT2Vr4Z++wk4sq6D+Iv+p
AGVVTs4RvOCe3BGFO3ppBKQ8s+8vnjFGRdqZ6I8tWEh2tb/tw/dYqKTnPhd4
ITAEz9dtV8cOKwqgQ8J8xqSDu4VmWcJHx1WoZZOBsqWS9IOj6x/ew0u+c2Sj
PXnwGu6epgbDcelZIO9im00u1sOigk+LaVe+de6PUrTuxiASUbN0fuVgMuXA
2+uNEFFN/Vm6RVKXxOfcMQdEpKmq0sw2EPeZN98ihO150AnfDE80snGJhdJ9
C+PTvSyihtcg+Lf6S6QuboKwPOzpvxqpYDH0xt8lB39MiT3qSbr+FtpKvrpD
R6rTWMoI5oVZPns8N25vSQrD5VfZIAhNX2ReNwK90gJzPPqk3SrJ3RQ2lGmg
QdskTyTqackPoWA/H40/GpKXc83mvbwIlPX8FWiRs2qUDUQ99BhCWQXz3INu
P47r5V2uI551CqIDwbNb/EkElpCxZwXI/VLrxMD6aeqVOMaTPxalCI8mZbjM
zAiCmKsKBirT27UmltuAO/DS9tBxqYnRjjy3gTFbHr6rWE035kx6zdUVoeKP
/GDNTP3D446MVnHR6eSx7cUYn336E3JSHOOGO4iN/Sym0Kpd29t65UrRZOLC
eoJhMorPhiLszEvhsARGryi80VwwQtaux3v0zKDahFykTHh2UOra2uvGe7I6
a5geL7j6zlrNcRaXl+exsmqcGHd+F29B5yQam8Zra6/0sPly37PtuFHtZosh
q7TlFT96TRviyzSJS5AV+bYLAQsU4V1KLDupyphHywJW9yAQ2EYlmMiFZqaY
3GV4YUIeWwqFqRg75WjeKC8WHXLHexxDyKTPNyJH5I3WTw4odyikmNhBIiNN
hHy4yR7dzUR5pJBxKYcnCb56kERwzzBUuVE6TPpJXpBwxSMF8I019NXxj/xF
gZN/YkpdWVsmWzSTvdfQygdvya2zi12Hn5VZFP2TAe2NAEck6W9k4QwTsEzC
lYGlaxBxX4ccyJo69FKb2e8qruoqOGXxEI5XwfUoUX07BKUDKAE878TLoDPM
6V5H3pc3Bw5Ipk4Aq9hf1LaaipyuflnrgTdUl+Mavk5FfM21jXsnBOyLwf2D
2BqBhO5CmQh1jXEyvMSUtYxES3+E7UfUDK18IEwJquJOhl6zKrEqYUwkkY9y
xKzUz/2XsAfB4VB8/EZePzkWTkzo7q1BMK1lC0bH1P40GO2KIJD5ja1hguE6
HzFrCoqMzFK4ionb/lSZv00jGHz8fUyAGNw06xhsFxI9SRFxAX9pjoJMfGUO
wA5/FLt1VIwF57IN1f7xOL4Hghri4EhtXItTON73wPf7Z3wLnLmXSz5Po99B
IWFbK0iTQb5qRysf7VTXWOMUeYap41k/i9NLMMtrwC+zNZm9vimbZF0RKZaC
ioIsAtLkxXOuv166hMzkxG/9/jyr4N2egF7axMpwnVpllTRY9KOKvGXojRuu
KyImce6/PE1HYbmOMyxc41piz/v6KD58eo9uktcLQDOJT0zZQeFdZVjnyMFg
Izi6l6jE//A+YwNmrWIcRzKWqOsefyqvUJODIA5aMJFdi8O6sqvD21E1g06z
L10Ngk3HAVRTN/ogHoG1BiRJcapV4XuvP8dwGrs4ACs0V6twbOPSPBrWoXR+
mpN3ebvlYQVIg0UJuvMFKDcBc/0CoDehvfSA8EeS63hAC5vBAZIpe4liAixZ
UQ/qZjOwHXV67MYqesHu4mnUgvPnSxmHSxIOHUBxUQZFTjkQd7++vWwxI1Qv
5g/B2MNKcN++vPwMhq8ZyWjGXyUMtFVGBgDgmyJqlcMgxFw77sDtplImYWcb
Rj8P/WeadRIFNnHPEwEnC8OCnY3LedDnHs1oKpnmLjHwvAWMU3/6332w3nb0
uAmrdNgzg8/dthIPSOENHQ5eC3JuY826HCqHShEp9ols3tDO0qNO5rjxjGFr
9zllSxqKMa5TtfqeRjyO5yo3EBPsZTmdMTzMRT7f5lAdUPQz1uKN95qcgvFA
HmZgYYeYQzPwXITMqnnCNTLEGQXalwS5jI5PQb0Fj3723UB4bYoQf1cFlGRS
ias0MhH9uoAqUlmWnbVk/c85i5+SRHUGkDFxFhs6Fb0UByvSeU9h7hohd1Uo
jihGt5dRs3NKA4ocUxnCPP/0nYL1xlU3R6lgTekoT/g2oSvueB6zeo1J6jgi
U3+7yEwp5UDi62Aze+PR/qJ2qNP1muRrtHSSGH7GobHflRz++NJg6EBfLrU7
lyH+pQ8mAGGBXpdlJbts0Z24ZW1iLHO5sDJPW8qw1Iv6ElpEpAtanGHqItBv
3iYj4c+/vB20cUD/OIZSpR7/WMEHoCcoidRnhGBYnFbTsKktnBy3VXGHzSKt
zMJ/0tw+ylkiGGwYefwJoMGQ/ydiMebxnoU5hFMIXZ6B4JbbefcQs5W2mJdc
1urzghf9QuPPhOIULfrcnj8Sxj42g2xDliTuFQ1e4AcbJDKdC6tfhoFPebSP
9/E0oJoK6356QovebV695zD1FRd0klJYprcTqM5JBmoD16GnoTMO0JxqND/w
mzgJv/decbC52IzHjv6D4CGaC4AGYQuVyZqcSbqPnLsyb5dvXQgOe5Hr+YS3
NNSjXRDbvMt1iU5sHZvJKKWYn/Bnn/pNIyM4WI9ja18MoSkFWV+n9aKv1wl1
BcS+tvWmycBnVkkj5J4TvOB5e5/v4yk8JkkovHZHMufgSS6JqIGo3/gRQXyq
eQMyuFqC0jYtf2FLgc0wtqnEpOQvvhI0v/P7IXNe6ZLrpkRORWiiEE2CsedK
TNsjW3D7jCRHlfp9LBadaCf1Xf0GKlWm5mwua/KOj60ME2IsPc16jrSrkwy7
qNVdVkrGGpZbjl2TzqMTeMi2Ek4+OMRDzYa4YiC4i/DOBnedlHnwnvKAlHDt
JYAdNl2OQV/IcBmlE9perURxH50Mykvebhx4oqpZ1bpWeXpv1iPgaAgP8Yyb
eAwp8FDufW6grHaarF/PLJBQiNb8RLOZ2qCp79LucHVQ0yRexx+itjvxPfg1
MBZdpMhZVkkbZa41g0JlsdghFz5r8MtRpz4N5Ai9wihbUfLMXcF5T0HpAN6L
gbaxKVczSqwCkoKU3oTPHrsBegqqnrdsA/zUJ5J6U952SUm0UrhQmnqpa5O7
wsC5c0V2SXg0v0/L5yXXEKltPuURkJDcMfj7oa5HCjahsQRePsrlGCTOsF3q
9PWg9EZrNlj3X+mMlNdTuhtScxKTFxzsJiliBBTj7u6ZOwx1x+rFo2n52+sC
gxVSJ89HOwbmzTHZicNrf4fuuPpShpb+ADSzE1XJSMDUklJdZe/8vvoESwgW
UFpT2wwBgjlLfwdQqusY3p/an2WnNkZdPWR5FW0RPo3zc/mo4O6dydNZ+LZQ
BDuCF4z+wkgUdALiHdnunslSl1M4QvI73HjpZ0mcRjfpzTLwK4LDb6stNYXF
Kvn8QrWqxOULWvxVOfvlroyWrSUaLexHKslnsHf3wU2/YfAA+K7I7SZmGuQc
81DqMem7t08eMa+860+4yu7Z0I10k5zsLWeLT7GR2kLhNZDo6mL6ZISKLgCc
zXMQ3UbV6gb7/Ih1mPUF9BsfQXQ7AI0Ww8HKcEznDsQ9UftJkrgxWTLmRK2X
CAuTvxQjPJcr8Zqqty9HI0yIoIRTug1d0PNpSpg6zmcx6NTVaQv4Vqgav6Gp
FIYIznvkWmyTLiTf/17uBVwpufUuNmiBWqCL8I4S1LnIHsSVcGmfb5ZD5wai
BpnwSSut0od38irBege235bdTLmiQF1IYaUVYxRdLL2eqKIouJwa91CYiD3P
6zgzX6mVWpR+cxda+o3ZWDEI4sb7b8XHxpc5tphAeE5AaA97avWr+Sw1yjjD
XlTspV17z3gJ+G3Jd+7l+L8UiNPllFqYySadG/dRu+2EioaAIAIvSEij1j1h
fJSGEHpY8Sl62ZkZfcDiKGFKz72uS7gWdEOBI+MO7Fr7h1oYAQQHcCLqGhQq
r6ndpFvV39NPHZmkmRtfU8dSlYPDNXHjK4LQFqyr39fMctEprO/YgE3/Y83t
13JLqVdom5pQGnw3cRPskIMRXgVTHEahT1cXXb61o2Nbm5Yo8rPFv6b90H/l
JWPglyqWZhMcpVmXIOwBZT6chVIm5Vm/ZeiEIM7H04f5pY3MNg1nEbhvDVAZ
Hnx6GWnxNIaqr0M4BMp+hEgwA4l3acSukK3UzvBx8fYwxBiTBZfqYvEN/11B
BEQLIMsLAfr/+K/fPZH5AdWTS7dhlD2chOToBsAga7zAfeFu17JLeVOPUcNu
aXJhwJt0w3dkFVvEQy92YGXctX08KwEaafcdlKDgnDf+GIUmuYwjwEPpGfmX
0ywRiGLQxARQrBM5McPE5B4iPEPiGU9rf20KbhPx6uhRGL0s/TNqw7VXKjKH
/7fCqZwsck2l27O0C0Hc7JMMkuOJqmRgNNtR/yevTxqDVMZX6tr7TFmrDoc+
ClBvkr2pZ7YAeWP1PzSdEqJD5fKwXnshat8a1I+MglHHCTV+aOIMPup/uosI
e38jcV7SAWGFsJrvMvDIiPMaqJE2kTOMM3o15iHk/ZTNQGXlrw8iUSL6lt64
/RtVM0/sZ2Dzrxm+J99FRJmOiicdQuduoKbmzNPbg7T4VAvrE0LkzHmGVk/x
lFnvo6UrsX0cMwznnhwCipdX+f8BHAKtu9hE6kYlm0kXqbSACvYsVrAmdClh
EuoYz5apcxD3S8ho9tJPdoGI8dy25t6vu3Un2nNZ45otNH3vbqkVbjPNUlVK
FcODd3Vxmc+Mv61398FPRpWdV2NwPYY4TSZwnX6fRI8j8bGypKKsot9gYmMg
OKsNpBwVeeP7IQ/p51cWVOFQvZ57wy2D360lA/0vRk7WEAXzuzI3pAlAf7Jl
xCoQoLgayClEptE0i1BIQ+ZofWiy26apaSx48S6VgpEiaqP88Vb+roWgdSXl
7fgoVqPV64133vwT3mx/X7g1s0wXXYCZ/LFKCp9mgAepuNic8IRVfV+pR52w
fOocLA5hiPZ+8ESqOGA3NFpmjxGkZSvE0+/Ur1gLCZh0LHwfEQoY0o3T0lyk
kYbIzFNE9eiomivYFC+4TtdXwZxKOaXAUoWk2fX3xQPHTDFts6yXzitTa3pn
1WTX3HrNlG0dcUvybdeeWGqpGJ62q3bTSTRmqJy88iIPgYX2TX9Oxv96s8H+
r3EQNx5EcSULbjf+ShsEtWKpU1oPe2VRySzaR8SQ0Pm7bBfKE66cwqrsgn4v
cVQrX40J4ERv9I2bngD8N6MIJXbqZKLB2iP2vgc4rpTFPoMSDQqHoLfKclkq
ARGXHJaO+iy3BQwkopeoVDAhy0dZZA9ptGtHibmi5Slem98DmQOfxE7CWYE1
u8V+i+7h18dp+EXWEQASHQMdvGzEjK1/3A9zB6nmSQvK8CN8HKOyFOmDMYxP
4OHU0ezzWpi/yoav6Q4k9bmGtpFHggyh/u14UKUOGr7pEoPrEqyMEBGR8Atd
0h11Zkhtr6AszPV24avaYQZUroV/8VRxnzfqVIZ4183yAJvJFwfjH9B4RE/E
cMbNyL7N3ktYBZ4Y7iZs282jPUqx3rf0s1g9Ur8G5Z1kW0OzBjZgj6YJoIcE
hk3DBSdHMnXFSn0Gdl5yFgmlCIybmSAPiWGlN+gMOEiICEmspXhtvA7F72jX
aJgMNrdrhRDk4wkDqzzLBbmNreQm7iZRR1G5s/UxgGNQj1dJPb+F3m5CSTtZ
BnTtMf7y+xBTdbMWzChNgBLA0SJiTyLlbMA/Cz0HtHooAMrLnzUyaqUAOwXl
jvAOBMY2SuXCYBcCwN3QLOssCPyAj5QOJiG0yu4H29NuB9gp8sy43fEORU7D
f3yoJGKAjAeqaxILxDPZzw1PamjYDa8+BrwRlA/XTcPAAUhiFWaGUHxX2OPL
g5w3d5aVLHTBl698zQrteaX6+n8lZ5xL3qQedjvtNOnsU/KCa/n8tbs/M1QH
EitOI1OFbIQmx1ed9PVPRlVWUqi8gqt86uazLiGZIY282iHW3UvbalYQStBV
nSw1jsz6OkM1l1OAkp/xkr/qKp3QF8h661Y8rBZtXtyab3nON2E1QNLLjl4Y
euLyd/p6Y0eUZOdITdFrLLuekhjgtPbgQSvX8ObL1ewAl90j9+NtyqrY3vM2
mL8lCB7/VX7vfyMg9VuQiifeme8iw4sxsvi6kqgLIm2u5IxzfKqRIM4qGxgG
e5gg7jsORwF2cezF4dlJwEPmux36sh9QFRGCyJky8JFDyfPJkqnN65v9yG7o
9/JvhoQ7s1S/DYfMjrpBc5o2d7h3T9io+mCQNIHMkIfO9OXTb4xNpfEGgY1l
AYIDuR1dMN4lJPUN6BP3owGWJTBAgZNlPDSFj20sjOjtIDvPyK3k0H+PIZoe
T1ytlFJVap4E5eTtSHKTyTE8qmjwqrTg7211874KhCTHZCtFGOz6flPRKvUE
9O/LkhorKKuuDcobSupiVnH4puDg1wRscUdEGYYpuTYcvJzRctZYtPVXsUX9
q9t+LloOpyn/KcBWlG57qhVQLSQgY2kSk4KUqGlvGvw+yLXNKl6dEK8ehaKw
3R4wT2SMZHczYFfGbzazGonCInKsYjhsZkiizi8qlG9aUYvMBSEx8s24V6VM
I7WE37+g9hoQQxC7SDveh/oqbcisg6lSmmovJrcWgmdTYWCNVuJS+JskL9xh
xFdRIVXYN9/ctQ+KzMIX+KBZ2khVeJJX7wK9ciwmmq4YqG5MUX2P6U3vfZhW
CP8SXh5N8YM93JhuMMsl5fUUKcHE3bVJnK4obDulXTj3QIpfR3aL/PRWNTdM
U46FHuoqPkh2cIghjpiS2i+G+4nPd8Z0LQWMIqVD90p40iwbheqRR4bf243W
S+6RT9jLiAEfESs7Dw3KAgfhldXc5Tce4vyxN4pkpFCyrZ0PM2rNrKddI9xX
6L92M1VEej0dEwCFuBjZmJZ5NMFhkcoRpmgSNvcmLf4CtlsreprWZvB2b2fK
rIzXpL8Z+Dg/1j045yXg952cjnhDjk0a01IPnGnUiNfy7v4snSghrw3lluzg
kguHVNTxlcXvZi2i0dRAeE/XObOGJoGYD2jqUgqUatzPmAYDSsiKgYKdD+nF
V7c7DuZ7Jr3Pdsvv5mlzxiIlx7XkqeqNPaU1/H0Aw8FP7ZFcenDb8n1XNrmX
GmMUMQHxWBJYFsO7Oq+LXJsghBmQQuK+Nkv9L1bwf+khnrWHzoOw+KGgVYpp
lIj0DAv6a7jLyx3tWgx4QBp6q9HBgVsAHOvaUlmBeSkPaUNdMfVwZwfJ53i4
Kp6ic7hlWS86W3V1HaPMo/M/z1kaBTsBjaHkQ/g4jCSuQToFppmKduz85mz6
kziAAV6w4h6SqpQCZli0B9HhcyqipBjxeneawDEqlknUxr1z7fQCDszBqgTz
qoPulnyuoUMLJ/uKWuMXghc05moV/pedAjSGpq0xb4u0+w+gdbAIDv0+IJwO
oH7s3U4n9sjWUnglhhjlRIrAb2ov4OBcKd9kVbZKZy49uPt3lfsNIQ1cTZCU
ARu5dBu48+rTaV0t/qx1sW/RaSq2j4sfM5tBx87qJ6RVg7N5sc3xC4wWoNLF
XaHsuos6X8ZuYhzSosedzDCs586NHDKcnFH6OMBxe7Am4IpRA9O8YdRphJM6
/lR5PxUSXVF7GNGtvbD68eurjiZB2Q2YvshGjPnP2z8vDIyjxb1PJ10bLnL/
yAXVex9wdwsARLuurI0Rzs+3u08ocVtyxi+pSaaGzt1Cl4xt5XuWrTSxiwjF
8Y/t7fgf/BLqvPcLXb4bCfSDAVYKldrhl+Napdp4IhxBqG0nmSUbfj4pjw4C
bJl9ljQda4wrZCXZge76nHef1JW8wi1JHuktx98SK0FjdTN7wYAnfRa/TSYk
G6MNcCWZSdTKcPINuO56237IFZ10U03VsiY3Y/K1Msocwmq0HqbQdkoTyt/o
mL0TGuSqmEF0wg87dWyoESF6FZUNr/BB8hwbUc0UKnZO4MPFU6LorecdjCfn
iss6/rtjuF3w3KY2AjsQaheuo3RSEO90A4eow2cdz3mxG/d4g2joJM4Uqq64
nNivtg0tjkHg3gldjhdDrC2Z1jiI9K+DTXTNLe9bl/s5x4v1xsN/SXIBW/f8
6+XY4WAbPgxusRvgHy2IrByUyHTcLAzU/nzQMuuxb7mWS4LnnzzzuKuV1ZEO
/7L7qt8/S+LYMCtWhXT160e+Tpoy2kkoo21hpojIZd460Ux3phex8ZQLWQUm
kebVWUSbDEvz588i9bzq2HLYDg6TpCQVEhVca+1ry6kT4T3CRxsNxRq2Pusy
XiF+cKhsBg67c902XlR+vp/rO8PI3v8E2YMphkkg9z1BjuJSXfaJywJmGvTU
4KwrOBc+0VXclQhxlp+HSBACTp63Wpd0WRFYN81BJr87jzGc3ScsBzWdSIJU
ZKBa5molemPhLsIKSNIw+DLyxJNZ8Cc0tFs32Rem3rniq4xd7+q6G6SKLpEQ
6+78dJlQkZB1Mil77OJKe3aUHaE7/pAbGp76nqWALvq9hfoFyBGSDi1oB95w
/+W3lSNEebRD3Cu+MnzQaxTQiD6pgP3WEYuBoh15/iNt1OK5iTYKpj/aYVkd
f4/j4R+RYxLy79FTc2zfUXg59Y80J6kl0el7csjrKwVHEpsuNAS+BJ6BB7Xy
JGd8X7N7pqAy+AZBhaa9xpGTYEVtuhY6EqbVWKlPh/kJ/QP24QySBzPliLHT
eDsaN2VnYvzo5OL47yz7fcVZxysqxMjqBpNBri6TBscQruxJdWZGcoWkVARG
cqokEf6bjQOFGV4ApPBP1mZXtwUdloj/nvmak5d2elYJjTqe0KmzbMMa5SJN
V+PPAsaJfnuqR5O8W/UoHcYAVPF30VV//90Ce15Ir144DDxFoFGL2o+VgL6T
7R1r6XbMfRn2/NWrdQOfoFG+EPK1KuqMv1FQF6+nHAnwoAPwD8BhP0tHVb4/
hntE7tCMK0DB5YXXpum0WOPwcvhDDiSdkMeyYXbK1VF6Gt9B5oTXZ2Fsrrn7
hzGrZ3Wvp380RoIakvIXWDVlk+9osKVMiQ3P1fhmnJcABXE2xx0eqVn3695A
YEKBCJPZ1mKJSOphL1qTij2rbvSJepVihxt+d6HUR45LHL9IXVo5j6Dzfa81
MupPalRtxY3rHMt2RLfd/uUCT1avaVAgdb2a+r8B018OkuCdCHIRADQEhdLo
9OVHDNdoGdXNEGJlft4Vgr+O1bD/e4VShirtCeOQoEENKqzg7B1vFSgFY1+5
Bf3Cw4upW0g9cT+mQIosk31DQZ6s6x0k7YgiE1PpmBk7J8ohwzzF5PmtX9Og
TuOZ5YYB+UJzU+VOBwvxPkZjlROHHPXDdYJ1dx8E2k6JT04SSIPm/kOM/Hs7
w9uXJ3JgKMpsjG5mAAAgq7h/pxpISP1eMZq5qN9xXF+PEqHydZvuC+PVpN+u
cd8NnqBdXa4pH/qsUOXi/hclImiBwgls/e78FpLQCrlkIWEiz0HBRSVi3PiO
kKiCOnqbSs8FN+IrrSMC/PAplLxWqS2C2I5XOYC6xm33uYo9uvbXuVuSnX6I
lWsPjAtLik3hFOdfuRMkptCAKXGPwUrdekVU+oHOmc3m8kEsrBcudiGJKJSy
2vyIYDqS+mmbN1o5BBz8PUkMq1o02oAk6E+MY8nSUGVxXHGvJu2IeE8cgBKC
ddy0bZlfE6zspfT/ijO6trzlgK7N5d3PQfkG1IXvjHB6c3TtfwbzVHewloC1
SrPZUb+PtghDh6BSEI7ZwQ8gpAaiUOhw6jOGGp/QNNSYnDyJBYmB+jNT74y9
I56B4J8yaoohicSrWezBsT3iuI4BTGivnkttTZBZdsAWlbSNML/DA5g9fUxN
dGU1bM5eoAM23Xnnz5MwUOdZ2jmcX4Xzp38bn1eONPCdqaBcZFHFKuCAZ92E
oa8dg1jSoTE7xyte36TSedYbcPXGrjFtafASfNsJ2pzlN4eFJORtc2LbX2X7
oYdjyOUemOgzigzbmLFKvaIwFuUTeWpmcmQdu2dBvBia7ubsX20Jc6AoqP54
WfydwKUu9ue1zuBRtYN7krRZ2bx57SVuRne2Mpn/+IC7+Ql7y0+UxXqU0tZv
w0+TG3cLgNOckV7wyKJGM6K3Tyw/hQDmrsflCuwn9hQVr9atL0g3fKWW6rRO
XEdX9mahLLkO4X/zC4cvEGbW8+Xcis4QPaR3eilwXsC7TPzOkOMWUOMgu3/j
hdfGH2oRkeQAvNcWtWPlN7S5pqIT8E5hAVMZJ5cG4DolWF8jP5VyD2Q2EdYr
S0djnDTfeCUhVrHFTky1QpWD2Rd5s0qpZChEcc/mk+8eRTdJ79Ien8d7YVTK
SZDHXY7kIcKEhQZ/FOaOKQbhqXYwDhB4ipketOfM+gOV0g2tjMiA6bqh0lDG
UthGyD5rCLW/W9UotHkOUT084DmTlOkEkXKGSn3ZG42xkXYYeKGT0lhiGHv3
i65HB3BizbSm1anqRZsQMh22FNy4FygAadDg1Yj+Efey8ltiu255Czf1kw4I
nhf4cXB3bBknddis0WDa6QQBQkxon76LnnoSL7rv4cPefnCgbfu617m2JjOB
6uVOOJ+3A0Qow+pTf0D1WrKNCYUcnSlt4DItYMC2q92QUGvm3Z96z7d2B0N9
P9w8ctYvDma3TLM7bxR+2hRK5M42K3uBHKhlwr88hefA+umQAYm8uFybef0f
ECK+lNCdh5HWeVo+TAMRzN3ML8evIf8SIRWjIv7Hy/Bes52F+jg+wRVJPf9N
0ShrRC5i0/dgVjElSdBMFe3AmhqiRnxRPJXHfTW3T/KMuRHParNn52fZffyW
KDgeexMha5g7CJEmcyUAMj84Bv0NMfxKeoL2mpBejsImCV4jXvLaElicVCOt
DejGfzFaVoTBT3MQtF/TkQdOKhL1ZBrbgK8DLDpcsaO8BWAIYaHFzNMbCuh8
213VHmt+NtKTkZbZZ07AFlvlN0E95VA9N4EGxVtrC+11OCryUdipZ/Aq4RGu
2Q9mjjGdB+IxlQxqKij6LCokhg9IaMT8xNbL6UP33P4Rfie63+6TPNJR3aWu
hNhTAH9w4/YW/7Otz9d3/hMjJMAzsfOaShB8UbJmAO+smieGISeIM8o9WmAW
2fc4PeAcxPRYatuCJDLUmggCC9fMrDS8HnK0gSc1DgE5QF4SGtV9tJtSA575
TPNSvm9Abr9RDuZ1t72lo3DvGgKrKAt16i8L+T+FHcCqZbcu/g5pLvegggdZ
vx937obf+JzVLrvrCPWEYz5yilHFRGDov2iP6QkIK7qpqbDZIC+iFQmdsd2W
PEt6ZtnxSzrIFKDgymfTIvljNKZ8EpjcurLjwdy8kNRUI2ctEvO17PDAohp+
M8/Lb4XaeLCWT7erZt9YqbpdD41iQ8Qtp544xLgNDL9t9akd2DMpuEWgyutm
ErLbj5p0xCQwkA/L5JOdSeEHZHw72tFDPy8KP5QkVmyfuchopzNqkB5Ypa37
a2r/OQqopseAzb80Sy5us5xKM4p8LxY0pmS31N4ozqnY2e7MOT8O4xw34XYe
ZG90qa2eCHL7A1/N2z7LNEeopNYxgDNvQe5fwfwxLGiVkjMnRj2hZufY9SHw
A6ZxRSX6Devd9vwzEMJBkkkJOfX2k/bLpaoFJXlkjOu0lysdMwwwIQiUDPWw
Lw1jUuMpaYHRQ5fODxpR2yIN6espjYAOeBHJQhFTEpH23nf67HwcHDqCsh3/
aXMtEWxaj+1+zi91+BNC/H2m4aicgL2i2kqvRNAn5/NHLoi21/gntbEP2CBm
RABTxwGfdWIvtEqDBDSH9NYrNgblkI+aOqcwI5KyKTFmm0JJ2it2uT6l18h0
uAWsyJEw/boNG75msOmijkLKCVm7ZreEVk+r1aAjHow2pxsJv3vY/66/f0E4
Lg5kivjA5Ip2tJ+efFm8lXopoenUtAQCOwLK/0iIfyCfk0DkFYvFu60YxB98
FF9UjFZQsy3BweLb8opmGQitJX2COdf00RapB+N4BldeKrHR8yg5NrlmqVtj
VOpyUtbE5dis6Bhd2IlDbKbLzyznzmDL7HT/bBvjKM9U/ikgeZGm625xLymN
F7UvESeRLfM0CmzgX7tEjml2R6Zxf9BzaeYqdkcZOt8RxER60eEAVAKuv1BA
EC48vEvnQ3+zyUrS/ycI/BKdddBuphklqIlsNFB5f3haU1MWxVWi/zgdK4yZ
OBlubA0rtzTAqpysdHuMZeE88ZquK5H39NqcYfzxCM/FP0A5rhiKR91HdNPB
W7LFURt9dQsjdfpfUXH5hSAombb0YQ/vo2gSvn/+D6RaywMqwbSZGs0+3YUE
P95AgkqGJgMIgucuXARed9qaYaepRUD/9EvaOsf156pTy3UOWFmgLMZIbQ1a
QE4xF9CF67qXju38iCJRlluBqMN2lVGxwZ50/3wl3F+wnvV9C39j/LTY5cIc
r6cR23hwk6POzscpe17vztdI6W7UqBPiC3yENTzOtjy+IE/iL1Yahihy92qN
w20PB6SbL6VjD7BJyf/cpm6de4Hv1QBBjSMXb+HvjWVUYM1oFdt+wX9L0c2T
HuMuBIc8GeTaS2KpMzrqwa0dMmFfN16btzvmGjRVH3plr7/sx9J6oLeZZ98L
lVrtqjBXq6DC0qvi/3eHnKCLO70NOdvnOJespLSJwENpXvjdPytfQKX3EQY7
825+iWuZijyDTd8EpLC2mT50Ko9ikqCrOi0RemPNBYJfgRkSHzoHRx50Ik7N
jK0Z9XcKFEe4OxSpT6I+4aDDBTUekRYgqfEsvXC/EJCAKmdVPPvn8oew3k8S
qGvwF8EkfWlandTr8/+LyYklzyV54ODNm8or1DILofty2d1TUiEDXBd2qP9Q
aLb37Z5AVxA0UBbktYS4A/tNLYTBmojSVPwxeMb1icNkxw8sqKSP7W7UOoiU
bBmAE5joRCH4NN+RbWLM2Nq5MqP5qJC7QdjLmHqawv3mCFcclhJyZYiST3x+
hgnJ6mZOiJ04hJks/aZvy0aungMHVHnqqla+KhD3gWZOK7mrScxQgfgvRush
wNg+H88qG/jle/iaGdi+v8NEh7ryPcXaoib0D0ZZSSqjKWDLFUpinpkeQyn2
H5ssVayx5P3XuKWIuAyBaoFS9nFMKZGXWTbksPpOnRrhbT3FKER2b+s8pE5t
K6zhw8FZBmE4IodDs9mM56g4P/nVA3zMtFOxm5EUm2hhqNPX/sLHp7Y6gdZX
9ZObj9KjFFUTxxr4xnoB1X0ASh+TKRogoXm5xAQdYC0a0AxHbd2gfZvU8T0w
EOUlk8Lrzd8zV3ZvUBPj6DOf85e+gvD+N1PyWCOUw2+dVVcLjDL+nZYI/4KF
6cLpfnjfqswNj9BkLrT7uyNsfK0AiPoyOE1yo/MPxh6l3BIn/RZ5DKZzc5Kb
96NNlmsZwsPPFDZc0oTs8S2ocTU0VwAeV8mWuP9gPqhSeee1G/uaqRVAztQE
g2mmpInme2yFO9i027BINaruVlo7Ng1fUjJdRn+M6Y0WeWucn3VjCWPhdArw
NJGYqae0CPLrm1q5L1791vTnVX2MLzL3OkK4K6zLYxDiic/bPR7TQQRF48wh
sC13X1DripuZ/DBSngttwCEZ8AzPuD6dLJmTpKyFjmpC30wEWdmpeHEmSFKx
I610QkeDgjh1VkvMOqUJ0qEGdP4QJA1tsX8Ynm8HiH7AwPH3+RTqbLnG8WDX
DvvtFd7M948GOXvfdKShrestrGFdSk9Tp5hoxNySPCYdHvPxkZdEYKDedYB9
sNtkRrdf5qhBTTM0CNCkU9+bI6l4OWXCUOA8dE1QwbgL6IV/n06X1oJsiBVG
QvjqeRAJ/iE/73nPEDOf3z7qLdYwdHoh3s9THIlU2eam74bZfLwA/tg08JhC
RgWikizytXwrvn5edIEQK95QCKLRq/ZAYavSoFQ7U9kMJT3zkO10GK4JhSK9
Ot79uGOU7/f9+cdtmG3KeO/9Acwi+epIcPJewCXYAmgwcoXN7QZEK57GwKvT
hXtibCnP5eccDiqcrPIGpaUlVs5vLZzLzsVyDyUw7rMuU2LWrpSCnsIDisP5
l38gUEOCewF9Pl9ts5cmjFfXMgXO9EzyLx8lbpoHueXvrXZkc7GRsNMQdAue
Cag1X5FB2+nt0HN1tlyn3g5sAd3Oks9fJCiwzW4Vn4diDMg+BLCrsFyWOAo4
uKkMbOF7e9SrbSlAZOdVQDGkT5Aq1wWGgM5oCCOehfr49i7qJ5asvawsMmlu
yMiezRPbmXdHG8mtdGwvcCFOdE8Xdr29F3sRsPzrSL6vUpNeoDqWlHk4ltcY
zYfGmUmPh7q073Cn+DzdBmVv0hfcE8PBIt4aj8PjFBiqq9Y0o+j5E/tNKzEF
dG0iD8EIpOHvSB4bGRHGP83baiCUswn7RSPQvlLg+KqkxRPKNh/vzl0I6t1M
ZxON9lp90Umw5HrFfgWepGvFf6moohGkZZhxkwpb00tl5Grvas0knej7gxkw
0O7dKoHXNH62zKRS+k+GW4HlxZyTGOSP3ymFEIZficG1SQvd5ePvxqTFXtpr
cg+jVLrpDYfSxkt2ywJy2OfXxTL9RBvg0FVegc2HfLgXhwtCdEd8C4LAIfdt
/yqJgdrtJJoTaMTItKdLVR7e6Yii0PjGef1aUog4d2tNwNRs7ZC16msEyorF
zr2CisHv1NSo8pcLBRy/BHvmIC/Vk2gS413x74mehYvRkYT/hWHW5CDmBLGY
dwoDPwRBVMkYQoiOWjguOESDSEIiGCU8m77A1vqFgld18YqCxpvAiOHl1bgC
rS5JYwzrElLcDLlxLJz1TqrvIejgz4LvrQweXPjeMQozMYl2gIzdqty/gfE3
nBhzzFqXkZWREn2wXOF+8CRWm95R2DaRS2dBy5g7kjezQLZlpzhdB+r5rDEg
tlR6YVTDgZpiDp1YoFLSgV20DmVYJxy8EFiWEmavoV963sQ38mXnbbufz7BF
ZZPloEmWpa8THjXUbOji2O125LRteYwKlc1yzwNl/wlWCb6mqHmFS7CxoUP7
QsJ84R+DduU9o13jMt41JuW0rz2mNLdM6kofN39Jcc4QYUtlHjamqU8GA7wm
l7hig7IpebdBCn6y8ADnhlG8/mgAhn+SDR52omiqJ7mEzRjBOp5ul86NSPPy
yCQpVqWmUXn8XQ0NTll5m7mqrofdk6T7YOwauMTWcgmud97Nt6s0xBUqUYX4
A1LrPB97oD+saGXR9ri8gQvG44kjcpKjmTeq/SmGd6HJPYMGsqse7dlI4OpS
XbKz9rP/SCno2i232Oh4oYyB9DQrSdXjnCj4nINnMuJPjfm6CarglwnsOV1U
V6b9Em0tARfl8BYy75Nz3ld6juc1bWJCCxdJT+jVHja4Lc1btZYcAQ2dVjK4
ZRYyKZHsDXu88xtuu9crvXDbP1cNNHAf6+Z80/zZfUpELp6FII2VdX2tGudU
csWNHhlUxL+e1Kv+MjIdglPR9PB/W4vLYl3Fmwn3/UiSEY/sIGSeQSWGWf73
sBusLtjS+Ky0UpwhaJNA9lcMvGaFDvZ1iIKrBPjWgBbszQPwrcfLAoQfK7Nj
CgahKAQZppJLK5tqXsae/99ECvCyHEGwwH/i+1WiXqwtgRwXKqvEAFKRuDU2
T7FLdwkAIz6bH+y6huCAcWFGtMymjiM8iAzuZZEAmsFeJTycSN6kY9cJwtFX
J/HzzlGiEjzhLNG85JsuSjITLTtWWB/Z86OfMSXcydr5S5LOikNvtZkVeUtj
qK8aKMqJ9TTD4oUPagg/MNYf8QAQPe12681j411uASJxs82eBA2lG5JbsejB
eSVti5QPoEtyqPIXy2g0xk3DsBfSIM9QdWNC1of3nFkjDiEwbxGNiUNKOqOZ
LIUW8n8XyzY5uzpllVZm50b5JJrTDanYjOYqWkOG3ZrLcDDEita0eZA5LlU4
otPUdAiKa1u7819i7aXa1WlUtvXHOpBSV4aCGHHxMTaUU+b9jCqbZypPwpTc
3ICnXBkccnOqVZtaFdy2L4N7LJNMfu82gjPKyWNnlmTml0WKwCSm35XTS2AM
p7CPk2cB+CbEmFzuz7VS7+7CSiZ7zK4MIH5JliXG2tRjEtwSfnISZddpjfHE
frkeFxQBzI57hcHxO0uwxrowvQrRz80EhYOJnI9JJQ/u2O8Q4jUUCBnIsg0S
MwFn6c4585AF30A+F7W167kRB7cbjvcf8NV5otU+rx1Yc8dYawuFdRHXs6w/
J8L5RVqo91Mqa71uoZNl2xMDrQYKpBWgPVQHHOBg9uZfUkbvMUA2ros1u6zX
LPSTxMTABALTZELD4byoNFwzKHEVV2itdYqOwd4vGk4aQR6L4u1Cv+aoguMC
RwbjrM3wyxaJsVkFYvY/8Oa4VPgF5JToH9f6ERsbTZZMFeycUkPQJnkJ2y95
W4vg/xmJHv2cklAcrmtj1hXJVDjx3q/xJCAYVOIk7myC4RTfwuEp0Wb9mO3H
c6OqvH+WWnYK0EmukSXbTrHy3YQwMwN2MI/wn9LVzZqxd1k5q1eMrPC53wD6
flBc6pITYCeAcD84iCHZtzA4Zks7MGJCzQBKzlTLU5JeQUYSrRm3NNQX79sH
a6KRlQ8bn773qSb7uBE4ElUBvNPuNN8WTj9QBGsZqIMg86cmiKvS+J1MatcM
pujKPKhIi0zuijc8yy5foFuB93lo/3Eg/6gVqPYwduj2ZMM2P5YDpCkOqOnq
K7q8WnE3Ksv9HfAJneT3YfHm6MV+e/dCJ5OIGUTDOK4fQ3ZZwFQPo9egUisD
6IFRI+FWBru8Znfo3nv3yzSuK+glVFEaYVt+xkLGH1RQVVn2+8g30CVKR8gV
DvKuPvoMkGBdRszop8wZI6FTgkMYCGFAkexTo5GhO7jndfn8S4KERz1115Qm
/dskOtNlVh9ve7Q5Y8pRiXgpWzPTbG9m2/nqtUolfHxOLSQe+83UrDM5oA5R
Qv1aNnjCZ5kqt5qQY+A7pn6o1pdeqaZpGCvTEQODcPDuBOutB5J1kSZ8GWZo
NUYnguEUZvTO+DwSDb1yjWSWp4z0IdqF63hRLBGp59RgABmn6IQbBa2AZLYZ
HjaDIt/C4oqUlbiicS+3sWPMMFB4QK/I1pygz1rGawW8lkaVJ4bA+SRuRM3j
YVn1wxfqLr7I2HXa28SUYgxEI3vXq05SjOApoARlkjC+sEFkCIQCfcgZvfhF
wJCKDgDX5+X8q2ysxirdDl31BOlXqOdNkOVyHcoG5WF+pJTfnNhGXnKw6rki
LvN8dVJyq9jOMoY0FN4aqzGk3Gz1rcgmVD56oYOY4zVqiIAsevlmjgNONUfP
AvUX6I6VP+dsNL7nJwbq6Drg3mMnD5z/KSkvctxY/5FgZnuUQkW8swhOvvoJ
pJ7mM1g44DUK/631VMt0nz4/cCt7qCI1lmRzjFo62DOGpXnAyPUhCPU0DMvt
Fj9UEuUfxm7AA5wSvuyVIdUrxuyWlmSkWK150qZPYe+iA+YNQpspLhFNzlIW
zpuNnqA+Jsvqe5/Rc+4/pVn3w0Uz8JR6zrhg3Vvw+RdwiDmBLR7nq/VsS67Y
/wC8v3sFPmCVlKk9d/sbUGOEN3wKUfJ3e1TX9I58VDgunObNmzuyW6JeU3ly
0S0Wqo+MljNNzxS9SpXtcCrqxEUvJRlLavQdJMzZCCin4EFJBMdw3CwtmrHe
Zj8HkXUtObWfwIM0mFrCU7IEUgrRo7Ai3VyUsvl1TrANCvN99uXMWuUs2EtM
Ew7OkGbcXsk7rAQwHevAe4oZ2sejVpbM3v6Aant44913kmAn37QJLXlf/UIa
fYPswtsG/qTnCKD27rjFhko7YI019yhLwVeRk/ScWrasqBj4czO3ZW3Eam5y
whuvyVkuXPV+SdCw4MULa1STTU+0a6J41a+oY+UwJ4cAAme5rUlxrwOGw0lu
HKIsbfQRuzhpF9J1ukE7q5/cHGnjaBUhaeRybXneh3wvyZxkB7VDQmOVwEBJ
8zLzZYk/J91XhecbwkQPsBeGmMowNSrHnU6qWadM71RwTOyCHVlWf6vTEpFl
7xRkAqSHcJBxtTkKpEwvW/e5CnQ2B4COfI8uxn+0949RgUBftsVHGUekPs10
dISPAYrtDVMkKpQGfUfcKqIWYZ3PobqDALKGQwrLwtFqnWHynQkrLSmKGO6e
5hLvVpLLeuIY7OMcy2PXThLVObMM8K7erQKTFOlDhtM0jT4Igfh4d82V2jxX
+Nw0qb3YXM0EbZAo9C8ranvYDdLYH26TLCKKidvGYgmQeu4zpuieVaKDBGzS
S1BSADjN/8gUis5oLkkfmfk6G+NItd6E4uKF2UUCr8YPRmks7QU2nYNABZJw
g+O6HGSQzpJNMBegY8hamhzUlLIyWSlkXTMT1N/iES6fcBl4N9ARDDSQvJpH
PxmN7UKGYFLo3QGP6XRpaXmcSjqqOpZ0tHTONF1cs0Q1oU605MnPczyyBn7w
SkBk8WN7mu6qz+vjRdQqZhNy7v8gGf1dma7GKFG2yJSFW0hFcW7WJ/FyKcpX
hjpXzxGIKcjUl2vpHzIhTIbuIbLOKTxgFxPr5iPx/V1uUqNUDFgI3tnC7KpT
VUcWcAJ9oNCzTOVRKNbxEKE5BrVOOs6GdFzVRHYau+RdGMohrk0gRKKlzLSf
+rf+vmR8YTuBEVqrkGzRaq8WYVUpOsyBkn327dQfvHOa4Dk1CK2rsfdKEmrV
7B66IkazKV2RVd2OnkndcQ02XkSeSsyHXviKGXU+g/9zFAY0ssU0HwiS8Yy5
BWHkaku+C2A3kfb21qbPjiQ8L2GmjZnt0ylpFM4SDu2AuNEafDSsiEMAHb8r
gdJ+Vv3XHbWiUmaxj5uqF73/vsBtvX3pBNhfmKP66mXSbDoABSONGY550P3p
M7UCFlq2EcK+yktrXn2FNldBWBXux6o6vYPQkXr5ekXHYDcBCvb9bXBwkwJi
JDSkWwqkpbJZj84CZ0vAFvKoue6C2QAG/XhNAB1pm9C0yz9I6zRHNt9Iblxx
Cc4xQ2ST0baecz28NO1PY0WFkKQDh//e3EMBeZgYn/FSuFrw4V5gNZFKj9EJ
T2ZMyJeB1PRwYDLRme1LnecMTMv0m2KBEARkM2A9r1AP1JQACDrgejQzixoN
y6LX+gfM/e7b2LgRVso+tnGdln/ouyI9STDtsYb94BQcW84eCchB4Wcni1+s
hpYm7RCUVUN36qWb5q+5YoVdAK9vNbzMDg4rRKFLQWYTCldeKngvdQRehdhF
pP1egNCuIGNiC3qrO277LjsGRntnWt96IubQROc4QUNzHq8Ppp3ByJUARHR9
v39XhLjgsbeVJCFao9RN+Nfq6cT9KrAOUJpq/PpvAzQ5wmrh3eCdZsBHcC6F
vPbzks9ERAr7oBzzmsp2GghV4w/iwWgy+sbuu+5M4mcQEoAKcsU7PzQE4uqF
umS5RLLF/PdoHw3JS9qwUWuLntGeM0c2RIdYvd1+zajY3dmY5snEAbWz4Bsr
b6om8AFn2S16zbFPbOCQCBd6+nigHaw89wZuuqdwpKt0cRjJBiJs7SOoCpT9
yKDE/z4AkPbs2iHnn04PLGhEfor3NGm5m9LqdvktJxpv9xkuok8pIfmAXnFn
pd/JnC1nbY2vvBrYl/MhCGkcyIgAPH9iM1q1KEPoYkuei/aYS2BOs387mMfI
S+EqckQPeWVMnKPLudmje24eUEuyNJXm3dPFuJAFgc+6cZjY3oaN4lewCopH
cmCEphSccjivdL5nn8ARWp283XHo1887kY9HcGPZ+xi+uAJeCYqZdLbBaKMJ
ewIvIo2EUrGRh5nGmrh/RSv4eYxhFVg0XbuuM9RAHfHvOzXSJLqOsCpLS/cV
2eiQLLUYYMKAQJSahHkfK8hoSYVL6ZoDKKzUCGtmJaeMAXcAwrLUtmtFwiPe
m1FnIo9Y1pxP0bDRSHbFM4y+hVxvWSLb3nYnxF1VMHHOn/fUf8XTKsoT9q/S
MJvM/pUp3tAH//DT8bucGpkpVdyXl6aCIdlgtxx0nn0e0iJpnuUy+mYU3PLT
bp3DPvYV23n1vyI3BlgOUvgqBYZDvmCGPV9jjSv5zxad3dhgXJJZ8l5XQtsk
BhnayrV2aDgdqOB8juqp5tZpw6xWuk8+HsZNzBVmtNCV4TEV2X825xU3ZywI
SBC5VZjVLd99/2bzmkrw+E/P4L/I/K7Li0Mwq3lhHuPz4PqudJIxlvVUmVDs
7g6Nn5drnBbpi7Vw/fpmPnFs0WTHdZ4KB+KgMrwO/yIeQZ/mADkevwI1NgOH
icEqQBTzl5dXdyHWOZM9Jb+gt7TS3MJA1VPy17Tl5hIg1L0U9FAHH8Wpfi32
63x1Najz6tIhNkHDbNs9qn93y2zwt96C8nrvxe18o17tEdW3s1trbj7ZXdUp
OfH7mVj2JQVNtX9gYqZJlrWyQIdZe5Fmsk41/pXz0kANcI2OA6iRnvBZxWZX
Fi4IYOOqNCAoIvM7X2voqVXG8t4lb++GebeTU1NAMCPrcWEayW/lVPdMS/Z0
k/lZmR8gBNMVZbrheCUbDPnghzeoqLTSfqgL5Rw/jSvJL2s6ZFZuxNC1qtGf
zKDPvvhSWzl7ospvHAFD4K3Wfe1kZ9TBSd6pmfx1zb1E1CJyFVF56iAdE5zt
jlwcIvPjY/M/imXMPjzy8wUdPREI7joZpLn/8QCRznMAFoap3gh5x4cl760Z
qRpjQ/PEzS/dIQWH5wu2nFT/zVz7I7vnG7waEIVA7ccks6thiRaFiet+Qtl5
cM6PJ8v4UZmX51xdR60uRRLYZF4xOuKWwYS7dl1OLGFzImeM13HOuU6NZ9jr
c3htqIRCLTsubFQ4YAuKGKPn5cm39q2lOy3P7hnuhBuXVzTs7+H95Py6yhtq
pGu3UB3GvcVui992ehPxqfbUgXcpB/y+NO6eZZto5WIZg1vZ6pCR56cHvpqb
9hpcjq0GjWjBahJazMo/AKphM5NKsaP3r1mFjtjeY+REwn4hk/5SW5VURRWO
1BgnqVcRXV2X1UkH7txz/BhiNwZbRWL/TW0f9Jsd5xcVYGLCA+fxUYMvL/fS
EYp0Nv+pIegLY3BZ0X5zS7su12ls9XS+dnxPwy2pzvxHnnrCq2/xhs9uHuBM
KSjBJzFFRqx/uQ8klAIyZz0sChwm0krY9QaV6WgMG0DzCHCgQO3FhHdGJWmr
qJpRqm0axIkHt6KyVGAkTrce4E9lDnKYKu2Ao19hkIPkX8ucFaDtyTD5zeFm
QzNXrQ38lIct7P5D1/OuOjQKtfOnhu3tANVkcNizYik44CZs8mAWySAer3CA
Ab5Bc8/KyfrOpJgVOChOoldfyVUHfuEe9trjSrE+1GNpqbQU7ykif+MjlUES
sh2YxXNkPWcj1F2ReQFmQpIzcBgc/EPfBJqb1Y+6eFcQkX6uqYd4smKcEUPA
ZxiYjQWyLhIW6AldQmRome3/ndX5JH0R+DwHKbKLPWH7Mi5te/hJTjk0/KU0
FVXvCCaQwpJxHbvAZlHaL5GiybZ5jG6kHEshvwxugJCSV7r5STjKEaheV+Nz
YnD35LQATSnN6YfXcdkFhPMY3SxZU1BnHQfb38IMT5CJ1QrfQmIo56FyZ6qM
WWwELoQOcHNl4SKmbcIPu3OMYe4xMmsnLPvY8ildygErVgcpctu8x2GSsZqj
0FPKaB7ueKdBYJ/b0mraJTRNb3NvEN7W5UKR7tuzFOF1yz7JxHrg3yikGltO
01CkqyxFwvGHOORCDn6ET4WPq2hIaDeX9yrHk5O7JOX9sIFydEWEe+l5OF9L
J4mdufNnAqVpKNXyfEqN/+ADGvHRdHEeSU3zYkNYpuMcar6E8D7qkDkDiTgW
YR6nUb/sy4RNyty6RXBXBriyl85MapGXT0X6xeDye1ZGnQBnesplCHRlw9mY
R3N53WX7F303O1Fr4a07u0wecn5a9u1ogOSt5iwoS7gLeLAQ6dcBrhXlTgWY
VgBM3KkhsFNXIOEnlxrxRRj8XezDOHXPvvV9O6t9xI7l35dmIGiSfz3VKkkq
taHopH4uKdzXoYqCHOXeCkaF4RKeP4M0ketzlRGjhOIdDE8UPiCfIVctnis7
fYqjaoekyY1+IEAZwjwq8U5peGqgzMi/jX7FhelMygpDeScerTUGGUPJZDCv
jg7FUlffhA7UKqzA7rpoMYAXq9ggWXTSITG2p22rIexI4TVMU6WKbsHD3GGL
Enj9SO8OVFrVo/Q0dq5+u6i0p4kFptoYRkhdxwC6btjfn5uUDwsUrJx3LK0d
qeEWKMDOyNkV/dU9NHsfxwZICP9cR5ww2BSU+X0BpiYiR2nYdS84Wjp+yCi6
1LyFwsTiUKX4xQH5SjBLLomZcNZHI6zu8ARMXkESNs1iPX9eEWhVnqhJQsCA
IqguW0LyhDqfBflJEC6WX4H7yHnSJusLzkQhw0aGYfqMcfjYh0uab1GhHemu
lbzoQq3Ff0hd2YzCeQ69OCJs0pZyNiyFsQXFsEBnLQcYQqu6iDocrDbq46rf
ihOoZmYEYcYBd4QaDkdssjonMfGvCKa1i3TldkC7AdCeglY/SEzb4vsRViEk
MLXv3xegm7ItobTFx/sqkAimVmpUVYOt34HdxUmFTmJdVixLt33atzYjx5AB
Vc4QtRo29PVj4sLL037W6WpLlR4VLUX/YlErqvA5M9HnXNzMlXAHxygL9N0T
Y1cRYeozY8ifM4VKvRvZXxQ/WMmXyBnwGXGl7f4qYMEWFKQvryxy5OL750oR
4xzRaC249XY0o2MAfVz+zOv9q+lh2EBmt9KSEVvNlH2JM4e4H+haEAYIlVYG
hs8oMM9Gf7Opgnj/QbSZPFWYfXtNxsauFrCAQhdKqwBmvobYUQUKrZTLyrfE
wCkpZ07Tmn6IzZfSDtYnQGW9P1EeHiZLQgGJscd85gGusyielgLzgn5z0JAN
aQB9Po66V60hTpZ2+Giho4NiF+dWpU8zez1wn58ttwBqfmHC9Fwfh+cll/FN
Nzqr2x2Oy/Josxyq0cMKCMR0TFQnyvobiCuiqfFI3tQK4Qd1xG4Dm2Gui/rT
jIVdba/goXShEG8VHKIwroknJ+vM9rmZUSJwEEVlIKtUtpdNpRFzGlSAf+87
JqIB+qDEy7q6y/RJ4dr/wUDgwheHPoEeZZHD0bk4vblZbs0tnNCJ/Oh/4vAv
7sjepulBRCS7FuBO+Xg2VNR8tocuLDL4z1merbTFQ0/S6RTS4Xw0B0yIg2Sp
sK8oKUQaC+8sT8Vb2AZHK3Q8ax2B40d5TIresAqP5ftnbl+Rmxkea65aeklP
88qGS0ASss2J0s5kJ6T47X89sshyIHpB+U6A+lh7s2K0oU2P1/fz3/SRPS5S
QZ7guZ09Dcx31aRWbGXZJS2kjkRagwuQRaHa7ZV7Poa/hS2Dgx5BMcrPxcOw
Ckfv+CsMRh99V/x9lM8Vqb7u1/88paFLUb7FqLPxAesvJxd/qG659kMwYvZG
dsZTJDmUwzXkPWhPHDEmeEg5NkBI5+fTXv4BUYbZL5MfOSam2lrSZPM+mkTp
pp0LC7oazxK2XeYvE0yVYtN2HM9OTZ3TEj+lXVqe7ksua8l70ovhWG597cJg
BLDGOw72nQdDe38ED70IWMDixsLJp48MdtGIrwHuHVJv2FioG1J9U2o32kkL
aJ7mM982HMBKR0bbzsJEbvbNS7MfICkGNp7MVxm8E/fIh8ZoYr3arDZuKKqB
hlTmUmFy7N+3wWRSoo5dhBspnBPkjJNBly42EH0wMDD3mBrgxOL/YRtvfo9G
2V/Tw000ilnIgmuUKfk9PTCpzzRaj3rurTAkWY+ilBtj9PSw5YyYEW3Fc9st
OcL6jRlejuAseCDzdTmHn0AwpQMKBEaoqNiD3J1kZ5rgN+AsvkXVMhmG2ZEc
RYi0t9eg720UMaJaVmfv/8CghlRagB4NUX1g+ZVB9+46SZsGwnQlqmqV9GmI
74PZq9dTP7OCxab5X99t+Hfe3uvTPsh0QlB+XCWt7z6G4B3rq0ZHj4JfSo8h
8m5h5Dd+B+k95QLiSydLdAJlF3XLJ1gAmRI9HFPIXihgN6rg8HLsgUjUEif9
G8z4HqAB+bPkf0ZY2FjdKLb/ZobKqSU7/0TmCllTcmMm0FnQDPZuJQdgEdXi
Z5lEZUpqGlbF68nT5+opHtIrDRW27EZdZjTPVuGDVwb+1n06m7uO5XpNVkdP
UGGGB5BOTcTsFP7mKeHCwDSrlNd/Uv35knd/+TT2rVxWFppWQ70IflSYMzxm
QIUetrf0kdt/H2CCClTp55F2zEVUuLrjU3mrJY8wJXsPFMPlTrjNlbW9pzQD
H1yPAoxNyx6O74fRzQEZBF1u0lJOvlpWxRfLNAB94jvYdbdPCz9gpB0k5rJL
3e13IQBFi3p4CLPadCtQtD1uOJ+kQjJ/zQHOCCVHG0435w1zkmun/4xdXWO7
BBEizcAiq/OQWIKgqtGtX7sw1/Ce/0h50TFUttwEXNicON+2xqCrmpSs+Fd8
R0NmdF3aMy57K+JdreGfm1QL4rS6tvY0Q+ccSmY+b0+G+wJx2xf9wLS4IWeB
FvlyxViEMf0b/wVnJ4C51wnB0RxfPchg7lyVkl8fOh6paNOqzyD4S3Vl+RHm
7a6e+LyGlpihT5oEpy/U8i4ORmImk4cw/TGGRZdWMSbeD7Bwr4qefwjZs2jr
kUFOgtvzae0UBTPDuh2TIMt/we4/H9QkPO65WyLvMdtTB4RKQEXhC2EdbVuZ
R3ciqZrsfDXwXJmITNEhwuJv4yWL0sj+HRmjnK6oqqnr937uY/uWAQpEAdnt
9KVyNDS7bgad0WXtJEBqxg+LqqlQlWc1CBw91kbsHTeLbu1T8Rlktr6YO8Bs
h5IO0hPefOg2QIGaZLFdMCMg1ayOis7tHd7vVNRaorND81nuOhZ7vjq0hNYR
BMRKFdfd9cG/CAWc2Xw60+cmeXS+3y6cxGmDqq+ej7AKOvYePkKEToNvMELN
Gg3oqGPsbQTng3iitjdzkf4MNSPE5dafMaZwhSv5nWgpfWk3YWJOnUBz9tVz
upgLV1Xvs8KlU3HAgmmiQ1BPd2yM5lhIBN5vBaEWdx80xAdpsKiAhVcp5J+e
ejjELXXIEfn0T3c3Xd6MIkUiPozle4ycgoiQAkfmk/P+GL1oSgRZ+cCWdcyN
e8J5Z3suUcssHMlum72GePdjti4tlktl24+JglhepoWy8g8pn88vHtO5RKYQ
O3MzR/nb+ulaSStOiv+B1Dpn0B1mP0k3Y0aYIs6+D4mSuqxPy9OinPAGRGwW
xdTPGSo9WQnJRy/JbGokdooLPfLRybNMxOZXFCGB3oeehtw2uApYWIXBVoM+
JyjgCZOu7AgD/zxnQtuBmahdYkWeScrGUu+8MSuSN2nXyoVduPe5XcjdUUVC
wgc59kpanzIWfYW4B0RKGITwL7hmzt5bT21cl0p2QxjEc3Rfy2IrpGFvH9oS
s6Q8fYrSRj1ARHrdfh7tD5PkJDgbg8AsGRj7TI4bccAh4LT7yBlw6xBc3HIe
jhzH7o1ONk9a6nnua8URoAdm2/0paCqSME1E3mWOqk8VG3EumvPOvkkOcUSv
kqNbcJ9/nNl5IeX26oQ0hj2SAtafwJsFbN7yQhKgkTNQwD9ivdffvyuCVjcf
R6QpKaPwyh605xuWAVp6NuAyqN17/eyEF8fiAlma1oC16WEGVRUD9pSox1er
7Cg/lKS1B4HLXKCsAKLt4dJ1AO4xzL48rC4Ll9brnEtYxxLgoDzTKmz+VO+q
rBgV1bA9MQ8uAtedt92xhz1b+CTRH9qBTu2zbw8ll8WQ7pLBMb9GR11qjZei
9IGV5E3Tg3vdnPt7GXT3xSAuFfSqZpGxA5cB++RKuNRKerld2EEYoY3H17fc
sCX5RUBQ1KTtkGpMaemHH40/C0Lh3D1QBD2bzOI7UQpMozZV8iJQscyW9I/o
xJ12y+R1czlKHAGrr6aWJV/Aks6sUr0Oa3Amf9JS6p4QLBfQuHoi11+0XcpY
BLe3RUqjQ3Icfht0VpmOrsYITypJvy6On3QE9wCuLDFfhuSv43wHzrkZy7Ai
khDqQ1cN4fDCEvenYOqf5qP7V336oN6UOoGgTPtNXr33KaDAXEE3CiOhG7Kn
BI2VjgMQXDK42Kz2/L2LSu80JpqgbukCbabWJsFpg8Z7ryYxeRESy9quT2Ky
NJStnGZlBvXGiQL2nwMm5ZKz68aiaGcoxoZFqs0RVDCSDdORDA0qp554htgL
96KkcIDA8jf9bVmNNVCK32bswBS6E1Py1SfDavvA9rFYupHT0dlt3UTyUAlb
CgWljQ7JrxQdSVe9ZVMaip0FzjHPOWyGQxhENdoFgpRMHvKaTjSG2JzPeP1/
+yjiTSibjJZMdtSicLBDLIEH45BYLiegfTv8wUre5GcYEzwdZvqA+Kb1UWb1
MqpdktKftp3ZDjukgXIhCPEfKZ8RUbt5qDLmPs6LLG4SY6fhrTUvAPKd1If+
rAOyhLxZTDlYxHePrWO5r4WSTWcCSIG3ftPuNnhEYiyLNI3xMjkO+jklpIAu
bgcL0BqtK/LHi3oVj2q7D7wjoCZdjGI/qMD1xvKWFWAazq3E7d9D7BczI8qs
0o4e0oefXJsAUGVOAM6YWB2tiKh1JhWx78rXvqqPiOI3cN9y6b25+tlREbY2
b8ey4hCjSavr89hQSu2Z7m46AiaQi+gvl2cZVtV0FX8qA1EKpuqvlEFIisEB
XAgcHs8gYfV20kBY7vFx7mB6OuvjGKAbIrfVVPmqplkGXTivZPAZtkQbtQ3l
26c1tujzhIxr5ARbhFqStRkY5EF4nBB6WGILJnpz5YmBf2GG/27MKlHuZeuW
CBy1VQl90darHFxwbTlZEDuvsj1bjiVQCEVUbX0MqXNnDB7ZVi2cDfX4ycJ0
qujWC0PYhyFL0ZamXic43W1nCeD8usSFR3o7oOVQaww3D6uVhA6HrGqwNfx0
0VrZVs+eDkqLR0m+3PWNSJjD7dyMhT2jix6ixLIPUYcHX3Fw7MRy+u2Fhmji
EzgX3qT2zVSSSEBYXqAYpdaPksFmT2AAGg/0ucyqvY5BjJyPDLccEvdH1top
QUynCfriXZcFTv/NzwqoYeUhEbgglNsUNi/lHPJNHC+W5IkkxlYWsUK5nDR7
chMZt8T30s/pBuasBGOFzEY9sag2E4/E5mi3NqL0ixfkmCP9x+o1RDQ0bx+A
pf3GrWI+516AHDVfxDTjOSbm9hR68mmFvt9wGuHUAq3pIofrtRMJifSJ+1j5
Yi0cwaJDhLwVOlf2WH8mvb1nflAeJLwMyQ8QFhiv4kP/b5Mdg7bIgyCsjsW0
im1bPDfLd7kGZno9fB/0SVA93d5+GzOV67gZDfuyDL2iOwfFG3KSqrPGYmH8
lJJAyhYVXlpFYFXxQK6dgRoWatWroliUxnn5HUF3ut0kltrbnLPr2pNF4sZD
wuImXkfbr8uZNB2mcuMLOYLLg+TJXWx/8Vld9hjru/ACO5SU5sFE/n/HATnK
EfQ4rhZVzmoII7SNpHox+Ykyx1L4IEu9BPc07A42mZ6sMwo6OAd4b10LRxnU
aMVeY+sr+EeY4+qQ4A5DepiKrL6DuBl6LaT/NL+hmva/KQnVEXGCW3aeG3ZV
cpy3Nb2HIZgeVe1uc7rd1Ux+5pxFYjJYrnAkRO1Ys/AueZvicU81dsaspVYz
r/MuskMUYW0xSu30/R00X6WLl0ZoZxj81Rgv2nXMXe616bqgCEo/jGlxec2+
hnzNSLViiZ3Irn7i0uUcfEAo3f9mZrBuYm0etqNziWBNC5KjSc2UF/0SHjoB
Pyx7bUnvSvvrrd7SnIefaBsMjrnqRdsoNZnd4RoUAraUGomER0EX91D6BFdL
MLrPV+rmJhcWrohKkVLeznvxvvKe7NMPBvsd6t56gcz60DZbt98wIi1SQQUq
O5kXA60JfF7Dj6nh8of+Nwi3E96/Hehq1jctU3Hf/txfZ0DZ/WkEWUYNx7LV
GdRrg1LKf+XjDYlLpLeJDtcUvJCeByoWx2scHZ6QiQxRhKzbIsCbjAVZWQPZ
GLSA9EDG/a3iIcZNmSJg3Kk7jSgW3HW0Jjm0ftepNtvhS079F0lB1ECmr2Nr
QgHI9K//zVYgu37rRuFl6AYbQrAv/36zhjj4uSP6YGaI30f4JlgTsqUQaWuB
8D0J2PnuO+CN8nw+LRlJ8AxoU+KGJbCCFssGyo+J1YZOYHpprkpkavTqk4VQ
4GrDRaPOSjMMY9QqZpwCy1MWY2dSE4ejxizUPZAC03+UYBwo6Deou4E+7n5M
4QHYvTP05SNV1xxVL81YHnHPUmbXlToPRLJTfT167UUsAgMTNyO7crYN89r2
c6zB7qY0TvYNwvc9U6Tt+/nhsRzZier944ntk+r1m5vGhMHH+cwWzCpkdVeD
6ziKFhy9SQJjevIYNJvz8JiCDzPAp3ekfWF3MS8ljdXd5bsLeyajVyCDtMWe
6IDv/ZwJsWbAcw9WhU9FYMBeEtqOOUPK4dRjrONSxikde3HRhgPOjRQ0/Qoo
rBQcBXBqo/g8x1mPUxyKwURluVF2JYRZBr+zuKsL8HRlfVPR1r5nMdiK6Z6f
kSCHms8l7BlI4r8rQAZGi0ztLHkRkM0Nqevxrb8J3MqWqn0kvLXUSwbjQvMA
XTsAuBAlSZy/52VTTVNKp4ngHd7s9naMGPXRUE1L5WViyXplaAJ2gTPn1HxD
wgjgnFCNh8NEkHclt2VgDViKwjJUy8wFIlTtMMrzJQDwDCfMKit1i2QB1MAI
RCNk2Rq3zzvUhfonDV61/eHGZ7QQ+lHblFfwiEFgx86A5QYXe+WZaiOYuiL7
+/3WbG4USpFvEDViyrXIup6wvT+fApghk+YzrO6+wPoY8+OjKS6/9rfiXuOP
kQZje8WT79ZKM3ILxkxYMXITShE5AyCUI/L38A8K060butQlq8vh99MWpPu3
bOBLwckFruD1xfiTpckKC4dwkCaa5nQ0tx1LVw/oB64PWemmxlNM/C/EazCc
3Hf6IUu02Zv+ElaXuIgIVx3hMsU8wmy+tyK9Hl4Pi600ubFv2CzYppPvAu1q
ITuOMFUXd2nTybBNyMgNX2RGxExEKg51apqrl3+397uvLRyJnR5s7WCHqN1H
aYfPQfddLhvkP+DSP9M2yiFcu5dWLMo6EY1kx/GKauBOsIeATHcBrarwpi6m
f/BMuG7XYIoBiXkzD8szLUOsCqrSUwmXffI7hhzNXosIn8JH7iOhkYRMzbAC
KSb4PIx7E7E5Ex7y5CbSbN8cxEe7yRZBN1CokCmZZUifYu2UgI/WCYPZKPol
FyY6lvnizAzUAzY1j7NrK3I9spEvW2wG+4ZvATZrKl2PDeYyH36q4hjoxUSP
sfU8Wd+kJaXqS4jt10DGUf7D0WD6N/0ev5VoGeIwi5hms+NPaTqOSAG10T6/
fwC3b5pjc520JDGOv5Emsx9HLXznTHaPqZJ0c5vJdbbKikeq++QsC4tzjMdt
hFdp74H9GMHq6Z8O/1xvhCeP0PR3KuOXgTHBVpPIVm9RLMBwo1xMaIZug/CP
UH5u9gjC5Fa7WDWDI5f0V6FvusRwinK5vfvpOvdo32I2CsGFs6UZ/fvh84Zn
bZ6JpOsnVYIUtlVONglYzTGh/SPMiy3F5gCgWi/cvdUIeA6ZQSU6ooenhBjj
yAMoU5SM8NjqLTitmgdbhWNiVQtWmPxm7mlnFx2GzreNJh2vNJ4DjgGgWKLE
tTgADp+OcRSyLdk/MgRjLgje+a+3SL3ZqlFaL9TqrD/9rYPDwcNkWT3tCwyz
juy92YZX8PoLHa/ldor/RrOcHq25U6ArzDSes4h+RaB4HaDgFC0Njki65ITq
sZhr2WIwrqFb/G41kLa5j+byD/fh1hlwmXDn47EEkeCblABF4ogfehlOehLI
N3iPxypkBT/BbSq+qSFh4PHF7ANuBog0OYnjxNwOjaktPiTD29DLdzGjzmFy
KVqAZt3WGONMrKzvSDe/OaxhfEXdvYYVY/FsIdxXXAzsdZrM0RqDzo027MaU
n0jIlJsEKvr3wwcOtRR0JhhBjGP/nePCjb/4dh7ojKIIsmnX4Rnko2XD/otw
xOJcNeuSTG/Wj0wuTUqYeJy55pYD380gc6mNdgq5rVQ+ESSuJik+hW/ce/go
kHlgEhrcoWgDXNXkLJcuoNYtyAtvGRykHV443BzCn7WXTpOll8MA9KH6Njv5
PhgafEUrHwZgIcg09dEz8YJDGF4z+TDqyvjxEyaRd6Js0WgzMunXS5I8EOpS
vA6EskHh9K1hG8y3sJ40XogIwmGAbuJBISsjLpM4A9QoG2X/akYIhI7xs9A/
BFxGa2GOFJ9j5VYJl9MqmXJ/iHaFSWzSkLmLWC16/ps28RbDLnN4vanHIA4A
bM4GCR7SKQmOnvFLt0IlLcBYOaQ1oPmbLRaPjLEyncfXGBK3KEEzrVGFzJo3
De7LlFMwhHjgHd32gFfHXhZZUD60Cy95G7xi9iG/7HmLGq34IiTuckr+g9L8
mEIGeTOa8QYZFaWUVCpMRihj1Zrgkef0DH4z6nW0NxU+usf+xhqo5vWmN1qY
h50In5edUg7B7yCdHW96oBAHKLyGJIF5gEC5clCRSaGknRC6yRggD5EDIptQ
EH0AmWcS4IsqCOftlgyzuFECkJnwCzGxeuK6fTAmP9qq8HzjQX7FfN9KNCCW
CicdYE1MfeSqk0Ks26aUsoRXwzHlG9Z7erkCZBFq/8VVZSeSTQU7n+awWFO/
36pbxT9CJgo6hx4n46CgnGyF5UaX2Bwt2QyhVwmf1daGcOLoJwItKNfpctgF
ZX355OYKu7B/z0tbHTLPYG7S95naH7A1UAvwSP4HJPZEoX7HchmzP2Ekwgxf
a901xzBhqf9okQFhcSmSD87Aq89qYJ4l47oblUzBXk4U1JT5rY5myCC0oyAj
NyUDSXZC6z4bsnrBI1zxlqgq3v7462U9BQxJOvuSWZfbB8hyuP8eyISqa41y
jkcag7OL8GlNkBtrzunNNqSTkGiIEMoQfSfgKJqLEVdcZ+dP4JnWJumNFIdT
qA+eouhU6I7Y5g+JwWwYayJ8IDAzGAcn7Wbkg36905e2dmbZP7q4avU1gszZ
AVwwSNLL3nDh9aMQpmBuRuykDZiP+L/v+Gj5H4ytACdKr7p8WL8YGasGEuk1
dr2SZ8tH3aw6o/yQX+v1sMbkH8cYkgEAO1/bUQu6yeZ9kGgFCIfCxNX2JFFE
y2EirTWL8023ZPeO1cozVxn261NdqGQMuNd0uZpm+zAXCe4peYU48nq6wRO+
EKvEs3fuyuRw3YHPJLGfmrw0ETY6Wg37ZqE4hDQcpKXTCrXCKyTi92njrQgR
nP6OZP5GNHbHvmHNYSdlWxlqGKppSCd/YCVjmfvyZyydqhaw6uY/Q6V5EiAd
TXCzGlILWIgAlaa+K79Wjyp4iStwtCLCkiufKTVAwgIVweR1hUo23RGaK4L6
pn3FldCenNcRmZ3iSSyuV2d6ZqAZZYz/cb+nSGHsOkaFTZjKtyNiQvocHPj3
FjtJVnk9tQa/X7mhY05SgHMesZoAdXRUzNNilKtUv1cJKSWvJoze0OATW62K
S5Ew39TLhbjxZJ4DBP/gj/jAYQi9FA6dyz0UB4+gSlwZtgvyRJh9+rhrBD1B
G5FCPyxGAl6em5FLsJs3Lhwet09HoM0pdvJ8efyfApPvi6ai8BwVfmIC1Whf
zNxRF/6hcHOrTS7kd/CcqZT8+AMhsjY7V2zfTZvUw6D5XDLV6RNRfg7ViFf1
Tu+yaOoQEMn6D3ZYU2AkcStTatqwl6NkXXKNGlIoArPmXJiOUEYKXjHhWdef
po3vTdDTqHJODADAkDJGv1NrnnyQtiXS+tHl4vTuP8fbezzA7ZBHGuDNAlKW
QNGsdouP8Ce7JVQ/9pyvb43FcswrpKAli4W84pu2PwvTsfjys3vFacoK6FUS
+rcmc/45FW1eglloVwzMJDfBsjN0KHFyMRZg6SL37kAJQ04kaDLY3P3E8s5A
DwmCriei7RVoMYxUPLj0ZLsNGO2WshC+99R8/PYnqcD2S+fTJ3iae7zUPk/5
rL1T9UMt8bjOE2/fTaVRjc3uuMUCIK5ya9qIMFYrgfzihimEfO8OaSXFhhUK
DQfZ2Cq5W/P/626dx3fPdaN3GcRwNEmY7mPHFfILfV8ZpyXuNgjb4Usl3N0Y
HiKLQgsdFNjF5ShDQZciWKIBIX21G3lt7FfFX0p6eJCJ/NoZ+QkGpJmiqcZo
O0MEtXIlgsEZ2Eal8fq3HB1A0XhjiNgIQU+R4Yu3T43aBpLlo4TkuwGAiQyf
8zClW7uTW2iC770GYOQB92f5XA9tyUIiGV6fip2FxKx1GvlgZGfEC3DQ6F/n
x/9roLuYgzG5s7SlOS4XEmAi3tUcsGIcN+QC5p8CtaMuHG/Kao9Jl18wfcgq
3l5f+lGeNZ8+UOcC6ttSMPzRtcFzeMgUAGuSBNYH+be9kMN56xSTfqz59qXM
4256TbZcOD7fX7BjTlDa0LR9kyO5fPfyQ8yE4WAj/WM1e86rspYm4/0GkQqU
RV1KypvGwmPKLH5VAaEcqtGxezTU4G0dOCvwRY4o2nDelUOqlQ63q9QKK9eS
THuDXCz0hvaQ4mnmiXRNYjgy6bR4vMNgPmd1dzXwV2B82XjYvOdl9NCj25HS
JaIHpmAKcIjviPadntBaCP3kYoW03B1Dgf5iWrT33VJMBXGIJAa8EaXYhClP
wX2NReW2uikzl8JsMGVeG3ntZtnUEVD5IRaBVWIShqrupuxTFuT0n9aO0Z33
3MpCcaEEAVLx8PunKOmRaRPPwOC2H9GhZ2L8QHqooFtoJb10zqaTW7AFm7y7
+eVMqSQ43nzTkJLZfRt52CeYoAF4hVQoAGDDnT4DXIXD8/u/GgleAw8ndDOe
FyYf9qSH5zlKffN4KhB1/Wl22lktHSfXxRbXHF2+jc/PL2D4CF+9HUN6P7Ys
BpVQlUvA2PL+3Q5fnMAjHovYPqR6a52BXBTcPXJekG9sknN4zmHdm+1bZWcA
0KYQZhEUkrKz1xH8AEcoFjwTYTg6tlorGMDUVJ4/l+BiK/zjVuS/BxARbN1w
t250jcjlf/i4kIcXSFl9+lU/m0IMSwf08dGQVrnLehOJvPRuZoOFV6yUMGUE
cOqRQiLGIWZxQiEy9wLhExz59XjQVTwqojy14wFREODIo1i6jKCJ/8FDfGuc
yxFG9f4UmhvQ1INTux13T+rp/hDYaw+8p48iA3adQZa017172T+213pOoIc6
/lnQ7d1tenjgi9hQg5NfOuBR1MrRYysFB7GfDJbQLs5/Z2akAECc37CzNZVz
2sv7/95rTSe7fGnvs1vCf0iC340XMfF9TbwMra9HimVxV5NFIumE/3j7EbRW
zSKZE403IOmaPGCc28pxMcKY0VTtgPcscHI/VHMUGvwuU80YqFX/s35iFQXi
uBuuA7L8ErtyTjkOgAVoHHsmLg8m0rojT9C6cxpbR4rI0luuYrdMVSGMMQ1o
KjKI95p9/c3A4nwEQDJOHnbyrlYfIt4XGq+cRhysVg4tWBW81cw9J4x0u72x
xHOk1Xo4Z578hdbrqw31m2VBFdKlXvwp2ke8RS5gnAFqPi3ZepgJ6QarNDVq
ikgJxa1/zYaHFVfHlQH42jTglbwfKIlis3WraO+eMVZUKbwjFrw0i5TJY12X
fNGGmOBGSPnF5qd+fJQFVZZtZeFonAEN2fMDFqtPxPQs83IqLhr0e/HZ3p0v
mpnAHRNJOK/q2862iDj54yiRsD7ON3dsGmBmjNg4chqMkRRpDuXuwBjqttp9
hOIY34APFaefsDC0aJMJMcPN5HtjDNs6RyoSmlNx7im8fiUlGqrSM3k/Q7iU
WH3w0iOtRkf/zvBVz3sBP/4ma7d8b/7noNpHI+XunHfF8sbyHl44bDHL63x2
hKoF7Lsndy62V9oTy16ifb+Fmg6Y6YkoRT/IQ45MQgu5FquZHNMSxC3cWtuw
c7g4yuYsw/pa6Iu251QUmCGlRG/Hfpt0ZdJpFKcj9Ro/aGWToOyJTojKhlo2
crpE8l5ygGzIFbVhKzApXbClmiqo4pY5zMSbqFqbosG+T/VCNDhHQbnfmOmI
W5x6qXfYpp9lqtMVJLIzNd67akC+KT/+cfBUUdNs3ca1bffBadCoSGReN9Ft
aSBNeErsOC/jU/nwpLfgPNl3ePiXcyA6EeSCBE6ZZxysVjz0HLDhYI4jSSr3
7eCCfflVEp+L8NeEPxQzXaBCVOsm4r2RVvg8XZ4t1UpMRAvV1frSP3rMg50/
eRqlEVu8V10r6gaybCqgdsjUrl5H5a+2v0yFlZdZ5dC2Qee6cyRSN3lqWtkn
+iBpNJgpDXPmQkX08EyxnJbjG6+X7M+YLWCe6RO3PCAoUX0UXE3nf85/kuVd
vYAcIJrFLkSApEU/UF0nAwmdrHGvB8TOnf85f/122MytYrfkC5n2FwXhEPBL
Z48ngdVF70uWzH1y2Hiyi3bjP2bV/Z5fdk/rVNAzEdsPEvErG5UaNJGq+Vpv
snn2mmH8yMDTtEd/3wp0SG6pfzRZU8nGAkZ4DKnjDD1aBHfUsgI5CaiNNA+H
llOIZp6JSViB+7yJNT9gzEUPivdNWlL93tbmkf8EKsynRiSAy7qWKVTq4QPl
3Ic4PwubYxGvev69KSfMGauDlb4zshDRxjYhtLNhkKk0piF+EUUvReabCcRt
4NsMhsB6+xAN9jlTFkZENnzzfe3WzOxn2du9/MXEvEmB3gFXRbu45A9sdtqf
FwwOm1/nksqM8RPX5mgdTQ6sASbzW7auL0MXl16B58HoXnhIUIrZKuAqUGBv
Z1UZ0oLLfvHvvmOuUha9UGBoKU+dsigsazuJe8PS/z0wwbyZZYbnHQVMo4sZ
PxENc6V/j6PGOsQq5t4hLESiyfEGWp4QqjaQlwywvXQylCTNIq4qlo5RQtBU
NKD2TJqJe27Dx8omS6J9QhYEA8aPlPqg4xfoqo3toiJa/9sEmMLES11QgqEq
g3hBROpLQQjquqtFFY98MSGR08BkfDr4tGvUcljF2QxSgTx/L/H/NxG7r3Y4
CbUMVI6ei0wJ4l5hKIX+HD7vejmtluyOcJSLgyPCqhcht/EgfN8kkUSPHbp/
IOgnYTqEgs61vtGjH/rpjicC3leUYmThtITiqhtoavUQHXLG3eQwO3B2CFom
8E/+ED8AkmEfJq5HFcK3SfjtAKAVRfIqqbvbgozHtovyupS75BHJJgHD5iSP
T/yfFY8cYWlSCP31QNCAganNg2wfQMhuSkhncxWkWpJN36Sutt9LeNumr9XR
3wDDFtC4oOAxBLBbKvAIZ2nVj9nTX7tw6OtZHwVQlJwTNM2fU/DCjxsxEyxz
Zl2p0zh2qA0A+T4AhpYwXP3KKgB/Fy8hna//eWV2hCNF27R01ByzEFCUpoCJ
gBFRJ5R5JzVvivJKZdq0CbmY+kIydjtYKySg4I9Ux4HHsjuF/WtpABIL88+h
2r22F0nn+jTY9SRS9OhoV1zk4EapCfSFz9jWpJcQuu0S7l2vR4anlW7dtuK0
Z2s2SefxRTbDWjD4GwGbmlJl0QNuQD+kh5a7kbYWBPjonv7Nc3uOr38NdaW1
stk06z9iRZufXnPvsJhwK09mNMBZ0sqNaHsSIBDyxmhkTXIEYEVEAGp9/nKi
pVQ+Lkik4OGKYKTDXqCcQxIMmdziDhWZEeuGYFQyXJid/OhHMBq7Tr7sjxmQ
yy1iiGQNR8O92uuGLv1RmaPPvuC07EsfPvIpGLNKuWPumBus4UE4pcIi/RzM
S+K3o28+peJT77ncnJH7gE5Tjkcw/NZ8AdpZaUmUz4paLEBo4FCI1HOcB/DE
gp81yZEfTK0XpvBFizx7ihk2DHiaVzSGqUgHRnFm67wMuC6/OU2GvUSBl497
04ElzzsnT86qKs5dn9Se5zIdbXYe/eQHYwbmAPFV8glHA9jk3kY86kEy4leG
RpwW9ph00OPon1T4/YzkTYANA5kTb2zutM3Ac+xB8r9hZiV6/jm4jcYsoq13
S1lDYm30AMdgNoZwuJQxyU3ZYzFJiYJEBYI52gfc2A75u5Yr2e6VIKlK2Jdn
Q3U1+w+hzpLpTpFJRURSjWf+Qo4SwEPNcCuvOwgixuBU1mx1KBnmFQz/N+sk
oixqruhTks+KXnXDeoWQu+46GoeV3zdMawGBCq33h2JIt/nXlsrtiU3lpqWP
pI9tbUZOrZqT26Ki9xUmVlev8ledIL/Mjyz0vJHxekAMsZU2+5N86wz1tvBn
vucKr/HFMnao6CcSBRfLcb3Ty3DkVGTbUobf7rx0N6vOjpo++hzkweKOytza
z6hyfii7kRb/jLMIu/b5TK/xGr7ho8m6DwesBkQ9fiXw9dWYkm9r2X9ebJi7
3Tub78p2qomThMY5+PFvoddsdXmABsVZ23NQItevlJziO4h74d2bK+ebhmut
nwmz62WqUYq1Ch3iPQebsw9EPV04XRF6iSOACDfHdPhfWh8ui3rcrLKIN0Fe
URAy5gsfCCqQYC8KpuJPrvE26Q2PFtopVH6W1XQzHgTDQS6vr3LM/ZEK7AvP
rcFg7umNBVsJd0CvWxERPLZ3QFC396zvUMs+T/pX0GWqvS0SxBlFkHwXm3mQ
wCEt6sgmI9h9CiNg9XaJbEmI13UYDQjLGpqUr9YgcwGu9Xj4qRKxCHzd0IZZ
0Yxrj07rR3EGFsPgdGsyJTKmcZZr+UCWaRkywylsw9gsiRFktPB/bO6k37BM
o3r18e7AcINhUguzQKnz8YdRH99f1hl+tqjnG2U5HfSMluYGHxeQFlupUN8q
w3t4cw/3Sr/6/10t4N0RcVVKv5M9RQ1wNTZ3ANbJeB1ZbBCjNlJbquqk3TYI
SPpzZFc23PpTnhIyRCrLANw1f2mrlTM91v3e1yBcLkqycTeNSzcYAS3o1Dsg
tetnh91fMEAxm5AAP0/KjAnObPfti7M/wZ9ai/wGjWq3F2tEClesIyi/SN5N
4VKViA4Uow8wYUEkajcjrLGpRpI7cwzSxx8B0FIsmfjDQCxI0VHT5v4MjrqA
CwTvvsDXMzlfpSlpKtbmltejYJ3AbLcMRK4qHFqMhEoGEFS+5on23bEaCy+V
9gOiJ4xuzXvU1hBJosUkz33PAXLU5YfA6cP9EcWLSbWzUSG4zSpzDx8h2Qoz
z49xPNAMTjZmZzlQ/0orKdTKxNUVYZPVDn3HHZlZxybhzyE4olWkO/nq3VEe
cT06dMJ2kF4WOJdTF4m0UcpGQI2Jj6lC4wAy34TMTgQoOCN8/G3FIaGEmx68
cBATL/3Nq3OKjYjq8/E1d+0oeRbaMtsA39vtpVV7QT9pxO0y4Js9nMlLGlsj
6qIVH8cRo89aqwTvThYKgoQ/NI94JuiAKSO5NGjz+h+0sNuV77tv8zJlzs9L
SIpp1JuulCBNHx+gYO9XCOHr45CaLwMNSMubXxUel8lYL1PnV2fObZnGSL4k
KRMi3YIAl5nVmF2dxhMmeBY7ET+htS52c4yiEXWI8N35ErjnBsgWuJrec3UN
uNxHUo3iy/9UayujiOLaZQI/5oJ2xrOwHUaJjgfcyDJyuze7dVTCf0Ny3dJ6
MHqRF01DcMglsNlhP8NBZXx2EKh+QtmukenZTbE/SsLs7JHcO4HBkAzM6iVe
LIbkqqvD36TJlISj9X6N9hgNRVMwQptKmvJ2Wvuy6vKJHA+wg8sgK/PAG3Uf
cZfHxELP+6bbwRc2K9gN1WLP13hBQOuopkDj4yoKRKbESDev8b/RoP9PwTQC
d32j2DNq66VSOMPLLL+e6gFYbhkgmx9ztMJhIsh16bMTVJxrO/m4vuBgA72k
A20bZmXuXB7q9O3MnxtfuZNLSVMeONb3N1JZwGBpG30WB0GINRvPTRSoZU7x
hzvkPe302OUu7eS8mEhM+ln3BOSB9dzONG1tpzbHF0qBtI4IHpG6PhkT95Tm
WI+17Otg32Kjp56rpcRiwHB/+TbBid3jjkE6O24lTIsCyQpTwX4nMohwMBGb
p9yoNvYAXgN3catP2c/RWUanxSILjigGH6h2G9YPP9MblywSCvYyRxFwYRU2
Hn0y2YLy3QBoutPMl8FTi4EbCj9/6gbe6XXr7PsVkEuv0sP36oOukOX5W2j2
riAy3Kk/Ml37rnQw4qEFs/jNKWB8hD6BdDYw5RUCR8czgTTlN+vg7G/1i01o
nBl/MtsH9x0BZcdXZmPO7GzBExP897h8HXret5CtrJHtyah/v2VjgdVuZH2S
jUP5CDZMSJ+MWzYAGkx/wu7GXuOgO5YFyckWy3GMRlefWMBZvTfb7sKOymu5
1EbdmA+vZVV47KiHlwUabA1Z9COP1rAs4Ish0UQKcpUwv5PEkVmpKkdifQs7
upU8e5ZPWYudVuSjszLaqxZJnzY14ZpHaEMfMc3NIIE+CZHAEyVZ8C//0T6K
3OkDcRMzCLjM0eM++/gLX3SCcexWlrh2iiMG/htoFz6m9YimxflMqGUbw+1F
caefiG2Ma2fMj/H+QKNizswH5ADtw/94A+z+I19lQ4tY0O7U9Zo4KpRdGut5
NmxAC/eV+1vCXs1D+VTgEIoqfZHa9b2YymuHGSjuJDVKOG2OVZ6Ms1f9Iv7W
gvQxKUzjugGsbsolK9MYRkhxEnhyFql8bRHp8Sj4D/kaznncSjwEIzWC7001
WtY6/3a11cBY9fpucB6MC6HHsOY/vnD/O27cMWLZtvq+hu6G4iuB5ql3FlII
nWRj5+y4slEtU/BtsYMxN97xwgq2nFH8TQgZMpJOmupA0rZ3ChukIUYiYUKH
afYbcjK30OOiR2Ec/R30x37Ejtd447qv5rW6DaJsKQ5vtZrrc5rgyCASlJ4N
uFCwOKWgQZqjfO6isDsOuzG6Z+TEto5Pfp25uzsk9OJ8Zeh7HoCUe8HLIr7i
acrWHDS94dKUrr8z37ZB1Q68C+Ac6arfDPLpjkUUKnoL4lXw0pK+GSJR2O7o
gtuqf52OyNr70bfgH8tm4JnH/unJev+rgyAT4PRd29lQz2oQ2QG9YdUIyFW0
VLmUFXhcFc4Fc0JGkZZpudkP05EzTrep4pXFM85sCUJ1gnTQwnypSkXpZsdZ
VgdLBHotW+et4MY2Dw8uvbI5vfYTBLeyiH5e6xLUJp7l3i6/z35wNmoc+UEh
62oOOaq9kNOEI+K+SV2tAf+viIPIg2c8TC0FE4hs28N4+WvGteYKNvqMIstW
ztdxC6tyhQ0eS7ZahIq4KIfDNI5bnFM1e7FTDOkKotTVK+WY1STsKzyF+cZl
xUwbPx+OEaOH+ol3GAXq8wy698CIfHBS+GdIZUWjoUccr5HZQM5ssA6CGD1j
/9Hor74tQEHfm0Rp256OK3e/w6fA0CMHIjLutkLsKt627IVi3OR45gri1N8N
7scBFMvLgVZiNfTNrNghoB7X76Kn4qeVRl3reAGzCz1VWI7h1eMzdMGCA+eP
CdLv+r46UQPHtGugtete6ueResrrKDyftM+4PTtps0DNRLCUysv7Li3HH9zD
b6eXG5Br3t8ierCccSEK//ppiEzkCVOsskSdxqLnqKqCdEq0TFJXalohsy8U
TFbm4pHrn19lSfmsKEcLcwXifn0NBSJtVAr14jTVlmteMmT0z+MNcXEiF4kQ
vvhntBWvXgK5P/KaQVkkhDEY86CO37LTcSzpm3K2aclMUkRIj1tAQPraxNR3
XsbxtO6bQV27hMkFnmGirizRtrsqBEbe/Kgq4O3ilBW/+2Wyss2x/vdeEDIX
XEqd9cV288UgbpkXS1Du4rW9NBkexDTg6l4ju1DxPVywnG9ejL2mxaNCWXJc
BiAZMKokuzHiHDc9WhPBF+QM41s2AjuS76rw7rVS0ArE11K3xM6AbWTEzNcy
DXXPFd1NYOZyy5lnyRDN8Mv4IZ4K2ls6YTe2III/tS69rStP5Bd5jynL3TvF
8ViwgJH3Q+AGGY2S+j+ZQ38kipK1UxEQnHaVv3i5h0fPPdv2zVRkGdboXq2o
B4KNFUmgsuwsWpCZv3ND2gkxmDhYXgqsfxAPmxrKp5qK0wQLxc1kE0PIzKRm
AdNzygjON+s1ymlETi6qClO7+ecL8ptKinaRdhJc9miuNXpts0HqCh3lWQ/g
AOZoeXfU8V4dHdgphQu6lXAUpoZ1TEtP05ElJ4Q6OKDAEEbhU6rhoCRnldcj
UubWY7BbqT09S9B3oAc51yTdJWiE97BQefe2xDM/8Skk8gpR0l8U8RufyKEF
lpHjrxdzDEyqYlNCZVnyVsFXd/XNcgdOHPWzj184GklFHOiH215FVevd3wbf
s+7LicQKxlAYOfkbg20zumsQSsrJGHlVdZQF8mlgu+/oykg14MuCQh+QPQsN
0CpYI/IN6Gm0gq443yMDHssZcCqYt+SXIl8UaPwWt+ZwTFDlOJZtkI2UaYL9
S+4+u6mJlKOhuOjswsi7T0sPSH5wd/s9o1XDjPhZbs/AM5s1kqNeKFKkhx3I
RiQ1ux2PS3uAiKzLagqwzRFLwFShYUniJLw0bTzXhtYgPqhv1riJ/8nbSkmv
zf4YLBd0uqE+AvIRB+D+WV/fSfUcWJGMaq7pv+Zi1kjTsGXafQaZJhOknI+d
UkXvjJ7nSdcp3LDd6VRO0k3JGTTIigi1ofiihm6cyy2Thkc6yAEnKB/uslmt
IPGP+ssoIiBztAXgv5StBu5slzBiQudmiY8C+jTiXyA8nIsv0B8Q0/Zs/K+j
Xi569qDbLOfCqw8DKq2jCi1Vy1ZMG1DQA/BwrUSCYAONzaon1d4SlyQu4bl0
31YighgMu0YhcHFhr0J6iET0A7YwBQEYPyahFhYiG1x0xeRl2RfK1knemge7
x5VadSNlUR+8aqBuV7OJp0hHxCdlQQ4U6Ajx4VxDEBGG2nkSNHkaCQ7fRenW
BAM3zWFOedgTmGHvUGglOR0FdLpLK/IP1Jfpnx7Uye/V/DcZrg7mLPxtXWXj
p2xXvCtx+ArMLqMQO1Y37iXvL9kvlZotiE6Er4hQdejSDqOQVFG3Mq5PhF/I
cG0N6H1TSQS4qewX/XUYiOTxySRaOql6NjXraos13dzMph9DkkUP9onwYbhj
VohINWX3kxlhirDx5FhbYQvDhqveN+NCk4FbaFJOsJOXGJIYWD2pSCUpWLkC
vlyHxQpD16gS44YfQXha9YtQaYS2qTylzoVyBfp7470hRen7SdjPHtxc9fF2
kg5Oh4eZKWrhpNvV+5p83eTkcC9j0DnpfGPKja8QShKdw5vLP5bSeNUles9t
E32aaH1NKRPU8CmtIcACGTzmcojtRxYFUHPvRz92bcSldppjyevxX2vbov+e
Q1bzlAjVsLkKXgA9uC1XHIOkgYcHVHyV8tY2uvc2M9ROn5QMIyMlH6hI2rz3
3zQHV7JaqPXQo9BGjphukeIETo+uBUgNtEPvpR7ERlhXBJylWltofxd4LVa6
MpbwHb491CirA8kldszf6MLpHmzfH1QbhmL348UvWVe8jPyb+v5PKRJZDPhm
40djRb5KmRSo3rQmUJznnAz3cE2RQWfylEY+bNeQOj40qJFiW7xxNE4fOryZ
mCloWkRqWbLJ895tYLvHP86GmGvdVkbVnx4DsdrA6ex8YxwCrNN2Z/4btWx4
aQqT3FJk3Al+rNqknCjVrJwZ/XZy2UT2GVsE3s34OkPi2Ytql8wHAjGPkQYx
dLEvSHFpV2iS9+EbDCq2c0vw2Z9qLyWKWWqfJ8qLw2gbETSpZi6XGMRvqjMn
ki3RWOWa8CVVclIpOEY06vazbsryFsFd/X33EGl/zNGLZq4hvPJ48BweWXQM
eMyRY1Hc/4m+x1amIS1rBUIuzikA6XHdHlLPrYfSKACIyoGWzl0bYgHdaEvA
ENWVEFHnDw4UmGcBY9+Y/y5mYoCvdFisPYWb+AzC+PyaDNNzL7sJ0Weo9Ti8
TmsLC2B05Wp7xYQKAbj06hRp0KwFLXisxrTgQkSPXVXZvUfo+WKoDO1OqBOQ
opkZ2cgYYGarzAzxgZDVC+jO4jhZzAgefZ3Mk38FC/+hp9EzW5PHh2GVQn/q
HRsoESlw+FcjXJLZeu0S8hLND43kFsqpdGlCHX+DHaXIlEKBNPk3VDiOpB/W
VEDnlA90Ey0JMSXFRPgGq1GftPq55cq9VqF/Wvn8pYskUQt81W2cMa+tEyIZ
AASNglCy0dAV+tsrrPvd3PouCYuNO5FGl3Q01MGzTM5td2uTWsJiaD9i50qU
XOMtZlFsTjmqsn4hG7oQOneSZpVc2ryoxhluu9ml26Bh+nHinWd8EAIu4D5M
indqABG+5031+MoJivBGvOCFB8WnJusJhtXJVTfG0jplPMynsTVI86Y/7SIO
xDZ2YDCm10i3bZQEo7GjsPZTNXo0kCS2Ouv/XGzFwWBMCb9nkDPNeAkZVLlc
r6OGVMOs+MEI8C2wGHJyAVRYsd6q/yRC+FQ0b387I7XpfcJfvP9SoLv+929d
Bi8Ef2KDoudfOgE/gleY+s1kJ2YVINnwd0ViTL/A5flY+nC0UBN2Nv8CHOXj
KW5gm8s55aapkM0OIJ6z7PhVKWwsf1xWgg9LqI4wkslttNVhErGTpCL59gDm
LS//R4SMcsgk156XHXEl8/8D/dsxXbXjrdeXd8GaENjnI/xGCkoIIUptmRgQ
P85hUGt0Eb3xkozdjpM/cBlrOBqPBRzsFyRhg/7T0Sd4nUl/bldiuCZiuYAH
gA+lhSssvk3zjPqaxpKLZZhtQUAyJ0e7XJ6YqZRQJwPM5oZDDdkom0xjHfVW
JVK1d9kFXOBUly3zeM3B/r5PUZhBhpyrlJxM11YsrIKVMpkEfGClqFR1wmp5
uISkI5RgP2Iip4DzTYD7/PuhRoDr8blKv4KsFxV0f0YT65wOpfaE4R+XAwHy
AWio5+SdUwDXPHlw62qmZ3XznMMPBp2n/IdqzSXuV+eQAUo6DjUC6fX/Ne/n
hqbaQzvsi167uHpsJovRMtheTkelmUO53vPbFfgc/ymd25RABo3XRcBCx4RK
bZxchtC4tovWq7DLAYFY4A3CGTRfa24v0pyUR4uQNZ3PmYr/3ex6c55fghPS
rSeRVM+AK5TQnRcljDPSBoCgb6sTSYZm9N4+azxY+Jqn0pcWBbooK/FvMv/G
Xqz1RfHuPM0WUmUofvYOCVKUwMA5OPyEyQJgqCFG7oB29LcPBaiYKBLNr9/D
WNPVkLa88Bsk2JRMJzxpn0rrzHr7bo6lj9ro61NM1Bbt39cvb6BKPalhrPtZ
o4Rvl7GAbjhJ+ikNC3WAss+TPU1roWJzjqSovQ5vzs7mI9tVqbdbXbmR4dL8
CsBy6Hujwvgql1XPBNQKkqETJjwdjHcvm/v5xVqyDoCfrGokATkiprlqb1jr
Mtxutke84i2PqKqFt/U+Ak1FRK2t3Eoa4hoJrkPo0Zgu4nILbO1uMmBDL30U
icTTjTwNySIgfsLCmZvdHhzFxRZcMPBLO2lXCo2yj+1XR3cI0W6Ct+8g7A0I
YNEvdoE7EMhInY4NrrulWZEz21fuLEy8HyohzQqT/gXbPJy2PpHUcQkSPRIX
n7q2PyqdESAODQN+0StBeITanAkE3C8G9+nIfXYLGy+NgB/LJrBf6RVwlW2z
y82JfXHCar30ArRNN+dc3HlTYnhSLrfJ7omGofUg626xvYYmruVjN144Rbrg
yw8LtrFl5CHqGIqZTUlhNSHErJqo5YFNF+RzsD4doIr2bew3l6/8ZO9JsMuh
HHUSR9LkQj4N7YeI+npk7s0Dhj9oEDQykaqTZYI1X8s0VB8B3dW6GtBJCs6i
djFmF1rXBi6ktvBwgPMB9u3BY1eCQ2QgDEqd3ICug6rtZRdSqi3hdfXWQHOM
BKtRtU0jF8uEsVqIrIk2ucynu0Wi3otOD+k6X1fyf2zAsDsDCtHKNdTRe/A4
qJy6abIOZMkcIyI6SGssYGNIKuEcL/cA0TqEpj3H3QHd5IL6JzIa7CVTTIce
Hlba1S0eAde6q9lCaODpgGiYjm0LhGWl09CdZAwGtZnjJbWSald7WrWpXtPD
0OGvPYqduraQXichaNA4QdusslO3AppDV8lsf/QE4q+yyv7Yu/VO8mW9ir1x
p8W0DDHtXcJooZMkzAtq9VZdxGQWFIA0IpePxMqMNhEHA37XsM+LPReyggs6
liBKwL6am9V2P3SXDUSy8EhawYxlLVlaBC0TrrC+B8bGmp1cmFwPs3ZKVEHZ
nhuKsHzZK3J9cL76qoL2owMOxIgcTHHhNN/95sxDVFYoHoB5xCqIG4aSC6qj
M7EBjY9QQAzeCa3OZk/Pe0U6DJQSb/KT3riaSJzuAgJrHZwjytljedHBAqZU
YRM6fSC5siCr6pD17TbqS8WmOCRsGlegnVBU715xGIQSQdfpBvd5AnkZGVm1
zQPt6Qo7LRyiuP2Hr258RbMswf8RYEmEKoXKG+C+2RuxbWcSOwl9HckqWqR+
LIX2FtGAZSQDDSKfcf3Y0ddZVZpaIBZ0VNwvwGKkXc60MP+W267FnNyhrIU7
ASfLy66uqhcNN+aLjalk5Y2SXQbB4AnpwD/DFDFur+Lo9lRLU34hNONSe/dt
HV2OEXuQ7DGa+7zK00Ahyv06NUOAr2aAViv57PrlDuVVb/f7KCmDAuLO/V8D
F+iLNBqj75jCBkzYR2+kyvmxXSzT8CR3rKxzUuDM69dbmz6SUFvHLvAwRV8f
SMXqbfOGbhsMKw/QVLMrxTDvEvejiil5bgcdOvfn06+47nr3QlwCaYfZoxwG
JZKNukNjdsTFx8Xnfn5bEUCxYHxNqF8+hnq1JInQ3/ICF0GlYaDDkbHn/Jsw
auAuuZCq0jbOnI1yqUzR9PufnNRxWugTckL5ubu//XYOilVuo+gybW6YM4u7
jWs7bAE+Ct+I8cwToqmuH6k3R3Y/KKtd7q5Dke1ydv6+X4XI+ZYaGYQTyFVg
gFzRxISX3eo/TOn5yQBiv1jbvt5jZV4CDU4CeFhkSde6BzcTxMK3Z9zkrDuU
QFABbhaAe5nMab0cbTPLjESTB9Ko3atMA4sb/R1UU9MGtkZzwM4b+EN/Mzwe
dQys1gi/3H4beUe9SMyw8VStwcBa8yWenMM+BnhEU0w9NI3tR2cSFBXWMUdz
0ivg58Ofp+LFUWBfZBWQ78w3bhfRDhVWJhrFPCtW8VOp0/LglRIoZUDf3RHm
fy1SuUhRAqr60VcyuhPgwDF9tp1JcTb8x3PXo3xtjr67AlCGL+dJ473MsPO0
EC8WqzU7t1wjj+rxnx6Ul2kxDxWe6HZvWQ3US76OxvL/imOlA5ZZ/w9VfbDt
8/UySI0OhqtIpsDgxaqQSnLp5gu41FBgzs/7WNMrOzqONysGeShBjwjyzNH0
Wd16IWxqAoXazt07UTfaQUa6szXv3pIlruI6A+8LHwwuneh3BUz1kB/fl4it
/8hgZxGwZcvkCKe+QVaeGKykZ7J69q9uDNmZZgYI14o/Gxj/GuPX3qwR69yN
QGEWIjrKNiTu30Rit0dajxkoKHutv6aTCzB4DYsTpjlC0BtBRAC9mzuiQ0Zp
5RO9rol1XoIkqNpWegq9lkupfAzOqbyVs8BXx3qnz5UkON+ND/1q3J0TKQhK
kgn0pKcCUWQN5W8h4mkvbUgSvn0Sc3YS8Pr4+1gC4Y4IImslOcOCWCfs8VLP
mIrn5Ik/f9vaqG7s47dVrAoqmRzlC555Mf/2lmz7STAwh/VDG7uIghBtFoZx
ki0K+G2a6mFmowa8Fpkw6kkisXTLgNx700/rUUpZNv9WUqKTbmqmT+ojFcA8
9wcuegCciyHXPdUQaKxe00DfGVlNTeylqAj3IRqvmJOwraDsw0VvOIzn32E7
WQNihnUrYU5tgGb6Nb1bHNHmbHroLKngy8EBZeheapX3gRzgB7Idnp2wpl/r
v6k4nZkYFUgzp/F3BYVxJmPI2//b3VDvYhSkfo/aJiP5FFA9G6A0PlnIIY3W
sQQP+Y70hisAaHpcp1foLeqibIVzgto3UEW9GW9MdeYm5p30zgZOtkba+HVx
giN0UtHtQlv28kDwXnZid/pOAPx725kDn/475opdboJ2mOWkbEQbhAVd1/7H
Tfs+uzdhhbJw5hSv8S3b2Mv5+TBbO4CukJ6oXpCmy1AIkv6ZMPDW4Rx5h+Df
zpRxCRZPFnMCSfrH3kozE3IQACEj5Q4V1t/ogXTo0hMmMSQKmHudOTC4rg2N
j8BLBsukehSpFz0YTIAhfEdos2ooKs9QIqroeCeMbsh0SYpVTM3csWYMMfIa
Xc6qRKrlpfBVP3qxyUseMn1wa7zC4+bj3MHYzeCbSYQnkkU652cigXH+CSIt
GyXy4tt2VUn3s1oei4Vrl50FJjGtFN0Pd5HJeSS3KMhRM3tSQfT6tsHI7Qzb
2HfJgs2CjrCjmruQI2KRSAM13x4xwITJLa5NsO0jK19kPW12NQBi+SiEs/Rh
F5ksEl34DGzZlTIi5f1mOVu3J08X8c6Jrbg7FT4aea5IeyXFQxb5zIWHjwIb
vkSgr0/6UNZcgA07aW2jguNr6cpr1RUXRx2Vm9T+7vO1nDKj2+OTjsGc3hdH
8HQAj/kctIOEHs5C2C+6P/7Mq6qctUaxZS+TKyhKHdU8RG+/ZAwnSO0vQEZH
oB9JkeYRfLK7j7bXcb7iQg02yOno8vvZY9fIerX2RBidaZFQ2qgIb/0hYlCw
Cu0q+w6mWW4SEsVebPdmkX9FZc/rR5R22CVSOLTytGVmT3JgOHLDb7GKokTE
NtfsdrZB3GCsl+qu+psi344dNQ2QR+xy5Sb/jD3ZSA4txlt0gIToj1bq+QDV
WqZbU7fOFuo5iLWDFBrVpbcZ0Iot/9+0ChmW5vxJFS0j3rWwB29m7R4uXuIK
HgA34tZ5J3I9H+ZPBwjS/7TD41f5QnmEwgdIck5PgljP1by6N1CDy00JAcaX
VZQMF+OLfoNK+v8WMtyQ8uZTQ3DYhL+8FhUtvm5/bEsoUZ7nlucZFanKXxyZ
CBHtrW8xN1cKfdmf3pduwAda65ixSMakCYkqSiimkBKDi6D+fFBF+3SifXUz
jeOdUL3ihyjdqh0ZNF+nkYXULk5R1eJW7qoO+w0F8bFMIcfQRq47AsCJWmNT
MX0ZM6bDTlzKMdiibH3Eig+HiMQBcJqPmSRjEnu2dhL1iFStaOTBeOS/h2gI
iMLeunxYTUjPdtTWTx33PsrQHPz+KfWnaXDTqxxLDKf9MoM+kBXJFhJmteat
ah6C7Z1L6itynNNT06CgN2TUgaqHMgZS3OBQK9Yoe0/hLimq6eurgFbiigcD
flZgMAevXVPDzjbUDDETXZ6ab8OjGePyAOs35o4o6nrxeNBma6x3wH8f2TLx
0FWNaeBA9N9BVxcMH9biku+U/LRMHhmdoWkKCaNSG5gEBg2UUMOS0fl9hinx
Vam8xDMsWUxfP9WvqsRy9TpnEMAPBuG9kGXQPUaXVqW4cmhIGJAqX99zOHq8
UVeVZ06iWZvf7NROT4ITl9IHnPFlYCWPzsj2PTOn5wl4MnSTCrZeCssqqAS3
RoV48dOyBeDadq2ClYEWkPC8ku7yEfX46M97mwYiz3WwNWCmVOQ7rvzlj+s5
k2NplYP1zKtI6IrxdXmdp5SvhOP/TkSiuSiV7w/zUKwobJZ2RCGntK23nzKK
nVU8OLa3ZyivUk4uTBeP/nkt/pZdHuCa78VM9OoNmPXTUCKIqBSAuDvjh23w
1bpXwJ8110fSfJfl7dn71n2cBmxwh4O5iy8MldTpt5epQHkuA+v+noXdDn7f
urIR3XN8uuIMoqPNdP/WhC+n6Ouas+RJABZFEcvPVL6TmK3nWiVn5UJNm93r
kwq8CfTGc7gm1Wjgt9HlyU6R9fvWunqy+aDjirpxV+Ur4a/+ee66gYyCVDxF
jOE+2jDvzREMPA0q+7g3k9u06TLi5uxRZOX/4wJoNMMxYbScQiXQlei4E+rP
YqVBLXS5aarpvF8ayD3yAtZ1QkBvBycxoygXFp1RZiS14FN5kucWH/FTXKFH
gcPqtwmOvJ9bqERzJe+cqXelAD+PBjcdboNIMoOMeVAPd1/wUhyrqsAoOZ5g
W5E3tJOzl+kPXDwVmtaD0WEVDqeJ3LhdgyuYhB8sBKc4wSHSAfszAmuqg1ap
mwyRNW5Ccrh6pC757fkowAfhGpiLgfJS6LCmOdlNLTPYeuT1CWJw1/8MoWSA
sMWVZGtkmapWybn3oS3p2AnLDNnEXMnRKZIgNqZDEkccI6te+fSmxLRh5P+L
MSNySoqS8I8hGkupWhM1eCPjR1b+2w8Kvsv1k2XWyobsfu9sVXBoJClTCqTx
qysRCf1d+A8CItAC33+Qy+y88e5lQmZpE25QUcn5ronUD4A3GX/bQ07ZiCcp
AabLSLFzKfv2atQnPvxdxfEk3Esq5oDcDX84iu92lBN6kcJpDZvuDvqdnhbG
l6TpS0KaKMvypETQUuBMLgXIBe+cgEQoGZiLa2I6XUbU6sR7TTGVNLIRC/va
s1aJghOSs7oiZ7JRDex70sEx4s7Tx1mnPm4mJ0xIE5KMbQ8nU7UBuw/kaRvY
j/JEQDac3XXdidJPSegLkpCGWt3bIWVkTwLVpf1dy6YTkpopzMmPbjRAO4+D
q/z25r0Yjenr9y3o4WlzExEeIMh8ZtcLCS6MGO9bhilq88ASVFO7QsFdwxFr
/vkP9SHTA+45ztwfAGyGKoJw87CzKnX+Hy0W7QLascqmUh11tP6ByenHPaQ2
GEQAQOfdJUUfGW92i1B7lcuHI12NB2pWQCZNjWGdf6v2qHCql21Vs7nvesZ8
Og+FQNsqspGPZp/Z+FPYe41UbKjnMOKwCtoZwE0FOUEYv5T8dUieQJJ7Gw9y
GinpQk6gJ5aULuTaIdLIfDFzK4ttTo6CtMze4xQ0SYRm7JsT61NWUO2CoAV0
1GWckKDxq5k4umFLJd6cgzUf62cVd96QwwGAqoj5HgZSI7izwG32PxkD3ENM
+If0X5JQ+8rvAcUKBc13PhiAv9tP/hlPeCofVbq0dCjb7kX8YPrHd6AefZYl
WGfHpnk0jIikt62azeO2wqVdFOohQUiDUHTBCR6rUaPTDhFsfg9A3rk/9BEq
djRmCm3oWfd0yA7+lLYKOdGg7FhScNo9r0j8aXe+4DN4p1m6kyqqhS9ha9I1
ZxwV29BJL2sDOinf2gA0ROVTDDvlWiQkM3WG8QFoDW+rSgn/Cx+hs4iBFUQj
XSWdp5F3DV0gm3tU6ev0TWLyonliPQoQ8QyS0AHh2yZwOMwiS3EeHG87AyQz
vo8v+39Fi9oXz7j8tULfxWqeCt8/TCJKQ4Gu0e5+SQh1uudI1mJQBkkF1+RH
wt8PI+2u134jFXkuqsTlJzdSHzWrt8P5aMBGHSt+a/I5xwo/V8NaPAk63htu
n5dkPB1CE5ea1RzXmuMTRU0oSaNH9SBTyKbNm7lyl6cZ9ItwwtEJ+VBjpBHK
vyFx88hQu5MLbwgMRvv9og5ql9TGkG5kiWm/zl3zKShanxgdKjWcBYiwIdYI
rzXtCOBKd07A/iRkm4lFu4PhhMnKDYnL/xL3hB0Rlb7nybBpw7LwQkh66PP3
OSQubs87SBTLQpYASLScGHO36lFc7EYx1eKkCVKoBgQhRrCvl9SIgXJaBsa/
rj7RLoWRnvnvy2fnuiKk39/kTlCjGrF76WdOe92pVgbM/qiOWnlUBhz0PeQo
Rk1FkxqLriSTj/3eoOrhCh0rQ1ZXDc+9LBKuG4y51t/v6GoSJoaBYhCl1pxw
HnJI8l7sgmMae++TBz8seGI2gEyLNWZcfiuXcD674HU6H34xbI2i9wHvEfWz
jhFEjNL+5ilyd+Kbp4b0sn9vwUvcYwebegDum2A9J4YcSYLJZ3p2AL9jiWxM
WkYe7shR4zBZOY1jRG2XO07alxgfXL8MCiAT4gJHQoyJxYpnzAafj+RH1fAg
67T+lFHPCqVywsmq3z5KHVfhdEEy2hdjMG/0ixZ6Jdf2qWVpvGC3jnR1LulA
9SDQtVT6CoNPJLUNq94iStRc3D/cjiZFMRWPaEs8ii+gCrNFY1acG+PyvAwb
J2bJCqluOICjC6qZh/s5u8too2w8qhCXNboaEWe0HP9wi70XbQUNoxse/MY6
NB3z3McbfK15hVowL1YixPWW5Lp9/ZIB7l2C8UkYSgMdfxbPGTDaXsge3zIK
L/JinIAObEiE5tu2vWvAgFG0v+rObgHAbF69w2p2O8IoGTSp9qGjo23yaVnK
KRpmAhZlzHobsLIZa7dQq8fFsKiHE/3nK2bIrdn8UhjmFBYTdvWSgKE3qdVJ
lqCyK7l9MKgjXM1A+jcNo4fbUUHUdjV2YN0JYKYyu0ISic92lvcNV8T0LoWT
3wdGEpSz+sLZf1bW72Yjm3lLtiiuf87aBa/iPzUcvtp0ugUu5GsLxRKLLtYr
AErFIybauDyWBgFk70/9mjpCrNn6s9sMLqMYsoihc5aQsxqqOsAIZvAtKGz3
TLj7FAAZkKf/DML42YipmphjXHuqZoQWo9zC7Vt9DDgZC6JyBGwXxuTVuiN/
bxVUbYdQOvJPuHSIkupPRUNdwz6kKyDAoNftLBIu/yUKdYQ4aB+Si6akyB0W
EiNJ/zHxcclbaDFRfKAmOza4h7dsovcnccxf+87OgZl18ZQ2jWY01i0SMOl3
D6vtmjDKEMlhDfhyg4NAsQCLRLtpnRaCSGR5sKlb/zSIZnNbNDES7ZZizmzh
m3DImwZ1gqIqvPFLnVI8W4RzN4asXiaAacvMFwhk+wKX5lDQ1H5mACcP17YM
JtMfZ1px1ox/a8xab9YDCf6fJ74UcxzG2+oqBuwv+TEKjUUrqb0OQuHxB487
58XAPAtDhNOAM62zFKNSJclXtyNl5CJB2OYVWRKa8z1hatITxcys7c/RvUiB
xISLU71bYLmVDTheLy2daEt9C8ZtJRxboLeJlH+TbDsaQ2BA5jXKmBPMwgAy
GxTrxzejoltRZxP/WegUUpzhwwipjb3ySRlaBAyubDQTwuU6ptOPVUXxw9mJ
2DrFOxWEcqoQOxcXsLo7kT9hn1WGCz0HnXDyOhbhRDHHifjYgmJiJaPyXeCH
yDZoncQ1EYa332SJ7RMfISVYJrVJbQ3qBDSftLelIFS8BJD3AHyiKzsOUcFb
xxA/u0AigGIO4e2GIUZRoi7kMmG5eTLKMuzB14UAc5dSm0+jYuqHXVU+dsqx
PZ3I9TXz5DdevFPX8oQDIpxbOVBjBLNWTjbulvKrLOhdzknBRgsPZW3jvLm+
HulgAZsWqHpx/k4/TY2ZT4wkRm26ZIoD2nABeAAx2unipICPRPdrLo05Bh8Y
TKJ3tRsSdUbdthuJ9pRXhKScv766bzgdzAKLBeqjRFBhu9EIlJR4SV2eD74p
cEUwqOVxCrEDh59kdHMonzYBpryfJc8goqiikTmzwR7u6KG8UWvQO7cSFZmF
dZqlMTZBAV1A66gkToXHcAl0MwdefhS3PJyrc9ahe2X8tCv5bFBhsC3rWYjv
UI604LPiDGbwiN9fWXiEaVModdH8RHU8cZHH9vcXKN1ygEhhyBp9A9AWNtVG
fSadzoZL1fMUUtz8iyemygiSDNuHgwd7ZsAcUU1JroJGMlhLhV0HZMFEEupP
vErcfxKi7nrKxPlhDEPr17+fCBT0ZXyMVOaeopnNkibYsR8va6XpnBuKOh1E
giHbMzpDyyDpUbYYV4NFA4bVdGnvPaIIVJbnGjr9FMDhsVXHXM3Toni1tZJY
1pOPCeS8kBCZRzFG6ols4PLbJvd8+r7PjEC1VoMdcficdzQjDNhVXus/u6+1
oH0O6LdG8aj5nPiTxKEikMx9NDN4UoxIpYVyCijpH8EDwDxgOETpDpW1/vxx
JM34FLd5EB9IAFFDCMtcCXdWxR5Bk++4Q9ckGcV6dNr4donSHAEdsM+L+h2I
b7NVL+qyMZ5E83am/WVckWXWhtlSWUmkiXvDuAFn/lIHzbC/PukS9LUGy+or
TOMrdZSx+WtME8OHcQYzSoo5sh6n89ScBR+B4H5YWFoODTqSov3LURFQ/FQA
IqPlYdJNzouah2XoeLUybK9x/ob/LNe7f5/YxVLS0WeSOkRriVpV/rAw7cbc
pAEzzrwHlRiDwJy3k93ZtrfKuUCOHVLgyD8wZz389h//FDUiKPi1TcyO3hg/
qRyqJ+OKGuVMkbkZX3hgSdfg/Eecvl3Y5E6XBgJ9iv7uFleRoCtL7NknsdRd
gCZ/BURNi5CDs1KjdsZab9P6k493LcR3x2w8Wnj7ZiMiCxcuVPVkWtTOJu7D
yLmTaPRapMFu2qdAFZ33X7v1Q3ORyOrbU7hw4gaqClLaDb9sAXWSFTo5puaq
T1F4eDTDdJI0nzIc0qcKD1g05zgQyLdgsoolIk0439Yh3KnCT3qUtnDuk+7p
LeOPFgWap+Xw6stYMIxFAPNGafMyXSAyYM6d3cZMOhVKmha/zOmbNaL8GH8p
E3ySHiVMcgaw+oaV7+myoLB1l3k4+zlUh7XV8jzfakpL0043JydhopCcA03E
FOJCo0fkxsBzn1M1/wH48D1h3ajltt8M8ADabl2Prt9ybngCqSckZLJzb6jj
/ZQe7NnNmlFYgMXLcHgzAeKEtmYMDgGSfbufgtaidDMMH9EJjROS/Lqi/HVA
R9pWP7YeDYl7yCfUW+jcI+JaKmP4/hOMkUQiGMpjiyZXHcjjCC3BFB7UxP2I
VvhqL0orZwyNmIaur1bZMFAvxYgXphtqYTpb16jR8J9RcNub4Pgsq/7TeKmc
P8vzw2hYEK5UgumCDXE3BngPAakYiBMUgotBtP0D4FHtsjgzMn4HmG6nRlmV
LLNI47nj3xPSiyQtTGFEu5+a22aI0ElSA+cFfVZ4uYjXfQ06cJyFx4ikovch
nlsUvvklchG2otIN6TsDogtfDPNaBxuwEAb/RsEKxcgzWJGMaMllis5WfYe/
AL41Azk31T36nbfCoQrxiYB81ejcwFjtIpcl1pR8pcQQrAktmfwTHxQEk/pG
YFTCzVTS+0v3DK7UnosaH5472mj64PK4sbGxvlqz2eQXdjnB15khoZpQH2+W
/0kZ3Oegt/5V335PztwDSIajOKcS67TISuZvnaw457Vjy7zf7va+mgdx2HXh
YKIo2tB8tMccR9AeNAz5NpKrpLPyt5ceL8xVivCnWnflXESP1d4+ntzEK88y
glcCSo1kjo5R6tyv1sLcDuP1prTgDEoovVqaJpz4kCj2eyasJWmnJ1kbuV5y
oEdNTvDt21Hp2G9ndI/OS5Slf5rpNazhaJ2eSz9bW76I3nrzaparInAsdI/h
rZdD+Xu2HIvuxmfgrW1Y2gverbrPdOV3/Ud4sx3WqCvCkHqBdCSavOktHePs
dmmhGqSh/ylibp4cWFEPpsmJTJRsfWsST7eEHX/lYUR8LRQ7z+lVANa0V2MN
TPRR0oLZGRR1+Fi50xWVZuLvQ80s8QbAhCaX5PrYxYOcOHZglXtLHxufZWYV
vRXCgKPBtsEDCGUkloVV5idZMHYIMJWtYH9BuY2bnMKxAXr2iQPBxBh628yP
e4u/UR59NMtIjaV8k29Qid/LDnQRDknQbP+8vvXFS225oTVrxUmfAivSkMXy
O2oe0Q4nHY3MiWE+jU7PmLHwqJ7T4TYivKT8XXK8goWqVtxn7U9PIcVHoJi1
SssGW8WHUi2tOIltR0lHrePeduohzte6DWspSe4dsupo9gKftK1cciCD6law
Ve4VH2SDEFLMt736A0Nl32Isfhhd7V4/ye8ZXbKdRnQwFDYVRcPpGolzO1xW
wghVgs4D1s9cHfejiWpv+4MKETM9geQCUgewbJVecuKgawgNCwoIGD3HOmiN
Fz2+keDNdyDjgX7fClnkX5n3bRjkJ20iB8Mv/0o6lL4Ekxlb8J77tg9TSfks
S0BjbJwrbXMi0rd7LSAY+xSZdPwa/DoYb/06b/tzqXJxpTZn+4d+RrJQOGsp
G5SjFecIm7E3p+UFv9dH7EoMTlzk342NrSKVYcLJ9rw7QSsPPFMSg9YubA+W
zZCR8Th7A7Na5W6fQDUyMGuU2XD/JTBxVnjS1g6AiBYu7uY8HXb+oFdtMsk/
n8YoEMwnoT+Zy6Bypq7Siihn+HdjIgfmOZ2Aq+tMi3FOa+q5W9OdoSvhon8k
sGdepnh6b26+e2NGx4HLzgn/cJ2+AupT5ihw8qOQ74/vEdP51dESwiN2/Nma
judHd9B+YcYjezSTOWq1QepA6Q6d44L7DrIunv/Qpq3yD2ZnNH4M+wbAEFkl
gCyP95xgrkzTUQdCkx82xqMcy19lsoAbGWSL7tirYNNDXR1p6W34P3m0vAeO
MUfuPiQ7KBY1SLRvDdTX157XhFaIe0VVfiKmvuO9j6I+3dnnYvHeowFxnGul
ohCkcvTzYIwQg1NOxFguyPPWLiY6oVho7rA1s+Wze59L3yiNRvna5G4egiN6
gQ6QUl8kubdJUOdwQCPcf/Iyu/c46FcUFfYSFh6kYIeZSlnrV8ylwBf1GacP
EQuQGXbD8O2pNolr/uEn0awTAOBrkfNOrbp5u/SfzRkakRxe7V7rZce1DVZj
0sWKHXXWcMV2G5jXToxKJSVLNsI/x4OxVMdwkrqAIlMlb9C6qNxmxpR9NqBT
7Os9SSIpqPUWYRDljwLDikefJCtfPRl+Zrph0oCY5TQ1696T/AV9rt4QtP5J
7Tu/zfIESImF/Bf2x0DedJlTl7kfKXhBWz47Ow5d2xwBE1Ha0IHgLn98b41y
1eFoDt6BgiDw+JE7xaD6VykaySz0aM1LaxsRfuzU2LBYIIrTIMwbZhF2xCCr
nDX8kouwo3i1u5KDsHUiEbZllGIkE3TR3FRhTGVLVq6AZs21Uf756zxaK/0D
OFTxB/TyHncROS6g/9FTrnisclpb8tXmYfH51pnPKGWvzcKxHnDn+1iCIsBK
xxL+PtsUlOpW0sLkaViGR/wwP1AzuGZU61jZGPsARV+DyXUCLk61n+IzJKLY
JrpUaBta0BbllBa7oPut8XOOyUo9pWiGvLMuC4z7DFXa/1Ie42SAx3f/0bRr
Nac2BeH7Ny9y2vRkMIKIQLNDUltGW8x/xY5LsYfnLmXJ3mjAMJyZCbTLOa4E
xpQ4KYRwLQgef95Ddzfn7jY6OfXbTbDtpaxwYh4LsC6YlE/8kKhZZtlxlVme
Lj/gPWRYkW5Art/bmiZwSWt2ANI1QCfIFrfQKuUzNZzwvrTQngowdO0xto1x
I1gXsgvc2lWdDgCrhEvA35jZaQ4j/B1uAkozr828W82wst7pPoX3dxz9avQ7
831kkKJI4ZtlXEPppAgVio/pBOA7QJnZe8pSawyrk6qqJwa+zsZF3FXoM7u2
9pvxjlcNWVrgs5vSMipUp0t0+jbO89+4oArU3bOtA7zgOEMgLO0k+w3qNFbY
HxZ9hHaz6nUcMhM4TzhqMCFz9SsTs4Sd/kCDlPGRIVws96p0hZUCpBVoGuxj
E9OPxPMbaIM1TPid7RqXVaLFuN7+fK1HEKm/Ylfg7MMEdRMnLX5/pnn5OK+b
NQHo1X4eEST8BZb8QQc37U6IN9fCUzFj3tbAnEDReXu+efhxR/L9PvrnaWsM
9I/uBFQjscYVsAI1zxL5sVklTWXrG1mslS510XbwU6/doD+ou+3xiudImpiF
bxZgml6pS5h+B2VuLSmf4ND7ZXQF+Y3s03xuHuUWCcYPoIbxmMdwFzRtqeNT
3RLkR4yVbhupVa8F6g4dTkla0zXScfKHOplkTkhqJZthVOrV5j8Npw1TA6Pb
HMAgnMIUYrEV7ZlzAy4IRYdd8CHompmUiWyHCROfN3JVobgs6Zu7/ELcOe3R
Ie1y+Oxnfk86udK0orWZYUze/BFzawc79/O72+s74qOZ2f80nJWaEtIX1EwS
jf4/jrZU+huePGbCq7DZixjEkpRsqXREOEAGaqSDKn9Jh2NNgvfpYP4vRSpA
ZCqkEgszoi0NkdRy+VTEZ/D8lCm1L4LV/ERmqet8VukJE6somPHIa4avkDX5
JGNMUNYkoditaovTpTj5Ggb1SjiiJdIuwlvom28Oyi0mUhuh2p9/s+tmFWto
hDUSNe+hpFodKxsBDPH2mN56VMfLyoJng4o+xKNVBaUoZPeXrMNr25d9nnAA
UPi7V7QGTCH4wxnky3lduJgcUAtaiNYKB7mrLy//cHVerkALCiZaG5Qs8CVS
A7u3Mnerf69ugkhPglZP1vCwmjBJOWjrT2PhbocoJOH+YnTTkXAabrtkZAKP
zmBCKDrY/jZrL6bGORN6CFoV72P4jEcdD/Md0JspmANMBNVgwC7Wz+i73Qcz
B4Mn30gRIdu1BA7EZVcR1HiFWRn41NiXViJ2OJDzligqFnWnOtqCf4Btv3XY
ZS7SGh7y9YwiimEYwtiXmAFVLWemeVUA693V7Grna9zzI8U8pp/U/ij91p5b
oD4gK4yECK4cy7OibW5JHe1lKH635drF06R2y0H4mgDhWsuqvrrvsTdhhOMw
ktcfVPgXF+JOXBYXcyTgNP67SyXNuw9NsxB1PckZYwbogBAFWNOTNyYarwOB
UpOx6Emu0zYo3np6erdsbCr6I7/mCWnnvr/4hci+47zpGBtXCfr+l4d3+9IU
LsTjxZ+PikL+yjJiZBfwaVoMwvCWxW5TrhO13PFFfHS98DY3kLU+dmMXbwDU
RYaa+3LPCgtoqpQCxDJz4jhWffZjFk7UzbG06MVT/LrsZm+hL26x1SC5C8U9
HFHdluSeCSRrQ077jcSDFRta6/qDF2/Hw//1X3uR50VlAms5TFcjo0roiZMb
I2NIFCk1iG+QK7C4baFrzfC5+vs4e3p3ZSr74Q/UWsoGXDkXYCD3JHU6wAOc
y7XqxE0pS4zmx0uXJyKXFkqZQBOK4dhVm14Ui/65AlzOU6D2HBIQo+mPnCLP
xWmvXW58Xs/pOh63YTFi1OnpE5tt6Mlq0wJvLo2liY1n4M7SKdyMdcOpeXYO
wcIbrAar9ZmNg8yYzG4CfzBIXr0q9Gn5uemKC7+YctTKLRY2AZp9wDLP4iw9
pduI13r8UXOipvQMG/5w2w9v27a+TTHYnjRQjJhkcRXrawbMzC0643rEoZyL
WDck1rAZa36/UkVYnDDI0yzckxNOigGZ9+tQfYPgVGFWEgkl0jrkLshJwk5k
4dO23XZ8OGOEkKPEdsLYUl+Wtx2Z9uRiIJ4b4PgCBk2HmupeRfzYbV3qdaXt
z0lKQKMET2yXDpVEmgA8KsbNkA+T70Jht4cBSlFvwQPOUZQm31upcD9Gk2jb
4lbcon1rauPuCEr12xRR8UnJECS5fTsVOydw1fG4+EkyU6sgQHBBkzz+93gY
wZWtJ+t+EVvKpvioAfV6eYRshnqvihcvZs9DRLKR9EYr9wmORylHQOrSRzNc
Kfuh7+N8WrPzCKaYqZlac6XOw//T0/Dq84hWcEhi0fwHIZ2zNHBugS9qXyeK
qmHZ2+2RJNJAfrQX5N2Ma9e1oXtZuLD130fcPLjz+rd4XA/yBt+lvYc13SD4
/y7GoiddVZ+R1CsE0WAgToRqSKkJQZDlqHw9CH/vrx8htRndqDzd0NojNXKP
CzwyJH64TswP0E0jwSEltKAiGmMDxZz0SyptmZAAp/84CaqjtAbgTKK8gmqe
Eyp9JrxdhW2YHkGIJolwt22s2nynU/UHZLoXr/tKLpCklw6EosX964scfpl+
jzl5xNtLA4LrOlL8KPkke/yS2SsmisMQVRAkK0w93kmVLzrv8SV/EVUS7Vcx
8zMY9DdEoRrvNZQR3QADAiGc6UY7Lqno27x0ZoUsvjnJZDa0y2dZhRU/qSkm
jU1GXZ14vaqfAe3NxFC2W7BSTrStHjWfhwJ/4XPpWDvEQMFtcZ+NuVfXtt6Z
nyX488bfbxL0f6KsxcRaSl1VAICkVRLjbs7gToJFm9u8OCxjVcvRmqIpsnE4
DgGmCdTU2+DRDD/JS2vhyyPMELBi7f9CW9fBtES2Gc9MB0/Uvwo+Ksynb3Tg
WwTSOB4EaqneWcUs91oblGurfxCwC1ExSR1ZwREyKQhOivZYcmlhMCMkX78+
BYDNzr7yBnudVukbT/QfIsYNWvVMDshza7CmrUTUoiGxVPqEIu38jAn92zpT
yFBAt/TFkOrGt+MfzdaaH8omAqAaJSGwc5uo8UPS/61BxkZeTEynUnPNz95g
u3aiLOGEPJwpx9R+Ph+1V8EYojqKpJ51KCyt+3Pho+BRqosyBcJt8pc0mrmQ
ZuTRJBikQNmlctoww7IML8aAOzmaUi3dJg8l7IjI0rnwNqxnpEM+9nQw3B0v
ILPa82UkoYQVzcQFZd5XnFIeRZBTMI184fda/ftqZIOg+vTF42VyeLlkZq5y
rIE3yBszadSEnZoLXW6OGb8H2eB1sKsChQM0bohzgiYIZg1yBpE5H5TrkNVr
f3nXsrE98q6VNVKOR2zPd35KiYchHuZyGVxCnGLNen8NeNRMlZWSNSnJFSb7
IfR3/2Zb1+fIiBU9cRc0tZi0mA8AGbO8TleLPsFAfhn6QJes47lPd3iuLU9h
NnnlnQJhzWnm/kwLMPfDFXwJ2dzRPzq25GzIPcPvtBga1gShLfC+t/EacHAr
Fe34DFB3LKdaF4ozGFtGGSvBZD3pxsa9elNLNMgP7rvIGzcoxCIST/QNydDn
5HdblFgS3efcECWuHjsiBoCceV7Hfr6RWgDBSm4CzxxA4KxnuSpM/gDioDfU
+AWYFk3RvxP3S/Jnu/aXr5ucKcCxqLS5RI4Tj042OeOzKmuatwlXTkPXlqMn
cUa7LipJF6N8O+TbWcHAQQK8lDbcy6PD/4bllXRgxuQLFS1+6TrMQ6HwMlbP
3/sjRjOtAlbHC2k0HZgr8bz//vMulPJ4QLEWxBnTOTJpxrYjAea7tHgqb6U3
ekV2nv85b7UfiRAq7yeqQ0hv+TMGPDKz5uvH8McWdL3+fSUm3mln9slbfjtD
yf8XtMn4P9rT4SyL4c0uXpVCk3qhBeO2y4U6MWIeCAmLLD6GC4CU9rOMgCYu
mQoPLGz/V6WtHzKVmmD00yPnXnOBsnM3rHLhVGBm/zcyuclDtUXFF0WgaXeD
yCzrIFM+owgARy1eyOft/HRqirQhj7JFokDNz91FCfx47wTv1lpIpk6llC+H
t+Tl9stEJ6qhcgWgiv9yxwfsIETVZ2V4DoPImHt2ZTBtCZCiqPI0U0LAeqA5
Wzw7rWV9qmiiPVIB8taOs637XXwcLadD3qrJnyGE3vGAVaSl8DISFegHTzfG
mgYVmEfYP1mCwUducfvcQoivs8uLfe69GM/TFbmR2kMrg2dgo3LIct38Nw/P
x2rgBof4vCYmwhvavS7VJPNjhSiFEqsU446szi0EBwd5a998l9c1uOuBErLN
amcV/VujErHEKZgjWaFFkvsb+2JFEaEJEKNr5mSNQAXsNhLBSWE4AHLTgO+f
0cVcW/rZLbVjF30U6CCNT1MC6hi/OxM9lS6ednpmUzHcTk/O2PZJ1z38zS1+
skdNcg2cI3LU9hkbAvXn5YvOGaq4rM847yW7VEmUesBkcARrNDI+AiUyp6Ok
drIyw5mUHaknmOK2r97Wxip4tIgvfpKTn64mdU9oPlhRn7I0gUH3wyyJ2H7K
w+LrGgN/GNUQwukHVRy4aPV99Ifo0MbOXIBGtZrSwK0gKdbH+8QntQf93g2/
ZPo8yV7PoTML5l8tKsks/La3r8qrC9n1qSXbplWbs9cKDQt2Rgrp5vCFnvB1
xfOdMmszZRrtVWj+QMnoYicJVGiCDHAPSqxkNQD8Xtyd9GYaaJYSnWXevaUV
qaVIMkPKcxRj/wnryb08i7K2bw2V86/NTB4PuueIUSxXIvFhu74XA7uAlRsZ
jcbx/95rFeY2EZrDW/t0s8omq7kD8MAyWl3XszT3rbwJMPsvTojXgth1jCnW
+3rIEQPL4i+NZ9llNyESJc+y2QD8XH8o/WA6Jaf6OBVZYdJi2tH7aYdnV+5f
MXQZZKh7UgF1TXzNDRUPLg2VIFREPBHCubEdh+fto6DWRK1vFlpIgn4NfRUM
lM9NgSWEU469T+iA/dNEU0vonv5/j1r+OciZRU1R31zbTGjRH75wQlIyl0h0
Yok+P6VOQHkh9aPFO8JivYXbYRBgqf+V5IRrGLhIEl6AGvvUPetUuZcFu4Zu
4zolZrkNAl0MqkA3mwadkhRRereWXXhkQtMYQLOtkI3xqRZqKHYMeiw04spT
EV0ZAezJ1lY7RpxHznJcdMAyNfAsExBty//XgrOs0jaPlMij9iacCdXy2z4A
DzGOJQHBzaXxhitvCGpSQo3h1vrgJ+IgvpNkJ7C9tC8bBe44Hmc+ukNERVax
izOPIKFu9hc5xaAobcqbwX5uynzfHb0udAsnXEf1VBYgA9OZ8Et4mLVwGjNb
wQ1ahAD/2HWEUTFWBWxjluBnzeofq2gse5618UAambrzsbIWZ9is73O+SWDp
3naqetmdIGEWxv/OSbSjmp9r7Po6AnfPbgI4Ky0U3leU2r6axStplErGYq1p
UkXF62SM7l5H4JqW6qMZIj6CEzR5XVlWtqNhjCZMJwnkndJBguJY4CIjCBgg
vwGVakD6+L9uD5n1MnvK5j0dgZmrZmvK+l8YGbPHQR+cBNq/yaBOFZ93qSki
awOjd1xa/csTCxfrTHU7A4ziBYbhd7N0IasGnLq00F4wtwtgPaweeyc8FoX9
AjkzT24v0J6Mrdh46ATq8Yh+NS04eJka0mIgeH0P0Swa6zp43zOCVfawhvDP
QVaYfXyrSy5OfVquefgI15KfTtnwazH9GaRNfugbS2DfwIs+H+JfgvC5b2Qk
xq4UyTbJVJH/X+4sskR6r7o3DeaderRQVlwH0CUw7M0690++g8hoIvz6SVrw
HxlaZYL8122OwvwnGU208KZTR3gAEyD0QW3ZpdAl6mhBUPyxgTfiebbWyepN
yENfwhBJoLm8n/HTGa2gAYAchwxRr92MFqw2Xr/nMYgcRVnePtizsMWzmQqP
7fOKtXjrsFTWDj44UE44HFqSh7PhuuPAFAZXrakq8sVcQtkv7TTvBwWQkzcP
cSES/jQNnkZ4kR3ziHK5gdS1tQSm3EfaXNSVFaGelzAazyBKvsFJlYxmQ8Iz
rqS9gTlCZQ/8DCUO0lC3BMe7xomrKX9SVsw+2txIYDQNJfrEgGeepPJCmSlG
MlEuxli5oOHF7dTC07kruW8JrNjwPqI9FCoZWFJflJ1NAj+aWtCnwm36XLE1
srZmnVPzrzQP/G0szS+kFPHsSOLFgRpHa6kMvWAjB1kJSOIUaixYUVfj0GzT
TBfucSHaYqYmDISau4JUBkTtX58XbUFQK6ZXuzmu+f2DX061bW9akYJ7s3xU
W5Y6h2iwlC4enuQop9NEXRcL5N0pVuac5LFHVt8OBh4D7AuNYjSR1blNKRQZ
UsGfTRUmaXk4Iv28jcrN2RtYZZN+O6LzYlSy34KKF/GyGbG+NnN/RaBQIgge
+V8jiqpN5Kp33zSVlzL4NjGYwWo8YKBErglJC6QVsCxQ61e5Jw6kINYSJ7mi
KgUUZGa6SSnQHdwHa194ZlRB7o6XenOH+dy5tOQVC+P2IEFiyVCF4pkKLQAC
WR1GUGNYmGWBs3AkptIQUew58+1kKoCq11AxiQ3kUqP4zBogxRyCw0FVVUPc
G+CDu5b3Kru9pkKfKokaSkvW4XgyOnx1RjQNx00YTFR9ZnXO9Cg40AWT2v6z
tfZRU+5ATcXTB6i6eMUENDeQBrq9hiFmUhjlDDmj7V4q3EVUPFxY3KNleCSE
9z+Fat3RhMCQpZzASEDen3f5wjzchFyZC5PYEHfeIFTIk8GjpkEfBcwaRGgY
Ih/sv4jl9Bk4WDUdEoUkMG2WJYzg4c3Fa6MipgiMf6/g6PIAhEPaSUxtkEBi
D/iNMNEIf6NDKHR/Vy3XD50sUn98myue9/AlqVJXZE9xxUSlTVrF4933ac1t
kCtjOjdXILpXhV7hMAQkhDq524kUvfI6ygLEHscyh2H9ho36+5dCjbdxVUfY
ZZXb1PK3zgRJdJb5U396+00ILOcPYGzZ8k9krAavNOxYk0+ZvnNS3dmKNyGB
g7ZRaJRfw+4EWNZ8VhTjGO8DZsi8eDFjZSym/0s19NlJn0/2v4Bnq5CKMdab
H2a3H76KzmX60NwfiaUqoatqXmX/KL29zMU8iz49aRKqYL8suAuEoXBGX4O5
g1WXL15cwwNsUWh2wrxTxMhbv2OHr2/eO5ehp6zGJTUQXhd3TBjLy4+zRyjB
xOf5EyGwU5/mxRVaScNHSq829Wrp5WLmnBPcd64cwN8+ZGUSH/YV3qERrmam
4kCMJnH6ZpemiWPIQeJdHvchrVN0cqYlvRyzQssNYIpFNddq/0zXRSUMWNLo
hDtOVNbsypuiJoA7aXCh/c5+Sle51LccoyRugM6QKgUmJYjcZAgXhASxK7sw
DSwcojTsB/85gxtoOeKIM/NzANVLULus76qeLFh+Ch3ncc9mcUPRsIC2e/Iz
MLYPibGfxRhChwI3nf+QC6baGsrnceas6oFh4iwCNMs4WBYfo4MI70ON+FNy
MVjersC0OPgBxDXppCsUoIkBf6xtNYvAjp/7OqHvIHqElHKPIlRzpj4HTy8i
LuQ3drEEv9wITsj6+7Tl5BXdikzzL0T0WWkf6hSPjg+jBEmdegUl2sIVwU29
jFk42h5o4QbtQvu+G3cQ4vE49rajmav1I+3dJNrCvC4tVoZbGp8txxMg1h6f
KjtLKTI7n4VcNKLBU2cXDid20YCIN2MuWE+kR/Uz/Uzz1TfOaSNa5yR0bD3n
2bkgQDgVfDnAknZIQ8vtBbXhNjo8dgpOGbGvhI9B4iGwWirsKvIe5kv74lfk
hbNhy4NucFIP1j2A9XGQhmgduKmYlFpkunEx8wnir2gs5FPWzKSrtqrtccoq
LEdRZJjoPwhC+zYav4/NlGzOU5klfslec3Fn5TDwPQzp3MT/UFKnpDNr4DY0
vyZN/PdXXDqbE29XfAW/tFdpPQp+vpeQZk90jpNchFJKrjnuGyFbMfSrtCeu
EwZZODpDKtezcLnEjTDE9bif4vQku/ybM2MWg9IQ5XpRNC/y1zBqVihqlaP6
xVd58mlJspYs5hGafeZO7ZnU3mpY9CyLFultjh3wOADkz5LkP8iMVOx9ofYp
/M/LnM0SbtiqqK8at1J63WRnxMW91T192EuhZG371lzBK7k47kPZiyAwPDgu
suwVR3bEL+hNEZP4nU+yWHUvVtsi4nZ0Fffu+oHbAsiDlEv6J3MsV8jXWdxq
d5nU0MAfQMd0wa67/RifkJ9byFG2qajJHIvxbqJWH0mQ7qdwrI89h6Xmn59g
iJc1fLacXUGJ/T+YleTElrUV3+FDWG/edrkyYvHRmBFxYFqsbYgVtJ+jvahy
N07ig+6cczzLz3H00DuxO9aEDBsgpukhIUqOrio0bXTxzrZEECjLKTGrIdmh
6mIQv4ifBzWYMura0yROM5x2Jc7tXisJGaXyVQXckTbXRFH3v9r4acbJnYIx
ebOovxUJtKp5WQu5JV6d87Xl4utytaW441EwFF9Ip3qMWO1dPhVMbXBIWrr8
qeCDckW9ZfVSVatpk0wpJisQ0rmrpxXqbZ74e4jjy4sqUZV3I+1pvGnp917A
iIM3X5bahUUkK5HlyT+9Vl0qQevqz4tvg0HUDe3TMbP3hJ1SrzpQIWr1lLKX
F9KN8y6IPMINGz0nUIloODlazmg27sFTOi5iPr82QCdgM2x80M3FFHrfoo6P
9BP0zKcENKNiN2ROZhS7Yx80hhi0h6ABv7ZRDI0NoSuV/EIZan9Twfonm7hA
fN5fIXEw9ZcEM3uMVxIdovX/G2SwD+qVO7ne8B88+wf1ZSVKGyASm691uUId
rMLYTXRB4uFqtHp3K0p0bM0BTVBLTXy719p1cnQL+CjK/2WhLez9PeKJrhBs
UAQGAmgMHb9RSmUyrlOScJelGcsWMQYOnbg/xLrDk+oIWP8jJS7c2x8nfIr7
gPDqzW/qTShVQHVlTJSxwyg8k/q8WnJPS0yVhXlD7lGxZOyyD63OMzOSTO4Y
DWyHYNKH8MZDhE8osdmUY6EoajkcCKzY7iOIvJc4PC3v7nFMi/8PJPQJXuh7
W8GsG8SLWG1rRunQ8iHqFjmuLzZb3W45+egVYIGjtHjZQDWxuGBmPg5sNkmG
8sYsbNTUFAhM4MEJ5hio1DCXKziR/5FBYWKncjM+Kv5O72dAafKQY+tsfZpR
OfwHokJMztknE5BbvteHD7PPGtC0+soj4oNTxuALwoY5MG3zq6Gs2gzAuzUB
0RY07PmQkzg3A0mIaHWffmJJBFJh1Vx6KcVAvfAEZYunk/BxPq0tNhcY5TZ2
pvA8XHhXwESJbV/+JZ+3nBBfG2Clu+F8ghmjB7ovI1slPjbx7BCNSznZqWzr
DDuOorRnpZyVkHJnyua8FyWxOqUobMas2dXAW5u4ETYlG5RF3pW6Gh3wR74g
QVtqKM3jXVOJ2G/DFOi2hIpnvqVU5PG5Qov8ALxb/heN1JUlfg3f9jL92f4H
Mg5aWwTFRYd0tRyJ+NXgoR0oRNs9nt+oR4Rr9KxjgYRmaA4rHyjiA0rylnuR
NpOWuINTITa1PlZ6JV0xhV8HpKUO33aZauHC/XIMr57hCKJgDtvRhfyFMw6+
wWMURUcAG3KqqWqOPpEQFZ+9pqF4jQsBmL8iY5gI3F8JnDWna06zPOtBSF9J
781Q0omjOmRi2WYvQJtQVxz93r/iihwkdxwZVKZ2IK9JWvQtCc9iWSICTLFd
uLELMjjwI+bi3KwuquvY9zk8A6C97HauW9p0rJ1FpUPCzB5UnE6H93cvCZgn
wzcmJPvUw1/eDO1p6D0SxumlIjkuKFx+lnpIK32DoMlcwG/XZl/ypozVJOYY
FgQr4TjfCxcczwtqK7g1XfWNKH120Mvpd4crnkFkUSIvW0SluNcvsx/X9Bcu
oE8mgtZznZTr8+6VsrOTQjxqH0LnBwKHMDJR5b+F8XAD7bMfmU+/TsRXxMwf
lyuniL5jd48zH2d0r400PCL49qVjvs/vZNEbKZDWC2zDFoBq9wOKzWSONPOe
kqpTl0tcXDJKtx+zi9Ve8Cy6jJLP6r0WaIwiQz+kHbN0JPt+0jilbH0+AK3P
vkD/EydxR+cusps+jDOj/NEJeJ3LC8o6uHnrM3ynqGCysAQ9vZO1BhHBzghe
tCCN+EXaiOTQpi049NcsYK3z/A+N1xRK8/RsylyiXD705SXPvTUQN1Mx2ouO
9hy2H2Rh/kysZcpmJVlGqdzKtt2s6DqhQmM1htg0Kree/qDWbth+349FTnYJ
CsQp7EVOaDbTCgP/2Zbexb6GpnAOhUUPLNdR4dj3aTB23TApkxeuyBnh84xy
BBarjJWt+n2c9zfxvGgIA22TyWvZ5br6kMxH0KmNqDcrRc+1CnIIRX5EPlc/
CVlu/sH7pXKgcLjxnP6P3djdqil6rqhAXf37648dZd4JqYMT0PsA7KixzJQX
quJHyBhv4Nf4eU54CATVLcyEOz+bcMWMtiIDAqzkhM6vgzcX+be//LlwphsH
nF9H4OBv0/SFAToOWBO1QS29Uz9xdYJ41TRb/pGX7GODzHM7AeYdPXJcbAd2
Em9aKEB5EJgsW1gmeDvrvqkOwe8XXKp6AK0RB7SJMjzlk5dSMR7Z3hIhGs1K
TDBiplNI22TNwUckDGUzQ2nwFv2yDpTDufh/U7kHe1Dvc8EU1olfKZl85SGD
Yn7TzQF395l9Hwa2sT7XNKjbA7GVknaxMoBhVh6Wrgr/XPSrGCphBDyRmxy/
Ueb5JbBUlFAFNuThDC6nBMPwk5CWcayY/V46hkrlJ00X8QSv1GS/aFF4rOi2
Kn0uY7COVu8ZF9FApgj+106C//AAnX2fKQ9/F//K1N59UVTCHCcAJcE7nZoT
la+Vs/KBHVMKpRqhUcnixC22HUUNpbR0ZVVINVudJr+qjFwJ/TIcSxhbK7Wy
u+NqLsEhsznBoEm1v3XOGcPlrhVwamDN884//rReZ+KsSm0fJe9BpjqLykCe
y8cIOldQu785g8zdeisl8m0K1rqD3sclVMmoKrnGPqjfl0k3aD9+wQXe9BK0
8w6OeuJ+IjmTJ3GlczJP2S6ixrVw8zAEwF89iDeLhN2IGr1BiRYwgiOuKPgI
WQ0F6OAKWIsH31SwUZmYKBDnnUt7DW4MdZlR5rxaRcmi+usRQZ+2t3iur1vJ
qF3CmJY4RIbHHhUO/rqeA5CFbLITOoErcQERhz9Z03sMhVUZkhSWGY+tydjX
bihbXSKaou14iIpU/qoiMADKrDULdYR+XffoFyPOMRZNURKM7SnKf8RsoaNb
u4Qy3WoFLd2yZpv6dF/diTWNejEWLKlbkHX36Ce/VtJiUVHXC+tDFe/iXfrf
2kG6RC7ESfw3L4Ezj/G62C03b+sxyhsIbxfPGSgm46ikPVa77rheYWIEyNn9
L5GuGUuYVv6rRNabwaQ5r3JhZ7h9I3MOszUJRBDjtfH9DhUnrX+QTCeL05cc
Tn0Gc/uACtDIrTwqPUL7cPi/AvOoF1OP38J6znp3Vei4gcCrkTwP5v2V3VdX
6BbM2c5VmyT5JhoS7mlUK1Ev3YuPxqYOndJAEnNVnW6Q8qwZ847AHbXB+cyw
Yc1ulxOAk2wWUNlp07ikAIZxlt4fYrm7881NF+OdHwudsMQNTNNrePeFvFV5
ZhGmN8/7VNLt+1bcIxx2wzfNZiqjwqoUWIkwiHJ74ke8QH10Eljdzye3wU3g
0DVlQwa294+TDQEzko0pB1lvo+Wqxu5x8RJJpmdOG8lmIFefDJ8eP2m8RQO7
cx0cK/F+7eZpUmtOIqVyM/bm4w5dfaHsTXjQaSbJzxH415Zg7R9CVdqydkAS
6U3VPLFdGDEAJNvcAjYBSzBEdMGkkTjrb0oTD6uu3ZqJa41FBnfqpavXH2H9
sw+VQxyQ1+rEZ51goCjrjLXljmX4TFO525zTg9xcchbg0nYgNVwat3hCJH1K
vUe25qm1Nz7wPZvWSljRcZXBn66d6Vpqqxos5jDECVIhPe/Nnutwwjpd68z3
4uNaMn2sTSAJ1VBDWet4AAGZr6Hqyor3zg7dxtnBUtv7Of0lQi5ZM3y9Xa1H
/GwTYrAuIjfIw15lUQXUQA20Dwb7PsJfSg9FYOjJiSrV2BLaNhl/fN53hupx
41E8xpeBeiY7RaJie5LJ2YHh7VPhtljqvXlmrAOgIUETudoLU0Ad8R9sTIJD
O0Xc5G67rMXOsYP6r6+RsYpo2XAb68MziWfZxPHI+4ze4hHgJ84aUzdDZsF+
VtpRFK5OYwXSByWy60GOAtD5TbF5m55tOqrEgk5xId+4Z0YUyKQ1TsT/Hyff
pP4ROrghUw8W/N4q2SrF3oi+zrcRpkrgt/pTSNJX+mERVLJbraajw7fSqIoQ
oO/UHFtJczqWK5JpsnXYwiy8aFUIvaSfRl1ID6GChaF6yPRq+ZC5FaLl8DbW
sIRKU/zlPuobH50FWahYaq6j1qDrX+P3wIrm/LD8selpVxplNhkQLE0jhWkB
/1YqkGbbU55gFSqwR7Ho2+PmXdDXZ+4Sc72CWQBcU9BQBKGp5iS+8scQuD3q
dK2g/LDWsgUNbniC1o9v2jcqkHCsOISw9cYTglaLmjX+a7oy9A2XO/XLixRp
sywvn4eXP2MFKdgtFb/boAMSi+ExY9UauE1pqvdT79vqofllvXJRa8tbITRU
WdVqGAJTHlvMAyJKGhVCmLuWXFSwIGsB0fcLWPZFQhQX4Hu2TXhbyDl6JD3E
jsMpsvIvcUCnxM4MFpGM3bQngxNaskBocS2isq0FUjTwcXODEPxQBGcM0sgp
kKEemqedu/yGvp7ALGGqPAkqlo1KFnmvQLVorzRJgr9SW+Ba3UaRdY70llvo
a3dX1o77cLKlinX6RdegYv7gc6mrsMvABWtnPtS8QZiewZ0OR5qiFR7fVpwF
TH1F+F3SzC24+HCswCQHfQM+3SJPeJyg4oztUTnni+qq7/oTYWZ/dthcoFCY
CKT3qLAT7LvShRbr4o6wrfnCYVkSRWG/1AbqVaQJczuyYzNyf3HLR+eqILj3
TBsBbtpTSaRCW8xlG7Ioe4maWxCRf1aN7bxHJeOpirtbKGHv6XpheGu2R2YH
iCI4fEYdy+HRig7P6HIZo4f+NdpAALaMgViiFsyZVz/8Ocwnobi5b/NypRiW
m15aEgU1ntYavtrZgaeyToVPHT2hmJG0236sxGzSbNqc1joqckLTm6oDd3V8
/vtNkmffRL70TkieE7QA6wYhcEzhNckxeH8wavJVZVsQ/HRGK0ocxPkwZsd2
+Dw6xKc2u24246y4ZqtjTuvZCBfLZ+LpYtIjL8MiSgPcddPb3jKEQOj18WWu
9RA3AeFbIQFWG8pF/UxpZbBEXeFHEqPhnUd2MJZJdO1weLB4XLEI7gCvxhg1
IfCiTU3K0B8yBnir6SdQpU4oJ7wRpnaJNDhx0rWQuR5N6J8rYhg2RZsVHpcg
y6ErD8gvbUgnUnzCwvkR8Hy6m4cd4QqYFm7GZrCvNAY1h0kD4Y8RYGZG4365
y6pKRmzBsVimJbM6LgpoZNOyGqEjkxh/WW61agjZilhMb9eX8+hJCZ1iDmBm
Jb0VLpQoyhbkSZYCvfYho6sdieyzMnjBafuSweoMNKDrtv0ktlFnHujlC98+
53W0NkLEfYRuDtGyIIBZiUCPK7DdWsHvny7AN1OqpiFsPWrJ4xB5m+avm1T0
1VlzWs1ysqNw44a6L8445hMdjWxSVruZBYHeVjRGo+2jMBIWKWsVjNokWCxx
/cIet9YDz4v3DtqRo62VpMjY1CQnEm/S9zXM8yZc4IM2vrVVCr5okFzlcL6W
Z9j9ra+urmNpETnyrh39IqjaYqo4S7NlGsLir0OiBTDOVYFAgQ5fBD7ySsl7
ix2/hAf5k6dOaryGd16qO6jrihtKHxQg6hN/U85iRdKHVHNlgw1HJqgghBm4
8p2GVvXHdvp6oLLpwZB7jc3BYrlH8g0szgW67DboDUTpsz0Ka87cMsEU/72d
jjoD99ECpVtI1XWjZcA4yEt8E2nwBolPgMQHFoEZNd6DgKFn2wDUWu9H5JEQ
KM70S06pgJEISzNPr68IpzJtSre3MJw+CA2eKZ0QNABRJCs/BEaEUMZcgHKZ
EjERz33oA97HGVjk2ptVy+YU0/M4A/CpcByaiIONTtfKleF0OC4XM6Or6WHf
mHWRGuN5PygaR4xuq8c1U28UDN5xAIYDEmtnzUVFMCpdKIkgxH7YF8ZPvQZC
QfHADY+4Kyw5msJeU7uENW8OSVi5cdSTcdfbTDhM4Ig9nw20h2rfhs0xew8T
uEdLK4EjIC5nyA9h4GCGDI9jLnU7z14iqpr7QaxoMl/cViP3yiIpS6WF8EVk
byWFoS6WA606RzMNADKsb8/WMUE902utU6aJxGx7Qg+6/Y3sDkpIds7HetyE
eiYOglxIpJt5lIIMSI9bENFGs42xY+6yYTYTE48N4L/bQ5jDsmiF42oEeknC
4zio1vNsd0OfOkUYs+INX4UCf8ZCQZotGyXOsyTGOifCxIOO8QppOHhkrpcM
SQS7zP8zX3AbfZ8ILu1W/mkIEpsebof+zLOB/UQiDdvabNegwRtHXVsuaW4b
jC1UtJTKy+UFGv7B6ZJP9UMmgQyvQy31IdhbEx0fiXZauKB1MZiviqaaLmNv
4FDUZV9DjLdF4yu5sxHH0yKn3oL0bf9zx0eQgfDSh811ZHdqObr9UarDapt3
zcs0xoeWjF22FsZctwkHqtOfG/PdAP+U7iErYhFRSZqcE0CMEzVaavIhVdP1
l+u5xVS1QiIXQG/8n5YRdE6afLb8PE0cp86OIYPhUw0AmIfbx4ruVHNqp87I
Yq9z42JB5n2wvUm3AqTUUyTckMg+e9r88BiPtM36e8s/oX4NbaSf0nyvtmjF
somZz62a6fuM7te3TfUfiOBcwwbkueeSTWpFMhvEy4XJYZyFfZB6OaqZwjYb
DPAkvEugvzhVIrdjf6JiFeE4pa+fKWto/w5xGu+uUBvfqsjgIOdUDysu6ZAL
QormX6llEV26Knc/3PJKWCbmafZgM25tALkh4cVITWNOFsLS78ru2TUpvKUC
p94d/QuMzTRKpTC9Drnxgp4x8LawIFSiD90sMraO3pOMKhLYt3KDj12F6lzI
PqlM4LxM/HUc/LM0HUgcnvySnPTfQ/8qNKRulTG3GKTmtXnaxrZdxd+9DJNc
QOTDA6TaFnYQ33zFNXKCKdA5qygQwm0a0Lo+o6r2PeUAoaoFFuObojQOtyuL
cgFewmMYcKEUvDCuqBkv06Dv/Y21lX++mWa6kTKdQr9IYXg+XIqyO7iBIf3m
igmmqYPNKHCtEQ2kILfXQFARnOBBSzQsolLCt6+KXBURmEKCvFfU24FeGgZv
f6MxcCpRgxuaD+l9f7asA8Rl9w360VTLesH2btgK1YqPuuwiBcVwyJxXGIQx
03CxWpxGqwW6OI97+aS/q6N1qIeLSTGcNt65HWI+UMXV0PKEy0cxBxaMCUmy
0F/995ixs2u2CZ5741EfR1j/LJ8/HGW/wFxOjW6IdaRTS8sdSysMMEMX3tWF
hzG9+wnGTc5ZIlfxhGuuBAKs+oflmi2meHAo8fRdz1QO19ZybPNJXrbVbpP5
9PTUF46n5KmOrVirZptl1HWBqDnc0cbVqhQISTUTjSY9HmoexxrlzUzcAMSK
ievnE89H7r0Oj/DZUPcONUZPpQZ7nVIspbb2BcnPhHPvo5zM7880yMlOc2s7
/UKTM9R/CdB6CMoFFRq2mWPR92wMDudsjuaVk7stpJo2+LlhIOmxWslrNzyH
WbZYQMjjcANjFUuLuCCacLNu+dX7jD/6DFgjjYIjDS6b5SNOIcmNhyR2AB7b
rs5jEjTSghioYVHOd3dKbzG6Fs0BJm8vk7nm0fJJegHe21exMEgASuNAxttU
cyccmlWokvV5DcebhulPSM4MSsOawph0yOPNq7tcmY9uNjuxYsQeam1/vo7Z
KpwucdyB4qp35r1gbZ5nBTRds7Mj88kH0yUAoQtwWp3PVxmvmGkE0pxVpbau
RbHRd7R+6KjDidshVjG19S4U2y5SiIR02ymhymRdkrocMZvScencBOctQwr2
zJUY82rOrTq5lA7Ot2JT+upi+rLruJi0ycgd9NhC5CnP2QQgLnK8drh2nn4T
8IhVhs7MQ5qzMILwPIUW5QrzP9BJtI7IJp7wUFPaPOQ8MXQl77ET7Yt4dItq
FTWxh05ATTzvDoUHPm6jnRTBf3Y3iHismHj+p0c6vNWFGHuL/DbKef3ONYa6
Q9yUBYKinQwfeDTeDVUAmCXmcpc6zc164TOVy8xD6YsibI5D+RJNNLu3GqnW
W6AOyLAh61U1txTdUiUmTBBgwoxYxyWvHm+n9VbapOcbIDibXiV4RoDNllt/
L9gX1kXfnuSRNEHpdP31WC6hGopCgveTHxYMhrgTMogNzNYgZlgJvrSvufwO
DxY7EFfEhWMC9UkPQhgzLcLPp5uYeV3uAJ8hznTWc8okSCUjiF9Qgl10vkY2
VMEWNch3bbPq5frOckwBHmJdyegi/QmwWsyPJN+LaxbO7+eL3MjS4t0uE5mI
ISzM5ujInwEn1tfU0f3QWrFXJMKlup0HzrWL4Qkg7kmSVa6Mk2SM2EnkwWE2
/82qYjPNWxP2v9muhGyyVc1i49gBd7um1Ax25hc0+qbKk9rTeihJFp7BkrW5
/0ZsF5vJ3pSvNR6q2QgaSfjF5tW0YxKtMJSqxHJX5T7PrZhrL+781iLbQrVc
ZFHH4Lg7d4GjYAYOA7ZG4+Mn3VkgyHlYZzall9UiiDWp9kIKT3TD22U9kogJ
wLLMCYQ/dWHxBwt8oSUpEYkIrShDV2d8lXzeyWP5K593g9+cDr5hN9zYjcfd
x485B8jmMciZ7WgsyS6D4R0aonX9ttl1wueC+emg5fGJfC+vuZQvrPyi9/KX
SKt32GONC+KRMICWBD3bOr7tkfLkaePGHz7gKmt7P2f3tHwG+ettxA8u4BJU
k87vPRK+yjkCw2K0+kw5P3t4i4W5VP8wTZHlMEFEuqw9g/T17FVroHW2v1FP
beQj1OOyxBOqtyjygewe7s9wmufyHX8MTRGQqXLlBa8QGdiKUiD0oEAz50bi
s4JJ0Q/bibIVNQnbSZ75coSeOlW77xoqh6qlyzkSbqb6SskL9Nd5wlJ1OOI4
o71f/Je4hYrtsJfclfTh88WxB/TLdAtCF/b1TvIU22NpkQBz6ctmebPAJ8BG
mVobhIDUaDlXfx1KEZ9sUMsf1S3FzwO7A0N/u3BCocKg2F3Tt3l2i+5zp+8R
xRQE0WeDXw+QMJ4wP9W+wOC9mOagW3MHZX7wBUO0twRLpHzU3cd6MrlBnZiv
WS0QUnZT9e21tDSh4XFIyWTEkEsW1RmZ0gExpc3pX/WqGbwmN6K4wMCtXtmd
lVZNaia/exuKN67mfOotuphWq0lvlygax49rCAo1UfHJxYIPll+7dwTbwMn9
S2CqiDaD0Fbu/sOlTu6F05Gyo41zvWuGadlIua7fjQr891wSrl/by47iHsu9
3SQOiFqbcnqi+O4NI9qasPNvMXyZT5o2xXUFwWpEwVL7k52v+1oYlkLjQYLq
5uBUFxhB9WnO3gnDsLrWyfMyKE4f6gfySL+2N1SghIXn9S87X8M+hDp22I2Q
59d7SMwPSaICssEHEns8uRwOnzI/dVqBg40PHFdbH5eXovQNrkxBWlxUxm9U
3YDu5jgOszx42IPsx8mTfhoIHTRWFe8RObeSYbJgjKFaf0z9wqlc2O7laAfL
fdiyiz9CNm3Rt/BEhSf/sL0sKee9zMvMjoCnaUcehNv0OKFWtiaqBTN6eg4n
x5EauMKda3+gfEHOixbN5YyUJrxPEM/nDuzjz6M1VEqftZXqa/QBJVtBvoiF
F7hQVE7bVMH27RZnSzvYYCgy5T45/9sbYLXl5PzvG9upst87JP65G/QtPElN
UG0OGgqMD5lt8oQFgmR1ZlluRoyurfAF4CQ05sWpeVGlkwFAZo2IoZWHNzol
3MXHZhCxBpl9i3tS/vKF5XlsKBj1e/kr4KP98azSqr0kSr5eAyBurOYKzFA9
nYttq7kkZIP6RMjiePiiI52BOrXXhdl7HACEDsdlYYJ1M+8g1wuoGTJQ0MBg
AjKJmOyQyoYgUOKooqH9Kq217XtLD8VA8gg4nhwCFZ+Jz75vZPLWYT4c+Q65
lWBl7bXF8UdZb2GEAFeWcvoNf5rA7D4nTffR7pm2k4sFe0xFv9aIp5ndO1gU
l4Q9rO8yaTW6WyQK8u/NBwuzRMvyOPFo/HC5ESHSpt4zmPnHR02BTVJMlnqT
8FCzPosTb7nS0cmpwne9XLyVbOyTndz1TryP1WwTfW3SLEAMB24Eafy7cTfh
4kKsolmIFIYEBL7+HFvf5TPpMBoTpy+GAwsU5psuqCDi7i3dWaE4hrZs9vmx
HGLjdJaumZuUfgFKjqsRxREiLTWhEWLofwL+d8GjaeBMP5cGLgGJceZwspCy
huHRVXtciXCxEduKn8JNyPapWZHyIMPyyjIwQhxxJGLOfONVMmW6JQqUWaqk
Q36pHQuP3uvJ64YyU7h0wj0we6p+pdLSgH4NpjpCUOng6Wqv+hQXKBnrqG0s
xeg95myggcGH7oAFqHDFvVQ5SRyjB4lMI+2ExFyGAvKkvPeNaNHEQPr6RRET
mIJKF8hyoRmURK0h0bKpGjU0hveywdG3PgPIaCRgNxIOK99sJsuby1oKMkSK
ZozDuqZozFtG9TOsNhmIweynqXzwmnqWphvhGtlsIRa2FPgaunzDMau5ecpr
NpRQsfA30r9sH3jI2AC9tppZlEn8f4QPXbY4kPUoQhZRs+XmM1IUlfsH/MOw
M1q3JEDFklsC4QVk4JnLCKyar/kyV7PeaOeh69j8RR0HcMX967LZGznkXhdm
ztJ7RqZI8b1QiGu0OUBD76+1KPjcaVCvtNKKNjKf97CqP2/7JB6WS06pag4Q
+0fNceRPO67Q2a8PNV5jN2R75dOuTIFHJkLR/v1x2VxwfqzmTTq4lyctJYKi
v1+mbZsBCI16iFnR20a1lX8n44Sb+kiJt/bsdWK+pTTMo96QsjZYyStMN6So
/fJEBnIBrDefUE/HyMKxjktA67n2XG9lenXtqwwfuKRKwCUFwVyKzVDssF+C
Xjo51VM0fq0n01JUwJMirZzBM/o7YxSIBf6O6b7DpUm23BimrWnr84W8ZUS7
2PC4Vw1smsbBAK+uxanXd8lXcmp2gVOpAnsD6uDied82LFYFz0NDx4p1tiTf
vxOLVyQ+Q7D/AXhvcg0FGbY8CoTnnv172xAcYd85p1Q2zxjlD3kWUus2Etjw
m3JVPg238baq1KJfeOpfC3lGDgn/lPxLwuHyPMydrFXjO8mvht2kkk0EvWJV
Q/tMjbwm/wZBRfmUgdN3l4XVa457SRgAnSA7e4XueeQsj8Bvyn0rxd9cp3Ng
60jTealEv1md/CxHUO37Cv+mZppuU8kJXhRdUdvW9iNhW7y6en+g9/bQDlnl
Hv53/mvCyN8kUNboJe0NRDkBEzrqOmv7kOKAt8Ccu6ncJUcNJjF7AD8/ZTYx
rFWeto7sq6Krb1HPQm/sYy0UwxbjcJpu1HxsRuzkfFpLphihLIxx3lKoT4lP
S37kJg77jU5SPXiMV5NefuMY4i4qDW7MOH1Q3wQTSVi8Y0w4PJfZg6rPMHcV
gkiwupbrfyoJqNO2w4xQYEbup3sr0x8QS4s5aGYt4tZxyujkK53xGYdCpein
iLHXBAbAJnq9B2plXn/bwSSI0Ss3Gsj1rpUJa8mbsir8JeRFmo04N11aI14V
iONAsJGA/MbUr+jyfCz0Kl63yrjR8im26dQoJFDKWwmJilc4d8HSaeQ0KhzS
55+beMbNihPCq3nR/ejX05rzfQmOKloJyUZkIoMeTd2fFWtsm7bDB+vDagYl
ZkeNyos6rOMYFKVGQDgMQH/k1HxwE07n0Aw0EzYw0lJOFuF1jgA+uC6R7T6V
hofP7VPFzRGU3gyoa+FOp3fKgq1Z9bt+UF0oIrJl59KIX1LgtJEMZQSZS7YZ
ZOq+bFU3T2Z/vP11hvxuvRE5LE6k3uK6conn6quTSVNL0QCcTUX1flohFuir
LJEGxlqc4lsNRX+iBRIYlh1nPgeY56XDpQ8A2ydix8mHcgSN5dYYzkvfCnAj
vkNobodYBCss5P9o2sPCENyn2QvGkbsLeEhiw8wG5OIy5X6Ja4TXQsUmYyGt
/ouKN/Qf3qtBz4IVO5Q0S0Sf+1gcVvKcdH0DzVYCkZf6ew7bSBRN8lCIuzif
v/6VK7urLnzIekMla/GyI5FEMJZZpn+GQ2xsvjoLLBrB1EbzkjWN4N2BtQYE
n0XY1lYV0UJBkyudH8Mg23lsvPkceZtMYQwEFOCiXvnZ5Nq/QbOHtcLSIpqk
QnnY85rs8kFJT8LPHx0+2Etap7pEylaoVQWROxJHXdyQ8BGEn0KDObS6kgmm
C0/kzfnTdePa/sNdInsAF9lP6dF/iXyhCkLC0ODGHGyLiWW/NK86lNtBEy6C
1L6E3lCeTZthd3WU0usJwklvp1tx5Y8D2vgk3v7jUKtsSmKJhTNKZmsr94Jo
TIZm4vy8r0UVA9uGMLzYEYWBwl7ksGWgU/qU/HnUQjeiER45h6TB5vqnT1l9
p6PjaigKL94lviFfWrNC4OEM2p7QEEbegHMLUYxss0Qht+xJ08ZygBGxyLeQ
3326gxQeTAUMR1DqnagD2hc53HgMxAz+I05tjFGLlKrkVJpRxH6qoWKqsyWB
dZlkfPijJDCv5OBqGoHJXFynbJeEAYKJP+FM7DB8bpNp219eSjVnqKF8LDdK
IIOedgZJ6Bqgq9zhBQqcKHMY4+PXHqgocmrXDhvi8WdEuwzB9Muv2fo77yj5
6sw16nxvlOKk/6h1BoEShlSGBxfQ7xNqZTPu+Isgbt3JwlEmYymalQsoOsb1
zhWtLaUM/3S1zGFehTUWvBfd2X3NgG5nNynH6X5bMOLRZu5jcFKWzYSyAd+X
jq+mdO1UCXKiKYw02I9XfM1e0YxVa9ngT1HuEDoT17zLPZ1GkeKSTDChE/mb
sT2nyPkt2zumWaYuvtVtmgx7vlclE8t4oo9YwoV52kv0/+jK4HKR4quVNXe8
jZAyq1im12AT8Zbwvm4ObNJLFuhgVlSLfN8T6RLryT+ee7v2FlmYJMTmURHb
QhHDvEIlfUnRs7osUjeQWtwBpc9DQn2CihgxE18DKPZTENyE/JXO33H3Y8XD
4dqMGHC3UzGkM6MytkleULFsB9yOMMj2VGddYx7FQ7SO+4q/YV2AitLEEK+Y
XAu4m+I8dPOTqOVHPLWvfi+TdpS79qwgF61vcqG9oetgRw/jtuMFcOAgUtQe
rhrau6ZccQu6LMpjDAzLeDkQH77y+JtQDJ8fbZyD4XMGtrSu+cs7vr+4Dma+
AoKJNUZbSlNtmTsnG3sAcjZSTUtXpwDH5WFQofgA5QffAb7nkXKj4Ink+Mpo
hiY3x7ZXhDhVMVDXwhUo2UXgoZpitTdFbmyU+oEBz6blO4COSyL2PcplsngG
Wd+uJvR3PZv+wSqSO3cXv9ughn5VhdFzqe8dwg/0pH+2C0LrFOpCr4Utr7Tv
fiVCYIxg4sSekaRoShcu3tlh3BDPesqWwNzPj5TKlnpGayiw4v6urpCa3C5W
qQVjSVS1SAA92xGsH4KFjSI/u5WHpQPpHs+HOOWHoGK5cOMR3X+IX/dwgasc
FOQ9oENVsbWLKelt9BuZoPF6XpXWA05IRQRC5sK9TaeTVoJ7ZEt7QMab3xLg
DDYtEYyXBvT8DGuJ8LxwI3dpGcCFXrGp4DQ9Lss3vyENyobzIQCYjJkeNi/4
xbBHtx32YIqrBtPEia/qOD19J5Zo2uUwGsh9yJyC7sgKdlMqtVb0iTAjR9c4
5fXpQQPuIHXiwCHdbUFUUxTPzpBrdNZPPyO+XN68TBSXoHOfDEBactgT5toR
PIAQHvp/PIsbQUqJu3cC5t8nQyg5ZHAjWwCBxqtB6IJGSIplaVOfO3qA5j8k
rI6cPy5+0rsfFBfz6ed608oprkTyEaxeWkLSVrmLzs2bZu7C6M9MRT+v04wP
rBMxEDm2jm9yqaYwX5FsfneQa+JKF/VoSylpl7cVT1nteJzPxNMZ4ZSqYmTg
PGJBXqAvfWxYQ/Tq1ZWGlJJ9zOKPApYoHz3yQIIrLL0LBnOPvauCuOPCkjm0
mW4V2GKJjHIu9e2fb+RCj533nZf8MynKFjVI8lvMyvipAREbr197pl+8Dj//
D8wmOY19QhwWtdRPE8xhiZk4hQHJgXxafuzDG/0arwfch8RQwtp2YRmbYNCT
5UE1At5HORsMTVYV4mzfe3+DGfv3G/hqMjBsa9wBMmTZI+k9aWidSFEAuQCd
cowZGkCvVI8jGHFbdwuwaApb9ULRlfBiCtlPGBknHrnt5dmkib27NhQhwm/m
z+WvYsX4lMYCOd0ZOuqTdit3WiTUEuDC/a6qc80yk3AW+7GohNR4N8+RxJ5/
hmgN8HqFFtdrB6Qe/e/AGa3PGuJYaeUSkMWRld51GFAJZuKT6F/GqqDmb4N9
9lAc6qd8UCjIqaTPoVvWOxCbVbzEBelwGX7uocpFRlziyCeSxVh3Dn1iWaTg
Qu4gWn8E7LUvj9ryFrWbXYA4AvM/40z7lvqAF0m1cymrFpz1QtBEnFSRI69f
btuUuMJtZFOX2OqQlZ6c+0tK2G20yazFDiSteBKC0tl5/AI7hzXV7ohup0XY
FWzl2ZEewwWHabjjjyKpwtTjASSXhWO+1C0mQOqJk7hV0gBMvS23t354AKEs
/9lmKJuvmAQcYjjspm/p4n5HO1e/cR7VErWHzKXM/KFzTaB7QTVU6gBBsLFZ
3v4c0IreIx3nw7dnQZ6pHyOJADN8NoIU/Ufd/SFgFSm0kMOiLER7GQ4JyXAn
LC/GywaW9v3G5OQK3+mkIobtSPDri2VriZIs7VxT1QXhdU4wsdbeMZQbPYKb
0uLNULiqweKu8d5y1hbZSGeGYIXZaAIQlmPOSeCGStlNJNYWlJglJrjNHU+6
Np5A3VmxksKmZJzIPJPLi+/CMpJhyBbte77MLoYdSQIo0LVfNc1639T+MvN3
RWHg6rtOKutsXnn9WLg6E9kcxEayKCG2Oije7C0ii6KJO/9tXMG3jIXin9pv
Q2+is6VuCMptlFcrcElbDx0nQPlbUUpMocQ+SRz6RXnKT6rmdqVuHndTVjUB
O9lXpQBmul9Xly800k1hk17Ksohm1lhfD1gMYQuVjOGN5dghRuet6MWp50mL
n/yeyFH3N6snqksP2iizy4axPPECGSxg7FIlPXPxuPiknkgiyjXsD7WR7D+o
19z4tePHsvxhPQBXr7pm5Hss/pYK8Knv1Zx5IUu5a4Wh651Yh5ciVMFOuXuX
BwpfdSg043K+Yzdc4Xpxw3RAnewG6F1nAaN/pA+vmXAy6Ya1dCuHPxmglYU+
sdQlcxbhCTZYncFDiV1by1Yt6ltSrEyKQ5+r66nsL46W8XZGnSp2hqoiB6oZ
Rc6kVsNUBQ+UytXrpahQ0TR9HgQvfSfYfw8C44/0KOvHr1iG6j4bQzvflTsE
eL11Z3jclSk5oaOMEpH2AQPhDUowZJrKpePOfxNCbfUzm7+MRBz9cPrupysa
H/Bddie0wqfWvpDaGcHOvg1eEX73AEjWCW+oa9bI4ZHbRN+2ZocrdLIGuPWI
VqiWrDP4sjaMt6oU1szSJ6/hO+iOJBE3X1Zm1heJJ0mBH8N1OldXlZKP9d1c
3BuieEDxWPbdDLeOKTtc4AzQz50v9Kxdhp9cJixoCu5w0p1RDl/Xr9pzcSc0
7OCePlpFbmofPrKmzw8Yh9nLcNWI/UEfsiLXA3X95zyMYywC+ogTKsBK5aVJ
RBzYqF2NcRb5FXcT0YswlCAfLo3lkWAeXwaaFg7jSHfygS6sCcq8y0FS0GhG
03CGZRAQS3HMXRb/3sYH5dhtLC5HAc6DOHbrfOAFbAcXvD81bX7UKcGm/CE3
gqh44KGTJGMxfu0JdX8yUvLRPwqbxX1YBSlQsGujkwXZWG3HNTo2X+HqFmyY
Za4dlkkSsaw1YpgdQzKxH8lKzxqnxZHtkfKqBS2I4dUi/lqYaUvIpwk8yyuJ
zHVYvu7/m4mcbIepKVC7hqmwCOqbve0qnn2KnY+ydiYMKcBksW/o0vuYTyxa
IdJ2GVB2D0CpuFzZtIU0sLNDEDjgjBaGqgOhAUmARXWVIu6snIxBz1SlxcKW
Sy9+FCvmZ2/pPi1taHu4fi8PIZ/anU4twDpks8fZcbFcdMmElaEBG2mBH9li
RtE1ChxUdVQptzty4vH6wnIh5vjLDmAJr5fF9Nkj0ox53cJKPbKIUhxHsFh1
mAGp9OfCTqqMWDbWfcf6AHfNQRnonbbZxuDdip6StEXPomygU3J1JHpCThXt
Rzjj7wWorpu1N9y2toEiRL+SBzIGkkP7FGBCPPAIJaGZb/Cb7Ls2dweP/cLn
PRfUxjbfhdSVyZGp8/x03ELhADv5E1nxEGplqf66UHP6LisbNO5zCniBfE4B
y6CbxPZe/1hHS2tjUptgrYllEyhsXEtLbW7aGk2DG6kyU6e587ZiCgFFELoc
DCUYYBlyMWfSfMrJKQahIjkyeQot94nsq6vDahhuFSSdS2rKAZz43IPcIKr8
YCCeyIy1Uz2LpBwDKaqnfDbiZ4zvpUkM+ORvhKU+ISOFE2UfLyBiFdVfJDqD
7/nD5xCVsCMnPpsKQb+8tq16MTLa/oCgXoxK9/cTTbE3tvYfMS5damco/rgj
b4mIqqQFCwNrxyJtpRWmA/OeN4IBeB4QbV1F+FYODBYu+saXzOwavnIPHGXU
oknPdLilTb9tkM+a1xuJyKxeTd23DujaRRuQOQ+sRR8hfWCBDm4bmkvsiTAo
NJJjfSZkEoPyfn3i0xwEqP3bTj6O+G1KYW+kmosljA0Ny8HwZCn+JV7hGBpl
DFE9No/cC9wio5pkCpqK+LOqZcK103Bl4I4oRTdKy/6Fr9qCYy//Lb3Muyrf
HSMPew3f7lsAOk4BFx1WaAunaaGvvzRZatIgT5JRQdbHJLMEiP8KwZe9aoYU
qA96mjB7HHlcDz4DieeegimXOmb+YcFi5sYt6DldyBsrlpDv2p5SHEtaY8eR
ydIeQNrxdhLZ+4APreG8a1gnhA4hBbtMJlFIV+cosfV36qcdUeudOZ9POCw5
3yN7LJc2cXStVT8nLVBBcMWzrwIAeumCL+SKUE/KhOx5khfeqHGAZOjzJtog
COSMqVsHpzzM4IYEbCu/xIV5m7HWcYrEj1lA0BNop19zd9yic7NYEjsOmHUN
jlID2XFl2EkkAtKWzErYDHFBcKfycSNptwhAU3hqgMFZ30yHOI+KcGu1iUYc
yIBAwPNtOfNvTIT8EYG2f3bKNBrGKiTryeP+ouUkYq113qwB4as46Y9+vrsQ
9EYkItYoVOCxB3WY9KwHvCfkzMlyu2oBHu7zIhg9IFyiokMF2I0BnUUG8iqG
inXku0sNdL8JwH7QxDE4WDPY2dRA5PQMNKR0uOWRtwOsdNJXLsZrv6vunoPT
xnrj+My5M9M1X0fNovDXOiJpesI9VSDjVAYe6KSeCZ+SQSLmUodOG+b6Ze1o
I87CJsO78GiqvyeFxhYCUXaOUhEVzQo0yqEWjossBJL0lEvSwLdOuY/2i3Mz
Sg6lZamO/ZySax5IBo4ILTcQIM9B6oYYB9+pnOYX5XOWzr7jk3PhRsl5OAQX
btr0/QKN+SoFEF48vnkIgkw70a/rd+QPf5xyDhwO9eSNPB1GX7ihtKudAeNA
kcna5/U0PsTp0LcJBRdiIlZTNv+OW491P2o1YxF/k07Xajq30gxNNsmTpzNa
hyyiouZJoQceWlESwA9qSifnJ8UIL+S3HsuzaI6XZzf8BdLVqfoBBu/x3JyP
FvsaALcqjMb54ZQ/0th8mQan56cSog4ygGTE3ARpkVWiDwe9yBp7K3ayt4QN
eQvsyPBs2+TiuVORP76CUwaRUJaAP5iVEORU72xrQBwDnV8HzbPiQvROM0nY
Dw0O1yo7kQWRRux/LwMk9oDAQnaAxh3Omluvmye14y/uybLA2z7y5zpESQDH
QmruHZ/nETcCp9x+ak0JaLFROkfxJLPXxKFUrWpKRUxiFSY1wuLYbyHY662q
BFB6n9SWdXRYCsYrsKQof47gLhWFu6PSuM7jCfy7LrX4T98JAyOTdBAuhouy
bb8VukGLKVIyArbt2SNeMowfIYLVUxLCc3y8XMP4+jukKzIyKgqhYOshIfMj
lEXmVdGXSFYZSa4A3um79y6gJOSemmBF2xRgxjqPlNk+mUM5wVE73JMECVdj
+OXQKD8M0CNVzBkP1kIELXBUpEax9vwUaDOQG2n3ZBkhRwtXBQqX2k9Apvdv
52aykn6nhNjO4px8dWggS2ch8QvACkblswFFBwGcvq3lgvnam/5DFRSe7j/T
eFwzSnsPL6uSCPSWBEzAutVd80t4BG+PqgGvh724yFCp6a0FzOs4gX+0JuuI
i7Ulfag14i3BQiAnuouCWz6xLSmv0WUesPs1ddyTuqLubP/1lGQcgsYh/zqn
jP2eUq664tzGkCEMAQSo9zlpsy/gAjQ7aWMZSmX1ij/Qj7BevmIC2qJb+CbH
QGM2xUNxVZ4se/n2xI/IPsNXE2NhjhbIF+uzjkVyPjW6CrOBGnFGCfaAb+/6
JdxJzVLQIaylvitb0mw2CKAOY47HHoy3t6qxZ8VoEW8NKB4nwblWhdZosIPU
LQ27VOFb7MaCn/6XKltnkrBck1Pn/Uzh9t0R1b2ed4GAPtuXw9lGwZGZmotm
zP0eDAN6XfsCy2xGgnhK4xNBPBtK2pMm1lBhIWGqGaYBPpD74VapT4UlvCb8
oUVMExdT+iUx2g7IAoc3JC9ve80fw9waDeABwd8l2i5Q3jNIl5x1zUw0t1DA
vKFoEgXdqSsuPEsM8Kl5EgEXHx9afXqFYNrFdNKb4LCoW2pukgrfjlCdCme9
orP9uqHRs3gbV3XBWMdP0SYRZj1jymP19WyrxdIhN+uWFPDz2COvW0ktJFAt
Xxpj4r9Ql+O/thh+hlbTMuJf9qrWgc3jTjQmhMfrJse8DdyTnZ0xbr5b+3aX
Uc1lxP43XT220aI6xYJFVDHrxT4VIEWF8PB4AhQD8GQ6uUNkt/283/bQL4mK
l3YBkujAF+zpsggI2g/ElRrg0p7ALQ5iT1bpTiW1HH+sSyC2ZoJv6K1eio/G
mG48lBGt8wBlktnOrb7KFb8cqBNS9SbCaW5KVkDksNcNC/Cf4+bKe/PJRAjz
tqDctqy3NlQB1N1VY0BxNAt3Q+9tgDL4zlmI6VTh9sf/CnulGT/tCEAKOvla
LN8w3HXqPJ7NJtP7+mkV5XXQXbot8Tx0ZMhSuTZSzjy24iarmDup4Ny2RTHN
IFAwzCXoQz8Rcj469atq+KS61s2MHnB4xug4bkXQKy2DCSKdBDFSuJLu/+az
gzlcItv/XTrytewxcXHTY9ryig6QZJM/82883bDuWTM//vlvZNo5NkvbDBUA
D3WcuAE2N6h5DhFQIVyBlgcW0jGJSTwFv7MVNV8gRMg41wF1wZAmbJtXW7Z6
uf/1aX42A8KRqViUrYhbFwsgVG6YLup+qqzJ8h9/RrVOAxvhYkOlZ2N4zlCG
ldC658BaxZiay8i3S9bD/9dQppHzmbKLTqha9YwH7Vn/S8Bo1l36yfKaPOcv
Kp4yVdE4pO7zdYtW4uyZt4Xv9fGfBc9+v9kAFCJBDusNsF2a926g8hJOvYED
c/zImS6xdtqE/BNbKnJ2/DdvshCr3c92dPBGzoz5dawLsYOtYC8F64T4n4dj
g3o8hCZc3QGPD/KT4k014EGY7sB2rtH1QhBndozm/o9JUx+XdMxmGwCZYxy4
uv8lAU7p5AzJW3RxCe814DEggOTaeFJSGArBSjTNR7L87EIns4aIKIC5DADt
xiZRzx2gvLlFD2aysl/mzGJg/palNhJ0fBZ4iSjgYTV8XPxKBhvJ9gJ34QtA
/FbaB7454fALwHRSpV9tMQu9BDEnstPPHFmumei5pZ2eyFViz7Rhta2+XQD4
TXjSMXaj1uV1Fo3OLzPYGNgAmuYb5QWKRn0G4rBof/p2Yg1CRvKcqJ6znNle
Fl7qjq3ySWFNqKtRGYmuU7yzjs4PsWwOT57mNQYqQCGvOXqhvZ0j0Xe59YMT
B+qfI7hylRYC/TBK4qlBP8LJ2hZ0NMQhv/fwLvYYozpAiB5w0X523XMQOMmQ
5GdgpNJ9G+MXIiLEBm4xF6KYCrSdIiVFUrhVisyO1VugmK0LvP7F8io1Hiiu
deS6X3vDNItlUvUk+AqhahaSk6oXF7ym2cikVwpWllG1dCGdA83Kpt02Td3U
Xa5qdCBjbCGV4xLL+puZGmZwksrMeDZag/XwprspRdASgvmLlhgeQw8yWeql
czN/qkDxbrd/aB94RmP7+WaJYdhSB9SZuXcJ9d6eKtin9bSf9OUbVOTXjrX8
Eii0rT6QWpkqXyNVGcAvnNnKYbJbUzNhvs6aJcyVsP1wUBs3Wwbo0E/ILYH5
OAmocYn/YXlSOyKo6Wfy5Dl6KweFUPr4Oj/OadOpKboQk68t069Zykr7eH75
Ivf9Lh0aPEbYzoi/0JQjfzpy8DbOSJi1KXcVcOvdbwcrXsY6Z+W1EwJOzPeB
Bqg215uUJwYsXE824hC9hgTK8AGvVuljs6o5RpKWt51nofOd9kG9PkLrQdO+
7cHrkrBwa9kHvUIme3E+6jEuAmBj5nqPVyPGKIH9Ta9TBvEig/lBzzRiXVtL
Mtd92wfsJWNnHgIP6P8JTn+F6lEFLWBlLPaC/Uc68sV1pMyxE2utKH5qcME1
rg5MoUjijZZL2Gw4Ul7JqGp6rBjVrRJSylYqfXOpNvMiDdYXT34WOxVJy5hb
JeQIsrtRm+RCwcYHAgtVlRYvla7J9QhRlruMhojQ0yfRlyNSczRO54f1RrB8
iYtn+SUEzJnEY7Sret32KupkbTPnBSX/HQ9ZUPFdvdxExNSF6Ix0b4r0KPBO
noAeezeQqKmiANIBK6X0TaHBLs/9AjwyxXnfMF+IYWFTLpOBdy4LkZxn3LHA
NzJDrr3PIIhmlfwzhQxnPvlylg4iAOn4rvyBPmt6K2UxcDqS2cebQSPxpxhe
qdAW6eUfBo7Y0XKjxNHEqqFBNXnPtyK7h2aKE2d3AVB17GLA+FzICbtYHxps
bIJ06XWiarnUTV7T1qaHT7F6E1CRSjsmpI18AaOp7qljcSYS80zAILJ17y6P
Wyw5Iyrv3akuPT7SADwJX9AZWF4wlrYQLA1tnuYKn0tzoTRUR5Hi90JpZm83
vcBspvSrtf0TuC3ADXY9VhZ/t7aLYnCJyK8xc2xzPv9YPuOq84u2XJ6qZSPK
Gx9Iibk+fI5EpyKrrRoB4omOtVAS4MGRO/x0EHQqw4qEEUon5pnh9nAJRIT6
+gIYMNn4yfl5tPJJodUMToJZFBTAhFdOKA+qJJ+pj2DldQEKHm1BJrY2uYFp
QQlpxwCs5kTZ4khCJNuASi6GhRK7GTTSr7wWiB+1EdLf+knlWfr206R0U3V4
MHb5fqJ4PfmqNYDD1D9pOma43VzcglT0Ibgix93VRo8cjPy9xGKHYTeGNuk2
DLLFlnIKyGaBT8brjTV8SdNvXLWnQHKk/isUkrz/ZmaaBziMOyXrUN1Ui131
4XfpXvEWNhMP+2HdPLu/OhRy9Mny8VkmDKKrMi8weCb9oQlZb1oE/3BYyLVU
prIQv3pGA5P4+zbCwRwumONDGvUzmkUBoLrGXZ+mXQtqmUxBr8RIU/JSzYAg
alWCEXDjhNpP/r18fpZBNmb1PkgGUms6FWj1vfQk8bV/8c3ogJsCmQefPLHV
jWYv4um2kw7JuKGgEkBrPVR273Dk8rk6UILNkpQ5Koize9rrMIT9Kwgzb4rj
Io0bzmkEZeuYmbKq8RjFbrl5wwiLxmtKwRLxVuFVMJ24+gHoh+VkQ/mlEfoh
6wP2gIfEXzGzt4dkUdo86Q++tr13aiLi0jM6vT0ccjsn5lnv6BCvfdC03KXP
yidMVb4OE07+AlyuzlkfDu6FNaNbu+80M9UB9Ci5STKU55bAOkdQiBjY8/c7
DSbi6OBsdMLZW0aAdadSgfbytpevwsFBtwL+BoqilSTTa8DXtQ8ObHJjFTAw
IGs/UxC8u7X/96+7VJ2IAN1WI3cQZRKAzeLZDlEe++hX/wTQkKlEpu3q0sGR
+fWNt+eVwKO3BfPvNaDmMoAoLfOHcaQYz26eH0ZTznHNWALVQAj00TaamPUz
ElcM4IXEH7D2b6epIgR/30OJOBxzZkf/rnasB6K3E9SzDETsd37+986X/JmF
sOKINq+DMJZPwXr8du0+KQA/ewQCcsrthGvy9NVFN3PbCW1V52tHm5emGuUh
pXhWEH6Q9jD/udikTL7f78E+bocOksQ1ER5HTf9w/CcbiNpQs6d7WiXecXG0
Oly9YW8LjzLGYLzETboQ2RjXZ/LbXB30awxnj3yusHDFu9saepvFzv29NuRK
JUIF9LI38Bt5GcLJ3fUshD4wGwWaw/+/ScCARBqAKfdoBveELiaKOtpVRcFZ
qQHOm264eessYG5Z8i+cDV8LrlJYYVlPphteBOX/j9nCgoJKtrahAL179mTQ
ELOnaaUW9DOLYLwIybydzZSp+fHeDrb55ls21Bkb32cAQ0e4I2+/mnW8qjZF
HleSj7WoeMcT2s0FdIbK6Nt0RJ+vLytbjMxejIZ2gTRFAEDPU60TKt+L3K2b
x1f4I1p+z7QweV15RIOLYb3XZN6FYk9skN5Ckox1anRs33I4JBIYJnGy5n12
D0n78BqbemWDD8WT0WnazLtOvVSqFCO+xCYf10ui2is9b93iZ/sm9xyBVYkY
dIG9tUJV874tiI9DyxgP+h8fWfHz+Ruci7FioTdR55ixJdvGDD6P69QTGjJe
jhjH4GZ2Ldm0Jy8wo0hQYlF9qrAm0c9/nKDg7WXzczftnokOpyO5OZFvtCtx
4NYhmKT/G9hGkH/NFJZWXGo6rzzYHAIq/K1LJpTjuZ64OY6IZC3iyD7HTTJ+
X+vmG1p9nhxVyB/L9QlETDu942wh1+vuwyt9Fya19q1AMJMhoow3wx7CItyE
o2jI9lWxbGpXgIIuVRwjAR2t/Hjm3pf0qmt1ziNMg2IvNLcr6cd7ISLhXBnu
NA2IxB40hGG/UXymCByiN5/KqngJk/pjbKr1vjYxWLsh+4Bw5YdXjwPlWbOi
RYLlmLF/J7ciP1+K9JRJIT6h3zQ+TYk2K1NOfgO8E2PLprnE6AH/WQEJa9FT
MJkudV3SkLsEzvfd9TjDJNxHgCqoyb1T/tVWLhbn6M4mRjAwMOUaofV/iecv
bDtz24/NCVUZ/F59md6v3lWDfVqQXMQDpnIWcvOBUClWVQ39M+E4Pw5xnWUy
qXlyPIGKhHuD9CO3AJU26MkyAR5Y5B0pcs78JQQxYnd8osnAaqW0Si0auVzS
swR5pa0ZmwJQbhCz0ImCuUIqGqR2lkrB3ibo9hSwacZppFkYVswm2L4U5p5l
QDdpgZFZkpfxl4h1jfsuFAGJA/80WM6zkW/MdR9JswgS0vF36DcX10TwqRcu
8G1W7wgsoEbFGAvDt2xyGk3jKAuvbMxw23UAbUQ0YAt/Dq1LSR+yiOKj+hC6
JHzvr0Vxx0+bFONnL6fKLGHdrUyuSSftvgucJoILFjx5+Pm1YZ+F9w1mK9hT
zsxB3x5AEwjJnQOxvdKPIKvdRfbGsNEgnnzdHu/z80yAt8sVe+7wKXphxbTx
0veZdsrOfF3lS864sRLWkhX5Q9M8w2RUOjlIvmdCK7DXtyGAF3JktBJwTbmQ
UJ+tN3/9q+XZxGRjSu5m+psxBFVGdZXkB6tcBfxFvgZJTCFVXa083wcTmsSk
ybxJzjNZwCr68QwIKJxsUkw+pSFBJwFn6x9Z/1X3ze6lo/BiZXu//a1m84An
aLHYAZtHeui+NX9uNAlEWyiwIgBU+sqFOFZdKBZEKY+sDe2eRl+tqmeDjNO1
vhzSWG5yM3AvnCdSpe/LlFHd5fYEGqugpez1YOaH73IXnaMeOlSj3q97pnBA
ZlxCLP8iVCgItY0X8Tf9Dw6vChyb5T4wyWAnjKyPc8UWwov9eRKkBclbK2JJ
SAjplxh/FNbjzch8BAMFvadc7eJlW3Bp562Tv2GOP3jNAmK04tWRSHjjkF2T
EiEmC4EqCsRpYP836DChh7exfnw4MrBti2nJRKpJKGXMxyGEeWcu+L+pV0i8
VewVVTxZoxuI9qtLtV3uemTLAWD7AXnj9S/Ht9ZKL7CTPqWcd0aejU/1Fz/X
aamwXS8qSV9PliqKBqbrREVuStuxpWJmfTvdw2fG5n2wHBd1KfCGqv9MDzz4
CEdJf2GtuTngscL/8kNPlzjOG8YtQzgA8Px/faDHzlK+2+3QESBcik17mekN
Q379Hg6W8GT2jITybvcs/4FQXgFo9yN+Qlm3GhmlpzMwLRp3Nc/Fwd20oAMm
Qc+LpK5XxuZMyXpOueUzHDY5ze2KDhVrI5e/6ybpZUmvEFs86mlupOtcoxr8
FQNeEyHqO/7JtpEzcMgaMBNg04235OG66+0rmiTtWkNlFDmAg8xIklgXuQVE
fgFXogPmVBEcH9EJlDoCfrzEmNgqwe0G/tl9c1guk1Sc67G2GJnHZX3v5FmG
NOeYEpPW6lg4UssRhEq6vbSUXvp4EHnZ4J5KrAnJFcJoZmbBZ/182sNHYPHk
kUk21K6Q6Rm9vQQ+4KS24nZuqeKsVI+kSFKZ2h3O90bveyYRsm+nTKeEWR6i
hcZ0l0paB/uTM4GdEAH7Co55x9CvbPz+h0xFeRiT6LY8vrv+t70SEk6Kw7aY
VEkn/lwGiLuwZjxtx2zDpk4Za5Qn53rhQIj3bhs8sUc0lE6uIBdcLxV+kq63
GPAR4D1HEUkz4B2BduDyy/JypAB2cF+XMccNdojDRLo5UmhVKxuf97CPJp7/
2be1/A/C2u2yOYyKdnxmkIudCP8xEmK8quiwdXW04C4xt4nvGZi5LXRLmxo5
rMSQTgnxsm0tHv+dTqJapCEJZMkKASh9zws/4XibcTJnb0YUxQDky183XGyf
Zyc/QXECzCvTb8WBeNPXAZi14u3Ad+k6OerHbnARfAbsUNMvYHfdUuN2tnDI
rcN7bla4RsgL8rMNSjwa+uaEM6hRC3P4/VZzKAi9+OTguA4bs3XRHrYI05zC
sA3MtPTJKUGPdD26Vw5IBLbGp1sh4qKEhoUW91jVTsmcbUNiZJr5c4uK98K9
IOJNXbsDm1HMblwbfna18X7G/p1uMebmQCICiorq554RhCszXOgZA6SFxoKK
Q3AKj3G67dT9hntJGWBnWe0TmlehxfRe9EprpiadvbWhDp52k/fY9TvQoD9k
wmsIjzJMtwyOCBiadVhMEZV+GsJjkcv37EuRG5auJnJv45xxu8B4JwNs+E6X
ZnvNLnHUIq+uFZVam8d8nN+UpCrwys71v3g7TGd0o4CgsoAH+x3hKMyFWGuj
0921vA/f9MMXd0FjfYg3QtsisxwlMbSWKvlk+Igm7tISCuEilB2Oj9jRM471
Y4tyBVHK44JOzdqe+qGDJxXReUdWxlK71L+ViHjP5KrItENRkINhNv0d5BbD
ZYT/7A2xquZ8oky6I/413MZjc5HDRMMNrnelAosj3Ad8UuGLfGxsnrrxzslB
GKtL9prG01c7OYNFJYyqGJzLrBMsQeZZ1+0iPGa0Kz3qoF/8YMJ6W/oK4C4m
QR0DmjJQnUUkYV5diGiXvD6QXyRblBoDYTpHnbBUgw5WQlGsuTdhnkonhklo
QIcPkehO3D5LOnz6oWaBEwg1bmrLPHIrRtQ6VvcUIE1OG2Xqvzu4syzUaH5N
o/E7QFHgpp/4er0uLYX9Osn7RrNbfvzs5yWMw197Ih7Ze+yEd7vIuuBEhf1Q
GtLmNMDobWB8fXiB0V4Mk3/wEi4KxhZEoVBuqPf3yHrtCmwIqQ0VR3ADDv3c
+ltPBwYXUeUkDVoBXyq7Xd8gReTaLZ69F423EjplCFp+rpwy8Fxs72hIYxJM
d9e7PiJO3byeYy9loOcQ+K6+pAxax/JLbQCaSQ6ZjGrruUvFa69SLqmWzIfC
ozF0hQT3cYKkIno+6Ezzq9Ixy4cYUgWum+zXSNHaY6EQ4YfptIVdTcion/vO
xakxNW7hutLpnt8qCWjmkrIVbz67GLnb4obmOsBso5yxEd6db6dbC5ftmE/c
VNnu7MAjv3As1VfpSmSyfrrTScDib1yOIBtjb1JE+kRTy9cfm3y5dfr92G89
5EZL8+BAOaLOSTCAGgAb/2TOPE4YcBOvi7eZj1pB1w/XqFT/kI14ppc8AYlm
W7sCu9DqIz2Bv5vYbyhfW6H9WgDkTDgtXF/X+/T/ciwboKs5unasO9jrvGFc
OAvTQ8tEBtvAXxOqE5jFVULlYu/lOiVLNo6sDcMzE6GIGakSb000UF0mLkmX
eG2wWLBSh+PL2d26TagSvwy2RPFfPmVP83gJ2ftmgb/vOmgM9AfUHLR6BhUf
RReAg+qcKe+yfbq8EMn6TunfRB7bAGesbliZSanTH2Sd29ITwLmiNmrpEj4m
4zaMv4AokWkOfFMDrHnEW0jBZbrdH3SqH66x2fX/lOpS7uJyuWjcQDpnjxWV
rmOFfVFgj0IPv3nJmNQNwtoMGvgibGmVVRBAEvAUU58KwGOBcEvgzjwej5uv
HUtVW9QFW4c+kXrjz0Lt29TIGh3HyaI0HtJQKkhzVi+VYKjH6ObcHEm04zkW
dg0NBWvIj8AxC1Q/PbDcGSLvMHLqqWjaJsC9AZypYhRgv+eb5Vp1BV7H00PA
fMOMPbM5gGJ7jjBCGp27dJxkVPNfKCKuwIrTTQS7igBP+jvz8a3lzJdnoqyy
RZoYewxCx8RqLSJPQJbMebks7rg/mxnpD7Y2sqQz12XGGO39IB5mGGIbKOgC
gCJ7VS/WAl28NRwdVPTI+03RkRzU8et0sMGtHPPMZmC5Y2cpdD/iwoBvokFT
XTNlpmGzsrCs7zT3oLWvSbfxWfCg09KI5AvueajPMU3aeh9xVQZsHddJSxc0
TNMmJQKpPP9bD0uZJCfJtZr/yNt+a+Uozi7fScu74V08qlPpgO9qEKRr5qNE
t847zD7Uf/OXeNGtYGslWgSrDX5Sk4NDMkYGK7hrGeOav5H1AZJAsrv1MPT6
5DPWg3tbAzJLVB8TC3CHA9iWezjHmfrQXUNSjdOw9P3U6nzMaGZsVMY+DeOi
gJTMQ/6Ag6cfFvBgp5rIcI5WKWyKxHata7zBQ68Z6tI/niLKZdL/KKgrmvl4
WRlgXr9URywar37dNPbpgnX/ICtsZfPKpcZMyLbB8SPlgQ8wY2GY20Zcg6LA
wUz5j+RbWXA08QqiCXVFuO6t8RBdGAX5XeL2yf/XNzo+P6+9t14rcvyeljDP
NWKfyeg7ot+njLi8GwH1rSVJAD9BSCYq1KJVE/GpEZbMGtuBrc08riLspPeW
UQZzrXPustt34MiMTcvpvgtLzN965+L103gZfLCfe96mGlsKP8cnkeWeu8do
nrjcK2p1UvNMA0d4eYOGCy0LsxQ912drKqbC/LkPsPoysHjGLsct3m8Gx6q9
HceLUJ6vHKRwGUDLkX5V3iA7HDzLN1cx8fhdNKauH9+dEYByk2UQakpQjXBa
Xwv9ceDT4A6qr+YidepOKZFBeCWJfhAo5Lds8LPRp8SNIqr2pYsLw3rgogkH
hQI5UMewdRoGQXohY50Vx09Ddhw1mWw+BSa9GWG8fogImyLVb6AeWbl4E7sP
Nv2buz5M3arGX+1l6WVVvZ1bo5+EbS+f+K/vptOz9xFZqP2joeqVByNv5MsL
7VF5+PHYQvQF/89iLmiFljkqVJSPZOQqfOmWThVwRLM6aIG+dBmQs23FYJkI
FP3phJwsvmLUilZyavwUyGRM/Y3RxVcIKOBTCoNWgZGqAiJYB0tN1dtNmMlI
sQDPG7XCz2uIv/XyjwVwku5hkX1iWMGlvO8A1X2TAwq4R8ZoHbKzDaHEIkdn
uMlEtq0fgfL1jb0sP1mxD+f3KrRzmYa+XhsvzNVJoegr/20j7R+8zy+H8whA
9S8+oVLeLjrM6TAhIGwo5oGGgmBUqdyTUcjlYZUDmgz+teYYs9IiWrBFA1bB
Mv6jBvhB4p0NlaIO4DfmDoaMxYoxtSdJ3svTGAb0xGejQNCRadp8bIRZp7ER
sS5YFCdl1X48E55yGBjDLto/5ns+oXAhZHO9gZeEp1BeWocTvngPuTJX7a8f
gtHdZ1l7EkO23ZUjZdxdpiUl0XEvf+QukvMKcrKbvLb+QZ0zO1MRgP8BBfZ2
976ZYaG3mEbVaDqsWgkc8C9Sy1W7+G3EiOoR9xhPUvb3PgAPrgmqHCzfdczw
uumQ7Orham4pTGoBXmBbGqakvzzIlFQ1+A2b+prqDr01qj7ndVBzjM1aXdQ+
sLYs1l8PqFIsdCW9Oz1Z44hJ5B6xwmIIhHvmqCVkhRHfANUJsd5rDuB8kpfL
uCxIOtmFBQ7m2wDTJlxC/ekffXjbRly+v0d7k189cUiHxk36C77FUOiv8iLf
5MIOFkBZI1kT29gd1IXmm/MKWd5NAks7yOYKK7gi0hol7AgNMpczczSKBJ3I
1qxHNNkQwhgaC/1wsTF4ZkwFbIxr8w/5NSoyY/WuhidZ/NeSTDf5UyF1nLCk
1hj/kH0JUHXuHEO64JkuQ/Vj0fzWBPZmp8CWWtii2I61fsJfBVvDHHXO6g0V
695GsA2Nt29l0qlsSnp4iwxNtgpQ5V4TCFMppFpxKiAl3A8MrRwzZ6KINq/W
itogbRXiIrUXriYCVfTS/i90DmaIVJ9xZTZWGi/hNQ0h6tz+o6gT7p5P/6nR
iSLqll+/hPjs9OOEwQ8jBiiGwsf9wzRIWgjdHOiFFT9JF56SuIEWlNgOeLr6
NQo9qEI5Ud1r+3H1mAZpoOFb1K0aSWo2G1wXBQeX2ioWFaa1d7/G5zxZ3ru2
jOk5TcRmZWfgZwoaIt3u6wQsvpiHdh6DJ1N3q2GNSBgB6ttBSPcE37vWcN7Y
SnaoGBjYWE0qvPuSwejXorAIeC1YOqIdBnNsGSpiBpcofOb4eBZ1IEsA0zUS
tl7SYZ7HaVblauRe4+qnZ0+o0ulzNOKIGC+0a4ymIA4CpsWFyvk/KS6LLjkQ
SCZfl/o08DYaDJjt4eWNFc1PziIHqiugAkSfH0la1HjRZTmXst4e5ha1+o5a
9FBlfXj9m2kFYp9OD2QyN2E4n/r7sBgBdpvrPFEgDvxGn5XB3u7w6l+Dh/J4
cys8e102SeZx3K5kbBgDW89PiURkOXSNfC3/atCXT/SXSuXZCH/wOetJeOnX
S3ICHspM0fDijBJ+OK/5TiOM2WSiF4lJc9V20rHh3NIRK78eVCMTuxAJG4fA
cbVbnOHnEdOIuAxDv4vMPIpQAD4i658vDupQG4kN8AzJWleY0Ki5FXAjfAPA
Y1nP/Gr49/H3DxV05iaO11jIeRJ9saTVzs0JMG8HaZ/YEB1ikAF7Jq09cNyl
WUMhqmdsK6pLf3Hu+CyhncqreNQN5KtKPWzLkHAiEwxJHKBtL7rPxZZvj8Mp
VJ+YZ6TJkFzYn+4NC9UKFzfiC/cV5m+7+DvZ4higpuGdjqrtOEFtosEh56gb
fIT65B8mzKMWETywhKFBNIcY38bNbpkYUEd9bNUyAar/OUA9vZHaHb+XxbFr
v6m2Vxm0dku6+Y+ahgfTV4Rh7bMTtJZx6+AictYadOBGcLugK3pRoJKgKkOi
N6m5+ZNyEuF98gqTWwqVSQREqPc89CGS1GJEfwSD5mQpOuUBtN1dd/vLcHee
XmPkZcifcColfn2F0u3LA/hRw3ctntIAPcx6ohylEROnU3z6fwb7laQMfeqq
l4kvy/eh/nz4J2fX7M7faayx/UpGxgBzJ8I+o5qGrp8lOUxdYP8eAUO5fAWH
DCFd1BhX9tnKM6BnpuSd+vyNhXvmQvvh8hfw1ADDrHTUjBTahdv4EyuQFixO
zUk9nTQ4s8AJmsJZJLZxpeSZULyamJADng/WuTN1uZj9i4ot7Y0FxijssDZz
CXMh9dqACmQ3FpJq3hm8PUbENmKFZpQFO1bfcXPJDaEi3EkSgtLrjQsVMuH/
MC9MDYdDLUqESTAP3yfP4c5qFjuboEH+9lPH1ZiecLhLXs75ayweprMd7vbq
L578FkXxlkaACqvkXDFEh40xBBQU99z2O38pYQu2/91v7xQItxJ4tEn8bPJu
I8QtKG3qBoWU0HWvfWOYQ81Kqq5Bp5J6TMLp8dXbkJLwWT75uVADwDaFYeTm
JvWhenwCbRQGBSrtS810vcmvNT8hsVTdC3C0lGhyxamQyziHS+Us9m9Nk3h5
IxWPxQ9AoycJG9ToL0ScxA7XMFJ5ziQsMBaKY4QHDKjl+e2gvWMA8dPE+YvU
v3xioNzZdmUt2+D5Yn9I6UiIalax0wuBKaV7erMnhkJ0IzrpInOHZd+qp1GH
zSkoHDcfwlmboNEgqvrx0WF+1zLsh5snJTaIsoLsEZ/fP68v204HY1P21Luo
vhPTceN8u2nuayLWHNHpPhW7NTYcC/5DULLlY6cju7vgYAX+PsMJ8us6nIg3
vmE0AHiL6b1Nck5ag+qixMnIwpKpc1Xk2keT6/Bb/VzQUfdLeBr6ValbH0yP
1vQEr5P/G96jZtYYXcL5LPmKe1Tj9rEUHu0na1242FbxEZNGRXkplaY4iwpr
Rt7TOwStN8+6y1MkcRojBjAnM7/p+6IT26NoDP9IVsEGGzVg8AOW++keuUeM
JI7d4b5F1/2JUEF6pNLmQMEGY+B0dBp2qu57bc9eVt+87j5YKYyMXZqi2OuU
nr9zuaEP2CNTGKwVLWvGLvnDxLAhMU1hu49WYE0sfM7pG9BAwzYJ6XRyPh9c
TKSqVnxETOgVN4UC+WAD2aRv/h5jRYwI1ItVBput7czDzoCH0onVMy+8M4w8
WdjEsZVXktgK6gSAN3vcBMac447RlP+Tu49N0CUP1M0i9CMl8wdHHRxOXHUc
0E+WxeKqSBNENL5dnwhmW5J+GkOEOTIBX7XZmwHtVji1ByYWioaTDUqQOeu3
g8SgHVkzN4UKiQinnVkGkfDbAYRVQNT3uRCVlqtI7BhDtSuSXDy9oZfh09mS
8/Tq29VGTUBwIuTPL/msmGdk8tznKIQMk/FYtZRtkKqWKdznye0WJj/kNg3Q
7EDDdL4FiX77xoTZL+1f6H6VAiBKL4BnbzQCT2NDotocm2Wwoh1h4p47yqyO
l9w1bklL9RRvdWLGi3qE06LXtkdppFsnOBD2YSVC+snG2n0dkpJvtcm2LrhV
v1GEuMPgkvthalojFVEFIcElCcRs+7DduavM9g63pgY2Ab3SEZl4jA3PPpkO
kC3l+NQi5Xx8UtYvQOkvoom0Mo2mkpwVCLlU9kMG4upOKFQqZX3LjLcXyXGC
Xp2HP/4ud8waCrZ/JjkFy64yjSe3eSqE5C6x9hTZBKyNlGhwD6DPDCNjDFkk
YvCHpquAiOn8NCQ8b0Vjh3BfcLHxprYzY4kqUWAB/rLQdJYVIFC5QHIgymsI
bbK8+p+c/R/E3MqgyZ2m+9eh7VAw0j8L85tdGOvhk8Qf1AYJA2CeBHi4yqjj
rJacXnJWeN3VIoNf64jr/zH1lFU4ihRjSPLs5h6dMoIFo2Xn3jzD8Z4rSluy
dcBh2SipPZwQfkgf03oAJOu+RmJCdCS1f3722hYC9//AxpeACDNUL1PMG1/m
Up6VAeAjVpUsAI1nMLJg+k4MngCyqGgNf2tlk/eStybQMXKbsbbjD4m8C3sv
/S7zmE9smyam+HxYuaJ0zv36yps04LWR95G5H9pz8RKM9AC+6uGmJ/D6oSsI
bpM5oYoSEH+x42LswTWqYn5GRxNYa++jpnzI6xJU5M4grcHCk9iCiXMULpOS
VfyTmufM2UO8HF2u642D+VQPgtShTtjiDmEG+u+J83feGF+oCPVNmVyHsb2K
w+8nTSE7SDGFMfQd52nqcsdYv13nrSJXRLpraB4MQY5H77KONzxi0pNtneuL
a8Yx8aab3e6LbBGjTd087xeNBPwtBSCHkYjAdUEJ1YbgLBInzvQWCWxnxrHk
+pr8GzLhG41713SYmaIPoUOa0GOj+RRz45YA3dAkB67TrGuFF05wKQJBxSm/
bClgowDEYWkQurUu5cVCESWxwygLfWZNepvoOU2vYwTJb7HGVgYWyEJSVy3S
FpPPJPJlLivGhzYsKB1A5PJzQsVJwpOQN+HiQd2AzNQMDKagsuhIYHWc7c+3
iksypQVjreCOCrkT/CEcma9B4Y1IUlB6FlgWjoHXEETqslcENcbj8hZnnwz3
sHerm9Lm04AKoG4WvN87x931rZ8BHUTg3cN/95YXjqyEc13+BDQpE/o5RWF/
pD/1d+MK2kTcaNOwhp8IvPR0ZpmAvGf+BjgAomYAybZZoY+lIykhWajFrw++
OV/hfvnTwNYyeJG7ULg4xTar5QQvq57Xma+jS3dvo1Ri9LujT3yz8X40hH8K
CiyCEuPsUVyMhOjXFXSf8/YusLIEBbnBPBuYyySST+pdVIeLX3Z9ODSzAUX/
ZG/1zj3qFyvEBnE62zJt+yQrkyLnD+tOTe69vBAWgxmSIOccSqTJ7YBbVar7
EdqsOMo4rbXRuATi2/4YMIXCvyperMQqJZ6n9n+utzykjJrSYkcFPGO5098F
KvTfTu0Dfk2ui2qR+76ztcbU9VHAN0hlIuMuYx+uymxBcZkTl7/bLU00bJJW
y60f5wn9/NMb+ymGE5O3quEYKbgt+qBDetxWPWQ/kU2RfZOJCSwjfjztQJbb
vrhL9bwRRLFhUzltNIirYL1fLppRvq6VOcirNOJydY3HHdjscBvoxFKsYe5p
fCkbZNZFT1vQ84cCH+dHraKvES2VMrygNDig09k2JIrKO8zj2q1HsLzWeiPG
vIY3yqZXcoJO0Fo/BcKdY1M9mWJ/M4Vb61z8E/pN8heJcFFdlWouAWhftcPO
kgnfKv1CIyWMhaLl2bWmgjnguzY2sJj7J0F72a8axoxvkQMmhary/pRZuTSS
//6CRWycnB7DoA0LF2BZLTEstVn43Od0n3Vf3wScvEJFkYwg0Frz6H5MnttX
8AKvTLT5Ujk5bbnFXIO8plG78kaVttWWs13MtbTx7X8WYHDVQEz14jmt+jCK
D4UlnIN+m3t3b/KMj+eaCCXjNSzPsnhruGHFdNiAODxSWtqw6/3YYEGwqXgn
0ig8koeRvsQsEJ25cKOSjBArKVQ5vbG0VCqMFrpVl23YNKM4sPMQVX/Wh9tq
UNJ5ezpw1MQGPgDOky+VQUgud131zLkpoBDUsIgS/dqsUZ+xmi9PSndX6ykz
RQx+D1lrARSevMca2nj7lGMmDST0+7WLS5VCUB9lwRpxCqHcmWU0ooLHBbFQ
bnQ0PV93HSopPvXHtvsT8q0NIL2Pvx5OdoYFl1yABbQH3QZwAJT3RJGRK5K8
7+BDSQ2vFiZIF3UnIF/Hthyg9HFPBrK3EWKzMnpfT+jxlU3zQOWPTxPnbqz9
gwDF7oplGVZ4GrzGU6hl58oafdWX4wwqh8dgppFjlKUtrFokSZGFGWNlBRtM
sueBA8hYzJMyq7UuXHpMD/4d0fc9+qJfYIYTrBzjKdFlRcXw5Oylr12GKr2s
IamInYTyxAHsL2XZmgY/nUZj/rUddsxCiIw7G/bMXLRkqB3itWxvYayWvnlN
Kjrw5nMlAI0Olmj5xmtrB/wJFcmm1YxRBZU56hfO9S7WxINqbIMdUPruTrlv
z1KX39vsuoIe4WpusWXpAsfioZTkLUHBEiKYfI9I/MWzAJZg/ov1YWRvigNj
A/mS/KDloH0pkfIG5rolLniuPsyI8T8zD1j2XAW+rLcf0JytfcXK5sXY8I+a
VLKBdOGEBp+YMw3+gPAmdhwXjhwunRdUnb0P/V4dzgjkKF3jN3zME6Fp4XLu
MsrpIN3i9d9lf5mPi15oYvc8/IPjqVzIA4DUMnhRMIuW3VLyrLe7jzE9iJ7e
DUHAQTzWIcdAXxU6fG+z0PdKileDAAizJeb6LcbNktdSKNM5julAKQsz1Rw/
PLXTRAWseOfdNl1FToMy0+8zC+O3ROABE1qA0/11q35sOnKxoKsOdh42YAeB
0Ci7Uqm1wGoySi+fVkpj4wSg2GR04mqGKoEiS4aV9CviuexQ4RMQRr7wlVbR
NhwtVBG5IHT3rF6iXiSlskK4mxJr+Ge7nd7RIsgPvUwWClXnwzCMkBKpGMjP
rVQ9aNRHPK+DBiwmVCkEsjkn3fWU4WNFhR17P4IH8yMsN43hIjUCaFfh5pVo
4QJkCJi8nDQDdr5QFJtTunrJg1tcoAZEvE2a+4kjl5D4NEH7Sk4xNUxqgE4K
7X2yxlU3nCQ2049OEY/vXq9qrhiwnccVNfIl7jihYV8CRavbfNEcLtyH2s+g
ZzMHxOdBrg+9ChzJUCgykl/KO8Ks/lcutD5OzbYVVpyf6vCG6+MZX2Zzd4ZK
vG1Ee72mxAxfRBwQU88Il0K3GRLMufB0ze02cQAiFySkSdLPfyoGsmI3UTja
yIhTSp79n4rVhY5E38Tyi39fX07h9Q3/NBek2wD3Jm+baQ02Bm+mJsT2ft+Z
VqEA0kVkWkcAcurgmEyYpLLO2Xc4HKQZUtUGJZs7ZmuIJ4W4PolQ2k8H/BNq
pRg6TfYlo+UfRyqGJUPgCGsoS7k7cqfATsroxptpxb40/4aHcLKk+I+xYdwH
748fiyV77jAZi39LjJjf53eiIuyAm5rdmWBBH3+43ge5aRFnl4QI2az013PZ
GOJdLZg88nG3zANi+2Tsx7FRYMnvvg/QF/PHeIRjNr10oIi7bTSngtCI6CwQ
NOi8Lg+MLiaqcqRhUJNFZj+10QVIyiFk99xp9IqQUVQwRm8hZL1WxOKU/9wv
KINhI1Mte4a7ABMuNAFEFvBAlZvC3VAdo7mg3fjfAE+I2CmNMPx5FNwnjV49
smvvtgnsaQiIUea0F1t534mbaRTikcDpA0h88mifK1nFAPx8IFP8UcSPCFeD
ibx/gvlzJkCVcrkje+2E8DgazOk+w8w1y2LL/wegUZOLR1I6UpW1BFj1yHL0
2brfHBgGEv31OeCRLghkdSqNsx1OkQYDN3eFBvBHXLZe/DJpSGlBCuRVoRTW
47fuw9Ymid+t0sJu0bSgadmN1FrYJ4w2Jys2pngg1Lsz6fcm/zIO3pA7rE8k
U/1/uf1uH/Rzaf8bX/yIJeb7iiXF75rPangEWBp54XPr2yhmZ1/SOPTZc4tF
oRROalKdUKq+5FgvYjENqLzuJn+FP/Nuh/dPvATtB2NtSm5RIfOChj9NxG1c
41/JiiApagRnhtK7VE+h/Eit8nuYJKG2AB4XzWnP94dEzmD5GcLgJ8BIdZPr
Re9926eskHXFFeSVIHHknFf/tQDptpJL0y1BcNvgZI3HDF0L0m4oKzcWCxph
kLs2u3Ivm7icSoJqWPh9cYnb28dkpcZvX29ZfYzl+IXjptJNoHTS+H6RNyZW
Ot/BZ/T7K2evk/HUMIAxWGA/wR4DWgjZtrFs42FASEa0WrHyHacqAD7moV5W
1tkn1b2pFQrk66JdUykKKneaGeafyUhUIcycyqAbWO5E4TWyov142b6ZqJSI
Au9xHoxLEEcSpBBLH0nRcSp7RafnZLn7yQaVqAxgEC06h2GgB2DOeIrsZu2A
eH75CIiN9btaje2uSbKA0rXnT07VDyQ9Ysdh3R1aDgWdlwMF4CKCLo3p/dgX
1H2nk/jfHiVmKs/boBA6a6jIccKev5axjrumW9m+bbPWSSo1166PkOpmDDK+
WPm5+bq6hkLP/pdet/h88eDxly/pB2ez034hwkYj93gLOO/naIrwvVRoukBb
mjuBfDES7Y/vV+y7j7kWsiub/AUnF44IZEm9zcQgz0dYsDFbOOSylZh79YDn
dbPlgWn6PSOugd/qZLlwQoepBAQl3RCulzhBG/4jjURUq+oml+uUFekZC1FI
6PBOWXnS9jDeEUFbaufgcdNH8uRTQYAGKt/RUUBUtjy5pOTjJmOYfQuG3VkE
G/BzL/l9wskmrnBpUcePTGLsHY4KhmiA2LLo0zAiCMoMmyby6pPD5sCa46e+
8PGoj23looFs4lWsMh9qXI7CrTT+6e8VNUKH7EjiKHrgbdgxcCrgfC2DOajL
RQPrwRoT+6XUppLPWHS0/etSbrnTlyRxuIZT9YdpcoHG34Xux635x8U/cYSY
vt0fiSv9GoM7m/CGPiHXgnW6ci8flaW6JFeBude6ijKZWy/GWhffF02fUTeI
nIF/t93z1CvH6zmYeGuxg6AkQ/yHY1uQevcGTjYcX8PeZ3Z8OS1RvdKALLx8
keQwxbyoGH68ZKfEhXh45VGoh0SgwNsCr3SixhSDgO3WWGzMuygwzIVfwUMx
aFjkMeQ+NvkQ4IUk85bOvaTWVHnVY7B+xm8HZfpOHlh45ANiJJHW+VFEutpH
jWNHoltDblDmmgcg+IOahnP3LyipAGzfiEGQj5EmADFrRrSAJTXkV2zXRv5O
8Td/6Y5K/W4IvNmo6zv004FvjyWS9DRqeoniIG3yiQtAM7K8yVN+zt97exZe
+PO6zFpoWZKdVyqE2emhqBGNOx9p4r2u2GC2apewRYTj/UJ//22cKA0ZIpeJ
fim2NrtDjeclkQog4QeuTJCpuVurPrvwr23I2xI61XhMo/zB26kK7eBUIhNP
CkjSR/BRBNOOXeTPZCgG9BEqN2+K+af8ZY8EA+8Tg++m1ldsAh9n0GExuO7W
m4rIT2/N4K3mxk5Eqi50I8WiRHQ4MXeF4NUX7IDOdK+XIT2VmCGrIuw1XGhP
QKErZ4AkRoXCmfZVWSbssOXQFyZmRJGFLm4C22z/o1CL4+yp5Fsp3SCWL11p
RC800rkpnFLj7zLx5lCz+hjMEmuEdUqHhqLHdeBXDG5b68cH03v9ka8MQcix
bgPWYpiGCTjJkTeJe18LJSXIbaiWGz79DvyRIhxIPKbcahEFHCPQA64FGGHb
ekZFRPKpSSr00iDDFKMrDiNBVtx8FvMrjTnJrOn0z7QHVbyER4+F2xaeVaux
oSH0UwbbKZa5/aFPuYtp24dNr3oZWOdFSnnuRR1nsi5ugIttYT4IFYT7W1Ys
PGQAKpnMX5ECDtxXBvSv456+oo+XE0wfWfdvlnE/zTznaSe5+sscScfzh0ej
9b20JELUcJDyz871UT5MkXn3yIoE9ETBm2UvAKHq60M1Be7A4oDm9WFvRQ2G
Qa58WCLUuaUwQlOpXSAgmfLOxuH6dqB4op/540I6qwm7pRtHM2SI5Sbc8YD6
LX0pvw/Q3beoER7jUaO8RXvfPNb6jlp9A0YKNLbgvF4mcTDgcf+DVSRTBK6M
zxD7ct8moL0XyyXoYkyJX8tiSOZB72gfl4cATOHrvqX/h7526O+OJFKWXC+3
52a8EZpsSGduwCgwtbNKxQFJgNeRLI8n3/O44M0Lr+FFQ3ScCCvb5O4Kf0c/
GQ4XnWHNKGvcLmpRAEp6OLZFRT8gb5iBmlG8npCgsF2kZsqCbeb/OyK4nYdD
jREwLMXKZqy/7yVFar8zW3cYx4Ys1bqiDFI8nvscTkSQbvyQzkR1pgSbxRMr
3ltJFvW6Ddkaip0hOlNsNUHGYDfpc4er2vK6NG5amTBefgnLjnoCQKY0+Z4K
EMFFaPrt/hC8suFPmYg+ea2JcSbLCcO0uIuUaVH4ihxrycpH2iNfdiiNVBrD
oYFi0Vs7L3sueQWXaDievrsSVMEXPvIwCiU5gKsGb+fPC8rqnega0+tnyNCW
GAIVX0IS+t8X2KsSTyFa+Q4Ds1e51SHz3X+B+N0MHEXGobffJU/g2Y2K+dbZ
tBDpAVZQrNpzynJBFLeN1BjKZdf3vGXJizDmIOCNs3Bgsj0Ub9U6lsDNvmRt
lczCryZbwhDEDaMtlOIo3NN0xAloWBdivBfTl7l5VF3eYGvZEgvtfF4rXcfq
Zjr8QyAiaNFKKxYO47MIXjNSc1y9rHhNn3pTeggDuqqSdjiJwJYPWMlvtXnd
Q2YS0fOcQOg8rQgFsiTvVqYKm4jvNIr8mn2P3t8socgps94fS2Bo1rjSjzmm
K/KFmX76VLd05Gl11DaOBEecYvwOzcyx7KAliqgp9XKPqU3BlwC4psa96Irh
xSuZoHh9ZSXrlUByonsZzZm0ozVftA/dG0xbQfQNg+/M9+ax6sIBFfS42fN8
KB4lwe4Rx/oze/HFGje6rXM46p+gB8Tky7zZVw+Ai90BC2mUdyEQ61DTTmMM
LxrvuxBLfnxdfm7OMOsJvdeLk9Zv2HAx+ZNogb6/ln/+UJkp8O8YVQY7Jdp1
mGuVsEgIYCkjmSCQQBax7IR93/TYN0xlJ74tbsP1fscTHHYpkk/Cxbu9nISv
o0gC56hhMGuaWKNaQqrZ3FvYBFn1escgmqh4TBNGfulgGlh/PxG11weBn4I5
Nb/oJd5FJjq2eXs3wsrYIzxwB4NCrFZKOlAP7C2Ii6YN6W5rk0sBZHy3Ap/m
ZSAmWqG6E08i00NtDGAUeZQblVRFszObOh4ZfZ6jePO5Qt/C48owQTcp0A/T
hfFja1bGAwqvhtEi3n3q+e0V2/hEUBpe8Z/4Nx6KU3rU67YDlMsEpB/2lC8k
7CD9UWwdkqULg7FihmeUzLNT/rVQrBAqMRRXvwYdV+VIkomrNfgogP75+bJQ
ZDyTpJnT7izxL9wwQD3PWJofbHsOLXr13QmPFIp93ZMGbuKGioCot/zJbnmS
ST+JeaOKJCB6rpXZrS8vgqv7PHF/Uqkc2C9zVZ6QKmOOOzV6RhH21aOFZ22W
ejJNgvU+C6PL1OEjWocfcca/l6i1kSMlQYiSGNU9u+cNQinmH9s/bBi7xivz
K3VOIRVFJXB93noJAYRmQXLaOkxUvbDrZD/AagDma4FumWoQ5zfPHpv3Hhaa
OY6rLqnE8wiq7gsLVycH3elt3IWQa5kzw+RZcUS9Kqa1K094cyCaIZuBEuO0
8nodFsbYsciaMdvbVc2a++Z+1a8IzM2FKC1hNP9UMMjm+5NSYv9jO0faH5/E
cM/0OA/yeUEj6HKVtwWFgolxpk7PODsbqd9qDQ9yRRwjP4OyAtEvT3nAsa0Q
ql64LVDY+Pit4zocrfL8x4yebjDCFZPmD9P/QhiRbIyxk7R8/FieSWxoKIDF
jeCnwNcBOfTt+42W2lKHRwWGXejn2j6LosD3CHpqGLZEf1GQyZRKlSbx3KoU
TpiE/5KPxtlNiCvmAXSgSnGr2voScbKlZerb1qQSuaOsmqtgNZ0v6tx6xGgH
dQwKEHZ4S3HxXVq/+G29IIm+/zO//MhyCRrncKOzFDmwPgNUJoRUUnNx9ENX
Ec20jxUWYNJHyfF37+BCi9M8ENxv94EgBwhBtSlsHUXFLssqW4Nj5DlO5dcp
GiHVFV06s2SB9xoOVPiM5pJBO9OMdmZDu0f0i5w0dLOIOFa/5Btj9eS0Shd1
SC8f8zRX+Ejk+8yCIQPYRn+XltFxF5v9AyC/iTeUYFizUhYsrFaSyTudxYiL
VWW2PahGWUw9p4z9I9Og5T1eK4Z0uTpq/kXyl+ASE8m3QlflNqDObHtyUkpr
xLysFIZYAtUdMzn5POdaKngBBfa62T2NwnABKLTb9WVquwJLKIdNjPzSxXcH
7xNWoZIBZCZTMTZWxzepPrG0amTxV6eakjGRtpd//32OPnHTjjVz+VTOXH+z
MhLrbdKjMBVE2qZkbCHrzP6I+2Lgo3ut/ID0RCxJYL2CdWbIiYV9iFqkXcDo
rAwigB6ZutLuNKFKA5X/DXY/aKlA7XWHae9G889WFUiCnR0TL1B8l9JjtDAI
PYQWZ0bYRvzuP2JrvUY9C39/PedvWOYCKIikKNKgplilhKw5wapO74GoaPRO
J4CKBdZ26n3/jnL5Gh8a/jTL+HdFcDZsMcesP9Xiq/nPj/HxAU0IPr7rUAQ9
oCSuXnzCxYOxEMsK1UV8u7EZ6od8fpI0SpqdyGFK3pf3OsisOzmScpNllKku
KnO7SrpH4tqL2rZyyiyqBsYEXlIkEZhEtTXJh1baAsCvJ8vl4iSb4td/kPOM
PW/+yFgHT1K1SAQZt9bsSGCj5u9+FLpfE8cAfYxmvTAUpz/CKc7yK6V1Irh5
hhkKKMPgZV54iPgGKmyKCnJGsgj7c9+r90QPS9k+OShVqrQCzj/5kgUm1F0q
rdFy2SY0xKhiv5Yz+YGaKfbQUEqb3XXgmMvE8bJgCiHwwDHbMx73DVJnKh+m
u7DM3bu0JLUBEBieAV1MlFkz4w0RLnRxA/kc54xUD6JqeAQsFBSYO7Ri6Ymt
/NCsVO0Qoatz7FzcFm+f4vazkuiaOB/Uu5WAc+IuqmzF7mEw4v9wwU73Z/4t
BILT6/h1rPNXQctf62C6ZmOjrBUDWamhWnY+wPw4XXMi3tD9HidNvBuDQjxh
lWL93+rfCergqvnGpwudPoRyIZtuOfK8Vy0uO7O+HeF+bO7Wf6AHYYjFl18q
181AqzsoMMN5YU6srFfuRdjR4UEOVB3o7qXAcc1QZbZK02fRK1kFQ17vx6F0
D1rMgrQF1jHlQpVeCz7Am9fVQaJCfoCSzyLxa+1UbkedueuOK8Q8GNr6KqQk
0tdMnJQRfcoynE0iVytkhxz44rerjwNyXMkWqViRGhz34IPF9OWVvJJrv9hQ
d2cZYpSKc8L7N6W8Lc2ptdgpsY1F4g6KPBxBhUViQfJ3C+hX3wlEgHJJwPe9
cabTZrCRf+69EGLejBx2SghPoADy8/QAqU7OI8nQeQw78rzX9CbLKUhHt1pm
+x51vrkieNjHqeHTcMvta9OMwtrDKH4j7UafC0Nvp6ynrwVtxIbolpJiQKjP
3OAvuxOtqmEWqNOnpcMT6sbxGHSay2uxbiZ670iK6nkmqEK1bwO+hXnl3kLG
JdM36CBnKqtFwew5+zIWNffrBFdV/hYwX93sdudrLH4USKc+QNvhmQTv+3Dd
Mm65UaVz3toiyleL7evIhmKhAWfIzKIfvFurYqvDX76yr22bOMzmk1+ht06j
ZneqF/NWV6OkfvizJch66WXUax9toxhBtHgQx7qjTlb/tpUvzoxMoBw8dVQF
uGt8ctDB4KutMOBgzRxQUSSgVqRejLr/GXWZ/8CFqmmCdYQE/NFsvgvicNdz
RoS6TJu8HRNzdiCe4dQohq/lpLJKJ5G5zETj/8yvylpMR8roeasE1oP3wFzx
1CgSEB9CLyKVKbFhoaj8Wnb5lyAIpvdUt9qHJHlIFf2EmbOasfb0tsgB5AaC
05E7uBvn97UMA6mBpJK26s66iUY+5Z1vrrSEKBNY6QMozU+VNBcOdgWh+xKB
bfsPz+9Bg1FZRdCWsAbwrHsY+x2IX5vqLAhQZF6y0HLYawKDWwz92hSLOv5u
3BioHgaiPzmzkIOJMkuI/HGHdbgEy8ohq8sjVpR7Y6BHThOWiN2i8Gp+99iv
phHdZCTdADpzpOqWgG8gaczvIbOI2vrALA8r7N/JfdFlGhsN50OXPLPfUzIx
S+ucHNExGfsQbadAKtpZz8s16bqc5306rh7Kn3syhXS2EE/Ve081Oxc+3ra3
bfQZPpL31AfkNZqpzZFy5LX9A37MHQjW83YoACzGMKEq0i/55ktp+lT+PUo+
owQjSz0rzQWsbRIi92CHrkVUGxhwpDVKgYq0pjJweassglrihL9pXNExDSNs
qCp1MS8AA6W8LnaRJSNO9I5LPSehYZ+7QpE5zrbvRzyPdw/sx38C9qyLSU4K
FlaMA6x5Iw2CljAm4HpPBU3wdCGMxyaIIESzsDYU6G3W4XRdeOVEG8Qh3mQJ
bfXXWgGlZhTmGeR4lt1dlQi6MvTgtEIf+o2PKzqAbtuK74pm0HHrChz2zWYL
HCwTDi9kt+qvS2pLrrw8pzIFtaaRXJ/4AChxHXYHGEWLB+fNmhEKLZDdcMJi
u7GeeEgLD8NN5rOmnHJO9QO1YWY8b2VyHYBZi6gAu04Ynlb8/whry0gVp2Vv
UVX8ha4I9cNY7m83b5h7yMYHQMgQq6FffNw75/8d5G4TKzBdRwj2rJJBG+Z7
J4ktSkz/T6Zia6WC4H8HYZt8gzIxIsMHV2t5dQCpnVcrNweUjG3BNCwgNgyW
f/zFs4JcVnA1W5wSJGh1n3tRp72lk1+6uXM5tovV2iYr9WFzdXpXHKPfmIsb
wTgIx8iSusm2aB92PiTD0bJm1GpIMIK1cx5MsAUIPc6W7teLzDwTEPgmZ/Rr
r4XXdb4x684XnbCxkFKNcpFFTVQX2HOZmwhEBkKlopUTX7hvz4rKmlBvdc7z
fHKxOA2puOOF2MEAaU+qRxV2weVwiYYJ0XBpt8zMHjtkDzZ40360qU5V2Tnb
8xnMwVF1zTn3hB6CAohtWnJN/pHOEnWTIpF54ZbZNT47oQnonF+IVTnWvsB4
eaFuqr8J9Swna/lN6tmRBqGULgtSg/SEWL+G5teDwthIHrr2oHh7AV7DIQat
JHNMFm3CJL1YmAN25mNTCSvcy8LDI5C//wzUj6XEW9mLc+ut4O3IYwsPfUsp
827EbX6L89XrjVqSO2N2bOeAjKUkPcPVUZj7/g8XQ6cHIVavL62wfWJmokdT
TqwNWJWx4NT4F+4bwKxPLwj9OIYbSfYPtHpRJfj0NQ9YJ14FzyS84jcI1oJj
ue2mzTjv6a3zw2FAI/wR6gX6YGimtdZpsg84SEUssIQZ5hjxJ8o1RuCEWitl
u6xsmzyzxucXsnwif0xVlDUDW54F+tW1QZsYBrMrFukNArk8JUcTeYiS9jIU
+fWD3SbsA3z4etaPAtV1bQE/emAVga0r/pZ0K3eX/eAGnOFSrMvv6T9xsMdR
oPlgSWpEUoIXC7Cke6TNWF15nYn33vktr0vgWb+CADKZiu/xwwUTWnEaHjf8
wTd9JDn2j4G080Depo9ewZyFGJw+i2ZJDZm8REK2OeAH0L+7jWsmmozWvWyS
P8QQfBdiObH15inrTCgG4I9Xh6bh9TyTT9wPXt9EVBmeg+75MadDh4gIX8No
jwOsNHYkJNKdKtvwIEQ7BGqUj0yeE9iWdLcCG5ogvwTSDwgYYp/vxVv+Imfr
FEJjCzWWGI/yap9pYVUIQ788PCechwVybGCxg0gCNeLbVU1yjKReWxeb3oRB
/72ayvn8at3RKCuuoS1aNebcOquZf/fe6H/DjGdQjDNOvMER4/Td5C0UUdPL
YYkWJaByx91zwenAuIIlhUpDh9EAx5lGzd/95GHcSnWP0FKJKeWy9T7nimMt
V9ZNWxJJ2jOW3eWqyDdQR2CVaYvkLAbH/23zHWmxeLDpeP0pOpffNkenaT3R
obR87yPutesDdTBMwqN9dgg+FJkfCecuiQ3MJ3+g6PlJCwIeKK5vrOfKGnk5
KLi8SQhmtOk6KF7sCLkOn7dnpYzxOVVNTNaO5CvQSJf5K4BbTYulddDIK/Tm
BPbLXtR+krvVh6cPy++qIkoGyVohqL6du2OnIli6JsmrOk7MS3I/gSh/ANLD
wUg3yBirqYkobo1n76I/K7n6wTbmtvE5Ss8J/g+B0edtq5XYG8hdC1om9Et4
ESRfWFM7BE1x2q+5gQWdrB/6oF2o/p9ob2m1BG7ZpHymezKT6byMZxLxu/Gk
9PK80YTonGhfO5DU91HKd5j74fnxJtIhojA8q4Yy9stTV/Y4yNGWw913Kojk
ydc5S2MADZ11M6becG/crxWRR9HYSy+SMFY3oLyZ2dw8bE2zU7/Ll3mX4S13
G6BUqrT8orWwN5ISgpFzLIrMOlUBaedeuEqTa8/YYYUz/umd9QFvZGOYnsbV
DtGODmoFxAzZsz+tiyelXIRa02ySQd9yZvhHRBN7/WauAX/jJVHONzkSVNDy
ZI4ENh5/6FMdWNDywfFv9OuLL5zoGlPMhad3cYzvvU3yoGH8ml3Z5KGQ2R1v
AxcEI0W9w+JQvD3Su0JAKPHksn2I4E1kCcGGmmhDtS5WqOjvUiZoNQBaV8KG
90bhST0yj7l8DKcvAOm+m+Ectv4n4YP3UO+bITFgMK0nl1j1M0OYsDzC3PPC
MBFJjMZ/jbXjtlyYxBkoWihvVVZQZr4h96Tz0JP3IjdDJDz5VceRLG1TKc9h
27TmfXrIf7SsEdlObFe3JZ2WkRKbO2NwuHq0baMyltYiKMpQaPtqpe9sdeqX
W3FFqQoWwgDc8RTtsLp8ZLDJKafCKHE2SPuapU4GDfJujt6yjW3xXUYexrQd
D/30L8UuqCZ0XlsgX5z8e/iXMDKWQ4cc3p8xZ5uOrKwON4+7Cb90ZxA0Ws19
uJzzoSm5Bz45+vnH4zxEiyR+Cueln1fT7n9GWQ8Hw10tCYnUblUuFUI6K8Nm
xs1bW0BF4EFvRPMK2WOOnrjDM/GHmB8Z3Dx5iDfYFah73hspybJ/aMoflxRz
famPgssZePzTYLQyrhppItxC5CsSqLgPTLW5aUcV/JVZSXeWBdjrYCHtxdYt
FOAtJCN+VFBDCCamzHdKMkMkZqCmq+dYciX4THOujyBPK87gBYmKN/SL9BjQ
2pVvhMeGuGff2XlXn5HJ507aQvJlrdPe9pG053TVRHQQYns33Zu9lcodBcvX
Z3OP9tubXNigngEo8DBQXK0/yC5CmFjYHyqZVxRLGW2jRr6rzo4jf+UeWz6i
FW5r5jlFrrdOzWRHxfIKLv1yvjcfaTVccxEmgprIPJ+c5ho12f1OjaV250Up
JDGfKOrHNh6wpsTGKE2Yb6hP0MTXn8BumOxnDPyCgHOlXrcj23qx/anu2PiE
sq6temgMxQmINdTvvuP/+1zYTwGn2qQ4LsbpVqiWucZ7nnKMiBYELAg9pgTo
1t3Q7Mjb6VrfaC5I+mE3MNvtm7ZP2Qo4ezMU+xIs8+7HWKWwejM8ODQ5waom
JHeQSDH6KbIM1fU9+A6N6HWGUtyVJGH6L2JMrSoV+g2AJ6RfIqyO8CH7Ried
yC5ljF9jmG2ZVjqFrwzL+wlOMFh0O5g6x/X7ZWlSogs9Wa13s2uwRDvxtTBY
1V8t+KN0xRu/x4fGWxay8o6x7l3E2pC+DH03ZE1gZBqomRc5tiXBGkHvThpc
D6Tdvv8iAPBu+LyClEK9C2xKV8F6aMRYXj2QUipe6QZERk1hDts75EygF1Jr
WQCCC8YqeQQ9KC4H2J0US9iqecDSyiduPhMyRjzsKJ7gmH/Di6WmvrJI61y0
ii5PwHKac5eEQ7n/ROAba3s9rooB9xC7rdXlgoEf6I3nbOHHezONk+N7nDK5
dxIXZAxc8T8w7PGD2dIEhi+Y2Ry+gM0iccnJS/spVmCT1zhLE0+sTs2uegKw
qjAjnnMdgVJLUg9nHaf25SruHwQbfKtqzF6Bd1L53IW1D0/S7LpKHA6Aq4pG
CTe6s46eFJ2FgH3zXCBIXaoVG58y0uWJM2pTP6xeboaoOkDgLBcbVP3179lp
+/zgrb2B/0p7uj1wk5ZDnPlKVIFA9DxQ3iWhmoDZjEbRUWwJkzpIYSgyThVx
NBhlusgRpQKsEkHEsprbkssGWI4VyovRE+qql8yVFL+kEvik9HXPEzmPkpiR
5Rt+Nay/TRTLiwL/4vOWTzPLrMhV6UZYFLz21d8WXsl5bxrMINjEIkldUPwc
tSImq5Wshqk6n9ycMBLbhkOPUCQNLDnVysUgjWfOL3aQh0Nen0b59C5T588V
2KxxKgoVeHqfNBiulUVag8lMgecpeylaiMP9VRiV9B33uJh/DpUW9PjgAAUa
kKmEwA//anfuj6wx8h9IJgXQBCBLeDiHSMUSd4MEUUJOrCpSmj0Mx24DTYaw
9eGDYd14Gfs11TxGaJqvBN0GbF4918xwy0aDhOBxP2e7XkoX52r7ljthTw1d
p/M2r8Qj/Yy/SLgIHA+Zq6YdxjivqHPcwZnoylN0nSD2mI1M6iN1M3xeZo2w
A/7tzBc8dBbc0OJG2+7h3BOzZS3Pi9gW3d+5p/7tG5In+hIFzWoMp8KJvjs0
w8gN5olcsP+sfMkVPlZDGi7aiFkHHG0A6xtcpFkLTAaCbaYDsBFrXglL6K9H
2FqEYHHTasFMjhHzIStp23md4kxjYmt8PgSxTQPI+JPNIqNHZiXMJdxTSEae
Amfx7iYSoer8VclQ+6BUYqDizLoMSB7b8gp+2NQIQLC2UAE1qEtUrOE8HJtm
pflJIgV124xkiHbVLla9W6KQ8TL+ETZe7VXWUD7tl5T0TJ24ahVtUpRmw8TU
UkgS/zzZI6XLAwOxRZ9jUBtB04Tux3cMcUGBlvorxyhp+FtUTgK5wU/X12jU
AsseNBMwrXbxeLQQNafJNf4pcoWBVnf55m+feUBE/pNaNlo3gJ4L4aI4thW4
Y8pw32J8o4Ds7kqfOtsQZWQiW5EVTCi6xuXCWVLm8/xE4P9ZNkUsp0aAvuRt
//oaEInM4/3WLHkVwA/ylKeqA3lpw2CkVBc/mMZG2oXjj38G9pIPzu35BruP
6DwJVkHvF/2qCF2NlEJvhfTnPS4fUKODdtyG7aoXZ+sjEwifZ+1oYokrRHI7
yzBfw4abPxaQP+0gKbK0+63/oqkzGjnuEV+fmmB7HcVJr4M7r9POJ/5AijcC
iOV3TiT/cm58VWJ6NRb+kYwpwWYoxnASUEKOMEttWz448vfOiIL3vYhP+hZu
a1ZVhhlEIxCf2Ak3efpgy9J2xgdoN6v+USGmP0qT4lTadWRBBJv90pT8ykBs
sSpx2xUxRjSh5fs4wp3Kyrz0YF2n5uJcph2B6RRUbohr9NgXHpYE8SijT59U
pZPvu7mw4EqQLaEPCn008IxU+0/LkoU/nHAUJPs8oJVuR6eNYR4QoDDU7vLr
CCzeNjFJpy8jHiAqasYgLvHKvzUwQROTDOZlqzxyE2XLHNOsW/DHuhoH5LN/
8VNheIEn0kSd5v8fB3pASqA53y9rc/fslj5u9isTxe09u07/cN0XjC98R32P
PFE41HkfUPUpyTCgR3lYAh/oWIf6Fn9qSCIwMAVUKDBhe/XtcMyKh1khSdBo
hqZqvormkDe0BVw5C/OMqmlBUeEkHFwpnxspmNYFR5YegcdGR9ANo6VPbms2
IlCRHRdpLw0NM7/LEJWu46hzot+SzHgVweYRaTt3vZf1HNH396erEAcmFE9a
JXO6hegPqc1GVyvNeZ/Ua23F8qBHsRTZF76FONnJnE2wSdfv682EExi4wndM
NKgMHEPEC8OfApOD7soVCMs3HMTxXm8ETgP3wpnjgOlWhVm5m8Z7uidUVgl1
xBupxJrR7twQeac0h8jEj5NgOazjL3k7i4WHD6EXaNbxwgHJfjn03sD60pDJ
qhBmxTNwSunaYkmBpcWkrraGu/gWzlYHmtJhty0+OcHZprz4RVX03xul/G9q
Qx0wmNLc3RnC5PKA/7Wms1SEnDxdg8NjcfWEKJLlA4uniJESFyy7YpoiWDkN
sznh05SROQKO9G/P96QA6igVGzGWKLKWS0l8AlT5LMZIDiNuwZ00J3buUyyB
yf+AuLyRNHzqOkeaxBGezrGilIsudfXYsq9GfD1IWghx+UOn5otApcL+7JRI
yI+Fy26y3qy4u5JwV3hXLIR6u2K/K8qnIW88hYGik+hTT1HjEohPpLUE+nrR
b3aGF+jHTm3u0gmwCPSvBtYmazCdROkLoluycEygwubksha//mRvnNIqfMw6
5XmCLVelcKoEljBNFcJ56EkR//EgolfJQP18WUyioNo0rO3fUw4f7xA5srqa
F2Z4DnTViYLyw9FKxhyRCC3DPVATSYgmjLgKYFSnE14UIT0HEGncQRwUG+c+
bDPIXDhPVNAIL6gyBuX5BI9cLYy11MTRTev3PmPCLRY4Zyv6KSN1pwxk7O5A
PseUENpuEVVlUQW7NiYBT/hy4qkKpJzGTSqlcdeQfkXuycD/6WD65Hnab+qi
gamB4XjrCV+QMEKUVyG5GYrEYksWii1j5Vh7/foaCLV7Kb95udUYQwoXh2bp
G/QyIw950xBa5KSZbCwjmr2K78liB6XUHeAM5nwkmU3lCsLlEkyy5vWI645F
/Ji13BLYvtGMiUKeM2eXWaWoBNOU4uizJ+9+M7uZWS+mCUS6plJXByI5FnCy
DX0w7CQIyhXgVy2bKnDXSH17ImD4HeXJ0pcAWX6Xjnq8iNnK/tUDYEPCNefI
f309ZMTy5+EZUOJsqQvBLAhUP2j2/82hR8nNFuX511PWKqCBllpqIXalJvp7
soguicxOevo2SIH5wenM+5o7AXFH4pyZ24oXuzHOaQTv4fn4K1xbyvk/GYUa
2llYHykBvwCLhvwbzZyadBf+J31CJU90UOjhc4lWWhZDuJe7pqiFBaeRM1I2
kGNXbKmxAPyLibWev8CMR+NoQarDy0uydq43MPcx4FrDzA8+8QOeYZpNmbPU
7uzz2mLAxvzOXJyElENcWCpnaIBK10mizLEwyImp0L1Gc8yov6Kvuz+mD/GZ
SW/ApNF7CQJpbNeZp9+SH/LVM77+y49Ps7e2/YUwdPX9evdrg+llxZp+jSSZ
CCCw+sEi4herLQdkz3wC0xeruwNdTBcVN0EyFwDHkdncwOPe51eQeJmzK6sQ
UsvdSk8NaCII3DyawJxu5E9pU65WM2IKkzifcM955t5c08YFBDztAtc2/0Jp
Ejf6zNn+pvy7T/qO1p2FMKZ+kaWRXywBe/9pYMdYsYiAlnQMc4DD//561H+I
lEpEJVSCtsE1e/U9eqrfkO0Hl0NSF0Nz4pw2qR+B4v38fhnk5XGEV1//YlED
7fKrS84XvFtvBCMTeXSsOUTJQ31Q4Jytorb4YAtfn9ZHCQ0xW7V8x13BhdLW
aFNWQWFsFDuMpc0qSyrwgej7I0LQMM4ICDj2f69EfD0N54zSpeI41Vg60WS8
788N+QPn03VA9QbblODIa5U4nE+7p516CSaYH0qgG3q92pW6rn8fyv6l8wJa
XDVonL2HNenuOS0NIIXvvmMlkktKP5TzP6RA3huIIBWwTZ6wfwHo6LpsT0/j
Fk6iGYMqXApOijtpd56D5/VmYn5w9zqbBAZpV1kWTgloGY2Sncj5SmgpNdaV
q55Ah7Sy5eCxAcvPAADOKTMRoCz2rlPuEza3wYcsaBMudDCiQqYzXNoHZG8K
/vdIZtyjVfTVnfL56X21NgMkVK/prFnqV4RsBo2q9YLXXZsilH53AMDRWzwN
/NfUA5UzXigXnk/U9Y8GgtUpUu5iDmJUJTEG8eq17s6i8YtXDeX/dCiN6hwT
SDZjgWygPxytY6+chiMqi7AGlZou79II93e1aHs0e0++GzqWK1wyBSXgVPsG
QI65gt8eB3bifOgcFoh51uU7e10IhDiYcsAO5VOZCskkGi7YIN5rmX67/+YP
am8OoP92N7AI/aBjMFBZKlkDq2U9lnYRcrA3BYn8IaNUW6bBnsMHTTW5h7qA
gufsdEsrvZVXSF1fyY7JY+SDsvPWFrAkBY6JQBHzw+gr2vF2RyzKVkXvHEGA
mGi/E3MlEA7pwmr48cc8KBSGOXBNnpe9FxxfC3S0FqAgAQ+pLcN9k1uVwWhK
RpSSgU4zGCfnTFPMN4p2DVe8T1fJrkvz1vGRwhcP0vjqwjZzOMU1c31r3JlO
cKQ3asNYL//d67HFkTq6I5wwVJSyg/y+PuM+nxsTY0/89maVuyaw1sZd9XUB
iFj9jtihCAg/Al2NVOZp+JxVSqkzrFM20J1tqjTbJ9vGsG3xU9bJgSVVe7M9
Kzf6aP67O00+z1ydRYivqMD1P7kWI8xpG3gOEIvrNLiyaKEeIvHzxh7VKBlh
mTB2QfcnO4DJs88nPeJQu/kZNbUSZmMw8xO81c4g7EK2j6YnA8UKhPL6RhIw
/H5aXNauubkbVy+HnMXk3UtiYH0tUKNAO+R78Q/Vuw39kqj6r7IVPsj1pYkW
RiZoEHXrUEzMQn1JJQ7tWzbws0XMmTwO+pQGp8Ui05TanqJURxAgxzsaQ6Ne
7gcAuLhk0LuJSNLSUoWYFnTtC7LQ5+m48G8vaJ93fiwoH3qAmwmBSoClwB5t
XP+3Q9//nTZn6iSl8Zzs8Ma2oiWoubYetRpBvAOEjUatCNprXrWERubi38/l
bT5AJxspufVFdaDchn7lUjkrpHGb+jy+DpVyUw/roMhwHcj1WGzXb5HpME0d
J3JIJ9zsMBHmpMT28qz3gzXwkZCWP5b/IK03vwF/b/OaXt/Qw9GWSzzqU897
HHEznMP+4W9nm3ihvVeoYmzeHebjjAnam4l+spSAMZNseOoeWX+TqlePrKbv
kVuoWyVsqDFUXYcI94eJM3zzfrwbshqMmF59iOingBRXUjip9PPTz9nKNLlG
5PDeMNmq4FsYtXDvrdFhh/B0ch1+UNNnU+81SyISAbNCtN+5OigpE834XPDU
It0rW3cseuPDu4tvgMyK/N5EZzKBAg1hPSbElZfaZherc41TYA0cf4BizVop
UttIUTC6WsK8N3mS8FNgNRN3OdxIGQcgsg7MtQ10Lj10hhLSOEdrpsi4lw6s
1t2ExlCZmyQSTgiwI1Gu2sSujsc/KNR/bB+KLgpyhEUEs0kdGXbAJJv8B7QI
a9gHI5UJ52oUUuvmoTkpUnGZ7ZcTHKxtzn9GiR8932Kw17/k8G2/vlkUDQz9
e9h84ueTE69l6RXel9jBFl3ije76/IwbYDftvZItEv22JJ9Kf16uDKcyQL45
SkUKfCgTYwDj8SeE/WsIMNOhfFYi7dmrgyt9RluEWuBUo9dZcZxm/8FgYUed
bNlhqDg8kElPZDjGl8I+wWLG+JMuKzIuhwGiLI3vOM8gU1G1/9BoQIOhZj2K
tdtsnG+sDxWY6WT3zMumF2uPiACyhdr3TRObAvF3Pu/mAm0ZpAoDiYf9pzt8
BpZ42uj17eN9FP+AN8U3AmNa/RSFw74tWEWZkZCUoo61G9zflh7stZHTK+TR
61CjFkcFR87axciZieqc56HsM9NPM18rn2m6hLKRvjb6llBRCoJMF6jE5Hd+
4j+bv5qS0omM3yNhp/QXun2JRKJGU3vKkMyYIWtQaGTfM7O0ottmqoGyRnVH
1mXNQ6CYS7bpFvu39rJ/YhTxW1laVBrF2lsT16jggo2py3KMpUZT7i7K0WfR
Qn0Av63xwcQjaT8aaOsBZ5Vcaq3H+hGB0ID/5mfoGFhEtoMESIVPhsrHK3lP
nrxVYnv3+qVnixeyte3r57PHNwB9dClEpJ2emE/eUeyATuBKWo61ekjOGUfo
l1uxZlstXVDqzHLusP6euuPFNG1fqmHM0DpQNylTl+h8Am+nmIBTS+7L6yXx
MTcXY7feo55bpxF4MUdZIzwiq02ueNJt6aZOBW3nkv+SMYEPVn28htQHie/T
ddczmKbKNVlha4/Lv5Bmcpik4k6KbAbrbj8YMfav90CpIBR5p86ZryaSqsS3
C7IF4HsHDnWfoKO6Wkwd4t691Bu0BMxhdTxS6+t+hcgUkDT3mtkWdGDHtVZs
P3oJKr+DYl2c/skpN4bPndjrLz4egBJfoyFLsbPptptgkRNu2Ey2ZOqd2h1i
NaP3jpsDubJTjS73tnojDJFYCY+haWTjCuT7o5cREoiMSDA4RTTfMGXSUpxJ
JzIQqxBACd3POvoNL28DHF/BAwUWEhjID3so750N95wj31y/xpf4mhpgoIMg
13Kjl+WSXrmb8IVnG3IWh2dXCXpIgyipnSIezPgjkX9i9GQsg6PeSRu7TRbm
DeBUutKtd0MT+8MK5gzYXpMbZ2iz3Jur44VWxrvj9ZnfJM2Ra23rKWJ+rRJX
noesGWAwPIjawXHPky8pyg3xxgltw0HOKH0Vu2uNuHXxbKVof1ZMhmMyt3IK
5HZSakPMT1t0cf/uo6NqQzsNi71QtvyHd6SR+/BNhugBw2ecyGx8pDFZJScQ
05iCk26vFjgDH7Mb8FAr7zUqdEd5KgUFtRCXRiJLxEbq9yzEgskncVhKSFCR
boxwdlv5VgseIOaOgLtpUvpHBipQhRN5DksJAp9Y5LuMvr2pg1D3R70uAS0f
iSASEHL/oDZ4y/EyrjX1ZugpgZDLsMYMkUUX0NEPDxbjrtLrWAeIwDOOz2Sj
KtVQAFDzszEYHB9nyK+jZfMRcLJHmzHxW180oeCpV0cVm/EKFWqQd1g7+q+U
msKURT7stq/0FdWmoq9usyUdVsIdRb3jOOq8k/upT4Ncqrszax0FbmwWtA7P
e5IEXTbLm0zBb+MCV4Z9GJwT142NIV6JbxV7bNBcSedy/d4LD27yYeOE7A8n
V9gv83EC+srtR0dE5ME08QkAgM+yJ5UCFUM4jCE/pfe55kf8d4pG4vxMe3Xm
1b/Eqe80c+Vy77Rf5RKUoh+zx8iGOjE7jArTYAqkZ2nJ8abop8tJfs3HUSER
8CTW4OlYYxq6eHaaWHO1DMNBPD5uEHUyoAwkAzk8CVxYvLVmZN4nh8JtVA99
/rJlp2WHVf9cddezhzJ37986RH/OuKplBMrchkLeDhYK8wyOuDQNw/s1wYil
BNXHVNEBchFe1IIpv8pdGPnGxA2Zm/os5bvuCcU9WFZ2pDDZVsONyWs+Dnah
yGDrIbxMtoTst6QOBSv1FSZtict8yOMmBxt0NzRZLVh6c551HfL902T85oBJ
ljjAmW8Xzm9y97u8s07qaY2FBkvVkHmT5Cd/Z7IkIHi9YupDKenX2s0YJQAn
DH6mMDlVioHTIJMaiV9mqUoyh4XTQLwskPjYlUjEGdthjibA4CxX3pBML7eZ
WS18k+6rhqy8qsD0dln1IUDCErntv5xQzxqh3W39EbTccZKcNJsMzYuI5ehM
ZWTc//MbVmzyKj6J7/oPGL+ChmTBywOrN757D51lyFxAiFg5YbgNqsj1Gtcb
ES7rYnxyCzhQNzLC8gZMp+ihyLQFdMQpLS8HwzxYpL2JZQK4r26zju+pidU7
z0iZ2KI700xRvilrZphC5rCKGsuEZTl+Ek1+lNy6w7q91X0PCleHttYs19L7
2qyRk4DjATCjBcDFITagFhYXX8PYw+NGVURvMljyppF7UBXCqbc9jmeQjGYr
QTut/ylAZ8/BVOOATtYQ7i0BueY7agUVtEhlS+kP7RYApp6P0YZD5RcwBVhK
dxhpk+QOXlDC4vQ64/ETRhJCibRnWqHmTCXaN0nMzTf51SOgvSdXEDyHvpeG
V3ALXuJ+trQHsveXRZlRn9ejYHGFPbCDJBvPEBgq7bLskZ5twlgVT0tmgUdU
26mnOU67VGpliIp0ICNmFCyC4lP/N/8xyW8dYy/mCT0zcTh7z/5K2GC8fKBJ
G0J07flN67A3BxnHCizX5IyEjzLKwApcdBdXevIrxSaoiGO9DaQGne9JYOGp
d/nvEMQ00N5tTZXTE3H0X81Bh3TV9CMu28vIOSr10/y0s7KMSNu8K/GOETAt
7kbVAV9PRNd4AP7v3dUCvX3AtwVKPrGNk3GqRCZexNTeT2CDkv24d5vbfwxS
40BLdTZ+ICctFONRE3Q1TJshvgPNCZqxqrr/57ibz+35XCh7xWfBdiFF05Xv
1/iq0yo2qmCLroZ5W9+KN40iLMug2JJ/gHpsFV3gyKiaqtyAF75HxPEETJRF
WnOlW55hU+OKcSFsD+QmHWaec3tGXrrVH29LO/4vDVRZn/Bhz6PDyq/kpEbx
b4fRjVdFnaT8tAylKGqoJIuL74iezhxVFLNkJnw/FImS2J3i2a8DGeBRdsRF
WhFe/FoOg0TjohlTfIRqf8uyv0FsetCR97lcYFEZCl/tRX2ydR5A0J4akBEe
ipHsaZ8ivLJR7swPHGLJbg0emKBUgLcCpAVEXIW21MZ0PufzSMw0KAU6Hekq
aGwmOcB8gBU78+GZ3M/jv+1lSajkztn04cfjPAFFsIj84DeAJWKGUwJowsxq
/p1d4yl1ztF70S5bcVKhTyrVd5+tDR7TfDguP3QxyBMe4OSgohH4fTs5El6T
IIAz/4fi3AldDP3yhVwbIYNrGK1g0ZhQuKShTmZL3DVLtbsIYtl31GHZQA0s
3oMtbMiu5EgKCBFpwRJFyP5lMQUykyN7DQpUnAf7UbVaz6PEwdHKy1CRpmaV
KlbZo56A9glw709s5vFCTcrjMXoBZmVet4tHuPSPiOgKM5kd78J4NBvCDFSy
kefmqLo4J7VKeogf9o63jiCqLzYRFzJNBo5TY+SGOdPTy++pHrAIdHK5yDCp
eIeuDSGQlCoRcJMu3JtNOdpL2Fpz4YCXbHGv/9WlcyRbhaanMiG6rR6PMkgw
OHjj7G8RVe4YppYikupS03ycIIe8tgkCISrHgeqLFJJwtEua9Qub1J/S3LKW
ZCFdwifZKI3HElHBsBDeSbMIobbCScYbJ/7w+zj3itFs2BNmE5+KcsZBMMdw
X4rX7I9gw6FzL0dRIgeWIXt5VmGSoBHM8tvy8MsFf07tsP1YCuO0GEErbPkT
MnLPjF3Oa4l1K1usaNKqiigcfKnLCpn+c8sHq25d9gB8ZdlvEdR/+XQH1gnp
q9bIaeSI7Z+LzQxdVPX4OKCKO6NS6I9N25hBAAtLM4vLv0lFGhyMgiJ2D67d
0TnE630U53ylhOa1ekBo6SojUfO/oCp7YE26Crj4kIOE6IOL2+rs4TcBf2xv
EJ0zThVeVqmmpAvmIQs8L9qrO167FQbs5LtimwHITQdVXMwm7mDAmeJ3hh71
GMLDElzQEWqbiAHju+M8Bnt32J7NKgMra7dnss3sLOCWMAQuCRzRCJZ9dWbd
WQ8H8o6xZHY6/YZot3Mo9C8J/Ae2iMfflLj+cUKvPYJJ0JWAKPGt0i3DxUXj
iLw4Q4ynZadtZaMTy3XTlqNAYQLTsrBfdqvy+ohTWi9SzmvPPRqub1j7r8dO
7sHkiOD3FbYU3S59V1HDnCpyOghuVdDdpYMYWYUO6kc5GWv8xSZ+6s+10yHH
PrGxjBAVLOaSjXph2fEQ0EYnY38wr5r/PuO7hpCaAxHJ4cQ46E12zrPuMsBm
yNLMBMVF01C8EEHce0hwm67XXlXR1PQSr4DFQdk3MLJBCxyf5m/CGXKwqljl
JKNdDuaVi2dIFS3DmSiIYO0QmGCeUC4K3oMNJyq2+EM6PG0Jfycg/ZOsf4RP
yBsrKol9B54axbyZcIwhQs3s/HdPUeNYJwJdHXuAK7fv9dEiCY4yJSAvC2gV
qtswEH+pGAVguya/8XdVkxgQ0JL7ZVuAdb1DQKgT66AiQd77VHO/gm2KQ0Z3
1Q2M8Tqg+nzGfkKlszle8RiqntpGt7FFiaW3WSJr1y7MDkeD1nUwcq8wvPPp
bn8zSskyZ7llTOGc6ezKCs1yrWRuaet2qNSkdfytAYzUqzfwypD6R0BbsXeh
OUJn9rhIEoLpRanroM/D3FrTINKq3yZUuqoj6+3nuMGbNp6HiinY8nVv6kTX
0QhZwUAnlIDHcoTbPRez+FCz7ArsLBegSwOQTNY0+eYjYw0oIvIdlm2SnJ6t
oNtWJoclqp5cTOYPvtJ5BRvmkdHuvu3IEciLpRrMJ/jt2hnSsUGykRdy6jBp
5iYEMaZYUOMOqtu7B3cGn1EOT2C9+WxLw5aeRpIjrE5PaaO5dfJuRG/qDLl0
5e0m/ESfnXStsnZfMsMFRnoT1rVDOU3N7C25pl1VT6kdzntzR2HEKa0STssW
6Ks+iROXC1lYBT7BRo/CcH1omfg7Go5oDMT8Tsgudc9Rngp6wwD+GeVFsMdr
sjf64Cxp3HOf95iLrbujsZx1PXvLUxWuD4Yfqh0gDohW0oWMy4hIZsoM20uQ
XiCbHnX7XhrGhTxmVvrD8wCs9YwUzJ7oTCgdWsGMDGyyvZXiIjtBtehUD39/
EWuwUbcS2P/Lq8djmjFOweI++J+2fkuHdYd//QLq7/vqcBgdUc7RUFBlFqIK
V8y3fu1PBz7kGhq9sAVYbfbklX5rTggwN/jwHPe+8dyakmD33ytw6YPpmaJH
MgStnmoz8mnzMQ+c2eY+CLGQe5ioVF+GUzXdlr4T3lDBrtkRVDct3C6kP0xS
OYfbn5XFQX0ZlDNWXcoz52qAdPzuBG9KOmW3XnkqiyaRIZMdWbbtvM6JVMKU
+K8DpDa68OfU3Hxj67Wne/IMe0rxtJExfup5UIRShvQekilIKMhDwnRMwc7k
MRbCSxatRFTA6YT4nffA/ho0360o/UFdpfXFrrrs+SfxrelLMEau0DHGuVds
SKYxFI1bnIn1TJSVWmQF2t2EopAGQlXBq5fEAI5X7MJwUX/1YBwuXczZwwMy
JaR6eYfmEFbUbirJnWiaLzUyZzqPDuyns7k3Oo++hhIwpJBHdvu1Lh9m34nE
T0rNf1uCbNX2HmwrgzZL+pF3gJ/UbJpcz8fzRgX/50KJUkJyzHaWm8gFYU67
AhzlG33IYbtenpjYZbkyz+Qp2ncQdq2ApNgla4hQiwg6ZgLzuPDzlR7hefYB
iwmAZlYgRuplF6WsEpCM6YfEd4BaWM2h8nehEGcc/GyD2uDmmSMM2VcUd1yA
uxo3sprV/yfdAq30+dTj/jSpKVlOS98XVS/LP1Y1G88zu+vbcdkL83OD1YBm
1281UcQSSgfDHCClTuR8JOjllNoAgXpA1aBskEpHEQa2k007Wd7AaWW14dX0
KIK5bPsACb1zL8J7GE+30sVQP7TjFCC96a6Mytfk4PMRznf9nSCRk0fL7+5/
v2sC9YS3j2mrnsjlUlPtPEffLugUq6at33feNz2Cv1wqBfgrgFCIsaEUGKQh
Sl3Iaqjvj+h2F/1DfTPeY3W2PpQ12WkGgxvlqC61y4SWQC5gm4d4+KVCWL5W
j2qNdD6TjRB6ugbikcDLX5dA90qPixTZeXvZ/Pa30We6aoFLXX0mZTVPm62I
mYCG0qevKZSRb28MKkdx+tlIlQBBZ0Zu/FbtdLqp2IFl00VA24BVMreyIv4x
NccxzMSqTG8g4wYegPZaj5mNQUorYDUbU8Ats542nxWTbxo5GbHisKY2wObu
tBTuOVwDB9iEyCqbzSGC11EY4h4erfpFke+ukzMssiSNtOjdutJ8zPf5MCaJ
O9LdbYP4eAWDzUsRpwy2w+b+0+hzsTMr2JLFVD6BZlf9jDbNXbqAecOn7+00
I2zmft5LIzPxyt6P7fb4SU09hGDHvpAsFlM4Me0X7Qa6ipDW44LxThBJ7Fn8
B7CEP9V4kiLFEsgMclfFvRdyHgzHYqcqmnVXSiLJ7HEQSUE2Ut4uxMS+vpzX
H9mzC5OeMB9IYHF4GuDILS0O5cqBmpzmq7syD+8w9XYGGmv6M9UEt9VQnJ+V
yWYCTq9VRfBbe/pIZKM3nEKgDirRr3z4W8pzqah7sC9l6jEZAz7BlThM9yPj
0F7sdQv/QQ5R+7C/PhefwD5zla0U8PUudXIzQlcTDG+ZdSGcVHYdNsis4O4u
wn/oGx9tWJURK1EDJQt8IoeWdbs2etDWwl/wbLRuqtXQGvVDABLLrFB2Wejs
s1kPIFy6xkQMZEBSMbsXe8QXBWW9KbbqJNt3dcQExhUAVjhJlhCsFQGB059L
hDgwiTFKy6c8b5+W98xcZMm8nJEJ7HgiXRskxDKBftf7ygMiGObm8iFqkFOd
sUGVRmvSxXtzZva4pNmG6x7c6huuoAxHXYTEEMe3X1FdAcF6Fu34+Pr44vk8
VttKXUkp/Hz/WSXwe7HGf7X88xXaruFtIDs0jmWAK6qghXUXCJA9+fBgLr+Y
gaDRuwfGaURtaqUcRwMWBTJOoLHbrXZjdgsd5GZpf3s3nfTKqUWbNd0DL6P4
KwswOK4e5wtCX7ziWkxlTyTXW7r6/8YRrje5j4XbSfx2lMY7nY38X6oxvtF2
nF8RoTD2hGSM5YSqG31FVMXzmxs51quLm/VmdL+2gMKO0QnF46lKbm1eg4r7
hTGnAddTSX1FzKEIHRlA2ymmEywLyUXTuLClaDyMucIDyQoyoi5mldnMypmC
ZESj7BsQPErThEVO+cjhjfE8CDsffyFHYCxnr13Z7b+tz0NOxTi77tF3O3G6
1CroJrgUODm73Sgj94NDqI9MzlTZxRy93E4hr5A1PJMI+lOVQbkFyI2Xk3On
zwLKWCAysvzojIBxyHKWmFMVurY0NUTsHqSmE8h67k/KtWyhDQLXPSXlPSGe
W7CdReYDLYwRo3SQYU56Hh0qXV1jbSXu/CF42TTHedosXBrZl+NAa0bzlUt3
fDyko4XuMNvORoLfSebggkClWS+HzTqYytQZicJePZoNQlNSYT5W5BGAqqvk
bfEocHwgmRcTuFo26P85Vjmzt5ByZ4StQ1OGwCF44AatTuNabUEktcHQnD4Q
zOuToQ36qZw9cOsfyuLK5GcBfQ/hbjwi4dAApEdFFPltXNY9J37YI5znvpNn
CGM/OlVQf9ZaF7U61gJWbuyfOjpPOLRWQCNws4ZHA7r5dUioexTEuRj11JuM
JqC3k8G2tKLpZ4A8keuBLW9TVFL4QtAwg1B23ATtf/s45xy0MyttXQxMYfXi
5JY8TvG5vUJosDic4X4fsxLjWHQQpmIEfgDP49cu/Fq6TODp+r5pUxLXTj5y
10uCH5AD3gW55tIS46Jicej6uK0CQI5WMpageM1mIMYtWNgJzRSMCnpCk1Zk
Sm+khfCKWK8msbObQFbd3PzLc/3ZV9gpygjkxA5mTrEbshsUb/p8x3Ol3YxF
JgBbIXCQfEeA4b5O2zSkN8Y3njNtGkW/C0leKNL/1B366xLwFds9eT9aOSwL
MeJihrekFksAWwNZ5f93/tZXWBmnqQ1xlHip6qIC4WqEPI6ehxkeh/3Z+6J4
+AZpqmNTLDD+GO0XmM5bTSfI6Mq81jA+Dly2k7wFuBH987qvfF0zEXCIWPF1
kC4N6WEJXPRLHTO5yKaD0QzOKlGlHsvDw0lI2rhPvj+QVBXpQMWE04wiQmMI
pY6+NVEPwv6q9ifRk+mi90VCOqR0TbPO3TiO+cKB51A5kEtSy5Pnl8BVO9xY
Iatipm6LVo1RJgPqjQk2OAEx8uAI+2q/r8qAT+EpWmXJU+GWs+pSpXStHTvK
qpaYzsy4uN0fHGVtyMOeAhRnVfrF8TkPoB/zixMMRQR1EnHBN+fxJRWF3rvB
if6VStL7II/J3Q6egVYuJOy8meezJSVVpI6AA99U7q9XnKNogNNajSvw3riM
yDbEy3k5uKvvh5V6BXF2M3T28c50cUk9e/FautlSqm5jO+YOZoSFKXDS70co
y3dqj3BasWvmlXKmZSrGVVo0wYma2w1Obga45xWxh8wF355jiZLOsgEiJYaI
vnwpVbxzsl/6r/lFindX0DS7Zj1qPpkYhUJHEcWEqp7cTA0uxe0oUkoSLgdE
O77M70qD2f/U9+Gk3EyeEc+w0iIuKAzFHgHnCGPW8hK/YXi2V1PBw6YyUr1E
C4JlDygINqvZvkQp7T2KeaxugO7CYBPEfJrp/tCwIhhoHJw2Z9hFVd//OavM
AwItTRAE6FO1TfF+F+M9SyYxtDwZLXY2oNIzihmVPsVk0uK1QjcATnouXDss
HVpCXJ+vrmGWduJJ2EKbGqkZ275u0ox05SPQQ3gK+qYP8xIceGCoIyCcob3n
TJq3PzaApDCv0PJrzCuHdilLFXNyZ2uiioM3g88is80qn+mgL+aGi2zqttUX
pwcI8sZDzKynzVpu9LprwZQuQPMDl5J7xZcAur/cUyLGgj5T343lUuRM60f2
sjV5p9RzSTeedXNpDYS53pmSwaSL7WICtZ1UUsgJEFPJ4PAp47DOr1lBXo2Q
liVl9bZVPmYhuJzyYQGeSeDFVz42Z1E83MZXrc57rEKMGQjifVFiLL99k+G0
U1vaNQ+8iZYpWvaxYBaGf3RI7W08cIXPcroDBPEgnpepYyOW2q5U7upVv7WN
CdkUssxijkmnYJjRPHYjyKx8wjFjM008Mfdm2g6XvY/V3zGZK0YLhvtqnxJ6
LNzwct9OOdNSIT5oZqN/DlU+Jd1UkD+4PAfSuJoHpe7GTC20k6tIX/r42GXv
NjHDYJSluA6YMm/fMBHNeZNlS65IGEsSJuH2Y0y3KhfI46Ns1dV5HkNH0ftC
jqn53mxWeYzgl3+MAI5NKxYn/2z2QALyPFaAzgxCwF0PG94ZEz67SmiNCGYw
Da+5SeTjK2xAxtOfij6qgrpifKzQZQnYc4HMqUVZqKjDCAPjHEuYy3ymdc61
sQ/Ku9fFmGKIo9nqrNcQmFHuT/Wh9htBCpl1xJvc8QT7icJdecPo3Yao+9PS
rHPCgsizTgTeH9iQ3zYYpZfvNjhIubt3538WcRjczFy9dz2f/t42uxUY7l9i
XRVL3kIGM9HBrsWpcvXckS0h5TVOqSX6Gc7sHyvb2D4DibVvcYuTGO1S/VMT
B+2dDNtHwhKnc+dMQz23omeJgF1LCJPVf5KA17fb1lE22I6bj5g4jbkr9HtY
AjcVqYhJnE6DKAZMYGj3y2htaPXPnC7eZW6LfR8UKK/cxb/i/kykntt+MGB+
MEZodGi5s7TBxqeY2XdUwJ8Xlvjh0m4Zd43Lz0ighzVmFrtGJt/eG6MmO1u4
i1a8P1weIaJFGuMBnduy3jtOLlmDiMywyAuz0J4OU41KRQzGcCqx/PzyTZd+
oiqJuYUxTSvNNiCAqjiqcHp+v5uFzAk9EQLNPsw/nFEPX9z+SGZSTtGO8pDp
dtXaiudjy8RH3k9PpkCQICn2SAiUfLLMtHzzYcB0re4dAzuA3eTkatUZZV81
aQQW724SCIl7EDjk1cInodhpUSn5LLdFMsN+LFpo4GBY2B7jeNESR43an3CH
hFKiuSbcMqDPo8lbA6ytWpd43ryX21P/izAA2N2Zo25RdH2zXgz7kORLQdwf
4RH0a559w5lcdJwRTivh9klTeV5CuNfT70pqE7gcwGFmXT0EWZzkscasFLQC
SVqYUIK2eFSfWE1OYWWkJFRZOF557ZpmMmTvA13e+pW/hD+dn8GIcUORVbEC
Yww2o+1Re2w/uw84fAG6U76NXB8pZezb6TQM2q69UnZ9MvW2c8NbH4g8QDXV
YCQANsRAed9Ff7NTW3BTx3jUGEM1nCl3Tu088vgWAJkvp30TmtAJ5hSjSGqe
6IKaSOaQTUQRK5Hn/zTi5Ockjrk599j40+xE/KO58Hdo/ksCe9zfE/jsJhN6
F3ifzT+pnfilavraGGttQON1pWlPgAEVxnKh7f/a4kx7MnQL0VTA/o085UYM
8DVLEMYMj4maATvYqdePpXQhcCTHJkf2I7TVX3kHw2JaeqSns2Mrlq1N+6le
hre1xgGOSUzKbssuigVLdqksRJ7PAwLeXaL4WHNb+CTKspt/Oo+YxKzUxJSB
hnuRPap+YOJyskyaj0LwAF98xB1qm9JNEwBNe69pRxwwmgoMegYh3DXupgdR
7KoxDP5g9qJG6qlCAoX7f9JZZN+fdbgXBuKI8NbiqhHrls0DWnS3M/tvCC3K
d5/9yuo8DgnxxC5EFMSaEbOhAYgAShW/EHetuqpPitUk0sq04PIYpHno5aR8
qORGvrYuArWuP2zCJAFOn4GpbRJrLQuQrGS2IdhKR/Y83oQ6zsz+ZM12+LHQ
W+VhGdPMBk21gHCIn/LdR3l5zZ5o8EvUxHHd0i/hFvmJkns2+bfD0BwjYPpw
GXPaeazDzUviHLYaf0o9EsL4r0kD0Falal1qRePnN6QSQV7wenHJg23oKwi8
jOBfh8M+KdY7I37XbqbTVE7KzKJN6vSlvoLC2oLW/lCLFGWBXnxtUyQqOal+
AzGjpB7jRHq51hQdc4OeAOQXseS0DkEGv3/t95da+015qOdntfT6YNpGkxv9
2Sd3gUZ4RNKJlhxlmwTdpr1B4InFvBJNU3LNxMHxwao8FbZwfmmqvCz0tp8T
EhBoyXLpU3SQOAQjNnzxVRtxd9P5EmvUhQuti+6gsPrFH1gDjA6/b6BD76FE
yLLVd63/7kI7R0vXjrs6fxoxdb330Swx/bixlNCDc888NpE4h7fXgt3DeQFq
TbkqZHmmBnV8iChC+wMmzGxNXq9gxH9DbZ3v357UN027u9Sg0KByL83yaBwp
wAxrpK/KTNLuxZl58myglXXCQftEe42ZvBOGDPZeQU/B/l5PmXJHmyCpWaFQ
XIOGif0EAamKRbqsD62xEmW/ilBgUC7f4i1s9OlFQn2VHNrJEl+1gf5Fi5DB
JQrFB1Yp/633wtSS2QK54z1iZXJwsJpTzBOmKqLIt5GC5t0aQsjKdneqCup2
nEeCOGrnesNSSRZWqrfYPKHxrgQ9Fc8Y1kMCU4sReL/wKXeFJPRYFw12qGYJ
Em4ieuiuYeGyM21jWr1nfoE8AOD/RpxH4MW9Pi6li5o5aR8txD6K99QZE4so
TieIs9tu9SZzYlZVqZ3pbzrIRlNeR8LPRsKN6SpGDvj59cABxAkncC7RYIX9
hr8WOT0daWAZk86oEt6WIaZ7sG+9P9jk+SN0Ms5MK9ZQ+iLlwcrpFwC7V7Y7
wa5hAKSn3JE+IimmJ75amreseIfw/DSRYh92LVRRsbEV/Bumsg4AcQw62MDt
qFTYGp1telb1u8QzDWMWhggicPIeVQXz4wu8GCCkAG5c313hEQlnKc0/l5Q6
A2EbEcmKKFSCx9r8p8UjLwBqflZfKrBsMIURKzHIcWuJN4Y8mc3ZJCmDUK9I
dP4Nwrvz7qfN3M50L649011orWrlWHumH5pMCx6OVkVODS5WKgXUXEfJhMPl
a+cVhjKe0FWSlFD+bUYlGheaML+9NsOyeFZC1Ckm1nIBwzypxj3Y47TnuRZF
7dqimDi95eqjqgyOgMPlVDdAiw9yG4SiJgdQed1BH6oHQ5t9IzxCpDUoLw8X
+lNo4VBHygClNsFu6Gbww31lp4MjbrNQZ2yMYxSq473iyosdBMYtMDaT961m
UZeq+spX+/GihM89CL0QQWkmEE9jUFC7kR49p8VAAVfX3K0xtgsDg7tawRl+
di6Rzwt4u6d6uocE04q7OdW1QW19mWagDGTIQffLHtAIv/uRNHT+aZ8DSUvn
znL5WgG2X4VPR0i+nCg8zG/ntdKeY3+tsoPkA5Rp9vlGVwijdTb4D8dAkFna
hh+W1bcvOZgab4Cg2SxWiNymteUE3fIksDOch9Z1j67ZAdb0fF/bmA2hgs0b
FHRKY06YrWbl5wRNUttFXIu1j6WVE6LBkTqLw8RmrcrDFYTEZeFbXPYV4Ym0
dsHxOs5ocoLySnbaPdJ9vSYU9DQ3+kNX8g5AaKf0oLgBxuYdurvCYs8MNlEb
8I7FMTwCoLxsr8zRzlDXz263wl6i7RoWd5Sj51aVUtOE3kqzrLuB8+bH91Ef
ifivIeDmZSYZh2IxBzgW0iv5brwnkiSmrseBBUa3UszMaO463DxWp+zWQyqi
+MgDHkfLiaHvJLrqw3b8sxVbYuNcGSwkCq6aMmFSQBt+0yhiPkF7GWPbJl86
XWEw7mvLWP6sduiuE+GgTFDCf8Ey/zgcvKUu8PJUmyMsVnhBMuaciqzfMLdE
9SU4Ob+aFCfMxCUfVTnzeGEDzN3ik2o0emzzsgmVuIYdbkYL5JU0icl/G8Sn
4pBqSjQdqykXvivlZLjdxPqGizoAhGZha6VgC7w7KIKJRR8UOwv8mjWK2d8z
4Lz7emOyHcn77N9rZJZrRdSQltn4STGa5kIaTFnvi1yhZDvycqrRP82aUgIr
DbMDzA+9yyKqzUJP+UycujDQgLY/oeOXrq/mJzm9bA5OsnrcxxWVyW7Djcit
6vb8CI+UKg/EQidm4yzITOtBVt6TxUQwuM2KO22EIHyrFOm3VekzMDFpwhGH
BfJ+Y2xYNo4uL2H784Li5xRui5Hdl7H1mEHRvq5JsQHLwd86edFBwIKbSyky
QdH6aLPhjmTl1ftl6XzrnY9Kuz96mIG7Clsm/zN1LisGkLF0qhlT299kylxL
DhL3p/36bcD+Ru9MtfAZbdl5bAoFefEmT5kEHR7gKWfwQlwGRBBZNZpoe2AK
rAaRlko1GXnSBcxUEgpMwuZIJN+gLnhFfJHFjBD118523Db69Lvna3WBT+K1
zT0iyHox+NDaGVim77jnzctL3M+H5/Hf1kvFO0+gMnJ/9iDkFkdVRDngHw0f
P1h2uiakl1C0JfMXKBfXq+QpQVqay6YbrnkRQk9HBbuVg2/kF7RoqlG58q/w
GbTvAHxLIPXGVNVRbDbhKCmlacZcONqtNWQZZQka+tDizhR90L+PFqKurD3d
gz73QCczzbpYrt8qMQVnlQ9hHKnJqklU3rhe3XzMQPywjHMVh4QBc5vDY+t5
cMWMmeGAgDbeoUKcO9KzH264mY+lwWfr5IMr8LnTJ/41JqFTJPVyoiVo2x5X
BE2XwKQ9+MYB9J4EdlD9uTBoBRDoQX1UqqSyXhYmAbPW9NDHJjDdESHHtH4x
hljX1l7BjOOq+fAwJkOW3Sqilg/5p2atYrIvnn5bBtf3Mr5mzY1bFax6qfYO
z13+E3q4YHsUWf0x+4IDvOPEyIYQ+kp4O8bbU7SsPrtwqxupJ1iS/jX5Q5OL
0anUgsyWjgJYoY3T2mxRWldP4xKAvWwC/Ifx1wUTG7HfQz4SZWYoCDKIcquu
EF4tDc+9pwpyBYsVoYcAMn5U3CE3k5Ltn/x5G7G0cFW+36MmWKbJ8//g44qZ
HCCMlJ7qQ2tafhoPQu4Pl8go9WrcibuEwZmRGGzsxuoD4R3S1C5Atzs1P/z3
zAVF9ntYKrtZKW34kisLnm5SsOpMcbpliYxmh9qy4IhAxYhQVAvO/t93VbWJ
qjRt5/wo953KxVJswfrSDlj0qFfswl8VqQYVEXMZIm12M7uxrTUMrKwrV6Ki
aDnqU+gXhq3Mle5INuSJr/6xnQ6MOKwZQ/xhVQbTA5q5xE2yDDGsDM9ZLoqH
ltKfzUWHTNop7DsagF6tHEYav6vBdxXw1YaWFcUGFJLLeEH/x+qdR0FTpjEZ
FyK2T0PJ94Qv5zSn+D2tRl8V7bJNJkIMCcEZ8nkD7X6bOtRVRvNQMsGdf7ct
uuQWZuAko9kCIfECocE+U7Z1u/xGDxeCibwCGbiBywfZnA/tqGOZtSlOo4S3
ioeJSQWjm+roLLncpf05I+X6wJCR2VBlu7vo0/7e32g8F8kSmodlnAa+cO02
1cIvs0Ru/Q8YR/1eEQRPaqZUp1gnhZHWQFXHIprZ78zfsA8VrjTywWzug6Zn
BtM31QWqPoRVm58854b/BeGqv9G22r2NcZQe3toRrJiEo4I/CjEPNHH50fdK
IdGcNrm/1ZZwJxxIe8m10AhE2NKDGxANWxHXP2iK+iO4KKHEqhpJSC/4pT9A
wFZmyh25D1ZiQvfHgc13eHA5ZKkEs4csN8dOqmaiq2i69eExr5Q8RdUzt7mt
gOKysZGlpKmq3gJODnQ33xBMIA7vHZsZuXe/3Ow9CirHQMfZR4U67YEF2puc
VBmZJOKNxsD30JWJYYH/qtaspkcbe+usNaCJenqLis39EzJiHmsn7apGwTgx
1qlYZNaePFECUKGUAMKuoSa57/O7tUlEgdsqWRikg/NZuwpVeMz8MJv2bcb3
t6KDOpcufR9HiwY8Lbce0nhmi2TtYUa+PUyxXRADkvOmHdeSjYguOFze4FSF
S2KbrwcyuffdYw+2LuXqDNsqGoYYu+Knt5jdzuAaDLbTMsSPtx//6RyJXAzZ
fF6U+YYd27Sa8PqpiyYDUt48xKVwjhczBibaKeYYWmeja7w9s7OTFC9pJLCN
blayUJx+qoN9YYkC7kIpnRDyHUYfR6PKGxb4pnDrp7IimuPjzoUIJNhBcZmZ
MS8INHCtRfQ0Gni+iVk/++yImbGtavda04h2/Erm/JsCh74y6KwcAmIWT0To
Hm8PbulHKC0tzMtQufODfWz+YlFpfrflA+xh+DOcE04cw0ZF9ZCvcY1jPAtP
ri4bKX/IALRgAiTPp1rAqaS6AZzu8VAulhhn+1ZXGc3SuMQSFmmJhZZGhf1p
mItss6GTrmalS5rSabYkhVTdvzMn1DsSid25zNpn3dOgteI5Y56S9hSPNaJd
kzCD3os8MCkx2+iE0PYtZZg8EhH+DKT8WLuUFfnfKKjMzRbRvsDW+Qaop+a5
Z9SvB0KgSreP02LEbgfiin/wMym5vDWqJ+XEVrd8kZKrC2CxwFgGFDrK24BV
zcQWAw80LimDyByDxsnJhRnood3mDdO4BWgTXQwUObQWDTaK4vijxqn7nJZ+
yN4faGyyXow+kYwaKG4yrELTHJepAriM9RQK32yxrSTSk5VxlA9T/v3UrBoa
3tjyv+ooMEtRugWl7dN2EajsEl1RhAfBm3Nr+FDSgO2nskPXd6na4R3HLSnv
YOB3W4K2k6KWTsbA2Q1QqJUtImnRQqVTHQdQNq4y3SnZ2pIdDPCE0QIjSzaq
5rwGTXFgaTdYuz/Z+DYWZSCyuisQeNl3dHaB2XO1mFSl4sI3neuxZh4ckv17
H6PoImkQzdpXE8TyiDpwNMoN9FSQj2PEvABilu+JvlbVozc9IRUBqvlaSQof
Kzkp+GEBX9vlO9EM/gW82V+El/SF78GVU/sIEr96K+d0M/kHkGTLPs/rY1bh
CSLPI25xQPPQUSk3ib8/pHW04DrGtazsEgoLbHxZZY7wx7oqk4CPofpYTXgZ
wiP08p/VcVMFPr7KPA6IKXsarQF6HahiDPakO04KWqf9cNn71VaG8R09DOlS
DDWMGJ5/zxqxz/J1HK3PDprbYOQLRoZy5hpFrs/Nq4Y+lEuWRkQNorEvrwQ8
Km/EIOOIMDhq3XEsxHpy2V1DuFoo5Hch0fV0I52EAKI6AJNyGn16F0458bGV
VvNW3kdCJT9gpUW2HpbvGwCUfBpWdNfnbKJ8fwGrw5WbE1Shp7kv+pHQelVf
Dae8O9KmlCKr7toDxcERzhPArAVbbAHRDr9z5DpTk67plQ/BHc6Z+qWJJ1g9
uDd2kMqPNYWQrD8D2W9Og/8vifNzsvmr7yPZbPWFTBI8x6ihKQTJcVp54MGS
aRfEGV8ogRRinWgPz2PK3wHngW91/QTNQVFxgU6voLR6OY0giUwH7Xn6bdWZ
Zu0tvdssqto3FmyI1PYb0TrvetgiQFjSgTotNrVsEALDNtecfuQldq3np6XV
z4X9crkfJI8TNLOjoPfMghOnWANhcrognhXKBhGOJ1UJFQOg7Fu7Bt9TWx1C
BRdP5yPrKYHxBwnMl/SE6HsN2a73Qw5dyQKV+zlOSdXavLo2QuVhngHEoMKH
Ekyro75lmE/j7RfzQlq2mOOAoCI+gjXOZQ2v/lzmxWWXPhGXKF2iiHtYGq9f
8YXMxM4xOcOZjvSob/p0ZMgoKPVdXVwPVK+LwXiq7QhMyK/Zb1Na6ob5CTH7
TVU+IIvoC3LEiJvFo3U8uPqFrhy8xiGLsws6P1QRIm8lvgHGgZGuJqwNij7W
nnXxztBpSGcuXbVOLQgjI/ZEjc8ymznCb/OoOQmTxrvjr1/ZkYATpEq5tx6u
dXEusCOyMXi7X/9YYPvJ2YwwaBDCqjr9+4hGxoAf8Tb2hLEYHaS8PNwYQRoU
1iq7yuDeavMsUIXiBGM4tJUvoBxAUIOwnWhw++5LuG790xKsl7ut3MEa5QvV
Nf0nGEFOaEVvJ1AXVt++Pz2jsBWchAmCpiiwIqs3RrtBUWuubbmM1Gwvf+zp
Hwkral0llxaG7aYUkSZ/9heIzEyBMjMAlo63jYwy3jmjdDz8vwK95jJz9lGP
QZ79GNxMnQBsv+49W123MDTsDFBy4Or8iNnJE9eEr8enB6f8J4stg0qVkMs6
gZhej1XJqLS/lLMyOXs2+F2jcPmZxbleWpa0xMUA077+Y+kM8LlqjbBlQWWt
Zswxs2IT/1abftNz53cecpOMy9UnZKpl/6Ve3uuG60w91aTAojj1xEnknUo2
NM0wKVTftjseK70YAQiMZG34GahM9Y9CJxMzBCZSgIZJXSUDht+mYn/bsGUN
TGU1dSDvK5v8L9M4K6k8XTYq02yh0maaD6Efl1qCCg38opAhQlhB/0tI5EI2
boG2ECTJnV3WtBWrS7Nj2tSC/iS+s/kgNcxeaxFDhLLHmtHYbTSyLAH0hLT/
Z0YY2qSMwS9GzJ6/79kz8aDDreW03cj2c6B84pn9ZRZ8rWS/pe3loXD2Z5PI
Nm0IPblTDZKh+kx5Fy8hHGbtPsTpkSlsys2sa1925LYYwehYiEMzsFJ5ZBjZ
/HqqZKE/0yZ2Kvx6q+pLn5eZALzNUuXtXXhOtMLOAsltiy8X//3C3O9nnH5s
Ulw0O+ZHYeEvWag1ulbxSnjKXOiOByackw0CSCgmKt9CafgW4T7KOpybH8zQ
pahYwOxVGo98/fnZqiu1CU/0UpP/JGl+X5dhqeE+QgSK3hmr9ujMCrLKdwPo
t5+MOGdGpBGUJE5um4gL81Xk2u/4WOaCvw0q3FBqTd65UjmDF+aZv98GlGPt
o2F37UvIrksKAxRShoScH0BE+etkvri9e0Izzd7ZnlqPj9O0hoF2hWG6MveL
yx9l1jMw25Mg10/RTAvGMuEP4mtTgst+oz23/o2P7yJlvGS/z4ApBYRHA0vq
wimlFvIsrfuBpaLocwqsLupNiwASz/umGGK8EQAmGJT/OR5zh92ZnzJ14Rbh
XVMPw3t6Ms0f9PoIdQZaqswYn7liva560vEBC85McV3Xq8Yv36AaKwaqHHSQ
x0BKlTW+f956CcdHVSg1383pz10FxefhyKsuSfhaJiingGi5beV5p9hoA3Jy
O1IvKqRDPjwDiwr33GUdyH+oxSPeASRvUuup/HVHg7ZNPJd68Qe0M0cDF0HA
JGbIxqPJH+3Q3BoniNK+v8tFkB+7GTHyDAnWfJj6aXCt64XYo4U9JcxEx+S3
TJyqHmh8Mdmfih4pycudswB9o00WMjaHI6uwbTAH8RRj7uf13zIBLlYzn/Zo
N9htdn/QiLJcr83XC9UaYtfn6ht/K57UWwlGjBPvsqciLAJqIjnnYybA0JMx
bqwqRSi/msr3XxzUsv4KTWTzfcVuC6kU4pUo23vNMpdKKT9J5dDmj35TlBjn
vJa3Cjmv9UKjQ2rAYTI9kRJETd/kBte2BIZrxZerKG5FzR1nA5Wr1+8ch9yP
b0HQpxExtvWmvh2Gvr7Btfc1jdEYalsAkmQE+bVWEVkefJa/t0zJJzfkGtPf
kdMIB/SrjYqMs2qFhkMwcl0VNM3b2kE/4/6udz30IYQalCoUOgFgKRs2T+PF
Q1jIGo0Uwf/wSvzOjY64PcNpmwpvrDSkCEW0yXtO1bgEVIRse23cPa0e/dVI
ra+KbkW4nGkVc5tKv6OuhmUVZO457rHMbvNMPzrWPoaiLTu00j9ieRyz5gCt
pxfT8iy/bgIams+nKU9uhodvx8TAPQyLAqiSJcGfibJTTrHqaDUyqIri+kwJ
OsZkgOGr4or5bJ6OoUJnaqH4THwSw5WOwHNek91WQE9q+wqMNy5bzTK8HL9q
4rvfQpos9848hJs6MnygGAawe0+Y10mlCeqbb6QGgb5vXBpX+ZwKMOzBcLez
QoZRVcxqCGnLmRqFEmoqjQvYBWSxiclA1dUiR48NTaNmvEef9MOxaz/FPQBC
RjEWXM54OY6gPHUBcZdnyQhlSAgmd2PDcTzK6gTTLMiqNR0pQNF6YW6P0JKB
Pd6I4US8FdZF9OZgd1bLir1fd7ceCixrWZHmHj08eGnZx+yBTTVbXjpgi8b7
N3V89ctwKDMYmKBw763LjIBlCIZseQbzydUQ3DOYeWpqYYhE8njZfJ3f8PNS
q0rRlazMSW5uksNdKlG4ALLFwShBXl/KTtUlFwn/0n40anORBGYc7uFOnT5m
3Jq9uK03xGphnIe1sBVhcKwPnGAPSuiDZAdMLLtUnihGSDXxFJfXq8hwFlxn
nd6Vmck+jlsCBs0772oboTB8nCd9IhcG5cyI3MDi69qej8kUDuwMUft0Ygt4
MkuOrxamyLJoE715noBM0b9ev5OkjRXTKUHINnFGDA0TQ0vl4OeH60XT6HPH
nLaMTh9XycqN6/0AdOxfJ6YxTZmtLqDY4QXyt1xThiIwV5RZGdaxdB/0SVu7
VRu8xjeWZhAzPyTmqgcwgb/2oTwbPlI9NCI/GD0YOEZ//Di4D/BR6zP3dRKq
h/pzp6Zhhix+f+K/czMwMJctqtvuTFn/74/0FOQ8p9D/Qlgc/gR4WPboun74
08NM8ZPOTMK/PL5OfLMIcP+3N/7heQaa/nTkXwXVAyAw7LJuYJJrG40RPR82
fVYntBQo+DC3uqEzRJ+b3gO+Kygbrwe15CYKw5KfmYGfHFY0OHCShk8jNZI6
9oP1iTHUfY3wstydK+XRSO+JQdAWahPY5S+4IGJdnmvLvelhtzyRK1BXVj0u
CJjTXL5Z//5ujeNBdsUkRYS0gpyURKpluwwjy6kPbV6rP5rLCStUAqDvMRHx
TXpgOoRQCxar1brITIoJzJN4BEGK7JH/2cehv3LJ5fZHPkMp9Fh64KMUsjNS
1Wk5DBx3JkEGIV9aRgQvBJTCaq2/wD/r1WsXyqlBbdj0Bg/Fal/G9Qg7R3av
5b0YDl56dBPmz3qmDWQb7EPibE+/sv84FBCjr0WH9gOX0OdV3HTWtyFDT7tT
eRIzDo9SpuPLOZVYTwfRT6dMYOJRDlW7fbzpvXrL0nBIHPzYengdLChetyR5
kW8Y2O2XCvlQnrzKb03JGzBwUk9r4TwSVFnA0QaQLp6QmVuTyfGp9BFDYsD2
e8YjUut1etyVuenyflJDqED3S4pTUy1GP6c2lr1jy0zRXbGZtkHd9gXFk8IA
paS3qZFCHXA+CWEdHf9EjVamA7+oKH7pnfSMW7DwKzdyGgRkNEvJ5xZhbe2D
FwsugGoo3kGiswhOG/7hnqMBQrMB67gtOM3iEP4Grrp0h65xg8HgzTy8CXDv
8C7jjbuKdUWjSZ5Ybg64GOaisZO/4jw9TSIvAc9IaBVxd4BeMS95OlFnoSUH
LfkjKOQ/GcsJ+/JSmQ66AAVr59nxX1jAO8D3Ssbe8d52DlxOWvOQP9nuAL5v
euTi+v1JrRBCKJ41OesCNJSVHrIWTbYISfUqPdY7KyO+STnYvBMOd2N/5qgo
3yAk1gyyUY+V8O4loDNDhQyNeie3b73OTeOJ2qSn2zCVkrE6Dl8fdw9mL70t
VSSv1A5q6pdkU8lejmGVtcwn+RroDhCW0xBuyMIW/sbSffzX/vxhExaWzKRy
7HhwGw2R59KdvgfnoGxUHNNthi2EQkInwfxCubrZDPiyskEwdgIKJeD1GsJL
mMgDFUHL7e1LMm1rUnJg9eKmpWvC1mCo0Mv1+giMSKwawkb//zmkr+k4Bjmq
D9sfTecFq4zgaLH0Qr0VS4rJmm7aAJgchP388z2tWQMXwXS2c1Fkk9pCGO/d
T1vo9TWPR2nSKSANTswcO28DW6Gw5dxZblKQmtzErO2Ae34FQkbyCr3nUc5c
MwZMfwid0UBe0uRUT7BRVfM6lAkXRXBEgAai2n9irCOZb4Bj8odn5RKkDubU
iR/aHvJdqa+GMMj+xnCR6HN0IBD7ItaZgYCRn81teiBnCzoFw5u4GJ5MER1R
LTPNokIdn4d5txhKNswpnZHXPS3vV8Jgq4bwGlEk8nchauwMmF2yXfNIbWWn
hF/UiX+xySCIN1CVVViD0Rps2KfQSUtf0z4zuK490XioOSLUqPHvgn2u7KW6
AacCltKaq0Cn4RWSkw3ByRhg72CyhNfbh3bZPO5pIppw0Gnkk5BHWwRaAtSQ
SpbpoWTaoVHBhe6Jm6TOqnZCIxSZBvtuVyxC5G9k0+t4tbc0jzWVH5jMydWW
IDbx0fk+d3m9JPJ0J4IByUVHgMGVNdEayZNcBCZP1nJYLV3xJBPgz6Pb6WkP
Es7/HVJiqnf0fXU12Eeow4B6x1xVuR+nZVI05kJQ2JSF0OV5v+SF7K+zHsBY
2kAqa3eyBqcTzQpngQVZ9zl8BeBH3nBOKPfmSTnPn+wHx/806KlTqWw7pXPX
bYtahm1nHkRmYzOXaH2k9/HYyac64IXahEpjz9kEj5X0YwKbuAMqAE4KRDS7
3JU3GEE8GlRxVdZcGfAQbBSzRBJNF3Y2BgBs06TOjISY5JWm96IlhxOyTzSw
fmSjIryTrdb6wQrhNA5xmwcLYgJqHiwhs6LTuORSExsC1Q/QY9AawGkd9hkO
e0Q17fGa2RZEkVmuACuNLwe5MLh2wr1JbN0nK/KmvuAwVH5dn4QWqB1eH4dy
miR0PauumpbL9P5yTsaKRDYc1NezzSRknPDTY3trPeAqmFmYfScr6DaaN3g0
x0t9I60pepkgHUjt66+CngFUGwtuupX9UMh01ySmuJ/Y0qOOa1qBNSr9eyq/
JMiQBoCRiv5TIwNxeKyY+67ZIRIHer1fZtXqzPkgjjQnjKPBqi5QNVNVf4PI
lX+ippDRZtzDP/wSvDaV78mHX8LHzbqM/iPArnavK8ZwijLLR+LOIe4Tsm6l
MKVcrHHrLEL9HRyH2ln5Mjoz6VExX16OJZUO5uQ57sHApde8QzMZEobMDS3E
FmW/qkNbBWACGD9OTUmboo5Yw2PKjYyY2h3PDF0p2oIUzIFovVXRuj3w5hPE
jISzNDq7Efy6ARg5ukxaMAEhLwQEyMITolI+Z7xu9GxErsyLYxi5E7meu1dy
fzohrTXDjLqaHfnWkXemx5f8YrH5XLRCUQeDPPggjPZ8lxXFaCR5I3BP1u2f
AkBbVb0Vrt+5wlA1BTUrIXfqrsxYS06nI94dozfXEg4+jNS2SD2J+ppct+PP
REbKUkJKoBJJKrSZVbqEUKHGObHEUWmwH/Ni40VkPV15BGlfWSZPu9AOHaSx
NLvC4hwLTvYVyHKkiubTvE9/Mel9Rq/BVK7+GsJhT6GY+jhb8lyScb/W0fSK
GvKiXVkBSPECKEYPbUywpwu0zkreK6i3OOCtjFMUy0vgSM26zRk70vrOLf0e
PgB3sksrSH7LsNsMMQtjdDpol40qtE1NixFqm2FPbUPsZeXWahCJWc3Oih8L
U3fYLocD2e975iJhGk8kamO9lFtBDADyNgaiJkvW5vz0AAiZYhb+a0/26Trt
euxrNr8wFAUpob9rF2K7+WtXf3+OdP/EjB9laF864VDNDqbT/JAnrXefLlxs
KGyB+cX5DZKlt/CzxI8bvB4J7NHt4yVja9yfJ7a4L/Uox76yrSCjnrCljzHo
9oUH09DJc2aFgUSq+7ihmlk7Fr4VARoOaFhLiWi10w1EmRGnOmxRJjWllIpx
iZWpbWqdzIbZuSVcXAw6K2Wb1mWwRpq5BXDf4KM63FiH6AzWQ8apHNVflAyG
F9Fb73ZAPTBMIIdK9WroEy1fU4E60cj2iVj/9gty/eqk7VgWxjsehLgOsxQT
ox+vf+boafsvLHKaSb50ASXbwPN7Cb6FA7HgHBSwG5igyjrjs/c2KlAV0SYS
FdIlwItFIIYrU2fDxvtiAm9Z+BvmL5HnyPM4zgC1tGcmRwyatA8UV+4LzMv4
OKiqKc3hy3gstqXimPkoS3zAZlfpVzYrsEPZ0XbXM5wYjkkYrmvtdRTl2S+W
0TNY3VB+EUsoYHyNPq7cGlS0Y0CyMDq46Ezr7op8MxoGR2xLE5ydegvO4tJy
CP9ccX3Sq9zCy4cLH9SoQre6PUcye9qeJYee78ccAGg49A8hV2Fo3hT1ca9e
hpg4sKbLuvhN3/MScoRoshdCvMKgIF0dHtyUBphzq3XnSok5BujU/yShRZDN
RWEbdKloT+rD3pmI7ZfUsVWptkT5TeP5NTYgzJqA5zs7lFfny8hw1t4LQNEC
eJCLBuRI9lHcOcOONc8nlfD6K1u/kl4ZEzh4pc2D/TuiBXpXFkSTiCcH205C
VajnR8bsFD53g3Z9iKqzPKAOhVCs/IkhsFjyDULMkg1FWOmF0sPWkwjzO2Zl
PKdUVxNgD+3BUaRqGJc1cNUJJkDPdddcL71R97qMRmz/l+jA4v23NSegMxGG
KNZjmM0X2EGgfVJ2MOd/bBaNcH6TX9L0xMb85kIi/XjCeyf6TqqSYTDtySYO
G8OIRMxDInImRnmZeawvJFM1z29oBAqJlRoPzKZ1EKG6e2wlKdETNLng/QAl
d0YV9RTrwddpG+TfGWZFy4Gi4nLTKiH2Y+7nrNwtvzXR/I+GY645kmyzUa2B
KB4nFlHeCfyqKxThci/OGTxsG6WV71mc5TQJA/0HSKzU65F4ohtvKbfmRQks
xy0YL6JlHHf7QoCYEYc1gBjW6xys3WFIEYGOjIMPdurvm7C4XJsnzSjruZM+
GjOfLKfy/+PxFQNWasHIRs/eBgoMiEH8pLGJc6cnOng7suGSAW16sfgJwTKG
JH2Np1QSzUcOsTw7g7lOdGa/E6WRBIzEz/YszvVhiGigKDn+QwilaHoKRrO6
QZo2ZxIYq0VpguL3dJ+dJePA++HpevbjWFEGYgScTvP+busbNKs9uRzXyO4p
GfehxWYyw0l8KSEl80iCEHqzY40YPqngJOKss5ihN0T7B1JJuGz+YFKF6NOd
LUuKk931+SVBpmVbsv84wyKaTvOnxZLoNqDIIzB5lay8Cx//1S5hJR0dVyXx
UeHHrFhwGacvcjvtKse12+Ii5e6ip+vKcxjOElT+2oj6U+2oYVjjbyBAeXvy
DftazKuJ5wWiFCMTfHiV5UgJFO50z9PfhjK00l+FaiAgySg+0GO1+hzcM1Qk
9b6r/Fp5f2e+QeHhPk/yYRzE4HY5UJJk+Gky83VVMPeg+JQwiPo6XSzaZd0r
ShkMjHqgUiriDgEzn63y9czNHln6kpDqnh9iTZuw2R/+fM9bMHjuUxBHsyyO
oQrYeIehK1EX1/YskKcBz3KZRWcafgINMreXldW6uz6Uuu0yva06oeaVqfjG
iKCnZmTPfzUKEtAEJlHNPLOBo4hwWxh3H4x8Pmur0Fw9H/Ss6trjWRqeTRkJ
KLVtfrliE/OcwXukAJhCQAyZ5cTufbHcw0e7aNgI1+uVSLof9uV5NhgphTY+
yS3/Udf0UoGh7lD6RHxL8HUZtA3C8dUpXRWn+yu+6NdVZKaFzhTepAy90R6g
Xi/+6Sm/T/GX/icWw3huYZEhN6NI6VnJrVzLwmCzG0p8TByck1uAioO2Zw61
J7Hvv7R0ExxH5ruupSS78cUEUdZ8lkGcvUOyCmXrgeUWA7AZ/z9Pqrkq7Mg7
wDdeiM+ElsqgSO4xhxvxX7EjPTyhqOGE8cJXuMNWqub1plxAInDqvw6W/ADC
iHNBQ7Ufd+WI/xpGIdJME7uVEUrTkmFRSeflSyLmkAytAvu2DFturx0j4aFh
3yPPFDlrWSkToR3YFW8TWHvqAuUjUsMSOA17NvSLA8iPT+mTLz1z0xKz7OrA
E+hCdOJ9KQrpwesoT2S1NeEgxNUW1NOlJVSTPeQY6Hc8dZ3JtJ0z7+gttvE0
vDV6pleitxkbVFEhB9loRODSbJaQfn0ozSijdUoj3k1e2K2mOlKuA/u+gRNx
pdP2hwYUgoUM/+TBuotSxEvPIkS7bM3c3LKgdj240Gmrr1d5235i2CNUPSrC
dbpW9qEry9TtSQPhowZgTRiB8LiQD5XN4w5919YEviYZqfAIMluJqtECry1j
oNbxQes6RXsRmV2QPvqiu20fpeWQJDEz2tfLBQtYWEpeVbug2ybtoRcbl/BX
jnAFZk9A3PW6BSeStpuN2+7Retal9Kme0VWdxwyNI2ubIVNtChdHFgBvG1d/
kgMrIuq6JKHkEn7dZTPtNdWR6vQUk+yNLoRorw+FvWAqI99T0vgDEtwcfLbw
UIOiNW1TXsoU2Qg5PzosWCW7bZABWvl64aKaH3p0nmdwO6j36l5l5q/MHFTc
Xb89UZt0GK5OnuGdnLL9BLSpmhn2ELO8TJIVIU/I+1StoC6zZEFC/F8AIKfM
aNDnqgmKjcoDo8Ws9BxCq1gQgcJt/FNUOvHY+T2u45e3/fMfyrRb64+NXn9M
KMt0MBjKluc0cQZbdd1aR57+17kPzt4IDZyOtLU9sQXrxhpo1GOO43KwzHpL
7F0tcPVpg2tHiMnefbPekYe7XC0+9AFLV4bPPIQrQIs1p+MYsiRCJfh8Gurd
wONeK56ouRUClWfORbssONWtO1BdVQMCipsgW+MBFzHBvwpqzxgf6+LGZLUJ
dtZtGkrUSixcZNDPDlvc7Qx7+VFJscz2NK1gBOxS8soZQpxobd1ekShMbW6p
0f9X3pKQQbiGIFKIKV6zXcjpRHitpctwZ/JcYOZEdjiNPmQzUJgSsebeM5nm
4JkeaocBTbyZR1+SKskAiBdbreJgaQCYVHxtLxdY7FmhJ9kW9lXQDyg67VVp
dVmQvx8IdH3rw5Z2HuTf0gFVKHgO5Eh3uPLez3U5JHuPwhnPeUwmoZrh6IXl
mmihNhd0iYqYr4nAgDZFDhdK5qtW4nCWxB6qbZCh7a2GT49mid4r09F/lgH3
CgzAzaBcooLAC9cwjjT4KDrQhjKM2ilV1VHTZT7NBJQxdEnY0ULtnm3jQaNj
e1XKtE3xdWMLkh13MwB3vdSsu04igQXBG4GdlAsPUxCC9s6ackMkg86HNPFL
VmXHyXxQ9/N2A6ICyFhff4rMzB5XVi3oR90f/O37fCcYbTL+xNYSFFoef579
0gmSP9O5DLvu1IwiAZSMFFUZ7zR1tErWPMU6XhhijDO3/H+cRzakTqDONnQi
5VOg/gda+wiTUuB0GJC9I2NPCdr5bFnBtjVwWMutyYsF75oJkyfyFl4RaMQ8
Go4mrKYB7ZjVgrXRdVbMcnvE24k24y0RAw9K4ovPgTFzvAehOIqKC3pAFatA
8klTW6/pafrxMqM3HGJxl1PqJ0QzD4sBzft94r85RgW1fJZe3F8zac9Iqq77
/jY65t29UZzMzHme914V00DdncsaHN3tAxKstLe6d4Yv13ZqcTi+6uUesQ4c
IWWw+qEXbPJa2UqmJgsxL5s2VX7NOwRM1wiVNbowIG+qw0Cw7F0b6fKklozC
BdDZ0KM7nzJA6ZUIld+MQiZdGTQRp8VPVim0dOQdbavyo61TuKFDrHWmLj8M
TUSF1QJarrsljrosDdZVHmPsv7g5O6YJfH8Mlhg+8+xhFKmRFhFX+ohjg6Wa
Ah0TZiIY5Z7vebna7oH/uPGJZnvKj5Iwx7eChPW9gdWV//3pDaTCNDiMl5WX
2h2uWPMBoaCUqXtx/zonRJK+4Zr7YctfUyD4nrvLIrNAzd5zfYAWYQu1gz77
G6AWwWo/CpkLXs5N4j4BTyqkn8fRJ1xxd1Bzup9+6lclelcFVSX1kZ19yuwY
iAKbEU1yslJVcfXsCdkP/k0axKvqAAQuu755rY/c0hfyCxULz5xda9uNRLqZ
QxQBHZVHwUxSODsP2cxPIARI1RNb2Bv5aPoHLAofnWJGA4vLwcCHKtZe3V/W
hFapnsOppeR2eGDLIyFY4C+5ZvTI1b8s9pqpVj7qR4St7V2Uk1Io4QN1IeI8
8m+QuhDMjpcTANbhrh/iJmPpLkzVpVcDfHj8gLuRu98YXFcS4008jdWNgRjR
jtzQ1xiP5HOHXpa1wxFvdSJ8GRWT5bf9DGhgqrvU7fjN743VJ3BhTMvfuHCT
JW8RKSxjJHJtWG8gNf2ejmEz5SASftpAaWP5v5XIUgynmZcfYqmoMWBKTIIj
/5J/lOT/d/fycJAdGs+ae+8NgOLW06xskl48z+TMHdGKBg/Cl5+qWQcCmd+m
7hjaGx0CmIPORFWtwIFD1qHTFOmAIdftFy3WpBUGSeXxyZ4s4JPfKcEZxdtz
puYH0IfpJdMIPhwfu3KqVGQT62qkjU2oSsx+c56zhMOTeSIJN6ThTPTpHhzP
OWYnDiBGgGe5t/j9hZIlWUQKil2xUB8k4PE5ThQNVY9zHPy/qZa8yR+hgdND
PMTMO8kfEnziqbbioibv1a1HNqN7x60cG99a4dKcffnSRjH+Jkt0YIEMeo77
SNgQfDEQwVso48gcxyk41divJ1E5t0B/Vi/kqAB4UPVyfzcSsidZmyXnduuW
ldMMbbVDmBeRulerBMjwZ7Qw4djfUY4Qp2tLxNWtsoNmHBjxNk66ICZ4RJ7l
4LjJ0p35OahTE8DTsJ25E2Oy9X0KQCtqRFLAik9nodP58K9vuAPT+ZJwFEgW
/ByIEASCjzFUdDygtV7Meq6xQa+A6l9d1/gRUVjxGCGzMporYuAA8QA2nHjf
4TnbDU/oQkHvNGsKJUACfdZeglfbEXu+BEB0jSCobDw8kfMOfQnbyXrSHfNu
KOa/a3+HMNStUx+LrFnJ+b9jZUp6V+1n93NxzsjNo0xzZ8m7cf620LByVVpx
i31SVKw6Hoi7wf1FB5ie2TjuBDKXGGH/dWwFG5L+XGnHNC8jnFMYD2nKQYOo
CTKM02zn39glCOpPP3M34C+Z7TaM6liGhdpk3QjjL2kpg3uAv3uqbTk304dg
Y9sOXP9xnCdIWIL1yUiNmUM/qM6mPvVcQ8oSv4Z6y3SwVkwKRPpe/YlkAJ38
WxZkMOUmznlUYccyRLtVrpC6Xmd979ENXoNCqxBGD5ESewxQQIxSxK9E6rWd
ypObJfWBzKxOR8TjY2Ub3XM9ptG+x5aLzq0gibwzFPLnUaqlhrHWFoOmWOaQ
6woEmwTRvuTo2Y9wVYv3abbaTaQ4VELzd1j1vMhs80ObUthg7FKZAYykPgZe
bYVHKFj0sAbDjQkDWx6gn1kT0PCBoUUGQrMJEztudtE7oiH3AQV/r5MOxW+K
p9+tIyyvwfVHARkmQdQIWfzfPh3f23IilI6cYCE1VTXVNhHODG4sJ3/aSvAh
O+GJMEOmD2PTyQRl3ZIfGXo+Utr3z4IGgZXuOTtWgdd5lpchMxa773mEFIWL
E2by+JRPBYpknMU2uKbs7qpZ+4SP6BGN9fuCWjH4CExhzYAyaODOIM2Rm5Qs
Pr2MOgTBF+kABzvCzXLsHttc5pDhmjQ10Z8t1+LF4c0O7Os+eKSB5rC3nX57
NJ/aQWcKC4nAr1ZIldqctvQGSWIpw+4305Z7ALncJsSzjLEbJw4DSOJzLcPA
JzCiV0SHgzQlax/1BJHgNFPYRTfgNBUNCoAWaMqV8Q89sxuKLUwdko31uVOi
n5hXL2QoGe7kp+mOqq5iLUPiXmjcIEwznaxqZtCdf2TlJj7vGURbYmEv+gJt
nx25uYWFoaWS9cukUTXbEgdHg3T70bc/SPxCZ97PqzFS2xLoXymxNu8yXAoD
o3bIFxhypBxRgGqZjpDcv2lIjAjLuhCu1fYTH0qHBc3S9adl76gdgSx0jWIy
Ezg1SQSiS8wbyzEQ9uNl7+MstcH4v9Pa7cLHVYNqPxt/Z5v4DQWmlFFBV7ku
RWK+XCedaBZu4Bx1/Nk3LhXVGHnnbEiFTGNHt3r199axmf0DkL1L1ewqtU8h
Jt2FG30vAQdbQLOpT8MumqTZaarFXLeR4inEh6ESw4qdNWN3O0lwRXtL8LTT
Tet0dzZ3TDM6YI5WH18q4WNHVn2s+ZQlRUiKaWojMu6JTHkOk7Ra7FlMutUs
qRuTgv3JLrkejK4uWA+QiIkvmS5uiiecneoqPXiA0szHI2hw6vJnIhaZpcV6
4UHGEkyO7jZqmqEVhZ7KMXYQryFP7YCODPexjFs60OXnHN+LBAqXRaF3IdLr
nH/qycRkyj6CRCVcEDbjkuEDH9aoJZttmftYRvQK/8fhMu53VWZXOBsSN0vH
NZD1CzoyiQ7I/M9+nG9mfAvtLFTs0ytZ0TdnCm780rXMngQ2Q5KBJ5WruUwy
/Ez02L3XNkZqPQwXhTh6zzzumlU2YQvO8GmQdokfoXdyu9LMFVjDokxuQyCO
ExsTWKWg7cYgIzporlDxUlV2w21U/Vkk5okKOfsjwhTPGAC7edAAMOT/j1Pb
YRBCLn5LBlYquOZE0BwQ9ZVKQl0wK0fAYlhDWwN7a+tmFDwzRPLhfltdpsc0
KVgAu7Ihjv0bsed33Y0089wthGTKxZ/jyzazYAukrZFIK6YnB3giSfsg0W0w
mi7WXixHvnxB7/26LjNi931BROasUKEoJ/yGZtgy5PqavBXv/XE0uYAf0JSa
Uf0TdLFT6E7L9kawCBEzS5y+J0NVg0IutaZn5dsv3kXOpU7lnqvi4wUFJAxK
iQcRLxeQIJJqbih6eWEjGQwO7MC0WW1TB+bFDfSgyE1FQkZtUuLgsJxxx0Ij
sGKUeHS2S1qklZ5Y8n1D+J4GazZf70egHXZaXLfaaYqSKYOrGqHGUNzmCFMD
8gus2JL5SXqpQxqqQEvOpYdizf3sCEMq1iBOw3X0r7R707z4u0ULwTTaW+ax
xepkx8//iz//glhh2qt/UB1mhYxtpuqFCWM2JG5OVQ8TnvQyA+3RVjB1p8Pc
eoruFoC4CT84bYWZwd0LuBHPYAxJI2D9+QJ4csxQaCbJUOobaXy2Gjn7QC0T
O6qEDqGcImU8NbnVWS8c4542psDMM6BkJdZmciar5O9j6F56+0vOV4kd+VNf
FQmEmscyDY98+HoIdLR1pdF8CkBtTHsJAGePMJ9xFvHXdOL9UH2pSjlnbYNx
9mX6tNYuB0cv5+b9uuSVAP7UAbxJ6ICU+JqGB5IBR7X2RPGM+OfvtNwDIGUA
okcHcHrXr2PSY9f1EVh0WfopTGB7n2jkC468QV1nFvebmsjCGqmMkoYdpTYl
atH3VBdaHTjQwLvXE6vgepPspZZMHb6LslHQ2LnJBG5tgejcsUBHWz+SrI/D
H0iMxK3BkpPCZ5eauCEYgVOP+0cGpu5aECZZSgXqqE3hcwlhNPXiu+vRu4Yp
P4qHT3dR8Qu6J4KwjX2Fn29oeje3OL6XERE1qP4w+IyT4oYKpzkAWYfM9AYl
EaR2WTiISU1U5xl4Evs/JdvqwQ4G0cceUTYHYmkxAGt07qVo1N92GmRBvrT2
B+W+HEvX1KdAMaSVYUHZRWunUcfs9yv02DE/nM09tJqnstY5dX1E/CvE8uBQ
FhSNGl9AM9JDs7/DsFJo+S1NYelFmFsjHth7pIQULMisyIvEjUB+vrf/ASxF
py/NlRx5ufobD4vp63wz79UantGFYkbJ/rdkbvHnGTO9IsQA45Xnl1mO5iuy
30vpUPNadWAqI0zH5d8ZyLq6NRTtU2meQGxPGnfsQSwOrDamf+DCaFzY1gGp
QvKuRziYXQ2Xj9VS9i3iIcCXFBS4hJIUBJAn3KlcgQTwaIu70gh5e4G4qKO+
Z5bIfF1nTtmiYkJECXsBvfWP0bDAZtgZnrXcXoB7zaBnfQ1tLJmqcQ7ObTj5
ERQuBucNjozM5TvFtajQ33MMlKw5CVp5M1QidZnwIxKIdz+C5KuEdFhQvYip
w30M3MFf1x4Oouf5fT+80/f3qFtnEEpS/4oMLInmnflDlpdJKuUOM6SCyvXs
54VSCPZeIrdlwUtfkICJzqhohvfLu85d75iDmhlRPZamL6IGKSxrA56t/ip3
5nmcPvshMhOwDAJitHVbTOVw7m21mts4m3MF8RzwvDmOBPLgpPYRnE+7Ir5J
g0QVTr1EoZd7VOABgDR12EbppaZPZZ//1INOWFik9vqDYMHUXzwoo1u1KuF8
AmDvaONRaauTo81onPKw4pvjN7xAWSpJKaBgEWAzLoVA2VlqvfmlCovlF6OW
kkifcmdiliwP6Cf0wtYx+qSUSYoJR078StLD0dGb7P3BxFIdddU0gh4ArBz+
OMsGX2wnOyrF75CQIpfpAMVE8sxcbPBB5e4t6kFUFkLXwtEUnPK2Xu/QCup6
lie9rHhy9OgWApQ1Zg44NRwGpnv38/bTNkhoJxak/YxwwOacThgw0JLbQQZ/
OXVCermvgMtLBJj30n7jEGUX6VoleB43oiYHAx5KcFQztdp0Z6P/Ame/mU/K
clW5QrcE/BGCimdSumIH/KUEtfYsgF11OLDc7TZ6jgIbWW/lYvu49Gzz2zl7
ecgJq0Aw3ENZkvFtOihpkX4VCczpcyPeufWFELqZMlRGjke030XyUg5tDOgI
68q9guQbWGobyfDNWGUTrREWALo2nShXRpUuqHt32RqykXcds/UvDes3+5VW
1HnCNDpayx7W+lgH3b1nw+1KUQyDYRa9I3OkQTmvHmYkl0K4g3mJ13Cu0VbS
ewf09y/hmpTRcmEooPLFmUn/8GGdcWhjx0ii7k51hmW6GbeVNZn2L2j+IEE6
EBDMq+EcWEEZ18Z4IFqmVMmwuABTRY38LBzJGWAJN8Mu6ytmclW8Q1WudP6F
zxNhZYhP7orU/oL6a7Kk9k4F8EinX8jNJHHiCd5IqMzTK4DYX/3fgKOew8cX
oGZhxD/ewG3B8xv0+Ag6AIUexgKXbQAeDDDDk2ztIeUU5hdXgtaZAs2qgV18
7G68Dg7XlpeBu22KO27wg7mwJmZz3AMF+lLs8nHLZ3++4f1QFLaYNq/826Ck
DPU5Ca0MEm5gUJ7pheYLoqCduZvLUnWaHnQDqRHA1jfylC6LZStL6sMpjpOx
9jZUPRk6sKBqSHhYTvgPsxFCKXHq+o8fTH+DANuBptEh1Jtd2TKKWge5X8YR
qBTc8cWynpazTjDQH9gDMrnxGhdpRzDW2rLqI66DM6q9os6F8fvicBLuOTR6
2I0m0poZQCqbDtEb1spxKF0odDaOpgOH6KSBW8/EIvJO5pcLglVnQpvaySKi
c8K4RSjg/PjYUnrIL/D7APS8fMjQ+Mr0Agl8Z+xJ15C1tAcWagDT+yuDz5pg
xh7Q6R1NlhM+yeKYtH19LsyodjvVOHWVzMCtyNxfbRsEJvI+oZQZMU9+hU8A
ddBJNT5YT9KX0GZdOa7MP4XvOQFRdFkrP9P+KZKID5U3ep6Drmh8qettFgaO
89uJotI+Bghpk5DVhzY4wJNcDsPmZ8hrmg/n3KcC9pC8GdlYYMjlNqClIic+
kUkcYbW4zUXcK5kvqdYbfEDwECGtS/YygX2KG8CxUKb3m44cniaxFhiE7qYm
r8sR4TvLgNBmHWwr71Rpuf4rdoz8Z1LNISvPXA2FBQz1gxccMk2bgNDRMv4i
zQaXijMD0VRvOsZ01vxQfpS8e6gxhrHMbnDhzwbJswR9CXcxfWH/GJb3OMmL
WZh5inu6r9FV0sj1hRwvaKUW0Bnd36cznS42HXSs7FISyjxNf7TcV5X6wnAl
FyTIiIcYU/71g0D36x+hDqOOwE49baiOe0PnZ62spnn0hvWlkwf3FpHpKQMG
X9CWb8X9I2cQO5UVYhM0A4P8XX3lML8yNi4163QwMnRYjKP4x6jf9NsdnaGe
9IyRnaJ6dhqmwjet2mLv1rzYMietOaCE1h4+uk/wPDK378fSdQ4Nd7NxgGuF
8GOlTwHzDe2zXEdX5mMkhM4Q6JnOHac3KPgHp4y4utTm8iB1v+5rADuBz3S+
XD/W6U/EiDn+xzFDxfOXvBqwnBUZ4NYkYX7GoguNKo0GnrbJxf4uwrwyfAum
wvD72jmzHh+jEg2FGfn3qm6kOr4naSiyiaXyA02Hzx1i8eexl8LBrnNQr3W3
8aT1H5bhbsBIlcp7NuIDdjC6sfG3VeZbvvJcJSK7WwwQkNimF+CjjARtfcsY
lmCF0gL2kvKieQbrglCrY7msM+4NoOxq2bb26wO8dGMRz6athJ4xBsDrUnNR
ofyVJ1wuGZTu8J0A4fO/sq0UpAW7P8C1TB1xPGYexEOetJvw3FjGmWx0ya8i
oSqn6YtbeUc+ZM5eSxuhT4JQglZa1p830S1HMqC4QaNmJZZQ73UC8/Xq87Af
N85NOObtAvn+5U3a0U1P2JrWxM0mvrjj7kZ9p+yQcZiZ1Kf1HR1PMo7OCZSH
efCo7r2dMsXvUv4mHThI1mWSPL3yVy1kAAQqc6U1CjZxGyczcZtffaBRcQQL
k1s6HJ5M3i/g5HgIQzCmBz/V9cwPrBPa8fd7AJVIKmF7oMj251AR7mpWp0Ck
n4II1jgzqJdmqdg6ohMW1eUqKeiGYcU1tioBck+U+BfPNF5iRCiQAfGXd1QL
/j/6VnLsdOJZnLRzaI5vlQJ7PRuXUodcoCSP6t9uM11jpkee6WarmDEsKoXM
JbFfCFQsOO2n9oxNSmcfrlnBJ0Zrruj0B7k6el5AaVbK1FkM0hHVF+pFr6kA
8kAsw/bpeIzzbVoS/fvrck7cpfViTaObJylpXDuz3WsWDWXRcQwc+jdnhcI+
Gczf56IACccW0slCFN7tVO51SJnTqPcoHwBh9K0smvdgQ+0WG84tElqjRSCp
y1eJ2SAPnLB3Nsxb5tNVI+WvAkozfboL5T87GcaqrrqblZH5tGm+2COYnUCx
Th7+WD8huiAvMHw7RLe4tNCLZCzVZcKg/T4/XKyHkw+6s4hojNQYjZ71ijvN
M432AU+o9SDVOR0HFPWcEgzNF6KQQ2KtUP/63Bm6exLIUmspF52Lb5ki/OId
QERRjGl4N/A35eHny8DVwFG1qfocuVoCePMspY05EAvPkC37IxLc2pEek6sX
prqd+RbS7gbm2WcpOlYnUb6yTBNZwGfo+6R81VYae2O9buygPmwueztzQDR5
zCmFOv2RjVS4wLgtcy5pl4YGQpULc3Upzq3BpHgfmNLUzh8gpevU+f3/R4Yq
hXRQtYKVKjsMKQB9SkzPwqkuHlgDyOL1PTP2AED7/ygHZ9WG/KDx1HSLYjP+
uebJOSr7QGZOw4Nl9GAhLHkaGcgoVy/9bGl0N/UPts6UxpDePcFgpGFOCAit
Ai+DtkI9utfDlF5FIJwEXfeiRxphyQ2OHezA1p+wEqgCr7EgaeLWicxFi0vo
99z+K8pTz6sz+74ZO3bx32oHiLMf++6ROF4Gc18Is63iqnS/1lz1YN3dRk6P
m+McJ5u3ybyivI1A6UlS96ep2GNy6UBTwtY1zlCr+YH9J9H+29pLzxJbSmvk
5USv+br3C2l5kLqSF1Sj4YF1msyhPH/swqS0u0uIT3PD2CskEN54qGAeZkXN
uHUtfjE8YeMY8D4ax24LheV9/QNXgLtaEaAM3/++J3QWVRlXZlfKcOHDEUhF
AIu16Qv7oEvVlnL1lMGpQDvIEp7isMv6+cETiPK/VC3qZJ6ztmhvZkAoW2cm
jbZB1ed3BQBzKlL/VjVxPX5l6czPjol3VjiixAPy4SXRLf43ZxwbNCPNaQBi
wJ9Hezj8zV3rvPGU8RQFtM1SmR7lyF/Y2uwa5nKSpZt8UyWhhICXEnDtclUx
JsBA+hCqFhSMcJgCg6IEaYh6eQp6IO0HFcAgbZ+cxlEuZBdNbSvlp3Mw4ZEZ
6Knwf7fKWjvJWt3b3ucx6qBY0F0ANjGvizJryampE0na4LYkxYUXTzaYgUpH
Z3P9vvtUpc3MWKjLO3a9gc1u/fl8qXktadJR5bmwWiEaPVgz8BaObfOg3WGx
F5pHUcCQ/9nZqL21lc4muh/VR6Fd+Kss/5SQ0eYetb24cuFyobrMJ/ETdQop
ndZDHObwEGXGlU6D4vvEq63E39e0HY/yrTF+0JooEELggEMsMAl/n7f/Nxzc
3JLOMyPv9IouOsG4uA01erLlkUQBsPlS2WrxxOd1cN/63vjPYqvvWXhQ1xbx
1S/4F7n/nxFbGVWLDEl1ICzqFu+kvij5I3gn8A4FGlzg6QEb/VYBSRBx9aYb
ciEU5LqurH+b1z9hSg+EL2WJGDzDOASJ0eXiBbxPrrIe7eYH5GzMp55ZHGMe
hUoEMkCaqM/gVXhVpMViuSMqq3+BVN6wbT/66Ec7uq9UTbQqT0hPxx+w0Tlb
o/SiS9q4k8dOyP6/RG9oTsbjnnY4+0irbMozzya4DlUuCXcweGRhd/QYAe5H
Wh71hGfxv8hSrxSyD3DtMOL+rdveBDQF8ruF3OS4CmsYhDofCZiSXEx2y5oH
D/Q75sXXYT3krB4UlvvYFRo0bVq/DDqPrH/3DOI0KDePVJxyRIeoMVNSvfeC
IUrPM5/H/S5tnPr1OJ4pfyZcF/2lnI9QX5AtDuR2fEhkar4rhXkQXLBLMyRn
MIjn8K2gKRZbTosaIzAUFvYL9YbzeW6o8FZNRg1JFvtxCnR/+b19uQkoYhi3
zNlAsCybzlfniCnmcalj/DFmCAlzfLAoqiQxe5qeaglrjERLrXHlgf+HXprA
ESPK3tFjhojhSroq4CByucKFsOzX6COESKqnEEQIz1CnxVP4xTFzRn16nVs1
QaicuKIIjwwWcnLEvbH9wf1R9Mrdr8NHHN7a/XThEKOQukbcPsSGynRZkfYJ
CtiWABojGHeiPqr1YvMdG3kZrzN3KGBYy4WWXnHGnZ32NjlBshgGH+AEolTn
J4sKLCWH3kjeyKKJd0pNk1uA7OnzEiUlpzRhIE5hO38GCtc2v0VVKJcJve8o
5NhAYp1ZOjQ/5B+31aJMAqYRf0uFUbjBjmq4RG/yi45H7HBgzXTdSyYa06xN
Tmhz6AAIDtfL8dBIYluOtz/9ZwF+E8/T2FQpSN/gdaXkWZGZ/dsaTR1LKZyR
kMX/y6d/9ruulZo5hY3Ppk4RhJohs0YczIsBHM6YtcF5C+ytFrmS9I9omiUt
RBjV5n7OTPLD1/KA0riGJOF12MqEygTJdtn8IsYjlgRPC95vxA7fN2XhjhJl
AA3Bc1sLrjw7Ing1K61Flaqyjj9zpQkSr1ccT3d70rmIzxVXKZtr7SPQLwet
5O0N/jBBZNyq0Ur37QfuTBsFAQd0RXSRDUDTR9OiGUznYZen5YQB29OlSNwY
5X/KNzw2flcuRgjkmOUte5xmdXtHddHpy88jC7NEQfRCco2X3RAqb1GD6nRt
UxuLMJAXrg/ZRV4OmsonAHQpqfQSCLW/jMl2zM8nTFp1aGBwSG2IidFR8B0y
faKz1cIxRyN7dQ8fhI34EEyFyAO8K8lkAbHrYpiNrHfrEzSZx5lHhnyhp47S
RIOFqkxXiT3CpZmh+rhh89oVCygdYT1RUIREtEHr7VoDHx2BObsltO9TRn+L
vawfmtUXrQuXyO/wiLeCaTJU35XJuj1CAn+8mNSKuZgM19i7iPaBY5xdf07+
eD/xKdTY+bDYsGOjnb4ab7gjLEtJR6cmC+zdvRBHkAIUYGIERXKm2GJFaQPW
FCMoqBhb7xUQw5saHWg3tMf4WdPlUHFZSJZTJb7q5HbRB3OpTi2gBWPHSXH5
4X8dfSCnWBj+SZcQgSEhfEEizQ53Z8lwe1adcozCIHYffuvB2/HnzXlfq1lx
Dk20Tb2gRbltc37iDEG+XRfJ7CoVKzbdD90FTXXiLAqcfuC6pechfVqfREit
8xuSCsAhtsxIxtKK+M7KVsMWfkAZaQ9SFqFKMPa7GQ/6LukOtd0wxH0RAnA7
5qTwyhi4lPywmyzxUQOE0t9UGaLszungJnCXVci6d6f5u56IbGVHBgfo8SuJ
03S24t7KheaHg9e6NiTYYU1O2Yy4W7LdlHda8ufM3/E1a6LjSpuPIpUSHVZK
S4VCCtK9+0rgd2UivJvFq30ilNx30u2moa+8EFMQm3sL2pvW/qSl9cqW87Ol
A5xGgMiiu2uzoivmrEFM9a80UyWerALyAVW2bJ2lV/diq9NiOJgqk0ZiPWKN
hC964w/KKWhydUXVOykXj9lEEp8ltcssWs2tpaoQVB1eP3I7wPiaKSL5i2Al
0nMtbFUO//uLR0nF3zFyf3WvRSfSIJHrjzrlEdQEt5e6Fo05bMWgWWQY0ix1
ZvRlF1Rb3eqnaQscAUNKqd4tWbsSsjayP3Np86YJdtFpXo3+S3hk+R3T4v3E
Dihsmx1mv69ogVNZUKJ4B1IkCBx3kyMuc0ftd5s+NX9iYTqfEJ6aOWhD3yT7
rHL9O1Ryv0DMKc0VNxaLQMa3+RjxeNYD6VpcDLlsgdOV9wK08dM+nZtXwRyL
dSmFBO6xx0QtqeY0mmJzfwdLnKbcAJXlpUnQuATXIqithvVK+pbtaKnnNjN/
ZC7AhC4vqFDaohVCJYCSxnn/P+ASiSEa8IEXe8RBuWVzM2WRw/4TR5VOS1b6
75Mks6SIekkkYkPQNHiX/bZ49VD0PWkGvTvS63h2uqFqmvMayg43foSTul3F
wFBkbehj2Wa+1U3WKSwFZXXAm9CrIlnMZJuL/+b4DhAnILTM2vaQwAtbPpqK
KzfleNjGn1v7Dnwo+c2pbIsaZFwXXOmfdjzOg3BXPAjFYvXafITXEVw8Y3TK
nsJxrjBNTbVII6WJchkSYhifvYY1ny2ZTVryrONErEV1NluG3hbKSX6XwGIJ
F4P3HfFJhFH/5fAvAB1n08AGWHt37Nf1jFZztcE9KNxvQLhGu0Ngvgkrhk92
Q5ZGs2YkH54B27zqRGP970pJKAt424LEtESZUCV+Z6sDlSvpzeY75EGsiZxD
aS3fIH2HguUZhZdF1IzQnw2R/UiwTbvPVtqdlkv2tJExMCsvtEtczFMsMk5e
XglsttyCZ0Qv3swJsJx8iUlv7p2hxM6/7Ve07WC/mYUYv8MvyHtPvzeGQQ9v
YbyjmR51/aAXJ73IcG73OOjTxq5OpeZAgUg8YMVTEmAx46pXQvvMZQOc7Zi9
Y/e6K9lRl+SR+vxHaJUnPGIWggUzr6NlYQnUQEzTDGekLkcrnae7UgXOuKRV
UIczHfEOVgIJVK8VxvRrBcWA8NqNSEl196gJtu6Ar+3H1yTsXSds/VVdm7rB
lg/gAEn43cIQrDdxojaf0429hGbLY/50AK+xm47dkMdv4z0m1CNIqRRoUvdP
xu0e88pu9IpSDI9QvKhiNjlTIVdmJ3XWGAMeGvjYCMsP+C3mUNE3ZD6sUpQL
ys12+Fx1ZlB0dyx60nC5/LOy128WM6IU5Z7xCfVaH9GJtsKUqUKZDkHHRy0l
18Ok/WF05DsT/uTAPtt9Ryvr6DF0t/cCu8U4QpgIPx1UPFdokL+OweymJxkh
ohNjB292TVm7KmSm+QiBV6wD0+hzh1T6ZVV0XiBV5NOYx6k2i7jnhvjN9vj3
lTX6H7SM9emgvXaZdPq4DivMp4Ox1Ly7XoBJ3z3HX2+sHkdep0MKNK6Rvnni
cgTc5QY39WgzmzJQrX4IJ4mgCpuamQmIwT/kbLQ+ojoMpa0YU2bSOtcRkW14
DkXFHLEIhIZneA9cgpC8PNS6oQTsSDGNHlyB58Z7NIFP3h3CHnprqzO3I4Q3
IsfYm+6BOJXs4rRGQYAPphiwhr6mDy/nPAqayo33mFG9WL1i4LIS8fzKlGBD
jkPQUBKnsIn3FNrJWEZD+mCaywNU376naILEKyhb4YTViXsinKnLxU1Jk/vT
M9dKtS8+UxU2k9CaaklpZ5XytmiJ3Ce03aDEZ5YhAqyM9XCT8sbEbMVeRu3F
6ioQ/6e4INJ0WkzHzZH/wOCAxxJMWZ0PjWeJgkmG4NYFvLy6r2RcnvCCZjIW
po2e5SAbr7yRL69qwDCjREJuDKOEXxkJ0RLXIb7gratElBDnb4VlKoi34zQA
1kxryucciOAJWw1aPxh83UyDs4zIDMMaZSf1OfhAsfmrnTOjhup2T+tfPI2v
D/Qxq5COm4M5qn+jHd/Fk5nnBEiKj3i8XRwWkkPL2mu+sCFBCaHsHua5aotu
gTmzJUt+mnb27hoY1Ic/MQ4rLKB0m6gS5Sf1fy1cMHc53cEIVdQUX8R65WLR
ofX6BKsP54gkq/Ju7z1re3zk+n8FMZDuVukR0K7Iu7v9+FB6+YlaksXfh/mB
zEZpDrp3t7bbn3X6rR37cL8Qw71X/fqbUyQuvMUcyE+A8kQyWE3Yypy8YUTi
LRMGROwEI4sLFweD9ElrBeUATktDRdvcumuOax1m/ibckP3Uawxk0+X/BPdU
LZzXsuHBIe/USSiGi1wIMTI5LiW9Ux5WD5XcGLE2I6lWd6WoxYo9L5kDVRgw
rZby8ne2U+zkpCumUlwsIu/y7PLEdimlhmzItrlXrGmXwRMpXDjBJovNAolu
BekcZyZDnkHU0ap6pi2WhDNKoZG6zpjc8sFof5yh7YDts5+b+lqn7eewCSsz
0ZQEYxKXYq4/sS/SmxLfUFGsgJW3bffb+tIdMSZf25Ao1kBveE7Yz1L+R80d
DJMKECEwEU8VVnWZUcmo3tyVHypu+z/eIpfrPGjlvAfKkfvgww5yw1abQoNe
LgGpM7KRQy2KaPVgLy+ie7zmrZqgX5JYLfdGeg9EmTGPM2HzEriK4yw07Y8R
g4p5j1ju/7jKd6YKlLok6R38QedwDS7gx+6h0mYnGH/HD6lXw6TAhd94mRM+
7Pbu6EZNFRuZXlAx7O20KgyL1tQxUyx5lszq6ldUxoTybGsOiTPTgCbXRU3p
TyIDeK1zbaAfEp+O824n2zldEazWtsDxDTyGPGcuA6y0gEQkFl0YJz+DNglB
U7USTs8qIYkGrJq0uWxLsM5Mel6yqXudtVWuExRBO38iF1KJE/KPsOSXMeID
bhZKBdhRIcvK+5/EzPGEB6JZvSjr4DwqRA7wbqP3aDn3F5b6PWblEXtullRF
hs6cs31g525+dccJn2wZdHvcWOqxFtVZ+H6+0kNjLd6IwTrk/PNuW1HmoIAc
Wg3QjRIhgL6Ot09p+WgQl6hh1WzpMgMzM0utVmpCuxwY8wnqo0W9dFGht12K
z0sxlWMzxRYquzsQiYIVWVTBy0WMvv9kjBUdM42ps84+it7eO0ds1uaA02eg
MgghtLQ0Ql5dXIvWnMmR0JyyKhYxtY3h3OIdv5/WY8SuiLAoAgTnjZYvSfII
X2oCSQfkffn0EYWtRYcy9r/7AeDqA/JINLQHal59VMDqmZdAqCob8Y46KzjM
28apTMTR6Tt+HZSTPrY9BMnUGEsU6GcCIkzu1CgK2a/AvQdUZlcD+QNjek5D
g2GIDIfCKE5D6Q3LdmIL+vaDyYQ0CREbFU4sQW/xKDyAXMdBvSl9J3I+rNWa
5jGR9tERftXWT6p6sWKlc3YJIHKK5C2A06geM2XrOAhlbmboUNhkNWmnR9Wi
eBLDvdikK8QUzwFiwOrMltz+d02cP9LlNhEk3rpp1t3mklEG1YqiIPyTjaJ2
IRHnYCy48BaMbr+yczYk5cgtzpBGhSrTQkbQPkQqqtJmG4lqAOKVpaQLGfDW
ucJ09sp6TY4fznrk5Px6W96OyheTV6sD7dRcNAWdDTh5667RmfY7sXtmXTTV
Ilzgno2P/2BD+X2bjMZy4jR9zgsq9SEpWzC/tnWAQIhSRTwKdctdeXS4SKHN
mz03ZN/ymXM3G4Qkc2xWvLk/E2rGkA27hfz4ntMyTsIg+6hn2rgyrLkX5++M
aYcV6LcaNk1R9nB08odPcL1BmB/t9WC+PNskfEDWuyQT/RISexYQOUH7yWtT
Mtz8vE9AKEMAMmndrMPm++bSa2bvB7ipWJNM1T+o8bVsNPzHs1vTUPN/Lw1i
EiRYl9dOB3HV3eRIjRKeEhVIGjlWdn5UI6Rek8+eBMy+9Jh1f7Kq2mVvNtwt
vo50MDALCFv+8Zt9NqciBik8d+EKoQ1ExQ3S2UE8ySdxxphv1BcyFB7aK67f
uVQzeaS5Nk51cTwMgT1SMvFgoJ+0dTmMShn96/Vq2E5mJl8H2zOrHeZ+oAle
Xc26KIawPqKnKxJc/T/wgWoLj5jIelCy1M1ZqZhxCUpw4LLkO6pQ6otI9Kft
POQ5SW/+F+cxUpAPl+GCbSQ24MKcUnzeHXtCRE5NOKmaIGYpgICmgjiZlTwL
sl6nSfhGaIpakC0654qENUW84LYfjQMKjT4UqhvGBDRpwq8yDGFXc5d29vFR
W0k9Id3VF5D0El4L/epPBy5DrgLiaRDn0Q0FDZXRttDhonEvZ0MVzAlCbfJN
x19m/UsTxYddhbYkw1zCZxF1mbd1erzoB38Bg1sIzlZ1NzXBxgQAVmXmITJ/
O24iuo9cSs6mpO91bATjsFTmnJujMyErj1b8bVJiDmXlwi5itjL63pJ/145O
9c/ReX0qHcI2Rycje30DJet1G4hUcXYaX9eDDIiwOHciixxXnI6FuymN1Eq2
WVk5ANtGOU97+eY9JZ17aAOApCNl1uXNl8WwKVfQkckuFoVnw4fIyi6N9gc0
j1Nq9ukJ0M/vjmA4uZi3uoKaC+7rWFRuJpVmNx9vt7fGRdw3J3lfJKvKdjcN
FvCRsriyqrrWGLd/uCBLmxD5oJJG52VCHTIBi5b8I42+QPrkSmRpbu80lBO2
0/PmcaCTV8rNvN0KT14bbNMa+zQW1X1247ZqIgWps6DqbXfBc3e5HChhr3gK
59YZqhmumaQQPh81ZF3fKeMv2ygzofXXt/elGsVZtF1OlQVQz1RtQMoUl9m1
M6JAB3J4Uf+r7AZH9Hc79J2xirfUzN0Ql03ghjz8cLdAMu1Y7vRPgkE1wKm7
0LioDSK8NFvckTutjVyEsNPUhT+i19d7cXA5ni01axq0KptCnLUoi2cfTNHq
4wMiAfN4nU5TxVJHAJagLVE+KFRf4Cr0EA5i7ylT1jts+aTBtPM2LpLPig3M
3FLgPdSbb3GPMg/IWqfYYLU9pMYK7VrgxPRwng/IGrZl7GOfbVngb3EFS7Tr
5c2G45Ws99UnsTHkVY2zaEq0TUYidvnqP2DA1z37+apJo6S0fxigIijKCzxg
SWQHiQuwtJ+tjdk3/TP3AqLOVuVHziiBn+3a+QhIeMiJBq3YNClO59qQ0Lmw
GtpMmQmqQgtJtPjW8g+Y2hRWJuExDgnKno+aL9VNcmZrI6rE7upshuoIQDc2
9g8eaPKsuSPh7EV6sLpXApXt5VmmNEtuNJrN2uWEoUWKvNONPlYS/xDJAd+H
w5opC1l3hZwR1F8bzgteOq6BuQpfZnYEpmzYt9m04UwWq/djFKw45XyiHc/+
VYrWWpB0sr+sEQIWTuYxZjjUJCNnrXxZvsV2IWC9a4vbSnmAsEoTfQ6wiSbP
5qyCRr92XytgqJKJe6Pd8soK/1+vQagxMZ02tW7B43p+k4qB9//2ZkSSB+qe
30zNEx8j1XQorItRV/2W2CJkP0rTonEQbJ2E/jOYYln3YJnSE7nngyD9Dxn3
5OFYUxp02sGLQLur+MhoLQlnNRS8iAaPDSIz7aqDoaQSjVVW4k3rTRWRCnDW
fhAShE6z++YAL1CMfR3DHjx4PhmxFgUV1RWbOwuc7C7w9jabzwUua+Xtg+0B
jhnX52kQZYPVTofUz/gwsyaCNFNHwFSubSv1aV7+x81htzFMQPDXfb4BdfOj
7XXki7RWJlQ4VTdapZxfCq+xd/FK9aEgljOFV3V97ThlfDNLKNUO26TbSZig
bqt6YMe88KS23XHyN2cOM6DCmYuuO4Voml3OaNxY9rTwevCq6NjFcAeNhyvC
WXhV9tJL9L7T+g/cr/Z/BQnuUMVeFuGl7AZYkX0oENMd62gdvz8v6f6FSltM
8aLIIV0JiCSWcbmErZi3Id7bswm0pEImAYUEStw5CvX6nFxv0myv/K9PWqRW
wEkY8+fJbpe2edO6iNbCJ58aWQgWkAzKwuFiGCcPjtuo+j6BORYMxwP3vTP7
ReKL2JyVTczsuBhpeV2pp2ZHCenRlK8Akbs7Nh5WvgYX1LVmNT241wXuUIG7
CiyuFwFb/x/hJl1maLvzUtTs/Z9XgkdJE1FAtnOQri0V7DMgZgagNs1dTxB1
mreLsvuHbqkxPBHr7WJfshwEGSyeIhRTKneMcrS01FRB39mkY8Jz6zjWEE5u
9eRVBoJEjsZ9N5Uz5TK3GRb68UqwJjJ2cImCsDlwQZqTKpPxfIvYhTIAu0XL
K6YDsnGIk1a0XPLroz/xurBXNbDsjSt0lyz0EVzCGhTiRJNXqG2aUmPQoHe3
oYMsT8MxgIUkJJv5s7x1UXgUZUnYlHWeVzZPRXiljZ5vME4ySiSeWsnmxSZu
aTWKuEffaa68bXcpO3Ruvbg3PrBIvRmUQZ08QMu0PGHo7GS+bwg+AR7JNugb
m90tfgycy6gA6U+8MNbazj7j04oBlfSKqd+Ldoza1C5M86WrsBOy5KF1dOfY
wIRgNT+gV+QbjLnhMP6jMnuFE1oYbxEMknbOnbTg2OhkAMNp3VkgDeHRSIHk
QPD1wXqZQ2ocIJ8DOkVE/x+MsG+l4h1nThr5L2VnsKkMa6/uWbsyRz0lgnoj
5HhVMS/QispiKvu89N/OQPHxOoPSLM509lJ2VS0JPLhlTeJFPy+NpQofadPg
dTUwBm85piq3QxA6emG5lLQFmtESjunU1oATAlftobDqeLpQhJ14EqF7W51T
OvnC6BN3X4YdVSA5pEDCM3iygtrDqwN+ziMkG16TXD5Fb6a/LExoYQuJuJN1
cCygX0TnE9fZHsKeB+maDJ0s7j71CIYn8eRJY8tR+bcS/krZ9P4AIB6Rzm52
qORP7/xUIiBi+qbLw6trD+R2RrNmPs+yI3y0I2y36Zh6WRB/xdd/z2Hj5i9/
mYN6uwchklOw+hyGCFEdxCxP4ERlFpMLQlk8TDVdahbycjrtjUFZ/OW++Q85
W0Xt5Ggm2RCBfolibAb++bpVlpfzT69Hul1iQxzH63wi4GKRcFMHJBocSCjv
5qVe0xGVT8LvqU1mJiGyll13TYTf/SK1LoRp7oveGBFE0GEQenyUrz4pPO7s
QRbveuLb3Gm4O5eenKCEqd7vEzDyPRYvzZCImmSj668XC9t3+H76ah/vxmm5
rdBHeLSFXqr5U5EXOoJqj1mEf/lAJHuc6juxBCmiApmtUi/xjg99E7N+9WIo
B43k9lAeckMRGVAMj1jGNADC1blU9Tm1i34u8Pzt4/kWQ8vRXzACdu1ndlP4
PceGC3+mzCuHilzyjctapk0U8rXiSfjrBlhxIGcscDMeJ79f+gsIwuytIX9g
WWBPhIzXYKfmiXrZhzijkwirlmFXEPu4wsZ2OCd5qb8utEjQuD1zfqS+Gyx6
kQlBIrEp2UMPrANTsJAcrplKLna9ijMq3rL2ZRBPS8kWeSdyp1hsu3vUjJlt
oXaJVanjbLyL7vx4gZqGnJxJ7k50dptTvdjnTQ3/EDbq36jjmAVxMwYfhWeE
00pas7O2HtkJaNcA8JmycfteOwpSB1j+/QLB7KCQu85Tu/fT9PsN4O5I/lVx
JtrM4phVh25XH8lkNqkGd/PdZvGneYH/4wD/0OcA5/B3JdcFZzdQikjTybP3
CyfjYLM+97HxtqvA3FiwFwETOM1GXQuYz5kRaQVmSOZdU3ggVST7pHTRkleV
th9hzV9fYwAeZxqnZv0Q2nNjl93jVjPR5ml20/vGWyW9Yg+Dah0wdE2Qehvb
kz8hRIfi0GF5CROjmT7yBghxiCXUEef+m4HsJcN8JQcz7rmzBdJjpxxkwE/b
P953Ch+YQHhXPXOMYv+u7vy87Pu2IEP44MT6M+6XAqcC3X9Okdo6ql/AJ2Zy
mSxsVVDU2e8w5FxewuLC850dKeI4T/4RXkB/7SRuPuon1z2HN0XcBmExDKVl
RvM3SMO0cow1ASlBCjfpBTbhqt5WxOZxgwWZiCyaAFVElrHcU173TeUChck/
+ee+1+J7bVYNOiO+wokP62d24W9AWHjaZa/63FVVEWs3daOhzqEIIB5Qu3Vq
onmhO3mlaDopgsPncJhRy8GIU//+6Z6U4qsv2UdiG9AP6mdopa086bnJL3y+
8qlEY77DMmqdly4dk5CGE4nCrrZBkORciI7SIWvEWWeTmBm059J9bpHZXnIb
WG2DbmCklbiAHMZ/SGsX6inGvedumVBgIV7xIOl02gJ3/4zOCyKEQbVXig/8
a43sq5Q8fmKg3r5on2sxywUsu7PqQXlPNzxk6cAk3/tRYwD5fNC0WzlKaf/N
9WKFo0UfTcUfmFfop40tKs35l/CIGgeHd6/z/0SvBpAelR9+W4OtS7Znj3Hp
h2cOFsEJnUFbFetmGgCBEpyLvZbsmZK8R1VUcuICecsyuJu4DtatVBx7oDLT
bRkJzwZzU6QYv2EdG5oEMND8q3vRuIAVCvbEZNljfFczhg9DXv2piNLL35TH
q+82XHgWP9LAPuxbAzRdGB3odDuMVJNYIj70lCFJ3eLuyiVxhqw56RT5AnWz
VJfpUubIOmqr9nBJKSQUyeCVfHLVDggrfVmqA9UHcS3CR5f9T2QLZJ+O+evT
XSk9wiBxUVxKcLOOZegpeQ+7Lm2195Bv6+WFBqN63LhsL7cj/2H6Nsmy9+cA
sYbzB4WDtxwF/ECMQtL+jRosI/7WCFgoaUaEliVCUrbgLuGXaB/K5qDMcjf8
KATy13H0RLL9MFHp58l4QiC5BkNtq/Y31hB9awIIfwmsOj2Y0YdEKRgOp9Bz
qVNw79yWfUz2JyOr4GmBJGW0QsW58zqH0FpT6Ptn+o6u7rv5/X4hrAoEN1+C
wV8gdqOYIpY9s65wWfTkLlPivzo0NdRAu+UfoIAFKcaBWJN0VlZfx6bbob4h
0bYXEU4U+hiFp8PbS3GRbZw3jA82ug3wPeaCRft8i6eyN/oMYxOfYsWkpLUC
KVdfCHqVXJNtCAQPcxOiv+/Z3+XB4FhDGMLzvvDZtuacUNerqmG+eWfkSavE
4dX86c2peRDV3mvw4IlbUBNYfODKpB+i6ks7MA2HV2YThCG+ERvOwNz1cC+9
ukLR+oSu4GIw/boNGvIniOt0QXGBXj3G8MEEkzthQsv8s68RLijcb0J8bj6N
u5cBZdzK6WyFs0Nv3lr43g7k1kZvvr2RwIKoCkxCKX9v4hkAB06OZy0wSXqz
hZtcocBsanTVjSZhIs9gxfilbCwsNmuNu97ztRrtSTy8qwqaQsl6Ueb0LiDh
2t2gyhLERXVerKCusM7BeWvAVt+ubefzhgOOdrmCocSJdCf4n2vorldWHm/0
2JsTLfsXSE6hB/31pfjNiAdwTbaCac0Gl/oPe4wGjMqcj8slPgE/fqK711yl
6x2r3PzrUJW1fdutqNtZSwQnVTDoOOwmMPzmxVIjCmedKGFMxadXvU8Xtb7z
VrWgxnrzACIiQn8DaPYEjzEUSoQRYPTsTUL9O8BM8Cf6Qo2c/ahIEKo/ghZU
UJLmp3PVoTTnR9MHJ5emXPmQeW+1dqtoIo204ywwUeOclcQ+3Bf8Yt0VDgrz
pJGwkRQQE6YMe5OGcqyV7OU/E0yBmu0Pi7KVcQ7WIob748UJUPLGianMd3qA
+60/bqcL4FBdf5rImF8GDSRcRZhTq+RldWpitQvRHTzNbR7hQIc+fp3Ri7RD
Gi9ur/c0CP3AtjbcAEZo3aKzvWJU9UXSPVyGhHOBGWZIpDNGLEROIGQwflrB
jdvEF/97Udon1l4i+WKdfNL6rhbkC3p46C666Fn8qiono8TR7bTTr5UK2yTQ
ULNY1lTkVk3Ka7+SOZzw8IYfnh3uAPmtqQ9UunLUGxeghrhab3KxC5r0RSj7
Hazpyi24SKObLB0AngGgiTQg4Rd32oEqpoz0ZVRvhiFe90Y4BmvoQOFtFbit
ULhdq971r+ld5KohXY4SPydlhjM6+h59GALDHwEY3y3gWRaXAO5EHFCjRGyz
UTJH7pwn+dSD2Fln0bWpMBpEpRlPbLWc1bQvBCh12UlMR0nS8iIBp6uKuou/
3nsfky4BBZAbBc9eJpGO+sPQKsS0mnElbXKhbIUsnGkHg6VYcelg6v5GL9ft
b3RVZabJ9s+uZnd6TiKb4vLACH2+D+F0csXXXdWF9Bfq6k995z08StfakhRK
bBt2bUs/7gtitZeMB8dRQAXQgBueV9yRGbfrhrP1BO3h0lsuEbH6Diif230X
y7GN7vgr2C3emus7sJeAoYyzpe4IdqmUU1K9FypBoXj31TO5AKDrpSCHJYT6
h0S9oCKgKLWxKHhAVkNJouVE+QGEprJtKDjzR/Oi2NfLvG8RsPmwqsOWr3ix
BFw5vGNa2JZr23evMVWEVeAGD+RTVa2njLu1VKhZkpabRMdvl9/LdHvOtCwF
8FLGzpYeThhX1sFj0qIP+uw7/WhUtxXq4fAP2XxZ7c5k48YMBcPq2VM7k+P8
gATIEyTyC+Y/ZI89hi+E7RIC/cf8q3/X6sxFssJ7T39bOVTUFWyZ1QmYZLr6
hfhaONIMGwlPC+QZkZL1VkMO6dASc3ifxB0YQPX7Cjq7aU/FiXGW38uYMcTg
HqmI4/urcUWZoBDJYAkhWl9+WE9HoMz7HeIKYzBHIt101UoFyzRJx/qIUxFU
Nn5eaj3UyAIll09P3kmRB1JxrN313NhCusjS+k69UgaaOiUw57O0ezqhBSNc
3/kFBPgbzq2d/WCST2biiL+ixlb/s11DoFlLLqTma/axdFijXsE3tWhe7NDu
LlSkfDh2yLOf/yzOxneVtfO5VgH4rVoyasGEnVTP7OWHjuHvpSZsfHOEhScX
F0vy4NPY+X1G4YemMLLQm4G6wmoKwId5nYHFGVwrUZAFil5uIFHnwHKvwTAq
XBBPiXHKh+TPMmah3mgJdxhhLHAdTmWVylDC1gcjMtJWz3Fvpme7jzKVEKyr
8QxIAmynjtlHYylvIJ1fh8ioONgpk+TWRb92hCz6vkntUO1xiv3siOsDjzZ4
DpPjbob8zct36QADaKDRe5SpySrwsnOBv3kJ+KURBRz1POHT2IlXChHJbtP4
4qOZSshJgEw8+bOJZz6sTYbj2ryDSAEbuN2Gp2JrNe5Mn76gDE9Gtji+2Rag
iTfHX0M55fnGbX63KbccpvSS0YSq+xNO6RLfcivARyuZN3E01WyNCKFyIBT1
hRN7lFKKYQOfl+alXM25ubkRit2fzKVGu+td+sSG55BQnHLFGV5ZNgTTvvsa
fvnRZXnw1zPuLpxOsvSG86Mxx0VqSKx8+h/04qZAagKNjFgWGfJHBXGjxjFN
OUyE+9SGNpkQEvrsawNfLj7bxJmfTTLdNpPe9FV4+x/U+MNf6bzRf6qfxOIy
noEltCn4l3ClA3LCs8au9+xhwxH0GP9osWKaqm+QhSIoyegUTUr3O0Kh19G3
FaH5Xl5Q/1Qa+uZKgx2JBzvVnky64PRFZ8R55bCVzV+roumq7+R3LDz2vRZG
yJGt2CWloStGPiX5Boo/tOiMv3lcSpvkXW0KJIejEpRASLcWB0TZdBR3hqCF
ZvoiDi44+HWKgL6tGp6muCgZPghpcazS196EDaje3la8SVIQL682GBqg1dpe
iiePmixd24FZ1xbwJTWLki/ehrOl+ajV8T7PYpvHmfr1L9n8sl285iOtixbj
Q0VQBQ8LYf+4eG6L8I1l5X36dcnmPdhoQ2GT0g7SCWeqAl1mbTAZXHfaJtnx
OVT9b7waKeVNFE26XmFWMUzsMiM4ECP0BvXZLClUSMuPLPPL/GVLRePLZa2D
a+COv+1yz7EfJQHaVLcL2MgZ7u9r9scnTxtbjW3GjTPYKs4HXdOmiDpiuB5B
lJy7JKgXjmV1mC4cglR0qQDR8pR25qLuh1/pyzHBbWde4E7cXtbODb0OSjOs
3EfK8VmSRlbqffbD96SwbbfxU++oy5EUsmeR8vpdXlZM0sS++FccGod7lwdk
LxE2Ej/zSkmVZgwkJukineAjpfcVI88OfiMlkVth4pZxYchktfCso7nl/K0r
aM1e0aa2ulXSmnMulyAW/augcaE/ss5hSHXEqgBw78PGdr9RjC7SmwNdGm9t
BRTqUYDdht1etAAmno0KyPEqVrOIOT5PGKZmP02tp48F30eyZqWNAofuj6PH
0wQtt1u0vfaZTY7YZCGRfu/5k/2t4PGHD9F/nvlxPjt56jXBf25u8ItY5qBm
+RVHsxVkpwtrTLstHBPhyyxBSIJTi2tllk5frg3Wigk6Cu8Gu9G//9gomZvk
A/PfEVAPowFM5jcOMBAJjDImdDwCSUCKuhUj06NCEEqzZEacANJi9gD0IwUH
h8fqt0FTKpoGJ+FGtzOWkRZK27peMBMSN0hUPaf+Z6NWnPxvXGKc4HRgJf2A
dRbuwpN8Mdu8UDSajQ+oZqbgiuh0AyJlCYVFWRoTS53Rps7F0gBiB++QOW1b
jkDvgDiDhNoqy0omdgtl8EKaQGQpjaitom6/gEUxFndAhftemv9lDSj2Iuh4
AxzUjvqXQQX1UYm2TqAtDQUrouVruV2HMCbF6m8Gt1c+BlkZ5TQlVePDiiWI
RuYMqMeKdUK2fVbqCbB+a3ZfkmkVZ30WU5UmNGJ1nFGRm0cgfEe5IMzfHc9Y
1dMgx5fR/+MpbqpQEuZNbE+Py/pXW+HKMhLtz2Gg1gAEIV0kqJGZQ57tl9VC
uE4qmA3tnkOtAXdQLTmxGxzlfoRZdjzoF/7N+cZihvBd54M61zL53nL9EHVu
WZFAa2QkNJeRttW7pPrHY7cK8k0tkR/8uIpBNnD9pyUq/QNcOYECRnnNTxx4
Hb9X2hu/1NBJzHV70WXoqQ5Xs6eHHtPMlDSmB54UCWEefwWMGYMHomxznemR
eDBs3hIEmNIfj7TFE81SyU05+iV7Km2ufd/cjAdaf2zNl9f1kGPcWgSDZNbi
hn3G5ASuxSDWez4iL+BZfLDoT8B6bdl1FdoXn2ohyV13M26lvrwX3ZAGbxE0
87XCfkKpvVvZSzohPJPZSH/nXV+3bg1PhTLyK8aHz978LKIrAGYM7kKawpuW
iQ+9BgrEF8kXUCFvI9AwJ2ZTo5zcccGiOfGEXRF2aR8DeAjful6fpK6AA6hc
ko87W9bX2RZi+3wXSZXZVH6mFc5U5OfJKxowd/PtXMLdanN9suVhL4UG223u
0/Ko0P7WTbnP2BKO649YzF/MMIWJOQ31S4pv7TSRW4mKvpoHbqsxdBHQdPdI
EP4NUSEjcIDKMcNFjQ2YWyc1E/G8M9nkKjw5QBxkBZEKG6lOlW2exHqWygcX
ZX1yMfBXbxbBsgEipnt4gfhdZZ2TQG0IYO2ohsdCHwyApP/ICK3yQVl6eMMb
3fNtUYxiam4d5yhZjHXyIrldU/iiAPJ1VGnW1r4Sj2k4y2SlxiVm55JuksJV
AP1/gToRHMf55R9fgNbfqftofDuy9deZwlae69KWaJQ6odSPpOoelX8DEEk0
s5YUX60N5jQrfo4M3JWamvZbV6RlO4oFeZXxyOuc6heAdZJMYp2hqFi91M8F
jquY83hkTbdGFB0kOMg6d3vEZEXHOgT/UitFxLQZNU+63tpj9ITodshyyOLF
z6dw7VYH06FjoalA20w0FruKaLwSWjQ+s8GFnDfLP1kZm+MZAiY0Yniu7llV
3Ga/rzQMiUxCacMfy1zO0pRxegQ2b/+8Xo4Kg2XlDgg61R1bPADzt4PVlMDF
Tl1bibYhrl2x4xERv+Gv8y3/EKBmoWJcDYvc4qWZRYsZhGj/RRXONVIUB3bp
1LWSbTmrfZDIiyYD4vjOaICzG4yagvSuFHdIQNoabuONTEPo7/Ud6xGxgtzi
Hb/l7Uu+q/bcoz937jGAY7Oll1osQMhReJbsBpyKAXmYoKcEsVrxflKsVtYU
NthFvHrogvKDDPkT2gp4yweygKraHbWm9CHGJE0RmIwhLDHQZIimM11tndqr
hUF2ULgV7l2AETDIQBKyA4W1uA+bN8NOliEzKdfGPAA2fGnvRiTd+j8cJI8Y
cDCY8Sp+5tyjzAG2TEB5tg1fsnlEnzaY/M7YNL5oCClpWMTSBmwDe1e+NtSF
39ExVPBwpjcL6jC01o6ZKRub4FI8vKpd5fkwITob5BDkea9Mb4zwdBhc0zYR
H/7ODK1wOm5R+yKhWWlz+gRASkmdqmOK4wF0uH0zEb+MPcAqCh0z4Ypr3Zl0
Y9yJJd3+xvQVX95rKDfcN5RIb/VhvnyCHKJBOzRweos/sMMhvNAfegtZnSLi
/FltZJOXNMIoB4WJwEI0m6tAJ7LdSMUu09h04C7sHcZQm9AOLMQX+oNZvIXk
EF2SPpZltaiuWkfIVJs90dj/CHnFh1JbWLHp/4CZ2I9VsaXV5CQCQm9thrHa
Xf73euqiS31g9uUqvN/c5A2kif5h0UznEwewdP+oYL8aDxKoq2dm5w37OxO6
ePPyYu2pl3uvMFkaE3wQL30FEJExp5klXZXLTGj6+PEls+Exc0v3yujUPlob
H8zsBqn98bazAmWPtKKem9nmMzIyucJKRp0UKOwiJhrnwmK3VcPVqScYTaXv
7WgyEdcNMD3mGXCuAwzIj1zMjgjypOMUULcgNsMJwB6eeK8wamEfbWeNmAOu
9zoiXoaP49VKLbHytbPFvrTtkM6YhgEvM5JCwJqZQ6JcGkaeliWOswu5149Y
iJ+K3P4e2PHRTDcOfm+cl0y/0ZFndm9IB5Gv33NU+Gcfgj8vQJR904x0ZdbM
UqwMHnE/bu1FXMC/DfFeDVGGMRKy++QwvTtocA20cV1vVmumAtgTWlocMlHN
Yw8ni1KBfKy1kf4wT0/6voCygtm4zgaYz18uzGGqNQW2EwHRLYWZDmmnysSl
1UlJ52M42Iabjx1rPiQpZmiOn7NSV3j92NGhCVCCbBiV2gZSJY4p43kLint3
7Pnl/tq7X1Nvs8jSsppZ9Fa2omq0POwhprrOiGLfFzhiE22z1OTLtggpRiT8
T3iz5oLDGQNEMuZVWj5NJG5CRO966hbAAiXfOHLMN6OBjo1V2edweGlLWQqP
15J5nL79HNGVZlPySFy1ObpeMybwqMF3v/Y5uUkV33pgo3poOs8mXMPTcT9S
sjSY/6SxTm6xQKsWLhp04RjDjTa/O0fhESmykr37P3/aDrMf9QFCKuhRuQGW
B+wPJKyEnaoNHprMO19NVnIm+SsoPR/8cfwJ3AM05uEZXSRRX4KhaprFcWIP
F+1F9XdBxaMpAze6uemf2lW5tg8j74/fpxCd8M/c4bnjhymjsfFm9E/JSAzf
6Zcm8DV3BLcQ3ynuBVPpKwq7/9ACeMTR7dk66n7RAiaw4QwLXfHgMKi4+oYq
aSinbMkqPWmBXUqMMEBp6yZk59aA4EiNG/E8ZyY7GhlR+QeqpGvSejQgOinQ
0XGvIfCYbQ1BbU+W/fEOhZwVuEBdTqILqatMn9E21t0m9udz7UtjmjhyUnaI
Vf5QSt/1znIGS5uJTL4a+V0GZU4wsD9t6mqxG1VqB6ZehP4Z3OHSx9yCLep1
TdeCwcgh7x5U1Ha3XYIFGhzcGrtKV5+W0TM69fghsoGphSGNq9CHZ/pyM117
tynd5P1GOjOgWRa2Qge12ShX4p970Fwv90Z6cnJvL5ZP67x0JnywfbsVIpCZ
Y8tFwlD6VXg7D/ZPOTnjxAhKMTykvRuCis6oA7uGfJ5agDpPZtITsc1u/5J3
NrO3Hs0aJpCFJhaii5Bvh6NI2GbkQ4bMeL6C6bC4fj2aK9lWt2sE8h7OBkWr
n1uFleh9Ch5pEqUJj8UALxdoAfsyXIMpafyn6diVTSXtINBFmr2kmHuad50s
E8L81jF7mEFdqHacbG+kTJ+JN2uCaXEvt6cyzjyXza/du3UJWrjsC1UTt3Et
s9XmLy8aPADUFv9wnGkOeCqgHICQe6TtW27xKG9wyrr+7PXpcfz3MpzUXr03
dFnRq6kVCUpVEpds+DWuc0GRlOw3en2p14bYo2pnXshD+9oTPj6+oCHpeWVh
K7DMw2z1tMryQPAbfDF3XA43MsDKUNudWyVYkiNE6erjtpOg7ycQ+r9U7/re
BqeFEWX0XNN2v5bhj3lxFcGzlv79nnLykhBJiTdainS7EmyACc2po+fh9WkD
gjOfV3mQB8iEc0hiG9GHYPT5MOdp7MME9zhS+wxEimwwm+HOZDCv2gS8B2gD
H+p2RsO8DzZpDcUsUZdFCT6aPM0vPFcq1sbmJLO5MBAG15RxhfXU0JccEId9
r579OSaGoYuSNuQyOEm2pwj0pJJ/ZGpq76EpNMnVdPuhmjXwK5bWqmlzeWZE
iyqVXghe6l8CZRkW/QpD84gezyDS0LaoWJvHbhOMpLaloLKj9JDAEBN7ql80
k7TxexcDB+KYykv7/8TSrQB6wutkdaxkNfh83hvwjCqfokxoM6yR4zVGwOqJ
a4FUvtua5pvCZjcQVI90cTYzuqJwtzqEV5sHWazIb15/2ilpsh10A8w0HBZP
Pc7ugJFvJBZapSV95WOXZVKYN3zb+gE4DxLVgfbky0ONM52TJMNrveqsx3dx
ybx0hT/B5jB2qNL11FvJ8Yzin14nqfok1cJ1YbrjiO8/WPTLBx8Ykfvb8zvN
SAIsDyoVI9d/H2pLYXJFpUTwX0qUTIQQVcSGBMqhIsNV59Mck8ts3SQrrKB4
OPUGqR9JGUKJt2krEbjWcmnGQ4GhYRVQo2FFojWNHkeHT5rQfJyrnjTMY5du
EWm2UiSPAmw9ZSB0N1/0jGm3cO98XOcFD5oxg6j/n7vLYJddlnBeqTSgk0yk
lSvoBvVW4H2lAtxyScrMIx3QXCRE8Zk8/7hPNQSqf8meAGg5PIs8sRw/M3G2
uJBQGfkLQkds/H7R49EWxWWMAcrycCfIyEtP5FcFkreQIXGq1sMHJjzDR1Wf
WlH5SYj4ryeKhSeCn38QOxJBVSS7rTZMqmYMAVKEvV+fHifYIcU8791EQZUZ
eWw441TGSl5YZ2uCDIUERkG89E7Fq3xxxw/iVC+QJcvyYZW7SCY0mP1QJsqA
RY16TnPQIp2DdOGHyyRkFgpZJXbkngigS55tbsPjYAL2GU/ga/0GzvckCEs0
UyEREsd8S/CFDE2CWWhvnIjblZSHEpR2B2rw4Cm24ZLanbzzhWvWPIo5Imoj
LMRx8KFOUHixElSjr4rgK4wroESlN4F38Sm9vJhhSrVnEFoSzUVEkWhD/Rjw
fO2aivfUKTednOjca8l7fZ8dJvZenxb08nI4c6iEbsjFRdgoIOIjkfvAaiwf
m2LBeAJCuiRJeiu5SEjThatg+d9Oyc+7RgBHzuKCggX6utu/cP6fG2u3HLVY
Ibj0dILc2P/Udfd7tezxoqko+DPeax2o5468XSISkD2DDXGf8zJ/PKEt1GJA
PsDuGTIXjl3j3mW7jvUk+EZdsYil/tfmQ5tD3gcXKjP2P9TRCZWhJXQmi+bp
UnK6e3ldI8mI5N+Cb31DoeqBRXgp+H+6EeuQpga+EDJkpkWqCgJgSbHjnBs1
3ODypynXFZArPAJZIZqFz8GSlWif3y1DiiybS5gSO3JC1iu2PINa8vpgj2eS
m/lPxYy8tlaVm2D9evHmogdLcAPMXOZWKuh/g07oITjgE4q6p/Es9B3U/Vo0
XpCUwaoc2kkrqshuE9qLRSWcuKluq6dXoyDchCsUxph8XrzMZgvnyYyVZdId
nB9XSt8HxmKH8kjl3cKq1EPGZ8j6xwn9GEQFhRwm2/PIMTC5VGqpYCeFwBi4
l7p/9fPO01PeBIqCB28RvbEkXbAbkIydn2mrYPIlHx/BAwthfdcPee1Kg6SY
L2LYMwuw+saHa5tAIf1FyC6NJnFRtIeRTxoGSQy1wCIR+gHzrORsxSs2sZ/I
/m0+SMCWCtz5am2RpUAXY/2BMxreTHdSuAPqCv450FPPV6kf58zGwFst5ov+
px6UTxlfU9ff91L/YMOqdLBPZwps++n3Y6wEnNl9FnVEL+3T8/NGp3lLt6my
ZVN/iERypu4mjtS7xsaSdXmRwEj978A2MO/XU9JE7CBWsPiKq/iAU2tteoyh
nEnWh4CB5ONlGEynom6oFvWfJ/uHEqG6RkGuDVUPDuZyMEZWGcMi5fmpv9Qv
Qxs2/mzeTR7fOcfcXfgu7cIc3ESEwZmNU+2bryqrU+U2WuRq99cuZKOMQn6k
O+iC+bIRkv1WjXWAfgNMG3eS0F1ce6lAZ1ru0VfavY11fs2KR3UZAcnMVHZs
RZAsudknhoZv5DOLETWcq4R5Pbb+rqM57zkHAzklCAbEzOYCVsenLFyrNpVq
+TwYRof1d606pIuqHyzCl5k4m1TwSUWbx9aIBnglo9qUujPLB/Hy8y+7oHED
VG3Gn69Eg4oId5i4Pyk09ugEqrRfFWW70lTusGtzMW1D115PMlvfgPv3ejat
gwqkFO1rYTDqgYym08HkHHMA4owj+omd87YmBFr3UuZF5Z35eyWODDRFiHHT
yM+ifam8X8ULWJmvP5ObMSoCAadvIKa6vrYjF4/2boNU3g==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+Eqewe1RJEsIqHfLjxYTxENISqObAcLvvHcua/ZVAMsTZcAvh2TEEf8luyxXONZd50oX/Nikhp3TE/jdW1uE9wf+ESyJg/+8kefZYA2RtYwbbSV95jMK8rhEh5fJnkcX9Yut3malA88G2TOBTqUqPubeg12rE89AcAkbke4hKx0pDyZUOp+NBE21SN6SYZ18TIcT/+NaihY7Tjt93I3EqLeEyJgm+WfHpaMy8htPKuShBVL+kiPbM2VkBM0AEkaKDV8O4VO8HswANCCrFM2IwvxaL31AxQ4McGyshqu+s/ITMnp/D1dmgwJAxfk7aIfA53UbZJhGH7dm6K1716phPuu1dxg0Ncr/KshsX6r8iZVQLnJ8Cf5l48FOVFTELFaW+n+0pNVNtTU+RN8CBnNa43WxyAarNeWT4EYUNiLW5IhXqXwD/Sts5L2HQoMaYtwgB89v5KAfGpvUCdo704LqKtvrBQcsDmV8qK3+pYfv99t0UMoZui5FOayid/SRo7siaQDCm4C/xKoUeK/jE9/hLDk7DCQ4SitQw4eKBnsIjAB35o/D+rNSnf4FHr+jaXJIpF6o85NGxOjqjpiiPsRtDWcdF1q25C7PhpeQiG8/N2ye18pYRLKy3ZrcMqUyHnBExjVysYT2aRUq3DGLR4r4VEazHEAYF0LDidoyd5cUYsU02Nfv84kWgyITTLpj5+eOolILmUGz4NRjDeV2pgpEd0BUlbaY4VflMNYJPpgD6aAkInlRrAZ3nkfpQ1K135tR2wM8imxF1yZLbz+ZWf8ZhwAV"
`endif