// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
xGH82XCU6WE4WrkwDF6k88THY2mWtLb8wvFthbRhMsCBNwyaWxMLoZVhruoY
MU0iiUd+zWuSptLfuNq405H01j1UFYXgqmYNJA6SjfqOIQk/G8dqeXXKpyNR
d25Sdl5f9R8+jSPartewvRky6cQaOeQxRId2I/uE+rvYWOi5YdaEfi4Zs6dM
4V5HpAPVB/z/ZcDd97IJl8qb4MpjKD4gP6UD8twqLoLa/ZAW+MQiOzMmWiRy
X/RA0O97EjnWoKN/6D2OvVga14E4BFbqkNQebtePHsUbVSXUK+fJE0OP91vX
cDhxEj4mZyMPMvmNkX0oleiwIadzTZpKSQxL10smpQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZiyxnMByXrvKzsoF8q/Oi5HXZt22ddXGlP34ggK01W3m9AHAAq/fwtazMwG2
seFBQHQ5fX7UJJX0V66ESheMnz+ntHIv5Wiyqwao0mlVbZPe/ERiC8TxXqId
3zELkJ01Bi2S6bxy292+K0cysFcAkOHdZ8Fib/gS/IGKUDPHfzlaMS7/WNjF
zyw9VKIl/1WMFwx6jjkirqoAX8LUGij8d4R9m0F5qquAix8b2M4EslGDR8nP
R4klIGwDKyBMTZo7gc9rOAc6OaqDF0h1eHYzRRJEdqyg3f+37pQhZR4wdut5
lf6bzrcw+2xnovQP36yARZfL8Y34nh4MbKu/TJ4SLQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QF3tvkt1lGYcdKSFZbJpAMZP2Aw+PtiR2/b0USzwFeoJV/HxtKsS4qR/jVGm
S7NCeS0VUw4Tac4q50a8GCHNTdlmBZjIb7apH2fef27LCoYLM8cZ5Xb91Yli
lMLHaV1UimuldORiWF1/FMPrLNlnAq9cCRjwI3gCHJmqQc/QowbdP5Sf91nk
byQi+X/2r/QCorUiLGmcFxmUrGxEhqZ8LHq1a8UZLqoxk1I0M2PC/ofn2b/M
olzhLOZ0fMvAmHml3XprRGnumEAEymVyxwSbN7E0HaHwbh+cl96hy7Oqjgw3
fQlBkdnajZnCovJ4FO3c6BvURqxHpkJrc5nOG+2eYA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HpteMyKBqdDvY0cOcS2LEoOBOFSqJ3gHAiigSO85gZZmu5AH74TMEWLy+4WE
PmDV+JBwdV0GCLwLEUDP5FiGWI3RAiVzR6S3l9qRbQeaLOtyae999II5jgLG
/8/kFQOrcdqsiqYQYpkC/Y10rwSv0f3YU2z4TJ3e/JHAb0ICVH1kP60Ita7h
cYB3a92B7uhmLuh3YJkz7LA8EwJsv3OshL6lMk/gpxRKNGJK0FEu8II5C26e
hJQCJdG9dDmJ9RTubWUFVMTUsPsU3QWZfdYmmNMxUY35gTZtqZ6FM17q51c4
JYL36ePSo91Sf5WwUrY8HwTKZzSFDI4wuLRO05MP8w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BITAPk+u3PJxHMzhalMs+FFE9ugPC4SdXCmlQMxQlUGpHdm7gvAa0IXaR0DU
HvFhdH4yvthVUFg8EPhwxN2eLpFGs8b6c9uKuumYwhXhoMOF8fPCO1iSkrcl
Mjzv6PSki3SjWCWGmPpollriUJ2KnrbFGr5yfP6rbeac1ZFnby4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
C+CUG4E0/BGIi3tnBJW/wNdzSPl7iUQq/AFHJyrGTP0sDdRqbXiyK/7iLsxk
mtJS+qa1MdBr+w3ggIUJPI9Li0hiB43Eo6OsYycXZIO1ZyFXX19paYrKshUv
si/7zPPV/b6haTqTF6HsVHAH1324ArRVoHlr4rtY1ky7rg9/HaXPps3vFlA5
8K8Si3TT0y3fGp3uljc6+LMQQEgQzBxFDkWQlCO2YtCwvdOHnzW4mSdP6VkF
QqSjEk/aPLl5lQsxQ63Bx/AqUX0pu7cDglctsev3sfiZp6Hi9bXqo5rt8ZDf
ZE4qm3rl8VEta3dps/3QzgLI6byPv1UJKJzb9alejRdPWrFaPJBZVYPEbr7b
UB2bN1kH3P97O7DQ6OZsJz6fl8gSpUt4TcUlE91cH4qaK7+Y2XuZT7wuTsAc
uLUJ+lhkCVhBqoWHbK8qX2Xf5K8NKMp0Jy3ARLti4CRrtML+KSQFnbzBNb4g
uAlEGG1v9zrHNUtoDpcLy4ou65WS5Xhe


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ipY5FuU9JrIm5rxCynsZYTyVsH6jbG+hFcipATRdS24hqgwmHGhl0VY/9nOR
6aR+gl58SHf5r3enNFyo/x2iIXOMOsnq3m0EY9O5iJkBOCaDgrYcmWPsczPS
yetySD9hBxXYfv2SQ8VivzKNla20GJCrbVWZRItQtjbGiDFjuGE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MvX/WO3LGsIlRaTIY9kasrr5iSHhS1M0d25dxqV/P3nGLLLlxlDmOfM1VhAj
1OLFdjgYalBBfzamyLGIpHnV+uHrGGGkebN2Xypq91MU5MpoQBjukuUPpmEV
J1NO91LXAoY7E61Z+dq3MkhawbPE3PzZWkAnAmsHQZZT5LZsyPs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 15472)
`pragma protect data_block
QkGh8MHmg1SF5zw0xpR/CQl8RQoJShLXJ+bUx1OPpajNi9mIHo5ev9KGFDNO
W33vB/mCJ7XR8iN/bZICtLQ6WmOpQmKaO6VqtvzrW5TPbLztQy0WXC5SnKeY
DHv5rdVW0Ey7RkS6oF8gh9G41zpz4iqMWB0Idrxg1c680P3WQA490/nhKXX/
2h0ltOfDQUkOBtzHcCJDnO/QVISSod2e/cgP7k0h9wG2/7hkpIaReLA9sVcY
DWJ2JbFyXeV00seMcQr0Lm6q71XdAt9Fg6uZ2NnXFCTZnJ4MV0ZR3iTgzm5F
41eUl9tTfMcztxWyTy6Vs6Wox04qjfqiLe+InBQb2TzX6ouMV2PI1II2+xqa
9adbiWQHF2FEb+OHFkFn3jtIKcgUtIIwJeKFW+4ItDRrJX4MQOvqV/yG2niJ
uxPs+kJ56cgr42BLuEPiTyVxvXwgbBf6Fjridf2HjZU4XrlTe+QcQOJYmKOL
zsjWLpcGSc1VMoBqEM0nMYiBnYO+hTxuzPYTq4W0cPkeIemv4l/bh1GeUCwR
JbvPy7uVOOP/CpwuMLs67NdoJE4lSez4qwUCdTpqxV4lmSVCBrgqIGs/cz42
xkNy54USv+UTalNBxfcLnlwAA1WXZJkvPtLfD/ooGY68lxvWBKU+bS8uflVI
3W7Kwb2gOvfKbD2N19Hut8Nj0dmj1uQcrzqVXWL9itm8Bt3UlSWDNNGRwDZ+
ZXIMG3hIRzbv8lOrVkavIc/SQcPbKQXhd87oV2uQrtfJdeepSUCdX7EC3fnm
uipy3DSmriJMPBkoylx2HoC6xjVIruZ0n5AKLvmz/gqiUUbHq6TW5RXMUuBO
RTHfw1bMVAwrAqCXbcKJff9zalvumXpyoXdjSrhHAJhcXe/sKLxfRa7oStM8
KyEQtk1siNGJIcnAMSrZXSBYG94mLIbQu2fSQ6YM9myHjGTMfBRTVhiEAVPm
U/g9XSA0RVa2ePgbJxWFsuDtoRWnFdJrhteouhhbNuGK8A247hnXyPECd/Hx
Cfc4mmuguJPIuRnuxy8cKolJvEpVK5kF9e5wKgx21YjzsxLO3bLJvnSIHYl3
rfQVuG4vJWu8bCATd7Z5tp8+qUM9uy+XYdyCW4wAICMMa21gHNsZolPJRt2g
ptdQ1ht+2Hb+3QTyyHAEA+aQFU4rmg2Lb19Ab1uJaEZE6uOG6XXGKke0snE8
okqO0/DzfkigcJAvNfzValMc6vheG6HRCBT6VcY8g+CBa69KB7fvXovs4gbD
457zvz8VADAKgCtUA3TEpjFbDjr1oYYQbdcHtS1b0HJaKVbsvRBCoBdr+q7X
el2FRdxXk+C83Qct08Qv83nc4VMAKeo85VQwTMgOKD9eL6TV0ShTMELt0YQ9
0OyyoCyH6FbBQEuEC5hf2LBsuAjnbv6jODGbCE5c4UlYSFm6qnzuP+WUiBob
vla9Nod7/JnjDWXyyNuPLcQjWQd7N99JyX7IychVUj4MPc3VpDtA4LoeIycN
IHdCDD79kv2pDV2BQkWlajAka7jZD9BZSFviV1P/4x9QMz8crd3XhFmvwMwy
hAjTSS/RNzr06eeD59Y6skFmUOwE1hWslhNr1EZ6LxxVX3NsqisA5FtQ6O75
XzZMx+JpflYqTx+E4rcq5MMU3rGHbih2bPjzvtQitSK2BOy0xQG8MDjifQkX
aE+PfCcWl5Encg/8v5PoXX1e+0WY8hbUXTWnWZx3q9DL4OHh6SAminJiZxAn
BJ44T/vLImS/2hNcPIGyRnLUsEhyONd2hmKG4Y9qtdMRjpnpzznTmZaOD4Kh
Xeun5+ahwdjq8oTxc7bkiCP+kZXelboUuPdWmdpp0etXSdpZZNEH9u1bqYaP
VueoD3llmkGQ1dC4NfTCopRJ/FKuiwXiDIw4vXPCstkm/TI5YjIfCTQ15uq3
E7gFtLJt/l8/wMxJMckuLRBFBfb/0OO0nBBnTjVGwqN+6pR8mvKFbsJfOQ1O
6Xy91IHPgdxPU6aTBKDzFn2tMGgzD8yv0x060y6GFjevAs9qw1BQIOR1k77F
uD2IBTBbjp0oWJxkbswpOmyByMTtyLFfk3Us86/BYS6Dfg9ZC0/PM6Qmyozc
5goTsiLhos5jOJDGti04PWTTDF2tMNM/N45nN+Gj3dgTKjwihVTr0dULxpXd
4BleHVmzomaLI0V0IRtVKLLp4+8BW4hXBO3IH9WpnwAB7x6Tas9IJQ0gbGqg
poPlFyXbP6uRzz2KHFbM2OVCxmigm/YsMDrmXAi9TyP1jgMnblgjmN6Irlx0
3YTy9QbTk+2Xq332dMrxxNZhkCAcOWCfmms5SWX84ydCn8il0OodHxh7cOLv
1xAVdTQUPIHMnY35KJwci134gkW9wCU/yCLW0ze0XdxaDYqtUf9al+5pTkYk
KjSR/zOQu+CRZe07f0oVrhM8qV5OntsBYlmskJkQ3j7QNejiSXvMEaz/YMrm
rfgJIKTKooiVMBr6EyY2FaXXEPFk7T+6YWA8uNeKO9zcDCylovkUTlCAWHHm
YxaZRQV0xo8jAQNj5T8eMbMWTpBy3W9ipidVSF7Bw/YHoKZ4GuyDqvyr2stn
5bSIoKhItgdYGN4OkI7QqHhEPUxxSXeViQVVYmycqmm5v89pmeLUyvpq7hiZ
fWVs9p8Z9/Izqmz8hG56JIumuqSVOZ0aZhXyzqHIegyD0a2Atq31bGym3If8
9DrBHdJPQYzMv8MIYTLsBcWcnHihNznd9B19WA1aTIW3mEe/26JM+JcR8yiZ
i+clKHpBdXntKUrGCtXtcSbJ+2b7pr/sfjfSm3h/x5KED9zTNmEsbOWcdMoY
9Ut3CpZ4w0tWHdLUlzU0QYn8ZmzLJy04Bbp8NBKqwSqYD/R8wjeV2KDVqGoq
dZweSxo9p9pKJ7xE4wCPXqR2RikgrGEFYEwH1ipuNylGsUw1QgXUE3uBtuYu
AyoIlTOt+L4m8sYxBP6EtU43vAuAec3FyC4OV98kyTau/xvrNzg6/kuMKMxy
5Da9ETa1wJykrWtbzDVPN1j6RY6aCmNsEFw/QMza5ipA4Dp3wYDk0leNem6k
wogWYYn9zJCW6IVI/b7zq1sM3Bk/GVyKAKm/ZIv4oN452HZ3pd6tRoyJcJ15
NH4RLiPHbIIC5SXXcWmJ2OPt0Hw2kFaeZ+9isxzkEHXceCfT/N9JZfCgGf3+
OQqXBuu9U3tJXef7AgWCZH5BjlbtE30uVzmb4HrFEXhJwZlZo/4PCKiX46u0
glH6JtBQgX0Qml67uSGM+9c3FjvB9Pe+2rf2rDe9xIP2F5ozUgLhqtpIFoFg
zeERqNTRH9zPUvugpvJ9myA+T8Ic9BDyVyoByNO126ebQ9TFwRitzP+dZz/5
g/R7nRwvCPtYR5Ni59Lg89GawSw6Xl/QiF4vbFvcUTdXvD2Y6BWeeJOONzIA
PVB1vNidThYlLJ3Jm+DkBALoHPwXr2z2sNPS9RiiwfFU1oOAcY0XBFkkW8dn
MP4hGIVW2ydLb8ijhe6fmEuvppPd2NFnJIQCYhRGsdUta3wMGkIxRu1GKTYW
DdTPaCX+YiTowLVn4Q2PTb7e+hSPlJ6zbaUlnKOUmrl2zNERqcmFaTDnY7or
muQUX3fq0CmBrzxS0CgFEGolyLhMPfr3hG8yq4miIP9ktU6oELgmU360HXCL
Q7eHJNKodLWDkGd+b6V6qHgHsjZm9jmMJXJ+476LJfYgOfJqd4tIxEjIDfh7
kpWY2RpMwyvP3+NL3w7yuXA2gIETyIxBN8ETmbwh66gEpWyut98dJbVmdElN
nmCP9Yy42DpOMeiz7ddvlp4QwCnC6zVFNXvMTfkpNYB9/1QzkGLb3TlXpsv9
GNPI6DvpuzYwSDBPOCYg9t+onIKtc11EvSbXYrd3VLAvUq1JtiQOQpyrPBvP
mth9jdI4GtCo4hazWPnIOTMlfBWucHxIphMe1qg9DQ08ug2lKo6sG/AaC8eL
Gj/yJjHPw0CWlBOJoQfwRrhVMA+sNgFjDsbzEK2N5A4eCReScs3hXUQ804ao
DIXpTtBQhT91gLQhDy7cmN7ndnqECznqSsJjDAwdvI5JABX1XrkfpNZNBmQB
2PZFj1EJ3Rb2bmCOKGXLoW7cungMMiIbpjguLnFaYu9XJHODB3cUjyesxY6e
vIw+/DGdAwe4u39gxcU+CoP4ELsuSk+o4e//EOnJ5rpl1f0xvY27cxr16iA8
vJ7STTvUmvpy5XQBKRXPB/2X4o/h9s7N+XSCDMfJTI2OPHWLAhoUpfINtd5P
P5bYXYTkf46XaMoVnRi5RDmwKxa9b2VaxMAUv2wly5UXBKWL8xTniaIkKIpp
OcIurVM5bef31eCvNTECGJfTWMsBnqpLBPkW4waEGl27Q4umOLw3YsDNZjDq
uXrpsKnIVWRffsEo5jWmGsKyBWsTzSA19iNtXWoPnyT1ImGc4zS1kuM2v8Al
GF9HlnTzIyru0oJQ4ojaQJNytYW72iACwh2pZhLs/1io0BN9bWqhlKhZveiK
IfhCuf4f+GgOkqiwegH1CmXkc0r3lYXm3q9FLZGrtUEfPgBfKOfV1lHVt9QK
tk1Yqvofk2cFYIGZVqqc8F6QrhVF/7fgM01Co54p0pGORBomHuA1b9BJ1So+
nxPeFWhT+y8SDyKI5/uKxMW2jKTsA6+Ru+Q4ocqZz6dJHkHGfgNHzsKZdmMP
IFw8wyi2XebtuzBZmWceuCBzAGXUWwNnyMElaVW3FTADp411oWrG9EDxKO68
h+k904YCndU/A6v0jvq7U8XJvWSgtyt+sD9UYncbpwXGUc5w4hxXjJrgUnUC
AaInFRJIcTMuAmIaZbLBJ/cQUO/sfOvZxMVwUnxuDR2sRxrnrLDyGY1lGeVV
u4mEshvdYWCW6ZKQIUCBsTA/gBS3kHSUXOrtYV+bxeuJwNcb69PCdVxyaMpA
KelmC1YXOT2DqbgPORkini+c05W3XhOUNlyaxMPSD4BmDUHsjoZvVEB7JZ9k
IsH1b2jmSYY6dp1OfNnMiLzsmCzA2iRzF+WfcYEne3VFluCpsZMVUoo+EKkP
5IrW/sgV+w2Z5VKKOmRzB+oaMKRaWNCXuGZFU3hqENwVYb3mOEY4VdjHcu94
bFBiY2S0fO6Ntpo0TzAs5rxEfUu2D3DhT53A8sihcxidW2LQ0rSss53pzGOB
2K7xuj8zaAZVJBlflHk8BSGNbLS62aDnd39S18Yzdrw4FdiEMXmxhJ2b4bul
ukTMG26mImRH7zxWNoCYCjH+sib8QKv5zIt1JpZl1EajX3U9PPYvpX4HcPie
CSparocHSWmgkomT0S/rACVCyckGifNjeR6IY6LZE4mLqyAgsK9TN3ka2NHi
p0c4+howkHEyfy4E2Q4tU+b9NH9/HpnY9PbTmeQyQxndfJvRz0SFljNsGkOk
+8rVFxx1MNHuQbt4dpbbtr2JsL2bJ4+k8oYH8wkay0bn2UnqtDFSlNCYZIhc
OM5QiU2pdk+7Y507hHwJJaA/CgkIZzELvCbZhIHYMWlq2XxjR1ODDJcb38gM
Q6b74VKYh64BZDkLk7Eq+Wc99d8IUdWl11+04wF/JqmsecovU83m/we43R1V
sGAomY+h4mHJbk42FooGFsgXysd888Rjp0z6TbngQks/wBgpMwaIfAzkKywL
274EEuZmqb67ZriCnftLqA+2LnqfDKHwpPFT/MFHWktsdTzmXFG0qOFIuZcw
yzQlMv5leHsbw/gHh8gl09mgJo/YCGy+GQdKxaHIYe4/FanYjwHDJQmBzZnD
UUZcI6buYhXqUxI/75VcxEkO4dUeBWZlmTCjhgRMvlOeQuh+PFM2zYjTI7s8
npfUr0cVJVVf+qukD1XnvXfZIN5WYiXPrwsTlRaPcInIapUbKk0GxkNYJGJy
pWP357WK+OnfDAGGIwvSvaDAsdqZQxffKXgLw4sfaO+p8geJ6jTj4kbkX+oh
AddHum+wdCSuDSBcxuH1N92WmgwNh3oYo9sF7OAlxzmivTJTinw66pG+nqnb
Tr65HT33zJ0xw0jNEkag2khUSaMab1insKLotZ+LNUFkILBLF/Xqwr5mfdpg
OA5/eD60S7lJ4L/lGcyk/kzDHT92NC4cspoKblO2FGCERpnbwjHRHfg5f4Y6
CVdJmtSxuFztwkxbPUKn01V0jb5rCzxWZRnalMs7RhrRbgQBV8y6yUIpPsGh
sxwaNtk34AHF94ZTtgN9F8rqUQeAAkKG1Dw7kkiEzl3d/9LgKxaMcfvQfG40
VEo7R0V7mcizg6tMoz1imUcIrz7AnN9HcUUPDaG7wi8N//hL4Td12TJ2couK
4QPajMtASAJ8kZIFF82nUFQSLwodq0jEfxutQj76bxBH2oYswGmrTVLaP9/1
6DJp1gilThWtfuMGgIFV8L/DGqGS9DQQTpy/2nlwCyASfdLh2d5TyUuqRwPU
jN7LFPfmIs1h53vqDzUcj3xoutxzW+/sXYgx1sloAke4yKendXI1Rnb9T+JA
btRVrvKjytOJI8c9kW1l12bAP1b72LGq0sWQd7RI+UPdWTyhu4isnYuzueDV
7B84oIXShzBF4A4tUrQyHFA4WMgA9j2NWD7fNhvYfAXRmLKbonW9fM5mrEV+
Qne+AWV8D3Fs9EdGu7VkfF5Mt9jSmBAo5tMbJM8L85Dfm9cFfSnfJrf+057l
5a6RV0UjFcPHg7IiiKofl6YmDa1aLa7ccjvjUE3zXFq2RafHEA1UHtd0o7Zy
P8YKCCuVdEXOf72CnMDnQUwmiLkB8pkMM2t3IEc28x9uRzwcW5QRY4paOfUj
TzkIRQtYZ+GMiNwoZsL62zWyIF1ZyQBfAqdM6twJCZBtdyabjz6O/GOm6LzP
2ToTI0EPH7f8inCjVPp0NUIIlMwnRHu/qeWgzvj6YIBastH/yPS3jlwvDg4y
t0N67UX+Wzo+dGP53nZWBTDgdWy02KCSib3uaixmfUba808O0ekjL0AvvCwU
yB20yu/IgTpC6te7+KHafpKuAktVX4PDuZgAceG/Fr4BKW+CcvbJQ/e4Jjs2
qUT3zGJihvn/D+CqNp1IfWb8yKLAPPNv8BEtiiiggZKy2ogl3N3yCEFmkgGW
YQAyBR7fNyCAtLNTPbW9pBINxeG9io8E2HNRtxAQh3bOYqCB6eXX5hfV9t5F
gkMHnseDZIJo0D1j0onbxeTZwYrxjC9W2o5aUoeKIt50o2UYAjnqsiBe/of/
/t+kQDNM7/MjeMd7LZIet1+K+ho8Ims6izGxozyZAxJU4Gs+T5QMqIKIfBMJ
EcSZG3iO773qKBtJUOGqMTeRZDHxJrcLVNZTFcd80oAFbwe3h9R3sjOJSZcN
4liGma7VPSFhPErC9WKYbMoh1YZE4Z99U4M7RtgPzsq5KGfi1ftjuf1H7uoZ
ZggH8NLUVj4Jt3xpn1ElgNRECybQ/hCuxSA7+tGalVFu2C51XPHztdU55hHW
6/zq8M3CwaJflS6dHOJbsd/oq1peAAtSIvCRKxgQo0EwbL/FWsIa/OJgjUG2
WzkQB7YWNMM8JAMm+ZX+7VNyYLK4aM1alqrrmLJDPEvc9ltEPpQty2Zw8+bV
midt/f6YGed5KTBtXlw7gVXFza5chB1xDAvgmIajTaQ5/W4RY/HWpbCN9xPT
oQ+i4WGRKSLsWjSon3V3298aXkMONza9B7w5QZt2Z4BPxLupmv9ICNbHf8J8
rLED9YcbNhekCjc9BAF9bu1iOAN8oyY00wU9bLrz3VdfoybNcUvwG8WyzGXZ
lUTKQwnNS5zzKgv+r5u7TRA9MAViUtZNASnRuj9std6FuRsC6o1lnwTklVBB
JSjoHl1eGD44r7bHVXOjib109EibAXeXgjwK/4CDwbkM6iTpgRrTKDAry2TT
bAlRnmP1y78Zmgidbvvp7SbGCpAW9fB1oK6J58EAAJMPqPyj610N2Na3GtII
4gabCf6V8fBf1/J3MuqAQd3+0aSO7qhnkw33Sd+oCP6ZQHX+4yzRnLW3LxdI
o0O8JaynVRxzd2gUbEj7Qvrl9J12eo2yv4Q9f1bVtN7ejHS87ttcCjcjQAx/
8DzGkCDJL8jRbs3PknDrE0Can6WynJHOarWdB4Oy3B/WUhEDhyKfNXxc99oB
qI835T7Y2RVizCaqmp6uNeUKKpxkv11HYYq016nmK36NgtNgeE8QaWEjCaNk
qQxOAS6avSOq0DffY1JYHDmSERqeIrTcu6mdGGG4uwopypikSeqEAKaYEjbm
zqXckYPwCmF2kJsB8qWUzH35iyrALWjRxJCsGRVioUnyGYNf04TXKy/uot5o
b/4boFlIZVO8cLh75vXNIRpgIANANmrDO7KU8xvgi6zUgNDySiM1H46iOWuS
vJ0/s3CyBDZSmvN2RPXVkzekWBqz3kmHuCtsNY+9bJlGYnng1SrG5axZUUsw
7/v4Vws9gGh1V9tCwL/4kwTWGaEVOsVWV+HU78MZoBKYXvguN2h5q7t05zRH
9v50qrEh7t+zb/caidULrXhbXFynwehtBUwZLx7ZYkNmkIlz4T+H7efr9rr5
MJ1lAbyebU0TYF28T3s3++tTTy47p4wY5SJLY0c1Gen/E9IUfLduX1iY2Tct
PvEbRZ34f5ePK6uO5MImCoHW6v44pz5oA3KdfurIR3vUsbAvf6mZO/1Um8u7
L22hLyIV6nJCcFclr7FrHouU0tq68c91jGWNyi4mifSy21/mkUeXONZjJb20
X6+Ywn82eutFNsMY0jb3Xh2UBNAtPS8zZkh9+tuILK68sDI6piFJKWuUpcKP
HKuXmxVc7Vus00bMr3nk7jJPVjr4A2aEG40FJNWGDbQGMdNEbLyHvygzQ/Ep
AOJSgpOT0ULVzW5vScpvhLCSMtTJS55bVR40A9R2+39H2QDLTJPtVgxnG38F
rfpAhIAXIl7zrNf9o/zKRgrK4mbGC7WYT09+OsIAG2OxVGlVXMnhc0zRJMJs
PRta6aTceZCfjKh97OSAZjkTTN6/2IjXQqe16xUVOsYKb31ef4rpN7OpkiNJ
wcLP5riqxXAQ7D/7qxK2uUhr6CepM4162n0d2RmDGoqqmKOrG0bxLQFZqVU1
c7RE5rYwEG1j94CB56w6Kyvk3o7ywZOL+0T88Y3zWMtEqtz+7rOtsdqeo6Vj
eijIaiH0OgTuxJVEQFvo6L4wzc8MAu0sfKXjeY0goPozV6fRck9l2vVSsifU
VbLhz5H45S8HlkJbiktVQ6o3SksrXFvNtWXcMH+jLY8G1aO5dVZh5+mFxxDr
1NjXpaZpUsvmkviyti07ucfhJbxl41fYoO3S3fDsBgjRtRREWp49tkaThvNv
llDlpjOGU5YOYwFxGbkd2lyjxUf977x98PNXdOiDZz0X/acExLdAESFq7CBQ
bu/kwLtETX88BTgg1Rc0PA8tbEPdByrnCyE4lKE0z5wgKCtCXdcBZtKDAfS6
96Z0m6ttED5R09MIi4GNXoG4GhioModMPF8VE+Q1QQpuX3gJrJSgzOfZJQAr
MiNE22jJrwUyBp0hwEpeJIFi/R/DUS2a1Mexqx0nyXS9MNR4fIpMdBn1Ys7j
vI6T+ONjGcd6evTkd/XfAKAAlTZvV93I0e49qDrgjto5mYr3tK0ZbFbkva6S
nxfVLNXP6RqAP++jhDiPg71bokW9rN2mKoOhZNZghhFZSkzvBPOFdMzRo2Qi
dEmSQc+RwSjzM/sLVYeW5XlA+L7GwqmYC4LFoeHIcdTj78/b6uJOwYUt71mQ
0HNBQf8YlOiCUcXUcKJfTxK2b1u75dWhZigVSF0tiubTDUe4bAGIsKJlDV3Z
sdZMOS53eXuHX5g2UyzCHwlZfKoljWs64a3tbhbsZH+8CDytkV8jjuFOveT8
XURkgJVm9sQZH6ZPHEgBXAjEJZN+XPmfq9lppxoJ8ADHphbwJgnlKqDNg2KX
hdSP5Ujr0zDM94PBfwTMNOObPqiTlTIauPE0e191ogN/Ly213nUE/NOeZPB/
xQLTk7lg0UxF12BQH3UmKTI/iDtXvoTZkW8E8TGlsVasuYHpCN/CqpEoIcul
vM0gujOzB6WLTpDEyFu2fazJznl/82/6mraFMWwftKd4ka5/vznhyTK6yGAc
6wjtlVb8cad6Ixw1wdUm+e41pGjPMs9zCtZIS5eETuDie2XtPCl8hOq9Sw76
3o6xP/lLUxXEDiNxM9p96s28IR48xZ6vk5TUh62hmXIYd6HKrtUz3y+4VCDc
FYOYBqnSJ91SWEwzRdb1sYi7PtbExY9x8tXk9BUK/oD7cbhVKbxBcL+5bRKV
iT4x9IIpjIPsjry29j2u+uYtcEcP9wJLUVlQLB/DVMlInbVpcpdaj6p5CyhU
j0PiiekAmiRUSChbmZvzJruge8ISI/PMPjZy5QpHVqmBL4A8KAWfI7Pi3CGw
VEyXePLUkTk+j29W9G5S46Mmx3qqB0Ox30Kv20LYL4fWc7X5/tJuGFUSo/FX
fZBBkzD4zY5SepKkerW9yH0WKhyKS8un2bdOVApXAQTZB6d+MyPKIGifFlSa
JJEmnUFYhoI0OwMD1+h3hfpvYmymNGS0trE9CSJKJ+lGDEmHr7O4ogYxjCus
/DCZpodaf5qw/2k7WXq+5aidJOXErjtQKi4ZRICYikMurqCevjLa5tniMQVb
ZADzfLoe3Ph4TLQpS5X3pZF9FAcHKQd+jYT8/iTRR4aWxWathineKdcEErFs
MV+705L3IaGyn4NcTsl/NbglXsiq2F0WwPbZsy5FYONSJH0mQPxzzJ0JBycV
Mg88+SxrXhhaLMz8v8QxfyVxIqaU9mfREjbD/sbTjveCO6wm6WUznzcKwHIT
Sanq1lcZ2kbDvQwVdx6QN/R0f6K+3ZzDG/XroP/8l+5iB/fwERzUA+DVZjuW
0XXC1W9CSpZzIQ286Ca1fZV7OpLvOD9TEPgfgqcnumnX3HvPv4pFXAtR+WT+
y0mg8hc5vO86RT6MqkWgmogW7O4cAXfBjiCaRen/fNm2Dee1QwAJjnUEJnfN
pQIaFQERYq3QJNrfzLptTxXjWgEdn0RRFhHSWSFkkxVB8k4l57tCz2bi12M0
bi/63WPC45BnE7w30qkYt25RW5X+2o45mjJgH7mhmt+ty8AREBDN/WLfma3o
HtBCUpkyX5uu2UN3VheVac43/+fbjywgg2w0WC6BRr7h/xHqSiu8Mn39T2G3
zzyp5BkJIJNX0X1cYD360xk3Jx8EpT+npokM4g2oezXaarUotQGHOOlKpa87
1hrZrtAAXDhGhWelarRmPgMlQ2KRl4aPpKkMScxaLcLromH3uWl6Uh3FRLCc
CxgZRERdM97TEYmNsqAgcSEnlFbMmh+ot1qI92gWxvILYA3jEFyimA8PbaZK
8BQDeGOrdwZdH29iM+SP3ziypQD8mKPv8dE0EWNQVhmB6HY/J3UctsVnt/xp
oOViWFQ4qMh8rKU+KE8NGbeJz/dPjuGOU75gZnQjHsj+zIORwiKuQIfYHSLv
1YCWOvp3issJ+nAKJX5T8o7s3LdHunkR6DzJaXS/eG9o2S0N9hRcPuHKiSw1
DiH317aT2LCOw8CQn9PwbJZAbadI5nK0kWaRlck/zdABhzx88i1a80zKjoAO
O6jVlryzpmZIi8OhkuIHrOuRzXXky2rfezfGCQ/2mtB9wUTFGcwq1Ltmoz8M
gJ1sNpW3ompbyFgF6VZLMluhRpGFLHdl1CfKMiPErn/fvXCDYxsiGxR7tXqN
aAK2x+MBCAzxNihRhBlOFXjkflIVwcK/FPDvq6nd1IOeGL9gXxzZc8QX6XWz
G4SVKkuuHtCnTD4Ieufr4EqrU2jyrmcEEzXq8b1QNeGLeHYKHhatrrryOZw3
XtlEPaX8jEzR7X1oKr/e8trsq9/PoV53FDnPuLbrgu4D65aCfcBgC+HPifWh
iwRgqeN3RIzteyXyUzQWqbu8yo/BRPi7DVu/vuoL3LzISIfLOGQCgjA+m8gP
Rk+O7sdPzecC2UafHBA2PQFiafDl04JUTYopZCGXcHmvKMjScQQKOZx+sv5/
IQgpRLlB+gvZmiYJzddwH2h6/+xvBXdx9YWKvOvglPE1s9nTpKhyA3WxZ2gV
9aJup1R0Bvu31hu+9hxzfnUB7WLg05yY429WmlZzyr427BvjXpsqTuA3g4AH
NjMyJ2322+xDWC8dOK5juSEJFWIuGD//6Ef2lmi3Ejfk7kym9Ig9kNeYd71+
urllY6J8/gQe+Zod5jzPeQoPC0NEZub8j0W2+v/aBnsq/OcFQv+GB+O955g/
bZhvQ8cKwF+a61xA+Do6VZOmVvoI0jEqMs9RBM8VpqElcMm3Rml0Wz9RmzTS
xCmNSdPdWY5/8WRyKb94KwG+nAEMU/4OSLaik52im1vs38WDqiZrO9pbPdz9
k3aO44YKvCv2XiEYthovOj6YXdhneE1iAl2Fl265xn/fPMLYGZ1wdtWdzn50
/yLxP/7DJxgoerweYqaycbjAOzrNeKBhz1AcYzMwyDYh+B8UCSOkfdTunL7j
nrSZBvtJ7i+FNx9uLsDFS9NecUzcWOZNuHDNTIv3dj8MMsKvdrC6bmU5Hu+j
R9dYVKE4GseryZ4qozmaO7kX3Iko6RtaHp+c9XJQBxu1l3X24RcM2K/mNH7d
PshGhPA5D5GkiGbHDLLjAdTp5+NpBb2mpScDudffpi/zKnPyLviN4FpHc4dC
SDTtER/ZO3Mouu8j/ISLLuhaQ7opTm8FxlbumEUdtx9FM0mCKxgllbr5EuDz
LL+wC2/VF+VkY68wn06Ju97OK2QN09zQIrhXQEk3G0TjsE9bhx3rUVegn/J+
GsZUIJPLMCavF1mKPyigoVrK4NfvitgV20L3FA/erKeuxF+90Snupx/xqRZN
Vp4rwXYFGzky6/XKB46U1VTqNbNXwfIGH246rmHed3BQAt9I4a4MOYH1c9sd
UCnpzOdzZZuA6vNF9xvYDD9nQ8swhsNdwh+dXUX6oB2GzrMdelsGdRQq+Nwm
xysQIacOywrv4jn8BPF5wA8o+/r0XbpjHgXSAKY5dqRH5Oo3cF7zYdbzM/CZ
EkFl5b0AZwQTUkI2uFJwGjCjVLmRSKUOEalxTcjiAS2xUzbqIoHiiUdKvpn4
I5pUukHXBceOeK6bUNt/t+xHpI9/AhpBB1qRAZbFqmbgy74fFNYmkdK6MPyp
ce7Ut+EjZ7xEZ4Oax0x0F4IjpWORTu0spYmNUH5RIkiSJol22FkaVK54jeAG
haiRQMrKjbCfsWjkjlfetUUHUS0UcU2sr8sULhr88jlQj0BBr+w7cBvq3cPK
7gvXahNTBIGF9266ozzM6gwd49wWey7TjVugEs5cemZC717NIMvbW68hO8m7
XCm6JIKbzhc6oZLEAV2+ItBGBOiVihAeqPndoYxcOLqEBewuuAndso3+3kXi
kM3XfZ+TKyu/AW2zFaKZONaOZbMAaC5BAa/4nezW0hnbkUKAHqYPWQRs5Glm
SLoNR/9pN4eesLeS2LBbltXyYQpX+e4F0aLTZGjf0wvfIXd+8HcCaQDwTrAV
bFmtXmjOlULkN7wsQAPLkf2x0Alq9R5kLRisnSfSLccihno6+OOt2YLAOs1F
xJQ+7PQiFuf5iaE3hBm+6hcaHqeirvCQMBzFLm9keVC5yccwBtwFIMlfljZo
GqEG2ujfcnA1+mNo9VIgTlaQ2q/SMlVrfUGKT0Uy6eU/e+abKntw/ysA2mFM
+J2gFfsHmazSAtk25IVHnV0tL+h/DL0kXu1xGdwT48zKMNqA6cCJ+kBqsEj0
rUoHBBLpnU9pITAPLheUEROixJPaoYZxm6l3a0ods70y1yqeJ/5Qs12cWKtc
pNv8EJMrQ60f4bl9QeTdi9FE3quTorqZQDlD4MaXkLKRr+V81i8masAfSpsi
Ca6eJLfT7Mor262bfOVc30FNVHaNcV/0MPAc1MBysUztIYGlrmI3kB2zHidF
Ga3QEKVpQ+nh878w1mdc/+/ggtogTfz8bC9efEIJRLBlOxzVQR4m4vrSleoU
HUxAboIpPPTl6qKDjbDiMOZifLdyZYZKJTo3lXBvgN1CffYHc59NAHpPjTl4
BXOr0FNFANmxmFdiVjFfyPvgJiT4bZWwGT3TGOkg/fZaapAgaQKdfNJd+jJR
vVcl8ADW/sbNQe66EOAz8yoSVXGA9Jqpo9dzGVT9LJnK2qrEbEbnAgfOQsZf
DRw4qKymfdebunW7I2Yser6hMVbqcBEpTnKZqI1hyVypoh+jmkftfRZI2jFd
Hnb4/ps+F3f3Lj/PaCSDZg6W+tu9TP1pCGqJ8Wv7h+ekknp33/hYoSznr83T
aAo/3HNuQ0b/8zhGCrkd4bxb99+0N3bqXW7zg7jW6mzp090KO8QFeRo47oC9
+m1DXCtp7etfxP/tA/24LUtiBAfZHM/ygRR5Dk6ze51IQACCk59S78C40L5p
Rp1UZICxRtxivIFbgiz1y0smex9CmrcVp7F2Qbspg9gqmaIpPYKbhZNgYReb
JUIkQjhgoYQa7n58EKhMtnlu3THFTn0mEqtan3J1pq/3iucesi6U3Q3J0rTF
XEcG8uJaMrMIIRLw7TweQY0y4SR9uB7kO5KtbmglqKOMez1lgQeRtF+RHK1Y
axbR4R8KU5jlejFwuQHYt5M/x2pD3oTAz5Nw6PANYG8my8yPb7/nhKeJAK3+
FIxU7jX1ghE36cRBRt0zDb/xhdn9NK6AimtkXcYUW40C+SPMyagJoe4NuEZE
h64/SQi6rPShAziwgpWAx913XSv2DDHpVAaDYd8AqEoS1rVlcOWHyHsDCR1A
d/uJAG4Iw8jWRN05VMkzPSXF1hi34rsbkxA6+kywqbU8fTKjsn7D/SPFfn4Q
eu0D2HNsooSFksuuoeZLTEXu5ChD60p0AJqi6vy5JaRpjaVKaQGJH7M5InYp
WJUnq/9sMyeW/5KC5yMkpnTiB+9ZXs3cIAfmpUmbFY4b+bryecEbGh7bjZTi
l2EqafhiRgVRlR9Vt7lVrIFu/OaVNSFD9Y/rkjhG/FEgbsHsgbgJKkEMVPDN
yp19hhh9Z+yhlirXFQTw/fkimUsyh6nA0jspjqJ9bRhNqMwTvTalbNVffDSj
/oXBOl1ErPxaAja9bfSt7x9MOuMnku1n6XlM59gp7tC1xSWc3IYUF+2hdaoC
PLDisC+jbnMjNiHsDrK/RszIRygytBzV6WjTvcrlraI/VroAM9My5Xyo7uVX
ya5Hy+iTJoBJZB3HNj9as2Ct3KIcAZtAzo7bfJseTLtw3uZXvQiWg8EX0oOu
qhhOQxvanRBQV44H92CYraLzarFZG+15sMs1I1UgP5K5CIZif9TLwDrj98FJ
p/ggxVsBD/7gxD02J6OKIVlX318/PxdtDtz96KCbZOAIuwAg/rN26pKAZxZ8
oF6qeMxozsXoPI12ri7Bfy/UZ/1AHd4V93fPWqm5QcqAZetw/l2Y9h5IWOtO
kjEj45P9QqyzVaGdCjDs0kq2+nGip6DOsdKE7SqxrorS8SOIaMONzG/tdwAS
OkWL18xcd/xFxg2ITmMu1C48zy2oMXEo6S4C+zwjskpncbBDupLActIoJIhD
8MMaWv61mSDDJUUgf+npb60RMkFZIoVkqetz1dT2frzN99oUqDG3elajbZo8
R5Rjq9/KcvoTM5xuOdZfjCuVzKDecsFHVYy+i0saQXAkT2iwjqb2KD7PGvAH
4FVyr86oYhDAK/qJxvvurC3KIF/TKpOCZUqXH2M6ameTh66nm0DAoBXH0J7E
lIl3asAKQtixsvGCj0YlunfZBlpn+WMxdGrDzRL+Rjn9WCwsXgKap6X9qUEf
ejHD3fY1zrG3TrFp0Wa7UWLcZkShRhf82c4dhwbLFkMTTkgGS4WzuKY9kago
RkAQi50dAsXiX47P1mm0y6jIGKqA5j7A7l3/zvonaT1GCuxUSq24fAASmpNs
QAKSwIJb3qt8OeC6p9NO8MoNqE6sTopgLTJ8oFDkYhJRjZKriddxm4JNaEm8
YuOKom0uDz943iQu4vJKryo1d1Gm2C5ezrCJSD3L2iePHZM+yWuiyQqfBrmg
CWQmnvw+enCnQR7f+vr9/Wg/rqTiva0obFWXjKrvyEGcZCx1zrd2VjgygN/e
1AMPZjVohoNwHhJFh4kBPrHD+Xvk5su9beggLeWrQoWKbtaQcljpjqV3yuAx
YdVmOoZzsaYOyLvn5xDtuBrK+rxGE/tBP12OuhQPYZkjzfoKn3B4qXdC/zha
7NnYihKUZtP1aJtCq0C4dlhQ+E65PTJmr9R6wc7qL3eIEY4nImHNfnJQlo/I
2RBzP8wN5eiUuKqopgqbOjrTk2/SNb4L0ty40TstdO4o6zKKB530om5RiW2G
Ck96aHEez1KF+c6SuxxHZwPJlmhwx5gSW0/cFcYO+f00uhVndHUNG9rBzQYl
owVVdQu9EwgIdrGLmQDqVHUzesetoyMJ3Th8P9+7l19RjrZHPUp3hVBUJqiB
2A2WBF+BKBdJDjqvIt7TTG/KHSjU1hauQOk4tKwE10PYn/jhdOy37ylh8p7e
ycQJ9Ii9TLk6SkhCnaE9N1LO5g915VBh/gwuQHM5fgE7wwuI8tIJ4ZVhwmGw
meY+oZL4DkbKHgDoMwu9loQxdtcEgBNnB8C7elKAfjORMjAWVovaxQ0FEC1R
DE8F128S0krZ56YSLFgUNfqogE93At9zRxphUatmqPAczkgQNy+TQ6YzSZre
c4G7MTU7osDcYN4qhmBMbG+buTTp0dz9/VME3nivHu2foHnc1AB+k7spv6T9
RJm8G9wq2B8WEsypOTR5vW8PsOm/bdCfXyPCplKVyczLlQZqxSGejZj/r9HS
y4B7tlsnpPjlrxhd437m2DFmo10L9mocnNjwl3m1W7MpNnbCkM31Sh/Q73kT
ez7UPB4KShfWU7BWVx068SqP74CreH42Rzc4HwwJQprkSdlg2WtPIWwxR95k
6y3Jv1BLTSAlXcEJ0tcho55vH5POE0ilmrKexM3/9LscDJAmyPpAmOzskjyw
OmFp61R3U1/BZVOsPKEXU7D8ScS2eRzvzM8MjUlZIktelBLyRbD9XlcnRcky
Av4AP86ldJKceHyV57SM8pN+1YpA79Ci9YZI/K6r4awt7cxN/kNJQNbHETPw
GpM+2mjt5DlA6ZYmBjHKe4P8HAYUikmKCH/UpnXVbZgt4EBV79EW+W7uB6oh
a7Y/2BE72B7tIp7kPC6WovVflTaPsDNzNBNJ5YMbbPzsRplzWITXY+YZ69qT
Kiv9CR2veHx6MYvq7NOKLve9KoKf9t7Qav7SJfvLIERe/NiDkkdKBBqYanZO
b6Lu+Vyss8t/CAQUh5Fek/cdTbGGbQuDV6NvS/lIIL7y8/p+tNgiXq3NW2DY
DKckcr3ZB/JyHZSIauFe1CUkYpcpqSiXZfojjWvYUIxa2dPie0zlnxH7e/YR
+a0VkXr2baxDpfa5ce6wTj4xD0zxskcOKz31kcRTv4aZ29xDP5OfpJOr4JAK
BYYSsTe1NiPb4CSV2Q3Lbbd5nHJNyxsvtkIptLvM1g2+81ZGeo2nMCKVSVS9
4BnsZkfUdLD+Gisaodbquw7CDKoIbTYEC4bDVYn//FDFaeQ6RJiVT6IRHuyx
pR2QofW3YAoI8YP2RatgQD6xLNuVHlokD6P/CVYMV2sYASrw4Tx7Gsrv39ok
2p1TadTqUikRhhQnOX+Q+O+qPWdlu/TEHUX0knpImF4sMa+fpj/u9+FQPnMW
eilFjqn6pGbFEscsvDxikw0vUUFJ23royIyciLtifd36nYC06VRgOdXIkHPm
tZiKJQBme3bRDalepu75hiIER9loeJ6OXKVtXPnEjtcA2NUywZsOLriLPLzy
ay1f6M29MQFjfa32xa4xkvzxgoH3W6EkgLicJZ4EdJzvJr45fuMEpT/B6dey
2soixIHbW1FS1sC7IR6p5sjK+HCTORppkqygPZ01pZ/BbaiPD4cuUlRVtSLH
VJz0Hef3D+K3Umy46SRghrhqrl/bIY3uZXQwP812t4vpjCe/Wl0uLuVvsek8
2HDmNduvLPK4GET6hko4zAWHlM46MEmrI1s/Mpy7xek/j0eAfr+drhfA1f1x
qXBauHGwiNYUtLmidTUpypfGcGbE17nhDuXDUhihYHwZDx+4iJOPoUNm2PfL
hXU/J7iu90WwkPSCI2c0TY3M/mzKKcYEbNXNwJTFKELPYVHZfhc6DiItrWdx
gpdnNl/junMrboGQcRYnHClWbbfkc2AiB05rL0EMVKHq6e7djGLRwFuXEuIr
Xt6y1d7tZVG9pmU6TWJjefqErWrpOyj1Hwdq9bmOLajrQKZQWGVrq54VFU4k
+/58aRoUNY+nlQ2UACAJLj/kgUYOEMmsCVnEJ8rHtk19Z351QMHwxS63HNYB
wyFi0GiHSPxx2OGP8jqlkAUElmAPWGqevwxWwBtWtmxevxuSuq21tEIH+3Dc
4cz8pvy9ffJfgHJ0l/XFGHZI8taC5YiqCwY5utBrKOfQiUqH0sSp6ekBu+eC
XJxkZ6VQl2BDRNbQvXVz2R7x961liULR3YkXjvZ3EfmX5K6LQamGvXq63UOm
UwXqbavqJOW6/5tQ3Vvh6+s7K9gbJaPCU61vd0p/YwUQB2kj9nyTUXOd78ZL
DuBGx6XfYuMbNONmG7WhK9o1i/WDbnVDUePtPa/ZcPtEEdY8/9LwaeP5girB
uAdkLAltkGLX19B2/8bG8r4qauCtj8Nh3qh4l5IKhf775rugy/Tkqu/x2WA4
k0qO4bi02MhlWUl3mwtMp9PqKPscy1IC3wu4oIUwv1M9Oio5qruQNDEJka5v
PIDXoN7yb9DVqmvCDhb2ihCurUw/Nc6u2EA9apEHyskpf6RygSWsQyeTPLPS
3pcbcYeyjAiJjnRM8Yy+0pSqiUPmwKIyaqEOgAH/gUJ7l5tIAmO6/Wlt8V7n
EhRUMKrv7WTCBQQk8mAC7vHVgKK2DuexBqFencvXiDGtC9eOvNHl7Vu7Wz16
Yo76fwxqxwIkS71ljTKxtrgCfmszSzuyQHqV8uUKOw25Gj6I5KB/QW9xs9tR
xloKaSDoaUsPXF0Axgb84XB1IUrbcLyZDlMpGBwUxKSItJdYatkC/tICOXbh
/SuSAwO19PMnlk4d9z2l2bgGcOpCRO0yrUmeus4fAzGEURG08m4mL6adwGfC
oiz+SSXSS5GjGI6rGN6kRt4UUvxXWj23/Jp495dltA4hSljQAUjW+2uyc1x/
DijVIlzUf2bUsNEse92K/HAE+XVew3rH+OIRbEt3DYA0oeyx5DAN946XfTwC
8tF1TSlNjv/ovUlwPK15Dd0t6vn4wMAwAVoyu5r6XoXhmOE1zgHQQGLXbR8b
B+KUIYDo3vV1tjxVM4aLWvjVo35y51iGAKfDWhluENgqG8M6nXFzM+/3mrly
hNZpQLEMQQf9VJV04sa84S/iHrRqnpdNImKQ6AU9CU5KWx7bCC4Ca7vuzBOp
Xi3Xu7mZHpmvW3LM0q3fKsEjtX4PfhL6+AJyKq/uUIcEKcnX2LxhdG4To9dB
gQPLwgmZR6zYSZHxImujJj9GKxlxSst8VSV4Gn1q5hoEvRNKWiF5pMD1Bs76
FxRVkoWljE+CP4JC4AaCnUhYkLJlBKeOAB9VQ/maQpr5wfU9cPcAtMFRQkcD
E+VgWxSx6Pii8u/WmzipBGw+6IMbm/aIMQBc4BIPV9O8FdtjlKFdk+CO+T0d
7OTZkdmly9IUxrAArosvTkynhDw/YEVQi57DmQAIAz04BXrnomiB2ebdpGgp
Cnebvp7GJ0pYJ/sNzOcCC/7zJDrUGafB+pOmF8U1A3UoKhlATAnnAvJLciNb
VU9kmzeyWStqIxbi4WG5ebsV4unTb1lbBeVFe7CqAzIwtaIV6RiRUkodYKuZ
s1OJkZSgOhPOzH9fFOh7HblsnpQ6YzNEjmEEp90hjNApvfDQN96LCJmirYjz
2J5wzGe9tNEixGNPCi8Jmjj7u/7gknq54qjXjLgFivlx7rZMf7xpmnBRwZjV
7RilpPQw5Cv2gqJ1Ge/zORMKIHWz0Im+wN+m2Iyhxr4ibBWO/O+GG29Enx3g
BBWZD9tySL08xsQATmWeiBBQz3ubTFcfHxzqCaR6XuftydbkjNxWdozUSceu
1h5XCuAXUh6Zi/wTmP+dTyxz/fLPZjnaHS7l6fXvoN2byRIWAVyUCvhvr4Hs
FHwuvr3KlEmVR7CcLvOY2xqvBOKdf+Vzli+ghcdA4yr2RMy9TU8uCEZ2PRLA
VvEemfLmlka9v5Uo3euN6sa3K1rlKPS1+qheXph4CRXrqL3RN7Cd2LHuJ6eE
J6+lyMPjeIiwYohAAdPou7fjsCxOpL7ErvDRzZhco9INBoSZj4dGz7IbRDyq
uQnX1r4WIPJIS6PbmfJ3Juv4RSBlb8LDGmbn5nr/FHJI6phclF/DintGwMGi
BHwtoizB5fxCW5rcSbrEtpy8LabLkT08U1keUkXKgoPMYd0hsY/PETBI8yao
a597RnlBf6PLg3XyEiHL9KT+1+KUt3HMdZPrGL01YsxxPQTCHV9oh/RecU9D
3tC1hi5fO2UYvnqi55CAWMa4O7hap5ipWDV07gk7CmgRaLNINidZp1Ud2c/M
m0hH+N+hXHJV2D/kYsVzsBre/u4EeqxNz+ysmGNzbhvV4G2PqQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzfs9CAantPxn8QLgwVjYh9pjcEFtv4mkgQ9AJxTO1xQ93Tjf8GTnW+aUUkSPEutGjxoOki9c1g2jv7l2TGgNyiG/jeuxHVcaGm4GdWFiFetsyuOhkox8/F7ZvrxF1oEjLq2xjMxsUwQdPE3T4iteFHwvvsbGMM17UA52yNxTR2DrXIjeVcucYlHmTuKFdJB+oDl9wJYIrXlXgmXzmPxfbd/MiDlV3zPkMdJ55TcUvXlrt6DbpiPXks4QnlKJYbJPC2LjtV68MB7NA1WifB3c6nGNW7dU5AJWvrfL9DSivia8JhPmmc5EAsXJE9HBD9oqFlz8oc1S7KNwpxNHrxeC/K1IS+PsgtQl8ye/6GNupO74TGjHPPGWkCziA4nBaEnbQy7K3qUWDtDsR46hUfbpi0Y0afJlhsaPJACh6uA+HK1u7G6YBBXN0SKElOzgvY5WYY9+x5zV9lM0TZH13L4iK+u13T1PhU7oGbpzD6SH1WMekZJ/XxmgLRi6s3L2qu1rOZYh4Eyve/s8kOVeWv0tsZwswly61hkKWyiBwHajaIVBXCOp5Cda8j15lNwZw9YcsXN64TjkhVrwH0x7u2HjSQyKYq3DmJNcXeYfEv8m8Z5l0C70xVayE1mDJD29stKiJJUSQz/eEVlDh0CPYySKf+eOAH7RVrdK43z2VPFdTwPKVyEv+8PqtIbL2U07cjmK8KREtp4INWEHRi9GnC/e4G+x81xYw19j2rj1RkgsSvgrmO+3+Crf9fxPphE5s/ry+zBovG+8l0cWNgH/ybBoFs/"
`endif