// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
F7I4IufMf4Iqq/Wml9mrrhA+7gXt748h9VWPIaQ9qC8SyG0TCwjnQTNvahwH
qRbuDC2d5HpmN289G42b9KjBhOdFEF8+czdanOh9RBodiWiqhzQZ8Zn+dS2D
GUL/NVV46z4U1to/sl5+AX7NACjoUPi8OwSObdOFgkGp+bo5U96ST9UKQPWq
79ReyjVd+b0SxXBfkipoOtRUUMmXnqOVF3OStrd4Ggj9yKvqec4xtxfms5Y0
CiVE1VesqKRW6TEgw/Tpib5t3KTNiq0rXKeIeObyJ3WraLse2rfWVswydUo6
BPZ+8R9U7MgdjHZGoTw5aVSI+M/crU4OfxFft2E2Pg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
S1TYq0Rj7DlQDEJLbB3svyzikGnqF/9UPqAAswgkss3lK5/mHEahKgY2Ymi3
tvs2w3b75H0GAjzugrE4fWizLI2iZfHxcot/Ieh3Y46W9pNK8xbxID/tkQKE
S3Nwsqe6q8hkl6HWlyUSszB+YE3N4Fhvgd19ZMWWIeE6XuaNNV4Te2dgVf14
RnIa6dNYOLnBXhMacegAxa2OoV0qV4xu7gI3LMHnXYcuYU9zvOQpEVrbzpHG
j7ifV0/DPXSDRf5PqPGbRiq3UYE9V1wlCCsjKlI/N6z8EPRpfQG2/ctSUyoU
lJIU5FIS8rYvyGklZKQ2P6oCfDucdXqQn40SR2PGMg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qSZI6px7HMbfjdccJEHnaavWS2pFhW5uIHiZBPF3ImuzFILJNuVzQmiHd+A7
U0SeF7aTj9XcnBdz3r4Nn01OkpbPN67MygIH3ppWB5HKpvwZS/rERilCsoyX
6aBonxzmQaKcyS/L343Jik2Rzl46O2c1AobTxAOa6lsdIZXDLlqUGyuhB06T
gOSebFFdCZ9wDk6WIC65o00BPWm6mruFJItg3fwEv6r94Gk63qjuEUSNdSkl
5BiheRm+vlTkVJs05i8/qy+/ViU+Uhk7N4Tx9Bas7P66gvDRCfqqrS9wtz23
6N/zwj8qew+WPCxHn1GzC/6uz/L21Rb8wsHk3lfCkQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kFR3Lf3LJx2DlHO4ozr5Imzlcc+2mNvM/POgSpdED1skFK08xS244COUg84p
SOrE27tPqKbS+SprbtB9RLRbtjT//v4TPp45hrcQCbgGjSlk1YeFgvsORyr+
sY6WdbKC/dsRSkh3l8eqZwsjL5oOfALPQuRbvspJ19ns6X3BBTB/vOkHD4Rt
ACkKLU3Jy7lt/LCIm+p7rt2+Di7Y/Xj63fTJwNRa4RFkzdg4rK2KEwvgddk5
pl+lYb0IrZABM3F8fi5U6Ts+iTEqAXusuyO7prIuZWQ6oucdEobwjbOUaqh4
jwqqpRu6p841Xuot8IM0NtmjpznsMYR39XhFW0APdQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DVwEGS/5QKlQkcUL+X/mzCH7SFy66EGUaSTVAjUHgMAgs7dZhgu8+UyRlh6z
of/7ViDPBa5IfIvFDzgAD3HmHcxxFi4Q2n3+5X8IEs2BTQcLVv3bdtkg3qyR
21X74NbC6a1YD5dXl4d0rpa6GoyIGpRn1EFWUVNV6dBp3AnFHco=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
hJclXrgxTyEtE+uUliG2viL1S9nyTwe8r5Z+z97xO47TrZ0tAFLE/xbraIlA
zkbVxLUCenHXx6eZH7TJhONuI5pmSol6gtgUyvkoV4s/iQQD2CXuK25MVaVY
828KO3htJs9Ct8KL9/gjAbGKI+S40MCzs3yKlOiVgR2U1EwDuefUZiPF84HC
8uE9wbDxp4YKjBiCwB5d1KiEHMVgomaThXiKJY8EpMvmZ753eYXB5mJ73PJM
avtmW5Av4NMMSIjAymi/cFy9KPxLGb66JUGVr24xKJ8NQHdDJKMkPrK8p7tX
eXblG2GlVaMMVR63B8biuCUVEJF79WvtQiwM/x1n21Z7l1roHfreu7taYu+C
2bxt7kNNO/fMe0+KhyiJcsSSF9aFdbA0qMgcxr4QcMYS2Mu3XT5O9pb5o9bF
GTK+ZZkhmkNijr8lshUbPNcxKoI4YNf7J1S2LXntj3ED7NpxsYntN+4L6EYp
IPpObYQFX/Cn6TE1wxQzEvdUN3M6i4eq


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gBin//jf/qrN7mOeqOg4EEmVUuB0EAPzMUC8FIDXmxx7651mJx82wJSNuWnW
16Gc5WsmOrFQVxpnIGNNceJt9v+ck7XseODBhdc5xftztgZPNleFgRe7KjGt
JlfISlsEebsQr58EDqVAGU12FN9CNFUI/jBDZeQUlQtM6huAp4w=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FDSa3giK+NcmSxT7ghbs4214OnXK9DrMAM4vr0Ol3xi2NMziIV1waAyQ9OjD
0j/fhC7hC+EWGVgak/qGXy+J71MsF/wiXkj7+lfhgS9VjMDY7IcSwhJMWl7A
OasseJBixGTY/BdUjrcghMKELiy9xAPfD5Sg2OjzRMCzi22QkHs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 34800)
`pragma protect data_block
DhPLGMBt1WsDWKS+wk940tv0Sh2n44gsr3g+ewwfFGuXPWyeQhLR4XD7x7tF
PvZovNzUGcG/x4W9A0r5Y3Y6EbJzCXLUQPb4Bf0uIa/DUSiEx8/FT3KJYWwS
R6BSourg+41wtTaHhF9zqW/vr7mLD7TjhKJzD8pzARPev3g0P/Td4pCfJ877
P1zBoiMO6Au9HVWV2OrSfA80wmSwNr3M/eZr0tY6KA219YEzTyo5wfV8K2q+
WBarGF3FbL2+tKgJnMmuuDghGQGAB7PuVtUaEKvd0hsEGCjqmXFI6y6GyewW
JWvAgkp0rUdGwHhnWx2Lq9mJb2w/5SN2+f99W6xBG7wBPYxN1CttLPjSPtjR
JldAiFPHb13fa8AnHSx77fN65z9AbAn9XMm3C3WRlEhxZLsTmiqtBSHaP6Th
As/J85O1ORxjJslDjB+CdpP9qbkm/lmnQTA0oDy5tUvBVQ9p7fjlkXb/Cwo0
4QP3TXJzUHPmZF4IV/5LZ8ggBhUW/v+yxt5B4+sUDX5oidGuFawFhdQ0trCQ
0r56fGwvQ0MP0EmV3J6perbCC7vSe3Jahq/+KXIsS3478Uc5OGsMBMtCO3Ma
gSoM7G5BrCyGZP5Y+CkdwiLn+Zex7WB/1IYZpbufkUD4RXjBpeNohBwDaolh
CXSioT9M1pxYoYAoio6PSqLsWfi4BfkPQ6crxGHQ7wmp7DTiaZv9PgShWC97
qAQ8hLSap+y6H5DvrBBl9OxJN6jQ1mIL/Jt91DQQ6Kfgrlpz7QdGOy/7D2Ry
lNCoCHtDqoRX1m3E1ZIUyvb73HagWJZFzoS+IgBcCpb26C/C+m5XZPj1JvS5
OXHsRImWjsKTCnqmyzcIMypa4KfOiOpXgY9GtkubmVq1R7SnGptv67sXSjPY
s958WO+JsOpM1RQ9pacfxBUQ4PKb9PnZIP2UAeGI8Cf9ruBHKQRdfpzYbjYQ
tgWgR1Oas4PhiRciNi6jOxC5qUKlcfu9010L8oz6IAHRs3yPd5d/KoOhKMHo
0w+Wr47rcDzRljUGVD8vTERcFYh8hptVTrvIxuph6PlRFiGThk+9UeDjShO0
Un/oyIsOOurNx1nUHo0yeeOF2ri61iJ2gI2+V1mh7agNfQDs6a7uOgqZy6H7
OZ7Jc3HbIVCDEAzdvxMrQVZLZD/Ha6IWaZlhg8gOAth44DdEb5OqqJNB+9i2
hvn1t0sq2xDjfaX9nHioAbrd9u+n3vUQorw0zmdBpbzzSBSpcNO4CGKAF8LU
VBblthDvsPuLlQ1l1wRjV0PBjE71jos8qWdlQnfXg+npUTKi7cDgh5fPPWc0
yFui+tFLdUZaFMObD22ODCK1VIcY42S4cb5Qs7wfGGvKaX6w5w4iMiDajt7J
onx0k22ty8ntPcL7sx2Alerp1pL+tl+5eSWwQyrfeIQLAPc3G4T4qZF46NBT
IgcTwes1gZReU29FnNJHFNeQX5nKL8G8JTsmep0jz8xjECHANmzA5HxKqjFV
UG5dzgslJYagpxSZeB7+lkEoZ7IlNf793L8osMsCEJvT8Qat0YT9mnKVcf95
kw7dMkdjQwt9qPBpOB5+7AhjJDzBXx1uFhqiHKZZKk/NH9v6AdLh8YhMay8x
VNl7pv02a7sifYnsZBa4lAtz6T1t+z5L3Z9Xi2G0EdFaUBRlLVZBmpFVaLw1
1Ery2ABDV6gvw33/p/gWvAQjZ0eWNrVnFDpv3UQB29l3BPwZ+b9M+VACcs8I
NKcEyDZe9u74xJ6V8VGI40Grx+0CbrIMB5KbwYerB7tIEVEWCQsgj1Hm84zl
3xqVIA6N6A96y5L/xvMu/oJuyxiQkxCrlBDFAySVpX6vOGsDGNa2Og1d0nvC
cbmXsw5K53Ztir+fisHp16DpT8G0JABi7v5UR9dj1gNRNLhxdh87u8D5NcxX
9qcUF184iiGp/KXskpzQ0nHN5nvk+SgmA9TAPzhqhGzRr3PJ8fLY6Za8ZfMI
iGI7dwOe/s3fikujdTgeqfH3GAqVXbRV3v2wtyw+Fh/hHzYAfvB0whocV/Hz
vInsYoiRDDRRkQOQ0wFrA6q7vMizSZu+gF3Nnlq64XSnQ65uIw8xw5Ihih+1
8OmsNGZLIC3sY/R5+ksxpuYta0KWdebK8CVgZ7zWmoyFjuT/v6Eguq3++GSu
qvzFAzAA6Ah34+FvSrxBJQMhU5Q4lfD/Ue+c1u1K764tKCv6o0tR/9XkQN6u
Rro9/eO17e8zjxVcnb8oRGDf9RWzZz2r5nSezY8smhYYk/4skpzXk6mTa3pq
wUS5h1VA4N+QWeu71c1Uow7YbdmIn/sOwxKkgC4VP/w2kjvJ9n2QMZ0XlP3o
PTG7oMtQ8r82pfxido+2gZ00zs+9j+BaiRgg1GXjPAroFwaRgAOxUTAsi5dj
yNdurQMf4sRk01UTnPpS51srfbyvLtUJxeVXlRQfK5pYKY78wVYmuZbfhxm9
5QcJ3gR9IQS0IWnxvVVqCRgOyNp5fggRHd6ZYD/BktuwxkdARHpU5tmrzAPX
YUnZqkFk3KQe8mM4gDrXeuMYnSoD2+hJSqn8nJQlf/dKla+muRxFgybY++7l
b2T6OHkWiH4+bsHMfrj6bGnVG12SIbOrtFtBICxfKBGRFYvQMUAR86PX1/UP
jU76UJugtnMX5L7Ys+NeVS0MwYHKaTANASDi5ZAt8Dod7ydaK/+84jOj/iVd
f58OdjbsFWZpTFo1ZFtEmpvODy8xiQ/4+tpaco30UYWVDxcqL2/6mgQm2A7K
MT6LESzDO6eISy+cpYFr7CPnyksIIzwxTDF11ISpbuiWkBIokkKrfp+ltC8T
eDd+tMZIL4qpeNaiqYC8CIzyJpajEj3yuhC0GdhekoU3N4pS97usFpHv28LL
XyaWmp6spLmw5pOuRcWORrCp27Bz+Z88gjGggYWU8XKLPrSVU7gPTCHDzYaq
ILTsEemTaEO2rIFBWJ3YFePlR06jrFkOuR31JWrgnJjtJzicOMZqQ33wYBpH
+JOd2F042adtVnF0IaiLITMx4SByO39wCHlX3lDnHHZuRtYrBzrDnTmJY9ur
meZGaRW7EzJWcOhg8Rfz9bNEsHg5sXYqBOle7nARrr1yGAU77hjogWWdHjSt
W3hmTApFZpGv4x7vaFef9b937zJLWI//qcH28UZQm1r1dxi3rtdDWuXXRGas
xsDDiLkDv5pGmucpPn7mqF4aMThXYQjL01wdhvK3knfKdW+hNdq2V2gxrW6i
xJYy1E1Rbbrx9ejFCyYpwQwtvFWU3238H7GYJ7sZ5/SnE7hTwd+GCL3EEaha
IXxwxdA3V7ZoO9Ph1NPWu/YcCyzjGIViGatd/RdXaJFKpLc31kvrZnDM/oLZ
8ADoJivbawIjDUfD9CZAeJfdveY8LiIxjKbBPEdNtAkxK/xLdZYKYCsrXY2c
KF2FMqzrTFzxPITLvD/z81UMyESY/stV2bhahBH93/4Pxbk5xNfUVPOjRmYb
u5kPt+PjFXGRB8BLl0r263CTRALE5K+F+XAAr7hLjk12/DGzAEVsi6DSQsNz
58OGFoR07erVisvjNiHxFMgqwqflmOybvFl/Rvmz66dgVZAIV2WD5q+GYQYL
7eLJKnbwJkFzwBucGTUYwGGGvs5GrO3h3cip6W3YkV/zVclBeV1x8D8D/XiE
DX+igIWKuSnhik7rBKNg5WCMr1PimKdDJoJKirbXpBb496pw5raGUZrGlnPn
VzqDERJqUyIb4ysU8k/EKGYzdb+UGcXQ09abUuyFiDGNkHou4JPOTvVw1Ymi
QGuBoMCKT6pfE37n1F8sAFGOdCmCe6e3aMUUP5+ctcBpkhDf1Dc/qWwwHeo7
+sOYky4JDoNjxAsB029bw8DDA4jdP74++GdfKwm2x6Pg6JkM+4F3SfXctBNp
vjqux50CHJH46qdiPMDAiFMosoe7ILvnzykjO/f6WiKDNl3zcDSeGl5wJ8Ey
wZxPxzwaRe9bFJACPqpnd8Es0TntwTxy37cRrbKVxICWUyl9dhTlEQLscCcA
IMhr7CBEZI/GWryzp49OoKseZkcGndCg4lExA1oQyPEExcP+K+bujX9bGRP1
QrAfFzqDPHhXTd7UjFQttZqLWrEurwYWtR7aNO4zFp/1vcnKAXfR80GGao6K
qzxGqnriim6F2f9StMIu5APf3Lu1lheYOWOX1vQc5X+DgeMvnOJGZ983aQp/
04x/xrKJnY/NOi7z2z0RWCTfGsLgjLR6G4SESYxY85SKY7z93AfMugmHm7VO
8tASETfbUaKGHzyRv9Cl6rcLjRxXgiL6UDFlYc1xqjpuXU0yePTbBpthJlEr
ksptqJnGWsBOMPACC7Dk/XhqFYYlSkBmotkP6kZIqbHLx/JmTv097sFVHgCx
4HqnqwVnkT6Js0D0Kb6nO57o520NeLeq2+4Uivr+J1NsX1gXnRhjhJRgt0yk
FBiOQYTqxtPNKKBytGYBmJaqh1Xvf2xE9qIoMtb53DVsCmJfL2hloqnaqT0o
6f5/a5pa35MlqHq2BwKjzU3mG9C7OQp5muF/ZgxVxhS0QYzfrs1MgH/DbakZ
5HKaz8EuEs2rkjzkU6fKdMRn66wj2bKQ1DP3m2b6YVxgmd9dolb+Bf0H9KSj
VrIO50+VNB9MsPOcNebOsxbCP5x/VCxJsZe9UjOXhZuqWZ6aCN4rKS2WxOqk
zMl8Wn+Wr+EQzyMipm19IGMc8UESRPr7UL2nwiIuK5H9Ulaff3UjEyCEhMPO
yOGbo9uwIIViYV2AYJ8jL4nxyKOfO5sI5N0vMj597S13AllPLMcUyJlL4gRP
8559sAsP7ZEVMvYtX1PmnNC4jN410Xzvhvde6/YY9SyhSqRWXXkbmt52pQXw
dHE3wBFDwXxQXvqjdnnUkwePdg/pfC/H7X2g5RZ/QalhfCTTy2klhxJx3EJ+
oo7Kl28CXK5utNzDecnB2PVDFpOB66QDUf4xpEwjsjx/m5dL0TPSMR9k0q4M
DrPd7fSD4vfL53N+jz6/W8TVI6mJlE1hZdzTzcYA4yoT2CKk5p9+btTU7xV+
jNRPnE/Tri2r1ywGq3+Qca5iGGu5+VmMsE7A7WNo9CQ1eD2k12C3pED/EGjA
yepqmfsb972kSgC/L6spaeCYLtq36itf6dWdRcqxshdRxM4Fd658zZrsTlkJ
lau8pKQy1aSukRQ7+taL8j8Gjq0ZLDa7RoDQ5c+g3YVaBoSDE4OmuZTpkq9N
eEXItRt5Y+SuNpyHnkPYgauvvztvYSs5Y7zIOxDqi9xmI0SFwdJS0Nzq23UT
YJ1O8G/+zBSQcgAy3kjmn84xAtnH8TjG9qjC3DZ4QkkrnHyD4xifHDsqXQoH
4DEsCOxQPzvWf6iK2SmmV4waWXv2PpDNR2IRrraNPZoQJiCu/FVYj4DSOe4f
DGGzzCtVR/o42G7j0SnvL6k/SxFxIFSkf9GGi2WD0wMTBcUdzaaDGwfSJihz
ShQ4mMYTtsBgR7b/wbSdJsRMkjq5WiSM7Z71UTkn3T2quNELOi9ffLeAVUo1
zNr8f5sO4AYYHck61n55cPZ09h9Rif6FOpoWAKiAeVzY2kaoNZNjjsWBVGWE
5Rct997ASFuK+WnAo/FwdZYFSB4TpYej3UwzfMafTw5RbSUybR7I27xvxf0H
xiIy8nDgZ6jBCpqgbKe0vqqBn6LA+KxeDvCOsp792O5QPYdkldwPrxRdz1cf
L4mZ4v1XmAZRYQevW4MlM/t0WeevXeMbzKWjJAGPt30kPu7kZNuAsbZ9uIGe
8c0LtinPt96i17ucD8nFakDObNw0AYqVKia4BGjCUxB/K5XGh63FE22pKsbp
ekw7nOIcesCh0QbG4OkoBM9uR0EClPTumXMBW9yrEZE1VbHaNFParITHB00U
Mn0Q5LKV8yPMYJNxZa8sfPo/o8MZqJTG+uNyNdcbmHrnM4aAnn2kRvZZpqGN
Bo7gqdiFh2xNE4QUJMC0Ry0l0JXIt0tMfbYAZORyiwUvW1Gjh13nu66Bw63E
/gUFWiDiW7wg+YOkPjvtd33iiMYBsrPGj7M0CNepi4+5og62M/aQnGhGQolY
YH0kCZtyDeVQPxaBcKSpYY41lUM4kub8FGpV070YHxz5uhWfwabn10184f2U
QerifWZ+vWWX39P6yQCigTRNiFCa7fgikGWgNpYkcVB2iiAVjDrb+ihKJtyw
B8yFoTzzsuZzdNjIMmEm702aJOzn9I3LIlgSsBsFZ97p4sAe1RAG41eyr+8v
9arnaq5v0+kQ8DstjaisvNEx6a+16XaKxYLbkyGbiDDkvVKDZgFL9oidC7Gr
g+233Y/hOrwXdPV18gJar1b0/E24F9MRNcNPbOy/sV0oLelgH6N9shBBGWCl
QluLpo0DOVEavlZIuGfroYWBU5q6S+OCgmx6reIRkrDOCXshNvgCCKFKyFqQ
HwQtM+e0QwPIq1pqvQMZXQQLPafSH72O8DJhyakl6aSFw8AO6U3HAbL7x+Ah
gVS5APcoQYiwKeMD7LLn8W712/zyKTXXyPnXwXmcXmA0Sllsfm5JewAjhRGk
8SuMyeod3JJyn/hx7A9MvpGi8VA37mQgH8Rw3T0EP+4EmVv8rAX6RnNOZ6yU
NS3kW/TNc0qw2+D24Qz6N+Ldf/jy61zunZWBtlEC2WXCds/pq+4vWLoIAUSr
BSVHLJpqoBIkMtjBhh04T8DLDYi4QFCR/AC9UGYPATjbvfHztrYVUea84l9M
CgilPawWCpv657+o0Krx2IPQWe2SL3C7cxoVW9xhLmkwRSYkinmfVut33Dw2
zuBTCOJcfxqVRhxnIOVu1zxUkRCDSQhYaTEweCG8307SheGvM04tUWTAe+G3
FMdqN3PNuYAqz7Xg4YbFBw0ayc/La4ILcj+2nCnBREW4OKq2Iwz7uH4k3Ewg
/mm/P5JgNvVnzIjdtoZgcf+DyYmvegcu8rkpFnaXUhMmiyv7p1K6a+mBStQo
WtY54IvFkq+a4oZyBhBmEWcp8mjq1dejpEldM6TUBzYjHsBZcUp3kGkxB3dV
YlmoB1vLsSnokcE2j5T7rmL7BRvxoVnEIO1mWnMSnUeUrp1VogHerd5N5aei
Ormt+v1f9cRWl47abMto9MLb1wXUjuYDiqn6u/SpOfaFcTPc+dalC30ripct
Y/4QDmwaYXyFSCg6/zqCWn7mFRKmoTa/prcU+TalyJVtMqwfM2a0wjs4q+q6
TJ64OAQzKz6vMBrJVlufDCa06pMX7d7kuUelWMw3qZeBT+TG7gOotqFLPwjY
VC0yJUzm63P0zyyuytpDelK/qaKmJnQ7u9G1ej6IhzhtklwbflapjxY+JFPl
BUq0tyw2c5jbK26IDn6273BZVxJlOUVKYaCn/DuSr/bBhHGX+GlN8ZLkJ8VT
+daeDxgAXm4S+yYgEc7QDYxxSlMkuSbbGOilw7tA7PnE9HmtvG4pw/NgwcSa
hmhbyOe6JqwKtkqbG1aBZnLTVYsVsjUVoE6n7Ns/buYpwXxj+XPPTcqxji4k
obg1Z6jc4cEna/w6+0840IZ4IC3fA/UPcJ464jBOZU3wN/J2NT0WhquiwnWt
QyUHpQNsFZzQu68wFmuCnKTrlYlaM40wy6TfEcZLFeA4yIEYc6SbqGiczT0k
tEpuYNdwR7RzTFqrFbPMpowU2Eedq5UIIoHpM17HwfXLkZwW8DjJEOSDQtIb
T7/8BIqAaz/f3rs2z5N7BgppjNsMulZls6Ju+ayP6utUavl5D3AWDDvFZtgU
N8NfqAMiVpH6kXWfo16k1hYmy6o8P40IQk2C367bnb4aP0FpZLHBtZMDV7/J
RpT0NIr05BxLV7Zj5IDXPHZqPmrPl61R0VgzpVGCpZaiVzHZbvuCpMVBCN3v
ySKMXVBbWZHYidzQHza+tLmm/P1LGklfmnVYMKQwLVfD+gc8yoA0O/ptN0X7
qa0oq4ebbioAv0V763QATX10uKQC5rfV+8OuzAfxZIwN6PT9Litl1/mvUgnr
baXnqmLQOtakPnniqScg7NAAg10QZDKkIeqkpGEFkIYkEYJHVHzT7rmUPPMH
Ny6CSd+6Njj5aajL1fz/yV7xSB6o03HBsfcO1qwCVBmv5cpPVGE37l9djhe7
q41mB0/v5mAbIZJUxvYeHTGir4MDPw+d4W54coKuciSvia6swJWyQs30c9hN
88X+17z9BOMc1EMXQuyoB6j4yTIKKU58SPrejUKYvXiMoJWltsCFOtD79xe1
cRK7D6/xE/2pjPLM8weNzLaGkjnQ+zlgHk7P9MCfeqhfg/hlH5niHjFUOcBx
9Zq0vQ31LaGVF++mL/vZGf6KfacrDkOHnAVCy8ktbCghPXfu1tyGaBSRpKWc
NbozfcCYO04iC472iZeUXgG6zhKq2DrqPhnT6H7nOTYp4xYZ+YjQCrjQ835a
Xc1vrlXo+63LLlm4dW5WoXh7RLSlxiLUmn7l6lV37mfxJNScohJmFmxGejwF
CsD58fjrBg9IOj2CyeSJ93OsM6rY3D/26XgiVUCZ+xzfKTvUe+rGqEL7nWmN
TuYjRhKsN6MbUUWfi0H52TMFbKvVPgGyDcq0PbviY2LegiNh5/HGeDgLIwBV
0mtaT5oIZEQumrzvk5gc3xJIEsJrCHc6QDTCmROE0njhG/+TNzPIBU2aCMW1
iGFcnK9E53IWa1KpuiZ+2xfEmMBI7E2ywramPVN7vnSra5hxOT8OknwGFO8t
HpAGrYRSrGbN1cmQAHpIPl7GIWyN68Ui5AfjKQ0zc/mK0yQbggAl0bIyi+5Y
iS2n3dbuTXlPs+/qVFc8RCCybV5A6NF1KCUJEkvP6iFVDGl0KT0bScUS2CKR
rE1gd434rZEl1t6ddiSflqnsjnSEPRvKZPZAQrlbNlc9UaqC/qoX/76WN+SS
ksXjKLA/t0K9xmt8SlmNp5ZGW+gQpx4xucZHSayfOwj6rmg2lQ0X1+9q3B6E
tZ3N/FfWdnszQGCYNf4OmJP/yu6dgTlUIyu7liIpvq1Olkq4lMPuVZ0eF1HW
OM/4rC7L2fpewT2ZOt/EE4vMRTk5yeEDu6UpVnxKnt6j6be3f6c0ckb70VE6
nlRWjHyg6ZUO/Q2CwrvFX5jVZK9w3qhjGaOqsxjtOTWzLpuRfCrdasZl7XtO
ArcZUF42edZifDYLIV0cKJIvrRT9YUop09ZvUSCg0I0ZgQQ8h8ZMjsItl97S
zCEyokdXAy9A4cwb90cJ+ftzcMTMyfEKwz+jhVGKlwJ1Efco5XwDzXXBqzZC
cXKRrVhflOOU4cnkLHxRNamE3hw2ywPMbuajYESzg82CoAtCE1TSvZxLY4h2
3Cx8eo+1yNdvYqHADdvcFgRbp1AeYS1apVWCAUmCkqZ5KUj8L2lSkRvSiOuz
k+HzeHK5p4Kwkm/EmrKG3Si2HibiOCJA4IBVCB6aUsSydlD09DMWXx7RCqkD
3L0OgqJ+a/6Yx2QbgWSjqRvyHPt+WUIuAQZ/5Z7ZHL7WBGmpM1nZd7n++1CE
Co+JDpGG4k1h0IA++QHaGJwyXU1FIL/ehPQx1TGDMolh3R/5tQfP0qkR/CyR
RWbN4Spfwxg9W41SsE6OU2uP+57r34xB72SqCdpnU2Fz/M/P3l1aiNCaHRUj
jMcgsEY91PsFacHYrA7q3s4ybJt2aM88W1gnMmmSVSopbZPAfsStrw08eGHO
V++7/uGPuY/As02pS0BDvGBEg/3N1YuKk+y40eKuK93ESL0Bpq9Mytysc4N4
yVvqIPczKz/S3jqDVGmAbFAMpXeORK0YrEuJCUIZZ4Xo8mr3g1D5wRaOxHLa
G0vc0UJmrYv9AN9dqmW2qNDgq1MoXVbwdOPqB1dExg7z/SssX+ktc5izY91A
Shj6FH4lCd2Gz8BFjdTB+BP28+/bhXzClDWfIYwk5TsbDD6BtKHnKDtvY/+l
nQSclP02xKq13+x3WWWcWmojOeeIk5zEAbMxg/bbXK2T5mFPI2zDgg9DpLIY
mOwF6FHfzWKAH8auhe/CXodmTfI+dRFeUfLq7u7ib6u9+NFPnrHWlWSHWM3V
LMFIafLMJIojln0rXQ097JdRcr0Uo/yZGi7BigZXzcIUbZTVNTqx51ukIMXD
ktTid6adMnI2SszhkK4EXK4hzhDeEFaSQw3GvFTI1fw71Ug416fzo34QsOri
ZtvSFf7mt9kXjjE3DX7Qzc83ApsstRR0GOseE5U/ol+e7tWz6LPfz59dLbKF
T0ep2qLL075fBzS/DfdzHpfMg/BQ394ysd+jMB5PGeoIT/cU64P8ckb6i56o
RwESc+GiW+3gzMIkJx0TevJhPOjaB8blbR3wivUelGZoS5AqoW7soLb69fsy
J4NkgDty0ItPKtYrr4WfeHhFLdfKMLU5VRYaWiLbOAFSOIi/TPmTlQV+XBV6
mHkCHHApJLB1lt7hvGGv6hEjoek62Qj22dYE8RgZ8b82kIvsFNpJF9CKKO+p
hPiJgb2OSYT/DPitbEWE7Cx6JnvGTae+rwOGiZOCamPDgpRZgyIHsoFOJpjE
uhl9o6Y1ViJNL/mgYDp5rOZA5kNLnV3noJ95Bgy5DQK3hMyDXEH0a45JGge0
naHoefYRnXtrz14xkQrQt8JFQ8xfD6BbHF3uv9ITbNgQhaq2kuKibzNtJpX9
e2uUUh6W7v6E6RfMQAy5pGW67su+nPnMZrV+nPelWtAh0ZnGrPVWquF8Liqb
fOey/Tlmz9DPO+aVFL2qnAor98WXRIrzwejfIjIKSzBuQ5mvrvizhHkoaHJn
Ua9bcUNC7cf+EoJrSg3Z9rLJMrvazoWyoDVM5T40BQK5Z5qIMLp4lHUUk88x
fV93X3Myq6HPr4kF3BRA55uLsmmLn9DPE0Ck+mw2TBKPM0Z5q6zQw7Re313Z
uSy1T3PEIdmm+OPtndGwuo4mhNcGX0a8rW8e/CZR8L7p5gm85pgE1NK4abVw
BZd0NloAVLkN2UyetjSeNj7ELBgSDJ1wJuRNfDCl99NW2TOJx8lLouyAB7PJ
PFpjBnDzgZaiZOzShdW9wJjGIojJdw3HSQWT4UVoGF+VS5h/nOciLIUN6/H8
PMTdPHebgpCCcw6/RsER9L6idQrcvp+ZBy9uhen8518mf3CKn2bPs9Of+uJN
5qwY77BXb4SxkXs5LZxBIxcdahvbQfO24MYyWsVDYIJdNiKg8K+69fEK/X3S
yl4b7hWfLNAzj/qUO+ED8zyuDb97RCA5XN/Z1Hy89G5jf78pki+NkRI1TP+s
gJDDZGe1VmymSSlCE8gOM/QzV25oxnwaa+wvCpfZyGqUMqUHYp6Vv/uKYZfp
aCkpULV1SYHXmjx48XfKBO4d1vy4s0SPVWU3Xm50sW5kiDiuJonujybpB7ZU
PTdS2nYy6hfnf+b+Z5kkyrNbbptd/RU21jLYJ5tuday88oBgSRY66SjyHCsr
pZggnPjOTIMM9gHyQdh7g19RyKMLFRCRrPNe3jK6442KAII2v+iG54t4NsO3
fvMybDVtuhsNyBZorjgOPgKtSIFF1OWEiFGmLGveKRCTFcmPCicYP3Exol8l
FnD6vyZfzojyFnMqLJNCIZ/J6sJlN4lxmkE+rM9ha/aRErp5lO8nRtjOkf8Z
WY7wZFFVZgwTwpIS98KXktCIjA9h/MzVSO/Uu2aKq1N/7e5k717WEJLx3Uvm
o2iRWAE3G2ij0YbBg5KGC0CGgbRgglc37OLL2Ziid7/p8bZhOFdDuobuNHEQ
v+xOwTR6/c10IYOV0aLxwCTD5TarBAm+fBUEdhsDfSRXoNRzm2kD0uzqtUox
QwdOg6EkfuwOXXdyi1w3BULmNBF0OE7SFCCZbLDqUsD7ZoUGZPtLnQh/xVig
a1coWUWF33lzC+azrdb6rAWoTf7GKYd/9RKGyIHXHOdG0OzhpH8QFcmhE0Z1
Bv9x6GHwnGf86+rA7ADymxBN7S+Lb1Wq7c9PSI+IzQBovIxLiGeGjYiOnQlp
UWAw//a1iBN7rVWTc0artJp2AZ7z02PVm4FSG0D3Bvqu4zElo4vB4bhQhJY8
Y7ytrpYBO8dAQSwxiIQ1Z4RVeMoUU8QFbttSHSILRdOMqh9CRSP8IR60X2tg
jEJ352PbfBKWhOKXC32opRTMepljHDqercJImZoVe657oR6LhsxfaXAX2xYV
VRe+yu8CtIQEzo7oIhEPevz/Kj6SJdDVa2rAeqW4M5DXY3qrrWSaRZOiqBIu
ptFFe8/yR+taH3TdQk344wunKEdeNkBGauJvnCZ7f3CVIicXhcqto/lxYa4D
64mBkDVWCI2HGx/unL/N9DJBcIO72zDksuV29+OxQnOgC7N56nqEpl7BLM4P
2fmJPyvdWroV7jkwDGzU9+MSogIYmVfMZ7wm1kv2jU4l4ZLq0HDeLs3zuL2E
LXphPAMwNbB5SujbbkA07j+YLWb2i/ZAtnzSlprkfUx0wcUGS2jGE63ZZM/t
mH2Avcd9e5Vfbqbtp2qvsyLVD65XCKzgrAG+ypmfwDjEHV/9J8EoW5b2Uic7
WFXsr9/limU8Py9sVlxmppW/OuQtsDgtmbplgvg7ZlTmmGoMR3PMH0VnYSiP
Miil7NUdo+wr8B2NDkiCPde5Kj0YTngZsuldDxwQk48ZM2XFF7f4L4g1HcN6
jB8SKAyUzopdkJb501ZiakoRqOq6mcmaYEsA2Vb8AzAbFFuXA8PJXA8DNzCJ
hnPX9GLsCOgTeq9fo0Yf/wIPLXHkBdydH6V8UzNh1IicwWFo0dMGWA/sPbge
0GHqlhMfHdsvVjzVv0j1ruTBG6MA9bJ5LmfMOLOFi3+DbAusbzK9WhIZcXGL
1Oj4xmWcqtxRs548mtFTc/EaL/wP1BJI/hW719C/zJ2KXch/2ETHmRjeKAxb
OSu0CqHQcUAv6jX6p6pYZCGxjJRQ2Iy8jVI+NX4c5RTIYlqaqAuf6uTT1mPM
6fUzsHSWEtrChRRuC/YBy8WQKwgKAB6+iQm9Ljqe90xzhkNyC6okzzocrpW3
aGKWvCCxf5hWN1f4O0fHbbYUiP9HNw3Xvq6/LO21BNH0uX9qOt3HkE10M/gm
95HL2wpUcuCacJZavzEgEN+Ui6DIkuPd3xRfbN6B7pFw0JCDWiBBAIocSjxO
9FdgETSfiWSaPbtnSm+F41yH1z1+TSpJVdpX6yxT9EXee1jj3ufsnLCylsSc
0D+iuHkWkyyTc/7d1bEOTWJFfoUpiXcGfv5xmvRT19NHdyP204qIj73tvKiS
rrkhctXfkbQq7HXAAAOACxDHzsas/VrffsbDWqtTW32RNAwOd5nke/Rt3ddx
IXASakyYTJFgB2mSQwvHudxhFD4Bz1HeZrxE6nH0TQTIapjtmirVhw20OtYq
9AcRfAHQOqESYdnr9dmBmTYt/QS8s/BK/bHC6sp69EHrrUwvr9CKw4HlM6Em
wX11B8aoQSywmIfj/QqKE2trhafbpJIeGFLZ2FOdrEvWhZwAMcj+xe0PRWhq
OPqLEAjJKyb+V6/Mme2KNpNNbVt0IQLyblYPmNqjYSpEPnPHmr/npbyOQw/c
jT2GLrreJ7o5vZgjtglW27rHpB9txVOQ8ud71HHn6flGOfbL0LeROYyPPYVv
ccA/TVRddYgnJtmBdDf2P2wr5q2xkTycGKC5FA4uzHKXgLpvBiOszk+Tuiyy
tjOdwevI6iW6l9e3uiAAyjvGwpMscIKLlcz4+SdA6FkJK16G6XyuustREPqh
WGR+OC8YebTGkqZRO+H2bOH3aFUtnU4jNK+Muk4fvO/X7Jjx/j235lfu4NJN
yCL1uvVlkWmpp5EnNuuXmf53kiePPOK8SAElzh6Ijwq46Lq2l6hvFz3QqDw1
MeWq6aRGocnYvlm8V18i2txdPj8IzQ2+r4Avj09NGDZBBGK+8eW/PhZ+T0wK
bQtxWQwT/7x12oVzH3mUaLegVqoqgv7fwgh+g3o8awuNtMukJK47JNVbISb2
Cxrx+BOqi6N09aa8sjeoKRo+7ASdae0tjgigIQUcI4d52woG6xfDcdnY3rpf
aLBsYUs01gbVAEcOjvctNuS9QUo0q1i1oxa0TkPsPrrSr132VSj3hEkwJg2P
tM3Jl2ByReQSenSBlUqoR/i2VNdcr4HQqiAYBnYBpZuCU8rinh9n6Bco+/N4
cMFoGttFmT+RZHB+d5YoR765BzLUTpygLU7JMes9LZFd06X4jT33IBdhkHfA
WUIaA0q8VRxUB7W9APJFoKydJSfMYefE3tJcY0jOyCEGDkX3+ua7aha9TaA5
D1ip9b+a5MyF2TJD4NhQESb6FBgfA4ejcHbOTGu8nFs19EWIfNWKmxsh88+S
vYXPoBRSUd3E9t7wHbJi6s1k23X9WmRxCwIrake+2EWoy52QXgRtj7xeBOTA
DUqZ21i3IzbfZ1VZP+l0zo7Y/cuZtUd1f8hhODc3IwUYfVDoFq3CAIMo9HlS
g6brlSkiJKvD9P5d8TNsevy68A+E9wrK7A2whyTi+UrJk6yDXmXz3C6pwCxF
0TVsrKgL0yBnpTEWY2R/j5xvmGaBQL4uCikDyVdRVG0VS2sCQSTYJYyUXPkZ
oEqcjNkVsanndeMvNAFDy+vjP/5ZpcflU/U4Mb6QH3ap7s1lZNmtuclCoB2W
K5RwsUJCU7nbjd490/5nKcwqMMQPG/TFX+1MpBjMGo14akAmo5gY87sPvp1K
znaoUQ2s2W1JZQVMq7/0IYW9Sn+VyVbXGYX29ItFLQvHn8fITaaAeTho7CA8
C535tP/oONCgeJW3MNSZtXLbcqRkX8tlSBKzSDgaShea8IVBmrKgTtdWIzhc
NMFdWBwdcZIWPtS+UKVy0tEBkPazw4xj6UqQvgdsJJ7hXG0wGw48zsqQmI+A
+SRGZHiWU/bDMcPRQ/4oJel6iBVibYh9fhIgNj+QZKLmPefiHltqM3njTTWb
89YeK/Q/cOvKBBArQDIreSvDbvWrJDYmYBPPRr9AAKlqMIKvAV70mMEzOQRa
uHLdzKOAFpJk5ToV1b+yslqkr/4Z9Ye6Tms1WSQqlSq2BptTq80PwNS3oFdO
wb7zjgkoo8WyfSaGb0c2GlsDYMQbBl0YZBq3TpoExoA+50foYFX/qFLVgoBM
IvK1TxzWiJonOJDPoBqGxA0Vj7DeSs8LMYHCYZZtek/BSF6E1E2l9aphyjTC
W3dpTiOhsFX2+p6HFCz9OJxNxXpzaR0NttpU14UNgToY2VqUmRHwVNRzl/9V
dZg0iv7YO4GpsEBPjDqJo/QCZEbCtYQ0cjT/H7qr5slyvDsXTUYwu+idUB+l
gMKRuszZCt63vj/dbU6Mx6ayvbMT3FPrVa+8ZhmGva5s4+9ZrD5CfmctVZYN
1wxCW69bmoafFpF6L9burK3hKCfqFzk7lVzEo7Fs0HPhKwjCTfF0uWV8J4+V
Ben8D2jx/Q4aJAxO7pXllQYJDi4XURLWJX23RYn3GguXVfc7x5od+yFDk7ZW
+k01U+DlJ1aEHBjN0PkzVVM6LfGCAR0Sdhovj8tWN2210HGbymYXEfNDzVO1
wHuxUWmmDP0gcPfOwMZkAIjMIkrFTJPQ+ZDUEFQ1M+GwGl85/WxK2uyV/LDy
FhnDzzPgp/rxcxmlvUFoErwPNK6WowOr3TVUsvVn4ee95FnT5EZkBy4+waZv
1cas3uugkyF1R5TlCwh2ifPsRoHbBWrIDPOthceKWPJbG+wJE5hjJT/LTSOF
JM813n046bYtf1ipF0wIfdwPwS9awBIVzWFP7GoLHU5T55ih5RlGLwVSItmj
c695gQ9tjwRFaWg0MuHPI7gLHv+2We2vgUz4U/eeFn/EUhF1Loy6suiz85ct
9LWwRyotSDvaZndo3fiwEQOyM1thOU36v6i3LF1VasLSLKMRv9Dtf3pCo+qf
M2FysWDKeNX32vr7xnNqMxLBY4hWWB7smLjyMiBfJj2YBjAQe4o2vwEHw2Wz
esQ7srRaLK5z7Mj7rtk2HooLziCyoApSJXQcO3wkUnCw4zf+FLKm8bjvFAOK
xbk6wOTydgKCnkqdZVZPyLL7+OzkZ613FzmBTPEV66bjHbYUCoW4DoCqpV8C
tRTY4EH7up2c7JnrWzd7G3VWDkF+EvM5iugRe77K1Ym5idBH5ZUEakTxgtsp
TTjEwLAE+8XkljSp5TymlsGW6bmdINS253Zbki1Wv00d8ThuAyqd1rM9OxAH
birSlm+8f4k3H1h7xx1KLO6qhcz0iCgVLMLv+b7nemJyXo9h5Ef1+EOi5mdd
rYLACJrqQt2oYUUIGeycJq0A+9y0JtSTcIngeK73vw5L+sOhmthjc9CB26mg
tRIvvwfBJd5lHLCJeUSlNBqSbCkiKUYZ3puZQKZoimr3AeHX0I2eSILm7LKF
iQVpbYymgG2HvqiZU7t4TPnLz1WRiMvi3UV20PRT0ULrrJEs6yxXlyH+bF3F
ugdmxRRQHztyuCuCm6/7Pb15/ahWCytMyST+Rvs1d+OYuIPxD0UmBLofK1h2
8x5zjNNkQ+OiI+ATNjBObj5CZPRBrKJbTPuo2EbGHcVxqXRfB1C2eaXKLory
fY3DHcMTPiZz+U5x1fX7XOOQrVyWFwTPLc4gSWf5TDt15Yjlpbdni2PuyYOH
0XH2xrHh6vYeCm437QNonlxzXphQJiE2E04FMH05Zh2cOsepW03GChuEz18k
OL1wbux3+gGYYKPtwzdj0F31LARcYm9KxCoz/SZl2kcqTlto5sYoZhWJVYH0
NehEZFdYbucyzk+SUXRioJTaZzhtXbybIa/wKIVrAaIkN03QQp/3W7i+VuSz
j2Xx8UlIpWrftyrYd3UQXgDOTC6B/aYpbiCcEkdw8zlrHUguLWdUl4RfYmUZ
kzJhAn8xkfpqhVMS5sVMSOnLkQEj84hZaxSaP5xI7XIRK2xS0Z8OIUQCxN6j
aRROe2haakJVgt7xHSAhO9vyVz8TE42GXC0SQ4KnQA9xPNDprJ7uJQNU1CFo
yIXd4i2uGqe5KB/u3j60o2JfXqRW93ynlpiykY3Eaacm2rqmF+pzSyKQpH6O
pi94DpyvABszwBL9ixiUV6nIs4OJC4Ts8DWd9UVYRAwITPNxkZlqhesNC38c
ydeaZ703o5xBN7rTivMCEJ0RZ579KJ+M+fUhEX2VRqbP6X9RDzHvSrjvWLkt
mR/kqK+/n94RcmOgsf3PEO5Jjdlf6igYRhkzMZUUBmqK5U5dyPrBnRwmETOB
Jccm1gP4RJeXG/kJxnCgsXoTa+VcxKucBYfTj/UY2Egbc9fq6cIbn66uL/nK
OcVerFTzfckFYhPcL9rfkpXHM/P4IXPyZLWleW4Av9i37SkPbVbC4hnbsDPB
6nMTy6ljG7pexib+PNov3jziEZ7TScSns7IFwP7fBPiVp96XgjUHEFX2YzDx
iVB74YznGmEh2lrVwx4L/Gbq2Q0ho8UYtrbk+ffcXhmVbLIl4UW1o6z7XJOI
oJfcBOAjV5WlxLTyMKgqOtOaoohwh9DQZRTm7dIDIh3g5eV2leu1EhTSvzlM
vhEV6MOZLtq4VrqL9lkKYakQbcmxQSBYy9UpXQNoT6+945Yw6NUaxlKfraJ8
Ej28OSQMBm3NbzswRUWm+7rL2CnCxnS/5vtMcRQaM8jYwW2Z8CHX/F8hBP50
Lm8pfAHOMI8Sevf7leVyTkbh7lMH/a9MxHfT6c6IOyPxZq4RSQx5vQCDxU14
2k557hiC2eJL+bi1fTA8ZPuqBgwOIYu57A/vghX4WUt93zIi3DD33zMeP8T9
Oh08+UzUNE0hbi57BgxapmNFeglZKFnAhKwZNjd2+2A6SOyRILmB8R8yRKg7
MVur+qM+rDfrbo+6Z8ANYYc/JPIbQJUGNHm0zS4HlM1yqjmICzU0I7shWCxO
nlp5feyUoFaQ2CGrHPXGS2crrhZqx6UMcqBYN0wS23ZSECbcPKRVFon+4wS+
8ODUM2J0FPMCP9GeWqZdpUqEjmo7vpTlwlfr1ySEgHU4n1Q/yq5Av9jFZRIt
NDUCXZ8OiqpPyGHDymewUHv6oyEDNMT1iu/PafrSAcu1td7um8hnRnN3nTA9
8RcxWVAq0/Q4Iesx+0oSvhWFqBcJJvS18m3MJ+wQgAg4q/6sRvZrOKdmG/6o
cLsz1b6k6FoDTHR9jxpqZ8FhfvOLEilDIl2rpxhJf1Honj79nMsulabUSOBg
lfvcxwwESk+fE25bQPTufJwW/9BocEud/FIlQSQOQVSkocdR7liZyP9sK/LR
RnqyCivgwtBDaFK1jYKSqisvQsYvNW9vTSvoEFESeSutRsO7o3IILlZsVagB
D/xvqg8J4eGkBvzgmE8+gipkgloPZ7F7fn2KLK4Wc9h30xnBXMGRFxuNrttf
Bb2yhrOHSw4ZCQRePhyEJRpiGu/RDUEovb7Y27iVfwLIuXDmffs4KSoywcGx
XKwMpXsq4qcYVadpSRNOZPrh7pg6iMV4UbEqvlhSXqcg+HyBxhSDLrpn6a/F
DMXxN+v3J2iCaiFIkuqRgX3yp0aZmtCWqOKJlgGBG6hjXTCXPwrXHyw43CEw
6NMWl/C9vNTkG/U6ObzxdoROH4dSF6hUhLznvYKoas26Ds1D4ZqK/9nHOU/x
vT1WV1x40PjNdNIrhc09Ud73JOHP9UK8KYITXA6qOIdtEXgTVlpA4vnXw3a4
oiXh4HwLWwjaGKxQGwhGUpzZa7DgaUvjZUb/N0aSAZ7Nnd78rgqIK5CSuYaj
pk13UFyrGhcX+nBSeSFan19C30ZhHD7C/qpbGr76ez4KvMivVYuxNEMl2ZVj
3OasZLtyhEucCrOdRDMUYs0Q+37XWy3XhT5vc+ZlaOMwyLogdjsdwVbXK+3t
xbUTOX1MSZzgNgpI2uTX8Klfonc535/01Ji1ygdy9nvx5SvAt1dGnpG/i6tC
LmDOUu+C7kzLHgxcHW0qYFjcz/nPZWLMSK1HqNjz8DY+lxvoxbsSmYAcXpQU
VwnjMCDFUnc4rzHNQ7WmhTawFn+HWwkG88rV+SGSwNelcTVYqBbUc18nrwf6
S4nH8uW8nsLbImRtVECCJYXOk0LiM6LXoie0jcvitEVWflUzTD8F26n+Lm3Q
lzGNUsCvBR8a53fL9NUu9vVzDxJXkM4CaaWfK/KAMXJEbCDtZejPyzrvNYdy
t2ll5dUt3NRLHp+WhFSq118VSkfGm9hfUDZS5zGjquqjnUvSROLVtI56yt3n
MYo5Nmbv2A1ogenNzu3/d6XMMqUaqFiPwewBHUMrTevz5S6G9mPKIq+xwBnq
GMbbsWFbwG9RgTopcQSf8J+uO91DROIdKdZVLJ7epB9YOJeuq+lstgdZjdI5
HaSja8t0bKyWcQmRS5QltYjzTnDg49V++8QfnzCKK0YdvK40Vzcj9+yDLZo/
xb2hLV9B9l53rejhfAP5dO0goB1sLYq1TAE+f7Ab5YTH8tCPKicYyRfYnPah
qWs3L0vcyxiwA2XzVIUQeK7xdt1DkVWnQpNv6kM0oYJoiB0e5ur28CF+2QBk
hhgfYNGzMKZzpAXjqdq4agVHPwawS4bG6fWXFuxKwyDtdZuBzoDB3v2Z7cl9
9RuWjoHX+l21qUmu1akg/+RwjpF94WuMZyJIFw0ENTbHblv27fPEP1l0nhjz
88Liv9X738+dM9L9EQ7rIzBLcrHvTsTKsjclLq73ZZ2xn5nJRW4AXd7QRGoc
ZEOGoC5d738TzsrWpx2r0JHwFT/43j2GTD6q4Nzx4sqYFVFMr+tB7l+OrNDT
zEZW7uWYITmm6HpmMj7RJH6mBBujrolI0IZ/lPlAftR+Er00b6EV024rOLag
o0IKls4bB3c2Ag8IrGace2PLGvFcx/EoY+oEC+CkbwjwBnjbKl0akX5zr7Cy
iWEwbPo3ILluja/+u3Tx/drx2J+09SFk6gtDXDkgRhJjiDe7GYxGhbOfikPp
3pgjBztG+ky3vUHIN0IqkG6zStTJWdhwx2+JYLtpqtRiIYdsKwMJI3NBgAsE
ZfQc0PfNZGQ6iPI7lQBtIwOEzrst8NiouPdaLD6AH/+u99tgL66VnWJq8JVF
wsI0YEpaguXbsN+Fuv+Def64C6rD+y78f6PX1RCh4G5egNdT1SsA7aAGqpiE
AdKF3XfksYg+3mbfSgNA/PjMdbVnvU9Iyq0e0xjnRxlxRGP3U7SDNAZnGzbe
tliYxEs0sa/YVyb+XJ/bv0NTu72Boy9a96z0H1FtudTg5gWsZvI8AJlfuwRx
zKIqlg62bdQsym1e56Im5hOvbeh6kXMroZI1v7JimeloFtd3Y/4NJ47oZoPn
AyEH9FF4VIgNWsjKjDYn2NXOJrdmx1dLgpK8xIVW4pFOS/VH+XGS1k3zGasq
iUTLQ/DXz/EIrML8bXFBz+uiTFrSxFpCQtyEPx6zcIv0mxMUuPUUVesUvopq
vaB05M2SBDXCUkm2JgXKj+t3PIO1nUsbaJwUrENnN1S40I3IADc5Y22lBniR
pDpBodLjcN1EgthfqLMYrNJuJZpeEu9k/f6U1fO4s6rAPqZW/YCaHBHHG7CD
ovXSJSW+kyOHeKg9zkJ0VhpdSALeLUBfjCdQSJTzNoRAzHOzmX8kC7XLM8ab
vnmGy/EQqlfidManm3hq+JJF3g7NflfF3BCrKkKKZNW5rtgiHh66MIiPpJZ4
b9I9zsCB9tnPmHDzREhX4OS/DDKSjQpIFqOo86wChLM9QZiRda5pyMLRs4e2
5b86arALxBM4jKfuy7/hipZ1ohlFAp2AqBGmwWuKhsJeGRft4ViGYAJVny+4
ZyJPKlRl0Ur+F6kXsjl9AABDsXizrNw9PWh7HELolpFTxjswwkynvutSPF2Y
c1Xt06Muo2oMGtYqo0/gfRplgwpTshX40cR7jIFTqKdYQ6078YfclL7Lp34A
OjLtQPqDy1KIYUVOeS7pcAjriYc5NFcblZ6vLLX7R76UevCiiXevYDU5jD7o
7B3nJFTdQ30DqrDc2Y/cn7JmD8nffmQq5gZv2oA0yeVVOFoovqarsDufF4NK
BQjgyF60GrKl211HlbXtOxDntipbbeRVIfsCkb5sQ/z0mtU+ae4CztkZ0pYK
5oPwYjqWNYYvp0odgKP13ekU+Nh0O5sDb9t77qFumXdDd4NRmzVwFwHVjoVO
aWJgiko09uqCbvYuFdOrWl9B5Kvr1CS2LUxcgUPn4fFSVIJ/KgKZmy0JZNc8
1kVFRRXJ+kcmLlOYX5PHTwt+H2HMVGu0jxWYDUN5TKjbCxg220V6j3VVqTvw
VqXFrG2mOO5UD8vvsqx3bz2hqOOO2am/nus+ReaHSF5+k3LQQEzmHvuI+jln
ntwKrIYcebdzKb9O1WNhLbHBZlS+5pwoljf+W9JOGSyZkdcNNA6UB2FZTNMb
hyIEkXpRTomh1ktPKBnxBzHUSBpGkqD8+rj/1YW+M3+0wNRliDvg4Fnvztdz
1UOWMDyO8E7SM2WSbAapnFubm432rmRK9PFsAc3Dg+cQra1GT97SGeiE3Rhc
+wkaScmqiZluT63DIcVFAr0AeaLdzYUCez6KSFsf+ElX42eMMogWYsyvoKkR
iK1XqnkBs8YtHXKC9o+NI+oRKCHxwpqp9FBbdRTRKscM5LmzQAalfm7bCnWe
TbuWrkNR2mz2GIZOEhKNxfMb1M5D1Ds02f1DRFTnyRSdTXKeZZD7n7XcxaPr
cc9Fk8hDOucRbOmgK+9HNmAGhyRXRPmVLYq3pFgx4pf1ujbymWyK6RWsmXqx
FKZ5FsAoRf/PuFLbmSZCDvsLxO1UsNMLLKAh9Nz22Hxc2xSfdvJGnozwWsQs
GP73y0TZ7z7tbk48i75S1qA/3YD11iXrc7pRZkmuC3/MEqW4Cptb9tuxOs+m
YpZ5aCmhiVm8SNM5U2gkRBJQ3duMr3j9mAnxT7rKswz+dlWrbseQcrXkPEFC
FdNApdsjBeLLLpKqvgrlEVJQIh+UUuQsYNcAgsGlYzBY349tkzMRGh9AtowJ
TGLCQ60LceSVS9EDrpZEmc9MCF6h9Z2mZCKjvvhV9teqmdktw8RH0IFKhWLj
k3Vw1Tyd8OAsrb4cnKSGbi19Xgdc/8nQAUFtg6jnrok9xVbr18l4lmj+lczv
3hfx4ctc9HDqHVpuYy0O7kDWGFSor2TWVKvjNs20TxM2pjMSzU3fkD7VHvhY
2/QJVArpX5XeRgiQcqUeGSv0uIrixrL9RY7BOZ1r/ghFljyULMYEZabHvabx
xJ124GsHocHiUKdWfxv7/PALd4ZTAi17qIx2PCa8BJXeehkhD03r/A0+tWc6
6SVwu11WqSfUR/8KUpmh9KgRvHpKS8g7BHKITmp8yXb2BL+1XttWKgNvGJHw
HmtU3HsCeleSGQaHtwBiPHdB0w2280p8+zvViG2l+Lu5sirrU9E+lfwEN2VN
48ZWMqSrLyM3xeGCOMF9Qq/blPJwvs3936x+kmJUM3xwCmNmq7dpOBHaUzvH
MD8ilau9XzhNYYScSdkyZDc1p026YQUy/eXKU1gKzZCufSUzZltHgealF3vC
j7lZUDBePKrzsjA4yR4u/B88/kCd+2tANAdzx+U04JIvV3/wUhdn7aNf6yTg
k5omHf2BtagbN9bMjyWb1FDhM3vtoV55ksDea865OjVlpJ4/swYu8mXsSfO5
9URIk71ZgbHQUZkMBpfYM7Rbk4OmlVOWbbpfVUvCYlcjLRhcONI4sgL/Vpy7
8Qv5N17xuIF4GW54TXsOJ/k2fVHQHviYPmwcfYXBo84woUVEP8vIqC0mXQ2M
B2FzxVJEsqIiDHDmHe52ARfeywzGl4L97HMJ8Sw85vAbs9tUWf9dMLIJuBFh
7hpkD33kfkRnp1LqhrrBhznZ4mdyfN8Rd/TJKkR+B0JyhC2i60SHHOqogMYm
hVVeE06hVk21VsIWMq9deh+UwyYNIX+TZVwDq0iSj4KZn6Wx+BcZGKhgeHSr
phZ+1A0Hc10tWzm7riC8u+2oUUAp0zDfpdYsrIx/bZuEC7oJjSNdyP9aZpyj
g9AILQB8XTmO0ugwv3VIvUhul4c+zq7eZfc4MFE4cyjGQCsju1juvUJlxIKf
pO1f9gEs9Ic9pASgFm4EVEwf9LnVSOKV5hrU2PPG/sPqhkSaffORsmaxdRBQ
oXDBO5LctOt/wBWqgFoRZJtbf6ldeidcEkvRJhF9UEp5FgEAfqBqCeqHzxoo
aQJSiB4Y/XNzAmnEeFzxSNXRWgr9NjsFTJhV0MF9bt/TRE5w2rpWiyCcly3e
h98BEh+vAwR7vCRWcb4mo8QSYSJXvEaKYNP415KYt3BK5a2VycZZjb8jIVt1
fKZ4wtgdLSUKMkGCcWK5Dwly9GCgM3s19gMSdCyndsUvZnKe/FjdmlLev1Ld
1hxZVcE8/+UDgGz8/S3WxnChjcC0ai8XOvIv4JlbC+OQQrjBvu24ZEByGR6x
7NVqezlpkDCABzGVOLZ/khg0umBeGS+f+xCqhkgqzDSkEf/QSZ8y7Cq6Zp5U
5F5+mIiuVzfNOXSqFkpjuZctvlShvLlbYJY4+ZuGEc5qAkQ3iqvOkfOBemsq
5Rc74wOwZ/EhIAoOnzlC/k+n7Bm9/69uA9rlUaFVjSl4oh1trSgn8VZrL8Rm
KD7BMg9hxXsOXmD7jrlninTFBHhzDuK1xDBBHuSfjW4R+Q3ynzj4ZcMs5TKQ
pLbap0zaHjrq0zRAcLJAF8thP5XDJap/uAuUAb2R/Sj/PXEMSZQK1r9CvDWW
LJ0CKIxFoFLxHhWZ5GfvRJAIPeZyM4G5434baJWV0EPxvqX5CYFRh3u6x+l8
NXWWahlvXbi3LZdS59LjJRssjMSG9LzgNwE2DuwdFEosrl9FN+Rglzu7ifC5
1X08/1biAxUg5sj2LuyjZUZuDatXGq5SPUh/FXzddhaWTHICXQZ/6C8OUzk/
pszGyI1CIDRY2bOE0vSv5o48kMBa+4hwqYM0MaJVzvDdnuG7CiFjmVkP5km7
d1ckM5N94yZUIFb8PHAVTBh05aCVa+yU7hqHJG8wLjQ9yBGuY86wwhgHDfAf
8V5UCNiOat5yWe/yFRF/eLk/RfVAM3md3+licF1GF3joqSFdv4KVMDltjfw0
2sDbLfqyNH5/s1jvC9d+qcFiNttWSRRHil2mdDKUvwKg2TyCvqRbzr8/kLQk
BdBSLHjy/6y8kLIYhJ2S28x8TKcLhwFWHabNu0CTTSUX/j/MnzDx/OpaGFai
7YMepccz6E7Y0u+EpkxC5O1ZTMH9IBNmf7JJc7U0mwvHqIBfwgvbhYNzM2uC
Sf8vjNaijCz+aZezajTlyJj73ae2iDnp4cBskJD/4xDgkyoT0XbpQ8lFgRLs
lqgsp+2WN07p7d3so3Lt0pQaIUnpmQy4RXVLTLf3jCa7PJ3AgE95at+oXdLI
eR4pQGXjso+g2Dq1saY2473MljpPEpAvHnBs8YHYXOaBwfYJs8HLtTEhozwP
fqgaBOf663iZsmKreS0iMUBPL+doroSgCmr2m5LizMnN65aJZapCFqDc7WfI
6uygUwFt+i3RgZFenJS+Ruj/i0sjMp4rEdY9OX4d1VHOsEbBTGiGUH4RHomI
FlzxxB27iETIGOWU/sdC/JPB9bV7qlnSLw5Z+K7srePTvNlikQwr2TGWWjWn
uxvC28l+ARVh8gJhwM6Gx/AUFGtLpwkanJG3x4oY808QJybcNA52JKHwxEvy
2CfO6PGlPsrMJnA5u/LkNiEWj9UiCveURE3RAj/3qJpQwIZO8BbzMTssrPQK
8vzdGgqZtLxuBYJz3ZQsKEPNHssTk5XclnZn8cGOmuT1AJZy8aaibHgHeJtS
EPPpF+vhnw94v+xXPz+Dayp7i12CCuuGh7MYwSO9D/43Kz+iRsCLBN8eZ6Dl
rWhczg1xd6Unf73SiEwcMY8nLa2gogqpbhpVbrINR6sJoAR9kI8ugfwEn6hg
LKcOIVCDsquzg/k7mQzTXhbrDDAGs/pX22aBFttluj6xy0RIZqHkAWapjWpe
9jZ5n2xxFTU1C17A68lGNSQTUUt+026baBfrWvO0FGlVHaGwfP8XPGl3qjoP
pRFFprjyZ+OrRtMVMGXZjHpnYW2VdqtshoqYu1SJWAQEKFkE2fqd++ZmpDQn
sffkSDUMYb0A6dQt2BdUiNIQMnOAmzJyzmgN962SD+uV6NbSOVy9c5RpmxEY
ajibuqJb8CFRpEsOg1ugqOY5W07KyzSJgLxcbc3MxEcQzpmOxM2Iq0guE4C2
4woFC1/yhgQzipiVT+dkyNrgwI0etOJxtj4yE8+ZGv2CGWMCmB9upJe9Q+9h
+2ClTYt9nhwHM+dBR+QIPJ14w2AItGrmjZIGKjOyR3/Wtu5Spqd8jzof28O5
Zf613LJRdkFUQCqzsaQPDY1h4hLYLGWPOwFD9uKW9gM/iL37/pyZBxvH+VwQ
4BnR8jGez5MmCFiotQCulUaRFw8cah5TeKi9CYdR2bQg5YABp7nkfD39Hg9F
SIj3xuU61QyxJmsmXB9HaJd4w6MxNh0CDfaNCJN7g/yGNuDi7hcqJP3ATvEW
S7H6OrGbW7YXu9hRsVYhSuLeQ+gwKtOqsrLAB8gaG/DFuI9lPi5r5+xKEcOz
rPBo/OfEIeZ6s1qpkb7ubMkME4nHAqc5HwBlJCFxQcbVv24LGXSGczPeQgqZ
UXy4A7eHloOpl1cwQJzvpBVLxkSr5yUaHTldAWrX8nlKmxgB/ZL4w8G+ar90
pHv8vKaBVjzodUXQ3z0a+GAwhkU2Agx3/8G8RMcamZEzB5swL36fQUBIZWvh
5C/Grn252On8wy4LM4QCWnVZv5a8y1p/2/+vk/L5W8VGwaDifYFlGxCb0m4d
oBjoxyrkwNAso+P6dAQmUAewnTdKFqUJED4UtQRAnALjtpvgtj0wL1NcyAkt
DcIqxOLiKsn+tH34oaiQotycSUpYg1A5rG5izIoWCFPunAFdYEU6vAPRbGR3
0hlf7vJ2v2YRWFPpDtlP3kQyIKWSIcKy+uKFrRtgDJ7qsxzAM7F4MWB11bNK
irWhs5YVK5vyvHsEpe/UOmXomvvhXmVdJuSyvkOqua3aerBwan/YmzrEDiAb
A56Y3wLXFZSlW2VAkhboa2+sdNmDq4WwA1xGNcPQfQnVW7kmNKDgPx7j1TGG
Fcjekht7buXo4AJgmWhIZ4MXK0bIfGpNFxN772xhuaMx+XB5KIwxw6+JaeYD
utdI2CvtP+67Puqn2hp4aL/wjcPLe+mvjTcqRBqO1u+R0uGg772aBzlqWpIK
0QMQrdnuxIk2MwB/pc3CeUE9zqYRHLbmcQ3M6rN29aMMwDI56hdrox0QyjME
NQPTMVkRTXft9HL9AqbP5GBGWL4hlNrOlj5nK3JOU/iwVwvABUw8dcNvNm6M
/qlYqTm9tDAMAfJkfgmw9GifEKrwshx/YTVnL8yrnACfX9TdbiM3Cg1wk0AN
cplWMzjx+6SE3wQi81MsNGjrThqzUVxfvcr1NaGy8JXyHDqyDlFLWCu+AruO
R9Hs+5GBSiB0Dq7lS/JbnYzA7zC1lsINnKen8Kxqt6Ygku0NFivIYn7Zgv/v
5sz2/upSe3UR1Xus2/im8h8SjB0lKVJ36O/YFy+y5lr73fOPMWo5EmKRItKv
KEhhcYy0b81Xv48bI/qr3jFYC08cq+pLiBCfjicImsJGG9q9aTWdtyzvoKTc
ezqhNqf/b617925Je6JMyeXmg8uSRJxwl/BATLg8eG+wxqJ4goJgI6IEWstT
JxCEUtdGl13Nwh278mscjmW4NmvS6/KK7uFIN8TgHBpIYU/9i6EHfgKvUhgS
eB32AjNxQucyxC36/nIt4+j3ds327UkKlpCY8eFLKlew+nJU4wJ6XmBI6br5
qN0wPWUtMFDmYrnF4orsBNPj+pYwllEMkAL9vCfmd3Z1PPJxzgg8y7ndBKQx
nME8ITUZaxUy/GZZxe/xm374F6lRxnJfVrMpOVRBd1u62gwjjJxbQCr65Gu+
wOb5ip+tGCtBbf4R2piB5N3HqilgOOpA8DUiVQ+xP5u6GIX9M4a0JL/m/DOv
c9jRkAj3dc/qZWyPLrn5fgjEqhb4xC2TqVqiQqZC4GyC2OC79nMgycdd+MDT
mLLeCQn9nOCuH4qyzqR8ZOOncLFmdfyqFsPwuaGhzqSVwDMW8wIFESOtTHtr
TAqRoZRe/iDwPhTOxhTuPpuYqX6QW1ReZjTSNIFxnEkq9MYC/Bu0apRrZ5Yy
GMK7V/TRBYL27FV/NIMYEUhHVMf3ZOslA2krwQ9b+0nLACeOg2Dw5KpHYI3u
T/qJ4DhXaegZW8br/l9RfEvr82eVRj3TWfyiy9gmpCJlAOZdSLUtEPbvLexC
K7IBV+8laMxll0j+rHs7S8x2eBwo45tJ98ZAkK/ipS5yDFcWhNBzy4vwEcrv
U+oEKqqiC6Ze2pBQUkuRTKECUNPkx1bOJz3dUO4AWry/Y2RSEhFi6iftRRKK
dOCt2lx31fkjhx4VFSIY6nEWq/SZuvcrUHlsWixsuJF82c2uE0+gk+8deZg6
dk7Bg2/tfX0MVzlE0zwV1bGCvxbSQSBWZ4/ZYx5Jn8NI3fqdDZC/O9PLc+En
xgOLaVaN8u/W7OszCHf/qbffplntL7TciPlAWyCOzlnR+5wizwswXLyQoJff
ENQXL710gy2s//kgoht/dSVVe1Cu2+sQ8TGm08DHXGkAozrGLJLNrcQFfy0h
JaH9dV7kongyvntBUJAyXTomx1sxHW5NqnBwwTrVDGeBQv9QHr+1M9LdwbTa
cZcOhbw9FGVyaDefKz7MHla49b6iF1rr6vaRWuXJEGHOtdlkcCogeaWsHwuW
DqcoaSrTgjre/C0UKo+BpTwKIHolr24XE1GtS7tDNbgehFTLaBw2ThAa/DHN
BC9nWqJkzYufKrIT2L0b2pNWxt5mq8fGwGX/AKBGV8M8fzFispfWUejMTsoC
7t7EJ6euEh0TkfFrX+6Sz1nmgh9lKSxINBjBntzrPNyV7WGNwOME6tjWR1XU
h2CkmoEflbNO1axODW/skgWCuGiQgASE0SNqK0hQenwwj2LQdBwA3E2Xv/mW
TuT7QwazAVY+ydQzzUgWGdvH6w4OrCYBpul/XYix6nsGPPcKi8A1YufAZUR5
BUCjY3HZ6guRay9T2vHBNtrutI4N+o1xWA8bgcfOyhOtM2fYiBk7ki4Zl+4F
OGQNcYK8ZqpgGKgLSQiOfhhAfnjLxUJb8SEFYK0iH9pCqAYp/9PFwV4E8cyz
b0oCIPrzpuF+UYMDMftdfg2/JsHbI/4FmJgRcsb66+2OcBCgxRLsR4H1T/pV
J4hE+VJKwP6xgwBK5wrgUicsxlmkERQB/HwSZhJMQIdVrmpMa3I6I6dbhu6J
epjTlOHMnizYbbfOK+BcuNBt8EsdRkorpSZUJLkk9krG/58Wb0yToUKbnavy
+G7AzvA2igRQ1/fkJBoOKBIY+icCYSeHuRqdrniFpi7/mDvZR9CTPKzY42qn
ZdiLHF1eh9LbPkZvECL+lW1H86u7So+9XDVIdvfiUT99MS5ZjPghNICBFugD
ojf+vrVxTdGr1vHvoHLNcUxuDWKOhElpvjSoXgc0rkCROhyIpkScbeIxtK0b
ZZoI2hKfXrmaLfAsXF9x+hQpu8cL5GUkJeckM8YPonOWBIO4ZI0kD4vEgX2c
zLnZX9nvWOqK159kS2Vtj/yMPa8BafGU3op2K7TXWSGtHSPZspOGJHiHxwbE
lwljt0v4wpfzPX4ePqsnnrTWIaKOUNIa3MdVIbGAdkFQ7uk8MVk2prLE70LH
7UgmpxrC7AolIWP9LRVyKqS+Sz3rIsi8yt/QKWx/aWSw7wvpMHuHqp/2MTeH
DrzuwyLrHaqAn+vEwvcPdCjkxTP2BvpxOfrsnSi80Ufv7cAoHfPnlrbA1VOL
fuD5ifVMaC0TXUv8+QFJkuyVz1yB5TDRE8w9N/F0pyVmXxBdn4og5ovC+zFi
Wx8yPpx5SHfzmPm0XFR8SbQzjt56pHgsXZ4pRPmVD9oo2BKcKJTYBbhNqBeR
eCF3TzUCkJecM47m9DnplrkHKiyIeIXMieSDkBZeHfmGi8OKcRWUCzu6fv6E
JL6Bc+snnaRYgKv8maWsktY86O39nRddRStcxxhBUvFiLHT6GQJtBsFR60FF
jbIOWIz0RFr/yH82QRu/b7zgXOCcMkGPiUE1O4fPg51qdiDEijPRYr5kDxfG
nBDwMb5+h40Kg6ZTD810Kjcpp05wPG5AB7lmQW6AAZQrTuFDjPFH/oGvffCw
akMgCn+vEnLkgPSpkOsFT9EduElgpMT2Uit91JDUr1GoOfGjdJPBsjvA6ymS
rcHiYUy3K783Quitf7tPUSS3tWSv2qWZWX5iaM7lOpp5eErXEGbTMgHa4KNA
xJYK4O+AtMrKnAshNDR8pQziQJkRaUVhBfBVmfSBnbqWhIq4c5qCQLnlRJjM
NXgjmJgVIuDF9bxg/Ufl7Rvyg00ZoTRWDtWWOuhehLmiKnvmITynyZqA77f5
EIeBo6R08bOs7bUHjvmbpM1DGNG5a1HseFp0tN2Fz6/M2MzmILEO77gA8YTt
9sp+S/lGueuvyTF6KgUuQg8Qs0xxVeQCqJdWdBt4E23j8uUqf9qrYf361xBf
f3hU5xo+ODLf93nBC/4bT1MfD1jZk9deMwSLbIOr8vk1SgxESjXAnMRyMOL/
wCRWP+J84Ky5sTQgbZq7OJfJ1ITb6E95oIF4pEEGKspFFYgQpaK2C2fM1/mz
8xfY97jAn/0923KUWytaL8QJ6tAxF9g82PXOR9pHCdQUDBTMHohmD1lFAgTu
5ZGhRUG9+vfWpMWv6F3TxNxu0TqQ5DGnrr7BrnotoGS2y65flN76kh8FHmuL
k9V321dSartHAGrXZL7oG8R6xFUVOH7BCdrm8MXu9JOJUvktcrF0sC4VF1R6
8pJq+bLXw2tPl5rkcPEV3BrgfqLqPgxs1RDPWte59LBzqCAOCDY3wLXJiXQw
CGVcCE5k2ewM96ZlAP8+VS5v+YdnVkooFH3J9FLpqV0sbrnTSpZtZ/t82pO3
qiRPD6KTCNOT7mllgJfvNf6Ywe3tU+Mju2u6ozGmGapkwvR/qepVYQIpyq8w
WkfjqnQHvcz08Jjm0UO8esG5tXZ+o+lrJPSLCIlkI1AQJJD3DpTwoZdJnxCt
MsfRh0sWShDHorXH+8Ag3GNjQ47VdzTYg6/JdUrhRFoGeG5J6SmODj5C8Avu
ESA1mG7rNaNoAjizZ+fYPPFheJO4++kiUmL851MtXm/4fFepAZliLHwphstW
H1Wt4iEPsG+C1OekBw5Z4KICAeT8ymHy5ahVHKvvmILuGgRd/bNB7tDyvKeX
VyNauM3/jZ1AYF2eK1Bbm8Jsdbdzhou9fKQn9giz0W3ky/doPKeCSjhRZFHE
X0/AvPfVBeHbSUqUr/UAUGjWvbvQWMNydVhV9RzdHoQIzO3bLIcwZk9TSAv/
BDT56cze8QJRuX1nuwCGHf+xjTvjHw6vH+bj6B/vvQJz3ooeFanrRIZG61sh
cb1HPZbgXI1HUDiQ1UM91yFOZcksZDvL8cCqza9apC22oTYFuj6ECYfKQqQr
zTqcB7nhpxsQcB56QbTNbtzilgn89cQRJ7sf/1sQlG516N69OiKwKLo9G00v
TeQtxVDOHcDsV8THb1icqz/a4pue8feQubRHF0WyrdX09AdFtfN/ioGgZrm2
sDFaSY0XTygb+XnBAAf1Gt6nsYETsiLIddJvc17gabvWEyTcAmvvKnjOV/p8
Kwu2mFFQyEIbXYi75x9PuypmCV6YZLBF36IDQQsWO52Tppr6pI6dLsxmxrDI
lxVMSMMsInGdqdkOY8HnAhZzP6M17KWbUr6t+qF8i6qxBtlS/Fju0cZwA7/s
tRJ8KVyrUAwrw630HYxl378wMQ7KQ1dS6srET46B748RSaxdhCHDzbhddvkC
udCZe3ukqtkfay2hLYrENhR9d5aL4G5Zne9RZPVBAI7pa5+4qEiAAw0zs0s5
c+khss4N6VDBfbaPJpi3xOAfAUWZm+reUpNmfvS+QJOKHBajq/4Mlns5C8w+
G8eS/Seaj6l/v0KHMSi+0S5E7fkpbbFysRO2Ga3l8JOuHIU5u+9OUyhFkhFe
zJXpVPpi4ZjfpS5WAPXC3iJyptwk1vnspkQIazHb3CJ4ubyVM28ngxrupslL
crabAIpISa3fGO8JsjlhXq8jcKHOtbvLO/wuROdHCiFTNfOy7vvgqkNnw0sa
ULMlKkqYGU3/mvWzuET3mSCEPVodsNCIej47AahFD4p5KISf6a32JJXgzVFT
FjC8NHx3GOuOLS9Z3bHIfHDcHwSXAN62g0xDfzIFN4xVHzdl4b5NImq6Q8iw
V8NrwjJp1gXB8ZR15ZwtKBMwyfVOiZ15nmJ8H5gNxbP/0Q9uUauNx9qBFTMm
Jm2mKZ1BAu08tqCT2KUFLXk93DTwAzJZhhVt9qDN7bNQ8Y4n8eiUBU1T8iNt
R+HOa06xSgYgTe1k0UT+roUjoqEKHaUOfqclsZb7lkykRv2xUTRewzfpkqXl
BKoE8tmaUSnHZkAOkKsAMx7/aPQsyuDu3SKvqKHgmQWiH8gpZ6Nyd0owMIah
GfXJRuSWXv8IPY5tS1HaNk/sNxskbQ3UrGEaajOq+y2E4t2c38jNFjaglLWZ
8ZtPU4s/qjaj/HVHnkbMXesVKabfOw+om6SOOLIE8AxUt2QmDl0EI5SRBZCd
CVIGbkGp2Zo4nbkU5UNnMc5BjR/s4CTaPb4aD/M7LYcsvDblQXG9jsg52hOX
EyfIZTL6g3RKDHW32E/OBFTDIi9dNaxxVFD0o17U3/SfGj6mSCMe/ZSLjHhJ
KIRaj0GVDuBMHZa8rs0Itm0CxK3fpcSqMeVPUw0np11rIDH4VrNVjXDk56Wz
PJbc5wCTqOx26wvvIg0KnnID5/8Avcgro0uUPNtlc9DFIlCFvAVxGj5Cp0T7
9LDWxtTLmDR+cbM5ItQblCDVcOXrLTYcsUg/Z2o77zvJa1NJHF82dwjP0MIf
at8GP0VSpTIlGLONPZ68b/ZwzNJbbGzoAfhe3GFaLkq0q6OHAnjwLzEnMuaj
cw8BodUVP7wXo8gpbzLLSDXOb7o/9w5q+l/dWM6Ko+92MCJ2VevVjtU3PUD8
OqNuYc0K5uy5sAKAwL2amIzBcgI7BFYN7j8Yk09Y9ZQOeGLLif/wTXSHiFHo
x5zde/IQeW+35krjd5rPOZ21jRPW++ZBkQ7e2ZOKrLq8stzc0oIdjQieIdjc
fYpb563fJ+tEYT00uiJk6KzTByLnMh9eAfpLT4TloSShlC5ZQI5Qx0/Ls2vy
nelhRYxTJ6WADsleNKy0ym/Fa1/eVkovdhycWH/Y4YOhRS8qzheWoVXMMW/L
J61ouLamvCm8BXCLxpVVwfatGACoTVBt0TaFk53wHJLHes+5OtT96Qq7paP4
gyLZBgjGyXnyiko84oSJPkrGQZodN6xTzXjgltGN1/0O/k7rNpnfFCGTGzgV
hZWIKZes69cZiCpOP7JEmKC1WxwzBh8c7nbRM+SvwFsP96dWK+yTPBSKOC1t
pa+u6yMVQSXyJAyHjapS33ADTYc69jSP6ub3E659DrtZbB1hFk3w/vWWfhQq
WbvMKsCeWFZOrHYfVsm2Jr3nh4yxYj/Qz8X5HAqhJNOghkBtYWj+I5xKmqyQ
qgM+weSInhr+KYWZdnCJeCp1Z8s4VFXrfUirI5+nuS7ohX8nJgWzxzzbdOu4
b8b9WnfhHbdQaeCxbs8hpPuUQHVLDPuZ6KaZD0MML9YpTgnFp2sFuWyuvCuf
8fk67ZYAssdqYbpV49f5rROXfBt134RUuJPnqDXL1PSX9RZOs1Sm2itoQtsH
OXuD13LX/JO2D3R2b7L9+BkzHFfNss8begPJZLnUbAztaDGk5JDTzlV1MhUQ
7xKjFgph/UGqBNBRWFnyhLj9Q72cSyZh9yJFmwc42VI5uPwFksfjXRJHP+AP
zBobro4Yrk+cBUqwdvn9YGImsWQgmb5P7RUeOHEgHw0uOKTFARLyvpEDFObO
VGP59knsyySnN/iHhYNCyb3VrDV4u8lZ6RB5nq41mH1IciD8kyCyP2rFtwpV
UzrlBPwpoiF2Gsi+nRFonAhNNZZOSTpAykZHzF5tslzWY3ZjvyYLYJlIKtHZ
vMDRl70ZpZyL06JyjmdhHHaq/3MHtWrtf/YTfEJ8SAzjFjKQ0G9eu75IyIm4
tNBak+2T5f4itp1k+zm5Dzfeef7Om1TMEqv8ve3vMr1jb+kfjLQxC71OoFj8
zKSm0brT+GPVNCtL+piLvb8hJ7EyzV0zoeztM1UmDyMPWzNkSW7Rnipx+3N8
MKIpUp12jYVE0tKOooJYd1DYsEjEk1ESCQQBekpJ537OkwaMI2WPVteNwmJ8
/6JdhaO2KaANqkrI1l3hGs0pnjuLZaNY5lrkv77z5EOkG4KT1zAkijc3pKLN
ilVlPgC9dTIxKQDi97ChYlgeIKZe2ETzOOUTXA1752d6ZeQ/HALrxQb2BmBn
42BK0DAnEllG7djhEfdbWZC6W7oJBA6zRJTNrIOrNRgA0hDK8XN2uZmZUpxG
Azvdgq3ZUyfd7mtXYWDlSE+0/NertnpgAZ7962bkVIVU2gW40fu56BzUVv+2
plP9lgb9uK/vP7OBSewehdKJczdbcnVQDATWv3tiQxuHKnqOVOu606W+6rtk
mYSRTegVSgHyAFQmRBQnNipyt87ltmk3zE0ynQRR+pOBzFDgv4vTe1A8+mmB
mVsL4c+/QjbOB143EnpivGLj6yL+iVKVg9aiKr7Qszk2BmEn3IympqUnPULG
7AOWHsLJFhINablH2aL8Fqvyk1VRIIBK+HkO/lBTybkYf73ZGa5t8mMNqHUR
JiWoFAYkqf8ssV2S/S6JAn/0kq9jKh03z7NbeerBaXv9eGrFdjAFozyHkKTw
g2699CqFT/MpksOxtPGccQCn6Y5H4xOXuItJw83C3KKr9HLyl4RR/2rh1bmR
PRW/A3aVGtZcKfJQtZWDWmTxG+OPJvMVn/EajSDX8zTuGGMpJtXPu66NuKNf
mRVu7SAQmC+WaAkBYGkLOJS4p9NQRKpu7Bivyr67HnTX2PoRh6D1tooG9U3v
wZMWn9qTpcziY8p07394qNCBPKUDxdoUy12g3K3UBuAJdMIaNsx5voMlJwKD
V2jldENgQT7OqPy7YyUCHtgpI4Ve8uvcQOWuMD7T6+ONIRBn2IM1TbfD/jb5
zdFXYMgUY2397tem4LARssZFJyeRrNaGW6opxXVA0wOvV/+nH9FQiKdKQphT
MIq3MecoSmxsMr00DT5IiITtKgcbdY9PnyejVSmz7tCIYsuHbDKGYdnTPfgj
FSdxYAz5RGFJyot9+ckmGdQtN+d4+PaaaUoHN7St0D7jDZtqSb3DS/uqGwZm
IzQq4ksoDynVBctq0ILsSS1RD3Ex6OKD33vb1SKekenxLaBEVRyRaoZGt3Ob
bjfevovi7oOCvHPS0/YwHdkN+oNqPRV3TrC2wD0aj0A+zk/bDiVq1zUTMEWi
afKM9Fe63HXXUD3MRlWBVyPc9KHeYHpunJYMIv4phPxaxpKwUVMWppRnfPH7
gb0OJu8EhANQlrGLRQ/Uk4IU9nFy6odvgDv5Cwxanf+4W9lTgT1AKHERgu4P
GFX2MgUhWuGUHVXY0pib3GoZjD+mmla1KOU9lrccMpSizTEJ1o7VeViBBVsQ
EY1FQO8gzncFFxBEJaCpfku2pB+Fz6n8njIcIsxfVYonvF67gW5nZk8WWLlt
UAmj6DDNCWUw4W+xPAAjzUMjFH+UeWA4qKlh2SuIigVFOwUH6saXMguMqyuk
03bcgPK2ESJ2rmOymLwXlUlo+arGHCNZNUs0JZAlGJQwTT+b6pb7hnBh7gpd
m+qg/270L3xwh+aJpIbnpv7M8qs4+o9VD4udYL9YbwH0qQExAJbQZBOZMOjo
b+14o5a4VTXJUoIVyAL3vDD7Gxh4tbH1nVIeeRULhiDjFHd5P3o+BC7OWuf9
7uEexST+/pi2ZPHy3/TlAvMM0Bt/G5XdQl+qCom0lDG9S7wv/lNHwKYWCD2O
d8gw/uIpm955tHB1IolLiuIsySMTl+3cI0YWiTHYlE0rN54qc/C8MqnSAhTd
NkNCynZUAVOn8O2vWyxs1ii+w2j0C4B2W2IzGjOPJW4Zii00LUBopA/q62Vi
oT9LklnZ5xl/wraEVvKR6yBDxlkZ0l5yqbDvFF91rDy7mndesdn5mttN8qb0
Fly4aHaxstWAY1R2jU4j86X1QGpfvjdAXJHNMglBJVD45ZVqoFx34f1LpbP7
QkUz21keL9lG48ZVOtgfo26FJ6X+xmeiACReUQ+w1D1A2Xt0b4Ob1+WfVWXv
NRUBPgdiY1CNO1iD4zxR27A5u2CcfHNFasiSMz8QG/kHwf2zr3KOIwGm+56Q
C2Vv6HeLFD+Q9tQQKw+mcci8SKYxBH0Vn9soQIneZA8jIyx7zwVS1IPuoCBH
UdPe2URDWVJmxajxuZ7N+aMT+iLgVxY0XdkFbdtNU3RBUQsBusMaYZpNAca/
j18ruX6FeqYfWnmRlDWJLoaY+ZzPi03/hIQBJqtwqFIqlbr63DP54GsoCo25
SM0xtwAbRjY8cM1Yn1NC8BCVhZSrhomBkbPiiAUu5KCvJMEB17esWo3p+zkK
9fn/STbh4XhvoBonNHlBHScc8pYnCH4nOt4YeXvX5kE/TI5gkg+Y2apX6fbo
VXzGqKXzgquuMFRnn4PBTzf9n4by9D9FJgbV4iVXAotvxfXSvJkFe3zLzeHD
3okNeskHnqZODWo34GAn9hnqzOpGptaH01y65V14wD6A2BllsyiA9Of2Pa7H
DbWFCS57d6NS1xsWDQewezuoKzOuMw3p5t8ZvJSOSYz1pq6lXDm9QBeObWmO
7vi9auH7rw2lEPYxTCTvHHjq+m5ptlUr0XHp4NbJjwkBZIjw7vcaYIdzDzAZ
dbEa8CoVzSfLRlMsmsx65jU+cjqpwFIhcd0pTQeC6y6LN09idufX4i+dEebT
MZOCH/E8VdCLo07Dak0lDMsaUvsQMGIF3MuVI151GQ6ztp3wYlbENZCckilS
3XDOTh3i9/0KPZDotd6iZp5Zw761/SlZKitKSpAVKNR96wG+EOGhO8LM1Vc+
IhpxFEwYZy6aPhhHVmZS1jPECWDmOt3RH+0FY4yVSj98Z9FcmdYKRYpcvKCU
3DVQhOK1sePZvGhxjqB5xDXa4aJhPwJ70Ii/LvOlWVmbV4KJI+tfNGrshUVE
vk+wu/A422S0FZn6YTaKSJ6dtFqzDw5z7gzIUjubdBMaCyAZ+KszJx/Xr6L4
sB1bgDhgtOhBnZyBQDxThEAwn6XBjSkCM0aoNs+3KZe2zHfqXFgBNXslNdr/
fNYPD2OWfV9xYsiqsilpsiuoZ8mRmoa9LjK+klQjE/Ml/ORZBf9cmxv9QIRv
GFbgzYfkDKMtCUZe0xVGtagyS2t53D4gXDCP969gmx8Ih/QY/mzj+tB14R0z
H2YhmU1gdEwYe6WIiWzeHkv5x2uXD30WVJyN7zlGZ6NDXbaj+qkdPWMxptlA
N8YLidVFGp6zGO9NNfAe/n3ALrUvYrTaDvk6N+04PF2oK0de6ADuHYRDwDA3
L9v2QPBL4eaufp8Dm0bUHy9fKA2JVCK2KTLGD7w2QiVXWNYsZ0ek0SQ5UYQF
V/ZavRRVB5OW+jch5rm3alOSs981ZWSx6JhDglQYMSW8iYGxax9SOBbGHeDm
Y98J3ZGJrzUBpV3S8YTviMoN0VWtt55S5nrctSKzrSzX18zvPzl/SZ7kDlJt
YZInewgw+REeQqSXW7T98GU7ItkBNud813eZHF9I5BksDy0PGRtrbEQjTa3E
fx43HtHJ6xa8bGJKOMRBQ+10g01pDJ73GwTwcQYMj18KkiAe9Dn8BnZC8V8R
sA1tCP8wx7YSZjABWjocsBUSt3cukdoeYpyRGia7Rmq+4rGY3i6DsA1XXP0T
c51lnK/Dp5x3mfzdAEBH17wxSWkwF2Ttj+g0OnGGzd6zS8csv1syb6gSyCWD
Fp1TOf7uLYXIfgRWLZmlCOp/hEBtNnCRrXZyiDxbYfMmzhqXFPrZiugjbmUO
rQjlWrHAAZak7BXi2uxD/KgTotTgaiIF6EFT2xbDP2GVQSUwJHRqMLGcEgf6
AnKHTEiCBMpW3uLGLimYTW9UMOskdRGu2eR3QV8+cYcj7BOGkgw4qlwzJXcT
7fmEUux0G7unNj52PhwSX1t1YVtuAZw9Iw/lUKYJbKzAkHKzxtTc7wIWS8dE
ZGQ7VQH0Wp0iy9ez0HT6loWclWLilnjBFPOnQnmGIym+NT6d8tBflZLsKgl+
6z4F5CbhoYN1Jz9uoRIrEKXw64ckfbpJBOzAatqmOxos+Lu6U7ovCx59pBvw
EsLshgguTfJf0wu0jI+r+dAHKiJyp5d8DVUp/NHxW4d+VutwZ2wkhgITFD1v
wukpoUTkewcVfU0KpIFMl+V1oQcfXtgb3LNB12vNtffAsx7mtAAH5hj1IDPr
R/ZVTBRvfiYFaMYvI43EZeU6ZEyM44+vZPxd3Ty3LGBDW2Zdnzm2s4+f1j6A
o8ieNs3wNhd0QgPoGHKAabuMM4ecLDak0p5AFOW0GvR+ry05vlJYWyjzzEie
xPwxFS5ww6t9NAH0X4qj/F3kXoRGdgjCW1MgBc0NXrWjGUqea4+WCQfIsmgL
cyRqtha2mEDy365vFAiM+OV2liHorzoV1mzoQLiM+QtphyHnDAV5dvpGJmWA
hSL/wkO2xYRPQNgA7QVWn2P9bCJLstyS4JRp3e+ov6LZ2hCPHwCy0T8OAhxG
Iog9uCnV3xbx0M6oVCRKrZ8atNvHakglE9aNLZuoHzW0nipdWQ816k0VPZQN
wYi/ji3bG3YHz5smn5CKg5COb+uwSeAq2P3pWH4CYfxByHnsobPU5T6pqnT4
AEHQiR2TnYewQzB9w00gz054gNSiPC1c+7ZNSsyxmXQpEnsJ4CaJNPXvojEZ
lUOvn7y0s7HYxt2INm2f1Hnnw033lxqOp6xoHwZvg6FJAEPKfU+JdiVNs5PF
qqLsmmjtp4K44D9/NjtrxhZHZQuSbnZtpUXka6kZ1lMKmQ/kccSwRdbowXKz
BLuvM7IqPqW9jekbccHwaNLLXIUeSGn/q5JP2Ju7+LQQFC30ny4FTvTScUle
laqo0nskxqhG8GPpLADm/V2m8qPRJS4bb4v0WHXZcN7vp9I9JBVw2EklebMd
dQCE2tG3Xh0ObxDTEDOaqXb9auDUhE8GCPbZ9uLJxJ+Htn9lBoc/gfN4cqYD
zf0KlLJMOLhK24P5qxCpiRppeRz336LOTsCVISXD0/+wm+/ex7PkynxWsJiM
AR2qWKRZhcsUOCGGJSpi82JcbnFz/lPjqWYVFqTADSX5GzLpXjwYeVqUsBKt
OI67trjABsFLj/0U/Y6+LKuWz/w+FdQ9B4pqJwOfJ7V8vYGWLdDGk3PvfHby
2EiK9hVM5CfwxKDYp18dvwvtBirdxTa3oD28XB2qgBfvWZhKEtvVPfdb/XrF
SVy/SEQ9bbar3g+W2I+DlCaS333jFhRM8vnZTbLyZ6CScpmOzvsEcf0JmX3W
8u2b0SnDp6RvlNwi20RnHvXxInUQSu3frvgEvRWlaZ18tsLj4AL2BPufvX0h
7mS3UX7Q6GaxRTy+az2OLxcyV7NhQS9ZrX9qnq4x3BUUnSTbOIIxg1NW2iVW
nuDse52KXHqktvCUhmlDnU5GM5MWpnAjAOjPRPhzNLk1AGSPxMAHpx6eT2Bq
aAfwyc/zFYO3W0yECsWYs5wOWiwXv2ivEPkYI2kcLWYdnTM0JZn38RZi865x
joRR1XISJXHIu2ps09ZsujEmUVSnReSYhX29KfOba4eoAhnWdp9ZTHMiIb97
3v1iFDj8DC0pSaIgijSfodh+S9T44ZYd/JSjub7Dv6iehIX8EnW400C3nR0/
Mwhy59AXmmqhUpGpJ0XTyCpXIlQStsYDz4Uk+bBwqHaKMg1fA3AHARs9Biup
3j67FFzolvPi4eA54Glb2nSq6q9YCnwo6sRjUZyMpmiPDesBovcXiiiyJOKI
unxW0xqaunoY0UeNSbZC8s2YeIM6SUO/09aNsICHuukb2QTcYvwlK99MZiaN
H9/ilHwNBBzrYMWQfmx84ZlGme7xDBr3xq+HSNImIodJro5w6aIy9iZtLnaq
MTvVUMhEfzrZTbSAQn0Qr915AbmtYuoVb+BurdM7vSwfop/O9Ro2LeNaOcPC
sTeaWZWJiwi/R/owlwXS1jWROtyiDT9Jh/m0bD4YPlPdlgMwya8SsNzJcxhM
2dHsG8kyCspBLFTF3ljEsZm9pkoXTRUgD55QRuj9+67vDTOS/Ygtt9N4sFZ7
0ydbIc5Ft6urUITZRQUVMeIbdH8j8/w4XTR8b/0HKoVx12NksOOHRiWNy2Wt
jBqN6JYTnlmzkp7tqA0KCTGfZg+vA1/JDo/RAhgvXSS6reSd60wu4GnYEIpU
bZUeHJHinh5k/NDmBMEeUv4c6QXyiASdfg8xg5OL/3Jf5S6brKVePPHYkaPW
70L8FWX/pyaUygwN6/azKHEUhi728vG8H3i2I06N5x/wflgHOEUGW2HMhbb0
DMaqAtY8GU+07mLz6f7CC9xoBg0vXiyehz/+F/mXkB6KE2Z63Ec9+t8Ebuua
JyYN0n4g9PS62zWl+KRQCK1IrDst60lUuP4WWJognOR1h54MOrAEL3zLK1dS
rO84P3aU/AVmmbdX0BfrZPqZCqkt7ehNxEi++8WJYctQ7E7AHZikfC/q+WgY
koy4zLt0PnANuCBZXIiJ1JS3RWs3OFE1+eEAuzWEormMwXUOImqzH5NBZn8F
OFhhImLcmDuWx81tpGSxOhXrSzVHpFnLTd27/+xbhbJOEEg+eyoRomeggPeM
ha/4/CZeXkmfd2oggRyC9dprGX9AITBLGaPWP/UtaXBeAPYD+x1n32122mLU
PEAs5Kw0lzWCrPbebehoO1gRAAzzeenqnctEsFg57YFZiRebwr2LtGoO8RLI
whBuIzuZDvhspb3sx0BFuYwEA4V2MJHejLitC6nL48Re6UKfGnvsc9I9DusF
91/ihcQS1wTT6N3w6QbznM7JFsUPgKEP07XUBri9GvR6yJgi30tZM2lJNkO3
YG9n+dPxPhhjUIfmyu8l8/wDSm/FIL6F3Dq+mcP02kRrXHvrucynja3KXJ2j
B/PllF+G608zj4ypOZoC3Xn6eSbXvb0GDKYUwqZ60u4McKBaBlIzil+/JRL4
glexYLesTnGvjGnCbFgdeVD7n1r5chc7qA0dGkk9svzpPipoqJt2aeHVuVmE
2d3JFrgJn/e/jkqK5V2WFKk2YRRNGx60/Vws3LSDrsJQxIjDuUtkRe5+x+OK
ccc+qmfYIItUMoIWfSd9dR2FgPeNfwMQ79D/w5xzqg7tA8TgmX8vbw805TzP
P0yfh00ysMTOI2qXRZsVdnOAuQ8E02TZwwmeshfdXqSEL5PDMFP2NwQb2hkD
jJND/sEwBUPMTP9oHfC64tOGk6wlr/a1KOZgyTWWlSrp4HUPyFw/aGHjaayS
1fdZ5n3vVmVaXFUW7cg/V2Yf6Ij/vygh+/oxn15eBXVFRmvUgGKe0Tntpaya
GqpW+L40LwC/tPdzAh43ZFXMyhepgpTkkiEkiMfkTRlfPNJxTBHsYoDdRz/N
9RmEnkrZ2ou5FUZT0ogj9zTfFMTOAVTx0r3nQ92JOKOVbP1pqvt1lReBjBW5
NuPUIbvL/xlwNjna+c8UtJKOTK1Tl/1W3Xl+eARfKcjhNO6qOh1VUFkH79vC
EVQqJNrHR3sxsHcEHzxwr4gG3WdiqKjxBMTMLpdQZZTS5xxl2N+IhZmInnK0
UTwLONYIUEup+Ao8akd4iVlMmHz+pKoqPLIvpvVEJcozhQ6uteBwv7krh367
O8qUZFoFt+DVj5oQLC2Zka0/TS2EVbgkHhH7TPP7Z6hZbQJifB1Npr+8WJjJ
HORDR1OulKAJJ0aj1cD8G+2XXttEmyNzRP4DFao7+Fnx/mXWqm74k7q9mIrE
Eo0/hdn5kyyyBJjs4mTt56rlxXA/zSDNbz6ekJCiv7UnvqXUer0WlR72cmIO
8yqphuAwVygMzjFK6IMJ36cvPVtqs/M/UURhVlVqRPY85tUyxVt2TErmfqCR
E4RgdvIyuWdE8o9hhIVs3FEe+tkgwAbXhj+jvU9AQaOS5f48kyI59f3PS3xG
xs/pdyzJeqQq4by785z0UXM/i+GQuerEHaXXk3VZB8b8gzQgvLF/pyXQencg
ZrkHbzTkRbw9dVGJFDtjhQuXRg6RIzcipL3RYxVmGrKPShJwlWsaspbnWdXP
yNezwKP3QA80wqdQylPAzZjkYz0KllC266oDZfe5hjU5wxXwrSqZAW1nM7cH
YrOCeh3y5LTRTK+47XvB3A/TUEefwWzLevNu+suGb16KMqgast+Yu3O9zPSI
gDQMWUNiLzhtSTJ/Cc7tDQ3q9loERMEdiQkuftYma34ywyQEXb/Py8st1OI7
wskPudhpZ+My+PFJ7GVFsNxdiHLBItzbyPvWy4eUwRNjrLnJFXpyM9me/xPi
G20D5bQIEV+ejUHewb0X5cV0wn3yyFsKBclqgWvMkV+eYth3Sa4TXVOhW80g
sq9Lb8QfZFpWN1SRrbDMWGvupgXJ9IG77cE9Vnkg4gRdnS1rjikw9Mbd5BfZ
yxGi+7kpdN56XyFBe7tx33PyDkSWD0Q/CdbqzTB7MBbe2QZnb2Lf8btGPsTX
qp+aQzGmIehbS3WjSxZ2kyyRy0PcfrSKCifM9z5rgLZuGZ2m/wZDE1UFpmaa
d7vHMJPZl391tTnEZ3lh1f7b01yWNR8K8Nme6tJEcSUC3YnKMY/2Nhv48ZLk
a4x1+l4IwRPE8dzX7Zcq5wPMZzQUl5XeBnPrAb7bKOXKI7ZbApMkgDZCQXSU
IvNRQnKMQ4yOLQS5LehNv+Tm7ckNSS4NEEW6ZYtGbM/oJlevAOBIcDXQFZR2
A1OTV8c6/d/rbO2sKGL58G9oeO40oE52e6qosFUsgvnnBSoEdtRP3Dyr04/A
tpppKKT4YxAJamb+ttpEesVJwK9kw8ym1sVkf9E6Z6CoGKHdbrH4K0YprSA2
sU6JP7WHY2ydAGkKcEJbfgVAUQ91CdBe7tmenNQj6I369E7g92rAZD9757Dq
AXO2xHSusCwMxkDoMZnKfTV2NhPGAovmpCohvqaXXl8qLY6/+2Nyr4+OfI8z
O/IBLdsTNyy5Td1ViB7QzAGxHzac2kIdhICYxjE2uPMNROeG4g+AL0ODks3Z
J7dTdjMwsPXCMXfPozf9iM6i5hIHx1GvpxZ0QCnt3h+V8tDiNSEVTOQkVA7W
tts7iTBOTEjFYUWDlZH7aQlwIYRy4zz/mwv19z1cEt7G0Cbhl/gDBqJ2njiB
/w0jT0nkh0EuxZUy+icoHao3hmPnJUilwtB0cUL/f/gpcQG32lrdZ/SSMa3t
P7zjoFakq4DgdL7o7TEvxZAARDwJoum0QLQC+0y7roD+JVhhiQzgf8dyPFWM
azto/XKguxIPl+vFkGJZr6jF/uhgBdjkQeygl7aiTN6u8SG5gtcGmyQXkpQV
x0gV+c1mrGKRJc64Qgh2PRXAEgRmoiW0pmPrahh/BQJube34l7nbkMXWMwMJ
/La38j6l1geTT2JQomRI2aDGejX3MMLerC5K4IMbvuDvzhtwTVrAG9072dAL
C71YhHpeNSEaXF22Q0dgkFhm0gHauRicrQIrF9PYvTie1lsOY9/YY/kSdd5s
6Sw0V/mWTFUfFQdajf/k4HiOU3AuscGhwQk64wB1srzdiqyLOj4w8HLJpwmL
g5Ot7p7jMzMya8+J2ZDSvNteQRscPGg+muS5ynd6duLuHE4bKpjfgQ/MJur3
mM7KDiCdP8SRRF7sn2UGskXB/Ous4ZYTwx596sXqiEkpsogjSsuyiBi9KHJJ
M54Y5/xSuQsx9UXY7FPOc+tDedY71xN1NkIMKhCEAXzIeuBpNcWKCRM8SZSl
1DcmHbJoFXGsA9glQP+7r4Wne12O2g7l58j1xvig4kxh3pWEjbGNJDwVPL2V
rGDXyc1ifjQ8Nvz09qmYwv4IuJAIJCPwqz+CiObylCy6r7xMfQ5sdFrF5xet
mKX8S8V0EJFb0P0+CQTmLyMBMjV0bq+iQS9nUI/Xr5btIKhUsAVufLruuHJ8
6gtjA6VqnOJ/VXp8YMJlKjtxs7EBBVNE+vLATrGw4HM08CvH4mDkmGC/Nmsq
B+NHo7ISYpKrwC6ru5SN0AKKm/jjMFLmZokYeaEfj/3/R2V44q9vSM7jIn0e
7qG2YQIhsyuVDUlqVKMzOB5K1D6FKx37Qk1uowDOALnXjVghZ8oSOTHLBreV
lox4RvmjlELl54bhcNubCkGZWBCgNQVllrc7jSwholQRyx2BpQsv5EXAMtb+
1LDX4ZInP/QpzLrQxWKxHZQm71p3lvvd7tmZbw1bKz8kSkCQ+NNaiP5NMP6K
WBl8gjy0x7E4+UPSqfdCP94OKBXXf8tcWesliETgRD/aUr7aXtMc4JMlgIJH
ZQajQCPZpxZIv+Cj8lEH5iplvhJpZ3C7EAfdqYr9JHtSid4czgnyR0Ka0S1i
qMHgteafuUH1nnLpTRDsgVLEC6/iLzbb0JkIM/lAaXbWjPTknY0C/r6fuhm/
EcYrnkojMbnJHKk+6B7KIXuDGH8T+fZ1VuSkdNlxlsgEziDdR7MGhIGKErj1
+fCAnY7Vj2g6Gly59wVsHkULGG5xsTtxcA3mKWKjxQnASW7wMxWjihh7Ez4c
AInPhq9acgYP/LPyF5nbbar7drg7tYH+IXWPkCtKomssabmXkxE8pS80MeyB
sxY/j7m2Y+2ojEvhgtr0aDVZWC6Sn1uYlkp2pPeqfEJZ+/vy1BYFf0EcvoJ4
H+55SFibzVjqbTZlCNppy0rHKyvAJTyaYnzH4f6J7kTSgEpXLjRZZ36bZgSQ
iqu9OOcRvfzyKWk3ink16x0RsDHmvVBb9PUM1ImNAsayDvEcsKHczi4xSUBj
M9RWBGXeEgjliZX+kAGZ8cjXLB0o+Rds2KFE0wtqulcVhcY6iE1ee/AGVChl
uj5pYCWTQP/SZs0fcdpTU4y4esVrJ1GQVn+ZixnCqF6KeB2OyL9Hwzxa5Kgb
hASvNUvC6t1IhiWsPqb3PO41bQMrhX9RZ6xc6iqPV1YLbIYTpg8VaTP0SYBQ
Tcr2E8epmp6KUeOlnFFLZX/FFXAwZClRUzcnGbqnEdglJc0wNJ3cUj1C872R
+zp6mstnL95LGie5HY2rwWvS6PH7r8HfNKv8tVQITfKqJHSYER8h1CBQbHp3
QWgePeAdSQnUaJ3mhX8hij+IS3da5t55cLTmbQS3QmBayPvmfjAgOT6cc1KB
uNQEqfmALdIJV9+awKUOROvcIoEBsmgBTRiLBpL9fbERn4H64B4O1Us8UFNC
fAEbv5OKa7XRghe0Qdk3mX2/4qUfW5XcizevOWvZ2acP9a2Y6GDWDnzOKqAr
GbAB1skKKCdKbsw/QsAvaHkjq/ZbRhxwfME+7AThG+95YtEC1S6QvqU67zCx
QEXFX3Y6+7n6H3RjFiueK4WIvOHISt7Xjn+ZxaxF1lXy6/u5tu0oH/zsKU4b
FFCSRGDd63cGfsS8eN8KPdOLJgaCzAdDSxWf0Kx8o4X4Dbxj1MklHSkcMELL
4gzEyIL44Fe4WylcOGBQzEH1qYCXwKWK7J6TWLDA6hB7eKOks+JvYghbrqce
P1dSebI+JvN7k2kRNc09+0FpcOFOz7QMdQffn6V2PDoO3dGBXbmQMgLpHJwy
K0sq9b+CpwK+7WSS5Sr6wXqiL/M3RoLF9+MgySXvX4rpZCwClYJKAE2OfQwr
TKdBSNrSX8ooSC8SE6U067V1D0/yQaQ4GbG0PKqWLfQUEDo9fWUcMSN0gHib
MW79mt/aONDFhGH7cgVmIkUjxduVoFbWi8CShUYllyuRbm4XjsMTOR634vmb
z2ej00FyXLsIGAb3qYtGkRzcDQosAkeESxlKMjtrH0tyJmkgh7nFz0bIcvwG
hWl0h+ISPzX0779HjLkqxFbCzvGp9a+WDaIzzmu+TXz6bnh8JqC4QPDsYs0T
bBcXymOw/Qfa6zMShIiuf5tr09IegJz1XhkSmSz57hyZhTY3Gs0snx30E3PL
iZGS41m5QbgWviAZB2iLM5flkJvBUDr8XzqWh293JJkyS0wg4IWTTTsdf9Xz
H+WZinwl9MXRduhS7mqrKN4E+jbsjZZ23sC/TdzpmjgvFH2XQxq4dKh7tATP
qObAXpt8NrHot2VK+njsrqq9VOontOKAbdEb7En3MMJOVg9wWJANVPa4sxH6
f07OeDpt0rVED4SFBkjJxqb40QiKqC68lSvx3Ir2KXsZyyXBWCKVCIRc0WPQ
b5B29Ar9B/xqcFG6Jp1Q6W0f1GMiH8PdQhQ7p5pbVK5+lib9ir5bGEg/khmQ
ukPjFF5fFas9oJIHI/bgY6doiMccy00dsu51/TrF2Ec+oPuCEX0ETWeb/IDo
ZbwzHim4ZQFDwYhRW14gWGtyyGmKLfNqIsI9oAJv5e8r9mMcCGhfohg13B97
FjdNk988+Qvb3SWu3+Iv6hhyqbbh5SjerW5xtUUyfNvvSwKxvgGeFzvthiFE
B6VjLqD0MW0/PZ1DO+UTBwJxpWLrrPDV3TX4t/da2GxVklUPpMKDB3HceiMx
696AKaHK2lw4eFZOWKTgU55Us0Yn+oyfxXsfBFqvR44w9SqJd9mhnILE0sZs
oGjT4B2OgjGlgSM0BHAbaUa7GOW9hFN1YTxDSuFRGz8uPUOiwVzw2ecF4U1K
Gmx2Tcnhl23KQcoTyciF7FStWwGyH7VRYbLDztOzk7DLfDfbahEaMZ7q19MG
LKBcNRREAgAAuHsJSe+m1hZ2t8WLslmD2Z7KhBqJ0tnTeETyT55OBq1uS4Cx
3SsUGHrlduCSPPE9awlfLuOi36ed5UZQqSxKEcjSURUVhXMU0lNYfgbNHhCT
l8BNWhf0CGUJ2+W/0fncwJFI5xjDvZS+yUtXr+MJnwR+0cyeGNVEbuseEKfF
8WulPk+1NdSdXDL3nQDaGj4JfD+nR+rKjab6KDHcMb/ke/1nNkQ3C5bjSKjV
x3FGdo9SVfnubnRNZ/Cl6aL9nPf+/HAuaNgjEVuEi2G7bKr2BfwF08kOEQuL
k3wPy2TR13r86YFTg4f4u15FM17/ynQBQpCMjYNnvxC8nzRjhGstpUeFE8Oy
1Pf9ZvrsG3rVhNpOHIe9NpuZWuYNTJqZ9nj2ntWb2yntIasi0Q5fSHW6SYY2
27VPGBdd1TEIlVrfqmQcDXDHyWDol/6Wqa0xCKBix9QucOnS181hOH0LemF6
gwwhdq5BUd3eFho1GcLkOBfJb9yfC6b54Ud6bJ8yJsezcQLnOOXfCXK3ay+L
TgGZKw/7Gyt6z3MfmJAq

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1KfGj7xfQTLEANB7qrqhYXda3PfJOtBCB0pDvqIje66TR3g/kpsyqW1arLdzLme9VFXJ0RHl0WaavQO/dVLbLkqSpzuwz7wEfd0WzUDKG89zhXj07BM8mW5jg8Vgm1qTBmUsCcK1uS6y9Bv74jFyUV7CUTDAH/6kkznCGFesjr8autzoGNfLpENS912TCWrkXnXI3sRyzY8jCufYG7j4YUo63I1ty8Fsu8oQh1HR5OlQohJtSQcwdnXObpn8daQZ/BOAEmqtscz55TObTDfxqTv4WOANJzRrSGl/BTAwrRYrzhZrZM4an+n9ff2h1wLb891sJfOogBFmC2oaK1bnBVCiJlHhSOZoqxQdrve8GG78sr8DHEBeohrS+1MpuV8VjkzK/yYtBWt42VHqT84usZr3JkJJ20ubAMM1Vfbf7BnJYbdWBAbo+orpYH838UqppXkHH7hOa2qbwkPFKJ3xFT5zoPvo3PIceAYw5UOrJQjr3d6hDtHmQ1JnNTCrSIieMT0GiFX5zy5QMHqAkMhXhJ5Ou8maeJo8QLL9xiQp0ss3UfQjFx8wFKIRLgFDZ7NjSiuhPk6Pg4qKTd0CyPlvKDzSkA3AmAig7bwPKbb9/nCL3/NyFWj6aMH94d202IgPwi2jRfpuJS+nYqCcSzueo2i7d/w7JYY5vaG4xfCkOGoMi9KOCXNWy5Mb/vZaLWQDTmh8Wurg18k5HzNBZLUUoZxTnTDoUG33bLnBvTcTurWKoFdAEWQBAgPzPjYImXuCd4+L4U0C7t3YClUQZjEJNUX"
`endif