// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
zARF1twe0SufJL/aPSrSMXHehrRwMhZl9LUHfAD6lOEaw/zfPEAyOBqzdPHt
8YNTHSTB1WoFaI63kH9qWQWpAsbecjdtvLJYjogrCG3pha0282pcT/wKO84P
M6mbE6dai/9lWSiT/wcjOLwK7Dhglqx+VM4vQzY58DvAY11wWszajjiOc5Xn
9lS5Qm/xkUD5JzhmKkG9FQ0vc1mkKRyw/Ps9eLYeCt8aKk+l1vCKdsuSJ9B/
sdJzcJC2Ywyz7YxoGeAr/dRS1ZPVO3EMYhTsr2pPJ/ycj9TzB8FvhWh5eJ8/
FraCkRmteN8Nss+iMHs+ASj6h4oPYUSc/GDYptOo7Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lafmjh6Fpnywv3OnoGolCfK49ZpEFtYgy4qk3SkPB8Fm92vM58pOOv9U2ZHI
w3Smvi/VNDo9bx5JB/I/te2MFFgn0y0OOcV+06g47UxZmt/AOYhqvraYMz63
5fDzLVESpa88Bg7BLy4P36EsLo8fciey/hcl9S+zos5+SYWcoJrj/PpndEO3
jOB927H65aAtFn+j3Df5tgr487c5E8l05HOnxoxRh5BQ2XdwiWBCK3X5xQSM
6OI9/5pSEjXI+ilV6QvcOZ6X5kWLrU52X0HS/3dXPvUasj6u95lH29ODDrrk
x3fuqFAsA8XWUSt8Xi2HJuB0+ngRLxxnd2vyB8CwHw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
uHRWRLzKScHee1moJ3abvXUB9U/TOr49r85gQaaqTzXA+0Byi8wNesn/XDs6
cRCmIpv0B/hAgDCuR518qr8BxCsqeFUATvQlaHCder9jhQDS3PGV6k77lWPE
iFRQQs4fXcjDURuoE89F3afBFEp08FvXehUxCO+WMWP7p6U8zqCgVl9q+sCD
I+DG2qRhu9eE7w+YT6mjl34X0b7Tah9Hqb3Zjn5lfdHGQEyPvyXqRwZkDmHz
twqDCc384/znvFvculRbvuqFFGq/zE93RA05p3jMI0PFREPHaak3InPZbZOa
7kvT5PZe+geNb5k2Q358Pz+IuS0kA347Z4eFlKKBgg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GpS95YxJFMCOc0a8sYcEAQwS8IH0/G24o4v5GD3YNj9COgaSAi3xwrvVH8dA
wLcChLj/s0yVnXvWtjH4na2OdRESaUUMbnnSSngnbOnvVwOl8+tUfpFl0p/5
+IVK+hcSwgzt6SldsB96eFZP7vhqY9lHmDoIhXfz9R5BxqOaxhsql48A7Qx5
zx0qbkMXhwWop/1FzllHE4DxR/I5kSJzl45d52dK/4MtS6TwWBQPZbXOka1N
yJhdTtP2ll7bWP2BgXDv/ygdPvSRpvApO+7UPCwTewUDnhSFMfQ1F2vDntTE
yeslz9J5JjeWgDpPz3JpWBrptns1Qqhy+t1FkIOLAQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rT3UT2duhAfEZUDUL/VTLcW8jNW++LZVpNKZEwGT6fgk75QvTFLuuwDLw7GN
GMeAO/Nn1Vmy+X0wy3v2vvuNQK5tUc4z+tEgSPaFoUBArsnbyek1XeGHeOaA
W8LhOSlpYlS8SLRIkS2wnUhsUxQfYXlr/xW5UsNg+OrSG1fiQqI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
NfJwdM8QB0ai9SgJ8xzwaq0r2hgr37YbXJZ+6+prqbb3dXXndbtYyrLX/wEe
IIX74dquNFc68GAFA4EuRnvL10r5ZT2UqEj3KsspccBQ0hEIhLvletmGuscl
TNTcMsivM/plZvBnlo/LNVmD83vi39tFbzP1W2KYWut0WoPru1M0hNdFGF1x
lNYUPnQPFPeFXF5EMktMR0u3LDIoFDrtBrEhj6isY5k38xeJjsqwgn18uZX/
rUk5TRl2mOOchwOVJyl9OvwSsHSlqISpySaK/bdZObd6x9B3OxY4ZD4bxskn
uWU8HkT/PNsDjVxdFqiIUwtHiZZ/f+W2ckTOVpy7+WBCCGkId+y1Fu4TLNj8
Cq6e3tVSX6gbkPyLXPqTZDqM6baSy3QTvavt5kPtgJWa9+n3vyT9Bbx0oeXd
6A9//geSwz6Evc/OOA9ok4GSEydvqMTdiauH99/T7zWRP/MT0SRiV3ausoxT
lIvvCgwxYk4ig65cwpOQJf7cmFBND08H


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
A7FLOPqZ4u/bMD56kdoh/Ga0HjySp7iXWcVt2FirA2X4i5pGq107bZ8U7f05
oGGn2qYBSoe6o6K6yFO9PY3Bq9+tyzJMUeLgIq6ScKr42maAvAwgAz1wfiVX
hsMwWJsLZKxJ47c8e5Ghmt0di5YZJwSqgfDmNB2X8zZWCXtqyvo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
orBv+idmd8cYiTZyBGM7h+FXsCq9HLVFVmIHxA9fcZe/T4Dc7mnA6Uq6vfSp
K9bCRokL3fXOcLFYZsln3E2GMxMmXS600N/d60Pmz8qSwTfv1JlbMvCURALE
RVD4xCDmiw+Bw56GJLumEzXJG48dKzXgamh7xDGRKJsup8+aRdA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8944)
`pragma protect data_block
QNIEf7DgMwYfcSkrzwI+KQfxbRgbHY7/FovPHXBZ1zy4opeMsfNNB7kTnLYR
iw1rc4Ug27zPgEBlMUM5lJFGtZYD00Jydg2yS42PxAcF/dKXE777lWF4Mf6q
g+8ktsuZVwGSFjTIHb7dR4TXJF1jY91/a8HkakCjZSnN8CoVt6sojrb3Nqck
a2Noxfjt92k7MXd4mrx6R7iELk2NMNf4Ys2dJSFyc4v1IYYuOubiVyzscqnG
wcFC8i2STpzxfxHHTrzHgOkcKfK7vb8qnGYs6CfX3fbeWikrb9ZL0xVYvrBU
NLY4YhUTRdcaSjQqgeA+TAuXPGJzXRuWNCF5TPCRbegX9wkLWS48INIRJ5+G
/JHfaUFaTl3M+hqBGv2psNPMlV+4+Hl3VCSMV8S45L80mswPPhl9FNZHspdr
PfW5SuKfQX/1lFDVkMIRUH+xBA0KEvxYnpGo8xBfMn8XvOqss1bct/j2KG7c
/8Gr68z+4XUAQKI9Hi3VV15PtWRxXj3LVMTHK5COp8aCGNfmwjUr27ebG1g0
pGt6T14WdNrBuR57nlT0MXW+EbJqNAg1tSRfeufjMGnL9mt5xyUvlDu/Y49X
e9G4LXDtQFhN2qNqu3+FCe9fryKrKv1wMcIh/RUDZ00PnInpdvDDoZMoF3g6
le73wSdkDVjF6mSHPuVDr3USYnoUF2z2egAjCaEUf1irWSzRMzYQJPiZcU2Y
HhZf9t4TGJLYhFWcLACBYUg93BROYkVwM/n517gxg5fl2e6MDqnCx897Od8m
JbPxoUjjnrL0d5Y7gKi1ruqrJuTRyqNZcQ4gTi/BoYww5QViFYxISKYoVBxw
Z7BgOwHVfWpsqCEDtSQq2+8JnxRDA/WfeinP+gd5YjNz5kSM+VPzZFKY56Wn
LL7XSkZMBUgCMb3ETNSDoACqv6aPqVbkXCGEeBh1b/qPGvn2fDlGUveEWzzI
+VDvhw9Jul+wPO1tC0spCacyEMeqA5JigraFK9bGS1ET48anxBDneHk7gQgz
vq7fmIItkPMWnVkJhujFdN2q+wfQumcy0rAfu0sWFRcvuGkZo4xITjRlezM7
7KPtONiiOnqTvSTjBx/XIeHNMG8l7lcCMwXG70Foh6hX9nX8MPK0WAcleecT
Smze9qUuBWi8PLd8zPUBZt/YhAwbBcYz1wR7gMjCLNWXTHsHMf6spohaNUqd
0RjK7RRQSSZLbOfI5NLlP+qZgyZIztBIcJHtksAVKo4EPT4AIzdU9EM1tccD
uEcc+amwf8OlRd3Qiw4otAbC6xhxe0DlM3u52qzaxOhB1YyGonGiV5WNQ3DW
/pLDrkO5qiq6U5QgPElwrplR01Ner+Be+aaQQozaJLcPjS9J7/rnRKTr+FXn
8pRbacFlCIJxaFFJXiVq6vogpOaQE+n7xY1IDIsMJN1vk6sWJGaa5ltb35Ae
8W5tOYzV1VFoJiSaLja6+R86r6QA+HeyoL9CayyVvkfVIXDKLMZrWpPkhukA
9yv6BYw6RuebkbBkbSrLHwd3xeZOhjDH6ABpR1oy4MLAeChtDMEg5I46FHW3
3ouCMSBqD81pxzqX9QB7W4j7i+lLyug5S7seTy9+taFfVMfkWtjbqXOmPABV
kLEVGP1oNmn9LqSxYurJbdERd/ONHF5IIpzeu9CKmUueY9gi30t5vu1QncKH
1aqbynoLak1nk8hCh1NlB4x5Vs9ZUKgFfd4eMrw9Zys2govBeOjF+A/HtYHr
F8LIdK5LvOeyLfJ+TmNu374ZeHUI5hzPC8tW0h67gCAnxf6W3F0ayoR7iq+x
5AAaTmGmtDwQLySScYaAuJba+RrE8QTjMUQiMSn8aO1S3E90WxXI/3nxKFoG
+dgy4zR/n5HWNPb/M1b8bxGqWdOyiKrn4fnFrV2jHFH8CfIBxq7LZFBI0hHy
06rlazpgTqgz2WxlnpEH+TyCKBSTVQuax60+qb+SjZBM3a/273vAtgv0vNKF
QeDszY86E6DH+Cw0u5vt09fLupqETFkwuaoL3tVk5gCb0Fm0T2kLG7CWpphD
6b2S+EGFARYLIDNlHSRH+Cfrj0vqJjxyvYvKS3W+WHOrZOeBeLYKqjWn6pkp
UpUZxel2iSbWXcstafvFDR5p/7xzc/yVC2R55H/NZqPmIvlU/C/vnzPVf6Gb
V7XiYRWCj+ERysjkgo/ep7Mf9PSmrElW2Fm8nECIzWspSQorRsW12fG6uyKP
N6WXcJFYy9yN6akWaIK/foVM47/EzWlsXghThXNAFo6EbLAHYLC+zdvqVVsb
uuNH5GjIoJV4FbHv6tECggaDhuIe2LfLb4VdzzoOrLmCwHZfTsPmA9ToYbcx
6/5Q+pyAX7Q/0bD9sDwEuckSrBP1VRsebQiMwReYFPjoj9601GmkaXQwS8Eu
qvVm8WP3LrS5GoL/aHwoHS+kqlt9wOKxwk6gJch4XLhpi6mDQw/VWngEaBBD
3eWdTVcdnd7WXSLX+PYZBVQfltomPxYMikscngVGy2iCHn6rGiaY7Zz3dtbL
Bwu6WRrg9bioIYwLPzs1lM8VgxTD5ZZMvcIfpxzyMr78tDSnt02lOVCwIZvl
4+wOrT9v4VcUz8E7bQYzyPtr7KvRJugxesQjfKAg1w9MwBM1AX0hZo/yvQBQ
aOPr0loQcsc1bz6G1+LU0PZgHgh3t9mrnyl9llhrM2a8S7drFt1Qo2h32ZWP
VJ+yaoGWYHbUXK3bDr++BDjtlvjPOW5Pto0YzHbJ0C3aIq4wEMzstSLkXf1c
P5mp0cray+RHtuKfI7N7NcPngA/R5gbdNHRxtOErDy6a0ju/dRWK8o4MM5BA
nMqdy8t6ioRZl0gYS7SlviA/GVRa6La71ja0zLJIY94x92CTUt2n97ySUKmu
0Dubv22mZ0MXbvru0CHZ1ThdydeBiDqjlm6JyteeUso8C9iEWvP0+5ILiSt3
Gw/Hnh2AA5tsSF8Ox0i7ZXtEa4RTfTe68Vz5IK0VQfgPgVvCDoVS4ItNsO0j
Kyu6wPlu3Nk1bVwFbzTLbB6eg2t68055HoGPgzuMbPVntnyEPChgWS5zdmPH
QRyaY/rrUSnYP91Mh5MROgv5tnKXKGW/ezP0hwzqrsie2dD4GhCT4blMkEAi
JA/suEAbpZX/xTXx4HBiy8MDsCUmQaWECAyKNZEJ5UDZVD4h1l6mc7ke1yiK
rFdQay7zlZ7h6UwBaSwRi3VzN7T9k7tdUu+upKTi+OhEWtlJrLyxOAG7i5es
npJfNVNrA1/YVjw/yM+iIOMLkXJGTkC4GJ4dfuic3N6Uplq5vRVD1B5BrAJl
VfT+YgDZ0o5RNSCw4/aq7slLFZgt6b1mdL6aSwLC3HesOmwyBbdV2H8rtbJa
Owc1+K67IqIMuKm3OHjyS6qSTrnMTdXpMD3Rpx/LBCw2+NEUY+XSYR9LKDxQ
8aZwWXDAfnkDiCl3kqR0bTm8RcNIDN3ULPrUn3/8VuO57LWD0+ODhtNDMC/U
FwCxpiWmyuHt6vmOVWS989PesRAZiMGp3pkW+i3h9xq1cRe0Zgz6kdS9+J4f
FNpM+H6GC4jc6Xa2NHUGwv2cMiN8BQAba0EPaApNIhZiqxmccgHlU+AET5mC
Y0F6zaNUcjd3eUnB0oXN4HXBw12zo78uXX3Q/MqRrYHFkw6xjF3lpti7PG1h
8v6SN4R9IZQD4tKP0NqpmkhRv29Pke3C1J5L2aOy784cqaoy9BZTt+pf2wpv
mCBWV6xCycfDBXgjQrZqXQSV9zUHtxtenlZMyhC81k20TKSHcebIPGm083mu
wMJ/vGaAvCib/QmkTE6O9fMWChx87wXIRzkqDyN9C5HU2pGVi2WW6NtTtvLa
ZMAqZovZons5I7SqzbjVFVAxzKu9GnZiGM6zWkZvEEGZdzyhRSNdo/bKwSBI
6WyAzviBl69yQvx6bhA9v5ESHw62Xu7fe29zytbyRly6CUoIZABcqpC8MCfY
4Fg7+oFPKxfyXUpnP6tQElDKOIE6Dk1sqEaikJt7dkI21mkWmLpZ13mc2azl
ld66BghQIbxqd6KWuA2oeCCyIcpEmjj1L+LMeidLn31yx/sHexn/kmnU/9hn
e33CEexDySLL3CpJ+5LTVcF0qY0hk9SrT9p3dxCRxTGzPB7/P6woEVbIEH3Q
ygf+FWBC17CNyRN4RGYlhUKVaSOrSkOezuMttVpC3UdPRSV8VBcHbyllT7Y5
6e1b2xcSNPfI/l9+I1cVpOjsI3EvB8RFyLUJOgQYwF9fBRFU1aaPGKKr7cD5
fIDFZaiWr8GVqDUa8HQYMYNupeCP9uGMLc0le7UVG+noH2f9ZgGOBFfTMCNn
5UtU8kLOyOxhwzk93g2jh2/VcX2JQoUKUL/Khvmi1Xs1GQxg2yNshUChDq7w
Juz7MmNpTeAOEQBHgxjYKfuTHc6a29wI/jHJiEo8v1Rcosl53GR3jYywvHqa
jv1SeMqqRIi+8xf0t93v6SZEg2kQGIGcepopW0lIE0yBkZOEat2Yi8fBqKee
kJnQS+OQCw2Idw7Q+37HLPRUcyVoDNzNDYLL0pD8iowP9iyeYkHUfSHMkpyP
2N1eu758ERUI/q/vub/BX22XVTj4gjse1RnWw23fX7jX9z8OOxjP8oV7JQTq
irlAYFS0H/Ds7vBHw/Y4d0FTs5gpUdUY2MJ/cVs2Uoqpy0ILEmf584Nk0ZnY
XW5Oh33hj3/DKRtJLAeBL75yOTTvgWYejxkT36BLnvbIgltf3LYWMHB3Egps
XApX0LLpjq3ufzF9n2WeyWRquGgaDg1twHJgncRdBJkD6fMv6YKCPrfrJpj0
sY6EFeeY8P8RoDmbqbb/TlfpaLr0H07Oq+KKnTnWhP7eDuQKdPdkhWXzCATJ
Jxn36vzC0D+zmXgh4OBkuKC4SE31DUshfskj6sDNPuTthzqpioIym5f3SPEF
uUyy8zSALH8uw489pBYQXQZS6XBMrB4NxygSdp7aGXGR915D7hZkIWFM2Xbx
+ul8mk6/q+3/jH+TGtQCBzY4BAn0rTcw5ZFBOxW6cN4M97IGuYosYHPTt3hz
jrZKy5gxfFsZb6SEaq5MbFO+RMwg4WVcOE1ByJqliHPAKUFgPGpYmdB5chvR
5snt+BdKJlnR4yIrx9CaYwklLwC506Nqt+4Qod89AVVRxUkJRAy3BnO8w5fB
M0i4EHEEIvfTTojLbG/2RUUyWQ5fgG7nKbFKGWhjIjhgOOVgyojanxydGo43
GxIE0EdNidMfotxQX0la4V+85UVnKqhXksAO7iyj1jo3Aj0vjMQxwgHCE9xo
wjSjmLNHI+h9LfaVYu7KJSce1kiZJpwfELmelyTTygt05ppLeGSn9JzhC0+4
I1gZSe6f6nsubyeVxVxJmieBpDABvTeUbKvqE6qzvT4uMM4Ww0ZZCWes6TNU
t0uHGcrZhM7i7qGPod6/S3F+qoNLM6wgS0FSV05GerKEJsGjiGYae6+d1MVl
9zhzOY7IiN2p3S6iTKgnaVWf14K9d2YBnOyGgjIubGzw8PCHIz7M3fNYq4Xo
HGoLeHbw4opqUSf6VpdFAM8D7vkvHR4LmjkIGB8es0PK8AB4NOlZ9EyS+noN
hHY0I2hBtBNESQbvugLLWAzjGOlNoD19R3WfgB3UfaYLx46fRJwm/SRuRg0L
8/9LmtXZqlxRE6O2SlMq020qW5kZ2VJx/At0Xh92IFAcGll96R0gWR1QAWS9
22F+CGY1W5/k5d9Ex0TpDkDOmp6enNVvoAPGx5SMrTBiW+cUatCmMQZN8mQ6
PiQw6AxNiRqq+CenYVkxOsjbTIIzEmckkf1jQPLK8fuverUwGsPdCEjXX7D9
GnelXgvKy7+I9fVzIjMWPcOvgUXGKTucN1Bs8c5J8ApP+q58r3GmvNCB9//m
42dyAkEvY3KFcPPvlpHixL7Y2RC3OJlqsFQqGORlVHQwKDx9rSSO4Yr7HA+s
sZK2u3dEtnUxQucJ3RUar+U38wX68S/7wMVyC6Tapmks32tLep8aaSUzTqPb
RLocL/KvA6cMm+Q/owGdT1uPbzV+GUr3OLFSYn6SK5PuyaFZy1MQcZTRtezw
6Hng9v5gO9QbDBEFbXx+GOC3ksmEjnoWTC3m5QzMCFbOlferBDIZklDgRamE
vVFxYLHvGwBbxjzHXpzktDHPfiFILi/+jqHsHAGpYWrowuk/RNIgaDmXVGQ2
CgoRAtn4+2igzah6vaEmgGNRDlFiihdqnyP14ZvFIq9Ky4OkMjJpD2xAD2rg
0/PQhAxmzj7nSnJTW3soS8x3CYZr3o9K6xvGqtbbFMBX7JgabKg/pJhbbGJH
rgswG9S7Jbp+NHLnNKLZ04m9l2RlyIrO2DaNXRpu26Rc/CeiOE1knYF+NPnK
HIOCxBGqmVq971DLMMppWppYSCGMtfHmAVWaogmaxLQfk2zqDWpF0uxzdPiP
MA3PMoqpW1bAWYqUIV5GUwue3xEvkacMXP1S+25znrYNH0yFQ8663njMBVMV
ExunD7kFiTwCBnW2qlFngOWjjilD8Qg8lVe7su7NkXqDYc7pOI/D3QDx1XwO
OxVUYnZfaEZsMUc+kjBkfgYn6BSeS+GgZk+F7mKNDJcip4hg36aZsgHqdca9
SNCSIW+NyuYSC9MG3anRrGtw313fcP6Cup1kObD698CyQ3sUCfA+Wr1GMWVB
susGVI7DwFsiAm9jRWAXbT/1eVEntE22q0fWYe03KmqnrXvaxSx6TIa44qwJ
rFsqzUe7aPePIPDyGR1lcH7OlgU84X0Jvqch9OpKwRRPJ2dD+/+ovcU7mfKA
qq4Yc5xmv1KwBvmfpg4ab4ao1kTffRDuotVmFJ12wAjVdCelTINLw3Dzl3+J
mwH+5sn90m58z2nM2gZ4FHmw2I7v8K/e3oOaVVoZMVwR3dKHuXQk1Z4FjNz3
J0767IOyTpVzYj6lmiHVgGLj5DvPD6BqCiNxocFZK8K+ZdweW2if6cZRSBQT
Xqmkhtci8lDG6Nw1WRLJy2AQTPXTdnlNpTWpyzGHJzsdtnF65zrve6YjmL5j
WFsvXLP7I3wwzWdugH6XTK3VWfyTcmu6N2ksOQgLCiK5VP3O4Fk62M418Czv
ypYhVmHyM6siWMdfiUK7skVn0rC4e726fvmedk2tU/4OximFS83YVFWKXZTS
ZDABlldtPmrgSgzDI8ZITOwFEq0o3mhrro1Uz+VLkmUVK2B2tCg2DHVASdZ0
zChsFoCZuLN/4KPbim2fSx54jy/Sb9v2ybGeo9Ttol273JNgB+wgG8c0NGVz
pt8lYWjM10EvxZD0JRUqbHKjHTJfSsfG48/0cMnWQxG6+bB5tf3CjTpOzJs1
rsZ9HUoWTa8U30cRerqjLUZzhrrOBRfgekIj7ArZYoQiRr8MY5r8x7Dtri3K
TjxquYJiiHRavwm4VE/ozL0p2gw9zfkYS2IlFCJU1Ha1wv15Wr+yCWwPEr83
QI9NUKt6TYnBlkPp0bnLxy+lcCjn3p4QCky2ljhSOhMyWMswCMp7yaZLwvzj
LnZwiePZu2B6YFiXBs29xIaGfy5U7sN1mK12aWHDy/u7PokBljd+zJH4yHp6
S7HXuVf6zT+RLj0NSiSXsFAslOfnzkFL6ykFbnUJOCPqhIz7ER/TNSZKRwC7
vrnPe2xdJV0nCWMQeUbfLkv0mU1Oim/GwrOn4XM8OSMEBwoMaqu/MMojpvqe
wBxe04xD4JqbsUy44GCel2tDJM9dRwlslfOIAZDdmHGfvH2nHitaY9Ps3jLh
vC/rpVw5VULE8iuhxcnNXRQcKuoPY/a5MaKX8r/0rTzbGND1O6dN2SrHTBJB
cJPe/MqmoOx2qBC5iG8JNeZ1dKT3wu5A79noeGQsxMPjJC0X5GRFAPxFF8KS
1WXrhIrs/GPFfT28UwY+6HIpRJS6XCgNk4CP9llFjZKZJeTyLQrnIsAUVpNj
mlf1dg64gArDWVcC5DOPmvgkMacgW4lzF8FmQGFSxqeof+r0P2oCeZji+ijo
viJ9B3WPjZRLXYO7KsrR+n0oX6TydCz6/PHqNvfw4A72IlTcGdCuYEStxCkz
LZbq0wmQyGRlyzKGywFyfHU9YXS2cvv5Bsh7lbYh1emkU1tzHNBNmiXdc/su
5OKFuHypqLdxQeRp6JZMzc3O5U0RJNDU2e2VBtOWTfhDsuokUo+UNdHb/SYI
sw04QVK7bw1GElWctcbibRnobhWNTiHqhuPvFyyaa+sxBdfIotIejGpwe3PZ
4xsGdFYYz3xvmcrPBB0KMZ+KGWP1fYU6RaI5l9M7aLjxLoUhuPE6uPdtkVzW
dk71B+c6Y6mqt1GpUCKdPyyuPwmP1u/X/859SHZwu5ZOvprH25vtAgT97+RD
tpdfM4cObOwJgNcXnZJaiH2Iv/+WdaBDDJLyEp9MZ2qHsL57bI8cVvHWWqev
CJkobjTFAnRWJFASFA3qRLcyLVdJ4mbGAA59jobxMBgEzD190IuG1vyOY0Nu
u356m+6TTTE4nXgzR5pgv2AWvGTG6F89pIhDVfmi1N/m9mkBEmqoUlmF4fl0
IYiG4NHC7B+fc1rhx13VATIxKkSENih3b4Fp6WFTjsZffiF+wCWy0lUHmLeD
uuiCkGjsnKEF7q9TMcJX7wxYyhbxloz9Yao7IXNQFz2H8KeKj6qDKTYvOYhd
fnCUewi7XaWM2ZcG0amv38tRf1UVzFdPyjERK1aSP0jq9D3yqMt3PZPJy1NH
mcv96UocY1ttmx8nvpqCuOwEWv/UEOJ8bGQRezE4PEWqVoXOB5Rn5VnEyG5g
/SV/ep3QdnZhw/F9X00M2n+j7Z2lpdLKGbV4JugELh26nF24Lv8fL3b+zSVT
GEprzZR/4Tf0NKoWFc/00Vn44PVACTqvSIqlTpRbVBmwyhPhVMKEYyDVWz9y
d/ikoKaqWhqdwwSgCPZe3cUlY+ddET2VkXLnQgigbxcLUc7AS5bg3CVbRNTr
rjUheIPY82T8QtV7bkKfblCMvm25MSDwyvDFhOF3uAP59zbVts9Fjkrl64Tg
s7sBBoDuRHU9LtjPqqLhPNZEBekZM27g6XM/V7/OyDzY1grL0nUAgYaSH2Ei
RkciDxJGchyxZqozZ1+/vcGMrLSIPhS11LgIUkubr8SOPyKC2ToKrCZptoVV
Bz8Bhh66mXdluIafqto05PM3aUdP6n6FxtfzfBcU+gU+h3epW+MAen2LQYEo
4Ie9pmnFdPXPBuN9jyn06fxsktb7mpwUInYfMzRd9mUx5EqiSF1HaJ2AvS67
ta6pSOVZDFNyBxbizVepXgxmeqAum/paiA4gH1BmvaWU89Szdy+oTmsUKXDF
JxCDvESBLeeb3QwRb6BkZLHMnNIBzf9dt9l5aBkTscFgdVSrmvZye9jBGzV1
Jmowz/bypSTctN0dYu2cGixhYgKKxWGwx3gTShG8zhiggTBy9OppUeQAOKc8
0UhNSyxq+HbBe+BhvmSAg+bJtEojlnKc/an9TND595+60fmkSAfRtarDpdsn
mdwEQS9GMiBycImrwNJNseklItmVfMTN9lYBXM7T2zbqCSEHq8LJmjcT74OI
d4y6XfP9zn/qKLhwnBjfPsZjZU1Kv0rm9vv8s/OOmFr0sceUiAeAQmD6jx3L
ZZFA513CewqTw+H9/irlSBqmaLF/2i0c7TkM8uZECmndCBeIkF65xxHHE2bl
aeWvq9qMri61/PGr1HnJzJhxnI7GkklB7sIoiptuCTqDykNGAb9guIPVuNmf
HFpDMWZgYcxmkn4duldJxaWtxRbq5fWDgyuxEaQmaF8lty7Hrif/ZF99iIw2
U4HfRZVt+MHS1hre9WCMl7475Wao39LHkPhl47Pv8Xb4WRGEHzIUGpbqws99
V8UWAvppmhV+wbPUOffXfLzeJgPTERmnealRRJbYm6qHsZBoKXx0Xd1sbBBD
y3MdKCOiq6B9OjxCKBtmIAEdttDENzfDVLdRpkbCequWIHIdzAkMAtz1ln8n
VcuygQQwDj6CrLF1lrP0SqYW+Wf8HsqOPKPPAL4POCvxtLgzqpvJGK2YVxoH
VNDqISMU+sHXz+rWlEf6zbMwqg835s0nZ5uZXR3OrDRl68nzcLe3c6KiAGzr
VG9ylpDfd+cpMaZpsB3RO8CCXFe3NdnfqNqEX3Q2QQxwfN5P+FiYcK20YkPo
eG6B3pMSNQvB2hyXFMMszDfLNyJKPMIUI/lOURhi89ogRE/LgS6ypHizpkvG
ZlKeJOU76OASXAuhuMt739B0tzoRZcCtY42FTwy09nSc63fBBVu40n32u89D
RFrp/FZ+sBwAmNbcy0OXcUw23uCHqcERAY5eYvGZSBnRAc+Ffnz3R/4Pb/o6
RpWq60yYQuWP6eF5vRLj4yuuAsC4g6fZFjXn+LO6lrCGpuXwvDHX1Oy+fuHy
wl5yV8TQY2fPkOJ0mGG1twsJjxruiwETOhvuBuRu/fC3p1HR885Cp4xI5K51
HFl1m6EleWU9g4We1hy9pEUIu9McDzXV03CQuTy/88B9bTk4M1l0wU0Jv+xV
EI9MP3gm0blbA2GrCQHu9yC80ipzf/p9YvgxXsun6EMh6FfW7O4TP8NmE9+N
Zjf5kkiIiNY1ggwHol8BJrrZKYo3abZCZi7ZeaLmTVrTFVm++TFLH80SMiWQ
odrqzPHgdTQbmpgQk8cs++X+Sp1T0qkeaqAc5YCS63zlT/zvtW56puwGXfQU
NRUOVEUs6SFQcnhiItee5U+173+Q8HYlp2AyV/NLwwMOYBAAGL9+JGT2JKLA
KMqjK9ym0+vm8Ardoq8NAapH6/e8GE47pKT4D8JPKDKfpPn9bRX2vIwit7cO
PTM+cmIQ/T4kRiRNZR2JNTm6teqdA+qVW1SbEJyfuKPiKs/uW0PUJ0brWlkJ
Qo7vIVGF0cqtMgMc9zhFFFm14ZaD+pV7QDfIZu0CMe6JXn/yb7NgwRcTIxr2
4SMDygjgHtUK6bg2Kowu4uakt6hn3ioMDGQzutlB7PatZ/qMtLQy0d9vZ4Z5
ciJAEbyjRSArZf6EU3wqMapk/YT8c8x3y4qg2pLwpG41dQUf3We1GQMs5gne
lnpPUhZP5boz5tUiJA+GMLVVJzhfwjmLPWkv88hvHzohs0KX0bC/4n9qTsJh
+axPUbQa1OjRFD05JkGeYLPiM/zAWrMaXrAwALty50mHYn53UewOwEPThiOE
xbDDC6g3d8QBv8dmv/SioOe16BiyN1Q9C2bic82KGVmyZIQKQvJvBi0jEROx
vbp/GvBXeUYQ+MSk4pEv3BA3ppThc1X0iuUeKG9EY1B/7QnfjLlakP4Vka0m
B/cDpjR5z1RegWFt3dV3wz0D87PV6TCsTIXNpGeOqoIZmjKyWevNqVyNtz3s
s9ic6JqQNhVkBirvGcjxdKHTorv//AoojZflDKZZO3DEVJySW4CVNzjBB5Jq
rOCV+Ny1xeMxC6AHx4hzldMjomYc0BQrP407sXh+/sNcQJsgt72EUVMKB12I
7eCcz3w8iwafsC2gK69ss5YTD5i89IFFkaoU9AI9ejw4F0ulOXUCA9cNO4hU
5Yp20X/a0HuJ1G0SXsQvI5FLF/VmpWijunBzpPE7yHLH4aeGnCy26R1bbQur
We7bTqQzXt8I1zWovD9Ru/vStXx34HH70gXGQhmP1VGecgz/grRq3aqEC9Lu
jBpzpYermKQrFtgYj3I1tLJxWPXF8oFjGazys+e+LtJfvcOZMvvNdiHWQOpt
crhJI1qNtDkB2PzrPXTNdan+ricrga952+PD7WelExVas3xcKyU3yI+D+/xa
gRYCkN4S4H91bztMSOBJlMA1ty4EBJXFn3opJ71EmZstQsPsl9wVPfmtBoSP
FJjvl/yI8L2g+3FDeXSvf83snDXFC3m898wCbygYlgCEH0PSo1pyzMjaRmJ9
39gTKCzdTB7FPda9utgrJToDW8CyBYh1yRXgBJ9Kf/YIyw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpejSohns9yn4q5b9FGSMpL559o/8E5BbkG29vH7lphvKCGDEEfMLBOx2TbG12LMO/JIH+Gs1Yl/5v8ktuUvXyzNa9XhjFK3/VmYm28CCDKrYOyjYfBIqAHuXEssxO9WEp6Jj0oLmdjGCH1DxFcjcZnTERy4HLTCUxCMIFkm/tNS6JHxZf6IyIm0OGelIox4YGouZCd/F/2IcPKjjFrdY0LqKlAop965f7+BEhOJCsSN/gEyeWcU+w2mJMo30Q1O3z1YD1GL1jhqMPn1eGeXNByE5ViC25X5DNPlAGKnXgK1ncbvQq9db9l76ifbP/8ku6CS8WqovGTmFmkz05aivtyatjphPRQ55BPC01M0pmhEPGEUnLSR9DZZks30EbOIPUoiC+SajlEbCbSRUL4EaO05Pk00goMTVm5iBZDw7WWOApgC/8Asjr0wXiwbBG1WpCf5PfTXqqqlJyU3mlPXIm0xwKS+wp9BKlwyBzUXQAvJD8BMKe4dbDwD6XUBMJXMw9Z8scLawvRMrlsSbsqdqfi5WvQreKNNb6Aqw7ORcgLN6eBdciThZ6b357BmgCFx3fI4AqNde+FK9LsCZRGpCjz4LqIbfCUlxpxqlAMFrJ2ByszoGqC19JLuS+Pbk+Eh0V0mmy13ebxMd4UU9owqBJpeJTTA1bfwOG0KnehZ1zNVTomvNIvNsVRM8/ggT9wg0r5ue77nEN9S+MlmuOrb2jzVvFdOi92keg70wWVmte64kDgx42Q4cPiCsLKVZrtzRdoPB8KXtYqCf30S1DqbTBu8M"
`endif