// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
tgDqJrk9EOnK6pS69/uTlxSIauHTF/xnLzFelMUf13unkEiBO2DuVXbRXOEG
AqmaCZCRR3UOUcJFTvU8HH4vl9f+Ht3qNjAwNRJSjktvo+OPt0VWptP2Qmlu
I04eHYwguAf4sSYcZElnzWUmUpAyvPtqfvD8HLV2eZ9jO1A7hBzKQPgACqm7
clw2wIM7ZcaKXuDyyzHNRwg/qzWm82Yx8sMzYO27cR0+B6yLIfUqBVduYmg+
vAARXbaaVPdBj6URGorU1nIXC72HblB+03Z2rphFQJxqilsfqgwwzBZNO/Nr
A+b9B6Excvt+46JIqGQ6411nWSNgNeBHZceJfAwYVQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nUpVHF52V999TmfA59Sr2sp9hPhDcnGYAQ11TOQkdhV5Prh865lpoV0o+ZUv
FQNUxFiBEKMhjp6iClpnA+uwjKVLJXlb5q3xvx01RrSF3tSL4UsLkt6wZyIa
G6cCzJerpkqOad3qbQ3s8aF/J9aANdH8b4GP0fjeiCM32lhxlJXUlw0xJ2xw
3HxqC0LWtgknR/QOybaEouVO9X/LODD0rMTDPdVuNUQYBuOydwFjq7zAy2j2
C2wNwLNCDH9H2wcxvl2rmi736Rok4qkJcPGF2epmglGW7XoFJFy+wXUtMi04
ykBCbTTn6saRCJ7vc/KbaAqWHCxuPwzTnZVq2XFqUw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gkehOCoD2Rtg4MJdJGbOM13NgQvg3ni9hMHPn8+DFZWH9IJrKodn93i7bB7j
EKm0lorUUrF+WmXN5kEIQq9EAi9LWZgRoDxHQdC2pptoluNNb7n4JRCVFANW
cpDTnAJQsWmpc5VfzQqem4iPgVYBT28+PGAOTk9nb/2MzL7Rjrlu0oXUC9PX
i35UJhOsvckg3oe+IW+u5egxXlgvfWvq2693AjGSatsIqJ+8mk8lVN3zwG8a
iI/qD+LM0hlhk0oithK2IanVRG0gmrYOYv7GKxwMiSO4gWWdPWDvM2I6B4aI
60TOrRuCUcH5P00myAjQE4qjofk8rQCYbXe0wscaKQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Vh/3GuV/uM15Sv/masEwQb/ot/FKL4AHsUXMVYeVmAEJ8JN1fLNhh62BIS5/
7kKs3P1mBMpMSQl9baA3DMm8QAeoDkmWtBeKx9sGV+g4Eo04fVrfukpt1X4B
a58W5Czqtu7ZcCtOZvP+gj0mDq3uuLw5HjLtV5FhgNBQkF/lMgnh8vPqia5O
EPl9XlJD+mB3rBv08M7YOzD2s7/VK0Tk20NvWZNKZzI3go5U1OIPdDJGK6a9
shYGqV4YZSzWMVAZSjQD1ImE8GJHLtuliedsaZgX7Fg/WHwXL0tPmrJC4il8
hD9LfYA23hxvdb3W4aDGboqIGrM00CVVGradOtYfAw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BXdAq0iRiDebWixzbjyqsXxgctOmkgBshkYAKmgxPXkHlNkfqkYe9DdzkS2g
HYGw4XYwRHTGGV7JXvcaM0wSJYzmOz/UHj3+NIN7oPm9q7DrA5rESAuTNNNS
wfnsUPbScNLpFI0cOmRzzux5ZC6mQ0Zwmy17b6GHAcnsPiEMWYg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
mLxpOdidUTc98lpdpLA2Yq76jvO6nBJ7F4wNZedItvg+pkLnr7Wit83dNkQb
AUT11bwaCAkm1p5vCs9ojAM5nlptA0hX12waS3JDELkFI2+Mg7SPMe2thoi7
ORZEl9sKBg3T6VmnxYbcMlgtu0IsjAgM7vSeNZNLcDJP+dF1cjBI9YN6Z889
yJbfKgRIw31gYKZxgeHoCGJ5nQ9l7i0rXMJE1c8S+//zKFmTlX5o+dUea903
dukwhPz26l7RsRzqJcUipYUR6oGoDQfmSPAtLz9JRfZXN0AC62O2vMLZXAyI
cyVFoHovCGbtGl1kBXWzklGvcDjYoUP+EotyW9uekhl7Z8yNCSEEx6yP5XS/
gozZbipJFk6K5XGf3NAy56y7uZ7oV3lBj8G0kN8gwlwJI+OlFZjCZReUVsMY
nGVkled16JRMTtOvCODToIr/1MzmxmXDGM3ZdhjiR2exfCq65aZao7x7hZY5
qxmU5MJW7vM9TIfNuHyHinbTR8PZ/DGX


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QAYKr6cZVj3awrtG4P27Gr5CeW3DO3XVDj1c+wJV9OqqfMhl9g7yZumkLX4f
EZ4ACwYAioCXoI5/fEcS8fMTti12zhlB+i7X+A4RahJuNOaka9Mkoo+/csz7
/f2zFGW7dN0OxV4jWLbj8ofM/syRGQXwyhWKUYU8Jm5SGboZ0hA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cQX77csUTe1ntFb1p68gQUo3f4K/HaVvlOKh2p3ET7Y8DjgTQ4//SxX0Ajv+
50q79HtGq6qlLsWOgapiveeEn9Vl52/GRet4Tau9sT2BNtdqCKgXYz6rkdj2
1/GHIZIUz2laXU626Iui3LXjPcHdq5y9j5zZ/UrHD945lX6EpY0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 12512)
`pragma protect data_block
D2qsiS4Rr9zo01mTQbuSqFuXsd592ttnhobDxnHKeAVaaJJSgMPW5Ee9lyq/
r+JkwRwdNFZvsv1Dae8hIHOMs8jDkQd76gl/tsSiTsuyPXQVng1x2UxzvPhu
fH5mkZmm1uLfqkoJB83J0OYJfS7ldwOk4ivC6yiQKz0J6RdzC/AWd0pzAS9m
Fz9ds+Pmp95MH4WRlKWOw74cJNr9wP0wWw4uMAiwWtMNKQ3CnkkaLszHF73/
SLAP72ms5PMlmP+IVGiMPIZ0gjT7FN61NApWYeUYeBQSuXUfeij3Usur3ezJ
F+47YhH0+UG1+TAhs39YpgjA93Mg1t7tSbekTt/H8O+rWzOYMaa9sIh+Q03B
X3N9VSklycprKEOZGKDbMBUTnm4sVvV0SpiXMbjSrifQziZFi2tivWHfLZrr
HLvCg0TayaFfVT5KOIppLds/2LuvEjdJJPIUeHmauKw+fAhTte9GRVJgE88X
Yv+BXE2f2Qmoivtfs7XxxDTFyoN5LcspjqteL0ilEtcdqjJGjyIptr9Nk7xN
hMWv6KQZQiXL01ejzwZy9uz4HcHsn0wJiY6hdILHgIfOe9WVIquIp4quuEwi
jnmpAz0WaZ1FpU7mdz1oJE5GkSehXR0niUbSYl/cKBSiRW0g+5XNlgpXCRbW
IYqGc2Qh4lscK097R4lu53CMHZ97+hOYb5wUmquoilcZr6bTBW6V0vwSbEf7
d26idGT3zSOVZDOLehTuRn80OK+FKNxPrYj/9GNK2SXc/V8dJ1ncKMr1f0XB
mrJ2KIAfTkxOkNWfWrJ+gpaV7Ey0dEpatfzxjxazMqIjlz2dNruMvUgZ7/8g
zPMaJS/KgT/qreeFySH8REGHdPgQ4UC3tiPldaBwC7os2h7fUWhFBaHgUM7m
FDPNDB0isExVhPVpPMK2/d9pYe5M3+5DBZz05bZXw3+tt8KHR+ORFJAINYFb
lTPhCQj5XbNzxXdANVV09Op+cC3C0DaOZ+yI0KqJNMxsNKS7KM0M8NfEPGBw
XYOKYeP2/rNAa1ewkdt/llyizqx19x26Izg+nvXlRBQkZEA1vDO4+zox46Ox
3g3mjB0oKK3tSQRPsCcyqafylHM0RdEHNMarIvEwgQjLEtqZzq7Dikh/m8wf
5J3Dq5+u5VAWtXf953khiPY3437q25SFVH8fCINS9zOEM2VeJYJ8HLbSBIog
QRHk8Q8eX+HL3gsDfRVZf6dzc8hpDQYARAnVgYoZmsnihFb6KnPvuPSt3OUt
AMhi/JC9Lo0zi2VRunVP3tH70KA96CzWbFY7jBqjVIROvebMZZB3gUDuTWSW
8dURCK09TGIngl3ZBHZQWwHRNvy68OEA/rtt3LVKgRzNG5FaU28N5dxNPQkQ
8zsLSHnJAUZJhVYQlOItE8QCGqMWCjeyMuQUf++Y7F5t/I2wyPNdan47HQcb
0qC55kTf4MXwmFx5rLeHocNBja8hLQcAbvRU+bRXTtxcY/qhzJUzTLcqWiDz
kj2n8UWK3vnrr18Y37nx2JrWLYU3WiDwVKResi+ZQcTLqOtjY3h4TJx/T/MO
kNsWvge7gY26TsSYndVE1t9Eb2aaNUQxDTYr3mDOuVyqQTysHNaNlne15efj
Zr9WswKG2G1pZcApBx61lpXEsT1difpNmR4Nc9oXKLqQpASB0hiXhfZFKGpG
cf1EvmV8bZjUOA0/So1maYcL1YLLUnT2DcgvFRGECegHWkl4BoBkgUIIMbDV
AUF9ZQ8rG/0GjwJ0kkj2gzbMhXrhV3WUN24p+uC7G4f0PfkfnOA0uW++cU7a
ujOpBLMOYHL7GLxgP82OApBNtOFOF2YUoqAceC6z3rQSdAXE8URm5YrViWql
EeulEPoctpC5ZxEuUrf1monMEL8X74mszDkiwcmokokU3BWIuvc2M4zCdSAf
gEaB+YEpdK43oY4UWfk5R9/E+0bWQVkEX6BokbJpWn2ZM8idjqNBlCmyJJoH
7e+/6oL7Y0Agu0Y/TVaRELg4Aeg+u4kv4TmWIB/VeH4gkQuZV9RDwpmK4Nfa
VGuIoCkK2Qq73Ic+fG5VUeLyxevLgZmypjvcvnSkja1REe/Y8P5dq9HQcPjH
rcSUjyW0bvOkO9dBdNsT5K7aDY/fTQXBKi//yreTvI0Tf7UGML9w70nc9uOH
v7cXMt3YhTT1d+Fr2TZrJ3NfvCKWJP8wbpz1dzGe0Mpktaddur2iAID0pScV
PB8Jkn9AJP3DJ3Z4quN88DDkF+YjFFnXncDqh8zTQND0sPKOwnZWhnmRpQ5O
8JmJw5oTPv/+bX8kJByMEg35H/GoVruwBMJ2AVFOikhJTbyeV3lVWwKpSNnJ
GVu2/jsH3Tx6JSbfZ2AuN4/EweD6J6cJPDwRy63PIAJb+Jf4Xx6ifwu7K3Cq
bZ+hmkHyYNQt2s+aMAtfMIDSep4lksw/yCQjYkgc8LsJTMtd+xjVBUPq0oGk
6LBluyvWPiZJJYzlBBcsOL2Tsq5DinCkYe37UJwYdPfOAzugMe8WsW6CCWoR
cVWjP66/C8MzJEy5cAAK4hPANm53RJ2qVA6zEsh3EIt/ih6H31a2wnf+art1
zOqJxBB226FxEr5nLIanBepUK3raEhVgthITfPaGSIR2jLfFodR3xqnKCkxK
RpYzzj+yGhKO8TXJIsEnYBdIAJE7ZxEU579adz7+WzAyN0DyaLBbrCz3pX8O
7wteb1J3vWHaPN2hN5QLDXrsqawkqkwCZRY0BhT2cuijQ82KNuMDENDoFT1V
DYS8pD+BVKkE+VgDuI8VJ2/ARx4g6BRk55ie4hopLYzdpddvVdfYEehoJGAd
JOrw3sKxKz81MqFIHb9PULTGJzSZuCJLkCBgdZwEDl6XojarDOHYPFx76/4u
9pz6Q4djTsoK+mxbyc/NmS8APXiNzuezXfpRvxK0TiH30AVopgvkt9afa0jA
sEntJsb2TwghmiCWTVVSx9cyzydmO7XthH/DjJ8ykocLKc4uChyniSrC5TRw
PKgtmIe/L9p5vJQxEn4NTfeobNvClvYX639K6mWp5YTDh/E7zEPkdr1PiNjO
UfJQhvVzOVlJPK1YCYr7L5TQHgC2bU7rkHY2PVz27kv0TLepxGulg7FN5C17
wvq3GGaxSKMIzCZD2zVIjqcg8E7bqna5/U9/Mz1pPi+VmA0CYmOk/EA5gfJj
4aRWeiIa+xFN9Jv+Q37ozLzRL79FYtnavv31JDNS0MQOd1T1xc+XAKkhZulj
zs81fsCD66dvZlkbvFwuxvfiaWiMesNrej6OcJutSKqqZnKNxtgmaYDls+OK
KppXuM9GZJ5+RtOb9qYLesZsewnbe502oevz+jIC+iNBMTjYh8apdKmqkyVt
RuHNAKRHRMFdqQVSiKFdlcrHA574r5GsUI4I866kUUxmLgVyF3XSbkwauOio
coiOyA2aCYin0k6/s769ui6ZSvGLiYklnyIrOnmkQGDrNoK3Gd6DxZmRPTGy
NxUYCSYqmxWmvy0ZkJyT/XQvbQ4skFgBKd6MrtZ37eO6YmMdoeqUbnPHbXok
jKPzh8Mp+zVeXrD111XJMNc0C2PxdvzQWXaBzmMf05iTBd/gAK5KOpPde1/A
F2viT4z9RQbFnSZbsqg8wVRidkZqtSk+0320lbgPev2P+2A0WmpYgVaMdz4Q
7hjvQbDK1Rf8glL/De5qxNJXl+4HHihVAhC4/1L+nWm6QoFiKDZQzmJt/h5Z
fZ7c+2nVw4pgri3LDA9ZXhz6ygM5J/1o3gxBLIlQH7HUXjoYA1YgAZV3wp6S
PNXJjhsOx/SGT5a5H5YdTWRWrJdLXD3EiLI+nLSwJ9vuhkN1mGGrrCXWqX2H
XU9qqkIf2y5kqMLbrB0b4Tyuf5Lm4Yhn+S/1ulmRp3jEpu9jtZjeMR85KEST
eSL1SVBE8msTzSkU3Arib7hRSzjjXxm9h/kqqxXxeLCDHxYq5Upi0VrtvVNV
tPklnFevFOFPqGcq9yv9A2gqZBhmd1qsyh2KDPS6zwj1qc45UEmPQFQVeIUn
EYZk1Rnn57BuTeGMWzbYGBcKxzXUkvc8Oyo613dL6+yvxR5TiNLxwcj51Kg1
RHH3U6ccf7WyC8kP+qV9OIcJZPtL4IdA7K6wmSXgTDoGRcK2/QMIb73K6x6N
wHW+tzu/zR5cbn1J6Hc94p2UBJd2Q48BO0r7pi/cbm7PfPQChbTy+zoGjXqf
UHZCxoOLhvbpZG0y37FnVGKxjJQpiYZCmeFynnYQsj+LWQsjr2qO1Bh0klX2
piFAR2Oud1jnMvM/YNadUaTmcIcJOjTKGg3KJ1fHQi0Eee5dqz14MB89KeOb
KrZvWebI8bgGHotdaLhdmMXjGuR8eRdSvc63Hwn4Ch1HyfP+a/E9bUpT5d8s
SqVnOwS1yQF9ZhwbwAmEjLhkV9eL9Q+gyH6zWGh57nZwt+KYzaWhpDH65BV6
DYn50yYw+ySC4Uvs5EOpL3lw7yckRgum+f8oixnIP+tSjsv+po2LaLF0Bjls
mChW9EQdwakq/ehLRe8Ms5VCj2iby4OCA/u6Ym3px526ZLSCOtQYmALxThYA
S4MD6AxGc8zpi/QXz2545emNjy/0Rwro/Q4Dq3uuxz00zqgT8y+h2vsEp8LT
cdlTV5aCh5QFrm2dKFtDQUv0CtXsMqIUApnblLdhn1IYr793tRBxRy18mD4N
F+0TE7/s2cHXrUWi/2+U8QrjVGaz2yaIUniOKcGkCawbO/kGlZwy/FApRbpo
uElpNXtYjs9d3CW/JO3z0igZVfGJ+dn+qcfNaxRiWPwwC60WAjIpnF7hZU6f
M93wYGT3Cuvu2bubt6+zwEA9pK0dSGv1WQ2rDyEl7TstwIUJkAVJQGpaQnCT
AvMbyvGZ5B+ByEEYl1QIZPy8Y6GI6Uai1VDiI96AKhT0ChcQyKhHTpwcFOVH
mhaxwqvU8iKpwkJD/xNy2/gOLhhDmQc9Vs5vrAoNINiRddt6jvBA35Ejy+e8
JRmnEJbuoEYpuG4yKhUoP7U6B2DxRdq5cWR60b0ZTZawu1eIbl3qRc5LHxW2
IScgB5NIJFTV4aXwXzUVwwJYrgCb8VKgsA8gF73pzQgQy2Nhh9mDefHo33MK
O7If4oa8WPzPd0/t/WczaGcR3XHeTO9X9cOHJaQ7ZPKSfoOpEI+UCngqHHl7
/6dWLJipoIPOaVxMa3Ni2RRH+pFD9vhXLqbV0BSfWHNcEf5aK8oGccPiCU8F
WW+jjPjCM4b+C+srH0GtIuuI19oIRzv7J79b8Gc5JFpcF3TGlf6qxhrPj232
i/BhXRiZbVxYIIvyqwAEFhnKvaXrK//NvkgN0y34LnubQub0KmbMjvV8Kb3N
Hol1XdJC+0jFGEDzNtL58BeCk04wqqVxheSCHoThAxE7EBSbgMD5thuc6H9j
4br7c6bnB2XewEf6wyPXlGpnfnPtz+ffcMZy0iN2oC6Z19Ia9JNkdcV2wCRn
dLYGq6auPCEW748hrTGAvvUcbx2njjyBPaTNrTjplkuhOTOTmAGBlK08rxNj
5yZHdBT7m15ze31QmXwCux40ipZWdWMbWqyN+HzPJJrAvUVq1FbD065jBXA/
JwijJNU9dFbYCDccxbX1Sw0GlSvAktU4dpXr4BXfA1Hajut8/IWWCxG/FHJC
L0kA+JtmMrKI1guNJV1Ek5d8hIjXpVW8LbOU8K8OiY3XWoX4X8zUeza7fxuH
VuHESe5RT8Cb6Io2i939AR4MhDrAYsB4rUvhK4N1Thtgs14AoB1Iwyp+ni1l
C9r5rVUTrRFDDXfJCILg/z+iZPaAUZYByfGYA9IYVGOF4wQDSku/TKb5t7Q7
U83Tg0s2DmDTGiWnhd6vYGaF+iiwt6UfnCxB6LEUu1ySyBGSj7Qpt9qOlMTw
xQn8GOIRT3RPGyzxWds6gm/skO7dut7hmFp/yXZatJXGvF0S5UEXmBV67fxv
DD/3wPl8avcobHIHimmgEhty/uTaclt2Y8ZMYejrFC2qvXYORrASqPKdzxSo
t+taKDQsqPUwBGFXVgBlA8ZntYmaS0LVbKzfn3MUh1o0TywUIHe0QCHbWZiz
4XK/oQ5OeIhGl+bvbRYRAQchY7JptfKfEcGod7fjSG4bt6MfMHbOwMzd6QUv
DQQYYfosjiL1NhiPXst4lrgj/66nxTrmJKQmxlK9cy0F+/VOpdA+ozJuLn37
d3BaRDfNVLFnloy9hCuZvGKRRWvFXI0AX3zcQ7HrVq2mS2Jxge+LmmcAMTaa
KPo8nJPqhEehbo1Dhg/gZQFv2iAFpv1r+dkRiQ4hX1/UsuqrsAirm/B3/0RH
VZvuIDoJ2vn7BI2GYeQGc/oDqirPb5Nda6CQ3LuFcOBiCdQFYrMnQw9HkoF6
5/VAsYfAE0K0qRvB2aIrZk1EYFOYFlr952iwUCwToGpiz+7wcN5SwbA4tCNl
bh+rMxKpJy9kQHey2/+rnH/iuwwt6u9JJvVxgjck1T8tzG5P9ppjK3ZA7NWt
yDhwuG6KhDjJmnCDs73gFVkpaE6gLQbVtm0hzMrQA4xdCOOttvkxNBLIg3+I
VXgJ3Wzu2HreL9IDaLJEMJFeZaO9NQxn9BLWvwqC63To+kFtiNakm651V8kQ
0tRsVYttVlPWhHImZppnO7kHY5sKcDCnXUeU4hm4O8E1EP8VkJoQkrMsW0dV
EPIWciXdlfQ4rQIScLEipf25snWi942xs+Rxm7p9cREd6l5bojEHM434Df3K
mLikKl3bSeHRWV9eUbi2R/qPYhXvKTaW8rOJKpPwIXdZU0KX6VVa35wF+TvC
1mL3QzeBLsaLeH+YJ3xXzBQ7HRELFhTSXWmxjg3zyV+cGlbXLofENEc1JZDz
Foapuw5EvKk78BFMIO4FvrjN9HUX2/gEgHO4JUpedNIJCUHvwoaq41Ak1QxT
nSIQRZuR/1H/KgRXSs8IQPBRlBD5+gejzTqAMr7vtsAIZlPCpq2x3lZiJaiS
oFvBCudb4+U2amJqnumBn9gT5JzcFLaBC+rSJXbGzMsz9ithFZn2i4ZP1G3d
1V8R8R3mVTSkXAk1vwdDV6sN7BtIYRlqKKKWVdrgi3LYOMVEt7NlLpc28xhf
MpD5xsP3jKmEcejvOFxSWIXV9Q3RSn86co97zMALBLCKS2TpfmYuwGQEfCn7
evxnHuJFmSd+WocbSmaE6HE/njhUGBV8nwWajlE/vOAEjenla8Ifqc2Irikr
WNoanAuSXS/IzzHIwiAB7b7J5Wqh/LlvAHLtDPtRg8791TY83A55BW7i/ov5
r+Kpbe48+cjMU/UNecH/5VZ0owIrjPDNdIRJQFNUB/hRGkY1iM/z58YsysMN
fwGooxY68azcMsK66xgCVOQY7J2LxxA6w3xIcLRu8pMuIR+slIDrHTUO9Hlx
Yt6duMRknbxyTmHtS2Jp+pJ6xwaXjlD5Gie1Jz8eX6hzC4DXx9LkdsF7RLfS
58fCkNcuN7Q+44J6EmYEAjQa3JeoSNjnjjfS/4+UFUyeDbrOrW/qh/GIFbrG
VVXdap4hqdvtf5xIQXg2Co29jZRpvlb1ZKDuAbSyKgY9wdOkQv3lie/VliGt
0WC1AkbIfcUhmA0xtDq2RPDhhlG89kLN3cWDCbppGqqci81segQJFanWVL6m
v02yWuG/M7pFOHAfhAAT/ga5NmQm1eMr2XUuGsF8kl+zg+IAWtABWO3jIj13
614ocLBXVLC6QZvoUSt5pZuszMN8Z7qbUvIFG6LGL2ucy0rmyP4ymohCjr8x
o3RFxT+LFdnKbStjR2/vqiYxvLKnhWlkgeV0OerjeoPH8JycqPzinqKyUWXj
aJXWBkaJYXJ4OaF+bl3/GsgXzSdyWPxyo1HrfeUPajdIBtn4LggXQUu+/pCp
IdQ8Br2yILO45J8ybtqUxD5tw9KbOktQ7NF4J1KA8dGlDq8fnn0T1t3xAwj+
cB3Wq/snhHohSknNhYe9KpHY7NKchIhsPMIumlCnVEwbNcE0KKmO0B3436dQ
vCR1PmwYVBLnGmv+OVomQ9OffunkhKxoEGziMQzvIrPGPY6H9OxrvMlhkciL
NAfk1G8Z4F7z4XabZRoF1yPQn8OnjSfrsiJC6eKEIIT/ygCX3dKDqbgyk8ce
07D4Ip+cLqEhnh1sFEb76sR+0vnR0tS5a6kBcgznGyoKJoiI696aaRSGYXkN
O5C7Xwr2eK3xz/YJzPNpgc1TNPyHEa2ZEtuvJAzpbzQSClv8F6m2wdtpTrfk
7Dr8QbzNUr429YIAkSD/XpLF8IgS0nmi3r5O7ORsLtIKWULSGFz2uLWp0fO8
f7sfumAypiG0d2OlzjQkS5ViZcCvzegS6aHvqCAxbJI5pFkuc3wL8JVCDZ/4
2ZU549w8KlkWAQb4VnWKyssQCcXFjzI9444LPqvJfYQiO9hjD7XWcHOLq2S/
oNsMLHNsAqp7RuwBbFJNMPdzBcx4uR7w8puaSHa0iXZn5cbXfyDjptpu9eAu
qpffmGgIzlkqc/U5aEk/vrYyx0Yx8YwWswZTRylD3SrTJA1ZyO8xGGalcl3V
H0aIrJxutd4CqgI4rnvLKZHHbP1FrPnz7oL6NFPP66rEs6V7vMXJgNLu2lZz
3R5eOBliel5WoE+3Y3z39L8ZEWVBocsz0VA5YOkkoWsBYoQxVMoTtn0LKJxR
njsKvBuoDUj3RcdAUMQsn9fdSRuYXnge4Wk2KRAYxIS8oDSUdudk2wlsfUi2
sGdnoluJ2wgJFVKkaCCYxgaAF1pLMJj8CYMF95LPMn13O2IcnPlY/y2FMoJF
MrKNd9SZNOlskhxCz7fJxQ8GmB94xprX7/ihpO41TfeHPMRVWsiU7UT9ZBKP
fbVBPIkOML7KyGfJXUg5WnJeiRNRpK7pPue+mUhY2SNNhTvNC8RETnJ9GIsB
3q0i4HIEEMD5v2GKbr2T1NQrH/h2FTCRqjSYmXkcmL/xqKJI6rgGSFeYbqfY
fM5gR+O0xJmlsfMryjDdZMK0f/gms59DB/5q8UISbiLm2qlavuf17HZRetyN
Xq9uXJv4XsGP5G11Z3sidGjd2fj5lBmw0iq4D9CDY3vyx7wbTmr7ymquEZei
gkrUyj5YJU9JRX18Dl/DpDIDmKJuWzY/cjJcKhclv5s5DSrfldMLOJVqH4o3
T2PcllICQ2+vLRr7XiSx8AR+spIhqiK7tiN8aoOnn++WqvjzqPZbmxJwyTW0
JyWdrk9+yK09QCwKGahz489bHqhxGv6cQ29/EuwItifUdx2tJTCC0LKzoLPD
/mtTovDCfMsp5Q7fgDTt61iQEEsD4xPmi/AamktGnUIcXNNxINbaQUvaN7El
nEjAGXqhtu9GndY4jv+bxp5vhO/hOp4hUi+Nx8qVliL1KRIQOzKbQkeNykUp
iXZ04u6HDxIwss2tiLoeag4veB5oLRdUaeEd099Nmaf/46QRBZ2qjqs1pfq5
Ud2aRTjzIdrfvHQGJBPpIwCYPfqzF8C4M1KXVZL7Kokn6HIxRFzMhwU8mo5N
ZPH6El1tNfcQUO0o/8bLyKt95R3XwbpB1nvspBTsPTYNqrJNmqYTWdhpx7Lo
FkLRwSDdcve5SieT1K9XWX+q0QyJWge3wVxMFQbFKDcHWkh9vv+uLbjHiZR8
q8Zn+KyN+3xhl52R9E+wTHWR3wtL7rHyW3oOyfzEPTpSgFlezwaV0GsigVoj
7AHWXobdLVFCLZsVVufbaymU9BVWc4dLnHNkz7lR7PqEupq+Xocr+hKoqBAk
b32GJikFGjEzSabiiu51ywi2I8B34YKFqU0QQYlJg9yiasxi7jzFZ4lxB5uK
JOmJhV7Mdsmsc+SWMwUUKU4w/0NcdLBytnbg6Fq8uZHL6M4fkO2GANDkicOw
c46tB2xRtTvnz3ST6TkwMAMOr9esrqH8UEElGhy/4rSUnHDMVAfCKUSMIyzD
wslMiqmnzAD1fPoplqVV3XKvtn/XFtAOjEx1sXrhoVOli6NdmHoY455xHj+N
RRU/48hZkMHqHEurOSm9qJaJjRgbIh+0AJnj6jCs4DYGmGWNAfP5RtnP7WKN
mKbrgfhFI4beIOLHqaGq7ZXwvWEHkAj8gFzzWoNpPHZTunrVlE4/u7gzB4tz
ufeAiAtQdiGGT5Jk9mf0BI7kYC33+W4KQbIOHcm+oYt+SaCqYHbBCb2a1rz4
79oTMT6VXwKEJ7kMix3yrJELFBuc99sq0baqCq3iTAfxkm3AE6T7vNylvq7C
e/lawRMrsor1xf97SsQjGVSQCk9f1EFjfSVj7qhvCjdQkBe38jJjmbLyVNj6
xGcG5POatnYUm3QKBjVDV0jULUb4DelKlEqYMJRnRfi7T4aZckAMAROCGzXX
VIjY4EeYp6Rz6RyICrMFK4D6vCGi25cnyB9lrCgZxNBpCFvxWr42TH+43Lls
AzYfnxFOilw1CBj6xLmqNnFPKCu/4yw+MxdAT0CsR5YEOlPM6xVdfGOr5j2X
9gD6BSKDerFrdUAtqYtTDraXO4GxExVLuwICzzOdJl8Lp4N0f3WGZFa+5Y5V
4Uh12V18513aSqLwEBCR9Z7/5jnbmEXxlrlkfyDLp1banlNHN2sswAs6rLN2
eLbQ0+75sWO8u0++5dGcuLI2qPkUzzHF3tcxik6z95yfikaklTRCz/Hl3k/k
qwhJZHJzHNSUFXn1jhhM1pcsB0rsLCUQMnRD0R/kyIFyPI23078dDutwUJFm
WfTGtgS4qGDwYSQBak53eH73e5kprBQu0fh3TryEAGLWpMFMStkTQ5riqkFT
L8pkUhGOqAVUfB6x9o9olk8nwJMqSBDXOhgQkXMyNN06O9BNx2dfWz0BC5R2
0smstckcmfrq3HUk96/CtWg8q6Ugk/e8SJOC4v0A6amkQPeR3HcMNE0hoJYj
tmKiA7k0VdxvuaCLrgRvReaPNUxauMs7SHPn0rGj7h2ATBTMff5dIG5cTAQ1
SP1xpoqrx4cp4x6qy90RAi+Iy+ZI7lo7aJ4ER10wNk4W/edJ2EgNjISOmiXt
/ekGQfZybKzvTCuCX7RnCOFAMmwwFM+nRBMYidSf1/MKmQpxmf+c7lqOy6mR
HoBEiQM9F7vq1fW/oQUmsyWWo9K4rE7I3J3o8HxX4nl/JWvZLPCDoMnvd+xj
iGpOTbqQIjrz2eL11LU/1xBPErpE7Kj6nO/zvdSdjzonk48z//q4kk6z4ZSL
Gek+8HlFlCIGTtQDKS4JW0LP2VIkHzgEghaa6KnAeW38L52T4XLyKgPUu51v
q+PpuAvGiP+/SjjSf+NEd/dC74oZW0s0QNs7WlVCldp3rDE5uV87MAJxPDlr
LZ+4EH5FHuStrYidxkv55iiJqkWouevmvICKsmjF6TVssJyCa/oTMR6V9DNN
E+Cmf/kUtaASiuw2t7lCNY3zhDIrH+h1YjIWuSmQnFXTT6fRviZUtZcjvk7T
naCnjVy3xl5wR8euUUozIebU2ka9jtdw5BXHUD8JZOUt2OTSkyRJaZrxGWFm
b0yT2FaVAog/2BOeCkYMySYMJCjSRG3120kN7nmsG5prLevBGDmt1dVKqzRA
ak+r4zPOf70hkMAWtBoxx6n4GRL0f8dIIq0VmIUnoveIAwJEIXIWTWdQX23p
wxxsCYfRmJ8BtZIpeRA4l5QPlkVqadVhI6efvQ3UhHOnemfIP9851vgLiEhv
ZUe+As2danbyFkfPQJGl7h1qcxT4kPPTpbnmJixT8II75M4qHu0XGmggEj/X
yiK63UCM2wX/hq6llDFkSou8b1C1NXbRJ/XFqB4JEO7PNNi4cwqFYAAIJaPt
zSeBU4vEQY7oSyBLnB8MAg4ic/lVQllJ4tuC9lDlQuSn9erGWVpxdXJ1cWoC
7gyASzanlK7gEHbTM8CNWxrud3gPqQ5iMHnm/Kt6FN5mR3oBLQGwULH6ROZG
IbqD1PbuBWJO1g014bJHzaBXZIV8HvFAo6WGCtZa29wuorCQ2QE+PPFO9F5b
p1zHCa2pCU+YewRGe6e3Xv2Pcss8+uoUMemJUMeY0EmPEdB2T+mubzwgTOQL
VoE+0hF7qiUZnOGmfvCXiTmEJKThbsNCgEQKVKz89ZCKURTlxudjn41whdQu
5SKu2AsBlv9gyIExNVeF6gJsddE8caDK5Mz+Y7f56wcXo0PSy0q6ontnt8uJ
2YhQzpwE01yLzhknjSqxSrqLciFtEFfXYdnci3r7yvGN2kwlHoHqjJJEyOaq
dI0N+V2+AX765o/nfZ4/AZdvq8buyHImmnNyHBeW/hmF2xjTVxmLQ4+H7sId
PPgU+92v28nE86RUuzBF0IAsLKdoVPpvgm3HX/YlheoeGQSrDiqU0ARqMYwX
YZbck/oNMoXA9vXrQr3hoZ2hxgoHsEWBzj0HA8eNCuNMuTGz5oIdbOgNKNgn
u6P5t0uw+pRCXLqz677Cru0x2USTZJv0ubFuxA3yZIGuhO3/ZaIwi3LZO05l
l2XFgG8p+o8ZKyPTjV6l1ExhnsNnDiidyH41madRmMuIXuA3G6TnIeR0YlHO
4Jh9gtrjFpleDa7hED6JqI+8Mz12XEYpsieI5LMxY9/c7GDkI6X/WJz7L2u6
VXSp5v1kLiWvFQKyjwxXwwmk416+JZduc1rRFIoE8NikuuTjpo9JQlgSoDJa
EXPKRykmV1mORULBksoiGGYjJgSUwy+VfdPqeXjb/Jqc/wcEg86yrklZsnX5
Oy3yQZ/cJ7C7nflgrDX742VZnbHTIfdvx+yL3xj+Gzqvs5QFGw8tAB293V+i
i5jZYfefVMXO4YpkMU6NYCjMX6k6izf4eiRA/V20x/lfK2AlMrvbMJxX4IDj
8IkFqE4/x5Zyp5+2YI9+O+B/KdyIAtGlxGf8naQUDgNhssy1Ma6ASTcnG5S9
LIWxsZ4SF7+1Kun3JjXM04MnT3+4Jhc5G43Tek211xuDtWhsh4oVejnADvle
vru0L7njTWg+S3rsSTchRbeNcwCPIMKJTqueHlbJTziMbKx3sBlFnfKIXukg
IRc6olNIkOv2DcSiVE6agcRKbJ0KtKvRHuUqCHaVGuOLdP+ueLJezJ01JVcx
TBWHDmQSYueDKOuV2hA0khElAH9OzpI2fQrIroJ+JCucLs3ZGihzELhZwkb5
MWlTLHxOEzOsRy3suk537Yy32cGEI4+vY/WzI9cxQleB6DDb0wHaaklrvI1v
gsQe1063t+RlZI+lgfAt38DukGG5b18OhO12c7bxfurd/vRe1qRfXIX3PndF
PfZIESJEY/+e5iqoCoajR1/cgBOfWSmysbAsfCIht+9Z8UNnYG9QHXbV6JXe
6MYSLDpP08hDKBnrUfmqPkAoRAQcyERx9mjIiMXxJZe1IldvdhGLGh6ITL53
iOoT2hhpggeb8V7gRzPN9FGoKYGarFAdQiMBt6fXnCoRct36bZ/M0lBkZa9t
m4rpBdip8QaYBjUQGpTleVHVugenewIfgynkka8yMtKDMJH6ULU5xj663Tw8
MuNKOoiIuidrTjiYF//HtvnpLbR24NmgUJNfm7q1yRrm1vXvXBqTq7/Qk30s
nLzUcg9EuZ++uZfpgPSB5QZE1fumJiTBQVaYbM22KI4k2XqKAJUlXVuwzmUO
cq7dHe7qNtnGCJvT2JlI12QAopV31yovglq/uy/rJnMcZfmTR+gM4scUWXgi
ydIG83XHliwaofE3U2fh7u+xyIz0iPpPh1ZLCb1iU5tHraLCJD5BL1hUZIZw
3Ut64G9GKY0odDjJF7TCX0t9bm9KtrkZ20UsaBMEAFsKrqmTnsCVETYpZ9gL
6vnNu2cH0015tK4o186Yj1bGY4aJJR7GdhNiUSDy/yexGXv24tEKBj/Q+7LL
fCVZZheJiF1+SCOVXkASEQka27N4ndBT4NG0v42rFryy5nMSgXekX02BpQHY
o/5vMv/m7Oy5TLF1R+DeizVDmQO3lrCMEAPz1pMq0l4vK0Ve2V1Mc1GooYTA
GHECyxUK2hLyJaCkSqf/ww2y9VjOFuafCOcE8iC1ernVj/N5Uhef3MzOG8Wg
sC1hPOdWEL5j4Nk+0v9VHZQQ6h1nMbUcAURsfsRGPxnhrSlCpenfa+QN5r4Q
o0MqPTvyBap6ZjxE5l8h8f4CLtmwVT6CULkC/RCfyEa5pXtHrQ/PV6tHouUR
wY6CI43IjafT5PC5VKTUMjgeCMdQMhdIAiLRnN8Lv6PNInyCB5sOUNdkIu5v
oItB1eJucjAGbxXDEi98WpLyIkPzJg8zML8Y1bocQvgeYxGVAgz2/4AtuQoK
aICrsGZYaEL3d1peIFRduWgN+7BqMrqwNIDxWHk/j7GgIzKx4tKx+2cJkU4u
XIxe9iGqpbNsRm8+X/bOoPj/WzgSZfcmFVe6oNNwLMHoUroCNBeY9H7GJZPB
RTL7mhAyvxbXtUJEdOTbDo45InJsdCiLf3ZnSkQB/nJeWvW6jvDICuz1Vn73
obRmRwvdONakkQHzLxb8SImQr4HXxYnGTnH80wKxrY3vX5JiLjhDSmVe2erI
EbzEsf55GoHRljLsNnxpQ5WYUWw86R9IRwFORTA82AMgZdiqbnyvl2d1D6Bv
0zbFiH9+em+2xdo1N12/EtrcL+NNEMRR0mFyWvbVhUqgWxuElmFOswLOaTdw
bjVZgEm9A6T4aU93iLo3zT5JBY994yZGszTLT7V3dSj8uWSps/796PBEgI59
9Yt9meUZfrmOTorR89cL0bMzG1FJ1zUSGc9WGhXk7B4t+jL7vIVF3PdUftyv
1Nc1wFm5ffvtb85oU/XQWyK9wIDJQ8GYMakj69DNCd9IIXQCYqYUZhy1HdsB
Kz85XCDk4KKFOGlrnVQux129rqM/Lhh5Fzb63Wf9+aFLNPkx9D3deYGiBVzq
LPU2wCqSKGk3RBLkARpTOmOfcePAWN3rZrcnAJlgFociSOplxFKixjdkx7Fh
Xz6eLZ+ofXCXqqhiUJvJtDg5Za2a7PXKLggwO1D0laFFI+Kcas04ZkqPOuHb
9e1800SKDbEffnUzbdhmqS/tXnHNqcymg9eGrrINpu6rhJilrV+VYP0iF5Py
WcMTb0Egg2zI0RCw0ncDb0nqyZH9HuQ6+/YZqQIgRPe3mnAclIVdrXt2z8XG
sQ5pQ5o1Rsa7YGsFCWe48r5pQAavwols3ToKVMN1GPD7s+j4Gfn2Co9dd42c
QJFBIu3bLOcII3wFvNde6GqlxrIcsQMLlowbcxxstdbntvSEdpid3Cyaijx2
RfcOmpahMLeGMXpqH3hxyEsiTS64pLMQHQ8kYCAb6UgLECvowBfkpf/FfJV7
XgCYGv4a1E9YIQ8SdfmY7lS+55W3m3BM4lMugOpqcZX+tlzMXMvFq7gn33mm
tNwv4ufe2JFZXc1jQnd15fVqHOW/B/gs6PDLOu8y6yplzm1bbFyOCl8oZl2W
UKvvjUb1RnChPhNT9aBZa9ftJTwkcGB2XlKRgU89XqOY6bWa3Nhw61QMOB2Y
5WMmL5N7bODkmUjCtOdjMg3LBWuLuwNLb8AJm4OwESIscVahVOPJSOPHj4+8
tyjTQ5kmmZ+7aMvaFvr2zLw5KaiZkdyX/ymvakzlyYK9UAQIV34hx3EL7xWE
MTu2cNB4L11bPzvbuNKm4WCVle4caJo3dA7UGQBqMD1nRpJqJ1g7Y6HsfQLR
2MKw1dCo8YmmdqG9NjDMBTohVETFxotI45g8jM5/a8lKp/llBpEJhRtFz07H
xAdpCTobwFil8v4Em0S0Jvgf0MtvH+let8MNB8Jr/Um8AOhk6HpVkZVmkDOj
OkIXrRzvWcpIulaTbO4QOYcQGLbuyzYo91ktOZZrGJ7bd1KAh4/xS1Yoiari
W2gMjkOSSAINiRD/TfjHpXu2yFx8Vsa+15F9qK5MQW3u8pfUbTgaPG8z+ALO
oGiZcA49nwOvpnRu+O16hqWDPAWHN+efeBOJYn6BHIc3qPf9rmTfOTgM9lPi
cEPKf7nvGwN4v9WNol+PxCclpYn/MxeApGWdOuitfATAbVA4LmCvRbgnuSj6
q5cc9zAE9as/PjtC4RAy4rkF+mX29UCIpBMgKBC8tXouSlrDDlscfJhuAqbw
/FMuCuwUIO90aiDra638aVpco1shmKHNkUq0OpuYsW1NeOs4pGK2M8Smw1PH
mcmSr9TGovplXyWTO55xrnGzr4m9X53s+InziYsHmyD02ZzPJ4nzXDY1TWo4
/+lomuMjIfplxh2GW+yLtxlM3M9N5KOfSAZfQnyo9f3d2xDAolUk20L+0jhy
7YHy6DY7x4eq9e5smvzmSM4hPchs0zZ6cCnEPGPy1IhwkVTSlrJTtkld5oXL
P7h1sIdJLQTpwn8mbmN6hZe1LzDABiUT4pS6MjPqaPhj5bhbqnUVbXtXjAuS
petgGZ4VJGNRXt2/zr56VEEsrSat5TWLBTh8+i7xdULkEZsnJ2Hq5Ev5/NVy
V4WFie6W2Y6JzoDBGoz1e844iYU4RiLFSpg+vJa1lXvboUTv4QJy0nYkdX4Q
+6lx0apQTMKRRUcm6e0j3AYhRbU1Pqz049gg5sFFXcgmm+6+GRtvBohKTsE5
uiGGlcIQH2fNYlWc2qkTmX315nrHtPzknuBflJWXxF03eUwe93XeOUp96cXY
7ZCiNg5PVVsKkVCdo2EpEe3akilY15YzH/kU0BzUgvybQg9m5UkV7BVHdMRi
tp8JOzQlNwE2CoOeaAfviAKXg5kp9ssHQP3IduUrrn16wo5rZkkV3gh6wTLK
kBM=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+ErslhdvWiWRkw7GU7ZdD34u00/jgJwDsTRVO575No3GS9wyZip5Ine/Wd/JIjDhghL9zo+m2+sWWKAmEWbeYeFmtALFPE7J6fB/g7xKzoWyUJkmtpBCO7b5uENo0zaMsxU1M6uyOYkKW63zCOHRNRRlmB/3+ANI4HPjfKHk/n3zvlbdX/x0HKpHjxAIMU6/qKif1e49gPR5D6xN/2dyahc/0RFzF8fKgTZ7tZOxYoY6/9trRF+xhlFpR7wxTPF+V9XAGJjBsYyL7rwBcp9axtj4VbmU1UxSVlP6mBG3cC7zqBDNkI8i3yDnvp34RNPi3goeIFmAhd4IRzEBvKe2EUqx+Cw2vhTcgy2lSW966VT62/88eW6+Bg4X9f/Sdpmy8yVDbqxTIRHWsN6fuffISWl6GELxgVfTxgBcEavIYyDKaosdKBjIMGwnsjNu2NcC5Np9ph7iWasb4XShi08/idVhKNczNz5JMJuld5t2H+eGYuSGu/ZIYQ+jEBxq5rA3j6D1zr8IIGxRurcKCA3+86NiIzd/yW6JmTSU3i/wcLivV2sMkIO24aPP/Iy+nbAwXO8paF2CVyZBxi98Fs391DfJ5WkshdD/WidhGpdTnxj5FP0pN3v9QYHTuQBsubp8iioJsH5xen6JS5OaOBV0AaHM70SD6ikNS0Pi8giGqEHc2OtMkur76+FM6TyczEgWmTNYO+ZEfsNHgQZSE2cE7u7Az5wnkDjHR6AKCNY8e4U2mcnk8PDlCqTTErH1VEACOrrSRRzgkdVSo+JZE62eBGBp"
`endif