// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
xCdUy1o0uLgP+j9DC8BE8b+CkG12YtRSTzMmzWu9CSV2JpsFUhuZU2A3Wgo3
39P+4gPQi5jfTG7mcs73B9v82ktjFzswu7XlU4IdWR/+nvoLNUZ6KOVHLpOo
tqy2p4t0B91mEnWNrt4DbzGJlQp80fsCq5apyb0QxoPryyjmJpPSY+fbg182
ydKV8AbeeomiHdboorJv0OC2T1oKJJh4ohKQNopQf2raAnYV8p3jbfzJDiGb
nw2mnNmh3u8LeM1uc/297Q0XNMoiZjJvn9v1/TzdnCxDTMs13BbX0aX2QTnO
hozIPsZZr4riohfwMusNFvH1NV6RnhNq6e4KQVVH1A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZtpAyQ7QYQOwHGuj7PWoCqPQMwHGDJfw70QzZFxpy+fVPoYIn3XZKu1QdqlV
uvSAvEn/KEbVBy71fSpT9/tAu9c+WmGO4kzAzNv2XhcF3yOFQuJWXFDQNZlP
dRpLVhCfBaeASL7wZ2uzm1c5SfDVEDr/sd6F5qJORE7E7cE51M1ld20PUQ9U
XWx+jkvWzUheVujfQ3zOLOxBdWFBpv5aWfo92bhO15MLaChABL0PZtSRMhli
hdUyupY1uEghHYF/8eF1WvQW/M/DGcYGmhPN9FPtiiGWK1t+WX4LNpuR3bud
BN2005rmT/yjJmnaAt9G5NPYpke0zgqAxJLHmPRf9w==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gmSz+3lcfBmM2VOjVd9SmdBA97AZYjRwcbGCHFKRT+qzq03chYK5aO19jOD2
alosE5Uj/B7F1NlK0JWWNeJWwPSNCSJcGzvuljiPcW9sGL2UH8mt4u+1V4jN
58s9iRdHGg5xVt1oxHHOjxC2U5AYDKiW725w0Qgg80HbO/RHIlTsArzKiP1o
t1bivaESQMjs62eUo6ivRh8fqHTJv8rnIlZhglt6N/Fk8lxc+cf5ZJ3ZasUL
zbXbRuJnwUuBxLbjWkN4GNJmMuPYlseZfqy/izNPzCxM54kwR7KYSgp8csge
0RakSH/ul0v1c51Rp/+3Sd72WtcFxJx7LNp+TeUXXg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DyQAYf7/z2EjPFjYP0yIx4tZZ/aXyzT5fmfGeVz2ecj/KxcdXjoxp8LjxywI
lQ9I8bWGVio1Ps80V6+abKQ6mcta/VGkdEfxjGZL0zr4R2/+glRRn94aQdO5
IhDa4ChUMJ4mZZV/yGkReUYTwsuQipDbvxJEJgi1bkyxCshrrdtR4fFpEDQ/
dcnptkacyqXoWmoghFB9eKp/X2E4C+R4C9JJE+5G/JbxFdyEk52DWvu57QQq
K6cVWotC1/aou1G0POLYU4nRpfumOmgHp/mqLs4jZh2ZyvyctfsFCpRRyKxp
j8nLyGqaSOrp4cFXk70cpTmIie4aXpLxtBRq84NfeA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YYgRRJ0AorF8Mml7EJ9VDtlQpdheohhdeldJ1ORyJn2QwzNfdDXweTx5NC/j
0DwQKR51Z0BgkA+upJLzuhnuxdkuwOiSblpxvRdKbzvASsnmTSJBlfaBYmA6
VFozTmHBcnb51+IGIl7szubPzS4jwOMPZodvNw3JYxqrAnHwyPw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
P7LNZOCGAIxvDQII2BmXhkruyJYvV3TwAvZcRsXiYNPTx1VZRpnaQkRvOrW5
gJFPVN0ScQJmMdb7bjYgEAsY2h3jt+wEYa1Ilf4gGvv8VE68BZTzDbl0O6T+
dGXOeX8kXi41ZzU2msaLp3aZzjhuznZ5+eEx60PGGsVc+bHDlzqpt+cXVJGn
SCZo3p9MLAcH9u43LmTXVoc2LWlUzner2azwNJWVZe21PAKEPP/g+AwC5yl7
rpglxhkeJL7toVMt2VCCZeqNDc6c5ZzxmdLxsvZi5dstp7krDzlcqLPy7mEq
Q/de86vexIfMP6pNQruuoLNvcqm1tHQj5r8DfOj/Vg8+gWeY+SR220KrMi1f
pJSmW29j6VoA4fCbax5EJiE3f4TPZEW/nCPWZA0qSSiq5UPdp4O5gFz9nLOM
vCNILku5s0j1R+nvtDNjkmUyal4uI8ztSau3YioxOcM1fA90pK3tnOOk1/j6
ohfkwTu6C1YffXAk2MYbNZesDZZRhU1j


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RXRhmry/5rVc9Tiqxd18Wby3YOUpWTM4dvYZXmPLotaJRqFr7EvXi48Mnbcm
oZOi0zoU+dkd+Zv7m7iAoQ8Q0eGelZy7/2ckEShOvfYpgbtyQH6H9UbiOAUs
5zp/8wWg2bTLddDxBM+d3YiQRMAl4VWYPJcNFhGn0+0qLiutqOY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fWJcSdpcE72efQyMjkpSNL4DCnMarsNXMWO+lKQPk8UAVynBn4wkj3KGsZer
FpxU/UbmJT5iSBA60qb1+AcAYD+Mp16sQ3KlEgsEbmy4TahVw175dUeKSTQ7
/pfKE7phftdmWgSEZWN6BQ+DwNkeladJ7MPl1chhsc+nzwU4o7I=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1264)
`pragma protect data_block
mOupbVjmD4F2kpcm9jc1UMgsCykvgCaQAApih0yuYXFR6FqGkzoMxAvaQzfH
bVOQPgZzKopC/2mUkM2ETJj6Mfu46SB1orqaMLNOVmTYd+D4jVTCxs216ZAa
FYSNd5CxRwRkGMwLbw2mGV4nfxegQNDoceiYk4lz93wFxvUmz0pZ82zl7O/P
O68DJxU8eGJVD4UW5pyoyDjBq0P00fR6E2rMDQJ3JxP1hTZIsewoxPs8DLAC
xsn3Ts3fadS3nUM8xGHpOG5vo6/LSO9g/WM1vzbROU4xPVB7ySJ5S5uiT34C
VZAOemro+vXljLJBLUiFj3OQDomyeAoh06P5psraxiYwjhi0QoJNKKH04u9S
Q0r1mW6f0u3K3/tShKc5PnlWVvyvpV3Pl+cNyiy80SryvpUEaUGuqzO60A6K
8eZuAQhTnIFRQIcQ2JUeInEv5o2CSaLcwTonMsN/n3PiBqxAFatZn5HLEvuz
JzdMBXr3ozu4BaQDHl43vNa6N8N4PU4bwEX3RY4s6PLJ6VAxtTFDMss9xfz8
WmEfQNLP1t6YXCASeoBe2B+0YpaZBxAPcu8B8qpIJJymYPhYKSb5VwvF9vgn
xNyrIofi5+aRrJp3711rdqdnbIUDspE/PLhPd15Tr9uuK/oqhv1dgQD2MfTR
c8jZ6J0HRe/2Z4B1l0P1lQtks+AH6jra8yB3eO8UwSwDi0PcDmKbP3KvJLUA
nnNi0tAxyHszC0ZMQedDov4+w/6DOoObTlIZ3GUX1Nx70gEgjFImtIJQhQU3
c44EVfKSZzWB7F6NxgOJa+4dk8F+iU23dsqFaxPWSWVH7IUWRUmigGaCpVKd
aVKSnyMLgqAtc8KF/jVbOamDdvsIrBTGFFrjzrRXtwJgAcczhu/vqGyvuMSL
CEnO2EaP0oUDOxrgxQJ0F/139l4M/Sl8D4adgfzrGAgyF2GT17HrLIWbnvNk
Yl9C/atymMh1NyC1YhFDYhyAIyuSw3+73LQti8WQEC/JdYsybZNwtXudwO9K
mP02GjRWVRxM30Jo0X/9yZrUdHx2ch7hxt0TX1uh1ZtD3LAPvDCJh9YUZsxl
7RMXrmRT4rkZKOT02RpDQ4KoUg/LeqBGzHo9R2/AsqCMzQLpyX4NcUZtUiXx
fprFgbjdyMA6vqIf0i65vGrz8v/U9wlrREIpWTqrub/uJe3zjQh3KVNgfOFd
73y8FapYmRfTpzY3brGWyI+P2Q1Rg1PIHd3dSWH1mddgp9sXiaRGZyKIOwhb
hIC3tqivNtOy5Ho+qFMf20WsoI0NjG2UUqsyObvMpvxJewP812cownyygyff
APtD3gjzUTJYBIgy/rrEq9bSBorL+YDaHrrwsYM4KH7CS+KtHijJEo0WkiJr
5VxWBKpG81LqUOIaUiTugiKNn0SXaldDnJAgGhXmyHqepL/wQphn5MbVAEYB
vKqVEkXjGfTe0Ijdr9mWN5mMFuEkdvM1gnj5X2QV5+pNbCkIgbujWQQxDAid
gtyDFuAWEH5wVvrIO65PUXFCfKD2GpaQuTZV9PIQXAvCwsA90eABJK/F4WTE
fLIX43hL+YeuALpKgixP04+aBEAKtu+hzebbe+JFRiCxp3i051ntFL4DMDLy
eb+HRrjxl+mv69vxXK8n6OktzlFPr7O1WnfiaglVwusowQQGCMNnUe8Bqr7x
rWGN4w==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqeTMZ1aghiARZBz5KvJcDQ+FcQRO1VcuBdybECJt3z2hU9I6p5GzWLKuGCqfeGNVXzuModxG1XVa6lLSSi3EGdRuG21+1RN5mkuQyeZHlPXLV4wg7eFz8xASQXIDUSynN9GAEFy5CS6kES45PV88grxzpIrCx912iwi6kgG9KTwzSHKNtuBcXp+4FIofKITmZG6REMiDQMeTLmSKm1qPOuDqM1/nY7QYjWHMpNBN/dvTPftfGuk9b01huNN2BiuGfmcbUrH+wo/IBS+8g1y44sxR0tkicIApKVNC9UPsaLfx3njwSfN2G7hu9g3BYNVcWaavx0utVfMangJ5KK3VrxhE0eatnbahteJFKMVPHyDJtBKaYICdUyaQz2XOVjWIl5gzK2YTVa87lZ4JPn8ML15VsXV4M2D10GamFq4RhyQPQ9qBsWIUckgeNPa5kPInDAhkzcrxczzA5wXcITqCsUhh9Ma3fV4zLFp+JBjfZpcQRwQZm20/wp6gBvhDNQqjTglc8mnPttedxEBHmys7yK5VCaFhBTn7CccwsYof70c8Sp2RoPdJcHuFGGxJsNSyxshfaeUNI8qqfXiQU2WdQFWiE8xAFuuW19nF91nngROq//D2rQaRb1rMsLraenb6vwC6kQNEXQq43hBNO83mT9GoeRlCav+Ck5hP7UQ0UdkFMNg5JOAzGDMFhiq3LTnIkDtv/mK/fFrOEkffE66m7Qq/hvw5AJ1Ewg6i/ifbMoo6MkhIChAQ9xaMZXDqSR5FgfbNEs+7oVMizwVZVGMG08g"
`endif