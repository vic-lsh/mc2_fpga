// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
V9zBBDBDco8+sjsD+K0wDpv//LhnP605fh1wcWPCasx6o+O6lcFw5coKPjbi
1VhoA+AD3J7+rzEkN5/YrzZNzv3EWVAWp3uFNbzop8rQA7gSJ8z7ilawyuIX
vJuyLrbDhQp7N6Gl0c4LulzBmSl+YutAxDZdgl0P5dacMoKtnVppjkQ65/4f
WSjPnz6VxEHqhNVdKUGmGxFRwrA1aSn5Uo6zTYmawonGlb/LKqk1wWoyV7oe
lZgMSH3nOR3jJvTcobt0gWGewqrlHhyqb4LRKWKZ1QUlz1PpMW1NEMoVqey1
hQ2eabShwO5h97fPlDNhWGvyKRxGABWFIbI98CcrXQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
imNs0iTwo+dwWKRkK/NckO2bCMk174KfJd4DxnCLX0NLnWLiFDRI5y11A7Ug
pbceix77U06M/EBiY0f/Rf9zfy87a6HN/pafvy/neCWBIvcadvcKUN3JH2+d
J6JOay4P9D6iZKrPp3IoMKAWbi1MPFG/aNE+BASMEWpn1GdZkH/RNx3dgdmH
FoOkT16wx7vX01up6HrinmjwTagbyXur7n+bId9mu8OnLutSHlNByRZ53nMB
KkASTPRE6iksWxfCh5+pftHHV6Skk2ibKM+bU28v768pPBSqhuKn8pVlCXKP
kHcGme8GvyNImY9dVctGSTs63fiM0dp7JmNiSkPETw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
k0noqnIzXgV7f1HSBwfYeJjHubcm0QDxfIsk3frSPouVCGPriQBX1rn9lqll
lIpJMr+n2sRfofloLmpORcfX3vdaMEZmAQEI9ckM6Dz5DqQfG5hBuKsFX/5L
jCOVmdO857vRWAvqiSG0Pw4LkByFNJHrzcdTvQIa5i9xAcBBRGqpBlTNhkNB
syI1UMHOsJ1IK0UrMFMxH5PvXCO17k0n0TKRFp98+w4lxXKWqWuxHpOR4o5v
2iP9DDex6SwMbPO6D9GHOjU+nfd+g49CyIiOWB1V19B2jMWvQ2jwxYdwl9ql
WG5BDa9SIojt9GKXMJqRcH8NAK7YtS6R8HX5AgTH+Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lMvWkueDXkj4SmBDXhMkMbO6DEswrPN1bv0mFOAqkbQlDaXqncVCiBvJ0N3v
UagoL3MyIotSR4K8p+pSdScJysq7xo4LJ0UHkOp+bkEPOVqcwf1nTQ1hYHbB
EeaZHbEJA6DezyWVbCo5vtwHXep2+HUWCoABN1p0RVXxcWfVxMMst71uE3WP
VJi9htn+VWtVOCvqIwo737OmyM9pfBrwwdnTPGoC45NUWU5Yyh4PmqpOfc7d
7tzInEp/ozWCaFQjNXAt9FdVN0kX9ZOcc3VZMB4q+uZpA7khNiipSEY77ld2
6/t36wu1XtMA3bcMsGnADzCw73wXwasGR46JLVoi6A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jHCrbHTPoII0cqYtCpJe1mMa+XPwbmcT23DuxC1dm0tcHWzewQqLTUqXNIAS
plYmYh6wlwNj9KTPG138H0IVzQsWzWG+TrYKv6vPrcfMbriuD2I9iKz9rPRR
WYhGj9Vw2zayCualXtgtyBGbinyhXFl9ebbFdeRswI4/XFjNyd4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
w/6ho0ynZawrSjs8ATw5Kd1omx440FCxC3U6L4cSnLtuWtkKaePQF9GPGteN
GUemzddP+fO3kIUlotL6jlNuveh7qysDbj3YPh1kq/40VXyaKyLgwcPtWTa5
/Nn8oiViWnbG7sGGyW0VH0hgfarN59QUcS7dKoQXidalZ+niBjfE1DwrEOEv
Xv+zzCHcTARmlgW0Ah9cNQLh4tTnyMOSHHSS+HYmPP50hX/5EvpnqImbdAN2
rqNx74NVJFSXPpUNfsKHcJkuHEpiPN3IilapoV59QHwuyf1jH8capPJdmRv5
RAe8P6nVNqV6Hx/YtSK3HjdBV8/jwOwND/U8MEMN1UhC8XQY8KIUQH1ZoNja
B5p4SgMsCFFv3t9SxtqUQdtwqLbYVXflh1Bna6p6Pv5b7nlFR7WrIulohGTV
nmn3CcVxU4TTGRQu+u4Y8rKL2CUnX6xMg1qSl8BJc00pw4BBbc8sh30lYu2P
9OAiukCTya91tyASf24RD82Q+iuEfRW5


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
L/9p7nO9DWf8fMkYhiOfVbtW9/3SE8Batq9hQDRFc1Qr2lp/DHRW4zvqqW82
/SpaeJo7HKu6LNNz8oWfws8ZXbPlGwGl5Cmw9EIQbcrSsR+OB37XRnzrW47S
hZgX0TtfyxY8laD7vY69PmIQKrzyDuPlboJhrnHFQJbwnElAV3Y=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cHI4AbolYhmIIA/A9iNb38+REjQ3yAXRCHJS4Xy8qrdduKSQg/ys+9uvka0x
X8Cg+K30jsBeRvGhY68TnHVBGqzWSS5rjcdt2NOTPJtQ/Cc8t1rzAi9sxuBH
4ZZPiuaAnuHm9UdK1siDar1fGY+88iCeoQwC592TI81p7lpEUpU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1024)
`pragma protect data_block
W/jVrlD+k4o9p/fY8Coa9CYyLr4jp+AFM9zvrNAoqRlvybrlJqG6v/2sefqM
P4r1WLaaTAeoztRxAsaFx/E7DY7h9tSJrOQCdt0swKyeUFewNDOwXI8jyzFj
SuBLxoPPxLZdK3wUKoaXe8jvAHN+cG0KDFe6guJSTwEHdxYCRxnQAkyoCMZu
ctz+C8OW4wRp7YVd53jM/N2wPpvCwFggiSPST6u0JBAUYJkXELBrJb0mkDoP
lzbhlnFw1KQG6Rpfa8VqIZj4tdrEt4XTkXOZ3UqyqH9OerolfMuN9vlRMfPc
Bir49PYhJw8xIb1QPxBXJZg7zr+9vlyjyJoiw7blqc/bg8/nUQs9/m+4vLdd
OnLIE57Nc/z0j9yIfpXzGHDo2E4VzP92zPhfmLLHfJCncRIlluWVabxcHiFk
s4wLcIQFP8PGkirZNh7vqxvUSH/dHJWuPoKvbv/bFywNhEmHVS8SkNTlvcgQ
TX3yaARnzv9E6WvP7NdDhghYWN7fmjGKfTget/EEAzy772T2LuwPSpnQIN8Q
8FSHiF8T418EiOYcdIzMl/IZqCvOKJK0j7Akee+It/kpSoX6TtzsZTh19VRJ
lcC5mQlHFYdBzvu7Oe7x8pcoKzw2gjLVFQ1TO0CQSF+LFeZrW/wg9U7eoOZv
dWcQvBdLIwvczLTqGuQq4iuT1bjOxr91KX6SS7AJHlv/NLFT04ntpIo0otWa
RXpIanzzQcgbcZJKhISkdK8KS69fqDBgWZx+aBkZRlvbAHxXyOjzuwr3nt9Q
cha3N5CemtP2IXAyFxd2dt8DvFuIwr+MtytmoiG3yAmRzWqOpUR81bloasEh
ac8DKnfvnwBdN/uAUaEZK4lKLahRx+u1nRALFiIgPRu+ZE/Xh5SwsJ+smxbt
n6ZxuscYABJQjS7d24sX5jPYt6v3w8p/LfE97MazRPcP5YCMUB020bACWDh2
i4qXznM7d759kObebAQLKsOUFdThCtVijpSGd3106LD7KRzXm615bH1X2t1z
T9fiPpTI0Vlt3d5MGVbRtQx+3v8vtlVMDWAsBUMIuZ7+KyoMb2NqC3SclKI0
EAlR+zlLRzZXxXEAeeokF0DdgBPz5MkEFJ5Fj/H9gofghLvyW8FHA+Ep2Tak
KzvJZ8A92WL22J1b2bnSIaxdSbMeOZk5OuT0LMaMnVoP0S7dcylDocdB67WC
Kzy6s8uT0mP4Abz3G3oXkkhE5wi/23UznSXuDK3rIYZS2u7Sw6HFb2XkDkO5
QUMg1Jb/RYHSwMGi2FO5OoYRo4ZrMTVuQR1FQQpVgzDZCG8j6/fHBaBus5TH
zCntqYNidA5v/4UxFFolW5gFva7gePDw+ma0fqFo/GJ38A==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqej2g45DvFwCLQsFhf7DEZYamtkqerxl2J3XesgZyKSIhbCRjaQR10Fw/f6RGmr/Q5txpgWpdo0GwgVfkftY1RBmHrPVGdOBmxMEs+rYBJ1/Umo5B5BVTs76qwCRNtdUCZNKfs5dCLsIkGwrX03SAS55IwcDGd1hPfmpll3ssilypMnK3ocP1SZKpp1F9SQQq1fJKVxc1MyY6zLz7i+MlvNwRCbwot+SvzdKad7g0YYz1Y5kI2JexLsgsQYuXcBWhdY9kXLCjjrgAhz9HlrpwCsLuHzJQyJm0uFDQXtuszRRJMUpuTVH4aec0EsNE/DcrN9M7dQOGtxPwT10BgxGUQnR9Ez+SESz+vPipaWOc7dyD2zZ54r+MrhRX1Da/z+qJN0MwmeNEwM85GZzFjWc4oKhIcyW2jtWWl24mxCs2/fV75hsYV/LjDocOEzcwAIoX1D3VHpJPQ17UgG9rlxqSanGe8/WroS4QjC+v3lupXTGFoU2h7k/JKYRju8dKg4VvumRJNGaN2aRYlpmpsGtmkubBIm9HWy4/bw0KEFQGn8UWhe5rm5ZGKv5ReQpVVv+eOd/O/84xFwPsJf6M1AID0K8iD77jX940S2DuHOSenVPiCiiWi1hPWISE2YriOIV1cPLbtfHz9yK8cQ6jd1iNzVzNnEbf5Mqs+lXEi4nLtWXwir4In1TRoOFc2+28H6wXu334Q+ktek/PPmdTtxf7+rlcVmVLzLD38KeMvwXH6iT95JYvXXoqPhcroL+PeE369cuWWSesq27yK7vdn9Sjai"
`endif