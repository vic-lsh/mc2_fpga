// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bTnMAJMCDuHjYS3Wpmp1Agsbnfg+pZF5MGpCWPuH227ASw313gk64gd7XRHm
blNn0NZh1PZtgQyMIq7wfkj9tahMDAYwbm3hqeQaqKNNicXoaS2XUP1RE5QR
1NbykdGR99hE4EJYOBTE+ApA7QkCEit9xitgZ7y84yf+kAbnSZsM8OmQX+SI
bNx1e36qeoxrC3vWpPBUxqjs6v5gQEkes0sM9342KhSpPf1V2sEirTtdnGpG
aB1haJ5b+KAmrfZHW+3+npWz7MgKo9BfVHD1PwSvMI12v1JaEN/Tga8VEb4v
mjDTm+o366BG0NSeWOu35Xz5tp/HH/H/7fN+josuTw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MqB6TZI+lFgc04umzCZhAD4rvjGetlwr0ZRB5dbgaIWU68MFRxUhvQWKX+C7
/BxKAz3+P9WBm3D5Xqt596yvzLM1qwbr7D3e7xhTUQG96h81hR4JXv+RqVgO
9ObRSdCaCMgDHx6o7GfF8V+0EeqjNkh2ZxcdKLV/pCFNSg+KEvZqTWxI4UK9
KOYZLKoqAPLbNfwrNCEmCadcKpChb+wVaX/ss9Ohjjf+uY/Wv4SgVwdROE/H
PQWs5Zc3pXUavsi7z4kXqoOmnDMm4E2PX3eGbVBT7iDJO8leBwp630M+9++n
TSq5HyRHbHdG7fpFqbH45TN+1YSuQctxn617X1zwSQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GNMqez0iA5cya+V2bdx9k4DfTXBCL+sZgyxAMQRu8Eeuz8/mrS+BLjfypgMD
7/fx8TSrswTNyubVnmNssRt9SPuiIN+BtZxgX/CRR7/9GNXHP1j7Kj6huLRR
Nsw6nJi6ila1sz4YJL/++J9Glpc8Lo2QsINoWjVPws87nDpgyRLHedYSezOG
/Mic4+Tm28lkjyTFccqPBvUjkJ04nv9AuY6y6Nc6PnmwkWRzSdKtBGOoXBZ4
GCWFfhO9JVdMf1wT0Sxdg8afPpf6j/jLHPyB92DT4hdeXS/b/oW0S8avp9rI
I+6SpVARL7y2fjweKi0PTDkBrwL8J1t5bXkypPBXIA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FPYVY65U7fvupZDqcxxqbuxIT12Ea3cfE3lo6SNFcWH0fXztidl7qPEIWsJ+
sloF5lH9siyQ4yg8SWgBFVyY0RhtBdkm038nGZ7qQL0/hkzjoCx8OhXfvN9q
xHvX6zOKvF/e0riqiOxGfXnSdlQXgofarTxE+5nAOajpyv61a+6ktYHN945x
z0xTmsqBkHkr21FYLH31c3IMW8tO8hoiMK7cBVGLDc1d24/GgtM2UTZtwjjk
QiGOCcyNrRpmsoOpCytyAeMbq0g2fKtuWj21qDARGAzM21+5I+VzZG4xeT8/
b/KxyjHmuFg7DlijufpU/Oj4oy6UomTYnM6l8T/rXw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fqVijeLlmEwX1b1sPx2CVaDmkP5peovJ/OJILsgcq3oXiRVBd1W/vXVVbqJ4
RI3cxz9GDShDMxG+1faCC7Xum98ozobdIEG+OWH8flq8BP6+lNzXjkNug0s5
yAPbrDMeGwLSluBhiKE6ik3y4dQnkSN4yYHmfiD/7wTuVV1GOIs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
QaJ0Erq0Je18qsKhu76FvIY/JSN7YQPZTDW8s4bY0Rk9jkF0Eu2ZVnKWt7tf
pnzfmvDOQ6cwOSTealCKCZ055eq5p+xTmkh8OrLpoahdv2Glh8xpGTBTfuTS
RoF6F1T/eZpJm+qw5AaZq4lqAEsUQ2tTsLmw7v1FX3wGN4xw6RSVhSV5+6NE
SAdoI/OQpWKKDLgqbIZBOJ3IjKDP4V5Z2vJt6OFYGdiI8hoj+70RujpW9TrU
hJ2up8fPpB+dmTd4lOO4DzOL97epFjtsvrz5VLYTAsiisU4cblcgg3i153WA
9M2dtQagqrQaqbnQZuyevlvGeOF4OPOVLxfIpkLwgf2zBwfRv+M1GglTq7X9
nyjRHwLbDuQT0R6UCTAKmbuqO4D7ar6yYCN15l/8hEYzaDoj9/YdH+bh/0OG
2OVaolksHB5qMnuiFTVsPfYhkFG4p5TBHNLp5liaDufKk1nlFMDnZDuNYE0b
nGcViOoyz0tuVW/EPpdmE0n+MRJr3Bhb


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UR4NyvkaPoEXF4o1ZRZrTq8JPJtCgjNHPcQ774TabEPn32Ufx34TUUwY9K+G
nuZMztCW0+P+8KuhCMr0yNaQoJStyO16h/9IrvcOetZ71xLYlcJB3yS5ZDZd
VcDX4WXS00lUx5jEFLH7aDa14XCVf5BvsEr3n3R0DRvmQGhY53Y=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fWSyaigJC60l4ifg76514qKpcwKOTeUt3jVJLGG2wrr9UmLxtg2WpqhMNfcJ
IoPEc4uscesPnCvOY4l/VDxu4RaLKoF/o6rkDn/NexbCF2fRAWDyEleRPqK0
Np+qbY9NzQJefggs9zSfvq8aKRddhjpmwnpxNcAr4xHTy+Bl+2U=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1392)
`pragma protect data_block
N/OOFFRzKa9hIA/ViEDCk3v5V1Drh4Mxj6JSm3VIPZt3AEV68GH1P+tISXJO
GNyt4Ar7S8pzkYMTWeXQGeTpd0iIKJWutwW2HlpXUWYAYxQAjX+Mm4oGvXSt
GiR5EElF5pTMAR8mBh69avr0+0EJ1z260P8PKYAlUOKHgsOu6UCyGJWisGWr
KySEGOgRwQabDQJEX8oz6wjs0NV3nDdV8QUctNd+QwpJoSl65Dy9tFV5+Rx5
7TlkUk0FMwZ6CzVKYhtRpjfZLY+AD3aapZ33KqbooOLZv8WzXJqKGgm1C12+
mKvKoKeombeKqpcUd4lIhNo25Q+7IDOMMDo0fBk9rXX9zVBh+dC0Gww7KOHR
lg0CR+sFyKDBcAtqLRFceXpop42y8ZYF5MsVVtzleIDx4m85c2EzzSSG51I/
Jqzvk//FiAgb7ezVluHuraHV+Ly7UpuksQB5dF38O1Yc2tZdmnwf0uY/r+hL
cytpslEnvr4yOb2ykeetNaHn4HY9jlfasx5+mjThpg325misY8j7ies4I5M/
RP4JbzKCSZcEtFJUuel92yDF2GL0TTJNFH7RJQ4vaJnzeZv85fJTsfUviOR3
dZt5kHKMHUe4Q4mmGXBr4Lh9EtYgl3XTzwqn58+PNWogDgDXbuFVhoqJWbim
c/tm8Kmb2gUl0M7MFTfizqTbFC4eqaajzwX1dTI2t7KUhWFqgw41jh4NeSzT
eFhCP0Zy5VxDRg2eeczKCjq4Izg43KNm5ZSIEb+iIiY9C8ecspHU4TEfz1TW
uxKS3POD2fz5uB2BFUGrHZEVZYHrQLZ/ct/55HABANWHC1n+DM4b2To9aovc
EZyFM61vWwsqmgtcyQiMsFzaBMYjbkFjWDYC5m7T6o4hIaQ8Lqe89U0GbvLl
CuRBjlbRZAt05ELTTw3o3Dw3xzcpX8yClxcF3Ej6HnMqptqd5/STruuRYJ7/
1cpchtW2Z3zh49ocDfABXwYM+NHlnnLAppP2JeOtmHjMrZfpnG/+IIw/HBUl
sPlDa1iU9Y0+2rhupA6kRtLTmIMAqXa1ImgOYrbtW4Bs6qHvuGaTJRJzIqfd
fY7u9ZdNXIv7kyzXliYsQOi9ThdKh6qieOoG21FlTA0xa17dNTlvzoBRgcq4
z7MZ8zDBSrzSbQIr0LgAZWEX0tJCWym9Fn4v9DYpC+N8Xc+pRm8Uoty7+A13
gOGGOxc6CDG+15dBbgqWSY2FUtPMWAAoZ24bDGOjmj2hdvmpMKNA7VHOLPaK
wQfXlsradBPGmE6znYj0bnLNgKLEFNO+qTVPVT1czCbdY3ulVyAAYmgYGWL7
qGp7dEwQF9rmfGk6QoouxXhuDuKGpePZN8fjul/MORk2Waps7Z67CNn2LAfr
gtLpyYvNeiP5twMQDrETmYWE2T0KJ+FiCYk0DMAOBPKURSQMatfXwWlOF+Fa
Mg33SuN2vBzLegg9ufMEXEMElvfZrm1DqBSx6yYZEg4DAR9lwtuyv6N59/in
B9qqhwoNKs871yedGi0vG18h/HY0Kmixpnp76JKeRweVDavLU5VQakIhO5lx
0o50bycrJZZ3gxdoNiw+fYWM/qSN7QWR6J6qUWXFl2hxFG20WH9gyiZ0ocua
pdTLM49e+2yxSaVE2dJ0qAjsYotnbbzCItytrmDTSELMOjHQ4nYxLSAn8jtF
1JU/EjzDPri7f03Xd27VGYZLdJAJr+gd81hqWEdfwKXNz+rFUGvbBMuhi4By
3smarDzN/t1VRYneU7jwmmVheT4oKQlZDqTOZcyOaxBD9Vpa0MA8pCRZ2wAe
hselXMkQIyF9Z52UDPtyPzi66ug7En3jEDyEbUuU3jvWraXuohyvzFN/

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fidd1oyAhusLLJ6+7Y4fW+UxvqV+8TisWbzB76p8J7jCbedVkgTXiBKrUzNVBIRDckfBwS/gk4qyrpXnk44TsazVN20DO3TdF1x8MmH2pGcTjxrJqgYV/z3UJLaYPiY1WrKUNRPOAuHkyYvfI5GoAsKohhmpB04sGLV6+cGIymx/RXK+eIUgAROf9S5AOXsk1U/Lqv4gR7i2yfj3c/IhJWMX+Ld3X1LJ1lp+Ly9OQox52EJ1DZdPQwcQTptwWMUNsXVBosc16pCsVmYyH6eDMY9HRBP7GVYDSCUPnV5iJkXIi5b7C5pLtSM2c+hXhKRz1kH7UTxWb9LP/AquI0AW0nl1goGyzmV5WXPeSphX8LUq5uoXDRE39H7rfqzKJwswuJIU/QsoEVWJKAod9F9+FVXl6drq+WGC1MRr0zpWIN/7gwF5SPoZikXxaTfcDbYA89fbkEFDiBoh3+kSrdEK6kZhppiA6dFatADYkBkJ3g/xkN54nJLNQRnyuanG6qSVsUEW7p4IcPlu+2Da3FufCFQpSzu1zRdI9Oa1yn5Ok7kq5X0a9sfp97k06i7qOhgtUSWuwoxSGSxmskE/Wj95ekGVSpdmFpGyZfXrQ02O0SwTltKpwWQX44uXZeOnabLTpyvBwwFIAZuHmWGiEHgrDYTyL3+HGP/9mOS9rhf+tD2Eg/FummFBqJlZZNEaT5bT3AkjQxfYAFfw/DuxtcUXIyybqYp2cIiN3GzDZb4gf3a3iL494y/BOEvdyDi0E5cVxxdPd12bhVkP67eqDL50bRk9X7qWzAldrsIIgJJVhI5BQH5DOfyPuHuZjsL7t7Y7ltsTQny2ez+CrHJQ6N2V/NGEOliQnA6DkFExT951KdtzIJPOA2iiuubhFPBGgJ46kxbcWMlqWbC0DwYjRso3cTbWdWyFAUxH4V9yXeLDqboq9k9gEP10t3Ar990mkM4X1Lo+TTR2G+f4dQR6MbeIMgZhmSaNpWF8gUdy3q0mNZTQ33TD5EMhFgn7jpSOb9f/"
`endif