// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZA90eLCLrHyI+0qDqyQ7a+JlAZ8L7xKTVj+4khVd0rCAWywixUDhFy6DJ2G+
oe9pFa+ol6EidRddYeWP/h0fcP34RuJ0zawGMeRhX6eWTuZHXJMe/ufqKjZE
D326Am7DWlNt6dt2WSc/gjfLUjjrlIfa3tHM3nM7BLmTmsQm5BOq6hzqvsJ6
69HF+rJtTWLJ2IhqSRZ6SnJIrsitFEAT+1bP3YtcC3BmkWY2F+vb5e8QVs/V
fRRYxyQjPDnlCCgzwAT3Eqw8MewIyQZ02qLK8qVVjBSTWOTm6EjX9W9PihLX
mf87DhxBthCIbw/0Wtfib8Zjjno652mpZR6LmBaUlw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hti/wXlfIXWVU+aBlbUjg52H6Vhz1+IGgbJS9CZGCd+wvQG2HHO+Vq4qzTGc
APC1iK3Oq0+CkGS6m9MDlH0ve+iLC8RDgZqhqoahWfbMCAJyPGmCpEepVtj7
A0k9avLDxHyNeJiL4A2iQTZi6LdjOZB3ItTKCh0Mdw6zsQ7pPl4XpLQ/8oUR
uwn473DjL4+TkNAvhmH9yWXjeCoE5glEhFdTmPBw7UJGrUuBKDxEHh47NNGq
nhZNM/GgWWiyRZVJc3lomw6KZr3AX1e/Zpzx+Lt5iDFNw6RCfhh4uBcuKdV1
cI+/PLQUOtNIMxWwf06W9WmcYfljmuW/dh+Atfkj0w==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RZdgCr6sc8kbzbDBm39XHVfoPdQLBWv+jx23bRO9VeqdbCppdtwu8yEISL8S
CdUvXKHaGGpXiVTwhYzhgB26FPvAWh7fbLSis0pZf5IZhaHWmFXCk7SxBm8u
aA2ErtoXU9tyxCNgUcB3G2/lY3blzjKv1NsP69ESD2E503WF1j/yWml/Y+wV
g/p5+G0HAdRqTJb545YPco3rXKmUrgzcuxw7z2NNJ/4oggdeuAhKaFRYYPZO
G5LO11we6/uFPhe2FolBQ14M5r+eCYLQFOHOdQqBx2EK+66bWRktYZVGmsnM
W3tOWi2eSCpyP/xCPpP2dcVcvkiaNkH2GMZYCcJBEA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KXBIugAwMQ7iiWLEb4nag6isc6Kbd/MQiA8PZbWBaa+VJKH3p0lGucFz2GbZ
YFa+BZX30hlh3uNgi9jAU0W+xpOaB32HHj2r1R31f7qtOWhmxq+1tXDOBs9X
sK0UBSo7yg573SK/dMEj8s33pmuINMCBrbkGOGc7CP6nTAJ6rZLEieLMFCIw
aXYnUmKuPmJZ19D1thSBV7IN8zcPK+oXfKDXI5lPTzhaWq3ercGJc87tiPPj
dKaJc8lVv0N0L8jRZKaJ1+Jkib7gxh8PlIRNzp0XyHDitOFlwgYdAbHlIiAJ
Cg2EqMewaQSaL2SQbm0fa2QZLhCBbg/kjtALb8gGVA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lHi4xH7XGNO/EPs1qg3u3T9dp6oBjuB5eqG7RwqD6JgkGdRLOi/hnWlmspyR
Amjsn1Ce4Kul2raFIIY16n2BZclWFcZCqoRXVqj268wji82Id5+G7XTF1MR3
y1C5UkGNQksNxnuNhFqm+oxWzbvanMJ8nPEhpM8TAc73reSfidU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
AwZH+sIaFlfQKVLHtgCMgiZyVxQNYkS3YWoJSNUwHaKh+dp2GFi1Mb38KgoE
3JhXeZFhg3RpolF4e39P5RNWPX9jO0BnnavbYbLK1VC56o0egKBjvamx/yNx
2k6tfQythfNyJ83d/gjHkZh5yv66xkgjOwpaqJmvuFQL1PHoY8bO6q4fsdEY
St7yRwhTVF2Y/bY/x0IOoxjlnGTZ9hkZVOwk3aU8Ma+gW7oDEgPEeRrWjqVx
hslpjc7TkRpBLJcfMnNEjmfbuB27U/pSvHU462OsHubhLZ3s+UMfiold5jk5
ruHPaxl0RmOoP0o6TTlMQUpg+Cyfz3Dgs5SxQvMlNwqtem4AFmilhesmXzVM
DmkJKFeUAjft2dRrNYXLiuZr7OpNNiWPl+QHn3RvlNojQsUJpp4tbdpaThYZ
FcBUuU4W1Zw2TtuQEZs9vLCOAZsescRKHSEEtllVSwkL1QOkPlASVSarh+Rw
ru9QkBSyHhn4h9rLdJrzjvfL4zjkakNS


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JNHnWqpIxHcSaonOD71GfPTfw9JCQamkU5o2BmMAwhP9ooC1tXhBxGVaqxt5
+kCSFxKC5Glove1nO4lCK4oGWbgAtgKiWLnrVWCpZKi0B1SiQwYM0Xyn3h4z
aTyuqFlXezSQhIx5fkOuwsyeFIZXmncANxZ3x9qGfoML9riQTmg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ppbZ/KdIyv5ERKnHDVqXxmO0Vny0/ebdQekzM4IL+rMUGqa6VM14HMnHRV1q
NJzyHC83rzfeUryO6vDXy/u7I1nVxea24vCByMRyhREIFkz2d11BxC5IHWc2
z5lt1DhnfE5DfbVhDUUy9FPe6E4QLKmVIggZDO+5VE5HgL+5E7Q=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1376)
`pragma protect data_block
SBbdTahZfsKxMat6ivlbZ6urZehbBcY7t0Pvbu3il0bGlMv7WywnXolzTfsH
CfXNnG0VVhvBtGN7Q8mevIfoQIOyv8VUum+XzmwqtO7VUa8u9nHqnro3l6oP
8wMUqxd6U6vJoP1AAj4VEQLgoO2T1AzMI7ZyToCRu9XyzM0VMwrVN34NoSUq
BR0XQq9gkvq+feUymAEZIpngPtjHgItXkK2HcG8nsobpHErykZsuXPqwjKAo
fSLiHnemMj5W0PVtagkMKk4/4NB3FH1gcj8wOgvvstGPwOSiR3nNG75y/znp
xgEjJEiN4/u8TQMm0msxPMoXyrJ8l2OGWFYm/eua7e+c2QjdkGogcssqfE0o
L70bASUD1TqFvp43jeMTSAR+7pJS0Zpdy4iD9sMzpyUVMBks6ed1kmYn6z6E
7ibJDNLytnCFgCmsxHURsCE/mRsPwACZhYbWPqb5eIWWtpj+FQT8X7/yu9mR
Izgni7dL+me0yug237NpcDdpkZkBd6GwMCTxA/QLUW2AcEY/zrmwmYIr13+D
C5v/MroIuMI0Nh6CBCH0YEtkSLzBakhtj7x4gAwqq9NEke46oq22uD9gL9FI
PfErcTvv2CRmloLdQtIcxf4daL91L4zGMbjzkhLdI/2Wg/qVRiZd1K40hq63
+kRr9HsA8vApusbQWOWU3SouhLxo01QMgUI/Jv/n+gZ993xrtL+aVPX2GuZG
wFecMWSSGJM34C6zHJP53OpF/6SeMXJVcIqvU416Qdtqt9BttjdJEyWbTTb8
6B8+6JCq4emD24h9P9zmhSCeJWwPaEKfxRzwSWn1KDXIY+YRjx+LWb/FR5x0
YibiGOU03Owx2om0/ryTLEpMnOmNA/TbsabL/6m8Nc3AGKPGWsLRRKBNuedD
kgjYVsI5Q5v3dlrki8/gNaxRvbFC29U1ir0DCnMXm3rl8oU4r1U8GDn9yBdw
RtjqhtCZuwR49GOoCX91405oiYLJ+xro4OS4ikHRFOeZpuVOV1lygLXWQjBI
IBzGT/vOs1rUHXVG7hy2zhA8vOlk8VVdx6eMUId0hUgqO3j2M92RFWdRhbPe
g464zbS9+G6U4Yvk8q0lDAsqHIINVMbPul1ykIM9aXaJ7HdUJbmJl+TL5z03
Y/GdVs0OAOEjwqqO3c14Lp3aQCH4fdAr/vvAKFd7a6FbGSCbjy5dxebysxoy
EOM8DjVOSJm0sM5H/8P1/+SXWKJTfij+Ss6Ysr/2vWfLgx+5J557K5qVSXxC
whRV+Jfz/PzjAdDH7KPinHTTIeIuA/RGT/aMrg/odP/iRPItY9iI/m7/NePI
AU1qPA6n51Wdif0J2EKX8ZoWub1bWXntUbARfHxvxWkXgCMQlVkdUtelTVc5
tSUCdYHMQcNqTrBn8lOHKanD6Gl8YS+QYX6B4bK2mo/aDD/SPSknZFKYi+mx
9AEO8cou4LwPDqTku/+IKp0lUPh0A6Bn6DxtdLDMme5YtKGvNolYhPS/6pNw
+FYEDVM8JKKX2Qi8LWrfrzxK780jiqCsHGzizGq3shUoyrrrbUb5z/gnaz19
BXwrdgYUeC4Q8u8WFC/v7SRf22CfCcGlpY9mT06JrgLWwf70slbyMQdlVEwv
tLsU5K1SApKXhGqFCQItwimC2WEQUk0yOgh4MnCvZI6Ef4IOps0xv7b+VWJI
Tm1DjsogvX6U0kiGcPzm99jxi0JPvX5RlByG/zimbKs8zPJUaqG1Kc4u1yqE
Qip1/q5m/GSPGpjmFr7wbKfDR/Q8LSkBQ9osX6Fo1vs6efp4PsEukAScHYPp
OtXci7xY+qItDw1DluTjozz9r8SwyYD3p8M=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqfFetwmo6SCVvp3iQDJ5qBE1MmQ3uhiZY+yz6VrAPoxjTRdXB+MptaR4aRJRATzPlF79uLDce/1miKjjCdh5ykfv8nfLKBfz3bTjyQ5gXgUgHX0CjPtJ7i2BIUhTrTGOXLTaQxOwQtq2Kvrx2JWMYMPfrYNeHFgUQKwHggeZYh9UuohhJf01LyCHU560kcGtQz4ao4QeN+tabA7AhUInZtJL1/GQkjpkodoc/CX+LTkSvgvlNC1h1i14uwJLeqjykAmIRtNJdBkh8dZlnQ7mBcdggBGoDkEAyAtE21/kZy469vRXIl+YcqLPrNvM419cZz0GLmWP7zVXekreb91ZLvG5a2d+KLvz9Cu7GWobAbNjCTgxmqNamI9uiGIofX6iL/Qs9r+NlE6dwEevKtqg/jWWglLbrRN+vmc1+zHRarM489yJdeu3AwN4aqvYaK7UTTU8eTyxlwDjPKxlTjx55kVVO3N4aNvzEvktEvIGyPMTQMm7yGGtgdsJNqIdDxN/9JPYvRlvj8wpAF3ttUVyd5Lhhf/nV58dC9ydHY4+aBgNAIIcNwiMtQjLBIImjLmDq4d1onT/m7P6Til3PB+ai1zfBp0s41JR5WJnaQ8r8U1GXAvaA2JOfCMyNz3pGiuWYFHWPY8s7eoPvWgdAN3Y64Bm3K+Puuy+QNYm10QtV1l1bZT/D5lTEuWxYS2TieyBxWBniE1OUeSnsXx/+Yx8BAaYI5YBujq6UwT5HedDQGsoYEXwp3mEiA2Z+x2Uy4KKxq326BRUcgeZ1nUv4lRelWL"
`endif