// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PXMODEgn/RKTdioat4KIDTOtZucv4mvvPi09quypwP9ceyPgEfABzwv5vrMu
H4BPYCnKqI76kAV2gXn3ChoVV6IuikAO77/1+Ii4JS1BR+xTANiesl3d86Q+
OLKOU68cXuHjyGCPgDcmfjfgKA5um6voyl8CUitCa4HAF7Q0aDGxeaRZeRMG
yMXabbzF+NFk5LFpOT5ShuTJQOod7FUg0chhiuQwpv7MO0wX5Db89y41BzHk
gmMyTfRDv60d9RYLKZTqevsP5ezq9kY2XBd2qcruPx7sb0ihlfqYoiR5h2cu
5lGBbkIw4PMZqHBOJuD+SrkqzQo3FQZVwzUmFziKSw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qjAK7877JFIUTDs4KfG2ucOv121KjVWx+qO8s1OJ7iTc858RCwgcZglXHAYv
RcQOsMgUkdqDB0X+auRmIKTIcfaQxHWbHg9gqgK9NwBZItbpwKX8WL5K1s1a
PCk/5Cm0TO+4Zg3x0w3XIStlWIWR95t7BTfay8WpJNv53CEFr/cfBhejAXS/
8MnoxzfwNWRGP6GpN+ssv619khwE3d/Dqt2QIspykKcN+frWUVZSkOjFAjQT
4qzE4irQO5sIJQDJsZ0bIkxkiWBT4rdPryH8RYIiUhQXfXjBbd15rcsgYzk+
N6ZxcrXrHSw6yAP3mgcsnRnbekwzmNYtXvB748DQ4w==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NpeO588b9hI4hrFtVYB172R1FHOIw9B/IuI+n2S+Z0fvEu2jDN+aB5DAgpmb
T41R2sS3CUS+Lnu7XQ+4xj//qobzkGqLpTQHHtsKKJUNaKCVwH8Bg+lbWZ2R
ZffURdB/tghUKw+yt7ltcSYFUy5iBR7G2vxS+ItGCyip5MSgYM56X097RibV
RqSsiFQYuW1GhuwEKBppx7ZBiMmouVXnrdg+RSb24UojVeqQ7iis8ncOR1+X
OnbMlBI80WiNYMtLwnUOZ9NHo3xwwsduOZkSzSS1yRs9byJgFXzG6nxYALaM
RQXDpy9ZK+25nlLoNs7aOAJGDoRj9dLbpsb5GcVG6Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
li/Plq/Ri28Kd/0FShS8f4zIrw3D5lIjJgAlQ9zNflr21KnkKsv9D5VlRZxj
3Da2rrhcvYuUkps81lVY8SXve41q+HMia4Vh1s0WimIeR3re07UBRDKDKEnK
tS2ZXcoGjJoTME1CgLurBM/2QUHmARYsX87pvs7aeLVgAFtX+efSWAHDLLPU
QWEPB8Qex+cKoFR6cEvVErelScyra8VmORxCWZQ1Qd6Ha+NZVl9t2Dix870h
5CFPNhXS7LokOtREtax1AEWyOqZsSjDN/zhmDkPJlFseIiBNPkswvzkhxkEz
sdOwg5ysVTPd7U+BWBbQrSKA5XLzjeVZVVnZkuK9Ig==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UIAHoJxKVHiWx/fnuxm0qbZN++w4wsa1HutLwL/wRf/9POWJqjC2RUDcfsFF
AW0A6vgFWZVXiDv0CB6ZrtN4N1J+LCcg/FJbT04Xo22wZaWcRwTanRVOAyKg
3yrOoixp4u9kX59kTSfMgDBweWa7uMcsrOBjjmQp7ncgX0qsGiA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
MrxMCucuamh8WGbZBgQkJq//SSgRbZDmgP9NCx9CW004mYk2Ohid5SJfH9Qw
8UoTofsOQ7m0bwlQd7X6IR0bXAd5gC9R+6xDqYfF/YFEHoVcpVJSbb+1C4DP
84fTyXpplYcfPcZbIh9wxYPKW658tVEavppZKRgqLfCcIRBYEanlGo+StpnX
LLPeUUJJ4sgo5kNDPKGrmfEMlxIr1nbFzoHtE/EOnbAV2RsNncA8PoxZ8Did
Sr74U1dR981qj/SWqimnUzc1e6zCHUaA2cbusZZs6SRO9Dx5pzSYa0Mi/0wL
OtEnDCuOxt9qxJozfCOI+CWC3Vvpi9e4C5WIHvmKR+2O4cMCQK3GnhO+1zoI
GGKzMhTzLvTeC7Mk3oBgUaD6dq8tPdHKzyHKHRDWC10TNNGezb4Wg4Sy0Yvy
UyqFZ51FQdyNsgkXByLEY77FPsiDMNKzDSgxn/ETh35+d5rQ3MB1FTz1eQYT
1IQmrF8xdLuPHdYQgjIqcgERNg9VkW+H


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GVIu92g99OtIarw1FD61lOX1wnzD+DcZ1rMyjTBMcvHtyMZ81gMrAGrPCi2p
KuRkXxqPtY8WxHmY8Q4lWTtwTss6eaYZBav4AJbKtC+TKa/ffhD7Tj8/5p61
Pl74r6YVPucBDEWO826HVFve0MOBydEHJHMZm35cboVyrQFjF6o=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qM74EcN1ObJSycUztvn7OIKQGkeQT85s0o155qAHwt3cuUj1jSsmoRS8IiAC
0Udi8GsU3wSrMZlqvw+fMCePERYcPWXuNsdb6U4M8N1M8rsaItwU4BZuLdp2
ziA3y7o/1dCSoAOpck7fOuVXfh5kaPJnyo5vBTV1fJlCb5BHxUU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8496)
`pragma protect data_block
u5rJNEPOi3kfLmvRPuzlymt1/7FxEvFAq3dVJAYNEP35N51jKy9Lj4sY6EsP
VyfIjtX8w93Ib+IX+KbdADKjNxr8ZaFWRpsiuz8Sv2/UNn043ufZR7pUBh8u
x1OpGkS6oLmmoJK6l465Cueis6XMd/VtKdTlrJWGdYGQ9zyTXqLXhC3BNEUb
OAIgzD6atupaEc2TFDmKI5VE8BXqnk9b4dT+sINo4h9cB6V0KPT69GEtxuX/
FyS+TvOOSosMiFPYyyuIM7ZMCkC6J6if4MaVUY4WInX6dOhuZEjvGFE6CPsm
CG6aH4XittprTA4/lIskrSRG+kOoz2/7lVH7nbx/FMymRFIOf9A6aDosS5W/
83tJZypiiAEWsX6nZ7qucyUMSiv19OsgbATGN8CiIiP0sSfQOuITs1Y76ce5
BnVe83+YJdbG9t9O1xCMivK685XbsmFGHKEMSnku+Y6MOn6bCuhc5FQAkaUt
epoWxJTFZigKKxH/HaH8wGwAF9DAbRNNeOb6+j3pzAGWI1M31+dqn/o0CgcF
BFLTubXH7ACz8TnZtX0bIDI+P7ZaI1UN6eBE36QNk+f8ljpFVvB8ELTo7IUh
bVOPRRNCfxOpoR7tnLGSRNbiWwvgNYY9Hl7nhVXWZpJR4jR+d1me+WunFKRo
fv6nItaZDoZtNp1sieK4jSxA/WpZTEhKqvbb+pJwfkHau3uhz8gRNHIEFibm
Annixi5TFqptcGlHYF4B2sPJaI7XLDVgDg/jNDWLwRU5mci3VNhreBZ8S69+
T9jtPvnQYKG5tMZ4kbQR7VsSS04HWXeu14cCmr95wk2Q12ZiOwRRzN+bxsUr
mZ7UMED8aisC1Cjm0T6/YRJ+cS+r3U4kpJa+ueF8kpW74oW0Bfh9CFqR8TGi
vNc2go6jcfduQJGFXSqAgg3mbIA6J/s5VltnmrBflEMEOjDYH4VWIaEAklXN
0ea+7kBMNjs8ghp6M/Rf1WTzkUZffNW5ejux1ig7wluyo4/Gzf3wxGeRoakq
5x6d0YxrWYCD882oTMalCt3n57QUV3rFYUb2r5HaXfaNIVTdjXYGDSRUjRlQ
3LrJlKLY0WqhCviH8f9qJ7I5ldEhE/H2/9LyWUnKohE/2jk/zR9P7UjxmieH
WlCR+ZZJy0IOJcmjzbMfRnzymIQv8vaVlfCuQBxcCrOvAsmyIu8N+cvfeleH
k4KfnnKM/AWf1NBDqiOCAQNusJr5rRkMhdojxU8xby2H557DpVjlp+CRwIiM
YFEivCIj2VRG2EB/GGI6r+YPM+SL7lPRooyCzDuFMjxV+W/9mwF3G6zSxmvZ
WSvuWBFagLFVbNloMk/NhfIPFsNVQwuyQ2OLjTG8ePvoRuh1FPK8/84uIR51
jWG1ggh1zEAtICywzpop2+2WGfilyLvCKdw0IGRRIbuxF6aq9HO6GZgYYzQk
Ba0fZxDLaw4tvrolXpYY4z6emH5/dFjIrRrFxJmJUUwBCfH56ythVd1fzqlV
g+em3RyY+M+rpbj1W6AcEfOvd8xKlKVND4ZuCGdJ5VzuGYmcQy9giqYG5xFd
82/E/x5X0Ub9IDM4Fm6okN3IzWtgfWO2Hz5OGA/dFaMp5fx0WmT/kTAzn/dI
oS9vEtv9LRXyiYufzseGhQHtbSOOTaZjyYIWFf6IMZiU4Qcd9BkjhfLAY4Uo
TvQgZX9zgEKQv4bBCoiiKXSLK4uES3NIdSslOqZOfLukVIgZ6BUOuMl3zY6s
gOVs3P8NmF7TseIoUzrwMTOufVy0KIkHB6D6EbtLqWQkfX/1LLfIdo80dqwP
VMC/6CULD9wSwPOb+TnoXAdHu41JKS2BWfZvbaH6YVdTtDhQdqElw/5VeKue
zRcQY0mM3OawCmaJVBkVqOF9DO4Sr4+5cGMQIXkBeIz20tglFQdd9i88uvls
c+SOBCU67FOpIH+myI332eKlLIx9avRwss+Y7sRSOKcnE/05OcbvCBMds1LY
C879AP8pwF2Hnht1jUAyqftJXoDBUtq3xTXKm9gxqxuQjVt36/yt3NBPvtoN
Bgd1cVmD5MtnyoldWAFiWCQuA8sv1WfXiRpXjiFOs3e5uSGv3/qRJXwxJl+5
rsDYvQJJ5H8fLYDkU+VsrJL02NmK6PnhBcGPD5uj8fNGdkWeuw9h+3lo64gi
WtxT7K0FLz5puHBGwO+xvO1clzNxdn6g994juhOuWyRVjWRQ0Zz+PYgpIBR3
pRYfSPO+NyHSrIzIDH4+Zm7yUZD4zVkDV8sf3xyLWEqNdFUunL0QM3o45aVj
6pS24JPaYfzLXrXSB0UyJwgCg12I3n/RyTuqpFiX/OzzaHUb8a/JoVS/UJ3q
mBl8NbDyk4WORqw9c1vNyNkD2YugPluMns/PnR8xudYjz27ci0DHDsjYHheB
qRHn0F+YaU31i/u/gEcSD4fe5VEetsWyduHGRM33C5KEQOQoeOahijqJTMks
4IiZ0auAgZ/3AoiKLr357PjJCeeZr61X88nWW/LFE1YciL/7mFcFP67UkPi3
ksfnEK0tyy3k3XiyvsgXF2TBph6FZes+Ro35nPX6GjL6DTxEUJJhUz9mXy1M
540bmVahqJA8+/zTAs+YT8YxbgmmObt6Sm3/Hpj3ftpWZ5R3Exs6i+XS3qCq
Vlm7ZjiCBpcApZjDlUbAf6mGekT1pAPeEGnplkhictjW8yj9ne6L0ucndCRk
HYC7pRmxeOqHfH0NSKsjrxlnEjVWqa6ofOSB0vUnjneh0FCfeXVvR9M562Cp
eDldbY+1nzTMQNqyQvjB0pLYy2ef/i/nsaYxO48g6+gzhiSihtRuQzNOpu4b
rw8brW5p9U5n8Zx95NQ+yvLaEb5JGw83ZtWIp1fcmmDazd/CO40nqDT/ZYiu
rwJU7bbfNLhyBhEoahPG3kzQPorh2niGAhQMdxnIajWC1pMrctVtaPka6X5b
/YrfChLbWKMmJt65J/uO6ZfVxjjDGTVGP9KMB4dyjJJVWyht8sXonREfm1gW
6RpE5xenSFzRXQdaIkzTTwkLRZIexllOY5D2924QUKBdi17S1AG20gC489dG
6UQYa9QkKw9d45+pVa7AgN0LYrH5HxqYgZanT+IUiEhVAQDPvoLWTZ0SUqCz
ILQl//5JoaONdD5eKL/YScZJMCzel9HW85XIiX+O/doFWui61+OJnaVOxHoI
iO7zNDD4xxBGBaXQMeBbuCZHjc0x4ofoAI9yYNudyImK/GkedODsQoQLPSvP
M3mcXSPHk6BD6bJ/IkWlV4hMSY6kqunoaDCWhcpiy9fHLYjGdxNLV90nO2ts
8fhPeBMsx29yFKlhY1o6NgeEPQAztwnSjNxbR7flcEl3BKp5Oc7PpI+VP+Me
+j1GNlo8uBl7dMZfCyxDv861nbSXi4VMokNL+v0Hr9hCf9EbL5q97+Gft0Mx
rESfGTBMEKVC594naKE2paKZzWWwACB6w4Q80O99AHnQzvoVy+D6DqpWmdDH
z980IHwE3l2UJ+2HHXsX1uIxq3vSfLYMNjzsvo8UeWNCRLEjAr2YUVycCYe6
ct6H41b99v86k5tAyx+F/gBHNAos3hBVMUK3Rsdt93jgrO4DxWuP3vBUBowg
lx+2N431Vp51aGMY7cMi3knXu0+hvCX/MJmr90bGvGevIAa+E0q0A1GnrfYi
zlYXaEhegvBINCytUauGybYmJmcJmnRR+hGNEPX7HH7S6TVGVcqB+4Snz63R
bqVoJh7dI3hTktgIUQDtIbMT4oCKbJh6jLMOro8FMprpSYsuO/6Pf68Bkqdw
S7VjQUwR8p/apyAgqXtvcqQRgV19q1Lk6EW/hpMCs6Epqs2zpCPsVIdT78td
+0t1qRGNqyxzV5wQVwKzYrzedrVi17lMM4Oej8kxxzv2ZP7wWBOoinIuDxnd
9/j0ShLe5iBWIV6o2wWoJDUALQABFGz2y6pjUMeb05OwXHb1dVExpFwTVvmV
vTnVeUQsoyDpKrcPLH4FiHJfSzbJoof7po0sghtAb40k6tiqra03gAJDEbqW
YxGl//JQQ6Xsf53oCTWN9MXKOiRL2Ows3moBzgBrAoH2MuuZlj8DeE/af9r8
JJYys2CVZC2JuM900lY6Zk6xOvTuHGFy8m7yPtNqTlUy4GZpqEUmXh3fnIjZ
9d7K0KkQqyNUKtKZGyfpa53EfV/2HcPv/+P5zIM53jal5lP/taXhIeMipA+K
lE15mgjAebVHfrsuziReHUMuoxKS0T6tFT1jUSkrbJGKVTd+ap77k6wEnW5D
eLZUx56eCAM2shMeBseQdf1LTMY+fZgtF/Q6CsATthRe1cOKHmleAE89QW8E
FuvVbXUAuMrcBW/Gexjy97bt95x9BMTAilc83YzBbbi0IKLZq0SBcb67ZfLP
ndjUfjwOojopk3Oqpa1JjqIqep21mGXx5pH25+lOSsf1NzE8SxkarWkdvkuc
ZlWvC+fBuFaJZXivEC1Os+/rOq+l2/Dzho9fphEHx2lf54fFwTaLVX7O3aIw
0qdFpFEMD6nIyQ3VpkW6XNSJHGtLbdkUln9L1u+ypVggoY9j47U+4GI/sEcp
dHirN5ZfpOF0HyVblp+p5u3nh+jXZaBRchaJftBPZxl7Q51R3eg9VDe0bUsA
dt/d7KZbStVU5T5Trvy2Du/Zc8WabNuiUR8itstPHUNpWW2lBQc0EFQdR2qY
OkkEGH31/AcyGqA7BhBUlaoTXRIW1CIiusFHh4X1Ced6dQXOBflRV0P3HHCE
4Zm6rYlvhf4uU7ipvN6dOekwnBrI3nQgdX88x+g3p0tm2yZHZvyrRsBqCROx
ZSIvUbzvb7mbSMf8S55BT6ZVZNf3hh8WfbZhJE4dEijHK2vHprefbJg7AltO
p1TVMfk8DFOJLs4PVgp+Ud/1aN/DfLfFCBo1rTtyezGZrM8lZ2Z9oMQGpqNB
FSAAjYljTxX1WKVcv1SU4NHM88p7AZrgq8iHeqguoSDn208qNzTJyHFXh76I
3Y8znMCzZlhZrno1Tb14oqPPoZGoygLEDHAFhFNTrN+0ay6Yf2wxSYaPTnhF
kN+WEfrC88aD0zjPTlkuE6dJ+NUTNn6ha1wjMSPG1c36BfuLqAAjRR7s7qPO
EvreWRzbtH1aI/b6Z3chhUXRxwOLOBQnDafGAGYpJvdDALDoqd3kEIbLuZ42
kuo6O5W5Qj0BjGBxsqc2/Sg5u7ZIBTYTy8F/ZYhqHUfGBfsmReWC6BuDSJUw
qbCnn3dS7M7g1qcgWTmKL0Tff2/9xEpK+Pmr5zhuJ9fHSGd592soDagGBCcq
gwE5yGZYjMuouIoJdMe8z7qe1T6RmTLV1vXi/iaFnEEx86e1M1NppSfAuhEA
7TDiJ0dJpoO/WPbH5hB8xndsmwomVQukt1s7wDM25RTfEpaVRN2Vz8HL3jlG
f8WKz5ObcIekFZvp45OrX4xDSbVG29gtokJNmZz6VpyRzajEAqIwa08g14v6
b8JhcVzTqVDYGVE0RIbC9plKdofwfgQe67VjGI/8VDCcTWOFuwNtbnhf8NE0
PZrLm52aMND+PaZKt+G1p7jimTLKIAhHqPcNYvMuMGFdLRU1prOG8V6e1MD0
Kaovbyn96r8hiXbv/syWsB2F+j8KVjKajjJmBT6rkfhoeKG5YoSLherYEbhH
tjH92tzbXeS3/p8fxBoFHcCYRNjzki99JpzRR1fSYHOBa3e6H65IXsHMlNXW
Rt2KbC0/gJMdIWeYLVCBpu877uy2vpeSUOfPr7EaiLCrfO6VD5C+QXA3fjUL
BUT4YYX0ZxGgmM3uKbz50wWjyMwPViCcN1idQ/jhlqdj2Nsp0wUA8tLRShle
uqcSVslifO5eAl+jC+3ggPYJmw+lsKo8m+fBvmGIpHcr6MievL7b9YbT1ECC
A774IbzWlPkTbRO9le1qPa72uLZUK1YgAeECV2Yrly7+FGbNKFfgfDg1d58F
xi62G/HtphZKjftsmYhgUji73FL4ftgEq0KxDXnjwifx4n2wDdNINRyDa3ax
y9SykONGfBpwrxKNuCkwOsbEAuNK0+H3fy++295Fjb3YTc2RIwCGE10/U+t4
H84HdtQo9QF/xpPdTK8G4Re/c6lPYH3UnELhgj9HeF4SUD+tiTYvKAbfKwmK
v+HpnZxFzWOMhkEq9dkX+nrcuUBtSZ3NbyuDOTdnfIGkCvloir+1AbSPFa35
OaQlunK/LjJOdgPn71ZZDjIe0FDQsO0wYIxuDfAwpFNpt5Vc7hxItnf13BLP
iBQrItS26JX7O8J6mIk8rhcZLZ1EalL4rnoupbpe1YZINRzfnLInyQYR/M8G
HK1XoM6L6cRBIl6Zm2eZHy1REtccS6gK2VcujXep6Dbu2+bE162YYJB9qKNe
vniOH4KqSjEOHM2mg3uU2EYUK1itLDSWSpYxsczQDzjaopf8qXfZsp8nWgpI
moonKZ9PmVMq29yrR2JdVIEKuevUI5imqile0gVp9kVp2nH2JizxBqz183sG
BTxZ+KTqoROLjrAs0GzcaqcOAbUZORLlrvaFXLkOegE7U5+Fo5fQgEXHL0+0
1SpkT54FxhNmGt4DCisPn58rX30e9TmuPB+Qetb+D6pJWhPzYoyw5+r/i2+d
53/InIBRKIdFWERWA80EWYk4i93P6GDeSxoGFgXgPAcsKSXGMISuCWGKUfym
dXmBK7mRZrCv7cDojnUX1IUl4tgddB5ii7+pWs4sppj8cOzL9BYAMa7FvegC
esNpkAAyxHZDDU74nRFqNMMefpwclZYrvd5CZCP5a993YHiAYsEqQMOow0wY
CATlbd7fBOJzqmSP4T9zuD2MiQHkL85XwWTQzdPDFqKjhpYEEmIgQcVIdiXO
gyrD/2SxIMiTj4XZNZroHas0QNoh7c5A3voKi4NAcM9p/YsZMaYEWHgbEpFl
s+7Xk0Xov9Ew4PdUSglDVehLJ4FkS//rygY08F9DVaT6UhrK3YhhI2fy2XmY
eirTfDn1ccBDJ1Y7vt+Hk82ow/eP8I8+fmhNHTX4TXAJrM4WwlnhhvREuj04
MdD7M2d3vbFGtsTNntWUmHkh5cIdjRNKaWvyzRwNfyCq3zBXR9VnrN62Qz/R
C+xcLBjpDvXYi/TOSpvSvoNRAuJXx9xDNMEtwKU/45Q/NCG5pw4G34fbGZeE
BtFn9VSYOWDOIwGQ+Fs+H+UhvQJ+boYE1c5ASOpEyFn59YNH8+iPUolFWRKn
j/Tu+zaoCEt2IXx0G0eph9C6hetg1naAvFOL3uTh4bAidohlT5MUUeo0h0RN
4aPozV/Wypj/BbYR53rJPmCyp6OjHj38kEzZ36UBeFaFU+tqrHfwQ2+HEAz+
GvL26SChnbiua+YR7jycVyFwOPO8yuJTGMQiBis8Ymlxl2nWCLQViYLv2oB5
N9LyxYUW5VRoha+HuTf4B2UKOVR4gnv+qTAdJPAkXtFVSFyM2AmjPxEXSUci
Uy3JdfNEyCBDyFzlQqw4utZS1NfY4m6uFrjVKgshCfpL2XVT/L01Dg1xo2my
SiBmZ1k6tYFF11TEiK2v3eJXFgx8noRBH5hcy+9fq1gHXe/s+RYgCFGAhxVU
jnpilrxTxTl7W8kyCShuByMV9bC1Lz09R5ygXIkIyInVgRwDvvpFtOL4V8Y+
e/dttPefiydXNJgVRYDExMrxsP0xCV7cotIQyYN+8kS2rOpoBCuDO381RiDM
dmPFDQzgoqJY4ToDmw/6B5XQOVT8xPfuRYbbifiM2+Z1sbo4Z2XUVWxEp3zu
NvZ/RbYcFVtUmjCs0pKqcBQgje14hUOrZoMyqv53vvUz6Rk2Hch5sw7bao5T
XUKHUlyY6XGnra0rQZsNys9nJHsGuH2DncV147YIJsFs2uT1bvg/0vGrTbwN
I+YGX5//khlJbu0HnAilhSK1IZHMDmP/LiQeteZ5Hvlrluvmqy1mDmVxTAmj
O0+Bg1qI62D0iqFWv7J0a1d9WQxZwCqkiwTMUtXDDjl/D+zwmuXobP9lVofa
BN2Fw/vIGJL61hwVHMjz9m0mkF48sDr72ORxnz/wpIgxirAu8Of+Y8bs3NDr
n2BbvuypYVjoppy2gHOTp7wFNxnO/DtAhcVcTuUr2/qjfDTGTW9irWtwZFS7
wXZyLGwXUn2V05iwbedDGLRtQrSPC01gDQDxdjwXvPWvevdR5BmV4iyBjNjc
ekuKevKHifnTCWJRPXHjn8gBgG00/zvt6tIdsGp4yLrMsfHMNBAOHmxg4tpH
/iI+WUc+qd0eoQRj6OwkYCwewFKcPgCP4WDTHgjPsn23320FcGNlqwl2jbjm
wt0vagcW0PgtftnK+B6gN75W/vsuFseEhFGOoIax3jkD0vglgAW/8ah4HSke
+SOdvDIgycY/IASXEz0MKbtdaDlTgW9Lm31DM4v+8Uzh8pbMaRxYL/bF9w7E
L5i3mMITT5KJymGz4csQbDYyz5Z4di1sxvlW0JjFFOsZP+63UQt7xz8gJ5CF
VCtoa5IFG+D3Boyx4aiUyXoXBb6XnBgm0s/2QvpU4TuXHST8AQ5IL3NofNe5
zjcpixDNVCqtGEe5HsgYm9OskqDzKism7LbVGWbZMzxhsfE4h5k0uSRf26K7
eThsmf6+3K7gWY0MH0OMeecHOloX+PiOrZgSCzN5RDgP3j8wEaLdeXaA62JT
69sXzstvj1RBfsFME+TgaGz5pUXPF2l3ko550cIldUZLE8eakO6Hxc0jh3d7
ZoxAUMk48nt4Xf1+vzpxYOXzywyKwpFAMAke0vEsnm4Nrkw4/8ioLWUp7j4c
yTKL79ZETrLRMKh9vCn9+ScxB5HHySoiv4l6IsavvlEIcnviQ6oofv664P54
/jJ94s45cUwGG4E9DwluIydTkPcQd5/f3qrKuNLKh53fPf63fGgJbdv68Jtd
gwdVEfvZG9JWXyXsHt/iFlZ7nfdPnXzQuI+p4poQxPvscp0LOmRbfxodhKCq
I1I2yI5SPP19OxNpwNqssirgPkBnss3Co2SiKP7Doke7KhV9wquNzYvVJfWS
UlA9LpPZFJirQkU+s8/Ro9xEqbAub57G1hOzObQz5NZpiziQMC+tZWCZwdEu
9yMxQTdw+/IIJ/0u7HjCGXaqbmBfqXSfOoxfOfIs+HpWz4TepXFdt+VuiRkw
OM2ffPMmqfm0+jmRInGaRshIg3ETLGWHk9HYYXAmmvAWecKPogLpKnaluM3w
FuFO6TS27mGnpJKY0sDyBma8dyJcekEo1m4OcR1IkFzv536RaAN6kkrlfq4U
SYK4/k/LkLElKvT1SdVnNKtomskEhJp5w89pwmECe34LGU9Sv982nJ7KUX05
UyEEFERbBBdt+dfcklDGjbu5fGs4B/w4gxxGKBpbEcDUOfopPgXYMMYAKw8T
8Zg1tCaAUBvBXkSYr0Po5vf1+xZP0P0wXT9rLqrjNI8mSQJ3mJ3o/mL58a6b
6fZGylaaaeyNnq6fj0SPNhBvUXSTjzg9fsKbvP6KwqidNkUN7JJvLg9rDygS
xmoUWGJ2ypUWRGJnI+/oG0eeheGxkiJHnY9PHIuZmQ3F6vvCnaMtbQahKwWC
auh54aZ0kj7mTrbVOmQlPjo6JTfHIbmRFi1CfdxDTtmBrbr4sjpYfHMjZ/t1
81Y/83gFGB4ZXb27MC29gBKn81IRPxLDGhrx+ohqGvmy9Os/bIV+jLRxVLpY
MHo9v/T8MP63ugSbE6Qd/v8odtL0EsN1Vwp1yzZjGc5vYckIhLiozilqrUA7
jYRuAJsSG8Dacqz72pg9aeTZSQcacmHDZT/y6DNhJNTcKCCA+dP8L/ChI17N
Jwm5f/wLea9qqoJGLmBkfLkbD18x8pz9sfgH8hB1H9QcfLS6nev55U3pTEni
If/7x2zPxOMeU3JRrus229qL3TVcfJbzV5Bg/bxzTxZ6PZV9VPNJpcwI6DN5
g9p74ZwTehj6LhN0o8JXw1l0mLc3jcRWhuXrdx1aim+NrWMxgSHBiyBTYeVl
FZPdT27+7amyU35bY0KEyxr7zVtAz/iaADx6Bw11liLiARatwdlxeCLCbtcp
bpuO272v856APwUFOzG5nalIDsmvLJekTQLG+p/Q/Ae78bHclvC4vINcsxfv
51mxZGCHooRC42YQp9uDRD3k3Cz1e2X3yDfnPzhXdM1m62ASuujQtQqMGDQi
7/g2C8+Rf2wmsH3fvLlz1/6uas3wg9gfBqsILuyX80l5FuAVzfArodD8/pcp
BaLSzrJqkG0goU9NIFIfvdguR3eZKf4IZlBs43/oNpnI/89D9URwBvUryaTC
/aWNqguGlT7t1uiwqDlDXu0LuUur2FFPDrD5RwoTyHL+0ydd4MEnyoaMfmG+
LMuOIbZiKRcVfhITHDaZs/1C2JGWZYeLgDiWgyaPYNwVQBU1y4Ixr2DpZkRq
V1UE/8GOV18kaXKa7Z2zEv87cB4YQIsdT7qTBhPRJHUiFG9emf5BccUqxMSv
9nnTSeCr6X+klaFmVhzbbfvUXXieScBx46QZ8ykaZGD8/juVTV9iouJU0W1B
Ibiiq62/7RkpHIax/SM8Gx77Ut/P+hJbzvigiZIizrGZhoDhaSblgzlRDgmq
g3vVaRCR8WOYnqiNTciEMXbrCZgZQLQ+YxJdNavhFP1QOKn/QigYwgh7vvAS
dd4daH5iU+RwXfVh22TG/FRxyKfSTi7QtGj8u7kXITf5e45TNPdCnpJz3XZG
WTG/PNlb7OhwooHQYP2AwSh9eFql8ezgWnywSW9QzUR0PnWAzYDo4CXCtC/o
2JtJEqhs/Tvsqmx5cwyWbJ4LOYGV3sA9EsWuP0rKlL/43AsfETuOkk2g/SvE
JYLvuYsknY4G2Horik9d9i2aRQiDJyI2JqDkWQfmRywqnzcENNEgQBGqhGsZ
tzljLK/v/wJ3uLqUtIypobFpWbjIxbWUrlnjk3bJl/T52DheLpDpuyLWIAxz
T0XTpCxvvIbUbWWUICgu5AA6yL+DlUG5Pn05gPbi43HCn++A7lQ7qIw+kvmY
VhvWH2l6WeKJMaP0dfd5S4GRWotL9rs9TNxysr4qY4KFcvc6wT2iBpiFnxLa
GjVLMGkzLm9lwj68/Ov6qA/RMfw0/mPa5q5xgEaWbEiCYEfQIC2iBWHl7M51
jXtaP0FoGpZQ8gFTNtRIkXTCwNmp8HSd4no8gG0v7N1OcVCxVwu8tPXW+Oa7
GTBbTbT8pF1u3wrvO/KYs2FmkcZ6mHYSaRKVcqJiX7tvyc7z9IdUh4hdqozk
zMcshySkny06Hv0mT67pg+xm5z9myWQGScnHnokPAi0jZH/1mgf4gmo/5cQ1
POkFYhncoE00K0/xtM62qg+GJDegrowOAmB5/OAx2zo3RcWF

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRze5br4HoWmiwNS6F19tGrlLC0tsJjRss61D96aAMRc5quDKbLHOUXYfbjH7V3oexRABQ+HO9UuqvQ6SeXkHp68KdDPrprjEKB532cL3Y6Omd/trJUS2kdgio6TdCndZXf1japZbxF0N7upk744+FY3zl/yyxWY4ebijqCcC43R0GRD/ifvnodldym9IQ7jZ11+KSdXzwfKQSSYzMsdJG9DVMsf+m2KjK9W/EcZK/bmjED1AO3KqLvsnfg0rMlwbf3FjsptRqPvreHlhoe0yjcLHE/BmOuV908jAHRz4Vr3jeLY4dsPsiaBADb2W/KSOOs38PfUk4G9bDy9xoa5ocfXkptgskVHRmH6/mKwvr2hSEbVtZm63x0mnclQiEsK/sTN+V28qIEEj+kYW6oEU3G24sciGiiVOBdN6PTvVYrbR6euZpT5BHVy+c8m8MAkaHCK17IgrZHj+5N3KvEYNGXJwoH3tAWhrJRTspMQrzBuCR67BxaVK7rhSvbV3C09Q3mBtJ+mjIyYN4xY4xLrCdMtqixxksm1dfCQIhVEQCZqJkkZAOq5zKs0iHNWIOpIZK8mLwxSOR5s3EGFE8vtjf5hXKByVdKknWZ3ztz39vrwvsH0LEiAKyRQvmHZom2JolaeVsvbH17ITQltQn1EnmWaQt599XeVtrYe3K+GGuh0Wx/73YUKeqCJuJ+fpYe79PlviihaYlk1Acm/WdNR3seHtDJBXTd+MKT5xd7HIjWg6x8r6W1InlcsuZNCGwlvT3R9SVFfq2MOxGrs4zQDQ5nS3"
`endif