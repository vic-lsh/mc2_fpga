// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
S1j3rOG1tv1IzP52WlqeDLsTOFFv/195P29uJ80QVNQndi0f7VQk0stxxtc1
wRk723lTEOJlnDtDIqPaCDkmfwr4CCbnw06yySCA6y8V+RRWGt/gG6WtE9kp
8OHaLF07sNeiyI23S7e6RfQAJ4ekWwoSd/zDyTvIRni3KMthS2oZnE7pIki/
UYTolnhAI4ndfafa+D7IwI8Ute5opaJNI1WkJbDAPhVs56za9TiMaSbJvzK8
RyaWYm3jpKv8djSbo5LeEDP65Hh60WUZEjYrMytF96lEdTi7et19yN5KikSb
ClL48OZhgbzNrBiImM3r+A+by1ArkpvYY3YRIBxNqQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iyXsYmbYUOYc1s/VpyLGC1+pTfpsDd3t/g54OJ2IxOALOs50rDeZ+QWLOH60
AUBszhIGxVjkyj2Ru54iwwePvfx9TdXIMGvEc+m+w/0LXn5O0LtoFpOo7ZXs
tMPZVv5BsdL64ZcERJHy8JU4+fuD1pLcDwed4yFLejrIiytPKJUK/GsouweU
QI8F0bVClXO/SzrvJ6C83V+FAbFeWUMhuZes36nTCsaakBQTvFBekyCUCJ2c
ZjVFeoNgdYR4MDtbEpnWnqAaKZNFy/URFTsD/JAIWlDKtkG6jYfRXZ0H+1Oz
hoK69hUpEwitlGSTbsTKnZCmkjXNpVHWyU+S69jC4Q==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PKw2a79Lgw8Pqj6K/sUr9R9ZnIWumAdYhdeQov38Dg+9+y2DC0exnamtUOnY
/XxRRIgO9c8eC+aWzUpY7p5Ya03YBCnq3FFlfzxAPLRVSTVbg9faB+zadCOc
zcMMLUG5u6Qo6r77jUhCNO+KWUK4ZTwNvozNBCamYhbxQGZwXKKvT0Y18H6s
SH+NP8jYHVmzl3xEJtU55aDXyksD7drSxk3Vf4zit2CTJ6eiR9tLX9QSoQLh
+JhN2MOU0c1FhvZd4Q7ibR7tABtiBt+hRfEK9gY+b+vQo4MYKQ4nbco1XCjM
UJ2yW7xMQtn4WodOtPvuchllathr8wrhgqGclNJU9A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nj98hDrB1p2wPhxevPv6J0HHHMWVwffL7obcMYqnA9pJaB66VDc1+PH6Jul3
efZoEKak9M3yOWYWerObqnfsWSfL+ct2C31B6aCLte7tFd9xZfuIaMU7MSH+
IuhJOszB3nG/RCOXAcA6qSdO8PlL6uvNyJSIwkJ37u1yrojxy4ZgzghfOl1i
psJC7Sw9bKgz2Py9KGo/5Tft5h3ARS5t0U4BWw1WVD2nDEThdQmTI8USDLWF
dUy2dAycQLUGwD2ZcC0MLjwpBTfJgEVbJS5vQwLwM2ON6gMX3lsarQ4xC/uR
E9qbQBRjPZuLzbZhEJ/tJe91sPHhv5VA0TiDHxdWdw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZSz6OmEemf3LgQS9txrW2nILq89Aepw51ATl7aOfG7UiR+87VS/lp771Oxfb
ywnQGy307Bm3umjXHGpdWsuNrICTItbMunfHud5vD93sXCv+2IsYa1p7nXaT
/k5fbvohmwQE3OjbiGXwc0RyIjDpXb+VUkFF8dbFzjQ3sCuS0xY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
DSxNV2aOL6XOTMP/76w8Hrce9GVWcBK6SfV7u6c55ftSQ545/eUQ5SbybfF0
Hfd+GVbOEJxHafvNbShlkdeh7X+VHNPPYF+0A7rUV8Vo08hMzQ2ei1zYndP+
3fTyZJe4S6/H01O6dpOZYEyk+lE4ePHzOXH6yOUVSRXdc57tREmv0fAdD6/u
xUNqFeELJj6dJleVzaS6ZLU0GnGsyYD+R0OjRRsSHtO1E0mLeML8mUS/B3Oh
nEdyVzoyAx7zBwh2Vk/4nLpzmlcrPBKcmHIYvjcy/jCbJOuYkGc5k8QT7jVU
ZPMoqQKN4dZcOo9k1fSV1z5v506ogHVRMfI9I6b5xs73VQKW4oO1QM5ycsiw
HuJWixs3UDsx9M7UY0HzulIwrJ0N7Sjm5NmLDzm7lT+FTBZnsH9tXJ2lt3kn
ZjrGX3jZWxyHqJ3WGF0czdAYmCy5SXMTu5uiQFLU19HZka0CuP70TKSdDKsp
JeccKe8PnARlGZNGya2APkvQp0qLunAi


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Xm4B70RCkT7CxMpY5QKvjYiN8AMs6OmaR+4Oh/Ft5IR0BAadIO9d8y0zuoXv
r2moapzLxX6UWZ919ff5dSYllrDxHuyX0OCTrK/q+J9xovtl8PcoVoblx9k+
9qY7kQfm/Ekpy7g6mpdzATfBNoR1HpKe5kIYcqolVEU6oVCthKU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sGZLimLVQRJDF4Yqt3n4Pgbr/IohgN+mYUGNl5+gPp3oACczFy9IDNAub1p3
tP/vj8ZFRz9pex2vDtxxbzHXSsm3HBPpA5oPWncwigWx1eVyAOuNphAv+9Tp
JAOYNJtQId/vZJwvlTlCWtYFxWFle7OOesPWf7n08nVRLCu8wTk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 24128)
`pragma protect data_block
xi0wKQD1RZEIrEyUSg0jPgfKhtlyep4Z1HZzcCJLejDzZckOpkgkYna/nGza
0otbPS3UoWv2B/SpsUEaxV44tigDZ7Z0OBJ/vQ+V+43u/EvX0Godk+gLkh+p
EfVzJovEeiK2sOoLPyq2wsXIv9a3UBMzE687/Rp2HAO2JPvABfyToWl2S7Cp
0Yuct13q1ox8FEOe8Rtvk8mWg9l9je0ph1f0WfyXe0UFiunpQh3EP2mayGki
4b50TqX2EYY6/AOgIQukK5j8DhZEuBlC74lLmtEn7z4G8edOZXn2ph1QehBl
FduErvZp4MSZ2X7s28FKe0hAfstntD34CSJyMSMM1cJKyTkrDOD6ZkNDAs9+
f0vBp58QVaIdEZkPpM4ODpxUPhyy3b4t9McMNxqxIfjQIx15CEwGKSsqGNnA
UPGDRnzJuLwkOAsFHDGiDcqAaG0qffb6cFNDXn4WSSZ28yBxjnjAPjUTXAwR
yFOR0Jk0WNoChzFfwI4JZDG0t/NL+u7BuwdXaJdfXDocBX0iUeltObsGdaCN
2EkKoh9cBFqHI3NOz9Sq86szEaCxT5UVUTXx2b8Vhoy7lLFA9MwtJUjbcA3D
O3MJps2hwSbgGs83TbfknSIt2IV9S9WlPgBPPeFyg84uHqCsR/NG7KxfcEVP
kMgsV70mX2O40keuS5LweOTNBpUd0qzyKBhsYnV1NB3udj/fsFrODh0BD6Qs
mSzMeFZyq6KDqJsKXZSEIxA9elI2kJpG+TYI2IowFqRf2db5hqZ6ZkxLkLSf
rEBlP7f7BE+TGhX7F+J971KnsGEmaiETHfUs8amomInexZ9rRdzyBr5NRWo0
PPYNisgHvermXmVmgxRz9Hh+llCsJnc8CDGyICF6vyQramiL0r63jXmLhdQ+
9Q7r9y9lbwwYjQCF/51E7fA2b2R42pNDyYpefeF9U/tQczVyccnQ7Js1ek3J
MfVpyS4j8bC22w7RoqhtGKWYS/xnxYyNQ8hvC9ZxIkUQamWiv4zLixGAXY0D
EDWgoV7RK2TZKgeWEJqkheri1r7/LGc1DGbfXyoBg2NCYOlNpFNZ5oW2IV+x
YO8wM5j1orimPE7C4vXZLiVhMy5QlSL8ihrmxHJzUMATddCGdnxzWsKuAOpx
laCqfgNhyGBNNDB/y0uTi+Smy2qDQ9GHdMq2OVj7tBZmbcbLTqE+tA6VmAK/
CpI/nq7z0YSu0fhLe2Z92Tu5UNlEjK9ckN8x4jX+Vs3U5P6Qtx6yiYBME2yp
8d83XGEgsUxkws4ZDnmgoE4EsCm24A97Dr4biKfqzJc6rhV7D7hKH2ociuYW
/sT4ku7TbN6yB4E0/wF4v6LxeoTel9KYbbQiQagS85s8vqbJMrHbOOXT4+/I
HmHbP+z2vfbQjS2OqupK4BbVecSHZIdLuY/bU/ysvS4EDVT71zNxnk1+6YAC
AIQSddEc56o1nn3RQpHg3nzYO7WA8bIc5J+yXs/sR6ozpJpNIQDNPu5AA/0i
zPrKhfVHv7giL0CrQi1YjWzaxZOEtqJ3c4BZrkAd1hQYapqwqX1LLlOmesIk
NtQZXySA4N9I2XDDQSnsoireKjUe+VpRVXGKd2KA2AVgGyHT6tzhPXGDkWyo
dmESQvyRc1A05610RypC3T3uOT+V+IM1eyrTIIKqc4jWqIkhuI3Mk8qrTEWf
T8wBqR8XBtHRIKWtFo9kGDjE8+1/OyqpvZDXHzloa0+lJ50f5QZUb/vkhPT+
vSDZD5M/mLc5swsAQAM1ri7ToPcMCKNU62bzuUi6XP5wnQk4HJgRd0STo23d
NuZUptDnUt3pGMDMu+xl++u0UIsT2Q4qDxMdiG2STfPVGuoQhDjB7AauQTah
55yEEm2kT/neU9ILoqbCVN6/ASo0uOK/OSE+qXXvgXeuKEdsZUlWZKAxgRzv
LxnUB2TlvrPLXCFQhOccxPlqHAXcYGmfwscfTVnRXREHmmKi2gz0I2UxzSKc
1XXDGDpjI5wMBWSMNbHdi8BjbDEvcKYaaK+qMyDeykC81nZFmn3ZrFzdNaGx
uHnKtA9nJcQXWP2txFivJjBO6TZFxWlB+Yo1HOD+mJSC2A8E8fcZC9qNXbKW
8k15LPh0M/iVC7g75nm6L8A13hSMjMxiaSksEKCRMP9I27YteTeMh425ZWj7
ax4666LcxFQWwtCW/htyvul22s6d0CB6g9GmcSqKjxcCbxhjVq0qEn/hcbCd
yqP1Rbqz4tvDBLNLGugHxyYBErKtVFbin+2BTeb87MVVh50fktqy/PoMJkLz
GegT+jxYsRJRr5F7UrzS64SC5jxHcfYhDlBt40SJIDP+22mMwyUk01lYL+UD
7c9xFf9cSDqspXEh9Qk9gJkaKdQp8Cqdfy4IvshHaCAGAx1qq8lRgpKjHs29
Q72QQGbmyhpsa+7he8QVFXCm9n49plKc9rh58RqTu7LnBDuheJEEjBoFZJxT
OuQsCBlwO1wvvZ6GGmiR7BdD2WVfGtOVZKM9GXj0lzwIFYqWPySvpcBp5pz3
uM11wymrw1UxdRngyTr2hAZVxLbAd49EULRtR1pWFU/zojqKADhqfYO+47Ww
VGFyd8nhUPXHjdzXOTyIGnbw+TouYSpCr3smnb0z2N5EsMLn8orx86U4qdb6
CYAhwkbbCSfVDuk19x6VyJLvLkSd9n9jSsAwdm6id3Jy9P6aZzgaJbgG9eb3
vmM7MkvTPGvUtSe61+ZcLfZhVeY9iEVSoo/PnWVRND+YCUJ43jrEeQIrzHRf
bUDym6BGWZaqpgQo8lvoLn4LZeRrvReB3ZsQAlEo1taPKa5AvvM9U/hzqqRC
/Hd0XGEwudI913otu/TtXA/A2L/1A5aqM0zv3xWF4SVQzTzTatrkF5/8QZCu
qx9dczuena18cCVWRp2BnotRO91Hazb+m1/fa+W4NlzJdiQP8iY7NlcblGna
dsJhTxq7h0AxyvPvPWhd9zPE7UDjjtTkUsBQq0OiL6AYTYlCxq77/g4H5pWW
RDNfT8w1vIjUtALOHVyaybmgAqnYDXl/Gz8omA081rYZbNWFoA7sckw3yb4D
o7Qd7L0NYzvjOkfFlpwFc3y6Rqoj4xSA/jMAONHtCMbRBQPlA4OToHpaM9s+
7aYZvPuRZRoKS8Cklboc2qz1XPjIIFankLhY1F2fd+cPHwuqcrkH0e1kVrt7
FD5puial+3snQIipq4k+/6ZWW1rz69tDL/Sy48X8V6d6Q9sc3Nj3vbtjC95u
pRM8JP576y7zg9POOlh6efcQj/atQo1v3T8YaVtmKyiPlgqn4wM69Ahvy8fj
xYG5DGnqu9GMRdPpNjnaJXGStCdiX5kUmAFuS91yWOsjmx+SoINZ2Kb3QD6Y
4Z1/VqfFLT7xVGriZYYPSSMe42GXF8FzNqOuYt5ySxSWMbLT3D3dSyVguElO
FL1/pxswpjxLE4Im+kHbau2UBnvxA1twmFc6WU8VMKpfpvWOlC6ShdQyI1//
rpbQv5ViZXfmlqeDAqZWEV84+P3hmKkG+1B8b/cM9uhjH5iMuGdw7qwt2lUO
7uFDKB/kiytyyDgH0FPdyekoZ9bhMSX2xy1TEjQhE9GMb1Zzbopy0kfrCke6
261QnbYRczRwZI3h0L9VLyboqZ0qhu63ExiYjFnkxhlGvig1jdQBbvJkSUz+
csiTWS/Z4AQW8bUF0HHct1OPgfbNNv0LgV/TY8MkhsriWIUKnpANhiI19gWW
f8O0mexsKFZJi2OYe8KnXJH0dLoFdSvqkboZdcnqDrFuc7K2MY1Wig/7xFds
qzUJnfujKjnxhApZgUjEiGIuJfhH2+PwmXtuK/NCOKoQY0AF49M8d6pbKarx
6hApFUL9DbKrdctTWEweBDjAyIV/lMAXFgTIM4mP5wBJ2W7f7du+s5Ld1OJy
g2FL+MrMxwk9wBOTeVwhy4A+iYEePA29qE+3MfzP5tTsbs6Z1MWLoEsQj9xi
xFw6ICtP7jzg6Xz5qcwKDS+ptCrH8aPSxvAhG6GcO5XAz9TSMv471sp2UUnT
AqJm9BWGQ6HrHat2Pp/2vwWURmkEgquTw9rKZ6o7M1q/GzGVHntfqoQDy0/9
wyl2LamlrJoJwCuOImKhY+A6E8Bn+8ERpStnu9xKdHOiEdKMOAX7MzWo+WPZ
wM+tcnPq8w5AY6jPL65hN4myfMjN55uIdIQoVMMMg1rfw2lb6pwq2RM5Asfm
fA0iX6MRkzwMGXb+NJlPR6hygztwGIso5wUv54xp5SYBtx3S3DQGRIgI46TM
b56EA32x09tLu2I6xsEya/dNR/h143mtE/SKaVB3tpZs4fkg/sL0/h6tDMj0
UZUSQeL3lJLLxfW2oI0rSbdcubzr7mzxlbUjEho1cJlb4Hb4A/HubGXcc8U7
YYcMhkAd5pAERtj3vybzDPEruGTN4o1zdvGyYdWrLH9yOG4EymTp2CeFVzgo
l6KUxZ4sX2ytqhGfeUpq5eZEckzfbBtzqEm9jEFsGh9NvYQYgs6OH301Xvyp
6NgDxGsqmwd9BTl2pxWh7MlHcpHHnt/M92QLiXwvZk1p224QRQE95e3H7eQe
wtUOawnJwgCfyGtaVtHmH/+VD9I5TQpsJePLwYyiTiDTrh0ew3S+m+CbOmJ4
hrgKy1Btb9GHPz5V2SEJDF22Cq02PmtDVKkGqctc5GYhlNaIVsDk0DdViqs3
Qmkf3rscm2k/v4pfob9aXMELD1rO7bmFGMDRgyKzBdbH6Tk2HnFWcKl28zhF
OPoZL2+8g5oYLmjtl6+ZtlWU6D9NLo7nyaabMGPo3H0PY2cpvVYCMqMen3/d
BcIEKQHNuq1OC4n24bh8I/CyoHkMjJjgzMXDyxrlSRueHWEly0b+u6lGFME9
VPmmh5AYi8cGYWMuJLMUzU2KP+H01GlGju6AHawX6kJ9jqA5YwmVS9s5u3qK
O+pjCRxNkzDTAF1yGg6XRhpRwu+VOmXzJIuTEI40nqM/XCD4py3A0uK1YIk3
CTkMo3Ebx1ORM05pS19V1tH4A/pyLkNJStp6shWGHj/WxgtLxjWRzik4Cc/h
1kAHv7fp24kHEOKf+ImimK9dc5BYpn8QExd/Kqt9wDLshWEig50FfXK6qNcg
bcQGyiOUDM5HHa5leqHuZEZLlgYeAUvfMTKMSFao3SEuIEt7IPpEip0nToR2
ixyN5BreBYg+A96Xb6c8VSGDc5zl2T+9kBnQypF9sJbLdMYv9AcZrqCB/SUU
5n3dOHeN0zm1bC0kw5+mjkftAoI08FxC7Ndvgz59iJx7dXlrBPzccUiXLhrQ
QfTJoRycemSJI3q08Q/FV++81gjF9p5jctq3I0EtDSUPR3UxDMpYn+/wb5UK
qy4RuGTitZ/uRWqMC9eY8Lk2xq3QQkHK1FYAEEF5yGlRZdIkaNSQJdgBNYR/
+cj+D86/dRHqwxAvn9XHbKdjuQZQiNxZ274cl1yG/jBUc+mB9x0EDPhnjPpV
ZknwsNXFfQLtUDejomUiPb1z9BhqijUDeRxl7yU/qEGv2lVz28aCspXCdCK1
ak1uvLOSdNOhgSw9ZNuWE/6T4BvEJ/nbkcKW+lp1yTiUHIHWG3DV7b+LtJoy
6WFtoy0+mBqcQ5909uKdGolnXx6Sc+YBKeESC1sJH2x7lOicBYG/aFLljvqk
UcfY5fxeaLdWmLr6trUoexw7QRquTRASuwxv70ssIdhy6Bs3IWX/GN5vzT8X
r+Watbuz7zi9ZJ6pFAFPxq+I1a/YjlsF6vUXOqgZ/ZykVbHv7h9Liq5cJJbz
EDZD4yN8vS5m4M7RDxemf06ifmMqZTAnuuNbfeclaDfQoW5OUThfaCQfBn/e
RsdMrj/7huEM07bn0KEyTNM9IlLDpG9RSWAMk9ftKvdFDYSHIX/E8teePBIf
fLG7b2CobTI5HJP6Ez+h4LwShKNPyt7E0nnJTI8I+CDLw7YLNXDa+zGvgx9m
zHCBRSsaLqNOZGuVRe1EtuaQ8ABhAz9kqlDcmLHOv1s1L7slKhgptFx6HYMM
hXP8aIw6Zueor3nMytdJzmK1dG9Kv4BnzOYtUcffbGt9M8hqrvwSDI/E5Hij
WQvw1gHnV85UMYLVt8b7qjct0UyzJkvHAslbs8Az6dmNsooF2qA0Cld6OFrY
t2eLRn5bEMRQj8io6T44mPJA1FcK96SG5dekVEgbRVf+jZCDMVKR6NsLNLW7
gEB2XAKg1SYkO0+cMCx7qNyrl3Ik1tAB/7sHleQ9iXKEHPXnPA8TTt+/ztDd
z4ZMlyp9ld9EoMRshclQGyxUqtEXbKAyTx05OcZavd5ewyDSSvEM119mLog3
1o3gDfUkYnB1QCBLukv/7rZM57CMMVLHn/3t5vXWQO+R8Wc/DXlxog5w8SrA
IsoobK4s1VRd2LAhXzT/d13CmoCWDYFZflgSGtTBPmFh6DF/y01RPjkGw4GM
6WwtM8XDO7fZ2afV5msVG7VfEary1K+6VNChmek0jC5MZyOVLAveaXJftmLo
2JtE0tSO6R66qV1Y2TuPiJL8Xwm6UU5ZDAIqZrDi9f1cwA401yDrEltW28MY
4DLlaggiBkZZed0GH5Q8TIWpxairMELuf3Ue2PqLZTBvdvj4ZtOUE/hWr/Q+
4AHKK7OlhkjB8/0kJnwvhyhTr8k/Xp9HmSPVBxzNhLBP7usBoFYIZj5piRty
RBUYD87PYNUzJqNr72BMAoEQkqz68sPq4mX6AddlNMqQhc/btgNOiQYdb40c
s40qiaoGHS1DpQrtzZHRNdNAjkB4WsN0XkcEWEijUVrTVF2FR7TOSTweGyEO
Qeq3F4pglCROMznoeEC2rxQq0oqLptHmvRDXsPEl/f1V2vNubQrQxlagLTns
/4wouTAJX9WpH85np0ruovZg6evFJsgGGBW5D70BKrpob5/Yai2uWGIJ37zS
pLGpr/j1qkYonwsYPYD+pWPGPbx+POjROE72brPJMR8bK9D13aSZazcft/uf
+4n6g27mQERu2qqZo4Zj+H+WG7PKxK5syjXibLKTIzpbQ9pkoP+L7YWYPwTX
vov7cTE8KPMPBR+cvigW9+WUGF+93LBHYTGEPG9lS1wipaUAHMzEHiF4wvud
teSn6sSXJNRaFeZcoACh+JEN+I4a7+mMKn+CC8vylJHA80J8IeQo7s42b4Nv
fptriTopurys9dX0hj700Xk/3uhmfPGb69TA1LD2s9KX/LQ9NBumb1+qfMtm
2aER5S7TPmaN+zXMwzLzRJEvuFEJFKrXJAzcp6jkYm8ZMId9vv38pqKXlLqc
/QtHO8N5ENil+6tDU/IcVFulivAz2XsFVK153vkahzJg4IWws8U8s9PJun1p
9h52EwZak3KxrTsh7LUsViZnAPmLJLtYTKDq5pjbOZB57DO8dbq9kW4a/TsW
gKL+L+/kcKMg6T8hAIk2MEERIdatyLfpY3nOTjj+66zqmZPtjnTQwMIb6IV4
9dkjTHrKJoaCRHUcFONztDcv4Kc7JK+Q7cJHrthXERW600EzklveBl6hGmZe
yEkwwGJcEbTMmsSG9AIyWY/TfspgZ5sy8m4b8lXARWseAynMEjAenlaxFaRf
RfGBjKN0DIDfH9VRaKdSDb4v21F4cGKFpQ1zKcwvQqdDqm6POfFZvlWbEX9b
LPFfWNnipNiImOMaMwKJW9H5ltIZzA5ivgbBqFGDDcYaeNqu9718qxuuAqHi
FX1Gozc5KmHcCp54hOHEQGDBvcrlOpZ6EFefh+4DJqcdh0raDGXZvX3Cvzsq
Qp7xLzf7wuW3HWMHAXo4Ms7Z6dijeHxFwfQ22zgPypoMAczbtTWiJmIUEov8
eJ9pLecVLi8WJuYFgpqvXbDasiiKmCornbeWI1W8/o/5qqy7uwXn0Z5wfcnz
YnmSZzfQBNFiEBJBbHrB/qS9csUXeAQA3mRIKHCJst7e8dhmNBxOF9aTRAQv
Los3BbvWF/rUlDqmL1FZh5AqStOEObXAzt3XgmJQs8Js+GeGJon9LFp6ExzN
i31hA4b23F3rgTildG173YU7lyMeKTGt60JMbc2OyZphXooKNdilRVgVOL5q
C0dbWs53qV8l/8D+rUG0ngAo3eIM9vwYW3l4aEzTUjkEpIFcWVlFj1qqtlfD
tRSyp07mdmOtzaGwC/+EKTqliKX2hF+Uh1UqA7/s1GD5PQfLlKS0JuAw8Glr
oaR6ojOqVNV87ulGSimT4VjyqEVB5RSZTnwS39CNOrRAs6iA7J/z+XBaY1HM
401wnqz3lAjK1qAao2s1nL/wX1EcKz58zOH8Ez6VINilsVeo8BqTZuRiUX8h
OqImvtNhF0qRfuP6CY8c6RUEFz5C68kG2k+VFvhUm077Y2fvnf5e5MmLkuEl
Z3iuAFz4cfIIGN+KbVfC8YB/TGyVep30OIZxLdD3ugEfpJfsnG92Vbtzm/Jg
K1txeuH//xZ6mH9DyjYFtmpfAr9eZbxv8JvUc+A7dYEBEVyp3EdVal1Q+STk
ElgE3opPGTYJ2waztoOQ5ime4Zl0oYgggjk95e7XRkJATYwYMOr2QSlTETka
1upvvPxGhzsFK4sDO5ZLpEam5iNz+v1FNrub278x7XkfETF7QslacZZYzZNx
VP0pF3HIPu9J2UfqSa+yynzj72AgZgJHacAq3QqTqURLs2DQXS7XRcAMMf1d
736rhuXyn91BEJbQp8Hm0beIEVYKtZBgpqvGEM9R5jVgx6u5iMcDxPoMyN5s
TVQuhoqKQo5qHGskkBBzvaDdURqDuvzo+VC7uoFUuI31pNFHTrIAOH5+2Q6F
nNzMX2uSYMHUQ82pO714iNRSKxkXeYq56z/kgBgF3bao5gK5gn/inofBMeNr
MSYRpOurI7XY/JdJy7PcjZl2+CAhtjCIbnk8+UlmHd4ipn1ExWXIyWSkBufo
WtmMPedS3CgDGWsYsqEWDUGGUC55MlaH1f2Jq1pw3n0nI1xm1iB4ry87p17j
3u01hSjju7Xk6VfAQeZM1XiYAMX6k1aRaSHPqk0Kjv7iJL538NeLvMn4rF8M
rPuMRGqZQqhJKLjn5wSGrOjSUFGlpGyshDEAGTXrdJ8T9RYd5yPC+P9aBioF
H0Dwf2DCYc8opYKhLPrYwQw9IkyTUWbBEe7xdwBYLCU+YXli77XJm1oSCNyH
BzTZfdtm1eMw+xJOwuaKCf7Wb1LNFjW6CpE2qFS1UIHQN7wOx1e2BaX3/SBl
9i4JHVDf5bbeEjWw3DfvwWw+bW7xPeuNeJIpPQhpKgnIIorcNGQLvzaBO2Yx
AGpMFER/OolgJb/pDAMtowKeJdhuiOyXtbNm6KhhzL5P1UFc5iJ0oi/PKJr8
0iMbDl1svYUE5IXN9846bBf5U8j1ajYHY7b9jFCnL0uDJv8dFKAHg0B+0+DZ
qFDN9A0rceN1yc7zy4yd5SZmViBtccBxFsGp/BbNieHdSDLQR/FYkPidkcCV
PmDEJS6SbM88DmqZOb7g3c/VLKKCVaYaqD4Gfk1p7HRI3Yt6DeoFDQZSDGS9
RVzx4SpzUAGrv+e1SwE8UdASj1lxRf8cHY96FF5mvO97YfqKhg2xCAzE0/9j
XSslkJsMgV/9prj5nNb6yR878yNM33LyaKrZBp/D2Gd6PF2TVn96VQ4KluZI
qYTq3/cZtSXEm5porUbBHm33giXMHGcSPELFQTl2yzG7QNNXb8/1pTqs+nHT
nDnT/qNOgmzFuuQUbrsDBRP+Tt2P+7u/pon+lk5ipk4W5PeS4rAQ6QRPdq+M
StNrqIXGBOoFBnLvmOsSqoph5yz3jeP3vqRXBum3CmO/Y5gfKeVtH+JkMwf7
vWfD/Zh7MHRxCRGYFUrtIF9/aOfDGRYq38g084ikGgyckoiAs5kzoFC+luxW
SwrYcWvfrmYdzuHZeM3v1yPQFdK0aTU4YzAxLDNVose4KLaXWbtDJWKGNY8H
iUqiBm3F9OLq/nV9qgrTjfZG5gEihUQAshuQ7rFBBEHAshCwwbV0tMQJY1QN
S/khAtlZrbSxQ+IWXEWT8rA7k2oBRvTrDGnbJST6nDJPctcs6m673JxC+H4/
s2geB8cJfNEvO+BfrMn9WLAe9iGT1NnjXmknvxmil+22X5i/wIPPWzCDtJyu
nkoW5Xrbra3xsO+hfmY8xUVE+xoOAgdd6PverlDWEMLDKGfi9Qp0yES+EBHk
RTfplDEwl9v0phbD+0RIKZ7U1dr9mRKPTnIWSn1jGPccjD57wAigjL5hzUTS
FLWH29pj7hwi/GmNKVdiWHA6MQijOm0rWWe/SvpyeDLjF7kin4iMOLkACDAE
ng3bU39F3BuRTqhYjZ2HrgSy8btL5aB4DxkFGo5TKBU7ycgb3sb53AOGVbUB
Du1daWsU0PLXPmItunjGflkb3ZLimsr0hki5liYOmzBhc4LY9wz7OXGinEvE
koywNVyEZgj5NbzdXlOvD/D6obkZ1H4YxDM0bg+F75FihwW6S81Li3n/xuSq
NAl7WpEpx0QsCGLD6LwENhlEUBdzj7mW1WYxIOia08MvaOK+RXmDV/sJtSeG
+FLd3+78mDqzxAh8c8V9AEaclupPfV+JFBkVhk7IR/Pw1FGBXKGF76JBd6Nu
stfN51IKi/kVeFspLBwFIMruxcyCNvM15xJOES9xiNbTrGXIYU7OkIn4qOMF
QFBZLbUySm4qnQ8uLy+7F1qoARtZOAn4mQBYpNjZSMr8QaxcEm4pgieAb+5+
NnodHAnRB/gHNZMCfgmA8saR8lij5NymutJJAOJO0XSO1zBrUAcyUe6YBLl6
fn3rRKcniP9rmFGD73pIYIWFyOl4MNRBgsEuQl6xrlxt6VLp/v89UkaNp0wP
ttjRe68tZsETIscCp5D+iW+QJEyPAG6cU53CEwHbioN3wN5DnGCd1e8ycOa3
hVRzBUzwO3reiNop4b3e/4mSsUVGHfhiykgLVIuo4sFYr/3Qk53ANjzmaAC7
Wa9zHDGonm4iow72F4swVw8BGfQcOCLnzi/LPuYA5U9No/2tgfmPmpkB6XWe
f3q8MRDELdhZTD03mgJzTh/jK2SfkpBecFl2VzeVV9yGSwo5Z62zq5MSWhEI
vdxy/B0ufOMDm1Dn5GQYD/K+X5t2aOb7Auf/i9DnvC8UeTVNG/raZ9Hb2sJI
0t6jfS4/4DUH4Wln+zNh8xuES9mM9RLrtTi2eA9EhxaRmjLrhicDTIfksqkK
GwjJttcjjoC9w+zijtAKnFW1jZwZVlQLhfQLdnkYn/PPrcSiNU/IS/p0deHO
dfn3qlUv1I+C7J9JTHPCdo5GaN1YTxcZt1/JoxeS/Ixd7FKZ17fnD+4SCwXh
oOZq5Riulld3QZTtg8Wpgww8gIe+8/Bj3dw0uyxoc6mnq6V1QjLq9SLQ3HyU
9ADC8oBYWL6anquS+6Vnay7DZGMB+UY55dXJcwkLiP3Iv+3dzWT9v1fE1py+
24BxTYehrs2QN62pXz0sC6jewlCLwohMjSkX0VV52vjID6nNEtEHmPPnsztx
J7eVbUX7RzHtBr699HEJYG9t+C/Ig/Q10jmu1BpgcWnHiz0BjQrL33UQWljU
m5SNHQaUi9CbThm7vC8DH5yKpq14BMI6E7eXTzVoJbyKb8ZVs1Eo5MdmRrnL
Lr6jCcjktIjSfg8KDfG0AX/C6q91Wio5tkzYKUwX6vYQ23S+UU+SffZxA2wO
Wb9lHy3UcDaFd4XZMkFD2mrpB3FgAa9G4PHF7xCm22/ailmmz93RijpUPUCW
8oiBuiYHe7OBJvXRXWhC5d4yq/zmK31Lvv/akjr8IkwbyGCbEm7FeX9TJaAG
iVsTMg9djmuPIU3loCSkcGuas9lhLu6+dm8q5kCIaeHZvguAIF2eFpq1h4BV
wPkvnp0M+GavW2OiRfPJFT6sA9rUR+LpDpuvH67Fiflaa7EwqxfxCVJvIRHQ
1wr2kt5HUwkJJAKMFOQmfyxsuR4g6eQxRc4BnMKf/a7CClmJRI1KB2aruRyP
vRibPCqDfEFhoU96L7ouKYwV9wW1wbO3vVW4/4NnwploKaIzSv49hkNP4O8K
+I3RrFyFmtl589WMoMtDUE4wyx5pGfCda8wHkWhygWh0i9ixMawhhoRpJqI/
7j43S6iQCNSARpwKBzqW7D3gwK00LQbSafH3oThrhcAM9mXM+HSHP3NbBpa/
bQ3Db4c5tcpqZGP1ZMHDLAvkL4FYHHOv01mzTMajJNiauBesqldrSAGtZuSD
2zS2l4hP923uGlm8MLLnkpkrhMKdJA2Z4X68R79eON8lcQnBCKVsSIl/JbcA
x7OmJaR9epLgvikpFPUXZz/qEV2WUGZUVQq/CgoDJYTQwEAmE/7u9E2bZzFK
+ZSap7NPEaJc3Zs+9T1QnKTflqlvL8SxXhAZJ9e3vAcwLlSf75fMZJon0gDO
iBxpLKrI2a15DaoCWjq7fRjpCHAMjS3xnwgf4Pt6PjHp88t074SODW2Mw1vC
jBAYOFVtDkZkr8qxDcG/J66OCCTd5E7d/W3Uvfij9e4tsGx4aaepPH8q5F9u
YYxaW5MrDoXm9Vifw4PuklgB5zn1YVvR32N7lBC4vtJZhereqET3SBLo760z
fDUqmCxL/Er1WHpY5Ov+IpHvK3X7tQyeVPa3DhP7FVI/UvX1D1CIbnqJly70
9pkQqomsVlEANeP8y6O6bHYhL8eWVnDixs1Lb8xX4Fdmcyy64TSbEbUZBCSV
4laGBPzOF33kWgGx7az0TobQ+cAFDyFHi8Wyhsfn0ArFshu2RGfqONOVC/EN
D3I3HvORDl7zGldURxY2VCfP0XQ8iuSkTwdS1Zz3He/cOL4c7mNTzOUAl9XK
pbHvTml9FZEuaf3swmj9zy7/m3qEU/45ddExdyNHomSnCQyyMyecKJbMG0Wv
XgA0sYVH8rsZsytZ8faYmwJfZrBTwgU5MuxCnGHRroqLDYQDW6py6+8w6hCj
jhVcAcnDqSZ4K6oqPToR7fM0eQgvaAi/frH/jU7cFqIcY5qfp3ZIBQAUFie8
njBRr8ycHmP2oOc5gyd4mt1bkmCaI9DYFn4aGa5RK/qAaZxz5RaOesbt3V25
+AzNj6JDoZg1b6XW69vT0s6cVIov7jnRdU2hhXsC1FCvDjrHoO/+1n39AHyK
o5KadjDm0GFcNgOYRnfpqicbKuUPZooytpnELX2pMfzXDRZzQxkpbANSlwHo
acWKWKw5YwR6xIxiKbLNAqUMpPcCNfIXIARkHf9wD2mfnSLNE3hsNQDjxcmv
XJMhjWdWr5I+dRMKU+PACNyhoDReKLpVEd2C0XUrv9ILAItLe9k/FJ8PlF4T
66Tvramql9bqMmwfuWdYcw7k15srdVxhcA0b6C3qcneTYA6OnqnW9RSQ1/QI
h8FUyXWcvHRdz6BrLu+PmMiGy7Jn6mhqYIqlabs26qzZElD2B/x/xPIK1rV/
0gBbF0MY9M6m31ufOJShb7bnOFdhuoJrb8kuKPsiJV1hKalI0MSksdkl1aaW
iekMyIGUDPveMXyDHi/EgJJ+Pn+F6gNMvg8DfVpifDchcfy8k2/s2U7Gqcor
gNwcus6Syqhw9iO5p5p5zN3Q+QgRCTtNi2QTP5BbtVSDoMcOHI7uL/l09Ss7
BP5YKBjJpMJCqwmaV84TbRionTRNDCv4XUCWmdRl+Di7BdRz3lUXXmJe5dsv
yMY2klAvLw9yhDZTfzQ1TA4oNkoj8NUWjLIbOEp2gJKOx54mhuDRam5ltf9F
DPpiE7DwElf27t3UTMsM7TTRIhJQQxVS9CO5/5tZNX/vIKR0Y8c9JzFpmp/4
qRLqdNp+slzBXfnGhvo/PGyW9TG2hfXvB9jcUGDAERMM1WCafjs+SQWSOMWN
1eCmjI3P9K0odchZ1S3tZDTOEdwief2hazDnR6ztA1EDE+tuvTG/dJwb1dX4
ELJmmWkVXhxT4NFHxykAh23ZvnwTI+1n/u7RbS0rqKZnCHkWNZ2GnVOzuqHC
uCapias/NH1pFSWI41JIzg9n7+xF4BLQuWqRCk77S+Ghocvo+jksUbbFR8o3
Jq3a3l07lj0IpKQRqwwvS/zmU7uE8R3Ju7c7MQCMr8aw+25yXVrpSkKdyAiX
13lE2Nvs74prENSTkCxcDl+gMirtbw2PkVXygrXM5LRBr88HMjGyPeGTyMiC
IGgm4h4wNzuelUWQiorEfao7/m2FDq9Ge86+8CRhz816RFki5NDcL8vHyyGx
zoQY5aN/EawlyMCpC/jNGqSLsIzadzfDc40UMCq0BDtM+pT+HPRb+0HnhFvd
MfBSkYdSKFYz7JZiLBUfpyF0qzDuaWUmqzCJchKJtQXj2a0fFhKy+lSmMX93
H53D6pL6lpP3U1lpT+TUVU4QzQoC3Pp7p882TpVxLzW3jycAXLQ7VhJq6v2f
eZxep1ttpOWKJ5VzZOUkAW1ZJg5/Br6FcDRh2DZpby1LBcI3Tua816Vt2E1T
qqS5qtIOUzrEF6EulSBih4l2qLs9LKkDLHv6B8QP9WOzcRx0aFFWC18bJPJY
CQ4wKs9gZ6Wg8LhtDBPldwoJT2971uhjBmQ0zvYZu/lsb/ADw+ZEt8bSgdCI
DlGUUgPbBpv2Bz6ZH+cxWi5FpuiqVFC2M1epupLoyZB/hijN/02aXg+pgNFj
ANOvRFhKSNMrT6V10hnHdlV2w3S30xvO7U4hPOTh2nvMc1io0B8pgHfYgyBk
f3Yj/ZseQOGr5k/2wuWPWb2YhiiGS3JUJo9r+3jCn97T8MuatlBOkKAHTiZe
FdNX+l82q4Ul9x/Nt+2M3xnrwyb90pj/0minQnOXf2wvVXj+l7XKRFftxZlc
bMe6s1MvAaVjwNi/CrF1c3j1KxccZuQ3MFi8OqH0wApHYt8EojVmP0VAMWvR
uWsdfnVmRPHJiFqLvvJ/Jahi+tWkjslJ1Y5Y9cGiAS8umCclmC43abTXBULP
aUfmtw2XUP2sAC93hB5kTm0IdmTjESV0fpSkngza5ms3w/O/r+hLoB/FLI/5
2nCP2NvRMwhipdnwsa3Ma2yzq0aYcVSkkG0qO+AhwWOAk8HDccgGKlm6677m
Tl6ZhSLnskzZXByy1pDzWrbaFM0wrA+lPiEFZxjXVBz2AxDrNKV1Q9PkQyX7
m1zSshvW/+C8M/Doxe9f/srxGB/OXFygmMRvXblZaoVFKxq10KKzsNTtYG+f
KiZtB6cSbc6VuCm6JLk8OdxS3XKu2M/5VWBzZIcVQ2F5A57BmzrdJ63HxY1A
oUv1cYw1AW4O4vcWMtpE0BhMPcOfOeH3uBoNWvjIXpnzhtDta46Mlf3NOJgm
1KFQGiZTEF5VPESy1UtMxfVUOepB3EFBvsj9zVQ8kdgHbK8XlTAq0b2+ufXy
VOQZXR3K9rk5ydvbm3SyWz2xxJB3Yf7ry0HuB651usNVMvK1lhyntlaUhB0q
eM3LNn4amucYzme0DGVTWQ7qOhqa1sJhKNMubJ+Ip4TJxIfvhVYNv3Np+K4i
JL2YYQG83F0C3Q22M9ui1K06xdlpWCpcEBvGfPWJXMsX3okxGlyOduKosZT2
mcDQyqfXmtfxkpfMNQGamcrgwM99Qn/ynGpVVFx/Fc7D1J8PW5xjGQ6DkmEc
4dWyYsVHAxAkNm4557A9lIkd1DysolV8JoHTc8qRffLwCCtKyet2Aqq+hBcX
UVr5qm0l1HcYxAxh0ZoagYC7mB5uNYXmhoz7NErUqWqlnSJma2Ny5UxXK+57
WSp4aM0zWY0i/Mmc+t+QP8EneORPi92BLZPhg/LQ4dUNpzmCUongsS4DsBVP
bQBpYh8IsbER2kEWZ6od2qDof0lppiVeWrZ7PgLy63vgRCWTNZEVfZBsSeca
36GJZBrSQ0FbXcqqFq2xUgFvJYHNldX35BragUse5IH06IYoZr2koUTPKP62
EmDw/kfMFGpkd8lcKDfhF6/Y3UQ0P3FM3s7fQYIddr7XWku1PgRprpMIRAnl
sVoeDcNUXwdw1P+9GOyT0Zn8iaGZd3U2Ijofe7307GsxdpfcP/XV0JLfAqDW
uiIJ7hs5yxEQIZ1qHIADt4tWZCfPvTURLDTJBx03JQP6FeDCG+vYHxfqPDjm
yczMuco8mBA2BbIv7lOnwvIrQIM8+7qfhmqKutMScZ7sdfCd61vVtJ/UatGe
1ElsjYV1gJouUPEc4RC0G9XKOjoqAJ1gZorxFni5K+yT/sUPMDjyUCmkC2NY
wjurgHIpY0ZhCIa4tA4ezSlB2rtzD/snFIvBg1OtJlwADkxHRhxUOtN5/iCa
D4rK9y2m3DURA6PZPxwynFRAqJUL9LOwpZG0rgR/5mxAENeICkSTUO9t0HCD
l7KqH+HDKTeYvtpqqViUIEMR326oR+j8WYdyM7quHbE7L4592DVn3TBoYOaH
OqzZa+JQjIwaGzKtjsHpgR1/urZDOCUUvCYgCqP5KMnoL+uixj0nUVF3v1uB
3h6G8fdeorcdn8oK2gcgx2hbyqUdCA/L5liKKvEtYB0wEUVHl+d4wU2jvuNz
3tDw1Ig6gShS2K1TM5ImPAAVf3jy6hajhf8ZZ9k+Rkl+jho8HFZHUcY+x5yh
Tppk9lh2wSfsmnquRuSPJWf3LQeIQioaK6Iq/ciMHrb6kyaG/cdrxIfjGEn6
pt/yTR/0sZuQKNSloM7zNak54jez7dkct6C5wxM/+6Xahe12gGC7QQ/g6LtY
1okoOiSv2AyccqMKwvnm7nnEpPDhi59hSKMIPKj+2iFKG43mFieR17T7BEvv
82pBFlmCOT4HEzZQxbdmTsJtN7nvaH7NFohXwnoH46cPDNhEAS/+BRFJm/Wj
CN5Y58qKETrzZPnSBjfKvKSpehuKzywn0IC1wOS2raN6+cyRVAn5fyWbqLyS
lxA/KsUGcSp9J8amha2+pqTVLtUBdqxwE25gkLv/vihtsPEdZN6bOesLr+33
xEsKSL9jKQIk6xUt1VfMux1hef3UhR16/0MrdHwBoCXYgfIVA5b8JUm9Ixhu
wxFdlUUF3/jpxeTTUpiw6l11eiqsxWXajE/Mb2z7mtpC8QCbk5ZZC0Epl6H9
liKT7aq9/KgeqmE/kZkiedu/qZnllExz/J0dLdsm1Hw3Nw3F7YDCDJ9K8Ap5
BefGRyPz81YO93SM7lccSvzgPKQoMnEr0swUx0j/qENJZ/ypaQgCwAY8iNBS
4cZAungW3sQE39ymj2H/tywA4hRXOx8v5ohtP19U9M8dSC5BHi9qNQI/LSxh
nmiAxgOKkjNGm9/gQfm/qk3ElQdg7NnSbe1dc3uT8qIFI5Dv5SQTsfyRjC/W
4mT9/biVIMffatrhsPpTk/iEBsKPCy7p8OijS0mIzMlrq1DGa1iCW5JiNaWN
cGO4vINSoYIp+LBtKBlUizWG7+EsBiO1hvplVgHojwEY+i54cyfH0t2XpiKl
1JgMyzjbEw7qgB2sxiXoGDIROt7GVX7UWcIoz9z0j7kLwVJKal8GmdousmEy
iNtO2PYRUiiGdw1siWWBrHe1kVSUNHIZNffbDZZh2MthPtotjJGF7T4cfNKS
iYh7vCxWfjvXJKIv07JRiadsBhXp8FZOJV1NAqCbF9B/yEokh5wZEzlVUJ/m
kGjLpX8Um4sX0gs4dTwfZU2zDtkU5rQ1uVOgCJCGkJRHxo0V76Lbf/zlwMQG
shBUQqErXaNfo7Heom6XHrj1R4kRAnotZ2hxn/mvuNdjIHrHqehrGCngasb3
mGHihUVMFQ+YTf2bF1D81waz2/WMGXl2ukcloIMKyPMzAklSEFaEBoIyLCj3
BIXAR5CkwBRJ1T+yDlGpC7V1e8OdZpN2W6jtuDrowjX+bISZ34tXvTdKqHyV
Mt5IVv+T4dKjF1RduSHT0YZsF0EX0RBrzxiBUOvttUQabq1Y09EQRurpUxAi
f/E0T4lHrFcwKiNuRYTov1DY0oCnLjUj53UiCp4Ro1qFahwa+sqDPGzPiBJY
GCBeKina8llegvoZigecPdWPLJscKvRHVLu54iMrFVQX1EnQg+Tcbu40kqAP
98gv7iyfpvhY+I08xTWNZqKvB7y8cXdqO97RPCZEG/H5K0GDIn5ftyToeCWW
akRb9nJn/lAinl3KXsvU2OQ3WYuHWMe4q+2oUUlYQin49PLZmO/CCmn5tSUS
/DgbLTk9/0CiBN1xSQPGcfNrp9o9U6HQnVLnay0YMKJc79x+QT/IzCN46ogM
uxXJRxMjFHW4M1hxLGK+Fiot9F0DJvYjHBnwNJ+JBit9lyNLkukxbNVNMglf
+VuRyS5hiNpyhg9z6MFqbY+R3315/1mUjhvTnVSfhAhTVi/cswe39IUcwEyO
w3GQP+QSbWYlDxA1T1lLuZV0YC2ZNMrHVU9gc6qmss7yCFH5AWi+vf+cZLcD
j7wFhiE6NKt9Zz/AfDhLO8iG/gI1QsJB9xEttieO0T95OWPOrA29Ii/vQPX6
37GhShZ6+bQWaaZqCFoZNzAwp/9/KdZma2GBNrd1NcNaYZ/88L9bbRKVSSqd
m5226xzqjcbeB0FMfe5/q1MzIuOF9a4XiWWlwwRbviwLWQec+rUoB+ZWCRA5
fKeNeB/pYukhx0eo8kKy7b757U4wpesmTJ2u91xCCus+pQnaZLKgIK947+hL
mD9arPDpmFfqPsTF38bi61dbbVUOT8EdIjzu8gC19bzlYz8qscax5wfb7y+W
9L3YKKgxWmTVqQw6KozlHTQPHl4o8saz57ArtE1xMd/Ou3OGd/NfDqsUSrjW
sKeLyj0ncOyrrX8vxlzsy0RxZHJ5ZuPNmp40Tm6UJdwbiWe+gItJOv3aOc+y
LSZVCSeZEVdRot7a42qvWcEeCniE3PHdxkJ9IsViBpdGMUPjsBiI3tSsv89b
xiUcKcBv/q9ZZpYVuE2fN/faVWwtgrICzTMkyAotCVBvYVTY9Zqi/y9nowxR
pOcKgB7OVmkoPXvzVs1J9ZQ2GbOhiiYEL3lkzSpEoZKwZXxWoIh9hEYqqZC0
dK4Z1HzqgdhNYb7JOcS6+E4nMFIAcnF9UuSisZ5m5e3LtotggP4RNYDcfNOW
lm3+GILQ00kZjbNbdEx41hwKMhkxU6t7+FFO6/YGocvFfxGUUBC6hApblCyf
mlKJluB7X3jtEqS8aMAfiY7un/bWkX5ZszK+619WtrfSferi32gCO4yV0+Zh
/Z8gB+zwyD6W4Av6mNlkUxX/9oEoIpossLR3PPOr/80vVHj7obIi9NgFwuco
sbYKaqo2rJCI12XnRLzJ5byVPqL93CXtxjLwU6W9q9nEeQZUU4oQkpXM//Xc
Hbx3YF3f1DiS696yWbciQDJ+qIDCwXXtfWe2Xu4/PKfT46O4uzfl7H9CbpxD
Et5b4CHnDHp68jtxvEizdWBOMUrpJwt6xtZXPTfuNatywSWPSLU6qgEicTii
Jez9rfq2m+JGsNKOc0B174jy8gafmBFSFD8CZAKBjohOSzL9GVeBSLLgOvT3
XNscWjKi+eJodF2UU/OJ87EvorxUQwNq9en2iAAayKntDT1Oi771gZEjFmSN
O87CZeomdEKcgsDnRb9RD8lX8DwmdyIAeEV3t60BKJzjMAZ8Ve0FMxhr/EFi
na/1JLyuA3yQTdoH0UOgMXWJm7vqFtXGkLQGT/OZesaTzdV90E5tcT28OOt8
4Va93erObAAZEvaeIUoVmW2n1hlKRY5Xopl22iVrQJ3Bod1t3wxaPvjiHGXz
JvwJ4M3+1KTmHNdAS187d3fRd9e6yW7uMi+PZ7pupaEptYzgc+j8dWE6IUt5
QfVTZTVJOImy7f+hUsF9CyuvXcyMF0wIWlpFhYdc3Qnt9T6He230Pq9ecrrS
fdFLVv9ym2MbMf22yurhXJR2V5r+P4OSNpRcveDiABsmGVrygMLZ5IY9aUw5
+0Y37rdwIyxFiASILFKSRuGlddGJISDxYD7tZycEZktEnaksIFJ3N/empvmr
sS8JQMw3lH5BNkkVV+D+62FM5AhIoBPmelNAsaYh4i+L+mBuWNaCnW3+RMY3
3QwGH0OPOt46uhGEP4Twp/Spj6lXMpuEb8uGVUlGf+VDqyt61Uh8+YVYzqlC
L8MLupWepw3BdytwlYVN7aI1f5Pybp/sc3nnQM5+rK/CZWepkRf7eV+2/5yi
nGPckEtp21gPIbecylgWt4pEjwEV/KZHe16t5NQlwgvzTnbKods2h66ak+bt
jETj7lO7Wl7jwZ3vnn2Y8Dunb547+sw4nVh3IUXnJmT3NyRpzOL1V1mYTM4E
JIshdvyOnoQo3/YYGzQm70hbsP85FdK+YbFuTrFhqD3IU62uW1kc7YFpRZaA
ZEETP+zoe1gdbBT354NZw4uC2TRt5docxGTAbF9teClpw44tX69Ef1MdXOsF
ZmOHGVIrRPyd4HdUa5sVy5DwMl3gDqJGT/1BPQvHXLwQ4AhsasyvDfEMz0vD
Ev76kzY0WS7vpKCK3AaBPQ7NAcfa9WRzozlUuvcgXNfOUsczDsn84t4xeLEC
4gRRNTUoKJD6zykNBbZm5MC0G9yi+Zqk5siWHVgld8n/B2KEBJepkiL73Jvf
sd0qE039/2ltQAHQpCY9MtsuK+J2I4mehDGRY1Op1llhLN0jYcmrfe9J0SbU
7XaSfQyj2QRkxPEkUJAMlwahg68tJ8bNRlhSLDdqRheB9VKlDT0n5hxRaBCN
zbg9trvK6mk31Nsp0e/CiBRWU7CXFf9YKsyp/bY60YUgMmuz1r2KtIYr6mga
7X4Ku9nS5UNdS8XlrmfJSVbAE+IusVay37pgTxMyjf28LQ+uhJlQ5Vfuhrl4
EQocY0lEUb6XBwrGWBUQqeq2ApRG7tbFV8GKB4acTT7n665zGDhdFo0gwvwf
qiMn8/9BG78RW/+w2whYar19rwUZ+YvVUmPorGgPB4ENs9UBzhCs7Whl2qnu
Bi4DzBZKMvsHjLWHfM0CQORh34Ru1pn3L4ksVBLMfK4yJBUizr03eJJehP/O
y3hBYtsJe1ibfp59q+R1l3ubuwDwhow9YhgI9gzYBtmJBJiHTiid/Z0ksLJi
aM2TqE14L0t5EZhMWH2F8Y9fBgKTCCrP+oG03XhEReqtAlo4KP3q6XogmkFc
mjbCrYc6/JcGRtW7hKl6xGeNkZonGDIL//NgsSKyIXEhhVe3ONYz+a8YoWtN
Q0sDP0FjGNVec56Iqc5b6Cw4vPc2ub3YgkUPIDs7iT1Sv5gABB+2b6f2dGD0
5w/n9fufp0heMVs8YojR3m5zbcvhMqIJSSnnyF2LNzhrWUpUsKRdU1Z1y8Pq
Oe55qvnxn1+3yDjg+fDZen3vwVg6DdmSQ31zAkjPp3g6UowKyrGXYFBSlq41
IlExkeQkrN+ZMTLtg3QcPkbCwkonwOXAgNqHZGQ+0RCk6ShJ4cfyk1KRg5Fp
GHLe40iLYWpiQbIeLo+I0XdsCyT/k8NRYvN8k0MQEMoz4qrNjpNjZi9QHa4a
3gUCMpg8kq1V4EDJdYYVHF9i/8AuYTsRA3cQfczSwLvTrUQgrM9zVgnDe2Vw
i/lZX51D/pZWSYDOYt6B2dpaAtFKYPn0Bq/dUioTFCcG+29gQtIieqkXpdYL
MaDYK6wV3gFdRXkJRv5+7h/f/+2oQ/mSUpAx4u8BisSUcV40lP6ryoXfz0Sc
K9JJUsmy/emzEiLhSuKq1KgTZ2wryyeWejlRRsrUDrbt1fkUnWBfaBydFOMj
H962V9SuK/y2ngmpDB6wcKMNkg+ym3VvGW92thFT5x/NTkQM1fQ7a0EuSZTX
ca94Yr5E/Tmaa2fLYjfGaNLMnTxUw1fYKlT7Eb9rFZ7bSbETEQ3hfpinjuLz
BrYs7UuQyirAFj1vlUyAU6SkOPyfLl3Nfz4mrsspdCxtyppvypAXQf63oFEi
EtvOhMZp0cjrJoFDuFJUC7QNBmlyiqjLVaqGqOihqx1r1+oNJMOhuy6BkBM4
4E02YZ9Y5HnOQA2JNsB96oGazPEq9mBgmaYSNAH9zlS4YWq/yWBtH1Sa8/LO
W4Ky3Arb31SljsicUOXH8V3MZAOucBtG8tikZOq2Kbear0pjELnLtjPyeJ+g
sJPg39lW6V1xRGOwmpHzEojjPz1RpI0opzBCeswRIGzu0lvX7/cKgPZ8Xmvm
v10eUFBrii/Y970vC6B4us20Lfdom25RvkBdBNdMKyN4QbTgrDtF9amUKngL
uviVlmYIiQFz2hT/gI0ldKsDZc553NnBa3x7SDSSoouBinatyA4zsRJyeH4g
KWiB55uMw/1Z+Gm0jj+wblM7/o5NeNpHkhV01J6yuQg7qwAoRIYTv8dVDOqN
6+mc5lnQ5Ii+uCNGJuGTy9SoP0i/G0rQl7b6lAcnWBWp0zxTp/V2cNdjR30y
2NcaqxlAk5paXpFz4ijrjCzfF8EHvBivbdL+C0Nb8br7GlfagK+qxqjgNgMp
GjCqNOYXMC09FWrMYAVvag6ik5SwMUWCd0+WxYhuIK2/R8SeNnxFtGZSgKl+
lMNbbiF9v2OZYwBOOq+eiGRX1dc0yY0ApYF+siHWuF/inu+siAAAYG5UYBqq
7lQKtlCbrv+CoyTARx1NPeoj6gNS5FecKDUlZJOdSI9jIChbOOGEMsxebI1r
L6hI6Mtl/fIBsAsYRaeSXlYPk8oO1B5OSJf6jR6khJVLuVy+JByNXh+zAWsW
yv6+mZd9nNB4A2EklydRe9lYAdxpgiiztxNOF0f9MICoWHC1jOT16Ai3x2x7
FQrwUmLvAeRxxCYtO9AHlv5vnVoVtVqIcGaDAoaBpnpFD5PP7+mD/7ip0fZ2
NeMl8eTkVlsz9mbZ7StqMRTLvBTF8tGQqZ+72Ke1/qGU0BdqWnp/fkVsYmlD
905H6zh8jLHEfzboAXDmxDw1b1ZNCTXvs3/lxitD0ojxGBD1W38NTub5BJ3x
KwoRAzAbq94x4swS4YZrCM0ZOF0ZFHfoqILl20s36NoZbZzu8XIjaG3CX6fY
B2SayVCf72hezi95nHlsBrrLiSHI0ht6nHCwHPzTr+U+7hGlFaXCzvSLH9D2
TW0e8mZ90Tmbb+x9VUIqz3OQESsvfshyxJnv6uklpeUkiBI+jEjYDw6FbZ7y
cLmpPzIj2FwYcQ0aoNw6kl7XJkNY+25qced4SoZw8fcw+TvZya9T8DsQhCy8
8M8I3jPkckhtIz2gJpFMCSZU+i0i5s0NAEFRhNpRSPNvA5fKGJEnZFtLkpPi
d+3EbIolih6uEROzjBcO/YZr2sgfq6xUqRIQKk8H13seHBSLK2QvUvUgHTWu
VCFIBIUZTSW4wd+kuggwYkEIFb7PhjlbjSUfvi7vQGqzNyOoXfbDAUdQ6sQw
l6FXrr/3V4+3xx/J/eDtoGzQ2KIrn1fhlJL0haqQRlzygBcKUMuf50v+SYcb
Y1YJXSm7OrqdU++293qjHJ5sufd0qFAM32AkN7RMEplvOUi/U3g2HNWjwI9Y
efTR+uN8ixtnHW2g/l12LUlrEDjH5pRcfHVa6c0cyH7oKTKkcCwM3y0zNseW
bEKFVe8wPTCOpke4FhnSqqPqSwfW9Iut8mOPLrzlz/hGQerulpIGdC+HCK7J
aXErSfsB1u1YQ6+OLje2uFvQ7kzsg6Fz+0hxQsr24FJ46ts1jd1PkteYxWaj
Ikp0wJeKONyBg2h7rSGtFC34XFYRONt8t50F8syH3xTgQr5wYzEZIjLa6o5v
CvrVnh+hBnVgGo9tzgNFELYoHRdRtG/anoOccr9nA/RapY4n4ZOpvG4+orpU
MXjtO2GT7AJbOa37teoA8QPQpoHDDSl63m8pI+DiclUtIhjR+sJiCQ/m1xQP
DMKvQktmbV9WAsOPPMyP+qK3yJ6vU0KQLLasw24V66LTYSNmFB98IMIEqcoi
3DczhBh6dAKul4dNoFKdjhigvRwOf0m7rLO9ljossA6zW6lOYuq/ZBBUserA
7aqmOQUZsYPt7Fmj2KwdQy1VkJoIF4MOsBKYgVL4eXfisODijMIEzMRECi8z
iaj8hLCwBwbpa4GkCFUkdbg1uRvFnb4AOa1kheMnqy/BHp337s/0vk0nGgf8
rvpKtou8J1AN/BLK0Ec8d9qTGtpJ3UXvvgEXe6wJd/qs/kHDI0W+c5luL+Tq
umuTlNaVhwXNYj4OKFcAri0fRo9aZ7IKtS5I/m048sexrf4bhqPqQltgvWiQ
2asso1HuxHG2AgqCRSJGoH1yqfkXchAYhsy/ZXIk3EsihNyWW5aV3RuEVDDO
fV78fUQqX1ExY87ZRfzRSpbccYMLcF8JJTfUB8FMwbZnMTSNPxZUiCCSDu/Y
ItB7VG+uNkXuUL2Wrnr5ReCjcxcM7n7Y7WJvzp/BgpOHLsZ1x9Kuv4loX/RY
V1RDRZtY28Pd9Lqbfa7qtp9Q3OOJMzJGpRjKcOusT6sDkYvQCTXBu6FnUaHn
zj8zNi/kHBK3jJPQa4T2tKbx3o2Wm6S/jTec6mpjWiI8K1oH4O9Ymuzru4td
BHV/8evZgZxpudA9GYPqSYHS3m+HgPxSuzfq0scqyGmeurfdWXmWh82tLjcs
30/5C71mv0ReD8fd+eDZFbej97BYmhCP/5Hmy0PggTodkiJW+4jVIhU71vbx
g5NWge3R1dhfjH6b1p0CJ7IUYyZ3FVkSJBfzm/eO9c25ZOD5roUkmc7H5USW
RuP63yHGP5CUoYA2OFWd8mgKFZAmaDCvf+U97zErwL+Q+vZrzKUEpclLAJi+
onJxe1lqQiLlu+S9q5bHiR6C4dInMhMDKBr/Y2nUaLaCYR3Macyb5onUpf6r
nrnrtlIZ7L5DnlrTwngU/yBBqSVrIiNUK8TCPoW7aCv8CjALYRNtY4Yr2bOu
BlHYUuz9jc4wTyOxYhrQq9EQi0ztgulFcQzmyTxCd9/KH0oXwEtuO2/01aO8
HUrCKC48gR2p4GdF95VYimgd6SyYcwf2zTQ+Zn91zDPtabRKRB9ZUOtaJR3c
aZewiTdDEABOK305ciUM6IIrd9yZuiP7B6Zx9BJlVrI7z/8B36jezIu+vm9c
Hg3ddEtHL2sjTMO5Oefs4TzKm2seLs/ZBXTdC82OdFWm9+80lUcaXNAS4T6F
OKDNyoNvK+xHDw+lY75ciamAST3W7vutc/WjDUIDYwWwFmUkbdI3ZEm8vmLQ
DFrnO/dF5qqKCUTJBGwUmH9tpkUcPv1Btf1IuwGznukwP1dBZQslNyYdhGnP
z1C24iO5BPcudBYnPA0nC/4rieiB1q9YmVJGLTKU63mUwnnnEKED1DDiMSqt
0ccUx4HAJNhnjgzv8jB9kOKQFZauX7dIVHgzSUYJm2q0Zby8ajq/7LetdFF1
VIzao4caTjJuoGRU5K/Wh0rJ6u37oRUk29wmZBTNNsGRUNIoXEa1P4GALL4K
NpO9JT59X7BrJecR+U5qdnf8n3q1Si9HU8grViUG3pzkv3KMc1xQ7aIJM9EV
eGKKtDrcbB9o5K4DBCa5cpNFVqu7nSbta4OWezLZoja/7dE2r5d/TgT7ue9c
EVp/8rRGPe7pqqMXsP1zb+dCS89gs/IXTfsMsUcz1CIEzQp5z/ngydQfpR6G
Yd8IGY/apd6yxdvubiueJ6Te8XPjyGvrLkFJ+nQ1uA2G09NEj2y279uD+Mew
sPRyhe22fj4IQWRQEbwYwtk6kMOMcLDztu5tVw5rIIhDmZyf5CQ8E7veYnNC
jU6GUC7WVVvDy2ChjgpaJQ5A+rjBF7FAOu0S2KUEBHowsk2531CkXv7YZIV7
kYJZxGcyxU6GiUOMQVGd052bLG/QWBA7ii7MmnBLFqwtldzztacABHd5Tfmz
47HwLx7JLjKlr5trrVL9+x7EjThVoctlcyQco5K/20wm34fulu0G67X3wVo4
Cy44IiLjWxWnpL9pohp6+oTelFXGIfMLwBvrI2t6kUIhsvttZnc1JOHjHjhJ
P5mIuv4/qLvK6oO3RSBB8UuXBVVbZ3AXSi5EQmJBzxeauWzz1CA4oYhhYHrg
zRb26IvyAE80EIUegqXeFX6Tbp63uQgL9CJyXMgJ3RvDfbuYzPim2PRDQTTL
mE5er/O2mA0VbPEqMlphc+3IA2rP/g1DygzvWTPtAy3oJrmT2Fxy4C5DSbzl
rS+cLLof7eUaNHUuAdKW90Y+mRt+j19VRr5qAhOZwoa4/s3XXo9gpKcDmR45
zrheMCN3aa8dv0aUV1uYKiqf2tU3l2DvjZEwOlDHxz3stFwr18TLqY7ZBjLy
T93kpq1veuHVe4ZizBx8ydIvVRzh2e4STigMuvILB/haxNg5vrl/PnqDS69Q
VgXXsj4ZVQ7VXFiJvxQtZCD2PGCPhCya9MPAzXFscSG2XACjH42hzW7AajpQ
3BO+BU2SMvHkyqDEbOmljdxlORmJvCciK+Hf/JPwOeVp0URdhdtLbpzVdt2D
MbTRP9B6ps/8JYXUCt1eb/9bKLL6w6Z99pxUr8aFV4PwWK0ZTRkBcS4o/qOk
3O88+COpGOagBscwkcFUxLCKMBFX+YAS0dhVZt4umJzgcS1H3seQIgmZx8jb
Mww1FZAKR9HnpEDf4Z79ehCxwFEpDpoRYLg5TwSiRhc/p/xCrXF6CHm4gDPj
bExM13XN0/WEXnFoON5kXAzKJk1hweBg8PZjcfKtHpdlcN2YumwBt20lZ2o4
x6eC9Z5zd8ZdF+HfY7hq3V01ahPT6z91xXS1xu/ZjZxfi9QtdfMMrNleDwec
4rClBuN0Stpc0MOGq7eXtgeZzYoWy8WD1xB739pQEhPo0WC0ZzbfiX8PtsDN
C+d129vaflVgPUmZqwJHrFNZQhXCoVhm9WWdIUSFOLeOrmKKhgj2x1nJ5x4x
ZSuKss3FhHxJrdOVRZ6Vi4Sij/7+bbgBkw1odCKV+J4IlySGryrLFNSpM0CR
9Ath3PUnq4+LytDYZjRTj1MKRKZNi77JWMRCz9jfxj3l+TRUhUZSb+sLEa56
a1SmZvvZtUTbQFn9JjhWnkgDt6tjoZY1bxqSCyAigjuCEo8Fw93noCp7hZEM
jsOELQlf6HiICYOUwaWhDsli3oPTwvD7gh8FkpgtCBa4D82DGLqdQWNNKMfG
HQ26fRFeXTZkfAbA08Gir7BBmoWhiYvR/OEGTC6BzgA1GG4Ivp6lzSFxPnGG
P6HvOXUselYVsxJnIpmtXOVfOKZ4l5hvKR0zliHnNTyk2dBQm5tWG+PEUOHQ
CR5FZJtI/NvGkW1DAScNprzRLDTjQfD/zrnUvm8hJnS6o1KJ27ZmkxcmVCQK
J3Ky8PkT/l7R7zsbICZH5xjWEFEPTMUYXbhwixkNjbUqKkNby+7hcwwtoJLN
NohT3fMKkEzkb6HDOEt8i1TmvTRXgszScBNQVmibTsfxEIV6at5KLBfxGXtx
r0CLRNKKHDPScGxTJYo4cRI0V6Q0fcswJtYfl12M7isciyBOVFwja4UTq75T
YSO6iUo8bh/B3oTvYQUm6uywfV3Q5K1sMszTln4GJYYDev+whhbkXnQAffws
qZ7kPxwbNL4+81oJ4oo/QR3On1vJVwAqRp3llHgvwi3KI1CefTA0zuE1Uybu
uOYY9yexsJzUFmORFdgZGAOkCwHztvqndyHtZ+x6v96sWjQ1VRWPWIsZVGoV
mNmSST+JCqBUetuxiZYCb3kPNZvYoBVT6MPXHKm2FLdoKztxYauA6Vz5f5Mg
zesvsJqflBVazer9CDKDnUk0wiX9rbCuG6nS/LecSc9Kr6h6Gqycrn9Fqau3
uAombBNTc4snsxsYHfOxfiwfTpu5tUwSFLZ3oKeYG9i1klN5MqADnZapC3Zt
N/FKAcvxuuUzyOAsW8ZFn2rmnQBSE5C6Rm8R7KDxPD+AQOECRKYYndqJNb1O
pubYoJTeyTyVLpU074JdfD8U2rxWzJKe+1J/9IAmoeFCiPTygHmcAwULfqYo
qirtWqezdxLhHE2pJk2jaTJa+mbSf3v8+1OlEZQUCv3MvHfsigjxY+fYSH7J
5QlxchsN5vK9qPpwMD02/QO2bOnfmpw6hsZzVnZDniJRXSz4vUsxydEOkBv8
LXjFdpZ8XG3R65WvINgTUq8ijZFEs7ABqIrSTVUuMA15W/hlUhKhc9OElUaV
5RqPNNi64ZkOXNvNQoayYh3FFDu4KE+3wx21ymMJ478wPH1PvAvUNHsrYqiX
VI9eIGTRFLT+vbzK3zfB/kLzMJGBJE5vDC/zFQo+3ltVHEbk/Yqo08nKEYrK
ZqfFT73ZzIUcWNO0B1mCa+WPv9kwn555PcOCl0tCD88vF4lTdA8E8o681dVo
jTKz/4fQG/ZZM5JFkVn+sURsDePNEzXEL8stKe1GmurhO0ZmkjDOed5/1fUN
PCWfWemoQ5Lnp/AET2K5luH8KJz/pq2DACD7uZsyzDoT3jKb038PAyniFMTX
NCVsC61Tk/dI3vnUZohypAOClcjGm+eZfwiXwFTos8uEWwp4Ss7Wu9j53TE9
wBlyn29q/a0vjJvyAqwZFspkK0yUyBKYZ8nIl6eokjjKoMsEvSHd+A5JrCcg
gxVhatM9nwyCLWZON/606fOGQzXFbgwZQlMdP22QuGUwd86O96vcksNyG62O
ouhfx4uW9akRZz2n8a6DPTobMokPiT70+IrzPMMJrfv5EczDOQ20Y6CvisVT
Uu2A9KtRwccznoRO+W1+xp4YyP8W3TDJyvXmMEgJBzGINtDzie1FzqBGP28n
+xr51nWtEay7hxinqa+p6TjL0a7lwDltx45AdTR2Y5Vx2bJ5w/VoDW2EDPX+
CsqTseIGHx0Aw8GbwwuM2wFs9sP8sVij30TmLHW54F6h5AY17DK1MkpeHtQG
f6oPFwW2sNHmpo5MX/fI/cMeDpQnwcgDPja4CQ8eOD1q79jCEPWEWtnWUmp6
JctNrqErTKwi+fh2eUP8Xq1gcBFJaUb9spHOd4XjHKMtTS8lJIhGxDbGL6Dp
I5eLPshTjBJoEz1gR+03n9J/cFMX7Nw78zUxxqw7P0lfDyuZuh38rIAkSPyf
lKd8an0EpRPt0HZNDps6anZYNVI0f1lSjFc1CzV/opx+8irr2v5vsSur0NKD
2PR7yYvRXylbNlxkFKQhpsNRRs2LP7F9S9jO6POY82k/X0fA/eG+fTaIoL4g
WXY2/uOZccwrho7IxPt6n3YqZDTkabVQIMjWGe9w55PURbO2qCBs6op/b4mW
yrBKIw5+JLLVwafjV1LzLUVtgUHCM9N4M5efekvP3d4Gzwsw5rldJOLAZ9UX
tYK09TshnFO349+xDDypLf1C1QrI+1KElTI/fMLSsYssCIvVYyOo4oKQLvYV
Z+tn7UyXZNUfQuvTOe9NJvFC7Lh/2ilg2OivBxay64zMiSXHdYwImV2m++DL
S8s5o7T4J50YK2M8ILhB+HTtQsykOaYQJPVU29SLozQ5626HFOV6Mqr34OfO
ptagqlqg1xPSec9t/WF97+AgXaRNc0eJTTmdC62HLjcdDPmXnCteAhvMiZGZ
3bevItDDpYpNu0KytQDlC3T/lf4kWGg/hh31/vDyD6hHx2rrwc194bLVU4tg
eTWrlCGzVcUOF65OsluhTe1TQD26n2I44+JWXsjzZBeAYqFM2oVL9f0rFw1w
zLSwNaVBsB1S6+bwiAFXO4hKy7aVTrjdaBtAwbgLvpYoxaWZj8JCUxhOgugV
Mmfh50mv6NG+qANKQ7SUHuAT7Ept/GUQKWix05baM3dPdN7FCVSUvx+3t+UD
0XKJ2avgXlogthewWZ8y02jhhCGH/moTPRb+/BWU7WniHo0f8WgCFTJLXYOO
WHdstmUQg5iq1LoK7LImqABF+i6/upnKQZl0Bwe1fQmflWXGk/wqwIkGaKVs
iQRF8quIhVo1/8Meyis1xHJ26PnNZ6dtubJNNJCaQaIu6qrbiUol0BI78Pu1
TsfIYPBj32Q8djdwePJTK3vV3E1buaPNqsf6u+xGY9TniouzRWWIMM3P9E3v
7+L9P3UHzc8aUYe3OSBYuosMxAQX4+QW8SNsroOIdi+SSf+KPKdd8Zovt1j+
xezPKOp6DexrFNwFwcopzjAC/8ac5zDq3d58kirkfUC4Dfljb5LTDxCeSC8v
y+mKdH2ngIqPKetStvVEvYojFoMVtmXHRlDb2tdD3AmDsZx0t/f4BEo0jWxj
ZT2qlhFtqtFikJdgVbIuKnpV4oii2C4B8A2JAD1n0po1FYmgDF/NF2X0JkNU
rF1q1Iu7kUs8zKgSPyymISHHUsJCsJqyJVn6zlJQPfPs+h9ayqnLBOW6/PUc
+TWtS4Wia7GC2qG/r0RdJ7jocrvenWdqsSuXn1p4PJNMyGgLfJH7xFmn5DUp
whcadx/KHaRF/EeVYC7K5Gg8aBuDzHImYi4/AxATwaDXxfc9ahb45kUl0BK3
+xJeHyqjIEem6xu02iuzDwVHR5Geu0flD4DIrEhOEvwhiyZiLWUBp5FaxJCN
XBkmHz1pj76t0imaCtoPqd2R3AuHLENbxLjjSNURd8UC4ac3GG+sqBLVivlN
r5ZFo3OrOKVSmrquTmhzhaa2O2/UA9MENMfD+PwT4MJUYWNFTkzdzrZccV9z
V/XFwTzR8iIzTtsBKw9X5PK5/PytsqEfODxfhGhPqtzlCsCwU7fnt593Xqjt
YtobC6unLjGeMDpWFUNxOvOOEpiHiFYWmu6AqifTCUmikozEuosnrZIEV7sr
owhL6R6AWN6QcWpyOIfdege9SDssYOAcwp6VXw1dphKYaCBOrUk+gBPF/1sU
ZH0EAJYEomsZVb5OIaSJuiiLb6FP5KlQNK6A322K/+tu5XutJ4/NGQ4Vc4uz
BUVD2iiwdlKZGOd5fQo7I4m+BkwKWLHzdO0Ro77kPPBe1f0S8h9TEax/Ec3/
qnVlJg7YowkOo4VwszRuSNbrxJaCSCq2N2ly71CreoRfpMG4DvwXjEgTJf+R
vzZ6jDAdyM3S48m2Js0oneBbwbeB9pRHtXdfPbV75PLLZeqVw4QpKR0Yo8Ii
h/LFsojUJOy8c3WslWxbUrhqGQUUX7lY8fm5xremGg4AXzBR1p3oE20vEYXt
OKeyFNjNsZvqynLi4dyYecvTDYlI7Y/w+QQ57dC3/1xwrEvlki5tj+EyYf95
wgmXa4YilwoS/Dkl2dusN7C+CwyP/mUDJZiNr9C1n6czDtlj5/IyRt60gwX6
AULwFZm6W61SSaspT/anB76w57g+EgYNSW5pc8BRIfoSe4SiUMzmQDy8SsIh
OnJtbHSr5AJ/qbxJfFDWr2+vTPPyDsAE/ncUWaZ8aq3K0TOrwb3egja1h1cf
MJQi8mld6QDExrKEJdOtMmps2vDfk9/vLnG1Rhc7knPfw2C0E8zOd8f1vBmO
W5GFevIIVcwi/vED/nAG8YiaxPNFl28xjzuMI0O77BCRevMmQ51U4UNbBupE
S+5sRJKKB1QNa6gFCRh2iL28AwBcZcmp2/UX8BIZpemk0ddLgl9K676mAO7n
sOOzC5SDruTS1sId574dV1EdhQWRlWyszPNnYjLDaBikRMvshA/ow+uC5Gt4
uYi8/9NAtRqjZTyJfUgNCd14hvpP1LadyVzgGLA4QHjBlXFWiNLnyBVS7nQh
diO4SOcd4G/gLvBMR8U4FOgLHm6DOP+f8hwTKpi8Jd/75a2VKYCenSzzpXjp
5vz69+Ttk18EWTjR/ltNGeowcyTgEG3e1WQdvQYi3BuotrGeyZSt9URpdGOa
NwSLpmJsC+Kf1QATvWiWx7lsdIKG+AlQ5NdUmNMMhzhRbJAoLgg6gb150+na
g9uYEeelkeBfkVoP06FITo28XVmU9tg3OHwpEjWiFoKEYpKKTxY/05D4TIU/
iJ1inAOSgPcTcMnf8H/F2ChmjBxNTzdUxyG548mfzIZos3NvkqjAlKsq2llP
KlkeWR3n12j13wG5mQk+wdZg8e53lginsmmrLKYEHRWGO1SDrjER+Rgt/qLJ
UxgdvIbblkqkEdoYzhAaya4eJVKbYGoeZJhBzKHRrfn0a3p3JqDbzNtWgLj2
9H1Ctbrhh62ljxtPJpM2ypVTcln1m/d152WN4C3hyyGw6xxfI2X6cR4x216l
e7qYdsKRseL3zWVTXtWO5fewAdX9TVz0GQPzvhRlINr+QhiarTUSuiE1l1P5
S9xHvvgXlIF+fUaNhvjnFPJNh1kty30kYev+fNT12JS4LJSuCGPYX4eHPvRC
LZnMoXIPKD4o+/BRnGN1bS77ntB/sSIARUSZDtw4q6hJ5fMK4wrasOAPUkxv
S4MRKxULGWvUdXSebu0RvUhbNsHx0EFrxgDvGhgjUI2MNROU6rA10CTLOtVo
VlACPC6ScTA=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "sTlVzHE+yhAN9Vt4a+7yJC9Gw9bfBRq6xv9kCe7Ng5psJnHruz9VrHCdetev/ZiPTJdBJQmffKsGhcT8C1xHmtnWp2phLrsA++mCi6ZvsisBHsXsEe07/2w+B8eMNZubT3xnRLX8hyEfcYoWZpsP3M1DFemdUhSKGBtblrC5P70SnbNX6tsPF3y1BZk1iC/CtfkXVJdvvd+neDISHf8HMgQ3zyVqVVLAWr5Qxk5Q0qSozsMWQthz9F4Lg8Wa60AsOXYert63uw13eAxN5BhjVN57B2wLabeqk1yTrzpJ+B4y+rbxTypVmaZ9hXKyFdFOsCJfcHm+RETiv36qKmXcCdqgqpkFKwFZ0Z8oTOFk2luXg0oqfyAmNn3Zj7GW/V+fU5sM6uXX8RGajbiFmeo+fLXVb1ziWcMUe1jMZqoXdLbh/r4jxT7iM22lngpACdrkcwK13lvpmEhbedVyUZ36qXqdF/vpNJf1b/HzgjJ0/VZQusS7SQp8vqtr8+QwcRZaVrXlUAGkTVN7qscDPgOi+yFXm+omsOjbJ7yzZvRsLtu3IauTC85DTVyReqCrKuo5zRcR8wFQi/BndMRAvZSwJup8APyCD1zucyT5vnMtsaJs8zFIKxMGtql/ML6Afi3r1mA63k4A/ieakUNM6nGN1Jx0RxBBQA7tJ1WCX2yVyYYON/hKtLiEhuxjvbBpayYpbg7GkCpmkXQyIymUvakzmizo56rv1rUWBAXDI5/uK9LUB3mCN2PFs1jEXgWll4sUcnQB8GmJI0xa+l2op+46xfHhYbO8/EbSIR/13QLp3Ncw490WJg5XRSQpWaMzca1HqIwBg0OY/kwhnLwCffJWe9SmqHit/3K6Nv0jBDHdCuFjEti+0jcv/3lSDeSlaYxdjlPWuQp0YyxT82b5UgslWnDsL3w/ds6uoes5Nc9alxYAtoRwlIN/bqN1SEfydWf0SLF+HmgzIAKLvdZEZVWpuH5X8kfu5hvsMNcOvQnnyjTPPuY33CXe4K0FqTwCbIT0"
`endif