// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GkibYju3MHvCo4XeJyStueTQPuIIy6NMxj7Az9MxD/uWudI4vcdeUWvsJMA4
YXaWXbeSTQ9dIDvnXGRdKRIF1/LzSNcCSnoTEVK4KTeDOVjb68+in/o1GCKX
YXsYUMfqd+0mUA26PJxykn81XzmUVMn9lBz7MZHM/JP8Bn1tOHOuwDHi1af2
rquRsAWyMeDBt9xJ+bWRG53iT6LZjl7mYRK8YAcim0sr3qP0ihTC/pcwS3XX
WcaPJhTamOfhzgXgl5IuOrVJ3iv1aLWIVN3sDfDgKExj2OXvv3iFJYlxg3pG
PQgm6d8Fe3P/30GUwWgQLzVw/a6Y0JAQXAWt4fAZ2A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mt3mQCgA0gHkCFX9pRB7Fx1aPWn0dweh1JfvR5dZYhPNvax4YHW4S56/y7K9
bWGx95EK7bkoZnRduzgmLiBYE5xsVNqJSP2b8u78fOVX9PwywjmsKtz164Ty
lFJazsXI1p+BgHtH1pxguQdAmr1Rd8Eizk4cCwDT4ljvY1ZQidEhOTk8ZDz2
mMuPGzVeyR/RUppBiwzSrcZoeqbxtD+Gz0qPciHdaz7DvZZg5zLwV8WPJD1F
izzNJj+mTCl0+Smv2LJH1JuEeuesdgbRcd+oWm47ROHKbDsIy3U0MdYk/LDj
0fSaqLXRb3dzoHcbTQ6QSmvu3HHE0xYGk5mNQGCTfA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OgQhqyOG9C7vqxj7Xjat79hncaL08uDXkipIToycZ7kyQek2iuKEIoZccEgC
2BUIzOQc+p2HC3v3dq+a57KKAZHACuM3LEExuVuQxgLJmP2myCFAU+PFFmCU
o28iNna0qVQPHxgrq26IpbTKRKazToJcUY4Gk5WHMkGGQPkpOBpNW+3FZNys
l0JjfoEcQtt4WRTTOwrDWKyDgrUBbXwt9nGfMkc2vbPP+eOm7MI5677mAf4V
GzLO27S81jLj65ROdlnW+7Czxh9csKWBOqilEgwcV/L14cexZTJAOUZ1cJZ/
yHG6TBeADQHJzh3oCUrxgC7Oqb08nVEI317wdyolYg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CpsYBGCuZiZ2ElOhS/dQrieT6xpik9gHsnk2OQefdTYANbMIJFKR7pyf3CTp
I7JdtmPQsHFEeVouHScmau2uYFup+QqxRdLmiAjNMMKKapkxBnt0En+6NEfo
6t2YkT0GLQV/Vx3HJO5qXGhTcEFaOPZPPUFmRREJeawED8riVpUl2WoABqcp
9hejYSjFtRCOYvwIeFIAtdW1VKVBzQFgLvA09c+QLImqSfqtwg6LG0HQFqza
tzTER49BB82Bud1RHX7dHQ1JekLrWwbHnytivFqwOz+jHPSPfXg0M7+W0SN5
ivOioIhVGNTBS7hpCdHjHZRuQWKi9uilfWQuUi+yzA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FD+BZwGZiGttzhLTL+TOuBAjPbl1wgcg7GCRleN5EC7gZq+UFcrGY7+7d6QK
1oEcHTmmDZ19kg4KaJx5C0tgsIYCGJJ2cbAQ+bJtu/BX5f3vEDWltSvo/YC+
aA9r+4LKtKwiI8bfDs27YtSRWqYPwC+3YleSVBuctiTZhDyE2xs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
TrFxXRDR6c/UXImI53jtXWxLvg/QvZX1ALbFGXBvCjvjry2VsaIYkmNEAgjw
1qQtMFxm+MyHmgpnJimBTaYUMdAtUJ66QrbJsmDLZ9eiNnjouAnwTmPj+ZYI
FewzwSS3o/3b+7APObjDJC5DTgZTLIQP5k5DmOes7uQPGVxxr3odxWtZfgEB
OrtykkvSzkpRxtCiBCIeiibTj0YS52n07z3p2ndIOdp51Avu9h4NTBWaTdCZ
nre68LvYBrsiBQiP/kbM2haoClmwbcEckV0AxBopotNWKRMFoNS1dHS49FHm
BL9KLMzp5Jriqqm8QrfycU7Z4/TzUunosbQnSodwUx6qoGsoN7kdYzWXTGI9
OjIrJTM9MPcyHW3IGazqIgGXzDM8O0+oBwh8rYj38vmytClPzS2POkFNLdL4
TlHnp4IAnQkHa/1MKUOTMhWP3v+gLy0WNoRJlAZik8WWqmYqyTp6GQ4uOxgM
u5itXs4PS7v+SJMmbgiwbW7ErKxtOEnn


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cI0THRk4/BBjMDSMjf4/cbyNP4g6Nfrpca4SXRYNNVcWCt8g597uOfyKBE2T
HZ1rt/+wtiMOkgzuXjmSDL5yKoodbCcNkTMciMWbcYKCgt5JsKOxYUS1dWjY
MgqTix0DN9yVllqoZUaLkVmm+icb6IHCX6nEn4v3elfbz066dJg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cZnB4/OfD3VnfBmXfQmYxHaVHMKXUIsPC+bxsmagWyKe3Y+t6s6xrulSpA7V
yftaZ4WzEHX+YYnO68xe9CjlTM3ORJWeLb2MWh7mTqIA3MLy0O3NRkfKXSMf
QXYtl5A6UShn4NPes9u/e16pQT0H0BJuFoEhLIJEX/xV66eB2v0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 18272)
`pragma protect data_block
SZaEXdU500ylr9g/X7+l/BgZ6UCxlKHDjxBedkW3HzMbHrpmSMCrUrea7lL/
7moU9uwGIdVYlNm7Sa9oyvMbpfD5h9FrsTw3JlFX0IXgb7kH3Qk7ka4frkDo
Pu7xWkjzCSllbfoRvkl/rKnqrzRqT+IS8O5Ea8L9yNH5NvU3nnxOCXwYzKeo
dMvqzapl9CqUKlblrnumFZRmb4vR9aGXU+50p8ny10jAIBxaZsjcGIB7QgnL
H/dKLxYZvtaPpkUF8AzDpB+tEUiu4FPT3gNscCl44Il/vk866yn7W2EHdMIO
x+OYq+PHqHY4vJHVM9DDEFJ0VRew7oInnrcI7DG9CE9DwJYvygBCxCIQMg/o
kzyI15hVYxN6AY8O6GODo3/Uagujy7W9ICrzQpxB9D6cF3bjgIA5Sa2VeZQy
F1lPqok8qIJp34VTJ7FnGziaK1hDcsPTAMQzes9MxOp6gXUJUk9wpjnBNk2Z
rqaCfo0+yCfkJR72aMW5YA538nVoRpfaMppn1T+2UOducHLRC13FRb/dUwfj
6etq1YTeaoaSiUwOEBChgLO8DAnoM7E3TjaSS+MKwwbQcXNui9ZDfOUyFofK
4/PUTAO+FA5LSBjOl3mjmZDEizhmRS+8T+sDUksMP7Ati2ERcY8OenPGvqYF
WGkp1gMIkUQM5r4hjzWGhAr7kU4BDcsTcO6fZp+lEdaq6hD4IHBeZ0e6L/kV
9+oGFL+dQx89yxZQdSRODe6HW6rmYkjQgtdwrpxsRE7GsO2LIQP+iLaBl+e3
r1vozSZdIQxgCqRRnMBRoMAQF8E7zm0lL3Lbi6K182xhg5Bcrfg/fWB23fd5
aFo8thiHreNx8ux2bAoccuj3Rb4qxqYB/o8Up5HHc5OTeSLWCC2ONfFhQYfG
l6mOq++RHNwn1IinCJnWSDukWXMeJqSBABl3HLtP05GweFFiFubE5bz4be1L
8lgUq02e/vOkjTXW3+T4bIpt2ngbDViUuJuVpGq3+Vs7qhWEGIDT2cyt8sGc
XVpDTGas5jDbqAvpm52mUSafaupK/dbBmaszQV/hXifcvBvNWnOi4TtKd9Wj
0Uyf8h4s9kh47ayVZHVezaPDHGFuVs3c+4aX1XQpXx+lkI+w76Qw13eaJPr7
WT2s910yLeMstDFB8bsrMVUOuJXCUh6NvgQzLWCIdg6ZRaDCv4wBNahkNYox
t5dpTDeaEpbmb4N4XlCScXpzOYncUjLIx33SFLbQPOpaWBHS0o9bp9ZZE5MY
J9aIkYbSPmNyD/NZahdYTYXAExRuRV0h3OCPVpHxn8p584VKE2s3b6sVOMNM
NC4cPjzg5maeV7J6wgUZb08eF8+jGfP/R9dMRbdJdS8TuobssnOEwAceacya
7pwGYQmYT1aw0USEEQXgEwnTUGZeDLfnZiqxqn4HG8Pb8MoJi3+qJiOcwCHu
uEaUIF+ac47kK8UPDzfTZllh/kIYHsor9UNuna8WgZjXJKB7eZa7tRhTZjYw
XuFT+KU/JP6xpe14hfw3wRRorhlPI0Zn8yEw+GkbEUZtnweOj48UNSbzqksK
jj7V73nTKiYizDbICzjNkE5Sr9gkRR+MBk7LcUJgwRa2fQLbBgFZjNRQKQe1
RNvZurCZvMeY/jAgSTgrhpsvUZtnlY+0L9tk9BQa3DyFHCAq9J0rXhu7pi24
cmGw5A0MhirJWRWtZkUcAYNYa09oufn+cYueFXrvKMLCT7zvieb9V9uFQ2I/
HQBuSIQZ5QIMFaFs1d/fUxJnY78p9AvGGlPKqFmDf31mXtHEGlNopn6LFM70
HHIohK2anMivIEzKPdxYL63uHFGdr7PzLaQxFr6JlMRWq2IUeI94oSgpRFpV
jYzMjKPJGY5b72I9UorzQkLEdJu7VXjP4L4iyJSkBvoopb7r+digbzdVkQdD
8B5Ao1H5CxZ+s9UloO4A+gB7/KMUm9+DRP7bd4r+xlKa6B8CBNuTgRyYuhck
rdwXfaYg9tgPlSlTEZKhmssIK8g+3fDAmJ5eBifZYbmOyLEg5gH1wc8lbtAo
JH4O+a1ON725qwTZYfepwejRI7Nq+zylwAeYK7ZkTrcPMXFMfZZJgdvLQAS4
/aQBxsvb9QcpM5vXEpsmBw2/I1sQHGe+48hrXn7+BUhMboLLB3ffBCH4TEZR
nc7ROA0/as7eFyfAn22WLmOd3R0Vzf5BDd+VF9aGoWQRrtj6hojW+4BU7mi1
u0sl7sFYiD5qZcrUKXpW46MXnHRGgef1hloQg+E7viBppPGF2W6kECcBKvhK
EBlJtMOs1sZyXpaQREvvxBpP4YqPXO57fEBc4ld4zy4tJIH+98D1c52Qwj8H
k0lVJcnewqaAHm6BH0OMd7YyhWZq4hF72zG2n23eYny2DBhar1AUUHEU92wQ
kjGZ0FUeVdVbadad0FA70sRtvWl2hXtVq4HrdMRrBcmmjYfxyHP8ets0xkN7
iUYFK4/lghRNTXk4xebq1XP8giCnlsL8XsJk7+Hr6Y6gIpYGJbbjha6uPxe7
na7smxl8W2rMroV4kQRzh47fzSRZq3sF9L2rggiFS1sp9Y6AOKoCYTNuX5GT
eo6gog7ijadsDL0eAFMe4M420yNt5i36+ukW1G2biDKUA5tAIbU8nzz620Qi
WxCR9uGQxvyYOg9OG0cgMO/MkOj6wHt9ipXcZ7C/goR0YgzhP43A362RzFjf
ZhUKqerQxbHBO0sK5V+8yPKfXkWBL2drqbBYZ96DnXaFNQCuuqPkm/yRuLDk
35nc1jQjdsupM/qWDnBeZ39HERF3XEDxmNh9esqNO1TzGdrwJhd2d+yK2MUI
r0qdFtdNNSJ0xKNlh3w2qmggPURgQh6TT6DLOG1bkyWiws29s5jlqwx8wQZ3
npotHXm0xAH7tebHF6PID3z+3jC/a16eUvy8yWZsQ2R1svogwWehacsSVHTV
LR3hlPBA35rv5BxJ2eTVFJZhuCGZXtfckGI8Otw4jHSlOYmbk+sq0ZrFPdDk
yQqJY9MsiM7NIY+/qEqTOJ2s59n+Pa5X4+heXasN/DC8BkZhqIvtlF8puXUk
Osc3XNnWOuB5SME0ug3udVQ6IrQJTKTvERfLOW/OB8NurfhL/s5bKxgmI6E3
MoCxohZJtles0DwNyRdS/q8rpu2tAcMGxH0pdf2d8ywthb59+tz6XivQ9Knj
uDeURIDWxhb7IAryjAfCP+7zESLppcWya7oZcvRRMCX90OPR6VRuYxK7vYtW
Bwm3Rk/53I1jsevUlx35MDTnFm10GvXaZTes7JfYJshleueU6jfZeB/8JQv5
InjILPcHoaaOglNnJKSHf224d1Vb6nWtfE58vTA7VPf48JKF3A5VtQ+d+wpk
vbI4bn9gzypqiAqPbWMCIXmrgMHYhoII41XfDIySpXQwP5Fl6sHhsCBuVk75
owuQXQrT+LuHR+/wJ0CQYeMCgk+UEQMi+D2dqm6p/sMbSPMvEpz4fO9QDJG5
HamkUACQJWFpRXV9+XhZp8NWiIDwz5ThBcwzvJtGoXOmeR3ffbcBIsddDtVL
CIImJzsbE2FM5BB3iyVbYsxdliJruGw6fImHAdqTxZX4h3i9270prxQsa/Wz
Hcvvv/P8kuLPoJ5Hm+ICiMe3pXn4cu2C6k6RGtBiJYX3TwUYpLSX1behkBAq
VVi7LNKIYgE080WDyP/bAHpuGzN3SxFnQyZR/zDxER2+LHuPKvyV/QFo1YHt
3Lrb/EXgj7jwrb+rmklpP9s9VrIXXmE7pYj8tCvRU1CfGhFMpSrJSuRUL8MJ
U93IBv9Z6ASfC6EhEQ215x9h5qjD7wHPCmweqBitp4SUpCniyAcxXm9sDTmJ
XBC6HfSgIYRdNXiO/PyUdLCCcTpG72AnVKAdDTMAOQ+foEaeaIcCXROIWlSD
uuHBMBPlYbJA+IVuQxCX/vNutwaKcAO278HwnE1l/rxJ150GU3Sczp4NNGL+
8scXs/HytaMvr38fAS33uwAivDMqdwJ46TeeAzRlU3cANmN1gyXfP3wyMekK
r0sLzh3JxbGocRUvBHH4nYUQnM+P1LUurnSZIPSoXhYQL2BbKYhVPjmsFJRz
4GocRgziBJ+QFZlpzr7gFVpjpm1T7XrJhtK1ge1YIJbrRSpJyHsveiQTjlgf
qjLSnRq3rrQliCdguUbEwQsmHYJ977ysnbhu3tYiD1+KnxDcRwhytaRhzvIX
pV90jCsxcK5NpGG5h2ng+MQwaMKPCwfVXYGxDJERKSdTiQ4J806RWDYph6J5
7B6smBAjUboIt4hBgEcph2PT9wBImzsWrBwazG+3vZyl+4CIQo98vmCXSqX+
Y9q4GaJBIzUrQyN4BW4jAAnIyV7+XCzOz4QLcbgCl/ccD9T3l00QVoWNyF3V
9IhPk3nKlQWj7N/xe+DIPYRSdT9U6mWn1Iq3eDrUVVwLpKePScfeYwmqrPmk
WSl6Dkl7xivOau8fCEG5n2E1xdbhl7BGFVnhZAJWR80hHDxZ913ZzByMKjJS
jFLefUAllAYJTCFJkAjLJGq6e1Y0HG22aRUQmSopT/nwReXXYkcZqyLLR3Dc
6HaD4Fjyw8gmmELPVprwPyQ1wJiqsK44XMSbg2ur0+bzVi1x6sD1cqWqxd7e
XX6O1OGa5Rgfu8NKab7KnwQ3xf4KYQbeigDrFI+EzCN+kw6O2Ns76Qh/WuGk
ZWTijbVClYoEu7HokCJB2blnbT6rySkZtO11tdzMKyKHqZd+GQKZ7j7ScXS/
KevkgCkIkuF2q4Wf4kix/9Ag9lkDxpKwKILc6NWg2EGDEw69O6mj4sg0Uj8l
9Io9tchcrHYPJ3OENe86feglCAjhLsuwAIg59H9PYVIqWgaoV4ISInoP9c1j
RiJjMTH2fifbWnYx45M51KzPj6xDc4fT9YNZZxbE7Fb0culUEOKs5tAtnAxF
P3cc361PFd9igFvMk7afG/sKtiibct6B6A42tIoaWkpMS7U6TIqqKXn/UZAB
E0WaGsKp99UXflAoM1AvwvrkVzIBnO58NWVIyfuWXl0UtYx9v3nnajxeT/8t
q6uiVVPandxTFHKBo0udwD9T/VmLckMknfh+KsAAbOBQHffmR6fAZOUdh8CQ
qgLJCENY3gr72mozeJt8fMsDBcmAUz98RvsIKLw5mwfiqjqMZXSUa0Rgg679
8p0OzvCw4AdQxQBzrxtbJA0csCrAMh5KbQ0JVrpx/0x993DQPL1kJSOdog2z
G8JpCgA+0IPP+XavMJOlgIBlsHT7w0Pypq9tqVz/V7yqCRRzp26twLKgvCpz
yUFF+F2YnZH2LZv8QUHxasJcFLjrQZjPUHuScmSgYCUoO2H5Xjqj6xL+5qDW
jNoKLRsmM5DJK4Xrtgvej0RhLQD4L3rASleTSsz1wu0t344HZoW0Eb0kGl0Z
vzq6hs3N+V961pvmRuEgDmrD9MW9fIJMtOv2FLj16HYZo+F2fcmGHIl/0wsA
5lKNBjERyER4QA50Q9Yhg4OlxUTVdkPh7j91ZlhKQvCoUmxqU7FgycQNLfCN
RIn99zMpGxUlG3p6ca+tF99f68sOY8kJooMK24aB+WwXmvCzaGygihA7t7y+
F76hGIDl1OlTu3u5p2/BDhxYKIFJKaEH8KSmkan9sUkAhU5lZRqwSQoWP4Q6
CIAaYSi4zMpQNxJnNpIo93I2fPXXWxYRJGWe16UP3i2oXX4dGKcCdv75QKON
b4LNrMOfGDip2GVB787Yr26PPy26RsIzuWciNLHJRJb6MMzYamz9JmYS0M2N
CiJzboVNDLX9ybDYihQ/xo8GNS68msACreYI4Xcr+DWxgE4+8faRIdrREdsz
Lm2PEy+fIy/ES0A44R0y5f/FW1raqSsHq9um+kYCpLjzKlNDP4nzEsMOolH3
CuSGtYSryvZwDgmhvadEGO6TIP7/MOMF6WGYDHcDbp1OHIANFJGxbrqtLYEK
U8+GtUEceGsuU3a15/NL114+0Ef+bvSzC3J570igo86Or4FkJ5O1eukN492z
gvg58mXWiYcMnxuknLVObs/1t9Ag73lCCKb0SEM3oKwQ/8QtYpk6LbxZno2z
JZWtIu2Gf1VlEbd1JiJEJ+OMBAjR4Y6Evm9z/sMMzfN+OJa+yPu+TZULimMK
kIcHehEd12tW4i6oGDMjUkBcVCJBdXmZBVdOn5p5WrwdTOwsoVl+iPOpXrHB
QNM9VxFT4SBVh3XKvz23s0KPqEqW6rwsSrLq42pb44Y1uBdAHYCjv/fiwEIp
ziV0k9eWS0rn3pTpTanHhhZXm9WtBpAxy7n9Kki92d0l2SxklpPthLVn3l6j
i1wlbogJRt1KiWi1x+3sM8oT35VI0M16pSPwRyMcygL0KQdL4VEI1CIYxygT
nHrDYEGFbwI/B6BEpNj4b6Q/nM6ehNiCQGVIhQtrNci8RtyDuoSrMG8pS2di
c2ttUBssZH3n57WsQR9sJLAdC1tl2Y4UyLrBScBI/JsacJ7VQAgEuVAr/kWn
UeA/yMN2Mg/OWlZDahbY/5O2cRg8kwT0g3L0kjAk3Z5wYO1gCiCcdBky7nkL
eVCb4N81aO3Z84zqiZak7xLNzIY5BA2NAjcNY/eUoAlGF1USFv75pY8YIsFK
gSGJ62ik6QY8DnZeoD8QmhizTdhgVqViUyiRHPGsGi85Vf0MA1Zz2ZmQpiX5
Dtm7N+e2bs7jRlKPbdw0T+qcAXXs/ZZyJDoZHkr8Dt0yb+Gn1seRnaqsqmT1
JAcURWLdzQEuENymdAvFNSg96G0e44ZhHexTBfjGX81+6fuZmJfWIskpSf5l
Vfj7R0FrDZiMqA6LcyQU6wBJwww8bM8Fa8HHr+XcfOnCCWT8m/nAzuZdJvqr
j5NUA9eWU09yHqDBzjrf2enPl/AbzkXOPublVq6kdbNadPbXLKoQ740AY4i/
RF2mymttpD3CCf69ao0fik8f6+y2XV60YzpOZhdQ68w/H0oMw0cFgz+bPTNr
erjGMsXBbyVwgwkToNfWNxrUuz9B1goKDuIH7iz88P7vJfQrqSn4JQwaHXL/
tvWSXZ223FZBJjBQ4R87rEus5wTCMizFSmvanHW5YAH0sVSZKOf+Bp0K6rcF
UhrjNKQRSsIA8ZD81y9PYVa9ZsvMDyGEmCQu3HjGbq4oEJbg0MKe6JdJVGGD
p01F4CJDBU6sEkFyyhl7nkpVZfsWsOy6Kyx0C8drmnSRBU2MlbRKjbVsdCOA
fPypVXThJVYx1g7+k4eduO9YwkNnr+1YE6f0r/ERH2YgmL9LzVwmYND/jKt/
Zbj3Hfvc37BmcHfDZdzlD34x2YXiARV8hDAJmzxhIONHK8HnHXw7RhTXvaLM
oqgjbbsZrBl9Ku3KvOKEbrIk7u5w8wrpqpZU58UrnQkoCS9SvP55f8mooa0P
GoZRkBmwAtoozYSsCj2DTcCF8ZBWXWuKWe6doy0pz1nR1ZHLiKL0ijgVAlfE
uJCccP/uQZlhqL27KTpw1jgMTyxGCQHXNCIs7AwC7a+8ocVQx2IWeeDeI/to
uo/EBaVSj0txn9oLsERYhey+YY4Q+sholiGy2KrxjQUoiDrkzrKNUwTynMAc
cYk0evLF32bW9yT9xLU1qFgNRkHCejGjHHudgAOxntDra7pvn+zo8R4hSTjj
sj8q8Q8W+4P/MxbIjx5fgse0fyNISRorDszgx2YNbCF0WVw3/leqcAq1jxDg
vVKzgEM9K18qF2jA09uTVr7r1H1zka5C0tPR9x4T2xigoWk0vKPI5U0swIq3
zxINRQ1U/BZdEB3SU/M7RsMsCcs+YTlW+eB3PlFcp50m0q08Hx2C8+dulgJT
yVP85DDo40lvJ8aTKvbWfAdToJS8cp4obOM0/iyJt9POCmhhCABNepBgcZTA
0OyN24Ghwh31rQFak6B1k5439/nmvOvdAQ+8wmOt6D3aO+YCQ3wfG+ZHr2eB
Fjr6CHV9a1ZWB8wNBelGdMcX1zQDqLN/XG7CMJ1lYqvWkmWb9w/A9FaZCpS0
luqZIzFVLOuPp6yF6pLWTUfBkXeVNabRiHhUmAdHBbC5ySym2c7L63JLTgXL
G4sC5ORpRT0Xb7Maeh/VycRgphyEI/e46a+oiYgQ8T/8er43PB3vkJlZ/2Oc
FCGWcRHkWB9/b0Dr386KP0FktlBmZGeUX44KFNaJx4UEikmzIQb9kNy8zpXm
wPXuDr2hSLflorSLkHMOy77o76x+1IIITRm2LfmuGiYeXVt2MwP9G7ahshSE
NEpiUJjvhPhBY49eNrLpFytq6UL/aOncpNYiCsOH1FXDg1SFEyHGU+IuvyG0
TYyT3439onlrU+JBILrcbRSqiuVYUxCncRMUitD0duyq40KN6butYF+RqzLk
/i8Z2YLnyJkCJf3gdjKdikfeYzBc5Na4J4ikkyP76S7tE8nGRFrJ5N3KVCU+
FJNf5F0H/ykoPBqsFNJIieGOD9uw12iTygQ8+JhKPRrqW3ESmE8WDA0B70IU
KSuk1Ef17tqb9HHVblOR3lCLXAcqwocabWNRYHIot103SfT8ErxEMYwMNHOI
HgLF2t7ocgW8ZqaSrbn5oqjxH64NfTedxABDJvAy/FrYb3+NJJMHqE2Yz9iA
6Do1wrHxkI8dbkNr7o7Un1JYUnanefU5ruacNHrTx3ziSFqWiabCwHyUBp8S
TN0r/IrvmfHlsq4nzQ86DlAZI4IYj1Gcbzfflw4PKgMFEeo5phU95rM7VSEj
jGmh2x4FA5bLee+S5XzitL3Px90MNrlc/5WvmOQK7AivB63HkKzN7V/XDE4m
vbzuVolKtXaNDXWyUZuPYyDD+2xTlmmvuCg3eTcc2K3yZUPNsVYB4mvc5f3a
6RAlmn+6xAK2V1ETw9EjwI8KromIkVPeqCyIHRWXw1ozsbHjoNAuvlra0NqQ
6DKIWYhVQ6jzzyJuNr/wNAXMk4B+frE24fhOzhdoKLLccwBUGcAWWZX/C99w
6rhHuEDNLRIjD619muWCs1CMJfL/AVk9atb1FsriAZ/yMRFAHyt7bzUL3twO
Sj+RUa86DJFjBMkIFM7uOfCvq6B0QAyp5KjlK2EhcKSbxnSkgnriFw6Si+Rt
D8hyRycRueQJnxmhRXqD4vgOTu3dOOmlE7y2VFt7FT7NqwOkMXXi3GO+MuG/
RGBYp59jfUMfFP+ZJ9kO8UWp7Nh0WRNS9vfTnrj5b/Zep8D5PyatUgKXmr/Q
AgdT5XtDgSxLmyM8UWHQ9ryQuHFM5PmW30GYT2R0MjpYnkGqY/lsa+2YNxzM
6Q68tTS8mMuHek/QyNY9gKyF5Y7gEYKpuUXagPw0pA891FolUpA4QlNgo1tZ
VBZJVNfbyEq2HDKZxDl/PD3hxcjwJZSyTHzlF8g0KVIrR5JivLF8en62n6nA
IxxeZPYf2e1aaiHxp3xjIRjmaYXLeD+B2wPdmipSim8eKAao97aj2hwV+1wN
QTEoCcSSFdUxkpshYZu45SJcR1r0v43mKok/lL/OVNbdkGj5Q/5C7E8MhwAm
+vjTM3jPbzQJ2fqxdy+Tp5ffL2ha7dLEfzvcJ0tTqogXQDS5vTjcw0LIxoOr
8h2sU4nTvO2e+ATFFCffHZV+AYvMWfrwVvpyMQLxEhc7HT/U5xRiz3/8vLKz
TGrg41CkqB1zSX7Kv8R4uDoWRszWA3HGmmTX21SDk6/KtrQ9Ajp2hk7/fbmm
ZCKLCzPF63QBA9JVUQVf/fpMgN/14yKuHTbaUJ+rUFLNmFPbjCCkHMoG10/H
4PmHJH6ySXBr3jswUoA++y6g/hdf+VrHKDhahv+TvDLuDLoOegI2MY3xx5LR
oK47G9GoBEOSKVDZcYJOBsX9CCT0l9eSYm8YVTYe2NhDCNQ8DH7Ch/imiOmm
wh4saw7uUG/U3Oj9q1DBZID3ZhbZUoIkRFgMHAeLQ1hPpnWtxnGZdvccqELq
4B7gspBy/UhGa8Yyvf0WtizfMExsVpyHyrvfVsdXUn+6Tx1amtJLlC7/Hdcd
bPje+rvtwD0YGhrkbosgXnQiRDouwetVXwh+75nSPDv++9Vz9hIRGHB/+izH
SF0ueAqFwynUFlZTjs2990mBD/66oBoUFAAD69rN4UTGd/tbaJqSh4SR60DW
HvvyujCULkLcq5y8LEFyiE9ImDW9fm4K1moVl98XYwxPsBfqB5Ko/glacZph
D+5p60nHkJRw3RrEw9PEMFeYKMa2FPhFKU2fYYI8rYmWGzIuZL7696vi02JS
NcO8CRchKeeV2aUgGi0xgLsbH13rshHwfx0gNSFR0AvEFI2elycKBbQ0isJ/
KZp0x+Lw6TGetPUcDRtmmw3amO1Qb8f/VGq8vFzx1CdlpHuNZXnu6y6Ne1mx
+LSRDx8cMWH6Z9yA5P5z/g5g75nwl+LvcO56WgPT1+bzZCW8g++wQ3LjUAcS
CZ/YHfRk95RraQGxbC2cTk5IofvKt2dNb06MK1NkgzBnayQAr9W04iSrEqrU
Y00jWSaT8dOu0Lykqn+n/4idrCME2EKD0KjI52EjN44/7z5kTktmdY1mumdM
a02JwxD/fQgll7qfZ4l1hkSomjX4z5HZZ+qazkDgnbs0/OG+sIDSBnqXBO5q
SK8CiQctHcoBi8ljkp0taV+eCuUJRpHAabSJmT01BRoo+V3UQSzgrY2vvR2l
M2A59zLEeKJ6f80IasRe7OnOOlvASC73iVs9b4ZfJfmWZJcxmLgCv8MhTRPm
xTIPJM+5Q79PsPyCZihhI4LPz030XilYw7BWP6me0HAMcJE9gwqL8gtooH71
tnqO5cu8DxkgbVVsJTIMJHjUUYuPtdlyooVaV+Q9gYYNH7+U0K+M1w8Oj2PI
mT/dIyNyMNVM9UlC22wVmU7K7aOn2sLT/IbBY1Y7vswsZYWydq6Y/ejwmi6o
vuQijzOeDn28UlEO5JvVjuIEsUhUnoXHezEKxwyukBtXG4h2XMn6bmSD5uq2
zXrSn89PcIIFrBieKxkF0/cPbwpEsDN63Qw3kr6eJTmXjaqiFCyQpWjr3SNg
i602xxzThIjFCu9+X41vlQqyGmn/jk0QMxVvN6xxe7X5oqaHQ8NqxTDhFDpI
PnaOcyQl6ARLKtqfgWhWgV6aBSoarr9qkJJtQAG+H5+1ZgefNtSR+r91oai8
t8TajrsSkrIJJE+TUfgfigEn7JqbxY5tAt2slirCEgGKU5rPAc8NzJqU1K7W
LY6Z3fKQ0WWT5PmWVGrbq1qiiKG9mH14mQ0J04IIoSAjEncSDhq9+nilcJ78
FeZ9aHHoIMZr+hR/rAGZWDs3Lx2tpiTRKveU7C2E8ETQ1rvNy5xopzcWTWBs
IQ4Z+HEv+478Vf6dhHLNB6SfnQzZssRZ7TrWoHzKvL91MpWij5Z1sr2eflLk
QLdk9tK7MccaIXBB4Lda7rbFWI3iDeM8vWWoqqJRinXs8bKF32fJVowA5U8M
VDk6/cawx/AcMxPOLRUqSMUXdzLBrZjSUZmLQ45HoRbbzbbPWwiaGjXdsOei
cXEHTHaikZKnHxpkn2YSEbMhpsB+quD10XD6T5JYA5MpohRhN9141q83UNu1
07UdT1RJ5Bv80sDJkoM1h4QwpasrE+X1+BLGnh3X2pX4N+dOGV/lLvjlPWGh
1Sr1DueuXqQwOt2aJ9A3Rw+vTcNZjVKnwiu3rw2ow6HnV096/I529TkHyQHQ
Gy3CrnIHY8qKTbOk+Nvn3M3t1ObZ1Oc8byQNlbNT7Pnc7xy3zcqCqz9flBvY
NiRYVhLdV6J3aFcwVx6LR5KCJUR5cxkufH3hapPrTtnXDd9x+FF8nE5r7+yV
BwRrRuSHKVOOLKhArKsSbboXwmE7Agvykl95XlONfleeb69V51u+WmA6gT6I
M0vAkLOwA9LGcK8PR1TN9v4uZyTDFxrHn8FIBpnF1MLPm0J40Y6wNtoWq1V0
xRPcDh32upg0nYxoxewBnOo4PFyF91QKXWFS1gSOGQlgJw8CmnB7vlbfl42y
OwPlYwDGPo7VBGg2OromYxPPtjCKiyWBXRyN7MUtRK7/faoq2izoxp/W0Fl+
HoHCyyWXpBzhc4N3rlrMAx99L32DtJ/gWM/NlpasphoNWbHEUY7GE3lquvVM
6Y89ip7gekK7lR5E7U7y5ZvtyK+/hEKglRJjOmQdsVF+gvszPedK01ReRv4r
1MDg8V0jWUsgcVHBRNUB4hKnWGUkjdKH1WTV+MjW5cepY0KqP6JsR6luMSU5
WDfzjTOsTJrRu2CdbbKh4YNWVWSxMbidjZ7kQ8BqelEYe6q6DHgGp0E1NhH9
E5XG63PC4S8IdCnEKgZNsvdvVivNAcjhs67grT1lrzrqVczeQDRsvXvhke4H
PPkhT51hiPD0iLqhLqc5S+XTpU0QiaNuc43iUXlz1S7oH/bx9TL5kZLqNx1O
W/+SZmTIBMZmVDnOo7IRdU/9vt1qzQAw6CClwhG50PCnKLflGK0y1x0HnB0G
4KpFcL4yyzvQEHwyoPnzsEU5NvFRBvtluYFWkKfsM64NFn+ZWy9ZI6VCa6TD
wS1do6rS23+RUyiApZyOjv3p7SyPFzG25A7pN+Xwox4ESeUmBkpHKqai/lLk
hcWoos8buuvi7o2bl3EHRsFWyrW2elw6HOCIwEbtdqEcI41OrCUmmEfhq5Vt
+UFEHqrGadwkcivi3ioSTTb/XsSjpnjJ0JDLDInGPEuDhe0hUT0jdkS2wbnu
puyt3IsUUPswKUnXaPJsyRQ6LOuRPtaL7bP0Ds1lHeCVaXjsHu5aUwxKhR12
f1+tNmuqhY6dsbt8aXPgFQ0gBPBIb8LBna1/WzA02+2XrCdKojKcXQgVY2DG
VWcKP41R8sWH2EMp1qZtWgZ7MSc3+oHr/vmIcci29vb7mSwNbwGtZ6UWjUdE
Zu/s+t+isYYMtihZ1a7cE3ey8UYe7QNVgLxYcYFOJLoNsNXyADfG6fTz0k2h
n/F5hhqeb3GuaGPLbdjSRhi2W6gvOSsSuXBSk1VMd9Yx4x2GKjAeEVnz6ZXz
VPLN0nwUJxVvlDqm7A2+qlZfq2FD+4yWVzcYxtOuOXh89G7DPr4/GspipCJo
m/zLtMWuOcPJTqGHJnzbYgHC91Lj3zTnA0AX2UUaF/rIoU03VWFSqrUoaySq
4PmHIA7qvpAVMEOcNwLR5OjfLbNRQnCycJrf7P62GVS59kcFMmTXNERasgDp
VV+zqWPGdqva6kt575qmrN/n+gO99zSxkS5Hx8+f0sT01TbQqxCOh1EfpRpq
YuzjUsd/zh7wpYntTaq/HumCtTBukRDj3BNKEEqCRm7k39BbbJWYWpPXvpDB
hIl61GS7rZxLMdhRYQB/YcsLFD7ym/3CegfX0ZEbPHTNwtn3xiaMawFsTQRv
UDESBosDxeA2SdwsbCQdy7mYGvZecr+eLV+EIWrvdAVc6MpADTAFibC++98O
mrht/C/mKUqWCqTUMGtr7KO+Zk0i+llVXDrZ3NHYPEFc4Ovm3nsGA1Y1XHlb
89I5j6gHL2ff1lvnnSnBcUBUph20ZD87oxZqgwFsXHD/ePlOEVRHkd44jtc8
eMdFwTVBAjzAKraTn6sc8uaDBuEGg+IapvkileHgjSj28MbOJfvvXEXszEO5
J0FtstjlwGLoKDh3t0c4LF/tZ6s6WZUvUn02BEOMhmBGUHBp1SAuOfobYlZ0
/NclX2/tyPqZfZrH8j0NzA3meSvvQundryB4QFKbqT7P5HiYGK4ERZnDJqks
aIdYiq4vSxq4zxXifTGBGoyVQGGvOEQX04JakpX3puLK/2bQVZNkfzBWvQaa
qr6tnmrRWYeQ7y1biaYW7Bo0I9+jm2623pmQOw8Yr3jwZQsqkJwqNpcMwqwo
WaqM8OKXlnkSqN4lDGDOTeUA4MIiegLAocWyMqj8HWDGYr5xpsDb4CQjVCIk
Di36WUE4vyVCk+nhf0sKlW8OL8YtkW7uCtDgxZYr6lyVLt0z1wL+8iFNMU7G
lFAGLUcrb9Xbu6NGs2dCn1fCL1frHjlceoZS6xImbR5cy80OASQ2lHnjlmfm
9M5jqSKUOi/xuI3+e9ROAKOKuy1dCGyTk+Giv/AADH9D589AugipOa27qQae
jV4MX9Bsd2H1HLD4D+VsPJO2t6aUoQmINL7Q+5buvP+m9u1KcuoTVoIRWAxP
6VQXP/aH5BBBX9SnWX4fJVxXG3BfRhgVp+rgAYeDjLhvBYiHrNyH4v4y2+A/
yCm2zmgGhQECP2CkgAI0JpKv8RR0phCm/D4sUC/zenzgC1XI1LOeESkPQuPr
PPmCw/qaL0W68VgJpo8xiQaCNqshFM3kHVzkiEL+vImyuWZ5xpN7M38xLvFa
VdDHsm2+R0+XnCV40Dpo/XjWV768kPtDPUUXwkNuKG8TUb2+tk4nX8Jw8j4k
nII6K8AaRRcldmt/XsqORtvG8aAW8ciWZgTguAilR3aOqgjDevrbREFRKzcP
PeOh7XldWOPH/GhcDD8ZfdWT8NmA8OT8m/iaPwa546s+zjGXswab5JuGDRWz
dEJjXw4GOsv3IfD38bDitVGGSU2YmOCX5vRUBWB1iCQYKrFRPrj+D4mdpIRt
Cu50JTQshB+0NbTnAcpIVjK66QcjvOj49mOS3J5FKw8+sPBW0VmZr4cqSMQR
X5MXhCEbLjBBKZhNgxmdx3Kc393Sh9/qPuN5PADZ+fcqo7Ly6r7BOUKtRfxU
olU4ktxRd6VA4j10Bpypdpb35+gbdLtfarHHoCB7DmSZXj3wu3zyPY7m/hUE
z7+DaQ0+rs64MKHrb0NXv4lh/162xwSQxUjCPUIP7hBfwTFGBrb529Qa0sLd
WfKP3bQ2PCuAylO2xT5vQk/J8tJlMeq3SB6Rn86spwzCaXX+XMf3YPbirFZl
EpkmXS9pyirbI6HSXNdMYNEHnQNVGZkW+ipYVqQa6pbSH+jc0rCxnM3GDBuC
xMuZY9m4YdHi/sUpAsDU+FWh5Nxsomr55c9Cz9hZnAisNbCkuCq1eLXXpvwt
YqdQaELYdd0Kn44LAe4IifghwO1g1hnQQBOHz1MvhTSTTnoagWiORhq1U7Je
8T+DnpQDN++m77hWSODZyQo35Uapuq2uDAK6vnnMW96KAD0ySkTwgy6XYywF
19KZmxnG5vQLKRmBbrh2x6agy/BRnWekjv9m1n8LST6ePFtvzFomHlRehySE
6Z3LEWSLDWmptmPbWw8Hb/NF4SThgi/g4vNubucsxlWxkGHcdGHOPPJvzqMu
O2aPiosbUXgBljbZ7Y9HaSbWvl7tQU6H2Iu0IaxUDIFWBEgTUWkURCX2rtBD
KiGceQAU3x0xn2om6KlalbdeSne4dAsUje+3lyoL3DmK4h+pJcTGi+qwd1Fj
Z4KnMWekHTonrWmlPzp5CGoNq8ZSk/UISeAb08Xr/fFvWKi5/xvBRQO0vpvg
mmXKAsUbD1ZePLLoNkegEZOnaa7HjrHjf8dTIzvfFMdpCgnXSTjYamxzK/LL
vvIsPphQVwN8zyA1wVDxXIv91/MYo2XcWgrTwGwpV8gGAF/je+SQKrV/mF9B
4YFxIXptmYqY2TQq8Izs0cl4FSZpqknJvnXq0kpNxuRm+0Vz3neitt0LZ6Pd
faIDmb0pbgScrBWC0lTP0itmOvoDKleAvVkIMVg2LhBPCj1O3EI0jWk2goKX
/t4FPLzGwuIPnfNKnIEbDnh41ML03yvMXFzjnI7DZlvoHntNZX3gEwwW4jhY
o+FSkv1y3DpsY3QXLW1olaKya302s/gLrklQkeU6MJUK3G0d/JWjQWVOdEBd
5XSeD5qz8VRcuIUQ6jeiIgEGuMFnsm9qBeF/W5zw69Eav5fcLT82dMaN5JDX
9gIEf5xIcxskWSW3x/f7VwvDc+avSf321ahgGQfYgmZ8preLD8RgxkJZ2ZE+
P7mHjNW3QULUY61qUtD9p+XLbCWSH2r+9OWruD6zPlo2MmXjVnHi4L/7P6wm
eVkQH29NTLigrriFaA8GUJ4+rxwmoykMfI5CL5f8rntDFEDKvQhtSZKP+ZEA
roud4SL0XQOWMkWGLzM0/sm9yEjs+AuNSpfVygq707rtJLeerUQFrA4R39r8
uybSrqgRcl8CIL3U34QzKG83qoX96kccnM0onDffQa3IKGwrEKthseUWxEzv
ZD/rGNDJ+V2BJgqyjNadoFuc1o/7b8moqL4hpnGyUqFzTtl/K3qh/DaILTvo
dK9KigmnE/cyWNaGEiMz/qrX+/Ks2GAaWFuMu6WlWVbSez0/psPwjJlOEx9I
ncunku35NcG5VmJvd3FKV3pWL/pRCahmZWowsf8QQSh4og7lKFNa2SYL9rzR
rc2BG/h7631DyMnfY9N23oDlC/9VWXYSIXKQdjf0U7ZR8UZWW/8lVl2BsjRW
9kCD0gj1qn661uBwz7MGgpayEWf1Oh8egn7XLsUb9EgT17fC0miCaXi/lpZw
VKYIKjEXkQh83T0TOSFQXeR4xvN8UDA/xNDmdU7O0vR71nAwPpe1Bai1z06Z
RuRlbAYNRZl2WtuNwx5RjWhYml5WQNyJ6uZCxTAqP2SjJG9TLjTZUGaEL+MT
CLyKCAv324DyESW5j+WLGBpTpr3PRPC0Sf/O1aMprSh+LNFeqFUINd060FpP
6ZVxZFyAsHkxhAZ8w3uZK1+dgugyG2DHi2jsIWnnQZRKn318Pyho2uOjL9Lx
RTac7oZ6FX9kmG66xKGvOUs/s6XNln6Oy4+HvdxRSPYXuwnr0iU6PHwdvTfM
uSi0wwzVE3K6d5JP/2xLzFUB6D/3AbpFDT1oGMRZ9ok9NfXp/Pd7L4aQD5MC
t2FSEOX/gC/VKT2q2rTELNrEivtzcnljfDlC/mZPAMaRoXNzvywr8GKlS3KO
Cvdojle+FywgU+cR9CIpfKrVjUrkrycWptcnK6y+RQHcmHgzKKtFDgC9VESD
sH4+x2UWga7yaHufsEtm05ic5Q+YzVZ+YXxTStybMxmTDLlF8JLyE7N2BkwA
zL100U2r0CMDzDJZFB9snfkzsQ3YEhZ5BClMNUSSzROqpZAOcbPGvzypsvXI
opvG54kmuRlwfAcI+kuHw74vKDZgyEwHuDtr13Sh/QbUzEwwLe8xphDNtTWs
7CHODFcWw04CFgC2RM1ypCBisB0qq2vzJq4D427X6Tz2cbaaQbUGR6npfKdr
yfR5lIFWx0b5uL04ORxIL2fqazU0ei02Xuc+YTZIvEltYPL/2u8o9nCkArUx
fJIWDFGP7zvLhwPqN34aSawR1itqW+71sD8/gk10YzfnAqQTawFtSwXILgfR
Gl/bgMbSJwiPTdXF9qdZq4QZjnshAJDqGsNax7NDLypWn31VZ+EWbrft8ZmA
ZYbYcEppCR+Ypw6na4SuMHmMM5tzrikszhfWBJuOsbjHJwHxDeQ/uzrpBNqe
EQ326u55wUA2qJKyClcGeqsWxQcRs7GBTnMA36Vrhrt3AV895ttsq7LIVI6l
2JmZa0hs100ScZS+l8OJeL1MzHZnKaZwcUCzjbtI9+apekHEGaScdSDpadnN
MnROcR3JY2u/QMYwx53qA1kjh8Kj196PE1p6O3fXByRYJLL9QgAxPfxL4/rC
4zA5Jr8iDPDbf96A+5HN80U3bUQULRsFjoNghUKw2kSqX2YjXY3PNdsPoNmf
P82jd7aAGiIrL2xXdwo0M3py3CplTMXQZaGcUkEFf4t4lVBRUqd6wPlgawl1
BE2Mc/QKgnA1WTkcngAj9qWGYz+5/R/OG5jGwdnrAhT0Bpo8zaUXjgB0mlaA
WQZozGwkwR+UjBOW+C1VwHdHty4TY5wHWdnRaqD6Z3dzdVCzfxvjYzKv1zX8
eESziZ+0Hjca3IoZAIAEeK8XTtvWaiAye3bih4V75V3Zwq+2+OxCXizmfhHj
24JD5X12vL6dwpTAE5k3/kBeNDixCef9OmmRk2O4UcsW6U0nw5JH0u5ErfbG
zSQHjod5KaQ7JKPu0nm2+pzBQjjCsfjwUTTh1a/KaKr8v0rsDdBJDmSBwA5K
QzPM604yWGiKEo22BpADiLcWORF8pceU6CgJo7vKrwMmRhVWRu+Ah5rQUgXD
XiD4bYMenypF2uTfUPTRLPSCUGYOeSU7OC1O8Eb05tkNVdmPesriiREcB1vf
5oQi8gG2fMvGy4tieBxP001PoNfXF+4D/wg7FX1C1d1Q/K9npkNAanmyoCYF
2dTeQkRr5pNEIKBLAmd4fyujlQJiEARdiHVFqHobtDtEV3wjkMJfBS6d1GeO
L+lXkUTu9VRds4HEpS03J98y3X03KY9eiCQG+n3nPuxpNiCx+dh8FvS5+aaA
emQcXES3VHCWhY45WYFykFLCNFz4jH2jhHSifqluUHx7YxO9B/o+6akOYVjI
d9SEB3ucytBWGQZ1TXVtYlSmMFZiR2hQM0zEZ1djaM2T+47It/3Ly/ZHCrEH
CnAse4ov+jIfGFffsUX2RHq1nu3uFyWCs/MPPyOX4HzqjxPsQJqop7WCWfIC
kvTCW/FKe/qI9a2eIHkkTnZKXILo5s8jb8/vpDRK/ozuoCMlV9umEoOuTeG3
Ccmqos/hRkjMbEuF0EaPdzwT2XOAnYspA+n1TIcHewC23nFwLO+7P9t2CNbR
P2t2pYzlVaLcLIsBCiqsNlyAKbmLoQlAuFc60qP9By8UlisxJfY2AGXWUJwU
UWIx/Iqd8aGWxVFAJ6nMH8whbiBOLOPnMr2Q0R+8XGHQUnoqzCZDLI6Fd41i
yInabVJRfOVteH3+aCpyMyPhKXWbv/X+E0J1tT4SUMVF0bdj5kvdaawyyV8V
1k8goesJlI1gXtzER1pKIvkNJ2ZXHioabUz9cqKtbWE49HHi7qv8O7NRIYyG
0pf1RqYVy0dgY1ZrNaiGaKx5rHlAYTl+W0Dv/4l3XkixzT/j8qArH9VRzvrz
a8OR+7+rk4fV1WZ/k2H6KKvENs4gWHwZXAXPI8VoqUFoHGsKiImvz0gH5GgY
6IZmmVtzw04heCg2fIJmXm3pSHt4zzto+xZoNH9AU5MHcOy/9UGEfSDITrRO
dLCFoAEDFu/nlD0V1RwGWn7vB1y7abf64rPgS9EisqWho/L3VI96eLxrFSbU
9Or6+9fytsKBVi7TbNgX1eeJ0MU9zsdy2GM8W7A7w3DZQKKDSt3O3u6Cq8Nw
3BQvuImY0J/ThasMeJ3BY6MfiKsD4qsJXhRfFC20S5Q7hVqEGMqKeKJPygvp
8LGCeX0fHpGBAOQk1L5r1L7LkHKRLPzYjw5oS1k6DemOFhHdFe/ISBUeJrCG
R2mxSs4LLUzoOd7DmJrZKA9H9tU+12d8zOmIfJ2sciOp0Paz3PuYGSKU40gI
OspoP4256A45c9fnI3HdvGxOWrJpMZHZzQBqqyGH9fYLVgpioAzdZVgt9QZl
v1BM90vuY1hVScsAxMRx0JJXzSzsFurtAs23TMEwQ2DIe3htRNhTR4+aHwnr
hlcgOVLniQmWCai2/DJOnuvmE4tT4ea800NGgygcuPTw2DHkTF2gfemAyr7g
c1HqxlUEoKho7CcIZKwG/ROjcPKrZwvP2GedQYfEPmqClSggMVcsdPYADCFB
LdQWCF0u64rStMF5OW7gMRPYA+o2Tf87wk+3NQ9GtXh+5AjaeyN2CmCtZ9ez
LlY7OmRTElSzkYTryQRJOw8dt0+9ZmC2X5PU9/K461JA4ShxeHTiQffT2VV1
oP+1jbzOoGs15DvcVqePNu7qslhKSWQzeK79c0gvtmnTH/9KDBpDZTtATx0D
QCupKlIYlNJQLYz4O6Da7O/4t0QtJ10IrDM7SxiXSuKie43Ro1QT6p1iGwd7
007T3on3BrILBVrXF7Ljpgj7mw+NIlODaQQHPTHL2fIhQL9bctQKKlpqjANm
f4mnZ26GH7eaP5hWm6Z9MSfBT6a/wdcNE/tyMzdgZF5IhF6j92YZHTE2szts
NjCi8Tqcdswh7IUYRSdodmwehEYT1XyTI9astl/+y2fHL2H6zY+sHXThmXbs
NXnpOXtceanFCoiJBQmwJmb5h6+YjvtzyI72wQHg74S6D5l6VkaNwbFrm5hE
95TfFcOAufJpMJo1nfRLlH6CJWNTKp+i3NDCG9do5jyWqqE2Js4nfKHdMdZi
Qez0jW4wG6IvDGbHTCwYi8h4leLD28C6IWK2Tv+QJMFew/UDoMKlngRutaEM
NRCSqcsSZnMn4yo8Ubm1vTvPvQXcKChp/++lRcJ4EiWq1SuEKQ+cMMsw/Cli
PYXzZjgXVKHFgk5PS8d3qBxeit01LRb0zGrN5qmn+6tatsUnZLkDonIakEl9
tZUwe+T8hCjhW43plRTQXMGhp8o+gj1oY0dHdKMQlC5gUhFBEI1CdtOpBIfU
YjEEp0+cuSN/qXYNIVU44FyMT8HDfNgso8YVs930K0g7Tjtz6+hXefs8YgsR
Btr6mMMjpGG0jSx0UJYTlyFCsDFNx3gy20lZ1hZhmHkgrFDLHyFoWvdJlImV
xzZAAJDfHO831No6LmKpkCZn+nzQ/lso0ZECvJriJZGUD8/sz7EffLUCz+mF
cdoSjmHRCNMpfdnGGUqusClY5E0fTqZN7uJiYQFNK8YFCWBgS712KHfUEjEH
PEO7Sk3UhLd7x/DOk3+/0xXP9cRHYgTaFPYuE97rVt6+qL6yUNLUOM7wovtl
QPdOG8Zw1MvxJ1U0e3lVX5e+TKaPENoyEgmhYW+BMifxSGe6lT3Qkpl05HzD
C+FEIxCsQCoUlLT4EkvjP5GUCQmx5xMiFf3w9Me6ULdyqyc21wdaZKU5Fvhe
SexlqSjciBaQkdbYDEZ1cMOEJ4VyhF20BIGScLWQ/iFCvF3n19HezBBExLLE
MKOGTZxB3h6pb6OB2tg4oStiSxWz3qIJRjstrtfpiCpQGxbLWo8JWAUu+fLy
fG4UXv+cEywQxdhozMa1YhEy+6vCtVfccV6D8zt/U2iIbGBz1d7xaZihGWiR
rWh73O3Pj4igwu5BeIF16/ReZvfdVxmi013jEIVSculTvBhRQEVJOLnfWfSC
yvzUsjKF/QFQ2DrdrnLuEfdCLaRecAE55MONmnEZ4N2kCKZRb9MX0foRfwkT
pHTnznVad6PXVqKqkGnnVPYAyvZq/hhZIPCcvsY1raUlhZvydMDX1fqu3xYC
KC6RtMHriFmXQQ9QZWgjLQ1W4CJBIqHe9Zt8W1UF5XRKw+pCzOaRXL9yJMDB
Bhcd7WQE4N997Mb5h3kRpSNvb3ujLD8Z3HGHJKH0BxTP3Fz6SBlpND5sxbqn
j0Nt9goUPSz3lLGdOxTXl5A0i7bN8z9xWAPAHbd+EwzIYmPqhYRh0Si5Jo2F
NKE2GPrbeNGYZETgK0tSaYXPS0q79Nu1eGSNOTPvfWGUKfk28KnvtRcv8WLr
HBKwLzTlwd3Y3+MDcA/5Sg7TQKVAM40ZYOv0Cv5l8lbnSpbAUysjL+DSe2U4
jEFsh70RQiV0p3YPNoGFhAZebAHK2+IikumGq/CY+AwjCFSIRAmxsXqPh8UT
A8bwnOqIR1qhIdrrZztOsBAEwgAKMIDDfrODumBgP6J20P3v01jXRQcnByOv
eSY2ppCISnIrCLNUhex2qmeNwtXZ7XtM22NGm/s/Ez1sPBMUs5o9hGyv9MDr
dPi83phfr0obo0Uz5IOTzkmZjBs3dYvWzwaGtpafQUni6i+Go0KwKHyEos03
D2k1BJObAYax7opEYC+bG+Qw/s6StENxZ5gxf0bIQAS3EMlnrhCG25qnhYXW
+oz5zTstL+0H1BNZ+KYt6X5CoQGrtv2cGzwIZuQ3fBRnyVx7Qm++YgQLEidW
32x4oCCW2qF+8NuN1p1P1uV1sQpKbEii+LFNeHCOPjNL7y0i5MPLpq5cX9PK
wPmNrgGwqToWoX2d0Mwzc79LVXkVOGlNjhgPTAxP2j0IiRkBRxUMVCwA5dj9
fEY+70H0jyrZ/jhngMawl9sQQ7EcQEHztHCDG6634iFvVEOOlZftyGLSgwPd
s9YJMaLpszDDIwrdk2473GJnd6BQ4u7CF76NJHIYmIdedzw5IByVC87p3hc8
vY6absRv7eHxgeTTcgOeqLMPZjPuvNovM8NpMgjf2H/s2ALE6OohrTVl287A
wa59vbe5t1yLx6HtQOTDxUDpjzFjWeeE4rSiziGC5O69jPV1WIkr2DpnGXdA
Wh1s3v7kSMU9gUejJlTTJML0wNP9JoZzkWu+qikfcDwr3dQpgHzMdBsLn808
LGsRWgHVLJNDlujms18ASRl///QCKHup4leNZWFwLa2Y/oJ8YNwJmZNveFR+
EZdKFs10RKeuKWnfPHqqRoWb15maYtl6+CdFbX8bJqOPq6ZTzXfDdRAesl9T
LoT2O2c0Ar/E9GUo3t3tjUg6HvK5O6dHCS9xcthFAB54yfqiFh8Z36Xtafq7
nBroNaqEeML/iXC3ZsbvCBrf+fiKi+xMh/F7JE9lTgF6dU7A7PYP4VNsKMK5
vVzCB0TLeapIcsHmeGihxhfIk9uam+pcWkbp8xskJR23zadd3P3ffQnwgH/Z
CwZnN6UnDHVc+mlFHefSRZe06oHu1kWtpEx3ZgHiGpnzjyILVeZaNNgTLJky
t+g8bu1VWkxkdOBchPWjE/Li2Cqz/HKHkiYapkcXz29lfXYA6DBbdgkJ4zac
djCcdiNROqU1S1jScy1EPe69hwl9Gh3dfw73AvAz4/6zNaEvjfG6RqOeSud8
Y7v2zofUyXHuPMamP9LluZZ/mWWP+30L6ZPSYEVKh0YOl/vWGsIne0CaMsYi
PoTXleDNuPCzixVKyvxq2VXwjMyxkvc4Savyi3Xyb4IUP+wYXMc8fbAZDk3f
9jqeUt2bebbj+mZeUQ8FpHvD9CW+usJ6jEs8/vdVYF5xQa/1YNkIb17vG9JZ
zq8U2nX5ePwRgdw2QxClW7CIAnFeZF1mk0c+jnEoHHHbZeHUVre5LLYA1+8t
icIAwFqmgkc5NILQm1zrVDeVegfN57Fd8Gkg/W97wdh9nqjP1b6gC7fklYVw
zLKqqkU8QzccrWiCQo2fUr3EyItfpkYQvJ48Tk2E3LQRscboUpeRAlxt1v62
IcFZ8G8D7HIZkMDRp7rkDHSzRq9RXIQGHqVh4rpDZBi6CR7TjaZ6HCQM3+BG
XiE1jUI0niw2fLsDJvMqI8ogPOpNBD7DQk08e+OSJNItji7CfpPdKV6hXNpV
ipflYg1djH/38IMseptpgBis0xpwpcinoDSOo6OqGdozM0NnrhwDo2IPtPNG
PDz7nfXyEW7Ovl+J5OksnMeZPf0pa4JZliRIriEDvu1JBQS//HsuZ986iZq7
sjE2/sCTD8zelxwB7fJLgARMRm9VssFlOk+UMtudNe+K5lNck/KOHl/PnF/l
wczTPgDSeU2qJaSOdv9nVuvXZNM2zOs49yu8zMdzAjyVWTHLv0UyHUWCZTxB
bAsnzDCHD5I6WyvVlPK3ljqxBCE3vRLtci9E/Fhql94tazLN/03zREyCpCDW
io6JPTPp83DEo0DP1f7jGsuBkmgSg0WhL3GlAsM/D+r3ZuSVdvmTURnUObkk
BBWa3hARpkNGADeP6wwnaicWyENz11tkq+E3xQRK54Hzbwmg8eWFeqAe/q/P
+KxI94to5x/bCSidI41SptyN1DJx0L678JihnHrtSz5vv2PvN0rjC/GmQTVK
44OVgScvz6Hw+ZnR2AiIIkkd1LwmyvP/LKxxgVE54PWqQWDYs87GqaHOi0CK
s6hF5I7mbiP0fn460/UQh3faF/SIy/0BkiG4TWiMSVzBubhSEg/0vxo6/507
ys+fQZZiGlEhXkotDSF9Y5uXk5CnGZmfuSFK84eOWZ2pXz+S2w9JH/zihnGS
Is7CKyS8NwW1NKWYXW2M3ifViNRvpP0QRLuU8SF81UQm7BIYvxVjGxnhhox1
wQhZ09wYzGzYn/Zgpkl3In3u+xt80qLJw98xhNe1jVzGJUalxE6o43rurxlD
a3SAnpVFjwEl+nmYeGiTI89fzWEqmxxo9kvwr1ZkA0Jmi4JJPpN1tjzawgi3
tSpUsBWEjZoRnZnnrsZozraPbG/9gg2vY5EX3gV7HVnvui5f2qD5EXZpyCHW
qJpMBpL9n8Uowrg7vw9WkIH3e08tP8pg5Ad+q+hDyaDutxwQTEKzGfFGWR51
NiKGI0Ae0Pjg5Sl5Fo67lQafQ0a/1eeMM5i2qTwH36NfAFNQA4+uIJg3PvHO
egwmrLp7jqY0F4cNDUMizVVLoiJ2ZGR8m0L0x95xFon1F5foijdWdQyL/9fF
zY41EXyS1lfMZ0q/nHhBQ4cjgrQyT3nG76t0GLwjKHr5x5prtjwhozG/GjIR
2/D4XtWMM6GbJE9jiP99L2LndcaHHluHg7JQxG1Bfof/gq5y0VRwVikvBC9M
jrUeoKsFR5LQ9apGRnm7Mz3uk7CdJR09LSqfL6ki8h+yTVXqLz+vBCfHIPGv
Gmg=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1JfhZcgfVXb4TmD95F4dYPYsdzzux/UC57pWitYxG7oSJcO2FelYvnsht1LpFop7jc/pm9gPkyWqWezmbtyRoZvgPzSKFNlErQXeZvp/WX2LLcC2faVVK0gkwBEizrp98RyNi4kXiyJZwU9gIIdBoymL2n+kQIHVH4EdFpG+uxNjJnnKuE8puXSSovplJ2vQDoqgrVn84BcarqHktwkag3ruz3Bkot1uZORvQiV6ys59XjwhIZfTCt/jHgSsIykmwXYML6QxHYSdhATemK20NoQsMCWF3eHu+MSCj65bQh/Mqqk0CH9fAhu63JEPammTnNMVdgs8U3/pgZNlmf9DCaJgE3MH0need7zn3R0bGmwLJmUwNaCLzqaFh6uKVQC1StYQJhrdiB0Wv1Yz/hb/gxDX88TGwnwQTFXH2KIze7pW4ckXrW3a2YhvBf+U7ChG394bY2w+GPs6J4MRfmTP8SX0Iazvj0EiyIi1CN/YUWqO0WAhma++Te6R70WygoPSimV8CXU0ogPSeiessFhkQQANMDuRQu/knZIURm0BRThkpSN3QiUSc2V/RematQkmEIWKQSj/BFWtIGhkUYA+G81cGe9XEhOrx7+iCffJmIkPbN6MsagVg/8ryfo+SwnzMS/bg/7CYCktaCm7XzZ1+b7JClpL31cGchrD2T9LPc/myfm7SwrbluQFW3LXbDsxkHZtVE5qipKTjQm96azudinRqOUM+jmW4VwzBEfiBtbM7zyF2E9KY6rQR3yQHW6SwG1WHqcMaJgSGYonBCz5TD1"
`endif