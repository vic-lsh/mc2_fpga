// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
X0UbXlbNTaGGfAQY0LUdbUZci0i2qQnF1qeVqYwyW8WZPRTMAh9jMpkO4HsD
F3/lpOZmfHm30OLZ7xOYbk1BDUnkDdCoTSS6IeFTrdTiW3UHzYvaHllekRyX
huwMJs6v18JlcYoV4JsQd2MwiLNbUB8922Is7kb5w67SzxLCd8Q3yCLFNdhY
vgbnoiNpB+0nfPgaDFJnEAfJXaOA8K6dvtx/TWg/3d6LqkA4ml0JHf+eXPhv
ZKrQD71Cqrt1wiJTI6qoVxq/Jt8XFwRZ/mzBtB3YzJad4Czr790vDzcyOqZd
OsUVq48lUjPRqBfsSgjCtwQEUMRWfwPvcRJSz+e9tg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hHL7huegeUqI6bGC5o6cg3F3SF7ytYYr7PnFmQucyZFGBF+YRDEROd+pKiVx
FBfMLsNfiy0r2777aNWcOObgUkX1AJRbbFw5RGJUE34KaZJZsCUaJR5iX4/E
r9qgxFq+M7bapQPdE+P7RBZ4qbFvjWeE6USSbutNkgi8ke9Y+2FUr7MFBxF5
k7deY5qv9kzmqgDBaASP51WzhqAEcEyE9adNMtz67OwOeF9BUKTzhqYKbbmR
nzaSxanWvTENSV8mzVG1WXpO5PuMi1Igi5fZn+0RmPWIXgtJDW6SZL4eEF+v
ECBkYN0pcfb3LARSXKkZWBXSkyEcbSP1pbw5Kz2uZw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gPz6fyKx+NGyrB08HENe+Wh9ALNejbeupmLg9ltvqQMRaHNNNINBipsBqTl+
C8MKE0Mh1KGX0G0aoIGv0/6Jurgzy+hG+mNjMex0B+4h9y8DACv8kuL1Z3B7
OjOuV/3XPuiWI4yunVAA2oOAW9O+UNgCHyfOTHJLdR9uTBa5iSXtBq9y9mAV
6lYS94GTOnSgrL4+XG+gRmIya0SHsMuYyc6px33YtZALYN+ePfFJb1dKWazg
l7H6ogZ/ob0M04QQzRAHgU66DLjapg52tFr/yvL8/0ljEnD+PXH0m9EatJ9N
a6RpNNuGSABpFN8hLGXLL4MkcMEwZN/+bjHbJo9kmw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AX8g2Ou6a2WH0DKQStpU2ETHftUbI+87QvV+otrNsu0hH6cKe5tH9sOEF4/o
fgCJEx+zby9CDt2e8PnSQnToOQBiBFiwAIcCR0yPzXULafEfdFyzw8WY19w6
2Rqp1tvxNNGRKqq1waD2DYOmOvuD+BlDKseHuy9R0KfmfmdA84UOK3FdYQS0
gFJR0VsHtY1zIWTFLz9z8rt55NtHmii+KyxC/QpeTFAKSVTboEL2hjOcmwUk
CCG+GrUCUQ3YVWRGNJ2SCVP/qJ1nNdwbz0vB2AfX+7sliPP+jEqriw18/4ww
0hLMH6DQRFZhZ+0LC7cGTQeyRcEg2Ubbf2yNzwIEiA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IjzkEnfK+uWe0GGyHrXIkwlTvizBps6B46hYtelHm9SkG4cViYSC8JWy2mF9
3TLJVUZTi6shUefeGenJGAKHjgRlmuHp68GkDm0eF8m2uhkEwXGCBQ1xk4Dx
CJVoBDfKQTIKKDHlmbYu7LxF25DmGulD6N8WUZE4JzuAxN6wc0U=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
pl4EdhhrlFosKZQ6pOYjtjwu1tivmkAxetMLK9BUmTc9d8OQd1MCxa88vxWW
4VRd5qF4hci7SLB1UHkJwysCyVXeyDvGUhAZLNxgIFf9vBHvEecKs3qAJKHr
y0E5qkp07aizn+pZZuhSm/jmPE9R0EXOA4j0J2XeIore5tpUrbdmC32+zAbj
Ikq/T9swxLXmyiKiScupXcPYsDYTGmtsDoIx9d8iVwi/oXrusuZk4JcRP9pD
AGV7T1gA7tuJFTjtItE+Fq4/GL9pkjblRMdrkWS6nuhueek5c/W5gqWgRUuw
HqASFiikg58RHuXaXWpijqjnbl7vhYXLHSyL8f2PETWC9j+lQsQAfeZptPAo
vf9m8PXPJF+Tj6L52Ah6BphKEf8ImyXl7EKJqOzj4F9Yxx9oqOoFytF2Cb3z
FUUTUfuUHcCmz/hOdi5BxGb67mnXes/JiCpDG7PXbZC6JFk6L8VPykjUzCDq
Th6kBkJtPVCq3lOIINqF1DOyhQU8n4Gk


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VnG+cttjxmAsjOKy4Q3njIZuKjCBa8HEmndjkvKb7k5nDHtEGRPul8kTcRHX
yUrxPo8NHLEIJJLezNSYVBPNBObmbA0iRd3+F1xOLAu/tcaKfbZaHe2hv/H0
5ST2gdBdKM5Fv0+/u8dRfew+JGZw9BJBaIyLfSmzNsrFh/7R+oM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lSJiPI4Mg4bFoOWGdL5LOQ6TAnsIO5VGIL/kPdvWEYP6D1MB4bZ0bOkCbd9O
H/gVka4p6vsAipltHhEEhOCw+R4XMTRCmUQS3IjNjGPyw76cmKeH+ljfGHJX
1XHI/9h+zt6zphjAL0fxtREOrbWLO3vISeuPYmDkxkJ1Jwr7mj8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 15088)
`pragma protect data_block
IrYCXFIExyCLSTD/GCcc6UKKJ1lfNQWdvXH9D6lZCzqJSo7q8AJ/s5qI06Ou
IESUsYELYCpoYfHh9tJgacwULw3O/tndPY/9q/Vgcj2Y58jYuSUGl6CPwOCT
dBbOW56r6DkpAvjIa9RggtRV+Ys4SoYG18QJnHc/B4MFs/Wz1WqYOzqh+2Qh
k1FxQTyquqQNBh3WBeE9HAb+4UfWx0xI5viNtuy4qhqlS1vLKmwZOYNsNfu5
HkQyZcra2TFv3hvLVf5pIoZKy5nHGMWzKExl3YEuUqVhaFtfUKlr6ybpA5gz
Imovim8iv+99lejp6QrPHiQIItioPeWBb/NUB86LbDXaouls27V2cobhnleL
ucdglZcojCP/idnlgmoSC8ssI5+i9QR/cv1RaTIbJIdj7L6YPYTB0zSXG0Uo
ZiEk3fLMZdoD8jvEmFhMmzLVId58uFRaC/H2hxkDW5iZvHzFmNk8byoNXw2S
xE0RKbc9V0qID7RcBnU9SLhOya90Ev95xszGhdD8zCIPRJ5B7XJU8cbGxwl0
BKM+YvnOlLy++V/SmfP9hPNNiFag6RXytCZ694sl52jLrKYMTtY5xysVF3AC
4D5dcaZ8SrWBJ332ToSiRqaCqvZnTe+H6HC9TPOkCvXr+6AtZ0L4xwG/60ws
kNnQsl415aM99AOVkUpk3iu7RdLL5KbFq4bns7z+csjEKJwamvneEHoyNRDS
kUxpEakFhmP9zQLWKanU6vMI+Hmlp1bKxRVvK+3VI1gDb8F+3/fcEZFULxIj
XLV6TyX0CwWGPqCX9YhM7Dp9gDaqyJlXs/41j5Ug0rDHdewfQ1L++vS89n83
D50fgrpMkjQU5Pzz89ASCiwyqOCCCYKT66k/MwraF7L3lrEeWa+6FrLbv//6
YPvG7Ih+TVBArBNMLJiOBexd7qF8+pPiHGoyB0zwcvuZhIGiCq+VzfkF+QgJ
UV7eFb+fnJ42c262oiCssGwA6rtZRbs2oADQtBHq5F7YGS4f1YEYfqirT2Vf
/lnrBkuRRlOMek34wwJeP1gTL4znDdPIM4PVS2a+8Gk1xP2B8V/wUGp5mjG0
kpfADQAaywMn16lJwNEW3mDrWK6B1EkWXcwqe3E8+OfnSmCs927+o7l/P68c
o/asx9FeDWnH/XQBoU+0m9K2Qm+rtRnestpCYD5ywTIi9MgGrHrdzhN0aWIr
uTfsg+yd4LGxSzQb3WYO9fqGWw/CplZfX/XBzWSik7scq8VkHyED+uCV1jdZ
HPd808ITcFlv3JOiL4bkcI6Cit/sZCZTwof3hBEqJ4Z4/6BjwpMzZEeRr0PR
DOMfILHEgwj6TbwodDhPyhD9mSa8/JvtKSlCGRZrbk0m4U0t5F6u71HU54om
R3SiDWBEqRofD/Musp+54eZTSi9hYiW44ggqvHUiTK/z/dqFN/mAIHbDaFdP
8pZAO/80JqflzaoNS6aCjipJ1etazBKfb11ZTwv84OzFubwsr1wmdPpZGt+U
ZIUmLyocvsQttNOjP6gNBDRS9ZpldGwInEBARcheXSc+NYoC2vgjVlfyI+kl
vexZgW6rxYB18IMl2jDuKsI5O1MnSVXKLGLbL8hqursrRIFCH6Nf9YSKwQrb
Hhse5PhX/e3ACMxCHAqEn4i80/9tduZfQrgLfqO26vbP3MBjQKJ86PNLI951
prbYFxsmIyX/kbwWzncNbTz1w7zojLC+Hf+5cY+8YK0NZwqquX3gE+IjuPD+
B9N8E4AQBEC8AfP0XIhdOKEn8ieN5mA7nWFE4o0o3zz45vEL7tqqWZBPpEYs
3yLCTQfwc7IinUd8Qo6hDxrTgCJl9W/+4wfSFo0L8x7+9cRLTwPAhnnrUIFW
MU9opIY9FvGa7KWXFg/mUHW/mAk3/ZWdkXFJxijkzfMdg/tt6E+5V41ZJEBj
AyQruU6dijnFOvqUmrwsy+EDjyZoyJ3/SpBcQ+pqOuIWpX/mshvSSjo5946u
zq/6JvMS4Yx2iqV7AstiNwmuYR7hZi7ivCWa4r/zvz5vctIH1B3UcQIEEpqu
gQ8LjgDptcLUpl6xZPQ25e6dMzB8qse/7F2GTZ6X/slIU3jrpupTdxvjY1TI
ERRB6QJCFtmDubvf+4pmp02IU7pZuf2h2Lz7RZP5g2AD2c13PrihqTctFpy6
ji4iytN48rwbEr8spSQdUXsZIqvzMu1/TqEBqpPLNIvoo9TAriVtzHeFoQf6
o8Dq6s0qvFrwTOXmFS8AtqBS9fhSC3YNUByrXjPxIT/YkQDwtEjKlFJD3o3S
GqDMwFUjvPjhTww7h1MvXYwCTPZIXDcW3OdsilHQwX8RToO9qc4+xEmTvpLw
fPhlT8Npv4CipTfhBgh0Tud8MgNa9L+bPoFoKyaJsroC8fk3rVp2zofTQpzQ
2DRaV9dGSkfuzJyuiO81Mfm2GXYxBCf2y4e3E3jHKvQhLCXWj6aQ6NZbx5un
aOByZ/RKgUrjEk+JyWGMzVTYDpacX42HETKa+nHX4vCIkz8yFpFtThVkRBKw
oDipSMTIaa0SVHUSJ1GyB5YK9dKdFBOKh8+SBeuEO0mCTsGUl2c+uWz7HmKi
rp77GTVrd5dZ8IpsVa3qgoQ45kvbrReptImQY/XXPHBnQYZsMLu+a3T3/VMM
zw1mB+NFv7V5Qf08oj0GdvtGzEyN7lAWbs0AyOidm5PDu2+qem0w1oZ6td9g
QndHf2WvZWjfPzCiTxfWQX7xMYowbT/ckmQtz9bdaz5RWK1ONv7ofZRiDkKl
AKzAtqoVBk4XdF7jrhG3ozVNgaEiTyv11aK5YU9l/JFTY2nvidIHHTOKZUCR
fDCyQdoCMISBe6Y7ABJNJGSourbM66FM7fzUOEax+14IrOHAh8v2XyLxXBqx
HRrXjwIom9CbrDsSiGNhPttm08oTLRS0uAFwM0flnC9TjX0RRMzcDHGWa2G7
krvYOh1Cl/CaCsmION+8xOMNttBmAeEmr8l3A93tSqiJyQ7VSHPp3h7bvADG
HEz45XdchR4tFT0IxB3FlkeZNHGmbsW08k+FR1C/NxiEgPGo1BTvV5MZ9o14
f1U8e6gl9VeDHzSPZP1qIj31YwmJIszn2Nbfcn5FedhwuSkl2oXkuf3ZC1HK
+cMPHoeNrTVH77ETXl66uLlg3GibrWGk27jmZ5fC1gYsnsryYsQpHsyx+sVz
9yv8NyJx3Xv5TtLGhrXHw9WUa5vuys70z5aoBOXRSBal5uxU6VwOG/qIEvIL
3Xkz+oEDAS5HyH87g/w2TMuZgON8MDJJmzCZhVEwhQfeGetQBGifWl6gzZBj
vBoHcZh0R3e7jz6u5cgKu0jMC0F8vJonya4fvCnjls2v8PHB/OOXL+ia9zbf
xCxpuswrT1Tz3S6zGPTAjM9+GaaaIh9tp9q0eO9MOtEmpiZnivjHrO/CL3LF
8SiDCRGwUhR7cwIchkpIE+VxgaEM6B0J6HvDP25jm319K/L6K6gYp00dQCso
im8ED9zCRMZwnduVOLZIkkoliN3c5Mzi3mRrpkrI+81PyKt9889Ko+zp4CrX
qA6Kpi/ce4dZRPMemsxj45p+s2d2S6/jAM9ix6m3NPYGso8luuELgQZmpqHD
Ma0bwKNOftLH4Hsj6sdszMSievkzVincftbu53VTDxxJwDefEUuIOALP5sGx
ivUTgoA90sdX5j1dSpQNCKwC9Zfjd9TSOSLeUVVSxMlq67rFcJ7DXagIclmv
i0SJHfv/A68QtMQxRwBpHl4/Qbe87R1QrpRtg4r9sNB9TZ7WaHO/I2UlWwSS
UzMKQk8jTXlkM0ADO5qWJg6+h6U78LBWlcJDgeE7QoTcx+CtchkVt2a+6Tk+
p4WbDuutUDbYabFcKNFhVGpH+Eqd93etZvqRf31lhjzBWnb95GZV5kVrSpNB
qAwZxhR2D5relhWyMWWF03c0nwNrr+gR7DWcw9g0U6O/PchBtVMgg4GJwXNN
cad1SrLITLn7tzh1tgZGp7UYNt/kfKsrlJ/wXh2zWpeC2CSxg+4O/+kTDdXJ
KKcNPgz1oDx3TdummhLTOBIP3z+O+m5Iv2FpHlo87hbw3KcOAtjW4SeljYHH
UbCyXguo+E5pAUONOIdL/F/475P1OXaWRbH12s+KM22XmKgGNFkGM2ceXJ/+
udMXiio+faui/qLv/LNJLuAi/wlxraiZybXRecgmlybg9SjVe6SIiqoC1fbl
t6tp2pssnebMctlU0Z8dtb2P7APwKtcBvBqm3XYLMuTGCaynV1S2cPof40oq
N1cLdcWvUnlSvwGibmXHV5Jf5D3WbQF9KHDktqPrDQcIpugA3vzJyO/KQ5NZ
nNUmsZJ2nVyORnzeIbkGN3iTRa48r1QSYZlB4MDhlq++u2iyqvMu/4xsUMCV
l1CoZhyPB9e23o9R/dIwaHvTAvuifCBJy5xi5x9NJE70eJbmPf6sXla52g6T
jzWSpYhOEaqKMzENYJqE/3d4B5tDBp28nwDinVyaFDOqH4OU4BR75g8P6Go0
4fsL+3QuUbabtkUQ5SrYsj2LDqpkoSZDuWJc7uYtGBtqA/NflME6WnkbJioR
XRww59ik7hBOLTpf5W0ngWRWv18ujsPQZV0YttaqYaClcVmlSt1pzT83/aZK
BZCO9WAr5pXa9p3sBmF9fKH9/ZXPpI5U29F6keuV+XUlhHUQoy/5jEArf7Ol
wigcslkoOZgjJpDRa7SUiCw43KJUjvMvjDlrFIXSQPAmp/Z/D5TlrrSuGxSF
YbDguZgc3nkPHC9YwBtCuV/ZRsqCq1AEyaUBtthI96FC+j3oY3aZ70W1vLE6
3SVeHJjPgI5QivX3J9xI4MlY1mTijqBYqNyltlxvoEp3s2TNJXNYdD+A+CAi
7UcKolN8irNonB8Oz79+BLLg7o0j1SlSId5PV8DH8E8chPbWyrClLxoc/bUt
7rUkJ2/avoUlyFxHR9xiZqlGbeQRSUC2ROb2b449Tdk9uJ6LMtVcetozN+n2
o/yrNupNatF7iHDTlACAirEhZ1esDNTi5dFBOeoJa9i21atcagx76YhmOQLR
AjVPt+ec1d0T412FHd9kL1DDCmZlMUp3NufvylU9/h7J65OF+p8gKzfVYvxM
kjJ+JqqeVhnZv5dZtDiAlhi2FPlNVlfxR61d6jQyO7HtNqBj2oJ+JBpar/0E
0ZKr2NUKoztRt7coHmbL512pyBOBSkHKeg42MLpTMbixIYxzdbutybVWFxkP
iiHYESr/S5fv5mVemLvy703JTMCnmAQJ/Ajco6Pkmv4enNTM30QywVzfreo9
BmhXoH8Yez3UZwiGLeealxeP5QBjBnA7KC+MLr1aUXU6b/rRD+R6xZYIF4nu
qIf3ggtB72Xulir5/D1vizCdPh8bB7XDE4NR+2NyiEBZm/8jZWAbRT0DCqNA
fMxJCDeQlTfarIZJIslz+oT2KRgphaSU/n6eDXrfZsxP7eMN+Q/o7Tm1QMBG
uceqozhO+5s1cfMgcYy4lDYSwCDoTOTHTdn5kn4SoPL0ChBezXsWKcJjYsEv
1B+1eoGS1MDgDLoNKr0P4FjWbZaWMg1tJzUmyno6aaz70sn633qB+eDjvGhU
BA8UO0/G2H5UbPEj/dArYmfUbjEpSr3a2c4XQCetuvqbpUrEQkfuiTrW9tZZ
9Txz63HlBePd2H9+b7uqYr+JyYpOkTaJFE2uAk4CDV0Z1wypyLs+6epEVos1
rxIjLSufcVBJ+2Jff7Glv8263X2Sk22ErMgaSp21qiR4BJLnIfDKHEuN1jlw
ng4N7KyH6Rs+XVYv33IFNujuVF6Rzw3SqJpLF+MT/gaSd7avPqbUp4yT6OLX
epY2bDIv2xp295hFx16rOdsmaSs0IPYmgNJeAws8PGdD26OzE+PxvbalMRd9
a2Z/Jw0xa9NUQmOYNGnT59gMSSCnv+LaAbsITM+mg416fEpeBjAMsQ3ocvgr
6eRRNasT6j8xqn90kTzzEgT8Qo08iaCRcnhC1qU2Awvqqts5cPTUeOxY0b8B
Mz0bf19uQZ+5Bz/ABomzmZesB0w1pLqEgg2d5a/dfZy8oK9SOzvikLmoBwS0
a9SpUFjubq/Hn017vrFtpNVU7mQG8P1hZJ0f+oaPIOok2fO0SXt03ZijF03z
yYCv7nlMR9RMYgXL17FtSg5Ra0x+yWEHd3+Xb6rhK7ZHfj3vcGNsdxW2n7Sg
BOQedO0HH+LpFsWyzIW5cfklPgWd2AB1Le9ofXWJjwpAXa2VBfd5sLDW8Ym2
4cEXgI0iYz+piKEtP+FD6pWx1m88uViTfLcH/0Hu1CBF3c+km2rky+YxxcYU
dg3DWU/803U4jrAwjxqvGVevlppO2GMUvwjzojkD+QJL+riGOCdcqXh6esy2
ZzoxdHd05Mi4L0QymDnW4d0apjEelxvZe4D5UysTmnNoGAVe3fNzSKwM69Uo
q1zmxkSoDUZq6JzN4PXYwYOCVQQpAEMJQdSMHxqPghmH1acrydbz6yNzoA76
Fy2AkqAR4hCcciLyfC+DkbizXegZn8SZPN1wSJQJWzwZbWFvCO4IZ8GpVEq2
+g2vElCrBzq58iWFia9Us4gA6YtMqNTg6Pxo+biElRq5vATJy+R7o0IeRQys
kmwc0O+v5WiXEDAtoNRdnxVJIMhRplApi6H/9DOcVDrEQNrNSFcSg/XNmBy3
kNc5pLvOkUDyCUg2gPmC4XYlvIQFNuyFYdfgqCcML2iH3xRTtWoF6KUA5hDT
iAs1h40ejQMVXiGvIQcVM53gpTl7IjKG2AJJFQTTKLoyE+l2cfk5ITpbIIsm
Gg5CmF0OjvjSVUMGhh2s8THdcRtNdbPTG7TaQcBDFh2MbGJjJw34CswZBdJj
b07EbRe/Wmh7NuYCQ81Ly9wXW6fAgg+kaA/OSQimkCbkCOY6x9E2Yln4o+ht
aTfS48lOTZf8QxPzz8H1V+s0KXeD11ha4av/sqIUC6sScLh8ynmU5iFctFJn
qKmCM7TQrAI4lI3hBI+77BqoY8eeLHmF6WhdPCP3KGKWe6ivzcefkR6OSOm4
/q+KAnAatkuC0a21JmCaTXfLr+P5HABwvbOLtPMaQ9MHyCrHOv7xm0d/nnmE
HAHHMSJTCpI/8/YEJDzaKJF8BQDkRa4dm1YYBh5RSmRzY04rkGoFE6eBBeT5
3/09EjHOHsviB6+A5lrlTmq7K7HFqdykJsc1Nb2UBjFxUaQ/Lsdarhb26dlj
EAQglykoQz22uxMRbJUejTSm8qXUw+TwZOqZMNn49W+hn1dFdpecqlJrM/uS
+tKsno7h/S1c+xWvY2br2pD8k2UgTHd5w6rtvdaKfUkS3uCc6dnFegxzs70k
qOsz/mXpcbRUhMxcG9D533tfXHsBmiY2BWH6SL99iP66852g1U41fX9KD3GP
Fnu594a+F0dGcwWzJxBuRh9u3YOKNwciU92OWlhIV9/9epPXVeZ9lQC2eQgQ
p0BilCbhj1iaGkTKyaVoZFoKfl4PsIFUfY6YlYHYhY4dARnSBJlo/5U2NePO
2t1Ytmkqwi+KBMfPTVDNmIKElku8/3Z01ci/rqko3Qcuh8Bcjo1TioeUKq++
0zNVBU/wJ4ETTHf/9BLHnN3+sl4aq0QGu4XrHpRaTVnECx4p5gf5OGWZZHb5
Mc3m/8Sluj16SlVyxqyx++iDmlJwMVqdr3s3WDdndXd81MrSmz7z0bIc/97X
V9JpuaJaZsgKN4v/WirsbMa/XgSmGwV5P7SV7Vm5lwKHhAwZUxBquiuXGghG
muYziknnGyVDYufN8ra8n5pXldu5+Fy5r6zxRovn2eimnm5j2AGDUcJTxdum
BDTDAmjs4E3Gx7YEtjP3HFuVxfXRfed0ZfiRK+3rNSFFrI5FheRn7kmjAjxZ
eVyjnZysaF/rr3yFxg2B6/44/fKCDrsZN9FYHT4MUZCfHHq8dIT+pkUoF5G2
s9O7e6fEMn+NsL2i3hyCrvK2bLVljtoIuhYFUeh9fLYDK+hbfw0ZwdG/jS4P
jka0kN4Su0D9G41o7ky5m1MIKqq6XmtiYWV0B7niBmxqSsHLJpfpYsINNczx
TBInJitoXrPj/wvRbPilqD1TUOGUNL7ed9bZkp278G/X+63t7lXRBaSjoGVU
LHZWnQoFRSKKWi8GE0atD7TFbR4KtjasmzEl1qoozxUK4pwo9En/RQ3AJHze
h73yvbNn1YaKlzOzs0bNRoqTJDhQT17tMbg7YqCKLAtGHDlUL/TI31AM8lst
pmXC8cHdHiuJt5E7IuWViiDqAdb/c0utvaWPLtfApLi25aqtlKygIJIK6Wfu
Nc3rETyO7Neup9u2l+cnAU1NK9ksPgAD4lFxjtp/O/qpSyXW5gL3OhYuUS93
LYGVfkSen273KSo/6/ShAUhalBs5DllXcTQeQyYkYEjyYm5Gje61EQZ7uKU3
ce/DF7ZQTqlRvmvtfSTnl+flDqPOGvvs3Fj6/03jB6zjeNLOWU7ZDEuBWdYv
3CY3dnN5RWAPxMcxXUtaLOpFlXuMsJIdCIsEMcbjPXZ0SKJp+J9IhoJB7Duv
YmNQP2FZtrBIJ+pHRUYwN6WLc1kzQYCYeZPgwmhDazsL34HySizTaDoeb/fW
Md8XCH5VBmsZAsSlTdXZR/FxBmZv+qWICCq5CuqUWtOrR5SKcauDYl7HD6pq
CZ2BbNwP+a447VRnIVolNs9yy/pQ24IrjqVnTQ6riGz6YkmNJlgxcH/EC4DH
2MZDm+9zWIg8+HgQxbt/gPeZTD9x5sDDv9pzJIzfjNLPw/Bevr7fQPYNlugH
lwrueQo0tzNMpUt83uFjiK6uJkaIU9J3XOvktDVH/T/PF4WAzIt6sU+vase2
SnobubM/cNgM+VzXZsGyl7H6j07DZlTIihRPFsrREN8bgjz6trlVzct9pOcy
1VoUv/saPgKKufTtXNFsVpRhVwUssaJHI1o+Vl9tzMvNu1FUPTnzzXebZQrJ
BwBUzJ4AkQCp3QhmUg7zR0kjm3s4sVUjQ2HmCg32Vk3GoVQqMhxiUYl0YxEZ
yUI7yUVB6CTpqY3rPjmEnMUT6w8QB7RcwEzLzTp1e6WS6UrtDb+CHSlR71D5
SLuw+CTiq8O6ZV5lpexZn38ZOHxv4TdbMWzCpKzDyq3Jh7jyfLRynKL+jA/T
4mwPyd7KY9eU7h3nGZSWD1F+o5WHtGAzE2adaiy26CcC0hhnWYGrNtn+UIfD
DKoUAZ9M/DLNPaoRhvwHFiNsirBRuBivZW5Jai2pQ8r5A4nvmb/TnOgrWf8i
qIIqNsHFMe8/sZkLOI5j7zSeHb8BN59/BuLbafTw2FUfarbvhsQS6RLZalpr
tP7ndacLXU7VkazcxTDGVTpZnZRJCSIgciLDJ15Fgl7N/5LH8oDiFHpqG/KB
QVQXCdO2/u1w2LNn4D9pfJATNrQCHQrUOW358Sael2cvwefRARTeeF87jpGp
5tXUXa62RXLWy1lxcTIvrrZVZ2zOo679kvuVweA9w9B73ik9weEa/qRVO4FN
ZyxC5znH3Whm3mCxVDSLyYEgxeEOoqYKGQ4VtKhTosxAlkDhr7pdu97v28WN
LoRY+2NtEkxhVokeDMqJ2z7DO/+q1umu8FFHcuN+kAEwHlVxH7DUt2qGQUmG
akr43Xpn6yfoL8bYuA+pD/Wo1S6lcO0j5yj9wNmRGXREh2J1deKqG1LfIJ3i
6D1xTjDKEK707f10NgJ+Ri2uHif1t1/CIuGppBXGv9N4LH9Dkp+oxPoaDZcC
Bwy0GmGwKaKFp/KZKqNvvsv0qwMGsnMCvyL22TPaWEp8Jt22GlKFtR3bvPFK
3dZsb/529P/jsEToygxEULhlI1qdGjTITlWM/CgtPqNy6zwVGil9EKMRqS+I
vt82a6OTeyIK8noDfPrVihZ1unLF44cBCBcpRddQpMd9Vpkz2b2PSvMDpdjt
yYav6JYVp6C4YQSPbqTo5hVEgAkvo3jP2Fgea7bHr+KAWnmzdnARsBbVrw01
SwS5c02Tgk2ITuruLI/7teMqVRwlutjPvYeUjRyNPCeGGBdxPpwfYwigf4qq
z5DVNxeKXdtIjETfeHRS3aUA3DzAOhZTfRQNOk4DCVJpPrgd8aYwxZ/gkBfM
fahvhhXz+bqPqDUwZnK/k7aPWPVr+nBmeXKjpF2XqjwH+DyRHMMaGitaCGMv
NnxbkQ0/J8ql4HOcfyuoURLbWuchRMMd5fS+j0S+mzNURvkIFGa6kM8ItMas
tJHrQiaotJg/VyBkdMMaIlL9sQryGkCj8/WfqEUQBWaJXdHXu6eGAwziFbxF
FRfe2IDxesiLmJqpUkoJPFDqumdvow1mRfwqtRJ2rZTA+DcrfbbQi9W8f6Er
az0JN+1m02g5sSIRZLdDh6O/+3362Qqg19cq/4BHCIqEKVK4tSkf7cUekDng
MNDeFsjjcNGqYw1NOXx6BRH/lznulH8HRHfxvJx5pL8Gze25vt0UTUiM1kLF
NUVqoTZ8zDgJYyQP/Npla9/AR+cQs+die99/OnBbfwoHiZpDRk018TJfTbcr
SHhSgB3vdlgdJA2DUKxW1GYFc6UQ52mXy4nao9HEm00oj0kVpK1mNh4nARbH
rlm8L7SzCVIR35hzrGn1Kwd9ZCKa4jX0YS9F3BaJvE5JvIaNTjHVLmnM9lyP
rc8qN+yWJMZPNKogQyUfzU+G7mCl0N672JJ4H/LRp0OQiklSrShzSP5T6UYa
hCEnQiYokQc3SMtpDrX+Dv8oW4xEH5uZqpT6W83R0v/9s0b/UovwhkRoWIak
k5QPAOxwPg8VWr9CQmEDQdlW1Wtr+VYRn6g5lV/gtPFNiD4eRdq08f6ABDxE
TtMLinLhmfvnaAwR+zIHSBikTnlsMpm2nctH3HLRt4atvy4EMIqeImYnDlmy
L4BNvn8KD07kbewiSUpxBseYzCPlEZ8oVgekSdDmf6Z9tNmgocBpMOw/g4RA
Q1+JphS6mxBGGJXQxiBcAbDX8kcT0v9tMZ7NjVhfCA0JRaYekJPn1QbYZpDu
wFuYPyySTMVeLmZU1v9zOx6U3TVeUDhwuhY7/nNoDZ4Uz+34rQoUyZF3YVrW
zgRVBpN3w5sSRKL1GNJy3tEnDRFhR8C6UlT1tYAGXMtSiahtABGXE6H/s4+o
L4/92K1ziFmZzMiOHKVu8dV4qrt0PmwCdUo8X3yCLUtlWfEf5QtxnEe8kLTl
nvxHzErzX+OwYP/qPFwiDpPkT9F8yy66kVgEHl/DpEi1Qyiui5+v+bA9n5WC
b8iBI7IIPcFCtmGZbq5LZLAJ8NAnB+lUWCg8Rf4Ilk3jA7C6x11e24ZIkpiG
XUunMnWB80w5vcv4KthPIwGeOqHtzSgsx65wK5q/18vart9AkhSHrW1bLzy6
dL+sP83JwGvAyoqzUvBfYxPNKp0Nc0pTuJzg0lHdrl8oJKVeHbqo7ZrEK1bt
+Pg1u0gyXUxESqosi19yFKKU2f1Wmr9YytpvLYZOab5WboZBNtZr7lKrIM1Q
olfYOCILLWj+p//5kA4AwuVeg/tPC5qpfSaJlUpRUtGQPja65nvc4/mSjtok
HJuZCu6aWlhMD4w1lmYzD01oSp1WQ5dW/d9GJBCX5Nlry31kS4rlcmqEQ2dz
ZIPgmhJm0Fdeo9keW+dDoJiKKgx/FtjRaD8fvqzj9ACxqP7mRv06wK/jcYNy
4ZLpI17MDhuo29u7DHYrYSUUN8tojMUAaSTlAI22CdRT0phuC5RwR2jwi5Um
Ox/+vq+N9BleYQFw/2IqeL2eBX2hMyBNiPrbBiKPTlH1YtJe7vcZnzH4rgSY
6uIUmoMzwAod18c218asv2yQN6r1zGZOdH5YUGKGqpJV+Ri177/Rq82hglwe
yDI3ejW61cHfFMOPbVmOcOKxBt862GmrilMP32dkc0AabaPBZSlFPjaKdZxZ
18bcDUclApG4fJjD8y4OjLZWjnkmdCAcSqJ0Cu0mkPgXsODHxt5FPAKOkxa3
l4F4iDl4fhNmOIetFlWs4Ng+MFTZ4kmhvt5rgD3FQlu3bdG6g8pE0cxSwu9K
pYLd5zuLhYcBAIa5enDGHUk6LmJ+qAVXTwMXP32YWYR/P6e0FpN81mC1qAXY
+8sBBF5a4vWfE2xNpRZf+bJ8NoC2u2a+76dqQ4xrk94Clhup60YpvxvYQ0Mt
7CD7kbhJH2EubUdNXohzlBw692hK5BV8y0UKOjBeXqE4z9wbPrJW4N4dDtZt
1nnGEX2b/xyvNLYbJ5ns8d2/I139AoC0Ai9TGdVqef9lKDksGiLYPby3hQ35
7ShzvVcnEEsMoZdCVeY5S3wKepu3jWqcuxaApaokegA62mQVOz5W0sl+BmT/
UyT1Nsax6cau5nnfmQJGCdv841XqRZL2ko3+mxKhUBVV7MktxK3dkn7BHZ+s
IuEhNyrNZbh4jIXLfVPBAyWzoemRdcwDugV9lU1E6jmtPx08eJUauw1822LO
qkVcWdX580/lPYs7BCBstza1Q2OXVWuChoVbp3ZyAeaS83KhIt7RJcA2Pd3x
RT6awSC7V3jzXZ9XGT2Sw0tLXDqvgRX22pigDKYb0b3xt/6VSYLDiYvQ7wU6
wto2YDNs596G6hT/oMzC9QJXeYw1ydOAyUyqkklxQrzGAvZZECWUk0dHYp1h
stvQ/WShk2BgxRvnIkd9YO6YsFLp3Qr6fJ8MKd0zuBvFDspo2u1WnEt6vOYA
v9G1jI4DZMi10eRDdaPoeiXR3QXwMY3IFr5cxk4m+zwPKL4/AJlYc5zOa91X
B/w4TKVh5JrDittQVN4xx3UxkV0hskuJJ0S/wCaMWMoLiMjK0J4FKh33ZeES
zNjFTAxjPgBrvYkIfcHUpp9uhiWmcbIxfBCWs34K3XJy+ysHAxabB0vxXVrd
O2itdUHM/FLdCgvL3Q+Qb5tibQr+tC1SX+D7M8H70vJXpAV+xm7x134wg1Dr
Qxym1fg1uH0a7nJjhcuITBWJmFSzOlfhqCPgPbdJr3jIEkytDRnvARksFH0a
xyX8VRxbOWk8fquXupyUb27OKV7KRYue1Ce/5vf51HG5u8/1DyuKjiYslTeQ
YtT+NSkd3FD1glEzVvlWmrda9MU+TXML0RGTSCjbUxoP98lniP2F0n3yx/w6
og9vo2mwri4fHt4icd6XgcLn7EdPQUbCkQ19IG/3fSD306Ejx3Eh1e7NyHjf
oHjkP24gxnj5YkM8/g28lD89cSgXutQg/KdJZ/nYaciRjRpViKj1zU0Y1Gh4
/uLwQZMiF3A2tZYOLt7Pl3SDU0pfsHcEFF84h6itLTaP6VjoZMQPew6qekH8
INqHhU9lJT0iFFt2nAcbAurY+Z9En5+nLANAej06T8KyajBPTYi17L359DHS
svtgzlp135LYZRs5sCuCtM7SvFBXRfYB1HBCzjkAmpBRf5fW/yzQ27x/rXC+
jcy1AI3JhvbwbW2PYE8yVvBYR/FRyFmcuNpjyGYeJjZQdQoo/ORxtNz9JYIS
h15SMir3hOCYMeW9cG9my1dwzQRyjpz4PXbUMEDHLb/1NKj/BPVFiMAekJ3H
VwLKtuJbF+k5A5UUJRuaOev6UeKremThGjFj1KP3GW1E8R59pgEFyOLRRbS1
f/dckipCHrgFm18UgMC0zQ8Hgvgj/SHCnlyWpxa5vxO9wsvhN5uvTuyueIVX
bzfkjl7diWQeRDakcpSV07U1IPGtM56pilnMRNkrZ3fCgF/lkObZIHI6eYJf
XR3poV3eyNVGH4OF8eBLoh3BQ9uWE74UFBSqAOVay3NhSFB0454FLCtOgBhP
ZUVyjFUTpPsmg3aX5tXt2z1uc77daVbtZW+WJ+3I3Q7o6W0CG+yk3Qaq+e1X
JsQoXwjXf/2MOYnP0qjvrMqJajnsAX0hCLUWdwcjxSoh9BGzf/Y8bWi8Bkuw
86N+YB4ojmSnMNidLEjeTevaBPrHl9myUDq7aWUsd8i5U2g0++krAfNaXWu7
AwByJzri6IOvAQAUIrCa1ukkVJrfsjPIV7TVmpFuPZRpQddV4hxD7bfYnZsp
G7zQvMmLq/uksAjO+XfZP12NLeYMYBWJV60NlxhahPE2oYMlB+ZK6HGMOebP
cJMB0OIAzh05t/v9NYnZt1w2k61o6o6afvP5ZligO5auIdm00GyyQMDKvY9L
kK9zdKiJoxBC3QkuFQi/nOw8WpNlIe9Vn14dg205AkN7fmeh86yrAje3k19H
/c4VZ0PN+k8Ui/6I/XYPgo0ZHwpIiiFCOYHkhQ0SZBmo5DDLLlaIOtL3UKYj
UvypG6LWQpwcxEUG2rrDjDIzYz9V3Fcbk1dSKxvD7a3wjHxIamX/rQQSxbwr
Qx0A5QomK0B6vODtbMA2eF/br1qVYlv6eT3H+PZujJ9opco+SM3QRuxYM8ks
gd7gvwKs1oe5tru3KqL49aurLHo29X1crRVapD63mMkdwH1gLDK3DRHcukRO
2+TyJrJnEe22itm4Xf7xfHhX6nnqM3+MFJMQaHmkRrivjoDCYP3NKcNnudw/
yllHcFWufrCs/cOQcAzgmtY/NMV8+1qkPtsU/86dewWENbZ6IyaH/4X8N6zz
0jb/JcgWT6gjq8GxB+8VO1XcYQqyEW4KD/h3Th81jF0fa426Xh4c+P2DC+B8
IVaUZZd6ObtQYMgVTLo2VLGnva9ksDArfJZFg8DSx35XL1PaPm/1YSsT1lka
NRr5jeo1++oEB+Olv0iBUEZUJsX+Ywl9sPQpdN2IdFPIighH13YuF/NaGZCo
Y8EaTgUosfXHFARmACgDdIhGdpj58UeGc2YJoyTWommMhiKzLUtUXGt222RU
Qj8uDe5piWe+CNTgSe3TE4fzyiW/xPSt+L6HEZfJeU6pGdHSoxT1jUKIsr/V
LaLFLX4XGqXD/hY9uSF/oNDbLfIT3f5VPe6HRnjEgBvEK8IPgYn3WjStMzPg
E4vMB8GG5XF/gUHSOhOXNag4mWSJKttDRIZdJRMXgrX19rJ7JJJFqiC40G1R
W4fl/yjEzE7FLdgrDfhHqlkUFyb1NqfzxQ+/wmGm+YuCJ3hEVzUMQ5zm794j
D/LlncRrKMAy8nE8VwKSIT0gUd2T9Fj+pb2H+/CQOmWkQkqtYufH50imwcOd
OwLfCMp65egM22DkgEAegs6F3v4CQJ/M9PYkRF2D2E0K+ifAhLG+1PPGUajS
kNxm++iJeRxuzqesKVH07L/9C5wGugwzFHNIFMkQY7Cmctt3DpAlctmiSCRo
7mubWig8BL2qsQeHbLfQXKkuSvQ/O+flo80mp42cp4w+B0Sn1C/Rz03CFHMg
4/ElMpc6morJ+TRVH5LjAzuBKlkcLzLDYRVRMqsKm8WMy7Sy9QSQIFVgQ1Qb
OJzx9I0CRXRW/NhIzeCklDkQKFgRvcou2fcsLPDrTnKJuwPkwwNu7bLtjFO1
tc5NJzA9umuDppdJCyscWZQLdtApZeuVDm7xvIfcxv5Q2h1YqMCPZusTs04u
cptJ93N/ew/KcT/04lDXM78a9aXxKNmRz15uHk9vWRRn6Qm7EXlO8JJwzP49
twvc66pANFpeqZir43hlkvurcf7vZedUYzPZuOI9zQG1j+1Ne/ASysCT3yyh
iimiM4c4/dZRnB2YyVWmhkLLtyu8Bopg5ZQVHpmNPRUADqLpDD9sfSoowPnW
BNmjunkMAyRQZCZn/H85uZYhvSdDy4XOkygdXp+ciynYz+21eUu8XABYsugp
h5/Uifeiz9buo6eGHEhQoHpVmc/HV6Z8zCtMOsEuLYLYbqD64X9PZZI3KXg9
7JwRpEIqwp0ERo4u2VhPog0y5XRTlYVP+qHf/6mYOfWj5WlCHzYn9uX/tqop
/yijevVvGPebQiEGTWWyMTdkQ7PaknXOC4tZDPiCIBsXz8CUPsjFKwq8Y1/K
Yo104DvdJBQaNBzlD9iZlTJna/OTH5+eri/eH7cxSTbQ9MgPepiGfB5Tuuvh
OWjYX/tIcziFJ1rMKlmMiUfD4s/IKCPekH4T7/A20yGpr3VQTTGwRE5ZBtnq
8JwmAB9F1GXRtofoFmnvu9NpOVpmIYaxb4Zs5Yo7AcOkcMzSbZ1/PLX49oeu
xKf6Pni2AzATNM/l9IiC1EuG21L5zR/QKf6d9KySzxc1GSpp/5jeA8GsE0OW
ZcyMJhyZVC10ytPpOesZq56d+08Xj9tSnqPYlDS8gMx8MtlHVXVHVq3DGQ5L
XWO29PdyjzSztCXr45oFLnECTDtO0pxMM0cEY0/o3qraGZJE5qCLveXUp79C
qi0X/TrMmL7zUJbH6fUXT1RAxn4jc7TBlmPzKR9PdWu+dT0ohdTNUnIq41Z5
YC5fG3lWiXCIWgF570CXn4if80vtUtwbpfcGZd/bb4VipAzwnTrvS8mlHyfc
+AAA1QsVOPMlhNoo1Wiql8vxR2biLBnAeyaP2tH6WJXvb56epM08v7qeGqZw
WeViOAmO5fefCVccssw6U7/WnpePysfNYErwKTY+42CM3YwytkmOKyoSCU5J
E7/OcAqQQffrINHiQMezVtOp04LQD0KfZXVmF7IdrKUTJRD1x+fl53KUEsJl
tvM1g4rBnxkvknMsnFLUR2wMeQM9R7vkPCj+jOAnZ86O0KALrAsPdA9uVBRk
4pmzDymXS43d+qtZKeI4//iKCYqEotRJtYF4qRHDXshRqFkf6q2MXAi5vPCv
1MMwduz+cRyly5YJstxgwH4cvvPPAJzpp1h+40UBAEh/TXYMR8zv2OP7SGvP
LbYRvMxroIQkWVkNf0Eb5jQ9dtMOXKENACwB+ufY20pbNe2w934NdkdNWuuq
ypjdFexbFwS9Os/whnKgThscFYgtcAJ4Ft0l8Z017WWaLZNpN7m93Uti9aY8
Sgvsf2i0NcQZDcu/GpiEPdzjPDRwrsavdsIeL4RimAJ1Y2eDSPUGGI+GWtFp
Ma3Lsm5lVDgJDNXQqOnkmKb9xmkiylRVBqAvcB2BGBamH/G9KHhQxxhCr8rB
RWGJhD6wFMlJrx/hbh7iKeE+9bQ/fVvcUf0w0ewyTsuP0r9YEokSRhTkF8kB
uIASY3bazNHkSY5PcxuckqcREIDCCEHzdALaXF3iEdrz/VYBPXcB+Bs0AKJM
LE6yn5MfC+TZAJB/s5kqnF7VmlZCjDYlrBhy6BE21tFSwq3wOJGbRj0O33Us
BvHvy1OdGQ+yLSIy9PeuYgH+jkGslhxTeT4tUnETmBtpk1HESU3mXgf/CrVV
+mkPByUCHgP7jHAUZI1x3gHYgUR5Kj9OTOmoetELgtNsjDkZgiBLw8cK5YRT
6EFdqrIRC61saFxj1wiBk91EFXuEeDS0KgHcRtuc4IMa9xPWe4/FAWz651fh
FA/O0AMSh0I2S8bU6tGWIBJakf+TjPZcKxobrgUpVcveukdPt7dC2vie0slh
e+NY7aYgmTtQ/Uj7uCorwjlNfzS7JpPvKBlkTwWfauzuNggcbzNYdidNEHAq
VcyFwYW+Xydny2Kh1L5KP2g2qIYNTIo8yga8rPaqKq9Y0mhjHGhXDuH+3WLh
yVG0BwLj22DC18f4nzSXKc0W4EilLBYq6EyyFTncoeI9dMCuOSDXvCEuML5X
LUK/5T2FC2Ty+N288Fkpr6cguipiP1RdHNItA4+PYcMD5YXsPlHfkdqaxZtZ
DdMHlUd5XkP2S+bao5PEnF6/gCxXWMOy4FbwDTupNmYYVB5AhgeycfDqOp36
rqv60rWUX5bawQDERD0Kg3yALTG4o1ry9M2CpR10uH8t76559taYV/YqJXm8
JIKqPndYt6emjeOCScutdC7rDffk3HWRBtYORd599ymxc2g6fZV2l9Iw9V9L
v/EbfnN9FEXSo81LqGYA/6Lu3hJmsJDoQr9kLkefMy3FthpUq1g9AfybA6NB
MhpK0hXqdfDCrgMYgxAcbQrpxstm+hAJaLnk9dymRDki+zgCueoTAKbDYHS0
2ArTcImvn27Ag+gOHQ5q+F/pw+CWVlpcNbuWOr2HMdhJlqPpm3E9LNVfd//r
Mg5xrXKg9Z+h5TgvlRYRBuxy+F2iu7HwJRNHHagj+s0lakgpDWAchoh7+yNC
1Dros7IGYNHxoOktPBxdXAf3vwFCnnPHm5ruHDP+vr+sF5znZ5RDWiaO37ZQ
FrV3wUuOWkaLLC4QNR0sF1wVajPxd9giOf1S2PANxvobgDxR12QEx9//7Gfi
fUInWjxq9l11Fi4u6Q1PiJrer5ixbKfH1RWIfFGaTXdtarGGXIhp0PKGwMxB
m1F7QsnTmCRzA6JXhDgtw1Hj5JVFeQi7Z0O1w2Z0ff4RsQxCnu9N4pdTeuK0
XhTGagh1lxxaSKJcrDJQfpiLbp+roCY8nTeodSRhVWgDuECEpMRHajjJ+tzF
svUFEybRgCLbj3YfbmuMmB2QrSoAzcJUDHJhECFbEjnWLVJbjXA6to+Be+i1
7Q9GTptNvOGqz+z4vSCgHfNxCkB2cT43S9/4Z4VZbrOHbuF+p6e8bB2sLChI
BOZwjwZ3YYK8/Z6ztLMvtb1myBTm0geOE36QiFxpC638aNVkcfyvbjzklEaj
D46mqIClw5nOyf6JjBD99wpHBvfJFHIolm7GA13M8mghKllaPxMv603F0cYo
Rrg3qdj4rDsd1zK70scS0ky3MTjXy6zfyf+aAY3MeyC4slJ9XegRgt3tshdi
TD5EFQ2iIjoyH9IDiDebNZmzaLU950vx6bK6fKKbsrt1kBPW/2rQAv61kA4J
jFjM4PmTXzHhQ7GlYqP7teMIWgVLwNHYnVbgS47LTzZp0R82N+IIt5jLVQJU
TZfHe0I1Q9KNDGb/ZWNpjMixUpe1n6WvfAwUpGRIWVxkQmo7PFVH2F8+7ML8
xjma+5IqJYF/P6HkNcK1S6Nh7dF9c8oEmNbcb8XDFZVYSM5q6Jfvbmrm3GK1
WPByhVacUyGQE4b/ed3ig1Ht9qiifgy27XbV8JJ6VH0lT4WyaAYXxIqJm4mi
DSg+Vks5vDFMwnyOqetry3b55Reytz7/b0eGhgtUmO9BF68+6rEiySukmniR
kHLchzHe7pyAeSy0bcglnMmhLELNUoYWQBrrsTzJSQylH6q7+xa/lby6DAeT
3KGD94H4aOaKYeyXV5fFH6UdSpoOIjWGwTXX4TBR6StQLxoEp90vOXF0uOHF
VMl0Gvx5zwDlHInNgiKnz/2ErACHLthflwwY9Wdojhi9NUIF3QVKY8Idtl4z
NOfTd77WTmXXbRm0LYupqveCwo+KFinJGLsvi8R02IOuugz32TsTMySeAuGp
2ezGLFwOGDUt65PL+jTJ5W/UJjQSWcOecmW/6fn6/ZmxLOA+2qX6SmjZyydC
YCx71mozZNnnaWEv81mctKBHagXWB7Js3hU4EXQqoPMajnFp77clR6ChALWh
XMlIRbYQoN0gQ0LTKsbjT5r9QB6tRIl8Ow3yDFSKScSrQ0zbJH/3TJBFQ0yu
H4Q9GGsDb7MetV2BauWqQ+lZZ4ZAUHrASHCNoAbCSt+s42GVKHh2703t/vnX
w/7iPfDzy3qBfxZqNTQVVopiisqghzoGnfxtRLzmGs8eEI82pBR9AoPtsd4U
ey3ka40pN+7MUiohTF9nFC3LmxEaeHB5nVeLchB1zgm8EkUbXYvHUM3jVGCa
CYUpwUfcs7csdMY3z4OzSKneGmkn+b/KBiYafN0zT0GKIu8xmab3F2AuKksR
qMpCe2mM/t+0pDM/KkWDUy1cIBB1DaTnNsayT4cCJqkYkiBvhTuo+10UnAtd
DOF0fJyOhfBDCVDLr/QBcM0N6WizSTubFe94CsJpVrvRQIbDRB2pViahZGfM
IRh67EEEV2Y7NI54DtT/8LYIarzLDaxFgIqA5D2HkL07AdZYHBdKSpH8YQMq
ep6b+76CrsKcbk4i6X5yqySEZUM5n/iFRPlgAAsbSYQ+ufXaU60yUh4AEnnR
77+EgRJJEU0zuxVc8W/GSkpq5FWIEXEYqPs69yPlRuBEB/7wwjxr45es2f5g
PoE20CvIiG5cKXaVvDb2kIuFprOSdl+za/PQN+mYCb7UI7Uuo3AQcdVve5ZK
mM33tHdRR9pJ6evTkq6P8cgbV8CArTUn7FsEYHBX6q7Mn4LS/For1lmfswBD
0OmQgyWEPxSwF2CN47R85MZnEL9xs1k7eR3AUul4TWJWfYEoFDMc6GyGQI3I
iTcBMBZoKzn0X14keg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "lK4MM9NDeLrdcSiRM+VIuNgpOLUAzWAt6nzBJ3Vw5tvBogzjtStM5gMJjD6PMmMyupOFzYouKIpJuOZh/11WnQBMmqEc6gvbtnHqfGmxFaxYyOv1rddc1B279ac1WEgUgi2BHG6DRj+tHk4+Vv2VvppW/Z9gUZ9e40aCxOYZZHwEVb/SJ8ximgD4Fihl81LOgt6U1JRoR0S/yAHMZXIkaoJ6FVEBkPAD3J3ew7MX9Exz4eTCaX2BwVKMD4Z/MOaDrtynzFnZbRi9WSvEhCh8oR9byir6kOnPh1zOy0xZulSiQN6SdFBsOGMZM4rR6Qk6MKYVndxL1CJfshzNQa7bFYG7qMnu87rjHNLp8ogSLlt6RTr4lQuPhZL3p8RmRQVkHfMXtetAdRnhIbU1D0d+4DN7GAZ+j6b4sjhJ1vp8Nz5D7Ndt/XRswEP+8IBj99EM7jgUeFr4Juk61F0vf+4TQaJaPzqY2n4trz6LX866fa1JoLMw/xivYkEMWrdp3nc+K45ICq4RBN4DMil+VnmMzPXyr5MFmD/p+J3YjBZhaCcSnwM/qC3zzflkSBmlE/gRHumCUe3leTghH1+SNe3CGHxBVSFJV1dJK9wuBG8NQlozfPOQVMjnS9Nb0usvhS8HGmBuwJ+LT7GL6O41VjtRuWYKTqX3g1LGgPCeUa5ERH2fXTGFAqxxzXWux6jaJmX05kdy+TUAWGS5LVsGLG8z20Qs7bepXliWgA+NmaO621vlTeny8HvCAqJkbaA/xbLKNeXsej1usF4ZjK/dyJJdsF3NF+rRJO/FHXmwm1o3jRRgLPVSCRplYYR+97tXZt/TxqK9KzLZnlEIhMqWRCoPezd1BPsgYMcFsA1vOXkacRf4Nr96sg+mOzif+0qn2i6/E4xZx3MswT8u4wOiX8whWnznZABPhKDXZLVjwDF6zFUttAyyGiPjxj5+czxTE+uygn2IYhHDktKJBmObnQX3JQ6nT9bkeX4DO9GgpB4WXBdkXFrIdkNTT7DJXVt+fVbp"
`endif