// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WGQ9KG7MFiE/ydjtBdYlCFNdEjeC0ZmSx9IUMV+G2bSrwQWi88dRkrRcD2rv
82cdgbRizhbiow3ak+d3lhQPuY7mmuik3D4d50aCT1ThQ9huGH6WwGi0oSpG
BHlafD/ERES+hSY3yxBBktzOwNBlVaJMadIFcvFvCNuY0F9CDZCLhadpIClh
dQX21Jh/+bc+F5Wrn5lrnv05xmVoeCpPAyFPuNLSMYNfdzVMF39H8BQLEqxB
FoV7ibM48y8FoIHiKwP9XALIgAHW5O6cOuQbDYwLzJ5CYbmXoRKU8kE7+Kc0
WT4MBPuCfblP2KROt5Gl2XeKMgxp8NS269URl1nhjg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iJRXF2/vSscLlrrJ1W55pRBFbjyzTnxM3nwdqigi4hvQwOFdZad2ir4avbMB
KrZys8fiYaJShibr6z58+NUj8htyUc8hlFXsIQXRQlYf5Mip2pRjrvebqRG2
h++Up6LWWmFVhYgiXIEL6eSeYiDg89NdLTDCwWyFdOQekh3aAQTKLem3dtTR
CLnZV5sN4+C+mmupgQohlhoRubUSwMS84ATW889TEbr7+SNWxHLpenSirRXL
MvkgY5ovzQZefNH+h4C1QwfYBS9bEzonv6GJdRHLARmfZ4vwmhkN1R9YPqFF
go6HqAHidA3vAGhf7YsWvvFqXu0Kgrli3sJ3TZhIAg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
j4NP4U/U0X+tYYqLs3MHyoMNE9bb+6HrY3DgDApcG6lK/GzP85gd+vf5zn0I
KgGpnaisy3d9k5seDALMFxlv5k4aPJsWu9qTBcLRg4KQhBehyyuWGo6Y1wMD
6O2HtAG41YiNt5eNXcJdeSnNcTDEwZ+IQOc08fovxkTWWmvF6xTZWnRPbkLE
DABVIEdfHOoGmuwHt2mwLH2Q+ZHuwvqRovbBoyo8qHoSwzRsgECLmY6/ETCW
8wgGEQ7RJnB2JGVluwg9ofnD6KV/MTDzu4Th9qPo3OHrJ5omtz7RJDUCmd7Q
KEmzuTX9EXFARtmBIf3n35feeodpFLeWA7yMnjE8XA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SJplbHb9yOBuwxjWhMhRF1UAkEgPPbZXC32LDoqxbZXa9xzyPTI/D2dyRbSU
T6EeB7ie9bFd/N1V7RgiCgBuD2Bi51SphosecKXY+6N+cIrXIw6M+ba+lL4m
oC7Gk3wjd1DL0m+O5qXdKOdzkZYKWENXtzAPjT+/g7dXLdEmsg9x2yrGOwfC
wqniDQEJlLCuXU5x3u713fiSzc9Y4OOMlov0ExkwpkfHl04LT1KVEXgXwOWX
aJe1j/wYsdRgRI+0H0/sSkCyEnXezpfm1pQ2/0Bq0RyQY3WtG0U6Bre9AUqw
I+V79DX4SAjs5EJ0pEkN+d8VsCc5xJWmH4CrlKl/Tg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tTNpFA/pCx8qcUVa3x97/103ivV+AhLYzIAqn09xokb1MPYhoFtV2S9H/99s
smXHUPezPWmHHiPMvhsMU+reFhbg+ESgPUczlOa/wCWZd7/BjWxTBPvuTlHB
mtmvHaeBnZVPK7Dzzp4POP07fTu7B2zl1Vsuok1fBVTRNdNZbu0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
KxC4KM46ysBhqHyV+KBCp9kdQnaZfQqwSmxkyYDConQMT4D1FbDntxml9YjO
/lQqFQCYiiXn/ilrdY8HXURP9bAOJo9CPKKLAnSLd12L8UWAQspGsc4Pnc1f
G6rzx/ZAO9LJm786esdGOI6gnx+pw99l/MakxoKG/DhPHFXQaTg4TwzLHMkc
Osg5AUTYq0GzB3jjGkv61VlRo9QKclWuMZw246vTpCjX9PMrPmXsTg0de389
DXe/melhbgD0IPt+dEc/iRWVuwAfsbYml/ngt9lOuu345GZ4BJOybGzyJLp6
ygu+0808I2nv+4FwgFNR6kJNe5WBLFgnMEdnAovLDAXtKWqTd3P83tVBSdqv
PEv+gA1o4iqjwRoIEoL26ACZf+9mcuTnWJfaOVqh1Q5QjJ1h8/cncUCkEShH
CObCqrdn+LoI1G8fT2eQFSN4t3DWptK77SiZUWqe1b679JVfz19juXV/RSzJ
CDn/Ve+zRC9mZdvAFLhyqoJyj4Y//n4N


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VbFiOTcUxW9b2wj3ccvubs16EpRZ2LaTdgJMNGWzPQj8fjnvpE9OIWnrE0kx
cS6Od9lHRvJgTZz6/MM1pwAjXpcr/Nk/Lt1Pg+IQvqgW3NkiEa5CoyzPwXXr
PQy0/aKQFxvmpUbn9/4QvIfKjN+ATZYTY/nq3dpezYxsB72jiQU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZC2g6RQ55vOs9vnm78iFfVkUbDatkakm4TDRmHnvaknPE+UZh+IBNNZtV8A6
yINKnugv3xyp82I65KCEgUDS0WcXoifM+ip54GAqqTrBb/j/Mc358eNlNYf0
uDM2e5/KLg5dexHg+psQKBUWbQbg+CTJEkbvMi30DXN7+SfwV4s=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 42224)
`pragma protect data_block
7BqGbadj7UUoeBfK031ZaCbsASTK1lildPMaMb81zrqBRYMR63vQpjWSCva6
KpQRnXICjfyBqUSh8PKAnXhyD7yKgTOaP40gjLLOe6+7rjVI3Twc8r0tDVGA
27L+bhE0ZMUbZIAQe6fwXC3TGEs/Qc3YRraN6iz1MLIeHMOJWRaalS76oFpR
yvkdvJp95QiX2FEZWrv22VbBAVLzidm+73SJaDfw7+ZJQdQZQjFEhp9Dlp7U
1TVAgO+80z2HOlyO7ZedtizbbItKCeAs0URyjD4cq5DCjv/ubr7V3zPW0R6A
Ycc25JtqUjFMHVwlcNTBEYMMgQ9PiyoVfSPlNvOhSVTxpPZx49VRpewx9e0p
pvIwSOCJ77w1sDl4saeE7kuFr7I7hqFAd2nnU/XN+Iyh3/Lz9SAKDjCONN1r
U46IC/5j61RK4OsB3ov5BmTRU/nTVzlQCefSgDjm+eIFOjTbAUstOZZNm4eY
KBsEDAfpTcPDC1gvdC1VBjSAsse00SU6gGlC3jX8ebBgKPgfgwRWZjW1ux5d
yFqDYSdtDgpX0k23gRMb/4yMhwqxS/37DaENZzf1G1GbVWeS4fQ7pu6nbH0u
KuFX9QLKp044QXNI/bkpWLEf5SNx0SG3KcerzWfBPGkgWKDQFUaaGqKFpDJf
vFqNKte7E8hKmxaJ7UnvBzTbewJmkBkXknc111nLHnIN7rLf4weAO3JsfLSx
su43neTWZ3lC3z0E2zbJaAn864kZtiGxNn9WrRYPKsR3ljDWjAnT80ZxDIg+
uu+7jKJtGas4H5pihUDCQUntlpVohQp58FBJEidLsJixqAQ4Yi668XcNp/oQ
FdaXWnI2+yDzLZQFwmvHHgVd29ucVuXoMklvRigfcbPXubu6Ycq7VvN4nl8r
PSya3l1s2ivZzZ2UxOoZO+zbe0RB7YDwNtxzdMr1tWQMxBjfmG4mGRSvyrJc
Y1vPIdu7EHaeEPxYNt271sPLJilcGj9KbqIk7uG7W6YSogmhgWYZjt8YxOTF
tBpXzurYv0g/+zBk1mLE+/2vvUZynwBn7d8ePTjDSJ3n7OHMZq21VSe0gJ+x
QoJpC00U9alNbv4W627dE/wXJ1bBmRbAQ+jjzcHh4oTPKwhH3w8yi+slgxng
WCMqLgWyvxpxpQ4TKTLlXjMsoOmmMPjWSH8MuQmYzUU10APrkYoNIQS4GvMf
WzUK9sWV8iL7JUcWSLqa+oB3GmPy5wUU+wXdmgfC062Gyp2NZdyE2cJJORsn
7LawJ54tmX3YT0qRSoB4O6jmUdmAWqNt3gIkkhfBjQRV2Su5BoQ+SgwGs/ii
aMV89X21sz/cRgjOxdJi2nw8rXcXDaU7RT527eJJjs7VTrBtWJGPKBqDNCYb
KDhcxz6JigY+20sjIfvhOHBZ+rb7ZtA7b19RbWUwslhKpDF80dPhSg0irVQa
jBsYaGZ5k1DAYDteAa5V4XfLHZQKb3/pwMBIMgP0xMog/qrzVU24u288/Qaw
Vu666wT0IupClITg9GPS+/xn9/OssuxZMQiEMSKPu2OEqYMh9twxg/bJqpNB
ZaOI/AKX57rvpISilFN+9mx2Zrbwy/yN1kPMF4RepwP31gOEOasu696IWIgU
Qmn9+lI6df27Udu9R6ejmqwD37VqoHKdXLi4SU69U3wOy90val5kBA1d/9V+
vHHDXFbp1RW+lBjQV6fsH68rra4Ih5/3GXL0v6Bk5bcz9RIpfqgH9e8dnIQz
j3Eb92B3JfBGMB+ZK36xXhh0z66IXGP1kKiPBEBe1lCxcLnWI5kKipN9nfJK
tFlIeHYdiTr3Sdu3XmniajQz+SLL+WR45ns0132PE03JIHLsxIFhGUQBSQGl
r0NLeoy9qfsJhW998iPt/4Q/ny5Wh6+Ju78Km4Xp1l6ttQJqG1A7ldB7/+Rz
J+Fx7NtmuR+86IELUref1IYL4IY6Iy9MK2stgseYPE/+QRWCeX5+EkqR02MQ
Jvk5zZ+8hsOkGCpXR7FSFch8gzuUDN4DCjh76S/OwzjHL/d5mlBSOkqN0Al+
LBId94B8IqOpp+TZFV6QoqrUPE5BwOmSqilRMXbUhT4SjMRfywpgwPxL7Srb
a2K3QVP1o2SkVMRM63XNOtuaeSSQVfvK0/RrE5tabr8eq9+/KAvaw3csRL1t
1rHe8HnUTxxIXKlmq9F3svALQoHC8MjEEsV0Tm4kGS9Dmpg449e95SlLZ33f
owsx47MkqjNEDupDTKM3IAEMX+7jJwCf54Or4kVuNRkomBEPiDVYQYE4lvBD
pY67NpWNIaMP3qjN6+qdnp6HSr7PlhiZVA/nYG+0NEmOvjvz+Oey3lXiELcL
R1tQDleCtR3depFa0oFLElo4zPM2BsGMWKCKCkxdkruCaYNPkHHBCRmXSjQr
FWoCNftEzqJk5dDTNTl3e4qTtEGm9I9rX9BCf69lLnRiZo3oveeb0BUx3Kw+
G7Q18o0A+XU9CmwiNgP6b67NnzAbXhWUp7yrVaCF4+S8ifgycOwXhf5bI4yO
oorE9+rImS0S4aWcJSNo2fdZ44SyCpFu+6MJQsECfyOodbPYclQ6zA6c41xF
hbXF7VwV5N4w6g6fPR2fumEsCopdKHsUPcr5MMpeNr8DrbgZs2KjjLqH6mzX
rAWNLR4uW5FF6j7M/L2xdjk6el2sm21TNOsdXuLpZpin3SPcUoQC7wxgJgw+
f+EeCCOv4W5SAcOufKk6EnR0K1dFM56YS9X2gQnHNxP+PZolmI+gEsrngsk9
kAA2BTOxMMTWNK9R1mlY8HUYJ49gPntpb91itqy+ruC4mPfFG4/8Rq4U63sv
L7hDuQjemWUO2FwPgxZYcsmjHurGmXDLmX3d9L+f5Jm+OrTN8pWDmJRMWaKj
uXGBiQ8gLN06iro9f9kdfmyFBhxhSasdlPHOq5Re8mZts9yLzoePs27jQisy
kIt0PvtBsIj4ReSb/CKecI2WZAWZtvNrrnleszalvYhicOupehSufMiTE4pO
A094vAvIuwuukme2b6lN6KDqUUZzz06SLom2RYCyOGfS4xaWgEIGZfKKNhs4
15kG+zhTOx0dJgyAInFFirDhevDX4/GPDpmAqMrPs2a+LSfl97FozF1aEDNI
rnnxN655GQJbBsls7cq0q//8O4uMTdABf3aOzgR+nDJy3JqilqXYu4JoekWC
NbdemvSU/wt2c839ejzS7NbD5hIrdvbnuKWbN6/kWth4jAJuVA11zLcKWl9z
Ti72V/YX+WEU7jOK6t+yshUl72q3NkghZbsR2xLFDZWZZYbVYV/tNffCc4JD
ZroibIH8Um10iqYUqgG59ll5X4t3iDKmVgwnWSrLIAf4ZJXbM5vRfO0/qKy2
Nin/eOxq2VyHR2xJ8HrDCiM2RaDkBoHQtzINt1d+zmDJvUQ4tYYr9jz0cgUo
s8djRyBUpV28UcfDdXqewwjHy8eK4XlUoK3HhsEOK2qNgw/ok772eeQMSqyq
q/8Ky+IjXLGQw6Xt3rGn0efQpQ3oCwkiTc/F+hRkayblbo0va2dUhPkbU4za
0RUL2tlDKuBbj5cxE0X8gWd9/yhkVLki+C4i4FVM9b334o+RUBOLiYU6CQdQ
bPAPxTBIsY2x1yGJI8MgYPoKxmqzv5oiBh39DodgjcUJ2Wz4ercYJGxDxhBR
8Pjq2m5xVo/qd7lmpLpcKZx9trweIO64UAgrAGOvPgDSQl2jVoD77anB2fI+
jw7CITfp9SvhS6UZmIEyDuW5AWtKVAHbd1lYRaOIWxD9cbVy8Nbp/wGSDEMz
UfNmeT/dOEUO5v4P93Ugvex+VyjXMoV22UNBc96xy/kqGMqL+gD3hMiSnEnM
xhsjtUsIlU3tFNt0r2GwDXn69j5hlCeZ9t/uU9APyXQ8w4ZhmR4bNvkSzYoX
1aULOIIiNSD6JuVC+QrKdngcZ/cWUYxXWXByhFcUbKuw40ZDHEaux2PXNodu
aU8M9bZBKoLZvnoQ2Fvh6kfgyLX5pnCETPDXdiZ1UFNDjIhKmVK8HUNTSY08
NLYc2/+5VLzr2XDXjXSHeh0ooI1kQLl/BvUKxkOrpfRYe2s3yb3JVYPmU6aS
9z38bWgFrn+gRAkrw7aXNCyfL4Eo8kC+wmshytsapnCCXZWqYCnTcH/zhrlA
iDR1AZaVp46hPSfjwCSM0xbziDY9KdNw7oPJVgCIZWjp5xjtsL0zFR0BcQvF
FDY7RGLxtPW8BDTz1yMXJVDcML2459Lp5VLce9J8URmoBkuQB2xsmpfpXZZs
VRWkP2UiIq4MP8v+8Y8YTdqqIh//ND40iX5ZkLZViQVNVC1SWRWUuOOv6SVX
PtMwtZQ/uP5hJlWEaXieovkJ0I/Qk5gDAUs3oU8MGZFZkfxhWyDZz1zZwrH9
xwGDfg3ZIVp+tq/tX6Fhpj4RNUC4pt+BDERxB9FgNTlcFmwUI+szRg6LkwM1
T5D9pJQXHCGvoVMLDnLaEqBVrcENyBeU7AaKE5Fl+VPU4nJsKBJ1KaqPpVys
5KltW2bd7TwAHwlxz52KHE7Ed5ggwQqEd8Pk822JtBGD1ApijnQte1lj0q40
NUC27vn+v7Pe2fRhxzYIt1wQmX044syRx5blxkg+oeyY3Tq1qRs9dcNfrfFF
VPtjqt2EY+AdJwFi8D+iaHSzfl76WbZSXEFVRz6TUlNQcqoZj+s2yQqBGqem
LgKK0zsPiSZIwT6FRgatJtIiyau2s+ki9shsZdv1tmeiwobe8J77+oUKdZja
gtt1H24GR0FxxxnzUmneR5hx/f3MRMhRLQ9us9kX1LMPNVzjOpbfu1YENJcE
rJXMxx2mcyn+Qn1brIOgjBCkCzxzcgT23Xdp8c9qob0ivoMg5esH6rmV5OID
HYpNgHrMmBoUT+KMR6WqMN3kl5HDi8SendaJA5DN1i16n4tUacowZXASrxHS
DLMBB5Hkhe0yZtB2mbfO5A+2ZefEvkz7luR5O8fwhE6nMDabn5R/hXd5qYe7
uK9CeLIbDYZLk4Q0ulI/4D2vJGxm25wFNFcV2X1qr2ZR0z58xDuvq8hw59Di
9I5VZEYIrE7TG1TxHPnMpLEdb05VGbKFL07hrMzxMRBCYpssQfmS7YbD5tNd
KQpqJWBVaplOz9r7+1ffeLTCn6dbz5bTAXJ1lAf1O+NlgLYvQ/NvENWChobb
LTU86nJv9+e9xuPJiA+DTEtKibOLrnyn1xjvSxOswXdQgqOpgSY3Z9JoR1Co
VobDH307kVp8Ysf5izz6IZb5okD0L/cgGBg4Ee/agg46lNQmAehHWSCsJ9wQ
WHOQHVgvMCgOKYJgNs7NVW4MNMWU6YYh1WeLirqxiQRh/PwQVntphRlMRemm
QKMjVI/pDr73FL5mzEW+bB79Q2yQZRTTRULvrE+Wtgs6WsB6QzVq8VHF0c7l
PYTk1LWOo6oSgTtPn9tCKs+jLwbKbL5OdNdHqFNGvexrNPcpBFPNONc9odFv
QYmU9cDYIksp000aOIqFdCcKBXeUafVzPqm9pfHc+y6+fD1lkQf3n0D952Ze
ggygv78javwcXOpiOnW7dcbd6qw7goqpErVwZQ0QQh+DUY21Uh/CKhAyUIX4
tk0++/qJfeog9bbSAzx6Gm/lC9D6drDPT8PJmiFappUarLZYJWVimQnDBTlt
OlO4reaH9+ySRPS9dxhY0cugL+JxGY0yCOZM+s6fp0oW8ZKDr00ssKxLOBTC
pgOKrYAESeQn+Ry7Cb2lpmhU8sFTEgg8rdoITGqgxn4ru49xfwix0ATHNlJ7
6WrFNM6OYqUFkhNGherbRZWHVJESXh8EkQt+xOJB2L4YteetftUb7oL17PfP
b9kInv8tmuNvFqmHUxClzzWC3GrVE0luHLhnSb//23f/cNP+En/Eun5QpJhp
13oPiSndDIGK/xxE4WccL6UwbwCTUogcqQ7ozAyyuAdIoI3EujppAkMCfG1j
iFj8lO60HEIGYbDbq33rmbxHjLubUOHlRNXQeOsjMFowt3jZ+y+DeeibTkzy
+0pcrsbeWPIQDKdB9HzDHKwtroR0FCS6vuHwOv3GZDQf1okcn+nRvn3cO+mY
hRDnL+9Tk3gD82etN8bSGVhGMX+YVXPFLiYdboaav3+prfoVtU3Vs1JB6TVX
Oge2dyCQcQF+7ZkNhwy1wrzficuFSS6gP3tSXJG/oof9bVNLdmbwAut9C37g
vZGV+Wan428wVWDkDSQj8RsfHOP/57MSAyncUtSAC8hgs5xju/lK+WDri3IO
XMUnWkkKzaYOdA/+Q89h2Sxy7M2uR6/1cd0s4e1XQwx6Gw+SeeuiHGWb9ylN
xK6GS4SnUb1OyYbgTCosf+YF8pXBuU+4S2UUsp/Svj8a1NQmP6UKt1UzE/fq
ZB9gW8TvmXP8R9JwclCYKnvKdx3LIxuCkB+wdy3/NSAoSVzHoRu6eoUJhohc
NbAptpyTmBWSNRJP1d7tL+uWcRymZJ1OHsN5Rt/Er+i8UDERK8kqpTnsSkTv
VObx2v4oQhFIEZqKZNvVzeAt2v6nyJvOaHZ96Hlu/Kfx0lWAUPHiJ0t92gxy
/fqb1C36Uu2yd7LpR3pGaqJ5vPONqqQRdpBnFSNwHg9cqXdauv0Fx9zCNq41
cyeXjbAh/0O9tmz+2z9jpxPRzfh50R+ThnwMPMKL4s4gR7ZWIzxGd4oeqFIn
FQp5lvqoBFPlmjIiZbskaXmQyaaGOSiRq9+Qj73+gyg9WLmNdv/zg/1Evl6I
Cw3b5dYWP5ARLL+rY1ESGKLUn1JwRfisS6ymk1/mruMVtS1NcpqqiM//MlZi
qoXPB9eBcVnjZLbxH8WHnCnWCAsTg9kZr+BYNXGXtvvTDHHOV9bkLXhAGREU
vaKUKxf9ujBgFsHSF3Dhm2XL/VZQuw6wZTaiHvUrOAUdKlUAzEkp5JGC1Xme
1pduf+euO8LafGa6BvrdxS3R4ikBm5xcyLXSef5hClqm6wxiLwHn1Q7IpuBY
9MYqLoBhIO0YpYMOfm0hg5xY+w9xPsI2jVn4RzXMec3Z8DPO4SnCdrYSJU4j
B3LnqIgHDrLnmPwl0oV1VuikznZrC8hcVl/glmsHlmZgq/q2UH9WNTMcjTeu
f7vFfsArmMVgmYuyCPojUzSz2cDoBm0akERCadLA7Z/YJ7UkjvQxQ0E83XoV
p74YP+kdApPQB7kZq4Kek57Hu8kplll3Bnq4SEwk3908yfAYyZUM2lUeKs8+
ZMPglmKKw18i8BBfHX8w6EpUn69D8rQ5jG8QlJpR0OwxuGyZ/wLM/OhZaCNZ
i4eEDxEmn9ybU49ZC24FOdqyHXbtw9CN288IGXaoBOraKMDGX+/NhWINfAZd
moq+qHULEROjguVQAnwKzMJPdtzkcVH9pSlJh6v2qBEtIDlZspTIKAgjc3NM
GZ9b+YoEGYcg/QY2QRBZt+rsPatCGyJB/SmOWkBIt/ZaiyjjvUwvzhArm32z
ZmeiTMk/IbgNNbmstq+J9XhHkAyPtGrIbTEg08Gml/PxTtgVxcZAqWq246/3
qaI5YZToyBtDoaB25YdbtZu8rXScQld6Pj/DsYKdIB3tngUG0myew0KeTl7U
KNl/SzhzD09dWXhQMArDHo9L9Ugaa1OO0wICiyxoS7zTagLioicRKbvP61JQ
V2myyFAtK1tEcxn+FrFkJ5HayRnWSZRskS+z7xp58cJkB4Sliris4Yb9pVmT
azkgvbDvQJPHycrfiOqQCoUb+eJzw+ZO3hCvDBL1JegbpMmAxK+fC5zSbLux
FOZhh5a1qAFCcQc1QAfeF3ttoM9WM6LqUYQ2BX7J1YE/1ROgkXOz/2+0ctnY
VBQrE9mbY3wgGdgU6fOIKz1RA1r1l0hEBTCuJhdW6HuSOPxcoVb9d+7K37wa
XBUSDnNQ6bya6qIryct476dtw60BqHXLoqO8aNBeTCikzfTa+6Z1dhlRVmZM
Zl0QMPhYoJrQBFme0Tjmx/xW6GI8F+ZgxZQ3rPgwMGilchPfDSLET/ac0AVo
RJla8NcRd6xNXw0qo8rS8MW+f/rZggEKW/OfZxCscCxpWL1BFD3eEz2jUjNF
Y/QCScZMRiI57EQN70aYi5X+POOaNrnVYeaDBSv4p+YQUG4bE1CF2v6HdG5J
dBuPJWsM+D+JWuLsjWgWcPGD0vyGnp/1Mbc00cNVYxY+gfkov8XMaROdwZNk
45Sn3D01hL2jWFRbBaSG6c10rD3W09ZTsmCuydZTNRUPHYivuQ2w4mzM100y
WTJDMSy2k0McvavvEQNAj7eQjNNlFJBoqs6OyPJLXTTghr9tg6usn/KtfEFN
h5LDyEAtm3qdhTJoUpezjTAeNr6ehwItmf0aSbfysHSO52QeEdfNwULhnC0i
uMXec06EwKKpEcmAA+cBhqoIGIE+cHZh9P7amZ2s81CfVXF0dDqTt5jkRUco
vtrNqtWbdX3NVsY0nlbgHPj3g/ozoE/Wbhprqq0WIQC3zfDHzcLGMEAri9PD
F7k6S9X+tsF0ia4Nlbiaw42sBlB9brun8+W9GftIPyjc1iAVaLa5JoRY6xfs
YRfHX2YPA97m3TmsNuPX4RPY4WEGPJf1iilHRBh2XecBFU9/ETIn1Mz+F7Xl
mCN9a0LDRHzyCwNxc6jsCl4yv7gNBj1osTchLPqFOuAtCHRaCSb5Q0oLYG42
PA9m8kfcUGUb68lnJNM9IEICk68C9hWKI9vI09WbZdOv8I/7bSXcIojkNDRE
zERtJokWEv6sfUTM52D1+ddyjaAzAdaSM/F6+gyYUAswUC6Cpj2RV4qERaBP
orFSa83dLFLjgmZuFPZrkcexZ2E4rBTS6Lqmo29r80a4S31s92/7Ky5g6T3j
bL6aJtINNa4RKlXStPojX9bqOfrzQN/QBCk/kOxQ+mzi/4EZhSIWGGgp2od3
/LN69/05v+4jao5/tlGZfj9vB4wfNZuDKHB6t8Yz9/v2o91i3kjU8mxDn0nD
86gBQ2GoTFuEXRs8+8LETUfj3lP/g/zY+cWIf1l838Z3quA1bZsSbwbfyZBk
ToAKjlcjU7ZAYDNmEQL99hg3obiAQByM3XaAuNnsMCF30fdqMT6D+IUsZBHW
bCbl+D4ASBEyECkCQ91SCAISPla36Bg3KsueIX9ZAIEhufDlKQ20Ok1AiOuq
lBIYXYMG2vWuAhECmEWg9iXv2yAHSQ7PMHkk7RGY+d02U44+KvIAC0QybFYz
ieS1+d1364Ad9UMa2rGOw0odGqXyjNJkiVy/V23U2sffA3F7jGt9t6KaolVN
bbXvI7qpwVwwTgj1WXMef1s+tkDBEJrBZ8YFGjx29SjW+zyP/SH6KbMRkQ5l
/ezCdgfEKiaNXMQC2M1Gp0Wj51siVq89P9BjaM3br1duHwI0zaDqXVreweOt
z3NLSZVO33ucui+BPePUGntjDqVrRcdiesfBzIsB8gKisPe7BCOBU9YfnuLe
LKiQgo+f7+GyaHyvrqI2a5TviARsNY73i+UQ87MleMBMdENk3KrycVhVpyWK
4MR+ZXoVRgDFWcDWsCBggWcxOOI2GZT3KeFIWUJ0kUCJmp6Yg4atsbcQ1lak
EE7ZRFbLdyVy3KP0qI6MJNfrXUnjIm1qK5AOLj7w+avAsB38ITKA2gxdgzXs
+gjYW7DTTHCp5fo3CWSkOrs79lam4seegJvwvgsLul30d5yQ+AmYJKGEfVOt
EP5+iElvJ2jZv1YRxS5xLv4uhju9Az/UfXH/3QA+d0TfZZfwvsnfg1/htaFv
bJtyf7HcJ8+ASqdXkqnyfh4A8kAtyhvN4KOMSOcHsgPNEZG3yK8xZWhWwG5s
A6GN4OmzIkHdqqk4NLG71SwfnmBn/OZNvkg+DavwXD3dRQAvQ2D0ZhtRVi9/
qYwpqCbzaypaI5QsqHjb8sceEBdox1osI6euTlTBfOYHy2b6xC6ihc4O7lUO
5EficAY6raL+5QUVT5thiIzWh/r8vY1b721+nQK1llhpQ5rO7TxdRaqblDCt
KuHWiKkEUHhthHlci/qwgX3euc7fVctKiTQZZnGnkpGjxSaVcAjfVj7dM0bB
R+vymKsMBzafxcly+q9JjJ9dtC0uu6pF3hMckDJ8au7xINm5XktH9H/w4dap
oL9I9yTG0143d7BaTUKwBAzVblJFL1mOnZAOMt76s8YrO+hsy7i1D5zlPyHk
6kwM3BT6qcy+ka6u8K9/Oi11Zy3o1u21idWtBF9g504Tgo8SN9J/lD7lQSAH
TC0cPCDMh7Ep0CCF3sZM2Xptru1e84zjM8okKx4JY2ZpIrQOTKArmCnflHG4
6uFLCxylFQTFIS+8vwn7efLXEhbZhzRrMjSXLqxBJUjhg8ktWK8edx2NlOuA
Fj3QQNUQmgtPiZdnpKZCzfqTiUQDviyrBObKPReYyTCSQmE9bsJx3X1vsq+U
/NbqtiqaqgncDNHkBM8PEb2D/7zOM3hIzVSQVKhOfZPUQkLj/TgvNav8hdaO
2inEpV2evVcOMfepVmo48QjBUD91P/zP9XyrbSRjDUby+YsBK5HaGOvH02zs
EUXRq70EMYb5wGFBbzyEwMYYs/MgJ2TwBBw1jjg9OeUSKcL/yqZt4OeVUk59
MI61CgC2LLfG9DSTlE1jo5vf1TSPaOaVy1GxLnuoSX08ZgAJuU1t3dIFDQvT
ldX/FuXBwhlhqv7N2RfTfJzE5Gz+ydf3dpPVDiHnJNFfsDwd7KUyiJv7DZO5
KP+6Rj1xgD18OSJvffHK3MXd0zYSD6huFDCYtF6zH8+ORuYPykb22jLfCs0s
EuEQHiWH246iZ5YztYuXp87SEea/Zh7kJn0t5kvtVUhdPnLihiaWGitcnscH
jQZ1Z0EBQSna6b9GTlaVV9M2hePh0GeO/koirVXB8LqIIIvlKUOnIBuh3Y4g
H9rl6Vr9DbSgO899BoIA5q0g/wwSjMTa+yVH6H6PeiSJ6ODEDklD7H/VQEcy
y2aqUj2dPw7q2PL4N5Jd9O796xWfLP+fJzTXr7NxCoQYBWiq3Dgg0zPgljsX
I+rY1w593MGexHPVXj/SO6SnBtxLwwvg0RK91Mzzj1PhVYtVeKuWHga4rq8P
fqtvMwHubeLQWFyfwDplTyM7FyomZZ69J35tzNRYFtPhnftHOQaOTVU9NAJB
AW9pfbEqsXHR03Y0Y4fdLskD9N/4MV3jdxek5ECFAdJks84Ww+q7IAncug+5
Wg/bMAG5rTsa+kB9gyymboxbsMatDFceKsI9V36P2/qb3b6UlE0hg92EuTcX
ETSYuveMPnFEi3V9Er2NqgINpfaxEeNY+hc7l+Yke3gGw3Yy49eZkW1Iztrh
+0qRRmS1CkWa+JtI6xBbtinCmlvYE98J/gLkVTIrhDPLF9YGu+tUDt43Ypu5
5X+JnVbr2F5QYKaboumniAxOl/BCCWYfQinllbuZiQihuYWdJNpRRYzasv3Q
IULvjNKt7bT9BioaJDKRGSmqFxb9hXJvNMPwJFMlEzl3C0SHMSTekifX7CWk
RR75L2OSTSVkneki9wfTXnHwKh+03eH7yoUV2gzds3M/kMo0bSXPkUwaaiwB
MwVER5knzfGGZ5sHOido2c75irO1fgzA//AxVPcsAfkWRWHrh71uPf22r7jj
n92h5Z+PICKQWnZC0BMl2Ig6/oA14cinz/2UXRj/XOgcdKg+2glH7tDqQy3m
giltPNq+t7A2LZ/cfab/PabzAznk+TV+6BMedCA3QZ2fdofyYWqOiAptDKlj
FVyoxaZu+WAafLHOHgfbwo4QDdfbeRXy1kZh/dVHGnawQMgF+YKZHay8MToA
GLxw40bdYKwAc6IUxWN4l3WdlfCCcjIzy4NIvzAJ4kvwiVFgudPW9XJhTegD
ZMbm+nMU3hTnhK+jf1AVS9kY4I+vcTR091gxuwE2tdBmc553KWH9B25Qxpzs
/6Ui5Sdsh9FhjE0wFjlO6dhwGYJkfPvUPFSUQ/VltKmKZRhN0KiJSSEjVuaU
4uIF+GlmLZ9tBLDrVs04Fh+D1CTpioTT/zSr5uZojEEA+9yDSSfsBS/x0MHl
f//XZCoFecXoTNT4MQ1fyFYx5bDPgV+PL0F7WIWF1jF4IjTxZB3GxfgeVU64
3w0KLRAVIpQc0O9rYDFKReYwPAkp9YChYaP9bSoqhEs6ADm91B3ajnie1d6E
kAHD9oiAOR73YCTFtCd+U7bEqkY98dVE3ej4pGowwZ0qdBB7iPf9gltb8m2Y
INa0jy2KDMA4De/eFTRgOOhrFGT6WVxSYibKHNI2qOdHZh9uUzk1HcSbMNAH
BaoggV/ZJV7ZHkkFanVQ6hl36yGJr86WrsqiWuAnV5kvFGmfWn6Hsu77YR3M
yM/8Ubpcl0EBlzFDHCT9RpvUtZQEjIlivvfPtVpkbcYS6/LnktqIp56+yS+3
3s1jhIYjtxx5LtATT29YqDDpN501VtSs+ZzgRgBbfNIoOn7kHnN3wAD7BH8a
aK7XC82DckiR9na65+oJLcY3epGcZ3BIYFxFPkZlm4L/2z2RX+1pt6YmGtCs
Nl6tK/8q8bZf5qMPdgD1D0+2m2SIlk7w+a/SqEjKWjllABBFn6bi1ec7R/vl
lbPyFL3TxHO6vw0IgQp1SZ4Uh5CaYFsJ/O9+zqXVZPOI1X3KoCPyRm9vbOFc
65+C3ZJmqOTkAJu9u/fPv7s1VgG3AYXdX4Way3zKJrIbPMYWh4n3JTiWYFus
91pYX1IepSeniLCAAvGNiHXa3t69XfcVoPRdWGh4ifScso+GJRM457ZL2BVX
sAbbII3sokvigUIl53tnfjsLMuItsgysskOALrHhawmM13v13SdSRBvybXu1
3HTp2pByBB/LdbCW5NGkPsZFNXW6TuMo3zY6oA6jaJ68yFOxTsSK/9cej1/G
TBnUrcoC93eM0ZJuQm6VdRcIvWYRNR2USDyJeQEmhtkDhgXb769HaPOg/WgC
2sX7WqBFdKCddR5EpdJBvZ646KuDAEmf00777W1bg6JA+upByh1hIyzmj4xO
h+JWkLE33lIQRh25UmO5M0B83eRkFnGp0HeGtiunMplssKIQATlf7DnXPOpE
/frXLv5Kd5Nxh2J4e+JZF/5IttBHzLmkY7SV/7/+GHu+KqmXXt/t3kbto6zy
gqxZkn2JJHfsDAyeDmBkdlg8Blim2iJc52M6/y/+5CgTrh6c5WHlMJX9Az08
j68wixWawoTE+51DzCccJiAmHzEEmJ/ndTTvYQstlZNPuB74APHXMRPNcV72
B5zo/CYyEIOSB2R+5CItcN4YnPmHPrKDIlc6z7XJHa8tD6MR2yjj1jmGYAA9
sOYp/x11lz2gt9u2vnv9eVKk1lTn6cgDgGTmHsyq3H1sXVo/pLRj4YXRlZXT
BxNoot/KJQqL/e+4oqPzqdKG4Gu3b8OR71AbfyP7I9TVpMH3sm8s5ya0f5RU
WXt+CQfM/hWP493cvsTzm8bJ8pUbRpyzzEK8liIs5FyeR+Nz6nn5evrC8pET
vWmQk0HpjLg/gjicdj5WmT1uRKrtRI/Ij8/g3X6iOmevYjqBgQTnvtC54Ly3
ja8mu7Hx7F6h5s4EP5aE36md9U/9ylNdQBau+IQVdejwsBwiG3azvSHSWdfn
S9o8yXhmQmhQS3JsXojaGy8WzyOguWBlqFOI6DpftUany0n9ccPvK86is+F3
UXLBWwZJ49lDiVdSsKzOSSRaYdFzwHDSTApL7Rnot9OJGa0jU876N/UA42tE
nUl0xBYuDw0yeqJWCPQaAiBdO8Y5ZQp48215kSG84czQAFewE8wsGbiBmbZm
ZWMQCcqONt4dNaOZkRGGIRefJolVkGlm/d0kl1Xt+zDwUxjp4QAi9Hp3baJY
QeRwV7SvInDstMw3RuU6cHFrP47gc9aytddFHS+55ziX/rb2cIrbvEIgL6g/
sMNcP2Y3i11xeegQnZaJ7Vxo9Q4m5/W4BluGmL/+sFT/X1CDiOWcS3x+7DmZ
8zyVGmfvDTaKBo9FAmmhSnXaCjnjpiLBZ03y9jRybjjU6NViMzEVT6BluJ9Y
hhPrplnebShdfr3m51XlvyHJ331B4EBkIc8jYKqn0w2sPHV0kro93BtNigVC
wS8nVwpvlhqE5O7ggQeUVFpiP7qhBYrTPl+Swu5lYKmxXY/L4fIU5s9auq/W
roI4CwpThiS22lhxoHDtJDBdNdZvf4NsPXgcMp4apaqqqX6Eh/XFCEgv5qKX
umUXDuyujcH0WwpO6AG9oaKhI2Aik016qvNBSbvBXwhz+OI8Kjc2kTgQQ+G/
ssxsQbnc+ipCdxRQm27Cxy6DzAWicXISPc9/Fb0XZfkS3H2BWLSHFPYCmvMc
o4YBvqTYcf4VdITcH3Dq9psICPO6pxdcCcLAulffuHIUw2TNMvjTWtFWhR+A
d2pphk4m3fvX1br4KLfiDODSyQLG6URZrsGK2ydxQklWGoeWxWbH3ko5kwcZ
626fkYa0i/5qnOri09bPAnjFRSzVe3JsVsItMSltRLbW7zrDIwhhbEUO1evn
9dAswzlcH+j7GrwtYjsML1emJIsZNke1Fb5+FichWuOEVSCr+dDK4jDAa3PL
XRaDDhMRifW/UcI7vOWNNA3N9IyeL+rCih4Gm/EfdOR4mZUQVFFqVo8dljnV
4zRZ0Ja/+bPzXNw91SAZGcRN7Jva2VcfHRsMx3EXzfAb7OHhSYikdqE4FXm/
9+WcwZOA6YCffsB29yhF/+fEHszjJw1qIfOZf8ARkhdD7ptssbxByo0NnQ2M
soNNFsD+87bC2ANfVU1ZC7Jn8xuPyFV4DCyPnDt093h0XvSck659GxO/ein2
tDOwPytO7+eZjss4Dc6f9M5m2WVjQwiA/lVi4srfnJ1myMFFQUNK+cYE1xgv
qQJxN9JrOUGOPBi71sON2IGeNfZLmLtvq0PzpMaZS50uEdQ8EDtECPZmhHSu
pWGvnG0B1N5Q2fOLg885sjwKBr3c2rZi2QuK7HhKUjaevCJfopKl7i1v+0dF
q/FzoEzUtTt6SNOBn86uekGFBjRL+1Up0c+jxMgDwyg59flirOvw3GqoS4gs
Dxuz1dv8Bteaz/JvCRZ2sVadjLzv0Oz7nhVZ2d7vT8j5+EGl8TQWY0H0/6bz
ULs+AxzFxDmBPSxasTK9iOwIjz2XWwRqv7SNcbmLAPyz4Dvmw5fgbKvW3wn3
/aJYFErlX/KLwSX81mISdiTCHOybnYF1nNNwIxMk/wG0rOKo17bvCM1swPl0
0/WlkyJhNeG7NV/1EiWwB64UvSgLHQDx19/qeuJPVvF05sBCxE03V+ndiYeq
Wgn9LMkS2k0oopXUuXhvXI1W91qxfi+ZAgW43Ic0LH7x35ObGpWZDh45A4M5
7Xg6P+fB7Vrp+Gxt167CgUfZkT2UqHhCm/D76jyctnEJQ5H5qFT3TIXjzspD
rQJyKzlQ3EMZugQUIh9d7NQooxvYPq9mGN4TbTGM9tauZ3ukqrmyyz3WMfAs
PymXkBkN7LbL7Vi2z9X9yCEmHfW9tv3plqk61yfvsA7T1+UTywsh4MlH+V/b
fYD3X6ne/ITgpIr5DGC+3pQ7RoKiNmpXa2qGN2ZSmq0HbfHdS5ztVLjLrQOD
SP+heXfNhWY1DE3Zh8iK5Y4thc+FuD0Wy9nQ0eWKXMsKGq55RyU8c2ITaThi
jWorKuXFv6uu+cLnZBIVap5cTd9XA2R22q7mX1cqofBzoKAgTZxvGLO2JyKM
D4qEHZ99S1R6Wl3U2dDMYZace9pkcjOuhNBwt/7yHys02NbuSoxLtSfL/4/S
pBH/1ukm66MfMUkvwdec94aPwnCUNgbXONFX1CYetgKJBS9tlxIFetHd2HIz
iDZa5POLyXC8YTOu6MGcmYYcgmSs97rzwcxYpEQZ/GP83y2KbGcdeUn3bVtF
Q8DoxZGz8gJ9HdE6yo1MqItwCn2f8iHGocfFf9inEGwUwz+K9oV/JuKfXSKI
uqTMzVmBMz53MCEkVecGqoKP2zX21kb+x210K7zBDfqk7nt8EV9kGi2dToPj
F9FhpsZOsoT5Br9CosuTsSUHJP91giLbQ4HkqrrffhL2G8svUC7/2nh4PCu8
WEEtNnFZQZTI/MIN9MnqqdUBZVzTP/8+v6B0MdzdKN3DvjDAE1fk8glj3XfI
GEHTifOTG+SLYK+T1tIO5m4jql5ywfIjRJoNWOrFN1J975+Bu8Nb8Uja/mUT
Ks07Z509U9V3vIR5014dtUABhHhagbNmUC17wjdwg6M1UxFuvgmQ3FyyXuHQ
DloWbr1sPKkfpyVzfEagUIXrBVJMadU8kLUXHjhRstCLwqPX497PS3KfL4F3
UcxXlhv2zuSINvsZBEYl3Pvd/QM31wuUa3azSKPO4n1UhDYBJ0kpTXNTNNQf
kyCxKh42EfwiptEZf7bumx+EYOzLt8XVgEtB1nEv20vCykP/UWngzeil1MV4
DuPBSil6OcjuEPBeuuupW1CS3hEGsHZVges44jNOqZ+8L+2b+0hBKC2bJ5A6
R2WbLb6khcT7uFOOd4tPp1Z82KYoJDHXrJuXtdFhUvHD4+lajgw6davJLyV/
+U2Gj4nymtgynkWtjUdwqLZDrei8ne7NgkLdWXIUCYFlKvEwI06q3/Djcvil
l22e0h0rk997EyPI7TQh9QPQmFrYwHSUYxpJEecGcVVSjqx1R5fxjs/Kf5v6
MSSp3ZKTPwh1TCohqWEVtGQnUEPVfJKBXrbYgpbwiZnmShHCGFBZWCVoIfvb
HIix14ho/qiZMiGuhEQac4YPVBZCizwbhltRIUWOoekM+SoIW9z3bWvmyEYk
61I032h7CgEtlBkIXkgkHZW7P/1EBzy3/znQj/AdFol5RI3TjIuzloUyczKa
vvSvMQfD2z8Mkvae0bbnjg5IcO9VD9ksWHO8/lklSrq4H2+REI10irNrtRAy
6SNLo2kF+yYjIsbQAnwvMLbMuFdTXR6QDZYD/dvInBvq/ShtgB8JPj+EcIm0
q+gS7FXoqjYBFpd7Pghw7+s2gOmtJYJ99H4Sw7hfx7ydwi0U9uCtafGbGHJe
jKq/rnmm3jjsGc02ue8KqiaZMyJ0/n0xJEnpIn+5VKOQOqldFJWmwhaGXAR5
v0FpSv+xQweIpEWmH7Ji7m2o8oqH8iP626oTRn7ILNT9/kl9RNusWHrLCcFD
l5cKz2BPa41X7j25wY0E7KwiKaoXjYS+3wF6rybZtEE9Dkb3ErnodfWs4kAc
HA/eyFeWpndI8cvfNZ7A7QgnaYgk/XQs6WWJEe0CRIyKwZxgmDET1Dzqtcz8
vvcgZvi42zt9ggOzuratIkWfOf9NJI1a8V7k4SVkKNgusanUydXJN27CvyRw
9pwyMsoa1JjS/W5DR8z/zzY0oY/SMHqj1xIm9Sj+k2WknfvbazJryGhtokiQ
ekhIDVwty3W6ifdOYYydBlvwu+ZlPeqOdldJHDfoxoGLA/UqWO6/I+7pXDmP
X7UZ3NQvu/PViKIS/wN5Bu4MxdFbOYckO2EzHBLPb3U6zpjYev0FA7/KUtCs
32umBQoFiJeO9HuUAjchtD4Vg59dV+9APr3H720uLJZ9Vk+8PIq6rQwcgRHg
7vMAtA7E74yfmVMZ+FsvYGIvFh4uRX9IySB0rOLXzA6PmXMzFdeBwm0iydqf
blg1SbpkiFVq4H3wTwPwAidNCo7ds5aa40U3Cu9rk4ZBc3rnMJbBIggFjEk9
kfRHsRrfwIG8q+NmHsioq24dZODOdQBU4NjpUTgnX7Gxv8+iLXBNH28JCyMq
bp1EFj5tQOq/TDeAcLk4PBjT8nDmYWdnNV7hEqXTRYqLdNK9ObYKPbgcVset
4kUpGcUdB5ERNj0kygT28uQI8iruqNoAUhOo4YlEpyuG111ySilB4GtOLWJk
zusFTolt5vCIYK/y8hbF8wmS2ZcarcrEKFaHM/8yGbjC2lWseqCgdPM7Bfjg
i60sDpfpnSI6HmxY3479GC47iJG1EjPB5KGZim2FE4vkabce10qbzr+QYhc3
YGfQ6F8V+599LUPkWUwNWWvyv5rx5oaqhR+GN8OB7S/AbTcqQLm5OYtx6Awl
yvWps4ZZEEtWZMtTmupcLEukkAhqmUq6ZAOoCmh/C7ZLpbRbTdNrbKFy1zrK
O89WIRjISY6J1aqysjTPvW4RBpr46Aq0FhmbWfJ/Fgz4mB/QquW2TkwYXmat
UQ0QvO69/MaXSRMA35v4wIVhfvpCX0YtVhod0SgriZ0cAlz4lnpT4rpik9WX
Ytue0VMTRelaWPSCjb2Tzg6f4I6PWXxBQMgWWWM6C7LMzUGM1qiuWrUCISG+
CKAll9gXhUZ2j8v8SloMF5pSN38w/APteu5fzyP5As87c3B+1O/49rB3mOLJ
jOl/s6WwQ/+hooSYgEbw0KSLW0X7N1C0ptKbV9E5cq1Mb9IKlIXr1B8TWXkl
JhXblkhKFNPyqF8m1PR+nhHwVKqOv2SQ6tDfkHDdcjtAFuzUhsbmCQSGvryZ
mXg8oFN+nPLBglB23fIa7QWsIv3o8E4Gdua2+2Lk6QwM9rWJW5INGrk+2n4p
nET9iffuBel5t9/Pz9MavMfouwecCVYvtaj87VcLf2g9uH1dCS/11xY9TI86
zQG649nhu0Scw3FS773vN/h4gunDFZofUwmmopB6KKVAGnIWAj4cQfudoZyn
q8seZq9PjjLTAVyOxe3Mb3QgCT0Rq9XJL8VWxW6+kq2ZAD6k0b1iCNSuyfWe
R/SytgiJD8xsvoqtA3crhfme04fsyFr5BjknlEcoUXaxoeBiKj1F6rTU3k1w
MMILRsnovL2lKk+mTBNmAVVtP65foSGRW72v25luydvkK0bUt30NAGWC5hFG
PAGYClo6Krp0r1A3sAVE+SO4+2zuOXi78OqNVShO7QWdnI8YexuUt1ImEWKk
Hi2w0tn+IzKj6mlE7dcx9rhX61NYnKXOeDE7ik7JT1Tyn0MQURBsB1tHmoUq
NhuLeVEPHhJ3mDOAsVlxEmuOYaJUz7dYlMYOTMSXjEHGvTeHG3ELlHo84frm
+MNuowjqzSn3wJDTmH8A6apL9mMsFgmkHNudnwF06w6Oespct/MWPTo+MtEw
su864ZBy2CJ1LbGVGCZJx52zEtDNRCPrLmiJjuo+N3P2hx8DjlI1+PigZuCP
IYSx5cXjsEnOevgpBk72sMLcGPjnrkWxzr0A5HAa1auhVsws322HICnaetbo
uKuMtWPVfaP7rjy4WuWI9t5sMKGpc9bKu/U0pAACUnDP7Po+HpUGywrlg87z
3gq2SfM7dZP5eYn9X9k4ejquV/++x5kP7a6QN2I1PDYLTMVh1NR/NptQTbxG
3Bu9T7Dy1jiKNrKlcKCTC41RKpr8ImdEd7eiLuEkzBVGhg2YSHr0ht+xQ0lO
j1wRemyEWJ+dxt0Do/4UQqYmaqjtZzX3VqANRYEyjaXWtY1aRfQ5pyGr5Ge0
sm+FBueXMZOoyqmezTL55sPWY7wgW8/aax6ZJ3cVQeWnSbuPPcFEEGTKmuML
odlTVdFocMpQEd3o+/59G7uiHqR0vsr+kW2sypNOAOMyyS0Ztj0n4Ui8MzOb
zVrEL1y+G+DHJMXDg2EVpoArKDRgkhALF803wRwa1hbakK1o5oRXf9GO4IkK
6q5/Tcy6NgvoUYf0ZsLTR66hL1EZg9xZrvy5rHkQ6YsSlIgpyQ3Qy/kqKs0M
Nch3A1OjlHDCdRA0pA3SY40B53FJIpolhjXd0omt+0+HsCrz3tMtrhzPLk3J
zoR/ZMCsU8Wy/ffUIWzODz9G7YHJcGu0SCQ8GGgmQRv/iLasOMKPMWdj0bsa
Og1umowAB+GbKVz8lcVvHt1B2V4PktntKIlZOVEhlc3pDY+klVy0a0WMPNxc
KgHStQlaHg65+BEys/yL0pEz0/I85HLNrYs/yY1cMJwE5px8IKTEkKA5x7Cp
LbVI90EJ3f93WtmAUkjo9Jgtv2XEQ08r9Q7EgMsR9kB2Iui3V6pjcb4X+i8u
Lo7XSpJH0DxgT1zJl/SzLAfUySQQPg0M8jH/AoEBW94Mqa4TpNJT/zf2umBB
cF+I4E34L+/6ewXiEB31PBRVQ0wHhuEyYGEtFflC5d1GcUiVaSv+1bLAt1mS
oxlqPPsLSKFMIxym5zw14q3lBAnNwNiwVqeIRWKH7MV3OlX5oWI37yF1KDJn
4udf5YC6qJJuelJhxsh1NY3F7to7pk670uCk8AHEV4fUq2alCo6l7G0xFVuN
JRt5T7ahIKQRyLsk053UJhd0luR5aJoyhH2/RcSHrZR/u+pXz1i3Cx+kIR8e
6/LNpW5iEkMurf0jtlFlT76tivgwRhJok2cmkXDoEBGx9i3Z0tsRbtfvYuNB
sZpA0qb2LdVB0KFDsbAKTRbuqVJ/dXJA9LglQSqKGeCFb03dnxq1R1+ZAM6X
ZGzxOb9Yev5fDWkkBTt1QWOQuoWvuzgTIxJt9b21fy8T1Ei4FrpZ5o1PBIiT
z9CWUUhkV0Fd7sxCkuvvNMLY1iNuqpB4r6g/S9nsS5SiWQhgla+ej+l334z2
ElHwm4WM/isg/9CRk2+QBx6fzDX34vUu5r3Ch3uA6XSvl/k4TERqrqkvL5L9
cv+wcMNcMa/RCTy7DXga4iLsZq0JImdG8J6phPdzKtfZcsKUW2VAitakmyUQ
netWTIaHk6b8oe2u2R4Oy1TEVmWp/rrKQawgASCvKSRwM1m3b/2mfbwAXKDt
SzdvoJ1leP5axW7/nik1m3CfbgQiFEmG26S5myWbdVMxCAODvo78EGXGY91J
S3L1d51ghvHpPLX8nH7RIxzVIGJbkzX/GHgL1TjPZq5o0dQUoufG3so+L+rP
QZkoPdI2udaSKSYThpSqgN/KRJ/mgQmf3m0xcQK7d8lU27hOop+A0JgBXZGx
CZMM8kj0B/ktCUGZBB/gWSgn9qWjVWabxlznf9c/oTAc0dOlmc0SgbInqNws
bO0gZ5TKAd10EVaE0XBphTm5kk4pnDdPirPBg7TtH5Z6iq0uSyNw5fwigBIg
r8OdIQnoC5z9tZhyTTqleEyDVUNahZ3ZY5yoTbuZ+wU1Br8dDZxOygJNrCER
aaW2eCUJ+ZKYpX93Wr85sTfUI5QP9W3y/x9/52jVaVgMVr6iHj13winNQzhm
+axblJoJ4/1bjQsxpYjj1J7IZRU7wB3aylRkHEbfox0jLWTSU26ROm+N7u+h
+nT/tojHvylBj+dDO3v65amMXGrbymGR2fdx9XKhDpT7jcaLtTaa27TcXruq
rf1cleNHFj8Np5kj6Ri+0esQNnXohFpUEFazMudEA5xnzPd6T+utbenh/rHb
MbnVE3Q/C4Nz1hZBOJ4BrIS2VVH6cTVNZBR+yuzko8b7quq1Hvn3vihLz6w6
+nosMYRAhCFcd3MTqceADNroCln51OdyBUReffsVu2Wc6GeM0q9eL6hpv0eE
txjoBdYkNUp6K4mOMaRtbczQIG8hlw30p7no3VfM0feyR42mZqxbKS7T5FFX
14tE60+TykItlMPYI9QKWZkXIMK1YSh8lV9hg91Tv8TdqcOBSI0KL7DQI0+L
4AvpjW4RkrcEXrC9K1+pYrYqh/0Q7u1xIsh7KwIpMhoAJZ9EpgduUYV8cEv1
CJld3bUrSnWHtBLHEh1AhXF5wp7iaulKAUJIbCTYoWwROiadWcid5/Tz1fgB
DCryNVIJuylyig3wXCb3bdywTK+HkdsKnkNPXrf6XaoeAt/DNtoiMf1t+zEs
US0Sp1JMaK/sNf2CzPBxdni88nFd005lDSVejD0pl/a69uu9TP04UY24UeLB
hY9ub+ITdnXjrUJRx9cAxM/0je7oIQ/xuUu01Zr1mX/CNOkjPEu/PwARnJdQ
uSMpX3D9G02Pbyyh8j86T0K2lgEEdduXdWN3iPZX/gwXNEaAAYq/55eBYfmH
iEA1suFn6ZHfq/anEmSsKvA5ZxIc9vsA/ffRpARfnpL3iOegKTLHyizD8eDK
xiyW0bJr8hM2ZqEQFdQj8xdpUthTvvviX2FzAtx7DhjqygzcSg1CWKEtE8ld
vD2/A/x/kt7q/hLiArGYFBdVsCR+RlaLsyi/LhIH8m1At1XS1B5Y09toupuf
cHLiocPm80BfaDBSBq1bT/2b62IUmwR9W9y/DfoqUoDcBm1A+x05VbMTzCZW
d8av2Rg0deEYldg4XTLwT5nxlPqdebXxoxjwA5tB0hiXejY3RZS+n+Fay2Jp
fyUx/aVsz9h03apU/oKCOXbOfUFpMjI8YfpxXdaxN96hEaHOVTwDhoHsf+Yl
YJtKjvKdYryK1H+iSFejh7lu98ols3QEYwNTJqAZGBlrNgQKFVDUpw33BrYC
FKbsMeZA40K6+2nYph7yVzSH9g0UImygn4y7cGmJUI6Lx7F0PBMBHcEl0Vw6
nVU3/Sbu6Jeie1YiU/LSpttrg0jffTR/ItIc+LHfrz1lgv0N7VBoJYstBl2l
L+FHxe5biXBTEgK/Xu/LccfAOmi/yrwTxkd6rvpDRbS3RzOFtisWHExQrQzw
j/Nzz8e0OBQRUKhSmT/Vfwr+f7jNT2j4QKBW4S2ZVD4PGwqn7ahpfMEz5aOI
DVie/iDwMNLGKcU22vXU3YW6dfLHGl78hpfQCx/j9aaDWEx/TANkGSBTJZ9R
5za4oLz8QIe59Y/Sg6OZ06gT84nA0w5a7hrWsXn+WZDs4UdRKp31b4aj0Qj2
A9nnDX4iJ76P0xNcgEnNIyezkUZehAbqyjZNT92N3uHGYH5atY1CX+wmH5Po
TsfZ+wOAuDvdDPFZdU8hXCaZQ2Wm4+RFJ9EpUrRYyRoV4Y3rltREs2pPu532
4IzSn3Y23xHvzV8sj+hgNV/hp2E0p37+AGNePMNF737AXG9pUmOj1f4A+LgH
rPHMAMqrY5RQKYRT9OtFYSCDuiqgUk8jrws5nkt4irGJj3QnTGro+DSTaHzM
dRBcC1rg5sTb2t3B4Rar9ZNntuMlPSTKQxk38F/2O/hbGIceWEgwjqpwLbIo
RrmrTqJm4Fy4Y+cJmboi0ImQ9Qyt2q1oz6MAMKIAZBGzEN6JaM232mUgxSy3
XX1/c8Z01OrxTZ1qRhlpeGa+TFpN0mcS1LQ1yc2xN5FZm57SqHemkjop/SDF
OilJbBQZJinYhZq/XL19facL/ur1UoGV3mq1+8Eno+SpUJlQDlwc4idyjgxB
6ixYKfLE7HgOqIw0hoNRpP7lM56+NiNkV7wPrF+C09LFAtWKNHkdi16yAIRj
14R4w7h6LMGjsoB56DhovR5fjOw9Kxpx3xVRRVTo3fcgiSnudl8racc2gdyb
QP0ckHjdFIE7SxhimWBNjFu89YclT5OA88LTY9fGRmLvxu/FwMKzQRMbSiZI
xv1OuvLjMB92IOaVsy/W7oCROWU2dUVSDZp7VXPFhLHbNTb0yHYq2BRsZnJq
lfAkwiZ6dDw0HD63pWWmVXEf57554JwVdHAhknwg64YtPGYCl24b6DKhHvqV
IG0reBef+T00DEfNSUyJQuKUBQURzEyOZZHqLOzuoe871SsGlUqe+pcp+7me
t9eOVVdtLp2wc3UTNYkuaIsxtmeJYvPFdBJRRMZ4W17G22XvIAmCXfkraIDh
GlwG2l0sPJE20mjKtZ9PnMiM4Erb1VFXi+lxxAwAuZx04Wkt7SEybnltudoJ
mjAoQBTONAPIJTkdvHgOM7CauJHtMCTo1uB/qklY5p8egCVlUwV62OhFHcHr
wztX7kwAf5SCsKtUoJygH8couPc60JDPSqppTDcvgdF39Y5xap4wk2MSYXkH
cqEpqEixfYdCCkjnvmobKMvUw4weIVyiJbcwnIb0hJF4/yzDZWTc8VF9vNch
KKEZcKashgRBJlHjrNSDjemx+zHXML0KtG9JxAD9WhpMIkeNnKe519tqGTzr
wz14cIyziHgr9Lx+0eBVFgplUiQ02xwDTIoJGY3zqXSH9FHbLgwGqxHjT0o6
QhQ9tgcAskF9erBGlj4cm502q7JXcLWre9ef03fL18XPw8ECTidB2utaYwmH
9wydocWIfH+YdKxR8XYYb1Qrzddq5/UatoHrkuZtPGODxpRt6SV10iOQ9vqO
ez0TFCs2bvTCCGq+jZT2405dI3ft3KVt7wQnGWnPdbmr2mmCmqGfmrbgoryc
7qQyvHiVB07sebZsZYPU6sVcK4oNF6CAsTvPQeg0ikA7OiPrWvW0Gwtcf1rW
SoYI/U2It0CY8ZFlRzy9GS8muqQSegBSd+rDRrPz6P+Zh4HQtXqomlvED/tP
omMXHgJzSn+m0Accs9WcL2lvq4rhk0/rKXmx47IzGEumPQfOHfj0bIjDyLDk
JdnQp6SUnI/C1zqvS1D+UP3kcx7qZNf+okivprWuVzET0uTkgWd6NzF0vcSp
f9Yc9dj8bM8Kencl3fgy3yV+c+R/AkoSTPJNFnwD/5t6fpn4y+y0/S89FBab
DzE0GgYeiqNGHbCjrVTJp26AgRG5abswh8E7mknmYy1/h17kA3lgXbv+C8v7
eHQQ74j45RgOt5Ql3dzVVMZb9IrN8hpQ/ka+8XXzEGrsxqscZOtzjUn/NmyR
Cfji+ncOxHzV72PPIBqgIQJ8mTmfZmy54b5IntCVLhUROtp0pe5ViZoHMzbZ
OoOGW2TO4RLP8luny2EQED7Ink/1zm7kssr0KOYntuu3XoyuFxtSYWtS4vpA
DskzPzpX2It4aUFk9oFpV+macPa2QS+tYh9JMU9smd2OU16cpIzDjmtLnb6U
v/vrlCSO8hPCU9xcVygkkQrmlKBA5uMm+73FZ++/59E9Q1/PqpauQcFbsGv+
NQn2GbDTQYd8WYSRKFzwZYKE3wl/TGRlrut11+nlXrznRk1U6toEnd4fpdOA
KtwKNH8FzJEnjNiTK1NgQwB6K4SIbNDPQF9fxKJGE/rPolpfA9plfEAvrpz/
3HaT5PyXi0kTQCj+WHq/sdLcUf5c2BhRGc0a1s8xnlZrI0Vu7WGiDVWp+gCT
kbC2XuExFbaoSHb6OeWH3Y5T3WaygTjLLj1EDBrr3S7jXA9FSWL0GFVJH6c4
87ULouJOGwkm9ZMPOCuSD7acg8IGJn4jIOX/qTY46lp8iTjxmwlCQBFDVmuy
FNn8BGmMlKP4hd3oykkiqIbhKBcC3TBXtJV9zaJKr7kSJdnmb+KOq5RRXNDk
rsgfqquZQC4m5eXg0fQka+NaAqv4DxDzm7I1joUN7ZPMFt3pb8GzLYxXoe8t
i8ZIoxu98P3HatERYn8ADirC/XxjAmQoc9fCdPJaVo+ChSeUHNUccAdtTsi5
ugnyXt7Cl7T321DnREOQIco+GMacoLjIqouVs/pVmMUmS6/ZZ1OuYM1uh45u
jBB7yIHz4EOd8KiZbceP7coPpwzNoKr/K6/hr7h6uPKU3wuNKDbqRKdN1Ibg
k6koPa2tKA87TIbIfQe57YlvSBYEU/qBWDjPuM/t2rkNPkZg1AIRNFowhuGM
OlIEpr4mlBw/Oz1s2sSIHHBQ+K0Fc6htcQXrcPP7+I3OVXLYhOnUaEmNhXDJ
yNTZZ17lPEya6VnMN2lGUrKRcIT8WxY9v2vsXgFpi+MB4YYmfHFTmI7G6mRk
dxbXlDg8eGM0ef0G9j4ER8mdX88r3sO3DcHAgoFnmDGzmgLHMO4V5dFy+9LD
bJzzyulA10f0ipLxcsCyfMYimCz7drp7Af/aGIvYuolVk0k7Kgk3LVPwa85z
AudL3vvnLQD8dB9+FE6e476OZ/XmXxhyK+Kl9SrDv5SjsX79Rn0sUGkv+qHf
TzA2VTXdlNCF6UHefbcDfasVNIOOlyEMTddU3ZdDTokwkMnWV5GbLHvLTG23
IZsWR9H2IvFsCceVJKffiXEO8GMFE1JaWZk+vS7V0NC9iZgpnzYctYJI9NJ9
0dH4EL5shVqKVz+M7Lt6IUh4YxEN9oy4qx/S1N77E7GdKy8uOKmxnq/1gtDg
uNOAfpKcC8gYP0rY1mNVcTxVUF0TdxYyTnzWp1Aph9DhAeWbd03W3ph2c8p7
hEecQUUSJLxxZef04auOG5lxX2P7ucaHg6Q/lGi+5uNSfhLD3t6k9KBVQ6jO
Sa9ZrFtDr1zU1G4o9PhbLE+PqGcOu6bLV98waskoZZ+tyALk8d1e4Ye/Cc7y
kCc1LT2tsO0+hTSRI88erIExUbUIbDvreZ49bFMteKj+sdjZ/Qn7pEBduYkT
jdGzwQHw4SxWwJrLozybLRBOzDKLJrq54dQHHhr9GG9Z0+WEJfUenAY2o9AX
zF7iMRjfwHFau+foG2pbt6DrhTuVLSK0p3irSMS2j7CNW0683qfGWIZUd6IC
1ZdUh660Amgj5UEplZzF3ay+zyefXypA/Ljgj9Me3xzF45ZjSeURKsDKZqzd
TudwiP3IEgTFThy64YLEIKORQkTuVlvWZoVbve7lLJOi5916DyJ6qteClruU
8gs0+8JK+0EmF+5WpcBRkoSwsrhbxTVjzcMQ3241ib92mMDB5dkz9YRLhG5F
EDWBCpO+6hyOIrcSZUDvaTIoxcKTtkvdTviLBVJPCcpA4Q77HMrG303O1/k/
DlMGc38V27AelYjQxhXWQn4Oi7ctiG6K3SD8uYqpETHnfBx7mUH23CTaPxh7
kzPe2xdBbjCXOjXIpviagB3XmRoT6FM0Hfrm3Abl1JZOKksvGWikBXPe59V/
TBVAnzjbEFzb6qPkLK4oO4aB89vEbuugBCDX6ramZkhuQVsWxndoLXuDbFu+
ifEoGY+20UvLo7B2BOKHiqOKE0qPS8iebKXJLG95XQgVHKcbTGBQNXhNuMP5
xavhxuPUeTNJJ/5opRgFJsJ3knWSwSHpzXl75IKx/PUDR9FkqDY/T0SRPeu8
1HtSU3rAQgFGsdmJ8KJ4+qiQfKsZ3Kvm+4nreKCWDwSC9qS0fM0Sl+3eeIuI
kTX90Yko07/2Q48MJLj1R6zuSqsc3lvTjhx9POa3r8Qj8IofSQyfKTftfDL9
dQ7wBghFVKSZFc38EhNmzFaScyQ6poXqKyt4p9a9lclGNRtHGpZtUN3dsD3T
WiO7qJetqCuQL03NC2moWOb7u5jzAclTP8xQWz8P1fyp3pRYccEmiOz7rqkD
mQGlB3rbEXroIPNZbnyBnQDUA4iDtPl+e570vXnxJiVRmi5ddBCADG/B4wzf
s/lOVJhmKDkR+esTOUJashBvpr+supdCI0Tn1rdZU95nzFqcS8vLAgAvi4QY
9mWieoIQ+fLOJC/G+YfIPWvt3QTvcheVATBJ3rtk8dVBkGH6Bx/PaAfgCBnj
ZNMS38+HjHl/aoXcn2qgKsHzrTtRo/zByNKzw6GoGpnsVSaiey0VV1UDzwx9
+IQvQiGPkwWuIzGCBfSyGxJxV0SRmDjEeBjDkhKDK7at2+NXPEA7Fq2bvnmj
YZM/RFBQZCWKLDKrtn90Dv7l7U63gR7vst/E9Edc2bOcwJEGG938rZEqoZru
78TAl9x8plAgeq5a15j1WgusxADv0W5slYHNg2KLUfhti/asHgoeyMS/3c+H
6k38/zeaaZW8xTWIP7N9MVGOEm/E8YnYGcpaUSyFrRtoQNtIllV4v5cIO0/X
aHmyw4F6628KUKmiML6CIiZF9iR+DeXuVroE3zgP1Odqt2QDUe9udM9ybcW9
bxCn44u/LWL4jjV48SWLMYCPPcOQOh7zyf6g9KmA+HgZAmMhxmW7yhr73/6t
E63rWVhdQ0jm23aGemjwKHy133V8QT5i7c43lfdfBSWwGOk/cY1s7f+9xIhb
Kekg1B79UL/E4AeBbljlzuoVNsY+Bj6nLF9XPkoRIGDBE9doCzCu2cfDENcJ
YZaRLrN7nTGcsAmU4lI1WjEEJGvEaAext0dvp15Nfi3/84ZQsAMI0Zdw0zx9
hTfdi98Ap37fMamGCscauzADTiieou8eF0LBOKi8Tvjf9htkJWrLgWjeRUsS
MFD+lrtC6WwZ8eF9ToBsGs2gAsAZQDSOc42E/mcZedwkImKb6yn+7E8C0E44
YetHaNTMbMVFl9uQXvpe3SAHTOsyAo2j7f+jRq54VsVnP5/fqrUdfvF+yHcK
RKZg43hv8XcibwqA+57on5NjPtD3IH2sjY83UVgsLA6mUcMyl8dlvijiguXz
VJg0boyleG2OPvfdAmGfmPt5wGXHdEZtEx/rCxmlcvdMVWCCweU5TBBie/A8
sPRJGKaFM8fxO3TcRLmszaospu9xhU9X0F8iEOTJdTBp3NbuvrSKFEHcDDsy
RTbUb1SezhZ7xUa5/I+7HPbRJ6e+LdmqZj+4VZK2jbpgHP9lvfnSu7pggzob
8fs3DscyafLQdFKF/GOsWZ7mVuvP50LL+bXpt19yX2hLtFquL7n1Y9O662FG
3HrCXiE+jKo4dZmLHPQpfwsLyoU9SHSW70YdaTmiDC/8BE7ySU5NDcMg9+C5
q/1z9LEO8VsbOiycKypDrCW4ui19gAeHdpxp66IpDICCp0EdmI1oZvkm7yB8
9YQXjpWOBcJVJzvWLchHrHvIZ03YT+B9JCai4l6nMhjSVHzjaNTXdhbROsi0
5l5iaiSZpP+as1hvy9wYCwkrwF3+PMndwBkZJHQLVHe+zEmF7Xf61k8mGnr4
JYdIAg/38IsGUQijPRZjOxq/MOKn4Cjma0fZL0LIu9PhcmHLHJBsEQhl0IIs
Z/ny6qJOcLiyzGYP/BQxPQv08iqiNYSQ9/GAC2osgXboHRn29B3/+a3s3zP+
BbMofwaX3I2GcL3ufvUK3TR+W422s7XiAhZPCgDVh5Cidfa8xqT8IQnFLeiE
pAbEWpi45564o7ZnRb5IIGXbKwRABR5rUU9acZXhTmCpx07wJxPBkDUzi8la
l5Mey7WOGzdhRE2CAg0b/340JAbgeikEGVwvYUjGWDcXYw/X8Sq49xAQUsgP
I2WxUc06dSU9en7A7r9vaTH6m4+UqkRzWvPVkMZq2Qa6RousH7bvBdseowe7
U0M3A7SNESeYkx0KLoK6lJ6Co5FfWBtUD7vXjht6/90MO1poW535xYm/2Qvl
03mb+NRMluKp2sd90skWHjuMiTgRE5eImTgxlh5oMlMU0A3Em/YGX70GlX0S
GQiQRraX2jVOjvvCoPIZh3OgmKKovLB/vV6hrJSoZwee0lMIuPi1IL9l3CVM
RJKOCMRAtBPPh3tzCpBp1q3occAygNOzi7/fXuEE86eCHEQR5EOVXDgNR0Hn
ClSlhsLAjqqV9HtgK3caz97hnusaQzJaWHiqySh6yimG3nCERcJYVQTfd9mS
w8p+uTMLk48S6DuATOGSXFvHdLTzjRt6MGJmNhYla3XJsqCsrwb41gadTInN
azK/ly6eVNfp3gR6IUBhETJavT9kV3V5mye9FmFVhTwWR6ZuBLkrApwj0de2
8LuUZmhxeOtcTmBQ908xp6XNTkFAshZrdHRr0K9q8SKl19TN7f9cZBPVmOE5
CKyeon3lcvfiTiOhRThGDuqpt2i9w/63mpmjK4aS9MHX7FfCblWvkrgOkou8
V/c0FoVyUQ0GymdtiffUPVH7pjD4ek5hMRGqUsyhLbTYyKTjsXEMNpu4FEQY
sLZ3a61hVRFR/7w3f4AuLqpil2PNqenhrkW5qSxWD2OmMAmJavumGUMZYkym
qVfNTRw5u7xkzrDQA5n84K5n50xpLRBmI+CHxnrv0SQhhAnun/j6SUMSqoY5
Nx+f60wwPkW0bwyk9aqK86dITmunyAXJDQ6RWD55mKvnu+n/uTHd6eV23ei4
+tlLE376ZuuDzhOMqmCA6qdYO5sfZ3c+cXyrCQeK/3KihtG43+AKQIDUlefV
qWC5BQKu1ihM6YzWrrL4KzvGu88i2CNJ6tLmAutKD8fc7/f+vHG47xZ4LXUS
x1dfyHhBL6V2tYacQ8z9LbeKi665ILvMyvpUL+6taxkjLgi5iW+XopfT53T3
Z/87st8uBz74Y/y+/9F7gdwAwWZdwkOTeKqtCWkK4k3U1HdUhlIC/XC7DO+N
9DWNI5WvyrWvWPyhKqKvSFOkXftETVkJX34AOr8VCYc0v5qGLw6b6MiRhR0I
49pWgXxdomLkzldI8qvksk95IyZBSuaBFHAZ8Gk0hP+zMmbpU9A6aqviEVbO
aOJg9Av7m9JtCT5TIvi5Ehm0dXdDHJjbhgF3oeRsJZX7CaxQANRmoWbawziz
d0+1A2d6sansmZ44PBUrjUv/crfHNKI4i1bUg+KGt/hx6UyjoSw+p2XIZifD
vQgwDkiITt+kZzmsqBHC8GDGnOlWpk9NF4ncXA13OTwpGjVUlcp+XUsyc278
TqvqaolJNFM8zwuC63+HuNdlhhTTBSJTvDOWxF2JATpeBPdeeP7P+asIgDwv
Rz6HF9kaHI4mvuHzw+dYKaUxPtP9SSHGDCdO+Ecf89C3rd7DeyHecMC/ccc6
9JhYNbX8lHiT10pOX9rwv9wh/OO5gC7LUYd0RF/9DgrcAvW7nEbveTRDaUCs
iCq32JpbxrEP7dSLn8vUeZ+3N0RzlMv5roF6gUYgy6uoI86vlDSwqEHwGPUz
9qomvWMTLELhUHDBLD1kT0DLq0HKZglJztsQ35MpwW75IlkYJ6F4hhC7+dNb
5gsczxEV64CdNxvvmYsYSAbMOl/UwMezxfCN0g/Awy22FgZq7CYoPSBi92BH
PxMNRAQVbI+5hi2V0+bHamORY2j8QD/12cYQRPJXNMbAtbVu4ymwcpxDxegf
qfPhh7P/l5buIDkthTddPUgAC5afnt9ChVf3RkQ15iz5NVjzZQP7LVpwWuCA
FZmL0oeZ06dGyeuvPCmWNIRwpD/7AM/6FoeTOaVMCZsZmiyuLkF4pdQG3DJ4
F1cUg6gkBB06nj1JsS0VuHHm1Rs9IwyOFHpYCK8xAf0V8T/hJPCywk1KYgG/
Pz/LMCXa1Wmi4aqo8CGh4hjBggIoMytfUC9c7n2e3asjsb9vcGaTM+Qmerx0
wenOZjxwyBBZ7V3bwfehCAggFwgOy56RcoZLb+powXL//9gAIGuGZErMzt1m
lYbPnwLbh/vVJaThWBa6Q/vn591VcdBdC4W9t38hVGCCKElV1hJ2wrIjX+aa
TSj0uKlJUEUGnWYTq1nI7KL5/u+doEIw65er9G35CL0Rh7K5r5pjrOIx06k2
BShaVc9b2q+U0zOOtA3fmuNC0HGlR2iEDFT5aeLqpfvRM66wMW5weOMBWah1
GAtqhy3MPltckAHPPCOQ4YbVn6t5XdwZQW65948ZdZB6b3+uNsFj8KGLS08v
FHEeQKtoCI21+3zxBpzJY5dfB5PCJrjWhKXrsuTQQgqAu6RSxzbtAEZu8Zze
3P9Yw6br87pdUuB4ICSQ+tL6AyMQ5FVU4L4b8xaUvObkVCrJXmwJP5OLV8H6
WwNR9nmv+FrmKkBaBOprFtgxVgsDDzMWPRVo3LdQzAVcmGpfgBq4u3yZd7W/
ObCQSyJWYFRg7mDadJ+BBff+6gOQ8kpLxCRxvoUQJo4y9/cZjveqbUvCzAUI
B2e0i6AsKxVbH3pTpCjjSPtPp4zRa70G27e4tbudbkVIzBonrpXJYl+Ygjxz
7SbnKUDlQQz/9Mv1YJXwMOnJZXfp+gLwcS20salIqupk6pVP1/yNuibxO+b3
EwvzQOlI3SIiZd+V4Ntfo3HdHC94h1f99ndKJx6H5dR4ey+kRyCm/2G6aBTW
t4Kt12K9jv/qMD06EcBk4usrdPPO+NgHhOqh7sSazaluibuvUDRk7Q64RmaZ
jKl5KXiBbbcu9ISjXK8mzYLonIn/uJF65gkGqeIkgR7ixdmJfUIjpWrB9zVj
LJl5ukKWA4pw61leAlEFlZdiJFrUG9XjiGpaeXTEi/xUymvD63AdhbARMT1m
GYQcAFMoet1Bl69UpJpT1dhPS+w2IRmzp88fT3/go36qhDBuvrmyRiTMOAo9
F31kyS3NXrb1of/oK9kLxHglYSVN7skqE7IXOvxHsT5dSOUJ212Cmc0JU+gb
sPWfAs0BA1+a1qgZo7OVftzholR8/rcMVCBGfKULMovqPSvmrgOHNQM2ODqa
broMtCG3qs1/gC74KIGMnpsJ70x6IwCyMRzJ4gxSG+eYrMZYCpZSRyr1t9rd
MvnR0h2uztVq8wqG51R5RZHilmIfQHW8e+Pph0iKk/OhYJgNpM3O5+dvU6xu
dV86ub02/3yy73ERqtPdfHnH0ujc9h+mss1t+j27ihnaE3rUosNEhOmgqHYQ
2hbEGUnsYeQRNCkyX1lUOWvKXuSVn0Pd8d91GqroNnXZInSa9uU7nnoX5UeK
DzUYs/RXvkhkNScikf3eaQhIx6hMuoGdbPE//wUEzdE5LK6PY0XilvgybiYo
aj9RXOY88xPfxAjFUjECjw0MkE3+GA1J1ZzFl3azTJgZTyQto7d8ZYBmF6yF
NpZ8RdrD4cVHdCievxnbRjLScTIlmtZDvPc2vP6zPOSzFcAz9LmkD4IlIgBq
rAI83psqlnFm+b/Yl5D4lSKYt5Qzz/Wl/YHLmJxsB178kieY2KaU938PjptZ
1cf6WYY4MK2j0NRKfxV7lGk4LRc6NVM9Mz2eBNIRd46zZTvZ0xq31NatLlZ5
H9zai/HGMqrfVJ5FIM/UECbOQU6y23vAyJtG4rDViUcO9V7BFSXgCreWGvcN
hyRmW/i7R2tWC4d0JYm6Oxh1nl5vd+oPqy1z0xOujb1QJP6NI1pMviTEjo4A
WaLLkD4qat1wWcluRYmlWzUz56zeHRnxGHIslGHnSbX5Kj24AWdJyPIHAsXU
Yu5+xGBYxadXeCaCEAeYcwrm3jAWpXe0Kt1p2nu8dagplCZXc2+DDAWtgcmL
++dwG62mg8zRe2/UPXR9lm6G41CYHbfXKMTHRl/koFYkJwRqF2lNGVrMT0vW
yfVG2bhaP+PJueX6kYYyATJ0oGEQ/lmcxh+TnC/Otyd1Q7yaEKVm7wM4xIUN
EYJmJ0TPdhD1ymgKskeBhZzEvuaWlzg1d/aKCELDvWFAsWIaQqHqdfi/NuDc
g+cbmpnJmhg1qNRiah95zKExKx+K4UO19hOy/5iF9dgl3sq16vkdjLACTNn3
y8ljg8/1ow7X3oUpzhjLBAx0j/HsIKgdAKGSBreK4ltloNYSQwnycxu4095I
R3l1POvkESk05eNzyHd2eaSxJ+NWLWoMiYATG8Kh9UQh9hd+AQJX0QJffcOI
7Re0861H2KzSQriFwI5cYVUKE/5p0SQjbpZA/fTldVZSjtPvc22x9eJ4yBuU
OtKFcD2pjyEkv/ShX895V8tje80Ef2fZ7TDLZ+pUd3VSB0vzCcFUOn61NdFg
sOdD+WtOu7CiiS7xCYdNK8hBuERjT3AEq+LDZz5eIxorvbMEc73URtgL9MyU
EMIDfWyDC7TIWZC5OeSGZ7VS7H19O9cfEWHuGmlo85RXUofiB3EdEIsGXKBl
XYvnINtRkS5KD1ewrxVs4erVgfcKb/MDk13QsAVzCkpPxD2CxbElDN7V4D9Z
XIg4SzCfZ9fTm+pOCGIenp7ewbtgbe0sDoaWyKKAyXyJiS+nE8LWvbtQQQqk
WmNbhwtbG8qZCWo4pz8Q7rEu92jyUkzdyr0LQLoYok2vj591g1BRKvTHndzQ
zAkun1CtWQ3maNcFmcZQc5WmHPWeivKyo83uarrQrEBDm/klXnVjgDrD4gfe
V0pbRpB2l+60G5jklYQ1lxPX3KjBpRvTAA7DZqsly8tcYGwftyd8cq4Oumbm
tZvwBPj3bZek2T8zIuoSyL+Rb2LEOhwcCOaMZjmC/LJflPB/O0s2RD+8IUmq
7Zwdv+0gBE4hnQvs3J5bjpdmtcAi7x9PhXuHCFZVn27WUNyu5xx9REaKEueA
uDyMSkdXSV0W4jJQVsOBGzOzlQ3vDBjRFo/oq2iInt9i8iPftCHhT/Sx89Gs
o6MXhdVlP3kAg9wGmTxq5vMbf23XiWb/EN9BecyCX1mDp4TliMEqTQuq5+O9
im12y8Lbgv8qnYKPvi7Nf5j0yPcLNRb1kpsd8KmbHZ4uun4+dI5QQWmdufOv
wUR//KZtXC9yW28bnexloZ/ueevU0gM5QAJGEmXAXTTQrYOpx8uxoiSaGVUu
Rn2NqQBpePbCqe8Qsdr0QgoDSbnX+Agh+LCfgrn0f56zNmTpW/IU6KNLm65u
D7iaEWD8p25rnZ9TlVsf/BOXXof40Ee7+ExC/L5dtrNfFaKZbvby3sbtyhup
OoE21RQGSjMO+0/8syBSGpSeFf34h+nGc/m2ryIN8gsNc3t0MhgQyVkR9lvq
W/QNE4gFZ6btiGo5oCiKuow2t+nml68BmeIm+ckDtykaZERnkE8yL3mUZ5Ss
6hhoKz6FdcfHB2Bl6c0iqPf+IxD59IrGuBKdDTZxL2Bn94V2gnH0jyrzrz6r
WrHNrmYMNREBcrMI7GqnrCqydGANkPG8uwf63BQsjiXX4zIVlVtJL0jsAN5D
YTzkvTdMsQlSU/Tn/gbri4GAmbFigurqkidcKjc284ZrKWcKqLOpXRi7rT9D
kuJXVSt5SZnpghR+5pCDCFJgN2RG4Oxjayf5e3SmIRZ3HUrIFXJ4BwbUPiIg
EtKeEK90XELdd4Bo6HutjgzuJDk1JQo/s7sqih61Xg2uUepqIkFVuvyvnMbE
Uy+hmA+aF2eSFSnN4L7577zbMbEiVzCcgOWUlDHgNN2tp6x50vF4HaxlHzcD
OqUkuOnWONwjRaDiG5zI9cnYX2LbsfBTCZ/o340C10jRWYOgrns48mZVQVh+
gscsHo6wWC+qSjS/iALoiyeiNiPFyjQlSd9CRTu1NC2/yk55iuQTlq1bsIOL
cBxcpeFf+55kKLiZNutVd6xZ9Zn8idip1rrYA9xNnxbLMaRmmzql+Uf+gF13
xHci/r/e04Oi9SifU2nJ9ehyhMlXeHNeDz7MmZzv6XCqoTBiyxZ+gBKoi4Gp
/VtqU52HIy4k05oygycMmRQhjNX9wy4est8+1nz2JBEQ3WnlLQOkF4SYCSuo
Yx9w7Jh4/WaLxSbyKMTxvrzykX4JBgtAAz2SNUpayaf38DLYniUTBuoSc3UP
Sw4WBs0hEDIqWsBa/i7W7HwHre/Xz4NisYo+2JYPIY2U48jHHYCWhrwLn/AF
mm2D0w2uuWM/yeO7+jlyxKv+glv/bJxA+z028qkcz06b8wmEav5HKE32IJ1u
8xmfeviOs9gSWPspWnEcGlfw1m0PyUGOkpHt6oM2kdFhY9XC44wenqaLtRQ6
VjTOp3Z01OuTIf28YUYAdfYXUM3/DckhOIw/hCmSIhLeE7qZTTw36sDW+SP5
sypeUS6Ip2bM4fDZB2ro7nEvjFsxjIN72RWvv8JDJGurepAY+wQod1OHIibR
eUkHQFpwTIaOOQaNdz7AT07c9JQ1jk7fK6lABhcVu36SudSbUE4bGclJ+xFq
S6vFg/gLRRlw3UO244f40CM0+fjqN9uYOvMovDRP9kI+n1nYjQcwurYvXKjz
ri/tg1V+vDfNH2wnS3HTX9K5qm2qxp4t28iiE7JMT0wZwlB613ex07GPzOU5
ynVHgzyuh/4OdSNLeOHbm1ZhWFLPd83xIf410+ka1Um7BFjSrtE/NRMBtjTH
mYtnIYHlNOO/05rKei27u1EGJ8toTyDnaOn5SUy79TCeXWNdsQePB6kDuXuY
CKm18PE292MfHgRX4iYRtY4BEkcWLWbEck0qTlPc3vO/JAIH47I+shPdhwGw
mbwb1yGEEzVZ1fPMRt7hsjsTjziEnU8g8r+c7rgMRe17Rfo9NWO1/XggjbBY
mFqXzkrfMX/q7IS/uNViG4TJKNkC4BzWndpHpB92sdk835zPbveCmjTVA1BI
16Zf7cuYaATeibhKjdGFNwtt6R8c1gi9U4s1D91aM1lcNWPXlqZ9ET/Vkmdt
VE1Oq2+MX1Q23W8smZTDBmS0O8L1LVn398sEeTmwiHMIBVpFhJQFFnDaLlwK
P4qMd0powBDYfhDV/KETh/5ClKjOTDh95f3W06uj8LBxsfkYjWNe6k/5/TRk
i5EKlCp+tIv2/ypqSpPKdh7SjXKo0VBfBSWv4hT1rSD/2pCvChOAAWmOx65N
jNt5o86M5AYsFM4qqmvMYFf26Xj+fz68/UsvA4K0YprX9p+PySbf68yTLwGb
+xJal3S6mXm/Fx1gLgsi3kIRWhT7p6zfGLu4VHLsjJRQJMKCWlHmrbrgbhn9
ntjj11HL839m9Ab4CWH5QYeU4lA1RRLNxDr2jL0Z73FrDw2Y87zSdszGI8yZ
8pajWdHEiJxf/CF1yo4IHyha19jIT4Ey//MOyQZB9QJTgCsqCU3oUGIBQLd4
axwd5AbD2uw26sNcD+cdaN4FpKQrFKoPZVrEn48iea/ZrsE0Dx9CmbB9Qxgu
Gciu9hFWbuYgHGDqQQslz/gQRoao8Pnfw+qnDinKoV27vEwtUIUkrZNspmjq
59celJzYYHWI6a2e932greGjMkXiCbhY+azspKEQi+Xa3QZ4s1DYpBsApz7P
5GAJSbZcUxKoTc7PdFrwtRIwk9YLt+8NnoOGjuHCtmIuxlOkQwlcsqhVDhJb
oN//1ZX4wEYnRXpH9jmJXISzdVUP1TMletJ9Bp+pmGdXlggyN2R+1ZEsLt+j
ANwJFsYZdlPsd+VtI9/G9fqRFcuWASmOL2464IhCaN5m77x2lWj4qIXNl9xV
ZHITzl0wpiWJd6RVkBftPkmtv01VnYjT+S5vhH/KQrdAEtgmRfNqjph149SM
c+abM98H6g7xPLbdZ5fMd3HyBS0F3AT9YT4GhghXJLpt31vX9o/IziNkCLJ4
38kZBnX2G+e6EzjUUmx60fz5ACKEKJddFM817w7rPRMbqeJAZ2r3uPukjgQB
V1PaeYSYFQbYWaJ8w25NUQvZ2jmUEuyFafqZfJ4M9EY6iOKdQOC+dVXPn4tJ
PQP73fFg4IO5sCvm+LqrcqY9Tqlcz1enfqDnVfhQrzE63Zk96UBPKYlE4Efs
CpP3q/R6jahPzAC8XsTRMnepcI2oLjkWN9dq25mG+1rR1nwEu4j6xPGo0OWG
r9Gl/X82NLrNg6KlkGn74LgvMYbGwduo94IgsiXjd5Gr2LZFdNDzgMBZYY4S
FCXWFbn7b7yZYoQx0qbhSkEZu3FTDTpCKK7H6QmV3md0WbGZkmAbb3S1UPdL
Lq7TW3oT4fGb7gz2Qzrn1hrF3/yEWPtqtvo6c1vBwHaqUwm5/4bbh5mM+9zA
Wv0zTV9MpLEYHNcoOw9NT0TmylBs2G1PtVecV4LyoYal2bNNv+JX+8g63ZY/
X0bmHfoxy8tYOBa5+5M82e7FVLssCMn39MFwPy+ZFupUoG/QG17MllziXmt0
pCRehtP4IoVc5yUAezNRAlVR8hv5OE8cG8lcqwQD9IOdZbgpfUvNQnbvz5a4
WPQ46m21EuNGo5hAXqQpCDkId52KBLnV39avrLfTsyU8v/vLCeh0XHiN8SAQ
f8cqikmLmH5OZfcKunB9g431klSqTqjtYpLqgLxAQb+Gqskn/xwhglk+R8Nd
m45+cV4nfVPkjjI3te2gVaxZSXrpAcOe1Vz32hsRFI2/3AcSZ2yB7PDfVsUW
qSyifV/17gAWNMrYPY2fQYSrnv35uEyqOA6ISQwSF70/6pe/R8AkPTJlsCWz
H5fMLT7pLa7xipBGfbwTM2DXqxapM39Tnzlw6U0k1J5HswxwkKck375X12QS
nDx9hS/o1b+mF/1ahotsvxnBFWWCMGNO+nKih3iMibaK+r6/HI+idPqYxTme
ja2Bl1enNzRcHqi4pKG8XCYR0nWok65UpbaTuX7uAM/s9N7cpP0iQ3F1tPFn
JxWmT41+CQJvvHLmRnZck1sVAEOAXDRDQlDLWFuN3DGnucwrvM7s4LKqMnI/
anSNweQPAy1w+rHcQd08oE1epH0D9tRmnE2cb4wPKkJHtMoNrqKoj9a1+TFo
ALKGCxQwiR1WqutjJkffPrCyuErqOP+Z75vxizwJU6PmJY3NLG6AGuAkzPoh
ssypQZarw8phkf9CLhhUYgM1h+yCTTB9QHE0IvO/YPacE4W4TCAhSPGctuaS
Fpic2WiF0HG/LRJ0dHFto6FcXg8UsVcN9b5J3Y90mgepOPxKpW/BEc/52YBt
aWciTJKSQE3HK8cUwG/Ayxs2Xj+ofqDagJ6BHAhyBLrQn3PL7PItvAlUSvja
ikK8wMrpVJcv7CrEjl5OfkGv1VswRmAm80mm8yQHQnWiIeAkE5/h2/7MV4Pk
A3oYLKk8FxpMlEVe+hyOy18Ol8EvJcIYA4oPjqKrBrF540PTW+/HISk0TrBW
s/E5VHk54PJltR+PtTWws9GG9uPiKpICT9h5vdv/dv9QQDK43ul214GvbmQ6
d+WUtXhfZb7JdEM6J3XaUrNJgBddhlQFewshGX47BjGoOX389WqCnPOBM75O
360paRU6L0qMuqrEcA0zrMZcUWPUni3MZqxVlEiWD+vAWV7jiuuXdJ/uI3zn
jcZp4CbhppPfY3YaMyJ7xK5RGg8sTWv/UxZ5s5m8PXRGTEzAaHMGNjbzMMTo
6Mv9jjdc8HcgDbri+cnCRKQv79ZNT6SyNrmI+ZOAFZN7AoXk38mu5jKRWP7g
qTXZQ6a6mbql+FLwydFn0n1eAt+y+tOgJa7JzSRQfLFI7G0PXfosvrdA5qoy
z+EOGaR705xFw5lMbWO+NNvLjygVnR0IkRvLZX/L4zRbR19282P2LyxoTEEL
RuxpXx1UQc/Y26RPEPosriz1+iA3RbGQXL4KIbCkgY63dw0fEJr7IJkpryWp
V4kFrXLdiB/CfJYXL+F9PlqTmmK9bjwofw+z84ARCSzRK0mV01JDxKWZcaeu
2BZU+8WgJW8WODUdvdx40tIciAcJAZLlkWzOnQLxMOmsK2MAdY4UIP6juVg1
NBZl7ycjxcrcKCmV7S3dGViAPrXoICNygrziqv+YPyxu3VLSXirM3dzpmX4f
ZmRXmM/1yt3RZbECvVD8XyKnPtQJx4WQv04dqc6pZEKIhQCZC2HZ1a844wvq
xbjRcnLTjp3pUa8IHGfDVwaXHQflVs2gwur9UdaRbAR0il5MzRLnmGPsnR+Q
EoBf992GFjw4R2ObsVO5uCpbvW1G1A6lYsVxWIvBsvB448nn34A5tsaIQCXM
mLZ3nSO4Zt6DdBlVdYC282HhCUmbMhTWaAjC0YhYXf0SVRFxtxZIvDZM8GLx
/QCX1ts+qzXJjY89DTowFPneX2Fj+wTwNW/c+piNPAs+F2kVHducOYNZE9GC
YXPRkZBiyhC6JIBCNd3y1t34sARual98aerLFmYoSk1YZaxea49q3hbwnUIn
V5huaxEwwdgwaWE/2NPZcJmDap5hVmr64lg5R3zzvqDygldTR46zaXuSeHoY
ZUluMKlXhfPRLTYhQXK8UQnEVfaZOzQi6YhCoWUNiUxCVA7M3yGVZbIpDD4Z
MUe4LU/SAKwdE8HPVuPEq1UD1cBxPXH//cu6E7O2YvezbqsZySxOGTfDpgzX
pmCEQiA0LfOV6TcPI9Fop5G3b3OkSgwdZsdgyiIwQWyNHewWg7E/sZ2WTrJG
GXKbmUAunLUc+VLwj3+gED4gwEQoBrgCDWiFDkMDndv/YLE9xap4vxveyMJ7
Gn/lvqW/RnQS8UV/JtwIx9Bq7Q99Xnb7sqTVemggN82+tkXZXW7UEPWoHd+E
U8CQeWPL1Jv2GngtrQw0qTTfosLUp8RH4NTZSkxpDbLX2a0uoYWkxVKUmY/X
XYGRQp2BqJaJI8mDKzgtDXUYvsd9t5A22OJmE7ILrWlTFoqrTunrZnDWLsXE
roU8WpxOpVTvkOQT64fdb6TZmh7dwnhlh3tNv6onB3bliV+LilCiDMtZn+2+
lrNhQbh98qGiUVt+YjWkzUbN+ncbzLHpkv7Fc+I56ED/KLABgqGyXB4v4+iA
8KAGQ9M1PiumV1KqSfSJ8Z0jK2R8v7Q6LhDZDIEyYWLBoq4nUoZCqso0pl8N
wcZSiaVUUFeJPApuMEBSdP2eAo+VIFJn3TlhABpsFjCTxpk9r0mqNq5lRums
fCTr2jcTuiEBzNjSKSYaDnGNHl3rfKoLkPxpHDTqoC7ez4GDBMlxcItfGw+5
cO9gHwpdwFxT5cFQ2hhwWoPh7Et4rnPOnl4gghVERJN0cVMKujJ2Li2NwVLh
+sNPecQFzf0T7STaU+tiMuaRY+kljcDsd06YMoy6wTkBMJquGlQ/giLf0+yh
FaCDl9N/NAqz+XO9jOZW5nlXxJP8Nn8OhSdpdNvBD+85up+q+QoQj2bOyhFy
Nx2mHhjdKZwSROH8LzS117cEJDMIY2Kfq/uFChbMznQ8Aw6YB+TspXPUUJFS
DY17/uL9N/j8kIUqlHTHUTw+iGvUrdISuwixr3d0PU/4UC9QACVFNhN0xyIE
qucYPy3Goaq9MDajmj1YCMPkkYsAy7gmq0MQvE+rMQ7orQCTFzcx3ZLKiIn5
lv7B9Ef8ZnEW4qcx/pjO2SGib3eBO2i+igFEJUmOz8uwBjCVQfSZ5G3kB8MA
UvjpQgc6LnvI2s/GEgySE41qWd2MlZvN0FIUNDjy5MkeDXD5++Clu+NIsmEk
oA6h3+7eXsxfZr6JpTJN37KlH+CLtCjjkALBjRVZgF20IC9iKcQbgTPZiQ8a
hGqNYJhwa1GJq8npcibdxatUB35c19R9FufvH51xFdjIkv86iFpM4lqPMa5b
m/ko9RzfPHCvXxk3jkF8VmcR7QnLN8jtkz0t+vQ2QKMLUFZFcrVTUuKU+Gxj
4zL7fjJWKL7BlxAc9xqf9Jput9JGPZFKYQzRvwmxqeTSfZF9c2ddFoofs3rh
LU05BL07ZElSGg9+Q0UKmcrc4quJSBKK9TVGY/t3yxUiwvPdpd3YsIX4EwV7
rZwYxFfOUpvrwFjpWWlO6ohRWGusn2ypKabZI7LuDcrgvwACOQBOIdTlLWpU
7fT50olcK0p6QeU8jGtgJm3UhSxIogZyfTca3mK3H6QulC9suiRukHYo82rF
1WCV1stBfmtiLzlZM94tKn64udflbE9EDT6QDt+Dxq9UqouJuPg4KlqJVsW0
knCzB6nOdXK/VphbV5Pn049rT+cSJP1TiroRO7hISTJulyC9HamHYvtDqEId
iFbCk1TuHnIUUt/Y9wrF82/GpbtborxwkIJsUoitfHdiv6LORL5qS4dqKfO1
2divTkpKQX0/cbnCAQ4nCUC/8S54Yl/d8vIWnhN1TvYKoXJxmVR4TfzvBVnG
+wCNlJPNIqsXORZBIPZvuuf+TMWJCMQgryMVJK32w5L6+GgqjpGM5+EhEelx
yTZ8yE+nTZiLTxlVkzqEyUfuKIZF65ttfxO4TeV0V+PZqzEMN3Xrbcf/XWrI
aKG7GCTl/IL+Pl/Jan1GMB4SGoMgbcNZAlrOMrl6AaTVM7JcvsLSXhkKhpmj
jzJ/dOX0QYgRb284GhGQQFcL/UtwPO0Jd0/MzfSyFwph05OBJuLOqsnHzs0g
GIjEG9EuAvpPIunf6s1c1MLM/wT7v/FArDIl2Tsqhnf2jT9/dUVsPyRVRv+3
sbKlki4yGz0wEXXDdhsL4XNdhIDYFMYpxdpe334dPGR5VX/kBy9bIPin86Vu
ABl+59uuU7ewG44VSKYOOS7TjLF6TFoc9ZWXiIzbQvvtmuCSp14VueOfn712
J0dft0pivK7AD3hOVR2OkbJfXUcwaY2T/S+LYkHGJQnUOkWS0QMEqMR3f2H0
c89kVM7CY0IWTr/m2e8EUVl2jwrnn+COxxOtkqdjY8xST0GJ6sFpnKTKcVnb
QzRs6AR0aPMqZ/9+SV1lExpxP6aJVwU5jupfHWnEpQBArEKlv8xeEU3C7fbR
5NTJ0iK8WgQsHOlOsz7Mlomk47S/HAD9m1Z5AUz54Rh958ZLeJTQ2fppulyI
T8whzxcU18fKrfq40NOVqKzqG/PjFYyQnDICPUpeX5pw/gKvKY4J2/GBovS2
HXUCNK7/p6PX3JV0HErwd5yTYDEAW6XJtX2y/ayVIh8N//p8LjNv8Ml6tdRa
UdAreTRm8yXZ0huizuWhU9Y2xZLjfk0dqnenyzKMc8qo1CruycafwqQBN4Se
9A2x0BSFzr4nPf8+8N/1j+7sKHmN8MOcdrw2Z3wTy98Inv1abCccyJPQqviD
ousipouNK5WRomv2K9g7w34AUjsivRV3kVFFwbYQSBjOwdjZUrVpvFK4CeON
PrpKQXHirlupr+AjK7oh/WWN2cIevMGJne3RF2hWyl17vOCYw1sgtXtdrGiF
8VM94YGnV8PImzuS7yL8kQnx+IjfWPfDixsAWpGb+AH1dQkpWfwf+U7Qwm+E
0xiHorNjNLpAxmDEA0PpzO0u7kW+7a++M7tIo65ZnJCFqRDiHjlAIhJUhGNm
v1QTMV1TX3WGeZYpAGG8NwH2tnURGs0ShX6eO2b3xUy54GauHKM0u9uT6rOS
SWkm+JJTN8KDiJpiixol2GnswXrIFYawx/VEsCu2dr0onwA272s1AnnVd7uR
R97Ek+GLvvmqXdijSH/T6i4x1IfDI6IefCb4mFAkFbaerwuqt9UlXdpXzQD5
Sd3LD+7bAyKeu7v5RczG7VtXM6NG4ePKoKDLqR/6vyTvSvv8NP5oSF9QZFwo
Z8qNdkAja5rKZK5Okkc44q1XTda5VZ5uXBTn5+T1AI4YtAMNe49P+vMvR6Aa
DcfHf/SU62EpdhY0Kiy/VlHv5CMbPJnBEH4J/4XtJ8eHlWLO8fCcxet1+IWu
Sudj6ALVqy0Uyw1yrABqkPpIzlAXIcfXXsihas6YoK1STEQ8H5C6B8+r+6aR
1tNMX57MxiLTj5YIaeWJSaQkS5kq9l45L3BU5flJCLkom5SVTwkDJKtdc+d3
tVGM8HhQ+wzsfrElnBRmdT/Cex9JGWdZV2+EfJRbE9WTv2KT3wZ1Br7xnBTB
3rZzXcM4xGE72k00NPGE6G8Oj/jmmQYAqNfD2apkCzgjZ/neHKq5LZhvTaMg
yV2pwCUVJIjbEzDtpVpJARgFfhjO/y0X/SnWYL/JgQ8erHEUKMWRYnHqQACT
bxp/y6h6Zg7NXRzY6HFl0CUjc+WGtWOBv1c6Ma96AqkoxkLLoXczIiVLidAl
HlbmDCrOLz663kqSHDZYvyuWcYElLGZoKBcuNSnxK7KagpEkKgswVjr/m0Gq
MvbXscCPwngvGnSwQ61EH9D5UGS5jvM2sz3CBxHsQt3JCvaxYZRgttzJ9Djo
jEETYY/4VIhVLqOjRZDfPqFNIw2fjXJJfi+aAbDyS0UjW9vGHUQOtC+602ly
cpnPv7SwqKvzMxvRyy9QF5f/1ttOx/NKSJrtw8YKfCt8XkYiVkDYzo6iAS1L
/9qWnvhXU92iVsFNhZzJXL4/6vbbpNleImCd8UETyAvp6jUdp4wp45qtadji
aTwbqT1Jzx6QgCxHRpr3js1sVClALqWI+6iXxQbRxEFBb0oqbdKoSJbMn+gJ
W9pc/i+X6Yfrkh2Rc2kmwgVLgDwl/p7Y3SWvhyoo0bcDfbmJjf631R6C1tzS
M85/6tU+UUvErXi0OLQ2ykykYT2tXEwbuvMj9NP0yvsuJ9KxZlieqsVZshRR
F1AsD3qHKsZB5HigLNoOXckIB+GMOiwioPH6ubhcc+J5cxCGFStvOcoyXhYb
DwaPJ56u4Re5HDrE5pacMt1yRoM89hUcX0z1UyGvdPmLw3G4xRuUbYBrkezp
ljwQQbQa9cWJtF6mTJW4k9huuRYY8PQQjhm66bxT154JhXZFNCmRY1XdoOxa
98WabaeVs1hZdg8cTG/HOLFPTqJfVVNo9UxuXKNIhtNVOuaTVpj7rAt2Dp6a
chfBb7C/mw1Bo1LcrMQnuAAkvVna8+aI0ChMnIItOnYGydfaaxmbPi3rkdRj
bl6T6x3vVSflmpEhFwpN/+3k5U8VOneevzHtz1WVQjclEV+DEK7OcQ3qk9Gx
heDnzCW0IiF0sjdPc3Btna4+vGZmExXe4vk8oTA6gjYt5oIHLLdPhSrYQOTb
uu67LhgJr49+d/jNE0PI7TMAFMQ/JXJfE0o4YG5zI9qPQFrobkVpBkCBoDcG
viPGQjE5bwMle+hQmpXeeT/9oSgDvJFyBglFWMhvZCeTWJMMha6ECdE1+IwX
97EwlC17tUyIQRhcIhzfoyuJb2Ff/3L350h0MsD8+gbq6uRgUFNnPRY8K3r5
ulrnszLFzAzTduNkFytTeaoD4r+zTSWEyXdw0kBWC76dGaMWZdXB8Dn13c/V
HVQgK3mR5HCQFJA1IWNt13184xupX439MCkpj5QqvYIlxc39XI2Xy+WRiyys
r7KOt7//DJew+JFj+fTVVsbLnACnrINziOWYGQRgPtncjlF2EJpCGlITo7FR
0ULmtYXsYQ5K+FK6/6ZbzKwH0xlyDO9VxuWlLiVBcKrcLG0HxKU2ImyHz7Ve
Yc5w+1xviQbEHqwnq9ymHoAPIyyh0gUWWiNBEb82IS7PpvKgPoPepocCTKk2
R2qtSBtGG2CsVzK7m8v3SDO02UUUBmBDSERSv5lNmW1ifY0ZNb2HfRg29BBJ
xZXzGe/YLNgAeMu/JfgSYQ9nfUcaKOHuhvBG7yIGoJuHuJUcGGoaGnKiM3iy
Cmu/oVFm07ugZngYlmtMRbAD6plqdFXwLQFVt2Tau+B4ImLhwOIH1Xw1Ip0w
YY3CkE82g65SpZVHw940PzCtC9v2SyejaWLbj6e4ZODQw4e3Z3Wy1zIIgS0k
IyUMLwlKGVQGMMVroToACxJFLyy04Lyq7eSU9Q4/6cvy2KKCwG53Hpe6y0gw
PVFpLhwRGTfvkeRJh8qJSz4bS951SCnq659Q9vymgdNFh9eGoWJeWWivTM1T
jnSCRVmtWtigzjc1ZcnI+Cj1YOZW78A6L8Uu3d7fay2lvkA1W+N+Mj02bedI
W8g2RzzKCZdALp+6A4q8Yx6uB1vacCAvEsvk6U8+lkEEY8g7/kGoFHU/zq3y
l7n162f9uPwHjXHbhja4U5v5LkoZHh7u0aQfanpm/L9pYTxbSDJPazr/zcFg
0qOiPUerrnmudYvY/GUrVkG3FWZiGykUcUsInS04b9Ea+xMu1cFbzHLUlqeJ
XSgRnMeg+uZ4+ldnXPZsoFmxWFFYXd3uWvoYyB69A3eSravjNZ8bsraFzjfb
ADPyKUeXqtBuwzuUPtb6WSRhZ2tlNXvfCS8HKNPRi6qsCnQlBDaF0MssmJqw
our9JjzN/e9SHOXCA930g0iutNLIQleqjKUCl9ri5RmFfWjR82EkibFZR2tg
tp4MHaQcnBwtvBMGa8WWPLg5J+qmUITtolChjhMDacUMT+fwzCMmi4arfgAV
8bltn2JJYNuPx1+Jbxq4PKNOYopg+q7CcD+9AQEHWBD2NLW7GpSFiKszkWgS
wQHCngwZYXCyL+LmKk8G/xTHLv+XyeGG/xl/YeSInopeq1tC9bnGHqood1hO
3DRtjzqX9HpXDjGOsGWfgN1j/c2SrL8cYheF04JmdKu3e6y0UoLYnSJI7XZc
RDwJboZr/TQzsuhe8ei289MALA4Z/sfwoFJ8hX3qZ5nQ5KHMBEMr93TNNB0V
+vQK30oPLr0NV+42aK3KfJSnec/JgBsXE3oKk5YgpJNIpxsp659/p5eolCV4
9L/mSNEUHNJ/GCEAppb2EsSm1scZsp6j/hbLN8DCc9Arwib9ppXQnCgu979A
LvmNRns9pCLfHy2eY4H9UFUxdo6gMt75uSJhjnX1NaiqNuVikPTA7sV34Otb
z3PWYLyE1/ceW9fUwBxIGcaiFF16THj27EAN3HV4CytPdKC/c+IRbzToCo+a
Z7hXmDBrlVgVyNUBA2s2YEx1wTR04FdHMXZ8As1cwmZntB/Mxk1WauQOo7z0
sO/hTnKU/yOQBrzywnmq78McspgihFUluUPj9TifTpfDaHffdPbCHjkvnmK3
QGoJ0zMgSqessp3xsuoAJkOkZE0/5xgaRnR5D+a9OLNURfhwF1aO6IpIWtYT
/y/YA9JY5KlpqKHXBGQC6jexg3fg9bA8dDrU9u4q0xK4IoUIq/8MAiPqTsWG
2eqn4noIEh9Yqcr97x78AsatGLb32LgyNt00Hk091DFHmGULo7RrOZCkwHgV
N1Eock7EEPzpKK7tWy9DiVDmnO94AHfhoJMiqYgKAnfvncfFJuW0q4Hs7HJr
/XzvVmA2515IntX1Wq6S4PCt9Srn7a0Uc64nW3/MNZ8VyyHF3kE5vHwvtVtQ
h5P2O3eCLnn+6JD7pFTKGO47GqUwhHMPuxU4OGeh9meDz+PIQTZ++P4E7WLX
PXfJi2NgWKysbxb9dTueVaDKBlz/R7SADUtWPCaojNTVg0bWkyosgk0LwWJj
FriFoFm4xNM2OCqdspS18ws+08MENO6zRw1YK4U17WqUMwK9X9Rck48MwGaa
ImSW18B58JGusPeJ5beH/qoIGXb1cUb+wxK9e81VEA0jImWyDyN2G7b4HvEn
RmbF1FWWU3yoKcdmb7zvi7rXNrttz5BCB/bWvWWU11atzOww83GHf3oQniTv
/sVc5lU9VH2GmG16lbnhHzceaVe2wjGeU2hm0mwt2Nbu/He94/NucuBh+zn8
Yb9JZZWBtJ3EMVEYcQMGrjg6t+YzQuPQ+TZ58NyFhk1eZ1xvluBeA2zxjydc
8HIp5LGTuwfD/bSTO5tBXHHFAt5s6Q0yC8RMlGhPU8VeU79kFkw1SkqJL91w
zBVIgO0guevM70TPiy78qJF+Pia4sQbCNw1uBiz+HJZgjbfqnWWy+4R816SW
OWIUwco5PAxSRvz4HlobDwt91SN43JhFDgibz5WcWqiONgKmCtXqjnbmKAXb
L8ioI+ehNO84q6ZkYmsxyYdHAzB//ENZjwNFlQqghbh9nm+ecq8ElipNUaiD
K3+2ua5X0WpPsGhdZ6Er3LNPaKbvi5TsdN7TXDRG8VXxJZyYCVo9sxWPmwBz
Y8thqabrUxtWCfR7jZVfMW1DlSmFFas3cTsAuLqLtq+AOmol3faAvUbGzxb3
1vlCAu+QRoonGqT+S/yp2OIE3xgBlMSIb3MIh6W+bKKwyJvHfSg3lRg0GMbN
REMuxTZwAMWJ9isBOfLJ4A+8/CkFAl+c8D75/bQ0Fdq8Vocxw2z0mFU/JhO+
61+iOENxIB7MDv4/tMoKiA//3KkEzgNOSOLWfwyK1LsJndLzFUcGNSRgsC0O
3QLH+PdS3u2EDpj7yRkKuZRe1XvtKheyQSGgMskPJr5yYIrIiz6NNs7GAmTR
N5fWBgHgV36X8PJjzH2QKSmwkhC0Ei57YO60PBHj32Uy4i5tgepHQD9if+ZQ
lLgHvcLIqd+iu155xjK07u/F+TzzMQq+C4TaPQaiyPG1r1Ji7+cz6Y0jJ0H9
TwLhAcr+oKp6CWbD7+WXjie8jD9msSzktONqax86e++OtrsPQdaahbA79Bby
rINiPiI5LHrfieSGKTS0NVkF1lIFjqLAFDknhCoV7k+RneTA2hdKrZxrW9cc
akI3sfGicr796EaYZ1VXbHZtW6RF5UAvTWV0o3L5EsJ0sGFDVBcB+Uf7KKcx
qb9EFLJiqVs5sveG9z/GxvlnvhLy6F+Uq5ARqttkhWwdSzxCseMa50tHVb8a
RzwUQ72IcBlzUl5L4krXFnxpXMytmdXs3lnlBVf14Flr9bLB/P4N11YTGFSk
SSLnoE1j/Kc8siPOrc+bLagrP+1IqbpYxRNWJeNC5jIH2QlOVj8nC1ru35gd
3whODEB4hTv1U/jGx9Yk192y98HyvEdwT7lJGYY8k2tJYjwn7//1K6WSabte
QJNazmleqJkkpK3IM7S1h3piysyz/H+pkcs7G6qcZIP1lZpWOB/OV276R1C9
uBw9hDXr8LEap87lY6UhNfs3kwhqdmx+uCvfyid8d83rGuvOOrxDorXv/vFH
xMQBTQSkzTP0MKbsFBON8JKBBG1HgEP3ActRnQu6k5Fq86IFyxDCxBEWij/D
5HMarQ1cfxbFPlPwnT4UyndvkZVMANxzQEaS4FsRasfbClt2ZAxyQAba6FXG
YqGFUbfgEy+Rt2hwK/9NQnUzl0yGD0ZXW8kH89e/L98FxPjadPmrwl5cIXn/
8NMJsZyeowuOCVugGqGTaCAQUTvWjo31xShNNmopHbo6ERX1OAZ4dGIfUryR
YUqhZnpvDZ/4WLHW+vm4DbHraPDEPMu6z5P5EvJ738KVklZLAeovC3AQn/3x
pRFuc6MqJuBGMZUtcDmjwppVnnkqAZe9CdUARTAlRNF/MsqjZ7E2zn9FeDlr
BM8A3BReCZ7J79EaP9PZmqh4RYKbDMAs6gQGccqJEpLy3pWfDO/0perfZVmk
B8N3Mg85TD4rLnFN1RGqJNJbWlm4aARwRVADqL+7N2EFDeyrxexc6ulMVdWq
ZfF/GHXhSd67kDR3MCU2/+dxJEmJ/j6/Y73VSZYoMtzWEW9sgTvQmJSFJWNY
f1FQE+OQk5LLA0tLZnRUkQfclRUjvYbXJzUM65fs2ZjSb/+ddMo74nhXzTdr
C2GsL2FB4P00PTdTqjWJk8ks1U3NWIiyDyb+zrQsCMcTwbfZA94ubW+T4y+Y
104AIPWoeFw/fnQkDYEzsn+ZDvo3Aa59fpBLIeguSUMLXXD0TJxCGsjxWc7j
gxkQJ7tUNRSmHvZfqcWDxVSr4PVMyR9sVGfe0TYkJUMR/MBoDCT9TVA0xeID
0HSnohRD8yvON8Vt+buJmxBESKZAS230sgLeuKFSgvz4TF2CSH0mIkBJmf0l
9tUjre6IlqzxR8PJjEF6ZIMXvka60Hq+CKJoEL4pNjiyKdxmMPSoqHvJVrTN
y9owlB/3P3izfQaMGDdARPzogZDf+NOtz7J4SbiK89YvNdMARtNZKpR0WXgm
PCaPEUDql80ar0T9Mn30+/vn8ztRTLzCaInCX25vSM2KuXc19qnvjUOcy28H
NmFU3O5N1UA79DMnQyiK9tv2CxaHxxo3svQX66w5h31xQBBpZi5prJeqIGj2
zJShs+OYt/tExlXdcrbl7oYwN22Bdgu9WuKCkvvyO3uf1VloNq2+IFBZbhm2
SHgsAheZgK+u4W1PS5iLD5GFCFOMMVaB6G9mbv3rnk7PULT0evJJrUnV0Hdz
W1hQgcZE/6NkJRNKFNO9GbSP112vr7Ph5mxJv3GrlPlly9pymu4ntH+DWQqG
Zab67yRyidE+1ZDhcFh3nstrE/UKulPbpLo3pwRUpCVqBMjs9t1nHPKY/mmc
bJNY99J/SOmLKZy0iUYZgFBW/g27/8WLSXrur1Hlbovsuz3+m2HzxITffWGE
bSZQC5Xae1krMfl7toO1Bm2uHu5kNkEEx2FkqSaNBTSRcZXWXAH6npeJJzdN
P0dZApwyn4h5d1T4/FxZ5Ubk6x4452CcEZmYyQksaoSxs3dWUhJqiZIR1zvl
vLotkRdLM04te8zJlVetPpNdU18Rv6NHU3KTerBk9gNsP28xUYouM0mFp8GR
fkrUuVtYqgUQtBrXR9kho6k/SToR7FlH/15/NAESYvTxafv3Zd/pA7p0EkGI
XdYZpNby9w20w6T0vJ641OyEbqmlw36390FbSXy8OcAw1rofGniu8UXQsjCk
z0H9cfCaaqZe2vNteGRaD6Kt0X5YR64ZimDt8Xl/eQjFq6fwFCnifjrmPM3T
sSxhvQ15EZhYHq+O5Yq0nTAady6zlak/FQerSQEJ7IHsoIV9pulzs39yTMu0
xb6mv7KcCmglKQTySX5nul5IdoL6o5HhZES0b69f60XGk06746/VGrsh8ukP
tH7OAgCLGI8pX3+M24V+Nt6OZFj3j8gU6OuiB8qwdn3z9Jp3Cd6KLLfHpzlx
RY40FHTWn7Ub7EOYT5K8ZiahGetQEWxzc7iiOpFk42g/ePuEMoWpp3VAcWpe
3lQvVUZUrB/9vjT6gSEwDK7sZRCHbj2J2QDGmbUNnFMeYf7zDJ53J6/izK5w
fCxktcbpBVqGI6DML7a7GmxdFGsTInYwN0BkA9OPn31VIdOf1xAhoWzhlUl6
vcVCxTNN2F1QRaQKLHYOqdgXwh8UmusyRdmF2bw1qu4bNl9kr14SO5jAjJsO
1Mv6T1SeV75Hc7kXO4PQQ0TLdcw4tPvFQTvhQegs2/lTOKWm20Sz1FgvY4WU
C+3vZV0p+CrIWObhzSoW4JyHYFWrSfmU7KWLwRhYvERbtE5JdI0iEtaTNBl8
kMeB//JaiV5LWBRkLrmjN0xiepinEuuzWU0a5rNulD1/57cRcoUd32dxUY5X
jsFuhWyyBA05wkgrN1QheSByb5+zqjKKFg2W7oIvLi3BIe/8LDo8juFWk423
FNCRbJSJH0NgJjsGntFhVdqMZfbbW7dutA7c8T4YfkPKyPF0qBW/sOSp7Qv8
dawWUGRCUbe5U8fsWJT0oewTPuAhbaITPpRZaPlftNFDzARij/c8Q+2hVsW1
E3f5t7ak9jfC3tE8/DJZnQSfzor33pJ0uhAe5WDWQ6jJd55m/2Sk6IbDZ909
XbxqR/dQ9wa2F3lLf4EmgTsWq2p+tLuGqWawo8cgJ96qqsV1eEHZL1ed6zlI
2xSfQRaUVbGrpQFFXmjfIzcifsBEp5gej5QRDnEkPb8STq7m5Wx26u3dbNzg
FDl0Lv58jxCzxYdWBaNsO7myS/xmwQ7qJR2mJfeNYen0Aigi/+OGb27dhKEG
ZA8J0pIB7L9Jm2R0DYVUHKjdfPVLk7uCKBxmdq6t3Xhl/p6BVx1qw3/HmMwR
x4zoBETZYfbbKSNDubSIXQayIAe7ppqPCQVWgcN0QDLXECAEbOP+her4a6my
rYreLM1akVH7EQ5W/KTq6lYMZBWEz7MGR0p+t+Kxfg1Sr7YcRW3PV8GhE9Ot
Elx0zWUb82aTKfS5NzCzRFWXlySaFi/QKufKY2uv5m0RBk1ZI8hkQNZ6q4PT
H7wQJaZKqtzEisJI2ug8CvXJ2unYe1vbu4/uHxhNLR6uBqTCJn47T5Gzck4n
CzZySwKTXsaluTzuyUCDLbmkd9SOQZHUG00fN4l/jeZ9YjK/U2sTa6ut1VWy
EoaIdwUjCWRVw7BPPxDr6ngBgsQdMGkj1XUIhIG6pXLddb2NOget69iGKOjz
DmWR79G64bXjpYkPSk1G8FwLda1tdyANULswGfl+3EYsm9iGCECjY5CTvyMJ
VdZBtJJBd3wXojMzxQZSRzWd4I6uxVGR784mCbyk6J4RhRV9zPiW4LZKDlpv
09e9wWeMxXzTd4owpYj9Ky2c8vpNz4NjeZ33fk66YZ9VlohpQd3eSvBl3qfS
sgdtcA5+4Vn2aMzExppmhJ6Z6KkfFMxM+16BoYBFLifhJD0d0rOLJOmZ3K9H
H7ziSxLdqrqSAdTMBla8ja3FFoAJueOQtR4Zh3LDV5HDalqOMsslf6ZYUpth
lf4YX/rbEQAfW2PlTvvFw9lDfF5arf6O3sgZZXYaz53UeIBMz+yc4PMiYZ7t
1zus/9tLqQm4n+AYYM6k1R6+x4oxEiSXNRHK+wZcFJsKnOVv22QCUuawsyeN
/zwW3bXe4oOxoKaQu4gemcUXOJaXKhDyExqyftPngUqxkA/UX4uGvP6ANOGj
grkVW/JdnvNxpniUCWUwQEWVp7VQ733c87ytWIF/28L0flwlM5jhp5UjCJXq
wM+KY6Ac3WNEaNBDCE4V0sSm/NLjpKd+5fkd1nNES3hi7lLr8YnOiST4e/Kp
XuP/tGqEWd0z0IUJsfoZ7TZHZyo+1l5g2mgnudCbIfnFGmhpgeKBTsNYFMlM
IYBqJhZkQqU8cQyxguxLXHVgZSIsoWo9K16uEFBAiPS/Of7kPMidJnGM2YQi
NCN/CEcfXsKynAQqQiGdFd+Kfu2Ey9h9TUZPZ9LVSchrSdsyW42jpFiFPm/Q
gitHyzNWwNA++pIDMEYz/H1+WYjv1nBmoQ608kmygeOZIzp3JmYA9eBqDn9D
WFJjzVa4b6REjBKmOQCSA4yeYG8FnZ32hWdfzQT17sPKqkiKWY64Tg24NWQz
ju+CceXeX4pwGDQQ/cTooRALF3FiuDVj/Wp33PdYZm8Nn78G2vPxB6i8sgEc
eS9CS0wLtWnaLuYAJIteZQxMmWzcr8a2q9KXW83VyQz+/hc7iiVROGWOfG09
oUH6K1T5+tkPI4Fq9ZaiLKAMsg8oHSXTF2dWpgwsPa7qCL7sfatqGxZowYEX
tmkDnQNPIGd6B1My8Yd+/LkT3S1kkBkrGRhQDA/EZCefbzocbVs1CKRUZ3jN
EkjqRm1YcR6r0JdBH0jKy5okg88loKyuOvSWoTeSic0nok9ay/wIeThLBxMJ
E6+WGPdRpxXckrN+jpx/YGo8TOESxi9L4TLbWd/BnyGHJLekpj85I0laYwiQ
lCEgviNspN70pG2k0hlqb9oZYRGY820OKeJazCpllC4zLH7UNafw4htvfAqV
NMtxshSjvx30+pD6QIdNLHC52fsEqiPJQpp0dI7AGnf6QI0J0FW+1LO0jwRy
prX1s5TaP6O8LE+2tDHkHjp/cuw1Q5Ipdh8KSUawmL6E+uwgmEaKgBdZm4Wt
RI0t9w5ma1AsDrVskP/Gimd8kP6Qp7O9YygFB2QztG9fC+Iz60egi5ZuUmUC
9gb1PoZIAEMgNARRBoQeKlkCg9MDSStqPKhHevl6ZDCh2/h2C6oYlBokEc+g
xPFVsgyvh/Hqn8ukkume/Y1rgqnRfAkYQrJ1/0CsvGww1IRp2nIRRpWa6lWX
Av9vjkXPWCvQ9IF+YS8/d6uAMXRcJdfovE+mklHHXR8EnZ8Y8kjvxGvBzmiC
HL0Hp8yIHCpFzAMLmYG6MkXiQg6zKbFdv1Cul59U9AwmV4UMW9FxmnnnUdaF
DAv3DMTKyBxKJ60dm3j4/8wjTVKjYNVCl1rGx39YAzIoifskk549mAHylFH9
NRZ1nxQ6/8XuUrPG1ZeOWzeLNTVtYEdla7v6KeGjCyK965w2Cs6iokyf0SKq
HdwfbxndrDts262jtNx7KWc45QXuWT1nkukGNJ11bHttyUiEyffbYU6Dn1b9
/vNihPSyGocZkpELZol7vEdDOBwBOFzA2R1xIDHWa7UfCcMTD/ifnJn2k2EU
X9AxdSvb2Ov028ZlYC8BKG9jnEZf389EPGuxlb//t6GjrvbbWj+ITSxeLnl9
WavnYje+OasoqYUZVrUKCIHd2QRdC5GwkX3fmeVVMbeYASg3TNruQFZYfiSs
jJs7bCrvhEhwJOIBhL5WUArRUqo+spCGt3YmPYkh68PdHayAi9Zm6USI7bXC
TdeBWHovvAs3yuTIV7Gnrde6yDUc3tD5CvZ/d0WnSYz83tBD3JgtvkVDic57
nY3fFvQPzH9Qp32x+vumOVQRiOcu4raGkRZrabaRcB0yetMbsq3pHUwYdHNe
SeWodaG5pN/LqAN2vmLVVy/r8ZeWOmfpqHBCxynPUF5z3xl7KwTPfn00COaj
zEEZYXtGWPZW1RtPO4qNtSzr58evpW87AMAM0zG2RfkLXi9ggftfZitEQnBZ
y8DAwlFiemXjQ90/VYnuXRe6tpY79xuUch9v3JtlyeUAT20AGZ1Yny1CrYrD
PtgyISQp57VVkDgdWRRtwKZhb8QV2M3gcd2DhiifrkduBwBdcgGLKZVRer+k
WIjq/kfdgsieolnCo+fvGbGGQB9qLn4vfGomqHX8uONS9yGVqPCy+5rrqAzE
x918AAHfKyJEzut6Ob+8UCNqhdmFi1B3RFuuhhFWnO6Nayx7Qn15pqdbc13d
2tBar4kB48LZVmuDan1THMpZ4638C67OaRw7tgKbC4vmGi9HALRFGULvPmR5
ld9b3eFbxEl2zYeXNkqraDdP/zn4QJsxQiON5HI1GcQgHlu6ypmM7J+u1HMd
phahvEJdv00jr7eods2Cjw48NVkLo1INdFu27ZZCGPD7mFJGlN5cH+RNz7qV
TKmYHSagF3S2wgWG2kp7p4+tU8P1FetffHfNgvTznpRgDprhZhTcON0OzkId
Qhvw8eNLvGz1elcTpkLgBgx0k7NO8EnMcXKR6l2anrHr5TUqb0R2IPc71uhV
DUki6/F4v/92nlKpbFEV2U3wQHSZaxXkZ/O9BLRZ7yPzwOK2Dwcbd/xsGqSx
k4Jfv04fumcQ1ibtBToutn/25KbueZ0tq+3u0xQGhpVE/O8gqkDF+jqimm4j
UvEy3ZfiHNqGP7B76FM/74z852PTIzTSwnUv+XbMNd72cAFyyBX6WGkYOb3O
ssNg7loxkjuhbpVV4YDWVoKQepHobYLrfut/VZrT14SGgZHo7voZkAdDa3dW
YZ+LzbASo/W9ih6mTx89etbMUkef48iGoW54vcKG3gjJs9+GZf3UTGSQOyb+
0WwbuPxRaS1FdayY3ku7G1FBVUaY+Q/+fNPvV2n+iv70U0vu+MrKW8VTG9ek
hB4X8O2868Gd/wHrYkKvR6mhVSgVksPK0oL6LeBDlZNSrtXK2yJqBckKXXuM
94jvBhd1uh//+/vnj7Oc3QUq9NpbYPgU1hjI+Jw3CFt/ZcbrFmRJjfLB4h17
SkAS8VPJzk3jEsWJaILjUD5QIpbUesRsL/vFreMpThIyQwOlKapqMytMT9x4
CV/TEvi194CLHpBrqlL2F1VGoXVLdMd9dzPGRs8ps/p6Qj2nMY+/B4m6Vkx/
3j33vezvUNKV3XZcTXiqz9XkuYhSW1vKWalXvWTKiBj4CgZlWbaGYG6Sgx8w
5zkML0x3BieVxiZzrHV6WAggpf/oWfTq8e7Lc8QV+ZjJMFt6FUBHDigBQNn3
VT2fxxQu1xDFm8e/bx6YPMzNEQiN1MQ17TQre2ncc2CBi4Su5Xqov6q9m8B/
ddLU7prufDG0NDjdM6jrNtyJ46MZXZAbbz6/PScYdRnNJpe56fOilfT4JAu5
/Z3DVCnVUt9XO7Hc8wvSPcLbLqS0/gLfJylqEVjCS1s29ugdstgiop93B73E
rTlk7YRKzbWsPAwGY7OEv7k6HrZwHsiI9joBHJ2pIayGnG8Opkne3AGSYqQM
EjCXa19ehNJKG7V7qAexwofTsG/s/p13vpMbAJc9vB28c8arIwlgBMlDTjtc
ae5QOJnJuMBqgq1OIJA3/TaUENON6czjimZxTqEBbOvD1juZhLmC+/aqWz/K
ngy+Yj78vfHRydWotDo6ymuHUKqzTTBncYZQaOF+lA6vIAs4+/QGhP345Xcw
7g4L3EwI3Ed/mQxEU/6IiNbbcI0DO+toLa1phlBxYFoyMDQxvHtJpc47Hslt
r6m8PXkA/O5BdBd1iGt6JQPxZ/Vv33LltfvS8EHPz9NQVG0NgnU05zX4D5sl
eyWmpdxNhRS+W6+H/90OJRSIrNY3apeya4RsyucXuj6/esLUkSUIaId69o4A
/Vc3JZ8xcSzKSj8JmGRgcR/jRIX37ZmICgvqfS2PEE/NSEnlxvsvu2jNI7sT
JIxdhHNZhXi37afJ1UcrfsKFRfdeqsd6LyJEpdGWjWJ27ycty+cPRLNAkfha
G6j3NJ7AK1HRuSyUJWHRhdgMWGo+qYbvt9iquDMa2S4CS3m4m+UouY7zezQG
EGLQrAjPc0L482kcAIPU4o5WBgDJ911Jhp1Neonx0HdlcmpU1j9mdm7ADLIO
UM+VY7QZK8FCYcqwF9b9jrlQKLdxZbxteInB3/ndHZiILMJdtBsAVWNNAFbZ
bguqf6HpI/Jwlhr9RJjN15n4gZ+3+3S9h/cWOOdwtridIIxAt+zMaA9nVmKg
2Lc1+3xGUyl1sQhY6FNtCHggRJN0OYS2NS3Y8PlYN3bycQ6euNU3g69MW5yC
WR+/HqJzoIu91nvtT9QbUagxhuNTRQ/x5aQ8D6+3/7g2VXGoH+rWsixC4mGp
Aw2izSuKk4mHQ4Q8uGAKmXl2itRch6OT1dZ8w0Yvcjttp1oQEY3hqFnEYVpj
iR4HVyz5PO8SI1Z3Fo1KK9HtNOesLrVha2wD7d/5afKOaHXnsZW0JwrVkqi+
n1iJSOZ3Efc/K3EccquRlVX7GijflQBBuz5EFLWnqmzd+GAVdpXF6rR2OHuD
E4F1Jhec4SdDoeMknaRznq4rD+vctsuVfv2Kh/WC7SBkj/6CO/lyWDpluIgJ
K6iTJPwy4C64eq5EbOkOwCH/EcdYLw9iXoIJXUXglfIGaKwPQRNCYBJcS/95
Qj6Dycm5HOJe1k9fmpY+n+yfM16A6wN3qdbpI2Iii5COnio0v3yU//cbq4MQ
QKMR8PA6vYYjr51AGgWIwt1mZHJ7702dKnwnpq/b9XN/oCeS3xzCGowleBmA
P+Ot9SlWGhu+29xwBp+sarcpjTpzuxdyuT5ey6A0dks5AO4a1g1elEb+ejZS
9+NbSQ3FRPvxJ1sk2P1LePGcs4dxnMkIv6MkTpUmgfrSw3kOki7hsarMs5zm
mnDhXH2uoXJWNjc6hJ+3z31lImGGRfI2h6jaQnVugOtYFJ1kWo3u9FAX2pZh
Ar06qQtbX3a+QJ8OQrg=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpegDS3XgEQ8TL+Mydr5D8TfAI0z2xIsHZ0oq0KVvVz1P8vxpmOXdSm27qHUIaX2Gj5bttI8rXh3THV4Q9q6sQwK6Gaf8OKMfprnIrbd9Et+c7ydEjCV5u4y3Va+BtinPM2zCSSONTNqhwTHHEqf5bYozKYPT35CrhN/hgUdKlVid/5PWuktk0Ml+bdlmwjiGBYRx92rRpSxYtl1xPvUkYbhFjAy7D0lhoa0iSH1+Af3Hqd1hqVTE32rJhEFIN0tVt+qeVR5sIfFLir8ddr0MvDDuQVi8KwNvUzseuEjG/XHBMoTFwAxv6PCBg136KIdEqonYEX3aXD+Ba10bDvk2gbsJ2QP0rqJ8ttY9GH3FzIiwxddLUQ2CZXZHWZ7DcC9NcUQ3AQxiQ5RqCc4KnkX9rrC3kYrDsqdQss1SWlUTin3OtJ+qlPXklsRc8BPVSLSw3lR4cMZneuMxXn9D+mzqyZ8cW6gxGOUP2I6tx7LFsZnRja+r5y97tpQt2Ah1JvpQR1jQmYRSiOBcOqagPSkYRq7rX535LR0U1ON6bInIOOO/2GoiDoh5Nsv9nJ/19pQGNCHCNS2RxJZulvfowLpP+JoTs0jIUZiJ91AgnG2SdS/SbjCIRFSRH+wEttTwLft1RqUjEaSyFcnfn11KYvZwJE1BbLm35pXG0n8f45OIQTvnr11WLBHDL48XdlyKeOl5XnzVbk1E/mMF/SNHClJbgh8TbfsOJdDZOPBbRmY27KCMk1I/5NngqdfSnTCYEw6YZDy7QMYyczs981fLY41RGgcv"
`endif