// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JiYE9RCV1SWlVz03ImWqzE+lZGUNGNG+2tH2TFN65rRHxKd5VZAz4fbIRvzl
/owvqNeI/Voh3C7PA2vzCUnV88vPyCFeqcRUi4VZ+Qq1tmpW751Ye5J2FaKy
qpM/AcZLoSmFLBtAUauv0boTTale6mhr5hEkNFkz1cPKJQ8E5OGmmzLLp9Eb
oNMc7xCYj8GB7BgVYWc6+DRIhFgoUFKsrmxyw9wrSFnfapjQ2BOloqK0eD5N
3mwja7k9bxCkrZ1tRy51n32zw/6uTnPyAPNREjAzxXILjE27rrCKEVHoYmhB
oosVnbV589RepjeHOsa2N0frlOmXuxiTh+gKT6uHyA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ccr6D/cilbu0UO4nUKJQ+l3cvJyC1w+mOoxHpCD0X8HrKfqHHYvBXRISBfrx
le3LVelNfprLhtUVlWqdQphTMeENoORIqzzbb3b44L3bHZx/6YV8MdVkRUKD
IYb2FMN9gs5HX0j3fFdCPuF0vZMriz3Zx9mtmGymmDHVHCHytGkHIoyDsFP5
iM+OITTteR0jhh9Jf9vP0YBU2IN15d2JxZk0u+cIwemxAXgjwnIVhHHGB+/7
5DBeuI4y4RqjSQ+pOeOAz4IpYPNpPkcRPbqgMWuWUpL493c40NuweCJpdL8y
nPB4FlfYy8RC7iukA0MfpWozZSrSbU56DWRYNGcmQg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IR3hGvADVknkInARugVcMeFBte8vPhRNj4iVFMknP8cwwIoi2jbV2OXL6B3P
5t5d1Kx+Ba5NXg5/7SeSdQ7yxQMjqbFmf44KFY76nTIw6lx61V7swAh7NHeZ
5Yr4pwPstmDMSyIkGHv7PeXHmu9CYzQJaqKAIZ9bsfUSY9RYg9cWmI3yMXfi
MlWN8aOVX7HxiLCEN1DJgUCQAuNJRZe1BnPXK4dm2GGYtIs9IyL39UorJw+X
ZOGUtqc/GG9U2GR0GvC/U7zvOCrRW6lSCnJJs2ltfzpqmyIjONie7FlY0opl
M0fuX7X9lJ0uA9i4WRoh3Nm5v6V0Tv/8FecEeJWj5g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KmI014EtL7jEqBK7Jlvo7lLHWCdcgH5lTwaHQ14tO7T4Bx/Gs31O80yKLvTJ
NYZ7yDI93zCh8HXAofAapLLxKbWXrd3Bdbpcu/Wjuk/ManCJjgqHvIJRgt87
SzBCiXlxAckKvOQNt72rDrLTwIQLoceLCpdeAYC38Gyx1HBAyRvp/UOptek/
eZtfMWMFgHLmHf6PSgxP24Ayl11Y+Evo+ZFRIrMGc9CmT2CFianS9oSM9xPn
JaDSb1SuJ1lZivDiuBOXYxLIQ/zLY31dYwMnw40Sw4Xy0QCg5yAtkF9hLMpU
KZ0Yf9F+B8Pda40NpL3qAQqEE0PcNInJ3zPI1Px5sg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
K+U8LoVjlBDPNvhN3npfv6IDVyJMp9WUMRE1x0H98oqWnfnj+d22vCAng2QC
JRzbIqPuaXjN4Bv+mFSBsYVFsRV7Dz7HUL3U1v7dtrQsaUi4ox2cJmyHcdDT
kqjAjEbDoAXWt2NvBoODuAlIekwsBODfHG9PwXndeDPDJCdDlJ0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
DPCG/0OO5Ao4Unu8tpW4Lguo2C+oabHuuUxoMVn4Bb7bXRJ4h8wbLdlzGCCZ
wU6OPmtDqQAc/fgoKSiHmGpQkNRQGlZ1d6UqTGTO715zWNzYickwtFabteVD
sW888F69SlUbUIsDHhxfBI5ikyK1m0xaKJIrpK3q+TmtLqgQIcnP18X9kIkG
njlUjl+ABZpWu+jLP0iIB/BXJY1kkkos3Ve7fmBSKHAxQK3TYfqyP5tT5U8M
rW7uCKKbS3Lt1pt99RSbhsaJoC2fq1YyeHZiGXgxKETF7uXtBt4Gu4/YXLvZ
QqqK/HGSTmVpQA0TqtIAiD/KVGHydJyY03v8TrJ7dE1wvZo1lPGAVYQpcIhQ
P/qLZa9nd8xMlqW3GGg//FFDflZXJNTOY0WD1zehmK3cWL1enpRPMhdbvBRG
gZj/RPEl03BS+ZteXbasB6q2nFVDzlFmz+VnuFQFHnA5ALVHC2cBjbz1/Kh1
zxPNbUxsIju6p5fynNagWWrdg5B3A9Ws


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
K7NFEQjminsB9ClVqGhhn95BxevMmzBXxKrLIdfm2sMy3x2mhIF/nReGw0ag
mnGYLuzTBXoJxSosJ/q3UBrs08LXEs646X1xcMzgUUyrS5bgwB5ND4xYA6IW
WyFLpmwXKp7w1+6lhtV9yzSFaCvjLu1+1rNlNlmpqrQU54O2z9M=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pg1Erswbl+EOMkrMW2CaKGj/wTuU7xEhFCnlnh2vjQIVeLZV+KUZXF+B8mb1
qBLt9Tko6a+PeivdYC+deUEqjG8Abqltir7Ir/2eB0wsyYnY7/ff8eP64v4k
FdffL3SyL9UK+n8ya/PULOZf0+sDPkGGSGwj/ELVbPXXBmYTQWs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 41104)
`pragma protect data_block
/jvNvheaayP6Xi2txKSAY+Gbl2hi428zxiSY6UDNlctZjBAxqNh9mgVWjBs+
G6q7uTqN9PliEemIhb6W6Oni6UUoit0FS2j81weNZ0mTRsiCHplGS5ZlXagd
Ie59HT9/T+i/Li/kvaqyOgN57GbCA128J3awlefuNL2SfDyzjIBLXsB2IEWP
KfQp+MkMZ674+3sYh8L8dBviij0F9Y/gj8boyOpwAP5n2SLIQGrrNp8S+yxz
U7yyI1JPd/GBqjSn9zM7xg9Da3covWrlkoasn9cDwzNDsBgeMTrHjzPjheAP
zp8M58j5tOq7KGfnzTLgkItgoROsiYh7FO5nXnBzOMGWVhzvyw9yfSvX5NNX
spaplWDEOREAlmN1NuJZQkcmrv5YnKhNQj0SrdtGQ6lGTuLfKC2wMZYYYr/o
B7NNDeZugS32pTCgYXNlrDIQNGFtDSKx+yuQlmaPK9NsA+c7jF1fArEMOE9Y
UH8BouHpAYL6vPACJzdEnwLLqdAtAedZ6orM0jqkrYe6os0nVqPCynKJ/azf
n1Q89nIZmcM7bOY5mr7b1VU1fk4yZDvctSazLys0+SeU98IArolQtyc3zbS1
lCYLX3MPSXc1uJoIOyf73nqN1hpdGxBIJqwPBgEB8kL/uEA00Uvt4g6vBsgr
cbZvnL81SQ3XNL4bRpTfNYN8pMTxtf80zAHH7Vd0e+VAz3D62h/AIkS8r+6I
5rm6j08osb72tOqsihfu8oqBfKziYOrz20yYCeSRIAC3Ym8ZZU93RiaB1cUK
HgZA8kLnL6zfORGHRkdFsbaVWV7c+2seS0dWxZGtYNq36ypdBtXLaFRN2mnQ
hF3phqrtIBH3yww4YPe9004z/mnBZvvQKS71xtxS7g7ZdgrTD7y41zioWnkQ
bNWpXPh7uY0g2ACjBfI6OQlDFYtDK02uQ31y75lU5F3rn2O92Kko5BGAUE75
9u+dBsPMcliXVm2gZUyeh2id2lUIjl6l6oIABFyM4QmAKMT1XOTc+BOHjZEu
3sGnOds+c53xpQG7lx5Gz0tew4QfqsLktC63sdXpTLwAy+NUzhyHSVQPLe1c
/gm/32ggm43nZuvsRyI9wH0b/qwLHoj6DAdhONNn5tiD8gPswICQPQYWWxE4
pL0nzcNZG3Z5gKlilSzazHCxKdHBxKPDhC+RK8Bu923qEcvbiTr7YcrvRiL3
AwXtahpgAfJy3PtkJPaIvqRF/mslD5qahSTZkW4UzwMwC5T3vKihEIUtQLgH
15m92dzaB+s6eQMX3COohcvmvJMHiatGhQVQtWzMT71RfYw/JaMFo0FHScMe
86OB67qdrFaradSYlLjuFGxizR1m1wH/8uw8nTUxUdtBnqeUZuNjOvo15Uxn
C+EvrSXc8FrTIYzVIhG+mCeFRasjxSB3l1tF3hqW/N4CtAWyorc9d07Ue+wE
qk3OwO8mElaP3LqbLUrfjOMog6gMVj6MTQDTFt5VYX6fssNrYos0LY4jlCvM
RbHjpXSLWOFrf9IlylZxtFdRDU9mN8iQ/3YzRNqz/pA+Ip2Y8KEsLeax1QZK
OnQD2JmKLWS2mzVO/DtwEW2ieBzZBYgQjjlzeVlI4eCbyY7HEkUecevOhVGf
efJMomZJi+nKeSqJlGCxbcUu8K6J9BfDwr99LL57jGAPK8FGjto4rVAZ0vb+
wPEQT62isNrEGQGXUL1VggiHgLcty2HYidDxkQKJL/PYgVgH8chJshIV6zVN
SPwbZTVL7rWmpnhlr6t4I3Hysa+m+LcUgwFjnaphA5vcp6E5fcRAq1fTwaRG
k3VXEPO5DePoYymoXukp47CxIlOFSkMwCQtbwQIO6lxyadaDxFdag2C03fik
8g4I1nAhwyTqZIxiu+zPubE5IpSUE0StlUnN7nARHmKyxQiL73IA4cAqGMeg
d0L1YKEU8ffz8/gNpKGAOnky9EbEFiTl1fsZcVGJTyTalRIz9LAJt++PkyCU
Nr424cURu8Tqv31j5F/5vNOg9g4U072eLlx406jdDhRmRKzIX+RmEPjp0rTq
sRVna7dAJdk2bUbZsN6ObeOb8GD+OnVzRxT0VJRzfq7AX3ugtlQGclvg9BzM
oXDJVQBVsdyTtQv/jNrBUCNOJW7bprNdIsE/Ar6hxtW2dooR+WndGnH/PwAz
DbKaKtrP1zZ5P1mDQncN8+v6jsAy3Lpp2Wh91BhTJVI1u94sT9Z3tib1pYQ/
bGLPwTMpu0rgYtrYJcKuJ+iEkOdTP8b3O8sA4B9a40PzqxbraZxXcmxy8R/w
GOwGSNNRX8oGnBYsrH25UTeEjzZ8liizj/Sd73W54BCwjn0akVoLQwWEbwlr
lENKCovvcaxRkglHufqdmC5AC6jaX6J4O5a+y0RLEaO86dhReQHtmfgHrho0
8JgBw5c8GKgtYdDTbQjHK4Po8pQMZKKba698dJbR4O5TGKWNzC8Ceiev96zd
im0IpBYKG+P+XeIGPuknZppQJCiYspryANpuytrWvstDBy1ugoj/g4fY1LLd
7Hyy5LwSlJt+SBPipoieP7gs73NHbiOFzNYdkaz28I3W2ugg6UiR+TPX4Cio
iIE1gBYAXhaTGGmKsmu8DsLzvDyDWoeyoaQhTvZMX847LQ7BknMCcdbQRhvs
6RjGj3gJfDNii3WltnSgENh/NsRCinAwHKccr9CgIGlWbXqm+1nCw3jxvrEL
9wQxCeWepbA4pX4HveaCNY4s7RhwYw8f+zLxPkK2xuoWTNik/eULCGKRgebM
JggcA98borKyaCy7N1c3gveg1yzzGT0HDWxMNORgizCKBT5LT+ZE3z90vNM3
DPeBc8GpdokZEoKo4YSet8K5NMlM/G14BzA4pH7oNU2hVws+/4qlF+Hf2tjy
XZduHldxPI5DW2+fVop+Ox9/tb71oyK+TziyluMpQ9LxgASRf42Xs0VpxUAv
/J4cehrQ7yRJKDdZIg7ta5j7tcokH4SHa1zLnacnwaed2/fgMhCBA6k9VPCH
IUi+HdUkgu89lgV+U6Ao3Nrg5mtnNwmmtQm+27m6ERRShwKngZP6qRrGfGfz
8WDUvg3jcS+5T86V650Rnina215nSlojlSsr0zhcyVmwbOB8LfrS/Qvhn9rT
MLPGMHs8GZqs0afO03gzo1JoRRER6HR85hK+fb8PDgowxSVk0NPpZtWK3AhW
ufnaGzBy2Zq+FxKaTW54tzC9wx8+q0rtDllCaztv+34Arw0mEFJnFEZO8wvj
VsdFO4BMvZpWPfJJyupkHlSNtDM7N6sPUtkJeHNKMJh6FzX+n/8wXBjGozWf
dcCzhiNIy7sgHNALTRIwpG2ErtOT72bfAfGttOUZWrIBMVEp6Q0iOiakn016
DgtJVR7VWzdGHE7NNmAqPc1V7LGaLAs/VmYCwxfN7XaB0sVI/KqSEoV1agCs
X+XuFcHC1yEHG3t04VPRX600IbHgqRGwDFwt258+euGWP2SE2F2KyS7joOXg
5E1gcEwHRGpgNRjsegVdnvzMEqNeDm/n61DuQjD6e/I/7TCtkKL02ZAbKxIe
AD2TYVqMzACBsbtDC/hWT3EakIkYZOusUIUffAjEiGd2MaS7MoMezHyVF1Ts
AoPCkQa4dRbjxwIRmjBoW33blZ3vv8Ccg++7jBHf82Ejp29t9aVf5uWfIg5P
MuABlvtI181aVDNh/93L88dBSrJnLH2CIkxN2cilaxtMOI4Lnmbq+cBeRoap
zdbZr7OmIiKc1Afv/x/2ZstIuDGwat2SlpCGfj1B0fJ+Sla5oIe+TchMaNE6
QOEhBvpFc3CFzeAJtkNdLz3EKLLu7S/TW1ESPVdL8sUBcK+0OG3KIU6gd+hc
PhoBl0khcnG5fBPVBmXjxaPdAsw1vXZHnZxyeBh1NgYryMOMFfoNxz8Bf6vF
IsVS5eDLzvP8CjhAYIp6rUSo0n/HG38JhcBCgs2AAKPzlYnD0ZnU+RW0+Xgh
D71EtbGoY+l01YvOdYES+e+5OToT57Q02KNs06LdC4iUz6cTjGrGbkLtGiZH
Jrv2EkcbFPYcpAbUvzR2oUFpTxDbKgVjrDhAb2y69r9WqPssvMwKqSj/NfqP
RZUnWk1WuqTQsMEM+yRwa/pxnLbZqK64/6EektvS56TGRUAKvvs8iAYs6ZiC
elNpqpM7nCxQbumMJPXdptpgeLSbej1wKXdU5cCfsrP86d56s2aYjubal1U9
I4PWfG15JHIs5jGE5hSD3Mp/9cUkAtaMJpKoajQF6V6nH780CyZRhWvedeWh
Bjjk54facX8MRWtyTYGiaVLnXLclE2ey9F+WBOi/mwK7lh/4mR16WZE71Unn
OgpHct4AB1UFMpCxWhECODzoyf25l4qoX4GleiAK3P6yBtPLGDb6P87XRA2/
SazU35q0BA7UQeM1vmmmm3lJ2EFEtxxHQMWeocNSNVRUPEd0SywLsHhoS7WK
b0fmVfP7mFoKMpeCgDMuAKrYkgAUrg8lh4d/UzBm9Ue/70Y6XVsmQbNq+EPr
pFlqtY/2ovKHh+w8vE8LH3cz/hrVaNTUJtrVZrYwcofoc8HRn0uoOo/FUpM5
623GdcBplXjgZ3cd6x1js0uBqjr46tLrIhQDyr8ooAd26Z+lDgJ8PB+z+CYE
Mdq07R33a5qjgBY3Jj0/KyZMTsEyUNv4Ws1ieO/OjyLG+YUwQRlZ39W9Qxkb
6xwEGfdluw0r+ifqPvGSb334y1FC734mz4kzUOnVlTCAbUvnGbOGIMcqeCRf
xMJZtcxhzGLEHUVeO874jltMLvywBIFzY89JWB0k6r6OXM5q7hL580o2FMKW
sEcNddXDEeX4fOG+RMwU7eMrahUsPzMo1d0IEcPkysUIqUTCUTEuYZ2r3kJd
4UCS9LlAiWOtfdr5NFp1SnMfttvh8escfhm+zGhqYHyaWW78NHTUsuYfcKIx
tJE1W1kwcv6LPiiOWyxRkaBPF9HovVFRoYWwMQm/ykPE6h/GmxnH2KU6jl9Q
5rVYyqetykHYBhYspqH9yZdwsZxkb16clGxVZj4HiqMzp4+X/JvDz79QRPqx
i1vt3QUn2kOkKBlQL20X/jakWiHczuXW51sVmfV4X3kVtKXJ3i+tm8/FB/CR
BRmltxUI2IbQCmP7I3RkQqi8TDVaOF4pSsqMVl+Rzd7FgNmi8Mbhpu4tQ4CZ
Ju0aiF1WZMUPf+SaEUjHp43x3yPAMS12i0WVd5w5RTsOIxjMfl6AcNtdB59h
VUnFDvuRVocza8eB0qsirmQHRzq8bm8r8rA84E8QH8yYK/m8nJuqAdVHwUBe
81cD5G2G0W3RHo2qy/HgP3/Xv3fqp1BzUS7PwmkD8MjC9JkeCAj8+YyDYxCb
rgm3kLNpDxL8zILPYzGn8NBg8f1F89vlZSGTQr/AwxpydgSfn+Ce39Wuds0E
32RFd0Z6GcuWFFNoNd3QSuTq6lno4L7IMxieE5djXyp6/bbghv6Uvxom3EIZ
wovcGC3ziNvelbYpzoIJw5cMvmndYlZcBpcjZdWVY20KDn76sBqgHvn+pp5m
qKwxWftHjTEt4FqwY1n0ZMUJOk6nErYACXYLTf4+kYqoSLmQoFR4LMs4luty
DdYRCFQ99xVHOk2tx5PXRl1DsFnbbuWCsyWwVzTu5x4wCmGW2BGuBlcplohu
2rpf7W2fwnqYQ5kslSRXFAxCoQlH35M66MF22CTMFeezeprQvtVQWtCuPqh1
yaqElYyhBIoFIHxJOcVUXlyCbUK9DQ9gu1FvpUSNdHP192i/sdaQKFsT2At9
/2jRt0Xkl03aJGCDR1r0uQx+3Ho6iufb0pHWiwRChMGNxuwPTMI8eyB5DmCU
l7fT7IYHxkOBed44PryX2XbkUJztSDiAjw/LPZgiPtQs5R/V/Nq+j5sqDqCy
Ln3NjuGvUf8nTsS2B47qEwW0wZCoU/nYfumh6iBfv1emMVr3tJDEdP5cMF+D
H3BCcSYvNTSrpmbmLWpvbPXStVyzh7PqFzfSPQnLGTxUCEpLn9pt4gIGMGPW
iBo6reGfQSUGLzZbrYI5FxgsHQZ/RwPt7G+2mH/524Qb4mZfBGpggslAd1oQ
I91dp2BsMrfH6nxQkC0V++rSBAzhDqBNeMfn2iI/rvgwWMNHkcmKvdiNBKjz
S7iG83WmkKwrV92gKhNGQOazEh9KN7/Zn+cL3rfIAPjtZ2SL5FLf06bEUiSG
Ri4eq+UskOgieMpacK4CAw7Adu/0koi6oGxUDnejYLOyS6JBdcUzQ6cDCcMi
qeGTlplyOQ7HuMvl/ZKHXDMJYpbVYtdj+qXGzFlhak9vU3Yyf8E010e3BDam
FrhnAjD7NhCH+Hp0sSe3kVPH7MT6m/enU1n9CI43a8qT/AsuddodQUwqU9UZ
KsWqkCsG+b+PqflbRq7AdHjK1jaTKSJFMoy7t8EkhBkIf6UxPOQzhFRvoRI1
8R9HOkKcvUpMA7ytbqH6CMd+z/hCkcbJFjjyX7NQTHNKFI8cUC+hWpvke5f6
Bj6pvKZMOssgEkqB35/2nO3eyNybC5uXYN2ubPcnQBXg1o8bwtQunGLxNMaY
7hw++yuEFAQEBd08591gPzMxDvPgtAILvY8m7CaB0XN8cliF08HPIz/xif46
vY7AQlnZC/2YC57VQ5j23tmWRfmnLVtrf64K31gsdGnzx/GBQONvHx4pjPIN
yA+JC6756wwemMU+bb375J9YBvcGB/IMpKwUXSsghK2W9dDxympJAEsLXbi1
DiIE0YBFiA0OqYYTO+LHDoLwbm2a3kkfubLup9C53R+8FSWIFPp0gfuN3Jiy
E2QgNIMKfCdF9oPeasg3P0BuWozV60IuP254yEM5JKTnV1OW2qx50n9v23Rs
gmCh/5tU67ZlkertDEQU4TlahovXgox/Pvk0dfcQ+Tynu52muiuYFZoDiM80
Fy239ERXufbcuMsB4ktcWA+uyfAP03DP31+9fU/78+xiBq923QYT+rASyWex
uQvmq2tXGr3lnmurPhhmTBS6SDEVE2+47nkISaQ0uWuRcKo6mWYxKD3OFE41
DyF+M70JxKmaqSs8SJ2JAdSAl4hAUyW6NE86OYkj+u+ejT5p0P7Aebs58VB8
0c6Tj/C0K2HnX7GhYm2inUj20TjNwLKLWsBuTr1T6eP/GqsSHsfVZZ3LOpZE
J5ahtBs1hd/I92B6Yfae5Lur3M/AHJmhTVodXA7K5S/BXAZwHmk7FyO+7Ypa
SNL3o/kmRRx+gax4jHIN8xcePHKjf57Pj67nhQjlZFrhWU+BJLyL31NCGqlJ
qPyuk+Svy2QV1mUsuHpokkkFVTnntXZBzvXBPBu2KPwLQ6iNaiyArLF8gQa5
O0tMtUClNO67qGrYZOlG2It0L+SfI0uew2T6ngXzrD+TxyOdxLkH82NPITKr
UHuJpzMlYoLK8c1Vc1eqcQ3BxB+MgaCOyG35Ko3YGwzp9QDAhQy87gEhKyl7
oS/3sb3kPyF+PytsZds10IRY3W15P3LD8gxY+fUezaO67Ua9/MkZseb+p6ub
cZ/0gZmI9A1iA9w/DoFAlOHWw+jWynPY20fK+ofVlNOPlOKbmMZ5J+bMABr7
sSaxLEX03eevFxhhsN4zS3XRALjWmx+8ZgbnpFcurNjo3VvI9FmAuxUmjz+x
kizT3sv2bqkwT92Z+mcQ2eiVlc0qtYS7gHzcHocEiG7MAk7rLhznmgdamN1t
77cDo3WQBnm6fdo1VuWPntHOoznUYGv33Zq6Tv7cuYF5CsDVItXYWHWdZiV8
Ro8N800q1HfU/1vhYUKhl0mfgbXHTmxzebPly89rhCnPZ8XwysfhlnrSeqcO
tH9vQyK046gjjtTmtWy4f9kcxhbQgU7OAHbdYv128tccuP4NUCmfYk7zp21C
q1mSFYlVvUgZbKUkwipxC7ooCKdZbq3QBEx2iG/D9waoF94qMkORtDRw8QX6
eY1njzfPB3dQ+z5XSxclBYz545xY3oiLl6rU/BfHf1iMQrLhyRDoCoclq4GS
Rxk69Y2xZyDX/Oxc+wS8t43d/SCLZ0lMOheoha8DhCjqPBfdM2meYyY6h4hp
soTNSXbaJk/LM3b6XHKUrMrA0orLRITmEm9BdOsioIq0RnbEeLiHP3H6D7ru
xPZpjz/Hqq4KNHnGdDZERollpjkPTsX0RO4uZlEGf9xq9hMHcQuQJJ85WdRM
Q+anfT18h9XENNXpd4SCEz3pF6fuAFEEe3dyUmKnOPoul0hVat6mSy+I6tLa
gWKxrk8F4e+QoHtUcurGVSj5mOysg+umqE8l+AcOhcGxfe1ci0fIP9MQlJi/
6zDv7EII0MnDN8UkWa4nljqWDv3XsJmZ8GNujzv3QyWJ0quyMh7bp6xs6wAU
yhi5uTVEMk/mi0B8kS7Gl91vhxNBsA2QwuocnmHFwzcdm9OH9GL7YuZbI9xW
LMV4M2LXYqG9TKm+XcBnjAi/vM/kEXcrTxbc9cHgriAFu7gCx2wNenTZY7GU
PqHKpNifuTlw7yY5aZKuIRs0Vnl5OZ6oXUMNVfruyIcdMQH1YAAxTf1Iw0Hf
X+briO6qMReuvCwSEH2I9TYaYiTxqkC9uuCyJr8OPJ1A/HjisivXojvaXE2y
X8nV6FnDmyyweLR/O51aci1QFqZn+wBDp9mWdduvGCIAak8yueiG5+wJ36FZ
WemcsO5M+9HvGU72YQaptmZAX1sqi+sdABtN8uzoK8BVsebqMsJwtw7yMO2A
L0trMBpMKlt8vEy/Enyq8dLp1pzhsJ3Lap6y1U3O1LAzwgGMkBgMWRV1iig1
n0/ltqsjh8vgQ19C+O0Pmyc5p7UZLD1temXbpIifI/pgJWG/297SpYV6bUE1
+ZZ1KciFXM7yV+JvSecPJ1pI0tlunNTKK6YqND66Vl1dPejhr6zIYAlGiAoX
0eL8a2CseYJqBn0V77TubIaJGwPC4nYELjR6PwRO2yAxqnmhcK5Uj3bzL2KV
bNfw7SYDVNBI0O/nu0a9ROEKX/taoTzE7tSVI95jzCfvg9yf/OW0h4Dldwts
mTUGeh8TN/LisQHAlc7UqU+kcHoJqEy3O0xalVnJk0oaYpPg+T8XcKIYhtnq
w7ZHljfh10KWFh6CJQQFbQxUH1ihoQgBheRtJzaMwAs5wN7S1Bdlrh6cSP8T
1f/hYczvQCg3TK26FynxXkKAtjishr6Z+lMRdC/17WMfyXtd5lSuGWq1l6xX
C7c5bJSI6uM1ETmMsGJK024pBpOx/BY72cjCn/FrWygBGZUps3FTWXRV7mLH
M+cEL90BBFvGocwLphs39zpfJ45WxG54+Y6bTv7I0P68jnGPykwmruds3onf
2TlqLmKEgZq62e89p9KknTB3g9FcF65nX7RDP7avg3ioGAj8o9jHcIU/t2ZW
+9zU7ptJqbu7CfTqHqFRb7ExBQ2NPpyLltM9BCAvgie+h5FU+TXjTW4+wrAX
qhsSGDxtYWAI47sn6ndBRL5hlH0ihBTNBJxN8Dxmj9SYCaC1exFIZJiGjtyD
9vpB5vwE0Z1SKoFdWo54P5Xm8EYjz9X8qKLWP9wjDW1ljZ8Q8jbDsuRoLKSN
SpA83RTYAgPx+eDTatIDycjrANie95qyPnJmJL7WjZVrBeq6TSMJ9O8LvFNl
NzYzAFstbOVzUbrGmAGoq+AzniQsoLmujh1b/M3THlVY9jrNEQzrY1uMpaq2
05GkjSQxw16HvVjVFyvgONaA8eZJHAxFLz5gjook4t6HHbZCEjnVYwp9BNkE
F6bzYh+83dq4zUYHzOWkQNBZvs7YAh8+MVcS8IdTKzLtaCT6UBvPX9OZjheJ
x3ppI/ob0YNyxXkE0g12f414G04674JQVn9WN9FVQATUvLcjn24eDr5//kT6
CASJvbRK1Tj4T3OOiYJrB20dG01o1/MSau3u2ZIaYM5L4NXieZJ5Wvl9hXUY
ZTOaEQPf9uA/8ES6rUPFlLiSHCOaJvn/OISwwINC7YjO5y6r+v29lBkImKzj
O3VxoDCGppOl/fa1QsCqt9yX/v8edl0pb/HSw0xIj7fkvBj2W9uddAtjEwcJ
e5nNxW7kyqVQ2xpKY7eNjCLELixvdJeM04Ywvv1ZC7kJOeY+j+HtKx4hOfG0
rgPlVWv6xa7e8+08OC1SnmiqHk9F6yKqbM74Iny8kN22TeVZ9GeS5rJQrmAS
Vg7B91LDbCHuhUaLEcZ3D7EXqKjmml3z8aB1Q2VwcAOtqnyX0+KFbx0vocVM
wMmX2UKypko5g8dDIlE2y98zy284/DJXs56wk4Ppjb0FoxNZ1j7qUN0BiBVE
LO8SbBp0C9+bcEPDg7CZXoQ0dRFiaIKl5l6hnN+tN5lTZl/31yNTzOC4+iVj
3bK5aYPKh0LNp6Ef275tjSFaBHscEMOThKU1bGSKCv3iUXBCHlFzXLRQdhrO
Jn0cU2ca4Os8qHCiGrgwR9bOIBSmHdVT1dvj4Y0u2mdgpBBX0NPqVlLbZj2C
TClilMRKX2Io+8BudRbYKv9lSWAx7JmhU/WDr5RhoON48lMygRCjhOQogNLL
XjcmbsW0VTPKkVsYxHgM+1N/fA9S7KjjUcYM+VebQvO7pVr2fT6q45jz3wM9
4CI94/+D4CmObWF2I65YtVpfE/BtQPMLcsgKy9iRDCR+Flu6rfnhz5sF8o0u
6SdpD4qodvUsDoi2fJzQBLSEfoGyAcTZJKTYuUMJpYhupVNvVk2DW6EDHojy
NbdbjPdyZMm69hQIBg+1wmkh8aJZ4cBbDZ3G/IRfclbLyrD/uysnl1xszE2c
fFy1PTeLMimQOKeefS0dCmPabcUAne/IywZtWBUem6s7M4yGWYCCT4ivnEO+
6ZHJYFf51KJ70AmXauBOoiYiBSEplT9k41ZQ1tZCAiLClBqlb/NtTIv8YpZv
zX3AJ+8I8yTPlFfHQAnZ1JAa0GhhXMBe144sQzTLzTdFWvxYw3p0Xq1EAdG4
/vvQHVUAgzSdvUKSBNT85b+uJQXIDiMz1gLEKyFdY64uSwnwTXKSeru58tll
y7qey7XYLu+ftcQVm9SMvBP42NMXYB/iV2DcVFQn94SR/KRjQ3v84OgdDUqt
Z8VAxmmN7jZTdU5z9c7rNUkMVzOdWOx1Cz3WqwE/YDME4/4yG4sIPQvz0WQs
LXRsqNEkZ79c2BlrHXAYcz66Sw+SrmuvN1LTXD6/eqS4ljEbjreuYSj+bBDd
eNRLvax8S5f3ccBWJxb6RzTBBsxg9qPm1YaynlhqDP+aavfNqYzynAiHBy79
JMuC0CXwXbwBGAdNtD8tmmYoxy5lH6OUGWnLnSXN1wbyo/QBgClSOF1y5ZiD
k8fjLIi5/DdA4b+ZHiTpf6/nUelGz5n17QPxYg4M6sB4qLvtG0jTH89qxMcj
1qCIZ5j1mej7tWu3ZoYINB4voAMtWVzunasJ1bUBBsL5Cgw/gj0hAOfMfuev
kQqi2Celv/vcuO0hHcvstcM1VjOXU37psK84h/IUgb4AZyqDxBaVUElbsHDE
LUTP1cSRf/Mz5doZSlBprx/0SHgbQGEhxSzphNRHQzxfyUdhMnFik1TbZMiF
09EpCZqsaCgA0h6v6EYZeSXa+jlOS714RIXuyFs+Kdnf/A/NRVH6+9loBMZ1
5d96ruoziCjfl4a7Srp3Pnghofnkj5N4ygOBxKTDcL+cSv7Srz2KP1Owoi0M
ygnzy57zi/rfL2DP4A0dlB5wObzrb7EPzlGasEB5wRMHBLmxRyAD7Y6ZskE4
f04eVaUfHdDXrlT7u6CIAxRMkgkZE5B+GKffIj39BmqzfE7i+074chHSmDSJ
dhm1qY7HyaGlUncjcEdmGvSpSbQQgKvDgxCegBcRB2WNrgN5dSCG81tZB8bF
w4n0h7RRficXkkG72qKzY0mZgWJp8U497Bxa54rU1FoWvK8Z+IfXkAQYEVnr
00vvMI0Dehk4KmYbRXfXxW2ONPnkuqIk5BxDeImXXOOKh/FS5t5HCWUcv6zg
3cqf6zGeTwzISCojD4oGUDfmoAwKmYeOch6VooTX5MsEEQt5xN65W9519r7I
b/LAiuT8d1/4D0luObf/WDVnN9qGBKq8KdX6IuWJQ986tbJSf3kG8QVyHHw9
Bq+5d/F+pzNHuNHIsEf4NCq6tuMbVKDxvn6NW0odLqpb4rEhNM3mmktTgkSx
KqCETCvQagJxgN6DofKqhVSK4dDjosEHlT3n3BHsm1mJ1sUMIvpUHFlPEotr
UtgYhx2mcorLzbXbF/sR3miwsa01ErQmLO8OXOh2rBZHQFTPzIDai/7nbhty
oBCwWV1xokdv/c00SAmXQHEKvtfhIdH1pQssMC5AkQ/LjnDjBKwHucBVOifS
DR5S8yriXl+5Tuos4EuDF+ZgFbnVWfv8NtfY2/+wLzbBUgmY4+yBsue9UrdM
/kEhchmeGPFo2KjrjVxPApBUXCXJX38cC5td+oZ9ePF8syLTS+piJgV9SzFX
KRXLh86PwOa9UXe8xpGLMc/rkcXa7o9T1gQOCwJy5fW/Fg83Yp2GxkSQ+0oA
AA/Aqx5Ij25JKA1YEWGsCUewmbOSl7lGbxF3TfKbhFIB8R1PhxJux2jytopJ
kx5RSr/DyASyZK6+tAu6pekx1LrCPA8kSwok0Q1lkY0+B232mLyXHCCHdFvR
/h4gYgHoXE3YeyM5BJMzOJWUNSLQoBP0LsNR5iGoXMRkNxSjcE/rekQHyHQ+
PQDS+/oU2cSoC6suFKglRN4zkdwq1HAdQB0seYwq3e6oZlQpv+DxTXx14xXY
Jgahzu67iqmDoQyk0WrQjVLYDZgmy3colGiX7LeliS9d2BWjuJx+MfSUC7XF
UbYBgtXoBxmlfYk4qdSoJXtK8pu32kcFEreOaEmtn1bGu8JXwrLBNX1NpAF3
by/os0usiolnGwBcmWGw4YXqf0whzjic+JVXc3jayWG5ENKcjogdB2xZdyjm
Va+wd4HD8TuuhyebTXSirSOF6oRS4IyPdadSW6ySdvd48oK9X9DDAEVZ/pMV
vbWvpD3dFniZVRR2cYsY/dP1PiZsivoHIwR2IvCbTlE0L1BdX+mWcz9jkYt/
8d1Qr+0sMDfUx9tKarsGP4ptnhQB8rXvZCxvZCGMOYhNDMKWRn8sj6HoPA3v
kYmhGnz9cnk0VsDs2RJKUFtWkqr3F6QAguoEigJonpRATAKaKMlvBiXHkyla
ifPVlokYNMYk9kL8ifYSTIUdtd60Bj58W/701V6LBGwvGhwevMJ6ReVbEnuG
9ZkaoBpdVMj2PMQxLERqDPuxi7iQndbFOlWzMPNL26jOKFPLFPNZDNqmUR4q
/Lf0ylBEh3XD6bNcUyQ9wFa6v5tKnvN7lSUbj7lpJixHIg+UF7u9XpmT/Exe
qGUSmZ5PxS1Bkr1C/MadrYey+y/Pc4K9df+F6iIYGSpy4ohUMBtC+tcerveg
HwRcG/whvT6y6qpie4joRdNyAY/a9SLnInI6OY9nJTDPZ8aasuLknlyLc7uq
RThLQZfMSYNvRNS/Y6d6HVl0xMe54omMYPCvVdmCoyTWewIqnxgs2j2eZIry
rSlFT7K83CHwHc6ydGaML8L6Y/Qgj/pyycKJ3OYHJ8s5F/9fY9KCKSYOL8qR
uwBz4ndqXnMCGVQdLwo1J7ZTVPxFIuC1FqOEwANg6rFbFnmje+Sg0G6y6PMR
kCc5tZv581aVjs4Ez0Rx3ykK01uaZ2Jd22hr/MMj1cEv2/MpqGbdQo9BPMol
VkSVOrBXDz0fHsGtiga4HBzuhswHEM+i8Q2smBLgwHpdcvXDsT6oSLMvc3qq
yQDm89iR/yCl+yydekPRtOn4rAXZ2KBXV240XXKaBa1TFOcu3VfhJdA+eV9m
06xJ67H04qFEOebsdwdejm6xcFLddTWZR8sPRqbb/aXbmPz/Semb1SpAES3y
GbigTBhkQdyhiIqp9Jv7IYIdG3aiou27/dSPTVbCL0qR/hjEyRokp0vCyZru
+LX4nd6vnbNK3Yo5YNhyo6ph9UAuQgwh8b00YWxjWi6fva10y2sK0c4Y6RzL
Mh2xqtE0ZxcIvueodcPpePx/0aQ5QqLbvRWuZFf9p2NGl9K+nmnvqGdkkBkl
qpwWhJGv5HoHbwqdnVWC7pagXJKxm5RSXEU2XSdXG0uevdlNR1YsC4kvFJUa
laMV+5rbrn5tSVlBtRgk2MJciYJC3Oeijc/1LmFMOXxwuCOz5LR3VaTVJM/K
8ChyMy9+Va7XfVY/WDuZER5Ldf5AlGFn6fkAy1GyKGAzJH3gqXUFYH2Rc9L7
7pxprOLCr3qqfCLqYpl+nVaopcxaY2dq2xt/oYHmj/yccfZzCldBhuyVR0Q6
J6lwVzuMt8G3sG+h70uRxrt8HwXsT+a6VXhN03iFME8fab07rVVV5M8Es+A4
nRDgXT8H48QZeX5u6SBxpY8YtvS0LwYt7Gi7FHb3DopQN1efxlXh7EY9E3pq
IZQxxnsqh1ZuS4NIk9LM+7+9qbCfsQJL5uXMXTATnKiix8ApYH30+Lm62P0D
6qJJA+wqRX9SgycykfQa6uesMw6V2yBRNb2cKEpbd5pyLCpIIb968MwHrKNK
6PpAXTtbahF+sk2Dt8vPmXKPW/bNKnObPQxtNf/xOrybAaRVK7BGEmaeO45p
WDxS9+XJ2GlapEHgbOb5GDWTkBPlB2Lj5yyRsf0UbXZvslQsGzVt1Y8MjcZI
9HOnNgbCDbOb5vjmYKUqil9N0gSqV5XrLljGgafthfNeGPBSHyUMYiYpDCch
oPw/Qz779/kavGV8s8o3ZeoQPSZNBdmjclhqeP3ILWiu24Qi2EVH+9+qDY+/
VXd+M55l6zBYoYuj7xA+J67FAkY9S58TPV1SJGVDVxrh570hUUsdrdWIpQkH
C7n1rdGtG41c2GHMA5UJ9Mas13POm59JK/YkMLXkzP1WTD99ZLvHNnFHS2dt
3f/ZcjPjxjCVYQvJ6V/9DWd4AoxQKYGGcPWOUyUVtporwb/THNL9vZu0c1b6
GzPnbVSsLA73HvZxLrCRslR6+Z8fmJ9l3UomHLmoeCotKoQ4d+xwUefrv6AG
lLExT47zCyxZ3sAaoF2ZZ3ECJEYVxNahQD8jS7TKVgK3IxX2RDulCsV5UZeU
ZbWRPFuwLnKDCL/O4j/00Bl23UQsnQuu/a65bkGWOlRRxjuhL/hwun3H+jR6
5ZZ/0WXhr2nwKEe1Q92ywZJaxQFz4Rbi0v8DIApzlvjdU7nrS0AUPrI0q2Sj
sq9ZCK70GcpdvuYg+KaO6hv4J23/tyhi/26RiBcx+KTZcngdjZb0HLUWNg1x
DG0wxYh7RLFkrTjtoKeTcqKCX4BHEDoDJTEQQqeE1v7BheMJDzxPcpU8tPit
m5+t+i7FXU6ceYu+RJ1775lIPbHAHfMXHusxuUp4sy4amXl0aHabPi8f/qT5
Qfe4oSmMFvHmsBMpfWBSJk23CBtPDVJiXnmOjcRU3MOSTNv0df6Pv86NApLZ
2iMVTfyy+lTbLqpc0/oYcQdWtGtLBi5JGlcZdkW7ljuFcpRVTCAaPqZrhJnz
6P2mmtNhoHGnym8sIt2XjzskzR3l0F5pjtI92vVTTbl6ozASqczCsfpdiyZo
svmSa+v7o3OCVRFYLDNHcPSLs0O8arMcM1U8yi21bAqupjATuFr65b/A1Aj1
npNnZQdA8DS40rl8jnxNwvIg3AVq//UKE5y+77pTAYg6k6WdDKwi9ublBZee
E5CG5zAOGjFfhXdhHe36kKxKSzRnKzE1TyHfc4ioL4z78aDXHcsVNVIMZ0DP
SPrvwTxU2AQkRBfDkBqaocfBTW+m5fPOqJ1iRkzyyq8aoIKrCYmZHY6NXOZF
QVuQ+S0PMUjxxPeLEcJoxHKm8IO6P/YiseUheuoddAQkWtTixb4GJuLLHZbt
/IqDrwbYw6b+nidZXz4sMZctM3RTZnSolZPSGIBXNKusk8HerO65qsh+JSKC
DCS2RIYef2N962tUkFYsBluQelLIOinGhTyIjA+wWO6gs7B9HUjuKeRA0wv2
KexZoLyT5S6UmX9Pn68Gc2A4+RrlzN0N8Bd35qYZRGD1yrXByK/vMmcWPDQS
Y3dCDparydQI6AsQd9OH9BNiWz59YUEZUakqqWCOZ4lvXMHBR4M9NfBCojbe
RGG36HapjB91wTH54pNMltOaqvUOMIdgba8niBH9Or4VRnn20QjAgmyrIngs
iHWWV9p76XiwtCJNXmk9MPj9gqGirAGQkkCcNwYYcSe7XX98JHlcTvytqE/O
OBfyQl7GP8oWT8t4t66msyupoHOQk+bS9xO5DLj/B53K9QSJGLRkYFU+g9Pc
9kiXyFyuIO2AAJYNZHsZT2Rwq1qcxzlm6canfDPi+GDTMNaroeXDyfNpNZLQ
4Ny2cvOG7vlI6AEHpaKoNjJEk7H+416MhOuInpHKKjXKxZy3WxPPv4kjhOPz
BSwCNqLhqq2/uQ2pJc+v2jK/oFA6uZkh8EdkgBHh6RoeATBMoPwZZP6KD9gF
okFoHT5Sy9VbHtTy/JD9b5TDvwVfOiI3Kx//CCpslz+7NNut/AqUR7qvVjMk
FmhHe9KBn6CDsEZAmKxZS4J1upFhjrBrqf/bPq5S+EynwNxan704q0/GNlgc
cQDspw4v8BiIEvyna+SIgH6JIJ5462R1q9glmjqDbSB3XZ8tLQKCFRtsW/jK
ryemG6X1s5dWX4YprCnG1Pf7XDF9m6h8c5I9LyZ/tGdL8PZeGnJDk/znPtfV
fUacyNLp3Df4p/JAEeWbGjFCxV9mPhQf3kTAi0y1sFMtlaUQV+kZEyDOw40u
JMdJAzZhvdacG7fgmh4ZayY6jbfbCsQOq0SBDe9oMb0Ra9dnIHu6wYA0ZZAX
eJqs+DOPoJnGvnxOsWtWEOo+58aC2yoPu1dXTEuuYR+HPSj5Ib1xc7BIuWfb
sp8MeXmw3DJ446+g1yX+tIv7H8DIAH5PXViJ9xuVcII4/ZdEvbOI4ATn79kK
roDElS8G3w98TEWDEofyiDmajdNXxkKpJvMq/Bc47fPWwLpir3H964u3Aq4k
fLVsDfTdwUUSZ9JpG7jP4T92FW+qvZxKsTcFiMlOl3q5ToC5am7xcfa8eRvZ
vTdMv11Khz8ADJW83vIk43/2p+QJZmoUtYCoKstjtBskUbS5ryZqyiwRJFHG
6M9X0kZaQdWP65/xkIAlR/JaXSRghDyJ52N87ZUrovBFxfPmh1zvtgwQyzE2
UVnnNoyqq6U4FoHntQGvNZ7I4rmdv8Ca9pMIz72RAfAUyvyss9SDvWJP5XSj
drvSYg/u4LFzaOaJMVPWQIiTDGDkIWVZYzRL5jjPyOytZgP2oOMDbKICXlZw
RSf4XfJyO5MYpRGLBNwP74mYTS5jdKYee7tR+4XNAQU9bddm8FVcd/ZLyOvo
kfyh///JXA6RjuPCdWS1v50h5ta53g8i3S/QlxbksJc6PLHzp8ZplSOlF22T
U9ss2LmtkgFSajFh8cX5EeXqYCqytlnshuukL4vSFLT1Vft/K2kiwAApxNjS
jCJXb/FqBBz+hcrBilVn3ciuzq1PlKZrqp08t6qej9nylIpDBKAJfguM3fvT
BI+TcMl1QrGyh2Y/CU4bcxAiJJ8lPKbV0/7P8tZcXm1sCKrZdqhxlaxjm/Pz
mIDQa3ScIl0zoxvxxY/nldsDGYB7sm6LSdrj5SMl4D04ShjSAhErHAX4TufH
hrOBdDFk7fpuI0bEcW7wSYERe2PJbovive1SfQk6oHtkQeY8rDAlIl8VyNHL
w428Twpa64yV8YYB3qBsn/jHBAubvmSsRKhR6DTTjbrfJUg/D+7E8uOPKXUj
xYm2mZUHRizEgPGyKkoGN1dd9BjJHK1WBD1nRMYHDCJ+DsJRUTK2AuLaC3IE
4GRlUfA0YGUNMkbYa8XCwY5FPZ6DYMQaS5sSMskSM2RsgCiiGTxlNZ/KDCAp
3FMSCNOiWc7I7fB88d2MtjDKSraW3yEMXtw7kWVYoLSUoDOP1y+OMgJdi9jB
tmeS9c/0lQjpy5UhuYB6IgUaOSNvYX2GXdsyVvVbDaTPmvz3/W186G2v9Qhn
SmPoS4Cj4Qr+iDuz8P8ZjFD73sMzEfwF2J6gkqRsnBT24o0JxP6ma3Z6G0qH
Qbw8efET5fJHOos54ywhH5N3/yMvY4/FB6QrD4Ll6EDPnW1C2rhEoF6w7nJt
BmUzlacDwH5ztFBFqjInDKK4SU2L/Tt1f3odFqAp/NuCPRFPDJredFkXSxEa
PH58z6EFbdCHpqYh7d2gCxYFrlz+uMWPlix4sOCYxFzSwWHCVqIOszyLX1GU
G+L7hvNE/Pt/qfP2OO9Qsk1Y1Z2g7msnO3CZgYw96+ti+cJCp3KNdAQKRhIz
OAsvRVUy7MMSKCUP3JH1oGk0H4c3DPoAI9vKyp9eVMOJkzKNrYkaE5EGKcpA
dvX0qQPayQOvRC/T7eqdCr2bdFaReFsjkhs7lKAChD5nWuuMGlmmxgcRkSJt
qm2fWFNQVYceOJKBbV3zLVNzT0qGLzZZZqvKffJdGFE19/3YOaROorxGb9+d
yzEpb1GMgxgmcAXvUHFkIhlGT+HR0DIjkp0T3IAfL4/BzDrkPFocXpbATlZd
Z8baXdiMLls8UySDvODm/PVhWyKw+pS4kzg4+T3ElKR4/gTye3AwkAV7F92f
RN5XP55ni7tNxzUD/J3k98FMIqO58GChIRtGpbujXkqvsvNyVef+pNKIbFL5
BO6oZ2d6yKlie/h9nEZM7B5/b3k4fZhyxy2EAb5LFqcqOjcjwq3oRDm2JkWd
EPq0JYBBBAFLxJuOyygErK4iUK6k11P41+araAOr/8sT4okf2twFx4RTEYI0
6kHrBmc53qca7UNXaCQPIYAsZMHj+an3p8OX/GeAum5u5DkUJfSBviPfs2Lj
T9LbvmFr3vB9/f2OsQxWse355gsEwZs7dkTMMy3AUbJDV+KLv3oNERpSYhjd
WEkgArBGCnOKL6goJzjj/A5byo/4DNVwYfBsi4UYnm5gKg7RGgpsuIX7qRFn
MwHczfaqMTSgNpA9Xq/N3hHEmsf62Mz4RnnLGfs+DTP5uk6Hl+bVFjcRyR6j
FAYWpDBijra9eMpTh2Uryf5YV90Ewl9VBf8CC9D+ZGeRlKAVTegyKYt5fzUX
a5hatgY7jc1Lm3X6whj0BRdG4x+bHVlDuZlw0zf45GkdNsyNMl6kwfLNuJKm
xblmxamjGHeJBCgZkioLl6hLctbXzVustGSRxVn0sN/8tS0oEOtHmIWOklRv
8nDx7UBEkyRoNODvxdk2qh80g3MxtL+TIvk8tbKJBOldw0ct0/xf8h6FXCVN
52ApqWUgEPFteL1xQMELb6hJvAsOqiBwWhbJqPUGZmKitcm3zq493ktXHvQU
sjyyKVG8rsFsXmzrf/FMNL4PyKksOklXzg/F+LesVqPMTet/GSZAdIHmcJAP
JI/IyjmrxJEW72y3BhOQ1MtHBO72GEN1doTawlr6tjBVDAYXX6o8I9z1e4lQ
EjQkUl/Op60BQs7NamVWQCnu7LRnwNblpdpgHhHBu95SNjL1hZKLlJQaVli0
+Y8ZcXzmYL94dbeYVlFsIOWlMFcR2OZoXHbMQTzmq/fptD7QXWOYX2MK2qlZ
/N8YwyLtHl770zpT4LkGuYHc592nyk4MBwo11zGetd9+17p5siRSCAHjGX2g
jhY1OBzXfdcXf5XBXzB4MlR1zyGpOMqFx4jnAtmLnTTYQIkgL7TDL4VPndOp
zQhWxIO93Qq3lX8L/MfL4v0Al25ng9SolCi5aoxv8k7XIVAX9v5kpTtND/2P
GdwlEchY7d/rUXcql5mKRScplptub+fY0NOnwp3pBAii15U4+e0xDz4KnWuF
frxUe0Dazw14NosEZRFK9T2WDLJoo2ZdYOIHholzJ91t8tUpmeFBZo0PZ789
9RXgO36CbzkmD5vJYxGMLjiXDa7uLjxvrlR6sV1LrRjlKmNpgiGfwSyI8irl
5lLW5+WhOaXP/9gbre4NniYTMTS/jX26m1LrnRhP38D7mKs4+NlxaFhEWiLw
zjNWELSiiy0sTOhWpyjV7sw7qY3XzbgbsNo/VN7ANKIUugkTumsXP6MHvR76
/xW7ArGP1jY77+8xeuC2qsmpnoCzne+SUYqRlMYwZBpoMf/9SaTJdVDxOV8/
uJYqSIhNNS67RS0A5Okm63teElVMQozkC3GtdpmFb7BHfPvpD+xrmLnnpQ0X
lRr1qAIvbVnrLJIlyUyA+SJLvc+s4+mtjF4jVx6S98QiuCwLcY+wcgXssxFT
hS+Zf65WJwmTJ2og61HZLWZOBwVZbC/3jgjmRq6exSlfarZwmLtFz7w2mSAt
E2G9NKk/yRVrpxnTpJ03tWp8zwPDMYDrY8ZZwLdaRCp0x3+ko6yvGtHAfSPB
JVogS0PV3HBOWXRqygFUHMUtPCOQHW6HAjY01iOQMC+rn22/gaAWGjDuiikB
FIMzxhV0u3QQmOKaT21xDg/YW1gQzcueVG1xo1QgedMxDkn/up8lSLFnPVnO
8n4oYRM09mmgNMihH3R1XCvEovSo/AqAgKtaw81o0SOHGvwKI7TruouKwsHM
ecN/2WnaWPk3tylVMYImxr2wqJKe0HBJyTX51jRhlyoniWJjP2AtOUQDhb5T
qGxJq102oRiu109vFTwJH7LaA25KF6XVHBLeML60DvotdKEkX1nniscTJWem
gdvUlNih0SLlznmyqjJsuPNS51MnOf7oWpUpcUEj5wrxT40QaC7HnYIhwIOC
gsGoRiuum90SgkgGyIyrt5/xz9aHe/U71qPjl5F1aCFegAJZz2F9TtnloQSi
94Z48ElTh4w4fWkCF7AOeG+by/ZFUH0O7GLnPSZFDkQMR925A35CW72CaRzj
5hBYa8NGEetgqY1lHExlsq0+QYMEXhn5QkPGN4ApjPmsskaUQNj6VPF1yioj
9W+02H1evwYuNRwRnyIDBnpSZfYZDvTeotZ4caRslN5YdtHYuIViAhm1DLf5
5p5GG5XAW8V1/XYHzhR9H1+XlM5Fp0LXRALWDQz4JVysh7AG5fiFG4z6gREX
PE2jqWiRpjRnHIn2kHYpyiJCNXfA+JMI3VdVfj8ctxnVMj6tB6Yd7WRTiU+A
aBmSt0B33GGZ9mh4PM+oBB5NKsUYyQ/vYYSP6TFfwl0zUFdrdu3zYrlBlWhT
ljPoSw8cmYDNl0k/Z97kuAdGqTLbHBIpsie4nOMhYOR7nRGeepsmGHZxzX/N
L4/XXlju4tu68u8jfInJ+uUNk5S0ewXvrNddV2enwcG3bkn+COqnexW2QpWq
vrptueeXyJwW+crU2x0I76oj+Iconvf9qWY2N8EjjzHeR7VCKH3gHYeplnYX
KySpDc2i0KihRVrJVIbAxnVStkn1qZaN74myFvOY/O8GpDQWuLWJWqQl4tp+
B2HvBOraPCyVxmB/n6pgFNjgPrF24t5TREBLlDfu+psJnjkS+C5CelUBai6s
EM6HTuWPyhhdZhZ04f03l50HYwMIXxDnS9hKlS+SO6052UECEubupSCTGg46
wLc7zJc6vOIDJKs5ODCpnpAP4wB4wjJWoS8TBDAczfv0KSIsucLcH+Etjsa9
AsqhKuFm5K7NNfDljdO83d2/2SrP0zsfIMv9RGCP3fQCT2nQY7fJo4ikdpDg
mB8E3itePnDOfyySioj6bX+jvDs/NLhDPON+tueAM47rSc+Apfmn8U0x4qMi
AApRJsjzUXfYat0GtlTWw40q4a/gSQjwPOtSpHv8LPTyFHLfEpmK4eTYWElQ
06sw6G44Hmin569g11nHndLmB0LdvFvzYaU4r2lCnIpu475KqkN6mRthu7Nl
hIeZlr2EvYQF3BMRcqOT5tYzlR3Q6iZQJIYAl89ZnH3ImDg8dD7r3HCGPrzk
zim7qU0oY/Z8vemhgyjJdH/yd1tWa9RoQzzlTo+McCmZPklxy8i0MQCe89sp
h2wm78+orcdXaJPgC709GWdTX0j7ZNu39HPQ5SB/tLQQP8joeHMNm15xZDFq
I+dTAP2qkRC9Ad6Ym9oPeTb71hMpDJ90Sn8usYQINjE4n5ey62FDu9y+1e0/
SG/r91L3DZ47jWLHcY9j3h4/Hq8DGRWRO8YGjOYEIRbtnkybDj4jcNe7Mck0
fIC5HA8pO5pt8AUvv+FfwpOBwLu+Xy9uJ8Lq4VLUCzZ016vyX1vczlKe6A8s
/Y3+Xb/IyOUUiEHSNFVHLb8KcgZGUKhyNBBqelLZWRLFh7dL6YdMk3wflepm
1JapCppOhol/iNB1BMxJfiDyBsAUnx6OV4DqsoCs7BjU3sdIpSHmH99ejjVv
DsUYAMkql1x2kcWX3htIV6gYYZ35908jXDBb15Qn37gq16uJAAAd7LpdOtid
BuObXZfXjadIPWNkVkNogzTb3viL4/vo311XjFPAghkUKsEZ98b71FmuOWG3
6cJbYhnhqFZ4TShF6sswlzMyFF0hrX5zdjO95vF27OK+4dHS9EVjSMbDENM6
XLLx/kQzN1SxtC6X+N4p2arz+QgQ5SZxgSLVU6VvetcCHYMMDpUBL0dvfn0Z
8uu4jTLVY5jRxQa3i86yCoNFgtWrckcX0bW4zQVucS3Yyll8uSLVCb+sfI8m
d7rqbGphpu/PMDBMrCk9v8aPaD17JrH8ZFg9NAdyiUkUB+2NizBQ5nTr0Uro
HfGHJtNeWvbN3/iVM0Ca8E4lZnJtWDQxCjuNMbwJYSKQkqho30GNhwGgDEpx
SDkXQTpYdrmyIuheOrjVieAEqxTqoSwRj1I2SJ4jK+j4AdVO3FJP4U60AvKm
ZpBsRWRfCmaFYdCuc4WVtuunbNe+qjdYQcSIgdN5kMfKvzkyxegScqJ3JUeN
A5Q8Qe6Ac62pcma3JzlUCqBk3TZRmSfOcgb5zfHX2fpUnuuTCY0QGefgc8+j
lN2ziFPRN5CeVoAY7D3e4nUsPDnQhwyJs4dP0qkDFrxCJ6J1CZPbWxHJsQPr
zfyzVO6x0vObiAxqHfsEYyg0HPE2/liM7o9YZkc6GWU7fOc3SH9iSWP2SKFv
/i1UiObzcl2qc7O7pCvcEOzq0WHFFU6b0Cz0J8D5EHbJFDNYTllVmAp+6+AQ
yWcp2qCktMUYRvtyEZglGec+wMu79iFotnS4WwWNCJO4Hbdb7LuHDkihejGR
kOjza0mW8PXDt4Cn1RVqDGhsaUzjpCasjULvdzZVKkCBH4JJXCuY404Kry87
Qg4t5Y9yDGL32LF3fE6bOdzNsgEwW0sghRVvNpmhFeG5Tyx56gmUGHwFjyTA
iYPgGc3Ly4k/RjFZpF8vd6O99eHXY90cOzUyrJonGyJJNi8Q8dDzq8IzVGel
/AxkrcLfiaw8bqq7AR2/B59blkOqtKNttVu/AzH9TwbHMYgAtSuePQFwELBx
8b0U7aTRRTyLe3OHXmSshuhyjvWIYDikj1G8xY6osjsCLhrZ5byicQQdkJVl
yRR/uCLG7wi6RAdXDp/W90BO7MViDamYqBJYyKGknzacN/iFHVh0tfm/Li3Z
3bF0V5eXrLCu6Kbb+aoc+Q73mhDIveICwYpwafIyZqJc9B6RV9TJfnHRuRHe
5TfJVW6MpZTPwMznxskf/GXw8fsbvStwS7bod0hjoXfqYkv42cM2PbEYx7oM
QEiHl2VcjBkmt9DKfaqipOqVYnySPvWvpK7oESaC+6Kb0vncIRijH0ze1Xgh
wAMpW/s5IRqMzOFLn+M2DztxSSMRNVU+l6zJmhMhl1zS/eRkODSzJ0nXtZIP
GFxss4hbdjAZJvZ+lhTp5B0T+SgqyUr/+YFt/Ib8nXCnBNP/uD4r16gDSjkd
5zR/3oZIPhux63DRIIVeNaibqV2fF4cd/hkRv2q2a6FP91PK1xLSlqTsOhpi
3AE4e832mO1rvAS6H1btTt/CImXRoJE1nIfOWvnwrinlI0r0DY7y97xmgmSu
np6O0Ab3zi91RgxeMa5dUvR4LlYm3WizJtQtzjn1Bh6hNy1qMfKE3UmwW8b+
DE0dKxPExWPRSZ4qzppiM4LevSiBhVQPHEdTlko8bzofKLLLp+01o8SzyT63
rNcRVko02nZTBITXKPn6sDnvbqCLkD3dT8O7E/tyJwwd9KWZqfpVSgsjD2pK
p/DT894oVXspAVjhoBF6NSb4k6qjMu09U2YAmHigVknC32khsI2UcdczsI6x
8Y9Ghu45hgdCYYETov+RNQta6bmHeFMDMiL6N3xSp24N91WriHogyMvLULLe
Q7HQrikS15fEeWAFSbKw44/uVqSTnixR1GNOKsg4InUFTfodxbbgKDj5pyOH
dj1V85uvj7GAsTB2zO2MKc1C+heVKCatBsBj2D7AseBaQQdc7WZBZYba9niB
WSGvVhD062lh72D5esEZ/OjtD0G7AoPieN/adz1oh+n7OZCfX7OoXY2Me5uj
pp49VP/iYWOpaXlwmZYsx+9cADazr+6HMIssv7oKEBGYWYjX1bpoa2aavGWD
oCvxz+6ecZ83hWmDjXY3Myrtq9y2mReEh6VdMMcnTsmNrkiUOnM1oNUwromq
At/2ar7TxR0xizJ1sv2Y+BPdAj8Ig/OsAr0mYvux+680llKS6CRVs9F6Vxbh
s8vcWyaeDei9ow2uA9LlkFqtnLraats0bxR4epxwoogk+/RSzaYxa2syixND
Was+VN9An/xDtn+P4NJQLhzclRFykWOQMX7x4emYKMRflWBZj3M7FKicCHCT
SLjYZ/YM/TjK9yuk47Lh9dP3G9LLP8JInfzIkow0bsD1703fIuHaIhGjWdIs
+BkIEXUEgIHFoPM/DoGDcn48nfexxSAWMwcbg1mytAgl6XnXKAAZH9fhVh0u
EtaYYQzXphVHOHUXCkq6wYt01ijLAh0PTUaGgN7IwO4jPyFgfEWsqn/6GzHT
oW+BfCgRNTgSp9Y41W59tFb1jJy+BzAgTmbLJRdaOg7SHzfjO16KcIfcE+XT
FbdOKxlOxRy5DdGW6qHN1BaVq1mdF/5tB8R7OT/itcLOHwiHxPzqCEIkdPGp
3tOUPetZy5jQh829bwp4sOBj0/RgUmARCOHv06LWrFoc1KO0Iyc4JcRCpXR6
gqGHPIjFyOWoqKnGGPwE+n9/5uRVnrVPlj7LyZcMG7OE9yXuXBG47MCmON9i
3zAQJj5gkDNVCDy5WS2qzX8KJKzOOnfVQFfxj/mZSxVXFQFrs7YVrUvmCjXF
YPmJJXjk8FVBExyxdvf47rxL0yNkhLSyuYJDqOk9xNuOyaVxKMg+ZIDRY4tn
qkoLk/wTymShRoly7VlXsHLgKxHa2Gsob009QrlYzqXJsAXaQtrc28yJxocN
Kqp9iJZTBKw/N5MXOZ8eG0SUQzDDJuv9B0nVEHbxspUReK49qncxg6HfAdPf
O6a1wHgxck9cphrnDdOok1560Vx7T66IRNOUP76FxlFlzNCudnwI8z+kXSZe
uSLHLRQu4XateFa5x/DQ355cVpPrbwsLUE9koyiUce6azQB8kkCMRPyT/sTE
d15Tb5BPlBf3RZUa8+BJFp/9g7tLb5NHJ0tCHFrjPqMDodTR4aGwb1AeVm4Z
ll6IygbIMUXavfFSFJNQyNrqRz8J5JkJEUcGZa0Nyqcyuja8ebNr1OhcruV9
h32GEtsTZ/qcEyki4heaGBeHGKkmkZOy/l204OEA7T1rKI+IdBck/6Sc+MOJ
AfUnn/jhUl5Z1E6w+vT8lblLbgSbm+zuVbS8SRqqYK6EPAYYZVptNVGc1zvB
AcGEfKnk/J6bpyQ3DCEH8GNyjv/lpNkLk6ye+SqqWVxuy6LCI/Xo4GCcIJ9u
py/rOz4ZTxIwcL1DZ5RKPi9ZFgwDWiu8wYok/PMkBAtOg9G8gTBjChrTVGxU
VdTPnQF/4Zb1xnNhVz7wcrKYnFpTclRh3jQh4s6J/kPgwfQFeNC1GUoW30LJ
ocQQHxYMm7HI7EUjuWBL9tmFbwUFVueXPnRAoMLcToE+HtRtBWOB0BK0R8PE
6JPKAUyfjO491ths2ws2tzsySftkBuR8ruVR5Z1lj9Y6joXEDtmh80t+ALDF
XhRtMJBEYrSv3uYp1XHRpCm9PQKqPPDAzGSFdkIqGHsDyJVL+AQ0IEhDQlpQ
OdDoN9PuiE8Jcjzpu3EDZH9tmJijy3z+GFgZELOb0KDKqlmH/5XFvgA+Sc4r
48DGEaWmWv9dnntiV6kIMc2MSooLKYjn82Wp49chyuzvkGCxdScDLWcwFe7p
KATZKryEPjNtusz9TnA68jJsG/36i8o4pb0T5wK+FDcanoQIPtgexL5U8zy8
keIvVF+NBx7JomJoqDgqsjLqcDQM+XUr7cr7clNrSyUC1BcgvYCNpNJhwutW
nzMvvQJyE5ZHELfAXImi4FARa0XGjco/SKWSIiePaiRn78oqhokeZEKOnhNU
HiEqRmUAB02j1rNfcwQsX2F69MChRVGtKLhhKX8oKvOW/zXzqNBEnmBOZeSz
nXk84d637Z0YuXJtyjJDB+vZVBOF7Wu/77TojO6FqseSTcZ/MswQC2c/0bur
jsbItqjGQ0yEZFYjIv8yQZzCf7T90xVt9GI/2AU4aEUORzbgz4OvoJacWclM
wZJ0Wi0ZzIeKVrfi8H7xGN1JQXwymd0QAmkviFXjQr1uZjiKOQDVyE8X8bu2
ZHlDfG+L7G4XZPRpI8cQSCazOWobmOlM7vNA2rGtA1XxgfzzNUZPEXFPRX15
LAOOCPiuBuTD8xE+fCe3hJ2kbF2q0+t0m9ayvzMErPwpwhO/fltty9pggvJ0
yoyN+vX0tGBtaiTUYo5Ei1ib+Tv5rPfBTejl7fWkp/qeHJb8tpZiuFqer0FT
AwI+m8xPZ7TwGlsqLED+v/AK304XRh7SWD7tS26AglBqEPdR5MrmzF/8yHyo
StKEna0lkv0go8eePdw/qOUw2jUhasHjsuuHhkqkO2vRK8z4A/k1U2hQoXW0
8etoYCpwjNJa+3DnbI+wlxwxRNWMzpgUml/5x7ufsGQV6xTU5GaVPBWxMBFi
Ap/npSc3sRxMfupKOM9Hwuue36c1c2d4c1q4Yr5LUKY7VVWwXl/RRgzAIKOl
y2bUGrruKtr1bkxEvbj3Gbhn1WSLs1nVbegK5HqHozwzYLPgE/0KJZFJN4mK
3jX8hpWI9Wd8LkzqQVXyqYFqRw2w+1gy2nRrsLf0oNSjUB0Rd4O+JbUVWf8m
FoLxAplgAfA5w89NqX9p9lFbBOkjXjUOwRwWsUZg6e/8gJmR9P4+r3UY270Y
2Wfa5MEfSMCmQ0H4bT2CGcsLKU4JCGuTt5ykuUvIM0Ysamne3ICBYZMK3VJw
67t66ef+ndqT7/buwVvq+IpAmHknI9IyPpFfH95PBMQZTS1TOxEZxXEuDe7l
7qTmBAOpuOwf86VSKk2N8L6xSlV45aHLUx+XfEWp4zC0Mr/4zVB5Kk0RPgiZ
jvYRAaRjrRtETH1IcSpU1U6r9dVZI0mwWiyv8aQlOhN81Cvgpb97iGlhdBqU
iAdazkNcowcKzomGMkZqn8/QaDTOAN0XA2AhQRe0suz2EP7leSpnACYKlsyp
+Tp1qPSlfAfOWwkln5VdtC0Il0dtdXGwjzQQg4Akso5bDkGA6ImMnRwaCr/p
6hkleFB5jVJWm7+TOaturkFepb9lDhCkFetAjaC1pyqAdF+7bifq8xcS70GT
fjxF1GvE5bW1A5RHE1q7wT2uQZNI0H/nKG7PNOv3y2YdKQgQ3siPz3COrPaN
4x8lI/IbdPcrNCjtFffH9GXtCc3TWGN2aIPZGe1QVBpGJNW1estWedn468QN
4Bw/asmie3up77uBffknNVXcKX0ETC0RbYxGN+OBvDYYPqvHxi4UTiv7N1vh
wOCzklUvSdfJcSiN8Xa2LqYKwMefEraV8t1AcuW/UUqykw5cRcbX1C95cni6
rKjrdGrxmWvNrtSGZ3kGmyxFXSC9/YKde9d9NeLVvupmPBZA4wx8NmXhTpwD
HihwQus+yVOGBwrnDwmswppfThxKypuWCl/DQbK2bkpIMNP8jTeS5RyNhLbr
K4tbly3RRNi1GiwWFK4R5P9yCHOu7jRQPGlLsb5kkpDaH9kae8J4YcEhV2D5
Q4z5ivvFOW8vtqQk5QiB+1B6WKsQaKcreDTmD0zoMSQuRbAME7Dlz9s1Mp4+
HGUxSawG+z7zh80JzZnonaFkztxcrc5e2M1U+ABmiJGPqSXdY62Ans4Tk6RI
MHkZ8tJvgsfuULgx0gNwB/fgModWYqcul/t8/XiqDz2pFXZu4CTCIg1EAe9A
+v0nWE0Bnl6BiBQQ2xdj4ze0B0QKNRxAdc3rGiis0pZYIK0jQHCnogRXw0nx
wwCWrJXSZevg+z19jGQ8irSK7amBvqZHOVKSjlbomWz19ufyY0XjG6PKYr2h
++JrWE8wcJQs2BQp2mMcneKJIFVTrIcG34Gt9K5kh+MaxES2M1UmXPsGusw6
z/XFuzOI3DJu50O+iXAXfd+Nqhae2SevMReKtsBRPuVf/Cn+YoL+9QP4OoBb
zzwq0BEW+V7IpIeJ43gCKZxE7+XkK5VeZT4EVeVFxOPwIu4CHXfDw4TU7B8h
LnkkU3g5tCfaImOMLL1aDEAyl8BQaVwKD2uDI7+HnNj0OrFschNDRJ2thpOI
eW8zAgQxY0KhJmr2Y0gYt9naEEm3J8LEXJEBCr9nVDLRi0BPaGFp452GBl3b
DqerSj78BaoDjyYUpaGwKFs0K8Qqg4Gfy8TLqFqCzFyvvoa+byK0gY04z+gV
hYW1dpsC0OAuqKAsQoCc6KFBpmziVSVZQTk/gJ8HWD/CpU2+RHBR7bde8c5Z
xOuKmx29QnlSDRe07kyPa1/Xjul0tcQaukJw9fTRNrc//av5VagijkUNUXps
994dY4MXdKoyijEV4zHmah+u7Pd2kqAr05Ep9rVXmg0/WlMuQyGGFFr5iXOo
E/7C654EY+zsLm4A7irTI1nuRKkGZ1eDZkTra8d2jnzO+4ZeOjAcGrazr9bx
WAq/kATS8b55AXns4eDEl3kzC1lIAF1/C7K7jlFiM5kbNB1S7L7jaBkryPnD
CQrplSe9zwLSnVaovWo6acmAiA3dkLVizSNSScZthrnyUHepW1b/1UhjJV2P
klAaMDWvSf14Bs+phudfxbhKN1Y7cSNdD10DYluzY+H7hgyz6YSXxVln0ZW7
K1rc9J5LnHOKln4+FbYbyhYAMmGy0jrIY1satpADV/AHpNyVrVVSQg0VesSf
+GOXv0TvR8bEz/WmY0ZTZhFqlprJMdrBcobJUTjA2NuTR9mzrDBlzQu0AW9P
RD9kfXb89YEj+GhadHtVJy7oTRde7GgTDNTip51hW46dxaUiixQv5f2TfAYN
E/6eQORMQIfOBg0M05Joax/NrtiAKAfGlqxM8ktRU57XCAMVp6PDzcslmqAC
7jwVnNRVzafqNUvaVcotS3fqggy/6+rCMJp0sBF9WEBhbLKVF+e0c+6MTcwk
W+98riWgPqPzb/TayBZg1HEy1Kh6wR0CTZA/usDirh3jlFS0jEuJrCs6HgKv
pEYSs5WoBqQjfhMszm8StqFBZH8KFdh5Sl5nttiKOPwHQZWHSnTGxUVn0V48
oMnJh8RMI8aTZZu6//H/4JAbphH+bXSBUV7GvC035xqQeMMMCy3SCuwd71TG
AsTRYVnQITxVQiVK4FJ1IojhNxXMcv1GO+iVmEhaM5GZFeby/tU1ugojQF5B
vdNFcAter8yqHaPdVCpNQ1Fkh7xibD/TF187e+Wr+UZEeADVoHjqQsRtIPk4
kxqWkL/6PHAHpgcIkcgAfjtNcxN2E5FtBFP+5UIsNU9fuKYg1MoVSuOYNrLn
277xYMJitWbzX2z7os/WqfVcO/14mYhuCgVa6azIYv6w2VugOf4HTJ3AXJWE
aw1+SjXWP/TDMFnLJeXc5/aliwD5JZXwBPYewLqL7Tbcs5f/O1kB1ufOvh3s
tjtWBKvzujzU4K/+iSdqXYA27jcNuG1sRdfe8a0rufEtcBbUHMKVGygG0xe0
AHbWV6CXuT1GTaR0NNPk29LM4e39G/bh4lGfJhgDNhvmDKcksEQXg4+PMDpB
TbSJF5PuDqj+EMdrDrd+YqdUkw848HvkPZInz4ja9lWQESsfKt2k4HrTiT80
S2ej88OyS4g2xef44FjERqdf1CWAROrv4I4T3fw5HIaGngRkunxlD7yJCuj/
98rJKGOang473/TehPLg4CUFO6Y4aouGXpttMBneJdWlm0IE5dlZ1XsYHmgZ
RKBzStl9Iuehju5oM6dGYRTfcrztHrpQg56TE7UkNVJ0OE4WX8xixFCxuCvt
nALdokQQji5fBqkj2MODERR2doXmqSZDXZiq3ybr1DEX9SPkUQOejAqK3FjN
87sHc6HOovO7T5ZVC9TDsAUfexGFUUSPYLPBfEyQm5Xl8Ew9/5lk6SI3vE7T
zh1i/JVD6biPu0WXpQAfogou6O6p2BZ4antvONGlMJWsoRjFSVuBzowokh6I
MTILDtoFO0dFqiQFuDywL+/GFckU31WDOdVacYWavzTN58x5IZwxaejstKLD
e+e6pK027nArCOOTgb1+UeJRkqXYv0xcJ/ZSTVGWAvvP6ckf6TIqfqDlwNPi
VJnIj6UM+Es64GIW2dE/PJdyjGTgWYE2O3eBpO13SvKoc1Cu9bXr64IA6ifw
iyASIVaabp2xQvQKzzfmNps2v9DJdh2n3asBgwj5dmLdYm9U8fRAWZAq5qzE
p34hB5V+xDQcKg0YIKYyQ7yDJ48JrwyLc5YIHS/++074m/maI0vKjoJ0ISps
6ozrb3208/nlYFRTYAflJDYkRyjK4pwM1mAS3hGg3MJPbkLZT6Ro9cBIYT3e
heSzbRRAF59Kh3ZUsdA1xhxdQYqA25vYdoXMa5xHP8sQufnMo3YgxXtMDrqK
gpZ8HXeixaBsbpDmwfL47MmVhygQKtH8Rh4tyceekXRmukr/dnVvNjSku+7W
K405vNW5Y9No2dTbd7U5LFPs6gPUyvl17bJCpeqU/2kBs/jMw2xWIaH6kV7n
lvQICzL7f/NggjqBDorVl52xE1k708TyS2a8CJxOYGl/fWpB1TBpZVD4LA8k
RGx7x2SPSMz11K++I2ImyZ7SmoQ6XDFKuyV9TO1nviSONdrZuvJJVOcO059y
APoP+O+BpGO6XsSumYenwmTh9Jyebh325P5sAumNfPuKJV2p56xR8c4K+9j8
njZL0nQGzCl4KRCqBLK8Q+giJlmcqGDumkpDnJbqZb7Qe5mUnC7qj53hpO/L
tQsDimrY1CE9X5zLtky9iOuxCo0sxrkPT9j5NZVkW0CZXRUilyeHEBoxGLyo
T5P0DGeHOxivM8wc5vcu/FkOYAWVBniTbRNVCzzEDM345NTon32qHsFwwdou
RTkmfeCsF2h6o+dlhZqaXcLoRoQ/CDd7Ae58/I2QazB7kKXf0e2tvw/M4Jsn
6kqCES58LRLbRsxgyOnWgQ+WGoJAyVICxNY7lh/jY8gC4vQt5ZgcPTbgUjcN
zXCad4KEF9azNQdGM/VGbcLC4kbU0jaYfUtsSh7syJEoujoV1mHd/v+uKX+J
xysYC0YPPys8AmKFL0fhpGSlDrCKzApg42gtHqopJz71iSZM8xOZV/LUmR1z
2vWIom1Jq6tJbcQ9eXfQIoVIQw0TIk8KCgdS1rx4XlrsGaQpNawsBosM6azg
LpCiPSciAx5n447SaLWXx2uXfCBD1/WqNt1eicaQgxv9xghVghiDnvhTN5iM
i3QyM/O2yR+NRmd/m2br/+wWFlnv8CJyNE1AStlHMO7avr38d2VdyvOUV86Z
IGKhpnNQsF4xz+6WMUSQMgg9F5j1IcRimCIjIi5SaeVUTCsLapa5hYcJevav
6mRBdq6VI2p5T7n9+Fm5zgnQx1ayNmqa3kuycmQmAUAWJXY/RVegNUySP+Z/
DU+1ZJin6AzKyQQ8R0LHIZjfZHjn2DRvhBPqwovECCQbiVryKS5rF96IGliW
hHQOgby4z1KaYZJF4JimEEeb6suNzyiu2Ivx8Ne4IlSyXvyf9jHVB9XL8NG8
nwT3Ln/xwK0ITfXLGp2SRneFMDuy4WZduHw7CvLRbCHK4wT8l+MKfmOKue49
Z3WnvAez8Q8ROZ542LzqFDzmFyUujTJKH+9WaFJaTmbwy+tvAX6d3VztaHra
BTu3SBO1rG02zkwnvUs371oU6a+C9vUYJsok3CNqzv9LOI7awCs9mBgJ/lzK
yiZT3B9IPeYFVUV1PVUQZy28Co0uLALcMPW1QzMGVgx5YQKNqU3yi/5F/06Z
rRhNWHrrV0wYVIkVtEpMQq13IV3gkvGjCoI6yy4kWpqh+kB0AT2dCkk50NB8
tV10SPwXK7q3cBmd2LKep6rh5luk+dGptiGHhmjNqQH8OOqM6ot9X8y+++Cu
psQLCcyBRtijkj5LRx0W1tN2t9WeuebZL1T3BjZPZOsLsf2AE7r2btyCv2WR
Uj1XBeoWw39KUNjmkGNgX8hFKz6p8nB1hLWiAeWSWOnW7jfNmnJmOI3P/4/3
f4nakWj41taaP0Gf54/1if7+G2mbC1HD8HK9cdYBty+8Yj1bqWcCgB+mOqN1
N6onj1TiKzDLr2qsf0eMvZuPYz1TgNDMKBU1OUf70KU/PIk3H3nJBhFJyu7S
puql+sk2ATJORnehy1XzLWLdiRfRNa2Goh5uJdQ0ubfdVk3s7ZpekcwIMb2w
6SuYRw0ERSFyM32/WXnMNNCcaTZ+GmqoogLtb34m6qSPafECSIoaaqImtX5F
/OnjxTRFyZol0IfAnPGCQaNBIaOUsSFkfjYPck1wadpKXoKy1Z82gHa4XBDO
+zaWbQbpVDWh20epBPiBp1lCl7ljw2jTsPre0rjdrDYgqG/c46jTvcKmrjVp
Pt204fgTDRRaAmaqoPwHSt1x/QqJVt1QpztcVNE0vICui6mMwKkKNYUJR/HC
hDxdpkTUZNWyO4ZMNsQQBb6uh0e+8dAZqQErKLvhJbvBceTxNbJrc33W+E3O
HM+cFZHOW2erJg+sd/+5b6CL0P+SMnq3yJ7YfEPLq25TezdSI8hTb7EMyyo+
4lRf3vUlv5K0hn6GVe1kQVq8fnI7rACcVqfdqOrmAZttRP6i50RKYi0267yh
YzDTwkBHkUCAgEZABlW9zbBVwcGRi1E9f6nba9vuAz9eylTO06cZ9ZTwZhJT
Gb6lwikxyG4AeuYwoFp4yHKrsShmvvavrRs6Xm8I5Omam1+OYwpurYoazD/K
3CW5AcKSxOqTK0FF1pjp4VEZ446CH2Qc/+lhF0G9rIBIo3EkTbg2v4IC9tgF
p5JFGtBf5B+8bZ3K1x6w7N+HVdYsgfvka0jYg7JeMCQ3QOMbOIbkIPhQajbk
w2wgbb8dOvcp3ttpOn5X2Xidl7l79RtVLgn7/E1Im3e0Q8C+rF1RGIHpSptn
+1vFQt1duH2bAM9ZADYk88jVYaFHBP3748jUASmWksCS2sK+33qnRDLJZuIo
6f8wZ8GsAz/1rpcidSwXfbKQoV1UAreKZ6mAisxEg9yTEDpmd6RomJefkurA
FuqsQeFjOdfqg1zhkDJdiacKybA/SLINqbHFT15VudVAcVfVq2d5m1bSQRm0
ADFcEHmbnoOqwJS+Q3/6P+1geeQP/3TFAD+vr8BVqkqxXKh6Uw7BJSLqx3G9
XhCLgIYuX/JWVo4/7ZF4OqeTKMs1l9qIcWJfEO5E9r3csP7vAYEErWb4mN+R
6ej8aZxur5ADMcSPzQJixTYOmq2vRbO5FOdw3eAgM1dvkhoC/dGJmpZR5PwI
mMiseKQxj6ebmXydVAkjGRCo6dLrny4CTd6S1d05B9SHra5347zUpYD/4GnA
et4gLg4fkUYi5lygZFxrSBtTGidPZw+i0Msdi7bUvc/+jLE7eIxlizUgE06h
v9lj8bdiYBP3jFbH8WCEe8OAhqX4kqooAHNBYLtrqts+XwxGFtiEkjqlCrb7
DADzllmlBseHxFogS2BZSYkBOrGiS6RE172NVxs1eCAT8O3wjRg/Js5Mz4Xt
T8iVMtY24uB2BsLxawulKNPytz792t2kQxMtN1RqtN7PPLQVpE7QJQL3Kw0d
e1zcu7vGLxJvhcnbZubc5AiQg8GC11N3q9dLgYagypTExKFZPBAJq/VYGR9D
hXrkMNd/um3yYkQbLr/SCtc8hfXR0Kh6ZgfIxCxR5Kh/1Ds6ofvAQgCStiN2
5fH9yIJ/6uD6H+K6ZE04WSJvB6n/SugTVkRzIUkXBjNq0N/fmgsO7i4z2fJs
TlrhRlVkm73sNlQ6oXb0CfV45RXhhNi/1j7QBHyQDkjn7dCKYv5EJzFbLlcI
aNjrjhI304JyEGjKh+CPvutLwBg3gI7rIplprX1VgRXm16l+ShCbHf/2QFzZ
AdGIyCG7qmni2C7+RpwMLHyarHI03TPJFS7bC9QuXX8pbkk5ktNpZ/zbWAZj
QUEdp3dFVBah2u8pZPRlKnQpMeJzNUvAtix1+iM7e8IbwOtyXx5hKxJwlhbP
SIHPPgufWsoxWIj84CtzAS7Dfr2vUtlQNFpm7k/x5heEIcB5cz9lSsvbK75B
o+I832gs50KZTi5tHrvCOL8bvzSjTI9mfb7cLCeBIavrbCAHnizbzJOnLM2Q
dSjx+/Za+YTtdk9fdltFQRD+70v/wcHmNgBfD9DerErTnMn//TncHhdcADw8
rhe18XjYr83nBAkaxzMUNeuD/6wEhf2pxsG9Yl/WaC7P9NI+9IHt5P41XbDG
rnX7oAf819t0KQtm3jtIEu2PhWd28cvPqP79E0kr5wDCHG/k/sbuBulaNrZv
xjiv089Bsz4u6zvHP7wy1rAi8byWmzSFfwq2DGck22bUkgKxYgssD7to2yvb
cUlUrhXL0Ta3ie4vpT31BhKIm7M+B9u9hth71SyuHpPpuQE+y4hfTuJagYOJ
EakZ7xm3P12b2+bpnEnr09GMiZRex5z6he1TCMudN9zgXmTX44DmPPAfJI2b
nvKusy3EATHAMNAjuJf8gVuagWjnGITsIfpVNtxHOZx9OeOGWWl3/+5X0Txd
G48rCAYlsufX36KdRswXTAXWz1Rs3wD/wIbg5TImc4nyZZZBtlquVhgIuSof
ctVfp3scdc7o8uOPOldk6QsoMsUdEuSCII+X/icDBrXt2WuOIEduEvReMMje
fibrj6Uum2kTaqwug2Ej9QiOdDJkHSVuHoGKmGMIZ3hnJkUoDsYl53QTAkNg
9Gv4g90LavKmSEzHGC52ImMu7WJqDnoSMQM6+mdJzB1H/7Vvzy50VoCHrRki
8B+L+b5C9ryxZ9AEc3rvOLhEou6ViH4E4FUWjgxQWT7NiuivDQ7JIZeKT2ro
oasiYSVLPIgJ9T+uv42CCtuvI6wmMQSU0+Qsx0Iu6ycKT1OH6u4+4XVcg0Gw
c2XDYqd2FnpphV7h66r/pMue+0rJFHRbSdwqtAFpu3wjbfTr8SUOnht2rbmN
oPNys22ZFosFkcWOvWmfAeu02TO9bU0QULhY/5ZuRaHQRZe/Epjmt1Bg0C/j
j6CGjfLuTU7TO59W6bMHnPBDPdedaoHsWgGep7ZCKou/uT/4j6tC9mi8Jb+k
gJq52ykpE0o+WRx5B/4XW0885ryUlMuWmctr7hsIRpTSygNAUEqSO4d9UkBb
/SWsoTPypYufQqC9eX2DO3juFw47s6pz438AP9ORHOiLMGy/O8RbVs0Vqod2
fXQBxJFEGqmRGJEJ8V1sMx7z3jHnY7mlbYsh5k1KR01EuIcFkq0JyxNxxHuo
I0MDOELPoTHmyJEM0Zuxm++I+vTufodErsiObzTvBeFk+ezUvWr5glxhFo6X
iY1htw/Sf0bHYbnW71NmnJDJ++oBXTKzBUvUH/tzKFRG0eRMafQsTZIa84gR
tkcUrQ1FYIV/dMJVof//GTpySph3I0IEc1kV22DCqAwKfqLTsOj14BIH6zPx
1QP/Zrr+BebndpRUqa1xMjWBSmUnJu5wCJB9eVbE+OaiHgYcF9tbrBT6aFJz
o/kCS1I8JpUIblHFs4vNpCazT1vUpaZOjwWaNXHUX+G9u2zV0sH00KUwP9UV
h2ObYasVzp/kxhm9zuI74ECVjOUjBfbXYLrukYhSguEG4tPY2VzbML994xT9
ywaS5poLA59VKjpj6hARSvrFDr5l8j4bqOgPzDw5qrG4VWPtN8qnblU111nV
uUghofSkK/6TMUTcCrMr6nCUJ8jzCVAAsXGMtDz7Y213bOtorsEsi5Anm7Sm
C00YEuzB8Y3AsLO/lMelKAupmlT5VShlsulp6+2L4yfQAM6cVtwLuo6607G0
2sGf32begRFqqhLTRaaY+qWczodFJzeuYGYPogBhLyG1kmim5bXKGYm+B6X9
Cyi8JviQgMCo1Wy/2jZMznbID0vn1vSf1f0TcoTOwOuxGeWwsjdTGiXe2AA9
6EpSd7q++I2waeqRKUk+OwjDgWQXBZInsg/Ep8v4hG8xiIhmaIanfDC1XcTi
DmCE0hcP31KUComKdk3sZnWkwJHyZ51XtX8A6/CLqxTRC7rcMd1xB5lg59E0
5lQMJa0BMZS+3reFm82t6/6GOe+RU44ekJT+qtTc9q9qaX/ezQwG1yvE4bAq
m4r+oCkPQqBkB63XB6QVieoyzjHYx+EbUcMuPaClCJNYxw9zfSmmivURfNMY
aVdudLivXMyTTDU7lNdWd/OR1Ay21zOI1DtJxryLb5NWVeqEKg0Ax45Z5Aj2
RPVpEcYz+N6wXWjdpszlPkjGf8t6byscvXzSBlYx/w4DWh5nfdRXDDVYB4kp
5e/GAuJMqsPWQxadnKdgOa5c8DSikp40vv1qH7QWnH3ZVn4/TE6sW+sHlf2p
No2Z4FH/ivD3bZS9U5rwLPWzSIypI/tf2mGA8GUDzshnDkw1/c8Z3E6M82C/
kML9E7GTeeAvaYHQ0kYrFF3BJF5vPLeMvckpJ8gQzuCt7vKfA9YMaIe4TYYH
BvBFbdgRW2Ws4OPh3Sbsy3oELJmg09C53WuutC+lC/LOG+p29BDNXbgiZyxX
2M6AtsetOGF1+xRM9t42tsVoDCe850nDj+/I+a1l7E+PiUAhZduOdR8JUvGd
Axw9g5oi/Niy6Q6xtRpsO8eAAF4RNVZuSoV95W90KngHaeu9TW9nutJOXtEK
i9KNyn6gwBsI7tkO4OA+zB0KbdRqSdokcKiDSa8QUQIHOHAyWVSe2znsmiHg
7FbPZLnF24YI4AOyOsQjfyth7cVx0QajUmCVQRbUzcKjyCQI574FJDTLHSUJ
Y9eCQAJ+yzJ1WK4wbyAvE/gz21txrGolqxuMwH4f3jfLwV4OQ8pB7akWgX/K
DeNhOMn/OIrmOzNo6R+SwHn+ywkwIJOBqTduLjGcqMJYxxpgYPpeQHQX0llO
b2eqM9R/ReHwReFk7fShSU6D4Yj0L7zwC1+7u4JtUtkfzbTrxYgflwLGvwdB
fHp+tp5nUnH0RZNdC8n3LdI6DxWrvCIBfJ3y9y+eSp8ezF+Xq7sE0nHZ0+eq
OolJVf7OK3giP0MRJaA+OiIhNnsTagKQJ2CedjRxE7Oy1ZL8//KipFcYuUkh
3yKvrakyQKDLcFbwwnqLD+P0UPrC78R9Jm8pwkUbunTphl6viQ7iJIs+xegw
rmia34ncyVIEGCizgOnTR28bqQxvXyvH/1Fo+1adswmfu8c5PBXJK/ZsjpAs
4brovL/VbfjsEG2mXep2Jn30WUkx8ayn+Omx38yyjUMUyzSFlsO/Eif2IsWN
UF0EBb0L7qBiCJFwuZn2eoCwNnSzVwnJz9G/xeZeeZtxG0PhXI9jdXedYjG/
sZ+190TCbnYUOtb2Nci5AXGMwQ864r5+3reQsfl0aivhUQJwVUKIu7xTQUAd
9TYp9bmmJxMCS9h+3FePJlCIrTTJV+zE2d7bsK+bF+CmF292cCdeyZHvBTz2
TijbXhhQM3UdCqSBC3tcO7wUjsv4oNhx7zKmjkwnpAoHYoJRGBtjuuvjkriz
AOnfa9jjN36OJV/3oAVhe5QGamAk8K8QbNKyqEC1OEGiM3o6MuXk9RHWcWl0
SeGNbzQKDyil6zJ9NNZXn3al7KwRHZy2i7DWLGUfmpZ/03vXuDFbxBK7oq1h
SWPsukE7NUtXnyfCw5h1drJnHUMWofOW4BD1QBPQQ5GjcU9JIohrtvFy/ANq
RlSGIOADKcnXtnYoXhHmkgIRc95qKj3av+8Db6Qj1wxeSLoMzZnIVa7Fuxx7
7wRg4c+tgC0ToPsRqc/v0NT7+jqGbbQXzWVQJ5veTkFIITt8rH0NYofLPkB6
K5ZRi5yhobX1Wrnbint7WIB5F9e//uuDP6Z/OTWj4D6MLmIhadL6Hw6fp+xh
vdYSKMnGKeMHdVvYN/Q5Sq9cd+X8puqd8ccoaANbAfqTX71+FADaqlSWaPJB
scePw5B+K9ikyHqVXQny7baavbWS1BG0paXtDH/5j8ROFjfE5GNN8X9Ky2AZ
dFh9QYg58zSwMlTGzGno/aNUnEQaeSAc+XdgJEBtcIBSr7BmMxsV5SwCEcIj
H/YpDEbfx3xS9PCV0ZJJ7ruCfh440Ntncepin0pwKRdx0n42DtEmZTnBHPvG
EaT64xtbGmiXlRP7f5WVXC8lWr+koWEloAIljEKHEee77ybnwlvwlE4yDjgt
1ukxZQFBu/nut7EbK03QQa3TzmVHts1NUoCG7uAupXglc8UjGbVyESjbE4mK
emiRLpcBl8Es3nUWGw4mEMMmri2RI/ZGkznzN/CCPUTmWaqGRESVa6LBO671
R8HN5E5mwWttb+EhSYqiqxCpsubrlTV3VloB274sCxhWdRi6uRNlcEcOyU/8
WW4SG3AONhF0AHQd9wgc8D0tXtZl6zuDasRIM43wLpgkvOx8mNo7kAef9njb
H4oFsfuoJ7eNqZTk92IrIn767WyTItaZ3MJeFkrDNSUfhqK08NaXuSLu8G8L
1iN18CLkamdEgeH6BQ21kkXT5AUm1rIQYsDSGwD/cPJHvs6OXYBUrr+voKt6
kk6upMBu0qAqX8TM0UgCaTOxpEakp8axLPi6GuGwi1YJEHcbaQ1DLmUY2W8d
sAQoOcrGg/nrxSQnJFtITB8o+Ay1L9iaj5LV+Cx2R8mV8OypWQeStjXVIx+/
Z1Ia2xP5MCrqynqyPrvftFgHDR4A39er3g43jEFz9uAqOVkMJtGfOtMGqLPE
7D/FajN1eZS4E0VwI4ZUY7qJX1S2ZVayB09vlrnvHwMjdTNsWthHVVDiT1NX
KoI0n2DMsnqWuHzJWm6svw5YkdSQi5uHu8FLXeRs5PNhRT8ylqR/+K697Btz
Plenf1TFh400LYC6W5+V35REUAhbeNBrtIpM3PwcFcbb029HgQea8huyad1n
rcEdcsfiR+FNAklSh0GRi9vOk/+lXl0vfG+PozG3rDAUD8Dmn+Kad3gYSHEN
UXux7JnIxAaGxt1cMyk5ymDhEDzMmJSSA05OzC3zU38J55UM+YYCDcHprn2H
n0+uSGoxsaftMvrtSQHky+V9Yc+jy8haEzC0EXO82pFMyoBvRBJutvQVCZ9C
oUch8NbVousBhX69lmr4MmU52YCGSIOhavud/m2X33CY0Cn1xBnZPMUaOuDt
/ucmf+r9N4XRXGfRQT/m2DtSPhcukPCLGbJrrtETZJC8VoEHdQnqzAOOEeZ7
TUVpQGZVSqGD4xOtWrlLyjVphNwP16ZmUz1iM/e5J+cDSQx4Q5gCQbyEL031
otZTBmN4wEecMUHbKuVbZSRK+OWfIb/OOcboRtFL1FQD+EnS2x/u98ZDljgN
dne3PRCOIld7g6IHAlTfIKW0fTmIteePhvQIyNMgKAlKCtx+7jcwD4/2bojC
OVTyQiWY8pLYviZ/jUFPdjSbcQSDmtqgvaDo3W4K5toY8tAlPNmEbF4/vG+e
KUin0xGMShWNJL/micfPAN6ni5EhF7VA7ofpsq1qh+66BaDwoMhpoGfTooEW
9HfSYk+8z2vuynMVqsS9uveV7OwxAqP/78Qie8WvAoF+JmaxDUS7whtsJmaH
YWXkZVIAN3aKtsDWXF+zbVFArAkiZsYOWyF445efh5PQxse8b1phGZj9IrQT
fb6DpQWO4JKuGo7zKGBFT2f59KFElW2oRqm2/VLf3H7oIIFsxCpbFcHg2qvL
EKJ8/exZuYU3Vt5251JJEZ37IXkKtlchItpYM6tO3q9DMT3HuXloQHzwktsy
rmIVGz/1OE1mCKY5dWeTpUM0p4EADq03TY3ZS3zGj2hWBXJI7puAi9dKGAbV
Sao2ni2+0lJzYpTwua8XXl1AYwaAFUAR29VvpfhitTLso5eI1w7DrAakWlLJ
zBEPg8j7DPmrANFgHYxHliV0kFoxxouj/61tym2n/O0qjiW55776MjFLlZB/
P9VFIRpK2FFlu1bdIV8Jp33UQnDUls0dB+uZtWKgpPscZlFgR2ZnopZL3SUK
D3RbxQggmw+rZmhfssREHtN5YaUl27NEMyjkequSHjoJjPR34NiNM44czr7j
QbN2cK1RpvWsCGBDhjGA6446g0BnFQLLaehhhIUnKFa5vgEYQbcOgyLFP36G
IjMyX0Hy9WMTmpwmcOsO4hEsFqse8ijUsR8CeU/ogWxQK5t0cOvtPRChhmiw
vqlc0S8RKFzECfCycqIYG1rqzQBJQtv0RHxrieJy4lHRNWwtDd5rzUN1bCbL
r4ObdN5xU6qGd+beONKGaM5rM7TE/PPb7WIl5AzpbxdzUJM9SCcV1jaLe1Rr
33R3vqdCkx4uFvQiF92VgfVjESeLCqaNnDQM3XjdSYBpfM01ybOekGvGoo2z
+12A/ePqmVdVKCxPKi25STjuen6SFHEQdcp4FmiSGJCLGztTqjDwP6C1Visw
15FXeVXbB3+KksNXBYR4LklPXuZtvU5xHbJQbtlSU2Vyf7FmGkCg/vBzaBhW
BHUqn223fO6m9DbGlyGm7wuLxUxjUxAhx0Bdg2RhbvyiWMi7uuKVIxRvtLy7
NbqgDZR9dSMqRf12ugEfDrnAEH9aDqifDb2bpGHgVilht0lImjEAWcGHSZzp
7KyikyqsYqU9TXSoIyzUJqvJ3wLz6t8KvGjSuVnBPfVDOPtQnXlUvFqePEJ2
hEBhBrHQc7sVCILvDD/xoSsVfT1jzXUijKOa2+nb3GKcCsQ0RdNn9qSN3lrD
3ICv8ImCLx7R/ynnv6Z1VWlnVjpI0gEfvtcR5EjTP4v160LFX92YbUS2HXEI
SJP+dr3pbvTRL2fClPsuDZ/ZM1vIkXkTf9m9EcG7AEJz2uBI7+P8ESGxEceC
sqLTpUxpib7RQeox0Vl+xlRnU7v7hDKAE7Z/cqpH8HatoEDJHbBbvLNAXtfQ
sTSpqARu0qL4zkwsDCiB/0T0JRNnd+uZJFevA5LOpjy8uujf/kKIkrf6I+f3
g1D1rA8ayMRoM4DHweiHHVtJN8TEfQos41p7OVPUAaKzx79kS+XYA8xpzQGO
8hBWsAxNZaneEII/OThWskPsfIwUJ54aUXxJbA+uBK3SAmjZ5DzFrft/VRlt
oyM4/IPRAhqqFY5/7lzPkZ9+fLgOyCPSyuEzhypt7cO/I5mto/IhGGm8i9l6
WAuLudr21NXFINfJyGXxmNUuY/4PoiHgh8Qqbtl/OAwcz+/lgGcP5G9lUJac
VjbL7hc/cT25P59xzR/QD0YJsZov7aBR7kkDTGkHKK9gm70xNYY+nEQUguNH
+TJ73UW/ZhwufiCxEtxDdSjrBg+jqejmCgt8qU7N1Il+noRpUbnufWBNPveN
xizNmZF2S5G6CHcSY/ig+rpySHTckF06sEegAXkv1QlLbCzwWoeudOSaMuIo
JZAiNlEK2j2UuO68rEOzzvOpk6BLUpvYdIFWQzbX2trA2TqT1IE8KkLdgdQp
YRGIoCu4NTabUtbDCHBwFIpHMvRJdr6rbBODoM1Y5DYP2vYdesD7Y32vO8Bb
FaT/I2i2PnVG9nL30rKl3Ym31CyXe7T2Q4OagCFj0iif1klfYND8L6Kor8Oc
/9fU3n3mXwIJt9yaLS32Uu0Is+sTspGFjIOC0/DlZExiSJPhnM+UdGi+ZaPO
fzM3mYOnpPMB7/m2lyxQpOhTAllpjauz+8cJLr5VQy1HA7Su0ZV+UYSq48ut
nsc4rskt06dzeiO9SSIC3MHRmSUPZ9UrQL4vr8As8ZhwnuJcC9m0kphDMaWm
Pdya7XZ/5O+DOmSfPdPK1QgjJ0vBeQUNxsS4ew5tQ/elF8c928gnXGU9Ilxh
JFFubH8TpEmfNS07GqVCmTd4qH5fo5KkMqfDno83yz8clih+E4PwRYFP0LOA
XF3C8l6b39M2KmRyIGVPWn2Qa1EKlnLAx8wUGF5WHTA7gwoMEORB13W1NQun
fNJgCX4izXM0RtUocnxZq3eYvyTOzqRLd3uj5ZmxlpTS4Wke+m478Iw20Bm9
j6dCpdBRBLu+GxC31jq0gasN4Cj1EYKgoM6wdcIZHNLPboKVkfxN5zgsoRL8
U04MQYXgkM3g8tO+MoQQkt0rLrZ7NWbcJaRikrckxii5DPHSOtLTef/zRmGD
JxZbL3RB3MGDDmmBXKlzr8MOa5DSYIuPgI7KVWwmB+wc+M6up80ZE9lPfTEi
1Fa+MnfyzgMEM8+6EX2mcpWaldJy9oUNaHnax5SIYyaGULMFx6tsW4P+TzYH
k2PCsdboF7ffIVmBZ49xkEXnHK5oiFeHy7U5TtcU92mghaTQyxDadcBTNhYW
N3tJVrBhUfn5EmpP+M8HUzo/jYZFeTmQQurILYUEZkv0wsjorGI/6q6iT8dB
NIXQv+gp21DLFMLDHtT7v7rAiv+u4olGvGC229K6zSw2fGqG+UsFVPXvpND/
Hg1ELhl2sKmUpneD+mDOEHF2YQU1Mv14M8NP1k5b2llR79hfyNQgxBp7lj59
nM+HwnGkqA4lrbE8PZaBSu5lERExh3l/+Ul8bwwEOW1qsAroxPqjZ4DRrj6U
74+yyKGNBM9GvHvhobdPu0OMC1fJ0yiUwT8EWbnnNDdRIt4zESrZ6uTyIOCb
eKURMNzzm58KkNU2D560Qgc5/IMlNw8d35ZUY3HZC2qK4LmWbTFFuMFMoKMq
yVF2u8EMKWvU3wF6X7sdQvMnwwqCJwJAvy9ju1o6yweWnj4TdvsIg7PPPj24
cVLbUlPgwqxpAZx07Q8NYHVawgnGUkY3TsLZjNrfdjTeMy4yjhTU8YYW1T52
GA2aSL63UYxCT9aBz+Woj8qqZFBcHuFEU01JsGB6IBOO1Nea+bLdKD1a/HI0
RJusXuTCsi5DkLdnL0KNym9GyE3KrmbSeWHxRV9G7hWRrbVcWI69XT52d4A2
1TYWapDg7cv1SXopQ/fD7N0m9K+oJeTq/z4OtONb/GXDGvKAitcBKxoIo8Lf
jYpuZuJ3LpBHw/X0kHYFqsbsWCrmK/y6Uq+RwQS53i1X6sJVbRsEBHtAhslr
3Zo1kWhXCDJ+RG9Uqwq9/bvR68KP4favR7tijr3Vw9klRrmx4m9oOSmapC0F
ImsL7W2U53/fqwPrbZb1csWM6R94Cw2WP5yTWlxN/Gn979UNux+x4HEFBa6a
dFO1RFJrcjByUCMhe90ScLAKNlb1g/U7nEjfAwMSZAX2Mq0EHHgYtsz0ggKu
fkCqjdMgdmGMKboSIZZzgfBQZ8IFsMXFWe+bjCA1ElZ3rJb4qN4nHRt188c0
pjdtyYY32W+Xv7hpEJUMt6p/x5p0Ag9aPmtirihKzstOB72qFxQaSo3sKISP
0eAgTtIf1SqzTmo4liERRckKTHFvwPl1/+Y5pdtwqa1k9PiLfbVZNEC9zxoq
4FppJn8WHb8iOdHJKCjQFsG6HnvHQMW3EDgR70Kx1OwZNGFdIJj5bUG7Kwn1
81of3JOdNX2q1wW6LYmpY6HkiUw5KeGjnv7BebMLNXL9fkJWHgtCtsZOf/61
g9UnQfors2ZhC/jhS/KstKzmnupss319ZtTZTYYJcKH6k0QCUmGWo76+UjtD
fDQ+hd4fPqao7vg5eB0p21kOcC3lE5d8CkRPECbhHlOqMvBhHd/6b78pRgGw
iwSBmuXedsdXeygh+YwNfgEX3phRHa5AMGYZy40YyZ2GPFgMiOhp5WAveoli
2FBqsfstofRMcOV5SJ06UsIzoMMCHr1HAXow5bu/V3Z5fYTPxfShnSOt3gvx
CVJ974cFguasLPDMxcgKZ57Ww6SfbzN8vMBVatDQqisLsSKYVC1iOiW0askE
0nmlsNW6tXrvPkr0wQGu2UHxBut9w9Lnis7QdMYHj6HmzaZXVKLi1PAENCaw
NwSw4uxm3nglkGyZbLjQPDOhepF1drIyt0qFs6/bKeNhY6/AkeTpePoJ1N9v
xxS+ANjwzVJlBEJZOPnHDl+HY65pxhtY89aZ6Fc/rkoRwGNvt8jvrUs9jbLz
wv9dAK4FeXM0+2D2lgRmoE6PhVbiGB4enQcgAKmcC1H6eRAQZjll21Q8trg9
miGmLX1AXqu4XV1MWH4k7vkCAtlhryWJNIXXUml17V7CAkngAgNuNWmJSsQP
C+FVfug2nElFvj5Xlu/PILHmLUFaDFyFNvo4uBopHoi/m2iVEEgDyg4EurKH
VXJc754vhfZ73SsVDtcy985iCMRUzuLjCqIoLz6Ue+c3+RyilBNT8I9apzvP
MUAteujD18dE+PH1zywXU38JKUrczoKD7eNmVzOL9rv+ZIW4DjwCR2Dhb0L1
OJY+wavVojR8U0CR7GncT8CXXUaxSB6NMfnoJrYACuLw/7Or6QG7dL+DuRug
cXoR3fs1OAGiWvrxe0qARB12z1hI54K5l/ltxJOX1/gFl5Qb6/OD8GiCFjsR
RClUWgLb0x2HFmpQIfAQakjWVG7SMre81x76c2zjrsnkkt/Do6VmeOpcAlOP
dDJcv5R+hBXUiBDLZmb2+FewVDRymSvZFf5nByMLHTDDvl3Rd1yK6SLq2PAF
7EL8XjLIulYgSa/z6xNyXNSzuTr7kRfqWGZQkoTc1rO11t+o73YNjEF6T3Ek
6F3Zr6qTHOxiJx590E1z86go+pxTFzKVKnQQvHFWoOlpM9jheiorQMHGO7Zy
4bm4U6OQ3RiAeNjwn3L4qGpcGtooN3z5BopaaPgU+ZtCjqg3/Ke/pJO1hEIk
yMecOR3XhhAbiKn2WMN3wB8t5jrNFl5QmL+XSuOIbs3HdYbHV6pnjIwXJfUz
UImEzaHPrjm7n8WudZDabw9VsXQxcx7vzAgCWA+unKqM7763MSEWXbW8Uh9h
6Uq5I+FH31aQpProDKuVnP15QWXLP8FoNJSXks55RkljyZRUMCHDPyB0MXCy
nrI5Y6kzfFMl4cpZST+l1y75HXlFWWvmW3Kk1TbM+W7j6tbukeI3GAbxHg6R
ZrP90RZa5ObMs0YH5QGTfax0RE7Ro3OUKtej+eiwkIdEQ+EKuNk0fwd0H7BL
19w7cYN1i0xK/N6UDmQCX8ZczBUd85d0isnq0nRYQoFkGnpxfxIfdmPUkYTN
cwcQpPw6bzUZ8NRpnSSHILnViU+CsnY6kDFlRED0jPHgTd3mEBtiJ3ZSOAag
k8i+DuE+URTDrsXx4TmYPeLpK/hYDGpV7R9nrZH/vIV9LNLxezwuMq0ojZIV
8qSNwIbp0pYbfaXe3G3uT5q6tNb+8eqMI5hLF0JHcL45oaABtCXzc4rN+5U9
9GwKbzk5D9ZNFmeu+ycMtyokpQnRvXkVlpKusegk6mc2O5cakuSsxx2NNBQM
CrQIbQcdGG3WU46XeJDI+2U8xDjtUiQp55LR67M7StGzJCIxRtms0XjrMe+5
FYkxz009rWpj5CEN2YkMkXeO/txlQveSoCLo4PY1BEvKlA/9ayOaYWhHE+7y
broW6PJ1tCfsMcvF8huRUspjKCwdMqmZxVOeE+Lq6Ejgw82UzEwK60QRFZo1
8JYsKKKmr3m4m1GJ5CaLsX2AytJRT8mwOqb0aVAm82e89u2nlxJO92az+WwJ
tFvLyAs+EtZI3ly5VYQvLTI1DLobIQ3WWRjcmV5SHKUjzwbXG8zajpzTUo+u
NmJOfWPRan7FXohPOs2XqWLZlu3ITm5yG9sgzRJ7rDLdo0OWu/uforVHP6vc
dmhQy657gxYOXvQ0jOzMgw3PcAMCS+8cKwQN+58EKaeeZqv0iatj4zYgJ2C4
3auGW5JOjU8KSqWxVxzZXMyRiz6qGb8QlJQJFejoS1Rzd/qkbzkDhOf4ELN6
0oI8gHVgpXKggMB41OYPq3W5jQjyScJ+ihmnZxJJzO7qIBFxlgocn3JDtAPC
y/836SNp9Cea/AJnFAQMuCRr+o4oKRr/qvDNDl/NH/RW3R+URwbWwdSicIJc
Wxqn0nTl+i2yXYG7RS9sZ499/FvHLvq9SRTHZO1PO5TaosEqTzrsPZBi+y9V
fQbuQEwIArqUJe6mPjtDDtyFSh5TO9pxT+zH9e62bDqwXp6C4FgW3lyZqgOg
N4vDZgmu8lkBIlfXWxqkSzLcrhbyKURH7lnQNAb4Qo14fadfjSFidwo0t9Gh
2bydquj4sAivKtA/hwnTFf2zDuFMCt0Fc7RIsffsKSTfD+rruC8pJB08YCY5
1WxGOIEbKAf+xrYHSv7Ey1Ab1fBbgU9iu6OvwjiptI3ym6GAffiLyPrcGlhS
OIW21piF/Wha5HD+bqp71z3Tsm/FWVmQKd1/BbI0h7w0y2KeZSsOAWIM/M/S
mvWshgKcuxOhvQXfADGHaaZr3cgPjhzWxSvuiqofxRnZAujxoaJ3u+O8h5Et
ItwwIT2VIqniUaRjyFa5ZCRmvl1ooK0x8BLZaRtTJYh1exv1fGms3u4HAN6T
unX8g4VpHrvo9xD1Mv2iXHNVkCCTiEONVEmYKqJbKdZJuxkHjSQ8hS+N9fNo
6/Y6rd4jwBwzdlIPb3hk5rmZ5I4AncPo1QOxRKR3XZlgQMvMul+Tnm4JMqBg
gC61oZ6LMOVRCu4SMqdk72GhAGJDF+Odzxg1Ny9Wi6JpZLsCpY6O8YezPJPE
Kgs/eO91Y+FVF/KNmU5c0ri1l5KzNQjwvy3IYerxSxkbxaULfRkPl++hR4x+
CVCL2q4GvJlxldhZlcCBAlN50Dqi6bjSdetyBCveKP1ss0itrF71GtTpgIwa
BnTmhHzQk4Qb6AXxmEeogxWF/tx1f17yIMg48CzCm5FlbfX2ND0zycMShM1i
lVxioLDT8WIufTH6ySZV2rxuS0qCh2PQfl1ZENaxy47sIr7TcdM7JfhbTU4x
JqRUZuXZDC/4FdkK5KGWr7kewiovgq2N+kL+gYF2X/QeTY5nG9UMQT2aq8p5
95gWYaEP4xgcJzEKq7y6ID/gxqJPeek1ElhHyC+8Qu8nOcQO3HtqodK0DvfF
kuJR1hBRkRUvJ/LeDZLe2SWAd4nc5HaAGWadMrvqY2sRTiHzBhdROUX5lJ2G
0uCwQdVNUzIlI/AlRmQ6hrtvRtFDRFvA1N80QK4+AIfxvv0I0SHrJnGU8dTM
X/TaQnFbb7zMh4avINbpwTcGE4V09JMLqd/EcoS9bUHiMQweCy0MN43dh+rt
yJERRWwKTa25xOWce3xh9b/fJ+RPYm6c53pLXArIIwsPbjFEdJ09Hedc+nqc
v8Z05JgwfQRPO9MiSuV3Z+rkKfOW/2QZyaQstPXc04UJe4kkOt2T9Efb1Cnz
w8AqungWXYz/I0rQ5udpd0NUAxnHBhLt+mzn4f2Xmxkrb+TlP7NKEO1wyz3G
dphGBkXwK3F/jq5opD2hpewMjKlQs/Q9jDi594Tg0FZ20cpaoDs5MnDiIzvQ
xNLkNPEDNBOxCh7rqWd4H3s9rBjggMSM8eZEDQLo8HUrAOUdvnQP8vF7Z4bL
hCdM9YlmPGez4WPO0Rgr1Xg7I82Y8fZUI8UFnGJgRCIobcdkWHJGfuPzjUgZ
IuGMcf6UBsGxMREU1AjSIEfYHqwYnJJ37ldujZXPi3rIrTJIyxTW9gnKVypp
Xt+BwMyurqiXUhNnGTWuAkRGLQx5GBOsU82tr/zU96iqf+I3zKDy3yA8G5Ae
7YnUQFP295Ov0pWGbWzVEG2aDzjopT8ZStCRBY6tbG11YOtzpqXZSoKHnqqD
wc3sCq7wZ5nCHZwcDfR0T6TEDtqsEZDIe/5+AeipGHY7W/6B0LzmyoEg/sch
sPLQ20eZcv1DvHLUzx6NgRYVTODylEJKiAIEmzRqLtfcc1IL89+ipFdTnUCV
Cd8J0mBtrdMw0mQNQoPiIJX097vs6fAbfWbrB1XIY9k8vBZHq+fLqWJ3yWVC
4dgrt1+Jp63zKOiS2S2S6sWx8Vn0ssp1UIOBVOlEeYDjfWdl7Ps25MqA+baP
0Wp3r5tpDhs/IRbNF3gKII7yiM0SYaAumD6WjL3tU+LVFYZwyNUoK2vvqxsw
WUQ1tbg0qPA9Wj7mq8l4wRlX0YqH9tfFk+evhlz4HEACb3OoFEruEJ1UsLBT
OjFcJHv8I8YxxLzdtk3QLwuGwe11ktaStON3VL06kMx6lSR6mtibZ2RoXSL4
s2HMO5BUDxnbVFWWLUgXVzurDGLyM8+22ZgcILV07tIsvLz0Rq/PdNH0d5Q8
w0RSfUehBB0a4XYbSNoIi5vkMSp7RcH/IJHvmSvpwZLTzEzWoW9UMU9wzEmd
eivze+pYPOKRCZ2pGCkS9Cy9+qHFWpL7ktbV2QN9UnvN8wc7x1lQtBArqvg9
KAx5guSfnSRg7T5PvymlB3S02xib1CDhnHTT833DXjB6lx6en2YathmNziZO
54gNbHE+ZH4X8efka2tsdm8qOcrmWR7TrW+xLuIdR770coO6WLjsJmaD3C0h
EhJJveQhtDwFENRWuxshgMt/vGqHZzxIH92Vdq896QYoCxKnpKfGWnpggmHb
STX2t/X0Bj5057gUERiyjBT/BAfL5Wc8528+QSbE7MjkuAS6+WHl8+FnkDio
BrLaHEmtLteVzJ08Y+YBXvtodRSuHdidQLTxIhhsOs5vRIfcqFPLb5xItTKE
0jkdz84Ps67kzeM0+uVU03+wctQLtTie597ebMzIFbKgZqwb98kWIccM2NyZ
DVEPdvZzcePjzT+EK/1gJsUeJy8VIktq1Za0+tfmL6r4DnkOalRXlS002gvc
p5oXZybyEh9dO3TRmLxEy74t1xIfuaH3xELRMVdgayRi3ml94dQLOCpt8k5g
XSrasQZZ3Ihocn/NiKsw8TIrKp9AylRhGBoCOzWexHLUSrA7pb6qsJCPKppD
BL+j3ZHytxFqJqZOfcS9IE9JU8ULP08ArGbvF6iAMcL0fYlvJ4eGwaxoEP20
UfjWssod4cBNLPIh6mTVg18fFsCg/j0unXuWXJYMU16GTanV91yy6eDTXGir
SxE1tkDlz8S6zk10KyWcgsPG0R9z6jmoxE9S6At05pmGiqPzOhzf8/dhJe34
qvz+YlanS2bwJZEH3hUlz63w143Qi9kuezvCIbOiMEdBH1KSOOfeFWsOBSdg
a8i+IC4Hiu7AZXRJQLmwcfw5G/QnqP8EfDwPFZqnHPoik1gYpcGqwTktnKy+
8Zf/7X9b3EnyArXP9ELkh7/pdtrtsQM2tKwuzNKEB1KB2cJm8mL/LOh/6ekl
0aACIM0IplTCYkepiBc2mV6/60nBtNHR/82KWw6xa60f+j7vZ0MWiYp+Qnnm
7+iE5j06Kz6ASKf0mz8A8elhMJ6HuvxbvFAg9Toagv1BLrNFCsmEFWjRzqgs
W3AAIzo2SzxcRaxaTHdfWobGaEgc/8Dp6pCfz2MKERohT+zxMH9b5h3VveEp
M77WemV6NrH46pOmaebnB0MtlbYBa+PrHv3EBWcmTLrlOfFJ4/C6zEMzQoE3
ZBX+ADIGWGiDRiUyfV9UaXrx8lHPA8ASIOdew+ifWPA7srNYUj0LdhAAuWVp
kslcuv6+80Wb1+FxJ0gaUExaxCBuOzV7QSqXR/fyEmItPXVpZjiuUZvXj9xI
sKPg0UEJofTLSE8wG8uhZBlHsrzcm7gyjdS54li3exEvIu1WnexLJR36XGnd
n5EwudMzlxGDa7lTQp8t3ueAv6r0mL8+0rO3byPJIJ++cV6tWXRuAAP0qIB6
eX+mPjSNyc+X/tpZ2eU4LQRh3A1cu9MbjrUU3vwa4KW66ndV7is/frKyYXVy
8vsJqaUMUyhUbZfgjzgUBdpHLE6LFJWs0nBRTvFyl5xL61vOJv2XcqGuDxhB
LS7GD9SljK+AUwv7MwacYkmt7CsJUooDxIiPUs5ILL6LbLiDE/5EYr6Em36Y
4k1Jkysz73z1rHtbi8MYjSIh8IzDttQqcDze3yZ9UQFsWzUtxmRpDMQPG6G1
6KHivuAwjZrZsHDd59n61urAkKnDD4VRhgCxTPYQ+Q+Ax4TTIBydwgL4AYh2
TjGa6327XhKUSBPeFRyJtlq5pHRJX66mz04ch+gSena02+a8NxANnzvkYT13
38KNW0j21jOGVoFNGD+9s1hoe3qeo57gWq0yHdl4M0jjth/mE8CGvisUjupj
itfCtWcp1HoISoKI+2bvG+FYs6JAHrdgm44h958OInHcRASvmRfRlXR/GIqn
fmvudN4yBH3mv9jLYCq1ZLxQ5DEeOSbd8mcxhnL++b1q3hLyDzGwXAxABMII
F8nyp3h8B//6blj6tyfFiPPDfOM/kN/Ne+X3j4D44OTqWOrR+XtutCx/6QlH
FaER/FH7C6tULGTlEbr0ZpjwbanLwxFBHU4ZOtHbEExvyDBJGBkFkQ/f8ZPE
WGHBUScClJ9KK36ydFck5geElx0oHigtdEZFCHyF4E8hFAaFJW8rJR7qnC6V
0p42TcyN0Teg2RXcw2a2AYxgw4Wj3Z13VwPHr3f6k88WJn01vCZxDCYfcrMc
VXbO6G1PLeFdxPUEwje7XFIpuEqyaA69J1lECD3AUoucrhmcWNn4fjcKmuM5
jrVAKU1t5OXy6dXffO9iErupypny6fEAxXEvtWkh19b2edoE2cx0lYiVT7Xy
HhoiUfTU8zy7xxyPxxVjfWR5Llgp7XNJwtkrXioeK7YxOuiarFE4pCY73AxP
K7srKd+8ngdUhL10UhIafcvc/TVGwvTIAOi0gK+O6FJxjYpAoRz7o6GrJykW
aJ72WVgKCTcdvSeLQkFSujzeE2o6CFZQnyjyflq0sinLozonK352U7+uxoZq
nWFxrPe7dkhzF8EObNs/dEHAn6VW17fwF2sMXSNeTpfKKf/E+Is06h3Q+X0P
ueFK45quanXTtXHYJtrASfn1zSiZF6oc+Rl1/Ab4myuoPVUFQ4HMat7a9Jch
UoCLnuXJ5KIwRohaVWsC5K/t0+xQSUZ8NyxhzTQhScjrvPpC9VI/hwIRvGn+
rV2GNYMrFn8fsc3lHsYcHM7nz9pdORyyiHmeojmqoQBErMfNGfHKFG9ST8ou
H3E5Xj4xCIqa+TT1tAuIHnIxyGHus1ZNep+vRIHCMtledrWJa3Ng6nzgxYCz
xYmeBRiw3Kb9ZFNpxzG9RUhWWMUmNtIEjp4enx+Ejritp2y/oDvpISXVHk0T
4jquzEzUw/+D0FyUehJnog2Q6J9bLMBTLi1Qmg25zOCoMidCmyXLxQiD7EKG
ZUr0YOvwZMmp2Ri6D79mgqdH9S2uO4Vv4fbhHuDi3LsS1ZAV25wtbfdmdcGp
Z5Pa53NAdNC8BhjZUqAu2rLHKPjwA6GQZm5mALu6SxdemEDBz8eRmw53Yjmc
zf5rt1sJehTgVRdACULd7mFlVmdVxr704q4h3JPBDZjd7JQBrbtwk8E4cYIy
uvnxO02Rxes6MH2DrTjti+bz8JWzGa3WyRWn0S2TprVH7310D8I8VMTwshQu
25DL6AJoVdZvKVJVXwDiYqTowNFMMFCPZL3zof4bb7nbpIYf60CWNSeJUFs/
RmekraH9IeZsGGDAO4IZtkFJ8dj7nXtGRRmNcuIQ0YmII/jf1+W03D3cSGg9
5NMOtLmIDt2Bc8WDk/Lsl9w0jIqpCt3TJ40Kz/T3+QQ2dI4VSXk87MtkBqpn
KA4UFM1p9xDSHk/tmbmeX98bd1NyrGhOliljNFLlHmoId57njxiegvtLSnXx
GqGvnb1woup7TNxlmBmX7RHMyzWtMHtW/ZaIYse8APZp3oavAYDAyT0x5Lu2
fvOJMe2eGVc+wa2EyQyqYz8661AZ4TTgIbrJvk8+TDPbBGu+1NddvpKN3rLm
TzVHryD++kUhGaXa5EbpNKiYWQYj9WHe12/yEH4ZibPkui+XEJ0IGpvdTftD
EQtTuIyhq9CwNlx7WGoAQhnpENrPLIkWvB1vl8neTT1fidqhS4F9rkb6nhNz
PAYekB7OPwQnnPKvBmmBH7PsoIEleyegwJsQoFV45N6RGCCLscpm1kZKDMRC
+x0ZrgwEiyteOk6MAJOh4PFd9427zPbzIS4bMntaTa+2IOC1G5Qd/w5w6awQ
7kgE6pvXxVq2CpBDg71KBosgyc1GudWEHlWsUjGnb5RAWKpolsrxY7z7ZPhw
0FEN6U98ujod0MTpDNKr6/qb55lk2rubuf4uiFxNEn3emjlsWWK1MwD+sM/l
VUHUs26rmZa0qKBLV/k4Kkoy/T6c9lFX1LSV7iNaMarA8z92H5LciX3yy7x/
qwJZVK1g3MdTxL3/IAZ+Kfig0GvR06z07B8pyCL37fEmCA4kLiBinqWb2/Mz
+i2HtGrEr5PQGg1cMN+3GqhPb/Pk3DNRqAeYEONKz/dM2FyGkg8AU5veZ74e
xy5QXtuLmKUFoWTB+ikzrXMXhgWenuJZ8Pcl5xl0KD5TRLpuiT786vgiZTiv
M0Tt3nx47rzmM52C47xWXgFQNSBzBCWxLJTPwwgaSYXru0s8j9MTlhzPR5MR
woIc7Fb3kzmq1hfWpGIgyUeWc7XbLamhUv+1YQPtK/WpFF2WYNhMbLHvJTVl
u15Tzv5ohJHfB7hOZrzEOljgODVIBKSyK4zZKXDjq/IeZe651hS+UVpEY3rT
ZIve3umQXQvX96cjrDLoKFdALHvqPyvXbCDrgo457WaMDUe1Z6Zf0DMWpxGR
EJAwY2knShrndpHOEHy2d12SYBNcLXuI8iuq2u+3f9rioz7htlZcG8399ldA
ErzSFOvOA9qnDiYmt6Um1snCOpgYJuMFOE88ksi5uIaK0IAtc2XYa2h4dCxR
li6CtUWAmxrsSAydgfx7lUs9cwgEeeGAL6vtpF6X6LAY7u5FjSxm5bhWweP8
sQqwMe0r0cH5ZQ6iNjY7cG/4TgglCzfh3dLVhZdqoAEXZL/drWiXPe1DGHip
AfIPvLvJ+P5d8BZDKnpKvGKItcF03e89VVwhVpPWHo79MXB2RZGD8MQi7dpk
BGON7y2Wb8LyzE65Qf2fmaDMJ7vtYM7I6K4N+p716okxVq+sDFx/G0/nyVFY
ENcc3tBoQeTlY0dEXZTSJ86nnKpx54yXL04f9ct8VaExUd/CLCO833u6tEJQ
KcSdm/1ozUEbTHnBj0YwQdPloZGviEgHYcR0N1zaS6ebqjtgsZVjrbIqrbYb
dDDGJSVov+pjoK+kNUfXvClSsfKYPOdTUoCzM7/6QNWo9qdAYVY/Lh+l6Wo8
Ew1iGvBuO1mLEeCl6tkTubPuhIo99sfEaz8d8eIRD56wp3UtHBwc5B8ZPXLB
hXywXvo0djq3yAGGB6fq+tzFoTpMeZ663AGqfPFSffCe/alnbTWsq41fLmdM
IjgndyUgQyitOLHjNzByorng6YA8vcvxRX2rB34Q9OhFr5CbmWXq6+myas2E
4STIHZKsyzTlvA6efzIbmohSbrymw+g05PVy9GWRvbhDbll+s5uqRyylLmqV
gckmIjoBP+qwnbilFdFGuUjfFh/p3biWSllOymR0+2NyE01Vq4rdU/jd764w
Pve7q71dbuiqQWD1Y+My5nQKSKHEmG/MH7ONAzsks9VALojeTtR6i0Nn6oBH
u5jG58P8S8iOXaJ5RhiLC80jwaVtGB7KMxlBu25CTkHmrjnVtJ+v+lavxILZ
XlwdDFhambq8UP/FgCJxJrDbvfrkbetdNQTSF2oaz0QqBXsKUAuuhsfdgc9Q
VagvU0W7Fc+FGq39yNiY2OIeQRXXOo/YS5BtMo+kLC8jaAoNZU65lSOPAGnX
xGru0zLDvRbQm16e15RsEl3Fw4hoize8+Nc9Sv+7WEJjGEnCbx/CNqtEHIC2
seolD8+VmNnC4UAi4wn8uGNDTRgnT52bUobTEkRGckUZaHzkVhk9XIgdqTT2
tYLMCzEdG5ZfEA32IcwiZzMmsv7lfZMoqE5kaV/AVPM4+3YRRcVjv2/g/0Ct
DQKHdGmX0MVakOfK80Wlbx3jWFq7ON8LqC0c/FIcRD2YXMHEOmt6nbvUvYJm
otXBJWMiagbtyej8Q/Vgehs2D9G2+lz1qzsdwPhZbujB359g65rABchwSmRl
C1D4zUdZ9K6Hgn5x8ojHPkq0yMlz+pe5SOqJAXqfhQhHSEQdEteyp3dhAhpW
0QiaI54zNq9QU4ge0usQY22Ft9CrBujbHXJEvCsa5CqLzKd/OwDF/NiVayLv
pKWpF9VSnRlrHFz2p97arl1Vqu7A0T5K5VZrMuXaRMXArWYk1CrbE/0Mngc4
7REX7iBABsYkQrQLUGmurneJGaEOFr9tjNPsqXw92csI14mdHC0s8F05o2mt
C1c5tdhNDmhQdup+vTEy40jv1d+3g8UxjP4ugOI4cLlQILu+iSKNMmD1PtsQ
vsh7xBK0SpENP0RrRDDcF/8osRghyPr+jo4V3HcRNEexzhN7ub51gyI/FT5B
wluiKXDc5F8KuxYydgegHo/y0OQQ4sbDyynR6P7kAT4t9WC4teKvDrHTItlk
K7e2e2sgrGZrfZiInMc4jF6l00iLqcs4Hww3fdFS9P5ZGnmXT53HZX+GDsUh
967fhBqGMb+JKzr/xPDb8U/ysA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpegedC2yaJwGVQI+OCOkVckZCMK+w05HMFBHtY1wQbFSqK/3WP6I4HggdosxN7E7AywfxsAx91L/UhP2d/MaDCFcdjWgowUBBHTU6DwIh2zHAZfO0Pbd07Cf9BbOMl8/13O9YdCrJ6FlnGPPcoUoCkVfnkJt0SKODcB2nNndXarWUXZYWvJCjS5lw7ZXxtwjKjc1k8t8fdYPfAJdA8fHQHJuRSEiTXOmfCUGAJpXPYXtIwlr0PpDpeJBMHvbJjeed1En48ZZ2BCIWYipSdF0u96fWvUuk1G+4DNbz0HI7ZSpElXFBe99idwCfIS5zLOeTKvNYZhwdCy/lwgqeY/n0ruu+Rh10/NTGfYZ0n2OeiEr7Rb/MNL5w4XNkwlPb9Igm5gxt8p9KufadH8hg1PbV85tMW1vU8pGOFSQlxuhsQa36+FPgQKCgJvWKBat4Sl4HNu1P0kHRZldph76aqnRJQR9PLA87mNPepv+2Wqpjog42IVP6Z+kOIXrTRbArOv16z6LsgVpWOGmgWnoL9/Re4wNwh8RENLpU7hvnE/QHTMW2G/NALx49j88i9NikcYt4Ug/LDDZ5NVcQRcXY0p+2jjayUiDqt7g3KHF+/NHVRhR3zzjBJRWLnOl6RXU0Yb5iYETGavHUmU2Xh+UzPeMrWo5ZmVl8Wq++0YTESi429vFCuCpa4gMUOZ90ESORaDIKD5/RG3Aic11Zcl6L4cZyqJ7a0b5ivExxt/jzUZJxrH8n2X6KiFBMmAwzgZRIn2puavL49rvRgFtle+e3lazDcxy"
`endif