// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
0ASrSflR0+YxQhNO2TPjdt5rp6pxhqmGaUMpq8OZCuTbWn9P2vmA+b2SrcEb
Beog5KA80np36jcBvIOGKlI5y1EFAufEZ0bz5AoIhlX+nbLabdQHR+Khmsic
zsQuUpcliLeVrA/I4yFylO0xY86dP68gxnO8IHpAttDvK5bxgrK43Y9J2WPR
spGoAQpoQlrOSvFULY6jiKYQ23GxcNEAF+RCt54paXa/NNU3/K/2rMcvVMVs
l/ldHeZwyrHQaRJ7PTq7YueZjVSjjvJwZnP9/HBRyJR8oYHfgkpOI6cSQ4d/
y2m3+h81Qgmrv11zXzKu6w0yrovvk6jSdU3mEYFosA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZqHVdpwQsgDqJJSo5AZppAB67o3h6nv9mRQRidDXHVGiqyO6YLmw4vPPF8Th
k28nDxuZCcyDBajcOyRvwTL7bBFx8nrnV7k636PaLW2tbOeZMZ/DmY4jaaWK
l0D09PtiXbX/Cnm0u3GZwI7KEKZy1Y578rX9XhlO+JOHzudJPgCcQRjEU3UN
ivPcoVxS5dVVLLz4C0SGmUkh+LGaGsJ0L19HzMCuuxxNivn6WFHSnfqHm+N9
//ve0Dn5AIbANeQZxfk0xKAtKqVSs3xvukfCW0it5UVWR01wi69q6wRj+Oz/
uA06jYhtWUeihq5wBQR9vTSmmleGs2wcvSs8pme4Og==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
L9FcDWdNMwYdczQgjl9CGjgRo7FysnJkKacWD9ow2GYOnbPlcLZigZJ+GAiE
vPYnXpoT7/gtBMgLMlv1bblWcIg5/69UvjumoHtRLNCxrPVm9Gfxzdg5uYoV
+A+c82O4vrlpPwnMpPWwy5QTsi0HnAN0YYZSn0doQvzrXDVNCiijhTOs334X
UEScX8yLe6c5CS4s8qa6XRjDyxnZ5EUSnhg1wAlSLXPw+ccHK4WwCXsCAiGf
7QtA/StDMj81MAs06AzvwQoXh6ItlHtEF1hPhYi5o5uaezwzj6RC8c3V0eN4
2IjdEHF3Ctg/gW1AgBiCiGbhdDjfbC0X+AmIMMMNQA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YVvPFeFWWafOzPH2pyjT2m43y8Iye+csj2pRlbu2tzBtjfLMVHzjzwDmD+en
prnFR/ouPsWYd2MVrzQQkh0dDE0k38C68wK9nZwv+lVIAVbUvq6MrkfiVbac
LqCBjUX0k2vv6m/B7jiYgHTcyp9t2JLYznKyaqN8rpv3GepA5VW5VGJ++iiW
6gazek1DHbHHKysEpI5i9ZNxwphn41zkIhdQmcYWDFrdgZoclT4mmQC+OVOv
L8BZxRzF24LJiL3Qe672PJTCPxlEG9Lj4ynm3VJfOs3gAesC3ZgED64UpeLJ
MxII2HMKdne2uwCVM4+1nUMiqfGvqdTUIdi+GWeQsA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FDoFsyr3K7afbQLlGgkOf8BU/E+21gAZWeKt7FB9yXscy5UGWNkagP0TfG0j
06NXedm/f1m/hrLUGfVGY0JxYbmFEEU/LzsVTHTl1M8xLMQEpi6KKH53AF7g
75WsbbTzmAs0vrOjN76KZkd08haZKcXonKvK73Lz5KOdfQ2RhiE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
uuQ/tLHWS5qitBbYyBZuA4gwaCPGthVct7OOzWEmOfSX6OWAoFDBiJbQUqPx
h1g2vNHLP+dcCUvrxwJfApyll/wpFNrNuDY09yJmoDf7dKj8nKj5ZTSRau2c
p3cXQVTS9O6pggYDNIAlTlaam/FAKX20Lkf4NRpL2QkUfBmAFRLpvG4ngrQ+
gXK2I2dfElpCSTgd6yuo2fpah/BSkSxVirdtanqn43jv5yPi3Jda6B1yHbh2
OUBMahJK+0xbA581knCloa8tb73mkXkKA6vPjl82qIfYJ2VDQomxu5PPN3f3
Umm+PeCUbOFK+M4dh7mvFIcJE2JuvxUSggBkdQ7vEhFvx5Y+7KKiIFiUSyEc
yFjrhAejZvwWnZudCwKtkCiXWfG46UBPRRtwABYW4PP/IzajkcC3iBF7CvMv
KktC682s6tgPGpWuey02YH6qoH9DhEaxgvP+cgIEM1IIGWMDYBJ1vPUCuxru
1voByfw4KoaP63vnMC8EcpBrOhPC/NSs


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
A/vo4c4jk8AW3tl2BtZNlhuXWFHC9t1tKPiTHKCB96sP243e2XhGpflB60Zm
njbE8suTM4MnrH7YuezuGmuMDFi93A+rPEcr0IK4KmMZn7hl2mbse5NIiXmU
144cKqUjuF1fQ3yco9kqdC/pQRIvh5p1crRkFHLj0lHubqf2Vhs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
d2LRZEkWdmcDGMG7xdeAS6XYhbfuR9yTWeD9LvZCOHYNfCTtdF4EzzUH5K4x
E96HB06hPewt79R7qSq+viCuc96fy130TACljR+xdGKS1dGsQCVgCHHWPk/y
w29RJR/rNH6D3fg8Zh957N1/YYNhsEsCb0pc6MEvcFL2j+/W3kc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1968)
`pragma protect data_block
H90njJUAcc0f/1R0SlF9RJ1L17J3CMpzNHQ4d77y4YbJOJhh6a+H4fQaxpUI
9SYnxIOLbJ8/tO2c0Uo7WdWp+7Po1Yp1aVpEsnPZ+At9yyV5NAW9kIuhEEkB
kR2eBCHWA2Da1YlLZiJJpg97Uumw40+UXv+/Ug/KYuHRj/jiNCZhOQmmSgZv
Z7/tfaGzNgHQ44Ld/Y4Kr/wq6wORatOjwpOs3yUP/ozriHTX2XX/bO/GXOCP
SMTRJPPObAjE8LGK9Frv1h4gOqzWNy06GjEcR+nxumTmunN1m8PbL2nnYU29
D6vT3qto4QXjGcK4vH1gru37uyTTKuwViV/niFHrCvL8kjg33cHKrbuIPkpG
0klfnlghMpiLY5fCICgC6a/G1PSdbfGlQU0kbfTNvlzozHfcdsueadnH+/qT
KgkKxlnZhv6BbLRjW+eKVHTrIbpZFnEivi1J3nW3rcCrROPV/82f3NPwUoWc
zpdJp6SesKMPaGTUzMLSnZlNSsQ20lz3rAGIQehy/XjJs+7Bhl7jx45r62i8
JFxt+8cu91U3o6sm2pDTBODNoHtm36fDM0rmDhg7sKEBGawVYXEJT7bRJ8N9
iY7H6/Yuq3EX6nI3gVMcMlffeJPCEU21guN5lJA4+F+J4YSH5r0XC5w1rFbo
G6qDXqXaJd8BHAsctMLKb3TPJoQpOwWd87D48s0CmEst5Dxo5NXCMT1XhdOR
MBymmdGOfarGLZG3Q/7WRI9iyqVw9Jydya8sIVlCmVPVduV5XPivuqJWdfi9
2tfWG5zND1REAVivDio2WQ5HI1hN30477XhS/DBCYW57g3MLjCnPW4o19bHe
2HWPJ2i3rw9jFKQ5RhdnJhtVWuAfwJ3D5u1Xs2yiIezt0bXWH6p37JnSg7sH
/jybfoJuAKRekFzJ8y6FWTKjhB0lQgHz/WIR2dDhKGgTuIe++CuEILbdjiii
GRvsC6s3b9/8ge8pHXrNKwz5otGdf7ZCQwFPNCxVW8Km4IaOw4uu3NwuD52b
fD3BGZb83odjjNxZP0/t9tPmV4ounF9ZRxKDZhKIFOXskYFjQz9iKweTitin
BCJeiiVAqq+bScSApuPdYRprzAg773165q9ZXjhZdn0vsrZRbgiJRNKKI5TE
ygNbGp6qvg9gyw43DhB4H7D+qbIllwzIgak569NMgRd4jDdKtJpounqIbk8L
eoNy86BUWYjfkMvrKVikzcBZ9GncdrhFl/T0m4NEN4US/q6IxC0v48P9/n1Q
7nWbEqxYP2DAA+F64f/FkpJqFB4P0NlhZMzlfa3YU925HsiEx6zxJU1kydHh
yVTPdKARnCTdS2CkAXP8q3fGSQz19wy+3z9M7CwwwbpVnpdufdRq7oEgjUBQ
p3tE1UyhJj31VLXRuqPdS3X37PNbkwDpKWa27gI/Vd+eAjAug6/TQq98yE5+
EHKvwzgqMDAIRDO9qQcttoEzR3DhPWqPu9zbfQuKknqRmc3LauIfYeRrAnqd
Eg3J5Vim4r9dzLgYFH0Wzt92q8W3JRn+GZAo8e/rhTrqYtDmYmyIXHSH6hIz
2GdfrL0OyIQcU1Mw2buP18jCfHMxEpGpGlYaCsTIJi7OfpGFYpmBO47qhOAM
oWpc/B9lQHpwlc3Vu6+XUQxtRo+NZlgCoGUeBs8re5qsf7mwLDt2Koc6N4Wl
R5mSQ++MZ8XEz9sdsiJgfUJxV09niAebA0lzvx3+yKLdCkYxmKRQX/OdyZtA
QRG6x+eXjoCoGXyJEx9WamFJfGOxRWzH9P0jPLDrUfsmNtbvOcMgRSJe6DP4
DKnL0K4AxLPGK4voLT7vNkn0jglCWSOcuOb1Y4MIMpBTueMdd9N5hacuqhmF
/mquqVoMvSF9YxJzUkADt0m6+WV6TtrayhSrUE/Rvhr0cXIoaOzT+kN6yOct
ZJiL0SMzJCawrM2CBotHT9rVyuZkHi+0W29kkiPXImo6OYGPtyrPqdMBiN0L
+R5HACuZbmxENSbGeT1tlgygKGTSrgemsepepvBOEuMSll5xMgnY9iD1a2UD
7aNQlN7nTtSozQA49FgQMB7Oa5qm/rpa7nYsYrVb5limYaB8L5wZgq0jJOa5
z3C+PbwdeCQPIwm68jDgGX1Qy/IH/2cRweVZ2TL9IXang9zlhU7KFFpwgbO9
8Rqz8sAs0mss2T4WTUBqrypboI8Px5TQEGFgHFWI6yCME9Xy3cb7YvD75kWq
pVd5mp09lz/OkDQ1/J3b/W2tZCxhf0QVzowLNwRsTv/TfgM0vmcCVXgnS44A
a/zwuQywBJvp7Z1/5w1ANC00IuvMOs5iw3OZ0A/t/7TPAkhTCahzeTBo1S8h
2KSU2K1OA3gKbY73UJjap46Zlkv9Av1rudulL9oZJeWOXdG43Qg2BCsXe7wX
enzQsY+V8gv4oSZdAdlWqq5ic7BdOckt4A2GVBWXbXD/xAElNaIrlOa6cyje
RijDhdvK/VTwFPa0I6+fPJhdFmLENCi72uI5o6kKoRSr+rWTYQSDY1eQ+89B
fGjic0Fi12KvAfbekJfm1Nw5hY+52mGlAQnT1QQWTP/iU20TIdDEZNOMWF3o
eM9g/rPNdEVB7CXRU3TEwdVnDj2zDGPJxWObzh7WyFvB

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Kttctzi5aPKQ6vg9w+1g45z6Da0UaxXtt50QPmQzmLiVao+5Qg/yS2eSRK3c1uFoxS+G6ngDcAKHm0LGGibx4soakCOjaaRTqJmqblCXBo4qigRRJU5sOpNJWGKfxZC9LZLfFjqN04HCQ8ah5FN3P2yNU1iObRgi2dEkx758LbIsGmsSUmn36d6MTHQGWCnH/AC+2pgOY84Iul0q5eg7DNO6RSxNOih+2JmnF8szbMPcfy9lnC60p+c0YvNvVakqxnEZcZi4mUwycdruk+WfbfzxSqYiGbJxESCDML5zjQ3lBZrmsnhjFc8J1+1SVG5IgRbeLkUlZLaEyNLayg1RYEp70cAlNSTEnE97C+DZHX5yzyRTcHEV77LkIRZGy8RjQffu/hiRjg8WK+ebk7xlm64DV04fJnuMloo/DVcFkRF3JqyfTR/LPZSI1dHJKt2rVInx0AALk7sBo/UI3J1xej2xIHM+GmOydWRUpCi0a7kqFwPoOk08nqgu3LCEZqXJCunAS1H946vAYMKp/mtZJfLBZZVIeV2DMUV+WHn2fbCpM5soib7xb7EnXo1bEIvdToxH1KeqYXr4XaRhbETNLtICY+Lj0KIHFhfnAqC7uL2xNlHrOi/IKP8fOeI/GLrIf8CqWuL4wXbeoM6Lf5pLivtY4MfMA82+0cuNmF4MidUvJiqWH45bMsB2KnRy1G0ikweh6LqfaBR4B4Qxw65ZOIDjHdDuZSJ93iqOYXaGB9irNeePKN9vWUeGqVB9ZRc/vDuqe3lgEAf16Kcpc68fUz/jN9sQDiwBJ3DeL8/l9qkHIh0ugHwxZMOgGzejSmwoxqp253ufZ8mkAKiA+449z5TaeunsOQj2fcXzXPsHwBKe4bzXr8hAmHRnUb833vOg0YlgA8edxbrYE+Yd7ym63M5CYdu3rBZ9cLjxS1y7OYTh++bVmZR2OHky7DArs68TbWqQYdLxmunj9WSENJM08TZNFBKvwmBpftKk8/+EXdapBsF+Bi9fgVA/cm1eLswA"
`endif