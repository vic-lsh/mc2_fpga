// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Jmh9+n7KAw7fGGUcsRo7YiC/Jg3b1ld86PzC6szAqg4IsTTuZSydjPf8syrw
F+3NoFpHOekCFnqb35Zx6D9nbfbTORsMAGoRweAXYMHVtuFo88Wuo8/vRgtw
4R6tXeJ18MEe4RsBkvQmFKYAFONsw587snGXuDtUt6qpcltmxwucJ+SQqOnH
0PhKMdDT6JZIexereA9sK88nT/0z6U2YOyDGR8cKlaBCA9gtPBhSPbvh8m6n
uM94600qJR+9YH75OBVTJ78DKKaztwNGEtW4geslfhNFHRWzm3F63A1Df3A4
aWKWtXdc4cVvyxO3tairGJdQQjwufA0GpRYtSrdIOw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Kuh/IpCbu9YMUB2GxdFilVSPSLk89KKq3FCa180Ie99VnEq0xWDSz2iEiWwE
kB7FIdXRB9XD4/EjNK+HOR6TBJ42VPp0BHorIcuyk1pJwv08Cc11AVRSyvvq
hUVHgnv68ow/hSuYyMznBc/w6Qd/vie2rx1BXvOp/OeRUPUHSHCXqgYtBr6H
BpxN+bn4C4H0g6AM6f6eI6FkcfWFgE2JkNdfb1OZbRqsN59tpppdR+XfXcnt
GfpnOhkrl9GerUDobMrZpFxsX66I0firZ82hEiTNa1ZVrzMYDOdzDnRrDtHn
7A+4fqXSDQWlhb7Tk2JANqVjXPKIX4XVvEl6rP7KyA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
tPj4VajylnOckomDLxVKKFsvL4rMLFfkVMMXg1KC/jPAwNsfk+mehnG0c/Ct
pVUsN2CezMVYMEa9sKpnoUjJQv/olumWzhHK2XpDj17W+NMzmMmp/wOoSohe
tRG176bITmPGsGQ5tcIXuna3jO8NYfP5EHFfI+TAsWadtxIic80NWDCYydl4
stCagGTZEdI0EEP3/dBKTjahWLviLHA8gR+ttDuG4xXM/hEytal98erbp/Qv
VgjnHfPNj9LfZFtLZ2V1ukKPhixiQO68jXBmoRtPFvbLpGeMIbBc87+S1uEG
nIApB1Y+/NZ8M9vXC96u53xnZVEc7mSswSy6U21nwA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LqrhgsNsxVJxonmS9Reo9QT2PxIuBqs+loNwlOsPlZ+v70YnOO3b4XqX0Dk1
eOONpnv8kTb5wDPwVEkBO53lja5VBBrdDIEJsXnNxNXhDcKSmkIAp5yENdCG
OnlQt3xkZTRxrgv+LlrkryV7lxdCD/JJRRUROGPKbTU1Hkf3lWrbdfZYZDZp
PwZAdHNNt1CrJF3/tbPfhZ2VK8idTM58aDUDXViw4BIxoAJe3gQ8x0GyMnUD
I5O/cphU3j1Kdb003V/LBSs/OkuNdDmiE8/Ni/9qAxwHSmQXAoDtg4lda9AO
qEVHF4NKJejwOv23CrMontoQig9PavVSmsUmsyzzPw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
W4VSeSvwDNsmBLsdqhTDRoE2Ud3cOBDM/qFPPjU2RuBjiLDagxApAFFksImG
Ktl2vd58coQckjNogtPh30QrcKXaNSi+AS4qAwrc9BLaiFBFux4vEpf2A+QH
hSdM9RWxwLRxt/nrRcDLR8LgkXqOXZr/jKbOG5q3kLSeMGDbLew=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
PqFAFH3dXjJfSQwxpC90Jxw6KUy1s0r0JJWh6gKaW5+YhcnxeVvx8Zw8wWtP
ry6DGqm0BYVfzsqpq5naVJ8PY/uDyGO3EsY6AnpzWtk6C1MkdzZcTOEoumKX
3hKShRZY0LkoPjx1jiMeDPHpNIr/VZqAUE4viDDYvR2uU79fuIod8viqg7dl
nn+33OurLSRB/inynwG0JlwdoBN62d8dACPR08tSCJZvGr7HR3dkyWrxcM6/
7XwfOHQUasTgVxs4pXolU6PKLOr3edTGV0MERGf0Q4K2GccsGhY8GKsTsiiM
8ieXCZ0Q78abdiWSfKaOGVIOk6W5XXd8nu92wf1KYVFIH5QSDeHl1fqUBs6T
3LzEj7egeFSi1NP3SRwqEP0v95WFC7k4/bn6XyD3lcv14YnB0LUcDwRxLeRM
EvA9ttX4EM3BcGdH6OEaZRabHVw+BqKSdQ4K4vHoj7lN+vY4aPS11qrqcx28
Q5sLgYQjQaOqfAPuwavrr7NakUcc3g++


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ipz5CyrDgvTy/gioWxyAdZpdCogLAHbKGjm3WYmnFqvHnVDSdJwD9qZwx+jY
PKzbBmfmyHVfoUDgsL65UuSCJZ3aVdDlTPGfDxGvllPWv6wj2lxkvl1lrjoA
d4ywyR9AtcgSHSadu4qcn034/JW0PI++sjeOcUudZgus/Vbc9PU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Yh7zOCDcnh77uDli2BEWNtaz0FtRsto6l7QoOXLdNtTd+PVJ0vqlkg1A5z6d
c74T3pytvuOp/kjCdWxZ0DMKVt8qetEG87I3rB93KOB/pjy7u7cOZP5ELHBH
GgYbPGhVNb4hSMgKqyvphYkSUCrtpCQeNGwVtagbNT/OCAwgLtQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1040)
`pragma protect data_block
vhsDlwI82gwruW56LXTNB2syxKs+XfMJkjn8m131T/CL8DCB0Ke2+d41BJXx
j1oshb3w51AJtXufB3+EReALkOHv4QBQ3DPuwkvZW4z9dQSIrwrfSoNyG+3/
vxKASBLi0Lqi1kPpCfu8GVul9qo68jAz5BFpuyam01HCEUcwbyjCugCcX7y1
55268Nh8chGae+76pIwJakudUHZofNz5b3dFdhaxxcyVvCbkEFLrVdCRTJDy
H4gb9yGcMZvIREcZ/RH/b+aHOWO83c/y8t9pZJtcfZ8fwd9YMLdhYVdPP7N0
RSUCOaVX4Oj4JcWt9M4DvCGGStWfDoR5M6f2+5YM0IpCvww+EWR/L8XTWyoH
yJP1EKnka8aSNX9fFfz1/2wpyWvsXM2AkE4zYuayS5PdFwaoCnuGcZhl+tDx
vL4Cf50O5rhEM+NQtrxSuf7charCQ5E74a85nXwKRAz4dgqnuThgiUcYh/Qx
lirLCP4c6dRZO59jD2iYTUDn6yBHqb9UIYYKN8CaYz2dJNUuzX8zNKmc9Y5j
dR6ZLHMjIQ+oP/yL4avLKn/Jl7+ZmopbZoPTp2j58uXTEYMull+N5v73Uhlw
/jUx036xdDH09xIIY3ABKW7nf8+tPZwd2kfFLw4JK4rNwZgg/914aett/zVr
/7cR2bFdfUARbnzM8jpmOx1Jn0hQvPHryMXZK0K2kSKDFYAG6lRvFCQcJhw8
ewHItliOWqzbZLyB+Ahz/eZK0LRAYlzcMuhux8FDbyzXX0yjUTSkE77lq+ND
8jQZ+DtoGUzpQb7yhPfxJUAHxmFeJfHf6+RXrVPevNDdP66EfT5+K2wtcyiB
osvl9GRimBzDViZkRKQhIdtqJTlY09MhYDWujyp98vh1Of402Dpp0IagqyzC
Z/9dEf3MfXyWtePb9YOhegwVUjmJUwTkvj4I5JLct//6xJunEtX2H239XcBJ
ZsROd8PFCyJ9lPF70xxkRtChmQQjbQYC4I5S9VK5E3zMKoGx/iz0qrtInQJ+
xY+1wfCke4aF+46GWbvvRxXamvyATiAQKRCsFTW4j2Y+qaRdhU+uYGePJZcT
nmR4DQJY87viwgLMVs8dzHkuZ1ukg8CfTuwfwWi78N3Ft2vtEGM0YvD8cuff
NzUrtqShljlNMs5655zQp7fX6yYuK83fy27xDHIwKFF+SJc3+PRPj44AWgSG
UGqbUMIcYIXNoeFq+j8QuMHfvS2b74aAvYYRpaHLewCqUmWXO4pAmUEWu03S
sjhRyOF1QGIJmtDNJGrtbx19SPHPdxaAYAoEHC2frfILRMTxnPP530PCl+MY
B5dYadYdSaDUCEX7eA/XOOPvs9wsKBvEwm3GiJq8fCPqwAqzu5WgLvxu3Mh8
kgACiOA=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqdkIRuogBWqSVRwsYejEMZMpDXx+AfuREsKpTAQgsJBsmRSPyo1wvk/Gg6mEsM5OOGPPHfEa4GU5b8A6f095Ywc9uEEucTpLUTdNh5FawlHGA4x8+lGvrwolOY11gGNB98aEZKxpV8SmQOsJQmqbqFTANlQvtuKlNG7dEEym6malpY5VhIh2IEwyPJXVKB8YIywFLgNbc353LGG9C/cCKwisoROiORBEYOGhg95jNSRAvVg/JYEyAXgi7m2DJlOJJ/z8oQugMzJ0AidrzF/e1xJoPk7D3Uw4s377crCB5dsSV7STzOLYq3qjhd8VFEMse5+WdG1LeQ0DtGnq2pTLqr19K+VHt+eXgHaHnTydJiv6s0sYqhaRh1MvCYtkk4M9GunBT3UbshoCt8oRHHlASMocLVNpAPMgrX//dHCbBaI8osX6In9ANbYjZPkPf1EUxMYq6HXoHCcBygO19L1kqdSyvlrqwGxfmNb/l0UeO3nihfHkOSkZhdjS/Zpn37rDLvBTTEMtfn5RRF4hp3lz7XK8yGa1iRZPlng/dd4jm2P7ja7oOsVj3oLxQ9Y20G5OFRX0ytlxmjlEUyewfAuviq+9qz1aAdf/VgJvFXM0Fp65OUlZz/HJJYClaUVTo0LnVhdI60bnR9gfS43lgEADyNDd9qPtgFWl27d3yHLGnLlT7Swm0HHGXcknIbn2TuR6CpRqQNkNm4owEcUtHowUgwOyVcNVw1qUyTSf0TB3S/UlMP03AwKTaz+WxK54jF/S6cp+XObYKzaUM1Rz+sU+OP3"
`endif