// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IP++Sph5VKItnoRyl9d8APM7CbSU+i81BTg5ve38WcYxVzkO4nk3XVYhn9Xn
19pUFBQ6LoRrqzyYkWxULOcXpcZkMlKrpeAGeJZ9BDriKdxnpA+UkMwjWxQ3
xA3niobcsrx7qrHeT2uYb9lzJmWL3btNsirwXbgbWuGP4mtAqaeA6XXZ8+9S
nl2GOSl5dBc7VIZKWBXtDvoyDIUfti1rlv941wRMORNct6viDOkqaJROg5H7
maYZe5bnzxLVqhYjzNdNxpDP5V8lbYIO9qxHJxEzXDayLPviKcbAaj+22CJG
V0p1bgINMlg4NEqW0nXjusbPjEtsRmpDkSC8pa9RnQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pvvLwE8IJDGXqpUgoP2tOJ/J25XVbOaAEj57wLzgTcQ8b1pMgwozbK7ohgKH
KsLxmwj6CHogAYF5w3mEP0FP5gmAY1OxIT31V3/WlVJChlAU4UQfPbWUUdDP
7C0DdHqv0CPuDaM9/kD8PiIBdleCfHQAl4UPcEvVw7DA37AckV6WhiKr+Z4I
gAvUPnjbWKXOXDC8m57mSTJRapjsoBoz+70+qK/rZTZi+MY6jZT75CAEH/Ib
no38spw+eq6IZTNS1X9oB8qOls3ts2re1Q1VMoOm21FKmehlKai23tdNgk1K
h16ZlnCkUfdGxs3uytgvtC/d9PeK+H+2lf8PQ858Dg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QF2A6VtmLOnMHE/jRjLefGnaKNS+zO8qHkCKGPHPqdrBHHZYEmTmOKZOReYn
4RDXiCkDt9tV5+KvnSGbIW47B5C9+IBpe09QGZczaTjwzfMofb62LCHrwNNF
P4qfw+/V3i1DhgpHb681rUXAmQpGx+BKk8JZ3JlGQskvOCyTsTWggDjGWHgc
vT9VqHzxn1nkZA+Q9/7OoccFdMe3r6oBkoTotratUZeq7WVNjA/9wxDVZVAj
L1M+YiVstkwfTzLd0jri6j/nu8W22jMJhNz28qFKvWrRq0Hn5AZBR5e/8Gpb
qAnwYsDV6vcA8lcYMdPMvOllRtOrauqeloPq0Xrtdw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LdCXyQqK8ffcnzIeP7nwSRjhTIjNIl7HRRQGKiIO71T9u3p9xH/NhJP+o3Y+
ayDWuw+Ff9EZ0niJgiN2TgdGIzfPN/7RrIPwZ0XwJu0VRsZYjBN3xK/rSTN+
OWvrFkHC11nDMxYY7cc5WavNHZji8LacUXSWRe5TvQCWXyDug5adI1LGOwDT
mfRkQOSnhoHMp6MrQEjg3dOZkzCsdlPsbIno2c8VVVZt5aUK37BYATfghujd
rgDgOIUFvrIvNhB2e/Gn+YbE+ZUlZxbHMNOIt5hiCOVKJsiJtG4e2T7P289i
fpP6W830r8ea6tcEBfKFngRPk0FCwYe1TU6ltb0Dsw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LFjsWkY2wNmCwFUIsr9De33b6HTSTDCFykl0B8zUloZLM/2CaSYwjT2fHDdJ
9sSr+EWqkoJullDNFsMBXSIOsxSiXDsKLsBZUY6xHKhjqLVnJ4Xl+T/kcpMi
diQcQ/3bBzcS+cHll/poDCB2Uf324fU+z2IVy/sN9ZJNOh08Bb8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
t9fZ58xFnEpGvn9v8k12RCPWIxDkAYaWgz/RfEEXLQRJl11LHxLmc7XmgVwH
Q3P31UgKFqQ3YN9Gl7ebxeNyz1gzz0euWEdhS1t9RargQdt8DmpRoi+M5Ozu
eNAAueV2rNTO9teGoL3l/fjn6PqQR0MkXJHDA2ah7MJ28l1OKIClPjrRDKLH
SlAKRmXfD5GAvOJ0lukEin6TxNDd/NQs81IFwqZX/hQU4NJq1bcfK9QvDkOq
41Pzs+Q6yJbGvJPZ/+SgAKTdflLxHyMJofRw3rxP42mj1ZAbfpULXvGswnxb
TLgjGb7an2PMO83/X68LY3R0OuP0AE+Fke5B+4qcg+tGp3R5pzb+gA6tDdML
iAwJ+hyr9Z1OExTLOhUCToaEqHy0imCnphkpTxH8QrUnly71W5SHNxv9t1+a
cUMjcrK6pP9T1bzwusAdhaSm2qW2KXItjFU2oKrc6p0Gl27gT3l0Gxie5FFF
D0CgQPS5G2xxXzuuo8e7tY/VtXCQDsr5


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GIoTT/BLTtdA2p6a4cTJq9+e7HRfDKzUTwjWNqp85aFCapFg+1B/Iuu4gdXn
zqIOVS5ElrLYRiQVWROssQfOlI4tdU0RxHiacvSA1yycPQhi5l+G44A8WNiH
H0lxFJcHEry8WcYmhJ/IvbW2ZCdb38aquDTz05zmUyQecg3uYDY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pndfApgldJ1iy+1Qj+z+oBjbsLSXuopFbnKcBC/DHAcp5ywr5MSER406JzCQ
gu/z8cbZwhQySgAJWqOMBhaZZddVD7VbSxEHHOSqawPfSIgKx5bnAqEV07ZQ
iTrI2bJK7BzIh3M9sTKnABQKs8z7ROpigBxbD6Pi9iBY1kh/6jo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 31264)
`pragma protect data_block
BnbxYHXHAFKOUEUqvPcR4+ucysfVRMIZGhDOaSI1tAr3ekBVzv6yxCd97laN
Pjsl9mYam+tWwU9rLv/dO77bxZq4OHEwYfcVO8myV4qNA/+HJFbpZZ5kkqfG
ftEeDhjjlPFNUsS0CzEGBMvLLLBGCf4ZbgzKaX/qpM7c8m1x3VSypACvGnr+
C0hdwFOpYNXANM0Be3ZpSnBGUfQ+BIgVwxGSqoC+j3CIaMz74q8UaOQKdVGv
57ZFZuGKRy06mANDMPdrAJPZe0lAEzEf4ttYM9qp3GjT6xKC6nVI1vyCfNPw
fpWoPKTyEGwaQAJoOy1ahvboXNberpTaW4IXinK1nKw/17sMRFDRD7CjL7d+
IxaBFM4zUC3y2PIeQoCAuhuAwJDKUc9Q90/GF5eIkrLxuEzlK2d6sEIen2E0
w0Tv9+inXAyXJcxsXOBbTBELSKycqb+aaImCbPymBbxAkEqj6JECoRrur4jm
BKSBGJHEZcTBGjyU0XwKzj2mELxSMUuM/A3wYkTFdbqc6duJOARsohNcqDlP
N5Id9ru+C27j+WNprNMh/CPVY5BEV+RnCoGT3KeD5NayVwLqdK9sfWRfPb6g
eQMoXbSRmqGe8/dVx/7hbeg+zByclDQM1DvLqLj3sMHjgirtWqtMTTcLykkn
7FHvzCzcOWkYb63j4DNPPnVXf87zePQAkdbt8l6twM1RBzTHXTLfTtFZYIPC
kFNmwbpVAuBnu57/RpIUyjE/sw4fEYvvNIYcZdHXrnYqxGlOD3OPfOjqoiSh
qdbVjNH+i/ProIpwcDAAmr91t0rMSVAdaAsxe7hu/uDCtDYShyTB5rSi8Iuh
wXjSV605mI1JqqkSI9C08h9M+t0tqXrFUrwrZFLP3YJFKqfrGiUFljchjbAI
G1TO2nWWspav/V17CgjU2giGFBjGgnDuok2puaTZaltXh2pdKOZYG6vNkhmt
lCOE73ppLqHxc+LEhbSe7gkcfT/d5S0AaW/2OxvjbMMFp02VilYvNQ7omRp+
mZyvdB33bH0YOdjAqvR6zdHcIBbdUe0fmW/sums2Yd+s8SkQqU+k21g12KpR
9w9X6KXb5iSgIIubd80OcIqi9liHQN7lR7+vyRdROiJL32jxVG4hDH03IyQi
15OcXLT13HDVp3z5Fa9Ep6Iw5lt0sSlGE4IXc/9q03wCjS5HZziPy6cq6FVK
7TPmbU8AaELHsgfh2CjkreNbE1BNIi5vzhKihbzC1M6K5AKyR3NwqLbJcgYl
lAYkOpq5MIJpBb5iGUIrToacPiBGzzqLGX3PDlDuVAbjgo9/OcuhWNeSnwW8
Fc9/s2QazojO5ihqmqrTwbmNsc4SYrAPNxlr/USUwkwJ4bbay8eErCk/9DXk
puhMjbAbO154hj8WrEAWTRdeSCQ+uj4bYqqCgn/YDJt13O25IVHhd7/m4j4i
EFOMQ84+5mccbOdlCaVJHxlMLdIaGkCw6/xkdbRl5EqbPs8Outqa35BDrmPN
TgMA5akubtsUUKQrN01eNYtfC2p5ymmTwY/QhqANF0/9gmd6eQiiOC0RHjG0
IE59bjC8eFMsC8D/75NsJsrfVTPET1lbejPSmJpPNDlKo4lmGPAl047ZE7kY
IegXCY1t2QrV7u7jKQZ1vde/iIzjdkBL7yG8b5G5Nd24QG9zLk9xDidUpBUF
8v8StM2zZCl6EJW4a+z/UWhN0C5KpyzU3BhlIxVBfEtlaFQRNJleTX3Z1nCi
UAsqf9lDeGOQQXDgcDsQjP7SyfMr+Cs8YiM3uqEAwqhM/TbKYPPybHT9g654
C8G9H5D1dDrlo05p3yDS8SU/MwpFDqvkJm7eIoaTMa8aw+eh57AgdKRfNftx
c01y64Yi/xGso4NB7ZDQsHmb1b+aVHPw5dA+kRAGd/qhaUR2WZTtoP6rSvXl
n3eDayp/Mh0C0iRzw/BKO8QzHo0ga3zJZxWv+QZfPZhfnidzX/h4rjZ+zFNJ
IppEmnGTJPQWnsb1i6IOpV4aK9yln4fjvN7aBB66Ls8aFHQXI5VHZAwjPtp3
Lv6MyYiMYGGD1rgUEaMMb0oTnPrZlawd3u2js3K/yXoY/eRLp9dwXuwMMMfy
2MwaEdbqAuIKT/oN7NEgW4ZJn+dtUcvNgy1gampU+g2HhJOSNM+Ny96GaIuD
qkl8/NvF20LBTIVay8hMswcCMnWsE8Te5yfZZoZ0m+SbKHTDhLghg80q8abk
PSZLDIRK9v0ddKl1+KJFTq5Rt1RZ/eEvXK6WDVv2qOk+W7M17XuyTDFYYCTO
x4ds1I8T5dSIVUGE4+rQiNp46NGPgfGyhqRNf1YXjNiSrarz4tlVnSBwyCf+
a/jvHQdiNLoIA1OSN0ipf1GmImagZVSRgmdkPfWPPRbfl6G7VZsdA06vV2f1
n8ULPvFBM81LDJr10yqQNs9iuQhl0ii/IwCfJiVhCUFfaXx7Je+4VJbGXDiu
3fbJSSm6fERzqyrtcp5vv2fV4xbbV2ZlzWEVQnKtQjK9LNzpjNReuKvyA2TQ
/TSls+klJSpByYkJBsnpUGs7NT45B/OihMXzndRHtF5pXE4vbo3YtLRXvH9a
cgr3uME0YfL07Xxan3hUZL5Ma5NKweKl2izDcwsGqMOyvmlPJEeujgnq4b3g
vkP0iMvaAth1Jf53Iaa+N+YTSQHmyHwmiCu91TamBFaBLUUWZm8zHF7k9fTW
zw3MHCLOPTwBOOxhtNsI/5H2Ty+Mw5vyOa5s0OLbC+7YraoAdnmGZmLmFrhk
s5Hkk/F2ST4Xt00vMKPSl5ZyMkzTKZ4viwYkWhGjroGP+I75M2UJ4MIby2tK
I20aOg729yNhrabbjVverqrXOTTDznElhCwKU3tEosaVsqoGwUWobWMcgM5i
7RsHH5tncVnQXLIxCDc8YUivWsYJr46tD6cP162eAWrcFWEJiBPco8GHv7z2
FBfFTWtjFRfltTQ1fAaylUyfpB/ElLqhtpLHE9nwtAuS/F5VhQwfJgjIEyyu
lYajEcL1KvC140nI7FYOuBk51j9Xp1Lpsar0nSnirC/rlNjoIPWM/BUvejGX
xwDLCqkjaFsqYUi7QLabqEIEv7DKXOfntvCQZBTdnsr6ZYc5PJHnpEpaqGOC
LkrewvnBEouSoGYwBe85R++mpKY3w95E4Zz6X4SsVOorcG1M8OpGX01x+yp9
/fnK2rwuK2Uj4lS2IJxfWnBd7V+SZJfLA3Ifnx+PAobpm+qr9yubzqepBApg
hqZ/K7nBwE2NCkwUMcjY+YHF1SChFfsyXo2DmQmakBxGTh+ZnqcTKbedqsEU
jCOiQL11OWS3UVcK4Jxy9YoTbY0TWIqYwHQ++D7vs+2xHQrXRqbpqcNBw7Qr
rmDC0v/RIyfp+EonmwWC/kxvfeY4+AMVf6CbuXm5/ttqNIuWi2RFptLi7auy
dthB/I4e1g9ikAVJMvENdkHXhLj3elRgUn/mIOvI9pgf+zOXsyidEyyHDWgY
UkIU9dqjyA7RNGxFWjRdcFzPOHSicUiLapj9qnKi0zGVFeDAGKfAc9FcDSf/
IKsSH0nImzyZY93IWzod3OhNKkNQ1/cVGw0gSEtqEKi7UuTOF6S3IcUnEuB3
gvCOoN5kuCwiW+beWI08cAMwDJkuSHqN+e+dA3jTtlUfFHrLRxTbSWjsA0Vb
JMFFI+e1ibKRGiWhBWp0qyWxSrSP8l2YfcCK/q0v/EdvGl4j7CjfjqPJ7dtQ
bYGz77UwRwC9FfO1WtYfhpQR6+bmTLLN8cB29Tova5zsu1//dfjmdV5B5WYA
9hkktkg4/NMZyAagmB1vgfKy47WxxtAavM7+57TQXUJd7qEkN6s1xFZqXIlK
dWlAYr/w7PEONIJAEXQLoLw8XeOLZ4MMxkpk/BnlQEHhd04YB7wN1U+o9ZmY
+lzklmm14Oi1qHa0g17WkM/2klRz+blWZMLlJDIZ8uj3tT9cdGtrxE+3ckwM
dwEf4Gu5ZV3+2qwUdyfxeCa46/V5NVlOzyqT9lhlhxU2o9cYQf0SlXKp0T2U
zA0Z8IW4ZWbBpVubBqh/kv4TgnG9cdmF5mWQ3LJG6hsMfQYV1Rt125h+5Em1
6Dzaod+ODfaKdt5qhPAJGg+435LgQc0rrJo6g+Inzg9q9/IRdnPhnOABEic1
Z+gdjQ3xRluR5TudfRrUL74vghSN3+L5b6iD5fFQeBtFB6sMstWl58YkWBdM
X4mxn5qmbpCjvvM4wA9ZlvRIkHqKfDN7l5Kfu8uEd1cnc38LhBm1fzx8TLWB
aSQMIRo5oTQ82uCUEB5bBHD/azJZ87BhYNOXZ+4SStqF/cr/IZtf411YL/pW
kT0GCHL1AxjHjq+kekUe61GfSbYv2L80b+AuXHSD4w9Y8tkfyrKvyrNtFeNp
9GhaZTca+fP7ApCYgC6hVxDaM6Pry9XiKAwW6fNslQBXGPYJ/ndhVFVqcpBZ
Jr0vJv6y9XET6cearE4ZEamcnSfNun3RuwhKdDIxvd15rGeKdFg9wzasWPus
iKON6VBzfvIhM2mvZ+doiX4eZ9cIdcLngS7hgOtz0kKkCbGwb685FBi3qj5Q
YtdgZHtm/jC/Kgumv2OGGeRON9N6ugW1s4di41YkUFbruAHqz63jAr+pRtX4
UNLRu15c6dOtfTBlFJyXdbNo8lr8fe+35WBpkMl237fQe6h8r1XmEgrBeWie
q+AgmeirWAKcH1ky9kr9h2ByQI2CVpGEdHp7u6SYUWL+oPTwcKYRjV15NFVD
H3LGO93xGpGAITiWB5Xuk8Whqg9ZX/kjsjwM6b5NB5P3bUsdyi/T3FJfIHfo
JvvBhURfQGi18EVWBu0zcv3T5YQ3uzvmm44o7qzaY9JcJ2+KpjlwSdcPitnt
LY8/CKKvRKJ6HY9vAR2H12uMjeD2XJ36dWIWGM6ysxwV//u2386tyftAXvlg
g2mfOzzQ1QXWkYaW8HgAeWKpoW+WIBaJGNCVGrUmvjYVgxzEcP+Zbd5t3Js0
u9oTdYOGdvNuu8sDYyLsy2jIZpwIJVPsLvVk1U6Od2Jngkmal+Y98QyyYCG2
FjZVC6YgRKFcxYd7NGmD/8wQG7S/2AxmlyvBCs17eItJyujuSENfWEnR6NQX
4TFAnhiIKU3+s93v6mzhov5M55np21ljN3QTXSLwZVxnN3DKBBWKcI+zul6D
0ipI6yjoS/7BHlSY7YDDxNo6dN9NXmexNtMrqi7c7c3ntohiZzQTsr7iD0iY
TIJhUUNVPI09cpHJneoLvVf+igXIun6bm500QznBXdb/dpxkAjnBbP5vJ+qc
S2LyShYIVoyzFoEZrdPyktoU++ry180PMX+JhR4mEdU8naaZYPdvd1rWSV9Y
mMfCP+tpwxYOKBvGsYC7FILS54XCN5jN/MMjrHeLi+BzRxSMiKd9VciTQEAa
BYd7nwPQ5DLXcMTEfTpUyZkqsUZnGOpM3Cs8htWuYjpC5fvKeEzYPHfOEwlX
eb/8PWAXWIfUMYXQZkg49EuoHd8TN/qgkL0l6rz8woyx6t0Q1NTOIgUz4b9z
d67GJ9KlSlMm3OQ6rKM54K+LkPi4e9ViD+SpZeF+kSrG+7u3V8dAhUrziwSH
DDTV4dvq5cCnxHkulLgN5G5zvG31DB2uGQiHPwNBjknkfQzq3N2pHJoTwbep
H8vEnG0XehE+3hEwTjo42gb8J8bn4USR3gH9RyMhWCMTdAXZnTL8y77L+zPT
J9/rqJX7tguNdAtNASXA4pln1ZDww3B3y6ZwmIzywZPwZE4KIHqkbBX/NCxf
3MV4WJhJ8AvfpjsCauv2d2wzLuJ5bW7BlhLGS3qthpX0zd6p/h93TpyvdNdl
VKW90/C5MijO7gak+PceJyfGgWBkqW0aaOHydsbcwH2iXwMcnYYqW3vhsPNT
XySpggmxfCNsoOnJ0Y1+JFWJR3N9xvvDD2KVtGUzQrQzpHbq4tY/btY/rP3s
hmDG806NBkGxCdTGTa8A7oCgSlWGIs0eYObenrn0UxGR8y/UVtigfxeOg4UI
6V68PMftz6GgLmPWgBSLvC62D3MsIUV96HT5rPSc48BChs8YBOxAFfF5DjgT
BtsvUb91aV1fnJZYpU7w2wzyFu6lOT6+hyxNxabkQfS7ME5XGZP93LTc1gcA
7P1c0rzO0pM/JLIY+omyiwX20U5/WKtasmucCJEewXAklwYBUyXwXmReIwdZ
jxG8uMBLhYCIrG52QVEzD4SVdQ/1tpQZgAMpDISKg13IBDcy5QQbPsK6Agdc
WYiahr1dPp6GnKgbiLBsWGqbqmFgKE8UuSoRdqEz4tpyqCy5HXwqajM3XdtQ
2F8QRwcidEXVgaPxoTEI40K3DYCikDKBHfEaWUwE0oaY9E05jzA2SfSa7SgF
NCv3H+bXpjKSD2ybo4hmLLUJCKhRS1oJOExwmghaNXEdNKY/x21tVnBqAX7e
6ClhMpuUTw4+04R95ZcW+xk64OlYrggcIy6uf92SmQqFOnbUwCVuas2wDnUZ
a3NGK4xnSamASrFTJhOKrZSWuSyOWtlKufOMgk7D1OWKypTCsl2HGI0nwo62
1LHuog56FltZ7mlrgiLFt8sFUHg4T8AePF7ZGtTDIrXFT5TX81gDvOfkbMxk
5GG6uQ2UJvDl3gvSEg5t260oQf8EoBd7EQlqWoRoaPPwZ2rWkz1Dzzhl7Ndi
FBf2S16hTkAPtDUHbNb2t325hu2rwK27/p7WdWj1xZgodz8XKtSJuftaDg94
vyYxkHGN/Ke9gbksz9jgpHfBrwxsbTneOkzK4XftzVPHik2SVF6jHo1wFUE9
HjQUrIbVoUI99gUm/2jPoKcZhVukOkbdrdRU5UcOuNxXIylsyYB8jwRORlPb
ZFqYurbTuNIGqP8HZdZSC6MrAsnSgCJAoGy1ll6uutyFOzDbaMtQ/5eL/NC1
zCW4iXdgZJ9bCjksSPop1UxtWEwncjRiuvI+co8Uj/6H8C5RfWJFflpJchGA
O0QfXhco7Hzoip2xsPXBVAs34kTCL1bn4UFtQtmxjyV5H6R9Txyk769RkCqX
tK7AZU7o+xrzh2UZRDRVAtj6FU0DqeOXNSMKqOveWqEwdKnc78jWnsz08DRk
Q1uW/BtXQmtny/CfMb9kq45iZDmOZ1/Ov4IKouUiD7IqrcDA19iLgKXacP73
NShkJ8S4UXcsdO7WWKQoXvZJK/SzlIFaxbBVk47mdDJFXBRzNzRs5L0/z1YD
QYc7UdU0oIxGV1kFKy4l++CRV5atsOfw8gonOwPRvpjjUajv3lB9kB4hfNdm
g/RLsoULvMFQZKbtpMkx0RKd+5u/mZn6NiCUb/5kbEnLD7EufXcoqqIGYUKG
8v9rVkZlG6Ih/IMmME2Fm90wIcMr52mCTON9mV4IaznCxCf3esiI4KcGuge8
GJHBzL3U0Kcotnyx4F86gtevpSpD/pyXwkU43Ywxk/4HSmPEiimO6yZ0MpZN
XdZQNV1vCsiEGaWjz/wbegeVnrfBxpWwZD6PoHiA8Am9xMVAXLeHIarajQ8d
DsM1ptu6e5pNiF5b0Gq5RBAY/jTUnhn90Xys8OA19B1k9t1jrGmpNfuH5/L0
YuHgjfyZCeDS4UElqEY/teCsZkxO0MAvuLzlpnAF1pTQFYPOtzTZDZFMwLnD
hV8tJDCIe1Vswh6uTPrRVtoooIRBreMP258e8wvo4wbN7FcU9KjFvQmZ8vds
mR3tPHSNCY7plzWX0+1SQ7EfaYM7JmY/hC2nZXOcKwF0Va2jD5GLsSBdREWp
TH1OyJjapuemsHzZKnwsyQScOdmGpZE1ghcHA/49bneUzl4eKFvm8fggJUxe
1HNhnD5rto+yIntuK9zaz9ril6G8N5aHOTqKY6BswwNMCPaSnGp9nsDIOlz1
Z6SguMYxtcaYnuzeyij7HYdKKiZsjmUIUlqPmlVgRzOAhMJIb7Z/LgL1a3iA
v4Q40TkDaLFWjrYY9nviP65rHQ9Drbft3DrhSCJtXshEBr4LZv83R+YbnLV0
aUnfjoPyxZNPjGFyZuQ9NNAum7FtP7HJJB/Ych46B0TBsvuDg4jTkIpQFo1/
pK2QXA6MyhD/9ylBfobOJ7giH1fs2IGAuC5TliisIu2WIqylEmrZKhuT9cWH
+w89pBI69XR7jEQ9NCXDjNEu8NaDOepgWtEcudK4gR/cbPrdWaDgcMYprAO7
zgiSup/bfsotLzDWAYAC4zOFcLYRiQtNzMOEyT06VJ87SMLLqjrvngUB3SB9
sWNb6a0MlZlK0z14ig885o5kWbS2eHA8OX1oQJ+RcZ8kHSIBp/qV34t0QxXj
+AqjIgDIQMYUbVA7ELgnK1Xvd9tFLe66rl+SXJi8VK+DGBBhX4/jxoq257H6
tAznCxz0tbtsdS291CleYXvfQ6OyYaO77ZWYp9P0IsumvS6JZmSRRmK8krI6
FirFQq5Wg2hQTbj1pWXU86f3s3CHcjBDCHGbhxKzQALX45qiE0IWB+lB9As+
i4+QF6702+C9w419I+dqCGjNzh3ZZNonCVhHaoGtf19F6j0lDsbiCBSjODHj
XGkPqW6TZiwmPpuLIa1GTZI3UwDOvhPZOxSQ1tQIFbQv6azo6EXR6q08tb5m
Rg7wMbRBcuvnmZTwhxI3wzWbHil0dL1xDMvmq5VHNgmPTba0P6vFpoB4LeSv
flIVT0tQAYHg/dmRvcdstU9AGU8kQwYZ8kg1bCv26/6kn84DCYGKMxbodZhv
3qUYEVFMjGm/jYKDov2eWW0UZk2GiUWcRWtLuMIqfkVk9nhHm06Hz4vSs2hj
7+oECAz/J2aEhUx+tQTtLF3PGbtgBsK5WhQJSWq2fYqSxPx215OBggsApE8H
gpMPQu+cONUY880oj2aaTW4KdrYGTtZ3X1d/5t5BD0KuT8dtPjhVhVuvObBg
Qe3TYk2j0HnwtqQKlM/ap5UTn+4OYg64X/WnQeBaObII2H3witSEzukA6c8p
bduAYIo+IHm5l42WEF4e9HB4Vs5hMcGTW9kKOUZQSlQa9E867n4aSXC4Ob6y
loy9xXZJW/SatbrNv33Zd/vIggA7AHX4opTBF7YAz1bJeOJAz8MGN97Tbyjx
1HRw2ojjSoZBTmavcEdLn2LdGTL+WZPoWtyiGpiV7EOM3KZ0P9k1aWq6ubhl
PISrSNos2lceW9X8DpgMWwmo0yn5mFFm2mneHt8qNfZOpzp+QQz8yvJYIbqP
ZIAZoz6+ieN4xBFzjuVgvm4Bfy+fH0JYeMLnw4KZ9FQ9sM1h1nV92ixSRE1N
HtXfTYc6GLWjAT3FDEyI3lvV9J3RgVJkMeGTMQLhs9QfGbA/BRuUZ20fov/c
vc6pm5vNVbYhOatuGBu+gpEtYXBpdFFicNM0wGv3sN+UnKKM4EsrSqd/SE79
ddXlmt/66/TELauqWZdpDwiLS/h2BXdPxMhSWCsNe/8e9L6lgIK1V6BAIlm9
CkspaQVOdekIxfg1P0e6Ju9iZ2I/apYmyBfHIZyj2fWc618bpHYWEJprYsXI
s652Ow3dM/c/Bl1/Nq6Jd7nW+agaDHQJ27J6Xa3gsGGgpaUltyWUzY9mHnXY
H/OdNMAUeIbMYhoouSE1Sk8wp0NQEl4bPxup8zGcwqtVJhOEfi3GQgndLqMq
JyQSsDnDG6kWQ0e/iqvyB3479hUyM48GVHvAioYQ0dNcPnHBs7D5r6YdNiDI
1m5gpaK1jrbOLRo9fczWHSXFYS+3s94P2GMlwcBfigcoAlphG5NZGSyy59by
YFtfL3qNVOTy2VXC4VBz9MQJYsPsS6v4GS3uwUqz2FTUcrqqInFIrVGGZbPT
GwFjfkx69Td9CbWbtxzlD6/bg4L4v/9F1vmbAkFiasmfo5XR6+bm47ndF/xd
pKpL94jHtecNNM+ZCDZOhjYQ+R7FdtfWd2LYUPOcjGzdTMU4xcRhBw+UNQY1
YXlo65wPBhpUB611ey4/5w2UiVGiEjqXjP2ZAqA1+TbAYfY6C/ngBx0m/BbT
i1NgsMiwYEUGp1U9kamQ3WtZEkOVmEw6GRJXdcof9KxmBcHp0PfCTObSP02G
VYTotk5TbzgVxoPKr0xKiui7H0ShhWAu4xPetBdrqKCzRNdVQegb7JrC6kuk
T5vADjOE6gWYccYB4gV1vXhmU7laOVK5qphF00KA8bAqjpGHs/TOysgGGpSC
zzypLOMXvqQx3bORZVx0qV96QIu68gZwJUeNPgvm+KDFpDskB8yTqWzQuTef
QB48HSTgB3OXBXBedptXyuoReJqitKbdmIqyfIJ1MsEPoSsF4EVgnJkkRP9G
yWrAvh4p18ArqEPkkyqOHLVN3Ll9Jp/fxbt0WflMT0PT/shCyLHs3Oi3YsHe
ME6598C3yi9etXDJDBqIbZI23uPDjBUFTkmVjXzPs3ja5Ge1grNnWltaRU91
zh1jIo3OT3AZMsmWellofUp1J5H8htJXabUO/nAxF6eiHbLH9PVdQ/pDCLrk
Y+DfuAJa1UeirkNeWB+TxctSYnOoAbSNRAiGmLF5EgFDb3rFx8alnDbkET+g
XW+dkY6L0YUf62MZvjh71VtXrV5NK/vpJqdcaXQ9z7cvZYPQsZHA/Wak4f93
HLJRf2T4owfIwVZnsrCDEPSYMDxQhZ/xmKbLUQQ5xUKsWE4M8k/ZApxelpFZ
ZEfX/2aYavSLlLdtmEf56PvhmvVP8a/DBF6PzlR53v9gXzQGA/2cej1MEMyj
46ghcwIQC8ia0XK4iZ/L0rEIiAnDXRaih9yeSkOHpMwg+A3N4njI0+sYIjj3
XBaA9hW+x+TpSqgJkt0hjcWfXJoH5y6xvgIVboW28y1YpbxcT0hxY+Sbu01p
NLHWCAu2r8vzaYf1aiD1r6cs+Bt1wSsOe2sCOHyIEVT/BrnFZRInKPjeaFOy
p7ePgeMz+6Yb9RnbLWiuBDNagkTc1Xl0+fhZUm2AH7thqJJdBrWrmBCROYw7
Wl88QwzwF0hSdexZfrW+zxe6LuFfZdIs0J9vAEwA77SSZSfRfAFcDeFseLI3
NJdAtrAfx08UQYxLi/yybEoJLVNf1CU/Eeynhsg3BmKmlRZEN7HVdAc7C6rX
L+2u7kCYO5Os1elAtxyWNmtkL//WYyZ9zCXO1A6/bZU9rIfnk/8zPRZH6qV6
oT4qaz3t5O0vy5cS3ISy0QOUme9qBDK3GM4uXKxwEclAfHDOl8H+BzJk+5/e
0XY5jmfgazjsrXwaxbAQGRPc63gnnX5tORHAmi+1qWEckSn7F7GRkzjrSooU
xZKch27oxSjPoTkH8/77nb2X9OxDYTh7HBSz/IthPV7MgxU36mSLCixYRaNT
FQ6wlY4ZkB1qTQV6CMC7n4PrTsiqNcX343GAEzNBe33l/VARqYjOEiYdzAo3
JRHon99h5y/CJqEm4R7r3jnXIsBrnOh32O9oeLsVFTpuV+OkprGUFXbsCd3z
ooxgDFlpnmhv19XvoiNSh+f4gmQMcxB0GW8w/JSVGgHic8A1a9XXktNhqh3r
MHt8YeVF9O1DwsYNV7mJpeqMPo8DeENjnJJKUbbnTAcLC0UZ5KW+FXCM7pCX
FeE6jEaQYOnLPcdl+RaxXs//ukVKrwGIoL7GFpOUsCGXL7kwaZhQItVPIrc5
RtM+j3p2PuDMmfiPsdeU0Lv+7W3D9uJwoyHUpF0JiXnq8nAd3FvMB4Bf/wvi
gvlbSAhkMFmKRkiaj+zqSZRN9vuQFBGluO8Q45oxC+PPhbQ1YMDPuAm0/f68
6pGvopOoN8fIqTgc+rqX3ymwFJsgb5W881pGX8cHGN+ccFJkqagF6N+Txd7q
5E473j6kZr6NmgEDY3MmdJfxoBuArSQUh3uw60YLoF29KU24Ha9/zWqfnDw3
m3wFA8zY1hAAT24g3+3fkrMDVI5RPDPA710jZ9puMZsjQAHBnnc3peJ17Z30
m9GeOLPTT5PwtGCN5anoMFAneRAA4/HVINe2A6me4f1HEOeALUiY8Ofn/0e+
PfpTanry1uNXm0uB3qN7GL0u0rC0XZXZKUsD6+T82nzsKPioG1ln/9wo8tJE
RiyrJrTdIOGK+2NFLBJyLrXy1CVzs4dn7Kw2z22161JVwn/csR8kpapv56nN
SeEYrHG1QMVhMMRmrqCiIAUJr71QmHHVAGSPQyzE2fjJIiTXknsGC29Ws0nP
SuJvyCBBYKXi/eNn7/TBhy1KOb1mSdO0TOMclUH0ibtr6wuh48KAZh9A+RBM
E0RMs5kn2q8UkeOVxbhccZr75UQqFp5TRCJYOERtMdrrhpvRkB8x1TEjogVC
FHEeWdt5zezeWOOHa1mk5+4OXPcoHwKeOJIiVaAE8rOziVOcXFKkgIEg8h7t
/jQQltm3jzCY+A7qA7ujCVbzDIss2hbnokwCHgp2Kq6libLUF+JgpywUdhRE
a7BOX+sTX2e3ojuwpdmf4/bJ95aGg/yhOB6+LSp8V5YRvsHDoY7lOlZHhbDf
bybpJdYyUPGnyMHKu2LWrUqBS+SJoQ8vsdXyJFtRx4NW3BVRSePHfDd0ZNCI
HIB74ny/R01pVTZNhGbmqfyO0939lXnFctSOFYwF4icHXBe8jnuKWLZ1D+5S
kua5Ge9+uMZUh2SeaCA/Lj/T8jhX9Vzk4Il3P1jocdU3sGGPk1qdxghY57fI
oEBoX6yLIT8mxUH5FLhK+5eL4xliAs/K9l8bszbmpu6fCph1AcMRs6JOJ+LU
wnnyijYS3yogiu2qAN9c55nbNqDuxBwiSNApwJkd+HeRuV5IOBBh5sPC25BZ
ualDL/ZqcMFFrwnYMxqcP2YVzmtfwiaktEbRs9X7NB/Q3RvhKibXm7Ium6AG
L4BkeUyes6Ie8jl871URufe3MzStjUABqnuJpJepzX+JqrS+tHD/2+pUKa2f
nQ5xnyWBCCp7uANkAbVDIVbBgQ7M8m7Pht9SGoNbAVnr212OE+ldH+7ohwrl
4EU9iDWtnq2nbnlAQgXLUcSZufumDlrnWSs257PY3mDjZ7rwsD5j+37JOYSt
Vx0joCDkky/e/WyV+CwxmIz2P6WNeB9+0YlbsUwn2+grqTJmZz49M40sX4Zr
s7KGbLwD4pUtysJ2q+fNPeROmx8W/ipV2NZhqo8dshZULIrCg0taEa70tMkx
3SU/dvoyrq4EheyW0jaGuzUndj8uAXvIW17Rs3p6CeVfl+HwYufjeSxsKBTf
2nvQc1szJjdsY4m91xImR1ZlFyLOAFai/Yx3B3Ky7ItlV8dzFt5MaQK2s+aV
TsFh6obADJ8IJPaG0IACxr6O1N8AJ0tJvheOkM12aSkrUeneDQB5srdFpDaq
G/IGMKx6dd832bB+DXIglNvvQEmwus/7t4+qouCLXy1XVWyXEE/EQJbiuVgi
77X8Kbre7wBTjUO4/529JkrHsN610aH82nCBcArxo6ynTzzecCXAO52f/whl
Z+2SH1SjlpC1Pc+eyED+ZQxcxh6iiKtN6FN0sH3agk7OKGK3McgJknrnAXnV
IYYRW2okPHAbPABhgQgTPfK5j7I2Hxq94rzx9GG4GH5izdWq0KAAqB57fSbm
dJIWaU3hghd9mY00Y3M01q6ppKY0IYE4qXXdzWvzWdG2Xk39OwOvH9JlC22w
t2hs2Uh38Sigdbc9Eu14yR89Dq6w0kwRAn1Wup7EKHBB8FGruc50yiCPh2cr
iqbnna3lB0UCDfJxAo1LQ851EVScKu+9jPZAbM0GmovmIzDgusiPj2zwmvCa
svZA+f5jWbdFQIHn1nvxkV7x5TfsT1QN+mpd/ZtMsZrl+I7zFRwgVMgJv1Ok
iETenarJlGODGMHBWgsChNxbHW/aK/iNT57Sn5+3X9NT7HGux+edmdh8RwkI
2DfoGM7TeE1a/y5M56WUKeoDyaZ5bGD6tllMEqHXdFpIA90y6oB27MrbHhLa
8SvYfOwQIpuCQ9h361M/Wx/z1z4mhlsqlhh6iRotBAWMGSYhrTO2c57UpdXm
O2p5tchzsIChVeM5R0qQ6FeB9WfPEBBvm12mc54I5u0JuNU9PLwlAGXtnSrx
lyMna20hf4F46LgX08IBBUU3sDayeAd2RPS2Zc4D4fdbakLIsNJYVcf0jx5z
nTXHRRjZNzJjhYXT1Y2smI3iiwmSOqYECo5429r5SXWcA/zLfk6tNP8776Zb
M837zBUcGC4mXl3hMDjLvemdd31ZV9RXdOP/LLqbi8EPayoYq2XiJdQlrS70
zmnqBdrrHgUdewbCQUxMqyzQJJbQR0w0WQaVr3ApYsz3ISGzbUtFVq8PJwZm
TjRx19ARrjvqeto/+pknX1t7UiWDvOQAUFNvEoJUohKw2970sakxt2BXwgNR
/Kh2croFuLiCS4keC8dD1U91hAM5vH81dsSt9GmbAx9fph3sSV3RB+q2u2QP
y9o0NOxJ6TH3fSNwmH7I6dRRfWDw1kuGFZ9SYb11Bm3loT395TCQKtExf9Ja
lFmj5kHhN4TRzJihQ9E1jh2EI5u4+q8mnIMUDms/xbsLTqKySRfCzoKV6Uqa
uP7wrwqqBS9I+UUlXcja/y1jAYmV4ATY4o6fuLkexTdHv6ZATYZYwaXsXn43
LjlAETzNdieR+7ZJcB6LRovzP2olAg6G57z/kVd/1FkO4eN1DpprkZy/nkKp
2IFdtX610DNTeEK7TXJVDC0twgEJQkeE+CIHwP6mVHuAvUy41U7H+7wLYsP6
Ulwh9FXbgVEGdfKPyQ7ZV4W+QRCJiP6VLvoiZyBEDKA6nmok0vZDgVFlSDvm
gEJuD+qNg7StB/Mcb7NW8g8R2z6iCRjRNeV1JSigfOQS20nW2RG6EJ+9IS08
T57S3uCuDIoJxYuBL6AO1/m+pEWPXR+MC87BMNAv1rppVLzqjAddcfCDVcQo
CEfNBr7f/WMCdk3HDFfsPViMxbOATNlaETFBEKShh4UzBDJSEEfM6VN73595
ugr8240sPlDenVY1ln1hQbRYZr2fLT/bKrKKoNY0qoa9QcnmigkUYcszY6hv
U8Cp397PR5hO8e8qnguXLDcS2DhdK4NYp09C7hrZd2msoUDX9K2OOsDbUl4B
MH7ULOP6BB/AO3cxnUcKTnotfKsagJXv7j1S0od8psj6eNasOWg9gTfWiIiG
WH+OZvCPViyuLhNymnqFHTrIOy6hxa3FQpNkUF7TxdFaT9yTp1h7O3T2pFSs
lN1SwK+5nGf92OdQ+cDIRrLLlfHz3Ybxf6u/Shv9i8Vrq2eTrKHAG0KnobP8
HjJTWSvA7REJaTkzAJCvBz3wA3V+dS90GAZKOCEygmjURDQjGU5Nuc6gosWw
pGNunXvZhttylgwNQTM4y8HVt+KIFWmuwFmu24EycO1W1Tvec0Cq26PT+IU6
VLcZRL9MvgWFle28F+mXqI2tz+RTJh9ywoRqWBgWatrMVwDGBiSHzQ44RYl5
IXuUlFWYJ/YtAs9p4HU904ejAkFeC1RQcZCGIDL29gf41k4EZmjL/2qT0ssB
8E/Dhb9LVEnpsreGnxGWqyrihkD8WTiHGs/+gp7KlsGoC6tuLrBOXPwR/AT4
HkOB/7q0Qug6CUxiP12yuuXP6bD7+skhU240EKol55K2Z1x+GFUTsZa4mJB/
PnIzjsQC4PQPlwRyQFNws6MTbvq3znr3LvUq8GP2+TETpoCEj5WLBsLTZnjF
IB0XkbK0NuAa6GVTXc6JekNepyV1SoaVCY93/uVElfYKikJhmCDXwxDZYVnx
6Axedx79fMipRX7CZGplkQRqdY3dFJeDzJHMb6RtcknsUNfWNtJ5x2sDw0uw
bvFTPA7S6+dOgHaddSDUVGzRuziFV0zUj1NsIn0Lf/nXe1WIvsHObFnSTfAl
Z7k596gBrttGbHgG5hx8GKFpJVMRFxmWVkw7fTQE8i/AsPme0TAlwToGDoUC
MnxQFxDkGl2LE9GaZYoHGKFLnX/BqCgbZYGnni2im/Yj96yULYlo78GzrT+v
+YC90Z+x8GpndlNONdezTij5CXFFfywD8kl5i4yae8N5O7BKDSnYS8UQKg+G
/JsFSOfAx4WnhYLwQ2mNtigu0D5D7rSDK9uhNL6zbkmeLYo4Nr4rNNjK7pOq
72GZ6+OqQv5QdN7Y4wQ+oCghQwQlJBrjbxg/72DHetICVVxxaNcyPGByzoaA
pmemmo+Fo8DKB9T7aZdI1COzh3mH9zRhxlNDYbvccF5/JfOizM3FAY76DOJN
/aq2lgBo/1BRJmcGRX1XbjEuLVyq+h93xlGJiiF4CnVrxctXNvCzRfPmysM0
TrWLOtmwlkLRxh95yrcc1KMHaT7O03MwBwe5UZMays+Pg8WP+TeIYCDAn7fI
0MZClSmiuSI1F4kPBZlEsMl3WMM7n9CdA/sZ57gt5SbY+7na82B2jafo52IO
Wiy0uTBV9kGabYzmYzCswXHKLQ1xd9dOIgdDMVlsVqB4qKm32P6CDLl4TJ4n
bZ7sWjFjN1vrzPMqYjyWg0TTZfOeK9Y9PhXB3q2Tdt9ZwxDrnMHmzdaX8Mhu
+Qt45ZYJlXmxsw+zv/ZJ/X6K07GmqmjkxPGKoTpmx8toPM7aMeFhe2gynXac
/0o/nE9VY2kSkezOk+u53Kp+PCnfI4ziz9iXCYvIdyAtMe2TawxLm4IyAD0v
WiH3EsGD6QDKgmcn+djlFVvePirGWqcAAw2yj+6FWevLl4fYVSSZB7a3P5pC
xfDlFSpLwED3z6Ut4cHiEy4RLXxQgixKTnGJccOszz96YkiPu5tvDkd7D+Gg
OCOroSNI6y8Nu3d6O2HsH/2rpZMKNiFWikXF9I/JmcZVyPScHfGviM3Up2sw
jgct2L9BcucCZkTMNHqNnzjYdWqwsm7HcqUkDocnjzZDJgd4SCQeO9SRHl6g
BLjiuZ0/5KCiG3gykvMMu/yKie9aosa0LR4UD534PRexnu9AVYlmjEk3zv/u
xcr41zzFibbXzCL5643zNf9I/qKN/+iuFuXILNs6Lfb0KS0qNmUoZDWj+lw9
btZfJFtmGKBJr8kvas8G07mwa4Vh34rwbJFPWUZdvxi5az6sD16J4/yhMlfX
mUCLQ67TDFbfsXpQ8oNZbCA3SKiWwuQy5SXtGLrMF2tzqFvAZjAthYit/8F0
oP5IFQSAyAxstTlbgTD10j1MxE12G00MrtOcMWDYqI6SKrqCrZbQ16q1hsep
uf4cvga6CluLdW6VtC4+Oil2Ry0rmVr4hhiahBSoJNKG9OgOVfBlFDVve9MC
iixtLFDV1ym5z4TbjCMnA6dfFjfPnPbantQFOmgTG0laM/HK/pxrdOSy9gpR
2aHXB6rbxV7kguO/+V/DKEUGFl/5eoEvgbMNbfUuwChhPUj9Boc11oXcyLQM
KUGAH/3YWBpa/b2hvooNzYmA3gqGp6W7qxXQNvqi8htG889uKN6Q/eSpFpve
syyufbKIo23MfCsK7icR+X+r7kRzTHEoo4g8bgaltb1byUe5TDcW2ScW3Yje
po8PQENXH8273Fx4Xp6JwPtNERFh5ILemOB1biQkwkJrDcsTAFkmM08n+7ji
zjXXAs3kjUQ1i3bPIF6E2wThHI1J74KeBK+7c9sBSlJrzP5s5OsylPUMIgPF
EPO7YiuCkO5BRKpdAvZU256ntEr5g//UsPEDy5Qxn6QJuqKEaPqsCOrorLn1
g6FcptM4yEW+HQZ3dRK1MmQU4GkIgvLmyWoUBHwJHkhiwWEeIX0k4j7jSWro
A0BWguiNs/SSevPjnFEVwAhmdGYUOraCpkL+tBh0X9ibu+/p9dQ5yf7jO0cN
SGVQREUkVt1j3sZ38E2gTWUBCmzXaGWZGMPoHPpvOQjlmjX2BKVNNpKPgkRH
MmfiYrffCVcphlkdQJHiDBL6cH86jMafuGuPVPBo2lUP7drl0zAtaZ5Qai49
k+jokbStBgTA7pSJDr1FWqAH3/ny2uu3bEjvqywz2Ts4b9hBr+RlVYwYN02J
fKBYSzQLSuj3t5S3rpw7B49nmsoGLGNCDvrx1zAXVK7u/zkU+R5mFZhh5il/
xQQWhLoM1NXo0KDAy6gig+fpumdQfvgZSo6MyZkCryXhyh6NvOLLgW6mEGHF
/MECt6I6yA+TQZS5nQvnoXCOu+jsDNmzrnVM+8/mbLBfH6NLk4aQsvopXNJm
dOkNZPyQIjOpKXEedoQkFu4qvLW/dSfq6zZfV4IZRvMUB00F909QO3J6EEFg
/PwjpHTvBXfVewoV+e4iPxRfEdwgoWf2jRjhJBcxxLqJB81wpONtyajY883e
czMQ42P2HYjbapHeqJjE/5Ob16zHX2IDruqGD5pksbRrNInolXatgqMwgkPD
KO/71Tnr/Rii2piLXShb81xuJBFKLKY0lzWuqkCogGAi30ppp77MSgDR0Cx0
gxdkRb4ghAsfvdrUMePz1KGDYbTYFIsHWEO+Gv5zi2JFxLL4L6+l3f+OG9yX
lSuhOiJsyuEOjX5bXuWZbgqqgeQXCEacn6TXGpXowghaOhrF89oFiOZGjKk/
RNqbPwExOcCrKE1sZBOj6Xck5loFaBm1klBO3avNxHjxmwvXELgtlNQc2+V1
Y0bdtUR0WlObZOgXkuRrvr+FpyZ4P/faZChHfjLgywBeTrCJk0bhupohigMX
zG0Y+kxnYdATJdIjr/VwRdP/Ag49U6dXLx3codMJNDFcww4Zw6ypaFsFf/O4
AdB/kI47Pj1can1zusUx1dpV22Zls0+YbLQWvs9BGq70xnqxeT/9RMaj7tbM
yBvNzPDPe6cYjZ0tzDBh0vIX4oEbMAaciRIEEOBthvS5mCx61r5l9gFzmvkM
4Q54nlhU5z/5ooO1BrqfuTxS+cUgT0MSyVWcRiLj3ZOuD4jPaGwKItJwS1zZ
Ibtqv/WNDZ4h7gwJHt4dOFKD6TwbyTs+IEkMes0lytK6/Iq8Y70Jm1rLzC/D
kBWrUhj5SCkrnlE9+yNwZz6rCzvrnz/1UoVbSuiPLSPXzq1yA8d78Z2u85p0
NLtt/sDdmxHl5IX/sDB5V1DTATz5HvkLBTfw9rtFt0seHFlX3oeQS+SwrrCE
+70iqa6DDOaEVLwSwy0/J9hfYNsuPFFEgAdkHl80A5zW5+mVE+9TJTSxrR50
ShL6iX5jjkjH2+BL4agjg/reIFEOaM+aDh0J22yHmKUBvFiYXWwEWkagaght
ELFYuAtKlrCGZ9B/4zxUwUHtlDwzGIuZTH29dXqgL79LMc9YmvsN7Ydwfh0s
EB2FolHU936CLSkPp0KLM9XfQZeClG/dfA8wjs4W0l8LP99ea5ogJJ4zHDlE
oSlDwm5J9oGHjgrE93FZ3XEy90Z2lppCaHi6QnVEeRcTIqZYajNioaPkxBF9
nZlhKYanJCcyH3bhjLvSOSNLqcKshM9npI/vuye91qPr2430AylwPybI7s7Q
9BI9Syxasg+xcZQ5sv8YbFG8nsTOZHOQKT1KXOuvv2BjlcVIWQcEnsIFkIPE
Qa2wPa8crsqnA6NVOUseC3AvHl2x3vMjoQ+kCy49ELOW1y1RrEUeJ/nz0aQ9
RdI4f5uSDLCeNYMzyz+byRxKGUWStnoqqseJjbNce4AO8P7tN4yI43DvjSEe
tTpE5Lcbw5HW2/rCamNWLRZ/a6sABApCT8HYvakXmiCc55aS7Z48mMIKBdAM
FOqoOaNaSab1uKLTuTGyrKde95FywmSi+us8KOKbo9h4VOvHyUvcFZcyOQ4W
26xp14y1fP+TmkpSyvxuTYc9OAGEWbAeKE/XETMIh1VuUOhY/s0Jj8F5MvXH
ikp4GmEUApoj+L06qJDGOBvX83xZWD+k1638knrgg50OtxUDTSCbfm5svQ8X
aUPcXo6KoQO6wPsTJl2ad/YrmWayARjryd3iC8CG/EtdeZrGrzpkpl3Tvd3C
84w1nit6z7qKnrrSXWTrm/WYsRgR5g+xqf5blDr9FFKvg+JyyU6kFSckh+Ug
ITD5Yb4osi4zyhDVHGUuzFt228IqpawUCqvnoooc5durVQ7T5o/u7O///Q0K
YKG8/KKGkYLQkfHodmzpRlsqjIdWdzv6FNO0ZoYunBNaAN020rL5qDBb8xD/
EVGy9eWjKCQrTW43D8P1NUQ91W9PFnao7ZF5fXnRlxfb9BU1ejpI1P+wJcM5
h7osMNsiFAI/MTxwDbghWd9JOceEMF1io7jhJkmt+SCDa/pFwZ759rglG4Yc
YYcFRC/ifbYPnaqqqn42iNQbRJBh9xK+takq9iRmkobl2bkjNqZc3se6N7ZO
BRyToQym1BLCYmOgOZ5mfJy0bsGtSe4lGAvQ5028XFlxbMbOZok5QEF/PWR8
zxC8q6m0Uvsjminjyd+vXqxJ6s/KRVFf0kKzyN2HCvHXexKC1Foi87MbRfYl
7M3wY0Q/vMZMRNIe4HElhRW9hA0Hrl3QiWSewVfnpSC5hmoP8rfiOvNeRxWm
0qHh3UfShZTqFFVp++tMdDFc3EvzalooEZp69e24nHo2r5oFXQLjY9dT7Z+b
7saW8tANNf5RCoNKYaYaUeGYWq/MoqOQjDFz4gXLrFk/ETfzDYirEii87HmS
G5MzLqD2Fp0PCGYnuIkMvC8OIvFmLDcS6qiS3MrdS9xLd6K+dIh4JUblQnjP
gvDUdVsqFAJ5KwKkoi/TR5sZZH1id3V9ikU+ObarnkNc5f43skOZbZtFYVZO
/tiZCXr6Ip2n8+xyQBsEr/lD3NV1tegkhr65WOYIjhoxgo2AoINipfND323y
2tb+aX4DIH4baoVLtC7ik4TPro7i8BGX4nczGGQBUfGiYhoy8jTbnTSmzTPY
Is3C4pQ5fM8ZDHDOPjC7Ty2TcnDXJSm3alSUXEg5OO7jCoLGX1rKKu1xfK5a
wO8EHF7RM36+aUjOJtbBXEmcnLugDNrONZWNN6kR236d8dIIyvmNPW1w2zMF
txohM5WnjhLkMAcAnjYLk0eg+zQvZmI4DYkBl7HAzPzUfSKai9H2l1y7eM2Y
usZfvP5Mv0NzPURVAVsdUhW9omJdcge7QkfjbK0x1Zc/THoB61Gc9aM9RA/O
5g2utvm/foxuJiznd+rk1YaBolz45h7+r04Ke6PxA00kC9a0pufSqvlsGfMG
gQl55MeKnZQE7WgkIzjoWkWqQ+EpGYPH5PptKGO1tLKJCeXPKTHXx+c/0HwE
rvG2fnNTwviEWP6B+dN+q3xWZIc28tyU6ZwZRVqh92IYaXXkdoU3UL30c0tx
qqZOLCfxZdqO27w/GK1N1Qujb/lMG/exYjc/EfS/kZYsRFcpXUbvtU67F8wQ
XLy66MTcJR/unjvsd2SEFqqQlTmYCxH2UzCkkF8XwEUXbCiJ7lsEmf5ijpRY
S0WNfRpmkfdSl5ms51r6Ga5Si2FPQCcUsOW8JPP0pwKsIOL7yq3IybHhmjhh
QgmkXYMr1f6c8g+BRStLr0hI66r4tjutarNI5RYTaVr89G8EtB/tycmxMoSf
CbVIkg2wbtXrML/UKvTSUj9ULmRWtxxa7EaCahSXKAXWHs7ZaTWWIDNgONrt
xBnIdMkAfKwjSBWJH/FFE2NOz9t8O0xOf8x+gDs1trh6nquaD3t7x6jW+k4t
yKjSG1FU8YkTiEigchHwuOFrBaUQhoQQZfEmErPjMoyaoilZ410wl5p5ritg
//tWl+yjSUFUH4/aovECNJ3el4VMrmZYNIilub38LQwZnnrId4ZwTPD8+RXy
tjcs4PCTlk1iSbuRD4nrqF0u63vUMhijyzdIbqecQ78G22BDTcvglK/msTm/
mwUW1u32wwDUZkpemFdNJsyVAkwLvYeWEZrUYXBwjO0nsxuOCPrJe6XDeaoy
h7kA1auuB2GSM+KZW16JqPQUgg6QkkDk3ILOdr75W8nC+f3sKzXI7422+vf2
/GQD8V7Z5uj07t3RIwISq/v6neAkASdqMzLXzCUOZpEbbroEdeXhIqqLp/kK
zOrddpjfjduRGYIqLvEP7EKj8IHV1FuFMdotODUbByvhnJzP9pX4msxsyQBl
uLRg3xC3yuhRBJwuKQd3BY0npV3mazGcg0/cqNEWydPcUUHaUXpfri1kuTQ3
Z3ihG21+9XPx61NymSm1ZluQ3bcU2tHXGEqYWCkPrQawRQahToDSpdh15HBR
94r50mYUQcriTes4sU7t/m3SNpTgeSks2Hyrit9bPVxXHeyAzvCldLZ9fsJs
2UrfG/GpHl/hrkc7ZKv2ufelozqT363hwn+SYBuGpJL3h/vAjSgZNIA8Ozxl
Us8ACkiukevouhuXuG33rpKM2S82rJxDzOBQf7QXMcUCiTBV3A5zRAQv6Iky
CqtBbETtFM4CmxuwZn6M5Ht8VuUFmZ8h8lJfOekRSI6EqipuBCfnYXIdMUDx
NJ9rQSJY0GHVUe6tU9UtkhjRw/Csh6R9e7PjcRHRZqpK0DfSnMW9R48s+Hj4
N5NnFbaZWR0lULE/3Q3wJ2rP124DfhdMIccKXDsNjrYEJATi5i+C50gQh++L
pXswqgYfSCvMy/3r0KzxuvW78ZFTAYz0gG8yeGcDepdicQ6q+rUM12QUHiDJ
n0PERFw9gqvvPY3y5eCxSYV9cQ8THyhZzyEYybNZlsLqDQtOKXEBRm372AmM
8m7n7KrQkCas8F0FwuhAsXjGrett5zWmStM8ev3CWo7iyBfZ11OAGztnIdqy
V+qv96dKSBI8r1APp6Nn5HeEj4dbx7RyfLdzgqhvLOoHTJCQfLViqAfsSAQC
lhD1IlnJLWciFWXT6qL/yKG1ZWTmf/dbe5bi9E9Up+o4VyDCjzdksyhxuiIu
LPvEF2r+0mqGrceb8McfQ2j1g7z8B++a18cATQxxBUgg/Ml2ch/DSdWpu8LS
9dLOnrDVXq0GTWr6Fmos0hk/P/LWkE46lUxsgXZc5+G49/lLEqFMhxcBbXuP
eGHhNVSCIjQDUmyyuXpOqOMv2yToeeni3Q/IhUrEdHHP8o5jfToiXtHQs/BY
fZSiA5SV2a1NSefU3++E7ZH9zF+3TsZEVvWsOgiMmkHDUGtbs5LX5VmRU4Or
UgwrQdym5p2G1rVmkDGEHFPP8djWEmQMpUR44VXuOYUhDHebCsKCULrYgiNk
PCy2ZZlP98IEsQ0M9IUZnMppEfAyeQbW7RATHZRvGQOHn8WnaB09U/TIj/7C
zFInqKo5FMCmRh/V1U/MYc/2RFrzMaeLguagtEBILlVAbyYiCQbu9WWiuAOV
HQbfCWIoJQ6P6ksVWSsi5MCqB0pMUA6nTNVaLCSpV75R+yBCWx0C/JMoFUDi
2PY3ypk/0Pq2nElE6Kx7wvaxwz7L8cD1PKULq6uwV4XcImBylR6G6aH9nBnh
pmoQ4AQjik3tnRQz6BlZAa905kcy3cx2KkmHdnSvPkjnBvMsWE8hNqdqO3w8
2h3xtAUHV/qwg6Qy0YbyRRbaxVva7GYigPpq0B8kdH/bQZ5DDYf2oNnTsopw
h5Ze9YYlPXAi6lIRkNm/HeZxvttxCx2AR8p15rYjximnNzZ5VY+D0xmRcc/H
59ORyt9//PO9kGtLp6IGWXwT19Qom8Eiu85H5DJmtx2xVPjOIv03HIvD+BtQ
7hr0D6+MQDPhtt0VUHuq22fwG/W8n0GnwAV9FQqkL+5uIGjvm51lpvO5XHcZ
7W23sGJQfWBNfLy15H3q/RzafFIg/mRefvZdB9ipeenQ6hXeZTErY1kLrifY
dDohhx0IFSIuAfafNS2Lau0OYR1XV7D+Vgovgj2AVGxdwfRRuiDKJG3UbUVL
VKa28LyCoGJiorUe2lsFATk6Esh1OfrL9aaZfJ5Id5fBoD1Ha/g412K12zBJ
LLQURzD+spoDV55k7bNY/p+jHmFFYBt3ypaCsII8gsJmIwumgzwxGfmR7j0T
7rNPYZl+qteZFHQPMODze2numZOZK7l2HcnKARLLgrnXjW699dcRIwA9n1YX
WayLU1BN9tMLRMYCyhQREdlpoIgQDCYCU5/5rNiiNK2Drfy/KX5E9VoKgKwX
/rKxxlq+TjTnDN9WJaEBKQjbgDzYt+V8tFja7sZLlZTy06G+GOm1k33hSDuz
HrVNQAeX5901JcFQlfkikz3ev5/6uQF8bsxPmxrSiyNKKm5Ppev3w9Fjn4C4
7oTV1NSS83mItR/B25LZuiwM2TeJ02Ho+g4oHAcRradFIsOYIbnVa0EN9CMD
+odVKe81JC6QSedqsFlFudHOeX9tXapAehznpWeGWEnPQ/olpXnrgyZxDxtT
P6rnDawTIC8l6RGmw5kgc/cIHkvWCigNQG2ZufRhfzc9YazF6Xiu1GG8T8rd
cSNMwq+e69F32/Zq3Er8uFZHx6howxhWhtG+yJNN2dMjKbO/MDKVOGEknehI
if3PzFmQ4+A0fBcEjsyk9Iw4OirpmdQIAtMQ81KhHu2i6B6XZ6iA42fH2eQP
g08M7+UkCwgToJWred3EeWJ4PY35lunBtpsDJjLehWBzr860OccIyPc9Ne3A
Rtgo5HdNtAX6t/e3zfPkRt2WnvLzUovqyYyVdc9fdI7rU62w/14AMZp3QjSu
gCx3SgoJH6yrVzwhhi1C+ldC1NdPceqLPAosxfGNlUT3y3Nupl0yGwQ2Sq2X
7WNNQOL1QXoIVZVq0TW8KyNLbraag6n9qVci99sMV8F/kXjMoJ23ygww55zP
Zrvi2kCuITXMSes5G15gs40OwpEDFQuBr5+Gkp+K38BO+B2afboPZjuCVbNx
wss5BNlEZwLVc09srHQQvMRukOlgqIkpAy+aWxpsj4f3K1+asJOzrKNWo+Ly
aNaQ5aoL5SLMwDxkoyhMDG79oe/Kt+MXGKgw7HJWVg+ZKVNuHLpRuBl82iPV
EK5snIbOqyTAywuJIHaBxa0MJhMkPewDUHkbL6DwvHNj5pqvW9krypsRg+qz
2Wtn4+hLJoRTFD3AYLTy/WAm14sizuESTPmA4KJfCx4er25A+b0k2+yD1UWd
m6ZZB94XMI51d4RHxWlxXRFWA8qvVAMutJcThQtbZ2jkM8gsLM/bv4noV17h
4nzGwIe0Ywcw3GnGk7mrP5hmezivvNLc6UqS/QfEvKloG/xtaErHBWWVC9iX
o5lEa64zkaaGwD8JPMes9ZXL7duEp4c+EJaKeiCpBbUCZtWCZQgAgdvozqNT
5h7+UwRpdfii9YUi5i8DAjAzKbWEOCQEzJX5RS927Fjj2X3l24KLqJ5q0iuP
MJfduPRmP4nDo2CcSrV7757tarLRSRz6ujr2WAMf6+gdv3ZLQd02HL/xTEsZ
+IRUzFJm7ZO0p4dM92LmXJSMKEEXZiqcjzfWmqq0T6TCnpqlG7pVyIm4ONEh
B5MtxXNjq4hjtj5IGT8h4rPJ3yTk3YpT7oSDSF2QWVMs3YhB9EHC83GC3hwq
uz+40stTFDQS496NT+0wjpb5lhYp5An346aATiIwsF34i/0bt52eH2slJs/6
fpGPhaOj/oL9f+XQmE2m/YvbJ+nKqNmIPXWB7qA+E9fTTSFyIw0pmTxQ6O2M
R9G7OfK3Wx+KLZ2KZ77w46b5V5zUGVvJoaDOk+m2/08C4oSl0GI2bm058AJq
nH75idY2x0XouLwZ7wL3RVY1dklddDE5lGkES/WnVe4ku68dqFgT+1HKFg0z
1MrCntM5/XuCLXf4oriljlEyBO0o2+ho2diB0qa8i+PF8nZLIJMtIvEQs8ml
SZ5k3/T6JFW4WcanzDFMfmiFLBDYoR2V034wCfWFmvCya7W/X4jPLonoosCL
Ko6ogAOBdqSUIAqfKTOQkXsIrcfLKgy50m7qD8ez97QGtJKZQoajKszvmdHg
mDgomUB43yNInt03JbMr5qNpZus5MKbvDuJ/B6HnCyIlswcqfm+17N4BrAAR
vzVbABNPAwfYyvj0OoHwq3lEZXCPkPjKEW+gd/cyOSLjXbQCXNAs7DqnBqhK
hIO6ASCAVgbYZecQJRtE8vD/xgo7MBhfUs/2utassXVH9Gfcqg+g/zTZiWoQ
K4wbks3LypkhrK6fGqxYX52NbMvWefDVjUIJNSEdgR8mPnYkEBj5Fs5iO1kW
5TJnC3tofu507IxWlmF82t4l0ULHpwVzOwv/qF/Q6j77qWLDrZ/2KcdgKrOo
Koa6rLMmXCAJxOopTDol/zSDQiD6GY1PXnSbU3sTZ3/t4LsJm7wq6F/xqFYo
OpjOywzXcVQZA4qnYWQxWUdCDyyT9b5o4tOzdAeKnMxxAnfQiogr9riEPouM
UuhaBhrLhmtEURP0fW3DhLf0a10lgMdl4/R6MHxhjY0jVnxOGPeHhk9Co5bA
z0DksayJGgsnzjcM2UhH9dQVY+h1RzS50Wof0WPbz4TrvyLDYp1sgFCYVOtA
NZvllClVwqG1hA8HaIJEAa/BnX8TawF4PQHDhcIMxJBdQ0sFM0oPVPz+TB96
i9WeoI5oXCijBsuOX6QQeW8dvDcc/Q4Gh/N8QKzlBgsSrC11GTCinC/oZlXF
S/FenKOjhinQCmTB2CUim5eMe13c6sD+EqBOcAE2Qvtg3fYXsOI6sJPfh1pp
4834qNYN5cmb6BTxyrRjE9wNjNNULKZ1yUylAqVY8IEbf+uMTXBjNMap9VyM
STcSQiSlU+jXneKkVW/blkFG6oNku7bjiRmirze2lqV81iOSCOLpXEeB9ssU
BV6FXda+c+5XogyIOcxIc97DhXL70hxWFCCg72ACRwZRveXMWsJygUCJ90gB
QndtAi/GYhWC42cd391b6FXIS2ya5AmY6I7F6WUJGvswQU7SKh7I/xgN+VN7
g2DsHykZaxhKxvdRp1UGyRdG8ucsZXHai3Y47x9naV00X6bVcb+AFkQ21/8s
SUkNXYUF76QnRWZwI76/p9RxJoW9BVFccJziTA3kDelbIRzM+uTRGnZv4/JS
dEqEmED411+qmWkbq5bIdKfWUyPhoPfRTqkZJWdwahcomDkuxbi1fZBo/PCB
Ge655FYAl+sMhdpFqhFrK2ETaNDquJn8cyHhEUMk47sKoBcETjSA4pC4CewZ
w+QPCWbY2oAsyRY8remrXmTdU5qAOr33KCLxkyAwdKyfYYBmjlbGQAb7xCDb
zZNw8zikeFqTubNa2TGBKeFAWn1lrhdLdbayAOoUCuBm/SuF8gURGSlS6++B
xgGdzBTB61+YUVpv8oxZXvrCNCMJF84zYY3q0kvGiStm+vRRjFjtwcml1fCA
LGBU0vGoJupI8gQlGJ75MB5JUIF83k1ndbus9w4Ipn3HE7vT2CTyooeQLdHG
iEHii1HrIGbOFtcvY1MTgoeb3K0NkHwg8Ne95JOA/05xcDl4AE83WD4vMkFA
31f1CBULFstHh0yoRU6RMxTjHDJzENfvjqg8EXUTg4ZFC/6bk0eGlrMvVyQT
0P2GBIgOKMJPt1i3mJjhHNosydv0Rs1gN7hR77xJRQfHXeyMrCjfwLC/KWzD
/MDLwZOighNSExxzNoJ3VZmfUhh42MzQrMBmgJiIf7wzhZv4loCUdR0IY1nB
Aw5eRfiyg80P3kMdDcOo+LEHJsDpHpPQQ/kRSyAiHfPwdBIoXP/pk/IWTXvC
xo57mJnZg3dr8x+QudN1Y9hcXS0hw6EdVfCiiCYk+2bscw7xQMuTgZEy1BTZ
d5o5tATNQ42JTmRNfMPwlyXlBOgJufQY0gFMQAoEMBgxhiwS0lilJ9HmIDnr
woLQS06F9uerX4SDXhSycQ6Hotthjib9h2Gn3rEfSg/8sYTp1xMH6xaPQRtd
rJDxfd66AEUYCUivPvXVguPxlK6i6/a+UNlqPYuKOfcOGL9Fuh2imjyHpY1N
X8B5pjmwFbtc0qIH1opcuIqECLt83eh+Ll65iS8gQAi2YivVfudmSGsBNKGK
WPFaKepD9qON3DJyg2Pt635Vu0XSopxA18LQkmYJcqSlgLYPAXIVqECUByLW
qe/iG+83OyKI1byWG7bvKmJvRa0ow6FgwBMe+MtNVjXJ3r2KT5mQG91elpvF
7Z9pvTsQm9Yswc/PWpWvoNFm7vtm2Wy64jpFG7SbvwEfWey7kTgUy7bm29bP
a0/0oGCHozqKMjm9uok/hphTERKhXWmP68bI3aYryCAa0JawMdu7cGr13EO6
MPvh+9P6wiZJyPfkg82jGGBJlQZIh29D98Hhx5D6wF6JMGubjloqoW6ovNUb
h46x06ipGTPLWY27+vAj/th3QXwdRkEhKCvvyjAIRRJjHSGZ1I8NYCA7B5C7
JTXh28/H2xRRfq1bvR8xamaKZc83qG5m4LbHtRZ3uc6ekjnOQ+4sqzzLGyl3
NikC/8GV3VL7PPFzWOG1gpT2w3a9N/o1bQe0KGzlSEyGXINww5k47iNckX55
iUAcQYe+Y90aBmwvYFFBoqZsKBzW4QGajtc5ivOChdbwMSMFox+oaiAojDSH
Tz++KohBFGuuDNuI8vEDyTmczrf8hkOhJgRdr6QGB4xfcR/ndFIPYHjZzX7R
pbPQaZmaKhlNZ1mhWPcTtL3C46kZojF5hVTcnJz/UxCJSOjJpKuAVCSFxnR6
gc90Oza7vjC0BICMDSf3O5FFkuF43vKmDiMkgpJMbdg1shXKP9HR1WPxZKzX
33bZHFCkVsMrPuB5xBxb3s9R1aiX7u4fMpn0GR2J2hxqpKT11jqgFUCK8AxC
HS5yVFR7oLhUPHhv07FYzMHlWwqqJLoZsGhHjNY8Zx9qxZeI8aRQal58p3Qz
Fb4/u6EH8bSVvNAUpa8+VutHU/oq0mMkcM4WQQ09AUVCkgGz9sJP5cl51BOT
8Ypld+JvTB8TqMoY9vkh2fm5c7et5ZrikYeuk/sLCEeRX6sb0SSvJEG/XbEO
Af9kKlUuVYVkd0RXNg699N8D7jzV7x6ygyX5pAaLxQWl6UPVKXFlkq4mp2pc
QhE/xmpJ+q6pOw9yIXmDqGLa9cKekxFQktl5wolqS82xJMLOZI2fM+m/CqN3
WW0K1fOaA06YXeuYQy4ImqGQxdu0PDxbpdPDyJpmwaOS1fsB724hxf74qoFJ
GZkOrxaI3IRm8HVV9PyUEMNApC+sNIjtnoxL611/SN9T9xOXHsgnqBlX3D/O
7MwQz84lU0j1/ngBDbMD0Pt7ac8OJ+HPqqZuAx9/n0JkCh81XAeGzw/xVh9o
wZ0s954dgFhaXQcwog6xPer1l1rdyFFXyg8k+Fx6XfKVAhw4oxTlgfGW7sSN
ZBvanQ4OnBB25QBZAsZfJ2FeeLDnuPtm1Sc77JQ5gMmpX6u0RsvBCb3pYsfO
j2kz2a3XwA03N1iwAL73yNGaB7iZRb7E28vJMr2i5Ly8M/FQ/g4iCMHy6MU5
wf3dJZky1vUeGaWXZxlUNbcnrOgoB7WzyBk/YyULnIO7rGs3areKOvE1giXn
a8djt5eZzaE2M0Mx/VfywEC6Xa92O2FatwzcKypdKhbiVKJdmhgMFaeScElZ
IbAV4ccSk4Bygita9C2+Eta65iNTEJDJQUmZqDc5d96TAMmosZalqsoYPPWS
Cri6vmNUi9Qjh9t+YVQRjuBWQ7HXWxKHuccb9VFF/ll3vyLkn2EklYRCgCb/
79o6GIGL/7sL8BUZIP10mErmZhn1TWynJyAvyeLM7xIh4OB7B6cjsVd9HVcC
Yfvmne44gnJCgivFFFPAJ5vhGbOFFSvV3AlckVKdSzml79meJmfB/9PKemc5
r7qHNmTHu2Kg7KLxCSx43jsqoMmdML6ssJd6dvUUAQv0L3QBTR0UgfI4ajPR
pgh+HgBuavL/J5v2blp2iDr2UP3TcZCwTu+FwJ8Zqa2Fm+xfZz+CDe0Xnkqm
mDUB8KkWKxKArma5eVwEnVPk97JQV15MoVN1o/NjsGAKHwOEMDxGUaRss8ZM
fWMmzwza1tmxjGSZ+23IZCViAUfQ06mJrIJEEEIdR55P6aNMyQuoEPRS8X5d
Zh/rbl8zvw3OWDSVkgRarEp+UqDk3vfT5aDUpESjrS1elQ0Elhl5y+Q27wj7
4VvRAj6/vXhJfca6z/+KAPh8bvOf27k82IeXy8nS3tqtpD5f2xPbeIYT9wZ7
sXGXpVra1bKhy3EmHaWW6G2vzERGpZ3IyuKcs+6AH3wlEUFu0mWeDlvJKWfg
/BlVb2n8zoMLBMpFCrLdnRQ1EyPtG5XDsbYMxfWOcLe44MQCMcu2RvoA9RGk
NWf4+1P/wHC8wqCmrjjvK7IBtgLMcwTbwiR1xun5Q+TsL3yxKAbeVX5e7296
zo1FKLxCt/A1B5H7jt03xt+7mQeu2SbVOvJu/9Fb2E01OPEdtbWtoG3QYRh2
xW26Xu+ygqE7csS1RUGIMbmct37FPL3hXcKUvD6XUhp6TzEp8cpujxFPOrZD
vFRcXW1HqJunt53NPmTTsJ3MfENgt21D9JfgVrqprAwSGaorhBsUoyX33CHw
K8f879leYRdBq+Ccjx8c7KQt43dtomypRQXB05MREKmI6qo4wKmkTZOex/T3
c/pwyAQK8Ptn2SkpA1x6GRFP8AUb9YsaCWYBfxx5eIiVX91jaGZaOng1PZM5
c9zBMsvqlUW1kO8E/4/OriASt4ITvxBuXWCh1jvpBshq2SgH7/DNt4swazjG
dOWwGq7wU8r4c1HfLtR583JlG5IDSy791oWs2j715J6h8IlLqXkLWWbsXoTe
yvZt6XiuR0wNtHe+wIg7BcwiqHqscPteE9egwcm68trOaFgXu3PZIVq2qZMO
5TC9myt0824G16EqBQ5XIqq85kBN0fIkfC6fTfLvnLAdhlzDOuytnej953pP
ZoZx3CoPQY0P953XMwc82U30AsaySpody1z7EoO1cdqlWXuABCThCvALrhzo
SaP5LIbzJQn5iZQMCyk7/SjIB3Fjy6Wm2vvtf5b11a6X6DDZ4YW9tlMJ8NmZ
i4tedO/7kbl3QynMIvktm6bcD9ISDxt7ooNaF6iQp26mMwC+k+M8vyf05cPP
BPuAbbIz+6lZZflyq7A9HujO77ss2cbTnDNbamn61it3UUDnh18OcdisJdE7
+G7+QAp73NVlXG6Zo94FBLDK0gg94/Qnp/qgLeoubb32yYgJnZEdXv4ISHVE
T0EfZBvYL++MPKWKre2WeGZWeIuPebBRn2UdAxwF7lQnlh5C7Ja4e6VkWuKx
L8WixX/JVNCck91W5zqHJ9tCdrRkBMQxpxXUB6iFKkusszUP3vKgmBSTd3cJ
HuqtrtqSQ/cJPIGcc3SMv6F8qnOZI+Wk8ObpfDM3/vEwfulr2uckAb4yCU7b
3JdUkvD1TXyJ8uoFOKowbbCmfIDyZpAPWEi/2cf6S5fQHdRZXUrUWb878RfP
PSFue38D2AoXnrj0ty3DSWohZUB0KBcTdRj2/F2EaoxR/YrGZkln5YgyxPPG
QV/9PFKC3Iik7Kt4Jmr8acpT5pozyYA48EH6SL8JIkK0NLpOEgjDBZlNKh7R
/AffHfLtdasVEJmxS95ve2tHVjXBNURQV+YzZglN4w9n69fby+JcRXFzlXPV
NKLCbgsPJCrmRrpqXf/B4psMQX9+BbtIucw3QeXsxLGt8Y/FzNoMMRPRoFde
xDHnxNw0v0G5T7dQ+t7UN01hpWKoXzB4HScRFxnCnLFj+2IP+ihDhDCytsCf
NY9SUCDmrqRb1YbtSEEavp5RlSJ/qOnWiwFHqWltGjTflgzuLtglSofBgs0U
UuJHnOsdLgSY2znwP2KnViYuJ4NZdB9q7ES58JxPDxF2h8koIoUNQ6/ffUGp
15Ex0uU9bJ+rjw6/oBH3jsH1yIocBQmNa7rDiJ9dr5fQnREeFo1I1Xzy9i2e
V3EF18G3QPO3sbHQuJggRs3TOZ7FtjeHtGKRMB4HSDMZWpsKr8V+Iyx1zZM6
Vwbn7+jyIftl4xcn16DOQvZCoDiuyzw8UOey15mZa02V3su6gng9uLoKMSFZ
AUSusvy0eR54zkhztPEZXcCNP8Wkm+S6u1UsvRrhfbW6HoQBAv0U0QY8Sy0p
JyuMSZ0Fz4a/vN+DEuTiUc6ReChbUGbDI7KCrAJtjMPeFPApDoScp1g9LOc1
JEd5gq/qq02wHsoG672hlVBHx8BYEjOB1mn4Zsx05AOnGDHrzHyrZFACMaFQ
RXXRZx3pWskCduZuGXefo2rrahAprh9g0SFpbA3AzWn85AHTmUEDJk9ZGK4t
fOFlKA4hBn1hktvyXZF117KT7ACbCJ3il6lvQykrgfRedICp9j5ryv878vYE
XbQsBKWUOnLeQO+72rwUv4Bid1hHe4uJ0zuTmsZoaD1OZtG1Zqc4+5RgHUi1
6ulwcWA7abkflHH6R7v8ByC8277vhqTITIVDPqfDDW/qNlg1thkE2Oo2Ia3D
bnvkyyPimjIk05K7SecCZJrA+X5d6MsNc6Y/UCrLQV9iniKcKu8/2TtGz+nR
UkP5TUCOaBxJofIUU53emSxiH4OWibpsnA0NkWcumF3eVOBy9v68mcniM6Rj
aAwvZr6GCCRZAaPzwQ7fpbwiI2qcee0LW7hXG+5aSJ+hRsHl2ah9gJbHNz22
jd5bn2B/lJKAjtNktlv3wBS+5zsSLDyK9D6pUMbOcXKG9K0KMgugF2F22zeu
ciZNcgP6fyTCmPWbioOQNGAfOxuPLK85RtPwQo9yYyhfB6N6NTJIQWJTY7ep
KZTtbXq2ahiX9vd5Q0Hn/+7NUpo0gK+rfvdwwNRKWxHzNlzI1ayv/5aL5jsP
N5GzE/1E6NVb4CuWJI1KNKhjUMf8g5ueHyMQRGm1l07jqyPFbhrbAgT5YiuU
RenmAxgmuyJe9CMH+lmrj9uUkXv8orb+gXQNpZk2KmyCrp5mCPJINTHulATH
YEvrVIvmKCA9SLN8gGxAYoBx8s6mMVvwPnDtWF5ULcVed68Le3gYMPO9sb0I
kA38dI0tHtpYBtRMB5izU9k20WJJGcGG9cxWB9Z2QKVbuJCyLizBrH2BBEeY
F4ARP9E68KGMtHdWjO1GWJrO8L7d/CL/e8I9/ghdd5O5wT7xkOWqMZ0Evqyv
7Eyk19zHYPShZWwQRbG8UYZ1I4z9s+J+F6wZyEF//i1eyRs1sW4RRamPwlUB
lkYnOID8oUx2a2IokR1HCvks+NPPgFVtP+4F1CpTovNiHfbXWBvJTn3A8Jfq
MRUwKo1qP3isQ/yJ85cKVko+H9NwAYWjYV9FMAbJhM8BZzGNSVbJ9bmkyFxS
M/F4Sg64mXPYtYGv/XIUU0XqcswSaCUrx5i1thREg3qaiIU6rlxU/GWac6EE
7si9yKOIJy10in2+3eNhC575hDymlu8vfjkLdmXf62JRbYxj+U06iNVJA1qk
DNuUqkq1X9qe2kDCbV8yy1DVIeB/jRrruwGZVVtDiK1p6SdyRxBO7Otlocby
NaTJHp1cVKavZ9vHJ2pbGgTJ9YxvcAbKQaFHBTaL2eT1vp7295UkZtyWh9cM
IoP9O74Zp6jVdfx9I0MhkQcmGE3x+aBq4DYu2++kU6tFPJNCzcLrP0xV93Yk
PjOAA5TOnAYkNM/YQVV33kNAInZPHqfoXwDcxawOlri5QDQ4N/7nOX4KZQwk
nWAImhCcS7We0uXywDwJ1WwN1ZfSV8pc+EIxnv+KM5IOvRWzdpMM0g0FtL7q
bgwgzHPryS6YBsZgxIyoap094IpBeWrzEFbOSE06ZY8L3fddX29kJv0rDsXn
Q4A+0IYvVV6sYUut+vcm4D/kSXXLTXH/x8nMz6wCJCPd+eK95CJ+zAQlTxL3
pDicELaPRfuJtww5Y3/9aAaiCNSZ06viS78oOv1UiQOX6bSeyyMn4xXzV9cT
yUerpZM/00TJ4zpxRxQ330Bl/2e25sbodAZ3v2R74g8PnICUkMOOtt2InoiE
Hx9ubaoX7GnU86Z75Qi7qo4EHD3dUG0FJ5X9qNCya6W1YkV1axOh+DkQBeKC
Ijk2zzygQfr/t9qtrpBOeZBZMMTAw/tAmNGNYGHc7u1liTxkBK3n3wFmsblM
CDManFv493Xy6LgUcAhqWoWKT5HzkTqHCqRfhdE0LceT9aPFzfj7gLvP4R5f
4TH0SOQgqiegvPwg4ONNyyq0PXNEVa4e4irjc1oHYmoCER3ldJMLAZZ2SLVB
fog5EJbr8C98YcRKWgW5PFSv6Sp0cNSmPKxc6G6MFUWdcajraWdWNcQomsAy
xssMS3/43NS6limR+vQY68KZ51Cnk07URIb1A+zcW1RsrvIF0PDOI/Yav/DZ
TLzzIuBposeEsTDTGI+kMxBTccPkvDnaykJ3ofeOHKfsEm0K+8XPv3LKlMgz
KNhCf0oE/H7eHTTJll2ov9M73a1Q0u0EZY9M0RmRWcZmrbNjR76+F8joK8Tq
Z7r4kVIffy3B8qIjYnfGjG4gYf4mF+Vsg+PMo7IKn3vzJc5XwJXUKhrBzoM/
iODWBi0MH9gxaqVlawpPoNYvpATv7Nzc+NIr782S+wXtMZyAWoGilFlyC7ja
VRcwC2qSfqJQDlQckGCMwnf0kgjSyVoyH1uBgGjhVEts8K4gZH1eZQ7DYw4k
NOYJCnWQNyr/sBZpDMCB1v8Wsfj/rfK9xzrSw5cAMLxBS8eN06dfKtV92Mwo
LasMWRhF7QYH1s5pEmn+1sF4ogwpv3V2Yj10iazYWNtcWezMQlF5zb8eTdyZ
HbVWESqVqagHOkDLDBgTgprZnaNHS6Knlm0wRfaN8nFyMdDiJVJnbglyU1gS
5LlnaiLPzWE/0Wnk2FaEjZlObZ5MElETAdKi+B/Kt5pMdhz5HiBzOxWtmdfL
iKXk3hsDJp6IfWZfFR1roKW5hsCNc0RyzarxirB6AdKMeImURgrizfyNSC2/
jOIu8/ABTpY+dKRqQ2fr5kVexMgeeFIl+mCHVZmhYrtsHo1CEYaBgIxCGcLS
Td6EByWDmK2zDxFuGfCuoFqWQoAfpmmf5D8QTEKMyd5v13n2RVo837ATQNoX
f0YtsQ4huCMsbGYEASq8Ux11mAPoy4+p6/1BRUCEQra2jhmU6PYcTQPbeMhG
QDwiTUVVJUoG9uWd7r2iUdqBVHjYxrMpZZmzcQdSZXkbF7C8i5ENUwmnQXXP
dDbtoyMbOLzLSRK9+uLHFESa1HGW1hNxbmZhc/E5qcEoGAAJ1+y+r8CHI/N4
XziwAUF2tIBqPY3n/hLltQaZyejdf64XBBbRuwNvhXnCtMZGF5JsejytRxVx
qvqP2qW2Rc/3XIKXez2cnm3LiYoCLPJQBHV7xtK2Un47X69BEbhq1fgHlCH6
CBoCraVp0Qk9UTygk7+4sEAq3lmzZWgLf95Wf6ZijgShbhFhWBUBzqtQLTsr
H404h/fBBH6PIGXK8emlaBYgdqod7Ahj3oU7F9OciwYNQMjELSHWLloy2tzg
dk37wbs0KJ4z++IkWjeRWg4h/6LLehtVyjWyPLFymNoQH5YPdqdx8joXsTP2
vRCejzu9c5XkR1tCepeXvGi167wIMVVqrTnBjV92ASA3YfcDlXE9UbgSmB+U
a8Kp4dCzWE5J1lo37xoz7/ePMldoUQ03lR1KCf8mhfpiI7DvtsxZwfCFtmXR
hGT22frcqvKyPEErYkS31TMVvyz3CKIiizIWz58uWMCy3ztKW799PNSO74cD
FU1j10jHvCcMG+0C43JMwI5/uqCtHgBveqCEWy9v8UO64zuB8UfFu86ereb4
eS38GIwT/mwYCgS1MPqJriChPArbnsfjMq88CIM9QGS/O36Cigqf2vRMm25f
FYUlaLksxO2ZNHayiRxvAOzb1AdxvMBzy4l/y3psjDIQapxSw6MK4Oii0Cxf
ASDZ60B8wjRiMiLu/qDqJ86viTx8eeWdxv8FYv7oFcSTulfJqPCjWsvlz2Lb
44n9jOpnfn2I8P4G0RvrIis9Vb0fniakDgQutPRhMeAjGnmutRp2FiTT6yNH
Jaw5ZmSN4OIil7bXz357jclO9OZoYI07ftjrDL2g0IrffHHHEhY2FKA1zaV/
0loYmO5YpK0mQAxhwnjRRmz9CGFhcJtNz/sb+uZDPvJtLaSt487mSxpyxYaS
xOzYSsbwdnLqebJYNkiQr1UacPPWAmjaViY0jMoRsmoNorHel4bGDEYRRLGh
ESHck6zpXO1ZxQp9WBItrUKDopg1oPOcnMFV2QWn27bZqOmYO4PPifJPDt9q
f2o61bmKw1QCpbO8I4D60T08Q+xF8jJZ7gAGGYHzr0MbKBECm57MhK1m4Xwn
tpimOvdcNq+n2Vz3ggmWoUZGcaUMR9wE9DCm1xm3B8A9k0Tac6KSq+gQuyMx
WOoLGz6D+GljaOx6Aq0Lo1z1BsNY+H4/7nPMTyjRPLPvFtDjuurzrXi7weYc
PjRt0WUGP8GOCq0fPincTEhJKfQKgVFrLEYR4jXxSCBH5kF/JFj93ab9tgwT
4gH7wsf67BVKOzwHA6s9CB8mngY3fXAUUALm9Ommg9AvAS8HX0EuPYqieUSM
gezQT1mleJZPoo0Gp0jgrj7L9HtMmh49G1+s2gPvQIAu5t/Rk0Tm6Jf9Lw+a
6GRS7btWp5XgY56tNjXsCnyq8T7QKvhUofurzTyP4l3UUobiifEVC6TFFqGU
7SDOagwnZZeDNLbVc2r8l7soFhjO0LU8FN+8ZL/Sp9n0Jz5yg1CE3nqgwTR6
DJ0kuuslRPWRaiChWQFun6EE4yx9jj9Im+xsSYgPIPXeXJr68fqJSv6h0FSv
/QQFW1UrLMiiMmajhPtNFB4sNTmaakV2lvMCLAx1gpuhvDur1PkjiR4cVGE+
CptHoOwYULNKYHwNWLMF+O7d2ibOGKPTAwn72M6qm3G4uLfLSc824aiikpUr
kmHcOVkMBgxrvaCSH5zgyqwwI+tOcxXWwbRyDXcdgJ8s25orAcYNSf5WTJ4G
pYo24RfLsafBXlDjUHvJb+LYL42vQNGXOyIrns37KeyfA2A8b0N/rCBgoRZs
BYrWGZ62AXBftV77IsHBaw2BlLoLg2K/KClbbaZTNGmg6xYdgfsP1sla11nb
oD4xGi97I2hyA8cQNRdKssJP3UesY1FlD/bMl4YOUKXqpxo+EZH8R4el58Io
SATE3VKIlG24Xjk1O2U+OneluL+Qok9oVIHBO0Ews+DWvSi8e8IiXV2jDlp1
PzFiFdQK2cuV0kKKfX4PRJbj16N8qEDGkR/BXnEUQBcUWWIZ2yvGnYTwo9A0
9ivneInQodTa5jcxYYyVlghzAWZaQyc8cXviAzwwF/LL0pkUgYGay1DH4EZf
RTIxWMPvCCF546BxKCI+TOGQKurP/T6fwSHKsZ88JoU9PtN8zAnc+5XgJvEC
jioh30Rb3QiC9bQaMRuLIBz/GpNKW6IMh6pw+MHOVMX0wakCJ3dgBCSHPoev
Sa7cXdVa/MfBPvCsSllmsNHmhNINfvxnsSs35tG6aam2lsknGLig1Qkb5deK
ZSepBYqB0BAK/zvCxqllHQdAgOao0WJJ0m1AO4mDNUM0a74bbMd4l9NwTd6K
lDZxPM3U74JCaWDT0OPyr+exXvfXkvWkjGMB2Ylctt36CFx1cj+uX324lPtH
2D+o9znk3hUz1eqX0OAnRZZdEsqPMuzmlMKK/bLlrI4SsGP3R7yBZH8414cY
KE4RCKVw5sbHcaC8s/J5jvXoHjGrhtaNPYZt8ZwBTmon5cBGiDylzOP8lX+X
jAEoE0V+D4G+ejI4Wnl6hDgtTdNw3RB+5XmMnbdXo9TlBiR4/Pdus/YjgHkV
Vk1L1DXfpw8f5YWqw5fe1OkMdYha9RKzrOySGo2smEPyscqB/snBYmXg/b7u
nJER/BrNYgd/dpo028DYEPojr8mV6zl6NZToaeGMGCc9ZGGCFjhk8rLNKgGj
yvLUy+NKUMUL60t/QUQaG1mQkbp1A6KHhB45NmWClE86uVmhl76xdZ/91ciI
qXRCGkOm0iHBeMyiS80rrIRX0iy2rCzC2kIbNiW+u4pdElBqei14YvVSe0To
5v2013Ukvt4a65ypXhFosTHSPW5nMEg58rXo5ZIWljTi2cSDAMInGoVbB2TC
bYSaKLFPNo6uEXFqAF+/IOL4/Usr7XWefu1fIpaeTIX1i+iEXzP8GnOqQBij
HOAT5kDyHLWEUCfGF9m5MofHdDKY4RGVS2g1TDz56k/8RT29+/MHZqIWgVcd
fIzfkOlCLxgzrMHWVozbdWOvzngCJ4oaE2lO6AfwVm4PSBSsXK8UWXJ55tAi
wM85krRElbUSZ0gE0FTP/IGLEblgDFCWtGAVzqwZDyPx8pa+DVbjamEU8pm6
XO9SqZURsJMNJNi2kzoIvzLZpYTLxuwSN+jsM57pfeP5EnLB69ypdwIcuxW2
3Ugm0PIs2jUyFD2Ec4uVZMNkvEPbi2S/rdwPuaOjTkHwyy35v43uE0P5Mgk+
sPlNL4HuYyRT+nO4prtc052RTVPaSas0zLeg8T6fVPasGb8D1HJAnDKNZ6XO
4UB8aaqYg8UM5rCbgoKTCI7mrF/PYZj93qwAq68XGFHB/cFLKYIxVZ5n5De6
XPjKZ5hSNcSJdoHHDHYJgvXLjCEC7W+4kGo6/qAWSi6fJtC0wv4udnedIclO
jgGG74hZWHbkg/GAghL7uV24ToBtWrqPunJPQCmwuoeJcu3otcv7CqHEgsJv
vZd+gBlJ3NBc/tsEwQUCey5e1hjdhmWHxvUhTLfVrwRFN12045N6aQGyFhGo
+/3J7HKsAD+qkCHUcjMdpkZbcPJZI6lx/gJIPKpUIkv6Iuo/Kfna9AN2Mb3H
bMws6tJk73WO8IiOV6DR6vmE76A/YudngFXGzIIjXqJvRAu1203XZ5eO5lLH
PbK3aNO7Xmke5gVIRrvonzXA6jcIFkQQE/3UQ6299M+6ttvBQr0NzFMDqQ5r
ENtTFLjjW9lp8IYI+7K2TV3dmACMicWXQtdeM4alD3fLfo/q1zuFuB2Xe9yY
ThLdp4I+zVKzbJD8Qdjd8Wtk0q6miNCgJ9rtBJbijYDlWDTQ7JRK6QE+Mlqa
Ckz9oFLMzA5wAwY0ePCe2q5LiEmMonBdGvr/ICpl0LT31e+yBGgGT2lWyZBT
CULENuWsJ7mQwQyy6awjA3qdIYcxIsPaowZYB9b8ZNFw4eFtPVW3g8+CQgok
xSY/RjnU1KLgkX+3PIFOBY/MtVWAukLm76JjjhmRwZBUDgaOy+cEfu5+N8jb
nm5LGVVQigH1WtSSrEkucxUXsdcU5pDkNQNtoAspWrZAH8PuYRiiQNX45Ph9
Ef+9fjofZqzymciTwwJvj2V/U2lOzJD4TrsDOUEU+EoEBvVZPvuez21xsuH9
Jm+OQb5Lm59LYTvrHrmxQpL+46EKpDztKczW7wa/y6J/PXoZqosMzgV6DNDV
pitoO+KXajKWvKB83cgBE2Ljzz82eSpFIQnGgzlJE2+2TQJsgGC1poPeP7lZ
5MfLstvNlPcjVaTaw0nAEMs14fNzhgvdVLju9chPvPa7rBgGV02NNeaSAOsf
RPFFKFXVkrzENke3Plluga6kEtLTP57Lyp9VMat7gnED1sfbbYpyJpdPb5a/
slrYhd1Xd3P1JvxXcMfu6ZchZaXqTx1kkNMVhqQJQhxF3dmbunNsD3CHpNB9
TJHQZGmqKku9yWJtptjOmU9EoD9TSps/8D6/nonYU3byH0Y+A0fFj5u1Tfk2
dCOtZau2vqeLp3wKyUu5SiPYc1l2Fq/YXRTFqDncg/r4Tt91RweSAd809PH8
Oc3VWTxnXDTZmohu+3ZLzMqkeD+spXlXilCKmzpAHqUKnwEkZV3cBJWugP3c
gmUZwha1YSOCVRM/Sk53HxzpWHXU+OTCRz+O+Z1Z3cXk1pQqTD49rd7MKdnN
sw9HNEdU3dqFtnnWJS+6CNouPSGuviy5XICSFuQ3biaq9ICWvsfWPQBr827X
ty7cTZa2+4lj3fR5bD7nV2rrbUq+5fcQ9gcEjgiF94V7OCZBzD81sEsDlx+O
YgZm2DhSLG6aA83tDeBL57kVnK48WCjKgMaa21TqLnK6IkK7hPJavEdycmIi
KPRFTlHTHikjqKx28bztpzySBqYADTJZA+JcwnP8I7D4m4PJrDkemr9KRqbD
V+O4UcpB+d57BTi5WycU9+nxgpBC/hN6gOPMUoxBiXNfPY79VMcaRqqGB6uY
/paoc/TfbzolyuH9j5zLvAK3ZBupolCFMAatiHGQW+5F5RuZ0qf/wEsMylvy
MjvKX63mlb2MQPrS0TcHLRNFbFyqy0+yHsHS0uL/02/FhPb5/vhz5Y44Gjh8
scSzMZkWIZypNKr5ocjcFcyIdFPGEAdp0FJrxyIb9eSoSVudLSj3FuIdqUi+
nqjbUMorS7r06oGXXQdJ4oq/W/PjgHbdfFpxueelwI6FKuM6JX0QkMBeynCh
BjHEXlzGpSwMA3l+1uYlG6n6M1iylEABl+OR8gtRN3gtnv9P71HB0JNWgdPq
5zKwU82Iyoy3WSW7aweEq4OunzhAF/eS+xE1z245NJZQVfC/uQMFzWVNHC1j
8/y+IihK80XyLtNgJSpBpRban80CKAVXNpuzo47xdetM4Gfwg5mQGcMDvVC5
xe17x54LM8eZ7KGg59TvyoHwY+lCXVcmOcJ7izFehxlD9kZyeUaycAaGGyDm
u7815Af7/apa0QBJRQPia0HhoIqF0imxP7i9EEkYeNdDPAD51nHnUOLDA05v
KoUcXqGbnj5+4s3m2s1xaDgL/dbbDAmUhEsASNCAPEUZ4me+CXffQJ6ekdjt
nJfWxvto9O7QTXyFg0dzDAShS2isbLtt0gojelK7FGbhz8EFWco5W1J2wfol
wZwvnWhxsIazlPyPGdfn6MGit0v5SC2BWvLi+DuXRFFLMcgNY3Jetgl+1sVA
QvaLYXVKTX+MFqTGWFFQbKlIpDTyzFXMNx9/rPG5QrETu1Fh8dZNuerJS3xO
vmSa0klTEVNLBxObojY/lcy/rkjbM/8amjHAcjM1+3TT6rlA4zFwMMFnXLF+
sy2zB1B9kp57w0TfjMnk9IVbANv6u2v8Iao6M7gIANTJlUMGNIVwTHt1TReb
o26c8y4yu35yEBFQZZjVp6vDysHsxrxP32Pt9Y9YO93xtrnbJ3zJhVngmtQv
kFfUfi//o5nfywGfSQbGVKqBZteqeyRvr3GYiZgFlBoJwVmqTJ2egfrGevwN
tnH+KdTS+G1FMHhk2E8mpPPKvzWET7pvS2Tu1cgx/3EObpsa0Jln3J/Zyoja
QJkEHQaxGigQr0kf+XFN5amuimZBJNitzLAQIqoi55mx4XvW1G2GuCBt0INw
WsoYVRAlwcwfW0BVHnLWU5Fc+MM0BVecBYoGbdnOMKbcWiDPD4bQsFU101ah
PPlxmYv124+7OmiIgzmNaMOt9jvB4GhW0aqhAf2neQnWfaGvPdwxMbJAoiRK
Q4R2pW8lwqyTYeBQJSfiUb7K/pcktL5q3Ze1H+1JWcqRNEF0KcSQCBiNpafO
8KinW49YtURPwo8UD81/FcxlotiInJ3u3vWkHBfetZ0IHNAOr0oLLQ2t5NPQ
i+bG01zS71siAB8ZhbK/Kyp6F9FRdBRBAEx0feZRrzm6k0nlqFbqAU5jpB8A
MuhXSNIUZXZAOApJwrMv9q4Cj40bjCso0Su9Po9RZnnT5eRrQW1PrtOfoy0W
ic4bU+iv8T7OMWiQ0muZrjqPffQkboA0ePzcU5Cn+CZ08Fn2djy1XRQUGhb+
9Dny8UOelMhlneJnjppSPdy3pPxtO26S4wnbh02lHaTypEKsV5Aq1zn2sFQY
eKk3OyhT9JEHcngtZo5Nr4gztiI+sfUukyqS9kT+izhVoxK43KR5B1HRCE18
GqxMLE2UBnkodgR6RqQifoUxAiFf7xrYn4j21ELch+Jkin9Tm9uiOZhgucVy
L/bj5U4cwyDCrwOpyzuIojrca2U0k607cPqS47RAFRKPYw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+Er6HAub3m0O9LNH9TIonn9pxsicqqkuAKswZelNs/HH+l5oeSINz1cVLKCvIyiFI3j0Y6Vou38qHSBoh4gzRuPlC6sR2XvDCt/b5cmcUc8pu7UMFm7UrvZMMNv5Hq27CjZ239xo+C2ubsvSaj/q0hOsO1I2Uadvg3uSb5+B9eukLx07YDQFliRmJpy5BjwMPm6L+ow2ZVeACaqhAcxgX5QFamK/UKz5PQuRgZCTLTI1cQfeVHCExX2e3V5SuP4CxuNHEa9aCD6TWDv/rwarFmWPRlHwfI5cqvmmVIezCgqLyp+MDS6f6ANInoM0yB41bS/+i2+hrap0BvYtPKcmMPXtpYcV1hH+tpyknFAwTRTVgDBCkInHZzTkinQyCmO7zxjWas5qqTikmGwVSl3nyyPPsvI0hR/IxiEu98E2l4btm7VfcyVCJ5toU7sUpAO6eGtfSwFufSku+/lleDkKpHorqcwBc5Dlu9DM2BNzRU0JKAvzlZdFJB0KzRTxAyXd2Td7sLwxaKzU8UuYx4iG3ImgWlogtLDIuoEBwz++WrtZNC8taT10G5+CsVUuhEFw3i57H3qoJ5h/vD9inZ8VU4gbGjsHI5qf9dEJ1liLJ/orZNO3TbcJgtM9u0qSJEF1FmvL9upFoeg+x9faVnDgZ1Oz2UtCSuIBLCNzhC7aNEV95sDHW9rlOochFgx7WgYOfG6jSJ1uKAw96YphzZ4bSUhCb7RfAE9AONpXMDJwlh20pJtBz933OK3OZL5Qjif2fnDwx4alkTl2gTWSW9aTuLlF"
`endif