// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
wx8W8or5QCjuFiMmznrUdHWiNZjprsHYfTi3e0rlIPlHxUJu54ik3JFVLFxl
xsCQR7lOtutzNF6FcBDqFTWwQZczGUca0ZYTPY0BU/TgQdwzUWCee/e12vJE
mKEbrk5IG2Bb3deDxqdgiLNLLSIEv17EAivMZKoj6jQPYsvFd5cf/nyagz62
Y4gKcgH1RIKvltsWvDGCLsF+RDlrKYvCAuXvRd1rE0XEtZbA/jqD9zkTnfGA
IxvOr378ftUCrImNOmxZOnTXTXoaK9N/WFGDpe6tGkjnIa0Qtl3nIhYYB50K
ZwD5quaxiwXo0XLNjHCZWDK+VvnaJMB1jmF7hZFYJg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TAP+RL0HyTNwO7pa/4lSg4crqwT4NGHWaEdlqKs5+ykKvGK/+T7u5t1KIxIC
A0b0ER8n+cAIV7cMXXkolPMICX3+7lyGqm4dHA01Px7HMu+SorLdKcirlmGc
MBOCOrJrRHuMM4QhhVMJnovcFIE71blvzs3x7Qu7pAP9ouNaIvyiGyrYoK4F
CRuybJr9RJec4kVOh/fYxgsB+6n2oUNBM0B4WgFG0v9pfnJ7vnkc3AktLLWd
51zzxn0GSdglps3gwUqHx5MK5P7/buuot7O3Napm0MEB8sTv9X7ufBM9Bjii
Bd4l+n6X2PsZ3kBej8yP+Eu7TkarpucdQ2W1N4L+xw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
vUbyg4/cU62ZT3PCI/3H7B6VzzTZAQCPsYdhy1l6hQeNz1goeF68qwZwjSgG
kNpgDMll9R9K9viA51zeIMf8tkEDehng4QtNWzaRXMv7/XMvlrVdOlGyyxN7
seVjPDuRfjb/iuGMM2w7UwaOHDrS5T07bcmMTxK0yihgQjm6Edhbeyp9bej1
dKXytl70v3CLe30OGIqzJn4sSr1JwJkbqpiRjdJL9V91u2+1+rnKMRzflGRN
f2gtQkrZAxsIFr/fsfe5epjNI51RigKZ3p6UIMCUdFaCzb6R5JEavmGaHsBc
bGG+RMeqeGoat3TQHLupCBSNNMHJlxQFI8E88lGgdw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dGgg3/y1H6XFeQVJO+nqEPAfI3g/G4qxVbv6qLYpQWLIuD/iTMK8ABh78aNc
ukjbefG6SDK/3eVNTZHU3eZ2HxJoviC7x7Hs+SJuPMB6s3xVFRYcCftaat5O
HSgvXNaWaNwOXhtZgRQOjLPSEljrP+lcy5a/O9EgTKBsyNAOYOjEPPOgds56
vo1eqHo3hN9njjFCxGbuRA9I4qQgzyl2YAFoP1p8jYlB0eW04gFono33MXqI
LZ/L2xvKIEaYFG/+QXypoAHoe1Pv9wzhjR/pEpOVNuESf4T+PPL6VjUq6L8N
jxXYQXrXkxc0Embn6yOyL5hexsO+FDCwhIUpgJ0ChQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EKdSrqvunE7PozajE0s1onk1uXBJSnPVrjvJcwJELY2sa8d327A3i7Jtp9zK
f3ptjCs3onwQtL+CP02ZMoxPGmXpaJ8fF/Uo2T22sTPaQt8JtdA4Kqxe4CtN
YwiNkmg16DYQHAdfD11qMqz2tDmcBKmfodg7sD3Q7asq1BJvD3g=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
CAebFwD4+oPj4QLHBq302HVm1o0n3zhTgk2kx5d0SVmUg0OGuM1M8pak1Cn4
rR6oJoykqUCBQhtNaZqa9BDuvgauYTlR+9UhMoJiIOtKuvHEOH7FLpNlf9KP
ZzrC46FzMKQ8sqlwX/z7y0VtdL/J49qo5nxQH/iyErDcG7wYNVOXQl/AmOKF
HFeV+NbLBoATmXuYju0MQr23/LfrfQ2HDBSNP75ITUWehTarQnr2Sg30sL1c
22nyD5a428433Mja6ZereA0mjAfdU6y30hdkzM9hRE3tnrrH7f34gPHKIb13
+AoZaw+jWXIbNPiTy0S1i0aJ1Xrpzr51eC+O5JDY9z0beBKT9nC0YAQqA4eL
A6udhHt45/19TJ3xMU4vx1DQhH1OcnQvF6j0tIZsY6D8uYthQziZI7TtKDZU
6pWZ8VdGBDI5ajKiMvtfiBZ/SfawmMxq1I3WWas/DF3V/xJ/PLYMd6/Mn9mf
yUNjetRyawmeEY7DVlBBNKpDFoC8Fet0


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aHdDfVLqRRgfDg1lNrYwQCLMrnfFjG9duU5TmVEa+H/pKPfaLgkQCssoqR6c
isbZpLif7WxSHchY2VfrdYbjGCOoCwcV0UdC/h2ZTjAFYk5omUSqNDNbkKsK
2cX8o/4PeOOXzNYy2qzDv9VEsHzI+f9NcJbMVl9d2EGVdmZ7iQg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KtRa41JlwqzoCtg7DNInQCAr1dmjUEO2VaNsmVbZn610LLz0JaAeqFGYwBn6
2a6O1SWz4/4v4BNhuDkUTwCFPa1fru+qiITmPaYul0ntoSqeKv7XuMaSHR/G
P1tEpNROSt1SNSlrxqUWB+JIAuBkU0wbkeFZM7mhJ8+BjCzL2yg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 26032)
`pragma protect data_block
o5XuIMsy832kkQYOvxJlhOq/Y76enH8i3rASPiokCQSHwW3L0OQGk1WkmgGO
oiQUdrk+w+ZfpisTFc7HBvq5REXlePyQBAQ4x6cRg2CM9IXiW7MIGi8dsMku
HybSCANR3ez0hqECNFyDNOgwxBWnOvTPiFb08nXOHgQGjOd/sWF2P7Z4eDTB
sGolOL0wF1bU99rrJtFUnecDnnH4lk5K8RoxPcQ5Yi7mqy2rCN2oUnseOUat
uvvzVNuIoqpRxyn2/Rd4qO2Fa7D/acdMnXiP2eTVuFMiXgscJG7KS8EY8hNl
gwEcjT9E7f8muGI16Mh6QGtOWq4YJi+qrhEeQsLm4Z+OH7zD83H/b11HXfSV
71uf+86IclLULw3QXv7iCp3dAl+7oDHNKNmTflXWczqGUrC5Bi9G7AKKRwjW
YlY+CkNcR9IzLPyveuLN3c/IyZUX6D3zOXPw6bMsUVDRV8oJ146m1njEHSDN
vS8zLrf3BS1yZmBGFklOShVX2B45/TScRoeOzgQZdJi5wNC7wV6B2gut9Dsq
yk5ZDBCkWulc4bzX+JeHzAF2EjkmYwDYhYRo0Om5o1gdfJBp/TCgx8vl4U4D
pHot3hNpQTXkmmByBYLCNdrQf6KGLr3R9BGce1biljXkjTt0AagKzbDzq7oR
dC9E3523ASYBA7R/J9sqSIGziPays+itU6MDRO/9xB4N3Am+Nl+7yhkocv40
T4CjOig5VS40SrmH4SK7e6E660aJ9tfvzBCkyBmAWrH3cLZidntbKRzNjwzA
E3lrx1UUTiJQQYA4fQl97NF1x1UOzOMETskQDxDSCaV7LCjS/eb9yXxPBnYo
LYcRtjfXB/deDDNx67sj252BkpHLouP39LMEwt6rgVc6Q3dhk21gA8gDF2td
TwcwG/rlcgBLyoAd+nbF2ZSrEgoT5YjmRjlhKvUaRcyj9GJhQ0Lip6RVNQ5i
Ejy/POUVeORUPfZ4+00h3yQv6qeBV7UXHEQET4Wx8lntrK6hTUSPuHRlRcng
C/QdhFsikHOgtAK2iHq4++V5UlcCcq9DINhEaodOPstX+fBqrzo+vIdUh23b
+KxEnSo2jgdv1uXVf3L30Rb2RVBx1qY0Q3XUninXwaYbhYDJVgdKg6TDzohf
ntM8YWLgA8Q8xfJM7FecSORcbDY/WOZoh6bosOBsmKgxUSIffK78PJ75VP7l
i+DsWxgRDVYBF6VLrx0In0qY5Vf/jKo3GwTM1hY6uBeKcvBLfy79DCNkoJCA
P3YnliqQEygZqhxR0si+1gdGSs6Ijusg0OPP03dZkVK05o+yVNYE4Kqe8b8Q
/sQOV3La5aTu9MFI54OdZ/0WMkKmBMm9E0fvK73dA78bm7KWPgA7PJPwVXR7
u7+1rIAIJ4/L+l6pGeN5qVoBNVW2qziQYPS5Q41G5ZLTrfyNVd5hm/Pjly0x
f5IfNFXK6vUDjB15Fu1faETiPjemTw3HJZtaUIj/HGR8a0gyW8xRbkLF2AvD
ANsWCCryvfmsglqn9lxXj2u0gPRYN1zpSskxSh+q4oSBf065K10jr6ACd6Ch
qkWLW2M2BGqmQWGdh+Xk0xHOpDtgSi813kaKrRiXUMmk0wtKPQKCtSjgSm/S
yMIxC95gCc4HumoPhfujA7vjf6ttreV+NFtfVWD5qpdvW2GCtLsBuCjvjRox
8HXLObt76D1AkDKHtbssgGe5AMxtP2iopAlbzA+/NoeTj2yYMUx+uOolTQat
fl5Ih/OtC+C8bYuJpQmiRntilPPM6yEOeBE1mic/vWHXSSyd76TELq2T6AVU
RSZhseCJhZ2sed4vIsHsFhFussGLivC8q0iebKE1WneMRINcK8RcC/r1NAPA
LPqmROTyR08BiFCqFRzrneG2vUrIWL/GgClQsCTYQ3YM7o+ebLaSbcxsSllB
0UDHksYtCWLe36sVVTcmTiWEgH7+xfUQg2dW12ZBqOtnrr23ymgxA1Xfp0zL
jMKLV+m4R/d47vo+IaAndYaXR4HBTX8Nxd17RNdlILdzjlncEdoAMjsJLzz5
ge1WkklPIsWIYzv+Ryy7x9SCu7bJFdpF6tVJrJLzv5j5oztqXYA2wl9g7LV5
kvry8dvJCANz8c8Bq6nPofuZs3Ez+goeaeOYUKioKYigEB8VMJEenq+Vf0kj
6y8z5OnAN3dHyi5mOchtrCiD0YejUTXf1F6vHR7UN+q0JDOJJw7m10mqOKoO
o1Ms3nXEhaoQzO8h6ZIEuVw1Vad9zDwYpddhzFqovs+PoKA33MDEc+bqPq+8
qmJ6nKBKbre5KPAQFIbyXUOwu+kKwHXmtjbw7u0lWYCgQMC+wZwvmFrZKz5X
7f3vQldCul58ELKuTqRo3wSSIFRWbeBtt2Ddfrv1fcDwa1DH4e3z0+9B3+1r
TbCzN1RziWk0Fazo3b8h9Twd5de24xjyH75Lhit5IzEWGqA6bkd5yTaImXRc
9RusGCTGPlLMEsmXISmGEh4eu2nvO5KMyVGc09u1JsTMyfX5VQOHscpSB7oJ
kUfVXTHhmfIC2jtPa5rirqQetdbd6gxL+6+LXSROPaLpk/SGCDVAxAYv3chr
OMVubEehUjMJWPDCmWEgk9fUthp91NcUDiFi86q24t6o1JUMEFDSVhA4uhUk
sYyqprPYyhOgR3as4Z1pn1VkMOpIN3gh8ydEZkIquFnNvJ1qyUwLVls32BrS
vyz1jQBTBqac3nrj+UXkyyR60jzsNTgHNcUuCRVikktWZm56CDRwF4S6QRe5
9FrnvIwnYxBijPoMJDTTg6QPVFjY5ElBU6+dkjWvBJtzrkjR5GjIDEY8PmCY
5nuNJfncJBAAZx/0UFxAs0vt7tqkrpBy1uOdgSFQFis8+cPo8VMNcA+0pEzr
zYVRbKWs6zL1cB2Y7e6i9yfuz3GbOa8mErxTY4glOKYrRIDvxQKsYHk1I3B8
RS7gYMRKUNW8pyngRjVCNlYDSj1ziUhp/ZjNTLEsjJ1dsLpH346dpOXJvbDX
ys58FeJ+5xGWJdbd7nrnWfBbNB6L1LjdHJkUEUEpvGz/8TU+JxexHwBZLtpw
UoQq1AuFaeGjiRbq8ZVcdi47EeKgTPvLaZG0byHdVpLtGU8RJYscI/IkQDH/
Rg9XD0DEWlSCe3+xdtCkRKpbkvJ96ZILTdIA9HIBNa1LameQv0+UtW2Fc31Q
gMmj6HtIUVh+6YwVzgesP+MtOyyqwm7Xy2UJiSgTQahnsHD7o+30jOL1DtLV
rLshhtP6MeT/2wtZffYs7s2ZVVr2l+1bTJoWm0WRumYHsD6c1FJzJN8cWH1N
JELxevIs0/rY3tDdv0lTjubcWio2yhDoT0rhvgiUTZZjBnel7vmjOvxdelzC
qG0+J2c6OCA0PW3q3F9KXSNZ/PZ6SUkLFxMpj6rg1k2YVDTf7cg2eJJ2wmx1
O6J2+Slmb7PLJMIVnRgAL9ymBaOxvoSLOPcJC3VjUwuaA2QULUi/etMfVOM9
EGR3G5P10HChowrP2A+r0yS1RxU1hV/7IvQz2q2vds/2/iW72OYsgc/NJPbJ
B99ESZcwdAmlYaX2swUMePLXEyEH5C6sKPXv/XVlsQwXpTuuRh9iOX1D1g38
Gu5sbzXq6reecXEtLsqgFJMt2m9FY7oHnDWOLfpPukCNyAbDQJyyvhDgQTgK
iE1dDn7Yijxrju09WuQoEmDe/xmExUL6VOjNZY7m7HNefXUKhsTvgp+W7m0k
Xt7q4z6BJVT0AphIRIBKuKT4BXlFeUJ+VyWJZsAq5hw62G72WURYAv7Xc8D3
U2AghURjFcsrSX7VAwqIhLSobMBeMAgLFyBr/P9Q5jlrZL/kx3WyNHnpy0fN
UiR8bIQ2g2VvN9Cl3+5c6VeCOgwCWzKHpNuDHLTXoj0BsUcsY377HKlcQRqq
Ex040uTYlWQzFvYfKlBcoH1t1D9RW4iUh2MG9uo+QfR0m4CD2qJgR+rv1Ap3
eJp/AKLR703fHBhvgbVdmNzKyfKVNeTtPZpYVUCeeLriZDM7McXNuKiNj6lR
NlpF3yf/7rMVghtey4NR7KWaM6TpRX9uzF7wWp0T/UOgR1Mm8Czkbd1p415W
7hPlRmrW3+nFg6m4UtHQ0qeesK8x1PfoeqtsBWbpm7U7TTVi/9tF3W2hmoVg
y+8xmmvi87n+I+5rBbqSYdoYLRLof5WgzmBWCxap5IraMgIqxkN41bmyq3vW
0jWK80NvA9+VkZCevGwWOg0ek73m4aVbnRGORYJyXyhmVu988todVgGabtbB
bJEQHkDq89hbWhfdGcd0iL+qUaHOxdYS7GwZ78SnGdVKFVRLHqTR2/Q0AZkn
TfHfZqWuZt7DJdhaitgu1u3o+/I6fPdYKgufae4J+cIarFtiuUx777NUZjn4
cbPcp8THSDvLorynw9wiBPtjh8N1SPqMPOYvabsdAEzs7OmFIN3I3NzISmaI
vcZ5f6cTwlys1a1CvHDMFKPwuZj4L9i2vzCAmUlvZ8o5rvXzEadCr6zptYog
vHGgDb/sR+zy8AE1HaijjCbqJaIo92yMWlqTsKoHCVhaIgQKQXWPNExNo+Ud
27vjWyryb0TXoqeX3gzNarGh1nr3fqgHXxkMZ7YfBiAJhJ6EdE4MaVgnfyf4
XwR03wfayFgNQR6AVdEAE6U3dlWADQunChsQ+GjILoXq+cAUylGyRu/G2kLU
U1Ukc1NQatK6/rHJkFGclxhJq4gTloztVvQVICjNyE0KfR5GI4hKYnH4uYPJ
57QZD79TwMhSSfkem2xS3NaJlZqfT5sKU0NKoXKeD2rFZOf1Fq0of2z+YX7z
7P0vzR/PRoNxlg9rLiPHQd8oCPhohYjhoDurVsvT1qNbofVJIx69kN9H/Ycu
wVvrfrm3W0sqrLv+qcmWDC/7Hy+wDFWOTTbwObOCfZY7XLBeEg6hjlBXziL1
1v5THMsPM6CvTasmVMITFtb17vXzJ14ZZwINzRxtcbEeE3YbB5kBbEprO87+
JaoAxDxtxTMxY8RaM9PN5r1PWmIe9S6wz1Npy4DDfqsCH4IKJGU0TpfjuTSJ
SarnMKgEKDD8d1XeEXNH78LE6it+2JGwGu2uVeM2S3Np+I0nPw3HXRzmv8dA
qRFdAXM5f17kRLsVUc4/bxjAv+JeVOR+DN2RQevlHfce/4HLmOxINimR8tFp
CB+PjG+pi2T5hUhs87lsFFQLf2ETDXGV3znJ+5p7BAq3xJDP2bM1spCUm9G3
BqXeTGjP3rVaTIke3vOkS3jn0UJterAuVCX3NSocz/TEvFbJ6udbmaV+Zszw
UNxoDznvrTKwdmbSVOUnTCLiHtQi00iT+1X6UzfTEEvRnb1ShW0z2s4gPNEs
OIKtQWasZbG/PrIcUXiMTPAbCGTJaxb7LS8Axde2HSG5JkK2lk75QuPb91Q1
nzoNuEwxfVtZmr0IGrcrDWtGlrhCuA0kqKJlurblBImzR74FuRcL80XzkfKa
Ksmh9nubA712ggL8fxIduv4VgWhVwhyeuIPVFyO0LPwJ0vENnIBt7KqAELny
HgZoOVqdYm/cf96G88I2LwxNQExXMXtA/WVXDEmUoBw9Yv3hu+M/oJ0vR1Mu
wwqPkHLA36Ibi9EH+rjLgb1nmY6LEZlzPZjAhT1xtVbGci9ZqkKeEVccApvt
k1e5aA8SeeXlk5z2s12jEMHEOPKilslD2VQ4M71sxFWTS0CHtOq9/0RVB8gk
pQXWDF7sijNsvq9g9FM720cYmUz4+/TlHsU3PGd9jViQR7bvIFyoVYNB8cb8
+Rp1l+8e4wmJ/PRvifAb7DMvVeqvi5Y1KPzgFfG45cZRfX0wd8MqAwl4k4E0
MhvV83lpMo2nOFkrxlhmmG+hwpSn+9PpfaApVa0q0IJV6uVKiq1s7JCkYyL4
9oU5rvOoQ2A+3W0kDvKhQgLv9C149Jq1QFvemrwuJAElA3wDaQoGa90V0PIL
YBw1WdZwZdtQmFihpEx/ouu5eM1CALkS9zSUHaDJbTkYhBebrwepLlAxYYkR
N9GDnoYNhrllxeDDgBgWiZDghOdYKCzh0F/DCzxFmsYYVLPOc49iH8y4zpBr
Dlvs7lcDZ9k3/eHUbTEVKKafUp3CT91zuvtk1OSKikyAyujaYNgUPCsXhmlG
cCObeBTIM0PNYYnsNE7NPVlT558HDuu9ndD7jJDYyC5zyTVo5PbTIYliH0B9
60GKUIYcK/8nO+/XFoyNDBJJHlLUsQWRdvPBozBT7z9wqR9OgCchGKVRqS7e
LXHlwcxC+giCQpBMhoICJVWeK6vw4AxNzHnsmkWdeSXaP0UkK/iasawL/9/e
YBTDGCp9a0My8GkpCsXsGA3e4rmlE9q+5hQEl7y1tfIcFTUfnrhKonu7UOna
h5xQVVYseonRfeNR+b4zTvEfC02Z1yd+jJMTWGXhyCZhpwCaO12JzAc8HzWp
V/SPN1cV/0hc1X6OagPEuwVFsUgOdr7QgGVIzb/s9XBZTLoBuuLaz4HPWgg8
7zZ6S/Kf5yWUJWtR1podW9QIzpyMBd3X2I5FDeXxkXRsZzRPLZHlgCihiZ3F
INGjkuQ3w985PDzcFTYgoRLgpLVjMk2XvxMqDBjl17fwNuNlVQ6NVzXBXAyo
A2N3/BVJwLs8WLEMLSYK+UWb1/c5d3Wn+XS/J9tyE+/vBSxvNIRhLDQB2kAH
G4pj0ftkFudRTKXE8OtpJfyNdR1wTActmSAmeLMaUqJyf2XaP6/Pj7hnhy9c
y+wsSwkaFJRRJDhexy16Y9aDSAVPqKmRbw7wM/TGpNPoJi8/JoBwJp8V8Qap
gj3x9UpZzRlPgb5W/jDGlwciYX/17tsYdVCOlH96oiiazNgAaQO8E6VhasWs
Qog1Hyj/yaXyjDe9mO5GWlx4/vpP0mcjsp1Dq9eoKSg8X5hvKN4y1++/6ikJ
NDrOd/K21iDlvu8UAF4bhTyaF+7cphjSiBt2VdsLQyRbakUWmAxC9kpHTym4
G+SGGDp+rOJXNiO/hYkIUcXIBKrB01OOIinf7F0wCQC6pQc55JJ8e0OZu97Z
U9t/nAedpqEAkPZ7llgFQqsGPqoQniYGdxElnsQS4ffsbKjWFb2t12p3IxuT
hKROMZo7gPyPc7IAzQjndy5Yy7TPKUSSyYXp7Of+nrY5sP7fgmMV1O/+MxiB
bkStl1aAR0JCLre/LcoPjOPGwrIW8oukBnCsQOZPshfDm5Li/UAHvmWjEaDp
I4yFmKMTvmIbpvmJx4slprZISgO5VU+/PAOFozeIxvo/lwzfipCwTRlyhVNO
r0OrTO8fCkfXy+U25F9f/KmwA5aiROsZwf3rlTIwpqCZ01D2LytcqHzgK4X2
vntyUK4T1xoDpPS4/OfxPUzIjZlFiJQcOx/0fdyZk8fBXrj+p+7XfL9Famkk
vIlLeZYFpg5SXrD7a6JGo2J9ZzDlaPe/2fWnhE2/5DNkoA/+bEIEVmlagqF3
9gA6UJuyFdaaHlfKY+sCSy9Qf50LUuGGTC5Rx4lpV29lrn31MCY96RQMMKqr
KTdKCSK3lzfSxfcYbj/p7gjPbZ5Bm9FKucHcAb6PMzbbvdNy4nk4QAnEG+DB
r6ip5prIN3n98aFk3ut/qwKollp5TtztMyh3r8hizZ/MpP/XwGibvW/ve0Ax
et6j6pGW4+U1ejvCRrYFqlQcc6QQ7CkP/aSXGoq8QMVDcMP4KZeBdiZQqzRv
gNIGmombP0FKfw9TJs72D3TD4+0yqIymWY7pFxetLaJpALmFu6N8HFZ6b8+f
MA5BtnjJE/UlHg12Sn02pnsrkbx2AB8KGrXvgVADDbLISIzKdqmSq2ndsHyV
eL5QM4oWn+MYYRwUOCYu/iGNCieMEL15wPvTkXJmriiL86yYq/U4b0tq/qzc
aUGwzdmySXdbhopRkrQlG5EqX+22+VVsShJ/tS+Znw5H0V9pOmghlgIcpqgr
A4oSh1tVbYocptYQ0K1+PMZqEwelcF3iSPBBfgTaehBnvCLmTGOiL7cN77oc
jSSua4Ry8yD4Qj/mlCF2w+H+uEDK5FTQGnKJQRSxTkjWVlmpZiy35JherHLY
CoO1+avr2tSF0Knr9SKsxkBJ5/RK1MlHmU/CgzXvQ/ZT9Qz4V/ntatm3Py1v
389QQmR2UisoVCrEhubAV8S9lhx/HpKErmxfQwmPASITiu/CFwNw/HrBUN8o
FkOPYQDGTMVPS4eTWinkHq2OwkWnR2vqJd9FA6WP4oZIi3M7KaJorkoIwVqk
rnkiaXW3rvwr1zFcng3HM4SiciEjXcRn5sstIGupDITtZvePFSJcUsfAsRR1
QF2j1YYwaF949CsznAcg20jgKgjkQV7389WC5v/1Ustld+HT74y6zPyQzSLu
N4c4ANTV2H+lyUWB1ui2kqpdCCCkFWNNXGx8Fw9iLDDlgYM3PdV6arLph7sW
CEIgLFADZAOItPklneASdG2Ze2u9+eCo2xcQXLR0a4Rvpvjpr+yClIfZk3kt
wDNsO6xHRfw92A4fHwQg00qJUSDdCMor7Gv5dcxVagYR2gBWDDO1UqLTAzsM
tfnonjmLZNQ3dNwNJswHktTQwpp8joXA6lFcoMXj8jGQB0PQrymVubtyC58N
09TM80pwVzERMaqDHDp4X6Y6JM2COR/lmw/OxFz6hvAEsFJjp062iW3T5/UY
LU1PCIRUuGzijsfzw31ha5lb8Ee8/yWRjzJ6Dx7cZi2jPtsTypqKs1fOClTJ
wC2tVijtTPxxnni1++kTnAGGa7cmB8DwMEcdEzUJ25TIyUNkbRajLzb0LRmS
5mFz/daKTM8DRe0vh4Ty4bGg1JrDO5zZ5sM2+BwDflynWUcDjJUt4BNpX64R
w1SH0ArrHYUSZsaiBzZHbBsrMaPs1GqgRu+/nNWooevv0uufCfy6Ogk84F4G
KlC/B+qYmxiOmeS3aEDG3sXtq1qwSLxp1i1Y7Wq/cRU2J0WnT8MVupnB4prm
FtJHIiU9Ow3WNCD5rfwh1z6jSXj0PFbPrlHNVavj2pGWy41QNKgtufwnOY55
LpYuBDjZ4ECOt4xBbzS7vpYtKEfIfuQmyd18v33odpT5omZ7qbkPk5Og6vDY
niupSdNMcB3Z7gD4kflESVN9RWFj0mGzmYuzoToBJ7Vcxq6f0R8x7D9Kx66q
7Kwf9hIUmyG9zTfn2xS+/WFEWP+Gd68jWmpzlepYkG49EwBzZ0r2KQHyc4/N
qgwpvKpEVfTSMTCmUcB831Wn5M8Jy4EgUu3/KJJHqr/74BpLcKfx8Xw2yBk5
6dHLB+WSL0gZJ9juy4SV4yWnZ6k82sDxnh1fiEQxXVNSO3RLl5xkVAw7Um1L
jMHITfu6ekEeOmAxXycmI7D4eeuDhH1lnIH/QQ6lLvzusT3TprhRbnh3ZXBC
iC7IDC3oKGzN/V8pMnAwJIYttrzH/TLgq257NIcJIP1xuroVLUxOVtfLWqHC
g6ycJgDAtvMqYkbPjq0sv4DPiyzifldEL01KVsD+GjpQQ7zexCM4fUYJPRrw
E/9ofoJG9VgojPz105lQMs907kE+1I6FOyAXhpZYK2rGPfYA1l+cm6ptYtB0
NPXS6yxeDYLJ+eaSLvxN/YS5djHML6NtAJq6aNowAaiGWWQ3+XfpckmW4t7L
r3nw4EWaq+edke3c/Q3CocIxifxgQMFHzqGGkPV1AqO9NhAGbA7fvIgKXNMi
vwqd4ov1+gXWAqdVkBe57KA2/KDxhHGr/X/qY25WTQVSUChu3o2eivdsZY6U
sgaO3Bx25884SEvuj686+xwTIZEBxHTfBTzFS0p1mTb7ZT5kyzyia8dvS8sJ
jAi2teBOjqFxZHhJcRf+BFcS8QG6V27pr/my8BIBUjMREW7HlXaBqg8QBawA
OjBRvgy8rGgkoCC1MzcjnuVwpNmiDK27LDQq0rLk1E3RU2qblJWbPmGnMe/w
5x/H8PTWN8Y0wRrerZNFQIi/nlAkZuTs7nRnN84TYL6d7KeKQBYVklvaVMAt
YMc3QUXzKk7GsRamxQf0RqfcwGUR+EIgZvJxCX5qx9RVGv07bjxDUdR9+9Ug
i73nni2d83CMlog8J/013VpmzXij7Fa5fxxfjcsgqnaBCZwQ7Y6kbRtZF3Lr
v2xC0KTXhc4jH5mHC4DmuGDm5fKCgJ9aUPFDP8m0ClcZOYZxznqpfOAmtbTs
vfBFwI7siSAsMh9RSpY7Ws4kZWlvh39/CRVOav3Pg8s1U+INOepLPtIrJu4W
xg9KURgQW7CCubcvSNBMos1LKA81xbiTHOG1V8gS2RA2EQsoX4nfF0pEsO67
5bUyOS8HWCoYloVxX6I3pv0ae2Pu4Lfe48FAozuhc/thmTJcedmBAN/vu1xq
Rcyx9rwmToU/PjcLpFWJ9crK1jE9K1owE/ojPb6lylWRCalbTiWt6C1M/ugu
K/0UQkUi2QDA3We5amaL6pZeLCjbkBK10rIBELPhApCpJLhx3+DpkTz11tIx
dWlzxWqBKmRHsi+a4NmhPzTIRio4eaJk9iYadzHZasEo4ETT675coPWfj9rC
keC5TUa/OOH2YNLPWLfu/6U0KdxiYMC6NsdJ9RQ7L9zXyTw1AakzBzIZCcaP
UdHkeqJ59SjeDqggUER34Tc4Ys0OB2hi85SOwfheRXR9/PKQXS3vVS0J+9CN
F6eqjVHfwS7KMwPp7Wro2ngqO3GEa2noZG95MMOTvgxfedmwwmmmQRH7THAZ
/mORUKhU+Qmk1CF0LB7F3Hh9y3BAAt0EiLRRS/nJglBkHpbe1CSLJ72alqaG
lDTGyrBW/VBQyaNvlwCgqpQuwjitcRRRpv5OXNJzT24FYpo33AYm2nyQdImh
vjVIql1BtlP3S0ZuCbnFI3cnnr0z+sbuYSdTrEPQTIyZ7Q+6r7FENGwTTuev
RkB+//UnynrjXnIkeAYyZl96lVmT+UJucid4VRNLat5FBUqsTBGiLX8ZhbSv
jLYaVg5sRcVNzyEiUcLChIelRZ+u+892UIdZDrtsQxjHDpGePqPSYggJqQHk
zbJNp2CfPHGv3ppCxjC0ZUZMe7Lj9QjOPuVNoVYIEZHXamdwxrQ5Lr2kdqXq
Z96RrvpdAUDxnR/GePYlPhQ5gSXYCJEiAZg8juMSs5S9quKsfti8TnA4kXKd
SgrxHL/S/N/hjelgme7Ce+ZYxrgAZeiebjRmpdoMP3ANA6EIJD9E3Z4L0XYX
k/TicCWh4o+xFr5Ql5mysy2va1Q3ZJXkg94xqsNx8KhdJvRw1Pafi8Xxfx0G
IxScJz1H/K0lJTKusy1v2Q2CQmyCelrJMa/1StMQXT23vg9UTr63hHrZC4hO
6nWKkuNHNWlT7chSPdN5ImIUc7ntdnnephgGhAz25nKxpD7WBFvj6TdW+aEb
pnyC49MXs2gZjAlvLXkCJGrM4tsZEjylMdgAH3R0RgS7Mxl3U2QDiXJs05x2
zUNMpb4CYGOz2oqPKiDEMJ3MgrTWKyl0qXRe7SQoQ/IK8RCA7xKDsxiynVzc
ahURGpvpC+Sri4Xrvo4s5tZ2CGWbDVeHMjFmfGPnV5D1M1zypwG5Efmor/Oo
4yPrdAtCDt2BfDjdZbvMKX5HMoGgx9RYBUm/eu0SqLimEw4KIG7AK1Ly15Kj
iVSL41RkYeLXrhrSX3L8EQzgSrR7Y5cmwBIZ6z/AA1qYJJHdIjHmE0kY7Q7c
RxQvLLApkadrXqJGhSN/LyXA7Jwspi+Ijnswc/XJYoQyuy0K0lH66+SbqV2p
XH6U0PqlHQKtkz6OzlD/ZjNgw8SwvdiOjgHbOazprq5HCUj12vO4LP05i4vc
xioF35sCBwAnfdQFlUs5IrFSOhf9ud7lI/qoCb5ipUACI8gfmazbvUNkydIh
yyCrloHDm+7/eehI/hNT8YqqGF3RT/u2JUavZEDcyKf3RHBerH1QkPVsLMb+
XfkkrhYKWKdgYncxOtNH28qqLtEESS6rslkKvHAau6/5HbEZVlmjPT0TaE4Q
HNQeRIJO8qhdgDlw+/5Fjn3rl/3w3CQENM9WlLewP2VU00Bcj4EAQ6iNiEFt
hOBvw4g1oOY9sOHEQwNKneoD/mUyElwcgduLbSH5UIQR136qytSTqqnr3fOJ
VcflVqPUw+pEL31A3NTtF1P85/KqpMDgYcJCfX/lTB9CZSn5WXn7FB6/LhMh
2+Id5/+sYNsYouqIRpGBDK0eivxNG5g8OlqoMzRNIswJXO67N9mvTQBP5FU0
FtALlT9d0YnlQ+Y8pg7iTkJi1fASXkuuAHfM78fjzg03iNb1nXGvLDvzKvD/
P7MMuIYmezwefLtFZApQe/BJCqqTa8QkHHhromObfqDVGtKmZnSQA7Ajhv9t
QRjN6i+tXuuuhHaoLscGFUuEGPxN9EB931t471c61W+Au2V6JIyjsF9mH9+7
PIu7dphgh/KKgZ3aWDT2F0FSE73A1Q/rNhWu5hMCkYv+DO3uoziG/4TlNIJj
Zk3X4yvDaNrh21Kn7g3YXQOSn2dHYwH0zR9GlBrpUpSKSgVF0j+jUqZNesmT
1VFaFVFkjyXLWAS7hn2u1PQwsj5gHfvqVxLg5fgmsaKSIWJoRn5U7/GkRqfa
btRGBUWB+hRxS/GVQuO6uECwbQ6K1Lx2NONqAyWxyFj+D3B6BcsV3l9U/tYf
oSX2DyYSSe847jRZicQEdiu+CShOvVlpqcdpu4yZQIlGhhqFMu2CYzKS2eBK
4lH3kvtqZTIOAnDob7UAhWK7V4cX6/o1QhssBkKlCbGHOZRHNo32iNZph8EO
2/IRndVzlvSIx1GUa+EUdV8xlqHaLn/l7F5NOJZdinB+61sqfT9s5xp174N4
ZGIlpjPwXiDfjnVXWBNkV9rLyQxS9x1cbQ7eTrMTc0wSCF7rjApM5bCONoks
Kao2ZNKtpKyqaW0wYnbp/fbSEIorfBFB9uv+vQVcJZw2A6eblJ2xEXO/9TZn
kerON9qG4HQM4Zex/G5SISJ14XVIwU8XwTkOvDxFwIDJwAwwGX071uxz9/6y
lUEUhWjgMpwFZJAQz7C85nEN0kB4nyvRxc8SFM66YdfrclmHWoIPbAVQllWS
mttfFnb3vZ2GzemGZE3QVDLaWFXPju154s20eU/NJL7vytK1z3JI5Oo8ASHi
0WWB/jxnKVQojUFtjpaA6rg8J0R+GfCY3qXkWX/G7dtLJ5hOZ2Lbb6pZUGdJ
vzEFlWb4vEP/gqsboPfHiWB1u92na1E9GMGfWDDaCbnbDZQ7YD96BOmdbT1P
SMtXaMOMyC6bhiDWS+nk3Y24lpdswmQqiv9JevnVmImKverBzQRviBzk9fS6
p3DuJ4U5ZV0m6hpQc1k8+EOpdp+3DZ1KlhNrUSHUx91HrADajv1OHzEos4vi
BUP1LydRY0Nan4JozSbmbGwL/yZmLoat3w58dvjZAJ0UX93BKgk0mNwRA2hC
pXZgD4uLh5aS7/DPn3LnQpLkyCUsLZAuikxjtenCyaI71qmKIWJoDkxx/qp+
lbfFbpuDb6z4is0WI8ZlOkQX9uCd1nECq+ag423DEKS97gQ0PwxIeQhqDBJ5
HKuz7xtE6LiSN6w45lqgGe26f9V2kd8so3OoMlm38gqFJVqVV/2pvwlzVPm5
76Ywh41rqy5KGnN+PX7npTPm5wz0NJDfzB3tvkZTQ51npG3bMnMmuHXfC/Pl
vGtfWqGVznNXBzVK7lM9kIvXfcNtrqzVMDKgjq65AQt+k0gcB6dJGx7rZW+X
JopQBbkf7uyWgRtEz+c598Bs+cTFwqSEmlawpzS6b5ZoKreHZsyFp6C0NtcZ
+vCJckK9sZhmCWQspGXP2IGIk+e3ltxSCkrn3DA5yZWq1S4M5Wp7XrtwUd0N
a2vVEAVMznLJU/yWlGO5aomQhA3oGxSKRAARv+TU193cZmhrhaDyTS/izRu8
oJgCIM6TtBfmObbmLAfnsn+9N/gH6jgh5y/xkiHDI3h5G65x5v1SUBD3WBsr
zU2reTxoNNxLEcA6jkY8ag2QTI95A4cCBFaPjlorIB1V7+oGUG8fS3qx6jNP
wIl7NPSs0VDJgqgku4xyiS1UKEM8Y/OOr7dG9l8uS7d1i7XJ9bF+5lxqzHX8
5FpzG5zwuDWIGBmPGCImIpB6/qF0RQAjD2X/o2TLEk+V5rhX23/qYjlIqbSp
zHq53cudfJy2fKbAqNIpHEOAyEPTPeFt2Ae1IHXZH9K2+cAI1qy07fFW+6Cl
W+KbF8qHyf6HmlUiQkLugahUG8U11F+7rVgsIL+Xf3Olnwr1HfmU0apme0QP
5v9/rEnO7a1EBPiwUJ6igu0O3l9FO8XlyzfJJEz9JyM9xH7WDJ8t5Gliw7iD
cf/34M+MftHhWTq8xV2G0zAotxea7qvNMmrnr728qaYvzDYEdRRvbXiPI9Fy
S7B7oJKNXKCmsVZhavtRCezjwxkPYieM5KqvPiGdYG2CRbWwJ83TUUOgrPzV
ro18nCc3YZLd4FSE2P/z77/MegPe/EUKKzpyOe5qKWSe8QnuURWhry+h29pI
M9FWPmXEN5H8bzJQt6CktcxaClD1Z90dwJXWNUdM6QW8VFn3GjJxx1HaoE52
7MBhGnY9wu2rexDaR+U1AvDKHL0i+2PNqy8YaqxrLHJbMlWwRLU6dq8Iw13A
8rlkg1u1rYQbS7/g+7/EoYokBH+fa/su3YrZndVZtB3WLhFcAEm73IXPhgHC
aV+b/EJJKbFtjnCUwimv9AUG+6BvyxfrzwBvnlDM/7zNJrnJdmwwFR0JIaJ9
PpAl6JBnztj1UG8QhgmOAfelg+hi6O2waPj+ifDhAve1oSrqHds/sVT53Gox
j7f5LfTYFMDJnNPCdGdtqsJUNzEK/gjRjfD60l1nUJnI9hkllIWPAAvT1euI
SwzVaUHWqrAfNWFzcJd7Q9xpgTd18jW5KlUwlB3EuQHAIAwBrlPm4nGkFxCA
027+g/WDPSvOCquWZkjegjP9sO0gkhrXKk3Pkoz7HsuyFIZ08q1OL6dJamOi
2DYriq2HYWoMEXvNR2F4mj75hckoUIvtO13lqrlilbDdM32k5IaX7v+vWhQR
TxZasGmt/tIq2lT7IsPfjZpsUwPVxmXxXbxLosvtLdrslJUF1HomibkuNGmK
jYENKinIKnh8WXCRpxG4/gmFtDB3bP32MDqT003iAvqIKoAKgCfIr8oNLuql
KzgYhzmixvLW3EFeWyp726hC4yvfpzIoppRe4WQyH8WILJZHq0ztL6f512r6
c0cuMDEAfyvhvmRAaj+aeCfOXHeP/ySZXbqGSHZwEErFkWOTyJiKwRIWBluj
rT+bbEs+DJi0K2i6EmRn4e+bTTDEGjdPALPsTW7UxleDD015+Beo+oplBtEy
WRbhS7QDo+fyJpDyalhglWkvtixV7q6ePpwQN3mj0a269KGu9+sPDjqQ3lVr
md0XmpUwRSQuHCIYZu8PBFYxXM19SQRUjBfsqJZANLoUpGy+H0OC/5wjRIcu
AZvfCYu/yj1nZHj+mG8TvvctaoRf6yXJC4ilOU7McyYDuhEu39dIJjWkppzw
yf32vH+bLKAJYfkyeIUkeJs8YI60jt4gEkubwqHHKm+eLc6/Noh4xaZWDJFN
yFoQVTqtFRoGOuZJfRcfBLmELWBOWSc/UztYJpNomYZFG5It7yHogtdL7f4l
fM8I63siMVK5YmpDuAHdV5R4xBLWAzcZ7ohj5HLmYvSFqHfYcVNJIRq8QIBH
K850A3yFF66g1uGEXt8yUjInvTLLi0aP2YOMQ+zaoIE05+aYKvQ8EFTjL2z1
KKnuv8NTWH6XGptoyRKvFNffLc93gJJIgiz1YwKHvs6qZ/pzfO0XoPuhC0Uz
cfFFA9N+E2CDMChQ1MYPgYvMNZ9IqfWjVUHoYmyzbvI2mcEaKwBGrB+ohlwj
O+Udw/aKgQyVWI8MLA1KvjwYFyjdqZb5UUUkTTBQkqQ8YtlY3xlhZ6E2et2I
t/Ds43FkddiuXNXPUMnqT11S2F6Qnb5JNzeH33jlmLtepbMOQkL1g9kiibgW
Yy7yAtUo14UCjvPAmrjGUfCGWEbNy0UvnhtNr620kwSj6dcbDW827H1Ykj+/
8NsHZMRwCLbOwqVHz9p3wWxGvWZVNyL4QUt1ivnKu20B1DB0sFt75k/nYta/
IwpD3P/rWZKIsmNnkp08Iyy8do4f5Wfm1vCV+DTYZENN544S9q9WQYEOlgEN
IchS3NlRTzD7+TyAic9TeRH57Pc1WyM3ccgimlllLsRRQNKwbz5R6WeS9kwf
VF9U2wOHsoZorQGztSRvdMET/6Rmw6udSM/2x/euy01JuQztCPt8LyFM0vSX
/s0uAatzUF7RLWfghCuwQeV+JE8A7TkhKAb8QulgSodzB72rqnYWJqo/y1/o
vFJi99brPspkPs+dKLyBGb2YQ6xYaY/hnlz+UnvwNJbZHHjp73Qa6eKfjdZR
3LdpjeTa09/IImNxIyRUNfqxW/tQOMg5RbZSq/y7GDUS1pM53v/lurS9+F1p
WvZuFqZDgCU+gz6qEG0d/WBsOz/nhGey8W/5gALLLJW6qQUUAptbAQHTRlXx
ZUam0wjiYkKa1vieH/0BxtUC64e3PUk9JGbruB+5mI8/c9KLWK4kxrChFCzn
DGVLfntyXtYWd4gR+KxO+K7ZAhNTTGONbI9JIet6+XvekMsEex+vcN2ETWN4
YidIk4RWriaZJGghXAYi13sEGyiUuyDgOM7qM9rGRAX9e0CJHkQ2x56h64nD
imlCOooXGtF/xW3qwH8ICRo6LyslsY4BKHYOWkfoEzY4128M0jd6BPcymU6k
D+kdu/s0J/NxcSBKre7UGBOhSH/VssSQj/QX0sY4mIJpaq1HsO6R7kGnfkCH
ZOI4JzLSOiXsPcr4KhL3svMbnn3/YtVY4+ZC/qlx1KzfjV0Cnc9ghNoWxZSc
jqpJotlxAaj9h65OJ3LlfLPVR74NbcaiWFuo2x8j5RLoSzJw7n8YLebVPt9d
kMeSReG7fOnxb/1UNq9uAa8DmTqRIwdTzEkKmUgwA7xsqg6JvWBsBVb8tzsU
wjGslPSScMZERy/KJS8GZMOggnxJ5VPR2T7Ys9ha2MBT0C28BRmkq6r6Ehj9
oGjp1UMR1L7KAvU5+gEgobosd9+Cjl/L13gAC5GGnCgHux/dXy5fmgoZdmPw
q3gmOR2V+DTkgKp+q2PbK5SX2rzH1fU1VOtAjAIjnSRjGclvVL8QhS7gD4iD
pDa3K2IBQ22UbORuNE9NLW45c6Gp+mXEOlDfkTYAZWPSBh7rFqRo4pa7AZRa
qaMjWBDDpX+Rsu+tU0VK3gCClH+Fjd55q8S/wDlbggeVuRLSL5GZDvrkplii
6MftXRHcQV6MyA4fzptKWjrjO/JkkPFS9HduXyvPPsV8hYCIfZ0GHJpuU9D3
g4A7QIw9tyOa7bN72Wlu0IwJqMqOfDuy5eOtmGSOQd1ZgppeLq2lRogNaPRA
fNTeWihWp2OuzZ6+riTHv47sqgdiv9qfbEffHWYWyzDC392KW8AnCVyPpK4h
ueE7KI73idOdI9Kna+Va9NLGxvr4bpvEAPtIePX3GrVqTdXXPtEK5oz8C0s0
uuv0xquZrmL3g3YL5+OINy7JW2JuTW+a3ggI4GqqYIf+qSSQyPojgYQVDJjw
dUBieUlAD/vK9cQ67ef8BDIhft/QjnHzpLprtr4mVnFGkvRckFXBWXGpRxun
Cn7dJynafzFhMeUzTMf5TOe3CU8oOlnBB2IrDWEwiz/HHRbOw5M1AQBnt3Fu
0QdtG19wSnQxUXjoozOLRgHh6vzknO1kSAasKpSlDxWat7RPOsJ4pHCgPFbt
qKNd8qyWQYMX/EOCgnnig2GS8m363FLCpdSP6phALGOVtfpuHTV1dGj2+Mo1
Ni17NiTkLvCsTwSr6hD8HGwo8i/DiEir2IpBWytgNXO5FOnPJB4venC8u3CG
cdguSXo0uTwzFyUhYum84VZyalfXO9pUYZphqIwmGrxpFh2evLps9ZDrkDLT
dzwXgHNyJ+pbw+c3rEgANRNFYGmuz0MeJHLhfsQO7HwEAQa+plakViTH7G/s
vuJJCnfusRSB2HS3VFp4pKMrBAOrV41eNA1BLT8l6Oc8ZU0l++UEkt+vYohL
Q1NmB3XvZ61rG8+GfEPSq7FKE9gkKToyWjq3zlB0cOKxn13TgHvLWtffgpYu
XA2loST971z7QyAuvjPoiOqErO719tsysLvdgK4WIVB0U7mi/A78y18LjlUa
Do9PRz3ZnoQ7RVJq1IRdqT69lQp4qH+PtsR9h5Ei0FVvCpfRV4XD1YJd2xWw
yqBNxMmaR8IDfE4sNjyvT8lI2hyo9Q/1HhgIPKQf/Uy5OVG983pKDZ2RUQGc
eWrogPTtV5C+klZTc1Ta8Rg+KFIS8DI3YE+cN0yKodplec+vmLC7YAE1rTg0
4kzbdFs7USbTgqvZdLV4EGsG3rErOQypHLyy7ko6403sPDqHPkOLh0jgbkWs
+SKMUJEaThwf5V33e//95W5AvpAZZHFn2sdVQmMXC0mLoG+AjB9+gnUvpZGG
1lk4mJNLCBxslixVucp5szhde7FURyzsqobAxA01wus4dv2v9+oDqx4LGctN
uvPV0/IoTr4Jvq/e91xU1gLqpnA0DOdyrPQT8wo6m6XCwRXllDj9SdwoK7l+
SNHharjV6tyJI7ZKlTXpIL6uJlZFvwqAAWGY/Z7LMxXw63psDSjFz5Btutbj
NtUuhVqrUOvUtvVd42V6Ahl0Wxhl6f16ltIR1WS0PmJEj7n0aHbBFcasKLKL
IAok+bK3qlFXk7RKH/jyDEam3uET8SSb9yrr/zhoX3XhiG0ZuQ3IuER4fg0j
+Xa0whovoYQtFwsOzujTKRaEX2tG8uVW6oXf3ikhOBvnQzUIIOWWfodEmCJI
ArNeMpieS6haR9gPWc6sBE4E0bNVWdq2v/o4/M072BuIlVxdwZO+3JBg/wRG
vnTPidsLRnfNtYSJL87wn23+1d+Aqi81TjB+Jvz31K47laL5hlfH6RDI3kXC
kOeR76Phspo4cmNv2wVpMSADTkkn+dO+khEikG9l7hD+HC/Wt+077rY9qpRv
MltU41mdvNw7s0Yf0S5le0IBHSmj8qewqdUdqxaIijYI1nndpHEMakPTrJUy
1pMU1dzInwJQoj69v+sNLaRIR5yRU7HwBQgyenTWZJK5gFEdGGKFv3YOBZvR
Gw8qm5JY7JTY0irKR+UiSnFtu5GN2Fwkd9O4CgYVkeM/BRyEYqnvK3sTUIN/
ZfAqCBZXuBTdiNPZ/MIucSwRAGrYtLQKCpB8IqieL/+qxy2HI4GcEbNGi8bS
V68OgMGjFKWHzLu4r43S+5JGF0q62Y6I/4HajKvhe3/mIlOrDVtmmVDOUXtA
Qe5nvF59z8s/b4dKsfONSdiExPX8Ki9Qlq+dFyYIR6d5LcZQEqZQqJ+Rhg0C
SP7Qo59I04+x8Dbzjhrj4+BGHRV2Lcn/RL5MmZZDIae6X+9K8fYZcQQcvlSu
E/iqBpGGKyz2E7pSXKom60HuaEk495W1YFTy8wY+ibNl2CfgR5VHluGbvsXS
IR2G1olJ9Ebziq43CacGTAUgiI75Df/n/13F1lHODwxslrAi9o2lMp1t+Jdn
anpQsW84uAFIwbJR+AUIVers573u+5O63CZpM0uJkl2H4co8r9xgVCDV7jRC
607RsVye11XrpMOEZFkO6OrY14mlOPLsQXFmGOl2sN5mj9j6A6f2Ibheimvw
/64xNXvZCZUrAoNs2qIvnTFsM9fM5445phYybwnlWMoRXnsAWP/7NABKjlOs
yKUNEBQ8ON0VV7Tezyw5j4ApF+EeSmvAJBT33AfMOhhQNcYBp36Nqw0z0lHL
4Cyi+huu5AWj3zlXFoBlOY4xpAZpBU1D86TMZjaEe9Q1UqezoaMrrwHe2LAs
/Zl320OjJ6twwum3qgd3lMvNKCrugOJxTRt36VL9fcjDnfrurDSsDjR/qPOi
Vyrbcko3QRTRx+gZtH2ZfsyxsQVQ7QoHmTZxPR42j3jPniz0I3QCnQ577PmJ
uRW7HSy74OSYkm1oIsReAGXBToq5RTZMLib7EyuLR3hIlMw1tgHXICUrOWrc
OKXK+fusVHzEgpTZUAfel9D0iMbBnRUbXH0ut0CWNnl0drg4MMimQUqqRYfo
FQ8Pms3509EvGPgA7WBJa8J9+8xbMR6g4aK4e4pkT7CMr/q5CWHJQvplpH0f
Z+41PYUqFbpV08eVXrGOP3j/L38/A4foFtcW5Ucwr7txiZWHrFukmibQNalw
DKStNWGcpkRR1dLW1+/WaObnqYzlXjYJItXoBLegxqqaD2kmRzKCDvMVyi6a
/nOMFoeYXE+WxLVFXls7oiqkKWBkDB4q5CPIl4HCq7905JSrxoT1v9iZ7V9G
2euUhtC0rrwckDPgcnyqHGDo7WAlwgQ11j2DvGQlMmgTeed4cKD2VL+M3AK2
NOSYRSUDlqHZE3KcIu+cyjCgc1h8mxb/9cp4nSKXp2SsU5r5tWiO8b7vT0Si
07XwpVd1BZvbITueMsIrxOba7xkDWZV7TeqK0DBor3SJeq7CjPBrhTaRqXTp
rJXalGSaipWXF45AdxdJMsZgWPTmEGMmU29pUuJNgy8CG46ix5Haj5kpsVHY
UALt4UYnzcnly7q7ZUXLfJTy9hlyp/TL8+90ckzwBBLFiBzGn0XLinS5L5F/
0zRnKaij9j2JmD+/EC32nU45JetwZir0mdy7Kude5LduGUIacWkhUxA4ikDt
ei1ig0eaPAt4i97Ql0rJjBbSsZ0zXt1dPjx2Ms/QhLCAtklytoF3PWECGWdL
S8J1RdHmLzlaRv+LZ34HRJIG9D6L2YJYqxQ8HAzoy+EPBccD6laIl34o5U0i
DspFOmFs1y+qEBhBpcPV5So15AAhwwEss11ltk9OxlIyyGKIw35btwQFo+Dh
xbkSAed9LDBB1iuWV6IvlbSVJnimGinLP7DuO4XKQTPhJP9KaPHjXw5DncrX
6knCeik1mykTg+chf9qbbL1NqEvTvEMAHG8oJq4mNn5W4gdFT1RR9DMA/RxC
2YI6WtAn2UmcQ27SAxGiQe7zlsP1UbAb4hcwgzK85yKhIQuSWyhUL2HEe2rM
mw1ASoyp7ovtnjniCR+f+A/LpF2M0fflrUFxtKj9uZIgedGBbGCQrhmBBAiV
nvw8p+BMbWwi7nAmXJHKUVIfqeDe3zdXsen2uBYrEUdEJMSVzHvQkFP1Fm2S
Pkq1t+E1Y8tqAMFTlvvZA5MdRhJpOMqj6D+8CkTGCwaxH6rF4IFHvvvp3WGm
8LcGAz2EsNZ4ubnuvAUo7NQ390Fb3ZqxPd7L6tQBnbPCydVAXjrbsy0KwvR3
Bz1h9Wpqaql+37gcdyWd1sSv8iY0pk11bimq5bugIrenLcKxLmi6kp8+70CL
xgZgOwGhUBp/KqmmdnDPyZfro2fQ0MLXRvewzYvPPKromKaJ2iVB9aiqq09r
7mzIuxJoolCOeC6Shg2kUeIVBOUYjqr9MQ8F58HDF3Q3BCL5Tnwa8VemTo/d
uwMGU9RoF7CkdPFpubUHR9ALAifuHWNy/ts2ss/7MnVwLjy4uyhAB1hU4A5G
6eklOnQH6tTU9ohxjvZVznyt70q0OlnuaL1b/i7bkzG7EDspwGJXm2cKT7Vm
CkmOhL0Mw/aUOCvBXh9hTqYiNwoNRf+U4Qk/psTZuWwXXWdWX94KU/E0Fd+A
Ohw5FZNTH6L9ya1mCJjGDcaIHMIsOQiyCEtMmf4qS7QcwHQTHNQE7TL06+Av
Rilq+I6+uuNLDfce2az6futMZBiqHz1egS1tIRWzUV2BZQHHfu8P4GCy8JQR
nn6McSdgAzyJWwVAFCsfHDLCyKJDoVI9XMdq9aL+OrIO7DQTyivatYnmThGG
rMKI6FQJ8EVYNgPnHUb4PSfglNkoa4Jkm37kw6qxL81B1MzYBhfk6+FS/yzi
aGRk+Pr3zFiFUQe3USSVrx/SZd63yx3+MNMYO7h6TnO2o6+mkM1g36lL//of
AZgi2wBrzjNn/r3ZU5w3fhkO4Cdxme5exvLayZh63pBg+2zmK44nqnZgl0U4
D8043f61LIkVqa3xqKKzQVFy/Nlx3Z3dGZwsTxYKJGKRCkLw80Yk83vowK++
cuUtPlnTgo9c9vnrXLyGhZbC8VCIspESX1HkWwKegs7WD5j46tKz07zu/ryn
whCqly2uvy1fBorRB7iTglw2UMGk7LuvtImOQD/w8+1KP52w3yRB117usgW5
BoURVNnxWtJM2K2gtDwCzpcNXyv+goZcv36mj/8mryg4p1cNKi/OVZbmVlX4
UHjFp4nSL0KQogZKAQmZAB2eunr5jGBA9+QCFKIeVNfVxsSGwG+GU0qBHppb
i5Twap7GlWBZsI72t/w707+08IEvncVM8MnjW2TtwvnnYDwYsjC+eXmcsgYL
h6rbKAZSc2DV4Szo8dwqsLCAoPyPNtsvoOumPt2X5ki6lPxTFMo3bQ8jI5GH
o6vK9LJh4cHLIspikXcA0xgHhNYNxcc/cjJbLwlCFMxgPVlNTiEFAr/Wu70F
/xMYqQGHunC43Tq/m0ZiLELLYOGUv3ExF1FtxfFVaafbZQ5Dw5o6+h8WVK7Q
FXNaSbiz1Ag1dq2wpyan52Pxe8LT18Wy0NG9AIaJrY4rjfvaY9S2ANR55LMP
Ub2IicGhsBPcE96kSS+OeOq/uUjoOqbxYVrVDXLxMRjNUOEh2PZow8Dj7lK/
GQTX8cqRVOhBORIM5gskS/OHAj9i9xcN7+IMDXt0HikzFPKZKXkNaLyg2vcy
0HxNQaqvEGo7Ji5gGaitIiRtXZumcy53t3o3+ZYlAnxSp48ms0y/84bkrMW8
oSfXcJpum/lN9PcN9m7pqRz4c1RlsS7EY14SIQ8gjSPCexG6LKWW3mAytApI
Th0CrbUhYgtM7tU4b035v5Uyt6wNR8e9RHKayeHH3CDRyDC6Wsm90gkYmVR2
Mejcl7kLWNw+BdHuiS8x6hsZ0D7GmzTq7zF4uHK3gokWIU3S2b4uYxmzlgXJ
2sWcFuekR87VJYiTAnTwrFTTNfz8jxMsH4mhLDyQpjwZFODv7vJYmg0l3+4v
eM44diJTEkLHPIRijvk7Bpnsmx4s9yLig7EE1UdBvkw4pScsUqbfzcesMH3G
y187itE5YdGq/8Do1lSINLBscLlOzC+QgUQmOUWBuv02FtOuK88uEVfeTJbR
6M4Mb7PeGxNCitCZgSAo/17Y1ySJCVcWflh9EmNxWI4U1Oag9AceByhtmtos
hUZUTOKrAXw1cYQ3+TDCr4V1b8GT9Y+YgwRwkp+dEPNv97W6wGuYQX4FmX/Y
wsHKiGpcSYcW0o78AtX/wo9xBxpl0g499HT/5L41L4U8eGp0RdaNW+IdNSZs
bt/lrkIrLGGUyVi7p+aZ9Y0BXfvjv3zWQtCX0Rh7GdcfydPaygDsK1pwwZp9
uNj6QUXB3TMLhjnSAmGb95IWjZCkotu37j4/JU6/ooOWpVt71sPxHSLZlWU5
kidQbU56FBseouh6X2Rdjk+llweoHjwwuISSD9Oab9h2j/+Ks4uQBZVrGBXa
Mv3uodN8Qy63rnbhfHpoqNoG3UcVlAz/KksEpg/VlLTWw64wH5zjnEJ/y+EE
41fQ7ez6wmk8Jmq4aw0XJ00F1dEMD6ZwdnAOGWkrRkYFK0KY7ryG7CeatXd2
I7jPT28MLechhTvhkP/jOvFvk9tKfUJIzU6NFmuPwAdvgOJg0Xc+Ka8H8qRE
RvUYtTLJ9HliXgYaTnPZ+onFr9tAk/S6IqhpjA3zVZLPuDUntU8ZcsFJ+vJm
TaL5oeQ4o0yDcUH8JWQcxKBb7N+ern5yoTLP3HiEvpuMcsvTiCeDt7w053WH
8YX7KZvjMg0H49UdnMgt2ICdluowBsZBylI8BZ/IbvLxhRcvYYitxczyW+HZ
iuEnbtpYf5MOUkdy33ckmD+eiZNUQVRm545Naw0GnpITckM74GFLRPJqOrM7
pLhFEzUlGf617cs3IAEBN+fUy7GByzUQUQPzlNwnWYSOgKV2c7Sr27ihnwO1
b6tNOd5TogZYOYZ72sxu41mJ5adAAsH7o0cRqfZsAlCJ688fIxRp5oJgxUwo
R4Sqp8ovEdlnsqxzE2P7E3YCCx8P7qqefrDkPy6kqto+HPePFnAWNltxGMD+
CLOkRSiyh/paZuADgcOhxgsRuxB6274hQpuxIlchtEm5TJWZZCbTvNMUSxWp
nw5VGqMVeQndaIdXE4EEYGNY8yTOVFr/d44LHmBqMR7Oz+8hVbBKy+7oGVSE
+n7eh2vX8VRHsj8OmUItki+h2ubHQR2bQHtaLxtyXts/hOg1WBFIxSYTXYvd
UdD4tO1IPTsG1FPfi5dc4zOq/DOoE10smALGuuc+R0Lh5yh0EKv3ldFk3SEi
Xmh/boZt5fRFdK5heWzLrCka9McBF4pZeHbmnNV/lAI+/2eaH9FMOZHrE0Cg
DICJzqqpkyjSoSjFShTmOcYoPnKusgw9GS/3s5F2LHqsMBsfLg5dTsxfRHnu
f86qhXOZxuOS+gsb5+wEvd6x+tLvmdv0HBgQuIk4tgBA38qqn8NJtWs+To0M
BL1eUYn+3EBWC2/XsiFMMjX5Cf1wKC/csyaNvSDOCZQnY7XzPbiVbNXNxewo
n/KIcO9a3y5eIcGsXKB/lszPgeH1Yf6BImc0MfMC2r7gBojZSN2fbAXbVc/v
aXT+Y3uNWcTo0v5uoJsr2wtn8Ut1vrKOm/3FRDKbe47gWGM2ZXyYHTRR8/pF
vEk7GD967c6H72meF/5VAT+U6NZEunaYZjECArk6JGeuGHvd/NdxbEcFU5UJ
UtyJfKnszPIyIsHgsdcwY07PXNLl9hp6+0iFZhogZdDcJEQypsPRpNg3rFYl
MgkAjxF+qU4vBbDwMC+b+2uMFGyLZs8uHcY61Htrl8czXDZoWtKm8p4yyXtK
3pQ3kalIw3arkSNL81spUUaN9pw7l3WttWpH6j5NmNj20CVXcKurnIW1/Jvs
Es2MSt0EiUGIR2IQHlFvm94JQspx6t2JM+GCvnFwrvVdvf7xHn+Yr24dKOMz
CYyg4iil1WkDJhW86wuM1G+cGISUD1OACuS3U8X3fOAabBphp/AJesVuu3kT
b8nzkJ2DHWqsG1WpypHVWf9ZUVgHCMJL7nCNw00DjM+qKdYE2MyqzJf/6D0Z
xlxqie+Gte8duVgOhZsHaDWk9SmtyBD0e7v3NFFfQacAhtrtPZMJhKL8FnV5
B6Q4MSTCDCYKaqjWO/anA40pposiuDlZHzR7vltN5CKDPji4cRkZ79mGUtMK
yCwVaOSHwmLVCJIN27j91G5q3qdT+y96f3jGm7uSVcWuOzTRlCkcMn/R/Teq
FXH+2ALFwd+gHxjx7sI6nEN+u59R8wyXvZqlmHC96t7Y5dZ/X9KvqLiEMBZS
2JcEOBRlSr86pdR7DPUOntOh9a4+vwT/QSqQosLOSd6FV4SMpYpRc3EVWFOy
DD3P4v5FktwJHfWeEM5sPlLFyYIXWY7xFWP9i8RcDf3apOlZNxD/AW6aiAad
WKc21MjYYVLXOY46hUXTTtT2tKuhwQ2EZdovp+xKdtzlD1cv37dxOowQy3Md
WLLfMRYQNXFmQGqC4G+rJeRfmUYQYzAMhAie2DZE76nlLpV+LsJkXXGHSfW2
58pXzX9fiJ/Kv2LcXzsGOMPQpDXd/tzLhdjPQQV2deyz8bunbT0ACtR994Ga
lzFgJ3YuDeMXrwYWAgptrmjAOdDTFursbD3pnEg7DDCe4TBH0QEbrzLu+UMb
n0zcTNKvg2YHICNDhrVrYANttrndBj+Uc1cwXkXjjtiDVmBPlBmjKoJTAtu7
FG6d4zJIVZM60MtGMM8RFobpt4zoO+VSrG5Opjjqu6C7pre5PNXYNN9w5LTu
zyri+qpEdtun+g5YxxgUFl5/6c327I11O8UcAhdNuw8LSEn/qJWgkhKu299N
j8DmsSCuziF7t5yu3bB0lwg2Tlj6+5thdDaSfH5oVc/GyEizZ/wvEyff5E1d
6XHlVoeQgZyYiUg/P3pMds2o8k7xFkpuRB0qUxTUgIbSvXSrsZUCJAci+suf
XhiLgluC3iUbBFGhjANJvlF5ieiy88tQkGpTjZHthctvlQSi5nGlTioIShrW
zCQAhjb14ybUCTUGYJnh4YpsVf8bw9wZ84NDZfJPPy7xmDfO6B1Ss/RsoAKV
JiE++MorVNg1wzs9IcJwJTclJlZEMi7RGSUPK3etghg8KYE3J/nG4JuQv14l
yGdQJEWphThkBgsWpmUQn0IOcwA3+qjWiKzGpJDE+0fREaifGUckvFUigmxF
NfteZruEgBX+UUi9iw2coPXH7scExg0+x2s/9qJ8C/m2mVMElxblyMuWyk6q
n6C32EYh3keXsDGK5qJN3egumG+N/VU54ZgrmMVywJN3GEwmcj/X78IVtGqx
u0bleXqEaibVpPGwhAC3AAw8tIbmSLmXZR4dSzdTnW9US+O77AsAEQTojYzR
apVsn8bXOOhdFL6nhdCHh1u1SPQXV6tKmM81ykGlXwtQqg1pa9lzIRWPTplp
EonC/xCqYC23uh80N0UYAOqRsoIm5OrDMSLwEuJAjcEf4I9CYe/vYvzvnXN/
Yte01Xk+i6Ce9KC6ptqU1gGuEO17/wiAheGBt88dHZChxLaNFVa+1vQ3QBFY
rM98lO5MmhMT5znJd7m5B9mNHRNL/AKgorM2p9o1Xp9SLNA/7Q6v2LqYrjEz
/BmXyIXvugvg0UQGez1i/jRxfJsgeA0xGppNIwRYC+NWUIr0lckVJp7zh9Xc
h7y876yA+thnKHUyikWd02Nu+J4KBjSq0Ksz4rslVKhPlTR+BKrerjE9uViE
tDMiuGDL6CWHtHLCTYdRtsYkeYA46QwE5eZ8WR/LZhy9KaeUA3BbiC7l3jZR
DxDxwtDRYnyP35KYQ7eFnstICteeZMI44nFzHeORxUiUw9i2JIFTVHRo2d0z
0cROx8vW+0vuf+iVKnLQJOcJUJE3DBysM9HdP9fHrB9IFvAY1z0SwaHAmN0i
lsusINOUJ/mJx+geEEcp3UB6okvaXdpsEL0rrhXdlm0UNLs33EacOilCu88W
VlP9ZQYF+wDNKAFLika5HAqie7JkYIB334bU/TYmGhmqsW+IdTVdVCkOjO8a
mdp8TFDyPyuzRTHO/2ck1ocFNW2BWuD7jwZKU6W4m4dlwtxwsUo3dFyEiUED
HxPBWUBSnKXV1TOg+hsGajDCY8RLKuexxNS95jkNLZ1omPtyq5xM/jNit6VI
tx262f36NVIPv3ou7Krf+hNvjxPkQWREf0dMN/FDoBiZY56E6I09HesjVKuV
ITTXaggohhZvtAehclcevPUIdP3fmirqVrBynopT+smCV6+NhuxVxJtkuUdI
kGcsMZEubgDuxl4nGOwP126Jw4GucWGHDpQbdKOeqxYHaa1JWMO5uF8jgOwt
FOGTxI0gFwbJYBcC+vZaobFXsSLdmIdhwszLhBsvEIkdUB7onCGEeykfKMhl
fcMZzUhxrq0iTRqZfO9jaEomaKk+WTrV1au3hgDm98xcYPv5c0GYUq9JmGd8
q+EOhLrgu0HtxrjwUqndovpOhFv01JsMOq7T7Rn6Xferdx3iOFttRP8Hl0KG
zGA3yCdQGMK8PFV+x/r+TjcRkODqsb77r03V+DUcJeDAO6HgAH7DgRZeAqt0
HaxyPNwKClLwJDyfb2o+N5lp748fbK5UnK30HQE4qLouZEpM9xA+LO70rCBf
Fq9nUIU0hKHtUn3/naGYSALIzpHhGEuut8NhfLdPSESQ7QD2QFDv2TM9tZ0O
G3aGdTPrMOtoCuMs3J2GEIJ2vT68H3ANJicudz9AXjUKWZLWHfeECZw7IXFH
B/JPqB8N48L867KyzvJ5iM9qYElc0wJ6nWWruDYh/Kd1IcmJcyGnljSbcZA4
jyTHB3jzLeUNVkU2TxG52YmH3L0ZMoOFK/UJ0N4zzbhM7ARGx0vOy/clHRmm
2U5gq8B01GJMCeiPFty62x77tFSnZs81riJXADjr+TU3ZQ21Mom4SjRFH+kK
dgzQl7o7C8dG+uvrsAA3L9kMTw733pd1Ak20HaYHupEKER++i5g93WYk+YfI
taVt3BZBn+q1DlJeFB2NsHb8Xm0ym1Ko9Nn+dHuWL35aFIzRdBDAiaf/jNEA
ondjItusiyT9YFC8HbFOqcpBKzSSkfn86KtSO3pQdHiNFYKd1G3HooZRsR7W
RLfFPLmXx6KATo4XElWyJXSjfo2EYdRWcq5Pee87ifVvfg8u7JkGUmNcJaLr
RolCSLMlZl4HoZDvw3dcNsHMxjxmzsE/e8eZF5YsR9yPehj3wpeUHFNKAZSK
9wPFI95tdqrNOQu9KGTFvUNz99Gl3/zUIWRb/fT7kcahO7zn8+f/X1e1a9fo
1K7CoGkY4EU0Xs7aoTrXjOIw2o/WTMUheVhVnHfQzoV4LLiCDSpWdy1NgsUL
NXsq3+wQAQcNsAAFL3ah20wqvFL00zb7AKS6h4Lc7wD/JzwHMXXoPf6UOF4o
43+7I9GXsu6GsgOBC0BeohfnxE61xhWSppZzs6CafF1I+xEAGsNQXoleGM50
CbNmE1mKXQgSEf7zW4QvUxQ40ycmDK5/i+4PA3mtJrNaeMREqletpbQMegpm
3SX2XYJ6y0tbpKBkC8rjisxnmJXiIzPOqbHC+mlIv2yMUfyu7om/+cETVyhW
KOWjpQNvRt2OTHhnbhFQqCfLjyLuXcabzlqwB1EVaeqi9/jnBdQ519Ies+Nc
Xx6HHzuEPA6BnUF7WPZ35j6/RI84w/ZuPg6KYL9OCIQMEoDGQBOq5Idgsu70
FXk/PQESUckVMC4+b4BhCMo8O3SMCK/mBMeXWyhaW9GH77blkcToD1hBttKC
AQx8IPls0sObYeIV26I/pKhZuq/ICOCFWp3EVwOWuvAzzY2wVXDSVumA35wt
48E0Khyu6j2j/apNtGMaXhQHzsFyeCpCjHK3OVhxlJyy5/p56672ea6LuHoM
r/cvGunqaeaj0XaY43Tav8FOEmJ/Z/5e/dFgDN1Ed51rYq89RfE23s9UVrQx
Hy9daatc4Rl7A8SjA4kIJ0GYAR6WIzTk+CxnBK8SiAT7Nq1QQuGQ8nzYnDrY
+EUvASeMa1mb9XULjdvlL7u/bkpG0GQYQCq9cxqVw8wPjrJ4QqBa5sjMCs5Z
R2NB+qtdCxr12XYRhO4vMU+QeVoZSWggRIQWiAvFFIyq5tGG0BmYefBt51Fh
Db0KSF7FTD83lDz503WKWKHfUrxurlVs2ucdmVHfEMk5UXEq+jGbiYJKMcpZ
0aErZ5ovnUXyD4sSUQ+PhvhVyr1Z5586joFPv8ERbC4hz5xWYF9Hr3AbojwB
L0dzf7LEkHZTx6ghAv8IxrsII34HpxUTk09nTRGLvOaVQ5f9CT4pdWr8fODN
GIBVkqv+K5NYTsP6Zhi09RVTm/cLcmcpwi6fvOyXRa5Eq6bXG4cOvaqEywqj
RnfKNCnjPqlACcGiMBw9BQOkPqKlhrm2+nwzhToCkcwvWm2e+4aXbzk46QeO
6n5LXtm7IjD3qTyHiQSs0468KLPfkkLIsggVnm6B4ij6pORiB6UTabAMfmHo
2CGnj48fmJWPY6Tz3+UXyzEy13K0pKZkNNF3Xxkc6IwQvQcQahtqAeoDPez4
9I63UNnQzWxnt/ivx94I/2P+tIZjrTdRk0NTp7O6gRLd1NVn1ttRBPu0x0p5
WtL5Dt+c29dbc+JvE3Eh4//wtdM74S4+iWBdFEMvjEW3FUep4ur3ufgiFjSS
Cmz69D1n1yGjGB0mf7/b/tDwIpGNLHaCh0CsOgvzrwAokbzNYh9K8kdtYZwI
7RM1u0HTn9fHaQ97hBhJNcDA2I8dT/PA8S97nPy8t2vdgrUZfWAKKpkv8lm6
MMhrqnzowAUu0BBIxNwDEvET/ain8149pMTYAagvNIFklSRzCEuyCvvr8Fd0
/F0HMPfHO3Q2QkZpvp+jBFVu6SO/lu28ovjLr5xmYZnaMiCM2g9lisBJDOdB
+baHV/9n4XoP36j/uvDDodYMvYyLtO7Oo18WdMi9/kCvrPmEqaV6Z6C30Zfi
E+fA6Z+J4d9i5lBKHIspu+1KCUYFp6JfwbrChPFaKFgUbThb2pg9czKjvc1C
2QVKQOPFGfP65fkSV+XcjHeAnjlsHRFnBsSEJqSBMukgv2ZKiLFA8dzE65FC
rJe9+6CxtjiM7Wh+WPjawXhJpV0W1C1dSd+h+2W0+JoHSAJ8V/j9CwUQ6Jmc
TYEuAavdI6QrNc38iCMTvbRC4kE4cOuruXMC7d4tcXRApc7XTuGJlwCxvzxm
BF0iDV2SO0oM3r7uQlJZmP5ZsMwGDn0WnpKmiVMgLwtHaZYtMio1JLqfy6eT
YJ53V0ql0Eb72V4enMZIv8JdnHikIv42UgrxuCSosfrpQVTgHHfIR3QBuQOS
grwThlHBB4Y6u2+FL2I1/osyGG9hr//116A1hGMKh2H73oNV4nhEWC4f+lFf
DzRtLosP6u78gUl+QPDtHb6Nknr0avrwpcdQOL7ifyKqPRirjH4eG8oQhVGb
v+9G1dGAxrV7l7UaJZDgyu4qrJFRfAeW6DUDwXNerYvtZ+M+crQ5x0Soplr2
ct7FeHKGb0gpAvJupepBbgvgToXHzU8d1jD2n8CMPhak465duXr9l2+8mf3B
GYaNxqBE7yGdEv8FRt09g0dA66O9j0P70kfmq1pDqZDz6orYJP4TwXXSzluq
7j3jLCW7YWRd+R4HbYLGxn6wbNUYcyVp3fez5btSEjliE9jQnXsbNaQpsudK
ii+8tK2V0lM4rwO7q5lU+GWrJ0AgdIyNsyiiNbGzNCA99yco44uyzdKEt8wv
Sg5MwTu1dj5+tFaJuRONyei7dm9MFIBC9aounTI1gmcd++1ffOzSTSyqeLrQ
CeAwW8IwIHQ+kOx8uyRmdaKXTenw8z2qru3RQRNQXQPYTclQ8pFGTjzC+mvh
eyqnzHI16hFB1wx+oS3PZqJHb+2uN/cbMVB2B6vlWiAZuVdclEfC0k/9HQ5Z
73DS8qRfHmj4qgvHcSVElV+iVZ8mbCClddRC4CTu56R+VZRQEWXEqmqfhaKo
bciCR8BImiNWGbI4a1t8eCKLSE6msBoemfaY4HJHRhGrz5Iim6EyEcy/mapQ
oKiVASbG3PQMUiUu4uQF6VddVeCCLynTzbT1C7aOyRRWTIFv56irwSqM/CZr
jT7T03tktepa1pRvOpnLivaMW+KVIE/aRIPuafTyc3umKMwbmcvJR1om/0Pk
QXuPm729fvDhqpxJYNM/xQ9uskXX5ITquJwlHu1GWXEurMMNC6somkQiWtfg
tb+5wr2fVZLu2raT3CUwwewx8aiZj/LZ1aPMPyh+TN3MhNTmTyb5YzMu9ngJ
jXa4y8cUszOv5g3hn0I+BnkcoweLDC/WSKflM3BX3Q2k1LsmkClFjJ1G29M2
LKUc44bXO7loMmHGjvxG354LCrtIhX5/die2EbsivSWEX+nX+Pua4JMy2/uK
JBZCdwENeWTpnmb2t44TmkERquA92mKGuUU1R3bAb2BASInjzvgEPlk+eJ03
cBy03MZpVXNjbdQw6VyhdrSV7YU4wl25rPdZRWfIXTwsbl3ttBPMuJQ8cS71
PmnaCkRuEywVC6z1lTlkz/pObyDmpGNXNPc3GwH+yJnYYBCYFpbXCp73qWTa
FqyHPppoEJK8G64YlM2rIAwQybnUkhqrIdb4PZNUqsosSyDVyIz5KOXl6mq/
A0oi28hrCox9SL9Xnb6xHbIRC1+H6aKO1Eh8cJD7Y8IkU5haGGx8oQQlJ6HI
Cm0srcxsXy0EiiweQXiKiag/0bOB8B9upiWDEJYZ5UELjTdRe8oNqDqduah7
UWwFirfUKXBVfDx/zFg1BFVbst0l6A1Z40xZnI8erCvxe1kGSm+AeHJP43v4
b5JU4B/9peD1xZi5XspO5agS577lUeJfohfGXWjpFCrT+D+4J9hLlbSiuLbp
6j8yrPc4TmWTb/JB7yLTsgMVJ45xs7g8Qh9+B88CsAf645YpXQ+RPv2HamPR
KT+f5s24OS2pWIZNodPwFsf691OJ892YGmJKDU+PtCNybv1dVpeAA9+UQ8ha
hUm66LFthEkUE/75l4nnLiys3I/NghqnDWjyicq7SV5erlm7WGL53de8pyXw
gEmXiuSkuoAMPw0gpq99gyobx/Z8S9txlPcCLSOx6gs62HBBmHYHj6Za1A9w
YzVBFN3CtuhCI3fYO9xwyM2HLNuula8aMOcbtiwVAF07htKzx24HSoBtCkHJ
NHcWHF2GGvvr3vrvFPLNZuLLB800JIj5OaPY9mG8jUdEJiSIQ+wh5aoBjzt9
23LJuFsoDpkOcoVsV/RWab3JYQTxXhnVDZnBNWWxvJ6RwjKAkW8d4f2LLIfe
D+6BTYNr1jzsnwSRSO9CbyGH/kmvgU24Hpd1nWb2Qj3F6MGHXesS9ep/uZQ4
bdGfTtRulKnYg7GXz2uMVaXe1dO+KRUeyO3c2MHHXa+XBd3o1Ck2chcxPtGe
ZbDJUp3cUtdUV/7xB5dM+U+xni4BiDUkYon4vWWETJ6UnKWw8UInMvq72lBo
6BxrNwNjpP50P7qg+gTphoS78pE7zNnWgNDUAxToFnFWP+oia2vU1IreBObp
g9/nxnJxXwM+QrQAyMHDKiIbfr3sT3NJ6+Uv8NWKCvflY0NiTHCAkZZEjT55
QsFQpHRtUlh33zxoRO6ags/g9Z1yAUB3ijU2GxBXxVVk8xwTllP8sIIR9ZCP
u37UEFzTid9sDqjYEShvnRbIsLtwsaOk22I/G6EWNFwFtNJi5nUYyylDPZrf
MuPlw5dDv8geXZx8z/yihEGoEMXL1eDMqX8QixawWVwjFaWBuXkjeqjRNNEG
+96BQ9J6e3GaYXdf0Y6gbdflnktP/20ftqLJc4vaXNlYLfDahR1OYOjV/wth
3P7czuXzNMW41qkjVT8DSmQMkuU8RM+JLw1LEbQDmBUALZhilInZ398/Mn6o
6P2U5EBeqr3hbV25EoCWCIMCcdsDN2I2N+gy27k6oHFeVbI8p4tPLSkhnTL4
hWlDEv2xbEfN812E3QHpqUF1fa7GAZRbOwFvsGDc8fGvLAZ9h50k6Pv3W06K
5a4dZbaqqbpVLAzSq7m8HlyXL16IewAr0dRHqcBmYLAf7MEbvcERzEnYt1Mb
UYxFWXmdy0usTGR55xFybmpYKf0D+cxHRA6IqqAnp1yjnUYIhrR+Uhbat+pi
ckERaCgtGHnW8u5B4VSm4HtVEwj6ZHjr1p7zlMUH4caYP8DMVBPyQa1AFgyU
AgsktvpCvfjBnCRvsReo9wZs/NV+MJ8LJaCvPyFetrOvZ238zNdehpJ1KUVz
CDz/lkVayDTsbzc1iE062XlQaOhq5zMt78ETS0wsTlBllGF0G64rrsEru7jS
5c9TIZqvWjuUSkJUaXfw3+CqmBW/WnfGOe7VDWtsbZVV72B0r92Y1OxFn+Pi
xi/te1qxPgYNAKVOMQqhpg9D79KW20nDCdfEy0Z2gobyu5kJn9aKTZrkrMUl
s0JV//8FKL3p2MWPK9sHFEIxrUdDad4R3zBAJMYqpKV+WcuxQmaIqipvElom
ry7az17/6yxwxLnUo6b8Eu5EU8Sk8K5ovs423KNFQxHb6vSAi0X9va3ryYGU
UfKlgNpxcVLMriBwSlXn88ph9cPsbnuO1c27VwXH8dQpbtBDO1GzTE4tFkDb
RMRL9t50TNXSJgNHl++jS+t4DCN94rPitBLoRX6h6u8PvzldRNpSdTtAwTBh
ck4wRc8bXIIldN8vR5zMxtrHoZf0o7TdLcbapAAOyZDHp4k6fGqRSvYCx10y
w92I4zTsOCx8vsMDjcbGf+zYMkRf7Mu6eQcHCS+rfdjc5+rRQjjAPoj2rYkW
LNTFvHjXRQ5FhrKvZaA4sz0oM8WSTDvzoDHy5DXhcwv9GcCugGaOaA3YEmAo
V7bUKYeEf/XP1r28UIiNB973yDvD0YPQ7ckRDA3afc0Zaqj3erWnqugCVZwL
M4WIWyIqvZgx5OlKUNHJrwvgCDg66+EylLhG3Oi/tzBGgccEf36+QQ5htL5J
C3nQ+zOgFBVagnz3omAapcL8XjWg4t6J70ySzR9IMF1QxGOfeiJRozlc8qk7
FoAc8DIGJIQlK4jw0pPu5bHGQ+InqZ4wxjPd0T7GqIrV8wqvHP5zLX4Eq9hB
h3YoXX86t8cuYV10xhveCJCRYUvaUSjvaOy7xsbcy04sWpI98pjtE7xA16mG
5qtl66Qj+qPFTP61o48GsoUJb48cQJ2hwQiLBmQj3NO8nJi3WQrN9bmRlhce
tPgBPhSbf+ImiRHjQUJlW7hImPiy6v37OhUwUfEKDUe4g3uP0y5t7OH0Latw
+2siChzU26KUR708kxxjAAd6i+JET7aGtisi5xKlryovS544sWeeFtCKTxfN
qBxtm7vWjsABSHqv9P6pSYMWbvVJmgP1Wsn1wzY9Xtl0Dqpte5xUrHypgHRz
5LVvC+yfNr7UFi5/QUgmSq5bpP86OeMwk07lbYNYbqrMLYmngaHkwF2xBzaG
sad5uN1SX5JXcj8tX62n38y4Lyp3Mr6T/x2x+NDG4D4XEd9jCgLP9VntJ0p5
HjCpHz3d+KM01m3DD8tecryJ2ensT0+bD7j6gn9yC930TDvTrYr7phpg2Lpz
jVq78AYoyz2iUhrOdqFeDnYpPR7tbQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "9RW93T28GeolckbYRvHffOsKFRFmORm+azyCUYhudrVC3P73ufaBfyRVMCXUVPfCA/gVx4qupGWo2/MTXHrbiqujt9kp6+gvryDIvlW8esKlSeDbKqIxzhLY+DL5yFAjg+mCmTKnMSoiZ9J0N0zgOO806IAkac+OYN9FbEIEFuaO+G41krhhxrcYAZ7qVX+m993ig0jH+TdTkf+bgk6VV++svRquWf4VNDUj099hz6CcwzVsmTX7BBLR7m+pJ6O48Gs9bUPh+XBwnv3eAL5AFt2YbuwpDzAuSbRrRVOgFXpKeR7R3zIbOPrJJ3R4/3ay8ZoJa3G4zzKfkE8b6AYlLD3qHa6HhO2AF3EmmjRKS8HSO26Scn1y9nLikFtMOTIftr8I12rtyoc4dOa7gobGlJs2EkB4TbHE2qgx8H9omOZAYIfushdkeHNdyNwiR4Nd5kKXzqC7/JGlPisrFAnnTZIetfBjvblU600FaTblEWe8AxP5QUna1YSVxYFDXRLaFDhx7xS/yjI8RGGWZZIUeqgbH7OLWF00ZDZIUiVunJFk/uBv9SJH3bP4pcyivp9/DnKrfZRUgxwngyx2F9C2/f6xVX5CVtk7chmJJ14Su+HRmz/xYBQ1zuIIW8/YGpwfQznl98L/Obr+hJHgPxwxFYmxNpnAf3i7yv2QH3Jnrp3Ctp706zLyR8rLvwDYN6nrKufRlfKiLH8AkWtWy3AJfO7f1GKZURA6fsQ4MwjKkrDVwYh8ws/ueopQtjs3RL3RgDXdckoNL2sFzaldwv5JHkVexXOaP4DmkSbHEZAfj/4Y3viy1kLVK3Xed48Mdn6tLlV/xqm88eVfL/m3aXmBfaeCI1bWLFIQLjchTKAoRcUT5eJrq3vbDC0l//neBe9jPiBG2WIepm4BUJoDXzDNKuMGU2gVQtS0kmvJMJrJEOi0jfrDLp1xpdTYAAdpSiycdsnJBbof6tDxPGOoKfI3U0bz7rFG5c+ERgLEOGaapH8LU3UaroSWH3qdA8u8Qtod"
`endif