// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
yB/NBv819KT+5lYGW515TGsEkDTSXXiBGIzYmptLCwpgSqNMZdwaz0mdBQkc
0Aui+WBLCyMFpQ6ir1VLH+O4JPKd89Omp8w2OQV97hH3Cy3g/Al7P0s/PNMp
9uqfG9mju9CBfIq2wAE8dvEzl7S36SOJnZy3q2CL7IEaSP0IrMdtk5dqzM0v
qfzX7BMsDRz3aZ+/2+aqxatGFsa+bkHgMG7mU5NI000beYAgeT5VgtLZ6zrU
O45DaQ1qNyWHgfWlPI3L2Ag+dtxTqcgFPrDa2Pe+nVIB16JfWBH6ivV4NMrL
Rv1go4a7OD/ABf6U0//fgLrnwOkLNlDiyBZeyf0LIg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fWf+Dytch2TlEPtnRi0ofbIXvkh8cv8DbDBV/q++7LImnCx8+l93wFDd+Bv3
/T9YLASfXloMeYeMWNlI/UvGNIXLDKut9LoR/yuRocwk/OdnEP7AKMbG/cDs
MR6ifZjy8EiqZ+smgvLNXxQ6pZd4W+oHNAls21KRxsJZEn1ZFsp3KSb9gWd4
Mm+kgJq8NwFmCko3HQbr0yIf51db0eCrfYwiYPafPEmzzH81QyVRWevMG2a7
qbHCyru1VJugW4HEg2Q7sOYXKRq1iX6kw2jj1slPRJb2C4zUA24K1Wp6MaMS
axkVqzQ2qQjJNq1un5M65YVPOrSG7tGWcychw5oXGg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
R+o/QXX0JzBeoBdhNVXoWapeWxL1r8lJXWaQZlEw01q4ungVvKQd7N+pH0dn
tFnzZd8ana+YrWefsJIcOK+jlFnLiYro44FrwrKAs5l+eoxLs117RJOLRRG9
m0plkXix/8ByBdpgJ/al+ejlBL/blAKoVoLwoMQMfVI1sYakhPkZULQ3kSeJ
vqev9jr40xFMYEC1JQD4jgsR6F4hWbvN45e31qhkHp6YsufDaJySN4jHSP92
Qg7scXQlNcUKRsi/3gsy99/rbU3VLUcA+8hfvku0vj9PrNjaKF1js84V4zPX
GptnezGksZdkYvSa2fScKPeU6jTm90+/qcehB7U25w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JP2TttNcMxO+/OQ81y1lwBTSHqFgLIKgUKbGXqztyadrVpFEJqfDybJH9971
LeYF1JomoOm/TqODoCdLD4CaOBW19vQ8JDe+ejevDgJxnD4DoHLFBaA7JkzJ
Pa/luUC7CFetVcD+KUNuOJ330WbkCua+LOEBOitqavFurRPsLkhUT4YhUOVw
0toNH2nW+KDnjQ1OCFSBpdd8jIhjJFmqhkfQudWV+I4/nFKsqNdDcJYpTQAX
+cAH9BWB8FPxvh8l0CXUHRUilY2b1tMsOUS4g3dT1P43oAwrwd2K3oNhWT0u
olj8PDern+XNV4E3YcWiXjEUozQR7dWiCZfu9ZLYmA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Zlm0muZDRYh+hf+DXQq7vj9SWh70iNAOsjGPithE/RycztAZScco8ExTE96M
Zh4tiD5K1dltnMI+OIOUydHhikmeqeFAkXt7LS6f44GOZgb87R3qfKOvHnKS
XNqjLbGcWrBib8xie59IZR9LR18+yaUQYAOvf3oZpg3GG4GCrVA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
mxt2o3mO6s2umC6dGFCK2xgkcAX9UxLDn5Tt+BZ0sIG961ew2QVBR12JIauN
fGuDxSChMHoMPpJOXaEgrPrE+KS6eKNiy0ra5Gdzi+ZssJOnGRW+9mQF9FnO
cH271e0evE/ffmkol4drvkA6DExzByHizuJtYH9UkCzjDp/I3pR6HdjNy5kK
U5dVT9i7ShIgJz8XrW7GeyMGeC9Rqf02jmeepxGayzrWLaQtF9pHsiNk2jLQ
P3oTm1DuqL0HyGQPzW92Sl2RlIXyhVozd2+U8ppCjwhHpwPy7VBF9H0kiHUO
/WePumFNg3nqmAIYGz6uYgwyCL86wgV9LB3uGdc/CwQmy2zTHUmOus5tbJIC
l28JxzjZ1DM0qgeMvoxCTfehry6NH+9LJrCrJj3mOJItJhevXF19e04JzLzD
FenkPJXEMlmhT34JOMtF2EE/e8tiCLwBDBgizHGpZB8oEyq4RUSAR9bQ2Zz/
Dh6csn9t6HEnzUOn3ZGI7Tsu26rOhKW1


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VbSY4WNcAQB4/WPI+gdPiHgulQKOwmdo00e4xlygVpcGUl+xkQF9PSg+8GJT
ml0b1XnqLgjtrZkiptzETfVfzKfKKpVah4HHQGYgNROu7cceB3PQiPOR/wfn
3VGcOL6KPqu6GcYHmpWnJR9pRB1ho1XEXvAMWzfqUMHUrLk+2/Y=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ooSv+63NyG/PTM6nMPgQcFK4JgVMxLs8JwgbIJSw2Cgn9KMf1FJr9ScW59r/
FUd1xmqAHIxynbxZTRZ0e5Hpzn0Vq0Joq4c9Ggj4KAWDFOYDz7Wi0y2cGGtv
OV4g77qv/H5NVk2+zpX0BSo+eFqsLxFTZ+L3aTbKv1Mr52zoft8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 31616)
`pragma protect data_block
pUum58Km9SA6SAZJq5fCDX4VqhDgYjsEjF6YZDAny9C+ukyRPQuFAmZg/1FU
1coFNJ/OR1vXJOGOVbTomv4QTIK6UjjmtW25NgfJdl4VWIUZ8Ybfexher2+n
NAon7K+h8mqVfbHGZAw+u1fULlxf6RfFZNTCBZzzyvWLJmPCnBXq7X9Ogdu2
+4mES2tg6iAIEAbza2tP63g3rXKHWq4bSjCZ9mX5IaFdH8Mk8SPYOXCoLWdO
XEBj4Xmljsjwp8N7Dgld+r35DTK3kH7EHXVRO/m6Zk/maPEmmhCtzWn7yXKj
u9uJeY3lnxbQwLhe+4GLXjUXc5AvanF1m0JzwO45DvULcORfUGZZBaUmLqIw
JtIs0H77FCpIs+PH7ugYvR3FVn4dVhs82HNvjMUhzmXvJiYTvYCpDJy5hLxp
gY9IY3XnVNNmLZn2kD25B2sGEirQ9DGdRXzRQS/qFKdsnjVi7R47H/Y7Zg+n
lF9f3j78ueDWeGYTWaLpTfOSVJb0f3SmSwuoDU4ROcuZx26kp30Tu8yA593Z
AIjO2rt4BitwNJeA72/qjq50l3fhYYNBdj3ap2hsFXG/31uYxmIwRKJKO9Hv
/D4SK01hvpFyopr9Fuzrl0Ox/F5xtiuIalQGHpxalKYXRJk3qA809U+sBQcy
gWhA8JnfZLh+YVXgPJ6bIO4uV4ab70pGY9AN0EkGBkld6o4rW+I6UpAFo8jO
7Q15+RcsaBbIH4WA/xbnYiE8LKdGn6oWzAtwcqWzn8WdBMc0d8nZnAeJufXS
NWBOKlxXmsXFtXOjZ4+NnG5dUx1RJg3dl7FOQ7CZhsRE6b6rfb16/q8sHulM
EZI3XdGdZ9RwfQJdj4nsq/0Qt1K1lphcdTQKwLm7QI5uWlNUDU2dMRTNnTyh
89yzLr+nZLPdebGXpAGbwWUU/yMm7atPlzbkFOrIuY4lspFXct5sjVeryHZg
uOrto1jWghTSfT97OwpntRY722DNcaBRwFN5UAN8uFnqctRyU5yJZJJ22yUS
ESGZyIx+5oSR+PJFgjWkYVUfOxhfISloqSG0Tw9Pv8DtyFw7e9ZvXhJE3GfM
pFsRVuo7xfxA7zIBDlgLhO+8HOF/qktKU+h79WI6M2woUfZYtnsVTAATiBO3
NkllEqV1Nk5Nxr6sMhGW9n6XLe9l94h5xJgiWrZQxZNoh1vvpTRmi/eMIjdl
KF8z7ITzqsws0QB1kcVsDau1xLaM+w1jdoeadhxSXBlhCyZhiFPfeGpKLUjG
nJGCPEeaelTbbm5gvgFj/W3fORRvKWEJiGKkS0npLoRR7KMlui+zwDPcyGpC
EAmdgfW5n36MyN7YPYQvUfV2f4kRQH1qjYhTfYUc7BywgxKhJj9JvpaJDQ6R
mjStMLfH5B+eX8QpXQZFFM1jMXSQk8h6r4I35Qc4qt6m7n9fHd8ihLw6VXCn
o9eUWdmbjG64nUCc+Qh+Nr+ejzV8AXbt88XO4JNoGknKEz24YggJZeys/XIe
Nqp4EDq656jzH8G5c2Q2gvJap0JIOjXe7vEIh/SA7xP9bIzxL5gWwKtNwNm4
Bk6a89qBIE3cJ7xnNhxD3qGlNR0e2fkgFJoh7dY/sb520uXw4MMvy0+KeZ3l
RyUyrM5Ojk0G96OzXdleXDx+1d3vLi1M2lQRUOIN004lyxYW2lIMJP56qNiu
tIeC2l4G9zGPo66097WUqb+TkLf5rGoAHWv0FYd6GaJheMePd4e0vb2RIdaA
ibIU5y13HDmmMwvfQGYKz1PjKq121C7X572K79THeEiY/i3wMDV610PL6A04
LkZe9eBb0qjTmmvSgNLiu2JSoEYGeMpRR1FdBq7OWo6/uyGJ9Cgpdlg8Piv/
BMWIVEdzsbWnFk7S+VFYWbOHHaGEEvsN+xtcA7g1KnWnTNEeqbbIeXyG7FeK
OpE4+r6ZqeEkFkcm6ORr4UoDUte3aSgL+sC0xPgZN1yskY/7kPBHFc7Z5ekk
UjKTHSbuZ+doeZHmvi+1+ZaOobplh34JPug9RSC3grqb+lRoNy0claTxraoK
L8QjDp/I9jWTsc5I33C88Hj7qNTlK1OB2eSInBxL037B5y5jefh7qZVYtzez
V0Ht2FG2LDai5QaecfUldav30lAYE1/GD/ejArnxz07NvRBVyzK7cpfwRp/U
ESiN9Qw8Y3jVCykhoTCbvC+T6OyN1iiJccwXaJ940dDBFvx29REgIiHETa5c
H/iuBhr2OOZwxy0tDarz+eFkBNbe7hBFIp0WaC2+KvBgOqhTwwr+zX8RsW8X
ZUkgPG73hjWWlM6o4fGeh/7+4NHCTYTUpIHOblNj84nYjROAY7rRIG/zOPF0
/Ud24MPKbI5p1IHtsQrVy8e3sUsxGX1/4oKTJ9I/92Rqc/jmdSw4+HgT3m4m
hPyFnspq6YAdDBUQYIE8Jiw/Bj99abjlw8P1afiqMWv5GpLkkWfeFc6Tffzv
Im0g7CcN2g6Lbbf5iaW4rx2GkKCRm1nzUIOcPptk9RZD+v+AX5NJISmGIUjx
aGNh8xDx4QOPEWGpVLcfUPtINySJ1qRp+5CsQ4UgzykbmlX2iWhb3Co0I/D7
vRZM27uYAE/rMgkAN4SwmNL6eKkjZw4NvWRy7iMq4ffkJffKm7smNFw6fij1
ooCgRwW5UsDkJvJzjQJZCmd09GOf54Ij3raT9l54rU7CfxhmmBUOEUP9OG7h
j9Z9woz65PQ9MfL1DrBGajox7z7dKhSIXnWV0HbMGNVDGyH/u5ZVyIFvU4yA
/q6iRFBjyMHTf+S9lQYKF5ebbE0qXQIZLuYypc2TAV6IrX6/R8baJiwN/eRW
cQU6DNtwExpuCD12A8SM/6+gymzua3lO/v9z+DLEcvWQfmmQLfn4AqfxbVyz
w2/V0ecRL6fuEqF+Tgy1GQA4foa+ZF0kBCgp5kLEKhTEYpfcbGcRKZqW95Jt
ZRVH5UQAOm756mLugU76ft3CF3uQre87lRGXPdxfsh7d9yK9AdrUkIQfgnLu
6MZNoKGinrIxaQ83RMdJYrQsdZNHsaSZk95WL0MGX6fg+4N4iqsTElx7RLfp
0NjzuSRlbw9HKznvHL0gQ5Wh/BPXNej6IqUTnZ1uqB84LUq8JJA2iespGQ13
fN2yZIMEngDDtt5asZcrfdSEg9ny2/v/O8wJprHRF/yE3meBSraJp+Tj+/vC
gqya75sTX/LYny0bSe4xg66MygFLBKfBAvi6ZiGDKqTTo/kJz6IxBj22aCc6
LJc65YmRO9B8ikNN5FzheuH9wNdorbPbYNST4VXk+pYYBavcTJiMEVjU7/kn
FlbMxJs0/LLru/YT52BAdFJOEP3Joas9HhonEMY2ikoZC+bv2cEzVJ3Wxhua
jlubBT2e/jguMmYEPBpt3zkrOUKXqFaBezq1YEZHHcwAQe4p/RMcVux55R+P
2alYAaTg+rO5zL1A5RBxf/ijdbad2pR7ACcvlLhcxrbbrGIq6cuKWPZNH0D2
6XaXVdx4FJjQr3CTfMZZDfdAe0PcTYR5Z0vB8mkW0IYCYlNFopMV6LjzVHFc
svBt3slyDPeZz9lgFgPRo4ufQNJJVLZpx2tBBtqSHZMEAcSS4oR9P7c08W6L
4212cqmR5PPqOELM5259lYTA9+m62AlJI59vGWd1DJ5ZUy1QGFJ6kKThOMJN
6a3Nx4lVT1zfypgkTG0SMkw5jSQrfrtsVh1oIo5j29TRIWaY28zXcifRzYUJ
yXlJcRt4nwACJAdIZfBNW0EE6jWOZGKSqm4/jTfwkeFeYcSHuhVNjcpVPONM
ttDXLqsDLEEC1jYFG+W04Z0UoApOsP3kf7KZ9ok4ilViIs+fkN5brqKN1lCb
uPi6syU2BWu1B3c/gbd+T6JwsUkTyxAqckjBPO6O+qqyG597PPIBY1+jMLaL
k/zKALKnYQLgvyTjz/pCUePIalP1c4veS9ixHYiMmw7beR6rqqZPKrfPeU1O
e8CJhsPasbgl8S1n8xzK8YBQwCklhfCi+jzo+dyXA8LLXFj6XyQ+/Ul1GgYo
4b8GkUpT2FjgzBxeUWtRgiCdjbkNAVP7t48O8c2IrklLbranH8M0gb1nMy+n
QUSE+3YOwX7FoQHbpKv9bSvhhLdfKxQI0f5f5poiTREW6n6ns/+uJcUfQa/Q
+w88hKMnVL85sS91TSazpFeDQtkdYatAkduT2UlJmA9zqypCnz5bKPGyZpFa
Jpjmp14AgaUU3gMx8j7SSPomvV+oHi6qqbobZ2W3Q4fhLU1o3YuIAPgDZ3De
x19FsGs3r/UG8tWVAUCRXAszDF6GUgWfTB5NmE1cN76+hJmn+wQYDpdNWTD7
ujTGfE6EfmHDGFCUQiC9iHvFemelrvLs+EHRrpTF62JWTDLtVF5CSqsTG1QF
ttkwPGh2UyRv4qfrst8VVUaDFiIvqDWzGW0fHWO+ONCGc6aJsyYJ1rnZpRuf
mFSxNXS7ZbXOxo73lt0zmE4Hrol8d/4rK0rE2ZLUbAkanGPrYuxxzhSpI032
OsvupyISngkqGm0nt3q4aZWtwJlFVUFNVFefacQV9Df7bXDpndT/DlVofTZT
u0K/qRGfbMwiBmO9me6Frk5hfxIqRJCyo7y4nLYtM5zCMaeXpmF2msncV0rV
JQ53tyNPDuWItIB/wXkR6WgEjfYORNr2FT87ceiC7ybZwYAOH3sT501kb+d7
JU8Pev4RBjXG/tQSmgjk+62QdF0NiiJ9hf9gythf9YVLsUC6zAkEQ2Shs0xn
e07owyeE3iP8XzPa0HvT2MP7AbPZ8wXD6/JlO3estgniebrSHg3kcS/Okz4K
zycYUbnWcIpZ1p1wjzvkEplASVjJANzLQg7swJO4tMGtLXB6BBszCNMznkUx
C8y5dRsj0QZiomIrvGJzxQyw4aRvE6fMiVicK/ZqRkmyu4HE0cXxcS9kR8RH
lYXSKQghiKJdy9XiqlVIldobAzJrSs4tvpXCrhIq1G0Ppg3jTqSdpp9SEZAF
s1WXf1wD2bP0VrsdIK+8bcDJ23BN7mL7yo7EfzIqxYWkx5tLch5+WVvP8JkP
cVyvlASwN1DXUVf6OsMNK8ilIyK3S+JA0xsA+U2Gq2U1q2n+N3VHrDYHjXr5
Db45p9kNZ5gPWiGt0+Hw+qHpoclXtVup7SSZfPoZVupq/aNhRjn57bn1xQ8q
iwCs4gQmuNOyMjEo9AsCcRNBRS543BeadcHW5p/mG+W+MmU53TS2H93h3vKi
f3AcR+MS/PxTIXDz8gCussStDwy2bRak82XJvCgv1iXOXB/m/CnO+IiT0wPx
yQII2mV/4LfH6EH1QycOdpAklmwS4+Jlcj9zSAn/NseVnlOnGDZja5gjcz4V
Ygj6c5rZ2t5Yib+GEx0WXLdBOdP08p3uFmzVOI8PgR61ss8LAI1+wBEzxswA
ySNqbhrXeo4XOB/mR4wvRPRzzI6+1hNi01HNCfqGhGrcxGn1/1PbAjdE1msU
GgFui6wZluBL9touin/TrlAK/j+O/NwzIe8o+2lUUZ5H81em4b80jDo/MEMY
iAd+WkjSLrAxrMWRJeDPls6uXchr4r5OHQ4fmIxgol6z/2d3IK6YDc0Stp6i
PDKiU8HNevsfcbsda0NEUyik1C8gfqU1eGKmuM6F7Y7mmJELlYLoDbKZ087m
kDrbpBJu2l3Mo5XIJEAb20QRlo2ZQtIMO4pwkD8rGHllfWPtUvegkhGv2dRO
bMZlP4uMeaBxuvryZkKARqfnGg5wuloavLdm+a8QkEdX0/nHojCvbwluv4ew
IVNzKVGEf6LHBSBKD0H+qA0hznsseIN1Z+OX4E7vJ6fCYFHpNwJbokcPJns/
OOg0NQ/aKwstk09z5NdILfh6JmpEjj897N6yIXwL+rV3KcgbxTVT95pJDYZV
h9AKY+OSOcyMVw+k1IcxpFSOpyWEvPkjw5BH9yGR1hwPKl9Zrs0ABn3UO/Sh
0YjfZaFTME85QsQGq5lSQ/o5y62tzsp8S/urwTG10qqXmOCOWgY40V8vorSQ
GLWT5KiguSL2gtqMusBnrunuxKYgK/AieYHKdJSJSsDC7a8G5rUfTMPYIzU2
iVzskunFdWXvpveUBxlwrBABm2rxGrZIxUvGzWGSw1EtFa9YVQDpoq2KRY3Z
uRm8grJP05xQ0Gz/Zw4R7TB12IGR4c9usnhRHCxNU1z4v5yACT3hJl+2uOc9
6Z396lbBAg3CQUHDxrne86tFrWT4cbGqETZSiyYHIiTi/KqGPeaUp+rhbb0I
fEtPvyCrOGPPYVj6k0mssZPSvg8GTwrhOvK5UUqS2tPcNXu83ouoBH+ydmBQ
SjBNLBa/m8FLiExBuMtWhE3zHphmTPgDgUg4/lxU8F2hVhvx0Gc+tahsucJ8
myF4Ws+BsBYQyY/eib0+iQTn6vpik4TruURCbSVtqqdZ8h+sKfWeHqIaa73K
na3/pfdKnXlo8bP/YZUfHub8ev8ezioG0UX9EexolYGVaHlEe0pFHilsEech
qnhqKvEW1O1+uU3rImlHBfPBZQYryvTRFy6WZTl5REIYzL8xVitUaoXah61y
VFDJKA8zt2YKpwMr4eOwbGzzgVtCAOk3HNvorzfP/Lp6RhoovkT3H/H0OHTe
UM/XDHjpAI+GZbvGeJp165eMUI51+PH4chFWjmbUZtN1wWltuRNAnykeEMLa
43WD3NFCR5Fgo5V0iZL7LUXyeXYpD5fes7gEPNKEUG+a/TMaWN6J/kXgwy+4
pQm0RNuWqGP/Km+PmNHzffzzpPRrKlaBYBO8A1ziQNBQ57fixfiaFqk3yjSJ
pDirmFqJ/vZ/2CE8AiVGIzR2o7Rv4Vjlm08xp4KF5fGZ6bOcbGtk3HfeSNpl
8ExWP0FjuRJ7fIVpoBF7qaBSAMpjEo8qZ0XEumsOyE3waVJJkWiAXPnIJpjw
3i+87RtQwAK9L8+wtbjsNNn8DWz0DnI/R0Wd02Fa1sBUdXOWLS4fZyj4j0zX
hMGG2k/J9dD7gH2DjRK5MqqW1RY3WEgHJxyor6c5BCB3ETSJsbNrprTzjRUv
CQDMW+PEB7f0B50qJTzEWmbbBqvGNupFHcODjq/WLkWUiQLtfT5itz3QVpgq
1u7oC7ihrMgaFDZlYmRWWNr/srinUsZ/WEyROQ166R2aedWCUxs5N2cCY086
hBurQVHvWc2tCCfKl2OuGAXPmwM2VUu932yvMbaYQ60f+Mvxz9IwRcmGpkBp
NBscVv9HTFQ3kRd/JIt0sgy+Ot75Q2zPU/rms6Lvv+g4JGCYGc0+5EJXTyn4
UdcZS9L2RQvFQuadi+kxhOtnL2N8eepd90VeEXzazbRY+1zmThDcHmoVAZUM
usL9F1Y9LTitNyLJViDIvcD7f5da9aV5+4g/u4s6U4PuzKrLiExyd3HZq6rT
yEskchhDewLhTLy+WmGcASK7Mlef+v8cacXZ2Tdgd8STFiVjFUgsW2kR3NIi
9mM8GB+suuQ5r5mGZAH/+zFOVjMPrgHKiO1DWocok4baj/TNSUiMokwh3jPb
9KTLbDyw6fQloHf+xeQoKvrlyvpATMeVrCHPNE7iK2+Ta7UOzSJCSsOqPWxJ
qcVla/n+Z06b0UPoYGTgrBiOhov1mstUzNvDRR8+cWuK+79PDtsi23Q0LB5F
39eZcl3rF3wWycUFFN+lSzDzdoC8g+YsClqKhtiI3ChLQY8+B6QTX1gv6IeE
9ErDDsmsl1PqDBbecJgnqDzPydsGd/eoK/tu+lO0o5iVhuJ6VI1fw7JGou3M
uC7XyU2njtWerLJOpSTqEWyMNC+91wcebWFdhmIFp+LOaxwbxpO0lt732ugs
ef4eG9v+ZrCda+GN/SE4t+xlZjdjgqx+8O8al8VfWDSxDAyuhZHxZznz76Mt
eMwDFiV/4T0UPI5UA5K0sucS0bl8baQP5zo9aeEv9sRvng4JzFrXg5cqWTHP
a9TWteH68Z2wrs+BhWd65HWn2h4EjLFDGdMvrsCy1Oy0x21OuYl9VVHrQa3s
ZfdETn6/OSaKxztBvvgZXwtDdCLXOa5KKIgNvARCXZpiFfEGZ8zkPF+68z6B
51HBj2fW/89bDwvncFZfG71c+j86FQsNsX/yFNT003mmArGsUvp7lQ+XTQob
3byH0NQZ4Tp5Bzab5ADZZLDkguRMRt6Nm7Hns4L+VFp3NSM6T0T6GRnxEcDr
SFtBSPO6gF6zt9gbhVfFufKlbhDikH8yiLiKikORJRMNWsnwnTtbIcp1BkuX
adIhkiOavngT+1xD4SEiUMsOjhMS9Ar5L3lLue82e5lUTOzfYRx+AP/72oRg
F87X0s3yi0ez40CZNgJMIvIzbMElzFxQpdWP9BqlrWeAuJAEe6AQv/yfSQd/
QhA+o9zwer0ebUYTx1/TLppIpk9Rl0RTOB04pqvFwvKF4Mo3ckw54C+IalbH
JPmEwZx2fNS7sookxINbAD2G4Z3twBD3khMkjV516/Wbu/M251zuYYft4WEh
JKzDNxdiU3MmTMPMxojtyqBRBAlx3qpO74dwmGdJ4aucg9EjvDt8v0U+1B5L
putvYI8iRhIITr311K4yBAneasDu0A2BB7sRIuXfD0PavaHfuWOUpczms9Vg
NMuszxjhxrQa+0PQzaNOH2biD5bF+UCBbY+by3rUvPfYYs0ycy2eYBU7FYRd
WICP5E9Ll8Gai4aI9N9aoriZ8gaZF/8icTxRFcxEQEmB6INm8ML6kP40+Iuw
wHBVJhRspswyeH4UbtKFdOhDvAw3LP0wp5EMdHzkCnDZ0H6/3NOOQoqWjzrT
Afoi6fekDYshk8/Y74x7xeNNyYiIuIdpU+5kNNi4KUNpGlhT0TZhCtFzii8d
gUkdxUJfEk0WpLBcTuWScUG5T74purL9plXJEHk/J1FtXdIkCVtJwvs2Y9bI
1pFMmih2etrcjyCdXaxNOjcpdZj9vx/pn3fnUw4s1sxAK7LWfmMg/e7fwHqA
L/XIJJO9/bdCLpgllYcyqPfRKZGOedrmCdfF8aavEPPhcsReFPnLEF3eJHm7
ccCzOE+kR6sSSKx1ehxZPd/6QQqlhVgAa5I8KvSljgsVcF7TMrBxUfLmUFlh
yQp0muW8XKhlkBnmKMRsIJNReSVmWD6/O/nRy0iOWR9iENnRj3PSpIJXzd/Y
o1clcW61g4G7h4VnAEOia24S6dEwBwOImRFcnkU3N+7rKdG9gAe/OjFFgEDF
ovt1ZDQp0kt5eWs0GykUdUIwgHDxcOYcZOcBBCWxs6sWEIRA30s4Q6MY/PSW
meZmgnjKj1hgWGI33Z5sUNn/wKDqJQrAFp5Uz9ry5qTLuIU50KpQ+cww9n+h
dO6cOBc0QFz/YoocfsRQy4xmPjt62/UJh5cijq76LCJvTZ4/QS28oSD3XQKS
CBJ0rk7lpijgiL1be88PvOfBs8C5MJ+D8oJySRFYv7qZreYPFMix+hhtRyTL
WMaBEhGy2u+r4Fcf2Zm38odUrbwQEROd9NvjOPlNoVR0ohZDlS9llU6/sbxw
PrZ/ifpPn7xYbfc6wIocDlUhVWKLAd81bwLEqE7R8HqaMQtmrjx+tib7oOue
i60yqMFrGQ0DAR2JmF2LzbrkAkKzSmS0ALSnibwPIyUwquaEJJc3Pc1Uz7wx
9qxsJYMlf9SoctorUMM5aO6kxYkCoaU+tnpzBrnIxiV2suBLAle1YQbatpPm
Bik36XpQmqqwvwEIhjGg0SwdbcPgYtYZuq9lzhsCDvYYf3MKAY5YaP4sM/CI
lQHWpTb98a0w6deec+9rIBu3FUveBmGoCVLGS0tPL3SMyC0PjCks7PycqzFX
V26hbhAT+3nbkEbN2LXP5iRgALvKjBu/0c5N8k0McBA8OXvqLgVI+qwGG8M3
5bsDFhdv6t6i7y677KkBYuMLMQ48KHkDFtaxQm6LMoo7MvPoZ0bugltCu0Yx
XVbEbDSCk205aYEjeMTtSYuCmHofNpXlyWQJqaich2by4ZBVRGC4RLIKw1+3
6hVWpXIMZrFb3RWDOobHeQ3P/cXDulE52wSaUUGKqTNMTlzVos8ru3/TMwzL
avL2fJdM5iXxCAzg7ipeYe+wsPdtIcxIfe8MxXzRsdXDVmdmVjc1w5igJRdT
53OuuV1GmicKLXiyy2wfSa3t9bY3OCAM/3kmbkwSlomNcTq9XtmgoIIJl09p
LTfpFHbSESC4Ho+JkG9mKJizhlB8MxDofvhDTOzt+u8g2nQwJXS+a7c06m77
CNrlZ3eK1h/bdN0lLW9IFkvKc28dOkafT8gxANCSlUfNLqo2qsVs6NMVjisO
gh4sfV1ICwz4+NDEQuK0LHlVfcUMHXr/nxWGIk27O8WQc7kx4Ev4g0YapJoX
vFLYh93xX4lGkamRP9R0ayh586duVsW2nemwJ66ZwGDw4+JW+1WcjwggCyal
dNQH8IS/N+tbzUYbOMQ1A3nRBUJeTFDZITt43xqtCjKZYIG3cfGZkPX5rO2M
Z6dcKRlYtEewHKLcBkqQ7TDykhzpAKwDn3SrEyLoXHFqTYzI80IHkV+Axn08
qSI+ujT60o8gatVpNqRHXqN94SzycDwPENpSL5+rXwtt5XkTxS3u5MBMWI10
lrDnRhyJUdINON3kX48jFhShfx5E+/PzSjQry5sxJiMclpET6X0rdGylCpsL
l3D3+pbcte3KayoIzwbw5kiXYd/RYl2oxA3xmcKawe0oL4J9nQv61jopoVYQ
cIzJ0+b6U7FgDilpsNhBHABtfuNlsuGLyXhmeMOW39F2Rjl/VFMzFzovJjka
PJcBhwoY59UgaR0YWY5vQE6dSq4G7g48DLkk6DNKKiJHCmQBVFz/zaYAJlEF
QRRxc2N+MsItBeHA5lwq6BwoVfXoqlmaWXSg3h7URfWXt5z6WE4CQCdSLLPV
pQk1kEKHKl+MWWMR34mcHi90mems7GM16SD1MljlCVubsudF1zoeIUBUyd8R
9gCU45ZZxmceZRvzi87KZ8el37hwY6PswAnkxnYjVjDK7/+Zjgk26hXRRzq4
OmeQJfmNHt7c9XlivtNxktnUL8vv2J8KkMGmh6EqDWBGcBSD84gTj6hA6pX1
H+q3Q/7ebrraZManycqgPt7dMdq8w9IMJu9mXtIxr06D07rZThPk1690DsK/
I6xqPGCbsGDYOGLPAkBO8+Hl0mOWVYrtyeiRIZkXPToHbul6pJT1NgTBN+pl
d+nhCMnEiqgyeZhmEeDOt2V5m3p7mMyTWTGE1YfTnIA5I6x8whj9zClmEt4Q
4tq7GWXXqeIQSDZsC/p3dwzEd5JmOLbwy/kL3L9mwoaPDVsvSTeU8DjjQNll
bAiWpLejY5r3vNywplbBTpAcHzYHOEyGO37UVY4zrxWY0yVqz2YuhecRsNHV
VqJElf6H1vLfZuU0VW2GuRHh6p5QHZDed0dBYhOJz4Ao594wRNC6rgZLyF1d
O6OunKGzezTpRWWZKBvHOaic+deO14C0wZ/UA+Krgy0DHpA9bQnkJDznf99+
Fw6j0zafmEHE4BdguMZKlpA/QkuCiKZ8ZgZxCC3/lUi9v2M764OCgpW1EYGo
hc0yA0EPSFG/WNjJTB6RdEN93CcXMplLj25NiFfN7/Xlb8q1tx+DoILGM1kH
Cwvvf2QLoRQOr04+Q6uAIPpb6dGCU/u4mx1xd4ZHwRGC0FZLQm1KrPIvZbMX
DuwApI1/HwQl3+9V6PAMUsvWyzcSZPF10vPG6RbRh7HS6kRj0MiEKMGRJH7R
1QD24CicsZiRzcJ7GLpuom418qIpv3DSylpOIazsCe5xE9w9IFdHjzrwne/6
cHUOBFa0MGuQOOMFULSKGdevq0VaEH29kP/8uLSrnQ6tVsUZjaKXpx1mD4H1
u+vnrKST/7rCiNpv0k2nWwQqK+pTHntycvCCIfIxzWlCA1W+6pYuMVkOjSm+
WWRbzmIWPBP7fvbjd1WohnW+1DyAkoDtJtMAsBfhavNICk30qpcMXu3SKRhK
U43vePnTsemae0NgUsjmQSd2RERpRYFiuG3LmKGvnHU+NSsGrFO2CY6+zwUt
vczqG+y0A6XZZz4WT31iV+ksq3EHRfGOx/Ca6C1KOlQS1gqPc0j7Ds3FOBbD
ux3J5vAoWNL2b4wlz7C6TWibMCv092yOshdAyq4UP0ZXVfbDd9qoh1R5UHD+
ZsA2qntBQVN/TNxB0jbjqKUfpOYY+1KCFy38OuSsyv5b/HJFeucs3tyjUUaw
W9T+SUQWTkqgDAd+EhRWimEu/Jj4e5kFNckJ5YACIF3uap+Iyce91150/Ct5
PsMiSMsSWbTLK5no5nfjUqRxYBmXLbcTx7vMgxk52vNNEYAPP8gejH3kvpHN
qv/BGFrKpUjN04tnEJM3aDynjP76zNDqyma854XJtqBNeYufWDbjjyhmIo+r
WCVdYEov9yDfXfhmDZzRfgA65my+SGjqz3G6kXtjkwyJbn9rD/wA0/gLfVzj
CPrgXjtc0lLWrRdoCol1AgCMhuNsXbL3zGE7ByKoA9Js6O9M/Qt8o6JwIo4F
k5FA79DR96YA4NNijJva3H9AMz/V6GJSyar0WutSFR2K1qAZO23A0VbNN9Mp
s6ReAPiEsANZLFbodUHWJrSOImZf9RC/WDdGe47CMIYoFChTWn0j3Y7WsDj6
689VmeNenv6flZf2S6pFkt7pr8HOsFIpQU6SiQK2omYv2wRJIj7Pg3+AEMt9
IW0YnjxOLy/Omp98a7isPzJhi7XK+qlreYrystkW0jOH1G8r9wVXaMCvaDnW
BZ9kVJ/aFhdukK8CNbYNZMmoBNFOn+ElH1Iwd+3Ho+IlZnIeMoogb/h9dvpl
QsJ8Jpmyn3UXl9poxoEgrjgjG5zURIyo7PT+awQA1M8A/C0DbN/6cYNGif3s
SncWhdMuU7McqducasTl+dlop+GM2+xDSmWgogPkh68KQAusp69K+toqh6tl
Be+iIGbjpALSEaQrMuPN0sIa0XXUVH3O37tYfXxadNikJ4Xoa2dLtqZ2GV9r
QCd9iTfEmC/IKe1uRalCYJajxK5yUloBolicy5eHIQq1GVZ0dy4pPrKxj8oK
VJ38i5DlU6V43cQblovY6ZxdvjKAbDkjm/Do+PPjPzYnOv8dacpzulmfNf5d
qCR36VAoXGff1Ke5bgxaAobo8QIlptfyKeGhUQBlZdjeUw92BMfT/MaCc8uC
6YjsGouBabfpf9JPy13taM0AQjNBJ02wF+grkQl2bns0lM6Ox1DCelzr5Rlt
J8JeVUGi+TgNm8aewhaka0UWmoWvcnq8Fj6jaW3Im2wPlQtstLSRxshQaRX0
pcljhVP6IKEfBnOOhB9wU9Ioi3W0wlIqpQtL4eAnXU1cAXnUL/uYbChKpAs6
5RLBHri3cuXS36zozsi/lH5Olu+86zFhaDLdJp6swkqSjeHD9IiaP6KxrO98
kWMEVC4KKe4hcqhFVMEst6JdtO9RuTB4f1q57L4A1A92g63FpINfLcVYm0bv
vtiDMcN4xOvdff5C64EsGKqGf8LwCT9G8BQX9OKG/A1hY+ZT8yxpAUoOZjb4
qcHoum8jLw1HdvQNqJHWfW8vX9QNYjrJm3xxIeS9Q+as12NPgsQ4gJGHlmFx
vdXpAJu4M7ReLTrEtJhBatkV9U6wDwfZdCH53kO6JKGLghWqrAokP+m/HoJy
ivyGpbfE1WyV0aR9QnNiQBzyquJoYSmGlmnDUP8VdWZOBj7LSVKSvBnwmAaO
/kHUqc/ifUp3ctrJpF3BTo/BKRPHPx7eCgJxPu+erxmntnn8KqEddUnqPjyj
R08g8vAyqjDzpUJtrubeaEpSrp1YloCVn2h1Aeo5qGKA8MrIryltTjdHK5TH
SfJ43n+zcz5OZCo2EMjIFWMFIE/os4ACkaIND0lXnpVv2b/Guy/XjRnrEM+/
kGMyD3ISkOOtjSU6FkpGePEXh1NXAzXX6vDNf2sIfvQ0VZOt8P1exlani3SE
lRijm9VidzUQGbZCh+aAbob0qDPaLmVJDomNDs4s5IlSTPIn4XgEmmtKWeUJ
g6gkGiHqghG393+DNcwo2TdTcN9xrXQW+d9U4Zr3jHH8eEHr7cbDJcgQ5KM3
/v27HHCN9DIXonzNjb6cmIzFWpUPi1V5PKFioXwAiis6MflWkHqItsY4aH76
5aW0bgAp6D+45IQVMjQSU2T0ZKccBBrF9lYRcjjyOeZebZX7a+lDcN2qYJZi
AFeLIiuPUPTThXFuOdczOFhWxukkVXkmRZdoK23O+WWbprfq9B6mxWpCUAQs
jS+UXPf+62A3rA2Dr+RLhO83s7AGEUgUHImwej/nZ7AR9IZ1uECTLysqUljH
WDpLgpnD4Uz2+y8pkPN2nHDkHZ8TV1Yq0pbokgkf09XyhSFn+p9eNUecJWTG
oyTh2gW9k/oaXkSZYm04iHxfc6oin25gz2NaUJs2yFvPSOX8tFTF+fHRWrJK
GsfqhUIDEUPZ5OZhodtJfGJZEF9QqJ2teqMDwd0eyyWgvY5mD/LL4fz3TIE4
rWIgLaOUKHYOf5YwpG4DLbZZInnpECbm079Yu2eqji4PrViDe3XTxSNJ5rhA
YZ53hRzIp6cVas3H7e3JnKeYHFvrVy0OMVNh9TB4QqdSw8OYl8DSNQm2r4Gg
pL4phmsEngVQjmy36caqFc+iaN2x2ZLIlecQqNWEe7Juj7Dhjz+58yzcLp/n
THD3UXLLBqbIlfcuPs4T5vCGOO2cRncBnOCLxPevHyanhQITxSjbGkhvafRj
fjJN/50nr+WE5O1qFILR6jPO3NBMf18RMKDPYgI4fTcarl1M82re/cWrcVIl
UQiyVKmgxCj6gwvBBHqWY+ilvD6fvIvJmCB80GpauAx2VnTmWlR3OyKViN+k
hgfmV5pybLFomFyS6gHzQd0aYdm9XL5lOkgZjB6xqO7r5U5lpAP5I5Vi+8Pe
oPF01f/lDgnS79H6pCvMghoL/24CVLPqKeIEOn+Bsrx61Z7HZze92HFsa7kv
yxMdK/hLTZlyWoRLHidKH8G6RGCKchJHJkJka0Ssxjx0cX/hPUFnAWJxfLyt
UARQbeZ33bvoDHlfYqbY0omwXwzH5D5JMLP3w0OAF/B6L5ZVAx8mTZgcVWsl
wBG6xREGwT09QyXxJLE5Yz1Op6n6a9QS0RxR2YN7foS/5a0j9m6jn+Jf8zVk
htKBdTwrb1BEdgM7me+0T1qMmWSH7OPX8UkbzwxnfKCF8/5LMu3iUKpGzBP4
6EHZgVJwDFnpthUljv9pFFc7cI4X04i9HC3Y0xnlqagVaw0sSqPKPxFZPoRT
WDebjutcsDKbCiMHKT8mL6/LP6brSq7ASuL2a7O78L5fnl4b5SvRagK3IZ5z
E0o4/4LcFmJv/iH/bTae6FT9s7UpGr9+WBrVrYeI53EnjWXk1k8w1B7sjZND
zwv+8VS5K4W+8M6mvUhyMEslq2KJ0jBYi/uu/RHCcag/MYu3UBZL4IxplqNs
oyVQmli37qndLqEJNCFGb/jmS/gJqxiG5Zaq8xAvDj/pxQtZtebhWC422MPh
6BhFDgKmd3YvRddYPOZIzfwJm16YwPrrgxkQErXqZ7Aqwlp3/xXDTgahFLcY
7dlWFW1K9je0K0FeZHSgE2j5isMtoN/ByZ6XKOJqPQNEbJQ5fh2reYczfwSd
VXh4xbrrEJ0LHUzr61yWsjLzEh5Ph+kLFK4FkeUEPMaJUOs4NBlFTwMD1pVu
wSHQ16cQoyuKIX34291s5x6dUf7YzYsbcaXqwco5CqxWTvNnhyY3hrFoP5LA
nhUGRswBdoqitG4dNLaO+14QAKDnSvWtTQapaengOHsC1fQ6FPaYXXJHrMWn
Y+oLfxeI2iBLVRtQtqAfNsjYS6PBWnnkijCU+qsrMJjdk5/KN4tCSOzs5bAZ
3Y0UIW+UCqqYyfHh71ym2meSbv/OeCVNoS9F80qlt9WQmtMe+0xWHjv/DxLj
nxGOPfJtTg2rf+ZAkYfwfUHio7jKF0pxUCeAxpi9IkuX3CH8x7ib/FsIMqSF
zimi53FDTx4aerfH9deTFCMTtpvJp8fn76o9lyeMSXWJyYb9MH1g9hK8/qCm
hIg/lb1p6+rZ09JbsUWGbSYYLb82eEUMyHav9465vxOURNgo/20RdYZOcOzh
rSaC4ZzYRNi/T6fki9+iNyRwQFa3f48r//gigvfb8cF474bNR/BvyyUL7jqo
qH5280FEr2pbFdukuAYOMMM/UEDxNd9NEUx2ULywFG5aX4hr9FKbFuBGvvrA
V/bRR6NIdoIqjj4pgjod2V7S7Qn5iCAvjwd/u+hdBMg3KydmqBxgeUV6OJw2
utdLCJbT8yWX7CgCWsoqAMob1ZyvO40M1aXRs7PYSUt6fSGrUQxvqw7clTyj
JatI+DxiIjVk7G0qb10MyEfWFEPjpXhBPzmpDWdClIhqhto0tZTeKn1z09rJ
xW7qSj78f5OiWycLV3S+B9Fqek9mP+h3SaBlT59Z4FtPCmNCOODQN2Wdm0oz
26iAgfuETp39jnfVNem3AWssWIty7jvn9f/NaC01pSL0lyMjZjvt4ivCfFh1
4oz76ZMIx3J5qouP4pWpQAyTi9lYo87XkyHsrZsFlrzb2b5jk//yn1TlkkGx
zifL59hiiK51bvLfsM0P+/iBQ5iAxlH+Cmw0Lh4ryhxFQ/tWvteSINR6Hp5k
Mr7Nl4Y+EpQT3rubz/yyNmq2E7jiRJ36aWpc4R/aoXXT8kXiiFGcdz4fqXYX
o7Hi2psxjTzdkAmzdx36gJd3cL4fOGBSHkrfn6iQT9IjjqyjLajsz3qZ0miX
QkEvsYtArXtEedU9WnExIoqVS0U8Qeir072J1MT8nX8vVAwMTqLF7T8XEea6
MH2KO1zZhbIAjA/YvAv1M9XjEF+NHExnkXESOi1ZbZ8hs+vmbbgSnQt/e2ZC
L7jZjLRR58y0Kp04BpzbarkH5pRb7YGOradwMrTWzc9ylIPYvL/CeM7NZ9g7
ojIh0u0kLF4XvZkVXkyFkS9HMBIpdJ6LI6Avj821pAF/T99gBhZygevpqRgR
6f9a12SmCxbitkMIKDXSEoq0L2/3IrEXx82PaKOWnVkX9HDhoB0yl7Y0qQq8
ZT7503JvAq6RCi9B4YlFKrdnw/bGQ7nc4hmzks3JR7q23TpXv2cg8IVomH4v
U0INqhqRIRygh64ytTcrZZMClKdUtmMiX0ljZp60iSeNE3FH+9nLKS+ovigS
CzQJnlfr0afwFLxxb3vFAHg1YgQ+o9kHWS6ryxxHFYpGEDawhqQi5YgxjyVl
S21f96sg+vk4rqVGjRPst41CoCpJ30lqQ3sLncr1YuwSPSLzjIjr1Bq+AczC
RP8lngmMjRi7dcoWyPbkpCf7CdCVlFx/I5Z6j10xsVXTD89su5WNC/s/epxN
MoaXtgmq7PEKmCJ/r7SsHXhbUNK0P6DcOUNfn9HTIsaSc3LUQ3nlhdRfDduM
xLK9+cgS6w2QW16btn12MIeQKBJdErq4ASfUaIJd7j+AYmcew/AV6slqegNs
+gAJM/fn7N7Pn1EnDuD65fnq2n4nuRufWyrtaFl1pHgE6ncrIC6/kI03fchu
e811zuRF8+phZUI0ILi36mnKUWd5X7nKVDXPK2s4oLln27ozORLnqoAJbxMv
zFu6OSKyWbpKZIAdNOIKPC/0CpFaKAhaZGlFHLyFP3xlPh4zA7T4Gj+y6PJm
h7S6IyDtcTcq8CJvG8eZ2JAsaMdli6HycoqSIj5YxUrBuvBNWXWKm4ZxOg2e
olCE/k82mE5Fe+fYGyXLJBxWjmFIQbZQftg7vUh74lc08//srvJhugrTN8wA
S4UwKqVTszCG0bvLCgnnYFTvwZqEBAFJqDFMvlvqRuNQjR9X1doCp1ZtaD+L
YeSZ4TVOd2jEz8mHMlLlUQ7PhtoQEmxu2NhpRljizplTeYXiN0M4E0AfUbIK
5c58C28zM3n83MSUgdS3QA3QjdgVCqeu0ZxadMJIl9a9nKDz30U7361/lA1p
UugCNvOPDprWurGomVm0hbd7CLqsehg/SwHhHDaXL56yo9ZMFrb520uwHVIS
4XfWD1EvezT9wbNeZLssgjiouWBGmWye+5XV5zxxJ1GWdEbLYmBJ/UgjdAFt
DQam9wTeft1NgO4QcuspUtF0P7pEamHyZoxJv1LeHNUN6BwvTpZwoy3TpvO3
c/hOi2kIsw1CJIZG+9HmQHsRH7Gt3Srm/hULhrm1w8EJ3H0E58YtKYssB59q
Fkv6aX/Zrs5Tc8hnBWHuEEqmg+FwdAhi2SSxRTuZ27174ft1xuAGKahDQwKe
0WLeFnBu1oKiB5FTlGxZmuk/B1Nm89H/gTl+5AAW9J7XqgDpLyWPBjixH/RY
H0DYwnTy6jlZnI+e/2I1h6GMZ8beedZIuc+NGXLD5skTFXJy2ZRYwXE+XH6t
xzBz7Omg9pgBeejIKpQbm1kVMksVdwQiWjvm6hhdNHVim2LCY/hzqipsxTQ/
on1lM9fKAQcV3DeD5Dycz4LWGmP6izC7ieqrKah3wBZ6w7jYi0WxgEBh+Z3f
H2AM6D9zt7N+cc+nbXoyzMB2ED1WcwTQyUg/2jMRAZMyBhQpuS0vgfOVfZUa
6lNwX5dKZNC2M/ol3rq3EuTrh6p79fybzehD7tyQ+kmyhMNJEsxTXNXCneAP
vqplI0bqGM0IdzKxmFPKrBsRtNaR5xizY8rQO6ZzhaBr1ePO//zq2cgAOne0
cFnlxMN8w5Mu+UVV3vncHRHkuwFxizeLgxdq5pXmh4tmE7Ox7rMyJBiSlgVc
Xyn7iiIEvpWlpiEBuYiRU5wvq5HoLhgr19fAO7CyUuFNCzVGnmpcBEp89yPV
6g/hPPi/XcaJNGexas15BHAA5Ld7XGv/CpcoR6JHOn1vY9ic7ejxWP4v26g8
Ain5by5jW0QGlHTT3vOIeoFY9sqzD/kMKoj1amOMyo6Lq73FiNOcTmoN7dFz
fAALgDtUN7wf4KJ2JXuyVZoMuKaeI6B5uXD3GkLQ/SV9kNQX3uTIBGljgerW
OEdrT+b6E4GTHonrWn3s7iLCvHl0iSsjuRH/Y7JqJbLE/Gp80xN39H20EnaL
8XF83HtAgEg8N04mg5zxJCJhkOiq5dnAYP1dG/lxTSKoTcJn8GwpFGRbzL/G
o96rXoVa0Gr4/xDGzQ/d8k3pRSzNOnchJESUfcNnz7EP1wIBAQ5PXz5Q0TvT
Z5XheEKlzHKP6JGiNLmzC9gbEwhUOu+6dznp9ot+HRWLGiyhkD0QovGEv5Ji
pS2F4hJg15so8XKMQRyaV9giu8tkMQVGEtKlPDU0ydKMWKdcMzPcJvNF/5vv
CZihdLElvWxIaA32ItxXaxP2cfx4y1GNDnSkL1i0kEh/w2rU9bxUlrEUXyPt
ofHeNIhPZcFtzkUXMSx1gwpWp/flTjfZwRFt1oiKumAqNo4jd35R6GQTN15e
Syb1lNuqaQwBq1eQ7ND54H84LoToLEH+sGhcxmO/rdd/FRjZlIhDkm9RGPyw
YLzntfH12zga2cWyAJ1zo/mRn1HR2bpODVRKz+7Tv9TD8lhThnsQG4uqJkwB
evzmiBx+a2+30mtT90JQve6vCwvDCMcUr405LEWg/xBuPupitJI52wAloFvO
uIEuP6LKIUuyeBHuG6Yq/AJNLhywYRGKKXJq35sZFafasMOH4zxsEkfYBbvk
13wsA9BU8vmQ24Teoy03h2fBEPUZzTJhPV8EnYNVfIMmbOLp3Y+SD40IzVCE
CPIXwWmZqJY1u1yKVMhHXRTY1JTHgNabgi0cbgXN/HRWS1ObCKUDenbgpLIz
ZdUoRGIxB/21a4L++hlw3lfwya/lNANJric7KYI8aR/qM1gX/DAAgD2AJjSB
czAah1cnN4KgB1FQn4mxQCI4/vR9GX+URYXfx+ygZ6757hpXtuG1KBXCU/kB
2bAx5VOcpPqSKu4/mPnUL95cX1uHT3guaWjuMyb1/PTSqgjm2U1aFJ9r+shs
MmG0yNRClZ/irFU6d0+T+s2F370ZHXKO20HjmHbjkt66Mxu8kbwwwZ5LuCxt
HXV/xLrvdjvwEI8LAH5tJyAyTKwzHI+yk+EqL9rq6PEZ2ZkG7u7hcwZWvVV/
yIYMp3m2PzBog9FiokSfKnmkcvXugH6FHuib0ziF5wHsc1/12FyAl2kPg9XI
+rL6PwJoNWvpwz4KWNG7QlMpza1yfZYI2al24XcizfIX8+RKpyvY20P22WEB
3a6EHf3IrdLyX4nQYrgMUxJn/evAz+qaX7MjwmJ/Aj1ekRu3ILWZbWHglgbm
lFK4eBIpiy4ziugfZGIpCQNvE/ocTBqQ4C93ZYzWo5jyM+/zukhix/oDVQiM
lBRA/YGNIOXNSBS/rf4pzLbBGQyfnhevNjpjWlqPdUyafjM6elwUMc8ehFyw
GPNgN9ZytcLu2LAKs7kqb07TwvThos3WfyeuUvNhT9/L1l78jtzXwosWrwTw
UrM12kGMdXOwe1pWsHlMLGGNCKQ48dwoGFQhxYVPkmVNKkL+1capMniVVrYs
4EJzypYJqIdZ1lAOP+RUfn5UKyLEX/elBHjvDyVjMqJjmzWTN9+JYmsxb7X+
GJQh7cTQ4+2bJ9cl3bwfMkVbqL0wkm9kW9dlvGS7t/Z7/4i39sWkWZfgefxh
EcJN3rEPBc99WKfcGtBXW5ylVp/DswAgakP4otvWCWeRy/q8646yJAfmSZC8
00t1/LYQB2xMHLe0mBfyjaE03NQeYAectZM3VplwT0KbZx3LZtMhzaA5PB4K
OlrsWyA2hk2oySKHe8+D/JOlwwxULiovzqPGsIr7ycXtYEghL149Ae6/G0p5
A9B4r6KilaSBcHgaaQZ+BvLpk5vzj8H8NlMP6ueiUU9s5DjHRpAeien/rK+q
8mdbRNOrMsmpCGa+pSNw6mcE9Qfjk8E01Fr4r6vodxZ3gL2HKfaZ12I0jvR8
gBpwWwvbstD7VFXn2p7P4/uR3u9j25DSdHnldiGEwc1xyNFl77/GHpK0UALx
dQdsnqwDsS/65jSt/z71gch6zy3Rf+HVqWMX56/8VFXO+hjGk/4gGpVCN5HQ
/Ssk/o2jSb+d+DJ8R0qUvs9n6eui6wVZAvbp9fd4Ab7MJ6mSGw/VbVj6blnT
iMsMYxnSxmIteS4ybGgLFdQ8yXZKCber6uQs9bL/nTqU9XTme0hg77OJE2uZ
W58Mi9S6U8w+vQLVOv7aLwX62BTt26wLv/XN1QVOoUlQGegPCqbvSEW7baZq
KuasYMdr+xlsXKkgby/Qa3XMHachXOCf523tNnUzO8H55FQ9xjEY8jsg6eWI
R/2q+Kimy9SX21u6UFz/bAKzNmTgjXRD1k3Fawut+4jCQ2/mS/0k4B0npYNb
QGGK3c0GCAFhaShQqO+7LYN0l2xuu2yJMq8gxynNXFHXroMPbAdHybcb2CNq
oAxpgaQRnvL+Tvv7WV3bgbcC59fWb+8ntMy4lQtpD/66+s9AVGz1vel5208u
EHdUbkKoF/Tgnu2pVj+kOpqw21ipOm5C67JAhqvIBfwM8aMYA7js2po2QOQ7
Xa4dWYAL4sDT/BWbcvfYuwC8/LXwad7Ma4HZyLfeWMAa0t2N4zYlLQ2dAD0p
9tZ3edIfEnUrUi+7HdDaR9xATL9vwR+wCjOPyYA3RrvKZLj4QFF2AtOeBSOo
YmQdGvJArw1NxVfk6wy8+x2/FlNUZLXuAG1Y/98+WoQGcZi0YdVzkN/hUpll
dfvnAxnKubNJeuBM6z1crVx9IroDvHHara+NYs/9G4D8G7TlJR4iv9PNQUKZ
m6AH7loWvC7iiCj5eCMe7iGtW3z3b02y9rjMSWxo91zeDSRynYYorHe4U7eS
dlMxEy+0PrFIIn6RsSMKTDyCkxi/2FqNFEIBrFVi6YLxUOv/ZFoTFUv67XVJ
VxuASNVgVsyz/Go1pOAF+lt4itCVDqhC4uhRiPlcv92rTObUBq41umIvy+0i
NqxgKiwUB44GMqJxSxWsumXblF2MXJdnqZqm7L6wfHwcAGSVOyR4sPSpDBzr
XSWjaDEWYEnsWE9AUTzhh4hL2w8QpU20+BUbsxooepl2YJUPb3w9syClaRkY
uxa3s+GvNxpAC0NULnwIBZyMCsZkXn+A7DuH1DtxIGNNEFbMOmANbsvs5LHI
/1GZF2J+z428JxCsRjwoRleTKuv6LliVu0piMtxSQy6yzJ3JHpl7UNdDTBkk
LU3yg6vedwB8YKydgeRng911/5Im9Ra3yUCUUeiuOGZc2dOvya6ei5MKO1Bv
7YdD0EQZoYpRJj3wMQNP7qBjkY4WmQGrMw+PCujhsO5yc67AukarF6RIGVkD
iukaR4BAUbe3nZk2Zu6cxxFeRWGiB6AYLGj6A5H5ScVh9xKo/yor2hGaXY5Y
3wjy7CaSbgs8E9ZzlYUGxzhtbycXKbNuPegN0KKVVpTYf+BfNNpBl2ZC0Y5z
WLMmja5IrgXNoFIBbyxoWSgQsGjdlyljKXRaelLS9e/ztp4RAs2jyrk0zIGw
E1lnMbD0c6gDOBi9Vunljeoa095SWsX96YSCxu+6ctg1poggD67Oolo7M9FI
Ovfy5Z4Vg0TR+lw3Ittd2wDPj6lTfDOICnoDit6rqlPb6fxpdn9qMiYlI0Lf
3/GXRKQ2WaDNJ8LSq3vQaXwaP1i87HSsY2L+7aLSl7EHZpNrcVO72YPPjyCj
/fUHiMLkBHVeDkXNImexSbRl1MpsSuYoRjc6v/I6scrKBJco4Ca4oVstBL5u
s1SY7sVVW5RknuJqYugLLhPWL/slfLYkFJN80XKq/EuOQS0k1w0nesRPc5v+
uZC8GGPTLor4xVFExVSbUCz/lPTsaYLQRF4pN+12muM0wsObiJMEiT8XGwWm
UFa0C/ltMl8ZUdGNiM2P4HPcTq4sqsxxNOdM46lXtNdaOovoQwloefcK4zwk
TgCh0IlbILmNfexJ+AEyDGPiGXVQKuyaMnFEH+WDqnb8XzPalG8BtFAit/km
VzPoRpns1ckVoXEEOc4l0rWu03H9M0yl/qpTFs5ZYMt/TXTNfX6b2mJE+fzt
BnNBn6OOraw77nlTcqT8SvNHg5n0cLnpOPfi+WQJdJjV3mnF1NDhuPJ7lyxm
Uakr3s9xjgkmxyCZ6Ki2wC1RiklWu4IM5UE+ATp+2wbR9gH98buRKtgoIDnn
pCVH/FbivT44jrAtDyXWtqbyXVM/+CjpEDsUD4rsBBg5+8hh3bjk/EblNjqU
dwPYRyBDdTa3zQzSNU8/Hb6pGXTfCAorTTFNiiZBotaQGKMspq0N6sxEpTjq
V3QxwHDOCisqLk5++gJS0cc2TEtYVKKOBRy1lZOaDCj8xdd38B3w8u7xSGqR
rnmQtI9YRat8CowOIB8yx3WfatYI5lbMMdZqtejJ9ah4gfOrca1fSASbo2Wl
rHdhVN0GoWrFqfQEumR3WwNJVOlMX7Q3XaSkwIwsmKXpvhzwfHQ6kDcEbygF
ooOmdr4O9cLQ/W4gd2uR832IMpcUUDZXTHSXV8G0YWxL0KjgQdJZeDvYtFof
QBA6AhagsF7g0F3P8+tARDCaq3Q4e0mP8bMXc/+ScIU77/eF3J9181qH0mq8
+RISU3KtUp6NsO6M116Glb8Isxp+04tM27NqBlSEnzcbqnD1ZHBKpemIdojL
H9duef+W2d8V8jh7lsOcC+nfzlGNybPzsurHHW2vA6SAa1VilgAJ9qj2xUAZ
wSYmYl36TwgZgtBW7JCNej8JHfbIWWlc9D5wSVjujyddebzd7foRbGCBXHcj
dK1ee4nSgnQ8iA4S3uRR1Jgithv/9Ew334kkJT6piGiEiL0CKgh8OTRZv/zl
Sy5GAqkT+zh4TOogNaxhnAWoP0EPxlqhZs4dPn5NVajq1Q+hPDdgLM/D2DFl
iy9ZDSdSMcaO0y0QbzmBKEcN3u+C3jZPLeTh5CPPaMX3t3j3A9OP3bYHgoTV
hH7Cuwg5+lA7PkrXGE9KcJuHB5ZysMpB3YcedBMnUBmlXlnIbrWSSsFMFjNc
k7x2uiqPtBwhyFw/Cet0I2tx9+ZhwU6IWI4ovR0OAtyq5uRJTx+7+VzHB67m
EmfZymqDQmkFTBK7Ymdtsx8jfB25pO4THn/xOV8eja7z9mjglxvKybI6Z+nI
bFpSRgcwowKBc8eTXD/a4U4eHWB7bP5jGs/GkvaY8tcWz69oqPUL4ui3UkEE
qkJLSkn0WSay4I4dn9SlH3Utr9I7wC+wDdpNEq2KgUJwArJ85f9iAD39LNFb
uTzCkzOzvYRpKOfKsCwOX9NwAP+0/YyAqR88s5bF2I58/3Rgv+NFUTsBNN3X
ACFnyzbb9g/XhtMSfMNYZ5qBYILtwJ5Vjy8RlKM7PqMb3Cc2qCIZzDkKKtwG
tps5P7inNO1u3pFeg7z6F4nvhrfrbAGje9GgGld0YrBUDsWsDijn6d+hhAbM
L4bbZN1HU9OX6bYtSh5efdnvD8RZkbATwvQ0IEQZVf3H4C4IyFVotlDjxgxI
HUgQZAOgPS5VMF3DDOcEmT+nsO2+BIojfnOwJApgRr2cAXIxYGQ8KOr0S2iJ
F5wgL4zFfDOfBZDPqttLAKBUCmkRh3Es8I8d8i/P6LLbQZdyibz9yNI1/AQ7
z78WHBaNTeOpshJArfXyYB/Pj4PqS/qy+bormIHXgzVkr6VArsGyvvUtkWyO
iimzGrsq5HiwbhQHF0SAaBZGDiWvZ4uNPe2igpB03rcmEisKLQS6/TyK+nS6
dnWzdG+YftNbZOeHAs/IwxixhwMM59Dy0nWUfk1mjAoTpxb9e99QGRpCAQGv
aA9QGCW7GEkue6MFEMK44BDfQC8jGaH120B8G9fFyDhPKSni8/1Ajx02gqGn
goJJNsACiSBDE9trAw1NWpRx0Xe1XkbDEimBU8RzLLcYeq1apuyhP0ymjYz+
G3mpNYz64VHw8phwoA0fZNF/ptYLyW6njGiBqKjUHZAfNMqb+zMIwphP91M9
z1UaVg/DEVVVvX+iAKZkc/hSxxKJPnfYsQ6Q/HLyr+jvbogqOxSJDdp/309b
mzbsMFhbOx5wG3JMVGREz0w3AjxseBTeZID6AQ6X87Q47wpgKh64k4b+Z8NN
2DQKlF0+iOq8q/pRQHKgyFNst6vGuY6rpfOOM4p10iXRKNWbnz2ZneCIFHoK
S3UvrBuN02dW2yTpTuAVjK8Qq6ExJIr7mcYArdkLbYTNAOJdId+F6UtXI1nS
rcznMMfbePS98wXlTf9d1hueK/8ZOsPD4Vz7fRBIomjmOhLsIbFF/P8x8VME
zODRJfpyNU5SiQ9IKGfu5QcQJiCf93Hv7j5yHuKhj0CGfWrX2L2l+80vllrp
VtmM8QBtUoeya/YNg5EZaKby6dGLWFAofXBmQytcSrwGxVLbcpGrhadM+pW0
ZrksKTqpTX/ET/qZTWTDJSh2l0A6QOJ9WVfGioUlCQQu6Oe6X49i6Y0AuqnN
zOjk+Vn7XkYtyP8kXwr/TWVCQoVe7HxfJPQ1UsxNp4v7f2dgrZse2mhKnTLc
hryKiaeOq2OK4Wu9mhhfK5skFN2x7wpq2y3BsH6/2R9pgJUCt1+9ROUMzYdC
bZJ9gh3/uLrIHQrne3qOk/N5WHuAU2uzJpwyGITgAJS6X7pxZCD1aDg3irKQ
zmLVCJZlbPZHEK6Rlx4xy8tZ50Mk8zb0BN2abhx+mQBaEBMTZhV8Kto6wD59
ZlRkuDau2TOPkrwNAj5ekDPOnVPA58FlfCMZq7XHqPQ1GLUtipu7J6eGndBA
sOvgRtK1iYg94k+dPYGOD99MMY06nmXVwplhCW3Qn9S6M0lvziqQG7hJyevY
inAJMJ77YKXHHqoH1nzxeBXUfNnujoqMTPZa69BG94FqKYCR65SbbHc87NR2
sdNS6tbIUCZmgDwD8z1N1Z9Pl67XGyBB5+UfX/w7xFYwqU6wfkw/AA/2ZEq2
r1vB0fVr6OUP7M7SW5nTtarJkmjHTCjX1FTMOSycTA92jkkIgWfDXhEBl2et
kMPXTAimbE9JOP9F7h5W0UR++7QbqVxrFD5BHpqrdfqKIZ/qUGyqcX3eOAZu
PNRRqXjcWzKFkDyxYQcRfHDAEh2dng+3wOkf3pllnOG1pKGucGw6s9sLFscs
Na5AD1ojsUSa7+NKxpfRuYkU+gMgBsPtjJuljBhBLCyXzM1bOPTEtlBeZqAk
2E0uTjc2IIyQM3Tb/TKnhQfFgcBMDkGwQ1+k7clVRz3igL8f5xL4FDmrldBD
BRVLKoRClRzFc1EM2VlLm8ZreoV1+xT1+mClupbOWIq3MfHjCCSXZIUbk36L
U/n7t6AwwMQtGNLjd6DofkMOrhrGm7Uh9Cyb22otFW+xOr2HtrX7aqM32jw4
FZVByUIy1RZhfdRgSfQRQor1xBWGu51ENMm6ed0SdE+goNdGUq/I3olDjprH
vrff66EeEuKywXNbRDdYYrCoiNjbiqGvCC/X+UzqcogQNqZMaVDOsE3V1nKo
ivR0crOSw5oZy2Mrk7u766ZfdpgbRszOGhnlam3Ig2O+e0esSOO3NtOmM88f
ak3tMAaewRKYDqXYY242wnHoMKYg9xZvluJr9E8rTz+YCHK//Sf4uJEpEaJQ
1vLoDSgEO9mogTohbypkIFzHUB2myJmg7O0JoXn7z1cuoCxMI3IobtgEWTaP
uCAu2TttRUtG2F98IDABKE2gzi4jZc5Y1J10bGUpONl2Ypef/fmP+6OR7lTo
KkBGOCfwmyxWRFCFPgAhB46Jca+beTfown24zOCTeipeXqHJzyZDQgLCRPmC
/MIDJaK3/uRewVTVnVz05/kVKdZjev4Sq0PmssO8MKbmLOpZQvkDKh8sc4+i
fhwvSx5ZZ+n5LB+zLPlI2v8LmQtWpq9QaE4ATVoskJ/77NEaRlAaI5KCHmGR
/2khknG5mrHTquRb7KiFqV5rqUBn2RCuJNLvB2BJKP4YiSbNnnDUunHWDkJY
06AoIuj65NHJnO/7ydmxv8KQJgPwY+4lhMzxilOr7jTHBHX505hCH0SdEUfu
/MUNpV0tym8zjYXnMzVOOV/GZTeOCHphSqQGuu/Qh7QHHlAHycYlUY2byyFQ
hEcjH6H6UkaDOnyeUj6yc9SSc0up9DLiPYKGkaMc6YSQjU0EP+QffobcSaFj
5BbHZlJB5iWnRVPBvmOSS9NgBeWWCJSQHY8KaGTfoyyaLF43vu3mTfNxVMwN
ra4UomjuI4aTGphyEaaIHDdwvgN63MEMI/IGmVcfpY0/zsgnTt+/jYdP25nv
v9ArXubSDzN0P9vTdcEzcOkS5Fy+UO8dRZKjcaeA3j+sWzGx2KiTCVm0Oeqp
ESMslimppsg0A3aQi7YVgzTrVIci8pNawHbBRM6v6mUgAApoxZioXRaO+8AF
0LiDx88rQkG1Ok81v4qmWXmVKbYA+wyl0JHtFAijDBnuCmhfpTnOiekdb++d
lPOPy0Aisur/bmt/a3q8lh9D78Nqv4sYAbOxqp+nN63vyjIH/RAZLVZ4svi9
ptVpAmm+CysewCWK+bM78HVJG7g6F7Vqvfhb6eNsHbKn9Hl8V0olHye2w7o+
yUhgC/f+tY9hl4g/0f9rI61UHEEwoNy4aHzIAnnT8DqOGwumT1JfeiQHJlGS
7rJRQmG4tl0Wu9yOTwHXVL6b9jF8VXV/bw9pENLmVSL/D16uJWLVgd4BP6o5
3hBstd1Zbq0u0MZPa8gSEsHuCKjsxzqHb6Vn8U6XFE/R5d7bq7zcQOFB4vsm
xI4gGYG8CGUH/SfqB+udgMHhejXYJuI3D8CT5jSxYS3ZBdq6huXCZ9tUcjXm
DEUZ7YoQl0uACU12eHscIFo7F0+ylXPaujbg2xItXVdZkthyV7FqAqiL954c
Z+Ypeq6c92PKYCa4i2ZOMbEuNJc2pUgPp4wUuehC7KLZ55/ZmZzv1X5bpQhy
NMyYZ7LK/asRO3PrOhTigv/4wEIykIIF38uDzEQpFMHdWPf5oJUYDylamdzL
mCPU8B/jIsqHsaOrGGceDDE8UmlVOwVx8mI7sF+RFg9IJfdexcqdUvPyCP10
XMEVkpXFc7eOGmKtj2CEkIIxoNqfTECx8m335n/elFqYrLAh+ceF7YTjRXqF
aKn4bJNyt2FVyoJqwpuJ1E1l0sS5uK6+ssmBaJroWhjzALAeIT011jE+gVrA
/6c/LSh7mutktNswtkF2B14Q1jxQaKzZ/087Lqe1DfQLBfYfGcRFxJv7/v9U
8IJy2ZqWR1iIvzEuDAObyMSyre0G4XmHnK9k1fXn4JnOW9pSh0ev45iqayg3
ujRqfybpg0gIVILpBFGlFkpP3K4E4zu9Bp5gtwv7g/Os8IXUVt+Prrt8jcnj
4i8JS0D23yjeB0ls2vW9mjoUvtM5xce4N/BzxWaGxhyuIbgyYpSPgCGCZLm6
2iIxFeQvwQglRXLbAviI2tgBqykdRuYbsrLGl7wAh0isYPhNnuDCRNe2yd73
tpKyaSi+gcITc6jLCgRb5N/P9e8pMdWfH36vSwBr0wupTCmrxDek1FEaijw3
Vyxeo+dDjvvfspePkKTkbO0YCqg+AZGhJ7ap3QrGYLidr0e0TgRy4YP8IDU5
MKhkk89xeSwXgtCPlHF+4bmtnp9FpbTp6326irFJ/ggYQ6SHDvIGhiG7lny8
OYuulwywTJsG1VK0qULR0sJUktyWQDVnN6IMKBn5kn8Nv/1HPgUghbH/2UV+
2ee6nygABlXX5AkwHdBwdPwRmqzzqfG9lPN7YN/O9HQLI91MjbnGb5b+RPHu
um09n8GdniABUz44GmZW1MPJKqeeDCOzBehPgOylYLylvk6TeRKQpiUWXPRq
Ux5LJzxHZi0dGEAU/nr8lJFrpC92RCIp3oXfC5tS0mnYsooMe/Xv4G8PqZai
gSzeZfIlJYWDj6WFX5ehvwBQjErOmZSsdoQF7jWK2BOguFos855vjVR/aolL
VTC8PZm3Mg7AV8mm2CYO64m9oWFHKCM7RVlK+umyBykW2nYLLcXRRqQ81aJE
d9F7d9FW1gMJJCs36YIp695BoGzfN0r86q88wn698cXvI6SDmY8rIfYUuo/W
lEZkqrf2ony6hjZCw3gyVCmIETQ3KANY8ZqX7TTz52DrTgvS10DNkPndVjPX
w0vFwcNQxI7UDjpXGH8W1COVqKpVn+HztlISsz4W9vhOWtD4mHKM5hgeb3L1
IQGFEf/ObVQDnYdTtzr4zvBYQshDrD4xLkBZ9hcDrEnxBJ7jJE3wkHM2NkcO
2jpw32zafGCLsUCHHtvbmdS9I1VhRT66ZQNhZlVhxsC6PmAnvDvxWzCc4JKc
L8DpVM4JLOB9uD4dDjGSrKRtmaRnmwO8Cx42wER9apYhwT+JtRkATk1WU+vX
aDaIvXOrMtHvTjr/ona8d3w5XiGfq7/Y2mdsMy7ftYFBovaYBESoVa8M0+45
s47c91EiiiqD9cijJyCiU2edXMEIbihHR5rM6v33ANhbof1FMaFhgDIHfbCF
YsvjwyilwTo+khld/T0ePFDxB/hMbXitgxTvfjsMQ25aX0DJ5ppkric0+AIv
c2ic7mDaMrKH96P9A/I5spqPWbnOz1Fr1/XinmM89b0SpNw4lbW3m9FCfrtE
cJCJjjWJ+RYTZpUZdndEH16LqZo4Qxn8CDci05bbCvzLV2SxUPlj+yBOR7O2
z/4KZ4DzB0mPmuVYGR0gcuSNJl+yyM8v39XYU6gTsLKDkRSlwvC01oRxeTMY
UhJw8dkmV/KzuEAnXMN0lL5JwAmE8ZL0raaS/gfT0lz2UEi66hHxuc31Jo8U
vfVTAst7/un5RG8pS6DX3wh6o2NjsfALILIi0YFtd4xnyj3afIVGUlWvicXL
ajy2ta2Th4WTs89jECDNtmx62mfOZtUG+JtJHxQqE9yySxcpb+MP49e65+Vv
jpIPCUTM2Dp18Zdi2ZVQq1mlcJpnUhCZ6l6FawXCsshBraHOPNjYswCU91nK
dWx6U2XOknsKOckA6gU28QLQ/bN9Es+UNwKp5V5/eLx2aC3qKWIdaC5qlqnz
dgKwyK17TAxDB5FemfwW2za9BJL5gtQcGcxkTodLfiO3eKOgys1YN7IIq0Vm
aoVFuZcNhgYtEha2lAV9dgvx8dCCufkUetkwqFG0NaJvV0fP/8We38NgvNFb
LPE1F4Ja+iMrcmKuIzqSmudnXcJSJ45pQ5a0rxRLdWzUG1B7za26fS9xRVqX
KoS+L8s03CPv0kf23k5rH76m2XGeYdw6CUfeE999NWHAv3GSU/Dx0hFwrb9i
46IrB3EKWrYFd3T65bk8gikJbHZZfMgewbMR1CkUQArBdXasWEp5wHZnbHuE
G9ZSl+564CXLT/5ZwJ2alHDoUv8hg0rZpGJomfF9//eRWqTXmCs0LDfyBa/n
WAzHhuP85D+NM7u2434D/2SmOatpVw6SdUPP+CIQ7tPw2hhlrlSN2r77fe7F
Cmino1vOv/L3u0tyVLXZJuWPmKYPXlniW3mPvxHwm7pG4wdL90MVFoviVbOX
aRgfOBzmkAl+/+E/dFTTfSFm2rwBhHs3wRB71ySJJn2/E2SE5Z0FCHeGyiI7
BkxOdhhIQyNXfnFlCulAE9Kf2+trQGFS6E+3gwdmVU+pDa5REVOKtXcbsyfn
NwkMFCd+H+TV7qroISyhc6+frAxZlxzN6P+ttc940TyQG+qPloXVEdOsOPRM
vuNZFa8DbfSiERYOdI+IgSI+chimDAYjodO7TF5sGg5mbkq3Bcy0RVvnTU0Q
2TGcsLPO3ZQdqlQj2AmnUSK+o7HGzRl0X4KL2W0fptaCDoWoLLGKAu4gaqyQ
/ilK1KqivxUe2JZxPWjvHxqxiNFSzb7cT+0HxyAncyi9izu5hTprqwvRzJiR
0X+LkCgZPhBChanoz6yR3fpxQFYdiSi5DGeVB0VXyDkwBFyIMFkpukRlIwaj
4glZPWNhYFRx4b2E65smXnsF1zI2HyX+DHPV1V36UDWis8US1oMuVztkvzYE
KWtvX5DCL/LewLZl7w0Qg2iUNH8sbkejGtzWkhJC2hRPYiim+JCiVuiM71or
d7nZ/oZd8d2GBjnAe2DbQzAHJMz2zpSiaggsJ4Qy1VbCtIzhyDCilhZuBjRY
NM6LkeG1ZVieCQMUxI2BVWzLh7gt+OXB1hFHqSdnSubEVf4sPUJm57EAiPJw
hnIJagI49Z06Nlk0eNDkNaOHzpCKYRiYFSD+P7AV3w01aplCR3nbesLD3J8H
jy3/Iv8aR6kaAmsJJYYSCiCI1OBUX1otxBKiUp+CC+vpkb6UHXQVkRuvCony
OrXCStygj2hPnZylMfBx64vJG8j/v1QTw90OydiqoGVpBMlwzqkuZTzfbUpj
8cMggt3rVWTqWCaeIQKjrxLpi1XRlhB4dY3O17+lMB7lb00p6aERChuXVH+A
c7jLPF+gxsNqw0OuHdzQc5/tYPo8XpUdy5XNVeRm/5igSgi+RmYz2gJLqJ80
QfbjCy4gFvQCUUeHbJpGUuMqTTTnpsGVO10td/zo1HjoqVTWDKlsPQpMBlv6
MvsHMudWDV0rE4QWLq9hDCtDSgIx8nsyXdQG5Iw+MZ0boYQIWKOvdYClkrxW
aRihmEqYF+dPPGSBB3bQBmypToQ4/DlVAftbE3CtY0SsQjWr4dC9Ob+bBO5p
T8/SowrTFedXZkwt4g4/0+QI/6JaMiAsNEMIH/nqZnLpZGTa+LqBNZ2OQPRI
7g0k8n6YCODQ0AUwJlDxssIfxrXhRxhueHoag7GaGNAyp1J7lSCTKZImobXH
TFIkcre39MLWH++NCO+JAtv+9lONynRxS010tfgel+jR9CExXf4mzGIBm5Yv
1V2jvVjS5ythPs/QxVohkeapgNj1L1yODWdtNxQbPDIHTxQONDNT9AR3osPI
n13Ke6BPK/PdilRXUnSWltTv52ax9H8DzctWQjL57TLnyToLMOqAs39jhEJW
yIDl6ub9zRZOFdc84cclZTyNdp3oBy65orKeI/PpXWEZPB+UWi9bdAJDbIBf
bEHH3nGYEJzyVsqu4LrUaLrKfyMgfxU8jMZb/o1nB1q+51gtoyNxEZjPB+wx
bum7xB92anF+U9EJ2F2t+53LWfO3R148AeSVWdXCS+mQSQGfRNxmdyNwKmL2
OSjTudODPWSVpZ/ka/+0sOXIRW7OVSR540XWQV1VpsQbFw7hpppOwmfq9RSa
HhaMVmGueD64XkBx9VipxS/eyEBVrNOi7CwevBDR2fV67odCMezT1UM8vy/i
3Z9++GRgkg4uZ8u0fJJmkwPWXKE2gmyrU++lqvCDsm1b8wjvYZ6vz7C9nYad
RwFJQVNvo4DgADEMZEbGx9ZO/1lnf3VkmILVQvZPcowem5Bcc/riFUIt5Rlu
cKlviGCkSlgYZo4sulti4e/6skvgx2QUsVhj5N0A7zbXsBufhKYfy0ntn9gF
7C/aKyNUUDjWlaa9mEpSdaKrY/hmXPzl59uzY9kNtk1UYBS3NLf3tJHEn1On
+QEJ/F166arT7LfFSH0ADKjIPviNhgln1ldTU6iFrBJRKJg7wg/AlIn7+SqV
lPJciWh5XpaKSMrRYZjPULi23HuDG47FfFROAXUJtDHjENJON8ZGHYana/VH
ayXGZvXp5BQVuceEau/UHlyocsBbVeCwoyTw1RgHS9NNq9SYXg1K6MCCyxO2
oOykt6k5R/22yHAZQxUle8vDH9o5CISp9Fa97QFoHstuyVVx7cREqV6rPPEp
I+Om02QLe92fVBzvjoMpPo19/BqYpAJzQQR0mghjcunZUN1XpJ+Uzgtysoid
MO5QMRDqxO9lyQhNcSpcu78Ao8bq2sFAMeObsaocyBudsPEsxYweJTOseBq7
afl3DfG+5cCTlGLQar0CeXs/vCi/FH5HvWpG1K4zTPRblo+hJSCv0mgmuekk
A8weHoRsnu3fi/1ZdQCDEobhFXE35CkMq1BMWgKk6Lb8uRKv0eAk0isEDwhb
vl8Nf2hA/rPQbdtIYE0RJvrbB2xNDmfhFVQhyBFKYa0pod6T9y6E3jImrb0o
qrzWlKhxNsqrbw2rNuoVyJCUlCBAmRcFrIse9QIeDlndvx3jHaxSE+Hu/g+i
WpFUBbFDR7UfKwXVTPSq5JjMEADHcKqjJq78MqYKph2oT3kzLqjuseSO0A65
EJRaUi9G/wUaYjjOM+LJe5WjBLnmOrxd+K1PhHSZmHN/J85Dgc/dpSP+04DS
jT0R5QXPhI5vkcbM6OGvJ/Scr6xiwZXfXNKOIZ+jhAPpWvle8Y2Vw549FguU
FVy0rI/cHLqUkJS+Lj+SSt1M7K+lxhqXJy7YfTgsZggTsS5YbQqqC3EbN9mW
Ienb46n95IHhJCzs03icXbB9RTFwX7ebBZ5C4B8cCWgqwE/sHCEGga0OxlwN
asDgBr94/Hs6QCZDZyjbFNB8MbTBn41ao8naTnjv1brL/vukdusBmAJLZY+4
SvyTtFGOTAusKfyCUmfQ9RMJfWDEB8xa9remaLWczCMxqNQONiKIRdN7GV7Y
BGhalBPORWwAA3S2uU9g0fWKP+MsXoExGfAkatEwKN5fEd3eviQVrJhH+ygU
z+1jOGXLyruGhMdHgpa17M5TkdwMiVKnbSG/5EC8GU3qNXWjK+i8oU9/jRB4
HmpAhux6ZCx7ReB8r7bzcYeaQDiYxxDtBhRbo06NCDWggTgvj+pPtuxDe2ph
EepAIQ3c2HXokIOX6f11zf3YY2k5qaLx/x1+7ougzuykiDbLd8Bz+o2VqEiH
Fb58MW/idjgraR+e4b7PNMMwS7uox46/NuB0MgLlLmJ8ZiH7B2u8fjmfIS6b
rS99Z+ZJTiOUoHuo+4Wl81IV0H6R3CXpGNohayDYYlRK77BXgOfj+mnomNgi
9eA8bWgs0YtEV2kSMNtiS42ThKLClqeJ5sLtzzoeeyJRXA9Adldr/FyNzT39
geMMM6LJPW/GTrzjcigYF7BrD9VTcaVa4GIDiVcfSFt4nV4RO1cEoRYK7fBG
4a6hEj+tBxmE+y4MseyfegzmFVtSInwFsBONIym7pS41FFOtdJtkeK0CbKlu
mMpalumKTgc3J73QxXMqYTpm1o03/lSGfRRkygOUnK9citK9/PHucJEeS9RA
VksaO068k0BISJVmbqn7TjkbJvf2XUoE9PeyeMcZ8qickKpLFrQF4Jj+VQHX
O0yVPSk1nTDGm9Sl2+qXTIevJZ0ccR7EWgmOqHi7MKkHI5a9TZXZ909SAcEZ
OGGlYspC34oUpF+QBybB4b+lw1GTEcVIxcUOAH1paOTqBl9KSDwtGdFvtL78
f38YzJ64hFY3J9+9pknL/qfNawwSwouxSSlxdOaXqyl9MqGGERoVa/DGl4aW
SJjfs7DxNXV19KYhn0aTRjYa/giPEelpJNk18TIzMcN4NwYxlJPVpbnduHo8
HeTTrSsGpfHDPsAQgt8358TE0sZpiHFrtjGhc6GaRfv4pejNikkFV4RE+BIw
5+QsaOqcbHsgV+NXe1OGc4z45IJEm7zh7tBR4RDCNo7UNvuW18s3JflRlefR
K1g4IhuQlE0Q8IiYYEggG5PFe5oRYgAifNfH0JBdV0jDc7iFuCpqeIYwLb/M
8Sht8MwaEalTtyBb6p33K247fXCCOLHfopPVNcOAn+/B9exNgGtR5ptQAhq1
DG6BT9axeBWlIpyKVqmDwlhzrVz2RGA8RpNKpc2DT1GUqOL9tdhBzlgOZDK2
kOWmvyzjZTmtigF/qRpQJAaIcokj+LDsynXYr4Z39OWoSDDqFGyHYAjmm4Vd
0qjn+DbDP0YcZa8CRA8TfnU3115tf+6FHI5ctpKOpsFPCK96ACwccziE4MwW
klhiIzunTzl8n5QKaMuPQ/BRJQEprZgYnGNFtLpeC/nja6YWoUcvCzHKKj1P
3tpgfMb9L/s+dDujZonu+U/oMUBWiaLGTGigLmjJeJQhAiA+EjPO07b5X6dU
QZSJMKwUlk/XBhFEvQTeXHhfJGZ3M2iZE14uocmvncyu+uz9trsyJzLmmXap
DymY8nm4pGOeN+q44DS5Y9yY8GP+7tbLC68nLA/tkPD0hlGmUrjiyrPZ/zND
0NwcKlCnbylIVSEEwPe0abp2bQSdNuI8HICyjkhxz3SWEPxJXIEdgQDDD8Xk
4x80QTyOSU3puGr1nIkj83DBqH1i/Bwkel2KLOFMtdzdppXxuTBHdxWvAlyd
EtZNySjglUkt3NCQEmV/mOPH477MUaTG2iq39frLb1AamLCmyYwNNAiNOXwf
GHBJ6wXclnzhKl1spFGAH47VE0e+5QyVmLl588b70Eh7T/XxX7OsgcYk6tGq
8TnNFhE6yw4wW9yhQNw8oPaTelQRTz6EESTZm5mPXvDrzDidFIBfbJpIULaD
pGQkq4KYaXefww1uqgGjqDyftuRX8otZu9QXaH8nBmZrm2ezyyk15Ot5/UTX
O3+IB8UsNEcNuI7lKmkuEIafLWIN2Ef+Q0euOYBkNvTBznLn0oCi9QLWll8T
nFhAvYsU1p+JxoOAHz4YlFQMF7uFNJERQGpwWfrPF8CjJlpFgCy17oj/R+P4
C/QC+gSiSzwdBQoUDStPXCTltTutYISMqHkUFHJzDHHNWkB4c0UWgxUCHCQG
IAggHz3Gi8aDcZobHRy5OJXbgAFzEt0A21PY4ChVr/Rs8U2PqkW5J1sM2C9l
YOwlHMb/yHfCXKFp3Bez24Q2QmYUODpZ1+eRiS/dHI4ggYrV2JBbARgEHdGX
/9F5zhHuVdcE1DLaNTIj64uciJMvos+T7uq6s44vMZUVLsLNOBUwZFTeZ0ON
bPjKpuHq+3nGMhOUTPzoQ2vtlnpQupNuYMkQjnuTJaFSBp5NT2be0vj+5+hP
+ZTMhxpD1yHLgO+NrRLPnIIa1jNqgRuYaz3GailTInM2b6Jt9UJC4yO3ytUE
nHQVCpm4GvkwO782xfgcZ7qWNCzZuL1LexJXjOc0x+2TjnQIknwWQa2Uw7ch
5seLPZr7LGqILQAyQ0EbvLwd0HRJZ+yrdG0J8+bXZ5t4fTX93HGT8Vi/50G7
ved7a7dHXmIqMZN5OeYzUgBnDuPQMlrvW//djJb1ei/9e9ZKp0ZmmwR/Ht2U
AUqtOXLOd5bgTpdUGTg+2os8P0YRavefMHsASAEkAxfGv9vsnx3sIziPdEbW
b16LjA0RPuHRrEtfNb74Kz7yv1JuGFC4XBS/wPhBZ9zHL+DqcTaVgX1jzrri
rMgZE7asNHKqHx4U25sZs+ytkDOjuui6T//2J/252MheTI4D66+QngQWL1BD
RAk9ArzuZY0D1ekgP1gh0FY7QzqVPiKRS8k3MFbF3a/nMWBgMU+mHikyWLbp
TYJpOIOurVgIRP5W57RypeE2dhUi/sfeo4K0u4+qtHNQpaWfT4yis4dAUBjx
atbNUmeAHBNSE3Dwe8kha1ngM40RdOy1owkMPuilf9tZKdfkEmQpA35v/QnM
uqUfiCRJmb9rvfjqIFa3vDoKhD+0jS0coKUsyq7/hCOjD6J32LIDJH5Kssd5
x99TUxPGGJFWtJsD8kKnKo2dGuAf21UZj+bh49/NkyVaqnvtmcd1ioTVJaYu
I4w3gB1YKWnQMz4Z0O4r2djpNDumTBUcxNzx9SPrXcH6Uvq35Fx5y67Dwzk4
zWATXHvWCPlDYtZptu9cjXmOQ/NQG0q2K81LUTuLDnMSWpTJb6T0ugpxS6F0
gPP5RoqmwQpNMe0jmXqmQrxM7mZcZ10fN45CVMqLakVp1nMQZ0Xnhaf9L1E2
I5PKi/4kJNFfYqtusnavDJqTvC3wzMXLeVpmn+DUw4JCH6cIxmn5hCy24eqM
LeDfhgL9fTlW5nxrcgFvFfP73Dp/SKigVxOr6ggiYd4uEkCVSkybEn59SfWY
pU5YN/K9Gbxf/WKwfZRIUJwe+NECIkTwlEQEmOfqKuWAM6MVcfuPisWTqD/m
c/FVDXrlT9eP+R7Z8ZaFuAxe5Vtpbzfxwq/JFs+LVhdeeJMTEIyLR9WpYmWr
4x5cLUotF/IeFVQpLZy9WMva2mB1n4w9FsOyphQMVm6xyR9RF9tdLDdmqclz
8P3z2SOJdBKhXYhSXcWRd8l+mzPmEwItDuYgKgNXgsz/eB73UnEhDlm8A0oR
DrsK2s/q37HADOrfonF+EKZnYjyVfA+nGN6Mln/lHqRANmEPQcEiGoOe0+TD
jrTr71Tu6MGlqdA+2oXfUMbKR1cnT+eJTNsVbc3oItu553uiUyowONffCrRv
qsbB2y5Lrctys5CfY+T7BdA4ucBZ8IQQNA4yXnF3GUoui2R15Ame2FaoRUfE
gymAqDc6HlomHzf6XEbaAZZN73Yr6V/IkVEOHW3artsL2v3cj9wvL4UEj1N7
blu9J6CNXO2QaipamJn9uhqmO0oOwTArg2/PO+JZuT1FO8KQFbkR02EqfqBb
YgM0dSRIvrgweRzmJcY7cUyFCnB0g9Jj9lj4x2B7rCoDLhb8FQzA2c1CA+se
6QB12DP8y6wdaYAYIV/f/5pgI2e1NlxTGU+mBxg/tOalqOpOjEbf9+BuV8th
YJU+JZnEImTKq1gYvb4Gt1oxWu2iHdnodXDOVHXV0ah7GEGX2xbUIiSoy/Wt
3LaGeARANfzFSoNUstoUhGvkfkIJ24maLWUqUIm4KpqvJtAPIw0/JtCxXpcC
eOgBRCHzP8KQ3aJAXRFng8K7ZUMCRBQuLP+KhI+eR7BWCXjuroEV/19mmC10
MV8iEf/76LFl0wJk4iHQAY1wvk8yuveBWjGXarJauQ0eovXPU8bRAwlfdSw/
LK2Q6b3UjXSouoWgOl/AuKdpkkfoqDGGI+yIWshfpE9tN4NGHR5PAXKxQRTP
uBbsFC1dI4I0enrqt1wAeniY4y0BmQdtd24klJw8yNvi59tVxRYyI9bRKw2A
Oi8Oow3JvRwNRyIr7bGDXPePk9VR3MH/uKa0lKzM5se5723LfNyCN7gk44tn
GbLcjZ5ll7XLERWeSFVVdk6gA+53mh14mX0KXiR9VhfX8xA/BuZuI3M3rPVV
R9hdSEX1rOZeK+v2yQ5jnb88S3FhyaUGZhpaxNgdD/IE955n3/kIfqRa2uPv
c1EDXCEVgvJkJQ17YNG/ILfTrpG9qir/6+hMPLddcGJ/DHbZ9N+2mQ52QvtY
vkDbxSS2WIPwIvYHcyVuNAGarR/XuG+T/X3HmOZtBPVnpcdcwFb0Y51WZG9p
icg3MU7OKbKhABkNiCmFSyOUtLLuIfvwN0MkvHAnnwH9lujkUUo7O4ZDL+Iu
fCrsGbaGYmMbRS4HVpvm52wAObjQt7X616MivS6f1NpDyrbhv0QQsaOxQRsS
3nR0NfP1Y2vKSKhMF2R4z38+PyWqXcikfVVRhETAUNd0pRx2EWyM0rXCNK1D
Dnd6ijHM/ux5/dqZqDvgt8EJB8Obcooa4g3dZ/XpweFjO5JdtC348JnvZMsQ
8px80JMMRFFJqIhf1g3VCK6qxEOrqUvxODouPenH/aRNXhmtCzxVvb4VRvea
TyjVywjJ5XPVapw+fsjjlvnXqyKY61KbR1yTdaADC6iCWbw71BZjv9aSBuco
vyB3glarog873Y32FY2Fu+aby2xARAls32XOA6T0Ky6xLzoXgt/00UJ30RjA
mX3QoVCwY5GXrDMxNl67pXO4Wm9Su2xmB0I/NVW897gqEC9Jg6OHTZeaAQUl
w83mfFyuJlcPLPU58keqJuijmpXdWOcb6ZDSkWUb7Az8rZbSEMdjjrNpdx4Y
IxBAPihdrZf/pm+MeKhuwiLasNaTXlciv0sNyy8i+kAJM7pz/BE1KXziOK0R
7ajUfFqnP+t3LPeCLvXGj/7Yh4X26bdqZlV1d2/sew5qJQX2EP5J3FCgY0s5
nDXiSD9BzmLzv1J+oRClY0jDSmf+Y1B+YT1pVCxUx+5yaOkOOl9teHUyiBvJ
0yfiYSdxsFw6S/gVzZY+bmzcHqoSWaWGuyCSKGouHqtPhYy+lYB/yElfgGiD
B3JfvLq/ZEn797zPHxIQ8NloCLoMJEMMshypMRTNzu7+Zf04BHb+zHvnGhRT
HSFYnlBHtWw5mYix8ntPXW6cvjESvC3yW9OQaChsCtcGk2pKGTklggO54mB7
zSLW2Jghl98OTIAfcCL90pEy5novxQpKN5jv+gsMolJDE3np7F55v7lEs4+f
9WWimrVk1JAux8QBNOG3OnqY8zRH2FwKkol2fVDbeloK2RBRDThiToNc4X1p
711EVfHvOUPB7eQcoW2usACVEht6IfruRGTGFrxOKb3YsWlvBhRBMWQ0p0Pa
SoNqhQ1ZZv5HdLDXRr3Dl59IR+C8ykrb5ZcPsjkn6w/g1P73tHAphfx71q9w
tMBsYt1mt0tNSV857bqFRP6I9+4XdlzjXOL7fEs5lLLYZfyY6uVSBfYXXjoY
aY2wRKV6bilWedN/uOBxuTBOPUBo7uH0QJvPYU6EsXsz7Bki3e5P+I3xt+BL
LPw2FAyxOPQWJkI/MiG+HXp8qoWHRCR482AzdT6Ta/fGyF61SxsT1Kk2nPLc
P9O8FpQ+S1kblbVRHx93op9+71Z30vITmG6TQAH8RDzertokIO5Sf8ALuKgO
ncIsHzIur/NvEl9RM52EqzInrLYftJaRy024P69QOl3u3/WDEWxDUiNrPsBt
KqtQS1Gp6ky2xvWvDsCV+EORmCaPsvMMZpKnKe+KprkUTPr32V950GqPQWY6
pfwyGgkHynfmDp4AmpKXlDs69bN23crWfOCI8nsXHwq/9Maw3LEa2eloSeiJ
S1INfM2DSici+qLLTJlyUL3y00rSBwSV3rWTUzAn/2fSwdM+rS+uXoTPdCEj
t3wQyx2vzwC7KQsSlns0WW5fGEVKZUyFeRyfLRe0YhGdueKwG74WDxzbDVmR
dN8bikYPHBONGWiiUTjhPmYMyHPgIEQErlRyP3qDgkN5WYojLHGAJe+foEE+
c1c0xAuPvh5sqAfFF+hf+WbULpKd1dmTnfWPMRblstJDoInZbPwrUxK9q0lQ
PpRZOaz+9+N83yonfIjUlAX6KYtgHiFxKo4DuKARSt2V2yLfwIZEv3XNflgd
U4EayNeq9AcE2YzXjESdApwIqb7uIru4601W6Vq1hFqdOi3tbFW5LjSB+58b
hHOMvc8VlFqbnHv7PtBQb+xtl6++4RymAaRFkjQ5DWjX75KgSWwCKmp8jc1B
N9m2sXSGBbfSl7qc0rY97A+OGxmrVIPt0qacXz2qC6ZHZmgG2dGGkqv5MI6G
L8cJqdfqy8A+wepSc5e1hhe9GMvP876H7pA/h9GKiy3tx5kJJb77hL7okbqm
KfX1NnS6t+SuLW0zTPFjbXUJ0iP/A4aD94UpKsAprCUJnPPNheah1RJ+XYFe
NVWsYBfMev4m2I0qS0LKD6WBye7wt4N1M358KDpcg1ODDUw9r3ZPZkuy0g9e
AdZ1gn+9877qY4CK1yRjVRRiLcF9z2qqr/Fc61q4H8N3F/9r6GCJDROijOiJ
br1knIF425w6ii2zPFHLU7JwUNYM2HuxeSAkBbRynZVw89xhtCtLnm8ODXS3
UNPlllNCJReBh+dy3PfPEoVp1FJ5iZW67OALOcRrCT4WyANHqo4O6dS+HPHf
jb3KM7tgtk/jW/+cPxucuuruvRREJhffdgZfKMU6XC/8N2Zln0sXycwpyg5/
/Mjnd3UvSCBfO8Yhzx+NOWTnt+uOW1oEpB46XT06S6r/aKgwhbxXKRxQ4eCR
tJb0gpyMIpJfytYWf915mzxdrjcsXTwfC/mMlLWNlGFUX3ex8L4FLDys0IdR
kgm8ewJ5KECBFzzIyz6OQh3j3iYdJm7QhvwO9e4DvEyGVWI5QFTMkaqoQtH5
dizf7VMjLnsbYgUySHQZCuNilvm/F8/eYdByAEtR9pgLqdiOKy5+IUxjLxm3
Uewm26kY0XlO+Iswx8u5+/eEVOvo1wajwmsnzwgwg3OJCC8Y9LNQLG2jnTzo
PI7tRltr4Z/y8KbGa9QIHDnekNr0eh5wSamUYolsocgCrEGF35JF2vogrUPo
JEBb5g9RUPjiqUe4E49BuOxLtu+D6G+KJp/ggJ9l1Mf8te4cNlxRx8lxi88I
Dm6q5iuAmKbdv32mWiQIjD3r49Ye8TnL79lT8TsToUUIOqNEtinDi5vdLIsR
BN1dpyR2MmF8RfCJuquqO8rtwRU23HP+SVCRB3H/AqasRsambD1jvEN0eRIw
5PB0y2K0xCeCCbvfpwrFi9qM6Plsq4ZCR9YaGRZXKmF9Lb9a/dQfhlVeZIST
AuRct8oztEBwZ4f0MkP7BpaNeaIO4w8qQ44jZdNJ7nJBMRCsHpCwjWPT7DkJ
CST5/x5Yw4M/6Jq9MMVhHdH8y9ma0bxLqwh0qR7ir/QA45EfYBRvCzvyRqv9
O6aVscXZfiLdJ71F4uuho7wZ8GxLsISCVHG2GbMuYqXAXa/Ie9F7+4o2AvDd
jPVzTvLFPS7NoJAPNxh046MkDSDIu5rdZE12Q6+Eeh+mW3iJS5jO3znbf/cK
axwcNJ/8gq4PD7e2wJWLGPDPz6goyLTzNE5Y/xzZkQR430fDeTERBiM+yMmp
Gqeyoi9/kX4NY2zTXeBTUfhPF6UGMzckPQnvFOfptt3D2m+HspX5rhnSkITk
B/1twa+DDOH/2UrpMD/7w7huiKLusjaFmSbvNWiPRo/tXh9WCUS2znbFZeqD
hTmejQeQ+HX2crT4frkB4kGW8XrxEC2KgVM/W1iuptmtVvoVB5i7tLvylASn
hxDOcQdOw14wY5vIfYeKVUPbC+cDGI2trB2ztjrvCgijZXswkf9pUPxK1k20
gL5jRcxoVZwbTtGF+xH47SpGx1oufi+qDcmfrOc/cTuhMrdP6jTxuE5IGwuA
tnVUdfZQyTWBdlOqyq+n+4/VkxOAQEpJ4tNDXdNRmKNAojStPbRf+vTGMZn2
SercxN+4LZDeO3YYNpLnNdD562SmuWlH0m7Hlh8uDkCDyPnJ9CafiY4atTSY
JExlBgbteahz0i/AmGl1jcM2hLzQF8li0ZQ5mT21gYNV7U6OgeqEHlzGx0Py
VqMTZjRratxOdoQxCMTAbFuv5rnBYEujFqlfJHQhdNQ/irB/FQ3NybKpgZaS
q9sP4KBFu9nQKEp5uDWWVhDuRkfYNmPp9j2iunvN+WBT7ZNSU+gRL+siiaMx
MaVMYvoMbVDF8u9IjZxrk3m20NYXajkah8LvIRqtqmXYTChI6EuwVgPqDJN6
4dG0SYqgfoN3cRyPxaFhtPt47WjzCK8N9EY=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpeiALHmJEi+qFaMF6O40WOZUzQbRj8ELdFZ5Yjr6Ns1loisb9yXbww+0nJvVjzIYWf7NDHoZQb9TweCO33S3ziIfxi5Yy8d0NcRGJ68e4aHjWGJ25L6fQnduWaAX5rTVBxAuXuE99nCGsH1bI85ZeKZCbdT8QADeX6gI5zLhEnlYzYDY4C4bWYPcwbZbFU9VHIjRdGRBOuG+4kcxuUmEUGOTVJIePA7ve8cca3f0DiXqBsyJZiXrxOtHh5nnlKwoNdNsBduJzkshdKsMHJA6X1PP29kgLT/c6XKBqsKfAF296ANBRNnlZtB4VHEpSQuU7bh7+VagcdNfBBP14B9vidg4cOQwaTvxiZ6FpC1TufydmxwbG9n86gTb1XPpIsVvT4OnqG6fBcb339UZnPlRXS0gRsTWrAnM9QqMaBqhOMfw3H3I1nWwz4PDA7LTKL0cTWoVZUo4R4FZLgSD0j8hOfSg5UsO9tiI2Oe7jssjmsWmG0DaxaYOy01v26fOwXdwm4NIrongkS7EBY9AZFISzLTcuaKQuM9Vjnhl3FY5HSlDHCG7ECHYiiT+PSYt9fDHLob6tlzT0UstuWSmwtywXH0/nvyR5Ffu3OyCQz57Wa3cNPpJ4EV/LShEtm2bFJx4lQp6txU4ksVXrxilphezDIHXw/A76Z+71NrwdcJ8QWLlY/eGUfvCRAmTq9JhCroyad6GdKbcU8YxxlxjdFhNZh7AvIXaLj5NBkIYrglqXKcgVtmYGRKaBmpJq50Owo6oVdYP86mUSreBKPl330utJ4kl"
`endif