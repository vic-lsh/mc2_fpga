// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cAQW91GoYmzGEwAx3YDJOLKjZFsTG0PGaw/9uDskjOowbSVg6Q7fAi5D+EOf
g1yU8SfCbepDT6NmFkMz9NGHFfEwecpCgKI7MUBrB6dz5FNDLFd/j6dJf+LE
j9SJUIfgXhQdkozxv0QvTbXIFzfsDQMJFkUIhaL9FUk8QLXhW7kVlJMR/Dvq
99o0r6ZpkZdErdgR6+skNtKqXQ48IL8ToKo6kkXx+taB0eXtms3aAsTvNcNj
C44VWujl5l3Ua/6vkPqxRpAujBBzNNnIJ0JJpy8i6WybDA4JzTE5Fn774jE8
nOvf/cuq9Hq7jjK1VMkssViyhLiPNGtgH+FpWuw4eA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CO1/h7TFU8DK5O2lbN9FK2EcHAufDJV8WTkg0J0MFTAwuccPNjW0/RwyatkX
QHwHIC6ED3a6U/2JfqCkXw81XY0BRSy5YAwAO9Gb4XBQz6lVxNAjxexro2Dq
Cjt5tfwipvfpNEo88ihLDq8qpYH94Gvguo6FBDU2aLcjVUMWgh/OLKQy4+Ot
FRbPbGDXU8siZ3Rj7lST2hBCZQM8QpFbZl4I5H+NHlVFJz00Hjn55fsmb55n
1DMNiwOsooG2Yn8YAI75CI+xOPhrQdiMHsjx2ZYQ4VO/2WbkH+iFUl3xfrdw
f1MzdlKL5zEb1I1BFOOH7sj+/RQiNLJlSXY6xfJglQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KwaXV5LoCHTo8aPD06gdMO5gMP1tj3VIf40DfxZ6u1vrF0YWugVxL2tR7aOY
uI2aRYt+W4v8qNPlEaOn3SJhuWRxJ18aWoVKmNKhX0z2oj+ewO+uE0UifTVf
1MNIhxNFmbeYINkbfB4v+YNLDUv5q1ZofOn59we+MsvTuciVMLapz3FmDhUK
EkUAIsvRsZfShItVMPdr2YOayJsJquiOBdOotBjg0p+Jyn4pFQgA44ng1pRN
3MEWX5AcJe0RuLyjybTCNNc5UTL5V6JofwiK2orj0r/nkZpU3zADSSr5iaRW
iSJe5MCy8djLdOIllGEX3WyrMyYG9mDAyAtyYj9hAA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
L0IaabIex0I3as3VGq+H37beHor1j25lc9CgIUk2+5DYI6te8gYkTe82Vv/4
JBBQkvt44QAb67Ug/jsJhyR4HwiMCX/XmGGrsiGhViekSHERNKbo3rwDVXES
+1p18FZGJxSukcnfKCIKpGSwVSETmZjAogSFRjHz85OCfb5fEDeSsCZdRa08
+pFEUIU+Nlsu2s7Ch+RyHy96daAj8f8h8+hbCD6hBpY6boZQ2NdPOVwItoim
XN4zUYJBFCHkifVg3UgE4q+UxaSw84wWmDM7yuGCgewxqLLpzj5wfwVTh4AY
lp8A3JCSVm7FJT8a4SERqzdPJVIH36yOb502i4Pi9w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
W2VsSaW6pJ6MddQJZYkbpk3OlkXpqA8BtVb5QbLYHRUzRyZtFH5bYTZuyBuE
L9nCfIqWbQNo8eHcASvQzAgKjRr9G/MJQzsEo/ASG2+oQ7mJULM/bL9f1UtJ
yrRD+XKOIceAdVZZgXM03r0NSdwCV7cif0F87LedmQCKlJZbuYU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ERcpnAAAsj7xZlSOHcM1f87zg5582VTukX8aOfiDRtDefxtTw6sihY2MjRKQ
cSrkZmgBpXjBwCZblLlf+F6WVQgG60etewish+0VSTYXybivnuq2WrUnXYxW
kInkFUv2wT7XeGastRY62xqNyZ5LLO1u+VJGKhDn50cNXc4tV6GQH0x72gzb
zyLl7XvqYaWCIKMdATo54OTN1HHg/cUDqZts5jhV7nJ+b28IrswKfTZx+/MA
hXOV4T1WcNDdSoAVMmC74voLp6z+CJaJ7zZlmwPs3IFpDB341tAD5F1lKium
3eXGOLjf5McbNdSioFaO3VY/kgB1UUgga9V+rGG3iikyGeBYToUGJpA3xtwz
3jgYSyn2jsLsoJdnYuCsuln2IgDX/WxWgBmEmfRyX6gg36Z12QMgToXXB8Kz
Yf5cpBGa4B1DQHFrf0nR74STOvDcGE4giENMWKm1+6o/A4GnXygE5RswtWiY
RiWN6KM0goTyS/7XyPbSoRwxmdRDnflr


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
E3sd3zduyA79QTwkbWRTSXJamJWuxejx+dZz80hwKgAv0HnKoW3b3UcP3oxX
mht7zkhdrHAI+uVWBGZ4I8ezylT8m6ktThdJGt1vY9y4IxTYo3yC2TqoF94s
UfJz4SdnSdgOvwc4pSHw3dOXUoHVG8MULUb3Juw8a9Mye3Iy2Os=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qVw8uggLZ1OVwa5zOkT/PHmsgFXNZUvNLCziLaXi5O6Jf0HmYJdhP3y37cli
6x0d3zWpy/o3Go7qQR/nbI6H2PT3Ua5A23U7GJ64eRrb5g+/2mDeEv2T4S+t
ZCEZGjP5bj36WvKAZ5JIRNcHvKntShyGecvd5R3LSH8Q0GTN6fc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 81616)
`pragma protect data_block
/Fcj/VH9UALkeQuGiK6Cu0IDW/Z7vohtnL0YCeCyMtULr2cD3YgjvLkQ5vKh
XEsRQywuvY4XqHPcjjQb4g1gvuurpNVEZaPU8zkXMVGB/lvzzMUgJSWSkRR+
G2Kf0a3RqXRWirvnZpxWmIrWznJGJIrH7zxgdtRjszBow/qd93GcWNNEPYR9
dPIjjNU65nhjwgapW7qrcA+j+g3HX5ubrHwZdLB3TaG7KsQw+SG2AiG8nQCD
q98MLhvOa2kjtEemDcJIwy8hHDn++xoO+yIgb9rR7VyFLW4G6KVU6XrvSqSW
y9RTAUcAJ+eZ3l473dgCDdoY+d1VOVM5u1xahAv7neovnL1aPZEbBRwjV4CH
SfLPdQ00+bzSp0/gPG+UPtfeozfawWv3WxNgLquchdfhI+30PCHla6C+p9lk
z7MCw7XI41wHVnaAC5ReA8f4ybeMpHZMJfwShnQoulBMzc9WNDVJGHH/CXFn
4IrJ/2Cc1NwmiaYszvhd4t2ZELs4k3Kqdtuwrwx60n90e6bGCjUVGrjiJHqe
1UE8rgBJIx6li4yG0VWSaO3trF2Vp/a+hdNfFeWt4PTF/d9WdLs6oYFH61ZS
3Mz8Wl3mSdit5l35Q7RwHIZm60TaYpQ6BI3y6N8rSr0RK5ohagkQiFG2gC3Z
qoQadKksnKAC0ItMPT15ejNIOKVCACuQ2e/pYcdT8e6qWlWzxGO8uJ/bxXB9
Km0YXX/ECgKtYv2iY0H6E96I386hOxWf9jf9NEPxJJChVLKXC4tyMa0Lqb7U
SsIDT6P/B9BX59VxRJYZkX/cMjqjaIgaopPI2fdyZh9POmGbjZNTvqRL2siv
0bbEg55S/MPNeE1RqPwszKtr2VB5KdQcx8yz+Q7o7JI50VnQKsrbfyEhAcI1
pwT2teKrMAxk18evLzOw7iW4f3tV5J8ffNehD2ckhlkYP5TLR5vXMZ9h8tK4
dwjbSqJTNAsflN5tIJs+kRpfH8a88P3Ms5BJGKwSpg+3BYv7hnY7x+/7RKAo
TjzzxAvtEPFIiLxMe2LsCSMni1CpOjc9dBioHw13pfFVq2H0Y+Cvrq04UMjI
+WT+oZRpq6yDISqWx7MC6kryiogkxGKqFl7nAqpiisvm8JP4ZZgYa7HTE0+i
krtR2btMNeNCiXhpuZc5T5gBpyHmkWzaBYM6aQLcGltanrD+KUvqVlPHywwT
SyXrr5PBlb/c3GHBb08xGwGZsT46+pggBI7U1I3gvnxNYw89lQ3WScGCIou/
dkSuyb9lsKtvQbgJmKeTDcvxVlgep4cyk4YqHuuokfqIW9Mqq7APiE5QDIL7
rxKNMcbsLp3nPazX5eshiwhtVE/SjeT7ew+521EQXwkvsqZPaJ50pziDqxBK
v3FXEf4LLK7Pv1JehbvOPPKFJImbevBgGGurJVb/rpKaUlm/eskB1MflrHaX
DkZP7B7PrsH+GRjz8fjrG/Ocp/shvTh7Tp0qg8WXtp5luV93NyJ95VKmVx8Y
+zwPL/Ds0kDJDGkM+2BsCA49wjLHSfnlD4sos6wOhgjr4zyadRO0JxJsXW+L
ipzAb7CEFh5YfjdwzDMY1t4GKv32Q8Kdr+LXeExYeTHXpUUrc2yFr04mk2Jp
8Rsh70bnW3I+WM81PsH2cQ0vYi/LZkfsftCWq7KhDKAa0nxgpapbQoeYpIvl
Sz35vRRfGvv0Pae6ertSSZDCwp5oCoNhXmaJTGilqvM5d+gna9RpQ+jBBx7U
ZB8updFtb0k4XCwX1ZQG6MraKuG/aLBB3dpZ7kZE4nKGumTVVvE8zmN7sBao
EGT/oxoQcAsAoVkBygZySKTSiZPFrwA+VJWyRc5EoqPdr/oRpqKd5cDfk88C
AWLWHTAx00TOvz/ZPij4SrMng4tiHb4kswguPI9XDuedA9EVjhU6wA7osTGv
iZJn8CwqD5/YZwAn5V6lzXMhrUCRQIA7imQjP6b++HdTt7kaZRfh13jzUZiP
Ah1YnhZsJz67QsDKNvSKk13NkS5G1a4n8UebDyO0B+lfbM9GQDSwI9ZNnvwh
MU0Vqqjt7AMM1eKxw81rduyriNwzWZGhI77dj3qtfWDyui60rPeboINfnOc3
Xbb4i7FYATXfscS8wPHKsftKyqKqd6MpCWvx5yT5UNci8zB5H6juyxUIaxa8
e7nkG90OAzN1VbcV1cqZuS1H5/mcMuJ4j14l+TaoPqW5oJwYWd1URPANoPuH
OlLS7IxQmE3dz7ptHt2W4TfovHdYMhcZehVdY0GJwlLAItCVH7EMm5GQnXyT
aTLVLReY6vlMExGlduEWkURCc8lVvhU+X+K4dwPo1jzxK2UpBt3CZ8vIv+F0
E3qLB1n+2EV7+fNrlvmyyGhuHETi1j8u8WiSb2fZ/mYuLaE2o3hi/vrLKljU
aj+eLlFU+IgCpBuXjKaWua6I4+LOLuRIPvjT1U4u6Lwy+0BqbdEhlM/6T1Qm
nDbJngpQkBVTt8ubgW5pHx7vVBDDpYUoqemSMbZlUzBTnRIpTI4czHfiQGhi
g3Y1fu1FPANtx2sIbP2EjrlZy5oDaA2kMO+xuTqK/pNeQz+Z/ahEfdz4A9W7
HGrGhHyFN0vCpCYPFZLUXGP2/Z0cQu2f/lvAqM74sJbIZEvKmwDNnS8/7w9e
aBiQ7y8L433G0VmVTaRmCp+y2jfZ/qGK4GdjC2NyXqGuVK7bJwbKarnqVjaW
gisYHKEU/21in7jk2qOFDPtIAjjrcZaNXBL+7VEHRJASyYQPm35SLCNAkwkf
jzJBSbFHv7vwqvIPRGcd9uwOJgR+HNTCmBhs/bnzm+hchdfKQZGKmkkSktYx
EdTrL4LRnk8bjEs75w1TSrW+qaT/JawoysdARIJrFUiM2pYOFmm1C6mMAvaG
qBbhrqSrR5+jdBN+ECi9UIeEGgrbBgN3ykNS+0RccdEBxVsKuQtiZnD4ZJ5s
mP7MQHzQXVcSlrXlqO3qLFxCen7ONQYEChwQVsYUqgqEtEt4nhT9RbSn6gJX
nNU17dWwynANROZej18KlY0oDinsm4DU6qyIippqzcLuV/ePWiDvpiUQoCcc
ZndxlG02VXSx3gOYLGsexWv0pwjZMPTtNHe7VBdjalH8c5k87dVs1yVsfEMl
mxBeBzHizZ82nIaPUv+nZLCT/cGJUxuzzhPGXPS/jV9H6N5Yc35PSJokJAQn
ILvojknpl4nyzWPNk79duCLDP4mZooS/ucPUlzJXJH+mMzYJAOwkDTIF/Uvx
gUBbrxG0sBjbq47Z2gx/fmbnEbtAiMgiOkXV6CYLQ4xWQ2k7PoKt7Cqr33AL
kz81bjja7P2PW1r5IZUjJqChkp/NgAG1qy3/ctV0F0rH5OijU9pHOyyC3Skv
juHIFqUaZKJ0w7fGHjnG+BAIt4pVpvSIsjjr2W9YiV3hDMGWlEFJc9fCzvGb
fv+yC3c5UOoKYBIjyGlOMHlsFCKY6pA+T8xGVrkr18YkIyHXmeRbhCR8BR3v
+lktYbyE5Cn7t2EFamlfwHDciyzoRsaDjwlx8Wf74u9NATpq5IYI9ks/znRw
AT1AkmftOtqvc+31uzfkcrjSrZtphUeWvu+fsK4sF8xtJWDV/2/L4Hgl9JH1
MC6RmkZ8RCAYcUn4GAd1TGhqbhX8Sn4M3LMv8y5RHKW6dZkH7Wja909gOxSv
XC32lOD69S79E1BQxEjGR4kk9Ifxw2gX3Wu3KY6zLO8LDkS+sTytLRsmNpwZ
LNrRAaESTYMrA2Mhi/vwo4S6cJGiPlujuyP7LYd/gqHrc4PZIGuglu5ncpgQ
Mr56LORNtmYw8y3nCeiSV4gSn3MUSN5cmdZFqAUI2sA0fcyaor75q8Neim/e
9eoFAP0Dc3ZRTtGMrAb/rXxPJXX4gB7EwiogQjWRG8KScr8Pa6x41xDo5xbl
i/6B9HmlQAlpKmb4IY0xjHY2vPzpWBm0Fi5uxeNK6eVCigpywJHzIIIfjwnV
EHOeHx8/axeMBkuf7MK77o7AS0bal1YxtATis0JdaZzuAMVGFxUlnBEuqCvX
7KvPzGxNY4i7Okgy7D7jjFTzgb7GyMHQqXz017po2hOcL+s18tPeQXrJo2iN
czAZ+xAW05K0w8W5bk4Z2goLrLHp30zpNmmuzEGCWTQBT0QzyTkLNTNcajl1
j2HH2fAygF09AsZh4RkavoEYV2XTIsISJ/4XdSuz5nRq9iVpfpWgLaQEhQna
Go005XyovhRh0RqJcXDda9bIa4aOGj7kAVsnWwknMi/17HsnzR6RvU2C1saV
4HqbUQKw0O8bff34qOlZjZqA0KyASdB+ALdIkfkWWruFfDXIFHq+zWjwFGIu
C2cDy0bcw5rPjinNYiZRZ1W7GXslLRHAeMBuqwzDyyV1C0P9ZwxpZUaRhX+V
17AbfFPr9/BTiKiK21DMSUhQyICbwD2YbFa9qVSJS71843SjH74Zx78t0ieX
4otHmdYWoWaAzC7s9eF+5Z5EfxfoenU10T9DTqJa7zgitx9BfrP5LRx95hr+
FdeuN5RX8oL51533oKKtpyuL2ng4JQu0cYyMO+D9aVoYfRBHUJ3dO+IIE9/8
NPz/4Ogm76Ozk62You+TASpY8/RRHC1bhbosasb4YZJbAjlNWW5XkxBN7U+r
IZPJumiUoAHwFa2m/3Zfr/wBdF74jkhjXR3rnthHy4dywi/7O0MfS5NzsEmV
ASRFfMOVu69EZnkyhyOKRB6buWcl/BTBkPiMdoYiu1Dm0elTGEr3kNPhVZnQ
Mwoo2obtE9dhkU5xu5s/p0mQXDGMI0E+KA0anhS8M5Ltjxw2W8/MMqll+5KR
c91gTGrarokopwZY2EPgw1SuhY7Y/lFakggLm+Ljd0e1Ki8lYpfeLLN+qZ//
oCn2ILxSo6E0IP0K2LOoX3a1OBEMFX5mnx+wZ7GPsAgM/EXlt255H8Mr8ttc
EwPd/3k7OJy4/gRVMnIicsuOLrLY9LkQ6uoxFM2F72zs1GGbaVXczdPqAhoj
XaSk2mlaL01PcU8gOsa+iFXLXdOKIRd1eR/0Q5/M25KMHIpoLdn5RUwF3cW9
P3KELzkgHshC1rPfbWkA2aZDEkN8QFlrSX44HwGccgU6FuP20h4j26liTShp
OHF9q55qzqTvEq1UODyQ6xbU99aYdR8dGOK+f5UicIqivCl5Ah6mNSUxeN4W
E5t0lRlDmm4UMZb8RNgeTagUE++osvfxIcAIkZVn0F3eq43o4mahrRLtmdI7
8KxyePQBLzPcWWTzjA5xXJjVkDGDMVffuOHz/XUpGB+l65rHZxq2na48KYKd
ThR+gqoiIOIIWeERH8Ics+urPlP9nUevBWevs/zrfIiCmhSXvgtm+8ytRfhE
v6sAF+F/A8hExQ8sPK8jEmY7V0b94oWCDKM73zFVwinDD+WXXU4fziPs9LTS
8yuds0nlDCi+wyQ2+uqhvVlKYCJDF27YibY1vuqsvrv848RVsDBL49wwFldX
01AwwtMoaTm4j4uaDkFGcF1/6Zo/rjh1BVH4EZJ0ua++lZRgHsZEDAikYYp3
wzxcjpH9WhZu6F5+USwWekQIPuRZNc5WQBuzJoeyCWL/5BAx+94rv+FZESZH
aBx1qpqRSOxgJmQAqoRisiqU4aqmMXOZ1KUukJkvxMfVbDnOnPUT88YEg8Nl
M2IX7WiJM6j3n24gnCJfpdJXPDBOSPCXPWz6121lzzMIMyiyTFX5F5yQCyN7
VYp2KixJrBG8PuGArfH/YLdnDgWOrFZB/GxOQ3W5+o7bYS057ZfZhImHYe7G
pwjZ6soyJbXlGOxuGt2nD/Z+zixYq8oJg+Ns75HkWlu6ftRZlVnNH0lUY6gG
p6jrXYVCEOaotIw4mN3XX/OL7t13eMylAbjMpZqgCTAaeX4qdXGs61bD6aCM
l26QHa4wVME3ruCLrWU03+PWXptTzUJaoZkpoIStn39q+lFFYmAGCnFqxP96
zqh1LOFQ5AhCRvAiwo1bDi6kKWWGkL6ov1vymFD1qslNLAlS5jmkPWlJWoN2
90b5Tv380RmIFmMvI8SSqqDmk76jd/UqfneEjQ1t0ApmAlNvt/cFEZr1wHYj
R8AiTX7ovc34WKobS++SHd87SUKPpH3dq9QP/uDDkMH3nHg+CJxgsBBwE8cf
jf+kGs9qDO+j15vrDVJEMu/phuh61F3am8AOIYG5r7c36RIc2L8OEEiN3x8Z
p9ai4AwwvLTECyGc44SlcHquoKswCupGrUy3oC7Ekn8zcLIon6/QT8YikQvA
WBJWM6PysGZDGAu4nR7li/NB7bd3YZ7AMh7Xm5DWkQsp9qQDhIZ5HGMygTpC
HvP5b/ylF4KbcI8twDk73iUoQCPqORoRP6jLny3YbgKsZtwkz4ngOCzUJyCk
uaStej71+JOBP+mTz5pIBOZgx+6S5gke6xReICXmMC8JuPA28csulqtAR64F
w+sCS2bD74ghN32m1gMQU5FxSwULr3jGMSUZjS9nrd5vh04pNP+xtpXlzsLJ
B1FWTUrWIcd8NR4x++RDD4C8odlTC4Wqgni+5adiCMyq/SfysfIRLuDJvGEB
s+p5s70NifQ85Yd5EeT7oVnJuFU53gG1duVUe3UynT2Zp7xAfWy4snpVVewP
ABE/Xe5m57ucT5QuO6OpPE8K4JxRB6AZW+gkO/8Cq6xX2z25VoUhQ3A2ZnMc
72+YE87NjgCXhUzasUW+Z2c/GXFgtOnvWHRZBMNjrc4mlJugKB5tjQexubCG
yFDG77JfoNUy77F6hxGS7G/mkpbsUUWjXGifWCp6cjo11D75wT2jZ+m5IcMt
oJc4xlz/lxQnIxJIazlFLGmSjKdG7ZmuCcVpDc6ZDE+T+pgW1tF7q4APtmFo
PsYzUAZdCb6qMOt9bTF5BFAqM19wGqJu5laC98OQ94qHieGWx3l5GJmw52/B
6zn0gqMdDk+C91ox+lIcTxWttaXXmK5aUzYEUAC3eppAi6uV/3dvwcRFe+LP
0rtNvfM/sVKPT+RxbJP2w0rYT7Eqoh5CXYVJfDI+ve+4UBjnd7QOIVS4yUiy
KHnQLRpNXSnASMXMXrGcw96J30lLxL4meV8BgFZxghE7cEQxjiEY3HUrJoLa
lcPfJcBm9Ukkgc0sjAeg4HICylSO+nxYXP5muDIZxnFHApkqR/BnTmLm3H99
SaKP8sxNM0ZEpI7CfLfgn7aVPf8nQWBLzIZqz6FtlDq4Xm7/jI5gEZ/a8Llc
96EVoagW23ANpgzTAchs57eyWwjvIUJAh+WM191daazfamA6wpddFuqIRc+K
upvtoqfAlAfRchuhgPyWjI0l83YSleG4wYrpVgoVDe2BljIsxblZt6OCC/Ok
eI6PmqSQAY6ifSXCfQetDtZC3xElFmQiD4COXszJ8aKSagEOEgLqX0pByjAA
OTgmnbt9WAjvi1oBSqJC+JV/bfoYvJ2DZz/E8BfB1J9HtKwE+S+z0HUC9TKs
0LGoxrtx+kLxswuJ4QONtIVHL4GNoXbletKnvpRSx7A3zfT6ArIe27HcTS8E
7G0CibZ00CI9AIYFwEknbpqgdPnDOpkxjdwwbcFPf/37UbYD8J3sAuNhahAO
zkPlQtzWdhz91f3jovwAOYEfT0rIBv9NIqFgtgyY5eez2xdptAgDxHIwKSt8
T2PoaKlhwUm7ggsltjOl3T3tVCjNLL1HwtE0bZBLi/YFLNN5Mp2upsVZhTTi
MPyWzpAWrUQNChcQgAPFreLrU+hJsouSiZxbWmBW82g4W+/Joc0RT2VuIAgg
KnLMCuDqPN2ExpO3BdQ8sun5ELmCg6MQv7FbY6hs1K/W6jq0q2mb1mAO78P+
cWYwOHpY/Pr05J50eBZNgBzhlplGEvvcDlAxUhPSULUL21q+5o6BD5CLaGpR
mzaKpXkVh2E3lociXH3YIrVhgF2MSFW6fnvR/2ENgSANf/2SKhBF+tCTCrbS
AO4anCuhsOxET6whvpDXUjLGHScaNdZj6clAgYwuHxT8eek0uW7PkkFBwnVV
o/BX5SMOKxGPuqFVS8QXh2Rogow0Zix45kxT8ZXtCZrd35lgHKHosDAdJfKe
7ea5AeK8+XcHwQ7CyHhboCGHzCMt4q0Ol80KN2zfIxOdqwo/IhIUNjV1fgXk
/pq0b1dW/r25yR/K/Zt/dLDHCyzCtqTdsg395AuKJaHtb5bKpZn4UCKBSqCD
WqmsOAXTh792vMs2xxvP0YNJ6RDiL2nd808bJJNh0al7YZiCzrMf40gFFBkF
LnRML0RoPYALpIf4dds+ABj8h0fHDvPGzRs2lowpWbaMY/453GyxljGdTwVp
FsLL1xa2vyaRDz2qZODEEEWXWkOh6ODdFz3ctE3s2ywmbZyOl4Ih1TirH/G/
KkT0X/d6ji1z8QIoXARijb/CQkkk8UKNZVtY21Sy0ZCTHsJG7WNx6KdAftAq
9FxFQR5EjhZmX82OnfN24JsiT62WMy70QJcfhHj8W8IUPLkj5+m+DkyM4/Vo
scP+yOwMPDme9Imi+0WrT92+5q35b3CjLVbjHLgm8sgvKi6Zz648Gl/GZltX
O/Y5DDu9tXCmYzNmDmsA9jvU/lD0+E+lri1ZAuHPzjKEbZ0hu3HAB7JOtdN5
rXDE+ZzJp+36opkZm9f5WJdRmDX3x6b4hD+g2BvYU4SLjVxpNOZVVIokf5Tn
LLePf/aXE4irGXxpXNQX6Vq2bvFrf/5xvLWr7q6QlFmxSNPAQICrZqDhrsbL
tI2ciTU3xaehWJQtqezE7VqS1EMTa3dozUSDuagDFM6BNWB8DEfaej+nJ1j+
6TauEBmNA6pZFUnDXZGlCP2O0kF9HQvRFn5DBv9Xnzr4MZ/d8snNqJdQBtOd
DTwm4qThrTcW17nDL0yv4DpKLAzGpkHQ3VyLVS+ou7S0emarY28mqaBH66CI
ZdWKunfX++kwsTzxg+xT/IXOL/eN5mckhtjYZtj2AOxWkqdLiFm+mjTid3M0
uFH7MKdie05AukVMfWJMtamLZnlj7ypEx/49MHR6LIwjluJ9iyEv4Y3rlcS4
oDdAmdM9V5aBq+uH8qaU2dZjWx9moMJ64gD7mlAK+k59f7V2AiEzoWR/IUCH
B/d09f+f0yxdhN/oOBavgKj8SWbIdxRbA/uCJEFRmW/B2agObuBKleXhOFOQ
eVKk0QQ6LC77AsCjzSQNyX9aQDc6jAvpPNGf3ewm5r2fE0CTxYdNW0bFEhyE
1gz86VQndnDdVNDO+TvEdv6nhxDlAr5hEvGLN5wAcJTfp5opnnH7+F2lBxyU
8gwfDIm9kj+aOnIAgwsvvHfYFy6Y1b2a6t+V0l1G1vwyTg6Ji+zRL1NKvZ8e
TRMxpmCrooKKhqNPK+0lwVZffLe2kN5200Mn3t2XNN0hvlsOkZgICAMHERum
UxqHu43Y2m4EwkjlByV7pqM/ddOCOMIHNSKarMc40ClpcUO7KjykOTAXEC0H
wZqRIq/FEwZEt4lbeUc4o7cd3WQu4KIG+KfmUo7BoeYkgdoHceBHZHmXrMlm
v05H/jaiJwcL/vGVIGx5daHzKQw4M5uwOVQB9MBC5kwfVrjI44qgyJQaGSIF
x2hDqvX9Z3BnnAzj2VLBtUb0xylMGQs0NxRY/xO6LdX1GUeYgZspl1mpcGe2
vKn86V8tsiM/jtcBPaFyn2z1MemDvI/+wlWY+1BWlPRqxXzwzMoi+y5as59T
dqvXVdrcFy6SZYssOm86ZfLno+r9CZAZA/Re8/GLc++C+4s6j+6JAK4NES7g
805Z87EeeLJaJBzNE+OrIUqGVRPgEHW6s6MvlUD97nYM8swCwRfHwGLooXBn
ThE4tDuUNII8u6qpa319eQjuAID92QkAr7oWoX6EDFImq+M0WDtMwlKn49il
JFidKhXO6cFjo7J+Ds2bcRc6XzEewoDrt+e/3n22WnlogHkz3P3aCishkYPc
02n2x5nLBrqNhk47k2n0CVZMPJ40kR78j6/DRhkmAzsfTdqBXEH32zDe1eRh
8qEz0rrutyyEFgx5iUJuhVXcYPp7X3Ryi4OTVyn+h3uPgKFM50sJEf+GIkC5
WY1bfdH6v7kX10QBrpf2Wl48LZok3mI8SFW+oMbyCWiadAAo5IxG2TniYHHp
U4sa6sVcIIUqtKI1DhgFVcXV3/vIX+1fsWHiFYPWUkUGYVEM2Q5okT/BVg4K
9N5+qVOYEjXtKKSe1GgoQZBSboJwjF9rvT+eBtjHvzCEDIubz9LV+UTe185z
lZXK3zx/e4ydXZeCQiygT+rDnR7nP64IlGS6R7L+rUN+5AaeVERRrLgWoGTn
r+5ee1o10TVCASl3+KphOucAYFN0dZVefjOYpJu/H7MyL6eTj7+J8vTlxwz6
w2XhFuLFPsHHYjG8qlqmd+q7rVXebJyb3fDAherGDpzoHcFRTKJvU8dgILyj
2rgayVqrb4EMFFJHQ4Dtf0dy/vqGMz8W/TcBM+IZWiQ5nXjVORxi+klxPF0d
5v+knRx95vo/gehKY7bnAH6glpwZlkX3G9zO97fXqm7q9zZA9NXWyI//saog
+nD0tK3ydyS2xbblEfl1wigZrP7w5zB0fO8IjNSNsZFDiufBLAmZZ/nSP2wY
KhkPgxY3i8FtvoUoliFFhgwA4ua83YU/++E4hPfD5hZVIlOFKx0hq873NJUx
Ba+olTHdyMaPFrvdIPMoBCumLbDUZGjOdkYbkBQf6s+FbtFJbGRhqLuJIsp7
c58zZsl6pr6kFgCK/MfCNK2Mp/ctlMfqdOBVTwQQPApeDWirw0I8d/ouvW/q
i5URyVJALBkyuNIlIbCbages6FNJWhBFDHv5+LHy6EjKP4JIVZve/mu3EEdj
6Cr1XmWKBqKgUuuj1yIazA58G2vT0BJcqtS88GI3icrP1LlqSA85/LWFRiQz
L1lrIq12CLTSWZYO5tbwzzTHfDkkqaiNHpsDnB3ap2Zg4Dvgk7MXzv/gMXJE
btLWRlZw0hpi/H+ZvTRYAf4QW7PMIaef6rJcEmcG+GqnyJS44d7Y4cWD7Uvy
34BWrZEKwcURkNXxsVpCDzs4aYlaTnFJOhCH5GqxZ5eCcfb6v276ZhCHj8Q9
ZlBn0K6kNDuZQ9PfUP0t/nVjHMbIOldIuS9zndNaX7+gn++o4uSsyS7UiKDY
aMv3P5S3A4BWIdM+P+II6kCMvIQNEcO7sMdITqosv07EgltRybGoLRwWdMVM
uSJAUMbbpjRT+rec1plp7zrM0MT3OCiuHzrXt9ygscohcO0FKXA5KJi39Uuc
UsX8W1UU/p3pfL4W7RBM9bjcYl4INlkuLvvCIszG0BVL+V8OWaFR7K7fCZfo
nat6V/JRQLqSx7N4+n+/xeW2lmXdZRrmw7zAJ3C5a3xiKQ2MhoSYUV7w840f
QQOdRX9L19LdNzAyqKm+hT+o1KClniwdngk3eZfRWRrJFA1BV+cMdWngxVwe
YmdlEkcZlO85tbD7tyyXgFJGM0AJjEWkEgL8C92g8dtk76LZc4Bmg9Lj7iwl
072OtFqyG9xXnWWcVzj6nnNklISk9x/LjCvH+d4FiL5JF1O8GfNBe7G3NaQ+
W8V0EwEFRr0tUm+zxUwumLJsC3zAd532n8nOa/5zFxwOkYtfnZjRmOrClHg2
F1QjN1Mt6R4YB4Kqs2stQBZWKO2wTy0bMOic44Psl6kpFnnrY1S6si9zq00u
vN085rPg9ZGUFjZ+aaq0NnZe2ib1hZfj/NjfYyvi2QL9pIUaBCyzVH+IuEst
vTGo9fMvPWVHHtk4KXtRLbmZWwg93j19HGajprkZ0Jjw4vmksBIVrMKCn13R
QXNfG2Y9qQfwhNhWypSGijoffyoYxxrNJLlv/+R+bOoPk2OHpqoGrEfJuvky
IuUr7A8wcr9CZ/zEPoAEa/rsfgLtl9nEjzxtiwvoVe8+ZIHr5ZSw/bv2JQ4y
DsZyNjlGRAhcEEQYBj0JheDIvpM3uay5l+uZOj3CiS13BZVIFfQk8BRbg2KL
NIcw58QNSHB9Sran4AwelwM0eCAu4L2qffQuy5pb5abztNDAxyIfXhj/NMct
gXkVf9XQw1EBRD8/aeWpOrIHkEW904GdEh6I/rGCjU0vEU75sUbq1z/hOwbE
J8Q6gbrmarrums2PrRE281mFFlnnjBBN0dE/LJvuKAXdHDFg5OoLmWMAJJc3
NnTgcn2x6FKHgmQQJQvi+wsh+GruvX+AahxGW8dmZKb5kgmHb7YsZQKl9pKN
1x2O5OE/u/eJTd5Y0HBQXYlBnLcdIHV1Bm7clQ9aQk8bnp/hZcyBDgKlyfJj
p7BxH1/FueizTp00H2/Vl29OcCibbt8n7yEVSHogtOv5hN8cEz+/5VReW/YW
AatllY/dIPgwXye34UGGNc+9YNhmAnZcTBsMWpOE+CJmGYaKnq9KEe61sq6y
O3nmxNH2PwAyUehdTK79YwcEq8suL8ThHAR9S3yxr9il5PxjY5qnHUJ3NT0E
JGuVy4JpJNPySGiMKkyLMkx0m4z4qB/lBpQeapx5YQCj8robSTiCbzHu2i9z
j13Uaj2K8dmbSk2g9KjzZbtUFUT6uQ9nOoqVyQ692MLSACpMXu7X/41Q0nOT
3I+kAezfnI72xowI/rRUWC4RHEjrBoxxS7qP+PAJR3OOcxkuCxmehlux+pGo
RLkdscab7IoTqy7f8uxni9AkCE0J4ZdysRkFCyQTeUzn3+NWwRQ1uWep/Zlx
5LSgYEEiZ7GDsT2J9ujDTeoyXrMNWz6lxAGTsRJlKOQWmPQCnzl88nghrA1b
wdO5gl1yH7ZSkzljPHbxodQMnP4lEZEX/QBqJIgEr1y3RUiXn8DZGzhVr4LQ
ZnaJOIiR1tZ9VjN1TZK/KacjkDL2M/2c96da8WClBxvS7hSST6Qxns1KHkiu
HITnn11Z5q1AkEaQ7VI4YM2xnnJ/M3LOX6T94SNpGz7i5kH0B4Ogm2i1L+0A
jdGmWe2NuwZUohIRAoK87Gd/lKFIARZnh4Vvx+xEzABf7U0GnT+YKg7oPjLN
wEf0nJ9UXzGGpG/UnrMMZsCrEc41kakXH5vqlbp7OZ9ZNQnqG4YeGm/Zm+Wt
rR5vrmtDgyvqEmbQGHafDjQWkn/yOdY1r+PX9cdX9IbhR71vIYFGKZEcnfiV
jI7NLVPVtGtQIEMYpE2mOqeehPmwiNdFakMuonVTZSZeZYGhRDPf2FfAgzf4
JQ7RrUoDrSOYSjgw6FxXtrJGYE3G9yKAOSUKZ3ESsad+Vwuenz7TcHSw84hU
KU5aw+B+z/lYhvvBUfTXMCAK52gXoFHmIOVSAxGUmKVyAiVpw1GlvuB/oK7/
PCuoxjURQLvFJsk2vKWTkeNMo3JtKcLLwdFe4Kz/e32i7LaMPtyFDXzJGqj1
PdQdgB/Vc7XuTY5nbwboBlSfa5cpqZ/iw6XiU+yiaeLYbgEqcKbuvQutyRBA
je5nQZQZD8cv+6Wy9ECDx93EpQXgKnBEzfAtwJrU9zH5QHt4aPPp7FpyUj8o
A8X5IQaZaxAXpgMB3PSseQB4IeQyeSIQygvvaXKPBj2ndZWB8BLTI/CVCudE
fFKbBboFFAghTT48PTV0sJP4Ky2HP1EVqcGIsim9fHN4XIag5146bZXnoqvV
x7DGp4XPeeEFqKNjJ2iKw5Bf5yPxou23UbA7tw/jXXDS20Jjl/fs3NbPLw8o
vMSaOtD+YW3g31JxA/Hmk8wRNxbeGKCSZTvznIMeKOvC1U3dXSIS9CJycJ5k
SXRAiZoDwx/9ZHH8rjSqrW7e+hKN8w5eplaSw92au5jKxFFl560xY6KMfypf
u8rUEDVx82/QTVch8ZXuV14F3TrY1e8I8XqNuoiBfMIAvyqfm/H3Gh3bMfQc
lLuyJCoccX7lDcYxnzF48V8jiZkFkyxo8TeOpnN+yJ1/TzktggVl2tRVS1XC
YD0SEtetvdUvRrit6YglYRHYGHl5UjOjNt64Cj+CAhTkDLhJrXfpKTW9YDRk
fcUEBKc+De9sOPl6TtXyDKZgbGtPcS1Vu76l2guCIoaHQuaDQXo8U0wg+2d5
lxcZfU+aMyhHnmI9/Rv/Yr+sunCMhdgMCtHFlCgdD0RZU5uN8xrmi1D0MRTa
zJC8mN/KYECENdotzTy1481440dJ8QRQdsqmXGBmnE4HlrD/nbE+UYWruBlq
+dSHUFApiTQEh8nDxItUGAhPospEIY0Twi+G35IOyFfn1IH7yfANjFe6Z64K
hWhbJu0jHiJ7KXbL+6XiV3Eab7vDbv4ReUy+kepwlgWP6Ebk0JBi88dxgZX6
vXhtEaZhJG+OUkOFsnLTjj374/WBibD0kwDa4feXJP9k5TulWv8Lf/vSnRXi
mkX4mvxNZZwJGU8jZUXGBydmhcqLFHXG/qMzPe8POFyIVbjJUCO7ZS2KPBOe
h+L9h3GJXIEr56nURHVIhL18mwfMxYyHP8/sc8qAQ9pn3voTrunLPUhG0+51
wYFyYfaCrZlC49yETGaf1CFjpCXDhVrtpgcdRsAv814A83raqM1yRv1CkZ+3
M0WA1W/7TPMUevTCRBKSdsBOKa6He8NERncU+mWTF5dzJH9sI1c3jTeDts/i
3spPIe+IPPbKEgD7dxW/d/HKjSdkXk9cQIvAkBqfJwL+98nvU/v5z9onnBBd
uzxbr0+OtIFITiJ8Mn+AQ+iPnwla67ocNADTVG7s6dJLnNtmk3fGHsNL+ZXo
bIZ9R8mrzOqEGyLmqSGveBb5MHfJkYLAxjMTRVwGzFwzcsk7OBCZGJ7GlKv6
0FpSxJBnvLVr0sp9HH6X84A7UAG8OVHho6kWxQ/5vHFRc6J7GhimubJ67GSR
FdVj8y18eG0AwHsonumd61iTzOD4y7tMVHWoJLssP+Zmkwo7HlLuPkb2A/x0
HHVIP8O5W3vQoJgQfUZojuMt9QeLwa0dFkDMUlJgSX7G0/FpVmqGv5q08yWR
58SFVuwL0AelIaZhhAJE7OaxvEAxgtpuHrplwkYbW2Dvs/u7yjlx2jiDp2NH
0MAQR3WNCwNWNYZhCKNEwiyAlCByOgurfqFwvmV8XRELmKhvI2lTWeTDGVV+
DfOBx6EPWW6CAHPv6QV91ZmDr9lgnFtTJKA+NMYXUUWaQQysTozlsh+isBrM
lkAwacwXFua+BMAZVsBhkOAS6bFvXZ702tmoG8S/ePoD35IMxUwHMpCJq5KF
U/GIeYrdMqZwAK9WQoz8qDiEb55ssGyMHlPsenmjhZtRNnxU/68kNomrhhro
upe9Nwu5q8ENYOv73yPP5zw0Q5+QVYQrGEm1jwkkWUTBYMmHFtSHLAlM4PZp
Xjw3E+X79j+maOIyKZmN1nZlvjs88d54tvz+SEXUsRd35nOJSsnvk6cYZ3zy
T0I0YUcW5gTWjbB18eEj/YW7tvTew+VnFwA6lm/IW5N6VHPZALcToMGjxcLS
HwQiBbLXf16diUzq4lHnITZ72N6K/WIG44NFNS6gSrgorrMWThxnpH9QPLE8
0y6/HtyIOyiina3VbtuwkVC3AeqGMI5LEMNVYE2JrnkBiK0wt8xi2n+YtkLa
/F6HVKtxOWiwsXm8gv/VhLrJewuYRj0TiVYbusHaoD9ZtYWtfqxRT2d/UM8W
+icw1HoOvhDlSXCK99lAi4NAkcwnLK3FsjKcUcWxZc8OK2JA9LwhaUrGh7wH
W2atEglBP9ajowIGpL4Algo5QXX+UAG7kIB3s2tMsIhifRiHgzwbUvpe9Bjl
GYzOtmxo9+cUHW0RSuRYhnmTNjwnNWDZjCOE9WnMl7WZtvc+2ZvHp+IzVXTx
YtNwotDUKFMUf7gA3Vt8eVWm9OtXPcwzDyfEF2cr7SXqfTs//G5xvb0pYhZM
gK2Xho3ErsEaVpFIcMAeNv7Ae0sOwtriTyYg5Kwq6TtjI3lcDxW35Yu4LT6J
G6Y1i3/V6v7bd6pk1QlK2IET4JcnKwgnYLUMDFRdC8Z9C6jKlQay0ib/TrfO
KdzB0Z9NwCo30+2XbAXoo/Gkupipw3GKx6ScAYdbmxkC69TodG7tRpeIZQ3i
KDKMgc6m9rJHwxRO20cxGBiEKxmV0fM9toNy0wvGJVc+ePJVGDt+FZG9qovm
v6qRWUjS6xj/+PaIKDa4lrFbBSIuwRPoL5cTobSwwmGH0baK0DTsQfl71FMK
KuwF7qNN7mYYP2YH9r63JF2HDscAFAL4hhj/Ve8P24QleuMitgNHuWmGKjzC
AWpnPrVMb8Thu6vcbwBo4vioc8vTsPlyuT9wPckmPqYAjl8jyrgRf3LS6Vau
kvBQqhTtIHxjHb530VP6Ic2MmTCAkqrmVofe7qeXvmRclRiT6KpoWz4VI6j2
TXV2F7wHray2ZvxPz660A+YKQdQJFzh2vEoIrXdZIZ8blAUDVZgUYp1H8Paa
6fzSLF8asIJgPZ6UP83S//E2QovnOwhOAhQf7Vc63wKYVZ0htYU/j9zgBPNy
4N+bH1MHUNoXdZiWrDEtTWKwCsdmVi7YdEatB7lu90uR0lrmy4oR91f1qODj
AmN//559tW/GTshInKz6ABRRJVjzanKiYLeY11TCOsoSf6WIVpR3qFn3U6/J
sst0AvITLVy8XjeKBm89jOVbIlGTii8fb+8wvWIHG7ofGB00bGfPEW+691gQ
08Kopx1d6QUxVZohHTB26odTFrXC+zacGIkkdMnTAVLKdL7Z2TkB8y5LajII
nT1U7Y8V3+zdkeDRWg07+N0CknbluNfQB2KHWvoYxdHZWGLdIpzVwOLTQsC6
oLMNfRFH3VL85h73oaQB1ySIyhU7oQ0fJKG7rxx/4jBjG2lKb5ick97Eb2i/
qzT/EWR3EsV+OB74qsnd2ajHPSpR6hxRgWxrKnlxf7MkPxiKtGMig9H1tj4F
oXdz62aY6chbYsKsrwZznnn5ve/LcRcww1XFsViBODxGY9X9utQK2cHv5Rh/
yeofXw1cIzXsaPD3a8bRBYD91sadgkheRhNC8NFhfeyLkEZLaR4/21VbXZD+
XZHXpGcMYgCUatwB/2N5eU4XY++CBndeR2DxTdgqi6f3DMpRLgbnLotytpNh
+GlntMadlazXLSilfo7bdaJRye1fC59eCULFZOf+LgNCU4FwfFCs7vUzCFKl
tNJ6dsY1G3QeT/SAVp/pmRNo+V2WiA+7ZXjvThfGBu30D8GOEmVRE9DQZPVp
wSYFbRItWsI+TjrCh9b+lcYkdJEa4llGJKjxPDwst9pzDELH1Q65i3fyrPz5
cyL19X4d1UxL+Xk4Q0lCUvV7c0CfPsuS2zrlSA1QaJ4Y7b0hZS3yo75dM8vc
84WkAQYAKRXRsL9igqQBvX1PflyZKdx87o5q7c+DAwBkTeD8htNw2XcBO0+3
fmdxua4ikavaHjaoVqC+Jp4fjhqTGjY05PAsl8ipaakKg6aQBmcRkOozJVUl
aPP6UMO1puHhOeSTuZx+v8/iwqHTwVCHDz77CFwLMecW9iNYs6LklrksB54w
Mnf94fiHIgN9vkpLU7x4J7kUvQHbftmP1F+tDO6w+lBuAKWK52g2s2tv80ne
/m9E4jlM/w9rkb4X6N2cUa12UsEn0ZQnqr/xdot2G1+XWZEb8netVpNmQrwv
9SJ9r3/OmCAJE/FnypduR2tuFOOqhkfqXAMqQLD0YlR8ysW/hL7CElGiQAkt
tRXIgDCmr7DMPzrv+CbwCcYIggG0BRa3/gQb2dXT3LbQ1T2j6b1O7purj+Sp
ULOxmlnZ/nbGoWwpNuiNRt2hm6FvhONdRQis/ejG2mJ0UYiSwTUgbRK4Nhuy
CP7EU+fzromT5YVzZRjNvIIX5tEd6vFEq1nFnFaxkH6ZpXGVl3UEp2/FfzbN
1aF7PgzTtQdVVOD6Pk0ho23Ot7SycI0+YAc7QRKqb5CtbXa6J+FXNf4manv1
tyuAFOHNOZbcw+q2Zy/pOhF+oEJYVjTFrUDoRlil4GU/rpoyTQRvjZ9yJhjh
4cv14Ui95l9ZvmBVnjiG5TdrUyog66HHapONDtlxh8cny5RJI3R8SCqPnjgj
xuNLtagJ0qB1hn0i7Xt+NHuDoLbVWStkkfXAwMW3qw9Tvv7Rr7vGkUf/FK/6
5+7RA38fJ4hbk0Bba/z9gdindHAWFSvh6aWO0trO7qGqQP7w5d//MXenEb1w
QtaxWFN2PI3O7FchoCilbyZtjMqH06Ars8K9ocaiZ+qEDziaXZgpbnBthmL8
bcG5jkTwUJe9Sywod0SGUcAnEBkFLpUBNw1A/qDAQAFRcUHHG4ZGiKl53YfD
RmTMkoxkDuF/sW6qKjcp/tNxP8Vc1aTlWZlcS+nuGKcymj0Lyc+ZOszH3PJt
Kb7Ej6bfIY4OkyjM48DDgclzx/Dg62iMch7qe2LP94HYya74rrJBmmM63F2X
SF4evAJpIG8TS0iqvZs3aoNWHFbn19auGmVK5m/JeFipv5E6ozaKHT50ymNs
tUUYmsY8fKHyaY/wgDOyXQkk8L+ZNcpCNLIqd2O4BHnGsuIve40braVisYqq
KEAwBuOrLV5GbdIwjONLAJHbsn7iFb4/0eiEQbCeEkg/s/NxtkBfqC/3IjOB
auzqcVFJn/cbOc88Pk7wbpASecVVLEHksmPD5AJrEghT0m0EHTDqB6ufUl/7
+NjVdFev6jVTm1mFmQn5QDe+Hot0p2rmGQuPYo/cxNE2S3u7g3DUzbAmo3n1
bhL2wGal9htGFupn36ofjkf05SGLVTWp9N3POcpfdeAIqtD99kewNO97Vfau
A+XL/mrROvHrdIDz5TUESH3kJ+MdUcDKBaSA2a5gua4gKaexe+boaWFul/tv
WuGCZiOH7dqIhXCofipPGQkANH0HMgUUwORJMgw53Pq8OT7sErDHHq+cm5rf
oVg+0EKtNynikKJARWLCVG4wU7wiFOu4k/ihtVvVpgD0idb3EG5zBqnL4srY
KX0DmPaUkS+qsc8LY9hDRcPmy5Rr6JqpjguAwhJyRQT6OmoDNHkWy2t39ZOZ
9U0Qg6qdNnsLvrzULZgimXxqEIDhI/+vhAEzgHBzEVl2bWLeJPoPgpK8p5Kn
7HbclACTcEHIjoeerV7kP0/O/UVTsQBNhvjvPs7LGL8wPMXaISxasx0/3Wwj
cNsqFV5WebMYz+rfezAC4CpTcxMctYvdGjDz/8qMqaDa/j0XnMoIxlrlBPoG
QamYKVH8RBvKWVjJKGhcttbCYvJIs08GycPjSresDaXP7bOgSgyzsFwpy2JX
kV+Ce4zcRMMda3wWlzAqcjYdnvG9ADCKm4d8tRIf/khwAHsAk0iWuATbW9jU
MBeLYvGjCjobAjWx/mLy64QPgbszln8mxQtkQzfsgs7CH6ni5Gah9KmAu+yA
gmRtBgPJmlzv8GURe2M4/mPR82ueCLoyp6d0Z/UfbBUjiEhBWNL+mYZTltTC
8kIbV+NbbXA7p59mL/fcNyYot2ottSIaFW6RtA5ufcnvQkAnEQvvQOu8QTSi
PkVjAS53RQIz1CMEbro4QoXmq9BLEFpTuMfsZLJS8GmTtBErj5AqS5SaJxgv
VwF1mficTzVs2VeGauBbK3N7jNTfATibN6wm4byFIwLmqeNfTSSdNzDgBImU
+vLmlI0lGsWM1t40/E+3jF/MrCmZEuiFplrg7ShxI/qOidS9cFF3ONzeDqV4
d3AxF5tmJoFxwMDIVMrmftKjTuhisKa76SzvfmH7lQj18aAA7gDUR/pDf8DG
mvCgCDvXqzHT7wk+to2/ulcS6t249RwcSZtKvUbM7c4VNYRWaqgsnZ9uCPTA
SYKpzQ2wGAeBpEAn4beW9/D0IfgqHBFN71r+Qc2JQyjh5a7zRPCLjAS/oIej
7sdjody66GmGT5wOGY7T621Dc644hKwRjBfBrzPe6iogJaSo3/ii8fQwpF7Q
WHVbdutE9PVlHvOxdqGegh5kd4CHKJ8mPwICO7DxK6GljzA0P+HoncyuchCv
DmxCrLmWRFMv8hFFf9rxopBABWzqSt7oMYltHcI+DSBpy+QlbMOUC2m0DbHj
aWZiUrz3aNbTmc01qpnZhVMhkHsNbAglY0yAlbpzBmtHvJsI6rmiLtW2ho5L
WWNnq+uR/rbOVe9rY7tx82nq3mjQ2l1wnKWKU1Rz0paotsvjJMwqUbdcrnZv
x14mnkQhFes7OJSZ3t037sJHvWXcaW2eh2OIYd2Ctz+dbVNXPC77lUhJCQAQ
5AvzsiocSdEnB4L6exMxV7KYPLikAxCz5QDNdiJZnZ9oEkJdFaOKHaGszjGs
ojZiSkgySfKIC8IBWMhR47nJYXdES1bpA4mMUG/XXVgTYS5sIDRuoLZTQxUO
zXm+qDgzqifCUoiDA2dSl6sLR0IiEJiLRPJ8wOxZ+kFlIsV+EPVu6M/nYLl1
dTPYNLOlrBKAFLPIQRknrgP8MbhzFxCPZXcb3zGqxJkaBXNS+TZulmPSNC59
Sf/62k+cKS+our9Me3Ujf2Yfzc7QvWfnrw4yWZqvVLvY//eIsMVS6AqGSu7P
sutiKnljqmkZf8H0da6s1WXbV5p5QfKfD3J3f/U8HPJ4QWah/vzRhR+nXqLQ
iE1WF/T1R7HJgM2E5oeHtOrnnEYQaJX9YDFGrw6/avYTJX0QuJBVmEfsDiZv
9ouRNHd6/cjvvEO4hpOMf3Yu1RQS7B8h8zCKUENEy684pgiXz45GkyaAIR4p
Xio12qAWJWfvI+wRc81BkJC9sQe2L5w96rGxtkATp0uo35udaAfUvhwGWb5N
volU/ug+iGTKQil1jzc6sALO2xVnyubV80BuR3dbMN0MvZM7geFY2y27g/GW
/H5NmBDwtjoft2VLHRbCRbmHTiuwDV/itaL3wMNX3rCAWSc4R8SY/bL7PbLd
85joDcttenkwLIsuTQw8VeeKtSEnh/TzOaAlcZuDLjQhWR6LmLGXBsggST4H
WQJiTI40a62OWaz0VgiC7Zpdqi4SBrlaFyX82qawfwNFvXSLSZ/eZ5+XthXK
xXig9LHn4Fji+33VAadYGbnGaOyJ8I1ScWA52AupDM2gG/018r0jVALcu/vN
7ahh1wcL16spz9UFjdPyd6WU4nsbd1WOJ8BMTfMuQng/EodJBQ++pox5kizA
U6+23ZP1vfuQefFLmT9Va0Xsoh42mBAKk7yhvNkKSpUGIVWoDstgzQU1n8TP
zKFA0GBgy7Cq+orQyNxoc6x/HrTl58Rtj+wuTx4lX+DEeKSkb/X6/QoTcE6X
Cr0XHn4pBEXoJlTrm2aNX4Caox0oqJNmiJcY+Np80JxGHXJr0/Tc6d1gMdDN
X+CEVsmbXnbrAxvEREarBLLxBEU2WjzZ0+C76zW2Xyt5ScDXfpJJCc2/RQDi
nmGpYNcJ037DZppYKAkODQ8FLWWBGoY6RM8n+CDlAMmAnlTr2816IboEcJk+
KVR7oBxFX5CsHEbvODYwbUEwoZEmNRfx1Yh6DswDbUlPlNemEIqNJ8KrfEaT
S2O97DBXCBy0FuL5JMMCRgwpRPvBms8KrIhxSohdRZxo/RuyiiW/Dm0EfQik
JpoqFSdXiI5I0PtdH9MhZm5hq1c27iofzTOQJFmJrs0mkGBnidg+9qdCFKXa
SW3BmUhSpOSPRPMAuf/GnaXRJvvCeN3GjrdMrSVR+4XCZQ0+pgpg19q3csgN
/Cbd/Kv4bXd15EQFgXn//QV1zyCqQmYlN+9025T3DfOZGlcAu+Rpj5ginPep
XXLi2hHUSmzFnEPOUAV6x04/RoWnOFGTMjJDfe5Lza4o2dcz0f7vzMFaxzSK
GB5Uy6cc9Yt32ZMLBKyPxqRSXxbqRo8wdzYHFUD7J6SteMTNTLdWoyAcVMvY
w1h4fib8c8A/UYNhw+x0mFgRRZ/VASdti+268SPZ2LnD8shUW1MZZBzhQBrv
LCfGIVJfD4VggewNCqM/ASgY3+MpCFwKXivLVayQSrX0HVt12+2bzQqvhhR4
xwNJy/Fqfbyr+UYJKH30gevZcEoSIuiBnrcvDF/A+TfMBaCrJ1OTu8XS9RpZ
+sNaEZb8sIMKNCijUUhgtQx0Y5MUV5ok5aXYODvVM7aUpR4O0JrEC4oSZtNg
mG3vdNpj/JgLkx6amuM1eRLU9/ZsgNvIasM65y1tVJpvq4iT1pIGT8zO3UYF
1bWnpJIvfl9ySRRF3WrYsAhx7Tya3ttEgTEZASrBz5i2Gv1AcC5R60NpUwDB
M/Sli9uuCKucFuWeMk6NA7YBP2tvwMkqEHImNc0FP8cbDI5zGB2ksSwH2/Fk
QDgPGH4lJmJX4w+T/4VokD4yTS5bb/0IzscJuSmm963gTZb/1eFEYPUSQ/Ty
15sgO7tuPfoDj4746qzjMahSqPtfURMWWFkEK6GjdYAf7cDEIxIuXp5KQDCB
pacjm4QIghCbKb4OI0onup8nlLPiSbZvCxmSFIXv7zfsi/OMAKhJrMUM6vXm
snEv+4ev7FLkJ/eAhcsXcb+bF3q9TZ3Pet7Q4T2ZIlqTvbfih2ZRs/4WVDE1
yw6tqiwmTh1VqVp+xuwcgchM+HdupAm8Kg9mkuGxEbB87s42guIaS/qwGqUV
G68/f65VeMbPFaowgIj6YN50W1y5VdRrWZ0O9XNiIMWqXh382d9N9jv5fGs4
D6foY7JTsfuiaYf9WXT1XV5MU4N1UvYd9lFFzb4V0QNEU+ULewEIlEbtEB0c
gFg8ZIkLVih4sPdA0wtOR8EZ754LXG2gMSDgvIyHX1lSxoSCHDOoRVHutg2t
TqTSzkGdTFPvi2+jzdXRjYYE8ZpmxAnDRWhhKO2n+oPZPQetQJ18PvT3oy8G
SA1gZyhcOmUVOimxLZt7R6z2fXCda3OURJWw4hSnckTtYRjICt1zUjJ/nRj5
elz+hoJn++R3GxSV7S9CbSDi569oofwwhF0c5zh739+9+iv8tjzvLQIwEIUb
lOZwzmbprW72sJI3pa8GD5jPgLw43naoDceK5j5UVbqIV8kGoYyv9Du0U1IA
koe1/twqpPbm+D2Bf9gadavGDU5pCZy7qt/uNdRx5LuKYxejehPdi25V3QtC
IFw+WyGNVBwEJe4BJhblv8k7cAo5LY4vakCNMBssm7X7aeAPWqXbmNza8io3
QCGLPESJ8X9egFtfv+MBWVYXCunqvLJwSWjw33asKos/YzQrUce8vyzEuTFA
URGipB9feQJU7n19zzncgjmZrSiXsolEVxmivGQ2wOXmmNh/e00FGC1gJiVS
iaB34dRdrYA5l5XPpxDuQ+FRvqj07HQ2cwC0FXQKfgX8tglRgGNwDWFm8CL0
FqY/Yr7mIhDZly/nG24IYHrwqGF5bBJ03N0Mnc5ooCPwIfFFvFKMq1Ul15W4
cTGQ+XTQpj5c4wRNxOHc1AYmYCK/dAnh7K6s5Pu/t0F4HJkm3lTttlG5urPi
TQul1x4u+hSXka33i+2FmlSmSfxvIxebYoTqldYFnpHSpZ0jCCeUvy6Cion1
9HbnJzreqinvNAZlHVLvqtDN0LhdNu54qDtNQ5trVnFz9u1nBnV8xwt3SvYO
J8mMOY9XLNgjw8uk+8jmxo/NCgTRBpoq1xC4yn/g+t3rdXFRgLt3c9CSFx7J
qVJj8vDxfLRVGhS4PgsNKBUnOmPmthOSKfmwkABF/rE0/6tnD8vq5ls89k1B
SOubzoMo3aeFOqVSrVWGPKXB0Tg+FjoR1oxitct3R5u0NKOALZbO0gF2zhzN
oM5kxB65M2YOycmohsIh+nOPK49L/fRr+kev5+WDtX5lxWekq9YRPPuRh+zi
Rmozt9woKcBf5jr1TtTktZcuFa5OHxi19tUhKfubCODkLWchoznqXE1UNvuY
jceTBcybB0kLkYzOSGwHCzF5HNJNJ+qFIsWWfderD08QzXZjkfuQ1xvHCpxS
7OFajjS83WssNEu9xPCQpgFYs21Z7l4XE8KefsBmt05QR0CpDb0lMLpSU/e0
G/dOfuUj7IawF0O2qcZeG+yaIlVxGmO2zoz47BvPpHkhjb/TbQqTe91A9cV7
O8gPJu0b7+WLU0BntoEHdo8nnG8cZ6r2N/gMOVys33+A/1Lz2423SziI49Wq
rjus0xbkkdJsPdn4ZUtbIuW0dsVO0FSM8qj4Fj9s2Ag5OmIS99tQgVJr/Hy2
G5k+FEsVhyiFLn4kkCwR4ekumlaPWZzpki3EAfWZ6vrBr50r6V+uESior5OH
DEZUOB1/k+uRA1vX+V6yV35VrbikGbiHakD6jw3f5V7ddHmvwiGsfDIf0AhX
syvtblxaUzGWkB2JfViIPPQCtgsSFk0fsXszp8lfe8iv4VN7xxFSqmRKo/Qn
1B+TL6+KO1FGzLQeHQCgV7gOgByhImJmXJ907Sa1eXoJ5twQEaKnFiHKRnN9
xlfodeJXUkFpjH3+ilFGi60UbLhohmb2Q+xnDk6Y5NgdMYEQQ7IJ1h1qcQwI
mLWSMyX9bdnNFZ4i7iJ3b73Q8Pu0Zko1AZ8oPGkjwmksKWlkM17vcf2iXtda
scgQ9wVP+6PXjPpdqid+IqjCk7y1yJay7hIpXz1Z4A0fioEPI70f9HG5zDmq
tfcj7LmcIza6r6YdluvreapL6L2hP/Z6Zz7DvSkMS3PSj0wV/PSK6yTNLtKj
XBc7Ava8mY6KOIvSOV1qrAB+napIn1tWiIsUVHbnu7TPylcxnUlexPzf15nA
LprFi3juco7noEQUhqxuuphgQ638WsR220CoVe1MU+pqRbw0lqVX9S9mR/4y
F2mU8Kgq5rCRW7xJMwybB1UT/COZ5icfmBdTxpYoRLRkR6cJSVk42AdlhDtW
XtGhbSIhlNze/WxeTLmLXsfaCuTqSeyFEwK/0lU+mE+iqzqz0cHkAWP0Gig/
D+M4GkHtFEc1KDMzwtWTrtHblX7V/WkFf1kN7TFZcDdEE4Gmd4J/pH7mh83e
qOmE+ihOXkyH4wmfKxyXnARmb9EyfHjYkXsxBUpp8Bk4G5hCCQ7gZUVyuDtX
PBMsiux+xNyW74kUpX5kqTaPRl9uvF1+2aB4N2RgQ5jCLINN6yAAONTRnkpf
PVFlSt3N39DnyjXQzwySY/ZLqTZOBkCMsSsFlHRHhe7n6M2eVRjwjkRDQH0F
FfOgOow9F8ef3H17e6mg3p7BtxSApdxqlj9eAw+vbu0ThEVRHCNpk8i6rQya
k362pJJhyF5Rf/1xxwg0ZsYwYiiIRALI+ZHN6hi5EsulQ/M5wqgI9R+u4T7G
rBT1IjGkNbKNkQoNd8M1zZYjq7MRhXVQzPmTD5Lj4fFJdRB9kbrXUPeyP347
4hVPvFE3LUsAYHygqGdQP7XzOq9wQ7vVrouCqUnr6X6qQDFOs+AZNmSHwlfi
DjtMDArB25jSkhrtQ/Cwd4Qk4q5juwBc1CNXHKn0f7dCD7+h2/TymBJR5E4a
QEFwdARbxtlHMRnDWMAUdnpgZAI2SRZCxoeHk/8AyeWYDD/HoZnOst+eGQ4C
5NH1jvxZrmuvYPOziI84k+d1vkWv0VWkKMN+mPlqloU3FWbVGfP/K4952l5h
JQhQQIvVSV6kKcyokoLfCSmkIkQuXqpMHjZWBVdGCIj8CcJTBv7fAFi/0S7U
Vtn+nqqZIKm65Yp2tTUDN5ij+tQqcBsRbiwCSp6EXz/9+ffxuSr1yDLMN7L0
513EZqzqM3zHawurbLdOEwX03mhnHIZGy+ywA6ys3zPC7StXQ4+iKEvDaGyA
qyJkv2Mv51RKlSSjgofyJN5TYK3Gufl5ErZc0MUamf+vnW91b8/9ip5ykprn
SEuWxKC2jnRcQvK5hNah8kM5EqYbILhY+gbq5aSS74LrMDVnhHPK10nYUO7T
KifXppgFZkUhmyeMT+kWvHwDuXTvx2+DBec/8mrVzliaFgtqLLKTolO21Yn1
XiGWhuQYCQIZyQ5K73A/0NjXyTTlU7KPrFQ9bKxP9hE6yYsgJgPmAAWyRkBW
Gf0C0N1eJ4jdkfbqzcudAr+okYZQk0wiy3YRaxLuPJ3ILGrBqvBRdmHRWqWf
vK2fwuEEKhfDmdeb5pw56N2oAEbA7R5YfA1E/rjeQ8dhy8qBLUQZCaPE/+Wf
4PBd+NtzFDm7VSBFWhMwfUziSXuhy9tdiT7v47blBxhCn0JvH+h+AcdwK2qw
MhUXOAjBE9SSXvsgistj9f19ev6IMW8zh74ottL71ltWjBxwMiWeRxYHeeQT
MxA1/sERWVXpRdpSbZ2jgh+RTHKRchox3eeto3Nh1teDVrgtXsJ3Ez4NLaK+
6w0lLArCYJ0Y32YSlzlBpOj3a9wH88FIDKyohsEhsxiVrJHJHAOWnqHV5Kxf
qoslwgIjuNzpiXej6akURvYsyEwT2Lj23k0B5WsWZFo6W80VfNBJqXEtLBrP
MRnkH1IRbRFTpXJ6en8oktNpSMdGUEFUzP0FmAu9bq6t4mruxya2iUFmAsRu
wVsaOB0VQj9sK4VGff6HMA1zu/xI1/rdTma0SHbYJw9u+fbQuVHp83EtIkIZ
Od9RraGkoc1yVNeJ5ZHQ0l0wmGXkfowBkseh1bPcijFL1g3czb/LYhxIzdWs
6qGs/VWbFePcFOYXV+xmrQLkL77lfpmvgAsxNfGm+67m1TLo5QBH+D3sLfu1
bvkyX1tGXujzObXKGO7qxL6pLX2AXud1aptPWXkG1SuuZKKr4rqmXBwhl26H
edCoz6wlXxB1AC1bJWFnamx+028fCWuhMBhkH1iHqbktaE8hMn8598bKm9uj
fSKMBLJtFVY+y8EX8HxnymAu4KU1xX50Qd1n6MFbY2r/CfbdCFnEXylVjvbA
+B6PfJulX/4ynCQV+mT6otCodqhdAI7jFUapi02sWzsuw4sJgiPjgd0q5Ap5
YMvCmNlKLV+o8hUfJpgZtFLBmawlLpntGycYDSaAsBmemp9TWHB6/vnHigEE
GTGLjYQ3Fa4abgSk1Zg7bmbrdEfEb4NQcBSYuoYfbqbPC+/VckANvVEsqY0Q
I2CTsHT67W4ruDjNBZcNOICDroYzZm7e7g/EjotMI/y8qaYOmXjLzgPRjH8y
YRzrP7pFM3apHkFaiWVyvutl4qgt2ntk5OaVVXCR//EeCudzRdxYqfGcr0Xw
Md7jMoDZJj28XvhxSu7sW9BdqkZXmNIg2VYcsZ8aDsNsu3zq8berRt839Nma
sAjgelRtcceUZdhJc03krhshPlOiRBRCSfKey5HaTz/M0rRV/M6Agq5BAqSF
zWCO2JgqCfmkmNvgC7SuQJZdHJPeJ4SauaIY2Mqn+uQW6LKsMNele9MWQWOE
PeFXB+7SlGScHKAQQ+lPPRV/WOE6fzrLZ8psk7yx/VyoiaGssRXOpaGW4vGd
SS9SH+5GY0dHH1tW71KKkKn5XZWG7tH4OZM5ZfslJX8l/9otxx0OLV87iT2j
CAvwoZvOlKnG4LbwPR4M7BcYkhxB/1Vjac50TH8Ge1NyyHlRiT72Bj41dVoJ
X74EBdoXh49zDtXftt87LpJC1fXiT9moFo6Kvl6PpOMVkSUz3EvP9KYqdhBJ
yqy9m9cQxusre2VXzOR+h4GesbLoxkRGgwwLHFBl44pUfvdZ19Y4yuBKEtyD
4aKuH7cgP6PpYImSTHq0UYcmNPYPdlLYjpx9qN3ayY5YJz0xwS4bXwuq0Z6U
HCPlwJn1bd/mVrht8p7etJlYZkqOuGnMSnmooIinT2Xuo33wQU4QkjiYlFF3
2Oi3Y21WXFE9s/Ttom13N/Y+qNSiHwSdW/z4p2HDjs3b2Y+D8xAvATkvF2Mw
kJFNOEEMBYJSJKbW76h8JbnlzQffO/YmfdX/pHBsi8mmJl7/29TuaUD6oSrX
JnuvTkxiAD9/JlYqRVTp/E7peGLXetAaIDC1V2AyKdgZZL6rJ6KniFvwDxbt
A5s4cBGFrIIFB4OsrELFvoQ/TkQd5vIcyYeSNkXuV2sFCO9GqN3yeXN+LZ4+
tPEm5TEwXYMlAEBJamtEWr8rcb1gTHltwnVNuFiLQhZpTOBJjsrkx6pC5tpy
GkllAjnWGixFmKZzhE6vqY1Tj3i9gLDeLjlV5KvJJFq/19m6HXz8DGwhFmvW
tYzK4FJSQaYa+ZD8+z0ASdGs1CwiOjngYOU3A43Dmpb6ibYNJPbY7zA1KUXm
7xwu8YW7yAbaLBFCqtg+7MOao9GVLMaPGNIUhuhEM45Ox4w1RZFsQ09I6IGV
/2XI1HPap1FTCe+lYufE92RrRhsVsbXpoGVaWQ8lIj/jC9Bhtgz/FypZsynx
eo6zdMwiq8ttIF8uMYyfN3huJgcOzkbYTyXEFrTx7UBsnZtfRzLUurfhb+Q/
6bCUmlzj3MsKefc7GZyeRjFMZBalJV+25qCkzaJkbJueGOtPkEpA6+Ub1SJE
Hv/siVAND2zi84f3MWO6WxTpVAn/vi7VcgVbtWifZ851Y18g7oe1ytvwCDGw
r4MOybklZXU4wb1eVIgVH6JTmaXKTypoeihZhOUN+xWrUcoXC9r++IyLH0cI
z5CM3iS/rhXDLD0ywoZuwgzDtRbeVp0r87I65Kr8OxQ7Ubfi3e0SuGXPbCCp
mVzxbw83ukoDtwo+dG1WO1xNBwm1deNgL4YiGPmiMHJ+1a6c+PLU8Wnkmf3L
a2XsBQKaWiWR6V6I5hGa/UkEKXk0rAUeaEqfAh6f1mJJO/oo+i9gW0vjxZc3
hdS/gCOkf6SQWyB4eizK4vBPlIT5QWv4XYlAOudV4Sc9ATI62VsW91de5uHB
JF6No1s4RhtH0j0gJdfT8TUsclYZyR/PW6k7y2BL8xQuCyjxZM5Pn3lXmdOQ
JpOjTYjBSwoy5WHhrPUht2yZ6e3EN+HMM99AEecW6kArnR47AzJ9QCn7AVmB
p22ZLRQU6WPzKkMSLdLJ74qZ5GT/4v1EKa4PrjKXNN6KwgjYEeA0St85i0oj
C9p2AToXLwZ+9p+jtEf2KRNKOJm2KmJ1CWPyFlBBFmxEtdit8I1PQEhIIeAq
nWEWeiAl33ZTXYNMfekA8gZIOLZK2Q/609cfrORzBAgLJUoe2NFlUORrxKYc
lphTkWVrGskRxBOrwTyALuCQbzOsh2bEejwxYxyPhZRCjxlc3QVhZgUumzej
5/bwZrHbSOnm2hHIwCfh7vxprV2iSJOw4O5GSE7pO5LsE+RnPf5HwZijbE3u
Gda+Rg016MMi7wShxVW1NgwaFxaYYHJ8WpYUnQfHIOX6uro8jugyEgefmqzV
LcJCn+fvL+P+8chduS01bZcozGZALjMk1hI0+wya5mazpeTI2nAci8j2N85b
NP0xUXdf/Ly+G+OM1JKU4Fu2X7jqHqmlt+WLb5r8IcI0TqXIbc2ARSHE2+RR
CoASVDnUTksrjPNrkI2JTTMqLPpDtBM7HlojDFSMpSqppjkvaCl8Fnr3OMRH
OG/5uU45d88CuFx9rY/z+TqekGcuf0jBlil863jXpaXmLwwBXpYInA+r9A3r
OPj8wZfUeXfzLnJlOxR1bnxmXBYpfQJcjo7MywExAMUwQJxSeKhOPQbzxqO9
HAudI7O150VclM17OTPjPFRJ0EngedP7461LOyzmJ/MfbXy56cOGjwbBqA+f
2fvKFDcBpOCuKEjeyC0D4SB92pXOPi/SaDcZ9egGI/J/EMR/0m/Bf6rlq0Ff
Y7KG1AAS1/Q3XzxqPI7oE13uhVbXzOcWtBk15BaaABYYOhzWy3ojFu74aOLn
0EbW/nu1VIWc72Eua4zPvRd84kdBo+x0tWc3fsPkCS03lqMlyXqi9wD12OPI
/FJKIvXT4KmjP2nkALyPgsXSm0dWtKyaQ1ODn1y2jv//zpAvPAR6Ld41O+Zt
Iob3KS4YChzKE48iqqoBa8IC90xQLakNzn1a6OMY0t8lhNkfrpu6ZtXEUaR9
b3MbPDwK4Lh6chr0wW5CsUIXgjY2A7XF1ongzepBQX5s+hWLkDSq5arkcIwf
XpV29y4xK1YBtebX1GvYdo1w7TfLjg7EkJSbWkugWroZpN5cE2npQiwCBS+d
yPGAxaSQx6X0E1ToRSfJ0uQcvlXqKRp0j/JaRg4xuNETvPRUOjzRCF7yAn6I
fMIF62LSJIMO0vkwSxwgZzA3EM0RX3lmi/BIxn40BRqbwBOWO227uK+f8Yo7
x+vwXhjAg8FT/iODiose4MNJv7iPvBR+BAzg0GqDJ9BNN4CobAumu4rO1E4L
js/z3aFdmCvN+sjhbNuL0o8Sca2ODEPBZImI6ru/l1IEZTjDFuFnU8N4n1se
O8JpX3yZbj/wAjtm5Cc2OCjAIGXYd6hCjdKj9kHHhKWLSYoQ8GDkpyMTVNiW
VQogYN8V0QMSFE0tYI9p68+JcnbMO/0gNRodujq3zfuTv4Dplw9IoAGYevH4
GR5nKXbgDXggaVF5AdoKt9IWfeUtwPV5XORuWBiNvFgkUdjs/YbQ69HWcSqQ
VZ5QP/6sLmicXQ8UI6Tj1WJhgd2KcAeaz6pe4WVNvMSdWvwSC+owGHELJu3k
UNFFWQeRWcIXiUoLf+FCou6ntVT0Xpa+n2gyBwRbHMUEjL3j9b9rCo+Tc9lm
bXSHd95w0bKLwPIzUAoDcRf9P6xLMdP2a1qja0peiB/z4wDjsCYaUjTeQzua
xQeGkES9QuXlch6nvE/2pIq8QkRKIxPVtpxWEdd6RVzNq+MDPV6j4p54Brr9
YT92hKMn9KBU/Fl3/+fxbL8oGJPTgQpQry1BQDyk0yZlcSIi+qrQzKYUsi4t
6KvnWi7Qb4A+KzL0Pd9BO0s8vuM4joNVfiyF3z9ka+5xuVHn/M9ErFsh+oQ4
yKEeiwoir4QBm6wNAIsXei03w+gZemzUG3E5E0p9ZIa410pqWmDoDRKhmP80
UP0lelngw4e7/GiT+imKw7VW4kepUbsohTPwCDecWbiWCUJg7/+bFg65dQy3
zeGDyoAaJeINi+gdYLH1xlzRfEtCaIps/5VoRiYQvuLDzIH87InGzJ09CxuN
WP2lSqfgIaleF48C2aREnn1C4xNyrjH7aH1EkDpGJ4yhT0qkPDHiFN5WGQvO
iT9G4N24RikpkXSBCOiDaQ0CqugfBfywsQXyw0RqTAJAMR9qiLrNIhuMZ12C
cVnBro9sVXW2uAsJX50oXF1iKP686YyOyofLKU2yrGgQpQUnHPD2B5o+My3Q
awEbAfL/IQ++lQms6brs6CYU3++OjytCbpVFXZcA+BMobt+cneAwWYGQpFjE
OijGtExTTAWTVEqPVH3roXAtKk06652DCNG6V8qBSq8HirmOecy6WomrbaYt
kj/Dcgp5W0buw1ZWXzL2IIhG1oysGHfV+Fif3aKhZzQSJmeW3mktWF1ciOFV
347TQvFWfMOwRk2l2WLYmSL4SX/kvBXigcLW1k2PFqMij2fexao7gU3F8ad2
x7NdPhMP/+KrBtuopCLiCQjxmzrIQDYXrw8DYJpk/xneNDokyfxf+OHQIZnJ
ObHcEwkhXzEd8Gf6ZR3jULdsvOcWHPUPINHOO+Y7O1dwNiC+Gcv7nQiiApon
W2WDLfglox/zAja0SbbqWKp13mNHaLxTMplsmeMLrtp4WWrQAMH3KM8C42PM
rNGSgb9cHnuKUVNSlJMnspCzx5Hx313elrNRzDght428KafvpYntvaBkeVF3
9Vt/zBJlKhAt+HuFvqSiDoAbrjKeLaj8i1SP/eq63Dkh3XOlPt1Ippzx5Y4f
Q7ZtjQZHgakVO1BI6pggReFipPRM34/dnrjW4ViyuNOH3bXiY52/gg8ni7/J
YV3VI8nn4k5fwB6WLVl+WW/lXnvddRlIprjSY91pxGzyJF3MSf9i8hiUDGp3
dabHOdXAXUYyub+2/uckCdNVhtxrTeYiqxM4b2tawtagFgvsDasy87MzGYA3
bmgFTPnUfG9mtV00X2LNUeAnqOhNTkLZJ3o1qWvYLB4V1nG9Kj3Q7OJswKLN
66eJfTUIW/JtsXImApukiACZgdApK/6uTYyuLiqRaQYVd3KSgK1LPC9va/cd
iSC5CwOMIypO2nLG0d4ZWCqhfuLzkodki3o1Sp3Tmo/i79XH22j6lBmI01uG
lFTJVXKaIZ5Fkrm2Bv/MhscWsxjQu8DR7vo2SYTM+rM7Yw/heb3v+OHMkBAM
R0qzTK+iz+zGE5LoF2U7SNg6JoQ41A2jeYgEU85coPXkr0tFIyMLv9C2oGoN
dq0Lqy2MDknQcr3uaQV0dGLDgw2K6e9x7ewaiRkkSKyXAkSm2qtpnA6ZhJpW
vSj8WL5zS20LprKfSoPYLRTCxL+gFMjtpw4VcAx+0KhXKCeCQV93bvjG0TVx
lyaC06pTZOLc3XZiDwnxQW20YiQIdQps5frnpW8NR1c2ShVM/NSWXVb/P+oQ
clZc/7fRef2/+WXqyxf7jZ2aHT1KHVZqNdE4hC6c/dtZJlCMqCWbtoMvEj0v
WKxcqCIZ/0+kGmSUZ/G+x35pHNeAZ7VOgESheshCuq6LaYeRmVkW6YIY06WU
GuiwOmXyCdGp7vRwUvn6qrHTS2vPx6vkeZH8zn5mAvsTd41+pDJV+Jf6H2mf
RLNg9bYSCcStmf/iCGi3blAD0eHZQ7eSsBbtx/nHrkDMPl//QA6RXC0Mh0HO
sXGlEbdXEBlKYzbFcXRkF/Xl5lO/kf3rySFD3FB8vBau5LvnK/9IQ7UmH7UU
zWBi82vzbIXF0KYHpg11pupbeIWHRLc1IE9YvehyJX6pOzBpBt9Vt7Kd8R1E
f3psY/JhFynD7vNRfyzkmOVy99Ub6g87qq6YPZAo69k0+HTf04W0hpM5gMa0
wbuQyBFh8cCGr1MvEv7d7EPoe/4Me2TMPmdGXUso5d2MpPg+JUGq3CsExlKE
XBaABOIUsYlu0EY9epMr2iciINJCjC5RWU4KSdV7ytXjz89uL0cd6SSZfgGg
4A0zs6GOHh6R78eKKSU4vJNghZ4jlk9zSRMVxSqAm4Guz03UW4BZSzhN3/qg
K0Szolviah2YfR38J/0NmoNqUjTCms71YkT8qG5JObqMug/N/19fyilkWfIq
FQ52uEW89TABgvB44vEXW0utBs2dKU4vdtovD49ZU4G+6DROfOmOsaBoCIyl
m0SmOGDj7AP0TYZahcXBKKXe9e+XYg+SA+2FDrWnPK18Md1+OIZLRGV3Yr1u
LwdxemB/hzf6glksuxOu7+mnMzLhaYCAjHQcevtmWk8NJoq3xT4JR/hZuVxh
ZWgGBxysbyQMkKzd9BikGSJhtqCAE22DI47pDrefm8C3pNmF/WfymREUUJzA
HyZIIjPIE26fUWkDn53t05P96K4KJzA1X1rsUEcLlDxz+VmFTvESYJeamnX1
7CYxeyXkKlVU0Df0RijnsEJBraNZ5aXWaycNOjHJ1P0p6HV0Q188/Pt7Oz0Q
zIqjklH6c7Z6ektWCM9AkttTgMdswpVJL7IuL8Mnyv+FOI+ExfqICcZtmr1C
6BVRFdXU5T7crTHcW9YfMGdLNwq3b7hasedq7RxgYLRzlRJXFTM833NfDoy8
b/8E13/+NpWAQJC7t2NUf4YqdurAp8M5SRMXxhutwTvsnu6gMqxOy5mzYMI5
LhX9WOzsXHGRMBfFQ/uXNVJf8wCaTd80GBqHKy1r41zEwEhT/8+ukz1WwIer
JjGTs8GNWnJ+QMIFJwRp2Qv8QNoRsCyTA6pi5zTay2CT0bC3OdXZjdfuphAI
gC13N2eSlT/FAMyElCy9sE5d8/woALnSq2tjCdEU1oO7k0QSOd5ooXCJOof5
Qh/gIoUMX1WaoNvkTta7exs1ySzBFy5MslwA51tpvspWdVou4lLG1ci8W7G4
I90U0+Ancw7O/pQifA8+xVuHfDhUsBS28VB9pZtbEGMx3CVndpKWvTCDTVzQ
NKwSQvCZDGu2f2neRnnlbk3Id1ibewwUNUJ/ujxBMZZDnIJtTMaWgz6ZCQdm
QI1oGgsEzEeIJwjNOjjmgDl/+JsPGRNM5s9EvDqTueTS4R0d42POGHcA1/bh
7mi6yGM9Jp7kz6qBu4mkVcsZrIuPN7qeMTW0FNKpTtixi4/aJu/tGLVXInlQ
H1QafylEeXj9iMBMQK5fLlSe4+eVbi6OHbwCtOsshm/ygmJmhkAo2kFdUx0P
FZzG3Sezh58EzS4Ae8NEdrWKPmO7PDbnQrnS+IHLZ4WFkPJLAw/K+D0NcLQD
ve2gxcfYoeWxm8d4A65VWEKrQ/ec1qg7m4K2Wd5QjlybNhuuzCZfHO4r/k3T
zoUqaHWU5f0DpCqYl9Tq0Gx5AXsErZYXgL0LfHG8+BpV/fREaEwqc9trRmCJ
xVW8f5CX2yB6SB0jInseOLa1CwWQ4mCHaL+ABl3IL6wYC7F9gCk97E6LQCjY
fOTyvUrPA1QZ0XdmIk7Z/nV/FeE4dI9/jhZRNCn9wRoyBGNM81GTu3NWItPg
CUNaDpKm1NPwXcGWIcA5E+Jtk1Q4E4xEjIa6f2PrqWKg5mTrPyc+YOY0UrSw
m9yU/k+uMaDYzhZA0ZLYfej4atmdES9g3+up+AxXmBxgDVVCQnchiOoDjbsW
8n/9fqncaFJkjxSrsCjGCJ9dI8uTztbGYuEcUzLdhaly8CCLdOV5xsGu7zHk
9tpmAo0x1Rc/lNUxkcb4/Pf+NVzlq3AKEpltJW0Ytj/2yloHriZi7PSLCdhT
jkosx10WsTkLWX7oybRwXqTWEYz+QEbBV7h+nz0B4eVoMQ3ZfyLgD76/0nEc
cnXHViSnr3WqJ2X+dsu7XCR0qhfhDkeRn7K1A1iBYNPuYeyLetU0QP1nOas7
fFizesZBW70fQlpKu1OuDu75pyCc1+AC2peAnp4Vj5la1CSVf20yOkYPG06Q
WRPjM7kf7qRR0sKEvDzbqxIp82GEf8DZEZtHSpN0/qQUXw+R5dVWPju9vElr
fYNPvPKf+zOKuspZr1jgDfBcfa53jucIwPNi/ovSguCGEEsocFPtpp5yvlRO
8qYTqHfLniANFTWa2bP6KwmTfe9kZF2A02C8l14Rpak7MB9ke9ZWrxIXdujU
SbykIneNBjiyo1+XcyG4GmVHKk/vu1o8mIVYqed/lhNq2JbOEr7Oa/7AY7GN
YBNA4PEc/ZNbWArjKBKKlvo3PrbXcWZGY8vlL+OcRDyVVPOpz0SQ1vMz2iuH
8osexQaW/wwPmwxUdSC8S1jVvi3JvxpkJBQ2qNDZ4XAFQYtD8nijn8DpRv0g
CtXDMGPvThdcq7Eu9+0Kyh/snF9tk5mjbCMHReW6Krg8K/EL/qC8eyADfGi8
qaqu4DwOYGIpybUtL0sHFKmGyieMjozls/Xd2ObIzvFaCCB7S9fvyU7CDbGg
fT20vUBLSA2+WP3frsyD9d7Vj4ut8/fzPw3buuYQxOIbwY9Q8V1wm4Cmxo/N
Axgt55A6FX3QPzFFS9YurDJ60b6v3W7/H50/rcWUhkpjAuRResDoKMpzKvqA
UUn9FVlDzTn9kiizzr65V/ur7+wwg+8XxfmDtZ0K4t/9F6Z0ThGG3Jlp1b6w
LWeSPvvkuQWShdaK8jH5xE/YjdW5z0U7yYK9h8WzlvcoGig5RfGKGm5TqtVF
Alr2bR8Gt4IQhOHcHgGpF4VVoY5tOHngc88DNLbdd01DfYdI+rPN4O4lgjVD
TcVrOL9lRlbkthH5zfKr8DvjRQoD6472qMDRopkXVzOcoiNe7Hw3vdDTFvcM
E9JXFmdKaZ7cJ4OMHE8W26Tad1HExXQJBp4vof8v/DenDLJFLlZoWjtcHOl4
CzKihcCBxS1wBeYZlYFylH2NvwjrmHa/nhkg6Fihz6LhzrOVSndM3a6ZeA5N
S5a18OvWsxC000hMCmxJfBIHlVhtlLAVUa/3odVSOQVR7qOSMkAJNprAUu4o
g055eRMAE02rD22AWd/kdX6F/ykqjoQURKbjf2Ot4ebZVj/m5Js2Ne4NyIdC
3tIpt/LYCVD5RLcuiOathk/lWlOya+X86fcN60LXGQJefLHwMOL6r7Y/Qm9l
B1k3u2J+kny2+46S2g4cRoy7dB5vo3+OY229ZzsIldlQ9FMzRshDdFSQpWl7
drXn0WNFaUweTgsW6KnWfrYBCh2jrQW48xRE3DATo+tmXU/uRRu9WjDS7Kb6
ZYrUZsSOVXttgQIaFO3IXwNh/ZOY59rNnSBpfV0D9BsPQxhp52D7jLv+u8XS
bF3qx7S7pdxE7KeZjsUMjxmhxan7PPzssQu0CmtJ3g5fnDEdA1m4KYil/bqY
j+QlSj0zU0iN5olyRsaidJMyaot5tWhQyAUP+zIjE+RU9sxuA+wq5IIybxDN
m+BwaDwxF72HfX9hUos54qZxWNZDrgj9BLiznDQFAQE1iDMvkiynt9eBXxT8
9Sb8DZEDyyjs+07qTKXfiiiu4pjfiyzV0VnxYNVjcaGoHvm4HuSsf96nbzT1
ddRxoO+jIs9riikX5KmYuAAuI0uiWQb9fhbkKjAtxc3DkkKsCP5nlX8/3etR
kAbUzwYenlbrJwKD1h+PC+rcs23JN3k0mR4ogjTySIo1Nt0QMbcJM72rxeuY
CE7n+iFfiGllpzp4NH1KgzjtgbCzm1KRHxKLdAAjx4F8kHVxFu9Qroi+EHth
ZXQdrs5DdE1q18WOSccFkoU3ttcCyYk2wyiOlLxg5PdxCskEeBDkkcwN+riZ
W+WvnLRLk9kUa9Rv/1mOa92UT4nIi0R31nWhe6Fwhz3c4gUuK4eRY4baWD1y
8jXZyXZCLBL07p9SZNsoFM6wIynKQ2Fww8aJ362XTszUj6WU7wkrD9jR1Mfh
53eBkvxrA+ogfUory7MIk6sG+QqvwZMlfREiTNM0XKgLu5oFFtW+d7hioZFF
fwBst4vBP0DRi3bBlZMNyBNo6yxphvwmNeUyFSdcRGH2abqYcMoRc1Yc4Xds
QnmZj1UkPvaGttHAG4KxrkxW3IeMc7O+wPDY1sz7ccOuONlZf/zV0kxTqwWz
tBXozXwEE3Y/gPzvMWJ3s8FeV6bn4Eip8Vj6cz5+KpF3h6LrRIIEcMxzn66u
2pjrrxeFzIm20cvshDRim0f2yA4tmbrgEW9k/R4qLwDgCMO4W3eJLpUidG4m
+7Z/ibBXVU5c3SgU3i8NIzVxUUpOEElO27X4w3vor/BaBWgszlqccpkxNomK
UGKAygiZcIPORW8iMskNPd1r6HzX/5ZJFZk2++mAj0ODLCHkZiR2Mc4b8VAo
sdhwZEiYn6Wx72Q3hOkluNesEh+qslfFsOpqZ6xKEjEb3SRnwLa8YmNx0yaE
HbPBX40JOLKLjeUilpUdc5YHFQCrSaFDY0vhfLsIlC4Pe3PN2bM9p24Ghxsd
j1O3K69OXs+ref1Cs1Glum6jSqh1FfDznmCoc2CGfUWBbj47+pjgXyU0J7dL
X/A07LwawJe34/a0n0gCcKgKJ5/uqfhK4msM/FmQN73FSB8Z5d6pPpukG3FW
Cr8LzMUUxxJfIzgI1EIoMPWmyKp+M2ivEOQlu9E5tjqZSRyHBGIrgR43t24N
U8T0cM5wQCCnZ138ZJabwyIh3GhtLRatvJSUScYRLS+gHxp7VrZClSnVcT0e
Ol4qRds/oYkVD/a1zygUGL+Yzg2+q0OllkE/4ttM8IybHXDQ5ZdoS/2+DLiF
KKYMXKVJBZVArC23HBNxyRu26ZXkka+TaMwxa7tpKTFOkBFTBcxmVN6LcGgD
vcTMnKvmBbuJY7e1YwPVaFlGr22XGbV+DxHvUfbcx+ZwJvAr+KhzSSAjfvQg
Wb6437Rp+M4jR0d+C8PPj0bVHTvcePJuRDag4JkicX68Nhn12BHkiIDAbBrM
D08f9QTCUcn1eEd8Jek5UmC3WWEnoc1MYOU9uER1A/tEguQdDdqL7C+DYY+L
OEIwCwHVETugsUpiG+xApSXHPt7OdvpJmmkv/Ltf8UlHIoLbBLaYEU6ZFT6O
wqF2cFm1S9FGu0wHwYlKtTFzrZEVKUevQh0dvGp8+kxkfMihgYfBWSooPG8c
zk3BcGS0Bh7tVEnUtkkcaLQhoEbIdL4/5b0CSIb7dLxMNYf2wjj8TSFQ3GS+
g+V/Xt9aS9m2qtiifR3a88q/cx7YApUwFoWEXlfTw8QQDb/e0+kdO5Vd3F2+
jPiRNmETkHL1n4xnN6/ImPzT/Se+Fwe+gVEm/RxH/NLlIurhipK58zeHEgaQ
hxViT38F32Q3RNjqMRp6/faUc7ixWK25FXGFEkWa0wRWcl1IRSuzqUja6acD
jSbOmt712BKr/wFjtNzk1AE6yjLUFQo+e5t1S+uEytq3Yb5ifNgYlGkYqfW8
SEAZ1XbhjuhVyEu1qZdR9aAJ1Su4WaD7iTuJZokKDREsCaE++sA3WieaLJCW
yHDIS06BqphfYGknZumOhfGLlL6Ni7/MoQlNXNpgoSePBZkNs3zjcWjJ4aqm
S5Fwrn77BoKjyaLLXH3wjXxW5em8RFagSYzt5RblOQjjBiysu/+T5u3jUz5k
P2wAn4GnbOsTMtfQxmTBz28uXnHxh53OSwotn/AeTbstvEWeE2hj9YrRupD3
lmBQDjL0Aq8thyAV6MCzKPE700+d/Ohb6hYLCYCPSCy5p5rNvLuyktNy253T
HLimFTVM14SrRh+YnQ8+lS4zVPcU1z60/TiAIQN3yecyJ+dgGFdBXPq7NZvH
d6+wkVjbZK0R9BctkCJVlLHPScAvQzhARFKePzWylZqp9Qd6/5Ok/IYwHmpg
n4jykCDH4I+O6gBnsoHMwMpLIXjzi4Xf24fNEHfc76O6nOrbsZNcvMSTERvT
q2X0btEh4LUDI5f3J+FF+p/o7/soUOKUlovrH4NaD8ID7ui8Fy50xI8BLsWG
o48JJ5moCZU4nDKNFmG54bsoBNdOf7FzK8LySTOT+zGbpTITvQHlHAKRNF/F
D0kvzZLSpFADsYFXpud22NuVQi/31FBe2pj5Uh05PItj2i+oQgKoi+IMYvIr
53nBDechVz3l/if8M9fRV3/pg+YyG2XshjbSYFL33+ZY2zWb513M4dPB4BxE
0VkSljec9kYLQOMXK6tvfgCowswcnz6MuMyK8wG5jcaRL7L+SLWsS+/R2YUq
qttNKcMjZiAfPjXxdgDVyIVczsUXgANdQmyR7uhoHaTs/AN0IkokTV9ht+3s
ns0q1Cc5p81LmVfUZQVWs3JEFRIOq4ib6/LRO0oL/3RnUei8ouhZ3ZECaogQ
qylyoV7w5GZrQkGwAJ5aYsipoeQ/O8Jla9zDUyOEIjxZ6kfvrOowYkmwUFcm
zG4U1IGPH8vTE1ZSmshk1BmpVdeRJ3djHsiJ0ZNu4FVQB7uu2EGhE1qBST27
3Sq98d9CiwdC777qWqS5JQ7RbwBYRxIUTu50bX25OrYhP0y4cSPvftKLu7Gb
AoCyt//gC1/IrVeZH1eBxTcaobv9Zi38LXVLxj5YZsUDHf1KqKXhR7oAYiOM
hzJil55TehORMERfkFhhYktPE7MQFVc+XFeFAUkT7ovAeRNqoq767N6LtEVx
9GGz5v8snp+hwIh8Jzqc5oDyG2VmkIYDYvIWM27hJdUACvECKy6tukQV9Fi0
Q4gRuo2DIL4KQLjGWoAH8dC1U5U/PZBIXBNNw2lT1p/QpEOyCkwu0lPLezhp
Ql7FAxMeoHF4ggNGNSyo1hM8Zn6EsIJfyXXyPjaTZMtGwEYTnGOpSZ+cqF6a
d5pMB4BzqeAVjr4k0L1kHwToGvrGjNi0FKDk1KKTjnIYfdyuv6oGiYU6tXxY
V3iFx/Nuwh1ITP8pzcaPvydj83DPVUzPTvewljEkZ2YXWy4Kk1rEs9PFiEYV
ASaea8OwTit/l4Ezv+gT0rec6Qh4jk363ujF+et5ZSfRDmvo9OD6WTxEOtMq
YHJw/76kKLSgQluqzdmUt0iwabWcFsBgcFhVRY9S2nEZl0LqB8AlP1tgTrTp
Nh9SCSscCJUHtXMRVUi5I30WIiTX6EGfIW1JZw5uXAypGaK8lz/gMVOI/LYV
6KkEhlJUlapkFb4WuvK4FyYGPceTn5yyox7M3xvDInYLWPrlHmhbU0rhDRaY
XvMhlqzT0fXBxpehmijXnnJgrWse/DJFFrza2QOxcQ9fj0L5NBia5adpOWFZ
NWsJSbiJhEide1J2Lsi2Y2XvtSskIUokkqmBeBah6UlSZ0hwIKJqIPK0juWP
5hOkx7c1LEc3ijKMWMigqHGVflM+Yj2Wqck4ntArOi3C2Gr6iipZYxCby1Yn
XMQqKbD7xCqMddGVLkQqVr5Pn6v4R9GSOWbiBXwpJ7BGW8lAzxZ5i4Ptnnq3
5Z+8VIIqqNtzu2V1MUaCSNfUaKlAlni/0bQNlpu5lPql+ic6A8mOVAxL9TLH
2vdimPJ/peYPz5DT6zY3251whRNufqIyd+50i9v7HZ2kLY7RbG1t8SF1jaJN
Vq1/mp4H28f7hUcqn3MJX3KCzFNbWhRt7xQP8KIHrg4UQOUk4IJFehyh0GfC
GqzbCQZGpPY6C/2tEdTlV5xYmjpP7+4cE26BE31WS+0Tkym6fgInecxea3y5
H6RzuM6gHI3oExyB2p9eeQlGF61D+vTTTq0040sEWyw3W1LTaYn1XD6RXag+
PZixm6/RHliGA1BN5D3A3WNddyR+6+3BBLPmk4gcO8lfMNj+Khtf8MBKCAbe
03Nq1i6L7T27qYiyuZkqz3uKPRSIQdMNIqiV5/JqIri39J4kMEO1oOCCjGPA
L8Fd+sCXNnVWeb9OFzJAcZUKdseMRdvYKZNcDKXdaQHn0u17sd/YYQ9CoPBq
v4PGtAsb/6+V2GtBwgT5bdmwl0au5zB6XYKv2W2FnmCbxou4nYqhteCf7ZpJ
+Hrv5jk5iXItUlsC1whvNIMB697h06sL0eG89Gst1D4su1o4DSdIakxFDy7F
UDsM1HepERiVtLJCiW1dv7Vzt3zUYFJpCiA3M3GSedeorBAEGFObjQWnKYOh
FXzmisBp8i84yMtB8d/M7nV1rys2AD/yzFVkMjJC5qdWshoTVaRSa1Ezyang
/+nmTrPKPyCvsi0WZlAyQe7sqme2DFlvEmmrdfAobf56BrjeFrHTlyqRWRuv
Ce1GA/eudSZ17CZHCCRnsqr/OdBdsOX8UU59Tfc9bcJYPziz8fzi98cbcRg/
sqtUziV2boJmVi0tQuOnApNliDi7pR00l+yqlkecwcJ9lOsqcmvGaoghfOE3
UfUjqsxY6X53YJddBfBs5zEF5b+Fv8bE5v9pwaxbNqIpUG/hgLBCJ8ZWCLH0
Fr6UeXGsr9KL6TXpxde3N0iMdkcFTMyPfMYJWRfXUzKZzXFfpK444m5OuzaP
RF128QNMd/XCp/oeCXlx8SxIhFrpgtRYdz8f8EuIZnR1lOdIzwMoMv0dZhHb
LkFtOvOr1QihopkYFL4N3yOV7yhurtWnAblf0HZNCFyELM1Uv/UCVzaervfz
UDbxfymeQbFTdMcJNdGkVw/d0k/pMXHAFrrN6hsJ6ktfe0x/0t3OSEwWoA6k
22ZhXDUXaL++UvooYrjkhHVrSuVOEN3XPbKX9CauBvkPPE5fWSYrpJI3HVzo
AcLNWeQaKV++PEF2paKkqWQdyVMDusgeyC1LQpHzWWVaA2XpFOpabBHdBRnV
Slt7V8UhLan7+Kq1ad6gX1ajGqChP7EvgzEAeCmznREP+DXkfpuYHf/MSm2+
q2OOVgvEWddNpJihQKPBS+rBoJow9OhtmoG5yQPFbcxJFGTbRA7OQl+E8/0R
l9bNdcz3IzFOpzZskDUUHtjtgm9va3OUdApkD5A2HEtOM4s+t3q7P6PiKdvw
KZJzexid1YkyNvbBfs8HrthC8HWCQzLSjG7+jX2fDjUr3of+kF71O9rlJxyC
6PzqV0FP/uuoJN37D91aHM/Moma9o0Bo3HPd5HF41x6PsoHoO/P/f3wJgpIk
htPNUXrxOzju2jSDjq07+/DbcxQ5BP3URc5WqfC1dmBdzPg4uUPD+60EjVUM
91wGARykuA9GcPAfDIEHX9Fu8XuyvwRbzwr+f8Q1JR2ILqELlaPXkrcQQq1j
7qZq2I3c4ZndNs+hg7GMOhEL9ov8sK0V6DcTxLuyB94KWwAt4Oh4wjuW9gIi
ZRY/StEbxsHYhdfRaqH55OtcyaNKMoN1qgmXEIftpjp5lMvO7iHYWThaPq7O
+Oawkl8Dy9awU61Hc9aAhdheDu/TsquzVG1ZIHds5/hMG1j3ou3lZtA4z3Yk
jJ+8dDVioxjbjy1CUfFD5V+TZoGHWCRQQN4mll0NO2s0XOC0hvwi7zmplD4+
zCiwfg0CgDdMQRKMuIaClTlN0qb2w4X6K0MlkBzQeG1xpB6t5ZqzE/Y7A1Vh
/Uo696MzEyNUybfEMNyKoFYqNAJU0cSXPNcayijvX8EYm5+WZNMvXyVJBZUF
MvrUHnCXnuNgsOAGfb6Qceo93H3IKRhZCYk02cI52jUDH0UGpRB6ntALIdRU
a0n1CGwTmqGWlCGspRKIkpTxIHs+67CYWPrFcfQu2N+8xIRmeOQPJ7Y/hmPv
9qJFtfwPqoxaVIwBzm+NJiTGGtGBRHhwMvX6WZ7YPzKbsvGys56rXK+Ua2cx
/ijDemiX6buQbnd9Z9eN3160ljOAdPHFKIBCEBXhOyafAPPK50hmOX/EUudM
BmkaDrCou3r5FW4HsOzfKN3vYd5OrBQB8pEZdZRSvSfRMmBZ6Q5VHpceSErw
cwn/cZa06xI1m+2pLYIIGAwEvtdWyLcpHBkGVsBeAzOqOmaBfdPArtgbbn22
dtNWZdoPMZGSJfYKWaTKm/bxMObuS/ei2wasEt+jsvKs+JCGz8+QgGxz408Z
QsUZtolYM3jqk+huxQ1VHEvGlsPd54yR2cebOgu3MItvT+gJCV0YZ5weDuUU
hzNkx18jGL6FVBaRLOasVsfD7YYgY/bxEw1RRz+pjK5vjNgJi0nQGUoS3QOh
GxNFAucEqEfIfZgdxSVzar5YlesZRuNN+D5pe09XWwLkH++fNht6UgkABIkT
X3XTXhzQuv98/yyzERJ/XPns1Q1fUkfdpCm1gEJ8nJQTPc2l4TxH2eJTOjsj
hKGoqgtMJQ3sJtbJYgAaVs+K366gWWRb0bBNHgAJf64szB+Jh3bio7/wihA5
4x8IZjColqdYTg4iNIf/F1JsKUCxucsRe4uOQ6kW/HiOaawXTXHjvNtDCW3k
+Is7YjT8K1C8bsyuvYDTRipRNS1nI9VG+ZxVITg2BjUnCZOcRhfSRbgc16Mr
qE7EmSj6dwolzJ7KNCMKnMJxCFwrdDoehSfs+buPyrIEgjyH/bejWBdS9kfj
9+APyPAj2erxvTkdi7C8si7CwO8aQUo8rAOMXcZzLZekflkl8BQX+khkLe+i
yZg44E9OmxsAMpjOHpb1Z2kAFd3fGSoT0uA5YczU2G8veCbLAjv0lPfePSkG
7JHDL0uI+waGJVQXZOskqbFi6fj/hZQcGuGqBwInhIxZF1Aqb+dUZ2LI5hXo
xFR0apBg/81BVETf1h7xUfFbwuH/THj0TTco/IJbX0PGXLnL/3AOtKEaEPEo
1WWtkTHdHRMTnvQSfE28qoR1TP5je3ogIoJv+fwr0SHhMg7XcXiyEOA9xYt2
Is/UBkgm9qtraKEZLTq1/4G5S8bq2/MrXPDKD6pWk+SqdZHvHp9VxcXRWBkB
mQt2z/01UxvzMDDfPZ7EoBsbM8po27fwTNUKZgbMLERmUp0yV9MIMxX73zK/
FGoq+he886gRSIHgn7ApY5YV5SFD24C3GvoWqqeUdZrzHqvglFsMvK8K5Jlc
zE9Z6C9MX9ndVJCZYbLOhU21Zfy0UmDyqu6pIFNpZmm/IMsAS5rDYWvmG/tK
EUBc+UjSic6Gl3YxK8Zr8ob65hNnUFBbseX8CksnlEGnE8UtZlErHXDf5+pj
rg7trLSUPnEfqEp/NRKM1RzWczXkr9GLpUOCnwZu3HUn27BmmstygqAO8WtQ
+T6KjiYMgsV2TrS9FRwvVrCNMj+1jKb86om6z2Bc2p5dYhZC6xef5oV+nW18
GgsmumPCeV5EgWtuwbnH/tXrgqc9MjozRPXbKsVsaMZUKZDgPjIQJtEbgUto
db1t+1ZuULmSi0YbkplcteFY7fF6QCOHKLHsMBnGDZlJAVmSFJSni2qB3ZM2
xfC+q0KqM3obIk0fJlOmI05LjqKKpSk2Kfp1U8s373kIaymEr/NO6XPgDjh7
w/XfYbghMBVt2dNv1Wb9/DMtEjCE1huqzN26KQXsGhJZW4cjC625FkjX7xo+
bfCWpDjBAXBBapr44mYi80T0jec+ewKTnjLjkcY+RxHBKZS5atDbsqRT01hz
8EfFI0z2ShMkGRcIWQmVam1AhlH2p+6gSrXZ/7gSmiVf6txG2yEcR5yHJoKj
YTMA20N0UqrwIks3DMaVNrGTPnJpavAWPXnuzJ/xXGAdv2q/hMN6cDmvNWK2
nKVNCgut5QmxrteMAxRK6hJS8OC4x0RZ/YJm2IhxiBPu06qPoWNOMW5Z72+5
HorzFOoWgikynbJCEbYucAenMNdyKe/rcDOJPoo7uvMrwE0MOetHZCeWuoB8
pbbODdmP6+8AaXuN/IHDf5ILkKI/ZnucWCNpEhelnuVL9b8CWAtumbJ33B7d
MT3DC2MruUP0TJtyKoAUhBl0LUm6UjuwZLEqLrk2Vel2TAFdEFnaK6bcYIsY
WZW/mAE9bGbexUc60la6vDUv3+NxY23t8zrgJwrqIDITZdyXIirgYF0iyR+/
MUS7mYUtZ30wLc1gk6pZovI9RVng2rqdzOcEFZITqcS1J49xagrJVzfqxMII
8mqjG6Iti5D7/7QjNvexQTwHA4qTUFlAeJn+VvYTk6PNWUgQqEO99SLXGIb9
67ob0GpBxIAutB1BY7HV2s6kXq3afo27HPRFZkUfUdhN4F92ruAQPQdzBkRZ
uuJ8z1cTo2ZbbmZMskRpz2uwIV9AdgFyN0FFU+FWLD8k6c/geo1mvbT+S2at
Sa4wV4R8JjyfNm1EPIxV1j0woaTKLlhdu0kWE3fmoiexeTYk+4Pd+sFxTy5l
XCRNxO2XPslAySBBxcQpwjvqAH4RMSZZcmdvNNPUBUn5SrK0n7KVLMaOnuIu
U75Ttnc74VTUegF2MUO9srBpt8cKd6hcfyLwle1Wfe/fUsehDpLkv6Hv1J3P
8TCFXUE1jFxF4puWNIJcaM6nc+klo8wdmmPHXQyf7v5HP8WvLvO9Q0bHgrpv
yLmvbL3y2QChKxhjSFP2BtrI7C7SgtTZOjIxmH4jJDeqv7oJVCmEQ0M9kxp0
RJBu4IWZmA7acNznvUmGk9szvzvjwUz1dz60K+gkMs2Oc7XRwQCLvdp4nn/8
9C+0h2krvP3rV3hHELo/2cLQlgQb50E7QgLrEUVOal1rzieEnCoECJzMvUsN
XO5KXiKdvxNVN8TJdSWrp43LBz9DhLpmecF+5td3R7VeuYRYH4yliZ81X9g5
Q8QJxPfFMlmPCFff4+3Ji8TGhcAj/x3fN7c7PnWCb7bKwWQdQa0QHIsMiHbn
8N6Y2eDWWo8iO4ImFclPFQdAFivcO08wtDtc4HwIsdvoannw2ZSG8ITt9S1N
kPCzjehP5Ig51dCwdZ1KE7JztgyKB3zDNYU/SJV8TIFJM1RLgXLxQiwxh8IV
Pz4wlFdRyFUMQNO32kdRL522uuLdlEOVLuTsCwF1apfCz8b1OJElwAVFWCQx
7cVHMNtISRk1Gt5QHQ3oYo+zDIJ47JwtoCfHu3r9j/21nYXap8LlKlwifsYJ
Jt0ceepKom77wir+kZOtAj2nDQzOrL3PMTIl65SanIefHAZDxRpc0mdiVbOf
MlG2VSf/I+mKr/m0yncEMJsVuLLe2KHLjLSmB056T0OsuhJFPIclUmqXNaqt
pUcLipXzImB0x1OljDfujAb2QCETMESj2JwmoEUdWWhjyhgoEUwoXHTXrxeu
cggqZt68XgSSt/pe9EDHDB5QjPxRO8rOTVp3cq6CQbNTpiRqhzTnwcxuoJfH
7oPoS5egjawZ2xwaEYkPTNPEdSYdoJzE4yalacVVGbCfThwd+uD9LV9a5lzL
jYD6yAlV0elZ84mLHhJ45XDuES5CYtgzVbez3SoVF3Bt4nOK8ESeJRZEhv3m
uszcHz7GB4C6gmTIzgR+kymYq1FbwcwWHhX10XEEnx2XNOm2IORIntjKhXnN
gv4yt/xjR+gvr5LFUI2TiCJ0Rf10KXb390NmTx5zIWnvj1BTgvrIMDEJ0yML
xuW2HM5jwtwACMmy5o/i6XFUyAWD7cwvQGSjchK6JkxIRZ2zRsBeVOrZTmT7
Qc20UyzPzZQQIUz0Jl8RJh5e+A2G43J/kFYhgLMtz9DaZ3DveBTOd3lNCgml
yDdpJb8/bNHcOPApgunKJlPJnovHFudKvont8pK7BGZ+6GSxZzU9ItSrjo3z
VtIsWsGacHM/ChnHbUHjove7fD9UR7nS0kxZ5j4uMmS47jA+5iURP2aSmo1v
q3EYtMVMNEQuY3P5nX74Ey2PzHQrzMZb0ppG5i0bFzXGqDUWPKN+dsYu5nYh
/xKK2rLn8IbGOCYm35GelWQyrZKNNM27+KSNLdtZQNb5kMVqAshn9Gds0Q9Y
wJqDk24j2juvj6yxxrcE/6qNBR3eRvrpZPWXCtjeqO4notWG3SqC16hehkgm
57wMBQ24XX0z3W13FIkgOqyU5bCg+KaeC4kAHwp/8zldf2S9W3kqUdRMXTsv
0FnjrfIl52k2DpLUBUL3sTFY5FCL1rbMAVWJZ0ZNLtcF6967vkEWIEvR61gR
VUTYPr7sHAEk/rM3GmpOvbSBSNCYkDNqHrRLjLfnSbv7WO1nApDQYLIEX+mR
K279ocZ5auUzjk4o1G9zKt6SOtPWgT4HU+AcTVD1y7tlwfDeYf22eQin3k04
qIT2MOJNP38rBwbS1R265KTjoV033/FhdE5rleEoy1QrPe3aQnqJBABwULSE
1NgLjRh+/h99y6B96OK5VpyrideNrzakKpkxe+5VBSwYORIj7dXrEAB5Lco1
khQIKQPqxt/UIls5ao2OVQIaW+shl7SiNNgGXaiz17atm88+55W+YJYHHtKa
1jWPjMtxtDi8fygR4r6j5dRPup0KoSwm/2ScI0hdojQgS29tA9lUYLkLgcIs
obAWUMzVSXf/6gyBTAwPMonJb2QVju6kX9kF/Eh+OnItnk9XzwhKmAQNoDI5
xW2zi3hj0TaamQQREF7QONJQjUJUcg8ZntGXEPyseba6xpH1e+UgWPl7ir6t
n+nrRsrOB45/fC+4fIpW5OhSuVIkHIu/oWHnivXsQlNTRcL3hQG/+7J2nG2z
OaiV1IGVLlfbTCS4eUigu3NmPCGIFYCNHE+I4lEldyLBWFwDLHDb4tuV6s0M
XXATHXC95GnL2dQn9A/aloUVLexe9YuPET/IRJ5djUBFdlWIP63VjJzj7z1H
EokLAKPwweTE5QO3U9hQJjHmYpgfgfSsft79Grf8cognXQxnjxRh1o9zYpxp
czBHwAHpY1qj2HcMrNTlYWSmU41voMCNPmEsXwt69Hb0uWvrDL5UH12PalJi
9avVgmcLfN/tiu9mjoYu0HaCx4DhIsbkxdDTxxU0GzbTG1yXanUlANPbdTMt
o1vVZJ9y3SmbO/99yJ/cYkXXQB67e9eija43DVbX34Cwc9F8Sh2x6bhVVNii
moEmnGzron767wd9JZzlUH9MT/kjzrWt9IoXbDPhnb3chwSPg9Z44UgQUyij
OCriDEFsmqdOB5a+2vXCR2qtjIwCPYAryO1o6aRUrbSq+0KUlUAsSiM8kJvN
scwnlaWFlasGtQ5+B5ddKgCH/Hm2uWXtAlS6uEhd8FfSNghj00tKJbOp9Y9B
7n/WxjrsAXLQMWKwEJiLApa8XwZ+rRt6fcColcM5giz/bH2J3kQgNJduFuvS
G0vouwU2XnAGR8kW7BNm/XzqB2Uufzn6Hza1qY3urwMf/vUKn25YP4zsZNP/
3fwTiGPaNj1CI8co8hgXkfy0UVTGgu0jz2E/yYVMCwmTDZlPFX4jSGdK7AQv
qEBx9opN5035/DxyI5bWtO15Q+9piQpBjAz1mAwZALfVUUzcqo8YqpQin/sV
J8TCTrFOXuo2gh5IxloxsQwd6i4LOGeyrdCG/Ec7+88poFonUKkiSqW+GtBA
7jRiFhawDVAvYUEWdMhAJioXPtytaWIS/uNxdAdXggTwAHhbCvvmoVZC5pgF
ibNd6iBS6hrlsf863bsTUInHHclkg9PT/NRM3HTYgwPwFkbCYXKhHMCJwlJ2
/8z5oKoeel8/H97BMA17lAIE428MBJNpWThx5agvgKM+JlLzhgNuJVKbYXfr
jU1TC9dWQRPDvOR2FEkmouVY6lEkGIFD+YKXHTvEfbleWCbbh//7BxUqZDkA
8G2SSWwRGSvIZ5UKbM8DnWX6Ew04z1qtjWFHBPWpTsSSmvzt7mkmsp1cD8Gy
k5sn4gcwRn7+mzFFZ2s5OFgkPmgcZ7s54bycvGQgRnss1ZhwcCXYinTzSWi5
h01PrUNKpQq2zpG4Rypdct/0BA1EpRZ95gPY1CG6fkp559bH+mGDyAZmaEkh
oAAv6iX72NXsIaKiviwpVXb26vexU7T3Wpij2InYTOqLAqSDBukp6mgpCjVq
KhpzctnSz6r6O4kO5I5AAspEqAaJPN+VPeYRse+wUcoe2oLU/jRJcilsc9Rc
c/44BZyXpC/h6OTxmPua8bz7VqYBce0YDKtQH4PDvZrixYkM/gTSnDXuwrip
lqwfQo2N2fKPzb6mceV78zs8ytt66Oheqs9SGoGlPeQUp1++GmDOVLmhc7gi
eN2BZm7HVI3XJW4+JkFiNdv7+o5jBbon06xZZ041wnJzeVls0NgRtDnrH/WS
5BeEnsN25caRLib4IjsUlci7QlXKiNr4CKngG2P+YIcZVYvKBhThIHleqBfY
Ca6Kaz25lwgaiWF3jx8Y9GZ0TcyDLNBO23ysX6iPXr48qTPEIbTtnQ6ey8w8
6qMbz3WVBPgtAlKijECHilAuQWw/dIUpf1cni7neXGeYnZfBD9Q1mVKQT354
H3n1wSWzhxCxyCCIk91IMtKN+7DJLvwY9v8LMSnUDmUeTpfa6Sh3k39hjoYA
pWAXn09IzBX8mEPirqb6/jJUi+kiAZXAdmALgzzHsLxr+uyTjfCSnfJdHz6v
COYoqOSK19D90rsC5xAe086IQhRJBpFnFQqe4Kt0iKGsRLpNBJqhmEeoFBwy
29eXbV+Juzk4afVKWXNuGpk3gFNAF/zhsNmu5agJiESuVPyPzVILtgmCyHjm
YC8Ut2vE95aJe51CTysp+GcXXAfHdPuWmpwNy8OCXB612BGlCMi+/XD1f+AO
7WmzOIkOIAaoTv0zcPkUhOZjHIAjAumbJhA5ooJGcIO6FxMRoITkQ2aAIYO1
BT2cvdG4MZMuoLEj7Bq9OUVk0UjqSvzcxSnVc98fRPOkfad5qI9BY1KyhA1D
2J+a4fVwWqJXLS/T0JdiphUm/crNXTsJD7+4zHIeSk41A2/URglkxNPaKv7x
yjydzxmwyUy38/FCF5GVjWP/jD99UQSwEO7TTCgf3E8JvZN6E6lO24LVfnDn
SaA/qSSawTF8kEKpy22nsDsz2g7GRwHR5rN6EneLYNLc1TFlZS+SXNyDE18C
ZCcltqSDoijAPhYzhPLa9HDzqS9NsSXyeCdYUjsulFgEWnc+adcctLX3WXq7
IofFY2YNBr5h9lW+V7KGPA3+azoM+21GfUcpIU8dkIBO+6Z4btAF+YSTVQrP
aLJbYe6dCgeZOy6pNALiKnfIL3f0gCD7ixLNEPCmam14Hfytf7fZ+0tUbAoV
xbWWV1tojhTztsHMIH3/RejXoIVnYhCSNlHKe0XkocKXi3o9m80jsLYDdvkN
s+qWTDoLuThzB30+AJNXry4ZXNkInDG2itzWwYRDg4JVDH81j0oMyiCH/k+y
jkF+UtCmGKeVIGZdgV5OSzxjXxUdhAqxeK3LorF2fn8He+/UDQq1rVsEAVvn
FnnV29Z9uPyMx/O++AbFeLIIVTfWFYAXvAV7MXN4YTQAgxT1SzQn5chNKEqd
kH+1Zb+cLg536LKUyqHnbBr7rWcxAWNP/KTCmZIFgiU0xgERdWVEXLPsi6u+
kejcseSH0nM7lfITyZ1Sgm53xK198CPJG5nbkER2T8oux3rpz4AYzXxAFNZP
lsjlUAvfJ94VUjklwgOPpunbfciWL8aQWJBDrOc9TzhMDpIlUGaD1fIjuLqq
yNcAhA5wbm/X7O+Z1DMroZyXaSQn2fpAPniKBy5BhCj2Hem6V+G5d7g9UDXl
US5NnHwrhusomJfkU7Vzk/PpKyEo3u6q53auuc/pU0x2I78EsCDZ74G8w0Dq
DDLI7YJ1HSKdEWQg/cAjzI1y+wvexp20238UHU3naqLXMTNuCv2Q7U/iimZJ
yz/j6SJ/zYVdfW746ZEqv9ws8cfx6fVBT3zx2WEu+DcD7VtBh5GYJKUg+aqr
96znj93EeGcnL0n78mS+4y7RfoSW6cP9uMkk7MdHUdCebY5a88ynVhYzN9wB
Ze9ufRKBnMztQ3b3oPfHC8tpYzu/75PiYUd+yVZtfuGZHc1rfZnXgvxlY/wj
TudBG/P8jAL7xM3DEWE/u8DyLai6UCBRIbvi/FMPhc3yBpKiA0yqHytrVa4p
LhoYKNEUU0x5lJV3JHejSPVzScUxaa7AqalwDm6gyGlH6/tznWjAHvi9cdKi
n4FC6bRiDTdNZ/KTae5uPdOtZa+7aWBtTXJC/EN3E/G5NItEaHCraXrhMKRB
LpCv8KV/KuLGLvW1e9qGEyzeeAxLQkgiIUxtJJCaWP9nVLAMTGHOvG4CbCD8
mNWDWuBUE9gSsAVDiL9QzEG4ZfpdbcvOdCZlm2Bl3lQL6mDiA2Tx7hfn6MEG
LL9yP2qL2x1Po0/URm5V14jCYntE7/t+GLV6nkIKPq2Zh49yLgNBGVM7QECO
vzyWz6zT4Q+g6zmiUoi3jIcEOpDqSsWHlGRRfR8BQHzSqxD1PqzcCpSW3lxc
Mu+dfFx6JfZuTzYxY5nZxC8tmn3yD1wSzl6MFZGV8PWJNgI+lBJtkvlS3Zk4
DkAf+pvGrdezYifM/9gdByfEdWglIDliclRF9LllPVRkDK3k0gQhLZVX+CRY
I/yPsTupM6jWY4X1uQDsfj3RO5AhH4z+SHuH7zv00oWvqY7UprjyhxKDTLu4
Kxg8fojemG+j9Snc+ClhGzCUrqjF1MbQqUMofMqdqo3Lx6aUDRMkJn0jlJtJ
ipTdV9fZEk8MAYGLR7DwDNbbJJRB0z46ht1feViLsWIqEVmUWUeQPHc3IWL+
GcF57RgwIPz8mJ+q2cqhpJiojYenirdaPjB/T06x0tSCzpnhE/S9Meb7SFyt
zRtRntqqAHXDJXphwpc6cem3FAxFHkoQM8Ju3e4fdL0gQ3hhve08HUQrCyds
p/Fb2fxeVh9UiyyassJ7aSqpk3+11CoYDIlUxgbUTZiJlOcmkNng/giECgTk
KtTRg4cnMhQScy7MQ/6Cn2Kq4EMmWIya4A9ZF3N1wqdEu01yGIrBz2LUsidg
UuPRdQVJ0BPAQJKLHxs4MDbo1ZvGhygDB9yqr6CWCqltXfgg8AE5fGDm2GJw
u8OhtndGcFrIcbMdznoCGpR5ygUO9d89fffuUEZNeOHrAyuiOOVZG1qLyf+E
fQsqJBdhQdIDzQBkec1BayIaqWY7y6KE2+XiRYQadb2Nb7pX5XMVivO2L4fa
X/N9XvxmUwiYJqcGcEMvesLrfy5+O/XXPWXqLf1CCFLDXQw41tupyQbmiRTv
mb2j0VZUmq+8wKo//PrUahjVF0ZRZBCmUN15ak/GUw1Kd5EA11mT/NCkswtt
k+qznKO7Q7uxaciXyUArt1l1vwLjFe0LfjSRymxG4GZNX9wlV4DFsUB71lrQ
KhIftVe9Ksfy0STP7r2mGTAAJ+JEM5tPxAMprw480zcecXLgrGUND4fde/3C
suHxO7j4YrQ86YPYVz1xecO0J7spQdEdKr0ypjUua12SmpGJAP9j/Aybf4uI
Ikk8BCaIdB/fpOhvGmj5FzLLAA9ospsHIi+MrRsuY5XBO41zTChPczx4uQpw
ma5pB3P1g8CXRzj9cHnCDpxle0FN6k/KqifXZ981+wdqpjjKRzg7t5pAuAnT
iJv+I8+bpMB5Qle8UjpDWLRC83VfRilL8pJnOrpRG/T8YXFf9uSVMjS6K6FJ
TJgavpeNch+mQ621GUIB3aQ7HjcxHsfMO33o1kybuLM6sgdOY9qXO6MgZkkp
p7UftNwAMyps5lrgK+1VPk59MDecSxWEB5+wPjVoyntOMI+ngA6qMz1HTy/c
Vu9sv/3yS3p5a9KO71l/0dsM7S+gLXN88LUgHJhyxP8VvWsrLr61cUI7NWXf
+JTmUBl9Qxjbm7Vpc9THxRyy6jf0lrpf2rWk/4KbBL8b0SR/N3Y08q8z8Q5x
Pj11FPbor6Tk/CLF6QvD9ishaavKnGCWd58awsOvBYc8PD5p94fVYs8ZIRPL
2GMxBt0sKcwi4+Qn8DkUmIXyN0dJGcB9LPoGkuOWTzhC1J+Yjzab8HIW8mtZ
14oZlwQZ2LbFUAS6F8/7q9W7hvo4qn8IZ67JVIWT4Hp/Xt0YzCLn0vrz23nh
FthOJn+I5rhKNIukE9cibP5iZhLhJYCMD3OlR77Cw4uhW8vVTwhR+Navlotk
991SyLKRGKZDmzWHBsTTmjYKxguTxpJ0Oekx0BYV+hN4ptWh07LNBXXetaKE
jQXK3QW5Pp+CRUHm7f+TN+W6zDGScipfjQNwXK3/AaP4+5JrMb24a4CPBGhU
AKU4lrxNV8TcGjfWLvmXgTV+0TQdV3ZKoywo4v0ws7d3pUJBSHYyfTAvLEVy
PTiSQhRdDaB0JNPwsnnQtA5I0R3zmJlgKLowFwkItiZalZwqN1QE9s0mUGzg
hXPnRM1ZI4th7xh6mH777yy45WKXhKPXVrftMhoXKs4AYwyFh/zQafz6NBng
TVpBZ80GvQnGTuDm2F7jy1RO26WVt2aE/psW2inqjsqElU9NcseTzysNwVFL
AsxhlXkYR8wtbl1xz0PZLWv+DiaL4BTFBTR5c6wJTmXuVyPZMq/xqwFpG7ja
dqJzR0dpfw/mub3DCF7JDUoeb6xsZoouookOpTZk9pMwVZwUaW89+vvavTTY
QrnFDGOjn+fwUKkdoS4do2S29KZx+Q2a8CIpyTOBBbef54jFfLR2e1hfHVnK
9SjcBFWaDDknwOLArhdS1I5AnNtoEd+aki6QhnF2TUvgj4/7Co2oZZt2dlPp
jsU528gBJyg4PP06znFObPbOiKjnJQsc/O2/n+IH8KglE3sB4dpasD9Q3KM2
NaaUIjFhkUm5jxreyW7qw2iaFHZ6NJi8rjU9JOX1mqyqo5OXqDcvpFL2ot7H
QSmfCafJHtoUB8RyrDJfjvXIn9NR24SR1981rDPc6FW8XWRnaEyk7TKT7iTC
rSdxDkPwcql7ZVuw9Lrbvw+uG9XTTzHIho2Zn6truoqIKEg7k4MvWamA7oh7
1RgpwNQbssNFANvOpwADOheUz7kYO14f1FNrPCtEmMM/YPHZFReYjMSXZjuD
ibEmzG3/a6aDPU41I2ihcjkgCUjhU/vDMO79tr9GczYR3DAbsFxAKS2lYrnq
A7OnoPK0yKUh5t3AHBoenRB46SOfobixsfebm2JPloHB6TQ0ef4mu2oWi0RI
Y0rTRONypiNgvPk5RizQIf3q7Xhwko5v+RUWBdgPT2lGqwBzG449HxMYW2ZC
Z36R3FnAhDWermu7Za8Y96cPz9+Z6kyichkXQu2cASpzTPkiP/48trMLLtFY
jmPQ4WZLUlmq1jNWhMxUIvQZTbYqEimNueJdqCfEDwETzfbXJxMBTO5ZX/kD
vCpvRpcL56bTyNgPBDMxIMY8fhQDiI/SQcRcEMRXbfPsf8MgPnadqxoc7ucc
2tZ4qIHPFUmNn0iUs/twrF2y7fC748oe0t858TkCILywO8VW5CIxZbOgXON1
RSJpovDq8APOZmePyKp0sBZPswGlgRw92iadq/JYuOOGrP9TdOCQOuTbpifz
7sRT0KmrcY8qDvNCkvCRFwBcciEZbwqhP7MszW6oZcGj2peXtrVtuhS6adI+
oYgsFcBzPM1KoPVg+YX6uEBSSpmF1NegDILCWDJYYyFfcaDgl5Cbzi4i/+So
cVLlNQk6vfG71WNdUS/vY+WrY75FxpGfUCaKXfqKMcno7PqBNNIMoZZyAX3V
Solvuyqbek8GMfExdZqFllBcFYxBlK2obDIXSF3TAcCgI/4IccTE881eeZmW
yzpGSmWjh+PO9Whr1qZ00vqbJWP+1lr2axr1BAMC4IVpiAkoI7ka2Rr/G0e4
vEbMIMzIi1Jt+m1LHTwOF15HRCMQcJoDcYw+prAGFawJoaUrIliWbnwFQglU
gjzKhKPDs85I7lK+aV+syXIFltPnzmAJM/SG3QYRNyG/DywJxjo9bxookv6U
hYV++GfyLz6E4LUqNX+N/TmFeUl018KylhxsZ7AzgsF/AfrAzwn18lqKtiO6
tvPYQMA1v6czgkATPBoTLdJwQKl6peP26eDoa7YQzZVK6SHZcOkZ8zKwI0WP
xXMr6XappxqQKHcuHdFsYCzmVgUsOkctReaZXmxuneEqPoiyu5jHkQo0SDwy
nZibVmhgYMDlpar9FFXhEqdQsw/NFmTfefuApruFQ1eHo4eEUd/vuxvW+z2u
gEa67U1yiMBeTgbsywlfcLur2X8KH9pS2rX4Tu71B2pcaIIJlCqg3dM6bgPE
ZPJl7leelLvVqpD83R/vw2mMuS5QK9q1qjzY+AsLTGYjJlp79m24OYguL7VG
zviWhQ8KBhRn2ygYTfjF/YAXH39CH7TOVUNZKA5teVUhhyDn9BgjfASmnKxv
VPDY4C2AXrZMnpUgJWMB/Fv08SQr/65WfxXgdE9qjlBIf2XKJlR5MKdyBoOJ
/4FU0/EGOQki1e4PhS6fq9EkJ1pGhBzGQbOFOyGErHap3UThuXoZ8Mp0lGj4
PLF+tRwuu+TYPLU4JYpGQFElPJhk2sud1H0B7+dZLURSmidFq4+cyCsB9JtD
Tr9OdcZ5Duy0DPM/ytN1y7OjFcHVG6gc2nPiBspDOch643TD42ClmdkTBWsV
QRGpLuk2laEfUTL6cqk7dEOfzjBgWCbVo8uvaFJwFXU1KRPWEYVBMguSMJwa
ziD0fekMWYjF7J1cahV0Ak1vwi5f2rAD7ocrpDYuoVx4tqt69A/h5NWqOKzO
FZR3jBq6aozogu+rGV1Iy85qLQ+vfQUNz3PaqBlDShnlpZhLn3sVN5CTBKYV
3g5vzm1wUdjxYUSKDa+9JTjTc2CbvkZgNgcUbQWGZI+qwUu7KWN7VSiRxF0K
lqIQwONiSBXUeW4LKgQk03qrlg4UXO5XtuFURAohG9+DZG4yWdFF67KH5kul
ny7FAVEeISccgPCXmOUbWgU7L34RlDWhBYbtAFfUioGZThxTg8sYaEWN4/YA
Fcxdv5XpWww/L2sESx4I+yf0EG/OdL1rbEycZqqaF5Cq/8zsQxx6CL4qMEDy
3/Wevu3lAstMUCRGOOunAiIyhOYEhUI7Ds18FFIeOfCjfcmzVmLOkzZf6jjP
F4Cfq8F9QYaaovHFI7LlfgfwfviLfVXBIIMbXSLCHhm6EhdVTV2GnI22PXE/
OE0VAsE+DuhqdYp4/ykVDVRqSpCEHqlroQbMZtAPYw1c1QSJLOiASniLIG4U
1rAT1E9aBNpVSQyqB6UzhRtAZdGqgfzTFSkOK1sXrsBjCyZrsN6rtPvvHw+n
gM/81RTq6eCd5v3tb577MwANNFTN8xbYv6IiEIepi27SR4Y++MfBuLd9NyqD
eXJEP3QaZjUL0GgIccecPHtXp/B8c1jbZ4OWp4xzqhZvQ4h/YDsDTK1KmFUR
dZFbKOBxG26VM4efhEllM3h6sdkt3/Uui2zrALnuspEhupzbgpLUVIRev2JS
fbV7tytb15lvSYK4bYlm1prRyE/bcQ0DSXMYnK6iHoaAmDbNgIUy90b/Jz+r
vu2RV/jxKV9z+CVl1KgjzIf4mHahW5pXzkVyLdC8uqGOWGacabsJNxcb9F7M
0Ea/V9CdJvQaDb4M/uoDXD2RX/vgSRv404Hoycj+sDOG6dcNJBaqXeozFk5X
kE7acecTQC93Gt7zkWlUq1lmY+hO+L5O6LCK729HK6VH8BW74j7MKl953lNx
IvglbnJUQUFSU2BXxsvZW+YAThyO3CZjcS4S/e1MnL4nwGOf24sTEa/yg7qp
6pzFEZpPd1eb+nR/TCNtZIrZ1SU6+RNJOF6KGbxWZ0eVAL0sKN0Ou4pJ2inB
yxQrFWtl+HnXjeB9yHvZliLHUb4vafiBSuhaXQMK2wlipmHVa932lKkbZ3pL
1A54CMG7CfVp9yHW+GvFfYyPoZM0bMqMrg8tsVjPUfh6DrM4ThZjRQkcNUCf
Vw4ucD9DPchUXr1hSX75lOXE5xuWKx8VtIg6jQxC4y4tbjMbcGUmfWqwTB2P
dL4aFDp7HFImWyhxIyORPWS9mNATnEnmg2WDpUEyzTH5yKT8ugqnRgNgWGwz
BtVgTN23Ue9JXxAwhhptZDSXfdKEbLPWNvcY27OenaT8Uj0YK3iLdpqd7yw8
N7kCOfxVpbl5jqjfJ/hPfWimerXePKoWvyS2SMRtI5ZT9OzY+HdjgDplP2/E
qcc0DZik+1c1lqPd3rn9S/CDbhvH5kpN1dZzTk69ZeR9dOJx+TPSqskd1Tyd
K706Ye4uaNmU6E2DEmeXjxAcdY9gtZOpIml/99Pxc0ATSuST4r7CQlBNSUFt
eFWUHcrABaVoBrBwaIyHjT+8VSKb4hyxwt+do6zLAJJWJ5ar+kxd7b4nIJnk
Qo3ym8zXt5ZTyMtF06RRH/GtsaehDdJDdNX2+gT70T+StxKrAV3cwrlNi222
JzpbtwoUWzGKKVfDcPWmVqDjv3dl2XVc8eFveo7J6wLsPI+YZFVeLU1f3HEF
/lx5QN+OK4lQhQJhwi8+rf0iPdnIx76TjKtqnmLT6/iQ3UZqGEP9BIfqe1tt
16cDlaqgta/Z2V+RprsJ0Do33/r/DPOOnwFbxqdzHSvoWBQG8m35QYNLQFRQ
Qz3nHgtpYyLFc+J+Uh/pD8CvC/uZh264DgOdfelmyysCfn5+SyppLDHheV32
iH1UQgIFZX9VXmdg3NLreYkrI3J2j/lISYzq1ARk+tRJ5mX3ZmoGZAjOcExB
I3z+4s7KX3edvzMl43RsQP+oV495EatcXPWvREv3SXmj8n4xJ8h/idA8/OUr
GeDhXn+2r1EWgx5XoWjvgNXNjr63ZohiZDIlx24fnctezV/2EOP2twXz7ToH
BPJoZI7Yb5jmOi0DbK9iBSpTIgps2mEPEXDGf6LSnqy2jTa9JYhPf6rUq2NP
MtsudD9G0zZoDTSLk2pQH2hOJD0HV/MaTi4MVaTICXryywKOdAIDbi3+rdMX
TSxXKJ09MMf+n3X7erTS2NX6r6BZzmDKV1djhjEe0Auwz4FovjJQn1ORJjrq
LNFwQbKn+lrBSZHCZ+Od0vaa1ELCk/SU2Jrt23SwFBH2QlJZwE6PBksswBB7
dRQEYiBNtygfhnfoO/xPvQ2nXe4DP1ccd4LYvwABKZEyyygwB4tQvE3UAmYH
00Y+a4WXFA3+XBfqKecrdWgtfFKtN+ZW89kVeVz2F+wCSK/Tb8IpYdd9b3hC
09oy8cxiI+JKIHGmCpklV17uFkF1M8J3cwnOksgoOOSPPHGJ6PKBn7yvEp9/
03Pg2ZTmUHtr3VA2+d7JnVCvpU6pgbj+UBX2bBL9PwS1DeytmQp3AVeIk7Ec
VVJdQTjPxXjszBQZlR9j5Xnwf9iBQIni3ldhhZffvtwis45mkcfKeTN/o2Qv
jMbBZgTnZmegJSrMGkbrlFJyDtPNanMdbFVaIAUUyK7dy7qk3UAX/R5RnkHj
Narucds2nik+SvrURBnzarbyjoSq/LXx/cuSZ8Rnrhm/VSnuOJn2Ha+9UpyL
IbYgxY1Gq1iq8WaR984o16vYs55vDlij7S3+35Xa6xLdexNwLEy6HFzafAP2
K5oZFA4ykmB4vmbZVypOf/jJCSgX4RF21M0txf3vvZsfUmkTM++xCrrKXNFM
JIA5Dn8gZhHyekzYCP42awheIVe9e9y14I966HMOrrfvyar6rkDNwcQZvLER
Kqkhz7z1J3qAVRs9Zu1XvQ3I/HUq74Q+NQ+H7p1XfMphiF3nciLWUyr8RVzJ
z+KhTcktxz/0YP3tQfbloCVfIEJscQ0HrPZVt5DqaXQzVUu9BE3iVaB68zlZ
S/lZb7W/qqURvlPN3wEll1iHK33MEnWroMZoerHlO/BSeUPrjiGLf93sk8eA
GK8Lr7s7xGIYsM0RMt4y1JwUe+T5RY67lbN5X8YzFVNek8sFAsIirGzK3VBg
/HdjTWJCno2GIEOG1eFMhypJxU6wBBkxt5xzyY2nrJlyaESL7+9hcPokcTen
Ri8R5Xepxk/4n3J+7hYrLC5aNwiU1knE86Nzm+0z3W5h7I8Rkpp0cywTRicF
VnCEUMs0KRong6RprzTO/m8+jAPhNGkz4Hi2Snu/q0+CWY9VcSVHWZPOBhDs
jEvAUkI0oN7JrmbVCic6ZxxW4NarhopZktiPQ4ZUP+3L4XaZ6hmm+esBQsUP
qXAwlA9Zpj+y/B2QEpOe0TLV1YHmGa6aRXNg69OlLRbaxEXUC7ovZgZt8yIH
ULW2a8JKQ4Kzkj7dgrHbNeggE5u7OkovPPMVKmCovZiq7jvO2K3UwEqogXf9
x6+y+VmGFRvUrXcvmZRBhiMWh9ag3U8D1gkefV6Hczxs0ZyZe7/tiJtajiMV
ZfKZJi0SzglspraiNV32HfZBkSj0+/KWF1zHawyPsnE83a5oRTS/h7sQWDW/
RvSRZwQSpuw1P/DWwauCQ9DEO93x12VZH3xGVoyiuuL7KWnKdg2wwIj5kguU
sAjtv3067J4y23itfhYfJFyNRAQ9b6ekFjjydVxN/1RAL83JDeo68kT4FfMb
zo45u/CXKA75IhpEwEDoDepcEJfh065Es7mLWJzT2+GgMUrig+RBOgCZzZ8D
Y8qud1oekxQTSU4GICptUobAG8DLouWxjuupLQ+GRlh+NDZcUPXZXPoupWam
qazfJ/jO8IHpD76R6ZwOe0EQF01Z+3JAyqHajZaFlFfWGaKad61tvE1kgCr9
PDvuvm5VsEQMh/UtiPfYWy59gfFpxtpiYRq9WKaNQFYUueRTBi3S3LOS0qyq
t3EMVBn8UgzEROyAkXFnCUcgc6pfWjVyMQ3zgTBs9emy0YJgjQVlkwycfXQV
5zeWdRZKQA8WoVLHGGnncXPAzx7jn6JT+ciMXuucls0/p35Qi9ijaxQpU9LM
6cFSER01s1lfLyD9Jd0/pRdADPSrojAskmUvMPe7hQMDrUPqlXU4SiGTSwrP
w8M83GC/0z0xjziUqT1YrQy+eH3Xo3toj9DZufd4ETTdKZ1XsM83o/RjObKk
JKNiIcg6pZVRjeNzTKWRQeLwlef9K/RZ3L3ON3g+zM2q95zX09t9fR89v5Rz
PTZndepGpE5ncOXQ8D7CUoPiNNeQbOV8AOJHAs3WQ4juvNdM1JORX+KjSAcY
UHUFfuvOKALzQtvITfBmWO+WPX7qMus2U7KCD4wyMRaSK1ajziWhWR07J3a2
NQsAHF8LyCe22/v/3D6UxENSJcxUfEteujglzBpyhUiJ+LRcMhjzt0Jw+v/c
b6r8rKx2kPTAChd/g6xAR/xt0IHK0MGcvIAbCg59JYFWFNQOl3ifm7bVafUT
PjOrz7iPOnVuP87RWZk925WV8UEJlg+85A6z6qNZzhyDlWJJT0EbwCyKhxNR
Fw8kYIXbZklihwWJiKksfj1LF8SYRE/NCF2lXJ4c/v5NBwo02Zx3LRE8TUAs
VstEnkWu20uZ4eqlzMZrvL3WqhzqduQyEYg/vb3zxca4dFIMVDbiibXtAp5y
o982eetZn5dVoKLMrm5usWwGERWQIPDCt2V4ObOMC6/cCI4V+RjAiBhicPqd
eRwnko7iKCDQhnxLYZkvw/TMcvz4pcJhltcIRSePQMmFl2hsFSo4O2X1cvio
q9TER55vml5y/b+uk+KjdR1NcEMwcmA/mgLK2UqHPubekdW/eHVKwsFONDD8
yZL7aXwF5vhaTjz87ouCVDihXBAMkwJb0kKvphELuEDnRbbIBozaFlYqKxwA
HCJDAQR3NKChcqRQ8ybSQ9ag5ckO31Z8mSaZQJjVz2dNJAb4UH4yvje6lEx2
LDO6nDMYU1NV5uK6h/VZwLwYpG2JZkYxZbgBaSxRfGUrgACPNxpKBJfvNjP+
gJt99Y0AMCP2d0jaif3yCgYK0EiepeHLaYzyz9Qy6DM3auldmuvYlVNo4b8F
hSIh1+0nww1sIdwi/GE3eMmcCBWOOVu6LYWDotvc7finwFhVOWFyKjtu5T9m
9Vh7IKP/2jAkFbBewe3K9fwQkBncvnlJ4YB1FRsqyFrpw5KfEQc3jEOcWqIU
tY0jYL9Qr7aiJksx4PGwdMWVvQF8SQ6PrcS0D+u/XwzyV9f1IFRqHVrjjDEi
fluJb1WFwVlkUMKXx7XGHT8yJ552xtSvqvNbGHrQluuKgIyPuRYlKUbklnI1
Pm94A7+36xpV7BE8j/DI5Nm0UcUkOrFBKkY+/CwTt21vTO+ZxxtfxDY/nKB3
2zdB0YwDokLUHxGWrgvllKXLrYD4uTLjOdGbPUci0E5AcoTUg/lkk6PJzBZV
yMoDbilUD9C0FV6QG1qWqRibn+9jli8DnW6lX+JbcMwFsPXg9T0TnZGTSAYS
CN9s19ds8xVbNZptcpELt0UoaEiPMC5lwHa1iF7tx1IqpGx96oJiAf+95qzB
oGC9cspZIe6KPdkhVko2HRgJx3bpwwDpG8+DSBhTKgvWtiL7fY1qk5ctkeIx
E+4uSCycEa8pGF1weBJjD1U/3udPegm35I7ewjRRSwNCKXT+yn46iRvNtJ3J
ETBL9zZpii1GsAchBEVA8mt6jZg8PFk0CC0TGyyB0u9JWLZ55epC5zlHo9MB
bRKvE7ykai+IjtgLICi32xraVCpePHj3AzWb7yVWO+tkykxdAblVhp/ggorS
uRiTzWs+qkQRorIPO2TdsRyp2Us5MRONKqlE3VWMUcRU31oedK1bi1xAYu1O
9UpFdhP+rjTDJKvuZPnWEaAZoXqyelo4ZeSgFuWkSEZAIYQtVIFsHW6j1GtL
1Pmu8wJqFp/I+f21S8M5M6WIGuVJvJhVlIt1rq82awkeQAJMQErTUyqQ3SIo
yovNP1Fw7N8A18e1qeplpHJUa8w9Ht5BoTLVA3sDAsTbbVPCmoyEb8dqQh6N
C0YG7ZBlorpcJV8xCaMHM88wE72TM09qpNbMMI79ZWoQtr9RRIoukvgGh/G+
AcF/t27LS+E99Nl05fWu4ikc2a+fw+zUuMbDxXByQ2nGxmB3rFA8/fRZcDQF
CqH/rB0l49w6u8bq8r0ka6YAUAngw3E8nnr6I7fHO1QQX4a4ecE48KGO1aXW
ThiACJ0gZaLBlej9sIzY5gK3tkD0wr1g6xqA64VEJjNc/qfRkoWyurJLiffz
HVe8QceMprOmp0Q8BlcumRR4/w1QTqIcjB5c1TuKBAyR4wGz+EE7WIYJCDvs
ufUM956fvEoH+4djgFqamEB1kG1jnlal+SkBQWMVTe7J5IPBKgt3qmAJK0Q2
pRIbX8VNo+bZ3yCQTh2fahvULzPm1rmcyF5DDQ7z/MsE+rvtFUW1SsK1/Ycb
UpSx+OJgIIjmj0vxbxZWXcL0BfYSgBim9582uWDHUZuJoYutLhXcI/yj1Hgu
ivUAS2PLrPn0Hsm6CzUidJ4H5Z6PV3ZE6gImOTirs7bpKx8yJ7/YEMtomzUb
3edArNjjEQ4A6hUgT7lbtcNwhxACdU35jbWzDENlF1H8L20p+swSO8z7pOaR
mBTUrvU9lbfQ2u9ai5iFh/DUblia7iMOwKUYOj2tflCJY8OR7jYPu2WSELFI
+UIJyhXL/WLQtURpied12SXDFsHnuZZ6Q0Kggkr+q88wvCFTuBAJXEeuIuRa
1XXJ9hmpdFlVKaCxbZl+JT/nZ838jRRL1S28oXZnJf93KpRlcKeBPDgByMgq
ZYPY5GA4N6SVgsp4FclQvws5kBVGz7WElmL4+wFcWx4OBNLA2l2iRTvDuHY3
nLWBYJ8685BgTG7CgPil3dPYdiibMSFtQ07++fieY4cZDJCODfies20+qr9J
B3ePFgYlJ/DXjA7Q3bGz2aftxIdB0bgPW26SDeee8p7KOluJOSRJgn0lanfB
/9+NozdZxmt8A7yd7uFNruDDFWEL3qc2r7JMHZdKKyzIdChEo6bqHx4BDO+y
KloJQj5NQOQoQrS9YKhRwB+TkvodwT1qgmMH5ZmdQAKsdEfSbpCo+FHjrYII
oYKOPFeWmTK0XW5TTch9bWVgg7huO5UL6AyyGxuWFfdGqtZrmeAlmz8t6NnO
wfe0J4mvxC2O+QT31oiybaI0W4HCmOZ1BBTHCZYJ4R79CnGzPw/1kcYiaFkw
yEzejTp4/26jmnzpfXiRqKSEgf94XfwgyZ2Wsrt57SZs92TYNvUebL78EYIP
Yb26NtDYHa+6GU2jt7dJ+STgBzMfLluaC7qrKLod5ysQi8Ayx8HIKDnMJhcP
NrkllmorA0l9QlhIJCOLhwVroFqbaanuA3UoJxQlKf4kCBpkJUeo7FP+qEjM
1o5hACh35rlZQtLdFlJLNBy/Wmdly2jelSmlAFGE4Vei5XI4PQdrFs01cmvj
WJfMz6TydkwAJZt9ukupwo0CpdTWL5nHgGMymTf3wefLk3w6nnYf4uNQDZof
hB2busnwgHArEfnba7RET+CA1/rzb+qA6lZRIJAAWpjUW8DaoUDSSjGMTBRi
LG/TSD6gfNC8DJHpmCKJQPtNUijIoFwgyHSjqIl/L3Wutpi5l0jwPU/X9ZkY
9MCbiA3r439KAqTymQ+pKl3OOwTq8LzDRM4Fudb5JOZt/22I6MZygjy05XSu
0LO3+3uSbfo0hejd4H6Bd0FwP8Q+bEh/RwT91jB2cUMivBv5vg9184P8WsSy
dJ/FlqdXE5VzEqAtpbRqsrXROJa1iQxNet8T8a0ZeRJGiKh4moT9wEV4zFAw
Z2bzqbYHuQZGHQwoRlfKmiUo2rBxG6//N2JY6Gn0pgJNxw+QW0/beoxLpXC2
0BvxoRSfpZwicg/QESNNDFfzhCgScghlSvDGmjv4bfNyQRAUaw3fgWcEe40x
hFgQsCB7h4BrPzhkwANJSm6EMVa2xXinVIKjrMtt8mhjTeCMeURSULMKPRob
a/t6O63TyCKZdl0fSnPAALudS/zX1lS6yaBnXfHwf7sL18Q6t+MGPyNfcA9C
3toVxK5pI827rwjpnq1uvR06VJXTik+AK/1czLPDVIQ/0GstrO7re+Xbz/9d
6mA1jzemWEiAxUKu0omB24orVRd00YHLpLeMezS/6+2wSsKpQdYFZZTn2uzW
M0MQKDT0beE+O4KTA/zO3YoLbNBjgWIO8AujeI3P6mmz60mHMhTa23TxFjJW
Q5to9lAHcrZwil+VbEl+VaqpAyuYcBqveDLrOvl0bI6l7z1DPQDVgT0OPVZa
uJUjA0IRLrXIwW8kR5GQ/puiwyYFVCWTkUP+wLvK8nBsK+hrshY1el/xFRtK
4nZx+EGUZxN1vUkcIXievWbnQzaPDdrG/nQY5x0o29B1oDopxkP08bq5Z2rs
hjZVCI3+3UTCFyai1yxN2StWMwYhBA0YKuv14XX9UA0e/9mr+9uyc4cDcMOU
WhEuFGOaUCaDQZkgjSPVJt0gYHd3Yw2um60Xh+bJEEbmsFl0zx803Bk8OsI4
WUmh/b/7M6Qu7gM1y5H87PpV5hIlaA6Op7Z+4lQ+q6jySHROWRlSq0pE3cF6
GdRy7X2+22OyGHIYv/4h41Hd+DTDLTb256t/ZdRMSI/r1qWo/cl9/f0+4iAA
8HcB/jmIo8uTpt6z1mfF1ojRp+QinJIfvSg0YIQly9PcK1a1G4wY/60aeJjo
FewoB7gLhh5ls3SrOefRoAVNtOGobseMMjZ4/FZlZ2LkNRv5kE4os31PM/5R
puuR3Yi+4yhWcG3huGBIXBUB5qyXhyDCjaKdrvkIF0Ks220UAq0HBLFB1Myt
lLco2T4x+RNjs/AINdqFQUBvXNwlN4ymdncFw1j+TDNzEQK0c4B////5zZxf
qJTwQ7enfrQS3hrcVWKDObv+dCcjAS4XL/T1O0lWdKthQMPZehmS1ZG+BEQI
Ubr9llD07XTYYSyrkx6oL2UwQ5VOiGCnvlejd9WL1Xc6e35MDvDh1VRSo+4b
ntvH6eCGlA0+/EVASKyxxnM5+MZKFde8m8OgJdDRy5XQW8CS/y6LPjZqhK8v
jDZw5Zm7qti+cSzd8bnAf0fjZgUX83LFwNmxPQuKJojuTtFmetCUACQELKgz
E2XzQx3AH2sxjw3oVlzsjW6QuuOSBmQy84dqzd4eaJ/QDKC8vAKmvOU2Co/T
Fe0KmxqdR7c2DTPAoJdpM4e3QOBWEv94FgfpuD3qPVsXJBVUphDPSx/AoyFV
MuGpEsadLR8y2Y6aEgpMtdnAzS5BFfDCf7z3EuqgMmxMEwPGhQ6LTc4N1MJM
nujCsA3WU3zg740pEZFAM7++TC5cfgmyHdMxgL3Wm9Iu3p+VPM5sEEcLm/bp
1AwzNTJUaJgOK3ZKFqz5267P2MexxP6UeodcaOehK9qToEa+Eyg4FPOb7oF/
VEGYylHmblCX0qF1ko0kSgymBMXzVYtEzEG7uYzrR8K6pay4A04c779arBMG
3W6R9G4a/JV0ApWk4Ry7IAsTsqe2A8qEWtx8l1W3pU7wG8VbXVEQKN2T4WVx
4JyMajOLyYMckxwpNXZ1XEEl3xpxQX/OMnzN1glaJ/BpfOGyb/lK3WzkcLSr
WynQLyQ+TaT7E2JCX6VUmA7qCwBu+yGWI2iublQGiP7Roifl6NdsTGfZY+22
j9Yj9vTj8q1yaIu0U60J9RTQ+4MwPTtmub6Zr+2chfSptmOk/8MojxyR5p0J
XanSbO0MzM4QZ1GZFH2aYheqWqQib27WT7fGbGH4hWB5UEvZGworM/V3PZyD
EuiBeZX2XUyBRc6QfewrhAOoYWr8sg33Q/5UlpBWA2vLYufkvjobkWkEQEpk
ZIFmmxmkzWJLifQHCjTBylsXQWf2r3hfhJjY65Q5hb2/Gg7Jx5W3ZLbdSx8t
gUxsVKNYFaFYaQflGMqPR4FBjEisfx5x3vsv+dkmnXBtdpsq66Eityd32gKh
td9vzohxWLawPeN2CkTt5sthKR59F5U3eoX6nlw+iDosMymXciyRsy0N7itb
uKg3ZAvcxAbo4X4gJh8tyNM08WIlrciCdLk9wBm1OUwsIA+unAWLltJMJRMU
V5DNyw3fudoMdtryZJPgvAtHeyM+C6cSw5jZv8sbQyEafApQK+7e2S19yoMZ
+duOrFV0lHPDbauram/x0YfguiRQcfkhkAKzW/pFqKgKbSgSagW5FOWU3TIO
wV4EyFxFo662r+w4XAtmBouv8VNjZjBB+kI4OWTrPgl/w+a+RtfGYwm1tlnP
Npo/bT5o+gT7JozloAa2YWcXI8NlxX7I98TC7lbA0C1/SMubm7faLbBCTklU
QwPgaIhk/DcFeYXvluIiqfkVAas2YPDDMyLrdnhqEY2JwdmWTjSSUHII4uxJ
pa/ynsGvxDUWjFDSryUpVIVBegP66CEwGijS7yaSR7ZG8maiZRfS9cO2Kf6G
CZb/MQyOMLlVC4iOM0I48cZxklJfImEm+vPlxn6XaGZBBkJcE7AThoX3EqoZ
DUTOobF/N/60R5h8xRmPRRcGZI7HjCWp82NdAaMCoMH4blIn1PpOfAFs5yQu
d9pwni8okWnn8pSo5K9SR97JbNqvoQG+bKZ+alBGUweySkRIj0vyOg2nRmuJ
1fYBSPnAaOsnWo+zs5SKANdZ0+InUXrpfGBaYQR+se6rnXu+wuBoh3QSFeBO
l6j6Yp4zeM5r7gO4PeZUVWHB00YDY2GW8/B7mDKVXHuwBB1ThYgg5DqMdG1S
G51bBNnQhaT43BEfHpdgF8ezwbQNFcblW4Yta95mhBMxQGO5rZ4HqsxhyhCK
HetMRpt5HX5XSBIdfenbcvjXz2JfRpg2knoe8AZmdJ7A5upTd7p2DC2/VkDl
EwxUMrdzaxcRm/dxNA1epqJaGRj0C3eEmUEg1oQFGEqb+kBUmzDO0pDC6ThW
NKRDJkuuYNFo+QeJlGGv2JEDD6HkdBJ2dM89HqcCYs/kCSfcNH6NgSwT9SE7
0RZ4H9866Du+YV9sIvB896qmRyvCbYK8C19KWUsVugxq9Z0Ic2/meivIQOpU
77xltYnaHC/fXyYqKgZ+QFaNC7ub0AZN95F96EcJ0B9iN4RAzVoIl945Ploi
8rO/pnWXL2WBe+bCWlQawvNaNYacktYSGnvkOR6+w753HMlKDqK54vbFuFnE
3HBvyxgcIeyeG8wYQ90o3gA+QdPgW0p1ubOcnMzutG6Gejt2duKrZe9w0aug
231PIUUYgSdLit7VbhFDFz3jXOA1ve3pWMUL8V28I8huuU3fUh9vcUTjQkhs
EHUWPPvL7w4wK6PCKyGqpfEPxj2zMazJJHX7gSBdva6g5uwR52bySKgcFeFm
v/aC9UfwkKetSFTAPVG2Kd+bWSwJB13biWgwNh677ucHmUPJX6sEBIEcWetk
J7BnivWle61nO+j0y0I22z98q8LosvNDDkwA720PB00bw/wE1tE3pPGB6f0D
zD9aGETA38mbf/niHiQq3aE6pG/RRSdNvIgpgF8PlRn6hhcLzyfeFt0GW6v7
uKjFbh1LV9/aKUl/Hkw2NiYz0TocRzRVmfxx66mGCK97YdzIC0LSnBWzxjuK
JSxSJXV6Pmh+L8Vz4nKsa6+333r2CzdWkOQpCJeSEgmDkf04y6JEAC6Kw3CX
fhwkK+V/BdCmtMkAy85DrmZy4uT5Exj9Ah/yO+I/Rg664YSnW1ent0sUoBPo
P8rStlHS2cuKqfSzXBTxpqf1m/1KyYSXN8AkYMxmWyixA/DPCHI86u8Y4/ew
SnhCTMTJAF7rzzCc2h4JPV2F6FCmYkjNCdfQ4xLsYr27ruvaDVD2wAVYodZK
DneybDOcJYSPN0CwTQi6Z+XhgA8seQX1t8mPDYP2uicCoUw2uCa4bukLeYpi
zOjrg8fOue18SkQ0Hs+sHrfM2QXPeFpivikCvZR5NLEdzqhpuUAZMlPp+iZx
RzFjgRAOaOu3YGTTb7ck74TsLLaAO+7yCsl8Cbkq0W+xRZQbmo+s2sToUR9k
RPA99BJtgYfSvj/RBOX4wXQifU6De5tyRUJEt2EiKfgL6fuCx7EAzPmXal7j
vZ55nSfTsQHvlaunDlwHwzmci85xrjTm1xs99rWnrTe6047vRmBa5h7fltyi
wHa4hS5xM8KYj8aJGyY8E+6jBPNBH3i0RIfwP278iLgwuUJYVo1GFcqJQs0C
offggfsQuCBn8lT7GgYvdZeTXaJqp8FVl4z/39blvrqKE38x6Z0m46tuQ2YF
+ui+tVbngCCuWcYb3rdg3SCme23d4w7GnCmioiVtVtOMe4n29gmZ9ju0hRDn
4eqoR2Zc+/l1OktZC6WHkE6WnkLC9a+MolLOCEQOuWDnDvkHggEaWcn+9XL9
eIQ2IeT2plI6bi8Hpr3Voy5TwYtpsHRn6oDY78+7oWXJU/mf5FaPVypgcR3W
8075r3oPImuYGoXL1HYYZEsv3G6sU3JWDMutKxxSkclRdoP72LpNLht3IMBN
LeY47YkHPgHCUcB5QCgCFRf3voF1HE3Yp1K2pT32yoPD3jbEKy8F4sx0CbCs
XRDNRPqLvWF51DiGN8CWmDEPWxh+M7wvozNSrpJQfOw5YInYUgqqYPXZcAye
0k2UvLzfK0hC06VCkpmfpt6N6zS0GLuuxK0peU8xV7fz7X/kKCIfly9kz4ul
ukiX2TwzkXr1MoAZg25kT4/2YU0itEmQhcVq7HtpgHEtZap3poM7zsZdvDwg
/xhPkisxm66kMMh/D/XNQdhQlXw5DL0vWpxStJiTUzXFoMVfHkhDFOjxZAjI
3LiGuq4Odih99VGxOIGpXG+rY/r6McgSt3fjsRDaIwjPzxr8EPokpH1i+56S
F/ZC1U+XWTncAxTIplQFMmMzntmUzN+hy6A+hX81nuRCBs8Nsw1cE2q12XBd
HhzDgKKER8HvkeuxoOIhQgpPXg71+Ojxc8XJsKzH2QfeUWTIgaCsT1nFg7P7
5H+kt1UeIs+YWQl235rnid6isHSyzqsD7sC5Ysva38DY8GMiPrBudbWy9D5b
z7QqY2zWdetEZhM+MsCCWTWzd0HNvWgpX3YCtefadxY4QxADEJo+i8PcN5xs
y3Df8T80ucr+nWoutiN3KHqA4bP8HEqAMK67IcAaSaktLFiDdmXj5YNx5BlH
5qUR4I3e+2TIdvkIV2WGncz7heG2QWTvwNFaUnTr2MuRFxCfJq0FYF1lJp+V
WjqBk0mfrFzIlnPt/pfRGePw0p2MOlhIL+sFCbrBARKs72iQN9zuIKOqwVnK
zI4RmMR1LH92GjjicL42uPZR3CBQ6LK6v5b8SKraaIcsRdDFMOxtq6W7wAAq
NX14YkkEC6c3t62x49TysiOxgh29wu8uYmtj5uvYN5kZeuqdjrQMjJYHVnkD
Y3RkyX/N00muD5bVyykbjpypps2DSMbkHFvUxgRzNcQn2L3JCTjl5MnLvvx0
p+nRXLPeA0GwARCUbng5d5GDZMQo9W/ycoIEdbyFd7kkR9rSPE2tEStkKyCB
twcQpSRumLu+AkdcMBB14qUvla6XZxnoJn6nYbqVRrn7WYxc/+11Ah4UGrDT
AcVmiBGDDjZfenMZqE82NmjVA8BA3FHaJo+prk9io99qyT4sQwYzk/fHao8G
8DhHgXncITR35uN1xOBA9y5zW808UokRc7yTwkQloqYR+j64T7zPD1goul7H
PEOu1h5wk6S0G/opEo2rxg9EcWsOs758Y6pD3CmQfSbUW7KvToAks1neVXpi
TAcp+5/84uA6Ye+Rne0LQyMlkdorX4/AHj+XNK/PXdMMd5OGjpiTqtU5KFr4
PCsLLKrYfEGJd3cfi9cZPUSRPtIK0gUeKC6pAzJ04CEc/b9mBYncPuNaAOk8
ue9F5xLMdS8aoB0VjUuB6ZEPl07JoHqE8vhw0AAZyC623hfSSsto87c4cUfX
HH/5+09u5yEiVzaZ61W1F9OHBVQTAzMTV+tYBN2Ww7Xo1D1yZ6l0CxtVwkWn
75U6p478vaI+tjWCTP8zoc158gTS9mFHlOeXmiKHRC55fMryqyYqvLnXK0cV
/3ugsPoNATsDLnjYNnptd1EGANG2gt0Z4qK1d8B4CsQMYR8RZiGZAcmSViwn
AuX0OZEtbd+0rfGx+9dlEkRzw76T4qj5s162O2OKfvJurTTySJ+s6/2TYROU
RaaaUHTy5BmnFJuVE3otbyoBkHjwoc2RlrbbtJhKp5D3t3Wtoh3dBaHi25h1
vdCNjc3gxv2ISqmKfMZPEZX+aNVVH9ABFAgkJ8h6HFtpmFVOiHTplOBLnraA
KiQRdZbLdcJhH0ct9QtH78u974r7vaHlRsJCPxMFuQeBjc0+QlpH4suR+wzU
gPVlVptUTwynwMp+LXAh3ohyvXBmFyd1ZrFbs3NzfZwaTMQDWTuhAe/bmm4n
EwmBW+IQAL6UAd/QBA2gDpxCUOIDC+pYcKpXtYDSOGOtvjDGgsj4++UE1+Fd
dj7iz67bP5IFfUBVeJBmQoSF+QkjCZzvxe48p8flXFTyLm1SZQHlzRHphPCJ
yjgOuw57Wi75DG23+aoAGiIXb6Wy5y4u6RibNM+nfsfK66dJPMo5y6JOCF8a
fkJUxhS/zSwh+pU3YueXhLc0KG7oc0CmPy5+fyjclqYM6uV2yTbHjbXnu89E
JaM2gp8JHI+xDLb2G2adKMkmwK1HJO9HAOiR8rJi9fDPphBR4Imv8GY2V+DN
PHwm036Dg+ACOcJ28dkhZ94sjS3coCZQqnt4nooc5KlYjwlPzV66QpI1qJul
60TPm35GKx0O0OoLZUiCOLHepGVF6tIV9emVeH0VJLAjtEt9MaysgRSTpXNP
E/F5o2Bo8KZTNw1gDsPuJSjAg5cqW+7fdyMi5zulocqVcFLQElyjvxsIeZ+H
G++b9O8XnXRN5Vw+Y1oBeuQvpmPZ5gvPT/YmX/UpllygsjQK1kZGUi6AouAO
doiiaSMc6uJlsSV+PLLpWiKykABECUfwEVCDHl2tg+7ULI5O5F9//eoLg/ut
f9EP2BSq7zjuzq1lVGBJnkTUgGkrSwyfvR225gIzdj0oID5hPOqPvrKvckjE
xBLKl4YQy1HgwfsEOE2ABvwxVLs7LR5Y0Egp04u85uR+PRffmSV5RKzVZSlY
6FSxOteq9rXvzJPQox5VIGwXL0cR3t7FSl8LbcxZoRiQeRzT+/azkaV9E/15
pRAUGvcb/sSVhc6i6GGaMLAXVHmCLrC4YM4VYXwTwxDsrkYgotaKPEaN4DHY
Cl6Lx12L2McQJhcaHn3jT0MGDF0UoIEq742qS38r2oRRnIuqMIYiwyZz7qZu
DrUcLcq5xwe7Awk8uJs/swDX052fEcYTgw1HUnEdS47yOl6u/Ddcmqir0gU7
t1HFjhWUutkA6fFBDz8DGaQz4L+gevpBnsMwr82Oj6+PKUOHgJJ+azRIvYoH
jWSb+dOsAh6nMUfYBMwVArNjfIjxtx7fhc7iBR4g+Zd2tnh75Csk+pWCRLu/
Uvuf/aIefXIVV998SQ2mF9Sh1Od3j7mlhuEjydHL5t3KNDVF9saBDDoPtLtW
KyvoHH2CCiwNEW0oSbHn6bVAXHTFv250ppsmYSyldJmxw/GZq4r7tj69JELG
h/ou0KjE5O5Ryy14RCzTlQVzP8IkuzRK/ty/oqNXuceqDuCMf30S/hIX/S1l
xzaId8cT/0KOV5wI5/5q1XqYImsQd1224QQBC8UerqfAkuAZPFXNXNQ6onAM
QhIB0tZFo2yabi4nHiHJHtHgDd0XdlRv2p8ofiu3p56S6+PVD3OB3m5cCvSf
BPfJH9wDmrylJxN6PnygPzA1mBtlVqRzZPL7aNGxHxNu2su5yNPU9IuBJQqB
DeCpaQM9Z8SK6DY4tKcL7jw1Bakflo331ps0NjB90/bnJyTPMoedPoEIQ7hu
F4bPIvLwHl+1scTw0dJHm5P0c7Ihl1/CkdDlTLJdODqgRWoAYca0O68b70Yq
JJyDHgHpFlMNr33DMkor9bpDAOFQ5pR2i/bdF8VtnnNcF+C1+LBm0Ex2dXPv
mVHhbflCako5Xc7EOFeQz8/UL0seR+MVRAOlt5FoA2F5LRss/sLQ+h8n7fPl
N3rapQlGuPTBw/CI2prPFrPNC3tW6UjaKW9USv4MuQXJhv5rx9R0W8D6oRuF
qQ/qepkxfFM862zGIno+VhvXYmn3J8obt8G/SweNhrXV8huvzFHQnIyXEPwu
HeYBQBdYo0F6LjnNzy+d8tiDYhqucsP7Q8nWQpqjhjcBKSD9heZkXZfhUGlf
Wf/4XJ2NZSXgq3qjBtuF27JeUunQ/YfsfV/C+V03BkriqRIsChM9oSC6NVFL
cRTIo+v9fazB4+LfXDdwcPtn2q3B7tmVAPQB3J3WfauGgSX4dpEdS1MLqYMM
ysckpLYVeTCEY6HP2tNGUu0PDJqLabjHWkmNgEak4/gbpYSzDwK2xEGb9FR4
oO4ElqtiNqYHDKIu7tp0+x4CZw/ysnk5mKd2VhNKggha3ZHR3B9jCMYC079E
3IrW/yajaCPOsl4k8JuTHbbyMaLmLey2ertLM+ssBHeltsqKbG1VGIgRj5Ok
8RpSt5uDTSdIwdWIqVdKTUxFfBXIwab0B1KCD2WstH+V7iNwv32tY+uZgtQr
1ALhCAB2qXkGBwhCmANM18JBBRpaoAPaYzBj9mzYdgI3DqPSiRJAoin3Z9sD
1TQYZd/kzafhn+QLtiiTPO+TutLSSydJuapd9akMdYGkU0NN8/241CTXdJsa
0i9uMUyDeUeHoMjsIZe/Y1phNSTUPyZHOUYX7j57vWBU18Acw8X8DFazYQ3r
KsREog7kYYy1Gqh7CsxmeUdpFAmnYaJC75Ww9kVAuwQKEe/9W8q5LtorvnlD
ka9KjW3EoEcm35RRDdeRGfyRBTZmpATwhw/EXpsQQR0nfh5nNVQ0SWXONb30
Zrlg2HIpMX/esfVcEMBsMfqOIwYg/JSVNmOvjl0bJtVHikmm1AEh5CH4k5t5
YszqmNWXJoQsdjdv4ALGNwfrQUSbxvWvRW3lLe0r9d7pViB9/QniZu8NJ8aO
+SYQ1ssw4rCW9q17Kx2/4UCzSM0OwfsCo8+ANusXEDia18RYo2n8aVPgF/ra
L3r/rHNwMzuYfI5gXe/t2ZUlQJyHp5Rw6AuRO+UpNDMT3ghG+3YEqgoxA9dW
he3gBw5FaP+EZLB2L+j2PwSoaRKFwMHH/Mw/nXgQ6Zp++/9aGMSf2lZaRrNo
0r7llAz0q2vmJooYR0HAbZuoIywDuTiNo/akzKhEpiZsH3Loe3ojbhqSVvjd
fb0CAdhqJI9LsbogimujFc6q9EbGCMuDxpJrD49fqA04R3cbyI85yj4ayGAJ
pwtwZ+zevnc8LFETrY5lTOF4B5IxXRP8Wri9Hh4aF7CcjsNb+NRyh9RKA4SM
I82EkAHQw/dcwKbQrKiojq1R6Xt4T3+Hiua1r/jQ3fa59CMBo+EeiFvW4OLC
WWTYdzwiHW3oUUH9lCF4b7XNwL2SpxnsHyGSwWbIA7KyIPPTJe+Nhz/JZ+1N
mMePXbGochSgpP9qgcH90IW5CY0uHiXdrCeaObeIkzaJ1zkqi8B0nJ/19OQX
3jLw8Hoq966pjgKTGb2VsYMtQ8guCbvmbQW9/AWATZfnQhz/e425kLdPOqPW
cxhaUtktLCDr0BL+2azsmx/7qXJ+TKsvPnHBkI+5nsrfiU7IVhm4vfMK0F1R
FmOBmvrD2OtKGFherFiPQJBgKZeOdu9/03NVXIJvoNP7wJZml1I9sHggFafR
5/9g9JhKdaiac03buthsNMvNZfpxI2bshPtTlTbxLeZpunishYnk3qDT6pF7
DifwrowvJYBCGQaYitX2MsqLd7Sj2tLBc8UajiZkDr98/yPgy+NTnnweVUl7
bDuFerSEYYVo4yWkBG2maXg0KSic9eus9d/5GWSxhzPbKnX6hkaex34MncJm
B2797+6EFoUIRw9G783mlTsNuZmbL/FgJ5+huXdnb44BNVwruJIsk3967z+n
cgdLyhsEV7Q7HtsU5SlfZ9vMViyxw1p/hbUTvw3pA614XO+mSxKp+ByBe0mK
feGCtvOxb2og20nOwzu1pjfHZSZcaAcTDmzhebAFwnpPObpB9pdw8Wpetmsy
ztW5jVaWjva4RnA+1Ux3Eat9pUa8J5PuO99VGuTAaFl67qatq2Gyf71IzxDR
QsNWQruKoJx8YHL/t9P21kU/eVnrHDpYWQBfhvB7VtSb+Xj7sy4D7UmdhWvc
idSF0N1eWn07v6B5MCAJaX4dT7anIePTrwuCHmq7N+9CIWjVg79l0vx82Ea2
Be5wsaC8htw9ezGDrP7vA+Pos/BTRlytjmi2v766Z22OUgOIKKfaVjdD8pIY
GALT0hhXlKJtRPB0/MVfSRlCMYfRB58T7MbChletxVTrx1r7l7YxbTPOdg7l
YhSv8d0VYXumSVfsgLFpVyjc0sWx/WYCYPvYvAeTMkrDp1otK2FAbdeseQkI
7VK+aO1zS62tSpDEzgowYLziKrXoZB1N3D/jbRxGqCsATlhcLw8h19Jc6MRg
PZcgHCRCMSjRypcxIrF2MFKRZdzCTZ30kbe4FtHIFdAzpg/k/fqTKqGyOmb+
+L+8XYlT1uf1duPfTPZwUuZidmatBmjiPJUQuyg5DmToEzoS3+GiXp+qi40U
aiWK8BSxpdgh5gzzD6+fCaGLqcuhdmVdjUI5N7PYCicKgSUVUNu8kvREggXn
ZG+bSjrqz7MwyfuNMRBTQDsQagBSIMUZCf0k9MoijLt3U5/q4S/qsTjp+fEm
xbIySuAd3jvkvT0YkCPBWlpLJpuuoA4vF89Y4Pq5Xwy/jGIBQuVyz8zoYaii
GMngIyUQrYam6iQsbT9tCSWImA7GK509vPaDkFXCCYJpUbskmurJMi2E23vD
fB+kgcpNYTVk/VPCtJ5SOhFIn9Nb8K2aarnOoQE0PpIm3yxiFJ3zr9IhfFa2
kM0W++7Q8vrabpaUNlcoCNKg4y44bDegU8kCTQcaVwCkduecWPug0IOB65WI
jmUMYn36pKlxeGswsh//wRa9Uh/ydjK2gy74msZlCpG80gAUG4IOZJxCPbQs
/Es4fJvwQIILoqd67caPZQjqOZsF1Yr4z8vxwKfjz2C1uXNO9gDX6ftt4xrv
w8FrEENXwLy3EbEGVbqaWYTVA+QZhHSWFK6WUh6xhjmuKxu/5WnTO3URWtzS
0VnYdjyrOGEJk8nv+vAqUVIQ31T1RxgKpDVC6QB+grqdviKHx94c2LNcj9Sa
sVzwN5ji2bWPOPoc0f3sbzbey/X7InKoSsn5YNgEw2PS5rRvQWiU3NFGq9En
4gMCGq97vSbNLIW1eA4eyrdpI7B7LHA7ASxGuln23blJb/v6bYIlg2gxBwAF
x2GPspoD8nEBwsvlDvNOUIyfRGYMhkA7qZGtoK4Oqtjakiu0s1rXYg13+H8c
ZYnHSzod/B06eiYOTXPfVxe0+q9nrvl8bVswV+MFGK6lvlkCFEXSe6XjLk9I
+WKRRftuCLheF4H6Q2KqUhUPCrOOpbt6PWybrBdTR9ZmaSi7caBasyAiDV7X
M56UVORJ4YwwhJf/DZUZB9wdntUjRzAQCX8h5jtQ3GvLIoW24ovByEaDo/cB
XUFzfZTUJqvnkOFQE+orIwj8CYfNlm2+taAP55SpeNQeDLGg963FkgcQ/9pT
6k1pem39qbXjG7zMZCQM9Dhx4GsDSc4vsR90rETJCrW5xxftee2Jw+USyLWv
Lue8KWSmW/UP+hiREdfkjfmfBnALN+3zTBwCR5ZpKOdWBKlq8olKLseZOI98
OeBiyfgRuGiv781I8VI/B0d8cztU9R2A0k8KI3GkIOISHabo9/P8EZfen/N3
cIhIS33msjqbCImHKNEcGD7Ab/+YmdslQdrTHL/yRKnR7tZRnwM+aD7bOl5n
HLsBvUVug0d3oK9AsTlukLWofqkHu2fmZ1LilS4bLOev/8o1uPV3F9lSH/mE
3z6EDICVtEMeZ9Qccd6gYFLAVvI96VeHzCGhhRrG7y0X7I6Nf/tALbiQLe0H
BHG/i1wBtHdygMOWcQmPAK6j72kZVi5PXRQ26SPk5fVhYubZj9ynV8mQYt/z
Nl1PrzaPxIKsDE6LoAS2wbXTWLsYR40O3cf0rMRWTa119jFa/GorURM4H7+k
+Pg+HrnjRYPbPb81BNXMv86Yn+AcPA3L96KVxW6ApTsRnzCu7YEfJ1XG1Wy6
TZ+CpuzKRb/TIVfv2wcl64g/hlZCOZMfkAaJ6X1RZ/pVANUQ8g6HMx0rztlU
/+UFP431IoCD3TZR+JoBIzwpXr1JRoQpAXgJ4DTxJLxHKyHLOEVL+HXMhw6f
Me2o6SjI6+okOM2qpNA0QbUmWN8t7wpFtmSWZtBNqhZRB9baWR2hCpa/aykb
kP85S88rxV5/N4iZf/AQSNp1sHFji68rkFpPOjCyQAXzrpBVwnBjkUNWBect
3q5/nJHTwPz355IhKnn2rV0bFKdCJlp+AIsZnXXkqJfH2cvDYzg1yae+/Wb3
3VqUNAvuylVy42HcVlSCLDoqhdw2kjf/9Q/HC02cskVpXtydkRlY7yJu8uFP
Qlu2rmAGT16WfE/tJKot2M7AyXeuPA4mgam1d0fSpxNhnxXeplYbGbfcIxWu
+yW59KouJTtjPzNTomKQm9B8jKuFVkn9YFuaFAJDza391+0pAE1Om6oAJPGV
xW8cFKZPe+/xIRvtltW7YNZpaOET74jXiv40h/UDn0ytRwddmS6jnrjTs5eZ
W9xNcvpocJATJszNjqfLT1wAH61yy1xOPWwNfAAcO4e1+vrWXyqjvwNamMKX
j15dlJhdqMnK17s/CM7dlEt0LantZx6gbSXrq0uxB0zo1kVxES3+1p8RzkPL
JH9+4NIC4I4HEZRWoQ+7hGKXqQ3hP8FIcE9h+9ZMMRWTIMSazL9pEmX2lqst
5tGurOqkbtlvTWpQ9raixWFCDzD0KCgS4JZwYYR5tqG6YTIhrcp38/xcpb4h
Y350c9PHsaxih+xXvJQ1v0cl7TRZU2lAYch484JoUq7VLCmqVJ9A+U7elOoI
bqqf13P1qLoBaO6iYPLIQFrhHNMt6+m2moJIMDmCL+/oYd8ILMnr2OWcigub
hvfdTD+lBGI7hH9ucUOaFJVBMekrt8T8z1lpRKcuxYP+0qI+/qQtl11XmXG/
4pTfNt2HiiYzlTtrbUy2JyvT4/8WLi9JwcZZsOmD6Ix+r45G8G+ofspi7nsa
2aKINXmtXf/AEVVit8Hnfogz9ncV8DCbhp4ZmclSyIuPjgdOcdIWrZeY/dO3
VRQVm5Inmn3iJEUQKNjCY78IUqJNxzJPfO9jN2qksEHvZgxlOI4WUqOcFIfX
taGiQtzXabVwtTgaKzJLqPcctTziGBNuq4o3jD49OuP6fctpVYCyQhiIoj+9
aT+COxbKGIvOfOQYMfpUxF8sK9T1uOUygRdH5q42pQN92ke3WB1nkTCyd+0N
zNxUNE4xrvboSMadGU9HMZtx+6en9qK9OrBi0eX5ZX2M35XrJj9cE/mGssSh
KNryDyMPwSay62KUNJYW+2c52d6F3KC0LelJtTRMUBOpPmAljLevL2c/nLtH
0jM92J/lrLGrrZTw6pKU2ntZ6XI8c9K9BPIad9vrFg8OZSa9RRHFKQOJWsj7
eO1Bd8JdJ9tRGfqMFQAzcpZvbhe2y/W05/jFXImYaSaal8//RGpQiPB1IIx0
7dClA0up+HOFgDRBXxlvHYORSeQXncKCQ/M2BKLcVxLQXyuH5xm0DV04hSF9
FgJ0z5oKF+o3/NGDRbsUSDV2oXvQG+oM0wwKtC14zn9T856EZLEd98Lc5tvA
aLNvvxgS856v5M5fue6vBkX8m5tBXmxdK9EvuWYiB2lIgFpW1I0VzdZvi1fK
bph97RO4DstYQR1HVOl7sU/cODe3O53aaYNJ9h9NC+kwYDavWLAVC1sbeMx6
d9n4I9/Z/1fWFfUw1xy79L90RlOGk6t74CDvigkTLfnnPCqiq0Tl2Z/EzfwD
b7cQoze69d5PigqxZlDt5dvCrSoO9p6/pJCSLbgkbTX2KNiPwermYoCtCnzm
v3f6pRlVEEtN0BnD2VAf5K6mMZJhntLx6uWaJeJ/7cQNZi/KFQQvu6JDA/3d
c9EDaJjbX2Ik63+hWpM7BBI6EmZ1oA3VIAjt3Jonmg4ydq8VUzWdUk2FdoZc
y+YJF0fbrI3bbyCpFTj8+bAfwlv+iVpU0FelewfdXUMuMX5dlLRIXIK4SuJn
IGhtAbQiiFyAGPLAHTlfbBWkVcx0YxoNT+by9E/ABuLuVxDXrQ9d9uUm1dMF
AERfM5C4KRS4DWfGiJBqSWZMfK0PxsLHURFTLIyFU5luUOdHLkQoA2fEGIzN
sN38orYbpXGtPVqHSl2aC7XFd7ZXHgwrKNBLMzDyTLv5YXYSfWBlH4KBoOFH
ciltTGhjNPOCSYmFe14JSJ4gPYw4pQG3p8ASsg3jiaLU8ZKZZ7o4gYRWtHb0
qEFYYqSHf83nVdjbR5w8wYwyQ0gQ2mxdPdp3GG2QU4WTxq5rTtIu++JG4REW
y4aclGlTm2NoI379yfPF6hxtCXY0urWdLuEWBfyHGJqaO8gFv/NeIdBcgVS9
tpLi55Bmm/qmLn120NH+8yjR3sZaYSHpfGOsed97eiV6AKkb0knEJmGwkWbo
nkVokvXsZeWIqv6Rz0/B6bM80BTAW/3q0QG5vFvzuKPHg+Z9i70PPNYhIqej
kAXQo5mf8AXir44wnkA2npLaokNfh5UEgn7By6pi2zjR9ISyhyXiAQcLtC7a
sE/fMqITTkIO7k+KJDMDuJrCrahXw1armQNbb5zOEQKgeHB9HSZjwqh9x3sr
2dlpOj5I2ua9d9kyWifslaefuB4iiJJSgcGMZaXgZFbdEnlxn4mRAfHu2cPM
uYWMlf4l2qjyE1H+nFINp6zeQEBnrUR8dVXRye5BnjWUHFSYAvjYnGut3J5R
RVaG3vs0yQmBE5L8ZUC3CU+5/NPK8GlKNxd+dp4lygCkstd/hS6yg1Cpkm7/
D4c4QY2nd8kJ8to1vElCy7oGj9pGx+bsZPMO6iQYe/B4td5osi3QpSlOApLl
vW1hn0zhxh/95d4SnEL61un45Iuozm159ERJhmJGp5y2Mq5lUcr8Hqd6PgOY
qNYJVfbsg/Zy64tgRMjOyhXli6+r9mPCHP2GiGDUlY/7nM6UeUJhfk236uXm
gzbxdfb1fTrrOqI0VovjMgPwHxnioG7BLcWYE9YimZ7M8lo6CWblwkyCofLM
Az8J0aogOjevkErXXBeBM1y+Ng3vX9VtfSgNcTBAYg8eftIC810AxAV36NDX
QJsvrVSG+Sw01tzi12oFj0yfvAP31I0HhectGT2gaPzY/tdGuxm1dCUM0KtF
16UCJGl2frK9TzghCVMdgBPObDjFZBkD7F73PqdzO8R9E9oKmzRnHYYJ79Hg
UKVlwSB02Ebt39DTekX7afBP5U5TxMiX5Z1RpOC8rsBqSdWBJP22jGMviFKQ
lU+VgyD3XPdCr8gWfI8W0Ts4AodKlnct0CWFq7hgbCvRw2uHcBBrL72JyqY5
qnjlhpxKE2wX7bKQaVYt28Aa7vMQllH22ibbjJYKMQkWhiROItwdthXCYi7Y
fXZtNWTQt7EgZn0vxrb8UkMzdkV123LJbR2k5PT+IkGu07o586L/ZKP30G4Z
KPGCitoGHnQKz8rIsMrWTpCEL/MIvvawIcdX3pVzs6wQlyEmkbLcqLC8xIlG
QQHYTGnqudKQHdJvIqWVpPoV5wB9AToKeBEG49qwt3ihKv6AfVNoBhDWK0EC
c7PMpvAb8Eef+x72DdDp5pBfKJf+hErI4XzDzrp7PGfTqtUtsHaI0F2H9CoP
iCANcIAspviAurP+pHJTjeixIhQ6K9u8zsoGzqEdjAhOU6g61AtsxQPR2QaT
SZQ2SLLwtsitOFORr0jj7wrCBOlYJZyAN6oxukz3bhCQZ39MhFrv5KzVGAPk
M8XaJiqcH7PS+XrNRFGwgqu3No2cM2sn33uGWhNSb6y2I85ad01fdUjR0Lib
NIDaMcpn9T/fX+I5mnmuf11uSBLJFu6ZpFbUNXpsR5EaZdy63iR2JTsHtlZA
XGcD6zKek7AefNq9QD3vv2pRg+iI5CPncCea8iN+tvf2ILzFr1+w1xwD+pyC
19eOMPQAdDm0eyDz7m0sooEyV0dSLhpnXhjs9fmTecBovDLgGVqrKPUHzm+K
P5CS5yiRD8M5jF8vd9Udq3Qmzbaru/sQ/IEJImjCFvrAHbh2r7e/NkIIqUaN
tzlxEfeovxPQTTZuEwxCFTl5lbAfTLhQRB+5Ow+rvDCiINA7+FIGMiUeCBjD
/YoawVvQAh477e/KbamjsKBjMoLbk25YBjT1NUsi1Nt5k+L13mcgKMlF86Np
eHa7q6MOrkicwylqfvOcksZSCxIjs4aCZR4RIwxek/AHvvWqoq1vQAxi6T7F
5zwm2Ji6CVhSso9afG531WEcU4q857SJ0LeOz76RPlnSp3a94nJCQ8m2E7MW
Jqxvi3O9axZPAHbcct6U+OYaBqAHPOgF+PqhetQqsO4awddQott5zxn2CvdY
4TRo39msyhGV9YoIfjUjAV+vTdX9jgOleOrzQR0rl7G8QzW7D9p/XzgQ5dky
4gs07Cg8O+2BXq6jDBVYgnzVhTOb04XeyBjJAFXrX98jsHH6EEhiw5PUiewf
YfS+9ZTnImfoKICHi8a0W3lXE3KkTAna6eJi7ndGyg8VpNbtUFSTQqRgp0Z6
JasQdnhN30/aLT3fd3g77eVQ9LQ4O6e+23VR1CXSIQUs2n6Gugf0Yur4z83C
fK15vSeP4w7R9lh2HYV2E9b2NUVurqIqyBd3d6SQDv7rh4M8FDWIj1sRwhx5
eeflJ1Gy1dOtpoZ1imc2BmHssrWiUyMTYQ5zWsETqOJBMPoy47ZrfCuwYYGV
bpMv7dQdalzhs8PzqRDTASRy2LThbEaVGRj2gyKZKzOjZPk56O9XjnHhr91c
R8Kc4DwcujBayh9B8p4PZgapsTZHDKmAKApnBB9oNs6MXCRzWxWxRJ2cX2wT
aP2QC1LHt+W9mFMe9NvzJM2r2RufMwbUHe3dKSnPeeCoO9DiKii8U5eCkl9z
KIjx5j4yg7BMH+XklwWk/O3BXYHbcEhlyKk1Hg6Dvy0PqA/P0d4m+GIoD8Zl
byLHlRlok6f75uVSgxROGTZVBdSG7L7sfXVxp9n4Q7dskTLmmyrymy1zRHFB
fcr3u5XzYsyOCqzIx5LGvYGiQF7PqnwRbZHmJ4JJ2L9gEGdaQq8nWiEGL86c
LBM9AsIrrRhqrEGO4QRQmyC59H3PkIFPi7i8VaoUOOrbmuomB3+sq+H/mB6q
dEB87UODJBxuvJnnSscfCaWp/ZbqltR2Er1jK/Noo0ifYDcfy0mzZXlyTRf/
lfmMDouIPnpr1uoroFJ22z8zXZTYrniZXfXGEQ18ydtMuCQUsiAuaqEl+2yi
GeEI0sNcKMtlzNJo/CMTm1GYX44WZLgFrw17cinlRqfRLEGEsU4vHfM07gLl
FEV3BXgnzvu4xN8t2EVhWkcL1brVqX83Sxj5bW+NKzDE2JjMO7lwcesTVlOb
DQkWuWSObdVBi8hGOZmmN9oLJ9BmBr+UCsG8e4M6HHD5DNOoAhyPoSOq5s3J
/ChB2QbLA+9ItFnJoBtv9UpfG8km5vEDgSlIzNRRcTsm1FoLL6e/27+ffQI2
+JzyQD6v5CKMqy/IOyDXz+plPu7Py5uVoY/mZ9HNqJkmSCmpZ1Sft5ZVVQRG
t8sFZkL6YJCBJbqy9642wM6CRQwcDpaEcnd/dWLtx1nJgTPHg9R4fj9jTI62
7jTOJNhQvdbf9HWc83dgTdKPEqZuo/aSxQE945aP29mklIWDKjsNxB+Rcqgi
yQCSpDyACdQ3o/IhvpINHo2OEYZhWePa87ouNWIuUDXryBDRtJD6T2txQ8hN
/ncDADpExGcEbjRmsibjXeOZkDpCbQG7EA3CUksmfrt31uZI/+oYJ+PB7nXX
aEz97/9JPHzDQdmRoTsO4IGMizYJzeNZoQpuf49qde+tEBRkeD/NMytft8M7
PhTMRelxd296E1Wuvezj4RMssXx82tpF+Ii5SUuPu3v3Mcyyz0ByFW7qkF3b
hGTYsKt1XDN/XTmJLoIWPwHpfpmrJfBlWPttIsnBIKjNL5e1sdADxxkC0VIT
ZP4IcR1dRISJ+eZoXSYS5sOljQcBc8Iy2wxDfJMDwoHrhbhFXrp+NTojANaL
eyVupbnh299h9kyY6XT5OJiwViev419pfrD3yVAHc5WU4uTknx35WD3jzOyf
WM62ysBGL1Pr+WlDrNyMnW9uYUhH6IiB3uqQkeQ99xXxQ038gUlhQuxPIVM+
/e4vtMTzfnWqGJ76tSi1p6G5YnSWPylc6zX8pBCoky8DfD8kbt9DCSgdhARv
2AKRDTou/WKhDw8GVtln6WSOwLmwx5x8nloZ923isbf226JZnNS4+b3WrF1q
w9i69gEhCWlcnsexxcgNqR8r0Dxzt6LlARR5nYnubTUOuLvT5qtmMvm0refs
MJN02Jyc4AAkAw14NluT/zJC/DUNgGq/oOzSrtxP8NObgt1kJuEHI6EXLZRp
nW/kv53dGZCuX8ky7qSbSacAIUVXDTOn9QTZA8+V3O5sRDtrJL9WJWqxdQQF
yxlOyhR1cMTmPhWHs+d9Uzfkc2VDnw9J1nlN4CYnu6RIl3L8ZjOvWjO3w7ep
arSLb5jxt13/6A4jRsl8SZ+Ohv3P1b7rnIYoij2X7NjbNTgJIvd+c5mYDsJ/
6SUiYx7P5ncDXTUwbva1TLKpVFG6Aq3n8/3GSGeLPPb+EdjbQ/JS9x8fMnWU
b6anQ3D8EZb81VxfCQ7peOLINfFP7JL2kG32VNsz0QJ8934BFwjGZ5Cc0lkE
sPSLE3XXDl6SOA/elKMGIuVoZcdbA8drfqhZaV0y9WSkbkoQF5HaiHjdFgw+
X48N8YuKWkCWXl362gYaYCzDBgDdqzNuoVJ8aY/1yugyOtUvY4baPxYApCSu
tZGJCDhr5UuaCrcDWDLZvycNL8gka7w1L9UHcAPH1vhILubvORhpl6Grs8vL
eqHo9e/bwCvSwTi10p1pU1IJ1CpjjTwUsiw3JrL2WtLXjttutYNCv37ZvM9l
gNyOiJ57XdUaNGnOi2IDIMwOBBYqyMazDv9G+Nb5I9GrIH2jIaUjkHdFbJrp
Va9me4MVTjAryMijb5ehqjS3V/WMJCiHwJpME2nWwBEM/mLu7wYdfQLuzpzB
cKW+VyAs/6gn4Z+6SLjqc1Y7+WilMGYQWw16jLdZ/KdXzm51cUEqG2HvspvW
3wawPFQB5yl/urG7x6Wy6yAKeejjFsKkjVLJtWHq2hlfNtZ2BBIV4PnVqyWC
PpzmZ5ybe7br2Oqfy9ubr8PnxKJ0QuQ+eDACLRSeEBz1CyGUeIx5r41Ae4hr
BE6WeTvaRilNPlUx/CngglgxeHAkY5apHQ/eFlBHaXGCkq2UYF0JKPgKUqQ3
RwF8Gu7ns0lcg+bnj59KG3J5RZOaNks12440MhWGYajBCNwTtTJbeYN2MCF6
eqEzvdxWM6XrOyfVzwfqp0b9KuTLcmIPbKnAkNHlPBYf2D1adbxd+5p+Mujf
HK4trl8oPEUzdwWTDkxfrh5orteWwoV4lBB5rmETiJzjQGZsHb62q8VZeaVc
kSexDu2KlO2R3UP1D0e0Y4Sp4am+6VFRLf0Exj+Z1aV3rL9gQ/EFlw+mVrWx
wm/PozSDY6ugCIwu58tp2u2KTyxWw/WRlfBck0ZUAFc7/z8Vd+JokR1uYGv2
6ACrR1qeVByTbVYnW3M2lVbX+69aIteMUukDTbrY38kn3aPhO2jIiuwCtbA2
kdrvIuvn9IltfpWTxOIhdbVN1rMZHfFx6qb6heo2KFxBIZchEHk1J2aUMK6g
fUTQ5PafxIrpeCo+A82Me0WYbV1pqEyHIy7or4SxDU/QVNEUyxvuo6G0Dmmt
8zgAiXZimAzS+X5HIGcQOxRCySun1pVv+Ton2BOgbCBjx11mJTwvaOSDWNmt
2i7vOpcvMsNLGElOadsLKJxc17Fw21VW/AN5yzCA+g6fohBqS/MQXlJwqTsg
t+fwWDLKLcCM8bLZIt5US3pXwsDAQnxZY0qg17UfblA43b2ytuJvREXXuwdq
kA8Gd0rOBPizLeG8mlu2VFgHvPiJ+XAhxKKhy4wUX9gAUM910pUyEuKkKpcG
xl1aWBzYDspaxZ9mTv1pZf/dj0spnnpRiHn+wlHrO0T3RMWt/nxYIFxYsk/w
mocn3qYZdVKZ0qusmZUFBX1r/iYyVa3uq2bhBeWoIvnoEHOFKcKmALcZuPtz
Ly+XO6cxjR0rFzjxtP3qQuuy8bSkB7QzoYKE+AzJC1tXs9V6TNTGclgt3UKs
l95wQw3npx87oCA8a9ngO+J0j0OfHg0bwp6uH3OkOsEyOewsB0lTPSZ/VgQm
i7/Xa6qNFWu52pf8pCokYHQ7lPN0TkcgXA2uILjYT/dDehLiE47/C91y9wVE
py3Ccr79gkmrYhpuruxpMRHKmGi39Ul48yCIEMojmv7BqXlkjcIXkAUbg9Fi
vVybaSAduVkKjaE8Onyy9AFXM/6rG0GadkZcG/LH1KIq2YZy4y3skjW8JNw1
fVVigeD1xmomrq4oASULBzsWm8p1PtQ0XCPv0P3QFaxc+hrZhdlIDTqxFpKk
C16rc5BYPjcZoHuHJCsppo/9i/mGljgbgbBq4sYXtR8cT31VuNmfzs2r7o1q
HWfzuI1cn3mWz/55UuX9kCx34Q8tgiFiOn60wUdzpxSpyDQqCenRqB7YefMx
e7Uni7h45fcRn8oS4TxOkkR6e8cUYmSR1WE3j80n9bvXKUW9szg508F8SN/J
wgHB+etWw/e8CMyD1kZQoGLZ2nnXTDyuEPh4so2Rr0KOyXzbROCsUrONFPiJ
bRkH2TEn+f7tHBmpO2+HwvDv+FU0QNgbl5ckwsF7pkshoNcvptPTaGETi7xk
VcMicLm4qnrXMm7EJFbCrLccZ+MXSbhGStD1vvUYoFph2xWNV0+uJTRkQvJM
sAQMORfBWSC91U28OsrP69RoCsJdyYdKyoQgZbalDtIDlyh2FP5oHUDeJM5V
blBTNbiD5lOTBzLLDPvD4p/iVnnlRIfhomOtQ3R2kwtgUAPPkz5fGiiCUTDr
+4JN2z+P7ADWZOeCEeMuYtz9j5S9gTw1Q4U4esBah21JS1bRMkDp65+dQ+p4
DYINmyZhxkfFL1QY4Bx9nJZz+rfXA4/z2IQO7jJ9O4Jz3TaLfFENKiLD26pm
cBrQEeEh8akikxj1+cHLhQ0aNFLK5s4y3+Y/2BBXZ0n0+HsNbQyLs1DEXmPn
uIEOwToozUPA8ZgO3YABFDwmDPsAsaGDK5g83JfuoWeMIa9Mo3zktDN2Jrib
V7C570DJGb9fE0XHNjBDh3YK1hlx74GQLLYhmQMNRyAxy2cbKe1iVYDmbsw4
WKoJiczg+SzHQS5kjnu74BFLFAwRdQhY383UCQ35DoagGhI+CtKIX45Z9QSK
wgvZcY3zM+yy7NN6sLbmjDxzyPsfbCE0wmX7wa84OPs/lDAK6uelXB2aMAUb
9zs9YSJJWrr1UG8IKAch5+Be+jvK3Ywn7XTqYAt5jvLzggo8ftdxJNSMK2Q4
hcN3cyiBHhXehJPfAqnNr+sZAvNQFvI9G9/nNyidokvFA0ZAfwnnBqLT07zJ
KLVKGo2ZM8JVCPhTJYSz2ymCf2ROXlXhpzD7bvC8woVNe77eg6ZXmYWuDuqX
qQ+PW6BF1X6F1roD03w4jHiizerZFCx0aRXqWu81YGZDIH14DDsJ1lh8iXFI
coZ/lnunURAmsZhJ1VYEw0Vs3LCn74J49LwpP46DwA+kPUYzZPpx4cVEmY5k
CjZixswq76c6az4KYZNxwGK4rJSRfBxbxe9dfz9j4rALwXjmrikdolNMF6K3
tGMi3RKoRJ/a08PQ5TCr+6Igko3AWZAP4xly/eAiRRNGL0j5z1BeX4Anejp+
3zp4AuXxWsrssfRn2HWuYV9N9KKW20CksbhXxmIjeAfwROrHBVFcltIb1vuK
DDTiMQ7xaBsKdn2uuMoY7ALVleXpGlivu7VNfDi7AELV4g2AvEouC16xH95H
qtHwXKz68/zFEqZq7KOGvkEoEnfWghWeNxjNmCz8x3guKMM2uWsF9WHdGhz3
qaarx4LrzI4sfnGJLalb7uxFe9iwHzGS2MOq+vlwP+dwpoDKG0sYsXfxppla
RFOmxdTuK8FjSX+ZPcXUGbmu4vg9etr9cEtqqElbmZlVmweY0XN9jBtmyDFr
680T+8KfnCSxzTszAxU7Bh0T36Z8Ddup1SO77Z5vCDLi8EXy92p6Q9dKyIws
59N9BvdpCENPV3aJKw4S9Y8u47xYNdVB3drpgduyfuJomMqNHP+aZo410oJn
EWz9KF21uApZj8iTWhInI9qCKPH115jbB5RWiUVTfQ3myKkChPOyY3YEaEWX
IAOFGjclMRzMRu/lXEPpMIJci4Vo2ZeE9ZYPhtVjTVIdqTo3gkIsWmE2PV5m
7WJ0pMmDB3ws42/v01PllGbt4V5iMmLyk9OnKxI6oP2ZVjiF+C6fipf14aSM
ZM6cnESC5wBZVfl0MhNBMrjVOQHwp+Lj0bvQ+LMM4alVts4wtqYtxdDCS0xP
3wLnx5fhcpO/p3q8uB/kxtEZGNorde/bqACNcAnsk1UW7q5sd4hxTXRM3HbT
GkL55si3civgETxA93w5ELVUcb0MH4S7BSKqAOF9VIVvqawsih37GoFs8lzz
IcD4uqU1gZvHJ7Xi0bYG9is1ZYTD3htnX7vUbd970W1RcLTyqhFFnd3LnWIg
4VFsVBzbegm90McLsYjAd+wQ+VdlxgeE7BZb/Lu3RpODkN/Rd3NUnt3Muut2
GHl+nO2/SEFDxCp1w6vJfQib9ktkZFhji8SgAEcO2kfU8/a6WM2nfX+jF82a
83sJO4SmE50scAk/iqRFtvq03QUPNeBvqlQa89AIb2gvRe3rTZRuOUPZUAwb
onjIw/GfmD7SaJ25kY+fBuUmTByZuVREf8oJ3+ns10ID16nQKheiBm2Gesb+
SgaHlMkUDlorr4paxyL8JfYxzxOGBI78IbcHkpTCfgYk3JwD1ogtQl2aln3e
sMWt0f1hNMD//NcsfWuUR+KbL1SMkxLGBGE4MMPDrdSUC48VYZ0vtYGSr3fD
a4zLqSgnxhglLT0lfSOlLiHMi+lZYforhF0ryqKtKrF2MTYZji3X6Kn0w6Uf
scMGGcg+CiW0xnroMzmgEcQsI7MWxh2ZaIo7lwCo4Lxj0f8ED5pbvaRvuzii
b8i+/RK2fzE67oolH6lainfHI7nkgldbUERozI4oXB++PxdtaafoPr/R/KIv
d/EIB6Y0d5uL4GSae5PK2aA0A6StriUaoMl1Nitb0WDsdGJ6jF1Du/c7+0w1
sFy78mTZLUh3JyOemk0aUEVRrt3n+9xLdYP1ASSlWasVagA/5s08QDVvI/D/
H1qqiq2RHvNoxkiJ4xsTaC2VG//RDyrh87YW5VZKgJP2fUqKOtlheX91/9sT
kqEQuFkVYPpBBgvms+tN7+mfT09xYv1hoq7OMqtROtwMf+uxubU89TqHfPi/
jAyUTutBTZmfUsMABQzcxjPMM37+5vyZ0XM+y9VHuHeLEaADgqIdfnCt+eAg
z1Hn3y7rapdX+rwxjWKjv43mULiorsUREMlA9D9HulmuedGnhyxBk3Hz1Rk0
H9vUikDlWLu3XfOACr56qnyU6fNzY9+sQTkYgISenrbv9RMBvb9Tx8DIwtMr
nK/25wDJYLMw6ObQGiXYP58wXl/KXIw2RxeEtaGxN6UQxByCZRsdcGXip2R7
HXZ7pEpY6vlC2mh9bf21tfMXTcB6aLpupaD8E30ZIdbF9FSl9lGONGVFDZNm
UDvw9T48GJjl8yT4iQezI+RIGAJdUL/0YCYmHJ/TAUy2o6aBxnEZWH+XxovU
9QQFHFj/pteR8wBUK+98dyvottIbrCk536/6+IGwj/Kse6KSZeVICKRBMgMK
4Ml/ScvZQTejpDWLRNmG1FNvzAhQPgi3OnIkAQg3nRrvIj8/40RNxhCPDZps
tbY96QNlYzzfM6S3xFJsByOWEg1GVLoM7aArwkdK8jaM0BaR/OZ7kSy1PuUs
VeV0ko1K94ofFKnhIIExr3KIiunAi2M3pN1Yd/OuTtLwYa54CAkCSHZCs6/I
fDjTHn9J+Cj5NacvQVf8QGY/4/9R0qJTfDeDa0dpuNZeuGFledqjLFtMU34C
k6zzhPUBUFUfsHkiR6ef6eFMHrPR8ircqbmwbGSVmg3hK9mYM9W4LFFJA+vf
K8vaSFNVFm3jsHIOhLUP60j3uhg7L4l8/BhZH1kJ0szgTplxLMUxj4mmiyDw
JQbzEwl02dddPX8GgDMLvekn9uHflBNn/N0b7SXhr7UOPCBtqZlI+HooErVF
MFt2CFoRV3q0L23pnA1b965Wc8+xtm8id9fCHTu5ifrA9xTj71HtM2JZVDBt
4+d4ObZDZtiWWACZEDfqzrpqy+ttZ0mF8IN24w8JTjegDWvg0xfKUj8stzJa
GdjrAGZ9YwNDMrGWSMjgMSxqJ49Zi014+kRqpHF0rnycWtg0/cBmgIzqgRKg
hVWt64xlzCqM+6e/MCCiDbiNmz7iWGMH1mKd45jYw1qS8Nr4AfM8ArYTJXP+
p+g77x1DHcMmxWImOcRGgbEwXKy3mGSxohB+FmcxKjAoWNdb8bYxSEWzwJvc
lsSvg6Fi7A+02MkzxtZMxPKIveugdkIncpiJ45dFud64s85VRbXeWFGZdRWa
XgUVfHz3z2I+y3Ewdi26SVHYxG5h6jpIudoaq9BukMRJ9fTb48BBubtxFYey
pftXTwhatPgqfgq4dS4i4Kj5VcchgA2XzMJaj3faP7oulMmKUr9xt+B8M0iY
20CHHzN/zKwF2styK83AHj1fhdMPRHaZCSh2J7IzVhMyFxhbueD61+KkQuBY
kcufdhIaqxSTqekd4PUVshCEUk1tnErCpGCiRs/f9y14Tj3R6MfO1tFE2bI7
wYrKNGnfND9tJUkZ7qfYylqToBC4jRguScsxrZRwwmVAeQt3lMZq2/9Qs8fT
3sMC41riouLP/sjyHtgKRG96p3hbcXRMCS50GgmysnVUlH1YaYVW4KXhiuc+
E8NMZH52Qu8h/AZYpXnKTyBylnRZKTMr8X7LxYrCcs9vtJQ7wVzTIufeCRAZ
nV3gYtmF9z5KKawOO9BRKl+9SVNZz5Jg4hMwFRIxSmEuY6vcPpgVtW36+5q7
3jrGnh2Jx06BIH79DWCtarndHxQXfKShmxa/NYncZx1m0aHqY8KFnnYfhfyv
6gsrJ9fejd57DX0Tnif5bgcQjftUoOtVDjUAfnCO2bR44or4ZvjvPjGJanxK
LYWFJYjBBorbRoBXf9cW5KZZ9pY9RhfcY+HRHZQQG4b8W4bm4Y+c4CPCLYHa
FBDMRO5vdPNC+v5cXy9VHJBai0EnjEM60Lf65S6blWoB51+D1jxT19UEh7PH
JaZsu9iarPvN9hgkCKYT42Rz2mi1nzqVnLQzT70YAJfeylwAEtWH4jCFdUUA
op8oQAJCe+Esur6PTSSIQtLhTWW+Ycosx7ScBehPT3n04rmeeqCO+jtvUCJb
S4a5jLoRoruAaHk6ROTAkAnAKWPtGELQqzifX7r4pGYhFeevOTVdCfYZTsq1
yXbzzFEpxsU0V5W1S8Ky1VLnqW5X57KC/jqlOyDIiIuXiHdbNfr/8wlXK2vn
iUGmQhrpDRdqkegrk0Phfo2mEo0CBX10U5WjJ62wSJ+JHvl1h5ARQ/rFiCUZ
ekeYvo4QRAHvG9jtzemSEB6eHKQ8DF6ihuHHyDg9IUO4R9mmUCm0t8O7f4Nw
asJoQ2+H00AD4G3mW8yfi7KxbxPl0ZXLV12o4dcBupMVy3MCh+S2KMCTZFbO
/6PFI8iNVbLUhQh0xmKMse8zE+CnrGN9aV5STFIYla0eE3YGiQCy0h+z9QxC
jB7o+HjUWz4/yeLGhwwCKsvj0Xkt7Uz5ogOCTmPhZ7g1M1fefI63igtjAhud
gNCSJMV5kSnPRTvg4+TmI9zXRwSoa2bKNjc3J/dLdcqAqW5eJSeRjFkEhpqz
HtNUCrIVUXHWqlC8j4yRNjUCaAiLOw5fMniuAhqfbK6oYGJ6SWBnRdP0KKWM
zQM1T04CTuhZnt8FKJSEiH88Qearb07OHoeYbFtsCGPD6IGt2GT2ABpNmdQY
Y+H5fZsOiGdbpWjMBh/XqiXKXc81YNbdd1quBzgTbPNFAS4OVSuKI7qTrA1F
10wTlVCqqcnFnrDvzdKJikMi52M4YRzC3Qt0jPiLcT691dS6+V6/wS955Sgk
iSrhocR+fu7dkv8j80PqxJ1QEqFkQdW2zPpTM0V2PWt1w/w9xs68fN36Cgxk
4dvL2yl002YwYwchox8XvamZIlvLy/N0pcImEV79h8bzrIZXngtAenviFAQ4
CgeIoPvQwHcQ62uX1YUIwUHCVeSGaAwdv3141zuQAYVXUGTQp2ffxx0sj0/e
wDh4TcW399e7YOsRktENpACTR0Od68xReXjztr8k+x39YAM/dBSQO3AJAD2f
8drEldUOYARiyfIHqduJecEYyRAEUnP8WiL9SaYjYvtr0ht6ORCx2AeVihT1
2gqd2UkVndx5ifx4EXfujHVchqJI/zngAXM9nAV3q+zrt/bktWyLxaAhCLL/
yQuWmuKILRKjeCqpnExxhI7xmaAGAWrKW5d9fS2Xw32T+onWKffR4l1Ewm5k
uh0nl+3q/jKWiNmLVYYEjcFlP13KR9GTYqAtpyKD3Ef9k96qIY+3h7nZMY8Y
PJYKHcwgVI/dppZSWvLdcbrgEpQftu+vBISSAk/L1RkRWVtO5DmxdtaPK9s0
m6VkQqbfXAnMBAPMZJLTS3n905Q1lvJns27OYdwHpyytGh8rFuvR4vjdq4yL
3vyKg2PWwU0HalvAdbJ7eQwq83NsqBBeZvvBUyBIJlooWDDCqr6nmj90+A90
krVgVWVhWBFb3roCh5HJGv0P6AH+bmxoPxAU9lQM2hJZNFKA7akKFOn+X5uk
x2FxPWjPrmq72RLw+ilnK/D7bSd3lumiKgDKTbuIUNHxqb/nFRs2NLPd9WW0
UIIG37UkNMf9zRcYPXO4+n4N1TRiLxaoTDXWTyEDYbOO42F4WomfCMLNj23m
S/OWBC+4gPIaVpBS6ghFGSXErxucqIgGcFV32IaUnMANdQS3WuACXsyafpTP
37WxkZHYXRwQaYnO8+kQ0L2zNcl9u9WCkwRxdoNCiX0SCZgxuhnLgL2dLOiS
aYaorMlqy/bcW35cD78ItaM2Q62RWMo/C/wTawfCiXEdHAW/4LpqNT9ClqSc
ZEXyQllF3xWIcOR01EsyivLo7/b/85cS+xmXAyNTvBdtFqHPPNgHHdwlmtkx
HW1wOJrkxdLnrLUsAr10L8GXiVeLFlZKXlW+QvdMx1QiHSjtzxssnvEAMZuy
dyQ1BvSi3tljW388PIHLB3reSjlVTPFVFRH8QQe3syzahc31mb9odZ4wZ7vo
qbWZrWz96oEuwNHYov3Eu40FxIe6SvH6wQcHoYlDEP/tNgnmKPwfp7bYinHG
ILqgyJ/EVjMPAS6XF/YkkXOV7g7mHT6GK4bSUXZb3lg1XRwxRBTV14ydlXYW
OMEnvyh+Qrtjkob+9D9gX4vGLDESXRxUSmFP3Wvwj/MzdYbadbjyhxDjKSLl
kkeottQsXY81yOqYC/zhq4aA3ZlqQA1n91aotPKxkgsCcRbLuL1j6hIjF5Lr
Owz7v7ZcLeghnkhe6gicGC9JU6V86olb++bQtsAeRWOh2o4EefIb1gw8C4Lv
W/7lZXN5PxapsBYy6BTk4LXOQdP2t+6QW72XUY1Etcxn36wpn7e69mvEnIRZ
Y48HTmc3oVEiRuGTgxl2M4g/mExiuhQn4gMwzjwPG8e78KP4EbpHW8grX7N+
YwWuIG8WYUpKNLYGZRwvYM8z0wRzDYkK9GLxmqqICW0nKPF9Zj88AmydQTGo
RNL5gkqE0bbFv8hAxXoTauPkELBOvg4f2Z0C6ZMn187HjTIMe7eNJOK5TVks
dIACW+sYhl36mslcpZpctjlKyDs0bfigqhUoNNvqknBaAPt/LUY6Sv2q2hIt
1Y85HXfXwbbLpKwCcCWujXZT1NtcEDxdmUdjHni+EsNwNUTUAwL1YyIJdCrJ
x77kvoJU+GomUbL1gYJwokbsvUDtpbmk6DtXddi17vSDCJcYojNR4JPEtJ/b
KgF444gJPhBAQmeaZn42xuw+yi8+MH2VDycRH3K+JHT0tEyk9Ui5zKrQAlwe
mKt74EaK6CC0UiqJC5vhGPA6/T8ycMUR0IT6VKKn2KzoAsX3qNPS2oQfMgBX
j1meCzUy3LslV7DnW6MtZrX04JCL/7Aep01mOkG8YXhZWqkkdQc4gqZ4OOWt
s41KU6IYBQ/6oYJ1IIuRxMKbmWQTx69OoXndgnc/LVizLsCZ6M/YzD31uu1u
emd914t6grumJdO46YYZlq9ogOyj4CbJ/0H9BENgxUAJcNX+9+mxepMqSd1c
bDKsIEPQvi5ubD28qCGBubxs1u+bqyYiEqV2/kH5NbC5D1sfcYKOSuUUmSRB
N1QHli0cxah+NgWhp9Bw4FQohX8p0OVJGvP7owXE/1pz1uLJjwJdmdCHTGKK
ORW2G5xCmXdijUOVbXFuvhFjJ8WgizNCn1HKuUuJj1U/St26CTuc7Vjn0oI2
9EfpzOsB3go03MIh34yfWKegHuLzTcK/uN3BH2KzOnR+3hUOOiJQhKoL1lNc
5hj3GllZSUP7jTgQP8RwyXPfj5dB8IaBm89YH+zTHiNBcPHwa2MSYXkVehJj
u/AdFDxtNUvmxMhlhxfb8YQEpqb2UybIieY1IUc/RLOwY01FFcT1VMUv9S8M
RTOTn6R/kXS8q/z3MFN7d/+nbDobyh91XwdGj7H2JXOJycdUh3+kOQ3MBKEC
neC5A+0JdfW9dOjeuvyklv+WxGynBEvxQ3pILlXd6D1hAKvAVDce8jxU8gcL
4C3VZd+59HtnNjtJzKX7xFHupw8AXGsk4P71IgxBd55jB+VF6RS5O2EZaXXN
xvzYgGZFqOtRE0xUc1GGr3/PJ6ByzeAugoYrO/yG3p7okrYQi9a0bLJf8Lty
0Fs60u4B2hKeKevs5BJP1r+1pfWzmyio8X31hPhF6mNt/FDIXkR3YWfyn4NB
iziZ+9eCdMUd0KjYSd33scZ6uRBR3i85ELSAtX1SASkHjrbZEydAUJnNxcVb
K9Tz9pInMHEVDHkmSXr5UxL5m6w1Mqj4UuCxKpaWMQ1Ygf0N2wJAv4h/9WJ4
cX/5tXi96K1WbDSOCMUoqnf0OAwutvaPfCJkUCKmp286cpPwX3baCAHKbNxC
hti2NyDalkl517tqmOtX6yrH+Zsxv90//QO6aIStex8Oh6X2YTNA6sJVeqKm
N8GLVQpHc6cBldWobEyewQo0/yNkN8z/ArnIT9FNsIiGndw8rSaKHLNm1fv4
AkdymMs31BbGCdElA+eom24isUJIQ9lESjk0KWAJVosCs29U+I5a7xd3Eatb
yn6ke7SMbt/RN57mYbDgTYQ1WhAGRhdxQn/Gs8PJb+vGG9w4sk6zmQoqBy0T
bl+FcAO8eDMxnz3peyxR94hrwMJgAk+F2218MMFpPiLoeIc73uBSlGQmy5+9
dNKAwRFn0Oq8iuUW5vdQgrFxoUco287P/0Q9Yo0NgeOIH5GdGW/JX+Ffyox+
W/EQfA/i8aa4sQ3uZ2pCHARX7JJvnLRtB22sFh8wT495m/O1PERduzpGnIgF
JQf3dker2+uk/CGaL47/BnRphi+tXbTXetDsCQ5txzPHChSplwbb7eqKpWim
BuvCDt1MERuui8/arpSCv3wyoJN2qZ1ehIfBIwkbVW5F2MFNazY2EUrQg6T9
jdtwhDbjvAadstnKpPJL8ogcgtWDH17C3hW/7MNpelmYfBG6MnUXQbr6FDQQ
I47ATjZmbcNcjeRJgfEwTLsPG6R+yCPK2pjq/YnbDVMKSqb9GQ5TxnTjf1Wf
COBq8vXqmgsF6BKH1dycb/CCwoYluiK271zJGgmgDsC553BJDKD+auYkc3k7
kfrqy8VAGwEqcCJVsL/YNYC9QkWVWP0KJssW3z8uZTXZFBBqj4ChjHFXGY20
di2+tvOVf6TCqi3IRx5NfoRqV845vPvydD3cuLYTMTe1MNuIP8a1FMe42z+Y
5InfxsPEGlJk02DGt9QlqUDYLxL/T7nNAy/iQwcyac/uisDY9EPPXBYSmO8h
r+8FxUlahbZBjVtvJ/hLm6WMYUljr0tWCfgJ2WOMqPa89gY869mnshL8VbuZ
9wEJR2VF4qpeiPiTlxnaJU9GAGGbuxuoZ/dgAvJ4W68J0WK7AJmG1SmGADfN
drCJQONbC9LTo7X+tLPkpYKCscP4xyqthO+IWyA8O4RdmtWuO5t5JUfWtFd8
VyxsTJjantwLazaFxdKoNhykV+0QRsr2VhyDS9qboFluidUCoVfXXIByGAJY
+y7ZmPYbQbWJlROUwZVWXxN0qoLGsK145x9wMNNYwt4y6stMtYmo0GvZrVP6
fQ2ekUdZtcTWg/HWbefJPg3DvP2ysFshWFrUoh7B9imattoNu5BBCbYdaY8i
BNV5gEWsGgXpd7OEc23WJ3/QCAK93MRYq0ujYjip7Bgn8BnwhRvSjXWCiZwZ
BVkrgD+gg3TISxJnVZ4t6nIaWtbBGCjMBVqU6hKG4jnCKqvwjUuB0tq4DotB
VETw/QrHJ9JTsozdlHVZ+dBli+Z+vgAiK6CiChiOcbRRUZL40OOTu/HVHJmP
FmAi4WfVh3tEDDiESAeCapjoMqkVRgZltsXR2yo/znIdNYYWXi3+zc5E7hGh
kdg1ZeOyRmheKLkmbkImPaSPblqMDw+ML3UarGyQoE6sAjdr4MB49ySHOGm8
qj5uzUj7VLNkunNUA+CI6JrQhblIVkH0zQcF11ATnzqfOjGj1Wyit6bOMg39
4bD/LVpCp927a/N4ZoI8bGgnJzCMyeDK4DBCvfTcPlYE+LmaSLBDYYmIwhBs
7iOwanII9cmbL0l4uuy8DukTNhyDACQ1iQhgjwRaLM3KfWeYrxJIjUx+9ksW
ejXqG9gIrjVsZyYENET5KKya9vApMfH4h6sfKdjVEJb4vXXvkvQnaA/2WdPa
8/GLhezndhijdTVnD63sEXzRq+q6xTMs2t5ve+dbK5VS36K/4sef1wo7JtMT
cQeLeLvt9VUkqSx4HQjptdvYB+NkEHPQ8ubAYgvZY8gqukwblskgHcQbgw4Y
oIc1PJ/amFOQ+pjTnGA9Ci9NjT8truLNgWI5zb83aEiqr/BvPxqVv2y7/jx+
Vb3c3oWOkDhu7UN8+QrS/6CD2J2fjF8/9rCODOPxv6h/iPogQDACktM6JPDw
ZqUi9wmrpx8wu+nUm+JZblFt+QqXw1yeKxFcmdXb1prQnYpumUy0ee93nS8c
RiWQHpl29hVKu2398Gi2kx2X6neyDLcYBC2LQA3ZQjVdFq2+3L1eY/CXK0t4
0BGKyACSgS9xa4CWeZloYB0JoD+/cNJV9nDSXZiu+xdtNbD97a/pK2+a56YE
MlvigV7DcPI0SweJorB5NIr6kj5nV7R+c4YGVEBv8eybXhi42gcmD7tHviBj
QFiWifFFf62uSoQstVR72c6ubSH3qZI9MzyvAHBTCfKXcP4zhs4w89Iu3/22
TpqjUdbBQZWk2OQJ8va184eRWLhr7Gd4Q0xnBK/3wvlL6k4v9xRhs2qq4rCQ
vy4rZIvRywtGseR1+p36Xko2xZQ/u2oCdOw2DmoOolTjDmhN6HnrlFLMzNVk
4OiBxLbR7ZLppi5IVnIMpMykuU+cxyTQVYcEA3LTuZ5wIqn1eKjLKqfWN95c
RZSH8cTuAWW9/lS0WaRfR61m/f6denYdI0rYMWL8EseAshIfCB/KvHRjO1ub
ofRykauUzbMT7MkWkdiSiW99mXm2SWdWVmayWaQqd7xTjUyR0hjSN61kzQfF
d951wvAvCgLwzZlPxsmCCASFmmmRPW/czHWWx3CIIscoSzup5yudiTfIjKqj
JoGTNnTVGlCcS+ojZhLMTM5mXpQO2umC0Ti2l952fwKg+S1bGrOS3c8MokuS
MAzcjFt4yzCDXvFQpxGvuG5teivuuAKP35JJqwIWHgpscZiBx9NxD5D4YgID
U5cBLjn0vmYfzX467wrlRUM4JbMB8QkK+C9v47x8/72x5F4qDWTbQ3OWqTEk
9piaz2DvTEqh+5XIfMso13ey2RvhoWLhkSnuCMm4rp3SLa94j8nbmJdgyqlf
cfQ3VjmWKt+8g9E2kF/3DtcvH/w5nm7jF9VxciYR1yVEykQ3x+zUwDL1ArXB
Nq9opxxaNta2ZOce5GLUW7uh2+IOgiLtTAin0F6fKrAOJr/tJicKNCS8ol2v
mKN2e4XZiuF7koec9x4GK/KaeIKwa0LNtGzo4d2lZlp5NRxTm+gSZjGOfZSF
5Fjbx2nzF8W+etwBEm/mNeaF5mo8seE0qVnmuqogclg7o6W1imjf6TXYq2qe
I/YUlLXSPIVbHf7JFUCofQGVB/kya37V52HLo2EBzzlnMGTx5IFqR3gAFsv7
KQxshm8ayZE4VNJced48ftktOAFQv/J9Y+KfWQeuQm4Ak18FRGUF3vt5D9yj
SxehEGR32xeAJCs4kqiL45zA+yWQHqBuX/TIkp0u5+xs0/rxYorHcpzSJZQF
eKuzPG1YSSlpRt5lIuwjG8Hs4wYGDxLgAK/uZHAlOIP/FYKgiXRUd3sbC9vf
Lt2Gsj1cZ3p8MmJYZ3ITlgo6WuOyxcCHLUjEAYkqvj4MBQNc8psS8Xo9G9Rn
I3xie4V0NgMch+c9M6MvqyiiwPMkb2gSA7gMZRXijMm9wBlYPRDnHQIrQi2W
u+8TFOQNr8+upzMPCZnxqjuPQPdDOr+ww3ie24974Jz4MU7r7UUBszHazSwm
0QjnT3iapatPNjMiyX1XYjkQKE0agM2aR4PhgJv8teobuteU0EhtprhITxJB
cf4n97OJtdOXTfngp4hRZbJqBkUfPor+pxsha5Ao6s6+7hiK5lfMdH/8yoiA
FrMe8WyNeTop/IuSqSWSVkiKurS/+VFrUyvVRCGriZjwriynAfa2e5lR3IW6
e9jsqMtRJWcUhcoP4tDcyE7bpj5+C38JGT88USXpLrB8dsg6ltjuP1UczGY6
u54zbEVIrEHYBS/YEwkIPnuCimZtdJf62u0G5CYu3KDs8/nKeYq8BPFRXsGP
sRpIVrM/nCbXK2tEllDN7iGU7KuP68EXBuIzN2k4uTueawxvXap7f+gtW5m6
J0EySQ4klriLdB3lpMDvaOsCXX3AUCFEmgEaZ8KnzOxM+Vy8goLi2XWMFjxb
dUvTVAKQq6iIqdTz0C6N+YEyKItM+ZPeeJJW7f9UAUvlyXgLTb0luuZo8GGd
5omaEj8bEmUWRk+22oS5ftmitXErr3SKkJuDep7WMBWz+NKjX4mJm9wZzStx
A6FS/zX51jWefbbYDAc1rElHp7425LW+ziL4a+35NFeLMtIYTzWuxTluovQf
1DYlu6uWeLArwf0oqSVGe/IAW46onXoNe6OWP45NdhqDli0NTbDznSYFxbR0
xaOitID6iBTlmkiD7Eg+xKUOlKCTHYLiCuZzrx17EeoYgVo6YZcvImyi5FY3
P5I8XuIxBlqYZVjYqoKOb7Y9UWit9QD+FbQsVODGx5E4YAI4i9ae692HlQJi
IHfzAjz5UV0kUw5adZ3O/ldMnHoVcfnr740Vn1UroCsZK/g2Fu5cuqDWTNzl
OXlNaJLFHMmaaOC6o0EvNQi640cDHj0xXxoojz8FEl6FNhIhV+gon4VBw4Xx
Mz6sdqO21RcIyzsdAEtigusk3ZlZKBbmHVXI9r9qS3c5E/KPi4hp6rbrPebU
pIkLze6p0RGnMp1i5g3j/IIKkRY1HPXtG/Y69hSgTZTaMQ0HgykNBaHgOxiE
AzmYKZKNk8hwXkRA5c7CJU9KfYG0jh00hV7TIEDGjBqdvwj7E/N9ZGtTpq3j
3Gu+K8Md9kGDu5gOARhHtVPgjzVp/Uv4488vAJa5lfiApOn0ganRGmsg97Vm
+nyfB9bxgnRRVx10jjiPYnJZIiGPum3Fo5WANr6s/CvvdSqqyDk5UeVcaivX
C/kTPCVqoteARueC0D8EVd+rO6JMQCgkA1inU7Ba9tN/pftDhvQuLU1wNNSd
aXYJW/oL/F924sZIaAkl11sXYDfXK3v4wFGB9mDTkL8PSsmDu/Sm8C+ZwPFx
exGag6z/KG0iu18o4rZ7Kf9gAwp831PsIaZXF8a6oJLLmTwKJw6qt9Qd6mff
A4Cfhix40FbZcWI8C3xQcGDXKNhAs6gAkrD3T5ptaefh3Ud/20lwpzi0TJ42
nxTZeokIggFGG2yoSTBTNjDlhcgOw26azuAAkcMNoAjVbW5moAp6D36RZq48
CuFRCnLtry3Cr3WwbPfMXPedxzbgyK+YZzINMTnVneXLv4U8D/xsUSQW4Q/6
LOtqV5Ybn77iLmio5ZRUgdQAbrKtSwSVV0zgu9DvU3QcbdV0VmBioUhgY+qh
N8BkXiXdUQtiDBqZMZsxN/FWc54rdoXOopPMwRByf6+Q5KEvkt8Wzkpm/LSc
URPMFUtWmqVS/WAPhv7YziWePacx3BEmml0AfE9O6mXWeGBahIemGUMmOPP6
nhD0OgyklIs+DUqJAzPhT1fEDnX01d6+eA3q8LhEFTjAbH+TpG++sGJvrbGK
97iAAjcuaC+FhFf/0f4bKlvZkkgU/AkWkl9/SWyYKY43lfmxhO/uZAemyc2j
cK/oFjyE14CDtmm9tSvs3rx1BwFEp+gAquY/JI981wnh94FkMvNK3X3N1fo1
tXw3ISVDTmvOrC74c9/wve/oe18zfK5v5IZTppZYKVczD702+E4CvLrNCSdW
2LQTbxFexRyIwL6EIEAlw1ApFg8fyKR07Zq4ML9fjiVMPCsOncAjuROy8aYi
KpLh5PduOE47JpJNufMLeoQV5l7lbvg/BeeMJD8Q8aIqSrKlxuLuGPyXPYmy
FmL4lC3s5jqwxt9+qTkVQQBSDbVGdQk/ZHiZrKqOUTqaBJqRJKFaCgBDG4l0
grSDlhHH/zvCA1f072flKTnERKSKjS3fy4eo91YLeCyC3egIpg0E7KxLJ/+2
xXmvNF75TWIxq0N3XOLJzXUiqXr519BurR4u1DSegg1HamUSPHL18zLYNaqn
VPGR5bkWVUhM/lYTI6fww4bWjFN0zC47HMV5qVeUgTIHhMlrpmvxinwATuYe
AdimWk1a0ZD+pcA+96rCQ3s95OngZUH+B1ne6tZ7nDO1GA2oxgLIGC7nCfm3
35bEPYQ9z4mCn8LD95Lt6dV2REKCallQOypAbbl0j8hSE5FW6uYrn92JVZ74
DGGEijvOzQepaaGD5d2zAxUyeTxQOOkXr6sB+FOYYDRryxKDFLAAMrg9gOyA
oQaKfyFuG7GeI/XujWkUK5PU8r/lUMloDg/ftmSfDWgUX5CYWeHlTHZELVGV
toEH/F8YA1Fw4vuqIGDmCUl2BSJyK540MWfvFDGrGFr3Gp9Zhs/wgI6GN7n+
RFQt5udubWePjFNVr4UqroTj2J73LitsCIqiR3BVDo3Wkt2CXWqSv2QidjVW
t+vvBNFHZOGSiUR1IjoxEcG0d3c/vfB9OC5RS3OyCVYQSU/Dat3Ydw19+A2N
XOY2vkeiOgBC5480v+UNlWaLHLQgfWzpeCMkKmaeXKumJAiUntQUjmCdlePK
cJTwvuqEcdug5B5TT+CMdGQ8XLQLzhAf+B+ZNp0lXV+RSoVkXfps1XnOwKsP
tX1GJycu651BpMpUXI64Ba1XqFEmHROV7TOtZcoF6COYf9t+E50kBJd7M3Q+
qOmKZaofHwtlgID8AM9mYOJGBKRADsK0HDbQAsLNGPI+6XLFiGFUFX0qaHjp
50TdQB1u6zFK5KTxyc1wcpVwsJOVxLSPTXe0LQ9YrfChNcyL+jkkkVhgOvaW
J03d2t1CfZZkA38iwctE9BcO7A6I1IKrEUN06r6DJ8jfyv9BMVAul/MiiyXA
DV7ygBKq3dTKF+gMIOxVBPsYWe8filzpZn+SQAvx63Sb2DTixVuhR6CkC8k6
PRpVdBzuoErvrAFNRlfsjZAL/oIFJDqnbxAGGLUgXQk38dDj4nm4NdlH11FX
JiT6ZIppH5Jxn72SvO0IEX/rGzuPn+SqNH7N2scS6Mslgf1kGkYX75vRXqgq
mhp1muhLUx0UhfvwFDj9X70IWHXCEvsd1PsWNq+ylOlDYmFnw3f2l1kP+S3E
077R+v8kdFyDeELDC7eCkTDVuOdUlQMu2NJ8/h6u8IIfAwik+IuWNHHAH+td
LWPaswdVkQLTxAq6VumWrzwP2eLdQb2ILgdYfTZNg7wsEdWrGJd89ek1Lt3I
iZ9OBTVlTWsngZMRmlYCM6MakWepJZK7qLJ1g8Gs1wtk/0KgE5thsU746Hu5
ZFqEYdpaNH6gfBGOrCoM0X/Vk23VvqCPkHp8mwhpquZO3eLP1HzxwGnn0r0U
oNNMVMy+31pt92AT8TNgz+i6uv140WfLZo6YW6vvZwU+OHItiJGeJZ/BMmSf
SMDinKypC5HMcmtSa91AQFx+4/Ry77KQU9CpHNo6apMeufKXF3/KclAMKf7u
bBvzaP3Fu4uyLh97m7aQ5IRra4jnLzQTAahmSifuhomA6Sf8ZI+BDGAySdQ9
5RzZE/T/XRILmOuJnfnh0llo/Ifp/oChz9WQ8OLSDfRuTBh9PoU52pH5UZzZ
kKwY+zk8tXXH/8i3ZAl7LVTN5Ey9p4mzp+z0NeRxl1mcymlLvwvryQDZn7g4
7B5a1nEqXpFr6GyWW18q9oQORb3jERfMMleedN9JDQIS1N2eOb7YqDavAh1M
I+L8ZbH43a0ckYMpabDArmDkD3lsdT4V06UVWvWhBPMt7hP8AnWQ3q9TklPw
0FpxsTVz5f+APhTlBffJFzYM/rh1qcpMVLa9Ai1sBOj/PEm1BgNKcB6UVNnh
+A2AApbj4rBMB1Wdo/06Y3fbyNRZAsnRSVbwl8YKmDsEmQ+3/lwm4lfZirv8
l9WfCbXVo+p64luC5Pxlm/Fvv0TSxYwkv3XZT9Zs8ezpGr23knTnjV12briZ
4wvCmetRv36y4AiGGoglqqUQAltfyhmMn+jQnCJU517SdSdFZpv0EHfdCUa+
9HyVkJCDav+hEVvkjjzU0e/RGIYyTq4RCd5/W/8gPhw0N617/kftSTXMS/hG
J4MJTuG7s9WA63UWBsC3e0ANN8PqtKHCUCexbgRzAMVAQoo6MDlTK615VKBb
bNzpIk+MS6wSqhjj08Kq5T2QagcW5OWHsfPTwzWRJdSHJcYCVgI/VrxJMugz
3emcMrP5raKt19a5pxfq/rU7fJz+J4LnyRKVtSQrTSZ92yp9nZsrKxXL9Mck
nDrO4XAIAocUZegFb1pDJb0lSgPG1YaSw4E/+S1H+YEJp6jWT4kAdM0Fl5kU
14VI8Wv1t5Cec2I6BRzGljSoarIFQV+joY7fXvH+LT8lL0+VxQ6t8c1kCFXZ
Af4meC+1wz+gxYlPQxaVtG7710yJnv35QQj2aut7wn86/xQ1V9ZT/hLaR2kI
pepuTuXzuCz94gto7+ghsndketlZAJQG9u/I9uakdHy0dbvewFp4Q6H6Kefw
clzwIGEFeeDCQOYx098YMSV1benrGeNJ4hxJiSLb6RYqYw6S8HLJ/Y6yovy4
tq0PxzElkDLIlDlKtirb4wJaLhobQ30J+Bpah4m8Hr9WHt7BuGu5/0aOcAt8
0CoiQmL7W3qwd3y8QUZ0t/2u1HBVQ/ca3vfpT8swahYa6L96ME54+0DDqUPk
6Ixz5THVAIltAMPO72XH+VNLLtkzehSzR7symm+vCwM4z3AW42Q8TF9u9uWT
Zh3SydrRdMLYII/jqHvIy6ZeG0pN+vqfvWxeUbQ27t6TE7ciuBtJ7yGYFek+
u91cwggT+0TTk0AKsWzkJ0J/l+S+52dw0kgyBP92wHtcEolapY8SqYKBI9AB
81brkPGP3rSN/A7Bc69SDqtFXF5Ci1BXs6AzjNhFZiNFNQzcY2HLjvMXFGQn
tj41TcpmfDSAqQR/VCpBMv4TokONVO0q3wjmRVtwt2RS5qAkAwOUHkIJb+sw
pYyNsZ+x8vlbSFXW9e4IOrEQw2JM6GNW19xDBg3AhKXqP0QWufxOewL/Lx5u
YoYrSEnVx0EgHv+XBPp4+xsxU8moVKYiECEp8+r67/CxAm4185eyxwAuCj8j
/+PoVJQL1GS4rpT6j49RNg/GfkXPXtPUm9+QMjoxJVKhO4TruEzyQpZonPMg
Gk9wIIbd6lBl50JjzA83FGsPDfJwMN5suLd5MDg+qPYf0dfar7KhqENZ1GKL
P9xZC3rvT0RDgHAnecDDficrVe1JtLvH1bMp9G2Siqz6wkdVEpheTza/B1hs
LXIjAU3AN/co4xdTKfWCxuQXe+rnkuQotsWUjsq4ccClXymFoS5jpSSaVk/E
HXgH/GY3B5jDRro26Ut2g+A6KbPZ+ow2zeANXQxMaYyMilZ/XlqHzEP8CyiM
kBy6twZH+65BrjsSCGJa0IKgqyohFSSwu6DZCSmd+AYvzb9wHdW1Gwqf478t
NSS2zGNaFd6huoXw2xQNHC/KZs+hVzGOV7DTi7s2zkalneXJ7sP0bI6yao0s
nqB+BUZZVAr8iX9QksaY5yxPEEDPyHnFDIOsb5Ixv8KGeqee4JaiSYyecw2H
fKC+pZmGP8auudfnNRhYSQOhVZK9aEVFpY8Q5S24NWFHu2ps7Myy/LxwgKln
PDjjyYRKeD/j9V41ylBCnfua2+Fji9OFRu4i8R4Rg7+qJfSABZVt6V55t9tE
WLL1m/fBWZtPBH1HE+CUS/FNa2yVdI2Tf7qQhGp4uHvQKA4QKUvnoRAUxIIe
3knc32iTF+ny1j1NAtpD5IZQff+VdR1R2RkxM7jYJaAXl9MY0wtMbebrOkc0
IVkwC0LJ0iFt6Uf3eMl3/gfmNBEoKdp85s8VjqHZbPBqPouaR8Bz9yIoyV/w
uBWrbbpNgssEyEGob1G8oGvNtAXArzk77O+gx05SDtZ6NPtGk4d+6IIcwqEZ
KCPxdypYw4y6imQXGNxlOXm8eS2o79ElqJCa3Dnl5Y09LIV1BFSXB6du4irQ
tB/qZAIkpeuRoVTi9Wr1eOlUdlxaAZuL/p5w1LHYozA4NbSe9hRpVRVyEX2Q
yBXw6TgBQECGGfZygskRODqsWc7gUEn12pGC6iQVL60BzATB1fjkr3aNG3sT
+FO5TXUi7b35+9YosBwqZrSHiWxufiHuWuhA3m8kPYF2ZpnHI8yBOiVtWsf8
6YsVNu8dTemQo6PDTyNzLzfx+VC39GKuD7MYj186Ec3YmQ7gJgaiwIZEztNf
ydH2E2lb0g5AMcdKMb1Z+EvgiaeRAH+1XIERdnlFCFM6uHTew9qSh5MOgfMm
LJfPPAO6bsACtHG5z+x/eGisT5Mr/dgcmvfVF1gllHXqo2HHftfV1mV6fbuN
buY7ELJ55Aq+4arJoLpxMZyflfbV9zFXtBzqmM2MKfCxIKFGSrrHx0bjMyP4
y26W0/YB6fUE0LHqB0nmBq5zPMH9/cNFlw8ubfVBk99Ymne3STASzk+c4w3r
ZIPbn/ggyF+msdBphc7+xP9ExwINu1+9gYpcaMNh2L8jqykbSwEooaqBBqQH
nEFGOchGWq7oh/asSRvJe0s/reJbE6/TmAz8HyTWoOguup2OOTQckJeA2cEs
PiOGUuiR872q8WRDBopdgnEb47/cou+v177IqbVzFFRIwHW6lFGe1EKC2OcP
Il/I2mqF3c72xxDOcFYQUvfEUyAFhIr/zMxIUGRQ7KfyIret6Eym8JEYru6D
208cbb7yNrFXMwSPvmbiEziMZ5dR2kiQ/4NzenG5+FObd1I836o2sS74YHXG
pOuxivPjuwSl49SNhaFq6ACaUXXC+VswReY1CecjwpaG6Lwf9NanjtwPPBBc
vdD9s5uiuFHnlJTgDBzq/fmLbYbdwovuQBj9yfZslxli/2Vh+3gNjIIy05YN
ALx/6rfI6Lf6B/8mTspoB2Z+s0xmItDA+IcDiv2Wa30cTWxpVOKHaoBpnqi5
9j2HxOq//XzQUr4Fc9cxsjhr+4DRv7dbZjwEcSpfJMlTZUsDrdiNfeb9drPK
Yu18Bmy83mlqSVcgs3WFdllTlL7FZHiPSUs9cIHwoBiezxel47mr7e2tE5iH
dFcXRxhCOWNgO2WEox5RvpzoZvWtVEN3Uc5I6/L1cea+ci3HaLLX2w+2L4hP
QnSlQ80EW1oLBYN1JH22txiPC8QYuyXKFpszfV1Xf+zT0OFuIQkZvUhD4MGI
0WuBPcLZmD865XaGPnah33lB/xvn8QWtdwtGzgPfaUzpLpXqTs58c7ieddpu
9FH2jlVSWbhcgQwJfpoPsVaOkwFyE0nDzsIbZj+bK7uawadT2GxUZxXR+h1U
MZ1J9E5utMgVJu5h69ybfY6tKWeJRrjBwGMT+QpxO8kD2+JTGwGgyCYkKDFf
KUx3bo1X6VjRHs1n4hwRx+UDE7JHaDd9DjI+1nhQMz875cB/cAf1zKM4vjoZ
YZYFx47eHW3+mybTT+kM24F3syb24ddmdPDhu6IfUB//1gcZE8KFc/PJpMPa
n9SQbVp/Y5pujGq4CdjbTqHrcJQ7MMqI5IJgvTekEnp2Xpnd/kvS3ftbpVsJ
vkPo1ArGcgn+99fAUD7BiZou8Eo/gNCvt3jXQHLDge+Np7GuqvR8am5jrcCN
PBVTxqyqr5kWdwAAiUmYQs4uN0TwWzYT5vf2I113Cmx/iG5DfckXwpZxP1Q3
JdAKYE/BoflIvIewVxsv6YgLANyAufNX04e+zUQfYDenEJZ9k6q4WDy9hIeD
bywSHo0RN3L7bmS8509HhpxE7Qcauz1cvNmVFQAt31bkYi5Rvg1yuuQRAjkH
rULoie0LqYtNfaEpsTRNSCBZev3l1UwembLVM0kpHDzNaOyqJa3n79qWLVc3
egxiq82pN1Q+LhjKpvO+rtBE11Z0Jqx47vLJLYjb1lTeU0BPM+RJXxQnXwVX
bdSXIw3uYFtQsE5jSYcZxtT/IdH7rPesPo0iboA1ryqVJJhe74S3ErVWyLB5
IiXwAKIbR0XG2moKN7zySdg9jdHth0HM2lwTwDwja8cZIx4YugD/x87tmGQh
mmlF4G59RwDXPCPf8Rf0e5zHvlDsc1oIc8yu5fMYNRsWIu0WexW5YGWJFneG
y5bQopqx1G4138ahMLyCAZkA4dPgkVhGt+e1Wa58PLOpYatoU6967kBAbIsR
duFKulmImAZ8qVWcOkXR00jQeFtzB8Z9Ajeo8ox8VB5FVIQXVXjxNWUjCtIc
D52wQGhJYeXJkxBsOJUsiOs+Yto2aELdCgr4YgZBobXO3LSd7rHGt/NtNTzU
BOUuZBkFO2U/iFMkaGSBiJIZoZyObU1HPwIzZppvKU2lGJFpqPpefXKGUGPf
aHnc0fYYnymjpmPThUz0SSxRGHEGliuPi1COAZ+95d6AVgQKYBtAEMt9Stef
FrZH7gBzTDRrA8/qkRToXWjt4jfIPs9u+lwjpb24VZP5Z74+Kk7EZn2XTj39
sQm6TlRsQ7k0tQOjBcOnZiDX73iY3TkweL1kxCKGghLCkhJLRReGRlUUbV9V
EPgi2tLF8GkUgaW0xDDMG90TIPSt/d0P9o+3k6hNAVOklFxAvOwbYY3Kcgn+
icYGwIlIbvJDhaK81bQl6XxWaqMcKugOWX05gYSLTLNkdoWJE8gTJ08iBr7r
Ca34+WODegnSoIoGbBEkpTHPqAyEi/Zrx5w31+VYKyS5HnwRV38s4YyAO5jj
4CGk/Vag2P3Ok437kNSIDo89aMCfWK95VznEdU1G6z6bUu5PuyhDtN7FfsfO
l+7xbfIfvesqUZMYWNQKepqhRUtoPOCx+q5efipcWckaucql+YYGGLYbBiop
dyGHlo/Kgtpj1LmRFJ1O4u65unzOWhBrnLl94qvByQJHzXfjdHCV4T6zTLpp
GF5qz5XSdPHvmnHhBU1NcfJOWPa7NSJv06RxoQEXbJAZ3pe8jnNmXb6OpjHL
WeX+BRfwL9I6IxI5MDXcnx3w8nie+OIrsV8lC4CzdviZvQa4gyj8Twcpy6Dj
+AhvJjnGgF/80l5zjfVaZFwOpKSaP5vdM6va8x3QqghrrF6HaUJtaEsIbpHw
DgFIIrVbMycLEDSAHE/2A3mYVwr7xhjILuVUpPwafOBDGVdiFFeEG36CVVI5
dEs8d1Pi8NssOVQaFmzR0Cvlk4MhVYwmpgPsCKm+PP+HK2OlKgfjAkh7P/v7
1zQyByD9MxdUpmXPDoAcnJNQfELdVeqxN07IXsB8C9rFP1vvECEdxYWPur0k
bueS1vqCBo+rEFVgtgH5MZ9an5m/oqdT1eYd5mO+lePKArmN9k3KQTqgbjEj
YG2dTTBcQEUImt3PocaT4dQq9ScL7tECTfsQ7omME5VmaHPb5yX/4I6Y0Lr4
VCOugceypGWLjvBeY9OtFfbJrfCG0fQnAR5xYEhkeG9B2UHdXReWP6TlcmYX
MxMtnzdndmb2XdO4lJIjPzraLJbkDasg65+nJPTqp8aMpCFVUJCfiZVZL6eB
A8Tsd6Y3zCPP7+rjuauCfv0cSy0IffGIrPtYAzfHaXw8RBL8wri1NQWEKJB9
S5TnaBhzpg8Q0qu3FM0KWeL5UFZLCDs5oRiwLL/lzQkow1kVrEW1KrPJva20
L0nnRiMSZyDKairwGePd/UMi35qs02Q5gQ0Cf6jNSEIfY46NCSt67GE2HEB5
PnNLqyWdHTT82h8tLb2ZWNVGkGuLHGxBB3G6UscHhsvv5lPNG9gr96X06jgf
x2KCkGfskPF0IyYKGK8+4ecW346o2BtoNjVy7WRrRz4gaOI1UjurHA04sFMK
X3fzaZe8xMGdpxrPhEkLmObpEB5R1B9dc0bgPViaXNs8ad4pnN1h8Bqb34Sd
gtvFMNWGQ048GNk84Up/Gfcny7w0eD0gfsWUabsomDBMt1jEnFeCdak1TndI
hccinrLDNh0MPN+MG4nZpaAQc+xyK4Wmq+zKiVylzOQv06vydQnUpHQp0D0G
7idNWvwuYUOOt0lgNbEExAfYYCKbkTFX7vMe4hydye19KhiuRoR4pQqIiq9m
xdFAk2dM1kTDda3Bcy9TJ3NMdvWGlaHJJlnJF5BqdREBwriqTv2ZsLIDMIH2
NY5N9f69hGC0ZGHr4HzCeTpHZBy/DgMp4Ui5FRjXVEedyVpufHGJrVxhOcFC
XzHBbpIoWCkqqd7janISvXbfjre8FWIBL59MnT+Zy5JT2GRrAt7hg9jaodyu
kk7z+KnhY9WM7+bmQ+VEA7ErF12AuwmoRg7LKyE3iUduer6tjH8D3K50D1hV
6RCRjznLAwSYkMFYboWO/YW8Ocr8jV3q+9zppWY7WLjB0tQaWhpZY/HkNKp8
q+d6HfnGcXBzes51wDz+hvsADaFiDhGiTLJeVRV9u2nXndG5IdO6IDbft+iQ
MQgebQyfEFDECPljPJ3jMcU0WLDtu04/ddtIta12ih9Qtjq/gTESyZI1XNTU
e1Ov5Ru7iVGrW8F+KmLJ00shBRzpCrjqNxOJTpIPIz/GFYJlsc8GqIP3Rxhn
SgBk5uRYiG5AY9XwlyTUESJO6Vix/u3E5P1CcIS3T6MR2x9MV3nqJXgovHCG
9xfMmbLghqQ2LBiIVYlf76p0IYJR5aCoJvsyybhKDPfql87/rNqmUgwhYv7o
IowoagNhu6wgAD1/xob+Qi3FrvqumrZzCupR3yzDLV++MbbcpAn898jTg7Aw
XGN1+rg9j18wvqHtEfCsOb4gYXAfQY6bI+Si6ZD6uXI4jCqsOjXAGUrc7K/n
oxbOV4KOYBX5qBP4GWb4TBugqbzToQBvYDAeg7o+H8wCA3Ldg92i63Y41/91
WayFvPY4Xl+q4c5oAOatMDrkvjwyXTmib7x1EvMHgdKbTHydkKW7MOK0OmUn
i8lDQtAsO9crMaRFk1cXbaLvAXM18fDwENIqzcPuVAJvjRSh+aySzY9RBHTg
q9bZu9IIBY8Bc2Jf9xtR8ttyMw4E1B2rfUlYRrc86ZYnMPmwrdkfXE/COAL7
Zae9e6cFllPArSw1iJYKQ2I/I2GJhP6Pomg//w1WPZBLaaI6MN0T60C6uboq
VDyqcr/xEvnGLrZTTgITjoLDjyxmM/DSZ0TVctMRGGFnBQOBn4v40iUNEieU
tb57e6hWWAuL5z6WCPjthf3O6ZW8CBwssESmlHnvfsGoagPuxldCVluCKjLe
tu11eHFRwKTOg667MjgAfCmNQgm/H4jaX4hk4LN44wgYSWbk15HOOspK1PLl
Jco7oJRRjn4y4VEe9ZlgOPY5IDZd+8f9S0+zkg/pMyherdt4RWT5mzsPN3PJ
Afpq1z7HBK5ftjFI4YZcA/ETKnMiAsMVp2JvCMmO0V+4z5ecmM1Ey7rMOhvo
RtD8S7b65Z0JBMTbHCc4kiLDtQ/fJkhZWiKxHk9AXTkUdoOMBomEhzOXIRVx
PtHwlJxr+iCmHHe3h9aqwkSQeajJRiSNyZ1qP2SiA93ZeteShvFw1t2Kwe9d
eWio1mgb24T9mBxQ+P3izx19RK0sFTwXkM2nv78kX4bsJfervVexFwYfuDQu
OYuP3uNkguQrxIr4DzgNZU1z/ckNiQETIez7EP0c09J1wKUQ6Dgz3/ZyM9SU
NXSHMLwPODREb1TE1/+3dtRWZvcT3Unlm6B7MCtePZo4DW89azwZH/3vrIXd
Zp8hE4UGs5/tEeL2IIJVm5mylvB8lk5+3V31NNS3NY95/Mmnvs5tgl/4YInA
79VIBItSvM6h7PVQ8ZyNUb4fhoICxaHAS+UWUPluHSzqymHKbG1QFeoxNqaH
IpGL44iXsVp8kRBTlHOr0xe3Sq3GS2oqMjVL8PJUK4yZwjUgnF/1xKtOxKpb
Jt2Rl6G/DkD5t10NPW31YFsHwwLf9Utvha5JCnuReVX8vhn89gfsaQraFUjf
mVEqFxEBcn0fRwvXvjIpIpD99/PLa2DU6EaVe7ra8+apuptiNMrAiJURDw5r
sSGYz0njPvxqhQtWjG+E1x1PX0QzrZa5yuUHkbGoOwF+f9FibZcZvCRkoTjC
3rckCV9Pb39ZUMSgRcJEQZdNbgZhw/bFXY2NLfzqipnZxesayH1m1W6Hk2El
/UYV/TDxCN8kVZ7AH8Hn7KtsOxDHhjMdc89sG45VzK2qKDd6vwAVs9rgKufC
nZbvKpucgNBCQl9lO34ff58L9dfFREVQ5vxsImZXxsKo0t+CTN+54a+5KK2h
UdiYbso8wIqXw31JlcLp2BI5vYebobUIy5gFQeipdKcfoW0nEwTfKX1a1X+g
luJQiO++e/BK1W+fP8mAS0nnMUZRcNXTm4zdqFjuT73p2IAmq8BvZfpdRe/+
jk7TLwmdeHGNwcOz2NkLtakGYVr7JFZ1PSMPkzr62g==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzchl4DhVxkHIoiQ0dW9yReaY62LuglwuWWUcIWdhkCTrh3siEAZfjZtvumThnzW9KO/55jJ8Y0gq7SOSFum8pwtTw6FAyGd0098LZiOlCJfN6+NFwh71G/JgNBcg6eVI2aJqo7da0+fbAeCx1kDzpnWtWvMtGGFR3MT9+FbAGrpwX94utUSxg76QN1Nfo3EniRO6YTZCeKJIU9vB7liJVkX1vmoH2E4twok2Fg4K7kjS4u8PehQNN7+K5DcMeeY8lHurH3zvxIKvPl+xRCnMwD6msbMGc6qbsjGN9AK9YR/2LUoHxDfo9ii++oq1DdQu49jXKWiD+Wcgbx9TGeSYKTxTTEdI9lXaxnFnjMYLLcipJt1IUv4TTAjRoCD2W4EHTKxnOzBW2x0fg3UmuUvKnrQ0jbRbtq9iyW56fEWaWN9Jy9PeXnMWlHFbwXq6uRcx9NzBEVvCVCDKtsuL0Kuq+7rYpFAbX3x6GiC4uCKpZ21ZZv8Fl3F6KZw6iPGS0zin4W3bWEkacQPBEcPAh5WmuzE0ZFp9PJiplZ3iK0z/I+EqD5HMZ2RM6VRqrJyjElMG66sIPz5p2ch39HUqgGnVzC8SMibqMrx0bIgEBBph4ggX2I9MkDRORffUgHdcai/gTFMJh6mISnmGuChu80XfJD/V8gXRLHqAs+unIfUa3LsuHg1hbEEBSpC3nS2lmQdBBgKSJNX8MBLkbLnxwNXAJzR18MxsN6bIm0rlIYolf1SdQACtySd0vNR1iPh2eeiP8CtL3MVXx4Vrh3XXjIynuLa"
`endif