// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
tzwrIUqAN3jZ6FwEpsVa5OUIa81veKyaJdzHSybq0wmDcHSTMge8KxBV+KJW
2d1sAbWzpElLLvd8CIV7vurT2SFv9zo3uVLfp4WGETQ2tta1XEzFsGIT7pnA
Z7bdc+deOc8ADJUDSwd9T+XYzg4drW8GHemP31eePMlJrzOxTCB2aq3blNEp
C15678sGzTxbFZUrT/7VL/4pxn5465c/sHBBMiwZxoUX8bUD/AZRDPpIc/tv
Qyure5lcs0ItMR1v6+Jz4tt4S9M9uiA3meOIncU3/Nic0z2232s1BdhjfFfc
W0m8p0KqfMx4LTsdyOQNlYVv366/PHmSF4GRs1qOIA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ecq2Ew3mlLzqlFN3NDk7slyF+8Pw/NIRqhLan0rKyIgy0ZjA4zR/AM0CROua
gIfzShz+aD1jh8h6/iptYQRxUrkiEunqFGyCNcUnW9IJAQSm6R0CmDfWi4k3
xNMdGAP8ZFQRZjCpvl+yvhKyeFxQcEo4UgBN9QxgFtifvCJi1UxGBQF2XoYY
VdT++MrNOtsg60TsG5G/EpEfI/UqzF6qJPEVFaAPaEkk/vHgv6Q3WwPBNU8x
BA703hrzjO7zM8Ye1iCvlMnMIVZC2RrHTg6cgZdfcpMxBCpZucThLmW4gfNK
/x+X12FqydqnVaj1tH6Eq/Yf7hbMie9U3l8zioY2Bg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
avcaXZ1EEZat/hA+uOqaCI6TyECmr2gkf+ZSFFg9zylkpQthf/ZeJSCeV5tI
OmyWFaQ3kNmz1jAnO56+krZotqFT77ROY3K2SY+9xjQh+5GkBTGBb0tWwECv
6GSQzVl3Teb3aY/qGe2w6OwCyw0WI29pUQJ7kQ+W1Qxpxt+7d2mfXnHaSK9O
+8iYGLj4am2iMrRqUuqqLEyoU2+3mwWgUCZs+lrjpjzJsXjlvMV7zHrddt2U
59YW93D5+s3/Mcm7DjdFORvRVCvKfGV0C9GpBwHoW7Ru2A0uNJaD4GB/26At
6tRD4vobDxUSnyWUTcJr+VnD+TlIQwK8RuRsWl+wLw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DuHPIjOngSwc/QLVs+pvl9x/L6KcPOjSGxNqMMDwdwsjDUDPjF3ZSKSy3zlo
hRaQ8IW5DcxvWADR93etkFy4RG1ObiFUjywGHo+dluobwnMLZbsDD8VN70Pd
Alq4qnNax/gQSDz5VEUIhHNsLrhuEMzeTd3gZfCJN3U3LDvo5LVSZ/rbwBqe
11fmfu/DuDn7ZcGPKMD4EiRMOS4j0AmkI2swfvNtvgj9TcGqy9z19fspRONr
V32uVAOYitSwwx+2Y/3Q7BSbhYMrJFvh9X4SDPV4lqGjTNmpwFWgW0cMDFta
0FmP9T2hare6XO1Ug83eIB4agOmqCGEixZ2R8KlIbQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
n+EQlymXGR5JOeWb2TgihJARw5Ar4DvnGipIJQD3ClfXUjt/lL1Z3dsBPLaQ
fucJjpCEPDJpEtzQlgQoKgElfA/opf1wU53PYYuB63NGgyrEgELGKDb5+HB1
M5wHC5NIKFgTC2zUQR+kvZHfrQpyCa19wvYYZ6HuMVPrBg/q5t0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
wMJnAeQWWEpP4zX3x8ZEbtrr1oCa3w9OviG0vk7TwQJ6qvOyabRfAY6RzU6V
QQllwdZ79nzKECPw4PM2HVEDYnqrULUkYdM/7IwbdLZ5fGqglIHBNZAMRkAA
/ltym1TdiKp31hpvDlHkUzjmUWF1/M3dUaVIY6h/ildCpVkVkVbjp/OH3oog
y3DZMkLXrJjSMlxc1aMr+uznoRHSdY6GB+E6Qb2yE3pECENRkE+G/usNK94Z
ymq+m6hhnfCDGeVw6DY6crggY8FBFW6cKIHsWtnUYqPCqPG1PsjTQM0FK/P6
1mOSgY7b/3b35ApqEh3ptYK2cr6Cn6yzexHIMP7jtrr/oDg7GnVCt09lTOxh
XE9Y4HXenQrKPDexjzUsX1rkjD671picKnThj8ONysP7wrGhfcm9iyb56XJt
x0tojoEnfEO1HwFm1QnM8ey49mbEJXhalYYzCBGpWu2R5llQCrU0fRpkNxQr
RPlgSl3yrBNNq6YEHXrVUVWaM9YwNij0


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
d6dSoF+qcOYz/LuoyGx9YEP54xA3Ta+gTCQvvx4Ph4xV9EEKuq9CkxDpFqrR
RHhPWDnLIOBqpU2A6+fvCx3OZQy3Dk6Nh/Obo42Iii7bwmHuRJrWFMAAPLfI
Bub9PFdBOoV3J5rikhBtelfktMIENH9p8AWcEaa6iiauJ2fj7LE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cIYjqcLsTouVXtA2I1eOMAC+G9o5obfQAVVi3+nTA+3BZo06K9cMLE0l+56b
VcQ1UiKpG0JUqAkTZybiRyFMme/7Q69/da4SNGPWr0sj9Ujncbt5e61F+4Jm
H2O+BzvblAkANFj81HwDfvSqV0muTMqxkg2mr43RGZ8rlTF5cXM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8496)
`pragma protect data_block
DsZemgeNynC7Da+/7GmMLagW2R/zn6191wZ6z59hsjqvW09QvrfAY4nyxfaZ
mVoCoeaI/7agG+ygKSp3IxnFtpV+y5vjcHYn2Osw//KuVr3tMqC5gcllNT1o
1b2/3UbULwtHSTRGJTJsL6zrq2dU/3FYbGM0Vda28V0zYcbti67udXDV0ZqU
Xdl78U+ZjLiYHLAwZVQEJsD7eKaCZWQfVu3JWH5qg8yeD6tvm/UN8nLsG8sC
L+Ay/CyvSHyU+Kv52+LCvYV8pN/3EG0W9JZ03wrdI7rcnyjyTQrZt53yf/Br
Iv6/wB03l7ldXzWTkiWTquK0zmyal8zqLGp0oi95rCvvUVqLO4P7KGPyIE4Z
Je5/3n5Csy75ROCh1fwGUwMUBZ741f25KrPmSOEBmY+0yKIKGD2iO0kIaYnN
IhK+fq6jvAMYJCmPpAcU4ofL2JOOyWRmvdMiCqqmWH9yTbzB/nnYW6DwLfE2
dIAz6jkCFlbiV0ksmiugAALB3X/OJdskbaURByT5s0gFAudXHLs2q6askY/X
DUII9CrKl6jTf/mSj+rJZriFLFE2BuzjnLZqbzE6wa2qKbhlwCfjAbpDuZTO
Wejdy6mhjM7pgosBpJygAcb5KiCRAtvfBc8QG3XJzTAjKS3vM3AWV+a9SFlB
HrqMvcD9MoX8bVns//vAzcat9TtAyPgH/nRggnjlEE9pC299lGmp+aBGX0WU
G2PBIBzLtLAkDAaGizu1lsUoVlQT6+L+afYxhlRQrKse/g1gFZRG2TiiYRE4
dYOeaDWyfBx02VNq01yCJqv1NBQZ3H6sc3tvWODdZfIx6/+s5EZeIScFj1Kt
UbiVZBy8UYukpYl5VZs0cTLmY9kghtPhUpQqFeeT6PlNC78K7mtYNRqn0yi7
7r4VlfnqPrnbgTxBPoTTWWIwmMEhr2sLv/EGBFvruq0uudZJZ1KiVB7sXyow
5jADY7wz6wUYHRoUYzMLlMkQ5XKeblPy/HVNSWoKpKgNHWOWrYZbexG8ZDqE
uu+Fb9neKjcab64ff96cdc4992B6XyKOGmTlj38rat8JR3nj1g8ZOxSMJZIg
40J3i9Ag9cc5M9jnoL0zbTqDqIZvDWe49FzTBCfByhliQvzWtrYaI1lj4BX3
sRRu/FynIPtWE1GHTtulqu2uSIegUALoZ3aO1HB+20VB7ove0R5YvvzRiS0j
bU5oLos7Qu9UU71N7jq+o4ouaV1opz94fElMbqbCPLYnoOH076hdrBXIe25p
E4bZmyk7pHr0vrVQYWgp46nHC1FWILBioJt2/rgPEdubL+naWmUZm/kk+XRX
PbUAxN5XZUtz+SPDlWvu9I0cXPr6i6YS2vq1eMlBkPQIVupHuLhgAibVXY3C
6LLvBt73BwsO+9riZgpX13ppTCa0aUVcEuCtt/5IwTey/mk7qoztglzwmru3
DW2yTxHLg7w6WzM8Hv5Tc6rMtnUbt4Ib9yXh+xGoDXtXls+n0QV3d+mPkzXl
03ey+ROON/umE7nVnwE8PQVa8sX83m+hmeILolI6I0sn3guLNeWUoiK2cRDT
UzChlh2yyG6++g3+WH6ByCW8dcnZ20jc92kBR1xuX1AaBpU8Xp0y0YJ50A0G
2EqOcdECGCkjN5PJ4963fqGoS3OClkpOcz8h4zXM9XXUU2lX9Ua/nEqGH11w
/29YGyMX1AZFZm5Lfvqb7mgCZaKa+t4QbeXnQsWBSdkxrbmLLbgSj2sIClM9
lq3MbuiBlKGFZqA3Shsj9d9Wu5u0a2jcjTdLYgKqknp0IVW05o2K0Io2tR+t
1TLp0WwrzzykBMbJ16DfzJtxaY8sKQeolfztPR1adQf2d//IuLADRb/0LZDT
kGe8OysiGeCOFLMKIwLuZk/92EOGiA253o1U0OeUQE8+JHpzix0OQ8d+eLjk
IdjG3n0BRhosCJntWl7Phl4Sbc/3v3uQpIC7Eutg9c5hv694jZ+27eavYJF7
HuwYFAxVJ3hDf4lI52eBS1uWT3bMhChHLl3LgrRbtAF6MCVF2HvC+3mK/yCQ
ybFb+ZIjmPaV/4YiYPjUOcW8JdCfWMfWuPOE+QuMFEJDoKD4urYxBHAbcGa4
nqZ94A5X+MBMU255u+d1hR/QKhRArMTBlanH/uimHrUo3ZnQgsJH13YkEVmk
3JmwcgE8xEq+SgvRpI42qJGPFBCOQX2XF6UHnKx0zPaF0tnFJ7Z+jiIeIDNy
Rm9djekLzSmnvLwCVJPNMLlddPhaPqq6n1HarLBJUXN9a4siLMLWKwGqexdF
txx+trgjy7iNDH3v7ZUIViBsqAoBZwrjYn72fJd8yzpmemXsvdL7XGMw8KoL
tyBQUlY8QWviPzYsI0zl/+HPGw3E53QRCzM+jVipb8+kkFteU8X5PqCyhGG0
ZMtKY9gtDCHBNMm3dj3xDdQN+dUZ0OUdGpWCxZ40oSv2yrZH+0V986mlnrEz
TpTqTCFJG1Lv8HPT9UzloQHufSiNvAAxWHFE4xe9YWuK8ojQs5ZE4FHgWeQ0
w6JjCwz9RqJDz4gY89ANFgdraCGMhxur18lRbi5QMTyMXIifdW/1Te/V7su5
cugqt3SkxDmCoMk2gdXXhOKzrjUsa48HFDaEMk/jjd6IakHPM2al4lElvfw6
ZdmWkWqgjfvnvNqFP6oXBmRgUUDY1ZV/BezotpZrVebDRklluRLNLT68QPFz
UmB5DGV54sa02tJt5dPIhEDoMLC51/Nd1Bbo5CN1npc2QDpHp308c/EKIJiK
mjyinuMC5hnHaKrlQwNYAeAA2olKbVUZPQteFktiY6YOPMEaAt1kVfjhU3gi
bJzAR8Br43qN7RotYNqg4rSrNLrIRFh9s7zckNV1mUA034fO7fS6OgTDPBod
F8neSGuJ80h4ptRm8xVcpgUdXVkDMMSoet6JwSBl3oa8LJZNi/GPtgh4F4I7
L7Bn5d/7jt94ToxqcwZ7aje6CLQivoCWR3Mr+TKxeTH4ye+p7DqtQ4Yh4cAR
09Qvn2yVwgMCaS0+/ABtoOaNzi2MgQPWhzwru7cwsh5dmYkJI+C2XBnYekWH
L5ZbdtPchPNOxJrKyFlNqzRg6peseWtU1HkPt6G/SsTZRd7xtZNM1c+Z/03u
xTWSNTDlIIxHBtmdI6jUSeeD5z/+clqynOOfdqFKR7zCFZLKB0b3pvSBJyFK
gb5CflUpeiO47DrM0vjcM9i0jlsR/e5m8hZzUtIIydSSJVVGCbZ+fSe3ljNp
4bShJzE7cSvl/UnslbTSZzLad75IQsbOFF/n3+rS/23IVFf5VNFExIa8oQt9
Sp/gegZE1Wa+UdaeGEg8YQhlPCR1ihXtASh2aTqPUzXVcthNx7E/vHiiz9pL
3GeftxOPHmO8M3Ag3dZvthMhGRlvh2xL0o4bbgefjvmgciaqAqWSYLK8ZNd6
FGFYhHZ6WFi8aOwQ5Q0MXGS3HmT6c98cvwJ/4LiFQ3EzS1camY7VYUb2Gb0F
3TqZgrWGxk4oOpv16RWCfotbKyl28qCpbPpERTEvm17IKeX3N4j7adJ9f4GT
oW00iaPj1fIyj9JFDC8Vl6FbqtnyoEwGwqLwC0fu8Cq7IzHFj8OE1zdR0vN2
qi+rqwm1Q749Cdhw/ncEaLpQ04Xy4ggUnbHGClaahU4UWMmYXVQtgnWUjHq0
g6b9pHBibktZ4b6yRl28gbSOQzIAxtBJ5wszRhmWcZgj9K3lyjHrk3D2F/Qt
9SuKYGawh4V4NcPSSCuARvO7bjPI9NUFcn05Z5s++rxFhoIAB7urMdu63obb
3ZJEoenuPXM7T059ekhlZJdB64YVKiIH0mx6O12PpTsM8ArmvPMVk/3tV9YJ
FqF4tP4JCCZrecx1gH1MK6XzkZLfarRqCVKHJJlzY/NDUWVmg4CKNZxXMCvk
LmHt9xMJiDsCRqrDICuy7rpM72riSVAd8jcKrJayQt80gwZLsD0oy3D1BNGm
afpDoK2xc9csYSDd/ykvzYu8nB7Fv8nS2SuKoCctdq1DlW6XZ0hI+3h0A5QP
DxldkTZX1conHDz8aGnCAc2pjouWbvTWOyTAcY0R2b5MUuInUEuALjGPfM1G
eBOD8Yheas1P7lhOeSeyoCSf4Rd4H17nUP3833P/teG8CvhODY3Gi3dSZino
1e+vp3pTPes2q1PfdUCZ6Fc+dxgfpPHQ8EIW3uhY1r2u+DAhhRR3fBUaqt2l
FT2/EASIdKrKFAWxOKHt2EIpziAyLuES67iJmoyhpqxum6E7vQCXRl9or0tl
U2Dclg7Vz0bduDpI/8rl8YCFkmQm1CTXoqWmDNuXhdsKPZLY1NjO/RKzS+Vc
FEpQl3e+FEiIXvIlSkZi7r/vE7SkJ3e6zbitcIKgElGg7LnHxuLZw0PpWbcG
8K8J2QkXPKyzV5s9dXE70OysMxgS2sciV7lxysWHkiOZLWGEtlb3rV4Si4H7
rPx0B8och4jSjslw5/AViBtimCsxgdAp1kIsrqJfMs+I9MRIyKieS2WNmbcX
fw8UcW6aT3+zd3dxz4cZ4kGaKoThf5raGzs8zf0V8g7w9yTFRC9xDh/aMPYN
o2iZIy547ukvSjP1UfMjhdeWdOSsFTHiCw6z5IZw2uo8c7EXHne/jgEEfEPx
dqQbFKgSKtVqVZTMOJLKcspk3QRRDgiemxQ95sIdgGGw4BoZGYT7JAe909U/
Hl05LP6cuFPCuUm6toa3tP6UiTyfUIW0DP+w5GL0sjgieVvu3t4WRvPRvNG2
OhyJmouodwTs6I/qGgZ0AcBj/CCdY5mnuaiC4BtyvK3R5dIzNJF/vCe8/jZ+
DqBswEq/PVmIN9K+x+zuWfYe93JinbphHAC3wLqeZ11jqpKpb57qXIFJQdQo
3EH8lobTz7z61J9nEQhjhM35L60K5BXsxsnkN6UJ6TbPlsbatnuOaEjZA4zg
OavjAUEVOgp5CwzbOHqFXlkExTWShbOa9TQnTTWx04KL+6R45t/YijiiwhLi
tWK60uGMElaRQI4O4mFm0XLwO67VTb75+OzXV037OV7O1e0VEAz9QvXLykou
mUUaqbSiuShsWW9okhDJ51lLADvh0TWjEHqVi55NiviXuyMXMDgc4g6h4F3D
ciCDsGCrJwXtzdmtAzKPM6mhwD2JYDhCnsHaPvFaTZGhV2TrQk7SIcomfgIF
MVcUL9M1+H1Es0Vih5X0YPb12M9HhE9HA0rq4IMaF+IW5adSxZ3+MdHkLt10
2W1+rvkB1O7WIqWOPzjjR1Thrsco+x2cbz7MIF7dQOa4/9vQaH0i8gL5kHDc
ZURmfU0p158Hel00+V0EcvQ7l0zZwCNtfSJG+4p4CrXTF0HmWyus60ZHgUG4
ODiakt2Rzst3bKIUZI11j9/3x7CP370OoFO9bdMz/w0m5l16HjsP2Ie52SFv
wxxfSA9r1B5cbY31pqMV/T5pms3vyrfMU3MFKFzW3b3MBIWZvZw0bDyN74Lm
UnLStSWtuOzLXChJGxgQl63Gxx8tFPU0TvywAprMKMqoD2XR18LG/HCZMOVH
owbZSs/nkXMerjikzElRdHebKjht4NJFIU7FaGBSU8o+pXxQWZ8rId5hVDPH
1L3hRyPHuwCx7J3Q3lbhEWcQq97KMU9cRYYS04pbIIKBeSsfGAa7/WUX9tKq
g6zm92x5fVltzHDxT5Cf5rFxCs4DfhLYM2Ca8FpIbr5Oa4MfHsiKlw/NJTQm
zeQ6rJDzi+ipJrQLZQtQFYNXtsjxqilLVpIM5uldv++6xevRBYR5ko+myWiQ
8IIqz0tWRYyu6K4/OWJckF/29ETNpOZW3rBemEwlWYpRbv1G8LIT2JQzUjFs
NEWStji4StkiNbOm0XYgP8ERAaPCxgXWnDA0ApjEQMcjQ+K8xsFsFdMe1qdJ
jimogRSLG+XUMh3delXErLIhXLO+j8I+xuPvXyT0QZFVZX4BnjpVD4JQu++B
2TbSsrKYGvImIw/c1oIb56/FZqq0B9hvTEBpRcZO6tPaJiNK5xQk3PLaKb3M
ihEhO93QeDWUVU6LBld1anpVyI2iqmMlptVUeMMVQiu12hGYDWl/+2oVsQRe
gqtXYTfHveINyf58CvliWpbcw0HSdvt+TJJC1xr1vZjwlUfF2PZR/cypNTTL
m/D48bf1yEy6ruZ/MFG8ytwtXxTLRWMbTyT19BiCsjOZ8f8ToNuETBbXmFg4
UAU/Y00H0IaHTvdYsKINbfi8yClTUGVhXmxm/+RkVwebm6zzVKTr+qI+xPmq
JWsoI5EjIDZtj9CkpSAcI0SLifvXbu0OZNZap9NRiHJfmms3NBBEmpQP3eia
8f4P3TOLljGg7uWDewvXqKtt+UMgL0/1hQmRajmkyOWQZgiQKpl5ZXs8zze7
yTp1uhKijstBRCBHPWZeSRbAtVvB6V7xRt42n5+ubI7VkjGdOolgw69Eg3OV
ofZ3XU+MJpHgphZGdjvlrBVUSDISRifSCUNCm1KK/RCIZzloBQs1yos8lq9O
5aIm3ANJ1cXZN6gzh5U5RahhY+9OJ7MYzZUo8Ll0fcWP6oRSqWgu/7yOkfH7
1eqds5LS0/0DP8uoqLw6D/TwwrFwAHda31EqAYiKS40Sx52obRcRKYqkV2cZ
FFbzC6nCnYHj00Gwb58U6shCgInTbmGJZthHtm2cSa9RdUNpzsN4G8xVre2D
x7SeR1Qsz0L56AxpeoyUIUPMiF3otGT4I3EBy8tlUsUQoDtwDiqXQNV5BWFc
9FhYS7VydIU5yaqBFs3G524aqyBKznHM7ZaiVe08FuymL6ebkyVPNTAJv7qT
jeiuk6xW38vIuR2fA3bdHFuiT5k0xd07Px/1wvfBHnU0Bp8uOJOMfkoTRnP5
1psy4fmgEYXjgen/r3KPR5BGLkFgm46mVffvuLWhuECEN2vSItjA5yRwNbo7
pBaicqHcJ4olB0yqqFBI7UpyGgKaPlERiCoCRAt5u4JIw/yfyWPLe/U9LBO+
Meabv2NX9i51GwSZ1U16FJeTdYyHnatGq2E5WHB9OUnhBjyCcj8xxk2CzKfW
mSux9J/oqs5wHICm2JSG5StPwFPJtuxd5h8lxomgBGoRyHfkDKV+sufaARe1
H2leQksZdh2FbXtPkcte+xpk0CmOdzjYP82kdWy2z7GbVwoHlCgxtHFdcSq+
tULPtqOSgHZtn7YDoKhihGen6w2LbpOy1Y3fyNKgMK4fY7pwQBoK489XOPEW
/jaWVivJ2rzsW4pzKeg8AJNJXu9femw9sL4N6ILVKgJjSet5FAItf1OObgk/
BycEIEBKqcNoAn6874R9gd0YtFY5OGoGVT8rzrX3CtPTeB6ZPBO7EoRE+Hne
Ie+KvWokg7LkejnlKx6D8f/HEpUEfAzXxw9pPTi1YhMjW0y5hIP8fIc+RCSv
mVVXIuJbuTg9ufSpFEt3zZUitPwaA46Olu7ZmIfHhLQ5ZdegRkk1MWiIXw5L
eJny6bBUj40FZ0n4N5K+MdszQysaaFK7jDVbMMu5UKwywyPd/bhrm7cEcBfm
3PUCrHDfbGqxaFopDF8O+xHcyVl8qMRjeOYiH43POY2GVlJJ9eQ/Hy6Vc1ka
lAd0JFVfDTMkuYf33wYuzDTYQ5biM68wFZa0b4s81+7ZNJamPFN11TudloGG
Cv5g5f3xh8qs2JFsNx0iFrKZjxP1zvKrW+fP5amBzyf0Ah3REA0qRYgNRNzI
lQa/r1H3x3i5Py/TCI8UQzQUPukJpsbHLyNE4x0hTPTCeFf8ZWAGfEoPhGZB
xCk2cff60D4UaB7D4Z2QTnYA6f+gDzBr05341Xx656ZXtAwQ2zItdMpMId7G
iPnEDmPvWOGv+NYuQCH7WuuEdHIUCKav6+8/vM9dBEGFAGYehgkvHx1DfzWn
6B/G6tvQ0iUnRdm14uXMT1uP7RZ2DWl/wMk5OJqhIz32UpwPAF34j3kdPwk5
5wBU2wTqKAKFz7gAViKjdjTcwLiDHgKrdWl39McYUR9OuNkAVfNAX7aJIV6P
CH7qM2CsbSDtcMRAp9cG6llz5T5yX3pG8/TCr27QdzGG0CQ3tX8QVDBRMquK
xhDOjhvzVD7rAUNIPCH0uHH4Vme8Ij6ZofDoK2c0EVg92lMzny7cDAnXp3m+
WtkGcAVPieE4rhGfdnal35ck6aF2rA77J0cFc98KYxdfvtRFtJQaKuF9yUB2
jGGFebSrCuPu0vr5IrluzfAOzeM3jWiW4Dl2lyn17Q96CLKjreg78AudFtKI
UjfsdGF1czQZM0leFbgWB7h4iXq4xll3LWxxtHpVIpwRQxxBnW+Ld1mmHes9
vJVCVpbstFYoRdF90DOrLCMKlnxAB8B4HB+scC7ixGx2oTo75StS78KvJeZY
2jhRoJzHQ18R0UR1iDm0GnKc6jE/5LCkDozLSH6J7eadjoWogtuDtTDG0Oad
JRKa+2aJbZZ5NFljJeU6AoZlzDh28hKgcay2sxPefSfRWm2lEkD3Jm3mkeqd
VtMzpzBzu1F4LBD3N5RKsIyaC9S9+nMWZwHiSpG2YQef71h6qLtlt78Tl1nb
q++L4AtNSkqbQ2mf1F0B5eCg7lZz8xZJsCxKh1srWGXJ+XZbSrf0LMnNOkD+
rI62IBzgKFeDDU2p4drX0DgYhS2QIvlOatgFQTGg9gX5o0XCjmAK1h4yBjq+
rrRNI0ckEuowGmMXbmuhOcncPLyxTlUSTnifs1FhsDELsBE8mgGzsOOXnrqS
sm4ZYuXO3sI2bLvIG+q6oPbkx2WmLSuMUM9Bl82jA5GO/05DNvzLhJmquM/F
XH76EGdNTE3Z1ykz7IZcCAJkn7k5JjNmYikwVnajgKQoPcLNuEGPrhjwpULG
ImsrjiuQN4yNA9GdojdVpv+/ESrYyqmWP28ta8Wk9FFtTke3l3J4wl6gnziz
WXP6PRQMHNZoSWfbw5hQRDJ8aET0Ug0W1+4xHx7Q4SsV0I6Z7m0nPy+4ZITj
V5WhVeeprpT2HhpRb0EFvmSCS6r97HMxg6frT5gsERJObgE57Xx2x1fwo6Ha
lStqVGuZ5l9JG35l+ZV2r9US709zBxUEwFcuIDyg2zm7jeIjMsvKBmGNvMvR
+tg4ZlqkojzX+xSzYUuxd2Ho5358oYB12OV+FIUiapjzTd84Ws1uLK0FCp0A
R+JMwMK9Z5xSCvFlbY6vjyreq4L1fDc866tnW98hJVxHObzd4QuvS/yM23zK
hRziBxTvYwG80iG4bDZsVA9uvOLrlmQ56orymBeR8S9TUHacx1kuuROyL+Yc
HR+Me92A3yyhxL/UOdk///yBc+fXgukloNwHfsWbcyyd0FnhYx9nH9SjqBWw
65QNAJU1LjsqKTo15s3gm2GmKybCwuDKOfhQNMrSnPGek+f2DPyvIWIB/JPs
+rQVfQT2EuqwTv33Gy+y9yRXj9pF20X+dtfsGHOr2XKmX9M5RZgGhXuqvjBl
AoHgMRpS2rsmr4fq5lfNQTnbCA9T7m8FMbq6k0lR6VmBiZQ8qBYAI982Y2dE
38UdMaT7SOnfBtow0pw7bFnfGiMTHDrWniHQFf5AsCpH2WbhYDDR3KAJZloG
A2NjlNP+LeC1W7uyfX6UU33TJQbv02cljwrZwQj1QBrQZxws1MyAOPpsg3IV
kvXv/21fOMLEP5n6y04jGqAjDAFyvXQxH94JHBIgSsNepl+lwDZri/KB5zV2
i6gutdDln09WphRsJDh84yMW6CZcuJDSUjjn9C3BkTL5/zEkhditq8vyHteL
z9K9rV3dQIzRrlVGfOuFRWN9Iuud4FL1yseQ4nlsSllORsJNtaxywxnlV6V7
2/5iNgzNlFvAeFR+zoih57RkYupctKXFL4W+xYC6Q80Z592/go6gRZGEkW6s
parX+IJILK2NdHnmh1piewjl1OPguioK9u032ce1fR4JSbh/N5H8cKomVUzV
S+tpczR1I7gIhEFTz2V/cfHZGoTn73WG0q7VVQHC2cQ9NOWHIc2FTi/OCyaM
MejpUh8nUc2FvWe4dPozCmGeFcS/kP9kzRvMB4fC1r7mNhMj30gzaJAoPta4
XetQde7904OI2gocDy1om+qLGLAZxx/Ugqemo5P1Iw//mki4pq2cUKwcn6Ys
FKsSJHUo8jxW/9m2TQl+3p2zpkjwymCOw7FA0HfX6Uk0Ps5yXrt/ETGAIc7N
BidkgjxmAEuVcGBmLsmBM2pgZO9vdxNnghCgUFUc+xtjw65Ro3u+dNzHXozc
L7QKVUomcCk2poeHzHVVFgwepnc5o6AtciNEwF53ukagnWLITXrcv2OxPnbY
5lg9ziL0x9RLL4ng4k4CWTz56NEn9SPXZV0J/wc4WVPihLYGSk2Bo4j1FSQP
mwzO380ueVQtAtGDibrjDcpIvg29sb9g2s6W3DceMreQmq4Phl6SjesXgpkX
6P3y3FnvQGgrEamyx9bpciWfifRVxSzC4E5irDY/RJDoKurrfxaG9hWHnBIo
+CW4DVkcGkmPdtbAmUHxd9gkfglKDSjaFA6Jjc45iMQhbn0LMYoMKOAFT5Rf
1hGV3lLCHpOcgeehgG2DXrGUqHT1rKnsQHmB70pQByLqVrrzgniUrIpc57wC
og3R/UaFYAsyWolm+rEnfXnQnBPEXdGnjD8Gv4zjXWxpD+9yIJhiCTIkefka
mqLzPCMNQKQEQzvrLp6hewxQSfrmm2bYjUwyijq2ymihg7egu7wJqPa2ZpJn
9Bu5G9VxuxecikUUNRaPkGcRT+AEs+vDxw273qB2q3FVi/qZaVWUMmzcDziC
Lav0YVVhAaz0pD9csnGfI15M3TySeRMLa2LtOB53Fo807mfvdIkBv40H/Mzq
j94zlto4poN3TU68OdbTyCty76KtCTrjRIYKs3ZDFlKpx0BYrsWv/zzbx2xs
jgV/RwB+pZbc7x2MdQS/Cc1H8wjRpzVS8zzUPCeWPtov//8CTwy08PY1Wkuq
T2J0LZGTQB3OP+Pr7R487ReUQZ2r9nef17QArntEKWMiuiPqcDwVXrIVLZX1
UFnYajvxcmYDb//E1CendZbHXfSIjnxnsziFDJmp+MXf3rr+oDInTfVLreNE
RQXU6xM/Kadge7ZdvnKovFQ0LtwmMTailMtrFJFN+U7uItyYObEPb1eK9jAj
0eRiMr3za1MKMI2DmNNAIHNt4bFAF1KHBPI1id62PE4/VQaKnDABRSjkB06D
uVHA6SMqg6vklCsoSzemXX7tkEZsel4gqKr8vCXY5L8jQY0MdEy1AW/vhVRb
RBFH552gABtY3YOgkjiZ5Rp3Ai4v8+30KFDdzcw1Cjj05FlQIBtEdNTUKiww
oNUDCSipAAkyEmMA/jY8pPKc86BOc+9d6W+H5RyHXrgjQyQT

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzev1VU8OeBWlBW9JcJLFnXkhTYtGubC62WRyRA82II7bJC1tB/phKemwn3wgnvX+YuIK9Bk7zpkWG4Dmog+Mp8c85M3Gpjk73KvZ/IO2i43f2l2bpxGvErPGNm9cvK73McrxMaxInRbzOseTCnUVfhzKJDh1GJ30B7dT1+Ok39dYz/JicrN3038ROLnacoHLPFsG2Msr/rpagFPevXEWmSWcMjiS3FpTbNiQa8neKlM8KsZwIUMSS1BzNuXQzV/bLhc9nYjFeE4T3zWlxjZ89A4d+jUCi/SngXy2CE+JpBJwvWyP0dbaHhUa/6OtuqqFCax3usrNEH2ZAnTV94OqmMZUSqxQgWwkb/RQgF1CT4h2W6nLTdIhOoAZm14pefmZmjeg5HT+ax2GHDMKa83rqPmbC6mlLcKOD+5kHN3t4QeClgRjQ4nVokkO7EkaL2evdfRiKfkmfCD0awpA8lHqfGd5EW+lWcawbX4OB3fGm1o/LQHLjqxkEoRXav0RpLZPkVA17zPFzBsDw1a2/r0HyWn5c9aEbEG+8YhYFQ2AeQyW8k0vAOMR0yU5ik+0OSd8oEM4RniQR6zuH3fp27NTwBxVuC3leMvWfA1Q04vDm/AQ6WIB/+eanc09Tj5XFUSeOB+QaIT79NLM5+mGcOPL6PqomzMY2Y64UaYsjI/CmJaFNzMvyrLYTTVnfL/hHWY0Ofl4rBOI9FHLgqlVjnAdQ8qYI2PfHEsayFGGqDues7cU2xmVBsHn2cPKNRQam9+WwK3b1eBb2NNOvP6ZeTAtH0R"
`endif