// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
W49ewJRc2Fiu3serFgCa7Rzv8Y+G7VNVYZ7syPYwVCCiPNRM2LmsLBIcBg4G
SSDoBzlFkDycvNfVxXGq5cCYyx+mpBhm4iAvfXiljjnUGEXpuMcISpzWelfi
rX7CONtxQrRdnpo/z4JA7O8zN+xhKAnqhsLFj5dU9U29/he3DVY50C2Ef0E5
0jtyc8qGUOxsrm5MXr+3Cb1/HUnhCkjk0KNsoYeAiX5OmrhiGHKkrZibgCCE
xGeB6skxjHno4nwEO3p4g9/hy+O/VYqJoNwtA6cyppPW+GfHOQ0VG4aKylhp
L3ztJmpDhA/buP0FUuQRpcI1cLUKhJOgppXyt1E9wA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
K0bgp/JbiRguTUtO/zqH8mGBpekpIULVtyyRGmKzVpqx1N+PMnJ0ARCDZxkf
7hb6fl/apnMppXXwKFXpQugTfYfI/j5R8jR7Qp5fhyh3cLcpMgnqgMoQg+2S
kqwsocEwZGPlAlrqyv6XbDs5vjgIPRjEmyPMVJVDhKRQRZZZF6WnOCkbzhOU
QpNySNTJc+IFGsWL9JsDgFaGMSd1wGgHOih9Rzt4DrEjyElRqBhpW6uYnj5g
iG14swFcA3F4i+/lcBUHF6bfEqfgiBE4T9DwjgSEaJX/+nufiuJosc7LYrCB
cBe5eMj9ZZGWNW4PE1e6mUcFgApz0CUVHG6HD4s4Ew==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oWNmtVGpwGNoI8Ef88SLl/q3uD2yiHIYmMCieyyDyOCTjaJriVAohWN9pVHa
SNUsNAxdwxH7xWFQYW++4jbxmAOojBRhtniZ8sGDRp9q5vHEEahSQ9z4a9C8
ZX6VWz9D8BL91XUkvFSx2sjCodnnCG56950zi0fxxoI/wPoqZAxFJiLFkDA1
ZVJIkjJH5xVVKYJvgp43blSjLbniC+fSN8P3+1RkGw8DqQtCDohYKB+4wnXD
oZFWBoD/QVZwhpUhux0y7jIe05ySHjAqItsWiqNNplJb4SUjREUZ4dfDAFR2
GhZ6qU/g+FUjWReEE6kz5W1klJ3OYQ24mb5qg5nlBA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
U1ThGv+9uwF2bRl583iU3KbeOAvfmAeYhzMe2+6cC5YUfzyUjEdMujxsoPDx
TdjAx6W9EnpTlZqv5ZR6vaw0BOaCCLyJpVDa1gzz8tn9OUZP49ZsRCW749TW
QuPNEAyEADhbJXYeI59yHuXZrdHD/7c/5IA/m5+uUJ5RlJVLdVW5dc+F1IAM
3x/kUwfPiuDTP0QRAIg1gYDmIOhQix1Uaecvz+s+plkBwRd3ZCLy0WSqgcAZ
MIAIRXlTBhJab/JiozY2kJU2pwUnqIz8tGsusaUh1/8EE9Z75riES6p2YpOF
RyagR4nBVJFVMvpg+kMRk0+RO4KCjSpClanCJXzfaQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oolGmlngBHTa+DY/MXd2IvJVXv+vl18t9eTnJRa4stRdxreRZutnuOpfovtc
4VPBvb/EHAEqUF05T6+wg8UzEZDmUQJrE/+Z5LWg8bNY4O6DVwFBlANRsbWm
VVF3+uigdMJ6PrtAM5M4P59z33p7QU9EBnNdXHLhekh36JCcKBQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ma1vXhxUx8PNqMITo+ZwwJ3JPm0VAq1O9SBH3Gus4J72JTBVRCug3EWHLZ9w
2SLcihAMGPIn3/UBrnrQ/W0RI/cIo4mcbG24j3q41g1a1Fe0SmGL158hJfUC
1I7cWEqDXs4Zh+F90NBrJRZNIorac3L4Et+l+Ka7YvuerPEj5Z0Jx2tUf8+/
evcINSHk9x8EcsiNq9cAgXW3k/vzv1fzMGmh/fDi1sA8NV2Fl2UFFW8maxwM
wn4cDIRmAT1hc9BDl3qsWFBHfDnvu1nFRdi3QfEA+5R4q+KqPIxb9OoxeIm4
IHVKwqIqgeS2SE5kr2Z6Bf6QzabLMz5U6aXtckBaOZn4hSanK1hY1lUVzC2r
bJpocUeIDh29QbaFDB0KbUMrSxVb409p4bvuKrXfqhcjpH+n8TgOUcwOuMiv
gU3CIGMarEVDkt3tY7nLXr/UEWlgzmMEJsK4rLq8yc+QqFOMos8EOlCCt7qo
o+5LTAU4qeW+6gskd62JdzGIfpS7WZC5


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uI4FvkIx5ZLxXdqnpMKOLHhCKcMwBBfmw/S+dgBdsw6m5oadCzinyeKrqK9N
o0fhy5aCgBvaP4k8BxViRtxzGq8yCKzgrmxcX/OGnrvoBnhCezikPQnGxG5i
6L/qYwDx3uADXd4/zqMxDxQBzaYELPQPTK8TwG7SdNeO/atfzaY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pwMa/tFnlgD6llV0iYfTwOQFs9WeFPEWqCfO6cOSMZ+6N4kW6R/5hb9xxM/h
GarKevFtgMuISz2Y5EQb8UelOId1ln/Ze74YLDIPSbOphFijs0Z2vPKfx3m7
a4HX6kfjnl8W9JpWSa9X2I16GY/aklHI0ugvWDG+m6m4kF+3BXU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 217824)
`pragma protect data_block
NJtNJkyIO2bL3svMGQ3lVV5eqouw9FrAiGrfQywrdd6KBWVP/4AsCxSEXqyn
+rJYJGOE3P15b1EuG2DlNqNwYBtxoWiUC1W68SBnmjSXT94M0NyBYHAHD5/e
QV69HgZbvk8aj7QvzNERarWtVNSGOeaVb5RfBanQbaUjDo1FFrh/Xc8F1jhF
kaeLpzobAZZs2n+wT9BIBXAY1sodjZ0q2xzDXmcusc8NGjKtoZ6kxrghebog
GbJqVuGql5NtLWDUyR7MDyfInXlX4DqL6CPsTdGIhJIeVSBJgDFM2QAIrH6m
ew0Z608F2eWEMB/45iK3V8wQOWVJExTxmvuvSe4Ur0ViMIJRIptDHHwVIGLq
Lvpuqd3lCCbXsdqJMnPRFQKVNck3xUJbXb0UojPLePsetLU8n0wB1LC+kizS
YjQzsT+Kqn1U/Fdy6PqW+dw/XHLEIOn8VMJBlx6UaOCjORkT2XHx8Ka7gsyt
kTlN4toTQvCR4/7IviWA9MNfMz/S1xcHWUdpYSdGtMMrzhVcP27OmIsofqfC
ch4I2ev8CB+qKoecogJxVvMfTmFCedzbr1wNvUm2L9IC2lKdOlmQBx03gHI0
aFQuQvGZh6S4+Te5QT/C0KSKXDWyfHuZjQkghIz5ZK9k/nx+NLHCi4T/W+52
sAqSHTHSpFOTtaU4W1HOJR13wpFn/c2CKlYNivR1N2Wzrf5jbODZB4vWouBB
JXEgVXDDxpsFO1qV3UAFeqhviVRbm0ocNw+C71ViSa0hd23pWU6/xBBLVFyv
EdJSEPiAV+KmOjL5Ijmm2g1eDzhjH2wQM3xLV++XE3Nq1gO8BD+BBR6GF6xU
ZRSdYoASeWgXl0c/hf5ROkZBVV00clq7VfJYBsjtVuQ9Awey53u4qDww/xyM
Sy8W7OWKRtLbI8YZaF2d1gGOPqpMNg94UfDICbdD1GeeoD8RxBZSwVzEAIRA
SAx9ElBvdHRaLf7OGvAlfrstkH9Pj1793jOzV4Mm5PqPKOpigau1J1+fKWf2
ajeQ6YCq7NQ8bsbWxkWXEqR0XduI5nee9wAPn2YO+IcwHOV0rxHHFa5ehwMb
TfoENUS9juJNG/PsKcGmd8+s9XLJkMjtdjk8gssV2inHpd6lTRZWq0784O8h
/TbFRRFBNEroBgg3mMe6DON6AJM6WswyaeD+2rbwsLkfIcJlaCdJTblxnVmi
wd76FOOjk00h+E5nkhCQGR378jaIAoo4ucrPXJChmIJi4tOiA/azDFDfpkRl
C5DyI75BY+0EAY4owAwtf1WnMz/FJSG2Oy4nyZwRHd7ko7pEMTmp2lIs15Rb
pter72j5Wrqjr99k3YiMP6VcrdD9h81mXtQOfjKVWkMAhVRdosdhKhY6X+P6
wv7tidvxjWd9LH3G0gBX3IWfdRLnIbI6V0B3d2Hw2Fts8L/JQPbDCxcK9NGS
Zr6vqsyeU/4C4pdRfSUND6q9fJo09UqaahhRoEIiWHYNjF8mruWbY/VvvLmq
pyV57/A+qToVu8BVghHlgISUW1lLM9UDn6M7DTseaQQtW5rUNC4b2SYC5Fvb
jVlADFKyoYFPp4I4PHcyGwEg+c9nSaxfFFPRyD6/t2OPICmZ+7dFbJWBbJ1u
jZLOpcWmop8COQ1lxGo2FQoDc/I6Y2v6s410uA4tbRzfxMJGFJR6JCJBiO/a
Q8u3oU5DG8YjjuwBMBd+ALiJwEoUpf9WnjwPRCwZWdDEvnUU2B2Y0CWY9GEV
f5WR6/muIqx6eDZU5Ye8jMsgjnhr9MA2wkbY8Zp1UYpc1Os2sVbigyneTPB4
4zpyZp9M1aNedKnASKWUS7ojQL/rHl36S+PCWIEe5OG5+21UFw/qxIdcCxAV
Y4yqHLl+YYuFe77Ky1YBau+RokmwzHMNDrZrtZkzqU9oFASXIWU4ePOZUaqn
npLOZi3f3rRBZmk5r2MrOf63anahWZRK/LnjFCgSM8rRltvyjs2ClnUNHCpl
fHJHZN0GVAz/Yxcn3S3G1lpJZKLLt+Cv/700MtY0f7kY/rPHs9F/1I0JuamE
+jHtD0QO3caXcRJACzBifAs6W0r9EOSJ2lG1lXW8cktOfW/4kMtJ4TKFMN9e
yirhc8aiUi/UeBRRJvzHwO7/ye/o2nCvn4eY2KIbzL7pRaGo1Bvd0TPuaRlM
N5Ji5L5G+qI75ga1T6k/3kQkV/kapItcXKICBrOlKB5etBPS5/HcobBtmhGo
JnYVUKG6oZoICIBjrkEdhwH1Jg7d2nVQ21aZfNFSJvQczHRz8LQI3+jU4F8O
RDdZaptHs8xu75cIIpYnrxW2NRlWVehj/j+tTnf4YH50YwWrk2Xs+3ariLhV
B/Brt2JSAVyF/eegqYPzP8qoxvlCxWh9iGJLYL7LbfbE1Z3rdQuDaWELWrcR
J2xTvocHZXXHLk/7cMqrT4Q07B+Kbv41rwCY3t9fLm/G3KBuTZRjAkdFgMMn
G52j6SZU5ZcFFQs8XJET0QxAIdL5uBtfUquzdLXOFCNIn3al8+hesb6y+CTZ
bvYvKh+dZsaH7xNa3sRhLBNL95v3dsh1H3kZM1rTJmhIktGx10x7GGI6mdBf
RR7Fd77uoh42hhAgKpbpV0FflI5YHiZdAFA61hn/dgDBBWScX5rBLCxUQmUt
2oSLk6sUN2wIomV28XjzXMieaCwNZGG2I8PlhX/noxWC9WUz6mXxxVMz/05H
AvWnYl4ak4mkE01lPTEF+yXRr+dzFMbvMV3e6DsTEp1etoLOfHrmYN7S5nKc
uHfQ0ivIgWOP+DqAKp2G/N36iX5KCC6fe6N9QWH0iOENvTOKqtMALCYkFB3j
6/wUMrr6JFTlijLH55oBmEzwlvDclpre4zQeHr/SBMWcKRFWIfDVPQTjwkay
jX/Y/N7nR3SC9Qa/8VeYE/eDLBGuBpeMmbCB8B9QTmOKOWxY9Tf5727SdBWM
p2ckQHYWgTXp6FW/V6vMM/+zusp2SpQBpOPaNRZxIJEE4CeW49UCYM8jd29N
60S9gTGleKBDtCkefjzIPI9e7xCH7hiB4lgyC7LUqF77+zg4pC+/x2upPnDF
KBz8bS6IVf4GDK5SGl/c0t92nrzMiw6gZk1yBO6/Swajn4fEDd8AGsfCTyEe
tSigVvO25BzR08UoqAAOGAgVZ4hjuBw1zZQUfzUmF4HGbhtwnpH+LfDuOS5w
PGjS0L/MwVXGnLzh2baM85B/EDrPrkkW933BJPk4syv5ynT0zT120NhbPaJe
IugJK8iUswUFDTyAyF5fnq0r63tIvHdIA5BGnOyj9WqsdaoHmHtUatLMZZEC
ZG/scp2w5IJ6fe3qpwGzDXe3IIOlNWFI4Mqxm3Du+oL2IbTw20itiBKAvBai
caTzRICUSGBDaAbDS0mp7i7P9j4zqiFJskn9pqSaCEb9Fkse9ixNTMrvswmz
Lx9C4IwyBBgT0oo5G9C0PDB6F4i6RS/inteTIdfPqlXk+L7cmkLUU4wrBoNm
dZAE9zrUo0qGEq37TkvlmSnPpYphxXSrmHTIiT7F6okYHRXT/yV59uWNod8C
Uc2WshSB5qC4whTkUKsrjrfVeQt4uMkbWjjU0Y38OX1PMsHUVSxtpaYaQBSm
bJHflFMWUVAa6qIi1116LyE5OdZu5LPQzjklm4Nm+CZlhb4OzTNfDlDz7OuE
HO9JQnH9SpAHTeZX31968MKyYs0KhvMjC+jPrLYuUxPPz5qm6NDCZimcMF7I
oAD7wD3si8RT3nmNUIwpt/lODoe0+Qq1cw8g43LXY/6+4w/gIdXcoX9ctmJ5
sU4MQ5iz82XQRY3SORVtMyNSG53JvJ8JkxKqfH9NOpVAlM5D7FS7XWcO/Azb
7Y/PC1MrN1ci/7N6eNPQdIuq9gDZNvQB6bm8bjfe0kGxLizqwHXkhX/tL3iq
C051QjX/kZVKdClh82w2zSluh3ERqehQ8R685OEmejJNoo1P8Kz1eD/SyzN2
wikMHSkRIsAMS28JSaU2H/0RYEM8pC36JOjyCN2LVfJHY+oxvOdRpTHWBWC/
fa1FxDOuzNp2R4jI1LaRPuvalK07YSCOLMsgZp/Vc+Corm/y6WbHjwVKPqo/
9IxKQMYOJrpToWTNPiZxHn4EvnMcMLopvkFZ6YGPCTM0bHf3dBUgbfBXAmWT
OMvX3uUVdeQJSdwtKYZ9wfH18NPh03bEj0SJ0CGZwo7j8c42yNKbhpGGzITY
xbpd2SwykcnPwR1YgGZ0B/vwRcKJOZqHWxxoez7K0jNbvKUFSmN9BwdkakYH
SSov8CNbphS6aw76AYKS0onru21X1aXhncu44Gbc2/eBtmLuj3fY0APFrg2L
u1R4W4CJI68IXiJ7dRhczcCgofpuskE1iNjmBqgY1QT2yK8tbQNXt+aup9t7
bO1sJFdEgtMAfLsJK+SsllVARDyCEjSItDl7zahn5uiZ5zenPCqe6JikIrTj
ubxJgj430pI2WGNoLDMjZqy3eeE6DbmDn4s/ehoZEkM886cdpuJMtt8tkLkn
h7vPxFkzecR0PbautYqI13rDmp1H0MZEaI6biY05yHi53Gp2uhVDMmYSZ/Jd
NosAE55MXCSDvoCGZQMn/+S0JUz1sbN/k/qADJKPb0vYJsKKn1gvtnyWLeLU
8cNgjk5q09hQ7L8Y6uhjpYF1wPnlzBRnLLFFerLemAPO2S7oz6b8CIxXWLpN
zHrAjmgcBmdlg4nQasrtoZ2e5W91AkFme6+mKpzBzpNdIio8G735BXaSdg4l
w0NWaEktgkOSRXQbu3MUeE0v9T4VUqOXHA8RjLTszuDn9bxb8I9wgSxvcRJQ
mk7ThoCNHC/7QoZFO7lHTei2y5Wxt2AWOmPVh1xQcIxLZVFPSJ+B9bzmQggq
zvPf4YIIqDKS5DOX/dKsnCwngxhKMKCKZ3O3KsXntZBbsrqqSIJKkbb4D5ox
ongbp/ZySyK2uFxIpyBFVubKlIOWpo0ucq56U0kQ6IcRGAAMx9GRA4hrgx02
JckaNgDH9CJFlwtlZuRq4UisZauGqUejwsbYbk9AN+J9XuLLi2LJvcKURx23
SAHgnffb/MTJgOGmxz5xyS3lty651FbCXhCzASIGPQ1aCe89DGRhtU/aIhDb
CbTU8AqgcqiSWDdWh+36yV+fADT2jTr+PXrVKVO54WfX5DdQGmxQ0XnbnF1p
uWuCMkf/5FwgJKkM19nGHln3KnNA7N2YQ7MpolxFyZxg2ibwwS8FJVLkUaru
H51P8YV402Uw5ZHOTFwj53zqdtDRqmZTyjhnSSovLJ6J2lWMVafb5Zdx54Gv
ZAbOLWhQkUDtEuLQVefSkHgpLTjFqUFSdnuL8VrkKPUMx76qzbUcpwVUXLJJ
oVMh21H0+2XrxC5ULP07EMMcKQ3jCuU1BbUSHTe+vdKIg354HwXjjvUZa0mv
TYNSUHQOdLXja9UDrbpcJ1IOMLApqssBcBddn8TxN0bWLFQZCRLRPu3pV66U
TJRrb1q6aybGf2lzDpSUOazM/ZO5BLw5pTs0Oc2m86yAhjWEoa1mehNN8pLA
n1h8uf+i7B4czxj7gbxlt84gYbTUSfdYEzyfQqGOTKWY7IEOz2M9+6pialyv
QsLAPckrvIjzQwOSl4PA5ZkwInSqvmYkbWIUxVPXC9yeRYPyXMBy3dUVZmLL
1yGcCDPUWcT+a8xN5rVEhMPQPwcn7KjmZAAGAw8I2cCewIcHCOQy1RbBxFTq
bZEjgMZzfmlC9WHWNE4OUP7lLd3xU41+kXXsp80vEnrwOOGuwVVkEbtGe8I/
b8V1/9Om+onGadL3MEjk8OH4xdaPGDSWM1IMDUMOS/vKpW+mD3oV1VKJo18p
qKkUpRteQ+ZCasr9Q5iPotB8rE99SIUbvwz9d69tutCr5izLE2F3Ay8mRPSi
viMFLDotO2GhvTbFWvi/M6SoO5eQj6o6EG4QfI/Xv+O1+mjSCHrSuAdMgAUp
SjvZGUnJs4QX5Z12WiZNZI1aFSgDr0uNwOPN1PfdyTptGDLjsqTSKNrotuv/
LvXu9+P6l8F0MwUnEI7KjQbMHDYD6sWVRMxCKHVo8YnzpkqFfcATL7R7Nf3+
QSxl92gna7gYTi4tOvTg7JkoOjBEGl1pYASMyTHjQpo5X0jYBVnDx771DqeZ
A35euHKNtmdaUXfsjZ0BBRqId4zS9zsVPvAHAOHjrCp/kj11Rdk0h+HSU2XU
DD/7I1u20mMgL78U5AauVmvc2dzCQsWYF07ylcWm4sT1z8tKvI5mKYH++jR5
SunZ85w2IgtwOGW5x+EUmOcN3CQJjVZmDL6fkZ0hEz6fZXkgrbdti5HUrY3k
YhNe1A5xNtSC7aQUg8wdFZhJZ21F/g0jYNEgXy8fxE0i91kO/0W3weGP/Eno
4/XmBBK3ntwTSkB4NH3Ndmb3bGE8auPFLrYuerWNkRVVIFSpXYlhZOuqXcLH
WDADlIrCM9xecTASG2i9oieyijUeN+kIhwdFs3cqMJVra4QkpTW55yhllPpD
6/ryOZRLxbSJqvc4hCGmZnJOqJ2sfAGYW1kX2D5gpL1/jMSz4YPRCEuxHbCU
i6kvRxGg4TNP832RQ3ILEndbw7G3ragTSevW56O/vLl/DIYk8tBeCgUdixot
Gfi57FeutA7dDC021pTGujXWcV0cjH9Gs8I3WADRNm2e8Jmqtf4+VJKTG/+0
+s5E7B5N4v7gKHTwz20c179v4ERLzvG7HhmBThKU2H5ziqomtHt7WZIk4tek
FCuw3PXZfwgT+niipu3Y4pFa86sVN+rF/JMSneN+GONWIA6Qx+o8TOO7yjsy
P+bX9MNlaQegflQoPrLUYANKEUH5kaPKD1Vu09B+cJZlayWUHwlH7+iczKeD
ERwMHMSoBN3T0dZu8NpOWzzIjHK7wEVeph5/tV830Qh2v/+UD46YAPHjget0
LrTGSI/e8bqVvSjMecHxX9N4RUUvQu8fg4awzM7lNpPJHVmnHg0m/a9MnsMh
zHh+2pmyOkyXofloYVEYRtsVLwptSQ03lQu8rluZJpJ4uvZeiu6kL+FqB1Y4
e/hcZa/Ttz9RgMOA7hjvG/cvHvxa2smc+XQi21CHKN7HxsiG6YE3xG3hyft0
c0yqGiuRyLBq7ejlQSPAw9HnWWaAS0BwoF0599dfymIRHxroV9BFJuWfQgnD
35GcV4YOpy7/rnH3nRkftyf+cz7M2kxfTpU3B0BmTEfrabz/ZNM6LSUIueW0
Se4YuQp7C8XYr1GDElX0bDom7HPdl7MwmbUnMxO1VQncDocYVl067+OzKK4H
SK7urMTM+B3WSY49nWPrXvcss4iChNO+beK6sC3Y/u6/lk35vRh0BUPiRDli
UdpspnF0AkDFURLKYoMqC/hAQcAbPmbQwO0Yw7GcVtLRY3nEFa7a5/opOTwM
JiBKiRjkIqn+9wis0lwXJfwHGVppFrbkHgRr0NQy0EtoU2lkDmCVH+br3ECd
8BmcPb1NyKafERELQS2ZWESqBJ0yijEj0Tu78yXlcsrx8EEnvtAuFP9u4Nz7
hvjOIyIDTTGjUsEVOzSaL7pLGOm4E6vmKmxE+fx/3hYVCRIoyi2qCwH8Hngk
K5TAS7qEaptpiVqs2H74vNms3nGPd/aajyK53ivy+0EJL6dqlcsV16XcZe6z
UPWGGk6e5L2Qv65OGrxIj9TLI+DJTu3p27dFSLB/oHLnoM4nbSnpnXjiHHsN
b7hqKrWmjRduQ5fQMWTf0GpW1UGDCDWQeoumVNmN39lR952waoo2rE0lvq5d
xtvJt51KbCT4A6yywqwp4FiNyaEIa+iFXSFSZ+ICRadrG9JxA1OBSTj1gb9b
5AAAuV8j1t+FMPH1XhpV6sg1+EQDnL8q1p/BCJkgtrpQmSK4c3LD4ckaCYyj
YzRqUPgCE7TyiaPqcYSvACGJslQwuRNYV9mQsU9Z8YQcqDFQzFdFfMyKXdvz
OAlfunOIYtDoWdgGZIlZdtPFxv/b07t+rCWuGqjjkM4c1u9JriU9Xt5LuNHI
58Y8YB1LlNbH6pLCQOJjGCAM6gruuVdNKg564DiBtRDdmIDss12uYfYMk3bY
brInrrQxGMHVW1j6sHsivmml1NQLMma2WXKKYl3NNr6iglSL54dTY/Cf+MEU
RGAZWLxG/51LD6xHfgzCmh1e0RX9dN9Fhu87d6RwvoBmAip8xYPw4k+Rdofy
G4XRHdr/j5Hqh1X7L0EA78uET/eY42VNGT6yAV5xVlHkyW09xvA6XrRonJfa
0bhdLer+np0ibJ1i+5DIRWpyZy/hDv/4NFnXr2NnEH59gx/67qFEmXUNu+yS
rkC+7gDjvHl/6hPOpAJmWz/y7nb0hHIkLSyfl1IOgQQ7jcM8HNalkGLbTSWh
GHaeVA6NE1QOLsHFJPoboQU+V6krn9I5h8Eboqv+lAis3TwQDogNDPxuCD+/
ld4PJ25h7ECt0qsB7C1dh+CrVoJpy/NPL+S9Yo+ZWTHn47cxNwI+3NVHqkdb
252HvC9/6kzLCubms7HYkxqmDfjVPx67pcrNlVqo+uSHQz5McvulyJP1L6zH
wcKWlF7Aqvk2PQJER/n/xlBlO5anjuqvx3jJpv8Nuc7C9KRaTilN0bWfb/dr
eK8eC/nHvJjGIe+sLdVP9NFWLbzbO3C0SM+7Ow2X3NCm3ponSfjicYGOlknU
Latg1nMe85AYgcUgIDAwzrz1qQXaxT2R3t2OWzI2px3bWmZpemnKtH3FtBCo
vfSp4SJYGXDd+sJEMC9FI8OmbwxId+rUV/6o/BvdjieiUepZGLfX8aRZ35Mr
vh7imNoZ18HDZYMIV0XZjhdPGPJHM8gtOWKkG/Ntilee6tYi/UUuCNZPaXge
jXMRC4pISUOkP/t/XY5V5j57kOndEcSY8IBm1SXpWD/uO40qoa9FKHi1lDam
pUlwuiAkOhIbBc+Neumu4IJ2NZE8oeweStyZN/tjHA2n2FnZ60Tqe37GNXJP
NhgiF8RJY1fjUxd7xcRwPrkDknnjNqL9z9HfgGWNiME7veZj1VLXRGFJissU
FGcpf31nqVCROXP/SkyMmwDMGFWnfYewgiWxTPJ5rJXb7G4Jxf0zV+nF5n1z
WoW+fPUi/W5zjqOtLsFJeSCaUHBEEOZrlQNHOKBiR38OHwkblptKESwQNXLR
I0y/uqlVaELgP5sbshgIhZnSPwp4EzQhzRZhJGdL7KEas1FbEuRZt9sTfR3P
Vf2/tsByJsVpgOQSQxvWPW7qqI+mmd5+sFIi/kfA/iNGwnwHUu8+IU+TTbwq
zGkW5H3yT3jySevDgHxh5FSFo8V5xaps9vE3a2jcm+b+0Nf1WMSh1ywn3vdZ
wHcfLArnsBpgL9bZ6mByJ4TukfDJvgT1if3dwCxBFSrNE6sYIFEg824qLeH3
/WXvlGs0X1NBWQWt3g8Kq2T8VcknyUrDrzrh1vszT6xK52YicXgG+RHJQlUN
MIw62NaBMdaHyuZdiqZnM/I7doEoGNXyvR8yODcKaUQ6xynhOjXup5tAAEk2
7C/JQbCipvDSS7RqXk9uQIV1jVNALvgApxGDJqashsevh+AG8l+/JiV0QV0u
sRYym4bl6xAuTA15pYd4uggH6UiJPGlrRB7E672X73zXT3EcntVbOukWsEIs
vafeAhTvFhRnG1ubh9eeFEMUX79uCXORhUbBTLP8kfdU+5vXv8KlXYH6ImA7
7oYqluG+i9bnRvFyTBRddQ1kr+3t3c0oqs3PmYt0Uk5rc3UWq2QaBIf7Nv/h
wo/AiNla9ihEJx9pLMza9ixll67QmUi1xCWKRDybA1HSQvufxL1qvbHdkwyh
AY8NGb4w4vuoUmBCUkMSiR6k5BbHUkFNQqnJ13BN4w4iGlFjLvxJcX6DCF67
I2ABJb1vWGcjQhDS1YoJbHSoRstPS78AjTQwpOe2CRW5OkiJYQUI6NiL66Ix
uFzv8AyF5xL4stFVZ9VlTr+C/BzpamOD+4ibmNwGDVasJhDwgageCwAfwLK6
E6lvb/RS5/WRPcWr5ZcNcu0Pcm2YX41VCjkLwqO12dFF+4elZg6hW4srTM29
tNelzRKQyHbxCqaZ4vRki8n96xj8UgTp5cwsHhrR87wdkJbZ7hdnDt7WmSxX
0HXsOMqj0h2W7e7zhsXgLPL0ANVYJVRdaL8saFjcA2FbysCyE1FCcmDXcITf
YUltL9jxtNR79aLpM/GacnqwHR+TVZaSQP5DjpIP0o3xI3Tm73bHXNgOmcB8
swlorPF1UR2hhR+gaQNcGA3fQQU4CdS234cPMZJ4lRLe43eHp32JWaED3DRL
RIf6jzhAEN3f+gD1K6lscycnR44w7f/EBZe3gkESIROhFH+Q5kfKxn9lQz1R
zrVY0NcZLu62Xg5S/w1CxCKD4t6ETg3pOJDMuP7k5Z25r2+LC+KTjUinhVGb
TIbwFwzPExaJs+tYqavz3W1MPMZ99flm0d50YP7ogai8SW9zxGul4c36QOwJ
fIronfvUkgK2MEk4lti8p2KWyjwNkblAG1+7FUhL7tZWOjkgWpimt0bjPorl
AgIzp4NrUO7orkidB5LfDhJWClT/efdu2qxyvY3ZlbGnYUdgb9OnP8g43uuD
1B5QGbPGYnY9GWzzy1DADMa91luljOcOZNetRQZJIEFSgLMu7vFz0S6lqGSW
QH+YgwoNVf09yEKLfxSS7lBw3/VMdE8ClvXB3TL3ytEgYGYck143ZEKHXf1a
RG/rLuFUHU9QUEVpa6UwjxZUty1qe2qQw0tR1vlu9P2144Er4jRrn7M7AMkv
/ZhhmnuFLOnq/ZmF497qMXRUkk7l1sgqX7DGTbiggkPwsoJh56/SpJJlh1/r
pnVJx4KOZ4PGhewgjlt1DeNAo1eYoUucscd8pLAyWlGU8SapABg9eaFP+xEW
6+CP8NnYMeRkDKr8RXpLao9JAuRVpr9HTESk/AalzieHfnachC6PeLklgxjx
+JoKonlX0Q1bUoRtPbLBeJY3fK9r5YHbUpKE8oHUYh8PLLgn+XdAifZPOT0O
RVHZ6BX4Ni7vWEDAYIYJ7gvxsLAiKld9CAbqMcYlUzY7gCSSm+TjYlGZJYmi
NozVoyHken+pl3t3cyGPdtGEZQTI0l/oJYe+eXRapDPev+tKabd9p8/rl/oe
w9pX97B24i+notSXp1KejyB7CBLBC3Wt8xUQXizNGYffrL6a/yQMm5TFRsRh
OkEVZ5nM3wbClWsstL7sHEbxlLbjjfb0f2BPsBIclVyTWSk9M2aweR4jj0Nd
oJG0c1xMhPfdN+KIZuxtz04sfnyVTzxtbfcidMv5xH60Y3Pz4jnchqSxHwyn
5slOpMcUYGLhhBnqT0+Vbdv9b72sTwd6hs1YYvwCR8Rkz5dil3xNFN03ZKZ0
RuIKzmMsPfaDy0P8VMET1dTwTeW/hI3/PRJczrn2zXB6xUnXPwLtbYP3v9KV
cK64inmO7Gf478/uXMCWCAvlrz8HjVa8FVCDyzVjcLK8zj/t/M+e3OZDvQ/K
/Gq8k1oWEU7Lk+qcFrNGn2iMmDzDjeKT7gj8f1Fn8zNtdK36jiXc2c0lzyk8
+7rskWzDBn/UJXtvrMVtbqCMkSiiw9bfbpo7CNazrXaWDy8dcCGy+eS/LPUO
NfJUCrMhYYBq7eOd/Iyt7kD12pISzfvFrWUHPSPEpqAAd1IgsI726E3g7f5u
fG8ijZoydGcU1RjQYQDf2yGEwcJFwoCkjTCfZEgb6Nj/rbBdL2Gn1oyY1a7L
FmF2t5xRFS160gEyPxc930Stx4dQqnsAPXfHEzCNsMirErUGmMVkYVNTC0Of
o9npSF6pWMbAouXjffH6lyylxx5ghcy21NPkg94m+zLzi5fJJKYN4PSibNUR
tfVxHyTG5tvbSXhqQePqs1KvBqt7dDxjpmavO+5eh31Eu0oOPqyTedXhMP76
43+bxV5uhupio3lfwajUj2UyjgVSCYoYT/vWFYXjBkkGBGjsTwpWfBtSUsvW
Ftw9Gq2U9gYp/3FTRSYMpAupyVcsWnBQMzSPRg7WpFOwlaQrZYMz9L/gZPil
bseRjdRSHNdkrAolaa8RW1YJmpYjrp9HZm+4nA3XHiGp6GEdpKTabWE/eCQd
dCNma70chbiK0ZvTXWRll5NGKojcBITCtQ96pDOLBLN9YyUafQewH9wjHoVF
05uuc0CZWwmSCf2Xo9cbBvCv7KSUs97vNnjIS8eXpaNBnS2RJSM+z/Ca8Rqb
lsILyJ7sYTYEQNVhok55emWvWzpEu8ltTN79LZgxtzqkSaxjP0WOOR89eF70
n36mnyKuqcic876E3EIkBVIfQhITjTsCcTvlK0F1f4/P3Fgycow4pNTmwemW
0EV+b+WIDvp08gW1haI6NlGMOuDzldFEqio6J3LXxZqu8Wt8XP6HgwAKuj2b
U00UN9pdCEcUWMI3Y5dt8Kka9uVZrzhzgeTLw4KZKnjqbi6+ZDG172RbWDgQ
kdWVEgWU6YIWf0818RBOez34Jqy0x/FOiTxyxh7jZNbm92TxP1FL+9z8aFvn
5wxpx+r5FY5PYdTsWQnieD3zpUxa6a33OwM5UmEoB6UNj/IUff17g6x422cv
S4y+ck13eVU6TYccpO7ztc5HhSyHOIaBNNe9QU5ODnOAPzkHpjc3Oc30QuJ6
olJDBDhXKjecOpiX6gmOmd0FduAKXh4D/OiSjm4IHQsUfjBwpxJHwpkbFqJC
FzRmf6BdpEH4wgxb/vgE4YHFYn2IX83v7ku/g9JVMNsybB4NOAnsFOSD/iDH
C3RK5d0W38qMpBMriJibyTQ1EQYfm/rVEcoJ1ije98iugonO/ga+QQ68Zp8C
VZj07k0GNff9Xyrn35BSAx2QhdnBQQVntZQxAQWYY5PNcIGXbMwhbFaKtu2/
E/xub1BhTUkGtv6JJSJinnAO43WAj75vaDLh3ro80IQrgxqUfKMiW58vJD5w
rmrKYLsvR+AFJFmXJvdAlJM6/bC98XpgqMX1pjzAWJzY9vhn+/vgk8gcvE2c
fG+uRJc7RO8hrDJXOWtTsYyY7oim/lsUJITIOwJx8MW+0jXnZtYNR07pexAZ
Vy0P/GKPspZEgRZOBuYREL581j9/GQtQnsF9jMX7OSs3VEQMat8i74cx9DBd
I7buf8Po2LROUb0+/1eZi8ObcE6n8MgxgViPBbn3wZ+cDDSuugBOucnPjJpn
tHD5ybaJdU9diaHSlEA6G72pbDC7iZYpMrWboAdsxlFQwQfrHwa1mNMRNOvV
6ieTA9zBvzNr0g7Rq3MoYsUmCR/aTMmhV6J7Jj9afLRtRCxKWevLnn0dEgSE
54eJo9sG+mi6VzlPpd1DLP7+g6Vt6D55SwJk4Mp7VG0XgcAsC/b+fzQ2+QDD
b0k1Xrwu8wPvJdHe6snp+rgr1TjAVColTitqycNWdMIrLtNmJXMEyw1D3oRv
TL2PVna1txJB4JOnvacBYjdnvnsuCKR3Xw468CR55gC7ZRzCZCNzfs8FO0pl
FRopI9r+EdCvMsY/iNHinIYDfpTzt4OgcIOepFjLsIzbvLUSQ9BUWoHTr4uv
TxxhLmCGQXxcWyRTxMAcgJc3XhUXPNB+hP5j8R0qMJNhGOJNqBemHHZ6FcyZ
cgPL13oK5qyvh+WgZ2Xe/IL64tvVMXBDYvE5gpQkkLhVNNm2rO1H37MCSQi+
as/2+v2eaf4EJ5BQNSq9JE+c8SLu6fz/ka5FpOdAbqbTNLC9NHlZQ4whkvDH
yd/O7b/y92EtxYAbmjcUGPVQXGHFGwpSZHMmlLhH7ouJCAVjrSQWUnDEzqsM
e6M3338sHLuhTwz//L4MU+lu3b+HKYUbXeC6F3aau3rh8XRgV9ITRzhaIBV4
zns4bnUusEAUBYJxKOm5koI/A2eHWO00DqsPXD0C4D9WWvRw4l+QeyxbXDyO
j3xNAoXkOwda7UKkOTg8Det4V1OhkkqfkAxuqpJOEIEXnlXexFhUHJTF0uLW
NGoSqF/BH+9evM/iXGXeKrO8NKC2IrcdKXwITSzwitJGkSobQMaLzKZEi5zy
/xEP1eIa6/8aHii1aYJEXUM/hPOe4aSGJZucYRN9dw+CTbbhPF4BkVZzqlrb
EJnBKq+FJN7m1kbOiq5rjckaQS6Qqse/nIg6Rc650TRVsMvlGEvaCY86LO2j
vpkXGfc9lc503yOJsahXsvZ+LbpkAoJlk7tgC5Bzc+It8m27UbzKe+3oR3re
SdvzFEwQB263DenBlXjFmM+yEs0ChfwhZu1QTjRbdNavAVEdLmBwe1NkD6gX
2Bd0Z4Xf1FOZuL0bmJYVtQlNCyaXuxGITtDI6SmIqsAcjU8kXYcE1m+Y85b0
KPLOXFwMLMd1pyWGiZjr5Hw3L5ARPnaE/3G0ep35NtTMa5zRoFYon8d8p5YG
RUTp39u1SUF7ScD5S4O1S+QMZMTGAJFAg/VPxzqehyMhWEcMTBuGLHH95lZy
bfZBapTAIQMUh8uQw6p002G9+OCZYWqMOVhGXUffvpNbCx21L9noTQ/JxFLY
N8JGYRDzVkFOQNnBHCf0SDNix2UDUh3P+c6TkkM3DeDN9OVWCIssCr9WpPYl
k2TNWfB5URg9dEtd/45NQwRMiPndE5dbKOvVbAX8y1gYY45nQUItCXUVvFQJ
Iii+20xia8Bg1hQEtj9NIx4X5KBydVLQGyA15GzNQp8OhvA2U3zHEVCISras
WqMnJeo6kaOo5dzjUdYPer2HyOFyRnHHw55qV60eAFsFaOtLwuYBT0A64AAO
xh/XYa6uW6Tk2ndhoYHnxB8bXRRUlTZXfW0XlOCH//heprwvcV6IU0tfnn0E
VVw4siWAX7izLa1mDq73eRQUDKqCxFFL34//lXtO+WlUmQ5SKXG2h6OGjSYp
1AlV2qj4H2AE51vxfCr32wvFBQklP02wWqjVN08yvJfMJJDQpkgp6splzQRS
d0c1SnsRD2qRPH62SKGNxv85u944VtsneleC77nzPS0BuJcB/vIaUfxwecdk
02X8xUQaCLuT0V/GJVnuWrJoS8lTaqd1F3VMes4CQ2Ol/QLy8XBct4sYc+kl
1OV0eZzbM0sxNv/h1H3gZ4Riw+GXBOPVohAKNBLJIYM4BGufeawNwmxJvxFa
14XbB1bNKWiwnT70BParAwnCCLPB3KZPc0gbVA5KkNJe0ZFZFjzRtOzxW4xG
SSN1WgjOlvh0BDAUKVJ1c+LAu3MitDb16uaFMp0Rbi34ThV7WEO8MsqBe4af
74n5gzueyH/UK+7oZeVey4emquV78bpiIpkV2O+ZZPR+C+k7gKGG6caB3FAd
fywgTs5otVbnLDfkzxy9ZfamYpXDZTnlEFwfZKhgRxRMR/EzE8CPR6plIIp+
kaWnyC7D5kmdhoWhNITdUIJcIoGj8q1zHTQbHio2g7AR2VfGzY0F6noI0/u+
orPyQps6fazsZDYM0PHQUIUk7RNvlrOWXwfT8YQp5UmKAmWTbRvLPxi3DX7k
6trGJA2ewzawTu6qN/XjHAZsDYve6Y1jD3GmPEKS3Ry0C+UpLzXabgA5mzaM
uCi0XRVYFc61hreJQ74EefVBPzaeoc7Aei8w86Dx2yCEP44NNy5Q+MQtb7BT
wnCM0QNnJjY0HuUkEV+m+fQdVFxU7wDllgG/PtA9+ijVt6IWYt+VBRvGOK+5
Q4fbjvJik6AmqmXXP2G1qeX7RKJjSRiuLJZ7dC3/B3NYCiSTNWVLMRdnvtrE
HhP4PZPXxTwzwPsxTlcd+cn5MC0vpJvqmaCZQKti8fn5jEsrzfWKd7vrIozO
W1I2YFl4TDO5ktWAYTbyNUeqSvqOHVT6PGYd6bqmSX4YzglGqKj74tVvI6wS
wBekiEigz5+dnLbBBl6/iUuU43qZrDH+kWvLNvyJRoXqK35pnNS00g7+LFKc
w8Jj6unzeGJaFp9lxGhX6CwejBl9Qhy3U3Zkiw2HHy2oRt9aObgJpZsjaZJ2
cKHfV7sSBDr+es4PJSIeCbbZ9ho1RRyMuM7Z9KkKYkJUrY/bVZXiYgxmS9sJ
FHZM3qW9xua6bGXnmd0Gpsup5GcdVyp1/jsntCI/E/bpgdNuf3oD8Ur3/BVH
POg14UIFTU+7KEXCb7O02Cf94D0Uwz29Yf1OjAQAM6NAYvJ5494klhtTu2GW
a1/CZ77HyvkcizZm5EgA3IZ9ekt08GbO9lXl2fsS0uYcKgrBfess+w7XEXgQ
Ctu6q1oTufPkizCkwlB0m+MRtew37qVxyjL6/V0KcT1S3qcmRjEEoJ1zB+rC
t5C6+4KB6OTgMbiDQkSzoXks03FgIi201zr1NtqN121c/B5emI/VA32lrnZP
CY1KmbddFG6kdPKT9cxSvIJm9hn2XBHn6uL5HL5v7LSXnUPDlLa1D1vZGmrY
OJW2qMDJB/GasPCv5r0Hta6KWkOGlyp/olB+/tblpHc7AGJkt1M9Z0VOW04C
xYNZK5b+AODJnqqkzOpEYkPTyU/4kOk3A35xF9QKUZ3/PkI/ZflxaOXNbjk5
GIk42dyatP0BUWYs2cCmgIo9RdgdTC/mi5GgZxRT21XPXFIQmTvyRkXoKe+O
LrTsO5R87Wty3AR+7Xo1WSCAXSTVJA6/Rn2bEOkwwXVeafX9+gFgMQpbPV2k
Dskri6oKblZE0+SB2GHZZ6jbhCGeHJ7JF7H1AEogwDJ107Z4dGQHapPbTqfB
SuI2SEY8F5K74R651Z0azl3lNOmBVLsbRPYwsCNJ38zN6ziDrMc7Wcuyt/xH
RV8Obtf2Q+nLlQqQoGSrSX9XbP86CzeaCsh6juqsnHsUo7qewutXCENo0Hq5
49/hbnSXBoHyf2whuGcN/ss9xgH0Ij7n/WXw5oKj3Dd6Gek3jyKTN7QDnU8L
9/x28ENkH+VGPYjCWql5E6RjNWyfIQSV+iXzU6maT/hHYOPiAG3zqHBKioy+
FzOWI7fNZFvt1eluq0LQ+qm6y5vCEMDRyXoMdwEWb8iSTVywn5v8OKCdQMET
BpNwFYxto4p6ry2CBUovHMNyJTj/BobWHQ2s+frCCZzQwCTgMIu5clzTYloS
OiwzGYcKzkfO+vS0j8JQMODI4I8ibrE1csPChvKVv7O7Z/WvKjKnXXSu7Qh5
ujkxMc7Gm717kc304CkjHqZIUdWeAK549t++RShWNA/EAjt95sK9C+BSPxmR
3Loy3I3Aqcroqq/WlEONEaehdL/IHcR4g//84v8Rj28E+cKnsUJMn5mflycH
aMmeDm/Eu5XVvExWtYkbqxGlgSESNdMmJejN5aNPP9ksNxMla58MhAJGgPIn
aIVaT16rDTdspEgH8zWUFnPk4UCKeem1qytgaRSZanFeVlUdPgaflnJo5mCK
R1QlgnrHZilBCShSz8ga8cZ1IRzNLtOynL8gGzk5KbmaYMW6DteIB/pybMES
TAw3T2OXOmBuF/wbGLhL5LlpPB9aro0xtGqWEMUs+OOXTaCV+Ogv5Dl8C/M7
EcIkwP/U5nqYz42F14PylSHNQDc+Ifv0dA3ZVaNFsV3aRE1mbN4CfL5dl/w/
f6XJ7ctNX3cUhUv7LaRhWdnJ/Bx3YR49dJwaPczXBjo6ylsII9w5TvFGSmaL
WRQZLnIolWVU3k7nqpgGPp/9AaFDqCRqxmLgtEa/ROiyXDiD8MC7MiTnRQIa
JEyoC3V2q8LS5R8U5s8aj/ofD43Wm9Ca29xn3uzNDOuNQ05OnjsFpxCAw4CR
pI4ZGfDy0u4zYzh7C/BeC0fiTE7jbz0f9uI27ajZl7ZfLA7boaBIhyduD642
QgNJJDyXWbFTaMopBZgVkeSw5SC0d8HGb+ys5kHFHKAkgg+kzlvlVOScLoLg
2eNbSkhLLUxFvSaQD9ObhYj2UQESOGW9oV/FGclrMnggdvDVWU18FD0RZLZ2
5ipfqcb64MIVu0Cq9PI/q2U5M7tGMZ9Is2PxWnUugZz0RZ2+NIFgw1Uunav+
klK4WovDUBUUYcMcVvVGINdO0QvzspDUFR6dyk5Q3KjEYKBpFDwyd7H9ukjl
vAnAQthfPPRVq6tAzDPQWdErNSVoCkBJIRFipSOPFa/EF6UU6X8eLdo/dvgi
Y5iGpCwhhWDIQp9TbHqKxd+qbEGBLQ9bP2XmSs5FFsoZh19NR0vsSlbf5q2M
w88uGs8jp1YctkyTXtUy+Vje22aXniIRuOActzkAAYC1WtuYpnyCJiAzBC/M
25NI8Gm3SvPYen8laVh/ZxL34/Iodqi2N2iIPpCKVX/iil2ouRkzHdtBuiSy
0H3Oos6GNKobYx5JA6bQInGdatnqon8uz5bh99WWejhgVi3p31zn6hfElxIt
U+EeRO84iUcm2e3S/Sr1M0WDObdyiyolmq3VRZfXMFysMklWHQfjkZWqsK3k
VN7hugfcXFKWb1E7NEHaLCohWOIn22IWmi9az9Q6YKTGCfC4rKkTROhtLWIQ
Aow/WahBm7OJhdI3yUFv2SD0JRDHE0sCF5wcViI3w5f2VVs5AMCeGF5BDtit
sMpO9/ZsCFFzMkWypEQOhcHHNQXYxER+UH8xwWwRlmzSjKP0crdFt3ElrXO1
l4o9JoubvO9n0BvxxxooLIGaFpKDyZvpIMlZE6TdGW4T0iGR9rBNC13akpJG
TQZ3xwdIHdZiye3BUPKcfjUr2dfV8zA3isIexHbwa+eaIiD14qpRncGUx96I
jumGAhVeDIedu2Yemo4rbM5nkjVD8TtLvhr7skvR4ume7HFmtOvWJT+qtCOn
c7KiM6TzlZPlGCLZi5mws2XNm9lP5+3ym5WBqiBOJBl+wZmqIBBTupLGuU4J
ll0vuVTs2bznikkMGYEzcP2d2taqCnNI9sJ9onDh1kGtz6RG2ijqj25CE7XD
++zDB01da+pkNllJ7GbjeRx2wge4Q0lmeivaMD0jTFnPJUX7aReO6UWwMqQi
lgIUDnqHxN1A1JjMmYCHA0VjfoALWkDzDxHaNtEI6Sd3CnTPpRuGluTHKwVi
FCvcYTqwwzyRe+KTC9HYZEicypO8+rdC2umWKc/EVXmrqUFsHKmRLvExo909
5ZOPl4GwmpRjnXrJLKQ7fkLJTuqmVlzPPnmpNA6NUGLuPAkhLlAwSoK65Jn8
uZktPFIJakWpNWUvjkOpFkbeaHeyqi3FCqK7k2Z2xrUE3kM7Yoyn7D395qJR
CJCvNLkX9O7yMrQnm29VdVVckdSgrAe2jqN4Q3zXmVg/XhH1i0fy/+I8vTmi
voKcC3OTiz7be3D9IIUYH7DXD2WhZ3n1fsctBjVGd77AatAlHzqytGXH0m96
tkh28HYaicm3u5934j+w1xnPns/tzPbtRQ3N+wtwRhwodvLc2r1ma88HpTTR
db7SRXi2fF4YThZ3QPQGl3SZqEpK2NnNlPocqLG1ZKvdTwqLi8//kWEuv87i
4w2mr0cmcXukR6lpBPjHoJPLMa9n1owyBxwf36IoxgpbvEEO9CT9VuXnN0TX
jhpcSALxuE8kas34YxqT3sY+BBSlF87l3mJUUkZNFhOOw/3LZc5h/3uuzjEW
j8bqcGtTw+jHQ3bXWt5FD+AMCEihoeP4mRMZlOeCY/ihz9pCOdeINqqmUnpz
67bmWXCZYZaZKGOVywI6X3iaxvBgu0PoBk4oluC/ypqnChQyYV83Aa6I2UN6
63r/Q79ANa+hikOobteNE10jGOTtP4VVY7VrhISAYf6t09jbh1W8jWVEc45r
vPIgU5zEhvlsi5783JoQUqHmuW27x7Q35hYoPrJSllZhiSKgy555/kR2l1uy
eZ2p3EMvuRWpJqZ05MFB9idBAik/UGXX4yD7MMvAxUoTtvlr0/LfzLbKYdYT
V09g/DdrvVo/pBxv5EO+qp99vV8k5qwQT2tMYcoP1KhzguO4bcMypTNwUe2e
5uT1PzLgr/vSKqLRtez+pfoXzcFnmbcjjQ4XF8HW3w3W9WXqWHIwgE/QK9cr
2I8DOVNZlVPmZSGOa/kSpoXWlBXZgNU5VcPurLUtnhWDYhJVSWtyD2Wh55nT
rWNyL4TQmiHCqDjQJ1ov8rqahuwav0UdkRdqXpsodB+WSAYL6Iv2bQQ/AOzF
NJujipAASeQi0t2zts2tJF3ReKTxn7Lhpgk3KQcXi8DP3kOSVPDGgY3kB988
oEBx0ZCeGUaIo/CX888/Gvge79YRYTetrD8uxKEUZ5KXEE8hA74qNseslOxz
Xa6qdJKZUFjhYYdWxTq25uYoWe6rvDSsVdUaOGTw6QKdFsNEfAmgC5nUqwoW
Ji86MdcGDPQ7gOPrjy9H5H/LB5M6gCDlwZkMbl4AFrdd+9hK80i7VJut8SwO
GTg2VNQIJQ7pUb9TPKcILZAcPwG0yvPa8hZfrJFVba/d+6J8H5donkirfTus
rjCEODz3pJ2tbeFtKfphuSJycBoMVRecb2iub2/kdN0Bsw6sEjNix5Zyl8ai
f00KoitUzJWlxpN+xG7g/0+Wx9Kl3QFgfd3E0CkhDiaZcBFjGwDCeI9PgPfH
j/+e6wEehmqQOu5DWXrkLnTvsf+F7sp2AbjQWFM7RAa727+BK2POLZRH8bpg
AQ9NJ7wSqOfYrOB0VwhBQr9iQIzIstUa2tBYIq2Qt53QGsPjcUlwq0A5h1WK
UIbj8hVgSQ8qXAWjPbhUObDfhAFMreS1qYdzKXTIPzVIbvz1bB6QAADrcf/t
RBmSdUQEq72ngT2BgKl1R4VyPjrf1MRLqMxmnwHvYDJ2LgOvFlXiur+JploF
hnImVa5W8kd5yATr1s61TKTxJ3TS0ByS8hepZTm4e/3bQRTeeqvRemAA1ZqR
f26H+A33hZ/FFjFSREDguWFHBwkuocD6fu5INPbxENN6LRZdQ9tQNO/gD7gm
SpNHaYcY7SkrLGPyG77h8AeH5foPDoZCrK/TFoHMmWaf+JVTgCfk4PIlBR5v
I9XpvOfQDxv1D27ZK8RgYwkXQYN9RRI37E51Q+Hiu6ucEhAdyfw9Gr7ATokM
Z4EaxOsjw0GLuY4hJZzxzDnrvEpzqJPLP+jVCB0yo3C4ycaUJR2YgGGDdwgG
98/zI0RSra54vE9d9sUtHTEzsyl/FhVLXSsKi7vMSs80g1fUuUoQRbPBCQkQ
PLYUfNgS82WWYHF2l+oQkb/Q1egOqLoxyMhG4KLD+UjesfScowqET9ifrZB0
1kqM839xKEo4rmqzFvGW8mtKrMtKTqMCPwunWT7xV6zh/1T9JPxB2ocXnNeV
e3/VBBULhO+8PBrmaWQq2Jp1YGvhfkbGQXMjRGwuVLpG1S7njpb8mMYjonaA
STvzUzqepbw6Ix9IffLxBDyHbdUCFx8wLnINKLymy2z9XrZ4a3TDzHZuYw7f
ev+PHmkQIQQRBQRve9p23ZTcOGABYMykg3ZsRUK/vPgmBq1i7ZWWkm2P79ac
0jPp7kigdvhX7gHR5Xgv7pNM76cZgyGrtezNAOiwOQ4qG3sRIZN4RephUGhc
v6nZsq0Z3BeaRDjkAflKAJGuCYPeH3JKvgAdfSrQuv/pq5NPiucHDF8DqdYH
d6ldAheMbIIU2SmmM9fjXMTeiYW4moP8ftno5VDIdhADpQP33m5B5dQxu3XP
zR7p1IXU3Lp+okPiSe7kov2dUtmQ7JzABiRAhDlCw9TE+oV8gHOh1TE7m17q
oQ6p1Iuwb76yGA1P+S6zFV2BBCUHJ3ELJ5ifnzXKvbccFSZXpTLWAuGFhIFU
1Kd+GuD1nimxM2zBGHjEOj+e+uszvVnUrw1VD+tTTkZEOqpPE3QRgzRrulUI
sECMXCaYxtDiXNiSNskRMEsmvKGNirUqmud7VJxRJ8hIpI1pMhIBxX0t2/1w
4D1sxwZRFGHkzOgg7w2qUoxWTn/+li6CPq88uueFKYp+KZ+osr1YI++F7/n+
wo5BiikeVSbBboIKpIiRAlKs+mirLXcDM5wq6v5unZGKdNVcq4Vqo/jlTfkq
8l9a+oHayxkFMD51XkOQXxPKu/28Nl5MnPvpIXep99/zSmo1ddk5C4EZ9HoD
QiaX4g/Ff8dRJQlI4X+VEVfawU9KQiTXM5J9KdlLsZeF93I/VKJUuP4DnaSx
sNEeVgNpwKKh+pvPyuhfR5YjNRV1EWhVORdNANk7q586GRRNz5LJw77r7wxw
XZ/MzoGbieTdhBwuU+ol3aN4POCxv36IYCZlw1BTB4Ra/gHkheExLv4ua/oh
tRRjvfG92AM5juGD9/yFjHv2brN3LGoBxHeP5eGFeBu3ipZLAq56uHNKaRzr
x1uvkwNCPSFd2bCLxFcqPxz+X8wscAo6t0VlUDkgIJ/e4AwGObI9CBeQ9qLe
V5kSOAJYcml/afYYpxYUBhucZSGTup7PfuOL2dQQ5P7sr9HztlJxa0nAAmJu
eIMS44kR8Y1FrcGIwESKyYzC+eqVVDCwgmKf740VLm+zVQi2wW8WzF8lLnxW
dInFUNEOtGow8qNshZxwgsJK6ZOUB6AA5+QozPLbI+hzpvbqggekZM3pf6DL
coFJbe1k0wp+OHzjTxzgtOjW/g0jKUule1j5JsvO11GS2GkteKfF7fNlUA05
E5BMF07OvjuwfSsrmxFcg42OeC97QnycSnI38XhgqjtePzK9C36aNW0isoOq
+C8SS7MLR/K1DvoU+hcevO9Lx1uciTFyEvFTKZvakhdb13D6hz5dfshhedgT
f1EXCDgK0VPC6fpN34RqHBUADRDFvvLHHH3TNfeSWcVJQ+uD/6VWGRS2kMAd
rUWF3yXcYuDCJTEDeHPWr4benY0FMUecHy8fJLhabJCnlA8CPMhRgDD7r7Iq
0sVBHNWEXT3XLI+aZtOAybPXHZp8tOz84k9WiY2o+UIAlbzNANS7ACe8eUCz
ufJIGy9rw8SuZerRWQ7JIqLTnMcCKpPLg2L09/x4PeImC2s4SHK6gwK6B43f
9J5HKyzHEz2xx9nF0wSHeRpdVdHQQjtjonjeSA0vqI1JoXneTm+7ub2UND7v
JuUjGDXITx5c/tpnsExRX6Xdpp7zGrsbj+pFrT1s4j0Why0e2Xxb0f6tczX/
gmM+F7qV3WUIK6D1tBnfLAfT9R7PAgDLRtjScDtJonE6EET0u1RD/NEeATwC
VJGJpkS8eJVeqt84VB7siEo6joojDFANFg4a8lYroPpJpexDa9N6uKmNQUq3
yT6r5YGaS6FuD0uGIFKEfrgae70agqWvZkN85FAylrAykTcztKOT+fwxc75X
u6NsbKF8C114fP1mJ5nXu4odxvoRlKgXb8+w5Nl3nL4aALRQbW/5+XBOtLbI
NM0a7u3pHuU+Ez/0ye/HNfg02ZQvWFF2nUZ/3+ETemoSGxDRi/IiI9Owkcw5
es69KP7xwNP+KjL++TnECTKLZvnwXVEW8iXZCV/d2NrVh4u2ohQOrSlzsHcL
eE7pDbQsUIu67F3jEBem3/uUmg2ofq514cFIX3YLt9x6W9KnhWCcpEkB72GV
dfTykSNq+m9weqC3ZGluypVgnj0Cxo2GSA4gySzQQ/YMdAg5IooSTq0Bq2Dx
BRaKivV6/NIx28IW9GOYSL6pijj2TckRBnS45n7uwn3S+8oc9DOIpGqZi1TY
wM5QcQSadyJptA60ApDM3AZIKsYLI/UBZMur5GvdmuxiZLBjZkfUYQV4ZmdN
Hx6dv3GAzkb00sIfYNgRsYoYYBb1j6665J8QQIkHdDluvohnIwqDi15rLt58
+txgjq64VXO7pNLvUdKBc+n+yeKJGt+CO+SeqmFVVsgejyka4taN4zVlI6lq
kck1xaXJzAm3kQ5n1/w/LVgv+pU9w5MvWb2jEAoYRNqPQFDDhvtrBanfblj0
inOg4X3y2XCRfqmdPFlCNXEHNrxH8r4f09i6fXF/A17QQreVJf+mzavvdgOH
8Hjd/byFt1g0REkc0VcHLfCK8wPfdPRp5KK1KOJ2UK3PyNoD6E5DyK9kHnVM
U4vyqjIZdvMkSXyqKkxZpEakPj20lreSvOz5rLmd47wycoU64dsfsA11Cltx
LD/99utdyfPhh0VCAYtGHHRySEWlVexM5pJk9lkVOGvTAKPMA3OTycYBfLoP
pwW7wXHV4wI99XV1bMt8c9rw6lEA5XFiaKUh2lPKBsp0WV5hMNmEq74LNr6w
iW6c6lwLruJ/iZvvt7F9LItJ8to/X3Wes2flD7levc4L1f/rnwbjGe01jhHO
rQhaxx2lWBkvu8j0zn2JaGm9trcpBlHsYsvyRhHVvSTgwZQYHzHwVZ7iIeSB
BDkohdjIjQsFHu8kgOYkrp+Tt7DXmGr6cc+TuWfd4QpwgBLDNEoUd/Uzjhfk
eee0D+VbCjLLeGCcshjk3HdcakArt2PNK9m2hLM/gnQRYmI3zFA55xKv4qs8
wQbmhaZjK8gmtK6Z9u/6QYwT45FEZ5YpcY+68BsT3PaVeFFBveQgYqbInXXl
7x5YIJf0O+n7JzulNT5IxQ208Ch+mtQ3Cvht/H3C2tjgQ1PH433OrMS7TeU/
iOdEs4MBAEtVuaZdM52pa0y9/C3gj0NTrFw6+OkaBWeSBqZoRUUBYj/QfyCJ
7VJ4Z9mA+s37k6kA7LUFTxWu2rCXaH6Vbhcbxgr0iF3Th8q+EER0XOh+hqS+
TdS91LhKliEJGefxf/Fz546l0mpNzgEspG1GNaB5IP5ldQzCVWBwtWYHUhPq
BTIHt8CNIMcE9wHjT8tfyGLqWQLfcReaKEw79+o3NkJ6ekhJP9yV9il0ZKcm
U02dpR4KoxBS9wAdqlys+we1txocF/hv38L0G3cM+fROxw+J9qWo1pd6RmS3
9Rc4shBt1otS9CPhQIb5I5MnB9S13sqyI1BbeK2omNjlu5247EIzI9ihvtTU
D4AEQ4gMV+wVLgufO5AGiHqIG0bCYGWtja6QbmKnTOsu30X8aVV1Rz2iEi3s
KOpuA+RRH4E5IiGv1qo5GI3zwbQtzHCpEcFM7M/2A9vi9KJq2JABbJwvBG+Y
nNYv/Ghi9cs5E+37ptXYDsGPJgj5dRePWksow5Eq7v4n+scIaQdzgjCEAm3j
I75KW4jOcdhA64daDIE9YNUoYEDi4TFAGeQgCiNeG1YXEkfoHYmqKp2vQPoL
Gk70aG8iH/bnP6ilbxpaL9WCCg0o+TuDsR8S8DmyJKG33IzXi+hYSXamgsZk
IOJtHqxhPgRYkZkloU1h1ead6wFln8EX2ZJSpRIi5XtulDcsxXPbDGpYuiaL
ep4vDC3YCzZYxJSpkkKe5lSXxvFC0Jt9L3StmvYn+DfsaRn8ZWRrgrHYn+iQ
WQ+tM630qhQkn4rChdTcQGbK1z6QLoJ2gohW+0uJTygULlx6aGDRKnaRekIr
/aCL0sW54NViLOF22BKm+Jw/DNsFm6A97x8PzNOPQ6KlVC6hKZkFWlx42k/d
fQHtmT45ALzgjXBMyW3vBZIMENlbhF9w8gb6OtBQq7bhHAST/+o0ESNZ1QkP
Kcu4s9W7puMf4ltMZkSYi46icsIyXsYDVAPbedxacTWZesixkkjBx887W1FF
Rb4dFjpZ4jFcew9xScUIgd0th+tD46SvhkH9Bhm4J+1sziuqdAi4Pd853L9j
yr2TxJhMQxVlsMKYZNJq7iD/r2J7jTtJ1Jc4nsARvc/S9fgZ1t1R5bJ18UzA
Eh/it4yzjTI657g9C+wiBr4aIym6qChfHTaC9pdywZvUe95tLSbCR4MrmG7l
2chBgUcKTm/E5cwNoZr0QISbdeZF3qTZvYcekcCLdbVBswcX0ix9tlbuXcVc
ujY+S47b16J3nnoOYWj09hP/D/nw6s4CAfxOH/YN8l9PiH8XSPx+hr+mi372
gqEikKqXlVbWy1/gVl47K+fq1MA4sxUH1YHWLXlfoUljfqafnhv2XPrJIt5L
WYGvZdOTsQnTr/pk6sUUWekQI8NnwJVRujeZylKHa6EVDCoPBrHwQr0FZllx
V6AdJw5ZaQS1b63jAhhKNLpr9hsdmbVV4zFiUXkjyDAhqYNgnJpecSlN/+Uv
B6JuIkUYhFCVc8buUtKQYGj34ONpBMc5Vs56Qyfi4rY5xg/vtPGlJT/XLdbM
W/oieNHqnIphV0yI1zu8pw5JxlhNK6q4Tqbj4xjFFeRJ4oH+rka7j8pgmntE
KsMPdSSihdRONH28XD02GsHbqLYG+ypMqK0OdycuE2moS1TiKpH48uWV46D9
b8jhh2GSK2dblkVjBvkze2WNm8tyRmXMgYKJX1WZd/Sah7TYgTZIo9xK6zDL
uKnrAqBeFggjek+Nlk6+kN6OEJIXAB4Rvdxf/0+1q+eQCuk59A8i/hEJowvD
J5l8soRyI5aBqHT0zw1Zvm2kJoxi8H2LsnffqN5hIxJR1MLAlLm/5KobsC5p
QmBlom7tZLVmY/Kc2NzxE0BS6J/y0SWQj8wE4FlqjmTHpyWedM5QUPcaH9tP
MrLGEWn6yYwrF3gqrswop7T9cgJET9l9/xkOJInqz4NwWywNYeMFBWqjTMz0
rwUEWKm0koffUbAYYxCTE5GnMYC0/MEliOroUgrLU25SXB70Q2CJW9CEips0
+5YwPVpuI53Kc7ziKAtDuBXToDFYssJ8rB8O6TZ3sEKncgvdjkpex3Yq6CL7
gVYRP+Lg/l7+XwxN9X7XsNzac7rGxXSIdJ1K6Dk/gHVxbm7DCqJp3EYa5l8P
aaQROvfNPmPjBnfLZrL4VibeJuMQiJVVgGa9P7yqkt7BopoeYO21fkBE6hXk
lslUsM4zPtmEVap+hxI4PH2NjcCbyd5dlSOMIzcl76ok6zEWvcHUzCD8gjvY
Zvl8zS3kj+bbKJUthM2G9AVpr+bdoWkX6ntZAzU47buE2AWzOkLk94sBu3sf
kojM4j0VZr45GvgtMdS/byHlksqwcrnfeCYgmKn0EdOLD6WDodQqSKEBKOcN
E58AV1NZtyaZAtzgGTiLnQNhwaGei84iveAOBi7boi4pDearsDkml/ILV33W
qo555t6CM5hIiTF70Npcz7CBe/MHF0U4AjEIjWxnuCigDaUTJGusZzUUDaDC
BGL9NiY3tz26EKAIg97QIZa+tioRiOOvxLC4FiHZQUs0xk82QxPqVQvlcM24
7t6Ws8/e/qcG4I+U9iBjeQt9zWnaizYViqctWLgCS5aFgpmZwbl6oTRot193
DTsN5Ei7b4bLwUcGPaJvUhvWn18w+Z9RCusZGKmIBxdfOixKUe4rmkXyn8ai
DnBp0Xhu6O0uM69kWhLGUpi3b8+iX+IaRO1drWVPsO2YkrJ3XdAxCQ9l5KHC
Q87l3Rkyb1B5AixYSZcv8OJc/R+RZ3oQDQUAyW/E+TUZZA2RfnFD724oWCaE
JLEHjIS+zrg4fngZG1rwme+I4KsLDBOpebMMDyC1DrzqSMxYx04KywTrtYpS
vpiUHs0kpQ7GPDaRtur9zcJwe4OHKIZ+ky2X5T842GBJuqt92fyALlAQasC+
NYOM4yn0H0JV1Hlu8co8eHlxaNmzUIEuBl5VcqkxDjeuMZepZf6OhhJWq3mj
+rXp44X4utdZX+s5x/kV80csLijRx6qp5Ce30ZYc57Fs8xtRL8iVhyMEhUOb
BkBfppP53RT1LKBdre69tB6JL10/43DY9mVg09VhyFKW1jRQYHUzyOzM08QV
wKMh9w6xVCKBBa9K+pOsrggjfx9Yhv66XEiQ/ELQJ0q6/NRnB4Hfn/bLRUPI
o5OHE1c84uvvJyDTfsFs8Syh55eSeyekajYRIqbXabNxb+Tdf9ZGgxCW5YVv
M3YQIzu/anugC+bWFmtk4KFHLhG1DAHgqVZXXmsyhWbwtfW5RThJ6VuSuOoA
NtgV2EXh3smg0/4ifATzfNN1UtMK7qpHXdBihWz7nGzOmS7ZXv0g1e31u2T9
jUdwkymdv3RQAVmWlR+LtMPSGJpZcZ5xoKL2W/BjQBs9ruXAfvchcDImkxLR
Uc0bX4O9/OdrtJVe1OUfh1ttKlTdswZbYK76s6GSptTv+E6sOh8cE0jPKlrx
qIgUzOdKOTLJVZVKOIf6uewIhyXL6R2BfL3o5FDnmVS2kPGSNbcaSDfyp7TY
Oi4Rws1WlFWP2d2x/CpW88Y8wpJxr/O1A1Mfefi8e05WT3xKTRMyBQZa1Ydv
j7JviSC9dVYkwRLzFt8VgTbCh9fQKMLsjNPbXNCrxm99SGywlSBzO7OPRaOY
WaF7CWRBOs8l/BDyHUoB1caw0NuZ714wlUfeDJvX7gAE+Czff9qdh3CziI+a
jh2+5cI/G/wfZRpQFV2MhBSMsdgJiycQ88RM/wJCK5+5RwozVqQzWCBfu9Fg
M6gMkKlhsT/TfS8j2kw3kifXHruf7p91NY2lXPQXgxJ1Skh4kI+k3uLW8Q9c
cvBDA/X7yIJr4D84/2zdxJpLuXcwcj2qDFSsF80dPzwyuJrF60kCYPeUudtH
wsyFL6toX6WI+fZZM0u9pLJZ0jM4G0A61JS8qmnjcW0TOHeKFqvoV01wHeun
bFv7UK5knQatjhruEXSSa9ToXJTRURlrTp6CgeTZgP682fj79D4tiXZs0ofh
mp8e5NDdB5X6/KLIWNp0SuFmE7Wiz7pBvh6vgacOfeJbXPhldNzG8gGDGI/J
eWfCjkS68vbybXjA7bIAaAdabQTjOr1z2drV6A56fooXFZ2ixY0W0Pk445qd
mcYBlg5JunBrRiMOvBe7CEgOz8Hc8cVhivzRr3uRZbFNAqX0uZOqLE1LKbza
D5u/bpeWUvUOIiVjzUJtHyQyWZf/tPlB9pkaJUwz0vCTVyZjIwDz3KA1FCMh
TXU2Vu1KeJBaYHK1wUGXxTSlTIBauZJ00uB2KQTYkNiVq+uhkg/rfDddDmoN
mQHT2VTFQrjZ3D1B57KfAJxHUgdSwE/z2e7CbQfNmvbQRDarFXsym03svJnl
DPAPDvIcirLwFVV5Om8XpY+Rr1ue05zG6HGPXvBEigB4sooiGa8OewVBRZx7
HfyNJuHFdgRTCKjAH7ANDOIjPyrLQ4hLD9qphb0gDy7WPfwoljgAoAM+Xpq4
ksi9SS/2LdnpIv6LYU0jW0gi28IZt/1p67SadK44q8ApXa0lO2lRKFOLyxU5
oBxJ/jfwTXq/WbQs9j3H7XFMz8VGwbOKs86GuZYWOGGclSltFkdwIe733xkC
/MnF8bT3bXhHmiJ9rC554aSyfZBGDiTRU+/eHcpwI5Uvy/fbo7cGmnpbySH3
v69SIIfGwH/6VDAMgNModtcHhkuxQDPedVVkwg1m7sQ+SHM12G0BNI13RyK1
T48Yc/o72ijbwFgkPZWz663jS7Dp7QurKJkkjKRXhOmFCg40DtRmMI8qrvvr
jlZDBcwyI6lY40l/Q45jWwFNbugz9mJV9sxOeA80PXnDBaj3kF6jrJINt8Bf
4umqCsscO1g3agzsx46ssdec7Wg8W+alLfvyUez43caweLqLp8+X4k5zjhm3
tsGNNuj+xi//nYFEgu89LI31t9fYhbkLj5VV6v9guOUrd2qU6NhwCho4/H3E
Esulv/XZSNS4RaIY//9sDoUWpSl1warrqn2CJ0KBl7IrUicQe3gSWirUiVti
TJwkU5CPN6DA8Y38RHdte6p4d0Z3YbJaPUElczfgsS1GSYhlgyFAMiiB5ikY
MyCKqOlqhUZSoEhO4sn2Zztm9kY64k88jFqUKuvgaXhCY+7TXghfXiODoeDF
7o64nWDgUCfUe5KFNxb/G+WV1PDzOlePWL079J/Pw4Q80RbIJreR6k3c9iYH
WPazkNQlFosj7clFKkFUVJTCj1/vJgtchbqp1RNtXAHbU4pA6L2OQfQeRz5R
oCeD1BLt9I89g7H4JGR8Dbpb6/HIBPfrMJUDmtHb/x0JUXNX0fQFYgYLkE5K
GfjiIr8RBw5VXgJA6lAfakjEVDlnzk8pJfU/67Y75TJpfXB8Cq0NoNnvJv/F
u5wRvQijENS9wZkFIwgumRW3v67WIJCopcP0ZUMtu2qlx+PJ4R09jKMAJGAt
Ljdm/52i9rnK6jKYw/H+OPbylQ5ixllHECUR5MKh+xqyAIgnMQYQQKu3uaCS
ETWtnF+rGd3Hf5jEA5EjL2olYQmMwhK6czr41Vt8Rirm5LIA/3R4HJnVJBcZ
Zm66uUSZ8agfQchdY2VHvT7x9oQeiS+cF5fcI5nGykDl79gIkqHp9pihWADQ
AP9WHOqYsGC4YpN5KUU1s4EdTCHt6p3BfTXtdcEWyLaCl1zdRPGQg2yrHSGA
SaOPJ7Me8RaumiJqZuAufZ3eQjNw0VCTyc0VZLxONZzUJDDmecDNNt2eUXEW
rjsbtN+nY89kLyqLt3AymPxvOVzpoK6rSsd1ewg0QlY9PDf8BR5krzPnMZG8
zKRc/2jt1dxSi5Zxx4lNxjtJpC19O3VomMWCahnFUoL1dLk/uNOozm7iDg44
hTy+dcnU2AgHwsYrx1yymzewYeXULY7m5Ck3R/5YhOQxKZpUzFIMZPbXj8dA
9gPNYqh4fNZoBNtl9a8j4E5F9a9GcnBfrr0JFHgOcLjBok0H0cI6OfVL/+5k
qOKMs/og8c6/CDl9X5w86bQxDWKuVkaCJNU7LCkaa3+xo0XPgicB3u3fH3vf
z2JFb5vI9kaL3l9IK+pHNWR3iSzXEZ5shlr51L9NyXGsiXpQmO+JaBn+X8QQ
AbYhgwDBt0yn+dvPhKz4CHXQNaGEl5uYSlbH6XKotvkL4Xqunzwicni662Et
DfqQSlAf4D7jjPw/lWhRSPZDIYouL6NMYaelHiTZSWvZrY+KhOvvfHEpHWu7
TG37VorAB7DP9LcBGnqSn+8Mq20lnZkzESgKJE7mlsAFAXRGgVHTGElm+e/Y
6YyLLKihJSStQf/c6huxdkBXMr/Z3h5PLP6LMwDunmTyxNUBcQC2GzWQ0wLH
LZJ5u5kK8wcJ+UyzlfYIOpadtjmrSeWrZQQ2pMWlU8Q75F9fIESGi7CWUST8
J8c+CTtf8fMQp/eBPY++UpJNaepN4SFCkvJmr0Cx8CMdxrPPabKBVax52VSl
48ASS1ZyH44rxZmom47rlsgKI9NNp9UCWTdFXN/Wf0Dkc/YkwRiY41V7LMxQ
9AOTepXdGu7FFX1xzRpc0nbsc1PULj1CnzlTinDWp85qaSOF2JOEPVUhdI3g
sl0Dk1bWwWaPeikVeu/w05VkXwYYZO0R3pTcAjxwJyi0DBW9da/T+BnAnkOU
ubfAz/LimeHXlh28+AULY5xLXEIKTCu/dtS10W/kYH/Cv+1a1VDuyF/zBkOO
9MuM5N/u307nJMXytIxJSEKlUYfPjYCAxsEHFtEepj5bKWYiRidLBk89N4Tq
UJ+Y/iMzr0LdCGNUfy2+LqBuiUu9BV4CxBUyB/U/Q/0jzck4c8V5dgL8X1Z1
dl+qoSJZ9UOLbJHgkjy7aqqWtXmmUOhE7LzxI2MhHIeUho5uSbdpMi2/JyQk
n831XOW7cscExrY0/1oGJ7BFl+FtEmBk4M7EHxJwvqwAlie9pBoC2LFP9J5f
W2aIK5Rea0mSlSFKoolXtiEgel8YnKTgQFSXQMnzN6stBGhHD3IzIzJmWfTb
/wdR985UokzRIh7MocEXVhorcYfRBzRL4pmb68OKo3sMcyt+6/9+wIj3eB7g
CSI4I4i7AdaPNZ6HI1OIOf6tjvjWrQbZUqmQMyxZSfyA5h8kCFyBVA5CF50c
yAzY6ChAgtXM74DMSQZF59bbQ+ZlJ81RlnRwKNK32eUSG2A25byJWZrC730k
1Ea7RoezZHB17v/+J7t1CI5HBFnjOLmN+rav6g/c9LDMAJb/i28JKPWBxWSQ
HKdIHBeKsNjfV2p/R4QBXV4iMqr8sVFg+5YgHIzJdcEBBxdddeq7QX52xudQ
wag4TuzrPtJXS8sd4XsgLKwOuwhLfSowTyn6bm5poSV1ANk0TzKBZS/RClsv
DdjGxoQVAlnR7oQLB9EQiqKmHO8lHCo/5eV7SRZXmB02ULuxJCJdF6R3sW1S
2C/0r/olfYMATQRDLZy3qYU0qO+we57Udex3XR8byY5bullqhhKbaPW2DHNv
OvTvxhuk4n6aT8jjUNGNtOCwPvzFuLylGTJ6jao67zD0zpBBDUpp6wE5dHaV
df62QwZRbhipvrqLNhcs4af0SAKQ+LnPnnCVDdmtkqdU0PyR9h1L+1YiErdU
uv/2FyLquYdP3iKiWHSKRERGG7poHOjAnuYheDvuEsQXSDtumrR1kQ+Ww86r
SMo39VpOQ5u2iyxfNwPtlKnqGJq9QeUj/v86jk5ziGeT46/fvYBUrbeYGUBK
KBQmmo1XuWK1fUg6StvWLZiSE7KMYEsYSJ1/8nNzHftJI1VpY5k8NXPj/1vM
QipLf7LHyCDzYQpbNxaFGsDZYCdJ3W2lNqkchIDBfQSshuSwiKkJ3P8XUbK5
QMZgjsqTqdA8moLw5S6ptM2+juocKLRRtgBpQ6aUHM/wdbAWd9Dfovwq8bBp
kOKR+1m7sIfxA1pIiEc/jFWq2/UZaOlryJf3I8bKqH6uc6HZkESys6bKOwcx
iRvNlfdelOcQVgBba4MvwFP/zuLZVY+NH5ePP87SP6Sykv8mVS4Fsl8bNK3N
5OBO2IwigELLZmfEu4I03I3GEs5hyqmqk5JP5VUfMlXj7/1wQa+7Qv9hJO8M
GNIb1ZRWFhiHzI7Rk8mBtoNDETXmKgeuh2s9Krs5r6KMqGYkQeA4vY0hosNZ
BxBV0pbHeglDq7nUCg5zv7zJk3JJVUlg4ZijD/sg63b4LAqQ7mnzgOpnj9Nb
UlTrCL0mGn3fQpqBelCzJBL5apm8u5CwjUTJ8kvYAwTx0JpWHicwlE9Ro2Dx
5b9+r7tU+RxSpnOMqi5xeY5eRrnSvwAmnGbC6GPuLeZj5ZOX00vQjw2roZNy
ZW/MWmSD9B68mP/fAK//TcK//uNyF8ytwrVL8wCrAbiDp94yNKZbovrabNqN
aTFxYkI18ME2BXtrNJIqSCjHUeuGoSzvjFgB2OfJQpXgttk/Pm2IYBLz3Hdz
OqijVY8BLrLnRq4D4clRedN+nZrZaguGvUMhcRzzq36/2569bB3Dn5YYAtV6
/MfH2laixrWHisrWNX42Fc4x3S6Cw+2P+VsU3Y31MmhzWRnMrH041wDPJG1W
XdCQTCw9tOlMs4Xct7F9eF3x4h/FGd5veGLj/Amfx+BtZYSUt5E/MNBY7fbz
pLHiVomuwwI9gl826tbPqRw9ul7qVxueCkZxui9xizBd4prX8jV9NPanGAOH
ipB3MpjFSahzTzh8w5F6km+PPQ1isnwsm+pSN95ThXaNDv+0VbaNAsI+sDgm
IbbOd/TVhfMPdo3i4+UPK0DWxrNUhef3WGdJcJorHXAx9hhApX8td+0i6+IS
L6wyweyy78E4rN0OfGnk14dKxrkuAAl/cR7lBczhd/lZYvkENT6e4QJIf8rL
W+D3RitI1THzcy4Fakv/DJmRejZqNewtN3ttTtjY5o4ufp5CZyxVvIcVdHFh
c+fscggEqSaLjOHF1WFdXpJQZNDahoNeIo+6e1aygu/2MsEqVAaawBqAnPXt
oWKJ3CwjUahSdbez0ZxU5EMp1Mi+tNKOfe/6WwjGM7RN58XOADBbgrBJFFtD
Xn72cchofR1ymzyUkDD3Nyh9ZagRBgSPGhyxNQzFEMSFStBboMdqAjjmVS3C
lxFyVHH/liYVm7IFOpAElrfZ2rW1D3SEjRmga0RLOvdbweulsgmEmtic9NS2
nrIgncyYbM9jINmBeHoQiFmu1qpd3TDSGPrRVJq3emqwYMP6i8M7PijIs2kM
92LZTYsem2MYWEBBKyHM4/AecFqwv5AMNcZ6E0+zNuDVNN/4ItmHAD7pBxGz
+7iGA7HusUIMtHR04tT+z52xtc6RfWZcHGXXkHjllBc50kGxrxsF5Uz3ITM6
gJGDz+ISGpiLqIoJqaPSRHMDEPgyaaxW8Xw2kE1UP2XrmB8RKob9450Kkx0b
Sw/pl66b5+YEoEMCXLgDDB7khR3n526bWUGo+iZxlxnPMYysCOa2j3h8Z87e
UFjYH7UkU43V1zTM3DN+h/lxd999mHtO8qyLuLdVAyUbkMlHC8qsh0qjo2Nz
90iwiPiLelu3yhnei80wBl7JYvXV1hr4g5OFFYyxrk2mzG5xDbAciIsRffVG
TfluMOVg+2kM/AxFfgv8hDvDINc7d/FezPUvR9JAHGguQGzJlhHQF0xPNPkP
hwHoaD1QGC3XzuIvOIFTTyuq1rgSHT51VegnsjzDtONuBaKK2kplbbHP10Bn
VUrmV5zGrvMGdsNvLj84y0cytS8fuyEAjx+8J4Q/307+jg1IjUq8s8YuPdn3
W1FAmvqJLv6VNbzP47F9Br3zS9sY/7Va5hhYXi64q9TSxDQ0Cb/wpHO/7tFn
b9yn5U/PcDMalFa0xqMaXfVIxR9bNKKTCzsfhHWEVDRAmIhz+sjsydqrCC0r
BETImFryHfi9YJp6zZocIcj6yAldmHeBQgryERnKdjt109TQzqdXnsjBFzHZ
2LFBqR20Z+LR2I/hiJBNHjPRnGWGxCnbZp5ya7iA7CbcU4paIkmSTs2ag53r
aWFI1KlI/8mk3WfPmctYjnQVPup47vPwnfjZfwS3s2ROWR4UlBP+zs8CS8oj
MJ+GRi2SvsXY48CdSBPsk6dt110dR2eAY6AO+R1pR6y+1VrJrjyUvH3Mixy2
xkcEGa2MgeX1u0H8LbGJCprnQJYsHAt/+WmwN/E7tFz5aZj6VbtxplemVsLv
0Ty7DRWy/HYmllXUfaiW/fPPZA01IAycaLf2aAQnEVbYQaSGVqBr99IpKZPQ
EDpbaWT70OyFYxJIrbxHOs0GpRnrVKzas5D7L9TNPF9rTReuDm03s95rZzqE
3OTz5IUJ+JUoMLeBSSliWyS4KoGNAFartaZQUsj9EYrCStPv5ySYFpVfhs6i
wdCGagNvcCm6Af7U8rluqVlA1iLpQnp9LilcClHqaTR0S/D9Pa1AHhZZ5YD/
HL9ueDxQwPSumFIZ2OuLN0gX4FFCtNi6g9BzuX8K1NMtD5NR8xuayAjHgEOv
oEz6MevmeA9C6tt/FzWgsJws6d6q9H413Taxdf+xEzkqz85Z1EWS4+QBt7Yj
O4EM3SF5ygXCVe5fN14vc2ugtFcFstYp1NfhFjJEOsuJZkdFep86TbiQdm39
edyHZm7+HBIlj68rS5pCuK016ETulPTAxP+TkLeiBpTZb4b6w50vLXfaLvCm
aETEdJ9nF/IgRNvG8gEjZ5Ub8xO0UHYXI+k0Gi5Fd32aLfJasLwxMVNxGfk1
IsOD/M1fXvEVD76q5rT/BTmPFhEEGQq2B5DNxwzwRuqr9v5TC2G15WogEuWf
KRi+0iqO8Yvhs+Td4R4uHbBvzF1vNdBcvU1dZO8Ppo6LwgVBMo2X7BW632il
mNTJW55xbHF0H5/ISnmYtm2cYmfFk/Asct3UjtbMqWZQ7Lt8d6+HiGi3vF5m
t2y5abjyfzH9ImBXxaq9kv6iSRVufdePNGU/VCaIudv82iwPG8PwjsuYaoLs
5B6dpHS53wJUWeEt7h6kAgfqwWPp+7Z1nEXfvbHGjF8cFF87d0hLI+2GHq7q
cXqJfWXbk1wZ+7Zx5vGZQtEcfZ4mm4nOw4SwsLN6VSwqdlcQaO/CNy7CaOBU
LqzMWZdOqq1/61Wv41pQL4j9iRHg2a1JQ+IGVq858jciB5bNbg5kVe7imsFW
Kd3bZ97vmP0/cULZ3kWYxbJWjgo7GwfkFCvDqFbqe0mYx04UHZZqxtyZGXO5
xmNASTFOO8OQeWVwxa5SAmVHVtt+Nl/F2/mdrM+erpK4iHgwhfOA2D4FWLgH
CI6+Bf95aoNm4VpmP7FKUjOyeB7pZtu3qBxN5X0Wfo6YjsqnWwGqezTUaJoy
E2duVIoRUvKJE85YNO8HUzhVI1jT461YzYZBW19OvvDcywsIF5/FubBYeNLW
q8sMsLRrjMEvZOeaINyvPoEOciOi+OKc0wNHuUX3s1KAyPlPDZElclwkXTgD
xluhpqidp+4OmLUZVs+Cm4uInSosWxKdJ1CTgHL912+IyVectBAJkKBP7vDD
w+bpz0lUNmQFuQmOZhizCtF/2T9Fxt9m4jK/vxSsNznb63Cr/Z3g5/bCSuZq
ZhYOHkrqfAkFlWWdTEB2jR17+G++dMI1IN+kkqqpDW75bFjfOaWmoppmjf5S
khJHc1Mg3fY+Dm/L5H+2fwg8jk2WTSx0x/K3yDLxuM59B0pynUMzm66GpDxW
W2it5AOTLykHtBuvKA5qu/pBCXdvqoelDEBGnGqdwBJZD7Njb2C4anqQfC3Q
DJ3dGF76LctnYPVl4KPXWRN726+2wNbgxYOGEXk9y4XPVebRzyiUga+aqE/W
ctTsDAiFbB+iu8K/lfHd330NfqjdV2sKlniMQXQ2ZOpyXDwjAoR/ySJmi+r/
yzw5PHZecKxiVWsJ2Qkkw/eMuTLFMiY11eXC9QL7Fr2MrMr7jgS7IPPhggte
X/iYRnSzeG663cLD7LGubYxvSqvVuHJmNGFyzhZzdBn2ZI2YXseLnSb6do5+
8oSfG6VZ+QI4Ie6x7RAEQzhgRbfcdqOQIwtvfWN8UjNz7Mljxv4Kq01W5rgW
IuuzVVBnVFc99gSD0xCZ6qf+UtQy3JYmVAFahkl7hv3DqA50vUcH187ZKVRQ
CJCcq4LxNvyD8N5aPIvaJc+8RW4v68Imp4rTkZ8qrEa5foN+fY6fJijyHIXj
BsnX1bJpkVRWQF4bdvS3tQIIraoCYgh5MC07MaC3Iqaswxtz4EroFdDXdeiM
SWDMOl8RdbtCj7ZXsC2/yQquyNYlthefpklUJ1oSpMaoojjlxaXtKWyCZDvU
0a6hIZm9YN//gJi+6K0RdrZrW7dan7Oaw7RokZDSSdGFYPAhpgoe5AtdvkRo
RONLL/2/1iidS2hS+X62Iic3IlYdjO3eVlwhd4+5dCNCQw1YFE7eUAu3RTXz
ydb9iALnVhVP4kQmKAdfDX600FERb8ksNwPShjSEcODpmgQzo9YPLCQNnTWs
is8eVzBDpetVlJjzQLoDXIazT3nDsBQWNdS4aMlL3Gs8+NBSsUduKZB3mshq
yjC29L6A/1rHatFbBJmo2cI0kjOqYe4bX0AA0W/F5XZmfiiwDxCxXE0LJdhQ
POsTeEg/U3mQX1rI0RC7HYJQ/7DkGr+P2ZNklyjSdnVuNv4ef121SNFdt+xf
teNoNmgWsF3runZQC6KlqmU9GE5npTz1QETUu54u/1b4ZxvKBFdaooPJsxnI
kS+rbxPXtffMoqj/LXDzw7NM7su1z5Qr6YePjoMG0HZJ3WHm9sGwBSPnP4VA
J21nAzTcfHJDf5pJSXcrjl/e8bQoKdloM3lmQvP3oGFadqcP86+Vsbb2t2Ul
gr57HPefGWnSYEHr/FWcEemDzk1mGAvJ4ylR4q/stmZotLL9owZBBA4Q6vwo
bQ8aZ9OYXPzWC9RJcJq/S4p1ZUOVhg5Vt1/uZWItlTlCOSq8XNJzs3QNql3+
XRUbppm5VMJXFBxei/0miCC/AlzagnGwqbiozcGNmLnMC3Lj9HwN60CjET6A
Yyxgi4i+dY86ipxrUqN/aS+WG8n40jw1bClHeujLheKvbQcS9NCDFBVUdmid
VNauVhr3gBvagpSxR9jsot7MHQHxrZkQca9Ols745Gph3EskuC69pOApk3Tk
QaLXQ6tJqbjlAZdG7E5snhOCEHQV77e7nf+aPTChqHgXD1cSRKJIcDloUOKB
KGL3s473BHFXQFESOp3azvfXRIC8vom7bP2crxuF3hmvDrg9gJHuhlDK+byu
DuVHM2HL7cPkRh9v/qUzURSh8LsYZ+tRq5kujYKSYWLbNHLm5MZLg0Aaz98E
mJC78AHiqFp6OHpJV1cwkg6GlRecPBUegY0Hyc+P3doxp5aR8xnxyG6Ddoi/
3LgnyhPoRmr7zW0BZ2etkbJ/sf2RhX1ssqV5Vg3RflEYwEQHNQVMCAo4AzDa
1hb49BOWF8+oA0trdbLDAh89r9/3CNjrdfuqbKGGOdrjOeAPU85njLTz10M0
+MG9JiqQ6yAGf87XnbreUVRjqEO4L2FsGOvS65bz3o/Bw26+QFCNblUGX/EK
stT4PZbkWHt2SrHjMRm/UNboXvK3ZagZlyYOQ+FqmncwUrgJbEXITHMj20hp
HWYANHnupKj4HOT5gcs9brXNznYmqOinfWD49FxGeDvswBqXNGtQpAViw5hn
KsFrfBtsuvR7TEmk3H152PyLTbStIKKnrmPg3ZLbzMX5JY3tFVFNUYTQh93w
a0qK0vnSN+/orQhHNN0wPDVugS+Pke7XpYFC1pDoeT/cvtE1OR0FKlo6jR+q
VAOaU+C4eHzoBfzCYIBCl9AiTVF8vwM69K3CIxV/DU50Vg1A/mw/Q8FyBMQF
5KNWLrLM8nsGiAdO6iKQQ8gZqcAqOS8iJgvhVPjdWYMPPwTaFSnFePW9TdSG
VSfQjk4dTfZLtl0csK7LjTrH/d/PtCx44anBvj9EK9QMskbwxkf7+cRQMWlB
P3LKXZVEq2zm++mokCjPJ064wZY1zghZ0iOAFm5vBc3hCaTvD6Jz1AFALUzq
H3J1wSIwenZbnDX0SkL8KqHLjXJ+wSoQpEiZlj1iBkHw0P8iAXi4+jTgHp6i
QwJrT4Zze1GLsyfR4BT7giQ4RjPCeS3iuErPZnWaTIEoRDyDZ42/NvO5+O/L
rOnMqpH2hHcwmrnI0IBk7K872bIC6SyvJLyyofBv6QoVS+CYigucyi/ho49f
9aaPH7zC+O88xhSYaVwFxkWH5dO4EYNAXPYD3vaqEwNGUAfHXh43Jg+0/Mrh
I5P0Arkr/t4V9XeRc4ESY1PMTQyte++mHRHTab5ARBwzAryTnbLkqKQKfR7C
boq7Dn9PQUjjK6weFosuPwWfHQfztD1ldp/wjCYr4ieDkZbj8MZamNHHZTHv
YHssOj082Pj0M6vHNw81w144couWXa1lCA+2KCdX8sHb1Y3gKn9mvDZ18Nm9
8gHeV53uIiqfsErPGwturKsWEm2gxIPN0wmQbK9cyfsymzX8U0t1xweemm9U
xi+vXSN/i2H8TbLWY8nsj/0ftUs6yeWIBTKXANin1Vv8G+gd2cZutHmerXVL
8DgJ36qma4jry+ho66QYfQI8Uteh+trBtC+ROmNbExJwwKVpWjtrlt+I6KXU
Cq2gghNLDis/aWUA2yU/kXVnT6vXI/fmsyzkMhIMqjzKdCGso3YPvWbcm+O7
cr2FCdd3WspGmsTCgLxYf9zxBplkry9lZeni78L5anPe2F3H4jZ9oRT1mazz
Da7qIoi5z8eV+jNwDpjcKrD4QqCuDzL4dPJjaoI2kUfuon+YyDeyBYrPK9fG
6ETvRRk3eb6MMMRK7GvfwfMGoRF1A7X2bQzP336TJpnz0NP+1Nhg2/GgLSDW
nSpZKTARcjOS6s8g6H230/baAS5HMgDmWvP8/Y/Xhfa8qgoqG1WW/I7q+Fkb
VhMAAiDwCe2BdAm8DFl4/4BiwLAuFe3wWX60kLXKwB0cWNPQhARyMM2NWLMT
4wpE/OPzLCTUfDv2Cvg7CuRvaz8SF71YN2U2rNC90PUk8QfqXgzCFinCWRVs
5LvFsA2tcfOnjvGgSASQ3/+rHNtq9YKQJkxlTt9t3Xj8CfheBFZyZQ9SqUEA
VefwkfaVUYvmxnYszgnmvJHsNmSdXAcufaV38h827PTgFJqgWDinD+tci3D8
Y9dgjlmBplBH/QKTHDA9v/hNtXDDxrzQ1cf4pywGIfgdXy15cdrFXkr9uL+N
1ZUdVvN1LKKEJhH3kytH5RkWVYXxfXqQe9c2I9GwWwhJUXDaAGdjcrz8EUKp
naduZStgL6pX9EFR4LXoQq9RuaXFlSpgKopiAPHosYML+3t6xCTbk6axJoqE
d4iF4qqffMnIaNo2YSFP1m5+k8WUWf/svDsd0o5fYVUYVLm9zSTYLPKQZCH/
tJwj3VIssAKtOURvLx+6y+xYqcPUozvJa8f+ohSBccWO7raQ0t+Lkt4EoEvP
O/Ar2UxLIYzJC9Ou01Wu4WSnUWkQ+kfxC/QE3hiCDGdgq5EGREf0rqxHZ99m
3Z0eY2EpBU4o4sW3V+4uEWmY8UeB7i1bqGiSsvqMHb8FO9KovciUjv0Qt9pp
569D6SyWjhcebks+I1ozQkvADI9tL8jAAOf9GTUH3+PcLm4Z4W41ipWY9s5/
VQR4pdtuJr1j//cGXmvb/DJr/OBJZ/r8sNwxTgBdRUbqpHFaf+kgr5wLvajn
4PIu2phTJokNNQmX5x7neC80Svee+0yQKxzI/M24NkqCbwiNeodBxtE1kodp
6bc6QPoHblT8Eiz+i2wNhGordw/sVzXo9F55DsPd7K84ocOruiowwDNCT755
5T3GrkVZvkUH1N8I3lKNLgAuIQ101UT0wF++xF2DlHpmuYDXT829pMkqLW41
zZvZtOuNOAArYBQ6scEPP3eVsE7SC7xHwR7Rklx4r2CGbTyVeERp3ECKrCnY
1YAoeD2NeQHRErK3kTVOEXtH1nOcmGD+8x41f0MOGlLspxIXaqngXEnMZCoH
SkRudahk2ca6EvPVRaYnPymxsikGjKeIU9Fj37fShvlPlogqdI3rxX/WD2Yn
Wr3to7F4qMbtz/FWOOFrGPPai/2UgIo2QOf8sj6hrVGu2LHHPivh/fy8jZ7E
8+YJMEEXooawPnKGt0VymJhazROGHdWv33tJtCcy7i1lMpmJsJAIV/bg8hRQ
r5G38NVRPHNbLWd+6SfTyZRLa0rVIz3mGSHynZnVS/gycruL4eN44y82dXaI
6Iyu4sGvm8me2RYqoD/1jXfsg6tzr7Lh8gQnPsVoubHBdTwMX6BjN5WSMknJ
TWVs65nYfy10EfAICkhof8M0qdjCZR1vuNh+aHxCtTi+X+MO8Xf4CH3udISK
WeuVbqdm5rKSW8Kys1QVgkgs0eDu2c8vkY9kPI+7zkP/IKea1e17Svc6cnVh
EIzSdKTW8xRK7l5UQ9mkchUDSbwndB44EnLYT1GI2MMRqA4jyQmj+cwgPSeS
EQb0b9ObapUQRGP3FYCvY2Tj1iq2iVm1oPYiKvVoeIGgId1L8GK0pJnTQ4PG
iEayOavMR767Z0ALvjlig+zDsTHyNVUXKhQ7BNJG9c3Y4USkIFK1WhhzOqlW
tYj2xLfCXbHUIHG0anM0xgz/oGKy0RYMVROw/Nl0BP838Y3XFeqTYv4O+zuw
UAJftQ3qV7DJF1J0/8OThiJzgZfAMIY4WpsDWYVChOJtPmIDIswMPOTaLT5N
NTl2uvWiVZbmKEBOUHnsjukpLoXFQUnFEGhfFFCDgUyWgNMT9LzwmS+2yI8M
+plHEnZGnPAMB42X12loR8E0CagZ673xsn3dnUp1k1TuvxMelMrtWOopMZ4W
bVGk/TmaRoCmoKIPeBfhbeAcRGHYsdXrd2HjxVZ07pb3f0WwEEar1prkkxEI
mf7j3cza20NwiXltvh6UKUX4fBbOuKpD9lBoaWe5fiDJS3+iVlrweiMaz1ul
kVW+fGYXvobQOH2zMkxE4WNMD0fr8e6SlVa/UW+hKwZx7Dup44JMAbkVUvwg
NOe9mt/imvlrzInysg+hKmMlqb5XNrjUg/GLZty3ruCI0cQnYEIuuFx8fLOW
9lGsEgiJR/IGrnCia5/6M2ZN92HEAh0YKiUfyMpqX+dfTXWZ/62kKLw6o8kn
RaHZDzcfRgdtC9HsvV5ELjf2WHl2S4pAKUIJ3/GomaZe0ahSRtMtjWzef8hZ
Z159AbBCCgIOKF33DDqqDIsy8dMQMqOq/HT+rloP3b3avBQzBRGCyLqcdiDu
hJrrl7WfTI5s+aLbWWhFjMzQZVGnKohz+524KjRDE95VMJ+uyy2u9RWWVwPm
TPVb0VUZ9TK48f7FT36T8lDQ5pBy8P4GWFPL5h+gpLwg0PgoZksDrV1DzTxX
NWHrUrdbNpho8uDnmbSFpV0UHZOKm+hjmOaQTd9FmXlJi9y5/OVnZ9vsYjm2
NuAIrwvaychIfSUbyx2NaqkUKpyn+/EfkzPUnZkeEhf7u5DEO3TAxNyUOdt6
O5IQUioXe5qYUCYdm8EJZ8SmBs5/xkY4xUtyE/ywlj3F+oSvf1brAu79ASiW
Oj5h04bZMlF8mj0h2f6sTY+HKWS+A80DhK3UP6U3sjROwAxBYcKz78Rdf7Rb
/GZg+uGQzyQ7rebZZyNgs3I26iP6dVeLWwGRynDmDlyr8C+/qu/mdz+yi9TK
CLK2JjGm/iM+hzR3yemrDgBtd4duo7yiX/xhJAppYGJk80zuHNZtdpucLs5q
6+yPTGc6c0hTBWOo+nBrulJ2FUU+BR7LkVsPbHxxWZBf3nOI4R2PjGgP2/+/
ajHGZaXSGZEEN50qWINtvnfHefmlbdb3UW04cDT9Zhc/8FFwCqJoCHrzqAre
MZs6kncV/Up0zlgEq6Q3czuq02yxR/pX4bXLbsX6uNLYlTSiytDUdnGmcBYa
NhHcICv+fWuTjWu2xxFkcN6404+R6zmE/zkUj0xjgsF6LsnjuqCHupplzZmx
icObEmeN/Dk3sYwl9hRLKcqhfbUals4dobpNXvIZoJa9GIaWcBFkec+UUXWq
hInCIBR7DVDvl4aCcPam2TfbWbKlWbC+/tvruz7iKGUfhhqY1jQVdDwEufrI
lHXodKqaFKIfmAnVIm0PwOFTrjGPvzteGlVYGNcNuw5Eu9R5O4dPsKt/Qpct
BBRO9xo6KCGGswC3UnPeUqFacaC77BXWQhqmSIHygMOgzLerjcxySfb9cjau
1Ym7qPZ1iN2OGJlfrnXwn0eywgBdZ2r185OMJskUdfBZgjz75mOLBFo42FnJ
8xopKrRjePW4Vl6c055z9Avx/Bgwwx5lF6Mba5GMqqNWtx/TJ4ShtgDqUN8Z
V0Yb9RIPJw7nQqV+KIlZrOTGiQqQYNXspss1uvG+x2PlG7Y0dUHk3tcf3lcD
C0A+8QtjSVzA+NjxCssG4i1ltBoSPtbkFCULeFTxEvs6G3NB1rIKjrsp7ckN
7w7o9ndg3Y97vrri795qgtyesls9VYt4IazPRsbXkBXNWso2FYfHtJmJCfJl
8AfEdjmQwSuE+4e9Vbqetfiv6HXcVjbz0oD4JgF9JJcUobP2rb1KuTXndMJM
BonHkQue52G8rs4jQSVYPAVXcz7YqC9eKCq86eyTfCvc8DIeSXuJdo33CiD9
U57MJA3PwODXMM239b7qwm3LW5CunOkH0E+I7bGEzlcgnBkmUI6I/m91p7ft
mSjrldPSqDwhpwOZUGw/kT1LeGFZjmfFpJyac5C2t58uzBBGj/GbjYlxx074
FE7BE5fCfSfifb9ajoFg+tb0Of486X7BfMD3Hs7LC9Ug6gc+JTkE07lF0Ykz
t5NqZxgYvgIelAWiQqxIVdFT7VxuDnwzzdTXCzJx9zMeBIrPiGy4p4Z6QSzA
+BVhDcAipyIQ5MBvEA8KokB1Spbki9LCYO3uwnQLyuqVdgZm392E53ZSD5eT
PVPQzy+hqvAIwFknPsIAhkWEVHQBNWX1dIOik1815Qwv/xY6rwyRC4U+h1Kt
pfNjNktrvUnJXfacIrSL/UGi5ioUDHuhqo7g3oB7mOsO1KtkSnl0tycF4GCg
zMHnfv+N7Iy8NxESaQOZLym7fvyKLGe4uvYA0LQPvukmSnL81nukKiM8hoti
RMhKUDGJau4lZvMHFsVsFbf4bEEQcSnYsCo5hEqbwYvGzNDUp/3Fqd0I3LFs
4ERYLboA+ofneByYwIGi3TazZP9DYRD9fi9U3COkI31fiD4R5C584SjpGQAz
wE//xpKxvrVLgJ8KWCgr1RJRBS9LtySRCU7cjS0yq6aVkdqm2QrIRpWSuuW1
nTS68HW3lnV5fP+jI6zPC2Xg1yVDkI4b7lGPXzh59lM0M0aVFHNeR4ZfXBQt
TUbxYkDIw/Fu9GiLkVuA5mXHWuGVTyIPey45KVKTejMtUkvvIn68r+SRkCr/
wc0n66YAtlKD6G5OQut7ib8+6DldDJLk81k1lwU7oCqf5QvB7YRdpANVQZ/4
++B1sthJx8gvd/UfLzVSh1WsgMpvNrnMMUgmxPLhGUAw4MBPyjkVdrMf+xyb
WzckUGirNiK3LFUJYutwRc6Lm2lx3HBFHxQl5NZvJiKXZo8bCqx5koo7sRcL
3zfh/Av6VFnhn/fcvRRsmcL48FAKQZGHpOAs4clZ4Yldu1ygG1JTQPJeroH+
8tlTh7VmnTiXj+6Rvb4cMbLqtg5QxOksMRJ60qEUWb8o8vypauF5Y5UMFSk0
tVy9P/5Pt9GTSeUayuOMR9g9qxlwUzmbQjtsui+d2V/z3KUqZwfsDGj3+10j
Ae6u+K1RGLDfdeCwWWQR+c1N7fkkTr6NRGhYL+V4UNL6J+1UkgbIPMC+vSCR
ogHACX0pr9PxMZRSCu55O1KsFSFJ7DDyqRrJmUmEb5FCyLKILLuYYxlxcr/Y
CZyHvzYq792wGjjLd9fyyzl9RJCgfGX/yeonqfFUQLBQZyMEJ3Bl1IqRUvfD
Sw8mHtLyCTYXt0O/Dbq17ytoaRczAAbvcZ6A/ow00U1bPEfbVjWnGfYSIhHz
AzGAtA30a4TkH8LRV5SXp7f8ZDAVNemrruBBBL08yRhDjrajy2KNWXWOONJj
LqROsFZSRLeCCeQPyIVoNAYglNVgNP4c0VV/0+pPq9ShAZfGVmY/HnfLeL0Q
Sg11DvnSjttsWB0giDBw2697NDwcBHzrOoerjphQwt7MtoYNkWWent2jl3Bh
kD/9QdBq+7MooGflDV8+NUVcGzy/eDwuNdt0ZiR+UqTDed1Ts1VaDilCJ3sW
Ekb2dZuRmF9GUb4HWmVHYsrv9jLutHBSGoffq9jaiHD9QVHhh7R+nbYl0nSK
uWFnkb+MpFCOl1+8xDprGRKpTSFap8KM/3O7bIABE9O5stWwa0i9Kuc5KY2E
GzA0M2n0IgUDXn00WnWotpSm7nyodoP84gWeNb50JIiZTzGa/22Sgu0gFNME
DPF4BbauaKIG+kJ+Z7VmuU9Sa/2ItShntf04L3Uj/390B/6jm7MaspLcn3d2
fwOdeiGNU4H2V8ackaowreMbt2gn3Kg1D9InW3Abd3L9viISTOYxO8WM8XOA
nmH6RFwlbi7cCvILfgvUugfPL7o/kRNAntyf8gq6n4R+XylezUcvwQVKNMBB
LWmdlWuH11bRJP1ucPf2nDIUzpqPP5ocJSNCsIHIqDrbnbrBcPz62bpnZxV6
6bD2ez5O2qzAmAioYz3H/5IPqAq3n51LFIPG4jyXep7MwXOW50qLKy0PTYL5
/P2nfKmDScHK+RlIH4s+uCdcTeiTB13NDKDME9gjDA1ExGarDv+5itm5rrdp
VWzabrZEBUOVDui+VC1KjRh350SBr1xDRYaC4KSSKwabPWPf5MsAfNRI0TaW
22Qhu8yEP8En/6hqDnC5mrYsXEknm8uFe/N1a0QVe4rtq2JWdJGUxL1/9zxF
o1asYBOxhtlI028CUMoPbmi/Fruz9+2v385Rwua79jgctHO/qazxJXoupmQ+
5rbjAVdxIwnf2dx13n9SssaflD5IJ0naSh+ZstrBPYqG2tnUvmIenDrUgL6q
DPBUoqZj3ktUXehpmfYps2m7LeU3AfG+L1hP0vviFm7XxNudd/tgcfbn8e9E
kjDppnZM7Mjqpm5hsB48vuv6XaTjUdpYaLWm8Z06WOI41Db/L5CC0lRL97Nd
1CqndM/UMzKgt8MN8oVk85wxZEkW8yYMPfSqiG6FaL+4KINBFAdQGu7mkI9V
NC27iYoxEjqK22SQCTTze4DjTtiJY4Wx9KgX8LaSX5LxhnxscFIeldrKBwRT
zksUaDBRk0tONOuW8RQUfAiG9wzm11QZ+TcOXllhtxEZ1twcycZ9OZ313CB0
uDXLsqcIQZKoqFHdLWFaDRbCrnUjR3Th7nvR7Pjrbbhk61v7GBKKjw4l8xtY
bqYcNBtiigLXNr7iFRK2ciNLW9zXmlR3k8OvkY2ApOyDyLEdQ7EZo8lXLK1m
dxdn5GCjLbqFT4CqC8ZDQGhYDEIkwJUnA80f53/lJ3d8XFa77a/Tie+XYKqe
RJ0tmICbkcJWYjXJ/YoMGvNXYnrFBAn7x73ZWn2lWJw/Ty/Ko8K+8tpyIeIe
Css9LBs4Rgn/2fTBXOrykU09IukkwJb5lLSnWgZ7T2Ui+p2e6HBnBvJPkvjm
Z1Snry5sLeDwBj5AN7mCkG+uVTP5GDzWPXfVLNmlvBowaU/tl/geK5PhztJh
qT9XonoYRVnvYONb1f3JwTym2Nb4MWy8IK/OVXRG2tvTnG8yEglzmzqvUoI+
pDBPjmy/fL8SnsbRykmL93qgG8AR+34JGwOPRzR7zrEQZLGu5LhIqBUFAEys
QEhVyu2Fo6YMWd28B4wE05MhnVCN7iN/gvyGSeCLcYSzz7LqWXcptZ+e5wXv
MzJ+PQB/Mdf2IiY7qyuVA4lsHuuFR0wWCk4rXiZXD0vjvKmv0tgwWZCaGsEs
mpQuozYKj/Rl4ippnCuEmVg0+hPJ3ZKrSDGnnqRc6bll+GPRrsyLaJckgnbd
0oG5gdySDqVbYGuP7vmZUcTFXHlnfXcESeGNrrLqdwZ355/cZMUexE0fmh7J
uyjnlegHmLaTCWzAWk3+oFoltA3JOlb/QsCHk1CBlwauOFfULdWvpHjrXFDb
yDt3XONVmZbBc2ffHErHBJN5Weh4GCOPNSyWS5EXmjWvg524f5q7FHuk855d
TB5IKbGtZ0id/9xVSprvI4+MMYf76j4UGztcQnLmMP4UueWvVp0bsxWTd7WB
0VoUtqtYRl7f2+xCAkNC2Gd1xM4C9iOEwHHTTUC3jaLNKIanK3HBukNECTrT
cweEQnetGvVCB5UYNn9CgsKQ8U2kK/YFSqnKkmQNJ/cGTu89Qagt3CkQ54Gh
gRafpEgQhbKSTVYlWH6MN7m1qk/XTM28kOMThu8WCWXe+hLJbKi9Fbrk/SZd
+nSGdRshn4fAJc26iT4Ybg620yT2Xa/xt1cCaBoQiQ9f93uNjfiFmK4cKt5Q
LAJeB99U+0X12P56yUbQeJLKcBItiSdN8gZ4bwzw+2I6DAB/yex/nuCDsnh1
T+eAkH2EluJfOhz7itZI0qllbip+a8efnRjG5XUy2rxBBIuKmJ5TlFB+VP2C
PkXz2FNTWEEVIgy1vh/Ftsseh9st23VPOf5kSIpAdsrmEB/aWyudztAlicrI
jnWh/ii7X9zNjWeWln9gigUBvAZsx8p5ZSvXzPMnfVEnBamZ5raV/MK+k5Lg
1FZI2lb9NLwS9RszEH1JIJUuGB9AvYfqv5ahSVIpBUTrNGl+/ECGIrOcTeS8
vadtkb0Paupac8ThXLNtfGlu0x+qMwGw+H77HJIyyBD2PBqygEFZLcbeb3/Y
LAeHV5hP5O3+sAi/EN+RZ2NpiSYz3S1qOydyp3R6ZOuowvSZwZ7CoC/2DXwi
2tbIDUStxhInCUEm/P+T13TRH5WOMx6CFnsDVRCuYhgk15oaxk7HaLegZgqp
JmcazUg0cGYqQCmE2Jf8TA43gHOdqO+rwjoL0VItJM9tiVv1FqTqbSTG2aVz
YCm+kYDD3VMOsPvoFX/cGiJhBEXH3cPiaEiDUmyq49RpRo8D5vpYWtbeBkRt
dUEpxqk5OfucH5dqWHt8d/0CcZ7ZHyFLLNmP76o1XzknPEi+QhUKNStsEbqK
pPOklaVufr4MKdUaDGv+Vma8hCDXWsQ36abh4WRKsIf8dbs9scD7fWnklRIy
fVO55NW3MTNTr3X5E/Dt18MF1XNbW0R1u5A0jaox3qtkSJ9p9uZdN6hcjSpY
RTcyu8sZ1XrhBPBWZp7ilR1M7IztHwyWS/oE7jx43qXfoEwFnUGzCELieZF5
l1Tx4qBN8khzIc3o+n8v79Bf850Og+d4AUO7b4j6VpY6H69MlceBS5wVPNc2
aPEYcPMrqxJ/8JmEPsV5+wcx1fRefojgN0JQm+ZnKmyelEv5oUfNAPl0BOIh
h6dklacZVn3SqDGuLDknXQ7RRuU+9JS+PmLZzoL/IN6ZIaw2iu6l19o3ejBG
QyWCWNtE2ZaT63WHhbW0rwHWIYd+yEPIzPrYZ+UpJDtu6cswjb1uz9MHgQHN
8+fMhnR60Ni/w7iqcayNHSGZ5p/WM8iKDjgHhqi8H9rmtdmZzBTQM3GoBb8L
Um+Z2rwL0pvIiN0nTcfFpc0wOo34j9JrP7bYYVzzWzJaZ1u8gkNWgeh/IcoD
v6Trb8AdgGNS9grIMCb4qz2bNf5ruY4Bj8g+h7N4EezPbJAT0EBI9tVSzAoy
2YWAwyeM4Kmu1EfM1IlZ8+DRZxZc7XC2NR9/+qh1RE61YIrnnbOUmTNlNoeX
1hQghMXjNucCclMtRxH5MJ8HqRH6MSjcZkv7go0a7hwiZCGrotyaWk4x6w54
79+XPXQkTkDf3LULp/p6PyISK/SrgVXyQ/kUuaIq78ZbP1+HzzKaL6v8cv+L
KCiPOiXwXD/1rXKeKP5jitZ0rJ2BRJ9AWil58pwvtArUhdRqFMvIdylSlgF8
pUX2NjsOeTeVEC3+5DBDprS9Vi1YFpkS1pUW0bB8XBFgJTnlRjSbb/+PRF3h
RuWqMQIKfkDNJTSaFoeXqUdLWQ3GOj4ELfasG8lnf5eMHb8PK/053K92TIZg
M9rbmvj4q8t0Hvx4yckI30JHCAo9jvU0kPl2mL3bg8Cst1RIREZnrowfKNvf
0mnS47qrm5tQqmTSsf/CQUsQoBvNumSKu+REDFVkbdPRDmUwb1MQs2RzNZ+M
Y2VZliZ6QCraFc4dxFR8oWvWQKRLN2YTZjdTfRS3TAoY/d0spUcHl6CIsCRA
INJHCqm49Vbecoll2Zvi82S0gEiWcHrAzlAfSbCaOk5UoU+MG2TFGEeVCTT2
JjQg01Ep3oHAlCVK9n3uAkDaYfqHCkwkDyIZrAFndvn0yk7wrWgbap2qXMma
vGA38PS6PI64vMMOqRWOfFpxjDPNzbgK9GiH/E5wr0UdElf2jRfyh1U2dl1f
EOL/IkWn/unWtQAk+JZuNyc5kqPc80eNrs2A3NuvrbsCciQxpl78lGm7uoXH
vWv+/soMtYPB9SYXjYJ3iEoz0w3eiyRRXHLxHZwqaP1C1pRYdwgNWXIjs45m
0HL7JCz8XMPCvV0sbwRqL/LXcApKlhMtjR2+cRRBb7Ca0SJ6wZIsMfPxF6Nf
HPgbANTBTtsPrClxthkFdHsK3E1a4mZLe9Ocl6p1++9QEE45v0GH5MSAINVQ
4qQmBs9Se9ns+e70tJKAJ7L3gfc9NL2NAMePwD95ul290uEUosYBLe8HmQEf
tWP8CbmsobqMmw8bMitljGdct0DAtkEAsPTa/dk+1s3GnNGuJHFu9H7awIiy
LM5UbQVWliN7Q6PzL6rq1S0+6K95cVtTPrtb2AFqMGAb/YijtQZUF4SmOV7C
I6TPHfd0PFqwmhvCSGpcUpIbZV869URYCEXdGc44gn+1rgYNi8vTLph6cWZ8
2o80geWUPK9Xk2wkinAlUE/LeHII6Gs6CNHbyIYbdHcQaWThcBISsNkevP5G
i3AH2IsHfpTlK5CZsmpxzNBlBNdc4Q6WTmgF5M7+LisZYsr+GeCbevY1m1vI
QLK+CKAdaF/5fyFZWxb4vwITBtsz//okwgA3A7oDNxV8LvFuYlppxkJ/eZJI
SQaVBXyZmqszKTjLQUtQP/bvBAn0IizCBPrr3vMwlTN1LoaJB0YW3v+OBR9Z
89R6ilPhny2qfBqDCXbDtgW8iEvwnDrAEJvwiAFxCKzLdVhr0cuYBkx7v76P
177NLCgQ1cwd+x6QKhTnMfDC6ufGtQsasTaggiuuzWTIJC3q2zaoNdrw5yiR
NKhr0s6ppK/wEolJvLRo5VIAbshpOdSgxesLiQ+eC9Zyf0wGsNWLONuMGMdS
FbpJrsAqjaUv3yMN8gE3mykfwRWiONjz5YG4gRPkfppLcRzhn4YVZlBYww1Y
G36WrRFQxadnB0Ml18NejC3gfqIbrtmf5w56M0GA8ea5aSzf1dquk1Pc4v0+
WkD3Ko6VM4Qcqw6Yfb3Q2Kd1JEzu4+gBgU+dQe9aborAAftfRIBYd6vyEVC/
KFax2MCsdesKtd2OCZauhQ5hfkdkB9BGcLT3b9EGdT1M+Kj7KOjKxwdBk5uW
hndYyV4EEifNx716mdivgKeXrmY7vml1HJAlIpsMUkGRXMnq/BXF4Pz9hT7K
LaoG2BWuT3PNCRaaY0kmrKeKtN/XK0vU9qLKoRJAiEKuf8sE3qA+1md/I5Q/
AkJNsvrzCl6zdcmFkDe0rwpnOuE/bt+nFevh+CEh8ZZa5f32GalNm9dM1XPD
9ikrkl3vR4gjobMQHXf4AAgOVcGXpVj7/kgHk/TL1sMt/obp5xtLSoYW9t3O
1OLJwJIQ30Z/4yjMou1QeXITm6MJT/0X0fqodDICPM31yx1/PxfEYtglIELV
ovncBw2UeNcB5QNRsv5dkILh+PW1iXBCMCThZ21iDLBq2yWSzF7C0bFkOfj/
BbN2F3bOiWYeRYIvdYbP7PYeRqo8UJ+Em1OHbrfy54gu3OdbxJkMbGpljl/U
nXPFTV6nSNt/dOTL1NTmvoMg17rczSDAPJg3Aa1ETw8hrYrOFF8pK7qrBFwL
GbCVMh0UaRjVM700IBYsRkAXXQdDcXHvMnHGL3TEFqejX6m83Wm6ORW72I3Z
RfbzUQ3PRzDw99ruGAwDdhf75E0DCu0nUbjsrMeVD8ar/9u1HqzxaCoqWOq2
THC6n1Vp33rf2tvY02fDufB+MutSV0NaZQhHg/HtvQhGcY9w6Icm36OUk3LJ
A5eTZxGPgKVXuEFuLDJVuiNz6Tia97EYFjlSI0uurK+32Pztjl7nELuD/Eda
6Xh64xuBkmE9jcm8GThRUVcLS//PjTlTDtuiO7mzjPbfLfQ/1wnVw1E2m9KT
34IxfYpAnfzczh+DPg/GyazjDN21eGEFVqp+LvQMtEhGlVEL41gisV387pW/
M3qE0OA5Gk5GoL8FL03JpeEatVAT0r0u+8M3Y7q69dBUjoGWOntTlcmvOqfe
0TQ1zMiJ9QFTz3Wxfe5tOYw7sv84DmDxJ6ldNtesL8b9iiiYyjth+Xn8uCtK
OseBLfH3jqM71trfFibbZU6bcaIpoONO9jAulRZXKsi5tdxFqTN713MGOMqN
V7vyXlolqx+HAbEAh5cU1dKBMM0+mhFsDTorvO77qSfnaUdfHVtX/z7YJRyx
y/CSOxWkmefEEaw9JzwanllHTDL3J76kVito/7/y4ba1JOFHPmrmDwDuWwpf
fFzz8MoJxGnxrndHP0pVRGQeb8Q+snf9paogx0KMs24XsaKi3JE5EEcvhVos
fI5gKLIBVuXK0oEx6bx4sv7frpUv5j97hlMnV3R466/xROJJe/hDZ/eOpMMq
FirEdJ205xwoBo1jR12dxG1+nREPREAeiPAtgkRmCkXQdgVD961LFiZHMmqr
cwb3tw68K8TrxydAa1b5NCQs/HZs2r4a8naG/UwrHCYCrftJwqpkPoCydyIR
YB7xJnu3zNsHaBUdWv/mmM84r7NgylwnXK33U2yWIeBI+YwWNp8VjOAJQmAE
2NJ5+FR3z1RhtD1pSbcCp6rAOoDIiyYJUhu/+5eETmPEg1OXPBLDgo543dwB
aykCE+MRusUbI3Oj1NFfBFb2MjFoEm9gQPtV8Dk1cp8fJjqsYM6RPh5rQKeB
Hp9RBRO1MYEN84ttsDPakZ0DcGa8e5zcV6Kwq+ZKDW3NXyJMYD5cUcNmWgfC
324rio4WhTo88SYve7o1SYcEnA962AMb8GF6KzsRJoXOGDuyfx01ZIjEbp2+
gBo+tyPCjRyQPsV+/m4ghIxC83st2sKSS/yyFEpIPlv+S/GO6hgbXnzmT9H5
8tdFrRDTtXL1Ge+XQPyM5k2bGARB40M2oBwwPCbow4tNdPUHT4thBr6erCgx
rpnBPJloVm2TAVODxD5SQPT5Do7tszPAOUDx5TnlUDbnQ6COhdvm+0HZPnXl
CHzf9wqd3SvGUoHVDNeRa343q3OYd9jLxSj6VfSwyaJ/JVOSsPY8cNzoppFg
5pPHhxglXppXRyMVUtzr690AiYms36IKSdQP9qqOem/cFkNyraFk0Q4+l5o5
OVMRp8J56CbysjiB/Yp0u5P8+4VvDvtJK9who3R9EYDqKd8jYLuac6o3BYMF
jWGfCPRDJpDNhVxbF2uBF0OrVPsEC33NTAoF2EmKMz0nFp5uajFqN9SKBVH9
Kj4da72qLw/4HJrRG9J4rWwEBCxqiAlZ6Uot+MkOfkILfl6qxWWGrg3ZKkDW
prGvqJJ3Lgwk+MJouZhDxxSZ/lKNUc3Y8xTlrna2fUEHwnVa5PmK560C5vQl
5N7Hp0tqdgMEb60uHSxFWlzQGR9C5TtePYjDcClw2v59yKZmTqWiG12khIIF
OG8biTR0VFFH8mGs7HAA/9FviBrHOlZch0BC7DobUofDUi1rm3dUeflm3nTG
hFDPlwnz+THlO7BYjSjsYj+6QUi2KPCmAywl/j1X9Xv4wndsMTKx4eryT5qu
Ui78oPjQ2XJYKa1Lzx6hS3PLPhc4iOhOOTgAwy5IokhiooJn+Y0zUM4HUM3J
wwAgAw40iL/1IweggpvE9Qo4bC/9JP9B4tkLc06GG3XATyqbFrOS3mQpwZol
mjN2Apmvj86eHU+kAB2dxhkd8ugkdiL0Pf/q7LEzBkXhePaiVElqCfAu2tFi
QsiklVaOAeMYZ/jW6TK7wTIHttSD7TKLJjwx/tvpqhLM27IL3DP2HcXWJ/jM
3pI3ZIjb4iymshovG5b+UOflgWBtuUu4/KDBMXBgq7/QHmHb1NM3dU07Dz5m
ouN6Q5n6cMUWn6cWV/lFTXWqSfCH9Y139UbFeQyJ1MJ2u+vYtKKEJpPDk5SM
eoBqw8ufFfT4zJxwwkUcGvCgU7Epe27BVHdn5RPFjFcaKXGa7jKw36DzBVvd
ODu3kiQyZYKX/lLpdXyml7mpBpDmsEuPwbZrMan/XbR5qKbRUEsOHPsSGQl1
IoIgerd0zcv6yXDB46ICs8IY73DoUKwQl5EE7r/ZXEVPf9dsNxJaHXIHUBOW
Es7vtqw3n3fk8kycdxGcHoueT/5cR2qAd2nytQhHpiLB87XZWir/9pBhslZ5
kcyLfbKVevNEvNNMf0XunYBkvprmOSwOEBMJ2ev7pMRzYIGl57FbxIBYRwxg
PyWQqY4oSITQAD+PGkCY9Vla3hqC+utLkqcLd0UtMgUHtN14nM9drEcsJKBx
Tx12N59dyINM+wSh2v354uguR23BykZknbX3WWkjuTaZvspPPYcsOg8xDM8E
skjFo+m7/OEBoocMR0jcD79/JLQ38gSpel+hgI1TBELZ7igORmwLuCjiqjgm
035cnu8M/QEAEcqeSbsg9ukNiq1bqmEmtDWbEkNLNigB7B91rY5uy2CJ/aR0
KKluqLOElCzm0anORt+XsR54TaSSf6QdMK6jAAqlqgmfAcCgZIqrxJa2fa9N
BZMOF4MOBUHE0aRS7W+gfN3XGNvQhxPP7p0L71f91T1Txv7pcU+NJ989jgM8
RC1Px1Z3hvPcDzlpyQGeG2XTgTw4FiFaBaDZvx/61Re+1k8OUBj6VAc+GHhb
1+/szNpLslVNzNqCbgT83ut6raZEo52yUm0UgbpvF/dMGruUHFD29XX/pPqV
v/A4IZDaXwJX1A5MQFXaQLRET8k4qkDloa6xq2CDdFtd2k5cB6Jfy3qYQZdT
ET9zSVc3nXhfhnO5yiNh6qG0tQQ2KwXUs6c62415epTXW7z02CnVHpqJo/wZ
mx3A3idtIMPg/4Zkltx6glBl9Mwz4GPwmb91PIOZh12gk+oMzIzWPr57lXbT
l53xevh8vpBHhHKltBsJBSHgEpdmg3M+KMU85v8djKnFTn5vWHKt5eTTA9oz
anRI6brxmxDRSu5KDiLWVQS/kf573YItuOVxSGsZtJTxk6P88uVCXD2cd8fg
KNXrB+g9S0xhWbC/U++Cz25I1VbLn1hVXU0ztbvMZvwCj6RDDan48PF1MIGB
V1kyVhTIzJCxe41ORUDgIwVU9nt70539YevBN5PEJivwJMNYTaMDtry8d9Dm
lDu290Ot8kPSoLOmmyhJBpJV9P8/dqpR0g/IeJjPdP8o9Mg4O9TjH1HJ0FdY
MsN0lrmycvBq4Mwo8rkGnhFCAprt0Jo6aXN3kQ6i5uPMINt/p7vvERYnjvJ+
8k5Ybn7bwnmkC+HkDjzbTdoAWU19E5QVT8jNzctARP7ZPcpXMJPWyheEwVLl
o0YqsLo8b8NKtYFqH23qL2vmKVytyXXVO7XwUD/TM6Ke+5wnlYRb8oclY3uv
bbv+1Yk3XKFIuyt0lf/+TxUEbr1dhY/WuSKj5c9ok//V0bS8RrP8jhAKkQdR
2Yfb+nOq3bpaTGDdFaLuD5mx1HITYx3GQBQ1mO0UeN8CAWq87WuZ0D5TmNdG
DmIdzPMP7EWrnXL43RW2avZUHG3qZGE5d4v5AiaN+xqDYb7NlgFkWOsz6u4W
5ZvmC3FqV9Cp6yP9/remHDWMm2m06X4vIjhyV7JUWrxhcufchFkKuVQ4QPZB
m4ybrhwxXO+p+kSwdb2jqdfGSIPBp0qiekLF/EI0DFIG3AHWEJcdw4CqG5dB
S9foOSkFH04YLa/UyrGaxhSl0nga8+GFDSv9kE0LE+CXxWMjQWsI7Inwhhtp
/1ZNAA5Bhd9EZAp+s9nwgrPaFfLq6y8Mxi6lt67P5HKpDLdixMz2vhDLfDYx
NRtnWpgfDiGJhj0DvoU6ju4VUmPB2fZ9TF08NnjT0hQE06vtqdz2GQsCa9Du
gQ42TdYNix8LAy/w4or1LmyVzuWLrdJHPkBGapXGP8tJ+D0Kw37A2GSrshEq
oH6wVpNf+HdKwCHDDAmwKzSA970LLFIG64ObAx0+CHTv1PAVNDH6/UZZxZ5M
g4wMyJmHiUfW79xUNySNs15XiMlABqGPwmVP14Ry6RXL5Xp/E/d/jKeNTCWx
6WiHgNHFcexZSXfmlJjE9arlcANHwfBH1SvLfahemnXuYXqQYSzCN7u9hBRC
k3y8mAHaMAB8PJlGFaJZhEYp9s6SQRrr46YAnXyyqzZwyPkdRwvc1v/ejaZi
z6ertP6gvxd0fuIgZ36ptkQeavRQajuhUpt8Csc2kgVl68EeYGs0J9oFkVW9
1ChbnhEEp3XQ78MG05bgQ5oF6M1F57jN77BsVmqr7cIBPo7aAcRCsp+Ua96+
kT3jxaLAyWDEDeyuQX/Vd1HUNm27FhGz4mTBKxF0REsGzi5a1nc97ySkBYfD
meQqHrqwGxaO7j6JCNMX5CxLHPfRcv8JBctesrfzeEsadMjbDN795fNg1EcH
fn+QVGR8F+EocWTrYemYxuyAyLvxRyCs89xrsgDHQ3Vy0G4IdqYLPLvg1H/C
hvIJIpZnGaw62UXSd4af1VREqg/Pq9HFqfP3oB3lKIcqpTVG4DuIEiOXTbXs
6kQqHyRNuP8GyrOVIYFk8JimDWFO27aKn60YJrss99Rq+B0PRgHiIvYsZg5A
Zx0xMyXN5L8a9Ic/zMN6Kjt7BzXCUz/7HMBZfYuLaML5qrPynrVAH0pKy1lB
FruXcnCAcy2VJdXiFceoUYxZVFAkHaOmhfwCVuAaqqWu2IRcRRYP6rINRKx+
u6h8hg5/WoQovx6Ty5AHOrwe3C7wMIXAqoL/wqFHI+tKP+bbILiQpFNJZKAo
fX6V2sh+oiG50gKD6TE4K0D56yrNbLT75B+zqE2dFfurX266BO0RuK34uDDV
9IoqvpLxH6blq/rAvCUMe246IvaHCo8EU3ijQvVkvlHCjqq24DJLdUU7bSvk
b7ZL1qwJ5qgZ1mBxbEjlRU/jUWJqkmtxY7TBqcK705MH5MU2TUYe7a5U5W5k
DCnfDQPO+uaBBTmQrOWHXrd3dnVH7Txqb/HLQO/OQvf5ScG5n17R3KnfZez6
7o2RJ3Qv4g7pGIgvMofdNu148S68w6vBf83zwqq6NkASeXC0hPMp+UpR39fw
hN6hu1KB5qm9ngUNnKzdOHmfWJvA+vomsoywA62oOOMP3+ZLiUIZ7Z896+GD
X1Uc7XyiDrIF8Y8+UuY3HlRWmeJKEXi8ELmTVJkfPrRrxNvOPxEw1k1bXRe/
E4E6kCFySbZXBhWyu+4/h/gH65meDH/pqjHoLs3Ea91I5k+/Y3xj1O1t29Ap
g7ooelT3ig2WA6f6takqqA6Eq6DfCTSC7r01/ZcA3NBCQUkxFAxbK4d4B3d3
jDlmpapIeMjUZ0JbK923CJeHD+9wNdfVNHK1tJF2Mvhg85BddcnWahIHZUCa
gLTUhXG0wLwyBxK/c0Bl82WiIUJxxr4M5zGGf1pkxOWo5FPQl3f4JURWx6Fq
perHQrwku/DRBqE/9rPdhu0NNGGx9MKz48p06HN/3NTbx5RXkeRFTkbzdVv9
2Q9VUO4E80r/x2faRCY/F9RA4llylvmoqMtkW9erJdACQ1FAjih8N1KJQTVn
tgVk3isJnLII+Zlupr+7iW4D3+CBDFB3ZuvpNLxp8rrHhN7/KrWIHjqHxDjI
WxlJLyKoTO2Xba4QjapGkbBGU9tyh0i0HAq4nZmB0cetPZZ7frwUdBR0RRqG
x7r6atwpHhKGitUPue9f8BiWs2/747McN1RO5laZI3/Ma7Uaww7cyStXDsPg
knlgw8HSgYurMUxDbPcB8Pu7lgzEmy+kZtgQjYc1IuTHmbmEh1gIm7BrqztD
0R4k4UUCVZr4Z1cK6brIz/TGqSXwRevSR7oIowhCWw/fstiQ7jeqgtVmR/Si
I4Uncz5yyxv0MwWdtGn+y50g374NP/SUkQSpmr9V5Wjrp1+zrJq7mFXw2V6d
Xr0spGP8Oq6f6bjxYCHiWKvxf7FQjG35khIU1tuGSMbPjxS0pDyKWXeJ3MKg
hwcVSQSF6POqxvnXWaR4hahiiJ6TT8BHiIvIgJ81B6AMeYRjm+AdlLFccaBB
AfJsHF7C0eIbRURrKM6GlUDJ2g51mBSSjyxg2d0C2yrEQyTOIkFUeeEHmaip
omZh3xAR30F2G58Xy5d07gCnR2xe14X2sX3zoaSqiXwKSM1vKJ9kfXUdRqLQ
MJeds6XbKz4WISH8qyIGOP0aM9AuHb5nq4KnzjtmGbvZ4nS0gifDJsGCFGFt
Sdg/BF2xR6MoJ4/wVXjJbtJGsyRAs+S+Ia0AJUKLZ+kFQrTWOSJASV+wToSz
wvOCf5bqfav230uLt7Pfj7Pl8FuFkd/C2S8wjqQMYTQslCWd2IGCZn7aW0Qz
Arnt5UtfYX5+T002BW8+216NMDm8emwtDi+IVd1qu1fqtdqPxJr4QB7r2jQZ
uEIm6IIRYo44QpZBlDYSTojpIrWVIYZZ55SsPS6kvpLYpmXKVw1jPBJ3z9cZ
scFknRkfs0ygvu6MA+ecar7BmCWV1qymgGWZREK20UAiHqmLhZCWBms/WmSs
+E226lrr6BBQhw3qMwrOELs7Tbd+47Z+3nj7qlt7c9+8GQVlTepvz1ypdIcG
HwrF21Sb4f/vLXVf9KVF5ykgFL2Bdm5HS1F1o/cAqywoOwsipUPiU24v9o/d
SDPyfynzwbl3z/2gW4KBkx+aa3QRnWNu7fwUSRp0Fn73PlROloGk/FoZDU82
E4YRe8SSnX0LAzrdXoYUxhL/SZXmMJpul/SIqJ7Fwja1E746T4M/1JtPh1Jk
T3bBqP4Yit268LEF/Xa/O/MY7fIsaF6faj1j/jwczV3ZLpPzRLKCHbgpnW/+
iWf/s6+1YRnvEk8PYu78B86okeKsoIx0+AGOXtdbDvbOl6WBL8WEMnTYBtLI
YHhBhMB09xv54TGEPYOpU4rXaOxvqsn/d35tiMbEo9lOplSk1pMttePPN+r2
9WRhKE+pdVkTC6hnrvZCPvNfDoUH+G/ztf7XaowvZ0/8zJwqXrNL4H1DTr6H
iPZkXRJPosBWa9y4j5W5FzD4JP4tGSrTNQEdYodgnv6tEmhRXY/nDeZeHXx0
erZTA6xbG7KBiu5PG0JOoodw7cz1vhx0qX0D03JsbyKZDEpliqNtVMdkIop0
byuMz/ZOBMZlIg+2GmEmyPbueF8TBOSbffAksC0zH/YhyuDDnb5zFAAk/o5J
GnEdd/MZ4OAdE3DWqw3XtqL10SDxgGJLB2uq+bF3Be/5voRwjp7wi6wbY9xl
gZiy8xYv8XkJXxPkBrmrgKpteEOyTyO7JqsfI/srQlxC1Po3lzDXwEZDyyOd
ztBHYoOW99XwA8EDAnYZ16d/hltaYkDhtKkX72jMmwAypHJIqE9L1Oh9iA0o
8cmpWtKZSj1KvK6sbeN18JdDh4rhHy+0KOUDcI3nqr22EmK163PgoO3Rk1Dp
k2O802HadRiYmDEd1U0zIeIqqxmUP0WNW+SMfqxduArg2RJam9qLWEpkNZSy
/EwtRAlX/AEika2EAIKIAH5lnCtjpEAU01b0Mih3sfpLcAnC0gZpsazeZ0mL
+/zSy62MgFb2PbMY5YQNGJ60P2DluWuXWtEwNBdQTjZN5lo1yw5ka1+kW4Gz
Ye0JVTyDaPKHhBd7UQbO0o2gGXGr+DhFd1J49m4yLbpDt5TSep0pZxUBY3XV
U9nsOt002RpumL/U4TpE1P/dRPZUFO3RATkmmKRuEmpZZmylOBeA5Bhce/tb
evX4OZbcHYVtAJ8SKz4vZxOuPAAgSaOmSNbekEHZu1WpTfU/tpXvpB6tGsPs
88TfEWDutEBFRP4pp+CYOXotjmwmKph/HodpLKKGggMn2S0FRvbIVVnfGUuk
CBYScixYmB+4ADoYNlWs6AbCrBEiRhDvGm6ut2HYVd4J2kdt1x33Xp/Ds0xe
yEpGHpf9b2mFMTJY8X2ElsVPxT9DSvsZlkWPoRilrUVxeC5YZBxCcVST7lvI
OWu/KIoDIhyJQ2PiMiek5P+dlk5gEKL0DH0G6LC/oW/M3uGqOjxUjtR1V8SI
6kLJ5weS0BDhJzZc9loY9lGbRwlPytOSFaCM4fzmwC8+40p4KeAuqSJwRpQ5
EwVYK3hoX1M3Pc+QgtUKguM7gzZeKDpd5DgOxdFA9MW/CXyvWsQoKb9fC87J
6z1T6KRvvoEtz7nB+WBSPoS068oNsTlpaAiNYkwANKdmf8f+um5cjeHtpvgP
Az7/ZO939QgQoiKpv+7g/+sf6fKZGzz49Tt2n6EwJ8X0EGFYO/nTVqO/oR4j
v6UfA923zg41k/c/jwJ9G5iGDV67r53GgdxHzP0alyZ8icIWkWDgOSZKQpHu
7OjZz2cwcqQjW60trGGsVaDuxtuoZ3KIvmARo0WZ2aKNsyDZRYmL0Q0XVRqo
Zx6Hgj20bYkNbN6BGwchu78N6DGUAqLSNM3KQSjNCE/A5/EpnTMj5Drc4TZ6
O1yn3JyME6s5fZTlvAKbcyZv5AqegKQkaxU/DmpTUHGGY9xq79Ttmd7awvoj
Yoe6C+4x5bvTHGnlr7fSfNYOXxZZP5gzzqyoi0DnDcJtepglxtID2mCXdTZ4
MrFeCWMyUISMSvAlLJ1MaYlAe3vDGr3dbTbdYT38VlD8iJeAaJoG4OA9qCcw
nckCGaCQKBA1NACiYLZWxFltk/uWvBiIMU4xw4iIxL5GYHRwr3exb6L13S4q
ENaL6oSzC7lLTR5j4JYgT2xpmJWOR3ZCocnYSk2ma/7LZKYYUpnx3gI+vWNg
/k2kwZDGUeHWDaUTPeK+GtH0fz9SDuY0fjmWySw2mWxzNi6vG7Isupr9H7Ok
h7xReo9XhHSj5fXcETRr9tIG8/MxM15tMbJgHmFqBGwJGP7TiQ8wac6NP1q/
z8qjWsNDRnKqyb1yj7XpyZhCPzGNpFuLB8bbUsvz+G7w0hJBLBhCcjgVEpKH
HDZPCVdMTQgE2U/OOHJJeaj2zRmDWNaHxy3nJXQK2sm605pTAa0WOFv0LnK9
7LgI0jbOtoYi68+mmDrU4M2Gs7DbZIFthVpTRB0F//glMzc/EbAr0pWQ8WfB
XXEhqPnNUqm9bvUY6kqBzpRKzldrHatEN6xUX4sog+h1T92aVT4T+5hcAnwr
2S+x8DvPlPkw6NXomTJiHO0+IzdPRXo7JmkoV7VbupPY22cIsqB8c670lEj6
GJhZG/qA+ZaggAWvdpgKbLVKb6IeJqLJ8Ks/XrhwNjTxnrkYgGH0Fnz5Pupc
vu95BSXQCCZjZuNW/g/7OAf0thCcBzs5e01pAPp0DpVdqMXjntVvk6TepGDT
soFQ9n+cfqzfLJPwQa20BbbdvrwWsnpB7Ktsu4ykKB7SUn/t9LvOTKicXr7a
DHkTV1IwK/VysKXzjbpvPuyxrIs8CC4Huep6cNesM6VEwai9Heigcgyo4+3f
bkjfd23rx2D8qatUr+VQatXrUqK1WUD5HaPV5roSAmlCVp5lHTi+atN90bcE
FpsaNw4wpPwgwJW3tgXX59NXvuTKbQQRPgrIHY6H2eoD21RiZWBaN8XQWJBa
ynIWZR7nNijEY/Eo0ZA3MwEURcUyHrp2gQmwG+J4byF5YiOb+RtUw+wxhWgm
aLdzuxOCeR6EyaLHIGcSIvUPW8jjJFXTeZyoIaSnKGvzK+lD56lcJajGRM/d
8TuPa9ZUUNAkwX3zqYrwLLqAIWwopIkcwnQFsNOOttUWw1XH/5z7mo6lWDOW
L/4exZVptaxFO1/Qh9bn2aIThVqaBGa8uTdF8OOv7WsqiymMZWR0gEAqun4p
brAgDXYDuwMvPTqBfnO1e96p5Kk+o6H4VBGXLxmDTGpQA5KsPDxSmc6C5M2o
2CA5+f6RsWqMVjLTSyVJMgTORKWVaAXIuIzISugo/tsNfKucgrRkRBh0y7vq
NjpqlobB7N72OTnKV9/KWpxQQ3bFruPr2do6wNkzdrfuyZFC1aUHVAZhmbA5
DfC/dAjUFGoLVGtanyPTqgJ+K+hX2CPpUr1IB1xZCwe2qlIYRZfVwV1lJd8K
FyM+53cTxqvrwXOwWB+/1Y/+DbbiLQREQat2lvyEjlNaGQWrD3B8E6+kalZN
J1qNrWCsUb3J25IBUTJda0teVjuPuKQ+zAKBrAHoXrwqUbCSoOw7O5YrU2Iz
6KkhkZMKQXkfO4camBvaR84YhQjapJagLXFiQMq/b3nboNXC3SLfGpHmpg7+
8QI3kYuoYHWrfSMi5d9DUwDkkur+M1fU+Mv4uoxYqmts6eN6s+ybogAn8WUs
29sGOkxL13zHKzyRTYwcTP4jfIFdO9W89UNhBNSTAkh8QtyWDLTJuWEVDeij
xEpYnpZXMeyp4sr1BHOzsvv0I3mdMjkn8wLvH1VKbaDKpfgEobN8FhjKvsgY
Z5kWK3ZMnlDltT9jHZVTv2K0ABmdmLaVX09Koc9YowbsDO1RXNbiCq7Or73o
XTEHWNLp0Af9y7uKb+MxclcZK97aAuHgxMXbzKG3E4o0nU5Ci5iSdOBjAcEe
4YchwiEKRavfiGLJgfsAsFZTfAFHJ1Lipa/b/IAFEVFjsQ7dGE+uy2qEAtae
BbmN2JoDo758tcceYu5koKEx9ZhezgfIEXIiuQEOOeigD79p3SuC6tFQkrUc
S/RlAiywlIGZOifYLe5w/x5XIzknBBCvRbbCOgD/qhHWJpR4ZdI+U8xoiV16
04EROPfXBX45/IGAkQ167G0oRUUVZUXUR/NpjyBbWcMPRhTvXzU4CNeM1vS0
IBmARYb7eHF4mXM9YAASI9W4py88NHbB7dHJQiaMoE3T3BfsJOGTLtaW0BDc
tVMh/7g7bR2y6HUlETHL4CAYPpwNFMUZWgwox84CoDDyXT0WOJflTIITLrR5
VVjF709Z7gDaMWCB9K84FbF4i7/eYSTMTYxXD2qJjopIKoOvUv3BHwWIxOe6
6XdqA67eamvtZGBqsJfcuwIk0+Q5fC/FwrVATeNN4fbHvYON5dWCAQS5hp1W
R9uAN6H2AI6YNndkJMMQRYQty8TokUqn3Ut9cIP5ZyijIP6oIjmVvU05PUaH
cMqp6YxdybGQ4fI3dCZR5a37pX1PVJ2SwajKiBmoTXAE57Ol38fagvJkaxVr
fVZ1FJ2lF2w/UEgVuXURkIPVZlQhO2BWCrBDWidOqSeAXqNrYqHixGsbiVcM
9QS8DXbzTvq9LLLpBGWERzV+gO1MWz7uNfqhye46CqHTOIeIgZPWmneAd3Vy
GBcCc+Nv6T0fnHgj+FFh3OEAkqr1Xe/VuEBulIyuSAkHSqRVyHkIVByKBmq7
AJeoiKqs2U2C0P4Jv54D3M3c6FQPsp9QYQwBd+t7ftDJ6/5rVZsamTP0JqG1
sti5/3+EnXmFqLvKV9wL2vgCi6DtNkQMwas/1iUZp5JXB3rFv0LV8CtvfpL/
BPUbWQE28cVsHzsPHH9uD1f9ak6LPm38JdONAgUSg5L9MgdQYcKu7HdOTEsh
cDBnUX++Oi+jw+tYTIc+oM16pyF3q1GifI6gNISGOGAEBl083eiTHVEp7Ecz
hvJEunNpvZmMXybnaZ3DQFkCspK9FLSu5V9dVUaaLv93yK9Oi55d+Ur+GO0Q
aIV2xzCye/YSqLC4Px0Iste3DiOGn3OUxQgNngJ6dSJpJPI7uKCu4nCN7J/6
xVJ8OvwwwvP7999Q8yRWgXSkrM1qNp6/7rYUM0GeSceWF5xiuPSX8C90N0O1
y8hsu7OR9XIfMy+SnxbwJxNwrOkkJ9DJ/E/TTVZyF8cSsPur4luRj3Paxw54
+xh6H8tcG4l76BZHcBxFtyC7vrEOPwlwyV66ji7W2wja3sQeDLitlX2Sz7Jt
lsg9s8pMWL0OGGL8YCFWXIbsvEus4vmzYtpKgqqD+jepjySDsLe4LdAmEMxC
t7i2KlODZw99lxM83me1pycdFMKILMJL8AMNyocbNl6kP4dL1syOKpL5nIO+
Y0FHpYZfV62gkHC+UcZd2J2DV/IplegFqL9VQvy0TibwuKLgkz9Duj1JCrzQ
9D3mzYVuVSDyEE4fkUgwSpvXY/DX+5oq19jrFSjgX1hZaGEfxslCEKesMd36
IQaKnOpfgxyYuhwRcJj6TF7er3LBniKBmP2H+GLfeaAhGCZbunPFKx+zFnSp
kufHOpV9MvBakreuBRkHLHEQxq6WGazivX5o+8Dhp+Z+Gbxkgl/Aobjl6fsg
QnwKoSmtpLAFYcRe+PYpWJf6Kj1o81XyYBY/s21rAKzAdejhvgb+QaIM/3mr
tPf8SvxecjDfBR9qy2kX7vSzOcZeFQ5yPYI0p/ahAU9fPaBES61AT+Rj22Ui
zp2ym+Zsvut5RipLL9hiDcni/HeaTi7u+/Qsn2fpDw0KCtP5AEF6sCJju+Ai
A07zMTRrVjVgQAQahl0jVYHpeBzIAFYL/jwo8i5/q4JNdQ1eCwfVdU8c0LV9
aiuA7PCyvmlsJmuAoqFP3I2Q8MOnP7J/Q36TyyGyGPTp8ycVgLaXmp7r6ixN
qxkFnd8zz61+xBiwhcFCOPDJGQASAY6sv69gJONlX2NUSveM6HqGC01b6tkD
4ridUBoHOsK6k44MaU0QyLVVIFm3F/LBUcMNx6t4DpOKEgXzL/34NewdH0YX
YTNvhYQ0QlEOUTPdl2/smYLoFAwM5FeFSZDkmuryunBDpDDiBSGZhobNLYZz
MzjQz/YO0/bDOeRcIzpKM+bYZnQ9DvifJdsWg3HHaaEr7KdLnQp80mWcKS7y
R88dpzvkLvucvrcJyZKAoC6IiJz1Aau2ZkuqSwCXlFvHOOshietjZgBEzCyz
6boRF5Pre0YpuupglU2qmGlKWbEA10fM7Lb9/Wt2p15GlFjooc2linwQHjpn
t/TwDsdA0Jq8sxGklY0NkQCOz6Igv2s6C7jq/p5ZAwM+FL4THsaQiTYZVU4R
jfEnJKaksaViFLR5e6VUQorU9ShRQwtvApjJ3PrqPYqRBxDHHsYvVK6QZbfV
wsd00ftUf5hu5faUNZO3G/PeYeShRQ1eCCJHbzBY5S6+wzjT2idjDSa/M8UB
AbnPV6IgLWj4SuLUW9jlabOYfiL3DDR+yLw32JlPab5rdsJTEekneEtIcZtd
LIxoO+sOCJDWgXzzPTPO1XyFdC+CZ8BNsw/kl1jdiCtoEQtZBRzRG6nkcvT3
nAYwHbViZhIjv8LsnnFm++1rLZsnRsgGn7pzzQk/EAxu3KYXAbKTRCCn8SOs
N/zXNPNoZxuCgmuNG3xmyllBlvg6JhMBEwOoyUnXN7z0IxmjG3psLIdojqaW
41+rHHt5LOaG6cjeY4NY/9wXM1F/5ERIQ9MFyMd2vRXiFl4bikSpe9OaLfXL
TlX02TlzHnNJEzS+ef1Tln4jv5x8GWN7RHRTUgKpFyKgtO4EJL99wuTgqfxA
46IcgpzYneWbck9VolYc+8itpUXoaPdey0zJyMy7KqkU6W3ZIYUbCypgflqy
MAUYPrr0kJYkbn38FBtx2NsXlHOmO9dg01UuqFp+V44WZiMcJw3GBJLdTyYz
kUlW7zctGcFBiFnXNZCiDKGhmOScOd9d/hXM/eOmpkKr0Rhm9d7jLdC6yreq
OSkSS8KKqPyKT9FDc93O4AKhc+3AOirnhX9VooEwLuYx+iDihCcEIYIpgu/9
t7YRdIFwcSxtGz26oCxriXbg9ohV2E1jqMXXvu2dloMCCFa6vMLGng4VVVwE
nJs0iaORRcbhZcUjP1MT/vAPSLvToFisaYJqg4jCpxQ2xb+dRtyeePhR76AD
jecRIuggO24eht44sSHA19gMYu0F1ituqTuB6Z5cBhvxdj217OW9KHcaYnEl
RvQbo6O0VZMoK6h9K+IYppK1dMSgcgkIXo166KKZu0XZtwL+KhEQ92e6mqnU
jd0on0B8avSxFiijGYMpn18yKVA1lRePFiU0AEtOHJLpE6KXzKwqymU88OkC
yY+6wRGZAf89drRO1C5win5Dea8KphgwU6pQv1hqqX+ZWHzpub+nGYw+iKeE
6uhlG8czFQTJipUzkwFZm6zOM/0+PlO1erWCymu+QpBMdj+14IzTek4Wda1U
MwPEWqeGuSta1h43acggCJH3aYJue35zJ3hSexSx7dwBdNSgBgFulROcYJZn
dLMh61rC4FWz3Y1yYNhNYaLMRfJUqHgguI+bz8maj66Q3jife+i+njNs39s+
YEVEeL3mqbKXl1T3a4gfZqPbcURHGIXInYUdi/m4dAU7q5GxEN3VzPTDfcuC
YlDpzE7DdjPrTFGK2AYY9t58wTI6sKQPPJdituKi44JhYIbTRaBaXIPK/zJ0
dmuDefRT3hm0hRu2fQh61m2tjpz4bDnYmGlJhvoA0XAG4ISJr3f44Y6wMuu8
ABRN93wTxBd/gFZ3f/WHj3vVzmt85VmbRxz8S/Kd8bkwtqPP/bs3dzRpZEl8
BeaTvgE2bXiDkYf6UECRHkLHScd/ByfDxlFDzh0R0Ro440K2kYTJ+H5lscnM
wLOch7aviQa672oeXKvTE/unu/XXPLFESo3Iwqqd2osedDuN6KOd2TIqYgVn
zJKuOvyf9ZcBF8/7505R9CWcI0f7mxQFiotwDdrAlzuEc4v0pZG7oT2AqW5c
ZjyI4DpM8Jsnu46jvX+uLKSgy4EXTWjE2S8LPICg4tg6+LWbDREwk4hSx293
EtbhlP6vULzkZyAhSkp9qmiylIQUbOpKiFY8ZAXvoqVapamHII4cY5oMt07c
LI3gmunQuV2+M7GNLeCe7c7VrsEK5XR+LBbrxlpB6gzqnRS4kN84KcY4fIBE
htBFjfinbnVClc4L5+pg3s2QWwvtbpp6HOgyVrHpLXY4hv+h0LyMsAKcv3pS
wGBnFbeqvYKcXAqRXTcr0kuTSjsEgNMQyLvu63eiR11Q/K31x39cvteqoyoh
i8cwyT8xrdH+mLmyHyUhmTicw6nKu9R9l02HCod49DLCue9sd0sYFeRb5H8H
ixGxhyJQPlIMLyTtC6d2vATxF8KOVWAvlzuWEPlemdkW0Jgf0I5eJDjM5xpy
8WqO7c+PBX/STS1wkUeXHgFRNvbZ2nY3KuyUwoS7951GHEqZWsAxnviWAgHm
7BPGdUXakJcssZMUfgQ0ONtIQuyPEAZlqVUSIpRhie/W7V3zt7aXU/Y6npXz
zYl1HSr7f96hCc2pHB5SGraOb6qpV7jZk8byCUjPjZUTiUis4cTk4KgQcjak
MHroSBnBKJ+O8nP0I7XenQKkeCXWoIcHVYogrpQNefAR4f7EHxFkP+x3Ekij
f1geiMLQIGKkiE4TdfTUwQuFOVOkUDk233IdkA7A7a9jQzDMuUzQxCGkpEnN
II53UWVuHyqGRzjI6ozPHIXqYCyzrv+whCel3iBdqxk/46takdJfyqKPVO8C
2fhDgRoutktpURxjF3UKLUUoJ2KE9WEzBATsXB2WxzmP5lwkGo3jnssXfNRr
ps3+p6eB8DKkjPj56fGMKxxtOl0KUndgggicEPFHVLTbD8wP/8h1zyKXsbST
w7+6UPBxT7snobasaerEwMbbAMqRv3bbXAgELBL9gwQsIJhHy2fsXaLXJ0oX
HGSIg8sR9I/ZBllYRzQSOKCyMPrmvWkf71GZG/tXkxAmai9zLXBiT+Sg7pQP
OaZ0d4DyM3Kj2qZ+pBh7R6+n7BA1nw6zTR1oreA+O8OL89KqYA7Ym/E214tg
z1fVjUBLnzPVTnroRNL0NtHAvXASuTkzxWZfkjvzp8Wbh6gvWnm3+r2wrOgV
xHz0ngAi89yOmDxGOAk0gb03nNWey6Ix9zM7hpXI9Jr61uQ6FZhD+Dw4nZtk
bGXOWYdaWnxszL4cUj1KDk/uOvY0s60nyoH1mdcUpnyGkacAkLtw/RgYBKNz
IrM7uLxR6CM2VkNX7TuOaGzgt2kUvK86MmMlagpJ8h6rGw3q3C5u7ywm2lEk
2wF0leY0tcdX6fGfQrtnuPEf2S8P9QzRN8OEVAEycM0dUaFS4nat1/TnMNaH
MTI84FsEJup+lryamLAaqMo5JyE7+OUCCJ4fN/cYmzrehubn+iXB0PhDm4FQ
te4A2tlkscVaoqQ/uv2sJSRzUyhsaE/5rXekpFRZBHHfVStp0BXggcTDI/9p
Hzvow6pGmYh2cYLLv6AWO3NadthHrI4/UhvVuCabdY5/CzBBLOsIWENMgnA1
p+MtvyJ9l2t1EUWy7VWiYAq0r3xdpn46OGZ2crps+weozmZTOQtNLNKElVqX
rH05865VpKix8KttlB0QzKBijY8GHbbY8NRcsZXZFyQj1lBomAyDQiccgqTV
9SKk6G+wvBRbljGJYs1naoUgw1QD47ytNL+XUCQe608eIyLqE9RsFlG1wgjh
lmveaCGYH5EqXALl40xG/9CsRG6ae4X7XGItSKatXLbHspdvta1HDbUc63g6
aD4PtsNVu8RIbxk/dtfoTjxQkdnLELIxnQygiTWKa6O9PX6HP7yDfZk90h0+
qc2jikWytpeYtjo9azlFlDn9cyC/3pfwGexkFQShhAe0+Y/zJjqKn3P4gPCj
3vxbFMMCTrjWO5fqKNcZE3jj5/yUYiiVzDpfONLIDxuGMb+tsBSKg3P0S82D
WYVfO3FSbP3X5OXzCs6K5AYRxG2leKilQk0Wu6FIuCd4eHTYDYLnsQy8g9bn
NB0JmTaQ6axmecTC3bUAjPJgoafoOqwQrP66DnfGHUjaAA2+e+Qvj75kXtun
d0GTkoVHa72xXnwYAClyJftTlrksaJtWgm26V+LqVED7WYo6Xb+dJwFph90x
3zn4FtwCB0ZvT3zPH+Yyjxyh73oUvItlNJ+M6k/oBnEzdmMUDwdQ3ZSmamgh
5b1gQhGRkrtIYQZ1eaGflhr8VA91Q/uXOcj9AwcBlVe/Dsqro6koCqrw4aco
hMgIASMgmjr4fySXodmtKJhEQW5yX1Sbd5WvYLi4GnOvf506dhXEMp1eXp8r
/NvE4DxMeBrGLookMiONM6zueA4MB5TStHV0P/emvXCbszKThAVVo+eUzqhs
bk6BtSnG53megWnIXIGVfuURdHGDNldHk3accO+U9UHZVHwRgwbk9/WNAIkk
Mme0evwjCtBcS/OxLaXtOCZxvyVGxVIA8wcoo4cAFm4YD6jNdTWBRGLdOF29
n3GE9I88ht1lw0ODiXU7+Wo7Siq3CqhFg8a7zVuCjJEa2PoIek1g6vfwzQRg
uJzQ2JBYLYX09b6I/k8KFt73sM+DvBoi59RPMjlPjY1Oozx+d5Wu3LJzptFx
6mErczhpPNik1F+094OuaVWL5biSOOkySiUuAeuk33Lz6ZeQSU8J2fga/ga9
XwvgDRW95GqPSqMks9zE+kuG1To8rp7UFtAIMmF0z8QurfQCZNCoOzoWgfXC
hz8Sw1+Be15+LcJW3R7ioVikivXlhgu2amrwlkEEG4YOxz9miGSdaFdLj06I
311XmjiTf8UNQG2QDZpxWJLrJ7Ars2OLFx4P+JmCSqq88qIaePzAmTrOApIv
qxTeW7tOzfP6ZKr5ENjCcAB1ivGZZZPV7ct6fdguj/GR/z9dzzj6K/5ZHeMV
LuG1fyfhXcOYzdcDq/KoRiCO9plBdGvBzO07j/sbpMOSERPsk8EIXU19VmUk
ki95jVeIO0eZl0MyqaWxT+jhKsrUZQaGMDBbAYxJLJbsAEs61PsKR2WsxJEe
f2iwPNoCNyNrdICapBdYGCsZ/mlzKioby8S7gIPvoGyuZsHwn/qk0yEevL7g
29P1LLSj4FLMRtgVtVDufTLCGEJwg2lyu/d5cuiJMqRwu4OOa8yT202pgQGx
O3QTjbcE+lpGWNXe752G9UneZhfnVnOkDioNk74H9mj4fbtDJcx0lA/G6zd8
QahBGKOAbpx8frYi2fo9Vm6HxIJAz3icY9UNbqdgHKhwkBw92MkzEVtehGJC
hNha9Ff62F6HgkGW6rAuO/uZLxn0Lpe5WO2cwI1ZV581gRtpSq3yzsfh8zrJ
VlR5C7QyFMOQB2gELczry05IY4HKAnQw1k+Si0r9Ps+g5VIb8ny9KX1A2F+M
cEqsf9K7oSWnOr8dl1Tw5MK+8LoJp4g3a3zDUmU9BfxRNhFOdBajS/OSB1xF
48+SwDnO8ZeWbxE3sFS7xDy+xU5EMLC+QYkcDz/ZhUxj3CB0q696btdllVEe
1Vv4L4a1o3LUSuyvtIk694RbvrDZI7vcdsuKW7PD/VJdBjI1vtzfGpKcrVGY
PQ6lM99rF8qwnpUf8oeY2fHJ3OzYkdeg4Gg32cFjL3ZuOpacuWQTBoioabAR
hNT4Y5c5WhShrXGP97fK/jCMocf1euWILnomlcgpJfuaD+vJqs+ncZPd47fs
S6dYvmG6oWZH9dsDW9Bh7+6I4M3SpO3Eoevb13qL8wpyXGAiIMN9QWGYwHFa
ijhR5aWIm+2/JIpqwXaX0YMbORU6q4iexIeykKg6k7NDJpiao055uJqPxA3E
RrGbJiR5Ga/pd0BniLUduOHCMMWwSYbO7Ix8/b/q+QGEP5KAbUnayZj9JGKs
k2pvE36SznHTRrEXGYVlkBZVc7K9Sl58p7UY7/12XADJLJvwm/yo3YuXqK9p
L5B5ZCg3YF9oKw8XzHKj/I4k37aceT9KKB6Sj+F02/uFme0Vta1yixyF3VDP
iqjkGqbaUrkTU+cv0SQpV1PVxeDW4Mhuj3LSstDnxc1sGA13nepkeLQ5AkS1
/3bODMIlCZdqUY4ddht7y1Oc70MngJFgsfB88jWUeJzpmz7/QC4ob1xco7v0
iNywP8J3kWyTvL8x4jjUt2VQ9tGF96vxD2ln+I7gJwNT36mWPtqmak0PXigp
IDBUNcHTMih3edsHYTHTEkPMJAxAnzOPp9OFh42yR9jQmOiSInzrQ1QpmmJ8
vN65CrLJ0nI4uTwqeFVHv0Um8oQ37vQMTTaOTkPxgJWQgVVBaBNhrU/kvLug
tLpuCRW4qGHB8GKY646icD1YhVm2ivJ/yqyTXGuYW3K4C21qVE4iodvyrLG3
fYD1kZPM1vxKsSTlo/VBlLjGwDAjZQrXBaWHslJS9oLqtxVNLX3lEUo/i16+
9WPI3YKgsMdgVv6d3YQQmdl0Oxhr78AfNybuR3/tGY9a709b0b+JdYGotZZ2
qQJN2V0wyB3Iv9FqJMysepnoh94QRhrPqFYfMBuh9jKrShBhdhJRs6q0ssA1
U6nAuuNmo3oR0DASvBQYBm3GsMkMB71K52kZmO4VqAXfMuHRvmkr0P/g2vR5
fhmiY8NxsTne5dHJaCyEmnb5IAeJuk+kmUeHyicHRxdHubZ4/6ylkmG+3FIg
IZ3eeAvf5DzO3xcwvL/hUFtuCNnyrpEEeFaSlil8Osq9TZDcxX2ofxFQGF4d
cafosCncwb5/DS9GcZ8pmyCuvxg1c4C1iek0v4M7U+rNQ1Supz2YnovfQcxm
ImmrgWF72rFMC81LVSNg2PHrDlRByphZ2Wogm7gHh9AK0TpoCEVAE38Bq9bA
UAt0/JuPglD5dvAl2iDrlCns8nwv7iRRzreqno/QpTS8xX4R9XCEKX5TtMwK
z7vD66G8DUiAd3lvTo/AiVE6NPhVqeXZpEHTlORpVr2SdOSBwYOue9czcXJx
DNigXegOvcbXVAxe6gwSDqtyd32/SmRF+XjndMUfycViiLmkNYYiWQhVKjY2
YLNtWxH12Qhc6eudpd78qwVfTA2aYSxfgYfJB02c5d6Pup5smlY7FnsFpRUP
W/lVLjm5BDchrgdCOSUXrgWVM1ZEcQ0fcrZWEngJhqnqm20rODW58x9/pYc6
X1N+NNdKtpkX/BSJvGEtLc0PQrWAhEccswZCHsmb0g+2IgVa1sdBbtgPWO7u
YmBUjcoeLvBh/5L8F12HGQ62rsg7r8hvuVh4JipD/ncffrL9ilNCsq8gYztt
DuWZPpcdVNBMRGxsMnKhh1d2+FF8FRAX+E4uRfalUTTKH5UAXpa7F/IhOFuP
B0lXc6gyIh4jFPCRXK8NE1uY5YN/4n0kBx+xjUxrDtHfeTRsBlKmbsH47LJT
h+LJ2sKxWZbfsv1u8eWIiVbcaykKlPUznta6Z4PosuMYcXvaW9KexHgv/O9y
HgIpgcYFEAIhP3eJJE2P01Mf6qlTt65GmvH6IAOQA0NwiqBgZnL9dvjAF9r2
ihyZoABcxGBM0yYqPbdmYi66W2UrpkTRUVkcNV06TPFEN8jiEW0j5Kxa9hBZ
vxtIb/Fr9mZ34aa6aBarm74i+fnXhzzDLlo4fFZ/m7WAh/I0uSGKQjPZ/02r
UjVA+fWufUpkMCvmVgCGQMZflXtz4/9tY5lMUcm3ytKqOKmtc0hVHCiF7cp7
t6ygv/BCWJJaHnXN+LWX/wdmkPfekHKQb4hJUkZ2cUaiT893NpfwPpFXM5UM
MtZkV7ve+joHW48rUuryBQ8bPekt1VvHdmxsbKnj7wV9C5N5svmSO6vYxDi1
Mzt6LY6oHzkslVAh1HSUhDd0gK1TShsuTvgytW/fHe3nALvYL8Q7grG7vLfx
8irvOzSCm/+7igh6x7ua5Tum+dK/+1BibtHsUIWmNng8y7vupDy8HQErI5Se
Ve+Ybq1JSl4WmoNHtvtQUlj75FbXcw9/DPcdiNc7vBlAMVlQ7+AXAa12r7cS
2C6LuK8HFN4+p+4OJ2dPMP7ri95nShQrKBopRE0bev8hsR0f+eHfbO7cfZFl
gmtpSpyuH7azsGDZXm3JPBY5KuR/5pUzgKvTmiok01+TjqYph2j9zQExliEJ
oKqgFtlCsFRe/DCNY1hcMpxeX9/f6PKki6ejiL7IslkmqiBKomqHqgDAMbO4
pgZKR3iElVuQsHoDugJEBBdOhdIlS802AsZwYyJX6O+tw9QwS6R7VYlYp8lK
TApbaA4JHB79cGUDZS/JxUgmcKi5tet4lRehRgXIxwEV1PRs/9dhskKohN7m
ilFD+AF4hiPth8ShxlP5yUuHl+GI49kwDqgs7dxQrbGPeTV3ugWlyxLkpR+v
E9xhcNDL9WjY+suH5EAwIrXOmPTsb+CM0wf3vZjp9R6meib0BGqAJBZPexJD
3jNL4ZJNWzrKeGB1S/LLiEHZ9QnRrK0anqosYczWWYXy03ZfLeh0PX1ioxjD
wR299RH7tCqQ2EbmcAiP2i1Ja/vlgzN/LcaXRzLNdgWA1hMuUHxkq7iyCGpq
/W0r5XfhM1Mz4BHM38V8gWZ8AbXkA6gSRv0usrnDgBua3ywLOEkRUkodu1xY
pA0KGUCCfzdA3BUc1dTsJgJ1hzJgEMAmuyiA5w6Xir+QFfVZ5eUBIivWwRYa
ZTgXNy2ucAxSX7Zfosi+qIHptR5Soj2+S9+d88xlRDTkAjzj3mXkFUW5VrNl
7IJ4N01VMWW/To/1Me1NckKSwRviuHr9k0snDzCasjAghud9unxr6aveCwpB
1MJIdtybTval9HIoKetugzt0tdl6LjiU3ONwL1YpSsdThUYv28TCA3oEzlaj
6xjBJLykHaXqx2ckRYonRjPGHRLjte3mBMdgMT9UZ/kCyaDQfdNNC2saDnSG
8oR+etizopVC7nQ+YtdbsX+KO1LzuvU5c0eLASDW0QQmj/Aeyaq4XORovQpO
3S7JDLRHeEA1Q6dPHR0HOnxv9tOjumZIo0VFfLCi42fbapHA+A2d0dZs6JJ2
lOUmZzNqKe/LszeX4PevmzeiZjBoLYh7yCadRiYpjxwqEiO80jLEXQElouXL
vIwhqkcDyguD5XCkwBMK8vEs6uW2h71zXe8KsJwLFiuUQKyxToBF3G5lIgn/
SRcJCESVnGq90ZYu9Y6XxPAwJwomDNmZFz9wq/WBlbVapVsx4q5q69x3AbcK
sZy3qyJAxA3SHvylHtJ0jP5l/C8W8+g0pxtizGRtcxEbQw6BcwxnK8o3leM8
AGqaprcLyXm+jspqRZIYiVAMvmRyr/IPAKQayiVXs+0vTbQa+UH4+dO0QHuP
ZyFTe4r4xFjLbxEUa2AE/H8+NfJ7cj3hw359dG/NqV79Vg+A8UzPVkzBdzQF
D7u8wN2cBIjKRuynxJHD2vuBMtBADVw6Syw1t6CbU00gJy7x3Bvw8gJIwgKh
9ixRnwTdZc8SIeus5K1nG+iPtMa/EkHxrEymf/ttjH7Ow+KBgXe8/RguAcq3
koRUuEkLbzG5rh9yI9rSCdrHwoDkINgtHECLrbw7c40UJI1aB/KGu/qEM9Nu
Ie6jwU7kkVFbUpP+z0U09qZA54ou3sh0dxr5bQ0E8RT0sxXvnEViafWZGid0
7WczqKD6UlVvhGQ3O0zeoWw6hEk7jH1XuwcFFoIta1rCCtr+fMIL0OFTLTGf
XnET1IF/PQAFpascH4RNPKr0RaDq+YosaLx6G9A1WZJALhew3ZsjZsYJhUgP
CX0rDTzyL4gZxK8rJMIQRn6C+jQmVg3I7r/g2nz5itAlGLW/mxJgbScTolFq
JjAMYpK5d+D+GbggQXe32tZfFUZjZXmC/TWPM5+qTqXLnIFzI4kZGWfepZ77
m5waDpBqXUjh2OyW1ZEm7IjPhAxBZV2YSmhH8ISk90rwOP9qcyTMxP33dgZc
0Q2/HWqddupDg2TnzSp1Ra+JNDZBDbdLJQkNSGBSxpJ/DmoZ4KU4z58vJPq0
gazJxvDS5JOMFChuzC20gDiVsICpIMo/SZCghukC4Jvoo5xo+9i38o++UW5S
ANQ7fA4F50LHmnJyawerltjmMuX51mk+9z3DSQsaIIS8DGZRvStcXKzptVqP
DCfNE3PcXrSYUmXzwdm3reEnwfe/86I6L7KI+tuiz08Omv4FcL4RUZgOMalz
VjVw2GAUi8e/mNri8U8mk31X00jD8/xRet+cMt14DqB1Av2z4b2g8XSHvZP4
l5ECyOrHu+yIqBhG8C+plQSvJ6p6foeHDVH1pZo/cTi9clKX5JfgsseCVx3t
VJxviDGSPxxew6ydK1WiVnNWDGHrodVTjcIu1o/aXfi4vtVWDXKuuawSRo1A
1RWIY0BHNtut3VSzV73pxAsUrIROor6QH3zGr6BRFgDN1NcGdHQdFdNWXP26
Z4heD1KQQzs3+I3HZ2AbTGJDR5YY1bIYN1TqRGSJq0T8XFl+ZUsbFpW8tUwV
5E9aM/A4TrLOBKWNX53ach8U8Oy2bfbL/IOpD50cSL9jbfVwWd0CujMAojD+
cvoHN6wFOdriTxkvofBy6dwQAeuJsLvR1sp0qw/pJmmkEYp9dkNM9WWcNB84
B3W4fIMhwjvLi5WGxVs5np7TBPD9WYP5nkHKq3U6sraXXA51U8Dc09GsPTjq
5mtQP6IxhgDEA1FBC9rlVV016oebh28nlyuQyajlHYsic9UK/v/ts1I0Fhn2
QtsdBxKkQs0z5E/H6ktYdBg/UKST+ImDgcbfFLj7ogSmLpFV4wYjgJ5tm574
iMfuiFampIS83VnAC/rx/SfXQ9qa3el6c30u2xNU9FC0sEysgZnIg/8gI573
dXhAU9h//F7H0P09o2Zl0yNyhUUQhML1TC5pw7QJg0H/odIx0o5TkbM/jfMe
le9I8QEW5aolv+qfyY7rzSQydXk1l3E0T7C7WSO3BCcQXQxq6BheSLC2S1kO
pGz+IS11nfsyISVVQAZfmzlaSuxiKxzTltwr08DstzE74YSwfpjzqr7Yr2/x
Yg9vd5vg2eh4/MWOWzv82rUjKlwA2InazbXl7NqxOhkeDMMwjKLZUwCZrMjx
tPS2+KmA0tcTTs1xpzCa7qzqeps3hINfvtBjCdYzSB2LCP26y1eQI7ufJqcp
QCc1ukbLNolPlHpOkKBgMBXABR8TmknvXRN6VC6pxfr3xvm18yHda0ShwKwc
xi5uSvdc4EbVIFcX5WQE6NWx0/Fs6K7A48bXQjIk0YMSZfj9GxxUUl2O2Qcc
uO/ZWLrsI/1UPVastA6M0ftQsPq60m5NPW781r5zxZUzUDWVgx/oLBRGsAu5
rNOpH0p4MxVHmtvy6Zi1MlkbrlxYw3GKRDcvXL/mfcFQhoiJzzNo2zRVZtlK
IXaGgf1clByzJfTHUnnVJYVi8MvT8bu2NdvUfIqngMO3l9NY2WGI4MLMR8eU
Vilbrh8i5fX0mm4L5ZjgXKl6MC5esq3zQj/mWblKxcq6MdiuwsL+9V2dZYau
tSoMIut/LHTGGsDGx5jj6OAGjsSqxdiMoerttokaPGquCP7RYjvp4aEoseg7
bEpmHphwnFuhzft06q9pxxh0jvJe09c8UdJGohcpeFc91Gb+p30X3bA4o79/
VfTjxtZ9AKhC9ZHYftAr4O3fNQL8PGGJiCTp9OjxIPgFoZF5oLWa8K+XA5xH
iaqTnevA1nTqd8Sh0c5g7/tavKZvrbuE5Q0T3Nsk4Ksx2lr9CxSkTmor4ymV
FaVumRod8+Dhw2neJd4/Ck4Ig0T6iRkVGjiSV+HynsM/jQFxQuxWs21H8A5O
Y/LcM/bP8Em7PFzEaVwA77sBttw4R8chbUuOyDrfz5fMbA8k6eig6Ow40HOp
W7oTrVdbAfcaDuse4+Jp5JeFdwbsX7tObwt0B3PELZhF4ePKEgk9xXg2Nnuw
Bq9jfycMnWDsu7pa4+Z42NSsxgj4onbilx5i6A5HL/8Rjq59RXIGoCbG7Wz8
w7cYyyLdiuDpoV7466b46I2/lzjhuQ/JQAf/dvXYZ6InovnlMBZ3jEfLZdei
R4yDPLsPStlNKAwTaMg94fUwLCzbBBbmlE6MH9dJ2dbb7LLsuG+tCMLq6gmD
oRUDfXjW+qTE5ixhsVfij2K01+2uqFY9YliRxctpjsnhiXbcpITMSYCglFOd
qZNZJ7xZtdeoIletkFxFUIH7F7y7drl+rr8ejKPMtmf8Yiay3Zjls1h4M9K4
S4KLRGATkTdDe2S4bWxVyhd68fS2t/xGVoqJjulCGmv4wq3fdvm4+9isOEep
s3zvBPRLkMiaprGnN1uxDTnLZdL/0vyH4MFv0OiKXtw18HT6+nVxGwKGn/th
gR7A2IgDdjheTX2R3ll0mhJgoWuC8OinMd/P90UGlKxRhGwDJ+IKJor8pZD/
KzYdT3xvnXdrU9Qj/5CVR4PqJUNhojHW6uWsmBcWPz6xMyiH/aKu+S8qMZwG
llPK0Jib1Zcy/foK/eamrkd87DdXUC15Kh5+v7YIiRpqG1E07FKZ6JAeH2Cp
AnNlvs9eiHzyugI6/BOrzDQKZvLSEh0YvoT3LrmX5vPD5D4kHyhrNcnLGRyq
68nDEMHcMNuIwWtbqCftDYBKYOxSKJaqm5hwJiY+87jikwieRJIGwOnhONw2
wP9jWp/ipJGoUIydLg9MusuzUvu+6Tp68V6HeYr+63XUYW7jpYixoqDGWrL2
6ObLu2iquFmRGVgJ7dNAnaqRcWypK4w3IwSE0FdxgGJ1gRAhetFE7G+hyHut
HOAic4HeYHiKVZYji4eI9MowE7XBmsxUo993YhsS1z4ZWNADazTFSOga0B3I
LDQ/jN9SN434qfhu5OtBgzcP16MKnRlDa9TRs1c2GS+ioKAlxu0XJRx4cBUs
OVoGkVJYk69YqYpKdZ16yz+Ko6rTHjdZVR8tfOPGQeODvMy6BG2OPUgWZLQM
kxUY9G20ryBbjw4aP8MZ+AhQmtAy8PnDyzqv4sBela9oQ7js+HyPjnPFXG/6
/kz3nzqESoQJ2KYuF9c6GjkUIXte/cgzIqSDLIeXVn5Wxz0Tc50wOK32cTQU
j2xnWECYMNHBChE6Eza7/t7O/VhpgN/95UdbaN9wE+KY4EsoKac1e2QyaXD7
9JiA2caEXdn/MvaeU6IfMjdqDZjHagP7oBgFyt6+/IiY3wk4oukngLEhSAd2
SACKUTkLrVuOpQ+sMPnSqWFS+8dfqpeT2HJsUztOcgDBUDjWX6EqUCgjWdCb
ATOIg8EpHhuCRICi+IHbkSG74uFt8K5N9huLBQIwB+ubOcxTVCbHxUPVxiXU
+Pb1jmZ8XqYFu/Y1jKH5Ymt9H2K2CtAjVnXou66AaGdfZFOTtGiqzLRk5SXY
cMVogerm87ZK3iMyO+TG43bTtooSiC7kUZsmS9elobVphKIpeXiMk/HSH9pC
3n8zvcZS/BPLI3/eGqHiysL0iMlI2fLekuzMClXfL8bkZAwxtuH300BWDesZ
Oqi5NIvuFPUKQ4bG1f17JofCDC/bnCQXqPLytvfJ5MfHf+giKaItEqpuYaUD
S9j+zlSmzggPSAUZ9oyG4B9EWBu/ZWx2QLwR4LFfyMJCJiHRyTgVOES9e9i6
hmRL31wWCZz7D0cfmzqGHez64X3rJmMNA437rBiiME70eLjva5RbSnrHz6ht
dfnVRCB03pGCq8dOS4vqN5lSJxUlJd/6P0vT3/CBwURcw7Bteu2rtFQzpWug
FmfY04YThp1gYXblDaqzoEqy1/R651MYC1w2IKnrhiCWSZslDqUuhzjaaoXy
MXwXvpUpMT4yFP/Ih3etSjJKGN2El+3rs+xMZ0ZrByGsJ8hw8ibqv/NT/vx7
RwoyQRbmn0Ml5rVn9GSOUXfIjyWdW6yUNxc7NiHP5I2G6GxajH++9c6Xf8d6
pKHCKnCIMQqZxAYu1fklSfDL+OCk/6OGi8GBs0Rqcp1qcIen+1jflGSFUvPF
D1F6mqn8srkdbfUNd3uC/9SjQKzl9wLWqaOq4bGg31OqecVt1BNnuoNgquDM
9qxatUVnlsgSD4uSvXKtUx7QNEQL0vS3FyLXDjJuFGimZXVeG2tL6y5b8yEd
gbBLUgpeW9j5g39962sICOlG08SUJjQuj+J3GDrH+5BU9mRjVY5GbCGJyPEq
j8IHfVjqwYSxhVL1bZfS4jT9xgVTKz6IIOB5Qu/5w4qdvrxCPcGcE+gCSSnp
O2np9pChkY9qLIPJ0pjVHZO/fMI5i1ftV70A/LZanzwgnUZ1hUaNwVARxSZi
5N6GNS75ELQUCFOeipd+ctjHEVwsQfue8CNLq89LLByRN6oVpY8NzDPkNBxa
SShiC+5VQiM6UzKOTjgopbzS2MczHSB2KET0zlnlSSYacxzhIpO2QmAP0Epn
bITEPxgkm07V1+eus1XsqQugmeasqaDmJ5tgPLJPODm+U5FQjzjnj03iPnTU
qxVZFlkxgO75S3xatsFb/In4ovIyHJA9Cu2MisXbLUvBSVjkKCkK0XXN9bVN
6QoeyJw36+EwMtU9rKQ6Cvjvc+Q32/3YiACyt+hO8K6Zbk6c5tnghkfvRYsa
oCmx/+a8V+QeYsEVXt3pnqCMQQsGGlGWf/Wno7LN9hHmcsctM7w6p2KIC6Ao
CYgI1Xq5gcGUE/qOdICYIbGQphwVDnXolZEtTa6Cl2AOp07ypJ4IdxvVQOgQ
Z8pVZlBqlv8uE3/c5DqWOxCyB2znGg/LETaBFd68mbdZhliFb6BnUZWK0Y/j
eftK08iBQ3Sd2Q9lB7PABL37qt3+FoiIrqimdbX/gPDc+iNDA8N9EozyK2S2
7lEzGrnOKrFG5eaiq0Xw0zJO37Q2sgE+BlgeGGvJSryfOocs14PimMCDELBd
9aflAw5Nhk/YEyV+riYd7zkYIoIXqkS4Z49+buBsJgMS4drDbJSsRD8wetgR
YB/VYrJllBA4wzgGhmBreehNQS8j2eehNTK84vB9EizKUI1P5TFs1nqeLuIx
DDn38/JXQaUtYYKNolfwWv/6GKlOBWnYBFIOqxZCLJKIJq9wJL+IG9NEIzsY
ZGNkmNgX8nxl8OlsEGqJWblBl5qdy6JWqRlTx2xWmVuWy1mu/gNGoj5TyoG5
rmUpfxCBH4BztL2MMXqLiLJ6qVWRslVQE56lYo3fPOVDp6dazatPAwB3e4E6
oNkBnxIzLJ6wvPC1OHSwrL6s0tMs+cqipROBBVvBxcYXPRQIKiS6heZ7Rm8G
jkAraB25sre8pQ/EzHFmaHLgJ8A3rcJF3LfqoJzLkTu8pNPoTLpbCEfIXb/S
tJ/JsU0IR34ht8wtW990h+w8IKt9dAIY1wy2E9t/n70zHGX2CMB4oWW0ZiUT
WD+QIcsop608ui+WsJOlb2CJDIp5noaNboV3iak+14InxLXT5GDcSRsk2JId
ihvzaNjUnD4b5aksEUDDWy2QJjgWb1CvgweS8jtgE+P5vWuL0mRD7+Z6MUW4
xJKKxT+lIuZoQ9fkV9km0/jmQE0UzJWLNT8ZV1czuEGYJXxmIIPJ+K61uvKA
nv9EYAXe7Zt9CpwuzUf9XqmlBfPpEyFUZ3Un14w/BpWYApHUm+B0Of8EbKbw
hgaC+rih71U9nW2DdGgsl7Hb5xmHnQZqwyHCkETVeLISg6R2Iyh65TXd3xs4
M7rI2c/alcnxhcyZ4CQ8EB2TvCSsdCRrly9xEmkWxm12zl+xVkZGTFo/RdWQ
FnWoCK3hH456QLXbvCuRfCkdUBJ0WKEoVmqaJ4hRnTua/PR55eQsk6NoYV9E
qbE073ggVlXwVp4vKFiFMuO8t3fgd+bxKW+xjPzyU96Txl1SblDBQIqSfhCI
2WcNV2i/tped9JfEwwe5LHAHup1rRc/B8HebZn3tegWStND53rKPrLp8UMY6
EG/iraBF8pfrNWXZNEYWiok8Bc6ySdwypSS0j6AiROFKHqQQn4+A3rEAZe7P
GZZh0PPka2k8qAUPW6q9kzmr8eTFdlvc4AH/586QLB70PbakWfA50bFp1SB1
KBq3uuanGLbN93BtpWH5ldwmFG1GxxO6Ngeo7Vams2oAgV6K+LbDjcp4HU3/
o1kl02Tm/A0fWZ1NCgQ+PkFBZn5x4V9uJPnQ0UrDvDAOIz62tunYWNg6KQsB
p/jvvr5iZFIpC4iMinhgNEBerpZ3EdALrnWGPK9fNhVLR5cAljmpl8ZzkckQ
fHj8rTfNEJb/AlBJAsAoySywgguam8lQzFjAMNoZqiXHugSkIOUSqnS+kM+x
dv59dLNsBrWHMlB3eFkq9X8N/okiJyymibWAQnpDuWpeuQ2rTRYoUy7TI1Xb
5Cuw8l/qaWB3xNnoBjPAtFMRHdv/A/cbcCSLbN59lBPXknzOo6qFu389BsR9
FcwnC2l546zRZEZAPt9vZ/ExYhCVDR3OKDl7JtJWWWeD73bUWwlrVUN6ngl9
0+NiqTMyJN5V0SPQEW1eLihIzl6Ah+2USNlm4lDOPSBCuxuHaiXPc+apdmdI
07vqtM3UCNGx2+PrATUkBBu6AnrfbmraR4kzdtF508mHsxQ3dJNrJqsUNbz7
wvPhDrRGjKS9SCmULIMeJ5F7dHJ2abVyl72OCH1TmYags4Aooz+UhDQihGdU
tr5204Zd/EU5+5GHQHzYW41y/dIufE8zq6u2SXjQqOnSi9LDfk4P58NGVtC4
cXgF4eVzA57Oq8fIiUGgP/pVHnSex1FDZemxtabadl7iXub65ECdz9c1OSj4
MzhxsQZriDSVmbey0usuM/izfhEWagEgLtWqdkBrsAuR8NUoq4eyP3PeDZa8
3BtUSS3oth5ZL6aO0tVZjVcnLGuYED76QU3lCN7yRWGw4BJUdyN9nhaZnPg0
tQypR1fSoRCRoSjSNmbrNms6OpIgbD/hXps2IUm2Rbr5saUIwOpoiiArbs1A
rNxt6GMydUFDyAiuuRhkfMMQA/gB0bPliUwUHyq7r6RvBy7Eksbr8w1jVliz
/fZSe6AZ3hK1HjqHMh5dmRAdrQLesLyTqA9rzL3WASMFObtdrs7XP9YluAcz
EMD7iMxX1BWi4DzBxtKqId0L7V8S4LpnwUzbt48tO3NOIIJfK/D/JQq7DQDc
eesi3MH6sGZ6M0pwaGklFyi9FLhFGgQFIq+zG3v10RgOBfLX1Rv/a6FNpSJO
UjqOmoHubWn9rnMSM0nBYYtWmxpts16/Z7RuyjhRESIgKY/BEcrAzGJ3gpUn
nEyqCEnMVLZ3KYMnBOtdcN4xTZ7hmzoFIaZcqgRZpv5Zm1p9xfe15eBRVbrD
NGUm/LvlV/imzNeJL5N8EsuCj1IzbKAOi5jMByDZ0wQJpz7u18pNWTQr8FEZ
VU/vMyTpeTf4O4ETN80Vu9qBxkcgRBuK+8bsq5h/nzUaO+bNjodHXFkY2HwV
UTNdBLtJrseheLMtFWSss3tf4/IJ3AJ+3fpv0rUbCQgioUiq0uXVYDBk3/49
iz4rfsrp9XNuQpfwTIQy6STxoP0Z96QXlDUm1ipccb40vvrlLZ/cwNmYnbE6
Wua7C7AXAoou7MKTc0jOfKgf2WDIKazb/vKgD910z0fkeZ/O30E9qEJMAlUg
X6eNYJaJC6b0mXP0/OMUuW/WTDBXySmarWfbhfNtT8oIXm7ot86AS5+pJo0E
sabaQyNNjt8Ccs/ak5V0vFW5FxzMclXrIY058ZK9mZPudGyk4nG/9vnhXUnC
CO13n0s7SS+OAN648/gTPy83Fb6OXjhxDCMN5Mm8Hmz4bO4/gFJHOt8eQzt0
sEGNwwkh47mecSPclIoUb8/s9t2KvSWo/lsRyM0vZSRRcV5jrdc4bCuo85wu
6iUFTMoVMPXIiti9uw58pndtWXf1j5zjRYkrHNKwy/zd2W+8P0VMA6sC3MsN
6DtZRBe2mYmRVeobpDpwt/8gUfUS2a9+ouGBrU62+ze8xkIiEhGWJWV19Y84
Vk7TJbdNNAsk6C5YkldVkwW3uCQgkOclIXYaYLG1ns1t4G4yNFwn7Xfx5PHq
QVM6Yx1YhPqimy9TnOvXCvgxk7OSwbG/pFF1Kv3qfYV+8fo8NZeq+z9BlfIB
HLaVHThGHNPl8W5o/AATaXgg61d7jP8D5Pz/UeVAdugaXfwpd42vsRxJm7o3
dft9tQ7ndPYb91osAy83hEHYXIPXXB2LMOE0Mh/oTFfBSr/mtB0O6/kBQPxI
P/HbA99K6Ry2xZuG8QpWKFotmFfTDiNxqQWZi9dbJOUKCTfvdFzEfxK2OfAI
8qn8lzSsT0tMy5XdRLeHpvIjGEmXFAv6v1DxrDx0Sgho0zFQF8bWVanHHXE8
avWHobEwYcgEwO8T/XQIGQtrnWLkzk041/WTUsoRm4/Yw51KaVoSzZgk/TW+
bQCKaQz0NRENZIU01xETUMgBUj3591IQ8j+85o9qNOwxqSLIZBmxa8jGfy/l
niSrwyitMD14A/OBMwSfxnsLeVcz5Z0/J5AeFba4xZPgiijHPk485DLgx9Jc
nwvFjF0X6aLfBYdJ06N8bdV9ZLbANgV2b+uW1on++uEx00uzTR3+lRYhSGKw
sRiGBb1l7a+/9mwLmLoeBaryb2K0XDkNdWTh1+xHCgGQZayxFtbselUMTl2N
PpopnV+xrnwhnOkcJnjumli1T1Q/sN19hC+hBrCWTxDvIM9zns2K4R0qx1xU
OWiBM8U+WscYnxU1aw7syxKFqIxUwmwKfF7g+4ilahFVHIuemljidFdvTltV
GviumpZOsv9B3jwQF8zAEk2pLsPdCcGv8ZMKZwjCUoUp0P02phSEVCh6Sbs1
KI1wV5sg0dG7IBapKcGWWqcav5wMTLRlRgUGxP4d/xaJTEc9vyBk8K8RwyAE
n+lMYcrk3yvmak64LlUaQ63W+tNnObxSk/5oOMBg4awo6AGROgQvQEnSBCdW
6wHzm3S1ufNVeMNzqbO5PLF9VO9oHb8zV37QBEI/GMRZzXoFg/1kEc8CR67n
hBAXuT8Txi6IsDDEt8o1karxtxYwnch/qJm1dauYP9ZfiXt/B2Egk0uuea0E
hSs1oNFkFjJyjw1J0baeT2Z6JpEuOvdGe5BhQKwvg9Fd+ANkzh4EGdMQ4hxc
pKsNkzcM4StDYlh8OZxiDxBsix09QIzBxk598cheTS+wG9UNST28GIurNY8R
dqIlYQMAeY5Vd0Vk3xmE8Zxs9TRn+xcNRjKs/L4NjvmoAuJGo11vny3e8ONu
DWiJYFi+nf25BruYITIf2v4TTZpw06KeA4JZQPqfHioWrOOvG7fWdlJIvfy7
xkZEiRn+fTcka2zGWO25B+4rhIpj+2kAaoi77zgnRj7ORyEDI7XrOnefeijI
rR6Zae6PfGZi1hgyKiz9oJHVeg2mk6MuCINhr9nN//Eb5hHo3I771XWR0Oc4
2+9/OC7F1bB9A6vOtToBAdDoqvC65Uy3n0jKwXso02imQHSWSN1TpT/6q5LX
qi3ZxBB5RhdJuZahD/c3vuWRszvjlBLpw9x0mS6fhv8vNpQH7wnWQZDc6l7y
DeZTYwe/s2YSjzVZP84G3EuxMTbFSTMT62IPOjxnW7NaHVJSBBB+8xLnJXq9
J+f4rcsZjd5hbxao1LLfv3iKPjdP9GK2hSsA0yMwP3EkUYX1e08rh+v2wdH8
pcs7AJf7ts6nOWKiHoToW637E3hcrdFC9GEbrjBModfbXScHLstSyf4jedFm
AQXHhtoBHRxHq7tT74ET/zVY7o+hJeuAS3MVgg3LFON9PHxqQvLirFfQ78cP
G6CmzsE9JcqDXXzYw8tgNlhudpnImTBKCc6567p/S9JXcMpO9TLoQRYr1L+h
fEXzOsfB2QVSg7s/hhfKNu906KcqmAB2M9y8DsJv8HWQhArLyO9t3bAPvX//
/WlB9fXukirKV3vRsBj4Xr/f0AvRfcIYzB+F2yd6609uJQt4j/rvitiBZsy8
SYTHSyd7EbRUKYBkBZeZFk9pcbMa2xzntvNEDxARDkVfFFxTxAzZsbE4+PWs
/WqdTZJAqCeFrUdkM0+yUSD8q4hFVWaFcGHjJhwwNUqWJTjPc9RQWpAcfTiW
1cjglzgkkAOF+fNT3GGEgmgZws2wF8MVvb1oyn9H9TrvlHtDNOxVvdEfRSaQ
04H7AfyJicHEYWC3zTw2IWhYYzbJV1mIJclpzQ89I117sVB2c2Qli9+cU/Uz
K2BgConrtKucpS+j7wUycETvO0LZcZlhlShrGeAiaBayVSGa77emmDD5w5tZ
MUm8wHwxPGapelsu+mI8RN7wHgVNep6mqnsCgBcn9O9aZZpw052jqu2bIYIL
tfO2ZucID4GJDTREAUKVEJbVDd39AYItJaGWeCOfP64kguDcC04Pd8nlGjL3
K0A9CCGmD5IGEQSIgwCRNkeHJKVAHsV8gLCJGBJskZfPxFDj70sOM+T6G05W
xL7y8QXhzWjdj9vYH2JcxxaM6lkXOXa8w7cssWyZG/EVHHkxFzmGfOFtO9KE
V9gGd8akA4BONZju2owfHTvbkDzR9opBh2wVKQwRD652/wyRbVWF2vyg8uiL
VLL55nQcPYQ6gMNsb2eaNA8AMQXnK3BKgBdSWDZu7dmPrbAavybckx2/vTlQ
7veuwRcjDvGfhE1EU/qtI7Rl+NXkExnXAD2Hi+mV1j70h5JLDaM2MaDuNw9z
2SHoLj+u8hq6EbrgGsDYc2bAmskEhQrypKlAMLTFylwoaSkUjyyKd/mDjnt9
6e/9rdHfV8oH0pQIBaWSQ/hTS1b4V0b0Nd+CzxeXPqChjBo4p9lclhSk+tcj
UEhlUMaCPlCEz7ors3lMrAAWFwcjV0cYtm1AE1BDzaoph5Idv32dvhD7ubdF
Q/gZH1RauWHmle2CVFcMfdJ7uwUywHOvFS5VW/CEKkAmFH0qcqVs+4HtDTgG
yP60vhoD8IwyapJtq6iy0RKFTrPzBVGzSZThz7rFsDkVNe2iYPFHlw6eW23V
L/VXxt3i1RI7UEmxZxfQF/cgiu87ROJw2IwmLLfQN6iij55784xeA2HJmQzD
D4byEnLlpZKdRAwDzSyFL031FyRG9R7X86aAD/ss5mZTyhNnq+j9wH5cRppt
7t3dkObQ2KsWtAcvxq24N9bb6rcE9z/DMDxPcAGb5CwOkHeoc+TZvmXoqXEk
nu4yCIJt8f9bGSnfHX93YLeK/+Bk7SgdiPd1Z6UJaxxQgYiOyRpemM5nYfQm
8viW//yDm60nbQ32eLwVPYA4CQCSebINi6la7Tm8hbKunRFLDOgyR/fTYwLh
m//wSMTYCX5PUzbT1RqUhODeOfZCbBEdWTEs8qvuJBHloZd8KL358H9w6gBu
QswLMphIipU9znZKs5lnzqzuleUAkeEtwdv/eohYX31/ntBiNiZOzUVdAKnq
NtPN7udQsu3T945+h+MsTPUfDPWKP33t4QEERMQC0CFcV2mGs4dYA8mjefdU
Ej8KkmgqWZ7tp0G0ens1Ms2bUtBfE+DBd/z7dcBW5b1k+ceTllF6nERw6Zrt
2fdJoHmBDiJ6GMl8L+X1oEbwIeM+EiG4XQVzQ32XH9rRLSZOhwxf1pUPc6XY
cw/v6sSm9vbIY9usmjGdgCzhx4VovZsLr8qkDeerFBv+HbqvQBT+JZt9bFBE
VMsP3wMRONQO+FRCRThHMAm66jyT9RihiwmSdQtgyFgDuIgbI3slWcs/AcwP
NxW5KNrAUNtd1PbBVQjy2LwPKESnlHDbFN724dyvT6HSCSHH2COZ9avT1+jG
EAUH83FxfBF3UPyOfDYmY37rH5tsOan0aEIqZN1YAWK5B8dMrDFTPpgoctEP
t8luyYvYLtj5xIMDdH6hGNnWliwWw4bTS1QO344E/1bO8GC/nQkiCO7j3A5K
Kh7mBOp9I/31yEPjTVRCMW5C/2IC9Bs0MZrpWQRNNsXQ7HTD5kugBQGlzfoN
omZpCHpix6SpxqaH2AoTyQ0XxE2H+phBmdsp+NJhYLQHK0SI5xsTzVjuDYQC
tpQl4mvOD1oyaTNmFWtrb66tNTKRg+qVr9tKTkepdyqarACVVWxRmJOEJPA6
6fU2G+EGSQY223W6uO8RREl8RovhvnP58Xkjj5UeQpZkctKWJsLD1yY63Cor
DY0yygfKOdu8Q3ARHOvG6ZhOgRZ/GCu7xABbfRYJV4Hbl1OXqW0NeWRo2mMG
L01m0/7diXjkEf0evbS0CVGiunAoEP6cPpec4SkWV+oLzAWJOT/flp5Zr40j
eZfXZqyxUkFMjPdpUzpGvIv03B7PhZQGW84sCTpqS6wcA2AhIClAlNFGsxlD
OADgIEnG+v/lH0AzrmTcznSRhMKz8Ghdxd7W6WfjRpMETPtxt2qyFMW27aoj
qd1NzdADvC6mmsgskwu66AwramtkcCLc074/gkb9HWj3KqRPPbFwITCnN/ql
2e+lIpKNdQFVeBFCSG5DogvX3yv/zGfwz0AWohClPlkTIYSkwF+omzyd+j+w
1d9jF8wDWsOR6xYn3yrD3XW4+a4jGno9V3PIT6MniyBWIFq7HX9b95sAKsbl
ZO//Rv2XCcZs26Wo3SR+2ppxFR4T+cGL6YUb/blWzHQXryf444cCJIie6cTU
Mn1YVaTVE98Llbrx4wdqiX0suWI9CKDKoMdygJ0g2jJGjMBw8Jd3lZBF+nKC
aztP97EhDb/SlaI1jLxLw1yJraWIAu/t2TNzM183rnwSfg/brdYucxA54gHS
q+ImpzAT95UesHDokTnsHHxTtf5yHgpDd/2/tpsTFe99Qu4BkTVKcBjC0BC6
ZwQz2nmkfZo2EF7gtonOceKE/BJstiL8DGRQN2P8d3d59vUpYkMVePw6cdBR
PJdmZWxo38HsdmgpjrtlCJ2tnNmh4JpsqlC559IMvZqCDrwyNUwBhvjhNzR2
7ToaClBVEQyfahMYal4YlI0wiYwAVv0uYHHSnvjks55C5Cv9hqk8TGHQCG5x
zIfan5UXPyBQA8IMjePktCw5jMlqwCCDx7s2c9kjsvdfLdUiI5gtHiFSVtOC
pk6eu5Zgd17H3rZht7UycSSeaAxC2635SBtJdeFTrOYv+Z6ZbYZaGobVLzu6
e9I758UAg9WkrZZlrkD/zLw/mMF+uX5e3N49Ir/NpmJ4bh0hY96m89LurAyJ
PGG+xRkrbU+/UZy5O9X361Ic68k5erDjMVBgp1K/OvZX2oIAM9B0HdshIkn0
s81hD9NiWX+J+hrSYV2LS7ZEPKtLNWwQVW+gRzzGat/3MSPU3YlODDfEnTMi
JfttXO7LhZlIReVGwyYUjOSFOn7LU1ILEXgMCudhC0+62psy2iKsJ6hxZTIW
2eflIvaA082A9Zb5TUcloKAwSrpPHUZHRByNW7ODFHO5OGd5tGNPVuqtPKeO
Q/riASNE8iMhqWX0HPY9FqGfQjZGEfyfXYa+9clR3bvfpxm88C24XiEJ8anA
duiTLWZ7K1l5bEM3T4y+B1dwDlVuuNYxVfhylsWs5dqGhki2Nr4ukZjCC0Sd
v1DdjWIR3wCzmoMielKjyDA+4PGrQnLwhqqZdxmzwpCgbPJLW9O3NRBmreof
WUDnX8g+jN7vny6msm9BtGVNrKWmOCMhrsMefXk2Zz1rlfvqNJCRlIwsscm2
1vQLFdkFvjwF/p+tzXL9Z7kDr9Rymo3KtN5uhdHa89UAp2pC7sKPvidTvmsq
mgqwdSw/nf/oiPhtcOznvtN1GuoslKhHU932Kz3wzHWuCMGz8Mgo8bM80F5e
wPxcow5jRBnQCaAzjhzE5CQsSyAP26zHtwImxrnbcDFaxsSDb22Q1ceKUGfE
8Qj2XAqr3ntvzAVpnmrUPeOAkvdYOnoKKOotGxrcOnV/flrG8fxx5zqMrLoJ
IMieEFraB1l9NBbTVRGzX+s9XV/WfGUn3eCUCkljvLQgtolIq000FDaPPRtf
e/0b2O7JKIjN6jr6xVbveVWVMOk5lquczwxsGvxGT28lIk17QB3m6DHBdoK/
pN2CiObW1hvjKBEkPnDzUxooVSH7vAvnC/lNpE/sKlg1TYvG+Jx4EQI47PPY
Me2B6dmzmizZw3P1dYQq7Y6OQn63cMVScN4enyEZ23mN+x9cQq1n7YVElA/w
xCdM2rdMq+jas5HkWrcJa+wbsulXLj22WB5Ew1QZnMGmiAJSm2aXy9epRPgE
DLY4qCJRC7S6RgidwTTKp3GlW2HdwbYS3k6kIObfFtzhBx8LNXqcC3jYnE6D
CDOkh3L3v6Bn6Mm+VRegUNFSXdKPdVDcwiCZLBg/CsasDM32MPOuS7Frzbhn
Qje5Q6dzdgdoy4dIEeYFW3AbQrch1m3fqi7xyeUf6kyuX0hEFvepbts0nSTi
/l7AT4NuiE3cdrdGgFTy71hicb6NUdJboSRECzX9VrlRlPPN+he9EXARbsGn
yl6yr5jaPWAoGoTqHk+LwwqpavekwC2OVw+YyOSp0TA2brPEFfV8h0+2xDIN
5/Gxo3To6GN0kKfcZs8+sGtpXQ0oZg+w8EgNue0NsL7pzl2GlmK4wPJOCrC+
Ry4DGMu3gPxbKSXQQjSe8eWMydqMwmDtUxkqj1guvQf7ZVN6mo1tE56esCno
k0m/GQgu5ECXypcpR3+h1cmwutxQqKz1/FNZ92wafN7m0apExgkn+eNQFOQM
BIyG1RF0N+Xxh/jxyzHIPYHv8zLs/hZIZLFlcikzz+v3mUnUSwYZymCOiE4r
nnI8ZCKZlKwsQtEd2DXVrwt2s7zr7TWLrOAwTNs0tGo1deQ0Dj62WpjSn7a4
DQd9FaCKqYKNCN/0x9IZUEzyd+OerlMEvzTFQVjpNskL3emepYEnT7YlLTU7
i0116+0BkCVRTtG4RzX8/NKRUre2l9Y6XxyrLZUWaGx1PGa9rb0Pm+nTZqeU
wU/nzDlur1bKzPsLl/ZybfcxzzgZ9yL1N2eV7ijbMfBJKpQbguKJbtwY7mZX
mvAAAhpF9xoSCPDy1V+F2P2YxHTozC5uIKMV5+3Bqxzuih8N2DZrl3XEYFSB
vZ2j8OzxmFEFyvEtlPGqwtK+6bK+utwKXEDem6UF8FDxObQSGDtF9uIiAIC/
NjtVmPH5GMMADYfaQPsFtNi1+DhccszCRzTSTh+DbyEAZRy68I2LOal8K731
oozxDwEnkRwHmVHJFArvtf0n1+YXEqWUu0tWgY0KFuOAS5kHFZoilWKHxJNW
VfV2eZoDxh0YscvEG3hu8Y2N2oQ4o05S63usXdMbRbmbG6esBqt+RKbzdhgj
csqtNdnVn733yHb1Oo6ZngqMy2w2RV5c8+zKtyafzMsLM+l1adEDCut5GM0n
60Toe2ErCBoRrOkGVjhR0LvvNEg2ILulXx16RhUr4MGnfUFSklPkNcdXD3K1
w14eEKu+L8aJGreGZ/tfyjKHchZIFRe+gPomgapeqpDEzbQr0qAMLqIpeMl7
jiKMvk1OQO8CeheAuA3WqcSZGGCYLU3gGXOjIA6uyVGpnKdsf59icK3SCfHA
vXjYuWhYeR/2Lyd7OgOuc21YqT8qrzqyP+guUbghrVBWEbdj175lZECrwGnU
eh3Y+Q/OFim0a+Q2NhHEdvIyrzu17hD5sojipBWRGEZuo0v5ujn+79NAoXkD
VB1S+u3Dee7OhSqVqg1hnIHfLAJ+A/3oWdS4YU4FUhnPJB5yL7NqiQQYpnfV
9LWQy8cHNwHsxqF0Ddp6fMhWm1IC1hOdCEYwQoqRlb/+sxaiw+VHlyBvc3BO
gM1HTjUY26y9YPD1/a5rBcMl7L1eEvWcsFKPHihGKak/jSwTOSa8/vAsoMZa
PQP+Mj+pwzg6bdqYGERAuEEY2RBQJnH34Y69huBkSDiQ2XPBInnTyK+VtAX5
L0tac2JfI6eUTPHQKGooWhnin+qzrRKWWYMxsRf7QP+9q/gn3BKR3bBcfw0L
/1UdXrYGZd240fTo559IrWFWFVL1NFb7h5GanByZW0CXrZs4InBcnQFkEUKZ
KYOX7cBHNwhrvysLKvezCbpZuWCPWXwUeI/tL0XaMWkNRYa0BlhVrtrYE6mS
Yl4QBoC+lZLr4ONKksZjzZr4jbFo9asGMwVNY443vXwlT//KsbxwtllKmn5+
zCyCTB1LO21Mt0Xzv+ewPWCnZx9MhmEpOiXxhYbQrSYYka5t3CwhzDgUmZAn
Pf0w3SshcPGKhMyagjiz2nbjQZ4m/WJ4Sm5TMskPS4WeU76uKCTQf6E2/w+s
D3ZSe5i1fT6lQvFjO81WywwVM/OUz0YBt4ttFsJCl/sP69T3W9tCgraRMhbT
s5Ao/5/UnB438rrpYhsNtZhQkd0Kpnd+rxG78DaCN98d9cFIv0FbJgiROnvi
tG/XyKQJQPfgoiiZmztanGD3VfSDa0F735IRHsRqH/uPVEUpKyaqINjMXLly
tKXBKZj/3CROUeZBBJz2qGOGDWaoiGY6okhw/PWJ5blA92N+SuiDj/55Yd2i
2xv4F3Ayv5+ipiyPXq9k1sPVvwgbgKUfHTZcz8s6r06pfWjeSpEPEfqunC8J
plfW+n4xFwWr4qkStSFfoPU40BKUpdUmKDTm61NrsWDDbH0qc27f+JTARVdp
L6IwNgKK6mSEoiO6hTapnf3vC0+kF3hWWCoeKL3bVFN2GVDEEHi0YbTgiP6F
Hbl0XToJql/IjgLNDnWfOZE+BUMqhh/e3xeKSAikm9c8bGnE32AY9oh5gneX
WPa32/4vUvsgnIhtr+NmVdaXlDs4a3tE5PmmNVrogNfUlA5ulARWniLS9KUF
FdKDfheJ7tvWrhXq62CPj/JsyCNx9Su33f11ROuhbiMSJkchonm9Ys4ynXJL
llDl+wB/jVokYRlrMIIAqPfsprqljVkpkElADwB1WVXFofLb17mkWLq+L8m+
vDOOJ9TMx5Uwt/P8OcCUS2UbamohniNGZezU18nfd2050GJQN2+Kdu8PyzkQ
/f9+kjBZrbZb+Dd3oxKKhaDsUTz5rIRDnzxlpnO/61YSf+9hqxd6Od0wmIRN
LBlAS2q4xXz5iy/bkIrBCo83W3B9rKAC61RxELJ8j7hFreDVAWQeh3ZD3P7S
nhqObTBlvlf5nfMJml4ZDqhZ5OBpfStoZxg+orvaF88Hgv5USTJG4ZtCqjpS
ND+UKMUSi19jpa+A62VUhO/uWOpXr2jRlhWyx+pc3IqhXupA/29PhQcTkALS
SsfpvXWykRZXC/pc8zrq67FRE3YYZseL2To64YCdXIhmr0qSDKD5FazmRvDs
iI9hHnemEEN4cf4ptWdBWMGrViNgoP4c3bBm5YNzHlDW2RBmlu6TTOPZW60v
/602Uw8K0QH1qkN+ejrVmoiFylmpta4ZCyl8ypDrBq9XGVV2OsQGd6gt+6gE
vQjZWDuAm6BXEyUZLh/dCL6D8xaBSocSr0SgAm+qVQflpCASUWIEgihS4U9b
SFIheh1DQEprrHoKUXDgmvYZZGQiIhS5KgERAhVXsxeCb54+AKBKbRXeINm6
RjOHlZp1NRLhxZF7mnFs53E15Fl8Gs0UxyWww+Rn3jjtbpanng8dd1NwhIsF
9DfqkfgrBaBP0ER8cB1SY8Cxm7v1WA2hW633TyrtxpMF3e8FwLJzQTCpryP6
9e1q6JZQSZLiTV9ON13CCm5LIp7Pz0GllhK7uPPuzvOljObFiZmp3iTeugZZ
WZhPkBUN+PTjK5CkvWQd2Yao1sNrF9keVtFObVXv0mqZpAluVeb7FFIHm0lu
y3gJb0YPG3H181t/KuI6XQpBALRh3Kcwk+ryh2SottLILIO0hg1b6mC3P3Wu
OoqXNZGrpw22CIB3p7B8EtFe1/h+dNR0HFXZk9Scf6qcopcayKh7EgvDfyKj
t9lXvikZ7G3DAeOMT5a2KisdMb1jKdSj8t7z9JKAqU5+HhboV8dFHw3vSQj9
AptZYfM/sYFdnJu7e49j9he9R5UMWjDw1JYnKAxAwT/ujOEFkHcnZ1RlnF4H
MXVy15rQabBdFoup2DYPhsSn4a8X05IqD3AtZ7gmbPvJVGw8zr/zx3AnYgmy
0iq8h0TCqaxpBOLNL84BCC+3OR4N0zvquZDYak9lUQUv4MDyTGUpqtNnioFH
AmSRMgvAb0/M7lK7FHKojAY2NfLX9T5iT7PiBeQjCQqXrFFO4cv6q1AeRQ6I
qyRpPOEPNNqt0t+2nYqPYlcHK4CA1i1kETJXuVu//Qsso8LdOFUtzAK7IYPt
Sxh8ZyO5Fy39Y7n20K91xVJZaZ8pWojzMQDyiu1JTjKS17IAX9BQ+7NsKBDl
zN8mt+sNjUJGaO4V27SWPglQWyU2mHSzImdHLis9wg04lp/lDyLZmMGzkE5Q
zBKYi0ztx+iNlc+gon7op0ToDynVyoJY3cOR7tiVH8j8KOpkVGz1WAX9yMFD
OCuDRN7/yIqYdpuDrDokGhqtRZndjdF93M9lCVu12xmFfUESqiLkleXhevxl
jSKu8bLsZdDSfrrySz5s2ox3yOgm4z9S/oRGtSUCgUOOafsyy0U+zV5pZA7E
mhgxecErniXWaBCW8eUvz/6gnWGGvWPG9dQXuDydkqxwAgFvyAgXAwJ1SrfF
Xo0CV0mSjEz/bo/5RUK7FjV1wCimHbn6OPwW0r8NKJVcVuSt8aBaCn0kp3sJ
j4pk639yM5fYTRyO2U4pLljWGYDEqEQU5tXBThGs4k89w0oLBlcIkafcWJrT
275jva7KLL7wYKbkXFNzAJqzQ+JGXSObFLuHnl1Jda7r6wvVX/kJRhUGsUnm
LY80bP9gj0gAD7upZ8sMcasFgcbKeMa1150uemWcMGgIC72eIei/I5aydOU0
vZExIKkXg1fvTt3CvLM47N7heNvJQNC7vlCAFncZsQxQX8KmpggmK5qVnMNJ
oRoklGS+KLBpX9V5Ti+OZWd9v4NBxDtX9OXEDh6KMFjpd0UrsTVoaJ4nJ3Y4
RhaXfM+t0WCLZsUkcOaRNbhtdocmVS9v0PJouhsA66rwr6aziB+jB05ELTef
buG0qiEgX2+NgCYRswrlkX3F9/qIWv5Y8e3/cFeljMflTOoEyqMDmlvl4fm8
/lBcEYsIm/P0WvjuiqdZ7zsEAiGSvKuDJ9igiwkaZgIqEku0HA/qNttAcPKG
/qU+IULatHNSiSdQOPVj5WFV8ckax1G30YvFa8PpmFdu/3InU9bvLHGdMA5e
0kalqSWRXBPM0zVYcRZCU/ceDgmGm+QlvNL3F+SoA9E4m7IJPJ4tuKvaQdn3
z4QDlhrx0OPgwMGOlx8kLVtVSgTPFlNMumVbPlp51BL0VK6bpv1c4XVZNBIt
l3b+KetzfvW3TO3350u7xQMNFUoUsym3SAXW92AEBAccwphrY4tfFpf47t68
uF6AT86mzG6tFzjp9hgA7tWhul/4kySPeYbKsbkME+NQCRmcls9lbgr+sOhV
K91TlpRooE5h3HDK7sqY2Mhrm+xtGGfj8bpgNvSj+4xTgzMAU2J8SSc8hy1o
LuJ1u/dwTWeREiyLdzC748NGHPvBioF0mjP2HQ/Z53CZ+9kwi6kq8DH2EunI
Q20FJFySTNZ6Qr168hChmX8PVAFX5U3bzUjyDKo1Dkcflw2pHniBzgDXHvpo
Ipcgu8FRtEo58nbP33okIB/sYyVDKP4WyfT/9qbtMo9NTGO9HiQiRQpTOl7v
z9KKnfglzHz34cuZJuF0Klzh1U6P+gBkum/reFmfLQ8hv7A36x4vPaU6rtqY
5nnr37YwKTo8Jce9NURHvvQ/LtLoXnittnDBYI5ElawX7+Yp4q0zY4SRFZBr
5ZFO+19lEGZbtK2XyKqtm272Z7eKjRCNyq4mVPp3diW9XyL2YzH4/xBJ+syW
vU/NfoW30y8tDBViEBlhHEdFYOYvb+Cwcmna5c15xO1sHno2v0kxb8UBOH2b
ZbhQJrf1Ow21KCTA6kmWZmuJhWJf7kzkogXJoNsd9ySMU6w99odcg78JElz6
h0wG5ODFMf2Y7ToM/MYws3yyICRxL25FfW8brbc1LIqSi0VeGBYWo8cwBD2l
DFWfx55HX9ENgv35sQvbDC7sV3PNHpLJg+DWWp8V6hJVnlPs3C/j1k6/ccIh
9P1HOiR8iLeO5hhG6A6UhNIxx4cJjjGi8BF0HP0I5B/oIsj/Tf89lE2xYtQz
Dc4csDm7AIxFwMBqbVF9QWS2ribUQUAMlRAWKb97BT9Cb4dbAIzitaMBv4Ka
aOvnLFYvLb02RLqkKpVLBOAlH4WQkyxTxdUm2uHq9SBV5o93Ltd7ItYuRn/M
91teMPd4FNrfbQWUaL3PLtbcNsj6cb5LrUoIO20WjA7NtJocL0p+qm8pUpRk
7GHY3t0duIG3rlGLRCJcxNBESowuK67qcKuO7I8H3LnYxfcgI0Galr7JDE71
fmdg86JdJUpse8pWzU1vZsEzWHhAcSj++9vNeZz8+0epQmA4c2nNtx8HJ5IS
7Sk8/24MvVZaVTTWFnJjJQsmZugUvtStFo/GR1i+FoMOT1jBKPWbggj9ZLrS
bAL0cnDuUlEEmXTP3dwlRznj1l8mSqbdRYsEIKhJn6sBxAUrBeBbCMn1cgGp
WydFY2dXsM1lCjrPeif8cgLQe7JjgT0quBREEEnwrsTEyaV1kuVfXyEIUU9l
5HpEqr9CYgMHbgm1sSFhAoXho+WLBgI9mfaIIYxrKYApneQZ1WT/mQJyu9jx
FzzE1o8vPTqQUorAPmEYfVcILjofBoVF1QAwD8/B0FTY9k859FcqsO7F9RQM
odELa6u7b1WR4+wxMg0s43ojLQIy1fg+Yg4SBMen2DTuLqaHq/siKGVFhab5
GwNeRzxErDdk9NYUKXQpf93hE8trBJm5v6uA9dYiB9MsALfCnHrBvVGctBKk
n7pYW1d5A9NK9yVVGO+/nsYGz7gg4ogc/9eqabKf1/UxICpyF/GC0weLwHHF
LNIey7Cf8NgDk3753zOR0GDoLMt2UmGyCwwVI00w2qo1fkF7t3ACY3aDUBHG
c8IJtUE78GokFuX2LJCvSwjjxB0VID3r4dql+PRlK7Jq1aAnURN7dORcTkVQ
D2JoTTAZR/rlMyYGsl5Xcy2YquzHJ/mH7ViyDn+QREdXItr9EwyeU80Bd8Oe
3Ut1QOA/u5r5lTAyQj42V+Lzm/3MeoMBw3a7duPafMxRmuERqqLZ64j0jtmZ
p+vcbXT2C4Lm2kRH6QDqvITBg8R+cIzA7PKv2p8dFTFtG2OHNADroPCQW3zn
28SsJ6SCTdMTh7S2vxudvF9JtORZm1DU6mxEUaLprFPT/gwB7BKpNrVQ0sbZ
InChzHeViDhj7Iv7GVO8SZ28G0jTKtH+eUMEi6KrgmLeMSsOUxgie78Niq9m
y+GA30P5G4uDggOM6afvWteUZ4uFFDLGU89DsPV7R0SfYeRTRPNaL1l2BgUx
MEhPi8W1ydTKuQmLv+ggboiK9+RTbtKn2jetNfhpDdChzJacQUXvcSyGYXtI
4fG2MsZzGymOX6wxjteJx0PEFv9eHiZRA2bMDrYmLm/w1jSxqkWLugFqXq44
zJmDMEcAu/SKK0DovxSyy8oYduimNN/FNWPJu1gda2g++ZaE17sLn0ZAtCi2
Z7HHN0SutpGFqrEMdVGIzLGSIrpXJcyfQQeKfewPMkOyoosWlf4bgGJdTxXW
/OFDSAGTf+zO0p+ko9Ay9ZG/xUWHpu+xvTF3fPJH9dSJ03yJIEEKECJ4CuyP
jptjiFmNIAuFOydP1e7Jfk1zp4Abgq0lvJPJypeR9mHtbK/Y1zhEz9A/bz8j
AtfL5y4ofJXtg9wHD+K07MuKOPSv/wylapeG8TxlhO/4a9r1K4gK8knBAHN0
DHnVmX8JKST3Uc9rE87drSwb17t3PNOUS/YBD2zUbDZnRjqx0lA3IqAjCfwa
iho977m6Zp1sx70wxcVmkBvtkgu4Uw0lTC15YiuNTbTD/M60tcHkbACkpO1T
Kay05s4sTRdoZvJNp8izaed1+DyFamGxFs8vTmM2AqLryC8aFDlBP/vXjx/T
KyvHY/lGypX/tO5OsaYbTmy8OgEZLGCuxHLOI9MV8P2w76b43hCkpqEx/cAQ
N+M4sS02jrThcpA73wURG0SrOP0FNtihHpRZ5I0xQWc9VuVwMclSdKLxHfzF
24c3VnYDx/8jCC7PEaYYBufMGIpWkAbAGyVdy0jamnQf0tspuzETGRbf2RNe
wY2KtikSeHkFSyEL1Z7c9PjmY38xKclvEtjCPTia9+SssjN/mUHOvbVR0NN8
TQYceJgF4MMVnLh4UIkxtC2smtA7EOP8A1SiR530l9ceZEt9pZP+HJG0g0tE
eeHfwW3wuw2yCkCwyx60g7UHM/HEp0guMtWfJMKpKOL5COIsqHv8VQF1VwBw
ZG/hfPUJmhuWEC20y5jpsRJzpgFDy2vaq3j3893R6m9m3zj00F8CVNUfSy2D
5xggcpAYptIyX3IIvVrmGJNRqUN/Px5HK6slFq0dY6N8m13mZuN+lyJMD9Y3
Gnzd00rvouYaBdpV3Tbw63azXBAwSPpRodVvrN/ilTA+a90BMiwLEVBW46g3
BIzEEPDLvJRB6bFueKcdnsFEMIH1PW9HD6LglzV2pselx3CqhfLKr4uhupJw
pZJuAF0OwskAxNa6A2+ab2o0AnLe4ragYtU40i2p/K1DxM22QMGBZy8ee+T2
2oLzvSOGL1Xz9ik7qwhKWsR7KyhbuZ6fmHDk9PVvUX6tk9R79vHRo7PF5NJG
uYSKb3T516MG16E4uell+wvEny7hdUp/X32gN5ssJz5m8OWvLJNKlnQ2YFy1
Yd2+QZCsWO2/1NRPMAn7GsKvpe6vJMovlGmyAb0AS4LegyqHy21HTQn8/3i/
pKuDW/bLwPvpX3+SCHUC9NOLxG1kNO/0civXdOAVt+tyLGXMQelHKNbB3gsS
2op1bt/zv46DLcwVekd+5S8s/LVc5cDHSPfHjWOyJzcQxVWwlpLduhfnv+rA
eK8F68qs2nlftuLZnX4Cas31IYJQtMN4JqYkxbOAFzDqN9wooiA4BAgH9aW/
SFE6nnra9SJF8Uduhj+2QIxbp+OCOPg3f6gQekRGDxNJxE71+u3rsmTdaYYP
qvdCtSL1eigZUQhGZhy3ZekU3QeQ7YuOOLObIpykOROor6QGPxv773FpKYgP
2iartGz6nWI0g7CawU6wFC/yfOArOllht319TTAJc4Gg6d0DA4DE4nPnglQi
++/4agj6IWA1nCl0NGskPxQnv4GHLr6OcpWDyifwIfoSOyKg9fdrNnY5dK5b
Mn9XjgPwEiNuMTXWVoM1reqp1EaM8/K/1J2R11iBHyqHjkrpXABw5OUBaob6
+Enui+8F/7vl5L9CQgxQFXDceNVWcCaCYO8ewv5RuuA4TbAP7IeCPQvu373d
vIwUVowfn8BfRfABu70eS70KRQmG+Z670pun3UUlP6ZM6gxs4qdOcFVSRGEk
WlFpFe2AMO8a8EJcQWqVztEGhrlZ7n9KyJYiZyL6SKmVuURu24RpVAnv8PjR
TJLqi0rB/Uy/BT/10Le+b03R5ltFPN0hp7AMb6zSREHGinDq8Ls6H/PfCp7N
MqasMdB7NWgthQ1XyermMSQgCi/QVD2I865GXOXcEz+F3QIgRwsrfPAPKaZT
V3xvLsKxYKKLUdMn+KXNUKToGsreba83Hk2G6I+Irx113QzKO17I3wLFgI3P
C/OCkfPXhN8R3GL9Ny7l2Q0IhzMnsn/XOfgRn3GqHtYBQayqYn21iAdXBMXE
6pzAGsnPWssKjzzEKFPc/8Xn9LJ7ldEJF+dSVizX2L0Z9Vwdl4sIm/ZNTwsb
bREXxTQjFqYs0FINKmIKVw9NdGahdoUlyl1xieUk/Fhk89lQI7vWidepGN4w
KZkkgV0G5k42yzXmbY3x9MLESOz12/e8/QhGkoE8tfcVkY8N/Q5DmdnzOJvU
96CwdTLUNYs6QvyfvG/XLgGJ+WLr6o8pKtu5rpJ+jtZWZeE95G1P0x47kobm
E1tlHqXKHTcaK7PkV23SsNUhOVIfWAV5sQ+IwvTiDhp5VrELEprWTXNtv33K
HHzpmhcRfhPo6hlUl4Kq85AsL60E/plGjIUb1/MmF3tfKcVoIHrQ7jK6CQP9
5kvru7UpnO89fA+fRdNjudNwFaZjjucYnFqSs+141N1G3q/qZUQE77r3sDNM
B6ldUQPzsmOthVR3BPHu4b4u9S4ntfe1OOSgOB1untJvMXJO9Fq7IzJJ/gdC
9MSPe/t1X/XE5wUsbiD8FWnNbnscwaEzlh6afGuDyBenkjK3kgFs6m43YRFN
+E4SaPBh7GcL18AnSsj3SKSYV5h22Ue3HD7B5AisWfsatbByJ2KQyZEefbeY
gMavgbreDhSU5dGZ3hBo0Nk7qyTFYDEnIFMsQrFygMEIoZf8pUow4g/A6cr0
sN/uqVY+CCyv1Ww3ykojQhcIjHuvslYlXl2G5MHOByQuZKLCfQ/4D2r5ljls
F6+mOmzgGJ84CSRC+XtIJVFxClM8EgyA90v+RklyhdIdNN2Y1tLu6r54sHFb
b6w4Z6+tr5uNSTB5X4Q3OWmlfppUWSFhbx2O4+n57g3Mylyfd8Hl8P8Y6Pt0
yEyXWDR755WJYaspLFaNdANI5gldHaITiWHxmx0rXIMw6jsLI8gPQZodG3Dc
7a7fHEchRwkH79yvjQlkhyjiKKMQn/iZW6UtLCsaa9+E4/vRFVMyx6Hn0jNF
UbJ+0s+dRMUQlWmJFRX4/g6wg1L4wS154JqJKPtjE6klzcXIGRFUkguDZH2W
40T827rjvwWA5PK+I/ibdCypHcQwk0tC48BEp8IIaQsKbZDQwMb+vQUPi8rC
q6Lvtwk3w4qGItKAQqcmBTWIYj95TgDvUZcpaLMYQnGLJBiuZeBUjkKbt5dq
B/5H4xacjt9RJimsVah1FFDbvzykWlVy0o285ystTEUFKprOLV0htzNqoK7l
OvevEFFLX6h2fuPVknMQz08NTLt632aQfIaQ8uBh/25tZNwx/m/e+97wHxE4
qL2IjIaqFASc/5EMtLnEUQIKBKnnqvh2BTStx1rfrFxJ6Jm+27TNHjg57iLs
uK6MaCX8KCwF19mCo8xiyJo2i7pOYDM7lY4wGqEuzps6WnXCNEMPsKBgSp9F
Cii4r0mWwV15wfHxX7nbIPzOdgIZkgws2VPAsAOggxKCNL0XqXfj94H9MJOe
MZaTJpyBxJqE/0FfGiTx03K+5RQ0ux+WNCkkVEG1Nj3DsWANhL4zklC9ymn/
X4Df9WqSu28Kp6PC+fYeYC1PLrqZSb8aMgjAQK56XaGSw4r6EqPVSf1N41eq
keYatb9lTzTsazKFlkJsnnHWynU7Vc1asW5GSBzFdnwNEnOzviFHVGAwE9gS
xv3kYPLEC1IrMkvgZ2Ube1lk5CmMxbDlgd+AaNTW+ZuZNZulJrDM5/441/LH
0rUYY+CVQLLc0BHBVSWXTGbsH4CHC4imLgEZLDDI2yiAdiu7AE9WOKFzkpUs
ESX1vGNB8afVPjuZ4zL52ZcKixxFrNXBP1dah025/lA5vv0a/aywurtwY+SS
vEsyU9+tG05OaxRl/KrPylD2mIS0ioNZTDtruaCN+Vdph5rXRA1debK/X/qS
TfRDJeE04gFG/kYUp6NQaXlMKEVyjC8xWAJSdAcSwTSE+Rx3Rt2KRWFjFs5B
+7rBav00Df+W3MkU82VdwBnhRsWmSnzD1f5TSOg3cqOUSVwxCS5yx6CO0dcc
m1ohx5jsWY4WhNCT73/NFgK9x0/A81qFUVOH60Rgn3NXS86rJ/ng/48WmrHP
XRop2LL2z79nZxbtYgD8w41TWh8rVfxuGdr+gXUuKGqq4wX2SKz2qo4on17s
LcQEfYlMo4hOIY0Tp3RsHT5rUF4EHJUxDHkClzfOhk5C0a9Y5TGROA4Wbq1H
ZjA0FT6fjWB8Iwg1fZ1igTpCOLL2k1AeFp9CcPe8wAQQc2JKriHBvgbw8uMc
t42Lty7zVgyVrEe/kVy+eoxbFWq94yGQGF/MGjcejAsLSXwzbV9YfW/yLkWn
tPWP2Kt7it12Q4Njy3TMSniCwoU+UNdTyt9pQfKhXL2fGLep6R2E4AxgyA6n
dvLb1xToffZES9fVxcnTSZYkJCI4PqqeXPaG5+evdCNNySt35GdhhdGJ/97f
idrZvIPD1W39TL2n0eBsAlr5fHt3NcSqd+0TuoU5D3Dkk4FzndWR8e5NGaoQ
IyLEAECEBqNPET27Xe5DhFh30a/1ygSdkkxhFo3CyWfj9J0C3EBKsmxeOyQB
yTVZhK5mAuDu9WMiuGXzHJvaB98zm1Qm6cOhvzeY0fhVAf5Xjx8YqD9ABSQ1
T+FGtsVse+gffZX/5F6U8K0cfvgwg8dyRgU8lkkKfDq21UcsU+o1WmYR7PZ0
rQnOSv2ccHy6PMQx1GbXaRZq/OZqmUrUg7WwsN+XeORSvG2Wq9EhJ9XyZQiV
gd3bzbvmU2DyEjgaszB+vuQT7l2x8wU4StHhAf0vGAgiSaPD1hnwZtopMJzq
LCGvWQQfY77ZVqxPIYtb04JXF3Eb9/iblkFK9CEFVV4suffXuLFe90Qw2Qin
AuFxn1N36yJpny9REXZK3gaL3dwlqmSkUwSlemK8I7oYcq+yD0yKuyZRMJBw
tbcpEEcETL3hW6EHq6YGUq7whI+JwHPOz7BZmx6p850usHppmryPiVJh06dG
+LC+ed9/wrBIf+wJvrnHfcp5/5LBiP1yC72j1C+cMLud70ubVNPleN+PQ9vn
w7htgpG1+Pj/omfOa6YLORS2kqHuwf9De7NX4zs/cRXwwgf5eoubTWfXNr35
FLwpk/iH2i7b9+9Yx2WQYuZOEeV/6F28RJ3tZ1arsNxmMOxrM93kQf3zF/wj
6rbCkQd0qZjHXHCnKHaRD9arAHJNwwULYikITFx3KNAgBYv0fxYhWXhzR30s
feDGHVyqTdV1j1FQf85ZjUQlZXcsPsG9HaXyvEKAhSdt9yhR9S6P1ZOa/eSc
1I6tAdppfDu1j7t6kcv/oM/VRXh9RfIQvt1pFi/gwUbvYC3XiGDj0jzYSMTy
seOpzuG/enipd2VB3tsauSXZeokt7f3UquMLGRq/t5VxX2yLjZ7IcsisKUml
N8PHPIBk1NeYgtbkZdsYfFloB2B0zhV4kBC5S0bKCVn8fE2WHTnLLF9m1+WM
jlUQV6adj8VhKUthpIRzclcd47MfD+/il6yIed6WEhSWbq2wjsUtXFnQHqSq
TGAFdsitw34YkdM6O+ldArOEXxkzsKllhTwjkJCqWmFy4ZQY0rb6jixmNJlU
ML7qvX2qSXUt3BkDicbS6jc2XeyhqkaYmksCMqY3gohpE6qY/QJubJrd2/kE
MrPtp1YV59e7Hc41mHwzNL+aMoQwVxIH8EXZN2WYFF5DQ8BmwD4wwKttLOEL
M8HmJMkJPYFtgiFqauNY2MD52GfClVcsqJqPvLtAu5szbIIWzvRNX2lwjcRT
LWmsyxXdA1QCY8/Z4tzugf45QKzbJXs7aghrFRABPmCWGfxsryUPENTKJ22D
jJYyKroX8mrws7caM6TrsvpemjgWOdE06zSCJ5FQupON0VfKl88vg7ZtlWBP
PF9ziqNsl3mmRYmG851qNJsG2tFBKz6jAR/t7gUOmdRpp0KkRq6PGnWYjTer
NKdr3AIUredN1hXE3oGCHP28uR19i9hG4FKgvAtYY6gSnOhwlBc9dv3rNrPT
g04dvC5A5eHgjXILYsxnSAZxj4PPmbueeUoQ93h/pBq+UY6BuX4q7BgII+Fi
8/OTZLJ4JDk3okiOg5JOXFm2TrLreZ74cBPTE6+wMCF1QaG8doxkZV1+2cmU
oWGCeZ9GgQ61MnlnGgen7IDs/hHaD9BqaHFXf8SbB01jrgFq3TppjE6yI9e8
KsLDxma+X/5efoe/1Aph5xekdoN4t7ZiwctUTqEozcCYQ2epCA3FC8Ny/iwd
Swi1gWeXs1YODez3xm/fAaznwBj56k4AykOwVhxxqOHF04Ojb0HC7MC4x41Z
wmmdNNLsn8XT5NAjR9APhnFEk9N8vu0OGQzAhp5fAYlVC6QjiL3+pq/i/121
uZ6RkBmXDo8gvcgIkdAoAonZGSXwDtUVI/Ldpl6jLAbQa4nkt1VlFMGKY6DD
xxM9VX+Tf4jfZ2LQy4+b5DdbajaMXQMOR5smR0z81PuoK35KwZhoV2LNEbOh
DwfVknD+l+zB5jmfLq+A4M/0EHelJ41KQvD8UBT1miB78ESKxxwPLy52Gf0N
EBIkR7YiyUfpCQQxW673gQeP3fQ6HV0a6Z9ZT6HSOkvD9rqUBluCuxDD0vxg
SgofA/+q24IZMouuHJNuQ9p2W0lWdp8+ubhxb7uzRqMMqImDEHL1Bw5F6NS2
vGp94pMrGTl97LoytNKvxzzuS3AY6E3rUJJRJp0eN6c17aySCVgGnWHOT7oa
NjLXoo7BBc/LPjxltfpvzCNAayYw4CdQF2sciWwTWQD5Gc0JVHKwVb50HxZf
lnSMBJQQ0IhXvCmTtgkqVYTz0snSHNVSt+ln603tEcw8Puvv1BFK41NVh3o3
x7DyBlAoaZX60tgdE0cxeIkm3K2ItECXYdFZOJ4I+F98Rxmw0RPzWy1Mjn1J
7HJa72VpusoC2BU9dETCXCD7TiCJUtEpjNoRlzc7VBvCu4p4LC1egeIXB8Ys
xxQS83Ymok0sqbQ1iq8mSU7cMm38c+/gjILeBRJCMRMGcHxNYorUOOdr2rvD
xnAGo/DQiOqebFwXwhANyjn5T0uOYGKiU//Fbtxczdo9G3/IfjkNUC6rfazW
qVYXjHDcYuTIJGMLcQWUWeD6vRiJ3BzgRXA8e5rl0EDs2+SKkcJmZgj4xuEW
9IHd7nHK2WEKWz7SQNSAxdPDn8sGTFFhLVvMkHQfRAhMyz3amapUxDDs0s8d
eXkatJs+6uMSNaQkwj+LxO/0iB3w5de+Szdn3910X3hw4TaN7ZRnbovn9LoH
KiVTSVxaw+S+Qqy/6BfpRlg1hqfhcvV15wBq5VXrYP6ZMozklVtXMQ8MEu3I
+Pe7C+harvRChAT0G/Xs/8smFGLgV8H5jtqfL7NdgF3zgQ0bclGHFlfWJIH7
IOHX+m0oJqEMCTKel7gs5SBsxG+zymMUzsLEYv3BWZs1O87sxiu60fHY2Inq
fZVM8Eu80KHs9JI8QkTlCvbmZgS8csL6hDuAuVahDxO+DxdduW00Dy9WWAwR
V+Fx75WLTTIaiZl+bRQCVtn4qOn+pvQ6uHt4XLHQPvhYeWyQG02CMeAn/HCx
TVtAnzqjVCcCjAsEeKXKxbcpNvUdBv8GIRc+y8mmK2SdVSZrJkXJ7gY5aFSc
g8048BYH3GZn0Eh/dfmw0w4r+XNYEbAu8ehm4DF29/Z6VqLY6eNbQDmK9t6C
uX9WzVJr3BUh/a/c5h6Qias/8L0G250iOlg+n9PID9T/xaoan1WY1TyrmnkJ
87CCnlm2qB29bo2hyatMETr0j2afKxVXyRJUthcvkP0VTTMK34ZkxgDNlqgn
ABSBUDTjT7uj1fjTFDScisqNOu3W6u35J/nfkIbZQ2MoeYFrocZryQ7r2Cfv
RZZjZoKIFJABkT/BxCRLHZdnTdvpkJj5XY4Wn2LZh+EBwHjibEurfi9nfKuJ
gzpOk1bNVa2nK0cT6CkRvh4F5C7uJLs6Y7VVzNYpu8im/izs8MA7cSt8Nf7L
t6HfLOpOFR3mAxkrgWsMhT9m3zJqqjA7xT4+Is+5sReBb2O3hfCkKTBtgxyf
2RbxtozyA4ugI/Mgd+7IRWU9+r8N1odKPzY704z5LHUHfLObgmuGB1bs2u/4
UR55m5lMsTbMoPcvs4PAQcvTEQG41LEDc86jf7pzG1gkyAYLaiNRjtuIZs1I
F430xVANJhqLGCmhk7VxLy/PVX4Dxi6H1y+OXgVxGuredAXVD7Tahq2ialLa
BpICvNr9yk0GEp3KuKgsgM2DXm2f18CRskOoM1D4W7rff+Zg+xFmnurioeIx
ByFLjUW9CWCpa825IugIDipMyK2+04unOPsE/Uwa1U/OJOMamSSjLYXhSgaP
SRNO3zQCNMYwpv3thkFQMDp5u5eEjIY+6O+Hi8JSU+0l4YgzDsWp4OMA40Xc
jc5tVolN1P+Z38ATHGHp4WbgdRGDSwivxHDO94GGZujINL3EEp9RJjr0vI9v
HhBPO0QHCVf7WCAXY81mGrNw3DYi5uAgXTgVUdxtcQu3BcdhjYAlO+YyaBWT
U8xD5EiliZZeyg1/HzHUKxNaZeUXXiKYX8pRduoNd3V+RHAU2W/OC77nb+Qn
NQwCXqXuqIb0u14pIW0fUbALiguIAuQjKcdFneOmARuxMEZ9x1phrLv2JNH8
NPIq3ccvMoyrMbN2W1Ke8nPuo8H+XOPJC01rjCFb4q97ZljKhRPXTmXNdiOM
sBKG4oUUCozDyl/C2FoD9Qbx63QZjWecNMIoWZmyaA2rG4isFGM586wSNwID
XeCstdjwqfJfmqvb3pvH+fJvHLVqvw2wQLCwp+B1us7Fhgy+FVnffLfwF3Oc
GdfAxbUI8Zpu80QYfUKIf7X9Il5oJ7eLGbK1mAgewzZrxYgJRroCiI5b0ZYL
psS3eEYJasmEaLUu6FCXytGCDo1AS71MRO5qTMTweTFbEoJoYgR1taAbMD2N
OLexijkR3OzUMgmzmrC1ViopVNAOfUP/73Lth/k3urXoA204eytuTW/dAc5e
zz/8HhAbyrZU/fKt6hwP4S1wdSsu4y4pXJOM0T81NU+Satkh92E7N+02SraK
NFBDcqDTuIud1BS7FTysH3//IbOpRY/88nmijQOrvW4/tkGL+jB+d4jsktcV
nVpGfq6lY48fvjL19R3ZHpyNKehWKra4rZiJNl2QmDC5hCrhUKbm3ZM1AWxB
FSDVd2qnUKUl3VySqYR2eN7/lkRM5bjVegETdpjQPI46K6AWg/xUl0qJ0obW
gziffCq4WWcm/Yc2vhenCEvSnbX8jXqWtZGWSPKpVQ01y56JjCo7fOM2EdSK
vHv96xGwIiID3+bHCo5v7OHrOECoVgtgv71MNhRg1C2MAJae9IUOgNfrVLLe
Qg/YA2PDZ3D2P4Hb9578hMCCvvdxEkWFSamGr0RDFFQJREmm/OxvgVEQ9udX
TRvwleD462MJhfMgMeNE3dGdsIqP/qutDiYBu/zbcHvgUQPWWoCRo96v0KsM
TA+OEXQNEqgTo0PjrO8ZaYme++xYSPZ0OTAW1kQVwz/TgHTKZRBmcA6Aw8im
GKPEA+x7iidZz4tl6rGDl5u+Pw2X0coWrU8vyppRQo87GPQ/kosrRZo2/qaO
MnXYQXEX1cvDSeayqfHzQlz5m1gpxSRBkD1MI7Va6DhtIfViYjWQCba2jkiX
WFzBwhsIIvMG2qK7V3x/J1XRNh/eGqovzXhLXBDn70waL/Dr63iXu9Uo8ppv
/ecPWZwngPrHkXomq06HWnrYAkOJLYkzSce8PVShCsDTL7czI6SSUmcyNSKx
gqDKEhUWuLycKrnmuN5orOyTO1B6l9RwAZEWZW0C4OrE6De28JJbyJP5im1p
aoJBwF7dOU4TRhdnD0/5IFEDKpSkTua5iWeZLn++3/9h5GvR8q55miGZNxtH
6xrT99XGRsJQ2EKt0FHB0cX2xaOoc94eGoT2pBh3ljhC+fwFDARG11B5lt8u
spH4XZQHqG1pHKxolDxED3rAvc6f0epAWYRfQnh+oMRp9BJuGkt8CV2q6i0I
Z19J9vtIiPu90Y/WkG/5D+ruVZZm8F5+p/zcyLY6tfaxZFAYuThgs3DaA46e
niiGOkPUXozQoIO9HtActNQXdq2i+xRyuOAzinovtviMIwkyUtG/BWi3E41l
BcDSqpY0g1xR/brrMLUipDJY2gaG8rGEfskVZW0HJtI99VX34YaR3nFddmkt
ghIhSIXQ9+ipRvwpO29psoyBxl4/9Y4OkLsYF0yiBGH2w7seQjf+5R2i7Srj
byb31vXUTL0sL0iMozvkFNzSoV36vmaUaBSjTwJoSeHU9sdL/NBpRRQP7xtt
/k04npkfOPk+Rwtx1GFuOEhE7/R90Kax18PkDEmQiUlOr1CLg+TJSjewsMRC
oW+amEZn2/3SW5cDeewPw+BxLCf0nfJe1z/9YVZxHlg4U1lQZzB6e8dDTbPC
LzERZdvgMLcUX5E8/89nIXWPWH3FWtXGTOaAxfIPu0qa6d5l7azp8FXKhhaa
zNNMI0OAwrpgzjc2YoLyYbZ3yYFB9mKGzD9AvNKOmRQ9PZzxWjEnf1lLNQ02
0M549clQMQn6pMMer5i/7ehvk9AR9SWbVknMZvShDJVaCfeodajpmAqYa2kd
9wB6024AjzJC99xoRUNM6UKKhPYKHEYpkFPXEuoTHuQ0INaGFyqfK9PRZ0HT
SEkEZMYd+0Jt4gGYmMYcz1qeAgLiYBEVW8OiRzPjq37ozjR6qpe7Mowdwpqv
RpQmvXtu+DUc+hR9aSuty61PSN8O3YsTtJSdve2TpCDMOdvdkpH24Tq19XMc
pMzXC+CcxvXohRzFk2rufu9qWQ7eil3D52ytWe/UYGMam4kVB1lrzP58yash
20ct3jCOJozRBejav3MYrp+Yz2Hl8hfbjd4N3sGnSHeN2gpf5no1Z1k5Q5Xi
kaKK04Ub+hKe7qUZMLVKvsWRiMjUluaBNJmXH2mqTz0OAjYqEuYbzIQEQA14
/QNdKPJjewwsEv4V9wbQTWLVTzQg2FjxjKbTifFh4pZ4WlZ/SU/6e2viZjhC
lbIW3gBtUZoVP1wqrkH1E/TBak7p0Gk0YItHHPel4qlSKfLovP5HEf6VAcaD
091p3j9ze18dPIflauMj4OwmYkM/hnClTOuJrGghYxo6Z5kYcGqIWZYrFawY
cXZwAbRFYvS27yB9rZO1I/YttJRMHJ2nt7Y830FMK760hOnMZ8ZH+TRsiAeI
wRC/VuwrAvEfL+k/W3sd99TXTiDw0tPaQeRnWuUkzdp37cJRPgnNQF6Zmy4U
hvB9UxbXMJN0BWrsrCNayhZX7hKBL0CrWajB4zY2AEZqJUVwEtKEHcG+XaC2
61r/IucX+J41X3mM8KjX4cWFF+VwLP2YjqdoPbAlP0c/qTVx6ta3QVa0deJJ
FjuiQnVQf8/bDSd5tatL4ua7tmDStZ6JJYXgj7DtM8xtneNxnrRYlBgjZpDL
HSMyplH/2y0FDOF7XIUrxuD2vXRzC5UcNHOJbGKdAC+HxzeUL5bE1iI2zNul
o4CgTrKWb3dPLagDn4xHXnTTB1uhnXOK0PWmwhcHHkZjVS3zZVYnThVPEP/O
xcgG7nvgwUexWipzAaltSpayGRYzbWtym2VCz2Z2DFrO++00tTA7D61uF99i
m5nPddmGAChUhrqZ+szrhuy28hd6xz2/4juq75INP+EjWwrC71AqiWnttvzi
7DuWum8f2bcqGxFK3baAxlQTTqq61fwrvU0LebjQkeKyKMKitABNP5rm+U47
dQIQ6IevGSOEfLT+Ti3597NSoaApdNt/gKM/TLd3Dm8oaL5I/kf/RHPW3Yn3
ryCUiEA0N088LuSPZ9aTtvAyN6uxBILir8ycEN5UecblJu3b0cF2CnUC4N1Y
t+42vA2aWXBleFTNfRvBN/0KFyRG4L1LFhQZlO2QllPSAGbUWL5U7GDPBNcs
fcDwEFtYrf0ozEhXsvjbmzcwceR+UXOXPjBZ5jsdj90F5jE3tQuPW+Xprub4
0lTVEanpWrrtEQ86ESD6re5mzg1KbqX9RuAKoGSTy7lZuaoxWajU6gKc5eNJ
F9KcgKRjqOyKivzQ+Z6/WNiS0BJwoCwgFZr+3b+nt1X2cQZWYZ9LBCxhoo5L
ErWZ2tyUQVd1cbsWSoGXTi3GoV2Z4G7UUNgDFxdP/YmMUBdNd4FJjxfB8jPw
KBSz8Zk3eBgJ4SIPKmC2ZMwF4nWQr6pHA0C6csXsy5LfR5ZG87wLGb+dg2hq
F9FTeu5jSVfHHzAHQfBWOpxW2x5WtBIQm0j5d6d0a3EPiWC7pCArFte82xa9
rW2AdAqjEnqQEm6S5UJjgaXJo7iSS9e4uTG1jWp0/wpW/Tva8M/bX5Iwm+/w
lCNfuUw+LMsH6ClCjXXfyU7mUjdWnxAxn7Uk+kxkOawGavqJiIyOyPEy76XR
EwzHF1YKOsPE0VBWOlqQjQhdLA0f9AV/6bu3wlc2hR1BvELOUfLetRN5CwOi
zXR9ZS0V/nSBJk7ftowKw7WMDg2BmLT//Kod4enrmqN/REMWhLrW8vtCHnDF
q1XstxdG7cYjT8jqMTXIYyLOxM2zQqlfZhE0zJ9Ufqw8U9o140CR2AEQuaz5
OYQk6f6+uqlk03GmbTH2ESA841yl6p7JCKqTiFUN+/jiNJLsoWjTzs3OrjTG
5VJMN6cB/lJglzoZKxURPtFg+7SeRVxT6UsRT7TghqiNa3acTcO9mQhpaDQP
eNMWCNxMvQS4giye6DB00+C0wLF7K68AShLFZg5BmdIb2fbbmMD9qIlVuebM
fj4EnJpJd61UskPhG1/d7iIr35cTU7LsT7TXR1P5qW2T/QUHGpB66vROVZly
/WgKkrsxv472ykUXeN/2Oq1fE3zP5hLi8pMXI/OqYh1A86X4d7/wKHC+0w65
qoaF6E/ZuVbXBFohXp/QYEhxWQb2AfZHiv1N55n2DE8Cg1EY+koJ1xGxVfwz
tMsUQJI4RFoPbiPKQkCQhrRLT9wi4HJ4DjyNmzo9UbfQbN+RQ/S2RW7R7Q2D
raoJUzb1Szb1jqy8r6YbmRXF0GLvHQC0puRoSjubBKDIqq2xKqbjKqg6aT9o
hDg6bWrU/Dx/WL5FgiDVzWynzU2xYKpW9umnS3w4XLme3Tcs5yOE1svYRDSn
flXY6MQ22fr1msBZcrXm+CH1xmeZeFSWnAW6vUBbrY1xdplcitp7lJwAI6/A
vRVhu4PFJwZCb3wGo2hkQJl7q3dj6FEignbAK52Vddf8xyRXZNtvaRKluu9D
4bQtdfOBkHQIpxENcsr29mUsqbkNVgTfbqv+syKGYB0Lb03VwQPWNbB/2cLJ
B+nS8QFu+jwn0Tdg/+nTe2A+WGO0eKKVdl3kaGZJQof3to+CF7BRlfG/BKz/
VWjPViixDxUmPo6hLH2GhUcvMJKhiyXxqIaOMSLQ+2FxeYraiZu4Vx2Qa9WB
JCxkK7CTVz7dhgDy57iZ51IauYk1wdNAEWm1d27IA3VR5qy+X0LQFk7ITv+Z
irRgUc/SAss1SrQVH8q5XC85VSLSvMZDAGuKM4uKg+3NlVu87Yfmx5MTrFWU
sQJX6mJ4tFDAAZiZ6epDzE3rZ/7fvTD10S4146uaywNced37VeSuqaP+VIKP
9nfz8Z59x1oKvZaELjbqLetEsz3m7IgHUdaaHk0bVl+pjUtXyP4xS2uZCHZp
1CM1wN+ypVb7TNvqfGetRNPuWs+2LNUnvW5UHPU0jARE4pqktmLZf95duF+H
Jnwejiia2P3LkFE+UnohH+0IDnVHGtUFD9oAa9il0kJlJ2zygXf6jRfqK0TX
TPLVh/PwF60900pCfphJcaiDcHBZEk8Ct3ZRDfQpyA92xv2nh4BSMoFGQrUo
oKd0C18j+EVz0VPrAmY5XGqWU5EcBbQ3cD+Ci+1KMAPG91P+Ty9epjIWFANL
ijnIGqNmthPmmpFU7qjVeUCOnYOlo3/yTcENg0D4ylemM1X5dWJ2lYc+Pfs2
eF+jBmr0FvS1nrlNe6TsnNh5Kxdv8uv6cKE7SxZg/JmdY1AYfxDJFEvreVPY
MRF8BJpc7nJ5hfpHyXuhqeMVI+qoCO5DqATHfuJ1/uI7F4I9GA0scxWrElCr
wfwEe6F5NoYIudDp4Rwt+VDQxZ0bTwADIcwf8JiTSswUysTnsTScmwK8reRp
5y7jagy0Q5vMKHRHFuS/AsGE/yeGQDhInPxn9mx0DdAV1Fe+duoHxK1Fy6Io
6t9xf3xp7NadsQztuYJHCLb9ezjhAk45N787366h5W3kKPvwskKFu9iTc9Vd
mmXbX6opAdoVzPfKUydo1kvjjydx2TNwC+UrNfyqFydg82Q2wCSbQka0rfwx
GmaZxw4KrnYK8SoOPJSqsq2NFsUG7dPASSRgHI7ReQG1xhQV6twnkjc2wiYU
/3UB+6Biu57jxH1ljykC5D+uqQzKJI7SVAI8AOYyJ+NXKPRZNZky8XQxPYkQ
+WQdFD8Sn5SGzDX+J119lePjuZQeYR4yD52HpG1r/5tRJS3Chl/4jHrbphFF
aCjHPuSBjPKbm03YLxeqF38fFq8guGCpbFvKs67ZDLzjDpIk5agmuAhYq7iD
8gryl7xEt837OclkQlo95HrCOx3JTq9ByML+1icaNMvczjkZMMnbQ25g2ipA
DbuzsSAW12009XlvZdkTBTQgOF3KTPddPYirK5zggGZXL5YAlPFNGKEUVoHs
3cqAYeDX2Sg3MNJmmBbeyFSuZiN3FJ7SS+atr8136CMHiRiSEh2retThUyKk
gpIdLo1pO06ch9ouZkOSvJBsEdd+wH5Gk3/CIMqmDsThhqfX8FF+zvM4olwu
IAsRrQYhVk8i/aG9B/Q28kPhAyTB73vDaWxdSiN2CYIVDYjeZupyVbo6QG3I
QNWph+lnFIs0wLFzYVKbLvR/O1BLKI6ErYnxG6e79ivlE10/ZwsIZhMGarUI
iwuZEX/SPm+780hTRlh0n5g25wedQnI8wavsoTJWiJmK/G2OoAi1werjZ7aU
S2twMeaNPCkoLrnBZxzAO5Pyvdkuv7lKdzCJ3bX9v61FFyw6o7Xc+72oX2/J
2jUvP1YfeTRE3h5VLY2C4HoBK78KoKzTEQ0IPZEe9MHpVJYOT9NZcSRwwLyl
L2/toAfQzHgaXb9r/F9bvf0ecw+B1xcHNl4smrfONHDhcGzRewOvUdyup0rx
lzLg8G5bPe9+F0diAGzixEecapG/OZuvDvE2FD4Rzj62gWNtoTdzoduuZ60O
7ycUSdXro83OX+fGthiO2ifiXMuoM/rkcT9KPc6baH7MaCkE8+xHCxNFf7JA
YXlq6rTDzL/xmpnibxNuFdNJbr9atw4CvRuK4Nh4yj+UyotXgamt4pF6uKyJ
KtW6ABtArz47VqMUKAnaMlg6I0WxUQHr7UVQmu1IDnj7kY/HvFtBG1qB+L95
cv7i30injvg+5KMmFFR5XHLOQcfcZpTscTcI0dWnVj6sAYr3JuBeF4X1jJXz
GkKrGvQuFDx2MQgGMZWHM+r01GkKSYazk5dW7rZ3nk6NgwoYLx71bON2DpDu
rfdBnnzdFnpnZ/Jytr00AOTDRpxChtmReZ7Y+fHYYYKUx52cuBIdMBbCLrmZ
YsJvPZfgCsfLwStv/2fYfNJRI+/NRLocqXCJK4YGSIXTaVt6zpBIj8HDwtha
S9+gfdRH9L2ye8cMlsZvVjE+0ku4PQSyRCtpC5V3Hoetdpm5lIHrxDQ0GLyH
ihXmad3g3AjdcJpHLnzKSI1F6JliKg7SFcITCU4lJY6GJnZDtWXC0+epptlX
oH1pEDOiLGh12bUZcVBHT5LTu9YtOkgv+ZlK5RXl5AjAkgBUhEVBSMJ8cnMK
rOFfVwO/nEXDwf1wt1GVLnxfN59/tJYaF5E5Cb8p73rnk/vwtnE0Abx5vet2
Zq6R3hdZdYvtHlbNR94AiQBXnKIu3YiHaN3vkCNrfKqAzvQ+l89pvqKA8mXQ
IstS2iPWMabjTMF8F1SNPLOtROZq7qrsPJwtTt0HjGkBrlqxfe1WCiBcYbsX
vF4BKGDLL+eW8hlrqUDQyrkfRPL5sNxEjxCpz32XVq+S/9PRgbmHmA+6ostI
s/QEM2W3k7ntFRxFiV79XlMO+1J9AO+OlEg7Lw97zKvxduG0NPs0LnnHkNQH
aqK42gfKii8MV+bP+8w0LHT2gmg/aEP71GLrQzms/GyadmIeLWEP+z0TnjHI
Duhx6ERlhTUZyY+adrULqct8wGzgXA6Yqt/nSUOLIv5Bk4LIw56lztYFobxT
qNnqavP6DjHKOXWOx+oP5+u+97M4w1xtnFLmBpGl0yCqYeY+XbjhwYqu82SG
IGPMbWqJF2mD8KjaGawaqWHm8YtizADAm8WIQhz80JNeugm08vaLcaOlwvnd
Ha6HHZ43HnIe0lZebc1zoVnoGOfFqaFZstvS9gVuQkqGI3+R4ZcLU+zjqueI
MKjo+MQDxpNmmL4K3f8EOsIkjEEkGOB25Enje9EcKIZLeNHsDwC5afAt9TuF
MUxxCaqfPp/pl8cRXyiqfP2A7tR5got9UdahCT8J/E3GFGDOdMYKEy14H+PZ
wVF7d4QsRcDe/4oPGTG0QznzYB/qj4osndi/zzuwqprjk26FvW3z1sXOioL0
7BRMTKzTtDrr3Z5FBy+Ozvji8KkQyRWGNm3PL+WUTTLuf33xeCeuGIxuj/NO
HWovBQQ5EWAidzfb4VmsEr/8xS1mhEx0Ua7lMlGrm3V2M74dmHtB47RFChrq
iI/wwdeWFKHqqBTmSTFsJ455qaIiewcjI3tE8eJOn/LDB6178XQzTWabClbc
dus6NWF+v1duhN15HAk0YgKwtAl4HJTQCaQGfU8Lnmhrub97gCUigxbl4HVG
OCsw98ZL3TnCA1v8xn806yLI6iKORf3geICh2teiUMDgAu7gJ/lWJLQKFB8O
JcCUba1wvjOfC2eQCbrBD9Iq9pIrChq0eaEVk1m6eZ8NHr/adtHFVXc+oWX0
uJKPLWpSt+qnJVTiVGA3aIvS5GBd6BZweaIP6gfkypLAj6ZNusly9Amm+sTG
id6jB3v63sZEbHuwC09gT8G5SCx4F6Dti+2HsDFeSd13LYxbZtNVyFx3d5DC
ahXFvxZANXDbiibkvz0GLjVLWZeYH7nQI6fgXQcxg6TvA/1jlXVzr7Hkvk0f
2oR9i2WD/NQ2VMfOsVXE72AgztebtJ1dP2LvkW8Wg+Zb1scHIyILiwq57Iei
AzeapsV0cdgzT7KNGAO8pulYH2ICg93qhNle00PpmkxST+IQa4g0Zx1c3zct
khbfLNlB+kZPI0niTuJfM90LG8PFTxE/zyNf1V/Oqnv81ArUTWWW7CiL0z1s
2CTgQCHLrhIpj86onMhkVaHVmCrPtuiYiEB9upsLirKbV6L9IDh/3p/skR3a
HZLOvGJu3sv7diedkms4lZ+102sGTZtJvekOoTIj7KJbG6pyFRXvMkCr/i+a
7xWDKyreTC9i3yFqiWK1S+6szcYHcqlBmjn2y9MirrSJFqAuWqaiEQc5a0kt
Hsk2ePs/UrWc5VUipztgwgxyuiMlz+bQ+oluooN3jwl3Qy5yv0PmZNL38+Ok
Z0BD8ndfYrvCJFDO5XmEy9xtHwD88jq4C5UU4gqYU6eueeGHoOz9vb3KH6lC
ytCFF9bAOgYjILGasGQKrrvUvOyrHCzdiQOYuW30BVRJcJ7bV0mV/2PEsi6S
cXTwr+3Ubsf5sDXUeYfsDw/4KoyQGx1fUOgXMawkSMqMH3/NYt5diI//Wu86
t1iPtpA5ayfvsi7/R+Ui/ZvhSskLzYG1e547Ud+cFMOzyfuPq6X9aQrOOSCs
jPPG1p0y33iUWb1qeR5JZcrFk8FDB8jjooWEnDc6YbSEhTXJ4KBWCZz8cL1Z
JOT9T0+kXeFrrQxxpoaVx4SVqOrshgwoosyZMXf4UFYg5lMutTkJueKPEIqM
WHU6JS0GlEXVnNPQ/D+x1Mi3My0X7U7a9zie+wnIVjE7ncpW+9XFZM1YFLBp
7cqYB5LlNZOaR6YX3jhlnIX05VEOjJ8CX1q0QLEUaka7aBB40RmoAYfQJbsg
IjnPJZ9DL+CNnsS9VFYLavVUfWqHCGfa0NWpEQJbFEDJXXYiIRgiHU3aEeMl
5aLDKcynu5y7oWxPL6aS9eU9Lmp6T3UQAW39Gsdyp56W5BhCJZ/v7Onh2+h+
QqZpHuHHGj+0cQD68eWHa4NvIKip+Wa2WFqcRfNzhNjd1iYOTpstPeaTKTe3
+cpw+8Ajt+WNXAgHzIWLOFFS+hu2aUqpYO7QherJBCnY1EYrAmcXkxJjgP1O
SCAMq/JEnC6sPsXX90H27z8vfE9TtmT6t6WLkpOrhZc+CB7oaOhbBLiY22lD
75sXGoEoCag9O7Gy43IQvpxsTbmvrtoZVY0ZRuSFSpPRMM6eBWa4ByJCdGq1
ikZo3xsTqsjKhvv9MhPbYv7lS/r/+RTXG7DaQd6ejlCC4vX2xdDUi5vxN1F0
PgIbD2crletTXp77iNTErEc0lwG1rPzAi78Ft9qVHbsrtL3Bi8GoD0TLYcwz
CNMIR+jpge3ee9MwPGdBN11i8agslxF1tyr4lbItuBDr3S1qiBMVTdf8U9WD
8BwDWtMGoMBT6D5Njltz5W8zLgU/nXabXlto4PGRGR628sHRzAT7a24D2LeR
AaueOBl+6CLMY3bb/96v44zt+7kFVuwWQWqZAgQA0TRiVoxwcU3+UDxmvzAS
Kk29B5LeZGWtMvjYlpHeyPefcQsFmJzpQkCDP4ttpOsxGwkhtWYiHFGUXzza
p2ObDfh2eD42CjcfLsCNJaG8MyeFmWUtB7AeXHUbcZcrrergSPaLrDRA0NkF
LFv1qVZT0xj33Qrsy/VadHbjwGWUWWMuVhoHkV9wQtnGZlLQ1JcaqDJmXYKb
3OJo52KTf7jOfwPlaZSE+aZdI8vNdD6cfnacPRQTx0c57iQr2c01sE6n0Nz6
upOF3yvg9mL92fmvjQHsBd3yuNLVeYkAwoVPMRBU4xlXHTT7FFu5YwQL0QnF
mw8x9wDJ3NJC3PSVjJfDS/gEboKUpQeIClIneR5kuNlaWSiuzv7J/reX5T0t
Tz4Fja6/4P+KIm4afDwopnN0Z2OZfTfEObBiUoOOImWzEqudgwpBctMpF95L
MdYgw1eNWG9l+EadzSXj5FJkCvOtGT/nB4J/+Rifg1LxswHNeV/ICvPKLt8e
fA0cKXf4BLxPQSi7slx15+UAMEBDByk3xc4xR7qO4NUP+Ybcnc+PRc49WY0m
TxcrY2tWprpRDujp5h7d9BK5lbg1HCZT+DqV7GV6XUqCOKkWuyg7JvaSWgdq
WbqDSmrzfrvLA950KMTjbnEDmbgAa6HJWgPxbq9CLaXb1X6ST0WNyOjJHCGF
eIh9rF/X63wrOrwbP5nLeYS3qxOscI3oVW7CLk7LD8w1W6rgiZh5PT1wzNIT
uRkEPVyZi9RTIsGZNMrefz4wLFFuisLworl5s3VZ9treLTgttTJzRBCkjp4+
FwwcmIvkyKOlHRP/kEYgfuvMfDnxxHSVNtmI3eWETAqDvi0SbEBeYMolllRQ
+DKlOLgsTSbDsfKUBPktdG8e/lgp1G5jXLNvvYLc+j36h7IKc+zqQE8q+1AE
jLlk0n5AKleCSx8Y7YD5FhsFYn27TNsUVhPFBMMVmrdVsC9qaFsW3GQkXNib
wByKwkK/OqlVhKDkHvuu5xCcOpNYGXW5xInYFhRvLsEhaldee3NkJ1VNWCkV
CAIF7LGUm5723GIptrk0YBkJrVURUEUGTqLnD+lWyK5+klcwlWe9jxzDlp47
+q1dTX9a6EhqzZNPNkdCBmDcba1Ge7VABGIiaNcf+0m628rDpJGrXTI3Gpyw
R4g6M/NLZ7C2k10bVgBKCf847mF1H2/PSh0zatlKJThLr+yV0fS1hvJH/wrI
Omtbaoy/FZOZcWGGZW1EYEi5YS9D0DumrgG235k/HQnrPaO4M+xQnX9qc947
rVdWs3glxNNVqcE3Qqioa3PvImGSIn9HgMhklqSb5/RUQotG5XYuj4pgW5I1
4KIBm744FUs+qOqd3DVkdCXQLgW/K3eLQJzyqn7PhQlN5Y5+eV2DlXJJMFnX
3xSg5b6aEzAWxp84LU7nZAQ/uopdF27/Y8oCm3AiFUxTaqsY+4sWOFZNrOMb
rTqLkbyS4pyNeMX2L6AMs48fl64MhXUhdT+klm8phKfAbM4erFQecKMUMBbp
HGMO3pEdeyo7NAy+TQpJqilIdVeN2Oo7DtwCFKW8KSXCsjHzxPKrcHan1KOf
7buL0xsF3B0p8IyZ1sT/3va8iSA5FWE51HI54Ig2Nb26IwKAtXqeHX0zyx+Q
eUQuAfHpWL1eq2ZlNhow32hQ9dz8l/zdNdohrrUXXRZF/bIplRcZDQLDbSr7
UQrMk+d/pOwCNB8mKvEcdpVUxXP7Z2DEqVu7zeBdrR/WdE9nWSlGOLaXFrMB
G1/FPwYZzNzeQrj+o59FhML6tr3NgV+3vbNwIBivtvLHZ1t7qqHVzHQtsqI6
4jOicfp2eBhQ9DkNTDtWmgi4W+JVo0X2h6nKIBPAIPhZEWyKy1XhKYy5csW/
bKVl4c1MDsccljsctWZfB/HqEvwiFIWNTQQA6+skfI8WfB1j/DGpGjT+MbS/
IYV8zSmClJgdV6F6Xiq6I4VD0qNizsa5os2CqQQB8xj6oCrggW24Okl+dbRJ
9I0RG6/ECuxseRTkIWcPLe0WMUyZQRqwk69jZmCiXALx5MzTw8c6fp914POK
vwzPpeeQDKbjFUNWklFLnQ+euHeMX/5+em0NkJlQ63Yh8G5s85pY75N9s6Iu
gnXUWDShTxOT/srhxHL6h+wUYdyfR5g7TlI7wvbjruh+TzONlwcqxFUr82he
kAy8FLz+nGwBzDTZWipUnvgovWYtPfv+cs+zJ+NV8GRztwRKqITFOmWM96Yu
uQAoAfSdyWIxnaVE3c/rW9JFgczPQXvyQC9I4BKuFqJrdm2UF2dc4cURg1LG
ecLbNil5rgTR4x28nbd5eTrjb6eDU4+ac4VqIMK+AOT/Q2FRPzT9o9nq22q8
MZdpVlgeTv/zUEv4mMyTWjVOkcYLTe7zrr5uTacpmPaoYTNrNch+a89fr4lV
g5Pkhgql6UNKJgSFZk+HMcHCtBC/C+GlOksZnFtuHMJkpYvW9dnWU3c63y13
E6RzChJUnaUsQGBQHISoWjpOG2fbKoDdXeYo89vmKYTLa7RxXFgM2oKudDgD
/TCOOwB7oYNQvJSW5fMEUH2Q7hZK7Dwy30ANqsDakAtCgobT8km5BZOwB7y9
meZiwz/VDzwSnhbqv6HkOMmzL2PzVQSmsJny0tk4lQlwAm9j5Ds2wg1Lj4oz
aVBp9rZl0e5qyCI6ep9ME0TetSP15vEk4eE0F52HWRPNezaYwUPPgAQsyUKA
9cZAhVSwgGa7cSmljrIh9YdgDUXBwv7XPnlQl5To3npLe8wd0gCqvV87lNnd
eJry8ioJWqq5oYI9AKuyhRyaXOk0kxyK+DYI9dy63CRxwVgh/5CVZScJv5Ac
EDdDFOOeYjP8b4cYVShFSYmiDUOlx+9RZRMhSldMPgXBeO+5ev7s4cphwJfe
7MkGUUiwqV8sdjVAO28hdXjiwX8+nvyUrqHqpqbP9l7WgJeO14O/jExtyvAE
g/vaEziEvvQkI8mkQQeMWvP+bg0tMbp/iAVAsg9tKhr1MVfZWzN6jS3zcZLo
rU32tV2I32RMXTpiTXZ5jTtg2rdLjVlFhQ2HwZOtzossgMAhMBaW25r2+9X4
uiR5dJSY7MzAHXP28IHvBpWkpUW+8h6se24nsCX4AnnP8IdbkHdErJF/hwKz
espSVckqSl6iOX3N52tYkPKQY0a+RajG6X1BgMl6Z8vpG61ms1WK1jajh5cU
5yr/IZ8CjlRqY7B8tsja57OR8PlsujXlQIP7uimZfhHvlRAmo7iqNz5oEXql
8o6wC2gwVgGZX27U4lTlk1oTmA3z3X9143h0Q1Ebr6PG5S3pTsitg6wmGs1l
ZPmIHy2BXNlfHBHmiff+MLlcLGWg0Z113Apt73spaiGinzqDKsCB4y8Z4Vta
npxt0WOSHzqs7R/FWXyjyGCCAr+EkDoAutv4cRwUhw2zv3EqxemxRAR0itdp
WzKxZihuQpMU22EYaXqpXeorV0OY9YAX/UJDqpDSWjgd2RiWfJg4xS8ja2rQ
f+Oenl0eHFMnVomcErMbuTWxfYGqGTqkJJpAi0wFXJi2uc8jSmbTRMwAH2fA
/CpgsbCM1sm0GAVp4f5teVAbsb/1rkvqKVhKs0eBDKzuC+Z4KhynOkHguPE/
lv4D2o3J3L+8u+bZH3kBq0pHRWmZkSzXOLVSgk2koLVlJ01EZyfl/YsQQ5f5
Ftx7bDuuQQvbTjf7xJZas1w7vmmcgADLX8ofkS3931WsA+GxV4HVBZvtk/9L
TEpRm2Sy17jMROZ9z3UNBAVQYY7rHkTKbiBjJMCIzRC/pOYt+pPnBjbFVXmm
tIgaMiWaXJV0d9Brrs5swOpkb4oROKGmInGhDmmAg5f3J6ikQcbAH0+nk9lO
aNOB+4Q895hHe5asQwVs9sdl0hgXTKAIEntmpVanx7PgCynEdWJ7588rE1C9
ucEP+Je9jEmXADe53PxgEY3EUWwtvwMVkPW+Wk6Y0lTCtd9b+OXlZsZZRfMu
u2LBFHIpVuy0ZyihOiFyGkfp5Hi7sXAQZtd+tb9fsTo60Pqx8UM6bAm72YF/
RbtZxbHFy6or1t7KPhRy2UW1CmiTHmCcAjkpdUuWgFhq0D42avbXXtzWqxai
kSvP6Zhx/cASQq2NdkM5Oih5/YJ4xhuy/rM/PTf72Dcn59648nSAFUsrGCCK
jch546rGPJGCEzclMd8Cl0QFM+Rjtp4ydRd8ZCuzZij1vLTydjYl2dX+Ug87
PBlVXiWKwpXCsLpqBqBOOHAHGGoptRnAJQURm13g8GMb7ft+fTisdwqLKfKY
V5K1/JMtYXTK74dJMUPZ8B4ASuPrLu2cX+7IjFO9m46wE6jBEDarym2gMM6o
KpwKUxI3FkDC3XeWpDVD2jSRnptd8+i5pdCoI3ze/PAYSVI/iD5LGgjNeuVo
DMScqLLI82Ainf3o5ujg+1pq1OgWnhE0mbXiSFnfckCrMChZiw8ZAJHsF8kZ
6hoafAPkTShkiQNRiJZyw/dkMS9PdkfSjFCYxOetX2kG1Yb8K7oJnK+9ct/a
rsqGiL6MgBglVaN6gYR6YpK97GIsivGY1O1KV42RpG4+EDiqkrrhkQU/gx9M
aHEzrZiM6JD2xqfW28HUlaw/yOrA2999ejfjt4MvM5JWpp7ttqGKFdUa9y7E
6Cwy4qbqG/DeoZtvB0e3q19OruuT0kq6atwbVwzLqMDy01YvJYD8qJ8aS6a+
F1hcWJw+q0hSGbM2V8Oz/sieEvzQ/01z4fePjrZ55rzniiIBSxVvi0CbqDRT
uYk842xJpD/FArpDSq0uX5WFbCPGfL6uYWPZQtUSvOEV9ja5N97/aWrxLk2j
AHMvQ+NX1fppx628voGCbEr1DAQyYANcmHZQ+GxRilKP9K9gNsSsf6FcjaHj
TvAqNUyzL5LFSeAW7ufa6p3OQOvyQCeiXkEmWlBe5q1tfqJZ+38xK+7FQIZp
odu89NsFoady/1lOomJZT+xtxRBY9bLdiogxMmPK93rOCx3P077zRDomNCwe
s+xO1rmaCUup+NekCqu0hu+3+5r6o3UaVPBbgFSTKijY7vqDRihcS4aKmsYV
0kiSknWhYUYhd30eL7d7VvLF8EAiX1htwgjGzJNpjri0tB1b5N6RyteH2MGK
/Ij2Ezu4ztZXzxcA7NyaQp+rKiyghuBkC641pV+v/4qb8STfM5KNbinZ7WkB
UaU8SIAk8gWcOUKDM+45WFGX7gZYpNdRaLIujjz5uWsq0e3byAAkcQnsqLPR
JqXTJfbbxJOe7qiIBbzGyWsp6pB6y7W736WUfGYFLkhDpTdSgD0faiGXGKiH
QCXjSixFzn4SkVGUUp33JP5Nij9XoshjHgVh3BYQHvhUSJX1X+eckXhTDQ2J
d5LZ6vSqII5hc2upIFLH1F90ma3NEMVSTo9ca7/f1J/NxLWTeBz0MRjcISdO
xYaXeAcxLuJ+sqgy0+LVpZ9YV07qXSob1lLjO/U6TNnTi3dz6OFkBJXMn3p4
VL3XbAdsIysZfAVmB8AW+GhG69PJg3UwyVogCHN9GPyaVutFM1kNGQssai1i
Q4zKg6NZKW21ZIvrsv3JNrFHl4Js1F97Int9poWBJhrbzZU8dX2Gy21Lkb0S
BbhCEMJmO2MloOkU4DE8bnx3Ce4ZvxOTyJWQ4fw1Y8lRhp/0p5XQRtZSrdO0
Fg/iyyAaFnTJNm8RLM3USLl2kXppNLBp4ZWTy7K4tNvoccDEpAHq1PxTtRQa
HX3g9EbRLpkhhOgYcdk/VDp04D1Bgow3oa3gntdgPRrNK7gVM1NadSLb2jBo
c72lAIUxNCbnKhRangdkP5YpUHnCUuko6f++gInEjmBkBS/V6U+rkWairlcP
3Ty0W+a/6QTX99ZXGdZWSoWv793veLkwVqOq5CjnStqa47SATFf6UnkYuEhI
DUrBm0yZVDBzyXPimgbFbOx79Hfsev4b2DVMcoRX2m8ntLBvzJGGbJOA6EuN
/GwqCOHdihL3kDDauXXpkjcGO2mYaFvEpzOtdtk/gboLrTVUJSTZ4mi0mg/T
cj6o+uW0t7mk2xJZkpcG0Kdf6QOQ/DByZqd2ioxPYkdspW1Pus/XoA/YK/Jk
qDwP9W+x5sS4VWtGb/u50kjMUg0gJCGPnLfyMnzOUEKVRrhCV38/Fd+Dq8Yq
0n4OvlQ93DAROF43t2Op8MbjWfgcYrVNVomxquOXQK3r+6PKbgnU2TGmUbq1
092i7O8n+fRSjfUjAGewt8d2d0clac2O0aj2ZoFLhT8Xt9dVu4oyaq9xc8/A
URU9GbIwC307san8swG7Kh6aUrb51mHi9C0szPHyWk+lsSBVbqwSC+hWXo5p
HM85eTp59WkgLj0xsD+4bFP+aifetXFpi02ViglhQTJYgFEG3WrtC0VSmkZu
0C5IxpHa/9EAXZsSR+cemL2Xna+rpcLV0LpM59ETjcpEUFQTp+ken8HCQ6K0
9bRJPTXL18gzTK61/VlwcpzquNQyeRi0TA0QXQo23tgiDPUrS7GsGT85KMAq
8wuuve+3yT8RHsXpb+GfFCPGy0FXkXnLI7D6a3U4oEMRVetDqhRzcfB4mUQn
VDiEUAtNvwkOenHsuWshojp0eQZ99i+/1FCzU3J29egB4Dnwia+TYnwHQ+A1
0FkcBVBufSze1girb1nQkTjRpocNansEi1t46yDGnSCBYKs4x1z0pg9FlzZp
K4CJUE8DPq1GVvEX7bvek6I3tK407giT/rLRJCh2UidKn2IiG3QH4brwyf5x
1vwIFBXFSv/TiDaAdjO2QRB+Bc6RxTtWBlQOrTPYWXVx7G74ERplUTaJlv/V
+f6s3IwTA2I220Idaauci/Eq6wrsXHdRkd7uxbqpXQhUVp5gRf+YaD2iSBOy
p5XICE32Y1kW2R1kWK8PP3z+Zv5sHGd9CF216sBcCuRNLBePq6uc8qDvri9z
gBmaZHVy6sAJrCbd7YTgwatl3UcPPbzISPM0zh+RcFifegy71onqTUYWpCTN
rIiQq/wulOCJ+OiQB6PZb0pRTHXX7paxN58kH2cJ9mcJlk+ENcHvXnA7p8e8
q5yS64CvS3OmcBYNoMT8Ti8WbS/ttUcrOSYoAGF3tiYDsWam0+j+Liq5VQFL
aSMgK/GyAffzAAJdTIzDGx4pXwuvRo3GEVGmJq7KJeGkq1/O0xf8FJ3a09hI
OEBvxhZKsE7qt6z1H0bR2QzoHB0P6t7/L+Y3BhvECurMZoou/OyNl6px0PbB
zNNK2/BAEDFu5kcq6ifI6kSj9FXZbNjz8mLkMkz+iQLBbbFiyCIGBozW+HDw
y9BeyaCXaYtqQliUDkqGKhAExCh9link0bIo+6Hj7qGvXYH1UDSQUCnFgm1B
corjmYhzWvTjHH60PuBhw/SrmjaZHPYvK/EUTqGEhiTt0iUzIUcEiBhB4P89
EmAv4LfZi+FMAjINlHq4CsW2j6E5VVpOWCEYh1aNGkw8a9vBvxAWQ1IMTgTl
FujP2Vyd18+4TngXMpraQZUs+ix4+8ZSFlXg9OJsl2MMie8WzxcZ2/TSJ5pD
4LAUh+eSsXT0i/HGSooiXDQtqgaSkSNMxhRECIEuKAFHYPR0+gEXBZ+IHU5J
wZL5J5aS2GsddrmJfQxjwpufnZB0C4cox3YGcmNd3E85Lc92f8h4asVZyqOb
ptFZVEd44V/H/NkUkRrx0dnO5aqmM2zhM+tUA+PGRHZzKNavSHEBFRhqCdNF
7n8k97zPxnCZXFozu0PyPibRKpeD0FWEJFSbR4qBcadxkAbRJKo2PrVifKUB
5uoTayltxCrPOrZ0U8acQu3AJyYct0ee5gMBcaK+x4wYYTIxOUnPk03sqr4M
Ocj8mEsXTEa1m1SU+wUXquHYdg1f1WkiZskkui5tQ3k26nqKRB5limXy2E1S
qlb4WjbbjvbZYtCbA6AYDheSglH4ZtiiaYLZuDwI7cS/AJyo66ndIOUuampt
+Y8bwOX8cuf+0ESXOPOL1FeeA2Le/9xvh8W2Z2401uxvxLHu92BAADVUuaR+
no651AgHDtnIihOgS84QfqS8f52vOQejYkCO1j8W3dnWbiGpZq0ktciwwX7G
0jeHJGMRUvIVb5thVp5kQT+q03+AUxBR1/5k/gLUEHeylcLmiWFoj8buAg3A
aXTK0hT33vC8iFb1HBNJC+3NZmCcVyhqwGC8MR4W0Cqjb376eb432paS/VTG
K67NjmnD/s3CbzV+li7LrW2b75KIpctmGPgeWAuF//DvE/CjpnO5hjkbCnsq
GsnzYGTGzWQ984lauvixZEcmnc8gK8k/iCsGCLgz2yudgA1sjMM/bimNRUve
Hdi0mnybwPdsmLoP2ajb3/B+oAZYdAMMDQTl5YNYyyItChJ9ZR9JA09jyD1R
7AhB+NT1TtlddBnIRIRsD31AOXvb1AEynFdENk4dxdtce0cUcXFuM+rkHyAB
noDwUTZ/ciJIfG3XqfJxf/YI9mNp37WPTZ1vsW3TGbfQWcFalUu5ka03PW00
cQ3aMWasmAlEJNBCcIE7Cm/35ErgYrwQts3i0in6d073xVAKqlCDYvdFcu/9
AVDnNC1KT7cLPGexBMFW4Thhd0Zyk7N4fg++wNx7nW2snlgjYraiTA9BRutg
vF+j7j74nlcPJW+03ld+1FZCb6lDMvnsKTG2LAoTUNS3eL/fvPZBMQuyF5tX
rKPJLLT8DZ76DiAgmg1HvN2A80R+R+7tVfUVCJsmeW/N2gOzLF6z7egdaM5G
IsdL919kzWCaXiR3c7wRiYq9KBK8tQVZZaITLtJfgSZyK53Ok44IfF8OkN60
9u8NzPuZ3rLI5ctwmzjUN7C60I9HWfa8EdLpeWT76Hg+OQMM4UOFiXMmDrLZ
QTnSqozHFw0TK+ER8MluDOlZJI8z/ncPuYJGxApseb3to9UjVR+lBO5uP63L
ajqfb7n88j8LVwPjEEZghftaVpJ0n3lf0DmarRGJAQKOO5pDgMnhIoX+qoBR
HuC+EGJiDlK/ml1S4DWMcseyeclvzSLVy2ARN/MTuWxlNTg7L7BJrFZsRSl+
NcLgHOMBNDFudcpVKvmZEdNA96OARCR6FMhxa2AWs3pbgXJteyAG1qIxv1Ur
dWIJNim8rc0EM4b8lr2eFcfMhgzOMIYKN+dyLamqC5tCKDK/caCiHS9eMh4h
t8YRw+vQw19dUVGD1n1SMWWL9hxvvKO6WzwRe+feY/PMmJXM99JFd+e2v4k+
I2pe/v1ebct3F+jf4zYKAXM/k5kQbViG2BWg/C3hPfQ69RB7ZOQlfaLZOgeN
CmCFwPKm+MQ3UfsoYDKVIjpKLfxC27Q2As1Xhgnrp5lqmYOkuisEx4toEISo
ScvVyqBTS+lla5cLihoOhlWuXBZ+zFPVd+lw0hKJ7NJhVCVkTndTn9ygVUlg
+WniU4eOpvJ4o+bh+KWvluyNE5gH39ZNzMhBrdM0tNmSWDPBBEn93TnSt5VD
E3yi+Sdvc2vikSxXjA1BOOHv+U/Ck0IwF5jQ24UNrXuydyKCK4PRoE7OKN/z
chnGiXGAQXDXV0e8488GkbssiEdGTzCrkWklwvDnShqJsb7ivME35Lp5pjwE
6Xl9RMqyefhQhCLBAvDVVhOAFmCcLuonvxtFLmBQnW9D24BxJSjAQGuBZjj5
BrXz5vt4jW3w6jMsKI9ccj7lWs8OXXmK42FWkEFEM7ipWtAVeQRIBKOTP+hV
biOeUNq0h4T48v1QCs+AL4B60o+GAgH0JnY6aeG7s92xW12g+dnqQwgNPUrQ
Q+91OP99AMggkdhk70smiQujyxGQM4Q/+/KNq6+No1BqoUuKPN7UU4a2+bDI
nurlctTSQ6bd1yVSBJjpKCagzOh6S18PPG5rLKMMfylB213vBmwYN1Ojtmhz
JYETvA6H+Ze/Cr1UuxRBe0Vb5bbh7yh4MpnO220xE+qP9LI3Z5JFiWT4Tqsm
14LNiHhybrfYLmARhEiqX3qPUmuE3J9kcEfl69sZfYIsBPdM+REczIZl+RzO
BDNm5lf5JZ749WZMxYmY1D+R4Crw1pKe8ys+z3QTPUHm8zq5aUCntjYLTUeR
zFqiGq+qsrf19mgH0wuS0dUA86gL2fi1gLodmcvoXr5F0Za+dJSNs3etzzbr
yWjfsc4xC4fzlcGMqF+6DGKMdp2V1Mu2l8Ht6qfRsRLFWhgvQAsXEVtWd/Y7
UhspOz5gCcUqcYI9gqeU15cftfi7xpyrTE0brtj26ygo/LDMZElR7Lb6yCcm
Jf9+Tzmb8UgLYV7MwRseOqdaXp3garRkLuom9MD4sfEXcFAERBGNKiJrH2Vc
W24/6wDDNlVg/Fh/t4xpNtE8PxaDjfIgOYzER9Ml/rgSUXTvYpa/GZjnm2XI
lphQvlNkc85pWdewr81bkI1EeLcPfsKjrlpJUcKspKMVj74Z0zfM7ruP4A5S
H76oxQ7jhq2/oS4NRGN+AzADW8sjqe5f90W49pkiYx/bT1O6nirV9u/cMk/4
I5XD8RSvisldy3RmtEt2P2z+ZRXn2ubDGNlVcLHGUpJlg/+QcDxn0yAgygN4
BaJCdmwyYyi3wzcwdQIHiImPDk83uzVPIyermXd/BryZ8FzAvo75B0Q7najC
EKq7y6e5vU/zAzBA58UbsnAnvuwIYnjyv8oyoRUew7uw1XMLaM7t4/4krXLD
hosqWt8nGuLmcIdHtLctbZZHDypW8hMJxEXqEnpvXlzbqKV4kQyVPOc8Z5mp
t0y5SdElqJmpoj18el9H4FEvrurlBKxs/jZl7edyay0O71A0Q4y6xpEKiENq
nJLV6CyiO8VOopYG3WVJyif6riYUV7ylZTYy8VUD+SHNttUdddSpI+KujnTB
yWfQ3wzdoNAmwC9uE5dvGqq0BWgaKX1iWshNRfyj5Mt1MN6MzzO+FOB7nYWE
xEZXSkMfNlW7IWciGigWhp7V3DeA3T6wyaxbZn6VrczAGS5Pgls54IuxMOjm
96wmXmnYa7Y2hxY1KusOzFPYhfNM/D/Oow0QWNHlEjIKq0n6Tn8t0/ZSejIS
dqowAnq2HVr09kJTJ5RqUr6tb78jRrPL/lxVxxgwHMBdT/e9xjbwlb+fIRsR
dwIHVd+ZHsvFpgXUvT1Zvnmjh+mnVFJ84k21z5lsDa/PhogNTVb9g0rR8gv2
khpy6lPG96gQjxUHpDMojeF7/rfMd4SNaAWvT0dsLabsPKHbrhllr85trtLk
wjfl51OqH9Ndc2tPe0yV56MS/meI1mfTfr+ueNBUbssjt0yUOM3o3swvMOBQ
LbzE1+jLJFP8B2uw+2B+UvUwqRbz4bO/cxfnZe6HMCV6UKiKWQxR/lhoiW/s
i72MW0zG1XRlIVCh3yZrByaSAYGlg0Tog+EccdYyC12Y3NCO+WiEpNRqn2BG
uocDR7vMzufnRNUGgVStW6eUrY7OljXtk2uex9u4fb2/p0U5OOFYHN4KOGpD
1fSIj+NdTalap20kvDf/YFmMTnhKjCbTBgLumPmPVy/Q1HyYQWlNiXr1N8oL
9nz8xUCH1PFamN5OAJmIQE1t9ntxrXD0B8m2yvJB7Sccac0jAjJmg+4FDnYk
Vap1Gu8z9P4Qab1A8AP5qmCFQOSmUvSF2Q+e/VGDjAVAbGY7f8t6Szm56ftx
MAsYX8x2jmJe4l2r2QahCXj5BA6pFSICa59/U01GlxHpQkmDGFWduEHXFZcP
jB9LVMPoeKioN8prI6wt0YeNJJPRYxxtAx9lhN4+UjV5geMCT/1c51jU5Hcu
uOQVxyKxzlzfvlx4+0XGY2V7oSFVPlv8dQWYFFvcieqKIzLWCIcK8uKlmK7d
rLF98BlLeLrTqK2viR/rL0X4Ih3konVczMeC6nMLAoYgTy764AIzF57ZP0b2
L67X3ModuaoA8m21Ti2jOGPok67eFvJ6dzD16jRI6r+VqhWXIfMYnBbQDlqI
AgmFvpAJ/4f/iT1zm2Baacvu1yGo0FFKXhWYGxvVpwcRMmSp/7UvTJHr0S4V
+X34CUzHywEyHciEK6jVSVMucPX/Slr7plxb6UsugmQaOWUHm8rtUIcd70BM
G1z/QC2n17Tk7Bx898ZTSB0nLjpbQ8HYL5+UQSdKf0+mF7xm+O5auIO/RjdY
JG378wq9Jug2+IxNQeUlVAloxIT4NV61Vaj4ZZWRODz1wdUrUBV06MVYwRcI
KILN5hKNoZcuA0YlzkhBII5WeSKigfHa/Il9mGESPMrFu1KXtE7dHaLqbhEW
PAloL6FyqjTObQd5fPjPfUjOLiiWUeeBkWhU0bFm+tInI8xrJTV04tyWsLZw
hIjjgOw4eAyCQ7qZi+5x0iAtJSDCAM9JgsR4/aO4XtxZ5QJgywSO15nGlRQn
0XOiVEFANUO7V1Gek82VjslNsD6Yoj7GS5TQWfBi8/Wo1kIsYkPzv9/fRmz6
BMHSkYt2cfE+QfrwwgDp0mYmVHUy+/N9XPAMetHYL6M2kTbEKpprFY2kL2Gt
IhkzBsi1V/fksVYV5vbZzFdz3YCtx0xgEh1ZpM1+jbMcpLoVzMrjZHqGAQ3s
5/zpDJ5To2q6SM5zWTTbr68G/emdvVZ+4DTCZaA0hpjpUFo92Zc8Ybv+lFFI
GvalbD4V25y6MLcQzVXADuxRhMa6DOsl0BrtERabttHCq/K14wV7miF6cKrt
jCBsDzUHhRNleb96JNiQ/XqfKSgWSRkp4tIaHC7aYB/g+dagt+nzUcBnCZlt
Jx68YFSk5p3XiomuXYvt4BEc06t88DoANr1s1S2U8RVlIAMst9VXGEhX//Ip
FD57SmaanErhXFHPrM6pzq5UCA3UO/YHW8ciA1abhKDSUvItMYrERP8D6jSZ
ZUmM7qDZvHM8WLMVd8QzA1y29T1+G4LYkzcRvz54NYTJje7SUAxXvrzkb2Mx
5xQLzcDQkwTjvkDkHm3PCYze8lKn6d/pv7SQB8P7sMKL99g5QRxKhc54408Y
5nEOVwIIlTj8wxklLf42zXkxKc06BdhjVPN5mgQEh6o9b2XDftUJhdo3wrDm
TUZQAi+oFGsSqM5xEtM0UxTLKyUKTeT8oVvJmYW/gdMclJ+QZiE4ynFkhT0j
cPUi77AhpAFqDUZFTxDGUkpkpgCzC71eAbR7d/WFrUETfMAW5+pn8XdsGicC
yyDpIkOlWJMaSwmwicL5anBXFIFZvQFE/YkVYmME4Aq3vNH2m2HnrXneD6bL
h3vGf1FBqHadFuPEAU/YMAccVsG2rVzTc9hCXp9N0+ze16OhjLtyo/jkWv40
PMmiytSW/9KYolTj9ESHBOyCSO62Dase+S32SSsKiyGfL/x7aQV9nRBI4vEY
SOVbyaqESOavlUJwiBNayrtlz0i53VFSWHxMeKgXA6F7sBeKbHvlyPJfJCjD
V/+7uWjVcZA9BAcEqaZM+R1ymmjUFyoQxjF7KsN7/Wgk3UJ1hvSXKH4KBCzM
GKIDGqlINRBPxnO7L2rZ1o5HpUWf58yx3cGtmlzc2HfXz1R2k0OFRu/XJcQL
21MgcgvmZ58+a3DEdJjNUr3D8qrbOn1DlSqbtTOC/e+9PWtag5LkiqusswZA
+0IfcJHHFfsYr03cKB51xb4C2ejFLp8OKOzAJjCqIsky6HkZ2G54EafrlSCf
gGVsmq+NaYmsUA+vxFaHtzCSWUL0zZw7ZLyZsrFuBoKZm6oGFocNpwPt0hYa
NTnJLz3G3lL2uhO6AXfLQ2nPdp8QFuacg1nT/4O1mxOhv030y2IkPsOdPdSt
z7G5cKJeXmd2P8Oi/8aqrn7I9jSMF6Z6NRlvDAOtVi/ka60lwCdXoAre9g8M
a0O+pBrmkbmeFQEvu9sO0FILfrPoRcyl6hO/IkHmG+m75j6yDioGSPa2YJaC
hQbRxz7lndGbgSouj3RPUc8302WZe000sXO4rsj9MaWnUjkvNJHXd6cOtMax
diKh5iwALfRmyg+/kS76N0j6OZ1Hbfv3wSTSzwMrqPuuTuwusGdzWh0wjhS4
7TPoNuhjnGXmMfMm+PW600bU06dzG21euutae1w6nxtgXHh7QgrhjwBXh8lq
1RRKkq0XVcKhAABTz/IbggvMtXEnY1sqZIlhV85vLF+wydoaOmkSfFyXXvPX
LCr3MHk+Y3txY1jxlOAzV2PzJAgSLbGcvNc7lbjfKC6HOyD9g9aVwdmK4lv/
eZXuB+PmixDmyAoPTnlw3ZQ2TdXm+0x3iFzQgIIUH9a92t2J2QYBA42ZkISC
havFtyVWCWUA7YSihoVCOahqWeXnAUd8kQne5GUqryeMWi6zKq5336JUrVds
fkLwdNNJmlq4PTRPoBhU2pFyQRmRIIHX+ZdPJPxCrIL80SeUC+mkAyEmJLlU
gZ/grVmTJN4Ti0J6aR/2pLhsrunJPOeey0nMnfZZ4j3Sh1FilVht1lWgqHNL
PUW88rheRcblp0vltIfO9uw8ADJz2iWZWdBOWq9fCZ+UQWhPQVlUIuYyCDlT
su/qumH6RVyoqabFZJhIq1MheGaT5+9QvKhzx4zPfL0amGm5AkPuCi1NgGkL
9bbfqOjTMXl6utn7saBPF9T8xhH0O8sPYeW3YPRfJdqAlYpv5P1uVlD2/wxb
JJiSPCtZskhUZ3nnSSrtFIb0pUMF/UsalKR/cOC0uA41LxpHmoBI+Z8aZs/q
rE/2QmqZo7OCMBUkNq3m7IrwhZ9r++huX3vs6hOLFNmf8RhQTheivC+2E/Rw
Jas3qJqmQcvPhFLM575eX5ahFIlOzprECvcanWAybEEsp+Q6Qfqw7Qnn78bv
UiplJ67vFYW64r12zokuYultzfuSBTYmMN/6v4r7Q7wUUwcXLrc2AXzl7EbM
rumCbqJJygHMN9mWlMXfItvgk80aAHQdHBj0KciCzt/7vgg66qaWMc996Lfh
5QAcIO5NGw9vrtZ+CZEuCq5j4NBz5XbOQ9TictjsETViamS7eveo7doXb5JN
ylMxXv1F1ZDmPP09oNVwyoEp+k7gOII6nJEkE8Lzp7vNN+YLaUba0zLmdteF
UMOljxIXfSwc2thcuXwBf6ATg6XK3u4g6vIu4mx2tZ1aFcri8ap2LJwY2ni/
nJ1KseRch6FbYkW2bSXYO4SIGQXQZBDnEWZaBLg4X9IrU7XPRvrf+W55XvMq
vFTg+iIqYTVrJIHGzl9uIRHuqX5j4FH0kVBwSavH1PO5bqYBidiN+57WtJhW
HLZGPyneBe63iN9iGYh4yTeCTV1zZpxfd9Y/jVAI9NyY/TFjE/TMqH1Ji2zT
dad4+L8oMYzb5ADufcPkSrz0YEaaTwk2wwe6BDiWeyPfhr8Jy9U5El1z3OOX
avi64pO/tzEGXw3IV1iDJRigI7zDQWvm6GTd9S9I96l3GQmYuctjhin554UI
z4PYiXZRSd3KopiLwJqlYqDeIt/8mAYakePueKZsGdsngdV6OCt27BGx0HtR
gVpvb4r9PoIuq3IxBPfyZjmH2yX159AildWqDzG5YSOY88A0DLgGgQQZjvMs
1LZBOeCTJcvkXMfSKQ3gZoKFBvDADyN8lWLyArnuTutrRWbxAdHPLdCm/qrl
+6oCkGOSuJJuZd+8vxMOoTowxBEBe2nihYfiXRrSFDm/ZrReOHBqlWfFiFlb
osGEg8ubjD9WAmUP9F+EJe3SkkvekF490qzw515Pg262WOKxQO8joe1hEGxd
P0OTW1cOt44KGbbGPnCi9DJnYczgYzcsKxoGVgv1c9dcEuoz29A/6LlI/mXO
+NpPWd0KCgIgm8aNoj2MHbI/XLVlRo1Liq4kRpMLY+MeqUJk6caj7G/tYtzI
ahBL0jaoTS+Dlr6FKpAGjHLguqrgMmYI8hg231ZluhySPN42ukgrtYuR0U/3
+gVOcDMt8/fy4WiInwlX+E2IzAtq1jLl4C31dSGLIerOdGv36YrtnxhRyTzo
scmw+miiolPtfPaefMHHwffkkT6I7wd/cg7mbrCEU5ExVSi6EHwa5VpKbCK8
kKyI8GPyD61cDn4O5tHoBtQu/ILwoOeVQj7AEHSbMU1lkcSRvpqMx09etVCK
sR9c2Y3gw3K4EpgK6E0tnWntRYVgmJ7AzKEmzhySOaT/Xb0ShVcYykOxJpOa
Kl+nhUiWg82HGtek7DYNRbhnsja+ZEVPI49bQA6JSW7Vz6v2fzW8QeSw7xPl
lF9/fB9tJCW7XrS2lK77B+fN7zyc9wZgSme+Kc2HByt5PNk9OLSqay864dxI
k6kHNIV71riSAq+jRJpgbBbe8ARGZIFdZwsL/x62a33U01IKsgxI69126zz/
mRX1P2UJo++/HufgzqUbL0WXGEEXQ5/rQB3o+wEVqDqptLRKyiDM7WZCZBLy
Abq0RJEp/D4d3VOIcbhzn3wkWrUB4hqkmAZRNQAzuWC2D6mRY3riPfUfCsIm
ZfCR+Xei/pUJRIzB4TeSUpzXWZ8lwv0+lSMRFchRo0Pmzg6U5xWX9S23Mohf
E2ROoHAoU+LFnpW0aX2DwqfpnMYXXMHgCK5X5vHCB/8Sl/1QjS9A7NDOxTBh
CDt9z1D/pHsJwTSJZkk3Ie3z1rx9IA3cUmg4tLiwkcxA/vTcFxfExGZ8ZmtD
E+wDVqsoVozyT+Bk9AykisKNlrdhZk49lQ+ghdguE6LKrzmxSlHJGimBqq8s
8OLhxQxV/aMSojnNfyEPrH2TlU9qJ00uMLVAAuXw2vcuv+sAR/UQerI2xGf1
GwBIA51bLhELqq2U6+OnbxHJNe18nOCO4ZZdiyEmaTg3hUxYJIJhbMDxgHAE
Jbyj/DRAge5xx+taxZUrh9oheBzSEYghBaBKHv/nO2wjpt/10il9xLVrWdUE
pCAH3YZ9f+QtDtpdOJQsGhGawT26OvPRwOhw6qnFA4Czh2SGSjCgUxm15Ret
ITHwNyDtX86J8lzJWVw0H1gP0C5Ha2e6QExm+OPA4BtZbwZ2i06Ksdnpwake
BfWppvBs8Sg35S3ImjoRB1iii3Y42mRP/pSxxJx3Bshzht56wKYJVJM8kSD9
doTeXfeEdNo8bpTOlZzi5pG/bbnaNQK2o9gLh7X/MLf0Ev1yLQRWg/RxqITp
zE2DgaPVYYuMzADVGi7YLU2ouhRQHRtL4ErwL6zrGNAyYghvTbvVzgH8mjg6
JPJzr56ACAFgErxCDVOJsVFUxpQYdfLTPtYCYB0PNs6Sunbm2qA2MgNzBQ4B
2VCwDtzp2hWyxvr9JSoixECGOchS+xueIBkqRGfMeUVcn94c6fFiWB7Q28sw
N4ShbTGzSejIMWczL6OIxiWwcdMYZuTYzKWfbnWp5k7WimIc/HhNTvmT6jIn
RkKZlo8wijR/sDT1QXqMjos0nhTt0HG9NqWx0KWiHy0ofueBdLeYoRDftyFr
n3rHtMLcHuNdU9OND1o1WgQ9GN8iK3lXsYgDASM7DrdwXpofSw06q6SZ5lXv
c4bKwu6eFB06a+ME9huzIEyg3n9YJzZwEgRWKxs3PrxWGvSluBm+CtnF2nZ7
cMM+jbKs3os8BhZHN0E09aD1n0IWkaR6Y0FBaahmSWZ+yWVYuUJWfu3/T5P5
P9uui8wH0wAn5qG6FYEN57v+GW1REV0HtmyUEC1pxi5CcZeP3fCgYrsocUXK
2Iy+DvB0iBLOZxydE/EYmHYRwc7iYpbUgP+QmWVTF6Lj9sghqjbC4mzvTYEe
gOeE+06UR2gM7jOxTNrz0OONuirHPTr4GCeGqEnPShHON94zEm+QZrHLaiUv
vX/0zA/y7zh160TRGZW2vYmdwiJO59Clw91473ptsDBd2j2apTgEAuVNNYnH
dpRgyKnqOE2yqiOA4y9gwOjQuPGrPPo6pD8tu+JAeMO4beT6vuGZ2Gb/D5lm
uUZM6kW6D1YP0g6FzkYvKD0Df+5ARwXEbbEP8BzjoBo+U+ZSpducxQkod7il
Z7wDOrlhTBt0Uqw0SUFWxudGZ24CzzfpaEL6m+7r/6cWlNCnRTJz9F3S3+LS
T4J8WB/3X1mc2Bzx7oqomfImx5Bdd6xPrRJ5uRfwBPT9dpbSDgZNv0/zBKCb
LPdBDS+H7CqJuYQbjshztQDCee9t9NeuMkRvUZG497f/i3mgzZ4MiOchPFR8
ECKnw4fvuvqvoMdUkylF31s/aM1zIb6GbYZ55tfZajv0fLi7KwCaTv3Tzv7j
7nC1zNtFNmZWIAl3TP1X5jm2kNw1Xyu35orQnhZPHP8vY6M6+us/rImWqsOG
QV/jHMh3EubVJ+AwiXg9p6xHUWB2a+6YCgv4nmGQMbePjDwKdGZnxRWkbioG
XXd9VnzB47ks4qOzDSTIWJKpmgJfDEfDmK2snI+O+yq8R1slRVwqqbKBq6tW
KwvN+ICElD8wRMJIdNWyR/mtnykVFuYlxdiGSzKZn85TFx/s4fEwp/RnIFXp
41Y1LUhNzblNGiktc5ZkQ54IczitShnssMXFsnIm+WmpfypJts/Y1LyhW5BS
eGfT566Cfv+dbQtJVfFF+zK+ZMD1uQePTCob18o/02YT16tpVvW58HW0epE9
kzV3ozl09RsySyQ74Cz/lpZ4aGYGrv70UKkDgnWkXrE++8XOSyOBsvshh3Xo
/ua9o6de3KEtP6/W76nmrQLF2U/jfmKsr8cFIPOov5y4+iOsrNu8NZf5FCIp
A+M+n6IcUJYhmc5G0DEDY+dPKL/aG2vWtpk78IFgo4gNDL+dfJSFxN4Lf6tO
jJMjdqyBUU8xal+cGomdis21toh2VLyeK+t8PNSv+95fkSxsvXYSNqJ0/eY5
hmlxId1Qapzwy93hgGqoqXbAJmy9q8GgyykCdXgaIBqFctzDb2VVCwxZM6+y
/a3DRZcEnd+5hv8UsA4LTvOBM365K9U6wizzxKRmygU+jklsVyCKPljvTk9C
G7CHT+xfqhhrgYbIi0rsZqoC4OS6/zbOusJ8u4e9BGC6sJyS9PNdVWp6/7wX
mKKkqaXooiKRfaRBdsSw5cnsHJyVliIvhWSvc15VqYi7UDvPgGlEcYI3/iPT
lq1pF6L9vuAsgZlWXxs/hcM/JEMc8pI78DpZc8aZYeCFPUIVfxdYfnj93mmU
9cJUPaWEO8nqT+rnITPiMah+AbPlLOVp8WjFKE19+P8tUGFhmc1ylM62A5LK
pX3FHNoc3N6RG4PviObqGVTue2m39cgHLU4yuchURiMbxmIJQLeEIH04lbaB
5XucczcwY8lsPw7jPPHeUhp8T+YXKfpMhw0IuClXzHifyZu9rleawZLAWe9W
EfisLGz5bRgSGbQ7KafNioVDX7LCeVkmsS/TbPtOaU5pZyrwVdowEvgEDyQE
8lSONa3evvM1bE8SN3O08wDxjv++hIZp34bCpcAlRU6wkjJfwqoIqUmW44/i
DsAzlbP/nBWznZh9eM4E6ETltoZcqJ1JY0+ITcivCE74t/f/hVgC6rePvyK+
JNnYtRyt7J6BfwBzPPeTbjI4qfY4clCxZIbwJQ+DNR+JMHnRID9fCIR0i8e6
47J9vP7fi3eIYc16DQJUXMjoBN3VZN9vHRN6qs7bJ7Ql9AXXj6GtOYx8FuLY
H9eDyiiwXfVk9zYJ727yJUWZ9gmr4Yk2IB/tRQmpsDtoQMBJih+56IKdBIjd
odrMP6rKqaQlvchTKZt/tNeKGRii+JP4nOw9HH9p4Se/HzoT3nVPMCKRRkSv
30Wsgcm6jBWVI/afPWiy0mWQLiwOTARUenmDVxLgZc2iRWRN4O9b5V0Xs2MO
qVDvPUKJoMeYQE6hn6gZ+TIP6Iuw1CS1UambJR7N8dTaJAX5iM5Gu2GIOLNT
XER+unfWnbfI5HTPVIPOpsEf39NIa6KldAHWGSGnyfP9KRcljzcL+Z+72K4Y
b1b5w9dXEsX1355FCHje7GcVvYPG0SWNnz8aYYh7Mtcq21n/41shZ1h+Lx2v
i8n5tZtI9qFy4GyUdyuDj6H5M5aV5LT2sg7Wys2egCNGAFZpGklRQ+wfWnFm
vh89Y732wWGf6yItdNX/+idwJr/kvA9GYOi4K1XF06UgW5vKY4l/wwXxIs7m
bVGFOszhEo2HsBUNHyUR1mwD1fdmvVo04oH21UXA7VQIX86z9tsdveNhnXOv
cpVgOzzRhmW+vEKLrL1mX+LtI33FncnnQIgumZMo0k6pETtDMy5whqJUawT3
V3ozSUlzvR/MX1BTwXWTO22RonlEyWLjRsMjVJ1imcqhDvZA4Wm1JO9l0gLC
aBq2bmtNYmp1kTyVLXFZR7B0gKQ+hLcLsdNwMLgG6DplYu3mpirlsXNbyvC0
PUFWtbIOJrjSMCanGos8cUFB+DA27I7wEVT78LP6hfkVQhJC50Koqn5vHxO+
mJQ+2lLMM9gsvl9jBumNyvGqYubcHGW90Cccne0mVhfkSU4YtErm1EtWkTJY
YexBUn7dh9yOoAWJG7afeFuujU1vomvnxVeSLu0besDhTzCQ3ubhuqfeKUKD
a6n5IlsLRv5SlhWkUjFg3nDeelf9Fle2XLkUu4Q5Nj0FBqMsOCAaUHElfBF7
4O3Y2YdYQtJQxibwILTlkNLKCfMibwqBC1wFR9rTJWYldnbfntNWKTo2A/gv
FCdkS/0CNQBLzuVSYMs5Vgj5OP7oPPHqH4XAnR0QS2T9ZTNOYuUUPCcTv3hi
cYXtDkfjWmJ3qQxEffL6vEoFUpQ3IU6NZBPk4clta/mCrvTIi3muoc/VNn3i
eeu2Bd+0xOYpaGa2JxXUAxFEm2z4sk0bl+mItHw3HYmTrE14fDEAzt9PeeJ0
ega6rK7UlTNit5oOyUdBQ5tAj31JlqDE4naySUdSoGp6+Y/5LbfO8v9D97yD
NFwyjdU8kLDCyrS1YyiFuYYGXazrbKlR/c2Pk4zPRHEzvyB/YHVvGgOnpQ/O
/YVwTe8G9ygdBnrczF0Vflq4fyZoQsdFn7Lc7wZ6EkbP25g1xvPm2KKcEYxW
ghelFjeIxrsBEN2UMRc9J0JWHprd4kbUAarFB3Kli9c69/ZWd6q+ko2AkWmZ
4P+MfsfN2x2aosPXFuhsxT4z+i95IXIssA0y2Wdv/9dxBaTdAZjdyp4cEmT/
ulFEGt6sBbtWCXCv4etbFntqtj1fT4eGHi8SWsT6gXf/ZaZOZXfSSajECrz/
kNsaRBmqaYJVogcuEtZbrPn69zMmSoUgVpQJmf/bRIDkhB2BCKudSVvLAFTO
BlIwiF/CIsKRjUS3CXkK1colCzqx/5JcBdGGyyCidQQNfYRfiRUBE0O0Lfjf
iRroCWjBvV/NLh0uO8aMF8Lx+cj2p3k7q+ILfwhK5WL5OZCn3lAVnOr7RMyX
C+2dFqqvzbzz5KdFvLQwIsiupf/1OnhuXcm0gyWoUfz7osyqvrO1Yc9MotvG
XaIRkcapuEPZG7F6AN2YIXGj57yCJfRtqK7lXYj3oaetKwuuFkCU45qfdaFc
RkBtEOYG7B2Ynkb3yQUy8b7c7VHh3rFd1yEnHng6MDXk+hQRO06SqDbBo2II
wmLPgWE6DyP8P4z32DXtSJsnDSohHyHtR9DlVEfxQjMk/f28cNrx1X5rw/mp
WGmP2dCh0eo2v8QBRtbu2yXwwq7EvINZnqDmawY9CTrWDtin247hxAX0aKiW
vfY6FpPiMz2Q76Eg14rGcn6bs9oBJ9p8QQZzPxPdcEefsp06JbUXytQddfeG
+CHQm30HoLwahjSZaKOqlzNkuo4iBj3t3HTkpGyc1rW5r7xoukL0NODORsrV
arazG1/NODoW2EeP36rwWl+OMhglC0oAkdieaA/ShwXOWzwk15WLPdLLiZSo
S1Li2PIY2UsKETczet6sPcSoF3jAz4IO2bHWF7eecUJxlphNJBOq/8RNgh+T
PLQYenIV0QrGHnihc9dYy+6kTBczb6Tgty4prPJUk3Fhekbp6AUnlFgdqKG5
rAeNxlW+m3B5VNLB6e/dJtITzWUldsgtu1XDmwd9QfCdIIbIgFThf/NjWDI/
W5nRwQs1rDv2MRQTSffQGLcQVL0OgZEJeaQI2pLaqYNLktaslVBu4lLn3+o/
ISqyTyMPwSWsY7qewX/k0jY59QrU2oY314x0KmhZG0sX70WXS1oAK2x1R3sv
6t/A4WWBlmaA8siN/B8y7RT2Vr9+4j/smcKzzR9LbGkfjjR2Ev9mOgU66m3O
HIV1rK3IcVLZapegOL+2GkCMHcQaYPipJ3I3rM3JHFZLTq7elytYMJuhi3Lg
Y4uwHkHpxMSz7HEfs+WbAPuE93o93jJFkjEyJ2Jn7NeJY2FdTJ+aiFQ+ryiZ
J2MerKHvhe2bACJqiGgNbS2/KNYRLFRIEneMeBD0ungTbXKK4KgQ5iw2x6wC
4QDp5DdqVGDS5JQpoA6mafam0gcEesUlaf/ubtIpsDxxEPa/aAOyfeffrNGE
/b1pbWTBfoiBW3hAFq5L7MqT71S4fi2WY3LBsCbKVfLNmusc8A1K+AdOlGzm
PBC02NbRDMeT2D0r39BmlIv/pR8O5Q+hb5PMWaTyhhp+4jLLG+I+EtjlByJM
JXh6xsO7IF+y+KK5XYWC+l3klYJeaoeh6GpMHVAMEE+BdRxIZzmwoitNZcFn
VU0KLgPIYqKLryptYOlLZ3SuOT3CZKUeBPE89ijVmN8fNJVpZ13OGRBMAiKf
6zbb2tmiyztEiv3W/6aq7tm1BfEAEKTuDV0ibXDprb6UffQVWF3Xdk8IsyCy
Tj8o0JkG1noFTn6ArhDyL2CHabTpNI2ytDB5FfBnBhENaIPaD+UNUzyXcXTO
Ht3F7RB0pELVisY33TB1kW8rdwpNI6MPgI0Hj+cqr/31F6TPatwbBi6fLC5F
7wWiZ2JxVLhzsQi9QZ4IEO7Tdf3XY2fEyq7e46qtbhme/lc2ZWnu+BBzS4Ck
RJTkbJLyNwQHjl6Ffd9J4+/ZsWmBNEJ4q+jjArjY1YekEkNabehvFW5H8Ti9
jl9quKAZrjSNXTglxLl/WOoy3lfUv9AwO7pYSMbMVmbsPi/nk1fPrr2MpC1L
bbDvAaIKZR57tCzKgXJzdqu50uJkXIo3M0bEfuOk4BP08RdvIvBtAKej10bx
acbBeh8LbDLdbPBwESs1fYA52cPeEi8axVQdTV6KauTp4/HCsYpKUyEIue1I
uOnOdKkilBasBEmuxFZg1d9t8uTipwl/tDjvUpaB6Ah9RuVqfM/JVg9T0ZWx
ce+9mn+PJ0ITAPrlC7QO/fyGj84NwKSRhVZaZpm5Pdmi/7J8nAUtneOCw/Vh
YGbUxC7xEYTyYzpld4OtI8NhBsKcnCNdr1W5yDhkEEVyA+h9uPVaaYaLUx3c
4yuFbLbh+zayvgHVkeUGOBgtxaI6yXzxciggEvT6tM6vvljupDmMpTJdSQir
7RZtEhQV9WiTmB9/PL9gGpfifVXuXC4CO3GCSKktS2Yt3YVdUQQCi/a/G0RX
uqjXhFgcgKKXGkxedPzrwoiX/HAGIGHkcHM/Wfy0pwHDLDqRgwz0oxxBs5qy
bWxK7tj2RYEnVtx0YWvIIsf2Jbxt5rJg0V7hwCL4wCHwy/c0mQ3V+0TyPkk/
FzjvWQmBCPEz5220i5VojyUGfa+zs/enyJV8Viq1mypwAo093woU6xDw518i
xRHMRpt5piiplu8nqIPh+q2Hm1V4uOgF8XMK7VXafKC0P4z/Tylp3HrvX7lz
NSDFGJVqEzi9Z4nPNDW7GU+1OaJ8ShOzqyAPjStg74nw+lQvOJpltMIlEBCk
T2sgyEcnJp0g6Ey8bpjjN1H4NfBJXU59rnT1mgGn5cW/WokC2AfM453JICPA
96hOWCzfU9vuz8vB98rayCR4sC8da5DRb7mwbUuoJiGA3nJ6bUwyPEksmduc
mZ0qaTUCjhhZ8PSTE3bQPlVbGed5aA0couqZhF3Nh1yvvaqQccnkF65bY02t
ijfOrZlY4arT8VrAUKWJJlO5vJCkZwEFqN+LyJoG7vhRaWi6s49Yi8qfpPQY
KBlpKG1zP4llUdrqXiLMXM6caEXR7HA0HVvSTy+UbJu6XjocHeAX1b1UAPJ7
Z3q2Qd6j5VKx2DTGPKWCzuZpx2uepHA9ZhgoZlQVi7YHkfS/bf4RTTb6UtsB
adQP6FZ4DzYLgJGd070dDtIwVSj6dt1HmnCicaWewvvXOfnWwOdZeZzF+MJd
G9jXH+oiEHPOeOUYQsx0gkvtaU7wBwcVzdVXP5Re3nscjQ+OI7RxsqFXRFRP
KZpPUKgVQSSumV++IlyE1aZ5YQAWjkXN+6of6rA1FTejuF2RLw8oNVvQQ20O
9dZzrA6uxEkpSrsIV2iI7EsbtM1OQOATZBynzqCVvJLtxN7iCJXh6jVq50oQ
t/+2p5d+MOY95FfgmZyThC4aUydjYtQ9aYTUlxUw7tMZ6CG5xTqvREoEb6s3
y4TQhVwDowCaRS9LmgbPO6mrXW9TxbeHQOwn86JQYBApwOVrvTdOcyoAOaL6
t/kOTUePlPFXcEsRgrjjy39U3vmiGawe1i5nf0LRO1/rNs7QRAoTC4J+ZFsX
lcrgHiTv2b6rcMlCFDWgGZ6CnMqC9b55DXxRakKCphh4RcoWt9yIVKjvyuBS
RVC6xZ73Ck1IvpsKix9b84Be2T6iivU/azrKeoaNR+sAb/KB4VPOleWblGPC
GhWE1Wm/OO76RnuFUqf5Ds0WVSRupWQYmsHHtTTYeUs09AYYQgS4cTTUMksw
genSBlXl+2qefljABvYlNUDzw47kIkPFyQHvIjf19bFxW+qVe9NCSWFg/CxR
X6aAzGQz7fIgZjRBiPIHO5DxmpzbBYco3MgI4v6ApAq1e+X/12mBDkkS/qpq
v8UuOVFQesyg7Li7aYZ99ymZSEJbAetRtC0NTD8TpNjVRCC0O/a49+cH3NL4
mix/qLWdcCA0HHWLRguJdekMAEJPoe936ugIjIMpi0uwGanKmHpmYuylA/NT
j7pfgpaifssryyrF/p/zdcelx7c470EJhsuJSz9g1FssNwpz0K/DQ+TcxCLI
rqEtcFoZGBP3g2XV9G2Vp+OGzK6ymjZCEmq/2OPveJfJ6eJoqe6YebgN9eTk
VT7iUYcPY75jOVAOxjgKtxto5YnYc8JGbanQWXHQtgi8XdcAusrOdfmfm7db
XYDHEZt4tBEmrM8vJrBNDudqsV3D0kz2Fb+bJMNtkNIBcyn1dSEAU+Z7T+T2
DVYUxK6CFf11dzF2ofd5L+Nx3VbSp6q1DvnftdfUMWcNbONKIURDoA5TiB1q
qkXoRbocgulwSlpI8+fcg1ExR0edElhsDnG6kt8/6O6ZYTQ02nkMWJt/sQHx
NbfnEyDhJeW0oDBlY6YofiYr38fQYHwtROuyENeIJg8KaTRUCztMiRAUNgRz
dVvaU1bzFOIAIwYxn/7pET5ux9RQ5nWImH8yybcYFzKpdPPp5+pUgpQIFmcn
v/h4pNReCdsReUCLdhNXOhXdkWytat0ermmtIAltWZsRDPVt7B06GL08Ms4z
N0zO6AXGrMT6GJF5z+LTZE8kOZo12pMLRss5NuiPLBeKzq7l+wk8Hyxw0zCv
H7xX2io2IYvFf1SDnVkqGNne3dLg8VgkWiY71zV1yV60kakd3il6KdrQA9hX
Kl8BwuM4mL5SrFtGWFTPPg7fgWFcCMISq/8DnJtfFXjaG6lyIBm1YuY6+n5K
9HQPqvjyEaUBDmICHXpFHS3Dstdgm042DgguwySBFkOp+ZbnwA3Jp59GBRvQ
qDTNCCgGnG96ARqYCvcM7kSp2WN6/pvqXX23DDOTWGCB2MAZjwZt/Cg+TU2w
wDjH1Cdr7zQ73yqCg5dzGBW4IJQbErCF5gQEDkh+vu7E4keQFun2SfRMII1i
X0FAj8W09acAvQK3SNCi8jiVMg7aVLjscrKcfCH03rLg/PmuUHKYLqMLaCjM
zYmDIZJXZhT09Y7HxZopp4qi3mdp+qzAK4RMf2mW2g/4MR6v4Y7MiGUjGLk7
XptGC5qOXiakXkhBCgxHaY6EFGa/tWGYiupmJOfVBwlmz6YQ1Btygu6QR1s6
Z6zxmodj7YuZQPhTdgAqkx7G8Z57oFw4e2MBNOhw1YQez127yZ2/GcLmLEev
jhdTv7tJ9Vh1uvWDCaCFVAb0N0J7Vb11vnFL6xAO5FjtZiiqCOgZ8J8VwEqC
1Qhw5PT9cQecW56NKw1otSyYHjVJ59vIHtiuHGhXZE3nrcNe2igGmhK99FOm
Caym1x8ulIvslRSsaGmaIdwgHidezioyid0E1mJeqS1oWjPQw0idMD2MRxJV
sigrw2iMkPyNpJ1gWRFCWpNPUv5BL1+80HPcXM9fYvrh4yqby4fYfCEVV1Ta
g9YAk02dd7vdNUvJW4nocKGl+eoSQ2zLBAr/UThT06XVCvrbT6MSnKyRGyDj
DdwV+g4Lys+1tW4Z0zbATY/6c9sbBUprtazZRZv2rJqncvgKa3yLHtPy6+Wv
QwN2gC4vyg7+UL+9r9HQruQ3WPCO5Zk6CZ5cLZcqQCSa5AR07v8uEZKD7GlY
mwKiNMqGiqOA/UGf8sDW0t7qDeSfM/eJZHQa2d3lDm64t+P/9pxTDMvgfmOj
jOWfXvxpw60ZjtVpfRcAuYuIM7oW7T277a34Zm6RtL1/ggnGdcmiTPb9Migz
V6PFINtSA+vGMgCLFEdPJE8KdYNx8ZMzn1q8EkU7CdiMwHZr0Jnd0etqcJmw
XWvhED+391N/IC6N7OGj04Y7sICOs8Y+GMNYdgoy+j4z+NgFLzMrwQ27aien
3Vc096hQcDusEq2AYP3bo+uhOXo+hYg/Zdl/llsDjnAyoPmpmUWM1tcXD/M5
59IvYgYqgnFjHHLWnMXxe+RDjh5dSmgqPvm4e9pQTJVL2MRWB18zxZkJSsms
swCCbQzySC3CfonbatS1gzqiI3txSU4mfIKRtQU3U4FM961htKbTsMvBOi6X
RgcDWVd9UqddWFzLnIruMIm0HSbCBZgwXKBsLSVhYLEhgGV7nSIdAg0goBWC
2I8CPgiLiE6e7O9nReYLzQXri3XjSKj7yjytKPP1WoHsHuykk2WhrE5kMbMS
w1EJ706rT70OsoXN5nHurWYIGRV1zFaXodFhcaMbByMdahcYY8KQB6W2nDLP
Lenxukiu2Z2Qoly+UAit4iqCwcj/ficgNEhoxzBd2hwbQyGG6d+5WlTZJWys
RvGLvvNLnZ1U0pB4TGnDO8QiOabLDpC8/1tBDAncfgRCUxAMo8HWI4sc2M1q
RMMYRYJbhmXXhCo9A+lxPUli4JPpJPZMxPVz0QsXKcPnbMwlgOA2WxKAOrfO
GC970h55hcmL/RrdhteGeq/yp9IxdUzKyziJXXrQCBlMD4Cpvd1eHG3pU78h
5q6rkIuUyvQBpUwqow9+mR6rbA6X4zQ/KOnGTp+O7dQ0UKJSSau0tFDv/kCW
96ZL0+r7paLC9FY5t9j6xwqVsNWaRLAdmi50CpcBKIuoKVx5GnwutYqqomLn
p960wiFL6RPGVHQX3hH40CA/wTxUPWfD71fR3vBMYefR8fLCfieV973JGS4L
CzuSUEDm9q4Yb/tIRUoTcYhbDlYBzMjgu1oS/rlO6uPi+Vt3mdtXhdoDQVcI
QrWw9WItHVsAVy3Q8GcDGBdhJB5RlRMwDxUxkj2kM63dmZF+zHGdGXkgYZ8y
cK9oyzwdrCGphCxVi4kIgpBECqiRoeSyCbISMrOAyQOY2vhDmbLTXeaFnCTz
FvW7HICSrbh9n83w4jwUysWyW1yqk5HOf3tJg2cM2C09XCzfXssNxqhf2mPJ
QPCZF97JGD3fYLqdjvMUCD+wpF8OVb0104oZOssg+37HplU54EpHXDC6/ddi
nN8Kb4rWJnP37+o18sdydVWSi6ssAGvKNsicHh6gMx9fAtfCp2N/Suy94CYz
7sTbKIqQsqfaKDzUH+VL1G9DAgw7gl2v2lORr17T+XXkVO4D1wHJXdIvntLc
Ode76HGajH8lMfz4dvkz6RQLOWy5r2k15wvGa+7EP6JAA46kFbbFXKWs/rlq
UtsdxccLxhJVQvJPNQ8refQgVHLOE9ixGzAePo3sJk3nui/QcODLufWM/c2B
6pNnYYa1DDvvpCJJ0C7tWEk+/3X+sjdZbj9dIz+49SfXOCeEltaX/w8E5WGk
7WRJ0rDbTPF3nqrB9DYmoAqhCk/oAX2Urt+6GhpHZntdkFmAHMR4ZK7OdCnf
rJUEYpzQKlCRAQuxbABGGNpwpvH//B0v6zgUbIyKAqLKZF3CLSc5LG1YTcgt
0m0Wg06WsStq9QNdVmj3Zjk9F6tfybZCmQeZogq/rjVlYlWcy/6ffK4x2UHB
r0kvDnMR3kvW3xfVDczfkUyqhaPXfcuZUehrjvnqxH1o252Qdzz4Kd4jJVfr
UUlwLUUFPbzyU+Rj7N05OzJ5mod31KrPwCpgWFBK6JoEOdqDRBe47taxD6Go
+Vjt3utSB7NDLdU8cRWY3BwHIhajV58Q6X6j7L1Vten2GawSpbNmPtoW4kj5
Ozrnslp3+H8z4ST9JQTEum4gDvyNxeBbXPn/yMDBOphcz5W2bbNkOZ7Cg9en
OIdG5jJla1wfO50W6KDyTu+Cu9Sjk35iu3L3gRk8RmR+X2bBy2fyVbD7KvGc
ANd1Hj8OpzMCNPQU0rc15LZFvMvP5BUDJNb1h51qkGl9+nfubcbtk/WcSLj/
EHlmWRaZkgPkuOp1n0ZTL/lnFtTWrho3U4YchXgOr9Wqb06xq1o9lwnA0RS9
tiafwSyt0XfPtTNoMCWetO8vPeQOPzTWa3GNVtjfmLj9QNh/HpzArlZoKIdR
l7AtcfRJ91Cd7/jMu+E10jaezPbFwNI98mb2ZxaqkXYsXCXpyWH1aeuheiJQ
B2Lno2rJMiiEz1frevk9QXnIz9lVJj0BzDn0W8iKqQQkWfgh9T0s8DJJMQpg
6PdHPqWnpksnWMd+o+HpCAxcD2rO3PJCR/j40nY5a8PgqqOAyRI9hlmhzrZc
2G0OAfR84NlhrlmfwBd/fYGva6ehdqoPQOSQ291ldQgAu9qfmAZaO99GpI27
ANsGMbvnTa09gmY7iJDttnx6SxMrGsBvAHX6Cwrk93OJPSRveZBwFo0m3vdK
AMDmzbo7tRKDyMdz6aC6+qPFeyg+SCPfFuYfky0Bsd2NSgUPCXZ6DdIVLshq
6mNtrXFmumujVqtWUn98lEVZQxFP2AryXRP7bQFup5uw2CYBGgoUL5w+Gh3P
45FYFJS//rprt9oGBo7h0N4e3d8vDbcBobuKP3qVDalNDzFIjU9no60fmWL3
1lwizn/y8gzNBcw32Ey3Khe5Msrg1dd1NKkDKTg+VDPAR7pjHyl25v/qWaa5
U7MQlMTisZIqOX9pN9oGf7bciiUZYKHqllFwSJWH4L8lOxsteXwnSdWuy3TP
Ac0DxYLRHbnvVCgTFF+8Xyis1AUbAUPPNpoyd045P/HXxHKoTkcE9RmfqjRV
Jqhuit+41ILoBjzzvnrf/Po1RCOxtqQSojnCw9uPxmT7nkK+gUver33dKPgk
ATYuF0sXAlsiZs3mFCb/Iq8LKV/FVXAmBQlaCWCcyFY/GBRDibDHT+ipwdj/
MQgNgSB6P+JDikAvjaSyPA38InnEzhpy8HpNXMEyQSvtvL4PNEE5scl9W2fc
M84/QSr0oMQX7vqAFxOJwRJKXTcVyPAe5t9MrHgehLdVOWciLyT/+fjs+maY
g9+PducfaeUNM+doS5MEqAoqENmkNmVu31NiFnrmGbMhsbDlbh79KmXXv/np
3JpO2UP0XHjbUbhJffCZXrToF0IXf3rqw2IT72Fy/M7UsPIMsTNPD4N7Jp2y
FxUTeZ8NNRXWB5xXdDfDd0VKqPiWhbPjjBwsyoA0z51jRZyXqyVHwNdOrmMC
xkVHF98s3gPD7kmoff4FqxYSzSig6gQ4ddx69exh7VGqYhMuhu6YLFD8OFxs
PaVcw4YUPtjvQ/Vee4lGxooY1UJnnT+AsCdun/CMaLqmJGzSN5Sy3/javUIF
Sb3GmrN/ATdN2OtHRIttABQrG8Fvoc7Xev1qP4cfIU73EnVL01cq+rvMyYgj
M7wDBCY/3M33A+mB2vFEv0yYJi8YGO9DrkI0a56ibq+GkXp3zNQvD1Mk6iJp
YIqdMs+ri5RX4hf4hYwCOz7MJUS0QDKVqLDmpiSGip6Z8G9UpXoa5sCROBtM
Jd0IjUQQ4H2Mvo+O8iLg6VD0dz6rlpqSG+QUxVtYjPnOFMBuagI0Keh1L6kZ
lYhjUfRmxenEgPuTvwmgHQfn5K6X37FavaxvMxH/O7CRrCK5DmBQmHPda3rD
j73LXXuLyHsx4ZCf37kSaLiblCObp8N/golgJ8NFzhP4A80eO+Yr2d59KYiP
KZLee89PM1jHmD9a+up+Q/WibeP74VD2/fJTdEdBCa8fx+xLtsgvxYyPb0s1
h4DePVCXOqkRIHPWDS+fOM2mJlrSkGC2aHBg0ikvwGZj2DYhWkH658apO9Fx
B3+Lpza9dH9kJ0nbu6CYwTTe3iaqkYzGtKs1CeXDJRdsccd/GcDaVsbb7K90
FecF7Uyk53ZU7peN4GxIXGV7oMd5kgg/9nfbduEhxnBq7Bz5+tfYYdg9q9Vm
aC2oONLUT6wcsGgiwRS1qx2100wYtC+qyqd9y04LRkpVMcJpYT6reE2hcX30
9H5Md37h5vK6+sMHLE6IX7SIMbwzOq6ZFEMx7sglCmqDycqlBEBjJnd50KfW
KYbPNnqezZ8Zd9UjK8kO8N15Qk956G2QRQaedTtn5Fj1RIF+OvQB+NWtRo6L
+r77Wk1syhCbmoIS2vZ2ZWVq/mggpd8dFDw2PNLdromwq10orgp6y/EGU20E
4WCGgejJAUmnG+5chnRhCRKUyNs5q2VLBvde9tDc5wWXbjgxZq3w1g5r7/3O
ViVTzKbBpGCFTi+Qw5wMsAPK148AVSQKuldhWpWXVmmQyZCodgmOqYFXnqjl
83rK/UaRyaOauqriBbVyfSqS3WUzV/8YRmPptSnKSuQIY4Cd1V+43z1Q87zZ
t/7Sgt/Uwmy6GquJdPF6gI6eil5kxyKqjzWRRn2KBI3oDerQd9jNHgovVqQh
LULU6/8Mku5vFWBkyx/51Awrj7cpexC6OU7BuAyy803jo1wsH1vfvxoJaauM
9LHH5zC3n6Ws41fharxQ+wEq7VoVc+jDQu6fTNfBHNMt4YOa8QnD0DGf1irv
babMrCr1FzbLl2Tn33N87CUZrrMSTTKxSasYZw9IxWYsj3ct5Xt44d166pJ9
RHhODrvRzXQb4BCqZoTKNJX6+zrP1e81gpvB/xbQBaymqnP70/p5/AMntIAK
EwPmN3FKx9RHwKseYxQNmUrJu1pLvtgU4Qqwo/48Xd/JrkrKNvXOGFpyG86A
6WHYMUJrYvtMrKCAKEYMS1NVK+LGa1OBZuiC4kJ2+M11wQtwWvuzOT8QhMyk
7gX5sKZ01QqbtI4hei83wwnmGd7uRBrObRZ8NZ5AQ+ASo+gyox9awwFiBL2k
YkqaB4pLROpO36IrxB+ZCcjZ/F7/w9ofsyfvsCzkNA5yKT4yipt7ZGcilDia
1AJM/entooOmy6HJAK1Wa6wnR3woXYlzWqvLA1kUbi92dyuC4Gi8c5XZZSqb
Ytnug9GbKT0d4+Dj1NICyLeTTwJ+se9pw6F5zJRv5NnMYFBHuU55F3YxINYd
hk5zaetAbV7JK7P3SZGn5t+o7AigIxPzJIa3F8MbSZNpBgtsn3rVWDWQnkZN
FHSpe2B2V+al5KjofcT2K2L08kmvOIgvZhZalHBee2yxDNPUZ4Yl8YLKCKN4
D8FF9cyRVezu8zl0KpNNF3ZIrpQFmIlar6PcoRUUar9EKtYemz1eqqHPaZg6
qAuA5duDhljAD1pHFZpz5unaImAR1Tz+9hmWG7Wt/xiwWTZlrCy64v4fZHyD
vDJTYrtGCKZnroBw2H//JozLfpuEBo0fhrHfVZ52ciQG/ktQ9eTUBzfJJeeh
RsycHHxQArkrzB6nDSKhgcAgbaoEgVHvLmnK+IPVbxBem2DHVxKZOJnk0MTB
4p6QLg2Je24zz4FJCXs+iGueVCP5BfUd8JiVqxLv7ZSdAmHuCp0PGcm8LP43
TzkluA5o/3cbhR2IwKxKTVDGR8wRMCh3BYJYSlyCK4ngV6gKtsjvI/fBYKew
XOCEx+mIiHoUwyy5q953P2T9D92kET6J6Ql/EQa8nVxMG8677kJ6xb2g6zez
xz8Kj/+Gs4TMAj6+lOAgy17M+EdjEq+VE/HXyq0KqLV976bvz34QWXOfTy+U
omm9zFSfTovTPL459vHdYV2yoJV5q3G49mRV3hMiKZe4LXEvzZCMcQVdruue
vapZwrtbvSqT6VFW6hZjrtmdEkvqGMskJIm2hQS631wzjOe38mduquZC2KJT
VEssPLEivICftblGKv0j0TuUfBTnXHt+vQof/w/KLc4xSYJQvd+R5qz+sBXn
0JSrLrxq6+N0v9NrpZYwK159pzHlzw69WR8GgXF63Jrfj6BbCgkfGRxa+zYP
TdJZb3r6crT5LtRFseavqtQE2ricDpnD/DqZkLyPche5y6DlZ7pKHfExgwAN
jREZ4+bow81RS8iiaPamSf+4IC6BzFYP0Py0s0fUImnPyltaOQCqOEhLorDk
QD9P1jxxJU1IEPOBHQ+sF+EbPcFsqqvGXppuxrXMf8uUyYGsDBV7oddkVyYJ
ywFX6dNdkKLKmaLdfNA0dl1p3xrSOk1pai2hq81Aj/uUUZjvUhL4MJ6LBLSu
HDR7J7VA8rn2Uw3gMe+3jfiRlhrBj5rqTLU+4Xe5h65CKmisubdSiZfKqZSj
8Zq6l3LjK3w/0mo7d7nyHB3WWPIZiPOXKXvP7eDXiyNa7EQbGUPE+0Ow2NuK
LStHnmQPX3rv1r8M6eT1YsOTY+P9LdwbtJQYxdkHDbY6Z/buft+Z0TySg8H8
NyCNbmsG0qJqmJTuuJT/P75/Acp60Ba0QJikPgrRyKVdpwOsEpScLqlYFkda
fCmQp2k1fmeGXqJygpbBRer5ZRr9zzkHE2EvQvTJoPb8SqMr1o4xM794B2mW
cP+4X9uj/pzDaQUN5IyPNTJy/NaNmHG3/7bAM83iP/3JRkGOlKIVVV6A8CCF
6LDnAUg4f+jz2AVFqTVxl2TpnSh2/QgcBOi8O2inE9PGqP1PrVMTDpYoDJU8
t4ioLXdus3HwVqnf2UrBpCApjI6ndq4Gd51y2yZ0Fi7/Ci5iOhzWTrSOmPsQ
as31Ll2vOWAzymu9R+56D4PYzNr1nqAmF/Ct+OudcsYRzIbeWO0NglCsDEMe
egIFiPzwKyUn0Asmy83RO2RRayHiH6bX2f3LWpunmMXm7quMlJ3gBQRjkvHH
iaZHkIaPO7UY/bdBXbhaa7VVrH6CdQ8MfEFgr9XZeSB5qBOlfM2vUUpNL1qG
At++7KbGR3cpTS2cyqgOhU6hLSrU+m3Qh3WY+49ELLKoP9BtXfWGkZRp+DoZ
V4Jl+DbwSyfbjbrn0mHnvBuYn96CbIXO1sTl2SxjBV/tML5LHtGeGUWwTJu2
SM/mArcsh2hitt12d832sbFz6bfOAypY1eXrKtucmjJiFiV+x1c8z40m4tEr
MuPHO3+tJ4kSrVr3YqmM97lUe6lA4DkV9y1ks3W1LmxV8LiXc8fRgZ8I0PpI
IK5IW2zMYBIzHh35AGC2JmU5Lqs7Vyum0t6IJ25osc8nX6YDJf2d5ByqCSgO
irEfbLJSJBW368vxeJRo/r5nQuATwNwcDnfAWfnGq/rOiK3NacEf23Am77qe
wrOABs81SaDaQeDqnXbxHTMGXwMUN/ffxA9Ew7B/X+QPqWIXl6scceH1ZtOJ
b/XLpf8xxNVyBGKbuzlS77lX5uKlmAmBaMR1+CcCZqZJcd6zSuGNm9B106yf
MvFsR+ur9i6/kiwpT3H1oPrZEdgv68MXC1gSVcv18ZiRPRfy6rFvnGpdav7k
7oLHZhr3rBshwO9rldvkvYKxNO3DNxLlttu0VHO23ISUlN43OgUbHjiZjkj2
CmcuctVu3Xl+zDbwqT67/m/c0lYfjANVjg3Or66f+HaDrlqWZSuW8jjFWfRT
etkhT+FbAKpZvbm+zpN7ewXQv4CRFOTMsBUPmg6qpZQM2wRpds+NndNJb+YS
70OEHMQKBWthbVAtSM8pM1WF39UG8D0QzcWJuTrd9dwtlpr1T3rOFxDtfqfz
NxmlgsuEV4yz4ZMN3+FZsE78geYYi/Q3SGjMJru68/uimgSiTGSRApmpUmFL
459+OI5qzWeo1/gR6vBHxKB2iThcm7gWLn2ZNJ0iDjn7KRHsTEx34Qo22fTu
B8F12arQK3R61SelfmbXzgo+0lLBiaI0t+KC4wJuOOWqlzNAAsaf1g0O7FhY
4bfDU0NTZt1jubZC+t694tp0AFWTIAtIcfWybV14HfW24FxMDePs0oZUMP1Q
0XDExlgdIVMk7YU7hh+vDIYYtFeYiXOtqW/1oEcGy1zczZN6m5pWGVirhTre
gPrz+z3lB18Khj7m/QeuUgGYrAS+kRZJo5ZiZpDL6l4XXOD2kOtgkCTaOWYC
KhMz/BjwTMJcYg70bfIv/Wki2rNSxVmCiEnL7Um3yemBXQQdDIByrgMDk8TU
+zAErivOp3AE2zZgrkbFICTJw9htIl2RxqAZuhW7c1c4Dt6sH8qGEwPLtmu8
hhu1vhJ9aTkYdiee/yh430PfYVbEVBdH50qLAl/QH7ZLaEkooyHhmb5h4vpH
2jVfZs0cCeWqTcSjlfY5qUc1vUbkOb05OAWw0WDYC6y53H79a0VQbc51QGjc
YKlVSkriVj88Fsf5OIGb1qPaMH+V7jM9kwrtOWN1q8SGF2pVyE8iWnAmAWHq
VLQqPz7UIGcT/x26vJJowYwwUY8InQGH0V5u+pKqOScXZs2Cw/uKKBMb31H+
3nsvCdEVKD6nzRk/nBI96BHFwfoWDg+iElOK4zTAJehb+S/up+fF99OP0CIU
TxRF7ItIu9yVx+rJ4wP0zd/MiD6E9z/dGqY+mq+pM7fZf4+a790Jy/CbCJhZ
c2w/mzGeUN+mCo7AkrPx2s/o9FJRH4AjhMMAdoXXzVqU4uwr8yctLXFgKQP0
R9RFAlv8t5ta38fgTkmWfukaaie38JwAu/br+/NUQITP7Hkc0DmNaikHSsMe
A8c/3im4KhpR32U2DL1H5+iBHMRks2whWaZUbaqoGMgYEs9p0yIFS8cQ8fXe
I1cCKb2l42Lg1lAXytYHa8YSBj76PLnHP4BflyudXbvQmxBRJacTnDDIPpDN
JvFwISfb8XfdFqS8CZatEbzvJDNhcW19OZq63doSwXcJSBCZCCVJY0RoC45X
4riWA4yH8We3dmFDIu4U9EWAbOzGfLfREg4f5F42R3ztN5WMmWyByseim4rH
1+vAbbqLKOXmCehgehu4g7qI5dNTkrTxSaa7opY767ndf9ZxWuG5vSytsuQ/
m7uHnbp3IEf+OYLf2cS9GLT0n6cFs7m5OCcsNLnx0YblXWtGEraeHpMBR7//
4/Rzmg+BAmmx/o/cXOnyjxVyXyRqLKVivxUr9AzjsYEesi4d5bi4a8ejecBV
pWU9X3zdBTDaBhY+xC011lIz2U8fZCC61mm7U1iio7nsApJSZpjQyAEyf84L
cXpxDwB2IKbWAgB8IB0V6cLPR7fvsoLdu8/BXyoKxWOl+btM++5UQ8oDvw/4
fLJzcJepZ4YP5QgqF/p6Dniw/Crkm1zNOdSxPV7XNKVE3QXRefUKaJLVoR/r
RMqIfI4EYWDrv13wTs4+VOteFyCgju6MoUBksM86IQXEEQx5cke8c8jxpavH
5boO/3V5wMo9W5gQ2sRBTii8RVYkFeEHHds7E3HC3bRrIUwoJl6I21CQhTNG
4ZLT4u8eYOiLdBKfUBxezjNko1IZuA5OOTBH+sk2WVuUQmIE3PSE1JZBeAsX
K1bX+lW4gxcmExseGFUC/zZS7dyjeiqd75xmjjsvHFaAw0odXmInUAkLo+Qs
kBbYlKOhuDiUZgu8fdAliRW2oLGwz0b6UvVnDb8jCrQ9gHFcRqDZiKojaJgN
KXsuAvji11m12yh0eHAwETKYWQzUx4uMSa6YeAxXLDEUUV0i8jg235j+komP
YsWymZ7SRk4ViU55J3oX1YV70rjpCnkt38fOaOAGyjYivCR96S+iw/4WC7A1
F97xp+4rr0lwR1ez9w2csA5GemPZjl5fMNrpwLwpvlhv3tq2Cf2bgGyWJXFm
IFw8yLA2u3BFq1MRQzniX6jE7U9QwKxCIQ4G9Et4qj5FlDGzsUc9zLBuzmqn
J2Ka6jX1iNqjpuKklerU9NKjPx7CJwwXHU6VBLS4d8yBkrrukBeq50jnsWod
p/2X6Yu3Gm7lMZ75rCgXgomf6uH7byXStN2p2C7sWaYtJwjaBA2dxMHLZfaZ
HaMRydsHduM0/W9P1kRbKm5/ijjMPml0z5MaVVh1YTOrg5RqoQnwnfHU1xDB
/HC6EzHw1AWWMgNVD2160mgVVg85VcE2qss57dygMWq2/8sUVhkpXofpjuJa
8eRgv+lTHybaxS0Ry6DcV0AJb1yVzAnL5phodwv3HQPo9SY5ctTcLJvO6bcT
oBLA7BTEUlTB0MBnXHCqYAIpGe1NBm8iIpBqgFXK4XpRBfUPWPLP7RMa3jIb
hxOfn6ynXKfKSc/FWGPQZphDGRWLBDUPT+bwcR+PSxgbpVeRvUVt+jebzLqQ
jfjx9Ug2itmh7VKworWQsmBSvFZxd2qkko/sXxJzKXCfiATRFO3Mv522ISaN
BGPjVxA6kMucc3udWDakX9EBDMoKs2jlit4kwuSHW2IEFcyin2Jo41Py9/3E
VJzeg7LST/hDXJlRB+BOXUAy1GxMIT6hTRBi+b08NZDbkuRN9woswol2psHD
a3afUNXLdlpPqgsS/J6ybhfNKztf8/UF+f2k44cDe1qxQ2PwvYdCKiWIBLRW
RUkH9qrsH4GTkxgkjYkb0RbrdBvJAeGI7srfJjXdXuLuSqSAb2T8aV92Z/HD
2a8X5mPzKPXs4rai8OLS02wevdzVwsNi4y06waA88ia72q97zI5YXQhJKA0q
JEq4A7mPi4tkVvx+2zxCLIWve3DwlAmcTMLAPM0rLLCiymNNOYkN4rWiXUh/
HfEdrIArdZOnaxM+Gc6s1CijkKMqzBhNkhybV7cHfM8kZHRosv/gIMXFLaDL
gKzPYSbTy9tMbH20uhVzvmYR76S1vehflgEIplvkrymYtpYxo6uwYObh3sZz
bswCr0jDbjzps7hlU3MHvpQpc/bApOA5Il4sLBAIPlLVxpay4nXCoyeb0SQF
m2XNZuchFY7BFloJNATNgmEmTlQVuidoPMl6j5Hj/mARu6OuU+aDBZNE020D
OQh8M+RmRP+zk9s+U/Fo40drxu30ugy7L4ar3LTBgPfqFLy9fieJ+sAgBpQh
zg5nYvMVxsWMf3Y/CKkIcrOURxnWxrr521IbUefFTdEFQYZUTYrrly6DXlVl
lvfmlJRqgjLAwI0YXoGIaAPofqXADWrea6iJWY1vHR55QL8I7E0ugxbv4t2W
7Lu5a7nqMtoigfgW3ygRLriH2bjyxXky2+FNh5RAy22KSQyZi4JFMe7JX6S3
Sx1sV6txSqtCRIgOBTrCw+D6Rd7XCrMI3Zk1pmNVZcUZmg/i9DGZdX4fpdTD
ECjsKOzqVwJug5TEZnxIwWyqhMDIOOG53xZrGSDZblEpZrYjnmBojwswVIos
i9CbcXzTPmeGxiZU9kHA6dadGNUU7D5jH8G0KQXuHQ7BO9C9Z/eQNlmi0/ET
9qFivHBz+jcEbcCoa898CqRIAjVyCCx0cu7O1ereaE0/ZczeKx3YUig2nJIu
B323ejo8GsYhDKA5BKsLZWKGN1w5cTrtoL/rK4wxgmvFEXTSRJob3tqvLs4T
Xh0dyZnOLibEepastPrtuKflwl8cjx+dsg7BlEirVw/H9QWxQYhOcIvd9d2k
SNmPw51RO5GPyhuLyEHkpk/cetX6MgB7IRlANbgjhUVQjJx1R+tHDta4Cejy
2BfULAespCcU/r3LMtux9BCOs5R3blfn1eQcBDEJcHCKLuV6uSYo2jQQtTro
G4RNs8TWpc63WlOzDTDrWUjHZdxLtUGowvLwWTSekg3YjxAd4CCCh7ctnatH
dFsHgIvbsDdv7O7RChziCtIWvGbXk1hmfga+kM8EB+z1nvCa9D6a01UEakkk
3wl6DSFHajdwFC0MDU28ny/VcdUbgUiR2k9M/9ZR6N3GH80G91yDOG1dowaS
FgW6EDU8nA4cd0gZN4ivesjbREoHfz6/EHI67x5uTe6D/dB9WkoMhYTZNx7L
ES+ZA31Gs2Efo74/N6ukg3WWvl7d+1O6ipfEk8vbjbBEaQYxa33Rh+k75m+P
QCL/hkIt9hhvF4mYLsF33G4uFNe7nedPerYX90yzy/Ue+Tdn9sy1CKZX5EOi
3WQdafgqJTyPjQFHrGURL8cSmfkraEl0wSpLSN7TUU5b7cfmIvqwXaHBmqht
JHWsrFw5L5GvORvjYvBdwSI2xWwNX4yTMXtmzhcsbHGaym4x2g8l5672z0Ox
ziMmsg28H7gpP+mtiHZoHsKsZ29lYgbL1QW9XNAjpIC9kuz+U9rbZZ46/0nC
QQquMCJva8yBH71dfRMGywNDtilXbn1McExNOFJmHobQYJeye+0MDBrDMtVc
VC8bldU8Iyt8msdDk0+XYCt9kc3q3cPiObTgqDTWCgs2sJHvSWobLqXV1nZV
K9IaB1csRK2oT4URB1m+hMmivaN6LfRYRTrqFnS11+950blHn+3rvxYaRyYj
OKATqCYshcDx8am//q8W0r/FwWhrkbzdNAdgLWV/gjUCxDoZtpd49rnUe6EA
zbbU3SthosfXdGC1e67pg8/y0wU7aI4gBvK/e6ifXVG2JskN340R/WMT2VAf
uBMtGfU5vL1mTqXhgTJOXYtNi7OY6rTwoY94szc5UXdOiykHQhIVE07C/6E1
QXSlY2OH8P7B/WqiFy/fMTYoj3OpEAKnP/l1Crbyeot9oswjT6wSJBr+yZKV
P+QJoUIxX5yBx1h2wHIky6CnA423Ne4NRXJP4TffBQN1uXuzCD/ypVyqLmmU
lcCeMLbYSVBYbRAgEk5JCqaps9zfaB4ed/BeUgaN/U5exe90C0DeTpsEax8w
qZa9Ein2fduuSUb5nlv8qBejiN5olFWasciP5Uo3X/RaZIJIAM/Ki5TFUGkT
FrJWTxOaviyKf5NiInrSZd9tajB6QoGmgIDeS6MqX4ju/MayDhUUH9S5IkGF
5YJlpOztbFT0T5GJnkG/NXsfy6seSBT83UNrw6z+0LyBB+7qZdx5HorEEoMF
XOz8aRVfSLBRGoDJr28NDkkljE/sdWD6uEuUmHWJNdE/44tTK6zRzqWaAJR9
j1/3+Db+1kLjCzZ2K9h/ZuNHtzgwRM84GgrxApu6y3m5M3Sg1OLsyTO02Pq8
Zyfis7ADHWV7tBu28elTvWODjq7BZVlnNxNLcjCL+KJppGNaIyNmoQD9DZ8I
SPaxQ0CagmZwi4Mborv0UlQ8KdYzymk3QF4eJYh2D7VX9GKg6JX26z7LQcgg
GaFWvcWwqGmqCpe075b7arb+21dEXdSxNSne1UAQ2zABD1Q6p+RL8bbfH/Pk
YDy7GBDuUcLjza/x8w0lJhHf0GQKgJ1jvDYOG/QW42SzGS8xhegYwcXjGQCv
3gL5B4lv7KSV2WgXba2OXSIHWk5tBv+ZX/KoNGl3W8++v5JDAJMtAkRlqZkd
h/2GaOB/kzc7VZZvlRR5ZquQQw6TrAzh7bOlIVxzvLuf6QJ5XzBfXRj3ybMu
iUsXcaGz2MWFAk0mdDSEMWmJzXShy+Ow3/aRrlgKgZT0B6qAhXeCcmwERZ8Y
cKbr5BtxYbBvKmhPS0J8fMFSLvoO7PTZZ5s5cU77TLq5gInmqhyq7SWBIwsf
F6VzFuGsaiJAKuDLtszf0j5waC5P0rjXOpbdLxshxe3aIsUFJMgq9jvJ5bGP
vBeqQei96KOziBxxmIaa/CXpmMTMMEp6IesBsUUaWZ/2R3Pmxdg+ZNJy5jWV
ooPPoseMZMCRbOos4OpKfEjJBHoGCuiwAzLuw4qxApldiGDuEzz/tnf0p1C5
c7iuJ2mb6Xpkp4nLOlVo+WdtG4UHIyXsqKQyf/XwoOBGqb9YiWdTSaK3Ffnq
TvblOAApd5dbCFGVY3QkfsaxtRWL5bAirC02BVL0Im5/VbeEGASCg362GDym
B6n6j0BXQobj78AJN69z2f/1M55uMg1qIGYgRApXhjAygArgK2C3NCua/PmO
nBjgtyiBNrAoY8QTBJKVWphNKk5YXFCO6UjYSBShcCFxGfL82XkQ/sOUg4Ux
BGFgNzOX7BElBvkrp6wDlOUzof/S1cLlyXPrOsji9t+Ys6pnSVd7NRVp3fUF
MKA5dY5ZQ5cS45jOCunzmkIQUjEyJzaLHo+rOz34XqwPcMxCN2Dl1TlnkPXd
7TYy/OCe5JLcp1rYuxBY44rzXvFLFG/CLTgxb5yKUFx/KnspGtXhYtOie6FZ
NliUnvvIyXW5BdUPmo5n3NmXTXqVJLyVKJW8MCpZ5Cw+J/iXu+tyDZdH2c0o
N5cqxMuYdF3leFS2GvKBnJd/WQERBR8JEd56Xl7y5qr3BYbMp02yLt//s1o7
FTxt1UzHmA7AQqGx6SVnzQ3ZxW+hToDVNGP/ZChIatTyiXAY0wzxxY4QATnY
vma4k8TIo8iMYsIxV6ce8f8J9pmbfuItFykYTCMRsR175TDoXOtdmXx7QTaM
vxPNtUEypB4fDCSDF9dwtAzUIZxWwATrjGI36aVBUMhYH9ZFMR4gKPFYrQHK
sZ6dlY3D+WejsAn82fNEXG9tIOVuNj0/JK/E9kKoIhWdgwhZkakIwVRrtyrz
Zx0NymbE+52ADM+lmlMk/wC7ojNm9doqoCXE8bZVLeuAJdj9z4Xxu6jZhr3l
wH0RtcsN2fYJ2vFmLPS4IzlqlFY6Kp8/BGigLyxv80xubq7i+9gh9OfXErGd
hrTyTFa8LEaQMxjm/RxGO7VEsCAtSbEB8iBn7a5FqlDmEmJA94I961RHMuYw
p+HF0+GR9Yxekjkw8czvya+AwchYWBL/Vrh1uYmD6/xkEOjOGf+0vJFBLtpH
BwAVp+PMO8/83uxoOpjNLvrykFfeSgMUlv0hGicF++AGpeCs8Iosd1EGiAMK
8nzjoBkEHPY1R66+AcbUq2O4wZaRPYYRRNx7+sNbsO/roqix80sBXZrXnqtl
bGGd1LW+WWqS4o+dN3VKagSM2ZCzeZhnF5p8//Mst/dLieTwKqppJHWo4Y9g
3AMpC3e+KSCDtpIfWADorO4DuNfkxLUuHGCzYe05tKyoUNjaMwUvhUVcgjzE
BzANJ3GtSsOYSy4tLsJxgYM2W1frXKVbl7n9/0EuzsiB/7FkJVgCOFLDZR6f
zJO9XmR3UeE9hFEQVLVPhoW2LekUHOxLRXdnIasn1d5YAXvoGRKzeQnrIb/g
6xAb5xFHjYOct1IM0rHUaZwrxkuxxCtX5J+kEqAKjkH6P4flsNNB6jtFZq1t
xpEyUrgAmZ3NR/3/KLxcmFUJgsqbZu4khUSJgLcQqR/1Cgi/pDbX5fpOhPxx
QmAHOn1WTrN/sdXHHuc90uPlsR41fsdMbPZE023J1rjFCFQOYtRiB1DnArHD
kxh5lz1TrrwHk5Bgdv0Lud8t94le1zkj0ZpL6E1Qzuj4pdPuO+A0J7wzMDT6
TO1KaBRafQU/gDrTNhm7UreAF60N6on/Kgi4A5hiUbe3C0rDTeSP5cbbfczj
mjClZLvREV6ZIlYg7V7Qtb59ej+7v2kXA+LhA7XP3f6b5sljiQxYL7+JIzME
1EK8THxvlrWa7tSRzMXhopOocimSkOi7jvH0gh4I0XWhKEMqk7eZmh8mqndr
BzKQ5/5RHCz+GIfi0wfgkL+xEFMyGIWmPl0tSuBk/6yGu0zesr66T8GO/JF5
ncaV12whaLqVrn3KwwAYFxsmhnjPLL5LkS4qx6PM/Gl0/PYXodq5gzsXgxZL
7NzNwqmet4+lCU3sPyyFwLjyEh4UNTvpqbwWh6yxko3u/cjmCFzZrXVVv0q1
oFPKcK2mHkXkeuhTmlvsqJ3p9YtpE1DRYiMKYHSyMZ4B/yCMkDhlshtZT8v6
x5XNw3t5TQajdjmElcK9pubkJx27NNmk01opDxgW0Q7DwpRnUcVdxqx+g5lc
hnDaj+dJAKGZBF8OdDveIwJbOjeVWqQ+RRE50NI0vr+7374sIhP5Y1sD9+kJ
d0GbQNaVo7PtCZdFkW91j1eXpBh+ozyjdvyYc7IiEKe/vMIKT9DzrLbBC2t4
4BJ2KkgI4Vqe83+284b7G2Ub5jiYoSCgYnBHOFuqsFd3rFBR9KYAe7xv/PzV
zej5L5ggPCjimo9my4pILm/EeBmDucaBOLcVb+B56VjvjRhEsi9Bs39GaUlA
0J6umd9y3UBFObeivzZTMuqeJpv+DenX6p0FCbbjyqFK3nowdOAriolsljTS
7DJaAZ8OxcvhWNSGA8Uh3CPf8xEeibvu0wdrsENV5DaYnORHI/2TiDTXOBdW
fLRUx4RxhqwjhxTxdiwL2bS8vUHttXyJo9VTKyALmtwFDq1p/uUfZ6oEDkIk
b5556N9DTzVLWdNAMeJ9ZXK8vEpG6+z9gIlh8hfUUeWAk6GZbKxHCAuad5Wp
tzmb8yyRdM2HGlyl3sPSl+kCHURMp98LKhoOoRE+hKulo9hGvdzFsmswRIGP
VCeSiJLYkHaZGt/e5rimKmke1GXz0vnIYQI4od78UFgit1HgwZV5nTH4ENHT
xpKzRBbEDoX9iaCbfr0RZmxMatLVNh5iuRjZ4kd0UM08EVKyYUSVMpnxbryr
hHbTCQemyGdG8gYxBfBXlE8FAJJLPU6GTHXO205Zimto3MtNO0kqK4PogOB5
kkyI7Ld/QiBeX96svya5DewzsyC6zd08BcDoqP1PuIQxN9ThsqPtwxisikXW
8tiDHsG2Edk+eZYdBBBPnrMYeV/aeTR412gdQLFF0TPDOYJDFIoDld+6qH1n
jp/Atr/gDW+qZvJOUaoaBJP4KO3Po4SnU8c4majeB05SfnEHO3c4qQ2sEBnA
sQg0/jHSeNt3hdtYoeERQvzWhIr04IhFc3YM+dEt5pqSMNKq5uiHvPe+A+t6
XJ5HXAlfLNXcYyYd4ntxWCp5CothOWLEwWftJwpUYX9ZiY0bMxC0wxWAkX7k
jFXLwpzSfQbUn5jvrC5ZIOKzBz7Hqh2Nt/7b63XsugbeoN3+3ZRfz+zh8QyW
nlkwYWKkiGr6ROzcyd+a2lYiqR85xizu+KScy17dqOoNq3Qls7Ooi0PGp1GQ
if0B8wg8EvV7n6FyDXuvjUyrUyPSJkcEp/Fwt/ngQZI+vSVl7AUUelcZoRxu
iYKh7jkkLccDWZKeoMYZjh4E7pEDqugZlHAYmTBd83YbjZF4h3yK2vvwx3wY
3Q2xtmK+fwHUybNa5FoBlXgx+lM6rhzXKyfOdGlnOLYeyF7TWsKRjSz11MBh
GSQQ4d3MtcD5Mslr3Z+CI4IM8TZOz4jGan/nVKYAg1hJ1vdQr1DSLLCBfUFR
E5VVRotFDZ70dJ+OCjmmvaTouPmoSltlJ3nYHFg67dys5axvykCOQYCkGi3S
ZOJMGrtawa4Lz7iI577onXqnPEhlsSzj1OnVAwCre+9maExqd0K2Ld/31Ff8
LU5uB7rIGYAtXsTS8EUP0HfUG/IZghbpTiN8iWOSdBvUaFL+XxbkE/L+9zFX
9xEf5yJ7QkpMOsXH+TR5b0Dv+YfsNsFMdIuzUd7/n44dMAZsTzyJwfqT0dQc
NMsv8mgqNsnqzYIQpoNnwkuZPHi0NIgKZbAOhaNJDS0H6hMmEyDDZt/f6I4F
SQyTfVhnHOrlQR0cTxi0myWWqFOM00q0jzr7novkd0sWlsx6ciyCY4KBnLqK
YMn/DBskLZx6tNLOlHqAH8UwiTxUO8bqYsi+LHj4lqFNmHI6ORHJY8VQz7F9
BpSUuBIxohyCeRGC4LeiSepp7mI8k8IHOPzz4LeQavyxZi6rwQji0rkPAZ/F
S2x08cRPYq2s4/ZSE7LQKq+cupalPN/MttFDsD+LnyT6zNcZcU0gaSORBx9Y
h15FKFuzVC/AEj9tCrVA0Ion04/8PXV+lGzbi7QfAblpUBU6fasLH/fC0b+p
ZwGoRJpa4UVnCAMPsgKtTjkDr6M8wXy356HpEioIOsIaSKOE/G7BpMvrG41i
rTCED/cYHzXxZeaLCYSJGAm8r6xqxrStb9QNjqL1sZzKeH+eAhLbwEfb1dbG
oSTyvi8eI+d/i6KiiIKMiHteaCEvBMCT+oTaZmoc5ll7FJHXqS5SZf2ltQwj
PxMHVD0QkNR3QiyS4bwdiY+PIiu5qckmGy9eLB/GS/YHB8d0UDbyddBIaQ0x
UG3eG07NfnMFuiagD40RSBhVqNYvSXF4u1f1+OOHpXZIau8Xx/oo+XyAxtBj
lhsY9L41tiwKZtXn+z551Cq6s5JscySs0W3OgpKxRqAkOJ0TaknAENRsM5lv
EzzKYJZrL5hUOH0X7ehJYMlP3aTkZqb3FphUNgILsonQIStEO7Vm4ZQNXCzq
Dq+/w2v4uzuj9kBSLEIXxKvHTrsijcILr3ngLg4PkYeAPuA0vjNbbcAyaIJL
LS5vCkqEUlqMD74CgCXXZIXept+b4z+ZOiMf5uHjipMqe9jBrauw6Y4uU8K7
AlE6q3LdbCj3bF835U+HhBJFnPtIocXMrul9yITfoLx04Ek+yHUVrJgUva4Q
qW2eFcs7Wjp1CTMXzcNUyOCRhdWITfEryEthHRn4K+7u+1NoXGBjqB4Msw2e
NSemQnbd2UuxeLPFCoTaMlPzf4o19ZlT1ON7lgABjD0S82+wSZx3Wd51TmNc
kY9gKmeeWXWcOcdmpo2PoXOolWGwiIKPY+95sErh6p1kWdlZ8b1xBHBy1f+F
QdOLcJC8rgGEMOLtP+Q8jhXwrXumTyMQkK/9ywAqeScIF2Bu0p7oOGzsBL7J
5lss0dSQswwNpCgAypqW9hUofdnaMbD7VKOVq0cKQNcYUikq+7T6MB5mR7cr
PqVlfj/oTzy1gthg3aeugpnHSlp1aq/YOHVe82rgRSfB2lDG4v6cmBD1+Tz6
v8qYvsSWSQNNHdefHj8u0k6Bwory/Ft1HiaybrHmOI5miyO8fMj960R6oP7Z
9uhL0iOY8ph/w1v07H3XWhvtMK2vjHCYQwdITLSccdLy8Fs9gCPjekOmCPgc
QggsMCn3Ab3cZUlzO1dGqhT6KJh63uDBPhrhnRZ59LYBSKvFFMazUGreddmo
ls38Gu7Uyf4TT8a1budA1CY1GN8TsW4/TfCEXsWV4SY/1a3nt4eAkNoiT/gP
ofEORwmFHsu3aZmgZF973g7JR09szpJQWHE/cvn205lToPDDHS51i+GpJoSc
HpQRBK4008LepM0mwHNx7XKGyljmqA6YlDaBepb6AzlxUnj0L43k9lHbrOFb
QKyx+7AoQHbGBbotWXU1nGDRYA2cgr/eLGjUPdIxzYfrhVg/fhFiQJpsqg+/
0dgF1Zg+EIKqTgKuylYCodQtm4iHHb+LdtdSuo8L9x6XNALdkDjkTzp/wvXr
vfBlZUE2sOiH2F7XhJ09s0MybFNyaDSd/F5kpPZSWxNtE/OYzGLE5GkSMX8I
YmdaEh9gp+vdQB/uhZyE7ONvm7lnfIehEpvCj08xbzWhk/mYutrzcHyqtahx
/PgrtpVRvuXWVyiLPTl8Y8uEBq2czdGQB6N+Hqbs3oJ8mRIUVeA5M81WrH4H
r2gdkzmtPfP0/7ocJ2MY1F0aDFL4ynWUHwSmC/DLuSjN+Cy947qjEKCO8IrA
trt1IB/rhUDpvFkdaoH41+aFhz5FyYbTSHYwHriJqPftrGWE+Mkz0FleDItz
98sp/Dj+F2kb/OfY6kR+jQry+X7O85noW9tg4WXDKnXw72GeSSt6yDal7sPN
8QAP6u9AbCW9QxXxluw7FYUZpiBbA1OJFihgudl9XGlOi9khQcF7mKKQFknA
FbxbhiPZOIGFYy7YDrWC5CB8w4H5VPH3GT9tLcDnqx0da0+4rwsaSdteqbOL
8JCAgEecauvtSeH4uD0zJPv/+ndoZqq4nNuiRi4Gerz6DZZuzPAm/5AhAZS8
4HAkB55WuM1DOCbF/yobhu9PUWMWWMmQIk8aTvKeyu6jT5wUrohtgSa4EKFF
3uKWzhSTN5PiOw6fIHESvNkC+TsK8bphLSjh2qLv4atkB7E3kVtQkXWNg78f
Ix0DbSJMEQQ71pPupvQWXR8bh+jJbpb9XZViV+Si31YpDlLF4t63P7xu+iew
Hwg+DQ/i7aGOLShNeS/As44MJRGPl6GLhpw3/JGlCBRVIkozQuf2lGJWBBIM
oSnbObrQwxIbC1FlrNBhsoh3RXON304rYfSP+TUy6EG6sPKFJI+NUmOW3r1w
n12IiYYstrN1Cnh9HeWrEGhYaIQqFywf6Gcm4i1gMz1meImPDoHvP1WlzW3i
PyXy+OuDsIzb5bA7rixW5UNtL1lwdONreEHO0tas4ittPEodEZeNSEcYHyr6
xG7P+2iLVpH0k6XFKP2qzQEoXPjnLuswbAPu9iRppVoRDzvjFA8DFilcQUJb
3a1Ko40u+WhO0W6MRhiMFblMXyO6iFKe+zKeVn1mXYqxLy/CWp8bgV+ofHjJ
tBBzE4VH/jdHyL/0HtWIHgfhqL5q+TYQcjyPUZnuqs/VDzUY95/J1TEjGOdB
UD3wBr3mPBe4VgqxLAWxD4Bdr5S3XV/tF/XiaaSUHlCRf8OjzGRSWpSZCAoW
/6H8V0KFoaXRBUJSFkB5Gij0pvpZJ3VAQjG8RGRL0Rme3GHsmVQaKj1xWY7b
S2CaqjCX1RDbaJlWbWXtBXe+WY4UDFAR0Cp9xXd2y8Ap6Uak33vSc4sO0FP/
2zPOgYCi8u/Fs8nHUKpI2KAl8QphTgocrHY3N5QkpB3e7uCI5T2rUvrh3okr
3Hp9DgQ4aevIn8TkNGuR16ahg4hOeVVV2NTEIlLONsa1FiAVm6lrVJMnlRQS
Bexyqj9db5axfGwdEQkRa0symhNgI6eK+GTRSzdHA+RAr+jAPjMr2nyx247R
Lb8Xb6q4lajzFlUn0qCEW1MG99kWo55NKwfS1HcQGp/5GKG6L0jvSSSdmks4
DFnxKY+qurg2cRdFEl2RxKgd4/NA8kpU6dliW4ttiJ0f3sfPeQmlIE4R40b3
QtNM8P+28eyN/BNUXX3MLbYLumjEyov4P4kbxwuPR1FdfUaYAN3XeylEyCVO
2rIAXn7yjBlgsva4k5WP0l/eHWIk/EQQgVSyxWdvKFN4lx1vUcJUSrzphVDx
qp0d8yXdGvjDUl9NWbapg6C95ztUEOpXWEkfSn1Bs8l/uODgfUw5SFwTl2zZ
dyjgVfUFn/3jBazjngBnBVbW2HUIK/po933gB53BYYRudA0grFyW4DNPOqzs
R+Pnud/VX+qYqcIhyt7KEraQnoTTdKw3O8QQ+kdindIZ+5a8r1z10YV21LnB
gZrKgs2auf08Gvl5eoBTGR97gLbYEELBeSR7rg9Hh8qC/Z/0L6zD5yVclHub
0XXX9kQyYrX/iOAkxZkER5GPnpXm5vPuI0T9WxQTGXIJ1DpiEd7ojo0LIGN9
GdWOqP5tZFAbPsS24K2G5teJbqSYdx7+I6kLkWrzXLKyicJJAylN5+4KNORu
IZiaIMSF44vaihzMj3nt5xNXl/NPi3h/kDxVWuV3VlYsuwFhAeK44N0wcJ40
0NdlTV+IoPk+nN+PMHJryndO6O+7PW8koPssfgR7jWlfxq03ef4Hq7jAV9bT
oxSfTZpZ718ef4Fqe5rElqlMvg15fgWGlTVbnZaJf95VgoiIDBtgssqWcE42
4cudReMsdDIGpJvFiT1fu1C+jublKXiEDq2guim7/C/pAToA7ntup7HSgfBS
Tiq6nC+BOaEieMfAIv7wQwnKCQqA2JGFW4Mo57rus0deZRctuKkrXke3uEsU
biknBOBf8kcgblFdvbtziwUGMyF9o/RscdKiLuAZLQtWmMsoFDWtyRnqOam5
fvCwKp2/CU+KOyiado7YGQ/BlqgEOYzZ0AOOadCt3TzGNZSsONqATpy1z8fI
n/tSe9iS80nrOaJB7j938aQER0pv21CngizzaevN4HCmZA3ArrC1VEyX8xxk
wOhe1b/H8vCEhX6VIWN0mmCEluMePx4CSVv5tDljDUaiO7QEwV3qdVbGHxCt
Y7NOuC3TJhKROPGK1yVRy9Wvgtxumz3Ta8hHU1TdFyZDccITeqkbZaQGRvh+
Cndd3oUlf5bmyfPMu86JBUagg04tl42nkcCgk6ONwJGRf4IwmuUqJqdiAkzW
dDCEuS/ngTU0HSygbpIfh0ONpYur/beBam0SqrblJSzEry05AflPHlb6XcuD
CXvy2S2jT8nr3DYJgjrjl16T0B78ftLn9kFzx2WW6hievv3aGCg8Z3HP32pr
SsT36N5dUrMqUBpTijNzZKrBNYLb186DYQyQlF4MiMlE2X8ARUPa/YhMhRPz
CyWNnvuEr8FTy9mioYZdjf1FAGY+v7TrBxvtU9OMgO5x0CUN9WT9xX+xAcX+
HRGU9T/Xt5pFP1fIfbQqZuRsgyE+22a8KhwUH2+fz9C1HFYc2mSLYuArkxP9
fFKGoEEmi9fyCyxp3C10AApzCar9Y8nin090GYJmuDZU2uepUvXgQ+nrr+9m
aWP41uljCTKYIvNXvyjDD1/CrUotjr29/MNaEusVVws5OH+aRuen23uE4Feq
NHVEhrtVi7/Y+O5e0mXiu7bjeS+oHdvanwIePqDcBP9kFSfe9bOj4e7xFPuO
zvCmkINKBP3hJG6CYJf/PMLW8ciHU7p94kPmWNm1S3FOpdGiOG/UXvyGucJ9
o1KF/j7+RVcKI3j8RdS4rYIH58XNEs3fzFuUtmLEk9gBMYkmaV3IqqXYKtdg
EvH/Ef276c98nnE+5Jd06y7E3PAZXymna7Ci/zVk3yxa+nMNW7ROnU8Xte3t
0RRXodPp81tvdee+311lmOtIL8UOIuxUYbqucGdez8M9ASLAUSSiUUFgaFbH
2oEGrTG1+3D1ZfVH0RgICfuQkFaukLjx87jthHH9lBcatNJQC79HLZI+MZo2
OF7F149+xyjALKA1LrGUtwk7K64Ysnsn9iQDx5P2mafIFo4OINWizaHI0z0X
ZEIYUzamM9XljLlCu4ANdkSBessz5d3aMn49h7NP3zvwLJarH8s4lvoAqB7F
14wyc+hem1GGXJu7uBsTwhV2JrBcrJQ10lWwZm5ZlKvOHM4Par89msjhW3Ek
msbB8mJALHozV7uQseHo50EA6A2Snd3adcCfSsyd5SgwzRF9LThbyeHZFyUq
OKUtwCb8AylEGx99QCeibYGHKo9XmpVS7Dz+wNcC8ZIz2IOPXqJJR0vM7jRZ
Nu/xO8Hh315uPDW3ulncx+B4qHLVtswGrANk1IF6ZSZxhOhmpmvSUm47HBBV
mFa76kE2a+s7POVAC0MxeCR6cOzqGas89X5mwYZ6/DQMAabGnBjXBWmDXP5z
ZVLIvhH0nlI7tx36isIl8IeG1Ct8+zMFqbchsSD1hF18q/24D7WFSSxxSqwB
AZucXlz9mkHgWixDyVdNTffZyyd06IS5gb3j8KSAn5WaeQOVxjugoiJz8hYu
K++0kFoZzGYCHMQDbS3nTJEBwFeiuWdQufKZskiF/HyKf2DuZYGzCoAKUAdB
dMU5gOuQ2ZEITmRqqFyq7UTrzLQ9dKFfHhWwmvPUVptCXSKokzwugPUhcB9G
GB4bQZflq6LanAI9KOWIm5trXNasxSAcL3QK7zLmr4sxSTtp1whGCj5GataM
Oh0j5vQJa1unxI1ftL98PRAmD49aHHJ2UwzYRKODul1zTDpQhKSLOweqfLo+
ID/qI+8EjK4+RSTzifY9Q2VokzmoJL+XFVMHOhyiF/5KwQn/wMFrGVOJPt4N
V2nBdxK4pKbArJDkjlNVQNt/FMl5W4P1uGEluMEptnasznJrii4/UJ42VQTV
/GGea0A04G6Q1v2AuTgYIa+hz1RV1prRKW8DjhWQBGWcNA4BK7hFc+1VD6jE
LR3HMInQ38KVQAzccRFKbMNO2TJTxrvr7Y6OJ8bwOYA10xAHILKi7fyfneE1
/A7Sfwa7nxYiX7JMMWhjxRJ2T1b/2yClU4WoNz//TvbZvqxpm0beCXNQ6ltE
+xfSimJJw823IsPY4lWdDtDCJW0s3gA4JP5R0u0E0dz/mo1gyUUjM3JIWQtW
Tj9oDyhpXW1OKGP7DIkDdi/zub6S7inMg7Ha7kTJKoDr4VFfkXce1zq4oFha
ERJ13FR8pUUeX8fJ+i6KtpYlEmqsY/XqxVDL7+TY0rVw4kXLR30qbYvdD0EE
kzf8Vaijm2zo+YBRayphnMb7SU9MboMF4mYuNb8JsGaMQLAdgUeFnbv5kFCW
Z6risnsajE59RMB3T7H6ygcElazgkSWc0c9PGqWR+ZkUCMjZVFN53WMNLu4P
dMDfAYhIsmf7iTOgaEcl67sXVyi22ZPRoWuHomSnLmQkItdOzWNt/Alh6INY
C22jrGw+kfmtv06e0X5uWLtL8a4QMswuUdlJpJB1Laf48QloyuHINP+403h0
GQLD5DjihRfDB6RQIC3RekZRjkUogn5J7Eoeu0C+HMXteNUm8ryjtj0JNaar
MfhfzxFMKuX34okowT289kPdhtp72QG9r5ymP+dq0+4rXYlTQqzOM8tk+O2G
Fx5/Z3HB4Lk1rtUt/m0ny3CamtcrgnnwY/iRj4YD23uxUq+HczNiiJVt/8eC
szTPPBdOmbj6e4V9CDH5laWVebSN2YiFb/HtMYfVjgguT0ZFL0ogaWMDoeQx
koORkfKqyGsY538RizfUrQC07ZZ+h1/b01uHebWk8SPQ+I237vCxAUYnIpLI
BFsOTPn+72BoQekHWD82Q/xCuXZCkRAB2r3EZhAzhzDalVXskoyFSRC98dKb
NKtmRxOx7JjiZBUazIOYqjE9qLeJTzK1dYbkmR4K3zxiXPa0HSnANRlnK/I5
8dJlJAKE/J2JrjGAEDnLwBAxpWADLjaqhZctseYIT2z3Azi3XjOFe5Srxtrq
q+r9Wf2ySYMrwLK9tUoMuzRbvO5ed1JNQYDxYwKmbxXkB8GNdwXkeBXTBTbo
7E4F+KHSxg2kp9VC9en8f0ndHh+E4uHtogHk+LpAGdRThjOU5y7Gba/twpCY
taprwu7yum55glILdCWrs8FXKzxNuyxvugM5XaLxy1x2AUvJI/2Pt2HzYIAh
zMTQ/4baOVJsMmJOlGX/FGFDuWHb5VzjjZ2zjPXMn1U9sjTko/XUCSxd0VXD
4Hguf5YQGse7XVwxPc97hY4o7bcb48M6nCuKb/3hsNPBWRXrh/6eULWo+Mwv
mHqvq1lkccAPMzQ0LnEuCdX1wy9y9TjlaMbkrZtamhlkwOAAuq/8hDF7FEQ5
1N1FwxZ0A6gHMOYkxS9+LNKtTOZ9SKldsx3nVyCu5aLqIBmVuE+2Etq5tMjl
/WojkiK6Dy5ftI8aa5T6zDwQCgvCA/4H6a3bvJ93KfZrdOD2KRSTbgqA4VIm
VxlenxeXHdD5Y+7EhPe+Q13cPRtAd+loxGcvM3aE4xSJAPmCI5WomRWaOFQa
TWKaPHyExUg2dY/AYqq3P11ClNAQy2kp5NJnYcZ4IZkSTCWpSQdIBks7dkRA
eSN+13INzwGu2VelD/ucpi0BkJv+MfkJaG4iamvfVW4yKw4KXu+yqdrvn8XJ
ZBpLXY5XYa3SHqL84Ffob/fg6hA//jGNPi5/4TZTqRwHnk2ndemNgP0fFpMs
UbJ5iAByERmLtpeoi58j6LmEhwwzk4EeZ6u9yUmo5vbwRKXBQwNeka6D0XF5
bxiqZa3OILEfXkTFRdAnDZUd5zLuGy/B/co3RpEZ+v9uJNSalIvM4v4lLwSu
R4Yd9E6GJrFWWaSrH+rYqPKr72wgbP3cIaGRxQkxdfH4SYbzSV5J7BN+85yf
Dd1bHh32neICsjWlknhUMdUqh1sQ3ScTAcpG2py+QwV8B4oh7pIQRmnbd+Dv
jrshA1CepJg4ueTC1H1YiR5/Y/K0HKTBdvd4CmDyNjQVyu7p8B9oPzhrIfPt
4JlVM5YygXsM+RoXG/1fw84CWPbNLbobXo2TdwcH5qvH4lk+9k8ixfop+E7o
79ISovTJns2Irv6rRXbVelJtqrgzcZWsrMtFMPFTPghH3f6q4wykyszT9cnA
rXny+eMzD2w9/KzZbOpZd++4dFa4s+T+14lYA2VH3xKp6ft2PTD7n3lSmsRR
p+OiMAHxXcZEvPi3ROBf0260LahlacIY7jJfXUaQISw++3IBd/C6dz6cA8be
pDxcacB65Ic4P7rGBg5uvWGCiz71EQgP0kwS4+DV5A7ZVZIL2cT3Wq3I8qoc
//TPWT5O+VMh/Q3v8gU/2XXCqs5+cL9VqctkqBjHv/I4h4V2TYXdZQ5TbWza
EmCKZmP0PGPFHXD2I3nuHyl8m2YTpJxtOtx/Xm5eAk5eKHugZrRTeNFmycv+
uYh4I/Rso5uU8bfKj/bKngkqmoDv5r2f4+Eix3YDoX1QEzhZChhy+gVwpl1/
LBPZ7spfRhMMhfSokMRYzdeG0lazZckiZOP95LNTglDQL5SlMoYTFx+ZJ+kM
D6ZoLs2VDLh4niqBqBXVqdMWV9J1adaaK1+3bhOHzPEKP9RjmqqvlVfYSdmG
pZzGup4hBr6yFG14L4c/DwW2z0dtFT7tUMnOKMLN7VyMeN1zpzGqpUVz4aUp
MhZeCTmx7LMWkmNKphA3if7pvXNwEqi2FKGMWmf9hQgWm3kZA76wRZ6wYJpm
PPdpBR5w8YfdXT8BDz1vjmmhLUpFqz+Qkn4IAL5YRGt5Axm6yW37K67NNz71
RqA9DtNNVdfZWi/M2njqYbq7YXKSjxqhUQwyUYznkJd57ShKf8ZEm7WCng25
wqgjm/Xh3uZdTLcy6mzF1Sz/5gFsud3N0qOOvjqBYGmAw8Fp0l6JvGodchu2
tJPoP1BQ7nkI5tKGkMh0TseIHd6BlaO0roUbmlNYiD67GqF83WAwiQbvXQD1
RZstnxXexS9iDqKcZ8dJB92heoruMKtFIGFR6Xl+1m2HPluexb1IikG/2CmJ
INaM64E5SethLS2uuLgdWQZjN0KZACLzbmlD9sj9yT+hlpd6AfmjAkTdrGtb
R2yV+eMeU6CBrCHW0e35gWe+Mt4fHH+KUCSgaJirE4oVf2ecC3jyFE1Kmplq
xYHlQv3KlcB6lNp0nA3QFVJ+7k/dGXCO2bd1V/ZbDal3TTFZ6lfmZToy2sM4
lLxOfA7CrA0MqSnFeS95oUeeYc9azPtC3WrTyoG/W4bfgM/ephJ+YwUt+w1g
ZrCesN5Se0kTKkkjbszROKop1owXBgGfvXBB96uepYheEwzaSzOEz62bQ7Cw
Ql/3Z9eSfhQqJNnvVfSy+IFyllHTO/27wec7byVdpwA/sWsFrPhnja34MyWj
xAHFtOZ2wj0Ww1nQ8xPO6TRWhZXlDey7Ji1r4PLj7bRfKyfUNA7ZYchGKaHf
2C8I6Kophj3dBTAg09PthBvH4Ne/Bi63G/y5lOEaR38tiwRInpwhhgbmyBPi
BxsJrYUSylLhzWw7ALHzxVmjS6Hqs5V9I+t6Wc4FPaiYe9OQ0zINzUSmOYqI
do1hwfKQAnDDuGYPUxbkjd/cPyTvVWQikaZw4/h0PuYzfQGmgwlQpzMBd3mX
/LldHHidCEZiNeer1JcgngWez3qpcnItP3axFP3wJWYvH+3/EnCQSQ+hlhz1
vBdme21yj1em4GVwZzHys481vGyBj+iA211piPx9l6b7VswL2Eu/7DBxuO/Z
mMZAvNumUjvW7640JdMXtZQJh9Mbp0bqYA16+7spSgGoLrfVMnoLXfPsDzJJ
XUpvFoQYGUBOQZOQ8+ZFSrCx6DQuLBmSJZzWPR34enIW04G7e4+4cubaPfyV
I03Ge08H0rUY7xQ6bKPAsroP/tlJZ5+LII9jBFecgOd5Fu6ZU4UhU7tstrPB
O7u/Ye3OxoJ5VOOy/2I3in8ANERXJ+CMzUjB1ZgcpQEaNLsxGlC18B5qgZzd
9lfnYfNIZk8ca71iawVwPnluTP+2YihojzY6Z6stZFFAQdnf9v1GSdiwKm6Q
+9T2tG0+U/V1qduB9bMbQhBtYEjDnd5kKNnyzgImbc0J/Vrh4QsfVnOIY2WL
Bj2bE5wuV+zF9LoZy57KQ/ITHjILs7MBT3hOsrwI+8p8MYqHCx7zjz/rptvF
gr/XIXjUxS7/Cyd5O5huRTxSdAs3IxNiU5PHRqxpOGWzqVXGVavV/A1f78ZE
MSali5Z2B0YiOQ43/Kd9hFGNL5YyjMCUm2ol5qniHqWrf0gEkcrPUHzzLjk9
l8WwTm/4ZD9qJ6Wd7/UthV5hl2prs+DosMXosvAKiED6ktEEG2vAj2dwySGM
8WreQt0MsBNFciTNcB53bKPBA/OEIN6OHgm+gUtJqR0ZOi3gH6xjY+oMb9Ar
pCCr0JtSe0MOaiEsrm/PzyFSbTwvUqgSoANRDr5+BbSzdm66Gsf3eeYljyjK
KMRIj9ISEV3p1taL1ZkwOQoVPtZoyII07CFRzhHXMCGJN/9AV7iD40ciA7OD
Qu/udUVU7DrpkckwkmutkzzD8iWDA20zUDDtruwoNShzSTuTbXBfARRsVTQJ
m34Np28lHGxKvgo1YFL4roTqNLamXV0KHvnDMqPrjIQN0h6j0e3t9zJDyTWs
5EIWIZCuOBLYcnatrsFYOc4xUHTIbshUcwxXPedLHRpr0iFoWqCEGYUkHfOG
PzqJ0P9bqvmkZgpeDiwfjVmdFadEGaAk3jGOSDd5WRT8S0zOL82O7cFs7DQ3
GsutsVbFqk+KSw5pxeNK7XKVr+YoXvXggqPiCSK86FRRPHhSAWELEJKhkyVp
snhp+gdjxiII39VRaT/zn5KVTStEMujWUXhlMJNz27oOdXyryPzfHYKma2CP
vyfSOA34b/ALbewDe7wAjusEqojDugzOx/h3ooANoohL4mwlMiWRoFBarL9A
H6sHh+TGTz4qH59C47l4RmZsejbDOLx7JOt6xPFQKWA2XC51+8oX4gH4XfkY
RkU0swn13bmZXMroDC5XQ2V9qs/GdSetvQ58q4HW/bDRhT/04QGG98d+sg/8
bzUC6GfwzbjY6iRiuT51n696SaHyCwNYHJzImdgTvvZKktprvtHNEHqcSDba
f8VVYw/opp2b45J+UG1v2tzI3rAjtzgvYtHTHnj+zeQvnqiknpky/0iBQ9ao
tIu62D/HSvXjEFBB/j2FFzx3tf6E+QQ+9E+xO/rR9pppMaouOPhEDX+kk1jq
Yc3TTILBFK8Jkb3ls+3Ny2WiElL9rJxH0k8Sgd8+76PPnXbH494koFC0DkXG
zhV8aElSzUd+l0fZCktqKS4HxRXIwTbUrN3/Vo/B+c4Cr9577tvgQiHx43AW
KRj6nGY7l+8AocO0+rB0+jBFJ72Fw0X3e5tx/dfNq7kuao2rQlYsuoVVk0gp
PKF7eLJFdn2o7vVbj0m9qZaMPH0MVUsyi+CLzZo3M0B783thl+WuwgFc3REy
FYGPAK+Utas/RQp0gVoJIbLCkSHXLbkK/OzlkiqTy7s1loChX2Ayo+NW4SYT
mDMQxE2c4uZhu1p0V8x/coPPDXfu4HGKRbYsRZrdXuUJtoHHK+yBXBXV4TAC
cT8kUGHXL1cSm0BgCYnQRUTn8x8JMC4q2xTtDCBokK+7fVxNC8i/uedpg1oY
T1lrykrHlsflTNiR8ck7GaGOXXE1XLos4Lb0Y93whluhIiZLHQaZiEeCFMOT
4mRcV2xtUVMO7tP8WYjqMHs82oI4V1dulj72nhdVzCSKtgoNYPNvC+tVoXhy
gceGqDvDDlPMFGL8F3LAmj+moH7a5gv4faqU4tU7MP8zT1qNs6ggmtu0RB0a
MArt1mVVvg0zAVg4UpSHErvMCDvO7oZZnzogdpLbi6M/zfuWq8pr3azhwexQ
sr430E1Ikq6XTmabx6bEpWOacL/DdX7+4t7zG5GnQ1yBXDzY0zueKF5AsxLN
touCM1tCYja/ZbHdbWSffP0q+1/+g74Wm8CKvEbhOthpwSyiXIvX71OLMXnA
Q4G4+5rAVLyHiNNCbhn6ExgsCcnmSC+PCwzpAKq0K1ckM+iJjXSs6voufwfn
W3H1VrGRc0eLuHYvvB+1UFmF5XQykH7yxsOWAu7i7dTzLRzdOINryj5gLyqt
s34E3rwpRpKTL98lpGCU15trOnukQEdWGiChwxFnzWnJ2rv19wLUUJ+4hxS4
IpPK87yCGHetTpSFOpfAPlZhhghErSzj4oMRt/CD/VL/RlDaaYZVdb26hINO
SryDTxT5bQtN0NKxtDyGCpWfLzZAa2iPT2p2GCWE/JRN+zOTmT43lu6QXUQX
i8LMhsIcNM+2o6f4RLM65mZ1KWrL1/xy9HduSBGLXBPZYSYQx99nlP1+om6F
3j6nisIa92sL7SizA6VNCuSKGSAqQbNY9zdmTiYVST7TJqXdOTN2HuqQxd1m
nhhM6pqeIS777MLwN/d7CPlE2+bv6Sp2hpmcKVW9d0twQDzcw7oA8Qr7jRw/
TNnNekE9aTlZ5ICRhP1eSIXv18gtkKkbseviZHsiRu/0zfzpCX6sJCymSPZu
mXX5NSWJc+w+GhmnzUX+b8ez7ISsqcQyZcNGD7RsO9iOTJwJDy6FZA6eq2IK
Rt7Cle+3byuleI0S/PY5UzDQK0QMIKZ58WRwOCstZPIXyQrcwbNT49cv7M0U
/5aQQADaooZvjf87xszVf9e0D+H/kx5c8Om4YtxCJBjMONHEwVcb7wX6l3Wl
LzWpMu63HdKhQzhqloJ/aKJtPLkK58WPU5mSxtXuqNZh8L/XNoLkQHrpqrfC
FpCbf/ZXgkAU3Qmq4eeMDtj8YY73zYRvWXghsaAOUnaGHbdaXMeOiGqXIi/1
H1R/3AxAO4jwWqvSWmxkkvElWA3m8RBa5ilXrEnVp2qq6yJ05VBvoaznAuWV
a4wg5hW/zjfhJ8VCmxcXF8KWJnWe5ZHDAzt0y+k2kGSRZSMxYXdNyDimLvP/
vYrb6F5A6c743BJ3pAKTg4XcLMo9/Bbgvntgv5HsEHUXTlgVvFcMx1gLwa7M
MQWm15hZSXc1HNO1HyjB6JZqcy3vvoWiKxj/Dhg10FfiV1IlVMw346kxxDZk
0Clmt9HBUU9p2IhfpYIaRDbbtadzzXoHCZRQlWbDnYVkf9bJAJ7Kog0aBYxv
hNOV38jtzuFzTwZAvU/eW7XxeGNBkd4Wsjz7XRPdosLxcLiFwoehNlB0qRfB
Ek+G99tJgltGNvkUPPBYocIJIpwHETEBy9mNM1NbRKl1wBfvEdmxFgRy4nNJ
uQQ97H5EJHokCtJwM18zQDI8+EO2AbX2S9PRLDHnf6ZNS7LJxFVIp+UtCT82
MUDWqHJjesBrIqas+imKDLAnfjrSU83S9KrR0F2G4JXUpdYl3vLwHhpsBWeG
eQ6oN+42cY1nixGBKA9n/rLkI05hsJGgw/GiBglgAjejKCVWgad8zC33U2wb
Z93UM8OP33gT5GGJMmqSBR1oOUnv2PEypFVP25DwjuHiprdvhJ1378FaK3gH
tTRLbqn+aWylAa2K5Be4//TFjelDBU0yAjDDd5gPg3mDo+//VE0ST7je7LQ+
4fEc7dwcotFVAW5tctkAae0jabhtpA3NriuxGg//paHcNOU4TN0W5YQiyLSO
s+LP4IP69uQNCKRU/Pihi84nJbyYPY4jLE3OR+HKpZs7TTI2/ULx5xBN8fM9
rHSqQVFm3RnP4gja4veFsvHK5vwRG8qtNVYOr8b+Q3pVWmmCYNbuhdaVMwf5
rOU+l3mGWinl9JFFoNS8QBSEAbQEcJDenxc/Eq9Lom9p9Pl6XkVg9vpmmBbM
IPh0nAhEtoBjD2sQvYsSQfWzo0aIN4GdXxhQcyasBlJA33PzpsCYdGp+3G2x
iu+0lcJ0YK2XdJrqU6XgmSu35B+RvPoKNXJcOq19j6sCTIPPfFNbOazGTy3b
5/VlmjQenrpkSsEKxljiBs9o0KOWsL9YDKudY8TCkHU5jUZH+ZI1uE5rzqqD
iX94dg2S8kXeVm28CI6nbM3vsp0tcyrdrlz2je4aoo+XO93rWoLECtcoBJX8
ElUe7VzXLrnTbTH6ChFs7hvk0/ZvHEAZdxTugjvfx19GEb/fEO0iAkWqJHIC
j8QxeMD+noSs+REHtah76f+F/HfupiPc2MFF6EgiA+dkiGgxvs5yOrB9F/ym
M3luz14S7ydeZnrYUEaaF9BAJ+OuRp3wGh655U4/VaMzeTuPVQ5YkEamAfqX
tmCYs96bXeOGtU+1rXiMT4YZ5uxzpNyGohk1JqNlP66CVVRASiJDV7REWZIj
hcvlN9Yi1rXV9HhAiGdHZ2VgctE7sl47VyovhDuGzpiLcamsAe8zgru/W5xi
p5Tk7TkmHObX5/migmqXdlvUmKC1xcaTDixaSAdzs9rsD89BC55pKcM+E1Sp
Z0SKMgoIXuykTLPZGvbuEvq6cq65J3U5Wq/eQB/mS9ccAHa0YdsDebJmLGmH
dy7K0/wwlMk/4IpRw634lwGLLAckkCwDUTULT8B/CkQVW734zvmtF4xPqCM4
kjF7HLBFQkMCkVTkeM5fudwhBbplXMg8nurrm5ear15FYlGOltzyR0Ythd4o
AKhmKMcr8ejDf4qodVeU8pFOUNeL99IlHSLSpFvC8N8Yz5Bo6Rt27YbOVXcw
e/6SrUm3oZJfbqFdT+IoHly2ia8MktSs82GiNT1vqtsboXymAhuYmYOs2EJ0
B62dbnDugZYjUPcFCAkZJAD0qRrTqfpV7bjAVI7N81wNGvFBPgy+INros3ib
jhL4pwRnoC0D8fpB/058fN9NgfOFFKN0AJGeKDhT2EDRfYIjLOl/rxRgDwt1
V9jdy/kC+UErwoqMt/5McafEV+HlUDqj4YZr+9Nwj8aCv+A+MyAhsQLTgW5Y
uxVRuzG7jVDB79jSu7CT2bzXhIpJsJQmE4QuUp2Z8c3LMvgdQNF67u/oGNSi
RtgGfmt4Hvk1TTKeskZAvrmCc7Hzj7Haqv6CqKP5b59Wk7m886BaaCqj8nPg
QU12coBMb7ma+nceQmb7pYrKiDIEy79ufjUztgoEEZVZkbEWidJPFQR/1rbB
rQOQNS+UBNQQich26Lx3dx2p8q4WnjZS33WwaATmI0nTxHPv1ak1rEBUDpKM
yOPBSX2bzmnbDJvwBaHYP4qtPZ9p19Y2UTej/uPzNwy0aLY6tOjYRGzpIGk0
7EoMVb72fePGAiKUSrE73+54f8v7W/RXN9La5Pguew5LnhnKNdIkPQeWYDd4
p6RCcDShYAiiubT27x1Gs50fqwiHAr2A1GfQh0GON7q5SsSEZitLgU3YXkDr
8MhwQ7P/MFy0yD7DJgw47BZ+fFQdSLQoigu4OhACrYeZYflWlZ356uORK7Xm
o8xIUHhEmP70hWlLEOXg9y6S2aPeWS5RKuzjycUxjDhuh4w6zYRA5qXpUbav
eL3XV+u1MZAP2ivvNtvB8zKvAk36NSq8Q4i6PZyrmsBSvkjTjudW/ag2albF
EdX75dqW5o4LuAU8NHe0pcyHrySbKksUCquj4V9vTFHGVB5AMAGR7QTS1zZA
hcvUbh9UJmF00xhoXsiRU06UZgFIMxTfaMCyoV8R5ItLVZPbJ0Cak5hb56D2
oy92xOJqZvYAA6iHZ6/TeNOnX4+W9YmfN8xqOLNzWi3v53HKjpZZMH/g6vDS
w1Kn4RJinqbXdDC87trSwNMSn2pnOicQJFEqVySCSOlwxoA/giF+V9y2FiNP
AMJBv33ba4JXdSHyJRorYlz4V4D8WT2joHMXHOlha/6YBugIbJ3DY2JhEQdT
gzdBsOg/7ntdxpV0hryl+02U6OnZgcrqIiJydLQ2Nr57Tj0EEdJfsp/DMxE4
TpSyZguz2blG25ABlZepULu03A5u4bhMfB5QAqC+f1kPyyaO64wV7IhIBC2v
tFfSa1ij/GdjC7t23SrDD2W5Ia0BBUTXrI6eK6XOwdf6i3VLtnx78yPnX1TK
yXMHTnhc3YhXrG8WMMI8LIxWUAsrFkmLqfD9vdKYQW2JMrIdPJrehWLfrovP
qWx2StmCqo4ASFVRzfK3ehsJIg1TiCLUqWsiM9hd6R5jwP7xQu6ZcYlhwUi6
BvQ16aYRanGW+4XU8pasTlq2+wwHlb+XA208k4Ziw0Gyk9OBkZCbztBgXsRu
j1CbndKs/iYnsNnU3pXU0XrPamNYLxIZo/mLBtSLRqutRuFoosCxIbnNaoNs
2kpELpp307x/qJsLWsY/qf7G1BEA8Pasp/Xl8CNGR2DDA6ZrRiGqBQWbAn2U
Q7SZVvWglA3RLmnr2SAZWh6QvjbeZ7qRT376EFpQSUQB5K1wCG3LDtVt/2dI
i/6h4MgwdnavovBy/sg4ID506V8g/Fl3tsp0aNUjUrXLe+zDcnxwMcbty/LJ
jlVJ2aAar5ylJivBAFxpck0eS8OsC/RvlcUHY4gtPiG6VJL8CammfHxq/LRL
oJCCdY9BX2onC0drzkVmUwZCWG4Sn/4L8w/sB7qK5KJUEf8NLVquT4gG0sUP
fESazB0wE2+3WlQdSIMAnS1ERJrVdDwr06m7iSxfTFjNAocUzU0tpymEHvfT
3risqEy9ThLePsUPxcOKBGFuLC5iprfAj1PgYpG6XSrCZUtcboERqHR2YRSN
3vozyP9IM7X/E48kfmUiQWdev7wOElbaP/BjoVX0mhsNnzA/FyZSXepWZ0F9
hf0OFMpKInumrmpvIQijJzeCHC3+BU1swGt/2UN4+Lp8WcxisUPGPSKNl0nc
0uHEFhH3uE2qzTKLrRLt/Rs9XJVInuFeWfc8L5T4rYSfa+qe8b1qskKZlJqs
/IqbpXYrfvCFQocHeyaBDRUEoCYbXZ5em1ZPj80HAPq6q+b/Aljwp2l/PweE
vjds9TLkew3Ju1BaOuobyshBYc9vTdZyLdfGVVJvFj8uq5sV3wsR997tUNlz
Qox84tQjEd+zztR8Yh97ksi8ZAdxCws6E4LjjoAhuXXXPQSUc45GHrKXVe3k
dwvFsYiiLU8xzZIYvnJ5qzN91Z7mzkLHbRSidSd/yABxX7LCdmpT2tlMdXyQ
pBmQOKU1OAL7gPlk0K/qDPduU8QUZ8LYkZXopvfD1tXEH+y2JDAkWri7r+qy
JwGBd/6V7IGvUJScUb0WYMutrvHcSb4v/Qx1ilqJR3sZ6JYXT5xcp8mspzRx
Ts0wZ31jNE1N04iQo0lCOoh2QJ3iMy+S6z1tcpy2eRUZFmxVQgrUTTbeZSh+
qvtdigMZooAo1Hk5sNlDhtvRwEf+fpHmDGmQUjE7pOIOSpq1ux47bDcxR3Nw
TbvS7ngOxLykpSZeNFHuNHamupdoukWOLJJp6ZHBi5EM3SSR6IV0/uI2DfJd
Lw6rZrn7pNJz4uE1dJ4K13KE4/ufILXM+2Mb18FaDH6XoJvPyRWoNOhBAjmc
HLxm3q7jlfQZilHWKeRbFuMYa3DdfZ8Ty7MW8txYsFJAO79vUwql2kt3ljEv
WpXQp0uBTmvOkVUDRiFdl/yPVR7/5DB3VV5bS6M/YYZ1wMH7r9wjpXi0axEP
cw+1Vc+/4l+b+HEMO97KTeVunaQQeCMbGvf4yqUQR6sAC/2+s9xetxk9eh7O
Dh0KOgcDjCHm9EQFvYZgzXcLoxT8+OVr/ayA8j+9+dMjJNX+9jG0Lt+Zaz2J
WrWISbpQv9hUTTuUPBcq2ijl1iTrO1XuidDO2GYnxce74T6H4yCHhItpA+db
rTuHMVggoMly7xfdNkKaxobAN8rlDkqAggqb06N32tGHUC1T91YQnqazEyGt
4jaxDGmdygGZ2tG+7EJK4OYjoAyr5w++lTDxRfmCy8JjldUOFgUCryl+qRbs
aI0TnJwta08nxHZctSsqtybH9Uki6vAJI0wRn4HhE6xLk8vYk1odIDBtVBUP
QeEolA466zIcRafDOPMo/L8lLRVDrHlfzSkor9xlnb7vqe0o6YHNRoPophfI
045ONIdladLbitp1Lsx28YKN9mAWCWFx2OhjdkZRYmwrDl93rtk2IrJbPpfT
gEmdPHxF0Xe+sYnuj6iF96S0R3etpOJG+eS/M7HrGvc1AfqCvQfdWElBIbh1
VXpGVzEP5Lutrrmyav/MVWMB8H9gDvGeTW1QtpJhEibGE4wAlFbDLsbEALjt
StggThCzTZn6jGLiMTW+25dBo/zIOa96SajsUQ8FfCFgodCUiGX0TjJplOs6
EptQ/CMbYCsNsXwj5jC37JNNbf06PrNA30X+pYOhQckYt80psA3xeF7eIDR4
Nn4RN7wzVZsxbZ6XM36C4/8EGLN8mBbDrEBAEVnZ/jNVbJuRrasb0kxq17Hc
uv5f9BZ0P17ZTlle/jTxztDALGefw/Mk8WBlrIJEKvvAJ9QRdGZ5GgIVgKPY
lit6apNUF/lMrAZkRvuz9vpFGKTD/4NMGqXCuUq+i8UXrwOi/y5ki3BoZKPM
6W7KGDZjsaf7bOYZszWhyFccL5VKuzlSn5sfGEWRklCZoBDF0TxtckCNwA6y
dLvX4vMQmZjOW3n1g1wnX60lAp5WI+b0WCSeo6VwhrdOmrOzhzQ9EiVJBnaf
drwvPC7rUDowlxzZXAlW7A/xAgkVPHc6UaEN1bCjUxL9gjbkkYR1vSoaXQ70
PUchhq5LfbBS4n02WOqB3ZdF1/gEPJtOREPgW8khFIqyAHn/PeFSrF0eFijH
UCQaybci/vYNAPWNRuD6JkhkXsyrvf2XHwt0AOXJIrfp/cU1J0X+CMBKxIIr
PjpWF5A4ZagAPE3cbhZRf4ubMGXv/aoziQXmYtQxIZJ5P2T9utyxc34QRpCi
i7ZSsPWZrNWu0M3bO2uwiqL/WqB9M7trDtWy0PJSwjUYxoeOpaJiH8ap20dB
Su90V+MJNPrfEETCAOT7SQ9gPY2z813wohlXY6pr6MQ4n/oTGrxTCzL5Augq
VXsMC7ttfBXNcQzG7EB3XaqcKhK/muPZ/brRKNUU5H1fIF8O3r1FqUIpdqOc
rLXDIdpkfXmrSLakbVr4tN8obnSJLdQOEzcZsgb/0FpdN48MAdA4SnSNq+A/
laktK/H6nVx621A8IKgFYm2CiwYAn6rebwdVymqlyNHqb4ZNaqNB2w6aCF8R
6aflhryX23K3pV4dJi10mTb9P5NzM1GSojSkfgJKi3TfL/lvLiiPwh2E9biZ
mEBzQ/aPNSbBYZhziZnqwGKOTW0kZjmMYmTYvIcWH4iKC1K6kEBVFCps27GO
r7Qwz1l0eMBaTTQ4wEAEd/LanQX5K3V8KNA/DaVASHNTBGE68ApPO5XRTqgi
YOaB0ENFFhiNDaCZ7vvisNQnnVVvLh2RPKYjGmakj0+dzjhalIaPB63n0Jba
a1rKQFo66nVgTw5vIMD/3aKKONy84RpjH9+L77qM6StVLSnhbcG9Dzz0T8QD
KlW2d60W5Mz/Q+++MVW3QHQ/YkpyURVdQ4F8P7eJGEffE4YkmvfBX2tjlnlf
Bb4q+RZTvfuQjEwC8W/TNS7B/Cay11/4SEk4szbwX6ZH4mzy2d5cXFiFhw1q
Ja6NYozoxaMdw7EfOyf23fZTvK8cFqWqre2/gwYOmYrmTwoAkd0o3Pjgtzom
I69o204T7ABbNW8kVIIc9PIUFTTfzI/Y0/md8bL5dQvv7pCinDscS1pwmxmE
Ml42UqtSUsSWGnrhwszDHM7lAl3qNuJmHi2vGcoWo6D/ghI/H6a/jepw1nG0
q0JIbDNkBBJN10cmAtyMEW+0UE0ovvdToeztL2qIbGnnrxF6KfDceGynjQF4
i59dcdHv/kGrKmKcm0vDUl+nf25qi4hjZHdQicimL48jEtFpPRghgPnVGMJH
v/AX+iNNJ7VIWknEERgNMAZwqNHX9XUcx5X/SEeU7Oecj4/sxz3WSz03u1wj
xUhkn/B6fWkqSX888hmnPMrTP4vY/28Kp+Z+JOml/F7V6PqKe+fr87s+OhY0
R6uZxooLgThoWqesZzkTFLIjGCU4PF0tTjhwgesdV8rmQih0AnFg7YaA7qwv
TUKY++7LlvApxBjV/bDNb2L82HHRUWzogCp7CsFlVW8o5TQKVGUc+9YQ42yp
dDQAvdoc0b7giB17h+VQZV0DiLJAPHtu5w75OVxtFPvKrH0WZttPHSKaeKzt
1R7SHHLzcpi44zUZCeD95Fcto3z1oVBIWaC0vaUn1VbP2l0ISD8uji+T3ngO
FenSgH/yoSio7bo62/wMnM1sDgZ0i+0VrC88SIYhGxgsDgxxhsDJNqkSJmNx
N8ytnZoMe/Ww7o9HqygwCEckZrMwynjSqI6diXRUVi2XWHNYnA50vN1DtSbV
hD94nLnSMiXXVDOSNHR7UxTHYYl0lBzDtg0lwQKBTaULUf93foJuYwW+v9FH
mQAHN0sJUlOUZ4O7S+ogQeLIKXAat4iSGlg40lDu97UIe0q18KhybvOdm9Pi
0ee2CNxKiSoN2TJ29f3J8umJZUoaQIg/DcJjxitpFRn+Ywtd2uKyB7vpIAs5
s8qWdhJaad0b9053CduDq5QJYDLls3oeeP5vB418lLTMsPOnOIhzKXvJIdel
NuzHhlkTbX+5j903+3xWN57tLBnBzkxuNIJVgSNixFjAabXzmdZ8NvyyqA/D
wuzO9jOa7brqWssGmtDKSvLALpG7THLFHSpDMP0MeEVxO78xOBKA9KCFXwUg
HBliySVd06ua7sGfBmlfolrr5+gr6ILz+ntqHf6JDaca+wpo2w8rQTVJR0yV
v81769Qx5vMO+pVzOzXpOnPl5QzxH4bXk78NTFZCiS638VyWGn174c3gjDOJ
2Vsji3KYgZX690pWm3OXteq1xcFj4m7Y824r2Hpufqd3CsZex+qyqlbpeNSP
yasFShy+Zy13li3BM0BnVamfQ7KqZ4iRAPouoZy37nIx1nFCPjktyalb2jBC
18dsGa5V+y/ZafsMQlPkuVw5+IU6EDegOgbRrA4b3jysMlY84Rmk/W2OEyYj
LHGHL7FMHk4cGjzNYnh26G94NZnH+YtAQ0ON99famvmNIo94jvXwo32EygmE
neB2j+oNqoDKUbQnKbhyI2ndXIJsj/l37dPuN0/p2CU4SehR+xWzDMkDuEVJ
SmOdT9CPZQNOQdf3uN0v73Z+V22bLdvkyxg8x3QZ2GMjIvkFVxrUDv9lkpqb
qgBV54EHFV5WxkDQx41NmR1brT1N7OHLqiSCc+TFbDhyqKrUWuG8D+byKA5k
M4IPXT6FdAdh00CYQiC9fuz7TvHbP3igdAWt/UtCMPjPusJvAByegBgxBY+w
Sj7CMDXgy92lwcI3Ny7tET5LHnietRQJY9zl679RtBqhzqA8ly/LCHOONGGb
hdNMh0J0uswRloCkYcEn8iPncrdUGpDBd6FFCcmDj3WwZFjLER30dHQWRQNl
fm/nWdIoijEFbTMKm2S9YarpMrjFAG6Pi6PE+CFVA5mdfoXSalVI8CbSrM0V
Dlm9I82QirNMkadK2jY0WkdwFJoDIzc1sjHwyRKrl2PP0XEBuBYGAUe6hk74
SA52SdoCPzXa7pJbcpeo6rT16I7sD4fcG6nmCx1Kf5tnikHWIcK2G5lmAZ7a
ER2asWyHKL4qOQS9IRUTqeDWfMiJRpEwyJCMUIiVlkVTnS+6vgXOpl24gcwc
yqmp1+PnBgiUzKVNFUOh/QY64AdQ5E0LDJua9HagEEbaSPt6DJOhwHhZUPrL
ZYHfg4s2ccSe7bunz/cLb4NjVJFkmlp0BGtOEaSDKrxmYowGLZL7ygSOsmkA
QD8mOMpyjlPUsSLT23Lp7vp2gsgWipvP/nYyXKRRekeykvYzpdwyQcURHZp4
LOQ06fhfjIc6zJiuXQ3/lHheo+d05cpG96Av+snp01tI/GZpXRbmN+VmWBSr
i0CQy8oFOy1zcYqhcZwSO3eQQJ6TyCxfpFI2TLlKvEeuNhMFZ73tI76REMgh
UKCUsxr5FvNrIDRDMaAtP0jM+qVh+IxT1BY58s75Vkp44vk0i02Ydy3mLFXt
AX5U4fXhlTLd7jt12baA2QCVTs4MtHWKZXjRvsmsP0IMbZkUjQY7pfFstvvs
65009dbkIMiUhzL5XCbvsRDY3VPihhRHb1CqEJsdLKW1p/yHEjLaGJ9p9hx+
z6IieH4611mAFDXBfBCex+mF3hoZ8v54hqks2NAfUlGRPtXGF122V2vJqXcQ
8RrtBF1KVbxq82cruV1FNGJiLE+FztIYhmbbRu8JsoXJY0iw8UFDFC0ke/y+
UhD6VGisFfJawWGW5Cy61sTVI74ORXMhaMLkzSY1De1xJlxJ3Sl+jkkR6GXP
ZTBJe0t45B2CfEsAmpFrrDxRfOFaf3dvn808fryNGyOI16yQDMqIngY6yDJ9
symakYm+ZVSSm4AXfrwku4DD88TAGxPTZo8VeckU41b6W5olTHwip4V/fZzV
tBaehgeKe8RVE3hoXVSUvWaPAfAzW0/Oma9QVb/c2WomfUFOhBPzcoyIL9Zv
5dGWIkeQ2GSwQFzufKEhbbspXHCr0Udjd544enPGFjS8wIsYLruEnoOLNl20
ryICej7aHsmdu8O6Eu0L1+0mPUFXR73Kq4pn296Rvn03TS413tPT+iRljb7E
ZRzKF/akwSXEmDv9UWuZ3EUQGipGL2cL5MbpFHCCO+fouFo/thObZ+cHwc3S
Tpmqzj8dHhcS9GW+IbSEtkKDPV6lzzd84KMeG27mEoylqszececCp7Z7pqpN
+8/NNESSkRYeAdSrrh5MPrK9AWGr3itM1uhXL+/zjeJ7Fh6xEmgeaoJs1141
09/D7s29lCZlAFw13OtutNePsEfKkRplFXDKHexYO8eQoE5/1DROANexgwJ6
jet7MQO88IyDLhsTxgoC7HiUmjvzrPEFPCrp9GlxC4oztAmXSwzf26HD2jZ8
BpF+w5NP/kvCOohO8rJaMtcwrg9UjhqUxWomG4tQmnbjAjfkXUOKCK3I4/uQ
Sf2dwPVEcis1mimlb/ZuYg90Mqtk9S0HpLIuMm/3NaIur3LIf9UFmH8SO45T
sGTbYvrlgcr8P+f+mNfkuk8c3G44OJ8FhB7dN1jQkpypc0qa8tvmj9eflaIw
uxPi2HHJBfn7NNtHQz/NBGzSIPAeyodSmPDO8mh++M5VtnNcHNM57x4JsXgG
r5MPxApf73ZMbqBat0e9vOBhtBR9leJ+AGVZBMBH3WSeIP9jaqo9YUB6xGZw
PtYqQHJaRK9kXP988ixnrqGeLniG4Unjjfhx4GXza2pNB4rzexsDKAH2xcOv
3Gmwft6j5+Y3+IES7ntm48vZuMBA0xeOI9yLQlCjz8/hrLFLc7yp5M7eyoDW
5zcYocJyWDukwZrKp2RKlnJ0VoVf+xXk+OSb3Qgi3dBaMvzRvMyejrFqEgWD
reYKOg3fudPOQ4Rc9ATbrRcmuLa9UCVEIkrCRsLeyDzeIc2rqzFrAfoBrjbC
JvtNF7a30Szr7T7S7NmptUEuVi3C3twKoHjCYG1O8znrwDhv2TbTsVBOLKgY
F+OJNSNSJ317U1JNQ0c2io6p+FeKzB0ZCXe5Ze8wtvXU0Q6M3PvPn1t7JYhH
U3tF2RyYTooOpyxPt11rSae6ouYwVwFD3ojAdHWT66wKa8HH+tQ8URi//O5V
ed3rKcFHBgGEkvna308fpplnSOlh5ufpDVnzg88hwqjQ+flLITAWhVOfQvaf
IYsk0gWT0KqEy1ptxQX3j0HT6Iui2gSKtzDX3TV9grCygsH/DMasiv6GOTHX
beBHVSQbiJdaSDMGNXFWum2ijaRqV53GKO393NMbw5MwrdL9t6bKCj5rGfsa
D1pkUsUajBRQF9hdVGNRNIqhrUa87bTriD5HRoFrn/iU9mKysooRVKexYdBq
JDJZ7OId3w54qLinUh/9U5acv6yFVpyJSyKLGFkXIWfsDrdoUSAxGVYZBiUH
b8+xYPvG5WyxTRYvs3jUG4BcHPvksxJHuhaQMdk8pHBgc9IPGThCrgYVWdCJ
45cJhs8ixv3PWrEm0NTNFeaMxRxDy+hZmeitNNsRyHMjCOKz8SOmbE91fJOI
lpNxDXq507Bevvn+dTmxk7X9D89qNKFXET/nIf6nGimDVspbseWL7u4h/GIn
wk6pTcuphSV+TwlrtczdDGEWtfqHaNuflK1ng9Wt8MLEAqkR1FczD9Oetth+
aUXdvioSxS+mSv8ySOr4Ddk82vJJdekK1EGR2N3mxnsLUreUVMaPhmsjgutD
BMdEbEQnF8phtI64yq2LTanG6HQvcjHqlT3aH5QosCFsIjXQ6vN4OwmmqfkK
QmP7r1MGDmQomO62zyxwrcMvITzRGE3yfcoLHNm/POPpzpOWLAXQ1gE1yRkm
mgU+u7acJORtjixtS0TU54ccfiO1T3nKAQkGTvy2U48BDH0iBO8N+PAoYv3g
Hum/5rjsGwoD/3aQ3Ita2qCgEjRmnlNTdaJRbDSXPuH4W8XV2sRAYmNkYv71
nCOJ2/hggt0s5UksH3ZxpqPWVmItuVR8D/2P6Rn/696mTm48EC5DdmVnRRVP
4kwhH9N3FeycrXgOgSB4LoU7XpRM0s5CvTJ0rUnIi6q/m7Pyl60EoEVHK0/T
fqB2dWchEtlweD//uNQtIzPpcTocd4MtGhaBcZyjoKlYg8+9FWlgrSAxxGmZ
LUsPvvHt7kr6qngPEohikWbZ7nE2m7lfg/yd4gmjp1udi3fDgDfW3kNLYA9V
MN2p2r9/51IiCoMlx3Mc7bx+h88VqWCASlcAS85Pe0mPgSGIO+S0fIL9B4oH
eI354xVCgaVmEs4vADDyMaSpBVtbBRowyDkYRIywHzFkRFao0+UzwG8uifBB
hCJ1b23dpNBMHvEVJ/LdTFJZ+QQmgeWyC6LFzox+512kFIwo/kp7epD7St9A
gnD8a1rtmlk2/VPr6eUQP96B6NbxdB2QdJiUkBAJt7hci8rbfyrZ6fjWwZ65
oTWeKPOvH9PuupB2sQPEpDIkdyzrSVrYrBwjrSirN3HTv9hXp2HZbjxE7zcH
r1cOv/zPAtZjlG7tY0MnkKqSoi7kk592+tBTXH6yerRuFceihb7LR91a6TRI
OxVq375JXT2xsWKJzQpmyMtysju0qodSjAxaBG81caAjoAtdZ2nDBE+2Q1I5
iukd4NHH/HNTP/p70rEwWkPp9RNaqFnaeYnd2kDtVGFp9MlAbw9inxBJZ4Iz
MUI3D02Y8dHGK3j2R3CXluK+upEFi0PXPATs4S4XWoeEdM7dSXs3huvPnOIQ
bd32F1znutd6Wjn+xU4uvelxeaT0LrCJD0qb+W8vdZ0B19CvxaaeZHVBoBeJ
B0+nOmZQjg+Z6Y+K2GZQljEmIcjlPYWMJaj0jI5nHleTdHy+cjZZBCCVQy3g
uv0wEl46pTrHlJdiDtdADCroOgj6ubMRJUGTAjNsmvhSyXNKripnrznNG8az
OEDg8/h48mi5jcDa85I49OgNMcIt2o6/FpAh7dMGrC2S+IoCH+zx0wJEXCzd
g5w9tw00dgqTm3vt+OAdiIKF051sOJTcx9n9d0of/yCNbNjnjD2x361MEevy
STYN35PJpH8wyEtoC2ZuOy5cZ+7qMAQRa1BoeTaa8mO9dMcfJH2M+VKJKl30
ui670OldLKY1W9MGycK1X5TkEGKhPwqEDH4/S03uMXK32Vo0eWteh5BhTcKm
vhM6mzfr0ncgoKg7O1jeazqWFzV7Cxq+AkYW3DX/jM0+jtWcb9myrwdpT+U6
qfCkRU6aGFnobHq6YobSthX33rJrG8QGtC9gfRO2dEqIVnU3sWIHP1vh/0ZB
ms7L/Z1v6/z3yAt3FxCtWmVA4hjysd2XyMNMoWMr3GTyhCiRLFyiLqjoBvHg
AgSWujVdiddoeSL5J3TiUSMoK7jtbH5/OtvkY/lpmyISnUIqPl6VXE97W2yz
gs4B2bBKStUYvQRFQQ8duwOu57PkOpKfqo0eOodOKSLxVd8QOcLUw0q2JliP
F9OsmOJkim6ycRNyzi07tCdUd/trfFFY+jurCjuv07aoS5LLEjL04Fk1L13O
0PNHJFxYnLyyc8Et/O4O09xYZ1TKicR2vaIzdWm8bsApPfaYXkUw/HGL+sbq
7iYb/t/pbEc088SHYoODvYXGo2208PqWDIX4SKqcqOUYfXyqh4gZXt3oN6O2
aDX/umbuC48t0ggi6h1xpTHO7m1HsRTFfJ/ddHL7K1AeigqU99Yb3E0uRIyd
gH3iu2mRXRoeaRe1ZDDTwHZmf59AE3sEQCeNHJyIp+THIavQr6q9j0CljjmZ
670+RUo1mDEjP6OMetde+3Y4JYyfacvc5P//MwJwd9Ro2JVmj7w5KZoETdCL
74JC1dD6t+Zbhs57smVBhCs/Rx808FF0eRCFl+K8UMY6u7L0VL7qo55BlKJK
Y0BtebHU0WHzDaAhaJYA90GemZE+gV3hlYHR9OZ/ss1AwFY6wLo5ZdEBgpB5
sE/3F7OEmiarjjTM9XmU1i4dZdI16ckeu3w2Js+J65Ch7UNToTf0bubD7SvD
S5kmaoccYhTi1jzz21/9O6cFY5HCBlNruVsSSfGvhoh/538ovkjpxciBjiPp
eRBrZJbf8nREsCCVkhAgNg/GfdlM4VR2GC2SB9B7QB6TDssWZP1W8xzfm/22
aCH8usHZDe8j5oENGbpDsb4+kj6nlnIzMKs7GpPHxa6NveZKhEZa778Fmh/e
ZMeDUGkJFMDmig3PVa80OuqynichZ17wnJhmbwRqREceQ+XIQO9vP564Hu5t
tXlpLxLAyMLDOSBLS9btgCE7K31dFJnzcc0rjPeHx6o+BY0DEwJVUIzW3M4u
b/+Hh96BcqU/9jLkeO27ds6wSJuz9ODkYpEopBXx/NeAuc3D1j6tpX/vadyq
xUl/1uE9u1wHI+hI0efUdzAu9pqq0wQHykonFIFdJ/FgQYL9Ne6xPNlxpTza
Y1HBR4ilwV97AR/IujhIsZM3dFtz0VC+6tphSMQvMC+dKC5Om7eJOOUa+dcs
kxqXCaLh2ah4SWwERNaU6C23bpgEJvLlOq9cGqBApeUyjBH0H+EDMdmvw+ZS
djFbLcXlokzAyh/ZkxIGF8maHpJJ17ZrTdlq9nZigeUtjBATqsX7SP+8kzn0
LYy7Kklk7p6wUipRJUSbHsN8NKY5KYNYckIJPuod5eSHgQppZqdWnLkn28QN
woLOAy8V/zlx0M98PwiIhmOjjiVt/0oknaEAyYpIHwD8gczvnffY4tEB0XVN
WQIbhRk7vjK/M1ZvVwdiXlVKDcJQyXxoc9T1JxU3BHLnZbLQ7zy0eO7yV6Uc
h2gqM7KEKvyEfUeXBnBQu2ARDpiO1vyJwVdW5+75Ya0LrZ/69v1cSp0w9Lz8
TiszCOC+O726fyZ1NZbKYDfmooSfdx25LC5O/Fn4jENpU3BdlfbdfH4UUN5L
5M55f+txWOZ1d6obekfH5vd6lsQQot7TqqiotJuOf5NUCOf+3hcCYqx/809P
ZUiiSNUC3pa1wTPeInRvhmW7f2Wzwu9go02v07VryiDESSti573/DDh8rSuN
GNPykI21I+NWK2CUgbrccIPuPx1Qaq+6a1lldKu8NxncaGgzMjkS8wrFgN2d
pWGW+vToQtNgQWGhSf/Sxj+R5XcvtlO3wrLItY+dqlQrhxe7vEtbTL17vY6v
U3iUI6MuhO/Gwhir2zKOcfVoL6H8m0rLRBRr00DRXi2zP9r7E/sF+wqBj8Qw
pK5TJ+Cvj+93CV7LSP1rgqcLv+9PacIFosI5aoIP637dnKyseH93qPBofov+
c4+C1ZpxxGroBOfo++Xg3b0B/JdDE5XuVehk/K80fTz9InFtSU9tz/uzsCRu
dqt8bcVcXgtmllY51r2VMVqq8hX4kyNUspw2+w9HFNwrM8rEAHosIbC/G7f2
ljyCagrOEbwdpdSzYd5zflXQEd0UHlasofQk33bmjEkuoT5YxLvIDxcwfbnl
sm8dQ9asFGVxZOV2pjFFMIUpaklHVPjXpRE3aOBoqqp4DL2kAF+w7M/sLWP9
oSeKovHRSQVuFPovqPyDThZX5IhjxHpUK1OUNC37PC2Go1do+y5nX2w7GvLV
1EcqiNEsDM4ulAtx6Pu2reOIPR7j2XyyoEYnQqKpkejO9rVxaXfFWbCT93PZ
+QU8kxWjtsMLIvjLBRL7C434eYdaxkXTB0dOz1elg1v/k+LjxE2x3pNYQY0c
zzJqtRPJ+29TvKBoJuT53xTAFJNQ+XKQ3nQFXfmKNFIxQqqoGHbr6QxWO2On
wQBEioWdIFZ7zmKsiNSyRbTYYABb47e6z444InHJGIuqrq5ecBJkidCtaXCD
6/FAuyXvYNaQ/tyu+Bh6jTp0h9q+QgDh3wRP4o1iAE55Q0N2+oCgxgDJ9zgb
5UxG3z3ydnoqWN/SNMbIzX/8TnACvjYqfhoOpygMyQigO27m5SpI8EYSwe+m
ACkc+O2yKbKMxxln6JVKs43IYTwhe1dzu+KlMSCzZNfeCTmGwR/HqlPHr+jD
ccw9QpC3FglWLHDIKLF/WPjovKd3HxHsBhXYPT43QMsVY5FJUEa8yhnyrH/k
06OhJyAqVK+oLWRoGKS+NTTCtpMYfUCtC/BKIlO6xyulcZjLb4ws8Qy8fSMK
BryQHfA8cN3sJmwhKJlNo1EKxnPl+CCkTx3cpGp2gUWz7pyGyOyhlC49jAzu
eQ3IWQSCk8ceFDGawtgasVrAnfMKeGZnruAvVM/gzlD6TqrJyOXH8ocB1YZv
r6VpBq1GXsM8FAFI3bFQcbK4UaprZQB4tSRoKfx9eQ815uSIJq9nVh2JLAPF
H4QHNcjBnfVswjierSS6ZDL+awFnxkKJFR57gxMgD+nha/nBUh7F4N343NoD
UKX2vMhBQS2+fWMNAetEd68d4FHA3cUcilMD1e1LzjuAo78XNUJuc/yvGaAf
Wiz479Ku4D/UhiydRE9arf6KZbbTgMWwyrg4TxR2UAo/qrzOvbdCQ0gMLfYg
fUrUXFLXbIXF4bn6R8xQEqdv9/LCIxONSpSe4pRR8q0Qxnrw8msIryo09XX8
wNyFi5Suok2ZjLCq4QwqBHTyWJ+UEDKBustL6OCBBRZD1O78rfLk/h+jF+W5
KjoposEPC1WutS3MgT2FWBO9FLkezMYou5VCsQ6/ZQR9Z9+U/A1VvLM+obqx
oHvUNYXXzIuBGCpQoN2Sx/+JPgUcKmZ96DJ+GhDttf9VoPvC44hJicsg5srK
YMbzEXILvT+AG5w2DqBagbsovwICxV4GB657genFnaYa1xlgLlaMrSEP0lhE
vAng6SkAB56gAbEBeS7g2jfGmruMt6Wt3/ePgyh01K2FwCoq5JxpHHpcM3b3
sHma+lm2Pdv94OGSXW1pWntFgW2iWAX3udAOoZA0n9SX9eWsQfENZK2sxwgI
O7Pkirc8Qg7z3PE3xsxCrb7FT/9hWHupiWa4VIvdK+JbCR3K0NQI2hyiIcGq
ih+VFIlANkddSved4xRLkxzamfqDMRzafhpuKyvNkinLMeFEfjPxMNfByxC0
nq8Y8goFNEwp9fpW4LO9p/b/5o3UzqC/qHLBXeg+DQSL+Sbu1PMrD/d0/bUG
D+tI/FuFzAqcjW4xDf2o2K/0CpRo8P88TwH47emTyZ4M/pItJpbDhfPVe582
MvuppD+GfnCvND7Buqql8uv9MYCumZ9Dt+gYp4U4DnIRFtAUZW126VVA0A6y
GfCWqG9vYGeTEZK7KXVAouNr7ipTpQaZo69Ievn3hdZmpHakBAjT0Z7Z2py+
ydt6YVSfE0Od8Qcg2RHvk/LlIRPQvTXJqSk9L8ywMLy9nzQsxQINggGtd0vZ
6Qk/2WFfgcxumiFGFwQCtPT7Hs57/2v16rdBhbBiMMsPgYkXMxP0iKb51QMS
dWaAQMyPd7/nh513Y9R3amr9e4+1SbNRzBuyt6ZBgBUS8wN565QuMj3DujII
4Ew/Ijp/+h3jubiFka1fWtJrVXOKfltqO/6x1Bx3JyCvPHHrgb3Hga9TAN99
7o9Ou4Ne94TgHJ3vJf0CEpu6nmqzPydncl/RxlmPVb3s/r8OPWLqYG8Dn2LT
oXwJYdS6HvxcAjYMQbtD1ahwXvxP9swQXB4/hrXsk3gHTquSHZ7k6IvY3sMi
n5Ue5RKCOcZLijg9ijkN1M2t5m1DEevxRAcmtfKB3wg+6biTn9JJeKuf1IKJ
aLCx5+ccA2pGYRPqHIRSMoVnjH/se91xJTgAM9bwhuNEHeiHkuQ+txx/ej3V
PRC9x7XOeuUmhtwRm9+85TyXYFIPH7KMjTPDM/flZqhmkIVJruh968yOujF7
fFYFVzPUa89EON3hp6ZonNl/Y7zfwDVc3kt7FYm0MTgsYZKkh2PYjfa42582
ChIGxjjo50rhQ/ndFJSvGjPXItwxVhZtsDRkd0jWIoCXQvYkWSgDWc+kjFcR
iYS4yf7VUAIgWEUPPpquReZduItuWTf1ndaA6mTcoFM/Vga8DWCWbaUJ8iFk
0jbEsKag01cjI4DAk35CS0+hSNO+B6iVuexpPpk16X8vzGWKEWH0XmUs2h7u
CJKoAeZLD5vLGmv0+rk8P5X2cc3rNwDV+Z/mGi0pqTcU9yGVcVuJ7InVG+/A
c0wt8KRNreAO7bAQM+WkU9s/WzXV8Iiv/x8brVO24sK9PrKxUohR5OZABgW1
2McI7vNg/igW0rdBnRFCpFOH9bw9a+LrR/5myozjX90u1WCy8rxd2jYTt3X6
u/cUMjX5rrRmyACnHDHZ0le3oFT13FkNHSfPrMr7Sxtyczt8caJ1PXn5M9lb
aOZ7mGfmpe2hIUaR+DXLUpnlqnEsMoGO9wa5bQa/K6+gB7hlzI/hB5cG2aJZ
xTHyedDOc+aVOT152KwFMJ4EcNam/vpDRXcgVXGsRe7VSXABB8fnbc4eMWg4
6+M+XlLDp2wRuUwyR0/eYv6xxckbNjS3j9Hki7YU0ueSFSi2Gxkd8XUqSlWc
3UzSDlFrvD7CQ8F+aCoeWd+PJm7u5ljNbToM5L9ytIoNFheFzePHuD2KQdkE
71GZ69IZ9youfDZlmZgsuXin9xHia+/VsEXQkQz2Ej9Erudzg/qspm8ISmNC
bK8QGmn0vB/nImR+WIBavm5D+jleN5SXHROIg1WpzXNXHwbv21wjqCi6XaWA
zMwwqSN6UFU6gTjRHwNbv/Y6qp83r/z7TZxe6zEKt2HEHLa7PmVXS947rkDU
76NzWnuzcOGtq6xZcunKsDL0HToNJnDZzZSUFvp0owGb6c2XvdxXwSNrMz1d
nA0zWNHvloriqOn6uTi1RFtWbB2/QcAyewDGR9h7Cm5sXiKVWshHxonzUY1o
rkcAAWBrPtwjYIvXaBSA04y7SdM4wUOQR58rJKchax4Qbh+PwUTPv4gj9pgn
nMezCKB3gSWk39NM+iY4jjU2VwnJTfJfNa470pkGKXkpTzrKy0J+Sbae3otX
rgnVBSWm6DOO2SaQuHeZvvIikY8v/Yd35UmK5xYi4bvgWs7NYAspDUJXjXti
3oGqD2ZSdabh4KD7SgZ+9qYMrBVZnd5gi0rkg8HqVFuehma4R66VOoEv6NO6
Vls8uImOZboufKPHUQsrhavqns47NC/KV2xMC8dnJiFxWoQ1328TmJ5+Ax0N
wWE13VqSlgPEpsT55b7/LFw469yFQYEq7cncRSIxXgGghTq9XGVr0s7GTxit
SzOFpUaCHZ2fcfVph+GqstdeIGmBDFhA81polpHW37aQV4n3luO+0habMepe
zoOL9lxHLq3VK72PDXPCh7d8+CTk+AcInk6CRS/S1zYxWHxNq93NnItrU1iS
cRY+3on8lkAIbO5cbA65rNtHfu1G3QDaIKmc1hQdoI33gRlrCMFQ7YCBQmKY
/Ziz41lPzhyyrTwdbhtZ7724dT6e/Jp2aBekqh5CK/cN6Z4ckir84KZ5pLHG
zkgkBrn02mNe1OhI7VH8IO6Jk9xsvuZq3UNmbKuI5qZFTrcfPIbt86Tztvxq
RxKUtu+YSw1EVn27wbOgQVaAgZZGTtuLoRvUgNMRcAMSx42rGfaNR1XT0TKB
Gaa5gSLdOJz2QtBg7leBtQ8ivPaZm1LYUYxNlyKpi0rA7VkiBgQKHHuhUcMN
FiNlY0iE7aTAgQc02JH/zeMq0pMiCIlsxbGGibe0FdY0bMOu2bsz9ILdcBPx
Nd1ba/vJ9Jek/eflyqC2wfJpgr/96n/jv5XzEx+e+QtNACv6ll7FV7HoIiCp
m9gW981LbrMJEzCxHQeF0ltr1Qg1yaoUq4+joDLPU0IF21YfvXWsubH1bP47
obKE7D5NQPWNOoRMv+xA7YIZM7jUuO7YQgjyK2zB/BrtiOukLIarjwaZ1x8L
BxI+KTSIZX3Ys9u1Ihp2JieuRh+2gH882eThxJjRAk115raJc4FYSrKMhYWE
hGKRZU6LIX0ltQPf6Gy1m4yaS1mxClDONRmpow+i9ufef2Gtpw0scnfH3jyJ
wv0c6y1mFSRFdr/muZ6Q78N0uIBGTOoRk7wdcOVfqic8nLDwVn2W6qXLVGm1
c3mfNPy/EjNLIaipD/uqoCQW3Xvu8CwJiDYkjVHWQ9JfrAtl0p/ttNN8eleI
YuUmOcGuMIBooKjek331ZPa1CaD3OGfqIcVE/CGV+6lhbisSygcEHZJGyznr
WLCjlQriiraNmpl2JVOES1NTjKg0/R5bmmmb2AQwpk7enEaNqSzYXMKVyu3J
ggRdj32XiXIJDGdpcMLTeIVFH8VA1jCJ8Lo4+kPgi5L2TX4Cgl7Re7Tsp0cj
3d1IRH+hpToy1G9XnVXuKUPtk2qwQ7MfKSO6R0sdxnD/7Ql0RM1y8Pe0cZLO
X1DeUNsNdnGyapu1VaMl7PU99Kl+PFeidbwFKWtSFp3hiG5Wfr3pqyRzf4od
VpzL2ygML9PqM3YyI5ZWgkkNrqyp6d0YRpUanMlew5ZfQMBDHdmDZ6KQdSPB
PNokGCYtcSra2U44+j6cU1bHpxC8m+LFYkkH+YX64/p+tG6Vmp/ry9cBgTd8
rBbAFpYNm5PK7/N3u7AnlFpo0HEc/rycX+O5I+lAQo7M007IpC3HyJ7LRPOH
cSq8XCngWHIRFi7mrz3ZxRP51osH1MjbSbS46sFdUhSg3ttTGbHYWEwuSKK4
xThOdvi3zcEydpxKiBi78lHsF0JG7n794rzhqyVkgQ9I4rsb8ipKl9c9HlBl
4lx5jUdVnNmWbpsL/196DDJUxTWSE7yxgXohKgC/s08vBSYp2rHzR43FHGd8
Dsb0oVCNCVq/txqhZ+gAgcujsnoJBKIE8zFG+isp1GDiR5Le9HXkZVHCn12f
EbhXndyn7CajNLk7XRzjDf+9DzWSgHcR/PTyXry02H5CxUJbDJfxKKyk4kEc
9JsUaxYgBj0+fdPZAejNpWcf1EVFsh1OHetlEtxv4Ol84xzlrdNl60h2cwU+
8c23txn0irITGyR8KHk8cY/6Iz2T24Ee5yd+oxmT6qPi38OCw6hiKRNiXXKq
IpIr1mbiHMJ7Dyf/vbzAS9XBeum9DOurHVWJ3ilGFJfnmh7xwDv/XFKI4daz
V4tDJ6g5d5+Ixy14vKku1GS7i9RfUBWhdzAv6hB8OPGrUyOqedgPPSEQSTQN
COgIBxDrjNxaoHzdTbgQEW5Qsi7mkRC22rA2oTLwCTJhdPVnRourDlwHjfQf
3PO6/k1CYZoiIch+2zo51BqrVunsE3sEh8QO4HvBa9ANuQZUaHCSdVAOQe42
RnUDoR4x60F/821IU4JCDAlEWuFs1K1mx+3YLhf6NVIiseW6ijd2xrBHahIi
nYfKmbCipLZHWj2xpAY1BfX2HW9tCCaDVIkhTR+iMb5sd3S7o9LSyGzSDpQl
JJZExfqO1K/vycpR9i6UhV1H3XvW7ehMXXk87h7h1RwqeBa/ugDLX6idxN/U
TeHJ7oW34F2SWYWL+NOliJbtpalgjvuB4VdUgGdGgz1KW7QbqppT5v0vhZnX
ekSIoBWzsrkacv3rPw+6UhxGjdvSGq/KBGlZjtJ0ewxlhncceV9EhZ1G3Omw
zwGqBRgPgEJ9tWzGpq9fEdH/AQ1LyPQbVlLptRIfLVDHN+iW51Si9eWUBKHl
uySnW1pLW3l5IT4F+0KHDt4Yfvq9UGqtczgIOWPkdUQXZ8IEEsYgyPi0rQTo
c5EcCyHlCJmwUu+f2d368/ZFsCJssaRCg8xLTYIJSvmjoQIRpObpEQXED0Xv
nAK+BEDLLWLAdmV6tsPCONmqkYwIFYF2krtzOm5An7n5MmqK8KLBxRlgV2ia
P+xrLTy7USy4wv/ed/KY/cqhjD6CSDUtOz0z4ed9QGCWUMVJEE3PtzwatBAz
oXVU4I++nH1Ra4En91ZX/fMkXt+o1bOA+Y2cDEQ6XUlmRs6BAQuOB7n6Kj42
LWUBIAWwdIEgXPguE/eDxYYASt1KxkVPf/9+Oo95OQu0sodsLpLiTKSU0K0Q
5uPL8srqRpFnSXaGJx24Txwimw8E8zPR5SNXO5wSBH0U+tlH/x2Wi0cs3p1B
82RI8uNz8FRzEg7VKngkoLg3WOm3mMIM82WTMpvae16LxMm+yr1MD7gZnPuN
2rJAvbc5rBOtvpro6BTI19k/i38dGG/CjxBn2M0RT975MzgYDwuguLyJuig1
fP9c4Fwsspm18LzNPoNkuVCrbuf2WU2pUHANdZVf31a8cesXx0Yzo78P57Nm
XOIQOkwYeJEvZT9OBeL5noZkhgZ6wA9RFnk0V5ROzBI0Uoiw5R3bG91Tt++Q
E7z4Z4HHESML2tkFSkmAgK01Ki53nqvnLBCmLXldQyX/NzV6Mq51f1LRzWpV
ju7JdmwlS6gu6vGSXzcykunlVh2EWqXvgYk+L/Zn0W6ARJNclZXzu+5K5cuy
FNwXiq+Z99PiCRZ3dWfmUg5ww55CQiz5uFjc7uphtdmBfiTCW0nCU5ui0iUO
dU0GtgyJbpd6eafluE7XCC/zgXMGIVH9NJLO5eindjK5HgmLx7/p0IIjtatf
uMw4cIke+zV4C4KsRy9HbsL8Fcej01N2vZmRQLGPXjpVXaa2eeZcZyWAXqoP
sRqP/3l33fXWhFUCw56peE3EW2Hy4gUKEI8/D6JxmaSUwjy8Zxe0Uo52n4wo
bYY30h7M4PaVp9u7iaAgiRUdcSc0RzfJLXvThr8GeXU1yFWPnSXoDCBD1BWv
1F3AnAH0RFMd4EPvV++ryzUWS+wXD0A5VHU+WCFVvDpYo2Fst47/41rq310X
hlT18Ajsds3D7FIJGm4tzQIHQn3skR1GYaqsJeBDsuSw2jFM3eMZ5vJ3v++i
pgOEAOaAkvwrxERAmhEzF6KkSIvbZl24mCCp70P+hu3u7YC9qKXWfeJNI419
Hwl3GaHE9L31fSMe7bJ9DEJu5/naYEFNT3iW+gh2O9QYuBdQ3Pqf4RoA5s6W
uBu5+MznGUT/QRW5XX1oyP2w6y3QHrd2zzHvgvU1MkmzB4+i0UzJHwn97Mc1
EaTsyFzuk5XcOutikyIxcEtjIOUeoH0He3S6PNP47aGA1eDGVyQmIVnkezqt
DyF7alEx7vZosWWqtiM6YvrstM7ZAhD0Mutj5nrjZZXN15sEGd8pCu8HsrlE
Tu/T0JpN8NVuN50uoykqVRHLseMA6DHJQDW46qNWgO5NiJ4zVU22qE+4NvUf
Jqkfp+sLbzs+jDi21a5ikKQoxvuUSwwkbTPXMmP36mQmeZe34vts82Bf5o82
rA8SIfOX0tnMmH359skNbx2LLLI0MmYU7ZXSqfwlFzy+RUSkliCwnpxce6Q9
/9H1/pUwmEEkNMgpTIOjdso6svuQJizMlKNB8X5q9fvrEPXvJSYfqXHKwYdN
jp7rZ0XsCkdDmVA6phnpDpRJAT8I7lkzYPvv17GM33Il9phBRsKFCKjejzrb
S6udIHKYBXrc1fllffbtAtsh6Sf+ZYt8fz1l8g0wMFdcvcO5UZ3Or/dO0Gw8
1ylZDZiWQXEedFQfobGtzrYmo4UFutRd2UjwtnI6lVg1+AtrpJCOy9CP3B08
m1T9iym1zKegSyasvnQ4iI2D1kO1xMrT93kDcodzzpZo+WYVCjQpT7QgJpPa
kUaAb2fzk/xCpQ0Iz6EBOJKIy7uul3xogLdfmWH5ZqbjH/jGCQ5BGhR61MEH
Mai0Z4271gQFpkY/vMqGU4Ma0BH9HhtyMDM0YkT0O9BagABBLdBr1nYynz6a
xq2HDBADwQLpgeDcnpZZ0uNTNqU6wcNEIB7/7Ji2xhwRD2pFV3iOwXQRnnDI
VXTTzDAFnQZsysyxoSihCZMq8m47ro8TI5a9l2CWA0NkCSfOfw8yTyTRMGWf
HtbWOR6qfxVTqQ/30xMh4yJ190LYAo3ozfV2CqajDB8d2DgnuV5XEcNfay9D
fVpTm+wdMTqZ22dAFtDEhWiem+MEPe+uNhIrzxp8A/YBqP5mKbsKR4TA/gdP
Vmi8aaX0e6g+L7qC3mi060BBEoa7ztkUbnx9GBd27PEMkKr55NooVm4ffnOh
iWu5JIr3WKK+jhU1eMC/CXX4sOO+WjOFn5QH7w6iexoQoorZhvN5yu0Dc/hL
0cNxeIExS3tR0DUzpqO8Fb9Et12jWdKX9myAT2jwoJ2NnWFS0e5wQcSDl5hL
AUbE0vAOeJwpcvQo3e85IJbpUAKxMKzzA0+wfz45NkqxYzyyS+e2WueHAkwA
oeQszd0JLSZdxvXsKbx1SRXH/kFE95DEyPOfH6WNIUcspEfa5pB2p9MaZYbW
eiLewfD92lPqbd31frKhjdzHDOuXcvxdwhVfaVoDTVWwJdTxznZmGd1tRxpV
hIRxY1AFVpx+jin5mtg3iiDdSwVfoOSDG7EwmvbAbUiBogLcxpxE7SpR9aTN
JAJiXOrsHW7rFT8IdFVu3KaqrIbXb2WguwvjjOC2uOt90HTr+jtj/E2NL/ST
KMkiY+Ag4Gv8abwWS4ulraw3lBIz4l5jhixcnIXnczPS+bOLmv0ff7BxTE2Q
/eGNEHOpjEepNtzxjt49ZJ2YnvcEDzHU3058DDEuCGSIoQFaqQVDfMHv9Ka3
z6w3xvo2ldNSDr11gNctS2hnkC3ageAdXS+0Jfw7n8e+BiOMNSxw6tZGr5bG
5HLnTW6UnsyXw8TG8BTtnywFInQG96tCRpx8yIXDpwOprPtcKwi50pmluNxZ
m+T4lJI/FgnkibowjosLfdYjgqq1sZ2JYU4bU2wjUdKERC7W4meLv+PNEYpw
hG4HvWYzap/1zPmIj2zZFCzyxf3odGawg46RmzFHAtrtA8k+O/Z9kK82pUT8
BU8PhE9ZzzFwu3n4d0RlW7InQOVq2UO5RKPbxCzbopdkM9AWHq1Atif3hGqR
tf1hOi2RuSX1EPVP7jr2mRB/CHb0KZi9L5JWCXY5X0+H3k36FAAIKni2dppS
xZhG6Na2H4KftT49y1tnBNgarYOebwE2Ki16nOnzqEF0BOKCBAjzNOE5uYp0
YI7NrmfmN+aDNXL5V6bIAoz9FdUnL8aKLLdW2s6Ic4O9xvmJE5TRtthZcT8J
UtNPgE64VQfJ+43tbbmDi9hJdFaGaM96YVERannh42ms9Ymdq2e99zb2JUmX
DxNW1zPmC8xkNj0I7Gr+/ibyzKbj1DJz/QkjaDTeMQ37vTjnO74eXeqahqkO
ecFlt/SsiTinpyKeDpgc8qvEtauwbg0fBV4uRSzf9IZLonxAFIom00CQ3JOm
JM0CadwYDBEyF24E5AXhV+xUyjfdw45983ribZj7HVAfkH4anaE+25wGtO+T
pQnWcAGEJCa5DIDw40uO9p23KohZXZdM3muSUcsOSgcGFsnwWAc8rjFkmuZc
30yuX2Funi0KMesJPPqW/it/5CFdRZv9unFtV6qZLJnZ05nH1YlSAQ9dbZUP
VJ7bR6VW1nudivWTy91re0zY4oeZfwxB5Zt9NSwD6eDb0RImqsYKECNgwazE
ZSckfkmP5TJfhwVxgmbJo7s9qdzbztzE2yjaENgU4IvD80L7ZUTocPpra+G5
/1hXwphRfemXJLbQRpRPNR/O+/d2rXqaj4l1SNpAWXNQ9aIh2gQJtV+uEFfm
S0xqTUu+Eo0pu3ZLBBb4/1uw14WSluim6PapyMzRLIYbNgYE0OXSGsksSEmk
7CK1X0DqPwOPeUPcThSO+KO6zxK1elFOob86k6VWBV5MFvZqEE/sf56i7ajX
ZzYpLhpzs1xxHJJ3HmOoWwzAfh7IjUbtansPjMALl9+1bvBVOZPyrdEE53C9
K9UXRrd7kcN+qXC2EgnxW5Xeov7x76bjyVmctNAieWLqyDfVQtHP7IJ2g+FJ
t5dIEwDRxB2sffJMeA4qnTinTWImKQqHSOKZ0TZrTDVOhpyWDv2E3RqAS7k6
nDkAPGgcs4qjppS2rbRGZD7aGkkO8s+5wm8oV7xSfX6o2/raZGzbajgB9kGw
sSfpU4FkPYOVPXMKKUTR3VORnNVGCMQKyn+X2nuMCS3A7SXI4ATCGi6pxNCz
QotND2Plaz/ccVcye18KotBhxZGRBKj/+PKhW5gDJ3FT3GKUTYMVQLE3owj+
tMaRFkq7WjJrfEiMAOkPormAxV3hPRqlCvlH/LhTcw++X0VO/WOGyczWMLhn
SCA/B42TknyamOjdrWZjipXp6b6Fvkv6yEB961rML9JHEC2hrFlLwhVZOSI2
mWdWZ5s9mX/yfOOnuZ5It6qG+Wn7Fko4UCF5lF8bJ7TOhSzBOKz5oy+sl9z2
s+FOwHJHtLejB+E755pZ9h9GQ51QggzdssZEyWd4h5RrEuaWMPq/JzCSZKcq
iKqufRsJcIVv2R4PZ9Ix/iXXJPq+MnYe8eqyr9HQB5I3yvVI2frCKuZV8Ozv
dwUN2hsmsEwDTbdpmZ5kcTUx4YvXhih2qLCFuZFEPJ8WEGTd/+2q6I3O0xTy
DIBBEYHIU1LMjU4uVJt3zq6VkJVmZvFp9NPeZH8GIr0+Bl7scol4CWvpVVY/
xN1xTP1T/5n8FchW48LvB6Ii755Xlxy7F3r/2hmdd+azGKO0Vbux511KaYj9
SEFpgOZZwAfQmmdLvX6BhhnUaIYgZo66VJGodpC2o0/R7DOcN9nE7GJqaFRZ
ZmNrf/jKfX/jD6q1SQWYTK+XVg4Pft1k9z0SfwQiZqNq9nYL0PS6RTIl5hqA
Tex7HEcMsVCsplX74BEPRlC7/NwccHWBQFLNDdkGnAAwaV0VwlYhZ8PWlFgh
VGMUgzMWYTHqpaVZFMWnjEYjV1ZXwNcq0es6kheL6ZU31UWpwTyjXHwoyWN2
IOaVpfjCyFK3vNnpBjVcxCFL86+5ai9ocOfXhvaNKLDLgMfO/CJY03IzpOS0
zzsCSOswwhTl7TB3yCi0b/GgpDgkUpdSoXjfEAoGd5l0+21hy94zK47AdCIC
0/pNOV7Dge1GqRX8APfuJ0XF6sk12QLRWmBjZbz8Coz935WyqdrP1bhe33g8
5MYow6sPMbi2ObBG10fAuBxal6dyB4Z08kE113cll0d7qcdRb7W8CBp+cMtW
FP34iuFQwc7YnoUfCqRe64zhuzGiCfVh1ioK0mhkDJQc2/qGrkdgfA38CPmb
hhk/qZxbQDXDP87wbp8IczQYXZkcmfJ9nTl3nkPJOkClK4dfnSQ98Dp5d77F
HjyMI9AfO26zWIKPbujeQ1m5rZPciuIuw08wlEPNh6waXWlbkP3VZtU9Vxst
C3WyKs/bsOkoNVg0Qnwt7oTkS4XDEf+I5+MsB9fp9gWRf+GttHcAlyn+HF+G
29ynLITxJWatUzyfVbGW4m6U1I4PNxxgyUrMxcsr8lsq8PZQ5OTVaewwaFQc
INaQrKrbrAJaPKC4d+1DYXGh8bhwL3rHQ4/V3dNysIlbqI2TS9v27dnvs7Bl
JSsVDMnjehcMLANIkpuj/uXLywMGtnMzdZ+W9YbetmqkNJdx+iY8neYKXQ7q
OwsKPkZjPFE2a13OYR53JTFOoSGPEZexEEEJfKjl6FSdIvE+Ra3q2BpjB1wY
RdMKM6XmRFqyXVq8753aIM5+OOevY727BAHbwZeOBlwbqoTZRzxMlks41Jkv
lf6Ft9bd9zjc1mPOEJ0/ZvE2pv/pPthdZLhI72AdFHWzce9OXHt/F1DeVIc7
1DXB2SETC9ORZlC3qemRFeOdf3TBZhk3RFnqswvVBRweYpVjM839kUdQssTS
i/c9v06Fa5Sm0INCfI8IhVyZzI56200B4LAKxre9uCVPtAk7pZkHoWoXvJTg
ZdgdRXKlFbujZ2jnaWBXON/71ZX3ObWty5+5rDxcO249B3a8N/RprXQE3q2D
Oy0bNLj9WxXXpA6YtPxBJ6E+B/bV4r0MUPt5qx822iJUbiVt4rm4M4vrruo7
c8ds0owYIc7diZDP3auiEfqUJ6Ae5xc0tFJJu3kgkDt+9IAO82/Awu1gJ4It
xYlI1lzrOxLxqDURoB1RQjELFAgafs8WbhQcLIztaOdU2QZtnPmLPtSXse8a
HJZar2EpHZXT86DBE7wGmrLX1T5a+AOMIugjdL9NUQxraiyV4k6W6T99PeNd
rB4jzIZda/xdMTpei+mLpToQDHb4O/DNRk05zD9HdPuW5163+/dsX6Tlfi12
/C+4nCLNULtEIDtjFcBLIIaYVGYh86LMqDOeU2HZ2+p5gCa5b6fRcHVnPorA
eIpD24RIRhFtKdSlG0vump7lPzf5YDaqbZZXkpiTOBjeyAjvFjXdXdpLDDIZ
Fl9LVXTZuksz9v7tcKuTza960YkkkjJ9zSmMj5RLtEaco13uNfueolfftNxq
mw9tu/mloFPPzm7XInTpcqd2fvXFtB0Ue2xxY7rWM9bhtu6O2p6DJvWzzI7w
Gm+5Pc+6WrbXZ/4dHsWGTpGO8bS4LzAZ0qiLUAlxjfcXaQBV4bbXLL8h9JuJ
wMVVPH4ZjeD/rg0mUC8Uxp2rXR+ReY5QjqpfuuV1Oi/7/fVGoSwIyp/ObLHI
ZMY//6QfMB8ct1jDiqfMvQNxUlXzdJCMHerGo/kmDap7+KmdrWIt2OaC8Vys
xQn9gMMvn4bHy84I1boHNotns0BIkWz8YRSQwU9IKatvg7KZWMrOVlcIr7Js
sCmm/LIIqV+BgEfFpIqspwT+tiUaGYTJS6+6NB3CTj0iD9ufD/Lvo464Sj4W
T0HnVO35jg0te7DaMCRVolyb2nhqN9ybaJ4cUu9GmxvPeIG/P9V97emSx4mb
x4N9vSMjNDwITAx/Ygwn8MRNpQ6lvoPRP3EpLOZPHBGU40eOT+vQAj9/EFXN
3ly1LY4jWZLrQzWgImh1BM71+wcmOSxlagGK7QSx9zP/MTtVYMXSohsODi8F
M149KtdUbB3/fbBEKK+EECOpzdvy7T1mbiVyPtdWZK+r+Bglbt5VUKJRLWdc
AFP9f3DzO+n9U4B4WTVwY7GwQ3NH3VOVZEs16LGVCdCAeLzONxZoI85czhHP
s1+rQo769ZJpqLLs71LUqGz//hcxgBxwZRVLqJhH6eZHL5NpdHQkCRyvSpKc
G5bAIWEUYqWTfeq7KRxnbvTn/xivSAckBi8KyU7/N075Gqlg9B28R5Atz3YK
fn/3q/gJQdZV7lr9al233uJueCizfZ3l/UQWtNjv9lZsVHm/t4BTMRoEOy8w
maChBoptvyBXW8f1DIRpztTllFOfXVH4B1v2BEztLIGogbXuAUODR/3KyFff
lgYaEKM9evUqhiNyBXT4Owd/RbO79yStvsnw9qyaHTtG4NRB7zu6yzcw49n0
tXTfvvNTfarRNTeYW5URpX6XVWmJcLD4OhlaSeuPKlASR4elKUMX6yaZsdiq
/sW1+GJShSUFQjcbFVi3RnG/Ixjy/AnDhnQvXTR04vuApre6NtI9lw1XKWVK
anm1scz1khUEnqvWAKOZRLoAnX17BkkioOI/kfrvKkxRtciQiKzieKCD2ipY
ptKLt5Fh0VOdfqBXkZdMrfqqYGNzM4XOT31LQsrcA+mbPYiW+fFW6SDqE6xf
V8mMGZxn7Iqob916oBuvlY0mDwH6MpZMNwytbAyb9Tm6pIRCPtW5Ah9vEeJC
24wmuQ5XwU6jWDytxHlRxzyXYlzftnKxhKYNGZZ8Qw5y0rng55WHGQHHPDXy
hajwPhF7V2LnWiWaMCojLYqnYGtVusZFb7ZuldCRkPo5LOkN5jHmiUEtEpoT
yyQuHVtNewnH8033pPb0GNl68WUJcc+zCt1p+VzX8wfyOuc5cCSI9oEqXxHo
iywZ7jpASBFXh6fQRnniMtG78AMAh7UvDJZKSt8TsLhavRSonTzu5tyMG3Cg
EKzASD/zNHXC1z7VFkjyL/1JLN2Xra7D/hnLbKttrBMpRrFSbuSzHma3xHNI
M0bdgkMg1Pt9hxjl/qor8on4aJf9k6h+BzV1nZaSl8Cs+V+TnStouzKhmpHH
k9uEYcmHNscbUVpOcXfFs255RvCXHgRk7IpFH/MS9tZtezetOXYAhNk/PkR/
5xshiaPRudYtH/HFoD4ctbtdiCpuLMDYLbCoMGFSSvDrVPjM8dO0PEOq4KWz
44kyH3W1O84QyJIq8tG4jAnF8ie0ZvPkwDT9DmoXF6YN2H9SeT1RgeThFLpO
BW3pYCjFB4X28STxYKVtIUnHzkKGEhS/n2Gcr8RuRFVKmZasxKglZa8YqjEe
E+N2X6ID5/fsxtxH1i9ztT1z6VrC/sK+sxfLSXQ1J/p0kj/6+A/+dtGzzZgD
nRqi/321U2bpDN2pNaNkVZcG3hu0S8B0e3HjvDRPz24EPZCiueLOKk1YzGS6
ggdFTxVJur7cSDThVA79c+VSJZQqnwLrQasfrzZId6MUb15N8cpxkM/i/BGK
Xoj8ly0Ao+Ph9VkkyHqCw6n7gZSYuVfEpLz3hH575eiRo/6jBDtYA6QVhdW3
i+WFsGNWFnS2unuHFDskv4ziTyRbR10rCwsVNOBGBzo22qn2mVZMFsME8ZR1
cQJa0lkHzP7CtLk4WufodnHfj8/2/B5v+aTEt9gkc7s/+NDzV5QBozpSGuX6
c5u7UZipr4KAfiBCxi7EpyeIOcNidjTjImjxw029K4upjMVVTXPVtVEH+dEy
ih4wPrRcm+6/fZE+Y2qENbO0q3oVk3CthNLwfrLXmFJhVTDzal/ih58Or2Sr
FdDYIkaDpFMh+CkKiMURBt7wTUepVxO70H/h93/HBQ/O1km3/nN1k5A3h3FC
/LHn/p05l0ujM62hpyfvVqyfaaUs0/2UGQO72CcZEA3HIlASaTobO0Yr4k+W
//OFTaCiGZTQF8hZNHBLkOtuHtawX6PDYfSkdNEDEpfgSmxSrAAi6tC4jKkQ
AH+lGioJpWgmxcJf2O5wTqQE/uX4ZpN7Hgapv8bhW4y9ESWbsJHRxaDysqp0
Ii5Q8gA9u/i40kCtEb7yUzJmDVbM+Jx1zpLZAStPEY2j1ckUtf9rcZu8/j8r
cci7qZnFkaZ18jaXH+SSmB26dc9FoURd6KmzylChXlN9S443t+h+nq6J/X62
knS4BKkgdl6ea0o/kBj5MRrspuLS+qBCrpIhBHSWJDnsNPI0V5udY18KDrBt
jmHER/kb6fsXeQTXnEQ/WYqdHbeV/IMcgwJ6LNHOdNvoSWUwSLeQlwU0vXI6
Qg1fQbz2hVobHzUucMKOLQdj5A4StzUWUArp/Zsfa/jISza+xSJ62ur3qiV2
78Xsam4M5iojzCX5qZcn5vunJLCob+m0hVaXen+6f+f9xzV7yf4mIm8cNUy6
Q74deQ8wISh+VvpC1g0E0WDXN9EdyzFacLsRoXnMiiVtSjb/YVJMpNjTQoa6
EsX2xHJWnQmAhR3YFzUqDsFiT52iqSoWNdywPK7f1JVmS7tv0iH1NlKz4Kxp
r1ROIqbOAM+XoQwo6bDU8eFzdDcf7FgkR9LmTmaYZnSDmq4Pk5mJ+WP8gKbL
YYCPjKmqmUVOTHWGUGN/8FyxyV4MCyhc6gx7ugM6Hk7Ap3g6eSZHLJZ14leA
rtwnaXuX9py2B3TuEXVsBPA0PxKwsYvO6f9NnK1C5z59u6Yxc/4JOdeD7kNC
fK74wg6kxPduH8sn3f+9EPaI0ehSgxKE2nI1eCK01Zn/JbelcFdumb9kF+LJ
sU/649T6TpVBM0RSqq7wYmUaW9v/WMar6me9dT4UZF9xcM5vYscqtW2lJY+T
hUo0oOAnpDnLfja49pGw1aSs4xsS1aFs2bPHx8jCYDZioBi4opUe/srbNXtF
owzhRPnZyzj+YUUoizkDnEhCBd7nw6llCSErunbCWpWZ6KvCijDNGHB6Hd30
KxvZj3Efy/14tNScSz0UEJJhjlVCQLU5227M1VngG/w0jYIUPq/hnogX3lvv
wCXtSY1xzbm6KIwcm5nH+mHrc6hYMDYieOC/8c0aoJrgXpQK2JreQo55O9ko
L3mgZCkD/jejOfQUe745doasN+HKnb4hd0dvul3RqtRzWQyUBWu3U90PNoY5
3qWKw9Qt6zfUYryckcLcIuL2ns+2uYFf6bz5p9A3owhRgdzoW+l4K4bjDcxJ
AVpY2HZv12uzwVCQCoj2pmb0hrgsG2IZPifGZM2uWhZoY8cAeecMfL2lVbsH
1vf+T5xpDMSJqClF0sep4E1PFs6KBLtvr+SLCthNH0P4jEFUDnL1L49ShFdt
0wBus5pUzrZBXlam9af+yjV+MJY9pdD7PB89ZFzazU7eR/urHQUDt1WRVydZ
31I1WfFt4aspsnp/n61oRc/lultTVpPMo6/0aJVaOAz+EMQBoECGs9Ti+/T6
Q2lAt8PC80ZYoNdW4EnQuW/WLtgWYHmY8DqUoygaIoujJ7wiZ7jrfDqHH3O8
Wvo1xOujMRgnN6Lb0cMelEUf1mbJKbifhrLtHEuMLGPjA5o3+G8+YiL+tITm
8Lc/fAmZJZM2AC3/QPSZ/Z36x5muJC/9iZGo+jj/bG7j4vAveTAq0of2gCej
dcQzEJIHROy/59ZRN1ZcN8zfvA27IJ9Zs85syV7xUadn1vEVfsrnepYD8MXi
ePhuhrZWe9c8R8JVEaY6Pxo/X8oNSipZihfcQpHI7ZFHWJhcnZaVicPpf2iY
MIF9ptOZ1qXUCtFDUZlgl/9PgyyXbZSDd+OcixTejH3ULqqurAm/FGWzu1ju
Q3aNV83qezJE9J3nqGQRsusJcxtd0F6/mPI81AK2YrDS/WpOFrKbJahfqCUe
E2Wyceml8w89Qt5vNKErr5rdvEhiFS+cZvVga5X5lincWEtmVwC2eODrYhYQ
N0DtXQh3Ly4WhtRpKjyy34kbhjCrUOOqFfM2qF5A21QamiQ0SicfFBHqyi6N
i5blAKd87oyaoDPSsh/eMad9XjOPH5EXBC5XaCDov/SbOEYWbSyQKBHY74hj
LEe4/gl0DU7HpECkJgHSAM6hEADb+KhlJd39eDQ9huMnMR5l26toDHALSeAI
i+QzAXSEQEqBAk5y9aGPBMlhPtR6+EyazqblfYum2PzVT3SNykPv8E45n74O
xb8/OeJTb2jDTa5ZVHnGMPDT87krQskCr5jOTY210dOBthJO/phyvJuxMiej
10Z3ufGjzrdbO44YOss3ObISZ8oarj/QLSpcK27MXa6ME4L11ZB7qFctAIRm
OXdmhp7cu1+9CsKN/670C8jvvW56+GUQza9DYm6Ntlu14oUeYNUknxfo7kUl
pe6hZpB2HhFu9tCcyHg+NjrHjaOxdOLUhaidXQD/BhH+hBXGtvJB8MAwfsla
1OUbu7AhZbZGEWTThbCLo1tjTnZh8fcz4AamZfiYYeBiA83afX7xbJz3nQrP
Qm8m4WfdwOFGlEatSkW8Ypb7fYDNFILrEG2G16yy2qfOn5Axbuw00s7wUXxj
g+szVZYlQOW9K2DlSpUT+E/1EeJu+K5ZZhynFGKGs4JO4fyTp4B9KiMYL9/A
JsiTFr2A2BN4J3BR4mhHWXCh0LPJ9Z1xCGr0nEgvUjmgOd8C4mrKPSiU94Jj
tos3hFecAux/tSc4fRQoS7CVsZbyW+hSeLrwgWI2n415aaDqfxsSDAbxCINE
XMo0OWxCrlnf5cdxkuj7KNb659tna3VGNvqa+Jr1Ew91AMJw4wfj06lk1KZB
rd8lL6IzfHe+coLCPIHNArsE9c0y6BnMsNJ5cbfhIRsQvfGXaXcelYiOPZRK
S4YB6DqJqtMnFpRzzcOMLf4jkkyl9sReB52vdiHvzIQonUXe04dSwYzQEd+x
Ce9hRKNOLv6Io96R7KvSZ+fecP/0FWFtzvt2Znndv7izv635gWGVZvm2CEVw
yvt7oznr9ncyMeFjbY8wC4/XjMkj6FGVIDyYNgVFTVtm55y8sNVune/y3K42
TbGsHCKHZC70ah4Y+RzzS6A6Uu4igUv5HRpHZjuM+2O8MV2eHMmMgtLu07oq
e0NsPoleyFPOKVSPWWf5S6ksUlKFQZC5OBxVEKQEaGiHgzzERpaP9yXwMHU8
Htod2TGf14au8ClSJ0WWqKhZYT95IGCIVYSyGTnM1wj86pWn45D7mUJ8UiQs
dGOvGnLqHVBk9RudC1pzAFFSEv71ny4gXHO2C0CfCAuxkNWtGY3v/v/Ul67Y
AqEnM1E9Ei88M8XKY/dKNAO2R3XUZYNRLmD6aviNGP9pyfzrDyWghMtffe9T
wWnAcbE0OcjGngUxZw+2QukSLVj5u5Styc4IrasQA3rRH1XD9+Eo3TPRjf92
KGeglJ4xIamwIcGB3c5ERWh7g+JVpgpQ037kF/Hl162jBElBeAAzvad26YqC
B2uTc+54Yq/kOhVUIVPYICKJsC3qKAatYquBzeNPEIJmwVvVAfHAd+1rHMca
DDvNZhXTNw7j6zHTrD9ERzD6B7vNvDAgjyDNbdiF/XKRPEv+jJd9ZrQOIY3Z
a+QyOdditAr7APX+U7rfHSWZfXXMuriyIHiYjxQCa7hC463O8h4/S0i9uOTD
A1ZEf2T17W4pQRR+mzixPtWtH4TPkxOa8FmsWPEnL9FGj4lOX+v3yE1eRL0V
CWBs/HW3ve23qMYvuQYjmolZD8rl9Ae01tIA7xyAaqOLG1C89W6iEn3vndUF
f1fLNIOw9dKGWbhBdvUJiWn4YEYp20ZOS6p2IoXL/uN3JTl3Kc4FkcKwY0EF
tPl/bK+xMwnpTyVq0mK+7LaCVLOvqTwvzOSLAOUeTp62UYaoUoY+Fw2Q32RH
Xs1qozLFpxiNeDntyHMj2D92yADbJhEeWsHHmQV8BQs754gFGOvV1F8i+2GQ
42l1BLTOBpPEDCv+kYi2ob4/Sc6SS1cay1nQgDS+d7IAXF2Pf47PRfdI2Z2/
IGl/hqpqWqed/2+uNVTM5s59HbZGbDJadpw834rNAu4vU8qqrBn4Ggl/u6Qf
J+k90YMQZIMjoispYgwKh0FhEYGpVhZM9JoB5osZ1Sr80dYzPIQ10GKdItNw
dmoCMZ7tkqD3cU8dDG0/2qN94wMDCpB6nyKt7S61dqmUhpE0O0nn8Dw23NqJ
necEZgOTHfx9Zi169ORff6+amGyD0AdxV3HD4UstAvCeM4DIeh5N0GLevU2k
88K64c66AcuScf79TabseMCZw2zAFC6RD0enbX16jsjhx9fxswV06vRYRrBk
F60+hLDO8+D5DDUzDoqqxl951jAh5Ii3A+liu6rMz+VLjhT+tOJvW2+/lqFk
GvoH/fSRxSsAcIoVIckQqItQh4DYomA8VIEdy+I4UWeFo5cADnhCqNH6OXkE
zFuB8oMN3QcGyXkROOCNoFWvcI1ht42cfNB3SBoPCl126oipkbjjnTYHlHZB
5P/3ckYL1t2EBHu8GW6wRJSjxhTMRvLoy8weWvARj7NcUeAIQfKAnkVbOywh
MouSeOtX1pYDHiQahxMJ8AJUyrUGaiKfoZYR+xRe1zWumHDmh/ktT/46nhkW
MV/1wZqHon6EDYpNz1r6pDZwpRPSEgsOA+0kbmwzHgsLb4/cXJNVhKpfOL2G
PehGwnk8/BeAdKrw0UWc4eZg//gsj0Svkm21Gh7XW9lliwEU6hId1PBzg1VX
CKhyrC6zkCeoqB6Qkk6wdjnVyg+lzxMNOsFk6GEW92kMuFxqiE5QhS5VVxBn
yCwKIuwpqJibzKmyzh7UCbaM6mgQgbCAycgszutE0v6yYYIAI9axQb4OOHbi
8fVuIpzBatkzw0K1Vw539xHnJQsTAOjiz8q0+Lqwg1FfliaEZG+myqkk32Dx
P62geDsnrBbgUKDZPqzzJYTAvPxUp/QkI1EeXiKbt+avbHF8FteJ9pvOwCcX
AuVyJPZF/K6866pQVngdDgHJg0G6+8Tb9bgJ5VXF420OTV+5PmxrLilWMWbT
62CVvCEu6t45UulVGN1tofdXwHd4YujKWe6q3pbLJ3ntWlkrViSH/fB4VH0m
fTePHzV4++ckRH+lL2PgnRKbJxYh6G1NmerNBxh+bETHGlr754hWR/IPmM3c
Ren2WPEcdd+oRJOAxIfyhBIxQ7J7RmlWtfWJGuwATI7Z1UBQ+Rwa9Ra2jwUP
HeX33QlV05wsfVgMWCPa25b2KErSEUiTtWELFyh3NslXrW+qDPzIuu7H/IYp
bBEWMV27kN0v87NTOneqdpfL7DxF/T6vnjzTYMP6FSZKU2TM/7mCHUDlAjyM
R9l9RoFHZNXBJueIVse6hNkI6TK8RuGQnShjsWx7EP51zKjs11q69bJP6CMC
bzvyIiSryp0vji/OjvPIyjykl/dAD77Pp6eVNktiZ87/baTc/gpNB9j/uYU/
RUIkV5eCyEO7LSpoPmMu1VlThP/BLvRrgSaCRtZaUmJOs9eTD2HreVfT9CdK
xuotaW7uJIc3eJMp8bpEtrhO5yfFT4ZUwUMm4kyMB3Vi9gAyqVHjaXcjH2uq
5/M38GnBVjOaBm82yZ7R5E7M80Dkc26/8a0Aqn1LxjMXQvCboJxDbRuLJGIk
OfwsIposgMvgU6/ujVyJyipvcz8iIq1ppm+WHAd14yJ6E/OavzdUtztfj7Q0
GNVXvey6INjpW2Wai1sx5Ya+V64JvVdij2oB7q/CX/HcfOAj4EEpmmIAGkJZ
o5KVwCOZwTtBSVSVM0RgXttVUZZFcFgVL5rmAOnJkGzNw3bid7oUnNp3KX99
xt/ao/JfJMQ93ZwAt0TJfxNrgkHiF43lnKHgwr1YCpVqpze5jSnHlsx+UrZO
D7TWKXB6UJZZYPeRzHxrSoT6GXK6OxGnNrvQLky/OdyY8DF/4AkX7oO6YAbd
mFU+7zmjyzJavZmPwrgE/dTehwzU1EC4D278hXtYLXgaDZYT4s+1cHuBR2oi
TQcdxL+l+z1WN009sU+gGDjzKzenRnEx9meFMyzCw5E4dAuFwJNV76w5Qw0D
DSRZBzXBoS7iOINVQ+/mvjZS/xdP6hcYUbry0I1o9TCe7GubRJps5AoCNptu
7qPmnBaNCAl4itcHe6MMZrItDcAkp1Tthp2yDpiEmV/E//D0med16AbfwM6W
kB7Z2Brr7Vwnf3ijPmrF6HWWGJEoDprvw3JLUtMljyUvllvKagWC93kReV/g
bpEGWSKQ8NKGcoUtRs/J2qkzAUsellglOlJi8h6dIKxob0s7JndDvtIzEKfF
LDs3Hba0umwI9MzpZfOLb7rBt8NE1gYzyZng0+ZChqLNfbGLNuJ9F3aY3BHN
C1o6coNObffc1CT1g57lc4p48lDD4GG5G3gV9hGFvBXSDzQhRZdkL4iArpK3
JyX6qhdXtTzgcKt/PXB0k+BXBmf/espVWhvUmC7cE/XTTI6DNpcq26vM8Or6
cgze1iBlcj4PHR82iY8nqqT+cqRP3C+jFUMvnG2KF1oU5x/5ilBSLhQu4/EC
+F/2ARFg3yyZ46BLsatLEWfNbN1skCyF2T1EdrkCq+Tv4UkSAT8Be215apr2
AooS/2IayHfWNH10jH/osz2/oD3Ad0jUh/oHQNUCNtFWo5AXgx9jexlCo210
ulRLMkGBTJQXzz6eyOCwS70CaqQ2c/smCi91c1O0pe8Qumx9aIkTqYLPGmXo
p17QF5chzsVc76IFUYVdA7oyRX9n7XnzpSnGWSkbzZx7o2sdZxJHsig9aTbz
h5hZ8CJiLFfs7bpV8XLu2LiA6WUIUA/WkYl3NeccMkqDltChJN8lsJRkk7Kb
HxhlexnMGu0SIoSal2hl8zEc+IQGIduRZBnEaD/Mclziu3cI6Heu3jiV08uX
P8WzSi8Fk/DAJ9ACzl4kZtlqz7AED7FNWbnAs+RnMNmRtJs5p3XsgtBrEesN
KhaqJ2mUjIsvyAAW2nutEp6lYxo8qbtp9/2/A10elxDCBSDd93+UB2tgSxRn
Mj1qvtrrUi77BdgJvM2jh6G9TnnJL2ocPxiWADHpmeiZssy3CTOGbl1bKaIz
mqxfAB0bvBN1w6URjpg7Gy8QQyUhUp/uYUZ9kE4cwH7szTcSIsL+/g4D2W91
YNysq1dYQMw6B1nSvZd4MtAJpAfsUmXO9/7NU1m6qs6hkTSLARHmhv/DCek1
ApWI9G9SAH775mrxHtcujTMWZuHc14DQyq2vcEasZvd+zg1cdt9y/qchk3wq
IGd+4xiwQQc0dXRIBzAKqU6ooVLNm98U8u7qN6SlTUz//yXgQ5erPgYxc2Os
4He6xBL+Zw61scEfjeE2N8cuAPxsl9dASKuH4tpVY1WjPGT773TSIPC75xvb
omqkFR+3miOWJD61trlVdyfUDXw518PWpmDK5RJgVf1/NtyDoac5YhYxJUy/
hsTa2mElzcSFb8dCMmADHzH59WtVRXiRlIyjqF3I6ahtKyqys/KHIrPF5uAu
g1bbMIPEIyxsGiv58DiTpYuVDAZLzEh6mIqGzVrJml038srLBXSSfm9aw+ey
8lQjU6mJHRtL1YhjM55Zi1RE4+ANpPzTq6o3gGObQDLdNFuyqQtCg61Ngu/r
lYdussXw1BmVSkWuRIuDVRn80u73whq+YJHWaeD4dO1pLgNHNk9V9Rm4G4Ee
+V9g/PFWCxY/3AkdQpbGzb3SYx1W03g5zK/AhFjXNA/yj9IwQcfr3axBEfAE
jsfp6rxrk1S7gWm0t5e45phZdo0qZYsmqwBBoGrD2DBU6LMzHwc0WRijeQ2u
u9qb2HlYfMXOEwKfGbH7Pcap8uT/KFSAqwMIYPWINfEbOZCB0MdK/ZIDUqnC
DzrFHWIcTkxDZaxAm7vv/6nQ6WL0P9a2JczKy/5UyMSfOICpxKasl78BwqFb
AlzF6EeRQWoggMszU2krzxIX/YhOLGaDQGXpgOKotyhmwH9DVdU1Q9GZEWib
/Uybiwy8cTYnW+MZzn93TodpGcRFEmAB19I1Pvqp8/aduji6ab6tJHNA2pUa
hT/LH1dDs6EznXJRPNKQbLTB1N3JkKSMEXU2wsBXaQaSkcl/VVdZ+W3v6v/Y
cupcN9tbl9r+LCAq2Vf4KaZhCNyNUPPt3Jp/ieP9/27TIJwcoHsx1KabS7yV
iPFAnw4XNinJfSqTlZ5Hd03AkfpNRYtq7mhEatWrUbUy/HS1+V8ney8jBGUM
QK/De8QvQ95Q/pctgYNPTRMinjZ9phTkgPfDshmfJwpObYBWj3yBRW7VWv7Z
3k9Q7Pp81ZgUCqAOYVW5qnwgl/XJB0yvJMFbE4+2H8DqpLgdzHc7d9508ZaA
PgJJACf4WFX7WRAyACwMLZMnRx/BOk7+N0x9IhxHCmn3yXGu/e4nMkXpnel/
Zf7uIigXdWhnochGl1FtBY1KMbho/dkR2TQZ5Br2qYAKIySDA94IwnfIW3zF
p/4gDGM9x+Sns4cQy6nqAxq/JT3IqRnBX+bOtaQIFYUnBVDRet6i0QllOulJ
9XK0av0F2dq/4/af5yjtRWwOzdZQYknOj7iBGki3YaHAbYA2AjlIjZzpQK1b
0QoIy3NMVI5gP+MBpdBnzJV0KBPWHtm5x9F8+ltBncJw9wIlpGof2N8BvRCK
lryLF/ky70Klv3IyPYwAcm/9nAB7Fo2fJurQSsolwIz2M/EhWUCLucpE1xlg
Qg1rm7CbTh7+DG+KlXwgmfC97YjcuPJfEfDY5t8wKbGMwl/T8Xadj3dlHkT0
l4xUlRJYL10vMHLr0Uz4EgafRpn9Qs5J3DTKJscM204Y6XYgpjhSUWXk9HZj
DpiSQtH4ScrdLnc/z2biT5JN9oD/ZNNd7OKumevwkOrM7Rgb3UuYoC6HwX33
ciTyF2BaLSl1KpQl3Gd+OvRoq1kD7KIwIDsuZDNWVyYuHFqtbHEXoDlhI+5a
u+CvKBdqmckOo89RbEBvnm1YDRoAyHe8mf4SJHvZ/11hdBPgMHNNOR5eXxJG
VJblymW+ZhIeZ7h5Qc73gozQowFW80xj2VYh715zv5lJ2WbZHx/Uemq4uzzV
DzM9ml2M1tAfZFJIwsHsJXXsVELSqHx1SgaCJdnqDVzQmuwiOVLY9SPaZn5q
HdHKlpitJ6RJoXql2jJcUNINJ7ZNo39uU8S79Z77sVIAcbsVVJ+iHvM4eVCi
5OkQfrhakoBnkzXq/VRSROKlwuA4TEu7AiwlEehpegcvtH42pwqFKm7vKix0
CzEN+nZn8Xbm+V2nuB/gLtyAyKb34v1MWMRnb/tYgg2tp+xYjEr2OWZKP/6i
T7Djz8065O/w9WCNmX7CwvO0W3VyBbt5+qJ2Q2GMqvPp7DHxKcCygEhdy73S
9AbAe/coLP8qbNBnjKFChnjt4Tp2TZsifnkpaVAUCksp9F1GYqsaquFLLDmV
hBW2BN5wPq6iXnIaA7lyDizGsuqN5sCcwk+abo05CuslvcYXyiXFCBj29vFL
q9PuBuqzXUkISwEljYUMA+im7F3caxAsd1ge2pN8I+BK783cOox5G5r1obeY
xbHs5UW9BOMcmqEKdcpAkTqwLa27OK7RVa496yA/YIIACqH3WrvP5w1gIGEH
GoMFHS0Rl4fz9pbiXaWuYlv9YynAPHNRVrLNxU9P+BNuzeSSODO4QTAxw4ej
tXOCTBOL+ewLPRWcsW2Qc3S+G3i7+3Gu1msHoKBh3eWFF2fm1fGOUhIPaFYK
0tmM1CSEa+J7fKwrVFWCxxHU70N8mFHPnuHQvloe1tiVZsMXJ7pqe6LIOuRM
TbQBqp+pbSAf4wErK4XmGNfCqp+8An0F4KPuUY+snciwMbLr/lhXfedscZ0O
TgX6tpkerEqUX9w9fTBohvs8upM4zlO2uTvVTfh5u5r+xWeS5Dyx2UKWFUC2
UsAC4c9AclyszoyOqN6LpWf6XaQac09OwCSJugMSy4SJSj6kyRl1AFqXR1lR
FLR0gpUYWRvHh5AYqWn/9qxwiCE6BoHDFFWGmnxWkYWKilofdtXkGgtbPWb8
QeQCWsoQtWzZcOazp6EbmrJiCEsU0ttqlywdb+SAOEx2wQpWgdT+49JiZaxq
tPwLqjHdDutntFfGQoDSnEibm+ONR3KG6vHUDBXoKtbXgD/6C2cVBw445E7h
BULEz7Gv5CbvUG1SlbzaiRthLffMjSicMbMIJqbX6bj9/96vXSc7YOpJlduf
hh5ppKkplvGpDprdBOtIcpD3rbzPLmofW/s46kj3fSPLtqn4E787fFj7BSNr
QKFDDuSycNnJKA1BG9bh53W2cLv5P2UOEPQFzA/o5/icG50hFN2hqHFourOz
PQrP34LwZ3UcGUsFXL7uNgB/r/IWOorV0WK2xhTTydNOPDRcdYys3JHT7kWM
atGFt7UEzk0qhl0aLDT1n0sx2shFQdBRjms2beVj1rEkctGnyerFmOiPWiK1
uxnJtlgMQdzMNQzGOWm8OK2nlHouFvozQlChHJj9yjJcKLy2UjCjbdEFfqxM
MLQwIIdVPZKPQHXroOs8LIty9i1STPGIdOUDguAF67Qp7+rcXOLCx7nI/wCc
Xw6nI/nVa9nJuhc6tqlM60PR5fjvPq1Q9v7M7NSRtR88klMcMiNh7q/nvTrS
hXW0bl5RzZTvetLDv1eOzFE1mDKnSw9PknJUBzKhnARpo5vI7ODCXb+p/fOi
fnqWSOaFV2TRX3RRWKFvPP8ZyQmuSzh8eGinZxib0a1/asRQsStP5tP1sJCq
tVcJKEXT8oHsTbbumQX5VlkyYhWblAJMjci9JwkYI4n3S5XE+a5WZ67cPa6r
Kr/5UbRMG0yiSr1THTzsqAd2CFm+A/tprUf3a4OF/bmUjajgnmqMh4KflBfB
GPxNG8bnnKMlEsVfoSephvTTmG3QlkHOBq48ErtYcXGGqKhgYxx9fuaC2eHn
/Fr8JN+vNBhslDVSf2AOyGmAnByAIWgxvarJnDzcGBx0m9GbxAn9nQEz9yQH
mnkR75/vZQUTkJteqpllFVsRn6a9S3sNPKgRO3kJpg9sguqBCMhaliZ0ZGZu
bYOYDHECFNoq4Dx81cojJF8KKK2uCDMRtlw+IpeIl0lD1U5PGFhBbLYg/5kt
ucD0o7b3eVD6TD5I8nz8JWxRKE+lql8mc7VLLDAMJI4sBz1FuPd/NSYQRHZJ
HznoCinxqArKKLDBJS7e4zvLTK8RvGWxP1aMSrXJVSFQ8HZaARY0e70cbvJn
nNJrw+RPuv8VESdXE7sgkRXqN0W0h+g1nZaDDrJwP1brI4S0LVB6yqWw6Fst
QTrbZoJMnx530wFbs0u/lwWvS77fiqdmWTqm1tNqrmwI6Hz0zdBU8jykanaf
y+tWS0yTAnwFk4DP1KVEnLON99tWm8kRx/qT4QJxrH2XVnBlcgvENIf1Tqu0
18pmmPw7qGX/eOSfPFY+T/y2eMSbi2/FaJqv2a36O1VOiM0ptVsVd/PJDyvw
ja2EQjVa9V1qmDOXljp7xb249y6UjkRRnMnFD9y/NP2piRwIEcErOKuKJ4lS
ked7Y3aE/jxWFs9HvGpxVh6K8rceOSdTi/hdwhCYnbnDdeaTQk7C6s6J5xVB
j4+W00QXy0f68Glys3zH3RE0xWf/n19mU4vAiO9FPisrP/Fy7hwzIkMxeXTs
fZjY1xekwP7a+fva2hNRyZIFC3lCAqOM/r03YDytBFTP/w3oaMQ5U2uAjjye
gbQvEHIGgXhG6ljd1FepuPYrXuumTobExsVChMB7RWv5etvJtV8gXWF4i5yM
cstCGGaWsllbOKqsUoN5sPsRMtOostMUA6oYLhx1u12dhkpLSbj0jd8/O6Tm
aWc+QQpXxUrVIVDJ3CHx+vFzY/hAe+rOn+D2SgKEmvs94ksjTbz2rd8yBEJM
0c6RNLYji0vXWU1kUL4/2UfVVJN3HapW+TCTLAqlHAMhzF+Fo0dKm5NlVw3g
4NXIkFWMY6VGDdRCAPOJLtXhjp/FDj9SDLBPCRztTS5cDbinVAwAbQSJ8pwl
mBE6y6qawYGr2+mHx54gx5PQS10Sqqtge1SHupEhOYIrxv1vbpgzdr5zxYd9
9wM95tLoyuf1aAd8y1uMK7Axa/0JWJb7iZPWjCbxzXP/6Z1zUKr6Rd+MkEth
X676sl0AVTwKldxMSBlopfk9yIMBfzCpjN+8qZq9Xwj6EHkwwfBwR49Eugvc
f61gus6uWHFH3lRSBowI9V/wFmkVUm+PKbBvt9Ft+JzvhaU6QZne7FUU19f0
M2VUtGd8qD9EIoLKxmlW7KcpM5yPAn5l4t3DHFcJTZDKuvVhujwvcztiIPHL
4FHE1vVxg7HktKg5q6jYD4mPtEXjiYqQzE6+hV7HtZYzNwifkoRZv29rpF4j
QBTAhFg5os5uSw8YSedMsSt3yCaf1e/RHIqTUowY8VKxLx+Uf8baZVsSG8E8
W3COdb6KjKOjrsQqbwc+LntfAlpJhji+BHvbFK+nWT6cQo8j3C1N1H+m06cR
llIgMRO+J3MYI1PQGWukgMBcHTzt8+j/39hNA3E0Cf9XYRn6o+juBShdT3jN
vQcz3zUyG5bA20s48Q+4zgGFCTYeMZT3msMT7xUyQp2kJuxpxiKPXuuhIJem
FDxffA7HHGyZEfLirM+T6J67PpfcHQ1ZEP91EnvGnBhy3ugplWsKPw8tAHGe
DcwCHXnvvqKgZ+RcLPt36w+yi4FBDjJiyFN/kF1s1L2Cphcoy+b5K7SxQUtE
FBdXlpK5Eypv1AelGUPZQomDrYsILbz4wazAnbnhDPSBMk9jj9IUJEYQEeiZ
SKjs/4Hm8mJRZ+SC6ae09E97VdO7CeeTAB7x9VfqOQnTOccmNJw0TGa1SZhS
Eq6uEFUyiZGEt+KaZYmwvHC+B69gJ/blQOqov2bzmY4zz5xkLeeLOiEeoQQc
1JbCDXmqo8ITnBxaS00uqdAJRRaxXfKRvT9bf++6FP/TyB6UpILpeRnDAZ3q
gwcXQgVc/maPdSeZbltRyb5yB6XW1sqN0VGYRE7LDFT10IRsEuplv50uRtqL
cSXCS5SgQROBvsA2PUONsYFXQw8Lm7VsUhfOQiWMasW1u1/IWmavfjOz6UFU
z9Ze3tdL3NWsvIXLjI1s5ryNDTICW01lGY3U2r8T0X7noAVSFt1kUa20EX7i
h7oQRMvD64W/hJhPCx5XS/lFptKG64d9jgPh9Vhz4o30Dyq8HIiw1XvNARS8
SyWHK/DpwiEanQFS6CWriiZdCiglLHvzF2JYqUGHGs8cXNYDT3XFIl2r2s0y
P0BDWc/RLz5jrC65Nu/rwzwCnJjYgsuyNdjzd+8FGfBeajC6LyIocfht3BWH
PzdusTiINWryOBXWJCj1uL7DE+mZhM0Pl37mKd0zXguCOW7vzwEpmu4v22m4
BYVJx0YzSVlGp2qss+PYKQChiyuWd38gbOs1sOxzojcIP2ujDdkRn2sNKTHe
rDg/ewzsNKI15CoIJsDGz2bfB4a9Km0ee//fU9T1r+eE7ggVKPPterQXiM6y
jxlaefSOoiVyr3qUke9KM+DJf0JUq8mh1WYF9YvfXrk4H/rMzLsN7m3v5jLW
o52X3Bp1h3QpVwDtnCnPbxGSiXUPedLUxV2dW1Fa4V2WWAv2NwiX+Vc4UKwZ
9KRDbx8VJy6CqUuwH0R9OEVRnLUQ3NikoMaNhbXlf7kPSW+TsmWrAupTpfV5
sAcGU2t53+LoB5ocYAMmIU2Cvjp/9qsYB2X9/SQ4DyLK7TsM3KZ8IcfKckBL
JIvRZDWqZfEcoPPcOi1gVElrZnHBilfOCf7/TNPz8+am0ti8fY2h2K0RLFTW
seUS5OmJ1G4oVt67HY3d4Ee2wlhFDMpM74Z9+2bTttLA52kmSe3Lp38jBMDK
a3ngDeks6iLCVrJtku70Mds3mQtV0JlHD4fSdSUKIaZ/A0TXJHwaLt/JolnU
43mILHpFVvVQYwaBOJSdSqfk8pQ4XV5W70/5qoLPuTcmzpfqeEB4U+mAWf03
dZ1Cv1sexo3Ich0vY9hjDDFyCMYmnPEcNUzpP7GtkwT5/bYk45IZD86pk3l3
RSpl2CSqEFjKcB3tb6SH49eUPdQ/RKIyItF09ZPVH5AIV7T5kkOJ0f0e1nOg
YdRnE0qR8ZRpYM3kfJDj/6vYqYgB8dxroAVAPnN4q7F37Yf62mZRSVy+3G3k
4BU2dKNXV87JkEFjryVbFwSHU5paA2GZP+cHPfO67tmWQ8BL4cJwozxMlolN
1CafAku5k6Py5ohrOEzYfarzqlc1R47SmBMP3O7cqqdZ5Mw1dYJI5zInGJGk
d2FtpEfTxoJSz3NhqqqXh+NJ5sJO4sS2GajfLoXypdFFYezaDSj2iHx+AhDZ
oDVBVntsfZw2D5OWFgTECgYBsjlUogObHpsH59ioupSX0JRdWMj3uCsWS7NE
jIM6jjL2uSGvA8ErKzE9Zu/vTIyyFJmG9FZqtYe9ELYGMWZjTW0vfSPegiUZ
5r7Gufu7hWCydkPL+GjLio59/P4Xw3cAYqZmaBQK1vZTbKbvFLMgnIMMvaci
t3q6Y3t6CHzxhSYINtJY4UY1RjfPs/wqXlNjANbgiB8Nerh3Dx6A8DPwD7zX
m0CcLvFOf0y9Y7koYTbdWXiJgb9gS6mewwic1ydBsofPGFOeIBZE0p/a9jxk
Feip81wu6AzKRhsqTvmxtdxVojd2MTXuNEXjCUhMf/Vbd3nK3hQqWKXF4MHz
Q9edKo9fRTXmMCMxOjcflksUYomulqOHe+OImZgVZaueoVP3TWhLo00GKPQN
rMAjUY3PG3bSpIGuMu+fPBPFpWXgqyFHVC4LH8HJE4OUEGAGzvBTWt2DF+8i
Wr2R0fcvFoD1yi91c9LdwNmjU6HBh/ynytCnrEhd4/Aa9Ci2WWXQ8VZXeIEO
BzEbzTPJUMzV7dxJxydIU4WG28ft+qpG+gKvs6Lc6xmxD0m+KyElUH3bsveQ
0DMtcjtI2WUeJXEcP41CiO4/UxQo+VaYkfEq4+rmOcSLOiksBqMVQ19mZoGD
ghm4rcBmaO501V253mn6mPLDslKycD2j+a+1hnjT3UkMPc/mrhK2OCfBZ6gq
OM4AUOqHaiKRuh7vtFUq9hhxvrT2YK//nZ+7YCE7c3gCBmPG24E65O7VAIHA
BC8qC8yl52lAAwPFYwsMvu03OH2MZnxNoYMl0CteitEfVca4BpvPMwRcArEL
PkTMSk6N6mGp/7Ww+czdAedWDQu9OpOADtSN/xWAG2DhbI8/ishcDE7xvROt
+KRthiLGm30jeGSMHJscMIH1SE9d4lkuoI9o/o41UN8OSIX1EQQccQF81kpW
CLEmp2d7+BSrrUEn5jk6sZMvOthg/PB1DgPYAWCfdAu6BtblL4G8xabPYzRB
kVEwzMw0INUdxRX9g85qwzACOOafr1P9sMeSVRQOZ14kTlWoBmjQKz2R9Tt9
BFGpbpo9CRSdnhaZC9JLBGnqtk+YHRAq5XK3S/kvGX5yKSLiIyjd3XXJfQhI
VqXvGx4bJAzBHMfAV5L87w21q2czGtCez9rFOpmCQID6w2QEQ8HsGdkZ2A4u
YV8vHZ2C9ZbKS4ytpNZZp1aRHkLYFShDiyI4d3gKmQR+Vvp51p5d374MyXoH
9DLMZZ8UCpEIW9XEhWC/1JDBGEGj+mJ90DjxUoi9bp9dAxCC3BCOz0PE8I7t
iyWJvzxqpNFxvc2k7LnzZSPdN9igEZUmls6mFMdkW3bY3ezSKS0yY3Xgn5Ld
Q4VrRWBzJhUEjzcFIOvgRhtzVLz8EUvChslor8QuhckRzjB4viw1eI8EHX7a
yIkbBlO3kA0OKLxzYWScvHIvcmcSyqf2bMDynrWe9H5PrI1qBnFVREhVEmz9
r4hueILJNHFJ2VDtXtjs38psUVgsINrc5r23i21opb6FW+yLm1Lm3Re4/K4V
VqRr3fWqNo3vltm3nGy6DvFNSJAHBO/6pCwNcc248RPTx5+QCi8/0gN63MDK
gQDRjnwhqeD+ugqytEgfrA1i7B+sUkgWfP1SzbwOkAns1xt3kXQ9ACG2Y2GC
NNPHW6tdrtuB3SylPQ85t1LK1SVxBHuvxJ5fSzP/UOdiPWLis6iZi8AdhP3G
TLYVKs/SkfBqKIwRolMEfu2fL2XNtg7yD30+yzIA0Q6Lccy11/CbUGxaYejD
wRpDO9MgnGvG1fdnnBi9W3d2zEJQd38cKpxGdmjbCGECVIB0V3lI9Zn/B2mg
T58BESD2KKhWsYucIkG8O0QNwMFkRE57ja/5aXy5dT74SySDDTAzbrGAqQvM
zm5fW0cVuMeCL6180NvUXy7yuReOfudorVvZ2gsO7z/yRONYKREaqmZ/d2Ld
bdMNQI80Lw7wET66jVOu7D2WGQ+TvLvErrHvmtSRjQzdiBS3B1MWRfvErDrM
MAjDMEEXcwsPAXlrXbKV/GpWj42C4WLhVKzt6II8S5oTuTphjkCJT9vO1fSj
eieuGvNYJfvuJ4VN86y76sQaTkJAELBHMWxqVPPbqXkaCg5yz7HjIz88/z0P
FZ/AgdbMnkW6fS6I8jhi8QkXQ3S+nY8+p3Q1WLQ2QZJU9vUvoLsFU+E5OZrE
sZd13JpsM1bGomn77kPTGBADO4XdIYD8kKpyDxjGG0973uCBJVKpSS4j2Kpz
tsr4aSkNd+1SgBrvw+yTvfJr1XbqXGc2ruH7d1uMOqDRDseEUXgxWGvTm52W
Ac4uPvzVaFdfb1otpn61d9HJinRiTcCTAmoc7v2GQUqkALjTmQX0ul4OTSlC
lbV/ZmlR/y/MDnFMdBmhLeeNZSDfbyo8V2I5bhCdDVRKjOD2ef6knlK+mSNZ
04jLAp+eY+KZYv0u/ZVffqI+GRGTlNNBWUkADSp2QvfWPTP2D7JQwD6bgxu7
LiFV++LQQa0x0cywemFwa732SmigRguqV2RC5Rm/rzunOYt7oph8wwhxwCsC
Sa1sg27zzdyA/xvS+Nic+w1gR1QX3Pzw2St9esVEDSmLz9KuArPwG6AGL3jk
N1JUFJjGAcqoFpHTynZIkBcFHh2lYLmRnwm3LqiLyXXES3/s3dYe1pCSnJ70
g1+gUbNyYs4QEWbuvSLyc0SbhEgN8tomOM5ejdvDWffGFiWwRmDJjV31wAfM
ZDz2WtgF1Jbz4JIl8GhC3pgpwBjB1DWBtsozxtmAZf8IFsN5rt+T+kwUKY7W
BAr5fzl6xTi8wMEc3ceoLhSa8VblNkWp3NMOqGqG8NCpfG8rrtoF/LPFi0/8
K2LHsPHvP0NfIK899bWbjm5KkRyXw+fRyR4aw+NZOPC/DbcclDxWt1C8B9Ix
PlYJhxDsMj0IF2jPQobiXifJ42BAPE+jO4ekVbkXV1pzSZvGhsOLxyhh1gND
DpyQTGTrX5g2zRva0919UrRe/FTfl1qQaIcOPQf9beuwesB7p8OkgIJ0ah9Z
FvZDjU/U4LkbjpC/BPcqBEYTI80uxVRl0CMmhYdlDwNjPggvb8lCtxLArtZU
tA97GExPa+yUjtM8TZm5Ke/Esz1E5lyXhCZSaQYoxdB8k+fGVEnhzoTXdB+n
8p747mE2goNZjaf9aJFLQhuT+tS+Hm3T+hSCyf3Elac2CO9yrUfzeH4u1EnX
Pn4V8zMXYui8v+VzkQakW52gFI/ZUs1g2BuJAGQlJRfrWTmKSp0Yftx+AJkq
99KLhMiPNP8PWwm4EGzEkm60NlF1ZcYR61LqtW8I9mZnXz/11xmNbU4dLwcs
L7GbadRpohigqMC1eggWwfGkhoMQCAQxrXhgBAeEDyuO/V/ZykpDJOzLOykv
5ituB2CbniH14Hw6S8cH+HrfYp3MaMeqLkHAO1MpWk7+sNHK+mp0C7ZYuk3/
I3b0c7jIEZYOhPIWQjCxujQpkjbu+xfDPdgwkImefqorMAcG4CuhgvMzWrH/
quiL9FbkvasPjQMLutGoE0jDmXvSn+mtuX2ArnCFeMIxGq3PNlBfVjiFaW4y
fTt44MkmMF8VgDY714yCz/tqMRk5I8Ws17SzW4p850fQYHb44NUoJ8fJYSus
2IRKpqGne0E7Uf6FKNGao9yMm8Og+0kFtV7jz7VZ/yCCwxLHaWBIwm0zA05b
9jLlih/Epyn8tqNomq/e/G3ZJfr+AYHlWRv3hK2ntz98NJ3YN11BQfjJRSkT
jLJc13l6CGKny1iD5W6BSEFqSUnMHAVKuDI4jOy7FrRYEwYwggQ1cNIsnJfj
bQWiuJ4/rbeq9nsBYYRqPZ3sGRhJ1uIBA6NeWCtXFpOX2N5ozU+vk+zxMdVv
QMFzo3k+bRQ9+vyf7YJGxGZeFDZzdPENPpvwv0k2D9O9AKbmVYiMYfk8ICx4
lPCxDCk7Oy17nq/DLoMGX7ZNKsbFUhs0byBLnIyy/vpFvBHCAxZi3Tzu6UKr
a9B8u577L4evZbbzFFGhGwbqpBEY0J/w6G+k43ojvi710k/DGZRW4TQKEq9o
t9JngQrsgpiG9neksm8K7EpIJXzeTiJqsNnmqJv7kaozOaxW1I/U0AFJ3Kqz
ONKiLnyX92NTQRarb7miNb3fy6gPerWIxbUukvff5grdc6EHxTw2QrJnXi/h
SAqPsaBx4zNCm857gYgxUwj4u7F+0k5QRnhKNmK0AlZMYnW7w5du5rW/qM26
tE7695ELrZrWaC5qG8SgzToSRMe/QdpRT1xO5ahWfEN2gCGkgf7gmHWigF4f
moNpJEd6EAw4cNT+bz1HlY5mHIvl/422PLIjLF3wpi7d5zFPxK4QGewiEaJn
MIrK2Dgkknrp8lStxikLcRaVZYlL70IPbhaCixqCrZeQ4pRXmLP4Gm2pE7IS
LndJAZ4TF/xDXaY2IGycR/Te6n/pfpKamtXVfByiYFiMzgAx7+QZQyUPLIhl
LZkHtEJR9m5kvQXjByA0e5DSkx6PoD4PVE5VkQjXhHl3akpfvnqBPhD8hlrK
y/wofIXY8MzOLGXq5ShCNUB/4cqtozG9Gdl4Hk1gH/u97fY4i7QDF9nDG/hf
fPrLqFVYwzWctuH+6udXrDuf2eF800TZqMAtTzksGa70teoz4wcvp3KeIqme
sRgW0jmNtbDRRS+LenQLQYwCHULp2F6dofUnXK6nH+s0pPmZuZEehYix0ADw
76ieFBBLEjDPJVwJWA17Jn1mUkNsdNcNvAxseDUav8W3+9TG59JBRkzs2nlm
aua6lBJoGn11+2riuK3vCaKujlvoTPF/DfAcN3aA+mM6WsILwX6E+RKP/cYO
ZEr9d5cV3Nq2KHTo76eWufAjAka8zDaRcHgKvEnFbIPQU3zbxXpw/js/xrI/
K09sCbTrEwsdhp5cK4SCHargB43iMd58ei9Ji19PS+frH0cwXIawZwX+jrDA
Po7lU7BDKfbw9uDh0wCm/7lfnMSlEeO9/Go0fwzkbvWCcnUP76SHN1+8ePiQ
0EY1xKOVyapnRJ234a98r6JGRlE8LcrYpmeEAeRGJoPCtG6yBzW01GT8A+ea
G6J7eRUXoMbXApz1kZFEq8nJS2VEAP3f2KbHTjLbf3hRLZGxWiz0uAIdI5Ep
aR0qKiz1GGEuoqGbgSjej0awUwSi6Ii4JwSeZUIZMbnfr5EaO8cV5btEuxep
nsovvQVzbdA/ma8SRS1/qHM+1E+8klfht4LLlFtnOiLPi2CmmF89hcfAIgxX
acww8cjX0g7JdZhtwCVujNF/RiRQb7XgF5wg5iOsS8OGIABUxQOwoSJiYWVf
wXeM88gWuqEpTF7jH7NDZwi2Y16M/0SiI4lQYewr5dI5g552sFYQ0Sp8veKG
ZXtk1P0nsUZa0eb3EovS4yGLThmxqM0y0227+mVDVTuqorVqzUI8uUxFW9d1
Pkb7fxiPPF+1/Ptm+06hN7hxKCUBGiIBagcERF7xCI2ckWhI6kvPUywWQ9IZ
PLuJSCJG8U8lVOS1PMdNB94Nzf0PiDVK84bbCCbFBIFRUf+bEOCZOrjDD7Wh
lw70SLl2A0qLYJFeQa+lAmdR6zUflL1CZQyXGuL7DM1A2yTi6zmBUANUv9Q+
Vj2SJWqaNTtzjXekU0KpP9QD1NRm2yeAbu/pwsNw/3giDOAEJ2JLMexDAEmh
4Ak6/T2biWeSSyCZHSsXLJJCE9f9bQVwj8OP5EmfJ3nVLvBdAwdYl9X9APyp
fvEbIKx/dHET2f4OUD2oLN+FAGo39jmKlLMulF1vr1azj7njXGh96CWK/7bq
knm3LRwFpXece7QDJDHe16y8RfOz8NwheWGKaBjEuevGCki1OoJ8OZTzcmoC
GJp671y/0XNl2h8s4oxOfrYwm0T6JfoJj3r3dqsunuvla4G960g7bG2JH/8K
4tSHSlGNWsZF/ZNKpjG3AknPbbk9JJph+JhtgTD4/aAmQ9MfXbrtCZ0PMV8e
snvY+sodphN7IPBGOMaBCJ1cMX29u4oeZIYmk/h5WU4ZOdpQofu7upFoW4E4
4DJ37d8Ia9ezrKXvaAuxOQVQkz/sokn0d7C4IQpS+2Lq67KaPwFQ/10X8mwr
akMYfMrYExLBgaWRNv4jxi6GDmskLx95mgqHbNO2Dnk4sLyAGYp/Mrc90E4W
jVz3J+8I+dfiiU6Tlp5+S4AZEhX0bHHfALU+XFqQJ3OjGiPVy4HcZW+auVHT
6XODCcYoelsrOxENZfgSnQMagdwZRbkJlH/oidjxz4zVKCQ/dfdQK1urZO4Q
Fj1uI6pYgg/OqVepX6i2QwdA7B73IM88f/Qn2KxtuNm0aa1odCgzVPbxKX4u
4hDqMr1XXq7+kPgy8wv+6xOZR7fk/SY8+06MbDforZyTwHyubODx/s3x31Hk
eAjXO30iNrDePsDDmBlN0n2J7jJOkt0/P7WjSvYCsnXMlAIfhMx7uB4lfbXT
R7yMCBE/gm1G+KBFemYxMO9aQcBNIOn7pbihcdS6VcT0EHl8ymi4lK67c20h
RLkj7BuY2+u641NXaFUPP1mANXmj71QJ1DbT/k9EwDEmYIH1zIqjiGZ1159g
3MWjEQDFpakhj+hzyAb6e6YI4JuYW/2uWgUKbehpdBxEbkn+3N4f3nUl5n+p
t/twpk4jXtm6Iw8i2PHAiihTPs56HwtMBhnOu6pQufUTTWMuoS/nvYGFMeJW
qaKWpSqabrpakuceQBWDcOt17uKQJaRnDAaN61WKwXBShK1OINWXTwS2LFJN
zeJnzpofgh4F1O9DOnfYEq0bbChX+xUhXte1LckRofs+rYiED5Ues+W4J0Ru
p3fnpSGr1kXl6/ydbVNzUvAsHlMVCCj+8RZmpWVL2bi8oFtqxE41tBrLwXJ7
xKlDgucR4rG8l4gPLKRf4h+55+FeQIyerbk4dbU4/mqNGgjmyHoxWCjguX4q
kwrVV+o4zu5/UvFploLcHmdypN25t1X/jnENnKlamhWYzQCqhH3qBgpG6wDP
KyegKCBGtfZ1nRZmz+Ga3wONik53HfsK0+9V7upL1b0EZHspfWZl47Vw4zzM
z3yocfcFogpJZQGknejC5pwsw8jmBOXIDM7qGiWDkDqf0l8BtopS6LOzhhTE
XyqWsz/d72DpoE7NHW2B/LaFo3551ojqk7wXpkfCyZahzJ6CCPwYkZsdHuS9
1OImnxtOrNYGCqZjtsJ+raLzHooiQCD1+3QXIPqsi8O0iGZhA7RL+n7lAvL0
Ncg58t/evmL5G+uAPXDCB5KG4rII9G8CsWBxqgb2KuLsw7GGBltc7n4WfOaU
X+mDMDba6cH1zWn+j6Adi4rKDZIUxvuoi5UmbWctWS0M78B1bl/12o3XtjxV
4m99Y+LKz4Lrn1TERDhe4rehsmaLitM3DM+zgep2D86h9zq2E4/YUhlwJfC4
3hYOufBhabtV7mlOSSdW4f9D+Gdi7qHA3XlYj0I81ZDhz8ambOInN+oCcU8q
VkZPa2fiJ4N/4skKBkUgcU3V3x//KB/bAdopiWSGpZ/P/pdDerRuon/hoVQ2
pX+iWt0QPur1SEYCiVMORlKV6NJScG4csCJUFLFGxuPcWmxQPj1D6Ek195wH
flg7NS0Ka1n2npVlypAfyBKdXfYe1WguiYT+Nn1IXAhmEIeMGPWWX9tw3Cm+
0niVPvDPv9rrJpw1KjMjfT7ZX3njL8siEP98N8ePx1qR/NrCAmIRnnAFT1yS
OY/arR+o+ZnBl37yslef6PGO/fEIZSe/RFZulXb3toMH0PpLVZ6j3lxJ2I2J
IBO2odE6bCT9Uz9AtrfXlGGiRY9a/FN+KUfQg2WZssKIW/wMmvGkMvam5eHT
j2HLiFS9CaOP6AlSkCQFmUt4qqkuEJU9beJBki2lk2ejTGOOQ10kXQ5d1SKx
qXtdhvQS9tHTiKWSbYavE/h/FMpNVhA4PFLtSYV1vhwukVeUc48VC3aaVuTc
uJZdFmKQaSyQVk9wQOuKFrUpbJHo5J977jW+Gydub4YWEW6GTz1chzoYmU9g
p7m1iIpX3FnOU32eZ+OwYkdWy7TyFAyjwJa69+L6AXkyhSokwpMSNnLBzAWs
GjBozpwQjUMw/QKPy36U3+qF35usZVoruSEoetOfoQSADG/CFIjC2N3WlddX
5R2JiB9YgF7y8C19NWTttEPn9ho2v3DTTdqm8dsPjhFIRS/6sNZCQuHgS4B7
3MCSHopdlFyO92LUtjbS/cwrEPpEgORBcGqr9t/oqycYBuAizfV8wIia9hnb
NBwxX8HIV0PH4jwBHNQrDQAM1Rqu7G4Uhab6TVpjpFb8lzZrJzn4J6KAwZPL
3/Y/oeMne6k6abQowx1Q+aeWc/ZDpVFoBSTWhTYn7hO0CfjnqdVud5LuQoOw
MbudG2/IFIgtKyCBlOmkPZKMAXGkmPDcKUfXWuhaiewWl5lI41RifrJ/SJZl
+/vWQlu7TlHHhnHK6WnKPtmz/foIxv59wz+zeFaRwqj00UbbWa0WPjSCPkKC
iXki1WSsawl/kg87YigAjexMVX8/3Of5NYcrC8Te//N9i/9aUneDCBB+alCy
hnY7Y1SHG7hvR+4m912go4NjuVL73IcoWkqTCjw7fD4X6Z0KDzUmLou8ncck
ot4R2coks5r63R27YAFYDykHrFZ6lwHy//i89jELDmkR0IAEaKxExO3ZBOts
DHpEPWq7VhPQzw/s/co+GI6J5lp87VeoPylqq5uv5JfpfhDRBvUoSZ1eHiU8
pys+4B3MMOOGNeUx4vcZXEaUVMfwhHt/qF/GEii57k+V6OGdMuowQ0JEPzIV
21XQW6Eref+0RS+9cdv6f1UMzrQWWdKE5jQNWxh2pDr6Ria1LRxr3vP+9tO1
pSFmwCBJM2CMS95uPAQWS57cfV1uM0seguLFA4B5EWISIA/rKwJEry39Ls+A
5tv4TPzsGVhLXgbN+OcnbQ0cNByAbAztROgZ2eTcknKW3Ch9npHhvmbiMVAF
X5azvKeq5VO4Djf1bIPosLwZvz2JDaviPUmKXVM++C0sfpMBuO4MT7EXDENs
Rt6XAggK0J0EEwzWxziYyb57W0Cw3kexSwCbnMiseCr0VJYm1ZBSFmtweadL
NamNsjtOyL7/adDuwrAVR/M+fJlX+NgpK4RBdM83dZWlQlcvP2EKwwWY7AUA
xNyiwrT2qtDxgNWexrhJcPus0iKb0qkns2SC9Nque40xaL8Bp9fIFrXFUKrt
zwZw2bqotYftU2++7hukf7er9fUxXHIFqOSHOO9mIt6bSe9Thgdxzg8m5/mK
C7eooXwgOA0jsp94157QBp5kmsTy2lcah7urJq7oPFs6yCxXIwYmYOfVl1WD
sl1ziBMyCjsZZr8EZ3zwT9W+E3PRmJFuK4+LEgUQ0Mz8+jg8jOcw/MPLy8IM
3IESF8CZPv8MELCWCYSZyuXCNTKYHmz4tRTIDcby8+dZgqTpvrd6jluN/461
5ViE1xyFye1dCITeDlcXVV/O9Pt5+n/htE/jmIhHxq3dh7NluPlVGknTLlxm
s4FkpjtsQpkb42SHPFauvHenvfze4MtRnQuuTTZ4WUmwwlUQLNlM52xi8rml
g/Y8yiPucdGicOxiQ1Xo2cqQkHQy986yqbX+Kep9uEVDE5xY6DdGkKzhV9KY
pZEv8pS9otTq8CZ3lbUYPpifgA2RrsWGmLwiXwZ0purn8P7POv74cZQJyqoZ
a60b+4eRhQzGszpW+z7cROmetkwJozt1/bvvaAf+jJ/mRgJbgHTAR67YMQYf
4qCxVAyo70nx7eaWeZbCNoMNgtZjKNrc0OSyq+P8uIjdnJKAhTmY+VfUrHd5
wVgkMYXYPHnol8nqCEMSFYxg9J8UauTnWcm8DLHr9gFQhwJiCPZ2nemhlLsm
+ofbWH9zWMXkUbSxzeAVV/LsQb2ZRBm0omHXSCszUsClog+vgbb9FvcPdfju
UL0FXR/XN97aqOjO9iK/iy9xrfTpJitr/fjNB6DNvC9ryRHkZZEEkc58QEx7
ckLIHw/AGuqsYwE27x6cd2jfPKPSkBIudowZ80+dUQxtM+eUPsQ691iatDHZ
+rp6H5V7Cp3vi4NJZ+cy4cq/tP7BuhTqrss/b3K+ZDGGhNj6xuK0Cx4Th4o6
tSoHAIXe81MtNknp8E7e7Husq5LLBFoRfeRJZZdZAmf2cxJObR7X26EAvMXU
PSOiajVeyNOvdWtY5M692GqGhKb5wB+rGbmrtCYuAyXovXR0zdNT4k6jH8Hf
OIpLsQFvrTS8rfPZWIS9OD4Vt0M8DMbpo7upJRqulEz/20ZLB5H+6imbCdb4
Y8DZT+HAEjoRqWgmY/5DUJJGS36tPrfaROY0NWXarqn/7tmsUZxmFpxmH0DW
VBkkzKWeFPD41PDGL9u01YtaXB1DFfsBb2ghAVit8OPUmcv+ZmNTSLi5FyOw
5et+9zcQKmBOhd/+cYVnM+2wlWtTCmdRwv2ydE8qB3y9Q1n4PM27v9YNQqCV
4Qrn3AwCG/NmMfTP7TJ9AyOuZy4XYv+8lNkvcfKMyM1WI5FhekyN+g8BAD3u
TKI66PyKJTJm6JZ7LrRlQ6eKqkxxdC4/xL5jUvURlXg6M0dNQGui+BRQ7WF5
fsHE+aaS15brlN8Ajx4BWp8cQlPhsPrwsc1p/BfCyhzJxw++EPk2U8AMSJw3
H7f91d6xhX2AwHrMPlCElACQcqtyfS89ywkSkMv0CnSWp+TA3S0FOUY2j5b8
oMW3UXFeVfyliWah1iA0Va4CFv3Oxi14XLPYOc7fglAjtl7c/Grw7pyR5kg3
+1cqPTkjAs5FtF2J0Yh571foWc1BIV3/v9piUmzQ6UMI3A0UleowtgBrWHtN
Vzr4ST9W4BIgpJt9LlUGbskqcip25kdY3XR/pWAjDTiwcntybw26Cu6DD6Ct
IkAYi/RL2YKG0wq4urL5elH1lta6cH4zOPtjbEFSDEradEdj58B/+Mg8+eGj
hmuRgoSZm1CUOiGfvtcSgFQJ1BrqAFShdM5GvJoQ4Xsqd8t6R13X21u+kxSn
wM8I3dFXnEv+G8Sw61SNqHHprXJFFaAFN+jzG7cj5IiVjy/K2s8L8qDkOtSc
eEfeqq5pp5610WnhEt+iVcEknLTTAujl1oyVOZZ9ixi90MmJMGtruOllSAil
jdDAUDv5dEB9GB2HZQ3taLF+T3HFtkgl4TxAiR5yHrUH73Hs7gQRUEkxzeVr
59Lcqx2Wbh67zWfroUd+3z14BQbEIWvg5AAJ7DMRo7excHGT6XU0WZKjkOpr
iO+LwLRU1OkHLTiQZRy8ZGyFqKdOmvKdq3187hOVUBxpXnyOTLwDQmEE4XmA
1uHFqrrJzlr3H22bAQgOqp/A73yc3llGvfj8cTcHdETgwMDXWmXMkiMpsze/
buzIMAHngrmORRh+KtpT+ZaU/C14gsxoiKnaZ2E3kglAhAyjiSIB3/kwBcar
NMc9UjOpdNQ/ZyR+VfKarvp0dXVLgEO/xARO50gFBdLu/cBHZnG9cj4W8EgB
CEqxkLcrNAfhnDBxHzp3jbBApEpjOTCcDJv0cdX6QvfC+cHIWjxwWNBh/FOM
bU7dJw+tGAThl5UWh8Ub4iocM/oCqQIana3qHv9ffmJ/jagt04Q21iJDVmLE
ERtl3Il8w9NznwSb/9/7wCboRJFpCGqWzF2CFPQ8f0jvSUZmfk3J5FH6S9lv
aiv+FHwRhJDOeyG1UwgSCYQWno98mAl565RROsoocj0xOf3EQTyLS2377xjG
Mj/cy52lTHqn+IyP1tlNI4LneMHdNi17UdNu7IECeCzLzrRw6SwlNfpDmMJK
kNfWIK3Ui/whLMvkzaHe37ZyHPZhz0wfB35MYniMPkMZWuv+Xo5+pKmiGHQR
bjruyZ1hUw1HxdTCHE/5qyoqSueIVX0W7zSx7inrrkqEnHhZaHP63Uhnn6zC
UFF8pPzcRnPqaqjVCG+DR0+GTS68cdkyXPrC1FCE1b1vvPZLzKhUH93mnGox
EiPzhMhfllBOa+/Z08TV8rjlDpLCv0xonbZyO40eoQgYrXWAMoGWlo5BFItR
uBKn+snSNaXOJouJze3K7eNqzFDQicmP5mFFLSeUj7dY1shrl9jyAPp0ByVG
mVP3eT+LRCRJECeUsLn+MUxRUvY0vFqHkNOJsr4wzpDIEbNa3MpuskCxcV1E
rSjXpModVGZtpq9byFjkAK7uBTA2bACmY+BrnR4//Il/Ng7rbHy0K6Y+frt2
1MYHIt2uEVYAbjK9frjpMzN7Oqkh7tmxn6CfMO9LGwnIx1rEoy+G3eAI+jx8
nhAZLF5XPAy+7Dl6YFV9L8bxSuG9iR4cvDzXUSagkqJWLFa40UTwL0MmCbPd
IhG0oiNeEsxgiALEAd+KbZh28gdt2sAGboEa0JcVooCRskukUmM9VUcvVLgs
yI6TvoH44UAdZ1KZzfd1AcDuFKr0zhWmjZdqM0r/c6D/FJMqGB9OcVBkuaLR
k1WNCZyw16G1W9PMQhEJuffOuuaXg9PUWweR64KL/5QB9aQeCQ6judmjlJNj
8lWsFSpwxMvTv9E6RMXSKk3MBIF8XNJysBT8FWyqxGCBrTQZpqgkiQkCv91f
Gp8ySDXJG7CjrJP6GPXO1BaMnAxbLdU1fdh2aMnBzDb5z+xJjAIrPGf2fujv
gZXUszD7dBD9rL+HzBLIqiH5AomRLvKH8KD8smiab9oZXdzZmEbnq7HL3aoC
mDk3oj6W7rz7Wl9otpGsHWGfIfBuuhhczf0VcmOl88NbqauPnMzm80vhmzGI
kJHvbWBd+3aVICdOqH5YXm0LHealGQpAwciwGizzUs27IiUM9gPqzsW0O0rW
7J3bdX2dxI3NLwNQdavM8UrMjB9H5/oxaQfWOvSmlyfvQWmJOnzlQgz/UIHQ
ZVBo1UeaU9shXlUhj+Nn1ZGZHDErUgWeQhS8AtoJnx00kpmlW3y681omRMZ0
O6SVkL8mf3NJFyj+cWm9v10W+iUhb8ej80VTFBm3Fxdd/Ebw0vRHk5rJtK9F
IjpAvj36HSnAuSTTjeugSmVqTQP5mlvbFQj5dzXtyLi3wfxb5FCWdWkgJmvV
lqbRklxIc2z6IG0N8I1SvTlPOEvF6579k8IlCMjNF/cdHmPoHJS9kJa7zhn9
i6k0cTMPz0tbRVCZutrXgaCrAi0bsPXAp8W4kduCXtRWNjA+S33y4UFkBqYz
yW2BCDQmqO7DWksGjGraf8GKbtYuTu1TlFTN0uK8YALP1dFp9ercJg1uGEpb
n9A8NmlNUHglzoAfP6H7hD4uu7HiL02enrjqBat6JrBnJN2MeM2wWHAoDhvy
mPamW8Oy+5jqam7w1VvsGGOt0ocXbCaqWKEOXtr4GJ16Zyl/A9K6N/WXcTe2
ziNlXzDY8O4o301vZioj9nbKqg0XC/c+NqP1VK9CED2yR2jWW7sVzNkFbQBz
s9bcQzNwV6s21X+wyAMh5Yv1HKXx5YqNBsHAvsTh7iO3gvAG9qj6BhQY4QaR
Y6TiOchzAX6VJqiP7jSY4WviLzuEHo1H+ozCChXzV9HUCyDROk0EHvFlaVJq
TiPGiNRAGxeSn4LmwxuGLKwxny8oCoHtYh6q2tGczi9GL92F7mDGy30ZhEBX
rS2Xhz2hUcjNa67rY2pskiu3ekT2BEn9O49K8IYYZp2PtB+5osJEiEA3D7DP
UYyb69W3aqP63mtatMTZLw0csU+MSm8eviUWvO+FHAbNyvWLfsrjZl3aMw6p
gfrvHikVxFv5L9m44kp25rAl275ztuOwmWBiXwVSu1sRbT69nEZWbOwVNLyt
W9Od8kPx1vLv25s23yTwfuftUTkPr1NKEyX3nQJk/294Ua1qqVYnVglXs9+X
/gT6Rx2OSguDmsnRTPZQtvgCNWQP85NNwJMIdHivT6GGmkoYDyPBbKYGi2W0
YrfN88OrovXTqhPsDkH5P3vjiWX8lRyP8JPXLsptoJ6UqaAqiL86GQ4LzhQf
UAdMWymK1MC622nS8VnCaHQwILMSfC91Cwj8opWAXV2ximNjLehU4hn7yXx1
oiXkucHUSe/IclnhlWbyzPXsZacXebnO/+e/jVXv4wXxacPj4VAe3alh+rC1
sVUhdNcvgmIp4GPKaVO1qXpH0qZ2HSSdsUGN0C33jyGm3otg1H2+zbBJ/cDi
UrCG9fV8o5ErG1kXpQ6GyNT9oyJo4z/cjeY3AG/EPWNPaXfobek8mnHSn0PU
fNm70wbwW2IHFT1pIasKpgAytfYIqgoD4hxgxe5HiICBfz9HEoUn4XUkVneg
Wn3WYYKpHTNOec9dQJXZ/nigmr+tIfy7TUQw+B5Lb03kJTWDhOOyLstisGnE
0lWfcO2y7wv2PoXcEL0XDuCjVYX5mjBsNgVQ6iBzh1QX6ka+oyTAvCpZaPu2
DbHwSPYc0MHQC7K04bfjAf4c9xV4n1YkSNb58L8WVbS7Twfa+c+ekvl8oybB
/bw3rvMSVLBDSXx3nbhTThKAY21TJDcQTVBW5ZxVvhcRMS7QxxQIvGS2+p6B
mAMAc4RxqKGgOP3ZxdyDx8ao1Y0QG7YdXmNt30yKcwQ5Rz9C0uJrB/DY5FyL
VZu91ykoKmicJAkkufcgTn2EEL5DouzUterfboRWNVdjkJj44ockXrFUcLL+
Wprh36kXQY1ENN8mvKFpUwBYb0JB7VRt9EWTb63OcME1MUBrGnGLL7UEe0nV
rjGhgBu6Q5OPB0fga9dpLwj7RGdkKLpes5ZopF7Zl2I1HAyIXtz2HjTrcsFM
Yjnp1+plY8SaEZADPyev0mD+dhbL8ZC2LWnZjwuP8+ht0T15vFj55+qk9lJk
HKdOHeepTesYqaLUYnbjueDBb7C+Fz5i3iF2Xcn0UOgDzSLoODe5lYJjbU8G
QSVSlVIRSRVD7Ep5qQnMNpRCytCeGfwnumtyi1Xaw+bLAhZ4/2Bo8j5sPM+9
YgWBVlXsavt8Nk61XSM5bvqUw7CJPPDCndK0GCnTPnFNAGS1T9y8frVKTHNm
YwW34vSoi8XgtuDiVUQqlOf13waUVPVM7X/6UMzdBVekp4m8h3ZwxSmuwmbl
Dboh9SIM6hq0ztjdblOkZRJArBNC+ZmEUS8h8CkqhMAfEWnWXjLq7O+tuB9S
zTX43GeyUMnyYqTTgQfAydQVl+4mXzBDjgWZkNQ9+o/quVS4YyrLbzoQ+DbH
5vi/DspEaS9w1Q0Fq0lk8WeOeHSILEJxo37/+yWLG8rLDQKO/yJPKIqJ5Jpv
DcHaRSDDoGcfyxCaIIRuhCLDkPMKRf8oGFtQSX6Ph4Ej51VI7wdr8UTY/vOQ
DxmXwd7DH63J97kTapsNsish7TQfBy0yzelhecbzJcc/4v/WRBOr3yy9rWCS
15aY2UlI8FzPakxXXAqH71VyE2vNjD6VRuDdfWlt86uV5HvG3aXMH3WmQ1BT
dgcFXEoUXgxbVLS9atdUeeOv0iyzEo9kctqUbPMyml8HadHtAva80rMHiNHt
4ix7/vFTgbytaG/OoOn6YL1IOOg5MoqYkpR9Ej5XdaWgsAHCSeY0PhgflYYO
ePnRt/XwSlv4UvlJJFRsSo2DSqdW8dTu5K5Zs+g4lDkf5y9FJxadxCq06p5d
YaCQVz6KdxuVSVCdgMpFqTnmhacftPF751bilWgAUhRGtMUo7dULji8+Wrxq
hojcaoxP4tLgOzz31pWQMlTy/lUxt5di9yH1i7pbbS36+ZZlbwblzxK+lQW4
VhBRg1Avhmdk9gSh/+PzzDzTqGDVga6txZ9qGZJKVbBfA6kWHoEyMJzgGsk7
dmrVSb0skg/FojcCfwDMSrw9jr0acOT3aV178pW+N2hKlhWsI5sgvMOuN7dS
uvuEWl7iDRLUli6N8hJsr7DCQX4TfgGwZJWL5hB50N9DStDI4z0vQAs8wj1y
zpAOM+Cs2jY+sUbvTx59WaIsgUlsOLvyImpO46YtxBSDV5VcLPTmWSfbhh9R
xIsZKE+WgErExPcMjPpvfPRcgN3sOf/13QEbFIECZ7l5zKMsWH6CtXz2hrHU
IfWGE47/aL723dUvtLm6IZMoco9/XVQiTh44SskocNI6GedvQN9aWbkLKW8o
T+0efK/odFCzhbNTgbt2ScKZis4rg2YTgDH5V6QQjuHjIyigpGKLge65GLDt
ZNMefT2VExmnbB0dzKGdv3zNneqbPDEXCP8P/vyB6Ze9UDoWMsix8vp+Cp7J
5e3QZn1/dZtxCniF1uFFWNJ5H3O23DGw5BOr6zKVHDW3dinO5+8U6ePdZDC+
ggdu64FD2yiJbmSUC8TYEIDJy3xOY/mkiqJBQkwr3XSEEd2kZ19Wa0NSXs9W
2LQyZfmef+v12lfr7ocyHjfU0eL8fHTfYRuHOCuc1yPltH9ATUtnGnavwHsU
R3Ls5TIiXF5he6KAtfKeI3RAYuHcMm8xQXTj+vMTlFRwIsM+YqCRysZV/C5N
hI+vmhGpPasQrNmixWlnq7Ra/aCtYYRpyOmGfFWJbYEI4XjG51/gkNcvv84x
H3CdvYlUjoGmqQcWfeCckEcMKHOuSpZ0MnI7BvBq1YTBTPhkfSgRGcJHiPqb
+ZR2L+BYWCMZi0Ukdwl/2BzVMs8yRrPMfoxn8UnoyGqJZBkPZ1M1hfGgNi4V
AUxmldQ2FsxJRRvrrEFlJwihM+Ld2maMLckOzhhFzkA9BIFp0f0pS5lNqrx7
DJPmfKhxq/TEamGD9PCd6Hp2kcoITvGSglpEYfhqZI770+WXQ+GzR062D/6/
TVzQ+R2JG72YilYwJGsKCWiZmkm7HVWPFffydTN/CvSWc1ei1Gfjyy2254cA
vahVy14/YLBytkIcBUr97IpOo1iEvB/78AWU9ltc7mDzIBUvLKVOluaJJA2R
lnQP5MN/6AQoDN1c9dQIJgt6ZHTbcztfU0N5uEIo1DBIz+5suYeEXieTUDD6
CU3mNSk60gHfwvSdnujOUBewYxZu/zGtId4FEbyqKbDPgDv1M/zjlkFdqVyE
mdpjU126hVQX9fQfUp8u8fP5GWaXpj8bVE7JvZvc6yT+Oi7hwq3n0CfiVLl2
DXQBsQujq+wSDDLT48/v0JLEMSIVB/hMYYg9O/Z1NQ5xwrqE4ySBNtiM0s1I
tk3fTFiD2zqHbzrtiI9J+AVKvNfjXCZm1Uw7q9nnEctbvgCFWUr2Oqpg/RbN
H4ypfOYMQNwZAqqdv9SJk0PxaZtjo0B/Wrhy09tRMSh1B2kX/OzRBf/3SUlV
Y002wM684mZVpgyE31RdE6/EccKU4niKCtVZ7c58k42482dwif3V/4sOec2O
vF4RyheaU0HwiVyfVjyCY2JAaO24MTKTJ844ZzjF3ilmXsMjM9hCd8Ba2mqz
/NC/pjPRCyuaOuySuiqnQGju0kGm4tfqxFGrY1OW8iFbmvOi7eBHZComQOIL
cQWxA0HJy1m0XUTzrHerUFGzgt1JayZY2ZsBKVTeVFA05Zq9DJXYVHl4xFCf
dKKiG3MlvwLuVHcDaoKLJ7VNIKatxr6PB88nKqtNfS6mgNy+cUPHYOtXMRCk
DJwGswIupeXbKtmxmw5AGVBidNGnH1HIPL65mwSpL1RBYKTinJknO6S7wZlQ
IUeuXW9sQN3Je6bquOgyN0WSR/FBRjUnHf552TlaF/CfLexRrES5SdifqdHw
pnrzOp+SUetdHQ21R2piGF4zMhYT45nZfBMxNkW7mHBc3UM+eEIfTGVAbIrz
BiS3hVJnNQwHSnReACO2b18FrJKOcy1mcdzvnk76eR6R/r8PSYp2gmMFXrhU
cS4/k4k1eZmLLGS7UEX3SdgyPfOMJqYm9Gb7nkV6u2++bQU/zlu6L1PjqOPn
xvSje7ImHO0C800hQPRtUhMVXwxWbzLS5cOJvVTLqRXigCTEupKNe9nQsQp8
P0DlPDYXDWbh6C67fNypm7x1U0MuksrTUNMsbwrS+OqwO0IDV4OgqXeBLz0m
OeOrxC9l3m3pjsvfXfol5p072kKw2UnpfQpvgB4qIS16S34kRqq2bVf1j/C7
ZcHHlw8W1P80N7mqQVSQ5amllhGvg22/jbIcGi1RWqX5Ikvjf/8hOS8tJACg
4ppa/aauQg0uLKqxGgmCcLDZCpyjdxkDXlsVTlbiubQGLhDJPkI9d6wBTxw9
uxMyp2uDQcvEESbHt1N/+g0jYjrw8UWsuj9nivmPlT65L1/7XgXyw8kYHig5
SzWSsia6ghAz06Eb8lI78NYBGjrzFuYYv5ExURng2+xDNF76w1RHg2X6ndew
9UuMdtD80EHxNw6iqyBGHt+Fp0Pr0bWRvp+n8RqvnFRNVn549Pozi7fS8fX1
LE9Jo6S3NslrLEpo2bwFKmbunG98lHskkYXluS/niHweVC24uyxCTgnUHCVF
yrBCaNTAWUcW6InaEpdE8W7LuZBye3/9Kx+fdAW+tkWlPf6ipFGrfl2uWA4L
1o5wbfoM/9EB3D9mnGmblFCYrq3ftCbReW0dy8klAXewQw6EW1evpAZTyWGA
jniXNU5k6Aw8geF3Z7UQnKJPEeMQ06401WTRo/tSwW7NJTYPRzyOtlGm+FBi
qQ09rbBUMQaLDvCdnd4END+zOHJTtEQR8MvhRZI/a4hXhTTMOrk+OQrQdjiN
l6TKHNTQPtWU7hMY/mqPw/riXaBsxyCm0MeUXBSYyb92EIswrofNHWUvhhZ5
6tYiYHRkX27K91VFDh5eJCzmHKOQaZIAhBiN5S72/RbWoBIrM0Muf7z1jnQw
iv6aelyaZel4OGHw+7/DsQeU9LdtncwofoZlmF8irkQh67jDvuyCjWBoKj2R
S2RsIOUV1LTJ1Bpyqs/+CCuLINhmXDNl5dYocG3TNOjbMTVSMsjiMIb99lG/
gr5ljX8Im1pImjnBAypUmg+X+P/IOwGIGopeVzIgA1wc75MDOxi8YH6Wmjdt
GE5T9TKLXlFc1wJmyWplQT49WbOgqcgDZOvFBFa9Neh9QBbvKFQ+Mlx/GfJM
QQHP7wyHLm8pF4P0Ut0UQdmy692YGW/vVkTUj3EcX0GgkUBZ+vzRzSspE5x0
47zHrO1khrV40PLwvwZV0s7uUorcI3Ss3VkNQTZpku3C0RoiXj2uEsS2Zae5
7zRZDwwThPLF6cC6S/Sq96j9VRivsJUhKCzRrsvWw3lMkeJ6yx3rwbBdiliy
QijeXkYcovxRNozuBExoazALbjzIFiaVJtOtnlvXY8ddH+xCawFaSDEU8AIc
MoCUP07G3Vg6UikeNM1fGDDBEpKavuonXTcU07u87rZYUhWz2Fkf0YzZOJOd
PkdbB/0GW6sqNeJACgR7tNeLFVjdckJ3Vf/FAO1vN9xojQ8L9JvtjbYnoKGc
68kf3yiO/TTWhpK1uvg07Msf3Pef2V6IQhOmhYIac7nmJfDxjqAq5KnzSPQh
0OG2nClNSm2iCdBlMx7z+M7P2yYWL4fJlGsznShybeLA9LDEdk3znuzOTmRr
Mct08KTaceY0JAIOox4rqjv2KbQpkHMyCn7ZMVoZDS6jwM2zfsCVM+iIInLa
gQF1S3dmZufR1qIcJYCbycq04CfyUHnB2/FMK8g/HawxMHkxGYGTlxfCR82s
HJHDfZiv3Fnow6Oa6z9eNmeCFSSSV955XlqJV9Hl8kH1EiI0SG9gb3W/bfmA
jJ8Y+lejNY8MW5yivpNoFeUdvIr1A7SE06LEJa87LmisNVHI+FgJJkHkgtTx
nkvcGLK5r+uAdSrB10QjGJN/E8Oog0fOVpS89EXpbllDtwsatPdQ+ubHDQEq
FmrrL5NR1Z+C8Cb9LOcVBuR/giKYi4gk4hfYSZ2tKwbabz/1jZZAfK5hAui8
jCHRu6921PGlc5+Rqwp5ilJ5IgNrj2lJ0jeLNI6FpieY6AOrPNFTbM7q3/pj
0D6sYCsvDQQzL3AnGj+SpWTI7sysU8taqkYfxF/q/VxVKPILcyJ6Zw0oNd0G
3ZF8Aw15u+ZaxYh+c0lzVAR+TG3wh9HvWo9IGPEEmzfeUPGeGogVIhMJayEY
D7bZKJIGlQqJ+GKp25uRiKSvbwzPJRieSL7cB6qFajf+zJoqzeIJlMBhdgBg
i9h3P7c4IVtV6YokP1VS1JlFe0bVQILNYJ6gGoYOmUWDtlEblaSzygtSdgJB
QQxRJqYhxzKXhZlleozX6jVvwFgo8YgjZaHP0cwUW1+YJYs2Ig2JtSbnlpKL
Sxgtw24JOvbE9dsJcWqJci+s+3GYBNRo80Utj07WpZfR0TX3dueOQ7CJ/Vtn
Y9KVZF4HF9xJMWky918gSGvwJIMbQhhkMPvgjbrIp6zALXdbKA+qSRVxJsp6
9sjFR9ZmmJI1q5Lw3Wc3D7a1PotdEu6GwJGyEKZ5E8EcyZl0dbLmUMMNuDrf
5fg47QRoBPSwj4OWdmeO548fQ47pA4WHiz0aUfde0C7afIF+zqI88egobs+X
OE4dgP4yuA8KrIMoTa8KOXiejr2+l8Y2s6Zpt580zQy1W/2cKPlhr17GAbeX
Iisshdsj5vIHXM6j8YTV+H3qAAt1qJ+Ff3H0sfExmU2RChWz+Z5p+/w7IdLk
8wxdeRxXgltfp5TYMYA9cp3zq5xQnQcDAByietaozi5IYTQb1/fXNutc5RZ3
Phf3a394C+RjVlGV2rIjOSW+940VhczR/5DapKzCBqhGW2VIEsDD9TUvqYJD
P5bz7aF9lBGuyOr0YOY8p7yoOE9p+MKLF1hZTtWPEEZOeVc5H4p2fdJva8V8
O7zqRTqoFdkk7SxUat7tQ5tH0G6xsfD/HgmK03b6AfB8JE020ydsfLxgafNl
NUrSYyc+y4NqHQDQ20iXR21hkCJPzSUS3zWr0rCdFrWHen/pgwdEvz+f8gtA
FwLLecAimmWVSGkoUQWydd8nvL25U3CXG6Wr+Bt9/EvmEY7XyqST4d1ovr3d
A08vUiFjUfAvH9tFgDUX1fgcZKdYzLRMBbk+nm9pjA++FVrzer+gEARk6xuv
5IMIK5STpgwWdJVPlaSMh5kLPbfp+06dV1H1UbcSsa5BUSa7hcWTomTcW+IM
em1nkMysDZSk8B9MkPDT1OppXKAbN3aCjE8WXC/rULGmmmdH62KZfVm7ATe9
6u0vl2IYxOYBgUF3ZHqpYRqnEzJedFqcnzCp7XemaPevZU3qjnbOHxlC24I8
C7IS/ANhi/DZ9umfK/9A54XFOMPPDRtnRLJFlXyf8dzTuqEEmh547UMm8Eue
JlO0fC8oywcudlJbbmo/0KM6DoMY0WXH5pBVrrPB2C4bxOreYrQYw3e6TPLr
AdLqQRZi9NoFLuMIgOUeeO0Qmr6s5te5LQJ079bJEVRsHVOXr/CnFrPq77o1
cBpu4auXDF8qq+ghY1P7/FTZ/vOVOyJA+6Rdbb2uISVuyA3NVWOnjM+vqCD5
Z3NTZtAcEfQde3Hm4tuMFpI2rpW9AXlfEs1och0qzYSyQFOnnabf3brzQVi3
xc7569ZDEaZ0yXY6Oe0piyjwoQY1pRAWX74KxrBCRXQdRfWGBIvVnZXHfKM4
ttinSoWPn56EhLr7a+UvDcJiCjtoQwxZzwkw8u/KGP4ugwyK1m80P2ylDwPi
heZVPaM6ak0n8CTsV7Fb1xvk/BqRZJRYA9eDJUmjJ9j//lgH/lwhtd8bJDZM
am6U793vA0JyO54/F55tygIc50WJGMdQK3Ar5eA/eH+r8Cl7x4hlYD52GXYo
DEnvXN/EjRtJ5b7bUYtufwfnEB1tLoASIFTzKGD5Pm5liFEWA/vBR6g9YQRv
JqO9dCALfRw5pGRT0I4orya12zWOOKaNZAtz72xtWl489ZltbTyq/XJKpbNG
xHtldjhOYTdqF722naj8YoteaQpZdYXl4G1f2inkb1fJEbfsyEaCf/iftqIm
5Ivpt8U8cqmzGjNUZbumaW8xOPMCqZIO4/l3efAQ6mNxzTUqXHNmVw/KBpNr
FUzgHx1ZJHcKDlO1OvUkFZJdTDhD6gXlavcz0GtFe+0jKCc2/rg9+G4CEsQI
Lw5phueISzZuq7jF8PN1W/AcqbxYUkbJnplMDiXNKDcS+3l1Dkgn3f0Ys6K5
98LyqRk/qC48b0VVfgSdvRAqIHyEI5CKxjuJ8NZx4HlTDkj7B6w6H1tyLQuN
xzCMpkLsOPh5DmSiSxPGWjbAVtveZG2s1nLGkYpm4DSyh5F8Taw2RCB+nQza
edFivXh0JNc1ynMkvnpATCqEoBHcHcYGbSKf40PTSI0cs+l8AMF7a0zbUksB
Kweymtor3qH2tbIhnJjZU7zjB0yk1TUuY7OfzXE4rxw+C5J67akbghJtucUA
Pz9QWP7b+L2qq8xPsUWPE41e+nDKKFS6D5jv7PEH7bPazzcoLZmVsMCgFE0R
uCm/puLXVwn/U9Y3GK7YFgquaNvPR0k4IsjUl1VqOIIm//B7dACC0xcji8Ji
4CidhUIZIZ2AOg2y5SvTj/Aa5Rn3dL73TuEfksTUk9qTXrtY6D3H8LVI7AZr
6TJkgQTNU8w40HtvgDbEf7/8/2V5EM1P136ibXA1vcEf9JzZNH+IRC4a47Ma
SMoWTpcG1TEngn4cMB+Ycg3gBWOHFTZYMlebNVxuU/PEG6mXsDO3iuaR0RKO
O9xRh2rqxPedzYbsZzyNSJqX8K2U7Bcfc4V+Xrkyf5B0w+SUCvv9BrPoPwdy
AvADEYs50FM6zSxrlRlScblVOPFbgOunyoQO++T3LF3w9iQLtKABEpfFi8x4
ocbJr7c/osM6ft+IMRoWOFaMML0cL40yyXAlYsmnMfQjEoz6BObIeRnB1uKG
VJLErE+4F4QqVsB4m49AlrFkDf/6HdXJzTsX9sfMUwFWOoroQT8mkZ8izW4f
m9nfvHSs7z+ODgDeKWS4yKCPMpwEKUfrKnCQAKBpXuAh5BcUKI0T/sllvh3l
EWnIvYu9Nio0iBybHhTzbcWbE2KPuN2oOLE/2QK2LU0pK2J3cbs8r8xP0md6
lurJVXxkpgAB1mQ1/wyi5uHvAaP3ANWX/vGrizrVRcXbdrPXxBHX2u3b3qWl
Yx9/j2vupRtIrmYR7Yvh/lpKrBkzCWOYjD4mnuhKocMutdQ0r+B6e11jWhde
eD4tyhPb/Bs9D2oxweB3q76MgAiDouSiopdtcPNGu5mR9FHgMNca8Pq2kqJW
usSvkCCli+OASw9Z1DrJrz9jpP2kYjFimR4HLXtviMuekA47EYL6018E89t6
Ui9EfSJKmp8+vnN2Y+7AWGcRHhWNsbU83mnboEter8b5FghPyxl54YXqy9th
nsPaGp4/nXCdOA9fr3TH1eQZNlPOSa+rSDukAHqti66tPIfROlVUPlCH4jMO
npakbTHWve0/yCEi+xfmZQT96CCYF2swftZwiVlWH7jj3JSvGc98H9GU3PYQ
q116qRXG7qe1w8qLwWhv3mAAV0lQREnFyeZycN2Ztd9wIFevFBUz173JltUD
U4eIU81s4PsFs5iuFdZvhdE3BnZKgS3XP0I23pY/CYvU1DgSueKx7L9qZYM8
U3WAcMiXFArLmguNC3jHHeg4xIgfdCkFUzsCi7a7XADAeXKnMjYTioFLWzrq
UVEgv5HQB+JnVE62WaCCu0pFwBMBsAmsreQpud7YU/X5mm+uEKhSI1Xqq32s
cuxQ02tSxWxGSnHTpg+Bc3m5qb5XoahXKGCydq2T35d3Ky2T7v5qfF0ZL8nl
ZbWlQ88JEt3/4skwqyZcVVj2fra3Mkod9EHj25U3nMeV7v/kPila2GVfMTe1
mJ2yHv0+wJ1pu7ZMypz0irXHtKIZ6ONwwxLUzQfwoevzHvIB7cSCbtY+7WE/
ovQn3559XRug726wY9sQODIQBVPC+urYj78n99Qr47jRzKl4tdkpYb3gFvH6
s/lQrTAqUxZtmjCxv5OEKloLr4MYLe+P+d1IQusqCh08KkPXsmHhB1TpVCkY
VjZU0dfPPDus2gVjhzjxcd8zSsn1ayyyy9kOJwUopQYzwcq1YGVb98UgvyIG
gCI8BlTgcPbc3jtAW6GkstevvW9xxsehWKwqIl2/duEgis37v98eezG7sFCO
rbzB38yt+yK45BO9jQADGrhwx6n2viTqLCteqcyYiJedFdKA8K63OpJy9+9g
Z4XZiaoJV8bnBCyAcChVvDaUnBHmKRfAnzmFq0drplE2RZZzWAgR9QT4nQL0
CJAcSphpVOyveY0xu0Yxl/bjX/2ehsU38l8cryxBcaUc8WF5goIFWKFYnS+I
MZc0cZDBPOlE4dVqbWk5s9X8nVou7K1u/aiD/2tt2jj/iOOQ4W/q/PnX8KSp
k1Vqsrhw574gmJ9M2/r9viJWf64ar/AmONDCwd7vdxfDpDhPV+4iX/0jbSH5
75slZIR0mDwnIaNqbkClC5XKcV3SU2C9jhzPVk89U6RLzgckJQbh8brqLdsz
BiZKQ62qtLpIwT8hGvLl1UvQju8NXyAJh3euIUIH5XBGNmriJr+XAAtuBPfu
GRh/B9mzRLS8aIkS6cIx7FicmhCkID+osFo2EgXavVqZuvhWi9ZHpuXgQUPR
TR30VCKVAP04WzLmi3mrK5t7ZcNuC5QDkzkHBbLhqAkuOMUAe1b2nirTuaJ/
UFnQnJUJt43hjZ+R1v17gXd45HX1URV0ZWIY4psKyQCwwxn0lInrQi7Dhi3C
NnXGKOmcl3jGWIVLw9dQxRDgjYrGKgvFikoLyzs7o9n25JXCDZKmQkAh1Wlo
3naO7Z8CqOH/pPagflrxaj47aBuR4sOmya6QEoifBJJ6dAKJRISVxY9mIopz
na4nHrMeFjSripT3tqyM4eALmn1vMfpjh9DRePquKtBCbhZHvJBmZu1JxgEe
c608qqgKVLc+0iEYqrBEdu9XhpZuW5XHoFOSHI6ixRPtuyb3pRM3MtyTJpDj
uIiXvahoIWyMfEWetYM22x1mvT5vPQ/A/mKEX1MZimDl5zQfzI7Os744kRCR
fZbHnJnv77Z98QcInEFni1cpI9Rbj6EipsbgvvwtBDiI9zZRcGzD4EpEk8J9
wt8xK7KKnYkB7Xv0yc0KpB3Kfqf29e1dH7rgA/KVfDn8DiR/A5T85i/lfSb7
ksNU5H8gzVc2ah4o/NyWyJfDKRU6L3xFl4a25sKBrvWu2v+fhEY4o9r44Kh9
uqqIc4/97aGIYx3Xk8tBB1J5zacQzC1SH8LGFR0BSNXagJFyk+DB/O598w/h
PxsAYftnYATqOjKF1hxO5Rs6NjvCKMcXUlNPf4qwQEt+Jm+kEbEOjpguhweW
9QEHDDucqmYGVckZ5+3oHvZQLocsRSnBJwunhqnkbKgnhCUDf5dx/M8bEXCe
6BlnWqCQOTiC7vKecE08FHY9kD4E2J2XbMT5Ar64vxdZh5WUQpXPkuyzSlLq
3PIFBWFB5WK1gLxYwRDz6OkAd8FdUmabWulZ3oonU0F6Jbv0+M4P4e2iCnQB
HGzBD5ZiITa6kEJv6FX9VEnGwnXdqwX6F+XiWSaaNC5Y5fpe0Y8eyRKdOTAa
nM6DmUDB0T06qnTMwg55fEo2ahS2ygVWWDWuRPyWRQTkrgZ+5tfv6V3Q3J6d
zdgvf+Y91N52W5wQXGMRPRQpLoqT5X78fYcvgVRBEDnkqd1S9ndDn7S2Swty
f8gRxN+FcwEB8mh4WchKbgvNXHaWqGfdoVhkiYjvWt+iw/vcorTtNn9Gksdh
UnmmXyhPBH8dkcPU1hRLhadQRZh0Pon7Qb1S/6qXNqZJvf7clAgmbiJvfxG2
YKQtQvnWgHeddJcaztyvShWee5pjB7aWmcVy9Szs2xYcFqXatxPGsuqb7CBX
oGRL+NKjpXnmKNMm6b9Hq68GgLjWi+ePCqEmjDytMs0TD4U/6PE52qtVu+SG
azA+Brsr9BXQWjG3CfAruQXZDD2MkGhsQK7X4vqVNA2YqLFxhUnZ8mfFcovt
OAeHpaGSrB/6HsRACpbuKx5Phm2x1ResB033Z5e1vpX/BSuoI4xhkTDYmLqR
+RIRduDgjQdGazut7GzBj84/5E/7Ww0zIayPNuQIQRDr8svS5AnieDUi4mRB
ky9XVqL4lBdmPNLrn2nEtMIl6dolmRlxVilJDr1nqfb0nbhgoLI7IWOVl+Qj
d1BnWvzE4vtpivwV5KG0sf5UlWYlpdvrOtQUo3k33EBpzqCaw+yXq7Is2f/U
rKJmSh5VtIEryWKiAFkfYcAHdMzT/8YrQhtSaH5QHhscxCbOdCLKgZPKyYE2
7wfeT+ZfReXOc1ez86RoIkdAaJ852E68mIvHlGdVz7V6UBHQvt7NQb97Goop
fPA/G9PyLc3WI9c0LlsGgpwx+14ZJoQ+gYaeB0MLx6tOk8gxfpQtK4b2dTKi
igLrDLukqsTV4jylbCSe0oia+r3lCa3AbD4GOPJW45zFc/S18JzVN3dMNrOu
ZjLhIkEYJbnQiv5hiPGHZpnqYilKywh7t4+BZJerbWn2CowQQIFNbOCg34H/
PZLWd3zz+vH4jusmqoc1EzXX4+Rse2DcZV851v9E8ZAaOitztyVa1R7Zyzlf
ULAmxGU119jzWoNx4hQX2Kc5Qz6EisYKcf8UoUVjPH+t1Jzj06fvbJhCXNNJ
Lq5yxYNygVfoXFiXtr1VEHZDkzd7gW2nTkCSwR2Ldaz5vDrqTeYvGkYwXSVZ
ixaWO+LHuEDRTN8qP3ZbybJP81pz/gUxS53roNK6AuFIaaLnhRtzdpTZFqWD
UrDVq7NWBPwFTLsKtKFRmxXuPxvGHrK2dE7VMixOp19NZM94n763M1DOGtvv
t70EgE/OMVHnvtsDHRjRo01cA5kAI1N0jtS4FrZtIHG1o6wJ8k06Evw57G/7
t1ZZ1UTFs3YPkWVukIzILijVa6/GyuOeKs+qdhWweINPSx9Nx38PaLOmkKel
l33xc4DUqalSnaMDwvKue1BVzM5is/MTKuQI+2jNu336lRKqUyfzmOGspnF9
oWfEzB4iNmR/V70jULter4z7idnb7FCStrIPJSV8hYxpinOq1b0jVd+3QN4p
ZtAmTC+3RICIlwzPcYHkgtPAD85RkN/MfY4y7+RdKkPB8HB08Pexfxbfnkkd
AZTxRUbeAPSG6kBp0Lr+C455gsV1SPVhOIkjxnXh8v4VWw7csOTgkTAyW2uk
lEiDBufU8aJ4y1fBAy1JF6aZoljk76qx3xFWzS5no2ilp9rbyES1OxBXuJQ6
ZMgPyLy+WmWpw8oZ/J4MYtpZZegw4iTHSZaLEUwKum+4LlT1P7OPTr5PU2Dm
ObEel32WHtiRvGdEm8eEr620KccPAkOTqZBkZV3l8mkPXNEP3aScuRGbNJDB
s/6e3p8xwW8YfFQ7kO9oSD5+RuAX0LCY82N/LvRkjSf48NqCRXzDPrCUXF7+
PNxadI/UoMNSZbH+cM6BTxH2SyZRyS0JTU2Kki1WFetsZDunyrkb0vHGzAac
83B5BcIl0/P8qta+AoLavgsyXIXDLMiZWhRLUrjZ5p9LPN1wDyOlsYTL94DW
igKIOLx46mYNmGCniWmGvr752pfGT2Ab9FE4kLRfWVFartgXt6fKHuvfLYvo
tn5wE5v0u/7OE421LcepbMK79NLlKAMp1o26W0+fnDubJ+FpNXM/5yGjj1kS
vagffDz6rXf8g00VrVxQwqJffIYMIA1S3Wl+J2EqW4tVIjezXN9iPbdpQ5Vf
z8xFynFFfRPnS/X6InP4R9wOdERtclrapkgW/epq8MDpXnC5gBc/qY5g/rXm
WkXS2ORMQ93GkKxAcr75XHQx0TAd3jXrTyBby+UXez/YYE4gWt6+xHOiuWya
d1R6NuxLDv5XI3bMncJVNyJ8o5M70z+FuQ81onxasdWMpEqAjLNHBFNYWLmS
amVofjjH0oz4LCOWezOGWmCz9hi3PV44Tlwpy4+L71ybKv+UqpH4iVZAyISX
UV5A376M2h1WABDn/wM6NyOP1Mca6gftiVJ3tB1azxjTZRczAOJDTv8VTZbA
7pwV4w15C+xp0niVmRXmYnx1TFa5RsM9LFBfGM6b9l+I2dlnEKrscNPPwjyH
gCIgAYhxIjVTCCvPYtfhPuQn+A1k5xi2wVcaroOjaXQUWDlyr8cznPI3WDCq
ceJcFux7M+2gVlUogQcPrrpT/g9CggRCKKN0NdTXyJDXgQUD6abqn+TZgeoU
oPBlocq+EHeNse+aGjtM8fvX2NTlEu8ZXZuFq2uLG1rZvvRkLA+p9ujC+JEO
PBFxSl7qy0Jx10Ts5Tnk7jMLr1TheNlnbP32s+IzMFMrhFw3Xk6mI72yrfpA
4LcdHKLaigRcRHAfrshQuAJhj4ecrwEI0hrkdxFIS3ZJihyjYYHho0/ym0tz
/lZJyWKKga3Zv8ukK/XvcOO+W+8Yft/K7nTUB9H2O7VvIqWd8qnaaGZvyvv9
mwrRskGQ/vwX89aVHJphxxcaIcjQNowpRGe9QgHuLqLtv+mJQekQgdJ1Vdoo
uTA/bfEdRIfFO/BfR/2SUnfNNLvQh29rmHpXZ5MrVhtTbQakBzX+7vCfZ3Yn
q8v+T4STmyQIzOfwklZkn7A3Z/MGNMHXhtAnnnPofuDOFrs8mzd0/SK/bI/j
use1vsPH6qNiAjQUrNpy0dtO6F1JqnZ4WLoNv6H6h1/aTVP3CW0ZZSfHfYxd
olzhFYEb54mSF5MH5xNEwrtCDhs9d1oOTGWblULyiIkrft5CsBOuzYHDoo9+
57iebNPbiP4ZfB+zZEh6YN5JVcWKth9ZujwZS3QbLHCyHZ//Fz7WAa/hTvEo
u32nmx7tNnGmjYJk5ssMktMQuci/DQ0i+cS9/KJBbCoAoP2sLUeky03WvTav
7dngN/WB08Il6Drb/6ozD/xPMhgh7/AqB7C0Uql8mbAXIRHpXS2aQ3k8L3TU
nV6fVb1Qia8GR2ZaWE/Zz8oldLwnxcIu+yQFHxajisMnF1TEWWtczOM+rgIX
t2Yfz1z31DMqa/Ze8GeD43E8+yBhBT8WQkP11nWTDAjIrBmVIrRUJI1SxSI+
9aW13dHjl52hwM2VseYnMYh9IuMXMU7pp2S0aY+RovU2/VFmxfGpIgOIQpEU
GBC8h0xEL9psJVPuEHP70snDA/IkExxPC5Bcs+m4YKrbYhSboOrOFNGorVBx
PqLQinzWcbB/6Aiui/2EMvvLb9fVXOxIb9a4PK70dEpUv7WewN711TsM3Don
PMg03jyBqjJNxy0FrpzVTjTiWxCSwfZpBoPpEFf/slFVS2+KGT00f3lBMLEo
6qpCdDg3OZvISu4YtEmSX7Z/4DugcIugnac3styhB8DIq6pPA8wwp9yghBDa
esRUrim7KJV8wxkpfd2fZKUZw3xhCOM4Ws82mwgPhs46KGpq+Qu+J99IJPzp
v45JYiZOMR5nrGOdXHJvcX532L0Mw7gYKQvn7T5FV5ov28NAZ0CiXah7jFEm
cyDChthBWz8fK/COnJFQqOFF6Cm/AMXue8VSrThIrg1EEB/dTfjZoywgC2/U
EivqDsRbBwxGD4ByrA4ZIr6GYKCJAFoby5pKzv624fn1VV0IEdoZIUkPsRV3
mFtIXC+F9z2tfeT1rA/fnOeOlXtDx2e1xIWTh2mjxjJHc8AiKTXyNCvANutB
xjOaXdQR9czx4j8GuNUdFew7qYFW10Apl3joGBanRhU833+7DM168noWZkUA
oYVvGGyeOoPLTSKTVtQGfcOxaLydY4rW2K6GC8/kf25PB/WkLuUHuFpG57ez
WKdEv6C+ny46VbG9PEc8ZZvhhaD9y5OAbdRt0E+eKqeymnD39h/MBN/I9FPE
1hZpyy1GIYfn9/jBvjfFtAOh0VmujN2Oh+M5d6+qahmi0xTlweP9DNnhPDfK
JZEeaVxrGYL3J4uNuPyZFjnvurh9TzoBlYrsJXXG76uNatbN+mA3joxcwAy6
O36HC0htnPOg2yjpAkMD68UZOXPlom/Xx3JIUaRBussmTa3SJ1JifZzwesd6
Kr81xv5OCJt2ynatRvS/DJIjcmwlCZppV6htn1NucpnHudqDwlUs5pEI83xd
64ZsdLgRDdrfo6UD3jSnIHnhq8Xqa/+GXf3AHVplmJrJGyzKO5bpv5yl9ztU
9tpuUIRT4z24uPu8P5LIFa7OSY/54ECT6or/PymCo1dbuE7MNDxwhb0p7x4u
fSrA9McQNFjzbzmzAFP9jP8jQmYe6IzWBup9PgsYqPXgFtIDns7otWt02Srl
zIITKPLUQf1hDwS7XRXiDgZHXORBFRcWBk/ZXRc6sJWiRml81udtnrsSKoLn
r8OIWVP5PzxOCQ8jup8r0cKIRbzuVFrQ+rx0IBPOZ/2hy0IES0k+teXuMU4K
x5wIex27zoKh4S+bI49lDaPQwyyUvnyHbZSpYtXQY8Jt9MrhBVk/BYLitQZW
HS/iRu0rpfpL7FRJ+x8c4kja7NlC6bsT9iVIh5qC17mJV8+S0YvnP/5kPuQe
uvAI9GejgY0YDYndagGB8+pns9GIx0qo4SR65px9YUF+5RYXE6llOUyzu8I/
AtA/43UFkiEubKOiu/ekP2CQbmwNGl5HBl++H4IxUMjrlbONkZUXj+81TbkN
DUk4KhJhds/rOJHOTfpT5CPU4Ek4hhH+oFyotL1GvgYgiUBcyntXO8Y6Xtzc
QoY9qnXuP/A+lAuZ8stv9aBSG/1O79wAX15uHyQsztl/SdIpaWRLEBq+9Z47
s4AoTKqW7vDbQS7mrMHtWqh6o0EI4pgxst45xQBV7T0MfZaJOo9uFViy1c+s
WZKjbQpkqMEx5gZxHdCWWHjpC2J+mkR9XKTt1KU2Hj4GPPoannNsIjKCj8jV
FYDry6C7yBN8RRnLqhopC3J5r2z6zKtwMRuCCUW6B3f7pL4bFirO6XlA0+QF
jToxzqARBQthM+wrac198oFE8ZhUB2W60p4eWtkctFcPk9CDNMpl8c8iZDcp
5tncAnjwwLREfY19stbuZbXF4eoJ/Nl9W8HPz4S1SrNsaFdQ8UGOwntwSp/n
GmMfWc1kdFq08RMyyHnWYeqKYuLAIsRcx1H0TG6XsO47K4cbKG0auhW7VA9w
DEz5cKuBFnqm2zHDOCC3gYt15GFGKZWi8hc8qmJ8dgNF8NzIpsANo00o2ciJ
YG+bT5uW8V7UgmLLpjz0KXAokXS+sKwcQywLbJtJzUlU2fvvlT57LvzloalV
+QpBCw104QIHKW4708j2Rl7iUNl4q0N1dj8HHH8VpU/kLXc8aTs+WQFhBb6Q
3/8zIoKmPjcYfivgeV/ugHWiBAifeRrGi78nhVxU8ggA3sq0OjLX6c6WXAdF
0pWXgBxXGIzYPnA9cIdwILqtqPs+Rwz9WVX3j8hBt84G2SHwhXSDMCw+HhVE
2eMx0t4r/EMrPY+LouWB78Pf2a1EZTlKQVX+Zh7/szMpZMp6287FUskljqsV
qAesphfMQmCfopTR9UQgkUWPqjUGqyq8Tx7dCfbj9WwVORoyaSJHX/pBbIxI
0PSTF9Qy0SiuC37YR1U/nvMFMU94BFV2i+zPF9uphbG4Rkw3h0CoYtbR/uiV
g9KAxUwQg3O2KmN3SzXQWHx37EAAE0/vMJPg/arHfhZUywtAH1BX8joqJVZT
RF0WULZ8VFTf7ZfXtdjMGFUvCc1xmE51XFLz0/izeQcgnv3aTFM6D02nY2QS
p3caKv8sLd/27oobFQtZAYUf5HTFJHvkut/2CntfYb4GjN94jGn0f8ogjp5/
MANVpKiyGWK08TbkONUY2U58mKsnzL+5V1H7mcVKuaGSyAG/XjO52w+iPW5t
GMtSNqMPRleHVkHWt28YEzRt/piBSoTpoqRfO4NbLd49WskT42zbkD25sToo
WjI9T5o9Xu4FnCUE9uWFAD3ZfIMoLu9GfMd5tc+2tuxbgGQPS0Hh7BtY7OPE
LWzNWByEeMxKftpj68Q5Im989TjDIR8caKb+USiX0UNQ1UKyScu4Vf0qkJb2
mbdvivhLUjQun/J31XIaZQsHN0OSBSX3BosEY/Js2mRrQJ861GArUmGezz7K
hFnvVUM4K6tcclLd4DYSe+A/xot7/kxyFCNB1sdVpPwsNHggqsaU5tYcgg+E
5FSO4OYEdLR26az5MmZJT6PdawCPs+/0UPHywRo4PX2NKG2RyDbraSVoWJmT
rnXpkDSi5+oVGhhLEvZ3NWboQuskC+OqlQkxkXSe0+sLB5pfVbdVdR8Fj4et
iN2nAH+hXzYLMa6t1RaSZhmWMKXXYmzzQn05wFZ5YJSUdFfxadf2lXVwRwcf
yFsCQMBX5tOFfP4nGGWIaOj/+dSL/y1Yb0lQ1v4cMaa+qtzLehuJ+65ExgYR
bQZRZzaVMgKfUr6ck0pJlGsX63pu9TEO/myvmlxy5IrIvVcxILW9zhxhXzmF
y8nT26ukXqDf6Z7O0WYlfbhQzskojRAFAQB0srmNxARfLNAG8fR1GZ+R3w9n
19vwA63dnjhxmchYBY3NIt++RH8ArAw4GX1yqjdZJuT2gNPMCJDEmvDIqQec
CmuiUGG7PFye/II37+/eO1CV3JiM+HV9wTXRCabvwSZbTQpinwmpXocwj9lq
Zn7WcrT78fOZLrmHThY/yoOdFj1USLZNzR2aYKhFqkOTM83EE3gvcURwK/fx
t3p2la+Sxs85IEBmgPEjNI9owYD3hz1Kt1TsOogNj20aG8TdpwRSSQDyOXMN
/XKVJ03drYNQdJFaaXsV3GB/KxyFWg68qY7NYb5PMvmCtzgmYsY346kEicHW
2zE0EtcwelK2v9Q+P8aWQKSO6Z3TSGMPcaTAjwmFTyFJa+rnKHjy3WKUFE35
AeP+Sr++bJv5dU8EJmF4XmrcYvtR4Ruq1geoRKp9lOiv56BNu84fV6f2KqcW
jpfEYo3NuBcmLGvG7OGAl2EGXb/TfgbmVxX2BvDALFS6dl4PLh6x82Haeart
Oxsq+1XLJtEUi9SizQDhb96i1IWcaJk8jSEpoNwoJ5ZD+liBxl3UWPLdhyR2
s8SLJWd/9ApA60/HTrtn7u1B2e+NdsmgMbLZJVJpPawjWJ2EYhgHdr/hyUQA
aMcidISurTqVkWrVu+1XCIBrQO9Znals8enXOiNoFC2jQro5hSrzxBDsTBYb
CMkGTqjwEvZARThFAEdLdaRQo46pmBzTooYnGGl1rD4T7+m/AGk3fIqt/rCO
yFIbNRnWThf8Ld1JN0rfNx+kMmF4VLdubvt1COAe+hFnJeWXpZNEVmxccuUI
QWiEs/BzGDqKRdWqDUB/YIWwv54LXK19AlvGU1i6XZUUD1otFClZpr3kau2r
srlOoOmdp42Lz6ESa/YgWNlN6J+oTy0wkvXro+UwvWI6J3m5P9z2YUTfgVH0
Zz3pf3Ni/XDzJSV+WvUC2yI46e2QkNUo/oTyBUpqjT1lOlxVMFCylko5rS0h
jyx38B2KZ5pb4NyZZDvx5qbZhiSSidM+J3YQfFVU9W2EVDGFeI0XIiZ9BheS
q5fV/h6rtcayeq/KOFb8z38pRFqvJbV5DDqsCsVusYzXLZLaXRAfiu/pEY3j
2g2nuLjRwEJ/jwIFzruwvsuWA890zBwq7hKsbVKT2grbXAJQj+wRKMQvXEmO
5aKZHxGjpQAM7pDnfT3qc5+i7dYL/f79lCL7yOkxDXF9DihA7GewxzY1/agf
Ahlvs5rD6PbQHIyoP6IOSrZCuqCKpvYhgd10da1mXJ1joI+bF/2oYw0GfO0z
Z9n1HZCnDrzrtr37/hySWg6IVv5sC5yqxaGa5kzdT1jTG7JtOY8ZuCRovntv
s+ABQd5mVSUYPjWzzDdXWmfuGo427ZBhNqcJrexTgBARKaB1uZP7IBnWqjh9
5PNTiM7ii5t0waADfaQ9t5LoE5mzUGEUjy38n2nXbOyGXA//wQlvFpvTOd+B
AmV4BTphnktQIBMtVo0csJdcOSHLWzMSqzenWi0uJAYLatjLK+pv34dIYvGn
nKQz212Lu6SlP8ew6S9f3+pp6Ebj0Yj4B2fecaujoPS+spRaViIs8ItgYnWA
KfHtdybV+A4v/KSN00EiY9CWy4ZZmeCP2sSWNw+EArBktx86tPit79vS3YOO
Av3a/makCE1eUFnfbyCNRsUDLR4wbVHVBqJ6w8zOQrEzSa1Y3P8WZe2ywO7q
ZE+9GEtw54IrkvrtwBffOxAnRvX8XBdjtW+U3zAQYMyHW9fo3eI4FqpPkyhn
D5duVoVgzC28dbJVH+65O6sF5uLptLv7vvaFzS/cHP/qEAPsS8TzGra44qiH
evO43pYG8YNpHrZvDkFWqbxWxZUZNGYwMfQXylWXEGGOU5/m438Y6UmvOzD/
L1ON7YuPfbJWC8R6Py0t9sjbxUxZBqqGUG3X9GByr9VqbN9Ix2ibC/6lB644
esBy0A9jZpO+qC6eSAnhEMephJe4EjcLav6SqQD9bTirpSudL+tcvNCqX2hT
IS7ZmkwL/BJNzVg9RAqGegxpVC/GVbPyUtE9VT36KL9cgBfj/7iaYveUCiA4
Y5PIhgzyB9VYh6HLPLaWTX+4XliwyRFRxKHRh/4gpzd16x3V/HSdt3E4aUnh
byMt2ZlMA19bAKQ9YeqNenSZLxuXPIlk4Wh6iOIKLEqy9+c5t2W8MvWa412k
7hUCyyXiT1mFmMMfYZlCrR+e/KB6O0YZhqVOoXcUKScdUZexakID0kENBKcF
4ASrYcqKJ5lw5EpBfSH2O31T3IgvCwNEFyEutbyn1dhrrID2DMYnpWODRhin
91lv1T97ovO0iamEXfHwv2OAkb0beeV1wZxuK4bURUyWqD/cnRVgNepgIxEu
H5qQ4VlseoF6L07GI1jwjBkoNpmvyOLBSVb6WwQrZ2DD70GtYVjZwzz8PZet
7xs93cTkH5oPZkoJu1vSS9EvIFY2N3bBAcxgkSoJqxxW+R0BONnHjYpwK9CI
ylRULpBq0kyXFun42AQzA8/X043WVo9NPSn6D+hdeeDkVALkfRAsH3Beb8vx
49mKD2v9AZKKkDOp/C7K9pN2WT6kTIWYocW/vvKOenmeNKfYNbNYkSsfpoRL
jAVDndC8Zj3gaZq5HwAMhvTHXhYBV6vUcVyUztA6Bcn4M2xxupPEFec4MGU7
YLfE1MPuVmDtc82VFFqVlSPW/Jag/ce3clyoAnIdFGevSesqWzFsn5C3FgtE
HKSJeMpdUo1RXQjXdxlX2SytUKiJCbpsBQVyuGPIMCQl5RfVdXwWO2TgK2pB
e4Xn0VAOABVAnavsnczEpWJ0Es2Xldn8r9ewj9r4yXTpoLSKtPcYywWU8ZTX
5oVTRoCYJZmuqvUNPVgZxqtxxicfz/t6ZY1OblAKkrX1OOxalIi9ehGq+Ozr
MzBXwa6gCoL4hN/hRHDhRNd3be/BIbx1Tz6PamgtJE+58EkI1zs89ZTuCCr7
AOG0Zn5pIhWGkiKIITE5Y5CLF3n8OEbaWtMlWlqTP1zt/+YN+rJSiYrJTOyS
H5Mmtt4ksd1j/G7ZZxWXU2QzSekVmwLUS1u84CAr8onYB09LhhGS3G9eQ/1M
EsrfpwYsviIGM2kuORqgevV49O77Ki3lGH+4/lTp7Bc/KlkbzNXLzed3wZOW
JRTdfefY2ZJtdWnHge0DA3Rldyb/wn8/BHVJAPJTPOnsPrEhBkEjfDhEGZPC
jdzm53lW5GN2a00IV17fRd7aA4ocUJcNylfi/4stGJWjHkYoOlS3paGBWXNH
+SndiXiSalmuwkQKppZXL21jyuMp4eUjwPp1KNmvHgVdKS/51gkWAe6QZv/n
6J4VZNV6xd1V0WqjjWZSE77nWa7DyDidyWqJI2rZS1s+7mNpPIsD9gRSdx12
NMxQUvXtxzT4yP2bsexYGWfZi+XOijizYA642RXmVpQvKLYQgBnDAyN+kaXo
5st2FfmAn0ABWw88pNhr2GQlc8ZEnuJ67w4ca0hdW5vPp5VJhY5RUQaoDxv/
RQBBqysqqQBwfc0HHr7ESfgA9VqX06FTqAeM855CXbbGyOfcaAK3AdSmnRiJ
ociCnl0EyjdjhTfxlag7XeAXNCVULDbZrTvVOR5urp1D17/d8NCBfkTeZ5Sd
Un0IO3B+wnCBa4iLt0OoEZ7v3/GAcwGSP9r2Gh1gAxcO+yi8u1kHK93mcyTQ
Us6duisH9AG/I3Pd8he4Mj+ALnMrJH9gRlSaVA3nnvAPjWFN/gclz3MmRyc5
DlsW/XJEeXVQS94UQR27tv5DHxK3/m6/u8JGXsxYcdL5Y2+SuTcv/6Uy0yyf
v8Zao4ZoSrvedyZbg3Ub8P78h2sps95qM+VvFfxethOW4E1ueILaywmTI3e9
B0mCwpZxbQ/kaj5Yms2L2VmP5gh9Bj4iKejCCBH3Jh1Yo75B8GXVgCNA1XSx
Qu/WBqxFDWPPgoY6JzICHZ0zEeQTndDEpr0oyRt+ngcXrZbKeT9b1gxjTYE1
urwkXBAHd4khQE6z9TZeiIVGnlpLuwmFzjtRXzZjUUfBUtdEqY56NfyMDGcU
AKQCd+L9g3Hwk9i6m9byR1gpC0WUORhgfMzKpPjPPa93Z9JqEqekrfwDDLMP
7nEUa1kN7dHuCOAN9nsoNcYV8nvVqU+ZThVFSLQDb17iqqSD8uXav7EMa/RJ
tUIaRYvQVovjH4/XHsCzx0BPTzpswssnIecA8gAtAcNnYgdn8kl8zSAiGebJ
4xHUWzhYt8E5nI7wMieTf4Fs/tJCEND6j7JYioxoK/fMMXeiYTgZqGAg6zWE
ZN0O4LGt3bu5nFoKWxq/lUSr4VeN+vGM5EbZsTkhZAYW4jp+kNT961Y60Rq+
mVFM14P5/46WaR6ykclBaqlhfbLi1n2tYgIspitrSVnkEro4TF//OyX0wx6v
lww0GxC4vJdD/dtdgJR/XP5oFhkfL2jjDM2gZey1ReadkmSkG/rJlEWxIoYz
wWPA7mOP6xyo6jzRhDHVgmTc9qbFZVIIlnOVxXVAHn0o+fW+XrW+AmQYsa6i
QFuT6MLgMmyJL0Nu/nC7fhYQyk1wUsSRtZP38Fn4KhYNIzBO3bJXlfznedZ9
Xm+P9u/PkgupwCRyUVUuA2ZkDgRs98G1Z11k5GyIsWayCdoEKiQT01NIkt3w
Lfh/QJQkSsbedl+0LlC2hSKczGnqRZVE5Lw1y7WpTNbUbP7V4aVxCuGDrwnT
9OxtFsq7goJDYHsvTqfVv5UPTMyzq4ELAS8UP1MHJ3ltRdeatF+LENzQACrd
eXxxilG9Jk9TT0a/fu2URiURSn8ks/RbcxVWe748NhSnXlNRLatJUoRKGJN6
SBxHbZ8EZzMQLNpFlW52n7zTKknZapG74KyUQ0dsYLebEzq7chF79YoPom4y
l1mGQ/FCAPUX2mDWOmoMWe/SzdW18U43BMBl+6E0IZKvgLkyc8Ok22ovFfH4
j8NQzrTcXzZspiD2nW0cExvJUr4qwpaE3bwOi1Ogu0J1QqpeRyrgP5v2JGPZ
fd735dOvuXxPE1DwgXgiTQqCo/3mJ+zP47ECQSsCZFYrzSE6c/KuxPDokHcQ
Q09gJ9yut9fTj7Us1nHhokfszhU4RzhvsCK0vrrv6rH2diwPga+kfhudMCyK
UcMv4ovNAZ9HRB4ACXdQ2wMa2dSimwKg8stkLyZ3h90U4JCfWMsFg5PP5Uyg
tVvvU7Ylyq71hYAELWBznkIli733RbjgFeN4abq1LjlzADuiAKZveMjib5Ia
3IfmyHB8AP5k5E2unErviWSPMiHtGZIWvLr9zqxMiatb/odyLnIyitJ6ekkl
HxK2PPgaBcLzuzKjAak/kCjoCJ32n8wYr1c81jArjufP5gxz0jwOTmv/p+fb
37lj7p0F9rs/lIT4A+zjiUEBSH9/v+myPbhw3OX627TfvIf2gckgadd74bL8
Cn3WwoxtP9/wKhSPbcgMx1t8EUN1dmQSQjYDPvWKC2hCsX1c2ZboNj4/CAad
zVP/bz2gElS/dX63OpSG1U5bjV6VXQykXN4QoNdqI69Syy8q9uRiCzr0yWIQ
eUaU86tKPvGDXO7soWVmkwUOPSlc+T5WfxW1Hgs6ABg5OlmyTqWcr83179b+
onSLKqAEX3EkGVIjOWApPkaW3zx4L+0BW+v2DablIXlYfrx9ED5eVsI3YOdo
sEl3vQK8EZx5KPohXzccyyhsZwXcNmfYuD63Oc9VCBKBpZ5eN9O9TIN5lT8I
5Be063fqZGzX/qgYK79EdQBQOr946amVzCftx09brkW5z84K8GrZ9+81Exd3
laEpCxi8CocKeJRtiZp8Gbh9bBUtWkKhZZAhZPzZh8OxjjTbmzvcbvupszun
twiqtH+6XiN6frxrDbI23togzZLdax8FTMOgNXVSD+F5/zuUGMSDm3sBwkNJ
z0NBc1jsCEg4pC/Mpqq/dWxZqtCkNiZoaK/eCSSgjqy1DgjRvmWrTZVq+bby
72ULCZVk4unC+aMazHx05Y3Gvt7obcqgucIyG4lt2CYQx78tyDnfVuYGmqbH
UdtmgEnwPxby42jCy6V+VqTE7i+4Vij/8GLGa/XsmGbYG8jr/Yws8nzJqrzH
mUNpaOV3HJi4iYqenoIhvhZf+ef5UekrrEXdbXtUrZUN0jEYN5hBHk/z5lyX
TKKE/5jBJN5j7IP8fple0jWnwzPVV9xz0KFQfB1EagrGCZPoqfDAbXlbSHWY
cP3yVx0wj+ZQ2DHwhTAlQ0UuK4S4SeuMZLEl+oFWvfLW69it2VwWTjNWWO2q
bJW+w0imm7EvUlQjn+Q+ndq+v85/PXWcXzIC6DTImyEmE297MqKxkA5Aq9C4
yUELFX4/dkyNn7ScVohQu7hfIe0Re9+/Bp+qTL7gozv1mQ0frOhW9p9+x4qK
rrT4NQPpasLcN75pOBfH5VOBLwsMwT2Yi4JeblO++LUwzwdCxWLe8U4o8xXE
0uVwOecCyDkOt5bcTfXjUKGSyNAlS6Xahfm6GpDezuL97423aJjXIZDB/4TM
5WajPmvYsoJ2JpHYUmMYgQX9oIs4ozlVGND4uh3jmSAc6YxBhlSdmT6UUHhk
4gc0GSguPgwIquKDR+s8HqW5yFbH/hHVSzitzoWEXM58B0xgQdxtBPFAmqhJ
RT1hUT3u8ZCe9Yw/d3fepfgitZ1l4U4/f9/EW+cLSHgYlUNaXcjdrCSADhFC
hOkIVvNboXntz1wzhfG94dTDw6FwHIdpIDbVoVzZ/lhhHU+8s2Me1ZrCtJrS
G7/XV1DgL1XxWmTRUY43VejB6/3XBwZ+Qe6OL45/oTO5i/RTyEu5N38NTm/6
rqZbLl88vN1SdCttWfSj+Ns8DldKkYEA6I2yW+KRlZdjiLW9eXJIN1f29O5T
FGwQLGg/cmacEhZnPUmyx5E0/eRzzjuDR9271rcjrEcxIC0aILyPP5q4Jp9D
N+EJEYZFYCKLyBSKrTk5O4B0I0/RPy7gRdGSj3GZrehlwMktgB4Jg+zTKKsp
Qc+Fu/wcJTyF1+HhbK3/FgHPt8j0r2HfiwwMLYSQ1rdCkdq/nCldg2saRI+4
tziCQ7HAJjouS2ytNBr53cNRUic2bQQ+caDt7M0NZRpC6X1nFaigvNDYOQhS
NYwRF2PsB1i7OMhJlf7RWMyPmtuHe/rK5YIWhK7XGVxYfLqAN3Ir1V15MZGx
2C/RT60Ir9Kso6jgOuTW92H+Wie2BOOW3PKUGmw7mJBPiksiwYxCNAGRqTn5
glfltTk/O9WZmBzN8bqjX3clvy16j+1BZ3xCqDavHXQBNL/lVAnneefixYlU
x+JD/sQCzOEg3Jgs0OzWkdDx5bNNVqpjaMLYNHOVGcEB937Eg9xKCDJ2vAfE
Omd16q7CkNPn1QA9P/ucOUANyNtokoyE0auEFb2Nb7C26IVPw0Fp+tjQVQ1v
+cxioXHdNEN2P+TJutQw6IT/vC4AcJX1pBfVCvlTsh8jKBLFT3HBuiEIWq1Z
FQPDC6yq+X/FcAqQwRrE+VE3rbOS5pTef1nQyUrn6zFqSDHnIoASF3UVg0xs
4griNBuPQYPaEzvNixcv71ISBQqxcxpD5LBp/PgcusjklDFE0kHmDMamytvD
ImLz0UF8WLorbxs6Rsl2e2aoayDEyigLJIZ/tyg2nswcpBbku0Vna5OJkys7
acBwjneGk9sEmTVp2NH3qEKe7CDPSmGRjTLCffzLCuMTFIyLjJUMUhUReAEK
1MNdR/haGTD3zZNcqdNPrjYfve3AugPCm0YLgRMxQfeCsTFI4ewm1UtsUcb2
Wu+YSoipUUsy5oL50+7wycy7xTLQZkJBlTBJDe7j/6xZCTXJiZXvEXh7m5Mp
H14VXDBmGcu7NjAE3jpDWaCcxWRdblzdPOBS2T6rahY6wV2M5duwK6uj6bF4
kEbzQGl/m5DrOyUjdYsiEBd4XRPBQvcoWRKTCT4XvEsLiDiUT1MpA443txaT
s2eLS5P3HXkTIyZ16xKbtlszhSqLeN7UhRjX5iuPlIS2zHXv7sivafj684qn
FbMcbVjk/Hu6aZ0wugx1aE7TSxvGgV2VldasmEBfgDyXPXhaXOssuSv8R25/
eY4N2ui31TpVtsi8G3J3lGaxIeVU1K8MW0ZbeJASsimUFNO4CxAAZBWMQ8+F
UW0otZ/L2GkOR21beNL8+TXVWIjmJpRl7U2j3zkZtZMgMKLTn7VFUH/wxEyH
gW1k8qtLrBsiLVUrBKerPY68irR99oTBnHepeamkxqTwKA+vG+CtzuN0GgtQ
bBWgaFTJiZHbWaCRJvvzvSa/8SH4RkbbHhu4AXmMY2oua5PSNGZ/PJRmvnCu
z6j7j75t4xfJlgTaOLoJUyr9jnNUiQPav0lsI6GX/TlP85sOeiOCVPqUKAwK
c2BJg51UlDrXev2q56Ht3f8pSZ3oBr43y9IzIw2JE2OONT6GuPppBaIu3MHd
xcRbpqJF3lFrnkaXVrXHP0psGEsyhZEUc5QzxrJ1423DHzxcRvceXMETJKaN
y1YVlJ3mY5GtekmOT7N95qgwsUEkMJiaLT+3u7KoQji46ZbZD6Jv18AAsOIN
dcZ4pJkw07GuppLVj85FF5ovYQENYrSDBc5SC807lavo3eToDyp7LduhMDpp
qksQqLaCY7gZc4zp+SUe2QtJkzlFZUHyunc1qet7ko7N5RRWGtCVhdXPLeC4
Q8bacMIYreCk463jh/b3J0JTdbzYAxw39AaVTS5aBMyUVxvI62DqjDtMvtqU
7YwTraQJSanDaGxkz+kCNw1IR/ksFV3//qaYEbE1/pWhqPYf5j2pi9+wMRU0
1ok3Phg6pphDiS0Sum/NXQ/UAHAsPxumPejqLh/AUfxz5Mmer7RZxttHjH3t
RT/uVY6Nwyo+hC3OvV+aMsvD3ZaCTbEDtJ7zTYNsXkY5JrZHHl+jGIbWdH1w
5+Kt0efw8ZHqibO0DABowEEC/WCbbkZ8tjDXWT8Xtf//tv5wjYAE5niHxD+7
4az9886fq0HHxWfMZ1gXJiq8nt7oj/029MLlGjwFMl16gmNowFz86AmOIjKl
OY9FXRPFjMtLiYYk1ue9retNY80Mpc0LACLJdZGoTjEHadsU3/gmQmfH4xE9
+uvPmF1lApdmPtcIHxouOO9X3fCAbKgkB05dSp+gJ5T6fNnSpnJrPAgGZgyj
Tl+KNP8SF0+/aSmScVVIjzN3fl7+kirU9yGcVubXnmZNhfURQStlEtOJzAsr
V2eLEzKKfc8q305q8EZBczDytjT+DKj/jzk4bYHGd8JK0VvpGUcwPDYhK6Wj
zuTVKv/4uIyv+sE9fvwkSt3jhD5o8ERVzxHCP9V5kOL8RGTbbQ1BUOG/Vu5/
k6vpiDT3cvljlSNnsmt5attwl9mlcNxvC53k1q/rtQkXI3etY5c0iU3Aidjk
rgM5VMlT990MwncgsjBZt9k5QExRv71fBg7iVDUdu6+5iAL/DmpOUPivcBiX
xTdCP1H5QDdwdlx3DaPfBfvxaDW4SELSCUKSUIUuieVG61WGS0ChLIOKDWeb
t8t6DV9SO5tnTFqzUlTsbse8fZZDkV4YybAjnW7MiW2nhkJZPA/58tWsHaXJ
H2tUcQnbiVZFPdjaRrckjQa8ZO2U3qKNjh6fndRbudd7jsS0HzUxNYwvCXD8
zUWWJZIUdO1mHlc91Rj+ZN6Xt4mrkJ/5M6bx3k67LB9UJstK9t+LxwqLbhdy
h9gaqDotQY21DXVSUIXc1aPzXcZ+uX1SvbH77t2PsXDsAs+lk27aV3hDLZ+b
2MTKoSEFKFa+UDGVrvMgAqMDIVCiE7X505QQEuptld36lvE0c18rq04YjebV
+AfXcOjKSCcqAMcdxo6luAHEbVrZuF6NRMg8NdnsiZCOY6tNBn3fROrzouEX
KoGXC2kZUmI1UFNSswBhoblFCY32kvG2eb4HkoCPTnefuXan9l0fKCzYgN1P
l0ExZZH8/9D5ehTj6eX9zvNgiZ4w7HkKSG8dT0VPHl+xFqfPnqL61iED83rY
u5cCnV3U/BKnKKgLYk/z7qbaDw6IGaX2VZS/ej8xX91sQYba0Dj8vfu8N9hO
w+GlsMcJeWkngZz4ynlM+LEUUXm9BL9hbYTImVyq6S949TzlammKpga0n8JL
ooc0daR4GbET5lcEddlUyOK4HNglBC/vivX3e0bYQuKHQyjiAgLlS657A8of
egvetAKithsxcR75SNWkHUkEqbF47nBcNzzYD6wCcIlF2xorNm2caBvQ+kWb
/6Rl98jJm4ABjZUUKE6bpMKaWHQuvN67xUUfxTH2SQmtdn3kEhMW/VPH3zLF
3LWWq/qX6uhMZO9lEb7rxazhzugSzbSd304o8K8sf+obRKPlLESx12p/aJAb
ltcKf36fqGD7PRmnQxgZTtdLR5CS+VG5LPq5omyo+A2O/jQKCIIondpT6K9o
gIhBzCBGYdrD7bdt/ItsXCV+d+dGRMQ5W3ZE4XaXAsutDjk/rsWuCW0bAD5H
iaSeHERP+mbKT/yLBpdqBuBRryXfmNnW7bSG397kId4pRvhPG2nULENI1dTk
RgcbEo0B9hpcAXAI7prqgbhNnW0lMRpiJbzM2+q60kr1itYjlBc8/v5m28Ev
w2J7KGXlmPfU8rXKYbR50nO1zpwiflmwkSPSyO1Z217RnLT+/W8BNRAh//5a
UldoJpvkHIboZ/UJ3hlv6zF5XUibxjxrDJGZFCMdEe5/w1knysNcE9tIeUFR
H5l/WnunK08FHlAfxiHvLSDtkX/UZZpJp11BC271zGJMsLedscDgw0SeXF8f
oCil1Oz+KVlMptNF0gnNiM88elzSVlQ07NtvY4gwOz2+bzzK4Qwky9J3ANAF
4diZOq4vYr4VkLZQQmcr30BohLPzWmpgNNwxcsR4FKZTAfZK3BORORTP/mVN
zujbsHSlbvokkTq3BKqXy0/6CPHL7BPw4ghATrpgKVifT/tME+7cnNaJT0Hg
tcM/93d1tH6y0gctHrDwNqe7o7O29KNmB+vCzPiYKZYRdGrUwdVQl31UF6fc
xjsZ7idfSchRlF5XxSBO7h/sZ5CrjTXmCiKUwoN3lZo/Kx/12XoHoVIfGW0o
yu9GKLyqZPyoP/UjBlYYX1//tFT4Z6mu5Jy4q0dFBijovtHKD423MNvwSqA7
KbBNMUihbqOZPmle6WVijKCOJSp1z0qZ8ISztjoVJzndaKpJ1gpnFlfsv5CQ
fDUtz5BeZOiuxFTdz04SsdMNcb/wVqXQAeoHbrAI+l2Bne0eMcm3ri56CjZ8
uwjEUW9eTe1P3VSAuTy7bBcm6scoDLLw/+j5JiatnlZh0bllf75g/EkV+8x9
TlTqqAtZ/2OJZB99KLOsfmpQsomBf9ilF2Rrcew6lXkJYGdPNY/o8PKY5G0O
eLdIf4+zcZiYgnPpx0dcH5qgfL0iPhhnKSsaIFPFh+XEwyVEJTiYBHzL4Ejw
+VV5W2VIKvpcsdQs7MnjeDX7uuwsjgt5Gf0fk0aTHOCWidLU78C7bXbY61lX
CAud0/9cSXWCpYNiW+9CONra+Ym2IUDBW8vYD55xX03RmbtJIb4hSH8LtjlP
DdGzsUTrup7wQSBN+apfvb0uhJr0VyyljaRfyjv2VD/oYk4sLUbHmP6B+2d7
V6smzZTuRIX0ysb2wNqzoDWXFiLOIY4jyi/SNDmC+IJ7hsTLU/x6UdoBAOoQ
kyRBm2KTF4qLZAZxO87sLqSv1McvBLLNFAbSB5SaTyhN5f1GupP/f7dQD/lB
1h22lpzQJPQxekkM7biCV4RLJXQmvmCFi2YM0zAVAN2YSxVVh8a8wk7Wib1J
QQvDU5vfcnOB/P6pSbgRCIisL47IXuh5cxggeWycVnVUhAprwZZirQXoFg54
myVpaj6fYMGQl5njUNc4Mmls6xwCqogaV6UzntgkKqt/p4aU/hDUtgMC/3DK
qA6S/hx7zZ9gFUvVwJp3zzjcRUS75ZIM/t+clG9crcAzGdVpFrj4PPz2wY5T
0RHIjgQeVsZNndQIbZKUCKryOORo9M52zYZ5laCVI/ohCRaNjYRqGYqG5rJ3
MBmys+0RKns+kiom1HTZf4NjhVQ2QPknDenArZddyCQX3RhfzMaR/+0LtqVH
/FRD1200xxoJFYjvjoXu4HC300zbGlGD3C3nke56CZzUP81M28FYMdP6sdSo
WAT/yUAyWLdwz1nxrXN64c9t2FHqtN9xkSmNT+Y4eT+vDUhLxcQTjrsw126S
GimKhhpxVoQCegss99FgsuVzeYcCrB690RIpzk/h3V/5E2oo0Z2cuZCeUn+K
OuaqP4iGRDakPznS5L36BYuV2cwQ2CkxL3+Mj/eE0kizucw69pjEAHjQArti
tcHw11d+b4t1YWkTHeckKFDGex98/7hh9+GiJdlhK0eXFtqv5BkwRIHnvvAI
YSycDA/ybcRRKEqtHnZ56SCrI6XHp9eKTXlrqsSFmo2/7m/KY6NChL9sN5u2
2GW6sILQc/wWc0GC03Bb3AKuf4p6RYhypNtkjBgsy4tcBWn9yYD33X/GDsIC
/hBIHKhMHw8MIxBXH45Dri5VMxMv7A3FgRnu+imLvY/h9S1HYucV0A7mO4nT
X34XTNOIA2RROdTMnCIQd2kKizh1hkpXCBIgQklwWzwLuclvvibPAfsFr+jG
vjWcSkdZRzNu7c11LBN3dMH9mKW5raVjJ0A3GkbkVYA0f+NoJAN0Uukgc64r
oDZg/etcX3n3qPBWT4ZVqBvPKA8ew/VvXQ7S6SFj1P44eboYvXqacyG8sLYp
C7Zf4gsJq6GKIZ+5pWX913sQ80THQtWDc6gjy8i0KDmxODd7uPpnD0VzgKEv
YwCUuTqkprY2BaJnmOJSP0WYTmbicpcHi2lcCQ5VRdJhSqF4rRvebhpK46Dh
EtZhNEJqq+FBNQMhHQEWbqcrMgNYo7ADzQVznC9koT9aQ+uTFp4FAq77ww9t
PQ7wfuGRYvmKqbuQYt3BkdStRUy6hQK38zNBMeeW700FMucGC3Jp2IkxChJw
XRwCMAfL1LAPIGGOL/wmi2G0Bks4lvCMOAkTC13Xzm33CDzhrhocOq57VhNu
S2KH8WAeiJf193YgOa4km14WA/12U3+FIfKlGATsNADFJMohGGhuLiMOOP7D
sx2YlUrkc3H25jazcoLwIOYtIZrRbLHweG7FfIo1w3MA21zbpp1u2PMUGoNf
ZPkFY/wGaRvSt24hKuE92tf49E3zfmv/C5LpR1q8VT1HZf0sOrFdxNIbXPl7
1qU0qPO06alp3Gp0KnIrfC2D//DHvp071jO2MpRB4LZCTHAuCGof3RkUVOqJ
ohxCdBu5DvJubfs4Mjujz4xwjtHBolH8a78FUUUEt7u5p1L59vlra8hHcCju
5louf06UCmG9Qzat6GPJLcv3qyyOG39dRzUlqBPUKbXa+Y2sfsC0UfFV3SxK
jxd+6bJAAmwSzFSbnuRWVn0Fi4juSGEwQOwi7GbR7MKkoVgUKlTBWBnUWMC7
05bj6A0Quu7Fe0Qah0DKCJ1PVNum+VZNd57pjiwmYtmbfLD0roc9PgOdmHua
YMRIPUObWeFYNYuDl8zeBv6k5yvedqFCXPBc1n6pt8Dg33RUvNZ0ngr9+V4j
X4gN4knBSCl57SnCk31pi8IrpfrteIhGd1u3lpoIBFlDGfaDw+axU3HwVKlY
m8LVj10hZjhdNQw5UwRZQN6d5uFLqmZSxA/pQnG/VMDCo6N1KvhzxU5TapBR
wrTy3VkrHfzu3YU95upu+aCrxbp83vQMysu+yx4jk0RlR8bJwdbn4K05OId/
WuyKyxm9dAMKfuZMBk9oopl+iWB0/H5s08XzScPWJBrBlVsHi4aUmtkwRMBy
C211lVjP0KZ4tdmydVlvAycWAMugu+qZv0J2f6frhOKtg+q61s4nNPrTYT1I
S7B0WZHQe++Df8trftVbbivA0gdWmyyJzTtddo+/K1qxrciPSMCxlHJY7598
8PXlhOo+jPWOs9nCoDpfYtFQxoNHy3z6KhulDUE6NOcNFGBKZuL0gnk4Fzq0
2Co6S/0Gtafs7Gua028utN3Pbpvegtg8erMQXWRK4C7Vl98DdvlWGY8Db+XI
3VD+E/jq0WNLdqlqdSQu5KJCuTx+x1RFBTp419zjfb+NHYu7+NOd1GmA/Xkq
cE7vWiA5MbX7hG6rq6t5mMf/8sYNIWPfelH0sMA1JuQvRKr4dueEyz9uYusu
3qdEg8IAXPHAaQDHf3uVj7CWg3THGOYhXL0h+9XerCYT8H3SAJ7dpoThZuAa
Dhpe6poWQh+PB4Mx/VUcHn9S2RhQGi8hiluHCK9EZojzpgce5vpqUZ0vrhaH
rgbvn0aUPKKAyYnwmVPxaVtDge00FGBI8U+G6leu9y7ZFcaTm/Htmssi4khI
ci/IkePLw3GvzeEgbefmFTwoX6ML7uPA1buaGKdEqtKFF95tYKaQN8LqbcMC
Ih73awKrKxuf+kAcTBthf9FaUmuywfJg1lbcM4mG3jamJhfM+NLketFpFSBz
bqaAiMT+GdmKg+LEmv/lK5BWU0avj/vYB9ysAIwjxXMGV1X9h7r+Q2ZysZpV
vNIFg2h09hVT/Cg3qih5BfbT7aBeo9JoMi0DOqTq9HwVuU5VqixW3GzSj00W
bNX2biTsk0QMM7N6Qjvl3HbLcYHl7diXEpwjkFbARWWqhz3/0KGmjTiOSwkx
1Rs2vqH82tFf88XELKcRYqPKsaIpfXKO5h2R+9cCOvyCOiXBCg5Q9q0uojxF
DNbgEx6uG9WfWLF5wifX4nA5wLn0DryOmIdqkEjtk9pwKJbinhM7yIp5W/H2
cdmNMwwPIlzyMW2vZ0ghcJ1BvsDvc6cNhS4ZDk4zlZaxYqSEy4ASzIKRgqsR
vts0yZSKb6eOjBtsB0UOPAKlnwLvosfKPlY9XOyZH+JpumTqP/AJ3mp0Mlal
Ai9OVlL63HR1lGfvtREHjcXeEDklV483/tJhryutU7CfPaZMQ3FeFM8p2DUo
aUIvxDXdtlUEa7CfTFALehKNFcxD+5zdDwWTDHk/leo1lWI9YByJNT/w/GmX
oHcBFamvuR3XCfvMv123TnVNE2MqOs1u7ZbnLNSvNzSPu/b2YxU1j+/4Xr3m
wSYaQpnfoVSyoM3qhAK9sXkVAYaJjn0loSD0j1YYoZaSz+4mAX7d6/TvfMoF
q9VJqLxW5mZ9o0/+c1Rz5aD7nOMyqCaPve3Qu1rcvsKBAcRcMuK2V8DMMCSV
tomsJvOAue5ciWntRhTROyXPGfi3XggbTTj6s9VYJAvA4qs5uwZXFLmqN99z
TAC4fey8J647DMs4km59ddisVmKZkyoDv53lvNaMGJLSSaOugNmjrx8Y6y1B
nxU+JIXAYozfJqiaeJ0WXnkYX+PZNWeJ6cCpaOlnJ7/K/2UlwlTJbjFjOvkF
eN3aBJX5/CTZS1K5nKU8R2PGWRrvWlHaEJe9Xxr1z7VMkdchZu0ajZvs+Rw7
tOwclLv5Qw+ZBjLxXqGo4C6/FhvVRMOseKFU+9ZCosBvdGRRxPkf1pqC0iLm
vZZuld+oMTsutkalXEdpepH/LDKtRlwQqSYJkuDIAoTmuECB8z5gCDcJWNTE
Pdlcp1nRgSlqE9ICXZpCbu4mebCde5/cTpuMNIyCijJQ3EzeThJsiokI6kGW
2LaZ8uHbpmgE3ecfTmmgvhJhu792gDtZvWtGWoVOQ2AdcdG+V/PECb0g307Y
xg9SqZbm5XCK6IM/2PLCafM3xGaU3gxQc7E8nxd9LepC+o5G/LA4YqAe0isl
LMCxBMWezri8SiXMG4kkqrRN/cGwI9LEK8MT2ga2hvWBZLD8sH4Pl0s1CZcd
MXmqbpofL59l4yj+hNyolJelDPBeuCHpxpmzqT4RtRRjx3xKmBVCsyYv923O
hYzz3yunCUJJRAU541OKvrWW0UR069IIkXP0eir2u0kSjiqTolMfwqbO/kGf
EhJie2i8N40SHiBfvDVJcsuIeRfI3vD1hxxWYdxTVnZwmM7KyuVIMnBLMIll
2hQAe4pPhLflbs0Xg8j1GAQl3p5YrJjB+Z32JnUc0h+klckHEZ+CEpjPK12D
B32ysrar9r2arQ5gAkbHF4JwZeAUeJF5mOAtjGOc+CZZv16j0pLBX88mDkXZ
KH0F/mB2J7XY/e3pytzP/SLRumotWANfUUZ/rUmau6N7qrn97D7ScV6nIVLp
y0oUHaCPsVXIbRcquXKiYUVxGzZ2HYGgu37Fq4I2AbHZCX74n/11Cnq2M9Ak
U94uIacImR+u86G3o1iD/V9ufTQeOlWQ1YtpCjNR1U+1rYiWKkvaxeJi4k8g
Xfq+xwzRzuSkraa2ker3+qcyHUrr+tdvnuymHs8OOf5ZdIjZqwepnLr0q66z
C4JVGywuy7JKbln8oirr3FDmGx5QYgIQon4mjEJckK7rORKLXKKkBUHTtu4p
DRdN7QnlTqfEg3OmY0uYBYaoMGYmy5OzU6CWrQrLMvg7zBNusaEA7lyI/I39
VmySRMqdSvWGeQoXZbWwL+9FjdQJDZ747hh8GA88xLGwYGtoBMUj/LbI2iEU
h1pf11eMmQyLo9L0Vpiyp7127KVZVEyT1ghY8Szua3CuVPKMcPxyfor4pz4E
BCNVU6OqNKo3epOFE+lW2GY/Tuv5wo8eQj1SUdlYwTKfwvoSekl5lxkklYTL
NXEE2cakHEaRxZpFllTOr7P/bTMxAZ7tUIzQio235DkgP8+beU40KTt9mJ3E
nc7cnhmPBMABfzEvK1vIxdyApSiQPAkqaMpDPkfff2NHnjMb1YmPuFUEhFhi
E5MehuhtFRIEGqBO/Yud3BU2Z2l79cXh8yv41oMBGWqOU5Z0BYqHuTtV555f
Ujbrj69gluQhnENzMfF9+L8qsRtVN6UQPL4unfmjR+y3tnNX3tY6tlDQ04ws
zAjKXUetNetcz9cTI9rhomcZQtOqejNTHeBkQ50uMDPseH84GpncZ7Mwd4RE
AlGpyg+BA7Jd2dJl+ejq8qM+bfoemfupWUlfWQ64+i+1hd9OmESU+my2wVaw
BmrVnh+fLO7EB1FQ3z8KUBrQpUg9YKbCFf74az1O5jeLSwQ2XwDh13MXQE/V
5ejJuwGAR9OYnsq4WfJ7fIs+1ILz6WIrOZmx19n1WKzgukbv5eRe2wLtgtgD
xV17Mb6FCWBiRvYtNBeC8UxXFpGg00RBCaiiN/vzfR347yZ0d4Zr83bANqPc
JRHJsozm+9v+l0Fv+0IXg8ypNM3foQgrMQVy1t9P6gapkWqX/8K7NZm58m0p
tU7JV3bT/ulJzqBTVM34ZaQYJv26D//SUcdh9ASxRq/YUP//OKjtoc3VQKmO
LmvQW9SVT0JARXkAhCTBgfykGjPKqjEPXZlaIxJm89lbcZAsIQUEbvFSQy9C
+88edLcGtmuQe/7HGSehilN1v3nIIF8L5mPzomY+hnA4mdgalfrjPC9iApyc
q8AdSLyGD43sd6g0PzkeJvSVwcUuKDWBol2dnQCqg4Azbo6njBBxPAbyhAiL
kQcAUBT9en15CnJqE3Gvv1sUyO1f0Tef7iiVrJ2T+96Wb3elglJMceTV7YA9
ryKZutotCiNVoBFlBC1NWRu1OIjfKRBhNMZCC52qebpVwxRuUnhSQeJCZlyV
2TOsvQ7jVYWOUuLd0dBVBDWbZpVSV/9Zf+FqvCPvbRWV0F5abLtU6BBi7zDh
GQ89ql4I2EMcAGG6x1DKqf3ZueRq7IFYEmlltMiOCx0zWSOe+OXnVAH8LqK3
D0M//MqNhruHNChC5vR/DRrHYkDhe6Y/TCcHxoagwAZr8btdf4A1mk7Xle2s
h16gSg2SSlCGObe+TFzGdHLk61Omoskss6VobhmqJNrDleTyK7msdT3yIcBq
nbtIR5C1i9rbBKbhxK2UlrTMwG+R87bPgdk/wLI/LdsZxVK2jegb7qGYbMnd
PnfF2KA5KPucivfcLsgw2Cq8HIQAeAYC39nmm1FZDYaeZSTnuPx8hGB1YA95
Nmd38hwI6/RJ9B5PiRs+5mrJSW0MAMYl2/9IHW/3pRZ+F9lXxbkQ+rK2aAmt
FIGQZE7gBorDdtHriMP4nE13PEzKwke+mNNuyHu/V+o/q94zvpsJVasqlII2
vIg8+R2sb2vbyUh2sB/1PrAzgO7dzvCWqSkjgC4Je/P2s5tFhldFInxr3Dvn
reOHcHtDoU5bPPMOhCuyNPYkK+ZkqwkSewmNrGnNWmTYcjzol/JzYpnB3GDM
mDI0yv4qu7jHDWjDkK6+76Xhey9+wUC01d/Fa5tKHA8p0ag18OdeN6+CB9G4
7vXCDb2irSUV1YCJaW/ToiAgXNxCEC+Skbe2QU/QzOz5YVs4vwbSPkSPHxih
3NQv4zG4IiS/+e675CHS5Jn13R9xZqKLn4wHqPhqwwgaZbUTJofnfny/M/3B
4KyLwMU3TS1g+Jomjz+nsSwxSWjfWjZF7zfPNaiMgnAE9pJ1ls6OJMZINKVi
zSkBYi0HqZhsKq/f49O4qSG6EFf51BojNMvaQL5Bcf2oH+qfzwY7lVW1Mon6
3j1VASu6ScXFUPfICAqa7SHV8P0UP+letnZkw2lTh0V8PpVo+Bf9xp/szZKX
ATBsny6pcP7l1snb9LxJZFHgVd76ngZe3vcBeVOyzAlCtLk0gB9sUgrtO2/2
KYcOziTVilQy7yyhavpWHnSf/uEuYolE5kkBZwkfoCEFteFT9uM7X4GbDJKF
FuNi9H2bPlCsFJe4IndeLLz3xuyMkzJaVRK1e7OqXpB7IsZX6NDCjT3fcjai
UkvzGyiqDnmFU4V4SXLqHOt65k0t93TJMRsvikoCUmhWirO+cQV9td0lGhep
SI/Gh82Q+UY+hErX/Avzwtxy5A+HucVq95nn6UIDVJa0Mo0oLi7TOCtPWjaq
T8GpnM041/muROsDU69GX2Y23Y02pb97fYfcZG96vF8odaZ7XOL9gW76gTPZ
Xiz4VRTGpssU5wIsOWgbK01EswdxRtAk7xRK2kg1l7xYzmO+8ytVB7AGKBA6
FV9/sJ5NmXPTM2tXTWNqRhgg4GSOH2jn1j1NJAB4Zzs95AHJlWoiC11Mkypy
S6RMVkUFvrrvGx0t08JSmgBBgwu2/Xpmg08yCmal+006Y1cfqrK4ZsqSGiye
zyAcc4BAYajGWTtJeUSz7VvDEqjtZRr8XqxNxSF45xrB+c0FuRMFWbvPEgXG
lz/0T87Hlm8WgajVTt9ezwi+kueOoTvXwQWeKOYSP9Qp//wEQa+bC66x+Bis
2aNCfc+C/7FOqYP2cC5hJHvnigUy5Qe+L+r/RygFq9cPix+PDBSngvQoBiy5
ferFNI05Nr9nVUndTXFRWLtaL1g2wzUJEaX5KQEwR3209JWZY3LLrWiK/sMf
J3Yz0YBgrs6hgc++Duevdg0Z4/HXoSDL/Ip30k9UVfJmRm/qpSxm5Qom3DXs
VNjvdxmW2zDwnT3eP/QKC5Mn4YvRbmRGy7Zu0wH00hmgAfsIfzdCvll2AMcP
wlmaurnSVgaXmVUW68NhOYiIwmIOQZyDtrLtfG1e5xbxANM8Fo+xBIRiNZgI
kybWsuJc/vU8v7JxvAippon+Vpa5b4qxaR6wn1oNehgMdr+D5O1mOB1rRad6
EeZ8ioiUbzMqtaOvxMQjVcJOvmSzEyHm7UT7IW785YstN1fusYoKeUmb8hF+
V/y4YNrGc1X5G7q01D9OKD/Wujk0qhJSS/azu4mrKR2kT3J2XeODywVOzFvB
7q234AesJmzfEu7zGIBQDqdGYhVt/oL/FDSmmofwE9xBnbU6oueaC1MuqFhA
a13+kLIXjYDxVGqCWeAlahZcc0vMi2D7uu74WLS5yk9uJSZjqFfwEa4XAmMA
Jpsg+s+RVuT2fK/1P+swTDL3/fdkaRYG8OOrjKFoZLgew6UyEH3au4pMxi6T
1jiE5Lx4kXYV10jJQCuI/pO7Xp+8e2l3gr2NuD02RlUs5l655K0Dt/tAwNk0
yJgkw/2R8XeBhtOqV6Jb2VmDpdoHHkLR4tHJnaZqXzT/PcRnMuaQtFw5T+db
45y4ZTjtLxGNAZLhSdE+f5Gpa8us43SAuK+q7+co1i8bsYg0l+UvfPsSnnVH
e/4mlY7fg1WaKKiK+77+w5WwirptVEkG+msFq59KkOPKLhQrc3CGaVA5x+ln
0Ev2pkI0ydGBLfMDAywA+jWetjI9wz1M9ON/RHT4JmNI+0hTmzNHhopm7A6Z
59/TxPMD38ey+hZ9I3/5tvu1o0flfvm2yc9lnse1+Jre0svKNdvjABZ2wtWl
lTeCKg6WdnpPMMRqn0cPUzZKriLr8jxIavxWzUVyS4cNppiaevJQrRfMfJfH
lGJgkUiIYeoPf9B5KdGKCCBeu0KeRJgHqG4HC8rxvZz97aJ39ZppdeZ+K0wz
cyJtN9M+c1Ykwbk4LCT5i5ct6Hf/c4iOkhlG/UwzaRSzo1IIQREE6U05LbVk
kXwAnuJiLlCbjNWAouDYmPth+LDKar4tAleJ0Lj1RouXc+eAiXsnvwzFP5oB
oY9RJFNYKQWBGeoGXIAAWJsaaAdMf9qMnCm977ofvmB4dFSKVOO/L0ZSoXNJ
A9PjK8y9ATRJHdQSIl3ku90v3JphrfBpKw9L75S1tnz4rRA6ASSky9muInMh
SojRl64XSUXCNaQJp8NtmOv8YwnJhqFOBDozlJQPb6jhZ30vfnghi1Xcggt1
+ZpJaBuk+UMN9efJ5jhFeFQx+rrVGF+F9UtBuV04l5QBaGwTP2DJeJRtm9Cs
xu5maI/btrgvh9MTNqfp/zwcaKWGdcOi6iN+BmUKXuRWD+hbwzMuqYZv8qHP
nh4MiE9940rGi923Bhcy2NaMZPxCKwQ5fXHb6aIGw0Tt/h9INXJFXBLH79rF
OSYYrmIvE8NfNqEYZG5yjURADQdhM8ZzFa18vYcS2b+OczRHwcbXnTAmBETx
jukat6/dZX2hlj7WM9PYPsjrh1X8z1sTgI69+lOzul1kAvJCEtoSt9uCdlO+
7yGwvrZRYp7p1LtNYnEEDpSVgpcKZCHuXk2dl7dxCmUQrLCTrz5Clt9/TPM4
b3AgVKrOkffe+Mr6wdyFES68P0wQvX8+Hr7xdEcQCuo+DuYyGvWOi9/GnGwy
UHCVJcs24fVbXqJUHAcDCaCYRVWMoA5Bml00oix5xzMUYznhCeutg+353kPF
mvqOg+NxYR5c+JaUPJ1S8QExhk4pXvVkdc1o0ZfY4h8g2HHPX2kXsfS/Af6S
Xg7MSu9MXIzwjDEWBRjppJPviZP7k6t03pM4gwECA3j2ABW+w0sc2POt6ceb
72DIIcqmvxjiXqcfQOGSXGdqZihlsvbSO9eP9YyqV9x3VZ7YFCDxKedQdrKE
6RnA4kvLP1A5w4EZrAFCBa1SwN83bwh6VeREC0CkyT+MrsfSUEfYRB+92Av4
cMm/fkpqjBmVm1d2OLEDvNw+QyeGhLFvC/MfUj2eTKifYK0OV8OyZKa8Xy2q
IwBfPJLSJTnFinMN2kEP+abVaEx5QZWjk3nzbNjFzVmZ0GwVLXbGJ6MCdA0p
FXt5VQvGggwLuxKfsCxxqHEOhUL8vqp1V1rRExoHSXl6bdRkTGH4gVCE7lvZ
b59LZNH0LJ07JA0Kyr19/sdG51FCM9VL2HYv0TMA0xp4Paf9fJqSD68rnJR5
oAG16xCnPySo44o7A0HxAqPzRfsg2fXbC267jxrT5SxjLIJb6t+yZlBeJ5SE
YLvGY963mbtXekR0X+b8qIwJ3shNPfDrRMpl7jwWAF1vQB9fSq9gBAuITENt
wI/E8cTI3UqtWHmbpQrikNl6xjwf4CyBdcss0QF8YHI48k45Rnbb97tewCis
E7tMH9qQoJ1BI2wlRddsnrhmVM7KZIGz9K7uuodnOfybQObNpeGlY04v5/Sa
oLmWYC4I+p0LIWJZQ3wj0jyS+b3fctXPLHdIqoSRKwvJ14sdX0UsR9ud+/0q
ese+LLNMkHk4AiKMdrCv9FsoGn5o4bvDY+Kzs11cxqi+RgUTrnKTB6UAhxjO
Bqiyqi5dt0ztcJp3ZHdVXk0c9Srugh/Y6RRZWdqb+1x1ItdoxN4YStjWv45X
UHRr+IqpqJthptu0zV/zJnEreZsaMzlv6Z7jlvqrNm0ZwEsjfwLGvQp4+0q0
psfQIDFqrASXCueicxvf8yo0itrWnCuP93PLt/zb5RZtL3qxgRVWcF4P8oBx
8KFHlI84MTIaFMCfShEvRGl0gi2PaKSxiOU/G2bb04brlEZI6L8pqYCBQtSS
U4Mx2qva9pICPQDG1CJID81mLw/Eg/q1Vqn0DmWUcCBR4BKhkVacAGwLtOYm
uswubaVqjPmJ+R++pqEx0GPc6ISx49gzwkaCFr2R1+jYfzgpMsiR2QQH+T3U
IXEx5uHzl4TslJjTO8GoHaVfFFWUJDW9OxFqi0/k2lZs9rMY3Ecx2fGtD+9I
BcZjLx6yoxKhIF+nA0cwEhf5PCSp/n4IO4VyBMLnYfjZUr8Exg8ZLSeCllFk
3MWTZFNy+UADB30VOeeeiDtUpPGieS/lscfg2gAb8VipfeY4ycGHazkwNpVw
D5LHENa+ACRuwnHzNGS8ol+WR3Q2ex7+mAy8Z2n9c5VVQec44W1gMPgn2Te0
KDyTyeNj7KVSq+LFIO15xeBc1vPqGCha0byvy8XvDqlr3Lp2XafDqxrwn89d
c8cdSTye0BL0XaCbCmNDdE1DuAFHVg/ROuhlwEQjQSeAFc0t+sRN7rdSk7Sq
cDhQeMbphOu/yUlCrwegY8V6/Fq2eoejIJOQGPcX9n9gmg7mX8u+MZNE0u5V
D7Ye3l5sRsU0p4ZwueUidIR9CQTxso6nai1Wnj8OzPWATz2mrTYsD4jQ7Aee
h/7s44vCIAfiZxNkNz4Sor00w0p88imxk867Qw5ozD0zVzAQfj3JunsTQ5sW
rtc9ruzJ7XiF0JE9gigKSCsmjZPResTxeCf8x4agSoP9eYOxe9169uwyz0ci
5qt8WjxFjsoWGQG65wzwEXz+fLdNdzblY8X4CF8n192am2q5pvLM5y0B79Pd
zdOpyZccPdNlgXdc5HBexaFx+GiNrSJ93kt0WeodTNIFXjUDovkuLk/9GkKJ
oGPWYGO/fI8g6i4X/nONXoZvYCuvJdUUnRwtWxGcpLGFbZuQmTpxw04U0FDl
SG9ilKynbWhlViQXvm+XInI8QKbM8V3eqeSiToZuqT4SfLfx1DaCQLtwpeK/
Qmt5UKxyOYk+9AkTmY8iEbfJTyDCICxWrlCPB/hvKCLyr5FedngNbuk7sr16
MONyLQXTCLtZbQ4ceSKsP0FqAYScSXFmUV3sPyRVMZ+IvJT81vWMYT5+S6nn
oIoPsDhiudszppO26s9yjvwc//Zb81DjvUPXSP24qEZ4utBZMJHdvHubAOtY
7ifkHb1vwLzXmU8PZgzSMVZGZ6bG5TRQUpSFhY+r2l2/91mVPlyry8qe9FZO
44QtMkLw+Uc4wOFZDdc6ULr1gOcLtVKxBLGT+O0zxayZSqwPmT4YRmOPISX4
rvtNTn/Tq8vdvElD4Tr1Ucy/pJ4A9ydS0cP1Z1DJ7is1c9LPDWyASO7R3WPI
nK40ajEGdMRkhxoofCDMT7nN+2+JXtwAhcWbhkvPT434TKLmGxcjDkGYKp5n
yO7DVjZTHCD9WpZlEZUi1/AzWDK/LCQ0ygchDJEE52KjX6PmIzDvwhS5dG7y
A+dyTGReJBjGhWembyLkosaQgHZmHZuxbqIhajBgNqBptkD6tcfvU6fFd3zz
W6ruxvlicrs+SWzTTr2sLxS0MfDJbeXC7yFWM5zgs7E7y0W7xaeRlNL5iQ2l
3/Eb/eUAa1mIvdJzZM1HCIRtQpEx9qOyopkasFfZWAt37ov8NYuRmWhV7EKc
Vetd+TfINiWJhWsu7s6pkDXLB2AW2zTmtiS949sJ5TFqoCn38pbKs/pX0aXT
/BV+JHv7j513eWTqKEmkflK/1WFSCqRaWqld1EIMUMzs+etiX9W0MWGoGT58
WYfqnzqGD91zmJ43zPFK/Iu6vExiFZo2xJAY+S4+KiSafRYijYKuuU5ghRH8
DQg6b6ZLSRkLnunWY09gegEFWUFLf62FXznltIXKmaLmGvXs571B+YMttUuL
uqQJnERgexobSlauBOh96TsgntbrgpHHpuEv0P+uulB5EtcftPn7REvzo0Rz
gWES0NOGtJExVS7gzBeDasry8QqFAPIg6KEwujMPpRFygjrlobMW4jrJuG1U
claI1ueIQObBS2MNb2RgmvrTEiw46lsQUxj74k+GS1VVfvAERsKaMPDXROdG
+9lby520zkCdmkdRVwehqD47hjaRsMfMCkYKnJf7hmoWhR3HNmPQ/bclRVLa
gC4yPMQxP7ylSfiJwF374GRjWf7KFX4dZatz2d3sIe99S/QqbhKqOioL29qY
uamxDgNgKE4zDFmta3zpNvnEak7VDZwzusECgN+U461UxJAV+dOaBwwv5AV2
cv6rJCOkN/8j6hoRborBKPL0MCnlbLk76zFjqQWj4RfB2pzoiSA5Nny9MdLv
InZENkCj75dZ4iLp0DMlAF5vQkSLhHTR1Wcbw0tdmGPLvHeT8ZFEyEcjvdZE
B8OJ6+YLqB4tSkQS45zn5HuSmnws+7wjWyzueBxGQSCH7NL2DaiwM7N+9zxg
wDqMqkJCgNyWkBx1wZGJ+T4XNwJF3cXiR6enJYbQpybIHAvTG4vxp3XIU4GB
OnCoi89bi2HnFIEJgUzE2rP7YpPWxCuT8i0wTEIiyHk0qZjgMZD7h/J1Uf+C
jq/9j7DOoAn1DYDwuIW1vAz2OPhLMv49+jTI7/q5YuygVnYfJqTn1vQI10c8
zRwDMQXW5NoWa2XCpd7qIR11srOuP9uRqS1urmVdvUo3RnI5TJBouFkEAgFs
1zDL8ZxG9qXTin3vqr86n6dfQ1g7UlXoV7e+92rFCV4jjhQUe/+gmYnRyCia
6rm64+zpi0yikUggPvONE/fF0WO722ywlovWY6JqMmTVlbphm9AZJ+hjpHa/
QZgDx6Kj6MNWnQ5LrxVZ4HbmruD0CcbDHOnb8i6MKVB4fWEb1GNtJUkOkG1g
tGyppsiUUUdIZ1iGuSKNER/SRh749rJdEQne6tx60JC7RbeMXnLK+SWeDBay
OuXqGYwcQQZ3wFwefcBmsbrmWeFlHWKjPQi8pFOdOQZN39wtiXeo1dAcLn0W
27vRCjW6DE2w6KYlkux5/H+nPmCuEE8WeJgAaitJ6GqtCegaLJcleoyC5U9s
YCzPpvgjdchEybtdL9pibKWOva8FGXk1h7Hp7b4LEO776az36mSOLrmzkQOS
K4dLl39Rur+3Zw3lKwuY8SRuLzwsu08TYrVVhDP9XyuDMmQCIWJSxFz2mqni
0vYJj3tOVNy0jueLSm2f+EZk1hvf4QW6960YUBCFn6Z49S7brpYRypXLmcNZ
1RBGzgs6Jj16InQ1cxs08tigHgTv60n9lbdukD18ayJQebki3oDJporKNS6X
YMFdvpMc/5OIi+cY+2bRgqySjv77vHKk/lyvss4E7AzyT8RoO+CCD8KCdsoo
h3Gn5LEkMFOTwrBGYYgHtyr/6lgdgC3aexgq5pvAL8atDwWkDdq3Xtwjdebw
JP1hw3JKVkEWm68TPpmaCyQe8AoHpPAbsPtzCDX5ARcCd+cFjXgy2hF+KQvK
1fq/kONGxITZl1/nDNTEYarQpnTz17oHX0vhxVZZ3r57RDojLOe9eGokkjz+
s7eacFvXwwAwNcPcFnNJG10KwGOMxTI8mFRoGDXQUu7teA7nkIOwSPakS4/A
+50BZxihziX+xxs3ymcInTGCqi3nmHW09b6yk+0KjLw9AWBx7BAi43kamITa
qhbalDidK0IET2EZTmm3p1pf4pEc9PfRF9lXiHsRwj3MRtnVuUCYpg1WhJm6
BUNG2Fi4x54eIkZHLi/DQuqq04qnm4BB/wH5P+v035UOkWKOLfeP9e3VAHWa
qg01NYIXjUiZX5Iw3aU1peMbCVvgckpDJEb5guV3v6lHRiaCytMdW8Sd4LdJ
fSZAQ/NtHMd4JeytU4tnlHkQnSnUJ6NqJImiSbiqwW7vieaXbWZVL/j8UNCu
Ta3l4nqSP0TAzLjE0Arg/mIkfoqcmcqSpHvw/37SCJVmC1wSMZw48E6PIMHA
DXLyWFBWEhFg6VZAoyo+Jtfx4h8kPMUi+8zUmumVzpwLk2y8aioMQyLdnZF6
vlTNVSbEN4G1W8NH5PXDgebsS5qlqDoIL/W4WJHXPAyynq64H80lTQxN6UsH
giYMpx2mA/QOyqJjggD7/vw6JsVAaaeq3GU3p5ubMOBrWUCh5VL97o+7QfEU
3KtJRJu7T0vuXH7kr1ah9VBgJZPYzRYGPRtj0sApoONy2K//LNfnZ/ZKHD6U
k68yxp8Uig7DTBt2bWmSlHRo+ux4Wj5QdkiLSzRNSLaVTqjUQNATrREGge4/
6HfXwFPoTCnn8Bo8qg8r2XZkAO8ENNgSKYKcozUXRjJxYI+QvcvGEq0wBKil
xjiGNAgpaZuMXHkhR+ceDFV/FOAnsgqcx3C/tpHhMBpSbG9BZTYEf4Z4k1oC
c7WXVlykxTgtXoW6ZFANv73peGlxqeJeb4Ru9np5XFtSqkzxZu3kWVSvnSi4
CmENUHgxfz87E8nCnUgbAe/qMzKSQQNL1ge5c85ftphEQrKY916VdjW3CHfn
4O7iVUVLiOfDzpO3uk9JHdt1QKGF62EQkC/9ALxTok0J+4kHy7uYMGmj8xCA
oEwIktdtC9FyVhvoUFTA3l8klIGw9KsIY+YdOebodGB2+MFwBl71NljmTkxn
nvBi5mY6MiwcwjRdV/lOFulY3B6MjPpXmQ0pBJ50pB021rgP3XkbM/eBoarg
j6FhreNGv0vwrYNTOJhitt4UIfDeF+BRqV7vVRFj4sBjaCm4PKkiqt2EuCs7
aUfyiDN6Kp+v8Ui7rx5JYIqci6y/BlnCKaLg1LVaVN4kn9Ny2+cgeSEu5Hye
nPNjVblCDxibJaz+8SJxctN3MUg6G2nGdkMHtilNlbSXZlDr9Wffwf3FW0RA
EqZsN0GHCVG7J1UeX0LBb3gsXjutgk/n/G8zLTw8gX0qTdW2yJldZpWMREsb
W7KjV1jOHjZs088U2JTZRyT8jazAK9OthakhCBjfeXY0AzyUmLUVGI1rn5+j
xn7eMK8qwQnCImn6hN0v3yW8mkgCSKB4AqCmfQpcmtLgbV9+/vuSJGL6KnmY
pMBM1lK3ogJw8iKHWd3+ZWzYEmkZLmjYNxTYTD8/pEqAYscufHZdFtOh6rmG
gYC/2EXeZptFhKMoQ/EgCv1xLEH5eMBaGtkDHdEjVNEfDSMdaHBQFk6LYVen
W3wTk4CgW9fabiBKrer93UxFMf17nnbzECAAy0QsoVDE/rs+8ddeqtflkT9/
SaJHMq3Jxki/WKAWycCPq6TNlULYRD1+iCE1KqkyLrDj3vMzEe0VFJgaNGoD
YWTmCVuno6Ssgy/Xmk5F+IWOPo6oynbN3JvYg+Yn/47eJq0JW4jO6Qax62Jq
ZZs3E6WuRXYRbgCKyWAi6ymQ2fOA/8REdWRzgCagGl7eOWrTtC1kXMjZuRiP
LAjucqMKeJEspSVTseiqhWm1CaYDHDunmYp1ShzSk1xBKfM4/GphY1OXZxIn
7JqfSGqQot6bVMZan/s4lsm8qRhEALQJEsPDg/TP9Vkn9zxANnYxMAx++yhd
4O8yOoGOugqYSSHoA4pMLfi8Dgp8psdxDQPdRnNhbxm2pp+f0v2vpGXBfYuF
c00w97p60C4D3kBYztozF1XCZ8vyFR+XZ7WLcnXAdsL5vpmXbEV7IWdnnsSY
233j0yaFaD28yKjoTDOSecyx4sk6C2KGoUVl1u/HRvpOW/H3OheoIjuOUp4v
Ual1WcNuTlb9nw2ePg3W171j3A4dMtjQlSFqNR62XqBGw2VY/FIzfI5fKMmn
ZS1Zc7kcdtPkJmTUJWA0nuXDvuD9f5IYr9GvkYperDZajc2y8smtZ+0P0O1C
2gDipQO3sxOPo2IxdSeBZ34IZOHOUkrRsfLUWoPoo/vKiO7UsnnRTvu495mv
2FjDdZOMX9NskoXim077rEme2ugDQSL+ioaOoU/U8D4IPsobwe3jCpb71MwW
1/derURzXRJNw7GWSSHDcqx3Op0Bs96gSM/HR8HzQwDQVlKP4l2kipO0b+sd
+fgv33nvSEUBvSvjm1ztjnbEOim8CWp6V6E4MB+jGfwBrSQuN12GwS+83zde
wvj/cR+O+C9/yvkw76NCPahOPHs0ehNxYJ53c905TioEcy4M4FT6HPvXvuqI
3ZP4FO7zpo67mSIA8UfD3rrug3aetAppglvBzgqvBEb5tFzH+8XuEu7NxdSz
2VZi/Ndd72vFjpxm8L4nDzDFcqYc0kPkCbf9Hvx1doDpFZXGbs6JHp5S2AO1
CY2Y+iYNNqhs6xmgYEVPw7ZcaITAMonNpJLrKN+oA+yyvYG0G243VII2vJrw
rVnkAZpLqAFjZYbEVLq1yOcvLMQ9uXz2P/rzOpfLP5eKTDIZRRk72183RXb/
UYQKTfKfxTfhl/Rkc1FZFvOWYpFr/NXkj/Q9EHnNVrpOj5gwrz2hb0MyNDsq
oqXYKloPNvzynoMQ1rVMio7VfnSOECg3KmQ0yEWI+IuAkZuQ9mymbJ9hpCVl
fXOSSS7AL0QSsurXW0O4LwpIk5R1WPpN8+tGHRWUpeHJbJUGtd8uevdpw4FA
aadXNk2AouaDVkH4aq53Ps27JJHanGPVPUzb1ZLP80bsPXSk1Mi2eGj94mbZ
3V6E6icFyH8WkHMwsEo4RSqS14NZ3GkYvp93+l+n4LpK9vSEvSTiN1NcxLP/
DWLO6s/ODoXtrhU+FjZBfXtSVwqFo8quykytA51KRhqNbnrGGWBj95vVxqCL
omgSy5obupwtXUEg81i6pVmcxS7G9P3rxMnRahYByoYSXe6bKBKiP3anOSZR
J/hyoT2uANkZp/PjDqvW2oAVesjkO7DylaI/QiAG/HzP4itbl0ZK/hAIPGQh
5/ocaqYKFuyShmDqBPUlpB2LatNZfeI5gHv5ihbfdz2oPwt6mNJblc63GzOl
DvdCnRbwQPJbKl6QjFHoNCrVFu6xcrs3sycsVNQlIQJL0gk4LkyOi9dixIuf
sFSNzEe3uzbttKD/OxO9rBXjicU3rgCEVToQt2ykHhy7wxzWLEXCxUfQBHzS
qlyQt1zvdd8wqGl67JUzSmQgb5tfisDOhibXbcxBj7b2vTPOVj0JgdfL8eH/
8AWjB2IqAMJvpxMozGvE+RisjUrE7ZONUAW05zYbmgzIuZntKO7CCniPeguY
K+h8/o2OErMz6u38BmLeUSi84hbgm9xSqudp7mqP6NkTFyntPn9ZNGxh+zGM
E6XzGk3wvfwiRYBorfWAFLQ05k8KF7bBxIQdF6da0bIopnp74TAZh7CPk4wP
sj/mxlqj0czNnuJ4XhiuTAKOpWEfVxWS7OMDZgASoHcJM3wY8o0u3CMrTM18
EFAxEegaJQZ1zS30AVq3Ym1laBzavBSiX8NdvQFh23WIkdAmp0/HICpmiYce
atR6nu0v4w70BxJjjvlVJxFsGtfQ96E0Ih7iDzHuhUCM/UcEgxjGVA3CP1Py
4nrmvuF9M9x8uNpSGerx54zcdtGwNuFc04X3TeH/whOfXtakDVaE/cLooi/y
dTtQTQpgK8TLJ5jnguiqWoYV+f1a6wqHFD2K509FaDQDvalckKYvyOBp2cWx
UtbVHU354bpEdwPLS1WzYvn/BtvDDMEjMdysCY/OFpynIPtgi+WILU3wtjGk
76AuLdDz/inGU159ccgmmqmjqohXSSkaDkHFG7ZjazPf2eJd7SwPVtQCF0Yo
QP0hUAg/i2fm/+/S6q+IFovU02XMAl2mtnMiPO/0plUB5Gky3YjsKUb3hnoH
IwOtBY+8+C0vMtPmKUildn7N3WJ8Ycqj44RTMboOzCn1LOGf93PmRqRJJlUJ
n+BeECauu5CY6NvozvoZeFLoZg+zCp3iOtRCI/DfDMPKbEy7Ia8aI7RwhncC
NBEYVwz9VYkfYYXritiOGDUIRL7nEghv/c8XHPfDPrUsR9Hbqlnk/FH5g5I3
c6fWYjOw9N/ngXEX3kJu7i1t3GpqgFfpfhbZw6czTdDCTrP386cqsad0VXO/
t34v0WQITp3TUS+n+BCE9uPmiAuYuOyrgWdfyQvJXbMiZQkAsiGRamuUowQj
27NGCh0zMba/50f3VGCDo6EJgnNH82gimUHKqeI/Ch0sK6ylIJ6xFjbZlXuQ
m4gfnrQyBFBrIEE6JHzCH0J7C0/fYbEfGuUiis+x8p/dE7OsxZms/6XHIiuu
z3w36WMp8aEsH9LmvYIF5Bnem8LT3h59tngIEmH5BtNA+VskNkIDXquVQLjW
667/OQKqSWNvM69sBINjU33JSu+LdOkO6iawgSN7B1gAMT3Bf3qq91tX7y5i
gkI/CdBzEB8YTA7+00EkBgB8il9t8bAZimw2zIdPKKHP1bUGqB81qWkdUd7P
aEuZcv0WI/Bkbl518OsBcQitkECln8qAZ/D0UzxFkytea1LE0giD5tnCEqDt
bkRJFq/Ox+3sKvs/wr5MPI4KHsIVoKYVHy8+5lXKmRxFQZYmWP8NsYh4kC5T
65/xwQjxKyalMpQYIcgXblpMIBgHD1i70B2dmeVI3dYzY6Ug4NVF7btN6FxH
Cy+fnWMKR2Uanadr6vZ5CWGDQ4C5tmGkwtpmAvk1d95fso/VedewGxO5lpbn
Pg295w14/6uSnBa5k8B/UWZQ0OB/AZOg+V9xYS4GJSExUbA5MHm70j8F9V3t
TJWROXdBk3Xh9DBZPJfYjScEXm6wfHJtqcFdxP+nDyD6sRxbb+rHOp0lobbb
Ll8u0TJpTFU1B6a0NErWNq3GsUPW8mdKh9/OG1OsNzoc+OBTVc05nOnr5gG2
r6KEL6LVdZLdpHERvyEm3vRZfSYPHcuxfggocwqfnsyJeIKU+3910F7QZD9a
gskYJRr88qUJiw9YDNBk0pyMgil2oRqAqLLYHRXJFnUqYR52MOXX3iRfv5ZU
jVnZALbuixPCnWieqFVAtUJA4zQnuITVCiz9b5hm0OBE0aN/c0B/ek0zoRaj
4kAio7ASUCkLby9lANVoqHha9uN5/YXqB4QNtLOn/ARC9djhfKoTz+ZX7iWs
PqfaG7DgSv95/QnQoakovn8SN61W8uX0NiDWq1nFDH/a155cA2Kug/Vv8Wk/
05kSXYb9zlYPU5T1VJV2JrfG9Rhn3PjkZGy53HUv/bu1clmTFPx95gNzs/Ke
tX5iYEfYUWApaPkFyDFNfeKE2oJytfXDCEEVZjSQf0+FQEgyyvwzTN5yi8N4
rcUbRTWRrQwFZ9QSCMVfJBdP92JkrCE8zYWlFWJa+QwGsdQUvQO4vpMmF//h
GT1VJQkoowdd33j7LNeAxgQAiCNupT0IUlbotnTtQ5akGj4cj3uZ+WZwnueU
2bdhpZnhrXxUVTGJu6mb4g4RsFt8L6lzXHSnP9hBldbg9TBPczg4NKV0Onx/
Qk6yanzdXJJJ2G6wTR+31BP1cAQo5jVHFDSPLiaxpScfGDTz7QBAAu1Z19zp
LLdrowLlP7og3+OlVnVB/ImZWlOA9/xvuwhf+93awTUB4MBJxMemhwj6ggHv
A5NPr+wCh5rgFMoW/IDZuhvwHUe00sS7SdamwKgg2B2Ywho+V4/eAY0FFdJz
VwM+ygyNysgvmi7idmfhIzkkdaaVMIKN8pj6yWs6wfhCNk0VO6Bjaqww1aNp
ubAwnlCyFgTik4e0rFeY4pxULa0zWo0JR00db7YI5hrCqYcyTqkxFkHFaFN8
HenAX8EKgMBG9hObLnsT/uA6ODE7JOhGE+nuG1wczGV7Wr/oe9ecuQbe5tG2
BDbyDefUriANhDyMWjL0IOsPYyaxtW2X6k6rlvs0djCotpx6vcBwSnJaX6Gm
hjSK9rcBb+OMRwtcpmqY8usPkUhCvQKMj+ax8Pd2nWJDdJBZYQlnAY8siZ+n
ShG7hVKwK51qpFFOg152k4tLFAWLSHqvSiqR1PZbFG0p3zEXpnh5eEoYflqD
hMvucwuPCGy9WOBHP9SvNtO3hxs2nE+hN5eMly+ZD+0TCtW3IhTaffhqTpvj
yw4kwKaZ61Xigp7hi7Jbg3vsqpoR1sQTU5V66MMMtz0R73o0CnijG5JdKKwl
YyVwEFDCz4TmScU0BseL/en7jCjRfIiv67HEaT2F0P+QO/ddJTg+5+tx1aog
QsyZnRRhFK5QCSzkAShOdyeNBjHco3M04N19y4CymRrIID6SY/DqI/L1vQ6C
22tqXbcXOdnKk/b4sge0gdycpuvG5DpcC1rgMLXsykgBK7EegWFjkrQJOZ5H
oyuqyO4394vnCmazybfMWJFmskCZfeVt/g6y3pes9PPBiwdpSGQWrz80EHYR
JRnCKnNS4U/w6F5JGmuNnEOh55XG13rNLFKNfu6OYSlHyJgM2DDTnbE8YwuI
t9P2Ji8OzyJvY7psTG+wJiqOsbEmlbzqjCeO0L201u/UuhfB1gYfTnP51OCx
pFP/Xv7Ic7//XXCVur6lgKqDbdOsskM7FR4SlA5k1T4Q6UTtkDc24vfxwJCg
qlOJcuoDiv438uTfERaCcv558kW0akFKSA+kwjKF/FpDIRApwSk2NBeVmnZl
ABrTbYc8G24bePAptBbuwA8ggmk6CBB+7LJz5lqiINj76mEvW3CWWfbqRPl2
YdpcKuGJSdBozmJmD4dY3JrO0d1W4QLi8c77VKmOrAyUE6bV4rCYFn3nEF+o
VEjJVQGLzwkizagrFJv6PUdpGyHvxz5V9v49zrwH7nmHjOz4VMqDVX6otv4j
A96T1LAP9Kb12MhKAyB4H3r6S9W3qdtfvYjOqNgjZTdZlnALRaQIDvqO7pmI
UimBwmBWfK3dWpz3pHqnLF9L724dY8bMbBDzJ954k7TJqGGIlw8z6IjYyAq2
+KhIwE2nnT8T/usejubCvCeQuBjmfKKop6E2fIDb507BNXGquGOzLbjVo7pG
GKRDoehGeHz9llk+s6vQkX5UyzkoEkiQYyaPLJqxaYZnJ9jgPge+VV/dsd5e
ILCk8nvz+gXkDRnJDgkOwhrrx68jsiSVb3qVcb2fb7P3zcw24IuJcu8oYLiP
elkoRj+2+R4X7OEGJICvtdBjRq+q4tUVjqLgIL8p1wHHGK+Eo4i1ckiwp08Q
dzSBxX+Xa87nYT3DR64XMD2alRcqwEhoMANLzGTtNS4KpLRg72M1L1dONcCN
DWRMK+KbxthOk7OaOpDb2TfmALhMg0VAqDRc2OlCbn9rW7odJkY5kpp672gn
o5I8E4zAJGmTpxoh/XO6Y9S08zyH86omh/x2IXPfhUnhtUl72i0JpI8B0LDn
yN4Y8S2EAvBih+F1D65iw4AMwCWnunii15FLCbIOYySBWWIBNLFtcFfDadK+
qMzBiYGgy6iCZktXFfQHfmNjL3t1OglssyvgXdO7zNj0Mhs/LGBWjJ4rvPAZ
JFp7qM2czmQOJgHQaFL+ev1BCYtqjlFYXCvef9CMNTCmXHgO0tuQz8j9XpWX
/OZ2II5JJcWH6MauRmTY+/MYWLSCkCtTVabu9Cd42DO46DvNmU/U2FbboZ0y
3W9q3L4Y4PN9WnD8rlfOppZ0xdianmOqawQOhsrcfOx49LQvRFD4GemGpWzW
ocIN9hLU8//DkQWQbPUm6gd2rsdXmZLsGfs39X22E2tH4ctg3yEs5VbGdzm5
/8k0b7G1c01M7FhiQvCXw4Qp7gXTIdUTMr2rb3FUzDSWIlBSnp+mebyE2hrN
JpAnxlngr8hUpVGPKbB3/PPsCT86UnWELN0Kp7ZBPIxmU/GXHyx7yIiAG67V
GWI6cMIotWp4lWb1LaBhJsDvnT1GjN03oVpH3ky/TZNYs9xxr5lFMif0ZPq9
e8bAPqDPz0SQwJ5cl3vHN4wZhXViil03sarjnjSgUbo+O/S4k8+CYOUa42NW
1syewDIHmLXbQVOd/b8PxgWWeTrP0KH+ps7jDWH7roOOgZlYwNZOdulkb2US
0RzSNbfTkcUWv2+9nPucx2YFzvVnyYqM2hrGcZ50QLgB26NN8AWi97Zrliff
X9M2pLJz7+MjFTdH8JhCKj+6/J5FbBrFyQLyZ0+zW2gXPSpNAkh/nDp6G8wD
huNw6+TzvqJ9D0BGoFP4J+4YJpzzZgcpHqVpvV27sMexIwIoUq8vLmnksAkU
MYX1FjssU76h6QVlIxLji1F9mYPj6iCj1lL96uWEYpyxx+IypUZByfk3KuWa
qTZ/RAH96RlbOXEOQ5CkVE31kNtNdjGYX/hzYoi7tImQjuVxFo4q08KjK0mi
nyVi4kAtWFU9XTssV8qz0SRJgqLKEpDZhk4Jyl/1eWuR650GKM1/96qCp5Z5
Zej2i8A9hf/vdndJnz6u3kOUEmc8Tm2JrAtPz/qT3UgD693qClT6KfEslhCX
chnILubt8iDzkhbel6FMNcq4wh87vuVn9/t8J2Mg3+F2qzcZiKXkA5/WIaD8
WdxPrFtRHYC9oygxocCNizSsFIRwF231iOlmghYTnOlZ7eR5gCwGGYRaHdpx
KCWI2X2YbogFdQBZZ+cfpCwzDFiBHC2JKbXtwBEPK2TFTpx3OwizHbPKioGY
em23I2Kofg5m6bsLHjQnNsMoBWJujFmfxefAnxFUR3vSaonBbrIkH7Q+CmXu
W/aVGXSqRt7aOpGUBDVbdsfwnCvwsU/nooNtsawo+KaR2kQi4Leaw+CAuKYb
Y4lslCMhUMuCdQo5Oz0hWVnJx1zDRhSeHgTYsFy5/Yn5gI5yr375z9qi74Zw
uBkHkfpmyMfGu2JhNzDJcAXuUDH00ODW3RlbAj8Bi5m1VtQhKiVhIiW9tMhR
q+cNjSF/agefYHjpE/eIoLXtlD/l0sfG+VyUlUdKM/y5en6HGIk1ehnVv4U/
QIHbHkL1RdRb2xEKYTmp0oOyZGykJRqJozhvxnFBV9X4GnrcwImjAIe7dxWL
eu2+ycTQcDqha1a+C7aHdVTprfbJhCbv1KbJF2SAaid81jwFBx9W7PeoWNcT
sbTUEFua8+gVKbwKTBGcJToTndVNK1V+pQENUMFtDMnuQt8icKJL23QNIJoX
4OAREy5vKs4/JVtWY4W4r1yVc9pY8U2w5HOgfVqJbrbLD23C9wdU71uHgYul
ePSRtv4QsEo445FCij71wAgFKD6Un/k5KUL1atEGhWZ7zzyYxImquCHmt6O3
at8GZnpzROqjAt5XMwOw6CsNjyoN0Pt4pD+EPPT6cSEf4/5DdF7UclSVDn1G
DNIWjTIVIlb9wbA8Je9m/I5zM+843h06wpHLaNLjv1ogMNu/dXs9twSkKfk+
ISpLgWwgC7FmNFGIXFOmiUHLdQ9XxuCN7phngU7Uto1wt/kmbnVr81SAfN3R
GxIWmpKfRwMl+VQnhzEN9t1BeZK+S2ufM9RVCBN8yfFpltCtuKyStTCpiWjN
zQQtX1jaDHl57y6AUOk58RaPszWFSGwAvdHjUVKcGn/8P1xAbfX8FzYy+Jto
xyqJyc+rlF3zVaP4/0oeVdQSq9yM+YAg69fIvKhiQCPDz0dIEDWELrTSyCkl
Mpq5uVExdk4lBiRdyH1wjkIqjweuEWPUs1VOD4B0/FPjUye5+t9pOVwsFVv3
V5esekgP29JD8wuKVubzUo1N0wkhUNZ5ImJO6MpnQhAiACdKpmkwpQHyGtkz
y7xondlgXr+Lgg+MxBbAy+Fm5wDbP0jthawTZV/T4rb9bF6dhR+sDYUWADDb
t2zXttoPpaP4YjZLKibNmd1GYhIO+k0Di5ux8kaqjeBeYpFj0u7X4qAwP0J5
ivMyMOCD5iRHZlm4w6fgFxXNDvcPu5YF2difP+OAsYGKtENG+nmTRx6ptYkf
7T6Ufj422JoIHOlZKUm79xA5DvseCBbFu0nW50Emw2mBBDlk2ZcM7X5EciaR
2mV6mHtdIn3c4mcwGc2UkI1vF/p/NC4v9jCrHqO85PuzW6c1KxfNoTftnE2v
BryRD6iciYYZOm6Ka4OdrXaVV1g6lNHOBPICM1pUHFKLT6DjJwvBa0sarKet
g1YZXNImrRmvPFO5doW+cCDIg9pva/ehda4qPHxcwD1tvtHCAtAi0TFyBzW1
fdhZL7rRJdknuGFR/eADjzRM+CFXFhIZq0XN5HM7Q8QLmB8l2XmDRvs3lF1/
gI1qXUCM6oAI8PLwNaAlyDxoFQE8UeCCswwlPJFlPGEFTBtXORSxrQPqAp+n
89ssIU7ljS9jgMecRtfGI1EaQSByvw1eO5hrIwfJISoi6cO/kaqI8uxcJmaL
4VQjC+gDwwHp0EsmFIpLaXqtckw2gENZ8m6HPeNftUGVX72pP3G8WutYeuEy
rI3V0hx3AZ7JeRfKoGrgHUE9DCNKZvOroXA/F+UClfDciMSpHpSSGB43SXWo
6ww7ygynN+aJ8v4uC/hS/roSdSIeuGzNw4cLSzusEragu8+HkNyFPtnkbaoR
Se7UNpn/rKo66rw+1JC30JDVvPp9BXNJnllsnCej0D7gOumw+TyuHo9fxgpr
O4h5oa5HsXZQ70A67uUElnzd+QXc+WG4yOycxsBVS2S7rkwWciEh47k32mpX
DLweC0YpWuQr+jK1ZNYdHFCc+6iI+1Zlr84bLDSdv9ZAwZCLHnOtexGnbOb+
DI9tfcsfbulsv1pbvyJ7qbA6X/LbYK6RepcGI3CJuI/sxr4nlmXv/yT/qHBo
2iS4P+IUaWIHaJRMIrv8J8k6ilfO+e5oQLsh7KESOWo08nAnAPP1U1MAk3rr
qXDgWeWo7WoVM3CylaaxxryZ+adSkws8ZugBOl/aZSsVpVq2GjnZJn9rw5W/
6A6i3pQARwSU5KemhA40P5KV6kAGLv+NHRJsxnFVToUlfkOqTzJU8/g/Tb+c
xgef+BF7JwvDK3i2/4duYBrxy95rR1MMlk+n6qgY/A9OfrHkwPscWh4FhUOF
JuUUDfMGva+CxMyO8e+4xbHcIpdcOXexODkKQ4oQVgNxrv1Xsaof8eMRH9Jr
XQmZUuJnOD6daobNL7xm7K+QSaekigcNC84Aix5F/QJ7a7S22xlIMS3/Es3i
o+9hzFrxo9oxy4FXdqgyZOHnnVNQrOJt7Q6GUTOvVDhP6rsLI2CxE4pSb6rv
jsyX1hpYJktu4jtQ/bEAwtacHHTuVXciITi13zcEYka+KCWTocg4IludGlER
ajtdvfeNd2ZyFEVWLa+fRwz/8IijJa5Ngei9zMzp3CAHTChkOglSxjWK7KQ6
pvL9/56wlJe6Hd/ynNH1JSdFczoLEAoAgJcSVCoe1aqF2hJCghvOyj4w+vDD
OrvkzrDEEiKc9sPOIJlkzEZHhd/rtmvpUmYBHQ3Ofeab0yA7ly4BUpI7dOgl
aLsyB1NpTp8B4Xfz9fymaOgBDOvKxvk74gLumVbJ65MCEbdXxbHmcJT87Wdb
73y3fF3IoAsq+T9JAwj9FPimJ379/LizRskId7dL20uYp+WH1N/j7ZSNLMxN
D/bgffov13yDhOwYEyqhN+1mgy7snWJJiVfYoL3hf6PwrXqbtzLhocZSgo1W
t9VqJFXPhO+2SKoKUluF35y0T9HDLt9jgpkO6JLBbsLfIcCV2JNfg82HPIiR
44P3AFt6pAiI8uMEQKWN8GSms+ILB2vbYEm44sCZZOOmgVmqrOUNa1AjxZqz
qLYoVONwrTuZqpU7JZsOQZ1LD9Lfm5GgDdY8hc5u2lpTJLSiJ92tEaQrM8Bo
+hH2WI/ARsHO0hilQV+8C518U6RwtS42wAgokoXpjt7U0cYETB1DmbiHxI8T
RzpYMGRR+4Ov5yoO9l/+IbKG5CjbfOWhhgYWtD6y1rsS0NARuaJjURH6HefQ
OCPYJqvXGBkb+sP0q7Yb6XV4nBWrLUwQdbeshtXLHZ9TY+PF9+eWs48m1nx1
qam1q+h9sBX1hTTbsIjEH08BT6726BWiq3+UOm6ZiovZi58sCcI25yTHv3EP
sK+R23HTJXRZJ9WBQg5+tJ8qyu5858fYrmJdg0X7vtvbC5TCc0PsGDhJ3fFL
9bjXwAmJBHU8QC1XE9Algg/tes+OvwF2kzYRg9AQjMufW5qZDRN/u2W+l7sR
lZNv0z0kAVDRN9pTHuthDOpB83WQJkjLW6Ihruel2Zx+2KUq/b/8f2/lBn3d
iHrfhPbaS0pwm3y5EdVsA9ADBeQwkO/zTVTMTEwbG0VPpocZorIEfBT9cC10
PIGV0CNblDPMiLG61ntglizuSdWlhDf+KYwgL+/fLopwjf7J5/S+7EaKOWTV
+opKsV9qTtQeYa/U2JUFNb2L5h1V3Ac9Q5JEn0a0IqiGcsbjNSPbNBmK2Xap
vkUuTO/y8bDgg9muAMSN9BRJKV/clZN/P3Z+wyXgzugIQ/GcKXaoTU9k5sOs
8DP1NPh3fHrCXQYp/2rK3cXl9foQgyTF73Otz3tZUU79AmTPIuQ08VlYbQWW
SYx1EAvfCNcMKNMREq55Zbgd9g8Mk8H4i/8QaVAM0Zn3vvwp8C420GcuW1Gn
TC1xzpclCscA/C3zJdGLF7Gbx0AE74XtmJWnZNxt8AOajYtXPfHHkmhnp/+x
AyRyySiADcfGVn+UYyiYa6b8EQR3MXpceqWim4fNRGYxKOjD2kqdBxEWMHaB
2TZjPxMjASOoWb1N0ViNQAivcMqU+m+GULus4s/G+AnOatqExl6LduqlMB1D
hspICXtYOc7UWdk1LY+czc/AA/hW5eQpyFVr5vuQ4Msf00YhswkkAoRciWbJ
FgLlLIR5H3ufoHCvGdf6eYvNJyTnYheyLnrRuemG2lxbUDZ/MgC3SDySZaMR
cvx5211fO/UwKJdfLl7b5/b6Ej84LGKcOK5mcAYcOuPyCD9Z6xK/qw3RDfkJ
Jkg7+T2oJZh/u9vcGM5cGO+IIs+4BLyLTqWwER8ehV5Is7bABJk8ZTNuk4oA
ELdCS1+qf8jLtS6S80mPVLkqiOPp3OPk7haSTRu5lHMribuaGkBv4h7OTzms
SFq33y0tbNQ3dyC7Lei5dRwUqLuobFzZortw637LmAMs/HpKhqrM60PTNKNF
OnA3ZSb+fn4OvRphAhocrMMc6x8tACOZgaLO5Q3JrAIx1K6TUdsVvWasZO22
vfEab81jOb7u/4R4yk1mtkrOCeue1g34XS2RQHf+Nomq5HQngozMKr1XRsUu
b1NbaRKK/bCyDyVGMk+1fAIfYi02ar2gVl/KKj9aHRwNzDYVw8+H/fRKlo4K
di8vYX/D1eKZ/3CMDcM8GIfgElLnHxrCpEbmmWPx2R52UkkS+tavI1YPzrmL
LfDBxkN3Bth6RC8BKxIIXNSMymlW7lLhj8/kdSFhl2YVbnXgntZY848zusP5
hkeRCHhRbLS7xw/ixtRI5aazYcJ9xUUx+SX2bf5yKVos0CPlLJxFVaQqiWvP
XJVWlaNLcgb2Ef4s2vWoXip36umgyJG9N2THt0w58Zzajh3gKkAxa7dLlJu4
3jRDVyIzx7i6315vRkI+scq7BzbS/KMSMo9m/pSVpERPyISg7t2KO37N7foj
zZ8aMZHW/+ojDdfycqYhyG9cBVV024YMOw5jTVZsgxvv5wPNRMC5qSBPX0Un
aNLo9M4+lEah35vgL0p5AIbg4O9rP6coawMMEt0144HORsUuXGujHas8hFKI
CXW6cAJrIDiqVjyU3k7WFRd2m4YaEujPumfV3rlLyRdb03FasxezubF46qBL
1rTLrezOl5mrKT5iN3TPxx6TYLgS1CpZPzIvI1VD2pyhvsGfdKHLh4SbP7+D
41G8hO1agiuWAvl5O/Ey8WuNAL80WSHHtpkU+XYFPY9NAIpGd4OLV3+ewtgW
LnBHWOawKLnF7BasYDL7N5nMNPd3s8NyXWvQWjd2Vzx0YVRA74JaxPpl2X3s
wnjk17IJWrmqGUPem+ZsfSm0n1RGeMeP5IsF1kt2+G44uw7YzIZHGCndjE3n
tuvwKJvcAN597MrrsYOFaCqBycGGlKn0sQsjZ2FY9mfDERcy0Gm2b7g3CYoS
HNq2whmriIAnzZ2fDPBwTy0KsXUEad0OuyiyKnYl53LQstZuN8nS3cVKzD7v
/8VjfuIY7f5iaxUzKLU+rG8BhvLPF/5EjIhZqGO0+7A4vS/zDyfNHenFU6lD
US5WLrn7dbikDQQ+2nPh1CxWD4Piuk+5qxvAQ+I0JuH3TvgxNxle9OhIZiky
BBB3VNWDUyXyCtwmGClAhfM8xQM0cYBzhQ/MKaX1NFjIkSOJqI7CnmJy9/4l
rfcSuXLMVthatAlMCVmwXwFgsLl/9iUUE/T9GE97vq/C//THLULfx2jwTUHz
anLX2AJg4/1NRC+7vT/futosyJva4w6RfuOCoKF2Ioto22RLOnX2Zd7AXEyp
b6JyLrzWmlSvJe95zb+wF/1LszZ4DLcyuSJdfGH7NauLj/lYsskYyJBdtBIz
PhnupwSpX78A+NbnhHZg43ZDJ1LNmbRCNtj3Ikvfjhnf0jY5er/98eWLvvyC
Pr3+8VYMMGDD1mEhKl+IqbYkcyzPIj8yJ7Cv8zvAZJfbNc5AqsBkb2hTDZpk
OjfzuPa2B4e4zYBnqILDHghXpXHcplKGoH4JQHNR6ctKn8tPL4qTQMKOnmO5
PyeY6w+GBWpBsj6f16z7xcQ25oZk498UP+CVj97YxBrQkm4NK24h4YpwojcQ
ftjZFpuLp4D7Oktgq7CBhiFd85zw9inQM3yym6+lnqbUWZsH43ddTrZZccAt
j7M4N4RMDvojpybcUgqdIscahLSOdQgO3qd8OWtjEQLK1jLd3R+OdRmQX1ot
07EjrEuesMOFu1h20kT/YIiUWSXKBp2SfvIPgM9XiPuA0NVdXTd336QHpX74
GKjjPNcEERzjrB5s08/i/1vNqtcECiWIKb9S5hwyT4n0A6s+J8KPjZiUIpgE
zUrP8A0dU1Od9iLSxqlsUwACWEg41N6xEY2sbgwlZRxlSYJ/0RC4X9bqj2GF
GR75GgmDF/TyCQi6gSzqRm5ezmHCTtyKoyYLlFrG1j1WAQxgSe3OAiyShkRz
OHeYuaKL5YxVWVSIcWEecLu5HTbJqj7oLlTqqw3V+u8Dfx+BDjSDr8Qwz+ay
w4YMlDhHo6OBNFOwsIDuCMFd13WD+UKqtvpFYczxOH3kZ5AZQTcqqpl8AqcW
wNOX0SeyLFMUxLT9bG3QopVUbx+Lds4kSjiyFQ+LcOWnQoGreI0gfZKtpCRW
1wFZJK6EilpyKm0JfRKTnuWvDe8+PjSOndmuiu6R9PeNYoJdkgJO7P919koe
MyJPTxAjecDc2O223jdCgODTIhe9zekqWt7vdaEHut7Nxd2XJU35hRpU2aAC
NNv3498RupIlRcnQarAYBHb+kOELFNpq3g8ULS7t+A+DQbspxBKCiaBkgC1q
4Uc3NzcMsGku3naGDs6akhb++yEfzQOnztnQYXyEPKayrVdiSucSmVK2oYl8
pyRbuA6AiTohHz19LmR4ueIV022so3ra1K+rbGbfFym62Y8pnfEusdvOZFY0
dhKVT2/KPTb6uKsY25rUu12Au/PHweC2h2mlgxHS+ddW+ye3qbLm30AnNVVl
gY6ylYQn0vIJz4k6HoT4pLg52JLdUWVVsSYLUVQNFM5fs+u7CqYQNFlufmDi
g31ILJAiFokpywQTb+aYvpgQOH/r5F4kC1zY4i0C1RLN0GOyoZ7zJ1OZRuYb
jxmFRJYkUBZ2cUAMGDiejSpUZ4UtXQVqiqUHh3qtKg06ixCAiybjPDFEO7uD
MIekulZ/rbSyE6WutYuduKkvtKZetiRT8KhghqZptCEb1DHVIAkq4fHhdz13
RxO7p7w+x09N5kWZHrOqavRZ+Pcx0Ebk1pBhpojUhzPUFOC1A07szDZ7qveU
/tHe9zxexhRiE4mFX9FwZkUYYvKBe3ixxUApaSghwRsWN1LQDVaV4VSDimvK
YA05TCkmgQ7WLgmKeDZlbJwEoFsgiUkodLK15P9TSg/EFiaBsGHj+pNFCKCN
dXBMVb6E7uA3FcA2p6og+0+uynn7Zn3GEAyGnnSvi43J0FuIDBi2CffuHO2v
jzyti2TKgBcLGKBjmm8drCRPvqjHBy2ewy9z9jaE9MK42AyEU9lHWptEuHEb
md6kgXGmR3OqsvRR0C5xD1JQlwmXBP5kFzjZlGfbjqbpscUOCJn9HLM2vlOo
KB/Z1YsKSKKn5Sntd+aYSteHI2Q4oMKBQs4+/rS2iws7jn2Ju7Y2i5AUwKz6
fI0tY05SbMHJxfB4p6NyhrPDQJnwJrfwQZfjAcRYz12p65bL3xPNMG8NmD8Q
75BDkANatlSH/pz078HU/xVLAkMXX5RR2nnTp9wtpr0r4DLzwT3pRROEiQFS
/lyvfhorAEo74lEnFAWz0WgV6/4AdMxUxDZLogNnzCmIkJuj6n6PJre0Gn6A
HuwxeyWGzOETfu8KluOsTBliobWlnLqODLUnEiisIJttdIjahGNINxMNM33E
SYeqFuvEuT6t+063Dx5gFM6/u2tSyO0pyZp8XendYsTAg8tjSsdZqNwcjMFG
usHCfNTeRgA9ymTK9V4tOHVeK3EoQNsnq3OBjrz3q0SGHhj2IbTTlrQ5WvaO
zlVZZ4lNwIl2d6wM2A/QBBXUSHRE2uYPVAmmle/xT2/wydDl1YiAkNeW3c5f
g3yfbhZpiAqI4RZ/VjfliwnWjMT35bkDDUcWZRKw8ZLlm8L3Q7STX+56ZgYU
MyuApKu1Gqe/EEIeXgr0BpwMxGo7Mpzdo50c0kFWAsNK1iCZ5o3yCpFHMEmu
ID+dB0anSqPvyKIw6ccXsaaliaxaEbgtJc+FuBAdm17BcMgUMME1yE+bNk2+
A/kaMoe1S9d6XBSirxeXfeZe9u4A2MYLDKNL8ubQT1cJTnBoHbIjzIc63eXR
4+IUjnzsENAWvaxO+tgWRAJHPnhtGBhp

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyK7N2hEILVk6YuiEiiApcfGwP0x/P9dU/ocHcAoZfW81Exg18/aZCycE9mjdlHPfcYIz6Rn0cSCQCWcf4z3VBZOEJB3rhLYYDMEtWwhwwZRIRDR5TcaD2EY+pwiMB9gVyIzlwiz31WJ6F4EI8s7VJHrZQ7XyeFp0jPO5wVfpvgROPbRyNznCL9mhJsOojh8C7tvi6Wnx872gVCMXc7pDXqvxXpZEKa70vCWTQk3Wmjgh1SRKDrwln4alipm8xiDDJQ9LDXg3YhAO5Ev1DCcezJjBJWivX6gFwf1DUjsXy5zaXdbD86J/peCxKSYmD5OxgCpj+AjvexOBW/FxnlqCdNjpSgiZqIcF0sbWC83ZP4uhIpe8xZ+aOkqYc2Xgfi0EHYX0jzGcqViM5pO6HFlw6zDmH18Ffutl/vlQ3GYFvdRPuM3b6i7Jpw4D9+nGktFCzZEmbTVFS5Iq539/XO1iQCL9Ph/IvLTSpUquuU6l0evLmA1Nx5psEzKah8q27c5Lg4eN92Rvbhl26U8hYDzeZVx4IBUrjoM1rC+JjFlQAGYYbnVJLN2X0O5GPXOZhzaUkGTSGmgGtXElEYltDUHqrxpyYJJegr+U36Ltsv06pTfzctakwOAfOASRI24FZYaZXfsGYDjkGcRq/9RB/5hQA6yqswNy5O78YH5LDOZqsIHtHGHcnSMkCHQR3trebTxrdgsbPBXz3Fx791zenigSZsAOvDTLNVGwJLOHZJ5Z3FVe1YxlA9QHNdSCK463izMNRSCa9bXsz+Xzs+2vGigp/My"
`endif