// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mUKz8HRmo393n58OyK/BP6E1t9BWsgSgZzrIkZMMlPWjlAaob6K1qLJUoUG6
cC8T4Ja5/xmwA+JM8zIff4MaQRt90docpCjLMXPVxxDbuFQXIL1/MoVB44op
H9oJFizFlu9OWYHuRMNTDmKn60XCVIv/Wgo1RJ3kZ419Q79EHdt5ZMJnTrit
CiOe6eVAX0BajSviIUUpvkEaCW9GmURWPB42zvZzuoXUaxgD0fFYOVObIF3Z
7DpC808+0tauKS7Ei0qStW867Pk0w4NVGt0QAsVbwj5rBj15gUxErSfoTfDo
/XjZe1/ekZwOHIFr2DQEunYIGWhyoaf40B7M/Mq0+A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jDKwLMD60GZgRoUMwbysV4jRBo6XoEof4aT8ggdVcRMr4awa44LQmf7CFgVS
M+21iOWHkIEd769tFil3ubfbn/ZeDTZO2yHABychzbB19tXZXdGpP+gvLKHT
OqqJg6dnBSVnMF3ZOGR0YrzAV1OWVkKqZcFqpOrjGSbZnfkA6UyEewlFP9d9
i+OC8uFSRQsC1FNXcKP/jFAF2fG738t6mClI5ikIid1nq7ZxpR15ipitnx74
2rEy0uqwDWcgp1LcDT8EDpoQ9PizazUGEqWu+MWl+FiH6W6Ph29eQEpFNalX
07F7pcAex293IQHZMvu+EQDYqNigGseKOKsuVF8ckQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JKUGQG2NvugRw1pxBbABWQhbY6o1XJm82BYYA1+Ym7t50/1MbVyx6fb+BBlt
KmDTE/kWJL56NCNMYaICuWxJyzk+s8E37f9fXq2f+kbwpD+51baMnhdpjkPs
fO8rrH/xX1YQVcrc3P70++LiJBqtyP+U4xXj8dVoqfegJJt5dPjfpFJpiGaD
T9iy766e2ESjNjQxThwEWGRFDQ6NJ+V5K+Fw5k4ANhLONl+4KRQ+N0/4kY4f
jxR3VngXwYH18Bin+YuKEpu1NGavXHGnSOC/5bJCPYJa7BajtT8OIPJfSJI1
Bu2HjmaWbjZblprS7tZaYJJlFU+x2bDvRwWyNH7lOw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RHD1BMsfAPBg3weZi7Z7ZpeB9RAVTA3x9kuZJSl0EfVGTY7igyimsWSRXahW
Gfff2I27fq7now8Cz8DAdOkfr6yjor5CfZuaIK88V49lWs8R4ih1jjXRPxj+
9ir6v/L4ct01UbRdAyYWNXSRSc1FJv2eHO1qhbbRB2VKiepgZRKiB1E7xL9+
iRJL3beCUTBZ3U7ZZIMWreDe12wvZyBl6S+Ehj1ABQvEezO0hVDor3EqNrC3
9PvNHHsNFxoPstOgoRv1U+dGzlrY/xmifH4QLB//Cie4sHvzbiDiaLHe5aGr
6FPwiVU50jUFQ+bYA+nujF2O50kqM82VaZGJBCbLxw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YqTfLS0AMQ5NYNWjhWKaYEczwVolqLWIj1j8yApdNsjGeDnbLy857G4rpLwg
pLzjGOdBKfzjwqzu8ADqF3rIR87F2g1DkPQjdu5BMjxiaw/gWtqRs9c4NsF2
QOXUd+HlJJm1cjwAnf1TncnMgDKTuoIqGuTYsQZ5ImFT7+xO3qg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
wvtPc0ovogmVCW37e0eMKiFRk2sqDuotxMbskDebhTG2iJdYidYawwcUYoP6
396c5FwhOUt0/LWxT7H41Jo6LF8i9hSZ7e3jdcMw1g9ISjpDuHtgLlVltvb+
Zi796n4e3zbwB8wyJpYUNzJ54V0fjX1Pl7zHh7Pvo/i80SJBoGl7WtjL7uAi
oV/+zpmJqmwzziDm2i+ptCOlVdPOuFzTVN5z1YuvUdocrIx+b49UDZ5J0Klw
2oDe/jsLkcVDm1V2vIrW+i6x7EIdnopY35zrpwuWDiIWSoskPE+e7QDsdURu
EJOj2M85OPX4LazwEe6kExH639FStoTzA8ZxJlKeJVn9yMpGBBeaX0X0btv1
/rocMGUFKL1FuBBIVCulVfnXjaNcFp24XqjyrFX//loookT6eouG5SE7Ant7
rdSIKderytYgcHiDETQFfzj7MYMKSlS0RQ9YAb9bZXH0WbqywFeEewdNeGNG
prlukrq5g1VLTSqL9Pge4ITAK3GU1NA8


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Do7RA2PThOdQINxhTDLxZT42WMkeEpW0/J0D5vn95XQDwm/oX6d4LzqHFs4A
3kRhECc5bdIrhOiNJ65LJrrwMHCG3bEgcecDOWni9OS+4Pbtjj/ydjB5nxuW
kfuVmGMAJMikpwMTQEGs3SoW0ddf6WohrOpKGj0fZlp+XE/9RHo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
O7RkLjf9NRXL68C4tMnWWVEWkO5XHxTqt/3jODF4ndTbOlgda/eKcfqCB1II
NiCtT6G6f3tDsKC7Dp/TdlgdF5F5Um7xIykNUIjepiLNHxz6ncSG+MV7Gxln
aK0ZZX2DyfH2VdK7XaM5OKVWTeFv3WTAL6RZy/zTuTdtj9D9ldY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9616)
`pragma protect data_block
aqqFBzA1P8+tIjJ8wH3qoXqsbmAQxXBKfCmw1rryR44zsrglpPJQwm6SH4oQ
e4sDG8ooRXBMBpzgdk8hVlxI/cy0lATOC0MpyeQk0Q2oIcS+wNSW5FZ4x9+l
WaGu2VHUULreXrmd4IAEDzS/jJG9PpkHpxXHNV7rseP4EaKFAEALID49ETUV
dWft3roZe+eaRMFetIM3xGBVrGOAfNeCHflUwT24Hp0DR4jwumHZYES9qMzy
IBA/CgXf8t7+AbuKbS6iYVrEsy7mS05YYgOht+ptjyTW13E7oTNgludByg3S
Dj9kVx0OqXirH2O33br+P+UveeqbsCQQOdFPGjlcdAmcQzrctsKwH286r1Nh
5GGI6k4FSDaeHzBfpr8KQr4WYV9BdgQxPx3UCNrzTieslkc8Jit130tQ4ygi
JNFIsvrWCEvhQBezp+IRhbyuq9z6FdONDMJX9f2tIxcLf7VV+8nGDb04SYhf
GrKMwEU5cmRJrBgRBYwbMxLlHU5g2kLqnd2v3+rVpNDyzPLpc3195Zu/3dyV
D+Y49aOwLy5LyAgQq6Ifk4SM0cVI/c6Jfk49aeUa3XAPMwXXUF+82X/8ixJA
1lfsSvuB9iZfdVUScurXDJn7P3BrqMlWZaFrhM7lnYidFrjpMUWIBAV59e7A
E5H+wDplNw3azG+SoMi7ra3RDhthlfyMIH/qypdvF06yyhb+d4h+uNb5SfNl
PttU2Av+FwyHdo3KKGOR1lyUkPWGoZ2t7R/K35JecIdiHGLrPzPS9nwrw4El
kth8aegyM55dzs4gKkwaIagFdfjXZFChOD+lVWhuL3hKJvLcvXV7MDwVVODH
GmtArSRgKI0SMOaKTdtcl6+ILgpRe2f1VL5O+LFGcDW2qtdniv96Ff0vihkk
iagfjUbIsn38+dHeh+DqQ1sMsXVF0fJCtoD+PyzFqmTzPuavaucv3m5VVBNf
DRMuvEfvXCb7IRgHtB8vKphpED/d/V5J4c7WGh3kuaLRcXWdOQpEqDtCksJ1
4DWoITRqGkG9Qs2OVDfmqrOfoK7QleAAS5PVNtbhJ/hlUtn2AUDRNX7bMjxo
yUDUqQu1/PsDyGoi+BzHc5SZeiMChiRKr2XUXHKBtIH8t5/N9Q0EUH6Hi6hE
77J/WcpcGNC2CssGylxEaMOYr9BoH5AP2PJVvEgAe6gN5A62w5vVILIpLaF5
+smtR/DuNeEBXE38r31nEvpCYguS6eQpw9v3zNv4WDGjb1L2A0w937N1fHmM
NFchq+ZxJeelo8t6TjBI41RruKeFnyTpuHPgBMazdzdmYnGi0G0Tff3251Ij
jGioxOqvl2nZNScVMdAofbc1+XvmSlItZ4AwDJKu/1UAtMpk5n8zPM3tHyef
uGYPukaBxWuT05TDF1TPE5Td+UZMGXeCW6o7y+m1kbubtNxvk1isyy0wXeP1
ikPsCtr2OYZAiMGY5cP9gAgxFsiRhrHeWjJAtqBDnVz6G9pwZubvwhChdNaz
pd3xE8e08nmt0oHcqqkKgbOkJbWIDdJu7tKvUh1hmkNn/lfXkQj2kJ+vzTfM
jVmKZSbCIRW5W280QNXeX0irr2IOyNbl0Hxmg1qV+GHiHhcs3zED3Y2nKXRz
GbeFsoNR25PSq0R/J/1ASMDQ4Oxu2Gm81ivo6ITJI+kjxBm9GibWK1YBNkH4
tLbuduEcz25QnsauyOAFa1wcH9U9vORSWVXJ0iYXcQnntRJbPoMcZcOP5ioC
RPlFRJOzyGqAVFmUqOqBH9RvEgcc1RZyFjoJogLmZN1cOiqs7uWRFicpgI5l
ndlqt0snF3KpJe4CYa2h/ZBRP0YHc32ZawI1IA7Qku79DzhEaeCo1HbnXjnZ
oni0UBjDPtGR6evsG1gdEostyLpAv/5YAJ48/ANNJlmJjM2OiqceUbC6KPcS
M8PKuzDN11tNKUzV88ampYJrjamRgw0uKrFN+hhGpZjnoBJwpqIV45O8v5DZ
U282Yv6bxo9dMkYwEcT2A02U8foT6rgQIARXf1YjTWjuMYIA2cJIwU7KR6MU
N9GENQ0hxOsJ3ZE8/Fxel2W1TqK0lOmP9q3mx5Nq6jTz3mO2HGqdaxsRFBes
03b/N3k40g7xN9XyqNG4iMiwx8mv5GmYLUuh7EGD5Mc7XnPHwohJVFw9VPyd
EOGDwH6QsIlbQx9/BFOYKDESvYGN5Pd9vGdvmC/6iG2E9Ni1NJBU896XLG8g
9M0rkuIuMUJJOQ5pQ17vURDIa8V4uDBJOK3juTynFj5Sf0iAjMrneVXQ9jw+
61O8GU2txh4wo3rdy0mmWZTetp0d3lNbJZrRscvMpPCN+y7P9m8lV6duf3I4
U+K8qBB341/6cnFKYAbnT9bAB8A7kQ0rMpb8aRn5o66nQ8hW32wwBftNgEaH
Ep+jEdnKrZ9yAbDejIDn72Pi8HG369gLKVCMXLux3sx3OOBqelbmp6vXTv1l
nvNUQe0VnBeIs6Mv6ZEPy+oZX9j1gkPZInDlnTKzIedwbKJP8WL9pJ2vqWCX
zHHEuD/QNpKuDtkfMZIvjJ0jSKuVMvEDfGlEBYsjqw42CcKS+lVz5+aEsQl0
cWpQMGeS425yzYeUzB7aafS+xFL7SJBDHj44KTU6dYwOCazMwzLOQ+CDf6cQ
OwfnguBRgaOzZ8EVZHw0jG15kx6vApXlifiNpiQJIrYuvGrNTrq6IZglMQMR
ZmEle3tc2lrZvXoZ1MmrVtEaAwotqwfmPA4aWIcehPAa7dvsG2EKKdZ5C7yz
6PGzc4b25ePm+3E8hbxFJ5ABo3YT9YWA2oC1WhNeM1LALolbnU3bGZWjsLer
MciEo8/ppLF3RHTkiBbwuRmAqiDuDaJp3149IoRDy1oBapMGv1S3auvzFRw4
T2gBMC3jldMo/BXfO54XYnaoRet76XUFRbs3vOTUSMHXZo4KpgHK22LL2zxr
ZJn+8q+Kuo82Xq5oi/7DSOBxF8qTout0SSFubfn0XcvnEOR/K8u8ZSoYdDgw
7hjwk7vem4GYnmqPn08hODcwA0AU4KEyrV+pjbOIUp5fQ8jxl96sAZ64Lpx5
BFfL6i5bTFf5bgBKhlATYxs5evZSVGaQcJDEDyhGo5NBikc9/wuLseURXyc9
Y6vwgHq3zCUSvyL8bG0TNxj2FPV52PecUUXzv0oPn90IjICCCdpQtqv55q4l
HDSzVH7JU4+Zi464X836fxhxtGwNziotPE/l1rA3U3apKbtO3kugs3KZkA2p
z2PM6NX+T20EGan3LoERazrHy0fKuJ9rueiDZqlpQmpREZ0v/MPtdFs4wDZM
r3oRDWYHn9uOnyupg9zAzJj8thcM0x1baNCbkTLU6915GNqo8QzM+WD1n6kv
foqTuYiAlgl+bwHszRrc4olccwWkCa2RL/kfqVYgBYSMnzJkuYXxyBhW1u+h
YqPrRR8DsvLGPaXqJgwIPHlV2I8CHlWWyZoQVZAr8fxVq+/Zqf7/Em0+nh0S
7qn7ZZ/9nzGgwYeevjd7ad+XOiBGx8tB3xGom69F3n+wAmI+qcnj0kmxEU0U
mAnNWcel1cHUPM/NbMUEyphgHanjffMqSdIec9o9eNCLgFOp3jUZ8ptP3B6R
Y+F30VHCnci06YsGmjn0L9YjsDmz9M+ZiegZeRvu+FW2kiNdEpYoPui0Fk+5
BGzFJ/8uEQQmMHq8zw+vOMb+Vr3i63z4Mz/F3kxJwwpvZVJDCk4r48iq8B34
LFsPtoEUfwGJlk4b7+BB8kQl/j4BZxjWsUnVN942+RypDi2it4Jl3LMbyMXk
kSYpYBk4ymJRGwDxmmhMv0Ct0TaEPCEZ4Qce22sWSMux0/xvBZ0tJD0xfWd5
0wEMEgJj2Ep/7aUeBazNM5dv07+6BouKUJlQNCj0xYVtbz2Q0iij8/WGGpp4
Anmbqw+ZnXAbUA63IeWH0aBqkeClxQLTqn0ybUz468/sMb5ZVFWbNq5I9DP+
VESaGn4j+7KeND+jGDDg8jArOZ5vzsCsIDRfxcgMZlXuqVecSPqD8PWFXAd3
I3OOvb5Up13CTR89Xedwk2iNyjnw6cn37KYMyUBduYYD0AcL+RAcupKkAzAZ
pC3oIT0drUQP7yuFD44BFEnC3GL9UutoeTHExJ3ERRbKqXNiLqVxBdnr+79G
V+ZxCeKswzykaVnAVVm4AfbJa+29MIvJjwdmIILsC4z8tAe9RFD+3TyvUPOR
WqDmEAQp4vMgx2K1GFQQaos2hvnHAGlIqa2BJ5lwDZJlCzWp1Yciv9SujWje
AnXgkvDSplsQy4fd05pN28UL2hAh95ZG8E3oVqG5qcaf16YJWq0IrzWGMHh8
BmJ9GY+Mjzic5C0WZZhPy04Hsh/BiRHNYvMjWsYZzlb4/Wvu0zG2cTf2iSaY
du88OEBy/cVUT4CUPLnsX6wPqMyR3+WCIiVLXk4AXssmSN+v+qzeQUdeGhHl
gK/JwO7facLObkz4bL3QGQN7UFkFOwz8YSBVhlFf7Hwg0+wrq7kzl6tO623B
in3vMJ8s+81tlEswhS2EpuJx6gJT4GDo5DOf/w5H1Gus5vgpMKKgC+wPSmvB
qtlBojYfJAmDC3/LxkCkNZw1cUQ0khhMI/kRVLJwLbcO2bR80eK2VhAbnAfF
cZ1vShDYC9Ca1J9c6QxqZKn5xRkQmJd/FVyS55yp372G9fLjOwumxWTsih+7
enyRPn6jZp9pKbr4npnEcMJxY7pOBGOo+Ja1yRRTKYQRXQaDBf7NavBe3f4I
1XZl0TOsskf0o3WQuvCescmmHS1J09HIS2rtyO0m1a4HKpTNwsMC4JlZI5UU
uiHVz4dkVLxyTGmqoDjpA8129q7MicpCV7ZfNB+lBGso3VQS4PRNI6Z3RVmK
KhRwy09TwS/vJeC3VA8UpJYIslPJTtPmw6pg8ajuzf5XcIA5NajjYmzwyPF6
iiL0wkWHSul4ApqlIFHIlg589mCQ9V1e44Rj+3g2mwXZqJjN5gsxSKkm44Ej
znHNqkQD5Tp18L++Kqjn7z66xr0SzREUyoCr2t9afHOIypTlN7TtcWbPa2kr
V8akHTWS/BxGWcrYEZl1wg6Y/AlqFLGjI+mF75BlgdlYpXdia35ZWMnHUTNV
AIP5icS7s9lyFNh95WD7X1jBoKTqhSPV4ndNiABEDMoIXiPaCU8cIVjpiTrK
/Xw7lVopPjCQoIwv9Mmw+rWmslVmKYl3gTZpdwOiesn4ANkpyoI/ZNo46NsQ
I78HtRpyZOcTmhNi5cElfcY9palKmpg8ufUHkkGh2mmbbuhSzQwoRkgNNla+
ydfvdfj4sHMcAjOicZAz4nMtUia8PxrJkfKbktyPtvGarjO4JOKHvmUWjguD
g8dPILteRBjNLLtTtI0dmXxs1I+YHae84kC2qfN1GWNa/5ibzGh2ZpybqFTc
mzttR7ad5sUzi47m7V4YGvFzSjPJyb1PX9dRrKCdQslYr388QbvN6xBYW7Z7
vQqSV7SnfEtFfnMAq8LpV0LtKCzLOBV4157m62ONZjw9Umos7JtmP2lj1Ijy
9VRBvLRCHfGrjHh7jFTZRQ9micMSr9h9ZSqMr3nHa+uAknn6qu1rE7kF9/Mz
sqf/A5zwVU3CHFlRCqywsJjqMjhztJoHV1gbMg/kRtIIY08rdqzdrywUeMxU
wVPJdnmvouTz72nEVNh3lnpaGCWPhx1iuwvaMZWvdpSeOmZ3lfrNJt1hf57Z
CBKjD1ww8dd4loneyYVWBmDja7LVTJNaSXQv8KuW4b/Ooa1Jpx5AGJEfL9tJ
BkzQeOnKW6uXVf7D5Uy+MRJylDO9zvSOgFBoID9D4DLJ70Tq7QwLWaAGALvN
CIMJOD7WqLy9cezCxzW8clEnufXETsphER6NaQV2cV6dcMSRnxrdk/csY0+Q
4I7dNjYjeaCDryCGhMypOta9d2dcEMwErkCJyzn+leVT5G+zoo42vN8Qe2mj
l/UF6sCDnCIcp0knDgQgAQwsG8y90oeFOHSXgVRb4UxtMxN1fB7ILwDSD8/4
3xYvmuADX34YWWXE0dtjUTqrdDHlMWFtj+L9aZBUfLHTJ7R4+oh0UImFaUfG
DeJN87xldmrPEuhCaGIdi8ou0gSOMxCzKDYGUXsFDsjtXEqoyn1Ver8y0miA
ss4brWuC7dQ3PR4UzfhYDHwOhf/BFIpkHQCigIW59SqlWMAFSJ/jdKsWRdE2
9q3mF1o+kr15QvJWF5LC2Up+zvswzj4LMLb+kLGDTa6yVYG2m65VpYaPpvsp
PCf/TD7dKpDeHrQPdQYe/IGb/OkIayy4U9aBxy5N9yu8wjLSE/m8oZmDp8ps
L3JIs/zpZItdrUS7/Ncm829NV96Ztt8rFuwNHuJEbTGIKW1D7kFvf/wQmAXZ
MDfK8Hpnay8W5qrqA2C4ZbGdS+m8MT837vYsR9jOU6UQ5RD/djwLwc791u1Q
kHTbnVoOM+7mD7WeqAHNyFFZjswOJ/+G87LeVPHJGw94EnXdUD5CM5AhMG5w
+Dx98s0BIT0BNmNifQS3p/3bVISspX86bgDZYrQOQtI0U/wIsvdu7TSVYZsW
p80n6932WCR0xWzMEzWdtT8QdlEs9okFVrUXtDaNbS0Pfcdo3avGLhIlOtPl
IwIOalCmlV276XYeRs/6FPPZFpvW1gjdmql+IoQqpj0tH3lWVAYmWMaMdreN
ycm1oT2XSlZRofm0D9M8hdR2siO9Cquc/qegqJmlJdawn/VuNLl6JmHAdnat
ZJGD2CAffhBPklVfac0C/yImlyoAFJdLzmdlxvtiXIVVI9q3yhuPrsrSD9Dn
X5imkqS8NJOHEPW/6qirnnYZTgGdsWJJEwHO4HsUG2Ekdpr1Ndi8oF8VMrtT
zL/71TLHvfIPLVoWSOQ8/+DEng5Robbynpnn4ZxHd0NRfmmdNVNEdbV18It0
E5APrGphQlXYNjs1//h9/NIpnFpeRXd/Mko0+noGA8DFAUImB/r3cq/X3R9L
R4rz9aCV6gkq6uFc+Xjr4vrKi0Wqjo7ZiHt2o/60E/lkf81oCoBq6gR4mlB7
3DwNko2vsFfpel33ImHHrKzkY0pFuDUMLl1HXRbvxJZCtCxisfUphYuL1GSC
ZeugbqpzFGmJiqWyD3KTCYIs+1H0gfa0p1eJ/uVkQdsBd9uprBamv6iOm/e8
OXlkaLwyeK9CZFTkvzwQ4DdPgxkcAHp61eJd/WyuRchjJSbHzm8HVFe5TJq9
3+ulhGheu8mY59D6rpIKG5fMme/KQfixTe6TQzVga9AzcHzRCzYkcJOQREE5
TFnxfao9q++6nRvbQ/XnsMKV64H9mk4o3ywvxmG+70uDFzLtwQkWOhwEs7q4
G7UCyddfBuh+u3F9JW4K+qT+EdQP62iqpfNEAJp9GeZShVb/DjbAh9PTNaWu
ygXizbSjxFPsffYkDphM+HLfX5Ht7wFiroxJM6urU4B6keVw/ZjZUdQlLg5s
okWn8R/TiOD5Z69LJGEk53Aoqg9eF8ju06tsrIXDKJ+wji0xIet+YCEGwfkF
s8sgK03RdM02OfbTQrFeJep7n7lqV5vNHf0McbRKEIbXt/cwk+Rm2kVa9yw/
By3oMWH52u1JvG/rByhRsuRXQZImrB+Qcos+DNEP+9jedQ7CowQHeiSuI/di
iektX5J9KSt8NDaJ6bS7IK3QFylYZ2EpUkl1H2qOvhQscrPTsI5BQnqqyFvm
m2yJZujZpeXzeKP7UCcNxw8mwZJ095ZyYfFMsgFTF08idQNsoQQVxogiwOZw
DmBYzAKXcTPR2P8b4AcPeaFZa0USnI1W11QfDp68D4e+PlturLf4Ss4O3xRN
cz3UpI4q8d+S+zmojeCdY5b6j6Pu/AbAzMQ1GeGcO+yhKoYhG3MRHPbz8Fgc
mIax7E4eIO/mVgv8lkVxuumvk1vNnq3CW+ENPByDpcXSub3gfrqR4VrZSRI4
uxxb3H9H2uqPiQJLoOioPRLpQZLp7jHLr2y8NHvlcigmphW8XjlPUYRRQe40
9/IyM+0mzqjheswQTg5IgEIgOniqz1rUsKdhWGhXfl3U9Q7pt1jhxvG3Smm7
8mc9hvbb6obi9yzCZkqdjZWCgYkHqSZGz2LpE1RMY/SF0y5FMC2OotZKJ6Vc
splARPpXG+wQ9mLNjdr8bTexpAl8NL0u5Gx/0E91lmzUijfkVCyh7Fl/EMdm
OuiDnT+TL2PYwx9eY9XuM9p5NxQiZszn72mgXQzf7XQZOOK6+ieNE4BRg2v0
s5/7Y4SnMm2KHtmBLmItED5HDu4OAge5NnUj9u/f6fo7hoxEe/9L6tN6fb7H
ZP+fWsnHwGK8L879UbT+QLjOgzFEKkheP0pdJCnsn3ICo3i5BerIlg1Mx0E3
Ic1tr3RGtLkWxbr7WEqgN8i/r7BQzdT7Vzr8Y6jcJKnLeaQsUfpfNfbwfend
ei8VBoGRGaDWNz65Nq+oxKs+bGzPMmQ6L/HiABdQSpiBaR3W7aO784kUplGa
FAy/oFrMhGieN8tghwbnu+9S5Fy/WvZ4h4MTGLxGd+Uu9eQt36gwrksvwATB
xEhnQagN/STkG3/uF7x8+ujR+OVW08pc5tDnOY/BGrJZW8GYs1OOy3azoA17
kbJQr/t5CKAjjLS4R2Ww6PDGPDCb3PRvS23YOon0T004py5eVKhcG4vLh/R5
cY+TMRYhCbSmv8YLFninnQ+F4iIotU2Xnf7ViT5QcKEz+p33sy3nHxBnx/QA
ogrdmBV3XMDfZ2IXU72hZ9R+YlsomGzHmVW8UDGn4/BuhG7I9CRU682VNDsx
RtLEvnzhnWuSjmbyQ3dxc1956yrE0C/AExU/LsPicxJoBbWkmGtMcddG1ME1
af/sOs3+kTTJeW54zsrBN3aKS622xppcNsAcBb61TtMBXeTyWf4vA8X1IZTE
yqNsvHtw0alHNw8dJB/UhLmq9dvv/EhVldFgS4q4ySKXi9sIfBep91RzCXUS
svXyUdhiscu450Ugwcd4N3g8waaKrL06HRtpECZHk8Wl/nPftcB/5V7bVMM+
0IitML8taa4UJ2KmZ32zKXfrc/KukrDb2npgYa+RFTNYzY3Fpqal8VQY08pg
UG+bfS7a3Hap11U/qMNed4iS6YTvqsL9UuKEz/yS5ln6ZM4dQXG2/X3OWU+u
bX5U9GHFKIcDlABv0A1E8Qldo/kRk+g5FN0YlU6j0bHX4h+D2g4OMP4rWgC4
vEWYzrv45Zd4Wsri7GEnUgdH6e+MEnPGuf7796kY/eY4l3Kn/KfVIdwziYCE
HIedFL0LgDTbch33LA/mpJDQJocrVv5q29A5xH0h1xscXSCxWGDEKodHD9c/
6RkivX90W2emMl4N8jjA1g2Y5FB5duECcL/jRYrQYqcQnkAe/dyFpJvzyCK9
T/q3CiqdHyxl/GJFDEeb03rtJkKck3SZECy4sDmPCQnHRL1o49D0pafwvlVi
fMZMSVIEuVXJyGTZ+wsNDJedQBZ7PbY9lPrwRRGp7OtZxORwXc3N6L352Btw
CkGhjxRi39n16dFMFy3xN5QGRvyn2Foc5ZlzUVJjkU0jFb2TrmmKa1vMPLLt
r/EzvEACjWxGWq5vv9Y0Hb2V9lIVDuDQRdRtSJOXETc5nuWBqaGdLwY1Cv23
+FxuQAbPzjfJfjXHa2nPxmS2vqOiNVwhpVI/o5jSUlQ3FDnSV3HqMT/hUHd1
11VQWtIsSk3vNM6gWPtpqIFL2JNv5MDjc4p37dGo9EWQE4FI+zml5vkkYeQ/
YgF6AhbQ1CuHlFspPJCvIcBsVT9XAiOLO2vsKF+6ZX5N3QnGtVSj0OIdCqEy
F72KToQSxPIMjHghChUXQTWPGOhng5Uy0ePZuN9bDEHcBmBQPdvoHylI95+X
jzfRMHqCGFJNkA6qBc9Fz6CyIm6A0kDjwtMjJk8ACpa9gSXXPSmIoG+I0+f7
3zUNQi6yAn4E6c9Me50Z0Ul5VAJmTjbCcFjXkKIqNC4Lqn/nJT7WnUbm0RaG
k1lq4qikcu6fHjXfh8hczriQISKCHv5CbhMx6dexE8DZk8FS7yx+wkrSo/O1
kO2cHrPh1URD20v1ZiU+C9w0BHZdKXOcXW53IaN96M63RRfFh3dvpm+xLgNb
/30LTwOWRbUeNZ4cKJ4nTq0WoBys/Wd4hucZh4XKHZOR7sfPcIJ0fJgrQMzH
NPTDt9l1/04WrH/1PPSOsGqErtKJ/lYAyBT1ARFRvm9od/jsHOPcN0Fk2mkO
A8Du1Nli+QvcqBnVxL+5gtzXmRMRFQQzoiXco/Bm4+gba/ENUxGgpQzLeVlI
s1NPV3TL8BowckgFDBF/OOIl1SmHuWrExmGik13sk1HXJGHUsbazj+/2fWQe
JAdd9EdWJiDSb7UYHWXdQM/RqRnS3tNLgECbxdkCbXm7CmyUbNWWV1mDn7yb
K4e7PeU7j0TTFG5b42nr2PSBT44cDwNAobeYeGXbEz2armNt8eGu3kpz+PfB
7vqzQ2QjFvRuZl8s0gCzWlCTcS6uSGYNNMCGquq1Br0FkRB8sKAe6BM3AQbC
CWrsvJJwmRgGzi2v5qA1KWUFwsf0q0q5TlCtE86VkVZyEVuk27Z4wh7GGWvT
fUtpdntC53vI4vYFCGrAQS6E169+1DqCvYB3YuuZIfh3ZpdGEs9HtwASxFcn
zeeKwNoMTO8NhkqwuRj3rqDkLLGdb22xu8qLikSMorRwVNmcgbEtI2bigLQ6
bXflXYGW28S/VB5r5Y0V6ePmIExwwfUr1Q10+z3aAcpfR7rtWvb3l69+65vi
jLQdjmt3ZzaX+3yeB9iNM9t45CbimlLBHX/pfaV2IMI2cNpxyDzWC3KY845x
ie2K13C2Mw9Ln/hlcLIqqY605XImDj4HLoAtQD67SfXcCljFdB40Z3zKxeUH
yfR9pT3Pi1UJWqDxRQ4ItHRCKN+AkCAlUUm0rWFMiULCCFUsPB5cQFei3gEE
JS4h7B8LihrjCTpEnF2nuzb6NXnQX2ABiE++/mMylqkuxBxYdtPEyfi5vOZi
ev2m1o+w8WWoRoO7EjTCvjMxgu8qC+ZF1W06yjRsO7t/4q3977mSOTNMcOIl
4J20QQotT44H9oELHqRx0L+41VraINTHODPEDjiBwoKFuBSI5wMFfjk4H1tb
i20NI1beC+81fw7+50wIyytqrKHyBEbnu5JPpxQkWXCJi7K/ODWSEfBYW4v9
Z/JE6DTpmGs3w22GmmjyyWPHnGVxwy7imOB2+qtYhg7iMJKmmfYtpppszUo9
Kyi9omJanjXaFbL2aa4XFKeW+Ms2YYwm6gLm/HzabgYXWlgovP7pfL2AG1E0
6IPT8oN5ZrMfIBgc8kSFxCsvmEt6VAerm1qrjSdc5EhLUR6WAxrFIbU2nQ4h
soK9ymDv33Ru4t7JKSJ5dH6DoHYTGKhWKSFwm5n/kXzudZXVH/y7m1mNQ3Ud
ScYVqCr7lEwYWQxuIAzj7zjierowtNU0f+r8cLm9kidfgtaPaI3REV49H2iD
DH3M9cZeBV9yl2TYrarD+gyicHTsWcyZUfPzx11TJ4GnVSDtg9UU5clwxDxj
7CyEG8wSQ0+Mle6HGS9vipXlrThdyhkcI7b7GW/sXfsfuSh1K2ymPD4/WM6n
7jlmUn1FtrQVZiqEkT1Rk8QW4rdNrjwCNKH4oJ/b2OdYIdLy74TAzyh2BINE
yT0aWhopd1FE9GsrEYrfL9zsO7tNk5EkSP9Nc3/9pEEvGxgQ8p/NiMFAaYSY
ITatVDbbTSIw5ckHT6G52BveWgS14H6zs3ky0VZUkEssJ8uGPDqJqVB6YDCi
9Axl36YAmc/c8Ax6w53EJHj6gd4IljWq80Xu/0Ar0vxlNDZQ0jyXh8XFYC0p
wZZEZsls1m6XywmMO4blcQgAqc/xDjjVXW8aKSjsc6McWsDJY0Ixtq2z+XA6
vYHQTyOrRx/rsrEEb8nEwaKX/nsZb3UYQZOpRFED1iTDnmXipZoYjU9kUB7X
xZg1W0LxSWuJkKDhrSD3K1OHt1r6S1hMU+e8kUB/j/0X/h4/hAMaqqY7MqsG
yS3ZTO57zcvxwcCKvmHeyvgu7jHWnf4sbnDqyiaDmf+Yuc4GQ3drW/g/reqp
8QxhQ9DT8/HzGpcZ250gfA2eMUuKCOwUhHRJmC4majlBn85Xe/okrus2CmFF
ztt2YTswqKdjwfzSAqjzN3mLoF8L49r8xfWbpp7FHT2Ns44ieQrz4Sz1IsKo
CytlxQfTp8W0RZI2wy6th3yJ3WszNN8wvjHs8yjaPpkrI3Xy53A6bJ43h2Rj
h2eBA6QXAUQbxIaVY8TtlRTMG9eL9zyfeYln5b1+LCXOHTzR3UL0G/4epecq
DCcFBJd+sCIjrfeS8rgBu6FBbFmY70eg0gk3rT6FNdyW2PVv8R2fFFOPMROX
eIKlnU5FWXsYn2UPzzie3ixOn2v7fLexidSXwamzy5OD5nvA5rVFGC7EGWwN
R++eaFI7Cq8et+KX+DcLRIrzn5Xpb6m9cLhtQuLryGEUz2WlprsiBF7xv7Ni
ARI4CdMglyKTurPf4B9EzbKinOGp1z/WuoiyXrYX2cXBZmc0pIwp3RJdNtke
di+UJTtvxG0KWiii7rWZFYxdAX/RjGp343JaSorPgCxOlTm3v8tVXvNszs5w
YWL//KVubwHzO1oiAZHG/+R7OomqyCeVzcLH4oKVmohgd9NLUMY5QvAS8GwW
R+iqWWW7edIWKb2WtFMObqosdxziy+QILRZQ8Mbu/dN8sE4DVHTYWDye4ml8
T11/k4wsR7SuMIEzFP1Ubw6NqCvki+a9LQTWyI4KF3RVAMUd+D/kVTzqg/I6
VO/wXuE3M6RXgxqD82ZvS+58kvSzd0+5oPxlnss5aw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "B40jvh7ud/ahkCWXo8CJP0S9JYnc5+J2pwOdONjrEnmjRzb1YpxBEP/gM90XdEQFf8e+9j+GJABVN1VA/EUgHmy986oXHU6n9uJJjaeBsR8h22iSaiy//95eH4kKFakRZgkZDqWp0dX7AUTwRg4vZKk0rom9cx0xsiuc1Ki6fTzxDmmuuNW+yyxk/luKJogixDl7f05H1PhFx3JTfD9y6cRFGovJ+RtyYHOBbLpk0wiu05wYKdmOMraJa/IX7Ry8eHXlSdqNm8MFKP4rxFPEijT2WQU3epYu9V/AsIDJtcxQzWf3F+6DLIUfNk1xdiOwVY8gYU4HTmqAjqHoxn6Fo3TBPrMDZ5X4RHWNu30L8GuDiRVtbSZEXBWzUVFai/f8yM0My3TJFZNGlwyc9qsDjl5ZMPy3NANSnPhfCm5upThfT12dzkZkiKbKT5ogX8ExqSzp67TA5jEI/D/TGG2Z3x6Z7XEnR4bBjSCRkxvGijxZJWfJvJS1jl6cObkV/eURYScSYYcIMOQNN76lpN2ilxlOh5ptMNNio7f9uOetNvmJu44uBgsLUfuVO/H8oR82N1NqaiIMk4ihp7uz8bmOfAeWK968s8WukPuLryu2kwiZtSaFVfZCoBsZ9t1j3fQyTYZZ6G1uK3PIu+xd4h5aKZbrbsFMnymTbbmfUZkdbcakzJpZk+7MeVgoWyZF+Q1dmdCx7ybWEtGgRFUyBfvw4b32DQ/WLIo97HNJgxzlksHTpICN9nNJAZK4+mO1rTSxo/oC13npd6mpEweEljsE08hnAsnWWCkk3Qq9MqXwnQPvI0f3EQF/oO7xlMBOKNOJIVVUh6In0mlU9r5r74ElDYOrnpcaIxHnvEpNJShaJDDakgauiw3Tr6poHVgjEoY7f36BNzIitOgLgFuV7mmQy8SCM+63t7ROR2zHytvcxM8ZJhy+yt4f25aXr0AlRrK17mnJfts0a3Puw6MQfLUJ2XJ2H5HIExlVOJ8RJDdeKhVcpGsOveP2p9MLR6LLG3n2"
`endif