// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
m2sMpnzdmS25kx59ZyKWLyd9j5N6krkmbIY8wCj/03wzTOOF6Vtbk9t2MpU9
wWW3QdlgF3LaNIdyLvLZKDBRWVCpxs1woyfIrCd4YKYHjim9JUb6jB1pgjZI
Cfb9/dPfOt1nVUwGmRP/CYLpMFw8MzX7kHnic4tWrEh7XWP9KVlSsDLcTyqR
+5wDJPNNwfsBbd/rC1G6M/QDcG5vcuhWfchBpdBcGAT8DEX43NmSnIHDlQ9x
MOJlbDnPb6fIPFEKgxQ7yiarh/lrN902V8U2nM80scE8RwZRm0f4kzdoQ7F4
zBLc4y6dP/qLNsGDQOLZLGpyekoK8vDgoOzW4Y4lsQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
g1L3oO0BdlLec2jDw59ruKaSmiCCFAeMr+vYjNu48zJAZgCNlO1+t2+F0AAv
0hID78jm7OZq6rmcM96OuhZeGrJ9nYsIEGTfDilVnDTIuG6rloZSE/ZT4eps
mq1JsKYfKbz77BurHB3rgcU3Dpz8ajZjH2Fg+dLIeJW5rIvMOqC5+teKABQo
y5/T8ocxZT905ABaw7g5NeIk1y1aXXE/uQbqzMu6J6PS0w0yKXL+93l+CtkC
Ix/A3cqJl1gK3CQRQrcZnJqwGS00MPPc3yOblOB5CU+UN6GRLxT8VuZo6BkQ
jGmnOXg+uj1zJVSYaPB+4AWtHEAytrorSPDxGqlriQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SoDZ5QMVEfDJC9t3u3eiv8BjDYAZZLXeAssg2GLja/nPsYtQ4j4LCh11Ukwn
XgGiZjBRIQuTOEWEIn8HwTpzJvPb2nOXa0qLpkxKrw6bPCwbYkNaxoaZhj5b
N1hpsOYN9jptc8MbrILDd3lEsyhAf2I/9aIJ0C2/Xv7GeijhWxHa8uYs8S0T
5TruiMl3KEFmFgQiOF9ZJwtfzYtGAXeu1xBaesEtO8ubK1HIaRJmy/8+YMSG
TbYtDjZpWmh0egQtjmqxo8ZoSKvDm/kp9fFXzaxwA387Vnn0bQDyfUPIKqok
6yo/e2cDp01H6bflY8o0EliQnJEYMosiO8acHY0uXA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GJNouT9umrQ5xivKe5L7EpuJ+q4+qgzIsMJo+Vab8VGk8GMETOlhwnMYSseG
6qWYvZaE9PKaLu5nLtdJzgzJatnfzbK62MMvVAav3aSp8+rR3usztY1Engnh
8jAiNmq3oVsEmSOQwj1yVQ+VqmjJft9GcHIJmd4+D2cVsDukbMKLZYHLrpfd
OX436VGiwz3dqk49mB3snmjTgbOQSKyGumW/uzIXtkygvo86t0FTQtk7Al7X
3v+BKTtGD+cgpQQAKQGDIto1s2qV4eaTIFalf854X6N8MpW0JQT8hM+02NeK
MWfFUT5MyQJn1ZRaFWPAGV5OHq2zrkVNq6RjyEo4MQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nVq/EZ3u+XhJljgIys8BKgk+Kudbev4twJ1Ia/YKJTRzUGQGdCtiYj1OTOem
7hCfDbesMFOtFGTL1iOGYvCMsJX9HelTxOLKdzeIpusQ8UIeMRwPenYy/Xdz
NVNdNPA97mRFBQ0iSHIVQnfxJe+tVuEFLehGZAhrr9ofuy4lo/M=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
q4O5RsTo6exQSEIn9gYcvpAsNmxZC4rTL5mB5+cGJgTMqTbJivHX8XszhJUX
mrJMApAGb+D30V84eZwklAQmI1Zw1219atErcSs6Ob7y27O7u+ZeWvMm3jWp
n8S1DteOpBhm+F6elEE6gki2jPz0NB82DabJZNg+cuKPLc4YqBjPS523/NxY
bMuhi4T1wI06JS89C2N484cuc0Iz/tcwvq3pRFv1HJzpAN8pB270hDHoVAgU
UxMM15wKbc7W/4pv5k47URILmXjlVai/Y6nq/Nz7RoXj2Y1P+Fwxjl+pCRes
dFwpGkbAEMn6KUKKMXza5gW6xz+WWaU/Yn8JFKq9LhOpOz1lbp+BQejUyanC
zWCFYxzlNAzuRnPIt5BdfYcLux7gWZcneDXpmu3ndrchFlEoXqMF39tIHjfr
euOm/il5n1shiJ0ZLrFc9FYe+aRljYnBQNl/DhZ1ZTAY/STET341EStzt7MR
OrTyBHONIpOejS+kAyODf+74uux+hcjU


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EDhoIUzQBCVyziQvBy3PqTPGWpZNbXcUSKy39DwOmBy9llBO3v2vvGxhJYB0
jiWv8om83u6PxNIKk8N/hCQOL+DFptKMksT4o5sT/UENIG3DfLCNFIBufTek
kV3laKMMuKn24F+Awh1vYKl4gcqSETtvJ8BeZDAYmdkHJFC6Uao=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
WyQ8s2nbSUaY0pnZXX0KwllvwqXCjvoFjcqcIaRHSj1QqCkFk7mZfl04PJUs
ijanrizJTDogU3Dw6jNsgxPKcpH/9NQ58pV/3aha9KeA1jx5A6zqYQ7s6Gxn
mVIztLXTHs29T8E2GHzwV7fVVCyeaR5ist95PsLaQ0Q3LYgk2aM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 37152)
`pragma protect data_block
UrM3mHfkMAphIXv0+jvkJaHYEHdSkn6GkcznZqHw14m1T3v+k8UL3S4qvCZC
0O5J5GoGy2Ybo0tnZ7F78RoWEutsDKj2s3IiFZM5bO0WEkyqhkKOvdf7slY+
qtv2MkUV8vbFLYf/ZFFRmzerUPo+T5Q3NbMBsHdUbklFnDyozWCOorX9Mi0w
1nGCblGN8XNaP/etG7J030466saNGdwH9LPB6QveFwzte6TDjAEgTZnc1J4X
q64gELccBsFWd7m2fIQXHpDuAaHpf5IRbbeYK/D6z1OzSywMj0xj3l8MUpuT
z4o/Q/QVVdDI2pHtIR3YQMCwnI4jhOVre9Gi+117ZbZOF1GBhcoHwURt+4ME
aWiH7HljiqWO1vLJoJ6MQ2lMvACN1qfD0vVp+YNf0Hiy2EHhBkqnEm3BsrCg
Cm/PpXa2ZYtvayL1qowzH/Gn6QY4rme8pukYtsrDXHdHnosDJu6FvDdT3U+Y
GtQgE8EOGE504g+xkKgH57w1JKteJdg0LJeDuXHbVd1YK6AhrUNDXmrLfhS0
vvCBXaDdTmvEN/+QWiIi3uCJt1V5S3p97qJomBaRfhV2yc2YA8vR25suZSAZ
V7hgX8vUdxKnv6C6oB30lsFRTm0V44KIO1LZoa7hn6qV86SgFioVSl2ICNaG
lAACsEwYbwIBwIMuzKqjouHYKqAFSxxvuaJsEUWpH5Q3UKdFIG4kz4XZL52v
Tq11pJ5xI7jsRilPidgU/XE2bAq69pVwjlZ68yfTfvC6DQIP+eYXdCiG78UC
Zdl8c6JSTpUrjqPym1fJPzSvECnHlexh8t8pKPfM15Rm8UptB1aFzPJyyO66
prV1GXA0NB7pcfyDD2+CCVgHk4eXJGlbhLWpT63nTTO8qToL5NgxI9Y610yu
29itWxnXEETn8wG8GIxz5UM/JWuYou30gvjYwy9mJF1PwQAPzRiQXm/jQCrA
rgd84Kqi2/+6FqTX1qHmew0a9Zc61sEtN2LmT3NwvrZCOycvpmYrAGVZHFwu
bWjJUmReaoMOaYzd6xmWj7TQYxGen5q2OEW6Yiqn/j7JOqq+cLsN1kxZ79cO
vSWr/gUidRMg7RC+FblUzMgRoVywGrzWobxintAfYzmJPztaGkHY6EaZthq0
ZEH2ldWkkGEpQ9VieC9skRfxuQZ3Tx8ZVlUVhz6Y6UoOl/k7DrHqyISD8qKz
m4sfpVXPT/tBM7SjG2tJ6psy7opMaILW1RRDJQIE/alu+py89RRzu1D0dyyL
qpZsrauOqulKuGhYkDcVqdTXpz6rhCa50k1+ilKV7KWbzg8+YQ8dLYutXcY8
wpDmOdPRjQOQu9317ri2jzcQUTBWad6H6gayO3kPEuidrFqzT5MwmqE4hwwt
dsUbYIwncZkv2Vn6KZcft3Ch966Stz89m9XiUrqk5wFZpI71Ee+XkF76JIyv
L/qGqyLnSFd1ijRV78bNFbKR5aksN7k9fUg4Wmdx44opNDXzH+bVjXCsy3VB
Tj7wrJoUVhIOLJzOhOx9S7CJsAsIbo0yzSaCLTSbCtvN5F9y1z9poPOA+kXl
O7HU2ACDTfy26FuvJc39yPGbYZJp83xVezHVlyUoctoVgWqpL9vTHpg+eozX
7BRgyaex7RMaTIllh1bY4orHDYhYlQ7nW1P6NvxElmn5ZZ7I3A0/NQ9srFoC
QE9TKhqAUgY1c4qn0IFnIayP3qQ4oiOtaPn7YSsX61WC9+KIMF0aB6aM7tL4
9IMs6YjEga6C2glj3XdzBAfHrcpELWYbTvVT767ullqp1TUMRwPcGUm+rsh2
Q99izdHQTz4unwKxrQ0sP7yVVeILPJuPsdzeOWYDJErr9AA93bg5p+YrFWDT
roUfCkq6ybt4K/nJL4JpJGSzS0GVEyn5zprzDX4dGbhecobYXKFqxQXj2Ied
v6zafh/vzocrrpHqzCvonltPpCpK6b7X5rEg9OKtzZB41AJo03Vzo4fAeNLu
cR7Tr9dlqu6bpJUAMVKgs/tl9W/4iDYrXmn1NtKvmRNnMdbIQOa9rKvInHen
QU7OE7XC9SokXGkt/l+7Yw1HnjaqS0nuD0KOf/OpJjoM0hYjwYJM9WGNXQiX
iaEdaFa6Uoy1IjKUdjEezR90b+mTXK/f++XXFI0MdKLayaRnJZf5RvJg5CLo
l7F1SozYGoLqkprBpwtJVKkbk+qWuXQ5jWMiu2EsUPfZRaVSuWNKHnQG1Dmo
s2Dt73qDDaeamyS8MvlEiCeCMbPO6+XSr6G8UvZpFsCxZiqvJ6thpUmeo3RJ
vXVwspATqrLPVDsCK2HJTu7O2QkrWiFFZOmYSqIzv+93aCUIqOqw/Mk/sK/e
kPRsijfPlwid6YbJ5uNHr/MHJOL3UUemxucUB/3ZMEg8tjBGYernBQ4CpY09
osuvR0hBUNHLr2GMVhNwSWNX9M4pXC+fRje/K0Z550MB0iXb6EcFli7ZDVqj
mEHnsWEI4O3g70+vrn4ZqXytVPIKqkY3kU33q1epXpxPGohtgzdFacYT30cj
K/RCIeJeBt8kLurGnYwPgoKUe5/3KUBVVp1PJWWSquDLI5g+AUaSINbiO2Bz
jj+ZW/EhWIJpB44AyWUN6JpDxp7zJLqhfxH4hbuiiX+VuqCedakJG8N6QKnT
cGG40hQGYdrJaSo7FBWa3i+xEXvBDXq7vgLpRdyMgBiuSgfIMdbsS1mFm1P+
mpb7lTY0RjWaeQfhtlRgTKXdWPjpJJZMp8/dxXgEMtRPuFixfypAJWp4stbt
hV0uMY7aUqnMTxjgNx6aqgqd7a+/sg+7XwRqiuTMywOrwcZQMtQycKNo7DfP
aOwQrOYQcJCV06xvrkirBYj4V2PNqAOEeLTXYHubjjOWc80qx4eSF3tpXWii
7DuCUA+cFNGYlWMoF1AGF0LOt5kcPFLNi1DH1s+B1m1YqGErVXEz+Z0es+cQ
/QvtnFvTtVYGI40FiWS/VnltGCYcoxlsVxS19Zz5+sF+NNFUtfM+aOUaGxr/
qLe2ByWj62EAt83d4q+Oku0qkmIhZIf3RZ1tx1XHDhnWVDhiAQgVmYUZW+yD
enZD3mdV9bFVV5MXdMyqqd1fUDeyxxsscO5KcMrIM1JDN+WuMvmd4QwplbJB
2Bk8/MFVXJpym+4OcFhOAi2RtmyIVOcPXUWu2vYFaOe8pBPXRatg/PdFnm0L
Yxucuc8y3vMvQRDxxYDDMRrKtr4vy7l0+gmwgAuj9gL9EXtzgJ7IL6mz7Iqe
b47/IpJtwlVyahSpWJbo+DouecAaKOhiGRlAZCq2LQWzfm3hsq/FRcIlKM42
6gdU3HmL9nqWXSyHvz39dLSP3tLPBPH06592P+2cdYfnIah0wkIj1NKM91e1
gM0oH1faefL+lVSe0T2rvL6U0dWCcxKkL3d6t3/0Sg7cpVhp8zIKqKGYRE44
HWgm2zsv184mhgb9c4oHw19xG6xSHQ+u7PPOKvZA194p05MBOTwAUfJLlPuj
+PRGTMrUIYToMK3vzgpMbdiRfuuW00rS4ndw3TBQoz2aDkrsOjjgpO37bCnx
BDTSEX/6uGbTdabvp1jSWcmpIw9rmSDNpw3nGmzLdvSlVoYM7aZ6+EUVn6K4
4djGqLeQcOyeH52vg2q3hK8bpcOguptZOWCp6y0BpNBIn86I1WfC7xRSfIQu
PCHcQUbLmoj1kIoDeCVeb7xpmUU+0jNQtE+yoFD5mFapXUWLAXPF3MgCfq4m
KMXs28F9Zuy5kisJZWfhKl8K0zPw4+ejHHW4RyV5o9RAQ81hfL0/ThCcwmsi
bOuQfbjR3qB/Qcjl/c6v16RzBSReBRH0jKHINMH+pNRVXDSJrxAY8B4rvTjQ
WiU/bUv/SwACif/R498TbMN45sXAZdswlf1iK1j0ofjk6xiHCOKRMB2f+/fs
6vauHidBCs1xEpumxgdBrAPkKchDtRNLGA1q5/FXojMvJSG7Tru4c/IHYJHH
O6hT4eoTEdveRSbJsCIq0nBk5ZvVS1OGsB0O2wYW3l+CihjCr7Esi6+t54wT
P9PbjLc65h0CwtIV11MPU0BkVOe4E4BlOe2GtfCz5M+cZ3aQXhvPQ9+hoyrm
sqHUqTV1IqIlGAT7NJrHRv6whN1Uv5e+X1hKNfYVcKCF8SypaqHm2PVzE5kD
4Y6Xn2vsoMFAmwC0XETeqlodklPuus0Y/7qOkyVIK2oFQiXcSDa/qRHjiLER
ep58nMmir7nVpODbxHBPOslFa+JP0sED637Hb9y3x1Tvjycy39pH8O1j9EA5
Qk6xXGZGQ8S33EH5d3nSabLbVPfjs1QWly9qxJuy+3UsOAEcAnWv5lV2wv+G
/CAIRjx0tuTIRipM0vYpfPQkHUJYAj3DfWSmE8IxxuuH2K/rsbe/V1bLZsGN
WWG6xNFChhvD9cui4SaBaajSvbOoZr1LmtArBEQ5FHeNHKSpFu+QZomJ7bS/
AYxz2cM4+9bpX3zy8csd7YP5mkw8Qra2zDa8qCFy/dsdW30SO0xl5jTdES6M
Lr/rzzDG3oUIAxbWOJ4lCCvqbIAs0QGuRymWePx2kMYDPipLr8pifGHqMbx2
h209yHT0Z+zRysBiziW5QDfecduURABXC6NPRs1GtpvccHL7ZvyWGsVf92Wl
A5Mn7OnaRIybm8ZYkX5pHTcKNKoFxTpQK1wIEtAmeynwdpEarPANWd+r23Mu
4OWHMSHF2HnoG2Uy3hoZ19mlGl5busGjf7sabz6QQzmwIFWyp8eGZxMuk9GJ
7DxdSJup4Q4Z3SpRU2G4UJCFzZ8P7Ty3tY7WyIR15230s3836v7K4R3l5M8Z
wu4Bh/LL0Bov/gFLi6MDA8OBZB7b3ZkmL33wLnCpR5o6qz52KR5+YC12Ohi0
ut05dXzrY3Jw2MVL2Sw7dPcFLTD+mhA84HCqiW7G0O1L03As7koYrG8zn8Yj
KybHlh13hfeBwoyFzviu/42H8B+uejAp3iCd15kEokHArgdaN2FiBEYAesGn
dB1vmJaxDGeE6vKCAwuBMVmYiql4p060YLocwl6Vr7QVMQfbB8rdEjeWb4zh
59CjVJKKAubochkmeXI1/CeHoN/4vmUdEEJ6C7DxwyiEuAEzcdEtch+wruGE
ufDcEzYPZAWkaXhiy0An8Ng/8qLCctU/SOuTKe9FdGt8oqiT/EQBCn894J3R
qfk/mPqF4abtqm7aQlNx9wJ7Ai6PXRLxgR3Kckhlri9fSUv+HlbldK6K+3hL
3T15J5dLN7nkv5QdduKh1kVnwaixbtHCxOa8kTJxi2XKfVDS/nse8eCGgGAq
szP4mlo/g2oZLsUeauaUxvqcQ5fu4sVZ6WGG5LqMVl3EZQRE/7kjrnWp72nd
auXDrxdGnqUILtMjCt8efawdA1Ap+bpja/MpeK6rQA14/gPrKerVnXWGGnR0
9Qyh/DnP/ldDt5wdUdS4HpPY2LHQ2wtwEYu7BkjGRxrBKYiVbKQaQgMScXFA
bK20Cojkv46RAtVD8ZMlFZQZhZuHs1rd6TneU7uT5anR2wpmIYELnEbNyZnz
KWx/FTdxQI2m0H2o2fUQZvKL9HZjZMswLefvncL8VJGnDOD6pQx2tjOv85ws
/qDPeCjUrFwD3oyQ3tt+NC7JcWnusTTNuRqnL+dIII5tJZcCEhGIq055tiA6
CHbdKg9vF52cpq2iTPhN9Vj16+OG+FepNiIRuNXv9YYJQRuXF5GNj98bpUBp
owdqf8e3R93E6k0aZitFJo15pFJaAcsqnctekdaR0qcCT7/vs0bH6pVVzorp
Fb+ey6O/O4me75Eq58vTRJrNmX/KrAq+sRjv1lcpdVFPv9vDJhuiZxUnVkTQ
FunF2CyNaaTwolAWENx945PW7m4QbC942L5/A4YBuuNZfDQqwWqpVvJmQMS8
VdSgXPs4/G69DaUaWC4+uX3EGSDWjJtQAhaCkeyZ7+L+szvgbMvitjOpgVjp
ueK9mgYXbklEb7I1h008u9ZGDEIYVZU+ZxvhIpCkrBww8PqQqZTs7TWRU8TJ
6h54Q/C6cRXbqmweJE5cHkY9MXZErudlW5DsTEmQ0E5SpbqZnHmLxOGglOUZ
8TOAiA2pwKIdATxmkr2k12OjS72UaBNVzqy3ZF+q1+En1VflViWS2sA7Dse1
H8ujEZ5NSoE5t9/LoGtYuoGDx97r6zGx3A4PNT0TykGmwVRC4AKBgBA5mRml
hOOiaNl/2PE0h9XWEMMCPM2G57tJTe/yIBAOC6YXAjyfZRx+WI+LlUEPw9sS
zMCiD+A3SET/ISxeu05dkdORbVBGlYeoE5i0EweiiULHD/Pk3dlMqfui18z5
6mrZ3SY7NGl1FINxLw9qFpZkPXK9MmPpSU/4Ibw+/lRPmZSjGw8C0LfZwsmK
dSFp3yqwW/GndPBlVIb4tqzjAn8QSrlOHKx9AdtHGWxG8sxFlvDvqznFoteP
crmFLzFU+gWOI31qVpfy7jtNTSNP+h6ngMLmb0VB1CLQ/Q5RMi1Ffw/vfpAF
pZAJg6Ib/LW/jU6EW4tsdDvxaiPS88QZ89xTbWQFAnZxLO37+FRpBstfGmds
CwOLyfWA3v4st3YeB36OzRBfKNfNSCLDVAKuu7OKwHusuoMEDFbmIzMKjAwe
FKxQxCCNn2qC/vN7IvIUVtElZfCZdPqXQL+LhpgYMqkcSKnYXXknDSeaL4Kk
VFnxmPqnJTZyjjHWamL8c1uvZwoU+/6tvhzNAH1OaUFYviV0DzPOGQKuaiu0
RIOlJaQ0/FeMnxsqgEUhst2qLV40FizOO255e/QB1HlTCJNA5dCABg9CwTMm
jFnA9WE3Uk8tnn40q4UfQAXvx5JUsqxmPOQp/vvP3Z++LVrSneRBq6AGckJL
JZCSbx1Z9XDlwdX29cuxtDqXxDOTqPCIWrw9XclvX7XwS9ghNbkznlbfT9gV
iTobSZP45nXxdO8wt79DwsCri6D17YojaaRt6BLNXQLnE+vGqOTHs51ppqLw
VdZWbID55+Kwr0MrxZXQ0JlM7ZN5Z4hLGD5ztMwEykxPxOuTcp26jMSC4BSO
dlmI65PgcY/dmxNa7lTeB1ldYbPft16iJ/lcaCLveogK7/FmaQCWOGpGM5E4
4L3QXwMWHem4rZRHBYE1IBVwoOVgVVW8K/x6ENqsCqK+utEPHYw6jj20o4RU
Ks5qBEmSgdVfa6W6rCgbeeeo+dY8mR6ZWbV22F2EFgqOitI8rGm/jqybUZAp
ynsGqqlosmT9cptLoa02QOFSl3NibxohBjoWqu7GzA2wartFmHHtqxxCIeSX
7jZTzPWYeiY206GGGKKnlJ6hbCM2d2rLgPA1GnaRg7Su7uYw2CKtyQRoQXzq
/7jDyROlH/cF0lKWU4FKmWsjyV/Q3Hzo173au36ygwYxgTkVk77zWSjnCmfW
7ooXArj3ee8ZBfUMB9xGhg3Vi9H7D8IYBmJJDZ83zFrVxu941w6gWK1LpbkL
JWVUcSkvxYKVZ4NZ1Jh2fmeDhm31a2bepFh7jHOp+/XNOPjRbetd9Usjt65l
2RlAbd2S2yQk9krIXM2RuYQ9YbcWYDmFbc+Rb/hAiyyFfWpCVvyV3zj6bd0A
m7cFr69+6nD7OrwcZeSteweWkTdxB9hetD5LEbZqV4v9mXRMQDV92iPutJD4
zEeNYmyKI38J0+yxeu6I9nDtiWQg3+MfzF3QpOsRWgHhoixbmzI4ECcSLV3R
MfIdkR6M4YV1OMHX26sj04nIYGXLo5ilXfmZB+fzSdWjTjbjB1rRNbaPCbZJ
8ohqM9m9Vwc0y35Ov9ydPgEETNFdxcCjvo8LsV2snls+Bu8r2OpgwOWV4nAo
kcvqAbPTungBnkTmml5GbuYECQA3EOWGf4NgiaPDln6PHWs19CkXOVUl7w6y
cEiORqFVJpzARkjnhqA2z+v4v0KcuM5M/1D+ECsX5YecbKhkD/JMp3jSz6zs
sByRW6+rpUiHWhc1g7RAhwI7cArsKtxeSzZxO+Vjaxioly43NyZ4TkIF3JZG
pup4Dk9WSJAyg8yhdEu/pZ1Bud5QAvvloxO+8l7iXfQzmkS+TfNH5sUpD9re
9yI/PZfqME4c4lBBFItiHpR5MYeYuWbV4B6gIOLOkCA/j2hAxPHn1pvq3d5k
JK+HdS2KpgAUAoc8KdrjC6hK4Lhtt70mqeqSfzrX8o+QcxbgQ5Ua58geDaT8
qO1oshdDn/4L3d9dl6QKmrydaQks6CCSZKSqbNnCMYOzIy6dFz0o9yducRuj
VipT6ovz9Kbt38GFCDbB5ghaCNZ0quvay/r4848aU7EY+aYNSlSn0lvCM9mj
U1CONfc+tXT5y7cBB7h7PpEQULA8zlfnlyUrkS8hxwilzowRPOidBb7tJMPb
yC18bQcro76XdPRL5XeW6Vg7xhOmVmz7DBrF+J2dslj4/sHTatsVAENXNz75
NSBH1r9Ty4utDyi0DTN+67B7g1oID9vNla7nClVYRRoJ3lUgGoMVwAk8bkcd
3gisWAOmA0aXDrah+ajmKali9g1YMvouuJRonDrhep772Fj9s5CrFN4cFPPW
RMYcVATFuxrIkwqrCURxCBMUD0ZYFe9OLTJZtFOQBUt3E+4I+S9C6lvXQ1tP
kyu09IPb00AB7wyT9SEa+dBnUZd8XaNsxHdY4pWL8VLvjvAMgalFhU2Ry2xG
0nObDxp5hUBGmAASokBQHw+0CyaxH9O3P/HrlpWbQM3PVlJ91vPMTzqNduPd
PcwMmc++n9ZP0zRi96MDUhtqCxUG7Imsl3vyIwzrL9GXmtud501Ng8MMXh6v
yBqApx4YchqJwGN6+p1s1s8EEmWCRBcUJOApO4VYDtW3nB+3F6kofPmkornu
J/rsVmYMVRF8JbS9TjmtNkZtJci4LYQe27cJu8nJ5ed8CzihcUQ2hXFSlCyw
idEp++PAVCAAWs+3OxNr/HynCQdMKK/AufPNpDUI+1CFN/YIr9hLqHI//dJB
NoA8yly48WVzehIG+eib21vYB+cKcOSsSQK0Eobkzz3KiKGx5uMRwfdnfc14
UClJmKicKXnS0vMSQE3lPzdTIbExs5tiAOXYt+w/z7F+vQ67C+/XYoTo34TH
RAt8D4/xQHZiTH/6q+A8iYTB4bk2C1+I6xRBK+VGc3I2dlK66cg1MCFzV2CS
JxL0fEok9sESWoxTWPnFNBf/SfdIVAAz8hcXy6ipmEVA6yVcaG6zktW6kgo0
AsluqfWlme/msA6s5coBQlMLdR441r7iUZ00oo2uLdv2E8sVreLNV8YiHLVl
OfwoGyN5BC4v1R0dYNP/PW7EPa4DsKFrhaIrxyqRi+Y3EJRkMmlH//jLscBP
NxPaYklKZK9Ho46EEGB3cILmdAVaSQQCXl85GRkhztozC2nzsDOKYDvhM0ZL
ZNwLuHWI5F8le4xJgA9rxHPzJNP5Jhr75aqCLykuGph2Wa8eZqoyAdHqWZ5U
ZIK96beEn3XYBf8boywfcRNc0sedk9cTXhTdiAkisvZrTzDlFPKe9DhaVXoD
hK4xUElsGhzbYg7zatN06JplPBcZwPYWcVxmV7wZ7p7ZWt72tfGKpjiNZMV+
bCJZ2ZH7Z1o8Re4BaB3aEUcs9hQXjdrOj5xFkx900KwG4wKnWvagAfTsAFeE
vnbd0RbXVSBFIx7jggjzeRQxwPBmdY9QzO7AHBsoWrKPaTp0TkqrvJLWRMrk
uA9KTfZG00BPbcy9WWh9esQ70Q94AsH6jWoQUrW3gC4tpbBWymuyXQSQ80XD
RywdmLF+naMjbqpsxCosb7AtvoQ1GuUw7KxvLjFACCPJp2F3CvE9/wewC3+F
v7H+ehj4zoZYQng27alT/YtkkxiFI/u4ZtAh0k9juzEGf0Syo5z13fki1ob5
huf2e2B62z/cenl7RUB3GqsbGJxzeoxKRrPhWYJ+ROPLqPUhHDXhxvxJ9vPn
TyZX0wVxtCO+SE3H9sBhHjiLtiZpJzb6Enx7miH+Qjwy40/1wOQXBXVB9mk8
dYfOzKs5BJpSId/7p17gomudtBXcTRc0rDB0bAK9A5IlW+QbIxJSK/LZBP2y
1e11Xpdl45MyJTEWkrXHBeqjQYdzJLf4cvgaz2XOOmuSQo9SHP2CkrryfKKg
UR6NyIFxnQ2SHpTlkSNByJh/5QxrlEeyL7usWywFsbEQI5EjpNbsxvvR8hq2
lBa7JdPNWkXlxN1Hvv2av6g5JIXMj5rDsUSC/B3oQYTf2xR3p42QHPlzOzOQ
DGXaK8nyw0CJAUgoOSC7FnEP8oPp8CmkM6yRz6TSqKtfBG6yKq/2Axx7uLR9
8Kt+jvGbjAZsxmihmuexbWFn1ooWto2xgzfQwc1hIi7/N+5joXUuy/X+Pnbm
ENwUfA+voBlxRXLFk2EiLOyzLqkisLiQHLTUlQe5pGOOu+wOt31uJPXWNbqZ
W0qSwYiIx894VdiFRBxiWO+oh645iOL1OGic2j29yS8w19Evyr7WaTAfjAX0
hQm6DsNrvhjQCyfJL8io9moQsLjtJq42IUlPq6zvFoFiW37MXk2wQb4ObJb+
5FmLJ2XOvtMopZX8ug1ayhzoH/+enT/Ew5xxv16MbJS3Xj2bqrPmbAshCE1S
dmEYxusQ6fiGSOx1KDs+3C4o8cCD3+Mnoye1NzPb8fDI1m5K+THjvB5ykQ0T
vnX0I4SvkqpSEIDWP7SMSpsY8iesqfwuLH4OyWatxs4ybkHeUqSrrD8ks3OU
nBcOCC4cHqIZWthm6jlJlvP6ddTnnVAN9cDOc7wxx74yWSunQE+NfS5LWrVp
91ZFT+RYmoDt4rlyhIO/CTuJYU1oLckOgxZIDUUW3x2WuOUVLMOtN8A6ZxtB
6nqq3DRrXDF5ijqBF1G13Y82rf8zPFA89F21snyBmbaSTEEPDXpcpm/S05q9
3HTxWXbtEoG6Jm600+dz1UCbSMl4pI3BZl8Mjqk/IwXJMcn+pjh7YWHiF6x7
gSlfStXGwIDBzigSw73M8o09d2/NdESo1+ByRTxdifiFkgng6oevVE17uVvl
JE6rXOBKnEob69VynfHnYzOKmcC7I6QncmdrGMMMT9y5C1HnW3pe3+xmmbo4
wTVAA+YPEQWDG/dntXZwBf1kaawkm+092Q/Qt6hhxwcY9A2uk4FDK1n0N/lY
lje4pVW1g6PC+Ss1On88tVBfnwnmrcw6lWEYtjXdsZx84HE2n2Nkoy02ziS3
wrvU/FhGpQRBHZa+6/mjHWGIOwckp82PC4wcEjxR6rumfpte9BkSiQQYjK4J
9ywDQxkGFR33PyU7BLe7HiDYiiZFjKFB8cDW2lIxpdU+joRXPGjjQa06qRCn
Qem8/V0OBd2iuLdUFpsysBTe4qirFc9flNjNIFswH304ptXGIpA4fBtvW+2E
Z/J3kgtj3A0WETzJ5gSrr1gLvGhubthOH9i4J/sHLACLJs7QdQa9QYXsJUOj
hvZClqOhbzEO3VD88AYOISz9EhhnLK5uhOx2Nyzf125u9vScAYnxfcrwnVQt
cd7e8NedZ97/MWdduP2NK5y9SBfuFIydBjL9BBI1jJYftDQ+3YZoVascPIW6
cfVHOGHKY1Ernvk6BmwnFzOZQ+G57fXfaNOPWTvBXzjyQi+sA795k+1Db1h5
Ovi069ySL+KGeTbCPwjYeFEuOrMNjazaDA5/DTMgM6D7Re/HWex/PVrUgObz
PvSQ9lz59qpkl4EFlO7/4KqHrsquPzJp3GAcw+/XZV9LlDzuYGJBcvkD0JEH
4ZVP2PChH2O6p/SwuUzpicFBzh6Tajw2GSagujRASI1yHPJsg1mzHm5XLBrh
25G8GgPlG/l5QcsL8WzA5osE2i1kM1i60hX181x3X4WeoKYY4UxbkEWnHO3L
+i+S11MadTi1cC2Pc65/AUerfsJsKjB6IH1JORg9wr7vMmQ8dt/M4FhK4a5v
BuhEtw3sws0A0uk8ISxW8/dAGLSoTWldO3jy6TFTRMSDXWqe3ZoCTvn6VNT5
omTzB8c9hrb6kl1nFle6LrelfwDGeo1heMfrkMH4OOVH+c9Mtcd0U2Px1SLu
zkimD+mIaYOnb0F8Eh011x9qyae59l7ERIL0mf0wSRoTyqZmjBUeuC5M0QgZ
gUT8XOPyjaT2k4QE0Lw6eD4ZkYypjpUNuD1zwYwR0EOYg3R06xFsTjMfcIs8
aL7h6qzWycUZZilBGrEy1gprQWJ1sPzHSYJgbHia0V3PurD8PCUlYT86Fn9/
4VLw9s7OcH3XJu/EEmojItMzM7EJLj+DJ82uyytxSFHcd0AFW98RiwcHiNoO
qpcuc2TFXlrbcbYhIHg723sH0zv+htuxn798caoYRBUMdleFRsh0x3NI7In/
IjcVhOFE27ydj+H5b6xT+MsdgIFXrQGv7iVa8KxQ4/FR/5e5rZS5QOT8KCGo
uoz5O1U4AheZeBW7FUOIkTFDYYuKKsty1cnxjRVOFmYhNsfy1SM9r6JD/W7M
7G3iyIJ4jDPPpGIW7JTnGS0+N01IvWCP+kw3YYpAJoSGXNgI4tc7cTNJsCeo
rqd7Etmi9FcW2bosPMPZ713yvoJPeG9CFuzN/pHEXL0wipSgWy1eJc5zqcZW
ST+QFOQ+/D6sNQ+1pPdyt1Z4ahIFa4itZAKrx7b7Uq0rlN9BXP5xnDjbq/xA
obtZ9Cp0pr6mElLM/JkMODlH+pnO8imUWSjozJb/B8uRudvMq/zIEddeARlM
PnS6HjJd9FV3OxvGBvEHuc1esjvhqpuLGgpVrnajb/qqzxGSu/fQcMv0yWy2
41nkdYBd9ahT8Rx0GzyfpdgX+epKfhR4BuDFnp6LBZmYPKZtZEu1P63AnHce
Mid/Wjhoj/oZTjZbQpt4BUM/QfmJwljUVCBJCn1Uo0EywcKfUdER9fK/9ers
mvONiJgHIPesoB4evsOgOYIc+0v5Iu4ZZSzyBWb2sDQIdi9prGV9Q18TQ5AQ
1QBO+dEz5ZCUTun3mXEgAZ27WUFmfD15fQ8bR/Kp2mKgs8zKi4Ph5/TQN4oH
bUQIWB7ZHmJJyPRs7QRaS+S9OyXjwtn5aeIvaTu5iRiTRWnrSIInGTrU9Xsa
1dhJ5e1iflNKPIg4d2rrZwxkVhGdYyVvi2lUxGGSBHVetXZK9es1QBSoXFQQ
eehOO+y+iCDiM6CiIWcygC4L7d72st9N2gt7KI83zOXccf9yNpH2rUw8fbYk
pIuAZNH+uIjDor92ymbxHIjSCYcwyeBFpzlCs2puRRsVl1YtE3CH4NSUNjxS
5C/j34KqxMtQOLGBZjalMlIw32nRHQhqKwYqKVWqwRa1rAozl7oRibBGzVub
vaPOU7eSWfWHcRRsASRkmj0lF4KTvwWh8fsFjZUrjSwHxrwCGyrDeCyOY1ka
6l2goTIx0AjW8eC3W9qp56mnkVhd8hHZPV+N0cj6LQrv/0BZozmem4yZ3+L4
4mQMdewE8YjMYWghz2qFauMFJKkVwwcFXK8NEDMbN+KSkq27zoyB6CXtvIcJ
WQSeqi8yZuvK0t/IyIB15ql2ftWpL7WGlS8lbftW2LNQfklwAYvPs5LJN22p
h88l7HPjvnMfuxVOe5Ts61U0XHZCzUv0qpPh4c9+vuFzGB7SbvjKZHxRmmpO
QNs/dk1D9NKoz+UJ/Sg1OAHOuzWC04Lkdcy9TAkh7EDJIlI4UibPeWgU7Vj3
xHyhxlFixs8hMdyIPYPDpOLHrREsUoZvwzGXTmpOLiAoCaBpbnTzWO4SAKSY
qDv3QXEnktK1R7JyphTfD9OPNdZWcHmVh0OtceMXhawWwZJNZ4D8CkZ1trr6
9fJ4IuthMMnfFhRe0tkrC9MPDg9ERx/qR4V7+kTGf32blVb7vQMcUVDLxpp+
OTbdvlNS2gI+E6KiOxpAQzRlaJcP/Puy0qixfm8JpQXhN3Rsaibpq+g9z/+W
Lx4e0Rulp7avRat0olLqjlpUUN5d1o5TYIo7CF7YE6GKzOvM4l211VUfvjU4
VLTC+n7Dd26mL6SNmKdlhQ4OnuulQD7hX8c+hAGlsgze0GNDKcDMthvzPwpv
dxm9fbxBIXWVQ+vbHGKjMc4Rp0tfSAPlwdgigI3hR9aqpgZZjoJhzHiKWDUz
3upzW8bx4PJ5UsYgJ2OLY14MHLZ7CHEqI3vR6ET82Ute5mPRTvZPlRC1e1SV
M2jrhQFz+dhC4hKDC5Kne09p9M64NMINEVVS3jxKI9lzaf2GfDhZCKZZyAhm
B05VVYo8oBtYMqDgCD2RzHIXu8skN26mFmqHjEZS9/S8medJN7YrwPSmHvdh
SspPzNpnJ24iGGfZJIceFeevcZrKdFju1sICghQEVW8j9sKMhp6cmT+nuGoE
5I3DCLTlRw/ePm/pdeXfgI0za8WE3gOqy2tjh05iK8og3NBu+/hx7ix55pJL
6t+hX5AjGkeGm75ZTdQ50r5fHQhbUW7bBIYTLBoCPbs3lwE+7DuZB759GtcO
cFPzqxsPRIMFezaNLyAEaDliTG8ZiWtdl67rDXpISVT/cJtGK85FqPbvrKsW
amHtBmze1q0PHKGv4bHB93Nn2HQoYiuBssRaQpoEdXF1RMWfBsPp72hTSxJU
ED8TrXt88tbWI1ndjO9RKrFe3+BR+jqmWomeU1TgPT8bJnMPMPvyhG1vnBT3
C72zCc8mcYEUeM5CsKdZbDzvU1WdstsSO1iKtt1L4jc4aBVVvATtCbJP0Jjt
Cj3skOQ524mUXv8zRde8NYfOlPCtmQSW8Q1BiUKY2jBLeFNI8UrQWZIucPlc
4FBBR9/zQLsVNFW09FuW4Gp15I4CqNM80L0rTlr0ZryP79UaOFSljZsWYNUs
O39C6rnIVxathehfgpFHruJD3Sd1qkuiHlTGIglxFtCGI0S5y5TCsVtYFLpu
MNsCLn5lNw82BLkyiveQmfHVHJ4MJSNyxCtUFC0GsL1ww8yI22R3BwIrLojB
+aduYVkLdQAlR58DinTB85SgCLJVL8J26h1yVIRk9k00Q/3gEJPhHfRA2K+8
n+4KWthdRRYGbhXaZxgGd3pO/0Cw0mGdgA214B8Q09H4dbaOkp/v1/bUVtKb
8Akg/y+3LROzJnkWONS+bk5EeCj36vClqE/vo7shWqFYPkUTOzkiGkqGsRW9
ji6o0hhTbd4oAOCZ3kQRHRJW0P3JLm2fmOiXscoDm2Eh0s70sNJs9oHXExEr
EzYZxAeBCPOJLOMt8cm3rQoEWEPHCgX7fHWUnaZpE70dHGsaxvBGeNRQrPUJ
2ke/Zw3Z+0KfqVtfqAW3wrB4ezCKKRfHDwl/6tatHZAUEiQoqu9djdNwc807
oqZXSJnn9RUK+bxsaXof0uCYGp0bpOLyEMS46125nWbMMA0v3VDQL91kfQlu
tjEBd3wVCOoVDD6tY2i/tCWSNKUSI2LaG/dkBwnR3wTmCY+WETNqPxQ1RXQS
8tkSPw0XejPwen2Knl9fT8EDAY1Raq/MXyQenZj5kDpSky4fKwmm+03b7hlE
6WyC2NT1af/I/gkycvgekjAaap6+B4EaVjQaRXHa5fVyjiAUe4Q/Kksucqdq
RyCzHwg0bTJAE2jDccD4aB2VoWpnyNcg+X546TosKZBMBPkRxTerNSPGERK8
3YXeKxFuZ+6w7i9B8V6gWDO90e/dco6jBgJOlYhDoqh+MdRWWfwXcNWWj1oJ
4SAtOJPI4hypIHl3nmkBSWXOrMaR5XZH9cPjG4Km9/rQRtEwkxgxP5LmJn+1
TMK+ox/yieexYd0esBtLut/ERZMjfZki9P5fvwaqG7AVd3O/QlkFf0skwFw+
1QO0kLrVrT5/xcyHjLixgshLSRcB2T67V+qe3HmOurw86OUOQFT76Fv/yjWR
niNvsieaPkEf9hUHvOoUmSB/gWNYfk44i5Np+qtIuIE+IdqT9R67FJGjGgGh
s9QTrJSLeoGonZTnSTBWWUYbk5PqV9UkW9X96nqZTT2JlgtT6miYxYWYPNo7
AQ0HbxWEKSW9ryGlOD9W9Gg4yA3PrTF1V0cqmQ41ig8UKa389H9J0vAzMEzE
lInzL/vHmt1geVfkoW9iojUkVLrmwZlkZhPgblw4v12vwwon96R5BCvIVDHY
gL+LHbSDtz9Ywbz96bVPEcBYtizcsjJZqprB5Kz8jzne2Dw23oHHrIwyFQ8x
eA9jlFbXVtE+pqLzJAMY6r8HtjO+U/htjoKchFD24NI2J+6FVDsDrj99aJhH
k4RMJbD2lmGCSR2rY5QXU+gdxk5GpQz3dOqD7uhdsUIcUT2leQV8mGMi+5F0
GDfTcLOanRP/v0/CyElVdzcI9IpYILwIYfJKtkh000/rW2hPatYrAm/iCLxp
9bgCUUp/Dtg20QCW5Hq+Ux8VLrWATgWEigf7YbJkRDsXQwfj/hb3WW1mHTnU
H5HJ7YjKkIiQ4jDppg2buZXDZHWn51nXEamt9NMgHng2NhoYZdS9HWrg0Jow
ISLK7Fqwzwa2seYeMLlEJ95kXgbR+blYylm5Wfrl556ikjq7o+1Ay0pIg8QF
FVvJt5qZZtATTxD0PImgVzK6yNRjQfI/cWlIBkN+Ef8kYKbaAqXjtRfa6Ahg
7nTo6O129il3QmO+rNSX332WnaQ80CTKXVJzkyxr0kLZxDKbHbZ3q66nyPhh
8orq7RyTSznZ5dYCccJZYrq2Mg3GQuI6/OLG7WJYOUPLtz8rj8fonjOYDTZo
4lmKCAVWe1ZOvBWxeQDrC2inLntjXMm/ibtKg2f+iWmo7l1jaow+xYecBHZK
ZSSA8+yeF8CHEr1QTDfTqxeYXKGFvNWrGH6HrTsDtcf8CrOJ4IKamaZeOZ33
+jKhd11ULmR8x5PBDz6We85Yb0dhe/Fr+R01FGzVvM6Xog/hxI33Ok1RROOu
/o3b9Lvd2+AFAs5otM/nzwHVu4Df9/w2s4yl96QYwiMRNWaz7FuXwLnIQAKf
0v28R3FIGFBjSRi1U4NS4sr/uw7uA7bGjEIO4qXIDvnVuHZtgJrjHVmmJc8j
/LY76KXwDvrrwD4gMTk3PwrYcJ2tnbxP/3uOC6Jb4RgDHqB6CHNceUBfMrYw
C1pOEj1apCcjIYRfbKEy5VaaDPZ3Aioc5Kq5iFBy5rh5lzgYHLjF/2nxuaDy
tOvpW4Lnq+8/u6dI0S92AY4BjL+g5EqGA3d2JARKNjtpf4KeFj+rBrc/5UkJ
/S+HuO4PFsNxbhATFIw9s7qR2VvOnFo9Jwc/NucMkalFNynQgznJ9CfId7OK
hN3JJE9u1OrbSk2NgZb/xLeVToFE5RCkxdiYHuVuMfHPubs9egQ2gjqgvPU9
hpANzBBMSqgvjupCSROOZiB8bwJNTjCf+y1LWa2B2bRtUKMcV3nVnMQI8NTv
VoQOE6mw0xiScmHCxIxvusccOfka6eS1MReiP0FTiKu0USpedkB1SbdcGdYC
E45h+CH2xAAcy5k+DzeTlmdmmfjU78LWmYJ8S6AJSL9zRFv1TYZJ0Yu2XwWK
ri1TImD6nKte/p5sLW2RKyZjmtvBG9AF4V+84ZaHfcGAiIciLitrDrlpNo2P
KIdn9inHEJBSZgLag+VTuilbD1lhhufgr9PoYu6GcDtO3uwzIuVEC6bhSahJ
bTyPU/JrQ8BNQl21+/TI16tMpnpuo21AoGV/U1ivpa1UVF6tnuaefRu2Xc69
Uz6m1WOenaSppUODiW9WVjYHeKMeeFTB0RA/vlXrGqjwI8pjFE06KhjqGNap
hW7T6rygpNrpUa5+cBZBpqZTctSxxRnMXQ2Q6E/o2/nzmgipaF9gxN3Borjg
gtaxNSyCPCir053tGX9lMViuuZs9u7UbWHEok0+iKWt0xlETybUJtAjdnFv4
bUBY/Z6pfj9Vz/qOHgZJP9XFP7TUmBWA8eCjevCf1DVd+F1N5nmgvOEZhQwv
O0WyDndsVOBvVzJRZkPxZAoNaHZ4gQaY49Xg2Xa2oGlF9gTAtlzaMS5LU93X
ulG7WXwxrR4hopIsTOD1CTd7u62l7TLZiRmwzA5AOzaUu85srpbHUf+pD15C
KE+pdJTUnm4Qmbs9QZzXlJGbYGp0ZQXz5zWogJf8SIIy1a1ttSFR+R8Vv6Jv
zlAywu//a63ywVnNQfqGdIYx7/tw5keln0oTFs3hpA0DZiJQ5iEkmJpqzsNF
Ssh0qO5exFuB0YtnSgV0OJpH+YZIhCjOxz7pObC1R53JuPUS1WFMQQKd39FK
fEfySaH4fJ5kPptFO53fppaqXJ8ouEPLSUDJ9kUqonNlZZ27q/zhowqUluM5
ylqvTgZq4xR/USxV2sP3AvYvBQbnqwGVUaZXZWmpdW+vuV0buytpOeMOFwVV
Q+zn+oziiv533h/xceDgP5X4Y/JZEMi6SBl4OLz2a0B15DmDBotwsRI7nmsz
G9bpWAKF7mt6RqIsW4KfbLJTDQFdGGx67QmZzxWn0r8rHARIX9WPcNFHk9Yk
jQG3omaK+hB5X7bw+U7W4HwDkS6WyDZ3DAtcHK4hO51g2WaoSngSgtspICG0
vWPmv/u6O3jKkPT+LoJmd+O+5Bg6E4JXEzbFGhKi0qCr1zALdo1cIEAoo6bH
5PxQ9ePy8b2UTSLQ8PEEZaGQicvT+AvfHXFdA0w6j8kPVeF4PoT3txuTrLi7
hVt9bDlvqv9ns7Cq/2uPgIfMRT30u8OjCHx6TpQYZR0RXLn/y47ikcWX9ZPc
Bkwju8uh1rmVoEIuhj9NTNoJhdg3KlnLudQJVH8GYDhqYdBJIEw741jQ7lWK
PpPhTKAT8YdEbe4zlxVbN+VTolxD409C3vMjWnPVyUfuZTQB/lewcwyG745u
1B9eXqM5YhRr/d5iUSAlMQEk52TZISHfcbQ1/fT7ppQDkyx2wNfBXaAhzy3X
UR3d4Qm6aEufybeHbdasO0GjnFM1rSpZYHZwmbr55H9KQdxFy7AttOTh74+r
T1haSAokc+GdAerpaN0wa1mZN9rONKMwh9uzXhrwes+YOsYNMzYFXteTkllo
hSaPFeDpzjFgO3CPt5nJnwnqY+rgNFeVnssPN9sAWLpnjVbNQB8Kb+kW89Jv
TxjeQ2FkV62J7lyBmjbqeC9TAjSIN++nCuq1GJr8YESeTfdeV0hggPNm1fZI
Zj9os4iyAsU1QbsCWOUBChwoksn2dTCDcQSpWeb0c7A70P8u8A8EPJ2zH1PV
8e89FsPPXWE5axkDXxArynV0pWKrkiSU0Qv7uda1oSC8E5ixPKUR/ePnfZ7f
U9+5vjPgMoQk+lfrqhtbFDYDPuLZoe4YpQcr9abqUJ7+X3T4zhfB+t6ZkuvT
P1QO+T2zoYWiQ51dVm2I15iVXlQDaEYNBJcKOHLvnWvGF3lGSj9Ws08b7SJE
Rq3ohF5DPOm54odjhfcpDQGI4qja4C4Li2YPa/XF5i8SDIAUxCxltTM6BXk2
O7OyNU0Kd7+Ni+NjhwHKeOrqYCXMkmclisIRg8wfDMLLAk5AQanrNM/lHaxm
fJvQhJIGZZSoo7FN9pjQYiS7tUxlIRQ+yr26UlhyhELDDUj+c63DoRXVvgYy
pOsDsi4gV6d/mDIBMTgDG0KSay5g4oM8UY/YKP2JrxKUlmxU76oGxKdK/o6+
t2lFQQtwFy+/cXEU/oRFvjfMxHkc2XBfZqSIZilCnWRZRbbLTGQTLOZXppRi
IOQdoJTxaSKgf43/HbEaYeltU5fjEM3fhEYJAQzOmBvmbpvLtsycSTywbfIY
IiyESnr8pNvwjcXgyqpYr4JGPM4Dt9LbQMDdeFO3TPggO6xHwg/mj+OZoeb0
LdbFvSZ/aCnAA20XVV6O2kMtomOzEceBAZpI9VbgNYZxaalPq4iIGJGnA95J
z/qkUbQ3QWrjezHfCU0dp1QVS4uOmFlv9eAxFm2Rf3IdJXd5R3v4ienuMWJT
USiyvl50aHgbso3BfMWliwOI3vlKrwbJrcfvdBkvhBV15dkjqCUmwOcdr8cs
0LM1cFUHKTDLg0afiTekBZB9s+FzYR95OLsY4GUKERtwPYtG5SNf4MYbUwIM
RKnLMfySBcAEIpRJ++BzngVIieHYVAxIFAY71pjswuDK5RExGRbzO0roLEr5
yDMKnLfLjWJWQdvtGvZKiStRn90A8im31Mm96Gz3Et6oesbbqtM1aU3d4va4
wWWJWh4eYMBX0j0vfHCheQjCCrVwXXoTeHa4XAMuWKTNo8ZGfsZwv4bg1jEz
kIrsySuuokhAp5btsaVRmUPAfOyzvqQLNopM1UngVrLiml/Ce6MXH3Gcq6WF
9d1uNf6gjS6PAIh3zPXlHgJ0fzFE5mqUIyfWdSthGNvKALkb8rFZFrEkJatQ
oUQMK2cVz6EzL9TcfRt5QTMY8jHfIFgQUuNfir3u4zYvMHbSvPHEVM6TPIdM
gV5LVuD12y5Sg/V9kpx8ZkuC2MhAsYdWW//3DFyMuSvyNjA9WRzHYifRRNpl
R3i2F83ygLwPb4uqhRHAWWFyD0NYvY7XaZm47pDjmbfA5B4uIcZG2H/6mLm0
UhY5FS0WY38KOw0F+Hj8fw/8TzIbMEtQG1DuujxbbEWb1nEL4FZemIMYpLWq
jDp5TUBVV60eXZKapVL+/8dxj82NfS4qS9OOwugIHh7wUHUijpGNssMovby5
w3bC7k3YojDV50N0vnvqdFcLG774h0liK/50f/pioOlKkxerOVYO0SDISPIF
F02RmuTdrclMQIA2475XlRvQ6t+ulvQ1fPY6j64CgpQe+JMbAZbNBbKaNQjD
TTBjz7IrLb3ttHKZ3/gd6fwpP9Bi7nDquSKlvTrutRdeqvW3aCNgJYcNGnkJ
TUK7KiyWgBuonw+GNwNTdI3K/yANqixtOZsKZfrbSIY9c88KuB0Wmkbesmum
tnHZWg17aVnLfBmEdenPqVrt0orpuGHPhdsf1uMi9w7wAfJ3xhJ7fwV+COJ0
1XKyvn/GNKMf8fGKQC4Q1U4zswMQlFi3cH1r5XPkGRFCmMWvBCcwEWFxqxGs
mpfZvrxqMzYJhlYnZ1gUKhRYE+mdlNgAiUTe4S2dATRvZyv6HOGi4mFGkjrO
efF8iHYUNIG41rpiP3RyP8UkbEI5DDHiAPwckl0z3cT1dqJdKmljBg7Eg0Sz
PrUeGj/kWWLnL3ixUFvrUDE11/p6cXgoOeYpd6xY2DZt9c51vgzu2oiuFBlz
+MgCDWlBPdSPrUVpaU4WMo9SG/ooYw7YmvH4Ts4ylYoVZkqOGe6sYSCzxgLG
OAFVvwtpa1uLpeBpLY6BXHmYKVZhz989oCZlA0YmseUufkz/oiPD5doaix99
jphEt3upP7/sJ77Mk/t8WtdHQWeuoARfRyVGD/RphfrqK07SMoM8zcGtnk55
jo3fL22aaFf0mMrlMEswKDFsxmX+IsXeSCkJLRey5VCbyUl67eEVZW7OanuD
4B6X/U3yJHAO+PI1+b7/XbrY4KfR9OwjH5L9mkK9f8BkDCXv9Mw4qrEppjkf
70WmsN79Y10x38T4QNkw0EJ/P7J8g2IMuY+FPOLPARyko1nVmINJkH8BK7aB
l21Bl6th81ZFov16gC27UmYmpisqoPH9TQeWKAkmsv+kveCr84u9VGMNWwEW
KL6wy8TppTAlTpZovGiIgKwRq1Q9GKFknBFPKpcSwUSpU++WHwIAzpk3Dna0
RYC+daQNsd+gV96OzWps1esveLPP+mF7wUdk7DkAISGdNDbbwKb8eKsGc54F
wpJX7Ly5PVS9nBs/WpYll8hulYiJyTZLomTSpU4jUrmYv6Qg3KFROjB9nlrv
aXmglsjYsK6RC6jkmqhNbyZ3UBnj4H+lRqSta0WjF6MYD2466XUNCSh3gL5W
7DsuMhABkicBBO7iTsYU3NA48f6O7OuOUN2Ni8yDAoXiuSlkNfZ+TdIsz4mF
wPeRKJ8AduEwx4tmUbJQg8gak8cGuYrj9KR0Z9AsCLOoaCKolRCL8bNhi64J
t2TXZiqsTr5fjGcLQ93sUFBJ1kCrSPZaYZL5ARJEEZFTrmy5TeMUlNV6qJIK
0Bkfi+azZY9sLZVTI9cg3Xd/rVNzamQqSSWRp6YUf2RuDEPh30aMs4C6ZgXv
ITCgyW9PekS/nQhyiQGqlmka1dI0jVwH9/oRGuquB/FCbesi/pAregj0Vg6k
mTIOxSs2cFPylyLWkbAwDC/6PjpDjpHCMGMLkgPZLCVgzQcm8B1awAA9qm41
UJjoWlDg4lrERawy+nrQK6mUjU1rwlTMhO/vJQsumuUlKU0vTxA+122I9TSY
HCUS6yiXSEpMM5c4EhV7VJ3SUL1MI0h66sNB02Q6yRTLCIAPVL0sNb2Sszg8
kP3bl2s0JsM3XDDTQHToHSihuSsKJti/W1fnfu+lo70TcUe07yAFZ/fOEmVr
aqpFwsA4TSTHm2nxLvt3dZEuu+RwT7uuLuFP80CsGGF1i3tip2aXVg/H4FRS
of5WfqFNFMlD42j2E+u1yD4NbLrnjJj70IA5rlFE9yabGDGy0NrocHSgqihm
8RSLAuFvckUeknHja8q1ZuBDaDGPQsl31dIkTPG+mMwtmNznja0v0kW/fhuP
Og7E0YJn7bOPfzYQf7Ip7VTi1RU5NvxswdAaVIRCkOYI5O0xqEqBf3GAza3r
eXkFwdhcPmwiX7SDOj5B9oth1K4JV09H6a414w2sa6uxW+Y2EVOuHCNkzBOq
MIb2j/qelohpquNSZIEHWwDFNAT8nZB3JKZ8/zxeJD1S9z356W9kAfmkCmga
TKhGFafm5O1Zvj+Dacv02VquFLHjDVqGH0eq0BV8jXD5C5quhRUzvAPjqJHh
s5KXwigSVbmkqhT73cxLCMAT0it7xdPOnQjuK514MwWTRmSk1ibVn276TF9a
hJMWI469jdFVqSpBz5L50NxpMI1ILHO8yHKyTMJ3jfzIYGcoEUKNU6hiI8ev
ci47DjL0sOc7NLUcI+Jjf1QHkpg6JsvgKMYAfEvIn3CYmFKYGJpscvXQWEEz
Z7qJKtWcQbB5RLIXYSZfp1GTttsL9P49W2FeVAlBoUC7wlpD/+w7OzH98lki
yxCrqS6ydm1chGw4oPMrLjrUVyVGad7z5TsAhE/ERF0JaxwZRkiTFcYaFdEx
t3cJBPHG7aUDeW40E9eRrk4YRUtswFHLJLX8zijtleJk2C5ktWrz+G4loGFJ
cUXY2UOZs/awSanBsT+mEdlLtE+27C42N/N74mJeenA2ToKgOQfM1LuYuNB5
kQHP9ieWu/YnxTA3WDzbc36jiraH+o4OylYE4GQuEhcpRjReRHw4z0kovsGv
gnndVE5M7sI/xNNCDhfnPJaAJGNJaPothOMbAFJtlYWYuqcq3HnH4roYhD1f
jtKOnwHtxpl0skvT3P5byncbV8gj0+d43vFx4pRvfkxy47lMwx42iGP3QvgV
np5Ltikyt6Oau0bL6AxlKHw04AAgLf3HvFdi7VMdGiM50tOyDz86yCisXF/k
wb6Cy6HB8++aCctOrAJSaMVHFlcwtJdir1nkgeeEfPnIZGqAw+ZuMuF0vUGP
DA2PMBPH3HVKOBoa94vX0SkSQcWqZvq3KVyq3VYSZqiq6wMSOvLtNHjJ+1DI
fIHCzTZCFPTghoHDePlNVqKlt7CwIVX00wETWqBxto26jQltZKXij5wAFoYl
dDTVPo0zMJzC3BGey/beQdavD3SaTJOsxkKD81ztzGER/bItO152mbzCC27N
myb2EdFWQfonjZ4mbihVfwTSls98BVgWKWhFlglUmbwSORdSVAKM6lwSYkYx
2swMdYOB2aW+SerxiUUfTbYcUoZ/tHn+1cn1sT2TvnJ40h3yId8F+8pMpWgb
wff7xfQ4dfUtdcWAEB2r9+hckPItaRD5WJn9AgwiUx09Ijo2dx1mUsMWVE+q
iGwqTDh3J4SUoeaFVKhZ0O1y+vbyhOEBy3mJQaFog5yeRQ8LpGuTkuEWvV/J
kIeedGeqj3N3bAvagxdk27TnHzZLxKq9TrymPtuHaTzgROySBOuysOFkCU6z
Ale9qBzpholRhay4vg8eCji0xp6+C3jeJQHjao84CHF307KLwbKl45gFcpPr
O9UhmPabkIdyGqCyZxglJsCipCh+PPMPn03Yb+2IfkjiMX0XGpfOrg7C08VP
jCC3OFmqkA9rwFEt0e3aZRuF4UvNtNvmZMOszGzueuC3zLuyVaV2aX59K2w1
1Fjqxrif2MfBxif/7c4ClgYgTirFjRAT3dyue78bBkutEljI6cSdKP21ri+1
loQo2pgP1NAQqALmW0+LEeJmxaLi9is8iVHbibQFtEGUg9UotxIsaZjkk7Nn
gsqgwL6eZ1UBcz5UWamYEuOPcmGtAuPGFXs5FxBcW3oTXTEV3bxMc777EyXe
t+hqZsxez67EyJ5adzRCW2a6gIpuhs5o4SfzfP3cmjYejBFCU9PM9+E3xCU0
t9ail8CTyw5iPz3QaO6LM6EpCoCg9Fj0el4enDDKvtHTWBtkgiPSNsMqbnux
0udNkye6iIeOJ1XSsrSS/b6X5+JKMJ7WPlEftUItxbAQiie6ypjQIDMtP6b/
WRf31Vp9gBv+/oR8gglZ3ZlsKWNPm6MisiH2ionrlO8tVuZc+xma6OO8/9WZ
o3jIIYJfR8pW/gUXQZtdQYXFhZA+AzAvHuxrSBDz0YT6UGF9VAygaAVWOj+Z
VdbNTnen1Q4cexqPILb3q2GljChNjxwqTrJmi0lKiRd2/DShj1diq12qR+Hg
jPLc0mai8VDrcqbALVKbR2YH84STDeozE2nLZhIEAn+vlX+E672vSeKRyiza
5BOxH5gJJKQlAIB7TuHAJIrLBSRxBmy5bcppVgp+h90z9KkcoZ8wT0D3oLoi
enueYLWoQ4w8BJ0RWDKlsQ8+cPF33RexCs6xHi3MsaxDvjlAlqIE7HUzY8wX
bSoYA8h+4DIEQ/wgc8cNuXAS9mCUM6mABKqj+agVstrSo86MbXoCPtkm3i8P
Kdu59mCNw3LB6QqOXpbU2JTaGoohIYfmCfDmVADLjC6BSt0pOdC7vo1mrqEL
kGRYp+9rDseu0rgLXB8gn/cjtQWM4D/WWDUOf2mPbTZFbG0GQSG444mCy1nA
DQHnFQxYl5T/p19XMxdDUTH2DHYdkCBlcCE97BqJi1mJrnljRRzC3DabbfeT
+fPsmUJW8k4AlefKF5fYycjGglMhfFs/dB79qBFRh6yiYKv6Gbpq9TuRHYsT
cRY9CrcjUbm5ztsWhdLIyky/kKQsoAAaYphVog45lQfDQu/mfpmF6z6a5kmj
AjzX8voQcS3bT77nJHUgw3UlRen16BDOscw2l943y+J7dOp6nQjS2ffTLAQ6
rRVE5/e5LrWSQK7dXnmtUpHiwacC8ayvClmmrMpYW1ziHMicpyVkhdsRZTLa
5nia+euAqukPFUcx4A3MGhoYzK15t1wBkoVfX3sAywF5x7kiipFFzNBwEl2f
at5fvjK+Xh3O17gUbk1ildtmAe6tbKiaokRjsHrGrHl9z/GYv+3sx/aGoOwi
EptvfEsjC7CN2ZxV4bYlhqqXm7mgQjykXTKQ+xmzR2as0bt0RobPJtDoFd/X
2Ib9J7IKPRN06/ngicnUJ3gyR60/wIH3unLA9t4EWAAO60Jix57K38Q0V7ww
6klAYwqKXV5phgBgDllAUHdhj/MZMWBq5kld2VeM9wQipzPS/deaAECPmgr6
GKoXvCqF+zkBSEOnQCAez2yRNI3F4EbrzCWqGd/19/+W0Fk9Id2TqUmRVJHF
mS4j70Lgbn1UJt1iWKJBWsMpEvCN8xAVCDPc+krRK9MVFQIJEdaqmvAgTZK7
dolvB1W9As6XXhdongDZQ0uO60mP50tnhHYq4Sy+8HNO7yPWGp6G/Je0c2GH
ypzduMS0wH2T/7URItKhg++2OMP7ptWF+J1n9K7cIm5ibVO4oGgH0HyAvMAL
x7VtV24swKVLH/WUnMUVv56O9vmkNMKesXk976juyGEhpdLyF6JXWVNXnRby
rs5BMG8NKZkcaXLVJhOXgMSb4Y9Tec6wWT95c9Jtc+03rSUVPYHHm4wAc9FC
gSukrysYAr6VMdi4Hd4QKS8Hf7s91WvPoom+afowKnRVCGIKOd5l02BpLPDw
+Emskr+1P6T1RuowpwmBBLEA5gfZ2VmEl1ObifuEVYkkJPllZmKM24lpMQR6
rWqPen2qy0Occdv8nQwNj32EsLSfoN7LplE+zumdKAYulrziQw7+tUVhn1f6
tmozmwT+GIGLTKF0mLUGHyKtZQE0jc7JKgksMqaNhlC2UeAkBMgQ0j/rt9/S
Lm/Nwmaqf8qK3GWOQbFJ2ooTCp0QshoTsTEREO4pXeV3EmPIpzFYH3vKMFEu
cr2pfWjaZ8NMEsEGzV8qg0uOIcHRvi1Cg9wq50Jaoullfz2EhxzTpZC5NCAp
pqlDLDMyHQk0SNiXQ9eoJJt/1Dw9KJN2wRIqpHF4bT5n6OlyAmXhgSzrEwjd
yeNKFyL8d83pqiBFrUT9yV/h3ahl8aYkKLbyBthhsQOGqd5fCHbJL18U/MTa
qI69x9pieIE6VxeV8xgitCmhRk9qUFO4ZDBlWve3Pr1gyP80J2/g3NV8BpBX
btojwjQJV/8e7DKA7ruMUvZYtpdB830BAPwBSRjJxTJ2xIU2gtjHG6oeMs8p
OcTQJpd6BrjFG5hDNcIFpULtrwaMBHv1n9ehUis7d+rpvZo6iFdTUlD7p4Z3
SblCF7Da1AeiDtD8HOxAr3bib4G7zAGNYJ1XTdxTJir/xgXcTZKhoKRl6KZU
rfdybTUeq2ycUa7Y3JQ+Ar6XuZu2T7ZI3174OYJoBtRrWMO25BnaL5SJkwaV
Rz6ZUSNnopwjQnA3F+C9SG7a1PygM2Png4a1AsNTva7GEEElnkzIts/p+efr
gIGGeCGd+dkW/2H2FaxtiipMEyinN/9hin2GK2PkNgQgY2JWZQ2k0j5T9jTt
SUrrdx9Oxh33Re+Ar5SN27LwObJw8JcZ0Hk8okkMic/eeL44SAnTxxqDx5ZA
KJsozv9KjiqK+OKXR6KpLxPV6WCNrDFoSA5U9XkbwpSR+aodF72gLsvDtDJV
IWLMB6A5dHMOCXDalnHCH0A4aqKxS8X0rSALTL1RZhnfbPVPSo2SzoIgDxkz
FyN5f3ntiploLE/qsW9zLnMgMF5UgrIjb5li0p5NU0CmPisybYP5tLKtRb/i
uXzhJzhIFzXTZP00Gf1D1twtkRvDBlAO7xOdz/1goVQN3oUWKiOIUaj+/p2Q
CKV11cTO/y+e/yjkhcpN3kOg8NMOrkZ3jq2kEbZaQwDBDK0hTV+tXWkuzBKc
3bpF3ipw6htGbbwt5osIpynA6PtLBnX0iW+AN2r9rRVXdZEIvLYI7MadQRwq
PoMJKk6BA3K3dKxe/IWm28m7t5E/KgMsD8yoZ2SvN0bfrCo9DyYkC654dSiQ
W1/4CpHvi/iwC0PuKOD2p8AoI5iK85ckk5cUena2/c0My/1Wr2R7osDf8kQg
V3BjnQrmF5MuCBCtzFD44R+56ArJ0aaN6zK3vPapnBSKabw3JbKd03ak3GbN
Q8BUgHa90AtT9EIzC1Usoe+OZM4Q89cpzwcKcZupPQN1C3EIlqPOj/fa8x7l
w311dvbfOH0mU5rMDVCi0f4rqWtRN+osXHHLC/JVuBVcBcT06q9kfgWZ9aOX
S3V54CUW0Uef9AWagOBvZMf1mKf/kLNqpz89SSFeTZE9h5vQEogNtGGydQYO
i3NR8HXWlOTGgperAPdUFBQG3CR30xkVdDFfEBqyy2+x3rbyS+wH3MHYSiro
VMKf546Fh5B1aIiqhDTQ7OQGEHkfY+K9oH1stvs40Zt62R/y3HlU/GUI8nYZ
hiIm8gKQ+5BWExOzunow2Kp/0KlGkGUN0KP3CQpFPPK8QD3sPdP9Ku7Dtu6c
MBEsCSVZUV0oeax+pKh2MOa1jRO66n6+mqx7IQG55HStY+ZW9ijDoDE2Nrdq
WxNniY2Ko79j1ONfWZ3rjMgk+x2pdni3l4RZzFVcmAUGunZEXp80vj3wloCO
7KSJUw4SQ/zuDmgg3ZHax9uR6PidtD37ovGv5tQDoWg9jMGP3mv/lQHVRjXG
fzGnNdi5nri2tl5yEyBRmIiiiDi9inZs4fBMRbxxuatFSUOASTXH/wzIdJQI
jy/Tr5jQBwA77Q03Or8H8T7heV7O8XVTilbzAm1ot9hk8Xp9QBHmDkaZ3Dm8
0RAjZkf/Js+tbNnOuUgksqNL55jrUrvqd7qXg5RTLf8Gg6spt5VmYGNMFQLy
CyY1LiHP0mPZVSBRgLOsu3PKGfRSNycI3Ebx0gOQINVOUYk2Dm1U9Z+bLJwy
XNaUUYrDXQiikE3jWC76LJzlT4KTKni8kaEhE3oEHw78cJ3PLiZIEslvGX9K
ZEatl6u/zOYLDfawcaXLXWrcW6uHitQqD3qJ/1oJIpiFRxBxb7sJUMhkjrOW
9Wujo1rWT4oeeYT0y0SY28Zsr2eMZkRGfUfUtIrj/kaOdmBBNo3H3wkR2B4K
hCeqKXYgKfLe/vZ6SMHj3bIdWe0CwtKul6eAi7ufx6GYNmud3EL/96t88Jni
3mhMpUxHw04zGs8n9PrU7PDOiMJxn0mxbEggrksri8SIMWafmCqQSkMSarch
jkVCipdZA0aAyi87pIc2N3pNQDJ5cSmq19WTChsQkoQYrHWC96ykjBg7zgbZ
7cnWqjbCFFYdeI52SDVA5e4RVBYeuFIUwdaHbaHPIWEvPyp6U2jB+uwrvo8e
IUcZHltgoocBs1vWPHAgEV7gKHFFHt4+VkRFsM7AflmqGI/ACSQOZngbeXJX
qg9HtSssufxPWvcgmjauLfY13OySEchpn82Lr/Wq4bjyXq1EpzFe9/rI20C1
klHKg0zIl9t1qlTxco2QjoaGHbc4OjVfYdaadMjyGrs30OzaWk+CtZBm84EC
tnI91V5NV0det/McaLi3awIqUW6HyyEq7PIGtZF9pdsNIUwbqg3PjxjR9Psf
UJnFGVj9QJcTgPUByH+OBY3KrkwyDIpmpao9EKFKu+S1ik4CgH7B0sGQOaEw
p68qLhI0tliPBeNPx5lzjtlIMC1oa0j5fmY6ymAIk+jes93Ha/rVeNlfkwy1
/658rMnzL8P7aq2mPRItGWVIU9IEVdHdFuVLbKjKC85zXGvkAK+69bjjHoLb
Mh2g0H/qCQkLTYbRVi/fChXg6J4McqxVCg6T2q1RbbqjhkPtOdGX+Y1Pv7xJ
VXg+oXWwF60YI+nhsMr38F1hC4hQ412vVaj57cgqJivSm5q9YwoGAfq6fzlF
vzC24OJPl9xeC/5EH+ScdTN4glGHS3bgoTR932ZWyxo6Wnd1RWDtfsglUrP+
d7JsGeEAHaMigdWg1DFfBi1hzf11zLmKy+nOArYpsjV8oNwwDVTar+O7dgaZ
/egKgYlUJNk3ysZa5wPNT/xqrEvpYaQxTmPx1hoNBDFeo/QTrtH+z+et7abH
MebLqY6tDJr8HiIpNvONO936bJIeqyaNJCASOSWijRDGIzPlub5wEN5KE/qy
eZR+1dhAdW67SWwtpEvtNIRTjv//JYckobwbCkCenFhPD7rC4qIwCMNLawtN
fG+/60HD3RaARpzQw6Mrh/s5vt+h3+vfMduVm+8dWgPcRXcKMZptSAzpn/Fk
c3RTMGTPK5cqFxfDPPQepnDoSNFNLJjc+P8QaZdeTI5ZULReXIBF0gjjFYdP
B02AbUy0kzHfIhoycj1/c6SznZwZpR/eRl6txzqlSyCdJreeoMrhBaaX3lF3
G+z7poSCPANuypc2Fas5+ejbeN73GZn8GGgJHv5DAWex4AEPSCERjFpFnOgz
BS7GWH04EuLOZCW+J95WS52SpvbhbbyA7Dv5u3Vq0QaRT1ylJr/iRhWfr25Y
nv+bKc4hntqUgm7dy6bwC3oIsZK64qPPzbaLnh/18OozuFThPiAIW1J+A/fq
c5st1jBQqsM5jviwB2NsOGyJP324Knekcf8J+1t6TY9Z3HTr9yxoitHT2ea6
lY9zJrI3G+FSpNtJXLgcRuiSYAhwNC/BjnMLiyt2A4M2YQ5lDj2lt1fwVVTE
RyQkWujWGShQy+tBtWbRclVjsZU08ZEhWYxjs9VSY/VbuzavWu2Vao/TJqPM
JNJdK+A6iX1aSPpQbodbu14LWuXJMinX7cKCEGczhYje6KMaDHzK8UcL3KxY
NDwGfHpfQqzazOnydqhL3dc7oGNmbphbVqSjZu9OoCo0MIAvWgJjA58gkLbo
DSkZlTt4s/fe79vzuB68MtC7PqM2JPWNbijxzX+rN2DnV3iwNcEK9nKAIZsz
+gCNMuSY/kxqLjOLNBW3bPQlyq1bcUTo6m4jKLOPW7Efd1K+sfDQocYJfa6e
e45ILB9+th7HoKmSatyYCVUIfZdEz40E9jPjoKyZ8N0LAY9huD6EDctqGKmM
YpcAddw+9pWUUTMko7njaAbk4zgU88RncgZszvytGga5vSZq8gDCpVttWj+i
A7XwTOelSHBqj0PwrnlEjsi0A2v2H0owgOKwj5H6VzvnEYBJZ3hePH0CUB4o
4dfR9YVqeVkptQ+Rh5By8p/Y0R2+Sp7lG6UIeCk0BqPXqcSmTUdYgZ3gjbHn
Cbqv/X4bXnJeaSpHAYA4lqpN6HsLjou93yeGMaB1EY9rq65mL5J2phECgoNk
QF8BNrOiqHWiOBMwmkg26QvP/tc2B7Hhr9b7uCxkXNeWDouPp3Amv69HlUjp
qGI201C/nQVJCRipY6ImIoWKPfm+DGbCPKFzUpjt+PYUYMZLEZ7wWC3UIHUR
9ULRLlgf5rhPKXkFSYDZY+B27oBgYToo2EiLY2Kw4MVyQ5fSzOTnXQZBmDS3
TKPkbhty7mLvoTK10vlqx7iQm+5ycNPZ8ZdSiONB4lgoVeYI5s6zOwQb3HzO
DAjBHIp0E9/aozz6WS3YoVj2EQIfFjPDMnVCYjs1nujb6uYHfuLitqGwxhpA
/JCR5aewVVwHUd07do8USuNOeyPEka9W71G4ScZd/coXSxzybZqsGZ9tKnMf
k+XLxFIu1AvPV0NxC0Zx7WlA74/IZjEi1rZ/dUD9tYy/OlJ552fBHl4mEDzJ
moHA41a/hG4KR+vpP93Bbn562q0VUTWgtxUJT1z7HIuqaLcOhonzfis9lMWW
ItIHiW6pJrMrvRZIoRGGF0yQoss/bUzJJTZ1G0jAA1FCyP4RzEZ0c7na7ZM3
eWnvbE8puqPnBAzBecJAHSRSMCfTqc/MNnyt0gnuX1iijjlu5Vn3BRTEfGpH
mZVZoeqkvSZXH2p4S9CBwrfb97l7hWLewQz0vNaL4cIdQjXtl0w/e3HIZCAL
rhDi/fltxjescPoTMKE17wnFIhAn8+ONhN/S0XMKAALGodxZuMmW1hm877eg
+HwPTWuDGq6BzWvYhW53KoFnC4IUceWhUvMdCJbJgGpU23L+S4MucZygV3ha
EjTvzJx+TdTcfdJ5r0Bs0QJcHjyk+kZxz+CwMDugP4DAnScoFwFeCQZbKSw1
/+MY+JFOGFK/N5sxwewywQYxo0tatGzfwJzFtl0Qp/yEfbGwPWtGFOqaYtnk
TO68DeffQJ0SeTvqhMwgWRfExqayZoypqkxdKvwDXEH/Mx37Kn/5sqwk5PAI
E7NgsqEtt2PUUKNdpagkjnNNEBHofZcJGF/M0SsqZ1XwxczOQl9BGE1NWsjR
TvG1ZY1y9eBFEvHytN4L8hTGsRURvUYBuQhCPurpal2WlywIULn8BW5DS4ys
uNBK3tS2lBRVJSTRJAJ8beMdUwzIZTnhTiXj1I7LmMQZVE7mN6QH7kH9sn1r
xbGSCUv0NEASnnz1iZ0MInqseeVK0P6zOrBSM3mYpBiATiLa8G4ftKJoxHKo
KF80GXIB1ebUG6hVoLW53uouEem3PB4SAxcRYjlLwKETtGB/ZiBK3p5Px6zp
lBKDJ7goFOgTZukbd2Qtb78YrZUb0QMTUWRhWfq8Tsu2X4I3Cvn47Dslh1JP
D0bbfIH7fxCQTz3auAN0TEqlMnVTYFEg8feFBGOIp7ZcA2Pzzx0NYJxtHjYp
J601VKQJRrlTkQ7azvzMBoD5vVzpdVpT6MtaYABFZrNr43VglNbF2ddygc+v
81YN40Nv4io/5njuk4Iy9DDePMqE5HtQwJvHA+TIjfjAQUI1yeZdz3H2BvkL
CwsBWT3klDsEQ23LQOLmh+xZ4DHz7vgyevnWCHTJXwhiimH2FG1oYzi60xXT
wwLPPYQKzJq1JDh1pI8Yy5auf4wgmF+DRx6OztxwqqqxAw30No7Qd+xWgzkA
I9sE9pjxWCSt0+3HNcrMmqp9tvxwKSCADzHSjI8ltL/p95Lrv5kPNPpgu3N0
HmkgYduq7394da9zWsybf9NLeiw9xxQAmVfL8KOr18iKbFjDwxSIx9L6uzht
dRpKPslDUOpVfmK8WioKhb5ejmpbAM5UIyekdxSxOTdPPxOdbfc9fvZlJxwV
uikevTd7f4wTmag/L1Vgx2cmvGf6c9d17IhOwMYPBijKIVvwIgaCPxvZapob
s0BjU52vKpujZWM/tnezt7DkDp3Jhm6ke4zqW+ErjMV7aGqT52xr7IJ+awum
tJGGy4i+zhCs7MJYZVypXzPnXBZGjMAkWkme3VkdWgiYaFyIJmu1IN/iqT9s
Lm3dWGs6SE4qW90ifQqKiJkQn/TizyCIJpLXs0Yu8aFig1pas1yChp5nMQ+k
raYHCzkHVQdashAb4c4wBBqngXCb2DFMZpywUsHLr/i4mc01AHNva3WBVB26
NFCMcNhoEvHde+AlAmgDBrmKekOktDkwUlYE6XB95T4lQgRN3Oa7uXji5Z56
Pl3X9LWrYhp9NQeqg7dDUZi8lKIJ2a8d+N3HD+Hx4kLcYYJ4W+F2imU2SE90
+Fs/tEPAnvpIT1F+MJpZg03vDHwE9bJb+TBKU08J17j/CI+tmjxZUWVYFlD5
sKMrslFbyRQ3jerHRrHpm3iMj0+Ujhix+zcMaLfphIzKVBIV18OMhfsoCyqz
qdziKbJ/0VzbXRVS4BuesEbNKre8ogNIJiC+01jCAKC4uL60lMYvxxamEVv+
CDcsDms9UwlysiwzfpvOYXtWblth6d2ewff7uNOy/lG6MC4Xi0HxCREf1XbX
378Cof+HzRd1hcr+0JnxdAgP99db4nZEU5RIf5WsCpHe/oc7s+x4bvyWqcj8
GBUhO2j538ZIxmZOmy93hhavkGecoN38Is9mxmRErtr/jaFnAf7ClpGIP2fD
C7RT6l2YOUWeKN38+R0PKqag4BRJ7mw9LGOvVsRyp9OTbAup2cnfXj7QoAAZ
Q0bR+kxN2rvblbbt9u7Ghuy+WeNRnev094qSLYHWO7nLvCYUF+8OgjgZNH8K
JGwNX/krrYkLJuJUYdODlzPFI0NveA2tBAYBcRXkhuF+dKIeA4q4EQGC7Hd6
UwJj7XL0vAFW3VHTlyInaRktyPZ2h3gw8yE+56TFMu6ha9YCyWtQeOhWvpgI
GPQ8hMbhlPLAWEiJu0SZth2Y/mKrHmJ+c6b3fbG+NQqx4FdTskU1NlKZjCXB
BJf7QhnktCeHApkSTvp+IITULidisRaNz6ELqsi+IoBMZ/cuQPy8B7FPpKmc
IOhnftespO0Sqmdror/w1b81ChikVnlgxqrWHu8AZfWlHR/RCvbrFjt7wAaf
yIddgkLHZfovtnMVpcpKguI3aL0Wuma5oeO2TkuoWQw4y1fy9zt6Xd1zM2Wc
JjJ25pwnalj4qG9h8lk2IZhM2wlvYs0IDgfcSLB+TSudNOJjhL/cprcE3DHr
pqFfxnYJkL00Zwkohre8vv5JSVJeVPKb9ado7ZEcmT1Ver+VrwxsdkvY9qEo
BZBOEYeX+13N0hi6U9EBl+tWCJVtf11Di1YMwP31x+agm+DxH8lPyJwXZwbv
i3JAIj2p6G31RNQw33+HlJbOv51iJE6qjuEZy42+r2Xw/wrR7cAANZILRCt2
uj2b9pQd5Lu6z2DHbOLTrAdILsbXhzEPBtWRcM8Ms91TtdIhJ8Zzq4Ga+4rq
GswqauL13BUq+tIvTAnRw0I5sxvoM4IpM5Y5CrP3qA1YQ5XzHhkQn22bzGh4
n0e4aVAzGpYQPRlPhSZ0bnMaj3Ww0xE3h/2yDNZu4CSnKBjLQW7Qj169K3W8
ELfdwlfrKEOzyTVQq+RQygkwiq7SDr3H48xe9nQ2VQFF0bFjoewRoFu0yL9A
IrM/GUeeXPS1YyKxgy0gyiwl+UuncpaaOBhKZVDcpgwSvqHeS9AXGsOb9w6G
uP3n5L+D5e8FdU6T1RT05rcYtbHQuByDyBZ4zqQCKQndHsHGj5zDt9DeyUpP
RBMXYk9erNnyG3nIA/uFoHoGAXChRytObf7ik2X3+6xcSFK+aCXUifWKWZBg
3sJAue6mtcbvO+LPpdcgo2M3vDUCpwhcEWN11Lpe2AVu9c9Mw8QjgKoqIjZj
5VuvTmL6wZg0QYMIbJ4jmVOr8Ah6GgU+wZSyNIwJiX0p+qK63Hiosiy6PkvA
ABm7IFx3mQDlBbFuN83ZKqvZusdwDXbwUK5ZETYMcBKo0dZV7jeZApSdgqkS
u0DykSGbJQx2OsMQS7Dyv7/KdpHileTAsxfIhzIuLRzVPkLSbIleHsxurz/9
ET5dafYNCe8SCUL1jCj8b4GA5J+woWyhEc3Ppwaz1S7x2XCQNaSr/wqquH6f
o6R6HaNQAOBgfaKI5DDdyoNXgUZ82eGVhdAtY8iomeRWSP3boLX4GguMJsY9
FQvgkqCRH5iVHigehx88b9U0pimJDBWJbkvm6vpZnSjNnS+a6cklS9FyfLuC
0Mc2+07OWUUurr1NFLlociue+OY+Ty4qTEl6qW0xkAiHJRV7JgQx4mWEnL6x
gLYq+pZztkgYsiVIHm1iCyV0C5IUd6YRl+eHEbt73FW8qCcfp8EeD8Mbs3YG
UWNeDXkvsfFIK+zTfE7Z50c3FD5MhmJyo7Wfj1ucAEqckhHY9dQbnfS3ujP1
XlfKF9wouyaQ8+1CWP0qlj3GEGMAlfUIaUpF09hcl0d31yGYe6zzHUe6f+/S
VQaUTGYgE/u1p/DdYmB58ZdnfkBxfXZeyVzDwByCSIbuczR5Qj4HMTYkKP+i
NKU5s4p504v+8TdjoXZmLlwHtNp0rruFNIk5dP+802BvxaZAra0YpXehlQu6
JFegufAUNWIqcRCIBCAkFm9vsHdJl+1e2f7YHNkpj+W65RCgHRRFQ4qBqSw8
h49pvSRYHbvO5IilZV0ZqTbbvKOdKBPo2NKGm6dTgNxqnnq5cgU9oi6DqfUA
fG1LYd7kaRiJhmbCZbh49eFEyssOYMBD4gGfbOlxc9kvPmtMRTM0JBOBZ/XZ
vt+Z9kNap6uNyMATEpsrbXQ1JyCrPx5Ngh+vUwC9lE5t4NQDRtTZu5GJu662
BLodhPq6ZSuYkSlcBp6eIby0/Ez3jxpbC4S+Mr8tQGoHMge83+4zNqwhL1mr
RGn7urT40UtAf+uCsT3hQlJSHahI+1S9Qk9EmaHiVrK+lZ84QhgH03pC/qzL
Ayvj852JDrCsFVvLf0IXppomx8VX8NETXmCtgbKTP3d7ZphCn62mo8CukMii
pYhTjNCp6zvdP0vZaS/nlG6fO52KeuyGcg/u0r6eNP8v5QEzsFH2ba3Qjpuz
yonsvQqDqyO1o+oCeJ9MBYmOHAQDRCugEekOpuP1qAh2Rto8GY2i1rycadgS
h7YFGhJpGZoxmIVgkpcdOVrbP3kz/0OzVjodkp35p2L5STytKYEZnTr5sonB
RyyA6puGRPE+hi7tGLlnvtwvWlyPT1jBrIO315bXlz3DyPZmqVB9kdp9eXqX
6wEG67mPpkHAXzJNFVwjIfrJGglMYVC6e5Rm+LbnPL3Q3k7b72cTE/FkH91h
aSCB7kVeFfXE1LLx/Cj9R/nLFsRuvhjMwFIhhn++1TpHyBcknwuRDATulbCm
gy++RY0BgYUj+uxs+KOMNnoOjHwbzbAlE3yhXnQ+s7qjQ1EapZ/F87UybYRo
Wrs11VMUyAIEIxsu6CPh8Ec5RIwTHfB0aTwwld+EYtGqXkO+UwlN7blmbLMo
lgL0gKIsfZJfWVxGXfRTNYRVUa66xmM8xdm5rSrI9rTO7hjyK9TqVv7fjZcr
X4VZPQfWj3/TrtFkq8B74g+0/cOm8/LQMzAF3B/AjzlLmbKul+ZBuzD47aE8
KJKZpp1vJc3CM1fP7gEZn4VMjevlu+koJCJt8/t7pAcp8vcnmhM446SWkRjM
nFZzQ2bIIk5JuqfT3dZJXYPjd3dkIpqy7GXlBr90nMe9cTicGIermvP2/7lv
JIODt8ASWzAA386YYGS+3Qglqi1El6hwZc+rnfBpAJFbFNcy9tOeVYlbGiOZ
IG6hTRiYEyfLD9SI1niU6q4vzGAw+IQ4gLN0FEO2r5BCA7M1834YytcHoJIY
Wurwmaz/+YRsyOQtdyr6anRM47wjdIHq2MRsW2cA32EsyAmwsuJLzGZyST8x
MB4makrFYM0zT2sT6xWQbOXN3jb2KnB4YJWsVZk2Q7SGO2Wr0bI9iqPhsexi
SU8eyK3HmwEyxawzuATBZY/blYeBMCXr0IgiEEORlJlPPpSSj5TDnnVD8E6I
WeJiO3JPutAKt87IQFeJIJrCVf43YOVOcJ0KWv4LODoIuz2G1HNEfVYrOAL+
JToGekjFMQV8pGthhPjdmhJH9s8xdqAk5DEXocS6Tcd3TaLUhUYdU0h7wwAu
/KkwIZoIQqROVOrPG+QHFP4CG8NlEjaK3g01Nbm/T4NhhKV7nABIFvzhnpcB
OYRmo84bSPXZ+0OQPVi7y+2UMJ3Tez5PeESGxsLslOaJ6Zvf0aGv2ozEdZqw
BqEXZa0p7b+pfl2vLoNrd0jiMitZ1wg200sy7NWrUC/Kr/kP9Jbq+VM0qWrO
U53DsXITNnWJdJ7OXXckQRquORJ+CwNGMqmyBxvApxe4WiG2KIqEb2Ln7ZAE
iCrAWZIA/h9pgBEicd31Pi2wOV00sBHmHdzBREEkoEx3+ecLQAvWr5LQT3AH
Ev1EsUOeKeGVpL+4PScrjc9GoQyDEzCBbiMShV7KNrx3x9n4btCzxfmFQ7kJ
fsBZ0UK22WR9XswXoM0oN6cZXOovCAJ3XzAZ7NH5tz9gMwrlXsy6ii0qLWgR
39G8TbijHYSQ8LxhyQU2tGud3yeY0hQeiSRIsZq5ndODz1oqFixGjCV6VbYA
jF/R2ST9zZWE4q1ToSdU+TA75Z/DyCCZAnC7wgLr/LpmHsJRdj9HjY3INWgF
TZEy2xV3vF9GrJBrviTcVQiyHl5bA3gRPeG4mNb3aF6wMMPPJWrDUdoLawvU
OSXuySJBkH4FrcliCcdmVPclZfkx1Ti655goBo5rsP+S0SSWmU7tDbXRvF5a
UnJKcSKgBUN0m7ue+KXWXboO1TiJYO08XTjweSNXurepKNfQuNqpk8uj4f1O
94B0KKQSBboSBQgytq96hy9+As4hgj7z68kuMue8yX2ONIrd9lxgR9XvKJtz
5ZMnrulngMQ1QUuVzRoRi0pOyryHV3N0ZHU0tJVl4JBXIpqzertVI8cgcheE
0PTH9DEO4In85GG6EkYLa1pjaj5BUGooZ/b9xfi7zHhCgI+G3stMy6u6uDsI
MP06J/Mur9p8cKqlkxwF8VzOoC6ZsyupoHXPDBry3I7Vrkpsqupvi7PQ13OM
FJ0xvypt/qmPEbOZULf3aNz7FEHeNK3WuvqJ6Mmita8gCNtZhF7RdgDSxzL5
47QLJE9Vox1zx2DkJ67lB7Ghlt+kkhgnNsT/83AH4in568shc9aE9c7+/Kwz
xUwQGkOSKWXcaeXUBYdsBcIYz5XqAP05GNgKkTMwbVPUI3hc4Mk/DimaIzCc
/yIGSa0xcFDainhpl/QALro89q08f0wuvPiQZHdJeHMW4APiFUPDpqst7qOO
InE1l0ZnuWaKlApzdy4kmPmPbJQDfCBp4LxxWViAvs7y/F/4fPYaU0KIqnRr
Vx/X1JE4H6mUV5AC7/jl7B9r+hntNkDvUeXiR3FsdfPc16pP5rcr3qC6xWFN
8z7XYfiFOZGPIBhP1wG+rbCrDxrKDJ16LGlt8aCFcmdOOtePAclvLH34VUTl
9DbUKTUwIjQjeON722e5socIGAWvOsBvGWmAvBxEfN9DdZOCg7y3xeX2O9lw
cqBQu19w+I9OSOFMBng4Y4RgwEjmvKQUhd+t9h7UsSHq2tCiEyV10idDLpu1
HwMIflzi8KmqrQ6ZwHY71lXzJXA4epLngCnis0wz9lAPfN+SFhiw3CDds6+P
jyRKFjksDvsqlJH8PEUyDsTAUh0P5Xsux6Ld/7RCFbCooIfhBeHxD5g2pgSE
WZLMgXY/+9IXe2rGiDi2JpBUrZi4LiINopTs7dXCmbWSnJBphqWDYkkirhMf
wCoeQ3xyfGBbSkBb3j+R/it+/7gy8+zJ4PVtWSbIuev2iklGgdWnn2H/uBDY
XCSJOxCJj5HqSHtemdMe/81aAV6mcwKoWmRk1n9zWgAl1CAr9akKdBL9EXZO
+3ZLbGIahjhGmSYAt6uop4hq5Wa1RSAlViiTCR46pYSClmnOWyhiQN6VFE2/
Tj0ZkavE1neoGStPMTO+yf5y1Td5UrXQwPoK8X+JyEs0hu9p5g0ZYsBJ2X0x
xvT9ptULvkq+3q/2hhHkAfKYbGfqIUTV1nur/qLnA3SKMYRBsrZH/gpwPce0
szWvhoge9HUfc+0dINThZjMW1/jxJEX6H2MYbYiXxNjQPzezysgEuMmY2oE8
5zqcdtVJsIuLINigwmlsyNzSXSr+3JKPj707bs+Xt3EydZq7jLu3I3xrnR6E
HyrOSUt4C0rFZKqfrHXtVD+DbByUzDYL/EI1tvvZP77HCvBVMjjD02MzSLCt
QgnGXrmvpcdc9EpPVgolIZ6sIIhJ9erXMqfRipMY1v1EcbOvb38Svk+hDY3y
8x04mqKjFX7lW5BrWmobQgAg2eTgJiBvmy+lT+iHbEKZx+4M70KI9+zTCdJ/
5LYB/sRcq8Tc8R3tY8MxbCMKAsTHjwek+BW6FzDYo7+gHCv6Et4mmKwl+oC8
IYsF+RIKvIKNGnImZ20Ne3lmNEnhlnXGEcOZ6bXR784NXOpeTb/H6WmZoXo2
9lqMgB4mfZ76L4KjXa1Vvpz3NA11DWBIWdpQH+7DA0TMN9zx7RkESt5zLwaF
MwbFsPyj3bpVTLAOsFbfLCfewGvAZ8d+fAJtbfpcO9s0OKRfD8KC7DYklvh+
ttnWxdETE3bPIUh5BLfW2w0bxTmxiyaDAOen1g+E/260gIyhekIMrWRixdAI
Kwqgck2I8/OqaiVbPc24/Eiz9qfsrllj7TkSN15DfZq8UBcJ9k8RPZrQM3/y
cPWW/Q4M6pJTx2Sl+6h3w2KuzmyTD2Vt9IlnB4/XKLvTlIcVEI7Nxhh7Fnp8
PcnsMm6acgww1q5SuWibEyIoI1dUlfbLQ+wuyIXhiXzrAmJ+ijqXMkedZbef
le1tmMY5MUkJWKFxJa8Wa8kiC9S4n70IUrqBLESzQl3BglTYuWJQF8OJ9uVx
KQIDtpnlCAdTUq9L0oEPxAhPwyuNBBafrHkqiO5P3TfFtB+easeqmGf3s5j0
z6kBjIBXSrMtWmxCFFly30jl3e1L80cYbR5AX5t8RZcOi5SQpA42sLxVTg5W
/UhwGeC/ixVq/2tv2hlnxQhLMjpsHVU3xokc411GIZ0ube9+mUtYLmAePqYh
RWrx/Z6jqwwIjEYKIxvU4ooJ314O7ZmcKlDSAM49AzrpWo6gagYOvpsv0Ja8
2GPYdiAkyIOJ7kmp1v6x0jMgQaOFtA7efoE5LYKzynGEoQ7agcV4aprbLxI7
ahrrFjuQlkM7HrdgZ25g8lBHuGs/qr6DU9aDzISyWKWAa3VbPyo0wT9b2ErH
AwJcJXJbBMBLE40akiK9h1QYRlptdBkBU5Of4GEB3Vw6nw/coPfJ/bWeDAUb
Q9QcmqD4apfdsUiplFcsintDCC0DSi29rOquHzYXpFVRoVzz7ae1YpBomK+5
/2XpKDzP/CfNk+hHyJDiGmItIXm8jo4cHTpd+E12nam29XLO15lBaI2H+qWY
XpAG6AUUDiqtsd47pUTrYosBp+XFIowsTB0xkqYaRm8KYMtGuXBHhV9tj3dx
uuccW3uKMcwxxaROSLhRyrtp4CPjnpnB1LXfjCgObofqY+w+mvUwQtTe6Vaq
6XwfZTlqfJU0mnUePPQNjbWBwV3erKcijAna46ytmAF3mTApw5HaAwQYehZI
IxpR49XTEEsZ8u5hERi1Cig2vRLkbC2nJcUpRG3BTAwT1KUk4jUIbBpDaQK6
AysL2fiIX0w6uTQJkcETICftcDTQ4lXNz92E1PHxY+ciuz/KSv7HO3Z0Pz+2
9zyYS53egO4PREro7CEpaArLVf3jXncP5f05kP80hda6i4AJ0z95n2zNwqkt
/ChNSooQliLDvFPRKZ8PCDCYj7o8H26TSv26YjS1P6cZ9sDSdObslwiD0wFb
yGY3zU9QDvHsFEcIw/hvbRBFhgVlfvngKss2n8FjIfKO/1Ct5qpU6p3OYE/n
fXEQ9bTiWGsqggm4rDDQB3ILIqppebXsCyFazWE7HPx9PjKWwGViyu49McCB
cgiHcOVg3CUUeq7mHqKNm4SzHTKKrlBNdF2+sKT/3HRzeUtrg/EHBBiV6ELk
IGT0crOU1blfdY3v0oE4ae08FViGj1sHk23T6TWvhTkFo8VlMTbJqZCMWg4u
ZJDGZa7VRGFM0R9PkuRmIAuF/LMnJFbej4wMekAF7T4aqrOd/y/yKMwzgRBY
h+MLa9IcBMD6v/loLtthWZnitCuqQHOaS3BKOmteHrJFGpTa2UmnIxc0HQp3
YXEz7ot12wfsVdABeFJYnTc//r3upyh16+DYV3PQMLeJwdUeJXahbKZw6fQK
wZEZtly3SA4ba1YOjCMWNsAfmJsXEWSKOBkWLKMUC2Hb3QZpZCyUxFTNn4he
ArrCZiJAI7XkILG77bM4XqqoTFa0FR80+2+2yaLjGVp70s4KuVXkF3Ai5Elq
XAmNvniS32EQsr8E/QrIJixVutFgR8fqf6V1Zyact6oncCAhQv/WauXrNN+3
CJnB7mD9L3XZr4uineb8VxZh1X0LQ5lfeurJAtKVx/6FcYHINgU3RHpw59qZ
eTwTbFGXMafYCzioadw/5i2Vkpvf7AGC/zXuzFqJ3hQPad+awg110DzY8Cpx
1c6JR34Smet8JEEgsibFOHshtEakE4ucQA+HnHZSUmyxrB7yRfxciRBvgOGS
xLSwrDAZSGWuADE4lhZClDGo9CJwV662NjQKPCksWh0HfaHIvbCXrv76leVq
ZEG7aZMvyUOdA/T7+T21j2BksMCvSPZGThYEFan0avOfyBbTSxLD627yknOz
qG2b03b42U9kWgIUrCGjKNE1CbxPV4nfvXSQtx9wX/8EyPHaLLN0x1YJCJyx
ojJ1c5c6oGqY4rB28/Rgnc1EBSnsR/MsTuZHIAmOw10KggFDecppo19h1c8a
eHqfk/BTQRRunhFTWn2+FQt0q9SRdUlKQAWOzSvD5jF9Ps+5p/cOsOlQihTR
vN7x+z5vnbrrvGUOI9rEMfG0nad5/fjL3SCyNuLtma0e8aTTQUOycNROMQ97
SKPJbrMMTzZUcq/qPhNZPkEHEMC1Xo0Emtm1BJRxQh8l02Qv4/b5BGCtDc19
6mgAifb6ANIto8W39cc3msDjSXoxqj734RL9t3z8e/OyNHx1GFXSiotSV6za
OBT3HpnrtqBcQO9q16dLkrUFblQvKCyEMemHVID2zDza0iSH7UdZLuPAYMLO
mQNmLqDVHHlBcoEAZLOBxrRfA+lui8IKncyEpB7c96dId0DABOGt+xmS90Uu
H2PsnQxpqUm3zVKJa2N5UkJSJqEmR+nUg/xiRZeyJwpJY24FP+dBnRrmzPF6
rPlOoXj8aVsRzWVIdRagQ4vPe9eXtu84tDr+RHniLiyrLceCkH2k1iP4ysuC
syzIXrvDD20OL+N1EGco3EVYOYtJ6xdGryKGqRnurHCdqBceJrow+WXBSCVV
JIXSZVxbW2WRCeelNn8d+mfViYg6HiNK9apJswPItJkN5WdhIH4FqLt4SaKk
IhEfh2vUOwrTh6ulVBiH4WS6K1CCueZAu7eRaLbrafRp+Q6x/hkEx5lLDEUv
mX3431brkDgf3JFwVFUsUdAUh831ocy3oTM5OARjzQVQ7zVWOycGDUz+DmqL
Njure0JoYvCcC544Y93nr0PYLG4cX2z0T9+PN+KW54nijgDoBqeaN1Nv4duv
GfcAZZwggxf6UQup4l4ybQ0ly8McDoAf32kCrIoNHZGMdFKG3e/CgnyGymKa
/7/PUwE8qh0gu0PgI/LLN+MZ4GcBxwXagaWHK6o3blyqV9utjSy0C+puZI8L
BtMBguv1hkmGRu3wrfv4uBmuDVe4Q2tPmvqkbDskchgCmWg/eBmapHDTklzk
lvuJIPu5Xi6+9AtPtd6wcmYIfFzlRt2XsarJIRa6FHl/8ZBq3nijSqxntMmf
etJbXIx+KGbSGtikqm1lNtreXwEB6ebVKVgzxhAHC4sHjVCrhPPlnjhcc4mi
ONG5z+8Xl1wC55+eeeDDOyEBJcIe0Kzo0qJvKipDe1vUBpmbEFiNMfWkR1Nz
3vl06vwugepFSnjdzBiTVkqKW6Px8Rtt4U7CzJB3w70WmVFLqEIh3s5L5Y8Q
Kj280i3JeiRMGnNaQW3SMR2Ptc9vKCp7XdEePmHl2a6L339jOmcdzjnZ01kD
bitatHxeb7HVGdnFQkfVUCGoehEDM2czikbf80eMeIi3+a0/QK4/0JI4Wd1I
yos7tYTP1UCUnDSa9XeQtJwvg2cagpgibJFvV/WGzL1iob7cdKuGLCwjN3RN
EssPsERQkQjW76PIxjipMSgHm0VJm5jxU7egGxhOQlflRK39Ntw6Ot+AYc3m
yMe0GV7VOmmD4hgJvbg4k4yGyNeoBEt1pZXa+A6KWMrJRWb9qpKOPrNLx9AK
lmmN9tAWyVFwCFf6lhfSDhnV8FGqacbMZqt51xO0H/dEsMAJw0EF52wkx/ff
xUH4avMOrOFhgDNB488XSb4wf9/mmdxNpGEFgvaM9wksrb5hK7s5WBx976PN
x+RMirS0rDd98Iu1Gfx1pdAbTMJ0dp1JkiWeZd4m55pLOy2u9e2eLDIi/GUc
pH9ewvliJMmGW5/+KOoWXzLhwBHzlpyF+SOWh6ZV2QGdG7R4XxuJkhzK4SGF
kc12G0IJNZ3nwyvvwgxtO95P+f8T0e2jD08mMj3M+9R1/isx8QcBopCgYZkJ
geD5laZWEc8tQUtlMNNy/AmCxDdluL5fRXteag5tHxwubk3kpd1sxVaaSgMj
jIB+jbEFRgmmBuxg+uJDVVXTJqwa+CMcLVdRO815VT6AIF9Biv+bwyVH8Ke6
6B47JNsUl986/f8Dgl7aXkYF4rS7gE5z6ktlraGdZyoxW17mKWzxF6LhRGcr
IA415UTW0+/7eSCizVSSxIaLvTUI+bMCWji7b3eDLa/bz450T8N6oA2N2wu6
9U/k/IAFnsghSuTgcQYcqG/KSTV4XOBL+UESiYznUM5huEKTts1NnESKQJjS
iSF5kTOYmXS+0abPpqsabPA7JXV8Rufw8ric2r9wCYtbKYERCb12r/uAOyMW
D++xqKQb9IbhhPfxgh5ePdfhO6itHrrJzSEI1PdfaWMgEYJJQmoeCZEPJJ2I
OOV1MK0sgjAg3v/yY/4jPWTMXktstrB1ptvlk47w74SakMHyTK90y0Z1h65b
SUVnK7+7xkbbweWxDjJhKvtDYQ46tBOvuw8MgQUAio6FxQBh0hgIjVx+0aLo
ZgrDBx5k2sFi5dvuU9Ys7JrXYDcuzZlha8LMrEulQR/zRrB4L8qyjapbPuz4
3Uga9BqxGRXk8h13a+F71QfctNZybjnjkrqHbMskyEfDCfpotV9SndA0Wuet
fIQX9/XYrm1dkx4oiGjRB9ErEtIMlmu0E+kQFvjvU1qR+lkvZ60PD/fG9uE9
rZFVbwPFwZSL0SiSOKz9USyiiMqlM3S91gOiT0/Q053NVubgONgC9+cKUu3L
KrDhCOyd4aNesV6irzSXxHb3awdyXQy6pI17zSdVsXxDykCwF2uhBc5adtHu
6botrsR7DQTcZE/wLDy1j/DMxCQzAf9QRbmV5MRKQKbVmQNbGY5/V3H840dn
Xj4qABcsm3rmLc0eDJw4a/Xs7HMOgVQ7uG37teKH253y49oxzd4HgTJPu75f
1+LFqL2Ud7v+2MwTYKkKSUTQMdtDjBvIuq4DCA5j9kCMMlz/MDAIirWzZUgd
mGjy1cK+Sz5HmjFlukKKSpEpwRuWA2edzQXkv3k39YaWfQL7i0qXFMx/IFls
ra1gCAq0mEjIPA6UAmxtT/D7y2u/b9WM0T+BfO5Q0pebSvgxqiFOaCGRxFi/
oUq+oF5HM7b7vfAhB146P+sHFs96a4+vB1VP+0TfOHEbAUjMS6IcZE9wMs4I
BSer3D52GuQCBm2T/dqJDa8+zmDKW1MOz072utV80Xhet0uHD0t90X65eR3T
HLCirMd354iEPa9QCgWVQKsdMXmqiPzJWmKUlC87NCj5njaLbOSf+r8Cuwv1
sJ37sSCYGW90qYEvH9SAtL/WwqKBI2lUyAjv8SV/OzI9f85j33Dl0LwNT2iH
OU/Nowz1Gnff75qChx6fBn9yIV+EXGFoIT81KeiDKbW1Lm17udOg3mjAc8jB
uTtDv9DVkYIe8NZLqA4r4j99OUGon7zCvJpmNw86fseqss6mmLe/qFsmZ320
o/yT7i/Vd5gP1FpWSmSiB/vJivFb1dYoGCq7uAzTbJhUiKHukwDiJXZgXHGp
AdS/fwoanZPOh55Acs8LEai/L6MM8zOFE30SfQcX6CjXsBgs1HlWN8I3hBFy
lAA9ybLCObeqNesBWu4JOJsmUxHZcr555ildirrDWEVTS2gdD3KZuyy+1J6p
/zCDFLxJNWmvck3UL5xDt1p4Tf56Pa3P4nE62AzvVxtRBr6d9+7UU52UxI7z
+bSPnW7UGyozTXyOePNBtOGUmsIbd4ARYBe0mKjmJjgD6TEigy402PQNpMSh
A7tomUfNWhnpALNiEXc5ZfjS9hiWLpwjsyEGgkzBQlPDKPPQ6HoxeaJH3Tl7
ALcahqdGdF/Fq0f/LpsQBjoVkwoZ65lEN4QZQK5HfNeGKKuBH9SLmneauv4N
OLxUGQvCgg/Jto95rXCV7pH10lTFYSS7OCoX60RWS+m4RJ0+OZ4csTmGn11K
wehFSvMV0Z+74cuPRhMd40cYfKAYlvXEVMOHaao5o7RVgvimGl1zO1kPAsYr
TB8DWHATjskJdUmgBeC1muwfknkVPnxAc0nWcAk12+tIdZJFurVTZCwcJGk4
JtR31IOAUJKV5R5vSlbw/AdXmkZflWmLwNwls2BwQBlSPDkSilPyeGlAQVVL
8PDRV7taI8tPwYMhz5+AorByG1e2nbbXKozun1CKkw87MToghwbgMUjfnuFw
FSAWe1HZKNBSoGjEl6A7ipxPUmO7hjQecSB1rr4aTzHyKs+QK+bd6wsStlQo
WG9d1HJyvSpPLlyWQ+cZG94vhVGqMgA7g4urWmm50I+J7IvA40tsrFY3BocU
u0LdIzv/g+nLZ6YdbbX9kgnwNgnRh3vvkMvkTeO6UR7k7ShTENE0o2ER4Ehi
g+mfa7YpnrSU2QH8JKCVAR5ly/rC/UIypOyn3hG8ux7SxM/Ujjx8qiV7BCVU
z+AJvcnjPGhq8ynOsR5uMONitNI7EpfEFQMO+lEhx8ZofRefedjznsj9+iCF
qLr5T/SUCQaz11zZNUsAzSx/SegELtcAa590bRSKX29BtKx4DwveznR1Ox6k
q/LkujGrJBMFkrI/ruRGzDYaEmOLvmyBHjWD7CMA8+YI5gp/4VAtEpAoJTyU
FNjNAnvvlutIVJX6SNA5ylW99iSmvXI6S/9D8Rb75RIKNJm5fffQratdErgb
MZij+aly4sD9vvSLztyy0vv6q0CIdlXK1ZWU0ZmHTXnrx+Mtj6mXFkRJ1mnw
jjgmNIUbERbKXrXWXIXOdlp4pAWqwhoBg4tYehK7RjxmA3wdOxmY9uFvdUYn
31vsmxkcK0glvbPyny6QBc9tRw5ftXU/IU55WNnTOePblSr2GM8IwzfS8gdh
UROEn7l/FDVmYpJHqzeHg5XzBWQ98AmviV7YQxiFiIijHUooPwJG8FwL0/YW
Iu1uz1svdpC19zSsnlEXjC4Fl64/vsJlH7iKopKDrkzqJVL8FgMfTvL0z/8M
dnR7YB6Wz5IslUzqBhV68jmIaYHdS5ZYrVXPNKeQs1UeOsAQoIO6fWERe84u
UgXysLsmwkL8Usb798HbQzXZNxEsqs9vwnfYPn/k6puQS3sL6z4gwqrenb90
IvJGWeloyraeSAVr8BdKUSydm8fsJxXs31xWhfEAddwFCD4HL58OuocLMTJD
hLSeWDHbnNVfmm5jZDHLDKTFByM4XHMk4E1ngv6TFHa1EwEigWG4SzIRXqpS
cpoHXmTREvud2X6yquDn2WhRIKSCu92LVPFq+U5QlqD3yRqGyqza1i14awWY
jQSyFLqdHLXw57tb2U9Vylv9ebya4BvD/6hS2BCB3NcSOyAshoqaQRRHpVdj
EV6CKTvtzB7B58gTZFn6uUAb7pw7uRSfwBn23+tMkf+/pSj7uNK8LLywlyXt
SbgIvAjQtGAJfoh5htygLUi77DpK6z96tveD4CiuooJtsyWJDvo9qjE/iltg
cT+xYQ2IrD2FiacQy/vmxgb5/SiNz6cvUKbbiLCCnan8H0KKYBzqRExLheq+
zb2rXt49Q4oujnzgNNG8TKZqj5cH3EwTo/Vx3LME+RVQ9RbjjO6f1SUDXvh5
R2Z1U6JUlW28bRRyFFEPSaMmrOnYRW6bUYPiAtsKUAMmvj/kLHEKX3KdGuvd
ARGt3xLlKrCs//ZCckpKjtohakOfzQlTZ/5lu4CFp3g1VybLQ/ZOo7CXlRvj
NlGPxj8HqHpWvOBb3xE41OYQE9zjye6o2K4r6V4+S1Ph8RaVk1cmS3MsG0JX
2BAHbR+blV1bAA93ETjKStEOgTTgslHMIkXq1uCZjqchHIMrd12AVFFCw9c7
DNFoRlhl3mbOhTAKYcxqIcDjRnwY+Xs+kqvt4mqkbGn5jk9qYUqUY3iFF1c9
eYrKvfEwENzG8DDJmjVnCEOjJylFOUxjM554hiPbWdygHnnIKfmx+P+rHmkB
jjC8R5hnlirJTm8jo8gzlk7o58Hoftr9+8vIhUeDFC7x67EB0f1KKpw8xqDJ
+eMBTRD1DykEUc6nlvBugnW6twHDhZ3xGmmapT2rJCuHRfPqwOSvyrO+u2D7
xXW632k+V7jiUwHXTgomvmtE74ms27R9k+J4IcPpCOsTQaOgxpEOsFRPtAb5
6fZD5+aU3iaKLqPzQj1jC+hKLIYb/J4P3LtAiTUXiO4pshzsGiuLnC9BfSDP
d1CE21A26/4E9qmXpgYRl0B+zTpiJDFiPrsMBy9TEtarD9dYLgeXb+DOf3eJ
LMHPX9b9wDdvBV9Jhoo0UHey5hcRShtnTl2eCRWwRNZkJXA2M+hlZewKwvnK
dnc/JKl1GHEs4QTrET75mwKGv1nEL0Q2n9vWL5zKDk+td3Kbl/i2G89NWSrT
PMxNDLMrCjWJAY8riL0kQzz6BOPlD6fd9h1JIubH3AfN4T9oMDY2NuTn3q8R
iXWTjhmQjYvDIz2N9kvuXpjs0SubNiBzWVV8//EfJunmbgf7GsKQJibElTmq
G/q1wuMHmxu5Hi6yLfueGErl1/Xr/iL04N7jiJDpAi0w81Twsjv7rIjXK4gs
JGlIbUKFrUaJvdZYEd4zBZ/e+aTVP+PdQppcEWeYlUVDPXF3+ZqJWyWSxy+e
iRySUk7nSogTZwpKMBuD/7RXvsVDPshKrMQO4ElNVL/brm5frybA/9kbulrF
y2R1aQnQb1ng8T/LBP5o3wmRoDDuFuksaEYot8hPynOYGgJB/2E4yNFGFlr4
tnDikFEv7s8T/aKnNXoyvb5+ksl7r/A3aarAz61eJ2CnKFHbURNdQh4LRrdh
D1gu3AcLs/nXXqmEdbc5Ef0cKAPyqawO4oT8hqjWQxyBRW690ptRR3mU38Gt
UP3xjibdhAuSa/YqTVzzDC9uwjrAVj5cHW4+Ji0Zxz9x3aRxAZ9Id6rW4bYt
x0RRJqZbaja0/H9cpeofspQWTfiCQ23KmEq0LWfG7NTD/SKwP/Uz7PHT0Pm/
jcZlHRrPrrlZeC0hlzTBCG2Nl4ax8Y1xzSbslGjynq7UXIyHZgZ/FnM7wr5S
bB+WhgrWz8TU4e2bkC5exkhbX1V5UGbu87u8XrJkN1XBF+KlFiN/RkdMNxwt
X75byVB6VPEbJr11wMHO3QRlRKY249Mwyr4agUEzY40Ah6RrUSvHON2CzhEN
01V4t9sFbt48iFQxJW+AfNy4Vp22FwgCbkTBrh41Y7t+r9nCsRj2CrXzIIJZ
72VpH2OuiwS7VxCDxOBgzF2dfrgn6Li3pgCtj4mNghEG9qFv/bbt3xxpQoox
N7UFCgj0WTdBCyl4AwPf7HvN7nnd7SA+xdFhfNzc9+ukCtqiOBTX0iRM2C4v
Di0vxn8ZJ1sWIqCprMvfTZtrSO/yXUGUp8Ak4fFlBmHEX7xZnaa789J4u+y9
v7DKLScOhNJGri7CG69pv5Djz60Olb5c1g7x8vVqr++N+ccmHviC8SirgsfN
0/IwgG/Fm4MjT2M7t08jcEU29hsQXX0o2cDIQSulX5unKYorZvK93UhJdQgi
CSfdNvNkVCn6C963539mvZdYbtaX8FiRHoAUkSlELJs9FWa3lVPmEckxrzRs
bZj5/ErMcFBNrYkYO5L/Qiw6CeBNp6kEChpILxEtz8onunbbSvazvoaLIpvM
UCBgzelS+tmolm8rcRMrscZxBWVQ+13BC2fQuh8HPh29O35W8FZ2dznvuMOk
i4TTK/PMJ+ZAW3mpJc6H/jrqquXpuMHE3F2mO4RAZ7NJ/PkbzoOMToEAgCAT
LxjNyfKBc2xzgRsTmOamJ6hvDV88JtRrG+nF7U4PJ8vKEIngtY2DRDpLc8/P
tEdoHqcganzgz4YDwlYS2tdSJFlbEvdJmp+Qd74TZzNTKZ7EcEufqx8h0urs
f8wEuP6w6GFG+IGmuCIMStf6hFivCJGL1W94LMbinCG7nKRYXodFvgN5pEJj
2zU+R8Sarz0s4uAMB49dViUxaMBQZ9rMAHclZzGS2WlxnQHy52DXQHY23MGv
KAtbU/FTDHcyMeqqh7lTzcqUCc1D2SXEJiWC3o3OtcmW7hElQ48pY4G1lwXb
5HHwMF0jpJUYUbfkGY77sZv6yUapy7Svks8ZfBxiPNqspVxhb3kEtD/5QX80
SzH9KtRdpxsiJFM4ciCH8UVvKuAdHfJGVj1oItWTqUrWTfvJfhxSdkh4Se0m
9SpjrZ9T5z4v4NqKk8iHlvq1o3cmhp1gpj9ui1CD/z1i7zBl/ZCeVDUUqxRA
NfXSPWmk+eVmLjwSPxAzVFXMUCeiFIeuTV64NjhrJLLEDUyO7bsN/OLaBKH4
D0WBCFwPSqwejjiWjUGJdyPsf1fmdy5bPoSa

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1K6KpxivisiIhzeYfH/b+2mLvtx5EXBRv/ucTCGRr962EDBNctg08CVy1rD8CNhOpnUTG9+vGSfEXlVgjvvWfWlxq5JXnWgycIPtr/dSJqPtAKMxyJWR2QcYHRqtsOqPaO5UD8OZRxlorCTSa03jgpFucqdv+mNjNj5Np3jBjYbgEw+ssCCQBykgG/ptmEWM+VbVeQuZMp2NEX6yjyHot+e4O0eUqJvx63W09zj96kIHW+yRKZjGpSa1i+pp1hQruiRoUny45c2s5/BxOO9SPmOFFMa575mdmZFtWw4tKYMQY+a1xNIbgArBhNuaDWfZlyuPnb4MfJwJUquccNCBdMYwDJZKWaG3I6/B8xcDcOcDYcYV4TR6Tbmzrs9/WZm3n5AItMTSZLoXRimrkymtek/OKRYT2dH3pGncx0QZqZLA38MZsonrNJihDGAR1ohLSR7rqzt5iGnwvykIJ945BSpkHx+IAeaemUSdd8jfk7gLIJSVntXnMp0p6EOCq1oZti/86vBTwF9jNmMcPd0HeZNHH1bBg1kRkArdNDppk1835uIgDouYUqpyHxdieeG/25Vr0G+hruQgIWru4yZAfz00jlaxpO7exhLFoARwgMfBYQ202jVXE4M4wlZNdpJzUMszuicic6jWF019s2bLBa2kCTxqqza01qDhyn0ukPOzkwH6JuMXj/lIb1wX0c/hwhTZyddWY6GAJ2EqKm6t5L1+TZMm1FxMvGC0B3OL+fPAoecRuiWFbvO7TYSDWgCQ1D0tV7kFn/zzpORnivgN2T9"
`endif