// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WsCC5/+ny3TqTFKyOFwiFGryxMeBEiAfsakH4TnAK0Ar5Xd+vcNLFnMxdGZB
yU8mo9tW+vrAs4M3vSOxYBwoNFiBAuuba9ZyP/vF8q9CQtEoFx+LYcISXLpF
s4ADp5TkMUacf4uxJULl39Z5So2QsbOeNyKIsTNxtxgLGJk0DptbrxEPcKyJ
gQwMgUFj0+fb41f5MWMJnGJAq/UgtdHRMD6N1pY6BnW3C7gpr8y6VROL5kQi
uNBCE8zgAh7tAT0yg+owrXpR5NoZGsMMc6Mx0WbiRYG8muMIvxwyV0ON5JQK
QPAnMSfMzJ5gudRnoLQEadX20oTrVbMe6iaf/xTI+w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
maJqTaePhGoH6yP7hEdZzQFnaYaDL4dYXtr8HLZ4bTZmrRazkQAvrBFRIkrZ
WBDc+BAzTpI+EUNNBJFYg1lWrD8di3RXOv2uZvzb3uXK+tXkh8NqEFIMTSDL
YW1cGT2UUul0oj/ZnTvBU8YdYm8bnHceloeJNwAiVrQ2nJwrDxUk8b1NZs5T
QPLZEc8ZwalavdM7WXm8ZhSJm8P6YOLtesqPkdaS1kmp2fpnZehOF8d7gQ1v
NxQLFa2vGNSSCbHadOzdNpsJ0AfZ1dZNhbJAG4oMssHndkMxdZOH8zMNq5lp
C+yu/4xR9xMCqamrFqPdFl+ExHDpEf8bvNHsJP5M6Q==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
sMH2Wqp/8AjOB7rFYOW1y7EhFjHRSeBjDzmQVRE7UgrCMy8F3u1/NpgEFhyw
2hi2fUj3EmqpJeBtdedfNbRo7s8eVA7lN+rOuNau4nR+QoSgRQd3V507gJWl
Ms0Sg4roSE+yvzUt/W7Ct+nvtZ/udb39jsciOEoLbNUztNSck9mHghKXNt1W
6Vbih4eq2aDASD0WUbyagLxHK3IN4zA8+jrlEqOewxkIT9BsOMsMmVyhrITZ
CUTUaTbpjVy9MeGvehiOYVUaS3AZ0WUTzvQH4LQrQ+mzBfUb9CtYG9Oq8ELS
2UrmhQJVR+GIwN6iPGp0tMNiA8I6ykZhZs3/QqbW3w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZHHxpRE4CwK4B2w2lsBc8A9Tsmu8xMg+zb9nVNQDrv7keNau9JE4/8QDKlla
MIdcshLWvOID2OhdBzHOG2kkaR9Zcw5rCflGR1c6/WvKl8o+DRCgNsdOIalN
IwTFKObZPABLYvDsqpjmUmGwa/253R2icaC4076F6Hrv8t9jAkHVz5FjSnQM
hCBrJkbkOB4lFXo8KAKHiiIAT7BwY4HDTRVRwlLV4dCIvsl0kuBhAok7RJpN
WYDkfAvuKYXqaTZ4X/RgHQxbCaDEIXwOrvgGjervmDw5GM7o0cWNoIwvny0l
wyWyzXVzFEfEb6GaUdke7cwSzCeNNPvg2DoAD4u1dg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Iw+M5y50YeQZiB1yHbcDk4+xgs+Yga8WBpadSUgXkyzxl+7zxjnVwkZQL5vS
k1WLfDeM3XlQ1+sYTQHUY7b2icPpgJB1BbFC+2gRpbD+giTznRGmkUZpbT8Y
AxMnZsd8YouUMwy6X3ze4xR1362/ghOXnICuNV41SUkClOI3nL4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
WfE8diywTIu8DMTgSUkfGKAl314gqNOeoocahBZ6C2Oc7kTMwO5vGy1LPHO2
FX0KO0dY8k7lA4jdp/McZ6AXvTc1fQ9Bge9/g/u3aNCiCGAoR/sHLMQ5s2zg
JIakJ74sBerhDmesK7QA2WDj3/0YVbJyZNunm+Kk/yKLk/0l9tCb+9/9/iSH
HSofpeLfiFOXU8jhgq+u5U+5xbU+3DsWZOWEPZGOEDSkrhFZz7qdsJ6kj9eZ
538omyCyHYirsUudgB0Lqa/372Xnaahzt3idWRsX+8xcf4SmFWXMBau/u6ZC
Giny2gSdnkjJdqph2vxL8Jafgz8HsINkpFBsqo/0QEnXKdlZTtsRBosj7gEH
3UJf3dAcSqZeYE1gYgouqXyJGGkvNIcSUmfkSXK6RvoOHkvJqLfq1dVKzb9L
JWWC8s9h6cjYhVMkATY8Yf2Jzgs5fT0079Ni6T/R6Vob1FAk5g0DO710RllI
/AZ+o7VpQvveKxmH7pXZ2dDZ4aMOeZZf


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RFQK+pfWOiRnd5uLGIsk3dbEc4balpZRCh/URcgCcNdEgIeasWKM1Dk0TYCs
J7X1xoEh+MiuThL+2YO9+3ugQ7hr4Fltat96DcpW5xG9k6LxkqGWhHH/aq6o
0Orhdbos93EqukuFIutJ0xJWUKUWFoMYB72C1GyrUjZmXFt8zSc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
C6jHASDnjIo6+iNUPVB+5BT2nUZS5gmhduO3dzHBEha0ItP35ak9eTI+vF3f
ezaRhxLmQezaAk4obnU8ygvhbTbaHcFjwlbM/ENQ+/nx4CUc+/EOfEEvMDVz
bzv1khRLiaJRnvZnffhQOsQrhE36vaB6I6adruVLCp1kMw8nRwQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1040)
`pragma protect data_block
ftojyrQDXlWN9qISff2DliKMULb+8e7DdGVT9+KjH271gXdKZTDMg9fD7Yz8
ZmFIXbtItQU0mST9IbpSSrTXjco3Qq72+njteAdw48axO642AteUlo5sonkt
dFHxFnKDJls3NxvdUyARYHDqiUy+ycVT50C2dbwlOP1IEXZBjTvxu0ori4Pt
4tZsSIBQFD6ZuUSL6vfFdnRFk2oncE9SwgGyS4zpLdfdLvLiMQdHsUfGng3l
fU3hAjbRRhsiDCbPUrkCiN+4zA+xHn/px/TlkEJzK7NQDJZV87x9rMGn4qAT
BlzCr04mLTD3tIU+OiTvXszAiOGeP6mqhRLO06kr8MTbLbJsExnU9+6ida2i
hlZym831RmRKKYM75YznL4W0Nibmbyi6Xyv8Vg4bv5rT/9V/5XAM1h4eJmqw
Kw4k3cgRbMfmhzdRSa1gg10VL4n9E0DpjZuxP9Egs1SNj7ZAK9tWBwxVyT6s
n2fR205UYC9ShSh8DczCI/XLJQ/1s4kyrDknhTEM6RRDJBL9Rf3EAVtJWGkv
yVdzB7/8STFisck9eRLUEY8EkkqJxF4Yi27QlS121IetBgq8o9YDtDjMkMEh
pq2+YjTVfxkiC153k0xgzDvKW4eKNZ0O2q27Z5VwnDim+A/CJw61B1hmN2ED
6A+7v3X+KxT6US0sNOIUKth0SddyzntI0g91rWzZr41sW/ERX8d2/D1zXH74
gU3irl41yi38TbaMRDbBrexZTyGF1xO9wsITR/HSleZJrFBuEnECyJmLv0qc
c+xY0XtIB2v7wmSy6avZqlTYB6L3Vhck03kQ6UGl4HAT3PjZB3TXMxIAwTpS
moClrrmBcTHHCQOlj4aiu4sRTBBOg9Xl6ugzz5OIz87gjgo9O/gCGFs8SRo6
6HHL1/EOegDSCxNnD8UNgvTpelb/AG9mohtBUdOv7xx7icpyR9VMFrS2HY4l
RUdinuv2ph8v26d47/GHzOVLpOb/uUFCA8W2kDTQoJiiAD8q8G3tOXzrjLX2
tt5hSEYUVzuZb9ZlpZ8jb8XjUMU1dDvjZ9yF0WAnuYW2NjGWjaLEsu2o1bFJ
wN5yyeqtZHm/p8OvWmS7L9RbIvd2LjgIpE9/iSSPHQy7ye9bjlkTl9X88kzt
pYf6obaWsoTHQBh02nPUS+AqVyXgbC59JHscVzilGkz0bgNgQ71Z2yQAJCmf
Aophl6M5OOOekLcPbIDR4LCAbZPaSk6pPbqsM5349jFWDlWHpCTrOJ7/Rw8S
Mp2fW1DBgt8uhLWgK4codzKcnHLuOiCsmmPFyV803fsXLhzku4ap0+sB602z
bLpGck1rALA/hUnFDCAlKMsNQs+ylABAvJ+i7F9GfxjJR8EOLuXsPRkl6RQX
9dHYVIg=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqcIdZOI/p1rrZigl8oGWBJchn2ElOFdykHOCTEHy9ZeNXXEKm7r+z1RTVg1Xo8O68VuoqeaSkEqnv7Z+7q4/xPcz3WsrrJbZlPr+7dTK6lYYrFs/fXToM+IOH9RDK4uCJls1/sZfKw8krbBXoFIpP2jlclXQ/lKe+Dfp5LLIBc/XBuE05jwQ4fVK7JV9OgDy73NNxiKpLa7/KDXMi/F7ZJDY07h4RHQ1elyBKSuejiOvuXCGr8SnUJusJWDBTZxbTobPvCGmuQgvU4xRdF/3DDrGzV6DgoxxsCaUsIBjuhj1A1tcbVLXGKKV7x7Dntakfd7Gg6aSAjetfMuyAsyPoQweawcix/nDjDFX/zoiHo6TE0UrWLptxdEWn2/EecH+zNmbdg5D9Y82+JU8MPZtD4bD+lJnlnXMJr8Jgroa864omH34rMJdsBd/HqOmjAm+O2ybVsSk6cGIbsdMcEgWTl3LQ1qSFRpmD26K5Zra5KgLquPIaZuKsiqoIUvXcKJ8rrACKYHjyzveb70OgXDyxHekmUjIj2CZ/k6tbzVlzicUC4iCQmYRhFRmYUNPozpOnKYOiKjsqswifKZY/TMQrFv63fbI5m1qX52QRlJl0y9kZY0magYSMTFuw/Csqg4jE8Im8jbBa2kUhdg9wKRc7GFzW6/5/KAlfiEpHu14hxX0rsmakq/qqOLvfbhvlLWaPnMtMc+TjaZu30ZsxG50qQtR3BG2cLvPYossm8d/fVXKbzXEqPhXB27N8M763BZr+OmwXatiAXUSFNyN/n8qHMp"
`endif