// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MsLs/d2pPThO/tiDPz+D1wmmujwQjXgBIiMeC5NvqPxmsMS32DjWNqvZ2as4
8xR2nmMfSpw3fEw/S7DdfM0GLwQFbNAjs27kPfEd6xfKHfgbteS1JEK3aMDz
LrTjmxEKGRz4LzuKcPN/n4l7sAZ/kUuheX9jDaAK3NC/FlmX3SnK9KrGqaW7
waIZl6Djz9HBfOS46/xX+rGFJMylBBiHsypLBpZ2GR3aHCZn8HHxJyBq9eZQ
rvzvGRWDAK6Db2VNEcfOZm16XNWAJgzVn6LdOjghf/zLGAG+gZ7efbhRaXrx
gVkYdW2hokDfxAy/1u99msfXsvETJfdH42RHKLPqRw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JNTKckUBIn8WR3oistDZ4VQW4I1uyiCdfuqBXP0U5zqSsMwjZy+uHxWWQW8C
5GfDn1gB+s+IPJZEdj5II1Ke7e8rPwef0YRIhNMqkGJPdtLkAX1hNlt3PNuT
hAAE0gG0NFtsi9tKOp5eBWrQUMqXnODiCap3uys42xK+xQfJZ3BzZnaWTUn2
Oe8Ia/KSn3XILo6ssPkOPjq6rhcg3hhI6AjcipFfMCr17jZuI1D/tG3SbGgT
m87Doo4uRgEn24mci+jhfUbz44CGrqXiBjOOW4dzty+VNeUhSOn7zGIxYqlL
WTst3WPttHRt1ZOTyIIhPZMmEfvnH8gbbops0J9DIg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qWXcXvq4VKln5VSy9opDE4gHTQerW6Xeos078e7tlOiiWs6DLUEnz/eZNwsh
Cdk9JtXORJ6BeAybHVupdwKcBCacctm+IdbXaM6S1/1hVxPqA9ImD0ncWqwe
5wVuxJkwUku5QOJ3b4XJ6CtUFz+ht4jLRKXy+UkF40mcHlnykc18w08j0ted
RmmgzGDr14ox9b8pknh6nrKRzSkbG6gCdQuOv/Ir1Xdxixn2s6IZa446gw0k
F83scw2SlDwLjnRsqHgTzL5B+puD9rsF3di4u2/b9q8C1EtI7HvgezBCZ0Ss
hPPmAsjfjAU6/PkrN916YA4BlmKQRlv5hHEacbiWKQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UrD22kzyjfg15x0n+rNVb8RzOHbCStCtXzxfu57Or1lU5WxJOIpwyBFgHZ6H
n4S7AglxXcRPYbj/5ervst6ow0/3dQUInkvZlbGjBdOOALnzZC1LDGbio+b7
TLXFdrdBgZyFo6gRwWqn2chA3tIvQRT+vT1qF/xayE0yJXk6D8D2FLNtl0ur
77/XuMZbrmLWbnIdLEP2auRHpBkC63L47gHLQfDEv02DbuxsV8pmgA9nLAJX
vH/XcvT2vW0kjMCP5SEb4hl4HCIpNIRcYhOCe6dvz74+wkud7F6MRfSDXmLc
9p/IreT5/kHon2iNvqJNVQLcMgjGpzVUevityxBw9Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HuZSKWiLE75sK77Yi8aoHiy+Dy1yCvXaDL/B4K/fleBOVDTynPZ5hQaPEf95
9t47wxje86vzobCB0+IrZBayKIUfwPkn75ZmJU1/KCgYp93VFE3fyn4C0TOZ
W6qIO84JU8uyO0a6uQN6r0qi3mW3/3KOGL7fniB8YFzP4y2h40E=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
iUPIj+fGozVCh5+12Ot5rznleodC0yDoRpyHmwpRDZ5N4uOf0PIbVDY0ljmw
r1oRHlepefba62oVmOVat3jM4WoAdsyC7KGlh9Vi4wxfofb9bblZBqHPFk/D
Io/ZrIdiSVc+7YQogNrVdNXXiz+odTMbgaA3CG8tVrnxHxnCp0l0S5X02+lt
Ejz738r+oj5STI8teb2MfY9/QiUCBDNYMisBylTlPSwPuUFDABIAyIAVJG6f
UoUokNPgpsz2mnZZZkqnXBXU5NKhApIhmFn5TPDmrO/O3U0Ko3w/8Etb8kCc
OE/4Yn9cEs9xToXt6ZV3cBQpZID+YucYIPmV1014Nctzi0FfN5c8hLpN+K9Z
tunWNzJvPm8N6xe/kbGXMmRWfUs0XcAv0hp0ZZHVEPY0sup4XBBVU1X71yqS
DMXZuSGCRz7PUx6Ylfy79lNauqdroM0sVXYqm46xLB0bWnTMGQeo9LLAgDFH
MZMzj1A3D1Z7WdrdcyOakppLc7GDcWKb


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
I8DvCwX4ZCQYTXA2/osQXgtV0uPg75DzZjZ9G4okfo/TIX0b4afj2rocqh6G
NddIXO49odNPibk67dz10k4Wx7IcTq5dwgO//6bpuTYVP0RNyaxmxPLctbHt
TIdvWhjYuZ9U319+0ZfJle7FbdUeqZ9IejglOiIm4RWvhjqdiws=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
flB5q2m6JgNJgbuZZvBZlYZmTwRUY8f40HlNc3itM4S0dS6gaS/EPZC6Nzh4
GelJSSaSAWy/XP8B4TaogWPWa94JMfmNPGYBLcQwUI1JC4vIWRvg7Qj8RRyJ
f0vQ2WEoo7x7nB3PlcbAzva7Mjl9aMvokcRxnIUpmwqD7y4A794=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 36784)
`pragma protect data_block
b+4kcFlj6yV8OwOYRURYdY3X3NqfkipRaK8msvWqkYCX1RVEKP5YNUiUfp/O
Rrto3s/w/Ps/cnduuLDZYG4hFkuRSCO743omFTQMw4VLXY5R8fF/sB0jqDd5
l52VXRR6/t1WHZaAZUEflGCZ3hibzYVr2UZceSkXFTUimTVixTTo9mMs6xW/
98iY5W0Hn2h9upIboYaEllKWwPR/J66AwOBW9LWBnagM4byzCvnJQRkOqzDA
JZm7x41VJ3RPu3TNaCajqXFwUuHohIGL02ruQCJUtluOTnIJS4TlGBFNDUYE
ukE3wPItZDWeRj+/KI4lDbCJwJ+aICwa/hnMiYvnn/sNC+JBIHIYt/jVhP1j
W/DlI5wtwg5vWVqtqeRQ/EdhjHeETnAsc1XJKMLNQjhl+oEYgpt3nicIGPVJ
GmCVqcn8dKGmib7z9bvX8Zcnx3Xb+tm8Whp+2ZaOKDCgs4HEkCB2FKDxhZUo
4K48lFhhXufJg6Or39WNjMFI+a0UkjitHtOTApKuaqfKmg2MQDb4ppj4cPUi
qEFfgoidNUyLlkHDSEutNVfj72ddoKy+xviPlNy6HreGIkzLumFNTjhHYtMx
Cgu+j3+xNz6O2UN6Ut8i5OxOnL/5z3OLv8zz7vJBA++k/aDcq581N9GndZsG
o0708HRdjIJjdchjTijwQkdByG547E8UJL8pTCRGKpL2d4a7wNJTOFcXapVk
potOUlNEdxdfIptDgxfnm3WaAm1YyjYihpP5rRHCTljo+m+ibf2vWNDWGs5U
03VrHlgUSQO5Dbu7FGsAWQr1FOPUo+URLJkRcGxBJ9Xw39yda36/RTErFdxP
2InFHTAo9dJ2ohO+C1HsrsUnTjQhomSOoM1Fc6jZLb8KrAletzer1qNL3vDD
PozL3uxMDWd95uon4vtkzqefYFW8Z4VCIveZUJANZaZgFbUa9sZmB2ABr1R6
wi/AZPNfctxD3u+FQCvV8AyojJ0kxnzpPkwNQt9byTcnhZfdqzbhDtpFKsY1
cPZVH4oLkQaV2JAF0N1nz8AwEFizZdg7gYgS8ot/cjMXbqeujibr9f3XflaZ
z018O6FiOAkl4G5LDGVCIUAQ2A9g9yIHbLAEZse6F5ihCW10FS5ef/ymemwm
77MrnWxFIcxH7c/wWcyQ0MSpbRZmFZgdro1bJK/YK9/a0U8wkMJQj41hAmDa
X4XDea+O8sbO27azzaYF/6SjtoJHxRvRm8JKXGns78iwfKLTRoUDXf+ucu2o
biy5G549GoDnxekYvGo805gLkILRUvCzM0Zy1BjCrEQo1NUNJWKEXKNR2LR8
IU91iTsNT+d/qVYXDpXHG5qix+nVRgs4RNm0SOVos5rPUa2/2ZlOr5umBJpS
/2zQcctbZLdspgRAODU3oNUgwyu2zXqbffTcbKPM6nZNhtFMz9/RVqcLISup
DSIVAzpptPMjsOelrzyA1V3O4hR9RWmvvDohUm25+X/aKYlT0woVpd8rSbQ+
d7Qdd/xjy7aqr0QpPneQjzkeOVZOKJqXV5V4hzy4hdGc+GZYccjCxL1IRmbr
NtnZVkS/mWQJutOKyWxGMhturqIuXqCM7/Kl3M4TqGeiysy6DHMd4W5mBv8g
pwLle3zuJ2rQu2kAtBfdl3AIt3/MV6f1xJEjkHKDxt3trX5v95uC84un6hPV
ncRpz/jldEcq+JVwieKNHFja7/jIc/FNyfP/NZNQ1x40G7t0mGkK8Eb6DpzG
gtJQGnaHJEQxh4Mmrjzo6toE+D/u4njZu8coqBqfVQ1r6M18njUanVEbM18j
8pYxN2qBR5I40PuO4iXY8rCq1vUZZ9hzbGVLwxDH1FOW8IBei/OUFU7jjX9r
44AkYMDTpL7U0B4a64BG1ngTiObcgwWe7HPMG9kJiQfYlWKBFT+aximwQRUG
/upvlWEmav1YDCh2tj4dzKK3BKxA5NvksUxX2DVDnBCffwH02NMVShmKkzDR
M4MzNACxjEKEILX+eoEj5R5AJBH4NrPNtWpGIbGFDnAVLAW64HI/BND44a+a
plqRZ6KQBNv6ZkAgiQPN3219qMvWD7kEodYJs7ncaQcbQY2eH52qh3VizqcE
y0KAS6WibDw6iWUIElXDDEcIsCSk15QPqmvNDJGw1qv9xfqOEzOQfJb7Ddns
cnj/s6XfJKA6cE1FgY8WPXajmqSJUVDIywZeCx/LJJ4SnnyJI53W+r1Y8GAp
TLN5V4B2Y/8YI0ovY+RzG9BVOhyWTW0qgyur+H9eiwkFuIK09r2bsMxK6LRP
ATvVU6uOSRq6ydNa8ZS1DGUf8dDYhBx8UMVf0CJ3uWDVsk9xgw5+iRCLs6Do
cL4QV8VvoiEQBCMEDdyqRAsa4GN2bQ2mpFjESItzTlYDMUrm8l0Xgb8aeBRt
kuUo7rBYeHmyFQSGsYMaX5QYZh3draAUMvltOlAf/UOA3BmfzZgqAclde8uM
EHpPRDNsvy/pWHTeMQoCpSOdm9RWenD8S4DeqtdFHIolgF1ZC/vmHFl1OD0T
w/ZDffSR73rU6c6QHvwR3g/iVQmhKxbmw05FYdTfGjNBH8hN8DW2uExNsukF
kWEMY8qHIeviczw1q+0ddBmIVr6LT2eDq6PFRnjSweCRLSnJJGPe10oTzHlF
otymete5i23kBOrKwWUvBt2FeFO33glBgseTUinTQanzIEfHuGoTfpGkXQZa
cbyksJ5K7fzcd9bg/Ot815ClugfFKiUlPKgBUfqvL2lY90InrYpuREkV5+kM
MFJXM5sdvz8Q4jooNj9IKdRQ9LPtncM2vM+dUpJzszRhM2S8rKiC72ASPvGt
xOiebILz39aCEeooPpLsGGNPScTsszjxzE+7B8tcH74pLnm+eYsiDJmmN8DP
9NfXj938MSiiike2NEH/lz/uH2UBgdqvhkVQruNn8OfIzzNGadSjaselrT8D
krn/tlIdLZrI83ErgC27c1DejBoGPBy3kQdVGd6juIwHSH10ph3tfTnBn8kP
DEeBPbpeyVU4NOmnoxGYCpVdasCAv/xrOa5wJ8hBMAL6m7aiBszqOJMFwv0W
6fAyteZRj0uPIKbqhyXCtoayhfjlz2uOv/wKUGLq/pjyD2sr6uibZw2kFuYo
P4RKtwhlbIgT3S2L7gkT/AeP3aaLp0aL9TCnp9m2+psBIyl9Jm7xNDj6F8zv
pe+IahysYofxwBQ/HcbYbemw0ORFGdvmsXLV1zFfwzDCI+wjHdl0ZYMMlHzD
6oKbMfIxnM4U67ogcOjraPjGqOeL9YYQHBm6QoSGULZkJnKnBBuoF6L24h8y
AGSF2cKWpSn0VhV6SW18/a2i7llbltC7ZVB4G7HASdoS1/qMhsNT7R/m58Qg
o04NFYh19JA42Emphbm3D19OXSBpblg6jW4w5IbDO9iKbol4ayQutlYhADJd
yU+lGuzrwtR/3LF3ZziwrEeC+klle2+CvSYXpQzPZXyae0pAlDq+0mUBbuiD
7qkI0yH4HiXSQWZLbDftGiE0+E7RfFptJ5wFtvsDLOY4KbM2rBO9z1eyVLKR
V6J409tfR+JtQp140PzmcLyi5NXItEGm55dRcDzdgoQLeOg/a7rL5pzrb7Mz
aKJuL5mZdslA1USj2tnmATJ1FqL0MfduPCDGhB4tVnZkEC4nbGrLyvqBb8Gn
VNuEZ4IFZglGqe1EXCnG/NnoSCyYLw5jhGh92gSaRgOpkKIkBDQXWCyp2zin
CC/LxyTv2H2gNYdn4FqICIb94BfqwFNBIRnVjVe7INfy+oMzakhs2YyJQQ65
VmAfNDWKYp2N4Pg/kGoIrXWosu7D8hE2yhnDrsFJnnbfAqpVC++Iia5woRto
P5I7PzQ0QJXxS5b/OnpsWX7zXN96V9na9nmJ+uQZ6xfu9V4+V+TWZg9peaNU
qjoJ2lmnnbLLC8ccFQWSqEzZ6rV315V7BUkL6Br/alGrYpp+30mudWExk0Pt
b70xFPjlLBCDxWYF3fdWp+PlgrVmT9rsTprkS9tU2p8uuHaM7lGrCPa+foa9
faQQpc11K/1jl2XAXN/V8KCO5c0qSVTwIwbh+mBTkMxQJDEzwTtI5hJIvwrR
2Tqm80CU9gYKJw0IzXKPY6aV9y0jKoeSGiTSYi4C+G+u9XuoN6szzf7z+tQm
YzLMOOfzRD8ECjbxnwj7iWu8hcmGYp1wqweq13ButztwqRsu0zi5RZ4v5mrv
AynGOc/Fz/qv6JorkRyybVa5uv78z/pz5qLixalQFJ5zWc8iKpj2wH8pQCdY
hRxkEHC+FSCixuIk1suTnkN/jyxmjSsAeEspzhrm26neW81lFaixDpcXFwF1
NmTs3YnBjqobuzylqCWcU9IOgWOSKhPgdDWvBpWVp0zGJD02/X0pWC1NrCZL
clNbWSFqnF+B6Dl5szbnQSoHRAwooGCFzFK42tWJw3MMpj42nQgQ5iTqcdQr
JHjQ8Zp7wzm5m+L9lxgLql41H348JCfHf+Y3qajvU/aGv+M0gsfwXfLdvNCQ
B7/4KxGvmRuR/Fp2z7DjJGkf1WvnwPghCDjCSiLqL03H8sfpvhdEOts5Dsu8
uMtztcK9PrQ05/1n4eNUJBO6zLrWqNToG/QxPbvJ4KM/xCwmSnNV06Zqxs0H
ecrOVCcoD2Fg5FDoPP7WvN8XfgzknGwFPnJGUBx4laXuvQ2jWUFtubouCCbf
11TH9dhywhtID7iSRG2YVwwxciYUbBPPg96bThehgEbSpg2yLmVB2vPjmdXZ
k5QFY8qX7l/VSRHu6YeSxB+120txzGCC0jGQxJ/vRogJI6KDEa5Z1V6Jwxnm
xsUCWZexp1SYVk3yK9jG4MLtPuQFTLOK2q+xBb3rGgZZZmR1eVodoHfh+iho
scGxYS3MngeGDa5iGwnGm+jlPDF/U3IXfnu5S853rT3gg+wX5+g4s1vgMzbc
WApb0vyoObz35MjLkw8nhZ4jzaCUlH9sarhXs1gGpMkBlB0UUAI3YhFTNv5s
F51RZOolEt1xgOJSpOnR5opmMAQYc3k+lPb46rH8g1uhQ0X0ohIOwhn2Uw1h
W9TT5WnWYAEeZYEJyRCR44McZ3QdHzpXFC1nqMAJ7OO6P1tKncsQD6s2dRRP
yhflmYkkt6OJDQnb0x0Vn1KQLMw/lR+HdZMO9OQieMHTqkI99OiEj737KlCM
+8FxfzHj4LhY8TqmjpIfOa0inHjh30/3e/LmwZbd4nGOG9y28Z0EqUwtcHLr
zvBSrnaZwEKqtA0ctE+ay1a4Wrs8gT88y2ye34Q26mLxYhFk2IbBi75sljHe
kVmOSwmOi5xsZXyBPpIy48rBRqsNRmXlHlP48PnrLkXA4l+PbLZ8NwPxpz4S
qbPpz3/L+ODgaJwCq4UwfeigxupsYU90gbGHZkC3ObwOPB097wUsLn/gBS6c
0rjmkLwBKPCn+AJ2fJMuLm/+wFh2GwXi/2tvOLym8S38MQpuUJAprEBjZeTR
8atTkwZX3JKjNm3zoAq7rdQQ1CF2Qk7Go4rDEykD4xyqo+4K29ao3W/uB3VL
HvCDdWqh4gDuEKykzWdMWEc7+8UbiPgXE6Mdr/ahQsAXMWLMkJulWU5Vu744
pwQtlm22icySG/KsmMRHPOOQdTZy4WvdDda2DljTjp3khMwy4v2DhYib17WY
AVuIL2tndYxvcSVL9kDoTSNiMk9hQ6Ok9FHeIgTIEpTwH22bV/86ux7CiQGx
GNvU7sLY5qzzuG13P1hmBD9hK3CcFHgvtnpBZtbNriwwL1nkO8mwyc+g6Dwn
jUejjMCEWi+FCWB/GvEDmSuE0SgU2lVqnWSINAHbQjnF5TI0TfhtsQu2AHGC
qz0lopLAS8ezOwXlUQr/BXGce7kMF1CEYJ6BUOnDeUzDjTqUraW/cdV9ET3/
a1I7eOoogY7r93VebsY9cR89pnQ19EdZibj7Gc/vf+rYS7h+Uzbmfn8xsWlE
CX/WBku5r5QkWKHZHuSjhnZpdBPARzKF6Hhc/0wlrjke1uQQWCPTt2XeGJyO
Zn0DQlZhUf8bGXcP9hagj/UTFnI0++TCx1FCJY8ZIpRcAx7FmVOmVCKYduZH
C3N78hXmAbUKQL+uQ7ZO6srLXixJtLfwn7makFtsnyI8eE9c164rCt1BGBba
NJYhvPrCBA5NcF2VHJ95H51vjXXZaTAlxKADWkmD9a7lB6jqHGhMvh6iLfdM
B8c/+q1IxC2LwTN7aq6Ymae7Hc8LAbylI+6S2XSt/D8WTFKHJSzaQf0HU17s
jyah3a353Ydc6gPiFPzJcAoGxSkImcG67LvcSYEHeJ776jo1o8FZ+7Grth0I
iWsmNh71FHYMImv7apx5Li8PCw4g9P1ueOwzc8tGID70+35S+KlD6l6L5y8X
OSqTe0jVrRqYc/MH52XhjHDss4I3+F8WXiqW0Rhv6WAGFip55IdBUjChSZXU
lApi+ytKd8WdPQ2Dm8x+/+2aZ7V+SRuo+VdSskRlAkZya/fP0B2Q3ymz6lzH
3uDdMDpY+xmvEunX3BM7OiKGrXKpraJDlEe77dO5pzEELdK4Z7ze3Op29jDi
dozAgKwjfU/L27+BeZYneI6Lz1mibHW+lcbFgcbBROaoAs3d1826tCgzjAlQ
+xMxan1u0bdhpgkUADk3UnFh0M/CHcGXF5zkqp87YxYzhOK97Q1tF4s2NPdX
IbZ12X7BU81BMtAkwspOwCMdazZK/XXsWATMcN5WBQ4HEFIY28DTSOK+smoy
5L+NYA9SUdGq8qNAPfmKqn6bFzqTMGlr01weXzQttityNVnpOzHzrefCpAew
dnYeN6L8JrLrwY91ZH7I7ekbEMPQOxp2vfkGBj3VcUrOJ9eCzFmyH2GZofwg
akGnj1sfvcfetPITUp7x6ISFceGgi5iWPkvuQ2s4GXoc9q4BIBtVxghl7kfI
DRBS49r5lyCoD7Gkq5JYBNMtvlx6xrTrlQWja0u1e17KDuwpUjurVPB2pz8i
EDfZZfClxLhy8+FsM0cJooMbujDPstrh4U3tTwGweQh/YzWfkujvS/IJtj4f
QBwRJASxyheqTtl0hNYT+fqRkB5A9XaemvbZVofUMvT9CVrvL8lovbq1HsmD
8LGn7qJmdNubsBdFiU0j36Sfk0qpRGPpxuLBQw9v7eKuGeXxiu7e27jRFbNr
SISdvWlW3YqZsv9YphazLo+oiZPDf0ZIJucB8DuBLQM8fCbImo2fwE8x3rB6
ORfue5zNtOEGzvBw7ZluBmqHtr88Ed8rVRfP0BjKWLEVHky8qkkRmo5j8XwU
hlZp7r6DjwMcwi+1ElxUgm5LvMEnzVWhYzyo/d4u8+9Y1zwuxxsuwX2ukX1O
TaBbfZILsjuw9gdPVzyZVmyxZlULwAD6g47zOyJahzDt01ThX5oojGwdrePT
PiluKLh0xPGN699JQ8OOGTgGieILezHUHyucyMaJPDe7pJfI9oOh6uRnlkIw
Qa9SCKcMzmR9uXX09vttozq7Id2Toz0m4ZgqCaDC2ClYoC4bYh9qy1iuk3ZH
NlFnn+XX/BdAam/mxGcmFFiIkxExYyMnjmmWLloAKcyLGfQSuGajnYyuYktP
Cv3w8pRnIq3XbV1BWYky7VZFdObkZhJUS7l7QMPeyosKj5y4jkDV5B3cChjP
/B9YQv6wKk+PL3q3z5ajcmPozMzNWXedqbcwS+QIzB/Rc6cALpsUFy/8dcO/
4fGGNs6r6F68uc1lRUlTGO4Z39zBN67z55wZPjXieXfVTgQrsaofa7kRjFfq
C9pqk+0NNYikm4jgFF0hblTEOpxzBbc0C7Br6YFEqjid/rsqkoYXGTthinJQ
0eOFBz2qgua5x1DFZHNyBAuvCpZEJI0RpwD1ondRToz8tl6ZTbUW0xU/s3zT
WLr+LbdCg+bCp+7Wa3SpLdMEhh+zZ3jc9QfQ5Wyds7QnSrnawkwVfQhHjuBL
vjP6wzY+a2AIldrfDuNZPrLs3uIjUSvoHsupBtdLLTamUasGE4CqGNQr3v94
PjGGJBANyUnIh4bHr2o3Bm4od3PjQypZwqQCbnzKts8xjbe82KaBhL6M5jyO
eCxepeHzlAS2Ag9wWvNfoH6zQtmSslJ4VBuYXnaTLBbxjwb7TeL5jF/wfHd0
hvMa8WIWLK0Q3W1u7+AUYFcJpxSQr0r8T1Un0CPAm114be4Hqs9hy51mWgzc
gPxNz6z6XF3TNVtKzn6BLOZIEEWCfHSL1xCsRLoSjqdYKbPsl7Gz4O8tZiip
6uIvDMt/JQuuuyjWxcc7nT79RS1iahYc3Ah5ZZXo9Jf5sEYDgvRc+HSmHCSH
NBDgoD1qI/JFn+SFK7lsYDWcKU+l6Fv9l0PsR6ZhIlYsBdpICwnvrDRFiN+J
vbQqRlDTjUgynNq2U/na9gwaUYGfdt7EfgF+s/tZXqnVSWlUtGhw0+fXv9cz
zO2+yIdJCvlMBjMY/Gnp0nqSoyio9F8+ZVnKn1zeGxo+o63gKfEuB73kUqXR
HOwyc+dir4rpm+vYEiN53H6w347JKb7Y8ghPiT6BwUZmFp+kdeVBd/51Sume
6kiwi+tKT0s+xvtVnGGpoSPm5zpQcLEppRse9SsOJThv4l52S+ClPbsdBgFi
8b0kENqW/kBomrSW3bip1CcZjswj+9Fbprt9iLd6Bmpp6OXXyRaY8XyE9QLl
h846ebMr5GLn/t3PbEU8olPoZ/tF3Ahj38LEXkvERzPlQaA/kIvdmpYXxa3B
zb3fvZhPLHVIW/xIRcnYNCoxq6MtiSVk/ipFtFcMXF25ZtXgYUGfrpF79T3D
BkF7RLOoQ9i+v2YxH9NUc6510P8WNcwMBMtnfvqtfV6qS78YsciJCp+sWjU9
2G+jir1T6GwTWixMxgcfUsIOeGdHKAIn5XdefhBSEgCVsDrqObzpxGm3+9Zp
LSYGBse2LEpP3I4gBybPxDtrA/ydwR01a2kN0LaiR/0HbbuOKtpr33AIpXQQ
M6cYnw3hDq4HUHf3qysoMIRWuk7xxbZemOWXgydTfryonQkq1JKEFpxnrkmX
fkR+Val756Ea2DwKAjwjtOmROSudGe0srMXNQip3pohZdwYAuHhEKEuWlcpY
tTxMfbQ2aQn8SnzMgwGTXubz+QHpKWp5xqrO1JreN+smwCcjgVvtPcczXYNz
Qa4dZC4DLpQ61o0SZPZehOutrcTsbUjwu/8990nJSXWApGmJAHxvc8qozgOu
GuyxladHrcjbJR3c9CRZqUpMX1+WhSlQjJDLPEnqcDl+0wtmMM8mAKlUOjlH
9hJo6N1tNZAYRJZlywS6k1a0B8tI4iKro2kGvKVo6K1LtLZ0ekNMdXfn9ruZ
RueDh7M6ZK383V47EIcY8t7N87dcoz8kTg9CyvwNEOaNKd5+bJEcncL60BL7
yaEVwvrrMZmsIwgs3ww44lZ5dkzaiTrV9nT1TK3idWRSe+WC4A93XVkvNCY8
v3hmhyUx5mQ5+FkYuyCVZB4BccuLxbuS8NWs1Zq4VVvNPFSL5vTrtpUxDSdF
i8tJOupWrrGrYvW/Joj52z4c2y25nG2b/5i6wGjHIPkZaG2Ut3Axa1VR/N1I
GPaoEmmXE/MlhX+4OroxWVCJ612DBUsizRBkgpgiQ8Bh4kb+5SFb5CEL1Qka
Vn2cA61A5+O024ZQ8JHG/7ytDIlOfSsC9D6PcSoSYIqZCeuX3/0ZWyCJ2eDh
QhN0Z5/7pqqiHTpk0hkHTfxknaMMyVz6O4bwg3ff0YSekoeS1vv57lEMJPsa
YpCu8vEHQY9oxWgE7FARtRfMpoorOz63NPGEWrMAcBOVoC02/Yq8UGQ+LlR5
7MtaGZnjnjVbU5kap59Ub3MUp2oUtcUiUb8OXCWju3I9Q/0Of5ETArMRGr5Y
ghHCi+wRVeBooef+WVblwwLzc0NbOwZfA9B7sRqEEbSDZRY45zWX1BSmIJEw
13J/tIVRf5D7r0SIgRefrl/TjtetMxBTj1o7snIDVnPCzURtGUlDOa340PX6
BWPtKPetVd4CXoumgRVjFgSEVh+QQ23Hnf4wysK6USOoZdAQPFGGSGprv7Xr
jHpDe+4fKrpEtYJHlEZ4gNT7nsRVDRRjafcnNUfI4nn3jzzJGGz9YQm/lXPO
KeSyU8BmLaU35YvuXs/SGcRKE59TLKWGzgAgfs8HeS7OqmyRtRDKHHG+nfty
m0v0nntmRRtj1PNCBN9WRVzwKLZ0Ly4QkFd0dVzHxQAFOIsGw7nX8WLnemyt
NEuc45/mrqN1lUCfHO/zNqdqn5XB9arPGN6OASZb4A1zoX6FzxCLPdnVuONr
u2K75MZAhQcMWLXMuEefEPBqPy5+qqfY9hhCGHKbzVfnzZTCfVaL8TaPP+gL
YeH01Bgr2jZDXaSxEl5dDDOET825H8emkF3XB5XRnBWnbvlwaBFYrQy6ZQKO
sDll5ZSjAyjgiqPLTkereJvxvggO21df1sVJx4hY4Z7Fdk+d9VMr4crZfGzK
zPI2KV8jRZrfLgvoYTpPp9UOaiiTIMLd6NHM+fZjOagTgQ93jCKTR9h1mkNf
SNOhJ0fND0FTSlof4jp5fwIJ3R8e6P+XTLlUgTVQofpLSTN/wad8l9qikrXg
o5WBJwKd2KFqeNrJU7B1GaAm4aVLw598h/ibb+ixx7rPxqum365EXzUzy1o7
2mAT7PLCeWcUZZbOpbJFLcvmSXRDGUbH7xiVqp/GBmEHKZtZ6KfSrANzmj8A
OxBmtdnPtIgt0j+Kf+DicGiKpsYw1+HwwTY1hf6uA1cZg1RlP+mF6VFB14yI
rMW82///g5fR7dcIqI+VIGD0pp1m9hPxLULMQmt38VHV5lceSgH1+II2DM9l
nj5smuTPklva7O2wYFsQxwI7hYJL9QxnLWbMDwDXrhF90bib1/7SJ89cmPiY
HeOG+YbGgI23WH32S7u2BbillByBOOrioJQO0XJIFMZz/FvwHHB2Ewpvwmqs
JKQsRKsQX62Df/zuhwCxg3IuXbFgd77rATz/aTf4lgQOBWQQeiz5PCwi/t2P
rbKXbTOYkDfp/YP9mkAkXbok08pdHLkewVmDhdoEapDpuiMjVKgF56oBjTT3
ECcGSs0x21yK0OfX8iUF1bBptXDAUQ9cGy54Q1oYqpdN0vDIAf68LovyLwql
a/LkM+9LXPdPtAAPlSmKKoEBFUWO+xbLavzQIpEJLEghO4845RFqjieB6K/v
0sLSWmB+0Pc0sdDaXaYbEfcSOAsJ9dYlaqR6CH+gxCwQXVOtExLeUzJc/gU/
NsDAvD8Nrq1ulSm4fXTTG3ebV/OPFIAl23tqp8GPfbQRgKBOOuPd4RqbhlAp
VX6jRtpnRRThi1E8q9Q2iydBkRXPpctRaDSLaLrppJu/AO0L3JXP4x0eBrAm
c8Zqp+5FlvMnAuYGBd4Ms5LFJ1UgLzT/DGz3qnU2KaRuXRY7/KBXL7wfH4/l
gXS3s+8bcJ2J8qJ6Ra+kJ9hzRAegMLZ8QPPggjB0abzS134EDiudQKf2JXGf
mXdJJU8gq+7mIzuQNB5yLL8nl3lL3epeCtJAVRP3vC62okr3sXeh83zUTGkn
5VvDnZmWii9kGWMFbS2Y7yb9QwLirh638UpMQABnuO/PTLJTSHTK79fWS1U+
fL2LL1KyC/7AFUFPEEqgt2J5+m+LyBkJ8xV1zXrVDVJIE0bde0sWtyPg55HT
KtQEtBvN01n998mys269/7m3Qiph4iBEooYUJ6XW10OIJ2igpnSf1Ervx25T
t/NtaZ0ZdsK8/Rh+RgZGK06p/bBhFA+Dp9MXjFWQ3VcL6oKmVvy35D5FZFm3
P2IMjVJZKHdMsSGvHQUR9ViZMHL3gy1VfIjpUksROU/SETPXupMoxCcHVjCx
40+G07cwXbnHvjqUOQv+Yc8dKA9gU/eXdjfc2Rl5NgRf8Q7VFqq0mqOsKWuJ
XTR5cTbuBOJDbNxyTRPpg2rjFtSfpVVW+qcO3TMd7l8spwQ7DL7aflQvcKEt
MHXgf9r9sk8tEoD4GjKFMQZoBoFzDScrOsRL7/Rr1C3+LOxxkWPJv5pYJ4uo
bDdwrjdeloQJv19uoyLr+xwn9/keZLY/6EJaYX6higSSWP7s11CgIjJSrogw
PmR4sK/dYW3JzSBAOE6Et8acSVhvMsRSp9Yn8vjvjvuO3m8WqaTbNlrw+79N
cZqF4ooYKhT1z0EFMzSObNQRev09olD2OcKIgIeztaxqZLNIeTPFzf5pHZya
kazC+970W8F+sveBusD68X6SicXlZyo4EQcXfaARs8JB+XjssU/H0Dta+Yqy
yfewdZ21jySQb2xq4OdgIIoMX83cVj0MmddKbhzU+JH5oWDCEdwTwARdBuAV
I/JB4GdgFtZ0njXWWIFBUbPA9blcAJE27B1WP+sVSJXHt/GQAUuFcV0T1G9F
Ce+FiM79OpMirLufywUESdnennWaZijtFqgL0h+aWDGRsdOPaaA39dXQk8kv
FXkJkEYuySo0buspENB4mIJM3wF739QmiUL2bwr/YXZHx5qK4k9cbMoT8lZk
m0JWYNpwcTLURnLjtsT4tnxDJpMIWSTjja+OFGkPKReFSBY9edhqNjjHLAk1
1zQQV1HzoCV6NJufQ/YojfvsyFpZuTZ1A4qNOohfonDVXqsKFKfDer6Iufy9
ROuWwf28D1GFbcHwDUgvK7S8IARNsTDYkKqoTPEokOzQd9HEYWnSxldfGM1D
STGtLd7GwQVBp5jVh8/9GqnQiY50nePenEhZFcPO0/Ccqo8PeBWOw2yDld2T
Yt7X3lAqfj4k1aG+AuWpn01VX4tlxUsSGvHlBXrerxNZ3c7X+A50wJas0lgU
pW/ZGSVrTtY6INRlJnbRLsWFMDCHJHkWqg4IHTIVZscHlO/+GSDHJiky3WV6
AUEQ8AiVC7b/Y66gPIqJRdC8dGFRR5xVOZ0Ql0AZ+2fCEckGz0rGkhki2e9R
uHaKkPqH36dVCfYNPkbWhv+xYPgWYFZujR+FGo4GEFK+piXWBAf8gWWruN2n
cCWqO1xQGFG579HSiZUomWvshBItYvJ8oEH2TysPsBnTiYjKCajCiCEjTfn8
7WEAEyoaspiAR70xEHpOFAVH/cdhwpJEBV6VzAo4Rr7aUO3HceiSyI7kJ1lq
b8OL8GTy439F4z5oAJ60TBix0VKkXPKokMz7If6PLYUfIU6oELPe/fS6ejNa
VJmLBxxzg0XMg1e4lER41RRSkhyQy1HYJgQbWCuXbFUXKVX5WZ4EJylxohMK
aoxpXMpZTSv5Ve8LKzQWOO8Wk4TPC9YnaeMbfXiUbvgqe2dZz8p504GfdQ1K
j1VWi+HGNBOiO3DuzwpYEpEbBsZta0ij6GU7Vc5Mim0WNG4/tbkT3/UHOgFF
C0ATri6kGirN75paG/6+fG00AYCOUvvee9GSiQ8zmV4Lpit+dat2pMl9+9g1
lAHdqHiNUfk/bNM6LhVwTPJVElBRPYYcZZaKvSbTQV0TBxlkTP/HXhs4Aw0S
fBttwy0GPZiFtI66qPcLqmaOe1wK1FGi++50kOpbzvdBRWHgJPFDrkiSpkck
+KOTjq4QJvJlM8mh1LR5an4HnHEj6tumI/mtBGnzoE/Rz16JbBN652cqQznX
555m6GOKL5EnWser43+rJjg7jOqTIHWtten4ZeHCgHLJf5B8HgvDOFay7Bam
nupohZcpnuDULdGyYqSO2cZ1UdbVnvFrFxmZxnEKcGkssAy0nLnbbrvxRX6N
QvLzJNy1WwsRe+8zGWp9iPVS/3Do2XcpZOJAh7/8xqH9zp/y5CVMVATjj6EU
C5e5XHa/JY2gRMIF4F9hMzwVcr2UBzBaOgoROeRnpIFUJThtktrQy/O/JPCG
q15Am2X9cGw30q/Lyn0ntHt6Qa9DsMFha/yv/MIK01KH5rJU8BW50f9JlqeD
fBKmLDgnhmdx6O7PzMCMO3BAuzhEHatpcqEF/q0OGvj9aaZ4ZJ3KN2Ldn5VY
FY+XUjc8nSSWLgMYpTVnCvLwQVi7O/tKQ8jmkEs8nbT12BXgH/YqtloAHVqW
ad31SxFduI/r40/2sj1yYwru14A8N/rK+9TEmPhwzK1NGwYZH3Af0xzyQWOw
cLR/pZTfRfkv7pYYn/cotpnP7gmLOPeeLZ2eU0rCJ/Sqxx8wJx7b1fdafrTy
9Gwx5LzCbfwGEIh3T8N/xveP+Rii4ljmclETi97/9gycq70H+fsiYGDzNoPR
8i5VGE54c8qFV/1YihvkMg3UyKsP2+hNQ5TUL2MEmmKCq0AkHPkHIVa0tkZ3
zZffabO91203qjp16TR1hsgXOwE3fuAgKS6nD6wUCdZwy9Q7xJ1EXP43u1eb
kF08r0MMr1P6TvW0CFXQZP3/dBkinDP0d8vwB0JLLZhvjt4qOLyZHYm8ImH8
+J/mfcjimItxuSDhshdgq782LW/Ha2tFv6GxUt3JZqEzV7aKfGisD4hS4KMa
x3GlPF+W7SFDI3Xg89n7bcSZK/svAiGVxYTnB4tSiLF/UmdIT//83rvweJ/J
W1NTeyfgslVBBnZdxG0EVvsxH3PtnMNiL5hVYnTEbScLHqzsHmuiOonKkuj5
tXGx723iIfBr+8La8u5NkEdSYMJ9DBf8Txczranu3reGfD0FskHJYw7byNzV
ZyK1SyhxwN3sH4wQZvhKkzxWgDpkX9xFY7cnqLmr88harjUoDBcoWGb2ylI3
ahGmyP3sLXEKaco4Bim5GJ6W0q8lUa80JXXopvKud2mk5hpyYZhUqGCTIXEm
nJYc2qOLHze99w/2ul9snGHeSQNd9B7XYP8k4XF+GUePCuF/cf286HktStnu
kILVWT32T9GXKZwbrX49xOg1cOhswrjWxgbj03V2XW8pVY/WytUexwk1eZzQ
6QGDYTze+4tSBtMMB4Vo7QF4u1Rn3HSU1up+n/mmnK4xP2IaufB0Y3ox+Czi
zQ19Sr8yBKCUVAuG1Hrkfx42IBCsYIEh/v5eQcwaKPUBARHsDf6yGaG5rL5p
515/xi2dgSWUP+8SkVLzUzzgj29uLmNhGW37ZHeIDCqcDM4vDObyLPc2fMor
gHzjBYZHJXp2D7eb7gL9tTdmsY3NWaZEvNxnNgKwPobB5dofJF9g1IpgbEPS
1+T/W3R5T3mRP5YynVXzPxSB0NX0QBFjYZsJVAXMeGXCktXGzdIzB748T24D
bTdc8nEiKDoKNim7pGRIHMCXM1U9wWkCUh23lu5lTiT2cxdkNReCKd3HOWL2
BlTw0M5y0w+WJ56KzhvzpvDA5IW/C9FM2ZkI9cjoVJzIwXQumPtusYUp3d4c
3qFKnFlFkvUKPwLaQzj6G33YM/QeGM3fmC+YFnxbMHF7mOEX/3+CovBDnYBa
yQdYxfqPJtq1G5oIZv5FaE5R5urumkPpCwuC+F8vZtSN6bu400cO5TzLxnCN
lX5pJU4ONPlIwHg590guBbEy4kuuB8QRo6dlSNlodB7D2CYLldpKYuHybcpt
ET62o1k0VSjP0pzZ71iCi4mVoRAGKqizGQNWjq3a4IIpDrC1d021+K+75mGb
rQiMdBLkz98fWkMu/1WamLYrz+LVMH3JkwFYWIB74lSHYXLI40Utlyq4PR0Z
0DAHPUDdA4w0DRhwna00L2un7CaHIljn+mekY817SFdLo0/tfucxLAfZvzXr
+ACvPoEXMhcZb3NRCLY1svhp5gzU3iLwfJu2EDbBH/yFoGXkDE74yYIW3cDS
lC6K/hJd/kewNYfF3VHWNVLYT+MCmYJCl6rLwjZpVdEB1kFp6E8ZqlwG+9zg
qoSl/VihVlhs5J9z7+29lzOHu9dOHqGYbz3IrtNDRDj6piOMqDIEsnRndAEz
7qa2GY+WtsGy6qB26PNBqqwD+wea3iaC5TCsZbdpyP58n42isFI7HAUo2xMJ
hlqgrkjaZ1UGr1KyiPJLiaRl4TeyTsOWWLhIlqBK66x7lt3Xt4IBHLyVVnmm
WAGvBNjYXkepBlYfkIVuvkIGrnFNRfMZ1sRqaE14kBNfoZOGBY8VjkkSdfs8
QEAddIVq3Ik/j8Hepyad9uddwXfgb20/CJwQ75m2WV00h0mAlS8zI0nzzb5a
qmu74v1lylX73BE4cMjRq5m5esVY3URCNeojpnQYrZ0iJ1GOkUAn9PzgUA0W
CtTxNmrd7yPAuYPWVNpWAjhCIKl1M6iK6TfhwNEkmJvI/NtRo7V2tEjA/6nN
KQQccQWpyV4AJaaOvfsrIw8+y46Mb7KUf7/b6vY9gpfO+gLV2TObtRkoaex1
GSSSvpAeM5QJoUoAzINTIpkVvaNzlqpRzw4QPDyhOBaqTbknloTk82GwgZpb
x/SMGvkyxPZ4QjVHQvAu/RY2x9CBkMKXSW8zE6cfN5JKBZz29cWsfTEN9Ehi
omfmdkgUMR2/Kq9a/X9XbY6k3ZPKbQnUpB3JNh6TbhgUgX4YswRGg/Q7AqwW
jW6OiuoZZuKmPdlYHFr9izKSTE+K0cHEpoY/vayoOs6HJOofXI+AjTQka1J7
wTfIXHuVKjLfE7LbujrDNYbtpbmGujGqkzpl5WmXPCo07rU2BYLi1F5Q535F
sy5BA8M1xiP02tdesOWQ6RSUaONjpYXeiOxllUo9iYX9JeVOxsZ87fTU/76S
F+cS7XV0hNzSieumh7dKINHl0NO4OzyULPI69uaL2wvN+x/RTbTZWtXAqq22
PbleHzh0136xp81Of0w1Iijkef4scfTpvP+ypWWL8K0YqkBZXRfhLshs6ppT
HXKEclWYsmbslGjurSSmxHlwKc8n/xqAwsHxw8R2KVSPpWklMeRXhTZ7JDtc
ZkzszwduFLP+3IJZ+6QPbdW0w7EC4rZxGGHkJ0MNtShnFIaEoa/lS6SWAHOj
03Zl8PWG3eMRQf7pfK7NjTjlYmESwM43YXFI2aGe39knZAQ8P56RpF9HFxlv
7Fug7Hf7pthxSPMdqqzrimnNLFUAoV4ItHu2QEiSPd+RF/Iu9wRXwZfXcrcy
S2st1zWNjUuphLCxbZQhd1jO1fXnfbmQ1mvcFR7CLIFW4TC2pBgIvygo5fIe
/t01JiYTUUIY966+sm6hnWdwLXhlT4Jat3ejYZj6YV3pfL2oBffZCqjuaojv
NYHZiERr9/3SD/Jnc8lkh4RqS17aREZ5hQgFkaSDjCTm8stp9te4MyOgN62J
5B5wkfnqW+H5ogrvr7CKWk8nPIocd0/IP1wZ5/p4zPGJMJZ3P9s7BHDnJRLg
0kkiucA3zkFyw5pfs6uWPB+KhxqEMhv0e7JXXviCSzqCbI8/TtYlk8KHAxUP
JtdHnfgFtB++UnOHlxURFUhRgB6R/EtSbXne0Tbuu8jw+iCde8Ni+pKXTnJP
0LffvM6qhblZMi5IM+tb66GeTXGFQWZwxtifQfo9oULt+rAAqtUpv09VtPIF
LCskfiuUiloMbusBDIzQTEU0Rai8yT8SLifD6BOGaxgVQmo7IxRs+xgTPocd
wzLh24qD8LsPDqTA+FXSZasGvDebOMNgbymeZf/nEDnYnXeY48opsggS9Q28
zKF3MM35+3aiM4nlQvUDOA8c0hEZKV7jGv7jZuMklUtD2n5ZFD9sGVpZVEqs
MKzvw8CBPsgUdSwL0IKz1s3CCQCw+47IsnJwZU0zJuQNlQI3gBweAr/Kaptw
oBACQYVokiuaxbx07BpmuOFrF0MYT0I6m7nOL1t2ly1ebCFMz6I1OawK4Yst
B4AVYt3aBfz+vfNc7UoB2onO9egPB92pEVreCjobeoRYU4xMzo5FGIULjv3n
ZV/zxy7OvD4cmXME1W7jg56jgBwcLOXKTVfl9q+1XL7rP4M1joCwzk3YDV0B
U+4TuA7bkDzhmZxxzvrfd00TT1kqrVsaBvZ1GTc5K7epuWLbiSlrMP2p4wAJ
NVoc+XV4uIt5hfIY9xZuqVpnZ7YBHvD7UiQGtd/t7xkdYGWKlUa2Ox7w9CWF
6tkpY2CjOLcLwS1GwJdL4HW6374nv7hOMOfZDVAZg6eiUKsUi59IBsv2p/nd
kVA4TGUgtLu6R8n2sCaV+oCsQABGipWSZUyCuUxNCsPqWjN8tAbAW0qHQ+aN
NgVEYK44RiKEJ6frYVWpTGrcRAy/F6RoSXLzdwfHklURV2Zjv8taawBs1C3H
DTaWcVNpX4H+l8wxnpocWVQhQdHBbOCdVn56EGNtlPjb9ULOhpKHZ1HymKfI
uYJUIk6aYH5pvJ94j7qWk1RKhPC5iEkVN1h05m3CjyMfl0YZJr9lwXsRGCUd
GENSDCD7vOxpnSb9brdyO5uDVmR0Qsl/xXL9DS64lRMfGnOdryO4X4q6ALqa
2H3AnMzb2gvgWlRKVzMx7Lr/x6gJkwTcpm97VRmTcwnGmJNv3vrW0rgV3rBF
1EPh1+Uy6up3q5baCP0JcZ6ykqxWfw2uBr9UMpid73YXSkl1cU84HjiE/V+L
y0TfdZ8oXCW6UOIC6IIFnIQJeLvLDeBu6nrQs0U3dE068xDEMel9YTkT7rXm
vKrWMKdqyE7UI/yfzNjMRNCGsjiB7KMcuow8QHdmXmQvgEaCt6o6E0Uv/W6Y
+0D0NX9PaBTh588JXwJHus210nCBeDkNdvfomD7vUBj8KgrgRAIKfevf0+vl
ej+VNFRHFfxxxFdf04XyvV3fuw52Y4ISbdKa3kCPbL5eMxKl0Pp0Dcngg1qv
/628glzR4JLsIHU2QLD6R7ar0hbZ74SbPureR/D/wB4lTts5ji3qdDD8Z32O
VlKUBgJJZ1AWGO9pkic/4kotEmZyWCRvzCgyqCgm0twwLoeXNLe6eJcxRQZo
PmzRdjgX08KWzk8BAHI0KIpFHtUFN8viZTOIDJZxxTIKScmU7Q8WFjwC21y5
v76SmZ3NBpobWbKEzhUrBdafTbDRZde/E7X9qMZU67WYVgQRZqY7Fy1UTTEM
SwkfJJJ/4dt+/sbdIOFNms3PxBVO4W+G5wlhkHl1myWkLxIJEygCSR9jJoEc
Mm2m4xy67afHrCeHJJNLfVvk01Dzvuxmwx9firWbEleKy41f2MsqUuu1UCz3
NRHjpJsfVuyGrQA3G4bCb/LPEu0uSPbQ2bVMlTPdssUmv/hIR3EK5Wek8sRd
DH6JqjXhoQH6Ud80pjIeviK3nlEWMLizKJabiS87KEwBZWPrxl2ebIJzAbRb
/I27P3tbkzPtW26QTTJ5j/iSkjnwL7otB7k/m+sTUhw07qfBoMo9R47npw5A
IJAb/CAljcSx7fogSXBIv6fQ1KnLkWj9VNtwbcA3TMO6lZ2IFZ6QmDmUILQJ
sFVU3vkTPXOYDmxsN6FNKWNDbYaXDabDCWpDcYul3lMDaE02bgjffJ8iM/Lw
QPH+6JMY0gLMF2hqlK3VuzY8QibzimqTPfxXOLJKbEDzM9qANIn4POPTQ5vM
wYZKxvH8PWnx0M9beSVC5H7RvVaodJOLRA6+wKGFu0/xzRBMdj2mYZLhddP3
4ljdNIf6PwgKPj6IUApxh+QdoWOQN+n8Z5YyjWPU7Y9bku6Fzn78UV0A7Plk
SuL2JwSlUV5OjplUg4x/eKQvjXlQh1cVXttd7uKl2ljHdM9nMMQJN+4vB0oI
UX90sFyqEy0XbTPWeZLxBbBZSKYOOFwV5saXuqxSBDwgsX/9GhOZLLDhzl9q
1pykGNnpzGwOdSPgvKqN5AKFIkCMCZ5i2Ft81wtNSnFSH3RcCet0CK86nsCA
7ANqGsfsUb2l3kiEnGTgYTZ7VZ7AnG0+ROYXjYJQ0JNVOg9U1eYh2NtfgCBY
uViNNTQeRnDvPbQrsN5M8WDJxzT+IIWN6XB4ZN0kt5sSQ7SxsosL3qwFPn9c
vJTU8XWLn/9kR8JIlt9JbIlvnRhFy96BuXFGXfSRuZyC0TJY3BdXqSfZkAjq
zbjWgNQpuTYc2ROVhfHmc/0S5ZOSj9J5BnhRhjsPVLOjE8tAj4YwZNG6l7Eq
j2cryxNjmAHrIa9Z0gwenDNDSugKyhNkfLsZ9Cf8H0iB2wvZ0NbiI+QHtuvY
avy767bIpoXfS5kF3h90yFV7ShY+lU15QqKlRguCLTjAHG2hO4CBf1CJ3zJ3
Q1WbSjbF4f2I75GyhX6XhwcDX5Mn+CvNfWjmG7Y3yetrfi/MfVCAQsxLzo2n
X5G3ysNDGOgQOJA4LboSMIGluCs06NjSMhXFzF3pM+ejYnhhFRAO5v48T5b6
/D+eOLtqciGrSAa66dCzNZCre/ZHE4bqHDBN6Mu+qzyJ+FfkJNaTn6X1z8+w
wpybHBLpbmshZBn5FwzlRdNUg/SVnrbEtg0X+vVNZXYWA58SY6bREQoIqdHQ
+wty8hOCuMNhJQXX4RXdyKgb5s/zo2PyMJJ0SVIjgC6SrHV09jhwOo8SPplt
5/YrHG/KIHfKkGme3Xp61fBBneyHvtCrleUdyrAclOpYF3gn0A1dJIMVQEnB
7JPeifwVLIH8AqLcnNQ3q705YDUXMzXT75sWjmny8Y1r4X7MMzokYuW9U8Ie
1Oviu4r5fsic1Jw4LZlR5jIbp7ZhyhCfREn+sd1kenjSuls9cA/cRdhdV6Qz
J+5gBjdlsAuEOiUHoYIikhsOywWT+GZT2SPwrzLlc2sOCP2yd5KdbTv3NnE+
RrbUiQnL1dUhmw5IYildF8oU7RZVVxhb1zAtFNYiQcgUGF8vMQCMpO1Ye+A1
thEfeUbi+tQK1ze8am+EGe1KoUqxQSioqdiCs1GDu16xCnGOsByBM9KnYpzg
s8KBwjJ2sN6fpSyvklhg+sc+uGU3HtVfGiFXiLPz2uLOvSCE1ZArGyUjehuO
s40X8ug2Q8aBph9P3Nv+rO+TtVWu4lp6qkdn7P+w45tZbOsq3fYfLVCqtP2K
BmXM0KZvPVUPAi8nYi+2SgI8RiZLwj5Jei7gJTC/Vpdx17untLvZQKtwV80U
cstmBXqMv5JGcaYh6t9FHj2E5akua95MgOv/6Gq2vKFMK3cL0FVKXGIiC53m
196tebzuaF7NC/Dz/N46eiozEL6fexm4D5ENV1y3bxS7NwKVv6a09Dl2om9B
ycwIDWdeouRTc0WffaAhAfj7MnyUrngscr64P5bD5c1v4PAaj+TnpRx8kdG/
lkCb+6vkAUD879sKB4ymFF6SfTKL7vE4+zLcIYSlkiemYTOWrarsFulqcNpR
Joeg8apScLE4oOlaW6O4SwvQk/y33va5K+EXRyiER1pXAMqfbZ0p9v3XnpGI
TtsH2QUJtjow70MXjqY+Mtg+vYObdr3Q030P2+XD1+RkIG6Dtqn/Om0yhpHE
QDWh6olcTmVAufjTdztk/dIcR5AX+tQIEzvhq60ERsEkwxxP67+TMJ+JOeYw
5SUNnmxms64cRK+lfXBeNbt1ZxuNp4fpsICd2aL3D33nVM4Efap+dLz10Iqf
KZCSld7voQ9sca72MgUfAPZ5JpBEN3yisTyFOhdGuyeELg0b7D6z0RwfkSAA
69LOdGCG/9TcMrLQJ5qbH/JAj8XBmHHMhMA3xjKQ/T+UyY1k6iN27AOEaKp8
LmKrg0iTM/aaum96hYfhQua6vLVBAcD5VAi/d5+lK2Is7MqKSC8oqshvXunw
qhtkWVPeeW+njm7ovnvRmClLZGiv2IZYQpiiedYgRiEmFZyeDl+nPi1YEsRg
ymYkNa6hnFEYXG57HWNkYZg1lBhyINGCAMWTwo5eC9LWr+uzBpBZIL19dzXq
wzubyhsgFTIgATzwsXk0eieeeiv5hC8LXlR+9QzIpZIpW5USkwyGI0POQfsk
NS+GXIWBacvCpi43m6zY7vwnkGYw1MdNBzl2zbBNgZ5IgWTskrbssqtEvyQe
DVdWTe7Vgs+pGo7vFEYK9HaO7X2PrWeM2dyh78jaTIkfGFubyxDCvrfD5bcY
gaooKo28SCi3iZNYES+9RKVV/QTY7vw9p2wX7HKL3yZgwJqMAYnW4CondcNH
RyM6wCO7DSu9e7JXz1y3dkgyw3wx4hJRl84xl5QqaV9EMJg9WTgsANXsx9Hk
riGRnGWRIQLZ4/fvOJXinjDzAK4JYH0zUjsrnFQsFO4sZfF8UVAdKXnyO0/f
KCfMDt/v+45Y2Mv1qmMwmSi3A+F0NBHEIInyj3M02ZfUs5m82OTyRbf7o5Rw
KeEaDBHK7ux/jbcYUdkXG2XkIzxso4dPXg6IkoBkfRqMGKBlKbGc+LLNHERN
PuJzvYPwxF3vdkFaW5ELQxCvIQg70hNPonZzcjIElky34ptXKfRrvfyjYy3Y
Ib67EQfmtn5SOdkQoBld2x1CQKGGsxTtu9J2cHYxWuDRzEYOl2ZBME9sAxlb
sbN/1a4McKr0aCF4m24jrICsz7H7BhJAgFaIB6Vp2FJyD/kU9ExmMfLii53N
nqhVhx+VPDZGr3sbCZJCGCpvl4lKXuuwMa9yr1EV31lXQxdUKPLjNdwQNWq0
s6Qrph/HOFoEB/p2jpgV4QF1JXtpHWIk3zc+La7taPAvIihgCodCzYvV+e/5
sRnAnHD9Mgnms3MUa4TOg3D5VDnAs5kOSHbFd//BqnnOxDPpuwQiLixMm6dj
NmjpDBaz3Y7N3gV7xVLLLrazFW9edtCdd9bUFZ08eW4jphMln/kAMzYjlOZx
EPRC/HUtos67tyZHU1ogLeXdnQ/8BtdmktkaWPIPjf3gEQsdM/7rU3MarWP/
MJM/BCt3qJzR0LeMwaZ6a4/cI+R2HrMpPiS1pA664lTVTghgucvY6Ycv4QhK
hZTQgrj3ft/ASqOYC8V5uOk8pQtz2UQrcS73CO4Rlq7PVOT7G2XS+8uo8NFn
xl1HuusI34yhaRy4xoucI2/+UKtty66lkKPphIOvXOyOn4517xLP0SV2QW1r
xdWzHxG6LU4v/YZecpNd2Y0bNDLfsn3RbzvVyjJJjq19oaE09JyFwWRGZgok
rfMURo2M6vZDECpBKdMjmOEK/JbGJQEcM8hFmy5rJo4+Z6B+m5bzv7BgjVnv
PVqW5AvlO1gqvARHhtPCbWwEyr+GF0UX5Jdk0f42xbHlkeTgimXcVoPN0zEL
GFduxJxqIWGtu6vpEy29jjOHmzSbMyaFfOn7xhhFPd/40lImbolpR/uDuTAK
4xbn1MH+Y6eVqC4wzNWmCTwi+OuPdwxwcZihkjaEc5KuJIcTRhDbFszGFslf
tF5P5syOxEjw7csPJwH2hj3pqSxPB+TtHqzreOhYyC//Hjq9RFyaKaOqYIgT
seSuxzlb+RZYtLcpx9xDxGO6CBBit4XQXmKuY3TOs3wcb3eJe7WLs9Mvb2V9
pRC8HbUwdWICzkw6OPy2U7eqyIlzGAV0/1uVs8e7eD2ru6Gci5HlSfahnZ2F
oqH+ZANu1A+Z7FpizCjfUF5ThH9FbE06mrw3BF5EzdCNupashQQowjVrLXPT
Qng2wvE5qiEEaThKMC2Pab4SeFveKXs8I0AedeFhPfP9ay9R7cvoWBshEOu9
lZkT0749rosElgCaw/mcDtTqVbqhmKhLFv6rN3MgFX5pAj697mnh+v1zj0yH
U+UHqluLGmjycHtAURouofffAM5eda3HSSWOb07lSm/5E3ISD7O2LFHlyYYB
5qxmhXaxwJXQ3nN7YlIpoKttJYVB5xdyMgpl3DNZg5q7aiRG8keDG/6edrbg
cV8tJlhZJj3vNkHTrtDflAWHkI/uOVPS92xgZyBt0YVeU/VySuacARxrMQYO
SdqcixuMEyUYd9DoC0utD2yM2QTVHXr9y4j39Kga7QPRG9Sm7pxswPqp+k8Y
f6mAEZq/cHUwxbetCf+MQu8BovFZ7eYZv0nkAK0T95ffOLLdfUnQAz2POVkd
fNL93epLM9jP5VUW904JT4kl9xj1hNWSuh8gOWEdJ5bOYmNf5Ba6QzTCoAvG
LY75kIQaoc2GJE3kkGRQI2ubcx20MoMP/u3R3rGsSPhneYgp9KL3exJgaNnl
HEPAQYWoR44hXZ+bFs76gn/adkKiX2g9Qbnb9XCjU6UZP4V7yYWW9NdHROQ6
UcVMZsWWkhP/6j3BAkpQERNMPqZ6rAsa52rcVJvSyF1OMhJorcNfhV2CoMG+
T59URsQsQ56eHWk/NCj9oKMfppCIoVeTn94PzV7GrJd4d5pMcZtMC23JlNHR
NwJiUrGQeD+eZi3s7nF30oColyRwRuwiTaaS1kH6K7fnSwOMKFipP0GXJ50r
LdsgpkrwDDGvflI0FPrOSRGEo2/m9YsFWS11zlPm6iWgoDJsdH2JpGa84ND4
MndQ0pqx5pyZW6pcTHH9x6hno1zm/WRNKJL4XuW9r2T3VbBfT2ZX86Pcxq5X
GIF5eOLbO2gkqS3RWXuAzLZXqbOvdn3D9EAMHsdgXrgUANiaojlvL3Fz6W5q
CplMa2tW+pWGuLYSq5y1iJYbRGkHtpfbE+kVclphMjqNwGJvZM7sMscLLX8y
AdQPCJUMo6UARvUGhoZWiSIaYvkqDxmfsRL8mLlnHAWJUXn0tEEJeunJem1W
OpHLAUt2uneH7EGz60wuMvkLik/mKEakWi93tl66m34bNSe7AlyW+7rs8diq
zmq86FTw4GsqRRRzw3/FwxmneuNzZECo3Btthr35Wu2ci1/Z+i6cK4SkWKo6
qcqXoDZAubmgZZEVav60fWlU+QLjepJ1wjOBxtH1ZcpH3tBoQABFPwlRuxLn
hyYfthzeMMjTbrNfJWDF86fH+zpoot5xWZ8A+MYMKE/JIYVmA6+689KDtgEa
eGgdsk9xTfxictid3/Is763aj5+Um6v7VS/QE/4rURhXnUbjmxHgGJGQK7iU
ckpbpHuTruRsBNFdga+K0W4qG9Ul83xsTtDz751S1eD3KigelGraQNHB/L/M
ia8ARqCYeeykAGYkEYR/nCe14EOu4AOF5MTAN6vAT/WtqbJ2r06ulggNyI1O
LXGhDncOZ9a5bXhBvuUzYn8DRgA4tc+Jh1ExBmVAvv6j7mJPgKPX0rflw/Zm
XTTLJuIhvPZy9iFQqU62UAT+byvTRvlOjmT2KL9GtCeqEGNlO3RygFWhL/yf
tzhPhVKU8k6eo3j4/Rp7rRcAzUFD5PbR3E30bg/AHknyiL4CDPL47nfJ9JaI
UfUu7VA1KV9SSeQPiHhaWE3Uknk1uqwjw3OGfBY1Z1I7p4l6GdHALlLxDOUu
bulJ1y1/WVAEplCynu2DEf9e2V1s1jVA26JcW0LPR6m9UDG6CK4M0m4lHy+7
DR60t7PN7p6/l/Rb0tdu4ve/MgzDyhCempXYMvwzxYHO6u+oVZDeYtCd6Au7
0r5MbnOScaiQzkxMeANFWNGoXz5Qh/Xs0Q2ASf05Xcv7ebu16vY0Eip2qmHz
Wx2ldkiLQ3ydZWPPRhoseD7rxM6KMQ5MTJ+bZNW1R7tO87dTn8o42A4CwW+d
MPJDaG2EGPvQQdFhucQgOznF5371c/VzNABNOK53eyUxLFoW77NBOgCyXD9E
Y2per0kdJUrvLg2qs+sCBeBqMBGjtktodidhL/0sP4n9+/nxvPzmhn0MnR9U
f/LeKBr3dpaimN61liLyvp7qe8aaabfrN7+vjh0um0FqpOtdGeAK/TtNYcyI
g8vWA6m5a8SAEj4PVlEFOdMsxyUJ4SjeVArNHIzTeP//sRCKobjYTq6GVz3Z
TVTVueF+jgXM751VQkrKBJn2dPHGr7VCSQFelax+8rttL9rYHwVcHCdSfe5N
jiGniGi8OZpCzEhr8WowYMuPTZNcMRrty+hO/osv9ZOa7tehr4k+0Adr/7GZ
HQnTqPFDCm0xq8X/r3BZTzx9KvWofuyo4+WAkrAZldAjQJTiigd6WSuG1P2S
AjOEVxLhp4bxxTRR5Yss/DJafWe/xC/rR2dKTmsopAgXtYeGCvjLtGA6aMqy
407yijnbbJDJu0Kptjf09KCh8AOBX64olnBJ3mk4ZxE0Yn5hGL4bzojURGkX
Q+N4izLzRNXPbs7m4ScWA1V57KKzONQyEwl5uTugAfMRlnbl+jgA0tvJVkJ6
SYB7faX07HfiXImro3IqhQDdK7xj+JUJrVBhTGrYXSIFT7DAaZIJK9vcmbk8
Te0aztSlvgs77728nPTlbXzrwATPywQVpTvOlG00xlFqSPtRHBc1wpNdXYIs
lFOE8hoIOeYvbc5o/F7CU43ahM+L8Si/s4LlSwh7rbs2onvldXRFsMyoaNIo
fp/YgFF64uZysEwAsZIBtmEvoCcBxhirJlBA7yP/Pnn3yoTViwjZuXsSalK5
S8Y4Z7WGuEWmU+FY0oQyd3muHnqxaZpntsG3XR18o1hNjnizAQY1Y/jbIhUH
6JD1q2C7bPrHnrjJ+3KbErbbVaDuWpPrqDlbRZ+TwIUkXJJde43ZDfq8EfWO
Ab7c+qadAEWW5jMDWF8JFTD9S1CrR9DzB8EGUo3Tv2EL+BlVJJgw66lpizBz
vzVwWIVIDzFonQUyOB8AmNihBUukE1T6ZZSCtaPGK1jDZxjzW8T7Yrv1cLKT
S3C1536oEkkZ4U0PVYb0yjqnoy2VMGdSymy3otEinWafUWRDriswyIgiw6Fw
rlsJH3CEpUDJCvOZKoLGJFU2e24PYo0I2arGrbDFbWdZLnJHwLeMcFBQEthu
f+CYNjbhqu+/Z+dr1G/F8xXSVbNKJjZWniCJGcaNR+50vXuVxVuP0/bSfdC8
hCbQEcKsx2rYyybUHQuQZI2RF5P8zkOgEfhntM9BM/nBTG/LfUwoV+lUHMxL
jM6v3Ibog2tmzMLxhNwWEu153lZFhQ+En/bZr9f+2JoY0rJ/IooogEx6//dA
ig9OoxZ8IVQIXhCpkuFEhkqPJ+ooAbhrFsKEE9PphTTBYsyyDhR2I2fZ2hJk
/GNn6gFK6wRaJe5e1X9YYaGSaR3HXU0iodyhVS5Jj9IPgarsYbJq06ccUrpH
2GP5CvO93KQDjzReNLfjUtTuYfEUHpGXREodTfrAeSop8hvLug0CGsC9VHGx
MV8USw/pFrmlwq5VCgBNy4C9MP8xG7UOpZ8T7q0PUDalv7esVmZjhKRu1n3D
1oatWo0yHjECMfkDCKaFL8/JR0pzJNqTgrOJpkhS1XfiOgUz1yIhgSfrToFD
1Z/GvAmT55Jl3OKOjR7uMZikYaeZWq4eRhaO/k1v3Xiz8ZnOWlJtH7cY2xv1
/9U3BYNd5HkfLtPYnv8HASX+YyujOVuY/5Dl1qUhzRl3UWbcWblWM2yhidYA
sEOA3mMq2LryJLbLaBxpnLWK3c3tkFJly8cAXelQCCSfwLHLAh5a7iQvzak8
Dqtwh9ly283kHZfK/g6lci7K24o70Bx2A0Ox3tpMpYmY4647zx1kTq+WeCri
PqAbFhRhdsLIi9axuzNQw3T/XJdmmvGQh0QZ+z3nALAJfzHbvyJMloGV5hlB
eFOzc1lFOyLv69rh77N1g/OG+hqaiyEircODVVHknwhQ7aZYoJXnT5OdqtP1
xoLoCJCCVDvI6EnQrbExSD1iCR3r3BRafNVP9/SEFBRoTWTRLZjImDlNM9lw
Sco0k/BJ63YGz4N4Zb7mmP5n4zRb9YNkoze5J5neafaP9FOGbesbBTPPZgXN
i6YjVqMLM6+yxvaGPM+8fMAj9z3FqOOhki3dPXftn8r0cb7WwkH224KUyDU3
o9qsPijAAzGgU44CDD4sRCddzw/1Po8f2TKqVt/WVuUMSa7HVDwRdKXrqiB9
z7dD2ecOCe1KRhrLqzZXAgBsnEpY054A2rwD/Ijr/RaQdJcMOE0KC3I5fzGr
fLSXYCx0e8L9w/wIHlB/mVfDOSUZv+FT77yBlly8weZ6lDLM0Rt9KmKgDXqD
Y8su9XM+SFYSdS/+3f36WhnY3orhlncl/P5AkxZNrXMUZACOhaW7Z2ARnbGG
ZmRtVR78isKEyrHPfgSuP0Yz3OfSj8n7eyr4y6yKTiwt8XTY89Ym8qK7lRPA
Hk8egLQJ0anHE92FD7ZSCl8Qx1iBtYGQxtmOIjGLff9Jr0rN+7Nz8+3PAloJ
Pumlr6d5dB+sCM5DB60cVKX8K9UYrwFGU08h/Y+8YP8he2KrKcbZf8SzS2tG
M2zronw7vO4lNcEhLzYZGfHN4nc2jjtcMjHnxJjQsK9/ca4Wubw+Zl8SbcH0
lGwIVJTn7Ew6Ro0G7JDRh4P1rQcO/Kx6K04WqN5jxUSEqoxhWEdVoTfEmgC+
iCxS0npIdQE7iS1afg2g4a2b0hEuiKgaOigAQBw/7c+nkY6HJX53ooY1t3t9
pOwaF7TfXFXfD2de9ATdNHJcAAr3Y5lPGMLB6O/k8wcW/tRiOZtxzFGRFCjI
/6gHEiCvmSF7Cd5X1WLRWqHAm3m2m3awpBVsuxEpN140aeeJkbiJKeoj2EW3
rXSY4sSpB5hcsaFHWQxT4LTh3ciAtJm7bkmRnYVPAmDTqKrxHwlfoFXN+Xj5
9sDSIDtB6fTtOJPoFC7lee9jSnZ3iY5ZGHR8X2AuFdyQbP8w7rGumHUErtRD
p3aBQtqBhMLDP2OGS4Ovxy5xLTfjl488dqBkkYe/F6UrzKGXzrVpc6XqXtSL
FoIFQ/EsPiSgH+J4ZIaaKeFNhnnxV2uuk4PeS4xNxt3JL/6+wmLjrLPPzG4u
OQCCXy55uZLsb4xOb8Tsju+ZsKh6CEOmXG/ryT39QpYsFQ+c6J7O4yKv8uYN
IOdrL8xpi0oKy++uUqpUPRLSXGDSCgz52M6qly/fpzAMEnmvYZvwlEU3lwxS
8VaiKtIP4y2TxG9OyWgOff6IHViwasYC0twinG7F3id372Vt0boHKiPFwEWY
gtJ5PkTPLBqiaOFe8pXSfadpbIyFOm64CCbmNoo1lWsQ8QWnntvvywfKF73n
QoUykXpcOxjiGqxI6HAfCVlDmBlZkAb9tlUreyNgNlGR/02GHioN4VBozseG
cwbSQJLl/U4Q7qMryj7icFPuYMPYbnjTja2GKowAFIHUEDUCHWMI+8L2/Dph
gw1eXMnl+7sXY1iNyly1GylWwGdURS/t9k78aDjMa2DDUKO7iNyaEiHG7f0N
Ngy+WSLmWQWIjR31CLqTYxbvSo8RTPOvvrLYU9lDf4eFx1RehI+ZLdDBdWt3
Gzk+B2F2wWi5EwtF8e2PPKBE9JX1lRZE8Kqc+lbZBkbS43C0VbxJsABNfBG9
upvq25uczIQ2ldoPupHP5vohNTPjoPcSqsjEErICwohXq5vyKXoQFJjBpWGt
bubrg4kXEGXXTlmL+yo4jW2EkcIv5kkBNfMB4Dlqj39SHGJJFgZu6SlKrkDl
hJB7X+q/h+jNsaHp5k8AJ75seyXYtFTk/lXOMKgEDh3XaGGEGD3cMUEJZXjS
z7DkoxBDQaPn8aNP1hp9lG2jeDaOa6eJT+GjSUv6QPXafvgi9i6MQTX7cNnP
AIOvn2hrnf+Pjmr/e6yX38VsWUSxjROQgAAaJYK+OM97eMGalDdNUAF4pjGC
fBn188HtYBHp2AWate1W68t+D0T3fx+i7pBo4c2dGtPLxGpJcJCgCjK0m+VU
rmm5oKyAojP9Izcros+U4E2H65G37yCMG+pFlibDG/7T5aHO6PwpC1l5BxCO
do9RgioTiyiZvxGfgy7GaMsyKThpmTCeYb6xtbyEP7PaZnktH2NNVexuVaHu
g84yyXjlrmgCx25P1ZwffSbo+151WtUC9gCgHILZA2fYF+AYauIzZP2rfpd0
rUz0B4G8lCX4Z+G1NMA6QLHQEv28JChuWjTNzSs5dtJv1GJuDGVLDrvXP4w2
Lc6j+ZTZmLY/Ane2zKCLHI5ajfkO43fulXmdLXS40kCtcLx5UOPiKeVckRwY
dcMnMdZ5mp52ohrORriWXFxX458UEHArtTN364EQDidGDzxnRlZGB/p4Y+P9
F5H44OSFX3UtKIPbMn62ePGgiNeBkO7H4jK1u+V28c3rGk8qrbtc/Ez6+rer
cqdhE975abWb6fix+D7CoNj2dVOTs5kby/3NE/uiMt+HHy1W+NjlslxmXgIL
OouPHi7Gh1OYujXawEwUM6CAlrjbli6DgDlVUP39S0QmnJQ9RhXV9L/rUE2S
FGBy6SRh58w9o+ShsVoGdsiHSDyS4c3IsA92aGw3sbIdBjIyOHIL3lf0EW2e
SBEc/zo1qGo6UMmWMnt06eO1gZTP9+CfFY5RsUBmlkQyQwzvkwYidzfQ1/iI
gMDFoWUp2XxpzXAJDTQEBT3OpSiEU5cGaZE/XjFx4TBumzgXpYO9zqFxFvtu
tA3fqmg3XV3hZCUWtbbMQNe7l9aukcFMxHRwEAr2Lm95ppGcDvPTYXwzxBOk
//OSA4ZTPplsoFgEASFMjaJRpX+5mLjYRGDLvI12zk9WxzcVlE3mObgqL91G
dP76JooZO5eCMFcfRXNRmzOdoh6RD3y8ZL9TtZULba2Ffd9LXDLtMV4uxo/a
GhsBOOEaoqlvRayPK3uzbNeRC2+gLPBV0lGCtGB4lyeWG0VHeZziTBeLklHy
JZFFV9UtMRE4eAeOEHIny779Enzf9U5WSWVIqMJZx7ryTs21boXEwo3f7OHw
ArHUHoanK4dyh29O3ameR6Noe8bw8mooqv87FM+Vt3S415rYF3YthbDekA3T
KbA7S6O11OMNCRv5tslCs+taf8VJ2A1d9Sht+lHgeRsOTRy1eHqWzbBJdR0G
2SjGjLAFnYcj1hhvqT7FghpUqhQyXSFUDqc7Jt/vvDPZ1Me1m6Ftq4kUw9uc
vL4fC6/6BCgksjLsfM8r0OXrNpGFTz4I0iLIdYWmTWfYsFhnmp3LyeoQ+LNh
TlVnN28dE762Af5Qfy0M0V42ScpEjn8Hwf2Bb0Dll00hyQU9lwrwmsoo7s5D
6+vaTZrzlab7tp6HhyHV/Xav1vgBbqHdCNhqdU2OKc5pvHWu97Oe/glp3AbX
QuNhcxBq1WKdByD3PZcKgSZfj1j+wpuXK03++Ns+H0tGYVroezv0y6vr//CC
jRI9Y5cDOGmbtU6LSj4O1+Fgo6f4IaONgzJPR9myPEZy9OqkDmBI+IGh2hkh
9ONTfcC4grWV9rpdqq5h8+hNx/73JBP8cfPFXMlLP/vmJxSLiYbWGb4J/zSQ
1MZoMLFn343D7ULmvI+MD5tFu+Yncbp0DSWXwKJrJpXqgfYYbfpmOlo5lLhl
Oee2fKaRBbvgCQ0h7cdgmav8dkkIKXmyGg2+Lp5q1Dy+vJJXmHbe6Juppcqc
NukKE3yMDsRODn+YquC1FX+oWKn94MN2PGINm9UIOZhsfzplpbqDTdg81psU
ejaFM/ETWVuHxg3QiUgax8ndYLJDS5fnrXSVx2TF3j7sDB3eQ+C2OUpe7aab
Ad1pu0ZXSlODRO094AjF0Mo4vhZI/fcHx/MD4Aw1xQAgRXo1tPM8a6wjMltt
9j47j0i1ApTlcv1ShNfQYMbGYUQwlDHsC9PXh/NIrg9V/5ZvbBRJHL0dNhy3
CKWZTND7bsL9WpZXWcdR8KdOLJBfNZHSmB0AYR9oBIK/8j0LGQ/cJWWTCNOu
cWXDHxL7Xw8jMDpZxkVob88XIS52Nc1YHqZEUaOXS2XuFdq9puhovNlDJgzg
YblwBY7orTP0PETz+4EaRMcu9CpwsJjjAa8z1vXKDg3B+WeRJvysRp1AI/U1
7v6pcWBc9DmrTwBxIhwIEt5+1E1qaxswLx0tZ+sgvoqwjhUiNXT6YjLmb5Uy
Jpx+Jkbgk9efg6T+m2gLvQ2gJ+OXXk3zqUCbAOFVnqAG5LWQ0EAmigctuBCK
P+vFUc6RUgQo0hZx7j3nTB7xrEefJGaEU2ctkSgNlBu1ctJuSbt8EY0v9xzI
sgja1h9kwXnHMg/tDkMEmw5KM5o6H5dR1HMBqwu3sJBl3gCD4AUVyfODuF5A
yFlZ1vDDpKDRQP6gs9yfZhFYM7PbwTa7jCNGfWqV/vwoEQ1H0Q3Ra6jxhJak
oFNhTdygsWUZN8cvcOPjrGJecu5rOgdPYkZZWNU2rVDPvfiiN/WY7zMSBuZ6
+n84xKZ67YHGbGcibvmVwvU3DCx2bvOWtZa/Otf0nxjn8/y24sT0FFCo+6qZ
kB6Z3rGo6gWL+aRykGLnbPX25Rn6X3qHOB5MTccxdWFYn6hBimTenmFHYCix
Vlahl77Lq7vkx3MlksN7v2El0LgHRh6irw20II6jEVG7Fu3JofyUD3gTFPGO
zxDcXJ5aPrk4XnyViRjerX5FAPYP3067aI77ev/VhJ9gsQTEF8NeZFkYi5j/
gJ3h4PyBrYa8/ESZk8NKZK9bpP5zJrEyevrBpf8H+LoWvMTlCnceFMQqSpfB
nUFbRyC5N2gBfP+mJRIsYt90/2i96LC136LFlSbbu5a/9fO/M6xX24XAl8dL
+B2ukUYCU9QGINEps/knszJ9LycGIEmC2ZciXeu7m+vO3+0TTn2jDfqjhkFa
uj7vviqo/J/22T/7KKIwu2LnMHfiLuHCTxvtL0g+bGrRgvyo/I4Od9ivOCCt
wC98s8ZUIMSk1L5pSOINOufuVZotfeC2urRDTMMtlX5bShcRIqHVsElUH5H8
W+CskpOgFnF+AB25kubd7baags7DzOeQn00NphRDkWlZ5pUX2ycYDsNHCxv0
UiAJC5VZLLkjDj87oiLn3Aj9YG+s5g0iMBBijLg5+EVRVjWEE5WcdkJK9tUa
Gh0AGimgyQB8IAGQ/9sDqAKarOXQKDMkaNKHQMLtV5FkvDfpYz2GZRMStgxK
shiHwljuwdBEVb5uNiJFTj6bnchpY4ksD2S2maK73gAHJax/d5Ff9W3lXCcM
nq3cduSItYAEmAjQ9sDFzLVmfpvag5K7ps/wRkmSxUPGrMPy4mO1Y/d1TPWl
n+AelQsz/f3u0fR2ze/cLNvqqgovF8858OSTtTAuE+FuJHtpAgYnOBsSE0GJ
8u2g2x+3iCczPuQqhaQJrGsCyDufapPpm6x8YWQSCqIKCALL34Vv3kS/NabM
YsLUkiquk2rAQZv1tjiBEP6SBU23Dpmyx06Sv5YfzPTfoqLbFGB5yy/8l4J2
+zCqtgVZPFlAL2rqvmX0mlUv8iFxRLQlovE4Gl9bU6dB6gYHSvnfVvmJju54
Ynj8FhcemEHwyULoYK1mHkGwDLFQOSOk6bUs9pUSKINsst4Zx0rgKWVOPXzh
dz7GYOXva/Ts4ShozokGQ674DiuzxG0eXJ6JClk12mYH/+XBZ0PY9fNM+muK
LRPq1AUjT+OrCb1jIcRw/tMr03BCzagUB6p5WNiJmJsewnsHHCzS/iqs4muV
nM2T3GOamiT6Il3HxSFAejdj2tZGxvVUqtIyKIaS3NEm+kyZZKUTpdI4u71M
Hor7xGROazIfdaUuN3a7GLvvDCGnhD4gNIzacnPoUFXwKRQvFvfKH3XHgotm
0rDC8wCewIqhGST48ydxL4BcfK7jeIzkE2rRzlXMFs9rwR5GAchl5qFrbr89
oN0dJBKb6vHRA5tNfzk6JczrTKS8+Vyb/KWuLtks/yVyRs1Y66V60FBchrEd
o3XZ5mhuy2US2uru6Akrkoiq8H8H8c/WFu1oUumt3854Qhr1ZLVTmbVY+dnk
f349IKPxAgLxa4itynpjV9SXCO9YZUGglc9rSfYqQ8hcSKwgL5aDPii4sxkX
EmE7QL+a4vMRgHb+YX4jPdXFykJpLBPDwdpXglwbbntB0CD31laJ6GbLo03P
U7ppDapNm4JxM0T5hdxWvzoaF2SK6dnab74C45I/t3WaF7l1TToujgmqMldX
NNu+HpJXW8V4P+Hi3L1jQvt0fmmc21B2BUIckJWiSLAbOG/YMISWgZEIv2GL
EZI7zN1Wfvh8X+r1aKBts25T6pRH6Gx/kQFHPmEfb78CCUrwlXQaOpHQj4rG
a6YQJ/MGOuQcI0Zrf9GPtKIKQoUtqtLq3YBm/PYWWUmqdcOjjyBMCJ5Wy+e2
NvfWmm+yUcxPmDgJJ2rLre0/ttebbNHjy7ffa+vcMeXK1NHvw6l2fBhoxr2R
8YDLF0GUOq7UYNc9Jib+m4b/KaCKn9I/2KCyZBLNwTG3FuQhi2IQjDYNc5j5
e/7swtCNV2YvNOe90EeBgQL16P3c7Eh3fJIQO/pZNVibadp5m+rVuv5ztu7v
aUpFWhoV4Ise2flolaig9IaPTRzuzeXGUoJv3WXhHy+nLUUCQvlqqOzov9kf
xGQnkzoyKio//yGPX0r7hVUpJmp2JuYBO4wC24wI7+lwnCilHA/z1K58mgd9
4PrKMubJndT9ViV7W6MhO1AOTrqoS756sDg2sebpbvX02oyhupGsf3EKE3el
9iCpxXGNdgsygGjWIgzt1zoMiJrmzym8QBi2IRS/t3MsjJCeEPYTdGGOGs6D
QeeoMLibGJ3KPKrMNnMEKrb3SXG+8MxctHq0FtYbKZSKGK1UlxyxZVh62ZZM
LdwQdf6jgXQ7cADkCJBkTHttHa4nVn+ObzkYG4d9EaSQKHtfqfPbeDSEIyiV
fGLyB4EH1Fu3B0qti0L+gvlCp5uUbQu714svPUY1Y24kYKzaKhN33AcibKST
fHN1RnrqoQDhjgaI6gw7k+N6LcL8uGGd9X9k5e0F6BkMGYpFVcslqf+1QwIA
XW7ARCjViA2acczJizmx1UQZcjCgPTeiH82qNAVZCZ3CNW1ogbQ4OiSWLbCr
+6uUZNn/7H1wcoxnVhNzZbK4GOqXO/6iKkzF44JqZTCD5Kjq7CYhw0c01ogP
1xdEl/kpLFC4tRt8dIyeoURPAqXUh53U4hqcg6lGK7yUJmO3oZ0Pphum38P4
ujOMKrh7pj8WPKW2jRIHncTh+7+9cw1hT7J9lZFkC4KNjxe2Qb7BJD79AB4k
4O1K3eMvcV4SZ1EHxN063ZbJW35Fw+wngaXQvfG4jRBKD4cazJsRMTK2+Yzt
QcezbLR+N3tfMdrZWYUdbrKobmkvRM2U5KNloTnzJn6EKmNxq1fXSuxh2FVU
bnDRp03fmENxLE/MHZGbZ4manaxFJPR73VexOArnbAZT2+yJmCswSGj23lCV
H408jhONdXvfGd02FNLrGVoD8Um7il9QGJrzHeF7g6hWr4NELdHFQ8rj3ar3
UU7yIA4yAj2C4Ebyy3hwvlFMbFN5pC48z4pWr9Bgxkcu/d8AQMsGOha31MCL
1HVMV5VXpr9TrpaElf/4u3DOXeXIA6eK4qggC20n0YwsIhWOYqTqjmOwjroB
ua7Uhkn7d+Pbp+AfqV6zSLl8qZC6qcTLIT/T939o3mC95PUG6WZoBzGXDx4z
xEwGXEartUCXVQkEFsqg0cxqRlvcfs4Qj7zv2bUIY57goLpFWBmXICGTICd6
FPei76vleGVIlPam+kusMjlAYOAjKA9sxxQZS+YC0xf9QbboPx/orpt+F50Z
J3WOsjJfZ74XvcdCFuMTy+si5573An64KV+ic7PXgFe1l0ylXDxF1KKGiR54
Q3mxfsz20OymUHPP71YTvwlcBUOxyqb9JSb3KmhzXKmyJhZ0eeVt26HiX4Oa
+N6zrQz/nQ1XZ84aso/IIViYsUmogvRxDKTNLJFIoh2oh+51vgIk+hFTnvv8
vE6hRPYLOHPI5aI9fXhqF2M0K3jMT2vvx5wpD2ySE2yZDOCfXQspTF/LsKV9
GPQ7cGkRWygYpHPvSJGpQCpBVxHpei7dzFOcuCiZg3u/v7+oxfAEa5YSifjT
9P4PAbbcuyaLOjEMSjVU92ZdtG9HT/Gsp1TDpJU7hkcgrPkYr+JeCKSa2hw2
2xyAFZnJLn6zodKwujJmexllZHDtJV1e21o+h87yZRV8Az90TTjgke1muUU2
EbHTInNiJk9imKGKq8QS5jOfzLCxeAKbgVDZgcKBsT0j1Hry7xj2rntJTxRP
2lYBPcJLHfO55jQDRemhjpx8ICN00uCgRyiEnypWLCHUGiZoye/pYKLYlr04
e66BaEn5r/RQGXS3K+ffIjj3jYuddBHI8pJsmCYcH4Zvv/5Q5LSRKkQxQOt+
0oXK+byaGg8hX0JNEZF4pCl81Z69yNQCAzoAh5prr8TE3fEdf+SVn0PjL/ru
rtoAHlKfIM78NdggVBheVK0kRmkxMhPeyVtX3OqE6exYHunNFZKx0GLjY4PQ
fKeleQQqeJmfygRSAoU2ynWqTlJf0MtT7fi1NgXNNng9q7mc5BDSK5T4cEkh
YN/bB5zKBnCzgozVPjEV5x1xqCbe0bxlzY1QWkWO74YcXHTdVnmaQM99SSEj
V/gf02l8xsLwsmmuEstViSJO5CCPgrOTef4YQhKvZCiJ3iWhHYHdKyXT5bBq
9vKN9UYAJu0KQSt8FJNjG1Ak9J0U5JO93jVGa6wja+JMkFKfqXMNzghExomL
RpgPCQQ+ZZUPdJYXCZpryu+2FMN3HSgApBqT4SKedNZCh5LK3b0yn4B9Lik2
kNHtSa2TqVL/K1uaOl6l9eh/PgqKHZ67SbJ1ddU+bvKPYDq5wg7A0M6Vake5
91kYQnzSoYoIEzSu8utVx0PROlEvqnxq0rtjnVPIyuGQNLel2wDFV62sY5IA
gJQn2lfYmaavKBApxxak2OW44k4oiwqzzNVw3qrJP56ad7NFpOOKy1ArOi0Q
VHfc5lZvz8qGe/9azx+nmWcsNztPFvpn3fSF4W64GiIhcb3Ie+nsxidB4LOz
kPKxVkKFtCgBIC4kQqPinPcsmgJufRXvcdEtBMvX+SwqWqr08FMpzybdTW6/
xkFqynugsSYDwp/iRUB04MTeExo7bGbM45fxn03GZiZUH9ongQRS2XIHZObV
MR4Q+tjyDa/WQhN2tRS3WHUVsxSi2ZF9CHp69qTDyVl0mbwqxibWgbklI5Rd
EbrUOaL8iqdRB1J5yK7VqGvUZioD2IXha5BdtgDpxl1Pkyc318WNRQrtIqEW
OeYsn/uAmkZoD4xt4FEzLD+ysm8FbpDEKpontm3xH9ETdv6UHwpNK7HT3oFl
hGun1WDCeIrDvWzAxVNfoxGjk5yEFz+pU3U0Qk0vWxQAQ2ZXfcXXwO0YsdX8
I0RtXM+pCY/st0M4zNTbAgMQOTrEzcm0yuDbU7kvo+keU8XXiUi8aWSG4Oc4
+q93EcL7nAYOGZaLx15iF3thxfZggeBUZ/M6PxkZz4Zl5i1ecZNPYt173YM5
5zEOgaFR+pBj93am281cwawEPHEbUsHT23rXEbyyxSnZV8p0FiS2UKakO+Dz
FSWPn5SEtme4CMPq1lxkdN7j2edfZCxVnD0Y+s5DcBHUuRigVSKv20QQ+W3Q
x8poMwVXNfeUzJWz57rTOVzhoueWAAjFYUuy7AJSSPVAvkziJDfz8fmyFSyY
tckoOxCUOaq8wTrEKV9KMdNTgsUSat65rvEeJPyy31/h2752A45qfcS3Yx1Z
JdboNwIuYiFrWcsbnVERhkPE987qnrPJ6yKK8tBXPiImRdPkiAlCPf18ezok
oNZ8dmhd3Ysb/OAA5sT9JNtB93q1fihB3j8SVvMkCKg2EMzuY1zTKiBx+uSP
lrsezPsNxXCYyXZWCUt+ocQvMJ0Q4VOHDxiPmErw0gmkEbpH1SHOunLCEg7/
Wcm0pJp6LZvJau/IRuJSBCH8MOJFyrU0VubS43W0KatcLPAZBe0ZEz0kAM01
lqBbrZQUkskjTPogWn2Zij7+wxX0dY0IRbG7AAQQ8f8H6V5gW26BnkaMoal7
PxuO2SDZN0p6TITjotyIIoOibcfIyvFLW2+yL1dfLiIm3GwTyG/ixsHohh70
6wZMmP4MGYSBMCE6EZHLg8Sk7U3tmuim4Us3v08aFHh0C307xmpS6OXbU7UR
NiIqmanEqWx/aLz82E3UhnNf9SieoiSrs2Js5gdv2Zxo8flGHxEgTXRlq7J2
3NEPlIUouQyUPnNnFxlfzeB15O6d+2zaBS/pkifVvKxy9sD25VL9Lbj5vx8A
mM7eygon0PkpbpiD2t4i52/nzCvjnpwnKskxOH5ihzIWT5mpLKVXJlwN8XHk
IoEUBB23JAxe1geLrGotFnWnPlSVVBpvR0/9XoiZ41zA5+UDSnCxY/vzDz+b
8uXD1T7/TJdJf1SKI1scvNNFpOxI2IDfLoOqRUcA3kue1wtkOURTTKWjbWHF
BXhTK+dgMC/GDPgb10hZ7pFHESn77YaRU8NgLb4ds62yuYZvN9IPWftBg/6L
2dT5rViQSTohUEGVnfIDU/Z51zM3CQ6a2UxwDbMRndDtiXyVSnq8HZsPu4SP
oaeesjAQXavILomPHHC8c9IRU8dw7+8Ngdk0ckftZKG+aDhhetAKMXx/L/ue
+sB01T7NHv3oWTOSxgPup0QlnU6P11pMPyXy6sRWHf6S/BkVmPl0LAxnBi5M
Qum8V5zlZAfEw8xmvuXrLUX/FJlQOYo5u+8WNbsRkQmxrwaMjam80ph9v0Fa
yMbHjJ+sjwT6bNRF0VE6U40Sd/dY753QWx0J3LSTNfmaftO8KoT6hMdPYLqh
Cy4jp6rJu2dPZ+WfDOLFJNzk6WhOc1TCXREsNNoEMFqLHGg+RvIlN+JmMHIY
f4LX9ggutvY7O1q4d2X+9RG1PDpb7d3r2c+dntRMd++IVG1uoIRMZNQX9Cnh
jSPXlKqxHyAHJ8rpWd/1dk1c3DfUz9RuOknnzTIQzjj6iU2v6S6Y/wDtbnPZ
JkSpAEEEEQeeWf7qzkVl5WL+u/kdhgQSAo3gmWy/PDskbe3FbSPWzvuZCbxG
INxQu1J77u1BT2Ca952vB4Rbbl1kCusbmpSCcg2Ok08InHVbANhJZIbSlDi1
rIc5jdH9Rz4piS0EGh0Htf8p9CAUOReaaxKBFGMz1Fz9NS2LM9wxjJcEvtAA
W2vt+fVDcZSqKgnOAY5+EnP0zTULw+Oomxz9nRyl30BPbGViqdUjj4dggbFe
2SkrZX5zlPh1fsKZefgmtxsnVYuRuveWTK8nIOrAgk0p03S1qNCENNhXDF2h
HRX9fZh+ULtFNTgtW+AeX2JjXVyOK+Fp0qGoHQLYL5gxx9bAvNfOS5i4nEnP
G4RphxWl/M9EqiwAm98KC0LWCdQlBEkEdBQp+wUgovQ2iGGZwpvTidIX8nz/
Wi5J4dq0ChcnPB1yr0zh2of7N0Pg2jpv2OaAaM8t4hwa8+gHklzgaDwcBVXs
1m7StgQJ97jVNlpQKpMai66fANL7M0JTeNO6BXBN06fE0N23M2EMs/OmRG1f
ugYR0godwG78rqDmMRbcLNa6Sc7Vpvpm/xy4SIqarlM/qJll/wi4raFf5TR7
F3U/Hj/RQ9BJnbskIYG534IVJlR3HNiSchfkCBfWj1cUHWkyDDvGK+Os3Tad
RiFiPpkGjKzCCnjvuJsIurpdgTysNJGRMulYj6UeBxuDy2pMgmKCs8KgS+RD
Dq9M8QZ4unRht1zLjCaHmQ7ZP8qGKTHj3B76ReuLpNCA3BAtghLUGCY5ZcZm
d6b57f1uarltA6nQipjLkkeS4mDC8Rc4h+QzTQ1EIGha08ZPcvVxGE0S6iYJ
lArEsIzXvg9tFcGPVgmwBYmIB9Qyd3V7bG82nAxzEr6330CyH/Vp0uJWC6fe
rvxRSalN5tCFd1HhDD1iU9zTjnENCziNsxjrWAcQNfCk+xffB1MQZI8+XUAn
Fwv3IYWwuaJHp6zwxWwKZ1Bl7M5eSjSsCoiAoT2ecFKYavmnypZrscsrZnHG
phokXppa7nnYSmSvUL00cmMcmHtOqtlXJOjZV9/gcv8KKn0AB397qRggpgqz
szwP4giak6wCbrPWmNmbEOcIFLqEt0U+q/pam1U+lzEwOgwVXRSmxxja4D1L
EjLkH8wXOgiSHX+CPeG+vP+hE/D+u83U4HpI/qHfW5ylP3JYPVj/5xLfKu45
K6UV16l/8rWiBQlIuWmKHMFIjJ9mQnqqfpV0BAXNur16Pp61BYyAQhIolyT1
vDKUVdw0JD7lXx6rB+tYjSUwLxdrc7BWiBjG0MzAXdZJK2qS6FeTDV8QQhhw
pCWxcKLc4rsT/TXfAld8pGyozYhcKHJo41EbaBKS8Yej82HtiijasnysO/Ie
JwDotGiwgqwAwA8wbtS/idVC3Da8qdrEONzC6xw7paZ9ka5hVgsaBIEJ5KIA
B3jjQAkw44yI7oB6UTDeQIaEeg9bd9GblayHi9n6XIYBm52nXWiMmbC6Dd8Z
TpaEPR80M5nP2UO9LlVU9rW4fFxhhPfgqCJ+ObnFrQozwapAKQ+wZxuJLDLs
RC3prAvv+lpKxPKdhd0uZVOxk6NG7onJAJxA97y3LEyiOzOLgPSya8zvHhrb
Ur7BY6+NQAQMLx0Myx0UQAWHiJ0FPvinutC27JUh4jvLWLX3F7NTF081eX48
+34hFQbd+fzTsEXh5IyJQo/wDwY/n9qlPYRxwSzt8HxwYdIs+lPaUv+t99Vb
sKikS1xFeAdnHHd+7gSoX0/2JD1I3VFtcZ8DIMotyS9CKyJWelqr6i/iMYK4
L69TKvpvHyZCwmDmBGC1PeYhDP8Nz3qcRQVRTFWwuQB+BcNqmRwbYLHkPJN9
Ui+MspNpDrHRXkNHMGnpP0aa+LfuD//GhndSRETG0a2bDCLE0WLkyOn7ZdMK
abq9S1qITzwCW8ZeYZfVp0Sonr03ql9Sl1rxAJ2Oghu8WzXJ3XdQ0mFnaywW
LZJvEcKpQ4K6VhDWEIpSd0j2LAuMRSBHv7jcEke8huDDBr3EBhtJOt1zrtnh
FmcSHgAlgi91sALUxDqvG94iRQyaXnUI2CE58bWIQBPDVanprs2UwMFaK24R
reA/UCS9TBdNwaFehj+pngsH6VveU0fF+MYr2S/cgIdO1gtqnwLqur51qOxF
zfTz6Xwce2olaXi1RbqX4wsHwRyULucZeYHYocX7QMzIC9zDN75pinQe2IUB
uMi2g1UkCIdGwY9Db25b0Qyi7tAYXI9ObwZUqZFdh1AWnjdYwThVI/+ZPNFy
rpbaq4JEyQovBf2YlLaKORJQpof4Nw/ChIjkeyP1+OWpWbVFInkf3gKePIX0
pbEakGgLzalhuAb/3B7iinqbRNkFfGpI2oQS5q+N52im4B9o/uwmByh8BQAp
aswfPjUrZMYVJdBLApQnEQVWvgxDJGE5zRFOhNLWAxdWPTjVTuMmeltR9guR
iI8xCIV1qHLKl8wyENBuGHcvOSqsu3b38E4uKBvB+hpA1KYzFg5sKwnqRyqH
97xTz/flT3n9noYngcXx9xtzHMaD73t+/SrJHxFou2Jz3g/be+NvYmKNJTMd
boUDYdC9sWAPEHn6wQukQzV6CzEiBbe2GTgmbt7kh1YSZ3XqlQxft1NtgRM7
+GJIJ3aemFs6jkMLBi4MASfykY2YZWfRzzAYxOYv0VDxY4v3YbbrRSN2awBW
J7K7C72QyoPzTXixv3EBEtRqTekwkOdxSBvn+uArIByhQzQJqFP6d4KyZa4s
FNipkDCTUWLeNiRkzO+57sme3vBBAx6pcK3ty32kTkY/Y8dBap+H+6jyDTYA
wpl7VTJI3e1NAT26Q+IhnUVwcc2qnn+qLbWPh0eVrWu79FQa2y6huDA36jB6
nR9XGs1Y1vnUZWt0h2/bFw4RGPjTVpNKsDP57eYJnM9qlFANYMapJHsH2Cpw
aKOjezbBid1UWcAQB7q2Bqvou7MiDC4he/jSL7mt32ciD1OSh+8l/FyCC5T6
RSGybvjTTL6yA9i+b0a3mtzMaHOGOCzracGNJM/OqtFNGNYoCfKUG/mqYPPs
hHGLGgcm1UBSFQ6ajCZK1qgB6sJCy+YligzQ6hmLc6z7ALFNrPHricqgg9h1
98fQ0MDFSRtvS33ibSx+pQZor3LydFHE/QsTOqtgavvof1CFl663HlM5HKxN
tMe54K8/VthIWBb9VmFapASout0lSI4ZBfQsNYtYe+UKX/DYTd1p4ipBB/Wg
KGA3QGu+pXKVBq7x6Hqe5/aE3P+CPrahoxl0zv4XyLkvxvAx1bqAoA/xw/KP
irGkarkxI4H657EYHH1K3h7MJPYcbvLfMWqCC89Q+Sr6iPirk30Ex5x7+YAj
m+YA7wdRst75W6WVnfukr33gXgnJ/C9QaEpvfB+KGnxs8riwg5F2xRt1gi9V
Zgv8hf0kCSe5K13w9MDcHQlN2AKAtk5R/LMxlk/6/7nYXaerfTpSIGZz5vyd
gZT+1ULpoLmqXO4HLtwEjKuNy4f+06bg4YGZ10PzITiEsmGxD9iK+/lKMDXD
gT5Erv9AEWUj7Hr3si0gx6gMbWa6uQbAjCjlMKqEDmC0UWtNw7FtxHCsXKif
WK4/JlXVsDECW86//jV5NA/+dn+KOfSK7+zFA9o9TZBFrC8ALQwiT6OWSJm+
GUjS3UiLojeQfdcZMV4vfufYYjxRW+XlelGau7GTcwHOeYdmxlTls0nF9Tda
sPEG7/X0h3mco41Pk9bRlwO0urwiYWCSN92tHXzXiCz17LJqEcI02BQE2DIp
T5IuhnUDqet3JBG6IsrVpWtCf31Ve1Rp7ciUCDnB7sYB17S0q+mVmyqd3VTY
7cevpl6n7z9Nu7ly6/nlFL/ibFN9wjXibAeWWAF5z2MPLRd9i2IZSOIkyvQ5
7Qu2zaVfEfmCsy3e/VBronjVnfSZ7hCaoM+enZNQoYHfdNk3zqg/3z4DSmvD
biiPWTxU0dBmUXbRbHDpfhrJPPU2GUD9tXh8F5vWOr/fcmckcvv9cxW58PQ4
ecXzQCLUDrL5DjkkTiqFNV9bPvIgDnqNsBU/VyiwOgn4nfYdh/AK53hT5sab
3Afdv5sZ7KMu+G4ZP3U3DAp8JSrC+wRcAJuSHzK2WluiHR7OL7in8JXYDJOI
JhOgUapfARpngzFXF79NSRY87ZaZVHZdeSKSSgSjTmiE+3uw4n/QvvG8KK2v
/q56nKnHEWFhpvTwjEU959VK4Lu7qHU5CTVppz+r+TtCngiCoc4lk3zxSzcf
CvLG/qUrWh6x0o6Yx6g38M5SHioUomAgwuKXVOxqV6vvzuga5WVCuwj4lP7S
eoLAs601xokWAg2zqcTQpremzhS+RkXM5cAYHWRfHXkXJtx60E1SOZ273MRL
6o6v6rqrX9l3kgV9uWQacYV3ilL1QKALhRVrQLB8kXn6Ss6M4a2LQd9hUtoV
hbczCVEmO0mJQoiKYX28zEhHTmysIKTeFGLv30UmUXGH7o0fgtyC8QbhdAgy
cOgbvWppmw+e0JO9wKYWmlyJud6gO+7G2Zb8sKSlQleVr5+JLmhlZ6JxrLyi
7BmVfC9D9QVjwfW8VIakxMRVAk8VYku/ZtNmamEGM3oEkXDYu8S1CWAdeK8b
NzhEpyCqZHaVqcZTmdrZwzGI7TC207OA0VlIA8STOPgwI6hVCINKBMX2LNrA
IDqZDFr3Au6N7Qyq1SvnLzC9DJOfCie8Ig6WGMYE9sEM9+h4vWfqfn8ohZM2
5vHOZjkeDQodKP8od/JP9/l2xZQuXe0MUu1NqvIOak2d+52a7fnaQbU2BBWv
OnJ9CLqAvzw6J/R7ISh2QR15Ad8H4qM95HKGvaoSkYUpFehu2jgxHXFsv91P
49q/JeUkmdmm0RE2MmeBJMNHyI3ZLj2Z7VLTxGW9fcfDKt85BvfmToNDskE6
jvfZ6cMxwGde1Km46UZ7lOjTVEg1hzRkLT00rOuU2BJ3lCu9JkbaiKa8pPQ1
K7DIe3xfYgQRh7XEfNMAIfvUwrsHvQjkeliVVCD4WKlkUPyyJX4L4OMC67lP
CGD2+HUW59AKb9CoAVVhZ0OuTQ9DS36BAJUsHskbtPB98F/lfA4WeqyENi7d
qIStnSOB+orC0WXWhTux4smU7XPJoxsKMlsvghGXAFMYvm3me8GsKqmOW0QU
DcapWMv8QHS72bBnXEiwkHyYcqMyGhYKHO+X3JPr916pMas3ykmeM81YJ9cJ
eTRP9vQakSSRduDFHxHbYd5oI9jXRs0rZB1HNI89SfArqiwpV1tBXB3yK5RI
McaUJJXHnxxeRB1koCsf//XCg3WrAQZmHJhgOeD4DA5FcECnWFPRsZVwtq55
FL8slF5qzmqfn/OdYYtQl8/G08nqjW876RkdoqbnlHpp7aDr0hbVbSE9x7Nb
pgWJvXc56c8UqOlri6HECa9xP34d6SKOkIfXn4zhZ6tXj4JCsqZ6G/sS4sTV
qeyJu8DF+64GK6+9y0wtuLUs4VUWGPcM28U8PCea69vwXHVxTiciHD8LenA3
s2uPY15TsebDlr63hdr+hGil65uy0YlTz9AULLLq2VlwkDb25th3U7vVTdNB
nfQfHQib2bplOFmoAEYmBrk1Kmc52yFltYJ1XjePT0nFf0xUNZ9h2rQJN7Pw
gUshYarWgIU+urYqLlGdpFXM5H1gO0uRyLBiR1c4LBJy9I7Si/CmGy/oNxq8
jSa/iM5exYYogPMc4zP9CZDks6vV9cOsPLkOTDdmslrgREYiFqiTzvgkt00D
jvbO+8mPHsJcvbbM+mwLL8HDPqATf3KNxJVgxGaYV+X/YykwxnPr7BNbovN5
cAq9bXmvZqt0r1NrV874pbvUqJx43zLIKZ9H1bCA3GWc6hsv18s+OaU+ZL9A
8bp+E6Ngm/sXaE4Z3tM6NcsFUMxKbh+7c0X43FoS6E/KxYU4xoe4qJviIsSI
+b1rnKFHQT+595UAcEec566bbQJOok1mNmeSuAtRHqhCND8rUm7MHrWuWMZz
3ffEZ6ktXdblveEbAgVrcj+r8/b1AwNDVP8VDGEJnGZZp+9YYQyz0DMgiVnY
uXWtxWKyc6ddGxw1Bu0K6v45iYn6bc8dJaAZWKBvPjy55qZ1RReJffprSwum
lwvJ+XKtyq2HQDUOQ7whMpJ7QLNAfMHEFgNxqqIFYhU7HAIdtC71n4ADru7z
wyCejtXheiC0kVrlYvgJLNFY3mAwlAWGCRaPr7tF3vOM8S69WbbCFPQPBm3Y
epy3/EORO2WNtdEeez+YqD2YGOq2C2aCrrwDZuLuJaMcdMxbevGV5ukff3U8
GQ2axYFC0arlm8giSdsOqZ9gY0GgAgrGFa1PYhCnxBOVxQmjY8MPYm11iDYE
mSSbb+Wh1gRCdYlfII2271SmA6rpyPDi/A5S8rCfwAJFZjAJO1NSgMwDMgZ0
856zErxkhKV2ANlgt7LHVIy7Wths+mWbrFQGJ3saXlJml/rEChODja265Fw1
xtQlwVlqGxh/Bz82IWbL1am7T4fGUd8uRRQE94O+M2EmHMd0LWKV2Hu0vehR
9fRoHrZn5LghNdQr5bRd6fGB6Xh80BGEvSyNQiACces+jOaI5PYfiJQVPSP+
LCDziswU0st1tn1fQBYgbDUyJ72eycF9KKl4lYynXiOSUqZYv6mbz/w7m7Kj
0jkOE4RimZi0umxRsvxc40W/yGcn5hQs1Wej665F+WFBodatONx/ugjO6nCW
WjGwzAMdWhaplcHK8OAX82ECHz6IyJzj/Mv4KljXY3ZaIiVDImwg56W+Bh3G
6uzwDQJjWIjJppz9XzawxI/r/jigUJ+pH9oApLbYBJFTht6baEJo3q4pFcXb
ne6L5nP7o0Z2zelUKvdgfFixbrFuAlKsR2ST9WkwIUklqK9GMepn50Z88Y28
HkxLO0YKawDl0RVW2SI8e6l+6Batoa0A+CcMsr0j3xtrPdIeUIrwRe/c+140
Z4QZ/3RL1JKnSBw89bX8+2ZDH4iveN/OvxEjCT8VWn6HkWSPN2ozoKvi4mOZ
IhCnQRDFVJsG1Mj7iBLjOW2ecWqrzSeVuCCjUUlkdogxFJGJ9OAuwkfEd2DY
wfu6q21poyIDKKMw2vLyfwDlsu7un1D8RNhh8ZAQUFKVSRj2LCqJPWsuIenl
EszCZyzuNHGZ5XFqCOW8pWJJa8BcLT2AhdxYBcGN4kbxGq4I7KEF2pOIXnO8
78GIijMuHz5uo086GJNZ9E5uFR/pAmnJTZVsQyTcuw77sL0ieYczFI0ckjQN
EdI78mVeG4WKoAzDdH8J5jC7+eG+dvnYi4M3mp9+a7ObGjeutDYjG2Pwtw/S
Asbb//xvL0viQUA+BWUwU5yi5EhPJTR1BvvY/0x513ptWWZL9hXblOzbufiW
dcM6rODMHJK/ExCBk0c4EqyQB74/bzLC7IJM2dja062wHJUmHYJiRQ5TuK8V
LFP+/E3+LibgvItKtREbCCMyAFum+BzWkm/0gqmoODXKl7IlCwhu/3iTe29F
TtXaQsxbuwCvhlQrz32fVwRO+q1YfkgbyFujfQ0/cu0iJagQCa2OV23+5aUc
CRRKX1AgV5lJEfqKx0SYID0imDwPNbnrihPP7jrN7AK6/StSZX3kSJaauTT5
R1pyvhwBoWfdG2WE8SEVljCYgSKWaSdUwwtG3RxVSxhDS63zSF64mqu2TOs1
yfZd2KtpBpoesGeuBe+Z9mUWQoy8YsFS0ugBFe+SxaSzFml2ZA+NqsM8jyfY
RRWnBi0EHT+chvJwxqu9dLuhKOteFJZGK5Yb9AFbxX0rELNi5Da2gUJgTwXR
3ku9iBws8DQwQhVpZAy+cSBwCZ0/zUd7bRN2jMM3ojqdaNaZglmrtSAml4lP
Zzpn5i0OdrTe62wR/wOLi9cC4hgTETDe2+TDp5ZmJbErkParxQGHoDy9DpI6
3YozlWOeumd3iqb+J9toq0X4L5Vg5sRAIIZYADNppxPpZ+AmIY72rQgn/nj4
W9G3g/Xl9QJAFRgc5nfigxLLKHfKmxBMYM6U6X3bo7FgMH6sxeB259v1TXay
iMIlZsMLOwbLyxxgU/MR8Tww1BnuZG1ee1629qCR0tGpo0GEPzLomyPcoTwU
dWJoUlFjL/z66/kbZEqYaWZyBtYUkI4kB+qHVVCOzgI9nQDZ2Cz4UTuORORc
3GZKFLNOoerFfgSZv06fg5oXGude4Oc73Sid50dLmBAtw/gVWTpQTFzvnXFr
E60gtavXaOI6dZhIAkavc/zK5e3QoEwbYJY8xER/pdwHLJNVSdO9+uPvzF3o
MNZ+JLVgRTs8sHD0UPQMzv8eXRVjeQGrmMf+wHNUIRN8RlEHu1hkJb/i1IKa
xlO5D9zPplzLXCuLs6c+ZZ7ebIWRPJkcgBB5qU/OIvvyTuLmBbGw1t2HzhCR
y86YyxHI71ww4kRmL3lDjgbPoK0mLxyLtZncujVx5yy4NnfDNzg6lFTQtp9Y
PHpm0LgBOBxqbViftlgkMcg1HEHp0rGJhQMJQKehKLbU8opduMvkw9izeLWQ
c5X1kuPRphmLxHF80VG7s6obUvZpNYvYmDkouol1Dq9hvjyA8rTAfT/vcDzY
hJUEKFieGUsXf5gAX2YQRwHc3HbPZRgWNMfrEGNTBRiHzceRkTDqqS6zcvGb
5NJBtxHxYQonBy+5QO8fVemud17swTjYqUKDftRyw/vEuFCXhgCfC1hRcavU
VKYp0GKHnw72O6qnPdgmMN/5DJpUxrijFvLIpBlRjMQy4Eb9tdof6REskYyT
81tPSlZ5dz1megmQNFjU4ZJ2iA3Gx+/PvS/4xsKLXy2/e6KLBjVT4YdSZ17y
R2Lq3f2wGbDC3n/TEb4l9OAgzqgi7JPYtnPVp1gawZNodkr0FDPV3k0pfVYl
ZMjacYv/jMpP2hbOe6ThRKHOUS+GATgWtGZmww9m36h456ylQO+1Y8+xqYFY
+FjHBtAKzAkZvehfUn0fLPxTrPB4s07G/XP6O0X9FrLCg7zyrUTQoKuJjStV
CP6uXnQvJB2Hu/PlcCEBUIRQgkCjaFeOmqNVmH1AjYkNiPyCzHg7OuhHHrze
OP5BL+a4eZ4CzMEhulG2iAbGVOdxMdBHFxHMCpDbACWJGPsuPskCreXaHvq6
gYYrc/Kd78MI8vGGqGY0Zx/nofKLCZhVcRs7mdSU53andd3KvaBJUOCsPPPa
Lfd+u9A5uqQS60tSHCR+88Tt70keA/7J9pUb1zjIg35ioN0ntVAvVWXaB/C2
TGD81mOAeILwHKeUOIzPfpSPu+S1/xEtbqOJwmhjlEQLFD9Z5nQVCGjP1Me/
tlbyG16Vy3vU22gIq+SoZi3YV9h/UN5mx8EUHyO/r3yvgvUH0OERNSQzgzP7
Ivnvw188yNW60wxnMnAOoGDc9sMt8gBcWtd3uq+ENw2zmZlY+dYa6ykCPd6e
WC3Tp+IHYYlj/JHK86hTH32+WsIf/X5tj9NDuo/jItOZ6TikickdXO5j9GYp
dyQSC8jkRNp0vLli8ciV7YrYGYZAxOK22VHpXP3YKv8F3Cm6QYazokblq4X/
4757nJYXVbg0OVzkZmniN+PbSlknLz0CB8bQZNedZHkb4jhTQVOt0R8rKYIg
ZtyA/JQRBhG1S+6ui5kLcwYTtwzxhpKAARMHlmwUiYHc95Bvxs0qveo7LaI8
Wvt5WITy0K/qK3gU6L0mjJ/CIuC5FXKP7NBIDneesGkEWk8gpFygQRUafb92
S3sVMZ7U0LdxZWWXnuWzXQGUg3iikjucMiJ0kSL0MGTdSxgJTqbhuoEv10LW
/d+kKDSp4xiSwGNbbNYVnbqb1dGLn72PdhoCOVe0iDDJW9dVKN07oub8X2wQ
4D5RspDUK3fBKSt3pfJ6ZoVBsdjyMfT8tcTrWj1+/ZG00p7yx6pRrR0n5Kv0
DlwDmsO9VY3ogYVbZXYWR7SZDeUZckpC9X+xGq08TEafLRRsq1LF6mR1hblt
IG3vyRh6kR4kTDJG/IimYvpZA3zFvgQdx5GnezX8d8q12r/Zh98XisSHslgK
YNS5I1KbgEUrtgAAKHdbNXd9W8jKBN/X2zFTUsVVGWEOtxXJFAPAYxIOARIK
pBc+vj1C2u1OszReFQLo9HnK/Aei/tnPJV3cfOJLWX7TFlcIEAIU8VxZdl46
B/l0QOBOzOyAdg3v2tMzgV8NqNr3/9Tpa1iJpZy8LBHnw37I1TQmuEZP8r8i
fa3CpKzumZP+v05ndhMgTmk+MmTZl20F7F8eZQmowVSAabIj4VCJuux3sbCN
ynnW3Z0OeDGB0G4rwGZ1jYJSA1SYpQ4VtzQQpiF1aTWXLS4vX3zyH7/2GuvQ
QJFTRgKStxC0uSrBXFu12JoCoHfb+tdVcyqdbkOQW8XBvpF64k7U/gqMllwH
mihkbcGxXuyE2dsewDI6ih4OlKzG6SMPRM0Q5c5ofHvQmImhzlIKsS+tbyPc
fPDydlJdZ7rRyi7D0cSYCjld6kJRkeEhkdT0zhTaqWNJwIpI8LaQTx2CfS7e
fjX6JX6ggliPVGTldRGVhgpJM9Ai7AsFiJ1/59AWcffN2R/agdClBAIaqHTA
mGIFx1bjlw1jH7O86Lgkc3Rx2s6cTlnH4XEtdCjr7evfebnbiOX9n1Dr/Y6e
y8E+VZiiW286QF2t1Nxb00rngg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+ErRjVjRl8Z6Y1Cn4Sa3j4W7m/WvvQqPULvZoXpr4K7hT6u9Nuol4pfX3KyMC+yLjopc5EXlbL2sXFvvlFyxoo3tF8dWPBbh/2SSJt/RGU7N5SB0lJVyOYHvPIRCdKbnoBJxgMcNF1/sADKv0HneYiv73iO82RVvSQo1FMqD/iO7jrT903cySfYNe27ge8qiVYmECEVpzw2LY7wgXAXcM4FCaYp5Yin5HjiRBX3XXLrEgqI/sdJLo84PGpGN8c1M5a3bTyaWxeSkxllKZWjQsZ98H+gyQUyG/BiPyHPbB8ZVh6aCEbAjq8XnmivFbGI2hqYodXwH00ZKwlRb2xDfxvNorxPK3zIzeVD0E6QaTpKE2ySOnzNhu6BMSq2dLWjzF1JQX24e4Ulct52e6VZj8UREpc2L/kY4GhcnbODaNULgc05f7qvRoEC5T+SqsQEnzyFtacrrJx0hjdq0eyR9w8IY4F2BpGlhM1Wc0DkqeUvZRKlu091/Poqa/TXIVUA97tKMSRaXnKD8dmOFf5dKuGGELM54nj3GRAVc2DGtVLj7N+Pg22qoZ/acIolbaiHfnsYtQ6ooFLFwiYM8lenySfQkyhhWhEGpDUpeU3IwbxSkuVtMs0tLv2Htnx/iYRDDR1mHrXv6sF4JhfXQFVnTpsWQkRWEzmO/X21VvO7MAqTvZABzg2rf7jOw5pCjpLmU03YT6NERWgoQEFIwKzIgz8kmb+uuv2L1bcUH/uMQVOOfhA6TEOKkJYeCY1klcHzJAUbiOtJ7GcCG7W5cFPgKuYNo"
`endif