// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KzkplKPTcYWkPU8wI678JU0Y8Tlty0qIfgVGCG40Be2eyHKMNziUF4lUmgFf
rZ54DF+wlVNto6g3A0sC++MOXi8rikbREAQJQ7cjTaSSXkXGB23DifjFO0dz
ZwgkSm5Dng9YFspMtijjC6n0x/cFHRIvtOXEjj8kIey/OkEYLHlCwfPd0Q7g
qJaZ/oM90ssbPJuyBdqZqVf7gST6+hWyLp8yXqFd30WBnz9hE+akJodh8XvG
Jlt2aDgQEPn7ZyRpsM5iG2nDfJLQXzJtwcckj//9H3nJoLiz4whHtaEWeVOW
gIb17XNZ7Qstl9R6PJCFGa0OOwcDQnl+0jzmYVVTIw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WcpTb9qr0+uZgkw5IxGJWLfkPyGn4iznhV5FefjDCV38H+mwkPQQb26cAsbs
fZ6t7x2cy0MWYffDB9v7iCviHApwE2M8NZZY0qxAQf+V4wE7Gygw4qDVzF1z
TihUkz/c2CPUG8ZlRFJ0aFfZjYOea6Rf1zhS1KX3ngQb4GuH2ox92d1BgahP
7On9eeEu1U2d1+fU7LEnp87AMH2M5zLhQHMJyY25kW9gjRxW+XSYtJs+nIhS
Mah0rsZQ8j7xar1uz3NZq7IN/RNNNknGGTgBvcg//RguxCAQhmvvWVDmmNK6
zqoTGHxOebeVGgXKMEPVY5qoKZSsChGLv2o88iVJ+Q==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pMpG+sv4X4df3RPx8Cj5WF6a//PQCPG122RCiX95ICzyJDKbWfduyZLwczlu
Fk+RY1pQBq6I3gpTCK8r0x5bovLmAkdRTxrwxuTHDAdMKH0YaRyNPXD7HiC2
tVAaZGnWBBu5muQahMKNilvxErJxo3mkNanovZH+YB9Gzndp6XmUgoNonrmb
AjYaKQknC0gBbaAXzzvjWXAxL+T75pp2KSwscHK7Kzeea82BgcMQaME9ajtc
ew2LvnIIx7uEwFnQLCiaXKUPk6GTx/HOKPFUSBAMpvidxihODiGQ3tXSG+3h
Zkigc0KtAnozh8r8/gWqdg72NJu02hIm2fci/oK/zA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IMAJkKIOkK0skL0Sxrg+IEOn0TU9p3OpSj2/anoZxMn8sle174nYpZf0DnNu
HUdfkXXDAOvECTsSD1TZYlLkIPPIsesvbyZqCTYnAHeew8VO4K9Iiws4XXV3
IWjOiNhf867Fj/c7U+meZyFmi5HnomnCmoFXOV+VgM0Mtc37ltH6cHIcWccH
veQ1xsvELaieqjQOuw6mbJUHh8VL2BWv7N2blmUnA1oOE5GItddDA39HN08v
uYb0TFf6x9ulRMKUJg3Hrq18joYf0lQplqJAVB9cjwBLPBYQK74XNjZu31f8
9gIxxAt91uj4cOXBR8qk4W9rgPhucxJ+ryAqcketqw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KNxBDfP3zPMsBDyUozxxqx3+Ui9oGTmDoZmILhyUVHmVfuaqZ2SurPII16b9
KSCgmDF+YKq9e5CdKRrMQSC6cu+Fg8D4Qkm9T5sIX1L2A1sviMIsHTmLRiDT
74tlKPrIZ9yC6xkNkP6yvkNJcIgYVuAz55Ce5l2Xt0sLCdsjA5Q=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
uRIfUMjUnFiOtyMBQrqvp88THrQeE0q3sfjjfWW16WqZ2Mzhxd6hSvJWFZkK
UNxpQUlDK6BJ8tc0fOaxdotZrkXruPFxUdGIs19mJ0DnpYYytZgNrNJdPN9q
XLvdRDGWMpZBRi2mCAO6TwONQb64xxkatXWGHjDnUczbQBqkeXqDz/UzOeWI
tcNjgqtmpXaX7IRh/3r7c1kOlrMMVVyv/NDHYtHO1dzq6gtH/LwVr3spN1ee
j2xqNt3sv7tQCkDGTXkFqFG0grG3hJkxB2ZAMAjGx3PfYzoivKEeEH46sCQy
9d0oqA24cQC/IExgR4pXk34c+xDrT5HrY2/YJ/SPIW0wU3y0tRs7dM+1WdTE
VWsj7JLG9q88nL8c3gI7xdiZhsWvjPo1bIhK0ZzV1K8HsLxeeN7XuofFFxYJ
EbMHGZRQ7IcOjk9C+N6SusllQhXZoIUxNxVVCFJCJQm/J4YwtkdlQv/8BSra
r4d7TCwEJMS2kmg0QaGMiu/9DkKt3CeZ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
AQOrHEzQ6kO0Rx4rusagWy4rMz9ULjYsHtGVmEwRfMzSq1USsWfq14gyj/ke
KLxO//3ox/W5LTwUTHMS7jBcH1tYwWVcyd4lza5TuMa/EAgqj0qDW0fQ/MKI
oqDFHAPKBaztRPobUB/gU7rYkU1uAw157UzDPC72kN3xyW7CiI0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
g5Gu85XMp1aDeXrUCyms4GLN2eQDr8W36FM3m3soIchdeUQmOsWvLluvr/Bk
zq2pJD7RcHiyAjbhw/HcxK6Yp/Wejc+RqMrVf+9pIH3WaubCljT2XWvxKHJV
/VbOs+zR7M7OwSEevGtAvG43Ygc1UOGSXTzkUWOkp83O7GjPAMM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1312)
`pragma protect data_block
CouPB20S98izioE96HcMmHXj6QFtPW/Pbm9YZAXt/VH+8FhYmIidIz3Naj1y
ZCt0oJ2U+Bjk+tN8EhyB69TTefT1A9LoUymf7FDApf2D+s1z1X2wH0u3DWMA
mo+rqTOweR8r5r4Y5ZhNNdgRWYRvhNlMPPomDPIPjP5RTN1c0yn90jSTlVaZ
sAok+HVQ0mqhHjTgs9LsfQtvrkcTqmMp7STcyYfsr0IFMkfzlqhXrehGJhLz
sq7/dSygSGBH9PV4HDpOjA1+gjTsWb5SQGQ1E9fhM2rUZ7zzXkdSWo52YKHa
xHH1Mmj5QJRD1QvHtB1HJNL6vLBUA9bNSHMzPZXYn1VAX7S1EOBw91aQf2X7
dOR4iRSHiMLEFlf+9/0znfF8NQgcAHDWEg1Mo4So7AordXX8x/i1Z8n9bOul
+sxznvBP2AL2wpqUE8ync4/0kCCJRfRspEVvFVPrKKTklmslYrIL4g2dNzc8
URUTAmm45eiac6zjbD5fq6b1rp46y6y8M/Gg1L9CpT2ooiRQUja6g8qp+o0T
7fjtAmKHL98Igz7tkefQf/ypA4PmrpdK0OxeXmbuwj3x9S3wM75dgeMW8pFt
BOyEq8TeezaU24bajj5UF79v7vpPM4Vu8dAFE+AG1I2LJReWmaJmsrflbCR2
cyRagMvymu625VCjTC7rGhOAXk2wygErdFPDyw4H/pj79Xl3qTPa/9nxbG1e
XedaQ6dD02t6AGa0KYVaUW5YaNIZxqmkjBc5Apu07hehvutjtf8g1ARLv1Vs
ka0i7tR6VE4JrlvLgK7r7Aai+FNoPuwDgE73PIJnYAeGaAcf5HYgl+CUq4yV
BY9xEj9gaHm8DQDoW2uy4p4j/qIeSG/bYkNehocRZJ9JuBrVaT5kVKfziESG
VZskBkWF/O978k/F2M+59KAxiB3ZhmPyWmti6U8n8XmXaAlPY+awzam8LHK7
DC3bAG0EMSw1Mm7CYs5ftGg0ek6luMYoci1xkJddc5Q9OTM6ntvJCy6oeLUW
RmoFxkNk52I3DUkiHAsda2PA5o4cMSqHgq7bXvMZ8XLaiVo9D6vugIMVIjBe
LSyl4ldSRqGkLe6wdq+aMQn4PIsKfYpU+NW/ljDPOx2b4Vsxyav83u6YjT9K
RpSiJdPQgKlMjwFIQwrZTMclPhD6pCfokxCYxT//CBmr39OlkBhWzIu6/ztC
qTZidllwf7ZonvajiEW1pY56FxyeRoqT5cmfyPLy/uusJq0RFB49rM+D2wWn
ZX3DPW3gWJVDuYCJ28fMMWLZIP/P7dHh411nCzdIzns7eFE7uCUPQjJOvm0c
8CTV0Y/Eq6IRRmi/SKtJpVc1MqobDRULB2bMNUf4vFtr+X9mt5ApiWnoX5SI
0CBsgUMWjqvPmXn4bKQaa/e8/9Lv6RrS1FGsv4ZK69RUb+5N6E96m7zMqJL1
XjxevputEsOyYogtAu/U2n+oX25I1JurVSQQk50rk7kD+NypUsg8NiEut6Ri
V3Xzn8KyMdj5A5mns0jIugrklMlquSzu+dZCu0afhs4ezKiY82gAxPZvOpCv
QHnk5IsOlBa7vec9HZYs4C5KFH0GEMsqBG9EZ0QNvn9cpKZUf3ytIDgnW7qM
cygo8N8ZwxT6yBWeZJmL4TP8CPRRZuCmxj2goKBoSSXgT4NAQPbniPy+KIeD
KgKolP73VJKZ9dbDUiqG1j6t8KedCofxbYAVvJbBoFWx+8j0bALBkTN0c9Z4
ZeXSeNSKMQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqft22P+pL7EEyVeAAoiiKgNXEhckrDRqD43fMk4xWLdUVk3+wAJqR8cANwdKQWqs/t+2VwLjvN5lmg3xoJteXxoqKkFG8CYD5zTp+JovXsu8m0Ou/XIWUTSHDHUwiDszb39vLwpzBC3A92hZt7P7g9wGj9nRidHaSIp3On/RLzhKRgRfVFkYdEN7FcrUpDV+o/9lSIXvnW3F7VpyTyOMyD1+HDkJNOHfmjVtHNo5THmKJBinMaZka2gqgrnCPqJ/TFLlwhCcYQUDQP39O5Xzig4Zf92oEumD8K1AHiOKzQe6+X741cj2J/dEWEBS0cuzmtq7+CJlUCcldeDZsWX2nJ+fV6vJluAX8Z/oQlxlFqwXPCx7mbwNRFVNn0kv4gw9tWFohDaz5rBF+yvBvHLX+D0s8DMRHoOQSh8fjTiY7vYJqMakpBMYTH2HgfYtjVMsnjsMvvORGTGtGQUE8otJXXmm5M7abyxNYoBRzVEMCh5G+9vj90e530OzCtTXTfx5tNIyLwUOf6MYvlljYSWmcQOkigoeNN4CI8AtIVAAV6geAhQ/uHobWPgvb9ov+FN9a35pog07mwoIkXqjtJnfIZwCjE1mmnJOEAgxw+QZ/oFG0+XKFXQFSQRZmWR2tavCaQnnwTyWbBGFaSlUXeyeuqpHXzXKv1VXla5YfmLi3czS2G8sVzoDo96aSdB8AYn/gf7dQTKwEpYrTJSaEzkWXs/8y+Jis3HgcgkA8ic8mU02s3QNgTaiHjiwBsc3JeiozIHK2REcaGG/uBOwCPAWt1Y"
`endif