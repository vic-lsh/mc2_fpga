// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lGGaaZWdA/RrMIMii8Nv4UiMvBYZBWGLILFbIswcoDnSn7xY5vEIdQZXV9Ce
9SY6qappFbKXagQ7Ac+VRe9lVV2NDIRacZmCytFLvFtV2ZRlZmFiSXPy7RxF
wKiHVP+dWCqkCZzUX/xxcdQyKKVxAieBM5MIGrn3nmSgrOOB4rRo+lRgoRN3
fxBspSyxtzpBSy7AEt6PehfWxIqFAKId2c/O8Y1075KX4/bgwBjcohN2RUKW
DS+qG1pHxHzSQJOD2g64PIlyiccBXMPU9q47sBp/L+GQTINV+/99VjVHaTiA
UKLfwvwsOm0qOucs37lopHB1PHNARrylcHx2VHWNmg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PPcFf2wKqitP5R6lyDVNDaNN2IlZ9Q0vuSiSTvdNUe6lEoB6P9Rk2YH5eAbI
8ITIKL+nL+NX51BYRNgoQjCP7pAm6hc52dqeYtfiQ1jbj+bdd4JN81k1Dfls
tGA98yGPpw1I7YCqQOzBJ/IG7b0ePR48cNu+c9jkMh9aK7WFUP5vEJQHiJYh
7tnxtnR/YvGz6nWOcibk1uGZnWHll4TugL2cNOb9smvSNdl1Le/OEisQ1yKB
J08OMYYuugPMeFEyAoCkOlJfVL0tUMLR7/8AniA5bqtyBQ4Duk+s067IpQF4
RKrsF3pvz1rbOojcugeK8WxrBPC3mYZ+Iyoev31Yfg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jKjJowAeQEIkK/EMU+7LmuXc5/+JuE+mYoSHA/CfWmo+aOl8VbnPECn9g1L1
UHUdx57BBAQX163KxKwQIk9Xgc/tuDsT8aB7m67O4zH3xteqadfbFrqxQ4Qw
arQ1P1KI8QAgchGMKs+M3FPXAAtQsl80BxbeRunclcOUw1YVVxO8i+vcozc/
PM6Pl3vSBUjdFqGZktwhEfloRBldryCo6Ccu9dvYSR9uve7dlxmZRDS2xW8f
iLB5+NMsb1pFWvZZFBUObDe0PdnFf15Tj2gBSQ/oCXeNUYl0FCDqped9arvM
lCpfw3+wgDIUjEE0h/StliPoSG8EedPUsJwEmrr+Bg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TCh7Te5p9ODi2SNq5F6El9X/4m1/Fn4jEjoqo/NSvFl0QtFGHLnUbs4UzU3z
fxec6YS3XE+dK1g+MAH6oSXye6cN5ksn5rMjInksAESbkfEpQBbprYbUZI+4
dU0wdrJOY9Kr6YofxnMOUTUaoSd/XBNf9Kgh2In5t2Lm7H5WOr8YKFj5zsKg
vp+X5FtyfneYsLIpr1//sYX6GL+wPFZC7sRwaGLD/dafFJJoHB2Wvxvnav7b
EWf430DtcoyaLO3GbBKSUCK+5/BzpPjFw9ykRWBuYCss4i6ykHp3cpPxZCie
WZxFQMn786b9l+Lu7mMvFQixGC4PHb7ybihrOjDjpQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
b3PhX7OnRtGS5Wb+qkgveIAFuTPa6w5hGPlmb5YELYqoYgkr/ZbS0FeE2yMZ
QVYYKoQYog0cMsSfqgV3QE7R/Z89xhi0HGj0fsWD6IYWgWOs/bFiu2sYzlFK
RsX+OllF1bnoujvkBYJ30bjw8YntLYzY/hrszDLPiP3W/X4mnO4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
BmBWVIIkvueF5wLhmmkXs2+iH3jfHU9nDKxE5b6s16VIzipX5h1879rnoJ1w
1VCXS6lhgZ+sgMjcYzwi8frrbgpiM3b+/dsD485pPkq9DgR1xLie6FbR0B0X
3MbcboNav1qzwzIu5CpBcGImnDJh/VBMMxAgVPXzdj5Xp7KE5Xnt5wOkTHhS
HN/736w7p9IKBJNmvfHCAFh3mb7bmKwdCoMNd4qGkk4hMnb6YC58pQbTNOoj
jVYElsfHz75JOFkIlCfLkEpDxOLCxGk6Jw8FvWY8aoNlT3CnrMXceIIAoT17
5bb4ay5K7C/nVMglHDhiZBmh9C9SbHI4tQ00fY/dUGJdrabjXYnVNqOyUY3n
WqOaNWX/dO0Wh949g+QqzBXaJuC5C/biXu6ySjcBhadMuUQp86e7IxDZI9bv
HwbPovFmhhcwg5KHH+DTXi0ABEiW5fO9ytVjLdze7C5bF95QCdb4SBARJW/t
tOz/AuTHUloiRNY0mvvdTzBsa7A4vbAy


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
T/NPsoXzVW1pNlrDZhsFwhGiqUjfkJ8+0P2Eu2csfdkM4yg9LkcwuXawM0Md
nAW13E8kxrNb2A7DWplfNH4R3vxIM9k9JtroE+d4GX833fZQo79gq4EDG2rv
YZBf92EgmjGQnYibdHJEU72VxI4L1g0FuWrYdN7ytnBFsVTuUVw=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ES7Eo8ZMfcpY/XqEpdahOf8ivLCDo0Vlmc5f9AC7qup4dmiyGdBhjIolkLnS
6EX1JJTJiYLfjificu9KP7hAcwUvp4+JKL9H+YP/uzGZERMKZupxkizYPLJd
LisgHRpNtlA5HmBepdvDDQJwSLutU6LaO8Ulkvy/zwyGWIeesO8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1376)
`pragma protect data_block
l7Hz0YTTaT3Y+RWSZA4FAYl4JGo3W9pz5neCTEUptLwBhPPWzCn19AsRYwjw
2aBMY4LfVe3IPavW4r1kKzuVeYSa44+0XoAWoZSF4Zmhq7n/a4vnbCK6Hm2p
yS3FiV0nyFwDBeA/Mc7/qPcbyveUMbVEuOHpezlaa7Vpc+jY5yU+2SYjPi6y
JkJs6hZRIC72kcmtv6C+Y8T7pMK8VTEUP7KZMver4+7lbtmK7mEiwcuzBb+3
AqHQouFG7sHfAEuu2RHN9e8YZF8rxfXKjyo3JZHH9xu8fxtb5GULwcJbkAs5
Hc+fZ0H7tN63qsiTzgItRtTEhvg8i6ZflcuYK/xsGWn8s7gWqo3zF4NjgMxH
lFJbfYUzj1WfSzWOLfQzDGdHNafHmf5sfucjKBWsejQ20oVxcRBGer0sNvAg
LwH55TfN25ZACnxR5eYb8+dNlPqHIg4FaC7nQ98//VtogvaMNu1d/FpU9O+K
DDmOBKBGyUjAEFQenq/NGlZwI75v0AFvFr2ueY+Ia0nKSI4ILeXlaXIZRV7m
BI9Eusf5Mu+qj3oYKcOfRfkrClzg/xtH4+5+jAZVZK9bBr4bUXVoJl1kHWNu
3UA0xjJAoB24TPfwy1nMSLIXJwx4h4mWol59JoNJKLgFz+FKxpyUjJ2ZQ+0+
4shbNDVZiTvYXtdb5I/+aej9p8CeJJ1XQAUyGJfDmpcxtmQZ6bI0SkEwd1Fm
NrcUUtmIxdicOl/K+d46M0Rn0qRc3+nb2AUOfBeXpmxAqwDnEp/SC+/+7IpU
lAbgI0Xtkgo1uFL11Mq0rGDDKwe4H3UQto+FC9FxZftWF0oKbvd3c4Ggr2TC
EOHl1nUHy0AE9uFT9PZXmbd+L7L2s+InmpvdZVTzb4Prks5lrOoyQQEuF5dv
62ktQL96urLfpJFB7zPUO05o7O+tDWTuLiSWqvA1CxHWgzQgWZk8KP7qFS5K
m70ZGI6h+Li+aSiE6FAxUO/tqQ0cUdhoZgNzp6ZTJxe6UeKGCjMZpZcvxOXG
D8JsLPsCQKfzbNhMnpDweNZfOSPjRtktJecmQrfl2j/muoBH0LccntzxWMHR
ZnuJcUrLsQosofrQMLoW42lh7tCW7oGadtrqTKtfZvWDi7n64XoGCaNvgWTU
U0aXKSKcbNKvuYrn543RTdz1gagRip/YLSnTLnKE7M3fjU4cNCwQrNohZanU
BOAJeOfcNpwNOZ8rTxviZRQx5V0FUsGZW5xRRnKeWzNHZYKojEgw24JQi6D4
QwpeeF8734GdzRQR4n31nG/T3dbMH2mDgxdrilA0srGe9bo0qmmOwwcY8si3
XUb+h43Oyw41TrhxXq/4mxFPj9DmKag2hicpnvVWpGhOz1bWy4B1n+WZtlj/
4y7qVhwb19D7FI1lKccd3iytM6e0OzS4G4fJtEg7DkzXFGrTMsMs2AEHDT8W
sm6bStZV+wm2sBxCiKw2Sm86CFZxgyqnNjljojxMVuHA3hNCAa9ITCCmWoL/
slsgoqDRgyNAbk6ucJbe2sZC9+lYM0/OC+EeDIVql3oUKMBwZKo/js0C1Icz
Yq1i5yxmgQzhq9d20SpK/gphnGxC6SgVU4gV8gEfsN6Up61j8EoN9/a5WLkA
ptI2oRcFIARCWhLfnKj10RqZKNFfoMKCVTzIJBWH5KTvQVeZY51PGFLaTLuO
/17SN+I9Fw5DI4bKNOTCk1GxoPIvhkZRxroqEQUGUIK6YLXKXfzJbHz8aDbr
jcmTMEHEWUO5LnFxuth4/hE4pjGZ7T+BEjjIWherRswoCodE5jND9b8HL6k1
2jNv4mtkdhxi2NHjIE8Kh7jUVhrYOJfofRA=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqdS01+BSb5BTjr+RkNOcwEu9rbyPwxYyGt87tR49hoMTr0TgGndq150qicoDkxYseCPIPtjhLTC97oE/kDNfNLp9J2ciiDtYYMzhcegp60OhE1jQZ9pvyh8IoG+X0ZV7M0zb4yeUNSAo25//J2hEl6vX8viR89IRypvrRqTj0ljUwlVVy0T46g7V1a83DIIWtduukV/V0d9nVIYfKUvx10msCXOGK53/7jAUQg1AAZSkQy6EyvES9IsyBta8hbHlhpX1xfp4oXiyG3zwB4qUGxKXoHVTImQtdOzkeCtNeW0ajcT74GTVByDtL41gpIujn7Xq8LAD1YIwwRFNYUkbLVCusnDb5/Uv2O2vy/NhHpxt6PzrUKqxEuBaYl0kEEiGRHXge00dnIUKZ5DVzFz3XDAhHdNMWfnBCAH5DLOzOzl3oZYSWK53YjfSYLa1m6Rtx+ORzxgTq5JTYz8pgIVC7h5jbXuygcp/dz5VJg9A6XgGutKKXNVd4vxkPr7DQTUqUQJlbSe1jzuTs7pw5ozkt2PNR3fDlQdkhsOIvEg6KtkUAIY8/7ZrTnF0mv30X1psjrm6Duc426w5noj0/npXX9FX5moVo4Kr7QfGbz6NKt5xMEkpPl1uEA9xb8m8UFs2nylF4p7B2ZJP7YR8uYrkQXCVXBF+wwek9koK39KoBQh0qAyh0yWwhngHvTeg7ptiKRaczkckZ79Jw6Zdo+nr0NoLnlrTfAULFZAhSh2eVtxhbplDAcsAQSTJveUXs23K9MnL3J+T1bzyRNZEHk1WiuP"
`endif