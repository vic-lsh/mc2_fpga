// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
0fQtqdJfOXshDhmJGKvZMQVs9foYT17vPmawB24/jNm79W6RSrjmr8vTKdBo
YHVAzVj5va8hlm/CLomBP5k9eOLem/aj4lIjxpsSY/nA4iMLyMAg3LaZDw2O
k2PC/1W0kCz5A7vpQBRyI4iMphtyjhtOa1Y7W2NYYec3igDvPVFYCIahw2df
ejLX82CSyvMujx7PgZRH4LmMxXv+DgPGS7wGNkOu/EcFNX6tu3GzC+BZWCRa
4ynGX2qw1aH36BZRllIiOsqaYe7Z1poBLuzxOE13EpvV4/I+4xUYJBqXwhVa
51bscbkHorDMDqscheF4JNx6y+QY5aPdBJKDOyl6OQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Xzd8Zu3mg3/PpJwJ0hc4rkxuGSg0bGHMqsaumQ59TqTet/N+H00JdmS9N4Tl
12nff8IMBUEN/47x1hkouPfUd4VXnMnu6aMogYJBHKP9FoxMhfGFdIQptUGz
sxjFpOBXfclxGGQvxtheNsWWLpvgnucWs2LxC3bmh/zQmgboyfp8lQOzGw7f
vfPoO0DL5az1pUXdejdD4YofX/LZUsQ18JgRdTpQ+erV2c1nfU7y3mwJEooo
Fty0oTEofM+N7JZNJPaJiJlnZ0A1P+kfVjPR3qh8tGaC84U8ZdU4m5UvUSlJ
kt+YsyGYYm6v5LFEdRmySYfGQIBnC9ccnxc1Pes2Xg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SyTTylhes3tjL80ojSXd2Cmdxalrx5wN/VH97O14kXLHfqIB93VuZm6jzpuM
rzDlz88YxboKiRnEI7VvrF8WEKsr0+a39py6LvkHk0ivDdYQmfITSzq6nnfg
ILcAKSvSRZ60uRt2VC5A9IG9rAWmwuX3cBJ05prfvdczNg9tcaXRbXRz3haD
hUDWevYmYRw14/ds4gYZQS5vjV9vHduUkRu+i10fbn3Y+X4OEksb6eiQoEp/
zUw3WoDQQzpHPIfl5xSKOGycpEQ1U5UHdqVfLkD7B93YVDmkl6RU7aKyNwAK
lyhohGYEgvH8MR1yR3sV90lB7Ya1bP9YfefRNkfKqw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
S/3KFkEBtfF5w6vMR4wBnBps/6ohGz3+2T8w121GGCVuzc5dHCBQY+GSIz6o
UM4VvgZ2riMqPJvn3rrW+FxLVq49pQKuMFL5yUVcK4f6OhrU1JvXTcSxPxGV
XytGj0lzByj2TY7nPrQFCRim8XdDKFIILtzxMKQLAUESBpfEU9h+GuZDNseW
b+q0jPc8JxudiIjXtqSWOswiJqs52BoH2HcGfgTQvxbvUHTHtbx8aTfCStL3
nsSLrTVJlLRmcbyRJ3D3Mjh0S+igkaisA0HqEfzZbqv4EeMymJJDoEdsnrlk
mLZW/x8xzb5CC9v/g5d8sQllsK0psweUoiXYcog3Ug==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TlXk1ldYIFNBaJpmd8HsMt2zX8/CCr7az2DOpDSyLpHDJUwwlKnJ0zAmuD3r
jytXOL68QOy292JRBE30N4WTqTxf4nVWnsJlJuyxxz/awGW/bBHjs1Cepnbv
4/PPq0XvwL29BSrdT5EJ5eIkzY+4s1pGFoGytOkJyjbZgGmBCmA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Ey3dfRDtljp+KBBEQN4UJP8PPA8oEiqoQ5s/jl0/90uESYzV/LD0JEJMdK5N
4vmwQvCiqbn3X1msfTo9+Zz7vVlWEIKxvvFNGlHmCrkCbElChPI5/fQOZqCb
mApC7+1ztJXuEmZMwoG9YWppEmlMOwnpke2sqi+MsojyYO2bRXvJ+yqLUfqb
HzLIrs4Fg0WzILCK3keyySxlHNDNWot9I9NXLrO4lmwSbQkazFTiQ1PUeCo7
Gye3iYtUQa0Q0J0G6KnOk0Fba3N5hMWTknSMr2mDUI3AkC9B8O6kAgI4V7t0
17pOXr5Sscgf1ikPLdYEYWZCYs5awR/pmkj7POyYYX5+cbNTuDyH/312Uhjr
NVRlCbMCzj1AsWsJ1T1aXrSbNm3DTp8e1jIckQBXSsTthPJSiNdbbtrOhTBT
dTKtJzEAZ0HU9XR3n5694+9ApiCDlKd/XkhHV2v/SRJzdDDaXCtb3mThZkmF
GulvHhwbdf2KFQ0nGNQk54txoGPQmciZ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MoNrEiQ4w9EdowpEwwLSvrv2LFXBR9wKtv9d0wfP8tUoJS8tj3Ij7uXR2MgK
3sVg9akYbbvTQdCshiVldKYx/SormJ2+hDYAW/+yYQL8Bh+M2l0fsLMXYAG6
IqCM62NpcTKHplTDGW2RcXpNWTwpEvKYzZwSuZEoiNEIEMU61D0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YlhCYhmxkonKIn2saE7oXwcnaj9Y05u+rY7SWurpCs/PO05MddhPHS0n7jtI
PuRB0EFf83dSK/gbew6EluvTNPpXTujvuUtvD5EwJut1Do05zdPvae3HIJWj
gMiEPcFZSud9fVpnIo9vAYKcYHR5w1iQ4m4FnZg5blNZXFmOEnc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 76880)
`pragma protect data_block
ltRGuzddEOtzfhHYPajaI66aMY3ytjsjmhceJAn0sSAdqSLbgG7/sR1cUk4s
0WH6E8MSWfJfufzT0FMU2a0tj5y09gYem6cv1/30XKEqnJ4wDY4hadvM9gXs
FJ/hUR8BZziFjeDrgp/wiQVd/weVv5ZFixzHKu5SecxIPWZ8AWmi3rfbyATa
apB7cKPJl6UFOg+5FNCDbLeZKbiShnHAK4AqZx1qGGYI5L959M8E79uIRmKW
Dc3QYyfBrQXUQme0z2l6sqrmVQUQ5FwCXvwHkUDESPWXetW3YPgfXiAw9K9t
uhY5AyWvQqv0tZA+hV60LfdQqI+UNW7k74jpw13LTLsIR5J5bRrPBbgmp002
kg1dTQgb4s6P8ryQC8Y7gPj3eVdogS3wHsrzS/fO+QczO7D7/+Ox+eZ7G4AN
fo1efQF12iWg3H0OROHaU+W6i7HK8TkuRMWco+Qg/lR8rEWEZDFS8lcyVgUO
lOOSipJs5ZZxdESFBWEAazknhtgQELR+RjYo9ZOpUPCyeyad1Fb9IS5unqio
VXUlmR3AS81qvEgQmS42ajEnm9JEnrR7gZDfYz9xKrrEUn4Fe/F3RrixrDnk
labn7v5yPZmS7B3Y4IirDwk6vBWVqbkAr12a9Yhfr2KIMR4HVfQSyfVtlofP
FQMUjQCCGcbbQra7mRMj5/4FO4yYW4z5pcRxsSMPZ7AdYB1Ujrm5XriRqdv/
vN0XWE9uOLCTXHkFq/wUUagjaCS1EIPyRwpN+6Vr356oIXR0nPLBj4eGvf+x
ckJiI1Ek0TZ/F5TA5MUVL0rY4qu/vv3FVuqvRngVYbqeHJpETKgb8sxaoJaA
sjuqdPreiSScvsRXapbO78Q1P5GBzHVWFb5HVNXrFjRMaiLkIqpLvZA3zRkC
GyBlMDl+6KcKwmFULrGGaopqQy3z2/VskiqBPvIy+v5ZlP3zZGvOzG3BKCP2
730G7roX03khTgPm6aff5Nvw3uF0FsWzFbNTa5ocNqhbbty2CdnkfViPjYve
lYLnpwPWJfrrVR5niKuNUEEdocFqmVJqKLeeewhoKD2FjvGEyCBSdjBd3kXk
LKUADiQgNHUSR4xCca51hFzOXGINK/C5q1uMRyJT+5Z8dUl2KHB1u4wBiBUd
KhfEqJHhkL1nIP1qQCF9eoa4VD1zZaF7w7xEDgtUpxMToPsrqk6m4maJDlN8
7ZA/i/joau1A6M1uhGWVXzZCLFVjLDTUjwJfhQLaEd/Mn8qRyT4A8/Xf3lHO
IYMyE2Bpc+/In+mHq/RqdRcw1RZwsPfto5A0QpbL4CWxog5CHQtT2xwuGRs7
qq6NYO4kNbshofZFLMFhzjM5KaOVaYnIiePFNdX9n7itc+Zt3xjROzBjlDTy
LWwMLr0fF28zQdU5nmQ2XtlP6dZwg0o/+kx4e22YiKSvvKIwdqBWPOgtpdoL
0nBacPQLq8JmQBbXQaTQ+hR7sV8KZSUDz4+2tepWdoe411Eq7aNPkYoY1Lc/
qowk2vc2y4qQ+oEuKC9gbcGEwZWcEq3SX9n4ipi9iqVcPjy7Rtj4XI3jkfgz
dKackbS83h5jEdFkRetzNMyRJZkDZ1zvxJgsBcoZWCT7xpGIWj8hhOXdeg9Z
bnbf58Xq4Nt4Glx6G1BOJnoinR91TzlG+fQbw9GlHa/o1MURpLY9UqiEfOY6
GQw5fHzTHUZnl1t/tzx7lk+oZcY8jhR6JxtMw6GStJ4o3asEq37kiIK02lD+
MKdn7JtgD436s/1PBcyvZ9vT2vFJwEMtFo+PAkSCGG50osERHidNc0p6qKqZ
lEQXUl3fJ4OY6GJgg1Rttoq0aPn07VF62FfCgekRPGvxhdzmWR+qHeBdMFPz
ZDTxjCHTR3MIDOItnQco9DMcpDQ4OxXv0w0MjeOrh+GqKNM+nYK/2Ba7RPh/
x91FpyOdhG0ZOzyrXB4YQ7/4wUMLGdKU84XIcA7VpXKAOJqli52Q6IcUeite
i2XebsQXDmuwaADX7pmyCPqUmB6iZmvvmnyzp5IB7XNar05S7v703PfUnwEa
csb0IferzK860nOdxe3OjNjG9ppWBFOyDyUUmXFwHyjnr1zh0TpU0aLTVaFL
J8Ewk6/AJLzcC4wzPuBmhpIDtde0t4kntWz0a6+FeaXgjhf29FQQDqv42cK/
xr47vIdKuix9BCivuKvuiQBtD9//N+4fmH7+lCm6bH+QCEkMO9Ri7kPrBqZt
RGYtWMwflSNaS5422yLXc99LPpWDBiJ+PRYO20sZBElaH/gmbXFcYxmOCrM4
5Jfu3DvT6T2ik5NA1sVUitiAf+LI/EhCsQpW7444+7wShCrEtmBLJlh8je0B
MfMnqOvITocStfGfZZHVuENCBJ6q4ocEnklzL/0T29TB0h+XYqlvqKxk+dmN
OJ/nk2n2/HJSoa/ImB2duou7lIgLF/3MwqvCjki56/4zc1pv6wtDOcXzymKP
is7q/Igf0HaQdPEBzZ2boHnVUXLCy5tgA4bEFXRPicKstaad0pbZhmqyUQYj
m4timGJmLN10nOKI5XZBNCI7EzuRUxhiZGXa7wj2FjeG/7S/5j+8iGrHzfPC
3pE/cH4pXqkV9P3q09MvOnawFr+urwp+fAc4MW/ZnEGa/lI3RHN1ckmfilxn
Qw+h2zC53ZOXE3q2rV90GbhVwGwwnXqwCN277mfce29crHalkymt+OfJpoGF
SpcNqQiM9E9nR44ktFH0ZOVSNXzQLZkqpQGfDmy+TgqEZcoUTrQnLL/S89ow
B6zlo3oEh2nUoMN+XQFflREMSk4lronGHkQIVh2MBwsJSylvw6gsdgayd4s5
NEsec0t8tvji31b4hrsfBSLzjrILQwn+erJKCcowJGjKGZwldCNE5YDMlHhh
j2MpadRvOywl7TuiqyxsBOXVpYNiKEtSTRrnP+HQsSyB/V0xRLr7r0GA9Pz7
fkdQnT7HcxS2sByzubLo/8giNLR99xG5+RNhyPFfB998ASc0yWK4Bwii+ouG
3kC5XM3Ph2o70542a8MfxSUL5kbWMlYWfzuwwgjqx6uGt964VHCv8JJLLgSY
5zUCZaOkLzrb8Tc9LyPhoQGtkXUG2fD6aI/EIQ6nrkhZZCg4qjhkHURcg68U
ENreiB6fKI+jiLpN1k5durUMxiZsyHedSdaoafzJ0fSfaZYMRAnEtYH8aQZm
1oqXV1Cr6+g/e81+lZewNrYfSvWXkFJUhSw1Kmmypb9t33Pj/ZGMDysjlmbl
/SqsJBFWdd3BdFg/kHdIJT74DrlV1BhdSsH9GNdHAmmtHU58xMLd43j6PGPJ
AbtSKtpyqMkmIse4FmDKZDPlOu1/4C9FAD1tQ2JRQ7O6a0W6bP0Hz31990gS
lrpstQY9F/RHDOnk38rIPOu9BW/vL1xJ5htxsDCoJEHvJqnF66kthBTEPUxv
zi1dx+eCN6zXNcultDA2GYqpQOak7xCFNQXIzvgdeiFs0ZfRrg1uH+TF+1fw
OwhYv72uNTXWfQBQlivSuT6OPg4Ykdv1LePKyGcP31BkyvOqBc0PVZYQfdj2
CrRNG76y1NMEjAbx0E12Oh4Kg6fE+qxuRDk3j03FKInNQMCuD6EU0mY92+2y
gcYaXtS7SYQLoEh+ULhpJ1gthlwJANzCgy5UFsOL02nVqsb7lP8bDzguvXy0
r7uyc3uGVYEV0LcCWDGu0M5quOsqzbJmsqPzB2pIEiefaKMy/l8EaDLJimA/
01skAic3bDhjWeG/6dn4E3EqTgrEvkiNvBWC4XxJ63UoBHalF2IJiXIsKMso
W/moCHO1D8oiec77GXlT5yRzCj1sem5WpiQ8vzJkAPqNyS04wQvkEgFKsSJw
JK4mZ0bPgdF4EcMsGA2yfU0TsqGef2Q49mxmpOWz72Qbk9B2CNLvMZrTJVNG
XeFK3CztiBNp3zO/u1t++xhsQfMDrUk/gvkGXLA0PaAkAQG0l+JaKEGW47lq
hvHNDXv9w6LtyZD8O81hI5uGDXtwvXBQE2oqpzZHCPU8LQTqQYZHW91fQjCr
thi7osszaWtdxs4P69iTodhI7xWnAahbwpFI9rKEHcclQBYf9cq6d9Hgbav9
J6V8r8hKtoEl36jdDJvVU1P61jQo2lvh7xgh9UMWWfkfOM72i1kwnI/xiNO3
EU3ENHa+4GGRBHo9ssgmXWcyIETdRhAX8jLwvltHZy2OHJqGNDo0kMS/BcOg
KZCboBKHrHiXBpLE481SLHsOsYDlKN65qDWIVYXa7S72PGwlunAMt6bLIUKo
1ioKO9LyDRJKG4+x7SClgScU4sg4dyxR+Wt/JyzgKVm24uBrvOP9sBP0Jgbf
2Rh6g4HC6mXAKxuSguJABOdEqzG465kkp3aSISnumQPKJEorABRG8J5HSvkS
wUnnC3DAEZzm36kootkDNolfnf2xnsTpNEZd2l28HV5di4FqFAzZ81DesZT6
sxKUZXgwt8vvajMwdKnvlhd+X6c+Rk/PZWPvDQCc9/AX2GRZy+3L6DzGSieH
cdeJrp9PTYB3a6gb/SxNHKOlksb3xewtLVtTYJ6rryvGnwFaV7OoYOOU1aHW
rMLGcGACNyuntg6lRRoNov3zQ5YgPV3X9g5rQzwtFwUqsLZmXxmWlDL2VWMM
AqNzoA/MZXTuDhriFJ1S9hMi7ZzCopcBDAQzDZsFwK8XpXNb77FgTt/8Ln08
epchKJyeiGldsEa+DmfKeP323StnmaJTP0w+PagDMuUL6T+ofAcKf3aQXZja
lmzzAFr1OEc148vPPIQjUQxQizP8es8TUHu3vOCorhaSVpXIe8Ttb5EvG5zn
0bZN4v6lGHPzs5Wp4aRdPi6I3IjigLF2WRVVOas9VkM6/Ldff5ldCXWcLqpT
bwDQbXRitz+xFGHFIzdXNOaRsY7FgfAMDgMr8IkdAGuw0tm+YiKfeuV/lPjE
ZXHMFPbHsAhGALOgpcN7UQhIcjdkDB2U0T3eMvXb+7w/ylJVTQ+KSJm5NlVh
bcjBpxgYRnJJNK3YAo+ABJ8bkKp5x5APvL1lw7be7D6RtpugYYnw+95NGrDx
+5pIRs/7oolH3KFDwsatQ64E0hDqL80W7RAYa6dbriJOdYqeoOxK3ghNL4NH
rEfl+iFoxeKqrhEl6vmm/ufeGoH7GNyIXmyMDb/w26TAKb1J9bRB71T63nRO
EAK2axGEUS0jv4RdcYWJM+ssE3lh2dLNu0Eyqwa+JgHcDxDqAQomv+vfRycE
GXObH/1FWNPSO8Fd2x0etFsvPiobQdh8tsvBfqv5nZdGWfbBIpx3BugNbWqk
Rm/8g2pt7yFCwsYJIiKX8JV6x/8QqTKfkoy11iG/ItBlG6Q/NuPKLsRcu7S3
3B2nxAyiqo/TsAGRScyvDCXSOt+W0+5z6tcwz30tJS1h02TaXBderMm+tnbO
xPorS0v+6CvxdBZqAJCH0JjnKjAqFUBMTXrGezf5p+Ig0/HgrFJH3Ka7UXcC
6AWxsENINRiQ2Yia8fuMOC9o7MVWhuDpS0Lg5q7ufHIqRCeP4P7PzT21i2Kz
01pVXJTTJrkmgXDE6D9BzLssdNRVGyu2MqetGprgwZmo4Pp1iWnmjaUl5qzF
ng+GSzs4peH+956chaOOMCXCBoh3UWGyKoONsAVK8a0jDp9+V8aChaZMAJHs
StB7xJjxSlBTpgMUP7up+TkOIo04rSWzRJZxDlokCqJcOxb0JRKH0VgQxwYh
Z+2JjDEzpB4ZK2fIdFG3Spn5tq39c7Qqr/0j34t0fUuL56Am1FqBcvCkOr8e
PCf08dDFBXXB7OPPtXhNgoAnKsQWRUzW2fU4dNLTVs8t61TFHyud+D3j3GLA
qSEdZ6Rzm9JCIW3bKMLZ9ttMtOBv+X/IYcNq9OcAYRU9qRjFUkD9RhWueuwm
rResV9mpgOS+ch2nCioDMIXZMOfjstNlm92bWCdHXosLyaOkCVgsRTRTGURG
itDRgSAu/tl5F/HwDe/x/2ivplBE9kwblaDKe9YRTUUcj8tISmOp9Tkq3mBP
6aR1LSZVvvG1xAJZgB4lRar2wjm+9NTJlqH+jsmXNwuE9NGxJOAXMcVaghzO
b/gxHWYIXXnFoEBtuUqWF7JcboR3h4NF1VAqgPOe/g/mfvA1ll57fN2z6AIE
+H7fRv2oz4zVaExSKApMw7e0dAp9d97PfrgcMJLGAoZE/hm5U+wCEWGZvXx/
5PeowK6plLWj8ZC8Zs22braUlN1yxzrx+ujJbRykpop2T/P01mBO0hAmpTNn
KmaxWNP4RHQgTsXdQsZZ8krhKSk9JI0zXw7prvLpo0dCVHnrQ7900kpxdyb6
fsTzdTXwpP2hidHue3bw41RW2T436DWixURViHO5qcuhKdm/YgkR3RkGeQki
BfvmJSjKYnFmpViyybZnu4DEhlUhLz9YyOlCkeQ7v2GuOYGI7f0CrPuf5Eq6
clDLb/5wHyqxqhRJHwOkhP3KhGVKvjTAd2ExA9r3dcN120e+HtL4ZN49QR8Y
XwfUPQtprOIeQSn2aUxyTxUSWDzZ2hFN7orvRspntLYuiK2Z3FM68GYl/IOb
0MS7unw5EwYClj0CFzdsRexEInhI2pLWaW160VyqYT5rzxb5SLjQ0cudtOHe
CTbBfPbKPty0hgsQ/HX6dG3S4XZKetXor0ATqUHuZ2sTvwc3OhLL9wTH68Es
g3UVzQG9YYAFJxzFn1RWYNcZAD5rXc/EynpVbEzaJYzetSHINqcONoZrVm9v
jmMFwDWwIeBuDLNLRMASPohAJK5qTdfTZWqBM1NrKZYKVyHaFpPX2zJVP9/k
9eFQBOwUu9/29gfgJ9AK/e0sdN9mR/a4MoJxARJZeKmMf7zsBIRVLLKYRP6Z
eVYmOQK6c4Jaj/N8JYr8cEQe3QdQ3M1VunzB41g3tinGvQ2Li1aNGTHpoRvU
ZCY0kG7ejE9HcZvRDzduOFhCI69Zsv3oxIMieDvLsxdQ3pytFxOEtByRVPMq
oaQlRPbZoIZ6HG1V4iMjX3zLKy5BGeF3rWOHU0xKB9w/Ia+/I5A/Jdclccfy
0buuiB+E4SFRmRrs0TNdYoXjy42rVYo+4boAgJzislOf0Z4w/p5mKT8rezOn
aAQ09i6IyJ3SLKXv41p7ZwYuCSSgfkK4NuTF7CBnjNflZyMrPfq0qCzqH0c3
lt8dXYi43Bzs1aAzJq3ZIAv0pQUxVFJyOlTnTjphhBzWmT1CLzLES7mEvb+y
pRPky99YrIZoKgP5L7KTsOcDmTVfoHpaeWoy99i4hz3DwQF+/pNdso822uwB
m4ZfY06Om4rq00JJULhsbZ7woJz3iuM0Z6WnJS3kTbUGAYDJXPsEVT3HHrqz
rGcx1RKYvk7HEaLO7EPK9oWoYHpMFDBc1+TJrQDt6CHMby/9KYtugmWXFll3
fWObqNs5L0XDXV8cbeBTJ4N8Y5Dzl0H10YowEUQDYsx4ZanUmGh9femOcsyo
XiefWzpGKUC4doTdli49BX0fLlK9h2VK0C4Y3sCUs8AaRYnWO641T7Pvdj2d
VYAFrwiPc4WLXPLDxMM6lSttJBjdvrj1cbYLsTS7AaDw12zC7pC4eYWwAGQT
6onrka4regQ8Ar73pggCPm5inRPj7IbX+jcisCwC9nCWTuGwOJ23lsw/mFJ7
JLLMRSkGZbMlfpvYJXCh1zcTbtjU2+CNnzQ/vp9Bq2mpsJGT9DlIsoA9YTOs
/v8/KgVy/SY2mSpZUxatMPDplSfA0WoqlJ285qradKckMPHBCvSDA0vVnWf7
szNx3cS5DPTSNsAV3FZsaEPhJi1qYcaymArimQohp6cJUkfXdOqTEp/eZTsa
DoDXSh8bTD8Fb6oJIvsNjopFvHGw1sY8KPGlnAH3HqO/S9rk4Z7Ne7cOE3EY
xtw9BBHrmoyhKn0yvmrnOTWwD3B2r84DIZxZUeHkiGnGHd03dMnlYYg34jAF
rC/Jt63PxuSbAe6+hQWBuBLmAMy7V+x1dCQOct4jHP0pLe/yskqW8ymYwiQi
+c5Hl4rVV7u4ofvlYR8nzGUUMBETAmlneXllreMIvXroHxncO4aK6JrRUPYx
AQo/v9olnq5XMglq1afQi4bxB/LtJ0DXwOsGmg0MywQv/TJGRRtTZGFv/S4Z
khoxVTQfmbDSFrrA85EyuwoIve2nXIlNuNzwTGonWcKFOZWd5BTQfFKOfC4g
5sog5ENgBVuryUkxgM4W4SzK1EL5l2NU3ZKS2moeo7xlmdn7lxT5wUeCRS98
dhYPEu2ZR8UPb1GOkWwfyLis/hYNI6UmOJt7RD7qPHJAYssXt2D4CNUenGtW
N1fN0L3f5fVeKysK11S38Xk04fYPQkCzFGVE4XUJCzqQ2CnbudmIvvOCm/BH
IDjc4129fTOqL8n24fXtKoxcBNEwsDyCcD6EVf54w5OE3dDP7nawe4l2KMil
y2AipA4cwO9+e2lRpq178tJDF+2nYQIbLfsRMZh1/294vNjLaqBoOIbdEfd7
xAU5ovpJJatZ7c1/aPBUKCQedINoj/bMQ4ti66GrNyVw7NPE99k1ZbA3rdCx
EJeZLyUSevz0M2JKlSTVSGaSNm7ZzyOJcujCQyFQCHfU1HI0auA3WEKPa1I7
S6TOcZkpC7J6kvg7035zprpnYCaq4sreOUXu53Xx++j5Le4IQKRMKO4etRMr
VzRILUU5P1WMxtoOmr5ZS7rsO6rSX/DYhM87MnyCJ+qniJrnvGyetdzyP46T
Xhwp35UoNUOjOYke5iiv7QooEOsnKGX9KW60PqdrMGQOaRYPrbotwK4E/Yca
x42cbGACk0A36sa5Fy1wxzKKBt7X6i8yBDM1SYaogchQ7okEzP33t2QFe8f5
/9CRSgAhPUGH9q85pgmywqX6p79Wx/sB9UvOgyP0dyXORMGIyBwsj2XMzlky
FWFLgteu+M7HGt4PtSmhwLDDR3useBkMvmINjG67NiN6o3blzMdjCfk9PD4G
Urt7f3uWOXirKl9LSb/Ohph9qn7y0ChLY0PanU6K6x+2sqeVxjhllX0RSfFG
OdlWE0/aFwuCbfEIllLTiFHz9B0YUob3b6qjUb2QcqicZT4Hpru7xEntAa2D
lN6Ui9I6xk/1sTMEMMyPp6aI2APMtsrU1NidD4EhzStHsdXI4kyJU3rF3/30
PGxzLhPdMqGh0ScaIpyQCSN6ViU/BuAPFHzpcbtMEyBvNvclahRAQi2R9wm+
7dOaOwJC4PG+ElTLSM+/BEHBJ892eDc0eaIrwYKE7a1zzWdiQ22UtOvm3HbO
eqPQ6tW28y1S1b4cpB0bG4v1xZFKkTu9lSzD/uKCWiY7X0MJCGI0zM3A+shU
KMdy1xI9OQfVNaVdRYhiJf1N3Iter/ssdiDZECUh855i8w6YtrA7rF2S+ylG
yKZkwOtHl8VaNw4RjhlIHhuJvZGlUO4uO4+MudgtUfJ/gUg+QQJSTBDhr8jC
7/cQxcKRODj8nm0Qum5u86Jd0SlCUYKOpKkZOIW8z3peliEeCKEPYUXHuTMH
aE8/qN42+zVd8i93zQI8i9P34p46p8TV6Ihpf1s7pJl9VLHiaJx5hmXzxybo
xhd6yFH6J+QQMSy0YpfPo2Ejn5lB/BX/PDaEwodFl1ftWKSJAnaPerTHiKnZ
3VUqRmvFPPH45JJsO5bAoLt9CuGF/eda3yNOiwRvgPie0PyGRQjcFu3B9bwH
kj1E/PheUOcx5sh4bOcLo+tRXFhJjNbI4O+JOSz00x/XJgBaDsKnWGoZ/6Me
pVpLer0LHfvySePlhi0omM0ZGFDTE2rrXNb1WnyrsTs0cUNG7w66XhNIqJpU
tFLE+aI5GP1g0pVo4uqcgT+/w6tbByqixBxNnhaQzN5Zh++O6lM6X1h8P+iQ
kjTIDQrmKWDbl/kW+lxDRzVxCcxC2xuohnDQBC3K/kLMyuRss6yfdjwS0YXa
Mpq7MVumA/pcEVG58AGhxWvWnIxnzulVBtGThX/FNqJYEx28wu8viabZ1u1o
jmnmHKshKF6mOHVmYBS2AlTeCGEhMJF3gMfNTLGvQWhKfRr3XieobMOuq2xZ
MIRWUCBwjoLHdKgWP6OXXmm2ZfkMNgsFkwqaxnOwb1bzN4/GGghiZl2vNfMo
qE1jf6oQ4f8acWv5SgotpVtc6SFP3eMv+5JdtM4VeSMP54Aa00vhuk+eNO5O
nfDPCBPHZ8OvuuNO5G5a2+jp/xot56p+Bn+GJ3X0PJ+aVanSxp+0jGRs4ZVT
I1i4cXB9xWPvfIty8BhmCHFxgVKrBf+GdlNKaGxyhDtUOsk+QeTzBJnMkyCw
iXv5h79/mrCBx15c3d3MPnjyVOJZBi8b67b/RztsGGmr5mQXDLBqNGCDbJMU
lAo7FtBPwN9tOeETfsGxNOCxnI8cyoLLsZCEqf8lh1LOXQe2rCHBS9MxZQky
hrmcApJ8dUQHoszYbw5S4AxweY89lQEI3DYuKsfXhuD9a913N9lbCzA6exZq
KFIb1v8cCh0BRB78qrvbEOXfCH0Os38cktzMSqdQAKvfD/czIy2Tc64N5u48
cZZEEX1FPx4utpDxuq7/4CLmrpV2/mZBLjloeUzK57kTVTuZSIOm14W+l+XB
4sPFPzB+X+BIf46xdD4HdyHydpeR8WaJYDMrbkjAXCVHqbimfHZ0AAkSFf01
tHUE0ESnNYz7x8mhN+2L5vJ1yfxOK5SKA4NEMJ8iBovNXp+rH1FiKGmwq5/F
y4KsbtdzYl+YItP9lGMJpM3/SoxGKKSN+OsBKd2NIgf/qAyk06GJ5grEGSgc
7/j9tMkaZFFDtiUhgtHqh03QCKpTjf6pzrG4wO67i9blrmDTGOn1fGziBml4
1wuVOubRD8vjD9saCdXEKhniV6vxHfnMbdQVJTlatiF8yWVtgesdbtReiLoK
tpb/NR5ywtk1LSQtm6fZJ4f2eoTrxGy+ujc/AeEi+SShcX4r1aYzyeG1cYyK
08OIqPyBrXDmHddmxP3Md0R6WKiVhXAQkJ2Sk93o9j/iBcoAvfQxp9CCVAAR
ckRkUAfEMVA8yY3Kvdl+BfPFZfT+ZZPPaRupWFouDIMHa2UgctjjlhASDQpV
jBu5EO+O38xCxk6WV40gVE0nl97VvjhS/6GdqPpb4f7y34D2JtT3+l6/yOtu
Flq4iQDakhO60hO3Aa/cU8GBbz6V3VekDj+R7vup2e2J6n+mu7KEmxTWA86P
8+FhnyRJSmOL3iXWXTSJ0/SMOKGCxgc5foAgL9bjO4SBKiypvHl+U+DfvbM3
mHBkgZCz0cHUO+DoXjHvaGDXPzzXKw1TIFf/5We1sBrqXxotZ7dXhdSEjX4B
GyGAM2rko6C2mt7WLt+M+WjqBqAGxXzspoGCQmcVHXiKMpRAlRO01NB3irbI
1xa7hnR0o8VdArOungIJ3vc1BxlWYrqfNiGQYw91LthvJ3j4vXVuqLSdrMxE
0PU4oUjVMP1WqDsFHVnPnHijiGdYLuVHQD3cjwS4G2pSsPLqJXPuq9AVSIxJ
naFpNZPHXqbn+CeD69miVtPFML38JESTY4FJH99uaCsnLkBiBHw0r6ZFzBb5
jKqNhgG7Fr/Y+Af10E24T2BSY6fN4ewmhvhpuJ/Yv4dXCFO7Wjx3OZfluwY0
VwaeKFznpsl1AAMHZndJrasfWadGX14BTEztY+83wb7Iv2nv0MGfanqZMlxX
J7Z9CCPwEK3g0so/7uYwMqoFjtGuG1p/JT2ZPJQbH8ID9RNPdwnOwT6TNhal
Cw0g1P3CNZV1ENHTXldOzO/ROWrUZzfk7abybmnJdnH881H79n8mbm/MpWl2
2apS5SrM5+QokH4I3HivBVfcVs1NfrP06wbDMEd3DCJrML6KaDyQmTsw8+xb
ZwlzCziDKRsaEljDijIPMxVWH9PUVPTLL5npPQoR+x1yURkj8P3nnAdBtarK
H4TnAeVqhvHQenvDyiy50sXwX0ztFt1SU9h+fW5Je49zI+FZoDPIR4XhX9WO
jlw3DjydmPFNK8mcFFRQcmZKgG+51FaxdBH2JbTI1DWWjzQpHp8v8VLkSIIC
qnE7ImAZmMYEzCaG8NAhK0P85amnF+xBjBh7m1ell0cI0OyX8SzjoIxnqvDM
wCKitZIbFSo7hr6E++f+EuOASSpTj6dwxBZ5Fz8CALZCwSjXP6D2Gub+hzN+
6eQ/kTVu4Q5o3GRUuQrk9N8HA1Vzw1Gf54UAQoDNSd+fsqRV1+GvznxZjdpO
VhXZgwsnayfiRZq04ohk27Er4eF9xqQXkRp31J665HTTrqsvvN0k3zePW2YV
Tc8+ZeI3dSYFW5SjXiboMkvPHVlGy74Jk2uuASuQEYsLzm+939TRhtBzas3y
r7qpLdXPdBuEDHOEpRWuMZKOeh2WL8fcq5/ZwiX4fBm38YbXmoZX1WP7X8x7
COU/k6MyyZEHqfxLqga3mR2JYdLypHF//PZQZu28JoWlMcx2OwhsQ6WclPCR
fAxUZA/hV/0Q0dBp2aWUX/EKg+dO9QC9QqdzH8WINFTyYXdErarCZJt7aNdS
NpNCSDDtYH8qJoBLswaEcrhC9lvvn/0rCHd2X5bF5Inzk4ESlR2xjqFM8ZXg
t0KfLup38U0MANSfylkVLUyS3vnbVq43ore8qPm6KXGfpE0XDE6mn8h+fJfp
enGGUEUqcJJjYaGPr/7+xpdY2hJWaDe+dNucOXY9nv/xbAOTYmPrWD7zBMdv
T7PyYesAU6JdiN7xqqCCnvJIFOmlDvfyWbQ5b/nXkG2Rj8DdkBarbgxeOuAr
h6luA4orND6KSMvwG0PKuAak13A7hp9ezB6rqqEMDkZOE6Qi2WF7uA4i61aB
OJxrU1MB+N/wMv2YQoq4fepRkaGfPeI4s/9iXw8BJrvuFjdb/Sle5NylSknE
oHhsMBidbpF5Wre3t+iTW08o8Nn6qxVmuABOiKi6apQPRcFgD6I8XSXr2wI1
DXRH1HO6c7RqgUN2JiBfyOyryr2wdmvPNyRqqHyoOsT6Xk7LChiwBQiIvC8Y
FcyC+h8V5WFkLIVRzBbXdogbS0zUlT0qBxI9WKvRvPxCY39RpkP87EXVmlZI
NNPiBjA4xtk5ctizmdytZwfOjyDOpH/iT6ROVCJPPWo4EY/vCfvndL7A36S3
1dOyIlFqtssIARP+BGU5mAHhkinheJ/wYkAuYyHShykE9Y1GOpRtVTUmeDLx
nDYDWQP4bt22WUMuiOVCMQU3nLhdGvhTle90GtG2YnD5jvGbJhTW+CSweDUv
aKwzxClNrgglIWmkdrL7OfSI+6PlBVIEuEG3e1yvuITC908zp5aM84aeOuwY
+viGt13OUmZgU8aUkRg7c+fTd183QREWDTQrr/j/eW+au6xO+XhcBXGt8FGx
WvfaPokRTSHSzktSdNRVU7Ha/UjXUuQsqEsA/AblednipGfDNks6FXPFMQ5P
di5BmmI50BHWJSnoz11mmLaWpzv3LCxzZeL1ZxwK5ICQ5MhGOJfZQR6DsOCS
OUFQHtYCGBmHKGwYKonXo6fg/JH/ddSthXYmlBpMM9E7q/QjpoRWNhDBS9RX
JU78bYAI7OkkKSizzJYVVbVqKbKDirbfkjrbLtfC9Uok6vB8Uk+Al0bNo2YQ
WPJ5uN3U7SIVf2Nmvw6tVy+PasMqsnewoUrmCQRdvvRymn98hWxb2i5Eqxta
NatwhMBlV5j4rziRI3KoqAxihM79sUBkcjy9+6ppUXQaT8gM864dy+8PUwE/
34HCbn8juG4vlsmyPSy0sSXa3L361Pn9or5+l4Y1FstjXQbHn9VG9uv1eB+c
uTtiGnPhsv6DnMiTwyfHZ6DK0oAKsfEP1D4CGfYjQYXpvjEsnvROO6sWzGgd
XlX3+teNt4Qj/FzCVurOwZzD7jlvlw984x0ObaIyf0MFqJ7Lzv25ghi9agJP
sYh53/OTGhxnYpTTibmvBAi+Yz0L5l1WIOZk8QEVZ0RXnGA/f/UH3FHMd7Jk
wRpf2O21FcopVF1AU+7WHbO1sPJw5HLl7hdDrCtJeePZBByzLGcQLOpK2HHf
VIOhXIUiJku08ihRgtPVRyHpo2lYfWOThZNNhzyC88GDyVwSsFRSXgBSO5XH
fIj3pOI9riWIl88VwPcmA3uFWqOx6AbTaPprlGsgumwPoQph6b0jAr9JxOsH
JKVPr/Idi57PkySh9FsZAk0hZj1uhCCAlwANXP0XWGt/1i/aHMenH+a3Jreq
q+hlJSSQzktridb5Rsk7GQe9w778FkO+pWK8Gmg6fB8/oWyb3VPlmqkgqq0X
fLmxZeWgNyH5l2M3QRRj8ubn4V11V4vxA/qw67R3qWrYvxDNzLG9VPuVMHDc
SUtUeVmw8OHdVojWFsZhpI4/FK8Loe9qxwSGLsumpFYN8niWUC68ovW3JgBA
kG4ozQhr7rYDrE7qxCubR5cFIYNKq36GnQsBh9IgoTEI0BLj4WVMr6/jf69J
orvxOJ117BRU3SylBK7aTl7CsMhIfbJDxXXfo0rfWxYq3yBkSQoL57q9QqNM
UgO301vlBUUpmDV2FhFqNL/cU7u/IqvJhQMdlrts+nDdA9h1W3LpikWV18My
MFXvrBARVBOjZw1Ud08q44HzVoTxvp52FG/7nqFvldSRum8AjQNmC9BUjQU8
2fKbFyd3YaLm+AqwIbDpwYtoahZf+P4Ynldfv/WrL8q8Lt4uDG0gmtBnhTLR
gNkTWZvFSnEBDx3kHjlkmMDkogjkEpp80C/Tk4B7QgrsP3k2uVVPRCDWeDJ5
hPSVFhRBaQqh5ktarskwa56QAU6iIZG3ipcLd6Vr7KUCdAq7zGVox5let0xH
s9Hp5TdjaXsJz0WZGLrQvvy2JEgMqBX1L9mY4u1yzIITWy9Wf9OmM1Xoabux
uLLW+9sNj8XkOVs7W32a/FBzlRuKjZy38aJgPtsbyx1AW8t9lh3D6FSxfyIg
gYZIiBo5JnyW2QWMRAfTvZ5D9rcpxsHjSCv5+0vtckE1yYTA/XrvN0TnU3By
ZGqQS21n/83e/Mr7opoxLsaPixDQJCh8PHQT515e1gHhlvI101uznNYqWKrm
zHL3T13T2pVTwH8tvRsf2eUb4NWO2oZVNCYNZKspbWrqMJk3vFHQ3mC+Lfo8
Fd60/4IdO3eujUp9dKYY2K1s3b0c5b8o0rxYl9imwcOn04LtRdpSHga5Sy6c
bf7l+i435XKWYpnocb/u+A9kUx/4U+xtQIt6HeiEx4IRui6aLl/v00kkYTre
IA8ZIZuyQaykTKwawdbG2q7p393ZNdaj41easxuMSgXMFJ9xHRKivnB2G79U
goahmVH1iVXiI/OUpng/X0gvbLAYZ5yEF/UXEK+ibMUTk2HS16hR5R3pI09T
6h6mUdyKgrxI+qLuWJ7CS/9a9DJhgz9qf9XVomzFToZbT37NuJzje4CUiW6y
CvByizPg2ITEFlPCGCAIhJRRFG023oSnXy5QEeCY41id9WrDeLPt+vbJbP0k
I3gdVngGKEunfsE/XxcRzhwZ1fIXMdrApswnYxLHBhZAdJ9hgKuIWlrDzraW
Yx4EMTwclCxxshSLZbGXHi4BZqcjWJ4gQH+OWA8HzGj1s2XZfwuZm/pyWh9b
KvwLhs3MqN2rysZxP0xUR4c9Yes3t2I7Ymu0CndfM5hph3HK5KZnfB0sCcwg
7Rg+ZSHrxiOhxqzO2eOZKh7r+fFmgGXqqoMEen8i06I5xlXLaVBWlQwUhgxL
94w5CKKE49kryK/oW1mV/KUoMnB0mH50SRl8QzCDjCdEhNpBFbEwGAJh8Lsn
kv7IExA3oJT5nfYLEIvJ6H7ph9HvMLDCrkRfD3oBsEj9UVWuZw3y2zPS34gL
88stNXtT9VjKm/n3EdLgZVtVFT39ZyPM3Lqqkj5nfpkhMUz5k7EC4oEdu9cO
VFRbijpNn3ir281ANKsXdSKK5PXcvNZ5ckOxxQ2oe9c5+YdysbZPUtJHAcYF
Sdl/BOXVpHlP4MesvO5SgGeUMcOFTC1u7D+C8d1DR2LK/DoMXyWe9xsLkYrt
t3W/ODj0Clpc211T3y98sPy6KJ7HlbGQzbIAdmLW8B2pIhnivmvzt7ivN4SL
fsByVzEGKwHaYj5xqDL2HUNkF7ijuzMzEmMNyvcaJfZMVBXmO6DkoeVcLSYn
aQ2YhgxMgPk4B4ZLsY4G1Iu3ubFtLcyEEyFnGxHot44o7R97AaKIldel76Zz
BIGyyi1/psCN38ykpLxr/XbVvJiEcaZeg44phfrLaU/j47UzQTliI7Hb8+02
L0Iqz27/7PQHjYnhjNBTrR+dEIpW8/G4e6QTLneRlOkiN4Ehr7Byq8LD88sZ
pNxgXjKiz7s3OvIkySwjuVA1C22CAvMUQy/Yj1L1MTfjYsYBtGqitsQCM4cS
vcPO9rll28IU4PCwuHzpFClfaOVNz04ayb7yCeqsgmM/nqlSrQkrmiIJlXlU
MMWmG5j4YTgdT+jO0CLbaL+KKbtzD8dkQBwBwiWGfx0A0LfCq2tP90Qq4Isz
0i2J1WKp7f8rQHqb9tt9Gw+T8MI/M7j5or5UEXpOgY3dmzZm6UqBNDq5fGX0
6O2019HBbSYRW6PHw5tMfDEXYNzY4dGql+5YfcpalWEa3zANZCl5xp9ugHvm
VkttZIaVlTCz0Iwy6yh+LlpS3YbQ7dVCRoxqjXPDRfFCMVRKlXtTy6JPi1q8
Hk/ut/xuo9LICup+Gggd1AYbUnuwEBlIL0kGbCyzBuaX91tccqeuxepqKTx1
Gp+Zp/vpiLNb2cHo+/s1YcVYgIdfnaZNlbmispOUinQqsEOWagO/TG0jfZ5b
5OVm25hFb25zqWRf2h6XWZ54g462P4riGxCzYMj4FfGJP/WSYsXPjIlZYgwd
pavk6LKannegVoYduoaPWT2AYgaB8KMeTRjBjj+eAO0vSLdd+yF5Kh6cWVfi
XGmI+vNfgydoNkxBz3sRdw6DoLMzk3RbsNvrKw1dXX7pYnTs/5jTeWXjTrGf
dFC78RrGL58fi8a6PGxPqxHFfB5bWbrQXeZ/DcSAO6OW9qadw/qRNQoN3QQV
7hDLbHnr+hd7h7IbHiXiqPPwmmpUnxlkh+pvfAZkOWD7/v5l+pY6r4eX9L/s
6uumutkneSery4atMAAGVe10Gyns2oJIWrHqb2/tEFh/lSe5ZMMuD7W3u/WS
6C+LovELxktgnyMkGoZccGYBse+KHOS2+BM0B5PubXRS7eM+cL3ztKYBGBtI
2ODT0/e1Ce2sveBdW/QtnuUBoGZmFNJUsHZ2azyQIw6tEQDcSViHYttWhFPb
ZaXX39lcHvTNqa5ppoOwmqYhyF4X8Ypv/oEEHBaE9r4wu9/da+vxwq7hiKK4
08Sut6ibgMdVBb7wp3U6nCTZypvQ80YkSkgCpVYk0YZk7STZH2naApOSlfi8
AOwdI2vWZU+PqUp7Pnsobl+KTy+RMhJ/fktRJeZuec38pvVWOO8FlG+wnRnt
l78T/T/0fGtVzSqqiNeM9XicW79l99LJrQf9oEBW9VLHidr38jTUshDnwku7
KVQlT8CSa1STY77tSPkU70OSbipw9nRWvMTCoSBCq+3L4ZGhznb5SlgSYyxP
9Gp360XX7ZY2jPrZGeV6IrwJwrQCUUyV4pJbeUG44mzQ5aauqOT0NN10CpyV
wYca++z5JWAVGhVv5HXkS+o+pHw6hOXT5qSMEWHOX2z7DYDZv6M37wNX4emU
Nr/5gDnvtcXLSi0G9Rb3tfRlRdjJNBadKpV7Pel//ifmVnD3VySYkJBwBlA2
Qp1UaC+TDM/CPj0tsyBnid2y1TGJ/ysgnXQlqSBn1yWPvSPpC3q81wSWUFCF
dftmACbUk8Qz2/++3O2+pRL3lF9VJv5RRPqkcbCi/YXrY6liURZsoJKGJYFi
MD+kX78oLukmhYYvOBxzWAiv7doAQc+2YDeGZ6Mv7k+o4kM42I1PB9OH+UVn
dOJxZPOuP8NaSWANGazc490IDIubOvaKU2MiOFi9DoJTjCQjRK8+ZZbfSxMA
/fjbmavjTGYZaQnRsx2Y986TO/8Dr/wajbTCH9UbhNU4aTvaqyEbkN93Ig8R
iqaXXfjoIbuzEBu3o0+jEIfky+c/XYhxdM06aIIPC2e6BLCo8VkRZui2Yzdk
nzvV+bs0nmvoRTvmsUFPyJ29R5Sm/LgpBoU0KnFU2cxDgxB04x0QTvttoSyJ
Il5lOl8St2q/KjUkDtCy9PcBg/txG7eZSph2Y0v77O1LXCHO+SH6Nb8rO3QY
DeMPaFn612Ej335QRsk2WV8ElhIj7c4benPMoLzF4lPDPgcsh6GWs/xZPmfG
yjb5s1jPi9UoXH1/yGL1lCzeY6KK4+HlosOYsKjwy517PsdDxWQ+GEOtGRFS
eUJL0Oi/NgfhKTW+7X0bs0lS3PshWRTAYzTSKHv3D//EchC30AeXjY7ohDIM
5Jw+YJMmECTl542AVD8hiaFA/jMBnRstEor4gd5oQQIBvxWDmdRrcxVzRHKj
FHoiJhWo9sYb3H2m8n9+vB39iqXNqqwqXj6cIHrdrt0tliwlsSnCPhuaat1/
cL4emeHrEnD6rAoLMOEEPQWTGwuGM5OnGZBH5GcvLVtBRpjrI4a/ph5MO7B/
mAC88OeJkFqq/30DMm4oa4oTaQiZIG9ixMwFPEzmmXYa7SEYgO21DF8kH+Jg
kO78LXFWMRPv+bmEqliKfRikLij4oK9M2HouwlaHEiaATYa+sHSM352xCAlC
GwCxJw/51wD7QBFf72TKkW39/cQy3SQP0z+nKjjApTQjHZgEyM8Q0A+KUEQV
GN1EU8hrTkHhasOWKJqFkSWjs/Izotc0r5jzsFnkD1sXhrVBvDdhKpbL317B
PLKWAqgCDkTMgH93BJMhw7HpPRy4vwuSLejHoIx5pMvu0AhGN3tQVNzHmzcG
eFiaGSDxAYdkwX0ytTFsUY/kithOW41kCvNnK7p5bWs5ZN2895eLkr+LviVF
YG9zhcibF4g5d8vikt5wHPmSlCYLrhckEFEv36pq5Y5y4aavgCnCgfXDC42h
ZCg/Cqc0wITdeA2kxLJd2UzogiaxkHDe2xj/ncPAHyEGnWqHJafRdmmIJZDa
dd+Y6WL26qUlwk7N2RJndDY9sbsX831u1KxC6Rb0NIBL4vS6hGajAL2w/ogm
LcnRMdGrT6NQTwT7RZoegf2cg/h1W+1xPbuZtKFlln9TFbNUzyTEmJhYMWP9
z141/FH7aHhox8cI0pOhnUMjl9Nb1KzvYakZbmzOFnJYShC/ZKyLrTnNR6VW
X+hemwlt94sU3TELQM7YanhsZlM64vEBQGmmRaE8jnQR0pRXJMBBj4inQ+py
8ZS/nBiFNQoRwd8DQBGD21lxoisE+CAb8Lo7iyQy4eaUCmShZvM/8uzbqgLZ
iG4y8TTXHmEBhkxG+xxA8sqPkc1t7NTTnHR469K3LrHt0LlXU/wqXgYizokU
jir3Q3RdJkJ4HRh2+qi0b/kU1n79f9/2/kU3TxaAQJAQGXYn+8NTrC/+yJiJ
68i4bWeQMml7QrQkJhbkCc0jJdqD0j04MVqYo97ff4Pe+jUVhp2PPjAGokbe
RAA3zq24wJI9QIhwojDdWCq4ZWCwYR52xnZDov2k/yOuzZ5Cl0o4O8aazDux
HuxUL91nFyESR3IjhVNj/az9LWkW4sFqdSu7BhE/vNJRw2+ApgYIjX/bv2vq
gEktVqGXVHapd3BADY+uefzhZsT8bKataBlLZdNzjRmbJKBRmlLxLtPuzU0g
//Do9knKU2Cezs+SZEbNsPXnWHjeefwUV4dZXCU48aPmkLVJCi31DutLk4p+
A6AXR/1mhBTRZm3iXu+MvkQBrl+3NYS5MjEstD1hsAKL96DIkAWcSFvZh7RQ
3s6MyubY3/ZRHJAMNzaEDpP5Pki8MzB9kshXB91vWE8Mtqxg+3MKz7rqqlRz
/byJh9YOurtm2vmAyOdo48w2peQItLduEyTwb+k1fOsMggSZ0GIfIescbIW/
Jt2UNYDpISFhNGLarSZjH9QlfJNnrm2ENxEnmCEzLOhz9OAdcCxo+L6LPMTY
TWHxbR6Qx1VVhjTMDm9bHp9+LiAATcq1gxQyWTT1Pj6RUG0dwX47N6MtCmv1
eeBHLGAtpabo+vadDp26wsB5p7d12jwlLFZ3u5a+wAa0amQ5zMEw/U2g9ZP7
1sYqqPLDDjgr155HNKa/hdXY1yOaeWDKS7FBuim1AvdmqVl1fgDu67aeTk5O
BgXfHilcM3uZnB2zmsCouLM0KckMhc8COgOZc84dLYqy6vzpcr+92BXfyOEw
T/n/exj90z2opjuyambIKOLOY7XB5wEQT64wjWp1z6QriYu0n9vs4UjKvkKh
WgXnSBzMnd4NOv+x4WLCXsWQFi1E2TPtvrXJq/eWd6BWOF4fnYKPFvGiEdLV
6oQHjiZuwRooOLYNdXIsuuJltvbFeFB4ku7QFFQWie75zdlRFZd/TOOTRYXU
suaaPfDYTCJ3YbQAyAcg1T0RgchrgDhncvvrrveSA7hh4iYufHotkm02EERR
kQIVcsA4btUIOiTuRNHZuBJ5SCJL89c80N/iF10219UaQfMt2ispkURbCCrF
xRLp1BYD8pXEMFhvMTH3GmMSfsloN3/YOc3Z3Goi+zi2wCs2+H2AhSjK1Mdk
zE8POT59jKOgywkMW2Sa0nAr+GctywRgerWh5oJvPB4HgXnmj5L8aWMf3wxC
IyHFaioRYfGjFL+exOmNeazDP2x2aUKzY3niNgod/0VgtHckalz7/4XBiqAi
cWXxVgog/krhUW7qmwt0256thLFliXu1NgGg8j8QpXBLWJFITE3kWulRvnw4
SDsdp/iSRyprPvuaheDWwj9XN2WWWDZC5nb1tDo/L/gkYKyuTx7kt9h1VGLC
6myywEwh0Yk54MAD8FH2P818zeySPqBRWD23IMDamXsm5z9Bj2rIzMczkZ0r
dVFoXyY52AU0uMTJBohKztqGLwJT05fLu0lHpUxrV4c2WxLDkQZu4faFNxWU
jZzi/dDRU+KNjN6pnFS4Lfzb+puDUV6MQ9PAlI4HMbMAb55Q1Hv5k8nnkLZY
ELLtbXvMHvfUuJiRiVmMb828JKQegZNQG4Eg6O4xYQHWjYk3t+sfAF2/+cKv
XIuWAyk5bjj17pQkr6ogTOO74U9+ANHkoMoero5pH75tW6SykRzJtaZWB2MF
ZKFa2N7jdnVRa7wzLvysQdu5dc/LCTYg2EB2OwZNCvQqEop595PGMF9g32Pg
7GcNr0xhTSY5WDHcNCku01fDzYbPdwLnBKbL3R+yS0qEKz8pAqWusEKOqcQQ
YgZlGC/Y+xWdmgahSYuk0gHZunObnMga57TFWIvhab1CJO331peJkLUQCcMv
moF2v/yn5+nO/UGLM2h4xnGPdVHTSbDKAbPx79nOb0DpXzO9KMB4WdA96xsc
S7SCt9wv0K5eNuAMMH2OUP3aKqOylx5Y7nNH4qpSZ0KwjBHdwrgmwmtWY+oP
k1GXr7CGklmC0NJpMX+pmDoigMHkLD9pLNp2hvZsd9ehBTGG/opKTWx3oaZs
TXQ1XO1KTUSZlytq18SjyF2OGxDOHuhk5eBfDInylzkVHSGrXBM32Zv9iWF4
iR7WJABQd7T2BBJ9MuhxCufd+QoJwguitwKnmMb/uQO1nFEZMK4/ldHAGiHx
aEBMtOi96QVVOu5UDPp/+StjW+g5aZ7BWAID1r66DfPCQeuO22wkTKl+YKzU
S82cvC1QRDTzqeMdXG2X/VrnsdHrsCz04DQ0yU08XyBde65+fopL7zlwpE0k
meZagzCPyM6GscESRv5TFuXynsXa+fc6myTKTDOQBwY405eKidW30xQjOiku
KVQL2xqnGf58aeC5jcWTErcaXXj7KmPdzDxU8P7KD4Z4dz1ZFNJfeh8KVmib
ryrPT89OAHRwdaDLRQSNHv6oFkBK7K2jJd0UpQx3rCT5xP3dNexV3r9Tutx8
geFjFFEaFH8WlsSSlwZwbBjCrfanb0ix0BAE1c1cR3dNlSIjB6Xfmqyoke2m
89VpuG5ubhTvgaZLlJIawqbqKSVrRmCJsvZOgue++gE+Yl6y+YuzRrDqWolB
ysNKTUYYwOS1xM8IJOU3XdRuWh5xiIYef2cW/2v40Jzirmdpv6jytCqSGMsa
+OROqnELvgCDl7QUqObdY9elLG0JdPFUjXyyIiNvJcowVSq4h7PrNTEZJ++6
03qxexCZMmlTUZDovqWmdlhP+SfgF1tYdLeoL7A/7Ws1/cT2MNMySe/qhbNq
PehVUwoaqV1m5E/5W7jcVI0T5Jrfbe8wRoQNkEQsQiDsBYlt+Y97EHNLUaMU
rCgRzsexn1hhiP+G/Qq+hchv6R3s7T7I7Q6fdBt3nb2C6dDsFLfgMOPPcJSP
JtM5mt1Sze2Ky++pT5ghnXu9mJ0gpWYFpeWxcH+AoxrHrdzN6JnwTQrVNdBa
COPD5ouLrrFQ7P79zEc1Yvj2W6Tk3XPQ5OItswk5N8sw/y/mCVISPUdsSaTA
iIXt69WZX86SbnJUuNGBbFazxbeKxnmOl75Gk616e9sqXdwgD1eC+1o74cki
OZMMv+CBJnSruBiD6L6T/DADSZ/Qk43w1jQcwVCDxO8MuqPj+XUKNBMiYXYL
j2LpIUqYmclKm3tjuSP45I+ynkYde8g6UQxwzCzENaV2+LegjhJgHNTYFYTT
A5hTz3zsEziy2vHAfEzVUzR5JW0fjTKGevujY72XGTLkNk0zVVVDSg+0QoHq
kHEcV+HBELStObzmKEXz/GCENd4fkjzjjaG9qBA4Ji2nyMxu7I1d8SG+gyrh
DdS9v5bupGb0F0uqa2MEiLUzy4iQ4G05k9mVUgpZ7zLxChufJs8L2UgZDFSV
MFQb9RSLu8DiLvBJTC6sI5Uu7jnTuuV8d7OHoT23Ahef3qv+7I0343dmGXX0
GBqIA7SwxwvDS94QXAm1tLb6yWn449zHtA3tZB/8G0ShHYH7jdnykBXhB0xj
zkDs/mQx3kJrmZZPBaS/H/yLdtVIHjdpfCmMoHnU+r0VhbaNnmdBeEuASiNC
f6obNsTxNDNbbTkVGThL/EjvwwyV/1186706XT3bB/O8ZwVfEqBO7uHBh7MJ
QbnT/RMon4fxbnl4yTbwz/CT6XIQVYCVoQk8qTNriFW6v+6nLy96iNkk9mi6
nV721d7pXhrgyGpYKvj+EZPVR+YKuBv89eF1KincOqhaaTYNHbjzEaBIo8jO
2hqSJvTCwneVx5Zbgl1sWDb591OiUni25Fy6BimFhOcDcziJJZ64yOr4N2KV
G8ksRJkMwllsYK0pUMZL7MCu7FTcfRico2o/EP3IO0a/IevE7PKjSSAHjp7Z
b83PHuhAtVrNJoKemImZ28yqeeU1nupaKW5ij2Xt6xHyA5FWMmKyfGq76tI7
frc4enmaqiZpDQtG5bQFFm/O5Tu24Pi0c2QmkKDpiJqcoOE5AvpIH0mxw54Q
l6erxWXwv7Ez+rcrTQDT87KYLqdDfy1NiltXMLv4ZKeR09zVYLlASrZmD9fX
xnnATpr0vEEtCK2sbpOz1l0KjPlFKPFsEvcxUwHFII0d1YH2Z+keysJoM9hS
gXKSRM9f1Hz/N1p29IUnqKIipfYIlTgnTYOSzR0e8uX4EqtWB1pB53OyXSzd
u906GbLjJVKiZhROcqZbfNPeHvAX5ri0u3rgT8pViLcM8kgoTu0c7FD7LMDx
TeFDLL482Fl7chNhauSSBTxQPsUwUrqasAfR5bwfQuKHzXE/BY1yIdEFJF/c
lHTUg2i3g9LWbgkPgZqMouVZIecuPZtg73HzqakU4Qs/uirO7Ix628hW21QF
hh0EDrn8Jq6pyeNELTw3UAg42+/HWvbswZc7XjxrAwNfYw4tSMYzZWm07RJP
0pj3mbiDyE+Shzqabd/pv+bX3NGIVFJEBpnFqVROavXx+ZFfryQMsgYmeD6Y
O/HPNpXsg0NemLvzqZVNtKEmvkYMlQ5KhWBXYQzwcRpNVPgnWUOovzafKQ26
PL4rRLiUUFJh9V+SUeF6Mw3rxgyaUzC6/Flbwp4Y1UaynDCv5gK7nGRCnJEJ
6n7aO1tnxRmaAO64AQMaXj735nKTsGwReM/neVnLRlPpnZDzqaik7D9DYTwG
sj54cAPfQDhVmVZhyZcSn9Fo3XffQ0C9LK2n3Ts4xHg6Us6+YedTTr7R3PHZ
/QuVOJwjITMC47Mj2YzDF0DHP/2evmTVW2eahgODsAoFb8TrSt6fgqw0FGMH
JmlIT1he+Dk9iNpdUpuIEOYvWiQbSnv9vC4R0umTSxamQfurIOnIRUNmgs6d
8WjG4q7ADWcSSISbEFQWS0DEr8nNL82fzbzEr0jJxM5z/LMfHTsoSV116QGq
gc7C/ei41lq4wLMWgsL3HxjDPkyPgGAeGlS8SkK8SiVg6SRBeUDLsWip0gW4
CpyMqUGpui/WHYdoxs6w4G9mc/+4XBaZV8WOu8vCzu43fmd1vUsFxnZh71bP
a9hc4KEyddzZ2zzkH6Xe00qbIfESBbEkCe3JhVBmovo4NKfsjNk1o0NL+bJz
BrDZ6Wf2zR2J+80twUloml+LmgcCLxu0toyJeK9aveixc/2tMNmzyBaWWEL3
6gYnaxUeFTMqiIqIKrCPrzjDLS+JgSBHL29HH4ke2lAh6pfizFgcGeZGb6yH
lPFYwusNNisvbruOLiEgeGKl8NCYIJomYEaiJT5cAD4rPGVCExAlQzq1K4HW
QzWgcKlG2n5UlzVuz6gNOE8mSbB2vHpS2t74kAAysxPNz4umpDuPWtw1iKnW
79lrvY2huWo9NtDtUU5ZxeAypnElLVWZ3/YKfEWv/V6NCEF459FnD4ChKniJ
mZ0HA7bMOSj5tIFbHjHvuhFTogVWf7Rkq+fNANf2PNlL3odZNN3ofSCzYeXO
CTR4Q+yVasMHLvbC+QvrsUnXU31GUWirP/UEtmOqgn2gP3xleEYYrCCXpGRy
PKT+G7GobmO0VbyscWI+UoULatWppPnywws+SfJawI4+v6qhORnTRXylZsRK
6uFUt9Z/BlzQgJSOZD2qKBdCOFhws/aE5TtwlCA8zdALupOS1bbHkJlowjpW
nTaxd8dk6+XxbsKk9OpKM7boPOxzNwXn842QmYzmvxp9/mY/ifS91ZXz4AST
SAksU4UMjzjkhTUYeMa8rYzTiw2QtizQqxL8BIvr3uFNhAgGXXYPt5Zpe+R2
q5FBtCGAJqZpulm5/zM1Aa+CQtZ6J67v0BnPU9r0JZrCB8PjnWFz/53CaUix
+UJvHXqYwVXtlcQCnINLHUpc5jIMCFPOXiz8aSK8a+4aOEuGRH3usIAotYKU
xr1zsdNNYGJ7yxn21+76V2nVUc1VwrG2M1faKIL7lkZgmLUD1KrcjyQYHWyx
PqsqXtWeVteUNFFVPYOdnRZKceyWz/y27q58HiL9lGxFTV9UUBuPk7QhSYC+
CVpr3YU6Z16FyjrE1AOuk0+lM0YtIHK4MG6DtJ+sYJvTKfXwv738Cj7xFqU4
RA6qxyrhgXi+4XmdyZVmxe0uWikuPx33EWko9TWIFD0IiZY9dAzjzIs1ensu
DBJ5xgoLykrOBSVewpsuWWAwAuU0DfVfI9vMzaCVoUTEoyPsXC+Qab8rdcC8
AZm3neJ2ES7Wll40fjy9/4kJzgSF/MzqsPOZAGaHPppGWkngbwZVO2qpb6DR
lsdWY5BNvmVTvj58bqSacqLF4MWojZ2rFafbm5Vn/PeyDmSCbaJ2IRKPyT1H
np5j2aD62/R1Nco68mxUJaacSWrraiEBIcpUWY/kMXB9yPJ44mXmGFXYHaVU
My6EbguyYhUqT9Hf1IFgfOhObIsf/nJRw/ZpLyTnF9N0uCxrdyFBOmFFYpGC
at6WliaWJcZUOuir8NCOyofAPOSivxoixT7i8cl6736zkwzUjbxBFOqex4Qp
nf2nSlnMkPH8+bDpOv0EN6EVFdBltwItNEKO8N1QQNonSK6MjT3d6wlAJpWl
y2Z5GtWLfKWlv9VSLE3KzSzqrxtYMtV2JBIoQSMPSla/u6x+l0eDiEMEJTPe
14MVCXJ+cfgXYLOL99VjrHn5Cjl/9yyKFoebma/CIQYmLKuIKu3mmOO15VSf
jlc/D3MSkg8YAGwptnHgleX/Ny4C/vH9Vvk63GoO0yZVpm+qjeEG4VBbN0f5
7OeAU6vNP8/23mb+XbBPefiu77DQX5SZvBGMrNzkwpg1NSWJmToTHtSNzcyo
dGStgXK7S0bsGn7VuQj0uh1jXTpoci2lcDVWLiaewR5Fhmu8rQd9kgvSdkx1
ZVOTYsJo3vo0+mMoPsO1lDf/TUG4ULx9U6uQNabCOzaDrJrq02UzlfP+cuUM
zzVEmlFa9res+DQcVYLNmPTdYWo0TZJpbiZFPi1wb/6KoJWwPlxRw6sDD//l
rsodb6dAqidYB+3C6L8pRb0zQNHR6ZC2DL6P2d04Zh4sGkswZqWl7kJkwE9s
boHXyP6NDRZAtiQx24eFH+noSIAFO0JGK3r9b7FZO8spuGUtTD0g1f3xknV+
hxuQjF+8Zu6EfEZG2j0ieZHo1LgBzU2AIJc2zCYZeULVBodqa5V3gX1gsRZS
pPN2xjH3wvZf/Jt3nAqAfdmCsJdIBDE9rVdq0/HFvheZpTdtnMscH6Fc9nH+
8cq2vwFOoKbCtHDegzTgj3rUpSsXrVIlHUm60Pz+npGBBIsFKLEX35FB4l9D
QkneSOEipm/ycD2C8AW1dt9vtAFxkBNijxi+v3bSKJ2CiEw1pf0vr/gm18uZ
ieCOtrA/+rZY5T2eSSVJL1P+C9THSXscZaj9z+Yk1DGfh+ufJS9ayeXuqhiA
bAuBbwVER9tQ85p1TAZebW0X4GgQnI0xoAQgB4T3YDgxnMyejzCOiYwGmeww
b1NLkFiSjz2B1JFs0JZHHplOqeXonDIlbZTt/5Wb4rqPTYrW+UcwflTyt1B5
w4tn6oYFxUYLKFevKPcwc2yXZAtQYZpqU0V4YbxaLaItqGMvVg+75wKZcTf/
tvj8S7X83g56izgzH4R5SSB02atzSQ50Qw228PpadT1+PwBuMcV8XknGzfwH
Iw1VcRJNLLqtZ5vnNpDnZaa9D9KAeMpoTz560eCN1CsVl4dorXc0E0ShBQ5d
VFrGSgly478taddX7alwmAIOK1S/qROT20c++aHP7GA6cUf0/HSWq/NWwpF0
RfPXtOctGjfwyX2HWZwfJCBzKNZQ9LLF66o3qBIhgcqDLZ4I4itU02qy5Uc3
IqIkDrDroyEghHOhDJXpYf9BGVjiP/AgUqqil2OUuE+3AjXl1hh6lLrK+yAS
aTwGHq+iP/NpZt4H7AgL8VkSJJPxqnhK0zVAAX3HMInvxU9a+24OwKVR6zsF
OCPYYXUg1I4RyvTA2CYsl/QDFAUmPtv5DK0kBgBbm/l9wH1YTgX2Tyv2A/ab
zLYF6VOdv9/lFIgOekhSBBn4pX71C1ByHNfp+eEfYCJqx8Bt+ebX2BvYqatz
oj+WYgRwBGbdVUWplzwAxpotP+W1GBhuFPpc+8bTDzed53/yt8EyXCf+7bRa
YqIxr0K8lF30BSuE3MStYzCwFnXoKSDJi5HHQukF2Rewc/KxdqU4WQsaWhiw
4w3Zx9tNDiPwAxi/oSTAy4w23lWYpumBipJX6z8a/5rzDytGwHy3NwkEEinW
LJF0YFYHVeOuUR0jd2WvRwOBWzRW3bk4GYOLVYR/JyZTCDVEoxShHR5GCnNz
GBhEN959ArHN4jNNWzt6fkgbK+HUbm3lzUGy+ooks5wALuv4PtSU++SAR/Pw
FXjal/zZAKsvzMFUzcrl+dcUVQ/flkvUQutcFFJTTKkCh7MD4xhXVCV2PQUW
S9NwBpTmJVi/80zgZxdJK3RTMLK49mLRAVI4+TlVtXKtkZ9eJ47u3I03qhHQ
QLTzPe6Bd69dYZUJ4pWp0Tj277IeXZBq4F38kIUp1pYFwZQrowLue5RaY4GP
+2QWkLKkqTivDvUx0CKfLMf2bUXzDWyIMJJPt685TgV9M38zSgBaROQUo1xW
qBVrwohv08fsDINhIwp4loSmNC3GTDFWlJutHAlm0ERPKPM9w1rQM9pf9nyP
FhBK0Kei4ysNJz9I268SYQfnK8czk+k89UOn6ZMf+7tDYYhoaz/bvY4EY+94
p0kvoY1Rwvj5ukCUJURE/mf5NMciXat4w1eCCxdb2+LsA9RQOFok/rUPYNQe
yriibXBd9GJCpCpuDdYP4M6qxfYAfJSiqLuCZuszYYIBKc4GKOINaMGEVIi+
LH5ul6A7ZetmmXC8gZJy5l5P9mht4FdLUiXbz1qDTqxaZ0VTUUTV3YuU03R5
BBaKpJYZsMH4Le8NetwnCrDYyyyHoI3MwUbvh85yWxCBIwpvqIoCCn3Sc1JB
0wnAYkXnyXpkjkBEZfskcD8j6eMnitDo7nXInAZdavIsfEpakEqyMHiMVei2
a3Ny/rYEpUzojsFLzNogdv3mGVzFrZgkZjxlnUUBArgZkdEvrSD8aQwEeaCd
gRXMP7fymjqafcOvPMF1/OVIOUQRnWdfyf8zcpZYRXXB6cCYYvetVzenL5gX
4VWtbUoWaeel8uU7aIRQP0oOdNwsYRtwfgjk7VeiUjzxcvEtWFHWFBfue9YW
G8oXWw2B+CFEunNTT4NIdfz4UbOgr+ka4zdVxXod/T3W7GYHvBG8qJCrTNU0
3pwuXIbvJ7blDYbNCTW9HARoums+rg4CpNiTrmIM5rOMgVDINHi/BfxS6iYh
Jf70cI1oKUpZZ6ipYyCJc33QYaT6JjkMfNaSQVXvmM/0QxZ26SseZ7HwduL5
ewTgIej1MidAQNz8A+ucYE2CXT4jiQBziEngbJV1WP9nmV8VPeTtY9FXCjWw
h8yjS+cCXPDeArU8FdQ6d6w5kYs95KGXSOObXEqzcwiQ8BipJkWHr7Wy4mgn
NP0GUeJfyTrX9J4h/JVbFm51G60H4QkwLXuoat5B1mmDZ1OMYiNlP2lGAi01
oOSb6e43kFVxZ2Viar7IDOL5x0Sq+g4pGXyoQH0q3/aQueQol2tiq1qenz23
xeTr730piios/ad2GUUjZv69TXJGG6P5Ndwg3cImNU7poT9YuvGekhv3KVYy
/Lq+fxSgUfUn6ykE3sCDnLvDtyuBZxQTR8qaK1YURdk9w8qmdYpJnUG3PD9b
m4AohtjA/4OU19AuS+x96xtmMfrtJZKzLOdd/3fWtjQNDgMd7tZAoPDo2K8y
+S8CqWmRC/Jer3TPiHaIl5HrrBMt67eWycBii9A/6AGKiXA1nyWBQ96lEwg7
56Vj1A1VvFbjx0qpxG9+10s1NzAHRxgbO16AUxaPy7SzHS/uuj5Lr7MK33Dz
dPjhorAlaX8jXRuHeUYVM5R+vlJOaHxgWAkm2C6Sn4MqaMpRm1F368jr4CrE
BIBthFHb/m4/VxZZY572gLYLjm7kElLqNJhkMhKyUnK1oaJUDDOoKcTPztu3
RyvoSS1/U14QENA4VLywOYyO8ltZGs3USwFJXyb5Wxm9hQfCzIGtL3JH/w52
us0aI2MhbTcST5XG7OGwUr4ZDmKdGJAKGkAzHGaeL+kxt4Ov+cYNYBgyDVFg
qOitTQQ6kj2ogALlVaKnXXNZcLv4ULf7IxRKs0U503Qfjwwl93jrzfpv6Vx2
GkBF5ALqlS95Q2fb6Z2QkaBmQUy9OAl6mkn9gv1Pn6wjIFkupUMyRMMlK7LW
KsB/EA3PGFZumRbqkR4peXdUbck9ICj4+w/BBw+S8j+O2U/UVBhhMZdSEaka
yNrCPXtEUEZSE1DdYOCLRjmFuHIsvP/GgqbGrE2HOpnIzZfoX6HRqVnWiqQg
bDoOOKIht5JuB7ZdajhfZ6V+dppviQF4cqsgVwwocVzy4BW/v3dpVTWm9kVe
iiqR/aKCKNj/afMdHnWhgNEgbrGj658mLR9V51u610FkaRUzbsEUy6ph6Tir
mWfRuEzx67Fd6elqIxLu9hcdIl08v1q8OHi0RpUSicnjojzGxng5H0LC9HeJ
nVNZ8hJia3oXjlbmvDBj7/zhfPHsQYNVVnR9mIyf+oAmzXAf6ksvbU+Jf9TR
U9DF2g2idzw/UjY2EM0STtiq7Nqgu2d8Jl5gyN5MrXHHC40j1wu4RNxUqqiN
1qbda8U0L1hkGiwDJ0/AoXD1ZD2/yxheMakwgdoRkiPagOVu55DbykwmjCOU
e0J+IxcUuJV8XArB6IDi3TjN4NpiIihhQUUYhxtJ0KULt/GrcvUxQxDYkyHz
eI+Xh3WQrFXTIxYYmnMhCfPCvtwkZAOerNVvj+5tGfk+kituX2IphHIK1U2c
wdAi924hMrD1Ud4+pj8vbeNjTPucBq9B4WsQGwkL7niLBL088hi79sWSDcNe
J0oIOiHysepee0tTjGDeIT9xrvCUfFcNHQrf3M+Tfy8fF0cSSAoO60643Xi4
9yVXjHtr3LZwkOHv2Cq9b+dbixkZU56ZLc8sFuMS21XShc9qiMZsRlDSKV1m
C/Zc/gVUuhE0Zc/VVU4kL7yfguwG/zJCYxPuVv18BV60ZJz7016aAf1QdElg
K9atWQqdWcxiYYinX1rPrt0Glvecccje6lsKrN+ZB0Jo1cMGyon4NEDpHD6t
i4ldqm4MUjHR9LkY5sZAixUIOJ+NKz6CixZyucg8pteKD3C4EOGnN+ep8/kd
NiRaUD59qZztDuVoPAzLEA4k6DzF8eLfcuNwWHwDsVacfqs8uCx4+4s/9iw3
pjCmlbqeyBjWQLz23d3Q5uATQiXPqNqfCj5+Qwq0eg2VOEkGNZAK/6FbC3kx
4+IokXqbxTXjAO2Gx8RHxv+CndP84ZjfsZaFXGxScjQao668QqqlqnFjKDlo
SWqzDyhjtgI29AUUS4kAQ9PmsPQJheRBosiHuxvL5WIAbE2LzunfXsE4rMU2
2fFMsUyDriEngOS9LPr9PbDpJbTo5/pfEibBB60ixLSwz0RmV8XetYIs76+K
uIubSj4YBkRa4QcKJFL/ActNJdm0+5USAqR3qlubUGtEKMhEBg9YEdTQ7Dh7
VN86gAvPqj2E98ZxlDwVVjsW4HZZE4/Z7hCHAxv8I7aFvidWW48+jNKa2dab
tu/uba/mND1VtH/t0bfgONv+IOZt3l92DOScfU82Lx2VJ4Haez6myAsRx8Xv
0Kg0iMII6vLXnlulJiVWyKK+NVmJdkZvMyv9wQtQAxQPDJjCc6d97hp3o0JD
3eEBbqxcj79al+3ZIyAH3SlZffHEireE+oSJbKsPuTGcG7FAeUQ/CVnx6hzI
FYLJCIjg3oORlyNpAQqVF12HvywzOJYiC1h3tM7DWKrcnX/zixf05f+BtOS1
8q7hwu1PLh8+ePPsbaaXZYlp93IOZPNTmkqfcsDTVnbTulqeb3tu8+a6FeFn
r2ofazPzuswkcHm+35NSdanz4/+FZl+ui3T/EvzUtc8sSBz1j9qaM5dqriv8
c74iubaxva9isSL6gtlTHMzTPPdbFcsamI60F5VZDc4adREncA8G9xjQwp8w
KspmMsjAn9bF8mHYEwv4e8ukkNuHkrVINtKuI2x3CsPO3ktV8zqO9juJEpG+
THYp6vK2nln0guYKisJxISrGVy7xHNMvAFqIYuHY037+NXpYI3cKeWH1ioDy
/Vjfz9UhtH9ZpM1ph2SuvJnM5/AajqFxWhTbt6kBXviFw4ocEpkFjS0wFZ1v
DzZSw0tudCZHiuSMO31xfaH564IfwfdGUuyN16mdM4urMrpJ0AKk3gIOaPu7
0tMmMj8O+yMpCRPRZIi61bjwv4vvIaxWFVooWKaFx6W2Tpzz9TKGLXFKvo8n
Oer/adZa3JSILRS7UP7S7T/G1G7oxaaA1Y0Cghq3mBbuI/5JgsbU37df/CKG
IV0VyokfKGMnMWdxA6abDVuj3ZQDtg3b70qA/76tqgJJdaFxi0sniFjF4Q6A
1UyjC8w6889uBVlgW6co6rYdwENT7Dd3in/D4U4198K6qDeQYbf0cPdJSg4R
NeI0yi8jtW3YUbN9LJtxm1NwFHTRvkaOD7kBHh0Qx9oCOd8tjcs3S5roBVBC
cIqmtkHntvl7TaSAv7qpMD/AKdwTC0S1sr0XIdMTEBSegMQVMTmYS/14lPIU
PYcoABfPQJVLDFX3tQIYcfn43DuWfOdH7GgHbuBgTV+2pCvDK+s0q0UTsJF4
0angugomXzFhe/mZuRxPmwLjYrGm97o3UPd2xyBxXNbCykcsp1fFbYAlyGyF
d705hLYh+dXq4m+rVIHF/lfpXDt/bbx09rteRyVy0LRm+DM2OHZzBLNA2ZEw
Kr1CTIstMNW9u79O4tVs2nM2A/XxwnkCuoBPKIlsaIUlApzZ93ZD4I2Pmjgv
HJGUdmx5rcCl4iUXvW0pQvOrHvRsesAD1etnWNUDcsTsTGlmhKjY4KFx4GVK
dW2MzHdVkQfMZkgsS0YvFckYgTNG0FLSkL+yUG2QxYRlpmpFA7qPqzGSYdtJ
jHOe6yL+63hInatr4aa66F7FT5DrxxB+lCkcfbhQ7EinWiDUUnVaN8ufbNPB
2XgsvhcBPhX1j7mRZ5NZWuCafdTvgJnfDUc9PnqKRk+wL1cXL9tl6/I/EWM5
f2b4Fd0e8hD9jVG87LI/Jaekzv8HDWY20Yrleq8zuL8pcCF813WyiiMsWTBv
8ZVUyWu9UBR+FoCsmp6SLZNEwUWDPBzJmXyaNB7LGZXyJaAIhgfSSVqdi6VI
vpEYMd3F9PQJx1tr7EHr8tXEfaRAGolAhFoBsq+ZXQB5DtyuA9wTFTvkTB3y
omqoq0dPwC6Qlv2JcJLVeDYTNFwWrH5E2v+ADuGTwYvM3B8PPMEHjPr41qEg
rn1UN7xCOm+cLLd3zb4rmuUdl9gtLMgPUKJ+afvAa0ykyR99kUTqYPRWR0+/
zyZFnpOoObogjZMY/RDMbgcSs/Oor918/KhS6s3dgp+6JYSCKtMGYV5U6byj
S/ShtKDBU3WTC/R/2PN6ZgaHqn5g8GCOItdboj+jgqgnBl+ud69aCo/y7IMn
Ah966yN1DmBEwp2iWPJQxgIFYnzS9a1AJW1Tum9hhDXa1tFYxWQJ3aKx3Xwn
CekYzj8r45+FVZcy+QRorrveTiRh8DpYDUPwSuCncSVSL8ewnPb4Fvnm7cz5
ew6VKD67Rr+IBLR4afpHtDwufjJlnV9ri8m7zJCE+gdTm1Z+hiLjGAqPuVOo
fMwh1pWPuFE7UaeBwMguVR5ZDL92k15nuPefs1f5xJ8y0ZGBauw2b4sbzqx7
9T6kNdx73029Cf6eVXXVw3cIUFxocOP5k4qkENnJGd6/Hd3Zh4eDFO4TOjwz
DcKrLLYR9IE4gisdrGI7IXdCjhPPQffZPJsJNmAfKvCqMSpq6CKYjnMuiKpf
YiVvU4WmuCA7XJnfpTkmTcFoNlD5/Hu74Bx+qCN67lD2e5eJp3wwyXfleKJl
sKIcKLTbs/m+cnJ0YEK2Nz7yYDkLGeaf43ZeqkPnibyo0BFyB+oJOarGgiyp
eOnJm00lhBzuDfpKlRKY5uFpV2AHFdnIVpETOyZixUcI7NMhrC5Fj/1iaEuz
Uu/RPputmyD39n2X9qoJ7kr+d7mDeKZjZPhd8zf8Ut7PLPs0DuACi9BnVHLA
iCLqjBMQmArgZjOKtjtzXRtOEXrc65PrVsopEMxblTL8DejRanafm17SJpw9
UZZ8kJ1sGk/NLdHkA8AzlGe4XquQ2b6DNgBHKeXREwWiBN2TpWQsSoZsjK2I
Ra1Wyty2e51+uWkdMfIXhNg2GUs8uWi+EDArUrhODsRJ1H6DBrW+VSGrdb3d
vSfgyMpMoP+2weHef7uEx3gAmnPH7lLzcTGSWKdUQMOZJeuRT77K6d5z0uh8
2f1FwKzaNf8T/4cePwgAMQAaKhnNFR4ovOl9l7O0B87VnZA2LmJoMMLfE7mV
t7inDl0FWKDj5mLDAmFjxtRLWz4ISH+1WO6/yV1hI9jWPPsXEgrmiC637rUW
kpMsZnN8IqiZ+IQoLT9tXN4UbxvgDGaCSHQToulx+dfosp2gRejXzgqCC+zf
cfJar8LjvpiAU/EYkLjTIqQWl1Lm7YlHQftCs1MImAnCfP4mDD6KVIAC+5bC
TLj+p0l21TsUkxfGBcg0gilqlin7qSjAG7/yKNqOquGMUFs4HLKvxx0Mq/D4
EjxlumJVXP7Z4m5yf7DYG+9sddwZ4C2FAqyR2kyG9orNJmdtwbTN5VK8+hi/
6qG45S4xhHnlvCZ9F1D8/buFMkEgg2h/iKGJYP7RyEyQ4WsxvgOkFURPbZVx
AwIttFlvocYQef24IuccmQBY2r/v98mAnnFQ/4VjaHC5s1Ery9T/041OqTrN
sQaS9QJqkO8f5L5gyAn87KB7zstL63ncU9M3ILYTqNoKiFAZuKTav954uO0M
G9cZgGCUKR/efDDChmVGDg4OP069IGGzD//ZsvWvr167S6xh34pC7MdW8MWc
FAeXNry7aj5osyDSqIkccZNG9oXVfT9YcGmQy5mdDsPDiKuGY3tOH8/1SuV7
AcaC5aGiqNYDyGIIhZY+HCN/p/0Bt2SkUo9Y+SU/BLpv97OFGtsFCd69+FMQ
bThmaG0rcrvzYdiFcloFnNnGc5sD4P6WvK+kXSg7HDr3nOPe/j0vAUgbu8At
nVGaYncGaYpeYJ5XT+TIPSjNUTrcDXzzYhjH+hOzeHUFgbabCQ1iCrkXFETw
JtwJrjuyQBgGu4TzzxRVemSQkFIhvSSySHXN7AcOMz2m9AX1YrTEwCZPm+Gt
rMfn+0h+3W8jFp0zqmUjJBbLeiKJP+zYl1AV7R2+DTlBGdSTe8m9YWRAvVVu
XAdNshV/6hpfP0RFFl+gRDioK3E8JWgAGneaRxFAG9wBWSzlXjn8s9/bQUKT
+eaMo8/ykcwz/Esq/WapI4bRC8Y+T3BYYb3PmQz+3MDk0DZCw+R2l25HvFeW
CCCfIyNYYKfqpc8t8v30Y8cr8aTGk//P/BKrpZ6qhgK+ojb3Bzus7aApklnw
XnbUtfrVpmKWApgSwi6mOoQdyv+PQChAqYKVrroj+YK1BRPv+KW/fgqAiPX1
OSncrF3IONjTq0WfSU8B56x79Pi7Z+FLG1+EwBp13JfjUaSVHn3TNStRWOVX
3brd42o/rO+osNH0Jjpde9S0vzNx3n2W+25wyMRdMN3wgWq5tF296Xsg6XXY
fkyyT+tLTuUBv/SDfFoE1JwPhcdFqL4Bk0zv55qaBC0dLanr79mGG97Bsd4V
d6utLTYq36/U/9Q463cg5ow2RupPdWFoYRszkLDypfjPwZHHwwGbwa5gVQ/U
VMXg5a2MUD+Rx1FqabK/3dXJLP0QxNMApJZlNG5wSiUuwmnsqrU4x7abvvTD
l7dYGkQ6/l1gh/mkj48OsqQil1xQ6Gozzc0C93h3wUSiFqNv0GYjww0Km1zf
A6WN7U0IKPU+iqRf4kS3Fgc9ouZVyNNQ/EWzewMJw6CDazq9AuwDygEipoFz
GgowGd73txOtSfbRCyz1/o4MZlZw4CF70AqItDKbwnvnBmOm/qu7xZ++M5/S
JjTXjobOcOGYWQ9y8lyrirXenwiJsgCAEltNFLtsnrM8+9X9ws19bVD4dzG0
LBRrqZf/vnEtwl2k1L3/C6lyiJHCGcINtJ/wWm+HXsIimIVqg4atJBoW9yoK
JGu64FsHgdiFu01HKGFz23HyGwpEA8gPwYAjSdoOEYHG86a10hdFPqOFJ9Br
lDSXNTWrov9IdDrtTOaHE2yXlyefQZE0sGNVSLTfXCbwTXjVFCyWpCTjE4AA
vAZK/ftJUCgBxFSWrpOnZ4upM1aYm/FSE0UUwzo7bjh7rpFdF3dWuj2jRLo/
wtBFzEU7La3dnlnePDqyXze3QnayjiNzVM5ureRRysjNQOSdBO/Ov5tmUHaa
0ZuuF3iKKLKhJ7AOiYYi0hNRJhGNCLpTNHuigUMGqXS4glhvFeaUJsenL93n
4FjyrFP9wY8nkVJW2237d6zeKertN5n5uXHE/qTuFVXf7k3e/O9sW0+9tJqV
/JMg29MWS3CSXmF//KeRRJFPCKBhT0UOl30LadmCyWzjOkclQZc4kR24XKz+
A7lS54xKafRk3942t4DBuk8pdWhMcj5uz4uhwlfQD7gyHW7GeYULNSXYjWpc
A98AWCKu567v+5wgr5Na/SthMD460iW+Y/31yPiM1mXzxWEvcvCWDUZAdcvt
jIqyMQjUHnyUbP34xn/2RQEEo9OsmrGpGJUr+xz7Vj46WWnroDhvi4e9RbiT
L5gf0q8pwK2vkBfBNZkHYC7Wrp3SGi9fd2x7XlBfqTRudagtWFEWP4nfcdJ6
6gH07JpWIb7LfF2Hp6AICs83JWc1+sbyLSgl/QenBs1+sa+TggN6XjKHGndz
7B4dUgA7tObQxqX/P7/+FZQVG++1aZ9sxfYDM4vl61pWjRAStP7PpGbZn1XD
0z3FFmX/AAFlyRgveeAkVc7wnq+AI5lm/XgBxWItFdR3FLtf2ZH1u+6FD9Th
uwT6+wXfItJPirg5N+nFSapx50Ru7FH2XzLCCZENuu4solrJkShw2cMF4r66
lQqLWjWFDerP1VHlsFnztXYt1Cvqy8Cmk9XD13dtfrrvjSmdF6U99OI79TZV
xfNuL77lFen/PSslTfJE2ntmXxqniTuAmWpW/xHSJ1dSIHVkY3cXrpfkE0Gx
GhIIVMw8BqvSy1gOi+xe3n6QfCJ+igIA8FvlSSB5t2uZPvjjU8IN7R/WnQjk
bNFkhqJY4mric+iR5CZ+siMiR3EQvqcSbpN3Yd/gDRLTK8NX9Kg6ZYGwIJvi
HVQWYGk5nDr6OWgWJdCz4GBlQ813xjAr+DWWemexQmxj1wISuryxjC2IHFlt
CXO1yFmQE7vXwlwi6u+Jd1RWYsk1tYknfmpJ6O88SisTmRqjo/kyYwCw0KAd
MlIlWWtJwvy2Gu29KZ53qpL59p+Uk8oqYz6ALu8Fa/H9MqEin5GhWyDDMRNR
4HwrT7IAU+WhW0PXsWzRNTZ3eoyyMKpe6Xe/lOlSHyjR8NHN9w5+Si1gCNg7
mPzBADiqItbSW4N14NCx60zGEKgfmzDZFdxxuMEILm63Tfc4MPwQxNcG0hCV
329wDPD+GbiT11r2Af7rsWIhYd8rjJ/d2hy+31I6NmMu0E9QLoztR3C4AG78
9Zh7WhCqCH4oNkgwG8+VjVzqsixB69X3JHCcq7IZ4VR2YG6I5QzD8/wbUVgp
LvHCddUb10SqnZF05FifQ8Le7OgHTzkjimFFdBqEae4V2dmKSe5fYZ0rF1ZZ
aEa2TO7m+pvunU3gl/EBWcu5zlSja23L0IZHSxjIXhwmNKZAj7hfuLxWF5A0
ujuZzGmpYl5TIDMpkcYBHT7mN0pVZ+klbhoVWvWb6XEA49OrVGZ8dyCiGB3l
KPADsBr5yeLxPVE8m2t9GDkZGiwsIXeCyrhzhu6rq+fzDophd7aSMp03+dn/
ptSOJVVCCosgYKkBT5AchcXUxovhGvqzZP+K7WSc3R2Nxgk5XKl27dMJ/F+G
n/InYkyhF5UtOVrBgisrO9R0agIhwH3IUgHIZQbt8AoO4Cq+q3+ISXtw28vz
VI/ReScs2MQYa9FHgvMuayQm9aWWrY+5k4T98wTUYNB2e4a2Kf5I8mTFuksA
3XX2Te2FoJE51ZJF4UXdUARuSvumbGXwymJlr3xiz07STziYAqKTqf5a5/Tv
PVBX3jy7b0bE4UNsL9fE1HI8HMSQlsESLIU92JRfTpzzEBhocOMMCUzCmpao
g5LrEIfxbBdQ8Ny0L6Ho4JLcKvR63pzjc+P68QlXw8Agoh7pAMPv0Ge2ex1e
Dfcz4CZRPUoKixin099wAaLviQ7Mpi1JkxNQPNEZzI2S4T2aso6Lbzph84MV
SNj0rVosPQNRznOeRKEPj+/V8sNYb97Mj2Ng+fRI/R0ZCio49dhB/x2YRJlA
vU+IPISpXoUZNKFjRKbTYnCeDb/cQIgLy3NmaJ1ouj68KbtFg97ypdGxpx/Z
2Waft1pxcUj8BRQHe1iejvKFMWeQXjt9CzBjac/GMvXLJDjylj0uDXYsd3Vz
lWV0aEWFIQ+oChfdfPZbdHzzajUHTbuwGgJQgMMZ3Z+0lVuYomCiuW+c9tG8
J1hLkJ3Bj1oMtfaMso5gBezHXSneaDhkaIzI7X+fDkoJ6Zw07LAJbbznBMe4
Kneq32FTDvccqc4lvuluKnT11QKpk2Ap42e9iXuj1d0fbDs8PKcFClaQWs9u
KvpScOOMQFyoGm2dCLN/RlXQ8YCDHaxnTrViDphTvwtRx6Y8ZIHOcso59RO5
B7uClZCwCJDesbQnkW8+YFBtW5319duykPgS4xXPpysNv15OsvduaBKyj4Jm
GNpXDyE7lKtICZrgbFpqzNzZQgHEmvHYl9ls1EU5Kxf8TV4q4MGrXxh+uhoU
rQZCqHuTqkPc5pj0MRTM9VC3ifLmj1fAznHbdQMAagtwb+KxWuDx6bNe8kkw
KPVL3deY2OFIIUliFSBaOX44cBZpuDF25FPDg4bskK7nmH9MmN3Lt0yNxX8z
VLTO5FGx/uL6c/kaDDLGjk24/PFMQ6dxcKjRS/yFyQoxQHV5Gf2l2Fyhj6Av
jVvsJQGuottlj2p7rr5jcpuCNpsTaHyDE0Eh2bNWL2+VDzJAo4af0XXWdvwZ
1t0p4AKVJ6c6ZvaoYzqqry8fpWAD3Pr4sySPyQ2RbkGmjgxTxcPX0Hx308lG
RCTjJG6U0eMovCyrbM/aqFLu7bsxXKLouEsaFIovYZEp93+oNzZlrE5On2Yw
XDPPgilyCGp5mF0Dy405VJsnvMzoayw2SjvjBlL9JkmD2DDSTYyZ6qFOxDDa
cFvcKeA/xbIuMwhb82a2kklu9/iWXKQUiw6SUTg5oRx4Qt0HZb3/t7kxfDA/
OXwsJoVn2PUrP4A2rvNLlxAAn0Ydr5GbmAcXCdEszGV3+BuwPhgdlq2iLGt6
bWoDk37zpg6SNFiSB+ZoqVJ3cq1Gn9mCsGdHVLsmyv1v36im9UCTR+K2kFkP
dxNdq98qVzboCDsf+jv3qTdokcKfHZw7CEgZo32U4zguThgVMRv25bIAG8zE
eLoNTndxvl53v+z82Zbr/A1qpoNJg+fhFIMaxmo5YYRhmyWHzst9Y2RumIID
WzfS9y2qqUedTNU/SLXhdltJCZtvNz3ZlocGYd0sFg8bS90vVXOfjcObahBP
IooZHq335oslDZ0zDSBxyh49ssTzuwVon9BXihKfXvt89gvCfwfT2bQZGo86
cJnLK8YX43x11q7O7LjMW+nZCwBOf7Wz/vyYsyq6eJfQ67M/iSYLflmeFlL0
xOVezEmYouS8/WfurId9/2JoAefqvzfhB4JonTGB0S5+iO0AZ8RR6OWaCStT
JPTR+MwwOMX+LMaHp+AvYF6pzuC9YZtNkCiCSGGh03ATveMyzLo9ZOcRtcwJ
rfiz+WKaFFZ7ZQNcI7rksKybHfemQkAPgEX8QPUmM3rqR9Jzh9IyiYyx4/RB
cE8SSb684Cl5WvD8hjBtkB30c4x8P4FpKIe/A7II1RgmBAYFEAGjz7WPrGWW
TF+rhLeMUMezXQLKe8QUtnMJvOOUmFbft4hppXjM9F74zZVidOJUWl4fXlwN
r26eN2yd0PLJ7R+GGgRcMBJRXXwjp+2cZOPO5MZ+hd6iP3u8zdIrOU7XqnZM
+9zoFGw58/MrDvgNcCKw5sA39L6pCs4pRk8KkpUHtLi1Wobm4j9daqYc4s6n
R4vzjDMmKU1hb0Scj0P8k3OXyMWCFGPDsMYoFX3NS1AyDlTINetFe/6Dml1v
Wh9DCp237iZtgTtv5Ptq0799MyBD5teWvYwgAc8TB0n+VE+VibVP0IrnZcWE
kMSECqO79ZYWg/PFmg+mweRPSORBjvojG7jHWE7Sm6D9ZyUhEiROMC3QyNyl
m8rQF6RhACnHOFR1AmThYnUssbsMRuAPlqwRglsbboENPQ9vTAArtgqw9gxO
U0tSGeyqDQrl0oYyaTq6ZH1x92AJjaaRsNsajuP6iOAZPOFPV09P4CnH/CDj
9VskQgZZ7dzNKATtFTDMuKP/E13T+SChV48mlshqIS+baE44XoOI8wpLBrQi
rn/uVYcZzbXsPgvUD4olorv8EqzIdaAdSAI3AO5Om+qe3xzUOXO8Mpi6PwiU
BEDMmubXEddCbfELG3DvEvUA3yidlSISq4ulZWpDHSlKLhYg1b38H/UTYD+d
RZtUV5tE/XpOYF0D+kkLD/oVs9Cw4uA3ImCFdYeJ7NRTMoUlrKoUu4xsV6Dl
RrnXXh0y331ITKXAeTLswWCajOTJb+px63CQk96/cQoDrV0V389IInRRed2d
8lAYRROWnriGk02ot+athso3C/pgmLkCpqk5fUAlF1RCjGY0IXm6KLjT9Caj
RJRrwmRKvVzV/WtQ0OSiwzz6o1++5VICydyVQpe06SX9o0kYp4dal13S3NBr
Z3rpGqG5b23zPSl19kmCQ/BkN642MQOd9dW9ZSinY92befuACzh391QBg3Ca
1vBaF3AaAV6jqcFYKZH9IMtidV7Rd+AZv8K9BiZoiv7k2g9XS0CcPFYSZfUg
LIN1OJCu1GghO5QH0/qMxBNUnFvQTJEFQ1Xkjfk1T7rKe8MSdDXwuxKPe+nd
zNJE2YMqplu0f4PvaCzIgSPUFUKaALmAP4ExoYcj9Cb8zefBcBrFHevBZvW8
sKrOrztMUnlijnDtkFUjML+IhA/mJBHF5f+8iaoFxBHvgS3OVnoeXj3jD8IO
LtasITG5w4Hcofu+La1pJod/l60gQjr1Eg9ZLhBC6mTyOoHD2R/x1JbGoGa1
tPNxMk0+hKyul3+ah59HnaVQzVH5eXJJ3ViNZpaQcVh/Nh3RlF3Sq88nawA8
tcOQTs/lBHMr5L9u+ZP7xwnfm0gZKFxSXIwMqr2KAATOUYY2y4jCby1h1va+
yelvLHcwoblyK3PngO/fVVQrFWpekRRYCbwEroV5p2MRSCJceK+30MD9kHzf
rEwLChkcHTh9+aj2mKwpstOcdOmhUJC7K9gm15oMxytacU3asTbRWodFBIBq
INlR0I9FOowpn0kejfK0LbkQZVYakuAYw+Yz6tf0TQdonxv8VMX9kkJWHqLi
KSX040lA8K5wzcV7x2v4L77EMBlSyxS/sGDBsrZ7sA8e8tNy6a1s4iZ1uWog
hVCBkQGNCFhahYrBrHxruIx6RdG2GQ5/MPACPU1+M7LgbNnhdHkdrvWMD4wP
YZWzS8rhKIPKlBHubbIxpUR0IgI9ARMLj2uM0Iwjc+eyS86bGjDXJhn8yWFn
nainjO2RD8RorkuZJebs7fdon8upzM64dY4if6rb6fAcUpG8ZycjT8X3Ah3l
L/yiWX9e61z8ZfqTqG+aXlreVQDByTsOIUR9yx6SuUa3qSU/eIphFPRHKCkM
JPRCCrcrEsubHzjUKP2nIb0x5vR7ihjoAVhhBUDo5qlXAcfOkpMXu/CZ5wdP
No78OTm38KG4KThFajL7spv1vf2C+POFlhWohLFu7Bv0VKZX2qZaYVOjcpg7
MI8moFPPdvBaDKTBG0SY/s78+P/2J0rZCqKcsNwcGZzrseVn4B5lsMD/UMnH
rnrmL5BVeonBfjeD5hxzulEK+RQszR3JY6b/B1wbf7rton3EJR5939jYrV8e
2V5y9OVpMCXzKRifNEP1FkGoQNJLvRoJCCw5TWMKdXQGEimTKhC4QUZ0roUr
4idj/8y1XmatF60mUV8Nmxn1/+fzIDClthIrQZl/UkE4DRYb/acwMlImJ31P
ZhaXEdtmgpdy/flbMLuwU56PR+08TY9iLef2uaFdqjeRzbDZ5riQuWHUASGM
tE3uow/bnoGQA/NVAvq1z8WAoaGm1Kc01Y3fxakfU8ooQH7E82Mhy3SXzeeH
qEMqfFtOykwNDtVHOvlzug8E7u5yhyUQb+A91SitGcMOXi4tXh8z6U/AOMBs
S0NB+FZEgCbuhyXwLfWHsUlEE6+AmKvLULCI2pcwUaDwf2g4U4/bTqDGrhao
oZ/xbW7PEf9XJExr8RNQRc6sZqa4TKan5rnIbOAMmhKAn2HFtMvYz5VQpX6P
dSFQtSLO1Wgp3r6Qum1SMi2CQetyK81TkCOg0NzYUDyWqveT8Dmph7qYjvZ7
DEqkVw7sz+8onxrD23FipwXXAxqUM4P/xU82AFEzlY4sXef8p4KZpWAFoRn5
yIayyckdxaNArtHnbEt1VsedzXUq/NHzd5Id2c5lRDH4n9YGlheaMX2XgHOR
Y01NqC0CPYLcKuuT49BQ1mSxEvkSlTxlYesEBEXS85Kz1LuzobanqBzEz0G8
W4DRoEyFpu/ku9vFNsmdWwm9C4EKVz4QL2Koxc9xgdSjQ0fwMOi208kW6jIX
KqrlG9bEl/K79sXrQ8CYtXQHbzHSDAAyMAguTZoKY4Auv/rlSwk51PhO9Is4
o7ysoSCBdkQmPiFOVg6bonmFA3euvQo7KKQK0yTJX/I9VL9lD+guxtIVTnMY
3HqeiJoysHYZg+1FTkZJkL+PUApEa942v5x7VbPDrFnXvLG+D/uOYr0R/c55
D0iqVkswFBwMT9Wy+eMOMHiJJ3IdZ8g+WbqlY2Wuj90WOu0rO7DV5TVYlWbm
Ir3FxQVYbjJqV5xgw0VVlQt6QnA+R1GSGLRtSLCBBHvHk+ewphgP0ZTZGywD
S2peUA+yPINONPErZ5hGfvPZELvBFpn1XtFS6eFJjXUMUM/JBfEOlQBjV6l+
AJgZZBeog0TViWYm9mFFN/v2vB8X9utN612a8P1EZ2EGNqaii1kt3vOENvUv
IUZvw9e/jMq9Vnt7bpud29lDiGmZMzBBaYdJk/4GYT6om2hlTWHe5l+n096l
/0gWCb0fS0599UfdPwloftDexuHbn3lULH2V3QRltNhnwy9qMqIMp6WS1ZfM
YYvpClywrUhF25BUww4cVD7zBptCdBXo6gkEjdRJnP9cOHfR7EkDYz76DK0i
k4N3MG1xZj2E/kfF4Q14V16OqAHT4HVjG723AhgRCuPxotRCVUtfTg8V1p2y
FQnHmuoXK3gFNv19zk+OAvgCyx6DFIUciV8qHsMoOqWcuAmcnSqLRXwL7ovl
Qf7LdeGvxwr22CGN/IXwlWH3byn5vCFFgxEoBnN2BAUST2ClBs+k+7HTFehW
dvLCIhoFitQbn9XjN2XzsyXb6tOfyvAsPVr6GWM4R+LbI/8XMnAVfmyam3DH
Cl/gww17WTrahHlyW1iCTGi58sbHM9i3UW/R5drOh/RQDq5pQ87Czh+B4Bul
KmrmNLqeX9ZEZ2Ac8M43qPr1TDOAJY4AmrPHG67/Pt1VFmYrCsp2XPXpOZl0
p/VDbujIgQp5crabABBGyKYhcfwa9AU07qXNu1sWPmPqgv1IQ7ks2Us56Sg5
4yFOAOGo8KbIHznX04+xh1KO8Jxp4dzmE0xJX2h3Rn9sktn68xcRiinxLLbn
c99ghuntuIj02e9rKs4ezD21W7iLqCrc8Z9EfZI9FftbIE5BeHD3hkl+HUct
tH9spfWYL67DUcRSeRGL/mCaeQJxT+o0vEqfuHB9/FH3tEduNEMyUxTJ52S7
gsnCvtoX9RqaExV6b1nIeLpUe2WGdDdQccS/f3/rtd0be4feGwG/FgsHTrPF
Dj7kxJrEYE8zJAUTNeQ8iZz8tguB5kR1LIA5A8OJcM+QQbre3KA/XJ7aF8cB
8ruoT/KNvx0RRuobBddqa1hc4YnSdkTacJ1juhwA0/sO3LSHkGGq6dJ7yVLP
VTV2Q+2xaaGm+DU/ondPORJpPQ1tgu2jeug4cWc5nLDokAakeSrWn879ECHC
kOc5xlMSbT47v7rY0kzAuU9erXLcp3trobmHvB0kg1whJyfbmRESqhLBRclW
exEIPXkeVvI6QCIrYWMjIjPnRdHUfFGLigl2QG1nsPfWc8XTLAOYsYXQaQ3e
FLJsFkfosfe42PYCaISySBm+oVHbguXXcoRWaPyuSH/QQ3sLH0p92CAUy5rS
qD9DqFWFNKdhoOU8rC2p6thID6i6ScwntQgByRT52hkO6Fq0UeBClU0aMJNW
R+wdj1UjztNAYmmRZ9OxgkpTheTUkO77j/ErKhSKp/sffPUxg256CgpI2K1w
KpabqznSWEWCyDcPbIxJ5jZLs9/ZuRBiiqcfFfGRhDB7ANedg6XIu1CWeRAh
iG68CIp/G9nmuVJNVxWSIAEJfSbNFFQT8Rw3eLIyQ2K6dDLDuRLKaaoyJ6Th
nW5pDUULIMCKTun2YbX39xaVSKlhrbLcwdicZmW8QwhRc2GtxlXMKaJtXX1Y
CLT+DY1IBP6ApUzXzniMne4lhfTzJz6Gr6iQHNNb9XNJGsZnRMyUkI2VF19J
Er8Lt2JicJdaFc8hKtRH/GvxncdpK8c+oc3caYSU/S0bJbBpUQuKlU3/5Oj1
w4x2S7xyIGoFQtG6qCMSZwET4wEQp2o+ixS+ICuDkYSX+GRPvzeKBAEVOhfb
w0u1GbMwTTA+1FFeC/5JysA0LIQg6yC9TbnK3kp0pYa6eyq5PVvcLaD/Mgir
LLDHtBiSYl/Tz++LkyNbCuMlXp6p5fAuxESZ84pxCU8b+hu5g9mQLol/Uvh2
0s+OMahEygTpozfyFL63/nwteDS9UNjPalbttjXX+2b95up+y8i0GqlgGlIr
RJmyh+xGQqXc+BBcZk6Oqtr1BNqZwj9hQTV1II/Ro4MAqAKZDwdRtwhcbMkS
TUnZB9fx0DN9WjL+VUtnOBxNlPVZ4lj4BaF9O8FyM4um/VNyhk/rJ9JxueQ0
datzJ8LzeLLmfC90wT2qCc2eUGfM3NwL+9Brn2HgcXUhMd8rBp7XXdlST22k
YCpbhm8cww7iNhJNJ0BFN94TH9lTnQUsQlRNgaptXp/1qx6dA/d4Vg7estd+
73VoTWMuKAYU9I0Htw2AnxN1WDqbxK+HDTNC3E+b7WM54jaULOB64ehnKTeU
xKc9q59j3nIenyUBW7PbfNhCs/bzjkS3va0BsuN6AQW5NnciInN6ztYlPWvu
lwPzC1Yj7BDWreoMYwLbaiJ6sgoon3a+qArVXtynF6ycgPypq39z1Ec+oMK3
1lLiAx8izHx4YpBO9azfVRcJ7rdYw53q/PC3aBgJARA06W8etaAiEyxoLD4q
/Md1rRlqGrrFj0j477MxVPkP08dpSkTVH4ap7oDeE8+4DlLZI3G3IgIHH7m/
5JjyikUOUQwNK2ROsxmZleemkX3ax72zYe5VOXTminwBTtmx9OvZonoYYa3F
yrQjk69Tyc9Yvg9q2EvhyjhcThCb8/2kU6cI4tvcS7QAe2lSb4sRPRMqDMhD
tb9rGyrf+2FBqXLt70twnxG530+g+5HolysijVMFdinCmxX+aYklcp7Fljbg
n7jBObLy3yJMmpTZBVilhjPLbHIGrzE/cAxi3GaglnFX5aQM6fGz7w8sSOQL
YUNB2gev7xMpAi67JkJ8dWAexyGC2Wik6vL4DQcozimNJAHTc2Es4HBg7poz
sFX84UrcF03zb/wO+h84f3C5aDpGDNDE7PkrXDZegIE2tJlAvr8se9h8fgUJ
HMcCum7y2fwrTxSX4aQYWFqu52B9xIG4Cxzd/D2tvUO6RVfrEG1SfEg3W6VG
iG64OB46POB8D9SoRvxz0DuT2Z/vsOsJIdZqvVfyIZXjvGsW6w4Ol6cE/ExI
WGYCkibE63RKbV6lxNRmaEsDARrq60xLS5A1ESpJwCiithhBanjCkVxrR8PG
uGYsjFnaRJDus3e6bCnO3dILT3pQTNyfGfnxCs9fCSzCYZPCkQcDiPGUuiIY
n34ttB07L/PyLjAQl88wEVmKYgfMJDY9uCHx67Q8iIDPxZMOTeETLrwiMq6u
aoQ6AkKIGV1m5ikuZ8MmvcvkARDjU0IYrU+ynzfJE+vptL1a3XcCz822KNaP
DYhYT123esm5DjpanK8/dM2LejAXV9qoftlNuyPkNnawNgQAhdfjXs4ZkhgB
NbLHR07C67UhD/rZO7dXVIu4Rvq/+HPuO5LXbFou0vrXQ331MLpUggg77rPa
bOD6kpwgr8Vjc7psfL7wFUDx/2P83sCOwxljIgI7//x8vQF5BjmfZHxLimVe
i+nuj8S9B7cZEhv7QvZ6SRN0oGmVANsBVAA3syLIjXdS8ZMbBb+ML7tez5DK
iUrdoCN2SXK/FKm8zvDHTXFyVgo7X354ecBeQ0n+66RsBjRXwST+FnFyXKao
MGCaprndbN56/SAheOBSMVPM4uVTvBhE3Mezuqi0dsEgxFU/7I8WxkQVHPvI
D+IGIbF0FeretA4vYyy9KPDA08lkAfg7R6xmtYyAq7KcD0yMOt6mRVGBcJpo
z8G86N+Ek37YLbI5yR4EM+m77wF4PNxeiqe21g9TKWteuXg+fE0VPbVAhTjq
UKt1IqTkjrgaE9j3jHzopOxcxGU6GijPRuQ97/tNpGEZd6vO5qEKsJ+6hC25
UOJclQhh9kPwdSShpi95VAcNhDggaMiqr8mRbQEbEg+LL7xSgpdJ/Z54YAad
ZGNZL2zhTvtPXhwTkjt5pW5lUSuOI99GGEIUHfBC683WwOFxRGMjSKvSulzU
YbFlZDO5UPFFG734AR5aKOki4bqc1V5yEwDqoy7KLBiHCWxz/OxMqL1d0J0K
sUdxy4xqc28wYZ++zA8gXOUg1YFOKn6U4a3NvBzTkpkjCqQvkJnXthXPRjtL
YobhkW2K1t1IPFVU1VtJI7WbapkxNvsYu1xgAmBgHKBL6OgTX5/bgIsVfbGZ
4qcqyKfWVmKdPaAwRL2W7N1bO2I0nwWrxW3QDvEGsAMTCPvUZz4rUPwWVIi8
4zjiBcCeOFWrvYAMA1d641WOjcDqmhPfLs3WuTJUOO7fnRMN9idw76fI6tJP
iEqFwyG+EaYYtYelL0eGCR53N9ixuboTGOQxO2KhtCSJLrSYhVxSv8HO/qVa
H9JlNmOqfjG+W9SFImNxHFM53njqXhlloZzgH69ss5PyJgW3X1mP03rsPvbC
NlACzzNVS1j5iucK9nZ2Ah1XIWaoTBWlKXKhAbTd4neCpeaw+ZDgUExTNCec
+7Ktv21FGNcEC1D6Y8ot65KWzlUYxQX7FomDXr080bla8xQlqnNMF5clxj0x
UorWIz94Bp/0upcU/eqtJeV7PpX01H7vC4Y+tBJ/LF8n04aeAp4PXAFsXVx6
QkkmtLMmihLKSWgf3OAZ/CqFI+rBC3YGsHDmKcSHZSH0Ve6ftiYIdgGaWkLm
yNDUr/ouucA1J1BlpJlN24qkHY/TwckByV7cQEY58u83emU4Npuv8XRx3FJR
zCmnwrBy+3JCiPowqR5vqvsc3K6hwJRtT+5nwOjmfjL+G9hk/wipVgdEn4Vu
eU/HrV8Gz8RZnRRgRJIdSFc34m7uxAyRmNa2SwbPCPSsyOmxCnq0evrzV6mx
n2Pq677PXEaO1QrHVqNR6sme07VLURzq8dHS9G62nUr207UeLB3GQGrP9/xg
E70xPNUutA8vsZpS6YuStMmSdbZYdvpbpyntz8gJZztWfY7D9BS/r8YO30U7
EWKCwjQns28PCP5DslAkjQdVSTzULFW23h9Wo3oRSAPPtuoIc7O6BfU2cF1s
XlmE4ijR4OrN7qSfE5kvDEO5HsAXwEd6SE1ocPn1F7ffGirW0Md30l26J93o
MhpEpB1gTSHsMgGUz5eIkzE0CaTZcBxRopv0bqL1qvcJ8qjqNpGoJ7dFjp7u
KGPqAF25K0RAuU/rId7WS3wQ05vJr43DmuY3z6JevhJ0Pg2pIGTyyyqOhphA
pqsVQD5WEG9U7eJQ1QZYxfWG8KUrfkuTJZGP9V1DDyP6ylZhJ2+J9AmBVh0J
32pPTJzTjvs9JwpIi7d/iqrUe19ZJ2VaZS5aIO6aOrCVlKqVQOmKrREz767i
Wr9UiLTxTbNNR1LvA8yTk2R7fwJ77jIbvR478/264kCFBQmf1eP6CGLIhZdR
NqkFyXxee4KqAa8JuJ5Cz2rQ45pBX5MNjQyQb4UlPPr9HI04SN9U7XY3IR5n
grgw5fJFIDbw2aRSaZUfZ/jsF7beAtp9quTaROWIlNgjQhPs9cWu+ryA93mx
lE62CeGWGsh6fH+p+xdXJI85U4MpLi0VAnPvdcnV6S8CJHgD9mWdT8eNFYSt
hLuxo7aKMVjNv5IOBK2qedt4WY2wQykE0YVqLIPvLLlm4hRBtoiYEtID+/u2
uK6iFA54PXEWM7sHTz00MYC2XLeE936q3E84XEif+fxWlvVglTiiu1Z2Tkxx
LFldFVwdNGdxCldZ3rMZtm4nPFRLqaQqdVHw8J0jZC5VhDM/0yMnpQNnAFF/
TkXrJ7S8AGqTOhR65en9FDS9EvGlLj/qlJCjSeAIZ+tLmSXBPFPZ5nCxjRf7
B0NcHt2QfDQriSd1najcUT6v7KpQB9gZdw/XlNQ1UpmcQYQWUBMpIEcaYeaz
e3TUR4nrYpWfX3CEQPjOgzFEBEcdCfJUCQze80PwcHJRjh6VevuPPX0ovXxa
Yf4gYGQRJhsT3R3g379jWcBX3pNXKA1lfFUUz5iBJJLCBTC6Hw4JNTThVZ5B
vDUYm+Qo7zOo40Q2hkLFOvwB9plCfzOGXIRAC1ylvIPsI9o0hG9jV31OKhH/
u0W34NjQdokHBStNbKXPYIwxZ3NZH+Hc4xlhDazFtArdLPf6Bl1UevdIhn8O
q3P8t+nbZe4KOx9VVguOriIOMmzrO/ZtL2QOeUZCMFZM1pmk6X5y6cUYOXa+
S+YQ/PI8QcBXO6Q9SMNX5IqNio2W/80IQENUMfHil82XI0Cz8h0BBEW2ocGv
F3fczIDMuBLgHk+k0nqzOnnbrWz3xues3GlyGACDGtQG9xUd+ZGFQ9xfGRO1
k3hS+lx0iTjl2yoc0pofA6NBHX6R+c6fpHQQ44iidn/lDjVDTPoIlQzbW71z
VR+qSa5yv1KiGLYgakTdsXc2sim4x3foLWKgdfvCR3jr72b4PRexb06GBBxy
JyAhwy5hzl5L+j+Lk9d+qVwoJp4Shyz7CBezl2wg1l9Aar4dXL6/DDAEOK3L
E3VJv0sJmsShQIKyTVOX9VmSw/AGFrlYC65x6T+bhdMAqY2TQvOVPO3YbNOv
cQRbmaivZOjGx8SihkN2xsr7WoZMpHnnPgbRT116fix9+eIw5IPHmxMIEeQS
nzsddvOe81+qfSPmSTzWFYllVqPexSF5gKgeGcxN8BeU+M+ES5Oq8VO5RKQ6
BNQjMSkddPAu/1NobT2auX8hQBOdwythQYDAInE2zrRjp6nZcknOVoqZzGAM
YNgQPyWgjViJhv3DSAVU4Z0A36xUsZKhjcFRRsSSgl0moslWp6vbta6DbIwy
GNabVwOvEtygTR9C7HWr0Y/EtP/kQ878ddFK9m23l3FyJcLIKe76iE0FnJLZ
MRy60DDLLjvFCEOP9OEe+6b891u1uXukObAKTX3OKv5tRGOS/zwyvA3rDO6O
yhfApJcRt84roXiuvdVOP9E7Ik7Y/0JVGP+BujFifS9/ZsurTHreR6gUJQ7n
w+TqRRdwkuePVn7CGOgx2RVxaenNwy6S5M5OUh8r0x8ZSr8iEi+ibXaVak0l
mbyeMUOs3d5i9HuGQRh8xwl+CA5mtJI55QDjTshW8+eOsZD0rzbiIukj0MGH
rq5JZlK71YiB88TLPT/dO/Rphmm6ikfK27JskpIqpCjG/eRP/6d60xqeDJS7
LhOQd/KKcql9CuapubmNbfvJC42cuBZTIZOOmh8ez35LwCdI5D5CiWHGd4th
52GcBERSJ6hbhcvYLhoqo+aw8XvZM4dX2unbKk5Iy5S8+XxZpKetaYuqV+xA
jM3BiAZCuDIG/6vceN1X6pS4HlB8ZBG5OX48s5FWzRCI5yl4JR2Bfu8CC4xs
13CqcAKoStqMsR1vcgmmIgSQC1DXQMpPfNekS2zUSh80tRf3PTQkvnezpGY0
nc8gS4sNaP/2UVeUOeTb47No3ywotlXeJ9iUj0uvMzO61k0sTsguFmfpdBrZ
EVQawMQ3MKt5ICTcE3D5zgWio6tGW1Ujq0L7YMaDUc7t50E1mbTrlVjY9QpO
N1xERcoMnldFoFpxxawepVdD2VrdoPJE3OBvdGh4xIO82UtQgnwBXT3ZitQG
H4SUEerPt8IBca8Ng4wAAxzZXTsKLzZIX6XOI8Cdf6iXpHYlvvzH5F54jh0w
uAmB7+o9VHP2980EBiZ8hMhO8knK/H6qKYFvA431jVGwOb7owI+lLXM7/xqO
rBxusCEq9XqIyjZpQl4AGeUxjDyH/bKyaQXiGcOb8LrEPNTlbD1kuoAxBQH2
VYRxIk6yd3CtQiMhtSW/Pt43L+mjgRK0OjIHzY4+dAdkPl6S1bnmrPQFh/Ly
NKmNZJ1ggzmI8hztwbdyhfpuufIDoOowvNa2HPmNFNyZ6Dws2JjPbKFdEOrZ
ARgwkNdVH955tH0hdNXEfx9HpXZsUx0TTwYHIgUPPaXgFHN2u8bk6Un3f3fA
gxUzls3FwGbWT4+6xuZLp+t+6ifw1rbLghFRwVLG2LlYJsUMOeLDYC2u4cpI
BlewKs1jaAcEeFYxsarsmlfNuIiT/k8lK2H2Dn4XUqfJv+jv87+FupoCXkgW
hP6LcRVkmOf0OpgCyQh3NqDW+U7IdSVuvESb84+TaJHgNZt+4CAUISEvCSD/
5ktwymbKboOnjpmAbB79mnC7RmMXJc758cha0FnV21nX7rx1KXpato084dqd
imhAq8yG0Uo12TfgstPKaIFt0J3tQHLQi3oGvgJzK25qEZRG2w9KGTDV4P7l
vOJaz7XmKe6P8ydn9SPS17GVIV1KSsxZ1Viw/XUToYg1EAXUUjas+XVUDzGk
SsnyIoVx+sskX3EejFqLQ5NxmQbFs16waHt0ra8OP9yWoF50rIq91ue/0ZvJ
9kcrdEP01mSBApj5/n6RugMyov/O9FEBJIZBw27WG2Kc1mGJtp7hiy016gGG
CkZ6AWCftjYOjnSi1e72d4ZJrbYBYYoZIzalSNabWHgAYi+adDjIBehvi2zH
h0RxEJ43ShVHpO8AKdk6rMRmnxATgdWtvNQz/wax3pzuHJ5+AI0/IR9Rawxs
vd5m7T0t0eywWZ6NL5JwZGZFp/XoBuF1NJACpMpNYxFKu9SshorqHrq6tp6M
1RXTAkQDiCqItYDkgK//RuodvDJUCDW21wt+RJCjCvxei1aNi9wlugOFBKd1
gASMxqdGheP45yjIrn6Soo6CoNQSJSf61KAeFKlxw8nEK7t2/gh6zvHQIqNN
Tyew1gFU8L4h/h8yH0w78fOP4MXNZCxHU1troRkHnj5m/6iTBnSrbyA0V7Zn
FGx/fRFe3RYSWHB5ElAvVh6w0usyJlwW9EvnwnVf4j/IVvNwZHuC8jPACVg/
CRmzvlPeAgqGMag4vZGeJAj65x6RXkYMfnAsAb8lgMjwo2B6xfI2PDGtAIyj
j+Vgs1u4uhkUIrgEp8IqiIjQsRNMPt/mYkTUpvx+BOt0ThCljw4F5hJMkGWU
kOJhQYOxXBlV93n2I6HMHx8hbA5rHvESl/q84LXCm0O+tWb8oim4NDa5yyon
LUhrJVk6uMQm7JrbhDMA4V5QwjZum9SLY4bzF5nmWBIDUXHMWYV1Ck20Q4j1
8VrRFsAIMSD+oz6CgBXEXChW565GdNFB1GZ8Wa7zUSRU5Szy6/L8MATWT40X
yiK3Ra9JEw9xDomOgrgulvRyO01l4IvYB2Vkbw+uzVeO1dv1S4+RQtXSL3gZ
daHH0jI8fwbFMGoJJKQzjmkRC2jeGdEOPxBEnC5bWmeEtZNl+E0rLyiJVOhx
Lc2xPMlQAXmAq3WIPeuX4oCHlNFucKoDZRE7a60e7c5iNrj6ogjPPQ//Xeky
KcIhZ7H2whJh1vWBUteKkskO0J8G/djBMzVE/N2ZCwOtVgSR54Z053CZskXF
4UFOTmJZ2VYQmY4qcIZARpxEAQ6eRSJybKBPdQHJhqwobBawFWmgByyqbkTS
T9nM73KRkTXs5cTJLJFGmf1yylV97fpdYFlKXV6MApFEkh9NS4RgK93F/CG4
jmZNSP798XYOvB7jVJ+ijCH/rk++lv+a51RhTbAG4N0AdXGAyznKbmLBtmpc
ZDLXuziRyZzTWmOQOspm5PuUQRGD2OHoP3+99pktPp5HQsPnyYj9CEdr3niA
+X0HRhUaQ7qgRI/HwEfy5mYMRK8ApBi57nKJRzC+O2FNw93kl2ulVjpom/P9
jy0VyvvABBS9TVGw5BbJLFwLoIggMT+kCy7SMbfe5Ltv9Y2XR88F59X0ThJx
FnCo6btMFWgxR5T1LiDhXcQL1B0+bJdBRy6E1VmnsvwCQn7nqdjRdhCLlNMI
3s9ehMnYOFKt6D4zL1NqBT+6aSU24Guqto5GwNwDKYf4o+aWXp8GeORlI3d5
cpNlggXNh2TZmxpB0CuTCy9ZfVBkhKfb2D6daXmUK65Nqt5RWiYHgfnL98Ec
wYDOJHyNruCkuMJabp1os5Z4kaJ0yExTLKezNJ7ba+dB1sFh/tXPHXIw1Z97
kY7uU7K03ZkxEzMMAZhLvpG0yj81mz5RmvRLXlEXi36d8xShLkphQ+g+2C8s
yKxtLuPYFz11/xSjcxfC+HX5zMNqgR3BkWl3GR+7/6rRhUJRoKaIVwa7RmMC
PKKoRkOsSBBI1v+y4e4TOe21DdAFkNMcBmko2TNk7wksrFQo1K/6/WM/Wqeu
SXY7/IqNA8YIdbsubfi2VSS7Q4OPcr3vC6IZbWN3cG/INqVHVrm5enm89a7f
vo4JxDcTBVEm+94Y6viKpyzuKdeckrtxdEURxGPX4IQdSzPs+KmM4D9LfF0n
ptSJ39TTCLEzkk0mTj6+PWAVxr63L4wD44adngbxtnfgQk4kS82pArc643ta
QstOEKFjTBt2iraYMBL2x61D7R5ZVrMIRflBO6RTG0loZTi/yE1rlmtj1xIt
7WsebaN2lABCm2YmYwcD3pAjCZxz+yMaWZmCdrDPEvD6/mTE1//ki875NWBh
FZEYKVapAPwM7kcAWN2Z8guF2oOsZn4SuDHotkE0/wteuZthgjhYHJGJkEGz
x0m+WPpwDK4+XEI9XoTwe2bWxIgVUQdrwzGL99twby7D+JPXSuCkyOzQORkj
C/OCq6yrU4kLo2jcpzXoEzntpLYPFPpEKHhu7vt9GleDnAuCcbTIhNErtOJd
OQnjCFZ2VxabX+DoEow5NKDGHtkmR7RiltyQ0xWxMWq0lu24f2pXDngVASsZ
xpTC7FiVKDddKSqOqSTr5K1lOPVbHM67prdhfVy/7L/cgTfxEdsCkkjN6b2X
ohqicAPb+2/hOLynPb+zH9ivGubljoE7ZGMgNoFJGQxA2vV/sXhDq6Gy3sUp
LoSlP7NHDOighULKMkNQgCjIEbEd5VIc58EKOzzAUD8myxS905HKOzRJrgmk
g6+Yz8fbT/QD+Wy3UhF5dvqXlKOHxjsxl7EXZVSbHmkgXDvKF1ytiqTacScj
F6H5A7vqRmZG/2nnXibt4zeLdmuMKcsgmeluoMq+0QGtgDgaXoTExAxr8D+7
cihbN8cBzdLvCjUbPZ4I8joNYvFkkNbPwCwAqgrHGCdipzD+s8EflsbaXrQJ
lI1wyEuKWzfoh2p+PhRLj94sYgk7/uLRY8EiaTBIHecmyS9ClXkTPER1pDrv
J+ViATPlw1lRg/AlUydcMg2HxHnByP+hloMGtzQzMSFwtscUZZuZr4kuBnZL
vDHmUSCHshqwn7emGrBxBx+TiPtEZeM6HtYc7QMmxiPo+CkaNSBjPupU6yJj
6cmJgSQQ4YUueDqY48WZ2DQOrDwljRQoTSYwrDWH9zqVSuqQ1OYtByAzKd8z
WESr0+TYtp+dK/5bh5tEcvA2JO/C/oPAQqx0t20zUUN1Cl4eTZx7eCPzmMdr
qvbg3LE6dgdVsYtOB/RG//P+Hp/aBX+7z6WCws1qGygjV+vBsyN3nZbpcf9y
JaVY5Xk3wqKe0zFBoD/6+STaFry3spzbbqFLt2xz8JNUAdq5x1s2eRLyVdPC
JZ9ZnKlRU+Y4xlRYXOxboLXf47HMvujvVgA4G6M1vQV8vPuGDVWzXbiKgIt4
AdV+/ZN327nj+3/9DZzWseJqWpFPYP7kVzSTo1GEJJVkrqv/B9hcCOuK6o4m
LXOCj1SPhYO+zqISnJ2/m7x1JtQvLyOnVtjf+QjJpn/I+W7TJ15ztoA0wHZc
dYXyDZi886mLYhevetLJo6ipd1+WYu8PqnBI1dd3fbbuBS9LGN2yI+9XJqy3
vgk6uACeIOfi04JKurfy49p5+lFYj5Zhrj2o66cH4mTHzM54/CpmNkF7ujgR
PZlZpaVSBMm4cHwajVA4F4x/WclLMiPCc9TtnoiZMRgwzyDCyYX6jqbljJ+h
RfFL+3ohZFySmebBSz5Vu+OYSbtpijfasbOolcaiE9qFBJoe4H3KAmVxxfUW
b1VfggxPZUZzBLR0oyq9WurEQ7nw1J1HAMYydb86RUeZa/D0SSCw59g70J1a
MA5yn6debIiQFlCAX+il85cRg/ySLWv7tduBqlKCvMrGv1oahPmTaSVbv7/N
aKYOoyqQjhhTIKsvVzQkSvyKl2icTjXrSOvahHZFzJjR/h7bCnF9mbIelIUO
w9nwQ7BySm+EiF4knAZEi0kHL4pYXbMDJ7kY0OxjT7vYIWHEhJTxO7z6lliW
2jcUyCb1+wUh/kwMcIMBMZEqccjCTAzYP522uU1NE0LT6SZjHGLYBVw4RZQO
GkfaDBGrrYAHgzCqYRMidGvn3JcV7Rtli4maRhtpsPLPw+qhsMxCXIl4Sf04
rvLxhiyKhiiO5kqyszpzUMvpp9t/m/mGECTzTWc5eTTodmw6pR4iENmfKU+t
s2p7mot3nELDezAQAYRX4iuhpldzEKWPrBkkmOFTFuvloCAeEuVSxGmhLi4j
1x1OBhBmsBTUp7NKEvbzCBkLoumFRQHswlkCDB/bbVuxsRg7HjAsmLGgfztX
cRNW/+NJy7X2T0hEbdBo7pPHK3Cw6Fux0Ogsh8118CTEzrR+48jR4fgbBr9O
BXkBt8seTSJOe0Hf2zOub7tDjKOrJMJInXWQVxNQsw+H6AHkDcBSLYxubF6C
CoNnrp7iKDkZIdyl+TNLRhPpbqHxC67rLjSvqPk4pzOjfydhYqDqXCKcxhr+
Q/UP2H/g10w9yekbc8rEI0kIACPtH1r9ZIptNEAPUXJUlI51jaOb1uVAW9qU
pCDarrcUh2I1NDh5vXeCuoYuGJ4Y2iN4NAbY7N2zz+0aKwxX4vkrMS68RAKn
gWy4M0nBY73KvSmXkms2IUwTNynXg5hlykEYMz+qRuQ6NMdHGqSYo9yiaz7Y
4HN9up5zAL29vhcpyRDOjQoGCwGAnehGc3iiSxLSiu53I4LYHt6+dvgoi2V4
6wxt9gVkp3AGu9G01wKBZtEbF2yuGkQpzLjS+mucT46Hd4g8h54CW8gZa7ga
jJW8S2you1Hj7pNrFIA25B5MaqT7xrW4yl+JkmmHMTzQmEXQKACdlgQuCIor
7DdGEHiPD4ZxBCJWCkJRIIPNdh+rLKyJ3YBS5LSjRYzM8tVjinLmzZZbNU/y
TsQOtFUtWq4iRobEdoWdhWlPXE5YOB9Z+4M3s83iTp6bO3ff7eUOac6+aK2l
7YcaaZn0QWI7hRLrpdyQZec1APQRHVrLWqErL6SdMy3R/kW281R2IVp+jtXs
qyY9yU6rcznzyKieyj2neStOFU7gSCH7Op0ulMk3LNc/P7q5EgNm2mLX5Him
6Yt78VuBZrANh89D88R4WtoOPJdor2pXMYwaB5aQ+IFlkLNefwYORCH9dlY9
NF4/9GdDpUjC/C56PLZAdL7UygpS54QztXA/kTE/TPrCGZQmzC+jVxC9A1HF
34KYPKeJHizrYOXNa1oI8yzAxpuP0r/RIPVaH0iIpx5W0RXsjE23RyuFSSOg
qo06y3pYG8DR454+GpdEmQ4jjG/R7UonME4AxRSD3Fe99pz/Yi0wCSPbNjcb
itRil0KL8nEQMaNjUqN8u2jDUATKot8x+f28ufUJ2/MWUcNg6zeL8khALMB/
T4gjBMwRc58/msJstncjjKdpJrDNMYuMZvYicdlNp4pbD9kwFuVPMmp2Vm/M
qPJuwPtT9qHN6WpklHyh7zdQ3zSxUKE3cW3CXiNLB55RW+zMjG4PURQCJYf9
1hK0Ag7+awuWrPV8Vl4sIOVkDP1yDjS6xGTMatNYjA7Y08/qCX6qwfWaK+fp
RTfsVfALS4ijBYN/jGviZtagTxSI30NG8gdF9d7apivvWIcqd817/oi/dWZx
lPovIKv5qc8CeBWoyArCo60jj+nw+bdolh0xpL26iW9iS4nlurGpmJPId0n3
eTlZdjWDTOsv39ATvPYuwifztGGlrfXU+zcgcmO/FIdGUC/UKk50oTeIu1U7
P6V4tqIc2E4Q2oBSuOWtXfvJvo2XV4Fn1n+sqvOcODY+ZKmwA/Fq3GfiKAjA
dGdjm74huTIBFJ98b9o2rjuUxT6g0Q4TIw/6UyjDhQ8Efw4BAul2u9/wrsJ7
77v5zz/VSPvLT4LfMwF/+U03wZijSTmvVbksiJh1cA14iAaW9ukU41FXqswz
U7AAjjUcxdv/k+I9Ek70fiUW+Fo4K7f++1H6CLvufmrEwVM2VNI2B40Qwovd
dZsM1xwuV4tjpbLS/oKEDnWgmw8ocpri+QCDx1qWoKMgl/Gw16ZBlf2B1Drt
fvZ4JabeYq1DksViEjJecbYWtfIt21QkGAtw3NOi51A/vtA96sVeURmrBixq
Bev/gC9u8n+sX15AhmyaD3vB6lQlTdIKONCWeF17IEsgDLYIaj6NMVF8SrGR
wuykleulxPNUZJNhmETLWis9oltFgluC8ZbHbleBFx2KIVpbYEZIQODtcGwO
TVv0oeVQLG9z798VTPEk66ekmYnNBc6hovFcaYi3wyknweix9riS9xzImitc
0srBQ/ytYUui/cWRa244tgi/tgNrjUXYRw76s686zzax6xo77dVnJh1vMu46
sUZIiMcXf0ce1HglZI7sk7sPjJeAKLumD47/F12sMqWZlu0iRfW2SA7fFct8
ep2z1A/m1to2P/rep2z1wRPcz5z/f8CWKVYp2rvFJoLqGSCzVZxTmn0l0Ul/
2MP0QfaEYPsrh7yDwrrHybjkK0JMbWg4lSsPXCqRXLTOjPgzJKTHDOBtaWAE
skgxRj0f2PC9K7Jnp4qNM7NwwRcAM7Pz9HPtQnYc+yqVsXjN7H2JLA6uHjrm
xMKat5IYLO5C6jEz11kxcOoj7RpTC1uIpX5jSJ4PAivPTOeR+4EmuXwaOR/1
KS8qvntiwbnRPbXwAZPyVwzfjNEovBkgrLvMAtM2ObA4eBouxxgBIFh8xW8l
2y6B+XR+I0aE8V+MAvrogohS6+5IVKZRk9jclux13PwJIOghgF2FnjQg49RR
Aye58rcc2U4yYJzWkiOuqaV3rDt1XtwHV0bJLQLSyyHODvHj2cRBSp5l8Psv
AriVnbdAehkWQGgEnrpz3S2Tp+4yjleT0TmW7pG7jtMSzxjhWP8u98ztE4fW
2IRkJjdDey4FBy5HUvKt3yFYqXhUvigQw45V7V6K/Li5BsrMxOcD52LBvjc8
/mOgSshiCMlcL+josrf2wiazTGIeKU4FaiIRLCabyacHVX0nHV0OhH8G5Opq
J6WiTu8q/ftue6dW6s2b3K5JziPGCdywC+6iDxV6+ZpVOnY2xnXpYKeWjDA3
s6qz9OCjsWRiV73jD2Uc43tMENoij1A2ui4LoPqQOh/rmMgdes+kbSUrWzm9
qIJriwrGGPESC6K3tfmcP+GpW7xVG9E60Kpdi3r1T3EUqpz/orYPV6Dstb5O
y/hxNDuxKtmtvrvl7BwXI5Zn2oXSfdRLgYmKs7wAf7oCzDL+Md+iNydCMM04
zjL5fHiEW2jC0nPkMtMUn+T3eH1IuSDA7JWdZglAn0DFqTYYwCorzPXvF0um
Fi0s6xvG8g5RBhBaFOVKbT5QlDNrup+R1Ta/biSqdXNyzUjIVlYV3s97lKPJ
klBK8TXCHbL8GpHtbx1+E9Jc5miQ8moSShTkwhFdysnvBXsBPAHrVGyQ6vaZ
N31G5rG8Fv/962mbKfpjP7fEiehzjSyW7P8GxAJ8+RnO99OuPw9nhlHLZ84n
YubgdYsVbjyhiqKsZIponIqbSUs5pim0nUhHMazc3v/UfGrbK30EmNNcRVu8
kPo6FzVJrokEEhgrMePgfnOUlK+f0T9a8nEbWSO9bMPXfs3N7Db0MGrwuCQo
d3E+iNF3vMPbiWZI4gUimxVUvTNNM1hwRhdS1KTqgroQb2J8mtFT5+YMsVwH
qrv7am1ZARIgFM2i8mpRu+eBphaj/WeLDWP5fh0SWZ6NlROLuLMmYkSJeH94
gPy6YoGaW1K7Lv1SFelHd2AiYX5Z5r6ifapN8uFUFzjJXobpucfFLAGJTnNf
+YKbOyZI6sZGsllRDifytM75VXRiHubeuG9+n7Ugtln+qNzCEthhN4+wGydI
mibLISQxHJ+c0LlIWraPLkW79boeVjApKB4Ydu/ynibeVIfFxs3r4NksGodP
HexGDprk+LLCqRmf8hGcSRdDEXzj/G0cPMxgGh85+Ax++v8CsIcJ2oCinTeO
rsMkCwMCh5jlURzhOFkqvtObvaWSb+E/JWtDGaIhfRKUETagmgAKGo4YSee0
vCTyKLagqQwwYzKMXmpsNqBz3axihhrqrWXVUJOVPuYI5QssJbrxDPEL0W80
aMYaN7Q5GR0jZNLBv2ldpvjVk9QUz7ghmgnCToUYNlx4eVHyAHyZZlHgg2dv
ZoW91Des/o8OVAXp03MhAROEAUscWjskdvy1QE0WW/91qYPRxjAxyuteWWy4
5PgB/7bz5x926seVSS4c80P3r580bDydNhaYYKzvHLyntiJOvyDz4zWXbDT4
kc+ZyDRQErWey1k5e9jqIJMg6LmXgnoaALIy5b7YYXIpMGvAl++0dN79MV9C
sU7KSxmtHVwTfanLcH2S4vROhskkt/kV7+5pi2lubSo5ucBjcmAv107lhJnB
YZfYOmFpLPep+txXWG9IqP2jt1vP+/l1AlFmvsCPjJbXBLHwOf82JA/UDRFd
NP6YvMonlnQ9bBszgoz5PdsjM1oPnZW56CKhkZALNPv9PQo6Ocl7PerMu2W7
yMYn+Ml29RW6Nst+PTIycC5odN/B9eh2DRlJlKWBVjqiOLbV5wYIH0rnHZKC
vtwghMZCEPzDek6XPyLO3eio4Hz/MUtjvr7Rr1pipDfpN81jaJprRvB2JGPl
I1tw3ubOgIswyykhzrwAD+Ey5ULJeKiZygVyosjwdXgbjTwleQ/v3mMKEbpN
BTIMFKAe9EWuukzWfcnpWmTlb8PDoO+nRB/58oBFqRadFB82GO9J9jaQig8w
5M4RLKJKs8WnKkIwcWhOuOswwo/PteKirjhjhAtSmi2ZU8ba1qPgk4X1zVva
VBIgbK3SEa0EREoe2+qbAiOYyCbZaxdkZSy9NuAalJrb8MB2tqdB9K/WFgb9
hmozbe2BVo03gfhQbtMAASqx/vHK0d6p72pYARN9WJltnvPqmvu1DDsce6b0
WU1I+Znyshx8Yp4uCnkWjsuH2LZ2cQl/I/sixYRNYYRA8/bn8HgE//9QdWJN
jqfsjFYGAmX6pFNjzF/sfC6tPXzZ4mw7zvb25uZuwDRcND9NUf5lFHfEtyqN
seB2EU+c8VufdUOuCo0Oallo0R+78hsbUbSZV6+d8Zvcelpk118Vrw8TrDhx
N98gTn5p7/Fk270dLDUMNXgf9dYtrA/hr9t0cLGgOscyBf6aTQp3UOMU2jmA
VETVGd5y+HImjraYH3ZNUIDTTp0SKoY++jENHQENq5wnNvNVfwKkCSkVg+vD
cDQJq77TAjn8T1SC20D0fkhVbskG5pU7VAcgPB5B5dTGFfWdWlM7BlSeeqja
dYWP8pppv7+F2E5L3dMuw7dByVHmdMpG+MNT49go0RlKEgRx4o/FFMEN3KFu
obA3HLlGlFftaMt3cjh1MseDKsjvkM0nbbLKih51Zhvf/IYckGBSNUb5/Sv3
eO612JeSiFh9gLwH3eFmm/r5WAEkO7QU3AcARxL26N0NqPWfdGmiV2Ob74Ih
3aQ0OOvRPrLayLlAe0FHfsXE02/FSG+2yl05FbU/jeUlDv30VsxpzOBiNDl+
xsEcCa5cGmSLZn5W02/4aczEBFD2C+9LXq3DmJb2mwTrNfiPFSjRuBTaBVoA
AR9NAWVsDD/uimwneF9HP40tvAnmtertoWKpxbeCh2jB6QLc98vhY6L/FltT
zx+BWTWExgicOnAuWdsX9g8s8DofnMKqDM96LgQobox5Bn1Kvh8lZkUYPRtY
0mu/mJ6kQKumKI7BBENAKr86l7/ltOtwyplGSXRQfkrfCYDbEhik9J8/T8Si
hmlGRtPHHF7zNdCrLikAimLWeFTeWwgieLIo5g8IV35RWTeZpA1Hp4RD6Bs6
xansl7yj22IEVw9sMantwzmn7ZYFQmVNSWt5MGfcmH5vWAjo+TGITQ3SmV7T
P3N57U0xcx43xMAtXuvK+8wp8HADAnT3jMb+4Lb+UVuv+x/uY+GO9FLL/jXm
g2nN470kn7LV04gKKH0QHkXAlUMy1jSJwg+okRnGRbCVs22/V+IjLkCXfUZe
VCNQrGm6wtbIhezAPMomacCS0i5FWHRpce3UTUmaxD466O7WqJpH2NGrfdaC
utS/PcV2+amuaJjg7MwP94m3t12VZGdn7JiT0ysJSBfXo/JwguO6SE2DAve/
AlfqoZaEf5CmBtbiKw2Gh9miZporTncep5bRNVs4+e2zdAGva2hyu6djXsak
MCHUFnHDtEWhDVG/UqTScDkann20ojqPdflJT42PdHdmkPd8IbDOv87RN7+7
6ThXgImhM/9Y1EecE6RdZ0vO93TtWYTPMadpybQX5JaxfAvKlTnQhNrzUplY
kdrn2cJMezdkWdqhOUNiS2XK3DENKy51i+0zfsn+tiIARxSOtgmhwuiLpfGf
auaFfv/TxGbG15FPPJOI6w4Xw+pNA7feof65gQU5XFXiDNXFH1L7JDJvJIjE
9ILwwF9EJYBxMpFiDI0JdykOMatpvFsEaHlTSgIDw3M96u+98fa2JN86Urtb
OX9SeSvSBmrTjVh8cIi9RbMIzRB6b3wNwpXoszS2LRWcXvKF9njUKBO2sdbS
LCL5Pt9x/v49lrySZ/FpmxTV1gGiAzkfzfnBP6dOksCiPs8klnFPF8fe3P30
8+6XCSSUKdU95OeveI5gSuX21dlng/kia6F4ZDCG/8LTaRMU5aPNfUKxyIjO
KjXg60LobuY5PIuLNPauMDqxWYX2waLNS8zrmu6+d6dKtVKebEKCl0atUQq1
iN4DvVyKNHTGPpxIA7d65UVfe6JGdRMHCTKfw6wXMASFVhdmwud+SDjaJ0DL
3cpuNhh7jX6IPFG+n4ck/SHjkZpLkQlSmmFebENkRSvPfAr72+yshcfJgp/c
Ij7TgufZ9muNLXw5Y30WcdDS8aVAltEDP2cb01smFsifuDviDXuqSv46xQxj
w7gvIEw4DRTkboj9UpfWsZbId9ljh9s+oMCSYVXBM521Sa84LbsmIg7tYe+Z
jm3hy7U7lzbhApFX9UkEHZtY2EjHK4AIoGGL5EPvX5kNMVzCrqPgHabAG8ad
so61lGHIq1kHW+zptz+o2y2KsqrQ77RpRaZ0z2s4or2wZS8GputkS3aMNVeG
GE2aIB8kLcHvCYakpEapTX8Mb4C2ISOYaoHYqX8czdtOLCutBQ2gEY/vLjKu
cYvZNCeivma01B/+4jZGPddm+CBURjsDzcD465EeU9X1OvKikHkYa/KhLird
2G/2rRbJLEsorBKaM8Xetc0PGKzgDUf2o7zmk/nq1AUyfaUPX9dNXuEN4SVU
6b86t5NeBAOtq0tn3DfvygEbAxCSCpbjwA88Bes89nQ1WfJV1Pqnsdd4H5Qx
V/QVRD/FjFLjcLzHa9i6Aq8EE6gprBfq+UGYomNWgGa/MvXsjlu87lnbpKXa
kAPs8ZuoLUBoiyeTcqche7lk4cTgLhX3keY3NjsneKP//XRsfYeQoHqMwlN5
KRFtYIEdC/ZBv/1IogTsbBtuDXqFlOdlKWjj3wN9KgT+RiXlesbderydHTQ8
vXrF7aid3WW6Lb3z9TkewWGF4MKdTtLPuKY35Y3jgCO8Z5Ua8LzTTo7jM0wS
IQgzHv2s8mIb+qZ597vMwnV7zyv+1vOZD3t4HW9i4x9w29HrmGum5CQJJyjR
jSwX/pCMWjrAH+seFWq24nRF1MZGN0tbmSbO0f5LcWkHOrlOtkwEH/d3fkKA
V+RnCKblto7YcwSiLdH6PKBjtnQ/NR3Y2GOdFWsYiPIu3juEWd0a9uNGvRgm
yKUCi71g1IEE9n2DCFqAiqD80znXWc2vvcy6VhK8R8mOciIhONeHJuddtT5d
xEuJGPyM0VzITGUlxDAvzbNcPpASWDMobliOfXPphM0w2FQgSU4aB7N/vW7c
6UNoTpCQZOeBOMBNtkNFKq4UWSpx6g+wxtZr5y/tRqdENNqgkp5MD5HMfWd5
fdxi3cLvLKd+7gRpVMNIw0kPT1HOvinWlwHuKk3wOynINHS2CttzKekH3ALH
ZCfHB/C4ip7YZc28WJlnc2gUyikFYtueNcLcWaDjKmys0gasKqnr4/vpth59
5G4agTVGECoEXW2YjpJCCgTTnwa4g9tWRfOMKnp/jRDuxqs1yCAfLUzbRk3z
lYcAka/pDwRJUhpsBMBwHd7OISqilIvmfNkOihVS14G5Ag7XM6NMMrEiejKQ
3e+wr5tOBJUqOcNfT4Ty8s45zfI4Vc76kkVKYMdsvP9sK6hyLDTGu0Ha1PR0
eMFf++GBqZGYC0tgY0ha5pIs5hIASlSy51+gYTyvDG3zbmvPRVcxByLXb2I0
D9UbR68AF4pRnFYszrM+FNFwxZFV8R9A4QnfrAw5xJU770x8gOmp1IzSKiCd
brsM84KLyxmXehLvByplVtfP6n7Wp8nEMZ3JrJ4qpgBUquPOusWLINIsVRms
Ed35SvQCsBiaoj0p3uOB9XLKOE8TQys8mE82/1y7+pGbb5IBElPt27amfASe
Q0VF7vwy/rPMoPutUXsH8hU48R6zkbhVbtXCRtIjT/t+xqL/nSXLycE3h275
l1/G4b0du7OHGQ2Qfdr4WmbCeI86YyfVdDZNLaXR5ne9//iIRIjsEaUn0SMJ
fBONFE0Roj5tGdYBJaiRKRDzX0CzZuGeVEFL+iXUfvu8GEkU5A7rAhSYFmYe
+rviqRQbZl3+5CgrOID7ndGYlqhOJ9fqYV05wGIOuantC1pY3eIgBkQrOieV
Rz34+f90yXkkerDN7/04a3s5kxd4DMnGLNpDfLZPboS5AnnoQtiE7c/DbOkG
xT9ftzAFYcYkUpHvzzXc7RlErgd2BROLjXhaXl/UPZ7vibegcznDjQKUH3JY
s1DVzfARNKP1w8b9Jv19JVXX+bg56fhmNdshtuNRtf/LMprRv3J60fmaT09m
0wClfGtpEqxakOv1bb1hkyXZWZaYp9y52rDbsmaO5PnCgkWNlHT4VJ6Oq+Cp
VJwLJbAZJ5odWR4MIMFAEPssyRyA7dxIH8Ii/zec6Ibv8MGEdHmqZG2sbH/u
RqaYbccLlAcZUh62oQ6XytfdM3EXB4U/ofoMD8C+js5hWNUTShJprwlpHe84
hh8+fYWW8Sjprdnhe1rOisoxDrcG/lkaO75VnLyPi6fIb9KcDwL1Hst3CfKj
DsfkCNz11zO/Ffcl5xxRpzU9tmvVICeVHF6+Z0cMX1ItpzNvWUhVLvM5gYGo
x3jgW4MJpmFT17AGMlWKpHOJ4J065icQmz+OCTi1BfCDpxKw2ZjtTibAmQNb
oMK/vhT5dWgP2XBeFS66NY63RsPNydxYNdfY7UHn4hAWDiltwkk19TqQBekI
9zAhQ/p4A5afOrt+o1O/MFtpMoDGQyeLGTGOmETK7Pp97qzNoP3DeXFEewSn
nGLQTfAIF7/AEDFyaC0x76/Qwsn0kmJCT7ONib9PcHdzzgjv0plVOL+uYp1S
x4fR3vAHjDff+H9kIyD666SY2K+0TMVfoPWPqtq6NMyCL38aGC32Z2qxWdxu
qupNjZ9dIANbMlr0E6SXy8HMjRMm48n3CK1UfKjk9tq35mOEsWGcAfgo7g5R
y+I8CwjONmBQsMZj3tMrBrAazsfKMwGd4KUixfq8JqVhzRE5W0Vd+4QJWwDT
B/OWFR6iFLgBPfAWNYY4r4Ib2pLhEJsjXRtxD4jRpIbn+DQANvJXNMwSP2v7
DasInpjJ+NE7V8OOwg5fMdUumauQOKKtje5D3vKKllDVwwqbsVuzl8noWttX
BlgK3dunO4sY2N36y0NZc5riCtaaHxVJ7/0b4YsQCrxuPqKVkPeLiRT5/83J
zk2UbjmUv41ka1Ol/G71WTkmkr9eHxWw+s4OOkLPgF96wpZgfIITP21lCaLv
FhWx3bfFcqdxjP3EX1tHDtKXDlIExjAQXy2FPjRFR4n0Qud3fafBt6C1UbmH
q9DO7NeSqXEbVol5QqIgImDkzsTDxt8WobkLO8VwAYBaCKBeelChEOaM8Jx5
K5ghSXrwCEjPXbecMZRX7IVxIHKf94iSvVquVdQVnW/7vzyeWAa308D+B2ov
ytLiN3IzorlF6yAnxrkg/3rOPdC7lANMNKvyg/Fc0LXY7/MRxSzjNKQv+sM8
Y04QKJ6GA7m9VBBuurn9G3zD81Q9UMNiFo3uILMgzgzgomBkB6xYkRp0P+6I
wExHd+lKvDQS6U9sZ2knLFT7q4w6X6vxxHJqklH+LUSMpMkWd9oPbAQBNgCP
tOA3MIxcBszYqQ3EZuPgrInZiRt5h15dGRBQmy5QY1IlSlB65XgHojso9gDL
2tYkcZ5CV8C4+npM2xZZVi2Ut3mQvYm4WBxh/ljtjYkz/7nZTqVp+9QGSENf
b7OXCzRwhonE0ztIEBvbsk+Xtr1her3fPTsR87AxuFxe7Tn59Ckn4ra2SsSf
zyLmATapVtanpJLB/ejgAoFJTLkF0co9Pf++SETDPWTQDABJxL3kzsUg7f01
h6kPQ89fObI3ltcmcxeTT4ZYS2XEO0KGQt2dAKCWtPmzwDwNuRhpXna9J13N
uSQsLuDAGYzbf6FPMfMfZKV/gfsFG1qBQwDl7A3Q3CWwzUTd0Rd5t9wZx7wu
f0IVjItfLNCMLkid4RTXN0v02hfyLV8zDgBGjUbs0A6R5sm/X87yxVf5XS0K
N9YUHPTzL2j6SIXxyM3+UE03CCcrLwSJ2WP5M/fKQa86+zA6NIpwEJ7j7kbk
I2CocZikrnQth2e1VthXmnkBvhH0I0EjZ8VDy+fgSx0zl153PLrewZMEhikS
Ze8o+ELPD5EBBJP3ldcu4kf7VZSagFgT7Zw6paB0T5bFBu9BIrLo8HDz9w+9
L1hLOgi2yxTib0PZupJz6p2oWvkwu5wKsW1UdG2CWh/j8JVHJN/lxJeCpelG
rSxlofXGBiwe4u1gkKp/ggASkPA4YmOxoQky3I/k/Z/O7oGLwWOIGj1mG6x2
Adll1BLSq60w/9oLp+Egconf4mirW2a06wG3sPqLIfclgWlGYJbeJ12TAinR
be6dRGfW8dai+X4xq2fhD8m+GpVFMSg0OvR9nxk84T8jesL+1OuZ4agW7EGO
VdRe1fw21pEtKAaaWt+FkENChvUO+pfYvgrj9m+DhFALMUWD2Va/wf5+b4+T
2bkNZhlzFyiLdH9dgGIYgehtngyFHL+DYzx/UQzQEjnXoCZ//fPwjQB3Y5jG
IIrMkH7DYVvBOdJXXEKmcoMRW/ShPUa9SLwppe8gP28BTmhGTxSQrSqvNTWa
5V65MtWWYPRww/2WE+q+5vQxfFrniUu+FT2xktiSFgUmQWyymujoKpJaHH8K
KsWu5c1QNwFMLseO9kQ/UzTaLTTHXJC1dQLC11eH4Us1K4vxd9q/Q/f0XlpX
j1KYlAzNrhRdSiYy+mkMDW0mXV5HLnXQ1n42Ycqw7bjv/e4ooARwMUDRNBEX
Ev/rwLg9snJZIMW2O0J80BSykMAIF+kUmhOkN9/FpwbKCbGnbUVmEKSywUcr
20fWQhvzjhcHg7sFUliUSwfhqpeehURqa8bI/a9KNsdk62NVG9uI80f8VV71
v/+ZmdOWIFoDi+ixmnEJoRq0YjhDBlmTOAJXhSra9OBEZE89EY9ZkZrZAF+C
m9JhBLM4MwCrkmOyKJSy4w+y/TSe1BMMpTZIYWVnzpgTSFuf309S2w7vGRyX
CroedgkZcGwwXHGoTdgj2IORZxSK6G56McKhJnWu7kRa5hLNLh5k6Ezl7Zmn
0mw4x2vJMUmLWz7ZWqQEO8hcMRQD08O8kpcBkIS9L8aY7Cue8Hp8QnbkIYdp
B0dm/Gh20E6aaBQWI0YoPC707qlfjjqEAzSsmIkVYwiUazFcO7lOl7nTNiHy
tobGNaFuRhajeWAUV34xT9y1C95klmpSGNiXZn344H4fbGzu2u7TluN++wYF
Og29SmGxWPjQqvUVfLsV8nclQ5CUU+y0iIRGtiJFRKbD4sWc+df8IfhLzHfH
9WGYyxhN7ixaj7b/fBOm1icG1zd1o8cvkC/pNPMdjAfd92CA5mtAORtbpRz5
IDpHjABcfVpbOcJT8CmVDymIUmtZD825cmmqpi4l+qy8ibI6MgEmXcs5p/s3
QLFt8ESvWCBPT+N2SsY1rF9zZkknvkyYhwcotLjW/gQHiyCaILPTkrJAW5B6
5wX+W0lIZD2u+ir3AhX8R/K+PRYMjXR4ifp8kFe1ojwqVBHywK6lnB0O+LIc
jEKHbip91GpMKiOwH7zNAQ+yjtgN7/xnajUZKSvPfHwJjsvIpPd/9fRGdhyQ
2UqgM8U9OohV9aEh8wWW3YFaTBnQhyU5fmq7RdDLlq2uxt+ngmE7JMhiJcey
sP6+fffkncVSYTYgZLUm8NdmmySqqzW3FswgOpDia+xRV5ua/d+nQ50otPiF
22IoahceDlGU+a8dbBeaSiXiGZBfxU94vsQePOFeNLHy3Ucy6kjpIjB0EBb8
3iqFe7+/qQhGDgib8MFyu/oVs/MH/g8/Vrp/ET0kCt5v5NgsooUDM6ppwn1U
0Y9Uvnp4N5q22ZnoC+cKsJHAitFLN0oboUnsS0iInkqiYgmS6y0OB7AS2DCw
QT/989Ogd7hM9ZEXgV65MqU2nfOKCJ737Js+urzWDxzSB2b2TVA4DL2hwhq2
xkvW8M6YJ5E/TEIcLhPmNepjWQAHjIfzSMemk0b8bpY/jOFxc2HubSQVIw9I
ABJBIyx92Hl+Lc+eEuf+PWjwvV0JsXbSusERx2dgiblbu19KnEt4T/SZxssE
IXVR2cB0RxR/ENgq/js2Df/M6BiVXt/FWL+HdqXuVSvuQp9vCtamRx+ZWT4V
ENZMB3yOjNiTyz/pWkKD7aCp0HsdnKqtu8NX5a6EqD+PMyEa/MlmXc0DUTdk
l8XNfE9dBRKZopgboz7ldfW5sMGaeyLHWu+QmbAKBxGRhLnRYNstNBSn4UW9
/t+8sGW0LRVMIyB7m3InftzXmLAuE+44F5iLHywfam55l8pNgtGPd4wSND0G
zoU7BSOcSI+UnSNWNhw2t31xdM2aLFTLo9ZW+ItPcQLrUlT83t5G6WNb5N2N
4Kt/EgpWKYTvx3IZfJXEX7aK1M/kstfvfRP6HLi0/dx3spH9cOCA2Q0CyEvh
i91m7oL/0CvhljXike8/hA6Qb6h/GcQ3rbskC5Zv4BHCW7Cid3Xv2UnHKIXa
TuDHKRJq7BSkMyGrXjDkryXtH6Cmdm0GvPgYSBXsaDggVtT74K3yqKFO3lHp
/pqUG+sELIDNQu3FOZFLGOdMUYfbPdunRp4/7Uv3vslAlc5wWEViNGyt4Crw
ER4FhGtnV0CaxJ6ztIa1otjQTPXnFXlCcR5M6qOjIFd9y4RQZw3P+4cpGcbv
t850FLfECzQpnDG12e5w/BiG45J7V2mRvBHscUDVbdlG6ud0ksumfB3Oq+sw
FsMnBOXcO8ytXd06mxN9wdcsa0Wh+hJ9pWJCn3UZeOykQVthyqy4F4qS5LcZ
Zq1qzTzFKdo2CjJzEiAQAQxo9LQd3VE6CwRSmdg0gqKQI2dw5thGI/6M0tB2
Ll6OT0YcExzptSeE6Lz72QxeO0lwktm4dqzEffkr0iLT1yk4m4Ct15Hr0mlR
CRphRMan5zxy6oMPx3FV3Q9wB0KBiKF/TMu+z2Cx/MKyPkZfXTW1NCdThcjl
ulIXuWSlOPFOyrJla3ONaDHqOXFAAFZ4+UCZyldN6Ll04Lkm7jfjpOW3aKKQ
3saJbpYQ0feDvd4eV68ezKvvRUCYBU31oYJF1QQJgNDi9Yk+ZI49E/SauD8K
QOnmIq3/Yk82NGSj/6zqL0n+wszOLMOC8zUoc1NdXbiLVaL1XCeGI+odrdhO
WYdqH4wzX+QApPlNpS18o6yJR6J0jHGe0ouGOaOX0aOOCOj2SENBDi6n23//
KH5gbl2iHF0SBYyaU56otMRDdULlO1EqVec4RtYC1dSuKIfsntLgKKtRRGQ1
QHLtapvHJce+Vf2+zxommOGDadCmcNieEa/m8WV023kfXpCpfrLdcG+iGFHq
SVK5rlqe5VcK5W5lxxC6/Jybw71DQ/bvhviJw5jasOFnLoXrkuvAO97IlI2g
YpRW1sR5XhjlkJoLp7orFPKPYzo7P7Hl8uwj6+dMulKD+m5/fy5zG8HJVa8d
c68vbiiUGOSMt9oNmmqwsd/5gq8IyQpjuw7tvUCiieX1q228Yey4KYldgIXR
Qx0K/efXJmV3AUA2jzeK4/UVw4ojtIgPoTY73A6kZuNtqHmilLGgedYX4dOx
kgNmU5t2xDQivx04VgCaNEUDbrwkFy8+EU+dsIA/EMiSeHPUCEGaSKCEvQQ4
byY9V3q1T5KB7UhUoqVNFAJAgYR/KqMwPOsDaoji5+k0moxaaju1V93GJ6zh
I0A5CzR8xff4Y2xWcpbHOth7888q5i33xlrMcKg3LQcjGXeq32nAAKSfLTHO
ehaYYGJY/i3DzNDBQzNx/UzcvE23bAhdpLvc/NGTAK2f1PnR7ykwr5TD1Ube
DjWVhxrWefCbUBadLmLwroPLJoWfH6eSKn3gEBmqf8KyB8jFCJWS5Ms2gzt6
b/+uhltACPx4oM/+j6naGrb+p764GrLH+hGZOzb1D63ln86sF47hjfBwAW+b
OQMGYxK49aPOcj7DHXuJiZg73EXRJ9xo1Do8erD/VFVwWnCpocHAAiUO+5gu
V/CzwIHIIHcXwr5tKUZUyjbpS8jX/W6X2Qi5ejVgU7slR2/zWZVCuuzNZI3j
RWtdXlwy8OwfrzUqne8LWxB26LFF3iyZ75XUGFJem8I5NDhNAIQf2ggoMnSQ
LVR/77CS58lZgLGkaOpw5nbGFzsWQ/uvf7y6nhB8DKWkawIo9adDmT1IB5JE
zet4O5QPv+G4FFtYbMOZYhJXebEG0qjdehgsDQij8lzbliBqcULQ7pkGfDBp
rB6IIfm5G0o0I3RMUZJMiGt13s5nJAXSoE/q1v6ErzZwB/wyzBSowHtepiWd
3c7Do4KLnF6IIfEGISP+WIvdpsmpC8vGef9diPmJZMxOnIbcZ8lqzTdHG7ak
Ld03vm+zeMtBkHWrASC5PQlAJ9GmrVjgXWryJA6N1/ZrFnGQABmhB6/Rfb2+
cdhZFMTgunB4z1JrcDMS+NMWBsJ0XtQcubwxQb+ELiUIYQvisPQ7i03PSVP6
1VcThJrQaNQ9ML/fKatguU6R5V0RJvKA70FpftIYz5APelUh+sRS5QbVvpYy
9RBM2Y7Y2wRq5Oa+xmFdLduupX4t9vOAdkdIS1mJeWzBalVZ+HJLiSFNiSWp
kHFqrkfgMZzP1U9c1cuekJZgfXEDySbp3e2nKtH1jp/bP+luUr/awKQYApf6
kAkJ+dFl+7Ym0IXsAh4+u8lxKWCkX75H6I7pqh3aoZE2vZydqmXQZA2sXrMv
Mbs14uFZZr+TI/oSXt43TFAXMgnzHztZkldDlCXFa4LN1xeDYXVA4QuKhlS0
lFLezRSL6kzJx8lPAioUA1vIPzBi9SyQ2SDNRUim4r+gn94msJY57FeWiagX
93MkLXGb35GEK4GW4OFuB5EiQVn1fSI4hU5cElUBQ8zuo1jxHga8ZJGWV2QP
HCa0NgtQdOHlQ9r/PITVyMt7BHdLG3yHHRqO+bqJru6npFBenmoG0QyrL3gg
+nptR5G8ZgWecnCm16XVRexgVrREqhA9DQjWenqgBeMJfY26y4AVXPHz3Njt
P28MFQe8eS2T+sRH+ZF2pjL/4QvvgY4W+0DjWHEY4PdvmC7cYfhKQp5l/MTt
pdj/7AUhn0KvhZBLzqQlTaD7GzZl7vID9naNZcyuGfyDEkr2CmrFGRKf3z99
nsLJ4EtSH3P0PfT7bHKP8D1lTPC3S4XnRBB9NvdFSx3PDqfxOp0aJIUD+q9K
G3qfultod7G6LVM4T6qMETjZLPAAKBUAdK9QuqaNDm8Um3JoY9jNLL8isNSa
1h9fwmUWv0TQnJFee8z6Wc3PS3meU994JyeY0yvWrxPZs9VFS9DtrZkKAW17
9fKS0Eg9YQ1zRCNyHCTWtILvUgo0nncMEVuw3yMMXCXYSirqypuy4Vt261f0
rciOj/rkLdG1st7VdIKvTUNge4V8ZVIi+PLe++s6W9avFxkwQLAjzldc7c+M
j9vndcFC/SeJTo+FYfjFCcT4B3k8YYlSCFLECyXPVCxS/IOKmIUCCImozD/+
enNVrdGWrGN5UXbewfcZ7SWyN5fMBvt1bZ2UL8oFOyL7P1sP3MqXV9mHN6oA
OVEsI7kBlfMsvnitxYiP0Nc5IdF65/lbWhwvctDW6jGtoFw/OOXuR74WEbxP
lC8j1hwKHKZSti0w+W/gyrIzhH7L8MZ9wFHquHZ93VDAeMEmLq2ox+RtN0Db
82DZpBh46cm4UbQJdrpUGxh2xCSlNaDX1KR6OCQTmf9/3dx1z1kJRoTdLtWa
J54uN57cbklUOz8BUKb/6mWzMKQgc02Qc0vJ+M2iL4uwv2uSs4cYJAeIn3PJ
cu8/qgpXVCFRqrE7ozTZElxPXMzJW4dBF+xiz7omD0y0INk+aFWXv42MxDGM
f8z1mEzBsa4I/m0cBrjjS3Ex+PYz66xNkI5/sQ8mqYjyLrNAyUPvL0e8CMcL
tRNP8wLVaVtRuaBfvfXsnZpTIaQ2OsdirrkRUpDzzErFwBUDOJZ6bG1N/5oD
A5wc4aQS8PwlK408mBeAKLmjNHu6H3KWbZ57b8BAC05Rds8x/eHfq7Kpo6co
+DZ1YxlWqVZK4qjdIrRuonTq7A12Iu3MT/c23thluC9ujupeakVyjkAzZ1pV
eJ4UoPw44iLIvJh6/0W/i5y9btsLDOapyZM7/sMpTMeBDJnnkwcKJ0QY1Yds
IciiYJ9H6K7YNfF5+dzPAOUye388YKoeKnrMTMZ1y/HzpwTbN2w+5zF0uo9l
0VsfxVUzE5hWT5ineZfKqnmFN3tGXTFy7C8QDrlmrJ8vRT5JZxY1QzpB5afl
55CYvCVZuKMcK25rls+1rG1QQDglEuYKcQLtrAXNokvy5k7qheSLa1SqH9mr
vW7TFm99uy9nqjilDH0CVpHY9du5LuA1bS38OwiYuwjyca8lMeDQ1aqrWTZn
OVvW9QxrCCzwUjgii0ZToVSpHBP5/FH6UriA7raGCd5KHnix7Kem4nXwrQBi
PKpME71586Ma5aZDjmteoXBH5k1OftCaWcwb0egtHR8hq4u8cWGMuL5+W/x/
qPVqHlmYX3p8ey4FGUGHR+i1PfgjH+NvlyPs0ZZIjtCs/BZRciAjzzm9FGby
askxFmWwNaAeW39Be4hfVYgEdSsiN9+cgV508tm8rQ9DnEoahv2SR0Nzn6M/
IgkuPh7vy5DrhdrwS0hKC0olCb/mPx2yWhm2UCQ9AVKm6LTvL6Dgv3mB5SGD
HNS7w6cMRuTbViiEm9Z9XC5YEff4eO7QQp7BzZsynDQkZ1NF3f2TnvFhrN5n
Y0CWDAdjAakeTOLhpWXQ/VCdI3Hycr6tlbmu5/GER78QJEzHHwS/BtZIpEzS
2WPa/ksrwrLo+27J3VjZUWI6rJevVbg2DRQfrl1FLG4p3xpS7QxyuH8LOGHy
chsIqxRgylm2O5QX4UWZWfCzgT04nUeqbG1c/YajeeHSARxptaZUmon4B3OS
Z261+7YLjAipYuow0xclnXR5S2FOIjLvGXqEWkbag46R5D/w64nfi1kOohSk
cj67Zu2wH5rhEIt0nYFcIUz3nEAjqo1eLdzX3eJAQEDMAPwBZZD/98sP+2Kj
amw25xTfg10qxZiembfgvg109xaUk8rtKcHu2qQiLfLF6T37jw7a5FVvcMje
ZmlBkY6QNLCDnpg5DDz18jwv3LqCWFfyqt+clSele2CU8PjTFODehj6W0oP2
G9A5aiSjZCC2dy6M1MQasx0Xse3J/ZyiRExig2KdAwQUGBddzCKwaY51MZW7
2Y0920NBsjFgi3THdOKBg0v/0dxEHREV1RaeOLvLKhSNw87oQRa3gUzRKxbi
tEvfCnjTyZRjs0BICPG3tdJB4QfWVbS2Mjbitf4/og/x7WC2gOSzuM9uvc/s
3CbvbaPJwVhU5+U9irTTNDyDKuvZSJ91rV7Jj4XaYvk9HNNUQd+vk5dsbwTM
LT6pJOjJBw9iW9oChFibu9BLI1zc89UZJsK/yOb0YXfmZhz+j8QcS7Qc5Flg
/xJajoVr8rbLYMnRaWiqcVJ9U5NO4rEEgMEmhQQQZlaamLkCtH/Af9ijIzbf
wvKA13Fm/68S5NL0xRc+3Q+VY4PXyeF9j6Oqm/0w0Toqp4hh+fy24z0UFjgd
IZ6oYKp4vURgL3iIWjYAWGxyzN03YxmckdIYSfw3sWIx+eFrl8CYiFDZHb6F
20tNXjqCK/KPJE4n5r8mWevipUrSkFt51N2yr67dD49iPbZ3GQ+uFHnCsqUg
KTxcHxWNSgCFBZEWFL0o2O2FeD5JJ5JcuvaTYiYAsJBJMsF1Xs6jqvaJwofz
FDgz0fSSlKzuGkIk0N4w1WZ8z0ix6WM0oqvNPDfRVrVT1G09ZCk6L4cutZss
wsGlX5+7+0mp96MC5N+jPAtEZfp4tQyEWJD1IETMpXenEi0gtH0NX6PB7Oq9
OrC1+YJfp857hg1TnMAnqloLuVNObR+P7xoaXKsgxwWtydCcNe+FXLY6viww
BgMINMTFnTWn48uKxDfPSHfV72xGYG7HI60W1aHF+jpErnyeAUZ+FhIhtmdV
k9jvWQhpVvbNWgsflgoUCMk7ntEVH+IKy9pF4VKBYOaiMrbXLtmmqIo5RlRV
p+Mh56btEjRGf9lasOvoHs/ZExNbg3NGL+77xmgN6Y+ZoMxrrGN2EU7rS9AL
89eYoufD3+CZU8sFf+3omOZFS2ehV9WZYRXX1yF2zoP2V6ic5miYDk4vUO52
SPpnWt8hjiq1BaIX+ijv9HLzKzie8udUJhn6Kgjvx21YZ93dW+tmUMulat5K
AIg9rN2pgP+92lMBN13CdA0FZ0Z4PAQDj3YH0no43Z124o3Hq7ue212hZNOI
pldhzVXjmmTwvpHp7dqXBUN3jUsP6E7xc1+jl4ObI0JzSst3wTcA0brWNPlV
R3PdHrr+ROREi4pk10TBWnokPgYMq4+DYVGbKpf86eJ/6K555RJpktjA7sru
jvuukMpSi0ZPsV8bVM1FgQZDUiiHe6vzqm41QkgDWQXxQ6kFJ+T81Z8nId6R
9asCTRMKqBeDVk/Bop3l97OZNK/PJUCx6BT3cIQ+yF3q9p12zMwHX+0Wiahn
A83ZfH0RXB+eooXa4gWGPwqdcIuRXpc9bgHSGURzpCZIqh65a3B3nfsZXIKk
oOyfJmhB+Oh7SB6yx8/LBxmO0vFb1K33ixQ4XnhdosrYF80/EOjOOkhOCxR4
QjjXgEyElCzPh6EHW0d0c5tRmOpcGcG0dSrIur+TkVko4g5bMpI+LhPwqc/5
EPpQxta93OV1CzRFSLFzqUbwts1v7Nsh37phuuJS77uTLS19yo83y/bnezsx
trQqnlCK2ntsQ8EK5W+/LKv6WCcT4tWxWVqILM/ARLvnxQPhF4KXz/mB8ASm
BQdOeyUg+FgfghkOA7Kccppio/G6qmMoveTRIQrR2lTm7ra3ql5H/Ef2b22E
Uww7A5v+5kOQa5ZLpkqAx9j7YRlaBqq0pyyhP1NOAe6+YYZ3Bgy1tjT6c+tq
tC3nc7Cz9WYLlAGRN+w7wWHUtibOSeq1xKon9ExXuh3QkpYA+LOxdqknE2TS
VZJbPTacimdtIogBDZMVZ/oR0oYTwMg3ZU8PPvipIj2JLG+Y3k+A3Ik/Smc5
QnG94c/lzlAB4i2o2CUbqvf0Bb5AOj8riQokuNhwPxjrIwjQYs6Y9EsgOUQe
5EaVJHYLShVo4f5IFY2qjWIXvYT/O/s6sxX6qMFhLtoF+vTh73wK+YvmVhLO
WAzeAvlvFIhWb+WMnoYpZtkVOafIB5tgEzz1W2Pztlx9yWsbTr5ddNu7Rkcn
5J2cTnXVKtaVtMB4C08mnpwvl9UU8F9H99Hu5+9nO+YMAgO1iDFX/nUVP8NM
W8a+o5uJLgM9t4g/A+tzsrzYMu6aBITzjM+6lAjCn00LQgKUQwX0Db8lAfXK
lJj6BKbuy/FkRLXSUhykWF3FolvytlGsfOTA3nR9RsKPixQormvI5Tsyx95s
KOLOaDeE/VEF3yhpzLBJN+3TSO8O8HQAGAEs2s/PBAA2aLDrleSSCCy899Nm
5jLnMb3mR5EWkBHcg190zab9chSHtY2ShYUrgDlC4hVXymLgKglhdjuTm9MZ
YAb3q26u6cTWaB3CnMRD10FZ0LcI7O1zgdu7MafKuRIswsSSD/B1qzFbS1sD
H9u0Z3TRuG+jVrB0SV2SLbQDMdIs7Pf9KYwRhu1V8/MCUVmcWMHFZcmKdhUj
q2uzsqyFYIEvZ4PgrnDU1FkvVcKQoi0uXpj4NiARGo3MqZQklWnX3G6IJPqH
SlL3qZJEmTVu8BfGKQ4KHFelpFT8itDp2ifXkCEMOdvIS6Hb5LO0SdM+zht9
pQfimKprhw6GQD4nV3LsAkAGyuiZrdWNJ7+AclPjU6vSU+bHvm7qLwLY01aC
Go/dSvruv3Tpnu8Tr4UkUk2VjbMZR9hCFvmGh/ICO/9YgAD6QN+1ME6PucLw
+fIO8SwVLB38BgulqUXjAuDtkYTv0jjnKRjVctNjdDJkdqlE9BKl9PYMTWS+
0OAJazcug5221da0sCbSxvjMtoce8xF3t6iTCndxE9Raa1gseL2sCP6jF+bC
Lanb8bwMTd1FKsdcQ3jGD8m4TqBcSLL2V3TYYp9nSf1Vq+vEA+39ObRfvK+x
sDM4QQle8BPvXz2dJOZxhPH7MZ+OpQ2rc7sTI86V+eu/88KnhUDsKiT0DKeA
OimYmdzRf7N9J2DtFMe9DVHtrzjAynphSR88srnUYKoO7rzPi4Dsx6ugdy7V
QHRJrgFn7MNKf6X7LGIV4oy3o2x/8XzaDCIcgzqnZhicl+7t1Xj5dFnvk6Hc
pd9cfbXpySyaV6hLz82Fu5gpQvcyPx4sf6w64uHW5hkMUbWGFCu7Es+Llbgq
p1TqDY/JJHmmMjFp4g6DfPlS1eD1SEhvj8XCWTV6cO0VKwHE9MIj6qsWDqwC
X5jW6tD2nR0x/1PBTBpgpJWQasHx78c7Do9i5nK3ZVI9VJAbhFEyYi9lP8Z0
sazhzWBjU8ODLTua7rrbvvCaP8Izj40YE7QROVuQdzREXy2lSHM8K4OReJQ8
0yWbFGCtg7AVGOBTjDcGHYC2yZS4Lfh86axxj7Y24ET3KjFHKvY2C2HGPGIT
5c9QHLTllywuXOByJd94NyizizxovyyUR1/ZiFBpSaxDYTK5P2v18wYW1KY/
k27aHqH4QrPHQZmKHV1Gnfilxa2jPI6g2lwQsIRwJS9c5jVHS60+tb8RwsHP
SlfuMao+cUeFjWVZdIqAVMn4lkfC/AqnJbuNpHSAOnSWgoxzy58BhWiTXcQ0
YrwH4B5eUhTbQd9cVK0t1usVO1xqrfobp9zz2pR9h7Y1XbwlvAPi8Pz4xeZ1
B1SYL+am9uUGOiLxriZCay5gPVhDkjl265ZinQFZFcbYKDj0zYkHFfOplXrk
V5Y/2eGruCVI1sh41fYI9tuim/35rVZ+GLJ1CR0zLFz6OGbqlSrMmxN3PMF6
HDQ4xlCQ84/Yhsu1GzzIaWxVPmWooTdiZeUB93mhVfcCmuyhfBCOm19COs4i
mx3jVQZqldsJZx1UPuKfuaIQRiCmmg62IXQRkLo8NauMxdDu6eSH/IdKx4xj
8qHl2FoCE92jbn81RgsfZ4ZNQeKJml7fmZ6+dWSkfVD5rLTekStgZSJtuN1F
zXZWIMjByP3q6UNA5aIT6Icrw0Nu67H5LKfaeploX1WPe7cYt+wWzYl2dmHM
TJyJygx6EYVEOYZZKoMDywsE8yAyBNfUYFN3m4gLmvMUBRT46C5+xVA4gAUc
9a0bRGKuw3E154mIhayMX3hzm1FOTDT6mPcDhHvAW6YORuVt1R1hMbx68/Av
nDzmnzh1f2sbSeKPw8b84jaNpKdOrUjPlLAzx8ESTDly/VM2Noi71cSPs243
MLX4E5/zRseq4CnqVJ5KXbqOtV0zEkpRjpsNrTJasQHGkN2ZsNmUcI11c9bA
VqWaHeMX9uiWona+dEd82c7mEe7jkwt7mWxNA7byuKZlptsdEo9JRRJkcMGD
0hVS+k9vTT+kZ+7zgflKAuydjR0oH864WTYPxVzIzsq3A+VbCXyzKNZaeY8c
ppbp8CkszEVxdTGWy7t0v1MYwF6HIPlnE8m2zf9aVnFbAFh7Ifrd0xizJimb
2vGImhLxIfdWVJmYnNt5P18LzjNaI5qTMAoIqiSHfp/j2J8wC8nyesrphpw4
is5+lQhAoj91Q1m1VBFfBonMf05D/lgcQsByDGzWmN0vsno4NZc1gnsFKCXH
hN4Kt8a+/iJwYFTspaq84Mvj2HxvCtycXfQpChZ3KenmaElwGukbSiBjBHhE
z17Ab6q8BaqILV4usacCZTOl3bNOIHcgOhzZwU02ptJuzzMfN0hiG4Z1mmSd
a6wyXzbP8UqzXYRkKMVVgaVvkudmslQ6OODNn+yokObb0Sg1mUP2HMGYwVjN
ni5bHbg3viKzYfvtt78ZzSivhUsFYzq/PQBwQjgEd6dBrDzL3Qzo/7WL+ek6
bqsnx9ZlPaJjXYJGMqSadt4FbpzklVDmx4+qQprxKQzHL22pdc/01Fuw4qvy
p4/kK8O45FeIIekFDcdTA+lxxCfcfJPbxWegbjq4PO4MGJKf4n3c47ZhhE4f
EqgZkRo0gAn4ZzGbHEANmDRMRGRQh7TR0e6htrrsUkxs9nEOapufNu65HCbc
zM3sh9nlAmtHSoKk0j1GIjrwwmfylhTevm6GIlunQbrJkgs/XkIBFYhy2YbG
WPYdDyixbbrfDHRzTAD2mqQDPwyXRwjWNTBfwuLWGaBGMCsaHOFAPS+A6qc2
E8UneEFlwUNuwQmFEq2hGfRrW3Aa3RNviNIzsTWAsXALgzbIFGR9zQ9Pl0NG
LC1PYE2+G3eOEDdEpoOOXkUFvZJufL7wVgm5nHeWnd9TALVA0p9KUAmpvg0n
yceONMHRwvL6chLyqCtLCu3OmjiCTDMPb9Zz2r7Wdjbxrol4t9yAs8l/ZFLG
P5kX2RnYBWQxE0YF6N9mJkN/8IlYsMimpTIWi4aoOBVkGyPF8JjQTERDzpES
+ltGDsv8ibkn3mUw5Da1R+y+3azw8A9gwlG5dtpU9vfRnw5TdGW44MVdph4O
Rq9gzm8vtUnIFhreTQsnuk1fTUeVJZJtq6QnN7kf3bgLQXKvmwjU5VjV9Zpr
9U5L7kHy9QIAv+5ceNTtGBbPs39o71n7vqwXeD3Fb2vwdjUpDgLmXlhF0Py2
EUsbopvwt5DrO9yXGl7Xris4ZS+0yERidNNAaXW1A7ymTANvYBXisGOYT+gP
gJkujdYavRrRhjFcRJS1g/Mj3uLJVAkHrYo24dipvtkRNeNiMh7SPTpXCaDj
ngnhTsNEmD745KDAXjXq00JHKRWF2+i0FU+jwp+P8JeBjIy+dnJeU0qnPT8r
m64qn5fCRK7BnGF0+y3HTJuCyGaJIKvV0x1ORdb8QSqYjFZZ7MdHYv+hvPAV
CoUtxvzgGtokVtEhyAbVwp13cPlNJRldI2l/TnfIqAcZUsDiqsxiCw/YHhcu
WeTPpDQSFIIWBZeWISMYa+H+WO5MpxGEq1FVdrnPEWIquMBB4qG0bK2UITpI
DaqPQdyEpsss0kcZZKXjVTQEAciicVxT1jiTOZ7gt3sXDXo/bCXy2WyqnBEe
lJxQ+Z5tPbo3kXR8shOgJ0IlI8fhNrs+8/fqYnwLbGjUNJuGsQjzxatKu5IJ
NP9jTj938dhO5Ty06JI5Kum/C4lV4OnbGz1w18NyJ43V+GXkkOHRVe0UbUod
xfdEizkFRyNJoiurpVe128N00qtoev7z4BFcKlW3EyXC1Rqa3gqF+TDxPTSm
liO+YCdJErm9i6p/cr6UGR58OIfKBTTcTMxFIi/08RpxlgYJOG3rKhFd/nFp
oGOiDOOGNHkHruGcRXTB1ctUThELgNsn5jMnMwMGrGZe+V/FfEt6i/bIVghx
sFLdqBtvy8QmS6wy/pMAJxu1tvPpb953geAzxdsFATDG/gdD3pkRI+Kx+gR5
Hs8IaamYABEbIoDruwf0m8K1EyAhL/vC7zrt06jHeGdJa8OBbyHOTdL7zmPO
5flJ2tRDUxEB2wd/39a8hgRFk8hNd8UVsWKCgMMPv0rn6goTc8V9sV+rrZcb
6Z8pmbw+pb9ztvUkZSjbzXXgF60fy1EJwsrxu6pJF3a5lzIfGbv6+l3C6FAO
AtG1S3/ctwQAPz/ukiJgbQqA8QyenAgGnabjduT2FjFLEDr5BMLu5YfpTJLL
fF6sWvPlikx1WngYHUEkk2aufkBGqzHwrpeeIgpKnQnOtnI63TejfgceQ0vh
HaOkGwnAuuf1viA4ePtQBeJND13UjXiPU1vAiV43r10vAtSylhiD27I402Ah
fJaWep0QTP8yXKmxk3kkoHeng9r54MLBHgymPIOWHhXD5k2kyVPpLKwZchzs
xIPa1a3HtUk2MUFYtuYY1WjS7WNP69CXylUjv2SFifsoapQukoZ1RcqYqi1F
PweJmFn8W9NMiXvowT9mbJsDbBCTO1XKHURG7U3wHX1/az7r8fIiOXpyMsDh
QQBpVwlxC/DuMwbTximITv0Q0lEDiaS27dECnhu7ec/uR6p7ftdbf7Lw3YS9
FehIbOI0f0kW7vskh+dMPwjAHCu2SiNOFk06lVHfRC1E+UgkFTg5P3soJQ0e
KwLB0QLqTiQ4H3wdLUJ4tap/KwqhrdhfuQFmHp38xXyB7PDjf9Yg5lZcCNJr
W0pd9btUTSGCHn4Kbo3rtQ2bAG9q7RSw0QsodQw6GHWLYpPzlaECmLIhjHdz
bJilV9I26o+eIFxaoL/sm8XzA5lr98M1ghSw2ZH9L3/E92yxxZfftnqvIp9j
ofCkhc9qkk1rYz2EzFybgJx2ET9LcAYaab6SJZx0dh26+ORoU1HqGKKv6qJq
xJFoKCilqFQXINOr5Z+VpGMz+aonfMSl9wVxUdtIdb8W24J95Q9DbZHx5qEA
8sc2LQrZdcEkpeF27sHUBa3kfpm+WNoTwHYsv3xlc9ShsxL36yj1uc9vTQnc
3VJtOnX466pceTH8f438GWmmVnUMde15N0TY9sZTNXtBcGro93nJJ5P60HOu
muVNz9FP0mqYyRD/+JVUy1Ev7nVuVCUlEhSJs9YfbqE5LI4ifQdKvUGqPY69
yZC2XdfI8LptOow5vKltQqhpsTa5IF16v98C0oqFgKJ8EbR9fPL7WM/f/+qF
BIsbR05s2aA3qWK8umT6Pnlq4Rr7T/l1FlzLCQ5fYwx05RIjPhdQs/LxgPAx
OZmEyva+Ki9zFhGop6/r/Qp6U0UHXC0CgCFat1u/55ASITdPzilSWi2k99bo
pWS26EJ9S5zoZj7t6QMCA8PhyCMdtBlQjnKxq/aWMCsSsdJcF/nreJol0sP7
JAgG/Lwuq4I/ltMuu9CSHN3Chn6DRGwIeL75MuOwH1S4/a321s6KdrODQk0l
zBlFiN2zC5yckkx2khaRS+cjgwF1K1AWOsX2P48U+eckNM6EbFUS/QEmuSP1
sSpXpzUS/IVGLQ62S6VmQ3904sih2/xyD94pEcZjlPL7KMTy5nL/ulEo5W50
xPf5d+GkFPWiVb2H5Y1n33iUSZFxe6KyHdK7aTn94MYnCHxc6oo2RLN5jjct
wTgyVRaemJ16iX0HuYwFE0fThnKgKcfAoy5QYFRyRpdEWyQtd1iX7MkC8lSs
H0eqwv65g1aA7618aZzimK/BG+UX/TxvIdRqeS84V7ZKu5pndfVx5bIWsXlr
w/oq9BVHrXEIGKqpCj+S0q5BC8EryNbxd6pkMnfOGwFaNn7cSOxqUyjhWLfd
xwPPdNsKyxEHlg4SOLDiVPEkmY4xleqVPRNZVFbqs+i0qVJeTmh/39W79uH0
UoB156WxFMmUn+rpJ0yR0kALMASGXASy8jbS1J+bZuKROzDXlD2IpHvTFTnF
POOzuwR7/kVg1fOp1/LqU06pZgC4f7NtvUOq5O4hzhEl9y7kOiNzIglDr2V0
3BMABqoP6L1+74fa8i/VXOPXp8BA22AVYNS/fhSjXWZVNTnCHtaRrbUeeAX/
7mLPnL2MFU1Syud1yjbgWZP0snJrrIzcObk9jdq+hN/cN6AIWD+FHMd5xkQe
W57rQP6E/qiXoSW4c9rnxFBjSLE4ihTSTF5kAVk1i3U8y/l7XPsdNSIeYn7s
6zuEtTMSwzbtDcH9z00vKD0+DAc8o6l+Hlh67TWEQkx4kKh3jqZbCfTR2Dnw
fffTAOqZdTOoMPQgztchGjzpkefbTR7KwOchoURMmBdZI3j7VdNszl1Or+L4
MWBBCVNu7kXJGSxGvINCfUAPeZoeekSugqmxBSyi554R3zoJIwnP9NyvMbuY
2vcKxHP6TjU4Mrn46B+Aqb/crk5KUWVd/atCAYKk0DRwuvspKY2V4QcOXZXp
FfD2b+Yft5qQUrTIB4W+9V9LeEycxv2eaebN+YUsAMHaoepiTKFdpKTRanqJ
z4qj81NAgZ4ovKAVb1JLM6PkEr7LnKABuWNchv6ksMyBeh5Mvb6odfD3txes
1sVy9LR3BKAGpS+87MPc0iW7tD1IxEcBQkaKfZ1+cqtLEe17boc0AMbHtW2A
EABi+YEFaeb5ScsAfzHqlfsPfgkQI8UitUa/qxZHfIcHJZHfZvipiUEvMUwx
Us9J8M53Vi2oqJ2dlvvDSUH1KoKgvaAzlYDG5FR/7Sx43oOyVKhQ5+68DvrM
zmhLbkPDM9a0RAaUkLluENidrtfOmf1VDtCDlwb/e8ybSFhQfoyPgvW09Pep
lia8PPJ3sDUJHKw3M5zoTfzVBP/cZArio79KrG4y7bVIGcaoSjVH9KUU35Cg
VMSEkLmf0IQha/j5P/qAZKUUZ8KqjVUbM/AMTtlFiuuTW/e5tcOAYHk/sQNF
Ia0N/sADoOe0zbPZCu+P0QnFSF1mKvnCZaGUtB7zSrKDqOPAR+UbD2vBcVR0
WWtyutYdZiaUZmMRId5cf0etWevH/XNhKgTyf7saPG7KFaNwoR+C/nsVBy/9
7/S3a2ysaX23pCzdJACSnIDXjvqCC0lBXoSlufG9NbstSN4WgxJt+VrIf0AV
wGWJcrXe2jB9lBGzfnuwMX9JA4122M+rL6MM6wbL4vHwgw8+LBrilP2/93EX
klsDk+W993fGs5S/1kmlj8fyjtaEsXtQ96M1EdKr9pFNAX1wRJUPv5ajyCy3
uOE0/E1gGJyAYAnFTdVc7B4JFJbZ1bzkkEGIZ3tsT/8XF7vxQIrg3TLx9aE8
2iJfP3XlT0OFFWsZM3a5SqnlgNKTp+1slSOGMYCiI/S17FUjYojalosRyGeX
ATTKZAK227Tf90h8KOkFD2Jg8GeWCejZfgKKRw4y2bN91WBvWfpxTpxK3gHb
C+ZCYJBjwFWE3juO0JA1+yDWCQ/CguPHP53vizJXa3E5rMd0UPlr6H28MwVZ
AvshEAHBd1P3jjriqO+khhI0MOmSrwfSAv66qoQRWOE0ZOBYRma8rPTtgCVv
FIIVxKvCEpSue7Xy4I9gBUgJN8mUiDr4/5/8IR2vvBtlCoN7biwfH7L921B0
I+1kMDDN/c9SsGHP7c+Ci3gzursAR6lpQJUCSv8siAlXlqYc+0QVXDtJOfws
e9t43XczrtjZTH0VdF6GgyGHFu+C/UzoTx0hRMwTGyym9ryOjpdY8Nro+hTV
uxGOgSUJ5yoo5lEQhoQU5QNfY4+NPhTNvYjGQgVtRWka+lIuUg958g5tuJ8N
OfSEXmtNDA52o1BmpHudQ/Nf32Np5WcJc8tJlDyqvRzzrXSOzXjoxowwRq9m
0WGU2VVZajyoZzvOUmE3jmy9hmbRqP64+BLPpzjQxKDK+AB24BASNn7KzVA5
NEM5ZCXszCxtgkkG0WFt83jKg8XMDS21U0xn26XPGPmInSrBorFaAZr3r4XA
9RE8bzNzYKEFbRANIUn2bygXg6zq/2zhF6sXvv3AEjfEekvw4ojEzGaiYYtt
dvLqtbaXoAPIz8R3FqfWUfnE+Kakfnvo7dKHjJkUpWprSeMgfTaNkHL2PH1e
YIE+X9AZdU9k7JmZ7fDbYL/b2yeTuMCN5uDRF3M+5CaSd5Sxkpz68NqXBVam
GRp3Wa5hIMxoE9bw9wmDN6KPmRuQ6IKb/6AO+bOw7fqrQQDd+U74Q1htzrXE
0Je6Zf4BC0+hASIs7eGMUpucasmPBV0ZxNI1kySsxQddrQeQCPmWXp2FGZi3
bssEw8nEtf8Dhx4kowsR942dvnVYTvwNEIewLhi5PG7YOKwy+qCpF1MN3nUm
TyZylsurU62rXeDT3j/YjsKRZE9zPiv+A71dGkCwOy7qUme2jkgC4xPebfvi
0/slRxW8EGRAjjdnO4wh2uEN6oiD0LPeLr7H1Tt0LtTzWiUscIHjp+q25neg
gyVagFhbZdAjdLW8KI3+kkJ0LhXYp18DkHxsyzohxdWLsp39RKho+vgLHhod
e9NuWe/Wuhgx1twT+ngEnSk0ABDb4kmlINsBvRl+chYmVKxu5ab85Vn966+3
XQSGdI+VjmjY+lm2GJzAfEmz/RBMukG6uqyflQ1w4hKmhYRyJlDN4KfaX0LJ
sbAlLVLSgVWnWFuUJ9oENILIxIKpkYzV8u1Sqapa3hYBD2vvx10NEBgHIsez
Xh6xP/aQPQ0Oh3O1h/EbXPBKU0XH31fP4nupMllvRwKPw8nTZ0YwZefNiFtW
MQhupwTXVSRgQOCqUm7C5BXg9EkgbdZvUR8XU4L8SKe9+U7vJQ3QvdQF0i++
Oequj6x/N2PEfqpntQOKxzxkJyHt010Kap1g+DegSDG21BKLzScd8CEW5XTv
1wTV4aPM29/K0uJcACDiHFQS7uCXwdH9C1dutTWDipbox70wImsItpANyQmC
uQN6Zp4K3hybZMoaQCiyacolP0y+TnsagPFOKMVBpgyWNZvKxtVJAHwUQwyX
adjZf0VNB2GnCPkQ95xtgDKTzTK6tI+cZabAHE0Ys7MCoJ5APJSeieJCdTBd
KxKaV+fIUOObN7qPrgg4pQAKVWw2O90hTLbpkzJftMXSYrXH/Nx93DjIGrh2
WGwairImp9P/YEJLoRofBudTgSruFfOJQjkC7S/rOYrwTNoHNENaWCiWwA2L
1UbzY+5uzpxvAoUmzJbA4JLZ7HRlcWzScG/xs9MzUsSUceoKAj5BJj4b+6S2
1HZ/ib1UojjcdJ3VJjUPdEu2gu70xqAdKuVA7fhxEZQtkxRqtR1+5F4RHwvK
O3nCKHOXJ9x6mNFeD53KryKR7ILRyu/XHP4vncZHotHEHSOUph1rSXKCbBNt
gUwlbSRLQXYiTCZo6DilAQyvasM2vkX+oEFDa7VGIUzp7R8Ic8OJX2PGpZYP
EBqCdgh/ZaetR6BeLlXswzqIqRASP7zWEMf7YH5sBGj5xW6M26xNSxi2jJUV
98Hk2CUTjtwChSEc4sPApfpz3OzksH03fFErCSVDZeFwhe7R+FIpL3+S+xom
26mjfPoCNsnEBXK6RtmrcJfwklXKd3Tf6l3dmXY09jSGKTCAsFdnx8XTBfL8
X/fRNe5PwwurT2Iz/VM8zylMj46GyUx1/yBV+liwIaGQvIMj3UaBKGVv5dWF
dFVkjP0kBbQcGYsZWYdhDTXR9mT2ajUzrlgPvM5+JX9pQY6z/HlyEiur+S5C
3mLae2+WGv6ZWX5ElXw/0jiX0EzXmUmCaTePGYELRWEjh8i7Pm0FmaosXcVi
v9DfpKbOTbcZrlaQEBO5MvLo0xEPJhZEjO+GcchokMpdUlF1/ZgxkFXUVxWi
HIaod/9zNjjn20FTs2WGot1wm6gt1kHSXuI/wLS8ThIE7NU0mWZwalIq2A2j
WKe/JHMn3sv3E3lQbQx1apnwwmq4UNiLxfYVml8p53dSGPBzWVw02WzQ1sUo
/yehDuCDjZgDDLQb1jXq17otsBWJNwvrqcFVhHqFs+I8Gq2mW3LM7w59CjJy
e8jggDaYoWGKLRZweuMc6Thc1Vg0m8sNwMpv/jpYJA52CV/8Waa17LL2zYp1
RZajUCAapaJ1Fg+SfJB4pP9dDw3qhaAWgiMvYeniSNYUMStynVMf2e22WRrN
B5G/1dyUXKIVJkDguO/sKQlhzusA6RgNP2QpCZOFndd2VoMdo1rbyNGBco0N
pjsvgAWICXO3oRqaLBSmwmGga5yQJ4PDOxiWdqa3aR4mVfZ5Lqo+/WpMqULA
NpJOKrBMBXpYMiI3GM9bjJjyrfkljmxCk4xaZBzDX1OTw2L4596JwYysG/Zn
CbPEv1IbNu8txTrMrFJzRtIc3X2y1ko+BoZqcxifdeJZbkCxe9H7gT87P1Iq
mHqRSpNUKNzwYS9Dp3GoznapRVKp++jYS3HKJMny1KbI+MHwFBFfCqhW/Rih
bGcPsCKYn7hhDfGKLKgx6iHXO3fRYfPguciBCkJ2nq7/E3KSibjvzjkvEIQ6
TTlwwOFGCxAfimaP9tF5UXfw/2OqA0LHZRZLgHF6HfW8AImaaSUMs61gEK24
qZ0iw+aIzWJOa5Lni6BjldCxtwzcq17snjPzQo82pz+2HvwpRy6YQ8VR1DMz
rRLj6OhS28GyXUk46DRb8d+Scl3mFiA6GDmO2ADSfnlmbu3JiTo3C/Wzrdau
OrY/MFFdoGEXC5XJWTfArIosKXHhbZGnqsMrUyUO+DucHqMMIFCTCO11KCqf
UACYOxFX13/W1009fuLBI7ERv5TFQLVONf+E0Q3h0XAZnhajAFjjBZDOcgrl
rNsq5PhcKrLSLJ+AfWAU9AyKkxcYa0rO7Su6om3qWVg8zSTVae+Av7VLeGmL
U+EDfoYC+Gdquze8Ddw1bkvpY8mi7i4bqmkECf3eC3YBsLkC8nfzLrYjRj0o
Zy2E11/AI19DS53NBbUB60tApUHjksEun8Y6PqVgl16Qp+DEG26Z87LAaFRe
P54z8Ws2/FmxBm4xyM9G0xUL6tlqZUIcqN7t2wrMySnxmUNmi25xQkdjfZLn
j1gnqmlDN1QA5XXHx3MhEZLQ8IMSNfRLv/knE41riWUdGbWBxuciZ3d6PFs2
K+ACCzWtks2q8A2d7/LB2D5+8zpmynh9bAP6fblORfVk7TQUwfGMtYzSzWZd
09x9jQghgv2RoqoI25CZqH9uI/DRlsEdv1EZezgmsWRf+BUm+gYo1NXUfNUa
BSKOMlvthQrk2jIPJ7rHpbMdf02dwYPAaBRkoYM1g+hNMKfpnNYnpRWEzs3K
CeGu7fDrm+pYzgUsmknUgpHiT6ZdPDkWM1JUWPPhTkou8A1cHv0Ik8fIF0Go
iJBGchAJ0F56UTTvlpypC5TxdWs07SlRyfNzSwbrYXGBtm0Of1bfIsKk6wNk
yuWy+jwDgN0mm1oq86WrysvHsxI6Z+3ScbEDGa1oWZeVfDF0F1BLjMwZ9FeK
FFQaX3MW/2quXcrcFgTHWN4VSe6KEV+w9ljGNJPx/yB8dq9ybx6Pao5dPvI9
bsJo4WkxYqRTnZLQXHG8hIHPMKrQICYSx/2jSbsGZPpuruX4I1bUlZmpvoaT
jS6gvj3wWKeYr65T2mMaP5i+kjK6VVO3nRp2XRtmTHqZagWlI+ZkWhYlIErP
wp4gKCMJO8U6f8RWEppn2NOqyC3KONkq+DgGLBxqITVS6izbrl2wTrm1QqpL
jU8kuJd3A+PTwvUQPprAnoOajieGwnZy+jtA5F8xoaUKWceOix1PAz2uRoHA
R+ivmIK/GK4x3/XZDpCKBLzcs4FRtoK40ttTPJTowzCVsVtFlzfo2XLOQI7G
ZSLUkCRfEJ3URNPL+Qbt5zo2ul1SYtVWwlB+JiUEJNKr6Eii4Ac76e6AlUgR
7HFTYEymvfhxtErmR8a4ZtHIjbvAX8vaHp9VhLd68iOwN81iORzk+tXTewIy
PJfxl+1f/4JXcsKw1sMmrQV5BJtSQ6hy+2TALI09ol0lc6IGVfGwAhXX7a2V
R54UkEGRamAF+VeYRAJWT7vTvQYfyQjdTI79QZpJfMGgtlClv+MMc703LmXo
2nOPnAP/DqNxXH1uX+5z22MornFZpszXQEp3cR6hw5LECE1k3CFdlf2IVr3Z
b1kE1M0/a9+wwzihFOzp3eEUI/i8hYViqp/pgFmJTtsTsBX6JzUVKVLbLi6x
esnBy/oV9uUhYg9sgupv08nVy1Z8Dy76DDgDFGgQSRQdq/VG8SNJH5Py1G0r
Be21l2+oTVhTcRcCx37NMhytuiarGmkzgLCvN7R9M3uTiH90Owzk8nI+QxlF
F74qLG0b54XxSZLIom+Ag6ZreKGOd+773Ao0buQvpYAJaEQW1aiBGMUlzWGY
S8vk4RoGsmtFnA91UobPRru9+GEQNaP1B3avkXtGJuR3i7gagIx4Tfa0WkA2
VG/KzYFRW3TL0UCGF8ihZOi5oAmL5QS9QyvUSQEY8ZFHhjjzUC6Mao7cVwLX
owqXFTgfOW2PMAMmytfyPnA+JP4r86FYxU55XoAZ8DZHAyE0Vs+QXsE5aONI
JmBEiQqdiZkEh9phaH3QGY/UV4NdlI7kYNn4TiCm6ck0v0FJB6BMoHUVrAQQ
gpNlD8FffQZge0bZupDgjqbpXxvi3Ox2VeQt8+7QOqr9GlCTOcBhs4rsA3Jm
5aoN6lSINqERmEejxiwK7tpEK2Eg0klYQBJQX8DP9w2nlKcUJmVp05zj3pDq
nRgCh3fyVCwQRJAx2YeEWSwDonMTt59ua68mFOuzt4+3+14GAvp/ejbAk5dK
/jIfSBab/If1/mJjrTmlhCBL5iiP67rv2gxE5NwmS6+8i7+kgIqoEhXWa84P
/ztX6yF6/12iVMziS5ENyHIQWbU5y60QnXSnTk9hlI3T9IBJRu6MDu1h+/BZ
ej1InO4w+9TLaa0Uhbjp5nM9+ceCSepf2TrWKmvl00SI5/D9OjnHAxf7Qeeh
RuWr/We5L0kEdVzG2d9+zOY4Y6hb4n3WXfjNr90fcJRagMuvX1l+7AOrAAiW
hUPXbxgNDO9BpE6GM7VDXCej6cPdrm6omkFMgSbsD4sVxRfSwB0TmtxuJvZ8
6kcPCOvbeg8O0PVmnrx8FAnAHNS1D3pjDs+psTy9B2D9NwkQo27EoT2PFX6w
1SE1o7kEt0Sr5hmSFE5QORsUWG7+HpYp0sqeNwUocPLrJKvr4gFBHtIeK9Pd
VjAdVt+lVKDc0XI0xi/veCbjql1MX6iW4YzjJbZmtgOUcxzHU9zuxUiVKyZB
93bBGLXIgCMeR4LUkVJUAgN8xm2UX8OYBBgCkb7pM8dWRVfDlC00Kp3aK8Em
VW2K+GT+EbB4sXq7ywKmZy92J3t4UOVlPgAR2khfy4c9pUiTiToRafeZphzK
eeNBPvtGzpRh5plwXPjO6kliMlwwwnW68coY+V67U5uhS/4ts6Onb1Z4mwnM
yjXJBrf0koJraG1dBVUldTKltEOT900imGw/8d7aRPvJ7ZZKu18GmrXtR+K1
Bpf/SaE7uf27gDoUv9ZreP4gXNqZRmIvxy9vy6tpwbwL/BkT68BUKgxEPB+Q
HWZSXIPLS3MUYYEE4F+IQxfgKnBkDGG02N+3r4VV7pe3ym9ZFPrDiItZ9ZIK
PwGp4Aeh0hmxCLVdkogdp9kNvKHn6dcxLCCp2834D229ja5U5Un733mt5St2
OIl8umqFlW4Zock5icB046935guQsOnZPFr0cB+VThCzVkNIDY4rn1MYYqjT
/7b2ZPAcgwiKJaOAg5jnUoGDE3nzfZxprqNY2u+g6AgBUg/ERCpjdtP28HsE
DYcq3unNS8WHP70IS7MqN+O8GqxfvF5qBHz3mr827Y9S4Tva5DqHe6OFAGuY
w0rp9mCs3S1YUZghaKcil9yoBZxsrny4411yeSc3K8VZCkDWokCFhNfRuRsM
bJBCmUSXQAu2R8A04hJnBp8o7fuGxGByluDqidiRjxhobW8hly/lyQiYZ85K
BDME36GLiu3TgivfO6zjOAkPMy3aNwsKEWu2E3V/ceadeazvUhzhBKj5B/Ep
at1paekxlbzf4HGe3XkO7jr1c30Q96S4CI3ePlGufkSFdrnOWDXs9t/9T24g
iO5s6O9i+uYg7C7WhetSDyHF2cgsY79vHtIRLJVM3G+NmZOQvBkYvJXs00CL
es9L6tsjMIW7FJs712T+RrEW8fjf8l7421M2xWiLUqFHG9Pm7UD6cXBX8/XJ
9wHQgGxqDJa9ccmI7QuZsKpLGekIDEWPw7i2kd+m1dogZTdJ/z+cyOUZ9Ur7
Rdm4BAkStthlWMOvfIVsKU1bPKP7aQ3nrXTHG7LD8CLRRZJNTQOIkl67FkNZ
g2mEkfIQc7TPfYsg77RRZdbDHN9wXj1vWuQ1pfsVzy+fIPUhv07CcKLmj/J4
bnOlEOYecbslGLyp4XzraLQ+kEUowPWVXKjizt3i1wygt5418iubVlDf8aDY
NilsDA0JOngWpL5PK7egXTpR/HVDo579Y0E9nLkwvElrIFlGd2/3DJr+irNW
6lBysXJRyJxrg+T/B5tErUj1BOi3vmydS+cyzS5fPldUHPvsCYVdLrgEUBuA
TxXM4mU7r5vGJbQQBEJlo+eoX1wYc1i0pNykOMJn6QxLckRk86uqo0NW4qwd
Ca6qcMHm2xW6mKyw/DZeQdPtyVc9WcGAfwlrV9YwHCGCKztSF67yqJq2Iamk
Pk/cuFXyb90Lle2vLB5LE7WRK3nwm4LG3/flDSMir0DeEsjDk/zkF02vqpDg
ahiiLxFOKmDIGBXnEAJqEjMcx3Tq3/f/riHuuyLLbyLm1X+hBpKxW978zJA2
Jzcl76l57OCt1q52WJyYIcJECNJ9cqofTn+oujcamJYDDRYgVTBs3rsYRZZ9
lG1yLN3dirWe/48EtXpkyO9BlUXEvnEZ9LrK1Av17rZYHxFATfEUFLOIy7Uw
DD08RN/3OhoCT5fEUGlTOxeuxR56Vk7oC7Aveq5FVCfSWG5fDzRmOZsJ3f91
EKdWrSiaC0d/qZgyrAw7b4ovQ9wGFTfhmjjyaceP+hqh5e0L8EgZVi236B0X
neo483xlyJQEfGY3htI50YDq/eSn95x/hq3fX+GTBIq0EQqPREPCXwTERntH
u3lRhdrzWtJAKxCkeLBJLzua+0PkOGQTi7G1F5KHGyfTvbqF6E6tBSkdu22t
ZddVOMnY0GhD8ExEUfus4IjroiN5tTQcJFPd0oCpHZpRcjy/pUKGKlI09+hS
UnN8rXbErNC0aYDuFx2trCJJA9UfiW3FXdZ4JFfxgqh9A0Onw7/NEtAMciMQ
zxv5olTP9YkuiI13G77FKOBVe6hv80C4ZgYnMftykqZEWDkn8K6qAucgt6Kn
l2d9q4cddT1mBPHRUE3rDYegGLvqZTv/Dd4DAEQQhPREwLO0rZMwsvRYNKSX
9xNK4kzt9UucjG++E5AA+BEN78sP6I4s3Rtl4Uaqc17XSBq8rS4EdD2PJg4p
5GMcNX9ZN3lwM18s5NakkRvaxxrXxTxUZL0WvrFTfoC4fqT0oCM5siFmhHdQ
L92OxRWF4tq8xs0PsbBuk7d3wDsi7WD078EzZ6Mo64NtQJV1b4k6H9JEru3d
5EX3UfwqiGE6qSxLbmFi9Ds1jQwdXxFCqaN1dd88x2NZq54ehrxCOqZvpHvH
6BOQheOvwdWV/RhJIUoB4sDO8usN+9i0mc8ZN6h+pyUtaiR3JFFmgC301UpE
FEPA/3xbh5YarrsQpLtL5F+Hd6kQY1CvjRjkJcpEER/fRZUgSCs4RJbJinW3
vgsQnJz79pFiJgra/dkjsGBgW9w2/ZYcSRQ+bLXyOBvslho4z0Y+5RFKDGWG
tRPXcU8z3Fgf7ES6iU4j2QfCZE1RKfjW4S6ipPQsNYh7leOmbUS493WNuqiz
zn3+FFJE4yCM2c8v2vH4cyZl7/KTRDPQ1MBsf2aSvYKWcQ8bV2ucqWGd2Y7y
6eqDSeGz9BcgVbYW0FlSekG1vBVtfWhdX2hhWIk8NbyMZ8wIe5PPBXWRS/8G
CeZvZ7rns3r1ohDH+nUYpFPT2dbNO4zTXyOJAuRtmtuYjFsrukmgeoG99S42
hBbw8XznRSyQjuzO982PbxvgWLuOYPF35Wh3Tx5fHY09TfR0rED6FCqPEQvX
Drz/Hr3JtQ0cOZQvsFC5RZdSNkf/WmvJ+n+tWKSYWA6Ltgj4W2Uiq2D7rfPa
4m2yOsr/nZ1GbOVPHkrqjo25leuSUKz47S07mFVH7w4iYv0CDQs2YwSurZWY
sQfzlh6IEufX1DbErtHEdZDmmqO4fEEX0GK+XOm6mFkXIDusZTKUO9AtneBY
72vC8REyBPo+LTe1AJc7lCEOdgnT9NtSS0YSIjx1K2t8jQ+dWe9lSrmtNL5e
WdHbnueKntj9tFoSHX9JnUUluHB/oXRcoVdXP5QVWn1iqrD8IP24hMPwidGn
VdIql6LqLagxhS9os53mSqsND06Hgy6cnE2IkwA6gYS5cUTnJgpWVWVR1+g3
VMyOfxPnJqU9MVmhvI3ZPyB9VFgrlJY/ch49dlv3J6IEfYWj0pCnIudlM+CE
X6/d4BD016sbFcxf1yXlaEDT5WZ2FlZW9qEZcKFIGdhYr5Z3FfG1iaA52o/c
eSqts5R8JojNgk+kUzeiHmKQC9Dywz2MjDNA/eOXDssfCKZECSxwQVQpaJMP
vzupPziCMVvQwOO+ygteLsXuZ6uzsfEF8dVJzFWTj9KBZx0NK4YtqIDktHkU
m7MKVXwosEuUQB0pt/antDfLTgd3/9ZFlG/coZ0+VFonzcB+Xb5aB6TDxJRl
lPJRuRNlYXvETruMOEBcALPrwE3eHbi4it/8m/Z56TheMmM08/KW6dJMV/zM
tokIaA8YZhVgpnLTGFq/vF2kItpecV1m8+YOXzsU4zYuiOfjZXD6ISKMgSWi
5toTNmOUORx0Bnr+p7fvj18W1W1ms+Y5vPv1giA9zClsnJssFdfs828YrzWI
qqgFOKhh8lnOdyUVzHJZzPt047vrHN/bmsFFdj/oZRXRs9wg/Ebx9A9vkHY6
fCezBs8TLCCNAbliJAtDEEX37O7rSoEJt0uZy0OWAY93NW8MbugUFa228WkL
roeh0CVhtcwusm+xCohRqKEmNZhV2qsvoOLouwHyXbaC+40pzjq5M2+35v4N
WYWiLGmuURIDQEqwYbQsmLeXLsXT/EPKQ4mPJFUyYXxX73F5sS05dQBlDxcd
nNx/QoOuNQnkTFLXt1jBIrDpxSRWY9WZgPGvaHKvg2kKmKd316PcFCqLQALP
i4Ln0wwEfAcVXdxkTw73xes31tZc6aF9233mb3E8rsdDMwJkqlHAli+mMmQd
QNiJQ+BgNEFILmFJnSs+HrJxTuwlDUZMNtpNRmrRA4St6rLty1jHh3vfUmFt
u1KAOo2lxOWszQjswpkF0BU8ibo4PBWga2wFccVeMR2OfH71Y3XJ/7r6IZQ8
TqSMcU4uzdfoX3esOE0wj/QaSq3upggcopM5VuqvxKHmbwB+/zji2cbI2qDZ
hTCmntVNtNAFvn6AoJpq4qqQ48f6cebvdV+vA0J6AkSCzk3Do2z/vxrJBwQC
8IrWkvPUHpAVMSaeuXHbUqggrQ7cDDdTsYFNxq5KT+Z24bX4tQpoDeONiTfW
3daV+lhweMGhRaOngecedLs+hGutP4zoqyPyrcCKC485CmuVqKcQqRWktJn8
vvy0vT6h3Hc5nHPGrPMn+gLAvy1WWBJi7eVwzdPOhGmZW+Cm2vo5ujbx6HYQ
wHXtEp9a8CsNhN+6Fs0quVOeY3A34Xo/E39AW8HLcZ67F+XYCpo73j0geC+D
Z+O2ewanfv8Ihzk9jvkxMEtpcPBkOLPC9vY4J7mmwYgiqLz5izTJ84Prr9GQ
jiQBsUpEs+hSbrrNlP5JzFlbUEQyFyfo/NSUdMwKVDyznhE7qfM/iKb9n1GZ
EweK+FP/Kz/vxXUliO3A/HQ2FL0AAJe9X1pavkSfj+X8Yrw5J5RH5RSAZRTG
M80lm0sb2AmuRtssdHb4CIH55pPg6bCINDG7OkJIQkYcjgsCNYMhZCiZmDjX
HHhJJrFURfNZL6ImkDFK3Jfa9OffRheq8nOzwWv0W2iOJHw0ZrBSLga2G7t9
8duXI7/xkk0Nj/btqV4ydAFEucnKSgzcCuMRM+eF1wb9wyJ8i32EsydGHofe
HCoMHaYpi/E2XLiRNSeLNxxKcXzCBRo/Xz6sAup5jobA7c1e9fedesgxxJR2
mEGUjkbakSIa8+OLEE5VEt/mvW/UWPXASReZFkw7xTJsWOFdfzOhihV3MRIa
IcHvzVXnx8ipAXOp9O5wKcYq+pr1O3KIvcefa0DOcjbPtedEf5gjXC0IGfpD
WNmkDT1qAU0t3vGRWycMapRa+0XVQX267CeFBkHywzM7mdqAsQbbv87CBzlZ
BnsCSuDg7P+FLCIzIfzfUjH/9pac9IjKcl/yCzM8cb6LZckgcgskl7cd4+7j
gBg4K52CrESv2m3X6udwRh1HmlxKZW10MD8oUL7744K00Vcubkovz40+yK4b
irUQ3XNSkxPodQuM48dxM+LXIionqeWoSx3GKvHZ/K+lzu6e1b+fXS0zxeEf
yBIXHRBbO298TJCpshcoXdLJjqgi6LxaLsN1bTjLihgItwe2/F+ZquW4kY6B
zOJ5gEz+Y6jZK0kGIoC8dWC44SqlJYXJ7K+Wz5z8YzQAgjhDUWvT8eBgpHaO
d82L0FgkKzaaPgqEShkSR9hhv3MXOnJC54+iplWnOPKEgOv06nUD57wL2nxS
WS+WJCehy9EuPQZPdFLJ99DrEZyEvxvP3/nHaUm7cTo9j6JxI3k+f3ci95iK
3nVqYL3WEo4RrPa/RuRTHQVGiRfobEnqL4Vrk8UjBTUfdvdTX5cZKxglWGdK
xCfv8aBsRleHrX6yzdtoVcc/xaHROM0/T8McG3vo6u3HxtvhAeuXV0rUQdQU
ae3oUHzIUUVLuriaji5vI1Y5+PaJDE7/z9vabOQbqgVc8XiqRx6J4Lo5jiBj
1H5q8Z0r/sRw55s0oXyc9BVwgAFLCte2EAs/gdZn1WrQfcb3pBZFFqgncogY
Jo6FAdp3HesIMUIrjVuCYKKo1x9eZdmKJDNdLOjxR94wL7SzLIdmRWFubDc7
ap5jV0h+/MRqsFfp3OgCIbufVyuTUku6MOQw6uX7h3wa8Od7JKgWzijwCojy
K4BoSGEzAKEQavGS6zBDvKt6TOnNe8u4u24/K+0obkStMv2wDFnOo5co8wYL
j6u317XAPaKcrBUcgRRg0AGPEvKpuogz8FtiEL0rd3M1Yfc0fhuzBvTK1Xcr
5X0KVuh3uPTkG/UsR3+urK659hdlLRPRB0gF+O1S6zu40m2F0LBuJrRKEG4u
iYWBpAC6LPvV3K/TNBYqCxW5kkV++yzAlpCIqNcirkRUZwlpwas+KcDHahPf
5kUU4+f/d20lD2IPw+xdDbwzJEQdfTKdm6jAMwSqshTUT7zuijfrj0eG/54c
rw/5yPS73d+zaGWxoyORmV3IsqW+RuMkQmP5LnQ6meaPBzlQ9xuSnmTWIFKz
CDJSGvOup6nQq35wphSDcjU8IvFzNgcVgqxOqcKbuYpbJqJS2FrXQygsG4Mr
U1SKmRonlit+OWYkZQ5ZR7kf1D4hHfcpC/TO0gwHxYfNdPkeyDRYTIYXZfER
DbjKvI55KcffbpjqcO/9qqI+Fb8CvshwlwH6X1CwNCZexaPJQazCCF8j0kHK
82jVTVbE4KlKTtyQ9Jk2CBZ09KmINXOUEYHvFerp9IN+/JtjFETTLbAFXaOk
t0J+8TniJamrBtM8I8ooQ0lRTiqVROHlJMfZ4+rUghmze5/dpaPznZNrRv38
48ZRtisJOogu+hAhbeBMFQFu8H36EiMhRaS+LtwkECvLIkkrMEWGssBQPxVp
G+HANzYXpQuMuQZFvfh60/JPJiHzZWqBocvtVVvrN6rRQyv44grmCpd6Hd4E
ZJSeAEFd7c3Dk03KtjRfAcNOqnUqW2HXuP2w+bgkwTMCH9KO3kZyA8ZSxNNY
Vb/5d15oIDrEQgdPYztveTM1QpZfipelmznFrZlq8P46OkQhAo2FitxmfTuF
EQ6KRUUKn5MbOqqhZCqcxLMo96+UFzBWMgbfXlBlA/So0XcVS33zrbNDS1Ow
9M6hHUEXVu/zthw7vwdEoVBP8bZzZTfA8oVDANKqDXjxKJQoMoGWjY0ra+uz
PeSP4lBbdyBn0pbvXmduYmu7UAocp1S2Ai/p2YQTj5lZ2MxEcfOaK81FrF5/
+XCO6Ta46GsvjldV2sD/S7NWuh+IXjp2SN2452v7uBqW7O7f6oSp7BPT8ctb
Vn+LkjD3aHZ3qjwMA/ZQPol60UqTzSwh3Sqv7sk219NNB9dNxgQlZpMeEiRx
vR6IQD/7yGFE42E7nV1VKeZ8zuei/DU53b4eSSqPvikFwUUSRNNngruyebqL
2wtGzLbRVmh61yIXWZhsLPMo3AFnPrSFfqcIePQ9lwnr88S6RGe8D+hef1aJ
qXzA9uNy1cpNzLONb8XQ6daS0WRKFE92YE3DxkUnUch4idTN3eqIr5KcmRVU
P2QTZzovsAj8KiBpb8VjHUxb/VPWrzXjvUCE1yMoeAy1BoopK09VLCdsJaGe
Le/8eoYDkmUToUrf+vMTMDDw6UexmfqOuxFbj2Tvc+RGV60gK/+hxJr2N4+k
XQKl2u5TkgP8/moPEDRAbBDRN6T3SRTsmPVLF90M22x9s2uedgehUNxOBFE4
7uaMP2JVjkIMaUr8FagJaluO7/c13dDs6a1F1C6gthpvFPAhQctix/znGn4w
tWxm3AeQEXFJK7RzElLJNww17q5sZMsnJRgmHfy7D+yuH8OCaI3Sl/jGAzQi
zkF3BmWfEaOHlY+yFoVtAAwUyNmdyMZqJNO69faYN0PI8xLnRIhw4Uc9ezsC
LfyfHOeMmj56RoXgSTer71Vx5p/+t+httx9EExYqPxvsb2DUCdLcfL9xpXsK
ydn9e5OfyFC0N9Az2/kWsdn4VtUrT68QcK62d2vRfwiKucoZO5DRAV5qyNEa
Kvk81/tmuMuzJZUkug2uLn5SNosfJFTubNne1x9NxSlHdthYaGq7NSbMnzbB
cXYLKJVdp+2guWEu3oTcbcpS9/04P5iO5P7Y0Fv0onzDiXv18JTYqr6JR7xE
8wH67fSdKixbWiqMvdrbifQmXajhTAq4yYboBOtQJVs3BEU3Mi9wiJEg3IcF
YDgXG7m5YWm9mBpZhejwkNIQfBlUXGYaIg31Z1vuUGWvvXs3MMlQ0Mosk0KV
1iTaySuSodVtr5DBMQMbGpqyoNwx8y4KVhne2/Aag5111TQds623BYEdSY+J
BQqEcDt1st68AMdSwWZnqwi+AalI65VxknJoVOQrvy14VgF5mEiJX0ptXI3v
iqrX2r6qhKzNMU/DPgsL0zIw/av3kHCV2QllE9pphzvvsaOT6kTNySE0Kx62
CT/1MwGz0wN/GWI4COVrZiIqgunKKxyUNtfwxWNWjEWWHmzfeF6eTI6UvqWw
3BVK/jS7wp1FUy2vIw4jsRiWzSLk1i4hdOEIpTM2jDngf6dI4tjqxbkViYkp
xCLnIqOTUNl/4oXjyhT48qKFVjYL/BDGr7SKS0Ta37dpVMO54pYcOMpqb5YE
Y+6AYiJgEU7glhWi8HR2+AQk3vQrQRkq1ai3CioK0/7512KSlKTQSiSmUDnz
7UAH1ik9hBmEoUPIRdAXi/Qqh4Y93sPrpmOMuAI2SbQO48/kGacd6yvmXqDD
RMbvEz1JMSsIebS5fWYzQDwCgqcmMgqD/o/SL5HRs1gWURk38cmV4QlLwkIN
sf6bU/OXGokIPcebd4GIpDOeu7Nkyr6aRlAAMbPpm63vWaySM/8CtNFJ+OjJ
79DBdGdwqgOBdA+ppm6fi5tHMwbSP1iQyfsLOc3ENwb0QRzGaGDiwJoK/dr+
XHnILoL5UMdCdLr6wWgcveZz6b4IOGqsYgIvl+JMqrwF6aDWv+RlJ6gc+oXy
R+bFhuI/ZyKoFdiFUzGWDdzDd3QSMHZpZyNKgAfhHutKGIbwOxgcr0kNUe+Z
2sz0Rg3h1XX/yKnarc91lOsMpiq9OrxTuqgEQzt3Yg/IzPARG2Q3HbhsHush
IenDrAw7uGrFJh2Kj0L1sMkg/gcOccfwAuLsWK1GcdNujWPdaxGcEaBvssZ/
adZmzoWj0H/hkbzjfKin6xDggMHRkWw+z6Cx/ySwWdqXVWS+GyomxYleJq8O
y/3kRCRenfzUAO15hi3Hi+vnuuUJrK9fJ3MytwVgp68smlm1QyFEqw7gddSk
wKc9wXFeMdAffNyasBa/C7IHy7014i2jbzGluU7A0h9mFQsdMGDPRJzuVB7G
tYiADbR37rRb6CvtF6/WqQjgr3KdEHS+drc2T4k2VKhT1Yot1UBpz8cud8sy
5hirO/GAsJm/HcA0UdRCHegi8srMl6tBILGEbqMgEAAWMeJe6+oZyNcrljVW
8WTZmyyWMaC0zS2navdt7JjMnH/mkiQWg0a3zCgZWFPD2vj/GHCchaGDqGxW
PN7z5l1A8QtiFrKLcQ3RO3oYRoXEJQb2arh6fg8pQu0EiqqY4Qxcku+vO1Su
ZILcRwp1XPN89Q+4kailqpRikPsF8YtQTKCOqNRZwPbsPvhpKMeskQKS+lGu
arnlfpPXHUdltcD40NwUaEI67UQk3O0L+jchLiX3Nf2ygzgv12rYXAHgNypf
E+be+zZlPwq/ryGgiQ8wDoLJjo+iyPOCN+EL/bem7MsLJwrrJEZRd11rnaYv
9EVfE5jwNw3umxM9tS9R4XTJ+w62q64ms90lwnox4eruKMgWaSSInvmYjtWp
NDnlmmTmD8WSmqDT8h9+twQZ/VnK1w1X9jUCegnLl8TLUn07kO6/WkbnIdQ5
gNINVceY8SQTFqkhmXPN2rPKhFVOntDVBw5mH2x78tObBWBtVTOzeIOxEaoJ
I1/U+JTqzUTFVP25nyoRfERzSJGbxCTRxuEWIDJygIEI8aO3+DQpld0+et23
E5xvCj0QgtPbs4YQSSBcBWml+IncswBdFx/AQcPufdIdcVcY9rlET9yYRuj4
i3llrjVhBIWA6jRaCjSC25xGwmhjF0V0VLKRO7fy11IHpD6tr2dj7So/vRc/
bedL1xLpx08Am1Op1ORd/T6Tc9/qTGO4sFX49QHPWyFfNRFpWraRw7EeEQ8p
2EwhsQ0zh//cVqijz5esfyWtw1ofSny40h66nHpTxTJ3kGDa/t6pBd6ci5vT
CaP+4mdD29K8fYfD/jRjOzDixRWKZ6FC2dqMIkGoQ8dridIjSujKF/aT4oTK
uoBXHJhCOIku9SevuCdRXyPRWrJeVRvS3Y9Bxh0UbuMY2Ch2FIkg07VyxAz6
OoyD/JGkPYn3AJ/+y/VNGiSvLol8E8VUicLcEtQV6S/9NJTjViJ14omuCgVJ
mLtVaWN1vSFgSEWezPLDiAAZpwq7ZArLlmD+4LjEg1QSrZtf4ZPWCVQU13I8
5fQr27yZj6Ru4P3Wv7koO3f1DLM6yUrBRZcGRSlsh8VLqDyjfHS3Nq5HvjLE
kyFYrlXqJ7DbIB/RWY5ATfN+npTGAE9HtA4pls3yUU1rvrePoKNXqg1irL8P
3u4CRyDYERtbTUKdMi+jG2JoLSdQmSc5Fnk3f1bx1z5Nv7oiem1zjhkmxlbp
oDNKVKYTMCBNu38uO9ckPMjucuCIEX0D7BL8H3XmFbHbrQPc7ymRnY0vx5eA
NkbBIjVP0qOVNEoy+EScDVjf7xrNiX3MQBE9bpHd0HFHrhZLa/O3nFbLOQ7H
3ZzMf+wQkEoBWPnQeHdqDnN3CHnGcri+43+s2qyB6UZPfljN+Z7ksGk7Xvz5
BbtjDvSKxThv/Iq8ztstnajkIDEHagbppZTshnN+bLhoCQwOejbc2Eh/IgLb
Kaa84psrEo0SfBQ4cTXtYKKWWKFU5Snp8cBQWkhImzbF2GZIzGmzJHWPFBKS
UJ7U0fBOA1rwJsNBePJiJ7nfc3MRdzQXPg57AJZ2Cu5q6K+qba18gqAVcNj0
E3A0hxBUa9AhXVKsVaSQHAm39v4VqKfK5X8qkd3cCGOJQn6knzXKtoXvAVDn
P3dDM/xx1JRcMkEeudjGes4KV7HBYjHbghZ03wFgQTBf8HD3Zwy9ChsrJ2jr
cya6RCE79GvRAGAGD5H1HDF1c+q9M+gFUYqIPvbMiH53XcWUBYNnolHaMgAj
abT7gZsaQSqfHAdLugdx8wqea1ZxrVah1C6ydPNAcBeAeYH9PjY2KEPIdH/6
zSg7xlCx4j8c5siPxDA02tBhzQ4XJ6WAQ9icklvJjySVxhXVMlEtVMrwst0Y
JlMm/T+YWtBkB8U8Z28ViMLJkOY37mQtb7PjnzfznQMYklafXdiL5fdAHvXr
wcAVgnK10z1gnOxumQt+MZse4yywwAIDBmVW5x5qiGt9aOl5gxFdSJjiw9Ks
UiFrUEeR0p42dVIU6yFIjrYhaZBQKjl9Trn64hctBalRLmf2PPw0S7/ADyEe
tk8m14KgWoF/lvWk7dyOovtFbR+0W44cxtM8SBxSnJmsFWe0dXQV8ipwhHjS
7ciOYWUpZ7/yW7zc2sUEBGdPxi1g6rA1S02W/wocEDuJirDsqO6/Y9PV4Fi9
UPjqRK7Y/IwXoERD1IRM8IqhjEiPW109TAXc8qX5arw/Xw/LS+xbCbdgx+LP
dhVJjYL9VAVAV8GtDcpLFG3Py/hqa23Yx5eAK6XPO254508J9jBe1TuhHxSM
kITdwYpOwxooIgOxx2pY8XV9cDFqblAj9/7l44cjlHbQcQbEAfoB/iz2lslU
AAyqyt7iDu+73kFdFqJMwPRgPLXxfVnDzoxR1DUCKotoKigyUWIvYfMPFgiJ
MBRsLtJTNO8oSelJIAWCpQsGsQC33uXifgrAAZTd7jsCkCAESvtXm4rKiAFE
KoRfxjRDFW0KTwBXYnQoCujCJcFTie6/yMIAaPILhSSEuo4Byf5xxanVzqlR
imuwF6dofwUNnwPzrUBvN8vVI91ZaxsqDbsCqYhY+mSilcmfjX95DfqUNYVa
vBRkWSaD36XYy9qdqCzF4mR2tDjd2tTLQpb7XtGYMs7tHe8Mn6k9l5Rzo3p0
KjfeOHo+WsqtGdPP3omd0dWO6Gfsludl45/No9sDOBcZO9G8dO256NX2ydP0
zgjm11vEjRabKCu+UX+KdeXyLz4Ka+GsWUU+LowraRuFfkqoQt0NpExC3zyg
1cpFLZMLbpw1R8DuxYai+aGhCV62TbRksNR+yOFufBasldSENgI6a8vcxM/C
fLcCXry76s+5s5RcV49ZxotHazjSnk68C8aCjWe4WZvihPYLm3mKpxqExX2/
prAH5BOeyyKht41YYM2Wj3uWB6yiVfZpFeZPPaeKI9m1KmczZLeTaH9Pwcdj
HAluwy9BBpQFGi11Q7J+jW4C87cAAWN/55ikLgu4tIF3AqhCEi41bOGkl1XW
5GcRwzRijzo3dopM/aQUGsE7DvKZcwPCujWUd2dslW3E4u9S7f8yiPSLCSNX
kZ0oil/fdoxCjsB8F5C9fkOyfOFr7JiWys+Prx1gy/lsRtrHtK4DF5pdMWiW
LkJOVimKc59Khw4EkanSOBXTrB8Q78o5ieazwZJz268qHiEP38LR1fkpcjpy
RV5bubh+1+iCR0jsf1e+XmK0EtkV3vTebZrNbZf/Gik8lqPqBtr0sPlQ/NBc
ZmKloLuJ0JFFqep6+77CsMadiiEJ1vuY4sNufPcgHLI/mepUvFDOBvcSPYvf
6J0YEUjxw8w9M0Gk875A9YdhckekXytoJrmfifYvuOsXJmgnvYSwekxzqmj0
LxTLT9hJhKFPxOKxdco+R/qWovv5b/lKb08trG+wO7kDHKHRYGztcCWZBmXe
7Ah8tZPm//rQr1LZAVk6KWoRmI2Ku/2WcMBOH1sqkpqYD3dhcV84xsNSOQqO
LhZ5BEl6nSjQRdNIhM8FpWJZIdQ5CavUQ7OtGvg4m3DgiuK3NwJwAwAY5Xu+
6o16dg6J/u4cUJj7JuqQnT4QXYskLXGuN31XZfQhn4UlMAht30zHGwZfiM3z
BrfAxlWYSrvHCR8e4q/8lIyWOUP61bqI7hqnxBLdbQjJhC4V4JEC0b8/A1HS
T5XxUSS4ZsrsIkMcP5u91QRYE/JoArNjvDnZGYxYI4xoFkMejDJ+1mKCf85m
twL0y3qUq0GbX47kYxCNnrA5Kv0KJjz1HUiSHeFnQTQrfwfdYiDAvgt0TeeD
J8je0Gr3wagLvUYwBVY6cYdy36rxooE8yoRv0cZUfZhwwBmaIcx7jUzXDRYq
FCrLYZa+6C/PXpYNcYtqOhiVfngzCa/ImOB7QylF9PTHLUQNa6Sycp45uxgB
QT9D12J5oPW7oVSyq7xmppXVoxU5H4JV4VbW2jDyAc7RaElq/g65edTn4ccS
xN7KS8jWYuItAAbv6h3guy13plDQ7XRxWMfkdR/Qs+Xrq246zvAE8gCz473v
w8HGpymsuRYk9V7sc3FeqyNvKQyzYU2XYMmvuvbAU15YFDu7+opGZHbM6zUs
0unjwM9OJnU3QPSoE7E2GfOASuE0Prw6uireQ0aVnldZWiyQZRW3PhHQFCeD
iIjnx7oEHgdKGCim6k0agFt4PBoWGIFjd799HFhk3sikXMS+OCovWkkRXsiF
cHt79lVAjL8wzB2WuPdysXp1GdHXJZbHAnfQ2qOlYHbIPvXgcE5PSxxR7ytc
Z7gzEEgVivzHJmvjgDarJRZH7KJF68wM87ko1nlewY18zT3E2Keb2czfcWfy
KBDvfWirsCsBDL7ZtUpZ4BcJOP59yjVECOyU+dxCuX9ihJ5Gx+JVWAg3+Lrn
zbkCoKtMJ6n3EQYqn93A1EqLJ0wSmafEdKVQ3+5Wbph3bXAk6Hni95/EZz7G
ZKbELh4pycKGWHqyPVNzc/lc5YLWXuIn9afgpedNpXvcg/Z0kkESWnL/9gZ7
/mEg4ngwTe0sBWDWnBHwuZF5maEMaXbrQCOk72JSJogdDJssMwVrAaemDRuD
T1HExaz+gYRviqILY2lY4wAJ3Cm9sLk16RupnjPVlCkWkWsWUQmaO3bOjrBH
ql7R2yqs9oYs4XtF70MclYX2q5UKF5uCj3AgoeFTZ0NjVo8UbtQTl0ediD1r
V/w2663THt0cy2uFkG/+Og2wIK5RzmOMSzGrfYPy1K7CZCXHiV+l2u68gMWg
GQwUzBfRrgAl7UGCUsVrGLOsUOjcvOD19f4Lo7LLEILBepxo/2IujHmLZuTE
d0PaRyPHpMcxGETnIYmKeYbK3s81pG8A60Fwh9CrNua7eqCrTVx1517dRiqs
v76F1ivBxEA9vzZIj1j/gdAdMrn+U7T9eE/sTjNXO+CH91ChaAUEZMc1ZnNz
9gSyalPbai36BRiG3T0DOHiht4oO9pijUKvvTBPjL5HX4t2q5NIGPLczvPxP
FWra08yCmxHi11+PMYwGgynEQNZT1nkmvF9j8JDlrJosfS7R4p4VtS/ZLBXI
Oaz2zPAedHItanNoAXVaKDQWJogJayLzG4GEy9FiS/j1qUz8Ud2iZn4qe0yP
YwLez549L0uX60VeeLGQMz5cN2b3rpv/7rFJ6Rb8Cmb6fwAIV6RiM0S9/SRR
4RW/5DW1tq6mWmF+jOSkEj8WUumqWu9tO3bTM/nhEcgjc3P3a7Lv8btykgkH
hyznLhuxcEyIr6wk5LU+or70j0BcCY9z9ZSQbmF74iU2qwqFBKS6OLArV8ZT
O90asmzVmmo90fe6dBK323PsVVrS7rF4djNiVS64eVdGowRYadz73sd9A2md
WRyxLuvA0omVNx0pjbIU76cThrs=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "B40jvh7ud/ahkCWXo8CJP0S9JYnc5+J2pwOdONjrEnmjRzb1YpxBEP/gM90XdEQFf8e+9j+GJABVN1VA/EUgHmy986oXHU6n9uJJjaeBsR8h22iSaiy//95eH4kKFakRZgkZDqWp0dX7AUTwRg4vZKk0rom9cx0xsiuc1Ki6fTzxDmmuuNW+yyxk/luKJogixDl7f05H1PhFx3JTfD9y6cRFGovJ+RtyYHOBbLpk0win8Jdf15cfT53/KNc7G8tl/vuqfhCAr+Og9JHrGcNQDS5hGydIlgv11+LTbikzf3KQesgEjssSWZW/bj6GnasSK2J763MAxSbBdjX+u2/4sAja4nOLkHhVsaMjwk4h6HSN0FHhZNwr/i+219cMy+D6jCGEN03Tf84UD2ZxdLPIDWKwxlDny0vK12Dpinrp0uvqd+hO15oJ/ndeUx43AAunNgZb+tT4YqURJxEpfAFD5N8MWbcLpuDZzZQ1Khd64rpyTYJHPloa4r0MVDxAp4QTUj0gA+10HbaJaWt9vPBQGILiCwLjYeYNCCUbyDchRu74Jg3hpXyiJEwYQfpyrJN8mUkXRaLWemXBJU43otHyRj6NVU85sH3QXPMJR8MVszUo/16ZrxWoJCreWQnD1BuYusR1lVLaryhELRREGWmu1HYdAH5ArPoR3TmQo6tI94Ljbccm/00/2ILbPijrHyQuXcs68sI1QrFQDiUwW174AlNPmss6zMCTI/Jlj+dAazaN1jQJ60GiFBTcIQ0hT/jzAsyTkkCfINmgXHxhKwOYIJayFEVAVOoWJNWGQREUV2Zd4JaNf1qPj1Gsej0dndh+LXCl6WXkf5bA9jRIOz7JizqyPVaS6L+VlvQgXamdlVYux8JqhCqJ5hxqTzUVi3apeXmn2g/Pw7QCD5OecX0g3hzygY9Df2axyMQFniT+h0d0PifB7Z91ck5Paztj1BeMaIddpacfcYT7jD9XtIM/MRmde5J1kZJq7azC8dQrCO7jXMKLANOKsK/Osb3LEMX4"
`endif