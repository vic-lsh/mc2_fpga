// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Gyf/7HthLm5RdPuZcvZ2QJLD5jtvriDgMCTXllgcr+AlthnSh5PZlHGps07g
Ga44EThpTKQZVSY1n7EDWCJODV/CsGv0MId4BNXZbroxcZWlIitu6acSI1LF
Ae9Q6NvP+tKSzrxxax8hAneehLrn5DCn+iRyHioOJfb4vI+NPrvva7QOgNyE
QaY+OdbtkTTjTH2HNQawhUxdmQMQfJWnj9E17erGcOR1/UBySZxqS7mZqQ1P
WOM4jkVu0xILd9rurz1gGWCkOp99+sq+y8YnnmXZCaJAPIP57tVIFzGeiBoq
P2MrtGCEg3XqQ5OBjF1f7GwSNMzkxQtULyLaj+CDgA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bQbEL4P3ilRm3AlnhWgr2BC5S/dTGVBPE+JaSD1/pIuz3VRk45YrzTebSv7u
KiPU8HbGux5n3Ec8EQ0c92+0gIt4ef+RE5htElmobED1HT6ll2zAn1SCwfRQ
8WF69J+zdaXGPoVh4afChfxyDVF0N5tL3o1REx/4Zihiki7/Z5CVtXcwz/9R
RizRRTYMIQsipB4GTSEhTyWbTQCQ85oSvI9WVdr0f/lbhqIylRdeUZY7besa
KgwjN/srDoDm9+6Y1CJP9ctNEDLYpb48I6z2pEuzwe6M+yZTsP3ZMkGN0fl3
i5tljLGMRlyd8VFwBDBvCCAUC9tK3aXZwDH223xEEw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Usz8buarieX89Zxipx381YaesJk5ljgwaIWZKPeKPiv+VibLyha4FPQeyjJp
IKXzYOWg6W2tA822MbkzgbFJmbwdPKJsay9WN+UYCUOGvS5pIjUZe8tsD3ic
owiZIwdJ+d7mKU7dGPajIrbGVaEmB7wNZ1yyeOsB3YY8u3kpnkQ+ecAwvBmg
GwX/dFm/083GUNa+py2+mmLJ3RHlk2LDWL8JmLx47/vz0MRh02RMCrRrUVKx
Ll7S7hlR9Rxr+ueiFZLpjVBBUbRrfMf+FTJqW4KBTvVh+5M6w6e14K/W22/4
G/xoopvPgOtqhvA51it344Rt9eg4rVplNwI7aC+gYA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ejlZQ0x8BD/9B1LfGjtGtbuZFo43i0s0FCU04KC21A39xhH0gnFGH8m7EJgA
hxWL8HULMKF13myhB5adx6Ngz9ek1AYx+p7dxehpSRdwT72OFgn88RNdKhal
c1SSm2064j/TiYj0IddEnnQvTTRGs2vmRidQlBKk9mJ5IxnMYFSd0gEGXbto
+9BOpAJw8sEsQM0B09PWRqulOJfLQXtWkBXbVnnz1Njcfb6oKwA4x+PEmbgJ
mU5ezuTh0nfkneHU/iODHYoSwvsq1+wF3P9kTofe5T9/1j9b41aGV6HydRtN
f2rGK3T6qoX5ZqHigP4uvRVV2LEgvq57PyOtkWk9dw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RY+HiT0vKmr0C1BTdibIl991h/r07gt6VIevrR7sKaE2VBYcsxydskPnk5cZ
ZafwRWKYz7hskW58VRgZ1Ps6spZVvpJjDor7hZKM3STdM8QmuvxH/i/SVY0h
FGj+FTyVZTnEfjDOYgPbCbZdKHjpYpYgsg5DVeXO4cOW25vJTWY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
hDYHA/Bgm7p1lg2cLnb3b5OTM7HUmJUxSbZRNtUIWEtZfvklJJjlVtF34J/+
W6XEmzgspmw9Wch7d6pIGbGiXksp5ujTzuFljewXFMS1qvJHCUYqz0Mg5tOM
pfkzPp/qzzJhN+m4/t3OgA0ow6H7f9/FYdI+wPbRrtUNPKWfHJiL4xH4EmJD
p1/V3fAyBYDtYZbC6Mj3T+KPY3c/5y1vfyDYwySZoBWyTZWZSGbp8SK4u9S4
0TD7jnFWigSVjnUA0s2rj0m/XWCaTziA4D6vmmkjm1FS/eju8GytR7iL0Sap
JGB86pssFP0LR+M/t7Ms3mOZH9APez3JW0blH1BGNsrVhsBqPaGR52UfBsHv
6BxpffwsGb8yrtzlysfeSWLuzfwePAXm8d3FiwMELDwHsCealZuTA2kD2mfm
Z6ohx26gmKU7DhLLlHiovpVsfwhpDvWlDz7zt6labcyKxw/YvAENkwyhncsc
Aav3Pv5EmniBvQLX5+sOrSRfP1mwCH2K


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GWQ2KZgX5nMUDfVeL2OK8iWwpr+mSz5JLQbaSpdCxrsv6hC0im0/LuphiIPF
38jVt/GfYaS9mvUqCshNqRsZnIcJYINmG2uH3UU2tLH4EmSjUcUzCy15pYY3
59f1tSrr3oHBYGHPcwdjWuIrEA7DtLEqKX007wvjBRaWlyaIvdE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
WqY19QDAt3qhOl3VZXt7R8+mUEr1IZgFybstQmHJ0LWYwVUGvwE3OcR3yR9R
DIqlLq+Gxy/vZ+qINlcx/MOMz8IkYaFpT856CisNVURT2w+66CpJ/AWmh53r
prDthGjbYF/6Zjz96IfiXCpNQtmCKbAJcDCSv7L3MwiQ0KhBSJ8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 22736)
`pragma protect data_block
C3plQOzC0kZU1w4spgz3fcYRV3xVITI/00iTPzyRMdM5gdaK6xgSgvzyq+Xs
OQjefR38F/hET28QvpsQFILnLbrcYzjCG/JXmFb6JIRX5ViUuXBzcZRtA3aZ
HDyYJ+1HdEwH3KUvVMl5tQHpB4zt35D1P69B8zp5BVaPJMmAFtUZuKQxj8Co
9DwXvpCSjNq3844Li5fdvycG9Nc6c8+kRUl5TQ+/j0NMR/0oR9P3uhr+iA/Z
sDBEqwgDw45V8AOQSnp7TZzQufI2Ah+kVd0jv4oIsLk8CVoJeM86zsRXXVNS
5k6sN82/HuCrPLwLtlxdIPLvpwmtVZ+aLVf0uG/KpZqmAZ1tR3FOwCyoNkGf
R8accizVEofi73l/vnXcde1LNKInyl4DjTx8Lz2whooJzfwuVKgnvFDRtAs2
W+/Ez3d6YTky+uyxCFRV5vYluVUHn1Ua2qdw+HbQdcJD/xT+JNE9apz73PwE
RMgX5e118jNCE41zVOQno0yG8Aapx+dk3G4eumRxQlNeAB8dzD+csNChrePA
Qa/1lktS1H+CQWitB5N7UT6BnvHdpez/CxStawyndPpDiuv2ivpFOdrqZTKv
/M1iu9HybRHGLL73921BYkp7Mqm8XBsJ+6e8qzbbjwKLumww7KmYXDQIF30k
fVYkpAryKkUG5aJ0KB9KxTXHZdo2p4fpZCxCKgCwjxDgetxBZ+yQqtH/V5VL
fwSIzbmWLmycxwlKEACYFyxaL0ejLN9lPMh2KN/Gx0miU4+6o9Ldg+CHkdlz
gpmfZ+z/pcXzJC4rhwuK/OaleM5ILR25PvJflqWHCdMuxpefL+uSa14vpcfu
1HaRScJMlMxDtUvzBd5ZFKUeYx+yLSO/2K5S9YVQcjJtazVaiF/WSTEU63Hb
PlnkXndoRvPUziqrvE/DD9IWNpHmuO8Ts1RQG6WFXgXSkmEgiARHybLqx5rr
UK1EQ1ToeWxkhrU7JVz3EfBMlWYX9XJ3uTncLdw26/obX/B2bzknGKYtinrb
SVjS6aD1SL81MkzLEjouaGkXXzCWXsqWwM3c3CyfBTm4jMAxChl3DCVqpFwY
Y3cbukZLJBgG1yaA2o34nuwEoTEg/Qek0WYA2XSQmE+cMs/hGIE86OaoHNtB
vOXf3iBEnjxZ3P+R5S2mSlHmEleLNQ4SFj5roEXjcnYD6gmVLw1OgEXHx3qj
D1syyxegVmQ/O1ylZYgjFNpo6xtixfjmoDYxjmEM9X01C6LcEYN8wT8FnpnI
/7z/r2LqkvvUBhEfgF4AtNAUVkH/JX5KswMJ09YrtrvXuHT5KXtXJlrtue79
AMBgQCpcLe/Q2rsNNPmxQ5USOLQNxmej3qCvx+Y2AYYQkr/Wm/i7FL0nz+NH
OOTjNrOV78ODFAApAlLk/b7Pwd2Xcq/YAVuO34KBo3a2Z+tq7Eqc9CgKkSkB
EUQem+aI7XerpjrY+jFJwvoAOnuz4br+16sOm3MFI2pCdt7GUoV795coi+7S
c5LhM2nlkQDbS/GVT2QYn/n5fGBiI/GhhXUnRI/kbkgRcg8n8+6rkMK7tFRQ
KL9e09D40Wi2FFxCMsuqWSDmgpusBCno0ggDwv//hIRBsDNHlqxTrRQtqjC6
2K1rRVjxfaYyAaGw7GWisJuFFpHtnzWGLyCna3CDHOfzB0XsyLXNSSMbsDzO
FGdmd4vlk6mPcAMJ+b0qu1Mm78qeZJ3nzWKra8nKhqFfx3rWUOW6Yy/n3uVL
rb80sYLFD5S9DKZl2GV+6bO55gDX5xucGMShS75OvsQ4E147xizBmJUtA5bE
1yDLTxp01DbODaN54hnxv+BZp7hnuYugfU0BHGVPDoB/dhaIjIdCQFLRVO0i
NBQ3oIweke11BlvGtACCSBjuMZxqTZqsMc283JiY+PlEZkfWlxzZDRMUmxUt
Qhw7nrlQ4dKMoad61vPk/YyGJheJ5ZY+SA+wdBU7PozQT8IPysBoNknkDRnD
ITq40fuXmWSVGb5bBuNAfDrkwYYZii0406rs1slCRAMuupYxPKz78VyaaeQt
jvsIRMXpXZvCyTTI54JsSiST0c1VBUhp+RC9AMSMvIVeYww017AoNEIc5nP8
7qcUv0wKAlqwfHyWC9HCDMB6dw0TCXf5/hAFpUynXBf7VnbCceSQHkKzV6Ht
n+JFws8nED09hlZH6PuJMcPfF+eIr2A61E/vWUPx7zSddUyGgbmPBq2HluUr
AYfAhBMw0JdsKAfd7kQI43hTAcDlacbpzX/zGZSdcdpxzJrSKKX/y9juYHht
30xMygJ7T6hlRihxZYu++vsbuRovTw3pWGaO2j9YSTNTW/4XbuK0fjJVE5hT
O4FZyhN7AkQi8D7Z2pwOSF5AymzQJxqWyCWMHGS4+p4r9J3nydmTJWPNYoh4
CfgQUl/L2FFfFKXDCau5ytcGx1J3CDbTCQ8M+j28hcdNjCgFRSFIGZYwl+b3
hE/6waBJ4ToRPbI8n2HIrMWevj0fxJU6CUnXyxtGstq+n/nBMP9tF5tjl2vd
bgebZju9/p/LR1uU1KhbtuG3CwALobFTxkeO4hhjAWpX7mYtc5/Sa7gelG1u
skzDh9blVbeG4hR8HWf09c3bevHUnYdECXBzRWtKIkbHolMtSVAlBN5BdqF/
yRriCWPmAul0gicK3JeZ0qeNRRCcmfQ8mcwodbfMzKnnlXdB3HAeWJlzf0sw
hdKJ0iGl+Xs09RkYNNIIQPGP5gf0xHEWwlb6CJtTNi7/nkRboc/OHwRtSptr
WASXNpUSHgSdm7prWdXG3dOONqZFYCCRmrU6tT6FDRBu1UrcyohbxAJcO6c4
5En1kCYVDNdmcEvVbAC9ySCCWlx9mVU1rKjhgwGpAl1JxgNjB79GyHFlBPsB
lX9VcF3Dn+mMDJjgduKnA5LYC2562mIufSOm43qxE791JuWcafTwz2hGmjQx
jAajdWuHOW5RRp+fX7Y0+Wy3PynAAl4ImaHnDcwqVEvCveCA50Osu+j5Z6eP
wS/epweRHDZ+7tx1hWLuTHXoAMNV0aO1SRZK4IBDAtOIMIuqJIJrQXdY0jSh
GFZ/BwesSs8vSBwe8wYrftHKywlOOx1yA4wKGrCNP+VWAFjQmT9mMRo4ZOfW
Rp15la7ohSd4S4n63p+Welteztd8eO/TjDHRBtruhYhjuSmraQXiWVUSn8Te
9zCoWp6pyDk9PNyghyuvYZEaMH6uzbmDnBs8JyCuUJZkcyXbtFtrIpEkF90N
tuBa04iI8VvXePPO6Udkvvx/kM+8SfGnA7NBRxLHs4I4Us3K8oHkhUlPqg1j
qoXzAMgUyWbyPWCPFzeCht5S2BBa6g+IsaSIDHgfjpo7pj25soTg8OVjDsIi
c9bdMHz+5kHv3xS69O3nbmKaBti0x2BBYAXDbHmO05YGTikODFJAlqiRe7tn
QmDntWYFq2iv1KySQolw6gnWkvL92w7gewUl2jySY96EGZ6nYE1pd4f6Dmuy
+jp3Fr3EvOUcIJcdwzio0yvODi19oVWOuATaFmjsyE5dQ87wgI7Hv9YTUvld
B+M/NnLytmp3UZZzSsgkCdhUpa1JIDPnJwsezNPcye6Y6UnS+0dLOmCrZxrT
Oupe5DsQ1oW5iwk27hFH3PPwgRMzl3lrrXl0+jVyScRCL3HIAKEck820wT0h
AiPjYruijKQWqSoIxY4+2suRmbDbLrIUXnx/d8V1wFDIBL/xbq/rAaL84mGd
7CI4AIzdbNdvHgD6gFZXtLUuPdy0SqF+/jRMnuomNUlCk16AMWVOr8zwbDtX
3AAPqxj96c6rVmYl8Q2UK5rdebP589t6bWZE2hLCpKhj896oVw6zI90094OE
lhMveEVbjQEi208fOpFQzwKRrmw6X/emupYp7OUpEifJ848JfBNyLpLnMD5M
fb8f53KTiaTb4Wh3V2tQ4QR/xWYCzzoSY+nmvw3B0T1Sc/AWSQMUqPg112tf
Nt4r83cE/lXjc/bUGN8n09iZgiNVSaCXZDTqL88pCsb0jn7dc//t0pqXqtVm
V+mxVrp+wdC9PFcOb0CpMC9ZT+aJxbnJP/yKDvyQTHZOL3qoyTjl3ZHmeAiG
hz+clYLx78t0NFAGLkP2f3ezPLwWED6sXYP0EsXLKtj/qRGDy/f2xjhtWIsN
8Efv2wWbafuAJpPKBvjW9iM4KI6WK2LzkbHW4onY0MHqo8byZetWT4EK+j+z
MXyAhWHP0Z2f6Zd/rQdvS4z1Km1DgBF1cLBFiSNcDni7uymbYHc+vE0n+2Jx
7riow6D/M8TUprQlCayFqqV2MkC/59tHtsnQrofkoxHTuNDWnYsw/C1ITlsK
LpwNVo+LO+xzV5A6S1aL1fcWcSCeLxwBS9vZGczrliCIC1C081xU7XQIKsg2
lbofuBhblSi8kLr3hgtX2aiciatzIYUl6AmLcs9yFNSCZzpLJNaZPeBudvAf
2IRw+BJNQqUI+loQ5YrkgM+3B8V3yCFaJuqVycoc9LV572lpNgcQ3oUqahpm
laoa2SzKKkIyKiBdLipx64eIa6Tl/dENxlweJSPz6qqjX9RvLedVsvB34Dpl
w6Moe6jzzCH7NSwg9HDG5Z/p6/sef9Zc38ukHrBMaVjQXwE0s6IMvAkF04y6
jbGH9BE6NULiraPbCB9S03X6zt0bQZpU+9u5z4lZoLYBvg7PYZGvvpnjd1w9
H0j0zhs9wIXarYxnYY8SUgQ/dXI273rmylYkw0uxl3BWwEMQ/hhAu9eRWx/z
JqUsQX1oZm70vYLijcpH2cowF6PnmtZCEcDeAGPIOyrZnKXxjldYywGXT/SG
ObJoQvvwbPwGcFcfBGVejANCOPEM/Y5FUiO2bDk4b1s4VRfy5YdfMet2pSkJ
t1DKpnySqhLQnfuo5d29db+7TLDvUgE0helOTDVLhIbf9J5HnW+umFmX081m
dJkFj0rfB6/Vpz4OHu6gUIyOR6JoRZ7BUTn6/ahtcV5wPlhnC63wxu10VKFH
vnRQXdkdAXg17rchXcFAXCYzwZYsoiHdD3jASadzkjXihzEI6EEUnVpSduH+
bUXmxuI/geBuhywTNBoqtynTF+ZVi7C/K/+DRpPDR5WovdXZ8s4arYl/viks
SPhhOYn7Tr3P4Vb8nKApqB4B1RS7Ol0ckdKcsPNq6cC9D4XejJqBBQcjIQlT
F2Ue+kf40Bj2PfmT0KtYUQFvfBNO83ln5W4e0UKYp27GbEiEWCU1Ez9Fby6o
KKuo70eDF44D5rXrfGnsOPjbAkjVw4XLLbJU+qr07rmkt0agrt5ix8h7lu2i
yru2ynMVSy2rB2lu2CRwTjosFshvv4fDZqdKfdH20hV6wqFuDGKxM0ZX2pYV
xJXbqprMrOIGAdPtSyi6UFEXPvEMJ5WfIG2rT94xq/ORupd+JcvndhPi5a98
EFMEgaxAogwOhYsFY0gJg0m3CMTeWyty4Qh+uFzoWVNuQ+WUr3fmP7xZy6dv
MAuiU7yXQDlGQOHUBm8R5INiFbkNmZqVptVFtbD7Iu2ZrrrgGzeBVP2aw+Ih
f2Zum/Komu7Y4O7NxWSAFLj1OFCw8et+ptrpBjypiWLQIO0IAfZUVSv1jsqm
bzq6oVt/efXvdo1Uw3onJ/+2X56p+kGi8DHU+dtX5MBNfNpdUDUGWW6tKj9l
EX0KzeVX/sAb41KiavyoFYg8TKkw13MQ8tnJvfUKKgwQciJqW3oZt5Wv4IRq
vt2Bv8gLqFs2XnTCkCyvLIr8jtPuUsvfbhWL3VaBEMutENhIBZ4gYohuG54u
sCYxvthQMGK69i72vMgvY9YReESKPUg6DnSj88PClNIX7alAssCVuTyzVvA/
HwVhpWL6EmATh9bgusCtoJihsyMGE3p7qDTVY/WrD2uJsOGwNsOH5cvHB067
4ovouU7dG5LEA6dFVMzSvJZ92rlVaPdTXK7OJuDotgPyOKaP7k/zIhrDQXB7
KPx0IXhPvGctp11qTbImmRJB0wHHjJNLuyIUIP6sWrbIoU0o5l8hufKEKjqX
CQHX06tpXKKEB3kO5apKYK5vluAHC318KOgLCBqHDHV4HgFpGKWNO3Xg5tGN
LAeDSBai5L/DN2XvUxbpv1vtk2Sr8+lyjR/aqhDjfhr3YF9UP/LPv9mw5pdQ
4tzYp87RUBFr7ZS/x2Ka+u1aoVuOo4fiiypp1f0dnpo+yuVuXJbYESuAWNBz
h6HrfZsaE7YPhwECTlX1uIv1LntgpWsHcypa7F+C5YAGJnptUVT8xGp/sOM6
eio2+WFqsWLk8q1Hm/OTiVGt3HtOK/sdspslZzBrhvVcYr6Trj5ty/qoKJic
LCu1bqeYLaJv51KrJi18i80LRDoOscz+HNYGOs5SppUgTH3j4Wk0qBEZg+uL
xjf+UYyAcpqqWbJbFduDHFwVPBCDLCJzR+y5N6VzIJsLGAItjZke/Q0n8Wf/
mCDrn8+LjEYJzubL7A7/MaB+3x52Lolj+EqLhEhQso+D0XfbbkRTLF3Ipvaw
wrHRKBeoB2Of7LmBz/SSRZWlhKpuMgcpAroMeSKB3a1KEdL0VHXAwjr5hsm+
q973gVLEDzCy0kDqDpFgfPl3EFS/FdEdxz8h/cK8KvN9hxzG1TC+EYdhccOY
R7edivTcHtgUpz83VF9qP+6At59e/K0rhT/0QRxQU+rLTK3bVIp5fRYBu9O4
r4keYTGIXXR+FLxzvHTQ97CAHaff2wJHnD3hbyqY6f3hx3XRkrTRNtow5a+b
hJmxqU3g2HArWiT93k1L839q+92k9LDqcdfX2Ne1w8AR9ssL8MqWLRbEhHF8
AV6mVIVOOlSVHEoHz/44I4auWjDODSfNtDpR+coNcg4Nre7/htfG+hppz5PX
Y2OiFeq4jwojWabHAinwtTQjufN8qFbjYh02OZZ6PaHcIrOnS2snTnN/Zmkl
WPKcQq1SQyD/ECv8D2rsxOPzlRHecg9wL7mRzSfE64x5ugWY8PaaM3DrZ3lD
UrffCdgzLzksOvhAI2EC5gczzjFslaNM9NgSdT5KeBikCDlpJSr+kPA5Q8w9
GCnjsPLJPyn6FOquaPYumLNZ/C185O37TObZaHDkHZ86W9Y2VME7oBPUcHlI
gPx84ru7IlaxhUxP4dlWy3qP0PlSrcYCQnxDxjI5I3D6re2L90oqetkk4x+h
tb15fa9ZriVjbnpED9hnCIJac4qfNu3F0os5l76zUgTJaa4RSatqxjnm81sp
X//yD0yGryRdnYUd5Io+Z1k+hZJfVIy8TSKt6SqWsIxHPOPglL3hGpl7r5Hq
Y2izf1iyGXAQlyQuv+3eAr2UiO1vM1chKlGsTLvh0SItZvUefK9XONs9oGt4
5SGxjkRVBs4rqbkUljAuCHFwho++rN3McgBAv/N4VCliEPIO/Xqanc1douEd
YGVvMaT003eaZQ0eig89jzHz5QmmeHauX0gXz+0EkAzLmf9b+L0rr+/Azo6t
PaLAz1gpUM77yYlqXlmGHmXqLsDVcFgOTDgydRyTJvuY0MAnaANfmOl3w3aQ
2ZaX4Fl4sVVGQw6IzpKXBMJUaFh1KcZtj8TcTdKri1+r2bL/4nBRXvlMOh4M
iv0e13m/JeroVDHccoWEAwPqe4tCN4odViJ94Nku72S7vdnrcvU3nwDFZdv9
6fcqSjvBapLtZvakuXCaa7mPF/+5BxMGA5Z3WojZhiU1uuOj9LnoRw2cFBD/
OdwiAFiVoW+i7KHmp8lyPn4iOirjBAvj024lPHe6cl5KUNEK5qHbQPm63aXA
dlkJ5YCH0prEMTqo2dKl/gEDutDrYDUGt/68IWeJDtroyjFUQ1Gnx1CHS8YT
mS8bgtu4f1u1lJrP15nmELn4vcWb6sGYjaSO0YwFmKG7CoHGJY+eTzIEfm4F
UE+2kD8ssuMXMcamqqf8eumTmBjw9ZCyuTQlhyNaT+RUjOACKb6UPSiFMsQw
kLnqgJ1yD1ihI/BNebj+fKpQwRo4VLNgJ28NQYMyN/Fx9GEC+dpH4CnGzDBA
VRfjjeuwBSj85uOggLuC18NBs5DfVYIScU6KrBHQViRE/tIFI7Sfq77ZN72y
QFzX7V87X4Lb6Dd+TlVzy/pmHkuKYcPmltPLA5p99nxAJ0N08ROaXy3i8TdX
ofko13jC8Y0VOhDa3zBTsVjmnbyFeoZMKRgNdLPrXdScZdaovOmbnacqW9bm
N4Pvkmgjtwev5t0PxGDorDTx6t+V6GFH/OU9xMcTRQostxHa+aMaW5ZbvfaO
9q7fKyvF0pwaofzYSkxmxwMSA1LEomT384WgCX0ClDDmHijKZLtRh7MIQmdE
YiOo/miJXMrApRQpo4UWd3c+tS6IACJZmfXkIUmleA5GtEFJt+2g8Knlspij
mxsVvpGrEARYTd0qXABb7xO5IR6gzO4M8ueTgubBMojtbdoPKjqpJUnCN4fS
f2OCCehynKtNM3d7yq7WZ8+un682bEDg77TiSfWcBWOSPq/QKEjoNjEw21/d
UNzq7RiiXvRRTZhnTKDcuHM2wvwfvoovngK28MxPprGxxba0HUM0SNYliADu
PTsf88tzIRJ37UwMPLY3EoFKO+PIuXZ45l8oAza2BG9wmGT+shKi+EC56gp6
2OdvGp4RlL6gciOrrSYmlbTuWlv7w6xqPuQ/WDQm4yA+I42VFqDgRimHFcjD
8aEbDWiQrgBKF4usnlAPtYPyyVIV3/+Htc7AqgUJxxFWT60xm1+o9Qon4xbe
fDxpSKelagjsbCHMv8lfZiNaZd/5gKuDUcdnwhqfUc0AX3eciklbQ0W7OAMo
VR6qcM1mn7Db2NJH5s6Jt9cmFBxUN4uod6rAfRG7V+XNndqBMOZI83/CoSdD
HEASzxl5UfB34GjBl9stkhn3EAnBrkJ+/N/Wur4ZbaRSIKvj5N6YbpEc5Evn
Ccb0Y1KvcF8Mk9bClnesB1mB2gxqZRgJYFJvHvMuEPUJvr0H2Mk+mqztDzHC
eiu4XMgGK7hPK+E62J88DhRvftns21iNKJGz6qj1ABw4UgOWdfomXdHh1e05
fmdu5CCC2htylbgFg+IcBxV6cHqUBIVaKYXZSn+8tOHGFQoW/sXXQe/fEjn7
0zAPzqumhcaiEgIAIB/RAcpynEJNq4XDW92eypASUvV8qFw59w6kj+miGcem
Dk/CDz2mjs1YBWscoH+U9t3twZXwc5yQn0LflWWuxzjFiwrhc0ajKNgaa2L4
Tc1T226gy6l6qR2SbSNgtnZz7H+ZYUAWHUPKLvx+EkOjz3/gHrNvoeCh+NCx
LSzDW27XSsTK32KWrDWxfE0BQ8L04ykc+Tnc1IV62DSQggxfGbEnVSsyAf3D
Orxb/jRzwDMImOYgBN7ZaSWqYzs6ddquQ2RPi9bppEHFB1jAGjJqIu9Wo26y
aqXvnx8PB7RzZYb+1vvmk11oDmNT9y4QAQWw5VpfvdHOEcxPR/agiBNe1S9M
UeuovaN6yLFm4w7bE97XxK+nkCZYOMHor5KlYpomsujujMCJUKANh0diWZci
VVBbgHnl+PyXlRIUoSd2ycT8X5whV3nSdEEL5c9NTtvINzV4mYfVVizUTZGx
t5SSkliq0RH6vqqqzAaM+YoQ6V9WCFJvRHhrn4qDDmeYRtoofwDO8ppJ/WJ3
W9K7W9PvSQ9bZYZN7+C3dmZV79aNcmY53GBiXaTz8zn9P9vRotjRq3mnmRxL
1M9wpGuplvf9jPVuhl+QfJOOC+m9P+kB3sFhVK7wVgb486S0pkPCKvqlgdsv
qYY9iWhxxcW6KIxAHXXRAEpW2kd5Wy3enLQyhVTLEGn4/I0cj/oDIW+A3ZIa
q5LVc3zpEJ62K9r1MqJ/M0HGS32sjaTwQtumiD4ufhV/FlJz7woTIcOcN6Bf
gyvDH/yxeCsgaj7B99Vweh/7qMzy0oBM8fzJT5jkKY5dwq1oD4q6dQ7WvI8q
TJMpJJ+tw2KYcr9siZtTUmmPOz9duBJxuhlOm6urjNPFua4+vpXGRSfnDlzf
4yF6SxM6yq+V78LMlPfe5+ilwEoygKo77jOERPe541iUiSOP+r6K9favDo38
bhPearv1YAHKRpugJZqXrMmP5jBYDVsboNX8rABKbJ7DCaraNDuKJGVOSUy2
mgqpob9wuIYGo4WgiH4eAtKH8dJAM92oydaQka/NXrNSwqykLOSiDJQNCWhA
38wonuowc4BwTYg1zyVc7vQo7Ao1PKT8or9KBm+mK8jCZFoQdetjwqacfh4E
7LswnWRZgKHa08OfXu9QgeCWRLQ3DICDr7tPrbOi7XkoEjn1XyxRRXzeoBzb
k5V50a7I0kJIMuMmlpDobuqq7OVmiu/ObYiec4Duotl3c15wnSVdGkN4TRf9
dzRswd4BUWgDGH6SpulPJ39OUo8yGOLA6g50jWhIsiEmFjOBluZeBZ1asmVN
5VRwRuyapPTHNMHX35h7sGBcf70JN6CSoRaGSYpQQuJMPX5jVdKVuzGtLgFI
ghdEnT+LbCTyrL/OQpHR4wdK64y/BlMP3QevG1m3oSbsSY6DLtTMF5zZd54S
ncDX9gB+Q2Jd45IyKqANSeuk9J48h+D6YHy2XEOYvNNeMAe1EBcP2RTfcvMc
5E/XFTUtcTg05Fb+CPvPpqn1ClP1lRIqbnc7Xh4tB0gFHjbQsULEMG/MGNvB
r9xqqEVLdBqt3lcMHcEnPIe53x1Y6oFqQ6KI2JvgHEClOZJtnnNUsYWUwOKA
Ba/BvKaTwmVul5cgCv6lGqGlcut2A+m0Z4bgzR9qo0BC8uObAwWqWTwpf0Hs
c772zKzN3qKssQWv+UAipst8FZ2xF2XV21jjhTRSefFgRuBhCj6vWZjFQrQy
w+Ev7bJdlBzG1rZ1HzPK9FAp3sHOgPHuzqQ6LEY/tgILKpqmmh3AHtyiX+Mp
jcdfRU5x10AL4pseNaxx3rcK6w8b6WhAdkuzj/TKaTGB8lQI2yI6Xcm6bBRE
FG0KBQoWZnM5Mf1z/Isnoyf5eCrPsQYkZzxZcDzCjMc1x/r4i6INUfHtST+P
2bTXdOI58d1EAWvbI06xsC1u+QZap3sXdJyiwH/QmXTQF/GfFlbMjBscKD90
qJyTwe7o/fKOD7YTL5WtJtUSE+Is4ctM+Iv0ZENT63F6cRLHma99xwRWFYuZ
XJCZObtz5maAyEZYoxFaMztjxvsrEgR5gPTeQHljmr3ccRQpP+uAgLQGaiHO
750ZeFtyqiMOIrXn/TeLsjzuo/k9bwG/cCpvyVgyX6HK9ceWtig+WaRPO4pr
NGhZArnZakJ874utIlt5UNkbUxlgeofE5JaUFsvf4nCm4xRyvyABwFQerAxp
2IGaAa/SC63E3zHGo508IeP3nhAa8jPfG8THLn62mt8CFb7cPG6JKGzwUK4t
PapTVjd4pVbs6jyi6CMGybdgw1FOe+ND26hUQi/N3i+AnS2Mn+Fhx9FhE4O2
P39GNXojAl6dZnb0k1J8Ye3SAwh3vY5aYmg1icBFJr4f7nHFSzdW7hkqbwQR
taEJfnpmGHArZnN55fzTq5aPXgLl+6WKt0Sir8hyPs4g9XOuEJVnv6Mrwh8s
SsHP2HrYfPdDggfwvccxZYMkExYrURlzr2g10418gEdnXVJNtRNS3bhZLV42
bNgiXaCC0FproLteppGS1cCMX/tzEpQRnWrKCTAMB9cMa4FKD8MmDxJWit+O
vYRKBAi5500KKkxP8PX7xxJQq5Q7cyLQZIpHvMC+OvOf5grsXMx4TocuN2yS
vhUAiSdIxzAN6FZb2r5+IlSO0QLEuUZAmXlYumFjtkYbn2cofAHPl6w+3IDA
wEPZhn2FpMLCwJCwUHNOyJ7QpKX1UCW82C62hHgz0tmtDLHv/Qu4SvrVS70U
WXiul/+Ce1MJFb8s07TFI3En995aby04lhIrfp87qdKSEAZx3FTXTMwnnbFQ
k0qbfXmnkqbepjiUDbhYNNFfVXvUBczsGZ03aDjMJjt2NCz0soOiFsmdNRBG
Wwy4fkSuKMu1FND1nwjd6kl3ZjsEwsIpLzG7MEmyiUlbIfmxWmMq0vc2BQMr
mmwx9Zk8s/HyhR/hVaTBAWGmC47I+fDH1vsAJaoq2XlE8aLvj8zbpgXzNtN+
UpREzdqeb9SZHDJPqO9J9sGhKjHWNRyWpD8GD0OFA3aU1xJOrGCU0c/m08O8
ohQY7Jy2Z1WXTZQRtnFtygclWohwBbptktV6wEE7eceTS4Kr7UGj0wa+XUOR
c2Q1GEzngY8JEbvHfhU01bc7FqzCVR68B4p7uywBx2P1DXmyd5srTDZRt6Cb
mq/18lFqx/QtbUP/sP6vDUAcZcCRWDR4BXMfYgYN4UUyEUAKZUz9wZftm1vb
Alit6J1MH0RJlrk5Rf2F5+vinZmhS0FIm9x5bAginKv7cs2cOYMdjo7fVwRH
PrkHPmqRDM2iA15ee6C/634Jg7x9NMlVeyDMynSUeU7t9hIP/fF2EEKBvdax
kOxNfcx4Y1RIyYhlTUwZE9+G+MpXr5vNOda8dliGVT6BjTkrt1Z6O4j8gOB8
bLH3JrqSlUQ8cTxqXEAWsZ0X8HQcBvSQTlIBfzU+fhxcQeF5WQU1eXLVKYyM
kFe21098hKUjdlnYDQMg8O5dzXsAt+hLoDwxoK88k6HaXfsz9fcwZfPP5Nfx
mG1gzf7pxVN2/eKxpx61GC5gxdtXTFZh/PPHSN96bGaI9WeDMM3n5fU92dTA
My2Idj3F6ZJmgb4YUO90U8xzR85oTSl3QA1qDdd6wxvmCw5gmfepR5QuDiZF
eaE0hQRQ5Zn0x7qezXTKe6uyiSWAHJIa7kHYU4LtU05Yo/6C/Gm7elAnJM7X
hWaZs8Y81VB2pykbiFLu4dQsjWvfiFegHb9tXJoYlfq7Pr6h2FmXH0VL3WRD
elLH1WNIdHLi8dPU2sMe8X4cmcJU9Znc+XONtNwzo3eFuc+rfA3H8i+G3hxN
QKWq0GH3gnVAvraA4xQhhW8nb9mIzlTD8jpdJGyAuJdrw9IPcOn49CkTGgq2
CoSjhV22FaWGqfG+wNNZyyhkyAfstrEhPpmCu6fGcabKJCW1noXZ1itOfUre
DruxuyvLy60pYf5fFSln2S2YOBOvezbv6JneYbY4Tziixkn+etj1gy1c/0dI
T+oXL/EX3BHVQqhefPlwdInlabfIQlSzC+4dIRELOqouEr08/W8cZqTBQLY3
fPoWTdBYr2m1bFUVFHNglqUESB+A8MOsyA+MWLkLAuoXAso6CpViq3zs0Fdx
m+ZoG9BJxzYLdyOwZFO90LG42ArKJMNiibL4OBMOkfM8j67nFbesJqy393+M
nr3mL/OOTxoC65LNdzdSt2hnAaLeF/l/RTjm21XwGcoh831HPCpdCCQPPuhF
52fmTR1tEI1Fb3EYb5LD2Xww/6KRVZoWJYdB39CX2tVFibpCz9YH45JDUl2e
+G6H070CIFg+idQ/AozLt6SkjdVZ31EgrfhDeLv19sRgaTZ3UjvXib+YWTrn
ki+ze8R0aVn63MKLwXdvrDFRc45CZFqHctDhB/PnujQoL/NTaQBxvOsrFphq
QCdVIWI1clIz+ctOW4KJtkrnuAMn34FBuh3lYfgRhGy9oLfzIyx3ABZTt9cl
NXzceMAC6e4/r9xaqT5abT1e3PsQWPqmUEJWp7bhJtbpnyKmIGondTVPHGqp
SaAbaKwbACMBK4IQJCSgLNMa/AvmyV2KbQag5tkl6RCjhDwL27OfPq8AySkC
Mr1HkJ2TeXunvp+t4NaqCbRwuhB//cvEMCQAWPlJlGN13nCribnhz8XDjvpg
RAcPjlVE5kaq4TLbohH2rRVKhZumpG1JmZ9R3yrtosnpyvilXMglXhgN6YO9
zMzpI9YabrpbVBJALjZLfn8pHxJ+LJlF52KookF0buyChU7xQv4qpJFKJ3zC
MqZVIHilyV87WAuMV0EjIywzVDBvAXWjqPO3HRUgsH4gxg18AiA4O+qKoHJt
EnCQr2aSKnBBRfUbYe9WBlS0rFvunUoSutgYtJVnmTqG7YEel0Yx35+GH9FK
SnqkrMJJ4tB6oq+HSOyZArrDWUemHmag4bKdi+65Z+Ze+q1x+IRw8vsTfBAn
ltbsIAPQtcNSqiUPYHT98BBJL9ATAw9w6urgExiEAslkK1YcJP0V8itU8W4D
Ess6i/ygJUgnxUf4A51XKGvhK0m/XDVNSTisd7YS2Q60+LiyHc991FkzY6dX
oB9/4dmuYLU07YBO3ytBLdn2ykhEOgzMvdlM31hPChhQzF/kmFPiIFZmHALC
Q63ViE2bom4JXwoKgAJNorCvZoUBGdC+tcYlCKsQFHJdDefRn6OZht2N7pt5
UHYwH9+FDGhzFPDOw4LhEk8XtXhXopXdyzU3Q3cFsDMHdwY8YE8kpUSq2hhs
P38EQFjOp76LdNfMmxwfbsZJSPFT6yBSlCV0KrHQdf0xpsE7QyGSDT+5e3bt
iJtsbXwL0tqczaAui4uBDNsW4h+x49q0Co0SAcpXJsraFNky2ocIRSX9PQ1p
LAra0J49B/199hOJLr5OIS4SyVRFTe3SghOa6PFVvamvvxQ0/eJb+wHY1Qk3
M2tULLMClM3YNlE7xdmC6lIL2v1STTZm/adZveuolOy/PA+D2yPMGPgsS9jZ
7m1R9Rq8KCIUKB2TTVlR1CFwNN0harcxxHylIuO0OAStGMcONuLAaEUS6RrJ
zcN/ylJGHhmtNYGLXBUPyZT8gokBUJcfOXsBswJVRf9gBKeaJjI5zzQS7v76
ugy7AatnZGdt7X3dMhXrTNFf8Lu2QhnrsZuTB513jxyYFm78l58/pGAqGGH4
yYZHQkMTM6+JFelD1AgVek7LUsLOSR+DmehTC1Ldeg/tJyQ3yZjPzqYDHaQU
kDyN/0MqvHv6lK5aY4pDj+WFc4HTpr2BverD+Le25rrDfu7OkxQKD7iyEK0E
wU/Ys5HQosU54y1npFB/vfuNHJVpr1Tc/vIN1Q9snyi/3/NevLV8zvhaADil
0s+5lfhT+y5rM9Rw1Ctn7fDPIVGGraWuP9Muu2vQZoyVo4HTRu2ojz9ohESk
sEznnkT9F0Z2JhHGs6hQMhwSPCNfJmQNUrxv1nkQixnS43iTwXzPsJz6V7uo
H5I1YbUSHGm7TfJzRMPoKUz+gYsTl91TsDcetvSjoryPGc0668wd7f+VlD2x
BUBARpWLReJSYIJ6VCyAMme1+ttX+K+hwEBHBTIr3wjCljuIE5192ccz+fzI
o8UZIeiDdif+0b1Ym2aE0ybF6Xlh/JzN595mwW7FoI5qNixJ1rCMNWFmVedN
1h9KFHDxgwTFH3uQfSkyeZ/S2h0RzqYcPIrxSrzbrKcfN8U79g/pFqDIoeT3
B5MV/KfnSl5hBFZqtfsutI9WhKJt7WlVbi+cPsmm4J719rc9oMCmxfAxPeQu
Uxki+b2XhWeuzH9K1vBgzd/lqA/iLiOlGYP3MKge+CBdOGdsaiqbBODtfggx
vrcH3C2+QigpgvVUyt8LWiZGlH5O0A3zU0c9Wc5/E4Zaot/1LIxNt/uWTKPx
nzwapI8ApOHVcaDXJ7r8ay5cn9P+vVxcAZLJT4iRSmiIahWmdqZ+IQQCafyT
5mZThldHishHpznM85iUxkvGqwGrUrLsVG9H5AKWCeZnLiZEYMbkfyd949Cr
MaTtksZD+MQnq9NOyntrJcUc1LNxdS1PkGlRWSkAVAIHs1E3hgzKgILsyarI
zIssL+h9OHwxRSYwyEiyvxusANMEGAP0r4OXUPZvZOUv/zlcZ4NTntCJ6aTB
JwvHL2PM5Ohz523B35tcBS4Ns+9caJX9TwPAUi576PrQf6ADEIfdhELwJe9w
76SYqtHbrqaQY4Wa83DEvlxbNAlJKs/1+q104/7BNAzXRe6Z43k+hrTLq2Pk
2TYNyJCW7FLrx8cb6etGlAxA6lj49NVGm9/wbwSiXIFXG19QVr+gjTP1l4kg
8n7Qc61uTjm/D48OCDQzkjFmsOK/9xRH/4JPFV141Wf3bhgcZdg8GXMqbZw4
fp+Tc1VKONayhDadG5n5m2EnAIznQFLJ9dcgMIimWErTMUQTT1lOF6TBl43k
TUWOselRul5SZcuEooXtpiptRahQWEvqCK2vyE1BjSGOW8gol+Z3HCLpdraB
ZMUqvdU+R41pJYc1sEMrgxEiC8h4amD/4glm30HqLMe3vnJWU/xcXh+lj+do
H5gQ+Bu0Qhtv05CL3+H674oUZ/PfuwUMiLtxMtTfFxH0Z3W68Z7d3Ym1jH1x
39CmV0vGX4bCFKYAaVZRuEtuySRHaa7utf3UvS5e+sDMT4kYA2b++MMlK1ej
C5Uw++Uv2gX6oqSVwH5C5Fj3uZlC7eAKye38GK536bQJLu0EJ0jX7maL5086
ZHN0llmojCqpgtzd6MFHaM2dioPl4lsgkGRBOIPvnQgHH+YSXPBiClBVFkam
nFC5oM4lDoR+gHujCe1udVan8ejZfsFEEbnPd+Dg3H0paH2JnLWtvbP+Nrlh
Pb1/OwtdeHYgen5l1/s6aQMchJW+quPmTbo6rcU0rc4NmXWsNeZkIlrVnJ18
UZisMidC6ACUQpoB/kNtlJTvcdH2zEvbmuRM4wa7TGr/5VaRXpN50bExKa09
Sivx/vT5GNW3Yzwq1JLq7yS2z3I6Gh79IU+JdzKk6lNpL/m8wtw6l0KtmJy5
UmXRmRWX5sQtAWPAldxHZ1aJu+kDwGvOKk5qHhvELZfldoXHngt8cm2vk65I
Dugsd2PTwkKDHrkBtrC55T2rtJIYPv/PU1xORnPeHuIDqtvhVMpGHobSs30t
xWPk8IHYqO39YtLw/qGid3DrR2f8JEheeOOB+yPNy2iMwIkq5F/fz2tiS1Sp
pzK2Lwm7HWubFnffqT82HuI6p9MOXic2zGAtp+sZ8Q503vM28GgyDoVGaUHR
mffilHCjxYuk0aN1PJGO3z/4KVmxIjI8vkLKX0sZqTRGRzOgH0St/MQPKjMk
Ux+tSx3uV5aOMU8irTDrVppdDGYYefIxWGh5EXreXBK9x8mx7QkinAeESgrX
OFG9XvS+yZFj40KnvKrIskWAT53MLnUVKO7RdjMFR38ZWTZIRlSjN7b5paNC
lmqu9rwiukRju7Vor8HmSdJiwSzro9go7qfr0oVkytOIplpnUzGxTvgXZd0D
MX+HR3BRO7TmnU9WwHJ3gyok7koxLIsGsM5eiA5Kzlt5TalgfEx28qkOjRow
gLz5jxOkvbPxdt33GuHk6yt6Mr7nMTOoXi7YG11mt8Q8DTIGqqmzWw/jdSp/
pAnGZ3cgeJIaLCCCLITqQBZXxnXMkwv6Ck/RK8kK5gd1/VyPYqoNFB4rMWF/
xFKV1Gdqz+0AJUM+AIWMFj03SnnOkLDN95vn9m0+/0Lp9rc73TR8wtP6tky/
JR6QdvnE955I8tk13Mo6PV/BGRb9t4Ue7nD8XDGoBcM/ALTDXfetD3DyQnwu
UxkAo8nZGhSRcsxIX4ScMkH4J4ek4HBDNoOi3O11nZRcj3iJoyChsq4r2+Ai
lwO9dSURLveMc6X9NQr/c/NLpEob4MvUMc3L3+K0fmtXFOngcQ0oUwpN4pS+
BI/vXwkkbml35KsUiaM/j3RGtaOrUNYvCaO5MXH85NEUIJmJozO9R0OmhF0N
FqSUF30AK7qKBdayz0kTpxY7RJsgf32Own1MqdsM2tW6Dn0wojL9l5ADt1Ja
MbaRK7o/dP7a03iT0+7Nq8BIYJQ9amRR1udTPUqX624l6Rizeblq3i0ICm4q
ChRJEZH+y6fmfVNRJgGINrgASknXNUhqzMmizQEmNfJen8dw0j/v2VjyU+lW
0igoOcIePcyM7Rx16emWUKaTvFAV3asT+S6sOXUt3Eqi4PIKeJVbPYJUEdiD
/Y/8dv3zLzFsjsRlQqV1KNfHtSLbpcNM5NiuavjGOzwzmBrxaUBiZDB2eJOD
r3haQw5c2vFGi6WH9e7prnsVUtX9tZE06VV3Xw414N4SeLIf2wO2rENkdD97
WecffUXMJ71ID0wy6EzU6GNYr/cAV2chf6Zti0eAagfMHZnXsKSf/IX1nstC
uNrrrVYxEDGnJGX996E34Dn+icaDfXNPZOjm4rvCijzxJD5PFNWCvl63FhMI
LKjeWyF3/htDq4VYaSWfjQTkNcHut2QZWYGjZUKKBwi4VnUB3AGfu5EoULrJ
EqgxjDZSZmX7AqyPdw7xMUXHjXBa6LFxoF96UmZ8U3os94XllIE2tnY8fvy6
lYWbAxcf4N9ZKKvrW5M97OkOUt3dC8O0T7ITRUg4NG8oJkj2ho2RChhFIRYZ
LuDT+moFeC2k84EijRHiLinrK3aLqJ8qhCT4lurTL/YUGgtryA4GLbk6+0cu
G3d0auybDDdVCEfLhVKN4MZHDHVPfZdvKWC551VPOAn+SvlW/x/GNyPw1DlF
tTTlERZrAfSwdvvYJxQNUOadEXQHhn9cY1AWBkryvKkSjlfhehgtBglEpPZw
XkidxsO2+a1vrqV4Z3IbgoyGR0X6r/DgotfaG1K5LU/ddYpNzLCz0WI/E6w+
LzBBWN8Cf2+/nyzccuard0Caz7i2hdCsgEUASssd9SyVsuJH3cVAmmKaOzOM
7UkB9+pi8JD767p9qUGN3j5jISpXVkieXYIOLMskCF07Gi4wjEoYpj/oecjW
njj+DSie0H+AA8gq5nd8LB6LrtB4IVITMsy1d1L4GNVzlFJnFcdHB0zxjp5f
d1eRI1O45NBSaKKuU1ZdN7+UOuEduEtFkJUVer8pRXgjnk7zvHONWjZPrBxe
K6v2bYhMf1wwXuDA9Bk54m1pp5nJPNE5CAzTBSUTjc6XAc9sI8uQHI4nQeN3
HNQaJjxaI3fe0HetxIsaGFNggzwqsBk1PdfXs8GKNjQsNyVO/e0gjHoWY/gH
JN6gLaPimYcSamZ6paYUvNLBTzZj6kJiv493LDvBs89AzDp3NPP60xZX9Y2Q
mtLYgHrApVbjAQhwE2sG+3anl3qEyc48Pnj9aPLxN3ZWC5KJf4YmFy6KCc8Q
5orfJhFYdNa0v5ZRY6ngAMdWPscpvMoSs9kJET4MSicsySNh2Wx8WhvxWvFP
OG5iXMbBue1Lsn28Gu+lyyi6GiEUAebPsk51lr6NeRgvJM7NJcOU0u9xR5Sk
4WuJnKBjZfz6tFwcHd/zK0k2rVT/61H28ItFJgwSD6tdNY7IFKhgwqZVHF5k
vo2X240YCLDS/pbIDb4z+zbQ12e2Mt5mnmSyF9H7IodlWDIeNXD8eVifltLH
5W2TyxCAXs0+A0X+NtFAGdWmxSnZ45prVHlmb7hSl7ynbraXcpu1/f6jRwxx
efp7/zQJKvyDxBKMVpm+LDQMRBbGmlO/l5wySSAubGJwc0uOuAF6B5Sxo6B7
wPK+S/uoeacktLw+GcEIDbMK60gDRQrmkAvRDWHG+/RoPi+2VbXIb3MPMz2L
KhN0uMiABIlx+2QMjDRU+weH4nvsCsAgkMWRvV21r1QxzCXHUj9wLK/odx9x
MpdPrCHnMTB4PtpG4ACBUVoNgdwbB9uRfEjE0WSuNt/CW6XhT32/IZMJFL4W
Th0MOz18VvYoUHs4+3WU9emYMwLUJPuVBvXHIGb1TU3iDP6RR4nxnvdyaZiN
TxDd+XGjNAWXZVrfsoVNCiynMMeXx8cZ3hMtFPLq0AevyUIC+RU2R7GIbtyl
uL00IMUkw6wJu2V3RceAwdCEM9d1U9fMg/nuIFWE/V7AVtb3xKWy0TeoNfHH
maRhg6QnMq46k8/edKzs/J0hwBscbuw0t/b0SzP9bNnHDQ5pcHDNrdLQcHph
CmRAQmVhSbgnaKWBR0JrsLzJxOoaYPrH4lqVbIkJT8XWB5TNFnbhL+QWTMBI
bI77TlOEVnsg3wQQ2F2s8SwGabKero2WRSvczFiNb8wm/TTG9KEi8kahtYEz
Bx4yUe+ayd43J57k5Hw0p3fW5/+fXVygZjcEr35luYaZSYZLmS5azt6fnaSW
RIn44LncBpLAinYy0nLjBFrnPpTj2JP85064XitqiDtzX7NAabvQIhZ0pbFC
W3bZJGoYbipLTstwmcgXirt8EgPS29oo9Ji6PIUmcxdUdaSfG+9dRtbB5GNS
Ca4ZQITPwu4KPE0VoNBx1drtUKcvEmC19RYD8rUql5u1UevM2yMWayED8Pw4
+WAhuLWz5OjgPAe1gwmV0sMX+p15lmuL1bE2V5WFcLaQjTwtCDs2Uj2kKSqN
ZksU+1+FzN/1QFgGAAhywzzm6IQjPXKeS8QcslEoUmwiUa9s5aMVSk5RyScV
cgRh93nh/gYL0eWwkBDKXG8vvU8ZFI3SosNWXsruPESw+feYKqYn+6B5q+lr
LTIBeaIARNBiQlRGZ8lURsPI2n5n1MVSmzSHTcBQ1rRdsov8u+LGcuQJTGZ4
RCy8leoZcR71PG19TmJUmzk4bQUhzlzII5i/YsSwnI8eVBJnuoyOOGq453vg
mngeugkPlLMGobxJ4h5lt7n6Hk4+Ewd/Su4NRlqnF8kanYVOJWj0d5FcmK0B
xeAfC9KkuBkKwdH6i4I/dtFIaP2XWEgMewOnxY1erZPlteqh8vBh+a3Vd55W
sORskQMyp7HAvuqwUP6Cht9wpGKxD7PriKm3k8QTE2mSgaK+I5DccVCuff6z
V3vmmSCNu8o6byGT9qBLVDF00lLJ9NUtbdEWtOkRJIupz4bQwq0d2bPSMP0W
er3fofFDaguTXHjr3UTKvjaiemwQ42x+V+/6AxsIX/0/KrVTKI1ZsvZE5mp6
xYA+7+FTjVeUQ+i/KSw3Q2aIkRnNsI1ZtNEPACgVf3c+qOQNY7HJ7JcO5qR0
AOY0pZXqi94XiYD8t9I5N3xMZ4NRJ75jSs+AeLmX6l6Sp25JUSx64m9x3tn2
Rv2c6sT8ppP0IdKrQ6c+M8VaZrSURhSBQ4j2MoKaauP7hVufpXRVfSSlcZk1
QRV69LSCcTaWmP+TM06ub0/OhhxhZyrj20znQvxmcfzzjQl9lC523TLHBD6W
UAqj+kalBV1WVvNA3LRLrpmlzg1t+SRFlcPWlsRsilBwe3OaOiYHRk7YcCyI
ekIEvpNF+8og+PL4dYwnL89tNeaMVYE2yVHx+/RTRE47kLHCmNN0K9XEIXz5
FoliorvqjX5TfzY6OgigzETVif04I0Hhorsnk6ogglTOon8R7nsK6PQuJAG4
BCFw5XzKWjqWucoRFRV5zGtB2g8eTMj4DhHmlfLWgPgqoRmwA5OGOz1zDSba
+HgXHuZddU5f95VVMOjKWztZrh79ALIyv5FpirOOu93FIF9jGzJShykvej2s
+xTPst7JuOl0jxKzt1ILHVH/jzBDB1pwNb7naodDG/Fex18jM1mVo7bQjMr1
lj581T81Uc+cnOr77O49jx+12b9XoUzXUtyrGROQWNqeLg72oiJKEzJfPaoQ
epUGA3Gsij9WN9XMapnbQURS5urVFw6ZSouj7OkDC7iSy8BZXpyg6m+tSab3
lxYVZ7URNWthTF1Gq/ne2tIFNh6r2LYsu03RssMV50jXRHcXjDnHZ6FrT5uh
8FKcrG1KzuPwvoqbkZI8p/mlQlh98RXxRBCdZ9zpiR/ZTHCJ0Cw5GTwrnA7l
Df9cnSIOIE6c5wamTNYUhqDE71aWBtDS8s3tUO7U7YabeiwDg2ENZUFTImAC
LU/rkKehkLuB4sMxo2fqU1t0mpNETgYMPf/ykaHBTyW90tIlDXAN1QjzKHdv
T1r38akxQRqesngn743ltj31kYAtwnD32Ui5rmQujaZ24/s+aSjFT52uAKSV
PfLB3Y0+c2q5ByayHg+YpIApFWIRMzKKtiir5nZ65DY2N18NKrdTfgNzCjUh
MIGgOllrP2YABiu190ZvLBtpVhBw3M9Jw/oA+5diqBhOjFsPilRwS/NxUKG8
dkZFsSPvEZCgiRkCqIsSUg0c6XAak6UhAsP4zHUKHyua8Ko83GuYmie01dTZ
pZrBahuAmIGDEMP2rqXuTFXEXvQi87H6qjOyloI776NXGMKlcu3k+XjC3f2H
vEId3bWW9LwIcoswu8t79Mo1Z/F8BYvKAKppW5AUQirHuN6KxF8QQmzEn66j
yYH/9PgcAS17dNwvi7GDeDMd1wFD1tR/u9TIMsUfR3ThGOVMf5QRLhvB9241
XJje3mux2mG6FAqhnEWqI5X6eTRoxCtF8c/066WV9tJ8ErTsGSm1YAVNSces
FJaG9mQUiXpAa2rTpAw26QeSjRnOaf+bqvAgcNZH6He26RrMP4ujFXLzHlkh
RcsKcGvNl1YxXyYexqr1UEhLKxZ2w8Eh5916Sx2khHK57sUD2psPGOcTretO
dfR16tbVWL53CAwgpNQ31T+gVX8WKiB2Q53SYXZ7WX80nK1JROYhrusbETyg
upIMO4hbADSstHDiblvgv5T5iOZNtaU/v9HSkaldQu/fbQujWkT+hcG5N88F
zV7hlpjvvhDsVBGDntXCtiEKTD6ZA4BDhxsIABYYiffa9NEBLm0uCoM/sgA4
wJmnBC3POpmRWJZKJaQcmmA2Vpgd8JV//cXinMEf6985oSWg0EPzlKrYMU6G
hUgfHv22FUXcTERxpyDN+B174KH25ji5O+/zvmCuYN3ZOJIXf95vXAkGDJ7P
7hl4vXIYE5WOfRLZyZ8SXuwpYXEEJDhH9Oj/hkvnIrv1zdR4oYaliSggqa/2
wEkboZaHPSZu+UPR7L0WiIfmW0t8y4W0ZfD2tMccKolkFkm/TfKmU3mmaN94
PBmr1yrm7lKacUhBk1YyHRP5gLLuv4fGXC2SPVGTCZKuC8jLzCrMdGfS6CNh
vddWrWSPITOCOlKJ50venr936VVfaeLWMfO6p7A4ce56kX2V/ufnozcivH4B
teVtxw2bKJX+vJ7h4NURSZNhFtTFrSx3hj3tOHNGXAjzzpuus+6RbrihjJif
8FnIZ1O4NLRbP/aSinjBctMThkJi36VtTA5JO+XEjuggGwNOvI3UwymKP22j
e2d/iwkTTyjVObhbzz1YzTUcfG4L2hhY0l/RSkGVNC7aeZ3ftgMhs9yopKFZ
AYn9je7CyVxyt461jkn6Vn2Aizd8twIdu9UHTaNT7v4X8ObbMm1AQbYrVWk0
uNqgQkpj1iXuq0wldzq1O7J313b3X57mQUB1dvR+MSXRME2uZ2uOKc1zk8hH
Q4uLudiIgxNRbzQLINLqFygiIA341W+uj40ZpdRB/64uxPqQttpqJeD8Bo7x
jV5p46vAt6tmL22RB9pq5jsm1bnBtxvAqdtoPJSUT5kCaXmvMZicDDsUIPup
RJ5QdN8xZUZ3kVv4uCPhwF4YCQZMcQrspYLml0tvuZrryLU9LL3bNhW1O9/e
ZgRXTSuIr/iK0ichTqHrDlt3y9QWtg9r/zhVRXZ7F7aNoltBUFd6t0vC7ofB
M7Kx7Lhs87+hCbHT4eOoF+03TERJI+uH0z3by+ybh4D6EBCs4ylhs5HfPvJA
TJJmNq0GCIlbV15OoPFhjw2yELvqAarlSu5rm4c5SiSO8vP9AhNH6sshWkWj
fIzLxotz5EXydN/duKovWXmzIz56PAu0hGUder8qb/0GCm25I1oqsjFBjGvd
1kKY4rymAI01BvM8noUF+fwwtC7XyalIDQAfo+cLB1qI5wpKbYV15dAjqf30
n9x+uA31NSMlmY7QIRPT2G6MWPsbLCY3HcLAmcnXm57iq47Cfg8+OUA6FuVn
A3w5eU56JoVLlPtUY4MTuV2coKbtgfk4JCxSXVOb1l16WkswjgV7xPvaIkHY
A9olDf2xLOU4H7QgE3RKjNy91ei8QpaCE+dLBEG7uQiDS0jBFPTKu5b1kSIS
kPf+uoAFQxof7+xKfQsJZAza4DJNvAxu55u+gYtKFNEmw07ErRIO6U79wn7q
3suTXSa42SBBP55jSee8PU2Ah/SO/p16gv5/Kq24Hbtq1qjfF0IlMajpTdDa
6bWAakA/PZLkVhqa0DlV9wbSTt4ztVedYQ3SmbiGXk33wxpJWoiAmVSfzuHC
CmELckJ1NIZM5bfBDvjk4/CU/FkWpx/i0gbmjD6kzanMJRCLiqXqs+vtuFIg
PQHGFnDLyNwQj55+1lunWBgIjZPGitqdEmy9zZsPYzZ61I9IcPBaMPC8SqWM
LutTGaqSQ9CqwM89jEUq21X9s3bs+SdEyVoeNlO7kgnjYyfGj66S7/Vn+0Rr
hFlQDLmPkUi/C0e4dc9fkZaMHwXFkkSsYQb2ZMAz6ZkPQG5sW0ByqgorEHve
QFD+POloyL2x5j0GPNPL8prRhhDz+jR6WzACqPH4iTC7q1b6VOv2zmOZs+M9
X0NMOXe0EeEbvn4v8tJopj4owjaWUEC5IWef/NCw41KGEHnoJIgOmqYoKDJp
YkmR4edglLPnRk9T9CunMOZW1/+sFV+A+bS4rjvmFkNtE7t21MpKe5Eubsdh
fer8ROmnVugqNdve8xJhrk59yIzxba5TA06Hb4LGkdi7AFre3jGhOKXD96sX
ceDD3xhGS9+dKSTtFtOIRpfcD5zYKZbovGswMatR/Cg9BFJRB5JgvX5i8jfD
/Pgl9mjlJdHDIxkaQ1EUO4/wE3kp6DlKD/BZc8QtqbRYQqEwwMKNF+B9vLbg
RiHc3n1pdiSnp//G0guLvS0b4maVck3LzWBc5kBaQ157M4L7/TFaVYT3lbhy
YDRyX13Fbh7rhevH+KJiS3wIlnZUUaHJiV3a/djxpZz55wBcYuAQgIR16Rml
6XhW785DiXbKsEpQjgUlBRZ7J2x3HjO5dvqYMqLsJUP1tfWE81XzA2l+VpIu
OkpiRNrKnmskRjZczJi9RvIBP4anO1q2aIr7kkVMgIb4WhJ3TEnW5Ys7oEsO
2vV56wUIA2Zh8Lq/YWGf2eK/qSBU9mI40iHa2XDV/n+LYPrPjdSOOwV0CseM
k1w3sTCPIkwmgJKlJI2J8GN4ytkBvrFLambVpsPdL70Utg0TnuPLadsOZDWw
3wiFkvBww4OHmz0Df1iRYXZyjGmGxoJEIyaotkkpBnjcRy9tA49Mc07Uc93M
pNBjfMWZHFRt3mV3zTerjd1uyiHaqlSa3bswpVjJvLPXIz5uTk1drhoZ+Fl+
msg76j05xs8T9SLAeVyI9k+GXLGS3gS7HWLUqovDt3Isn36fQ8u8sJUyj95H
P6H39B3Ry3WsEUy76OCG/SjJ50pcmDfoiWUsLA2TYeHd30yXg1nQ64vGrbeN
tFBdpwI+z5JddqAkB6/U21TkpXWhnJxE0t+21RzTLKMcNeY7FBkIdMuGFlde
CiVu5KEWQP9/sGM6EbLySjEPwQzFXG9DV5wNDn0Caa9Qg9xWnciBzYln5uRe
hlnJJLqAiAZDNzYTq+x/uOyb7kwJidOKLGFMwZLTMg1YvCaisog1ALdduE1r
wbFK+peyPtC2MuLkrc4nxEe0yd1ul1gyLDSvsPNuGMFCSYlrXfI4BsZM+f0m
wKC4Gt/XFlJ4NiEKEVt+JakTQsORo2HDhL5U07nSluS4ICgEBWfwzOjh/8sK
6OAdaJ+CwSjZeuCtqKNkQn1AVK0ki2ABB+JoCa8aPkcFLPbcjn6aWAnhlz1l
KLeANVSq+lX0Wb+qBmzdm9DvoQ1mGiZjcy9t6tOdi2hsr53U7IEFLoybhm5j
u2gr3BMm2Sp1NRXGLAJe435cN09RsXPUkd73JQFAmbWrKDKUMDAv0Fe3VHfY
E2/Sm0Ks3jv2tb265fw5owIrOV1hIjA0aadV+n5/NE7s5VAE8PG/FV6bhmLn
K2v29ls2nnkX9PezgZSp31FEBDS6GTAljuQHhjTpzhPA+aGX+0zN9cPBjCHS
Kv75S/KboAiavBXifQqo+OqVev2MzQFczlvuh8pXzvUEesw2sonIDiKQWSR8
fnaY6Hbm1FuJ9hRcT4Dgj8sWtJQ3ta6XMHbec5OwT8DYYEdGOe4mIOJduUa9
+r5ECWEaaM5X+S9QbeEycGSLJ+d4vZ6rg0quI56ZOHoYemj0lxaINcVxsrRR
AKiujzBtTp+DyrwYjldbA9NcTAP5VLymbpgmjH/TbY+/ANpc/iQpmZuaGefw
hKeqIoS+o0L/syJeb7Rvf0jWNaPBQkYzm0W9diIMku2DxZYcRaN8kaE6FMNb
gLdtMY5QRBwVJO5bh2K9i0wfe3dC+FTn6PATHMFXG9H51ETFcJmOWGmmavBT
eSOB9bitkByshQmBFjiPEwp+emuRIsFwdmNtrYSnpOLrufH3s+MVMb+knWzw
udJXbPnZYgSZatg7EFIMIlI8eIQL5y6ABNDEs7jK5UGkFtqB0wbw+6R9yUPE
r5GGvYPWAW87b6TY6jASvbjKFjekO6b0J27AnfjB1LTNuGpd2yfrOepdpofY
L2YX8r2PKAcBi0/BjZd07Z/6U5g2VLAFzemmqrDkaf6DnQGehi1Tm2x620w+
e76AJzdYqSYhwYF7upUj6NHrjNW0myxMBVAAf6ehHSuTQAZFr63/K/EYAh+D
AZB1UgZzE6V1i6fxPRKgmeuXJ+OX5c2pRLi7FiOkKuEBEEM6oeB6gqRGoI/X
w4f42Y7aGd9v8CcyGH7/D8TNDvT5gbf7p10PPBLlOY/1xxfqgS7a4t6BYKMR
yJdpX/o8JFYdouPuAHZzPigycPPYqKjqoQ1WjM8Vqyz6zJuzppK8sGOQxYhK
wRWcFhkajPu2ZsjF8Q1i5Ae2IkOhT1rtm0WNL91vb/rwordCHjWZSrzyViq+
mlV7md1OluEbTvHBV7Db8zub/IWlWABGw9dR7i2cNnccfAhZuDvfhl7Opcc1
Qe2MWEa4qQRO+h0g+bgnFsErxlo+HU1REcOsSa6F10xTK9J0eKFWcyC9kWmH
bIWB1mqvCNB285+p4xuplxZRlADepEq3cKBsXvyS5U/JiPkVpdPJb3M25Hxo
pe6tuUJvb8uZfSbNXbYs5A5foF1YECW4+nAhlJcGtKacV7s9J4Gmc2bMkR6O
jLXqubmubhQeGzT/VWpgwl1t7PK4t6QB3qsHL/oRfXzgvwypwydZ0AYUri/e
QZdVjCIrmi+ku2h7FZEQB7zCO2Sak+P+OrladaaWo3BeXM0S8pLG/oAl1HnM
z3AlcEKZYOMvZgWo/DbPLAMs59zzkpugss6rL/F3q5k+P4Vee5nFjlZyVRyJ
GHtflni7HzqbdqhoxVckZl+HpCAsHEZ2/xGNVe70hxxoQSAs6NDmCq4GtOjt
l/8J3MyE/AA+Uoy/RofoddB2W/2Uimug4MloKVX7RetFlSk9S5JEUM4QKxN6
3jVlaGylgZQ30D31vSua/h79MFqKIQ+uOSfPN/xtnHSOdWqje2OrYTsmAF2F
cgKlfQr9v6Sqd3t9B98FEAY2CxTNmceAmcQjd9t63gbuTHqZMh1ZUJsjc9Cu
IrDeF0JNAZ+UWCOfXmBDtK4UHxT4vtkBKNPoUxG29Ifs6c7JNtfOZGflM+MG
4F2bpqtl08dZEHi6gsk7+XKOUjW7hiYBuYDqnFXTnQSQp5Ip0eeyb9gpLE12
azPq4he00mGjPg/Ep/J8Tlq+rPtAfiJLulqyr8waKWU09mtlKVNtfhyNa4Qg
aB3JhlIdEDuRwKwVCpBkJ4zSdwMTWUmtq+5yvPcgbGzlUJ4pDvQmKkA9Ggyn
QW5x3m2EizRr1aqfn4kiQLlw2A4zOyQMKv8regY9mHmk30DA5dOOxWP3ufbj
JVlbmcbzaZ80vhSPlgM/tYtYTF5fsH7xOKwBQJqFaCpaZdqcHTaLGB527ybs
fInap1Jij+upv20de1V8vR4WtRzvcwX4ryBjnnCpI4iTpLIrKkyjozHwpLcz
fQzZYvYY9U4WSH4oelmJFP62tzAN0WtarD5f2ldNZ5ofD8bbQHioYSzffN9B
abI+4YC38/0cnzOE9KG6eBnfx2JUuX378jWMehNj42TzS3ISKgaflgefCF7l
RLkWJCH6DZexG+Ke7QL5uHlkMCKMqaWaJE9jk0U/d3Fuhg8C6yuyABXkNde9
EV499MtU1KQJ+QgB5i/wAyEgiOFKUOnPpi43G8i0B/NR073Fym4wvetIA2+L
Zj8ZD97dKae9zj9OUPN8xdm5iY0FUOPExFX1yfryi+fyj+RAzVjwsw/DcgnE
N9m+0UsbF2d8jSLGM3dPgrCIDdtD4ikx+gak0Ph3v7eOEGw+bz3Yt0alZN7q
8IJ6q9fdgiAKoNhWiwFKm/sjD6FVbCIWpSQ6wrEYLzP2zUZsfg+BoGRNhjRm
W/Oh3RvcMssRdGXIs+goFC3kMS0qgKboTrl1KVDYRHY18yYxlKiNyTznQZUU
ZLGGWbg3juqw8qvpwCGWkYZmp8h9VvYvgEhugFu6Q8ZQhZRodtoF4FkbGTug
jYkEM6yQWV02bYr0A+1saGQTI0gFTgDN0kOQxFJoZDyeReDoZc2Bb6vpyhpe
v8c88VNzpFSfurmijQMGbxUDHVYjV9+Hpd+1gQsCm+znXorl9+CfwOxWPd/0
aenb0h3fLccCAZq2F97FGxPnQ7hZdZxGDU6kWNkN64tORdLVNOSWhXXc89Jg
9OjWxboxvzftdO42gL5/NrzEMEoO7jXpJWFgwAEDRzL3Ue5gLbIa1MFX2gQN
2Kn0oWS9alcVquBMLdqDpwOUTtpqIFFgevI9vfjwhzZVJdC/R+7w2JHe19tA
RiiN1i0tOYamGMe7QBbmOcyA295NijYs4fR92WFX2cZpkLnpQGeAa7QIIPV7
UYWtIodEdjj2uFcWERc2D99jkImgim0JSH4U9+Uj5Mb/CRWIW3XP7e6DJSM6
v8H+vc6+C7LK97vE6mbHajgcWafAT9icRgKSBDqlrXwMCyX8IbLBaz+GnODU
UzCPCQDsiA/jHKpx6+6jTHo78Vn4wx+14jGDkHlKbutcYLO6Z2KqbzDyYL/e
LcqECLqvIYGQTalekVAcmENF0KyK/FsvHOSPjQdkSEfHxF9w5jdSS7jqt8JW
qbePpTPHu5rAsdTLcnrmkzT6JHAqI0TZNnW28Yrkx7n9mBvTO6TzQOlppUsp
1JUit0xPHJnRUUyemNXyBFkvYN0GsM7NIZO1XNCE8ilezvIwTkambB6g4nzv
pjRgL+NTgmH3F/tx6AQBw1hRz1tXOQjrmGtFqNjRWxRLzfhJKaa1i8gyTUGb
Dq3hD3EpZ7BlpS07voKgfoP02RsnwWO3IBM3cMOiuh9ggmVlRQK1YYBKLkGn
aizW/N1BlDArOSOW0e0X/xxwossdGfcFQaEZbuLxh+a4dZJk+PebEyWPVXVz
x+LGw4E6ZIVx9bSR2yuRT/FFKz5miWJ9BnHv3vBavMflaHM+2aT+ER0pJ78q
H+rpp2xtEl0b7boGjypsmipcSZM7ch0badDj3o5EdDE/zhoWa9hT7/0lxbTX
9JgbQ4C0fYi0Ms/fB0NWhjXwV9tcVrFV4WqoPsG53cccIzCmkKp8qPthUxh+
NxBXzN4PzOs/XFtqcWLO0uH0trs2ylhnbItqf7xMZrRX5rVo5HPHjgePpyos
6GAUnncb27XTgJHD2z4PHjDtXPryug5IneZh4I2Ka5mz2uLPk+3KMF3PZGHU
+HJjyHZ5wX9AEQMvHamxsYyDyG9i0XK0iiKDjsDHYHOquy+3HtW8XT8lIeuI
RSgTferjEtfEz5oc5Ll6pVIQN8+PyGviQ5z2T7VVaZSA24Dk3QTrZ0tCOMKd
pPjWICOUUrmIBwlpq8v1kvfvbe5X8JxT/yUhgbBFyuvQpW3m4rZDtDqVaR8I
7HysKlqyW5eO84J9ACYwZ64Z9bwB1lG+wZ2kpya8QxEdesvZ28XfMjzeLv/g
efy1S0vt3eLbnXScpO6lEur35PcMCjusQ002tSHp2TIHnUAqN9NkJq4w20mz
11XP4N3Fmdn0/PFVneIVsp3BAJeamMJX/WFcpyUhdM6iOPrTAsZvRB07oWET
uqFoZS6et59QD+Y6qyBKqOTy884uoMi+L6kPEfgSyd9KJpHpJ90tUJDgGhlA
1zk7CjIF59KqcOaN0/w6MXDt+P5Es4bx1dwD1Q9fB4kcFbWugMbZvS2F2IS9
MOY0Uku0VtVKAkF35Jqpoka29d8UFWQ9m2F/7edq+cbhFnae3RoekSx9/rbo
1ZG4XtfKKqjsNQdl06OFmXqISHjb34Xx0tQSP0K32u6HAW/mBfUrgZuw3cax
65mzBDS4FomDOecwJhk/1SUPBakxzhdc2cb1Q30UIfA0hxfQJiwjDzTWWLU8
ya4Rd1woeNHftbUjzmcsBsFxkOayvk9BDIw01YrRcIXhqIkxsdpxMxVVKnjE
Ev/a3i3lBH2g86rzP839UZOf0w5hafln4tlXH8QocSFnLcCovaXpJS4tyC9Q
lmFagjqbvl7pwTE7olRnZIQwz2k1G8JD6rxNvTuYxcyYwvn5possbQW7EUnQ
d7qvJdp0IiPOT/M=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzc6byktNjvwFKcwYum3Il62AdamnkVYoOH1nO2TvdKiSDb2wHT65vjsUldffqrpaYKvU6kgHGjidZSCG94n66FgoyxJJ9YJIXzqrJy5qXXcjorXzgs3+xPrNB//Fz8T4QfEH17HL/gDXhowo2/9hL2mdmEK5bq/Zg73OmKq+yclwNs2sfVmIWJUknqFGtHRq8N2xQCPvePCBRPDqjK1ajLAElsa/jIsE9mHx+hsiuVEXQbWtG1qa0HZO8nFruvOhz0S64ZN8kIo4o+TslJ7r1d2GQomOhQrbdo8JjN0MHfMH8ySZRpkZqEc2t5kJFa2Xkg/+Cn3B+bqbUBzE00gfbbf52OMtiHyNba2EEkv0Xae0JvaCwBBMUJNYSRb+dtL+/0OhJ1/odxIq6k9J6m2KnKEZUOCfb9ThiZr/hp2wt3C9yZ44Fmkj6Hu0DeGJ+KETqBC8+ei/hzFERX3lecGhVIxl9y7BGwFJt0YTHOEKtomvTO65dj9DRNFdtCNptPB4DQsnSwHa+nQgfYYxhV5E3hc6Gko6aJzfQNKREdKyk+XEAbvQw+uPXwUVsdyigV1VNODUZF8RV1147949dMBHYK68jqrX+bBQpor1/0lumG4vnNmAlsYe2zJ1hiuiMPiFCDQy8UloxRtwrEDYKDQk8JTgSgSeTIWciDy97P8AjPcyuRKAD+sN7D9HS23O1xpN+KO1FUS2kMxx5LIPZInx7Mm/w2c992Eu3kMtOsiuiPFF0GTi9RfPca6jFeX13KTfjwJzzGCFgwfT6eNlpjmRG8H"
`endif