// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
k/jo0rqIT942gssnbadml0wL7CcLHs1yDw/CgbMdZDpFZiDi9A9m4X7Fnz5x
zl9fQTYUk97syfg5Sb0Hwz7vUw7vhAKzBVllGDq/LBIzpOJmBYuEjOdv7Ogz
bcNYuOHZzH/QhE+0Rh/EBaiY0yse6HpRGcVxJ/j7neRecFrGj8hhav3kWCaT
4iPw8Ihs1XUxlBmKhK1IsqmHXpfgW9cWE2wjbRWzQpUzUNYbV9YMTRxM5JA4
GFHcyIfz2j0PR0D34Z5WepQCBLQww/4myW7WX4XPbggncJ6BiOVNEPyj9lNA
X75einWc5O3smnCT9nJPtdCe/YblsNgGuztKgZZsvA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
F+Imc+g7Cl50NemAOGa0cfQinxIpTOhJOHBmmP23pimvUvbsSLuxEhUKCcsD
n+ZQdvk83sDO2fBVeCf1LxitEn95qvgmxZ9fZmcK/aTejPVTSx/Xo71SQtwy
O3uwzfZ89X1pa/ZGuZUUuYCd3bQYx6qagm3IdL9LA3a69kvYr/iQJHja9aFc
64FjLAn6mqhOpV0KYR3UP2yNzXz544nOOp+fRQrS1U7CaU3oA5NfQCwtswd9
vdI6lyjUPhAnoOp97+98E6PVL4kW3k/0dEVKYy2l8exQMM2GzYOBiaVzAFXK
FbFH4Xlk+ackdMFEHUAhPoL53iSP61CPVFRLsN3K7Q==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mAP19RxMtG1G38yNfuKOylPeK8vJQ83yoqNv/vm5eJwwo3mzcmxu2QDhr1Ue
T6vGsKJ/q6+JXH/llQDRGVeA6lXvPn7/WEWDhFit0d882UhLG2pYBsbEHuaZ
ftm4pUMxvQX4D2cz6C1J3F+/wt9PksiWliKwGiMiNO1Ca1Xm4MPYlka2PB3p
X0Hc6V+IUHspxFcNE3e6bCvMj+yqsisVXJuMlbf/hGjx1df4MjIXrOtNWyZd
7m7FqoE7ahi7u29TZNMCWON1nOlCfMdMFKj8TmpXo8s5scZvVcUFn9U6mdni
n11399nUbV+9GqZuE5wdY8vkIckfXvSU9/N90/feLw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
e9j1ShmaRR/2Hus8a3Lfj2lcrP9QQW9WyJkA45WONXEIW1WcjP6KBGv8qZNB
3bjqpt8981ohvwhtkoFSTYp9ENk+W+l0p8mhf/DsJxXTO96EjHqjzfOENOPu
tZ0y5dDuIlJ2XNCnwxLtv2ioBJ1ZhavLIiKiT5MtbpGSaHOXMzY4Omj71JxB
2eDTum9ogXWcHCNB3ZgJtiFjEOGm8BDfUyMFczdExB/57ef8NL9yeyKuEiX1
E/bYJChvf2bjKDBv6aEqo4JkO2CR8lKEOzdKuJhggmGIcIUtIt35eeZfxQZh
BxpS8IQcbzGyCCONfKLx0gCZ+4wlvkTf79K/WSK6hg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gILeXnSE7exUtxlkAvlaCuy+TY40n/CD3flGnI8762B3TFPPO0fI3qmZdp3N
5igY/5VhGlcVGHNb9IMVrC1T93q96oWwxi9b0O94yXa9i1/Xh+DVrol2RFG7
qiRKJMSw+RqbtzyUjHw33HBuT26y5qRV+ObdXRtt8qCrckrOxhM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
msC9kbhoMdn2uKLJrQO6nazPqnByLXOUaXBnr9wult8NWXmu9r/G/yA639jx
5KBbqMxpuS3k2NmnTNlXnYnNmlYWnu00WTSU9WWc/g703tFEK4sEI79Jp5lr
VTiy8f3pPSnYGBS2FeLWBbw2GBt3orKfO1HN84AO25XcxmgxxDFW0IUuBKBI
25uBtNfY2zYBY78jo2tEURkIuB1PcLaP+Eu7kCu8UpG9VWA994UL7F0tuhBH
B0D9TAzu0caFxY7yCZS+cGfvxC+GkFYoVZ0Tt0iZN9ZycYsqyPrzol21bA2E
Vp9F2N2B87CFFnK5KEXpUz3so4/OBiDc6/w+GC7aViKCNMe/AuK3bX1wkXkV
G7HdzBDO0J6ZayqlMZx2qoMurrs9wwvSx3bUim4OI7ProswDYcACmG722prX
H7f6EKtgIgbFEXIGLjLl5MRM+naK+cNoDzSYjmXwdDiPBwZ8rGHQQpzCkZxl
FxwxK2xLyJ6WyIuYEHmBOBBlYVMLtE18


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iSYkjZg2ykYhYasAbaD6mM+Iwz0yOSXCa0fGPQDb3yJ59ANVxtPHe3lmp6Ro
MWBtMrz0qIOljDxDTigOsoFZM1fGSQxkbvJMZ/UfU4iKPXQM2YjBKt2RIbXp
GOuKSAGzGQdA5+sGwZ3KGu4LEkcjflFWzU46DKRnv7sDNObqaCU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
drybah0ggOrZJRwFawVyjfsRDc/6un6g61c5ysPSjf/j57l+MH80RzDAJ8Oy
u/XwQlGdSzjWN8pjv15rThmIcQm7SVbqjxKeAcb1g4luu0JEcwG0kviEsmZW
RRVXZVi49ejb5Rzq997KUFlw7IOp/D6PSFfggrouFco39nTXsvI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1312)
`pragma protect data_block
e3iMfuTBmUMshS3PFt5Iw3ZmCfMI+w7h8Eqixp4j2L3oL6nlHbfSD1RNC7a4
06yffwRa1ySaZUKpu/fFDDOwm0HDkyd6IyFrPnHCbwyKg2OSZnXiclfjbGJY
+TgHXato4SaIZtf4DC6BhbURmzXkDNgp8VK1zL7kBFOfLipS+k3XMAyyL7U9
xpArzCLdVoW49Zhhkg4X/3Vfq+pDmpC2Q46KCkbIc4HHIAoh30jwJ1tPYqm5
k727h7Gekum2aO0c6kfJeZP/RpIIujQMlxazNFePUcSC1I9qfVNrQ667BtP9
aGDKZtK26kO0JHSU/jHg5k8t5HlvzKJbf2S8/zPkKgdKo/eRG9b4qf13vyPG
u4hQ4jgCHb9IXeOAT9JcMpF82HSqjzDvFckPNLUzXq46SaTK9SqoFe+8dsjO
gR7xXueMcBxAwkExpDO8fDO6pfhOTtkIY5sgSlT08hBfggbX17TFcWmr1o4y
fjN8DSkEfk/VFs0g0fV9vyVUyRg5yXo5cAWvxx1z79Ef/Vnyyxo+f6FpGLJj
hSGEi98eQBZLpGAzm7hFcfBmw5LcsHxHttIjMn93j1yBJNdhZz6vF/TrmxUh
yH1nX/uKPV/qjHV/tptuXegF8ejwagkwBRePAKcDKCixIF31qVl/5U/ZzJVu
k6vgwD8CPZ8UC0/EcK9FFbAs/6N89lDnLnBtxnqVKaSgdch85k6wSWV81a7/
pFdThSbfNB7ll3NZjYlwfF7WGttlZPMpjLgi4voH6WYh7vuazUZ4Ap/Ad56f
4olwbteTca4ZaJOjuJlOoGk3bsXDkyAN+wKl619IqnISZ6ErAIqbotPAL2ss
Cq5anafOtz37JpAaomE0Vpteh4aYhnrjL+8ngkNgQJMp+61TlkzJlZJWPUKY
0+5sa/trB7FZXQZEAmPw6srRdlVVBKtrP5oQrqxtAFEFu1QuoX6qVp7dbybn
202YL+yVXhgkjliTb7Sv5tbZom/oaLbbsnYESHo0tmt8JvOHchpUe7gVNw3m
pwOafboVteC4DQIVUt32zYjLrTDCJRyphKp1EiTsuu9NbVYoyGV2nd1Fkl8s
lSbVytvurtgOIQjJADtk2ZdSrLw9DuXWklv1SsA7b3+ua0YMVLG0EK46xpDf
E607W11ENnHKAoP4Rwss1lliax8cDEwyehGOaD5bZBilbdcnNovimKWuTe3l
vor5jzIbuaNdBJQnDPekSq0H0dBaHdUSq+fyWA3VA/0KhfD8woz6ZWCjsu2t
E58klLkSKcLcxIQCtg3TtZUmEvRUhi8gph/+s76bvrqW9yByW7l8RUh05lMr
LSvfWX1C16qYKf7DVqohMg3nCv/Tj/x05hwFvfUX68QwJ0M+6u2V0mkVu2vc
hy5X3GtIFSHLr/ei5t7oQIuxsljGk3MfYH4/q/Wvr1R3Qwi2rnZccpGh113x
m4k4MQ6k/860xssKF8wCmfap7v4psNUP8vctLjg/NxbImfpbVpwUqOgU/4R1
+HlULy+tIp9yRbEyAQ9GhVFgp5z2qaLE8IhwU3GZKDa5t6tFKU6Rid3Tt1ir
UWZl9SwEW2YKU7Tol+g6XrNdW8uS/ez+T5vtqJe6t2ns7htzHcrznV593Nc+
VA3C4NnwmXLUe6SBkyPtkQHqmYcWhV0zd3K6RrL35A+rJ62cabRmcdCc7MSl
eZGMZl5+S5gVNkYWW5WRuJqVmdeLBLQlje5cSSduWLr7LHeMRIg1qrCEp4hz
dV/zFK6sCQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqelRvBNv2eVlBqbGylJVV5eSm53HY1D9LEFnQHRaOd2gqcyf//XFtQ3rNOtSHjWHC+MptTs/rKBPzCvPLhBTVUYyCpBw3mX/PrXucbn4kxm//jmThZGnAZHmqK7x6iHaJp5+jMXQruwu93b2FkOM1gUdIWnOBFHs4YR39AX1JZgc6E6WiETietjPBmsEPH3xz4aXJTXyWbXd58pH/dt5LdP+hYUTs3ketpsBj8twVw3U8KMhnntI4CwI8oS+7V5JnNC0cM9a1KyCn0MxKBEugCbRL6bUDNldVScKKZulx7K5h/GNWidMJ+qQRRS29AvWm2HLN17nG8gOqnvqw7V+rVb4K1QUMvjR1BKQMBhPsGJK6aTbfBJmqxFJxQyQRnrQp/WfONFWg3ENd0cRar5EncDs3iMu6yyhwtUtMzcGYnvp6Mu/w1/tEGZ7mOwPIfqCbcZduU3B4mjySnLiggPv10gJfE8VL2NxKduyrDK37Rdw5rs2Q57hFM0T/297D6VhxLyVxewaskwxHiAEpQK87p5GPnhxGgLjCknBKbImZ71/hX3jyQ1fiBaS5H3OlMa7RAFuk6kf8RVr2Xo6rlzzZ1gD2STNkmcxf9sJaY8CLLLAwXP4s+QR/4A05EqRBsZ1KEX8r23WAHlUBlMpQ+Ee9NqSZiWkHginu8fRnykCpdW7SP/4TbMJJ1ZfaPUEnM8liPLWBCuStN/EbG7LR1p8UJb7BwYmmvZTuIgqp79vdj46L2McX9rcMAfqhta7b50NtvbtWU17QZKCedCBQNLwiyg"
`endif