// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hqtpaCZVk5AULHVJU47Vac8rRAxA+XGVLikOoGVjAuaf63xAICqnW1pVXEoE
wXeRrPd6oaWcd3cSa+O++1oYUpVvfNoQZEHMR/fz3FzkFJx9dURWi62EcTGc
rBtPfVm8TRKoJ7VO1om+o3+DLQwo9UGVhMUU31F+ZaW5zQ1JKPFBVYmJsLtn
rNqV+BpFkJYEwrjNhHOV0utObqauBtQyPICpHVIwknKTOjX8In1Yu2pgy5V8
mR+0gGB+6SsuSSSQFFF1O/Q31qJRFiJl9GQD19YjIAd5KgYUgSWti0QKaylB
g2HbfKV2kkb/hqmcSU0IlBleQfPctqTIkeMvqkJ1Lw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
N1fgHk2ZyI7SqVX1NLM7nNWID8iseA4Wyp/t1w/jDzaLq16DBPpY/gUfOs4x
h4CuWGoYSP2JJNL5VlZmD3rz6OVIprS+47GTWbrWVDMQhU6GRpZ2rUsqFYRv
UMUN81a3Hc4nHppPVdEZLaTu0+rZqLoCxn1SWg6jVtsDRAv7FWz/qvjh4Np9
pSHNlyM8fMKkW0pgtmEpOC9X5dNEjubE2DZNCasMd+DRJQdE/7vSQG+JEAeo
omZUk7W/B3v3OpX2T0Kwcpyz6R+0raPI+uly5MqIduICMSlpk2BX6sa09olB
Pu78uYWtBH5/U1CvnuPVsDcKm/sunmsiHSeHQ7lYEg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fBkOfYeJ3lnCi15mzCVCkCFkyy9jMKTdjE5ZHwKXxAD9gdJ+nHMj56lHFdcZ
V/1E1tRSYJwxdqWLgqJfnv3kqpEHZ3utQ0KdM3o93Eciin9uTuDnaMd5enEI
32uhZlgvsl3vPi0llSoXv5FqKiXqkklUsyVqhhzauGhzhPP82y/exYKXEJiQ
Pj4GALT8AOLOdTOjUCcIID64aeWLTYmILXjVm8Y2gkfcw60KmFFj2MKiGea7
u9eOe1IfATgENayYEQIbPwB16nPZxmJBhEcPMnWVkQHJpRRoV0MeS+Ejpo0V
JROexZRYFDiNxI4uKCImERCjAAgzFrearzVIlyNejQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RdYn+PIkGtxVGOHq0RO/y8VE52WMJmiLDrlqvm1ot40YP5mTmEuiEfMndTg0
WzdnZji7Vf6yMeEsK71H2mmFszLjSAfHHYRNBtWl3ZjWxrz4trLX2VuagW4w
fdJh9BS8hgDp0JHGSscU52Sf2UuyrD/k0Th7OG2G7Icc2f2tZg5M1fXPXPCF
7jL7QWbpoYxJPW0cV6dxOucQnxsAtY9AwdL002On/wvpGKVF/NqbZ7GDLtFv
UzYvW9m+JAMYePtbLwjAGXJmyI22cOib0F1YmV3Tg7ogelw1xr4Hto5zU/7p
cKwvVkSG7qfaV6vGMjJaueo7SCcLGY46rT2lnLpaOw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QvA4lCc5sWRW4c2VT0FTCrdG1fRHOoalRombPwwg4d5ohyNzAQu5QP9mLtgd
wYd7tO+WoR8bnyDczyOsHpNbMkpzIsMgF8kNNhV9Ud+yQMuMwUnod5jjhT/g
ipNWfyHLrR2MCUZbrJ49mla1hGxOQa1sBFxrTyuvo5mCPsUKRLI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
mh9aZNSBsf1wRXkpL/ZZEAX2Xbfk8tVLlTGCdms+Ld2WFHBmzFZtYFFL3SYN
/kylclfoNWVbJTLjYAxzcJpuwIqgdYtV3wqSooFxmMnkeRaD7p15yC6bgsnD
cS1Mqhq2Qk4GEul1tUQP6MH2kod8SAPSmkW2M78H8am7WULPgEaMujA6Fewv
NwIDf7asn4VAHdpJ43Y2Z911uZjFgbI5DyolvF60yoZOStO+1EwGTTxn7tvh
baqLkvMh7ho85mnv8KZTTsbQC9/rY/WINHkKcBN9lvdzJBb7O0rxMM4HNV2+
MDA8liyZxkTNSoUXof+PbSwdK8QYB0P7K8B03ZxAdod+bCFa2n5fzV6B64xd
YEJywcLUHIkYvP/T1CT9LJWzIaPGrzLA7VRrXkWr5Zgl7vohRXMkmKuiIFMC
Hth7iK7otyzf/Rf0HYqYVhZkLAAA7PISmrJdfT9gqY4wS1kr1wtIynwUe+WY
WzeogsvFEYyoFV8i7w1ipUU7/jlTTOvo


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
R/nl4A98D1gr8UnAwfArSFojGP0buf2RzCyQMrxF8jrBhppB81O29oeT1k47
Li1lv0HoKqpdcplKqbgvzGu+HY1vgt8YjuhYrvZqM0V2/tgWkJeJZagfQ99L
ILSLP+Hn7V/M9Jgt66vQnv6el07l4ARxQXNz18ooLHVBS+irPYc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
r44Qy6dkkRKi0HXEHuUsm1NxFNnM+JGWij0apCGPMHGVQWdCGwdddAl8auiv
UJK6Aq1H6cztq9zXt5QgKyiGpJkaoiKyGSjme7iy2KFIKlifV0QDn6Je/MGy
TXM9piru0DtkmB8486xHhzw4mHWpnqQ7SjeYediZDeBddpZCegU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4288)
`pragma protect data_block
Ly7VuxBbHF7Cgx3LgdNBhnmmU7CBqD1VC0PlSXWkrRedHKNy2YOHU3j3mfSA
16SBMYgn1CjAmIY5afk2IUNQiQH+siATuzOQ7kudUvBh+VgawbwQFeWaOVtd
o8W1JaNDRrOJT155oFhMZ9KYNG9pdyCo92/onS3WWmwIobrtAvj1URzVmbSY
5jnjNDWv0ps+lMR1hpZmCU+9S6HtMHiG9X/9RQb2oOnyGXIy3A0IE0/mX52O
7vxFvwZ6+3RtFoc7cXDzUMmQkXDlP64I/2ADHo+rHXrrEYn/dPz9FCP4iLLN
l3bjWM4ORPC1j5ZS75J3zeYM/AtDM1qXrU8wMBoCd6t2em22ESbYYUNjN9Io
uyhkT22bj99CxFHXD9kP31mny2ACv8tWrhgH6ObTq4pcSmp62XVKts1JLDPm
ptn/cVVIi8u7vWSe9XeYkrdaqWbebi2y2ZjNL0p4IdfPIPyz8BB1GpeBAWtn
WlevbraS5Q5tYDSm+SJV976g9oAQ9ZHIdpJYCBfHkBIkf/1MQbQwq5ettM2q
QKQF7qrxphKWLBmxKu0WD1yYlmeIMT+aMppP33wOIMdUR0wal22qr0cg4SF2
Lx13nzVTy4ss32DCbXkFEMi1GfomkwU1g1kVys12rbw2jTkf/+KucyVAfQ96
Vy7H2HjJ8S2CTa/Usde01QDp94UuoKhDStfHjEnQlZ3daklBRry9a1EVrMP+
OQSNL3Z61gNu1/bjCA0LKxcUhFzd5x4YIG6uCoA+0ba7vXobSsraY0Zl7fPr
S+wlr0Dhc0ANOstoID+6yo10X00tHaCDquIl3y27yHVe4sFa01YJHr2UyHFy
DN9VTRvtzf5EQWC1jcHVPay2SMwpt9Wftg5HYqNdqgBN3NltpUWFEBWlxvYm
vSJswaIKNbpbqBZAATxdcxIh/G8TOvXF7nR7LOiA5Ahv8ujskLJYb9qNar40
eQYF9fdCJ+mUDX9dajIkx+vVEH/xfLXve5oSw01btOUCWF75tD2kMCG9UGbn
58GM9yWpQVuGqOpSXIvRtHEjuhGK65y8GH2lrhGqQD7V3fO7YHNCQaR10aiG
ZRoipj54bM9Ga8HqPuQlwXGZuVWAIub1oa9+lyTRnREe9nDMg2z9ZDHvsKOk
Hx1OIRf4A7CjiZU7kFIXQzNYBFEtUD56HochqyjVeHD3EtTKIYyd4mYOhG1D
geghYHE8QQ5El/3BQC+K47wTyVcKF3gpbXtkbiGg2egrIU37vu+P47Kfz70t
CA/WNZ0funn00LyUeorrmmFMy0ALZR9mSyQhlWPsZzdFCImfRv8s66CRf6CD
GIgQIbEeTnBwdsdjZII1LHPiZO5yIJZX/WN715VpTomphWinl0HeOAKcuFHi
AktKsnBnsh1OpbaK7K5o0ObWsgOiI+FystH4OeOC1PALLqS3Y4bzCVIy8+pf
uJXP2iHlAAdXdN5Qs7t6UwhHW0E2PfXdwQpfqzDfuMNevfZ6cPuFooGYkO5G
oJtaCEfCJNWarwMGQtBk6QaiTg0VynJz4ydFFQdDCtP0N3uebqouG412/3vg
a7a5U6+nhUAbEH38QcxMJkfnRMkyf/cS4QQaYYGhE5R2uYta0QBDk0R0VDmD
uIrbfJAHIZ/KUkLBo9J5Mu0Wln3rIqLNHtewTHozbaAEtPAzI5lAtcPysKAc
SNHsT8AmE9zCFWuFpN0CaZ9F2V+ivtWOPyZWhFpjNE5QuWaZCVb7N2/aRAl4
56K5KbDctYaWiQhh96Rh6cs3sQoMGfxQ6W4sU9iz/YeVLZ7S5fTo4GrlAYLz
PenkXoc8g3NnA0E2nXFyAFF66hakJwcf7Q6e3zyhd04Md53hTh6IXYU+r7O4
fxryX0X4VFk77KvlKqJ8fKehCDitQpCHOluDucdDJfeq18jXc1g/+ideCrtY
5HcrVrmSfChVRDstQSl40lbZmxToLpBFNLllLsoQ7wbBCcRisOT+vhaS/gWU
KZyCJK7H7IpNQatkjM088xp4ZRbZwH18kitv1BheE66fGXAAPe2FdLnDSkXH
0PU58E/wRQzUfpXyVXiPkywmRPt8CbNiTO/+NWd3rIVfXGYTeXfUDbhSMSQL
uDsw/NxdPGRmv80RElJLjdzBCoce0FCu+Y4nEI7XHx9hEDaNcgnKVgFTQRbA
OQ7ojMJyFbDtjpy4uz3C0A1KASdEEblpUi2+HT5BzIlcbjr+J8p8UxVBWCgl
VWas8yyAsvY9FdCko0p93KhAS6raeSn4fYOeHSQ9xSEVr+JCC6q1V5rDQbqT
gSld7fQfInq3xl6wkeywBv+gS2Qli3o520g20a91S2IM5xHUuv2OUwCu+3Tr
2nG0PAd6b8P3zgN9ggd+tN96UzARetJA15juDl6e9qby91w71pNGM9vfYWLZ
vKFM9tN8bK/g2/UtCa3vhXT7cZr1Cesw488Yw0PrJjZnsTAI9EWoDwG39KsS
G3ruNQxij+HdwFS+Xr3I4efojIaPw81EHGUc5ejo4cqOLMscGYWUnUQr1TrY
yTQAr6SZw3mK4UeHwzExP+mAVklM9JkaSnk1TrDWKsUbS0y6ve8Fvh0wjpDY
uIHbHIEAo8G9uq1zwewwfhpltPjWfdx9ygjUHERJNkrBrNzg+QxWbXMoxwVd
gSIIfZxm43Vmu6ekaI53eALPTwmXdnGsnF0nhOozgWuWm/UoTwTiJE1LHkwq
/L1ljHZhNG4zvBlMPOvwJ2N69bRUw2iiEtwb3WJH119cutg1IaG2Z0xU6f3u
OZAldeI6cH27VwLiTfV9jPbunnhPHQVPi5ZevUNEoV8NxDwrfeF2S2sspLE1
HwTRGnz4NxSaElHJEYSufr1PEXDj/Ua+gKdsxwDHvUoO9U6ry5b3t5DiZCrG
vBPcN/lEHsEtfr2XVKlI5KLcAKiICT5w2LSpshaAw9dTmuUQAlGufNqwDPG/
PV68DvIZxLJay00BPaQMZSk3oNLXAjW8s+oRodskwJZeojOncnhU07KUUlDQ
RYYpNVNex8lRu0EbQZ4AsZrnn2F9P19vZ8S8aKUewKMc15QMD41tGryDRCfw
pDvHcgIrX558pGkKXX3xw+YWi2L2tEf6CZP8eBJUygw4c53Q2k3MUwxaLOum
5zkvsAQ4dUe5Z7c4GGnRvV2QN38LcShsE+PIYtmu6klSND7/FKisHqOymNJW
MtEY9B8Wf0cyaN2L5lyo0zFREORv4jWb9u3mIJ5IqkEX7uGhO3cBHEYic5Ww
KGLHq94DxDdn3idwaT7n9O4gZXu9pBZ2jDifPixJfutJ2LMfKb8PIPANa/L7
i8ss6OZWcWlhM4W0lJRswgE0HptwF9cmiQvZOnax+JO9UlRGE98UfxAKoTH+
XTT7veP6zKT4TrZe3wGZ3wilgofrMFiCsFyn+9zOird9KA2M6NDGpfJJ4QtL
fotmefG8B1kepXeMWpa5NmzbTEbtwhWkR1fTjiSII9QjfOa24PC12a6A7uXP
kL0dBTrC8j21dPYVjcpZ1QumyoOg64+1d7A4FCXBuiNibTfmIicy7E2qc9jp
rUQYaC0PjO+bkb1fERqB7sGiiHpQbgeXb29QCI7gz4nfRm08g22zFk8VAeO5
Gt8EpkEy6VtjquVduLxE9GZ0F/EBWDm6ho2pceFFbRBufETV1nG1WmxqwjVj
l+mOf5N4ZJE5himnYXjsXHdATmES++/iCjh+NApQQAZYzv4Uozx9KuSdcBQM
h1jgL9fc5P9UWVp2rGPWyoh6ZHlqVyv3nPNqu0mK/sTwDetjUx9+ryp1FTbt
h99pPZ28tMRzua9uXPd4BkC2DtaSqU9kOm6fT6W+CP/NEuIgdkwNIcdC8Uym
wRZhxZrFqYyUyaBv2W6/QX1YVTsjp7EqUVF8IMKxP7asZV2Xr90oo0tdUPdZ
2+OxbJ8uT1L8LIY3V7f1fLJzzF9nLR4zl6t17tH/Y7eb31bV32h1uWadRyG7
8Pkjy1NsWI7YnzzNh10fxnloehqrY8n6lVdx4JCRPEtErHWrkZVqXPHeRmkT
N0hYziPlCu0GoQWs0OvQG2DRlmL270GQ8LbU9hVcrI7SoRn4LLsaNOSfqEpD
0JKrDO2d09DOih4khkcbC1MrKknOIETAlDc5+dwqi6XrGLlPB49zvNmUp61g
IwRw9nfnVd9RzJcKcm8RurrPfw9E9yeP9DEsR1//t3kXM1n0bB4q78b7+05O
e+dG4nB0CzmjRxVwPAi7wTmyNpXhWBzm/3ephO5mDwtLXBfq7xLr0MxBrvdz
JL0otnEgnyYh7ryRXYhJJfTRtc9XNTpg6HOKOb0S4lzJvnEwovKZTzNDtHae
waqIqIcYAfeihellA22vxSXzhY21zx3qCbTuQm6vgHa3mhcKkvDzpNBbLitg
MkaQYuPtgkpEswWE5kelv1TsDDQek78pCy4fELVJ83lvOt2bAHxluMDgmHs2
06qwjQn3i0naGV4pWkSNwsJwJ0Iq149h18y3GxlcEzW6CF5ue7J5KsGjGnVb
i4/5QVaW300DHUzT86Nsk7Ueaj1rpQNWkiaKnth1A4LCSW0a0HG+PqZLF3ld
8lg4+HcgedKnBlFWiI1BPdl0Tmtm6GqPjCSUwFZMmmq51+xpS+Lah5NLzulQ
WVdrgvtHiiETGgDFgLIRtzc1kA6/Cit9J51jqLs7u/6c2Zw4bAlJKmRbp5CY
A60ga50CPGEXApcs7t2GikIQRdaVEJ2uBB+b2GvETbb1sZyatIKk8LNkM4FV
9kwmtlxkJbmO2Ai0CetSdTdCLFUCz+GW6d1fG+dpB43bnnHQUXM1ylh8dcVn
sp/1IKMJE09BECsfDoCH6evw5dl4gBM8ETkL7sAKhYdLnBoaiUdXgz7OrpTE
8gn+jetLlBzb7CAuDfZe3hDRIMqt3Ua5HSi1OXiKB1JtTJ30zvd+RXHBzxeJ
R8eSpSzM/GG3dFTd3tUbQ98nuJ4qOpVJszsARfrWnhOC2H/eqFEjNPZqy3/l
LlKiiaCu/uYtVHRa/YlVUbtYfZdiIHT/VE7gsa+gEjnOy412TD81tomcXObe
NWmhGWbQJnSeSsN3gaWEzwwgrXufSn8O9y6rTKrlbWjWjXRebuFxAcK9Qf50
opkw8+9FjeDQnVaxpfSQyxfW7XWRaTkDs8rvkqmUWcgqQRbzHcpdkGmnwl3s
s7oXVxDzi/mLvZQ5Nw1XBkZPrcc31OwDzk4tIdd6nAafV2czH5/KQud2uKC1
qNzF/dNX7qNaNPt7FjhoViPqx0Q+dmap+LcO5dYDTVLtc1IpiHhpKsqPg5cz
K5VIADBaycJrAqd7y7bNKOGWm2Wb+XuVSH0mbPrX0zKepJYzHyOHRSco2Ix+
YUjrUJ/z4AZIOdVkNf65Dp6M6cOoKraiIFA+p7YNVY7lF82SmchnXPs7K6bk
FcWOooMsIZP5b57WNqQ+63adx8+idRWksoTFKadqgniDGt3QRyIZj4/4GxwZ
Xq/PwIKnVkPJZPNuo3z67gFvE2j/GtJTUeh/4Zhl0YxOeXKU5+pMlQ2IP4P4
8KVaNDSr4gqhuMQAfKlrlz049/2joiBLNuDuODZpiuwxaZVv/5ZfHd44/GX5
OKq/zpQT2qgHJB3XXhsEG9Z738h6/gHcGMkcj8zGEEzpJ6Uh1yWTXajojTUi
xhkzcEAmGGdAjUo0ar53Z1kYhZFyGIk0cLt4dy6J//3O9UQ1Fn1K3RCkVoL7
YTHRw5J+jg7anVaGjQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpegYe8tUnS+AGTHQIzuXZua5PEz27OPA5K8gASlSQ9MDqdt9c1EhEH+3pEMqynZBbQtX+jkL+1+1hDBE9McDMkos3MfInpPNPDXg/qW1pnMa/17+lZxSf1H47uFwEUgfl40iOD4EOcejDmo9OPTO/zUqhqd3d5K2uxi+5+lxIPn0gsUYn8O9XRoFI+OB4zUS896K5bgw3/K9JBAcu2wyJGI22VkQm1uoUpHB715BEtpR5aVn6ETV4ia/Qr/opbz/Pzo3KjquJeps4qpijPpPTy/p2dK89Zb0C3qnaJBwAMaD+DGim7P+zO/reAbRgOghv9v7HrbWaV0iWAZ5HJxygANE04X0LENNIoR5AZKvT7XREsriTQibkN7yONVZtgrGohlBztpvpp7yesm2ezHU0mQ+ReSszSHxtOTlLUbjguQoa1bnRKFAk2/V0cmtQIgaXEBQf32RWeNrNFq0tf8Lrkeih1SyMrrfkMWzaxXoC6r594dOZGcL18JwvObVFAuf/MR62LQ+LVZDRRLLlGt0oJ9NIxgURrxcsrgQOMrtjUI+88WX1augqa5TQzMg0S1dsXHff4sjUOrL8liBcjLpN1/uSpZc0I/Z/b+UjfXlDzbU8zhRHXxH2D8KXaXzEB1TnKiVu2GewmgIBfgrB5tN0gHBA2MTPyoXELLySinT/AdDiPRL0p7vPSMx6MG/vdGZtKk8PUYWmMJF26Q/WEnnLmH0xoTBY6XlqhWe22RsK5NHBMSAoRnpkAX3nCMeW9dByPVqsGtu8HF3AO4YV76/E2k5"
`endif