// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
K7CV83iORS5SC9cfk89ItWqF1MvZ4QtkYjtHR2+oRudtT96nz+mSQfN2UFPh
itE81JlByAyPCqp1wgSH2ZuY4jq3WqtWusqbadFGzNBTK8i8T/ZhDDx7v9bA
qA2WWBDktLX6kZ83rJXVgIihn6Mc3Nw2p4C1x+icWJowlTgEhfrJfVVmCIPq
U+KY/fT5afHdbUQaZPEsrN81w6YXlH4v4L2UuRFulTZu25PJqd/zXIlA1Alz
kIscD0r7cT2R7hipkNeksbvo535oWAmaaGPXW8w4C5UlFlqtCvSTnYPkF9oD
qgpYodqvd6tiY5jqXcXj0KfDh+ImaJkVkcrhjmYnzQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DTkgtpyHjxwTNx2RbUPabSQxrhUhsb0xKU6DY90kwku730ShF6m2lK6UvU11
SBZuCWmIBMUN5gOveWN1sa1Y9vfrmC/Zezb2gLoO19tiy9qjw31NWGqSaFT7
6YMlqziqjR7qVa2mfMjX4TX7x7VZTX61Rf/aOlbdMOoyHBl2Lmv7dksPsfmp
7es3PQXJD8a1tmJW+Gytwba5aVB8TDpJOU/ODAD9ue24jYBzG4C/f0YvoP5r
8TAmU3Jeu78Z2MTGXeB5OlXMWN468d73R56RgbrzdhOvVHvfpKDnF6gLzN0o
E0SueA7lWsXUJkAVKPdgUmU4eisQ52LTBvd0XiFirw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fD80X5emicL6X9B3MrcibUqDlGiOTl2HvJNu5hgWlCgAI/jLL8JZmfKy1Xu5
7vuKtzTu0TqSBzaBsyEpgwE3yNVF0dd0GRbVpbALm7R19avohgr9G8QSKeTe
BxHs3vtzRquzMkcma5sIe5DgTl/6gJSk8Chqey4zxTDJsieWGpyqeEtqa9TV
fPoPdjJ1aQ9gwHU9rFGK0dGmx4nFaLGwkGNXUKWDLFbc5q9GzgjGnXv+s32n
jTu93srcN5vzQmtTGTcYPxoLq+G7zm4FFLA9LzU/h6jVseEZ6yqNF3TUvARp
ylBPHKp8GEEKM+0JpNIe2EcAmuqHCLcWKEwf2+CZkg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OWdDul0YfG96WLBbGGRh4jCboUnFsFKy3l4RDp1IB5IJsdSMCykex3wv+yfy
d8JR0kSzziLoF6pZGI984QC2LJ6XO+tOtNAvP+hxmHiG0/H1nXzv3JkJvJH8
TVLNrGVqm69ezmCmYsUnepOg0dvnl+rNCob0z91s4SlrzCJS8NzOG2ogWcux
vt/R35X8RcBknzwpZXU0/cjti+WJfx0OnItcDx76CuoF7FVwQhoZ3maEk8a5
KFqdVzQXOcsCw6d8EqyrTyADIi3iRHcXwKosCVh/si4VqKCKCEY6Vu007CDr
a/DlGk6eQ3bGqBmYy2ONzjJcbJlQbNUxHUf135RR1Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
f3NXA55vb5Mgw3AYGIUHZo3OC3LdO96kX8DF03fwLBCGAjGBp3O2AhrQoYo+
fs5TLRww1kw43RkVWCn9RW+FeIs4MX0lFf5fX2Rrg7jvO3v2mKYWevupbsH+
UluczmBl8PR6W0UgxSAd6Czkt/OC6CeZdJwMAxkBBXsgsGuZ7lA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
DBQENuZH8JAUE/i2eTCn0LWjmLB/kWUwYH9co/In9pfxkbYcq1vifGSy21xj
8mCnnk5jlGKEgNF7Rrg0u56FF9cdNZY4NAqXppx1QCzIxCVN9INSjax0ZyPL
LWQlRayC+G1FUGEa6OKd6HJTOaX0S4uBoWrcWgvLXVqszwrjsV5yV7he9328
kd5SuUDS2oZKXQ6kHXWJ/8NRToKcPVrSvFxpgdnbW7t0CRqdWXDpt0g0ucZT
PJsd61aJxs2iVdlG0/uU3cJInSG6HkAhbhiKR54RFjDEH1o3G1PD9r1yV8qx
YgDy9pkH+P1+SixFirwX9oAkpgZPYzsZxh2WoM+UCz9OZWukBK7+eqYsfcyU
kqYkOQ3qU7BzxOQaX25PkoCZoJfYxxBwhR8fIFjTuqF8l/WgDWhozYAlPiHv
CVMiK7Yk8DQ0dJG3j72sIYknr+x8ap1ar4cz0gsm2LIT/7wuna2vjwTcbnMG
41axKpoZsgD1Fhhx6HwH1LbX5fbeDV6I


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FjwxJ8oOTFOz35yu832ov+Lc5JkST+ruirXnla2ghtuXkbfThtl1QxsLE9/d
xV5bfB2DUY54xh5dYJuY6VQmtQUpagCxcJkazpVJnxgz2qgUsDvLTPCuSDwD
iY8QxnRksFj7K409lZtjIqbczSTZPbQw7LXdzTjJjlZjLTdXlIk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EO2S7V40On6zOuX6P/o3Xtq92SKq9E5sS15Y4UN/QutOj21nEq02XGENFnzI
q9blgrm9BuNPc1nAPpmHWZntd90BgXPl3ICcvFl9kgBn2CSCV8qICW3cNIhP
z077XHHPcXzV7WpD/9eLZFXDml8CytnJ4FX2wIU7ZwjeIvaMJp4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1120)
`pragma protect data_block
0RFMD7Krl1sVALi+yIem8/cuVs6Nmas3B6p0o1dC8bxic0D3vfV+KH23cSHM
k5URx+JhJ5OBuVpYncAJvQv2lzlsiwRkNVCTij1vIq0ZCPCens5RI9EPz1+h
TBDE3HgzpC0sXqEtYUuBHafQwPj8Oluo50aJZyecnBM2hiIO1+5GYjeg/fwB
Ys7W+DHKLvOWjFPEyAWconw1wbDFcr7ncnQ8infZbP7ijiVe/+tmvAoJr+8P
rYAixgRjqTflIJFn/2gNMhZIlHpyglmvcKik9BAWhGAsUapROgHuDTAflZje
qNPpKK4A3ouXY04LTyiZWWQndV/GS3TZy5CJJXGc9vKYCuvlPFP56xqko+Xf
P9+p9fIYnMJweHvFSFkwd2wAaBDAtydhdo7vaB661DkLJ22ezA/QJvqiLBOd
lRZ9+ZRVoftTtw5sHF1mEumcTQ9NqE6vUsG8YSkStcfy9+OeahjaQU/19n1u
VcjXkaORA0TcZJJHHx1sHcNc2wR8E75IKLbxVm+2ad2cCebaBKZU9NjJjVK7
tNImRhx4ePDg0vMeumNA84Lc1gcZCnBAscWEzvWBoNXiUSTzVWfZha2monw3
bNM92gSWQlgmi6VvktxsSPwOcQHBB+i2UrsuzFM9t4wj0ihIdopjInbWWlcf
KSmA96ibJUPo5+Wpyt8CNqNYsBZplDJCUhZCcUTacsx+mRVXfUSnu+Wpec5B
JDlnSYYs4q7o46MCejRBX3Nca1gQlYlkkMx1JNS3KKWNjix8+wdf9VNC5zFB
JqGSRfycVwXV2Cwe4rYFRQq68BUwPEqHm/BsF/96kGXrO0h3r+wzYYJCUd+d
nPwiS2pDQbmycPDXxwP+gUG9osIrFQngl8Log60S4i9Z/roez6uHHnsju5qg
qY6aXCx06mgN/9XzEsCps5NT5MfAKi2aawAGEzdblrG6rNgboO2ERbglqmOG
GoA/gVNRwmImn2+53VlxIuTJeZmBKnEhoHKDvpoRiipWXrKudmv51TBuSwUu
yRFU82yMoJNv97HS8pRCXZrde/wSkhnmvdiwgvIk7YZWggx3W5XMjgJmgila
e3oiqck08cdiuO45TI3yrYDc/RVytLO2p88fBHtCzUM9BmApIeXFd8pAs/uK
eRCXZ3VvVvPRipmcKli2MVyMAd4BCOJwoLjjV68nJoE9TgXwcC76NXYCIxtN
lln4bIXsCr5RSc6aFyoSr0ter5otJffNh7tPxJt3OcfaBwoyU5x1i+BxfFGx
juxy0qsCMtRnFvty+uyD7E2qJPIfeARjjmvNlogYsXzwq84Brq6Mc4Jr+QRK
aMvqwsE8BZL2JpZK9Adiu8OoLxI0FfzvLBtyD7nPYhd8YvMsB2rydDWc8+K6
0yldZlZmYXyJBzeXmaWtqpqdjXZUbP/j2aMngH+Aj927IUeLdyAdZrAOCllh
/11ixe51watbqkPKYIzBm38RLW1FVURrQufeCY3JQar7LCM9UUJ2mg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqeLEBk1IvQdtoXsOHmYL0A+WTSL24k/0R9A8oX5T36YcpgR3L+Z8vBPPXIEPTMac4nr5cv84WvOwmmutROCeAKq5L+1AxqCZDt9VSD+/Y4+KPD/OqMmRfOieVtdsbcM/uF3W+iGLidEazjNFqR8Zvv7W7OQYj3+oKf3z6W5IrkEgtP02JXd7sv2isz/3aXhpFYVzJvS1lYUT9em0pdoAWiP++KgzcaFTjx9EpQ2WBQ+DrXCSW+G9FjZlsCF+PHA8twlRK0YW2cqMgqLYIbQfEQmFTd/Rnz3+2lU1eFY3lLNW2QFj+yYWC48wLJqSO+io9hPX9gpoN306fdN1BT9MxrwFYCDcVMTa6Buqj6nfUw27R15Rp3gC1aMPZ3WXXchxVWlKng9Uz8VgHTxoOZdGgyISRH7kKghdqi2Qa6ps3lZLJDbmhtiARhuEa3jIhO0PctaRdpvuHXfkEkj0nCFU9KYyounEB0kCGCykUGJ+4s42dViQNu1/BcIo4Ve6ps1zhj1cJ82R0zGDOIbp2ZHKoM2hdMwJlJP8zJmunDw1hIVST8hjK7VX/81ejuxpPrHtDVqTl0Ax7ShI+wwvOVDuK5DMt2mxZqHBeAFinsbBCcNIKTc23+4AmTbZXD0kz+auM6lzIpQFGgAc1EFW/QFdKv0kmW3PPmFq/FymcBdufhkgbs8PBXpZ+k4aWxu1QNbq+CdQewqgTkTOqWua360v1Bdu/Qtlrs5cHQZop0GhL+cc8imwNn5xGieyCDPdxLePeWS3XS+6tYDI+tBEMcnlm4X"
`endif