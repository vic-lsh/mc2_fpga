// fifo_8b_256w_show_ahead.v

// Generated using ACDS version 24.1 115

`timescale 1 ps / 1 ps
module fifo_8b_256w_show_ahead (
		input  wire [7:0] data,  //  fifo_input.datain
		input  wire       wrreq, //            .wrreq
		input  wire       rdreq, //            .rdreq
		input  wire       clock, //            .clk
		input  wire       aclr,  //            .aclr
		output wire [7:0] q,     // fifo_output.dataout
		output wire [7:0] usedw, //            .usedw
		output wire       full,  //            .full
		output wire       empty  //            .empty
	);

	fifo_8b_256w_show_ahead_fifo_1927_mrd5iwy fifo_0 (
		.data  (data),  //   input,  width = 8,  fifo_input.datain
		.wrreq (wrreq), //   input,  width = 1,            .wrreq
		.rdreq (rdreq), //   input,  width = 1,            .rdreq
		.clock (clock), //   input,  width = 1,            .clk
		.aclr  (aclr),  //   input,  width = 1,            .aclr
		.q     (q),     //  output,  width = 8, fifo_output.dataout
		.usedw (usedw), //  output,  width = 8,            .usedw
		.full  (full),  //  output,  width = 1,            .full
		.empty (empty)  //  output,  width = 1,            .empty
	);

endmodule
