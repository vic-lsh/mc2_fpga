// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
uAlOtiQqkIttiEHbUNnSRTwfn/ZB/amrvxMhgocO2byxUsbfogQB7H5JxXo/
nOoptNSL1tTS9cLLcqRNW7/ecMk0mrL3nM4nsTfZLZOxnbXJnqiO2rQEvlFQ
xBZ2sOSaFdlCIDKqQq/OTl66TxnX8EmQhQv+eWyoxu0mXaWpm7PaoP5P+ug2
h/zIGX6+YWU4eOKsna8BtL1SKU/lV00MNFUTtKL72A1y0hq59AKPZZIchSBy
7S9xCHl958NmSigCFRaUSsrWa3If1NaXLHOsS6UjGgGEv1Np0xtZtz9Y9fY2
CLy/C45hCIaxorzjo/PWphCwXZ9Eex5PCEyEIgboyg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Brz3kMbK1FLS3nzt3TaWjdbvK+dB2GJqNkm4lcaDTXLPT+h4SbMfQTExb1Y6
1LIMzFymCzN9wQJ/E5qE+T1nF0pg56pwDJdgqYY9CKjLIBZs3GZHOhHLX2+P
QE/EstBTA9bbc9yimMDYsrcSciN3W4NU9vmoU+m0L6mFRMExdQOuXUTC52X8
j519erbnl/YjJ91EXKSb04uZpjcgRITl6LTyqPKGY7blwTuTulNmXStVOcMd
GFTY2hY86/wnqZGp2uwVJBE7o8/6Oia1DWV8WbrAl8TmI9pF4MfKbvVG2rNo
MndBzgnLLrossK3xXP/aJZuoCL0BIULV8CDUjc4cDg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bD39OQ2ac0dACSe+7QdmdKDWDz6vhRk2s+9VBTiw6I3WOHZBi5Eoel5/Sgge
3RvD8YAJGokWrzFbXQWpiZ0HFO0uN4JUI1vfeSTFETtGDxeTFVQ5T3GXXJua
thNeT0HmF5hvAQ+XitUIL+ERL3+PukupFwMKhHy1gwR28JnDSfyWTgedBiQs
QXbgS3HG8hBtbm1cHqli7lshX644OuxVnICdcXNeGj1fBw/QMv41GwwAITW1
fvOwviiJPN0N/FgaeAwPVyiwpcDMR7+eKgFDIe7Oxr2JAiyZM/x6+77qMSlX
CD66R9FtjMnqRI1nQXF79htRGE2wuCLMkhXTiHNjrg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oQSRopBV7i4b/JzMI88r5bHgP4x6R0K/3807vODAu1Dv19jBKtYsJBw7sI1T
VyGFvRZgeSd5WyjJOEoJ8QHMKdf0NFPoD/xMsesy+MeBdrfnq+GzDq96mR37
9GF6jNWVimf0wPNzp2XsAYU606O082ap5BmnCeQ2zmFRVpvb8FzpZQNU0d2L
7IcC6x6TR2YenK+t/XQEZbdusn3+v/UPgUNd5P1DsZVB5MEfe73jMOOvsJZS
DUvKSCkAk5KCatOZoUiIrNTtSzt++VxifZvFS82/kFuLgVz8UwYc3ZpCmLw2
8Ng1/X6zT5Pk7YJ1JLtjakc6p5OGs+xlOq1cTvgN0g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GbCJI3bhJ2d314iEdgGrc+LZT+W9Tg086SrRNI5k6RkifXktcYIsh6agAZHk
gzCS1rOFmg7zvlGcEIcR9k1yQ+HkvlZTVWQ+kaT8GgFWSNwzU6AjlShaBmE0
45YPwGZhXkMOKpvS59QSj4gy47BIuLKz8CfM3zrqk4+l3/lfJ1Q=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
pzKnIDkAhrf8blI6NGNtiiNdWPL4yB7eVDI0tMPHEjJb81HuFohT9XfkZ0Bv
hFLuyVLDooBRwDI2Oh3OsEQhFfbE/NkESkm6Je4xie2XKgFvHypA2jywV/ej
lRgdMOpfEvABWqZSpA3yFBTO9kWCebBeaNl1V3z+hPR/8NQ70QNuZnUP3JVH
2d1UYmwxNPiiAix1Kb7espHiAqJXks4vSOQ416n++csmHW71su+Vf2GHgbwi
LWFp7Ra5lXHMUhudwl0ak0pKPZZM67XiQpZUyKjxTbv+p/xbEnxQYJh53Qp3
SAQ6ldqNaXs092eZGoclKWndjnU7THdw8d1pnxDKdkIDN4iWRJFlS33sIBLj
r3Bop5/obf5AfGDK4eQnvFpUyK8+HdZEZ1LiVr+0NzqJCtWZYSwddfQBr2eJ
CG1OypOYgqM0S2nHGSWXrML8nb9Yc6kLvm5onxnnLqEAnmrkdXC32PwcVBvA
LOfSPghL1mASxkFGy/GlWh1IXLnNh2Xn


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eVt71zliUft/iS9eseURtSanm2Coo3pmot8hAQCt21Y1hv2JwLnaukFsljT2
Nc4E7ryQ1a9PzVzBGdsXuXiJViJl2n8QAfkcVAed0j5KIu6O6GbXUVZIGZFO
f6dJnRzsm0isw++pAtWHBQBxtDoE1kic6Fu0SImlUyLyPTmb7i0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ONHYjh7nXQCu71Vh8aufkeWV4YqMXskDLqe8lzc64cRAEQPKLiO2sFVyVIfj
yz6esCFXTuIpcLYJt3/iELvkTnyThR8EUSJy/zljDYvM+/jUw9Aq+GlJistd
3nW5ud4dlbh7QTgkyHghKnzrG8LkKb1hBxl22ft1hgZHwcfCsYE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10864)
`pragma protect data_block
BIcMSX0mZWJiA/C0Iv1tXomTNbPKFG52NoGtoSlFeQ9sbEw97L7Ios8cknSq
UmkdeQG1zjnHwlNopEO1lnvgcO/vFGmv5GYdE5biIMvR0w+RUstw/mvg0/ja
lfTpiiQb917MZ0CC6XpXvLQaaGNVz2X9HaWrb/2i8z2i+RuLv9ZvygNsDtSI
LiJ1Zby4Rln2e3Xx6UJF7cw+gAO2e1tii0+9hFe9+dzSxRPhc/ZaCakB/Rpd
wMtHvzMcpmwv01kwaKt1/+ssZK5ak5VjHsxh1rNUXXhyZvAm5fAEDfyhXqIs
hNv2PHBE4oAYc8mCvfLLPuhqFaMibvd7fH9DzgTUYa6qgPjVAHdgQhTR5sBs
nCO49EVCF+7VLmb+CuXYV9PoFpLWfPqFIfRrplQh+bW0Sc+y117QolChWCBa
U77BTzZU84/Z6yErVCmRUVjp/gjUKXF8BJxLrna9botiUPeAWR3ftdl8SfGd
TI6Nmh+39mBzI8CLVF8nWgvi1vjKuS5zlSPkf3CwK+pkYuwevqHJ5iloA15M
lz1SHJG5T3NRxP16B9kiDTVxjEQfKBGq5d75iVlgnIWcokpiCd1zjU1Fv4K2
YlPTZSswEA4/MWzqawrGIsh9+YOiAIvXlLwKZWKwA/zo+tLpKkAviwodjx9Z
o72o05ONBIYpqrf8Yql55McTf2GMrAkDPSXrIbATPeV0xSXgsHdOdy36QTNt
1gLXG9cP+G+EQx7YwpbNxXwOK1xd9pFzF/p7fwmADv8AoGzGbRTypNARYZ6d
HjZZOGBIvfvnKlELVTHgQlxMTjDAE7YkXoNfZ3C1j4xlUs5By6JqfDvcN9Cr
N3I/tnP8AX4pg8FWH5/xbzCfEhxMIjZOemJAWs/P8D/b7Th5m2I+uN/wIjIu
KnE/t6K5dGHdrpX7I1dWbl/7BxWSi0U/NAeXDlmDecGUfo3QiL6eAfgphXeW
talvgf7FxVkiMyVgNNjomYWNhOIHanOM+qBkjHs16Qi7T8vfocUvn7x5ll+c
bblmAqjtfWa/nSpeBgX6/CpnpK8qN8UWPuitpR2v7h8RyXJNm7CruGUlvlLo
Lp93IwZyvvVt8AKbr0bfCafRyoD1sSaksiLIUvr30vMdsC4jyYDPlOErRiNB
Ucq64bN8HV3+LiWpOU2hv+hZAfyvTq2qhpzmtFuMJByu+7IytPI+Ri3P9+OJ
X2+NJXPxKHcKOVbaTS5x3AhuroOQdmLSF6gydvEbkGVOYPmEgCel8BbgbHsm
4BQQtl9Pazon7GvrbnhLVjU+Nf6MNKbqYgOFwKG9H4O30QFgjWB+SDsawWt4
BD3buBhYYEJhC8zY1xQu6cT6PNED7874/VC/oA0cMvJZE79PgTz6+I37R3Ya
E6rFmjJQb4YLZAB7hgZZrZuWs6o7fSR1vD6Y4NCqLUHjWiAc+WqD4GlpQ8dv
07UIF2T7vwu7xV/Jk7M9HvgrZGAn2xNZxXIajJ94heq/opmMP1NIojnGC6V1
7MMSnRGBQsIMpBhlr0nKb7btgMf8LM7V6O7n8O8ibjxLV6kvyLqZK8vppKkp
Ts0Bc7GX3JmEqzUZH2xShE0bIpWrafRL36COH/iZrOow6DetMJJ9+Z/g+E1C
PQTH8JSChlzr+yRWjcPOsasX0XinBSMC4I54C0Qq7PoTcOw/A5CSciDJfuni
LH6hIy3ToHEvo5ydAGEn5RGxAH5dFScddn4dBHPognLDqGnhCnxq/GXBX51L
mch/vVNhMotXYOvpBAvC8lsmpsdmNNTSr51ExUoxze7Jm3RoO2KLlL0nA74D
DTwkLwbEhCq+XIu3eqyMb4QKCBgYdx+RMs77vrHS3vevdpM6LO/oeeTjkoGY
LIiOGxaxrPyIrF2wHZk7n2lafzGe2A0Rc1anO2bk0+6Lp6rk1mGjCMTiKZfg
hFQp9mSny2+rXILvXptqzljKbuUoK4spqz/P+/uDlZAOsBS8ufbeQ/AYDEcn
uSUHxLNhq3GVd3HLmCL3DOgEGcEA11xCrL8zL4o4tdSbNJs3Izm64p2li0Yj
8I5fqxr2TGYg/3zmiiG17xPd62Uk2Ha+YYA2n2cty56yjlUHd/ViAAH73woO
zBPTsMSiaGiFdYToSqeSiLDT8V0/aeA+ptDrc5u9KrYsyKR5Ve88fVopgYVf
HMPAnmcRgMNMeiSESrVhWwEYSjlKlHiDeHBtWCR7B5dbOIiuJpUAl93HoDKN
VhwhQSg0KTFePDswLptk/iR97qH9msl/kDodQnaOhFmGNgiwI2Pwk57XAm9e
zCAL4Zrm8DB2e76QwW1br5sOIF7AP+JP6MC+FQHelJA9nszfFwBqY/CgdxJM
lihKisiYZShpZcBlkIwwUOCweAhPMIETmKQ1lAoepBcaDntc4hfUK4AAA4iH
89/gPjnthAcbHkk0CTg7mrCbmvhM+tQYjRYCbHY2B3POJIoA+9DfC0bft2bG
CFDcYDOWAmMc+KnMRt3ZMoHyH1yJxbW+kqEgm/w18I8prIsAHpY5YkTnwqjp
/i1EwrnoCIAtVCMOoVzjLtztwX0E0ken1Gmm/zI6w6hdDZhVwqMIK31RNvy+
NuN2SYtnrzOw5nNUK9Zxu6RP2xttpBQL8Pct1gwtDNHtpZiv7b496MhCutdm
9iTxkLniK4Zka3T7TIJY0opDcxYqX5V1nR1GIInGZ/1Vo7EtxScG2Fb6fuAE
zw+nIqBJQLx/S+OxQo+E+ka3chf9x5yo1beriVf43VSxa45yj5Dbjh8qfkLe
tpvsWwQ+p/KhYP6snZTLZQck33cQ1BvJTx3riaXeKANnMlRFtkOMN16OWL/F
gYF6oCSMbMsIUR9aWC4kRVgEgXlJW366EGFdygBgL4j6tDRx+pZwFpTi1hX0
1BD4IYJXcrwmhZV7mRb4WrnyRtJ5rzmXcoeXODgHzJoKTTjruMtTetd4HTdm
wawKiWolojMeK6BR2YGO9CqbNKRzII9GhdrePUIzHh9oYmPmL/HKjlZ2PSCZ
vG6fuEfvCqpv/Oj2AOaVGIpzGhQmKoMqA807tbL6kel73CXchTQKpc8JcomU
9hxQI3PoUcSsQQX0xx3iYWBYjYDKcnwH9DmGDM+JEa/zRYjw5M2OBonMa18b
tNiF5Xs0h+jG5OMN80NUS0qkUpvVZ7OAW7/qFSzMTAxSsnsuE6g0vGbEOrzl
4eEVYtSgCWAsvWJBhXwHeaE2ocax+ID+Z6vgSjV1/YKM8zsQVAwtCHgHssqy
v5m81le5l8nS3j6E9anSuwiJDvHz940q9QpzaXI5+1i6RcXDa/cHl6yylNXB
uqIh4X4isx3dMdRbmhmI9nLoyAd25dU42lcSon95PWmt55V6qFKdf4OQOUtH
bO0rju8yIq+ErUm4I5D7NYU3Tixca7FctbartwQWfrANJZCYK6xVhUYRkaSH
t/AAWC+CKQFoDtSUldL2Z7TnYI3MpXgCuxZCTwb1o/ntZbUH+f+A7YKASgFp
PGkkVjbqCaDrKgVgvYh58s9SZRMHf3eJWCOKEEASM9Uet3/JJr/0Dd2qUx9c
eCy/U6WRZhSjsOTfWee/E5MxoczZ0W0m4BGEDu295zi8ow643ifro1cVDWJ7
moptPGspzuNawwAN73TxsuAgjhOxXlDzS5/kGCFLP8E+SokkvKu+gF+91Kvl
klla2NU61QL6IltlF+cUF4BcFEc9YZx4HAHi8vVq/3ILk6ZJFHj/q67pTX3K
R5CM8o3j621lWtvqvGatrfII5CkVZd+URiEaItgh/OerFB9vrl6Gc++HgDse
91TVj15p9o3MsKwewuL3ZGzMjwDFW1pQvgsV/gbT32cQPRMa8fYsekHfsa2w
oHgI3q218qUiSxxpiP6BC+jiCFAPLbFYs5xXx4ZCZBGc4e5z2wPTAHK5m2qj
Ka0PossY+l5JNHc92uhfgY2oa6REK9WHB5l9IKED0jLsS9LXyex5TpBkOMsG
W+hAUTGGnKzZlOm4XHEro2BniK2PjhA5NQhYkCzh042Q/1XQjg3258PFzNgP
dQIb2nGbskHU5FUIY20O1lDQ7fuXFbxxwsuk5pPdCsjRrqU0V6rQ35lahBuy
eV7t31oeFZSymI1nING9GNBVmHNQWLa/FWmppx4EMopeiOFhUT2yVeSgauPp
r4dtTJqkeOogucygMQ7nZG9iAWH7VkkNKGqsQCjyP2eaf7d1VV00b5Lmmuqg
RfPTGCIZF4yyY2DcCilHqIFiUJLnreDy6L6QdjIcP6NU4MUeD4shA5p6UyuK
UHexcyoFdmyq9mfHUPfq7p547VD4fSbHXuqYEx+nR3EbOWMPpNOyK9fUr+nN
PJ9veVmhi/0hE6x4I32v+j9zJq+c6Lv7ewYETJid83+XDA8mW0vJV/3+uDb3
XLm3H/6HHDcBDcsS8dHphU62qSU8ZlViS2XGQTpld7LmYUIrYDhNbJvDHEWN
fuzxX95wRfzwzX+6RlZ1XZ9O8vpgwLAmivXAacW0aF77BcjaU5ZuKkmThgGa
kuklTNcGbPZQX8xpi5nkEn8MxzT6/MDn/DVInab0PZRgK/tRAAq6kc67WFf7
UKsjiFh/4UiFaebcjRyrNJpFLOCB5o3DEBWg0xNThxiKE3udcTa2f6J3j1ml
4ocW23EGjDuAZcqAR8pGELLh43r7ZCN5IxoNY/nklYUNDrg7J7+5Grw9rzSe
HTH4L8gxVwIQ5zcSsfJoFOj+bnkGoGe7Ee2BtqMHwsr68PMYYqQWMNxUrKEj
UBpGvFS5OcyUvmh71/qe+/Grc2n6FaopyRgVYqTPGxv2Y+sGZKZ2vFpLs1LA
38aOcntSI1N/bb9WL4tv3ygus1soc0O5H3vBDUa1DjM3s7r5jxq9cuy18WJ9
boBd4pdt5RmLP61H6ygJdxTN9y+XJyTM7vxuj/941VrfAkR2m2OWmNcAIe7D
lytYasNnoTk5ZVbd2SHCAbIYqaWZT4dZKgUvnO0pLNirLYqv2tJY6A0TLohj
uJBztKIvlbxy2QgvHgh6VeO8WrEmJNKiWg+axJ7/6s45UWH0t02WsMBfLhXT
0cVdPgjggo7aeNRrRbAev8ajNXYmm6Bkq2z55ln3l5zIkiSJAyuqLyCbClbK
1zF0fD+jN75BKC3KlIXuZmB515zddrqJLhWsN51tdNYywrgOP8qlSKYlOF6a
QBzM51s9BVBXgBhnE8W+hHk3k7t1KW4M6FLGvQA1YpKw41YH4oEFDYXfHTRM
wjjWc/neo0/g3GNqkuE+/cCf2m5jR8kJ5/96Q60nqDKCLmyNowGARYQuFOtM
I+WWL81/GqtxjWTQHXvfjPx3BDskyZshxSBSIf/tvMwkjVeuwZhYjC9FcQBO
bae7a9nK6hr2KL+UfqCzvOY9wNIfZWwAp26C0ND90PB5xKrhHjaxvFYAqfRU
Rjc4FPbKdRnfjgvWbxG5OLXV0lOm8KWIG3t/h7+72NL583+uUx2DmmBTsRfC
jN/CpeTVHaN+7LJJpZmkMb/ZqUl/nQZ+w018ucnv1zgcCbMvS8tZ8/dRCUHe
nqdPWxj0SiP5lLO2c1V5MATGMr3qDhgVXB7wM8E1ooqvLPE4QJfE4evqqZc3
MH7+7UNm2/cTZbFFTZmHaVf86LzwZyDLWtLvRxBFl+f9H0dIPEaT5T1rJ/AQ
ib2z29Pc3oeVebBUjmIWBRsoCwTV+KySyhIOgp1L1HR1Lm8dzIyzRxi6Mdky
Hnjl0nAqo9+kFIR76w/x1ksHPvDQHG1FuB2cQLrPiRTmngigINAcMpIRRYMH
n93sb8TAjzXU4VP0oygb46A0S9lj2J3IgHcGVhoLisnnyd4wZHWN0/jMmVyV
xUd/NHv4yUhzQHuLDqK/Asn+HHCDGONLJiE/G6N9UXqsZareohNMMVS6K8WQ
DrTFVODuFubSrVlul3V7ZRosRvV7k/Tm5opY3dR7BFZR5QFOBIv9XK0EjcCq
1PkVN0BF/xu4xn/lirdJgAejDQ1IjdoSvMqULoWE6St3XRSFF7MZkwbc6Yxf
zmKlPTDNA4FlWzFISyx7iFoY2Rk4W+bG/RFepv98LMOnTHeYf8FLlzmrLZqz
f/dRuCf721yHhVIBQO1n1afncUKcLL0sV3m1JaVje2BvRRWF/aQZOFGu3B45
siv5kdRbW3kVKDn6rUIr/K3lGH2/YdXf3wIbhjY+nUfhwrYf8m/jChn4tnIz
xSxDhfBo4/CtkPZUsvwDuKKHHK+FdITjUcfAGqpNXg4c/jogU8IWNQK5rRs0
YhOmO1+mqK6xppK8DBe/pPRIfUdHpCfb3JNAr3RzYLffsOGFIctbWlFSqfno
/3RN7xK5SIcRTc4jNHBUYkW0TNKSufinJrzH8H5AsZms1iU3ZJpz6o1cW27n
vu4sALpRDmRYxoJzjyOkStKUED9rBTohrybKKYYGX8XAw75ZBxx3lzDOxH9T
JLavOabYENpfWC8Pn+J+GF4/Y3HF2Elfxs19ahVk4ZimV/sAWH9kX4ctik3B
4N3aeOYPWXEFN8cr0WoRXybY4NV6PHYUi2jyhhLMLUyMpWp68wQKUhLvq1UX
KzZvRReyrxJ1+UK3s/rn5JH47GawaSNh4zYXpdyd2rwHkx5WTEZJ9udwoudu
QpQwjyd5q1d7+r+Pslh+DiSz5ZJIHfvrfNnjOsrEo+z0EOBzNBGRjVZbRLO5
J17BlIHkIvIClv7RpNJWR+fv2s85B/zpBSUzPQ3wJH1NA2hiE7NKcLhC3Daq
LBJGJe7BTOvNny4AfiARu/ZdcevrsLNyYAtxTp8vyNDLhReoSaJ5lE7VzCUk
I2JrD+DBE/j7BTSdsmhZHb8vQzl+2RJWOn31QIDkA4s+gkUO8uXSdPurZtbp
lqgYpfUOGNhpEtHY7PR/7OUb4/OQjH0ptsI5qlDVTgqN2umw/IUl8Vx/JnqF
lnd6vMRG1oLY1MM/Zz/XOeSx4JXzikx9Q2ugps0zmJOS/CFl9fX4x3IMabBD
fUEyjCFmo/fu1PIC1/oO+LZAvqpGFZJ1a9zovB3qSwbgI0HLWCNjai+kW6Gd
ZHqIn75rOqHmYshWmuyD9v7trv/Sj1qqWZZa5nDKe9wtPhWfQmsel81gBsmt
GbVIxgd1NY5lV2RBy3FZlIhdvLm9UwfVrcaOblkHhqKbRUBIOmmwZpEcvFvl
SLvJIf3FWo1Hu20GpXsFGSdZqLI5UVL9PXSHYwray7SA+Hgsxs6LvhItdYiV
sfvC0PhrQtzaIipOxAigDMdxxEULTawyP+dZ0QZ633Sx3M2UkBNOBa3qrdrp
CPcwxQHQXehLo3UwwQpvQ6qsOruu8FZx9B8tf1ofXwOCMjO8iFB/WP6C3Dai
aR5/0jH4Q0eGj7UNVm7VDH6b8tI1NfoBUfoCEiXhW4vnnghvtfZBBrFZs0QT
eCtX2e9o123Rc0dKs4V2oaVpjzoSevC1e7ngDzLVbewmSMyGrbKquAtIdFiT
orsKuJorXB1X9lBOTs/JiClE6JoSeh/+nPbQcqS3QFPWQTE0YjAtc2YRxO7K
ZbadQ7eRlwThiw5oXoSjxpNYJow+pT8y9kMmlS8a8TlcG95Yfx02pCuIyfIp
1Y/BsxqXjxNfswjQ8B2Ud17hAa+tTSXOz1i5RBdkeCUi1cslcBdBuXpIgGhr
8b9zc2zr/qRq7knDS/xQB7OiXoBwZdNKkOKBwHR/hfw1YsAgc0N1bnabIsQb
y6CSt6bmwG4KDI5pfrxU3uQ1mkuC6ndOXmEhb3wIZSDUJbT3KjsIwct5ZtFB
GZxmyz4X96sQLf/i0TSH7KUXXktpeb0URHP1acEI5X3P6ExR1+8h+RsbMGak
Vynv2uCIAf9M5J9wXB0H2oSWwBbQU6WmHAb3MgMUcjLoCyXnEYbxfF+VA4IO
llmbkNVJm6uwiwIn7l96vHs0LBUjdaH9xjBVzC1x8L8T6ARPS330yPyh7rHn
kWPc9hGkfk0l/9mYC0ggwpUA64CLDHHHX+evaX+239ljFJ1JRzUn36+u+nBT
51TIO/vkRkj7seUP3RO97KYgIxNClrmP5tzFJPchcaLiyQtGKoyyKeH6i25S
8NjVZ//RgQSu3kWC2CTIvKMBtk20zq6e6QY9En16sPJcLUfy/ILREw4kFClC
rKeQDI0OOdgWmnbiXWbspjz46H3EuNE2xAoa23NN3v8v2PS5y7mUhzl9v5Se
vKDmKjgoQnhAUIHTTcVCbQw3evH4kfFjdTFkjhkIJSnSSKXa/d1iPkJr6Y+o
P0UATMWLOFjAS4OluD89MN+/z5GEXBg+mK9bSN/YiNanapOPRb9GEcMyzHOf
0OIiIC/Jy4rX67P3A4kvr2XetRf/ZZEMfJIpbEyrg4dlB5GNEcDNW95uM2LT
YDn2JM+thGhTuKDUH/6jFlBIDRrCj1M4tO1G4BpKjhmzGWd/zVd7eeCZBQRR
wAdFvaiD4Gd8CQesOqDtMZ+0RkEbmEkz34ccs2RkwBWcP52cSD+kwAitwFNH
/e46qaMeHBqchbYUB7eRUgyFCwIf98iRN3FTR8bg0uxHms7/QtQwFI7vSxBE
SIjr+StW/TpQ/LJuj//+UT9CF0P5Tf8YbT+gqy5h82foToiTYAGuDrsq1QQV
3dVlg2rkKDQUa3RRmibzMeqGXMVP8RoxchhOtBUD+4NRmVzILpEXe7T2gneF
E0DsN0XLiFNWISwHLlyMpkWMoPPx2VAbMTyekt1b1HWvHGDQwx3WeMM+KG/R
t7Xqrqzjtng7y1BamXcU7yM4xFvrixeFaHqCMH49K8h/BTqz8etNHhMQruhE
k+YMkzKYAWtQp/pm7R4o35DEsf/JRwkgsYnbKpniObnFGStBnxkcaXTvarzg
svYiqaFvK8mhIDr10btcYBSQLRWCw6S9WNs4UHGs4sEAe73F8dMi+dLOsSuv
3/ItNbqmrPqCMOAEMFJhXYBkpaLaHMmdlNKWITub+vkpl9eGmv++GBUwPgIx
aUnyiCVXSIRVa4/TGMsDke64JxND/Klm0qsLD+PQgNnXQcklyNRm6K0k/Pkm
GQ3M6VbxArTaERdw/TtnHAqAJKMju0DAyGWBtf2Yg4gDWDQ1t3rkmMhDOcQJ
WA5g9YYMscdKzlhuY2H6975smslC5NYFiBgu9GtJ0vm1Kst6OKAURIj2TqDE
zW/ywjSy68Rz7IC93YycGi5ZK+POJ0pbx5Z+llnmnF7dveLUCFRIuMux28so
BeFPstKcZSwU264wrJ+Tw2BqmmJXanK+zgNA+rOe332zMwYAmPk8eMJF/4Z/
BintbTPDPRmZXU/fSeQIoHsI3t1CLrgDrHS/VCkxbdT6XJ7KLna3aKZ0zj1j
H/siG448KRAanx4hg19ZRYfEHt/8e7B+3Kd/1pkC5x1JN+9eazK31SOrSa5y
q4Gsd87InoR17mIxuY8to5/Jq/vGlxLjntwQzl7PeoTDd5GD1FNaWA8rGhGr
I4Cghr5I8pbYl405UrjGCUelqnu6NrFjwYW2FZMDBDEI6mdSKZEVSqNh2lqU
PHA6lnVQblWFbwjAMS+x3wWgkQYUgpuWng0DUFUKyfOC0Zpv7DZRNPa7Xv+x
bfwLgYJ+CyvPkCAppgXpXeXeza4544d/pPKvP3kN4AdZ2qxWyiEhb/9fI3Nz
vYIlewjZckTaIBCuKBB4TAT7Nt9jYO11izYNY6J2D1uLt5L4LEIIm+COJhfI
07cbqsCXpmGF9PPt0RSV4fsSUpXjm+4ovijMA+s8OMmxspp7R47UmI77dZrd
w6NOBMYdMrScbnYG4jpwtM70UIDNHEE9+7bvfF+gymWfqFGlbSnHwXAMCMRw
AzBEHNxbTj5KvG7SmHHvk5JiHqB8pM0s6EcafO+G1TWCdNu90uYooL/A43bN
V5VYho7AvxHK5oswNnAv8iHL03Vf9/Z1ggKzIiT3hup6uijwNkim5GPyagWa
Uf3JUtFShGNCR+zRi0Wn/9prCQcIEVTdW0Ed0wbQRHRfB154QbRj6W033yUQ
ht13QpA5FtfRFCMeeCXsVXwzfNVEJYfGvslDtM433Q6kH6ICVXBmip2bjAyk
N27opxfSxU48rPEGpXqfUxVOJwsyqDP0rs9iC5CKWOhLv34mf1Uss/Jr9LWU
YomPdlFXss8QwT3Cree4N6O/n+eNZPi6BXMkdFsgpT000aJAI/grP9wv3keY
6JW4fQcmAyFBweqke9W4O6TtDQ4AJNyk/gtMpSC+JonbmewXx8HBe+B6Ytnf
jf+neU0yE6HL83wCZ7vAqzrnjImhlKdaebN6D5wGIyv97sohSZeQ/9j5dYjs
T5sHBKfGgEI3iKOv2B3siF+1uPtfXuGSUYNHKVJ3eDArreZPlHzt59oRAJMq
29SThJDR3KDNGqSptff+uR0cr3OxsXHSmpoIuzAPBilK+Wq1ra/Z89Rq4kcx
FaH1eiUoI1lnaz2kvBSCMW1HCUgtY4Bahcnqf50Qv3ygafBnpTtZ0eJQN2LB
taDSQczGTy0uPippgybC6JK02xstbjiiCHmYWLhuN4EB6XYGIjmh12+Fjs9s
WBivP4SmDkksA3augZsCu/Ppt5BkdfGEZPH4uINVqGz5G8/ziyZL8N+oHcCK
2tyI3bQ4PAdkZzopCvPqmY8xpCB3NTpWf2UIflbOsmlgPnULNGHC2fKwvPux
6J2qyoORi0alW9x1Mi18KR1WeO3ltmVkyoHCSIznKqf6bZISw4XoXT7rSxF9
t2SV9cpbeC1oZICo3x/6etPQUAKiTYCE3B3lwq8BtCt9iO2H8BVKdIduJHY6
HPV9GlxpJDIoY5WaAOTq5Z7SYisa5wovlCR9/S6ibR+n2507CfCBUjOoeivh
fXqr41RtE2fv3yH0v2EO/OnIM0RgDdO7Rz0GArfV9WKkz1rJa3vYdDPke6kG
gShbf0zD5bD0NWS6PNVj5bR+bbUpi9M74Y9Fclt5trvmA20Km9Hx2VYIouyV
BGCYOOkWobJHR12iqPwlmy5l3ezpGkvCiKHOXG9b9mEg37/Sd9YV65Bfwv2Z
Ulylnvr6O7cX3ctSiIy8poJ/c62miJh4bBuxSAkbYHHkSVuvkVkl3N6bfj2s
RCzRaYTq4YHle2GSo2O8FQk/yYjBp8YBLRKKIgWDoKMnH63CRE+9qe+G86oU
tyPBOU3ul0Y/u81at9KjK4KcDH4pM+lh2nN488pyLCR5ZU0BBseQ3MDRId20
MSkfVWYzIft3ppE3r5Nuu+L62JPwDxYdOnIUKoaj5Q1pBeLFTZkK1Yr6Of5N
tkEPTxR7nB5Q8BgqNuriaxVkv3fxhvuGx430fte5MdHGOMwjCvqyF5G4cZBf
VdphNyDvOW5gjNPl2v4sS+L9JQ068xwyAYSFJtNmZulm33msC3osEW9Mazf3
NNJvanoHtPXt26bDHM2YwE7iSSTWzA312oDTOOcsLgDPpOtPQZS4fPPXfaG4
KaOtWCkSLung8rfHfiZMu4JI6EpdbAFcFjC3biKAIxhYF98GOLiCWZ54VYWw
kLrn5lfdteNs5xBmuzn2WKaqcq3SQQ3p7EhpEUiD1bQn/GMPSEDuCDev2/uG
vyt0xCJaWNUQs/zHg2KMsiKzt1F2VzuzQisSc5DXOXPlmGrMR6DRPg95v9mf
ep/AmrQX+D18SXx5GwgJ4rv6+9pI/W8Jlu+M49CK4GCNSjZOeTJuSzY0OUyy
oofzBfi743mkJP7kK9JdPIpZx4/njwy9YcQpWzKr4XSGVSzdOUxS44+Uvvq1
Yg1kWPz1V2APJhxdxdqZWTscpKHwGqRCcG/4zFYZiu229GFL7uehrNxpcdHF
1Lbku7hXjam3vw8pNImXhUKNK9/bKd/66q8ux8WW2IX5ibIzfUmKwqXv3Meg
SsdMCS/7u2mj+oPch35oOD06n6FeBLLsI3Uzy0rPZI4ohiMWkDecEqzGVysz
2l8hY0Bn9I2cT9WaBgimVciSn7Vq+U5/KtNPHt3HTZmPWKHp7oHqdSvSfcaH
XEoJ3v1LxCybJVSIZeMifuQIHaxlBhoBPyOSomMjTVTv3wZrJEOFYJIYmVN/
rq08lMKjw+5N0FnleA1Ef5L7muz4W+5jM98hE3v4/A8Er2hZFm0xcxiK2lus
kMchG/JIPHNIrcolp2sRUZGnUvg0qq+6iz31TRgnWa1wh7GsQveB2r/UwfYf
hAJUTtk8XH+HA2u2Odu7HHJGHQuvp+kAbORVLr79Kky0ywGOHFPHSG2YOPpC
1lXIDG8Ze4qXB5v4CVWQLIioGlhM7HWrMAjfhi+KUovThkQtXj7fpYghoXQC
1odtUYCTp9JNgUwF5H4WHeHHsaFgK3RpFOEwtJf3LV3OojOJJyze0AiA/vPV
18uI5trEEDYoZoaIlzW5HlyuF60cOK9yG6SLdbHGGJSZvDkzlm2diuZaTHCY
QOPLrGus19S0GlYvsem0oyRfPVgKwLOx6ZP9OPsRTElURf7c3dJ3pnegwuK5
HTu+1NO1mv4t/Oo7zeMnzqbunfF5edJzZLiUT0zitr/gsvBGYFxZDyVkb1OW
daU7J4RZxWqwHOtZuMr6LsZ/GQqQsnPGssuRU3JC364eOIL4MDRk64hTDxNu
NOFBv9+mEa3tFLXVzNb2W7mtAnGovuiKeFU5pysAy7diSQd2UTpP64H2+yu1
pxMCLWiar7YwMb0QXZNOfrSf78NWL3I1xktwTE/zxZJighjeULa//cB/6NNW
agQVHXQSfSqMlHGPsYSqCcgyX019S6QL73OV8eRY2idJajccu596Ow3ss9A+
q9ubgqrY9TAAIvLQ0n75Ucc3pcNhHL/BbtbCX0LyEh1e+oWbCs/woUh4Qx01
3ok0o2NF1lMi36p9rFHanB3utBJ0InOFMAIuXoTk1DbQshuSWARyhkKxjS4m
5Uh/uxwLQTZfmKHBJBWxGu8oSVcytQO1g3Xvufw3KYUl5mWu584vBFgI6AH3
LBklQghVtRGTFB2WDduD+jiM2exTwbpda6UHfuWdw9gyztomUav2Rfcvoami
O0E+DbBsABDhDfz3sM8CY08guTKjt8p3te952AKM1ZCNgtTeNDQ7BnUZ7yhk
q+wPCOnzAFTd20VhVDjieA0WdKe5hbaTi9Cykt3YiPklngYW2KqQJYylugHA
xi27GaKGeuDh3JlqRwSfT8eErji7K/eDJe/2sOzUXSzgXwiDsxNlAQMxAidr
eLUS3XBj+mIT53uyCkmtdRYtqBc3P1Xj3P/s4pTsak/F/rokzoovzts0DRkO
gG3aiiogBpUjM/h8ci7SkNs7i+g/fYkHKvGH1vQkQL3z4q10MIjOtwJq7scr
WyJZVfhQ5Q6qmCsoCN1rqinkRC/KSLhri9y2tQYMwWyMvMiQOsWP4aCOeGHU
1Kgpv2RGyhj9B3gZyfjxpKD9wW5xhgY3m2D5cPnwEKC3hMZJ0vsP2oMAaEg7
GrNbt1x8h/2q7SJxNpX+km6RfPzt6Jk9gXyfLb03Y4Pzly89VLnxBFho74fF
ra8IBRT+A7ZnePUUkBBzrqpvUwL1FKGB518ib4fQWXQxK+mcREVd1+cB9A+P
VMaCb7g3m571s0I8vCtoNN3l2b/rDhZupl/aBBq1nNtrOvhrRrpDXAUsE/ER
6XYEWyUhLKT1uEojsShJ9t6ReOS3QtW4ZdpRZDsYyifSM8dF20N67IsWFkO1
hiG/9/gzXL1mjY2FNhM58mdgVRNIquBfX/FqgYLTVEWDBX6k/xgCLypt+6rX
PmTmXyHdbYT8XrqlMnzpdG7w5Okt30KFlbRGDOG1pgfqdJ4BLeW2E5JUEWDK
nxnsKEHFdWvpEMfxPDpJbIYyGomrJTW+ZeLi+R/RgeURo9dRoBtHP6S76XRP
YCjw6xUNRaXAvt8lJ23tadK1acgnWU8YZt5oqh5rqRbzhRmwNzEF9Q6VbYx/
kSsjdAleRwGYa8ODj0xvg7ZHbazDWVssHrJoyshaUvFcI1UM6cCcigQijeGn
MwvBnTOazOEEVyN8XA3Eom2z6ZIFY3ZAIHCD33zKY36jXodlgdmKWBFMkzs3
4eO5Zm3w7ISLTiPE4iPbiwa0iM4P2p6tcBsJbE06doQzo5uITqWqy+nob/ZM
D/J3dZE0l3zBQd5/FYz0tpApj8cVp/gBEAB3cXPMyX36ifH/CHlU8rBkrSy/
AF89Z9zdssFJYOH4CjzkD9jF1D5uK73jNGtgzLX8aA7n+4bUJei+83eNEft9
Q1gu8UGqUYdVrAta/X+MVmFG7te/fxjSJ3T7y0uqUtcz/+bfU2Udj6f5LxXQ
DQhkIjtPnuoYdeln/eA8N+VRdb6Y1RdwYQyNLh/TMughB5/66MBMfVFBrTrd
LKLrctBAGj16ZpMIqnpP/RTheA+aOActOUI4KTkw0oM1q8UuZ4nHXvjUtq5r
4feIlRhD7SVPs1Bwu/YMGlx4kdm/MpAZmkSx2743yTvQw9skQLpou0xfZj/F
XJZzvDcBHXRgTj3oOA2jz2rmMgGQC+yfI2SXBBp6ArzdsI0BBnaAFu35tcnK
DHthH5p5IXgaT2BGn88YD/DIkA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyLTh/DWoqDcFjiSLCs/3Zt1Q6ItF49/lxoCPjEVeARA8isHUDxhau8cHbV0j6P0fTR2Lq4gXUOVDwUafZf7leGUehJBQ3ly/n7TOwhWiEGuNytdwK61bUkfmibzobPmzrstTIJG8jbwwAcK64QvZ4MSW+7+pQE6AGim3Gi+nrbDRW6cBaa4hgtXvyWBsgHiUC3YHU7n0z5sKeqs2+bUafuT9Iej947/SFBBC3hthyDvlOSj4RfFFHZhn1E3zaebaVv+QVJps9T21W8vm+6aDQEixU3Zse8oDlvRY4v0FXD0StHXL3ERV9mahecLDLsBZFSHVk5wCdZZzDpNAlEWdECyku5sB/OblNd2aXk6ZenTlmiwPiK9UvIEptk6UlnvgDUBVCzDK3HrrXeKbHAwhge0e/y52FecPtyyRGz3gvq3ZRgMn9c0qTS8PI8tNoiI19skJC+StwzQVYGx2GRm04oCiP8JOBMZ570/KAxcEfawFuu+EoSF3ZP/GRv9zvHGLdwZjQ9t2cUVjUdDRzTZTCaeFwXO5E3gFVzvCZL7hw5FaPqNXAmM/s1Vuulq3LPChA7yIKyMP4fdmIACfbRRWW145ioIwSvIlL1BFo/UqUmuT+WDWJx5GMwdiwpghHThYfZXekpxSZxTa5S8S3xKAG1/rQqVxuv4W0kyyzoDHKjHOf4mGcHshAfZFhSFLSMw6BTbmtmgeCieC9/keowf8IZiqgYJFJOiAqHVcGmJy2PPN1NWqw3YhtRKA+IJhaZIomcAkYFEPO3hslVqRXtUgcwt"
`endif