// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Q0EBtyQa4iW+sXuHvmlCcXsB47LOJeHiARUs8CpJp7vZZZB1Mx85UMQd7PmT
EyCNq1lkG3d6AJaeFU61z/iO2r2XRKzSMYyLdBhZzUpLVK7bMSqdkcqFCxvu
Ptd7SAc0WE9i553PFtM6AS5PCb0ZA2tzYsOzW4jO2rQ5IQLazUd8uAXdjnrm
lSmuGdMjnFeLLbwev2bv03091vKzCy5s8x/MW6Hk5mVjCDj3btOvbwBUCSL3
w59PA86QajBpihwEzShKXpZaFNrZ1wtAQIXrAQnHehL3qf0a9HHxPm1hNV6n
lWtmUF882CO0EyRzF0K3jGrYt+uRGS6FDJklszReJw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IvUeLvlp/5yjhF0HzgTMSCpsVcVUbLoC+R2qFRObxx8QzZ8UdRLJjz3/Ylgq
xxw+X1VUAxQRA0v3ZmBLF+1R8MIO/yaUoCHwvoSJ8HocVY+LzgmepJEMiro2
02pj1yWNunOcgWIoQC3tQYeyvLvAgISEU1sed72DFCNLoUudn7LKO32RYRpI
2vbueMvHl13EndzRBGRH8T0H6kwDkYeO1xyPDrNZrRDMKKM09Cg7EEVyIcTz
RiZ4QQtln0WfaSxJiOxiAdBipwCgAweqAg0luuYrXpv6Zy1EVVqXX/sjuqyJ
soGt/H6oULl8sIMteqryIxOYaGKwPgLjRpBfGjy1Sw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BBgbYepA7ee1mJnCKz8TUOpjegi17Kqj59eqGudybK2QPDtcqf1f9sYrjLW0
WtushORvsW6WMCKurdWFQpaINF48OxLmVq6Gcy+S25GHs7ugL8LwRh90HTk+
m6nyoclU5CESCUXAgzDX0Tucd7nQ4N9xX2/SHdsLILS8Ks5aok42bMJ0Y1pV
BtK/V6dRHx4MMcx80IMXCz0H4YoeW752bQdizJkoO7jd8U358+TkiI4hklc4
E+eG4Pt86dZoIGW7owUDhQHvqFOG2xbTpgSX6/Fzi/eNWblX4QEqwAvzs2gr
P7/J0w63aFj4Fc10+bn9BsJydLavro86LP5y59XZdw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Yqj/3rOglpZza8POUO4ZmNqwIru1evLakoC9AxNvXmxNj1U9b1E0vAb/THtg
UINKLbthIGg/SdRtl0UA+e1wTCFdw0pNdWuCoyfuPbt8cEYWpJEOfaTT809S
RgvwT7nJT3DcQwOTmhejAPT55lLwypIlbBwjHm8gihybqki1vFbrYUPoWKQV
KIiIKuhEjHDbrVabci/iArb288jtBRH2o0mN/S9rhTd43aJbNPvgxYegUBZi
Vva7UhJK5sNQuooaECWmxYqV3IXq51TsfpW9sn5JDIvo4SWw6tBarJTl7nYn
1lb8F2W9XZosvGD+MCb1vzdldua2Y0jnAHJgArTEVA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JBqsB6ltqPVhGw5bL8k1pXg3FT7Kyy7nMViFhn7wHICYUt+HB+oHoo5zU62y
4bbfvUJ4kEyWnUXLcQ/YqsnCYmDm7uNzNb+qeYccOzbUpn/L4BvufcqwLmKJ
E6PvfI/0yIwlPEwkwEuHviCY+7B1nz0otWs90qqM/IIKKl4D71Y=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
IaAi9o9czWeksvR53q50Zdb2xO/duPCZ7rfkH7U0C7EtlaspwKlFZ5N+rUjV
2gG1lEpDpXVnv7jr7INb0MCp6ACzkWd5kt4TIbrXb6Z4y3wW/tWUCbdf8A+e
m719iIT53QYbyV11XP6zh6IFMlAoO1kp9eAUMTXTp7LJb7Sh453WIpgdmJHy
8FdDQItg3H1a7i+2CoxXY8XGokYMWz6YePAkJ4nGGLMRF9lW4n1DFXRNthEZ
YUckMDtcWvuWkIccIjqJL8NIJqjAKKDwYDe95jR5N/yzh5Di2FU2uKPraUGy
kbln0ckT+fjA3eYTRN/8/oazTiDDA8jRTLJ09tsIm+m3DPUiwa5w6P1hjhQu
zHdyWmy88XEuM/m30WChdxKUd1FfAzF3l1e699Exu0kwUcPPccJ/Wx9SxD9v
P2IZfx+mswG1K32KXCHz7Su19pHO5ExAxFSZXx0UotQwU66gH9R3fvoioCsf
XcCxZHYIX5ls5JpQMMqzsOg9AONQCyUw


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dvL+gIaG0wnlndf/hqZgZgshOuYrLkt8nzDhHOypvDneT47RjYdO1Natfk+g
IuU5PQfvaQp1jY63qeYbI0LHV9GSe/Z4nSPOiuFnpSTPmH3bmb2aaCEeivxb
hhqITTkLue6J7hV4Je3DOl3qL6Gi5MhA9C2XZ8YLco+Rts/X4YU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tBUSS6FWH7NQwZaloYl5BCK9GfOeSoO+xii+/SjIhP4lKyZm0XP7GzdfAur2
zJTR7gOZbzXUsk1i/5k/XuKt0g8SwjE43UjXKQtKJZ2LBrLJl+u/sjiIqu5V
WMdZmGWY1IyHfm6JJmvIWb0qQ+w5uQ1jYMiBy/ACKSByY68lhLc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 11792)
`pragma protect data_block
pxxE00qVf3g47uXC7HvONjBKFWYgZC1SY9YB4hyivViCubCpxH5dREDafe/d
rV1sCi4zl80tvA3w3hFqJkaA5IIcmnjSHgU9YL8AV6mnAEo/FPh5BwRk+jYM
UfjASWKyEdL9zJIiZUHcjCquG1XNvp0VpqJePSKUnri6LGww2repCk5E+61S
SHpk5viLV69aPmdSsrZjqEXqYSDU0qR7I+kKTtxffTDVyvDB+R8yFVNkYThj
UcZ4ls+BEWN+E/Yeu5J6kG4gfj+rjQqg3KVwe4py3NVhHrXUSt07aR2y6h4/
e22pVnotCCnPjlFmtfShdQtjduI2aBudzgy3jCirhArwmS9iBqX5CVr+bHqh
6X2iDWfoh1H4Bz7SblDLFnaVsDLaQNj0HhThe7cPZm9FPoKUymPfiwbqw1j8
m410Io56Afs8SXM++/8Z6hD4jSRgTaJ38Wl44cA5jkeCgyi7XvdSibjtNEct
PSr30BQeCym/WRhviir17TAqC4kqaAnalRYA0V1q+HcbxOVkB1TwWztdgWaR
ZlJ01jkUcnX2GjNVEHSwhA1IcazzDtugb5/GSKNMarrAtvPGjpMem0Gm0moh
dLO7q9pImV39GOljKd9oG2j+KkVLW97FX4JOCu1y9t8qWIudW+ZnlYxwxmZM
w9LoHl2kLmsuAUY4eaAV5Ztw3ebMQWhew0NscaK2D38OYpEsEqKr5Cb3ajEO
Z/RVESRsqq8DIXBrbh6kjUdKForlL1mV9ZiYMaP6fryFNseHyEWz0VOW1wlW
Np52KenPss/scO3OZ2Ln7qckCK0cht6IgtuAkY+xiXltkSo3PCWBx1wvOx08
tu93kWsz30umWYvA0Y+SC/rQJYSQEAmJxoSbKNd/nuaxRZphYJbJzJ5MBOHT
uL2FK8lZpZhb8jaU/6lT2TeE97yOsx3n66En9te910lscojiaZxG5Nnp2/F6
hd+OIlYwUhvZqoyfW9d+OrPaN9eGjjtqsqbQDZw901nJIiatTkq/YHJ/nlK4
sVBsKonLDP3pLUiDORSOH4YpcUbWwVuRoOa+B3A28C6Y538lbFMkW7m+JLFN
CcpIIxM/53VxLQ9dotr1ezUVMhad96OECiq9F+bAtGO85JTa/qwqT7+UW1Yj
j4jHuo65ww/oXtkh2HBqx+DJZVAMChFM883sogN91fY7WyUcK3DMTapJLGr4
M+FL7OXFhmZPuOO8U5YYnnsZDOjR8cNmm0xf9ZxAOwqmE8B7pvXBVqUZHZSk
K1j6U5miN7mRb+aHBsSB0OLVF+FzJW4UiZVKCCBu4gM2omU7aJTl1ZrF0IWS
JylnvYnvNJjqlwTBG+WaufGBTRFM2IHs3jcg/Xg5j9EY4b3FwAUIWiJ3ORkx
rogKsFdpREmTvPa4cAUzqitecH4lnzKxX4LW0nImoX5TapH8VHQZ2voSX2Vi
1ntnq4ZPN7Me24RqKYtJkBwKVZP4b8u41iwXEsEfq54R+UehB5HeyHWhb2dQ
9O+eKSz5k8cr76AKX2B0ytFUB93yhkRpWktYqCKyqc6p2mhe9pinBDFoVCM5
z0F+BH3zr0CAO7vJrT+LCLOislG5RmfSv0aSZtQlrnpu5czFAIVjgOQZQFLg
KNMx2b0znzeYQKIPqOTTBA/Pn2u5MIQAmoicnEf0i+1Rtj1fzp26a4cklNZt
kRJTm7KpScEJiGhMUM+Ku26aP1Oc5xkoN+JdRo6LFcgh2+LmHTVX4iaxLlj/
sCz89e+I85D801omR7XNKr9RiHCcQ8tiVpobCmb3LA0jHFvIxeenDfkVju7y
gLrFLIq4NMxnmwO86FnOgKDwH72tdOm1bnoV3mKyGCFz5bFtpG0z81mCTQN6
8H3aCdI1F0GNyk6ti7ERlRcjWX0mieejoM1mvKxPpTrHtGIANj1Q3IpgUQdA
sUKhdEOS0JX44/Rxue+L4xoj9bQ0Fy/RKWh37Tl6zMXmqlTkGXM6Xtn4jX0h
hLSptOiAvB6fOuCBc5zz03HtTy5P+t7zDhUnOfRmpNmHgvh+EjYrD7L4fmcy
Jc9JCx2D0XffLkGBNHjU2/Pge91fVj+T6idOmBS3c7Erqsqz90ZQSQniGxvB
Gcpgh7iEPHs0FoOogXNnZA/j00QbyMiB3v8l/ACkJ+HrJSbPOA9GawpjbTIS
vDGL18AhQO/VT9uD2NDLcw3KkS1A2jDCgobYGlE3Yl9P6d12pULyJFIp8WXU
EjDP4G+HlRr6RAlt7Q6pzpIX9iWQE50znNfgEyfcgIDEdd/TuhS2H7qkETB6
tuA8S2msY0azFvIr66ukGvBGC5bwYDXU/rFMweHpswTpKYTODGk1ZTTFeRBT
z5B9A8m+pxY/XnDK0NRypiBXVz2+xzeYQ9mAwk7ODQ0yedLifZlF0nHUD7f+
B4eqnCM+YVSIcYdVR7h1NPQ9VLx7wZM+r4goXu7HwGhlc94coTHI7tOwJD83
KQ4GuYBEVZh0COB/W+81SEDNtMxQ3SsNkLHj6v21yowMjZzgwQApQhKjFkBO
UvT3nKJ5dM7jbt/kcBJyGBzgZk9kVYaHuqTbOagdxQy+pzTP3j8b8itmrtnc
nCpahVDe2ezP39/uduAYlZQ8cOjmFqnRwM03D/YLa45/A8trfcDgfckRjmUK
6DYW/WdkYADpA3UINIoDC0lnk5BwOAZdFM9is9+njlK2KWM0MM/dR9piHwsE
lb26c3Zbujp/uOufj9u4nLfKIJqamoCW0yhfAMWX5TxNFw4hE/iDtcBAmP5V
Da0kNF43eLiYtFFzAKMGiUp3VGoPx3DI5CwoAfHWuq+3HKhiCkLTO8gtWQxi
4C4wx5bYeZsO48WWXrnt5OI07IbnB8MgktQhtij/vx1tK6DuQThXcMkL2w2f
ezx9/dgVPNXysaNkpfnPWGFPMWQ2GMprrrYOMoLhJYYvFac/4zqdBImmEovh
vXVTiz3bkzKst08zWO7qdn7+dNsOFS3uZcO6JwMUX2KdLpFgve4W+asI63p4
sNiR5gaVI3FkNbky8Wspjsk341lbV76d7T96I0PYHvU7WNE1kThN6Kr+ZBQE
TvMQC9glerp1mTbmzI5RwFRAvAGrPpoeAz8TOmDveJ4bjfyLR+4XDF4F31sQ
hIvlrZm04RYXvMcfJRsIfPnvu6Lx11EhF2XpdMd2zbcaWhDWGTpZkxTMcvTw
/jyTguQqwg+lod1unaTIybUsvO1kJ7hAKEnD1hl4hFc8mAraCguaVuPZGrfE
rMuv7LlDEuOPetEvOKOD109W1MED7emJ1geycGIcelfeq8UF96DWtTfYnZ+E
kTvSeFZo7htMYCW1l2R9vLFINbv6+xxERZdsEIzyupmlqZyRvpZLSjm3yezG
/4EP4pZq9gi5uGNXJZ3CueRzw0JAukiH7QWe1Ajg7ebZAC7I7Z+zfFUerW+6
cuY6t60+xiiY/hCiKHKeLv2/88plrgcTjF3OheIVa3hCSk5V56VqPXXHwa7J
bcODHJgtoXl5H9z4A/0r4cu31sSzmwK/TnzhSbVcFeeYFPJXpXW0T4HjdclR
jTZn5Z2KvRWihzN7OhLbza/7y/Ix07k8zjMTyKhgOxQkCUkZSGP3yDRg9nag
zLHuZ7VEX8hhwCwJWnwCK5l/z2N7ARSOXKi2AGsdjFinP14gty2MYOUi8BuM
pwQKUyMU4DDb9zRr41zksuc6aoPkBLuO4SUgRKQq6dv2shJvM7Eyl1whbuyw
+fejiYjPRAQPEr23Tm1mUeGpRZDuvDZz/MlySy9QQoSlvS5NJ9Cw6oapEPFc
LM/1ELHt9CVxgIIcDJvKKuZ/tLcl+S9XRPpK2pO1FVfSwzrAnOc9jzymXS7f
Ba45aqvIeOYxZgvLyOQzCtmXB+DEPuqtQIY2QEMIPy+tViUBR+n4IY5bycxb
uvsKy2Bv3w9ZNuvnRo56BeiB5E2Xfhq5QpR0NtXOpB9df9HfkPThENnI/i+d
PLrjNUtCN50fNpwR2AFfrjAL6eb3pH0uPnZ2MS+aClpcENJWApPAD/rpMwk2
MSObMx/NyqAnUZhrqob89ezNbwSmNteUhv4as+2UNQAlIKieBq7zJVOtgk1J
U713Qp+H38ltLWqFph1tR3fG9uFN44+BSdPu2sKL4BjDziB7VWT29LAXldI/
zPAmdUujW2eI/pcfdwWSp/QFlro29wW37Sd9DF04VRQNGVH92hpQ3WfPTPov
ipYVRWOWtd2NH8LI1DhZuzIirvuDkNhEeK7kxsTih00+MDKKM2mQBMD/XnUF
owmF4diSBuwjh2v7uc0Hy64961VtaFRcNBbdoIQSsObRKcT/zd/lZH/1DoXS
yeXQoey0AU5JEO+G5cM45whvo/p9VTyx0GN79/LDDssBGsD0zS4oswASvhei
2kkfPv0bVA1P1ubnH6j5/odzQv975JxyUWADq8mDMo1N2MIJzipxaZPTU/Yy
4ARjoUk7yFrcVfAabEANr2y3ET86Sd6Ppu1NEgkImUMjtpIn+35t/CxWnECK
J/S7yp+rc2j4ilixGIznbNv34Gc6Qdszuu3pzstXpr5/4Wj/kRAjpZqDo5Ti
D9Pjc10eXknzLFFHepDBFtp8LOYofM5cLMJcHzRxMXXvb1GhxTdLYKZ7nAhE
XO+Le8g3X/P4gLp7Ic93jiRY7ehJrB4Wb0fHwvhi5xS4yYIHRIFA9x97rk9g
I8ZniG4ROb7pBllooHrL7JYAquT5347Mkqd+SILMa4TbJXhbwZEjDcEWDtyB
e41rucMJIcEm4C/YAPtmkhzdWM57Yr+h0FbnBiuwFAh+tka5dPe9oWif/Ws/
bjsM8cQ1xpVw5+9MeEUS4WiIUossP9oY54gdi7W3r7K15er5Gene1yyu4rHL
N/KlGs9Dij6QsM0Oso7Ho5ikPAp9ivVaeyZJmcSK8PCdKFg/rR9mcyvyd49h
IPQACasZrQUyZT5Jb9ursB/u/z44XF+nxj/H4gjxssfSZ26rNE7pqhITzeMy
HGtvBpfi+Ulby351lWEVdkGZCeuMi6CsvrRdXtvN53wkix8KNhyA661+jTyt
iYs/IZwtjWv1mOnbqbS3QoNNsE4DZBtOxrHs8J3ueHwkTDXYSkLN90Gxb5S/
y+BWUlL/DMVwiKr5b273FKZ1AuLox55wa3mH+kUTNqN9JT5BUt6lUOwe/pKm
oRptK36x+DraS5eeSuOtkV+oX8PhfcCEE8G/XAXWhfZxygKmbLeMgHguhPBP
kHgPcs6dSjPod+ZCBR4YtupV1/UEx2WEqqI2SCYliuoQXe0VYoug5jZpENI5
Jl5Bt5s6ZrMC74jrCJJHAdWMxDL/wlVmxivqKpY65qMZeUCHkp2YmdVP6oZ6
m7FIcjQ9vUqa9zDFWoKnu6Q+zcLTv8YtiKKtsPwob4VMq1EoqPC8yrnSUbIq
qra5LbWKrl0pwCPUKdbzsB8zOQqov7R61DKIZImB84dVuGd/lNOuU2aTOW0/
w/SsZSG/l7GlncYfz5wMQ86wy0Nto1gvYvpU8Plq5F1n9OTU41Z8BKCy8GkB
8jGnq7hNFe/io5mCt3xmBEtLWqjA2g6DR66Vxl9i3+8BzLyRVeXjuDrTo4yR
036/Hq5IXlWcveiSxw/6jk3gzar4yWP2TGFb2PtPAhXmSii3aNVVhWvPO/+C
LNKaVNtX5i14qeXFgHyF6gi6fivBz6wS9/y1fvzBGClNK+NG38X39dUd79oA
37nJw0v8acIjJJruOG5AHa+9yezNGuWbE/F2k4QWfhwr50nYrcjBx5yycfLz
fcQFkA41MokOEoUB8NE4iKOw1OzGpXRgSxA4jv0mxVEDNEKV4sRni8AppIwJ
oq0O9tjHX2tjbDmmi319l5XO0blqakBamn1qxWF7sCNkGrFCtvfGpzuJ9XcP
cj6ZJlTwln3wtaJ2SbbeDhZS3bRmMPIR11sCK1LKRtJLCcUUelayJTE9u1Q/
1KnTn+7Ufys3DlJvlwyBQwRhit+Weo9JmNgihOxi+cw8eu+DLd9qVg4gOR6m
hQIjTCKXmHQ6FsZm86pRXou6N+51Z+BgzpdnGBzQtaPsWh/L9mpWw7N8xW5I
mkN5l2Ea/mEjBdM4jW8kgvCLF7/lndmNsJ/SzIqPv4iDaDceznFGs0kc9a1r
N97zpqdTXfUyYjRQQFwK3lRjP/7l2tKHIKB7aguMLLnnnGE83HMahZqulYE5
QDLHnVCNR41oFGRN/pyI16gSuHUrRc0DJCo+NFwcdglR2HvjTKJGn3IzWo5g
+lAJdNDzr1aEKcMJ09iheJaQCIKEtPxR7wFqWPoaXCcPGQO0PO9I7Sc3EBsh
KUPKn4L64thSqfqYYeGbdxx4gr91dLbIsWL0v+nPN++leMoMmy9uG7qEP0mL
Tp5L+63jnLAblMeOktrRuFE13RO9RjLPmuqSYutjCfW6MkYyilctO32WLSnC
aMcStSGXAX0bEBT1t/8zkjJSaFXfd2Iqo4uPefTz8Ky3NNWNoJLvqLwIiuXR
Z40La3rRUL7dMtR477qCTHaAqclGMZ4aytSNTpmasz9df9bFtfUFfrn6WzwV
eKVLtI20DXiC0jZjao4MZmOrEG0YxVSmcadS9J2bDxyRoVdNGEhDn/rhnk88
STTQjNoVdEuR7FYPtnjYCAO491iWnY/vWu2/dT3hfUYz0aJ9cn2GDNbcIjXb
kNSzhNwmgZ7misYr+rGk9qrnqqgsZrEXtvhIvPlv12lRViHqv3OgWS+G9tq1
oAwZY30mJwdghDNgn0G/epswFH766ECStz3aZxFzC8RWf68dN35Y1wJO3Xix
9GPxR/uK3qYu088Op2GwKCcmCNhdC6fCh2zAPru/V6QVtsJHlbVlOlCAJL61
JfkclDQzS0dkJ/5Z69hs2hqElq+N95d1dJDbKFvjnNFpzDiT40NbCUeEBgof
MYtP+uZkx1RLkHKC3w2xMFWKajTUliaNdKjARFZ19fEIPOZRhbK4Yd5HVfH2
D/WL+RikF0g/uaitbfMPlNEz+9a9JIxjmTbFqT11kdJgt42qOo9KInFG/d6F
PrHZn6DmZD5vH/N4dgDADWOosK5IS+AdUmBEubnVbNEysAUbexQIiNCLHJBn
hi2vyiGFKU/JgFhnceAzA/C2KkdAO7G0CoJ8Po4dZB8o7odzPCbpYI5h7kxC
wpcPyYdq6+nPXrI4Wvj/clBJELIp+64dt08n8P522UhpR8vclN/k9ZvwpOhz
LFCGkXV13j4Xtc4TVvLCn7uVMy1/cCTgQ7AnphpYQ+rWPV8tcM1LyldV0O78
Iw9sOwgXLOpONAb/C1pD9AR3+5h60g4o08epXnfLf82akprVi3Ao52WhLU6/
Lk+EOtuBzJ9JSzyBoMK2YUnzECN+olfh1xLe5HeYiuRHV1drC9HF4uENDNA1
ByTPBHBtYJ7Fh54N/8BwlYpNRaybi39EJZzn5T+39l0YzkFNZWrxmXhfa3qA
cBRAqGxQJ7O8FsOgLYPDHpNJ/MbwmVJTkHl/3rikOkWvgH8yF9xFdZOjZmBi
qctbp3uF+9df1Sg9oSlNHreo60b+uqWQRavAmYfvm+zltTp4WAQNQOy12b4v
ifEUyAgfulTRa2ungMhTg+5SCWvlHRVjSA4jicpzCHvEHa1F61ADk+HEooHs
aLVwDX9G8g9hfBwp3JQHjnG+Cy2eH/TDqGta+v9SzftKulMZ1nLNFIBu0k3/
Zkonm12BZVOKpW+UGoBgDKTBunSP4ficPGLufSOK9h2GWzT5rArDjA39ONrA
Nrn15w0IsbETV0eNEZ2sWYH5OaRQCWHg0i1ZX0OTfh8ctE07T1aq6Liv58nY
dCecQhEiLHN1B+XDW9Dcq9/eKkj2xtHe0y7aBFfhCJpl+Vc6p0M/iN5093NE
G3RS7Uz3Umf3smOUYTxcVXxSYETih5GHj6VlktowRpl1NudnhMDxFNb1Pp4+
shGQ6zVeYJEKdg7qWO38kk/lkMnl8kC7eQkABdZP9l7jT/uZp/vBpvun654M
JNiJ177cj6BS3HoqpvqwRRRXkcyIO0k/ldZ5X1hj7NHIPtiGMd8W6SnenphV
dwrt2ejYcH0vN833IBgNWENn8WRbLiLBwDapNyPcRJcvqyvgW99onI7IQD1X
2RZJvTr3txHZlxOtBXP6SwBr3FrrJqrf2b0+zq4RM1U5NK9YqfdF6YypnviV
5n+7zddQK/H1hvbE8mUiJDL1WueE+kCS3HHKG4pB/KH479m3pC7iIdpiZZ6l
arLHmoCYPlFkSGddavCnq9mAALevilUMUtwwX4k9a0p5spHusuP4//vHsvZN
VGsFsxOGcBp74slJS7K/J38nXtVcXzg8dcUO/FDWeorR1Ypny9hDofmsuINz
GJj8lyqMBIP+7Y8QAm5dnjOMNAzdrwIB1IFMfzJNsYTBW4ZAflv6JtT/BfwV
S66dZTSlg7qQz9qv+UzKjDZXUgjr2h8baaVoKdcsmmiTzYymhNkg/5METhK8
/QkaZ1S/4wDDtVvaCpInQxyPOLbgJ/REhzWA7S8qGG436pSJOEV4daOi06NL
jqgbGoLxnYZ8lfxN+5jTyn+Yf35ixN452tZFOK0A81OanfousNp3ozJEH+GI
inGreY5xAgBtJj9HeWA8T5Edhjq2E0BvB5mpraM4VQunfEDLjnzJF4ZUkAqR
KkVVZRh5vM1M30xJkJaOp5AbjYdY3oh+8SAEH+UiNPUP8LjG7rkOWn6hHzfw
nD3nZtJdTQyNVkG00SYBfS6cACe3F9JsqbOEwBesKwbqVeyLPb1ckqFiNeo9
8ARouyTvHY++Cj6VO4iJ85EXIf96srdhTkGFowIyJBPSt1qznk56iSa9fuQo
0XyGYp1+h39n6HuX/3y24W1NHUzDHJFLebVsc5+Cu6+Ws2i0+W1cMw65OjHh
wkev//APVPmpiF6UzUpm69TBt+z1dvmLvqEwGjdp0ll51rqhnxIs5XRf3UiE
BG1cDsdPFJy5SpyWj2R77AO9cZD4Lg6GJ9DMdzR9Is8Mf2M+RNhDno+MWA6Y
BQezGDVRN5XmZTBImpjWEm2qPdRTKOTZ0AEgO0Q4KIzI/+4gUw93P+ZPY/P/
QkxgZcjkwoN6hLFHTLjmHTIQE0URvjEIGydpS6C8qPZVtLHBHLZyKIV/y1o6
s8FSXNiXZQJv9Su+juWp2DCrXTSJbn3jLKGONLqQ0XtGIWwI1Cy/IQsiQnMH
mgDJPDx/myhgalY3IdoFSdr1+IoKU5nmM7fmiyGtlj0WS/x3VSVPIsd1BiKN
lSPvflJUxVZ1qBemQiGSTHZHpXcAiphNB3y4b0k4TtH0NX/7+rjZb2dldKzu
7javxuAl9j2zSmJq1DdTbbaOvv8O7TPnZaRzhQPUZB6HeQk/4yYyWgCVMcxJ
vsUnfG++VGkrgEFm14EDeQE65kWnQ5nX4hr82rE76DOBoj29CNx3TbqflEh4
6DCZYQrXSVFk4wsGC8VABHqmvwQ5liruKDv/f2aKqHJEVo3KWa8oN/7PZDKJ
rfj8gi8FgP5/2GFFGeKN4xjeqi7p7Iwm265f19XzfMJFbNXZOJcdP20bBTGo
9YzmDA5Bc7diFUs0UHpLi4nWUPG3I1WDuqTbvkhTSw7tb/d8sJI55Wx346wu
l04UCBQgLQLoMGETqiSsHn7MG7WkclSazVZNNzFm6H/QSsnSndsO18TVfInb
/zhT3hq+FUDQQykSN1OKYdpEMLmxhOXmdtYOrUNz/vEiTjxkVtBJjzitFR2F
aq1CWWPHjx4SsgtguG5nH5zuN2o0XC9+kegPlRSUk27vPHahYQI367n9A9NG
1pcoDy153tlAZqIqA9HIPu0qsF4fIdbGdoj6a6bJmqNERZeuMhVsNEtvYsEA
rF8u2cswBFF34pyQboNxBZNHQMsqTMFVvlUoojYNKRv7iACMr9BFi2u+8uqb
W6JsnO+rsla9Sf5vJKqcHH9fiDQsvHCf0EZFfJOXFEn8GJmKVePNuIm5b5PA
Dp6qBGyo5xeh1FxeJkdlR18Mp/yzYxU3cw2OEVxYatOd2Dpr3eqHwJ5Vk6/t
EOPIbGofLy3jIRb/ZTRaIqG9Bsggj0LS7bdJ60r4bMAyhUXQKaRz5u/VApRq
f4wf51YGkGajcG6l6ItUQWQi95slLFcZIl1nVAoaZ8AO/AHqAi4NXoOtTHfq
RIwrXbHnEyz/fs4y1VlLwyc/HlE8AvFiDHE3jVrD++Le9gp5I3NELSpeMPw6
4WX7ObWyxuNHOFbgSXg90h8aHd/sUESf+vJTGgJVveWgV3YuNi1+90Z2hxyr
kJ7gh1cU6fLJmUY1Ahb+xj2+eaXXcRO0weq+2uGUcyPjBtCgRF9trvhdB9UM
kFHHjdobsMWcgt0TFbAbI/Twe2V7B9Ppmwl8Gscbn9i6/RBglU9udruPnY+d
p40a9f6m6uNmcp4PKUzjAtJj3NckEovu0dh12Q5Tp2ipat4IuGdDsMHiMJn0
qkFXhkcVSNfSU7W5yttvlnWqZLWDZvfeFVFVPs3TjNBAuLm2rToyUB1NwRqY
hO03rwP2uo9yZPVnwAuB4hDlkK6orqXdV40vVknP2xlSNt0JgwlwMV6a1/p/
Q4E39O6cFVpMFVle3R4kSDuPWygsqNd5iSvhljgFA3Etizn9fC2W2xy4nkBD
hmtihWM62kTZJE3LC3pw+qeTRE94aG5uWpSkJPxSZN6MyP3vFpkh7rYLNT+Z
Z8p19GroxV8M2E3INtkHUShHjKFzkh2GpapiYysJ3W79yvpsTCD+jKA5UacB
CPBus1UG/5Dfv14W/1jbzSKTXeQSInjY4OQwjnuy7TaU+p+zqFYOBwO1OHj6
Mj731MoCGA1uhZQo1eCQRJ3RBp2Q1Jnrjg2Bvm1oSEQGSSJkkHTnE4UCmvN9
C4tYTKqHTbf0qQfQa6YibYtOMtbYsCIfJH0OHUFESQ5iVHGiVuwinkVf9LlB
4cAZ0COYtpeqLBnVf2+lg1yyNy1a63D2RY/ctJ4+pXGvDgvj+1T4b4oESXpW
A4Hju30kkR+Ewihfqq6KNnR/nz6KEV/eifnA/ZhbRRMHQmoGg7K9rIfTaYVZ
fdLsDW6kxywbWobEPoapX0vwTDSZy/62FF9KPK16aIPRJT2RxbGO/TMUXHjD
cosf+ONeckRvU4e9akOmI+M2mSdsqYuoanLnliScO6/U9QiWbXabPGRyoxo7
xjFwm/BV2T/i1sB5v9JXblpuVSNLC9mW1K6nDN0WvLyN0zsuQ/xX5G67tj8+
yDr5bhuzYkIQPcveMMjl8cORmlAXUDqIEiR1MldOrfJH4aVcT0uJlZMnC7sk
xVigydyQ1MpG5uiS07RJ7UtDPzuMplNm9JGvhw/yCNWIwjAJNkWjxLH7LMNp
2bg7Mr5+fHkZ+kExpnQ3EO/2/oh42LYE4m3L/hUhP01aSue2KkuKJx7fv7kv
1SjTTN6kWnzouXTJrcddDj7EW5ogdDN3egDh4xKRSEHlvf/T9qiaFAhvhc2d
QfSeq3OF2es7YB+do8KKXU9Ei6EBqNSk3A7gE0VJd8lFbf0005UCUuMaDzme
NoYeKoKQjzLZ5SWaAoXrmA1AsVVGUUPwqGbXAcLfMqjlNIWLPXZQRmgldwvp
5FhQym/5ssMLWn4OmucVN7aYgb60wt8NhEAA9FNI9oTxc0QOGEBtzecVRxuX
do8koJ7DvX9X+JtNjchmit2TYEUEqHu9pj5Vmnc/2MaxkNtQ1fCcuBSWKZNm
SRvpF4hT8irSTUtHBUj+RV7Z11nGfjWp7kmAx/TlfgHXGFjmt5z7RMMv00SD
Xy1Qi9Bj0YxKroOBmidRMMToHyGeo0XC4wrYEP1vGKH7TC55cvpFOuPOUj/m
4tpoqNlfNe9R/ZrN3h6S8aCLkHg05esIoKI40w61BXCREVn2vi66t8LS5pLs
Xml82mc1fSy4vdD9xh+L+hmh2fe5YNN7hah5ABhPK6qmmR9fjA8Bvdj396WB
2a9xNwGOxIW2DS+Qcph6iWCwiqrbnAyUo7G+70ITd84hY3lnBgRc1J5cR1/u
WeluK0tRwXEjvP966wuttH2XeRd0i4t0c11h25ZuVjwDm0OvFRONxut05WFI
PBgvLnN2dJmsaVVOhMO0tMzoDwWk0NXieoCJ8wSBOAfTpw/h77j+NHlPp2AJ
Sk/bAt6nmSFcb5m0MkeZsUBU7m+ZZ4ZxNwaOPuGe114Gn7LLFJ9LMjmyTcYi
L0VTnpFvkaumxEQoHEFj104LigWb7CKWFK3BTvAAYaTutvgyQDJdKOc7vw6O
u/J7eh8Asszx5kdc/9aAbgExXboh8fm5GmStS5huY5hU6zB+cwTM3/Ux9aoO
PnS8DbgQBmhl4tJRg7vr4oF4Fsn7MVOerpvv2vPF5EDsEIWDDsLU07mH+5hr
uqj6XeszCA08mLr4ZK0WCG8ESyodlrF+/62scW+oZCq26N2aIEIaejYx+3vX
EsoHKwwPcXSVojLJYW06CKA8W/6GI9u7CrLmL5O4xYkK6lUEnfSXCYTRX1y7
bMOovvOpChKdVk+mVwbEzXT05Rr/DQ2osm0KAojbZ794mj4/iTh25YVl9ef6
1ulIglooFXzneyCM8WbbiCOm4vCcpQMpdYFr96BRZOtvoGhHiGP+KgwWkgBR
/TZPvwITwHcB05nPNsu75riXYJ4F1nKS611D1IHqp89afSSfwNNThbg3Gbyn
9RlNYZvmRHEH+pPk561MjH4KLx9TRKgHoGD4j0qtTZGAjTRZKAwHhjtvmVeV
Btw2tH2zDZ1MmtNYPfAVbunNJHJWId5YfX9d7hak52R1UNHdUErPxdMpmCys
FWoh1SwX8ANnhc7UM8oJh0sFbnkHay7CaFxI/6vSMUjNTDc7vW22gWhzJGh3
5LKQICecejuoSMphXiJP+NzmU7fEHx2EgRz8YOTVzbYtybxfc3INjqpez7u/
5GXzAJBGx0Bpm3OZ06lL59vTFnv3HHL1orFnEEzvjTkaI+zhSQgYdwZczxkK
mzneLMgvwtqgh/UJH1R/YNQvtfHaUYuakkOhawHK0KQV368s7jv1Ku32aVQE
7jYpiZk/cg4HugXEtfyLE95VNUtB7iGULsDf9TSlLlpKsEWoQZN3O08Hm4gS
nKUN+pszCZ8x1CZ3d1S/4JQXGWVtXqGXfu6SWhScycBm7ZS8D+ZR2P0D1T4R
KhOz0VMjbDDeTH2wDRRT/O8CeqRU4KiPxV1ZO9cvw4hV9EnyfjFH92lzQLxY
f5QJP1GF2+Z68TCk44NjUIO7MpBcVn8IfHcmCq1ZEWap0CAJGOd2NUwwg37P
WYUiBeurxcm3/fxGJ7Jr5E90ncYRXPOuJ2s47B6Rc4KPC3lrd/J5Vd9usoPF
EznvOkEVFV4f3WGpNkQK44GEdbw9pCqrgs+8RdPMOMAiVHpT0VO0Ir0pnyDZ
J+J5M0nJW4SjndBVmdgB5s0D2+WdK/mqSuaLxssx+ERqs6CKPbRMV3viUtIm
k5nvNV7DiYVhniQmRA3EJUeaQXm2qYkzJxqV52x0mXS0MvEArMtpmlqHCBEp
IkO+fuWZKcD2SQWJAfW+lx0PKzNcXROff+rVYs4f0TaAN7Q+UZxwq2ZK+LvD
wWnokc6Aue0D/eDijc5mvt6EgVJQ/WtfGF6Cn1i0A2m3rz0xOcckHho+tf3b
dBjr2T5Vo9+J428nfTV/q7ymcEOXfnmIoV2+2rT73Nev/plIeJBXt+Xnrjj1
3X7si6TIKgjCeFGZbH7/8N3mqSeGGzSSPfF52gXefmqmJKRpSSRsj6mhHmwX
YJz3MPR1AQBgE/z2998aI0IQbzt+1ddrP+v9wDOryk8qWGeM+rhC4VkjVQKR
5OvqqnahV2Q+Y88WvPMGqMbckj7q6QCSwrvexDTksgHgbuaFiozTnA4Lr3WN
C/MIe1BYkmon78ELxm8CgqVj7yb+vNMlN1KXeBCIW4LSTx0JAW/O27u+KtcT
cmYFYwBrkMbyoDQhSnPTHjN3YblzSRWJNcR4Yy0mRXNoU8Pr766K3bk7ghyL
WLY/HUh9HVtFcz8MK1R/ahLuwu26gPeqHiLVMxYk/u0QYJsVeN/GhtbkKPqh
E4/DAmX+Px22c5vIWNCrbb4Y24Sn7Xk//co/sKBFxEMhUvQCUQ22DDso/Vzk
QojOQFzT4NYEH8Ptka/rmL4lfFswzv2f866jOH4ufM9qj9jAkHJKVPIUr1bm
WHK6ZBu0m9mj6Y/ILXN0yLQeSD1C5hBT2qe/19lt+IvoDqKJWGse6LEpOVAD
VItAkjUd+DM0apVaW8BI4tJnrw9evkdlj8+622/lux8HZ4gCF4MpoqVQOtXN
8QaeBqIKEkgLF33beBYVhsYMUvqv/dzNodxj6RvkojDVFenGj1F4R06DlLK6
5JHfNsXUHGZQwUFmhy7w/q5SeLDzmGdAoflHf5tOzfZX7I6OW6WUEoiHQBog
ELSGO/2CtPVRxtACkzhahAn9/bJHGNe1skh529uAkAMSALZetB8RfgCH9uTy
u2T1CInFKluA370tRu5CzcubxrRwK40FFO11EipnFV9NA2F8ZQBx1i52KJUp
Gxtmg+07+qNRde7pab4Bj4tKWkzITrVNJBw7R4MUJZsuDUp6nHlCLg8Mnmqx
ZJRNaV5UirphesofxPl92/Ei3ME20BGVs9LPi7M0CWS/I2zhAn7/TKTVDsxQ
qRi5Cs8oWW5mj3IpXUpKRE5vC91M02pR2D+s60xseszch59jkX9LU+HgHdvf
RZO/VEThgzHCrfLYTbUmNCHbFeI6akRIJQIvlqsd1C8SnPPX2BV3n+JcTVd4
1gKkSzAvgUrNy4+iP6dKMR3rp9lcoPwxmh4urhow4ovrU0EVkSbBNOqIHDkA
tx4oIJRqLpcbylzLQBuNKr1mnp6lVxYlRFP9RY3H5TEi8IaHvMCvJomIrfqG
UkdFnOsWpWJv2gog8LZ+IyTgr+Dyz7IRxvYwCBwbZ6ZFFjofc+QyNZCnQMok
FtUfm3QxKHl2bbuUPi6nvatHpUTm7PsWn1O336BlcYQ+ipTA+lsFRK4qae5q
Rek87buPRtrP7kPMcGax7MrrA/0fxXcyJF31+AWkepzfIUJQhb94B9kiSIaW
vo9rYgcqV8I3dzoPWJXKROR+lD1WOg8A1YdQVQLZzrvm/+gQbfO4/EsfdSfT
YGTOVpjGL6zeWA7PeM/LQ/JO9Z0Ni1QljFH2r/o4G8Zjk1LmNBrPH8qp5oGY
5WShU9Mhww1a5cKnAw/t6yjnq6X9+8Pq7ELQFXzbYp+lDvpEGhH32SUvgz1G
VzIkAOCwDd2XBuXApmimPY+HCn+11yOTKJyj91MzzErayfkCLRYG+RTs5xU2
37f0Sr8G+JSIZKqqDr80iJQ796fv4XwD5M/03j9eUiszuW9isThRZ9Wi1xfn
vjQwE2MxdrKS2qVzNjWYyf9gsPiSd8Kn5HogHTiqN2GIBuGinmRwFjNDsfrE
Vnh64ymKO4WwlZ9jOXFgcikhY1RNLiQAY81Jv/A00rO/+PUCwtySSj8a/M8b
vp/7i2IapbIWwRvHZrfOHayE8ciWu56p9lGzQP4M+u1Nr8cawEVvsZoR2DD2
QMHCFwUHqzJOgsE9t/IJXT2w5FI0Sni7qeU9thmX/2CZGBcZVUrb+jwhQ9x7
h+m1j7AEHrZcdlfJv9iBc2Rs5QeAFnYA3lmd0aHY2p8Ez+Jok7qmLEPC7XD4
JyoKC4Kfp2gMEjMyNLd18pLPzmcJ0iBJ1YOOr3asqHn7lh5Jirn6LruNcbP2
eIw=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpeiQ0L3KZLcBbuRTe7VqDKMA3fnqiCSqE+1t7eBZ2A0wnxqVWlzta4wq2HG1nEifAKBfTlzycAV4JppeFCZ7Y6R01Y66XHXCtt7AcadXUASSo6EDSN3C8vte33uFNI5IlGLpk5+ND4FmUBbEWFuenJgJP/NITv1o629TQyWZ6v1qlBOUpynw19B7uyOyUS8O4k/2rlZS9saQtcxG3gQ7j1nxnx51fvGjzB1tWNPH+5D2Lg0cD5a84aYSnkW9YiFvJkALr/jOavkCwni78SY2N9Km81CPnsHaNUz+dHNGhry1+BUGCy1GEwaHVMcFPJA28IQI7QRPF+IwS+8JjdvaCxvBPQdSPfz8eKnqDz7GO6HwOc5rkXvYrbDFWGaCzScDJUtpV20wx658LFspbsB8ZC5cVRw5ADRg6Szlqz1vc0+IM4ksNpG9TreqpoEQ9PdbyoahIeilcWmjWOn98kOuGxK/Js8RGAr+YecPpqBxW+BQYLCxsUIS1t7acb14HkYQUQLv3zZWWQgWMSIskAjXfP279dh1qymfTR9lhWmtzVRjgc3OA4tqawOxAvKApkMRRYIO8Xfa8JMzEw2sm/TiHVEYZQZl8qDUKuGLPFExQIhSOatCzXdg3N1iV8P04mQdiYyM+2DrU2HuXIsxgwGMVpqZhiuLXByZM4T/iPqfH9VX63YQPmrOa+Of6/p0ikNOdAAuKoyYYS9Sw6yCmutRDjjlcBDs2FuPgdb6jd9SM449rZniDsPJk7EDiMADAv4v+TolPKs8zZoWyc3LvikVzzte"
`endif