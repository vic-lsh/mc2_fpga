// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UxR7DrbZzCqqAO2dg2p2xxtyJ8TnmbhTfJNlWO/6MgBH2YLEy2ZlZ7TAIzXw
MNXPVGpBVAMlIchnjfXpT+ZNxJgJmb6RonYupNjG3Y7eij4xkQtu1bvqhkSO
mauvLf66yGCFxDYKG1YsVt3/H0eDPQGZVbKe2h2Ozy7avycnnGLgcnCxykgd
6CKviRyxgk6+3WfLf0HJtRBHwtaDiKdEtGfqJbU54DT5ARNdfQX4Ss2RSDi6
KU2HVFlw2jjFpmA4Yzh2Cc9b/4/vMgQ7ECYCI+fmWufKvgaIT2wHo+ZySKh8
psKgGz9xbtTyu0Nu4ik1sJkaOuZSq50OUv7P/I1XEg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
frEabpr1fRc+Gbc0tcse+tdDaIglrB7FRMZ6+8XzMeV8jMo/sAJbkR0oYM7l
QHscJdrEi9nFcxnQgcSOmgajiW89cFt1JzZD52y/TpqXMX0XGtZCm9Lxe2SH
IbryVW/BiyQULsQgG6GwO9hXZxxJAyFLfD6pkczaeTFrhzYqrEvw/xW4tOkA
BJHKW/bosTBXVvnuSUKfuRkGtjJ1xHvim0IKXz0LqS3jYc0dti+kJz9zysiJ
djD/VfakPfXHo9SSv9FzTgKN28YCybCShP4wJhJAIlxEE1B1lObbD5WudvL8
RpfPWz6ChPLlBsdwprpK8jqcgwRk8FqpymsnOkF+ag==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AMMTxyRU01waeojlJlXIYkCoQ+6Xh1+uhe75z/OpchXtgF8lvHeivcvk5mCl
dTCLY+WyPul8dQJSMdf7/kmfSgT5E+ctj9AneOUZ8D97Q0z3tRUUWwTPxkGf
TSuraCBf3lkr9wpreb/lYsugLZRRtKURzCCFJza+9qtUCxFuyaiEMKIMseSr
bHGjB1THis+X/g7pge0ntf6Mh+y/0Z3KRPyHAFkg2ch5nfTF8COKdp7viatS
KJR/OJ2TEsJw5AOlwIKsvMulGDGFEiQ7mCGNWrv8zOA/IuWvMEx8zgtHFw7c
Xu8A3t6SD21pLFNT1AF5clTR1zCKXM2VkXeMztDQQA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oz/OM/0tw87UHXR4B8Mcxb91O5O5RzPavhN6cfSAjrv8cqYb+TxWKashqMYZ
tyyMi2XaWdDHJ+DDH8atZSUbc14RWrybR8eixV6xDPJV1Mnzi78rhiiaH2Gf
4mfr4XABP+qXnJvbjJRV8Oeg9T9YuWr4Ox9rw89C3RYDfhL6vmvhTfDOrhXy
iW1RqnnIOwwwU/MUsIqXzvbOnwjLxd/27OEf5hIdnV7iOGQhkAtmdTTs8a2U
27k3k4UTC/RxuuXi+Wz85sYtG1GDOd8OQprxwru+kCs+FbKWWIU5hkie8Hwt
sADbG4nld5bX03Q3f26mbvYAvvLltYgwz0S0f7MymA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lhxL+DHNAtOnOn1rXlnCQ8ZQWXKqjkmvSYya0AtUV0YhXv5NOaxDkU2iTWcm
GZIzPfzABRIL7TxVdT7GlcAzCa3jQYTER61gOVxGEujkucJs2YiFlo6sSOTn
5OYcSxwjY3NP7DcwaPryg0JLfjbbe+bQF2L+BbfGAN/Y/+loFA4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
OIR0JK3Kde05/Av9ENhSb50LeuUeTWg8E/Z8ohKsfKgJenyrxFzVVyCMZosT
QsIrsqfPyRXujHEjJRHPWJKXUd+kG4Bvy52QowUeWs1Sk483aBHMbtGXhnM/
hBSDhPJj+PWsCIZFxD76g7mhTLWh7kTW3JCkp5OkBfCvvBwkgJrKPXBez84U
r8dKLKFbl47UTKRxq1vy4ySNMYT3y4QLTjda3Pe4Dxh1gsJu160FJIxk6KCT
jzldhqisUCnyz+yFctb8lFAJTrOROqBoIbzgiSNIpgXs2q2mQGKM8njz5YTM
/ZsAI3N+5wa7jQrjx7sR3co4tgCmAoI4UsNKbw6vlG6aUDeeomWQLFHFDwtE
aF0jHVYnQFy56usxfaWvAmnEVwzOrNPhe5MjcPwHEPgxeqRWtjnqKLJBDkdD
dtI3bRtAH6Vqi/tNJbI0F5EV0QnDE8LZciSCqqEeI/rRuW2Ant5zUd+3FrOv
1T3cI7qPg+TG8IBVopKNDoxhTUNmP1l0


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
upuJ8mjYLVp4xfrGXS4rUJvWiRauP7qdgMVGUTblNhSxhLNEsFlkypZ1CsRJ
cQHgMC+5z9lyhamHtKZLQV3iqALWpUHIGfhrLJAT5U4wUDtYGjGM9dsm0Uc5
xS16m3y3AfTm0gnnSaPwlu8dkIW99fQhpMCr2+YyzLkdhLkeAsg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kzsUGjUljQkwLRJzby2f6e7wgzr74KdreDLxgJmZTS0t/jzM7ufcbPdx7U4R
kf0MCtLjLkY1Q3Bv00a9nFApVcWF8wisWQCITl8zdLFMbRullaI3jg43At59
H7ujK61BPqiF/orXN4aSQp9OzDzn+MNrD5AwGh9Ti+aTwHT0NpA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 34800)
`pragma protect data_block
jDWQp90u7Ecpyxy2+jna65VUW7j+3jydiO/GL65lWTwl/lciuMuGf6/wbAIn
UjrERrgUxjl4kNskDXIRaPPyynod3HTpg5sf6VEHJ4feiLvtnqovKRh5hQoP
I5TyTGyzAYYW1WS9di6Rn6AXL4ihgoa4/ysnKIkfutLm4Wxn18X/vfWEHpS6
cz5P/522xXCUHhzWEf5m46tXb/w+U0XXXBUtVxvjjWFAsKUknMkcMC9SJXL0
nnjGm/tPNlugrKbkBAVsOLvT7nfg/IJpp36/VnF1dNJGAZhc2nA8kXKc8g5b
GckUk9Lq9CsXFD/daVr0JLicNs5VmHrIGQOvGeK4yLVZ/8N4+oOsr1D/bcT1
gEEE+l+uQQjZCVkgFybZXM1cISSv2fa7/3FUONHXWPUnACaFZ3KM/yjqUH3f
kQ9waTPmJgiLYrBYevqwWvQdA5jrXuo97YIabRZeDru4zhQNkDInJMGU0QoX
47ECeLlpRrp7yDsu28MG1GlywUT9fA1Fu7+NAzI7TyonQKVnexlL1Fm6A3Is
Aeskjum55C17HTusMaLCbGkdfUAEoSBkJqeBpZT+Z5s5EcRZtI9sH/QJ3jeT
5HUjEjrtik25nS7FCesF362973ncMnLfiJx8e0vORe130A3fPw/bmZSa6CN4
bu2SFhTsNlrS+xY2fGk+MSlB2ahUfAhHbS6vpAvz/+67ueP5zX384axpPmQX
iPCCeeFMN4BOGm9qte/CdvuzEZK/wktqQ45uqR2y3KzXRZD5/kHj0brLtRq5
f3Xgts9pDv0Sz3k6kuC+yEC87tDlbCxjPE9psOWeWXV5oCjtUGrIZczIHOkV
Fo7AfVeKD5uEAWDRRSlYqrbkHovYwsfStMUwyg9ujwtXbjwgKYN4dpxacv9z
k5KMYvZOZAjY+Zp9wZSZNltqJLjxE88O7AfZCTmiYCNpQmgBk2hRQBcCx+Ge
5At05iubwjZTldLvAvl8jQpwUMtZdcqJGYgfVMAWVMx0om7QaZPzdC8gQcAY
cWfg4R7BFg6YNiw+37b+AlODUHvh5vYx9FnyjQGzcyk4IRYstU6FqiVdW7ux
gacVJjXe255VQomPQOYGG9eeltjUKKF6AEW3PCD0cEgYyZXgQwaFvqqylTq6
4n3CbI0lOuw/bAwZMrHHjH2GfRCwKel1hAEE4eH+oEjk5qQnIlXQR3VXbiIv
HEvrAeLNKWBnvrGhGmcPbQlr4hfCM/qwl3Vq8lrYoCBnK0iSUUyU1ODQSgmc
jX8GnbIsbLypaSNHNYTBH4L3qqviYdae072Se19HlYdqyV2nH/XIfaBLzOAv
AcHcz4Pu4xfRkV3+R8Hq6NzBN3lew6fURrSKZhNtUz+fsbLtUiapDsU8BuhW
aeEwomLHKi6uC+viaPkfNK+RCCIAZTBRPSxyN9wXsZGwKiLlaMRrX53n7v8N
IaWftvIF9ODp5XIfyFzlm0dCvaGpSbG5HSbcFpU1mu74wheUQkMoodSMljfw
q8j/4nWqVJg+5ldSxlaTyJfEKJv76nCGT0nbivtMfnL3XLwkAdptgARe2Elg
38GeRBlQqEleglfqgMmhC7BdYbeBoxd1h1O9x8DDW2/w9cdt2mQYlIdOizHw
4IIPsUNyOR6XF1u3LNP9DYkB8wCaN6j4pRljWZYdgiJyQo4aWiqV47lRUD7+
dzUzKNKNsltl+pVSte5vNrHyiLhepPaF9m3C2Q0dq2pKvuF0ejaPvx87SZxS
iGJD5WotpWDaGHQpmUMje28O+85ebd3aT4IxClg9h8ZB84L5xAZCpK4FhfZP
ADojrrHXBHH90dqpF5iCaPsY3LlfdNG5AfKLGNwYVrniH9u3KS5NqcE4noiT
kUXw6j8435qDlGRCe0FI7A1OhJZKJSvU0nOWtqcLGCkdadL06qJ0J9w+Sret
SYexNLmQaGmYwaBcNpL/bpbKyxCPwbj86KNsVJo5hlMnKkTQ2ldxonqXoaOg
MI92m9mrfiybWV+eKURj0Eoi4uwA0nLPfo7HI2AEmwdMWEhG72rM5Dt9pQ66
3pB1KKbXu95vx4ymY8iuLfwxfrkNZdJpf332xerWnqiUSq9BHiC2mj9UO1U9
aVlUC1olRhiOIZBcPEXdaiajtmuO8EKOsNcTxKZlg98q/0Oe6A6+3/0rBXSa
UI3q4glg9axtlD7pnhZIX3eqeFyPvb0cinjTC07l+Q+FCbcw1nk1KpkToVBZ
OQ8UdwQXOcotPIYJEWP9jWdXZrU7YXqNGS3j8Wj/Feu6SuwGRIZTgJ3cyjWB
fUZBbM4kfJlCWPcUg5rFWPiNVeutwXWtopUlnSAyi9ZRz/I0CQR3Itkuzqsk
NOg/UGGYr08LZSArAV3pt/X+0Ry9/kDCqGRjXHpQ5CRfgDyDiXjXOzChRxaf
n82S68nmP9P6yb8hb/+7X0B2TStPjxmZjE1KrXTsBWQW5EnActU+TqFmSijn
SEpWL6oc5OlbjmaoIeLGc+advOQE3nCJOUUUfovS7AGgwLA0n6F5iEeApcIs
gmX2EfLxhQ7syg1C+rAEZIWpCCa1gbvsEWme2/9PLMiCnUVi0BqBkPDKlLWN
SjxFTUGazOk5wbhM8t9SHOQ0DNWxSy3W/91jShqqe6rWcULYbYkb5sDnMI8+
RLqL5mzx93prjmk3oCi64rCEo2NPNR3SuVc/EydvG3haqOZkrYR+VfvaRefI
SvY7gHW244Zyydpa3COu3u5NoBCCVxZMqj80iNBBIHmPyulo4kYXRI89rzvN
nY0DA6KDh4YL+CeUpBHIb96WkILyEWrMP9e/gQAeITwxKP5zhcnxW92RhZBa
iDknu5ENbEtFdassSvehMRyJwtZYS86u5NqMWOcXT1Tpz15E8YnW48rBOIld
rtCaOKCCkh3bSFoLYZz8bvurr52617eNQ+v8I2bkSfEoTLWT2ZQAHRms9Nq/
i5Ii9qrTPrcAd5G8Pv5D879bfOGJwWIk24gArjRydyuSiz+uXk4xMBvQ3let
og3eeTMOwwT1GqQ2Fr+2jz4UygA7kGzwGZkX6EvvNZ7QGDmgCf5urj5qJl4u
OPjTkXQEK1UzDts3yGM5/2GLniU6r+3c6JIMAaTvmNZgKu/JwtW3n/Si3Eme
HwAgjhqPZZagSyFL0DQKQf5aFUjfShEgr0gKT0d0UDtBLcHj+XK12ZD1ZmG4
AiUqEc+ynjKeWQEtXpnGNn9ATHq65C4dKePGQfBkoX/bAMdCPRK07DKTNk+s
kp5DuvcHB41RtMB/5kp7wEcWJ+c5CIoCRogpyfN8lnaL3zYVoXZWv2Z54pna
7JF04YI+C83y3dum1MVsyP/Zu43TXq0AVOTSileYnhsyQv+j0WhPYFQeLf79
kqYFA4WbpmiWMpnB4Ws9YUOsWr9S9xHC6NJ3zsiIUREe7laLHfqxS2vyd2mh
lWKcs+87HT5XB+ukTQ6PiHVrQe1+hwiDFtg+SH/O8CQToY9JBa8AW6k33JhI
esZc456xhKmWyp8uD3aohKzGITshi5ddbepv7HydGbph/2bW3oBZsWMzSuaG
3DlMtg+1/1n4wtx1AbSNo4YRqWx6sWaRqpzF4kLrRER1pyOxSFubVKVDKqlQ
XqX0+VpUEnjVPdI2PJmPbSKrXwBoLwMjmbyUffsOE0F3p33KSauK2EJfuTV4
PFcE4lxyFcAdpv8zO4yh1WV82o1RPRz9OsL78F56ZxtuF6exk86Dc+WrjyY9
o1gVrjxdurr0bYSBoRnKgUd2q3PmZxvdk7uCmlsJg/IXAVB+X6noUlxBlE+D
ASouB0YSs5AOt7LNEynZxgnO0DP9Ivtk7rvbk05TBmrf16zfi1bLLJPmYB+F
cIHLmeUUJ8ytRrug8TTpp0MVTgNyuim+S42VBres5h0Op2AyQGyby4nm31cO
lnrf8fsPeFzn33N2eOU3bp/QxAaENLWwl4mlnEFfl8rHQIg+cICSE/8y3lFN
ZTNwYztVpPGmJlzAlniJ+KJu1GnIQoyZhndiiS98s3FPsh6Frx939daygOaL
3Sr0/9lJmQQeMAYAPDy4q1TQr/0CDdAZ09Dn1gYw091AArQv+udWNMCggrSi
41/UrEoTVAaE8vJ4Sxo82xI0dUrBCaJnxlHG5wQHglQeONuIvlwJedB9ZZu5
pszakrmsqK1cVQ1tFZw55D5vnSXat6X/tg+huHFglBFNtsE79p9U9HpuDNLa
5msGep1urqVsqphGrqUAGjtl8RhEvH0VWF4sMgOQDvPcxV5bfdPKEhAi2Gxx
5Ky/pDYWNzdzlMLFpdrdaSurxbY/DJILHmFq2gU+mOIuztbYVVX5Smx7OsKW
forba0zHpTT3nvo9nBi7H8OZGAIv03PB/GCV7TDctjQdsYrrV/qb/eYS08Lg
fyYI1oToGGa1tPJJBgmckpE2y4/9Zo4JvL8DIyCxyeKTfaeBR7jsPO1/bKyw
FE+zTp7aTWwTr26Usk57HaoppcGGPj8LDy5LEY3zQh+tDpn0p3iXUMFvTthO
JIgxl9UTiysfTIoHeCMCdRZ5TE5+Dd59F10GqPXryEzFjtf1yeyWLk47zT03
yKRtOPxSIE6/+HMgvxLjqwsqchr4i2CbYORgpj1Vce7zdWM4pCwJ2AeoYgZ2
S6Q28VGqJhUPpffEojI5ytpo0j+e7rbaSaCoZZ1bz/hEdIPAcxYIuoq2+Pia
0oXQJ32ndn+KNARdeiuOKYtcIW1wffISnKkOBM73AZbHenBfNylUpUY6vD5d
ZSPWR1ev3Wi2fxE9gSgu88XeVy0eJOvc3grTfpkEytdBmGi6paOSQhxOgL/3
Qy4v81xpGAWgrVrUWs2NlQ0DJDcSnovgqaRaKTcu9G1slh7lNxoKUHHWFkdu
Nq8BWSYtOcntMyr68VeDQS8d/xSm1LG6xsZU/KL7GEiVmeBs1XNkBi2EC4JT
icEo6mT1KwmZXICrE1GHJU9a4FHTryTm5WzdaRFKXRAZpKzZKDKrZa3oDx26
XrKa/m/iwELnrzgehBfYslT/Rdtc961HV5uM0e2gzf4029ZYd/0KyvvoBYlO
r4y+tKeb5dgeHz/VWAlzb8q44Eq2QZ/3j7YfWV41BQ/034AS7fVHyzRB47R9
9hFCyjTeLLeSSLkCArwioiEmuJCf4D3vjANrtvojTlH00wx3bVESny1Z5+mS
flIQftrDcZFM5+V+CnKCdQRqPrB3VVGYTkpjjzDmOPqztykmSFaNKh19MHoi
PWvdfsEEAMd++OGpHbVRhkxlhm7xIe1MeGvXkTJGTVrHslkk6AnpZ7YO+YPg
pe8smTHCTmardEBF7i9BGggVtRqCE8I5xa8tLA2D1WDvM651DYDJ7lexoRtK
QgyghgZ2LTzOJxRrcUVqYGvBqh515g+cYgD6apdbv2xL0Ud5P5upFPj4E3r5
64um2KxfX8ya8fU4FIQTk+PGNtf9t9KIuNXG0vfp7SFp2+EsA+JJbx7zX1Dw
NwXu87hI9Tpu+GIMh9MSTxo7VOtQQNxkpImirZTlxZeAPelx5lE/9BcHPuNs
9QDEF021mPRL+/MPAbKGgADNZCXu4PDnDcLuHwcBywJUB2sfcyTKEUpaqZY7
f27XggPLgNBEnGVywojyKVz26rJMAXWb6pixbEp5LWTsGyXxExpywbbKxDXq
AYQ0PVa8I5PobINja9/a8XvEh3ncPVg0ja1TQWo7MND2OO1bGRx2NZYoWKiq
BNO0NXNhxOv6Qq9tUUtJpzWk1vaeV8A6WroWau3H+uoRUcq5Op9ndawEQTea
lIeHlIZtc3CFjlKoG2tBuo1kOnneg29Nxlv2EioME2kEJOheMZwSS+H9zYaX
8EM8fPPCBruvR0fRf661Knp7tp+JU2QQZDVvdqueMcOC5et4xyWlgawdgVPF
7VODj80RjOYLECicbH18Gj8x73aP/AOlXYfiIwVQSqtqPEbw2DMqeGG5rLI1
52oA6c9hDoCwMUL3Yx7vI4sZ7wCQjqx0eYO43Zn2nipcO0zJIoP7L/U1mNfa
ZENNt6FdSEeMC4yClFCO+Cv8G0WX9CZNZFNCDaGxbVfHZdE6g7u34+FpT9yd
hhlk7ZSRrphH0FgkT0UZZwU7YPSNL5ofCIC5RDRa/xzKC70WhR6QOTzhLFry
Ex7Cv1pM9s/f7lTgcCaehnvKMkfrzWhxecslv6MU+rmKBJKPLRax5dqR/jMc
bZOZvDPRXfpQvTcMbA24e7r67UEtj0i9m98D6zP6VmkU3ko4HH8m5JpJDq0I
8fRmfrGkqw/Z8KUEf4i3odgctE3EibbtbpKAyhEzd3VU7Flz3+yYHqzlIFky
rbLOUkWa+fbELKVs4lIH1hlU0vGZtZEq4FBgPOUuUrM+akB0S8h5Kyrksa9I
h7ezZ8H5IMbrfUjpnCa01F5WTWPv9jhsgBojdP0kyzyTRvZjqafNvOPjxTj9
l2z+DbZwUwG2jSSTutD5JB9AD9qkHSFw1+NmVFAAdGvOuTRlgm01s9T84Vbe
iZTKjDYC9KWbNIEXP71abx+kmim3j2i3nedTJIbZbnzqDIRjqgh9eUlVJqKw
1WZH5t2ALAfW1B0JaZgY1wyRXpiCw9udMh8s/BhwpoeDOV4VUD7R+T9lmqa+
pvCgX2cDS9HglVb8kJO64h/1Vl+kJBJ5ijlbskLKcSCUA2w27k1DeQ+szdSH
9C+yl4R6s//JVDmBDG6sSZ1YFnN8xMuNwUssN8OaVuhAr+w9aIMELQJJEkYc
7akdbmm3mISmqzkBtJ6U3WbV2VZPc1TA/ebq1mUrNthHjK3dNxyI2DfmAaRl
WzJeWEyME25II4fzkrHB3YcDtF2axWCk+LIPtjivOYH9Spa1+M/e1s5kvson
bZUlciEo6uGgwbr7k/ixpw1sfHZXBsm1Gfmtx082UCm3QZFyhmmvf3Nk4DT3
IdM6epta6DN+rlHlMdUrgbd+GK9A4pZ+M3JpsEgHjh8hUuymxHE7KbZr0ApV
/ddQ1mJLnEyKjBAn3428cQSn6FTuAOVlxPKClsUArvn97mfR/FMZ1FsmfS9s
vb+QdLqw2+Y7iRmRsiCQ9JGv+dw+/MiTNPOU3HHW4M885i7WI2ZBNv3CCOLg
sofe6CP0jkTRNmrvXxdL55ZyMtyz3tq5Nwydu2mASqVuql3TPRMBigY1bjs+
heh4un77kOl+IHTu3CTqjzyLHnxDDgC93P2oRiAzKXbeB+Ftgn1GxLWmnPBt
RBFmNcSvtsCylX1eLGk/aVGTdrxyxOQ4BypHr5GbWSRaG9UlvwflA9nB9wq9
tvuhm28FtWljLEj6eYwuBzriYcHKBsJABrUGF4wH4uJV4Y8pic9x4La3OTDI
uAbeB6DW6MB6o3BXrMMnMhJab3Bs2tAm0qTpoXhFWslcD0dWTQQQ1n+u4ZL6
LoNIuY9pDLbtEhhZiEl/u6dZD5zRJ9yGjditPOjCXKCheJ4hTFYjnlhnOHdr
rKtHn7Tih1DKMFSyRyclwVILMyLy6QJgyvuJCmywZxscTfz2V1bUa8HnDn3/
iaPf/pp4xGjXe5bjM3dHDupBncMJfxWDMPcdzX43bRsmDPmwVLa+VAebl0Xf
8+gjdOh5uHcnrpRef71ESxNhJM5/ffNnC0MWgMAVp1+bFRnFPWXS2XqBTKau
64mUx5VRhMCy0xHwi/Ekklb2coC/u1NL1H/xA4Kk76qqQtZ45UbANBbAzwdU
IhH0JcK4hhUTVLVgAmQXgNaQezIJ2cOHz9zdPcJNP5t6L152P/JhTapu52uG
/I2ppA7NNuyG2bOGOKD2cOddVFQ986x4DQ05ImYOikQd8zgR0Rw6+Pc+U8G3
uRz5ombfHQqxBr+McpF3/UdDD64cQAhMSr1vyxox/EB/fzaLus6kpXOkjslu
13lM25wo0OPOKe9bM8lzME4RUGPhFvE4YMGKZZkL7D+i6YZJ/i1oIkYwvQPI
dSALSxIuJsZRNLOOzHjo4271B9BkMU2VhvWgmzo40kqq6LtU97w3wHrduvDD
mv65bmX/cqvC+ZbZaW3oUGolNyzaNWJBqLUL5uOUjHKgYnUjaQjAD8fFcWdL
7B/6og2yYLO/dS/6H8ROZiQrca24hPCyF7EW+t5YutUC/vMI704MIXjqVQMK
1hS+dEhBL90L1F50ePP64CCWKaHqOB+X6hh07EE2PtoFFR6cb3QuWCaqjO9C
fGbjhqd37gANfzHrHWTNPGNNZ886nva33/0OalPyOFdovswtfPeQ4vk+go4v
0Q3QWyITn52/wXGL+gLMrVVYkFeUoMCYHa31+tH2HqgbidsyTo76SJP/08rd
khEV3Eknw+UPF64QpVk5i0G1VwkRg9AxPRxwiv/LbnhZyduXQGWbKtzsnjqh
oAtQcR9exKDoghTunuy8vcoWJED5NKmDYaINARgLHuvNSccXn+l1LvMfFMiJ
ZmdssgzpXsZnvW3qWkBEluvPTzuPlkifwPfucQWAdCDlNXnsSrK/BpjK0mon
rejjeg7fU/M18PVao7dyQLszGNaV8/oikGYM+VEBuhLQGHrt1eWSdOeFt9CF
3I4KIyzI0YqBLVES+HSaoR816JkjCm4I4DEfq5CG86du30froNb3i47+o+Z5
vaVPb+UkXoZX3cNu1yEfP/WWnwY6doW22xnedZRKPymqw4+NBiHd82yoPMIL
hO0KKk9jKZjKEslSSmtbBPlKKF18hP+aT1C07AK+97NKcTvb86/62vmgeTgl
ytL4EIH36TL/PSXYT4HHQANsuW5i/jpR16EYsjl3SN3FPbClJpi0qEYX6VKs
18ijYW/v1ubfH/RVmCAjOuoAMO3u++zuMcnRQX2ND7gZ7UPa+/D7B05tz30A
xCzYWZ9+yoU8jnNSPbgEQ8iN7L0f+NCfTzamQLkHQ1oq1tG61pHjKSKbEE4U
zpjKxXjpupMjJXf2i6LThsgMFn5KD3JiD6iW/j0mTX/wBaUyXAf3Ch0xuKGm
NvTXB6+bDalUQMP39eLW+GT2xX3KSDNve4YyyZsGoxgqpNAUMBpA9MHjfpDu
vb9T5MQ4/Uw4JrhwosaAv8Xe5t/1bJTLwp6fgIlG6ChsZUqI9kZhp5VqsKZn
lipF9k2f/Bi4UskbWBBNoGORDXGu89VO2pAmoz1krXe/oSBWBH94e8hgSwd+
fxXDryk6jqWAmHh2TGdQDBV2oXc/Ee9vWsRyoklniSnF2Wl0j+2RCXBx7dhO
gnFBb7t12KhqbFXg9u+yg52Jr+h4WAttPAyrJALCG+wYNvalc4ORsnHOWWjL
7+e3YZ9zJSFyD1UXhwa9DuD1LBGnITV9LicWuYqzi6RcVAfHejQYC0HhLGe3
gMGjBKezvfmmHIAOPxsXsNqPqcrTFJq+llvckuYaaNd3o6NA49BYv35L/59C
lSLcFeje5aVVLfzEOHXV0m7+whaMUWCA/A5usp/nzSb9eCtOeLJ0WqLBKWmo
/XRvBXMCLuamAUXSZKwwndg1+PQz255oCRlst1TflVTrz1R7NA++brXKWyyT
q3Wo+aqZo6Kwt7y0RaqkKtqQNmv85bFBxeybqT6DIxx4le0BIChDUbuKJcFq
Fqq9O0aQxOB2W5IWm0Gbmhr/P6C+nAHIgWyTaP1Kyt71d7nW/U+KoG2GCi0B
hftXjjqj/pRWc9II+iYNxdclaR2yWaIcgT0ZGbWeabg1lWZ/ZTgCg0F+Jd+L
TlezZkZYGsvvXFIZKhbDDhA8lAmFbptIL6qPTHdD/pitQbK/OvLfDzqM+8cy
VUA0MNAGu3MnqJTWs7/S+OC5BZQoO+CTTJ4T1uDqipYHmCg+s+LHw5vV9HgE
W4Ib1BEyCkfmzzKERt4KcNS2cmGsqJ9qMPc80BT+mAv6X/q9ZX2oY9KA9GUM
XeQXCc2fSx4xuAi52k8QVA7jI90zqbLqUVQUz0/8Ju82yBqObJfNqjHpzVPB
Q49eRfFDldJutAMpLTJr9t4qXzQxeLDhyrNmPwLwV43YtJPjrCY+w1lBfwdd
Fa70DHJoyBo69LjootcpZEB2QUKZE9mPxGOL9yd8+xrwn/tGD2yh0uLSLNOY
emCFvGetRZjXltN9aQD+XrKXCckxOBkWpLWeUD3oLzJnudqEU6wVKDUbDcMp
ud/oI2XTxlXrlu/J64/jBkdUNNmV+pKJ98g4cr1kJvlcfeoQqXfPC7be0O+k
sIPgFQkQJcnKHi5PimSjFxiqmPbxFJs8dGZNdWcfe0PTUKbT19Xzexrfg7eE
+Ot+MXW1gBFIm2u5xblHsv/Ch+LD6uesj6rHK/5LB687YygFW6sVvRLbvPet
+zd8PSKwea2LfYRlcDxvWkktTEfoguqb1IgShCnuC6D7eehiie2N2vPGZ2xv
VihZTMIsAi9fK7uQhsxyQgZijSQMOl2gPI841IqAO6jV1bc9ELU+kLiiYK4n
+02M/v5D3u9nX0DCfpJ/X/Z1NrSdBOXdgM31INa9JpnkI7Ys/amew043p8BS
sxwyReHWuJeJIwRWDJ9BjsLXin6q8kU32DKFtd22l/D8BYGGjDW6rYkLYuO4
P4TR2M3l8800eeJWPfXq4J8o2tJrCkdViAIDuVy48c3lyBBtuDp21ZCyZpI+
5qgMdHvZc09oGCJXPZZGZswALI2pE8r2HS3EI6wnMu0+yLdVYeSbk6+ZCUjK
/YHLoUOrwJprKBetuHLSeInaMakZwQgg78/3yINnE8om55UtqzUfiZAER4EG
YW0X05DKV1NONhi4ZH/fU+01sNU5VPpWLKFDXobGKgwddFVBGYP+WrZ2aftB
Zaca7dulrkNw6z82pBMsgXGVm/3lbUf2BCd29nMVuljkrphjtUYWo+aMyQaY
/ICC8MWdJRAHyF6aPOY0JAhHU7FJ3deXI/dGhYkGo0Q0HlhFPjWDowqoEURH
wT8oQSXU9hnzI0IPof8EzQV411wen1tyaYVkK5hILit/uRGzEMT0HmOvnf1l
DmG2mR8CA+aYLECOEKfjsA/VGl+4hgzPTTa5WCr6XDOEfRIFcCH5KWMaBI2q
40p48OJNDbJbS6j0RP5GoA3ke6xl1Un7WOMpI32qf/CKxHyjnIRs+hZQ9ITY
WKPpiJIvWgrRXsx4ZV98i3ZKk+AxHuCn/u+taG7+dPeeFDZT8DDHZRYo6r1/
PlXxIIj0ju8oU9X2R0yDfZi+EgTVfd39BJaL5PYE3SygRmtKplkRcIcjTmmX
J8KO7GmMd/+WsPChUUMgWwK3dZiQExBmQsgvLHdI/vKdFVHRo2MjMLpaW00v
GpCNYHDSe9hpvxq6Zjgi/C3Nt79RoyYQHRONc8FFW7vYq1SZirA7kNzlqaih
K5510A1t7QLb55ondZGvyUF7DtSZV+NjX5q22cJm+sR6yFCgJdntSuYrBXPg
bu1wxMCYCi/k9wVKF7t4JnyKpz8IoPDiMymPJHpuDFYeu13ZftyDsKV45TaD
CnMFdgTY3WK139SRG7G5gDsmd7PD+Xno12XF2zWJtf/ZJk9PEzpxRU04h18n
9sOxlpzog13i7K36QnK2GEcNf6e45jiomeo9D8UhPB0h2n2EwELL/eLqUWFd
HyRnWXcj8p3mO7C+meFlgZo178i/qjvgbuu+gc6LjQjXttmzh5ZdRRQVLoJf
kpUwb0eHWj87zx/e7WeQTw5RtvK3PSXPGpK2BHSLrdY5be6+09lA3sTtpZpk
rUc84jWB2q8Mi5cqSSUEMfG2WY/YcE38B7CXwLPmlA0rKXnpiTa4fYaI1NyY
oyeXaZYMsas3jkOM2YFD7ZS++HpeWAE/uHtKTzPaCRXQlteaeg8sLaAZ7h8d
wLhuAVvSZno7kqGWpaOOgXHwko0BgLdSDAzez34KKObKA8t1+coQtiPjJflz
q8GmsxrtCHXllCvQhcvRZC5S16AtqPI9LMZbDeCu4COn8NZa6jTDnsXZ7Fn0
4kFMxSdEMk0xILds/CGpOWtcfIGYuKp642MMDgx5iuwe+yTFPlp1XBGJYjN+
afhL7qqduaH8Smq9Kj2xATMzLk1X34c701H10AbOmm64/92MYjbuJsHWBljN
uhWZp4NhjFHV51urJo0cSu3PxsJC1E+rOsy9glMoTfzNQKT3+tHzgmgj0ts4
PypVaBS82498tUGmeQW9MBkwpPpVU/9m2oPCNRo3kOO1o8Z66HdtoSg/Rm03
/fhuM0RhnJ6tgdPCUacm3ZqfZxaLL5BTn68xu45QMqfz+TwIBo4ErmC7HIr2
qAbI457kbWFzn1yQsfpH6eksAJ4Jzs/9wo1QLN/Stttztr5anE2I4ZmCjHT0
zB5qelXXS/VB1ymtPsoG1Qd2BO0wRnEZctT76vqglvxf2DluG95fL5IYzedg
fSDXYflrNOJnNV9p4cWGzDnYZrfm65O4QD43M5aH70BuTUHvngTr7Hh0cQSK
j1fSXQbngtJX1E0NkeoQtBERyz0sEMNEK6EnBzoyhRNqZFHxxDjXSPQOO7+A
1NYrrFM8UDWzOq/xxAbf7uvFwxZ2DlrXC9YjMgbf1wnMEGZdfcGPpUPUjOM6
DB1mFAgisiCltxjNenGDQX2f3V8+swl53vy7AOMeEzKlwaVNAAjBqtZTlmhj
MBcn9UPv/2dNd+2109yoyIAN5Dua7jzSVTcxeSW2/evziigg0a8rTgrBtqSy
PyJAKkzG0sH8738QtoXmXIrHdR5a3nc814QVDD4BPrj8GXO451aac9jCA/LC
yKoiumyHytYxqfXGRjQGL/oWHfzYW+smxKgKnfGWPPN2tD+2vlNvYqRTssVP
ngzQxZZHj/l5EyWGiqEhSO0waz5aW2hFDLxFuIlz7fMVBYPXEHTqfoRfgO/5
o4ko15s/icqY9MGJ0SYHz7rkFIrN34+JvYsx3q6Zmmvco9Yv0gpR0lxjIGbv
4BJlFYGbri7sh3eMjWQ/ODyCYUmxIMuXc/HE6pmqMg8k39OhSqtF060x5Jp3
QlUajwYdZk6CrcJ0eGelBnFZzHd+F21IuiG9ZNwJelG6n8I3up1gNAYUrI+J
SKc7W3tXrrJGptlUvG9yBpU4/CwuEdGHAchlczUzBNcxhPX2FoIsoSTJxC49
KbR1BPsCtkHW+TVW7KqLAG/AeSTwiue8t8IAsABHRX8y94k7sQvDDbbncIIm
HizC25bj2wtVBk6ZX5fwwlwncE+IuxVUr7gJX9afLofUAufZCHhxYrl/F3O7
6+81nuNRVGr6Buhqs6cELnacIYHF3Isl5CPJTxTzty97Yte8CnBkEzGfyqZG
5HNiV1urd6WcLNwnhOfJwxnCaScYPyj0BChiira6IwbufyB1h7YlhzfnjiM2
jO1l/Qb8QKzQSUeGRIBuJZG39ml1FKPu4+iKNrSKue8nETElE4WWeHlq4MGW
SJkk7jCSPDZb9M9A5gGGe2BcWJeLNxpD43n7I4yrDTjaqJhOoV2YBK06/LRM
BeSfbI/BRn939zWY77FsyV7KrQEsR8f1OQ0Bg0ycIQM8Y1B4tFaEwjxXEfHG
Tx0WDb09/qcQnpZCLjyxrmNRWPFP8eLR2voF2KET+F/UM68/4gB5hytzI61a
knsneQjMcIFB6IhNYRfF6rAa27oCc1w3IaqcncrqAJuocP7kYjYZKG1PkxNI
ebLbTrQa0jlpRd881a0p3jl71/Z4/9+I8AoaiWn7hSKHRMfxefrkkQeVJKbw
eJbU80In8unCZmki8F/vk2LVufrKRweFt+TrzPF27xqFV0cl0qp4MveLM4tj
5WmAtYlJVpJwbUEZ4Ai0MF78UK+0LZ8uxNgGUaQdv0sbOyOkhyfkf73rGzXA
RU0bigIpdwfuUjSPJnOjR6LIK6kn4v27IB2RlgsSNyTIqlFaQuAeGwhpuLBS
W60mAjXqDWFev13/xXn6oHyP3TwnVC4f+zj8mTArfAiwaBEyQH2FLt6Y5In0
kzsUQ40CQoR7hxS47FZH4/KvlLM84SbzrYeOyvZNbnlsXu/aiMW4Ar7wqWyp
6Ozt5JcawKif4nCZCcZ+5dqZmkkRndQVtW0dzbVOn/ph9ZJzlfd90QedKzN0
7TXu21Zh1JZhwrWHQ6uCvpap0d18lbc4Kb6fX6Tkzi+i5QwyxDBfa+Qp7aII
2VU2f2u8y682ul8ZeOy9vSx3N59YWdz/GICQKNyFXE5zhfOYddb/qCTGM91e
HKsajDXXuWyQAh2a8jlZTUNTuF+Xhdft+F3rSxjAV0hLfMcJ7V+XHs+bxLym
RORjbsijf8VUisAogs+AfP9s4FAnWMaSMcIaSh6S7fqysYlxxUygQI4Tlerg
QkkusmSW6x3NPG+qRTqNQqkZMCECDNGJlMSk92PxwOY6z2jpuxYqlAN80MPz
iwQRqx6qFHoio/CGe3XiMW8js2Blv7UsANqiZfMLN8bv94BW6eeb/c8lRlyj
otU6SNU1c490h4yyNeyLLUrMsZqzXAVZAOSYeBXMzLn+0IN1nX62RDpjGhWz
MFhGMp5oQsgAZkTLOxz6EV1hLJXHAHL/qcDp8q3LJZauHZEEbtBK/4Tokdi5
bG6WcROBaXXCtbWQPajBSDETGLagj3Tzat+BfMSkmOYHiHA2IJWWIr9MI0dn
dnwIn8RNgOURVJwsraCoHEnhoD6ciVK2I6DsOBFFR0ioVHN5M7JC5o6WDiOO
svoW3fUc2KuJSNsk9jw/tB1WQ6TB/99txfW9YCg30q7Hbl4JoxNe//FsyTca
7CXXpYkMbKZxTYtMUYd5rVO6O8GbnFN5kXK6Ww0FmGpY+OLBs6FzGDDCMqGL
9zw0z+eFzUD1ZkNGx1DQBrBhVYfbKm9ajg72E72L5Mpsr7cmiq8qvJ6bj0h5
o40GXKECQ3FWLDy0CozMW9kQZKoaNqkPwLN0WQFFHYXzAAwx265tDUsxOT2x
RbaDieT1fOioYTq2SXMH7nF9Uvb6EN8ZfgcGzmpEjHmhJJ/czkkQvpqVQhUh
E7WQuTmTJWYPITpCU/J8cIwPWJcRyzgszMSNV1DqRShU0zSif5TdMHcv7YBl
SBE1Y4h91rfQsQyHjC/WRKevlm46HLQhdzJViWx7fzF7jQVKLuMmfyYrObdS
S5rgAdY+0JvcVKfIALib9nogd73Mf4yxl68uu+RXaZp0JU7Z5WJNNOsb7Isx
EZe/w02P4tA+eetRXXK7va3L/5awKNCiD6CWu2G8caZwAui9HrD1KBTdfvw2
iKjlzdGA3LD4envDeSwUMc8BALaJQeBNg46TBn4fjILitLmily2c3NpVbLFG
CDghGUviLglhVNxClTISnIcFZSQxIUYEpwxh3960KjSvIopXU3eYX6DdXbHT
jH38jgOPyH9XPJxEOQdovGSG2pdjB3/H4qku5y/BxVx8a93I5gkD7EWzl34v
Mfj9cGfUL3T2MyIsp0mS0DVReps/PEXDgYHWszj0Hld3xbxAFRUglS82bej6
0NlYW2Rc0FvYMAp+/Rml089BI6MFpsiQdhARcH+MX/GYeYDz68rTsEsyGLae
gG3rX0RlB7WpBybTH5fO6K6mBR6ALKJbHufWajrQaP03IZl5P26q6TsUk+cC
Dasz8A5RHhb4sjraxpIGTVtBFbAc6EV+rD3/6Xg75QgulG32klQavyKaADZB
hXlTa3Mm8ttSiucdyW001pJulttixUXNJUSO1ecJjJfXn+QzJZojh788kIvl
txxHO5NRGwLun2cf6hl4m2t5zY5J2lNbjRYUECQwNV6sDfn0B93l7oGOCuq7
p/2iyhDfXol9U7pUHwIGSSS9SkUNVStREIMXIcQBMo9ko2y7eRqftjIG5hy9
cyGKVg0q3SmnCxhZFP5emIQZjhWsulo2nHtL0dWJIdU+Ib2oWe+jut1KqyaX
6dg2tJWugDqXhE3uNzmAdkTG7J0hWEmOO9E1xqaB6tH4V3jAajHltmpredAQ
RiAoVBYK/dHKXuFHJRMu73LuBidnFm0xpYwV0BC+BYWQ9rIYmJGG6/Faw0Ry
gacJESJqtupfqU9QK4F1lJmDPkiQYe8gwBCIosb8V2uzSipRO4gF9oXCFArn
Ba9348sfLoBDfMevOfj2D6OIZjA4dM1Lt+v7a+80c17XWoFDJBmMIxn3VaR0
RR5xvYxgt9CCOViYK/8Yd4LA5lXqfDBU02JjS5ygNvQRmyYplD0nTMwuQzr+
1SF7I41u31A3zXsk3XS/MMGUzhDPIS9ik8dbConlECSOF8udP8FPi6gsFlwk
dARg+t/2xmHbWUjLRRCORbCf2GCZBmYU3+e4NNZPWx/ogzN6Nmx+GXoHha2h
Rg7CCw7yZXoi4hoI0l00Q0zzKQARTToszMGdOBBprhS9EZNzbiKykqZ6iEzz
JhfaAFbGdDeBGWdz8CRvgjSUZnuHDxLcD7pxsWSEDIFQCWPZVJ7O7jYHhdFG
5B5+cn7JySF+dLvCL4pvJ9USznk21Crq8PDSYojvnBcrjxDwmC5Ez2MP+Gm5
aiKA/R+GxtyMet8yxtgQmiLoMI3wwMy3bAfglcrUXeLjoXkJK4e6TL9JvK6R
LLQzFtJVoBc/oQ554DKrn3bynUit+nhhULHn7/XZbucv7qohCqxtXiSkewhe
SkmHs/G34PB9eP4EVwRoc2Xo9EAJIugIiVdKjkNspTkFP+i1jpDqaQwW5a1W
WntU4YzrGiysejp9hvGow9QfwezZj0eC9WjBlScV5WNgdW71j94GsK91COsd
LgnN0/IGVIdTCELeIqayLwH+ovFm5dwF5+hIXB+U3k8Dg3qq54KfDYr5jfnE
luhwH6Ymh0TxRh0D46HAML0ZZc0tokL4DNeFm6Rqlwq6CknEw58MK+/v2Wur
PGCbnvrkA+UFTsC+BM6BFy6PQaoizRu5RNSNNSylN/xlwqWhixh5EyvLzUZK
Srna9E3FasxTwAnGPvjLzVWpshGxLfsx9LDDIUhtli6QWJfbw+D2wOBxw3cp
oEdACY8a/kpum8W1Xv+9yXsLqBIPz82M8tx0TcGY/e50uDHqx71GHKJwDeXE
jGuoRJ7E/OaeVqU4Lx9DFJvobbQ1WSu7CSP0R2+FOsTuW9YniCk9bQdlDwYB
sNvw9xpyhnIW4kKU/2JcFHz3sy+fNCa3kHoK11roGh+TMoWMmYwiVXMvRgEb
DFcl1rOtmk+m8b4uaP1aDwCJr+WuAXTBlViuv+fM7qmUtM3jLdbPpRDvfNiF
K8dcyOYP0s7fmCPJEb7/ZSY4viwfQ5tG/77FkGuI1P+LFHjSJAZjCdWsJpkq
3RTsjl5QdKgfE6S4ov/eBvpCBbcDZIqjtpUAj1f/tK5kOBGq7FFXXFJ5R2aF
NnipJd5mSrgpAmiPctcSB+j/ZE+5AFCPTT1KddKU2C57EbHj4tT/1liRO89X
cs8GJx0KR2YnTX7MgbppJmhXw8B59VtsBa3C2qMN01qRw4jcdbGAy/pY+TSy
XFAC9GC2zCGED8AsnJHW7r0iq6VPONSYlMfHIinZVApE65nnIaDyDWjUKO+f
tapASft4ldkHTk8Gx754HEsD0bYgsQQjfw9xyl+pR4zufLb1arV+zDEeK1ij
YMrirMtbmRivIPV/GettN/oe9Kb9qrVaSxJWIq2dSPqHknfvlo8isPLkGSay
FQQu36/xVAOpCNTntph29rjQsNcBy9AsFkAnR+oSqa+E1iLk9PI+KmovjoeQ
Cq8TmLhh094cp6UV2he61ZMgkJTtRZ3Vy38LZyTnWooUsrUsjkM+Bg0hwkrc
Ac/8GLq/70K/VCKj4gBxtJvMoiXgcaA0uyeJjLWqnN9icfb1EgaXVnXEVBuC
g8O+aWYCH8yIbT3tqCQeo4x02GPuIwIk0arZAybCDnECJeR5WR66cn1qnze2
vnQLj9rF5K/ZaHJVML9eOCvgvql1i5Q/SIiTllWa89vw4KFha0ue1xh4TFJq
ZukXNsNmhJmDWcrUf9d1hNVzvpKDfx+etnEZhj5pXUSZWIBVUm+dojILtl9Q
/E6A0jkjaONVnMkut8W9vVTM8zqW3RlCGDhdtHNu+eruFJulRIPfzDke/JLi
8s1vxWprPnPXpT/eakcI6QbzcHxra90NKCQff34r3nH2fF9zS1IfRiz/i7sK
7S6515e2nx+5MzqsCsfm/d0R0AOv2vcpBZIm0MAGq+j1xH7ccmYoYkacAOow
ANhQzqZu+m2TDsKdW4EL3MAvj9fWDE5PkwQ2TWQHLNKFOQZs6r3XGSmaKuWG
QbUEnkogcvRGYftbYmnCtXIzS3R64G6Z5T3uQp1CpmptOG42E64AazOCWnXy
hUWYTJQuquDytLX/fWBRgGysbuOF8euv1udlRftZVtJF+vS6I87q1AWZyl7p
dTAx5lTfsg8FlqXSGTgNEzxeCLQJvFyNUYz6BzX0OhCivulNSAEcc3G+AYk3
fL/9hwJt/5J04l0uXXxj7uHtNK4U/qXwNjo1Gcj5PcXGyq9UYX6nM84tKPZb
sWk+TpldOk3wmYxiBKlPEg6cfeanJD+d3d7pfQ1BsZIOMaBcH5nbl0FmdJW7
URiEP6L8AKyf5TqFODFEI3KdvABHf43nkleuXJ3h0bknhEjjzmYgED+bnHPn
I5WrbFUy2QIQzE56j0fQWDMT0mVG6iIn96DDHWONlgC2SnF1kuXmzlhgQCTe
GRcOWhxYHFahpXui5WgfZC5z6TBZ4wqnkR1Z7bN5vjo7yxwBWvA2QFhsnyF2
K8ROYUwHxULqAEddRUEcuB8rhV2ftosk/gCpehODyQWquukrcLH5STWfz0uQ
OxuVODS7AIbDTSyxxnCKQ5UKwrOL8NDQp369jfQF0NdXa57hu3aIdTOD6Ae4
nKWGp6Uf85T3yJfyRe3Eu5RNOcpCNxhXxrWiiRgZFa8tPcM9Sm+E04AnDstS
1hzGKeNg5yQj5wXkwJ7e0cKONInp6nrNEqAhsp4yGLqbsI4PS8igwUAlFwuf
YBGcMluOMRnGDI5s3z7StTrgLjupo+Q5KctJFnriE+6w0QBjkaPxHB93str2
WhErr7iPNOoe1nogmCihSR34DYAw9GAuocyBrRLLSPIht22yjctD1P1HauGz
iZ5xCor7IDbaaZ3Fw30XAFYCnmYhn5y6TLvncXvIjU7SQMqTQXsxBy1cnhfy
YYcdgYjs8S6dywB8qpCk+Vmw5Ube1bXFP/qX5Qk9k57crBXamCg8Phvb2tta
f9ZB9ATaz7VPsWK+rMpFd/uOebEsRQ4Sp/lUjs6/tGXeU6iimEyJE8Sq/Vt2
kSB7OFWDn5moI9rGikTyM1byQY9cX8XOVCmKIZGaRmXbNAxs/aa2rvv/a5+n
1Md8Uf/CDmHpE5B8NIJU31g2OPBUtaEszT52Sz9kDUaaUSGbXjGwJbJTtM9i
COoEbqOsHd/FjlTk0t9s3/xuY1jvDu7i03PbzEuGpXsMn3iM7JfAOgZBzj+s
GqZ4GTe7qBa2yrj/MQuDp7iULg8mzKxCTaYWwcEgCXbXVTqiCz30w+8MEy57
exUyxRR7pP2zI9sL9iurl+Q9JEreV0esXo9Ed2Oo8waoR5jFpYgUeZHUJY6p
Ep2fTeUDcLa5iAe2RIlSxMgumWCJZaxElGe5NzwQ+D1vuPc+6cWn7Nd9gtYY
D/xkTkhWCeDHthYpWAuQ1bEPQiE2gDIMU3cTu8ppjc+70icdKYkbo5eJycb1
5b+FH9vJ0rQpJRXsVPeiLhrYbdoCI9MplD2xlt/fukNJitbdQnTsMi9pFjFM
W+S+LyuZF6S7L7IRUYvJ8O/mDESglLnOroJddjSTCmODFi/eWtSASzqiitHp
/Lu6g86BH0RqlQOIO1JqW8F7mBBL6vSP0OLJPARj4MT367H4Q8e2t0oJQ4Zn
4mQ+tZSKZACCeEDMR4jWrLf9v03psssnyg3hOsBe0Ys1C98tM3wy8IMTpQAw
5s0E+PIWOada3X0tEZFsZ4W8OMI++dOPiCbLFSa8sawXRGJbivNGMil+Tjgl
KroaoioAsZC6miMxEX66RsZJ9WNXVOtg0u3eoe5kvfB2VQ9gB++8ypRx+WNG
48Bu4fildmRs3v8fXFICUddRMU8r0H8Bd6fVpxaFdeUohCJlYVbMvrfaeofp
0f9pUxpCs+Sq4GhoDpbaQRqv2e/3Z5qad182SmtGDl6mioJBFsuYYyut22Vs
iXGu5wHzBtK+nqlnPe6Dv2q/LmNgTIKdZWwcuYBO7o3kBP15G0+7ROchBQSC
0rWlCS8pv7ILEezeUGLTNNHlJlK9QORn3d+LYHcstbqPgX6Fz8N0WdZVWf6O
8mvf0SU/oInt1eUiel/0vDaDzxidQA2e2RE0sd8nckwYw/50dzX+Q7anzgNm
Ei3+yrk/hYbgD/eqh29Uu57oa8flvi5YqONPrW2YfuAW32ScO0X22E7NngRy
QI/6o4Gv1H7iExS1ryXI0LYxDY+hghLddMwsdchLbKyfyTFnIQjNKmJatRbX
MTN1UK8WqD2ccntWflg7vfbNVSkEv658zOXHQ88xSyxvYLwHBXc6s/KW7sB3
7hmseQbfJ+vRT6vRTRbM/HLRNLs7ZiOwipfcJAXFZPlCF5oOceDPpUEfvGuz
O+CLyWjTC0nw+u59NBmFYYqZnbFyMnNt4h9vG7xhXTJYGb7+8VYxaR0VFNG+
FFON1vblfA/8t18QNrlBQ2QB0WmOzj0D1xDbNTuVKnj71VAACdzoIcsEh9dE
ibjIfGmrvIFkAIhvFb4d5xxgHqu9M6MDsU05Q2OYVVyr/E2dRwxziGlMw85F
KX2xM5Pe9vsEhuX8hyyukoNM8UMPqjCtUtTxOXHdn83SOM5HdR6bMOfP2IRB
O3pO6828IXGGC+QAohwk+VC8TQcjDVHqatqmLi0JQertU4CMpb0tuOXEWf2l
jn20ye7gDZ/I1+8WVRXfVKXCkVdlb7xz+t9Cis7epc6ot/C2Vd373d2o/R8H
09bbuDhJeFdtPYCnwdeQQ5ySFdsIO6f5n/V21HhdNl2CUEbrprcwpByivzmZ
vB8eKjAboGROSh3iGI2QstHQvsdNnT1hen2FU1V26ad2l/IZIRW+bTd5sY1O
KPftLUbOJwZbuV7K2HyAYytoL1HNKHgbUNLXp9ui3hmwbhQE1cCQ2F1uxr4X
yQWmcetHuW7SJeZiyjdWWMzER4+iZX+ZjXF6JC1RS+WVlY2HqdicJ1CMYFvK
nXngT7uPFxNekFxo/ttleZEsIZbDMjw3t2+kHkLAeGn4ZwKSEwg/c2iReTPa
TZGYRGpSQHnhX58Ev815gKIZjeVWLPbGLS7/SSeb0PdxwS4i1pgCb/OkruTI
spoxX79J7d6q9sJ/MJfckqz6yNuzvmYDC9QBcPR1xfCOPvc6bsEH+XTtjIE0
4kXTrXkiF5HvGmdvr5nXdxFQx7o8aLkkwQP1UBcpWOUsEQv5S9K9eQIDpMpL
nXzvanRNMOKtV9bGTDoDyzWoaM7NROxUf7tSONRoGk1aK2p0dQCRiRSHKXkv
Ohahvhg906rK1TdSL+IZG1JntvoEn29CM5p04T3Tfr58aLeIiIYMlOb8R0Y5
eN60umj/IxGdi/6fv9zI1fEwzg7kVWTl9eDdl8pfDWQQpbSNYQ862fNGn6e0
xXHxXiZhYgQi+qu/5IIwCvehJv7/myqIk1L2LNMDTt7ec0i0DyZam3O3OmLL
ps3fAPD6+KQYvOy5zFlOi7pFf2JEobyPMAXXUFJWbs7ApW1ztZAhMT2e77ta
LFXDZIKCj03lJcz3C9dbQqrYZg56f3ngNS8ZGPPgipC1OQkeXfGQL3Sb7avv
b4ZJ3GG1MNHcZY58S6I0QlBIk918beFHQs0FYmiSby5gn1/HzOB6/NoG/5aV
XGkDjrTwyuOossqtxliHLX1liSHUNvMPqSxwU1W66hOmR9ntfepz06zpiGgt
I//aOkaXxHlAjF3wusWS0Ukh6f58RUaB3xlSWoK+XnT0183SSRn94gMNvrHx
FblbKexnnt3jlPY7N19Bo5gJVdmqvkGBk5PkirSdCHyLo3q6gbBgHsoxS/k8
Kk9VBHtggLv8pYVy0p1KjwNSLFcmVuAbDhX7hKYWUTI5L8n8QIhqaGPp1lTi
Z0L6hfzd2MtZ0LEHbpVTWAnYsZkIT5U5LU+RpDbNDnKbeS6mDweNtuZKc8qi
4+r059tZAOG7gDL9BmGfz2Pg4C2lCl0G8B0i7jpW0fwxlm/ApxHkErcA5IUp
BBqvi4eM+/wXk+ruHPW1lKhnIjUJ8yQ6fNgaOgmFPhn5gBcUCmdehqZl4+eY
u+xFFaIsCWuT8Z8CCAANC1quxKIGWpnhzNHCLcXDXJlY2OFWRqNbOow6oyFx
z8IMsCqz8w/VQjdYJptvUgKH4cCtBHOVxVBKCNzSwxnWSpBtJQvypKkPoU85
rt8drq3KjpC3NBiaj4cbh1kCrKVqy+6b0rz4ylfdMjuS1dde7LGZ+ycLFyIE
EHYGbI/kiZuA0S+nZREsrH8yBMTRHMtcdx2Ja4zjydE06Yd2grdGFJynIt6q
g1fzgHh1be4MIwIJOv0/2ZKlZua+cav1Xy7Zncq9aWJ0IWVRyvrtHTKfcqYF
0Ji4pZhnp/Uy+9mRVffsfc/JgHNuHpnd1a4uXto6l60IOneCgJx8MO9A/Q8e
lCKkezRHbW9TgOzgOPGwTAIBqJSdo0Ahm+MEnDFt9mb7q3lIxnWLECskepRP
PtC5xKwwO5UbBrgmLgZY75AyMmghQ7NTdEq1fEubRNYTSfNemoEaF9JjSFFc
rMagIEZ2v+jbEwzL3ZTiRrNSeZJSMW4NG0deCSHqpaaxEtDobjnEPMlJ6SHI
b2qImBMYHmwt85NSLco8utBBj1mtTZji4dwJLm33JV+n7Fryvo0JPVdf7kZb
chy6wOfpwTBC9wfQrCKhe5/mDxOAZxdtHyFUxxtyD3AT0Y2q0v1SlbrHqxas
psLtjb3zBQiohiTQNTNci/BsV0hgnGKgLrZNJS5wotl16U1uZVplm41IjKua
GtSrcqRgGTXlFJfrx+hB9H9oYmEum/4Ze4Zv9WjGTaYgnReqq5DmKkp09KV2
Ln4LV6/i+UUBR2ApUW0WeroZx0lrYCirJ2KhhVOSrB8+HjTC+yZvmUUtubJN
I9+PXCL2EzT0QEsxCLqwjUm7Wz3CVISa1ye1L+mgWqtzFyLJbDoxR9ucGxUO
q10/SymrWiU5K+IYYzBpxZqrRzFfhERF2u5/15ivW7oz3GC0EeGSQZiaZnps
SWapttCbTLE88w0E2ZGqniIV40ZQg/A7pl7nc/F189B0VjHaWZ0rxPOH06Y3
3XdejX5cRd1GEj4u0t/8vJal7WxrToBDsrFgFYTpk6pGAN6LeF0rrnCcbcG/
dFg/jzDsw5LR58xUOcZ7Ud8O3ygDeh7HFIUkYqdtKJ9mYjyieJrQUOdr9gA1
XGRC5Xui8iKyP+Jy/iQAYSzbppo53ak6fsTMv/iyOljmWA7Ie4BFta4DLKRQ
079j9Omnw3VU9hh3mDvVCpFMuT6x8FcX2fBD5kdW79I/nzdz+USUGnn8W/2d
4oOx6M3PqF/s+R3qjNv0cKZU5v5S3rSBhgSg7C9hbKLLsBtwIPX7aQsaMF4G
fJJ1tDcAqEAUf2l9vl0Mj5820kdnraL950x5ZRmN8/RGOLXC1aWOzWlfVeAI
sJkU4ii7OTmZjq6dDo+RXE2ZCCcuWyGbhwpR3Cg/vnGp6M9pEYc4cm+KsN+Y
Uu2GAT2CcmuJK0xZu4tiEOXA0frctcS6YIkyhNO8jsEqbSxvMeduf+Xs8fGf
TB91f/Pxf7thhjx0E1UL2NgK/BE/mGg8OsVl3a6pRb7cmiGALLOkbBf9MgRU
4Y3JN8hVVWHSEKxUBdXYMZwBIB85BoB0jQXfDoWU4s7NzPkkuPQOTz9+KXIE
ATAka1046oK/MxcEhahjpAnzVjDeLK1+TVJSwy6CQX8Zq+3RyGsVK1GZ3zmU
qPXzLEw/IK2mxYPXehgXUdq2WD/8Pzuw3NBkAEYOva9hLfs4F2DqTZBxTR/a
qiADwFcNVOKKJrIKRVAMdrDxwtIyZxkfBMssJQdmH33qXx/z8h5wc+/1esxo
qlFKy8Q0pioBUiI+PsC1quXbCvO0pG1Q409A4wz3RjWGllSURbdm7nqsEYOW
Jdn5p0cXPLguDxyudcksgUxjNkQTBS+0cPWkhcm5MjVaCPXjGt6eFho1GrLJ
u8JRqP88MQWs/HzIom5XHSNmWd1Kypdk8Tq4VkzWoFqRAZjFtIBr2EqbZSPL
Cppn6zcjGxSDH2bO+vdj7jVBXNgNUWiFYLX4n+wAH3TF33dvRueAoVGRYpyg
3QbfcHqKYCcEJgnAvpC63k9yDlptVEB6y0h6dC0I7vpJBQS4BmAivL+Qxtbs
c6MLX/qQ58VIMZmtejpu06UqTVlvJz8k8mR25qtWi4PtPTyRxjmCm2dmf8/z
4aEagJN5uRGB3bXWHETBBT197pP2d7lEDgbpsUg5il3zi4ElSBtl18Ng68HQ
vBEy0xIk2DcHF4meLkFBAw698XmOHcxxKLedjzq8WCPI7bqoq0B3eArq/oQv
xBIt2c1d7ILJj7tj9Q1U9VOoYCUktK3HCNwjEd0+1PwvbK2PvnNkcAJvEFSo
s2FEJ1lecX8vuEYEZzI0yd60mO3Q5tuOyshKABXy2L0ir0Ge+bjGhPCSWqQa
7O67jNiX3ePxHiZAQw0PkpGSWUETOcdhSu/TGogjh8pHhBErux5zRc3ZM8r5
7GfV+0ZEPHh/v3abUI+1pCXNyxEKnrnXFIZmpSF8QBDEQf+i899RaLCwGJ4b
xeCz3gFKJGr7ObkW1K/5O6u/4NnxobCmDLnO5/0NWUSn6XciuJNXxxGOf+pO
5ALxpxGXghT2s089dRg0D5bZ0zz6bVDLzXvVivAUwuoaDT8fGw7vrHWPaGxR
TDD9B64u8HwWjgpF+g6wBNv8roV+5g9GD71Y4UFHUTLaKWIyxWepzznSS+K9
dALvtyjEuQMXsfS4mlq8TPhOnwR96RqSFN4A5zwTBu3OybQBls/8JwmLGTfG
stY8Wk4Ej/mBr+d8pR73dF+CvDshTn2XVi1Za4Om8eokrJRkqo3dBsB/gkFa
BX1Ze6sYTW7VJsLRzzfcFaprOfCH6DjvQXBQqaQ0BVd3NXD5o0zMS9OVTkH+
Q+Y6CsHbSk81nEStpzXTUp0cKtGWlytjPUnXimLGsRGzvddfZO2uIPGo9bJx
8VqEsYYD4mhiSt6sjMAF4Yxu2tOYeJdHO/jwfWKMlmHaS/FxEMmDoJ8GIzY8
IbrTbAElPhiwwf0iQRC5k6n1sT9rGLXNKQ8PBin4mcpvuugIikwYWa+j9fd+
J4W55TLwq6A3Y4xhJc6HNQwKFpnh6GmTMxtr1o28Po3ZQU54sltK6yxnuGJb
Gn4RxDIaHq7+FgH0dibDz9W6DF43i4H+USaiu742yt1PJFR+jjNmHPwy8UGk
cmOrDGuPuanqKhEJvapr8slAHi8tn+HZvghf5ehoDXpXnwh8NBqpfA2CVfZ+
Q464uz/bp3RTEg952f/NlT7SG6h5CpVOPCy/trBLkWqT3b3H0HKB8nM13Pav
VZyRirj9AFuikBGokScO/mjd32x+5GyMhome6DNXjxSVIG4E4qg9tMEgoZEZ
b+iO77mYPUMQ4ahP7GxR6eJ/rOJhGvpQcBXOuZT8ekdOt6PZayKaBbMUMELh
zGEO4fnv7N28bsaxWx2qeFAOwHVRhl6zi81D/ZMgNu8pCDfQGJ8/5wUCVMhO
sqzcU653xq0/Lf+hCenCRD8a3Isdi4lbTJxcxLA59P7YA0k07h+s31cD0N8+
ykNNYWbH2mAoqaaniJH8hapPBkgygFC9CrlcIwZI/+iWWi78o+GUWwrWUd1A
j7N2UIFIO6uQkXd4fMhyWseAK9DfP6JO93KPYROY/LwmzG7d8hNOvgEr1Kce
w2ayafUqcQCag659ecvi6a9OIRZ0gnQKf1s1ptiMIRJwOXF2AFffqcdYXZDU
YMx85fg6M/4CLYhl324OxsGb0iHHfLsqn79l/f380+Oec5iJt9EMmsgIcZSV
7sTvblFCHvPt4t4SVGjZRZ/iEZZj3mT6h10T8otpts+atFkgJ8Yu+ZoQF0+e
pC+t3KPsCp49GwSxeKqHniujvDi8HbxcQrpCbUtVP1Wj5uOkFLIt1+Q+KXbY
8oM7pn959YP/9JgQoxQ3pXYFYZr1Npi3n/jcmgMEnjLVSMe9w58vLD7Mms9u
gDSTHQzXWgF2thUrGY3MBMVrUZIrDDW8T5S42aXfTLaHQrjt+il3zU7bfpfl
yz41AwsNqEK0ERyPCpeW9cwZdT+8QLmlAzkpLieo2+2MwXGI2lMcJLCqU9qY
N1LNDlQcyTeRbWXriSQM1CUb+fEsAe/2TSMVsT7SgKzP+R+dD5SRx8d7y2H8
81WeZXXPdELKxw3oA/qwFMdHGcIDR6npDVi2gjtRcMzfmTGtYtbLXORaFzgd
jhdBfELYG1NRYVoUupa4zSolkG97yu3HbrM7KUc8sg0Ab//lWK1XkeiBmDYD
LOxUOJ4OvdmoNreHwA/Rt+9VKn2GMzhWbuV/e2OHmRgaZ8hAUBmjCVe8k1gt
8srWxp42pt2PkelBhQhrWm0NDwK3Eg06VWiw5Cn2TJJ/E1zN8BLsd0xwX0gT
9zmy4qYMM1C7u0syK+Hgzx/0exfxqi8SHpTa1EO+bvTx/OQKRg/Vv2fQdGDN
crOGZV3XvPvPgXB12naHEZYMOwT7b9bNJBq0yRwuv2XOFFbg34Zuj9W+j47l
GMJ/wY+MpyZXPcHow6GKZ7TqQPsm2x60YASVz0/ilZN0esB+g2yF8zj/QiV7
tFuO/ynHgAnYWFaPPjGdMDyW0zR/eRQ7fn3HZLZViBWNKvCJq0Oxfr0W7sfK
uQii7727KzPQuHQtmI+bDBHio9OXarCYJompdNlrKMGPOXLcmCrfJa8b3Lbk
22ILR4PtlXyUTz3/BgwbERPYUpFdjz+kKsUK/9mN34GRsp2xrZgHnXGtO3GF
HPv/uUyIxCSGIHnZtF/JysmeKsQD76o8ShOwklsRH68TkzqU6y55ecMmQ9Tc
IVptXpt/C8t914ehp4H+0b2Cgj6jQUG+V/Cc1mpIe9Dkwv0jUMl+Ldq3P0/Q
1fYHKamihTdhxcYLOEmlhPvDjOY8iT/07qRa5R66nKpDYdxFX86aNlpb91Kc
ka//GUgJG3H5Pc3wzsOXBQDFOSSIncrTMSWr+GPEIhUWecrhnjL8JNN8SZO9
ekHuELahDYPz9BoySELiZ6SO6rW/UPjGSafM26+vNbkhgFDxdLcht3v9lMHs
uUssw3hXWcKge9gG3h/PW7zT9XhiyJVHU/tPzEdb5vW0K2TiwT5kNwtz/D3q
028pEnl7HkF3bJ1kq7rsmQScL9gAPFh0bC6cJZw8bL4KcaB7gVgRjhZHyxr8
xDnamx/CAxwrn8l4BUPHbpG2gtgqAFc44unC4F3cuuPanYuZW5bI+Kc/cYS6
IY3fuI/Ndu4fMKbww/OTip5dKimH11gx68Kn2EZYOvbBAhizyNf0skBV9Kcg
B6gEEFxs6ZWSDm39Y+f9iaVaz0D7FCcxTublEXsMAXHuSlsZvJDVuBTkYJl/
+r1qG/EQ4/VD8ww5t42ZCa+40/+MXk67cw3fZCCB1bWDzDLJKhypfkyMxJ1T
ohUUtoR/v4WQxJYR+/Z9Ag1Gi3s8vgiEXQvHN1YQHPnCjP54j/b0yBRgh+HR
lOTcVmT+0ZwD53kqD133uNzek6NlkPkdB/E1YWUxyimxKJRMntPsWmdYYQnE
lCHjAeKoffEKgE65mopsQVvDClne8NiTfjSjyRD1rsXbx9Q+/LfhFU3OgS5O
KnFbc0XqmnXKzGZtg4KV/+AfN/KD6g+4R5kOjyUAj6H8Jx8Av9jsnHsRC0ft
up43VYmeQXiCSo9vf+8eahTybqH7HKkZmJDJPKQf4E2geFaJUO2YIFgDnSfd
9jIgBsB3gcEs2/quvRlQi6H5vlmO/bqjsYm7s1ohDbi9X2ca6UMMRLfQHEhI
65VW13xpF3SvRxwQNBno4Bu5RJGVIL+1Sm8DFzek+vUwdAG9OpO6UBxJNJWV
vVhMoSRu5IOTxzpmLQaHAxAcA50HeWv8vflvN0DYGS9ZO/vRrBXky6kiofpt
RKlMNzMywFHXqOYfsGetQ03zUNwF4+jza+t2AkOzThIItV9bOS1UtThD8B2X
S6y25quXgfLp4tE83FgkXPqdFq0IRSj39gmpkKts0UUWoNvMW96v2o9nlmxh
2sGm5qlYmGZdKPDQuSjWDny9S55S/eG3Tz1wormNdSPJxkyjVCB3Bl+ixApm
Unyf3EzrVzFv4BzL19jh8qIMPOp8TW9l3+DJOYEaWp2fGHqff3MxJ0vHLaZ+
WHU21aj46YM/6a6G6qbaG3XoqhWI8lFcvtkz0ioFQFV7lie6iZPv5twNlSI8
vE1WpAtmOHV6ZBx5OgARqnI14vI9C49SctiT1QQ/gbSDfoC4nT6lBRPkSrDX
oj1G6T11loC3+oTNBdRmeCZFBvAvXIR+Bwu64L4ivLOwzVsWiq47iXMW4jug
S4h/jMox0xnBSMDf4ptkUn05twtX5MwMytAxKRsBs5CHl+S8CAcPZ+HWfCKp
35Tnpk9bagpgEqlaCj8xV3Y4opTS5sg3NLBsItkxGuJMpIigZsfROtIWDsKK
ZpVE74T/PHrn9Gels4QuAkKZn+VnBh1cegv9jE+Yet+rbWJ0R8c4znwZdx2N
fgibj2HpVD1ueQN82YXvQyKwCjr/ieCAAztsHkrksCgTVDDWZNV48O6hO5mP
pAW8TwESOMxXdesvbOZmODlu7A70X2Tgq5qchlJewbgohwm22Y//O1VLtFLS
bXSygppmDbAbERH6QKbk0WCqUNL48gEbIBIyxBL3RVz0aVcJORrppK8nZ6w+
7iGkrlGWp9drqNspOkCBdmbS6CGOgcXupUzJXG031BKCyLvb0q2NUx0sK0vi
SYyfgGfn0/cc4bels0Co8dwsCl0gw5JD45XutkVPfp2Yl9hZMeTDGXceqV5m
CHCwSKs5gs/HWKyyzcMAZdqqmK//Vb7EnzEhxAvsoSxqCckDIvVFzuyhCa3H
fUvhmlOS7UthnPZVWPYpiFwNe7oHvCy6LB0svzVTseYLPEFN5uOaYhUX+KlA
WqicSKSi2lSWU+MXhbq377ZATfgWPMrLI+L6fpUz9iYBkjKEr9tW5xA95vFy
frscPu2T6hmdKO8oGDEgt+1iGhSc57bk4p5Reo7+SJrnWl0SBGNtDXMtCRLO
NiPWPcezxVSWLWrId6qPpoPtDtNkIHDOwzAR9c2X60JonfnotipqhjmkvPA3
HbN/NGksgmmva/IfdHmoNMZ0ZwXhpjlsKe5pLjvG781fiASDO4k4ve9ZmpMp
/QTJ/UrZaJ/gG6+uYnCCNlvIMU3Wl7pjz33Y3SuPPZ/4S3hNKbAF1U8iM5qp
24ATpZaVc7zyD5oV2cSJOEwcR/PzFzBabeemmJUQTgNPsUoWEIWyHW2nZy7S
JtL3txTKU4pgi9aYQVSMcpmkqOa3240w7mBsfwPPL4EquSkUYy3gWGmol3yj
/KFR1r2He+pDuSKSyFUYloJtJTF4Elh9c9YcNpoI4UrfFzQLDe6jpA6P2vcN
bcn0k5HMrPmdN3Q5pKqBvSNCpFn9unrUUvkigi+5tfDE8R4u9+tQEh8WdVk8
DmAd44BcWh/6ZrOUbjK0fRKWPiv5xGB6cj/+EK/C+LAQSiA5jn9VwSuQwZyo
wALsPYhYEnzvPWTB+8xIjHf+vH6KN7LRQFUA5Do1hK0sSbKQ0lNU+ejKF4vr
65m8ormE8Xz6xSuTjbbb4ebJIO6TFMfBMtCkBFaSN9aPh4LOqLxCPRSOXb+5
LXKfthLL8U+4jh/yHaduIO9XQ/12Un4YSYQJf9ujlX7h/Zu6Jdrg9BJUTzXg
2q8suvkJkyYT4U47RLAG8dwMJOy0iBAsC5ynByXJ9Jx312qG3GhZDz86Ss5v
LZSkXDPiWywJ3Ui2pka3RMUu/sYUpsIfFiGHbk7nuy51BQIJkuWdLrVLexD3
jUiDk/CD6eaHGVqzlWRaDCJ1a5uewGKFziYWCogcDwbXkAbQfuhX9ZdAfQhO
v7laUE99L2y7UTOZ03jYZ+bJt4z9TQNfVduBs6RQ7JXXQAnr9PWakn1z+TE9
3wWdghz6eUmnjFjSTH/LKOf1NAx3jhjxZwZfbrJj+9ZpnAfJ0iX096ekO5ay
3JQ1EjRlevOTe4eUIUH0z8kkPfz9XbjfsXZBTpsWwbxn8kSpJZpaKfbM+y88
z60PxROUv2xuvnrocIVTtQmac6tO1xcp27nPhvwe2CnFlXaOSxETlWMgOVA9
4O5mxciMyWC8OyhPKVVZVSYLsr98Y0llSfbY6gu5YYoQldTDTTLvUjcHQIcJ
iCLO2Fbc15zWftMN/Kemm/+L7WQW+ry8zJP7O3cpSGTMqxT6SMfRMEowDR0a
QhBLMr0bxkNGjDBYRc76jRhi8npfydnCV44SVfExdKBr/NGQASDg4sSEc+uI
h4lTVfrg7E/nNRE6RKI/koA6QLa67aC6ZfnMYCY9Rt6Ls6lgMipT9qfG/HED
Rb5wpNAKrQFTBhHF7KCwffI4e3WfCbVtnS3GxS1Qme4xRcKO+PeYq2GLEqJk
7pNvPVoc+c9v/RdjkXriGvlwuZBxodbQUeIi//aBoYP6pv4dzVEbC0KTK1Da
yGIHV7PLou93v2tUCOBRo+GimKYPXkbvRKeamafMmVsXCIzqsGM0jpxASylt
fdJbIwoaQpv26B3dZIZBfT/PvDRFXIVfRpL3wQdZst4fyaMVaJdfaVuluwxl
jVA4L/qZvqXCkNNU0/HpaSpDHJU6IduLLVvtRXm+iAIItUqTTn3TGq6qdEcQ
y9NA7dcFx+S/1yKlci6RF/9mscRsE4iXREIc57cbjv6rEGjaIjOidlxB1JbI
+MJLj44SDd35Fbjq8F09GGQkuFWijdGxPxN3LwYRs3/PsxgOhCIEVmqB9Pt5
JE1/poabKRhCIAEEkInaRKRDdpZuMxy/loMfHMLkuOIOI323VSZXgHCF1ev8
rji2wxMIQAJ0vepeR/7MzwT18EwM7F6DkgqA5/jFFS4WvL346SRHRBVTzkm8
8LZ+IOOaSBE7aXn4maBB7LqTCESy6qlICZYdaEms7YqlQXB+adnPZneBducb
ECTmNtbxrmf+qlFSOQFvbk9rOBTrKO5Uwkm01PggwPmWVbpg5Ks7Sgqpj/7E
hzROz1hxDb4WlZKmIXam934AO0hTzk7lwnuYgzxXdN8goegcDWRRKc2zVr/A
UreVOzfoDx9NwzMtgebIcpuSVv3Tdw9BaLCOxUU6UmLUZlt5cBJQr9zZM+rI
N5FpGIumZNz5u55PrBiKSq2CxTcdKhCwXf1CEcdASAGpfsZ59D64sTsM7hYe
vaz/QOK4/bv+kZU4j5gWcoHm5Tum4CNL14VHNssHN9TtmtxB+3C54nM23/iT
x1yQSCSK5knxXoN1fwfg8ou6rpu+/cz8H7p4QCeujyxHemvt2tGN40rucjBe
Xyvhxz6GB9DRo9/7vxNUKuzSfjqEWQVdrhRZ3dQ4PlS6GuIw9H2joZXxfQyd
0SQ+ZY7MVpA9LyuGJFNT8R8CWIqX4ayzyRwwOcogFdcmc1+5tW6PXdCgSs8g
ErtolTswtWf4RX8rMuTZx/ytnn3rRqe3MSU225TXm8xukgshvnPJqwAgO+zO
oob8i9BsZhrR7fh5zOU1KiLJeuLzyYsxK+D0RKjV3Jl2PRpCTmg9s5KZtXnD
tdx6jsJFzTZhckOdE2L8roOzoTrdXqDZ6Hk7TDID3avO3BjCOqQM5hp1mcbV
slHVtO6xdNdHY5zNYY9zHvSk0cvMefQDM8Bk0UrGTCABu2cELeyKK/+IMKF+
GiXCVU2LKIizL0v6ppyUs7+rKDMQWzESBq2sTbW+ytmDWiVJng+hx+Hi/kAs
TV6hkAUEygEAHHNrmrKMd9WPIZOneYsgv2Qwpfs/R4QvuJTbhFCxmMcJSZOF
EOraOxWhziYYnBFKEkm6jyrkvH+ylS7hcliDFTpNo69YH4Nzf4BfabpSMnoG
utLROvynguukOoq5OvFlkNADNoBGK3AfljCQwu+hKABGD4i6NYVMLkLD0O0W
TRc+X0/BnXg8EtI78Ofqc/MEf8iThW0TJL9AjRpGsP2GHzGFCeQUTxrawwhn
mmkRqL4foshEA6nB+JPVBGvWPmZEHOfyxbQgW1Dq1IcPOQ7vRjbiBeclVr80
Rclj8vYMiAnXKK281nfWc1iaCN2yTOBKtyN1HReMx9LAk1ly7js65aYiobAs
/x8rjkvn2GI/lrw5uqHTg4gNfnDPIAdHttvOu8kYXhbQmtLEvIu7tIm2q//F
b1A4FYKNkwndeBiQX8wxYGmEZkL4Al4lPCvLgrbOLMJuVfJ/wns5ijEMWMne
FQLNjCPdsmx893+Wx/k2eQi0cX4dw3cq9Of/6K8Ut+cUP5/9ekRoELqNIauH
awh/eXSNbxhOTCgIXFS731QR8W2Z3NbrFdJgRlD+EZSe1LoCCFE7jDvJsZhR
Q0fpkW5tfwM5AVdrCxOu9lsZi3XO/68OQ/ygvbhxyeDsiUvZEaDicWpM+qG3
TvHZKHECngkagf4Bm389oDVXkYDsYr6cmeR62zAlcRPbnxSyQTYh5iLxDaG8
2DygAShng9beugG4f1ZJOj4lKOPNkOwPrQPfwFqEmde3kc8GuadlJn4TxuQx
6QsKDIgurBb0bx0cFL7uKvJ8c3EXQxdGVbpP25m1sSW6w4bL5QUhtRDHH9TK
w6U+J7YMTtjtB1JPdKywMHQIJVCeJgxyllrSKkJWsFq8GaPBI3JnhkORdKaM
s/Mlr15GWnZm+9685cGdgNNHYCG+JX3e+8mUmsaOIylhQpzDTv28TQPE9sCK
IfPJkK5D3hi2YiTlx/eALh+Ovft178hQ69vHTTrlxs5RCDNXwp+InFfG73N6
3AywlLuV3x2wbquJfC8pCosublNIG+Bn2c+2+QeJtEOyn8JsP1aWoq6Ju5Hi
YyQ96wtgKLOZYhQWZziNP9oRL9CDoyhB4OwSnVMP5DMSb+AEcYxsfonLrDq7
asgBIASMvM4B7iSzTVh/WtaOFevYT1xzVxOuR0jyLbTwM5vronALBL/FRNx2
NzKPv9nECWJbpnWPTWom2nG9TxRelYCKkCrZQS/H9m7ty9AHUBj9xURf5v3q
0V8deViTpYPq00iK0lzXWOYDlXgHrVgovdy+9qd8uTFsNLJLtUOUG0ZX4QHJ
kZ5TJ4hVl8Sk3BjkK6R7gSIAimZv6sOFbqpYrwdqerynhru9wmFl5THXntfC
1o1W3XNecd0CIBzq71VLpbtMAkKZRrcH7Z7Xyjxr3J9IMnt0LIwCgxC5tshB
CTok7rfWM2HTIDbdrVGIhF9Ay/1OCtp2CDccxwmlkWurhvuAZOyCzq/o9Lia
TC6eYYL+oxP6Xwy2nx5dqT3SM3bqqVZpj3f3ffTqOwNnwokqEe76ZhncH4iV
Ox+sZOldrgwoppngicaHgnx6YzfxQ0S6hsI83Wx2oy6MEwOJbFp1F2KxBGAq
20KWuBq4srlacQw9KhNDjEoqGCyBex2tJvRWSdhY31sooXRCCXphxkoHWfEs
JUEhK8+uMoXFXemz5co1NOJVa/arHWEW3LbHMrrKbI0gY0WYPQz+7w+ZyPt/
X8//pZdji6DHxsiz4PWquWk32YetBr7w/bFMMVfKWKs5yZXSmkTEnpkzeCUA
sV21p+xZRh0wBcKnqNC0G9dynASY1EgzGacEimwGmrqCr07dVlqD96+7ZchX
D2hIgSdFEvQE9levc8541tzbx8Fl6L4wk6WQO+oKrAwc9FLLiB5XBZbhwt6K
XpW5/IQekBtNpg3gIKb7exKbvaCakFh40cn69TTowykZPBHHGLSaypOsUoWy
6kL7x+N44mjigC986I/3wOfuWWGxZUMwH56IYaDJAohNvT/n59/+LkC+rtYA
VviMlwh47Z4+qnGM31RybWp5JWSvUeVq36lEpKQg8hiq1Jrv96Z9p3wpvD0Y
lVZFDeVKBE7NAErySgTI33tOMBxjQFL6NSJtwepT8oXR9bBI5Yxr9lr9ozJj
RpbdvtMB+04vJeTcX06K3qolXsgHNpouC4WoS9XCG4UFYuLRGR0IgpzA2SU7
O3H6fI83rYx+hb8hqBklCOLVdY8wZ1MQXpS86R0M2sBva1pf3qw2OiL8YF8L
A/QNSoHSGRr861bDSjQmi6Cudb5la/p5OosCLWEfWa1VJrqvIHnMw7u9fbI0
1mhmWGecF+vHobrW8ya0DZuqMZVpeHgE5zOV2iYBnwmek0UkzF0JeHySpnyX
9/9oUYARvkUfWOqJ77CtcrF2aT+FVrGP1LUXfDT6nQOs/Wj6syRKN+UbNNhz
OMbDhxAnyz5lrWBOAwTcU7+P3ECm6VkoxMgLPhBl/Z97g490DW5fdP4b7v/W
+GxK7goxqarvYdDQ4oPXXJb7KrPejZCTItAbdMDo2TrUbDPNoHBQqjXthioE
Hj8q/OHh8lmVURddbUlURFet1L1divVVr1eEDNQOA43eg2jevbN/K9xIwz05
7tj6Xx9N9piNhVJsx+3LwfAlfv5thQ/mUv0zgqLDmwi5nqrs4XBKIcuTI1s2
YCgl/KWOjzt9wJBHfY3+fVoXCvO4rai69l2Pz4owOnNR3i6To6QfILGft3gq
BDFVd52WUgsQeZvNpGdVR2g0PaFLXF83rHHyUOH/T8Sb4fVnQ5IL9J+SyKQN
rjfLNAM6Yq5nhjVHyUH/qVZ6ASOEc7r90SWbjFWv+f6RMGz45Q6pFcxrsKPq
GAdzO3cNqternMwEYSZsvViixOrn4bqcE2kFL4okfHkz8j+Oon35R0OLQSkv
DV9fJI9q12GWqnqBAxFjhFLUo/ifu+59OBTNa7gWUPC8E0Z/1FOZYbR4ButU
KRGaicfMsSszhqd6UuxFrGMapc0VnPH57bKpLn7Rhk0TRFsmEmIaFfwJsCX5
+tmYkd+Df9AhX+M52+MT6CzYjKvtA1W8Kk+2BhQONQifVkztjVnQfa6HCk0x
sO7kpCBIMfso3tIXhgLjzccUpfsicfdw0wlSLih08VxQRFZT/2AY7DGiMOwd
x04fh4n8t1AEP5IaagBRzyth4HY/3Ty+dXeUjSa4d3L3Ya1QICbRUPx88s56
RkOupDsBsx5XzEt/TmtmP/3BURyW39EkQO/hhuLM/OWTVS7pQfOstpKIPB+5
Im9VK12gkMAplC2qnAwEcgDHoFRxurpwnDH2goObUvwmKyMD7dqqgOBkpXE6
56Bj9liJJU11qsg0s0QwKHkRzAeAdM5KDRk842dNT1857l5dh1lfk8mqfSsV
CggVLqLYmjvxbz/gXQGv/3zn3a/+ivVsV6weJe7q0DuOlStNnBfw3GbDCP30
E0buv0LR4Ot469wXhcJ5LkFGq9m0gPUlzXkkuoMtackQtJi2MB8NYD5lKD8I
W8EzVLSzNbAbqGOXohObWrtX+1agKcCeAuxve01dabZByl5bMUAjbmKYJny7
tkNt2aXDdFyPZMnkJGUmEuFBx7L4Hdj0xSdfCx3E+ZGKTeKwZv1RgPYyGYtI
zzHnmOIS0U9nfbE1PSfVsTvTX18f8VxeKs34Hy3o263RGQuF4n9CLXGPuiIB
qJrnufqelN6PO2TAufPZeXZjr1YN6/RfqDmyrug/5tKSF8zSqbeAq2MUfSDZ
jvZeylmzmy2p0feYZNgl/K/hlbb3fUqo5Ud9c+DO8j1RQw2XG6EEGwMpRx0i
Vb/EUZA6NGjcu4rsu/4zUUDpNuuA8mkLrQmoRONHz4tOgjRTf1m8bGoHmSjd
s/z34q+JJtXt2BuO5zWMEtBObOhbBTyfV1tVG23NRv3IdN1lAGC9EOPsGjDD
RLs2Yau0cjKimjPZ83VCqS4GWsmsOVVr3ptfGV0aAu01mIi6k8uJ/BtVCxY9
Dx3hett4d6IdvvktWULV6zHXlP4ECZ/Jhey3p3MFWMnGdlDiQV7wFDuIQhx1
xcZFTYM1scb2Y4sZN2hFkboukhzysv0YN2bx+wr86W7MBjK8fsuFNWVYDkFm
+wbU/EFOKv5uooW9OycNvBZIyyWICO7QWC3Ewm7r/c56YSJ5iFTEWqJMjP9n
0dERe03Gg1J9bCIhaC4OSpDQ+gdv9dZPrLJrAFHMrBA8l4+BMKn1ZVMJtOQJ
BQwy8Q/iwxIoFFYBIIyoYMHEndV6LvGjf2ufLjoXK6BRuZ252LMWhR7c3U0N
q2aL6qJ2YvMZY76zNhtLPhIhb5rzSOzXVOiFrxdJ4oc7NPgilAd6iRnIA5Md
hqaGqRsm357+DY9pMo3EO4SRanrlX+s+XBLyJbiZZMNM9EwvbrIT/JGkcPKx
PWdQLwiqGrnCy5APebtLkUDC4YIsBzX8uyHD9dlmGInbcZGqTiEyO5RYf2xy
Yh3GZ69qxRapn9v+41dgkoTyt6/BYzE5APBBkFk0DOH0tMDyCsZSvGgN6ZER
3mXyPDIbqVEfPp5wMCELl8JqtHEMJXSFFCmG566agNTtf6oJVl0oWeF3wQUg
wA8d8npZqmrv9n8zdEcMYltvVgi10h2cHwhp2kdcyjBrxf+Nf49F1J7F6L+m
dcX1m9yzx30KQqWpCNXqs5iXh6tlwMRLgX21G1X0kZplsrGn68JA6PnVyaWd
PfwVnixXEPSb8VTw63cqnXTwreSLf6sd7PJtuPwXUOvHGBgS9PLhiS9oIzNu
deXHlza7zPaOij7tSyDCvRhLGEzO2Du+MkP/M6xq4yRV4fkq/rn81cAJX1Jy
cP02gq/Relf0q1rNnBacfQCnWNLmjRB1BhgDAQRokbvItOXkPINIr6zpwCiK
RBO8uWNvOIqhOIrjhUe/J1UDZgZKKiqojMXrUrrCxUhWcanyxjSzGkIkTjUT
7ojYuvC9u7FsyOHG8Ux6LJniYJI/3fgT9aT7bGfWflh8u9kYksGSmADaixSO
tUD8vZssSXpgzYKioYyB0+GDQyytEp0boxE4b4BKmV/nlMHbypp9uN3JEQM+
W7+9RZ0dVWQYrx7GK7bWbb2oRIhFpvh+s1+OJL1yybH+AcdvqmhsfbJCVcJT
vIAlsLn9aGt7rZfcm64Q/l1mS2QVR89GXbJit64ysB7s/aXjj4zgticpMHZy
BMxXogdbj5Ve1RIc/F5YMhuGqBs5Zq+lg5V0KfzTsMkNxQ8jvvdOzwpiWGMH
4yJi0qe8Ks4VKYVYcDVfrUmWwEhyTqIAcCZrLemEoMKwMh3/X+IiGA8t5xb2
cKLywa0pxZCpWo+0RE7939zCGR8jczlmcMWJO6gkO8dxJeHb4g5vkfcW05hX
VbXvwrvnjHMV6AiaitgVlxuRX15I01rXTjLN76onDY3PtxLZ3FVtlpqfY+U3
2Z5x7k7wx+/RCDto9HP7BLBe5OTCpF9O4h4zBB1izY6cZTXpbOHeWWjBkQLL
tPbTY8j6PecUU8J/GoiiEdt+lsUYgDvt5DZovT/WAso4uJUEetZvs+TE2tff
TQvLh4XtOFkGAXU/bLY5y9OxpJolAY5NdFz6FCBNAGm31uq8WOT/my43HNIT
akKnGuhFPmTSUj2H2lPJyHjWgNzG7RiB+BihHxmeJol9kq7feWrunjpD9HR/
FvXT6EZvgxpzzBhlcUm/ulOZ42uv7i19s1qZoN7GfVYlP/5oMRacxC6Panu0
m7uJ2uJf7/qqjzhxkXDXoFCzDWXjKvXk+q24d1ZzvqbyLKC+2kOOeFwRcsQS
UGXfk882WWO+tMIgfHnjtDD3ukTn4Yev/UBKQgocKEcXyYZG1goLkO8HwMyt
/21nKOKRUs4LED3bqvuCYVCiHqWEk+IambnA80tiMCrqxwKMHi7T43MzjJAW
d/Utz00kcrPWFOx/Hj+183cy5tyD0AH+cN11ylhGCIHyP81mLQZuTetuHfAf
X2rffKZE/tPcdZ6SDHuSlIrYZJop9Uq0gcFIg46l41lzkjo77h8thPGsbSWQ
3hH6ySrZH/6oY+MTa/B4sW6oqjppUjpBHyFbqyilvukJ3aJQojDXIWEC7xDp
jOZWkzMu5VEn0Y7Aal5b0lt0bZFBWdQS6K4xkliVRQx36J0VpCLgFeaG87Xg
z+R/OlEgQzBOcGzuSlvkOTUYigCKj+xVazK2YRAqhObHzAaeiJl7BcJJ/0lK
4smylZj1wQdLLFZCzqWOBf2XmDA/ewr25pX/QK99lp0iBNKfg3DcENCZckDb
fEuKokpC3ryKWMt+tzkp/GRqS0VKX8u5aqOYg2JmGx84VPJqKe5LXso5heFd
W9Ja+DYzngJ/SnDKeYx0LF5ieoa8leW1RR9QyqMg7Fhatfs2mLpQ4aHykgVU
Ru665anIbEATdehhgX9b7QJy8ko7lALCHJmwl+6jyfMJdMc6uzlL52E0q1bc
XNJMdNhwjcjM5ZJJ8/+0LQWLOCmsiCYVs8XKHe3x/LzpCWz0Klpe4Xp9wy74
XBq44aXP2FLpUM/Zlmj4Tqr3hoxwklZ+Uw9v7EFKkbYxQBQyI3wfqOhF6CwM
O4FQh/1CDfKDmyVt4SaAHZ/LivWYWae6yOQGT/9ac53X2MrxtIHMjAwfHGyu
XR1mP8ymY3eYcbLQHoBf24jg8qZwScGn4FjL1s575Ilp77aN0PUpYlfwrD0m
RaRNGXUPwtbskAlOJRG7O6xx9wI50bcQPCJ9gaQZp9Ce+fJ1wgL9rOdLzjFY
zKWyHxXkj0MiZ7sPMas5DFD3T+GRXRSKKSJY47lMvmDMFc8K1WhPvbfIdA9s
KpYYx3oNWoc99SwrCGAViUZv8eiDRJk95ora6mI5teRc9DXI4G5SovBc+GfM
ntfyqyXPht2qkCeTllFDOo65TOLF9soFkf4+Kj3FucIE1ubKVveqvIOIiPIV
zNdoOYKlS4MiqgUpl7KsB7M8Kk4/qDZgjtzIQYbVWcYCQHGsemGpq1rF6ujb
8SK7CQ1Zx6m8Ysfj5RvKyFDWhu6tq4aZkVB7v6GdMSzitWZqTkt3LCGi9dMh
t+fRZUrQ+MXWqQVc1jIpNniDBc6iJK5+WE63iaetIf62USH3tWGpEuyiO6j9
+DFBF6O4Kz6YyQEkyXB1Z3oXKfDsSylsw49If3JRT+f+OEGHHafE+HFhYuA0
e2EUjp954zfql19y/r7cClv80a4tcdOyPQm9MAyQutRzDvbDSirU1+PX1f1F
JM0mhTB21PgA8t/PCopTXvI/TdSIvlNv1ZchJEsQyjKEkt5YrfzOoLsAWfbm
7CK4A8heJ1jlvKMbmr2ycNUVlRDJUFQfYXRCySLoatAWNimpHnUTPuVfc1j1
b+vtuPKmnjNe01bWDgo8AdX14PqL10RF7CCK153jjNQ2a7TOQeXH6R8s4fRk
l9RVJOxhj/TXhD0TanSjdSleBTl0hh1o60yk61XkeNgoyeJHO+of0uwMaaEQ
Rb7p7zBprGfo/nwfpEsV9YaYMyy6NmLPWI22kS4unVM+oothI4KZ/+U4cSJZ
5NzlD3kwxlLQo6T4+zJhAN/QguZ81BXnNqR49ULN+GfCOLLmcsQHYZcKdwrH
qqpufEU41zeCJnl2H3iuApvlSg0lrm0ip2i0FQh12vzMEE8oXkv6wOwNMW6c
m9gL7cONjs6qYXXSAv+7eVN5yx2giWDwZAQ8fC2a6EdQKuWc1KgxY8gaQ+ct
Bp1BoCLlKKILh85/AwJEzMd2H/ADU5d4fOQA/cHN4H5KgxMbZJl27sOlbSBh
24yunCRj4sHwTX7Hzn6SPl/mnctjRo63Ofa9Jr0iVXaaY8t+OzyqQGsvN+hO
ZDC/oS6/LuQUWF1HEM/N6laGtUo3EmusO53x0Yici1Kf56e1JCX+tB+G3c6X
eFo8UE1KWnPfxoXI4zZ9y7MG0Y1Q0y/wjfING+duVsE1D2mG+eHIz/atJRBm
HAZBodow19tJL9YQxIQ4NCC1rq4qdsj8mcQnoAwa8UfobdchHEafK93AFbrj
QPtE9KA+C5qgOf0GbPQl1Unib8SqgeWRV8VlRpKrGwb9yROlNFw6sakPJMLU
0E4ldOELXXVBPFSogDKv/rCVNkpl1xa1kxBmNph/mLfSE8Df9CQlYaq/nt5Q
bVnsF9pPKzCYBAJkg/qg9koNCNrydYr9BwOES/lsl2dmKRy5SpGBggbr/8Ph
fuf9uk6F0UX3qnUrv80RmXLW4pHsiDuFHkVotf0AhMjrbav3c6LIf8OLzblK
vDXqAthDZeemFzZWIslx/28B8G4qyQalJZPJBmmnk936fQN0rV0gEMRBPNmK
sxQRu/FyZ4PBu2w7AMlPkykL/nfiyLKpAS7zuE17xhx33ZOY2yLLIrzScm3+
wacg2PQt3VkYyPYQsula+2F3nkTHT+DYFinRuZn4wlA6Azsc6wZC0Szu6yHi
gHG9NStD8O17//q/hNswo7OTmrt300MRFRMTED1bOvFySO4CgR/Zho0vx73b
uJjK6Wda8Eid79kqAeczQO1HUG1W+NGRIGYHj6Cjs2aM7FrdNzmNvKMn/UX4
g0xGAcmZMs/Yd+gzxFmVzIiMIm5Uxhpm2Q0lbbi2Fe7sbWgXrXY2vE4NbwUU
S3z5iSooVprGjV3iCM9osB81utrCrm/fSWPQSy6tdQcOf8hWw+x38OEUr2ku
8yMd7INPTF0Ng8BOMtisqGtT/mJb3QUP6e8M4UioLdrD/jlbIbWSgwvDLV/3
GW8djlOjM8NRmyzwRh58qV1qIh8kUHANlXnBsOw2xWHyz0teIdBwlvTTKojw
uEDEAJ+q4BSvBPqGT+1448vvZUOalY22IXZkefrChwQwiat2T6Xy0eJcjVsP
CKZQ71eCReHFTin5y6jRX2dL718U0+mYlL88s9m+0VUuDfXMPKKY99x0DVs6
KsSkOYBz2EO7XBM9Wf0qi3VZ9HPvuZuxgWSeKRHOHrO3x8fK3xGAuSLzdU67
JX2aa9QLLWC2+rLPL5lmYdAj1CAJ3AfDfbgHeXiGFWdrFHiX/SMjPZp6lQYw
IOxzlLK4m7SRTAYWf94wFccEN1A3fUtgvdw2QYcELc6+Exn7CLz++nbyFI/2
0hIjhmsK5TolZgHeaLh9XzmjH/G/o5wFXkM8nKTZPJMdDA3fuS+wFFpK6/PP
62DhLxV30HbOqpjogltqHoo9G3SHdy/fmawsgBTLu23VM5yAPnB0kybQJrKt
eFwwuq2hlNZVhcjerE5Bm3mGJEtEYsIzmZ0lUS/M3q8hOsz2ISRGBC0cY+mT
ZIY3hU0/8aV2BKwLxnl7i83oQpGdw6v2v/DG3G5lfUMKz5fqd/tNxZhVs/7R
d21I3uyGO1IIDTkt47DR6nTaROzoF01IajvTtdlsGeuw9HksIKAaAmf0XsYo
WFhIDa9Uf8IczenwpXD+32TqaiXdAK1+K36TBsc9BpHccYqzOoKEeANU4XQZ
pYwyEKXrK4G2g25oTJd4cj4gdNqs0eqvDszGlH9NOZjxfcp+zhpDrC14XNSh
xQjC6NF94IlpWMcxnkqiBRdf15oGa00eY2eg1ItcXRzKjrMsdmMp/s06gKcz
rA5axAJyUcQ/Koh8CyiXMlr4wA0HDpwMaqYnXpYBEi+ht1YVI2FmWLixI1DX
fpvRU4y4Rgm/w0bAYKSOhBZcQL6VYwwOhXNdL6zZgzMEiaxoNLwhKvcwTfy5
70Xq3Wgfu5abB/3wC8/s9yBJH/lGkfgFKJNHYqLwSXGA/sWtp0sAuLDuebfW
PUd3Ka+Glyrgf8xSkw9xd5XwGa7Ac0c62S0NclBt/J7ZS0pk9XbpxC8WHgvY
JSVf/AD84wcxTCtMF6a+pWTlvj3q1gzuB9CRd+paE/GY1YebHjzfUmlI56sk
jE2Y/1OU9lWT1tA0M2MrNO8zvsne23grCW4Src+RCjWIX7HH1ADzdLoao9G5
KXVvvJ3aX0y0MX6PgJkxYzNs5WO5t7HYc7k93kw5ByeGJbxR1NshNTzqmVi8
DtkQzg1HhilMnmFq2AnV0tg/lRcxUabu6YggZ8/YPpnWhNi8sNC+73HGAY6B
wT1xh2I9+jLHLGwhtm6ra/7uVqM7kQdaefEevhvNctUjYbRVxeF6QAjZ80jS
OZp7/oYF5CwjrCGFdwVkcCvkzVdtFk0SOouH9xQeLiS5cJPxJolas1XIw9VG
Ii+bqQB3uYMAnKOuoUfId1YhZu994cinIEvknL9m09Gtt/PurnrAm8SVvD3q
/fs6sDUYDYuxT05RpVh4NnAr5u9WGa5GQE3UtFZTaQk8CuztoV8nXZV6lPD2
n+y6OATVpKPYPHjMt+zOsHRjQwtn8qMacFva7jIdU1vPnhmpPvlwl+/0TB1G
w8dd3m5oI77TR3lxcb4oevAGzXyXPD4VpIWtnxV5QqB0C8t9TKfcRhivMasz
sgC3d48b4bp1Ep6LSmgJtzikVixrvsZh7HNPjkHl5gsBaFaZ/xzBBF9qDk4g
UW0ic69AWJgYnaxLOqWCcH/8g7w/9lmgySgRhGgIc7nOVtAr2oKNo3b6dNbR
NPl0Uc68fhC99+FrFhcjUvOpFPXm6PnpkCls7iswQFi7o8VvsrH3Hd5gRXsJ
ysAKur9VKcN8S0u/CuM8QveeEz1sVytPVeMaRQqR4FfKBHurHUHxRrBdaehK
XDSzY3vYu2vnn6q6wsU1nbgLuWsYG/7kHIk7u/HJYrWsSrcDRAWsMF/3qZgI
3kHI3XASNwMILUXNhoa0I6FkT3lxNF6ZG4UseXlDI8EAySu2V1SaeJE3Xt1U
FOiXh/L0BP95elc6C9kdTyNr6B9/iz5TueIIv0ncCRINphS9eRv9nCeS6uUX
fYj0tfIz1nCjo8vTOI8+R40NgVNpNg0me94NgdhUsnX+9fA/zfAuoz73T7wJ
gFeV9tll+z+1mgka/vqRdUpGtvMcwOtsj4uOpYC+vfrbNQEoHkRhtmK9zK11
2GU9q1T/7omE34vI4QxhaM6YuDj2IcUCeWSnU9J8lRxxcv5i9W/v0fT81gdE
8C/ioyUcvkA5byxsuBuqpx3YyWMgFcMhIy2jrD6nHAa27Po2OGEIt8JpStJV
xLgpyVpIAXQWOeN8XFS5xsHFzWk//HAE0xRgd/yMJ+ivk6GXsLvtYsoPcIep
BlqdTSo2DmLE3LJIfHtekIN58BBObN12x1duxx2CcOGNnZfiagZHpo6PUAEG
DMAp15g0FFydlZpcKoDQpQrDSf10piuQBydSisRBzqVEqAlIk+p5HdQGo5in
2bcwZfptSuILcc3oC0PXLgTlqTLx6veEaGUGsmZnZw678zZMrUIuSBj2uicX
pdZnmtkBgGbxJyi73s+Fyqh2igCvkFE/qmBbGf8TSrQw8xekruZbQDCDYp7n
kX9rM4bSlK7aOWxhzOeHb6Uxc9eOuu9/Yp7cNlMNg5zWS9yjlfhG5TWk6ISo
HNDTlCio7qAkt3DfteH71uBNOtN9nebmBaVRkL6YY/dh0OtFL1RKrGZssF2c
VHN6ZHpqNApUT7JQ4rzzF0/QUK+hnGDO9S6ipeWRVOfkdfVgdQcR2Xrnhhfb
b/fz1cPh9eeiJSIt/dviivFujL3fgkx5JtyISUsXGfU7mR/mHlB8u9KKZnfb
QkpFmoROgeDPz/Anu+K5PdW7fj0fqqBzqha9hYPtarBzkXLH4DH8qjiEhR+o
ycjG5FedKTpWNJ6LCdecdm2KqMT8paFKjj32kvIjSTvRiZkwRNap/NyOZg77
mC0qK3ABcvEcE7Oh77i7aDi4Pwb5TwENVkco0Q9G7CCGQQfYJWJtBYoDAZlE
wtKif1iOXhlNFPHBIjCxrU/KEuYVOLBROMtF9t0E1zzGy3e1A2pV00+IAq9y
9W5Old4eFLV4SzlYDBiYeyR610B7Cpgc9ZXwA8yhAxWmCjEp502tP41Tx3fB
Ahz3f+TFUEB6l3YCYEXijSBKNCZ4uH3F6Db2uuYRxv9HKKd6gZOy/KEHjezX
9HuPRSJdon3pL+io2rEBQhGTKMuZCxVv64nkVfPQxFc95qe/0Z8EUqFqHW8v
/oY8C+pmvW/2D+VCkd8+F4XArCckdMSiQEm5HcjHJwDF0S8xido/26wjNgHC
RIIix4dVipTKhlOe+Hk30NNbFw+cdKzRto1Rzlvd/dO69Wd88jNAOVy1TdAp
4oc19gE3HgUm1Y9c44UXAv1z4Fpn+VWI6Efe1/LQGo9SRbvrKIZJSqt+hDDv
POZGmQThRL1X6BK7aeb9XjJw3DuoY2xNTklTnLiQLG56aocG69L1Ig/a+EWP
seSs6WtTDN7M0uAKxPWdnsQZa99CJzL+3/O7X5KxqdTNdm0siX21FlPQT6gf
Dol9NfI8iJdeL7/TE87ENrJqOHmsofTO4juu2FVUXVTJWrVcslu7Lywe79jv
tu6M2M5NVMa+iZRguqehdNxiHHnaG5+C6xZmV0bjJLN4bzCcHgFP/go6qJS2
QROks1ICiEveZk+Iq2KanI5jjOURXCJVBnuOFgSXJmAwGhQpiZpZXw3Wmahd
jH5605oV23uoGGrQ9WmqDwl70e2DGxm1zP+ucgmMfvct8I/A00OWXD1Ew41h
CNpDy3WQwbV9K+epbjkPc53+4ESY/5IuQ9/sKM2Au5tx47AmeU+fWjRlKaSp
v3tRYxLBYm4k+nqii6iRQZ6y0ZMD2HPgCWvcjWGxIhtyMzsLlE6RBj8TfvCT
GAwaliDCy8NPLTZmhiuv0mUah7jn6ges92nvMu31jp+KZ+N3YV5a9XPHeuoN
GFFW5QC7s0soV3nks75GVog8Hn4ZH2XXXyQrBSW5QeMIREjOWUEc3r0mKdkn
L5xx6IvAHUdZb60m6OIRKRVPasVvq3YRiEdthTeNr+rdKUypV1ym/Y696AKl
Y9gjNN+nkSx9tZu7RivDN9z9KR+cfzn2M4nuj07U2C17+xI6dVpg5BKVyz8p
tUikEHSq+Jj0sRHr6lL9/Yn0rRgghH1N3Iu9MrxVTZeiz6F0iGpzufFpC3Wv
E7nMk9NyL+QZU3P71xHLIu6eQxNZxK3RJRvtcWeUDbhrIz+xc0b9kt6gbyjo
cKOrFJmiUhZZk5zu5rrdewSLzVF66l90Dcazj1a98oOnEx63zT0yPeG7C3fU
U9+UxvKjGZhECBPdQN77tJApzBbbhdHbRcCiYVeWh17IFoWCl/TgY5+H0vU7
mnD1QpzV35X4WR+nh6NUkC7bIVzY0g/VmLgZRbyZP0h6B3V33DGy6jezq/qe
C4ValjPaznyBRHYcKkEp+p9U8+M2spbo8jBWnqn9BpSz8lfZzxPRovh7Z4hk
ThSR3Oyiz2JXX/DfpkzT8OEQmhuJyn7VM76YdzFup+PGg1wHiMpDkQBQDxUA
h2L9aPppc+54DMibq4h5bdI3D3jE1PurR49pPHzuaBMnHr9huhugpPoHKmhJ
SEcHmelSReLH4YfVeeqEH6CEjel1WAx7eWhubsn9UP/zGQ1hFHqa6J1rTDv8
1p5FwqlDev0OTWEdYSaZP/VP7Ab32o/YPjsnMJSZtl1VmSM32CqcjNgznxNG
W6WhMZakWt4B0iOGWZPfgAyLd7xafHoMzFMqJMklCv55eot5H7ruG2URFcda
anU9MXQThf0uS2GWFy2GqU8zkGPng0NKlfbuwIZWXP0w7zlE3Q91kGvIDBJg
cbWXM21EVOW71sFWuzM4QJnbz6RKxGNec6+6ajWXejdLxdiUXdNp27eV0G3E
PvvGvLDWv9AP3N5mLvFo/AaUx2xwVa1sB3XG3myRuBZJmty6tEj84Bps3RBw
kcJYI9P4BNzEUqM8GAlDENU3E5W+E8KhlGgC/X/N5VWPrtkWVWCIqW7TVehd
I32eB8wrjImUPyZ+29c6d2U/YxrJnyXu239JoNo6YLxU0dE9bGxMNzLlejWb
QGU/ejiol7N+Ix5Vw/Lphb3KGSrymHJWzgQt/ts86KWzEjKr6RS8K2wfDTtt
u2L3mepshy0G1eG/Zzn6lpZbDUezRpUF+aXm+/tJP3xntXvEKXL5dVTNc3+Y
oOgoGPvhGmKj3zsDHXbS71h/0QlN6eS/eP1HBRI6XqYLrhRZfl088+DIhg3V
44UamLej7FKHMVuoKWflNAN/9SN0FzrvKv0hd1GIAaDm3EdTB7gMu9t006/D
VfGAKFfVNrw378DQ8Ua91HgL8UEwnz1JLK2hpcixorXRIfumzkx5uj91dnqo
9nxM6pflkmIkhindH+jGuNMl7n0p0PtdgwHnltV06C1R1qw9h6Dw03LEUsI9
Eei8nRh6lXM27q16P8zGj33xmdXsV9uhrYlM8sXHJ7EtRhFNf2ApYcMR4ssD
FhufJjFzH5JrcdzcxRlclJe3uFOeKAsyv77NIFf2ydH+FCkh47bnWAgGY+4l
w7o6bMQA75lD8rLViUZHmXDcBFZmBulomRpGsMK9KuvRa46XLgs9Rt/5Kb+g
jbvMy4NZQiRGU/frTI6/zwB+NkqdrGPgGSYCI/R3zCW24BbC+u1MTVVUSUXM
o1MW1ZtGerU2xKyTvdot

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "sTlVzHE+yhAN9Vt4a+7yJC9Gw9bfBRq6xv9kCe7Ng5psJnHruz9VrHCdetev/ZiPTJdBJQmffKsGhcT8C1xHmtnWp2phLrsA++mCi6ZvsisBHsXsEe07/2w+B8eMNZubT3xnRLX8hyEfcYoWZpsP3M1DFemdUhSKGBtblrC5P70SnbNX6tsPF3y1BZk1iC/CtfkXVJdvvd+neDISHf8HMgQ3zyVqVVLAWr5Qxk5Q0qRqkN5ji6TFlckAsiRmO11wQdJiRm4jh+7cBW/zJeXUl6OMqcwyEZMuU/29oQjg2A1J/hznazFDhyqwQe38GdRgNUBHo6CHqurGPChrl4jMRopOuGFs85nGZnQ3Pln6vnDWXsjpJvnd60IHUW6VO/Gn1SxhUpiRVSv1T2JIO1QqaraIfCeVgMJprVoL1jW41pZPWG6vZeg02AEm2oSOaG5uirxaOoYZ40pRAlXYTdq5vsq7kX5J0d9oky/24zGxcdVMBx06q15JADNL/E6eDxJcLmUh/xvkqAOAIOUfM1gtak7sbwKoy94wkD838iSyg7nk86qYIaF9EEGKFcTYukwZYy6+rtO1HRAAjYy0fPkDHQBXE1V72Bg/Evd2ObTmmxpL9BzKgBQinRrTwSDBUgsE2+01O2RHaRaH/Y92xvocFGmQpiahdL7B/iD69g4s/DPaeQs4h8/SCGo7z8Mh1cVutV9+RlPJVMdeAgYV9Zr0TpUKkcvIUkhAUzDT/ei7Pi78LCCxylgZLsAbIQTGN57wmAiUvz4SKLP+q/IdXV49hbWbCACEXUng/UVJqdvKNVhY92uaeo8hok16+5/oYD6aUt2mnxCkc4cVBQvJwm11WobgBdcdKNa9RtwjmNVucWvwaF2z/Mw+vlJJ2SIJ3QqR8q52faN4KbQ7BKi9TQRuUH7sIEr0z1LV9zniJ8+EeVN8qG1AKYUd56maERVY0Zf2MKYBPmXWQstG/+y/JTSz33oFJ7E2ztc9da0cxrBYXXisJvaWowcy/arqy0XKCdgc"
`endif