// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GzJ2Wjs26K9pOSJmCjrb0jAj+N3D02bK/H/gUo6NSTsdtoABra7T9OPOSETe
8uj6lA+1gfnet9cqhorzk5MuY0b1JkhOR4AI8ZF/QLqy2dDdj+ycnFSM3IVr
lJIq3MTbSVaXwrZkHK9AJ/VFwD2TdA3duz5yKD5JALWdrK0YnyDLJxeeKlIZ
3fu/0M/Rqd+tz5dcLRD74OlLFvYuG3hVR5z54dQsSWa8ihScNBzoTUKyNtu7
nOFMDgLkwYu1njYABT0LfRWqv9FNsZKoGOWUup6eqbrxTI/jxwTYRK+917vM
q3J2EV00D94PgtDmr65KwWpK9NtQxY6EkYKrOrzI8g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bUWNKYUV/823E1UhMllfBZacVPoi1UIKQGOo4aa0IzaX7visL6OuPZhSQmFW
jgnSeXlye0uqeJhiX8ZHLlOYZD6wTQDejTLp/+OrDrzJiALaa1VGy9punwmD
65ChH3rEnypqEnIVgFOGJttpXZZJkEUnfAEq8wJWUtECqTzpKDqpeNUGkbbO
STBoMl0csHS4gpTB5g49ugONya8f1fCUHktiLQ5lrb3/8TWn97MYWX3jyMYO
gjyDKw7zsuI4GBqTG4U1NeZP3p1Vx45fY2vV4pBe/KpNXrXXvbxHazR65qrX
D5YXAEOYzkEIMDnJANkFF4d+9+9Fhpg59vt+wcspMQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
e1Bq4/nR0Qf/Z+KxgJboqqt/5f7vMSgdyvbDGvNyK4NzUgOa23eBgR+SWyTc
CMuVFETic4oea8doVeKXz0+aMCuidLRe+an3VximS0zXqEa5JPXzZ/P3n7bw
c4xQBX675+Kveu7pSGkB06GU7JffdvJ2wODoTfqbxO0TMcRXWJ5P67veJ629
5Wk3JtJ3ZbmNV/kMwZdhRVC2wpbLRsmxow9Msmon9qrW0opjTZJ+3y575ewX
6Mh7l4D9F3+SxbnZsvzBPpq32MHgH66hcQwYbX1FqWlsDAdn6h0LGY2YwOFy
/YzHMmSbSb8tOqfdgC8uG5xa4IOKMv1LQ1KQdl/7DQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Bdq006g5WT0zUyLGmv5TRNBr0dMUHZofHYb2fW6aNtoROhmMKKoQ+rZYZ149
1YvIRoLcyD0gvhyxBmV8S5+5FPomk9Jch2VTOkXpEo+Yz7fEeFB6wKu0i9M6
GsGJKxvnXAh0WRvJIiwApDdt8G52mRnHPa5o6fef67s0XDjhJG9dgTl+x1fa
HwbhqKy44xiy8gzmooCCocvqsnn9IYhZfEBB4JsdbcfvYlUjqf8r2lX41kjP
ye2zlW5fKLSDxu/8HWv1QH86roz5/wFvS2prssNbpHatzP6S7qaBfzMKsngu
NHgBSN5d2pFXgFsRJxY2HwumsC5ReC5jkrQv4JciEQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
J9VoY9UggvDeXK6/mPMGeLiitHLOv5M69X3OxqKHvNN0gl243BZ9E5GVyzqv
nR6Msk5PQQnkD80o5wGNiZB0NP67/TfOJ3si9ZlEauq1o8XLFTKLf9Z6WD3Y
Gz1V3k4exiNNk/BRU/GlUu/2+d6uW3vu2toGjc4Pnnee8zojfYo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
FVJ9GDpu8sH1rHGE9SiS/4+VyOAt9IGAqLrQPDAmsLxSvGpX+kQeqJ5qfkVL
/Cf8Yw1oepYMVq/dWE6VgX7iuzf5EPWFCh8M12yj+MYk1NRUbl2xHpBnzGFK
y90XZpOhkS+X4e/HZwpBzUm4z/+kVISZ90pW8hnQpTODVIS68v4kKPzalq6K
0GQmDu8SYEjILiUvglN54zBY4GNS45lstOZKEMkZsb5hc4ioP8578sPlw/XO
Hxfaw6FTPDoFHdAxhnKDpZg1kokbTTK/oPdacYCUKzNSt95PI/1m1EoKKLdu
cqTMFDD9edXHDiOkj1Gv5Y9KkPNjF1Vdt5/mwDcW2iRxRNvE+8UoEiSvs0QO
oXRNU85EKkQS6OgdOa3L3HS8SSHhbp3B9zGNjwh3R0Rp1VkqMvFSqeSrMGIa
MX7PWyzknMgpQ96OxEkX/j4FJhzX6/ZNlO3vjhjnyRGoFzea9dtn55MzX64x
Ir0XgsqW3kA0SlWFCN/ewnUNpzdDZaxu


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HPA+Smng/MZsG25T8ZlqEoXwSaZaUlrYKbpmSE6HZvYe/pQlWJleR+83B/Ur
r+GVfd365FtCrPjGWp8mQJuheVY4ViaEiCPvDHbdFPzJ0Q/EaVkKmLQsesmC
SZhdnLxU86RR8zIfLMAEoh1J9b786F3aqa+tYLKr+armjWveeGI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MSso3H4hfq2iwGfJqzcw/Hk/Mp4ag7+LreabL3+sST5YeBKhxhSNkDsXUYiH
Da5Mv9h3zPDXv6x+255/iUf+ajvPt0wGWAAJ7TeT242LNqMpeEQW1kIKcChJ
DhV8lXOfdiCWoOF0I3Ife760x4rMjY6IBYYL3dAAZKOqFF6F864=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 91264)
`pragma protect data_block
ZrBBsCM4Yol0QDplq557LUfznnCSuFpm+fgU8RSanvRdaJGH/KHDGv6hUC/6
cxcTl1AQmIi6WNCmcBZkbKcVtY0hwhAMSmwVnjnqUKQSsY6EXDe1Lcp8tWjX
gCdvSvJLynv7+YRVd8F/jI/ZOtyIvg96jcVb9ebG2fYnDQ3tf2/6ZAqztNNE
qQ/liHQZTwjlPAfHz1F9uzd9ve7vfAvmAdayR6i9wo0lBjP9sOv20cnHuKb3
3RfCzGwx60ItdXpro+PtAsYzMrtX0mHE8M4JhKq7aGsaMV3Qhjz1Fioy4Zja
lOWg8Krk4qG+O+0CkcxEMRayYwlNhojtaQlVFzHti8P/9Lx2F7KI6Q6f2Q83
x2xbZFJu1bnayLbb0T6pCOSqFVGXs/rUoUpTwMEypKLG3mxtEqdzhT88KHME
7xooPL61+aru+sgYm/v5kh4Wv5I0C7MITGSvtZFJ6x/9O05blwiQAAjeqq4l
noDpxMdVbZaEFUNX3Pn9b4ByewvIiU+o7gCh85EJnQ4U7yqc7q9Pi82/4T1p
V9hcQn9K4NiAIosKXdtrtOytOpSo6fYlHRycLoywLS5RHvVKxAMgyUDVQcYs
i1+6cHpiSjKqDh0goqd/J25SZ5DCVp27EqgNxYqD8xnypM88S/t6oj8kHgIA
0t07HA6/RAwctkWNBt4Gtx7r0P2C95r0MUqiE53gFU1Ijxj4zr780wRcUATl
QaE9JUJQMdB5Y5giqY7BZSydWeLxBwNF9NN2qOHf1KTXVieLAHJZg9HaZLs6
ijJg4uqcdwy1gfWf/BeRHCH74XXT8H6eI7bJvCr5cOuLLK457PXDuG/3cnRh
qtta2VHrthY8zab0IfTTPzCbKJDR3gIHEmuhekLCUDfIuvXmuGZHpsLsU9DG
cWTIgymOTPnYB3WI76P/gb56GLXcszrX1Z2jFx3CFeG4GLGUqd4MeQ+vt2c9
PjZurZjcv/EMRn+nPmYbyZX16MH75PxUTBqCn76cg14h4aHK2BM1NztXw4I/
JRoAE+1EYmMJu9zzPIDCDIj0pYKTQGplb8S4r61KehvyeA8hhFMLnY31nzHj
5R2X3UUOuMhOMuEz9JdJjlnrDH864dia6aO+gcRWl40Ltgnu3XNaLKCSqVk8
IR7v+O0gbmofPX0EEGUz27neKfaDnfA7DRzvlEzW7fPhXELXHmMT3sATQ2jG
2RBuJm2ZD4TanoeUSi9/5xIrs/56OpgBs0+FtpZWA0r7s5GZ9K+6dmggtQOu
l+K9isAz2/0+ID7pWeAJf99u7tBj7sPa4tCZHTIcEGhhcl9PuRJ+1LSOcbpx
hEdu3a+bpfehL2OLGTdEzpnlkEDG4aDbgf5Lyw4jRwdTRSyaOF5GLxsvUt60
n92Zf9xo2QKq6un5nqqrhSomcT5aFJZamwr9R9NqiuLwE0i4idP71g+K83L+
cdYkdcCPnABXhLmai2+7S3jZfyrnYRju5WvSQrekyaop+x3quWLAOfuGLHzP
fHWkNE/1EjSa5s7zy0HObTyflc1mKSy/kn7PBDkOO0vjQ7V6WE2lTDuVKs9C
rbrvAdwjCDnzLIL4OGo2XrhdHlr/ffnw8K92hkKz5IufrLvQepOMxpKFuTyl
SyoN7Q+Sd3XDhuPX9CstPivzRcYy1NTiqqRr7YFzGJt/GtPETPWSOBmlONcv
/2Y+iuMM9Z+xGedXN36FjDneqSq+16x6Iu0FrKok+A9/qKkZTFRy1YvjfhJB
bpT/PqNwCyZNAbaSXu6hdheiDkQ/hRcNHFFCnPVp00VKeGCksry+novuOd16
uosoa5wTniWtjxQKTKkcxWrh6FzzFJReH1o9LUELIuLs6bMkJvsm7tGpggVB
WhxyuAz+NK1HwSANTGlVVCPaY/BVY5J8+6a1LtAZBbQSynlC0vHmnJn/VNNb
PyS2414x/Lp9dduuW6lMmkGd9pdf3i6W8LQtxdtvd6SkWBxi1KxNkwIoqpbH
6w59Ya7viy2a/rb5ASpTcwKTDSkdc+awVMAbTUuyegBWhY1vRqRp6J8pWEqh
pLpeP9RKoOeSGtq3Y1dr34igm/T3W8lpmFhR9NwUx8znsnd/Rj5KKdf0rEao
B8p/kSXXQB+ZbUO2ezOxxSCxQfkFiNyHi+WfqJ0GJV29cab+SjnwPvdBEpDS
LYFcLnh1icS0fKT+U05fWze7shAGcDC9yww6K8lpJWRcaRBVSHyUFV6sEF58
xdJ6AH1CEgLDVGj/teicU2Vg6P2K/bdGAAB1bZ5tzX/guWqrZt9/BhDNuSBb
4/V4xSNykd/xwjwYIogqNjQcoUiB4R9sQdZTqgZxx5AAKQRijvgekgd3d5Wf
oiVPuJlnxQI1QS55OJM05Ozg9aebveIvqA7Fe+IV4a9Mf1ymn/AJSvz4uZVB
UjLE3WyCNT+GFeDK1R4+JpuNNKEtn6gb/Ud4N6GjlPpIp1zhWquJq8sKeqf4
1LqsbnemYr7eVjNlXOVBK0/b1IKEeUQfMds/UMG7mYQariJxT3zSLL172lhw
5PGDJ1Z5dWoe7UOtEValnrqjIv71ghucXQJT+a48DHNNx0yrCmCctZ2BD4oC
qd/OJyn9XnyKxQF96JYCvwKzoLsmKA/eIBTc4ACqn4r3w9QZZbKosQ556dik
A8S62Tes6jjNyuEi/IGnTrn+x8Wqjmj/ZtjO96rRe1RXVHf5SLOD6cAKtic5
ZNxxeqMmIrRTzCFIsaQc4nMDwzqBhGicuAAFaMOi7L0pmLEwL6rMEQJn3KUd
3igew7PuEi/+EI1vZS89wD8yUUkmWsb4ThdcwYHEKqCoebsOFHypy0nvnxmQ
wL+dloeKtG5EuyV0vqrX2Bzjjc/R26Qlgwh7/G/Qgky4/YETpLAh1xRqJ1UM
WGtN38PXJnE1u54gxApcqYK7PCdGiLqLc2PZ8zzWNDlcmgyuAN8uYGHObBPQ
qtzIaefHrs+30kDIKgTbcip92l67ibHSCNy2BhdV7MKI775tWq/1IJ6hWh2s
6hifQhujlEbMGNFd2/O8ubcwQy4b/JIVW3fTYLNyYNFYfhMS+A9ZiC6B5UFq
Fo/tUeSgG9z958hnKwqnIzmlWrLwKy5SamDIkDSUxnlt0EmIC9ZBwuyr3zWe
bS5r9ECs8uxrOZsIbDEBHhkPV0QWN/fMqbCU6osoFbdU1JuYr+97/1qji4bs
Blg/jHE7OJghDYVXCRmzPizaiyBmp4AkNzpASC0kpBIRduxk9B1XZ4CARQ/Y
6EP9V8/DeZTBZARilbvs/qsG/7NpvhJdSI9YsX4XCwhbVBbbvwKTUur0QSsT
837aMxE2awYXUGcH9eN0Vp6lfrzhQkocL9a9evfYc8eyWbhLuryO4Gj2Iis8
5ZrY/YFkjYd8ZMd9OC+q+cPrgpszGMMG+ztTjiEwzatNmGpd8DeMXskqZ7of
y49b8P2rXYXpd5ysBF4X+8tl9IbX4Xc8jT0/7cxNXg524cj8zlGLFF+k5KIY
GU7ZqNspVpUdq1OB8thOT/10LqN7z7XxWCT+JN1L6vjbd/9cGWuP/PEVhZdD
F1Jt/euGnikD5etYJKG9el6B0OdiXiqA73WdRgN75bXRLhH2FpNEwewMuE3K
ffBF7IGGa9YY9YFR2lZMHAWpmP+jSdTLBw13HIEzNiSo+w4+ykv2kHYF2Zw+
LrFHHRY/ASsMnlX7QyFyCameJNHFBToBFB4yqyf29y5QJ11vd2ey6x/ovnK4
+kOPeW4V0/tfT183DXGZvy6/bU+XhAjelr6pfb+oaMOcXsZy2jqn1PkiLXgb
CZEJW0W9D8OeRBfPKp0tVGlyixR0KgTN7QwLjG1cZ0MHNQHfMljzhrhJSxJd
IsMp/tIXBY6HOX6scO5Ez5lxq0NT7Zmw1qtgCEHgPN5rsqaZQZITC9sCbPpV
aKsneneRjbxSgolIArz/8tAKb3Y6sTB6Vym8NAK8ifo9TaL1HwGEckpJdpue
9I+e6nieHAtikwhNGGbT7LiP+sPYszxxQn7YlmRxwq3R+pRDmzWpjy9IMQlu
ZnXJZ13X0Rj7iB+Qxaon5xBeqkamMZuS5F5K2Nifv7Lqxp5nGfVZmnw2DXzI
B5EmvPdwkuJH2ymO+KfuKTP2VakMHNxU2BPdyCrYwOpOS82XF2rEDoGRSxTf
LfVUZ7DOHOpT9up+bb1YfLOyieF+3C2AOY/yYrC0WOwUgHdMBHyum6FreXqf
NPzbo/8bfKCqYDNFZzpJnfU1+Tsg6enU6U5KXQ3buAEp3KXkmD9vekb1LytQ
Uh/pZ9JhlcR83gdhyfkji+7dy/Zj3kjeWHzg07ssa3UEtV+p8bKsEmEUdCu2
487cnM3Be0ewPRwWH47eFLMJVPSkLgbHtrQ1gjIY3f9BsOSXWqRG/sM4KPYV
s+ujCXUOLe+HdM/HqJs/M6dYko8BD6numX/vwqEcEMOcijP5MeGFYXNLg3i3
nEQ8f0+DpguooSl6WuKp88knbg7CW52EmVQQrNTNHlDsd8JQGjbttuT0NHml
6JkrrLXb2O64aDPWGD6RJPfk92VYaKpr+8GYftNoXjBCaVlzMmr6jsECZ6Tm
jJyhT2vbHG2hfrFrLpAvxEdpFlqmD76QSnCgliN/mymKmtgcEgyUorZ6Msol
H0gZLqVWTkQKeE7DjRcKgJ6HnkNXR1KkEcPf0vDBDslX3SbHcfhyGvPEu5Di
dsw7ENFyDvVtCQMC5uwlkfAefNjt4Vwhl2uYfeZqzQ3kOW77iloWBR1/y/jP
Azz1H/9iCCk60ETZgV0HbeIGjZaiIqndCIXzHLpJT1xIL4KZgJE8MJfoWKsn
Gnf6q49OLpaZ9uNtHl0yFCORlIRc9iJD8ZLsVDWwDmHzCSS4YSfpp2TK47P3
gaUNsfbi3XQ0jKQl7lWHSx4SWAlbtgrsv2uA7+5OI6Ol0lJ296B2BzJqj6wd
ckJmNuHKhiDlbS0SuO7sxrx+0wAQdKkbPVqRADN5hcgjtvsQOGcruPn0lkTS
4C1KRkMdhbodTXqsdHDc5TyhIIWO7FQhbsP4RByPdX4Q7I5UyhzzhPDBcQMB
yYlm+VRjp2RvLoNXluzXlcPd9cobt/0MFclagvcNgtqfGl4kBh1gFU1m3ZeC
nqc7lY2Hx4lyGfZpnaRE8EzKH/Z4WeQsHnRKMAIbmNjJjMoMa+CFnwLefy0F
aigNoRnnGdex4yfCz7mOcB6hNWea6lw/pV+ZV+P4IbjqLzBVD25HKN33fPgB
fzQriLNYavPEI8HpJt3naCcvcxuJ2aWG472SrN5+SbhTaZcprgG27s41JHll
VFmDKuYxKJgdl0tkCo+hrAT4MXKXu58f2h1jOYyBA/MRDcDYDa7TtTFpp14F
Y9h54waGFXgCJN2GiyGxU20f0M5Z487L3LYp7nC6JpY7rpkJ4/2L3TCsxgZG
RkEEkBMxVGQBAtRRXdLmO05jJ7S0RhZ6erMKcsxlRH9afCSRivZm1ChJC21x
HgXfLwSrMRtYG6veEr3a488XuGtEZfelS6MJCzTEQnrWp7o5wcRGrJrJqON7
WXo6jridF7XCOL8bRDkMFQa2MRzk1LcBkBjci0lEmrSVioC+ojLxXJt0rlJP
swFgNebetRdTH2Evozdk4JtGUNF2UoJ13eG2nT1PS5YMnwMfl6ito75tRgeE
xnNXNYvKzhi/A2+4t7UWVYTv0c7j7mBPx/2DoN3yCbfe3hU44QPjTvY0d73f
XNMR6cReCx3EJjp6ZPt5WvAygH3nCUaOaBBYyKZyN+MSGhBbvflOS6Ev+YDK
UYpGTYw97mQlCWBHDVm/zoNq/vBUMkIm/B9Tt/wRmvtacsaSVPNtXQLD1aHE
NDGEActmSLevZTVCA+CgzYYeVm8wkhBBdxj2ZJw+t/e7AaLimiyRxRhDXD04
1Gd/yyLVrxiju+/HUcz/lPDqrM63Ns6zcXApE8WPNQ5LJTBg4QPhrbiKLkCt
dPUQklVUNvvQvm64gIiWgrLhecwDLxwlPuM2KoUqUStOVOPUGqx+ys4Qpsdl
8pLcvHUPxHkrLKhZe/Bxy86hOPsfbCzy68vzmkA5d100pWOK6eRSX+wjqDlU
/mrkPz71Wuz3OtojZ9eyu0YPrjNEThRIW9qdFFAS8rt/pE7bNuvtVv0qjVIi
dqu1u32SXUr2c00Z/OUfeHQN6LZGQM2EC8MbuXvSxU9hdHHfQBXwHVsghMw1
EKrivJOC0tyxKa/tSQL/iKrKXmuz0cce9hGZWG2aU+nyDFqhxMEya7s4x2xr
niNa/bJX/+/9NWURm+9z43BF4D1AVF6WiegnSewg7GbXFfJ+CUpDRZgrQ8wH
Ye2SPU5NCYHadZKSbBgI8yqaAHGE07Te6wZXwFILm6oUrY/PBV4cXjjGehK6
YicLTeHncVYyNzyqKTIqagT5cFq+s0fDEZweHb7kljMTtSFH7xLW4ddqRr79
7+LcifFFv4QFHNrF3Mfu0v8FhVGh6XpKlBxGrB4xIMjYysFtqz4w+DeuZuJB
1/KKeBXvOywwpIgjUg/cxWQkh0556wiv7OoIxXdFs1CkST3RjJjhj+5rXXZv
YNh6WIrn9n+5KcNPryhsaLFAHx/YdeM2uq48Nirsevw6v3z2pO1axl8H6M3z
TQYFYgA66n0dzWe6LGBBRQeSqLlyo36qianLXTu5zFz34F2d7N6KWgLiEtgb
Trizfa66bN2hcXgEMP1+Y0ZrF7ws4dgL+K4CyYOD9n33E86BZ8gKizIBofdo
T3LjsulBrsoAkQLMC0zFsBpDXsaAHFdPqUPxvfzVc/L1HMj8FPUIeLCtnmKI
IXGeOMX8Ad/UE2ZLO95ixGTp1oNz0S+dVa+lXAS9t6Qla6uo3oRedLUYHokh
/+K1QvVQdaj0kB7NFzpWkoTSPNr5hvImdyQfYbBpb07/sxbJWf5u3B31rsAs
OipZ7LQWq06PsMoft/wC6j0je4imxn94gNZBKtH131BZviy6otCFsNH+qo9A
ZKTAi8hQGX3/R8WUGIM3nolEBvZ/YKnfzputKByGkDZ0z0mcCWDTwtVT4RZ4
p5f535NO0c8CgsreBk3Wobii+WwXBsRfYY6cVJlxgvxm4rWP96IXVkf+H9ul
DindOliU54oT9bHn6pCesl+SwYkZ07MKIUTtpcSBdhI0soEjPn3HG6uv2KqD
9xO0uLB7EJiJMrn9Fq05hbJNQpxsZqk+50qcBEylJPheoFf1vClMmVCsZRUr
Z6VfAjhOBAeLyzCLZlkwyKHwLV5VQ0RGX3H846OOi1skLyToQ8FUjXjZKsH0
g16B6bRkHrCkKXeI6YiTWilzQsfB433AlUDbySORy2xHwPadneVdTgIv+nvv
5V81k78g2XnwrZS4T/IfflRj5ADpXzy96N8jRjgi7TzfaVpDLtiDoGOPNaMY
z+xs4HQgKp4L6CHMV8ZSJDj9PdjtLnr9FhMie+KZaKcygjbaNDFjENaN870z
o4iiBv8Gi0+pLeO45ZRlODxIy0q5YOL+hAP1QOId5PFL9k2ZSplDFECU8Cg4
0Xgu56WJTpHdJSOatOrrvn3sL1xNvEOdrzc3fxvrsqNiZXgKCiwD1QcMwDe3
BGM+YwIDfUR5MKPG8uknXWPJgt45xHwUoJI6YB7Whxj7QkYaWZZVHJoKQA70
ceghSdC7mHYxjACz+PUMnt0Yaks6tbbgzMrJcFR3yuV/eoyWaCJ7VEPRg5Vq
d8W4fn7PDyo9kT0BhkVPHmmgk8rYQ1ylV0fsIzxb8pGFTPO0rVldVaJnLsdl
8nY0ZusbgOuy/d3DlVMyWwdfmHpmP26Blfh2AB2woldJb8tj3il2iFo4dCJ+
X1VYFel6GDhg6Vd8fANupku8XLGFn8jd+pndCkbTA76HO/L4DdO5tnmNVEtR
GSvLUTbqDfsqT+ASe4iqvoeq0FgwmmcKqyDnnQY4av1D6fYCxNOBqaGfE14X
BINIvDBk4eY1XCzZS4uHbE5ttIJxvwSnTwT3vnaO5wBbmRL69VzSw5CpvDhe
HnBT8IffPWeVTWILtPvCGDBGBXyAgHYBG+wokllH4Y5qiPZi3Ixn44VTKNFz
2nqXDiPUnqM+7BKqpnubdgvo0qNp1+CqMNDxTMi/uPbK4+16gV/HjnlIa6nJ
wwxOUTB9KBo0WlQAgVtFm74xoYUH6gIFnf4gu7M8oLeLAo/TJAeKIABZqzfj
I6cpL8l1DkmsoLzHYIJFjsbBdyUM9tzzt57SDwDxYYSaV1DtHnRq1QfZvdcU
68xDOeKQ0fMXS9It5Ravwi8kehn0WTCWetSkh30+gnTsVwUvPefdRkvQcFVl
BXqq2YEFtCOWumtyOOU+cq1KURGI9xBbMVfkDoQapS/B8Vu8pduZoz+cQuRM
9brmlf/8+tmUZWgWdjde/LyTetVNfyZ9jJV6fGgp8R85K4bVG+DxfGo7BO1s
ErzOBH9c2krlrIiOWF8IKZq3/1f9Srh6Cz1DV4jVf2Ce++YpAnTohWyC3wB+
8FzorJHp6vICkhtIydzmOsYD8MtrUW/DYU9gqUiL3m8y2tbKJfKyLjearm4K
uQQicNRjHTzaaaN/61uzKCFJPPh038U8AvYQRB1y5cVP+lLXorlk6Lwu8Ye8
bMeKa0e398YPtXR3cjfJZJ25Rd2la2LnkhpH1ikAsqq7gfove+RGAUkEdHo5
VQvb1rGsdlIShuoSfotPGXw4C3cA6blZNju6B43pP1j6YGzWDHxWYVZyk9W8
RZK0mUz50JI7Ft1zpM7EZLYXdwBA8Di37IQVfiztUO0u58du6U/RPcTdIzDt
bZmR2yL5C7J2qa+VQaX9uVyCm3U+aR6NAK6PCGIaTjWl9PjlrMF8OjsoBDnR
QMq0qtltBX6NSgi9rhFaLD27eyOAa1/k0y6aIVD2YpDThkK8GLE8urFaAva5
shNni4LO5PD+ZJIttmoGxrW+6g/iUvXkY/sl9sqM/oUcNtAQmy7lZApCHyEU
/0CBhW+1TPTkcR9WzeL43jZlc0spzElTsFqn7FEx6LWV8qbE9eeiVkHsMu3K
1Ms6GqpqiyJCxRdVoNoSPSUmaRYiPdbmmenBnOqzHAT6rhx2J4bjUJXZlRlq
J060JvaQPqa9c18Gv3auZJEx5TKji07PN95Cl1nAy73KcWcCLK+ewSAtw47Q
OfLQwLE8te/rOoBySQqFIpvk2JdxNDWsIXL+atEejiGygIUI+YBxkPs8APuC
aEZEinuHqoQld4TFdu8NjWmpHMudx1ntGPx95M5R54N1mcR6sa6fpczav8SJ
v3EZOIrs0TUk+Fsr3Izdk1x3KxqxhaVg1XhJNXZNcyeDpzQp28WXeLQVx+Jp
a+mbrgl/m+xXsxt2iSG1Nl5eSIHlYV8AvIKyj+DH3FfDjPge6hCaqEy5JpZo
dIcOtak00Ff+lZz3HGKyUrK7GwUeXZtOeK1tm0LBXutDxEATwdjjLwqOdzuB
AEwE9mYfQdH2GYiO6AvgfIcjWvUX136l9s3vX7jks0LxKLxvJ3KhwRBwrDF0
GmU85360DXUa+aTM84PB07+D3HQ2BlX+hyeZT3cZ6PghsHsR72JjWdTW0USA
4RSlXUW4MWthBs+ueVkc/ZilHfigOmF73rQ1gPyA5149U7OTCECZDKC2oLax
Gso74SS3uiDoiHfWA4p1aMDPwVY7Y+YWZncfdNfV0lSf3jpJdpfTW24wBD6Y
969M/Ns2G+QU7F2129QFyz7Xd3G3HJ1NEN9YWnL3G19v+Jokvfad8Rq04djq
W9fW8Aq0OjBDD6MVOQeMzjOA0S4fseZ7eeqMRR/QFOuKLQxqOdqh/kctWUhk
ByhVNCb1fUG9Yu7a9bBHjdom5AODKavYQO4ap69whT+PgSfXTai0IifVTmya
V+mDwCTDJ76d2lvkyI+TM/wL4tIxfLtbb9cyxoWjiggRAgsB7e64Qdwmes3m
0wYGz1E3rS70Hyqnb1pPbZyoherV3Qv6VYJAYOmBLgTvgfddGcoloNkvK+io
Y9Zh+be4Cl1nGJDnPlGKxhCE948uabTXgBld99qf4aSlAUy3Vxs62pqo0LkA
ZGr9+ZPkiva4HnoICAJ9rHpbKdXW5DdhXvzkyuk6kit+6rFYge0n9Bca4Ux/
fyxaUVv+/oYut5V+VrA6dReeXmj72rAG89tVb5cJfBy3BPwR9Xm+JxGMRaTD
5lE+R6yHw9YQuWCM0o007SV7rsLg/ftHToyllJfIyHTe5YC4iizp3EUU7qzd
uhIkUHf8JrQFPqJWs7pFVhIknon3zB3hj5nJ8Z0wQ6KhPYhpB3Xag9Nin0Bs
DodDVoUFz6BkVHujN6f+4rQZHaHgZtiL4S31OMHJDpHqCD9Yp5ZF0n1D7Dy+
aPIpyZRLm7Z1F1yKjX4Di/JtTEEkEQSc7tOTStuFuuhMS7hYzvF56yqFbyq1
6lIifqadKlj5PWWwRegPAWqGWWy7h71jAIQws0efwPFuV0xoECSnSuqaepvl
9zJCRFg+OZVWqMCIIwU0jP4ouLrCPkPMSr0dpWjqzEW+blcIK8fkXGCMUAAy
j+Rp0uHCg/vMqTzwO9eoyPR1otuBYjIgYt+UbHT0I9mMiO+VmsKhe8Nw+eHu
YKMDEQL0AXHxZsOP2sIyAvbe+3pimBbFSXnKwIognUqQbXVNTV4zVxvRzIwy
0GsOWaRcbKHzXcISarR4yCqYVopG/n9+mA//zglpi2QkBzKfEAQhBHqgI9Hj
GKd9Ym6zbHnVSGa9Pn46Z0yKL6DYc53mBe4pxbm5nPKfVCazlIkEbWiCllTA
Kvh9gBjmyk7I8mC4bMmqZXi/7NQdl6fD7Vok33QP6WvJ/mB0vUwvG3ZsPiHA
bvwnzm2ec1KkED8tdocm32eCoSKbnDLKegTYjA7F4fp4lRvtwxoPM8t8D/o/
hTzVqq3azIRHCSfBLrI4pgWZuuTEZ54Gdiu3dWo3wi1Mwg1Bg6BwSfPd+eYa
94Mhu8RJBfyC5jYECeGxaKgTYR68CTS5c5MWxIbuXvDJlQ9GwdfH7Uv5wY1r
pYDTW5AgGCyxNnmwY7mimb8E6dL2hriHulSs81vY2bcGjRBxXaXAMRawyndM
d9zw5l3ghbZOC0rX/6fle3HdC2H1L6Unzd20AM68Six8HM+kbcU2XDOm/loK
iRUA8ACYB+0V0uUoaUW6GkgzpoV9U0rAWI2gKtZmQQXRHYDiWHXJq0anY/AD
QyPGt5z0H+FBQB4roTgQRAdj5mIFjaNeVZfF4bUPy6Q03z8ugXcRRRlUtNxJ
k5DGLVClgToCbYTq6EqDMtb3+VOcNJon7b51bUIx/hdceIWGRAuuFYzKEj7j
4LIKJDqoWfX5iu5em1jpjrtTrvw0ncPCQFIXOonTdpU17zrTo+juf49GFw3N
40nopkD/c2UxjwmldCki8zvxOx2gIJ3iMKNfP0extcLLKzOI3hHIIvA2U5IP
KHMDYuXKA479sEkAnrzOjYGuP5jePAJWEXHwr6sqeGgJupcfOX9qdRbloKOM
gSOWplTndcDxrscVGLqhyHWMAC0rnuQ401022yAow4z7D93mBqPW72s5Tpp9
jCJcsfqHQ7ZEb4SyR7qbjSYkkFWwwvh7LtiGnIL9VYmrszvx+cDxiCA3h1QV
1JA3pgJxH77xZ+qC1SwuU62nkHTET5zECroVLuRv7aToWFuLHee8ah+PjL1Y
RUjBLyhYbxuZKU2M0BImvn/0N4HAagiHXPZOmwp/RWelCsG6klfwFiUhloLq
t3bVcxpPKYXZKefuLmKyODS3mqALCngchdUI9LStAuySoZTWOybRhUkUeni3
LSXUzcnyCuf2zl+On2hKClpADVgZXPeZcViLQWk1ZxDYbJMI3sPXBZpOMJBM
m+3r1sMy4so4H4PpWvMEpnXeWZGuvo9osiPHw9qGw50rY3jlEIzi+sxsr5ZM
5NapY2YSSMiNP0jaJcF/JWYlYuZOSdexrHpKVwT0CxRY8J7u7rQqm51dEU8T
v8sfT6m54C0eZMjL7F+HZUyYmsnFAAig59jQnOghQjsPjRoM96TFdM2loHsc
V+bPoprcZzWiuiLXotVl/qQUY+FF8StzwKTfS/T+OrSwXFA44Vn5ZJdu38ZC
IArux0xTH4kCbyHBUYo9bLXu4n0aXXOKw0qxKxGq3cKaMMEjsaa2D64FMUGD
2iw/vYXRxh0kO+eId8ggJYh/KLV03rE6YSg7fkIIRmYAkOyWujrJ9vEmZ93S
AnMK2JT1uK9IztfQKiDXIM3jWUUN5k/UsC3Wy/+BUKw1+TnnmqiIgRB4CXfV
hiwxZvPL1TbgNwzEHJZ17zhojC0vQCCvVOeOGGKKL4SrTJWQs0c9+9lrvFJU
smRxmke8hPRuShC9h+xY2B+OBQJS/0UYt1XeabJX10OaeK6QoR+ogfPlsaeL
j4XeVYny/HSb19ku/n1VXexiQkpw/+QvNJ0yRvvfU2XaLDmBNKw8o4w+0x/k
O8kEHAhN6MuFJEggTYsI4fGyKtJiWk+GWVC/4N3VcUF1VSMbPdOatRzOV919
dwkIlDuOzQqBPhZEfju7zANnDe6i9U3DQxDE6a7YOgF7dPKFTpnaq50LrDnw
FDTz2o3CNdW15xvhCB4g4r0AF+z6Q4Yaf3RRj0AOxIZfIcWTT5WG3o8ETfDj
9sFcDGpHWomR96l+hIQzwcs2+UsIgG0njqRPGy8wy97WK8jKKeHV+E24zt2d
KZDZ47ZNkCoaqCp+dGd8HOHFmYAhoed0k0Y+45T44mZi1C2Aq7T91T3wrOlp
HWvGl1ZkM4+RgzzTIVL9kZ9Y62PRoUvCCtnRJQzTkooDIh+tQEPjF8NXKtTM
g/Nh3aS27hJAs8QsQZ/q7r3G4Kr2cDkxlnOFW6W1P9SBFGt6T28N2tnCxSiR
qkVSJWSJ9G+5/0yfMplLFvx77gwit1YkZm0f3hfIT6tl75NzhZKqH1uiZ+p7
Ql18yJOeKY/s2eodPqmiusdnRcbiPrewY4KXvoO2IRuc5J0EfmvrlHD6/Udi
BvCzjwXPMiKO8WTyEwP9ef+xBXfmjV6Y60VMCEXBSHxgGbbjMrRIS5muICMS
gW7XiOLyC7kXVV1lpIMx0ZFVkN6Aw8preVU1FZPpLfMzllEd3CZzUqmD6sqi
ucxqdcXo3q/zzoua8wcc+JvgHnY/kfmQTuSi7UN5aV79hdgaYTDA1xOGAkjw
CeDBm2SMLBN3KR+lgjDhf7gBjGMQ8Xpaxv2w67EbumEI0K9LyamOnRCMm4xj
OePoShfrupnd0ElSP47z7vsnEbKheaFIXMHWem5T9KrQmCNa8vQiIeHviD2f
1vleQFBFqtvfw7/Lag0Hb1UE4vyXtJl7fZ+DQEqszRBEHSIl30RcAnaj0HJG
wBNTYMc2qD/xhzK7COaGODgO97j4NazLbzs/wWV/hqgf4nDCH/8Z1YEqbYfE
vsdk+Dl+nvaSZ8rHEPB5USyWD5z5xHdxASoYhmBdPEEdGoanF2ixgqwvCUsJ
bodQzESrNYF1z9aQiWOLlAgVR5CvvPsvcOU4JBoyatuAEzppbT3amXihjYj6
Smf92QWOMOMADOEI/tPYrKhJS/YcdXYzBq6YU8V7uHbP3ZOxR/phugHqVqEF
2p2XFbYq5GNXQLWf/jQm4QaG04WzXj7KmusELdUiDrZUY+aGD/A0acDgACL6
9Qn2ITBvqdnkCjJHigHSnGv34H64CPZo9x0KA1JFQjrS/11M0Z4LeGDdcL/7
Gs4WT3DTia0j0BSAjFEH67nfQq0OeBPzp81cOjS2bK8SvLYrwqxWZ0PljQRs
1O1BANqt1kdLAljJ1zzk2vgazNr7yg8MAf7W8TBHnO7yvvG114RNBNQ3AHnp
QTQa7Wch7BFa1w7O7OveSoaLa77ags+S2EnJQk/090qSXsHCT8S/Dw6yjtuO
K/SrW6Jfy9WdQifiycCykTqKXQWdDuQIzyCGvhjClhrHXXr5p6mf6Ua3HkjT
xRe/ATJ4FPx0slV9/6eX2ebez6QQZ+7FIOuSCu7F+qi4AWjzE8WUO1rJBrao
dAClgGVVKL6EWAxXtrqbzwG3K681s/ugulxY2h5kFtWk70St9EyD7z3/YFew
2FPjhNeYOCKLmQRc5iunQpouGS1r+6fMcrxP8BZf9LLufimsh37yrALV+egC
hY0hUkT62YpeCy9TWNqtupLvgeofalcVwXbpHEsAg3vCQ6W+3c2ribQOZfBI
1c0ZR2mBUif4qDJPjhfOpluRN7fEOhWqzgnjZ+Y1u3pp/UmuOsmE449BEoRL
Z04jkYM1H8MBbjj6XvBP/ziDRVHmtORfbg9Cvnm90av0mcLJSb+PNEbSTYmo
5bHms/mXOINA3MbshkQHPdVhqzaZUo4HbYyStzRd+LtLywFcB5J8l389WCg7
Zb1w7D+uKSS4ib9WWtQFRsBKmn1m/yS8HZzklcTlxW4leiCAhzVyKwWI2z7G
T0V3WHv/nOzHFS10rJQOnNEzO1IsV0DWXg3mi0QipLP2Od2AdAQw2/L1fYX9
KG26BL2Pdm7PILk4blwLktFu3FO1VtSSWJTRvXNxk/UV4i+ZGVsqLCRMy4TT
Z+lLJlgUJuLemTdxvTUuWcrsGZYdsbnsDfiCfdg7tGPawj3vYuaXGJKdJmPD
UeXmxcyl9YlI8EM4CVNn1/T2oaha/TWTd8yrWVv9VGpBzz/6SKuU2F2EDKwB
GcDPsnFi9zQ9MWbzGSzBuC8GmDybJldD+R7H5gJJ5rSILs904jJZASvnSgu4
MzcyMl35q6sYUki6gQYaOAb9mSMKYHQhD9TSYqgbT+DrDp6CY+w6J0pp94gm
MVtSjfHIUueTTAPux/V0ofY1S83cq+hvSCtW2uDy8EQIOHvPXiyaHGPxPnpU
TkcnvhUTLxmxuez1+hmvjpUK6YLqg/l2fRG9o/Sto2ADoWKt4H6dSNeIFp+Y
VVgk7Yy2v+wXiNuuF4k6fjoKHjk+hYulhsk4j8uVlAG8LC6r6Hlrq5Q/N6ny
86UtlkrLiXHdSn13nWgs51PqNGEXJQMiFU3TeOQ02WD6N479lIkWbGP8nJ6s
gYuqIIy27B+IchVFi5wZgOtpFnG84UPloFbLkyyXL36nspZzj/HYn+BBrdCE
pKPeCy5JH+P2aKxlP0WR/k5OsbSNGWEU0FXdJJQjSZXrodSYBMlK3+w+MbJ/
X46Ulls9GmnA/yVCCDPLS5dcTsAqh7mER5+fxoJt41L8AnQX1fiDIkeWI4TF
+V2Sm7R0/v9OZ6y64FJ7JyO7sm28KRtTmazk2BNM/e7Z+RdOVOmg8vwLwTKU
/cUW1lTHxYWH4YVVFmX0jhrTJyh5R7CU7cgrQmYBU4t5xJytZBNkIDnT9xOa
0JEjlyxJm60ShhjF+Nk5Gs923vsT1PCV33Ux/aJ0FzITqN2Xm1DZrQpdfR/E
Fdiqnw66y3ddYreuuBDM3DwGq/OH6N+oEA46XjuC4k7DY25f9nb8mfHMQdMo
sQLathwV+8qjQXWzVLVTF622wp0V8RJtGS0REoRZ1L0hQskUqSj1CjcwpZWK
cpQWZF/jrw/nmYEfhu1NFWhpE2HKBKjMoxZQsNBbeg9ocZH386yutApSAi3a
4rlLK9vN282hNel0hwmofTIuBB1jXRAAs0RS7oDNRfHDy53PLktIXhOEPMoc
cNBmQ/3C0j39JKGyhkLQy0qVf9DZrLYAr6r+wxda0gd3Xq0vuXwXHm5uhiSB
bnV/r0OvKWhSEo8L8Xg76AeRtXpZkG9UZAMBG4TnzDuy/DCaqAbH6cKe4C2n
e1UJdOfQOcTqVwbf3j1q47dVcoALxOi7d9eb20/QihzZGXTOrFnZBe88bt4e
bmIcP/10jxwSScCXxL8uWk+/3/OS3+2XAZvYZ98yj8wD6Hhb8EBHdApCJ/LM
FVpezcYoM9BS2DXxcgUOKg+sVOjM2PvTJbpO3qD/fEyoXrqDosmSpqwNQFN4
s+NDkKtlDq673MfXbSwdpNQa2QLBgrLTC7SH4K/S58f72IWXXVnaMXR0lInC
pEnVaYblAF+N1uSnninPTqxib4lTwuwgxwdsJoHy5OCRX4sAZjaRFJBb9P/f
OdDRWjsDJpLCNyaQo5ApnVP22Wf22F19iDs7zsd9eEaakqSguexAHOOZB4g3
hBkNoFnP5Nl2H2g5Cj5Oqppv5u4vVGDHoTtFlR1KvNdXhLiMMW5YtmK3hkts
+Z81LmgJmzvsYPRxlnEue+sodhrXgNq2COJ96RAKzEs2+lEzcOIwud0W4mxt
QVJf23wxRJbN/G8w4mN13O3EydllvWNUZVEqZoHZuVc0jzjE2aukSdGIXie+
dOKN6DwKni0BMzEfouf7z0h1cUBa+5NekPHeMvOgLP8ebeHPPEOR7+4LLktr
oKDrZv0KYDu0ZSoyStYMzT4wCO28UUzt50wDWqSEkP4/9EvGNm8AKNtINmOP
cf7tt5S0olqoIDmBq9W8dEZLoHHQCdjoa8EGp3pvdPYfuilvxzV+Pit/hMuc
1hjtsFP7jgWbn0kTBNeS2iTmml0XqeBgTWnCAnumtzrgdGifRHbAr2d/EZk3
EdZWDHTudCerN3nma+x2t8i3TP+k9e5hH2lx6q19kQwZBXrADP1LfRko46m2
QC602uqXc9V3Wx6V13fR2On+BUY6g4POdfcVEjqI8WNdMSUFNH7km9XNOgfE
kWWj1wRyfg9zWCIwe5oaccDYgpPTslP/DSJV/bmv5JfEsTS/HmVGIrP+2e6S
CWK9eGTvddwfeRHG55bOM4Llan6ItSTs5C12Ce+0avMtO643V+vGVynMRny7
nBNkJ8N/5AbFO8vw4cZsPZyOvoMjRV1HzrHRGUTSy8fyL3rd4C5sns3eVGTP
LWLDKjQ8DDFzJPUa0qzlRzeR6SW0dE07dMRtwa4+eoV12O5PhWNIaT5/uLeP
dGbv4QTRcTHaGONJCZQQvYnbuOrt/BokBKcfZyMJznNBKcRk5j8RNMwazZ9W
sY0rZVEwph6Gpck05OLCpiUAvJA+ZjTkWCvsdEZtVzwlkR81YEarhUmdqWaS
QVWNdx0cx/8tD8HBG/4kOreQ8D5RPS7BB+eub8bh59GqE9w/vMHAACjGH7A1
6DoATboABSlBf7CYlA/SH9hIH4Fj+Mpm4/i4QHxrunQMEVhO/2SUe3z/OvxF
6kt1bCVJ4q5BAkULIQT5ENVkNSV6Jw1deyNSBYaanSqC0A/gre6E+86DDEKi
Q60xsREXbVa6sgJE5mO848L0fNPtc2ED0pAse/ZSsmYgWVyB6n/HiR5ILBR5
JPFh8s5HG2TUAIHl1llOQAbRkSKVBMlJWIepTrFbd8XHx7E5SSWOnaaA4Jbp
f9jcBGPX/LOYo2zUcA2J2uhMAf113BjJowGOYQ2W33+7Ooh8XttWbf9sRaB6
VAIZ1Lg5WRy92ZaNIQ9zaV6PTAX8DUZzsX7+s6N3azyIawif/b7eGHQE8u29
omTGcThiUL6rjVjjit1YC/AOsl5/dIclgkUTZOBihhHZP+Ba/r8yf3hDAcUr
mNZALz96sgKfFIj43XiZGTI1N9MW9cgThIzZ3sP6VuAwCMoymHr+eHJx2uak
LlceaJQy5o7MxglnLPEGWrgsPV+qLOdm1IodlU2uJGPHyE18e80ikCYXSigm
nGfNPo8trXCieayI9lhDLmN6vEDLCJbS2YBJAyTOGQx6DLDk/zVqnBFjgVhd
vfzknNRiCiQhi64+HqoODLP5VYD7ybPigh1PTm11LaGIwlW20VUm2ElWQJjT
SIGlcyIyHeRELYD8Z5RDn4/JcX/qlym02uCaeowcDPKOTOApCUq6IEJdbORE
FnBIexEz787GMzLrQvrgSCfQkvtkvNhtcb/9LoZqzyb62DuvZ8ZZEDcC3vtt
Je64Sx+JpWGknpxXpu3eY86qT5TtfALfW72faEt4p5gsTW6it0sAy+FKxlzw
ilGDA+4NwjdCOG8NV7er9vh/svEUm3stRkTgLQlm98gkBI/t3EBgvaBv5PFa
RwDaaJveoN+/IA1yNXdM5MlS5Vo9esCzQcvy3uYzLiCLfuKdByJb4Dh/vuUL
LpeC9GYELb4nv0CxV1JyAU5s1ldhscWlr4pT1i8HB7k7YW6GYtxope1ad2lM
lDC7/MQETJ31hAL0grRldzwaiH3EX/lfVPvvPbheut3LNSFmipp2Ck9Nz6mp
n6YlMNIxgn6+6iprU5tqiHESdbK3KpgeP2th9BmvjY3hlSwlhTWdk8paF1ZH
78KXTepTKPtzU8aKTb4VGCvAmZR8R435Grid2o5qEYwYz4AMenB6o2gR5g1Q
WvzDl7xQQ/Si/Oc6mhla4Fl1sPxwoXVjZn7Chzv/J35COZ+EomaB2oqtMYsn
BBiyxaAKMiWr6w9dNCKGz6QMG+bgceqRyRFZNNPJZVg4UQBaWM0c5zbNc7vs
HjBwfLApg+2Vr5Hl/MdqGyIBKCsOJbyLmTngp3e4GvIn4Vik8yMIj8/tGnF3
yLsxbJyj3ViVVR3wwxltAdr9tmrguycILiElmtRGEyf59dsV8cR8+wFmqUOf
WyoRfTfgsrc1wthmxo8R0rsR+SeyDznNeKz/0WVw7qwzfi+8pA3Vc9obX4Yy
uWT/pXPqnO2kNn9IUOH/95LG1NPJ81kijTj+vJ3zgMS8iRQcSlXDTwahNheg
0jujLO9fbpUd7VOAe4apy5NBAtpVhDgej5Dyar0ZKCRTAgDhkfZ/smN6kzZP
a/c5hpLYOtcailD+2s8Z+a8LfVOQnbdBUC6Hcv5iB+qL+PxrZw9tSeFxjPqZ
iO6UEe2w0cIA7P93aCmF1xioFFmLv8xAoC6JlLUIZP9yrxlCzUbTeb3Q/8Vj
So8p8hkt9f679afC+QLv2lcW1A9BXKQjIhP3DDu/4/fKDz+2oF+4OY4xn57E
OzJFlV0tE+MSPKU9hVP+zSc3YXpXaoh2d1nRvTaCB87dKVOVXdETBvR71C18
0rxR5OBAoNR2U/SzbROdL8lTdlLwVVn5c5ChaNZylPuHU6+Q4jFTXAquROjI
BBqC9BHpiG0/y0HpzHMiWkKvsh3YbLLzB+E5yPW+2LNARhSuscO9hzH+bj2X
M9wX4Y+EcxbBrph4wf+iMiYsl8sT4o3dg0i0DStsPYyyoqKKCheGsO4tLxUa
ifiMn+WMEpV+IXpidrklu/Z90Czxr9UCffm07mIWMwA9UYKoV/xOIX2Smo7H
Xdtlhe++QLaXvOwm4RojS0OLt92dwUyAsGo9CamXBgGXFCYqPD15hdI6cE2Z
wWXCt4RAdh+lBInT/60290frBrJoD0Lh3yv8rUk+njfZZAbsmT9najsPGJMm
Ltv7t9Y3KIrtJMr/8gW4mUEHqRdk4+H6OBxCidFSaYujp/p99ZE8cZ2u1Jk4
3Qr+MJF+wtvu+X0bd4Yf6XviIJ1TXKtOhTniNiHOLRwkITluqUerPX3MPv8+
QXKZgrnby6E305CfLi39sqSm7CUZM0QvCw3YsDginC7BjINOyQIAv8wcUZb2
PaREUs4//Q8ExFFF6uhFKYkAoXUbGKzHyCGzShGyZ5z+hjT5FPdrD+JdehoS
3RgHE7xYJw1eqbezs7JyaxADHhjLz0G8j75UHMu6TpKPv24pkhn/aAtsaV23
I4W/IW+b+6DeNQR9CHa9hk12st8lJ7qATuZefrJCNpiySilOO0qZzd6TNYM2
47yuSKxd7lvysjgZovdzAO+5qCy69LQBA3Xvun9N9fexRCZGx3VNJTyfjqnp
HV/VtePtiW0BlScvJRi3e4YiFqhxiFkrVe2srMh7h4rhT/L+DTpPD/8j6C2O
B8+Pu7Hh6F25/t6mO5HNx/XiDnPHifOBr3tsGChb7VUUyjc0iS1Cp6QeejWo
2EY8DwFKNyf4PdaME/0wWOpDxDUrneDsjFI8XjNFapdkniGjYx0fOOX0cMmT
52JWBTTdO4VTkXutNuDXBzYWjKSd6XrzXKPGWoqs34CWcMJiatQ7SelTefQv
MdD/DU3ByqoEH1wg9h0jsf3fZdK7DBddXWl5Dv2Pp+bTvEHWxWu+4uSxLfDY
QK1xY4SzdD37eRX3hQ+wwnUMIq5fCZ7ZNV6EOGyx7Zz+TnsvXQqKIzjmSyqp
gL2TRUesgxpz0zAHpPkdgKY7rc3nldpPx0N4YdjABHlaOPY3P/n4cuKZyd2d
Mevsu+f9nlvnvMg4NKhqz1R+kzI3OHECApvhoTNxuSP4qsvj4sWE0v3X7BaI
1o77FjnTLh/PBOgKuuJFZViawKz6wYMQRA3TQqM0ElsurnswpMfUDYXDiawU
qdl9pEnnyl5k3a1dvC2qlLsRyF98bh3Y3fQQk6IDbq7R92jYTEv5dCuDST3a
uRCObL/CMtVHNMixFbFNnmnVmP2Y9GSY4UfLXRRRfsDwtv9b5JNw5kTXSzCZ
iygBcLrq7p4I3yzUxhFfTFLNcKVag9GCv0OkRW0VDRMFWbZpFTs3rkOIKw2m
Sq63pv4XmzZLsx3u9hLgEVnbb+TKXr607iIi9T/bPl4hqRrKly2xWp2Whkqf
fUHS2q7mJHxTtbJZbOczG9L/7HRDR4qhnKCyU7d4Nf6D3pEjyUI0cPdByj7R
8/5g39FNKUOQkbPYcD7fLqs9KoWFTnoslP/bG0Alwh15caPij/UCHcZNLPlt
S7Opwp38EG7O3kWpJmif+C/PrR38FHmb7LWprZvzM0WjEPeHC0m5kOeTxclE
SAZih6UlT8DhQ7jMHZkw3WtLUAxK3zANu0ypbkVG0FuOxGep3M2E2K8bq0Mf
cY6k0CGvWo+Y/5TdyQ+eFKdm4TfTUnptmu2gToZWrn9oDaXU26C6Aft94mBA
najRbizY2BUN87SRG3nD/5EZFeAQjwoko9rVzyiYz8j3GJob36oJujWMeCKx
XJ4NG5BYKDrVOJ89cbIyH9p4Ah6qb6p4iJGjN8zE4VwSTxTYjaFs1kONTVIq
i1OogXPUFIUBQWo4QBdUCtQIsjUwbyNfp1DNqdMMj+guVrKm+AjDpv1Z65co
Wz7VuvgMWp3lV6zigAIJMiSNkfFq6U2PHH8LyBVvQ9OZqaiZZeHBzB8er8f2
K+6qa1VA2qQXnKk2Q9+e2WQb+eR+Kmq4uHykkwFYL8BNce80T+PSh/ucKLOS
B/59NkXvyJIrRftmTv4/9I1H/TVLiTBa+pYhOBzJbLDvWt6DtjS4riRlfckJ
ZhbhBX85mYVLugqiv9B59hDviZYN9qMEwRkwhhv2rGIAdZbKBqDVeMVYAVOA
TsGgafC02ikn8cgELMR3UeY+YykWPKc3K50fgU2asUaUXj+LHn34gaEp6zqL
i9R6vEdQFWZdD8ofcZoiynhmcsPNGkrem/S1RyqLfsg2yqhmhCx3+PEfJMgj
4vmzUCG9RwXiqB6XRWTXIJstInxeKfgBP3mrzGKqRfxYSTxapv4t3Hg/B9dZ
Lkn4C1oqrCoBajP2nfT90SeANZqytUnnrhf4+K3L3fb9BUZE2WpVovchPWxR
4cFiCXtT2ChRcRqtXDue1sShrWyFfbaT12ptiVBNDn8zqSLfAFMb0y8XTjV0
UG8ivFnpDs/n0Kp31MqHZ3waCml/4X7roHZfsxgWWHuA7N25rNopIOe5Om1I
siWmJEm3XWcvcrn6WlXGtM3dz1K29m7LZdXTVJi0FXrF9TKh5QbZFnXL8Ayg
neFK1E4wk5zMZSJDUlpHHcDpKoVffIvRBmX37m42XVhqcY9QcQio4IrYlTWM
AA/INNlZbPNB0Lk7F8iCX9aYEVlQpJlthsc6JpZld05WAUM9p3HLm/UQ64Ps
zl1z+SbzbZjqPEP7l5xp/BPJ2xT51kq3v6bDmPnyhA+wZHj1IOkT2q09P6Kf
VBHvh61D5YpKcSw+Zj+KzdwKSZ3+XYW2fi8rAgpYZyjggHaLT72qHEYUU5Zo
+K0WxmUb0qarsfKcK382473vNDuq9+8tLOjBE8oAvqhkvg4KxnAzngN1xZaR
1QM8oumJ8Tso6rlYsw4nt1Zu7fB8b76vvp+AC+b1rkePyM4gITsvP2XYbtJo
xTxhezdDOfyYgUR3Wy0jfctYq5m8ykNq+L29FmzH+DNbzb8kmJn/wwLcFcB8
CdBmNUV47ZPJ0nvDQiapA4/Gu9ljJu8DqtrJ6wCqZ+eJI1uCPvYWGPbppoY9
XuZfY5gsGO9UYSdhp8fUAiKQQsrTT7Ct8gbYSvyt3D5QX/EUyuhKvpCLIRuh
Ik29zgK5PmSTq1izP6TB5BHN1qzQd+7WOFJ9/TdYTAWcq/0pozS3Vq91Cqni
W0Ud1eJxBoUgjPRvjpx3r2UMTq8Es5d9gwr2XPj+aCM6ZGHQ8e22YEUpLOVw
H1GsTYy6ZzMUfqP+i+c2R9suXdTVj/3QuJMxF5NUko0nlo+hFNRIuvSpJrDU
fLtqXkLWrRmTQh1fsazIwAq0ioAt4x4Xk/nMgOZ/ulWaM21qGyoYGvqvRsS4
4H5OyVaP//IPCDLjZWFnhW3ujD8qjY2CmmbRewTlJ4rgKhS6k479/xDx6cwW
ETj/Qk2ymxs2BX38JkyI2tzqmne/QgOQfiWHDBIVAKEGc0vSNDuisl6eHwS2
hFBcj6sItBS1ubasRqlCKeLvt3ygwSiwYHxyc17Van38yC69bT0NGDwbHIFZ
Ir8HN36fHZ65+vRzY4gtjmHIg1RI0OrZH7t/FMOnFhYVxmG082jS+u+lam1a
cqUMkfbmjA82NpXQ9lmC3CbajGIahg7LtvpZbeMx63k0KvQGam0Tm9sMOh+5
/RpzqH7vuFLTee+CEy4OkRAa99j8MU5gotzKXVfUwXBUoHfII0Ayd10Pqh0e
MaQRqiK9kZioZxSRH0ha/ilMWpoOgaHxo2hu5RtSoFEyZLeZA+v41l+BOQZA
AFpQZ2sQkI55TXAQgPip9I2Ir0XLcMRiDwQ2mSfgARgeIjHr2gqSuUEDPsOJ
BjXG+RwEkAb3Fo+rDSXMlG0V3XfVaa03pm9TZFLr0WVivNcD6+l6ysw9dWQt
z0XPYVvZ1QsYX3cbIdCehldfzl6UrRDuYCuLZm2l0j8SxEG9hy0URknQkmFu
7K/Ra2hzLfdn1ccEbLI5H0B+CAu6cMYL3KwW6tqryVNMxR9viNYkF+82KE3G
6UmUBwxWTIyzrq7o/2rcal9YQsX4sG1qbLNarJMMM6hgA0w4wvu2OXP0A8T0
vhxN/AMNrSka6iEp2sW3KG47x8vFhOULh8FmUyNEJFpzbjgZgRVli/SKCW2W
t4mr+8yWXWGVNcs6VqL8hIYJera0CBRKFxh/jrL3DswqZJ10KqConnt/TDUu
vTkxqVSKUCcMkhXJpQr3JzkkvVN/dVP2vAFZwu2KI0pUcHqXV1IKbAGxQWdu
/u9IY8lE9oj3RoFI50nUbeSwUnxgKAAUWtwa4D4OrwgYitgT+2i8F+53gJPq
AEKck9vYBdAoxR8Gx7AIVc2dpeJ+Tj+i7TqWJwxzx4KnkAZhfC8PqtVPG7Ay
XuFuCWiIu7QCzhGt+4pZrp7mad/46mbYqnY9z9cL7TBOOarrww3DOohP5Rt1
iasJ/YC7eza2FbfNDLWRuT19/Auj1Zu6eXIVda6s3g5ZkWWs7geCG/mafTKl
6V3QI8+6MoURluCGQj/DHkB2aCGvZ/a1UJkJMh2E8Og54edb88GIpCpvwky9
wviFy79lyM8a+IA8Cdq/zjxDT6qy5etRl616BuCFGD9IVnE5CFLqFDC7KMqC
mhJvoofvv8M/fgYiyWJ8SiBXPATx7GdS8sqV22hAaYW/OpUsfvMIxfvp3bBS
7M9TFwTH5zJyjauh/Lz2HLNr59aP6bjBZ2mr9pQJFlEpQQgia04Zfu2ciW2G
8v1WoQ6ZiuOgOXLNJQAwJ6Y3apKUtrbhgXO0BrNMoWVR0db7M4wdNUZ+Ndt9
iYT1A5p3lr2t4l7m3Vx0FeuyWQ/Wr4QcwC2lBUaU/lL29dUV0iqfHmql+Z6E
VSqp/WGosxIFp1KQm2X5Ez0B5th04PtjqZaI2gO99/7lRQBB+cAQ5DwpIvS0
equ3iNFqbe5nK0EPbWufG5KnSOOjwyjIpUpihG1Sgc25fDmNhHspxb25zBG5
VYdGQY9sMLbGXkNkiqRl6j+XyM4jGswHK3hPphvTAoWduVxkxKoAzA7rEEmw
WoYeC+QoaooR0++EzasjmFTUVdKWS12ukoBP2CtejyDck1Qu/e3H/HbFbFEI
bJTT0yRHAhB8TPQOzVUq5zFaoKi2ZL35QyzPEyM2nWcE9WQwtefefcIxQROu
pMBsHYAdND38uVzdCC62mRiPZVIlLA7tKz2DuaG7oZte1ZBE1fOcYpaABOLO
Y1w5uqhS9vyd5MK129w6jCSYRhc7aOL6f3Q65lF/db45Ki4KbNfLnA3G5tFK
QaCTQCRizIh6BQg/MLmd9FKFk8hQuzP5aGDrBHczx/1wJY6+AeH12ux8eo/f
CqkraIQdeBOaUcPtPjfXfqnlIGIDpYymPuN+S6eKfKuyR+DuwwU2VSJuM0jz
pGSXLt11tv665ckZarNW9N6hqHRTIQqUb6aInRm29Yj3uue7TtT+Qcchgvym
OVICSYCMTSIq/YcwUqdHZx+JerYmV0GwrnWmj74mT55vG0YKoqqD5Sovo7fZ
SDCtafZ3BxOSKzNsfUpjSoEsCo+cXQI9QKzyLXyH33WquAla08Jnxyq+8hom
ft2E/x75TJ0Z8sIu0QK9HCvbx80CAz2cpf0nHZBw4rEeQfb7fU6/zHGKKXxP
YMXwpYLRN8d0zGSiLoNUXvi+xJ50XTyW4z4LjmBOX/0BnFjw+yk+Wf4u9ING
TBtF8Z9VZ76BLxiryR9aSR0rzz0pfCs+RDyEDCyEVTcjh/B/vUWz2zT2EsDW
92nlCt2gwKyiUsZrvmg5MyEHqdIlzD1c4KKCh0Mav0SitymGB9aj/ADeYeSX
RNaSGNR4Qc8F0/V39PuMMbZ3KDAJihp4sEL8Ohy2/HJuj5c4o4op+bEx/Cs+
bo7R2YOu2V92OK+rny7U/T5X6LNMunGJjC0CJoEGRqngJ+FL9+Vk02lxd63o
bVE3pfY8Txlu96z05y677e9jSALMqdFPza52CX95ya4wDUxpn/rUfWo6yg1Y
ec/erWta0HomQXICzH6xZwfO33qNc0st/5GAhaVB0Q8T2GevyMO74sanoQbE
YFZ9MobGpV7hsTbH7LtDumGHLxLdsZJO4oHEGxH3mCBJdXvyLxj6CwPXGFHB
in/jkGiNxAlku/3iQArZKT8rOwSnG+hoxEyCdn0UIDDf3Cv2YPX7xQ3G9oXv
IOFLYoQ81ugnOSpR472qPTHGTbmviJozL7NO5P1fD6xEUI+IJtXdtzQIoJDH
ws+ckeOpfTLpfbUgRMGfPO6tAYUosKm7qQ2mAzQhnkGKWO1gPR9q/eHV6tsq
FI84frTLoNRPx2ZSEqvAZghJMGdW4QpHJ1NHjTkLXkPul/Z4tT/wCzS4XxyM
EfROkFN1aopW9LOMeM7Pgix32lLhI8OGDkOkJcTA76bX3k5XIz99SAHD2tzM
5QptUTigzss5/sZ6Lf9+Knjkkkr0qzk/jUE8VIzdJq1oYWf4P2xlj0EX06uO
987mlpyffqsgS0sC5McXzgyU8WO3OPEjxW8rgPQux3Khx+6V/P0/v/wYzrYL
Ljnp0HhLaoGdGZZxYCbAGq6g+hPDkI7g7E4uFb/uEMwW7Q6H1Bir6CUJRc06
b0mGkhM0YgS+fURmVzMZtdeSarOGcqqLJjz2uWQzyjPYIZkE0HYYBxe6dUOv
fr4ok/+N6r/T1KDkPd2zlSvSewPOvMLhE7rTwMbDpckOw0Qb761Cy8JxHmxI
3iSVEEiZiGgGSPwQFt60VQi5JFFDLxo9ocNVvop1IqotQOjFseM1yHnovqYO
eqsMeZJoDwrM0t6K6aTjEn4IOEL1PFwLq5WG1l5KQTF/mIF6j19D21qANkre
s4fw4bRlzVpJy2dhtY3vZ8Q+u9fx8Z2QUB0xf92Os7WRjfZk6+8k1C7oK+Fy
cPs/bA6TLKhhpZ53OmxiLfLN2mKdNzkMaREt7b1ZcR/1HczM2t7OZQB2BixV
XhoNjGDbi8RnQbLvMZhGUFJHU243G14ls56K26MGSAvajUr2fsG4eLDgkWD6
OZcPyPkSN/3R8BJNfSWt9vasY05SjdoCsplC1a9rrXDjARvk0QtIUL5HGBXn
LXjSC7KXfA3fquwxzpijBjkZ8aE+eqx+uxn/Xf3VJQiqq5WXhZv2SBIKaXzt
XTfHDKhLnKc6ahgBffeg6VdPKJ7IrgDPD0MOsOMIBaiJsr/Vq49KKYTSwcqU
5R0MVYfHMjo1CVFW1jHVr1E2YXzlmOBsBqHk5W9Sak7aX9J7yVAp6TfZykzm
WDsJlWNm9C4whtcYv9spPu5CXn9eLLc3t1R7/U9QX+EM3K8hsB+xb8IAceUZ
DUcUlfbzGZGWgqDZX1R5kfUMsCZZvhsvpVsRsfksS6cM7PfmCbSFZQZluT7/
7WCnhm/zJBi04lgipcVjrfV8VAdNQlfrB0eW5hsCTEwq+AfMLVipp/WM5Egg
LskhCAf1BUp0S/gCOeKZdb06dko5kKsTnMCgnVd7KHC8FKFZeZ03Ly9/MHG4
8qIcBbOUPlAi1jku4Bown/EjrVCqpeGv3cM5mZnkUXh4DZ/sXTehx2sfThD0
UfLNiR9IjAGjXG99+vrLoUtHRGyQHiIU5V/zUzSXg/fqUmWEtuIemwwT4f0a
69biZxlgi/leRW8YsO5rgxN9lxd5j7URQBIg5TIcSgPHeuCBuy2y10rxzKtw
OheYe3wgZnycLVgfKi1YvLjx8BWQFujHz+SmaRzoPCK1RWp10y6qAXOfF5M0
8y5KNM4BFnkrYRF9gn8gnXaNgn5YGXd7/IeqVafoUJzdqtAzlWUCjcouTq0u
wocW6gZgqENJp+QJ/qXAFovdhByQkiOP8zK3wfM/mK4UYK36F4l2GC3mK3Ay
2TI+g+LsKu3tBVEqBfsqHKQraTR6yzJemDNUi8wFCvXiHvxUQgRVU274Nag3
Rv78zkTdL+WaUQXqkqyOcgSy5tUlpuiNzLX4dCsvRWxw/T2vfK//JHwYq0Md
J/KlZY4DnIZBJ4v82CfQsga/E23tCXm3y1wH7lFZIbHobbCOBDMG8GbmqZhr
7DuXmPCkbauWgMn+C6idndTHD2DZqHdE/bdpYmv2ANCSp3OdULEHatwnWqPs
vErkcuRjE6mea4oMk3jTm35YTebPWl0V4Lxpa+tPfmNrPHZuaBVuokd2NCUY
czsNgWBS5hVn+613qdC/+w+M005ByswDXwi0jRg2QQqRP7P6AOoN8200up03
mndH4/+Lvca+fIXheDF7VH2PaBtURV3h2p8hcihFI5GRvlS0Dznlcu9uSmEx
Qf2lViobHbUScBuyg6jkrebYXXL1NKoUI86xpxMHV5I6Z/RosDnw1i0vGK7k
8igVXRd/QzH+mcVEb26PXmRU9pEvWNzKa/YnkDHaPrXxH1QpZP0PW0aAkwfu
x7OuZ6FfJR5DtHjfdOoIWCV1olicLXxgMtA5QZnN/8z9qyVGZrwF4/fQ/UCS
bpzJXLsRi5EkJsv2orJ3Z6hbY2i8fauIjUG0sFOFl6J0kIlS6OBNcJqRH6YO
mP4QS9WTF5qVCPX0pWcc4GS7qjw/K1kIua0i5kr4wYhugn+E5MFtw+xMXEgZ
5YhYYEwYYbqUUVXqIoXXis+3nnwON8HWtsNzYiUVgUmGUsgcVmdMXldNg1RO
+nVsobXrk0hRbxoizlC+f/LNRwjBBMO1r/97qabTLFGlrG8bw+oC9pXjTXrp
Jzshj97Eo3ZXk9ZI62OhP2MzpT0zq9A491Z/XSe/+L8XGvG3nZx3jYKyWTM3
6qonURXL4+hZXwvlbxRzMHh3OP4XJKVVOv0tXbzCFVhQEgRYZWmGQP8+xiU4
SmRNxbcJn3Jvyu3q2kSxkUWrTEQLcugKxKb2OGHRWl1ipDlE+sLKLVOZ4Amj
w7TxpQStsLvHGzRQ2uAR8yVkzSlqbNzyqgC35UNc9whMv4IXEoW+7ZJXscXm
cwbfjMBFFehGwi51b7BM4OzeaYxqRyCnozTHpzj5UocgSnRqyVrcOCDZixlj
/It1AwDv7Y4IOb8ztxuKpLMpBFqeyhuDHLTwqC4I5zVi+sSvl7SdVg2gq/Ge
3uJBeY6o6xvtjR29uzQE9pTsv2Zu+g/DApH/tR6ogf1VprBbb1/mqnqgnXxZ
+WRcTY3C3a7phN3R5KOvy7UfT/vDa+79Au8aJkjA/3McEUU6RPcbiI4snVwN
IN7jfHGZjjUFIoeNtYsn4T6Wuc5LZNvsDISGyeS4JCtHN9oOXYQIsOrSTBHK
EqXIQVQ64tMIjcbDGH1d6Nes1LwqayBcu4KmmQe4Rq5C93cbER6Y4gko0HMv
weRFtPJcWfTaTaqVbOi4NRgr82NC1l3k6F/ATDJHd+PpOdKPrcHQCCsL58jO
YuknbfgGRck4OQwM0YvCwHxTigr7qdJpSssB85bbmSij4ayWvaXkBCdzDJvV
9COal6x8NIYsnqkt1ekLqVhO2kRsseaB/3p4thVAy0QMKNAlL+oHG4Tpsonc
kbMa9W5UKHlkRgLf0Sy3ApOpfhG7Z7TZ898SaUfsFLDpUKK/KLip9JTygMZw
8B8pBlUPkiA2mf3uw8yxsUdNCKKlhZD+9OUu8eE2Z+GHiQILckhjDF8+8sIh
xxFv8stdOV9Hze+QTl/1X11lKzvqtxb78mjRzI88VnsqEVQYnaON4Gc7r7UJ
WaK+wghV3x8Na4YF9VWdEyF7DsF45ibhBgg9eBkYexHPqHsym3hI5IA+KoNy
mEYK/N486Y5cjEvWPlX6svwpEE3Qo9RABvQyQed25vdVJUQ7FKNvse8e7xt0
umPVvRNMH/wR04glSPxazok2i2maOn+034BTBPZU29rzSr2TkJFiU+x9bD85
aj4poYIm4X/EXQHoN8wt42FFcnpEez0umrFLOpPjlUr1Eef+LaVtkA4X8B+G
CAT7gCMsayve+fdt4OdVxLOPgZqkpRBJGE6sFKcqY+4mUgrlj5G9NgN/f3kl
fvmnY5SAekZIEkxk4WiK6mLAh4nvddIFJRnqkgjPRD4gwkWV5dYkxW0IDKfs
xhZ4nvATMwdkh31EhOfE6D9eCcUbmXUueovuUjYQN+Fc4IFfplUthG+GNG+u
qqPyccTEfDcbO8rHkIhknk6lq3m4+qQZhdRD7rUgsALKAnnhxn+pONnA+lg0
hTNSC+nKYl7Nhriv61pq/xZZtofbXJmTwIzwBmLLTTIG3MT0WwznZnN3ei0k
pJ7TpqGWxFpKH4mvyElesmWaBS+H153mwcCm2daZwK/3VPsXT/4YmgOt3ElW
oviHot0F93Xint4S7hmqdHFMwotqnqhwor0RVVPTip/ZznLgMTkkUIbR316q
22s5kqtgRVvavrUONPjTXRFM20X0O+4aT567mYkA60Rst18sObLT+Ryb/PgC
lTUxAeHQxxSlT07upqcjlBTp7Palx8tUrG7sUXCnF3LNnBincLYRkZttmnnU
o+f+2GH7G/ETekBb2IiFxmi4USlcGl+IX3roZQ+Cymw52wMGdA2VzdsaldaM
iyM+0sz7PJiwhEyZr+uwzTKsa+MpkvQyQYM+ItRiaUtphIhhIR6cjfIcwb66
DtaULTe1OZZb4UIPv1DX2FZeRMMIdZ+Bd4Ey8EOnuw25MPniJq7n1OZtHuJc
hvZmZiqRJXckIMYRMMm24HJ8Mu2z02aDN4Pckxu/Ik2bk9nUM+7pyWyJr0Q4
Jq23VJzhsa0q/Or2VuOLFt3efifP5bsW55o3FuR+qdElwaSKPdqC+ufNDjzS
Ud1cAkJrWdUrrk6CNNLOgvzNkFhbD7dtJczZjeNH5uCwZcrlr025i2/bH8Nj
gY7CTFxEzZKjv5Piei/r8OZZINyKP9ocT/t2vGPBhxqDXMIPjKbcEci8e8C0
ne14jXFY0U+PyzRoDryAWw4zkaLZ3RONiRKRPz26Gft1nvezs2886xvs8CiY
yB5anSSR4RYOpJ1dcetucNFv9u6zrNRtlqLFpTnGoFvxk63HTpLMm3p2fCt9
8buYYeEhDSxLu0/mV+VUywmkWr7depFWakHG/ETiR2czH1//kinQ/M3QexFP
qwhlR02SK3GFI9lnpwMTJi4MPqVu1mwn9kM3WK7OcbuJ4KiN6rbbjTU21tUY
nyneak43kYVPCdnzl+7FTwThSIWr4qrxsmU7U1LG5uTpk8xv7XXuxZXXrNiV
iDYPb5g79XQNlDlRB7XUFow+aEsrZAKZVpu4IJo17JQVdS+rkbvUli3X/0fj
uIqhWO/usdemzumuRDQxlhTjd5LJkszOc9bI0jwaWYWHUgeik27QkBiIjEvg
azN3z0r5JeuzC+EcIrs/iGH5gpfqzvKYDcmsk1ZRyEH2Uaxmxh6BiXYEFOvw
EqqQ+Y46Ziv66Ve9XF6dhNudiFvm7XP3sUx6HLISzmmtan8cs0RZv/FpheQQ
+KiG3m/0zyTIl8U4eHSbeq92WRUWATrxoMLJJaqR0FFMoiKP1awNJ+fUUaGs
mVeTJSopQhwrH7WS0m3PskG/ds78N+BSwRcBHpyNTku+ln1JanaHy2oxZ5n1
xIBQaYxQ/ssIf/xmcXbJgZIh7FpVXo5hQ8MCFSrpLEqtigEKwenww6EvhLtX
toCPQ9w91D8mo0K9dlZwJKSmi5uDiZdrm3Uk7nSupTVqZUTln+A25lyHz45t
yyP/sUcSU1DCn7Uitg8X2gnwLQmqpR8uhx3u+oSO/kA94jYib7GYZm9Jwhxk
O/Utc2uGrIypmWGbEkwrVMYOQ7XIC8NAf3SlAMHJy2aeAJHI22OFDBVMFB5S
Cl36+8Y5louWwbxJKu5OBBSRE0bUBCGo02lua9P48i6yxfUvmab3MSRrRb/U
Y9FkrdPo9GeIIeoLGcICPfIELgvXsfxiKh3kukumm62zCHeTysCPZQ9MJso9
O0wdzlQTY5avLTIZOGLmZZsm4TyhUzkrPsizsP4MJ3fBat3pUpNNlKJx9y69
QvUiUXSBZrzCELk70PL033BmqsQwe1ZNjP5cf3QfOenjZIiwvSJ2eXjjmCoz
HcZinhoeOr8AGTV6c74rWu1OdjXXm+eKuHgd5rXhNimWd9pQLtxiFIoNcM/N
SqvbZp7vv+ifGjpSE19Hws3Ead8Umpy6vACB69I6DsZoV404AqyLWUZ6LpZD
j/FqbqZlyWV66fM5rIOwDItKX/578LfWXBP3gY07LU74aTspGOL22Y9dly1V
Nxbsu2IAXl8AvH0t83A/6nSVhGIpVwoVnlj/H7Edqzt6ELqyjWBpc8LS6LT5
+qMAXLhXNGOw/B/q6lP85hnKT/HmnOYZyINPp3eZVkSk7/PSufozFeBzxXfk
w6jJM9EQfsjN+zmfF/X9NDVBVHLKmqi0Ky2GCZkO/H2SIEVYr8MzPjaEortr
BgkUqkiUNxxQ9V9fn+UTQxdbhUApsIdHc+sNxJoBj0pE8qhYODq1tFIRB1oN
F99Eg45tmAvDVaAaObPqfBcXHk8nhktBVlqNhDMY2iWK+JqqDgcEcl4WLYgW
No0NiSQ7LmpLz1mFM1nUJ1mJOEenFwEHMfi1UpfxjuqlKuvzmJ18HaImTAXL
q/gOZepiT5Y369sRMowW0l68+b8v5loY5KkiWU3okTvOcAcDP8GVpQEFblOF
3hcS5Y7TgTJjvYYX/N3PdkXRod+qBdiLFISkO6gcnmm8wMQ2nWphD6DwGOoi
QaXtiHw2cjVleRhqY4YZTeF6KT9bo73TPVWgdspbV8Yob3+TqADx4BJoqdZA
2Im+At/LqGlUYxU0YktuZQcVUJXxKKkUyFkwXeHDIKqs3JWoNtaPcWagE6mq
MUCbyRd3t+NOWWUbz7F84/zNbtqTWLfg1VB9UvLB02d1cn/WSn5ajzoywxpz
0VDoqZNJbJvY4IHtjGtJzQqLM0XlTgOfL/QSXJcpksz8A0jnMpePqzfb9Oij
CauzqrDUY5KiYSUyM/hQc/aEyvKaWD49vFqaRLPnMGw4k+BaZOyAbfp0Xyj9
FAqRL+aIVaz51GkTUZ5bStORtxvVxHclj3NjAlWnLIfdR1W3OupWAyzNvBYF
ogA1F6gNoeQoudT9DKed9QA/ILqh8suK7BatiqrlMJwWZtS+QUk/lOS1e8Wu
UPr+FcJXqjrviz9lmSXnwIvlgM+CgOO1j+OA9GoscBpjFUBGaIsQDCbSEXs8
4/FfXZhsEY42YRmQk6bmXNhipypLvCdYvTEmp7/0VpyYAr7pO+Hil+7biVTz
t54ljA3mhn72LAWnLwEMmpYhOZ7tAnCD1D3QTC42P0ZpoT2Nl2b+m2tDKXHX
ALzYDFbJr3O3i8AEbs1fo6v0G2AzVF/MFCS+dDSB/3fg6LCwnV2hE2cfzBSU
Ux+vfRaK/zAdmvk+ctaJxAGD4IoxsB/o5mLIl2pWX0U6k6xMkHhC7vp/i4yq
3cmTbAgfAHdMHj+g3v0OW5fy5rImBq2Sgmc8Dxm/D+e9Nhb8lu+k93N87Kz6
4GHB8KRL+6ba0ldCp2IEwQTChGbRDUYYoL13cm6+bYvxQlC5sP29rTLCV7dk
ZEDvM65TIDdesSZo4sFEBGKcDe12JdogfsvRCYeEl7Xu2w9q8tON/emVJbBs
SOZsyMarHc21tZgxCpTgEtxZgugdhPt5OcVZOnEscS2uOstlJhsw2dcKEIFW
mca/7cXa63msm5AX2LtcfArP4o046RPOqfFNdDbnQlEpeab/jaloaLYtML0p
VggGHQTwk+yGc+NYbsVDiY6gnfJgsqDgQrKZdq8cg0a7WOiftXjYDcDxGO4C
TVlQKcvUnSiKo5VFY3RNodnMbeNKkAszZ8BtoZPJNITSidOskJZjKwkN4R90
34TpxaIemnXStNGey2JqfplxlVZsMxk5RrBXUOnUE5PAQQAeegs2hSlh8131
tQlfTBrCmShd2PEybsxey0LM0iajniVtmtyn/1tP1KI7Dan0MoHRNSjRqttC
5F+R86lfxkfgAd/ky8XUsVpk7t4StmAH/LRUwBS5pobq9dTplnNwJg+jW2NX
+SKT/AOWlOWflG7upFLgIiWoOVFX2XuH10EgOzxufx23DdDrQcvEGNJ+UXsc
6XudQa5cz75akuoftVyDTKBHNCP2So1nHX25bjbZJ44z6iivEw3yTj2RV6gN
t6tamupFpr8MgEiX0bFtv9l4uO0Zx0wODVEpPSyVSgHVaIoF2dP3/HeO+ERn
r9OEUmB9Q+inoGhI40Lre6ex+eXJa9pmnovKks7AYvyy43Mgwxk7LEbsJcHn
bBxzUABSVe/pMdMb2aIVJyb0oWjXezrCuGsrsNVxQ5ZbQlPGBC4KUkQ2cfja
jd7JArjfn02tfvW4U62W5fpi+RgDoQo7E1Q+G+pLQsAKIfi3dt4v7b/0aphI
ThE83VoTMzADatEbLyUmKtLckvrHs9PvCEjFlYpm9a/XXkdzjUqb7YnvgNWY
E9QqX6F6WJS2c9JTihXUwTWluWHRLKoglgYcnlE4dVCpyv5KKOg5zmJ0emU3
5kaYKso5MKKW/1HhtdQorRgyNB8NQc4p/LgmgRSmJ9mHb/UKZH8wKkC/ppqZ
KCEt4DPeTvZpxHK2e/WCkpXIPOWl3j+5fHfKSS0jjYK9F1fEljCvPJe6mdQq
95IJFgEo9InQ/HZH19fCmrhg3Tait3Hm6E9dlhY/4sLH3lX4TC9a4xYN/HDg
IkGM3DKnbLmt9EXn1lba08IgxNIsD+RLHyuivwuQbvdACrD3e4qG4qtWmFIW
5Z4MoPGCDCGwxR8YdYCWZK1uqocrnW1Tt+yyKQ2s+LXTWB5MyF2hp7CQCnpp
PRbVGLBQsAH9XgbHZUtTXfiCn7c183jvVZdrAYeV4W67NoRhPWEPTe6L/orr
ZW6otp0kLxWzIBNgDW2ddFIBMvPlglzUPo3Cw6sumG6ybyU8iIal0IFSthZl
goTB14ixLjHxi1ULNduWN0B8gTCTSkDf6694+CDeN4FCU5rRWFmt4Ta7Zkrt
EfLzyVIl5TFB0el1+xqQt9YCUm1eEtfFPaoS2HhP7x/94skNiN6cafFoOesW
3xe/TT4aCOCzI9KH0Tf5t2RMFUepgMF/ih6UxsrvPvVNVm5oKZJiB06xT88e
jBdi45J0SB7dTD1NifOf8PO6DkdYmVT1AHWaHBTeUE3WaBAiBSw5uJEmHS9f
anTbUrzqoITWepDusOq+Se35mzFxnQVjbg2SGtKjlUOPPKnsoKu1b/mYZ+mN
lfkKKio4f6kjH9eAV5fRm0JaFePOskG47wjQytALM1690B2FuVCSho+qhV50
5tvuhG3cbaPRLoNwhwYLfm88s3UO71ZNYaaqc+S5tDlSNBCgAOMlyf1Faril
HfpSklW/ZhCZXKy6vFmxSEdIiAIAM4b6BNORGjLlfUI/6r/qtmJRPoMqC80J
kvpOgmz4MXLZvW26VxKiXiQpsBmdpKYaCEvZZJJZnn5/Ii2QZ0h5W03m2FiV
U2MuxYlvy0QKHsQDb3tk2bpbR3YX/EF2HYF/X7zKuoImLqw1hrtQ4bhjcJnC
R69w/ZRVm2B7JGA+/m8avP1+n/VZR97MgGzIJhpZP2bWLB4aIrUU5JSgXwIE
GZ5hkfa83GXTeeQ7Mfyf8C3PP44yINH5vD0yxQ4kZtePpf4u8XA7GJbBWAir
5lIkqSKn8a0kGbpwvimIV25jFFCa0x6xQ2t6PxptVJWvDsp358QYplPgPJeS
Fho782axIbuhWb9efslnqodAKZHglscrZWUFlF4g5AsgLX+bQpZ+rLJAQdeG
GqUEtR24uS2fmSSTczVzX9DKZFFztWYn2vGf2k6RtD9hQx9OtXDPnH/06PER
1vgWGLvuXqInWlnhHGsy3oIM1p4osR5EcWnC187k5Se/ibMcAo0jwtsUGWcI
dh8ilXwf6/pywsvzv33ZuMrVeJBYSvYd3U+0nAl/OP59FZd2ywQ741d0KARj
0n4sQpn69lacfpjqaMxVU19yznVqQC4vmg+fYmDu9rHgxnOlPYPVe9aAsuMA
7UMK3uIHNeFURmQyDK7NJQhiNXAZZapCTrRMV8x/acaei2VOK+fz3ZCRW1L7
eQt0VQINW41cTyE8GfCUKNWU/ScGd2B7jO35t9pib2jBTfTctoiY0MVidQp3
FXe2kbxMjN0ICzAfY3odz5elGTa2tfGa6/JMNBNrkZVKH+QymqVpRs8Aetc3
uGu+9EFFGN7Fk/Nxg+Iv95QxYWO01s5SVm/uqbiYsJ49BSQwdkvW5lXCJF5Q
6wnoTPx7HOWdyZDEl5vgbcFeUTKfGJCO9/jVIOdSYondhGB9FTOF3Ag0Mvt4
6FT1k4FsfdWQvn9gJ181h/3fR8suOQyfpbWviEx0U6/Fmkmt/BF1vffSbyQx
Im4mDXj0C9SAIklTF0QTKkP+pPHcUM3hJ0u5EWOBKjMlQCE4kDgXrNolv1Jt
GUohyZZA/DQ8kwdlWDp2bJ+//WFfwz51m4DPHZYugQi4ZUwFZVgmD55ZE/KD
BsvQFgYLd/AmP0FGiyNCj6ULhIB38PsWS4QjPkfU8Nk+6yKhoZGJSzFR6GVN
oVbb/QaVDr7PuAQXDxv+2xtsySrGRHPgBSix5mT5HWGDJiMQHLwb/fcpbud1
CZUTsspV0/vpLGv0er49+RGny1Nh0dJgY1NSMLnCAsxlpPKtOskA2kjO7VJG
fyYxGun3zIoAVBgM+tUZZGDiJxASEpGlUz3zyd4hB09gX6TODQ4Lwb1Tc9C8
zS5EXIRBf8MfDTT6SxK14NgsVzOapc4S6kV5t/XOn27vUgAOT9N8zZvD2Ksv
kTsRA0bNDbE5G/M0glE8BYCu8UQ6H8yt14efrf5bOLfrZ/vWi63JFMVX+33f
4t1vHULeyU/PwsM00iECmupqJ4SF2ZRIqh6kmQ7hy/SeJiNMkB87k99phDfH
8+WhQ20ndwFIfR+RqIrqrDeL1VprdaqPRFI/2ihGsbubP/RaA6SNa8pz+8Ry
D8tkRvlXVIE4AHYh5zJdHrRKRQ/aJm6j/zrVta6dR/mjw3byBDJTQqzsrluR
3QIcIA0FvEjwZh5rF+EQLYXmd4bpLwCF6/kcslwltHpjxNIIBB9UXK9tADq3
sItXZv3M4TsEy67TwiPpd02SPdpB9TTB7HwGNJFF5dkmo7kSwAL9P9dYq2bT
4ZRZiKt6Aax6hl6H50dKxDXl577Jf6S2SQUC8PHvGYED0KlC8vp28gzUcMJO
WaRh+uInDwaJzd+idlGyddR/wQXKJYa66drs7yYOll4UjMFkVWFnpyr47GN5
bh8Ul7qrStDVGzdm2kX7RqbyZW60tLLEv+Ixc9rDAhohYW1qOx4oepkH7327
wDdKq6MSWVeb51B/l4oLF9assZeTAxabk0WWnaCRIkDRmp88UuUe1ZNcraln
NbevygsaEI+lkSrA2brTAj4+BWj7TBoB14KenCOeA+RGhmtnoh+Aclonjnza
wyQVcr51OHcQWfYV/FIUMh71C5/0VWlcgvgr1eORIKgI19QMfSQdjmCZ6UEx
UE9FF2Jontr1t6yJ07E9BlUy4fKOAzYmxCAjsI6MIx6WxqCizM9WDsiSJ9fl
jXi0osuwYYkf7fwBv6nGggfACe8LqRpzKWbDEWF85zpUfbBq7f3wIRcBC1A6
pJHiXJ2mcjrIbxODltMkHqJ1d/v09UQLl7PpTNADOpjIBcmAZun74orISIrC
+42efscDqZYPQqi3vYfrU0S/X2QlsCNXtBh09IXNhRgzxkAC1DP3hiZ5hIEB
K06L6PyBf6MDOtz0NVJ1zkw5XUsPqWfXIoCkWB7ul4jTuc3qBWO6eCGyTdIh
37g6hIR1gDAC7IvRqVN4jyxF/kiNNUPOn/j7L9kJJX6bp9PyHok8uzuJSn8O
Hy2yjKq94skbJCF/18oUTC3s8A1Kpbc4/jKeTUmeFGT+H2FcHK2UhT5uP9Kn
bzrq08ZKZ1rmx9BZV6+e/hsS5+4C70AG+jAdhIwq33mh3Fy/LMeBTqX3NSSj
fMCmIj+7ScigJ95HmgFEmTpvxO/7ccfFeAsZsLGOOA4HGDGjl+8C4G+NrEQs
1curyNEFYfam9c+OwvTNWWzRxitXosdfRpJ6ljQtkmKl2FwZLBR1EidWrF+8
1vmqs4elDavQrE9g8bxVs5DpYee5IFzuEn80uLZ8YmCAciYh3J7Iv8o21vPf
ScS63g6JPrIkkRTJ3EZgPDC9YUdTXtaBj+N8hShTPp5xsP88WK+a7tJGSVSJ
w4G/Ho9ARKy9EHaIdqx/02tNen/1azXDQfdWLIrG1xCKhAbySi5mJFlyf6NF
wcLAoBlYxJpBYB0XM46cdSXOXZzmRbLBOvmjAx3ViPqbzc5g+6ke/8Cxpghr
dwgRo5LGUkZ2RFO62sLpECZ37UWovYUh1+ARAuyBWGYsCYRjwFibn3t8TJnh
QwzcEw4XCfsY2Qj4Z0QcMTA+crajDb+XPJpk3HGbr3wIAsQAP6FE7xW+GvcC
FEJzkI848zpuK8UY83o/TRhL8yNd385x6XEXfNENbZU/fulrhxhFD0eSJB9A
U92loB2q7txxzsdyuoNtch9zvHzAtLSkW04j7c34y3q9kJN+pSNrPAatUAE4
hvkYrkaq6jqxckokw29bC4msZHLIjRhqjPK2nhgIQv0oXQ4cvHNgFp0lCY2x
NwgUooppXflKWfENbtkpLuPdPhQgprnzni62yMpeX72XduoOP7/us/OOuuOJ
wDTi0t4C9Q+zctnorz8l1zcqmVETccBDkaggKlSLLrhhFGmzJkMeUKTLTBNO
3+maVwoucpX8tZbbEbMRnxpv4PTzJrt175Quzdi/C+OJfaygguixKRA5K5KA
EPdjUxT/5ozj0YvCSalzZcephknbdOLhMmNPl9bFcZsu+jv/JYt2fUfZM31X
ZmYPY/HEh6JP5+/80waHtgVD4FsyIZzuOskfuApp2pKATNbLpwCYDUlw62BJ
RagYHU0X5Q6kPK5M8QfAgmFkkFe4Z678BBka4yWJl/nmdCrATYO3/p8FbeHS
kMxafVveJA73vXegge0SIXqpwc5APZe3MvvOH9QIpXkFKLtvpZ1lE+urkqEZ
RGhbpixIE8RfYppDYpox8SMWoh2WJyNHqr+09BqHWr1JPEXFbGZfXVmsu1dr
gNMDygzUSG1TYml9P3tm/PP4CgjhKqMVy5GxG35op8KR8AuNFBMqjgv7psm6
aElU2dnuaZIpYsAv2KdmAUPmDtPFxGO7qLFpbKzOyDmlQYH7yW7N3AxK503g
ogavnmvZ8zBWoRFd2vbsUSZowRWlm/iNP8yKtCMUAKh9+bBS9zV7cB0wrn0s
ZDOJ5ALJ8hGVHJtEYJauHDWW109bDhBQUnMaIY2nq/UGmmSxYYmy4UOM9n47
qQxWABO3sRW1QHd4wIQ4afO2/VQGw9xMzHjCo7iBy+WpHXWyK+pzbsbTHmrU
yG0bOPnOvdSjENSzrlT27OH/Ert2GW8SWTpQ9Ok6lSseRNbdXVr+1jft0dvM
ZARaq8Udxor5sjjqVjh3Z+xRIlNfw4laBUp/xxKO6QacBmcpfeXgUQh82y1t
z0RfQxKjQ5DkGZqVLgMDTQTJyI8Uao3a2KbK96QcRyaPuuFIPq5XUZuZfSsb
68GsFbfIKOQGfzQ1M73JKIIMzB36vscbvdW1KZB/Q4WHo1m/uIVYm8Zljki9
4ejGnSNv5nDO/nWZ2v+Oe3nmwXVML3ouXDA+RLMpkBf9d97v14s7lUMMThTu
zhMQAIHYXs3qjzTRZWpWANlwEcp+Nij7Oubh+F3iA36EVAp1BlB7r+aFukBM
wNi70ghBDF+F/GCFtw31Y1e+O7+BOB/ByDvkHzPDcly3i07e/qpewSXkmPrH
M5/C3732TX8tNC7Q2zzHk5I43RfmYU/wEfySa8cHKDmYNcTHeeFlAZNMozD1
FSLP1eH0Mdw+TFr7PjVgZx/cgJ2dTpVPVnHlg2vEfp7FDYnrRzmHwx21btJH
pIgbgBRxAE03toEQ3rR10ZgMrevY9FCWyTQy2V2uF0LY0pH8/IPiLmb0Mq1j
B40aPYdpclz1ahYYy81EwQFFKI3ZUXC2NEz4xSTTehewjHi6JPKIZFXSSkHf
TrBFCmJ0zjijbOG/YGgoR9Yx/86IXjNCNIUG3gIRgf9qG3LUaXXlAwHww/ac
5Oh8Bs0l0UGAXDy09mkZ8/YGm205E4j+OH6mLNoxCJ374XIjUcfFkczC8yG3
4B2QZXE8ziisuIxEbyiRk9gyG/0X8XAZQJuBGVE+thJlrL6wgspD3Xa1cJne
T0Wlumlsg/YOneccxbv4t2OmIFoBA/rYNv5L8TluXYuwJR3PrxUpVAteA1rC
NU/6WxUuaBYIcy6KtYffF0iwVSzogY3/hu+ilV3kZBCIYFKbfxX+DBq350nD
EvjPktBr9lPbWhiClsSSgcwVpoTuLvi36vDAud5Vp6uqQvIP3YfbgdAQ25jf
tPKNUHmL3MlUMCpZRby20heukmlBHTFpt80QPaUUevPwRQTYXnvFuSgNJlti
ISAf06tHaIx8wasCCTxddTu4CGMcm6Shx0Ed/Y6PDkgp0mIPds/1fit2uuEK
pQfgOGbwPXRu82hPlerJkUbzpRcZAHHROTyf1wamMHtPC3l45THOuanYYoMH
HHxNe34thf0VROAMylcODSKu0CGvg1PW0puBJm7lBIj3HWy4ibR+0OsvIUff
9+GDgi7I+qV+G1iRv7Au6wvmxZ1G6v1ptV8EiuPXPQYbmMYoGpYZCiWll8xy
XSTsUI8vQ1RXehQfX3oh61KzwJpCZVO6er8yPStKKxF9RuF+LKA7PVETCzk6
Gh3oclYekBMmANkv9hXwvc0Wuljw7UuVaif4MFUGFrQKeUR7WcMsyoF69VDm
Emg5TayGBInJBtQRtwJ5Z5L3sb3+nXYmwievObjITz+H/bfPoGI2vVD88mcr
EjkwBcIdYA61EkXx3RUq2WAxMOek81gjyO5bEc6hcAkNaaG5eu0hpF2kgW3B
AELYBoXjluYtOxWMo05G+K9tsnqU5Yk4BMHAsjbwfZ5dCioPzosJ8tIAjhuh
85JNFmMWWAhHfliPpOd5+twcV4gN/FYNikKRzUykRSRxsWDClIO88xWhngiP
e71kGo0N2CMi5778T1FQXc3hxrhbgCC/E+CSBXpGpzCwBFj0Tt3AKHPYDvqY
oZffs10JYF9l7bh0ppH11aX1A4Wupt1faCxe8Fay8N5GlDHSv3gxeC91Z2vL
hcyGZDjXR9mLaHHO4vek7g9Ej5SrkD+ceVss1gunT0OffeyRIl94kT7M8FTe
1OFiDDY4LzU0eXdk7aKVKTk5z7SH4s7F7vWwnR4sShT4slAkpPFpn9dD3IPC
TVCJdCpbR2LjlOLrthW3vHIkxwffRVSQBJ40Ql/tNyU86Oz291XXoLRWfi3L
ZqsT57/hp5AEL/qfeFD8WOdU+UPwXhub1/nW1rjWby5/vO7X6zjQy96T8vT/
Qns4aJl2eQUsK9dg4uMOouiVOwBYa5vulP5zTgYeOaMhLwTz4bgGCWfvHoMu
1MIffaepwXCj72k1+iljsu8y+HCh2PQpKb7MOZPnTAmzKRfZ8/LkwDaS10vy
4NG1aXEyy2inJ+PYdGN6R1hOGuOcqOVVFgUF+6o4zpSGDGjfyjD0ZqPd9rMm
zorC22GwGl59j4VBuu+f+fC+15rXeI0uhyJXauy8npU3Pn08kXt+ccF7me0n
WrimQkhjDf3FCm6Fp0rbuc16mzmxM0d55koExnFtuI3SpkcMxEfuc7fwArof
yfaNer9N/PRm3Y8cTkOQxx4TVrkcxP8f2DXzlBT8dsL8YJS46lN1BEscZ/r/
hj6eSHQCfGWDuaTyWE5F30B8GgvvkZ/etinJq1wb93K6/MGvMYs7CPQu78qH
PGpNnYynJnak7h686a3gxvUN00kqHT8pLWu0zpiKKALxDnw3EFxRl0xvxIgM
MXvu5b09qeBhwgftyUYdrIM60tGG34oeH/jDUTsdWuL8FD1kype6wN1lmIV/
SCKsd1J/jONY6wdkyKlJAnCxxe9xvgs9d+ll2ctSlMiSq9hT7+5ju77AYppK
0gESqV0zYWsIbq8XmE56GTy/Jm2vpGBCk6rHcqmlGs3M2tmJNWLqgYsth36u
vvZFRaDl6fsODK7PMQSMSLzqiKg+rj3m/86YCs+nM8Qz+Y1FM6FKfYxjvrjE
b3ewyp4dTBXW4YbmI7k6PsQoOF0/K2U77KBskikoI3QhMGrCmYV31ZkOtAIl
ih2YX0bmbT67x3dHYA7P+3BPYzKCjLGftDw2+Sy/8MorNab2mTgS1tjz+aiW
XTdU2/ZBDh0IWJKYROAbOuu29h79IKJaLCsn9Gy2De1z1p17ohf395IYHcnR
XvYiVc8bEcAUTo2QdZD27DE5Mnj3XjfYo+n7dMsHUKD73lrPdC63DnyLxxiH
Bt/s2c7iLH/ZbfKpNL3qd/hXatHbAef0riUtmG0xNv32CRIr2ocNaG7uQ7zE
40OmCsuX/lW24IEHAYJXQ9pb9mN904jhv3wB/wW/DcBVL1IL8WrcPI7cFYAh
Zmez7hPWRPp4+AtFYQkXDR3uS3v0moT3kVXYlxVNRnNZ05Wt+b1ESv+iX4Uu
UeKZkl54ozYm+SYn14kvZfxx4lAj9pvgQzbaGIqPrhs3e2vc+SzCtF5Hsj0C
iHa0FSyKzDGikFzNQCwNqpaS1ooe//M8jh3uKmCeK8I14IlzlzapnpygSdre
nFV8sik6pDdLUrtED8KyMZKNOav2P/aTOSdEG3rtvxQ2uyDIBQt0xfeJrtMz
fT700RIRb0eLgvBt1wwob6ZEBd/AuWTilTIkeXGZifEezQUUdWM/G8D8H6MH
hWFzqAHRJkBNBS2rdoyJBE/FrT3PzHvsCDag2erjeM7wQHqvojbPwHfdkMdY
STtXLvsTdy/GUufueIDpg/ZQsUpS9O7RGXcM2DtshqKwNSXPG2OGAysV5AeE
A3gxnJ6mrvYsXPM8gP36E6oo7umDVBKHR8yPe1Wleu/km0KvwjDIZxE/jqlW
ud0/9zo6hZydBiYn+JJ9lDj1d7p9q2zwbIDkI9Z4KtJmC44SD746z5kvqpsg
1gJyjoaC0BQznnZEw3S3RkNoIzWmAkBZ+gW7JIAlVfhr1e5H78q4qmssWEFo
VqGg4JcGqozW8828IK0X9aeTeVy5LB7Yjrx2ak26daYOvaq7IE5RVg2fEusw
gfPApnV4PmexI4LeHd5Og0cmATMKICw1d4ZRf7bZeColAPgWwUCTyY3XA4bX
vesUyjHWeDKqr7glcqdclXOqhoRh/6/E/p/HYXE0ITDWGBTq3DtfzCtzyLas
m1YfiYmAfpCso4AXq+7Fhtq6D4Og6djGZbbqwCYQ2A9G/BHOugJG12121wRY
Z+w9/7nXw7ya7XGzgdTUg6zDr3Ej8wHVi5Y+geT/btDKwoBClyrD59pVuGX0
wlyh4vLupF4BauLlzG75LQBibtF4IGZ7UdnJmHM3vvlH77k8RWP6CGQRFUuA
NxkjNQ98QXpyPSnztFL3mdR3Rx4U29y5WAnW0uM/PRHETxJDA3Xl8LWKnc6+
M9bccsC3FfJmBXy7go5pCT5Wk8zrGpb9B4c3Hef2jWhKMrc+nG0v3aSVKYd8
2+mbeyDIVjlYTOyeniaTmXtGdbxNRTQgjV0JXa4kGzS+n+PJZHfSvP+RLOud
PdOz+knV2eqb6F0A2KFsqvMn9eveyWqrDkjp1eN8c/8cgSGjZmHG0i8cRABW
ZstScfyFoMH7D79HaRMU4/9Phu6k9EaK9fRuHRC5xy5GdND1l0JnCpgCrrGk
adthoUIU9HR6kQD2kEapPEa0EaOO9U0x0B/Q1PntOBK3RWn8fBfVojecg+67
ukOMBh+4pQE9oVReb1q+7FbXfg6BCVRMz2+EDctHIpYkjf+JK44rIzNtA7Ex
KjgrqyG0xDE6U7PE55CbFZi6pA9bjUX5E4BCH9aMxzXpNRbzFllE8XWG//hi
TQRu1Y5rqjZXuHn+e5kpWyaVJiUZHbrF+glFZKBP5bw4wCdvJU9YCV/IHHks
GMmC2S4c5Qs9MQ/+zZEVPHFJRffWuiUYKZ6BCfRjbjl3703vpThddQGVC1hF
opfNafXtgS8CqeSy4O3uZM8afJv3r2p5HjWbZD/kTVaDCKMmfmnM67fJ1LDY
4EoiLZ66518L7wBbh6KyIpes4VPBd/UYB4nwwLowm61VD3I1isk9o3h4XsWu
8e2LqeoqFcAmp0AZyT770gcDl5LOXNEevUkFgTIpnDBpaAtpm4rh9fowyltf
jQLzRNC6bLXzavu6C10V3t5n2LrGH6Tl/tUJUE1v6QDQtLJupSus54BlLXud
6VBbELUpOTmODs2ap1P85x0lEgHgJIyJEJ7syMBKTfhabUatKri6BnMxwXg8
zjIP8OFufCJjo94iIwIf20zbG65qyJ28EbFG6Vqwrn9MU+FXqm3acq1cmxgp
mhiCEnAa/JPnubTyBsV1KJQclkX/Q1UKbWAaylcGupPqKB0gsa5ZwILO8ELG
75p/Hs9OAxO+MeLQ8a89kVT0aCXOFA4AjwxVxd23iDpbRnb45E1DNPkEVoym
KxFYG3SftNo9HPB42oRs9AqQfQHfTI+FsdB/ia2OqnO65/xJNZPKZqAcQdYJ
2GleDB5U0OSZCbfj3syuMETdYWC9ScjmuiRrzs+XlJfzGuSr26z0yqxNY4mK
mPEEmabPvPFh9un17k4dwUhtSJeHkJMhRcYecgLNsYGxs6dJIUME6c+Kobws
SndxywIl9QnoySxuDXdPx0o4A+k0cal5KOKwKcVWSbOlY3wLfbbnReYYogsU
qxLzCgdm1VVilbxe63ZFn5cw6DC0yvA2LascMNbnjyEFIs/W1NSJuMk+Tj0P
ELdfEEx3X3ZQIheT4VEdikBFbIYTsFU801s2j4dOnu64i+rmTVmBCpKNlk2i
R6VXqrwtFJOoAgnv8hCGk9IsBeiTSKqO7VAN6PJ/+FjhO5tlp8+oRb/06YCS
xFWCqJg6div5HVqRtlrs0kGwlYnmxHeP/PO/dOd4SitJN5pra/FLJf5htagO
/I9NjA1VA5k8KAVB91ctJAC4AuDi09PHoOxto+V+FCZLY1WMMXIqCM3QcxjZ
vrYPJE1qO2JFP6qqETn7A/StIaMNqazVeC4t/vVw8TTZawbQ29aSnco5Pjun
UKW4w+VTOra/4imVm1eCRuMHGDHyc7JZ3TMKXiOurmnRec/x4LD9bVFbslh0
CN4yesS7yUX5V7NRTgG/0bW0b1eA4QqhIo9qpSveIhhfp5aCry+MU+yRUox5
LlqK5XSv5WdlcnBRBz2s8zUJmltQQkw1/yAYBivLgO4LX92+1jrNLeG8/g40
snd3W2GDlccYi1b3Ci2wjvIsFVRUazXcuDMTk6UiMHnwoM9wOkImIT4cXOc0
k1PlweiIrNwQshFIl94ysLvXSJCrk5N7CMm6sXQYBuf1/2PybW9a8dnaSS00
9xAT0tOwE2yss2uk0kDnEr9a7TF8z7+pW4yxZem7+NFlCwWSm0h//Tzt8wLB
7CuQIuYQlxiD8LwmpGaqZt5VLFwGZdNf2ynagiK4vWfp0iVV433QNzmFsxVp
qEYOixCnIM3BLN6K17TbG/xvcn3lJ0vmHknPEX+zpMBB7KCCSbc0XG1VrwaD
S0rafdoruuW4e/IrLdxh27qPcoXzxJyOxEViXyfcAw97/Wf/8YxL6Wcq4TGn
0byx35KqfbVefs8qC282Rct41QfVAMoox9NajjFVapOdwaI3+Aji/JJMD6Pb
5Y/vYs/EpKAOvXu0BRbv+4L/x6HHwZgmOaAICc6zN/jv5ATNhxXcy27AS9OP
WKLjpcL7cS8IsjRsqbag+oQPgzvhVo8IhqAEGnfGlEOAnmOoQkL/HByQ17AP
BGTqHLPijkF8tK4SgNosZnULpQaW7LntPWoMsr97XIx1Pl7fozCcOgu00BYA
HjLePujA9RVI+orRI3FRjdacCUTMwMqf8qw6c3yBabfRU9yZM0LBAUZoRzEu
jx07eq1vZYZxvtJ5DoCCnKFoCO2NZfJqpDgQeBJZwgBhG8hjIlLPO/TkZwGx
u8O8FDf44MeWUqGrEvqFmr53vZ4sTKfGDxXIaR7NQB7MvZRsl4ZfO4b1Mc/4
em1WYT2gPot3FbVO8p68MFfrPgqpL47XWy3d/qYNVnbygBZir6QOpgJlXU0/
yXQzydo1nTYypa67Wpj5tP7x2WO7iCosNAbfkFyYn2alx/AUd6VWehmHhQ+Y
6Pa1sRNMjNRjWySTg6q0Mcrg7HYsMYEK2Bay8dw8a8WRHdCLGeQH3fnlMEmt
HVgm89VwhAdL6CyLrDfhJS8EFcFQmiJZTvzeHLKV8M4PO1He1+hcyokD3pFA
FsggxiwKzCGbr0KuEQTG4AW5yUxMwt2mK1om6U9vs3nyjb9i7NfOvZEB6g+M
s4cYYFmzMwY+6WveUXIIMOPvVILUC7SwV2k24Feyr/VTgxl0vJxbNN7rjQXG
g7lX8qzn+D1kmkmzHryZpn8qqyMLmC8bQZBz3K2a+jII8nURE8LtiuGiV3aL
uMRq8uHUHvw7nTShbr4YYun3lM5cWo7/p+oPTWH1JL9AJl+AhrYFMzxyplI0
beeTAP1SxcLhXHba9GXk0h+NmFc4XuVovtphZzfoLjB0h6oPpH+Czb3JLJ2r
yY/Ovzbd5QBlw3OHMN5KFsSVt2KakZ6IBRDzAJ/7qxwd31smwx3x8lAX7A2H
ccxLP1e+NLGYocptBoK4l/aUxzQ4i4Uyv3lISxTmFbDTSiiYpxfgHzzlnekz
KdW2Q9NVzId5SAK8X0dG07t8PoWvNuBrb9XRp15f55Oa09dQ7z5C4TexfWYv
5Q5O0INVLAHDiate0lARa/a7o+Ax17iXvOA4Lzme45kHzdwnhIuRwWMjFJ5K
aL99qS4eMIgqSzvUpTZ1xck1YJUQmP/cyNWKLHFOIPVCMLA7D4E8c1vgxATp
8kh97AKNvwZkZNOkhSuKj5Z3b3l2iARU9Kj8RR3kF2R4LYis1dqQthQWe07O
uBSOooSe+kMP506voIeLe/Sf16tUz0nJFW/uk+5ri5FtNuB8OYVhhwFlRpIg
AB0F3lWjAysIeZc7Gw4sP63Ucl3fN2xsjaJWOi+uieHqBT1SPDOYPmW37fpA
I0wx63f1RsXLZdPU31/YkTx9YnlsdIa/s+GliryXNlG40nW94/JTXKFM0A9+
s8m5yQ1jwv07GsY0H3CSFLuN0g6hmKXJpA4sDpAzM01ltcg0G/CihBGDi73c
uaYwhOPER71HHgoUxBaQ65aY8p2ovuqlLzcPgKnsWhy++Wc7UA7DYVQFKwJt
JVj57ib3zxcOXm6XN2zIP8eu/OF0cZNPPgy0uxK/FmZ7FiRqCkvWJsRauHOT
FBd3BaJjAaBBNrwMv/oVObz5xM6xHYyUTvAPr7T7XHV4yqHxigsdDNB1UWwl
ceQLgm+MkhiVZUPkRU/YbyD/XguC2GdwjLjWZLR82h/NmjMUxoKzpomzC0J2
rZZwk8nnnGd6T4+U135vT6YNk1uSiXi5Wflk4DAXW/sWiVL+/U8Vcuz4sWad
nTHghrfYCJII5KgiR6nqKosPJm3tTr4EoqF9YiAOVNDi+OlVWucVwEJYJ36w
GAxjNL9t4qSUj4JMAxFrxekO/lTZeaa1Ivh3E+2YiLiqfnUu6bKU0442oIs5
6rQiisqAX7UCcnmBZPohEsxnjpUPYaNXACHRYLcbTnSMqc3kS3L5yNtT+hZm
ULS9MlLPclqZEISXXyijsKdeuutUX4pY27WFmdfUh8VwF0NQhv/CPMvWrju7
qxMrSZ5/Op+zwTcgFqKkcZVqCFmngtf+xpTUbhsaRx0TVmI2q281+87Nc33Y
7PU4eGf3eWOXhtBx9HCnnoYzZNGwR0cyZ1I7QaQLi5Kk5pHPjOr81B4ilL9i
vgpRBl85mr3Mlu0RglWUYabMigHNFVV6E2lgWrJ/uQ2AuIPnGSVwUauYuJgT
6dWmLeBmS54ZGAlrADzjX1Nb6Ru1XsCnQ6Q5A4DHKmlN4frVmO5OtteaHMY6
g04g2s5qvvcNBRKz3FgQninQpAaWr5AWy/N2PYjTfsC7p6OOPTB+VBptTtyA
QnrxJJn3/lFMZKrwaj2u+uGQNZM5wDBe3RiEmB7pWhjo9Wb6sVm2CTISPxiD
KD6gCtZieoNRrfmvqur+uNWxyKVV9bWnRHgD1UnD2Pfxwjb4grP29fOWjqMH
6LbcMAcgVgmcBGwnoxHAPu+HDjOUYV4XrEz7OuVU/98/lFCuSxiMoQ3EQW04
PlGEbbaZ1nta6/CWYeDw5xMAwTutlQ9A+JdHjuS4rgjBhGcCBMquCz3qhRb5
L8p6uaDLfgOk2sjfMFEO2f6Gutnu7DCEXsLKaxbONO2GzQBRwiXoGKi96+6m
EHwLc7sWf2dg4hmAld5jK2topU5/Zwp3uao9JxjCGn+BVBYWrRuAQE72ujZF
TaGGzX67TSLmc/lKAvE5o/2y/QPfHBJFu+vBe9kd4A1aBRiIdeL1b8okiXt/
ASWKzBzjWaFhZup6Uq3RynaaEKnsroQJox4gmaQhNq/wS57uuPdsP48SggUi
r3O6ptpncAyDdDbOJXdZHmGzIU9lHt+8OXUIgn5b2J2nU6yZ+PHc2Xx8EZx9
HvevtEIqUJYxqLpfeYmpTb2LqUVoVI0II7MGwg5Dzqiegj1G1Fg5HBlL4jkS
Zq5n9OBbwqiZ+yiPypnrPkqMWJh2K7xE+ffg7UPphfcLPoGTHwdsS2vgr5Ab
+m3aUIzFkn/SfK5JF5h2sRZtA+LI0Kc6JKH64q6+zxUN5Uy55y1ChbIXXG4b
2yA/p2+Nk4I0VjbfJqTBksTmDFNKWlaGPVnx5zo+cbWT05pYQ6yWugLdhFMj
Excl77QupNWGZz2b5Tn2bdtWKtcsJPVkYYwwie1zO62kIFyj3yURiW3sHBRe
I6eqKNAGyuibvLbfHTKCpMF5oLmjz2CNQwM1K2DxX6YzsLfneuJXevIEw6+2
K5ioE6YCZtcsWhLL5ZBdHMO6XMVPRfXoFwixMxoTfd9m5hozTUgQ6ggLH0xS
TfA79uvV8lT+aIE8PQBa5NU0kjA8cf4jT4B5msfT9pgdWeJvCxCGkh3uP1GF
k+zLurc9+xW+a8g+hgXjkMX2+FW3kG2ncJE+tgERAvKezPxRS4h7mT1ZdFDs
LZU25F+5RLUp3EKpR/lR2KZhuA49/ILVtF1zs09P72rfRk2ew10heIuRx9za
YltD/gwQ4eExTYkLQNhzHuRzm/QG27CJWxeJwOuG70/zQWq47guIA8D7MRSr
vTC+3lBjLwqiULdAfQGAZ6kCpuquvUuLP2OEG8k++jCt0tESChdLkucvQCA8
QfX670GCaupjpVB/Ct0uc9bkqQL0V6pjYgol3mpkV9NChNqRUEhZwAgu4XlM
qnUr2r+bkCvc0TstEkrUe0I7y4HNuBzT9p/ZVH+1/V9hKJqlq+APj0o48ORF
+C2funNi9m5kprE/XMRnJvhN3zL8uRbDCvTRDpLyt9APHTAAqSnbetbfi3lZ
jbMb/2YEIq2w4RoPr4DDn8P7Lwo5D8HQVFSlOrrpeCD0uU0res9dSoXTr/oI
4WyuCk5lOApWHEJJMZoCDia8dorzTFqTvinGLszGB1ydgfyRdNFyx+WLSmHw
a8z5mlSkrX1fHnvGXpYsmT1Xotc4zHNDRs6ATemLQ6/cAnRITIGAe1Lo/7OO
aNMLXRXx8+9MsJZQX/q4CM+zaaH1DXqixSD989c5HcW0SHsSEpFV+oc/NEXc
vWN/BcXR4MH5fPLWvzOrOOSS0jKAR6j6TRA/+yPACNTVQ/VeQx8bvpdtuoZM
xV4L0VePZaTyJOARuJS5mfbY7PvrLEWAF/zzSFObAkKeN1msqyYfSCBMLZ81
h1vJwE2CWkGA/9k2+g+J6cG0Ikv0Rn5Xd5RbZH7GsEB3fyxp3vLpWv75Bvsh
Gyechm5k4wQtEqMQGrtnJbRRxiLpd9GFOI9+GLxCtotaDmwRB0B5IBPU8Qzh
q03mWFHq1Mva0xuYsPuQ8pBUrGbYOJSI6STbSUTLYyQkm3LpsrYPdrPng5jG
sRqhPNnY1rQ43DsLjqTPX3tv6/TKvtlly6IO3B2QCCTLZ0uKE1m4hZB7dbHc
Oz8n6yQPaDSJExMaUHTSe6kzdFl3Kqn1Nv9btzuenRwSnQAtFYPdbOWhNjt8
MEV13H2//vhwpCTaRGACv9jrS2hr5qsEm2yF161uq2PC7hi7ZNy4XmgxaEJf
fmG7cNpVZta8TOvZY78/IqGtWthljrWcfYawu1wPPq1QjtZxA7qlYkxviDJI
ZR7MWVCItduJm7vSxVRlTT5aXHVfb2iRIYUleZJGbFm0V/rx7sMhXhI0Gc5Z
L31mFOjXCR5rFCKgBAo31dST9kGdPDV2ES2jhw24wRyUquZ9aN7V9BeKVOPY
ZH8lUkGihW6s1hIF+ioTTwqSS42PsU2QJS5rla+U4clRyklO/rE4O+lU1MCX
r8JuGVJljAqCJ309LW/2XfzyQJc5/dYVw9grbmZruDvfZzHV1trMWGuxLab3
IrzzrMDlZWTKd9s/vLuyQeDeJCIL3Vs1SZYFNzyYfCWY2C64R5X/sMVMSVVZ
oKjktHaBRVkMZQ84Zlzc3B5I1Hz4auTVWojDfagqCGBS1phTX9eyYJuwFFmW
rLLQBPatEFgiW89Q38T+SzU5t71CZYLNGLDfiJ2d4UHSr4pdFvi9oPSEnAO6
xiTFAZMh8cH7pR1BXujHODyEV4S01EQRVetoxXF/I39cLPXKBXPlNdcnbr0D
ukIGyk5+9JskxRCwn11L3WhOGmxDcdN80US+XnfmdyjBFbhdvo4lpQlWmUAH
JGd1Pr59VO/rzNRDYBrxUnqSDQVRDDDB/CXO6KRQGAaLrN+z1wFV62w0kXWK
yBC2I/mwQENlhxM71DtqcIi3+DCWb6rwt8rb0jCfkV9hK74/tJYdbk6nOzBb
KjvUsICQqMPGlg682xqLGBEZu6m2cIZZniU0ypQ/Eh7j5US4V57s0jiS9PAp
jtnJiWtHjcPbjxXGKdCr3Jwzgw/OR8LRTsgfH+qQhGBlips3X4fit4RKTGeo
gWiU8y7zsXWpYfIcTVnFsgqLgfLYq3+sJNqsfNUEUknkbFjBsou4v4bYXp57
5HRpAuO5E32u7uYeXM6suLzlHUBWg6NJLtSRQRfIGWHX4sbEZB8Nb6CbwgQp
F2oXiUQii7hCcZwTCgdIXVKzS6Ede6WLQzn0jugiLiaGTecXf8YD9DMgWWgj
iODidUHUClHxDaXbSRQaVDf+e/OyDoPb58PqzxYtzd3FNHZtP94mJbdJuih1
b5u8c83BRsZZmnJQy8MQfjdyBeQxDYzAQlWtOJbDVVHxfR3GFRFvhnoSInva
R/5Qs2+CWhC8zxXdSlxVuBcs3nicwwUQWed/4+945rDA211yUFEAkwSM1DiJ
ze5hY5fLYRoIQjsk2PDb+zfuUw2b86Sx7gzKeaDRiODLErZPcrnU5ShfIbZv
AEg/KyTJXQccC5p1egEkY6mSCOQruZjHTD/xqs08iALmTD7u8TdTpRnpF/Ho
dkdT6YEGWUA3xTu065lxkNfLQrpNtr6DW5Jm61zHY9SqioDTvSwxMlUzrrbL
XTeYBTR+a9dIrCgmcjT0DTWxZ+L64Huzw5RcncITy7bhCB82ZmipRYtQtX84
qK5AfxWnMboqxcfMI9nkktkBL9uxH0BPCIixRk9wuQi8Ef6qK9r9sC4ZTSCD
TAX4mEHiSMq2RcOPPEBU+orQWCKtAMBVDC4qgrtoaMcdeBozb420wHh/zlQW
oWw301ImwFjwd2Wv3Oey5YDlmmjipVXut1R1uHsSDrQ/N4ljaj0lh8tTxqTJ
0hugo470P4xYB7SQP7MlvqasMkcVrKYlaw2MRjDSIuHV9p/maM0oWC+YnOw9
xSYwUQqdEaK3IV3ve7F+l/6EhxCQi//lHi0F8YN78bGjyDFyRDfYQxOD2DEc
Jy3zZxlsoFLUMPsBP1UUYpZD0WbtSkX+TXuh/15tmoUi3VKOdw8MShWYfgkP
lnGuZW5yMlfEbSvmzLDkgj5mUBLeONb7QvvDfUD5O0576fCG2u9vKHbE5q8n
eEUsjwetDLEFbzVNDPQPjHbj1wRV/6oS02pJPclJne1+2gePRx6ev4QT428i
4a5W/gvbXus7JtvhTvE0mxJZfUKg51Dnt2FXs34lSPiw6P1zcmWIP94C+f6z
LuKpVpIPqct7D5xKRhiR8f+vIlRj85IuV1IStJjyWhFsgD83FqizNjhLgCBM
fBsia3ru7Wv9ZdWkmR59kP8U1+6RXvIjWQyhAFPK7ZRDfxRFHkua7Dlm9VJ0
AMU9pDlfwdUDN2/RyX37kLu+F0FDB2CweZ0MJ+IR17O+MPyug2WBEAmSA/iS
bbKS29hEv0dEOPHuVBuqbdUCPVdLUJZiHjVpaauq0O/jGlRkQa3kt0X5DX+O
s2jwUvWntsoy4eUCHdeaGecr7mjnya7fnE/cXcPardam1AC46cKaX6dydnHg
rrhL7fQM522zN2DQnvwtGdmwayIwDUw858jBUvmzk6AmFLstgj7doyayktWG
0sX5CtdhnO/PuX6wBG8+H38kPa0TGAIqx89VEfZ94oWgVZCLlRbEYeMcOngW
6ao+l7/VtcJ3SMBaKX8snbbLS/hDVXCscRFd5xcZGjdNr2oS4zbk+f+QevlQ
frhOQp/ktCWOQjgzsnu6Sj0P39r3d8f+yuJkUIfZiVnZkMqYLLTjod6T/MvA
Br1HcPo2GG9Q2Dvfw9HDg3A0ptbINidweqc5+eCn1xFR2MAqVSV6WxWNuz4q
nPzbxtosN6j7TPox35HmP6b+ss3CEGNKSWrIn6l3y0xbFNzLujKkfVs/tNkP
xeSPutcj+nTg5clp7kyrN2o697hB7/YZtSpB75wy6Gzrqa+AguRiPXoQA3eN
d2gMc1petmDMLkViwtZ6s66oR0a1F193MX3qutIxcT8dLaXmCKSfd/wDrWEl
7XED/TaaEaF3hl5vLyO0KB5wVmGlVtB8v/rk66nFwR4/7x/iw6edjr9yGJGj
uTiqIYZEdIzq3T99gicjugXMRvsq+M6wSH/Wuq5qMXGpsQ1ERSokuoQULCyo
MhgHrSnI2qHyJiWAoKCqQhl69/WPWT+bd5oaj/BQBteA+VczJ8YQMsDrSOo4
hiDZoQ/E1vQeleE1IEGcFS+8FLxKfeOWrAuWb/Zz7ZhGcASqNUvHkCRYY/zJ
6NEt7SA8ci/WfR5/vccK1H2PcnkB2mr/CU9dTpVwjex4e9R3ybAfy7iQpd5B
mCkVGM+1jPw0viyggtFro2mMQPXt9FTZH2azwlEEFyvX3uA83LQmUVZJE108
ShyXd1xILOkGEFeCQjrK5rhbnj5OfEz8LLcH/xsbsU39rj0+T0PTnUdQ+Gaw
5HZf3YgS6zczrsWtMyo5P+LypVuboL15dDUewFkmnfemd3qDmJdWd2v6MmVx
2TRxYatNrV/B/MHAPuzA+Zaay4rXSpLJUHm82iYOLCI4FLWCO4FAVegFEQ4t
SKDz0Uyd6Pj1ljPrJpkFhC60kZegqn9iBHF9fOhGrUSAepvIEd7kEKa+9NuV
LW+xNcqvFS+LzSEHpUx/0zyJyZ+xzORfU1eruyJYx8qWMOfBURpVkTAG2J08
BWmlXNosDJITUUwzZxae31/kk1xJuzFQxuQ7urs6/YDToyscoLMB2vBliKC2
4DO0TCRliRsTzHkVLbgLaAcYeUyrJms9HM1DQvQ1DN/whv9OkL11CZjz/fHE
jhjPOgXD8aRa8Z6A9rEBLNj1OsD7b1BYkr3hVMgg79hnA5nf4pAKx6DHUgWh
9xy0XSFar0qyg+87lJ8m8SraZuR26PhkpYUA8JkgoLmESC9p8nbwoAQyoWvG
FVsU9x9wko1Voq3C6u7+mxkijvbPIKbf/g8ZpECXThorAX++iixOHpkm2IDY
ihqgXPSnhaFyGXMYpTn7QzByf3KR5ZOhAEyonTGMa3ESuvgGx1wtGBDSIcth
PSLyJbl5KWE1D9FdvM+IyejJePQrryfzotzAecRb2giuhmUNqEAu7A9wUiav
v8qVM2C5AZ1STls5/ZS758slBCo6+GftOGMHlhUwPq2a26S/32q7J/enkyMw
T3k7Pn3S8eXHv483HXf+kh1FmjPGsR4sqgskVfZulzbZMu1xViO6rkByGbX4
C03V5uO8bsYFHHZT29scqAdjq3BnhhWB97xckWXZEUDfVTqYxqGllfoLNN5M
lNZX0gwzhRpdoBG1V79VBxJUcNgUgZh4Ge629KzsBu7oTsmETTOzT9DuB0jW
EYJ7ftKQ78Uxs6GOsDlkeBScsQ2X6TsndmzEd0+R6qh/Zh5udpOQTyXWKhf4
4/qElppOsAUQpDzyAcoNv3lPg30q1jUa1icC6lPgPJFKHWrQtX5yira+s7/M
dfhrpYqOydD+axjl1pVpmvTX5n4tMnTQSudH7vWNp000PYpQnulx41cnxz+k
ydl87j1ybJt8ZunDRJw+Tz2nR01x7rKj0WJd8bPwOqkWT3CuH2cVGiJk/kev
j6wAxIN1K2GmTMdIqBZFhAtGZm7Vae8XJbb+hRLe6woZ48nOzvXx9xDGFS5n
Mhvx81mOVM7JfiEocyNz3kMf1ea8P+EhKOarC/DA6Ed0P8O3JOKrMTmZdASm
i6DknRcv4NhbcTjIguPTLOVmX4pqF3uN2NMe9/vYxRlO+DldotaevNCRoRjf
3N+JG9875KEpFVLzjYA23op6Fr7aK080fcclBlTpKbR/lpwpW+v6RIUZXzuR
krihei7z61d4BKE//5f1z+8GULTiysBDWiXrIhzt5cwJI4Po+BhFhJQfgOs8
s7eoazAOebDEyiMnxI5hlp8c0l4ty9h9Si/2ES2NQrFwypUVuMyW76YDzpZu
bO05m66BPg3XpsLsTPNyEB+dqrCabEjDwMAF3LVjlgxPgG9uervXP4llwmFp
17hRNAmt/pylOUxK2OE0KLztZ0fK9cEvUkTt+ogpAmSyn0/xb4dWHuRI12Uy
lL5D5J9RPB7XvFlTWzq/LU85CvownD8wD160e8x2/xp4fvgXyDTNJ6LnReEb
e4kTKyWHV5BNOXJkN+tpqKHLZT9s71Yfq99uJjfgWNX0mFohKQ2yP0lDB5su
0TTwpqOL/jLnOegm9ktlrSoh756BCy4QdE40YSnM+dYR/pwtcAjeRs5d8+Yp
9PoBINNIP57MlRZN59VGhDMep3uAcFVczYh5oqXwhg52nXiZ0MpuJ98VVQAs
mLFfYv5aaNwz0D9AdNavPXjj+PZSwbytmO8ZZ8CXS9RWdFFY+M2z0FCqbbo4
hLEKbjN1hu+BrWkih3OLLYf63PU7xoyBmw2w/XkAKTwhzN42fuBsm0DNed45
HkzSV6HAkOTVR1oeW23G0nNluYssy3XfdEM69TTKareLRWDuOpsbiYCN3Mv2
bi5+DNuDg7NDQxCJ1Z8kHcJpq3GmVYhwK5HByRbMt3yKtpvPA2BhLHhIq5mt
K4D6bLr8scpyqp6faPqfr9cDZe9kcP33hbvpns/bUmmW3qyCTy78v2KpjPNl
akJY62EZSj1NXxqUyf6+tyRgOfKVzHfbMmbDPL/Xb0nd12HSc239tMBoGU6z
7LfvlzJ9tZMS+FkmQOimWR2+k1HS16FwHkSlorLPaWG8kDEJo1QwfB4Yc6hy
/YXI9daqgyLsVOOT9aU5dSLSh9P3ipMFMox4B3BT3oVawWkpsDQF0RjtRhnS
VQ2zIR5d99Jsn2/uCpELaXeJMPfNgo/e6vptT13I0uZIHsYgL3+GIt3cmtei
GOj+EdKxcmcgfRYleFe8E4j18du1QWe8TsHIyhR29yJHnMHgUmb+NaHY/lR/
VTbxVCLuHoxmFSMg0Whrckygr2PMMYMTGa42rQbb6gTuGgVhHIMP2knqtQRg
k0yVdZedOQWKtkHP1Pg0tlU3u3qHzHOQVF0MMQhirS3QZoVLAB/iybXVheiI
BnJCuSkybkZ/4IyITxsOVEYluV6H5KkjUQxRDdwjwcwiFz5ZC/HKieFHgXF5
V5DgfEvvO1vCd4QEz0iGyYz+C2Jl7xjl4TeOsBzNYLZ723T1Ng4+eUYJICTI
og6fpP7JoN1ioNU9vD+9LxaHL9Iet4iCtwl2ZwC0LLsJBMjqh9EJEKZKTNtb
LpehvBdHsgcoeTBiHudduRkNhltdTbFEdDQ4QVMLA15FGEYxveNG8eBLmS45
MeZZzL/wC3kztNWxgx/r4YkSQa2ElCUcWy+bjn8g2BIhILvn2dtBDFoLTof6
X8BlZUkN079NiOpB97JKtqhsAjIBb63mSZpdbZm4FpWry2Cqt9uz4bpsCrv0
UGIZfu/v1zvHK3WtP5t627zVkR7LpqRG2+3JSLAIhM/ZCtoXuKGID61isd/A
I0qMa0ij+XDQUeBaTSJVW8FFFzZX6afDRQ/06E0K3OjfPgZwDL/NBRE+mN4J
Uk+IXhWWvA7S82BHSP76euaulKXh9oVSJvAllLrGhKiWyB6Ww+2GAG3VG8zw
8aB+ymP2FdWUWm8sZbBqeL5OAcUAp66au3Ph4mPl1OOkA3o+ypmak2KMoxks
iF46RM6vDG+rbVhjKkz9pg7ZwtYyGlTOnsU9/3EuBMt3ZM7jFZ1V3jHmzuwx
9TutLrwOyK3bAZ8qtQCEPCssOCb5q4mH93vBqydBhUlKy/hvKPh61XbzPv5W
+s3pWNtf22kqqr1mlKQ4ocha49xdKnFiqjVEz4D/aNtsC0EcwzEEwZju+tIO
vu7E1bRZs5ppbrKTQ6C194YXvHHk5s1lhf7+0gO3QBJtYrfzZJOT/TYt99Nk
B5m6WDq/AA2v0YlNhdsVc7FIC3Fg/9CSXROeuieQYuqTa40KE7BRIvvPTfqK
xh1m1+qKygk7oNTnrBn+/9AwHSCxteRIXbaQYnJfa36u8+UidFGILyofjS7f
DowekUm7JzXIr9px3Zoa1HY4M5gyqFaHDY1KeWdBrj2NULdTYVqNTfngOQDS
Vtf8nOQEgsQzuCJPLwGTQlWv+FHjxaZkBHNghf7EjU6mBlFNcIFroi8J3AIY
VyxbogrcBipktGjH934Lp29y2tczi4j4XKF6dqv40jc5nyQv83/gphMqf1cn
J5co2v0qRN0OpzmEQGPjGVNmzmyOkECjlCAMM5UK9bdzMHXqS3BKydPLummx
Bc7EKztu0Qf2i/cW/PSc0PvQNtaZXWQxujzYI3UB1QF7+udIRBhhdj2VOQ6G
SwGjwQirOzrGuOcHRFmEYeZ5RjbgDlsEoDXa+0d9q9DKC/0BuEbkZa2ZNuS0
5POtmv4HM/Pl8P0I4uC7xQCdFqAinPgKGLrNQ5KZFEMFCuSzVM2MuBm77eJD
oqNfZnI1ZkBPX/7o5GjrQxa8VL7ZXsCA7McKwaigmyZ2dsJD8ur+mRnsMN8C
cAxG7G2JbGsDg557NCG/IfMxoHG0I9sn5rldNNUb01tuSvLXxmfUaf8ePTb3
0UOn8CfnBcrN7xz/RYRj8uYVtwFargHZS2+2OtYoRkzEZeTfQ8DB0wM4Po3k
k/xs4vL/fzZlwILEwtQzXN/HMnBtU+uMPw5kcOBp0ICr5seAxMrx35zndpGK
tEwhWLO6bGy2C7E6JLr2RfEN6ePGrIvFirxVXgjsHiW3lQ7WUsdXVyRIMKG6
2VoUalozHFIKyvEWDdlY5EmPH0FKMxMmcc/gUVyk5McoKwzSA3hwPYm8aTN8
15iyuBPihIpwRUtUJICykM9xFsuSZURb/IQf+PZ+MoDFaZzdm3iw7kgiOPZ1
BcmfD4nWrUdJQGkStk1XlUTrNuJw0JyqRfBFwMzYEE8Nuo08gilk+4K4AxqZ
F6NEGQtVK6SRJLf1X5rZ9cXc0HUjMY8/uSkn7Pm/i3LZovfjq+LXzMzYLST0
TFtaop/9w96vzuGYVYsyseV6jMJEIsWuLdCsazSc2FPUdO6cipH939/kKnXw
xOJGbeYzjRzUVbIGkoTr++y8wUw2xwhTYkuZlkVM2kWhS1+gwQvSBvx+hWY0
o29EOvRez6cJUqf+/L4JfEUdBoiPndBcrc+emXJBJPTNGF5keYOY0ctmaTHs
eLQJLBaLbmOkl8bwt/EGelJ3WXRGA2QQiMy0OiOsMy/EJYZ6xbRD4ie81hWJ
oAraGCKDmwchdtCaQIidgHGgHRGq/jG71ElmwfWq2BaxQHEkR5l29LlfCloz
wNKxj5pPsAB+KTM5ZAIVqrVKU+pbTYHAIgUnzg+KyiCNASjAY9OzArwllD5r
iMCIZkjdu08Xz4Y2ESyWru28Y4M4GaydrIYdqQvpU0y9kvXlldBJMEu2p/A7
scUdk1leRrysTjCKdt0Ax/QQ6/aoN4wZkD0kh/p7ngnIwSaful7RnH5eSCM/
JQLCebjLvih5nL9ssusbEShAoibfucW5RK9D6db+q2Y9qOqwUIdGZ+L/2+KM
wBVKIrIAmeEtxIUM95b58KQobunEaJJ0bTisP0Ac1dJ1w8mxjY6LMgPkfSYx
RrP8NiL7mKvyHXIo9ogkTExiioef/3w7UNlPO9XEQtrTMLseBGg1LWYDBPTI
WxY/wIUNJcekyndPsc8VFr8G/WHmKJdxL8JDAU2wL1w0mkDvxyQko5HHLBE+
3lN7LA6JTFzZVw+JRt7GTPx2LXLZCs2d/+3RoxR7stqIbLAb5umeVqyAF/dx
SmulQsbXgJP6rgZ5K1GM15ZXRXgZKYGKlFuWAHeekqcjhzF36dgDp6YYOUWC
ezJM3G8nnY81eAlMwkInF+hjfs8jFCvD16l1jVIamI2rqaBbpCSqkkaAiqL4
AF41GrRLozT6obBb2F7eUv3K00xsboHIwIhk10kp5Dvt8PvZ7MkyUuvdg4n2
gjBR3wcflnxPlbGPTms9HS8zxpNkfdH2037qlIK/EHxSRvR4njOIsPQxd8EY
KafrZblxkSWBIjbcRknbJyQNHP44OZqMxkHPJiRkWY5uHBmr1VwUviM5D8Vo
awwCWyCJqeIKaR6b9dZ+jIUDiyTPM470ZPI+rJzb3rPcKGl+S3T5C2xrGXet
MrZxhUGpSjhbflMSfwXtN5/itxZR9K85Kc3n+SR6k66f+lrAEGmK+suMNFfh
6itiUHpHyGYpKAtCl73J8fUi/K0SKxhWIKtJqJA1crR/nV+yUJpqYK9bf0jY
JtSBiAjxQyVyR/VBshwDxeJ0wKj9hFpdbzC//NZ74rmShcBQwjqE+zhO2HJ1
rO12fnqB13eyQg5H5AQcsq7d5E3q6wtJsTkR31P/cBVQN/Yr9rXinFhyPuGO
nx6Yo6gg5iyYm09I/zanK8TmH3w6Jplla0e0AzVgazImUY7kwB4QK8npHoWe
+lB64eB4L9eV7i59ARpXsqboehspwsF6VLYF0ivSTyhsFZubyZLc/BWCqwT0
5PlF4WvY2pw/2sUUqTeOFkc4oqo99XJ4I4KZm6AmfgkGZvAWFlGu0PVdf8Pn
PnQyRUWSYtGy8zAb4JDR9MFZ89Lg5OY+Ap2GbJl2hM+RN8kDSs8k5KS/SQj4
rINKLuJyJMmnEURysAV7SFzEOEQfllzUR6yxf2oce5qcr8dNmRNRf6TRd+zo
Oa+M4vy/XTYbXAVux+5FJ2HMR988XMPdyrFTeO1I7LgOaBAmaHCKt5GUmcny
JdL1fCtgPr5xHlpk4VN+DG1u0pJsHmzmBhdGiNwmgUcyYxudkzmX/3f/5xNb
MPL4uHjbZtKmgfsD8ihrI02ezEek0zl/nWLCY1skn9QRNgljVF2wGT6zcDkY
fzi4c/Q9EfF+NcGAi+GllXsIYTJW6VHvLUp8jZ86AYMDiE/dblmtfgj00zEV
NGJKrZni1aaoAzWJJ3ZrL2aQbmqgdS6ywATgLxhrgftFaXvQGJD31HqbDyLH
29Bc7Mz2mqKHhkra4owlLkkDgbQAGBeZECwsogXwBlieRKcJa6VFQpS9zB7w
nhxUI5Yxi+yoSasGqr0wUiKJkM5rA4OMyRrSsaSZnQxwxH+k2lIMkh2eT+OO
YQahHnWsY+6hrJqJuMtGu+9osE9Lq6Lf1On4FueJmhrnLyOgbXG3Qo2cftI5
Kvg77y/7T8bgnCOaXwiyS2Yfo0p0t2BpVagZ7LBViozgKGAoaOrGLzph++VO
Ybvz0Psrk+SuJQ7FcGgJ5I99/bqj6d/cr6QesXce0m+yICdnBoXF8gv8lODZ
autzSDGVgbnvoY5zX022BhI0rXwfcsKwNyQdZWj+8WKhXSn5Mg7uJvP8EwWg
vunWCnWbwqOuhXT0t0vcsdPd2lthetCNpBaUyVC7bs0XaIMcOirH0re6ZBE2
Pzt6dJOJw5nhgTPoN+/gQTl7ZqWPzl2ZFCR2tlC0Hcc5Yi61U5IfrOh9O7A9
ekAZRCozuCO+xEYKyPQlTIMmUDxqmpOh7zSToLP4SZTfqIdyES4uUlKcE6ZT
ljnKYFiHU4qDWyJO0mBUm77xaOJzaUYufzBMCSkMiTaNWJ6N66oJD1/ZfjGb
aG3en/BMQVTw7MtSWbu0GlO0OGJ13pUZ21lehqHrofo+3e9yuwo5CEcPzfoN
WEr0OqrM4g6cq0Fx3sdi6cHVip9eEACWZ8U8fHxgsqCm7tgnVPLq6l7XLqV1
yAsAz02+vvfb4eulFrz47h3zKkV4PpoCr+FUX5LgVV331ZJo41dfvVQ49EQO
AcUDrX9FJmcoR3xwXd7cr87vfkJeYZHUiV+SEv8t5ejUZhFepO+cOiOsUxbb
sw3DtTRv8ZLOXkd/xW3FAZiWVAqjOpn81qAC1OduEp9FQlXu1Fqv+uCwHiG6
5+njEu7AcjCjLKk0Qc8Fttev+NVL65293e6yAaRrtYzQnODodxaa/xq1yUax
LwPVF9Flk6gdvxKUgMqxSempAk+zR5rsXboZF3K7eUC/iqYdhW6uLdbZJ7YG
UgGAGuQtWW467ACrKq6+Xf7STJ8+wa+IuwYQC6EYtqzfUw/LkrlfUIG/K80f
h45iRwEwCCXJORpppcwTaG0RR83pCbJLK8L0EyWLSBbCMrM9YaO24lPWR8UH
x2WMvMLKoyOv3HuUp/ALXZ1Xe1SELGiTXCpB6m1lRKVNDHVvV8QsHsWEbdgj
3BjsiwJdn3WD+3y2AAE0UNI00QhTt/M8L7R3m09Qx3QSkrKvfqZimBOfDNYu
9joOSlPtXxVEIsPo7S4hE7Tc71qVJ6MGMIcu62xLdkGsEn5AvLXvJ96ggeRw
k2WDIU7Sl2LiMABYlKABtdndnwWbPkS6iBVqQagoMtLluZsLDOoCbGUYDxQ2
A414sA1tI/slEMOp9eQs+ACUq0ute0O6l7ndroMQ+cTOfNa6X9iE+yrBLXHS
Wt7/jOPFuD4VN7+eggV0H546bgxKLjMvf6976up6UX6J+rMLjdNqrv7AzRRE
PrJ7LOrf5Bcqi32Na5SCpFemtbOQTz2iMhR3bb22dcolmn+NAIlh03PdVhXd
zAa98GSsAOUpsjH2hYdQsidAtNRjqG71OhF4D9YfIyaamAujMNjEdXhJO+nj
y9C/m9xyrF4UQuBkEkVdh5uaPVwYPXZniaG6zrwxNWHSc72TQlCewOBKLMnx
jrH9f+3Iwvu6btbrV43dYP9ZI1Bdhyf4pBEfaRnUwpfazC4eOrl1FkHOh60b
szHEivumT2YxtJHTxV6+pbVjK5QG7RsXCsXC0PiQCmJ4STxuZcWxtHoNvHcO
hQxnJ657RecAZLlbV8y6qWeMQ/7kK8boUDrg8XbOWywt5OVxs/5I+HLTZj7E
3hlydx6G3igenNs0JgM1ovRjhE3bzfqL5zawj4QkZxTJo/ZWspAJBLzxGa9R
Cn/c1WciWKA37P93ngcPwJurgSsj4BwwD3TwTHBQTgeuYEK2je4wz623Ei9U
eAoRLEY6CZDp88ZkrhMMbu54uvPgviRg7AO8eWn51p9c5HIYpU3iuX1M0EyN
HQBYVXBUiZTOna4PrG6qdui4OyrQnTfcZ/9+1Ct6BIf0jIyBg1XRq1Iiw7uR
6BnauQwLCo7GNFAWbTvfICNPE0jRTXaCHLav1PYe71s2yzOH0GtB4dZKoU5f
o29m6jBOKifTtQtgGi/rRybBkPiga4PAoGUvjUvJEDhdFhN1hdyrV+Ewf8Jn
k78iI+52ovMhOylwoasShQE8lepm7ry5sDTQs8xyeCT6ovAVhbD3DaHQgO0i
rJWcCFa/UeN8mwDb1+X0Jx9BcfnYY7+UOaG+It/tDzxn+TX7qHefOj4gtEuI
Fe9SKGDiDoV2k2omKIi+19kHeLQldOFql9fOwE5YdlPIRGVUqa2oPxGeoLEX
V88QuqnXW4KbnLLNed4v8ckzEHJD2gssjz+XsDduPOcjeZa+mTfww5P9b/mo
WLBnr0gFMbf2JWPa+7+0OI11tUDp14Z8tVwz81vL9zBG7dfz7wzcpcoDidNv
zWIpXQPKzTEnwZKxTVPrdTI8GmO3RVeO9uVJD1e8P0y5KjUM0k4uddgRdUfM
XBhDsj/Heb1Nt+pTWXecYbb5WzX5aG0AOfP9LnIicA++wb3ugJPnQHYhtsjh
NDzr/ZWHbOUiKFH6c34PXg3nDWAiYhQ2C07j/ui/qVePYe4IvvRiDjH5R/cN
C8uGXuPODfDwdPqFKwgl4urbQC6qn8PLqlF4TFlYz9EZphvmhdXoriyaYSV2
yaLOaY6SrxPFdAhyDS/ZP8pVKkA3A3D2uQYY4+6jBueoah72bBxDtQHxAix9
ZkgotOKkjVE5/MWyhhBq3O2KjjQtBGkhBF1kfHt2No4Qsn17JJeTXuIWD8lj
7qkj7oBEr+lUreqL/8taIpchyUanFjiaTyl5MpDm4iJT9c3F7rNnjnCGdVYM
2heDvJW6SCHANuXFRm9NtJG0y8FxN5rWHlibcdn4hazISJn7p83HDfYJfbqY
SApG/Oz5eDec7MdfQ2XcBkqaYG7oIYlBr7E4geGEvtfPzxgFOiKVKL9iahDI
Op4rXaymr300esincoGpRTTuAiUtl7cZyhEiHzarv1oszMj6iiRGcxYTZWH/
dADl10OSJrXb8GilXvkX5wlxYLmxzUyZlGubbe81pffzQD3d7muFbrdg4kRP
g6H7t2bg9tsH8h9SPZfII3J9xtPATkDGrM0O2zSsuw6rCKYpr3W/uA0RqGCy
pxzTXiSR3smaOQJMcAYXKPg6L6N/g4VjltatA/6/fyRR0Eosipw/DWMSc4VO
d2I7rthB+CTjoU6JlyvwS5sfHZfNmRclmwpUZVLfZDNgXxXVbs3RJK2V2DRE
xVHrUAOK10KLZyjZ3gAedSym95u49jSFpy/tZlXjeblWPIWa+UDMKkFmtENB
Z8gWyvd8FxidY31luWNq0tGkJw73ZWXzuusVT2MiXqn/kx1ZHyGWxEycZO3u
OTxktQLkLac+Jj3BqRJgiH/EndD06Krgugp3D+1foEanWMBHGVivi8MlS5yT
l9PJyCVr9dZpSTiz51+MTP9rsgpKW5mjvo64/S329OEaOlMJmbLfNRy47LPV
MQfTXgOPSZiouGRz/vXsDiuJNlfSowhhiEcXGuU7cui3u6cmxaUUr498Wad8
TX0fwCt+oyxEP/IqCX3tHldu+9eg0+GBnLnJcyyUzBj5osMGmKiqaQs8ymIA
tTz2smw09tnrXoGwnYPtb+ht0aHRf4T54K0MvUpifIrXjW8taB6r7ExmoIMi
HhNG3n89B5FBNQvfLFcT6Su7pWIyPV0a5G9xlnVD2bvm9/fwY4nuhINn5QrO
r7MRJharFK4JF1u2DWimKJx7DNMpOMoRuksrp/ZaMJmF57FTU2/4b2LnQlZk
XQ7l8d1Qz+pNb2cNGklas1B/GGozbI3z5Z8uVTVe/QP4W29SsZuNrazSYYfO
+WLVpferMFRDui5vjIxescMIAP5Dfj0lIK50xwIIZT9jHnmHegJMGICr+eB8
s3lv/Rq47kuStPzBzrDxUE4QmFsKl/9c7PJ2SOLz1BnvOlpXfXBUxnD+RFje
pP1gksP317GGlyg5bB/8WINycNug/fhN4OUSGTb7zXvLGYCxLY7PDaTt3ydo
XZVlbrTH9kfLkPhpV7Vfor95MGK/x4Wgz0uXfT/qloK2K+RwJF8C5KSkRF5q
yn9snXI5YvXBmjEe0xgRMNyYMYbLrxyo1xPg/3FdIuEabeSA9VMig48bnSCe
ljXnjxjV2dIZuF5Mc744gEau74ujrvUGsO2+yaykXHxC/rX4hVBo2tZUMioH
9G3EeSY8YLWRyfZKIdpexOSrjYwlGZrVW5ep2ntcfhGJtx5cFS/PJwfh9U0k
h4vYSRErt0gDHM+Zo9tBgzT2dKHgKSh7JildssMGH+Y5l8MEai9hQwXthp0N
djwNZQbTE+J0EQtb3gtTrIeSO/WO4XfAt3mZSoJxazElZ4BHhHp5qYZHEHFk
+cKpnmy2qR0qe8Wk3xXqxhZAzxXuI/KIJFjf979vczRP8K9Rx8aclrg5DaMw
UbZWon31oh8B2lAnrYfPr40uZ8NC14vpT1dV6SEAReRQ3nADmPTq2TZiUi3E
qHU8fvO8j+lnP3jZZz0pabJuF2FJw3qREG3MQXDyHe7lGY2xMTzM+QFyvA5f
0IIg0J+gk1MZDmVqVmPufv+LkfwInaAkTst9XwPsPej0Rr5DU8JHdF0Jx1MF
G+ic1U+xR7Qfh9jbqLN2tGacjbxkhjIqgdTuFY7n4T20uEh4lxMoiY+mAhfT
DyPNfaiKe3ROSE+uFXl1uyUgpOBd1w7DdQefBiASVbXU/O/A3NksrWYU7Qxz
+ffR3T1T1Dmm541o4lCKB38mvaOg8VHietPwW0kkbG/E5mbhIx7+Zc8Ou6B7
LXYZFF25Q5TKzmDR7lHQO70sCPOZ3zL45Q5VjJLqBNuZGo1rI23B3wSwkrwZ
P5Pe1dGq5cA24OPGiX3BC6GU9Mg1crdgvd+Q4rmXyBpPBUiiv/OhGKW8Tiw6
IA/mLJkWN9Kkh6BRfLU3e634utftqr5qqlpkAsGh6ClNS1q5cidDmHp2gz03
YTFdJDRBnBKd5i2btJzMgquUXXGveALMCa93H/x9SR0JaqThizKRsWOSrtqw
D/Qnqzvrx90hVqazjCGuVcefkJxwZPS8HkTPWELFICecwUdmS0Lo6krRu/Dl
hKjAs9+9Nni5zyRfvfupNooeWlvpHo/6FSmvYdg1Vc9tLIYBl3oVZas9dH6V
TUiZXveyO8g7KMfPHGBkDynrrrGdUabfuKss/lHBUO61ebtn8eeUCX2I1tlr
Y26qhiETR0bLu7mKa2Bd06XJtkAhRqnqOHFGiYdTI2IexFuc4tlZL/j0shf8
RIQKODKVhNUm4JB7gEzNr7F5cFiP369NI7BbMV52OJ1dgXZL9BsXnds8vNVg
fRkuDkLsl+V8iqhXsSsSB1qGnObcBei4yh8YrheXQOmNBW01OIuHS5vivIK7
7GACoDZqr0nrb7k1kv6rxdmJpqUhvGbc4mlGGrer8uuv8KxtTSIpkYbcFUN2
dj7MYaIY0W8eLuTg6Ag0UG91ZdpiXSaB5Jk8OOuc4x3lweeRiOkTPm+5kaYV
Q4izndRFUbdYRPac2bMnR1qXdoU+kD7DKIBRNxjlpr5Hzn+arXpbnuWcKW/G
mTNFgz2JbpCz5q893gN4exk4oXeIK9GUiFCxDGt9uFXt/HmVSLLQrGE2gy2g
45HePahNEHRvA1LLWKhrrLuf3zNz61fzKhGm7sKwMvargXklF4a9iYhkfS1M
UoKxL0mVEicM4uO2RksuhZqovLFqAeA6YJK+Hb68s+/g7MHDYBvQjiCmxVAW
f1j2CreodHFJH1ZYr5+QxsQzehhQwCc7TljhTCWYpAawuC4zMKMgwIYTjkIT
ycneL7Bf79y/yPEBMJBExPNcqOV5NTp6zAfQKNL0SlBi1WZ7lmmwMcwa1x3y
1aP2z76x4u/b0f9xfkqdOaGhKu0yfUCq0rRBhD118JKMW+1azoINs3tfZPYV
tHYHv4+f+QySCDQ5QJP58n6n8iTaVxAEjhCs6YgZNjS30na0l97Scpd9VlsF
ogoGxJxZl/R16BRB1RaXzt+GWyGaxlakHkCDv72cSi7l3+u0pi6zQ9gATwbP
HEC13RAbTnxFYqbdgKhDAzeWzfv+e9OGX5W2bMUWJx/N+hFpdYeceIBAr5II
CvgASEePX5qslkr7hjASMTVc3l4UkVW7nvDKKAbs9wpzXg5pOcZM81EvTW8+
kJhoEt2uumLgogwfUAszxU3dOE3R5gvZ2XFajSi51mk8fNK+IZGhYczmaGE4
guhCPNwwkShUab9Et+ukaSLhlAN6lQ6QmEk0Rwc0BZs3tIkCxwW6W8yHYQYm
JphnyyTfkxo3Uw8iK+XTNCmOroojPEHXQehVXjyZFJkxjZKhbiwZkR/jR8ot
YZ8K+xPcDBzISfp/w4lBQ/FOoH2hbdFj7VBr8KPaZELnybyMyAqgEVmrLCTJ
/2Ngzy4ctGeDNVOZFRChBpaJJSd7JxpOPvhJje0UXJEPjBrrZlRK//4oWI4f
TCzDb4zXzzAq3FN2+vljZ5QKLTN8Bs5Lrj+ipNOF1rhY+O2lpT1wARtaDbMC
uGJhMMMyyui5JbFo0It+mKB0L3Do2NH6MgqX/KJiH1DN39y9W7+kL4fAdhY0
of6ejY87yAQNh9e5EeUQH/rfjDgbon93vtYWMGSklRHYfk0D0Zv1L9P8Vuy1
tUOMiMOqWwfYxDTVMZoX3COXdOfY4HJCwaL4iGgNxRb0DDV8u7TvRWRPCrCW
IkbsE+bTP8UuZMvYTmfn3FAfHLZOocXVRWfmn5LTMHNa9CSAUQLtj6AYL8lk
rFZEA3oycCejtJBG47vZMg/YAV4Jd8JCUlaBKUiHi/Kd4U4E97uVxkzf4IVt
/r3qHUzHp1blJbGceSv+vOKx9iJ4OBLRPGGp+2e3CBnmib3rJQKwgcIkeXb9
snNw+152rWjQfF9gTUp5bVZ2np9C8LKrGtgJicq8qQ3Abo1ELe/rAlHg6+Zv
rkVUEgLRYY0lworIBsumFToy1i/lvCIJgtH/OpoXTqZWv3LztVsWCfSIruVK
N0f//byNVcjOleooiSgqtOlRyBiVaGaKp1KNFR/X56EdJPfAKakGEfUhZm9J
NLV9N+48sx3RFCviaexfUemAtbmBneADGUL9V4EsDF/k3LQSbdILJ9h/VOIc
67JzeHF4t6yr/TuHOgY+ZhWMb3mzloecI8epeJhWzE/U4+wsICOrAyjz4KLs
PYkrcLuVHLRGR1rTs+WxUOi8W6tSwwU166T11zkJEdlZ9cBtQ6dHSt1VoLgY
gxF0AyAbaLfHXEifBUnpHn+v8pUwnV6RfLgTXRtbbvUzkdmFXsZBtv0CWehI
RB/Jg1a+FoItf7X6AonLYSM3OJCTVDsc1c4zezto7OHk3Y1q6r2X6ufWcXIV
tBYnljsMnXJE9ZAmQOVYA4Qfmnb94spk3l6KrGwfpaerXg1mRYgAu3ozc4+c
E3S6dX3jr5Hg9uI+wcD93oPMEhLgeqHlWD5IwnCcXaJu6ahrZVNxVhnsnCKr
hFrc08FYFKZLFmqp+99cPooYIDUj1UsYAs1SCcTMm/IM3eW2o1c00AToSYRs
xUdJ33jTK7iMveqSNpa6mTgTIvCDRVGAz1qeWP83nFzOAJY6vPER0b3fcbTG
Z1qjN63aaPwbkpbpF0Ia13MVwbKx/J+L26x0ifSmF7CZVsRyLaK66UybMn0z
IJmEWV5YeW0bpju+gEp4JsUs2UwYxIZN28U+uauV5Rn1Nz2deo/BAoU7anji
20r8pk8Al3aYgAh3Y504Moy4rq4Dh7knLckun4zh1/onFiuHe69LfnlCEm2U
zGfU43tr78hPhAzwtcN/e91Zp8K2YfCRw3QKeiipsPGWjsTo/Dh/6vDrRWr8
Ds1rZc9MvUSof2Mx6O8cr2B4KTSfXjYhA8iadpMheUkQvnlIHKP0CT1nuEWN
oZYQY0Ds0hRdr7orLNqzWITB+AG/Qbj7Y3j5smQOeFXyzc+BtPOiODn8X8CX
r1gjoeu1PUK3H+6UkzF44wDK3j8NP4vdBl9pV6mf/C1GA8WLLi6oVVybyEZ9
zPgK0LrdDQeJBHh8/DsOsINO4/gcc2VAY/fQoVhCT/Uahovmf1vCuH18DhgI
QMi8CwQ30E6jlKl7BJFuEuUZZFHHp2mLSPOk2IRLm/nFG6yfghhotjAp8upK
n2FxNQ+XdjHPWTgSPveL0x83GKuqaL0T2Q581N4cnpODLyX8FQ2yS7gHw8LK
hbue8gUTPP0fVbhcazGtVCMITGibXMkjF8AocJouQv8bdtCkmKNy0mDYlzsU
ChDNNhkU5AyzdCEBUpYd+8MfwXOtlQK/SaAklWugJkhEmBQ/9oqWtwBzyPaH
YWAXbW/Wbfp66nrtuCVc5IJj74skADl4JiHeSzYFsqGEEG/m1fQipH+Cjpp2
2b69F+qWixE5/ixmVz0g916jI/C+o+ZU/iYG0Ji0ZBXGRAtB4677ozNh2hiC
zUJNoMuUcgpcBnQTS0HfJpWJNIdunkfW1VbyUWUcGceCQuu2FkS8MKONYZFH
AFA6XmXMdEOp4fNZFTeq7lZmucUCSjGTzQkxjnGSU7JDpcHLN7kd443EY69G
bqOzQyah5FfhUIOFNx3S4HRbN0uRvugTWokZgTd8qKkMkdDSGSMGHzYxFAaN
aBAntdZWtZKx66EBRuU9vALl1aE5hJscIOIYiXUEYT0ntaeTVhBZq7vSSr9a
ocUJ9RjzXxzn1D504SRlR5p1qGxtkOkZQ8QZ/4KXNxdyaS3JEW3AjSHlmCCo
wl6/PUqVoVgZUdD8FFgjqwzd9ZkdJ8H/LDQciwef/st0Br96D/XzazirhDgc
B2avH0F8zXNKogQl+fsqk2nFRXSShwUW9u40wLzt//NL6FJNkLoA8OE8pTHp
oyMUmX6p/7q1QqD0h1BzphLz9gu6fxp7xlhRG5sBMYz879FE4Qb0OdnuuOrW
/RAyk+5kRVLCEOxeCXtOks6dXJncAvstB/QU+LQyETmkDOagocuJWpUDkmmi
fJRp9y/0reT1kmJ8LxBpTWsUpy7cZ+yv9SGXfhkLHFrSInSRmDh+0bSVJv/Q
RQ2Qd5DBWXYlD70l3QaZZCWBt/0KnsGaDWgq2Dyo1Wu94tx5ms3SVo8r5++t
5i05OO+PNsj+VXuC2BC7eJwGGKqzilcf50OZviSiwnur1L3PQr0fo3XF2b0J
l6TY0OFxKD7Sw7yvNaZNcXGI8aPBF0/mwH6xoO8vxyeYajYQPLLBIl87yPuj
Dwp+2kai6kKSpMTsjlMdL/uLRCDrdX9vc6lFHno9quIxDoKDcnP4zeKKrRxX
ulpAFESkBu6WefnpB2R6jsHJFjYpewaDrxdA8dRIw0lrdYrAuEqAZ9b6xvb4
ULUkZQ0LEb6ZY+9pi/5No/QRI8xylflHCa6kLJaHU+7yrzCRQ/HKfY/0t37h
tiW+i3DVhXCLlecTW0Hm5BSFhYvotPwUCE5fDC9zn/SKwtqxWNftdCgUCXjP
Zkfei8GnCobCzoKXqS5qKMF3g1XN64OIIP4KkvOQwmO227oHlnKI01URd8fY
Rag7g3odR1NMvGwtjpyMzvMklcYZtEJKnU2xes6X343HuJRY5ZaIcWFi6udc
BOlfzmLlvnH44XJYseOMo1F28xWNrmZx7xr2Gw/2mCtaN+9cYBJM3FM3GHkB
AiNlRbaMvOuYpF25N7TWfqRNbS/RESakvyimtQ4vCEBq9ajBooq5Ze2ZSoAs
WqrkvMH3pSsoGR1xek32cnbU7MAPcmU/1hj4gAC3rZhFA/hF5wKZPJoZkjDf
naJo6TORZv6PKRCmUFKaFOx6+OkfsDeq/fwLTChZjdH3SUgAqhkvix11qDHk
nw4ldN0EkXdn4MOoYOH0AAaPFXhiXyG5dn+qjeV/+6jEozRKtJLjWkXlOsuA
unmGrgk+J+FyWmmNCVWRM17OXy6glK48JRoeaFqe/Pg+KwYjENg5sVQuGHbJ
RZdsQ2N+r4fi+NmNK9Riw7peoNsViPE8atVfYefhaYLp4BuNbD/pWjtVn3Uy
sxP23ke16VyRM8VOWGXuCRLIaJbBH1JZ5cGRdC50etalbtsS0Wzv+nKhl8vm
f61z9E6KQFRj5KTGogJrN3Q3DWYgo0qULwV2+QJBD+TMIevAHuc9tVc2HUCH
2f77LIEoTYkKkJAuD+ZnFfraJt8hmosBIVYM8+hk8EexhDh5TLc/q/jliB47
pA4eUtE9Jb6ZCdXvHDUVsU7Ni4rnbYlXh7og5h6jFuQ6JtrwLzrKkXwos52k
jbeATeLeJtmwjNypVWosjX13PDtn91JnN+uDQH1zUgXVzaBbKp709c2FALht
11kwtdIx3w9BzST23+Un9cQ2pWqgR73xbx6icw4Y88YIGLQXWdJWnEQLu7Kl
/2Q38ePK/IbOMIdfRJQBpZC2nMM+qAyjnSdLGmG/pK0gg6xZ/MxrYw8qehYk
b2m+BuXPhDAqXGkISy8ITrHDlgLdGLAQgNOOIOvwpnKFfx4Yr+6abx67GWPr
wtoNFUTG9YJsU5Lm+J/uwWYqnMdbynGIA+AZ9HA5EflZJm8+cIJjh4zOCHF1
zBzAL8WtuAYNHVd4NPNE3bhSvSCyznFZW+Mf/kpSYGUgQ2cKq63hNqOTu+et
HTT/luIyOKO/lTF4JtPG3AtToM1ch37WuUBW8oizSP//X6/s49p1xLASCe+J
bZpbsRDx9hF9Jk4MB36oIlRe8quLLAqtdLn6phmsF6ZWUiEbc8BDFZDZ+09G
bXMfq0hUD9ZGxoGlhWHExeQH0kYssNYj1yRbjahn8hJGWRfH0a9XVJHFoUXZ
/bN7dOhGTgvgaC4VzcJ+egclMVmWFpGTX4ubmO7E83k9Fa0cmrUXSC9wgE+f
qVM1U9xf6IYECDsFU5HysP23deDZq6hUsJC78geKjx7KYLzNFS9g2ZcQgRux
ctX1IcOQcYUU/GE24zpexVynElQPMvVA9fD73uDXnBA3Fy2BF/HN/Tp/+lQu
FDupo/dF/+0upoMgCKDR1UuKH+fCPwSrKsyqnDqbZ36tpyMQYZYEW4LieQVY
GPTGuZ6S2m/HnVbNEQb6ey+4tdzSK6ZL/mUxlUpnbBT2GUuDSMVfxHUnJ2iy
3PKxhG1oXpIjwKlMpOLCprgoozh28SEYow4Z+0ZACvdFR9kGk9p7Rc5muzqw
4JdRiIgETSzqR3/bKzamvx3alWN4xPcOA9ylOnVsM3hukQB+PVf6uw6LWkUZ
leR9Otpx+NoeciuwnNtoBwsdr81ZMyGxaXQB7d3kUi1Cgku/ewTLGeBqolsy
mSaMqNAv4BaUUIR1yjxICUOoZFlh5LF6yO8T7cE/GR3uHabu1hE26REIyl6k
LigP+zrG8wtM14IYC1uABbB+xVroczb8ifqmxmWoXDOlO3VwXwCiiFiyoUFP
uSAn8QpoE80GY7fqTZ1OnaZfUYs3FOIW3kvuwI151D3QKEEI4qDG6QYp/HWd
LHGwNfeEbJPMC2PjNWU6ERbRxaltp1+agbHEkiwkqjv6Gmree6oiujLddpht
tp1UCxTXX7bU6aomR/mSnHh4yIFN29H+8EpVOG87Bz2IcNtUQ75ZUAwDf2Wi
y6MrXlPRfRtEUA4dGf3a2bmXpTMHrwzvXmel1ZpdJ5dsi8r2yf69FEXXYzzb
UqgARTaHO6jCvcNoBGr6U9P2MrCxljIyQhcZL+3vHqIvzKaxbP7cceR8wwp5
aRNNjGTKOGMSKyp42ex4QWDNxNNkJoLCE4DIDoAl71QhQQzE3hIrEqrv1MeW
O6h8qCdCJ7uShlbhIuZ7fwvyXM0OyaqT9mWJc4stjV2AomfyWBUgGf6wmAlc
lI6JKLmmtp5izJXGXw0OF5mY2TmAoaM31P9kF8Nw2NtHaSIQ/EAtDmP1gzNT
2qB5iW4sxEYCBejYZyvlsemkqhnQ4dzMdp7c0yeoodSEhQQOMO1xSA/qRwrX
Qd5Wd30gOoiF7EHXIvPC3n3KH2S0JtmsOuo+3KGkZ5A+LnWRXU+q2jL8x36L
S/fZ/0qrFKpIlTsdhgtzppC9bm04qUHObZMkZ3Wn6TatFU22pQJ4WBqG/syB
8R/4BqyrfzYsBI6fF2pzQtv2htGlZZ/ZkJDUIPVUl8lZf5CW8ABJTfwH2K+q
NkLFTbniKSUioiPJ9HjG5+vRobBHOwVPhjNKuzODgkGLax+z08Nw862jQQR9
KY8Kr0JOl3QoU97BHk3F5t4KFJoF6Eyq4kmTVFWjTvLrezQSWKMbd6y7Xwfw
mwpb4A7G3SxAUafT95oKwGCMkh2OLE6BBfsSR0nOQFhzIXYVy+I7OlYLX+RS
6yNHPFh2UytBjKZ0KEtSZkFZFsxBHedFl1AizBoklD5zSTty6DCmrcnxRWl1
o0C5axnJfBcHVSQsSEGrC+lmfKu6J4k3W9Cpzg53ZrzD4oMDftf44nWmTSZJ
h4U/ZmtsF9ca59fUdqFFwc5MpeTFSzXiKveyqGVy4vJJEBMeqB8c1FFFoLpC
LJttzQy1ea3JL6ycPDzkKu8i5XLlrd4hY8c9O8gHm/+/zM11hBLdeU3Xtto9
jS45H1ZXctU3oqFxo90HKDVVWdtKoht0ZaSWkOEOoKt0fhfS0dgHC9jHJ+A4
3czH/eQB4ILFSDgNB0CBJfnVfdmRIfRJGCpMGPqdH0bCDFBbLKxa9H5nUKpl
pktvbr/C+deExfJEKTpeYqQ+3HT8X3hZzwicp/8gLWQFztTsnksMISOqiawp
AAvMiY+u32Hc+aJD2uqXzh53DQCLxfiTaFMv0wCYrphy1iU75g0/haFV98eL
XmLalSNSp5dCfvlOPgilgcq8yBLp8VhaoBmexKnjTZMnfrozJBU6iJJ4Bmrr
Xq4hn+Ga9OzblM7qjtOMrkXkYFzx2745eQ/4HK4DJ6e+72BOMQABGQtCQ2ji
NJmFXDvemd5+EIfBywaXKaiGeNoMRzXPcZYQuGsPO65eVxFAa4RQESX8fITz
oiAmlaQSRYaTxc5mWt5Un+hcGH7AW5r/NWilTBCydCWPIZer1rxp7AKezhRM
m4ej0VsAmfp8B7bp5LVrfBn/7fcJftuknxNx9lKqFYmS7k8i0Qq1LWQJLPkr
ngPBZ4wH0GKM6/91pPA8+nbQzGdFWVf11EvalXlyNnhxpIDlzL+00XaiMwXb
eVg7a0SUBQagWSigBgQ5O/qh2eQMD0SWniKsqtOGCROCxrSnMyMdI5kBJ+7T
1k6xrm/boUXtkpqSsccCygJkGjwA7sNc7ipBIUIYDKq9jcyC/kf8kSK/MdWo
TnrmkMX0VbVA8Zw5yqrI3sa3iQ5zBsBKhtoJy/mIB4f7b9Fr1HofQ64iyd9+
lrMmj0NNanVwsO8fajEFCJlS3tMzleTfYYOCouUA2uxn+Ce4JdMc3pCyENN/
RWYmG8MI4Px3sOOYIL/U3A8LEDjFD496gh4gPdrWSt0iakZtk0KFZoGDQYax
SJTXHslpUctlDNA+xkeGfXdoZrq+K0K80XovJmKAHzIj+Zf9ckQ3QeQw4QrN
xAnx1mYA9U/DFSPGJT2lqMqqhmb1EZdnIZXRprW012pGBl1QLEHwwi44DW3w
beFCgv2/bG/KrA4/QdpG1btt4IWMZ0yC6PaU6WC70m8at1zNei/M6dq2pewg
bqNsUI3U6NPvqvP+T6eFwgxP7N220k5E4wJ1OHcG2zvtfg30a9VyahRB6Glc
7fbgN9sSknPtb9e+trXP1PoOqLXvfvwZEi1qWQJYw8kxfxtuR4Eqikoh662x
sstd2kWza/Br0R+dP2GzjSmTRz7TmbjcLqnauKGsOTgVd3dgG14FrsLppOd8
p08JyLPvMa0jGWx1bdspesNSVt1y+AZz6/zrR9JVRHBU30OgxY3jnW+KeIRe
JIBNdnP3HMTgIg/oohwE2VECkyb7+MOZkPj/8aFgiLX3jgtjZLr0FAziSpjp
UgtHrZxqg6SxKVapYluKUQui2p8f81All03ROJNu4p9dagjjRcM1flgGcXpm
DtwXWX1i+nwDteFwIQ2Y21h00OHc3CtnV9l6n9Z6LBkoSabQ3hgDirIxoZxF
OMGFpMwVc3MDg1Em9q3oFzEKapz6tds6lT4hkpkiS/qx1zTsI+vYWWTsqZ2B
YSm/UnN5bIf3s+EqI65G8UnrSmFTBHy/WJDaNbvgvGqYOsnlEHWB8mYFmKIS
4T0yYBxSdGbRvm1S78eWCLOTzddRC0ecex0k29bz7TQSJVqVgOyqOyrOzB5p
3+nQcMGmgFQOgRxOj9upAjLqBy3SOfoHIjyAYCflb5+9xyXaBBD/rUvR6zG4
BDUTDHVhptajkhUToxPBzHj1SE8HkjfGbPu+C9foWK6lEXQD5uUvows719w/
0kC4t8YqMCeoqARiiwDwe7KClSmS8gc0D30T71v9gy60f+Oyoz9fsnbtjTO+
6YaQ7F93Qn+k9LBFrWb0MeWrSHQTmwqY3yBhagx6YEy4Byq2khviWPdyrJ/1
T4p7VXPsk5LCNND9SBwZjLVaYsMjP6qdOZUiXl+GQzKcLFz+BzCYkjqQ5WtK
FmIlzZuP6fe1gOj/cYZCHCR6G0hnxSf59SrCQg96lWcfGyZXhyN6+8YYget2
/dbEeOVY9GFLGkZzPSaikgL3ECf+P3uyjNQKGcBiKcFAZPTxPcNa7jXxAdKm
CXsAntnSJJXEUhU/ZexnoeC7QZ/uACTIzGzaRiSTqmerbo9L5cSjr+fz2ex1
9ebhbh+Eg6RR3lY0jfxmuDnVsR4KThss1EFFlrL7ggHGM8UO1rIHRGkyLn80
ePZ5fcUrWRBi/5XkSWxKiRelTMWbtBCsoN2PscshC0DjA+5TO6v8SZxXEGH/
4xS7oiPr4WEKOq1LpA6Gq0f8HelzK80D/fFhCbypS8/IMqIYHtueKO+jM8Y3
LGJqWFiOy43FQBcoF9G3iduTIQvlf14Iq53zrXsihsd3CYv8Rnp80xOs8PKF
PGPDkD/w91ouQNxA+eckP5pVpHH/5yfzy4ZFxGVK1C7JIJkBgewUV29FIW/l
+L/0blI2jFXl51ygwh/q8T0zKqZ+CtFun6zwcv1mCSh9hX4gxdNVxxGPuuOL
/jyL46pzQTMn9NXGBYmrVmzIHUaX8v9R20CsI+JY7gNg+E3J13KDt/ZgZ8m2
+eJ1WqPnbZY0EOwIOPU0ZXgVgaEBaH7x2lTC3TCn/O0QsShemGsW2ssAnFc3
zwfBDnAc2y6LPOg72uyf55swvebuWzLYBaLJ4KnHV1jI0HRtkDZxiHepHgsJ
ujr0zkCRxC2aiA/sCW2vncHJYIYjz6dD7LemsYHi8l2+bdHAA8qHEpxt96gO
0nFQTzMP9LpcmBzhQKB2pfkqJruWzjCTwE1bcZZZYKFALOZHF4SpZpZDtxo5
F//LlaSwJ/2LvlgYtIxDOMyI/6pgZ1qrlRf3Egz895cNdMaepuWofNQw+wEl
JOyd1ncKBlxVC0mokS47oVk8WhiGXye48lUorcQrZGUI9+as9WYUsmcdiPr7
hwKSZh3RIEkt2yP0Gj7KZu275dpJntwAjGCpHX6TZEXEF9VANaoU5gHBgnPR
U7vbwtpeLgzvKodpj7Ni6UkBoCw/PG7c44NGWq+26Z+GIbeBFdUz0NadKot/
yFiQqyY+swV8VFpUN5132hcAQHRaH/KZJWHXmZCmSRqetzpXrnUERS6Q3tAI
v3qCjki5WY14NcS7V7vkWTycnfyeLX6SQdvCg1UYh7bFpGgRlu5IwD2IhHm+
xHebXq71+7X5q5SFfTaHcJtyOcBB9tM72GnMgftCPLQBo7FHYFYhoBZvIhKz
RWsKcfjvZnp561nxjKQiHnvus+JxUlemM0FyiNuqBr3CV6Vcr9GrllpDX6x0
QvK0VGHTVBDIt2BGISsWTgwhQ785w4B1ZFeIdhDbRePcDFFCUAXmx6hjPwAl
DFqv1ODL+BteT6mrFsQ11kI3uKgs1X/E69QooHoJVOwn2ZMetiWhm+YZC4r3
GErUtBgUQB4mGjEEBRfK7bxU95HmKrDZouBv9xdgP0TY0CWoLYml+idSdlpu
BZmHgp3LfJpYWvIp2X7ev8a6cO8v6zo6QWK4/hriG+EGE0ls7JNfRMUwjj4o
hWkgxKabuSQdeC3DLyKbSi5i5N+j2DUoNC+6ZpTSsFalUn+RoXPNwOfocJWQ
s27G80KCg/+nsFYlcQPg/qdMFxpZ3fpWfENRsWqo/ILIBrI7G75mJPbKEhj1
KUGKQroV2Lew7U5JDN2DvtxqHu3GRyEtUJIReNuF7CLlZ44SAGPVjxp4hayC
m2gIn9lX2vpG4xxOcEe3N3wHrgQtC/vAmsrBS+kBcRSPS/s7RNonZ+/UAFYJ
jcts8F0C90256racYHqokVHcVrQbgxxErWPuJsEfgOeREjxaU+TmOZ2mPONi
eHZvHov7lK9GBvQ4CKtCspXW1K43X7iIqV02GehxdtAlFJjCrlqgQNju5OgD
qFf3ixHBgzmq+t7gd0jdqEwpstq3yHJQu1fvBbXBrud/2NrVy5uPkytO9Vl0
eQvThQGn2mv/tgeVJzIYYZdz4cbI6ZGc/OvJRBidsiedhRjqzXkO1TdMoO5R
VKz07LH0tBzpoylGSRPBMIYvM9gWNCqbgfh1ZB6H7/z2yUXg/EhuOPtNh9Yy
vN+K50yTaLYvG6aUJg6DBUPUNF0JootSxF+aP+cWq1XMOdWiobGgfoGYFpCp
Q0PtCvXPeC0cESvhy7iP4GMm0Tq1LNwlY2sLvaNFEwd5RXCeHyDWFmn4YDGW
8FmuYidVsBiv9NbrkZ2VO/avLgU9ytM5n2duIvLPebe6jmsCCSiJ4knccMQE
bmusQMoWIiRKcwNZ1s3KCC3iEmdI6g6QYqotmwu7MaPL30g8uVPi+Vn6alDH
6x3Zi/belU8ysQsJvgU2XovWvqa55hFvMyELStRMdQrcrkVf+b+kQxTvxmiX
h3M+J3Wvx//CT39oWyZh4B3pzWJDjsYJPf8PsdwUocx1+bLP/0CeexgVYxdN
UBMuXCXN8ayCICUIdnFFPJCAi5y2ydoOH8uOQwe/gqJ802r4+is4lTQVFIPK
U55/Oz0nCoWxmalmhvppTCaddqI3+abbULFvNzytAhfjkyroBqCn1nBq5GKy
4LkgvwrtZpLX7zAYsTh7F0mMFpEkauGXC4eNOKGA/YdVWMy6DV9ZnCPpUycR
KjggT0jvxo59wPklQYND7hpaba2D0tHVoGaXPxh/J5vqgiDhqjZBmkEBy+TU
K0UsgFFa2DUnXDp8x/iuSPSKcRF19Mw2iGUa6D33oPiNgE0CPZiTykBW6iDx
iI0wDqxfig4eLyAdhoFxK1dQQSspqQ1WQ3f8WTOlLmzegksN3/c6NVLdzLIx
53pXxpce3CU9UlqFPdVTyEoB+cr++6shl+eZExQ3CEw7tCyGC+xPWDESISwy
IHBv+IsO0nPRV39IN0jXbXFMsPmTwlPtpLLUFaX0vXYOK6OgJngvIbEu7EzE
lFwGyfQ1ViYNi6MI8Qmb+Vy6sAtr/+aL+DmdDLFwsBeu5YkuL/q79DEaiGXR
tU9Z7fQfyizQpU3rIu95h9m/fRsF8pm+DOFi6siDdgebxOLvKtRtxQV32wFH
cAn9G0ZFdwPXxGr77uLSRC5+jvq6jCqKFtRZRHFJ+bfCQl0QeMc4ZxNBwmaw
Fg1eBziW7FNqfOlw9FW9ITCr2DiNdQzC/c+mR6dIso+Uh58K7uL/4JH65MoG
qt4cWs+aiagUpJBWtyRs6z6M3TSGoKsfhZqzIcGTvxI5esSx+cHjjqLXcZUJ
vJVfAajgmP2H/ZJkwEzaXeYM/7ZWgLS3u+FxOdBdGoL6YhrGtk0EAWPvvBHP
vYRzrruZVNvMPgoWmRghB8tOxNGPQPvibD4VG/zBvm+vqhQg9wy36uPq2+PZ
Ocv8CPXHG4uw0Wuon5MwRWBHqFEztYfhn3cu+Z/ZSbTnv/a594gNQ9OcjZdu
Sx4c4HUTWk5RqrqQQVmna+I/99oY0MYr76hQk6/K0Nc5BtpfVZXeuHdtNSYa
tSe0aRyCNoxrT/hLbS3+25Ew4JFjH9uTfhNbCLo9v1wMswXSdfy2f0gvY/d7
iAEFWvgVqyFlAUSuPvxmc5PQHTJFfSuUGYd5/Ydakj5h33mAcCqWsFFaHC8X
vKAHeqCJUP9QqlIOpOA7Rn6LvG3OZIiPP04ViEfk/wjp69KOmqIlh4VNMOJf
TTa2k+4sJtqn1bFhJAAQn7IX9vUpDZgxM1zD5144DIusLGwj+QvB4Pmpqkgh
SFLcyW/cj21HYVWd5BTcgJDFTxxPVYXy9pm+60aTf+6qgMmn9nE6e5HukaFq
soaK08Mh4heiDwW/PoHdQ4dBY369L3K8VHX1LQDWvpXOdUJTcc8rzFutOzxH
nRSjfuYZa8ncvD7ZTWejEoRnfAYpTK5sjfJzIVOqTNIadchcnzL4/OfDlU7E
oKk9eQsZPV5PnjE96q+doiC3sgX3paPPIjDdbPYNpc17+XhVPUWyDqys8QS3
wmoa2/6o413NE717Uv+PhSf1CBGaO0ll0WRR0fGDNvhRWa1ANtsdtm7ePMTo
VtLNPgRlscPpQH5uktegLRPclNEMTiiA5LfFrLh/4oFvfidDWsVE+SFU80y7
nt1+ANxW0VG64b+6jX1zd2H6H6ctowJMas4gRGTKZConRvsLRjNjI8ivFjbP
XriL8E+arifEFuVDxINHvMyXXB9wdlaIezROD5uX1Y5DKhqZMfP9S36+duhg
fsWRVD77S3GtjVPPq/QBHPutpvo3tozxzMbML3Q6WODeoX2OY8BnOaaUFKnZ
hSLgYosKg+Yl/azHiA7CT81+o15C5q746UYhQV+B9lsxnrU/DR5mq5n4nG47
GapYo6MtvUS6YELHwPPoZJewxGn8IU1lgNcXHUxHTCBAfPSS+3mUx0jzZoNy
jIoRa2IKkbsSjY7iLQcVQkwZhz0D4KpEhTkd8MHZu5w/TCXR/2cNYirSYD1+
Nrk3jwxNdCQAC8ihOoGVwabZKTgeszRqtw4HikXQnSmkt3FcM4Sn/iJuQG7I
SdY1GVslgBitWPFSXdx4jyginq5Xspa5rshiwSDOcVAW5Kf/MODosVA6D8py
kVQAIc9nRVMAAoHKQ+2lgbsfoddQttII76Maph7PiWDILZu11+VsYZfQAwxK
tk7vPR0SWEissaCP7L+MyFOVoCP0G1FhfPFEvnFZDjONXq6nOrNeZTheXa/y
h0i1I9Gwl3+HwXWDcyB/sC7LsMUm/Qjp2KzIF/LnjVO06eYbey8qZCdSMkGV
VJ2I/5d/BOaMrGLq8rESvN/E2S7sTWxQ4QeeiVxaU6GS5ZFeH6CloMY2m3HQ
gnjCQZShLxfnlGp/uzmzLV8FNbYEqzITMfhUvSKZt5KJseZgfpZvmDFY2Or3
t9cSO7eA/M679Y8cx8L1uOyXg1Ud+IO+F1Z2RYSUubkhAz3Yvb9H/CZ4VEj4
oYr50/jzL6MEEtDN3Yhzqqgwx1yNL15fIAEq2Rvyal/JbmcwQUPiti4k0u3g
o2aUdyfCivmAa123fgnsME+NGQnyZy0vIQFx5MYgfhWf5aw2zXGrYLzYW78a
g93SzurO4m1nfhwApyKrJLNBjGtBJISKKlttMkqUFeQotCv5u3DICz+jQgZ+
jkvhCTEErCXRHmhCEm4Gn3GXVnnfy6+glcUaLdsezbFtZNRZJmiZPkMPD3ed
0XyRiZpg2nfmgE0rA00WAz/JhZ6U6mM5LqQE+zgFDczC4YyC6uf4bEJu3AXd
+ulmNoBZS9IIp2KOEQre3e8DnK8xAZuwC2dOVTsNvx9CMZNcRN2LUR+iT7bq
xdf0vd6yIi5IOUO54iT3RGRTl0KVoE6okEM+Hy22+BgAnHbAEJqf0pTsDtpm
aJckuNvvyj5IJv8YcOBZphAAuoPwvdS2XHJF5AEcfrDyiXSOHCj//xVn1VrQ
4VSfZGft5TD9xX0dXKfkdQpQeiseXsZYZ3kGiLPW4KspYkUBHUoMV+83TdOK
NJyvUsPFEvRz2p1MFN69lC7DZ7UsJZfs4Xa9eZO/hQZyaC3zoWqj58Lx9FRk
4XZ4uTXxT0KapwzsSSnWK2U4JXATQhGfQ/C7lC1bwiirD15V5CbSPabKRY36
o+tpbvmR9MOzNkGFsjwfGdnnFvCjG9YQxI89cOWI3juSMBZ+b7559jbGRLdS
vZZgXT7bYewdhdtu4z+e+B1+YbiNl+xB+zjUoWHfTqqdH/6OzIfWgYN7WBQZ
3qzIoHA8x0a8sqBKTtCgshU/6V7uE7VaLBQiG/ve5Vp8ND6+CSRMRn+Qz7Vk
G48Z/BhkHm64VKY8LlIWVFgpM6NoD0BhvKtKnRManZarMCD5TsjZt/3uMjau
wJyuj2gvH2W9yK58zT/pDSSkGG4Dc+uwD08HSdzgWU+O2gsyVBLYbJNtXdP4
P14SI6bChCbfGSBZ8nFhKdRjBLjEE27rmfL7yXVH0F5ilJxv0TLVydVaTmxD
XQD9W5M/j6HUmDNIb3ZBo/XESM6n1lvzwp1LNRuqe9TLsYKBfjG51HdzT4In
3gcR+Bp89fC6xPb0iCBOoGAaNM65oK/M/oYVRRMTxeJxEhBopuvvpcB+NiM0
tYS6JO4WcjWapFa42yz8fBccMS62j/fqKDDHAsCHuuETVmLcsOmPExW2Ph13
+3eTYF3fZYeJHSfNk7NDsSsTVzIeS96dAQNeYrcJj6rwzwnYr+B9NIvpfnHu
3a7ITo+Ewit/PU1RltgOpt5YufEOVoiOGyrOxWpew8Xgs67GAZiIIOC6eU7s
yvxn3+uxaV9bCI0LyVPrSLXlO9cFOAz/4/QiJZfCqiwmXfvSSrAHW5ZE5MUu
w5JZu339MWpAOFGUA7/XQMFeXYurWBU5i/mKgj2CPe2kq1ap9JnETTboTLBM
iIiF5pEIXCNK3WtpKIfN9gZ+wje8fv6EcKI0up5NJDPMonBO6ePM9Uaspn9b
3XC3PEw8oi4tafizykztW43MP3mklrAxN2VQC3Fknhb9Ncf2TMU5rxCdOL2D
WXtfceLhTx3i1+8Lc/lb5ZpAUYnY2bO2uBW5+AX/PzBWCs+fcfj9zbnD0PmJ
TOICOLwgjOTg6R4wWlaPxcL7MchueJElgIYBpGs3MrFtHy4J8djnFA+a4cB9
1EGz4rldhGZIfHs3Tg0NrzOC2mMYchnv/oDgJlxfv9c2RKBFnmFeXnJXOWql
L2j5/IUpUgJjKNROut2w2CPXTr+f56q7rlvV7P46dmiCc+rWCQVWcI435L7u
AmGbdLWx1UycZ/YPwN6Ul/YEZTCqBj5GNj/45puYD0/PALgwLNeWRjeIH47d
n8jjzRcdNXE4oYPqLX4xYVLYHxNORBFa6PKgSO9d22G4lVRvR2j/+NCdnVAo
Ej4OS/qf0IXsD0Xfe63kOOvtSZay97gWhxqjjkMg17gTimp/MyjSDvulxHJk
tnYvYbxdloMTFBpRvZyA1D28i212e2KZgI3/hMtKe7Bxi15uXRsc9CEx16OA
5DrJ4cKnsyhdACbKC2w0hoVa+c9KSqDsuKIUX7aXkoPhOtjCruebqTM5T1J1
RAHT+PfoSxiEVWV1hObO53IxX79aSX6UhL6m01ADVJOHH7Sj7bq2YxDrAwVa
/Ssc8r12BXxJF8FsgyCfVqDU9b+TxdF2OpWaPNmi1y2HZ+O8yP/R/SGA6gVt
5YQr5SIOobrJ7FzIFVft/+JuL986QJtFHAH9HoBketZMj83ST1y45VrJ3CA9
zjvwlcVvly6PQJB+2q4bpCuS8NAcVgLSVXaM+JgSpwWtdEqkMJ2yyQNitq1n
jf7QSffkMiKAPCKIDLA3JxQb1Q+nD9NLspbKl1J623DIN5xwxHegYOhy39F0
r9+7h4fGehHCbe8NmhPJsqhokaooO52BHvQhe/9T1f0tNe8znj2sxQMloq0f
VJNOHhMQiObKJ3cDx58ZPBMMQBOy0ZPiCaeyzIue/VivkVoHmjMcwvKwvVhd
2i+hhLLHLvNuM7F8uIKnH3OcGzsr8F73fJ63GnfMFEBbrcgzqWsXIpBUA8G1
C2MRkYmI2QPRSl4UsfQwbkeHYbu4T6i3t809V/NOck/vPnXBKOQrIXQRQ8q7
TINkpUTKc8JJUllU9QQMoCECYQO7GGTMcZ9dONuKXvE4XrrBbnxR2mCUcJzE
daEri5QeVFWJwgpKqsDwlahhVQyBFeAIZxmJsb1p5J74LjXnHGQdHhc5EuYc
5+Uhem/QIj0Mpxj9MYnOXpf9wu5/whoHDkiL2gtLhQsa27hGh3eqcdUTDFT9
mweuyhh9fPH58VjksKOG8/rJMs+A5CFuicU2el7b1Y867Qqb6su8FWrNMusH
uFyYySEZZ6sFxJ6GEVSUTFdkhqZW84E721M8fjvy5b0fBXS7BLa6Ibr9JveG
joNrmt7reEh7SqpJkcwba1Od72LGItfUp9akF41AOM3AuL8OSymf6LlrSuvW
InxvhkHrDMMkQnv2bJLihpSs9Ay5cf33ZrtIXGTIcy1My43u9XKf4Nix8kxX
AM6tBFKpOWhDaA0NM72hWSWP61XqbSpzDPTqqOM0ubVoXBMZh9FzSFJf7EZV
jpnU8DXGN8YS/5J0Z4/V+CoYRd31lllaqCsuplbPYbcQLdQHeoIAuspdLcJa
AyAwJD2T5Nt4fOZhVIKlIfstitjn5ISqSMl0Zdwcj5kXzFlMbpDZVTek4kAK
L49txDhT1EuQmCwKya7Je1qbiDvhXFr/X9xwfN+r/KG0ZrLz3A1SvsdwCmgV
pDygK7Gw/KAFy0bkQsOEYeCUoS5kQJt+74cOkwWB+tnCg3nGP1heRzJsjknl
xTs2KFhkMFYyn3jRQacEL7siI7K2pCi1Zv1GyVSgngER7Qxp5/9WN6UA1thH
oFN7vtjdamAmW4d5qoYzguQ/RdZoPf5p/cgM01hqgyfPAYZBbFguBbyHViD6
a1+wyPI4hRc2u8mWgmbIu1ydJFX+RjzBYAA5JUZu1mWPXpfK0DHskmGV54I+
U7N2SJVWiWXhvYgvZy/pYsAYXw+aejNPRGkEA2S7yoY44BkBKvdhkb8Nkw2h
wu+TK4iTllTarHS+nmbBEQgFwc9yRB6KPpWEzS7dbFirwQ4p/OyHrNJO5dD+
q3+pTuAUh84JkY6gCd/6M1AbXEfruxuP65AWJsWievYtjjtDrfhNNV3KgQy2
dNrTMiMhGrkS7piaSJjqBcv5kwG2y6lzS99RdBJmzbmr3elQhxQh+sFCbTNv
JekChkqzhf9ztSzZN6bhnAVMPO2Vp+dT1iLSsP19ttrZcz4c7K4a2yRVLvIH
ZTBlX1Rh/0BdkOChu1s8IszBDz0loV3kLJHiCJmHLilSFiZIYiOsKqd+bNzJ
E8EPzeLvBb11owdasSvoiCiHdTCMmFfyt6guphMC610EMJyPyjl5/Y7W7Y9N
/ZZiX10vMDKnlXcgsS2Vf+MQZ23oCoD6I68OEPxUDhkWXb4eAx2yhsu4ihrZ
UEzyGbqGHEOa4G4SnwzUNddpV5/ZcKveMpJm3IC7JWRCG6FCX20mpzaMiy4j
uKD5wizzKbl9M2z1Ye2PjBV/ipIwMz0ejd9FNKvRvd3+vro44AZ3b0r7RZu3
2ndBdrVREzS+oLdzlF8qQe9xqFxsknJPUtrJAjqJyFEi5G54SaL75pz5aoUs
yCsUWmYMamKqypfpbAyRIKy0ys9GM2vx0omrj1cvZRqwtrg48sndMCgqfmdM
GL+KVzRHKo5SIAllZoDwkHx6SRV30dFCelx5Lv/Sc5szqNkOrU2plCrSq1GP
YJcuRgDRFlx9x0/5CMKh7JYPkUP1kn4Cs8D72GKp6tT7bXkkqjXThjeZyloW
Yjna6G93YobfkvIwAFzGp6bUMCs9UizLhxsaIpsIBVKAeeD6lD2AFCE+QcOV
48X5MlWX5FHOjizT9R04Nt5zg5dBkGpdxiarfD8afEGSDWZrUsZ6FUeukHQ0
MUx8VopJCy5X+/RQxVJCkwbD47Qk1+NC+aYeH57a1r7LU9+4tWM+touCg0QU
XSLZz3djIuaihJSJhsWBFBlw2M855+2NSOSd89MrhAf76Dy+bIAYeukCrefI
EMVJow1R3Gz2ZdCsGM2ebyn9gBcL0JR7c7hkj8jwSyOdP2NT9h1yqqLQusu4
YzMqIQvzOnyTGBBo+y0HVZcjkxp9DSfW3ghjg0q1yIF11+K2mXKNgDwbIFIm
d9poG+PovM0gC9tw7VGm5rYOqOBxtpeIik9NJ82KqKNa2qgUYTslrgNBX9IP
XTEsxRfEJGQornC+dE2y0W3LQ2anYIPgxZoLgjNA6soFpWPw7835FubRixsE
qMO1olQDjVuCjF1oBkNMh0QnJKlPpomXW4xTgV6Rs7HB5IVs9trO1xFZSwTI
91rmvw20R43gurpSkjcISuLqn8ZvF1UiO45sjPikbKT8v4Hv72u3a+SNsF4w
1lrfP4FUya1IwbDHtQhVr0mosWDSP+pbjBXeQZLbBzmPLqttfFRLW7Renwls
9fkpkN2xCt8nUYB/XAJaw0jeO5Hq2tz/n2aMaU5sE7OugplbMqCneymoCePP
gcnmP6vlxmxkQzcxHQmzWcUQ5n9dNvesuNKFOdcy0U1RgfLm2RYDLEDqWCH/
wA55Cw18Ll2HnKOl1aNo/jsmuaTAZd/TICmL5Islm9jXZF1LgT8PAQb5XbBN
pdH9Em3K+WNf7fcVKfO42pYhxQe6scipPaKO0kQBNk2/4g/DyEN3hrkXt7s6
BjV1tsMae4TXgiY10BzrrFi9m1XF8pt5MbR/SryFVaCB76ATVlYIc8JcZAS5
owou6HZ0um5tYRWhfcA1iKX3A1g4AOuJaJVtuuCj7gjM5BDDh6euXH0ywthi
u2fHrYqLSQESNQngBpY4j6fDurvCGItGZLTtPoXY9H9fJbyDu7KSYzAQyDe5
Ty0vPJIkKW5nOyA+yJwXjhQrWozQIqtxLlP1p6jvJD3xC6na3AuTUH+AsIlg
D1nElhFVHNiONQHQYvYy4O0B5cq3fSJ/XK6Jq93Ac6DKi7UpG8vIFpzcgw3D
meYHrqlsctCQi8zl1vQxP6/7YaEfyB8vfPPWoBH4e1wrmQdBFRy6OoYgINQT
RQI+GVxgzrj8ofXQkPlW1/Jh0oMywrdNuaxCCLCffYJlg7NVuhxdw29qAxcn
NZ784eU22gtGUV9YGJyN6JHjvx5xAdp67jOH0g98KR6Ax3lPT7sL7zC8HWSw
UKLLs8vBHKVDoH0ArYj72GzTf4qgy7lUwzgvJ3B6LJfnOh4w1bCaW9y941vR
c3nJ/mAOhnjmNaYBczxRD3djocFhpympyZmN/Vwpm8rwLwLXL5CGpZU60ZIh
oZhZJS2cNsMySaFqXCSmRSTOkeE5NyDGYAiXfuucZdc234o/hfpP08wg0YC0
0u63Xn/H6Jf80/v4cvaLeEt5clgBMk+Om8+vrCyA4NtgC5xlPV27N6trJ/Nc
gJVF3JdOOFWqnhWvoRJXgrFlJwmX79lRjCCc/qH821+grd0/g7iNiLizldzz
bikR/Q9HndTQtCbE1yVBszYW8xXSSO/OjGGTkiYGAFKoTADkMIFUdK0rJSTW
rDfrsBl8cXuHacI/ff3HJKrNl26mvnuIJYGY9VQlzvKaW3+R8UCQUg6qXFfm
9pN3o0RX8w5r8pugZ5fPKmISf7tXkTURAEV8RbVkkvDfaflAIA3mq8b82vo2
BharvkSATNWXj0B8b2MDUt9ZRbxWn6e+N0g1muK1nS94EwR03Gr5MSOzc0iA
4b7yIoU+83zuZSs7WGA0mei2OIVHnq7VVNMCayVJqvEiG8Omc74d94+ZB0eC
j4wtCoyeZMuMn94EcY4+cwj9RJ4SenFy6rQgobiqmOVueCRGzpGjArBEwuNn
8iMKdRp7rrs5y1k3fPLyuNAThgoC5fb20kXZ9TUlbSt4DRfJbjgwJGLKn+ZT
QgMYPzcUY3COfTUbaP9H9HuFPdDATFVHwFLq9AiIT/PCTiTS1koLfLIMli4/
QugbPmnB8fWyUd+VrR+ywn4ejc32bKs+jr2zUOSyFzUprK9tn8gN34eXQlzU
eYuRIa/Z1wrduQXwB2d1ioNRLC/jBHq9dYl31EHOW02UXTwd9hNR5BQ167Gi
A6aR9D7GpIzPFlruBIABq6YEmBZ2sZtLE9WnT3whF3PFuTi/4+K/DDJDhS/Q
fGFJvrdUtkuKYWRhOwhPpB0fyMUkY58aHH3BaiOuMZDR+D8lrKrEJpAhmrQT
5iSVnXf7RVXectvH0Tq5veleDSfCEnA4ljxQTQFJ3ew6P0VpVHAqkGBSMA/S
YNYmNr5YK8ySQG5TLlFNw+NZSlgYdbJrDBYv4gf+UZNiJ58o0Z4yQOXPdhT0
pWNqg+ZIzok4SPBRkhu/Zroj+xU7CcSqS+VIkfFz4sI3nBCupsAIIPmls0vn
i/YIQciSTaz2AZHP86SyVdGgFG1QndhB05BzAGb7f+HBrXKiYM6VZj9EXtp8
winW7+ZJl8gbqAD2sanMdDL0quNsR32wpG6bT7UDodN7LKAyVGVHiM6iEkgA
kZHgoNM+a0C9VFyEFYaUH3GMyzRRkmRyGh5z/jxk71LUIQ2MOh5rEY2jZNN2
mtanmoMCGk/vtl7DKEyFk+XNUytsUPxhHmzMTfq/efUsg0wBiAiBZjEY79gp
7+w001rOgGT/6ZUSreEIplJWUqXULuskLqJmyIO9xUnG/2Y2G90DL1xXvVSg
u/a9MyoCaY0Qs1m1/nsI2vT4RMoJ89ONyLja/YqQEXx1z7H05UNhBtfi05zV
K/VMASKMPHDvKfQ74zfjdlm1ERiMFgSnJgrjOj6adhdygQYb+p+NATxdAD/7
bhPw0a2rvi+UT1EvJrN+mzVPMhk+YFjkZO6pBYzUk8k4puLu7zIq+9T4gMKB
JgbI2zmLuCj4uyXi3ceiX6XUudc8yqGvUbaw1h19raO1HgEOVv/+pTNw2uB5
D++r4nOmYRUY5zp/6Wgd/YREHBTckjc7afxxtNEtroHr/k9lnuQfBVf/rBiU
ZoEQv91NcX+a8vEA5JAXQ7YsEuSBRxlNdsPiXSiGWspBkfJ2IZLI86r/cTo5
UhizumBcIcOP79R98QsKJSWLJjcxPN66GAoU61ztUnxGC1D9IIQbv65AocMD
7o4715B6zz22/m9+q33SkMQ+18MU3JY82TS+BoIsJjM1xBlcq4woMSTIvAGi
kzOsKS9SCspO7Erk9HPRymUC7NIMx4T6AFIYKyeGOqdoWnhpchkp8Kjp28ep
HkQxLMhjGWruCkQfljmnORxoTKGVEGShWI2pKsDGsf4Ajl7xjASL6SKKGqmO
z71h0EWxIqld3WZq1CFTXLcs0wVFZSbTE0gwZoR/l06W2M4mKDQMcJTl+LIB
UmRwNi/tmKyHbsdtKf/pGwOJAMNFhILXuDOmOQHPH1QLbQYk1KwtwQj7cyzC
UP9drMaZFRCBLQJT6Cjg9AkHdyPhbDEetlGEO/RXi8EeswATQjt4pStJ4a7r
fM94tf7fSqi3+72A0zxSnuevfBUBQ29qyVXM1feHiX4DlKyvTl63G1qT3mPk
5cAjDjvJ8TEtAYS0aoY95CuGiId0Bx3qpotpo6hecuACX0yEPG6rzzYBA6B5
em8ppT34GFGBGV/LXA14++igDei7BKsiNEJDdZxk4HyjMe8YWinGbyHeWFYL
d4Co3bywBE8Uy9wFjhEAEKVjYB5FKKEPXjA+qOYJskgjwl6nnlTMZhXji8r4
bPB+QEfhYvYdSRGemho7/so7hlIE3q9sSqQz0YD/xMM6hLfKEA3yYaMFn6E6
K+QRntv+Ls2Rw2I07SrfOU6xz3zxNvy/Pzx5Cguo3FIvLWIcV4gwCHgSPURr
iOx44Rr+oW5qyZ0xPqRx8SX9DvnZYcMl8VLbpUsu7d8xaffGJIcF5IIiFC8d
glohaJmr+4NVLluSPWXiCdThVOIQfMheHQyetL0lFMxFU//0u5QZ0zE+hG2I
IN8osGiu+YyEfvt5NJ2u8nfFgnRo0T4EBfN6efdyJAw+ci6bJ+20CRrl3P+u
9EHZgKNCFdOUXL0SIeRJmVL1WyBT/raIaMKwEZIMbWYaIj2nHnCc9FBc/cjV
jPitqOptVhgCeDI0/wU9IglaABl3x4P7ZdaMCA2UpXn80mIBhk+0ndym01ez
xPGZTCJVreWOLOjew0dEUVdDxZOmTfyMj1kkhN55QJpMRclTn+eOLcjJJYLd
QtztQan7zHkKbuwhMn3N2PWDcHnNtTpOl6lpzwAR4qHOJaPdTN/24fdpz494
LOxruYZzrkRzmJnl62UHPu1UR2TQKB8fg5qymL8fXkS53j3oPQ3f6eRIbP5i
VFueF4aWvWkeVUyycAEWTDhBZgzvcPimGyf6cAKpEUnrNLgLvb5fnUSLAduQ
3Lp0KzTI7rlIMHrSvrPCAnG5kbkkS9TxE9m/ba+0McMnM5uDM526IsxD9Tsc
HckBEmYGLiWl/A9tzwV8Z/adbaDVjEvvyfuo8kGBgkosCfOq/xjcFWR8QkN1
BKdVQxVCUytdWQhA135SOpTqaBQXmKBzpFxmKZ00Vk8M1urIoVHN3fu7f5Jq
A0JQtJLk9OH6AVEgRb2Wai5pyj9fZdP+XVBaXb5PA7Wv/xO0KDABb0/2Lf5r
H00pfjza34JxzqG1uokHGaSb9Vdu0FaWvvUoTYUX8xXeQnaR7suD013FS0Wn
IuLTPHn/eJ0ieNpbHY2eL/JP7XeMQ9p39VNBIxLBJMHi8p4qci+mP/JfrcsT
bO2AAjTJzFOvTqIPWF9Xy/65o6KVh+Ioju0qOdDZd4WB3h8uGYxAYFW3H+RL
FpgGVldr+oBz1wICGyTMC+lbrCTE3u0GngXVNJPAlAWefbputO+kljMjUNZ3
hmfsTXzrp5n65jXEXeAmulYM1QwkUr9F5TrWskeZmQtbduPu2VucK3V46QOR
/2uBhffkbPD29AI5FkFEvU33StYh2ysCCg/qapfFFAmajMEHE6A0cDkIeKZ0
Hy/6P4u49NknkTHpxsIvVwOzs/NtSGvdCVPbp1YDoPKgxyN0kt3pzpFD+xvi
O0NmEXgfZEK8aPd+eZjx4VFY9BVt5Bv+PKW6NIvyDn3lvWh8EEhnJNdwmVcv
sA6pz9zDcSP2f5s1n6e0LS5IiGwyUKNIvwNfnX7kbPK9zH95QSuzlksoOuIm
FyedtAIHtWVrsdURPrazlQcPdV9Gv0VJraHhQp1QI1Z6soZR1zLYKeHZfl6D
dSoPe2a4jV+C5LgNgca6vwJFPh1hUQI5vYDnS1+kX7tmcG54s9msNqOE2oam
p5sT95Hf54X4Y/3ZLWvzzCI4p8rkt9wuYrQvN7fCpUS+5Z3mIgaqUWoe2B6r
kVyCKItHtPrBmY/FetFcsx1klJdq6Xc6J1qokRA1DrFGnuSHrOuQlHDqtptR
s5hm3EnoONFNmzBcpB0NSYtr4JV6DuZxd0hAx+iAAzZGnMriuLrA4rapSXme
s0dd5lt/C2LOtARQx7sf08JA4/8dhpzOdHi78pjbbwB/FJMBH0OQG2uHLLgy
YOoh+QXoP0iJlGkGXCSstC70HJxxsG5BrU9saXmjBBjsXGriagZsOl51uayS
x2l0GRzQZ4GIKD53R91GfybzN53eoG5YvLD4i0diy/TuRAji/x4+FWFAAxhH
N0FTfYrX9SB1z1Do/zsa+fzhsCoVObrLpORHupjCP0769IYuhJcEsh7UjEwT
8wKihEUsVdQXQDPmpG0VU4QNRPTtStD1NQuStAZTwXDK9V+Dm1wkKivHehbI
OXmiK7RpNwIZN/IIndO6m4ZA7joAJ6dxFjYp/BbATHEcQKSF4RnZD73P50WZ
W9OjRUiyc8uEefMEybm3avumy5f7dDabzyI/MtUiLAQoecrkCSk9KCAPX7cX
w1CwBCBmYgi8H9ZXbWW5QTYJrchGnbm1ktW4Yv5Ey2ZC33YGJUIKIWBYhfCg
BkCL3CBjdTXiOHjV4UnYQ/n8YcuNkC4+eaWxLSO+ferWeLuORj5zKlmho71n
UgPTdK3fEWNICc94Pva1uxNwePHTG+6yUQ0XCyFO6bjuWLcnP9OvGJd+7AMM
hOdS/tWw5rCgFd5l/sM+/5rkylGwnhz2LOSZ4+ahjiI9s20SaZI2Z9ThQaaW
XerUZgKr+re4GtDXRXRlKPXCUPA8WWkCqoOIXHGjbUBuQwmoE9lEMz77wc7X
oo/H8X8SI3qZ+d5O+/gcVjLAXFFSEiV2DgwTCingeMxtm4Ly1FgbT6ogqKxF
yaybrq4awHt9yz8/uugJgdBtWPWdlKU+XLaGgh2FopMpaS7RUzw7r90KUDbs
RpQ7bDK1GdNbM/EB7ZALVbVrQlI9Sw4WelVBGsnvPuFE6tbrQLrcGWgMImJJ
6sQabzbSKcR7qr3Y5hiR612Vjwc1drB9/bsT7xD4PIycg7DNQpIMWqhsTMqw
Tg7odZ97KgwQkaqkQVEGxQzcC+RXEk5widpgKbsKUq2gsIt9l8Ej+GyDuikP
o9OjCdgO0mr3RzjsbCuOsRhOx/yeGUv38E+QadjOs89KF61KxhcU9d/9qpLN
Skqo3J3IpNSOLFyGEo5B5DAi9CMtWJjD8936LLU2R4z1aCKqD+gIf0qInzc0
4EKRR+kl7slpoVbE9PB754VWvW1cZAgOo9lOcMkFB+WHPzV3QtlHHA4RSUEp
8pe6twF3lwCecjfw9F7anFQb7FE9fKXK3QhGsntGVScJdaaqQriY4UJRr5CN
nZdCoUwfn+VZTf1wmU2QQdtaKIDbw3UzAp3KOtl0Pn2I1JYXaGEaYKQLS8RS
oK3uER3G+aHP76TQ4B+QEoKQtVqfVuUDUfTw/DSK6Smy9CuAWSZ0iXj2wL7J
Rj2scDryZu5ybSU+v1Zr5vgEhYGJNpXkFkPuWwKfXwTQPcj8nyA1HIEnvAR+
BM7PeguyAk3oXunWMdk+q1ab6jZPYyFXiLQ/htTPLTnB/fthDwaUFL6e12Go
kJSxe7nsS1qzOGWChaKn5i3/CADCbITUnwKxNhF2qH+GrKIwxyQQCF4XjrCf
Vky9lhDPFFvF5qbDJK0Gc1d3dt3a8Lyuaoyp6/vwatOlmdTxwMdhxlUbrHBZ
FkbiCIEshKM7CycYlsaEc1AkZUVSMr7ypza+AxlvZgXWaOHSlyImh8yEMyu6
IJs7ANAx/Soyz1aXjerkbF4SY1cK3fPajIRh3/SwxXnO9pCn8utJShTffmQl
QpBPZHuv+oIeHZKUZE9em5t2Ldg6njxq7XvHYax4c29o//jPLo+43cXGY7vj
//Rh2paK2UcMBOvhu3Ei/+G9X0YgiLQpf1kGT6WL9sSmQS+A6ASSFuNC2EzI
pCHN6iKTBSxcXZcWjL+yEkwfw5AlCjsNvSYAJW0+uRC/nlgbbux6ct8CUKoR
wpxqOZ1iIbl73ocxFdVfKwZb9CHMynbcucU9byyLe3aqqLGjm+72j1fOBhAo
KfJsn3T/4UF3SpsLxxZ+ddcMylCldxJCAIh8qz15vLDeloRQl4E10Vh8FOBq
KyW9lJA4r5Prg79bjVTXnfGAQgg2d0HwnK4R+dar7t1lJZ3c1r6LiqREIfem
5APf6Bb1qt4f4x5UBDsGmwtcqEnEi4r69mrwvobKEDFhRm6QXuMe0xx9mTmp
eKCHZcK4m1DWONg/lZqwsKkHg0tw0/NfCfR4MZ1OtqEWU31TjMRaTXEvoXdl
Bm0pZpb7jkpzY7oHygz91ib0gsErA3GG80peRMqLy0geGlDwBkpKXFIBs9HN
mqxGpwWzXh5LRL7OluHoAgsTPkPHWpFaJS6zfh3rz5z1gsR1F4SPrcQxBzev
dF1gRdcNjG5B/maVlBHNPIBHru+jXuX7UtQfV7aNg7f55RktL/BWWxyTq/jn
ErcWHeb0lMkWctwYXymkuezvvzgEMkoiEr12UwWbgdBBXOhfr0Ofq+q+nfbc
z+7calll8eGWO+UBUTJUphNp/Ap3zOxFaxHQMUtkxKCwaC4PH7/W6euUCyVF
FJp6lHhhOkP+6LXrPbVCB2aiN8y15lJD+o8/5uP6NxtgdSedYR/H+c8fAFXa
CJeRXASqKv+0Dd0MkdUjyLIiH/GC/KZgICT/vz2eQr9P6ynzGOdBMo4OY6Ca
Xe0QYjjd6WYSN3wICM7VIu9V/xvVZr4iijB6moSjaz8yxS8goCMSEtxWQrzO
fCSTy26NVE5zmB1roFQczHtkR+D+Eph0B8G2kiL+UsyYXpWLnDOz2/wbjb3D
zKUdVwt2Wm4BrqKnMby925F//dj0Qsz3hurSCdnS1e7WuV3pEdz6lLks5wlc
KT7yz/l3WU0/woNOf2LG1RlxBvb12Hiid3hYqBOP4sYp7z7nB1wOC8N1I5aQ
0R2Bp8mvjd0V+1lky2/NVF25joows9DL7Pp2k4klwktu/e6yq6i9mAI3cr8G
Y+gmGTVrxwRAALlyDME1oW4rq86/N4rzAcY4tUHE6nulnlDTQNvAQfnwu1Ar
XshfsdPV5Djrx4gkhJ1teKgE77+byigvFL6P33l5+lCl0MTHaqSjGRi9vcUM
XCyfW4I5+Nnpfet0gNNLiAI4uJW93vt6Nm6EDAVPIh/6uLqtAEmUrA93fkvQ
q+yngu4UQlbArnxQtt7Es1bcq85Qw6R4hZ4FJz5BkWBFxB/qOkbI5cCJEHty
1UFeMKU8r9qmbomdnSonLj1xtYM14Gkumq5dvz0P6rX7aKDC7QqkAsuX9gEQ
OU0U/x1KCaTOPh30qQ5c5HH0v9GK7NANyZDYnRmqpoUvZ2M2oUrY9SxBMMz4
z3cZkeQAEhCU6A0qitZI52qrFFDnC1EIKVson7NFZggFzJ54g6SfFRAIfva3
I32bclDHPlcMIiB2MfjR9Q7FVxlvUYBo/jICS7icrwQbUMPLprMrdcNhBwXO
2FMruhaFXiwhTBJa5p/Y1v1UDguf9ldZwTzuQFlqfb0Uxrdzdm+oknSoBnyc
DJTwNFJ0Ubp3kvpYXxiEI3MgumLh405MhkKBKi2EUqZGgZyMlvcPSXhlbnU1
jXWFFnAceGmr+CkZHPAuHP2H+jSVWaOCu7YbBYqNb/8Ph40cslGTsqW3MQrw
/HHk3Sdp2ladzJ/voSNGsxcoSnIRkg7GQboSuZkSjfCS+M4TTBLSTLBnsQlx
BwBZhfzhNXiTzYYNz+ByWdHLQ2v8HZzUXqbwLDom2Ad4c2a4bdaRDaPkp28I
VMMnkGbN7qaDjxwgR+xN2eKBA2PPOdPXvC1Rb82X6ZRxgBdUJBWODSd+BMGK
bVUT5/6WgdzN7qxfeow7hdWoiD/X6k3EKbv0WkHcWuST4XTYu94FvttrqPw2
cg7PB79M6i44UmH5Jm54+T1cSeWeuogV6sIGGJvD4m2+V0SkpYFG1gTXORGM
X7EmO70tGcvO6wl1SFCiiRif+Vhfm/W0UwQ/G9tf0Uih/JTAziCCROnwYqR6
65SwQ06t+N3Ycq6KvIicDRS9sB0fcbgz87S0Beo2e5oXupCGjbdBgx4NOKst
yYvRGUeU3KMN1xCoIp+MDnUxmYU20Y2up9zwKHK8PkiD+HT6jHIqiSD/rH+F
Og3WcyAkrN+V+KfymlCtfrKlz5fX2hqnbV5jt2sRkkA9gqz5w4c2g/PaAqyw
qmUt4LBwVqH4glzA7MSSN4+Gcs1iMkOEtgiB6n0sp3VmKE1RtHGYCJaMn2mt
Hyvn3UzPyxOk6RAQurpXxBb0zvOh6bIIatVDbgOAm4zLDIc/h8HSoLLttO8g
sXsnPCKH6nzSN9d70WnMtdsF8q5uTiPZRFXeYZPCkWXHeow1qSo8BlBUPWXw
hQ5EB8SIF+Z4eB9FEyVa+ZutLvIEIukpxicOiuERh671/GJtsP/vTd1QZP7L
za5YEX6wcYz8snLR4yCVyo8WDuGwBNaw0JrakAo3XhZzsxxl2Wu67+oEUd3o
gzg1GKIs9Wi2hmw3SvB6AjQbQ/E/KXnI9uOoGJUwDxN27ettyZJgOJO0419T
2PDQ+Y1x0T1GWZ9RqFYNNI+zL51omGLqRM+hcEdy1mQ5X+XmVq3GyvOMPgXX
V2gwyT3ECoka8K4yyGpCV6kl7WE8PRuWdrSNataz1Pf7BO3SZEL7EdWxqoXU
jKkU8Nf8t7WnBfVFHp/0NP9YmCVJjNpBx4CXyg55xeLcCS3szS6zy8Pp38Ai
3/xsPqdsM5o3kUhyOX65ACCeHlpb789CX+ZajePTPMHD4a/+4FFsjgDT38XW
FJKe/H9lnTtZxOmdPgWzPLm6RC/5XkNZsL0Y7wQpcmrM9Zu0bw0ZO+Ax0LSJ
i02atx0YxRzs0ubJZWtuTjpfTYX34IYJUh1sOqzmAnsD0ADPhW2XaW3MZ4aM
/Ng4eUNSXCdCIXk3kBAg1uONzmUTJ2Lb27vOGDQKb82crZVWE2zE18ddindu
fPBTry5oORFwph0U++QS3uHWfpO8eFmQ5ZjIMW7HKZJldoNJkPzGoyRHJwZx
J7cO+mukUdhne+5P5QKdCQS2Lm7HhnEnRw98vzUcgakvrRSjRGGbdIXt8yiJ
9lacdg4ZhBEgjZejTR8YiMOKwpmGfLGmeOGMQD6I8OnQtqJB1CBvlefltdlH
VQScL4oXu9UIl+SzZSqyVfmMXwwVIs1sKvJ0K6HHYJgh2e+9lujGpSUg9mA4
0VNn06CZAh/8wgbqzubwwrgnAasSB7vT66/qZN3vTe9I3NQRpEGj8ALpivmn
lrkdcP7VIuqcYoGyssZBExMB51jEttAp09ZdIfdTmUh4E7mqBmd/DC7gdbPv
1ZIjT9gRu7vmEu+qLBKU4lE85yYeB4BxOdrhnrA8q1yWG8t7z0yU98j22Aw/
SLjcmekUio3xl8u2rGvVda2TCSwM0lmurDB3YSZt3SIFS7d8X6UIO7VRSIj/
UMYFyc8VJF4ThEIrfE4pBzkLVu0wn3sjSHwHVyDmoV3/3cFtp/zORoxp5x9J
J9m3OuCP8lcHNSKz6K++aATDQlxenWV8gLGu1Mf63x6yTbP+7flQjN9XBQqs
olqJE/N8/qK6gdS1D6ZEykr4M9e6OCNqBs0BbRaXi6S93YSAoDw+x9SjA282
BKE2PEEQKokPUfNlx65RRKU4U+hTRe4Olg0jxdyJjEK51rtYJqa2RrW84CMo
pBHG5CDMxWAanvucS1Ufj1FbvyCU6izc98Qj6CT28jHYNrVgcWdTt6kZSjpQ
OiyyzKfTFAukHbFbXt38Ligjl7+kmMqU/Rvv63VhMajstjIzKMr9TG9xatTf
9tEtagkzA1rDgdnNIeBvI3H22O1ED/s5Ls4I+vdPeTL4XpnkHL7WIvt4ELUJ
IjN1k+ch31rNA1/+bSka2dASCH3zCCQA6/WC6VWsH92EKkYNyrqNgNyk2RyX
zV6rfyVJSUE2+EZ7zv1kMncI5WE++tEAIRlpjahqhSOexpgNyHjncWo0ZPXO
NRyDSUWOUqBuSqQleF28WKXhV2QKe5txGnqw8sv0ts9kdq6TF/QD0SaxKuxf
m/a5XlMAZ/iSxD+ConZzxKyr09wRY8r7oAP1YF2WsbIEVWjETp9lWxf8e1Yh
0zX4wVUp/pZ2/QZXrap9rVRg6BpWlVevDGaftlyoEOZ6VHGnHk5n+4tYR1Xi
MMmuTNk6Xpndc9zGsdlGmmG5L9Yxa0TG8twwchbJpQJFpvCsDk28Xi/xhUow
Y805T0IsE+FGa1ShFVsKF2dNio00I9bDyactgqB6bSh8S1F0IfoWeFjKezRP
S9ZWzMpecmEI7EmYFmD8zwSu5Ixf1gR6M+SRwW+W4GtrNmem/ojzs5DEiJh0
q7hJYhgnThocFVbJ/hq91QkiITSLOFU5skxih5UyTztlzZYigs4Mm2QS/BG/
HMOs6AtTcbmKb9HU/QUiIBE8pRhuJZGez6/GYa/6CtB1DTBpKLsSILO6tGnm
Of6wxtOHigyiHbb4OZOQetC4TUtPDzCKg15Y1RozgR1hMa+8L4f5FCH1B4Bb
SuI7RKuni1eTOCgdXvdfd7ual+R+H4tUbLS3TjO7AF75sJ4qu8SmyxeO4GLf
/oWzXnHIjWOsNCJae7Ie00wmJNdG8tfBt+3fXHQW0Dg1/o5yFWUBZ3TZ56xa
HKIQd15IeRL+R+WyGpxArxw2m4z1SPgPBn0sSAceyw8P/cm3IK0EwPcxn0l/
gT/g2V0XhxMlrci3mqM4r13XKCquqnAukbDYcdFuckQjWydpe9U+HknoE4mE
tAO12LNgJQa1ICFQc4xqZiB68eNlizGVT+FWTH5XtgFJOpL1ze+6e6DFQHDO
YHy0luEB6H8EMUWvBGW0heRVQV6J8ledW1bAEd2NZGhR/7rczO7qloz3JjvF
orI7vzzsq/PyoAKIzF46g7OAHFQ4woD9lXo6uig4J2LBc11n6fB8T/EU9akK
laWuByysppVAGDLXFSSg5f5bC/Io+qzAUmzBQa+Q5Yxijn/ojjg8VKw4VAfk
Cwrtvr7ztL3ssNfn7Bl9mGseJWAQWQ3bNKeohA2WlZ2esKiJxN8aRKc1goEi
RPjCtIoC5/5E5kBL6X/KKlSmNUrE1hg/z2W08PEFH68n3HowxoIaIcEsfIaa
v6bRV0Zo44fMdZZ9Qyt15tsj94wD5zpFLU16zfB/hXJU0InfzudbbKdEPzKw
dTzST3HZoLRqoAD2/8sVHXQNUpkxrlO9A3GYZeQaXhUYWxXHseuRvbIDOlNE
cuqyG8Hd2StTfLfm6magxNA3ekUUpylxPZs4Fb7xNgywsFFCC3T2IJvRTa6l
RW2HsRRT3ZpoUmsWhQiR8nEQJ3DASHuSeg4MZdwDB/4X/JjWHv2bKyh6kHrh
UrEWYIRidnS0TNG7VAStFagwoOFLbj2xUTj2ubQtfdy6vnSRUQm1rRcvsOSF
pFjUr3PNmt2xPdF9jgvq3IxjuRmdtPrNBnrTlri+T3uUjAjsBCFsbZRGli6g
YiNI9UC+LKub6hzd1yRyIL6Dk1nqdKPCKhOb2mHx3YiNHvezvkgWQM2wDpJt
TM11ycGY4MnxRzhF7Tr3zrYHTv/iGQhOlqOoov7BkPrKmD2osGJZpcNtcB/p
WXF7PQjvRRuaaPrGqxJbkFhblNWhhpBY86gB96PXjqq1lFMClr1gQ/lPJIyx
6r7kCXFdM3Y8lBKzYAAI+aAo1LIbziyPX75EjB40zqiGx5CwRxhKXXnYiC6w
wyplAxnOdYR8Yh0ocK1fDdDSfNTz8Ol8GqJr6eWo1IlkwmUrbsnmctQei5AZ
yx7LJ0kQuK49ClTVTCeGu31DpYs5HkypZt/78gW6ek5Ta9cuB589QSuA/6U0
NlcZxcmHs+4VLzLArZ7DAZzajtZ7oa9aSc/aRh365uFaMzvHjbicxc/D3fzx
FjhlWpomcDxltSgPbf8lA/OPRnOTACUfN4F37kGo++E3qV5smhmeozITN3rA
9j0E/vnTLOU11dcHUpWnIoRngIY8z+uK9ORX35odXetOMw08or0aayi+RC0k
V3Rg9QrbeMB9zPVeOE3Qf41q59uREJHVPBt8NUqXf3W/PDR1NeCw2ONpcIt+
Lv6jmT4C78apFGupX9nPd9Pm/4Yp7AEDSgZvVq1iPoGPmWb/Vv/wJ3QQHa9b
qhzouhORYvfOhbiospEQsIYt5R/SDSwcQ+OalYDDWHrOOoER3sjOyqyvbSB7
RJnc6YhIFWcXLJTmqiXEBUh3GIlr91LaNMyiYSNplvZnjb3qKoKGNRd8QiXd
f3SfGs/kb3Vm9YeO+rrzXz2eteKLV7edhlcrHpsjfr/wYSQBMn005DfgrrvX
ce92d+/CAYs6iHnzn0QloXWCLOZhWknf9yRXKtuhQAHsoJvOO8lbDEV6gMcr
rT08WlV3+tyvvIrxqf0bkcRoNb7GL+AvSAYCuY4h+8FCgTcQXkTdEytjxIOI
c2zvqT8+AuEl5UafQGYuyL2+sJfrh81WiAGMrwWmgASeydbcdxTfi+27E/Rq
i6cvCzvbCPOF1MiPusioJMLurfOzkz3tAJxsna0BSNyf+i2adXcNbMrNHyyf
tCz9o3AfMCTYnO1n0d2Q8heiISjFJ1m0s8RneUxilDTPpAuc7LyfscnnHrf1
bk3Nk+hZnmfMfkc/dQmjp68Y2ZI0foF9FGRFnagptX4K+QGs8at+SYu35vH2
BtThL0CyL1XexvvcHWtoGkgJfXlkfiUXdbsVWVmusjYI6ppSRSvQ5Un/g6xV
D+QqqDVJPjH0Gr8bOMgbyfeD6PtlEGlV2fBtpdWYcW+9y7AFFlIqvc/XNRV3
tYCar7FV/vIGFGkGmmZlUZFZR+4iyL7nDad3p5TeaE2YfAPB6Xx4LLFUKy0/
tvw0ppzv4M3T90nlJElcl4DrgYwnDv7ADzZ6I5ZX9vH/O3xwizn0K38NgpGA
uszFijUakUKJuwwFF7/7tk+yt8TiuV14MyJH3laXpOV4UO0Xq996tMYKWfY+
Vf87NLJV+cCtpx7/PR2SzR2BTkGCGseZNsUHCjz2/qWGjApP8XAiwF4w7t8v
3ukY3OgaGZefwkKu0cPyLpY0kcnqZOJ4asL0YlIzqib1g2cVicLp/mjdjnb1
tfCwdRp6MEnGeiDJLDnHaPgala5iuWOtum/hYic5Oya0PooJ8KxL9EU+auyN
JpPwNxUBtPiZwGI+f4dvSqngX6xhU/UoZu0uUHXbwl8ua7w2rYcunjgszndc
nV3/gP/VhHib2WSO2pRZGDoM2PZqEx1XXpe/Lo24YNRDsAwU8a16cdHNyQku
v6/AK24q/U//9SYcPKYi4++auafQr9mynYFYYYbOY2glzpsFv6yY+dGBfazQ
EwvXoFhXbitS0k4VzbEY58PyW2lP4ZdA+dj4uPMvBwsv3hsimN3kINvAqvRU
EUqcGyh5T+/tlfsJ6g+3HUiyBbsZiPHWXxZHC9Oa9nyN9IvZ0ZGxIuRuuFkc
bcympSMTspCRUOkLd+HaBvCKgrOKJ9xSu1Kl3gKej/nyhBqLGZQ4byzurGqo
fgqamSHqSIwYYFnpHMG9u6Bs+RDfvRiJRRDGeiSc8sn1BW049MwZrOCZR4oa
np9Hn3aApZJsh8wVgOMCZAkpq+5c/0p5GB5CMVfkO2TBXr8zwDiFixHEZ9af
Bd5pwj87PquIDAw3bYLT9w5V8iXRZ+P+yj0dFzhREEf0/KOdGwNGB1AuVpW/
8tnovixdFSpPSHFN4DvpIwuAAmghSShTW5amwkgkAfd60YdLbAZKM/pHU+KZ
9ZNgggeV9v+VLKBtcv2dJIDJyeCq9gi7wYLScsVA2kgkiR22KwCT5fwXBRKT
9V4DJWOsStXTPYBGNQf8WZxQ2QxiuMpkig5Pq/ICamhVQRpPLr4nEwmwqZsR
IVi/9Gq64drY286cgThDg2TmNBtYcjW124FOHdu/bR17w9YojWcNLdcZZw6v
4TJqAwzO114MsPCXyPX6NGdGBu6HYf+qwsSHrQX/hTnY2yDu++RErHhTIT4i
TXfnmBrvqnbV/dtPLfnbz4z77mji/fvTueC9rzODXsk0koT0x+WEA2ralTd1
xfwZUkbWxfuxrWN+skRz+YU0IJEz1f6WyQzwKPhedLXSLfjTDyBMeW5grdaw
WegeFD8d1Zj1CQS7lEYDHeuuxO0PGGCORuYhcFHef2I4COuvMBytC3hWLrbg
ps3M0n2EVu64NZSKIcauHcoRwZoRZKEE7gMx9WH31t5AsfdiTuzkx0qmydml
NF2o2wwMQCJmBZIOUIctu9KZ1yphkWXhXzl8YGsj1Gg1IDwXfJ9FaFVBE5la
9U3i75ybj5AIsnmcd6KFOyBnkcz53kv0DB1p+n5k8p2PhGL0eXA9l7oK3lRP
0Eiadc1zkAvhFKRuuyfYyLBCIpvzNOJBmYTXSJTadz2X+t7YyOkmUFXj5sCC
qQAD616c4L+E6Mf2xJvL87ft73nS7Rv+ZjdpfCReL3do49O5XYEMlGG1me2z
dKfZteNejTnGxf4iv7KhaxwxzqtDd8C74nVuJBYLU33UAfug7WaWqexQ/BUn
LhwSmLG1RIFoJnWn0gYQnL/XnEE+DIcr+krLWnf8qH/KpkiQ8evjqYSN/zXH
YXQGwKwvHZq6+fP3LkaU4WnP+DQplktcftBfHBcjmky2YYCt3bbDbGg3keuW
aa8K/Zp8EukE8etRQ3zXb9lZ9Pp66M3wRAM5C9mNjIe3DyhKhSvRSkii8MC4
WoMyqUl03QWmT4hE21Lu5UMqO3VasnTEq9gKH5PHtE7OELn6whTxkHUFnB8E
4km6Lz/xOnImUBX5psb2AZHV8xR3oXFa25mDU+zS920wjBfaYYuOqqwg37x+
MN9Y65inmaW1/F9++i4hhAYm6DtRMzH89vzKW6rCWM67C7cHwz47tymeXMWq
dT9voXBLA3uhCH7LDdiSgFngSr3zDXUFqnFLKDFfNGc8GmBH4rqrglKCmBVX
PpyR28k3UpEJ7lhhra8pwnFkbbdADhY7Su2jTodu76qwTIpufwISS/3+TGIa
0quM5oWfedjUZWHs/d6ANzOePebaqDqVgB+qhO6NaYzUQK0/BZ+2Gd9twjVW
UjnkIWjJKV1KWnX+d7dOQQvu/TW/kbVeOIpU4zDkzTuhvpG6q6tfjLToIG7/
DLB+P3ekLNUgn/a+DdujxtJNCuNYonv0nrjVowEcDVv/ZfTRPn+c7MkYIJpa
jJ5+xq2XxMn4Hv76B6fN1VZFa0ZY1EDuJWKf3gGuY4S3JNzROTPdwHBlLkrK
19N81OEMBRbtO20jMc2tO0K8vI04P9OAIcOeOntmXVRlQ75PBz1hFLkJr/+D
G8fJoeYg+ZvTX7rEjU3qknWHwflqzTEyV9Ta8wV18SJtwnAvQ6u4/rbm7G8F
yJ0Cyqy97hR/qvHLeoM/SemklyId/XmebbfLaOfgChh48X+AsMJW7GK2Tf8j
vcWkggN/mlnh8+W038rTmpfxpTWROawnUldkGIUvst9jZwZjfepxMDMapWQW
KFw2oOUs0UCEstToYfHm+T3jvfJHL1BF3QUaK8GTjDY4PpN6S/D+PgRCNGYP
IQ1Yrf5G2QVEmzQuq2qm+1mAt9/etKptYX5FK8FQHKl33wXhh9qxXVjOtI+s
PeJSjGQZpprKnBflhhZyzZqS0Y8ksCZNn+R99dvYqMeg4wJVH6rllc6wbJGQ
/REvoMshZrgJbZ7EbRx4lS3wc3832NWO5QwWzIXYsODQchVT0cN7j9hOlXcG
Cxxq/i2XBZZ08xde3ejTL7QrAWhXJcp549SBYioNUB0IffXW0DdembK4yDFT
LDymOpeAqY9B8RginI1k6IV0q7JkMr9Wr7gGblJJRiRFA+9HWHbGKyL7PIML
yu9bgvqAd7Y3YL4lfsbEsVzpMb1y7AW3oD5wIYUNWAfnCIYkegSIp3/QlGTe
uDHa33zow/r9PZlv7tWgulhRY9fWRiO8fgd1eLAoOWKh1/d3cQNQ4l3xoYg5
XW6VuK40J114hvjQ65nFf7L+bcxhLw5PaJq80NT4SsGUUsQEfdkVVltJmufg
+D4OCZrDEpGcqXnRGQ7LXisw5o/p7g3r6I+Zz6VqDNXFx8qVaZxQUg1rh33r
jUnlvzWwJSM4KEs99Bfps0kAZ7Qe/pSJiLT3F4KFBJtzU8Swx4ntqizQDUey
qTZNsU5aUna3JX7vikyMIVi6ebIxtieSgk0syBAi1k5STBsoKCQzf1hisP0L
+nf+6u49dhyolfEwmOyYFdFeE6y7gigyKz03QXrCf+8PZTr5fkEq/JhU6cSM
HnCeAYpB5gN3FjXzqOkAm9qxFozGe6VzzBWWzlaHi3RigUD7AFiqAyZ/K8lU
ss7kQ00Mf0YKWNXaGcXAc6NOx98CFlfzLW9HhOk8yfaApEQp72yJ86pDTNIU
g0quoTqfOtGG9EH/M/1uqSXcTl37HHwOc2pcApCdpe/CWASoOSiK7zeR/VLE
q+hIAm4SkxpxAZbI+vRnQGMklEVAaTxnyq7ENcvP/7Sdlrzq+mDPlL3BXY/m
PeleQ170xNHWx3tnypv/ZBVjXkgw0L/qMMLi/oQLvC+q9fXVn+uoJjl4N4q3
zZEP/VE44ObF5ulQQa284lYd5wS5x81+HhxUzpk3bLPZgqKKT1ZGQwZa7zB8
bNP9mAgYgpSLmxt260ZE3p2raV9jolaztQ64cJ+H6Agx1a8FgrK/1++X3vk6
LTYyJ3GSRPKRZDUEhtqYQ5cXC47LQQJt5WGVJB2XgzlmctZPkE6YKSeGGLBl
jm+v9CKgiUakppdUENw6Ey57vWkCcviAeL2TlQr3W436Ep6RwLsHffItBS9n
C91sW3UcET1oiGR3kwG516DLYuQC6uerPMu+LKlUipBt8iY5BUurngqJJwYa
9WKmKB8LC31H76X/mfm+stqhv5ERmrFVKWUDhturMvkfBZBtVqGmYZWtMbGC
bg6Le6wFuGiXqvCiHLcWxybO6w82x2hO+6WtHQ82f3GyoRZ9U9NLKU4YjW+r
r1pGobIW+az42XzM9gUXkFt25jKC4COjtqpba0p6eyh7cyu3lfbEOIbB8V06
8wZvOt2FsQ73K/OEVmBB+pUWC+3my4feRDh+5Y5Rvx0FPEevzvNeh3hPHRy6
uuHdfr51UfHhnLhlusSTxGv+iU7WRXoHRY++zOZzlg7Qgi9RHMaLz2bVFsRS
JP1/MRM9mvEbbRKubNaLa8nK/hygbSFiEv/iBdE2b/jp2ffBhh/qOhkFnRIT
vY1pcXi91dUrDWwXTazYnd8EjKed1kdJjj9ChpjLQ1wPzjnXGipTbxgX+cLD
spn2V4oAcoLlAi592X7hHzwXj+xGCwl2jDQEQE2VoIn5A7HtQ0W7QJBa+iJ6
E7I37CyuBP7PZNYNCj4K4gH8/buVChGRZFqYHgfY/8PeThzJ9Ztiuiwo0G27
YDEQakM/BooAxagf/WNveXqAIi7QAM1boeVUGq7fygaxISoNnsCsXKzKKer1
Dg1jwm018HkXVd6HWh64Oy0KJO6d3HOtCqEg98GcCpFbZzXHJg/0yqpz8NJV
STZx1RtBpORqZAtnnhVqdbnkkWX9UJ0cboCSVD0btCp1njUfxm8esJsdaMjC
+2op+5+IUQs869NiCRlLi/Rq5sQkM7nj5xMnxPZRU0ZB069HF9ZDrN0yiwJE
C8j6ajCHm4SsgnttCrGhccyKDMkDb3SfmIPQHkyk2+XUcsWVbOBNGryeZPA4
t7RGNzs1q20FhCRwcM7BzhR9NzMvU4LHzVAlFXq6w4lDcLEtUFGKO5LUROJH
eRtgLctOgJ3/a2TJbzav8ydcjs0fHTSnPFyF8b5yX7MUfxJRtAx4VWiz9U5O
4YPRyRNhkhw5HWwWJxkh+L9RtxM8uUFB90Ed17EBdfObCRo6RMogqVhBvVZw
TrQQavnUSVfKtZtV+F136jqG2i8nvcmYWmsIBCpfYzJaX56/cC1d6bKMHFMR
KL6cmBnRhW0R7XjFV6OEkKnJ0NSVbvNWZbx6TiewsI84N+Lw/1nre2i56yG0
vrb7NL+McJtQhp5ONt/P9WwwzX0wV2/aQ/4rMPZbdO4kNb+OkfGfUj2Yd5Vy
49HEZrvp+C79lyo+hoA/fVum57Mu/UNDdU1YpycLoIxhmORytIcLmTbtqFgF
1akDljrcz+W1Ou/GDmp/9p5gcxXJOd6WMR/4+3c3RKF7mfdIGirLl/XntkEv
G8FlPW+lp950CePpBvLaGwVqmLkB3K4IcpkiUJSHxhNOOsZZ94eDhhr6SUUq
2/IskXvHTAhxgg95h3UVe5Yj5lSlk25a2eNcHRDOC3TDfYnyW1KH6cYIBMDz
NiOwmjo/HpKZW7i442aN8AuJRzUSEgKodxPtZp+UE7VeTphpY7q+DGYe1cL9
aTl1mRLEK5t7i9zeloqXcrscEn3n5rNpkomC3QYa67kITy+OEKa3ynNfvbkB
0QfHIdiPullCDRaWs5IJih5ZTLEcMpypSBnkmOmH5D+5A9cTu5RXp2MSCFkS
vsuR+TUYyJTdbyvBbJV+nbsaSZrL98xFokxrXUqXRu24yNE3syP4u9o4LZV5
ga9ZFbHeytt31m/qhtA9/ZhGcy7ssK1BcQIhR7cXoTgj2vlciZocs5hhHHeW
wCj8y5ts7BUOkRyvL1h/TiEeKCzv+BiIDrHfyhKvysK75CG1AOW9zCZJ41UU
gLCt26B4hFHAyxAUZjqNU+qLFXNafeRhTcSftphqS9o0Zx6PY2lBqXGSW+iB
xfqqy9ruZu0uHv8OCVeM8V8ny8FNrirMr4C0MWpKNsi7FF2N8vkX5YYvxscY
4f3zyE+Kd1TeYiSzHwoNOL4oF/BqSJMB+UaNip2tfWufI2xa0T1wh1C6sg1o
Gv3ViFW23WN0+dIUHSRFKm+9UvlJEHDN1t2ZKbMOc0lyjC6bscemAleSibo8
CUJBs6GwoMmzC4vPoNqUY0ioL0yIuJB5GKErOwaXwwECp8hIFU2vj7b0T+Oq
0STThVnq6iRnsqgeRoInJm+L5hBuapLn9QK/vVdGCndu8DwOceFwy1HDX3hA
Wmt8zd5hrtgbp2eanqbZCMGNO0kEcfl5tLONIrxXeXFxhqv2H4GrbkVQW2GL
+APmI8qnVZBt4EsCrQQu1XmvfRsVKoPG9iKxQzQW/QG5OFp8tuW714SNYpBb
+I8T5fgFex8eZqoI2T+qEjx0IE62XnzKwJvD/RRkKK3XbQLw8szCRZoRRKFs
njtbIAApZvq2Rs4pLkg+EI3mMys/4JI8o0sywszoua1F4JZVDwkXWYjiZd1M
Jxb6ULyvo6dE3VIMZOsBbyMrIPS7X6da6b760b3wtNgk0HzD7MSNCBWuA0k2
PB8JiR9dna5ugKl46pRPp0TG8VyMOT4dpe1djbAx2vMtzltnMYe0i8cz1sHr
zIDoiINky6LDOnF7F/0QNFUrlgqPOYRohcmtwnAqr/jGG9sbFTUbWONUxXEU
xkOmT1b4WEnOZQNABIHBzzYYk9b1TazD4oHt+JyrJ+rdyYnR+iNYB/RHIxy0
EQfkVrA9qv08GR8W8gp+V41zJfuGsl49t4SihydxVetI1SvnG3UNR5l8/B5G
qEASHu6gOPRXb+FqPHPNo+awo30CfEUaeRvaAh6nfcTZYGnNN/f7i7fsyPOs
s+ZEr+KXj1qaUHJ5mqjhHGUuW/DuukGq2Kn6MiFxgvakIB+peqS3IDZUFnjC
xcNCR6aJLVEuhWBVq4I8HSPfFnW8cxHjykoy/eq/RV+JSxAyic2ogyOQR5Dn
AviPDODOX3itko8MDsOaJ9NYDJ7jnniI5PHZ+/Sw8WEcMfQV2PRoKUH/PVfk
hZtE8q83ovFfIs0wEgZpA6tu+TTASbhTVHCV2vXqbDdnW8AZTkf8ZNM8Bd2G
JfPaSirxC6IW2auNoGFs7Pl0HG8cu6nPQfM6kdq6kEKNZtcUVkur4nsyYM0+
CTtFMh4p69+Rcdkohx8eeTyoQcxn1+WIWiStFSMgg8DndZZO+P1F3aMGr2ZI
xPBGq1F9OgLAF91lTU/tz+XABstLpwYLXssLQU+PBOTSb5uigZihxXLw1Hed
Gbv27XQUxMmsxbXZWz0+dk/weDbaTdG1hl+8Na/08ZOBOg3r10JBeZ/AM+qJ
nP53zKbnxgnGJ0YmC9nsuXlKMVul6kdUjpy9JmGJQ4N1NpsaKR8xJtzwbgkW
4ohJRXC5MvcYQEkLN0T4XsjIiyPLuD1h4DDcDzGE2EC4Y7BHDTO2U0CJewmY
MuUi/E/dRO+fxF+2JiS5S8sDcQKcOijRmtNZApuYtAikzYtAD8oo/S09rnUk
YaMvojPdWZHWQRg9HjT289VFB6TTrw6DBEOyU3wvxGzs0tsniNeoqJtfMHhM
2RDY4KTrRkDpPUmAVZBJhnBM6Y6o1OXeRnIZoVKlC1Owo2So8vi7k4pS2W4r
ykcUSV3ZIbzFc6/yULW9HVYpNC5k9Xp7syejsXXd32OfcsNnYzcX8iR6SIrZ
wg11I2t5bLxerxZtddv4GrK0HozaEn5yGB5JBkATuuulMtJr2a6nVqiI/5yH
7Nlw0EhKlXNgjBowrUq54SKIYH0Ojsvqnx+eS0ukPFGybSK/vxmiNIped/iq
kWS+p1zKJ+ZUlZ76vbMMAuViahV79d+2T6vtuzymN/gaFTpbsVwLePzeQfyn
QGzmOdtaUWejHviSuuj+/OqqJeR9mvwDvrnjC1Cogms3HuoSBbngl+BTZ1x6
+HFS19qm9EXKtj2wMeG8iBiT3RnkDMbpI5XlOH5Oc7RRS7H6lqKEkm18BjPX
U+3hdLPXoA5qeT4I3uO2jXf9galAM4xji2NpKG8Cl64sXCQB5epsQ57JnC/j
V7Tszt+zMgibcmWLA/eJ3bVhIm/We1X44iM0Hn7pPzzDLpCn54SiyEBtiggH
kFq0FLRk6wC1CyHE0HjF/ZgJjKdsXwCZ1IW+4WTmVs2972brP+1iVmbgTo5T
dTwUqFXsbniF+xUu3M8DEcx/NTPMG2uOtWOvLJYwnE5v4d62kaEOiIHoe7nV
29bo7uFgwPM2BA7nXzKpo2B+nAK3jKS8BwhNXY8K+HLsI/qLGCk1qyyFXhEP
EEohOUgPOi+eM3k80elj8SZmraP2raco2LylH6a9zToK5s4MzN6WT40uZOJ1
9zM31hMZDbgbOx1wIJ/RpQnqiMRY3SlMBfJ0THxXibAr5xIuAoX367Pb60Rr
O3rd0pXWXTq7mg2kLrWTOydVVYGtgDJeuwju7XXd1qiEo6s4wMY/Q1VdniL3
+5enSmG5z6cT5thhzId8m2yLgNLjPAJlaEvE6w4Ewvpl/uRejATXeul1BHjO
VPIAWMRXUVPpZhvkxfE87Hv4kYr+NmMmM+iobwvaKdpu90QlESl3sQdnygpB
2UdD6PUncgTcFDmQJEez+s4Q8SEpR6ROZMnTPptvsWBlrzPxzHIEmXo/YWsS
3O45p9dfbJaO50HJhOlloOw1HvsU0aCGNCT1pBDqr2HWxJRwj6BBPw8Taz4f
rHfxXR8NvYxygg2Di1i0TprVbPjaMO6beANk0VVKgSFiK2POewh0dlT4H2rC
oT0Ym64GD/iVKXMxdbGCmEaqdubiTSKFqdLjXge4QaVvNvZ/1JV0FroLQ+Ig
UtRioeQlp+p0z3xUWYEiEeA/mTFTdMFAE5AyFFgFKkA7Gwi2wglHWOHQmZMy
2OUMxKmMs7lpXA520Nxo2bSN3QvYs4Azm7A1Id0CduVe6aR56/Q3MI7t+zUY
l42JRinbIvsFAUd88TUpCKpvSgyuHoKAI/aZ05cWiCIDgr1bDA2sDZdJuEWl
yIk29NmRj2cu4lh96jivt/fI6VZZna4FzfvF/CS8Pwc7E7vY5r4WByQxUc2/
up2xFuoJ5fJA5BJd5Zy5j3v8HQ6up5Cg2GtlFE8BkTLxeq2NQcEM6E/Pv+XG
O/t9ShMxNU+wsH/CkrobUyN9B5jREp6Hlys9M8zuTFCx3iHZ0KlngoZEHjCe
nku9EKRUV4J3wSmkeWrOrYmPkLTUEeFm3lcyIJDWc2Ykngw8Q27HfBzT3k12
mksQP4BJiW/XP0OaDq0jhgFVEOpnm7sdzBs2fKcs24pOyXA6EmanawC3iGru
KV9GhzN57mEc2hNjYFSunbZLn2F2h3aveksp+D37SgeKKssos/bqwQWXd7ZN
loYLfz9LIl7b364dV+EbHYZOJgtzJrzFU7bp++J17P5unZ4SW06VjiXU89dW
nuTp0hex1cuGD+d0NyjR4DcSKtsfURNOgUcRFhvChk6Vf+0Au19p9/rc0bsJ
vs966duM7RB+RcCQv7jx2F/xxKWo2ns+bF6mrG+y7PsiQvfSeJvphBmCIyyT
5Y3HeAEYGplYJZzbKnQKGO2011qNugXXxQQaDOJpqslOHw+j6OWl1KmMXXqz
QgkvJd63XZwhwecXPyIVHm+Z/LKf36T+CHt10jq1imkYsMSBNJjjaDX9pOZ4
zvQaNTc5wKY6LVX3SsMszzHofE6qZ/Fp/9u5jJcpCdcTc1qDFIob0cqyuMNh
sOAi3GWQ/usbAmzmJGicAoqgxkG8Y+XoqCBWoibI7AyuSJqcFNdKqNSAnT6g
uEPv6GsCnpxvQ4IWJWyPDgPcj0+5192d0y8VkWaDmbMd5c0UNHKXp7chSwgR
ANDuySVK2YYZ0O8tKCQC3YtlvVrG6T2H9DdJ6/bZMm/NmsC2NZBeogR2uLuj
Zv2HD0Et87Dv0fdIYURaSz67Ozo7BeUU1zgmam7JJwUo0W0ZoFa+QqcO0JJ3
dB1rbHFdTlsH/KMnl2CU8Bw7cvRXyCwB7+z9JfosusERD12Hq7iJcQeR6Rpp
AS+QC+2DFLoGXce3jSkyTew8ITnA5uxpEnzC2CBNf3YXxghFOSuoejzsxGqy
fWxuM/mvpaE0QJOfJ74ailAhiMRoQenPEdqExFewyyePKUP/Zt2PqoIuQG+O
y2SiJDfnaRORPhjBoNojTpXMpLGHOB2M64TODTMMpWj2Gd3aJCYeJmIHR8Jw
RWlxd2weHTlnBa7hx0bzUtmxRg2jLi4m2xV6RwhUFTapY6f9HsN39/wGafam
+crACIXStV3o3HMSMSLqcgdP2LKxu+Fm7fVlXanwnsNzN/Sokk+YLmwEJ69K
oHGFEMYZWsoHvzAIQclJzdvouFxtaKmsSWZVGZ8ghqn+n7Hz72Wzrmzbrf1U
2Cg3bK4sJvWv9Yb4WJkqp7d3A4P8IWzukv1DqC9FD9XvvfG4R6lGvvI/La0g
XHBsgWGHsFcfj+BFgVNZ4IMvYih4Oox0pk/Pc/YkIzGLsLWUxoDY2H8pQysU
KIN7Nyx41bk+0WJQFwZJS3SwmCQeLnx5IhjpOn45GrfUZttFH/VsZHAJl1ue
Y2ns5qx2fQShJwggwOi5yn8KpDCc7selhaaXQBlbJP1weofjUlP5qJ6NpOSc
H6/h3D+7VPGAZueJ9FQjMelUiZDBXQue0lp4zcrBbTl3ZgcQsP/tdHXun7BV
DMFFVu+hbR6EpTs5+H1n86IvyT1kRzciXCXUCu6mBZ7a7UoTVbTYZer/2Zp2
nP/T083EZGwezgMIi/Px6CUt/gzYMzhs45azGLOZQdA3ReizddbOIgGCCT6O
o6JW+pPouRAcedcSseDwv4e6M8+l352oc2+zWLFXnMJ0UqyuKvTJrqNQwIAS
yLi16LiQ1QlFkIAwM3FkpG1AfPLSHsl5VTiK6NtTqr9Ht5OKIzPSJji9QWa8
rcCUaAOULP/ywVlth2iywHjRDvUZKP5yBpwryfWaJaHBXR+HMwrFw8VigtRb
Bk409bLdcfvFJqmzIzBPXYms03+ePvwu24pUXgow8RP6DIfeH+9usdC4y72E
sMqPrTMDEwc21L/QOqXNn6PafbFK/zXKxb8hzUZi5JvQzn09s8q0hzyyZDxZ
TqjQ/Umk1B1IPre/dsYIzlGbU9QjNrFc6oD2teq22w++r4XeFZtlySODgc7D
anShdzkL0ZGXscwbXbIUJcruFkKKmI+An3btyrfIREqRp4gRwbJBw+szlw5Z
OYEUCWVAukzAqSUuZospOAVF8zotOXIkRELzrOLGiwhkf9IrMjCEfsjyIVLg
zdC4m+6idxGVoPofF5rQb45o2J1TIzRrTx+XQ0I1ztVXvBq4gniS13W3oa/U
nSO2Ww4hugujnnGJ3SY0t8cyKQYgKuHQp7BoeCBTMjJqmcGNgFHI+qHUHn/+
nxiBIcVCfuHIpQu8JXyp0rKyBqOAhr0jakOasivh1L0PYhonoDsmdFXhBd0G
IRpNlyy/2dZHSFVY1Vc77YPtsDSLlDXKUBGjpEwbCNujKXy2l87Q0SJSeKH2
u16ZVYivVZRbDAN0ZtQm1vV0xLHXV2mcJZauKq752ujRFCpZePABfk+Ecc1k
v7DbBYpXwwZn2Db63PAy8hfvSNtK84tVUXh3xOgL4p37pg72YVZzsisNTRRc
Gx7Xn3iDnRqEiQOf5r/333pX1XSRmqHZ8wnJ7U2Sex1LvaR9fQz1aI1gUS9+
/eIPWttny2H6tNAkGQv6G90VkSTzMJVTb3Me+30+rV/uHEfPf5dzJIttTiIk
7/r2TAiAnrxHbWs19ydqVtFhJCe2s3xlUY2Fwq5lnwTwFQyAAtxrtGYgGV/I
4zD3y6WW6kVEaalAve4w3nUrvnaY5OBAKk9v6eQKzPitDrfPrH+oPg4mP4RM
SUjevmQVkdzICYBOxirCn1E+k58S6q4S7xiRCeK9qrvNmvraLizltHNbF0xO
UuFzOJStlkAfE2Ogr8QaeXwZgfzFx/AYuRXpKrWckWURUBK5a+BvA9HQjsoG
69osFF47KdfHu0xkAc2R5WyOssgsuVez/EVU1CaJgR0f1o3eLu/kxqT2FutM
cP8AJXk5IVFAZqg3xjgnrVEhR9jtMR4li0/qO7awxkwirMLuTvUtX1zFAY6u
YqjOa2z0f8oznNUoE6wnMLPwA9wzJOEjOKcgAA2wVUL+u3cNFAvU0YYGveK8
1QBSoXX/TSmcNBRmPPyQw1ZchCbz3y7AhEc3HhC1/bCefRJV30lC6UDIHdOe
83j57ALy2M6g99LJmhFVHfjmo2veEBMUZOHo10bkotilY0VM/pZAcQ78UI3c
YauMkL2TLskqXWKEbEQqCjGKwqYnsloQr6QrZkFwtOVXUd0G5L+vOecLLV85
BAf9JF1HluP/kc2IFFUcu6Jodjee91BGGb1h/dtIN5kZw0h1iGzB0yDsCdWL
tI1tmnXo62BcY6yLhg3GeY6V6C6A0TcKL90d2cl7KBlavm5ctdL47QsGKyn3
mKWw7pI+tUseok8dxsMaA5AKCpHKH/VcqdtL1pWbeOeqYhBV3lOO91/brN5F
OszbaRgNl8QFdnyoUZeRy/RO/4qHggFpD76ZfS6ZU6/4RX3jel9AMPJHUqkn
PQefWPswLBgtJ9XzVYrNHugUTx47OcM2D1OmXiycrUoRLXYTxUsZkQGtNgsq
1dU6BuriGR3iIr94ZCBIR4l2o2Kj0B85h1HVaf65vayHcJlGFH05pngXyQ0U
NZp/R3VZB/F4V8+pF+Cxy7lhUNcuXH8fIBw+O9g91RT5p+f5VpajkPupYwC/
8ooMvlA/DzCbUkFNjr4tiRN/G/MpNEcvYveCxsRhn+DDFW7anoTLLVeb8q8D
0fYrojE+eXR9vYorGuzvKN8CZUSJ3H/no8/zFyX6IMw7CcWD44KhH8omQ/5H
gGauUr+EmYj/xt+J2xJxuWbkGGGi5vTxftNyrX68mWYaO/niruUJGrSUnPIz
mWoEGSlQj6WJcjxG4kytmmc8dHGAwhwfrTo7KrHE64BBwjDY5S3a6sJpDyyF
aB8qJvRzWoo/rpYw40lzlFlQo37B6eyXQq1CPEYbp4znuUv+DfZqzWDJFid6
FzLBmDwwhcrL4tIQ8z+FRANG8l07fQ+euMPPywu7oq57V4pelabx5/kwk46y
vHXK/CM7UezSvvUQDHQt+iajvFF9tJEPvnqlIb+jMLr1htJyL5hM1Jf2chCd
YK7uZ5Fe+vajxtB/SmL2CHlz0x11qQfuyj7f2gdwI4QKIMWBd2bfjphy8X4g
uG0M8jQUpKnqr6lNatrcNDdcwluYU9VZ42tkt/5/0K9Jtj2YGQByMpz2E524
Ed5Wvr+tjnZV75Buy65/p7+D87ta0v5WSE8QXzJmvY/cGM/oMBYimE3M94Rt
yLFfdQHkYthMr9yTbgHgxezerd23mhqv5VWRsWsvTvYLICLkRt4+Cttk31kU
Ux95EUZTCWerKRLtv7p7NwYmBqFZYn0+JQKNo67Tr2EkyImm43T29n9cTnIT
74QM7u5UAmSc125981eNgntG3cxqIoKoprOkMEHDoyYP95Qxb0zVKOgB4aYW
7yUBxr2UH2vIr0YEKv3Kmcxqir8JrJeOLdo1f1q4V+Rg9Hx5QL/8gyG1cijZ
oiNRXcMDGMj6wQNXVhiAwHZxxzoWmoBac0xtDJuJC6P0MmrCVcbrTHtMY3hH
N2BHwk2Ks3RMg8h+4G90+Z995BdQfiFOO+Pqy0VeJl6muPKmCeMAaMlsigDg
hnoxioUtUV4NmL+3BTv4TsLHxphUNDfvE8iT7MnLjNdCwds8V6Xvz4e5HKX4
EGEFr6SbMUTzPB9MdjHg/qHfKdKavSbUUqQ2IFww1nQTaEda4WUSBfXObSZb
D7qpFlLqHIfhRVIv2D+eJl2Ch89qshtlt+NHasbXkwOw5IIxENwot9pdVm+I
GRbcFXEa7iDgDWEkY4vFGv3Q5KEYaN/ryxusTQppOFEXzc4bvw9UNb4tojOq
f0e6U4ndqwZQi0RI57U/xfj8m+pzbpmU23uGdVSmd7qicQtXrw0DLz/XaYVm
uSI3FWKjhdIK+l859yzUdsT3+Wcnr9xyRdGTYh9q2Q6lko4gXRYZZjIAvj0Q
cIycSxIwVLPMbq3zktEsUH5LO17tbziTfuyqseW6g4Axx5UQFOi4FAJmSZ7p
MoEtSuS2nqb8oNLR1/9oQrsfStTAK3/yghBPbVJn6YBF2XKPDR5urnpTEbzy
XpRRcN3VcJLHnSshGy9NQCAg+JnsoxLFMzpYET8VrTeluCBjvBP7x9EkX0vW
1c6NtcaMmU3EwUAeR4Tuj/zbvPSMmt2UPRi8f2N0kUv0jCm3nl34dTLqR7lW
cz9/UXmCkuK7/eGYdn6Q7urKwo7ycOFbjTOvrlsIRh5FIXRDKBdUMJRcZ/qo
LqjK69pdQYIaSjFHnPNviu6zLPlAiFYWZsLvNW1B2aUUnxLZhnbG6ixGA7oA
qQMm/58/h8iWVBhcsuv5qxX18zlAqKwi5u6RPZn/O4z0oEi3EVVB/E4lnAS/
ZNstWQISyukLoEqX2/EkP/dkbsbecblhdd1D7ctpffb2HyF8PDz8T2ZBuBTh
77OiD/G5428QBVlK1Yh9RSB6E+XgH265tqnUcD8Dr9bz00H38X77/6lng1qn
fVsSj1muk7jDxZVSCXRfQm+qWKMeTlcdVKVdQM/UywpX4ox4Z4QVAt/9HFBd
bl3jBnD41JOtFduiHdR30M2vrClQuv2K3F2NRfU2lDUjmWIXaUrt7ftKyG+I
94BuTrxOKjh7RppaWG1IUr8gtWhsDx5Rad7tPi5U6ZVAwumcRqV8wBG7RHkF
V3drnwNMF9pA/LH4lIyDfK93p0p07ZTu0zzP1Wgh0YUbzfOFa+f7BmgUXMrm
p3xIIUmsqTIgT4aicoKiqHRpXGrpV1QhIfDTFuf5CuIGaMZ0FZ9S49oYaH2G
brHVAHDwNf6DOlSITuOsNHZPyPTVDSmbHPK+EigtB0BWjwi2WOdLGfOkCq/Y
2h0gNHPMn/YzbfibhppBWMRvLzYHZjt5BUXmtKhn1db+AHjeu923CSA1+a8t
YmsFIjqFqGWakJeLUH30Gj1tNR7XaBloRlUElGwTiRIcYOpfYahql2ffS/IY
3Am8lY2kzU+EgTxMZSqM4+/kNYaTuD2SfEZT5IhOQMsygGF0/zYyUEp+HCCQ
R1dID3tbqoAV9xzks7YpkpxK/bk6R8dQZzOXssfqEXIK2T8yeXI3Mwh11qdu
lk/zBqK1hWRRqmz4v+5exX2sb5KsMl7f0Lem5AUU9511h4a8qRP9wcdTGVdL
KwSh8sscQLYd8p4a8HXB4mar/9hfGOAiyf9Ws4uUXff7LFC+F7LuFH26o6ih
rTIQhu99fcyoYvAjVRzJIZ6c1p467fqQhaZCqzA6qzju5LDIdh+plo0RxbDk
ErtVbzS5jVkL2+DQ4K9TmoaNdJ2JHhWcBkPp1OAEYG+NgI0LvCybtEtiEhR/
ZYZl6W03QBnYBUIQHIf9SQx3j6pYNBGNr9lAtAk8VgSoAIqRS/cXDlqp1yRK
Nd9sq0lf94SJ0mlv9OeQ630x/eghOC2Br2Xe/qvbLook/ExT1ZhBvzBk826D
w4Mob7lYmV/vDc4Da0dcIHaAkCvo0gAFILfzuXc4Z8zt3XAzOOBz6KR1XfsL
wfQ6+x2P88WBdSWgHX7X83Mqb7pApBXTcMu372O7ZXa6pWBqroOh3Zn+T1Zj
Zhk3Iw8plGTCIAVQ8DANCKwbcsOKTrZTIXTesXRlaXmbKZzTNWl+21dMgmuF
DyL4WcGKb+MSgzkdZfi/IFYBB7Rym/tK5bBaBwvccFCQFaGtSvGq4yK3qrN/
RDj/gTv0Wct6JoRg3rcb2Xn/AKa6igUSFwWOy+Fjaw3txYGQNOn9NaKxa8yG
ZMsCCH8RU9yoQ1qfinOtPWxozltT5RGNcfZaP2WyanJMyU/xW/jR1as0y5DC
mJ/LBlWRo/Z1LylHa0tXWCgA7Wd0uByQf9n3LeQR4ricuqA7gQqbLq0qB5H7
tg7yzetcAv/xmfjK9XTwYvTZlmT0ltXuH3gGUUl11QXmDjPo2UeVBYC172jI
0fGFV7jV5Ngy3JrLBF6Y1sABOugFUZWj1CP93HI2s2tVjnggJIRNvIA93Tw2
0pZ2uZNqsOWafXbUFJ0yFOxOFv4wW3QZIcMH/TKUMyQ7X6iuhJTqQvRKRN6c
6gowJrztKwHGc2pEy77ipaE42cuElNdzuXJ3fGVITrmzntZ3KMpuyaK5gZtk
byIdcYCIq9XpcL2lKPy/QS+i/VF9Ibw287o8S2tPUQNnmWNIfeU8c2GHydZb
B3IxgsN5qnkBxc/k9BmBYtvyqI8OwXMXbkW5szFSFyRtOgvEhso64e44ufF6
9/F+smrwe8VRmVyTWTV8MiooSOx0Jqixvi1p4Nf6q+JDy2Xi+Cy1KnjbhRPj
PxoCe3GHr3kuhLmcTXLPYTsZWoXLpaw8D05T9/OPjlIPb2NQhNk8N7hTPaPh
Rc4ScIBZ+40H96X7n3jmLFbexSdHjtEvN6zgyT5UPuM3L197B1ZkvrgcKTWs
CxoP/HCGsZmQW3QaNFXAS5FlniKsyU6KjwtP/bBeyU2vOgTQ7TC2+IlsUcgK
8KCcEkdpaIaBLP96xdAPN+qRPgVXkGF9dACcMEjDIYNbWvzVeXAfMAXDPMh6
o3HkorvFwaGfCvSrZWyvvi3eV5tG+TpxvUPdboJVjNLKnwjvhHaHJirmOVXu
4iSlQxi3Nz1ydy0by3ObzTUL7VRTmtA1dfEK+VS8/+YBBcGcIZaacW77keZo
1BctV55rQXN4D1jb/qQ536mhcbGY3MFZYNLFpEwy1yaB3MqymwPhFDfsAyEH
JhdcGqLjXckar589IUb9p9Wwt50llqedk/UFiboEHsf8CV2NDgXP/uZvJA40
Z9BPOPcxeAOG16Pj3YjY83PtGUiN+GBFBwKK9IU2QZ0EiPbY9NLUHaQIIBLB
Bgn/tRazFs3U8/LQSeepN1QCEjOfIVdsWU8cH3jB9v1PGwI3wMcNj+oVcDWr
pFltK0NA8hqx+zTdoZyce+6ZV15G/y0I4UZeAqvb4bicDOn+QGyWYP3X30OC
bRF0ymkYcxE2iwwDggIo9nnn6TnSKBywLoCNYr1s1c5mxjZbjKAxvXNd9ORs
o7tHinbG42AysriysfiMPEtCEmQ0jrzrbBQsK4ynmVG44uGoRmrRkaSsWV7z
WfTcDggisQMLvux7uB5JxH9XOmt48VSPkOk/nYT+Ixoj29CAAbpzNGpyt6Vd
imZ25MLt5Y1VMEhMShM271sKncBH/1Nm4nKC75+RH7/0L4zMHhKs4g/S5VMA
72LHBc6P9BS0OiAOgF6MKHruYrEelf7j0lJyzhr78py/7W7YRhIXByr2UewC
PcbEiKUQBsbbz7XyFGSW81EhHzzfvu3rxiw2ZeSTGae9de5XK32yn11UxMsO
GGS6jSQap9z558cwB/OVwz4JHriZCWU4toHmeZ/z2iYsncrymVoT/gAuuemS
TT5+PsUKGk0UrDvHzJBKldI8NrRI/qZrgce47pPTrW6y81HavFvo9vUu+fke
/JM1gZplmCNYMT7//4v1zOpT1c/IiWKdMdE2gu9soFIp/PeaLwmjrpaMRoHI
tYY3r3ECEODFBlZkL1T8hU9m9O2SFBZNxN4eMjGNWURt4Y2aAcoLcLHhCTX+
uqxbvkgP8bW3bHF1KJ6v5On4uXfnUNZqtodEwf1DJE6EKQi5zYjO8YegLwwe
50tGCvBzoBuwxLvhDbePX3kt+Tx2d03Zpo1RpCn2cIP8XSBgw4N3CNXlDTLJ
tXyUPP4geIUuNtWlvORdHE1jhCuWbgsewhzuJhQCJD8SrAkKnCm21MmFA1b7
XyrOSue32xUk58ekNztAM7CZvun9HHDZR/JIbKKFGnRtHdw0sijiMpgzzBr/
P483pfELkt+SifodwClOtKz+eXDtmBbvlaFT2ZCKH3ugDhavNRPpz4UGseyM
WJPGwr8oioNb/ucJEuZ2pXrgFfsFV2+TewrkiNZubLxuNul+tIpTlQeUFEt0
xlzOKP5mXq/7Ftponx2rMA1Toor9D2Vx/JPsWDx3ddmukVA+kjPJN5dDHF1f
zqxZHmsZJ45XHVlEIgQ4/qPh/KUNflXEwY8Zl4oWOYHBxQv9ZdFAMQE6kfue
+X94LmU79nuRJN/9BrYK6s/AJ5QYpFyz3ubCD5+4yvlKUM1Whaf5XhJoxelG
Se5jm6dolbT1mLQGKeoNnpHtFIPdptv1Ya6sC68Zaq19yrA6tqsZ/4OYyfxW
TzDOOB4Vpxk/f8KLPwN86EEdWK5e2/oEUdSqOE6saLgaUd/l2sLcM+PM3P//
WCXM0mK1U9/QG4zdXStpkvENprP6oQkLtMU9cNeCr/kcrlIoVZ0j5XHKrPbo
StlZKqsNcyDlwsmHkGuxzqKm5OW97gS7d4RNha4Ngahc9I1IjWn6jnu5d/Uo
59hka2/KrkfEt546qII2dHEOBNGmqhukHWmoNwHYTvbkIr17wRyM1IjEOh5w
y9qY4i2jzvTgdNhEuNPLx1afCek71EjUJ764pgp7vu/LRJFngAfgzPkRiTGB
aOlqPB9vcLQ8rIpKBthRmo5RpXGcVlwEeolH2v1vgadM6P8JgqM3AveZJ+9N
oTcUHlnHcjEkv3uXcbtq17mt2YvkGoWJzwkdFuHlHGx1RQzRID9wTz0Bm/te
2q/yLlC2ThA21qz1w8Wsn0HBpeQVYd5iQTwHrYzyu1ytXbu4oe6kbMB9CZoB
aid41rk6aLtk69rkFTAiWJ4vphX8shuLSxzPM/4+M30d26DE70rL4yH7JfGi
AvhnVj9gt69/mOrSMW8l604el+sg2ZpvkljdjG+XGoUOQ1QluIKAUlVetqaj
d+ylkW+nvxmdnVknFiLlO3erFNd4zm+fWHna5D4mHH5jVUcODUj/anpG2Btp
Lw2z/ZAopYBzreHZ9Wa1GPgy8Xwinv10+ia+5gOcZti3qQ8jAcWCdgWbFBBY
32jtPtBtAnjY2WANyG/B1ImehDFGXlpTQoGM5ZNIEgIMKlwQneqe431+TJsS
38IpxsMhRLw3XbulJc6oLjOxUM0Rn5zW5jfFgHp2Uq+PebWney/Q/AC9lwhi
ql5V/6PpelD16r3AivTxn5Tx/Xf+/82eeuO64BV6p3ZlwlFQn1rKXdr/WYJW
NFgxykuxD6IHsAWEqNgCakoEkh4GDRVhIc34UBE6OXpU9fD32efq1k/xfiu2
mkZQRu4oKkuktC97EDoCwbqRpLGpa5t15oAGS2GMo5s46VuPyzfXMOJJp/ZJ
SxzrUZLanVsEN3kRTuP0blL16EUN6FZTotd7MdWTMkdvl/FX98m2r8/6nK9G
VSwe8Bt4ri29lGVG40hUSjXZe2WdWh3TPRuGlROXsF0H4R03lDvFYT6e0QPb
UJbh/4xej1StTvEXYNJ2JDeSXI1Tl/LQrvTkTZlFRgYSB9p7gMcUC+X4+SWc
lI/NhHRl1wW7jneG0D94DJAhNq/CsHpQdb7SXKIWaFqHwdwecFg/ADobO2/z
CSP5PNpjZPjdvZ5nvaSOrSjX82LEomeBc5RRuAdiQERtv0Kulh0aTOftplKo
VxxrdLYN3CPJ9kPTHj8xI9Wf6rQqsm/O1uT0fNyn6VbmREq25yfJwuNCRCDS
iy1q5V4UC7ju3kQvqRVnTSHx0MjeGn6AUgOflfkVHaCeupQ6M20JLFShpXwo
h48L9AadxsO/znmTw4PbrYjcM+zk9JLYBeV7heBXn84CUzoVhpYwr3hQkwhd
bh5/Ixl30edzCfDrsGHDncgktjtllsHyoqouQhjDbJwhpRK3YK5ieiCmTGFP
xXYAa9MuXmlkU+mEDl6cXuUQunHRtiTyvNYEg1//0MjMJEp+mO8aEJMk15LO
JWt1hbOqg6jFJQm2VCeGA/w72OKtWR360fKLIT5WciFgW6Jv5ZBXZ3vbli9s
ri7eKU96NZoSXNavNUfzVIPUx90BUTVwRG2//BYFr9GVNLauuBCzzR3/Cgka
u9tKsuscfrBmE2TN8456CObv3/qY37Bl9/8fryT+PuSAxvpB17wRE0ZXX/C6
HxBQUFiujqC29xXj2Q5qGEFGwQAcbRQrRc7UBeL6P3SzyC8ezRGCpoHs1kIF
AwPSuwvzDDBygxy91IllzfHR8cagXqRvIz8lHOw44oQODduj6DL+ZvPkTklB
pBGo7T6aEzwL9+0U9ZmkXWtQopw+IKTfKei4C7Ms+Q5DXlvY6gZ9lP9TNUW3
8hD680rnh5pugLkYxVTIZU4sakTju35o1qChST96WAAocZjId4yELmJO74pz
olULLMXQnIP6jAYjeHnJ8Xd8JlaXsmi7Q4J3nKlUI5frH94At5VFgv7+hfXV
nk8nYlb8sxeH5XHY3FWHrToMPep9W23xKP7jhYl2rhOciS+zS6nXWuEmnSUc
ucAqeqSFb8iYArDYVtBf8F1t9T4cfZLvIFYSYnxrRvQTmKiYPKXISAsmHVCh
0bki2EkXmDVzXlx1ZXP1ygPUX9rvT642orHsKmTok2JNIg0SITHj9Z9TGxvk
ABXtOUtoP1iiPSbMKdB+TbnUPlznd2lbvsdmjQ1ip7oyqw8Rm0zyuj5Jei9h
h3Q6fhWp/GFXYmFatfMaleWMc0f4zw8slL3nqpl8nTIIiZGiJs7S43so/Ddz
dwcUWbjWMKiHhNEHt7Qq64ulOFi8ILcYKzu9V9GgTAbr83Q89ich1PEAwiZ7
oMluWCIfUK5X94v+e6Dosl6L9W/BpC6dgZ2oew+EI9qJk6X0KFv+zj/4+zDX
82dhafHD6psqScgLhrCW237Q6fyZTN65t62XjXT3UsQYrignMYmxj1qN2zMW
vLGnTmbXSbAIw4emtzhkpOgqURMbxYRxszpWWwUB0g1SrJ1gF+BMMtJpo970
qZyfOdfMjQiIBvy1djNGhmxOZnjNnzc1asz2cJcTc39qfEegV8hUbhQTqIU/
aVao6/gWmHuLyynzGCQQ2lf3z57dOhtYmkcblfw8mp4E/am/xnvNsEEkS+yS
TUoMLf3kfNANjpbFZ4bm/sDdr5DHgi5B1iY7hc4Agt3UY5BeU2wq7Ixmoc8Z
RxI1qNZXY9pfoXMAX+bU2e4PpB+OHbZ6ApwlQxkR0IUDyn3hScIPOfB5W9xy
ZHOzzEJPWZb9qqIWTOtWf10g+3963s6PyNv+yrBoCATFvfKLyQxmWsLfXETR
SRmv1Qm4fnE+gYbeymk2Bfw2I+cqYW4UHDJ9KJDpmUoibJkIx5vO6zlm4CYd
waqU7yafqqpKi55hKD/dSZpmGA2esI4WLlEfhW9npZG1ztdUfO7gQh8aaNdy
SPiCYnifIxLuGg1clkS+EbI4UnEpWp+5yqlmf+dou/XFpjfuNvJFYzBe3/QB
LmmwxoKkcdlAX0CjKDFY0615s6A4XUCRO+KYJZMvbcwpeUj3OjzOSsCeGKnS
H/UqEQrWMQXKGoze4ygcICItqTO494bDY0XUs2zAtGwZTZlNKqMd3HPEtSG7
BIUqCn53xOqXqWmiPTL2wp6I9DWx7yt1EhV9UaXHCDxPnV4AyHDcioZ5pU3q
YgLshTsAukF+pmOTUUw3hc5DBdsZRv9Xx0I2TZSarpOUGtSoPJ2NBa79Ll0N
4IpO1M0OgHwNGI5fQpVsFdH9qP2mWWKEWFSXySH4gmDpUJaq+aaLdmngbk+1
CcV4e9+tbC92ML5CHXc93UGwHvAS50vHBe8V+gPi/2S/y37UIQmSAe1Kylfm
/8DxuEcZE2XFxXQf46RWxb33FuOW5U0XnGDhYHi9zOaFZ+3MBdzKxtyaJ3y3
R7aJeQl9R89mGk9krjvLYjTA16c2zXtC+a/ytvxoIpKsYfmAPdy6c70jsYiR
L73o2iTCJDDGH5D53TjOAez8HC10Jpkwo6L7RK885m4oyBHfC8ZL9uChnAJ8
hd+V+pRo3g+2W4kjMfOlotDmOa3DoZfEEBiYwvtCi3j9iOFcI6H60TPMUjdI
729v7ax3hOkivFUKoZDNIVTzAxJwUGg1Jbe+jWpCkVuf/Pq6lz+gPBEZRWYn
MtWqNYHNY4uPLqC1OPJk2q1svX/VrDPfwV/FOnF57lY2y8DV5TGiEfugn2oM
pzlO8oxw1jRxcKvJ1sxDBQRIdRBkJAd6jTpSy+SKrOT3OWa+QW0wDgH3+N3Z
f3lVRenAKFQ1wwfMS3An2aCQsEnUopmfcsCPDsdsN/Km1IJrMsDXE8NtJGT2
wv0qF8RJ4Z9a3EtgwXSWw5cfhWLzSFUM9HXm7HvIMBkRQx2GRMu4EgLQ0G+1
FoSbQafGvT6EoztXUMJVg0TGuJyn5FfwmYrgaSQtM2m8TedDdXeouCaYdV8w
ydrzSjyHMVUm5xOONv4EZoZK20pFxSGzgfaj2mH0RcrO2kh86531uyMiVIon
lG+ZxumRClmeCnqusmyP7KKYSPyP60JYZ32mYxJyrGhG3ZQ7RuEoQ2IhYrS2
cdsQUNRtn6MMyiSHZK08Kva6wPp1hau7oZ7V96vP9fHiJCq3GD5XJSZXhzjL
XLY+72l4JObCekYJXSwMTI65BSk2xIxxnn7UVOuljOBbYaeElFeq3UsB/OME
GnrDhVt0mn1Wv+B7lShiUfvjyXOEA/63CRU2laUY8gafMUxAtbpDVHjnW5aS
uIJC3j8mXbb/eNb0KaAwpx619OnxpMS5D8EowMmt7vZHcoHjEM/rJuTZzQPt
HaSqJ97DnhT1Am8dFFcR/4vpyWmSKn+/Vz2kgsURiIgrhDbb8WKB5nzHE1iP
avPxMfMZAS7AP5ljWoAN77LduiEAxF+7b9Pwsw6UzoJYEdD+Wls2Y7j4kQS5
EW+6BZBYAMFTYJMK0DHrqWRoaSBgZAMxfp7sbgSzRrKXaFYa7Z3zfW9mdDez
nZkHpESGCmR9tPY1M7KHzHadXwWptPOSpTqUlQxjXKlv4UPjw+2+eO6RBYKJ
kEtFvb5TyILejxfA1d53skqqs/Je1/7lk25gz9ksR6TKnHH7T6M2eb12wBFA
cctxrJ7E+cmcADReKYoNJvPDer1A/2y+RNOao54jQ5uln6KFXPztmnsTaIzg
UfBE02AVEytmxFSnXiUqsLLcRz9nsW/48KzbRh45Y+AyM01bSU55+A3b28Xc
5sY57Xj/tGyysOirilUoe1biKB+MUkKxTqNbUpm0zHL62j0An1Z+xn+Xq1Ec
Sppgt3RD5Ks59eSy3bkSzpd0nIA0ydF6tTm4AIu7eXp41DuS9oqrBA/8aB+H
J0oBbSSrCKPPQkh3iL8lcxMHesTDwWxag+u1Ijf8iopA4hppMeo67+uERbso
C0H8coTTAabs5DvWskDMdjWRFxx5YWqa80eHgVGktiWzQzBcHg2DHh6U1EMa
skU7C4B5QSXYEYGmO+qRS74Q1SDt43fu1nGZi3FlIgo//ayPqD+D6WL26ANJ
VFV2i7TZ7n48zlqhH4gp6BHQ7eiv/hhOBFXn2kGAVFM9Ka5O/fhc/gbhdKbe
5QFhXrCGOM246OF6BE/ru/FS3iD3FeSOAXWsleuNjjVmzmcwCDtyUELEWH3v
Ic6fUtcmaNrwyi29Ljj1kCq3Lci2DPTxZPcITMh2NZXygvChwVKMsEDqOuGP
ZugnS06e7AqnVS1Bch21huCpRa7wk3Fa9ayUHcKYeUCryh5WzN3ozF8dFUpb
9s/WqQFrYsthAGJYPbEn9rdDtN6g89ncYe8ndQv9HppMtYeBi9u+WiHxz995
g4GEFf4F2Nc1HD/RUeCLfwTnYCBqgHp1psjuYjpXKWRK4IXCoc+A7dk8Mhsw
yXVSRERZ09kiaiymgDURX960Q12ujF49VJH0bqkKMW3UcNtoqifb8qZy5GWC
LitEgqAIo7yKX/6Vmhd7mEnlIbhVTawQNyV/w9HSo+O4PEzR+njJol3rAHHc
V4fr1as518w3YqJBS7UluSW1m0nqRC9AIu2vWOykRmdRRV3B/LhPb5EpEaCT
rD1u5ZjYd/EQudwuKWAY0GZAaZmAXhy+akhuvG22CpaPxzvEJkRDS/RI3Pqt
0F3R1chlKOfGh75E1rMArs5SrUbuCh767ZXehybu5IWhGKe2u1fa6Cun5ZX2
8OcYFgRA5FhNORs6i/lvrHLs8LzdxXAqLqpdcSz5Hqmpk6TkAOfSQ+xA4Aig
FahXuGfJQNjr7uc1CyvW5mHvvTk0MYpq7UW/moTH84PTnIBPtDZ/3m+0l/J9
rXc2WZf4f/AZ9tGuKxrwNZ2vYWa8pKX5DhOWmPXZgFWvPl+xHSWOs1MxD6p6
f7NerJqa/vO7BGLbpGYmMH9I9MviyCqiRsQtGbbdh1AT5kRlroIxH062wCn3
OpzsWYxWeURwoBFlpbw8DB5gv7YMltSiB8oip2BEoQHh53ssxazr6G07jQu2
uw6+ZQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzfdUz6hfviDY9CJJCMnGjU3w5kMvfkPf9msLydmDOWZKn6ifcMLV1yLRLcpH5s1FT49E3IilxcRr5KOUMu1Bh2tPFIHuhf36821PVLVFX5bo3EmAQ9noW0Ic4cHSmdMC7bkfMiFA5zwYxeZwy9mT0LKHhjMuYaFdR95YsK0XnhqRZT0MfSXNNZ6qUsuOAsIIwuDwbZDWX1v4DgrA2+EfZjpgK69Rrxv8WBUWLKkPTenxYF90tBn+naDyEsIiNIr5euSo3VKK9G4a+j2b5BisxB5YptTM9ZCtIGejudgZ4LkJQJ9J3o96hSJG7eO1QKFO0DCfaksm597/+n6oebfLkgGocOkBvY+ebIWkk+Y9Se/gzYF4i+yUNwCtO99xa1WDNrrat0pX3S49c/Ad5RF5nSkBreMIhAtBss7/7KyI/b+lnHTHUNJ0YMtRzyoDYhi614Q6k710Bwvlou3nDsawxIJyjh87H+DqX7tWakHZz5NMoAc2l10MKxHDPD6Z91smJfycBCX+5tmJCEIHFRuFzQLqT2tA1pR5nq6haX0J2nhycnm4+C7mGdU9opM3lSXBuUcPEatard06aJgQwJYI0MA31ZnsvPww58HzQjVtWQbxF8k9FxVEvMhWmRwR6Z+0gRoiE8QZMNgff1z0dSa7B9BDOmVB3h0k7qY9BlHD1SCwgbff+NTVq82NvPQ1MFg09cpYm2hdllRW56QYoecSiDFkgvbg6uell6c2j7kCaaXZqGGSRd0IJeEZbNaYo8CtlSOkWEul4e66Y3VFKuTGhOW"
`endif