// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SN4+pu071nKAUtTm0LokQMevsIz/hnBIJji+U583Zkdj2hgH1XKgoerYLzZP
veIlX440f5sRqeXFDK10PurQXF3pW6fO+X8D6yYfGzrqNKIKOF7rCtnkG+Xr
TnFMDlSemtXMGXITfSyrwGzRUCsnkazoInZXexkCSg0w4Paco2DvmHfKz8RX
xJkoxCSdOQx1WzrQA6dPiDdKFscQSDPpGb9oO/x0LURQ9Hl/6w+FetwS5TWj
j/jP4OatLpanyLKVwo5z/4Am8u4UTMHydiOOsDYVS5E5ZkgpYHP2nN2QdnME
MbmmzDrSdHxsByRyZQZZ9N4QaU/oFWIPyHyR4qPahw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HdpklJcGFtCKPskykMqohWJ25zm3slDhMP1q8dae1W5U9jxwO+qwMoxDSH8l
F1wNGuJ+fdfPRyDqQItC8ACSI4zSG8oYF8OW3yK7RuFQoysbLpSDpENlyUpp
cwwn/9qyMIZggFoAC7VlsDkU0ra04vL06KopffWQl9hUQH4SRq++tLBT32qd
Q/4nYGaYvOS/lxSfMFlmkUPnIqFclGoMQ/gj8/QPwxboJeoxdtWn1FRFuQUr
F3rAaJMT96NJWo78GEjJ5U18AoEH9bvALaYG5lUWgvrD7kGCnYVpt0NN5Jxt
ay283cTYYll1pLSwlsvhxIVr9sO3rbeOL9HNGnYpSQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mOJUZDUkMsUbLfD6+UkCofj39AnDyz2MMGQ4muJm+/sKLx9ekGBrSnACKgO0
ePa69E6gez5jEIbCpQAqJPzUqUI0x+nEjxt74jy13ceYUFC/Caf1bU775BH2
EQcAgJU/tA76KSH3DdwDpQSIRyluvdpe322PCM8AOsWa7n97EaPrtpxfZqlw
uF+pyEin6l5tB1/vy5JgenZDc2HDgrkjTMAo+Anrdh8qBvvUn280WOgGgrdg
VIjc31+GsYN4AJV/rBUGzs8HAoMg2r/L6+weTV4YGMdWnRcw+ANNn76XE3Em
18iQpBexFPLlHhMtBfilcgzQrzfSP/Os346sW429/A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
m5+jdmgOqgRD6bmHN07qtLzlo1U4ogjUO/UYLS7FVGrsWDzcofLbiucXvTJi
mnTh5apRh7G3jKbJ1p1Buq9oqX4MNDPZ6pZHC4R3Sbccyyi8wUXcZZl/bMAO
RABF0hmypRMFwhdPTA8rkVep0W4ojNykszv6Kb5v6q2ejt/JpHeWGOFCibHy
xcdchJVR9voTIXLXjIMLEDlOD0GxK9K/6/cEZU9395b6IDTrviKWliAlif0S
d2LFXASLtuSd7p+HQB9kHsRdpy8H6P36odEkYNfwOdB7OCqqMOPNTzlutrGj
RiU55j+Ysz56PsefVFhHQZA9al0ysDCp26pBYycC5A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qw7OvSxieOUuJ3C3rfIkiKZFlB1vp/L9a9rXv3RxaAJGdEEweTZlKZOGYS7P
YFu/h17cUkOmLjaRIDB6gHk1UFvDJCZZe9c0XvFMNtc8AGCL07MWlVf9aLiB
Duvz7pMnQ8nVzUPcqsctDPvzKDh8E4uQOW03q9I0itPeRKaF+mw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
QqcEJmTQdJt7MlsGz60j0ZDdw8u/c/BEfevzM6jgH54Wuepic4zgLuiwuyrN
lJMTrvA/nMsFTUxjDf9QXN4VNnqHR2B48BL5biRaR4PX1uQF8cbYe2wRW/dn
U8Dl2b3zuLDyzYRKg467cDO4m5UxYrYRR84bdaHb+mycyLdF2hBjkp0xSYPj
F5OSxuNxj5oe+G2xs0GybX2XJuQiYn6xdpFsbsEZeYJZjQUjYgg2fjCV1NzC
CvCoQye44D2NFoz3j4eWsy+zPbNGsU35eafGVd00XLZut0DIdp3CGeDfJAtw
weZqEw6xuxiYdwnOVQ7PUEnSv9Xc3aJ9Sq6ZePV84cNYGV7EKa0T5m432SeZ
s1ofVFbWVAB3lzoQ+XOO+ws+cQ+gb8d2RNTE0ndpMBKOHOHkjr4kkCpjU2wh
kGnXBW+Kl1yDxZYHU0E8QcQdIGWJM0chHFrX9AkcN5Hr9ygOz/TtB1QOkJnv
IDy5PwGFzw20eT62nIDbw3qkyNSJYtkW


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mRCS+E9yFhn1y+fpGtpLNwF9YDjtQT6xeUzzofs5dQyc5w/HuD4Z1bmkwDPV
xg2lF0KMrMzFaipcyCY2jrbE9cimjJrAylk8kNcBox4GUa6SBSgQz4gMrHLs
CtuXOFR0PpmXnBOoLn3gmABLoH1v+dSF4xoNUBl0sx+HVE8zGbE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
CvVxle2qQbo+gEz7CSaa40QsaUmoT5TYJY2TNuyE0GNdAgfcpWk5bOXzjD+/
5WUdtWc4RZeRpM4FahFaGoxi/ZkKPcL+TIll2HrAUg5EYIeM7rMeWC7EpH9E
lC7OnOxUvEoUoGPVq02C+cN1Qlg8oRpA7vzh0B/r3uOjwdxxjcI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 335776)
`pragma protect data_block
wqXnCyE4UNRh0ySe4lxziQFMDFhgn2p7M2rBdDVdMBOjSPEVMjm7jCSy9e8S
DA4bVORHVTECJvUV/LHCLNvoa/MIdNvuIPUPBMRJQRdTNLyU4cIM75ZAGbyj
Cmw2kWY0jVbGrTcx4GSKaD26JCFF7H3PPEHi3X7nCi+bht5PLbpcM3V8gFg3
Gl39KKQv6/z2qVDb2SDViKHj7Wn3BQiAyN3G9zu84Tug2E/lMM4qFN9hSPu7
LXKLRO563bhbZ4Cuqnqwr2UadrhMggUhGgUHN3zo26VMpB1AjnF10GoJzMKm
SeNvjE0DlWIEksUmLTWlMHJFnI3KG58kCBNDwk5Lin8YmyhhMq8VN91PBY9j
A+dJbDNj6VHWldEUDmm9cKbCYGylXHBjDw8BRVxKxJNcw0bsurwRweK84A9i
pTz/oSPp0poYQTQRS0jlbsC9SLnPDNr6XCf2ySY7ag3dY7q/sdrdeZZwg6Is
QDtrSKCm2hu4fZU2PbjodxiPADdKQS7pLFC8KrgMltiWHPsdFXdssLTLSUqa
d14DV0xAJzos6rzGOgPP+rkWIAZKSFkRgdMvjLapOWMzf7gx//u2lSISZp1Z
DR5U/8MU11Wdd5HR+CsnJs9SxuJwKBl5QMeKRRJZJS51dLsdWZqQrrsQYeuS
UaMbJNvtDJVlEIuJhmjcTkLNmgaMQRBTwhQzn9MQ6FTs88XwG2mlObdg0v/9
lbgi6kT+90uK8yUBnFxN6UblOLhtYsVC1lEJbDy0XZ9BuKkrp7BTojs2/ILp
5Y9shmXZhb4jTz481dGxcL2F+nS2qsM9D2j03PXzVfLyUiWh918P+PuGLRsw
RQGfFLsej0XNa9hDKw47cc1tv6+5a1sCL47ZzQlnAfr47fkdz7BJ01TrKuk6
B1tAhbeBHoSNLQ9OWz6REfhMCRXUk7Gyp2+9R+/kxTCoaXuQDnXxUSqOF3hc
rrsD9N4RfrRK66GIv4ywMsgJfGT75wjqy/XpoyV0lFeqQBkOsEC27ZBIiYHp
UwZFbAjoZ3THCpIu2RPPYINShzztBh95vTK/AQ0iKxGargfDygjlAdYnNza2
39kLiuUoVyaw6SPPN6X+KcPqaC01Oh9DYZTzk6USGjKBQdJXAiQ6vukROMyb
2PiAUCtMvqiEDlnjFphk/brNqVGkU0dyRcBBRtmZIZlAB7vuJ0p1nyXNCp51
8xYWvMdWo6BAY3y/q+34ihc9wbB+iYOju3kZzg6GZP3Cr+BlKN+GCFkaBfvY
urqGXIr/eaVar1cdZVDoURaY1tBifI+fTVSNhQ5Blx4nbXMcW7UkeGqiula2
2YAmvfPy2JKoRJokWIRjEv+azWBRF1aEx7ltv2ENe42Su5fDWyRZkg1mfts6
nmxyvX4VovoMbzz8LBi6gG+e6x6O7iBrjHGRVemLfp+JqEVQTtqtg2MY/5GD
9K2mSltV3tibeKyaEw+YBiSR9X3gfyFr2zxqFnDpcC6PARen8rM+4tEYiAbc
pqL9mk5d/quJP3zV0kPTvy7Sn+Ir0C1Ku8xOjQpLzKuu/VtC3ijWPZuUYbsy
igGxkjuYpJvIc+nPjZVREMQ+uMx4TjA82YVTdDSJAQZyYe03ibtlYvszZrzI
SbijwHKq+qwEsMQpJFFVHzKis2mRlK6PhX3ZN5s+KXHOAYlUfhtQNfHsWuZ0
Jqn719HdSXCO/svn0LwHh5DdDScFzGXAASqYXEwPpw075Ij52+sreoWK70/f
RGW0NTUPtTfh87yqAs53zgL6+i0yqBL+mSFh5NJFP60qe58fRnu/FZWz/gVV
EHUDBt8+XL4YC3Uw3Icv07tN+DVxU9bb7ZxgG5jXfJ5RyIa/y2rokCtOYkOq
bEOkRAadrGZgTlGU0Tkb4sskld57PefU05zZ6d1SUYH2yX00sq+DNHTwUQNx
Z9Hxh9NpNoldgT88czS1Ub+3bbp94nIVbpS2cx0CjQHYApPcNMgnYH921WUF
xHBRwGmPHXpw+DCZdbg0ObRtbl467j9nd7d6OOys8RHpL2BsE8HFwRC18+uf
bdUPmI7DPYDi8SgQ1IPWCHhVN/V7Enq2xZ1OS1MAfaxMRzSqikjciJjmNyeO
SyGG5UIImm43BXRrBmyHdQFRLtJaR4NqYHL1O9Cbs4PfZxUVgSFWui+2jHq0
jdc3eXjv7D2QjAlCDveLC1pjPAupX9SXPTT8L1R+dbI2ewnSWNtAFwARaJuI
j59kZa/63RalYmgSU647rqgVEz7gEvQM+v547c+nifNOcTurbT2RbkvDD72f
mZ9xg3wyCK4ZgD/FqwkfYyplGJccOb77zn4oHlMRFM7+mH07EYbgcRiyaMlK
1qwWCI/3aTSfGkIJIH7FxkXZLj9X2PpWf1e/VFGpj7zYQtI5Rp2RFgZDwIhd
Tf1WN3SsR1sB6fhEqPgyX+5t/HiRHqw83qYIEqzTDhy786PFzsUNAyVNmYrC
BMFMaRd7UtBaLyiGLxYM/WDddU6PfbKz5RLa96afSM4CPGYs1JNolZz+Rwz4
i1Se02zh3iDyvlR2D1wNpNx5y+xlMRqextXnB4z645tAHBdkxUG7rOf+sxmw
wY2XaUjhWp/g5UYpfBOgPVjbl2CdFR/G42OMODEBXhy8POQ+ryg0vEkcfNFn
R7ON+XZ2tiSNZC6ywhT7P9ulV5tBUXJrufKRKmls1sOHHVjiwTuwqmHzLJUK
S/+koiLmDHKezBE2LGTd0ZGxUV4eJoaGv9Mmd9MTMvBQNM2t+snc/nz7XjCG
3wtBRXND5orIKUdCrgaXl5rsOf6Wkh9o8rCZ58hD/jB3aHOUX9nJSvXgvNkL
NpEek4Fl5M89EPcxFhQhZfJ52GWkjuo6wnUVU5A7qRhEDT4G1xMe2y03vW/z
byAaCABKtRW/p1AGyIr6AAzQfISm4pcX8AQTO/hw9J27NnG0LwLBDrIHlca7
hpkfYm5ESbgYlLWA0CWTc48OxjfzTcfoJxcs/PLSQeV1ZVxIwVNgJBVNC3ws
EakmuB4Q4T/Y6MoVEZTD8gYG4yKqpSAqh7AiEdd8FUHf02S+VaU8C1iwF8we
lz4yHmAAuHi0qB4NTMA+fJFYn7QSPHBp5qTsekB/IDbcRuJ0rPSBj7OfkqoC
hREm6ceC3aqtqKJM532sJzKVT37cO0aDzVlyFDznhF4Twl63sRJ3Yn9NdNi9
RyDmwkHLLpU2vD7FvFya7UxRDd8Qk2zF32+v2BDmjwnK1moySWzvvgb4b1mk
Qg1Bypk7PzgtUlMr6q+ydACg67AkKdAUg1PomNRltFuC+m13i3UmjuisVA4e
+JKmivAOXnlVJoBQJ5ErCGCkvz3Q2qk01+0GGiRY6NHGAf9URReDM8UeQGKD
KKJCcpIQ9h9QjbUzpME1/UXWQQxFgBf5SJTObh4B5URRs/BoxcD0x1t/hm9B
I2PPL/WFsFZRv5UeY+7rvhqOUTxeHuO1p+83FZQTFRaSG6eecnaQzE3Q+wgL
xqma5eyc3OCDsYyOZ7q6QEyGGYdeWuB6Pgd7pl4FKq/970a2fUKg0Ira6FQP
RfQyQPx+EK/4MtUKG7VFC/G/itaUUXYwipz9nN6T7Zh81zD/TB3ZcCPLpnyN
s8YG5ZaZh/1GASFIsS4PWk7xw85zVPntsVumr6pClZBh72TgVVSKH7thDYmu
QcKgAPpNywuKHvKjBx0Pz0ZV2BsafW+W9TQjO8cn2HHNzUmup/T+TuIK2/xG
Xz+lsgkQ2+fqgsJU8tVPTJrineMIidVXKqYEBVVp4kVvGNGMeARxZk1sqj3u
2W8IYo8bKLZVBMU/fxZh9Z/tq5bA5qSKpFhjYrorPpiBe7vumpuBbH8zt8Tx
1c5YU+t66mTYQJCdxwHSxZ+cL2jzjgDb72EcFLJu0yLYsReDaPcxGnPDWIoZ
JwYaBYKocasPpGbnTlhrNc+cXECxKll7fU6h1z4wxCyf03qgJoi2Yzf1mF1V
erFuFU9KF2OvqLKTZL1CcbD3ecDXn60W+3Z8qH7u8Ssl4txqZ+rKD4nGUPRr
T8Nr33fcZNHNi7D4QCld+i4kTvqs2DYYvoztTgFN/VYS6A+8vc5m1O+jb1aU
SCCx0W9ghCS8j0SqSyuK7RI1rJqFKCuQeyRe3xw3tQiHiH/g6DSgKs4g99K0
nBAKdRJcx+z0QIaoJvs3yNr4hQ77fPnDHgAZyXNPq75Cq80Gbxrf3fVjCZRm
W4W65Ds7MquKlGa5H5V2QlfxsW2NGUIBHbsgi+VN/T7wcZEwCB1wH424wzqK
9EAhdhUfIoesMx95y6v9ID4pJjCdWTkoK8fprNcVGGWGyzR32Yva5YZIJtzj
KAKnXo+todIa4S2NEOROeL4cW8vq/mmlILdaXcsiBWu/+1+FPUZEWOvzdKa7
6e7oH/tiZRdzpC299QGax5rsubUo/zthBEFY/M0SU1J0XATWJ1unJP/rkb7S
HJJiZctqWHaLwyb6YyiOEZ8G0o74hFhCoXfQbQWQCqqBZaFkfgeyu8PPpYjG
+ffVnWUxfKBdw3ojZMRX6v4teZ53/dzWynkC+XhBsohK7a7mLMSETzeXmXBs
ADM4fwmJd9Xb4vlKhybwaPRT0NKTOApL13f+1LBa66qdRs0Vxq7z+bqL8A+y
6KLcIACMBILKqepExdld0pIdpohwATlZad1RsDNNM4Njyc35xwM56S2JmG9m
bN9WJWU9IZikxq4L5XNHsKQYhuqUocMNQasfL3V1F3+oiMuds1OmDtDY/CNT
XfARgLMlSWHTtVmuB8YbrxPwsY0iIUVzXNlzQRtHqpe7NneaWETHAdz6TXsw
PprCD5tThstM+Qa8jd04tWZIyXGFY/kyteiJSEf8+ArhplUI9iGDaSI+OxHu
sq/VBKtsisUBQcckB37u5RujSjORvsnb5U3Y7dJEZ07cfusz1wnMJXv/7Eq1
6tt+yMwfeFkbBytffCqYe2/S1/HxMD+dqSFA9Cvb5Az5APw+Y+w+0WZIQHAp
1xpUcDLFdL0MIwL26XMikc3LwJ3DlCEJzx2kvAdQpt/1JHUPCbSzT2bd6SCa
NCkuZS/pHXEXS1iJyVaMQfhDB9U9waTGooqydZDV/g3KypNJ7u/h1EVfIb6Z
kfygnmmndF/ciuTRNtQQWJv+6XGyOuI+MXyot2ZH8Uki69izDXkYpNhNC6jX
pVyXHyCB1MofDPxa5l/a5GgNJLOxwePut7sg0duYscC35v6riHmSXyg3lOSS
8GQkH7VFove8vQfXMAtAi/aYrt2vE53f8W/CboUoIOHUGdg/Xurh6nbGv4L4
ft8lLmBFPyJFsp0HoREWb7ydZAxDJP7IuN1mCRnGSeOPo+g2uvDy9cJCvglW
JB7k4Iz+i725J8VkoHkD/wPHrXK0roAQILuomolMSwPDsd2t0FSUsOOjUqYE
dWo2r/2jlOf10+u/34jS7DNMhkWw4hZKxpb/enbdS6sCm4HzqEWkdrSqLd6O
AyeMOFHuDPe7X66oxQXSlAFRG60YkrPUEQBtvsIw5chaattL3z4zxtOIqtkL
hJPfj60pPKtoQeRSxmYydLQ0UYQLQb3LK9TIWvYAaB/2ATMF61uNXKP6bL8i
CB4m71yN/Omj99RFq0E0Xa3AyoK+hFln2d0qWeW1CJhwie+oR0qjgKEjK0e3
NmYice1fkGsotc+h5zuonemvTYs2BrKau6GjjZyf4PfetP/539gbmioomzDG
EuwxA5FuPauYFrJ0txtEoZBGhveci37H3Rt6DShCGiarz5tiEOUDB7OtS4TX
uEeHMxvs1yJ0ITuoTzyiEpp+bGlBuUWMBq5PnfyX6ZFJnrX3b/kkccMudcQY
e75ToEy7QcLQAcsyLoHfN64lO7yiXZWU4g2u58xDaTIwcGnNNcOoJ2VwCW/f
xyyq+wo3LNnELDnWMuVrSJZcYmohIwxESXVTGyyOtOcm9qMtMUb6xwWRi3g7
0FQ3WNSvHdNhTiF6RlvWkGxJAGdr6Fqklda59HV6MLpIKR/XYCS82aC5/hDB
ZWcmlFABg/HC1q7OP/d+VhYOdhsWtyzRDouWHNYal32y81doC7ZQDFQvkj3K
1a5yaWGepiUyM2YU6EvUXurE4b8Em0zJN7UYFB+fcUdFLU7vprxzKDj88JuH
kyMDA/TOodC7yd7VkAHrjArnBcID4HfsKRNF3DYzVXPD8r5QNTbmxk9XDL3F
VxI9mJ271qm/lYFI2ae+ypzvj4T0PLWJo0Ffarz1rhCSEM+2L+obNC3Pj9Pd
JFTmXwYPtK6TY+A+z+ZAdz0/tlFLndIo79r6oUKbVcdZXbfqkw8oiOpxrVXz
HQnMBC5VMEp+QmDMPRkg4N7ncGg+b8NP4b+VNfWUsL50B780wqHqZLOvLSg1
KCbOikXgnUw7bDhuSPQ1rwDsD+XJcUapkLsQJRGsVVb4zHZgnPTnbYsssLF5
R3QCLvirMb6ljG9dYsd0PO/BbpMt2fHP70qqFewAi3VwlcSp76nXANCx77WX
/SqiXJvvCdfTy5VMWGl2o/kSvMGTDqHaIoRIZvITvW77DdmwLDlcPc++TZAW
RQiPfUh+WdUcbDkbBKA4sMByYrTN5VSxbCvNETv/RPb3yG1cZGK2jrc8os+D
0E7KmfXmhiz10Q1IbexpLteh9HIr55q71/4wNW/f8utj+cuKEDaEKwr/G33T
oy6L5/PhKTdbqJwpK+fxDX5NsZLlDKfWcGWDBJXk4CI0vrEB8GIj3VM4C2rD
2YakswnTrWajfLvoppqvAdGwTDLTweB1YqY9i6qv0GmE8MXj4YXxz7JZI0hI
M0piq+d7g/qb2C83+9IcH7avPRg3ds8Zkrrugp9dKZNUHR3yx18jFIDh1Skd
e73AsINhEdxfjUWBashpCgDXcdYYJ7OA0NI3ZOaGlV0w35MZkeUUn5XYXmFs
xgAZOzWiD8/OMpUNhX7tqYSeRIMWqoisd8AgvsDXKukv70XQQ4NvDo5IVsb5
OuI/KRjwu2bHIOnJMKP0NTLutcQvKv1t6yU3FPZkRdK/e9e+Wny+HLP/8Mvz
dsZKlm8gPC10skDDuTlMqic2hbIbD2MJkVVzkAmdIYPhba8/t0VqLmY0u80U
eAK0Sm8YqklwEwpz9yOONCi5zPFSSynbdq+TVyr0NkdX9fOn3Mchi44Y6iht
fgpURbyvtR5TCEYztDJip+TmhVLQCQOyoBBDrjC2vgTtvHMhyo21nEgmHepn
G1L21jQDFDv4Mh6D/Rx995lGXdIMkihm0qbMLsVbEiVltrWsyDsnr5wmlAIz
YfJuQn1dFWi5sB1YeQdEgnQt6CH3EEqHx9CI+21ulbHRsO9HBBdr9V1oXKlU
PQfGH51cH8J348dXqRJhfSvZt5m9738Gz1dMwHUqOpo3AfeRbQKGy/iwl0Bv
vA9rUIXiBs2OQFbTMu6YUurpcZ2s3q0ttiTsxdUTkRGJjgHuuyegJ8pLffe5
xrc6Gs/QoL8FcAkjvAhKOPMqS1HymNHHnBmZyzut0o64yFffkznHvki63LuY
zJtxk/jYTxHI4iirOHepDCrntBwYOIJCRzFxISx1Iq7FfMIjhW92R+Hk0PyX
YkRBmL4mzcvEv6z0KRkvTvph6NiJ4i3sIMquhI+28a1DC9wm6ORq2Txtvokc
rHh19FNW+za2EmfDUKPZ/Er+VVXUyxYAULUmBzsPq6y9a6d+RzPkI7uYrYrN
mzyuV3efbJOJeuksJMM+B41fV8cz5icdGc9xps6cYRfn5TQEgWgcibAd0jWA
BjYpw87YV2CySh4pboRH7vNG/8BEqAU3XT4NUDVzeQZDcvn31xJMTR9PJbCg
goAcfnmq70HjIP5poOPwFhYbnQxoH8uTUEA8MXgi8w/futOg2/MKVvzzSILx
GrKWYgQcH7+pvR1GpkMnOcAIlvvFKX3POGvnB0Q/9o/HEAVQ8m93wFjmvNRb
RcWmi/l9fIZQgvWVHZ1YMDAto+gXUNe7kWyhkfc3QPMugNpyrgxeQGjUrPM8
k6VNmtIVo4bKYNeOxHSE8p96yNvZ2IL6PFo6IrD+sKjY7iyQMdvOow6vdBVZ
5cDAvUjN+rxoBJvX0Wt/EUU1HnME6LFTaNAARpxIOcSro1flNh0yRfO6dQ3X
wp5yj5zrWEZtD72Qmyu8CaWW8ITAPuIbVont5BO/UTITEvSzmRmmUJM1ZE21
/UN7O0QwyljDjsJ/bQCL8bKO64DU2Xa3DLFaJyjV1zTjeZt0qptulVi61zFY
v8FTwViAhjFnVkOM+7ay6IpcpG0mTUo53zFV+wRSeOq2P7xdi/wTUbjuOW3f
GYUER5qV7TZY2l4b602vaKUCt7SuLrbxEKzUS/OsC30ZuIthrOGi/anNzjAY
c/cql5SGB1PDpwczWyf4zw28Y77cmUupXVVW0YJPg/H36TcIsvwf3s18uuQ8
7y5d6FvWibNUVZEx0bnm9E4lHnCL2WAxMANuByiz1JN5Dk81NPKaRxRV4s0L
LokZHPOscpbdkDJkeUKNAmCz6zyauqzokClLZFX9BOJEguZLfVI7kIxqZaf2
ckNjS7BNiamtsTbar31kAdnspR3QV2d+cUmXveM0jreHx150Lg5dT4M05mb7
nRwLUN57E6EYaEHAxgFDd03t7xtbql4xUp5njO+f6+gTVWxFYQ5tCzN3fWsh
BxwdAJw288zIQHNr+EJPXO0YpEt0OjyUvuLevzV3EVWkm6muvvGZdkuOPlZo
y6RGORmjG0pYnyl1HBUWRpwSwWnbtq2f2JD2HYdrpFKd0GRUYt5MWJAABYQ5
Q8VQWyoBfxAZ6+jbsuTJPKPAFnw6J/afsYCJ6cs6FcYscixxCVEkgAQMJIvf
L+W/L2LS4ENJgDRw96KhB3U6wWnw8z0c+pP62TPPMUWXrJ9E5oV2zrM/5Zh/
CMXggIBs50lRCzqDCBUN8TPw2fkNnFH226R/zkTBXIA0DBAD45MAjOSjs1VO
KoJPe6NlO70ZlUnM2b3Hy3Vh6NZRpeolT+sQ1B+iVRb+lN+PwE/Galnrjd3j
muc47K26jhEwVjU5H+hQnyIvxnsfxFLbMyA/wxl8wl2OJfSszEchADCJrGoI
fVhs5kNxGI0pnRY5p3TGDs2Nxu1FGT2bEqtu96SGAQJzIGGfBI6d6/d7F6og
DkqNvuKCFE9GzcykR6goi+F/AOgXjdOVvWKgdYvm9i7bGEpU1Qq3o8nc8ZIU
78aOD0S37FXrptnslSqyGeTpYqpXbfGsvqodCBL11XxoUyEXD+VgQ6s9qyb8
MR3eNpD02HS44GiqhiGyrrQiADFu+JNV6bWSnqNBitHnzCcFLeHx8hwMHKoV
ncS4AoFTkSlaK6hrla7C+j/2maQlYY68I7zxxPYISySqfiKO18/fe6BP+DRn
VVe8v1RlBiHN+RoFC6fwj8fEMjqG63L8ELJApwqj4l0aJyQ63f9OOk7+EyKP
LZH7MDbfnWSNPyVks6fkZWDUrXRwM50ic7MroUSb73W0y3zfzYOkBuTLEDqk
NqebCMO4R5B9pJGNTBJPjQK0GRE1jaQFWX599vzH+iXPonfdjsa6LoqEETOS
E2ykAWdfKwe4CJeINO+lxdpI1vt2iXLQQwc3UMKOSQweek7N7z6MaT9lmf8d
rEA4CVtepI0M35Zn9yhEeJamAzqZTMXgh6IaiqvOuKQ5TjnIGJJQpFDO8ttJ
zrBlmDpCMRMqoVgsEjbElDCytusZ6rJu/ldN+Cucak3Z14cyJca7TeQEGQHY
IFYuRg3Ob/U6SHcW7BTZkGPFtjahdza0DbcVt9+WjREEJk8z3lW6WJcN1Zr9
ZpsOZ35oQk6MSml9xQpRxBfAFOS9R1LJzc9Wu4O4ja01f2lVTW38MhB4FomF
ywQbmqlbIyQAf23fB4YG+55e9cqeD+idQo1TACdxqplKlK1gyZs+6w341KFA
BzAe5KZeaTB9Enjxu782MsstKXFSftLmo/OQ10KS760/CkUkKdlJ1RrFI7eg
3nc68nmB/nRoS2+4/2BxsrlaOxhcEo4NRcXIqoPvLe0BK58lio66WWpm4rQS
Z7xvn7M97bDPcXxdqCR3WFgsyGV+Pr4kaHk+q2y8RQ0p0TbbDfjrDbvrdEzO
HUzmOX43eUnjI3reCIQDxY+qmLGpg508HtxsaqunIpuSQHSMdLAAT1TCvso2
wdV1vZFJESC94+HKelc4BzmOj1rF8p6GKUbocE3O7SWtwdTUGjllDDL4PSuk
GZNB/KHBFnr39V+XC3r1jirYyTaEYiujzIHmkoYboaWrTol0f3effjps5yu9
3lLH+PFce1mMxYfSbytoVu813KR0i9tGJtU4/QyjDgesFygmO++Xy2PYaGUo
R7cmk6sbQDAhFm84jGZoJVNgSpN9IsJp9R2r0XZBcGDsPvNU/QY9pEsT+K7G
KNGCaB5rA4TJ5RPosTCYjABlC8eZ931VHJY+luoGlBMQ+UAxXvf8MWHnjaa4
9mJMvT1n+swHrJiLr98PbKpMNl/330IkE7Oms+wC4530HZ3QrWsOfrDCw3Kj
MJo9SRCurORe/X+0l68DKhLVXUw12pTcP9P+rFB94txHyuQTW7y2vsvERTvI
MYfOdnQ086bwIdcO0YboPFD6B7q1/pc+igxiitUDFfKYnV/H1WK1qF3/T11a
nf11UHY1D/M3L7yYvazr+HHQ58yaqH2e/7fH8o0tfppPbK+36hguKROX6E6l
sE52TZuIHfrO8M+RYSFrD2LWL1Zf8R8xeVLRTGyGwrrIQBzjX/szwioozD0q
Xtj3+ELY+wy4M7uPka+95NQAK+auWDpzmL598IS1GHq55agwsD0OVNtcUpcB
avrDzYfgqSvZcng6FBJgVIDcQvxmyYDhrm+b45L2FQVXgbyTJ0n++PNJRXmI
5JxvHAhhVtKIMRFyHYpRddQU/JafesBta2wlsiMiwgSCkVH6GouqYXiqkuZI
9kG36ZTrYKoMX1QRVmwCVIuCkcb22CPnxj+EBQfBkOSor1gnfqCUvv7X7ARe
kZy3mSVlLVD4WWGfUWeSzV/8JvA+858dNawlxWbhCNdIbGgloVqvXjCoxPes
ZZB19sAdsnR8KGQgnfF6e2ENJRJ3YtoTQ9Eqj9taUhNjdK1En9/gWXUQ8D/q
YeyZPzafa9LoOtMqTkyIi/sz7ko6n6nZmvv4BjPjluUzWBoNj9tDVta9lLs7
pvFrOQFKxdtONMi+XA6P5/lP35KPFdIXt4Le+mkvDwx6LU59SBkHs5e611u/
mueyOfAlKzAVVgYnd2Lkfa/W0a5JsPYoxURzVAawFYpbiKLnILTHStjpqH64
g6tJNgakI8IgKbSvPL+u4cuK88Qst3ZXFH4BnBLopjsRDpdQ5ftR2IE9hcq7
OyUb6HwOAfvzN7XcBPPHAHG4C8D2YTsYAkQ9jmPNfCIwn3x64FLo4+2V5ihB
4af27YCtFb6EZoIvPIL5H0gGGKlzo5sHf8SIlDwdlwDC01beYCx0Q31lEEaz
ODSAG/6P/YZg195HSHhZJRp5C/Ba1OxxW1SWVEbQUVkkZhtMISMfud7+O3dO
iVWyTJSQ4+Tgw3S2AGjrL9q7ZQ+Pfs4HxUrDqh+Y+mmcf4ygJXWM0dTXZytk
i1fvFGxlLUCrkVN0DYuTJMmGobD9LYJfFpKELvI9oV/vcMD2Je0UAIcP57j9
CYIwa0DuywBHEEiht+2ALuyPcyLMKXrE75dUNBtGaC4tgF95aRgDQHdCZM8k
gdrlyL6M8/JDyGOBs5JM01CBwRA5GYrOoX7d7+EO7vvFYyzAAnbKPNFQPFQ8
4G/h8tEVLcDkCzh8+hgGl38urIaAW2y/EwZBedvbZQW35spx5ZXf/ZRPa/Nt
t2UD887cZAuAIkOLl4AIOOLH5hPIgYK0djNUQ2MiAXpvKROKY7VscZluN8ac
WDp6X8ch4I6urfW+qOfo3btJUzFf+utR7C67Y4suKPSXBPAZ4WID0UYW/wsN
ocF9Z1oMq79370AbUi1Ip4eAThqOLvLXwewyxQdsC28nUqbFhtRaJIhDusmL
wBjAnSbcPQMqFrfSJpuGcUqtQ7ABiD9GPsGyzkIxq2DMVLRevc2VBzhC7IMb
zmjQtglEGMcg7ZWbn6eMD5HOUd0mTQy2tGzOvAJJ91X4FRLbWSRDSfrAoH85
0ctDCJp8ax0OfKXXET2ZEsafy2OCLWP658/RODUxMITFdaKFI/TYIiwsNc7e
7TKRdzONJgLbm39WIUTsJszCC0JEwyMGbdnufnKASgcOekHThx27VmZoEb6V
Ap9A+pSd9wjCdWmMak1CCCdEXsOIHBrHROQkhO4BG52rJkvEYhvWiouA3rCV
ciAgTiOAMC/xgQ71U381LPrcov6xDyRmECYsIilwzEZuGC0QRZC8eIc0wk0a
UffwO9lfCMCgBSBCNSskK8Lgc0h8rP7I6lwo/VMzN8I4DmKvyACeQyFFXYt1
zYk4i6WIpy/aymFlB0OArT0FDwD9RWHDSKnU+QqZE5Y9Q00BEpXJTancKxIU
nsb4sQMDyIrVBWlO2NqgVni67gHq8JpDdLmS/WBKInTOHb/kXlEVk62YD+qr
2q2WvO7lq/DvP1CVkUgMJOvDc1r4SFo6fwS0DVNUM2ZdqumsHl1I1HnuF0Rg
R9Z7lap4HElhwMRN7+/z8ilyktdLT1CYCYal8hLGDHvSwugotbZ4rKX7a0Mk
Trbc4BS9OArJ3uUC21Xcemi9Dw/9aRh7sJABC2/hWwkmKENLEclyEJNaaZxC
iIxWRjkQztcphRr/rHs8/UNJqBFMQp56oLIpNRkoQ1gGoeXWTDhjmUvHD9YV
koSb3G1psgEmJ/vYEjcIq7+VB/zRXFiVNz81kiL9MvKMLeKVfst6DzazhsWK
S0kV+2RDrUG3bKQiRs9gwIm5TK3h01jJfWAcABEX6CyIpQ/shIFF203evtIf
WF6pqRX6dtEgeKSy6olnEVW/NXeKMyysY2QZTrD+SpAWPYaD/0AjLbTGX6Wt
QLD1i6Xa9whcXKa/H1QgtrLBxmNzvLSHoRpHxuKdeQQPyIeyrlaAYxeuV62P
5sSZVcunbrLzMTPj6FZ+9npdFE24lPfm4xd03IoAeHkoSECqqemsCFKZsw5+
Elht8wHIDxBminRp6qjkS8WxJzb5qdCBB6TJT/cb9wIWjyK2qI7MY1+1My4z
kfJhjGPKlW0Q+YkUxnblH2OYq2qQq8Y+yy8yjhxSOCVOJmxjy4AR9FC4Xcn9
flaa7L3/y8KIxQ2u2qZl2x8NmDSHhR35OtyYarKGai6jjbvRk8YSZRrzEGSm
QGARG4G5fV7TrPk3Z8I0HrKDL6fEL8uSav1W6upT7m66xRgzYWBCorcSeEGS
7KQQ1ytZC2xjSKv+YkGkdVvpq7n7naNJrQKfByokkeGy1DOKLx/p5VFbtgB1
2tetiDbOFUhU8rCg3rVOoOmjcl2yiM7iilEGS1h/4aDFBaylzwXdUucqgHoR
LSjUv+BF1rMSfZ0BrZxvXQr+9hiQlI+sXkOl44e6hWsoLBIWesF/6Be2LwhK
SOw1rEXq9tfRj6cFHAArFOjP2br0IHX4g2PXxxGvUWP113YgJncNjMHVbDdH
MUpxJlZsnrlojjzkU9vO36Lr/kL/AU00LUUlkZ8iZdeKpQyl8ai2JIHPMwhx
1dBXBg+CEc8kK1fN7TlhZVFTZAxzgD9R60vwTPU/wQTbJkWMtltWTdI0XXCh
RMCCh5rGMWh0YrAC7Z/Xub13vXJ4sse05JallECADSLNHZRx3rRURQM/sZVv
VJjvyj9NqmM0bL3m/RSFnCW/0L8yw4UMZ9te1nmYklglgQ5v9fj4Xq//9fMj
+aD7pz5KXJgACHxs1d9MgP3iBLe5UUOwNAzJTabNxr76Qsk23ze9fa5pxGYG
9UFO5c7uUsYXO/4WWTD7qp1Gn3rk3JwGFw3SaInmWbXspZJK0sg2rtwwQiw+
PXgOVyqbvt3t/aEvbEcLOS9MdBQ3LfdZCEj+I9fpImsPIppIBaeMtSPCA2Eu
67NjtSmCyM3jaHYiKucvuqxHOkSdVXSIP4Y36O+B39dXP96DwZi+XiJrsqSg
SHHbC0nA6goQ/J79QEXDeYsu4KKq0RvNcZTI5xtfFyBI7KUIK/+kz1GSjfjb
S4i6b16dZVncpiZfnkN296uwC90thzttODOk/9nCC4OewXj4qo652UxMmYsu
gcakhs8Lj25TkwvB3ww7ATNgOtG44vpmbYnh6nXRPGti8/N7RBsnXQHgg56j
AMtBTSpoZJre3tLKMoE4zjxQBX8WqinbeQxwWPUyeKG/qKWgnwKfEVSfHK3v
hb1VbUCtuZZL+5NDGY0oUh9oPeUN5t59M8eeNTlRkukp92pw6yqzVbaizJ6r
WtwZGyP/4rJYoAEhf4BPYmJmBDjRTKomE1p3YUVe3xbTaXQ47iyzQzVBFuLa
8ZtW3YFEb+kzC5dU1TsbDnZ6m+Q2mEjMVwVX6uVX7BLpKpm1OI1tdU4cMb9l
Uepd87MEQoR1TkjvodE9shwjfIm6rnDvqrXsoWi/TdzlBOQ7+dAVGf9zhMXm
CVKOZ6Tw4IYqYfpzhXrXb4ansjXfvChHF4a6S1dUJWjzQEagF2wYSs3HUiP7
5vbuLLGu7n4AljHcMthaQT6atdH7bXqS6gkf9TI8zUw1cOnwH5qYCEvoGIPB
+Snayu1uKUDGLWgI7+Iq28vpmQ6YT5rqofqz4HCwIVTNs+fBwAxJgIqDriyZ
ch+9qa6LhUKrjiqfAoTozHIC0A1vljGhlIk5ciJQuWNSN1SUMOEc6JFEDeWm
L4hiN1Zarctdus9NXMnqNw+xlJcmIw/kXEIDUbsmDqsS/Xa3lED7yWd2g99m
K+Pf8XDozPsctawbQNQEGZhYHhSA4BXdicwhdhZM/CX7XSjBmqHZbrz5vOzD
FO4X78NpUCDiHMRpUvb8tL6a5qElvEWJSM8EGJzrmlQCYPJlZ26P7ZJCoNNd
Pd/N0ZXeDhKiI+lCD66/VF9ItRxcf1cquOgRinrShDIXM0qKi1OsZsdDt2uj
khvSfQMzwbCfU56suGfdUKl98aa/NNwMJk5bQ402iW8y9skbSVUjScJ5QOfA
XPTH7kZhFz4B6puStv0ers9XWXI1vOdOb2c9zgYMOAm8AiFhX1WLEPXrtP1A
oaKQu4zrqloNPvqBAVUDsHTwBC8eGfpH6PbguMUc72CaC/izi6vRXuudsOuo
5cA/svLtdI+wkvnUC9D8YDB7uG4r5zLeP4g1/nHVtyZ7OxgMt7da1WtBFrjc
VmP9AE6wem3iwO/QhwPL7Jo5bokZWfEzn+wbbTwm2svTFH8S0FCvfY3XMsGI
ektUWmtwVD6kNXsWujKsriSHIiqydmQFpLnY3vE4Ze+r2eZhT3IiqNQFIgGk
VOfo/YvLR7aFLtgspVY3WL1y+VnHP4c2NKkXMmgF/3JPb2tNhOVzxvwAgbdv
21CtDrQrG6iZixcJi2Re/n++pTDnJtPIYAVnFa0CZmCWAVeJFjsemmmCG/1L
CPSoMSBRznDiPy0ofMhAWmSeyFlBprHyV4eVQRJtZSWNDHg1cU+lT7zcTbzE
HDg9m0c+Pc5XeCrWW/gewqwLUGYXuQDeowr3nP3MRxHrxdktMW5Pr5OMpZyI
nHvWrQ75AtZtHESv/ES4cn0CcqObEM5mKsZnAM3C+2PyRtQzK4dgJ33WE6+A
Nkvod9UZGrwHCseTMPDBV/B9QLuPIPChmPsFo0y/FryLjwX6Orlec40izh71
slCAXODk4B/g+bBhWBX/1/jIXw9910c8fItTCKrqaXXOMEIne1lJCuu2qGGu
/g6HS/i7Y/+fC8b7GWyIiZngOmJrU+Saawd2SLAYETFc+kFLRRIuAzsA75q+
rZvRPPcfMMdqoGMH9zAZo3/crpEPkjuwj/lzt1ap0HjGTDX3I6QStyZBCu6V
iUNLh/nUghqbaM3B2EiIOTvyDNod3a8m/epLqoYHZ0o4wKhC19VzvgAb3eW3
+nUIA1YpSkD6bRVc9RUjTXtJjyvUmDlopMyjC9NMgYELSD4q1ImkBV1Qlwnb
6TAAlkfxjfPIJ3J4DtaXAswLvCHz0BQFqY3NRHNDrco5UXYelj1TGBh1F/Ii
8t3ClJPeg0l3GipxMB0gBz5Rq7t7N6g+vW4r6Bac98XjM+7rtmtkuxsrDKpy
zvHRDvzy02PQGco30IDjZJi4DG4qTaFNX7cd/2VnZS+IPXkGEPJaqcArYeMf
84RCVeA6S4kD5AK7evI8HKf28RsygcXVoWI2CPhYyi2EbvjwIBcxdA5Hnjy1
e+EtlJ5S1clO9u3DKWbPNScrYY8rlOWVE971Z8XVwUv60Kn4utTIXzHg8HcR
YZwF5YwtNKoevCdQFs+azLoLo106BPVcsyi+JbDXq7tmgZLwzLOo/ahZtlgs
GROO5iYBeKPMGu8pb1w+Y8rza71ELqfb+nWoFaBBDJH18gIvkt2lU3MSQapp
RFdlkjMKE1aKmMB8ORH2cKP0bmbRDOP4HcBV0at19nvF9gii98hsGiSpyNXf
XFHi/Npq6YEme/JUQ+8/Ftuuo65Su4CSm4O1jzIaehbfn8fEcfWsNOVexWIn
Ej7ZB2E42JWT+PbzmiUqW4ZR9gvnRj5aW1lmDPrz3sjnUn7nviqsyG3gOSR8
P5+A4TM07pXLthpxzUb/oDzRYIHtidVU4jXyGSBu9mZxfXK88Px3y31eUEZE
sR8iuJnqaaKrM5+/wriIR6LvWOWXggLulNdFTgPDIQIdAVSmKc1IJXoOVpvM
RMuutkH/IHk+EaSkEqaD0RsAcXCEDoZhxLhnA3Dfr+WOLeaSJUyRf/qrfHT+
PgDWHtXxHBsm+ZNukbuXiUjFO4N06exbi48/Ds31R73Bge6WzV7v1ktyYlY8
o6HKhT/7oq2zSFP5FcfwjSsCiae2Q2zfhRfpSZYA9NblZHUuQhS+6FFo/DBe
55Vdns2IsKDyAP/ja5wtXbAfD6x1hchdqDwf+NFTrAP4bRLAJ1Lg258JH5/f
MHk8ZIZglfxo744tbKoGwVy/spON+auxl+k7dt7GZ5Rtfd0wZG1WFrY5v61h
e6PVYU8ru+sHHOTLoetDVrG/ma7RIS4NZ87GHHmD6bIN6MWV62QdO1/CqwY6
u9H4d//QDmwuIicO96XiwGJ+RTqrjR6UnXmV3vniGxz0THt16WbJlhk95hyj
wMikt9C9HPrlcDC1bbDsICzbcG9QLvVV12SfjcNerfYO1EzmGhAjALyUGgTn
1iTfVAoxcrRhWfdlWdbY91ZBTjdK8uZivJ0jibQuLAUCe1P+HQ+s8Q/QaDm/
NuEUdl+Qc7wbgZGdJLLQqRoeepel11gK+E2p7h/TYXoWY+S9zz/B25vQ8oJx
KpxZcZ4fcW9vv7GKbiRyDRa+PUktEDAgSsoacO/LNrswgTRmXyf+d6E0SroW
r4LxpyZgo6FFyZpEhEuDmc+hyoz0lkDh8H0VqDu7CcPKxJajjkIlFefg85gz
EkgHw942PNtL2NdrzK9NWEZjBM1WbIyJGfMy+zG/J0jYhtaVWmq2F1h6w2tN
if7ZbE68o72WVtqce3CtksVUqWIvUUo1qbatGkkFJjLOQD5ZaNBfUXsA27z6
LLfhmmI9dY5ugos9jjlVvx6MSslZLVKhCTSdcV/q+FmzILuE03VJV9ZiDkFm
5H0/0lY4VgI25GzW2qb4UNSl0c9TofQ1MZd8LuLyDK/fYvmom2qo/KntS719
wXIjpesO6ggjjTqozFWdpusc4qcv9Iucaet1dv1qryvak8V6AahE9aE2CQTs
C6To1SMYVueGdVSEZ0ATCkS4eicSoFD26b8ItVyUNve6HAPsHW1w23dy5owX
CGUQemmpGV89+g4WEGEX4NxbZ8jpyamDHxvJVSux1e9sANXY7Ms5hoWaQpWp
lD4qwcu+lVCZSyM0NuOjAxGN5XQf5+pmBXogYyXvCOm3BoqXqm3M2fIHtdlM
j80zm2I9wnTDhy5EXMYTi6MR37g3Xv0NXA4yN9V8Xh6snD+8+EL8BnMG+de1
uEggJ7kWHJWrY7HBcc+9ToBqxiTtpLAPnaIjRD5mK7FsR4aFlDNeF2FRRPca
swClKRftW9tEXBY/Gr3vJvBGKMEQ34vvcG77BGlaNNB+QLGfmlvFPE8DQzCB
YwdDdwe25IWuKcgKJKDYmVx7mjPN/Lbb81IIb+u3ZPoG9v05wUgiMIgYVA2U
c/h3KMrGiXObnqArmbF4JSGySFbuS84aN17R2GDOfvZ7MRYVi/2mvbxNQ68I
8yRZ4WQkbmrUUrjtUZmExNAKCHUZR5bKjV8MU1jpfzSuY2OmKNs/sPoYkZqc
9vqc09a+U5zQHSRtgk7hUvAoTyJYuiFLgCyVVeJNIhtwMsZEzcR6ggob+sZb
mPvrdhNQgH/WE1YSXHeU8lZoHfOcN9gUUjfbddMRM9EEFnB7fSyd8U3m2Iy3
DAGId/xmeLFjOXKJyWMb8bNRmIc5m4FU2rwfvHhgrnTbSdZP+FuCRM8gFYDQ
4GKGL5mTDswKdupOwuAmVfuz998HL5yyYYQKBVYLnN5M+dSMhBZnfmciiozi
MPQSM16fnpuKSa0CSxyEB0uJf8nQYFHGHcJPqOihtIpBkFOJSNAwhN80Oks/
WK153EClrOwQfwYwbg6Y7MWsgyDRXJGGNcbrjtA+BvWdev8rm99TS076jQMJ
h39LBpU0iWAsgnlRKwSbL2vs0H61R4cqYd4/kyDu4uY+JmE3rdtOQBKGD+RJ
JQ1gQcVpMx7Cg5uXenWAUMhwM643LqhFikp60obXiPI1+jz/ZLwsaB1wZ6dA
z6LA0cdR1+/kveh2MgVxxqLOYU8CZjUNPaOwPJiW3Rhuhbb9iBUwQRlp2SoP
u++fe/cukxYkxhK8W4D8Rrr9VhM1KbNlK39kr3i+cCHk9MIzv9r7SXhUiHqs
ei3l1OGfUtBZfnDFro9J71gmRNdfK/b9ebIE7BCRUliHwKsS9mayEsx9jEF5
HezB+XESNSz1hJySUWFfRrgAYEmrT52+jFBXwaixY3W4BO27lMscQRjEGJFv
/sOYXRx3LeBF5eEepbhPospVNzC/BL/Rb6ujB6qcOo0yfN9okyZCbbQweL8u
/LKdMMzgypEax9HdXFvkbne0eYwR8NUrFsAzsUgevQPd6t3xQzU4j7L8Z1eO
tOwOjcV5ympvzPiiwTc5+z3lzUo3CZmE8uUmcldms49w2HtOBqzS8RyYZf1c
eJoib3kMauXGHVX+tANa+BGWGj7ta06zT5iaBtQbNFuddNgS6YTr8X5nZmTf
WbGln+FP0DUfBvMMqLZUBteYgVPiwF4K8fpngRzH0rf5pFL0QSPHZB+mwL0A
+iZSV7n3SQQQk+FPJ+lnmgr1Mw2Y5r63V4j7a3MJ1jv/FiIMUYQRhnbPNfKS
Ed4unL9oZQJ98rxyzp0TanJhgrp2CzB2ZbZmogyMQ8F1izTJHB8QB+DWpBR7
dihMVpBXeQhnG+iDSgfAgo8dGcCY8nh/GhCVsiQ3hYnJmYcDp+oC2R2VutMz
zWHA61zLxAMLbVgixa5yJYyvJ6J974EYeBSJMOHQXOfVaHPiufZclCdvFnr4
EArS8UJ5b0ZWm5D1OzlzytM8M/Q4PoQ9gzmYQYXvoRhZ2Rnl4ErGamvj46me
KdgVVxsG0P07HSVhTRnS19CQrG9L1QGWnhIuOFM3tT+wxxRQClclKwdNkbVY
hA/gy3vtZFDEpD4N/cKxMwNPne9kxxEGFYXwi5g03Z/BxLSnFz2yhX6WdPPI
x/QJmGWzNY6fhP4cYCowc5XDXbALRCR0oMGhqhg5+dmzmbXoFnneXXIXekcQ
doMFDzg04nlSaWoLkN27bZvI+QI/scM7gNUdpLtawGuPGbHhRMqBUP2j6elK
bTjwHSNk9vkoL2ikMYGNaCRI1piO0fKPauajWUn65PyCRPxAgJ+mlJsktE+Q
43ht5j9d8nXnwYEfZZHZhx9YXvYHSiiLqmuegRgp7zJOPR0mMBxtqN+NXLlV
oW2cW54TSke3GtPBFcH/8LPeozo5DHuSlGb+HwNmysiph9AgC8qkpj8unWtT
s+xzFb5mx2JtN7Bz4k91q2M1wI0e1Cqcm43mZmlhFgzMm7XYsaYzAFwbCWVT
gkdPn18JB+Rmdp05NgCuB6x5tGex6z0JVGmITGJl31WuRADLMgHNAWAhmJ3I
z46+3EkYiCMt4ifD5F0VL4vKONnESSAH4PskLY975uWaWmrBi2uPvrjECD8a
+enMtqAIzp+/kaj3BLup9GEqsnhonDNOihODGjpfM48t9tkGxK83bew/IieC
zq/8yfcK75s3MaBFMPZkuQaE/uCv3gYKzFlkhyTFfirjBmKaECxpov5+Lszr
MP2Nqhc9dgH1TYk3OV4OLurJxUocDjEI6B4WzfW3+53YPFQjDZ+lH0SRs+si
FWmPtd67ANy85Adz+dib6tf550lQusLk0miwigSTq2y0l6AuNA5Pl5UcKNH2
+AZqxpd6A0YYUV9PSxwM+Ka/hQU/tCiaIwx650JxvxUIUmFU0KZaqQCKwpQo
Cypk1mNc5z+U14h6eyqFeJ5NfuxIqiF9cKPnXBbbIMkGKOP7OkDOJP/3FgXV
xipeI3kX8E6W7h8Sf8NuKBBRxIC/OvDJl8IfilDd88t2sxB/ayNPr0s7Yd2X
aeft6L74h/CFezLpglHKlirzqP4ItCLUwFNwZZjG7+yquYDP3ehYEP5nokQq
Qm8wDwFHKKiFGQ+s57r9I+NVdnjc1uobKoA95pUyAcjEbDzfMRHLgnkzvDtg
0hjDXFOjP2fFptkk+WNcblPafzCBFUMWrqeqirdCWqb6U/t3FimaZrTuTSlt
VlxmKQ678iKMImCHtUpccVBlcuYpM43Tv/vNXyiE1a7oUoOwNCqUuWSHq+1n
Fnz00dI2rABOE0VE7Y+lkyU37VRFObEga3f/Yg2I43bhfxM7f/w97a7pIDRh
/9PrXWqLh1puPqN545WRhM33gH3SCMcBlMj40K1hWtVvPD49yJ8GPFkxikF7
fg9CoKgM1uzKz/wP2XljapdBFTrPJV9UPeExRwkirWFIZgjkfAOxNcF8ts28
uhOvB28OLBZqHDZiGkV9BOCaiWnQiGyl9Ll8pgWwskAZ+GZ6kC5dDUE0MkI3
yFrorbgzVwafNkQ6BgpTUsNpX4C+31wKQEga6TbtG4UE74bWmoOgLUjMV7H/
LyjiqJvOcY04rK07Dis8UYBLNcmn55GBKVMqt4xY6iu7s1+e5hTDpbLkUYjl
a69kSuotBKYso3lB9jmAvRiCxBJfkLL91i9oIDVZh8y1wZ+a0siGDpbqj9uM
1samF1BmYdLab0r6U7vmKXFr7zPxzmahq+TH0rJwa8yV07wokkVVjMwQZ/ZO
WZ8hkL2GRsRbe5YELCc59lNZtG3bp03MSxbxffG+tixLkozPjDM08p9h1oFd
CrYH5pw6Ksgskm9ALMuDfBSCTWwXIGzSHXAC1KB6fLcZBuu6UVTDvkvH6hHm
kgftz5/0qT1HQ7qKHw5+ptEuqiF4zdZF4WS2VNk22fQBINeiDsevVjdK3TLX
Bvrb0ipEyvfF66LzQiJuYiwbRjgWQtNb7FdNbdAhvtrBaBLaRQT2j10Gfmmf
erK633h4869HMXu+60PEjI5VxF+PUh/34UpJX+0RLhUPeBEpTmXjckdI0dxT
YZrQYd1MH7ihWpEMLSRdaNw+GpNBQc9bssR2wSY7XvSg0AuInV66pJ3Ef2I/
C0XaVd/Q1xSzo+x1QEH9OA/Wc/sT/Fr12U8MoM5endb4KnN4IbQ7BueeMZVH
8Ra4gkB21aKfZQDAtUkQQgwWHDqbv8ELgesGSXLSJ6xTgmOL7hi4KrbJvDwi
5ABOT0PqCMNHjto9ERzcQAKrEYWOuDXkAyD9DH3Sy2cgmyDzlEdLxa02Mv0w
eHAMmr6nUS+LeGWmVsWxs0Zkk9rL2ZHDJtdgMAuO5Rt6OGns/GKwuInyeB0y
3Uv8fAY0UmR32C009t9+l7jAaLFBtuh32sO/yFwqW9oBvnukS1h7QKXHCV9u
CqzknHXjyS1LrKNup2tdJkQ+JpvxbQ1xeq8DnasnKIR0Usk8wk3B51zOOyjX
tupK+BoRGxB5qQdhsJGTbLZpFERXcn0sd5p4JOTD1pRv83VdcSPB0XQd/SBX
HO7eXN9Wol3njl8pKkyur6IvoPC2tqLo7I3949AX4KeqPRIvP1KXfNB/PslC
+ddlggUioEmvOHHaf/BvaXgm2YFQ28pV9+3LlFkJaQF7R+T1mBfpEQYLw/g8
rXyVM/1qABD0hpSJyUxGKFvvZzY58oqB8ivhuUTjKOEnnsnkwTFLKtpGInC0
+WmGmb0j8CT8RwNTIy+YoGas1ove1N2KAoUsrLoTIUEP4ByEekmSl42qzYxb
aHZfrkEjHrCP1WPF+LFqtKPxVkaTqwpRixmIsyl3GVfT4xNt7SpuFFmZWQFg
Z7DwJ5TIUN8r30b+T5y4EuZL5E7DH+pph6cm4v3wSbqW3WbnWkutsHGaiQ72
Yy2LCGWP8fADpagj1f+NePvhlYV+NYv3drVUDwtCfHDY95vHbtMGfNSwByf0
k/qfNhhChl1X3sahoyimR9rKwURQ+NYU0vkE47+5Qbi43n50GYBeUMCSTpPj
gydhcM5DcuoDFMhE0nLpJ9yk1479B1EWw4yJTSHwspGBsceWLuYr3kzfDlZm
4y9J/naRD3+z2LdLopFnDcbZeuoFaRxcUQQ8XdQUtWbSL4NwVvZyjnOBDZZH
w7gIUBwQvA3Q+ibOBiO8cKOEVqGT3kyyMex6/XipfcntZkltFcwYC0owXDZN
ETHWtcNGn6oK7gPvNCSKY+yUTFc+6Fq1prmDcgvcH/ms3YjhHi1Gxv4UQO6k
gaH5rlVWTvZggxE62kpR0Fz5tQaRc7Yq8tLHwXzAUUZsmTp7SrTPOzL2S0E0
z2OxvRkl2UkXFsd3YXum/oOhSUQaWGkyxzgN+MPCl3chqJIJJTaN+Fd6j9i3
nclBEQdlD+aoMWthv+T8EeCJphd0eE9CEl2sVzB7ORBqEhJyb6YuwjA8BcHv
T2aZ8W34WfsL0zZnHvwBoGIHgwJurq847gwzS/RzXMv5s6gUTibuq30+h2cD
WX0Y+kseGEmlgUgDrdhmnYwDNGrdcTRmlIqrDN/uUYrmC7ROrHMEUvQijQgh
Ak9IZa127q+BarM/puuY57kX7F+UY/50hLnMg8ALojz/r88HMaj4P0X0aAej
ODmj4Oiz92rRtx3q5kHJbipsLu/U+H4H83ovigPhpadkQ0rb4SAYcd5FOOTC
6al+T8Z0HsTM8HoHgpaZqSjCXLtieawAoeU+oq6MXw9uBVdujJ/3HoGYVeUj
IajxYK7qy812nVbrOJrla33zS4os7FaMgueApEu16YNHOEu88wLgL4f9VOFg
9p2bYOhL/Rho6RTZF5/1FiFtlQd2dwEZiID2EoH9KU3aXLoZXq9PHkFkszwG
MMqesJ/alFleu9qyxFMFRuw69WiYO3oRx3cI0n8DjyPEqkmrUYCQRNt1CPhO
VY0Ud+ly0WRPBDu0hrVqSXPj82WztYNOaJQrPw5iZ4XhJAXkL1pgdOnX6PVh
dIbyRxU6cDMsn0I2dx4LDuNg9XV1q4pQXNrT2/BE0i6rk3I+AKjBFNanBRIh
jvRsr3uth7AGp+DTSiSLVCTTkT2uw69xlnmDeE7ZHblDk1GqWu6jKDgIkGRh
7f8HjUp0MxD+CcuDW2ojuszZW9InoAzB9UVhDithnRiMSc0t9U3WgmjMHair
bA8hF7G3ItdChaOE04B3km1uoxzRBYH24MdOIVz2mM/LWkUgJDXRZ2heCrBi
uwfNm2091MWQbBIpnCbki2I1YXewGojfnyD89QBedBGon5oUWPRIMCtmwqKW
fvwGA2WlQzkUwMvpawvrpqcRUcBXVT0cDiTc6881Xl7ZVhjQMT9UTka8EgmO
pk7UfbuyrSqGCm+4zAutDsumSlLeU8AR9F9sN/0Ucqr325LanNWDr42dbTNJ
QecF3DC3nfsNo/GjYJ69m+m5x7lSkdVr5Z1TQLdhuEWlYlw9vP7zoeq6edm0
FZrPCQ388CLgLjmHnxXYSB2x/UB0ikloHRoeL+Dy83xV5IqffWI/2sBi+/fx
3jvx0kthonO1JBbcmjwaGV0LdV7O/GHZcpFj1BNTTLctR/OsnrTTFHgylLtS
4Tnh4Sq76tL7P1cMwowFHJrov8zojYk3+7/e69D7l/vQE6Sz/NiWi1FTI8wj
/CRFcaYaLT4Ls+gxUpEP1Gvrc4BBtuC/A8ZVsnOHAOGcUFK8vpYtgtzrOwoA
HeYac4sSDwISlrpbVqII3zdK4V1vOFdBTPquBIiWZ5NzjU0pBROpUTGxurDj
bebn+lW7ppA5hMxfMzyV07iEI8xH1HAyV93bggZQh1C+AfQ24iKkWOeku6tM
nFuRrU7+2J/8wkV2nDXwwJP1+OHFr7M9voNIIzlg/brhHfAleQYoVHnGqqTC
AJGwmkApa9krmgSc0xs1OW/4rC/PYQDj7oqE7lIwdGEmlbOP7Y5Eit1ZriP0
4aiaeX1jblAW7DT4gigf2JoII8pHB4YrtYTtk7tRUNM6Rq9qeJr8N0KdbaY5
Js16jwZGDPrb20dzKZAJwj1HUXPHuHp5hw1jkQE7gvca2LcH4sP5hq2ZVgy7
8TwOCvZAPrvL5NmBkQUHe8bYfhMhYDaZfApGX55ZpfeB1NWYikA4c6CgauTy
p12Q7CuY8fpEPRgIZ455r9WyPJLgY3/y4/jUs8EoplmPcAriwgYLybn1GerN
SiSwrnSCuDix35jUHt/hZRmwFLj6sLcG6/4Qao4A7l0o+yWvAh3bYkPvWZNl
ADSBbYKWLeu4rQvlRb9adTlfGWolxc/UpZoBH/LwKGHUTFVr2FYTllXYPuxQ
UzUFc+j+P61BMV1roz6PmyeVmhSQTzO3ZH3dSgIcitewnqRAEIrOLUR29JMh
2U0H1mdM/qT6caixsNqnOr2/Qt81umaBaWpDzzgR6HjGh32zlacvQh/jHzWI
2HQ9KtbDHe/K/wBQcSK3hKCi+joxasMeMokGyM1Um9Xyoae6WHsRQCafBHWL
oEiOnlO+aI67Fg9uyUSSHYcxLnRWF8OtyHDxZZAFRhBUh7YZQtjYi7jqZ4LZ
fp3H4QoFYLWt6uziIhsjpwI+P+KnGKOExZ3Ay6fsKqmekXRggQf5Uq+UGH7N
OTuRlf8SwPno/0W5DF3udw4/4WfNkDRfvZtjvJti8/mJxej780n5HmrxH/d3
O9txqD5zaanMdXWe6Vnhrs/vOXbmBxszb6XBIVQ78bt+qpecbAe3Bw+uuZcm
IlZ7iMppG8nnVoDQiwbMElNlM5QfIHHcI9fCX3EQXzVuwjVr10CZSPZJVWZ5
wYBclkLeDPMXlYADJ+P0M0xZW+FdpHEn17+xmysySWmaqDBsFnWtPGbZMIuR
aOvVs/5I+PexFf1ScdswQiOt0EgG9n4DB6fRiFyuRh3WhSuOFTb9vLXE0Lbc
stY5wXXI1CetQVpXoh+YbJi5kcvxkdYrw+eXWAtIZkgi9FODTKtdBWdxJVhl
UL1X7fu6XMIWapbrVpluH3ayULFLlW508ACpHxYLNueld06fCdhrobFcJBNe
xAV1M9rSEolrAQhHx0mpoCWdxKrwUUWOEX+HtKIUTl9sauwaKBWyg5i96uEb
piyWv/hZNxV/cDC4GdtIGUK4v1+chcH3WlNUGgQk7DLnZL3rxgB5GclIPHD8
952C7hefrpr3ojMPRFoeifzJbK1KnEuN0Rt0l/h4/sBRn6r2y4/o+GIzhQry
Oiq3BR9w6r+Q7jptXQx8DgG6UkLuVCWEAEUBqEG3fL8Nu0EPNY7lj1A6+2y2
wF3Qbs6SK7V7UBYOQ9bmVtdNT0o63OmlSMCXmQPfb8dUjOpedNafX+oYfLyf
0z1SFOnE/3phs8LCWiQPNuqWK5GaUW+tOOIc+Xn+0IZP8QlaN70Z1fhVQ21N
gxgK6I3cD4uEHu5oMD3+p/LuVvjYhnTTy0VzoX1Ru4hpGaWqMmTK9PP3EZeA
+hKT25QYek0IZW5LdmEIlcEkMNYacr7BFJ7Xy5oTRDHD2B9IfiXHLnr27nMN
bo027Lkb0I5VIfM213Lbbe+/jVPCEb5Tgv9EzBISOG/A4lTgcBQrKcRFtkCu
7P0qOZkyGbNZWXKtE2SFMatHW8vGtkMJVkum1+N874o8O6be1P/w+R6baL5I
KiIm5mW2zF9fiSDY+1Ws/Xe37SAWLVI15aFxs0718+/LyG40m50NuqyvjJpe
xSpfTPPF4TlPF0nyOIk/MUqgPnSSGaQKrblhr1zsi+xEdEj7vBxIq8lKdZxi
A7IjatWy0PONJ4ZFSu88mCHwvngPjVywYFseHIVejI2M/aTkIAUCG/FX2DXK
pOuaz+u0t4dAsCrsoO+nafXYCRm/SWFjk4oK7hT/bCgsZbq6Ualdv5gYWHcP
5Px/6Wq9htAr7OtMIBtYS2f/MiH/WkinR8R2Rqb4UEW3wQzl0XUNMSvhIp/R
vo+dOZVGSIbg7zieZ3HNPno6RrLprVUM8qWtKS7VmMPLeiz2wugWaXtCutIg
etyom8H5s13gRyIJLij+/hjptq39yJ5cQuVSaUHgED4+eZ5/GTgDbWQLRfh2
xUVKdlwhil/4YVLoBDJyWOVFI50pgsn9MRtwJQsCuNnFLh6OQS023RRtG2FA
AvHpyCcpSpecXriEUnPjHm40pU+tCyf+JcIVfrg8n7uf5kS09HD/W/1SiW/y
tAqZCHtf1Er1KwF5gOkFcvDAY7vK4myIMoMDhPalXASWpCb5uUwLufyJFXCt
9IPU7qdMOdKytbYADtEPHM99dcT/8logEmFvFWBOvwEB6P6dgD5ve0ylXiJS
jmyhFDXXjg69xJC9ri25WdGBZ2/QgqG7IBk8CRjd00lPCog/lIbHDbfPOzOZ
nJ902Sac3pEgWsOypNiyKNvugVHGM9Trm1uAzQZBrgO/LAZ7y0KiwQJkeFDt
HegRP98rFcgtJIMUmdmUNdrpdNnGk1ZQjdXaRrHckeWaq1RJ6xdE4A38ep4i
xbPRxoQsOh8lIIxN2vJ5KuEeuDXfjqL06uuW1QQerJjZaJtuDD+42WTdVeEi
Fe3fHO+KVK5FxpvztJ1LQm7LNU8Rc7P3QYU1ak4PD/aW8cl+bS8nmBtkc1cb
Ii38KrukVYpfzMNBeHJ+ny94UupnM9XELsS6R+U8LEGvt1OchJuGUPpU5cHG
PgBzodUt6LriemQRV1ZHh4XHfsN3ITEY9ehyCJ1OT2DJ4LGyUc8YHTTAeyfu
F9USmXmFFZ/292vLPpyyIG8rHVqg22g7If8TW8AZg8ajERsvKflEB1efMPUu
eKyHsgMzH0ZRjxKGCOzypTIuU/pnksGqI6W3JlQYzzchL505+j3pPVbPMcw0
F2C17aWNZ8Dovt9Qi6AwT/TFXjNRkp8TmdGmeNhdhJdk9zBL1Jr0gB8Lwk28
ldL5hUxuCZbyKWBs9hTURlPS2MxIZHKKg1l+5YiXx5z0yFDywmiRLDZ9Tolw
ia7TnZz4sJSSyw8I2PmKzXlG3BGRsnoDwv/vASnCP+slbu9pLUcA1mURvkQ0
bXPyvwAkGiCg95Z3wlv0Rqwib7HFY+QO3LK8bzRJNkkvZwY5FEdQ1UcKOLZo
atKYLuVGpvTLu5UCIpF3qeBx5vkoIL3tpDfG8PXo+SG8e/XgM7WfXOQumaU9
XoBqSevjBiA8CAJ1yJzZla8HdH5f1NrB0So0eXYw7MTooyvL9sadFPe4T/yn
jWlIZY+AR7vIACGUghRhdy1+gIJm40a/8vv07NrK4poDcuBgqEMn8EeHIDBv
XQXorWBEGhBpyyio6tqwqiWRr6p4rZiaNLQ+xR91oEjUYRVaQ4G044uVonwT
KYIg1hOxhTm1PHEEJg1XQbSrjBrqGH9VzDVbqVyVeGOC3DKj/5CRt85GcRHT
Hc7l2kr5lZhkn2aW1sC41s6eFJkmor/KzI8E7ObkWPnb1m846gTquax33oSG
LZ+8KP4GhN51D3j3DotW2FV8geflyv58asVHXI+gQbtDraTDGUCGqk59oKSq
KLzg2T4neTtlTrNCCk1o2J4OlpDq7yxxEkA82/X/PO62ioIKpWNZRDXx4f2H
gvyIi/0NmQHoXm2GeonLCVM9SH7P6CAsJqmKpOs2eCIDYnSW7huPEkHEvAbJ
u2KPkbtSroxvyRBLmelc9YCzHOsf26aEXET+fd4Cjb8P6tDKlc5fqq0XswdG
AJmSUZTUAaeSIVVmbytUkEGoMh1q+0eS9VOaVrQletMCATk+JQ6nBPLCWE6b
ydd51T0vhx5VsOtc8SbylCIrsX9MAFzqKIRzFkffTKIWHc2Ez5GBawdDT7qD
o7YQpKRkTv0c2DVJ0PF+UxoFhnDT6Iq0X8I5RreOptKLJ3x37FuKQmso6GnT
ui1jty+Y98yfUapmMhaniZ516lHZqxsrwO9l73LIRBGCFX5avsP8R/GWIbKn
6ayEQPEKDdSUHxaceVNCB4PbFIpqfWOq3NBJ1Nl6A96pY042GqJsgeEz8aLs
bQjNagTkPperH4EnsmwgWJyqmtWMFyva8k/vahxDQJJgc20mTIFcA2JWvIK1
+O0qpYcSra9KyVe5rYwtFYA5hv0yFL3OsbCkQaPiqnKs5djHpLKERJqBi6vN
RMdtkIClQVXXL5R/y9yOFA3R+qqQDxAOdrKIQJc3TbUWGbDczvDPIOPCWGOE
oCmjU7086zVABNvqrmyGlEm58d1cO78hAs9ps4MS69XpvRq3EZruyWyVviac
vF/zkE23rq9yKw/Jhun8Yh+sJIDBBoOeIoUhah/nCe7kEcAiTdg6EU1zswYp
t5RiFQC+k5OyjHTlVjfGAhFJzQXaGM9mFP4Qia3YXpsubqoXZ3aUnQOkPv8/
+JhjrjHnar/ZbHod9GbiipNsVwVoWYyHBzTq1hDYMS9R0i2hScZXe2HUZ0d9
T/9HV4S2f7rsCSPd7WUypT54FWJoZLny44/mWnxqlJ/PyhpCIGFUgU3ABO5O
FyQYCUi+LrKoh3+wWuTzDXZgBnnAk6YVP9HWXSlwKsTHeAmXA68evaf6Phed
zd8v/6SGb4TRpYmxgiM6WfrmCMYmUPDWlF9GvlUIjCt2TqUfn8wxQgjzRr6z
CEKqzssU2def1NaZGx5MWZDz1vptHNYaD8gMVOTYCtm4KQm+Yn/Wu//iPGd8
DAA7tMCCQzP9Gh9yoHKk6UE5GmigS3TIj/94Dc5slibDROevYK8qtHW+HIrL
TJaD2TRwYEV0cEWkVZbhsWmW0VZB2Lww2J8rFOZKvGXbzg10UXBDonfG8Ird
KB1cERTOoQHaNseYqdMGTnDycvYJYH4NiuAPON8nuzVWU3y0HhuEYz4wvY09
DnuRQa04oF0oSg+sl5IX5K26pSxE0KEyRS1tZfr6imekuLyyhqBYQ4/uDnIc
2wbv5wm5+9PFzSNGF49ezlVE/G0kjWCtvgj+Il9+iu2jw+Cw9J1S/N0RGWxg
1mKdNRSHUhfJ4MhTkAGLbmplz6sg2Xox16MPEOVwxt/m8bevicZ/l/uZytrI
jfkRhV3w38KNo0m/M/ndPllTc6CX7MeoVCgOgHLNj8B0WWFQ9Uoa+P6Mvj1J
wbWaS6rcVGDmA0Mlkaasm951b+f+I5mPaZ4ztYO3fqYWOEUAZ5yff7vZ9KpG
CwJjFaPANMJnwOstds+rZZ3UG1eZWa5S9RGZnqAuY9V5ZJiiXSX0JzUtyBAb
DGZpLPLrSL8UOlci/vspbsP2IImJAxOl4qxGGKMc2tBL8dF8HXRLZnSRQW6G
DPCn9vmtTc0BKgvFAz1PI6lo3OCQgiutiy6AbABGiDHjZzaDYbO+n//5cZR1
z8ysanJcT54LFVw7qKY0/1JC8ZhGvy6AspllV0U9+/b3z1MlvHohgAN2ucon
wlFrutxM6ZrgG+DjLVoQl1iKVFGul//NKPrRkHuwS8u8SX8Z2vTFQeyEGpIM
lbFgk40jxDga3Zsu9Mchb8kI75wE7thAfnGTOnDdR3zgi6CA9/yInlOD+Aa+
qPbhfMCcVJuj4BMQPO7ZKmujNoLZusqMlnmG379EIfGNP2clgPzMnjhpopkx
3sbRieFvffeMnZzwL+7vNHW0/J7Nf8IVWKVUABhGW6XkgwsNIVwyT4P2tZ/i
xfjBWRI6V97oC5NIoXGkFt6i7eFWGp8c+LFh/60KJQLvfV8OG91zDBJue59S
pauuehbKAC3cUrQOXiLXQFMcEHdI1VV+PKnBBQZpTh18nHQa4x+LaAZtWImM
54SUtIQPTUJKZBeYwFoieMDafTTCon4RhHufvHakmSRaLE+h4aOoiTUlM5gv
c63kcJxu/eEocWSj4Ix3tDY/ySgv9+XPWD+Tig5E0iF7p4mIZfveiCKBqJyf
8O9+UY31huT+FmQpytrvExLaQMxan/ToccJDjTeLqbXnZwEJjQ9gTtIa4cL5
ChI7GfbUYBolm4Mo98mnkVlD7LpDJNoEY13Co7qXcBcyTqS3NVSY2q1ptgVy
5MyF4evBuJ6BSyLNKhYVSxUo5gBMEVkIXGiqDeRwuKECToMXNVmplcAi6GFs
Z4jAZJXcoB6mIkR7ud5HWcyT0aDLI3gRG9M8/4Ic7P8V2SH2l7HAkCVjC+Sm
bhf2i7fDVn5b9uxuKWrPyd7hG6gWl9Os63hEDinxCObvQVWi/TAzX2ZvWMRk
Z65xagPJnwE42D6sz7LSOCVWnuIAK0nwfEc7dMsd8hG2JOLcr9KnOIVldvIc
Z4UIIuedCIzKVKj8ItK3CUz527f7NqV5RaBEhnBM4/t5k0LDyJK/wc4xGZ7y
p3YdXfUi42e60jBrbyATg5BuXbfv/AqYF4Xjeb4/HfSz2nyBwAY2OGdtQHtH
GpKtTa3Lc0YUE5RloiDhTlOlIC7r0MnJ2F4MaLln52N3q5AqnZ2GZWqO37/Q
RdZJDxw29Dl2pU7ZGVsFMAQ259+7SujPDHB81VtDOrF2yQmyaIcq+JMO1Uek
3J2oH5H1YetyFtP19qmIWlaNC0xUc7U7sLJIMXdGya6u3NQZKeXDGwdK45QE
n3VZn3yZD2on7xj79vFjMg3ZYb8jZb3J5RlO7rs3uZR4CymQX3rC6IsGkUsg
4AwFaeZuPYZVt1Jm5hl2dFhCCl0a1hffixbzciu2GF1wkxmfYGWGcgTtJGna
rpqD3+pnLu8G1NbZCbcRC1KQk1SCAtRhHPq1KskVPqrpsaUBMOsMrndSZVKa
wH2nSXKaFz4hduE5HFI9Z8zmU/EWq2V/DfW27zU0x332SjCUl8epJlkos/Us
PMDCuyxq2Xw7tQtU7YgJehTjQY1pQNkLT/iK6J/uL1w63On6xkvuQGsNhpo6
GgJq7YY/NaPw/EMXxVWHTpSBuLt9yFcBEgSYRsoG8zW6rcmIZbg2Ys501NWC
pQDfVG+CUYhO5H6k1YYMFT6vhVICpKzWfNXJylSxJ2swX7bdFRZB73cQ8n4C
YzvkhEsfwzGuWEFNxCZpYCbSqpfyQ6kziUtmyFXVrjAt8Km2fVfxFu9azQUq
XIld7q/CgOiH0rjYH/BMGl+V4ChQoqTpjc78HE6mZn7uYwFC4LM05zxb6NyV
Vr1PA6AjfsVCSjdnXzft+t+afRmoWpswM2l/qTQOnlSpV8/RRQ9po3pAup9P
NoYht5CknfVgcRdqe0MqdDwaBMJ3YQI6HFhbPphD/IxGF2gmfeXMXJAvnFg3
R2kKuaxXrEUop/uOQ4GZgF6OsbfG08wvUzD2nccEksANCXj49vjd+WUEv/2R
q9JHXzpiq9r1wOZtqfa8FMmUz/OMft6JJQdT7oi0yhCcqGvARzB7ohsZ/CAe
qAfVb9IR+vCcHRHGDI27LK0NiP3vmdA9vAsiGwO/ykwW9Mw0dM7/uqAn/5MC
ClO9XOWTLF7KifyZ+eKkiu03VJ/JV+smoV+9LMklnD9ZJRCjIebKh+YrM6iL
FXHQKmlCnKtpp64e1hHmMc+Rq/uGiCJO5Ko8Qcs/tI0IuPijBxzF2Ih1ai2M
8BdzNKOdsS3jubl5mKqFa9B5jkxSCqTSW0z5PoXUf/7troNZWCEX2esDkcjW
2FBzxh32BlJ61skRVztOFOcFT4iEVlLErVcWql3ATh2PfEoB/Q4x3x3I+Qi9
pt708/h/CLYpil59jY+7z0oTryz4e+G30NqLtlWDD76UhPU27XZl5bT+KObK
aigWoaAOUq+P6fYgY8Y6otBxvLH+QLq8V4EJ7aIKbRYVfeAP6uF87TuibIMc
VSpMED3/NAkO1A2chXLQ1R6me2HNM/IapIudw2H7D5vVN6NRPTyeYeX/z14S
D5ev0YpHEe8gZ4Yu1aiukNni5/Ht8/KUZAvImjGxUq+Aq/wy46YWerI4NTYf
WTpggFHGGZI6BRF3dlyPQc8OzufInLaJAM3Q3hjhMnEEQh+Tg0a6QfrGb+0v
QVTlHyVyeEiHp9CGq3gvkHQAJuEw9o4ltXgGOQ5jUNjt4y+P+ee13TmEBZHg
wC54OTJGMdGOF36lf3KNV3lvge1txo8+RZZdkqP8+PNqCGYNOCgMNpc6end/
CZS8RRznI7nj9g4x78EaEcBsMEpuaIcVLxCIpVxqNZOGtRN7t2o+ZU7o7QAz
4W0wjaL+AI+9/NC2+akrRa2VGM/CASf4w/5+O3m4beY3YbyHhBEl9RcOlVuM
8pusChCzXic8QVpLnE6x/kn4M/u8OUGMOCdQ4EdkWLraUisWaR40SRfFtz2i
hSQfRX7jmyvIgSlG9kBXk4XIOdYo0o5KTQlJss+A9BEPltexlZXNdJqR1Ktc
61OeF6espYvpiyjoUBZzTfp87KxO3/eP+/lsjpsv5SRnh6MUVsXPjDTYZE9q
FHkeRSqOnTq4UXjoae60gXVOC+Imd034nFxR3gYGKXR1oGIf7koX+Rc/DvYU
fQjN9iYICI9dAEA7VZ6pWdSmLx6JRQS/ePcyQiDGCD0C0MjqaaTgQ9oOOBFi
KdbSqf6fP2mbO4lKo/ytxiMNgk3qcfYByZAXJ38Pp06Pj7w31rWP+X7XTwZ/
ozVqmyTb5rXxWCnEbhbC839sUfbHb8oqkJv9ae2UjAaeNBx+ijXUItZTJ5du
IAhahP0nugPuGudWoJT5BA3sbRfpZpwYRm8Et1IHBDq6ufEJVrBfwoXMdb1B
7ssaSGHrl5if1Dgeaz/0hRFWKx6Qz7IeEhOhtBtIr+GL7El1gfizPrhmxyWR
Tlp1jxjlyiHQhmDihsnkoulI6/GBvC0WByTeX9nZoPrBgAHPDZEiJ0xGfuSZ
uk/yRVUto0lLJ0Ov1Zro3ntXHAWupb4LWWGLr+yUdcEdtLVXGQ4JVZFLCiBe
MRgj3rRZahs9adGkKjLR3x1nqXHslY3lxgQ25GC9Kl2fKlu07VhrSgq4PR4z
Qj0JDK7qemkMYnPBPf/Ky6UZHsPgmC28r6Z1mKVb6jx58tYNJ9eakvGhwXg1
459TxPBfvRPtEFHadhuUSgp4YOLn5ZPncDHav5JNh1HOp1G6XUWhojsP4PBW
Iv7kPGIvdjZMkT1jNgy9IG9285APDI7M1ZAgBqaVcoyOiu4AaOS8SpGPSr2Q
OsW7B0pJ5cjS/vpeiOeGTZ9cUlMBzFRA0JvC1Bb1Ziz91M5YfKzg0gZ6lE0X
wrHmFtnj4rnKFe6+hLSefsGBTkskTmiWrnF+hbcQV8KDX59eIAFnTmd7Rgva
SUFt+nxOrif28ze352WD8jrvxLJW/i40l2MFwdYc8ESAOD/bHoTtoM0B4leU
qgJbsIZMJAp3fJqDJlF+m+Ug1aY0NnizsXC9I1BMtZVjEkLS21JJouO/gpHj
/vS3I+9ssMiJ9/LH3lU3EiOLo/9hGKZ7mYCvfUlv1WzQZWfbwzfJunyp0onF
ItaA8+2o6H1PHxytbDknOB3UvZ0/GcYv5HmYiom4MWqxvYc6Z4SGBQjvHDkz
S9idEoeAX/K3Tg2jWZiT2aG9TC/Lg6MfCFilTwWZA7wbJ89/rvMTjdx1VF14
Sbn2ok2p8tvECTBffgrMHamEU9clgCe8ARA3cEiAfb1aT6dmP4jbhyxzNQZy
DwTpwaHGujK3Ptlw0iIizYSQ15YlGltMTbzDQDaEiTFB+EGoM2nznDcDHrO9
A+4MQRGLoeHWG9M4KlPcPjpqZApRfO0WfSvH0sLfidpUzzzAg4uJEHYcjoIY
wF+1ArBRTZVCOfSLaPnlgb56Fdi7TWHDxul6qWRd4tC/7O6+7jwYNU5kccaN
UU1Hu+6MqZ9SSncnHPvuusLYO6JuVJGhcvFkghvU0R2RzSuFjf8SgrtdZONF
nwfBzzEiDO2mlDWxtr2URffrOaq2mcZkr1+rd9mxVVjSjUaeJaaTAn8jHwlq
5Bz3JVK+SGX+xTRDR4O3nF6P9phDgYiiKuraQ4R/MqtG2pgjP7X8Nj+T2Ky+
smdzK8GE0juUX8bAp9dIQ0T8827LPzrnLx0ShQ16SDR/led00ApBR6G4Rny3
VBxF5dkb4UodXbiI4WgIgyeTKYwZK04qCwRuaLF+x4dgR9YeAeFowNsAMiio
e00YO4h7vId1GdHqjyRWYVUrmC+lhNVeno2l1m8E8TyXwSn22/SIQERvAAVr
6RgVr/z3sCKl9jP4x5gxs4szheBCqI5C1yCovyU/M0Dpv1RsSJVM57bcz0Qj
/OXE+bwxVCXhuXtKMWO4iK6oIU3dyLwxdtQ+C9Ljx77i+gg2THlonxG2nnFp
/6ZB5MJjKGS2E+WLcRalXOoSss7W8YfBjYfzFzL2G2U/yVB/OCaFT9TmISXu
Rr8Nuug2CEF/Zq35rze6twVEg+CcLSHBd/9vU90lQh8KzZPemd4jucQgPpIU
lt07DFH/cT/f9IUA7Th5glkGmzvrj4Dk2DlsH0s3ur5+33TB02CSivjejjLC
Q97y8iz3Bq6FLXnaTc46RyfXAeh9h0vrQ65oYTQuZQsqtbpSogO54A+/wlBg
KGifdZC241yqCLPg/pV+z9xDqXV8kWjNfze1X0Y3WBouv2VBPtXUPsXeGKRn
fhuNUXIVklliS6ocTaFN9yWFnsrN94oDw2lPKEvYX+MnuWgIyIjhcF3zZ4b7
NPwuJkOODnniz0GQ+S3ztQoPj7V2gPVvX4XuVjsr8fu+MKIlbL61NcWQJlrT
5RYQ9cBlks0+2MmA/p6qtfATW/Rciobd3GswxqG2i214fWBc/ckeXPfKRFHC
t4YEK0c0obEECHVvL7fLq3D66oS6E1NmbyUdqLxACljaIPE1V9J0invoUIfC
NpdVpfjo/2lLcb6nAtsG8a2jwBe4LH5nG5pUFfIDRKD96O6eTP7cPfczQJDi
aj40cyaS4nTpWFpiPr+DShaZ4c7O5pYVowWrTXt+eRyyynZH4ea09B0AW9hV
lm4EzsV+ZrHFCVK/LCt2R98Ww9q2eddjn/hAD36swm7acePjwbRvjA1GIbul
M1o/K8vZUsT6cCHq3YhTAYU0NOu5fE7ZdD58BA9n3ZXsFbOBWGDWSy0K4SLl
Ze5DjyabAXPyav9tRfCQVgg54wYloamqH3euP08j/1MMcbl3DYzW0aWw07qP
pecnOWj6m6JAXxneGarkmBsXcbCkvwcnK1mOwoKsvUgsQ2i0xLL07Qw8i3CK
qJweb9xhmm36IytD8d7r1YLqxbLgJiIkZNZvJGnlQVLZC0oa+d7/bEf3RFEo
QkZKVetrlkMO1fJbnsBzVVYRnL7ZrvAa8y0W2JEGQ544JH+PR+hkF9DkQR9v
Mf0BpJAViW9Ovrn3vub5O62PsRG5be03tw5lI2O2DGucMufHyRY3W6ei/JrR
aF8tF25ZM3XRqW6PqXAq+kTSe/0rXGzXms/ACpI1/RonvzTqDdaAp+UpXNmo
aBr2yZhno/0rNIC2LWSDpsJIfgVNEY5HSQwGUGTtPBG9QTR06EGgShkxpdQD
nK/TVswFAr1f5Iw9gk2n2addG20UAOy97BzfE7NQZ3UDoRFYfk4PzLQpOPHv
AEVKJlHJsKDYqTQHuranShOlySH15Va+7O58ZkwLzUxW7amnb0UFIH3X+/YS
i/lBMMese6739l+lZ4xOW8EEC3tZonzR1/e7aKUjCwkxH8aXN1+Oq4canPo2
Ev2zSjRO3ewhuScAlfjUVY8H8q7nJJfFLX5j4yC+47nQWC4Ad53nHeJ7gyH9
JqCq+VK6REydvfn9sqnVgBkh5RUm5I2rtbq6HOdN2JVgqbfk3nRpc8wn3D22
aEHAp/VpF447pDHoRmkbJAL75N/R3rCipQ/CABP2IXa9ZHZJmUz+TBV0Ylbx
WI8U1PO/chAz98mERYfSC8IrKVbbHSPZrpSm5MMBcQDmy1CKHmDGPsNjUNs9
LCtcw/XkOB2tXYDErHyEUE2W5j09zyRjMIxCkBOgxn0oCk5vsDx0MdWPm1ii
DGxM3sIy95fL0H5d/uNFl8Ut9DPWqN0fWL9uiABT+YOJ6qJYym62/rag3nmG
YhaRwYIMZnfHBwFrWN/Q3mH44QCTZ4ce9rKHBXWwcXN5istIJPQoid5RolBF
B4LnH5+BCGMa5ZvgiZqfZ/cOsUjVkBfO9kT8S9ttrCyBBhXCWHt2FCLbttcH
9QdZ68z51JJbpCdMm61iwRxgTJRWEsbOQcTclr/WQTb1T4/iAGGqvH3Ud76o
S0V+Eur8EYjXWdK9DxFjXJRdsmGT0yFTij86SghNgFJYZ282xh9IcFKX57lt
+Ugk5v2vFHOLncBbD0egtEndUFoUoWvKBpkEBmfp9gBGFiW5NaluuELU+2Rh
56vA5rUg2DelsTd7WBmRQsy0CdCenrSqYdlCCtz3+tWCrwPwhOJqqRTgHffp
zu9MusmVtRQhlCFrEH2CPme/7dsTnDv6JOAxBt+cHWAVFrssjFhpeWhKQeBZ
sZOTw6HZ9OJZkhKvLe5lO6FSBoEqj1zsz7s6TtpWPfzm+26Q0NMZeU5hKCbW
hIaEgddY2eYwYO/HSVVHR9vLtz6G393PkBLNJQXXmeZ/T9HTW2yDyCxF13Oe
nM/Z8W8QmXecXYQRuzrRYEg32UVS22C39UGnalq1Ur9goibEE1zFcVVZhuK2
oruhWVFd6Yr/PR5TBtVEaxpcj6ef6Rg+yuAzBeFEXhnVJ9KxejO2kgVSgxFL
KgHDjgNI04d+/Sw9UZO6Rim/CbZ7uvzgxPKrQP1PDU6fL7DiTnXL8eEMRTzP
ELoYrQ0zO90S7xxbR8nbDghjoECcgy0R1iaYb/PKcvC32WIE/iaNT9iXcDsa
d8ziCgZw7vaf4jBVydT0fq8sLoHULDLTzbCMGPxhDaCnlEBkqVNQ1EK8SD9+
0qs3TjRsq0Pi3udCRGOHhH1Joxq6dYGEUzECt5D9Ce1JdLQG0N2Jx0IrZdqT
RmGi7OZ8cdUak5EofKr16FcaIDsHMRuAFyFyDiB/OfCPlVfrF6QgTl8H6OJU
kYcoc9yjGg6l02Odj5Xcuq+fktrY69CM094qqpElVbs5LH3eohE84I8g01Xa
18Dgi7FTQHYsgAu5u5Z8ZevPEnk++5zsYaPMPbVmcYKkiiLjspMwV2qI9yRw
HvaLtm/X/jVuAFWC3Xl7s2Sq7Zp8poOfnPzHj2p9b+EQWqB363JSNfD8LUlt
dte7TE/2bAqq0ipyN3Q2Y3rToNyQ6/eW178rkhbi0csqqMqewOmZ97PhdZo8
dbOowjB821zhQb53iYv+PxmCxEhk9/hATm/00vXso+fTo5UlANb+0yZIBLib
dSajO+7108PPXYgWBFkrW7Lu1A5aeTvUErVl+6nEAcxz+10hIw4mtZBrqllq
h2GUFmI5kLcMTkqtN+muZzDg8pf31E8N5L2CWVtUKLj8RYSgZiKpVPPgM4ID
liiB9n29S/JYR2FH5qZ0PAR1xFBcByjbJiW8CcZq+Nueu3yaDYzqAsLNn5z4
eDW0QCoNc2KUALiPwEZetP4VptwiFsoAp5ToFhRwshYYDt7oWNxeAJFrfnyb
9Tqp1Jh3+UelzlQS0rfXT6DPsRbIZyzc8oCAAl64NEVf7nTDUqu9f6LDo/oo
vEz0Gb0KOAzHf1T1TeWxBFja1m1z9atb0BEr1Hw/U/UkegXbZttdwnrhZLKl
2soPBEFqo1NtotNq4P2ThrAAsvAjoGH6ACSMXVDRx8HaKehA/veY5XVlbCQk
mBnyGp5bEFHJ9zgRN2n6VjhX1NEP0N6cFrWsaIgESU+67j7kMRK2h8uDi25X
Qm8oyua2a1MtP1HVVWGLfXXIn/0i4XwRPk4toS7+3vh0f+tvcjr6FU4CjpXW
f7LZLUqNTN/lCXKb7z/9WNyIZRUgE4OOTmQEUjCsSAO8iD9Kl9omYTt9cv8J
uJfY+hdWjM6b7xor9Vk9jJpHpU5rJ3L6LKO3nKI5jY75VJRmAJC8PpCVkZUh
uLsQten4qTvGQxuB1v0c6lpFkV7zCatWRnUr/K7t9o7Ht1jK9xOqQr8JVtnv
RAKY3NTRQSpL7JaOCQRJKsApJMRx8pgRr6xUui9F4AdUhJJeSYO+XqFbObHK
Zx7Uur3+zzNl+VoCSMxyF4SPHdFPCg9V6EqYD1YCJ2fIfqri3frN57TdxL6x
p7fZypgFESe2wvqcF07n1vujpTEUyTGQ3eXyYKcVxyOTGattXdR0Lmt5SIij
13KEkdBpttmx3XNsyoxNODcEZBQsysVI4Cf36yHSjFPEjLpWJzPNHPl7hSGy
7gOXPe4lyEqE65cNRz2H1bMnoxWsG1gfgHr2SD8vgJZkPjZvrReGM56aBrsl
09kimm62A3+XRseG/QEzJ/a5Kfavb3xc9vY7Ng+c98uvuKLgmmemdyj4bqan
l0bZ770paq5aoI+lixUuno+1yzVqsBRbmYprdk15T9cQHwmrO4DxKzPglsYA
ih1e2yXSzAvTu6s8fZXCf4cQiJOBE6fNVyRNnavBbuqCB1b9np4SGy4j9/lB
UCV8knNQTS56l27MsD75QFXceLYMQBZB/DYPNuRLTC1u+aNFKTo042g3H10F
3ERCv80a9nqyZABcY+8wYbHwe0dxCh9UyEM8MdAusbAMRSuR+B/7oR3uWSLa
jUEql3d5AacDGr3ndHgPIL9iVDJg0vNPRJL5T5uUlhN+DPSQNUGblWJI3rxg
DN25yEPnZqt4mgRrT/skw7fuFONdeaF1hFLKitG6hu504eDXZabjKyoAIvVP
dGmmVsBYQW0mOqfzD/0sGDnHW0TAvxAN1J/zlm3keRXDJcZNBMYnfHxpdKRy
f5MEQq/0ODBqI0cG4R2NCu7lmK1Be9DDL9Ll0bNOkol+cjTseH0qYQz9BJCB
Kw4QbMOap0Q+8Jjt83Q25Hq+6Hiy+IahBPXIXn7BozENL61I1yoxhC+BnLaS
Xjd6+KDOKeuVHlGiUl5KWaHSkS2vAg/1yfZ7PB0qlvh1w1iDHxer5Aw8HR43
nVmKD76MIZLBhQRIIRYryp31zMKnnN4POwahAc8HlvKZb91f+GQS2pFFqHQj
RGaaLSMK3WzerxLlxYN/nK2Cvti5RG99Sqlgkn0fnHR1mOlcGYmJ+c6aAIR5
HcldXzujNlF0cfxAKOaMwFbMNi2zr07R90Jxz1kDHOAisfi0reotzicAqMDU
kP7uUob1gcDyaxTdyKYzbbT/+vCugTCMj8NasDS7S2r2dXO+JJ6BTMlLZwTg
epzyfDKwGgsNoulLP9vTVsE5o679q64dDR+XfP3NIe+GyRNRVd3cowt5NU30
kzQfgDBu/zGTC+Nt5ZwH/lAnEkhG2ubOpM3P8qRZxbcncFoMoY42pg+vKvy/
KDbyaMOXPL1v+/k/yH6mpdnxD8YD8pYyGb9S/XNGQZU39u7P0hmmRkwtdjXX
+QjOsODQhmkVeJsa/nYF/HrZgS4NhttD9vAE/VOlapIS8uRu9RdPlwO1k4+8
MoVArGN1vuy4vOw7CoGOrRaL567rtf5WNcjmWH2NmacUVzMFURQSRlAAEWCt
A7CCK/FfBPmMuUUIMfWI9s7SQ2wAu20EEA+HjX9AaxaOTXgR7SGYocMFbT3X
gpPEnuOOHkVsq8oHKwMzWGnchKSPa03uqp+Uk4KSRn2pyjT0LCFC9V/j0vqa
Mj2NxadSF0gHROnEPoXlQZZgT7toqG/NcATOWZm0yrlVs0BH/2vorJvBMY56
4QfHzbP42Ec9aQH67Gm2X2+/RR9/uYAmOIwDHIdR2uEr5hW5zswyfBUPJ5JG
fjv2kz7f23LhnaAn6PYzmQJFBjkZ1WGxsEzqo9fMcK+OPN2FxiIgYBovxvbo
DSymeIkLGiLIaQZNj284VlxI3FBKm+/7+ViomKBBFEcd9AXfG2p/uNfflsKn
3K6LTtux0F3RpLkSswfK2T7UQ4T8OuNMCchdPut2Qu4hQ6Dz0PU7Za6RUWzW
eaZ1S2Fbw1T8jjVx6xeOFjsz/B6wWCc+pk54b+YwPg888JRvj3fViHt4PdtT
wzrpCXKcaUwTzdfhISnTj8PItB31fpTY1EG8NrRp6E0QF4J91pFgl9hS9B1o
s85NNuCfoVv7lSxd1n44pjkMGY/UZE+LbXEe9Te7MS915wYzBZkkhJnD5a3j
DQ/whJBimYkr2MT+GW0fcy3yoYfQE5FaXsr4TlhbL4BcStlZUY9ElXBdxtRj
Yw3coy8BaRVuXAa5rJm+k/hWazXiV6GxihhgfH0q0yh/Z2+vVyBVLm91cUNh
a0hVv63+YoGnQf5AgiK35y9nsF8Bwb3g8CwGnV8rtjFqX+ogle3KfxkAiKVh
B0+M+xecwwAaa9r36Pk2LlVBlGekRcasYTN1Sd0kBCv0a5nT0cLscWMa2qRZ
e8vf9bvu+apCjuovyHRHKZTLzpeQqtXu1ULp7/uQ/gVGuf4mgqTieug5+UUm
F6f+MYmdvwBv1jiFE0QiI6FNqOB42b+pOI9xENiG1pT7N1FuBZu/xBWQzNBm
Lnt7Eye4zP4S3gLQT3GkgnLIeZgAOL6PHdC9KmeLhx7MO8T1G9AmBjtPQcHq
pv9pBVlIswfKbpqp8mZ3mGyk1jMXyjjISSErrXUcUCZkxu+Aaejd9lJITqYd
A+BNO2JKsoj5Y4pMM72l/2/qgR79OsVXUgGy1mp4SZtIbYOH82cyVtvxNRMs
zdjx9Vgo4rb6IuMMyAzKsEqo17HjP22g4qDXHUzBZzo+n8EHJDXRj9bAYUVI
rLQTF3XTZL8DxYJpF/l65IuwY55+a8LMenrZ9d+FF0KBqKnpfg2DxXI76Gg5
IWJYD8P3ElO0CA7Dh/sw1jZiL3TPpfKg5IaYxG48mNIvBb8IfjOsxJxgsRX6
C4aIPgPvRqTSaDYfyPvNt+3Tnz5Vr5n1chH1cIanH4Nvwl8NOWdjELYzgxOt
RXRBtint+UdF+k/4SOgivbhD1G2TYKsxYMmnbcGtPAdxYT+6AXQ6plJR7BnA
Aeyqpz+Gch3qh7tMABPVTtyhQpa1nMhNrM2090VU9w3f2Daj57gRpYfD3JZI
ik4+w7Ae4ZtgQDiPLkQ1TF8bbzUuO9K5dGxohumF9gqiERrwGH0wEn/2ZpKt
OwAJ0GT4yDZIufm0wJ6uwCklFa7UBNAmAlD0fi5xZq5hPHCAxmn77jmi1pRY
X5GyQ6vfMA5qvnMX1yw+FRuqTYbinbW28frx+B8vRNDvkHfAQHUE2dK9Xmpw
5h0iM/x1LhJek0Q12COpZmOhW7DRGP4bmWuawx1YzngtKy405WCE7keuY+ly
3wOCNaK4O4F3mhm9aPl93xsQvsNUIRPE4095H0BvgTmY5LENuxcIKZj7CmGs
ZTMW9AejnoYvAVbvfmtUV7hHgineV7qeLlvF8GlXKoDPIUluxphPHRdY+ZJG
0liwYD5ExcRI7LgbwtdcEHZymsLismT+KI0LujEJQf+sCKrxlXPuAil/CjiN
NREYyISvTBd6IY4MYrRnU+LKuRqgoL7Dp1hziHMY370ywc0XGYMzoMm17hKL
ZNXUTW6atDfiMztf3JzsK89WTbvFsKNJgrRAh3bgwKT07Jq4pWa3CeVc5h+a
tiV4rshWoAbL1F+IIWQ/QRQYZ5nrMxzEAukp+F8/jenXuzirPKbU1Y0Orf1z
bhfVrkK0+UlL819cuQDkNXlwcEcHkrCFpNa/wJRnnj11uT0GMvsykSd+GD7I
F548skVE0y1yu+ChP4NjH/+osU3jIztgELHHxgakA9Fw1vt4DeVljfQHHF5F
C6hEnpzFOv9MMY9X9NLYEy0WjD28fwLwJrg5DWUIt2c3osFFpJ3+K1VAWSad
4xa1e6eyMszIfziK8HMfaDHEEreH/cGQ/+x7xrLOlHVngUxEwxJGJamhNU1b
W10uj5XQB3tGztu7/2V4u/GEzX2rl7+L0h0O21PTir2YXpgXFRo+dRryPbab
tEPIwrxvhFq6YVo2C+sf3ZY2bjTIeaeMVyMvD5dQ2lkezBgXi4R1nq+MUm/R
6u0IPXJrNW6KkesX0U2sjR5rxeBsmI6t+dkLstcK42qWqAyHTN8lsIDEfRj7
u4l3fjK40lc2qpirMKyZPAvmbHJ/iGLCTFTaKVTOZNNHipve75iKNUW+eSRG
DPWvtw87XZi25My9K+CTQmeVAlH7D1vjf+HBl39K1GmMv8nWLtG2KL827yRL
5Bu2rKC2zY+R6fnlIDhvTp4GVMih/ExHeiDEpz+6eUkRhgONI2+wONfMjH5s
9YJ65ljGGyL0q7tgN5vT11HHmfg5ZtM+YVevlNNkyfKRRbSdCGLdwJyYj4j4
Sjo88demdSOChxXs7D250sOsG7kAqR73K4IiohLz0Fx4WknJU6/jP3BE+GaN
wxse/x/7tpngOv0SQ+Kj9Mq+gpvBz9GJYlxqOze6xfGD3+1SxZFd4DV7FVBP
X4sE05XWjO73p/0tLEANoaV86esVyHHPiQjn7keIu5wsHTa7a+bCeYLUuh/m
2mIGNBSQ2hqz64SgbhKTR3KlSYKOXgdXpjvIXEHl+lWR5L34zrEmc47+8HdU
jSPCFEnFfmv0ZQywn8sjHF3ScwBEsnT/3QstwDiZlBl1eME9EKLtWshPxEg8
9OCPkap0ZXv6kwxwfPonPxEHlERLRdIf/wuprgJSnwnm8wdtVBJD0pIGfbpv
AOZdJ8Hz6kCJDZU+ctKJlew9SZq4/6yfQU1iojkB9R9PuQ1DF8/PxdWgr5Qr
EvscjeiPt0MuHGCDBPTbxh5QuwkVOyAZsgvNt79KPPrwIh6uewnxioJR+mWc
zsk6tdX1ZXmeqLqO9fSyK7JRqNA8DQsXRKZEliZVTKtjc9FptanpJ1BurcDN
r0/cacgDwUpPG9tmEdQuS0A+8J9VhcuQvKs5F3I9uJFH73lEcdNCy1a4h0ZP
6yCzTq/oVuD4k6E6RUzToXZgIyExpOm4uzf+H79Gzfg8dPdr4u3Etwf7CuDx
MSSlDhiklg/6QHBPlVJyq5U7VQbLttnkjxwbNE9qodR74KqFeeCdFzuKCJlP
ufmevxcWpw9GFedJ9rGKQ5YneT8Qibb5V+TjODtF7+UXelro/hgxE6Agk8sY
pXoJrCXo/HNohdWq7bnphYP86snFR/46t+2QZQ5dWwB2ENRQM27btFn8gQM0
P1fiPWJ1N/Ovld0MQ5Xn555ZAQqYoxbrCC6jvEYCdLMLPPfFi0LIDVfMHYEM
waqt8fY71Z7wZJzlrxlq9p8TVJ42DfDnR5eMBK9i+jL8QFXyJvEmmD2tx9x7
2FC6KaKmqiriEkUeWmnN3iGHTtzUqJFHM6QguBCmgZSpYrhJg8P7M/FqfZ7v
gkxyKVFr4pVIqoqKF4pDY2abzzwMAzfuDIrpAIQ19KDThU67u54eNgm9f2MQ
lziRokvfEFb9zMb0UH6DR6Nci69diIiI0V4j3uxvZZ7imYmhMNXPyOFD4/yV
wlLIj1AqfZBjpp6Zgiu0mdexbQ1dfkm+Ib7bOmHW4oWXpwZrhoj7bo23+FP2
Hcxltg/4MIE1eWtBxh+abVHaP79j/rMf/TPaenB8La3b0cb7uJ8UZsymH4Os
5MJZ64TksHZ3jbHIYW3ouPUFEQdH9/+Mkcuy9FQzbj7/KLFpYpjMxix5jVVV
tNXF2MU/nUTRMNSYnkcKeI3LZ+EV9a4hcB/BMDaZ0Z+F5bAuD/oRNiSTN6n6
y6YxHHFvUShCnCpz3pGzrg7qDhYDdjjc9aZf4U2jns5TzmXTUTdfgZxlSCBr
Wtccx9j8KiWWT0CssYwQEtgz3X5Dye4Dhj+/ZGAzbW0xtGiEP7PDZBRP5ET+
EzPDPmxkGE9Qe/H6OO3Ksy0XB9P8PpCjnd5BkLsICthr5dGCgPlhGjWDCEdp
fVLKuLA687lcWlkXvgXNTQQQZII6wZQIkBpZVGER7l2jMOruuqKEmmMwzz6e
wvIOKC9uQLQImco+bCqftH1pPfMLx01jsmnycbdb9TqRkF63RakbEsxlmkO+
T0XgT6eelIGNOGNpAWuvWK38Hioe6USxYqWM5VKHjtKq4Bmf4LAQoVAJSBbp
YqErH0KwJE4b1287qx1geyHOk8U2iEpsSh6mW794cvH6Uxgkn1c41zd72qmB
y0F5xYaomwcs+4+OY0JKIuyvTA5YXFGruaiCfs9EicxEL+cgK8fJQhuFwnkl
p0MoYi+t5+Zs9wlo2y8kOfZoeL/BUXbpnZu7xuAiUXJVUKYcrbqhWDgD48ek
SsW9QU+ew+4DKrwt3Sr70rTgo/t9MQpNLCIJDL6wMhOSVxNzbKWoePRnspkb
cxz96i5UTRLfliAr9iL4uRQ8Yzk1nQQ97fP/AHU5WWDxJrrKri6hOV1PvMYq
FoVMLWGt8kWAy9bKPNNSuateisd3Lb62f18D/AM1kkeDRCYvvky0c4ksKsE3
vIVXgBgrMVuPPks9Ui+6kWIPJDR6/HaFuT1CkT5dnyM8fwT2P/0FdPmbWu6K
MiZiWiuBFXG7NKNIpu3zBk/n9qRn3HzVUCNjCtabj38W+f/WiOO90VJO+Vy7
1Yu/nKGis2DAVq/r6aRXsFTQwlLbjY+m39NUokOD/VcHoVa4zu7Hf92P8R4k
ZFU1LCYv0CMyhtgxVBpdUQHqBGNTMLDEanoNLPO+Pr3V7edM5zhojm6uGYSC
bErronfBHrq2IYDMxmxfx+xQDr3C76DyoRSdbZVx3G25rPUIsO+tnbT6bfLM
uOkiADN5lFP9qsWUqiOWmtw8fOXpOtfG+ZCkiVRffat+m9uvqjceWIfJlqDk
WWbLatorQHAApm55tj391JCkmltlliINoM6Thv3O1+tGe6Uf2R+zrO8WZXIY
5Ece0f4EhFxDaxZa5gh2i9uNpFNj+yZICzGwcWF1Ey0+VKliMvg4TMItSo4r
V+uvsMQsWoAabwjpfMyZy6dpF8P66rhm4QCmZ2X5Hel320FlcwdlzSBsCnRX
86VksdFpXzTcIT+JsS2g1xNxA5eV9YBSec7OcAIpmYMHECM3VwAZ1LNocRui
8Rcrjb2KRIp9Pcvx4XrG6M+QoMfM06TuBiJyadeyvoMoDEh5dsyOusl2NLIu
8o66PDYzZvRq6fLYg4mJ7Sq6pcmBVO/qeAph1e9aO1SS+6Q4TWc+0MR9L+oJ
7VQWUYVD+7dUkGZ+svmOMj+/M5DPb4LntCiDH0au0mbdfRlLhhLl6NlbItT7
kK16OsSdUZ1BPw+vHiuuMnMk4yHiPwKwJiSOlVpDioDnlkZlPV/Wp5Oo3mJG
m26NVDnXec/ff3u4XYgWebXX3KYo9fUA8DIvLYA2CJISdCrH379j95b6jTAK
+1bEuimXAagsOzR95NsuCa6aGhR50bYw6mMZGBHnD5f4LcCwp773sw2vjtVZ
0ZIcXXuRaaYGttflnsHOqTs8GpxIV2MxZBc5K2CqWjN6xkEI0HwrZEfvbJ8Y
p701akbtRzn11l30O9CufKy5GxO3Pi1/3AyBixN0/cq/HUqmfUd9YBFKv2R3
sNQAOOSnmblx7ell9GJWI+FmiEAcoiQM4kOIvL9htDJca+iZKcOVjoAbphQx
5hxpIWWLhP1EPS6cSD3PwUA6yHL0dBYNZsZB1m2ok6jB6A4vwJQqPV9ncAA8
PacVaG6VnBMOSI+bCCWI5WAd4AsVxHjkh48EDMRPu+cDYka0UTyEhsS5kLG2
LafGS0w19d3hFnKadvXoTMYfenLPiPRoOxamLW2/grEAIO0HJbikxzKBtcA9
DT+7NSZtKLxAz6FVhFtG2xjLZ8Hy5esYU+H+ohoZsT7UTdZSiDvAlTlYkzxP
4tKRtgE+CtSs4xp3zzidgCUSTV5XuKCoJp7PYSkwDwo+NQ38pM/en6sdgwEJ
Qgy0hCJlTN+9PUOTqA7MSs9Km84AMZ65yvCxDzij501p5yqvNAan4DBVHZPZ
kVXqSvjjBCb1hPCTdlni8m84tW2rTmGBqZnEtkoqJ2WBtUgA93uaiSnhEJLr
hqdDmzuRJRAoGQwU3Q4dLwF4A3NW+ALQ8OE5gh5QLRXPI0ylFT7OZYzvQwb4
7zRSaik2bkmp+Z5JXRZywDDgSu6t3UI9rnOK0JlB/QOnWs29Yw6p1puHdWXY
tbySUrJvNyhPO/DZpgGN56228eg8U13i9FhbObmx2VFxr6XwQP0ZHhzLCQFq
GtGj9uGwXQkkepj1p1PcMN44Kx/yzy/IMl5e4wyPsmdNYygOxLYzUdZWAiah
SGf7cpgPc7kvG+HAoxjihrin934mlkOYIWPmvEKmhoYt6G7tAaNdi14M6Kkt
s8ndTaDroMf1PvLsYcQ9xpjOuPY0R0B00h+qNBMkTVQYD60rMayjRjoLF2O0
IIEiuLniDenC7YMDxoFbeb2IN2Uq/YR4L5dz1JR/9284mzPZAY96BOk1t7Th
LE0aYTMMzbfexeOgf32Gd4q9yWXQSmz4/tzcAKZDd3JZpO7iNHiKlL5kr6fR
szW5Oh8wPg57X65FvheUL5ogP/nXd10y1QNApI4TU+1jTI7RCNcN9ngj0N+b
tT6livWWBBalAuTGDznLEyhYwna7244OJAYA5/QKJ42eND3re5UVinoq5Ity
f/aPlyw1zeeYGuChgK2/yfG3e3qq0Mc9MInV9Rwap8Ejahf3Ng9gUDvxTxkA
QdmaRa0OFuR9N8TB8IZDjcMULjrEkW+rFKb/ru1U50veyWLXz6qHa2aDFLZt
oNmUtOROdOSTbyMlzYOLo7Aqu5h7+YWZstGZ8YFnsZuxVnal8XQlhIx9rc3W
rZOBFwRviyUfVSh8SrvVsQt3uZ8Yu/y0RS2C7+P+bcfzZbovwpewEzRw2Yb7
a7KC8KoeHJB9qUyzNTNnYOxGruiYmBrt1F41YOfsanf39O1cqcINBdEJ4D5X
at/3ktn3tR5+uMwne1ZQZ9VzzThDniiLoA86oglKjYAfhSVtGsGa7wuDayLN
tLnWo6BS/E0znjCku5232bsQQPlTd3iqeF3L9yLTTlLvwqlplqEN1DeNe3KH
raqY5oKvySHh4mNSdg5ursC0kEDbmdkR9165Ij3lqfux7hp/uzgSO49ODrep
nuXW1wCYrAqxDwYiKlBzHpn2zaT8rocllrND6+A5NrN50hW97qpvPcWwx3v7
O7cRBswPlBOSgYtR9EpJVxrzg3aIwdl+5yywSZtiSLo2lyqCLMtSkladLG5J
GooJ9CKtJMu09F5MgeBfJBnM3cAhsofqz1YWjJxMVJmGqNJcPyVjou6mOTTW
fN4c+eV38LFuSs4hB0YJvuaLT/lh41IXEupVThghNUoBMaOHC+0wGacHJGzi
h4lt90/ONGANgoFrY8XlFSK3aMQKGtFQXehonhhu2CE2ohZD5fKVMKPd+gh/
3T/POYV9DpHta4OtyRng4f893VwGC854YVDyB14zILeyejUorDSFc+m73DIS
zNd/1/WgJMmFljNLvIgXTlpH0RWrQ9/8i6UgP7sAJbrUlYU3SGzkyyvWWwL9
WTrWddIfaPTWOckpqKxZSoTgvQgt77fe62DS6eAT2unYM5JYP5kOtCnAmDOk
NbHOPecljtFGUcAY7u3lzIJjo1FCvPQnUuX8Mj4G+3EmG+i2yEztyTQVwzwj
fj3/Lc3CEaJKMqTB3YQbqY9kWlLHmJcTc8LXnbcMEHbOYMy1WuH/nf/soLt5
kmGsygg9QghlhDrTBZV8Mo6ZChbEZ0dEGzH3bbTSnmC0AblaLkg5SZnI0rSs
/NNmOjyFiYOvyIob64CtN07VB+58XQTKZpPOiUb27zpalpAQKUkJCQHC1Vm8
SSyV6NITw5pky+MEXv8sH8BSqjNB3V/MoEUubP0moF6xjWsQnQSJZ28QcAOj
vvcLttUrvGZapC61aZ33MfzTOWvOQGHyNq6HC58gEmH2xDP9Dx5S51HD8hRi
mQc/4yb+4z7soszy5NucvBn+/Fe6pRO64WXH32lyFpJd2g10hRDgJQOvEhgL
QwU11FPaaYmZkzk+uiH56kFhgA1//buoLAwU94VQyEDebuD21y9xuIlc4HnX
0QiaGgjM3+HMgx8n1TAq2nOsDlhgUXrgiOh09VqEq0y6UhgjF5w1OsODDLEd
0mj3bbEIr1HSRLHnLU2XAJ0sM72FIAC2SFPHz2qtiojg+bg0GZQiH4Lwqu9U
QhIpgWxyQaNUCgGQ8cxvvJJOiaqYQ5FBNwDENL1lFkPhWedtRljboN6nBLH9
t25GwDV0X7yjr8YmwgyGzRVNh6ou5ZyEkEfLXBRpswVm5h9Dq+pT1sc1YS/b
xjLP6uj5MXYGOMDY28UJpKhURdWf4fh5uLIdAjmaM8jEMyR7KnkeNjmYX/Mn
NERxBAKipguXgAQqfxosMl5a2cbOYysxqSZSGKjryQtGiIlLEqYvDsZuGf+S
Xx5+woDL4Ta+k6XBmbFMj+k6Co5sQBFAHEbNdv/Wyg+y2gNbXKyge0B5KG93
jLtIqpIV79Huut5hT7GV9yzMRPM70TFNqwCPUFAVT1WpGN2Gsgrenap7UIZV
3Y3U8iriWzLnTgCVIjoyRUJ7yH5eD6le/3iV+SnqPV/sHORIp8ZETMivPITm
pVtkagonb64TmFWMH5D+LXN/20V7vx1/T0EBJR3Dmmk1GQmXhpyyridIDgkn
Y1npQIyBfhDlPGd+2U9Fglux5b8aTGNe3pmOYBUVyoCEHyOJ1zwBZxM1miB4
pQSZwsx/WBKHduG4yKIiToPGPNcm/51NN6L5A2EBHujStU0aQ9n+OTAXaMCH
M4tJYaLvuNtAOX120ICEXYdfpo5Nu8sLjBIWEH1Q74nooUCAssa2mCURZUBR
uXdU+8QO58kIyMjjIbJNB8yvjOKGf+Duk9XoErJQShTcD2m7kSV12N4EpS1K
StlNNgGy3Zj3SAL0/Mg0rgSJLNt5OFe39YygpjM5FvVrcex4zwxWzQEg3rAp
xUNqQ4NHofDYn3cYd64RszFbnS6GCEhKtErAZAwk/VXc87Hp1Y5o1SKRNl/N
NHnd25SyJBcJr1DUvL+xOi/2VvFlvDbfa8t2LYZvtbLx6ULugFUoTnbGV9/p
UjzQ/t9kS/ZiqMBRf0sQLxCB+b4orn3r8FY9P/jaSnM/V8/LmbGMAXVD7ah9
ev0qa8yJd2V1oJY5p34oqbeztSYZfvgimGgNDmPyJTCVPrryhiqRWj/smyKf
oO1qavUQtp89kcuVPwRDUZEibiv+6+2S7xf1g3JgY54CFRx57+JsFsvRzLbS
f9HEPyDjUg48ovN+lSgEYin1gMmY6JoBInY9sq4SKXwTzhwnfvnEzIJs2Xtm
UpZoa5PbkM2sTkUsTPzNXkyboAj98hgC20Wc36qc/G22Mh/Y8WDoKos4PdKa
iH00H4omxRWw5DmL5hUT7tDdk1wfzVmigTjp89H4FXqLREFnr7R5Yihlby0R
izoyy9cKbLl/uNp2ssYZYM5UvlEtgRjYd774BxkfJdHt9Abye1V/TVw3jLrV
kasv4BVRs9OGLs7VizmIFgxxePIAe2PSXJJAh4s1DmkDlPmKZht/vWksa18U
n9GHY9zYVynixq5lk1JB/GuqNc6+8pYoo7lPo2fU/6Jm30l0GN3K+CCGZNPG
WgywaeAq3AQJda73HixdlemtTt1AR05eMAsDNnYtzp5o4V98d45Nm9bi6KJA
p3OlDwD/hndabDFZ8+D5jCW44gwPho8JH7LqrVS2gwe81BhzjD1ZL2n6gHf3
pxr7j7TGc/SrpGZGEU7fA7RJhSqz1ILXBdRpL4Y+yEu+6ixxOInTrj4CBpCs
RICrif3/CO1sUaTk012WpL9AB7TusFWG5Z1jR4Lq+FG7JXemom8DITbDSGn3
FMIkD30wDIEvVSn+Y/0nHHFa68VGD3LHvf6wmlqmiK4JLBQe11uRfdfcGPMJ
NI7GriJdFliPs0D/ZLGU3lBvSVsPrFhFtfLqX73V6V8hUiCvmWa2Bl7aHq+A
5YYBFyW5qgwGpdUQHvFCSTmmEuLbitJbpZ3fo1E/7xZgP+FL7exSobVSEE8g
WDEsKi9e8N9vH73bwOkVa4vxy+BEDSjuMrNpdUHLmpVA2P7I0ocVUcdh3d9g
zZlBGnQR+M5jsLMebQjtPANUxp1LsD4d9txj5uscWoQHjMqy9EhkdF5iymWw
yxlxlFIqmMfrvd7qMWwZK9J4M9lclpEWyKTtwEKBlxKTvwYcvXIm9UO1kFWs
bgbeObVSu0naJKkPoIrWZ9ERkXezBdEX+YoMMtdGypyv+N9ywDbIMKkG37/n
w5jMw02Dd/lMlN9hT/Wcs5Qb7zW+opbIgG6g/lqQaVosncznVcwEli4WM0TQ
vHh8f16ErhaFiFYHrOD/0Ax+QdUx33LkWvK0lZBUT8IPIL3E+oSfarhAHuBy
KY4Qjrmlcmh7jjUQzCE4TXA2r7QxL5EvDXU7Go4YWYvrFsrNNhCQFVowuxpV
w1JeHLyUAcuC5z3Gvkytdb74Pp9GNjstvhRTf4yADGGAyGqfMjYpnvSjcMIC
fVMNCnaFgzXzgUxiBCHBFi3eZQK37I7cJKwjL5fcXjaziW8mbLDGIYeidL9f
41MNxuoSw7EWGYxW+/I9XJy0XkFeq59eIoVxWr9rxLq6Btfd7+/9IjqpkDPf
vLoGSCpCVt32CSB3fC1/chAcPVm7TeWFw4UKJ/SRYQ9nwHdf8MuYn7xvl1EG
ILIco4HCOB9vC1ehqrRC4U88zusdG9nQu+c76zzWwV5gk2Rx0TwqU5Sz35dW
T50B/8RQFaABguoUMpC00rZkVZnFwSznx8xIfmOn0U42ktHEP/1yE1JuH8aD
sw6lRSF+iRa+X33fbecMxHAlWoXfm1LqPU2wSD8MtMsKCTWyUYBcZgt0aFU6
4nZ8kvNl3fTjE/LC8Q2wQKm4TDh1VwT2sxt9eaxqy+hyWjRrNtprNn1i7Z17
BcIvpDqE/+Jc6zIWRLmsiQPzbatRU1ZCy5IERzmAjntcWFYAgL2z0j/WCT2I
QAkI3NhW/yUEVG/7Ia7MTm5PdN1xR4n5C/U7D/IeFBgTmZZhsQw8Q+cMWB6L
naORYUk35EOWf2Jwamn65i/CH8ugbmQ5cBsyySPh0jcJ0e4Tx2c3abLG/GjB
xmrfovE1291bMwoVxoQmRrubnin/aSL7VbjifAlFqQ5knov7uSjM/oSJ3ddZ
lM787IRbYH+5lr5TSaSOZq8JVmtC3+Pbt2jwrRfjxAIXUerK7RCd+fQ6TuGB
FqdGlcrwq9Xo7X7SI+DDEQT/IuU+gIueOsUyg1r7j9EAAbCKo0h5PL2AJBgI
B+GUsLst2RgFxHInda4+Kztkpqnd+KZpIArLX/Wt0+tZ/Q+ryKFalBjh0YkA
uqekuy26s5S4INv/sgBtH8ShflH5sKNMd52R4kTg8Q/IUjccGwe+6di5LaaI
e5fKSx8kTC+fDGS9XscPBG1HOyommwoiD27lj/4m6P9KfxDBSV6yVgO+sC+U
FaMyTafibgXXShbA8qT2gNNQ6GEeR5pFpliFYRkqmpEE26ZNwYtAaBnhZIK4
zBQKXxWAYZ1JZZkzg4IOoBfStgnxg2y66fF89BYunnXNzC1zTNNH1Ua453bK
xPYsblQOU8vGs31irr67OH78deac4VGSR6IYkUtDEsiMZ+kCxDwHfefZp1Ml
POXn1QTxugu1941GtpXbGpOqBWInNZMnfTkrna8EF0Dxr3x32qunWzHxImr2
ZJyO2xWiCOOXyp5TYSzoSl5XXc6PJoWeJ838YNDO7VQwMg5ETNWqTz7GoUpy
DtTB516sVO1zn6+oojn5HhIUInEAu/8S/yK6cXrGSHd1DRiobzshz0LbS88x
Rz0hFyaFYw5738ddIkFK+S7AfbgqAXLveTgdbqIbUZpRk5AxPaeFHOVFIgAs
3AZtX/5U8+0HGs5sYFF+P7Ddl1bFSHj4DH0kO3H2NRVo3RHX+5JVwsVouMFp
34t8+rhyx1LBGMW+ux3sOfwH/b4rT/erCpbPJGdlZCSTuYo3MYothVAxw/PC
q5vxP0Luq8hLTnxzJydKOfOvtOfwbEfkxiIY2o+CyZ9kyCecgtdnFEzMxqNV
bAvsye/dyRnY7OGQBQQEzVOLQAPxJWQ/Gofmug2OAh9YCx5eyFlZtyIXI/2x
4TDgKmxDCILnfAdBHrJuxOGwCo+XMayOm+aTb44vRQVYDJyYaZofA2r59xAF
irDo7Bn4frH4FzypW4slrktgvZnolfdLmXFwNUnhO7YnrJA1LKhDE7D1Enul
AjWyB9r4yNE5JPEJAq8AReXSwHJljc+Smhik/yRcpxm55Kut2iO33ND+Ir4K
VceHkKOhrVl2uXfTbRWPnq9Ni1M29XIBRXCpRfaON6GdwbET6OQ4gnsAdtxE
QLlX4fxpGTgvT8cWdRVImxHZ4pfoRk2uCgdpMdOqHvYmRLFYLtfljAKUFemL
iOhJqB7uqsO8iCHr0izonYxYKwLNVwkOYrvA4n+E0olWY0iehMOgiwmsUYKu
sqclf9HkLcRS504FLF5510A1tZrLqHSAdbNoszUGCr6/sxG85Jg1euqHFKZZ
cdZ2o6xpCGEeFrZapBNcVQDQrRdxu4SJNCslIDtlj3u8mwGNY0cqoN8sZUsY
4N1wFaFnYsn+PPHACV/rKv1O5meXiuFpp7el2OFmb9dB9s2urDbYLLtfaI4W
zRw6x95HpDPDItPhzQevpqNpou1Kf4zoFm7DShcV1kj82e9xkHJhPJu4neCD
Ui4Nr3T6f7sPbQv8zTKnhlWV224/+QrWTjUY0E+pJxrHx2QBC+MAtcFkp152
XTsOlPIE1o8uEpecFY6qZRWZ1CmG3YqaOgVHSbgQ36S0zV11AhLctWRp0UYP
/8KLQLvIzD0SIwO9L8PRWKAxw5ihaoeg9kQYiwn4yku7I75zQy4Wqn8SiAkY
qyCo3X2T6hNoxHn+S7l5Re6RZlsfkjgdaC6EwOXXxeT0jIG1jckQSBw3TxkI
M49FarvGgbWCt6/udXUJPpAmDJtq9pxXy64T5QutVnS2/peDlDgyXNZN0naI
2CngJBT2Hja1ovziBT9r2XUo2ofWL+Usc8fioZnqBDZkLsWTLZ8YN0oldVvB
UmeakE4/r5vWWAUFIidzaGAuPECVUn8POjM+2e/yVJRHXHL5DgsGeDndg2VQ
8+boorcH4VF8u7Z5ZsLYwM30geeHhSwzfe4BB7s1bWp9JYZc4q0ulUNg751X
oxYYlg0ZviaFJvkZ4vmfldiri5wUBjw2+Jr9aE4sCmIkR2rImeLlv8O5hMkR
7ON6ccrM4gtfxjgnGWq8BLzFvK0peS9hW4sC0tIWYd+j11a/M0whin8r6XIz
uaSOIGip3Y/YHtojK6EJ1ewsX8e0LPafgVj/v5D50OSIW/v+AVpMFFmr/3i4
AQURHbCCzJ9l62U47+YtzNT9I6X2s5OJK86DenB9QUSpqL7EoUUGYTv6kRsF
x0JxysD8VDdOtGAQ/4XaVSKreXDz/RS2SWKntin02mR1TqSpMAddrTQvgCHJ
bgo5lOaXDA4MNggEYbS5OWNjM5uyYZmoHPe4UjfBM4D1VM7FPqAWl/L/xH+b
fg0xHM6wTf782Z9ELgABPwy0eTPSEMGc+K9ugEpuE6X79IntCAGlUe+tk6bw
2PDqcHII+KF6u8JiXu1VRdxeIkffH0ijp8hiZGCFKs+6YUe0b2xrKmTh68Tq
qePWCLFNKIK8zSMUFOWUKMKYbZpqKBECAYQ5hyDCkWZw4GSdJ38ljouoRC8T
fdZev9rNxAL1YsnxnD9ylK12uWmekdVKNovv0ALmDzMMHCflitkyBiAYzfIP
J9GlF26HcAsEGIsmWLy3PGHRllpTh4MRMld5NAPVl8HkZDnljeHdHoWeNg4k
14lxD/5IYLU0YmpDdm1lAS3lhKkXWyPXB8dw/IaLr8DEMZIRIfcCp+N4BCVk
KswDMut97jlDJNcIQEHWmaom4xBnKjvTkhtkk8unjnmmvBr44MNtibSPTJo1
QBbfyNc3y9uUxANaEUTjCvNV+K8GlRkPD9NRjCQ1ujDk26Cgk1bH5Gyhk79P
vC8hA53Wxo3K++uqle8LowvkKmUno3+WBy1KTtRpWbs8F3VaXyTCkG1gphv6
0JIHgb0r0KAxL2EbFjPGa1fhu0EhVZ/vPURDNAmcTJl1MlyBzynkFwEbgdl4
UqWjgQEFgEyo0PRmgdG3mtCzF2Mm95TU6XcIFV9dOBaB33gnmDMshfAKmIvG
WAXWRy8TB6U7qpCZYGxUEJE3n5HqArNOqnYrUh3w3EvXCbav8XSKdbic6Vl0
l1QiFvgdh8KFjNgameesTxgg4AaGbuD67qBlvmRa3AhSBf5Buu0VHFE8JkgT
hzOl8+RqzXHWFoUYfdb7Zr+YfS7o5lBi5GULL3S1NrFjgPsfxqFHq9r1D0mY
7/TKf1b3Wb/wpVXDUMREvdkjM1JBnS4DWETdtrBqQVmA9QmZ0YoM99vlFfbC
4xuf8KBE+uq7O+VPuvzKfQyPOcbzoQFT+IfWBrbzmV7WNDv6VdiePc8SUV0g
zV6QHordUmQtE9z8hY1IplY3y5F0C7sn4V/xUT5hU04G8ACym0EV58kB6lAq
dUdEsOuqMIKNcFb9wRWDvTaTqDetoU6Rg2KXdTKpgybhUsHf5gfxO3Q77NhR
tkuugh7xGlQaCO/x85jzIeuOs7jsiThZr4Ra/Qyw252OIfBvMWG4cCPNCx7u
iazR7PZIH4gwv8bUGyPIX7pCclOmxqIv5W+VAuHLmVTyp1h8Sjksp/ZeWHrg
X1hud0a5yFQenc/mzTQEi45q2FHKCM0y7GWif83HIq9rUUq9vwP3RIP2nrfU
/2eaXr1sdrhRZMw9fRXuKVT87OtEuSa7KpQB/+LzEXQdo8PDbFjK0TGfPqWm
BJVP/51HswakzgfUGcrBunC9vq4ZkZw/BTZPO0PVG+Agts3PDqqMufjbmiI4
/IOfj1r9DqQe9tXO5yMpyULvs50IomUCWkgHaxsTvGBzJFB6B6iE8RSya0YB
ax7Mi1kylxAJ0Cww5VLA5Z799Upjtfu0VlWSvZDGB28alOjK/iU2g3vpEgRk
h9rNjb25xnX2J44JT5d5REPBLfNNHkc5yErbOak81BMtCk1QUeDxqXoXCzEw
8emne75yatFSorLFkuak871rsjny4WRlv3BiZmxtdAy6b5tXuLbaCX+Xli5s
goKXylBauQP30swz2AnMDyvvoFppfX+lGyAaMTzWQ4t0mkJyLHH+VlIlC14L
ZcLBUV8n7cDkTilEylT+8RLFXgBEdKb4tCFxLyk9hnATa1LybXmo6H8PfmAK
QWjiw128Gkjay9ibylGo7HJVoQY1wHSzg7OedOTdP8TsH6MWytHca8o9boPJ
wIas0VCf0bmfzoaVkBP7JH9PWEZ3Cla4QAgSOF3b9bQ1klM5WEsHboNYHwys
ZJERJa024U2T1kZQ0onm/IgfhcetOWhgBgTmvQxjAVqFcsJ5k1iy+Ld3eR4c
wFl8HfL4rZ6Xs9I07tlKoguTwu9ciAXbMy/xSHqz+dsxIGKRKtMkH2A6oygd
yaskyZ3/WP6ab0V/robrIRKfGFxVjD4hQfhEw9VwZyeh90qPykQ8V/W7wqVq
XU+l5oNTqedgoJmWeAF+Z0aLS/Xwq47aZrwjS++eCBCIMcqMISIMFzOX960m
rq8nnhq+s9RXT6W67QkwWZltR9vYgkEDzzOriOMKJByRPnS/uMTb25Q36wig
g32h47YehBuc0wplRvoXrjw7WYOgMN4IZF6dwx1gV7fhdfMZKyl2bHeANK3X
5S+1pMWw+A743waNq41XhZ9bl8uO76Ml2KL3Xu+qQ8xbkvDfI/33LLZU5ttx
7UASWUZL9uKhAfMJOW3bA3ZPfm37vWb2cpBN/JnhY8b0DT6EmSMzLPSReBrK
HXYueWVEXbxagu0yAxsbEpFiZfjeBYm3sL0f0Sc6H/vBIOse3vzoC8mH8Aon
5xhEFLqWrTOJrc0oqsJPPR/xw8awUPClFJUCYq6jEIdTpaTCuhLTaowdYtc6
ZRGH7EW+u/1dpn4S5Qbfy6lRRlJIXtdBfeNzUAZaAUxqMz4twvvoylk6Hr6l
WVgmyN5U9N9VYtzzJgpO7HVQjjWXk3Iy4sde1mjiQjiEpqdqkC95HtiaJdtv
QZUd5V6j8Ry7bTnVS/jlM1BrhMt63q10t/Gj9+7H/HXRwLc2v/WSvJnIBYIB
FBsFqtVDEDprIN9Gw4gFidt86ICezq2XoPLtVYA0H7qQx8BnOjQYrofe8h6j
BvnhcrZwEW0wIFijQiAL4wz6vs+fZsWGLr8XCOwyEoqAflVL6XTsm5X3Kvvo
TazIUMslh8i+bEA2kNQtKtHSpDnI/YrttS0a+aY9BUPz34+ARer6vDhAprpr
Tx08lu7jUwqnUV0vMzWC3F0iDNkT9wYa4eScMJtHCN2p+gkXXEVf+USeyzrP
xy7MbX8EyL9PsAImcV1uSRbDDhJEJC1OF02/JfBA3mm/NlbQXW6JssDVcXSo
6sKPdAKdKQextK7nIUJFrNw+hoYx2DrIIFcfz6L/UsPrAKiOTsWOu3jWHVo9
gDOL8P8piwkagtGyly19yI3yLtuRgwM3XTdE6SGN+U33GEmYZ/+RYGhHK/7s
w9hs1AiHEL9BJ8fgBCXas0usIs5izCYMCiWl+MM0G8xsi4AsBF+7jGViHeNd
0Db4P3WnKBJCgeUCCytR2eTn+GHxqR8aMoCPorLvQVEdmhen0xydYT2/t52h
9LGCbICrmxwmDTbSGqWN/lt0rIH2slSM49+qFzrzhs28mJ7PgmZky2Dqffi4
qzN7j0PlGV4FnSdySOtEzwJ2jzEB0q59m1xBAXmPRF8wrIpSwD0vBnNP4rIe
KaK40ntbLfPXCwrgNrY9CUURDbsg9ppDPSZ0eKVE7dUuQ03n6XEo7yvF5Alp
6j0lrqZ7x/9fK9LZqwLTu4SB4UN6+pzDEIF782PtLSjtmv0uBIB6OQlK3+5z
CKRJ3RR+Ew99+VH3TQ4lKyV+uH93fuOPObwlWg2vPocr3v++F8H4+/naLexw
WKt+UaGZ/VLt7u64PfQj4XoM0EzoozpBh3LCMtBdebq7Rzt/P0tMOLhZumpn
BbI2RAWRyYZFkAlElIw44seiF1YABrR39AfCdai/tpw1AZEM/CC6r093QkVI
Us2z7RfmuPbmZjRXAngM5K98xz/SSKQ7GleJ4CzdRkxfc6i2aBUJdq5cj7Ff
8CHgp5XOZnEX5gowk5sqeDSEhaMPM/NMO3nY2PEcVrjR6sTKTMine8gz0QPm
uKobZqb129MgPGSONl7tN2m4QuLudmnYVPtRi84vPTmUtyxJ+Uu48+URZGJK
95S5xH4o5cMFwa6bFCUPswD5V/0EpMBnRwRqPUlY2DlgEze9JuhZOIn6zX5J
IvBw6bjop2fK/LmmUtTi0Vcht8r+WmpHEyLwcqVBketwuIDCcRb8DFLldGdR
5CIYbh2pUSMW8wkmr//SOE7xkcwqnhr6jq+Pu02j050izmHSHVRmoW/Qu8t3
j1Nems9Odx7IO9tq6/0OVcLJmLzqLDtKVI0fY+CxSYyaKXopA2JRND/tAyS9
db9DiRQuFbQjymiqxqEeslfEDnRArF5LAPlVYBkaOdoEbnQmUXcB9OBfNfu2
WhjAKnetF+yT/29L0M5Ar+JIHCTXKQNQOlbOfMLgoBGopuaMY9WPun2a5hAy
M6v3KZKg1TkKZYh09HxRDwnBdU7REOm+fa5qP4YsIrllVuBqDLrni3QAJFBl
fmIRGeucOHMRny6T6rGsz7noowL639ATsDGlq86bTm7QzjnZhEsLiVDqsMCI
vxewTzDy6JAxiOQ7CaPtWIy8MzH0lLY8fiP7CMqJ1lU3cb28vNB3DssK3lOP
PwCnmgghB8RbbA/H1hwDr+hjHmUd3qXl5Zcz95jiODaTzHfaarLa8Bdci1HU
9MAiwFXOI84fmPdbn5pWb5FE7IiMm/LTO8VHQA1oG2eRl7vxEiaPPtj1Jb6E
WkO5jVP9fJ3hqnBEoJTkQkofnGW2PD3Ymgam4KusUo9rw8+y+7cts0TCef7n
sFNgZIOUV4G74dffUtz9TzDg3Jc2AENz0sW3E8cjGcZzVJ7IPFiynLgF/bNm
gjZS/AW0epzG5ytA3+7Jcpz7pre/v2ih+xvpD9oNTffiHVlIIs+CSJbQrygU
EIKTm6LxSmQ5gEMx52E1PfwfPPjjqTn30MgIudQH0Ie4OFyaW3tfIEN0lZfI
jAr9oza8li3fjMRIASFP7kd0ceMGKa6738JbPvVaByJ7V3bYx0/VkxDYOvMW
AKUb05BLeSpG+9Hn/J79Ty4J+ztH7tXiKG/cyPNnUgzVphfM92o+m2F55CFm
+BokXwOC5ImWhV73+Q+JVT9nSqCIDz7f+i6m+0Sy4Uhplg1dPyh/dZcI5Kt/
jPKrevY1+2Wc6ixS9MKPJmjpesq9dxV3zEiDUMr5f4c/CdAeXLo41tV2stbV
pBGF7j0lYb/KWsRvnT+BWsi+eL9mrbwanfz++1zj/uylGhEks8MmGxgQFv+Q
l4JxEHwzuyLQCsPabCfB2DJ2/YmrZNxTmu9/DFODCBEd3WyAEc174gV5Vl76
LrwpbTHeKDOomz+I/inUd7AhbFnxhV2BnbV2/QoIU39tnhHJ/VEfkzdYD/l4
3qnrsj2gZFXE0m06PpTChGL8/glZf4LSaB8GzOPuuwpLnzHurjiifcymLhGw
06uYW7kAX7cn7osFG3l9IWZiz2hZKwIY2sc7qwrd+fQadC6H6W4P286wh6+l
QqS3T6s7Df7D1UbnTF+9rky3AeqjTLXGUIXicew75AdKadltMV9sjSHEoqoR
KvZ/shVOifCbbBC1ypLsVH8FrQ0lMR2ksPu2VWtjqUQcBUrtZuS+0sJZmMKX
geN8c1db+GrbtMJT6097GSK13nQDixCL89kUrGjSkACGv328BWaEkLqa7KKp
0aY9hjDSSV2cGCeM7LBVCnejN/eioMDdBT3HUVPytT39pb2fBdsbMX9wvOiE
mS7lBZQeHob648fbQBNTUNemMi4+Pn0nV3jwWuw6DmfFnfgACpGYm2kNJZO0
8795Gzq0T0Kpd6BlILZa3xxJQZBEa6n9LDfYIQOKbLLU3VhmiTja1Wp+j9Kx
PGAZIL/iJEWb8gty2xZh8arb17L1nEl6jue3nyLZYJleeOO3xYFUbDuXk+wE
9Tns3fj5lsep0nDoyS4ZMHpnxQmnTX752M1pkWq1t+Df+Xul0GTK5QnZ2Lvq
VpFHq3oXDbVhcdUXiemKdW7+nVIkE3nP6+A33aua9o3JmUPH0hf7IF8PlPlK
8DzDhP4sPt5KTzWs7RlvQH+Bz4PVBBIP9VyHll30T6JAfh4g3JQgS7Ub9fon
b+dBEH7pmT53vWodhyOACCby5fGKdPUjmUx2+3X0kzH9Y7+4DP7nyBq5o+8j
+lwPr9YnLDdlQRJzlmHo/KXmY0wCnXA4La5E3At3Sk6IYN4FLHuIuuSOiv7J
rVCfJOUDST+sDe/UM5vT9kbeREWPYnQ8sdPehpPDEDNeUTDRRaugSk0P7DVZ
pA67Eh6qK0ZYygkeBKAzqehADpQwqFnvFnwqmpv2O2A8zE1UZqqeaVreihk5
QMjmSbNt8HAsi3qgKDkdcrAgMeGT/LzAB/ySvuU9036M/lhspWIvc7/1X9OO
svnAd1TlBuwSgjWDliOR8F84z9KmBjZNORO/sZwalZKLz/dTd1pV4nFESz9k
LcxaunwGGAU9Z2r+yEcQsFlr6huDd0u+Lt0qGOk+zUmdXU92X8nl6YHEL/Vk
r0SspSYykKAaAhcDfvvTttuxyY4Or3IMZyBQ75dMBZEEWI8n6pM2u1spxD/9
WM78GJYxT3n0bFYH3fE+AFwGMouDiv1zz1f5k774aOgqfKJntlZLnk+P4OMh
gKwgcEF4JIC0I6yPyVBb59BYzeIQ+eNrAeCCFJAbox2PhlEsfLjs1+aq0Lf3
tg1kpB8YCWhXludoEdEdNoVnjolm9k6f5O502LOxVUER2cCDmHaMknxEJe3Q
ERXNXDIERNfRqFEkTfRV2KCyF7B0O8A4K+ZHeCDk+GTCYHjUOGW6n9Ywj/4Z
KCCApVoPp/nhT8M77x1hzCBcg9KHdTmS9gLBWBil5qfixWBuxblJwgnfcL9C
q5MhW8PVhKiPOrmSnL7lDg/fbutN+OeHZ2B5T7iEAkDSVxff6Zty+JMnw6PT
w2tHfQEEWD0h8x9Ca2gWwZiTKDJ7SB9dKI5CVaiy3fGnQ9mayUw9iQ0MLaxy
fiwOlqeNb6qUGz2PYzly4oBV/bwpQGA1ry1cvz2vthiRVc30zpBtqenvSH5B
J9NA0n10Y5HLTpStpuoPDgrXh8xz8ItJuXdGCrKB/kcpjn+aZuUcBBdVV8cI
1fArgm97FRoLIWrG5hTgkE8Zmeyndlca3JSuZ8UF0GncprOSw2geDSAIZs0u
VZzERKlNFjXfLiz7IilAJwyTpfQni0xd9w6EMQqtlBV6tEtCVuPCur4MOx32
OYn0UgvpSpeYmYlksBJGeQbLeMpxTCMVyrqeHfwbOhZZtYO+mCtvRCDLZgNj
BLk+BkkHMOzUo1Oc+8A9uoGec8PDdF4utCz+Jrzvqa6Pngyap3NjECBEFJND
PqMDUFC9nqOb3G6Alk1LXoh/3tcg+pl0ZTWd4VbBus4U1ZK+dZXgXPiAowpn
EJ/YM3lMFrFAmwp1hUWX0B7cS6V6qc4tDGmfc4jfB+rs7MrecUmdOsDEoOg+
XwxKou4jDRrGDHrzMgLlMOoo5/oOtqZPjNeRT8T7rnnJeflnVP+6YAZxkaiX
WIGv0j7kLuK1jtqhzurVoKo9q/3YdGocL3kLuL4LjGyupUN159TjsgVOhiPL
9Lx1xtVtLd9XR00iOApCl3PA8b2PpGp2n4WsrS+QOsmQXGUgsfyzgCEq22fk
F0LK9Ry+Vaef6s/2Qt6nc7tsv8cQf2XWlayRhmDht7ZxiEca8FIl5Tyu2E/U
bCvwNNmJmGLgU/3g2LlRKUobOUyZO/GS+t7PYu9Ulp2hCqvIoKdUAYbLT57u
TCEvZ6CFKQLH8bpw42b0vXzS7TAHoNHgrek00hpnPN7rt2RjGEuoeimYdBgf
NSMyKYeL7JOnDduytgnw99S9RecpyK6mm8Wb3mlcWuz/nVLOvHr4udbcao2v
KUn+y/uJAOM+8o2KND5KLoyxQP8g6PmQq1DdwxqXD/k2pmUnbuhyca3Nvvh9
Ra9JjYT2J6ocp0BJR4eA7YP74BbUrGXwLtP89xx5MOhfEHgW3DjJ4PlkURH1
mYGd/3h0StK3HbR0l45SzAJMUPwN9dpvCkB5Nk1X1A8at3GD/aKToOLyAWsR
jspGI64zNBBmvF15yFMEZ0tnGkvX0iOt7Zv4FSDuJn+EPpyOUFdLSWzVP+wx
dfpbPYYqI0SV0vTgWL+vYjQlXqADjYubsA3ko8y+kXAEd2kc+MG80FKrDz05
DMGlJB9n1WQqyLsyqBDoUUetEflmv+yr0O1J+P05UKmmg+bBa6TqvxsEL48Y
fJoP/KOyi6l4/2t6VFg5kGtFAd/fjEo05aKji7HjA1WgTbZNA/YJ7tJIl0oB
LyRvwceamTgu+iefxNcu4Tz9Hq2CFL+5UtcfAhEGSj5ZKo9CXrC9Ab7tf7MC
IepDsWc2Oy1mpPhS9fFs5/r3KrwoXgmf20QeeXf0yLkWyzyydPn4zR01Std+
IFI5T0LvZ5sq1Q/eAXIsFXpGd87oioq6wAMNlTqohYcjI7d4it/1LTLmr4fs
91jtj52qJvh2jshzy23az0qy5G83oKXuTP6YjeS1NJYt47u1qM1Qme7LmpHJ
g5YiIPmFtzNfqeH5/O1iozc248DX5IGCJCIHnAOli0Dkami7/mnkDJM/gusB
Jt0u2QRKPu5f+gAgzLlhVPIJogZtSx/nVkSDR0lTPQftzBNwVVhx+uqfRIS1
FLuUn1ZFj7YRsPYGmZzBBuj4b7WjftEVRLRy8FJLUW0Z6prRWILSPPwcvoZu
GntxcePBBwdCqnDYOwBstpDJXGociQ1KHKSOCBIuJ/2KoIfJAXoZBVfOzupx
jXSoS13g72RTushQWyIPugxxLe9QF+jlOnQYzpCEvT5hVJ6NSHpi8gXPj7kU
SK/l3ndSEJtxWDpjOJDECttHoa1ORWdDhVJliSpvr5ptOqqxQvyTB3tlKho8
arQnc/HTH6Am4aaqLDrxfp9IlEfgrEjqbRrscgnEXNFmMrk3s9aO8Wj0toI6
OVbzCyotzum4rRDT3PCUs4SEmLYn9oxtbbZPJZ1FaGUefgXXBz9ifDkJWynk
uNXVCMm8AZIW7iEzQh4StUTwkgDm5io313VxO/ZOnxtF1BEe7YYztUJo1BM9
BRtxy/Wq4oNUZaY5jLcvPowfN9D5j4LZ7aF7Y79OvjJJwWcaSMR6jUA5Ma7n
01DPwmNvHDlFEPGFRDk/VkRZqMsZJnpJEFlBJadd20M8QGD9hPnvJoB/S8cc
qJFMC91qdLGIKwxpzA5pbmoZEIiyuxikBEJyQDEWfhzz6noR2Ca67izZXgND
J2yQPweSH8UCWmeZZqT9+OnmWIP4CyteFBStrLW7x76POZB3nlbnP60r659C
Fhbw6bmj8RCUz5LBnnL4UCtKsGMhgWgGaSqs4Xl/TaVZtvjeIlVGqpzTUQ1H
DIe7VcK+fMrYg5PTZMaZRKoAbnnczQteV/idW84krmtp020HXErV4WDhingV
tuTwmSjtPh6LyGMIC882tLupjqtqsDa1ZZv4/gIwmitLb6wDlFr0KLqMeuKR
3u57QsXz0hz88PgBAKhp7+WrdiF9UiL2+CPng05LUbjqKYy5w3Iyx25Gc2nz
dAGD47i3Y0lJVI4L6XqFikO6SZuPfTfVVBIOinTiXfr74HT9A195rXtsmdLw
/qOBoqGx+KyRoJSMkcbOCg6BLyQCDfh1Tlwxv+6J8h8M+afwmanaV1LO0jYB
vWOl/Gi4VovTTIEQzhh++FhRYwqMJlct03RTsR8hn6K5m6zsrgJ+txzxpuJP
cn8Z8g7SOLM25Gk4WcjY4XTg8Mcbix/TgT6UqTsCxUtfA/XkjW2puJzrsxwH
KbwMKcyCQc2lp0+/p4NKH5fQMCOYHPzJEcyqTTilC6jo9sTb44SKGIRYWSs+
p+lu3Zpn9aYEsYedCo4/2W0GFSS5xQGybJMW8LoUmgASHwCvFi8coVQYn/q9
yrEN2gmbYvu6WcfZUXQ0KYY7ix8uoXU7Ey/iH6Yw4csPc0RvgqlwY0My314Y
chfbOulgIC2zaoTBwhxG2qUUN+PAxncKt+JnKsHzs5nv3ugnkavsKOyARrAI
rrDSDfBYXLSMUHN7KFKZp/B378jILjsxKDSjwf57LtD89I73EuIuKjRwknzs
KBIY4d2t2ovzvFvJRq1ut/q7PAFV4bSF+kiHcvjUz6DtlBu0l7n07xylqVYY
SP/tF4SwDDHGlG0yi1ZF0ITZlMB6Eum+sajztPg6TX+kNh0Zu0ZXertplhkl
2QcGjleRvAgkJMCgSokQGT8qFCLLhK2WaD/pIh9t8dbsOm+1CEINPg7Hi+Uj
fnaqxRQzfc/2+z5wFvTkPqnFCY22J71gODVob63m7uUMlhoO9NPEe7FhVkAq
d/DVEJazg8F9A1CKspAWwpljgem95rPY68SNZ0DYx4WFC24CY6c0UHBFdAjU
yyBZx/zpN9eet065VLptXL94b71BoPwaQvkN3SSWGWQ2Xt44PDJtUiebaPG+
Dj54EOruIAaWwopr90B0oT3QpWrWMNPyYg/RkKYkQ00NaAn924sTZV0aJzD/
soyV0xetETFNr8Lkqy+XqBOZ0awoDq7HvTYOpwbdCoHzGD00Fr4LcF6bn98c
EepGO9rtaTsvSf7TCVTfQfRd+gyMHyC1kws451NAsNzTgPrv/NanAdQJeN56
2CRbznX3TfwGmcvROSryEMs0u98g8o525U+n3d79DHR1pJceQB8N7KfY8sy2
Sn4rKLXigZPskMl1IrKPSrcfvB4Ese0O7kmHCYsuni8xUtx/r5GQfo2Tz6Rr
s8D+nAvuFaJenkfMG0X8e5in/M7nVPhBLbyYNojA/YgKRO3EmTnyMBEudHof
Ruw5pUB7lLrol6yjDNGkW886gegKJ+pruLtRlqWC877AXLKo701i9bo4N1fm
cjE3iXq2Z0Gob7QLIaVRhj/fyBzQXOQfTkxPcb//+SSjiVV8JR8YtFhBK9xJ
4ZuoHX35SK2f1XuomzmUBAE2hfWrWl3jTPdIFe75xWtJvLAH8/ys+RQk1saw
7xVsVBsCCD53ovXGRGKyW2Q10Y5GqunOc9v8iDL5UwddxpzC6TjTisDjTLax
8mvsMpFoouM7ZzyhePR6/FjnHsalMNP7CrVrYMv94501x3vlgRqHISVMdVtd
+9p90JtdbZ6BuvpbFWl/m2kUoinACEYiT4Ne4TsueyJrmWNh3TIuqG6bZ2Dh
x5aktWmkM9YVT+S8KmfACq7BJ3S/jPJvQbwZx2lRwU9PjaraebyihUNpbsic
AX95MlgYh1Bloom3lcqU23EcrDxGQDSnZYl1usqrIGNCpmYT6ls8NOo4o6tA
P9lNLlHJboGacqBBljol6F9nFCImTzBoOSh/uC206EfpFrkL+q+pg8XOHRfu
FQmY0vqNs8Sk4UFTVSpF/l6wcbkS5uJLBt1TuzZT6/a46c200pp6x+hd8YX5
fkzH22qOEkemMC3pJrBK8rcm2a3+aWqnuxTlRf4kTTewJoakJI2h30BuAT0E
r1Q4sCpaE6Tzc5aL9uJ9SyJLP0UtAtlY6eDTazOuA9nyW340oaErt7GBNb4S
AAw1D1arZ6nRxSxmdf93QsYql/HkRgQGZdah2W2GgPExWsI2CAZKpaEuToXA
tfWHfD/PuNEuaPoNZhfjMcaoavZrvR78xjVDbteipSs8/mYMO2jNJt9rvNEb
nZZwCFydhVlVF9EY0N7NiVHAfyvfuJu55AmbBqPyp3XyKGkYP1pNBp+zp0Va
wQZx5WeLtCUKp1LjBL7ZDU31RJDVf7vaH6WCc+PSfaA41ayePC8bM2l+jVXe
H7w8+cymVAZ4T6OSDYEDPNwNe6A+QxRxOpNbyy5dXHPYZr7xPdW3yvlS2dr3
O6Gw5h/G3ATQPiOta2/fmd8y2H9WMH5ZymNfPS/bhkrst8ED3aIjlPH1Fkl5
lWDB1CsJ/c5tebruYBryzWJNgI8WNKqAJud5j8vGGZFJORt8LkXoLzOqXqXr
k2aEwCDyKd7aCKeqGSIFXQ6gB/aAhewKC0MI0RH+PWpynwVJcGaqOTW/SEV2
PzNBskuHd1PITZH0TIAcyhlFVgqsmpa+tafLbQCRzBnNSMUdRWB4z/0IRrc0
kJOru2vgGJ0tGMFtNXULOELsQOdhchbzIOK5ORZ8YBx80aVio7HfKrRUygED
o8OHAm/iTJrTxkem3u+rhiZlJniZXm3Ucy3Z6w9C0rC79ys9+R/kXT2+MfNO
XC5EchiA9j1fCVe65OBQGzmBm9I98nVPbstSXTQ4JPQkf30BW7k37XA0goc7
oZJceWEekPs0iFZ79UMICyIBBqEAHxrhPICSPg/MUDO0VnZ84LrlR5oHvh5f
xSX6OmzJRtllknTtaF6JIT816snD6q1UC7X3r/Rb8/4w5tp+tOx3qZepuGfv
CTy76yCMVisMptmT6LMTuM1NEMLxA2RzVRY7int1GLHCxQPswFSvlE+4dG7d
Yn5d6rnoqVxB60tBXMjJ2u/Bg3XNaVrsGn8p3JzFAv83SRinpyGoWpBkkkMO
eFIDytoEgJHJmrA4Tn8/NUt9x2kdzoF7dbdw/E/v6ZAWZ94oeASrwWvtJWz9
ZKVhVBnCbRvhtSl4g8BxD9z1toAO+H9S7yWC2Y8IvQtgytSMyyTEWVqf+30m
3eCSIEDOUlkMlkszhEdexjgNivpVy5hBAbMQEtMgvHPM9i/+KjgZJqpwb6Yi
cSb+QS9/xvc9n0180HB4tBfrZM4HWm3dMQzp/L8Xm7GQzTDh8n5swsfRu3Da
uRL1d7ylovuYQcoJgSWRtclJ/xiek9fDslugMp93vHO5mWznIgRrt0loC8T5
/o0duc+OOt6Xtw2K9Ow0QB+RygLjnnLJa1pP4WkZl/7IgERz+YRRHadSqcha
KERPOgbRCnq/xRiv8H9oEvY/ATy34p3+tufpLtWY9lXcxsGCBFyco+k/Bo9U
eUMnfcRF+aCPsLdeBZZZGv40X0Ff0ygZ0RAbl590QoHcwytgqBjsM61w5HmP
WWjwARlgiFbIvhMbz8BQ1AYKRL0CQHbt84rN4os3qnVD8C83kfTrKevS2owP
EwFEqcTHc/F4mKUaLbWizjBtAfOoDH6uYT3qwEmtjD9avundgm/GZTuC1qx+
vFXTaIL9wL+6O9oE2hmiri9vFJdtdy2bV0X6C4vYcRxNkxuYq7GUUq0Y9NHQ
E4pRB9Z1S6hCFGeMh775KQQIwtc/0NjdI6veqooNm1bAsY1hLGn2DXmDv7C6
j+FWpd4LQMn8MYkj8dgKlv46uCB8cXyaSptd4/r8fTFdywBbET2J1mI91fif
f37CzEvaW62FOxOAx6OFrqOrpvukLHYERiCZhP2FnsmIzos98B8R67p+yQnH
xUDJXhMWhSeE4kaVFfArr9ymu5B6a5e/TMdEAMp+slm9dh4dzz/FtOFxz3w/
HIVki+w9kvSe9i8zKtnJ1TuDP8+Xp7JNmo0UWYuZiTNFDINboUynQrJnGpqC
eF7gmLf4nZFUy/GwR4Ww4ITmWW6cX1UOcinyObO7VUYopNjdrtgsyolecWI4
xmlSiQT2leU7iamO+1sGWD5ncruVO9t8gdIke5zu5s2ZXQ4fN9FAOd+wyUnE
DvNfcUFdTdpISxRM+QmWs5p4U66e4m7KKFmvzB/7ZsWPwpLuEI3Vq0SgESGT
y+2QKcqbMRDxozFpJMZAfSUIqYPg8tlQ8/KoP8IzyxI3dY69gcLgShBQaP+m
5+zujIlWO1lQ1fpZCmL8yAk36nGOtcDlhmQpo10JslNeQI41524jLNWOLj51
kZaKGQbR6o0RxXqe03HSmmFZHUauk5tZ2GBOgEF4mm+G1ZzfMHtBhBUJB4+B
ahmzY1gM8qb59WbUp7756B3PBn9MWYUSDaukavTaeuqT36xt9IOqoGjZSVx6
qjen5eYe1SODTrGyYDQDtrnPUvLXq6yEzTRjW/uZHg0i/Op6iWPjTHCg5fTH
WWwIrG99P369koOxqA0JOV+df0ZCfL3zCysyjWyghIL/mzOCmCr1PUaly3T/
qeTXyqgR6kof77U02Ee2XecVvTjwYjUGk74RpqKKM7DG43ovZwYAfUu7VSvQ
ZNZpLGYYSx6ecICqQtJ7tqbuL/AxnLh8W1HbQG9E9se2cIEVVJLeYE7R5Q+g
2cFPBKjaCTvLj5yczM8koiw0p7cnNyYvX8sYiNJXwVIbJ1hA8AzUA5BDrWmG
ZmUEnTfANMwSYdlvRZsdh1ylr2+fZP3W0uzYezTH4gtv/S+mPs3KatGxkTfn
HOvZwjhwiLtdCoy0cV9qc0tQCUL9duKzYlZolyIuEqOrxrlPqkdw2UPjlApQ
iZWv0gSOhcqea6VngUM27NRIw47Ojw2Jwu6EQuApg1avzEVopUip74sadwz0
LBULYiv85uFa00nmKaeC7ySF3HOSOvGfm8JXh8l3KnxegiUXbGeRQ/rpI1vu
1eDF6uLj+jmMOQ9tCP84rQH31G5nqJCUcRu/tl1Lc/xIitm2WVdcHvv025Pj
qJHG51soUumV6X2JiZVovqmHKDMBvjV4F1vK0VeR7kj6DurUY7EivaEuofb/
Rx3id15SWljRiyRwU3sSp3uJdgUpdid414drq605mesOm09gVzN6znR50fN6
5B8iBdpDVo/JDOuodASvSGpjXyVdOoUPk5b0Jc89oytZd8dSOIKRE5hClPe5
Yck4Klh2CmanipnQpeyi9C2sCh6bP+HHJ6+j3YghDOfOaUKMidTBgXdeY99O
a3EaJkhfA3b6NJQPxJ/1JVoLCACjnlyKEO6xjQnAG9CXwHp5AA1xmel6xjfp
PEo6tm9C4RCUPr456sXyDNHy3zjX8Pk9nzr7Xj365pMISMVQuGp5j6Ygyguw
U4HNDax1Dzybu4Uhr5vbC0pk1pRMGyJglSZZpWfIqZ72csoc9UwhoIYaVJcJ
GtSel4bYTLQnp3AkO2IopAbUrMZ65C5Ld9Vj6VkeLWfCOLQptzUiMDokrQom
FNrUkoVmF+yzRjF1xL2elVpthdlOiMrgpgW3Jc+M5L7nyxrniWObEag09+64
8QdbjMLfZd2evnfSeNutfaG3YcXkADeaeQDafP0AQN2WXlT6pzhdcc1+BqnX
BxHuU1akb7EmhfSMvQO2wYZS0L2vX9v/6AKBHhuHQ/lQIa3qGnfRYHJcvBBE
pl8HdPjqP1P5r0Eqs0DI1FAbER/EaBiUDImPRGzgQM/PSctZMObaucFYfA3L
1OmoF9CvLnxtvWCJ+ZuVbkMOoTFZ3cpV69c869+zU6KCDXiyyqT10iQQhhYu
DhIepfF1QziEsYh+NQ7RqIVKRsfAFrI8Y8abLbFb8EBktrgzh0mX6swaLZq+
BKn/NFVQE2VdqEsraoHoleyDXjSTBo4ZvRNmJK53DFPEubmnrD23KP90HpuW
G0RC80vEG/pfSN4NlssFLvzzaep5P+3He2oMpw0HUyzYZGZcyjfDx9dw6WP2
x7L82ZA0HibmuSNn+MQwrz6wgkmSnu6/aKftyRETODdR2CUgW4MsuLdu4Xfs
5VsEuxTthHGY5V3Slqkx08g2Cu6G0vhx2It2BQfyKOZIKlx9x26ebouYEZi3
yXvql2+gY8qtRzanUMQV+k5buKXSo8jX4sokfeastYC4NH7V6wnojTWShBGz
XHLGXMh3taWu+4PpRV6Sv6vpj4w6IkVMcTclxIwkBThcBdAOgvBg4/HzdUGC
OLAnGVXhKdebFR6mzZiNjS45RBeXpSBrhR35NyoJ4yvYhH/ns5qzjxq0gMOe
BxUVP9FfMAInFgXBgOpqTixeTSNz+XThc4CWcoRP9pqDzpdHKzfY8AcYvhq0
foPMEQtI2JmRHCBD42KUrX7xQeUseNMjv5pe1VL+afSbZyAFeJr4B/w1Xsef
+JXE8d5F04qhPAt8s7uZcoO+vQp1xxsqjjo1v6/YzdwFUanYeky1t80Fs0xc
e5gDhmlAdxs2CENFMyKoW/dRgpgwKxVfvumR9s4A8GaXqFVtRapUTVVTc4Hd
xi5UwzTj3+E4aEqaCey47IXnllnJvfKn+m9Jom9YtF2qnFiGNpQ2NLAwSvmG
uSD22NJHwDKs8lxCYK4cz7FwcLsQC7FjlvhMqketXrZQWLIc8YlOheRjIkKD
kqy/LuQAqu9S3GCbPphx/ifkIeXU09MCWagXo0w+ZxjNygmbZuPwzeE/OTYV
aV4J6U3apnqVEb0JOf1J3owhGVISFonbqb0cG5DO/g2Ua+sn15PWh9pAJdUx
3cGNHnVdcF5d93SWI24Fh8iBAc0Z2rl+lcW3GGHt4Jb1fTP5gDRhieLZe4hA
lj2PvqgfOvrsikc8uMsYgJORnDqdFv5dPmsRkzvc5Ttnqk/08t4oHp6jfZdx
LyC250TOk9UO9Nzpv6fq09udMgku/G0mIt1E/TdLjrOklPNs5axpyb2uXMbN
du2tmB56EmZLapVE0z5QF3SPeyHJIuSGcwu3uBnngmTQ1IBtXdMQJInhdYuB
arrQazJN7wOgUSj2QaO/TaKiOH+q78Wu8aAcTmytA4/M7E0GuWoSYupby/Iw
iPChiyi9iZp6CIofDaOIXEfH2psppQqmMmylKxhe6YirY61brgNctbvz6SYX
DWyaahUIuxdb5c7lS1UW3ERtNoRf2D81k9iVaJBRJ7uzT1+hJWE0C4Lr3U7x
v2n0ItWQIMiDXuZQVAf+5N13yv1cWZG1862KGGdcDcZdUp5cTiJi1eeUUElA
JZRaphMSk+pKSAaAB8cPiJTTZ3zXiiPzwlcHsbvjKsAWM2GwFazHmCJp4ado
Cy38FVM1u8nMqrAagIQShBrIHakC8+B1rGwA8/e4gJTBmljzN6ypFOcgHFg8
CJWQj7Pq1jdsK5jwowKGegqs54eo/MWDan/eqyXVX657OCnt24RNA/V+q+tv
1q462wj3jpw3MCxeJ1XZdm80NGD8+Qzt7RkqTu/tVF0Or3P6v885wYu0DobZ
EfkH7xNoK9ozsUaoBlkhzfzGB/vwOHu/pE7BV/37Vc4vlpoIPfRxf4j6C9wF
7CuT49HEf/ig7/+4gkAHw1kJbUjG6KsP7tAwa7q974X+qdn4kiDeKYlcP++f
O45jqZzvcHWv1ZiBjLr5obqJguh+4CfD2lq/euejxhPBu9T9PCOkPWesVey9
jV/m57fiUHpQVDedddNBqzkQKWgQ/c4mcTaV3XfiWf73KyaZeqZNv3wIbg02
ys49WoTMNAXsg7V1DKxn3rzB3ARAlw+gDMFA05mFESizAv3ZAtU1qqs0kKY4
m2sMhqaVLeIW5fAovNCLvbhJsSOGJZrqJ+SZddMPy3YcF9gW4G/08qXvOVR1
+o0myEf0g/Y4Npqt7Vd7qXpVPcWZnxASFK8RlhDQVcQOPwpdEYdmJWIaLjBw
C1iWT81uVXiPfgvEipwJ6ezgauFisWfAmEJ6qf3hzCKl9MLSr3w2dm0Bo/gm
dCymPIGnLVKvZ5Ac4RN+nMmgvzMvwkjjyhQQ19thHgayE05EzBo+m7GxOYts
1yuJaLyavxvkQXRdsSUCcrUcK+ONcnuFSuAn91bC5WKgwOQ8mDdjAOahNiRV
PTaarAesH/EH5qBmQgcfXu/697KXtzb0jSB/vjvt4aZ5PIeeSAZf25MWTR2K
9wlPV1wONkZTLXKamGjbJ0xKmGYlEoOXsfPJTqToJR/VUfuDul+P0XiZM3x0
rUDkyoUBn+Eb6jhVf+eoTZmZtpJ01QBBSwXo2Kdr9XKxdvcRXOUwHJu5o+zd
CUK2QjszrYgrDRLVmTwA1a2DhuJ819NzuulgaGdiQQGYJWXt74OZCGeugHdi
ah6epxdXsqmHnhuGvOrqDs/AQHHZaxV8qtVoJb13KFqlulzLCwz9sydzckFo
nj+jfELmZ+kbtZeXQriPnTP0QUfdD8O8o/fwmIixzaQtjteG+KEYqniT/pHg
z5Xn1NwWOyHiAdoHZKY+yVounMd+GaQC+VA9wPDRJuvAZ/zpMbkCCkHnho2D
1o1AiBMH4JC0KN+IJCxXEgmHeWsxGQEShg2LK3A88NEqEdTAXfOqSevbihma
e/eOq7wOq7RNGM2GTOokffFxrvFaiXsKtM+/FwsVbq3W/onpNBaXolUrbIpd
SUPV0HppIruQnXtNbfrHTUo9Ru/n1W7y/bFZrv6ECyPP0SxV/6WK1BCn4G8m
C1E/3yOyQuIJ3s4WWdSFfFB9x+NWhI3qU8sCVg4u+rugib6axzIUeY1iWxlg
Qayt0vvq+nDuqDB4R2ZCqQZwL5I3hjzw/ab5MtCFZdwtemnNqOeZa885SfKN
hYw52HlGc+X0EgSDvDxRR5fvIDe77RvYsVVM1a/OVpK0hqF07V9on58iT90v
TH8WjgP9pB9ztJ68GhGuHGKPNQHflXqcrcK7A+wiRKoDY1i7TLU4IwwoXTuC
FbaalaRK/HMfyt6pFa+Ztpq/aRk3Lb8a3DhRvEB/i6zN9+Kotp4PF31WU5dX
dnyXhKOqW4mwu3I/0XypALh0/u60OQCy848VpEv2Fbe+MgRw1e/glgWaj5fz
0095r+uJ2k25h1CK8Y3dNK3UobWPOedzjfVPIX7ytvfLgqBcR+aDIU96zjV3
UlgzK8l58wiDxMCCjXTl8rs2yl++UHavM0pj2GL4W52v/EDrptFNBZ09Vu4q
TGk3OzJdv3FsvvY29YUQrkV1HM2jyrKq3XqFLAg+Mcac9aVZBx5vZvQLe52f
KwpXwpUfGYfikuLp9aeOo9zshFE+0o7kemxgmx2/gJFiRkWH4K+O0xSjGuot
TA+APKVVp3h2qsT27Yafy3FwfgZT4VAsZSj6VfYfmb/LdV06H/g7lCEj0xAb
fezshNz/WHIWzTTpwW/aLAfsf9VoUwncr6ICUQX7zLqDL+OmP2b02C9Yv1J2
Pc1LyzVlcrJ3COWjzGgtwYTQ7Vf35cXZEWcpU/uxSrnBnPHiIafas1FVuYrv
MxghZoKvGlMQgtOB1/IfxYQNEnEULIqLqmXw4sYMZjkkPPf2rOjXByZh+Yv5
uMJY/Pd04o2fKcUlSntcMKyFLKOhmuXLfuaDAhPJ7YPgy/EwbyG4hwTxp0GM
CZcUBaOoCZ48P81OBcLMPtcj3FWx8zlzecn1rUcBe3nc4CjeP+Iqavx+mw+V
BsM4R9UuK0VbO2w0UIKTP81Nbh3lKFHUfgGdzAJNfrMKGhUumDyfWIHN/Q3o
/+bpUiSzQAATX7VDRZldXfWYbxD0Yw2toqmZmauSKsU5bv13ZdrJ2NOgZcVS
cHWrmF6lRMbJbAx7/4y3BNi6brkQewJulwaiNQtoJpn/iMZPbRhCl5k3KD6O
kyhRglsXu9joZm4cEKVxoO2O2IyHDAjT9riY+64AqJvTLty2ceBM4A8flHnH
yD8CcuntZiCvt2m8TNJDvdRNqqB4iBHJJFMulDnJ9U4wm+BOHvDN3RwOZFPJ
jEphQUN5S9VYnQnaIYgMTWsOUuAGneN2x3ykg/IiTtUiWwLWMhIiZwmaknuL
679Rkonplpc1JrrapAesfT/AH68Gw0dc7puduA0kyj0tlT1HB+NQbN0G6fSK
ojonbUfolbE88us73yszzDQT9bKxrpsgbUhD8DYqWssH7v5c90LjpZjrtnVO
wcVAqsJJcAOdhf7dDq2Emxpgu9EjovaS2c+GvpjUkCJyJFDz2/u1+t2KV1uL
Icel+x+quP57PP74ETmo7AFLPypatXwRJ/0zFZzNWZjR7OMwwxDv1SI/Yosh
IFHZEmE00yP0xfa1jPxjR/1S4UKdmooxVCas4uBOtWTMVl/0899qbNbl4R5n
5i/Ytc2QEBESAEDKm9uYuuyGYiI/aymLwsDF5GxOL7It95q1TSxSRTB5fP6a
QtSbwQfw0CCP6ccLZOtQi6gGX54yjQMyz/aWQTfXHQ1GR3ELkXnLyui+3t8H
qa/IvRLToYLJ37Vhf3BsW2TbR2iG60K6S4aBE+sEEuQlArVlCgve12SMVRYk
qPNOYWzCBSfberz7mre5NdZKj/svtB514Q5EkrY03ogoTd5xW8rHSi7rTp6a
/p8H8dQqKoL/ZNB3aZ3MfgyjU+dIWygJt/OfPfkocqfzLA/YzbZLsk7Nztpz
GBEACjzdim9Cufok6RBRlvZejw+wkuBUTPVuHPp2OllYKGyJJ6BKvADx4Jp8
aRkVpnaCRRWkqP4PdBNHcVPQsfB+gwLk40RL0HmV/14m7HNcGgsGcR1SLCZi
qOQGu8491iyJuaS5iqQ2UDdoEYrLWGRtLcP4mOvmcyyhkTdK0vZuIjmoqRwq
2vtTyhwRQpYPMXY4mzdCEWPp5VMk4RN9Pe45PgqU40P55uc01em3PhxLAKad
qx3Z68Yr1j663mjFnfAONvjjA/PzzqqMe2NkthgX1v2AQqwGfAECg9h4hYiD
eHXAftaCrojqC1yWBiVMMUha2licjsCw7RaSH26CPoQh7GARCcNkJOel2Xhm
6dk+Pv74UdwKHAnkHr62GYLF5TFwqhC2tG7P7tX6uSw7ijcnhcj8jXc9cOX+
ZYg8kGl4lTYLvJ16NeQITFcCQlETE8NQZYNqWMwot/G51HMslBlLVvgnjWZW
2KHq6y68yf+Zhoeglsb6N2HmnXLeEVUVyzN5LRZXpbkfbKtB77NA61d95xVn
sJqBIDTVmQ5XeZLFTbW5fiTsrgFneCMvvIc4f3PXuSMAV9qJlcqoAhvmHxGP
yYCqdvb/zb2dctF2HzRhT5rf8l/b3y5dmYa7NnBPAp26JbCPqepdpqfXgQWv
SmPCgSpS2v4FiOcq//zrr4rIZnSridE8CWxuY1vfGEclduacoJzrL7pOFz6k
5vhUkUdt5gm26qxW9JLBVlczLLdBYturptvV1jGHnNalXtF8cPshvgyGkb5N
Xh6pgSVKWW+5eFBrFA2+xR330kpw+Ldh9vlKlB0qiYvUfBsi0ZcJOZRP3MJi
iKQHl5kVah2i22D+GecZcdAYsxWQALqadoGHq/5DvnJxqi2RfwbOgHf2DCH6
I0Slwz+Sb/wb1HAzYM3CjGsEGzSvDLrg3/EeZiroDgd0DyFktRN6J7uI4iPX
/8naMVvK8v6bNE5uR4Whv+xlbA7/f0LLeE/uHKBOKx2gndMeRqP4eL6PBhJy
p7SRh1Wleb5zl8zaqyY+LBX+oZ369Y4BPRWNs3pAPOIzLrSERnM5ipW2Grv4
wtzxvzjWzlHHRlonWZkjYnd0sHI5yySwTqmDrSv3o/bc8+tARqAILHtF2gO/
55g+gQLfHl5v4tiL5BLhTn6n8aBrvVyy0F5xsFYuq9ZItOqaUyAD30CtBwCg
QF7l9+KMfMe/+sk0IsXQzC5u4OX44qvLaJiaVqtW4Ej+6eXZnnOxm6VU9UEQ
QDmfBbhd+COSQcnkMFjZvhNfS7WCepTxePmu6NIi1yBwIZ7GmS/WPMePb4Wm
LeGL4/z7XsG5ob/fOzLWKVXWYjNtq7vbfle3OkqMSOxokfvW38Yr1aIMNWG0
C5qqRRpjyHUcm5XsxwuyI/3+seG04nUZOYM30JsSDf/iDI/76QMjxhxyp9QI
rQ7JrGT2xA7MJ3MCf6xS1WK9MV7WPMDBU0pnKXzTVtDmOzKkl0SWqkTvQZ2Y
12TqUZhVCXUiJ2o26p0YkxZpfNINxUgc9/NO9dbA4PRtr0c5aE1CLA46Cb/0
1alBNsAnMPd9DFoJWl8OjWyHognf5oHgbQ206Tz2dDaBF+RsZnL0ihFuEZMe
upeR1L9HcZFd6I4WT0FBDMWWwxPSXreg5S5uwVIrNNz1BYJb7IGzsQT+ycji
fdlDuNYlmGeq8IkvTdN+zuWHsa3UXKWBpcvXiDhFloo/URd0Abi1hteUegdS
8CXtdo+lQi1Uss8YJnbnoH7fjZ13uXzRjElhhU6rhzFc8S3DMcVwf9NLHiI7
myfht+04t1vIhzYE8y3MaSBH6i83INVBWtC6+SDH1ir8vF/t2AaVukJmf91i
klfppHJWgrzXQ8NHFZsyM/kHYrrYYZmQKrCYZiPJug3u1/3TBnY53Ixv4Gmc
Q9f8Is0KhazGMVgBcrV9CD/dwfySAA8EgMyNY3SL5VIRovyA5qjPu4x19VOu
OCO5IGylKgpZfsJCMlDjyZAEn6635llLLM4gDznzHeW3ATRH63Fvrq/yLLlY
Pn9iuoyh3sJB1DpmLuv1ZdCXCNtAApf5iS0p66CFwr6WLmk8H64x/fb8IUbj
OKOZ1w5yKM7oogQ91Lv4xsZ0hqJ0Aa0hYoNPnTO/XnvPWSi3mYD+TuVA3rEr
BzCnonkCqHxqMT7UgjNOLAaK5w1Md6faxNXwIRSSn4rBzP8dtZSSHbSVgSED
t1OwswnVNCOGn46fm7cWCK8C5FpNVQydafeO/szrdZO2sjok5Qi8jZ5lXNYQ
wpXYPdVmC1tODD2w5tIGggGo5LCMCMtvuDsYqkWczujJH7jolL/4nSfQNlnV
Cf6DfFwFbjmNlU4MPfHhIDBlKub1O1TxA5AQCzlL1qHD6F/lxYMyWSR67iiY
9nsnfjdEdnDYcrwU19UKvD8adIhgfHpVbhACCcfiPRKnQ9DuEURkM3VpUvhI
T1/1lN1YRBM7TMV8csjQOvFHqWP5zQMWHCK+M0nIhlEBMjgZp5Uv/Xo+Q5gU
YEZPOaDFq8PiFVcH8Hy+3UIFCq+TA9ZT6juHQNC7RocFpI2uXeSR1OBBAIYu
sVR5e7mxoYtNq2tRTxE8VaDN1lzbMDpN3CPWeo4Dixx+UdK75nDq/Tz51YVP
kdS5RGgf5CvKfFZBpwBMd5NESTo89M7ceqqC0yoOKaqqKF3S3rL6xuz9yihm
WyqyvuLbPkaAg1QibLnoaQRgt58nMCzMBHJUkc6C3DlrYqhnv0f+MBuCMdvt
/DjHW8BvwIj475MnZopvwFtcQCyVAYJ4VcfJvi4CDQ3TvfRNe7yfDA9D053Z
TBe5E8y6Pkt8ISjk+VkCl4xV2tNSMa3Nq00VfELRX2q10h+hBBDOwrnFyavz
bWLSacdWKz/AvY+VGeMLyU0pjjsYpG/i57Q5RRh8eKRPeZsBxMm6gGVd3uSW
4rG4EUlRiO4MCuNS1l3TvYJ9ikhpnrtkOyTHIfRmz+2G+G595YpZ/OzfcWxI
cw6hW36cICHsLsRNAOqRq1o6T7XsMWTZy6wyJMeh74aVJ2LmwHIsj0E6kYzn
jRHjuYo4hOMfbQyIZiCwQ8V+KpsqKjvUUeLXUETNB0XiTCH06cR4pejzclxo
r0RUtyVNpCfO/C35Ij7z2heXGy5VBWfE0oo/iWxyIbxCW9wZSUvxKKYEpp3d
KyNPWteojRJ1jy4xMCWTHhk4BklPZRMclIZqO7/DZG7Xr6PC9kUVZS+oda0e
+QS/nq6rYl1GEMpugweKriChDSO5VMFgN5K0t5UfNSDNJUc9JoUpncjSj8nP
lksMyAk9yUDh41PdpAuiwC0TZ/6Xdf7wUKZcZyQ+UQFXC/c13krIZ+dEJvJ2
fNhkEzpXOLDqrEElRB3AAkPyakDJCxrsfB7yTxSsKDCRe2PX3AVKafsE6Jd/
IAEv0fQVsr2THBkqTYq78wAs3L3rCsJGUaOBSEMoU3FZyveAMN96X5aLKYFo
M8UroK7YD72gAhefnDr0avx9sX0qGE8RyERGD/WkkJMtmnO0Sz3/g5GK9wfB
+unXu4epdq7Q/yvzq0O1hXNeQZGhNnPo8DT/80bd2OF/R64r74niaZ0y5Pjx
TVPP52xfwo5UvFjuUq3kQpXIJeXMe/8vN4xkuzhOLSm8eBTU9r6w7u3zN4tU
wyOu8+PFVFLVJTr4L6r73hplw0Gb61kma0fMFKoCZ2CClxfwLj2Z3yiuYDPg
TpujR2Qfx38saCe2ccbblet7H+xkQuGHIkzv5ZaF0y3XQr29rBME2qlD5se0
HMRrpb8umFaAcxLF6d++UKsjVb2/xspPbVFX8TF/PDNl1eTSYydxochXWsGc
9QAWdHRy/jfqi5TMishkktBzyXj4VLiV2czBcoMEplYAluuc2ldzpFNxNyIz
dj+7Hc2DbRB8Mt73A4D9FHgNPtzepLuDbFyPaojMSVfy9GQZ2xBVC1ZhbhA0
ciwP7kpJzyZOqPcbLDFoOV2vPkw5hXi7Lfrr5SGwaWzUYBZcFXkYRh2a0Z3V
HbuEIgN/bkE8E0hf9XLwqo0l+LAAI5FWUZo1ihBb74EYdPLCdRPHlRqrWYxu
B+YOIyX2iYYzpFfbrmdrlf+SaPuII/cYhxp58LE21WW1HqrXAv+lFy9QofFH
c3h1pH+DpwD45yeXDEYV/5qSybv+ghvcGGT4XFauTnb0xiEmCq/JkySDOZWy
nJyKDG9c0d/LQKhQlf3jfZldtEmlaBAGOLdEk0QTdTm9PTc1mjh13fJ/P+PX
HtCWaKysWEdmXq0UQ4r2bIjZqUh0tkSbjB0S/gmmSP6sMJJF/mHOqncPnPzY
1XdbjBo5t2A0A/Mcl9yWNxz9j01HZ0wmdfXwSEoLFPfm6Uxq2hxvwQEXQ0B2
RfuaAnwTPl8+7S3d9Nkbd4Sk+nYuCULxG3RRP2e2B3yJ6JSMCJANNc7/+0Q2
CBqGo5wLPHfuprwBFnOTpQqX5e+6qPooidd3Q/f/QDBgndyf8KdR/CnIF6uU
NOZe9O77QZTT8CuTpmEBt1p91En3QO0OB+cpB2U3a6pMbtGcRKkfz5cWFpEZ
YES3DENCjEoVrI1YTmURaFtqGfFVSu082Xa/o29A1yo0XiXgdlq6MwIPMvCC
TqSzA8TN7b6wxECixomdXZKPjGymOtGEl7VpZ/jRlqflQoD/uc3Zhef6pI52
SPIAnclTnLCmotxlRA88wsb5qEi9s2bI9I5yMP2wwAUjz2rDQ4fARSrPK73Z
0y05oBp4Fymbr188MPm5BU/c2jBlKrZkp3jtkbyh2Nb3l+L1nAUrhp+yTi3+
zf3EW4wLDwEPjdeXsCpaQRrEfGL8V7tdBf+oCP+Bi4rTTvRUgABQKLNM9Lt4
5XEIzl88T9Zij+en00Cr2ptu+JQ1FDC89gVjftd/46eX+DrPZnswfo40r5lb
bzMPY1nTyGEr64tnf94m3LT1WOnjfiYsZi0ROOfBw56sSIKL9Pm1ojMfelhQ
j0grVU4vdICPJOihlWvNvJ9Kjx7J0uyMiOgHTyx/ytqHvIeUTowcR4catH0/
oA2BhNaeF8xJCvn4ey5cz5aTWOwTQs8L3Nfk0x2WfZ/0VoUg7BJM8M5ImX4k
bWZXnAdnZZ9pJErcUt3IPIZbg/18alUPVYwB4aMUziPYzhdcB8vr3ZObYLq4
beqNcjRWdCOZS5o0K9ulxq7dSgnc07ReAAKG9d7Jawn+eIXXZ/2eGg9tlfUO
DluR+ioYtx/9Ng3YWDy6qzx1AuTeU0GVHv6LAVpWqF+55Bwi0L0iCjITEWyD
RGNQQS6ttU3wQthPoE1KhHN77JgspAlfI6hBeEvtoHgq1FU082DNrZp0zSKY
iWkqqi2AdG+UfDnK+mM0OMT3XWjTZX2I0cvAyjHY/nDuMg9OSpj4srTtNFd4
xkWkfRLJ1YhKPZXRpYGa7mCYC6RkOrwKFc00CZzQGHT04lOT7O774iSgMFwy
9gP/7bbls4mPjiDhOAyJzg1uKI/Ia9U3RIbicrNf9NaiuZpGBSzM6ZQTl1gX
6RCLaA6J31SAyg5/zYFI6p0mRE3WYs9HJVQHvZf9AhI9y5WLzG3K2myap7nK
zpUbdxBoSEOvCAkqBjgHRMC63UM/EO6lp2trdR7R8+teBRn0/7dU4Md6/0WI
G9ze0l0xGNm75zB6j8GuNMezfz6IOetqhREwafgnzsgQ8S2RiV60oXcq2vEp
L8+ABpexuOxsS17IcVUptMHGBBBVP9oUEotbnTXOqyGTnCSVdfgK+IsIIJcs
/Wwl5lI1ZGCgs+IveqyODLIQaayWfZMd7/+tBjmYQHqNYoX7E5j5khGtYI7j
VoQQP469Z+0MUu6JCmKytDPVH1BN4ImuTeDHv+yaQ6dRfFvHaIAbl9MGsxgA
tgbuvyktb6vHZlUrsj4ab2GLKwQzXINC6LpKcn/il3lZzQffJWKnPRc+hrfM
f25zuPWsGoLsfZodFy+k3S8H0ruG975gRiIHh/teqAlYsDk25ig0UK4II5ie
OWSfyIh6/u6fZ4sellcGWr3glnkpjeBAFMgWo238h8T70B9Nsgi7NPwKsSXz
H2yGINh1JFwZ0sGd1jM5PnTP1bXTlr7fVRV60X8lv7sTfkZOYrMigYprHYzg
ng4/AIB66l7yifMygxZVcnA6SrgGrWs+uzIFdJU+yLUvIz4XPEHd+QU69mtx
8Mc397KaocggGgGgsAruEvBL/CCKpO9PCB6afKeUoR8IpRV0138gH4nTzN9g
Zr97TeLoNyw1aNSATFjL6RrlzpRb6Xc9EgFz626pc0WGOdCQo93XihU9J32a
8M1yTxr/eSKbCugJrvQvGZ6UAsAESZTsrdhtca+f0vVq5sV6xhjyJS7tb/Au
Rcy9k6/H9SXP1yx4o/apIY+ITRAXK2jQ2GtzueBtMtD8ziTLBmmovvUgd1Na
M9jPIGYtV0mJrMwXbz8Q+FfkCi+m5/ejxJAFcDi41ZgnHS0rw2HtgtRpvI2k
obyipNWZl1Lj/vwfmC4aSChvfo4pr+FWXdol6oW6fnpDYszS/cbnmyRcXjLb
Y5JpAy1bcbNfAD08pgYEP+YGXeJ/klbDcvdeiUnscae3qJAtSmLXFbHtQnBZ
31HZzcBmXIpJ0l+vmihbXGhoXwu2QIZ/0sKGIzTJ1SvJRe6kgqIINsAIHzi8
rZjZdV3FiQ7v2cbh9F492afIKBhWJ3rxylC6QAOlBaofN3bm7+0aKhqnbSAv
bZCj8klfKuVC1zaT0roY6dPqRGaAvsxEW8l6fwBdWQsggQjwALGidt3Nfiz8
KIrqI7NZbMPQ3fjkux7WDAI6CC+IyXElc8oIRVW1rGG8hKCp0WFEJlWkZCDu
hUfRAQa3+GQCkgvibrRdYR/RdvGXtyz5AqQ422YM3MqU8mv64OJIT+tFiNJk
hwLHh0AR3tpFsu48LNwbPmUuphddtb/338pD1SwkozjpRPMiPpx0IbgOQq88
iNqftdhkadi12TEwCMVTopukws1PaOMVzfnXVxV7O2oC7fSR8UL/6vQV3mx+
k/2OAufHH3VijumvuXpcQAlTwhSD+FCBIflBFLrrQVUfapycvTeC8C09gkpP
rQlSryaNR3sVJLpBDXPK0DmKPF+BD8mLbdyaMPI9GAZhs3JmIcXM9fPnjVxY
itGJhIIL9X8cOS1DGfna12lfvjU77WKAEL+ZtGM3CJAa23WwBvqT/yGU9/X1
tLznIPCZkMXzNQ9geftZ4zYWpUNuypg2575rn2131dDA73KGYJ15ZRWoqcsA
WzSvaqucRNxnTWQQJcZosFsGgddk2Qfx9olfmvI2aBIrmUxtfpBXGm11GUCj
XHj/7cuqkWagloTJnAEJW6v3HNf9aNR2RO9ymxn4Mk44K5Ft7EIxAZAlqF6e
b51EPb7LTCO3hZJvvG/yZgVOU3tzfS9YSKJ+7NBzd+tqALRpzNBe5QXzkMPb
UTlWAjW85GHrd6kaMAH7ht0JD7BYoAZM9DN1r/L5e+6VY0aojPiB2qhZ+FWE
ydPhCDylpLueccSouOaPSzJ/TbGdC11OKxZWAXkXivaT+ylgt0PLJJRgtUoD
1KmFXfjBQTSYLwQIaS0AOGEKZNduR5KbWkhiCMC5bSf84S1ovXjWKoJXQXxi
9Z8F2E+WbkXHZlLUXAboZayc4rFKYNqA/Oukjc4CHYu2sk1uSBssVAFw03+D
mUra/+3KdNTfmYtFeXljtU/4lSLQr/5EGRlyzjZSbZ/Iaihm4Vq3oVZ6EPtW
vEuntQ7viDW2j8uNsPpwQd2kkBrw/kUJSD6V2ZcBykLzC0QqGtufiDNTzSjQ
88s/ZdYlWnRUHDrhsbyBd9R0Bl+nqUphfSVHOoYxArKr90nXW5rRUHkT8jK4
nqYWtzrcH6lguERY8C94RziK/VYKBmSO+bM7Tu81BtDNVFN3mNw52aWu2K5J
tiV7LBA7VKMiqMysOCly5/Udp4ySnvLpH3m8uiSTZiGslyk4NEc5EMmgntmz
3tLjbYc7CbVjMndqw/jm9sbfRQsJC8PvqY8cNhJyCUofrLS66rb4S4mWwcJt
Qlm9q2SmcHm8o/T5O8BZ8HXWVLseAU/1TjsC0n7hlwBcJP23n0LE0f51HJRP
s/mJ/qQDX2Dwes5XR33wiH/vH1LzSTsdmLc8wsvE9oipxKQXO3qnf67lKFse
dTtOGrV5fn0PHIZQ2BX+iISY3VecT/i/KLL0W68Kxa8OWOcwnycrc8BFfHqV
GI2H5vCUzuFjCeqhjiydYdzN3CRUCFj3m+FPSuNBxfQCd1ujeA3W15HgS/v3
dG/w4ELlRWlI4u0Y8Y+/PCAnSNaYDVM4Y1Ny76B3/zWgGkJqbTyPGS7dMxnx
ZwKpaidUXa34UWBhIGQrXOQClPYBTZdaLn9t8Lktzm6SfOzq6rynf+YihDef
TFsX3QVTKFHZ8TutckI86fpfBlZ0j2p5rK8ALNgS1jRuM9G1Ns/q8Miz7qmA
uGvLIGnDEvtzI+oJ8VnvrYwH/7DtigtmehsXPDOKlTL7Kow511vhiSo1F9FJ
zRZbp9Vt/78bva3vDQhXtXMeZyLLYjZqFklG6j+9Wm6L/PR8Sw/WEhmPgyw6
1KcOM9kOtqsLyw1gn9Lrw+IApCepZYF22e+z9lj60XYUf7eIWbiwtp6KE6mX
0Jt9H3a1Oh+XFQ4JOA/5crf0SEgVM21xTbvz0Wfszybym3jOnRf5at1WOAwz
F/LDHIhdeIHNG1h/itxKacr1dEOGxzaAzDvnktkEsgrUirtRNvYPvvXZbZeC
CJrfdpWIVkOo89HT3XPopjCljuDQmluSsCUQCjHkKrql4AjsZWDwLxQBNOzV
OCPrZRA8+Z8DFssASKQqckCeRyyRdLODWGXPPUa9iDortTj1LNMyETfcjtiO
V1j52BWEMIYQGAiRsK+oS9WImFWSkA4xIToLKWlHsad/+p6fy6SAR9Lh74jZ
KuDxZ1LgIEG01VrEmbTmJBPlH+KWghM+b2TvGvTXc9WaS21rHmTnn3K4B7px
Nc5OjXb9IA2L/zrzBNSxBE5gp8SgV7zm5yL8m+J0e34obu8b2MS24x85tXXN
k0WcNX+rO3p6r+kx/AokvzEgZl+gGIj6NEkYNC9JX2MQTMtrEsdEdKL11VOC
Oplg3dK7Ymz24zdz2DwEDzf5BlR6DMroHktC0z1x0Ic5WKwIm1wiPPago6Pg
IwBXqQ3IAiFKUUes6anxCCpOnBoVjAcDjHRtYDVhxVVAy71XACbV6TQejqOW
jRkZEuR69aoVOMTH/gjzLkarZsZ43wHfszLkIks+T+0jVwofqrWtjV4k2toe
SwkEEUNcFlsIYUhz4/FqIBNoEdF15E36/UDHP/bFTJs86JJ8IgZTIEOFLzf3
uxVzE+Wo/oYB4q9WUt8cZUDbA6+sqVBDrr8pv3u6bXadA3+Fc5EZmk7sCRgW
v90vwa9LyWADPKF/xoqvIuCUCcez+eENrciaX84Vms/Q+NsJKA76LXlYwOAB
JdBjUwXa4S+ttzPfjHe+cGVLkizsKjiIKY/oRRf7af/FCiDDHCA+l8MOrtiP
w5KDEd5LsFH/CwHaAvLypYtUFhV03ndEKR2Ic9iQwDQ2g/f87fqdNVSnWMqc
VWN2r+1py6oUMh7/Bap1wnQ1g/yHRYpT67Vz1BG00PaYzvIcx5PZnAAGmDNh
Ot8ZxmTZNyOTFuZeJv8r/L4fgJKXPaWxWrXwbuUv++pB1powPnnuVgqWqAo7
G/QPBTyRqbI8uhT/HetQP6tgjuc0fNGlyByPXpyBPBQcHVT8I7B0rSzz/xzI
YJv5x9Agtie7bws7aDAUgBvYn+fZOzeGi0OHikmZ1va9jozniw4/g1utIjRL
kTceOVufOAnWxYeP3LBJUc+i28y5baGRmsSyBwpHtVXxhG3kgoE5BESyIVSh
rqL6Wm6tuTNMh2h1fWxwNxKBobbvRvBpQYCTpxWfM1qncZgqIOLZUou0VU2l
TZsVe6wMiysXp9EtqQ6Mm2qcShieSc5WNFOlidQ0dcaYH64n4nh9gfMDcbHX
EA6gIoOSUB9pmd+LudWIdgUIaTd8oUlqe34qXMnvMsUoYF09YELS9wSYEtem
6Clc3C0aZe1oTekoAzB0u+YTtpuhuoQfr0LQk5/YIUYgJ0ZQyRWQ3Ya8R2+3
UdPBVOVqNpb1SIkSagbgM4IpTSaGxPG7JhN5+tAKIGgi4KovVcTV1ogZamzk
klCUkBmtLgxBRn1xed3qGMiFrXfDuyjnrKl2Yo0nX/oZgYr13djp9jVsuNo4
bKIWx20w06Dpq6n5xd6DyJkZnWPwGteceNAPbio3S7grd46STsACAbMKLOcP
JWanK/THCh6A9EHizileiUKpmcG845UB0NnNiEHLUVKyI0ghT5hyHvDN7xrY
IT6pv+UEl1D3xIbRuFCRJrdw6+zcVP7A7b7A9KLxRQoAHpK9IdVCz8JeFD4M
vHWe4aDCGGcIUdygoOZff20MM20HgMq4eCC+xZDiLaD1XXxTF6CTxlzE8ehb
l4uk0GHSNxf0+yapa+jbTN3mLNGAYR4jzUJXAvdfhuZFhCtK+L0gTEBifjtq
XH25M5AcqfYbOZk1dfVKyj8+gQ1mrL6nESw2q+EFLbtwdgGrtaHhKJa1LhGV
0WwojQGUGdeYnNmQbriGOjRWMH3mh2mGMp6RSGVt77vbCgjxlYrGx2wlboT6
btzrsnd8CxZuL2tN50tF3pM+reTZvIa0AH7aFv/DKmVyuzZme98du4deWxdM
ieCsdaHxrJIN4/g9fBfqP3pgEDOUSKEGyOd6fP0TbvsVq5NPkpRuM5bReTxR
Axy4KV3l+ClcBNJFlp7ET2NEcdKeDwNTKq8Tad5/SM1YA6V28pg860CL6RLm
WdBY5O746qmDtpy8dl6irmn/f7qJ8OyGki4EHRlCwzn+ig+RE9cR3vRM+EmL
Em08rbg2r+yhWBr08OmMwXMEyHZsRyCpOilJbx4uxU3uwRsbRlZkbJDqzO1I
q5PFJaRaEB946p+zpxE5eeVOB9aqFWPp4aQ2iiLWf6mB+OCcZti408TommgY
DFhOXDpVT0V7zGJEDWYtbtUD0DLe2FqoIh1TkMmZt+UoQST0pTpER4+RUyKo
+JoW326dKFuc/TgOXXwMxILwJP9VcKBVItHgwdQHWTSVGJMNxIQObTyPj9Ti
2CIs1uGWMxvYCtgjfbiE1GYBkoTK2cXgD1raOVdJR07thEwk2Qb52C8nVbuA
81Ok8eZ8II2YLpvUSYvbeb8roEZK+7S6eyyCSRWc976bO+coUtM8TZh4N3V6
PvQM+ndlgsRmpmuBcMolm3QK2HCCQFSxcQ9iFn1yDaOF9tugNPB3ndYB26KW
ppWTqk+qSjAoP33PLjWJG5iW5GN8zLLgZjkeYUKX6wuT2XIUEGy8ZaoIJ4JG
D3gjnzXqjWgKxULD2JxZDMf3YdG6m5+SyDmzyjn3lj2vS0ajGBb51rkNrT05
8DYcCnjx21JM+MgpPgf+gIeogGa52nsajXGUewYBhB/tyBo0X1CL453Q8RAX
3fGpTxssQu/j5J+OvqdBy4T+WH39FPUn/fYdOTcKMm+7r3fhQidNsYhw42Dz
HIx+vGUzjOwMc3gAsxJChFhNzyzYEBrsjH3lYx06KGSWduIEyuvWxMo3ut9I
UFqUdc2lhrsek8w4Ng5XXeX6wP6wXZ+zpqDu9I6zpxSPYJsBxAjDHhNYamHD
qeXYW4uJpNR8dZ6zAQuZEzUorkMxevPu9tH7OappKib+YexDdkaaR8xX9Ovs
V6jpeR2OBZ+BTDV4vhYgu4jOFIv9PyY3RWcgvBlP0Rb4VrTosLyrtr8Iwmud
BaGWD4j+hpQplmlHSZ3esahC5ZEP+Nu6EDmh/sc1ec97lpaBbqP5vyOc8iTJ
8b6ItEGfWOkAatIwwttX5SLOP0zhY4R18N/SKQlx/OvoeVNNYu3GiWMP0tm2
cLP+u9OZppwOQjsL/sKFNqqG8RvHhQ0roGzMcKcnNQ7+R9mYKqqfBcp/OKgq
fkd+Pe4Dfk2g2yBHxlru98qEBwjw6TjIc5ftO7csAvOV9jIDNJR+eSoppj7z
gLbPQXUMwcLm0V+4Y873xnOSxuoDHrP0hHiCPMLFfeYkdjJa8G+0EBejptjD
5/vV5Vy8cfSrLIkaDawOgpBbthGFy8zVhOtq6nmbbs1Zz+zSCvO3DOX0f9w9
RaVzE2SH30nRtl3rJxcVTHZRoTtnsQYyMJM1jyW7Y2CY8oRY0NQg/YGOL6av
cFqbJvpo9vdZcWFqF77Ewi5aNBUy+tfGNK003W3fLVKQ77LmGJkJkFqsZLI7
liD8RYN7RtFGeR4rYG9+S45SolUpbGO28kXfJsbH1QXkcdrHXsZNXiuRLMAv
xi/KH3FmWEOIrOgSQPqvWwvaWir2O5nlNUScG+qGFGkxagPscE0jHA5QHsD/
lCXjed8IbeXF8rcqHz8sPWUkUTXhj0QBAtnP+Mwyj4AWmq/pYI8Yu553GrgQ
Fuwh57Ve1ve5QB3OeBPslLKA8N7cU4K8aM4KPnLSu1//vpC1c6UX36J35aA0
a93abQ2Rj2NA0eAMA/SXfpn9Z8B7JHUQVj+qb+90fBznSAr60dO+1g8aa5M5
FNVlKJ9kYBg+/EkiGbALXeTOHcuAfxskOnzPu4e3kQ5C5644ybdDOu0x/BXx
pOv7ozkR6j2/c/N8hBDJLK0VZP4bd16BSEi7slbmmeoWAsSidX9feoMgVy62
fNbLKzPdZTAibU9n9OPuMfR1yZ6nXg2X6R3LHiV92TGWLEm4eG12HiE9h3lY
/s94p+OtcdSCrOWAHlOOtttwTdqRN/gOw36cjwOY2n9SDu3doCcbFjv4cJQn
olPNAONGaRTK3an7gWDHWopGM14znUH59N+wgLoAoTpT27FHZZJbeZlnvI1i
hLpUWq0Farmjnhwv7ptKHM9OE4SCav87evNe0BOBN7kUTcWhDTLk0zXlYev1
KiUGCtacCy0HrWLlKNFHHiUxHVNsPft4eWoCk/iocaJUtZZ6W82tABOexWs4
LwDLyaMGq18OAOhUksKnsPpXYFJf3ph29uybrr5n/qBp0irOGlJUW/65G8ZK
5iq7MmzhNxm+VxSVXZBnnmhrnFqoevMZx6NEtBHtksysCtBTQ7PYMRxOp2zg
RGujajNosvI0y3T4be+omrZHIk+j65eaQeQ2vRn+1CianT5ljAIbVGgtQ8vW
3GmjILWWAlHv+CdJb5DoaG+NBZ3b2vjVL6vGAbaJEkOYXsOVN+0GsP1LLpR0
/9Z2NAmPNwnUI/fApMxeTkyUL94jCiXmGvCt1LFdIhsjes1XL4YjozTekAz3
kSDSliDLMX/U/SDIrLVud8OH/+3dTy84UMF4+hPAAn7tNPYpYD0Lv2yZfhVV
iXzUo/8DKG2P3z9CdZkvMoSRQQ0KmAgBlUrbLiOq/wvd0kGU+tQ9UxGD2knh
IeX7gVtiJyy1JvhdxXK9UPjHmlApmwAHR6YOfC7iwx8JS1m4LP5SeQa/f7bg
a2s1lGNvTuX5Hc49umxfksjovsEhigKCNgwazh3WlsxA/+v22jDTxgNswDdn
wnLXL8LqI+yzYQ1TrX/YVRPFh+v84exdCMODzLOJVcgGVKKTVuaUQhj8nuOA
bbIsiF8vgY0yxlt7HSjcjLe5ibvXWNPwdpHENkVUNxIwSgSX68xrX7TcLJAt
7fiVXUAE4yFcrxdoxwtjwwmru7OogIyJJ1rxCK8BUkAUzWTtzAEhVHCvBF9T
O3XcE6UMeUTxKBWlgIKWscNIF912AJ11q0/j7gXVUE3zUZUzDvDeaHEe1+Kr
yrou8khAnKnwRZemszNaUyiKYYGq5/N3Qsj1MNTuhQJ63b0r+Ic2TMDyB7kQ
opn7whia34PfNWpC2BwPBb8NGG+ahRv5Ch5ZxyKb02I2qGHWigsYLwdrP+QL
PX8w8bCteFoanEUWTkhTZ02nGuAjwVuTJnzVF5EZQo2amw7ZEuoYu0WXYGcf
CLF0mkW5tWmdMomoRw7Vm23JHk/iCs+UPE0jcvzmWD2RQTTU4kAW2FX/ZEF1
4YxD41IgrIpNlg+O7052wxKrCHxyxdxQUq7hA7vv56qG7ZqLPT7+FEF6CmIL
V9rY1zwDMKC1zVjo8U/OiLAL2yrwVTzKhhg7BBESrVH3eA2oDEsHeGBgmy1L
Q463oPAfcp2W0D/tgIXmDv6Xtmw+SL1jUOgE+i7wsEid9TDdGR7UrGGECBal
EhqQpwvHOxRIx2OEmXl+mH1/Tky+AtewZMm7dfSKM2QCXkIDszBY0L6uGAdK
BJQ0sR8GFTrkEucYwjDtsZBVVkSZElkGn0LNvwL2ooVkjvqQTxa1h8K9s8Ij
ganBRTE5mEh5gcRqsnC84ERdHpgT/Yh27C7Q9GQjiOpLq1VFcRGNhxNdD2/Z
fxTFmKxFdLH+Hkg+ZFC1HO+IAeI7Y9dPlCVIFtZ/CcNgW53q1Y8YT4aCFYbu
ITkZSNn6y9gP8NP7VLcoFUQAyJjzU8GdLQ5YZvsdMa+1maZctUGpax4qqM7Q
MA7ST1fqzazm8kdtACcB+civhrMb5poYCKDLiSBFZpUBTU2+LtkKy5yrYGEE
ek6pSHkei/DO4fXjalI+tAMDDA0hb4R3bVrZ6HenpIKc5leDYx4/kHhrlV2s
b7txV2GQcTMc66RCYvp03sxZ27n3lBX6htvj3tyVr/omui7iTys1E3hBrs9C
YNseDHIWDi4Wl8cp657Z5di0wRv/ZyqicKicjr5boUE+DV65NaYkwZK0vEnf
VeVg16NXJPtXJAYC2Hlrf3eXzroD03v7u7f5jsQVU2j8h3ytxCQQ8hN2yVdT
63TFEgdsd0TlfHofuvEIH9Pzaj+xM1vjJ16BxK6IboaOruWJA7bI+4jJWl2R
e9twJIrHy2srIREC1WGWuOnAQ6+qZrKpceIJtI0XBr/gG6XClAEf/yG1xyEV
+f6GE6vW+ZJd3Rf++KCaSCsjqgCn9o0fktDoSdM1UHyY6CJSwZ9KayFWr03s
AT2bflUZmW1kUUamyfRfJUVk1SBe74m0/5e+yAZZoQ7nBzT3wYF4jurzCZv0
lnxHnFNCQLjhZe1X6RjznFKn4N1e2WYGX/s5sRxehmb+hseO+gCOpMeARKqK
DurCV3GKj1keG5js7PMtX+a2f9pjL1ePvHpj2obO1CVJEIZ6OVbqLGT+NTMA
W26GAWTXRYfrusufSecUsSw3SZDyXFK902+QlbR4CphEmvHh6QzjhX/ph62b
JlUSmv94sNjRspsbqLGqwqeVDcW/4sgPNwqtZy0/xcOVzGeke299zN4kJAWz
ykQKdFE/gwEttoWS2r1Etz74cki0uzFydcGfEoJV7HrfsBLskXQceaDaB+oN
7EHjw4yl5v0lMyCPtmqSMlZNjEJB9AxizN+QbcVQL6YFrUpX50fHeKmW7rro
9AcavDxIi2p1QGIjzTyttCS4zC8T6sdq8LQ6tzZbIDJgpqj0GgUBrLyWX71k
U4JjdTXDkrdzoODjGYjlEHKEad70sWexJrp9Zm31j301tdU3SSetAihUmqYw
lbEeQyKqVvRPzOPqs6FFwmoSn0pxbuRk2/ww5+V9o5zgaarl92n5PW98idYL
WaaAPgz6JDEQcfMxw/xOfP59ECuH5LhyNLcOKopamfd8CW5ikSd6lP6D96G9
jKWubP2t1mePbuWjvwkel9EaE377pGAuMIRNTauGqn8KRJKoZathWwQVrWIt
mLoXYJvJYp4asPL5PB2S5O4n9D1rbklU687mwZaIN5VSvN5vqJdcW9HnsqC/
7p1kK9mTIrUn6GlSFMDW5ENxc2UArzr9B1qH/lqIRSIJAX7z0GQIq06qMAXQ
zhbSuCmI92eeGWgcOc/0n8gC3XcD+3VpSmsJrV5LbNLTVhggNCIYTNNVCQR/
sV0IMgyv8EJNKL8BPUg0642OE2/aSdL8PormOM/KMAzfgmLv7R9djpYCw0aC
dWulB0AyI1Is86i0W50ab2thjVXLBNVNYkruXepApL4cQd+8u2zLDPmt54zQ
NBltYLDQzWKdJXKUAEmGW79rEJplfujjSrvL4wWNP6/Q8ECBvjzCnCeOlotg
QIHEiEx+vcrmcHREyyRzN+U3eWCK22uSK263Wpc7V7HRG8nRi1QmCe0t+IJn
VWirRXiNhObIVJ9a4At43fAI2tMiMnkc78Sx+XYnUvwF1HyAp/FApbmeuCQ3
2031bnc7QavVsanj63T9xfX3VRZsxonet0WmK8vixaT5PYekhLhH3o2OCx1p
cM9nT9XGLyWVm1wD3klogUvkn6yN3i9RGvwTYwCj9ErJhkvzhcriYXmocUIB
5qm+p+iBJxzsWxSa/+C73FxaTcskJw9JwNF0CmaenDSk+wfYe72EXNxF/MMz
0k+oTf/y2eNf8mA4o+XuSD3/Xf2nu9L9pmTxevnUrBHl539+KC6hhcQz/39o
G5M9dmyNr71JliDfZrJpJG1X5DUPma8hNtRKP7eZTawNkyBljcRlpcnIErI8
re7+Rnm+EchFlYopxPcB3iR3ovTmrKMnbyu1gW0WLqDyfptmDGmJtuzI0jSc
2/SqCMzoeomrACtNeh86VCwc8fW72XlLyP4vAePJW3CHt9gbNhUd7zGkOq8h
T4iRDi7K1X1mGIxeKRZI/ZHSonOH2Tpt+ZKWjs8fBKFsrbayDNzrbugwn3sJ
KDBU8FcC4xv6vtWijE+Alcu/M38gHSCee97lzygiwcQKl8ZwVSXu88V1EELu
CiYCMVTVwCGe9cjQbwXR33V9QcJXJiDXlR+O7pTjgSEdbT24z+/oIpvAtqui
SUAkVhPrQ/MvCWhGo22Klh8QvBz7qH+l6YMHfIGFe3eg4TXjNzHCWjVAaug0
8kbat8WE/FP4x0IzxdU3YuDF8QK/sKZzfqw0WxVye9EGWxqhnzAQuxa/hhrw
dwyv1WNXBgLOgxHDk0CQmpbYEPrM0Xkp4u6YGG4dRMmM6R11fe6Z2hHO3PDH
xmSOEevzuhPxXVZ5BGQI2KA0MQIoDNFJUuI9tY/AJz36fuiE+FucEFoysY/a
+bIuWfdfp85TZO2K8jBIMeradZVAWdr8Zv/YE8F9aC/jFs/1q7VvM0bgCPvr
o0BnXJBy4528bpV9SyO4gFPPUfDY86cGBG+JPmqPDtXesnlkkd1Z+ojmsEhv
oWgw7+jTgFdkbazU7KXwh0QD0wf7LVUFUcqY0SVwh5FbVBl+fymcUfOvQDuo
f92qfv3y6fM/HvNKJua4HRasK9bIGewpylOrT9UVbSyJ7GGNIQAHKgsxoeBY
iqYFBWqqIxl9WwXVKKIPZwoh3f+yKbKSb6QKTUrAiRCdC/tGxVxeyl2Cv7m7
8fVC9Of1rB8+KEQ6nNK8osidXahYU8ZWqCjheK28rzNgUZZitvvEBSTi+elf
KnIBgZVRm6u7JByAtJ0uWmLgUg4j26xojR0bQWaPbYfPo4bPXmADCssAZd85
eUA9XztumMcH71/7fzhkT2RH0B2Fdql+VsU+nhcYtlzjM5arpHh5Zm81dKgc
Rhi8uPTm6ctVrImbwxVBDe07m1myejRiOChUJ6m5j890RknbxcRFThEqolSp
x7SHUfU+XhcEODjY0KuIfDY+wvQPeJnjY++/DArqvshZSyTIJcOiH3QIB+xj
LtM7sLCWfV9cxPxsiJzxZ76LvyUe/h/XeM6sYwn6E9aI7H9hORWTkMLP5sY+
2liM+CeXtLU+X+LJeAf6+SlIw/3eQrF/acmzGvwyj/ZN8ogaTNM9UfWTzqTU
DRy6G44eOIPOc+C+tIxj8VGUJN3Xg8G/5O/Ct9KlicmBHvRPC2A+psAw7u/3
3pkbDFZyh1MyLGuxNQhlL2kWfN61QOMC/TfJO5llhAx0OPEMAd8U4XvIEb3N
Vy+HCppR1laxqqHSB0Yi5eGiFArXXF7aQsg+HwLEtSHUbZSydS7zSxStDZtx
g/xH6G1CNXbjEbKlFGZMcZVq1rCs81VsUM+GDnpuqm/jf830tqPoFcfThm/j
Z9H2qk3px0js1x23lPR4JmIXNvsi37keK+GnJPqbDL9V7J7hCOba91n7W+vB
56cTerH3IHVgmISSTSAtBdVsgPnEx/rM+KqdmsFLh00+nBzBthX5zEhERbiZ
GF9Dq0y9wu/O2pdlCPVOSDNj9YPO6gvFQvuyq5s7Ziws5EVy4HRy0Hd+Tubi
PKsaHR/uYwXQ2y+Y4GhJJQ7Y6A1e1Tc1g998jgvLUJK95IG34iTi9LTLAsBU
VkXZO+4jRUGgSOWQViAVToELRfqnMpY2KgJZcwYiKuQyt5ryHjhaDeKJ4WFf
jlVA4wXlNPJw4ToOj9MFqhI8rVdOBX1WNZ6ryuNbK/w/TB3Cuf3AqN3aOloA
yOsvTBvpw1IrQedhZZooJUW7eJKahuNPVKkeT4FtohD9mi2qY2u553cWjcA9
4aHaY7Q0Ovlwcmx/3Li3KuEiGmSc0tABXYc1zkK3yY4EQ8yBYIkjPCIuup6K
aH/XV37nOzel931Kn/No7b/7lb5X8v2hJUdDzSGR+9erzuBzYm73xWxRf3Q7
OQOCF+Xei7V7cWHAu4w04WIZ/xVEuq+o7ed8FnZACRYuLuseuBpXihuHs5zb
iDrevTgbVl9b0JC3JEeGacr2UEtk0XAQE1wbsG7s7dXjAEpSCPjzzqz8KQuL
Okxxa2ceq75Xe44okpfqvRN0s7bwmUSqQQvyzXoZE4z2Yw0sSEXqR0wb+S2V
3K1k44hOu7CngGGUubNxe0lK7LugJYRYqeD4NAPWApKK82qN0oRuoLQmsc33
WZuLzBPNZf/PaRXB3/XibLIbjLvBnztN1+3J+hGL+M39aQiSQeOUReCaaQQZ
jbB7+NGMb7B8xO++rHDwy1Tg17rozwq468wh6sNeYtij6FCcUxfYLNB4C3Mq
W0Fk8DdqTG64S4EvsNj+H4cauWJIuawkd6DvdVqhXs0XRhBzi9FblvinZyUs
lx0gH/H6jvARDDkkPZwTB4NnW+syNZgPI2LWCQOR7xQTkiuEWJgsguqNWsQg
09C4fL/qbLHWOHH3VWzYjNG+a0u2kuQbWP7LsSVm6unP762Y5fU6uYPNwgrh
oW8kdXMeGWZP6oP4QogkHex3q40mows0OCDrx01uoDxLnVMB+5d0URqYGaqQ
vU9sWyLWiFO4gNwa9YPVgp1GIH9MxYs6i8Q+AHR0WQIxTuOhuvzGTCC94laP
xHyjUFzrZLIfIAaeH9Os7xFa3BvAENFRSMO0gFkMVqwSDP0nRoM67390qrw3
SfC8gm7gD77hVX2BiwvHsiPOEdgxEfKzWMD2uXbMUQOUlhLGmm8o3GW61bHV
ItS0fJ9prxDnRUsNar8Uq7bdmetLr/DgO9K2R9/kxS1/n/7SbxmFx+9MkqsY
IfhnhMsFH08qksTxYR3h2u4ef+Bj8foc/Z0L7ALHrUsl8NrFVTJqjnQaEDdf
z86m2A190MnONV0no8/Bp5yfdkgAn6j2w26XsBul1PI4hygFCkXQrBy52ZA0
ebvEjHMlr3qAyI10LLnvLBD1UKS2q18uL+sYkfXCNL6lLmmFKGO+KX9bDG9I
utZRxLqPinmQVV6Knc3oEi4pJ8/RaPqPa0s/AfnmbOzLC7oFwqrErD4ESAJ3
moJK+ABOiBz6RpoW0R37NQSWidXYD/BaFykvF9037WutjyNrS1V7teeSwiLH
4K0XHMEwhOxdbVeCbwOfYk26tg9RPHeo3KbBoLHUeyY3eR7okPuq5ySGBMJ4
MieX0b5aQrr2VV2rPr7oKebkUSqVNJhjkaf4wWNHUGGjylNt9R7/HNOmZ1wo
Y3/4t2W7wwfH52qp4uMWWGRStP6T+HJd3qBM7k3DguJzQq5XBphcqDmhPjoT
7P++0QOckkx0Z0p2hjp1ZEwyCTUES02s+cUr+cuQt9oZF2ZBbRJ4OM05f+ot
OUJ2P8fX+k4P3y/26rGe3AaJq6O9jmO2a8F5gelTd2S/iIZra1b5vM5UhyGT
ZJ+n6ov5Qpm7mevoO7ZABezoKMN4jN4wpT2KnnOA+cl82g08DJzupe5dsPGH
8AdvKvVp+LtyV3YeqyhGBICEOW3tQ+UwkvXi/FgswwxhKe/8SjwlXFSPhyAR
VViqBC2jkQ4uBV6JPgV9b4sv269yaa+6HY6QIjs+uWlhOFriUyfDgdH8Auq1
S5UBTyoABPx2q1Of1auJq4VQmmoj3ku1BNPTzh4TyBALLvc/rkVmXDPfKQfF
4tqvSON1tUet8UmjYz7onetJJhfEj/fm6TT1D0FtLeduLltZgFmLVwO7Xu9J
Mny4SWI/1FwNMt1mTk19w/bnEiTtltYLLjmo8HSKS5NgY4Js/OmNPRtvUwXV
GOunw67Wu/2Pdg9fo8aeEQRNQDRSn/EvHA9ekUJWTriEr+8wUDnVEotD0RiF
P/ePzedeHsq38E9SOV6mKCvFBGFR97RNS5DDFqWl7voG55CAIMzgEYTARCNX
ho5vteyuVVNq/2KpGwo9RhHldc0FCUW1Zfz8+ASx8eddt2rqBMsxZ4NSfFgI
9iZ0zp5MlxNaD4KljmQP1xn+G1gpVsyTKEXtJep0KIY/2u1xlJ4djjnsxbHD
XoB9yes+GyWWeVwp7GGnAs93YrQEHrtt0ESAbzgjX6+p4UXddndyfiOcVP14
riXiBSkXnqdQgbrOVEJJ6T6iS6kHoeX+ieuy+fa8BN/g/w7ATJQfVc0Swtsp
v1WyjECC3N0jFosvZv49EBvAfgg17sBhrgcItb+20LNMj7fmrl9MT6wn/2W3
E0Vtji6m03LiUMFb2LGm/G8C3s6/GSuMBp1l8GqSrMy/dXQTqLvpZ5x2Bg4g
cURqPj2mbXASVN3jnMr7Y3Qso5w0BoXrSYm/bBsJJJiNvtFZcP3YPF52/UUj
ZAWSERYHlRBr5oWDHBXcbWvCxz9K8cQT3bsyZdfCbmT96QHI2yW1MBGlznHa
zfR7sDq5pgPFlEe0YTqEP/fFmWJSPG2CgM147stXhU8cpw1KxsAETP7MI5L9
G5UvbJfBoBlvid4QxVeeqF+Rybtg0w5QBlahQ+m6UGFH3N9jufmyGqOoeoaZ
R2CY5jXKo9EfXJxVNBkcO5QNx/qeSv1A5PQthZzlHVOizM6S0S9PEzdoYLGi
1wL+thrQyoMXUPi7LYnn9BdRZGhxGLTXX5ADsOLbgE1yOkujbW9s5YAsebR+
O/LFHEBI2RGomo26txp1U6Q05RFQdDBMriRyDJzZ3j4kD5/nBF/GD/2oIDwp
Af8srb4kqf6zzhqci5eiSb6IsElyCl3HVScJ7cK1FJehroFPTbePzJvXyvQz
R0D2CPHdPT4zoXVEL41jklV9m3cnpiEducsxddAx5SBYqIVEMgHQploNPoPJ
R8nlg4fx6dIdgBmjdjfl/0DDA3aogLvjQzzCCAsgsPNWbW2AcFuiw6ZswL/t
nlPtJBSMuEichEB9qIz1Anzvn0b4UEN1iriI7OG1bB4qkbT0D8Pa9sh+FHWn
NxZciwzv/VjuiwSc2KSYipemzi8nm/l9YONSoDU63Mg+8n+PEqLvo0vVCf/g
nLBTaCxLYYfBXTgOGbRwIM/0lQAvjufIehJT2gDFTbyRtngUMMI/qGhbTSkb
GWZ7Hr7W4nvzAihUrx+ECGI+MdVKmjYgtPju9HxAjDNiQqWPisUHOQOTyFiK
pXgxcRTly81Y2Y/kSpY7y5lsutiI8fVN/n+d25QQiUopuwmaEA4VbR74TVNC
sbeZUl9sBUpzjerGCPDXfPZoSCUKnxrmL3n/AOAGA1VyNLimNx2/cr7SH3ZA
yF2ew/Us8SkV+M6Ne/KwufHGlz6pmG5eTCra22q0kEQxbdJO7KuNsGdoDvMw
VxVlQSUEIsMR7BUa/dc9gX6BTFaJ9DIIhibPgt53u0sn5r7PjEEE/8K1clpK
i7PgCgHrBlt3hHNp5qaHTOtsm4534TyFPYcHyVc4ovn3/kxyL695cBhaDuIz
rsv2zq40Scy3VjRnH0DKEX4vPhWoUgAQKWEmhcymb401Jm8MykrBHEcK05F8
Nm+MvpKGGEleT8Xc9bfXTGNERKiQq23IIGMEAgHew6iHaw4QyKC8mITBmYG3
pkfZR3AtIvtJoqjKgVj3z5819PdUM1rxCfKOUD1OyZoXoI+y/B+Xz2yvD8ug
wwTNsVcSatYv6BD9JQJJR/rJNCm0JZfBEyYElE5xj+r+usfI11cZNV+H4ocI
8XFTFo2Dh/xtdL6XK4jCv2N6aPOGslDOZssb+20YqQ79F0xrOhM7wB2J+YTk
50QUBHM49fq6byUI0Ir2GWAFz6jG2WyjOg3NcfjP1XLThehQQzrUh1K057md
ddX2XgpNlpqdMnsBgdrrKw0hOwORvnPx8amowGItKvB4hTmwP8B5uuv8P3l/
s3QUsqtCipwEAV4DUj72Waj/vBrnVI1Ikb6etGiPQKmekNGpU79QuHFBK+FD
rSvGuDlCrlP4gz7UWqhru2GatZiePAaaTPRuhwmMiJ6yJMcIeXyPfaf8y27G
dygQea4EtDVG+8D79xCDLS/UwaRQJXips+WhT7VUUUC86czeVJ5Tb7gbpiEp
vXp4oyM/0E7B1qTZiNa5PXlKysk+ub4ifzXAf8r7RVY8ertlPi7UEC4N9kYi
Lu8VPAiRJoTafamgT7vugJ9hNYC5VU4wxDCVoOUpxL8BF63Crh+BBpNQ2D8y
wUMWKzXRyVW9iZw4hLMbXJTthJXMp7rMbO0K5jWmzZn6aJp5dSicG3CWouZZ
BPsJXIY2EtUngsb2w+N164pt9nsGSs5AdAty3ZsXNlYJw7jTdA7UcWYNyWUd
FNASWbmszrGhYQdWNG+KetOk9syWsvP+OBiEueXTD1gza/vKz1mFFWk+wz0Z
30idom6FLLGNKYQp74tec4PVY8T3lcHDYpzSYBGXQV1mqmXDvd538hWRDLN1
K1+0tJVQGXYWs/9DsbaSJpj6Rk5ylcsnuwZ/a+f97ylAlTucHo3tVIBhgdWi
PZjAL12XCQmUq4hy/7g4yenwdS6aXvVGcz1OsI64xd6rjfAGUk5nfdUWP8FP
SviHlNiXKl/WGjJsRjZsetSq4daPOuhh3xw1B+60YRPHQDvlZfdzLQ9lhAj9
yCjDxMabzpTVhv/uIwUtWcD+P7sDPZeqnOi1u+mVwCNk5f0BBh3c+3IkdYlI
pCl1PSguUQ0TAaADaeqfLlv1L9hofk1BMDYSTSyLfpjWGXrMarBS6/97iXXO
HESZcwf5285EJG9zVmPG+msQJfmW+0UkQDGoX8/qWaE/SKpOPkoUMm8CxT4k
k7ng/LlluDDYTvQwIgHLsGZ5hVzzDiqszsw7LgWoYmnqXMewohnFcYF0SCur
/w93FHxFnLsDJkCebIkjeM0121hXt4aC6gL4YxU26L/TAgEwFPWMkGMaU1ut
JdQH9aAY3XOwuH9BeFzE7Mf2OuAfcfXGLBcma4ZrqGKW6x0ayQRjRrE7N5ri
eQthMK46yOEYXdLgXacrwdwS/+MfKS0CJdgKBFTz8MjdYJ8CFYqK7ffthFox
WvTvtXxPCsyr5RNqAt1LzaaX8u+RUQ8Ge25L5uVU7gQICJeoUPk2EZGqbDrv
kce0eAaGbF8m/59j287SVTEwe3qJqjNDixeuK2kqgkM1LK20vSZXogGxwnOd
1g0vtj3n/WUdfPnJa5JFNsfpvfag4fZHs5FZb1+Kbl0nVpxyqzp7K+G+F8s7
pe+KC3D82x6T6imsiXdGsqfnHXPQNMw6mDsC6C7vBMBzu/cGkfMYG75E131L
p2dWHgTfj59oSlbvGmiRTRh0xs4GUNaIVPi67J3V2MuZvDRpxu6CBuJiAMW2
SQqlbqjhSTKqc/+bw04t7Aen8cUZTxTsCHAyY60cVdppGl7Lvi9tQeuqs+VJ
NU8MGiBtnpaYfQZPsQqvjeWkbUm4Wq1bsRhM9CXTt+apEkZ3nCFI7nGZJjOj
mzbbwB/eyDfm2zT8ujjZtqamvxpuaZt5XKBern8qqP1e651KYI1bfOdKCi8l
YfHG0PKiPlXi4QeR6SB155wZvH75X8UbXckItkPKndx6kSM6Hut0TvsblZlV
EHABwx2C6fpKnTw0AdPafbFWmlPZ3alziIqbvNU5x9wEQjiJihM0ct4YF3+0
Ul8fynGRHdLu/nh0JN7UYtDZWj9hPkxuFQ8Mi0GH7vwTeiouDzOB+FME3XRP
Z6iKL7KLlqK86JN2mmPjrbf56fb9zxMV1EKaT/bKLgSdlzBgnHvl7KbjSYKO
ol0iJruMesx/i5Kgi2rnqm1tM/KP9jOuf7NVVI0bZqGNawoB9okWQsD8dedO
+kv+kuhANKIVkGT/XdxgxOtO03IJw8FGLMCwesXq5+rklkpl+FnTlbArO3Os
CwCJh+USuuV5M48eQuIFZAr6hgAToB16K4+0cydEdzMNPjEixQrk1BHMHJEV
SBsl4gKNVTdJh6Kk3gdOHc+5xiqlOqnRAFZ5GG3ERRhE9Z4hzkumTDXgQ4TG
D6qqi/W1Clgt7d6ocFo+wkc7mmmJmxwkSk9RKuIZec3tLJ/w3bFoiDhkaBZc
tqERT8R8hgm+BKqZN5SsCfGFFiNPQ/1cakZXcj3VZF6wKbs9BMCq0WcIQpCn
u8EYxRfi2p86cIiivrE4wsroChfYL6SW6BxPxWVMuZvw9M55xOKHNpZ8DcJi
w4o2uqaD7XBdKFnOII/azErpf0cFrYlRDNg3Q1xclitPLPz4FvTebfQSofrs
LTO5uiRe4Zq21OG2LRcpMJobIcFDRWTWLvGjEugYU4PQEm/mDN5olE9K8lEC
zW1jbglRcCq693MFFa7I8Sld7Xis3SS4pbrx7jDbVB8QvZLD/giiGCGsED0T
UNvRa6U4g6QBhbSE9Kwmh1cwf+/lnU8GClAx6hvobL+wd510n0RZMTS2Z8Wx
Tko/ZisONXtojtgJlWn9NksP7rzvvN1nKFj0N7bHUutaSYLu+KUCTbTJiI7H
wI7Q4P28/ISUFHBw6uE9WXN0xe3QU+Ek1IDi6pl4MyVAB0xws7O86Siadw/t
7XITzfbL/rh+T541gv4htxk38SsW6gLKerNPE81Bu59ETNcOL00SRRNYfoAm
EIz1NtWhvxExqhLoNdkRfkw6fa+c2ewk3yZKGoziRh+XRPOpGcf76vGp/zTa
ltbPPF2Ux6ST6w5rrYeV2LdUJGaCrm8Ml3/mzVYFFwDSnnTKVm4WHpDES6NQ
PnjKVvEBorOtfrCItVjYIpSXmCfM/Xw3CmnTBcU7KvP9Xt+DCrOhslCt3Apl
FaEL47A4T22RG/ZKtB7cNf/ghnvdLe3zK2yo7eLdEId8vlsAhNi225yZ0epZ
QcBm4el5zZOrsVV+e4t98KCgRyZnOvnkDlqZTPOYFBwS5XgHmFIinhJuKKam
lbh7Q/uINda4SB5Rw6V7qDf+hHnsWUsz7EXrkwIMcsE3qXVj3hU1q+g0OkHv
m02/87nmvlzlRwKCBNPkUH0z7jG552L5ov8xZY4wg0FHZe/0EHT4ax1FLCh6
J6iA5J2flNT4hlSstz7ss8+Vtoe8YPhh6o0T3k/kZVmQvQiacmdxf3KoL23L
644F+h2gUo3fwN5oT+dUq8h6wzUKKr0aifvhHg3i8HbXNQ/fU4jMd6xePZI8
eUqUg3wHHEuEAfSEMeRnMoOn1lKxctiZOFTcNlGvJYdZ0d5UvGSB6s2aaqk2
2TEftegjEd1ddbW0uEUl4xDhIZHHHs+yElG3CjWGnA0GGxZYWjiQXXcge+MZ
H+66ITy6hWtsqPNrvjy/NV+hGOGpicGprc+cOsoMHCeQASV2dgaiJvj0P/4k
g5GkIq+vi24tuLZIEVDv3Xolf6MwzRwp8I1mNfZv8wM3Fv56oadwTe0QyiPO
g4YQU6KwWaumWP3M2OTr1g2UH08XgG03t2ZuffvALuvqX9f+wcspqRGE0SR1
uvJsxAZXkwAjjuFvAYM6WSdWeQNkBtoo3Zmi2aMKO6hjzavbCOIxIjKo5igl
bAsx0tWc8vSP/rmq33jPPUXizbM6Fnye5AdroPZtTJzakXPQfaT5REKMSk6A
Fht002rJyrYzuWVjlvC2UjTQdWXe5WfhdwgmmKCiUewwyfojCcaloRrjyjxq
G6m15S0p8WtpLB7hPN5ATzagXQG0D0Tq+M4crbf7waZZjGwga+xoOyCS4u0l
pdEy6pWGLAbSikagqcuDEvirzlcFGrFQBv8GTKPCuPc9ooUecsKKi3b2ywKC
wKpYVjGuXQENC/vcR0gOFLZDKgJkqXfkU80sdSmKBXtoh0fRcwuFEA6PS6G+
J8dIww6CFJOe2+SGi6muDDlC84ULjx/WptsUGOnpWtM1++QwO2eo4kg5Ye/H
qIw6HssR1N+oktbOOUm+NDjbMvcX8Nb9ALZQbGIHUdp6xxbM4pFRdQlFVHCI
Dzq0SSUzDsIPp0aVMdELk/Wft+msNJqkHWa/MYGiX/KBxOF0vqTKCpl7oV8k
8D0XOV1MySTlXGAvUHhefURCbiTOtDZ1NDMEEDAo3pTPU0CfkxTi394C3x1E
zluPXqZzyNGYum27ZPe7Mq8K5io3J+OqwR6GLZstp5aXGJi6Qolhm4VaVKcY
CWHETI6tHwOFXXIPyeTP/EvT1HRs5itW3ObiFfwzqA+84H2KXxQy5MkRs6eQ
UmsWSjJGw6/yCw+gW+vDZvdvQbo3p4Y95aasrLFyyBKTX2mXiaKhy0oTgkxN
t/spgNHN6wXi6j3xzSROdk+OBEWAz/So+RjGNFhCciweGrZ3SOmDagA/oWvw
oXBIU3OyWYNw9qvN8PEagjPpTNhskBmTm2nE3hxKd7EDFI0TptAaBvgeDRGZ
wZLk08pXl8GByNIp1AiefZ6yXUs9R5UKdC+Gt3lMLGv8QahJsaYMhpzp0JSk
VbymWhLFc8tb9QFu35wPHeCJ6WrjPIg2BNfKZ7XnnU50/OUDwpjRJ43NYB3K
tsa42LS/4XgTKUw1Z61UqeHFYdC7ZLI6teNmaVptf3pzEVpACHty8qeDrqry
RzS5CZkqVTe2jIkwgy0R5lFyAnRws2He3RlwhAHMss31tgWcvPRAslpLKJnZ
8VfRMJdKBRknVh//jDPNZmR3So3nIFZ8VDhA7/S1z08FRPFPSmygibkjTu73
2+BqTRmGhT+gNWOlRSsMThYMCkSW2YTf+Ymed5bU2JunnunIBEcM1R6i7dSo
vIYftbCi4t5Jj54EChYawA90csUItjD469xyM5dbj21Z7m37tJQsY/gYM/yF
MaxtgYW5clbJ18P3NTnHkHo2sjVO9BtlMtGvjWZpVRa4Zy9ahiyGdAfubukL
CWyFUhzUarImByJSFf+frjyx+xNjbcxLq1wC+rjyZIEqsXNBaJ0FmXk6ARqs
zgTPA93zqOljKdMgfVPDL/RWiyo8rEoGa8WN7q8lza2QPSq7xJngMlHClAPS
suCrNI8NiZDjeMZf/9xJJWdtHtqR/e5jenTSwf1MCyVPQ3ibogau86yg9Bmf
EG3Gxh+tZkYrY1yfiFSKpDn61+06cM+bdT4ZV+1ia7MxkklH1bQexLEDFpkl
RaVQA4gxicq50XUQU2HYvmbPg6i/afmm/P/keUX+VQm5Ym3xhUqFDOknTox5
w3mce3NVzWVOjMQ7YJx3H2noNjgKdx3EHhlmub0D0EfyB9BXBnx8mcb+dbKY
5BoaEGK2QY3bUxQb7KduWZEirIViaZ17dgZJ+anA3ux1ftJy2iGAl5xkt+Wr
/Mm7/jp17j7YLyVG3PkuHpPnT6qonSB51VE+fXX61Nk6bNnqfsnY9QOcld4x
EFQ9nzy8sK0cf4W+ycOaDFQnkXSUYFMZw89DTdbOl/23kveGqDQmmV3j01RE
REyfVn8ANhjWBps9cNaDGCdgxvVo+uA95XCjG/n6CezGF2TvA6ybXLjtv9qA
5rKTxFnhxHWh0JPM7onBhARk849qiNMQ5hf1aO9RFUXjqflEnIxMYhAtINpp
4hl5w2aGVlycsDs/QvZ/+ELKDaKGJMn9wbKrLNkv0ziitDFlv4bB9p3sBaMk
SOMJBC2bx7tQN6j9vXA405jAfCaZb8jOSG0N1hdsjT/DdDqztYCw7MQN0y4q
xk+JaOVgo7a5B4NucSYjf29Y11vTKrR76bBZPwmBCbKbYgO6xxX2FCj49yRO
03tu7fwWGhsyweizMy1bzydi9nd+aC3j76CZ537yzViX5jqJ4Qbbdo/TNYcl
dms04BCPcrUwNRRgUE3drj9ychMQUTh6a5iZSBY+UOebVLMeDQ9+v42d9tmK
+8+hbF9nxQ41mNZLXwKU4/jbnbwQV6QiTcJCcJ/2zk99t4Oy0JNHGEySqapt
DkXtbZhg0qC1xp/4vJ0KKql1lhdN3bPSCmLbYnpS0wqXXIT/OxyBx5UoLpwZ
iMltB8Y9k4nDHubE7iBt6KpcYbqz5oiLoHyMrEENgR2TdjA68aVE2KDqGu+t
O4uzEmRP49NEhjuOU0pgjnRl08qeR4tr/n4m7tkdtj1P91Abvt3Mcv3zLOHF
NCaqGIw+IYfQRL0WSDjkOCSUmKzCE3zWZe8UNb+i2e2tdu4wLPD8d/WRQ7ov
Y6azxr3rNEe17pJ4H8j1jxyTMN3pREgB3WvHD5xxQBk2wDlXrWtydxT3yHBl
39ZCS7UKDY5xl6ZScLYXZ/iAQSwk2VMVc7Kwje+hQbkYG3g/WwxVl3IdEwr9
hk8ZeXH4UI9SNWpvRbO3ASPV7OJIojl3bUNHo7MzTSXOYLzFgBqPc9xbDtTF
gMHkTBczyscQ0iXwvMCXtsy4H9QzNcxA7jACnGViBlwwuDv38oZOhyuXlG14
L/V39lIfOrLNR0wJ0ppTLwn0kgOkAf74JRBj6RmGntKpPucuj81oBhUe5Rrc
gL0PZHe2ZxLIza3y+HpGoYT+UxcUYRLhLdmSpGHFp65QxDkmkETPDgekwHr8
ELdwN37HnSUNBMB0gUFpYSyqM8oWWAVFMGirb8i/c64hGWpFKBrX2jo+Wk7y
OG1eW+HkbdYyx7Ujh1mhLNdiy2tRLhZPnHqXJAjWQWNvT/ww9gj/t5IwqPpc
WAl4tO4gKZy5iEZ54k5OdU5Xfnm+2IfL4rLmQIrWI8+u33fS8kezhZh1hdh2
WnQdszlhcL20k26ToW1GfndtIlqH8rCJnKqi5p9+aRPy8nB5ADlSXby1yf4T
lSzaE9TIE2ywVqSGny8PNEbVjwZHXI6dIWCXrVlHNpfP93wLY/HVTNsHehRr
C6E8xA6pF+FBeEKnAvSHIPsbXQkjpO0GzJCgujHBLUZW7dFdpFol64Na+/Jf
d+9xTAaBOKfNhLO4HO9KSdGwwhMu+NLtd4A67HNEe+b1SkkFmCpQz5Oooc3h
M4rtVVzisEFeAoyrlnqAbkFbIqCocgjapkryC/8wUk1GEfY05wsk55GdRoqg
5GQWXjEyi3egw89x/MFyHf511sS9hNl6tCwUdF/Ubf1xqQOXHDZwGIJx0Enk
59FfNprmVg6zdDZk8NviK211aj9cH9SPQXvqU/xV/jBQrqjW9nCsHVqldLwU
IX5UVf+AMxhAJUx4GITT2W4yehRAMtXQBUqfvBbzEaObRRXhSecRiYVHDgEZ
uoK9N50hNJVTmkwix6MDJDrlTgAJg5ZHE/sAqObEEiKF1kP5KBHyyzQxvLe+
eaqC6outtTdNQ1/yT5Ont322qCm53PrIojyGw/eZvMDgspNBh5ohqr/GY6rX
4iy76IQQ2/oSrS9RVtbzii7vTnXVyIx0ZFtKHYMRY62+3QZq14vsGd6CoiRm
CcBKlmuWM2nKzQZpfG0RcfZvoaCJPF/BW97rNoAEiz5cGsf8Giu46kHOC5KT
h9U0rCnC153Pjro7ZbsGbE789tJogIQ3CZFUnRQ0HjtR3etqW6OmZFwyCLEw
PNuo53ztRMaY88Dd2xUXoYOYWgIO0WY21EC9dVYYNJmLj0wKJ5NhkciiM8KW
kDU3gTpwYDuGzWT/Pcp3Q/XnG9lP9ZwOEEG9ou6wdllGfbWcT6trZB9gcVMJ
/4J44xrL4rVAo9os/OaB/bbIwWrSkISJMCAirTn85cDY3ZdrQIvWrXOVj1YJ
E7e8Z/pGpDKsXbjENBIrE2syPdFhhhm7PCHUlBSbJ+evnrK+o/iT7KIKafzu
d3gLds8rg8D024T7LK7JA9xYvqOPg4N2LL7leUbMOHXl7Q/KaBPeXFDFpVPw
m9Af4/3B6bxxc/dO4A0xDUkZ79SIoO1B/3joPB7gWcTQTvmdsAeMbmq27S6i
AJgOdCIjZk/dRUxVcKc3cUDQ1/IxSLyvOl5SSRTvpUL0B/rEYhRUdJi/dDOv
2KCakj7HcUgjuE+PtI59FhvhH+HMJuOFoyP9BT9iV9bWy2b46ca6bu2dEi48
E/kKLSqpV7lglBCqJkSPQ3sSs9VDgMjl8OUVtZ4FDaRQyXzX07hloMLUJOzz
zM/Dio8CYlVA5NrAYGNGS7AgVZwnWds7ZzbF3d/bxyf4d3vU1di1gA/Qck7g
yPpIMPRlGlIT32XyVnW8xGeRhe95RJoiot4fq7FEeCN3fueivWyba4Scy0VO
LVQdduwYOac5A6YGYawUq/ZBSVarcoY39otYEFeGDrjsm8MfSo1qlY361Gm8
CfG7jHqgGYVgy04tb4/vMB8CW1eFNQVYeyVZ89GYITzdwGyJXD8dUumulFIh
KGJQO2ZrFaeP/kQkyBbfJgcv3diOCHb+gEqfJFMi7VSgZUmVWtx/hEOUzsTx
8N8D39uxOO31zSf6GZVtymEuI9AVMI8KC08GJVtjvjKZDA6JqGWTPWOtfzV3
GsC53UZlsbYWSsbaOivN5SN3CYEb6JkN+Ze5n4einoBRIewQc4l0jk+NiSiT
dqO0O980NZW/g+60oE1X5xBnCXvfT5aN9tm+eDxSWqdvcvoyD45WFNGwouRh
vWMJB7Pj6bRvfh1vmUEd56gf9TNsY3IobfGYrovJcxHy8ZqxkvlVmJRIrGrQ
Xbjz9jqAU9WPlIijMFmDolUxw065JPzIetgvNKWUlfmVfKtgdzbC8GISz5mE
pUeROYk1WJB6mVq5qlqOpxgtOX5Q/JrA15nwdMs9rckAqaJ/oHvAQ0l0oxKB
bxXvXDCPUSS7/1lqQEX+6/NaMGSTfRmWYTf277AKOU84REtlKIs7zyau6tjy
FXRpCQKSEnWIpmRPn8NNgJtuCmF4d4LIU9J+6ekDzc5TCD+/ilfHb98tQlXW
imCfyWz8/P9hymZO6IChqc5ZPS1gRHSldDTLcHtCLk7jpX9l9hbhd0qaNcEl
+rSKQlE9TJik/HQNGoPCW2OTDR9cmkEBgktaBrWpC8RRjqLS6bxOaXVnTSW5
EzvVw7zj9dIhdydNoxSyjl0B9AXCdxYJHMEgNmWoMKLZjB3KJ0TqRnM4t0ir
Ycbn+E8BJrEKGeACQ1QCJc3muGJ28dW66f3MSJNTjEz249sekMN8gyWiy6Uw
7wiqgoncvN7bDxoWOagBTGhlpjepd4xYkjXIouqIctmAzFALh74NuCswoDWZ
XS3QFsnmY+8qszx0bdRpKCbinvQaKPCWEfcfTmzwyzYQYV1Erw69Vvf9bh4m
dKL9BjCesp5EOCwcFjyCQc0EWPDCeAo4XyIafbY/UWp7kLivv1UnBJIFtKvK
YGoaybGuQo62ANPCiJNcnSqR8Q7sVLvUz0jLadYA5HSIsE0ZKKlk10a4ksrh
BubmjoLFJm5MKnvaWb4gftbDH6yqkVUEYW4acOXvxN95sDx8L7ssXg95y3fd
DcQXVX5uW1a5W1VRlOGsxuamSxExXeRa9jZgMHGGTv1Z8f/6CCBr3qMvM8XG
7ULwIliE7HC8Amtpz5A6woZbPEvekp5i3CFevp4lTjV7jFvzBlFcxx9g6OyO
3W9TXY8+Q+HbAw2NbHfQEfhYoRkVQXMaUDouMQR6MMdA0P9K6/7Kuuzf6T7V
rU216sbDjMN1rucjSIwwn6kfnE1uJHAKmtlESEP6jlOvVkk5YprGnkI9ouuX
Mk9JAJ+8WneRfNPGLM8SlgYaJVP1cif6+cB6SnROYF5aFXp1pbzoHHwUqVGS
PCfb3r6l5D38M9IGAJD2TDhsIWUf0nXBvYr7UCPtH/XuQBK3UWSy5orELeJL
jDc735r/7RvuGGJ4zln0fbPjnnI0ntvD+9K8gzjj2lrIUbCc9xA2gUDkkXUy
yv/T3E1MwYav4fhiYpQemdEYdJx+AJYe1X7KdWOFpAQt5+yspAtoPOKzB/Ui
CE24jvBuuVwsTnaLU0HgHCQCYduxWtH0m59EViVc/vpzR77I4CHTS3V6E+Gr
c9V8q0InUafUVsLSAwGuqhqWWkVYN4kxuhliyumIklVJ2Y1lgLLAKonBU/Xx
jtGf1fTsJVWPVjlKmja2KoC1wjrr3sOD0A5TTivtlGuxiX/niUyNS3S+ECQp
a0M2Sj6XBF4K3IQaPvgg7XWOh4LtgzXfgE9IOOpoq7f6d976pcE6QT4BTmJf
vCCUu37jtYeZw/T+aQK0nZdUJpicsjJ3a0potAD5YaYsbytB+xtLqhRt+mf6
8hUg3MA0CBJJIVlH46P/Axw8m2CDEUQx/8PXbBGkFxF8ddngQFY/axcn5RnW
BcJm7asvFDXz415Eg3SzB0Z7ehYUe3n8hNlFIafANUaoSGRYzMHJHbfT7A2Y
6Mu4vdGHDT+WoNffo7qceQXj5M+mf7nzHB5yPTes2UI3rDhenyGYwpSDM41E
0OBi2fZUFT/NEKAKUHXJ33LbNtiAOeTABlaPfcnwjHZDXxD9ME+VIWOQhRIh
lAu6aUshsbKryNoxUFeLXPupy+s6wMSayuvfXXZtqP2s0iwfBBp4OQkAG4hP
/aTFS/vGJgg2RMJ6KHLJ3fr10ENQEncDugZxUtUfFXbMpi8cPtba3fBaZq+X
oKaJcutIewfvI8Q44/X1UCPRsNYJlGTmb4dogfyTVOcI1EcARb4vU9F1WakW
kxq8Z7sl4tRWE3rjubA5D4oojrLX+IKRKDPuRvkJRZuUGnolwzqqlYaXaAY/
CbyQqMgcIJsf/AS0WDx+0qFqWddgQ/yabWAlW9UR1yV8aU7xx2IkRQPa9g63
8s5MQVi5wv055LE2cPVWLteXXl5nbIRowy3ZRuq3dQUeyRV1fLId3vBhawaF
RyNO7u6sc6+qdRCNysIfYDs1TrQOPd4lckPTYLQeSRDninEpJPISCDtW3ijs
sWdk2G9T0O5+N8xJKnp0PCC80iAtXiAQBwtAf0pgv81dUVzTwSFYyuzTSg1W
WnHfyNmmV42BTZpInpucNZj6BvcnlKGif6G2bzjzHVOEHlla4rWB3YiM479p
Sro1l9a/nBw/2z4+xOOvIjpIE2VuI7NGsCFun0eDYx+Iv5aKMeZiXageifdm
nAhH3egZzGvA1XmBLx0B4TxkEAHVea7SdMNeb4OSGyMJbkAc4aj07/jzPT+L
L1ecq86NtiEYfyX0WjINZ4OsipZgdBuwmJWBlnF0iWVCIRFyye+tdO48+a+w
uslP34TVF6RvuujhPuaubsQjABzOXt+Px4AlnNhB8PtebH/XMCUG5Ks3h9KM
Fu+xf0LVf6wYugPXIzAdJJVEtTpPpWieweDmRDFTqWVbrU3d+jWcY3wUmvJa
CmvOXqtrfBzn/v11qi/dHJIhmmSkvotUhLfHpPhRWDJHAlCQg35fx23KpsJj
XyWQoF86s2GnFf9N13bI2wfJsBLziqnXLoO2qIXHhlxYoIFJTUf71mmnQRJ4
1OkbH8UC5TTRdDIjxYz3cYS4UrpAwC0DRojy3A1cKQADxeD9iqhoRIF6+VIB
OP7HWKhBkZtb0fJaYxA8jhEoz4F7G18SdC6ExqItjuf8qiiN7yyyiaIiSQEt
BlptvosjQ+pMVCGHP2Kx+cY2fNp6HLeOKTLHEwkDbd9gpNG7gJVolq5VKaDJ
zXAbs5DbGGZofQZY4PdIl7C3mo3NBMGmLpx6Mv/BRRAhgbrfP6gDsy/p3JoS
bzeT3ks2igEBYTpSpoUHO4zCSTh6lLiNc9Dbfa0k9vwL/bAnv3Zagtyd0qxU
u3+uEEvB4HnvMsGfKhppliRRobfkD9GoaXNz4IfaK0lgerFGSl3rUPT5GU4u
dO3c3wURK/tAVPKqT+GCRKm0kE0HjIl3nzTp45ekr5WZd0egtNQVDxGf7CIH
sO3Y+nGcGsCVRVqBAXNdDk5YKMcj2271+iDgJx0gt2gpJTbiIk5PDjm3LyMI
Q8bkS3v14m7uPFb+p+smxHWcR1tk6xbeznJaDiUYLdhrkUBpGW4GqS8u2z1M
5MUPdgx9uO0JJ/Gy/Nbg48JDvuvRv+3hyaUu4CdEA1S6Y8qOuUW1fo0AO0HN
Pf+94M9T6bzZXQjxZ8iQue5gyR9RVgD9OJw3hVDxng/jmZlxWzXy/HF2j7+5
Z2xz05v+UPOG/T4cwa/LpIWHAq7TPLkUNZPeCLsJj7O+VBD9s7fjuMsYWDjZ
pci+ybDO1ZN2pxAmpDW+os6OBUBlXUQ3MBjlFvJt5cigLVScEROt3mwjmnjM
cbKVmY6rAKyVkv85wrzHCskStHAr9uLRsRVzANe67Uxbt63RZRgKlY0uDa5a
0Acizos2bGxI4poK6B1IoCgmaK2cyI5kPfabe55aj3aw66gr0BMpQCO1l/eT
kSbGGqzAyY0J1gl9b+SLCwl8ZuEM+MddfQYNoSe9qmbNxTTSv31eB+yawj38
g/PRLwIlZFcHf9OmBRIRMl3PUKJGwW/2GT+sJQH2GGMFqE4nzS1lHxb52kpc
bfl3GrHTtOOe3iGunPjyoCxQzIZZZLWXPlUxYvonx95WMnRoXfqffohKfS/S
FAz7l42fr6xq1fArPiSwAjK+yPIIFZ/so39C2cJ21DceigZRhpaPMrwaEzRy
VRqCoX5kPh0hRWDqAv81xVSigGsdJRzlA1RXpim9QzrouvGPbFBO0RN5VTOZ
DvX3mzX6XNyF25UqS+/j1ut3OrLSFiNnsIDE2KToG9Wq97ytrS8170jQpAZb
3n/5Aw0Lii1w+eNeIa6yjgZ4aD2Lkf4JeZTmTgvDO6DbKRTlvhAE1w9ObupG
397tRyUYWAxa9ne6WKVNrQUPexoAu4D3jluZwjeSyq3Re7PdHs/Ie81vck+1
JjWKGOx20KJoFcwZaVpoROBrwEiZTg/PdkBj1/u8u+Ergtfc80hrPds+aQ+L
wlPHt2ffLGQG2jDPPLzE3fwXPCC9XYWsg5o4Pbw77HNuVLhnqKUSFnvHeCZV
GeNQb7InxJ+T974mad4YoOKKloxZJNTz2vmTYb8imA552puy2fj8cbSrLxuD
RhHsvcyOsBHcHD94aTU5d1pX6a2uPfEUoq8lU1pJBai7JS2reNpIPskGBK/l
Dx5LccXoHbflF+GRhPHKe5Eph9ql35bE2xzzfukMyQfg+2/GTbCDLpcnCJCl
Ky6YDlc/xBpPoScuf4EVojzPsp1KQIgg8NMzmfC7jZKjWvvHvwBw1JyhCjPg
lbriZfeIXbWrbVH+STgEKhfkmoN3bvSm5GA+1+tiwsj0DpPycxHbZUxLZlYh
b5awL5/TkycmnirFtqXVbX9gGSzeclHa9bX0noM6MPez3l1TRuT8NhwrNZbf
kPXxqv3gh/ZNiKuoZz4Odesig8kSDXCQOEfOQZaFHzeGbvvFzxUfr0ANYvjH
795rYjsh5U8RbwwvuHBgXfixDEbZuACAyzwDo/URPLOnu04Nw0/QW0aN0wWx
mRMJ++eD5oNCCP+INt0aUg4BNL3I/9vE99Cvhcn7c33o25s1h2NMErFmhUSt
Ma02rrzTIQR0AAlOxJLNKIX3elfPwGl1dMEefQPYm0HL3Q6M/MMMz4104ZUo
dsj1MDY3tGsNn7uxSbeoGk7z84+sRbSY9bo4IU6BJcOEHh6y8HlAanh/9c7/
dhB3ImH1Nb0deTyiT/qGfUENkiRiHGSzjHwvSr2aO863sEsVOw166W9V6BkA
N7fNiojFnXpy7T3w0o3VX8hp9kLBUgrZE5mWj9ZUlmxR66UMXm14a6TxGen8
knKYp1sH0K+nsdw3IBOVsqv0O0ke4C9qB93TrUuPxz0S+uxGXPrf/2n9zT8O
J2gcsYbb0+KMULjJIyyhjr6xtHJHwNlImXJz4ndEW7zYfI9j41vziy7olntA
jfZy/yeaumb9y2grR/Bj5SBO8tOJePVUew7RsIKM7HN3l2Sxwl12AAH2PhkB
7vU3XVW42HQcVYY1B+/bwcBsbd5aXegpUoGbRqjtmo7g9Ne9G2vfMqN50ANd
09MJ/UaEo6nMOqkxyXbU8HRmrMqpu8obHE/wyQvxda5/ODLIq62TsMcgTt9a
RtaNJVb6XcpY8tNZwjg54R/JXFU+ByTJY6Tlqufhtz6Tv+fxPUAFgm637Gs8
GIsschsSKnpSjzfmXwa3yv6Pl2TGFq7hLVTrbC/T6SJGkHV98PonUu/Qf2uL
3RWdNfz0XX+DWDqf4EIKghMq8Q0o0C5St50zJw+uCih8HhnjFccPSDCR0OvM
Xl5EGPjXSzwsBVqk8aomiUEDIq99QQ/uLkWbF75vfnp0KqocvzzFPk/LJDTF
lI9BuIm2kV5pyyeQdyVrVQyyzxhxT6rRZmoA6yzi+AoLGH+uCRZTBtjHLHq6
fi1oboEPxkhTSO5XhgvOswTqCbY9LKbaE300GDlBWYzbjyK/O31ZyRVIVT3n
oXWTiUUyxNrecDMtgLb4cEXE4IFVDBZv0YoJnEHhhUUJgmP3K5G8EOKaRfp6
pDlFyseCm9ilCvXTOBR/qjwh+lFRAxtDCi/U5VX5KPr9w8ROKXylh9NFRK8b
Tx5qR+3HR/3OpItgxiHIVTAg6+uyd8QBYmfPSvR4L98gWm4I1xCArAccX4xa
mvTYHySHGvpBV25YLlq8b+dFOjgiOUkmlBE515aUvW0FvpV0178TqIwCDqoj
dy0fvIEbqRe8kbnue5xK+hgoyiO5Dd7etBRbemcn9oyagLK3AsBSsrGnaQoK
wuBrr4fyMXCl3lCqi1lRSG/oAenpKWKrHHmlgUSK9r7YU40m5/3+mGnUnCQz
s4uRyj0AxLkXAnZtMMTrvqQu9OuB5VgNEyu1b93whhOvRvvtPA1V4aWMMpO9
ZV1+LVXKjJYKIZExvSFpnIU9vQl6QRLj3zieOZr35Gha0k2a0+SxI93OK1Pc
T+gsBXsyMyB28cYSyaS97YQg+4uB6v867WkyRDDPPN3Y8nRoFI4gJbDEX26H
Gn9UAfgclC6WAZ/bof7bTQb0UeauWU5mwJjvxf6P8J7mjEb6vMCU7dtlH55Q
IIcn1BXSy5OndeRbhwJ/I754s9kZM02r9+TH63cUyROEMhadaqVR0jcScdYh
X7i2G+r/jwNJsaOjM/KpDnjZGcqKKB7oG4qjzdATSXFT8Z7LwLB7HT2TJwry
aGYn8qPUAEGozalSf+XZhcihVkxi1fBum8SYuJNDBtZT3qOf49RAoXIyjwTz
koJ5W7bY7CPkFOJUlltdvGf6oopUv+FTgywBQz9r4uEcWud3CT120n1mKJsF
Jl8L0x9YLgB6St4uALh+Pek6YaLuFRrbfIekgPcW+Fr1NWHUXt1BlTlm0dry
Lyzw9bbKGQmH4Cb62mh8DdS8Yyd8Pc1P+tL2fsF5WhsKqV99l3Pe+6KvpJ2B
EbsK4IL7YkWEBvQ2rUHlrBsLUAeR1srA/qoz+jtjGF6TO0KiRz+8mj46+XVG
j6fokcsJwEJpgcisCO1noSjGdkwYWZRrbCzQNbJQR+yciPITmebdKqvIbv+C
FxqHp0qr3Of6E/Zsic16pPx9OhcBWUXo/+9BuFZAkmoXdvgpXC9AN/tMJU4L
bmO9tlPn7vRM9NY75WxwMzTe5smEk5zqMzAa+zuPl+5uVguzPYR8G2SmB3Rz
00huP96o+jyqjMJE+JbgaG1Ivx2PbeaQTtDCfLKoeNgGlDKwkdN1mtqlREuQ
BVM2zzpY7pwCtf2nJn99e1+om2Ry+m4CcsuFvgj/lRi2cudJ2rhQ2pTUA1Hp
SRqcfHgW4saV7nBhH32SS69P48EOmMG4Ote4bZWrXCCrXg2mMCCKDiaGBrUH
3k5J7BMU00tfXD468kba598OP2pvX2zy5B6znRWBS4nFOfD51MMJ3tzeF3za
SFUuNnTVuu9zmiJjigPClonHJJ7K0Z/Rl/dH+SN3o3DYoKqPY9fRisDJQCEK
lwLDo0lbFLcTNyb68RkUY6BE7FD2o19lcaqDtV0enie9zc17GUAUzc67pTxB
Wm4ZxDuGSChWzU72DXbLQp5EDaWrdZ5VHscwGTwBt2BaTsfk+H02hpO1LBnk
xb7jZxmh9MU1wgTnR9YgsB2+HQakSnvffrlXZjVb3Fp9cCr5PPU4qFFDf1z0
SvXGnRWTtmBEa3Oi/qluNiZR6oPYIHf28A7ZtEAzaiTm6pXEq3l/ZB2sBIEx
DTiEI23ToXA/FEDSSpF46S1la/XG1Py+blE7uUW5sFmIOG+st9+krT++jioU
Qqx2MjUu/mbl2K4f2w76nbGAKUw06IV9E3qFWA6iYBR1Akwki9vtuTmrh0uS
ffk6QK7J1XpZaPN7awgXHnrB5T6zRtnSQvlnGuDiMum6cT3orNaEklM67zFE
APsPIGJBnrdV+OW0Wi3Ifes5y2jY0XEF2qtXIxMNO1top1AJuizuqKsVmkRa
c5nUA63vCBmXDFT5WkdVAJNMlZsZIIpOnlC68jyH4SNwpgeu4UwBXiu1RE6V
vxIkPuDawJeS/RKKkz6AZ+nZWi8ndmi3apYEcviwNmZYIgvVDtnK5QlTMQYG
MSoOuAMrXupLDOYI/Nl5RsqY/LaMPeeb00KHAIjlKDXywmCSJK5H1lf/ew/b
7plf9Bd2PTB2WAZZWr4MIPQMq0q7Kap+gCXyxA1msHFve59BwujDeFEO4sKi
UTecl6In0cZELnl5mUKhtF92hgcGUyB540uN0xXxIDtg0TYYpsYtwDDqxgcg
0tIidiv2jwnTegR67VuCOdksmh1sj0vvKsJWQ8QMJ/YCUbkRr2h1+pi4sHAQ
srzxIA7+RcosuqoPZUP5mFmgwK46UVlvKg0e+qgynCmw8g36MmnZFqgw5r7I
FTXA3SrilkALCXZi/TvJjTonMIe/+aVcJ+mIqjvXoxKxlWRq2MurX0zep+IJ
0pOKRe5WTlW4VXwfNFDTc7j/K1e9W9KkgokLChzAvggJN/6tlieJky4Zpgzv
0IAn6iU9ZP0eBxDPb4/rOXlD2ZuAfBB+W2oRHgIfwZ3REQUfdJyT4hll5qiw
FaiZDXeKQs3ZW00OBuk54XWWfKF0n170Z1mxIthXpykA+Ixc4Xjm/aPmUHZd
tpPg4hFEI90RSEbZkPTtneqhMHxaSAOqDJMjXoVk5D5tJyZ48pLeTkGZf7mG
cYybidvj6izU2+K9W71MgbRLCjz9orj9Ux290K/7txmLDhgjSJg5+zWnmJ6k
a21gTcCrwzL+lJBecSFCwtsiUhoZCyaVanxb7yfIWRFcGLaB4qHpYSQIPbpl
MLufbxY15fjgoktaz4uXbSRZSPibbn5mfOJNjHphSCaZ3N2BP+ErtwoaHWJj
uiG8slO5ImGRknS8LP7s0hVuc67feQ0LmQb+P/lQg7WmAWb3fyg5p5/WO3HB
E8cgqc1y4SilI4HnlbTQZFtcDXfqv5NxmuYbpkZPgUW7a4vQTlhGPPAznI2q
fgQhT4Ua6p3HdRFR54yY8xO/NsktxHDBgO2Dl+BcFd1s49J33eLaEdRXrL2q
4dAvUI6Ag//vMD5Ixo6hqq0vT0JaySu6zQBcOYS3HDkqKs5UADbypJt6N9IL
InzFs5zK2l3+MnB48VcZgdwGuY8uLLxpANGitfTmrJONtkWZhRjYN4Oq+gCt
V03iouuRIIgZExEAQ81Nl20vN8UklK5KBLfeTDMec4SK+aPpuyU6qf09IfPM
YE8xXBIpBhcnlhtpP8P+EUcZV7xUPpnV03ucNwczNSg91XaF61q1eyyrTQrg
bYbzt8jOVP2EkN7GYZGB8Vfts3Ak6mur9M9OB31B+iCNxX6j2FTmPbvKyKIt
rI5tt039/807yDu7o7Wr4tEPe7YX0i7Y6hzH6/dpDbPhgw8JZUf4Q3bDzWXO
fDs9AlAYnQmQaEAx+BjQXrSFWix+7YXTSEYwnXZUJKT0xRK8lB+IHdlW1D1x
qqWXbgjuNzFye2UIUQguumkfQedP24asXBmQGFVuQynXFTqq9yKfHwTnf4tU
DU8jSOCCavslN/673gJ6zps/W487WHgO6N8Z74FVcuVJFgBr4bVTI1v/npyC
rJqUexJfyCAxai/ri2FqWGptCjyre8zzlivDy+cWNnPGDzIq1/ZnzuJ4m/Rj
V8GbagFQbO0b0tz7b/sfGuY0P0PgNrdDys/UVS1x4Ud7XlfO1Qo8kbdT4Qdx
X6PJF9lSaZ9jiYsMOLqPsSiRKei6ZYIaEP09N81NDXmln4UgHqx7FgeySXP+
4iBPmC9d98OmVRwfjRrWooy+icQR0aSAvPhVGL+KVzPjN0+nDr8x2BLzbOw2
WY+OHzDSIfc815IGoXTtsiaYh4ujl5pWJ1vYWrewuczFf7wLLad1SMwEfhWs
y11+4yC3m9CPKIOe4/pJSRND6fQ0KiP4l3+t+coOxjxkP4aXK9XXv3tFBF5y
J4/njbPdnY6RoKoTjDdOjYuA8nYVCZwd8m2YzibObjekBfesc0jjcn8imfnN
SV2eOn4cV5slyMjZWVYKrfDS1YGeoalO7c7LhCDUFE/RJ6wFs8FaHjtyOgCZ
z3ROPLUM6Y5/b+L8oyZz8Q5PPzjdKlu/whuN8xZ/LI6JTMmP643tQXXKrK3X
9WL9NumhAWgBerkbJCQlS9WpIhUMHqLcUQT90zDGEkVYoYADjhUQVmefXJ1P
omef1XHgOjq2+rg3VkTK0PbGmNXJ2Sm6fzAJ+ipRQB4HtW1P55kZzCAC3T/O
b9l7SLdzMmm4wgEKvONQXU7HR2H4/uFY1zP2UIga8TMLJF9fjhIy7i1eZei1
WVsNHkikvCRPpPhx83WjcRc57Rhlk0H/jOyb2oIA2STOrYHEZJJpUiebONzp
hwCEV1A+SFjihfaNzbsTZiBKez4Kka+sRuQf/2gmMrfkw2Hljf5I4lu2X8Mr
q1G3IZYL/1lBVV8FLoaeNkKZMP6CyMUpWxgc2WxAfpvjAg7XKl4I8UYRpqdF
fFf2EymmkhRWZsq0X216tyq9HNknbzt7I5Wm1Cpqp9r9OjBUZK4fD8AsrgM5
E7POjBfDeCQYQqzXwrTAlBpKlKKp0i9QAQFksRToDIvmeVDvNU3/f6Ecr/p5
PqZK32DvnJ07Fhk4PE21ORlXu6K2GmjDMUMgDOudO330EI9Gu2+LOqq0RG+h
P6JiyGT9yx/7hMruU6lKwByUhkPD+lZirIthJ4mSLFhKJEvP/s9IYWn1rhW3
x3yylzDPATzccABeN7GQ0xLtcsJDqAd1feju2VQR6aWmbCVs+7BE9egkxqka
HTub4iRAP8NV+r2OY+qnJwyLroHm26hyyMEpeCOg2TdaM3nkDE5C9kBOb341
UU5trf8CwuUhJbbdirtVlwf0PAxjjm4Cpw0AoRhLoWZuSy58u8F9XcONFJqP
b928yZLegj4hkFZ80RD3KvUo5sAOPNnJy8KtIPdn2vopojomNIovJJC2jT2/
ll088F5clBWoo3k+CMAWqZN6UyTq4z1P7YsBG5KgQRzSETPE15rkkH4N9eMy
5dP/yuqzOjfVb0NiHUo/faDyizxYEnaS6RGLXIVSknG8CXMCkRGwCKCzWLig
PGMoCrp3QaLfxXwtxVlPwCR8Fwyf3tYng0aymllJ8eXNrnGzcWe8O/P21eoK
8K/fEl/haaVBkVlcs7vXqv3GFXqkYYlU5KiXy5yUPh3Z+mdh5rvfP9UdwtdR
YQlRIk/cS+6I4g1dpTOyXNFO6IhYuAba1XzmeBNcJLxkhOquS5FeLMHifmSu
sprx8VeyyA4p1tgKeU0FUVExkx2CHDB2whiJ+pjleb22VVI9MKn5McJfvyaG
u7NlJU/b1HVGz9umLTcfcB8CtI6mFEoZ8+q1d+f2WBln8/l1cfDoX3Xr34Xj
HZY1QHq9gS14XsSBj7kZsvcGP6tJQzOt30OZiWx8whjsJZXCr+fWwYxeVnaB
AkL74yZ2/Xxy0De3t0gdRgWmWvJd+97maKoenHzeB6xIP9WWu9VkEp5bhG3h
2C6i3DLxJxRcez8wqzMSPVRoN/TELN2sZDcjoxiwxrki0Kxn1n1+RR8TDGOf
iPE7K4kiUzVIoGRziSP5vSy9BqBx+64+N8RvSGp31ni7KyTvnwyLRoMw6e9K
Rg/81kvSxfZ0nKhGugzL4qu2kAXcwGmEo3TRTTB+hdKBssyCxa+/engJ0lJZ
BDCZhc1waJjfdPnMN1iSodOU0RTxJEPeWbDbund/WY6QesPgLM6YZUVZOkbJ
pjdZmBHOJLPDiRS/PW6p5PKx1Kwo+INfEO6+GE80hcRC2bK5iBmRJHalNehE
rNE8SS7mUhHbhQ5vdWNMxQjV2HyuzSqpXS3QOQUYMzJ4mU28kAwNlE7nBr4k
ft8T/wNuWOiQ2+Yuv+Qm64VYRWSSdw1Se/x4v6QLKFbLn8W3DojQoL5c4/dr
H5rKHZnZeZrCA49yhSQkCpqzNJArevfH0D0dU4s+sR7Ool+BA00nmw+Po5nh
+fn7jTfoOJZJVQO2oHzzklj/Z0QP2kAER+yUzHBy9NtahG+3GiuUMzB/lvcP
hkXRd0qO0FAGRqrtDkeE+5W36uZJTCM54qKhF6YZRdOdNm4x1GYZNih8vGpM
lwAbV3oDclxs8P7cjdAW9oqTBa5iHHhK73WduTlp4xOi5bK4beuW8VNtbSxD
Vk91QZslBdhgX573Bi9dTFX8obzr1vQU2vgPgAcjxXAd0X2W7+kwmbEX8ooU
vOg6B9rAiD0ZVhG2VUgLp5qM99Pe/kxP6GrMWYzuN9Wx168yMEhEUZrcB6VE
JKr6rKYrXyLdctKg3gDew6+iiK1T3JX/DatDqhoQmYiaDc4q5IN9RYoLGJTE
XQMKVwiZyZIglIU3iv2zcoV2O0OH0jy93LNlWoFn8IKBNT2iak0UZbkGQeb+
rJwRuXt/IEfdlweM+Q+zt6tDi5BRyreL7MeUCzI2+txcr0L6lpHgb+xRmPMz
73GFSb4S+jP36rfalAhLaUEv/WVi9ybEWGEpRXoixzVUBbYblLW9Op0PpzrR
dac8kdif3C5zKbB2tbtWKRl/nAM2fn01asltzSw0PSBHQ11N2Yd2Bxsi7BG2
gUfHaaX5YFSFF1b3A0p43ti9xwIzOA18ldVtvjau+MSs6uwweM2gvqOeSeS7
JWWtiLB8xnIwu3EKOjX7EfooADAfyd9hMJnYnPgbCK+iN62aK9VCFpvZwJmD
1RT9u7TlRKBuTL/lXT2vKxH+T1aiTby8JpIYsHVT6XCeukWNPRZEQAHWqGkO
PrH69j6G1XVd3qc7JnQLs0mDYL+OjkcE+70W5TWD/EDD40VAPza5L3K+VWz5
YcQUSiK1YeSjcIp886fkQPe0rFsPqssjlbTEP0O3q2po/bnOQkVPLzJmB7r7
yHh1Cn4vatEuQ+yD37Ip0JEu5/LMuRf3nhjaSI5qQOCJDUC6h/eZ+/qHOWuv
bm6pFVgorZEClCy91kd9mi5BYYTmmSoppwix6o7sXFRJKSqG/a/qTcVDGKaJ
sK8mOEKkbaivCBpiAWjG7Bw2VCAv0G8sK8aQYQImk+4wdJw1s8mODlQQuYkm
TQc0wWa9NeQFAr/TuIuuWldP+OWegdMFPL5gecKaOWEMV1816B/+aXMpzi8z
Q0R3R67nyLw1IsuJI4RvptDkgFGRliw+EMdDcpjiYazd+L24VAmndGimvfA6
0vfVejRia0hrG5JvpkdmEnzZlwk6ZerhM6vYd9dMoOhnMZ9pWHZoQl1fWa92
OCxP6AVUowFTET1ALUhtQgO6NN2dZnmKmRP9xHTSVZxs+64pG14W1r4V9WR6
aKRBKt9JflPcv3GSaMI+dS0G7v3v8GSbpkTmY8bdLBLJBnPDy7yCGu8u15St
gZjMGTVGOdFAO2FhrBNt1057qBIFI7UP31f8eqTZgoM5eoZ1XgD81GvjqrwI
UctdjM1CMBE5VcK+zb7WMyYgumJJyqff6tDCzmvTGfchXYy8Q/dtGJ1H/tPa
CLbUA8EMbSPe4EXANPWm0g/C1zNe0OQjKAndCnzKABLbj9CfLNxPAz9KSTUt
9nkUhU0BcrHJuAcy5fl2qQ7fEQusB+EGeQHScLHnEMQd9++eXMOH4FQjhM0H
GmRSofXinhAhiMqsYtTBvNg46sx/zJmROEiqVN8u5V8lyoN5FHzx9IEpUNKT
8Xl4x5KEroLg4vcyC4iB9WG29Qov2h2YzkET/5nDxk79Z87v0RQi2jl2lxb6
Jk2N07xz+pbwoHSQVds4df0nV0SdVDhDKYaqpRCQfslNcE0BeA2Qu8y3gxTf
W6a3np8SHaMqP57lqNMPeBarvko/as+67TvV5hs3nT2tvxx0DBoFo7kvLH+L
qosIdqipgVlkjnX8g98z6s5wZEeeR+x5I2BbZlQDycmarL1fMDsh6S07UexM
7iGTHezM55ENQ76xOO07BCuBDJ29ZzFV44YapC2EoTObU6DDN7q++62h0RP0
DqDsQA8SRo6nhAzurWsejIp6Tdt8V2Jn1OZHDX4Uobj+TKwT82B7kHMlgjEj
26/5ehK2l17EEgTb5gnhYF7q1IqwW9BID2eZ3wQvbHuCYT9Dk416x0hamg55
aK/AP8XTKNPL6vL0fX4DLJQ7bordkcIelTXJkZZmtUni9VrCtNEBMMrEUwE5
WxBVjH4BQX33V9EzS6fXrpTpCgr0cGJqutJzW5U97dBOqHUpNvraQMiin/Dw
Q/qp3mBRH6UTY5JU2Ji56ipFqo/pWbQFsDAThdkk1od9zKqa+JTNGSmCqsiY
ahHLNz0YfvY87Fah3n97yRTQhDSNtMOpm6twjIN4zCoknbb6ZC/ucqZDoHvO
dgWRUVoIU9SVFD8/yJIeR3kiwyHxJPcBARqDmU/ErroA9KrOsIbcsVFRgMYj
BLuurBhmwL+7XN65U2blWXPx7GeP/7bHPF0NrC5jPUw3rGogVE9DQ7Yw7BYU
jHA+PbpoRr8mTulAyqdrf6PvbZsO72JSwadGONUPmxS7IHFzX8jX9BeP6OJ/
xW7zq6xvoKRjMUA5+ujbEZuUyXUvO3aygwNm4zwYNsSBH8FUXV+1udc07j1w
BHWR2ojZ41ayOGgKtn6dntxj8y9QGR11YM1T5BaNjt2oRgVfTJhSSpY9onDR
r6VRvUh/Q66IwsWqeMPuG60ZeDmesK3KnBsKpgEIf6G00cINEE74IVRL3qjs
bow+X44iDLPdtxvZRNH0vk5kw92DQUCzAVho0yYa+v2yHTpADcog85QRzB3h
KPhPvmg3tgMRxcXrAU72XRvd/Wgf+BIQDUzpPmmiUtZFzlWlAlMsb0qBoo0G
MiMMT91wmRZM7H1OG4wUDd4wT6F29ZKlXhq9VcPY7OgJyshfEd4hfNxFKCAt
DpA9gfhZuefb4RLkk3zXNTB2IInQAqvz2YA/XJsfBKoZxE2n1KDW2dcnDjnm
YMLFkMylUtFHMC3BZctAizkAnqQ1sYEnK90kEiskFBxdnXHNYUCR06Y16vwM
PpbxpYFxJ4aAwVicisbxye/tHzE5jbiglneC5zFfV8mm/AlZK3yuzP9Bv/+n
uGDc+AJG52mEk7vosKxD/VZiGX05c8sN8eOg2h/Eyj3gw0fJxqaQCv755c7V
dU3lAGnSdx6AwmvozWk7uPpKtOnwbfFQ4glgVPmiNXusBX6GjRTe/QQPGeOy
MA2GURuloyiBTA7iyb4F/tM9WF8TfYthlpOWkiNd2e47DT2w6gx06jvCESxe
0YlgWKLg1L/nDSrAYg0DlJOjOeCNxj4YNdHkWEvPh5Af51TuKsVuYKgOk4cS
yJs908df4PF63ftf0W9MnW+nlwkeigiXeXtOmLlxIVVQURx3bhRvSZbZ4fNA
ucK6WBH8USbRu3MpVHXkHZNr2ZJ2qELa9TrvqdDNY8sPkz2lr4RHeXUu9KLX
aDuaubyluMfQhXVpW3cQmIWd7mmyITXVOM5DodsjaPJTZDT61ztIGlKdcTnN
c0Qa8wXAzqocT5jWceF+XC4wfW1T63bgvE/7mw7aquKfYS0Uu64ZFNLT0YDc
RjWISQWdf10Da7nomEVRk5Zq3qcOTuGsPIo3mjeQSw/FlfY0GnnW5URt4PUs
Gbnka/zU9IoLF0ZVqAdOeSGG2w8ZSibHJEv7oRADJ2CjEACC+V8ribpAyPDm
CbjS+0slt0o5PTrA7PjjJG+nTd6SpQfnRkM8MdFtIhfXG0fme170fXEFITpP
GsA20b7YW/Gikpf3eVov7yUB8TF4yfJXjBADYE9zWX3pB4qJhzvnm5tefzjG
FzkLJ7P4rQy8SYz+DA8CKb6Wr1I4C+6Iht3AJM6q+pV06PjtapPxZkMS5uYS
T5I8CAeUBqVBDxElv1+0GprGUK9NREhXR25gfj72anePG8OtC9fm5W9FofCY
yTpikxQf3tozP6YkZLQQCrGjA8e0iODqbgy8Wi1l14/TRMaqGW94HhpVDWFx
apG4UPtIADYnMOOBLPiK34qg/lvhBTU/tYs9gxk28Pdf3LuR8wYNI3yqr5ia
dwGy726UON/kLidv8kVIan/LJJynaU5sSBOwYZ3tvvxB/DZ/ewmtb2QQSf55
T5nT8UEucMBPTFtoMbXj4rooXQGoLBNwPNbkMiKfksa6Tm14YwMtiRpy3xlu
KkCubE4bPW09pkUZ1+4W/Zm5RCyLdlk1eQIoAnOyJjXlsuX4DV98cxGtuwnW
xiR9dCd/2a8xfvHMkS19tZ6upMOtz8h3eLkV1gZ0XslbzWjDIT0fZi9VbMC8
6827kgpKcAzCuq0BTeX/M3/fp/VocU0cMXAjf9fXhXl0Gv7xzjOr1P+mFPK1
SeTeiq01UOL1AZ2E1Irm3YnQGh0CkTFXpX2n9/sHlPnMq2J2Axm+IbCgbIA4
DYTusJenc7mQOl9sAjJoXklW304g2z0sfYpzi/DlUyrQCgn72eL9sM22DG8q
6x8KXO0La+ABrGs1b/KnvDuBkeWt3EPvW+vGAfQV1Ld2GjQfs2eMQm5FJBDH
nEwc2K+l2ybNFEZFgKXUKhcy1hbFMT2vEoSi2QVZJ904GfXnJeZqzPaO4mMb
Iggs7yp2TJiwI5J00TnoAsLrJxxAMO4nDDZ6ysNk0ct4lYjlkxKkq2E/86n7
YlcCHX5wSBBLvvMiR+/ctVXsfhW4hQnoKcT8hGTQ9ySCX42sdFMZmUkVEi5q
gSCVcmwwkmSkJVdZNeT+r1JD9r4bFYnuow0FKBez0PLvKpNnQLp+3OGJ69o7
paWOxDgIIAOCcNm+uSitHFls8vYnHVxzYPqV7l1A6N6I7n0eR7z2Uziva/GB
oFd9OFuVz2ReFhLQXTVLV9pAP0yPqRKL384pILjn8r/949atPjtWmI1qy1Z3
108po3lbzBVwPJxWY0aSX7ARLk+GLrYdLoTci11e0ZGqz23o/NS6VbhapYAy
NxO22wfPPhqaW4oGPH0dXyjYQswBNM+0jMkbkOcdB8YZIKu7sT1YU61TjVPR
BhPOcrrpEjUJ2FXn3JZnFUy9/uHLcbIu/Iyrmd8C2ODesjFL/lCzeQ7jB7Tq
BVSKo32NeIWdl0nKfxtDS0n83dI3mHAkPKB7nNTtsTyY8AmsSzLsANdg4O2B
7VAF1TlVVdFvdjnpDAsa/nMWwTebIpDS5bWQpa2ElqG57AfJC27wSx86Yx4D
jX0N3FnhzmNOKP8OmJu4sIGJnim3p+qI+5FSjmstFyhACo72dCVufsbmf/fQ
k1Hwdj8uJji4QBgZOu+Na9pOhspLae2nzwYQDFolxxevImP4NnkSMr8hbMKI
ksN4/dvOKBtjVLxydUFSYnoJusj8Y0Pknc0YHuq3C2p5bkl6dH2Sg4AQJMvW
1Yf/+cd/fiYTzvKxAsdC4vbnWtWvqrkSp2+n53Seu3LzLsEdbY94AsrpMmUR
d/nQi2Bci+oChTMhjVquGCwKBbXIn94I9w6XW5reIY9TPwxCDQLVEb5YdfEy
MVB3pZPqR890etPGOibYj2iUi0UYR/88MXPlZMatzrYqPU55PqJuHyZ3AAEb
oLSEkjs/bWIt+sOXx4jSC9GjhsD+btDt8haAzG8fFl+GMKTLsJmCLOYFSACu
ymSfdmquE6Su6XgOPI3nck80F2NN0jgJdYEDtBgISeLeReeWUYdr1kSR7VjD
kEagAo8GRMJldl0urUVSwAMOwaLBNk9evJ848fAIXswLVPUdU5y0RcKeU9rs
Ff9clxbCFbTWT+BaU3bLhnY5rt1ke+P63hNnR6NJAfPQtFGAxmf1yRRNCior
Nn3q8NyGt8JDc63FaKeLuFkPY7JP+/J4U7quG2puqp8CJJWZUnwaGlsB1ZYX
GdiSAzR/N4jxJ1yjGvnxxvD6hhGiTYtMg/hhyD9bSGEvF6U3SO8ogrW2zygV
OJrHfyNBrgaSTO2ZZrcyw8oF1Xyy0q/yYTiqSIlDFgtMEHFkmFJkqpWkJ7dG
KM/GxvHzjLH3Y+hhkzYZDmlXGBGQp9wA5zzw4uN+l91iwoiyj3PalgVcKa5W
4w517hj52ge+Qlx6n8rlNRyDmykl/3/FOZohNj/RKA9+k8Xhf/rDz7dCFB2H
cDP8d7OcIME0EPTmYuv/yNHXOo5lqOhsWjXMj50C30G7yGclK0EmDdf9xIFS
5fd4zVehGCwCfUGeAABa47y1at5aNoWQlokD5gydcbril5AMAXGUD9EKwHyq
VcR64DwgzKzRTdUfrd779+Gwq2ONnELKyrDhiCUNdjUxgDypL+/QxTn7T98J
J9bc2kWWtP81l3eMUwDjSnf2EajbfhRAz99fpo4o85igAWf3lJ4GlgvhwfJ8
85t+MsLGDDgjpk2g13n4GXLV3VX/cpsVqPWsJAnnYFebS3fTqqjfy1qoX6kW
UgL/YoA7gtKXWB6aoVmt4x14Ap0jDaiWca3iSNux/m98xiTSd5RQ6oKw1N68
9vRL9ioRCMap6XrXRSFW6xjkt459iAo7oSfYr7Cu/91lB/WHiyxflEVaIooR
M6f2f/Wwg6OHf+W3j8bTA4wEDUg3bNd6QLw6u24xCeryhKnJrDzqEKPod8aR
9jqotl3HtsrF/7DtGohfuzyiU+rflAwEvhd0WyKDWrExFWwYlf7+voXmdz1B
Uh4KDQl4sB0UDNWEgbcGm/V/5gwiADmzraGNHZeJCIesNg1WsKIa8tUiqSMt
K4VV3vDB3wfEbCthaP8jdC3Lx1FN3jKfU7EEAbevwywmXxXbWni/DOP+CjVm
Ti0dir3xMIlxTKnPo2HuIZLQOsK4yo7FIQF6TACUGh/HL+pLgY4uk68v2ho8
JIpd0bNaaB5yyWt5xMlAyHIHUDNXfj9mI/+ULk3x8EuU6u51/1FGSkXkFI4A
FMQqyMMpNASBveY6/CVb/EIIFUz/FlcC0FfDXdY+JBhybuw9XKBbttv01ZS5
f9whEnDBHBlrWPGWMqThZIsJ9uFPMxnUxbxye3CwUHK9+RGkLoqqf5fkydDV
saqRi7iQDmjyvRE6rf/SxGwBGVysEWsiZQbGApxC40sUqlxMhgCW1Aj9v+w1
Uxc35OOLewWyJkFdLirRrP82ZlWSgJYlaynB3cKXLZvFvapbc8AO8aoOnawj
Qm8vFlD8RoCZZZ895QC11TGAVXA7ypOz7YdXkoc2s7/t11Yj/Rs2h/reMjMC
tmf1vJ88+EYdLWWJHZfvP0SXvtcs3oplWZje43f6rwY3AoH2qYno8Bu4D0Ky
JHY68wvwIPD55vNW2glkjaRll5TuYYyN0OdeC57CnZaTqvSMZQWCveUPfths
F8ejOlSQB1WtBaIbqBiFUUHZlHDR8zR194o8FNZVrf/KJ4NUjcNiLkOa9+1l
tzwWOZX00L10mR1mqR47kNzusy8g636uKKeK4UcT5c5K2m7cfsmCeabcgGqQ
sOGb6c+OHmBJR0ViYuksV5u6wgEzyS8rvU6yrBf1mYQBA3/YibnXWyupWTVA
sBJPdR0yKyiLA6bQ96hO5sfhLEMPJT4sZyxONEy2tipaWyB/xtZzgDiSHDVG
eSe4VpUxnMwpav49iN+ODNwOzAfon+ixjA0WmhDTQhvMJ5DGIBu+XpA5QC2A
9qCWjytrHSKJDS0C/LUG4IK8Jxn7fGCVVE90yQixeQQvWLnJ8sTnRWwzqKdN
NVslHWxPLjcW3HD2C6GC7S4fJLZbtoniFFdGvRFjeFK9qEEzpyYsPswfsIqo
1b8jIB8DnUxjLZOrASZTxdapGqFYqzYOnBgzeVeXgjC1ZZaumZEar1qNb7SI
vVfTGnLuy7kibSA7GVUzbW8G7YDpnmngXPurAMxqyqpL4v35SuOq0HwM01F6
teMggAln1NelYRf3nM6alPou1td+HzovMLkQo2FoRIEnOJ8gWTmgRfbwlrrG
I0wGvSrtFI/XQ+rbJwAaDu7QvMU70Za4hFVwyp/EVBJnAUjO6GzIhXarvaOF
zsqgyqmuYcGHNb95doVPUv/Ory40zhdmzqp87m1h8rlrQYkK7p5o1e3fzeqy
tGqASHgddRP8AywvfwffqFfJMDwAfsgoMTVhdDroGoP2LSXI/XcED3Iq1JmC
J5CkQQudfv9A/E1Mn9ahYud0bhZQ5kHtvykYCh6lQ83nBd0qCaadQwU6aPRy
ZnVHsjsseyd3wHaSL67RRrEg26lFBgHPx7+MU/nRKqtSpz3m99kd0qwVtl/h
fxtnTs35ti7Hl4KBRoeunS0krBtklxx47Ka3z0bn2/SjmyLFrLgXKB5vOuLw
P/5ynVyJvaWYtKgZpixbkLrez5gA3Btb505eVrx5TDKLQHLmZZd4Hw/GHiIg
lzXMLqKdrUg0+YcmnPcnpUKQo966MpYJ9ltPSocwWh51YfUShnGw1RDW6m+F
HHqVi6gKwkErFNi0Vl06AuSPOSwqUbpsv4BfKjreVXHKBB3bS1kt+4m5n9AQ
moOSsypf3OQT0GmOjJuL32HUo//bqR78gE3qW50Hg9NEBxm+yfKSxGWfLzQj
nrTttvJnleF3MfBPxkMBug2NktzZ/suNcqkva840x7C9DOaD3IpJtd7E9v6c
FA2ts/OuLgmzOkyvu4ewPHRWKbQJdc72BaGmExqZLsHsRHYDJFGz1bl8IiRu
L0qfj3WzKq3O1T5mGf8XxIKTTLPLwI3Q27K21odf0/S3gTBQ9kjfeyFNsjUv
GiukyNg60ENf6SAL6K7qbc9if6+xuIVf9A3RYghbsf8dU4OZqABhS6GD9A28
mNr7pPpfbP1M9EB9y7u3uPQMvHar3kUDehNrsicC4e8JfwfKexvNN3GO7Rs/
v41Y1QzE87SuORusrmMp9JpGZ6DHiykPPro+cpN/Yqdo/lq9ETZChKC1JYLZ
WCeSeLHXWdjVdQzonhUSlov7mFvfbscG/gfXHuUD0cn3d0F5wnrA3sHRTTnS
WtMt8/AfhaZ0TooSgIY3ICrRJgvHTjbBijfi8kgQ75npabb/vjOu+ggPjHkN
Qd06UhCHXIhwH3qHhDxSjXGjWCNsZdb2pXtdi4ulDkqaDNdjFrix9OcACcAD
aflVCxytV4Y8XFa2GUbIge31RJpnp7zNDPiw4F5MND5R53kG0fATBuGACyFK
T7R4iYwpvHDjyJucjPJc5GnK2G9LACGhY1c2inkuKsfLpEMDkjC36XuCNogP
+530kXjhzUpSjMU/auXwSuL/OEKFjAIwBiLYYwdSSfj5JQjUi/KKDcNg+/i6
CBxmw2K3tgS6APxEFIm9PMK7PXDpiCuC6sSXiEAZQf5wqnEbWBLxH5z2w5hN
iZ7neYongpPCeRacf01VeGhEv22ZruojrsQODsXTam0B/JKK/4dw5M5PjYbQ
hros7SiTAIAVfTG+iHXd1O5l9fmJbGg122Z31nZ7JI+W9KRL4mRosqTxGP+F
r23tqvVVDDvmh5mx5n3dinOW+Xh0ggTOv9wkY/49pc6PYi3fi/zVSv3CwRKK
eJV4BhBKjGCZ7f+goHuQeaXqpffN/BixibOKfGDcJK9KfhUsy06MlT+bMX8B
TAK6Vb27Bl8tiYxBPmGdw9GVAAdL+DZoRk3SOqpiSJJczSB7lstb19wtfpJk
/Oy+c5o9tYdnMowNsShiNH69oD/3R0hy8Qg7Z4zfXrQJjzYXx904CYNgWaRc
TyWRShel4wWg6oLzggV5RQ2/MevV7Nljg4Ee4ua5Ea380EEewhskgMLXTeyX
XP150X0W+3hMmPIwGTOuqvFV8Aoe4PiG4XV9n3qvc2UKHqdmQ+cseD41kLbf
y0c8jTREnM5bnz8fxyByQqZV7O09TfACq881XpzIM8MICSaQKJeL+9tczYV3
txLKL+cvupCXY/S8NFs1GRjlZ/OE5hquEM8R6LfQnldAAJ8LPux7baEQz2TQ
40W2flyrmFK9jNWc+4NiUgfbMZZFwdylgPiLSlPT2zOwSDKCVYbWR0lfDPA9
r2AJoYKacwtMrJt5KlFL4/Oeny+urHeXEKOViPvm4dOtyMsqpwO9d5zosfYS
Esu7JOY/vu9waaOB9pQU1DSyCwS+vu38TzSKBCdfF8LS36g/ER3RTE4jouBm
z4LfteP6+mre20RMTsPmrwZkTRTcpLF8NINa1FSBcb92GG2AuxPxoEghXPB6
c8Tgzw+/5daBl6aDbOeJsGKsA/5pR9FkTIcJW/1TcTszf4z/t4JtlbqX99l3
ZssueTLUf6pQDXfLxbnj/qdHQYT2lnGgkCQMSzgXx0582ARm3zSiroRdDsbG
S9FjUtbKR1q3ExOwa5b3LBo0u5gXA2LkF0iyyqmzvLzw8C8JCgPjWWHWK6SA
W91kfq9ErF3aey6oBB+vMYY78L/9KdfxyTnnncYHbO+nW836SdwMq5gcr5MS
K+0E2Ana1XGxghhLyXUzfH30glvClHugWDPx/mFu8znQckeYMrcx5N06ehIx
UNzKw+5Yy47dP/64txLtjk1E6SWicJkTVRo4RF/j5WfFx4yiB3/QDa50U69C
LkBbus+dfOEQb6k9CJYdKTdMbF2gFJJ/K6kbJzBqfcBjVtlNleJofFjrjn6X
P+3o0Okgpz+v2JLfowAjPqi3ZuSvoCxlgGnl8uXOdAzs0x8No6xxoWN9AYbK
iGngzmOcUDVyHfawGMhshngayZyK+BngJa0ZE2e9FhU7d4oN3+3O0lXzC/3S
L2xD1/aqJjEW8DDxiHs2L5yrmLolN+/7JuHmau5xRo9ABtGVgbVMlI/lhm3B
u40CRbKZ/lq/i/pDoN25Zb69oIHDoyr+eCDwdkmFqSuFphG3zKyJOmcPjosB
0ET9EbNETtoMWrSHk/YtujwTTqXV7ygXsT5wCdlTr9lzM19siiDJUvAp/xLk
EEo2f7B7xaes7QLBPhhuWWCdLcFPbKznL5YzoGukFQGdzQP6PsaVHWqMJbGD
XFbXv6280P/RgAYAD0VbIK4PKoy/sJbaSMOsh0A5vosVbknmhw18Jeoyx/4e
rz/MXcfstl1/jMN8dxNtpjSNR7u/KJqcgwZfTktudV6BeB+NLJRT2XWeYBnh
uyWK0L4s6Qu4Mt/1tF5QfOH6xOpAzFCJIisweWXuiFbXDgEU3zYrygaH7EwL
FF3ks73k22lehShZxnUYHv3zjnp6dhi+EmZDPGZIw/wSrd8+W/6MvsUvcGi5
R3IHMo5503mudD56jiExWqY/2p7Fb1YIx/qq4Fr05TUNqmfj2BtOpSBnuQkz
jB5yePPsDRvVCkHKtRUF+/uI1csCuzRre9BZlGEKaBWQ7nodUrfCyE/QJqnM
xtZm/uQJy6fzFmQgzj4WnE9zHzCjfZt1sdRE3Eps32p/rTT644atNsvt6DGz
HwTePQEkaMvZg1sZLqc0jWC0QMoGcufUR40u9/5d14kQKwT4q2M3VCe4tWd+
Fre2dlQtH7AWQdqDmxWm3epE5bqJ1N4QTAKnpCcacICocPs0cn9/RWGrEdr2
3/ID3epds7IRXDJNAA9dXQLouW5rdgK36OMY00fkMVjCFJ0dulJaWczVlkQP
FqY+Oqn94KfOcE55SUqWVO+DohumtmmmAY3O/QNsogT0Sl5bw3JXbMhfECxk
2AB12sIivS2cLJrJQP8qiDBF4rQHEpHqwDxNWRLNxZitASgtaId2dfcfF6Kb
N4fFtzpU3+7vR/bYJzgJ34Y+vjN5hcA4qw0zvOFK9Yms4v7ojcccK7am+Isc
Jcc/VoSyVNTI4vPuldjJG80A18ovWzxj7Sd7LtCdw2a+mh8JbjoTiEE2LItJ
Im9NajQpMf4yxHXUlL0UX+qd5WuRVm3OB5n0ec0U/+c4XBWHeQCc2Y5PnKGO
dy4w0PQfIvE0VLibb827lF5X6QKnXZX04kxIvDE6F7zQRB0e0LSY/VpCoLbE
IjXDvY00qNoK+k3EG9pHYsW6R+nKQoR770gCUvQXG3NTgN8u3ZzTfsZpQnPH
Kwe4MplJ9RrbkWeI/uL6Fofho5tvOKNObv0hmgSbLkekmli08LGpi9uNZn6k
uaNeORkivaeKvaI/I2Wyolb63aRIGPCzuCcOmPtMlEhOE0YT/v8/0Bujy8gi
WuzDW5xsonXfNG3GX0nytRh+eGSp3Bahbwe2Q2YTobwZ9j6XJEolXf6cUvJ3
ONr9ktDdRsIWcnU7yIzsB2HJuEWaeHLSgf0h4fEwzyRRSCrAPWvlOHibHBNP
zLquwIC3gGxcKdIKe66zxK00J3xzxkEupqN9so1SvP0/OFMZfb6KqTN0oGsB
z1H1m8TaoKHjn8EkOPm0cvrtmg+c1sAV+mcRrM7wUbgB6bElcF+XO5LBpqVE
AkXnIVF82c5jh2ONSoPE58lGsPOk/3gu5TZZ82DVSNw38p2reMCvSJjGCfl3
OJAmY74/Vc/0wajwZOl4Casn3ZEyQ1wvRJ9kDEA3sfmU0eYgyP+byYD/2d+r
turvarQRX9JZnJv/EC43/NK1/7yUocpttqGtmmvkBSkzrRs4STltw7z218VA
/OOACdPbey9XpV+X8NHGqPlqKyF44X49bd4GWZJ603drO92hwRGMzdyF82ZK
ZKwQ5QO4nPsXSpkTGZRg7oZx4QdvcDLU7N11xnJUew7+W0c44JfSYSvaUgeZ
6MwcrLyM4XnoSMMfWVOUBt7H/96nnkAHI7L6mBmLMTXDT25Kof9kkAJsjEri
ytY+3e0yTPRv2Xqn1RGtL5A5SV2wnPO7p3b52hxNZRjPWkeds3i1ub/Cs6cl
qkC69MgyTC2kBFHYTQnGDLVlMWPOC8HE2XAwdR3oJWGGLR2rMWjOvK/Aypeq
z858/M/6dLNg2W7JiD4ZmTkcBDYPZK2ObJBzhfyCrAT7ccQ2YPzt21e+honf
A5OSmrGYKPbr7ug4uGSncc/33qkt6dkUIp0vn3LrmOivTh2jJLrVtF+C/asz
YnRZX/2P2bvlF8PLPt/JLvLwNObiBJaqewLCKWH7wHi5tLMv1yE+F2EOzj/8
qcSX0G173lPz6u32apbQxFQc1FwJxNzgqGVI21zk+iuGila6aGnZUCencPw8
8hjf8gGoUXY6rc99sJEjp9+hV2F8mEOj6Z5uhOgqa005UxmiDCpLJV+XeFbN
q3pPfLhKWQVDZFJT/FdHQiSKsFaIlUpCwglU0xwC0LGbk0hkCb1M0Ani7cj9
7cE+wtfzFKnOhB3N6/d0Ev+/B7jpjafMu9qdWAiulXqP/LMl8dj98ij+LTjI
uHOY0Kwf1efGb5xim2b8efp6KBNBSiFZZzQo9MDqE8R8nz/uYVIn/eRWuYLy
SCJgARgU2DQAe84R5Cr3hDmW13AJ97F9ixBqWaPb0QLojsSNB0ntKSYzLXs1
nKwiMHQpIGwEV3MG8Dqwu78zzEncuHCppbPmWMvTBO7TgeXYCzphtb6eL/+K
9mo/9cNEhrOccU0nxJfTMf9f03c7qB59IbSoIXUvmqJZFiiAnk0pGHVlIjEp
V9tY3ptFVQ1NqfY5MWobiI+TrcSwPNVIFsJRSxhu/uxQJtjRTbPlCSRkoncS
D/OjMtgRsM2D9OtLhMgSEeGzcBoSHRLsbWtBW3Jwk30+q20ZMyYk5EKFzPMU
sK1IxlXVvq7V2fjnLUWgvnkdqgiMCHkY1B2uNzFf5GCgTotgxM8moGNNaddj
lyvzHDGUOxWXAuNzdfJXTuIRLeXhVOxNgFPpgUIXyWH1kWx8fSH3OwvItnH8
SAcF7E2Rls5RA1LQkcFvmmJViIrLp3jcoz2lPMF+W6gKi76LYijZGwAblo5N
3rDbwIHhcDfsr7A/cRy/GMLyfOimeNNPi92qMEW3Y+2Uk7LvVNwgHe+GVl1Y
PrBQMYY5JYHJH91ANWBoPXd/8lzOJaqPHIpZnopkjToCe8ozkR/UKXz6UFCj
fG63ugBbCVtoScef+uKnyFGj/SkUnEeplsK0E1Gvy0EZ4vZpl78g7rR2XifC
To4NNtFDm13WSJ4hf+uUVIWy+shR2tb5Zrvu9HTV4zjHYxBWYjG14zmeQQCV
s9jTljXAkFPE9YMW6VwroDOHZTnbamo+97fdoOboWIPDxF4DHWslNRuaHIJH
W+hjZ4TNc/ZJNh+FLQW+fgGkXlxAkWMcijlp+If2JF9zsCOPKhTr6jOoVNox
znDx8NBwNqO3o4QfwjkYWpW+fUnf8dyXwrhZ0cSSx4wQ61mSXevjxrnVIYTR
Jfm06eNnOEpLtZBFOEN/12wewHMViBPXt8J/qkj9H+LBO3gydvIyikqD28Vy
9fMUtiwlTU3KD48MGwINFwgtJGM2nanYtODfZCprFOtiw2COd5bi6yodqe/w
GLlTY18iqpmhyBe37NNfUhy1uhrzxpdEUEj2ScAgv+g0jaouYjlUtVxDQl0S
qPNJwWCBWIiJfapBXjI0oNjMNsLDO77B8LuPBDdmHztLNS04OVx6q36a0wcK
4krLtbsXhlpAvtcBw96b6Nnxa/MF7OVU3m5kZ9/53ooACDa9b17WNWmvcD58
cWOVwetuRETZTDZkMlJvG5O0Bm8yxRHugISY6ojPMWDHEki8+vvqnI2KYa2K
6b+kdogYthe1Wb2Tfwe1WWggw9XJwRRFgb+V/OBDuc9/vCZ0a4k1o4AhdE2N
GlqWXu4Hs/bYQxJFANUGHGzjlK+K1zOsUkJDmzWvXSafyfJNlhsFn/ER19tL
7/e+hXFcP5cgNLdrCDP1dICrWEMIR44JbQp4HEAlqC74c2Lq0txwwyGL+P0n
KMKMcflNGXxWblToihB12z7ZXCFOu9e6FHJtmNeZJtzGd1zQXZBS6Z7/k6oq
H+fQseC7sniI/NYOwLxLyrcQzKhZ/9PifkxsOjiH9bAjAfwtjiuTPp+ccYlU
y3S31AGAvsDW7fseP2np42VmEIukfNagCuZnz8OOaxLRaKuipCLRGMxw0Ptw
agKJUSoNpotaTzPhYu+gP38kCzCydZGighHLUo2J6YS69ICPepvhbj/2JXe6
i/JDOdDbqX4sBa4/d0ANXEsd1DaOcPCItnHMsSOShRmDhg6wU8Jo+qIGxSK6
AtTrNEzndgaSo0eE8E63N+wYXH2bNQHnezdishnEiNuDWzdVYsrSy+I6Aew+
GBzjLHbXPhteBwMKgDLrqrGcdeJbsUta4CEQ/2N+FkCghLnU+pLZjzkOwUQm
1O06MAoOxLWbUTaGgNCD87fqUMUpZJMMHsVJ529Zgi1kLdVKdibKJ2og5Opa
hKiDmurN3pEwXXkVNLMrcT+zkX0gjnDMIdFlYKiEH1yYx10UQZ/BC2DGWXq+
ns5spXPZ7Dge0TVLapTasXx881RnNmJi51xMOO69tZpZdtkSyEoFOiGQfLDJ
+MEX35iuxnxdzfHkaiVC6iToFF92jmAwsZEE7auezHfIkabsKEXCNSChxStR
5mN+MaTbHqHHzBHtTUlKINg/MkRAkWJth5wgeYdtbgTfcnUly8phEHwSkruj
5vrSRb0Oe2WMjEUIdYLVqHugDTb0aov1VHroZO6EF6essASyU4vAMAMt+gjC
D31rOkInL1bW/dx9/Y86US8ljhE0gRQP47N1C6ndrtzZLjfmft5Z+VcEyoW+
NVVoGMeHFj8cdzcZb9Dzwqd+8LPVD/K+V60aTUEhUtwftSTOrjgnBFzrxPGi
/u0eiBtOv+B+9b/i9D2WoIgx29/GsZ78eekjJajRvZgNMG9hbiTmdaGM8io6
ZbW7WY/DhgfzRAuFKu+sMlntyjLmtCJSZcbwf54JqVNT2YLYlRWtPh52bB3d
IOHatubyUVV6B1F3e3gkLhGwzh9k65iCaSSPkfcuN2ibCA0oMBf0yVcvkEbG
hNM6f2ws3l8e7m/k6WW6OvRSzF+dUz6Bu2b2/K4CR41ZxQm4QNtXaFEZHTw1
bjd9s/Vnt/feDmA3BC6JZ2hXpQvI/+33j2pfCitaF5Eae5Ga88w7Wn2CmrdF
/dKOHBcAaCvyJBaa4DUsMC0JHe1ijaP2EDVULvbtEcvw/9BDyRywAW5HxMNV
VQyOQtoLy3CSsbwRsx1en9HWsUAk8YfhkMJSL4srNE0SxzUFQnKj/ZyWWBjC
QLOg1ND2rOTZCsptmUqqR9u+1q/dsMRwDQ7ZOWaD+mJTi+ffRuAUG6aNx5WM
C4R5WCGKhGdX6/iDNuZAQbNdi/65CJ+PZLkidvzwu3rR9ssihtw/GSBqMS+L
7X0cAju0pBjEToEoG2ADUdQ+wJqujbwodudKuQro1J7tyVBSv1bjISGT7sr+
XP0k3gyPEbrSQepu1YI3ZM5RIWGHdh2ctfooz/A335C1dHS6O7Po86njSvDw
/ANkQSYdW5Znx9UhqtX6nRR3nfIQFFa6sZ6peBBh4Qhk3C2aEu4vHweQ6mh/
eNEJ42sZ9H67QyWEJkGS8wjPWUMUo2m476NWFyazsHKw6D6LvrwTefbD/GKO
wGbVjfcwjxfzJx8Ehp4QC63gZ4krp9zxlL3qzPWcISt69beXFyZA8hNnjOJZ
cyreSsyYEyqSc7nbDftih07JxOQxyBObEcNH2YodFfgZIbsXSwslGuHq5N18
Sv+m1dPhZN9EUb4Tui2LJGOETKgYd56aEqsx5owXZFFYdQM3RSHZ2kRbtaRG
s8dFdWkgcijCyYJo/qrOquIdrRNJQDj/Urq9Gus3UXZt+o3UIOedH9NPM4mv
BOQKFfaYkCNBAatZsyCSmoGROYMSQpSsVkrDMzFTQCXvoT52VtNtSEeDpm5r
PqGP6kEaia3ci88N4I5EO0vM7jsYTdRL1twd4o5vTPLhSiw0iKvPOASGUbbj
XkZvwqIrMbTRhI9Uyw162mLMS7TcNxM2o1WjY04k9Y92OWo6jYgbOKR7YZu1
+EPmCvLklStlD5FLF0PyDcdtWYlrUExvCqYRKbHpdJy8XON00QLD0pzsuatZ
pKDZ9ml88rfXP8ZBiIS7Y7/7jWxvaaQa9PHqBE03ydzvf0YzaLBs2soYaNLq
Ecp1QGuCaGRRsrB9wiheZzj+SsNv5gga0Gd0P99VlCXkbcpQJFxEpgofFNSe
wsYAXfSLMpcCh//Rc5p6LXEnR7vPDhY8Z3nkfTmlvekXDsQxnZyK6u/O+PVu
pla1hh7Fs1sZqfLWDZ9QUt7ZoowJKqVb9NFHEKLAkR8PIuNFz8fQHjswkg1v
Cz+XUyytgDLcuw4o5H/Ylq8aV3sopuYAgwM3z3ifQpItJnoLbac9GXVRssu4
Fb24Q4u9P3zDovv7AuCzVJAguU+jRdGoPBXmimMGhe96hMtXsuDpryyGX9EC
fVepmWR7kPPCSZy5SLiB5ujTwSqkrWdkaykz1n8Df11U3FaubUgE60I3T/Ug
CE9MmAER/Vju4CBXi1UyTI/hZfihOzJdQAd2razKjK/tnOblOQgMA1tCa+lE
koDpNL+vq9oSwR2iMDVlypqpm56wZ2bszyP8QqgCYm+VOfAaq4u7kYaRHNSn
nyS4FyWtevsFvmkKTsTfH4mv8RFuwSVnhrur3ysCDZlXVJFc1De0iGTP+/w9
6YwRJQ35MI6YIktvo81YF2JKeiY4dnexTD5RZjFViitdlbQ0Hsdsu9PVhj+G
aixXyzazsFDjyzjnmOkBHkmDIedyRJxIoZgL0/psc72TXFX03Bv/I9bJk9Mh
89DS55YLHshoUVuaMH4BvVBs4dTZae99CxTwpGrHKXa/1I0gfy1m6tTL6Xqg
zX6BUQG6yvCCOWrrIuciW3nEwN+glENvsNXlPMgvqxFRm1te/hOe7ippUf0E
By3wvb9Uol+Rbz7XUPo3bRmFUpmG6pGMRZOKJYLmKgNiOxxvj+ofwPr3OC+Q
boiY4QeBX6OcBI2lNxwmo2ZElollvT1i4IJ2/qcI99+yBoNVOktZRKt8s6l8
mP/384SWHVvhX+P+QWBIXGUHbh+3A5SEVj5NllfIpnpdTpFs6iR2VndXgwZA
ChyWWDCZaqcQaq+WTojHDlzCs+Z2wMKm4qLF51uu6ealxKDQXpiGQNPJeDEi
/OdsPd0AX+uY5BzvNRqM6ci38m/nCgJDM0FFtWY9oRiMqHvjc2CxuUE4hXlE
Zf9NQ3A0popJ1dsFu40q1J7K6ay5bG0g1hvPc26DmytJtXIwuT4AcAjPuF+o
NTOjjpx4dvAA0yBV6V/8H58aO5PUYbC9NnRYQSllKh9P2M5vXwIwAFxYzo7V
y37I5BAokips7pdwdj/wrJElf9914kFJIFs/ANrLFfZMQpgCsnYK8xWxv+Sw
HPQ97yf/IVZCH9An9KlP7fbQvfDojBDw8aV1VfeeL22XEhBSAOFWz3RK2iDv
pX1HLp0ds5mbt+lOJA81pK/+x0RFp4hZNJ2BxDpr+G0lUWsdmM7XtqGYlpBu
+G8/+Y5j07WcuKmrCjH+vQ6Or8xWcJFMb9ILnJJ6LIFYl7pV/SmCvNkcvNOI
AD4GS6zTFuv+mW0o3zjZfcOcxW9GaaLKEW91U5+oZLebhI/ErM7tsH8LqusM
H7/lSs9EI4npu3dyJ6nxOmgXIjM0pUhTvTXOjJMGIBO0+ND13lgVFxA33wHg
6Wc+q+u+Z7YIYagdoCUs9oVIPYikoHCb7v/LrcKs8Sth+/Wkf7ySHtElFQqs
VxvkxHkrFjLwxW7Rp1xJbR9hLUhYV/qZPHAkP6exE8hkQlF3n1iVBRrwTUKZ
PjQVpP4YHi89a1tQz+mb3KhhIr+LTACbpacd95jxSz8Q2cLpWNnDXVfuOefX
qPuXqGRI3OMfC9rxJXWOR13UcTyyN3GQQH5bidSdWjbV+3LthV2gDbBwAVda
HXZClFXCcflrsDYhbQTi3ElNSjQ1TTDhsplHur7im/MRlZvrpCmgt9kNpb35
cwXA/KSF7AkRJOdv6w474TCTs3nASkZWNyo3He37aREUz7Y68b0LOVlYEn+M
5VcuYneKK3DoFSbokR0ohmE6eGjxv6NnFN9mozTyXgfvl05yjsXxoLYNtQ5G
hdcDIRRqdVq0bwwavQQ5QDQFgOO8Lmt+TFjCFz/2zdvjPCJlYuM1KQf4Meoi
rGEHR3ISjILtIDajMWyqi3QEiO3BJrLeO3z+RbTydmwAe30zeBgQUj0RVMvc
QOAepbA6x+1S+xOc+P5S3FmOR14tIP63cRbY5VKLX+QLtMm7+xgkAYDJatPH
CBCC/0UdBgJNIIN/J7c89cluJ4r6WRi1/qqvZkCpHEuCbHw9nmcl7UUQ3Rtv
uVBlvtDUP26pkLsderIjolz3kXDZAKe2A8H1lg4aAwlYJ0bOj0aWcXDGuDvV
81pIuqIrHaTUVoKb9LF0Ua3ZnusvKGqfa54Q0909eZoxTmY6rRsv5tG8SUCb
HA48mfKNii+XBEGYzhsZVhWqyBEgNDfPA1irPAJ07RnoFM1wOSoSopQfreQB
agXZB1qcIaNLFdncV463XW5DSSc92cJVG6bt48caGKeM/Tq8pSqyGUm3JoaJ
4lIVDuYVetgv138hk9WJ2f0nKtulXdM9t+qyRkuud1btAl5yl3eM1BY3FbHE
GtZFHKGqPTZM3wiO+qmZiCZelelMjBSGF63dWQJG+9JidQq/KSxlVA75ryXZ
Mx7YqcCO42U//E1dNYR0in5hOHJvFrvbFZETsYgxOtkczvJNMZtjYYRhk3IB
027J6ZDDTyvpi73msrW8hHFM7PFFPYyXG2W1kxJ/wE2jzsZrJZMh6sj2PjXc
KjSriYSQuoHmr/QRlbVawUCU43xS4PeG0sCYnzYXT4U9FNEuGwjggGpGF8vK
SeUs8td1THY8Fx2DhwnU5DpA1LesMIefwR+8tNvfMWZdRx9uXn8wzjGrox26
n3E3EwBiOM0QPKT7g9TaWUDdnKiHqzSJkAIycXfQBDObv7rrQkdiqQiAN6Uc
pO6HfkPQqriDYIFwqAzJuZcTih7d3WbQUzvR4KX1hfj971pDTJrXrQyVNl0q
MTDpsc3B/evPNZxEglHT2YoTEo8Q2APGPFT28YnSXDhukpsWug4t9Dh0PeJz
89Xlxiz58NafNEYm9KxGQqUhpKMpS3BQCwoJqNG9jmrBkluFORt+RJjF54qs
+/SE5qCMn2n1A/iAldOsOhqGfR8u0DPQKVMty3gAYjt6qWyB7mDm9/9Y2VLW
JrznYettnpIZQK9n4LZcG6kKeeN3xTV+Q4kYWfLuW6XQJ42d1aJ7Rx3A8S/S
tc5y/9btzVh682ckr4Xv9jR+thGkfMBknBU+ZTzQn8/gxl4/gaPbJ8x9p3iB
ruW0pLg/4rkCeSA5BkvNZcvhRBkVY5s2669so+KxikRQWLw3Kaago8rrOf0I
MQy0/xyX0PH7OBVTClKnUCVTkafHue/Is4pOCnq33qmw569M0riDv1ALIIHS
mcZOkDyKJBgRImWEZehDxMljPj+syoBLbRPxojVQKakXFfE99HpPzjRf85yf
62/1d059im1IwNn5hmb83c45FlKv9YVDcprh7GyZ7n0do5dxOvAxVsW3FY/9
TwuIvksSmYd/ndjm4gOBcIyyLRY6Qf0tu7xYlM1Qr8WEG254kl+n+FxqVp+F
YXZBHtu+qgoSdUk7QtuzK2pthxbdngKWqh77Q0RU062pJJTgsvBqpXE7b1p4
2x9Jo7YRtosjg+knUreHfil6DEJHBJzydxhPCxMw6SQ3ZRzcmcg9luU8+lOo
7szfcMwuYYr9kX8uznA2gCyGrdhcpukCh9A2r7ji0GrmkLWHXVi0dwTFxDIT
yjPb3ovWLxGOhKajNQO+U1fsJ5JcGCPVi+UgD2q9194zIo8L8owssngJkLZh
ioTQyfGnczTkg/YhcncVHqmB42E3xqS4RkCQVex9KF/zI8zgKSV+Vi1zb1rq
qpk1Gn90TzthpeUEHX4LX18vkzYO0qghpXUOmp6CyMkm+7FwRHyJY1fniVJ9
OZW/R6ZL2dUGlPAaFLaxDaYNDuItc4EKAnF2WxkEk8s6+pkQ09qN1DL4e5bW
W+CfA0SN8kUiyKjj9N4pJWMt+Ma8HSFRgfFg/FEjkHRxqRYUOMiNcx0/yehM
doXTmtrWR4hWFJwBoLwhzFROG7MEd7wwKxoDasndfGE8gZztuS5KyohN8HuE
4qbtKCDuV0Fl8JmHT+eAZLU7+h7awEXoI3xGRqld8UjfWE6tzkfvkHomFaOw
Y2PCp9BY3Ve3PSDRKXaa64yV67KCCi9DatMHNDvqfFVDR7dSnuJtB8egqrVu
wO8lFhnispptnA9mRX7/trY2HVki2vkEbCWg6uLCNkTJdf+q75A6jW13WIKO
Q6BZ6qVmBoXGZxdYrTELewQ+JRLIjY0HU0oIWdqaj65T6aNHnfoogfsECYtk
Dt6fOOctXRNLykLZmhNsH3fCqfujXX1fq5bo165V/bIIAe4riktNai3p+siw
7bGPalBRktNF5yhiRacGaJwFk2t2X1YLafKFFNLaaoPu+wilSWpuNRatyerO
7ml9kYZu/Q2Q6xe4gt2RUI5jH7O2SXjSE5hmBv7xuBPx47/H8cND+1PBw+Xq
in3w2XMIVYH+piXf8hU3cjfiH+WExIqZmiVNOvxaKSkWxwoNdXIUIHPaTkVF
ZG61q8jhuGu9g2rqBHly2NEiKWoywoSVBqdjxS124LR9U8wmO/V/TCS2OySH
RXrIhvn3s6BsnbKqHta5jNiA18Qf54pWalQtJv4kSvPIBnWvZBWK0VnThZ4u
fL1WECNi0ljkWNYByPQjbcoWKH3Fvy7VgkXE3zkXLzeJiCeC74LzQ81vB8Hi
CHO7cZmlfGMhiHgyuC2UeZX+YzWQQshfQA3PA4gBm7M/VBVt+xhSkvEb5L/k
KA1Ziw3fFC6pLQLuKj2f93Et3i7vJJ5kJ2MprV2345k5K56oujibYGtGgl4Z
1C1uXlVJSQPcDlCl7iwwwayTSyX5BxO8Y+F6mpVgbCQOwrPy7P0NbmQJkeH0
s2n+bRUJhUUuI94B1V9Ni+bPzWCfyleuD585IMT4hxutmZM0G3KvX6ToX+pJ
l/wdDknqhjH0dgx9EhCK6AaovfkLRZHowCTXqgqZXJFFyznVumaAHdRHH+5w
ctEEZ4S/oWVQCF2kjIeYF6e14LH4S7S8Oogo31WQqkAccwenJ2L46KVAy7m2
WGTP2xl6vcWUvQ8EvHIcr8szdzALeyRPQf8kdGyOCi3YVRN9hbTS05yUSiVC
lbgH6WWHwDqf0iM1M/vOYZKFhD+ZOESlZD2CBRhTtCWozpJSE5LHC65vlneM
JZLzOthjx4ZtuTLjN0h/OrMo8QBSzcHxQo579MKDlpUz0at3+KEfgZrOnIT5
OL7tj/ehd0pjPRvzABsObnjz1M7OCHwDMHzBBkCEnT0q4TeMiRoiGuCp+TWM
SLAnmWnYPqeFfkU2WAP42wjkPNmG+cNTxYa6u0lH03bv12EGoVprvy/ZQUYW
0ykCR3IgawKRt8VOfXkb43vyBaMETRe1T1QQOuYQDELL/elwgtTsq8tZKcik
rxdEdOMM19faIHDopVRv+6uKJRUhebl3cDgXAe2IIvwjkVV5ERQ/8RhY+6V0
n5tT7naY3SvwSCKy0/135vhjqXS5zcnVpoyolSjWz5kUwFTsnrc2JCeTWvi4
8gUiAwXFwTWjRZhvq1G35TZt31WIOhXnh7rc7rX9fZyo5mX6Q+07CvkpwwBl
8JwYuWlnVHNv2tngpSK24qriZbzS/YXAFya+dAbMFV8HQIMgN5qznK0O/okb
yETXcriPzL1MvypcP0IH33o3rrFtpiz8gQPag6dZvI6C0vW/S+/zBHZypU0Z
IxZrYfH81EqMmCUkoh7urKtjpOXASvp0Sw7UXs0AsfG5TFZwyGlsclt+TTV6
5KtD/fBjig3dVzffF7bEietUmxJgfC4Gn58QPqO5XfvXqj9zq/JVN36DJ1yf
lQI+1HA8U8ZBA1AoO+pBMk2HVrdYh4jbsEYy4uF5EjU2l0NazsC/b8HE6Oh8
fgzZenifuDlYmsIXpDPG7f7v+m7Ys+chM5zaTnz4AQKdFdkpJNId/6/df8yV
sCYKtOawTu6yHSGNk52jxfTTzj7ds4lNZoqgaiL4VCE93i4gA1jh7c55ZLgq
/m1RdPvVLaV5E9WEC3yI+PVtgC3cGFDrBYkCqZkkNPlGHZNMnSbGoM2gQc31
ge06FzqC6V9Eq5tFRhZZh4nR/7MgoxXdt6vnFVVo3dCd0wltzrsCzUV780Wg
0Rtecqj2pj6Wv9pezyQ6iTtRZI6E+tMWB4pSkV/3NXDZan3y8N6Hsr+sUq+q
VTtk3e5kD6JWO4Zk38wtA4sbB+WATa30iNOWctlEj/AnJ3QUft/oOqbvOVGH
iPNpkT+srudmquJYG3Kkx0djG2kcTsRCGQ1U1drvQ+ha+xH/2dYZDklZtrB3
fzyIwHfhaUw/JW/PRPwAjOPM2/mC0p6aciqZMT7RxJkjGZZEjMmCy8uyx5D0
4ZXuNr/3d0lN2uZ7kFTxLx+IZ82UWtQAHfszkKcI36/5GGuqps6ZCUo4HWsT
pc5MQg2unxzua8kqg5rEbzMwwVAeTXqQOkGy3dneMh2um6apoIxkI3NldSzb
GsPW0KPwsV4F0C/Ec625mD8ndpah8kjkXl7B2SDmm3VnFAG3sa4dl6DbbPMx
LSQRxyKEYdR9VJRnuGl5FKjsfDedLLdXTbnZDuIEhy9BLgrn1PnePoWtUMd7
zRb6GWdv3NhF1/QnQzae7LiH27sYz4F2SgXdUFymI0xeEbwIvR1DdGl5+4Ju
I06W8AYZPiwQ+OsQU9yhXfdlAItyGhCzReEbHbQ2ivpbiPkEB9s+YotKT83G
uA6HMgb13T/NFl5MbszfD38qURdASBu9GC54xJcWq1p0ZQ++ARkgLbVaUozG
CQ3V9erGCm0YPm05Bwf8fXpp3jPn6GvvzmHExVIiodDaGobS1YwVG8/JxGdA
xlQaSY/w3Nu7hv++u7Uu9FdABhYH2luO54/Nb7xf7/bA0mu5xcQ/a1oFl2OB
318qAzQuVBOTLIR+3PtXSRzwhlEAFlvq12pc6smUHL6Nf7vb7X9kODy3SYYj
utL4392YfZwNdFrFIn/29FxWhB+QumGJ+eu228gYvzL8wWHjH6Eo5I5WMlHm
4mdqfkdZi2w5dHONEu8x4WraKtMRi0ISX1+nv6FbrK9ALWhvgjf2UNUEPc4X
E9W4qLohZh3c1R4RYVgaonkMNVq2nB0qrzoBpTAxR26ru7q9Vt/VoYOny09l
A+P9leGxPdkptNiOgbtpqq5SVsfbU4c6hg9u7H9RlaiiGnuR5FEg0raRx3sR
HpmX8Q8cpZ5Ss1AP5xNkS5fmI06Sk6TXvp7pNj9dkchsvaS8VQx7i4O0PIxm
v1oN2OsfsOi+cHDRDnTaa+zsrDwtBWUjENpzhwC6XNHgojdOOjGx9jTpyZmW
lkpeHvXkbZU7/8iW4GKBzreEKn8VS49kIkEDcsKNMzDRR2Qm6QrUkKYTMhiQ
Uoq8Gfa4xqXxiPu8YusWDH0hIZOw3FZFPc2aTHqWiU3a88I+37oH4mvGbkb7
2/46ZuGpe+cOQXPV1fu68bADwVhlAny/ODWU9TNxbtopEQN6mf890Xhmtk6X
tftRq5eH20eYYPdiA4hCpd+ORNOiuRNEhwQDyWoyBor5hBA0zPWwbEifFFQP
J3UkGHFLt0UwakPiWjkMbu9oux1/mfDJnauw4dz2oMr7L0WfW8wrPjJVd9B2
DFm5H/IpJS6vWlLFtqQKgLEqU9rCpwJ8TFDV1NRXpjIq3iLZ4iU1SYlEycR9
va3YzHfkqcxSrq6vYUoiVbFOwMYlslnHaoU4Hyw//h6gaaHhVJYMV4DJh2JK
XxmH1GcRliyWRIdHc3WJ5gJkJSYW1bYOcdNlDvN+haBgFir2zWzTnnD/lHh1
sU+AEOQSy6VBb5baVZ+FPmgOppwv2RcgNO1rz4kX1TUBAm6kcKtCTK8udY+3
TU5CeCL2v/gMAItowHzmHfYXVM4ADux6dlbpu8OkQPLORcU5ZWTtcLulWq5A
tY8cOn04r9kML9v/E4T/bRd3TYqXE2fEWzMWV4vdC+3qMnMwL3CS+duiuaAO
ovBMJG3ki37FNwp0b30XfC75jBFfKj6VVeItWIe2F94vUm+PsWynw1LAn5FR
BJn8QHfqAcZhqSWJaEc8owhrsYsoKT7faDO8GNq3TTH04VDGj/ejFSpXew9p
O+JgmRgGR11HnVgaWR9ygjDXiQRjiDDTfq48iyoTtaI9GXFJvhkytfCuWMw5
TRF63uFJ7HYynBeiFhp2XyqvQAqDdgo3+7pdbaKl7aLKCdTAxjnt920+mle9
gDXqkulo5WbXWhuaPTY2kzuJuBX6uI9SSRSfkFjZulu7TN3J2ypZA6bv4Ak7
giGDZ0RfuYMsugSFtPuH+H69OKbrI1zNUiMZ/tJkAqIY7pTl7Lq1u/q1MV76
c2T921rMd9guMunrhMuOZuU/ye5829L849Vww7WRBAWQ27J3IiJ/gDFf9co5
I5OQgX7kelqRAZRc0UEZ8o5/bGeB7im1x4b9s1wAJkJqKFXWqTVFxj2m5b+z
htyJFFUs9XhmvfgnKz7RdNbe6TuWnDC5dSyvM7FgLHhpXz4ZZWfdoOYlfZF2
/y9jBv1Yh3CLWNmKcfLnP2tzS/qjbSyi62iN+4RT6K6IRQkZZRqXAmhXAZlP
he5t9zOKlvd/2lw96kJJJHMIjVFxgnOmP8XhVxPUlIy0azW052Tcx86O6/nc
ZUzTC5xHCiagdII1gj04plhaOax07N57f+PuWXAlTII1FQmVm7BvtwRZ5mxT
qjs7gvVhSXxCytJ5Lxlcts6NVKtDU04JOFxhn094Xc/A7EFtUrbpB6mv6k4B
6ZNo5SkX2220EyCyCYCJaMfG+YFv/zlN+vOSA21VmJLIXacx2eQLBN393BK+
RbRF2NNRSfGjglaPW8ECYldpDHeiRcsjyHfoIpDTTHx5uUPuO266K1qVYjHZ
zoe3IXerDmf4iYAbjlbrHDsQfBeMbfADFPxgwyOfHdYLRSecti1UdJ7WwYeN
XMwlDBmwW1FzIO0JhFDF8kvtJ5/PvbTz4emvZUD2bP+N/Mj8XWbCBngKmSON
qRBhnEGj1pPnilGDwdyGFCm8G+7nrDMTp+rsmHByIsexliXPZPp+g3l+8etE
xemK/ximn3ZA5dJCdo0B4jB8RQ/R8SXdD8CUfbi8vKjdPU7AC7YrAxnpu6Sj
QAyFO8uhZyTqFgSiwVMVQ0lS3j9qC7QyuNILqNYVxv4isZf4yNbtwG0NZXnK
NZ4suhLHimX6iQ1dWAlvKwrYVmvxVUEPyOk+jVCBDcekkE7D6Ji/d3+zEWH5
mSnHR8KojEvM8LHgDTVkHGRWSWijMJPOhYdMq9egDXYoPEElXr20LvS96Q/A
j/Wa4//uHnyY3FTogaZkg6y3gKOSCiN2vhGvlgk7HnluyUhwQB8w7f+vcoI/
p/jkOhwTpH+cC4TUwJjeK6V4ahBO0oIEX3p7XnehSFoLt4T7dNdmrcgVhKYx
K7aGrR8if7/jteoEGClBfpQvR2jZos/P1OCTCI7aKIlYSjngyRWzhBMxFRVu
i5zy2IIqhD8/wW8EwgIsL3hFaxhkDjUvL+Cv9RA/V1wtfnFwhzfnL28W7YN5
ETPwa2Y9E2cjOZj6CtCrvBJcPondsWQu4gb97Jdd6GpY978G08l6wvjgIrGc
ezW83HiPQqtOKrAFUNzAhmWYTCYEiet9Uc7KOLjA+xnN9rQ8amI6sq0XURG5
ZD2CKge22zCIdfIDocd+udjYyGPtJec4k1suGUyW2pzDlI/mUydykAcuu6y/
WCfoOyYa1BbR1A5SDvVkHz7j6B8CHHo8MqSUj/olHDRnKwjd1SFdH5TNdkO+
2FKAW85JVcsyfFJ8/ZYAkbLQQi5R/3wnfk+x6V2YCMUeRVacPNbljeS2arKB
CNNv+KnOHWr6gvyxKeAmhCIF4XyjczhDmkcLI/P/FFv0I9M5QfYSGn+5EY3B
CTZv/cnt/5DlQhJkJtZ+bIUjT9Jf0LYWFHr0LEnfGnVQY4KChsKjQ4JyRWS9
wfBxst9HqINQCOaIgJFWsZ/LYKK+BkkPzwJ9Y4b80EuxkNaH5Y1xASyv6KT9
KRQP68mD3QGcb7lZgDfXgRYfnULukkIT0MLKfMmfsiGCCSvcj88jJGU7utEA
8vxSdjcuLql0eADphvkHwbgSWY6TnfhqT5RAmSAOzjXOVUCnerEDWmlihBaP
kb01gEdWK7pqc7UhvIlcxb7AZl5t+KGrE3VzzMlb7f7UAZ+XtdxA9GaN/O9e
QMoerfare/Kvgxs4g12rwmYH6nwjIghdTIpc9sl5Jl90w79cR4kTQ7z/SgqP
yR+tl1HLKj/qn/7M5pT+r7Ihg5HTr7uxauPuhW5x41vuKiBkmWduW4fwYwp1
8C9+TMVOUanhc8RQVAzLMfIzikvLMhz49NtQSsUmymRV3vkDj98lagrigeLK
yrDyWoF1IqnOSd+kG/dSScYpmfLO6/OOggvz4/jR2FT+4sgBpcJscTgR6Mg4
PEl8rqycQhZvgOgluSwOevc7BplJKYqpa24z6I6X8y+OAOMRUSgoafh0d/9r
Ho+cjNbG7oitaUUvCwAgz+nUNZnoxStU9h81gbpWHhnhxwRxxV8xCDEcl6Wc
ljZkQ6ht70qwvDdHmXZGBp28DNjZIo7uRAeuthdFAjMG772hu5g6hH90dbA0
B7yrqa5LfrRTKaW+eesjoCFbYWKL2pfPDLxrjnw9Ji9Ap7KohHrcq2Yt1Vg7
2S4/crFHTbRpT++PobnnwFaFWEdseeMSBX5jIoRU4xq8Ag3JKTzcTkKzI8vQ
hpj5K1sl5qa63aLlU1v3XDaEIao0G1eKV99X3xuV2jNq8v2fHy570jDlKin2
2UzwjUK2l1n4eB8MiyG+HnK3XgDtzGgckAeDwBil1vnYZNd8CdR2aWY2BxdH
j2gnuM880IMysi+paFypEp7FA6lpTYLbAdbZQcqx4ZRpqh1sLQwvtMxZpTbX
YzF0QG09EmPbqaiNpUuftjH/r0+TUUweIqLCozcUL26Ffi1RhJfxTx40UViu
a/jEHV2NW+adbcVOk3rJ59ZNCvNP0NO4yui4IClePz7UoXv9bD5ST2ULnQhL
GH5TbaIRjQpDjQd6cQkTLrobDqPWDSVnRdWuk/StTgykpz7qGp7+QNqDQaBS
O9q0l6reHBwupeF1RIdEbAlNd62t4Egz8y6Q7WLuuS0hh7mN2gi9ejqHkjY9
M8+bLBNXv2XF1W+AqocO/39rzEVTJGzq0iQWICB5vNiPKx2N6HCnCRPUlwK9
G1peH0LNCjetCe0aSiS3fv2aCjJBp/HqE8HrvvnjGseobcuYn4sIaYhEbxpf
IZxPNSSBPYccr5OVBUqsi6xSCmnKf/XR5ikp9plD700hLaM2CrUqUqd3hs2B
9f3oak7SEH4EFHrq8OOMqgYFB9XzYUPTULSZwa4cdR7VBT5e2jRhd17laXDY
ADqpNetMYZlyPK4C1ywK7E75YgengmZlQtFEZVkF3V88rxslVldtsZI1ECgz
fKA32lTyxr0Ql/ZEEBAxJaAXAiSKT7ObXwXVc5IWQs0L/xmuCYNR+W6yfAqS
PhM8i1J0q6qQyoz38ss93Bd/ghtJcD64V3UenSoyN7zc9L10fGq5X9U31lmR
vt8avAIXNiU7/PEd+OEHNNHYgVXtKAk8hTZ3L2wsCV7DiD+G8QHktFaltrGz
/1IH9dgabM/91iPR/+oEa7hL92AeGKro3/eE40GscSK6swCB6eUfKv1XdG9/
fPyZJE+flQBIl9ioAKV7e6MkP3gtP8ZAzwLfrPXTOfLjvYTrOUCDIT6p39nP
yfgVya9UOCQ1PQ2YzcSlw53Fm4QNjaNeawxFlwHuneFVnNF1GkgYAhNlHRRM
OA/KZZrlh9Ox8yx6Cl28tgVyCVz1b7BeOjaZ4k2p4weTes6bNvK7aO27nVJS
gAJPSWqQaiBJnG0wTU+fRytg7PElclBi2ml/aEZszDLvl+q6GubtTDSAvnNO
rvnkVN0tQI4pd++k7ywqPL796oDECX6gLDkUM98gthVV3ybRfhSmunADs6Q3
zDXXqlI2nCA/SJ8tzHYtRh2lU4S5iDgujCbJ8NVRPdFDnHUo7dQ4cir5JgDZ
0Q+iQz9uk7hHPyZb+Gbnq7MRyRCWZQecJ872BkAMe9ozI75Pc20hI3T36PvC
ehq6r0/+qzW/2YR8zq5GmmtYJxDOPN4rmQwoGLMNB+kHEnE88RWZH0/0Hdkb
+A3sHfPw8sFRy9bssnj4eq65RXNM/CQxSxdQ5Xp66YZMxtGZ55f9n5KvPRkn
OSZgtPnpM+D2onm8FqzsyAQgs21gadPx/3WQwyqVQUR0/SmVRhorg/FmaXM+
/eR1rCJuUORn7EDxHjFRJoet1vUr3+5Rg8hvB5B6wHSczukwBCClyOnfvM5U
RPGciDSXi8wi7e0g6sNIIFxOjjH3dxIfy/EGqvV24N1XYbQlWqZdHoDgJntz
dhZ3wdmuIAe93vx3b0LR1l6BqS38mHYWtjpNr/TPrhayIklrjQh24mq3+kkG
hDa/jJ6d/IEZT4FP4nq6a+KtNVdlikr8VIFtLgR8hoYEFofNxF0KFpxqqShL
AV3Q+S9hnvn1iQHPm3coyF5vW7phBJXKkdVkVwiU6oAIvJ9wHr9W1uCfNc4x
ie63P4yuEeSuPyOofYeKwn/wJIy7hV2bJSOTfVB7wS0Bq7JYHrV0cnVam3PC
kDiGnHT9lVlJCiMP2yX1Om1aJ3rVjqlXAMUBPARsgE21MyPJ+R1aVJlUpmTd
vaOG6Dkkqa1irks7/2ZVx7PN/PDNFDSwFcObBonyApIqwo4WjKnn9mVIyfH5
OdO8V4DUUa3cvMmGn/Y06S+goAEGtGSmcsi3f4VJ1jWe79BbvI8fj43u82P4
ttxG4ClobUo/mnoDWLnXyt8Sv/KKckRSfK8z+J4nGuKFLC9nXP3JjwckvOzf
xRMsRSTvy1aU9X5Xm7oH3K4FC9bF0p3I9guBFsq1oOdYZvmnBb2gZpwlrSYi
ykqPDzKitklmDOzUsGVZmorUt+BPbOEVU99QmIhDxEIZHL/2NF4nulKIzIVx
5WQQDlGvkmAkiETsZMO9JZfPuwbtqQRqInrqoHFewhz3rthahUI8Mm9ONjDn
z+cjEPfYXDyjR0I5RSK8Lmc40yGQiuuY4rG7r5S67nPmetcqLz2n/qiwiXjX
WzwjtLDkMgQZ8KpcOkUO/3QRKFAvIhkOp2dGOtHgbAde8GpsrVzMX8at1wN0
Jv1C+fkfrhVg9c9wTM6KiK/4kQfA3HRAhykgNLb+2XDaS/HvKmUnZVk4je9k
8krxxfkh9sipErDymiLwfUd7rJZ5sciP5MN0kOMNMRn0c07Y2zfyHjzcjiOS
rJnBpfnjcMQDsrdFVfTeN164EaF22xp1k3jOYEbbjvpSo1bPTDQ8XW1hVEt6
KenFYRM8bW7yFJZwrAqCciYrb/h3VdSJJpCr0xAFUSDo1wbM/Pe1NOB7kS1f
IYsS5zdqKD1zDPtLo7DRCWRQEjDtQQj/uIRxTdxHr0DcUpnwkKL9sB+SkxWM
wvj4M9i/z2jTl2BR5tDhH30IKTNVdDFEEta6OK/aCFI9vyI9PLDRurBCHkrs
UllW3EF/rlGhLcSj96iva8/gCWW6vGwxvyh0b6XK96HOopAoEp0cjtwm+PBj
fIUEPFdh3/8Lmvh1HqrTye5zUC5NJAMTrTrcncXMZwLEVo5Iq3x7qAxgdKs/
FGtHOCvPWDW05Lvp/c2D8Ig1YwrH4TfNRpxFscoHJT3vvIrdDOwOnzsMuNPc
skRKplRhsBb9Kn+1kAF8H04qOtrPgg7ydm6Pk61wquIptpw6ZLBP95zxQAvE
leSxqw24+Wn0FyaNeE70I79AwIMN01ZCAxDyjrgwCPdyw14TsWBEqYFumXXI
Pra9beMn2LtPfLUb7ZC3sjtku+BuFc2ZpjYvqsRvJEfkQIQq1kcaEfPBJ1e6
9FpiQbogvrk1YDcrXkENLHXW3HQz7yYdBC9TsF1X7zLrFziR3ysSKXTx3DWO
upwCJdZIPJIG1tWqAVCinTIwAMNo0eUtl1ByPwyFTNXGQHbZLAHG5ZS2q3y0
cX6mSUQe7hu67TcVMUsh0k345/wOiCv6tk3V6BwYLO/aY9GlgjOIZc+tCdEv
A4ZEBm9huzpwBnvrBmCuzPOrtKOQmxKW3CHDOLkh3kzaSKyoa2wj3O7MBzvB
PwqmFzUVj+Muj+6kEON/TeLZAd2GU2RFxS7TijkMtCRzV6i0phqe00yBcQ10
EnTUL1Gp/PghAaqljnUzuQYrjzpOcDe46C0jEQV1z/HgDiZ/z5G6ZsPRqqx7
1e1TRtptEO6OqOpGMbi55Vnc0nfgT1ESizAZ13UKHRXmdWM8nkTGySw1yVVT
udrz/EYylwNhD0wFjinkmMLk+4fSfqgOtrLbOlGd97cOJdch+gq4x2cJeNaL
bqrlOkJ/ieip0J3LxP+WGBliMqDKzx6EgeBMUSlIDFev4/jZ/xfpDseTHf9h
PhA2uTh7wak7fp2DtrIzqXfDt/RqdmSycY3yw+O7c1DNpMMXlsRYux+mAQCC
uvQy1D5CWRptTHP6YEMciZz2hSogf7oKEDjM8tr2b9gwJnya0CjXEBR6yDn2
qrv45rsi11OigUC8XjMsHG33fonHW1EVCoabpMuz/kCsFweUB7izk8NJ+34P
oS2GZ7vtVVJVi18Y/3+cqIE6o+9B9Snkl+N7F0HwE+BH4F3gJfQS/4SWUdG/
OeXPH0TR626lYIKMMo5+NZrFayMSUTRfH37Lcd1ImawmHUAAdHjngnrBzxCI
begqS/zXuoX+rSUZpstwCYapIZRVyPcO04BwJi4q+Lp57h4bK6uhBDtJcB3i
+DAPW1d0qYxElTKDVeIDkHHg32Gcfj1zqHWqj0QgcCkgYIUEmWld7f8N+a+0
FeqK7zfK1MXT8QABuYMjNGa6dJOQywz+d5jHOqaeROpWAIu4eqs7YAOUC1Kn
kfbC8zpvwRSOGT+O5OONXKTRBbJlS84Eu/KNk2mJ4lbHaQFMIXneFP/2RwfN
oDRzBqmu/HgpBy90lFbeQdfA79WHXKJNUnCEtrJSLQ9ITyf/Jha0agzjb8Y+
FNwM3iN9O7BW4R3J5Aq0lHGslT2WgRL2LpEc9PgYV96HJs8MkJR3FUr10j3C
fzZa8PuV50NOxnFQgnCpVn9SuUMm7l+iJ/ncWCBktxVR0iUb7GZ0HPxcg5AZ
ZwJdvK+zGB7YD1KO38JTEumAf4Nv+MCrGJyRYzJIjLsOP3sjzaPRCgXG2R22
auj8cLG9rtB5upcZ46QKnlTirgHQYbtQt1jR8rd0jh4vz4KwOuMDqlCg7G1X
5LpVC1De4jtyWUSN6rN806+2qCY0ofNisG/XWR3mRUtRRQS2feXkiNJMMjDi
C6Erout+fqKyXts/YNdc/YiiVp1IOnwsP4Zm2Q009RnJPhlgBYWLU4cdP3Q4
jaXinM3PIndc+SDtVTLh7TUnVVHhUXxLZc3ltaVKqthqOvkLvg2ypKRkLiin
OS4kYzG8oPkycu7L2qxD7P0vqZBaNObFsVCGoOe8VBp6hoT4LdHj2fhCagEr
plo5yPr4oDkrlhQMVZJLSa4MFkg3RPvKyPaiaVOHTec1RZzoqyEn1DLLw1wj
BZJ1JrcwboKqtwUk8gRGYkk4UQh97bFqqxpQ07Hrihm0dfzpg/QCNiWXPqdy
Os/vBtnPAjEwx5R6qMBi810fjVxETfLly06f+/0RHmLQaoZXNqMzzjxVNoRg
nCM+gK3OgOTcLcokQnVL8m6HGktPRDdspMgu1xndbBa1W02nbw6YZmaGUP8J
ul5Cmmy4KCjcjNtOllUuE9QNrvp9EUqvre5l+unDymgswTpK7zY24Ownce/z
bhAJNL+To7QF0n8vKWqjziw4I592FzlIc1fCSD2lGj7HV0Gn54zQR9jNJpsK
3SmLVLWTpu1kE2n/Gzt+rA5W3mW5ji8n04ErpEKb8mPvWDKT5Zdx2UVVZ0l+
isZmE7UFWnZ8Zc9iBj53HxrxgSFwIuRU6D5011Ppfv0ukIn7wwfd4rMgiEu4
ztMZmX0cH/WJsxYYnTuFsrfi4wo8gol78sLz0lfBFq+RAQ6TMGSaUbiefCWI
3o186tNfYbcsi2VoOdFXJNigh4/qkxaANpozuwfxCmKHVfp5RttXuoGbLA9E
tRKEO8qkcpKg8fJUSwbiekX4ufIB/6iWXwMKvE0bAex+jTMCM5ztvI3iDbGi
NhLQui9lltCMuVZhuVWyix+KnMCvVr81SMNu5ceT5TpVqiTV8lCUpSDyB0tn
uZwruMptgqYr7Tv3meaf6U0HLpH/QpQ0rm75V6ootiZX9rEjBVD7idv+gBoJ
ukpRqNXzDAe2SipveNR5rqFra+UA1u1WajQYNYjeHCyhg2V0Aa0VYmsoc663
0PMdakKCuLxMNA4FxWwylF4+mK9u0KKn0F05BsXORRkRwjYADHruiy2nvV8F
xiE6wjUP1Qr03C+tA7aZ3KsICc07wBq8vSK5gjg5DEGtuS8B5jvk0MZkudLt
3eJbqkOVPa0mVQtHePgM7hCKkvZVFo/R8OUMekzFl0rVQINSuE6+vW8hBZVm
mvNwAvK+sUFCv/idYCvfBt/Bg4vhSuUaMUExHQm4E8ty/eUUOpN0C1K5qrZY
NGpvnQccs8aLiXRGlGfYoJP2Qkv6Qo0WjSEYmdAb/d6vVSFwG4/8JUM4Pmn3
AVyyWroQCwJsO/gpgxY/ixRU/MieoHBV0hnzl8cCNYGBz8jmvyGM9H0/BlBP
R8OFl4PnVY9tqF42YjeAXO4YbHdWcZ7ViFvyEnsj5GP4e5ovUzMio7je9sV7
Eczc3vEDDFXbsoGh8gYpNeBtawHNM0bqlU7aDWWq0oxwFDDdsnlP97LbxglO
NM9zHSbkeQxfnDKd6BPvUroXLHseBWMqOO1ZH3yyIcSBQ3MJyoDmYrq+QtQk
TSgPzCQ0yja6089kMynWbH43jAmgvcSYopziwEtd/zIZXVRRC8kI6G81QCcG
JdQcvxCSir6FVZ7eP4kZEE1VXdyMG+xzpGWJE5eukJnWaQXs+S2e1VdXzJxw
TEDxU5pKqjc7ktfesDJ4wtlS4SmI1B4m74zrOkS3FRXdXpz0na4V/6kVdVGk
xHhr243e5FANPp7y9+J9ilOpfGyxjFyUEdYuSoQDPQfCVtvCADTvyqGUuSLR
bqjr9Jc9y7iAzN79pu4wSxx9CIJcyFu62TPdW4jhkT+rmDnzwGcXzSR5NmL7
N4GS/UMyv9ayQ+7MQeOErunQipV71D3dcrtN3/v456Zc2toHZgFrw0GCuiKz
KmN7rX8r8febMf97whC/svagMSM6yLmKO6Iu9x5UAArGv4wWmEdhNw6M2wB9
gVnZtJdVyB/6ABugM6f6AcPITjoKXtOIwjrOX+u1VLcPf4ZjOij5WC3BKhOK
hEGYk1f8bRY1bc2jbmbyRebIG8l5IxTecZtQWiouPDFWVagAFBdKDun4Lniz
72yZY/13cp8PhfKBWqGlbw6NB0t9L+8GT2m/wmnRlxJnbgWyZoeVnkGS2rEr
M9uMfPo/BYpzVPFaT+kmYaf9k3ael4SEdXuUY9qpebxkorCNa89fU86Wbq0t
iEMoqXl01Pd5Xiz0jgtbQNhmAgneQ7PcChKWm7TfKyZ5+1Qdw4nBo+FI80lA
AScg/hqpI2wdXMs4Tp4UJeZIm/PaOyM9W9WP88UaRw3HeGzXcA6+w2LITn4Z
xASqalaXhdxBJiBvePZh8sb7x9wdKj7iK3cbziWU/plfW/QR5SW9crbPjlZw
KZaliWeEkLWxmH7VmABMD6gYaMfkC1ACPo0Tl8o30kstX9nfrkNzzXiDXGU+
cmjtC9dGjc16t69IAj2d10876a03e2Q9RIg/eCuTSNIAwY2Nm33kkBEKZ01H
lsp2Kqjahmu29f5UMoxt9pmrkCD0qb8R9W06s4WhyH8E3/MYuqQpIiIosLRS
12rOiZTMSr88xq+y2mqLSdh0ZRPSwVedypm6D4ouckkQLG+ZOZBmixPGgWSh
3P8O+KHvg5YWHf6l4dCI3/cHfK3T07onkoZpzaptayjeBOt9VqnTcPMJjzGh
OYTow6Njr2HgStbgVZLvKE7qIwAU7xYUL2uQF/jghURBRyTnbuoWph0EGuJG
MZHfQqrL4DpUPh2lM4XJJkvdxp8QBPKofAxG069c4odykSlDb/4RobQFSMgi
8X0jmOGERVZDBCRL346js1J+cNrW4PIfBGBspEVbsK7H84UJwL51OZAr1JSz
ZirFVmhASw9Wv7sHZ+2SrxiXnKOZ5AJ+WrTSbJ0/Z/4KzAbE82DVdqTD0k4S
7qTF/h75O154CV9SZRxVKjJXoVmXnZQYXrceGnjdpCY45abOI0x9ihn+iw4G
ytrvP0QW4dSrmiDmtDAAWDPDpYIcjz408VvxOmxjX1VfZf63gmGk04IU8crw
4CnA7qYYvPTyCSJgkddxq/3eYASHIoY/IuK1R4FJEVUZZVMxmEhDeKq6+xsf
fqoVVfWDepLgbv4fh1GpHAZRKwi7RRNTslbHmFetKnsMXuoMZ1va/VIuNbq+
mN8o/KftbaO8j6BjEDm+dsGbGCN8qOn9n5QM9z44X5UW5F6KUHYnj02NkdaM
fTK7GzTd4KOA9Sx4E9Owpq/Z0UoYm1K9M/T4c2+hTEfT2PMQgTzmfmjM7cfK
XddQh10OySypHGHQUanHiHUZi1ZHT914mm/rv/a/bn2gJExZyHo9bYgXf0iT
mu1qm8UQU1BZR+sSRF/etvyOl8X7c3PLGjPapUnV6mu0TfpbA1W87CmQor2c
L/EsCTtUVagQNdtnhaNCMAgiwqfejsIhYNaU5qNCSFLeH1W2iJ1/dac699Hh
aMFWFv9FPI/ow+7ik2vUfMlId5sAdgv3IEoGnqOWevnD9yFYn1FuAX0jziR/
SCAeP59ZQ6+NCixK2MyzY99SZCfHXboqpcL72FrVVOkEJRWO1n5dDOujOCV4
ycvutpNVm7qMz6JR2snR79jpM3cI6aqqYUY8iwD1vRE+V4KISGdcR9eGwbMd
IL4JAYsKLMeToyOX61WjZPDI10AbOhbLGjOjDt+LXkEM2NF5Mw2Zav6oHrYF
1RJ4fhNdAgv+ONKYft0DukTkAs8ODw3DBgsf7xt0a0kHtTQO29iqZ2W3meam
CJ+6+uvasD7uYoOfcejcFVtW95GQzF/qye2NwcS9ez7kUOXXAli5ROBlgqmR
TebVNuq4KK/4eCPkcNzwcL4p2lOA8TpfgLEj+OGlT9KYrdc/6lwf4qo93XSr
e7mPdNI8clIBELC9/a5wxW1jbI8QyROxB3G9MKAdZChegmTQyVzDcE6ufCYq
bH0KXMK+kbRA4LPqDlu8e3QBoxbUVuZTmuIcQ/s4XomHkXoWhk/cwpyRIYm9
VtvwVFZ2VN3q2rkxPsPylk1uyBS0jIpcFZQ4WHu+yZFfM6CcxK/ETrhUystZ
ACZCVdoWt9MJdl9A9731ic9bxaEpycgSr8kFq3XwyWpXhVAeRa3umweBgRt3
RiaEITxXUOsRiHSHCmJPuSEJUfHylVc/jIAars3nbJiVkmkHQZbXeEDwZyvd
Q0ysQAl+cxee7NU2xxEfss64SCUxsH1PO2dwte64xG5ja7hmbFFrX71l7rDK
UeYEvjU+6Nig5Ccd47fCXwaJang+sJY6/R+TVdYv1GWpmJAonCsG8Mu+wP6Y
MhKoC51cWHB9arWgGffEt4S3fzGflbgN2tytfsRLgt9h/LJquz2KdfGvPKVJ
IIXw0Oaq7hWIDyBcZdnQdQoRHImFE17GN40Ys9hthlnbFH3dkl1l/iMIsj/B
/IWeMYY5yunnkr0oo9WQcANbJemgLIpjKV9uipkoOU3g1UoTdRKTwVLMD6uB
0HxP9BlFH0UZxfLIdMSSpNtDFs+YsUEBskI8rdvl0Wj4URaXyh+kHNkttZU+
D6SCwqcHFYw9lfS2AWIS4AWs31gn0d7Us1JD8N9+LqLSMT73wQa8HLKog7f0
kiYJBNPR2v+NaPVhW2ppJ8LH0wVRW7IL1Ly4F30Luhm68AX8ITI+L8iuiGvm
y0XQuSZrXL3qeinXNpDwnwpLUS89pitrFeQBnApzQdY/slQbjydU+LBqr7So
8YAwse5jVAWkkgD/p5A02/GLqefL4Bu2+cIKzNsvb5fN1+zYf2FIP+AbmpQR
8gCHzRB8+CMM1lcbb6Q1UW0yeTtVI6pZZ/B49jU0e3NPFOEeyd9b97KMVhEw
+Ge/ZjDuR9rqDwwtKTWbpCP8VHtoesUP8TwdoSj5g/cHhOUSbdgjCc+4f5+0
X0nnb5u6vFTUdmCBJlBGkZoSydTU34xNWNcYZHEj2ubyEOj3HfJBxOzW2xAt
49/PyvX09HfqJRyVQSYsm3vJIhTVhaBcY/0vFY48+UneJRHjDi0la04wohHu
azkuuM3ILLHZU4eMTrhGBEe4aFgIivGb7G15CwYLrOXbKDYc119astNQznqN
+psr2/G5P8mKLQZM4/IlR02RQuimg+0u8G+6iv7Jghs8tvYxDgwInapznKen
wYdIyfmNXghEYzinXDRLmdMfWDsv4lHVl7RGHw5su6LGQC5XQ9KKyipWK0Uw
ebisOOyX5oVDuBZt5tobROXGgd/GHJHaIGsvxj/RFyEb/dUBT9rKzqkmKIdd
GOmpmabZN2AEnU/0aKUc2uMMSuPo0u6IkxTKD8CYfajuKYZOEiYqIYSD9HlT
Q571m7PuZ/AdFmSoOZjcuu8AcMVx7x1XvOg4QRVHWHIG048NTT/R3HvTKW3g
OptUAnJneP3nyn/Eu6V3HaY/hISv4kwiQmptvQyRFuI89GmbOPp6/3cbNTpC
zZcsy2L7LKNdddHzftjVB49VHhARr6arNC8Je39fkgDRAxebbPx61Uzh9+Yt
ds8N3EOwx0PuUZh1/hxWxQ21j6QEmG1/H/PGVOTQk1zYHciOIC9xAztKSYXC
qWddcCtzSsZnJe/n3lQJfxPJVt7gv3C8eXEZxXIbyxDhNKd9689NjAU28clU
BgHQUqeVE10//yPc3nMJMyD/TsOSl/14N56nyYVq+G1XpvPZhszzunxDxTQf
NiAeXbsUSldr+4P0HSDXxpE09UYyAG1ugdpgGOVhdi67Vx+NtOUwlfDgpaGD
l7c5DcY2gCU044zBZDllbPPOSOi8+V3AKsz2p3UAkOYnrS9832ROXr4XnOuY
383ytq7JADrFBIJYTBA1plbL0V6uAgkmD23udfrXo+TFbLI/TPZYnrGDq/nX
TWljqnAp8ktZqglOlHZLR2PNAiovkNFCAp46Xs/SJYGHeI/MRlDwlw4MAg73
qj52uo4CgJ3C0ydqClkAx/tK77XEskzgnY++vbc8qzneHznQYoQeDXVFP1U3
ymvsBLtrsetthS/wRr0fTmntSB+s/7OVGK1azNFXJXC5MtLZQIWjkmLnAH0y
xXvAMvyVsgS9DSU5szOPo9hjBF2QYrh0k4UDFku4T+eRFASX+OgRzh2JLf8s
zjQcCAryu9XWwk1MgXV86fwIpwtWmY3oiD9XLelQoTqScj4ZshHFeHps78sB
eI3OAhVxGooi0LRSNFdVmzigHSC1mJm71OifcC85RQ/EvVfMI4OpBTZFj2B4
rns3qvWNPOspMwJi4ta5W+TJw9Z6OoDeqFIttNA4QZ3fJHGGnuBSljtY2kxM
cxZQZjDwiMaZ0TUvEW2Ve+AabpOh0+5fKbBMlsZIgGbV841alQBI1GRXyu/5
ZKsABoLOAC+6Hh8YnRZO+CcynSDy0OwiFedM8WIjpIx6LmpIlUNGC3soKEya
IrAxUuySO1RLP2b/r+1uRuyRPlIBIUU9P0WkJDMmYezk9W52VyzRAJkz+1FD
fH28/0sKIphTseMBII0Rf0TtvsQVeU7MsIT4ze4RTGk4KiVd0heVMVeT4vgN
LcEvifVS46s4mv6qY0ur/Cod/GQ/QZYqm5gxuLIVFKRuWpCHcWAjk4pfnZg7
1N6iPPFMdZb84YgsE++ujArK6fPDnTpLvzQLeT3hnuXc7jUwwO8e2UMywan2
vzc4dVm+kiFrdN0ZzSLcAXEJwasWd36tigNa+/cFAM6s/LSIaf6v1xaPVQV+
OB73jGh/0K+udTIIiQBmqIVOxh2k5sXGMO+NsKR1eRi1j33jIfS4yQi9lTn4
5dK1izbg/dwgzljMo0d9eQhreZyb/O6s/CQIeqKXJcTplDUOF7t88ntLGQU7
oJqcGplUHvwDDyMh4KhpxIZNVyYg4rlFuQ4DUeH9GOqkdTF5CEO8qaZRfZ/9
eHHLB2jmpgueLGe2/MdypyFcY7NyrFthYW1TbTPYXP45OcPJqm8aqHfE7JUn
sx36nxHXNJ0nmYrLg1f3ChdztLAY8tEzlG5dedHNknfbDQsFe9d2+ntrrdXq
zt3djUOUKm3Euz9gJ5PCVPsAa4GaPh+CrUNKnVem+BOT+YCZACTwBqlcsFR0
TjK1hsEIlFlptCKy3mUCQTUDMvDeAzMHFzAFIq3oTmNBYeHTp9faWNOAw4e/
Pa8XwCE7GhD0EwrH3D00cLvumXkkrtUTQx14lRdJgo6X2Akg+jKvF6skrytN
EgE8PP+ZAvKtm9HKNnRIWuEvn0q0THNkER7oRMabD/TbMxoB8Gxkd6vNySsh
I+6guTbRDokv/0lyHkof349Ezq2kjwc/C73tlWzYrc5vMoEWG05ZzW+1lB3m
7NAic/XTyKEs2y8LCNh6thYfaYMr+YpJ2+rzZ2enQ29SFtj6nBr1LTVJ8ARo
NmZAu7cFVfO8lY9oeevmcHWr7zgMaoo/hyAi6VJjAvGoRJDXhOsUdIdqX9nL
JENzMHR5QzzJVHRqgYJ3qNej+OlRjZwQhag4QZka5qzhi2awHQ9rCg+IsD8z
GL4Fi2Xn64DEwM71KBVUoD0ydAdrJ4OFhrGYi8PDJo6l70SoWCZiZelFiebh
3cX/fO00nmR5V0lXxDkm1yhipc2IXcTT0fo6jR/ODdXC+z2g4HUVuKt9uX6g
L/FGMQ1gBbjvLbH4crWi4+zwEOYlznNMZ/hLYVBINtD4SA1MJjNb9S/zvxq2
xS8iibjY2sYiIdHbT3x6kGZZW/UwR5JqnnDSdam/W0AmbDQQ/LcQtc16WFh6
TWvEcrw5FgtgX0AHN8wZnn73HMdf0n87zn/6DHjqhkQxpcsXkjKdh5gSUKEb
zBdiNto6823BHdQh674WoeaPnaosIDgnn9NUJK2LTFhkNYQkvStzR0BMlGcs
V2pU1m6sy9lalYwcC7oJ9fbMB2F7nND/yfdLSULSf3nhE/6jADcUKShoBPjw
i0QUQ+d/+u8lnikdUcK7brkuPZCnkShuz0vLVdj24sQnxrkDBzxHS8cXTN5W
EYBA1K5+wTU4P+rFwB2BiCHtdgxPzocbfdu5tIGQjSUIUonYjW1yAkIsheTX
Ltlt0h4kErMQt9yF6311PRfaHXmzFYuFJQp6VOdZgecVurQqTPwE2f8jrU4u
kFm0uHPVwoyEdrC1TmRQpYHXLSiiluO0RjVlAtdKqLTrO0ZB3kGWQ9OxrRIW
CDyGONyUmUI4wFcNE1S1fmV0fhCoW8dgEujPElGo0hbicJWmtfrXbOKFfZuA
2zI812Q0xOGQrkHOJ177vuk6dJRvd7JK5L0okmnF4AT/3yJDGIhodZUFNRQi
Vxx5AqcZAUpsqrlPGYU1ssGMkVbmcc3QbnuuUoMfVMGk5QahXQGJYYj/mXWP
EpXCZDT7yeCf+rD/O6ONe0dRHsCCaKd/SAs2pJpHYukzqI4GZGlBef0qrFiF
uSXPyJ3PC7yfLt4If72uctBA15OhYDltpmZkklMMUX0Qfbd/6fojBRx0k5FI
fxRNmO3bsjahnnZ8OS8o3QIpTLUvIDm3x7oPD1CivgoTZ8jPIt2/+v1Kntss
savqxGChKSPX8tUm81pyO6vp7No9i70vRvWcmsPywfjqh9IkggrfIzzo7BgR
cynV3lgPhkJAAGnqrj9aEb8Jby8DSQZR1HuA/gfU5RE5KUkMa27J2P2w1wNO
221UJEN5Tih54zuW+1+Frv5lHzk0lE/rafaL5QRqjXs/FhUBZpwQrOoSVCuB
6mISUnXVD4kMXsbtRsUKFyoAWcfZTERIzHR/Wh3JyUQx/f+12l03oFliLRRl
+a1MkoL+ilcJnDVOCxOcEJjwCL8Qfuqy7FpmfsCGM2tz6FiDc5PMzRbd4s5H
Y9/Gb9OvmDCyXkP7btmXS59HVb+0xOHVn80OHm44wabkXE33+HPi1aKDIxqz
tMBSRlZhiujNn2MtcnXF8csPAx21q9s50ST4J0nv9CaaC63QTGiG4tYXRAtz
COnnM9UqVYlEu1scG4o327nLo+DeWu+OOfFSxxEAp8sXArHGvLy5G7q8QA8Y
EJJ/FMYTKwOga8B0T871PKdN+720Zd5WDDCngXgh0HBbplU6D9356AudPCFV
UWC9GsB63Hrlrzq3XPbzJYSaSF2jhYTxKFYaOjAlqcU/9bcbut3G8KEDcs/I
dGkjJaH8myPsZeIina958mz+VImxofc7lW+tKN6ogtf9EchPUqVcjg4AdZZU
Z5+n+r8oc9lAACCZLrJCiTX9ZnxwrhfkhNJ2OQbCc2JggeuY7VTShC1240Id
2W1qqe4urQ+SF4eQzlF3B4l/82wK+lI2i3t9d0U6a5b1jGtruIln4FZj3rzp
zT+oyoNkVbgZdscFY9iPM1w3HrnR1YKTQxrw37G8QoIRW1RYF6j4RuzkBHba
Dd3f0T+3Wx1DxzoSsCqSaXlGo2exYDXM25dQtbYMrLOeE69T5fIU3ILvbxy+
o3W+N9sXPmgDZVayGayYLr0ECiUz7JQLToNqk0Wbjmznh7lpTY9dcY0EFw07
BIYRxLgPhMmObvw1xfDMH4rXrHYzVObeG+Jpo2ix52ixBps2x/PZFjR5JReI
iukyyLkxKTwTkGbTIQnqoErwsKOPUy4kCy+RfKD1tkVL/78wO23XQywlIcP/
sxetBj+1QWHQ31b9WOgOGqsnuP9EggJ90hswmrTActsVyQP1HvEmob+gxda/
4G+fkK3k+lI6SX8BOecKLRgPzDh5t4Op+jFWtm6W/eHoOHo7fikvIr/zcowB
OLJngLZWBckQZz4rpgQfFDhTlIH0beX7dJKa7jg2zXb6MVsUWMsetK5gWkXh
QxHyxCybYTvm0CsZW+WgNmhD6Z7K607FUUdSo/5twAuypmPe0D6XiT24FPdc
8YX8qcAV514jzMv2xIYBF1/d7/UfPgY9rbvstjlvcTvqNHmb3/rG/GNXo7B1
tYRblHaulJYQ/ivguY5vNQNs+bozi1xsA/Ubd/7CegNVKW/GaljQ2Smi+6ht
wLhLhBtPTkT4jlV7gemgXlFVm9jmT4812M2XfV7ynZSU86RPvv6MOqKacvUb
rJTMjIO9K2HgC8I7bYLnRdvWlNtbs3eAA6F1Qgd957LKvSPYxmB5AojJLTuc
SlfJM44VN7y5VDB2DKxLDvWB8C2Xtcr636Upp+W+yO+uvHjbejPsB2FjYGV4
JOIQtk7ugqI0jb8dsjYM5uPAcFqQXTY0z1TnNox4LvDxyzMZt7i5myrMDeeh
N1denvET7S0p0dhdpSolEzV3IvylilUkHSqATuZ5GjNsItUCo/BWoO1vZYn4
4bLQb7MlUMubJOugDPKZ/VnW0qldTL6zx3+h2Ydbaw1tLoELp67lti0e3HvD
wVGvr50sPz+C3QKOyrTP2nTUqMfcsAjY02WNbJVO63Vxi1dWy3lbOFoPcWzL
f+Z5ekOXNxDqNaQ1yRRk+tRoMfnyuBs2AQ8pBILjwJII853XtlC5Qsok1GNH
EPJ3FRqpN3VLr9DKijVjn06mMehvHlKzPP7Wpe6xb2T9azYHMRSvUSOykyEg
EfNmxNnu6jtXTsvs/TKS4YItl3XrMkqY0MQWc4BR1r4R7sjRdATwbLiu+vLG
CUp0EDyADMtc2XZxH6Fr3TvG2GvVOi6kLU0HL+QNqpH4qQSXC30z52e8LBIc
GPdTXtm2B3MhuAAOEzgQqmIYOW1C0X2eu4mFcZZM5TA2XcngEMpBWmOQskZ5
CgwWBzYvk5cQWVjoA2UDidwZeoerhic0pZn+wqGQ8BwWiBhLq4gSClOvMdAn
g70zHdGdYmJGU4Z+mmoL3NA1KdIUjAOKAZZIerR1ozTnitPBqBGAr3nPUkpW
iiAEOHlBY6B2lR9bRzOaz217LLJdPxQjhq+HNO64hXeUTvoKCHOLfG8JOA4t
ycaAbFT8SpafFxUoGCO6tpveKhqUzIIDfwAvpNyZl/Mv0HKQZzWUvvtCV75j
Dl7hwnz5szs5OG5s3gHtHYt1vxdkrnPU697TCGukB/RyTM19cUs8o41GWI9k
hb2xYnnn0jgqGK81Yb+JIDMJSloAdn/tA5mqFS2031nRQayKbSBAxzpzemfX
gkcgXll9qAxqda1FaSl5xVXHEm7aCparJmRVl0oe2YYOCPzL7rueELlsPK2O
QYmlEA+EARp2OtuwHHoDYXg87uIlMAfYhPKwHZcvxRYZFg6q+EikL+yf4Y8W
c1/0P78SK+d0ss9tSymdKruAlQpECiB8rs8JnWAzkg7cuu794VNYTnNQ2IcB
/GLBqtJF2alGkXEtJb91QclGzIAdzuFmourlBna2rBb21fQOAALJq+oT7g/W
Bda+l7PiVwQ6rvw2/+2UxqzbmXg3iFH5ZAQKf8fsLa4/u+qW33wHy/6K5IjO
R3TuNk5ivGNv+1181asu8bqiN0WfowRdUFSUUpF53RfhMsDPjJZ428XeIh+x
QDWsnci1d9QxgUklM3giU28ZOgfzdKmp2F3/CKr01qbwZCL3eqspJi24ROnq
sgZfOHgQtxv2Pkebwd/Hy8c7dAijH7jHOwfiJhDVxEUB44R1Xy/CicLn/BH+
vEPGcdWh2Uwhb0hZTIiI4E6ymisGlz7qHmRDSRpxd12d1zUaIb/3bIUKLnX/
IOpaOdt59hfkpuDnmicoi0eK7gxPncKFuZ702BR0TOlMpgDoMCquNJPPn6tp
rU0hsLpgSpcSLBpFnpIq0ovd0NlOMUFRvX9D9n1+4EPd3h2ORGgcVEXecJuu
pzmczjU1x55xR+BRpT/eeSY9Em1YhFTMRt88r9ZR/W6WMkaiA7AWOBa0oLVJ
KTysRG0bCprKtZ2uYz7SIspBcicwknlXLumN0zuTx5eR2hpH8eRLe85CG7nc
zxVmKeYMy1IyyCRpfB+9SagRgWGUnqZyuzXDnDm1nV4gqMd+32iYsdJaZypL
kGo/DjjkBPoORZ01adFv/bAIRQBwsbtbkNd3O0AgJtmh1rIRhaSi09PEYFMl
3sY/zhdTNyb4tHR7H9Ui4rqqnK22dTIGM+c/2CxoWrV/mo0q06mhFYThP+P/
ehPsWxqm7pMSvtyAxQMBpq0DDH2zfvMjyW2BWlZb/2tX5kl8TflXfErqAY8P
7LgnIQlLD5qv3MnLypfXVa+slURB+f/226CTj8DtkGRZhpCGTXsbOh/LTmCi
uVyPYcARkBlOxsoLZ2KHqoU2hZjvkoe47KF2+uF0eqTrJX7dbJN6XieDnvN5
75/KEE3OnzilxnBw8Tmp9Cvl0G+pGL4XIJa7oHbB2+9KHRxlxmQgli6+8szH
T7OdJCcxhJzJSIGzsI0O8bWzISf07nY7uVimfqn6PWAO7b0xg1QlUumj5a+o
JXC9uTBlBiwjeB1c1nlhB6X5/seb/JAIdsctp4mJQioRpGo34LuoHxWQLXjw
Vyc/0MNI4sbZAz2/DkRFKWpl/tsnAgA5+fsJ1DeffHSAFY3pSzVyV2IxjySt
ve2lddoul5ZKNE4Y9OYdEHtddHdCcR6J1Qn8gagsaC28qTlopAJRzVqj0Mru
UjBvOcoulswOD721LUaYhCjqnzfxVj7suXopawgEmO9OKr0HkzVu4ZLZFkKy
NbDNRi7ETXH09jnR9M64N5ePuMolHAJ+prKz6nXjAQlS41Nppd8s3F948bV4
n5aWsvt9rf9I+OR6yQVbZXg+sBBaid5GdZTYNHwgtA/df5BkOG1DOwIxb/mH
Qz0MtfdmsYiiEhVaOTjDZQuhI43CjE+aX8+Bj5jkJWRKBN+HfoKSPQz42F90
Ef9LRDQ412fWJmF2powAPLuFOHGJ6F6bvryygOhvO7WGWUuHRfJfHZLaE2g8
zIdxbMD2ylk5SUEptK029qygob1fz2DJ4DHqqndlH0LsaBuKfbyvxiGw/3wG
/KDsM89h9PnjQbLvHbTYpz07k65tOT8PqIwSojlij/bxl9gW3lI/m4KoWDzt
uwdRz+w7WSUQSxzYID3OUClzaXKZJ+vWr75eTD58Gcej4XtKJ9vXatvgbHDk
iIW2IEQz7uNpMArrHSOcrZN1NHM/dgmAdBjeSYHdlVFnLKnKAx9bF0Q756cT
xfs4sEkpviCZnXbj2So14YOVtsx81korfj1n6oZOsKFQIq5qUhUeFzXsGbHx
H16AIW+Cc5EnvJCYcCD5Cgke7GlFVTguhJP34KpKD0SoAPONcorC7WATU2BY
fyyew09UzOw6q3l7T6itDbxwGNNIUS5kSG6V0U63HbGjRwKw63FhINKG+KyM
IKlJ8Gr8crP+SXFwYTWIvDaRk5cinrZ57KcPC9pJ+WHHArolkrTV2KbQCl4/
i5tQRzTasGH0X4fsmFTYzhdblOSQ3W6ef29AfVOA8EnIsbU4nCvmaYCezebz
qqmY6c1orKQ+zFAj6P84t4jtCYjkKPsk3xwfRsrR0hvqt/VErkzkRX2PaFkp
aif7ybRw+6Egqe1Nm+3CnnDGeLFVYJ9LIiTyxdNZHj8JXLDP8wxgSsvDcu4t
+v1cY73yO+oDSQDfaNvcZ0n7xcVYFDxlQ1Bmrl2VyU0dtp27iMSSdj4aFtuG
w1TTf7j5Zq83wjHxFUewOq/U9Oj5cows4bA0IDx4mD81wZ5W7W2GiUjR2wxs
vHirI3k4VvjOCBsymo8rC/PzxHiN5Xjnse2Gb7Uh9CvuM18iVGDluUkvn1zd
NXRUyodcpMqBNVbliKDykw4fkaX8A9Z2cvP3KGddXf/xg26SnvHX9cV81Mql
iMMsbsQytvofRiVI0aS3WM9o3sG7QuZnkfkSSKk/1C1xSeXCEcTuPciE/cYq
9WFvAuYIdzrt6inWMqMU0G+FHgkgtO/4yDbnp+RzXuD4S5HKKhTb8fy1Djx/
AmxnTCSiIbOQk+oWij5gVXTRfVHmJBzr6Zzdm4TwBey8txu9yvVSTtpFf4Wn
v4JDNFya0DBecC6bhYifq/xpwMfppDrVci93n4D7kckMXKSY7SVvwhoVCQh8
xC9P2nGKJDg/ka39cdw6jOT5h4SwXv24V2dUvy9tS2Kk49OacdPAWe8lmB34
LbqC3WE6qC80mIGKCYhNjbL4JG9z/3psFrXIW1kgDMIFF7wsjkz02QsFc1v2
FqdBrI2t/vH83Lr8YLvrJ5D4BfRcSHE3BYICPeB1oyx6ejwWXvgSMd0dA4PB
QP33yxmBHd2ngK8LQGT20G725ShJdDuYV4aDTZOXGi4MzqgJktrrAmmkSMQT
aT2zNY1w5DcMZh9hDveXwIa3g8k5TA7A/Cm01YSWG+AeIX3yzOVJo86PJ240
yFRhZOx9MPccPNfo+9TcIMUqRWDKirlDiiN8WeBSGC6WeWEBI06ldJK2OksY
YLgxhrHTu/WqNYp5K2I+1FBTbayLqo+sb7+IZGS2BTebP+Z+pytSLhou654u
iXVWNBvARwGOBe6DjXzDVFtoYrhCthvKXs5Sv2R8BDqWZ9INULbNiUfDD+wp
MfQ6IcxYaSpewzq2d3jxICZAWMj6l73hwabUsVhL0h+xpe1FPx32JZTj26+b
7vgtf99FH4tNwo/L7bMEPPmLDq7O+mWxqQthJqiMRz/Pe1gIxMsFFx3H1M7u
nUjIblVn347wuVC2GD7VC/vH7+uEmRtiSEtGLFUs0ux8YhMPoqKP5aNl62Ot
XqHck2xhmLucg5SNgXsvhpcI28qHYKbtnLRAhHEooYfG6RqguzkjhrRx/BfG
3u6CSIZCchltPybSC7LlSR+uVIYveETkjCOV2nubew8i8OPA5x5+BGbYV7WI
L3vUXQs4Wgj5qDZHmJvP4y3LXPHo0ice+DyVDV19atEgZxlbsNSFmP0XCsCe
fUXgmFiOiAApXxA1fxIjefek4rAmdPhWLsq3s68O6sfpHhJ2wbsrogKWc47b
KEtxjTK62YXYlj/A5cqHVWcCCM3mLaO3BUp514iPZDx24k93Y0+2f6WQRaBI
81odqoixtUy/RTwuEPovmkK0ll7lNqqtXmiLCzqncpd73qAd2ARxwW/eU0j/
GpsOhP3DF+fdyFHBnm5LZbo3H46YCCuXcKHmvWLWqAIqYukMUlxTqVq5vB9E
aaEjpIaDj5uoRz84peVXHZ020egBIe466vKLnNNduRbS964JO6EY4S2LYSDm
KJ7AuMjDFz3izR5z1Nqz8Ni6xcqlmdO1cRfUt/3wKRaYKcG4ur02VkOwYOC+
cYz0dV26V/EdpvsTvW09sbinvIOI4Mq8jxnvqcO7a/fhWej3t9zs/xsbUBgT
CBsqnA3voYuk9IGzc73tDoyx4Dtc8WrNwCGDIK/w8a1j2vO9fGEJUWHTb0b8
R+MW34dS7HSDq6ojaAue6Xi0OaFhh3t+DlNTWhCTFjnwrd1FJvuZu9hg94u0
buy7PRZMM6lIYH1JqvunljU0UDvL1oAjQmE2RVcKce6Dvwdnjq7R3X9+MgYC
WZmHy5O3alQIVpKqEFRUzd0XcZWSkabcqbTALGWkPCxknWt/rMDHPd1/6tPD
YXqu6+k5TNmv8Xtuj/FeYpDP/HZ/jMhcQtgRtYQKwv4G1TSWvPohdIHyrmYQ
mFVwsL60bqdLaHqcdrTYtFeHAYEKfA9OsQ1IDmlZDzxxjpEuMG0hbtdgfvFp
u4ddEB4aGFrqFjMexZEyHWuVBsQNGQNz6Ky/iqblOKP01dzkoU6qxZOjZqOq
pl9lAfCapxQDvYOTxkDoWIthHWfHyPuutAle/rU6BuImjLA4eQX/YgULylBu
Wjp4JBX2ilV0wrg7U3FdAU1IBYnVbHQIA3Fe5EBrwiYEFYmB7yHRRwt26pRr
QI4dSH7d1xzrWtSn7VfI3wxEeUvCtENU5clsjOuSHpttE2ZNL4yRmHvVJFt4
kF6ZjggGFJ0H43QIW3zW+uuK6/dTItPI3aLuEfIrlRvd2xuiQXGaZWmhgKk8
NUPG0irQNkyw54Sg/6nNjOxuAfZlbGQK8IbQfqQgmB2mvimXJSzJkMJ/mi+o
A1ylh3QFalSisaPgo12LxR7roxr/UKwjYO1mqoJs591KO2ENxmHaCssVqup/
vTioInvSJwKyyvtzQuUYcbe1jCAb85frtakENt115rq4rbj90XuXrjwmH4uy
xB7GJ9+RyrpkawDPrNPpJTfgbCp7VaWSEJftnN16ZS0q5+F6OQo5Na5C+JAk
0m2zCuLDF5bPVc459oInjbPNThr7QUEr1unoU2+kr8YBSmZPn+UjJvaPNx4G
2pc+8c9Yi4PYhs164hKgRtJ0ja8FGffzuWha8ckVTd85HKaTjJA+Up884Xhn
tNqTAI1MK+oKhZxLOgZigml3JHajTd4NZ+ac8PeTKiPsP/lk/gtRvahxWqoP
ny03k056U7hhQaCnE4AWw80cmKlfiCq3P1ZGZ/o60mT5AYLIPy5y5O8oAek3
lnySd9/CktyKZ0LUCvVXZa88ZHOQ0e9aKat2bjBMwFLyJYV3l1pmpSqdsTNj
vSdz/XAkMiSRmUvOuNX3au6fE0XvnhZZAFXautQBelfpcdBE4ebE7CWoaFj+
pBDfgtZT36e42BNWKErJLRrmxHwh5MgSpDzIMylaZDDyNe8/dGMt5m/BUmQ9
DPL9sBOAWnbGyzcg+HwWfuEkQaH653Oj91S3rnSL2GtMvn9PxkHiQcl/Oj5c
od/EDkbtYJbVzZY+4zz7sWd+xnDe3EHYyGl+g8JfOYa9w/neSjJeMY7NQd6k
tA1ikzINapksdCVhM8U1XxBxLRI99rpEVRpt2jmf8PrE9btKthzjTONTNJoP
Dr0WmligegK/DoeN4dq4EWcQtn4fflqz1sTcBOLp7xQjj7ah8Qcao9rXqObw
wveTREMNIH6Zh7111XTrJmmsyCWY62JZh8xm1czNypZQdm+L6zJGWJ6cUI5f
1xo1o3kOM/TybFxNMInCHblYm/DejOyQqVJsfdrrkDN5yHIEAiEso5y8dNoP
LDnMxaWqAiWVlYDczzA3Gf+XX49NR6TkETp/J+gRfbEOxIYmYMBnNtly0IQE
9EYKLxiM13HCuYXGyazhWOo/YQ0/jPlTrLdminw5uL6dWTwqGBh2vP/3t0Kx
HHO0OnhLGXKEleKB90Tgs+jM+S9scOCmTikCek8NyrPqG2itGKo0DfEWuwGF
9UEz6TMPuQ+k8feEdmjkXRO9BL/NtRLjV6MfuRMFYVlcuemW3rjUpBYB90b4
9FG329Um9SVaEfRez0IrIMJ3bzlAF0XFm6GYXGVbU6xMk6W6D1pVoXQ9z4Ep
M2d4JOzoenr7a+EtFdy5hgFKRf6A2VTUQVclebQMVSpqcaE7fVE05kcAFISK
IkyvccOykPBx/mOE+6Ksp+TcpONYTVeaKQ9uBNHIgyLnK20kGIh8rnPFWUk3
v3WD9bBysv1dSB7KdyJFgdQmhs7VWwCQLE0jdKf0M5Y7MnoiT0aE2gqSDAXh
NZ0bje13ArYje4ylB08iFk95k0T05nWiqGWJ+4CCzoeCG25MxGTvAGWYpDrw
CXhpw4rnum8lcq2EkpD9+g6Nb00anObHL0dX81ulOEI+BN7EYmhC2IMvU7oq
MIqz5ODRW0+7qO4Z5ieKFPS1jM7Xj6EnvzGNAd6/AvZ70CEbYmZcgpydKsPh
5u0a/dECaB+0bd0+c7RchHEjr31GWx5gEdb9LOYiTCs5kVmGjJ/uOZUVKW7/
adWdkr/JWzOkoL2RdG5aUBFQ+kreEWBbMRg0qpMDLmbNK7kZGcOjS/8ccDF/
HSvmh9LAn/aZ2lTXQFftynYI5ACsEgABBmfbcrH2DGraph81bV0zTMVIfVKF
t3nQfQTlz9g5BHx8PI3OgBJPrwvDuUoFOENjTeNgXIw6nfXJaYfr7whcRvWi
/1j8pNFAa+qiRERp8f5TCC+S9k6Ns5buviwlT8TxeKM4OMhXgjI8jRxwSvWK
OMU+fhCFDYDmN43k7gKJPJsVkrNYHv65fQjc8kp24vATBQxM14IJuqt8Kyo1
7bgB6kkIDf3MVmp9hpK36zsOIIqmwII4akxlpTeYFlbGONY9mXWXfykToK5V
oyZBKxCmdzIVvun8f07XTTpQzU/EsiUWXm1JeZScYuqPQPqxDWRYKsl06xi6
WD41XGdPWWPfD8E8f1hLwi5xPpj+ZP0CHRUT+WcAhcp+DBQwcvoe+cbsVBKK
Zucz58vKIviBUqLqcWZPQ9OVX8YbnTEpECUo/zP1bP5l0SDbjNkECNVWatcA
YZPVKVMoNZvfJ8a+EWKUH1rTfdKOJO6u1xBn0vpe6kNzmylYiTUI+S0HWPeQ
ue/RuOAzBL7miAmzUVKPcHTFFIukJPdX6kxA4k74QKk6tct2eANZUPVr9J2k
qyxOzcShfONxiPQ1N8jyS+Qqz9xWoH+q7ThB7Wp58AKRnnvrovAkeypTFqiU
jHonQEFYyla1sRLNGk1Wr8G7EZKVuUj2mLW76mkSzK2yNpJxzsgiWS0NZUv6
AG6szfLYj/XW8DXrunMGe6Iytp83KGlCI6InGD9APrZEstpjq6nlMzWU46Uv
SrFb8tpIgUBulMHHRgmS4JeLi7nmi3tiBMdDsUpyYkhm+UNDdrQAleV6d5D0
PtzAoWidqvaajjdIBDnrMiFMYdV0mMrBors1xFvDlj2324jd5rJcPSyCM7m0
Bog1rujDVDZm8xoOdbU93dc0a7niNh9jTdtylpskAANr+gwfe+9+6G/1Rb03
qmc9i1AvV1XHInDXqJb6tHPSe9s3ktn4KBmLhHitBuvL0OSq8ToSwC43f8wf
R7mekyr/kexwJhLUVHTQajDgkFw92nANzkQsXRXs/68/IVIHce7o4STVvRzb
ijWNc1mL4s9QFAaLfM1WIqs1tnNT/HvH+6nkJqwB+N8CU1IuV7B8Dl0jTHdc
9pSYWAhh90d7J1R2ONvE+tF0qIkrv9ZMPpLIYzFZUaSphXvi8LfrLY1WlpBb
YPCEpHHPSvHd2+GTC28mBDilVWhDwjjFViR5Fz19P18x4zS6SKGDkP+0uUmw
GNFZm5QB4o+Wk2FSyjkdNUJ+sPIRJuhKr3mv6aloN8J+nHej/uBULs4pthMg
7ZGp+N0ENMwp6PAEzOLQ4tRL5m5fadqMGSzLlZgCYhNSUKcIlOHonBJA2N35
qyW++qTfgk0TlAaEUchxBRo1TEpw31XYgC/deF7kg2WtX1+VHL6vssRse6O/
SfmTuhf9I7TBVTq3frxTv5vVnqyd4DE9u6sWZxtPyhZw78nxcdY9wwGkiceH
qnYc2PH2ABD3vhzl96j4aP7KVGYk/pO8V9DVelcjE6ERmw6YSsAJk1vNgIbK
DutSxbQ7Bb7Vgb15Uqt3EbDBEwZuSugu5h4zbhKeml4unxWqpFdqLUnFn410
HTUyYxsJiUdka2QbOJZ77kVFy6fDPUYwa6O6JUusK6i3W//nwy8otfPaABTk
r00/qO/YOujzRy1hA1lylXnsOkEGNulTQ/1q584jcGc31GIgv8TvrSg0io8K
fAc4BgayUWweu1BDfJ2kIzG1jT4rzu6e2whByl7HgwrhjnvEkN2v8cNvICvr
yjmBIk+Qdk2x0+0Fg2Tuq0z5wbqFnlm72H1wJzLX0MUGZSb2MyZDmfy51yyQ
POamj7+xbkPLfJG7nECEjmvSJLtfXvkRZ9LHJje3a2p2oKjVWD19VZThLPN+
bu8tsmyPZTkE9QvUizEJ9Rpdil84mB3iYXWEe3v8+gGOffuYXSWWP1nf/pe1
8snzg7cZNtAow06eYT/I0CJ/EMIxXsfPhf9blqciwD0YPSJUpyWCSr6y4Kez
n/U+YQVtLLhBRakt4YRxjmPkCccS9V9LZZ0LUPve2fDrL0TrUDAb/gsKnXmd
t1JOfSZX+R6sLHyFD9Ln2zI5bliGK6SVl+dYleBU7M3iFaySofHaDsSzHNXG
oCbIrPBF7Vo2EzlFVbkRt8WzepvmxzBzHj9TDRSAHfTgRb0acPpUG3NV/l+s
+35vcll4u8JYG0dcSMRtLYM3qb/lBe9OkthV3xZc6fTRGbhvKpi58PNIonOH
DHWYSC1a9RmdlQNc//EtoUPGK29wcxQMLBJ2VY+qJYwm/e3GHOBw11z0aMmP
ukDnTjdSdH/oRZMkIDz+LhsilT0BwSYdGVEBqFum9LdcNmUzEDxU0wM0zkYy
weXsZvR2ZDWKMnNBrghie8EytHxaEDnfsYUsghNzlVYvt78nyujjZ9Q3Pp33
K5P2dveAOf9INzZ1tFqESaEt0gRonzekS1IkG1NauthLt3p08y48+IylIcO9
JLJkMm8sVpov/plv5wrStm9fhQlPKgbaWjypYDp3bVdChiMSZKnshUQRsI/5
1XguqZgz9PhhwdPi05f3AtGm9YoDY8kyNUhuehNNzcvuToZ1OX3HFCv+3++K
iuicyWUoIzd5uh7G43lCNK9J5PUqna1+xLi18TzqkecSTwwpVjzSwd1yenwF
0eluFWBNAktOStHIVp29CdGQ403SIScDvFMXbSA70doRxco12mXPIFrXxXIl
aV3ASy0WTmWuiDP+/SDrKcK8SnaieqpGSDW3xQQSiXCB3kDMBj/sjyoaHXDj
CQi3QY7VIXX2K8FjJPIEAa5TUa0PjhLUI28qJ5dw6NxlGVf7cnGmwODOFn0K
bR0oWyQHS6LszljX7dx9KwlSoqyjdlPe9ibt2RLkILFEBJTSw+0HV4yw+nLF
cBaXsqcDptFo/buPw9w2r2d8ELDYEbQCQXlGNGMNpe6+lWXsaGyM6myMpb1L
vpoY/AMVKw5wqmJpkPcWTyufeOqMwxBZ5G7RY/yrLTeTNWXr17LGhKyoJ00p
hwW3EZvDyh+pYs4cKWDiAvD7QMzwcdiWl91X9k/U0KuSC+0eHm24lgGCiEWI
84m5NGIIT2DxoYm0LiLpcptf4V5mVUIv4z42QEDsA//kkXGdM2TPXiZaHo6f
KmqnoZ2vZGXtmXc+5PcwBg3CKciegHTf749WttZRXyN31VkSA8we7/9LvkXB
i5jeH72aiEACcABr3rOeLhRtOPgcYDA2pynjaM07pU3wAnu3cOzZou0USdJn
n9b3C14S9bAAYVDCZCaiJUpSbk6v0Ova5qdRnbo7FAN/If/M0C4yTYxCXbGt
id4PQIrIWqJwEDxVjqqj9sl0kaWOAcsCnIBSmANQUUHKLoJyLmzS3Rv1KCm4
h/jZRqRw5+OclgiAIaxT7i/un7vMw/DEdX/OxGk7nSQLh8OyruZu+MeujHp7
K8qOHU974eY5PQZgCAB9c0Ku6uooaZAHO5H52ginKu9OfRAxULm0NowbiXMu
y3LHeu+TT9SHqrtjxvshXhesQXrGFyszCksDwdg6jNyO1aO3xIhq0x6Y/QY9
7yiS0wSOXSSk5luoq1SI29/AK6p97iCUfBDMWdqnAcle0x0zMu8W27qQazx1
8irPxGuphkNIljznjVsB7iHXMYB/AZsZhXQGcvTdcaPSEshZ4tYYVKZoenAh
+T5qkOVrr4Ltvs7NDSz/t8TFw58CIvDXg7zMYZQr/QQq598fFERDjBJav5sw
2zi7ofm3PJQohhTYgmFEbmpAzBtry14EGlRwFACwpuaBUyvhPkAyjcgt8MZ4
r5omz0YQXBy0wSy6p0Afiar5bWR7ccp8lb0Cff71ewdqYkDf/7LAbdxvGi4P
72i5HWU6GPMNblxqIjRkaeBH3dODcKOhgpmJww7wXF4M7F06OpzkVhNqFkFi
gVDcXCYkWGpOyVSQJ915fhfmE9723NIG0FEMmYOrHnmSK05ol9+v61RxuI8N
AJIKXpl30BU4nTnhHJ5uLLX7T5MY4oNLppe+CQePIdwHTFdQP2M+4Ty9b7J2
1H6dU/sJLU1L3hTPFAHkif6dr/VlOsusuOGVd3VedUY08t/cIy8JKjs8KE3O
kfFOcDj82Nv2CDORPRKBhIgoqhh7OS8ecCo8dV3XmnOKV5ersi9DeUexMvbJ
jKGG3kQuMQBf6krjePnT9s9yEnAhN5Z2sCCaUsGxBqBJJhAzp3JXuVNZfYVq
SqkniHB9Z2UVhQvTwzwNiwzfklCkfaEhTq8aG4l78mBYmmnJ9xg6THORKR1h
hZzI9QKKV3snU7OFmZGyAKs7H7DSosOby54ovLq4nKk4C35UP0rSLKYDPMsr
+SAixNniG341Bf20EsCNdZkhz7+7ieqhPvRiwM+KgZ5IJcsYUwFMsvOX5zyN
SmubT1tZNbppaCpb6U69rgo2XpE21+eLOgINUIPi12D9ALGIW+cdhnlG8BRm
2SQPvy/CS/tuOBz/+YhZL1aFelQTeQSr8d/vVWnzydjnVQ3DVKm4bD70Ethd
YJZnW6OJrLNDzQLzlHYJrrKHJ3ZEPh5P/QTKeCe3P8c+XAq6L0Pv4TRKfCLD
57OBQygwGm+Pll9y38wR5jyGuqEIBSzKwhOIe8u5vx/kI4XoUnLCmUgbjvk/
IbCH9m/PLCRClmKUOq13OYrRs0nHqqosJehoDAvYc8IgkNK3w0kmo0aBJS+V
ykbWdSAsdUMipbpTSGPJ97KEW89NxUfZ8xt1uOJu0bGshabJZ8ikKW0Nzc2h
areT+1TRbe2t1EXwrOQwn/1xdAqN4qCSsOsxUUNSsoIlPY2i6BL5TPVnf74f
uoB4BLXg3istgRRBPV5Zu+ZEzgZf2+TV2hx514iTc/mkil5/q8DKODAt/GBH
DWSTt8RCRU7rHTvRRwiEXuEFTf9QIudolwTSHfQGL74I7x9mm9qVEX6Y8aL3
kG1ayx1nqVtwmw/wgVw+5+Wv+iNL19xwGCZfze/uFWDjOhgOE3gJOVTt88xx
jpO2SCHhcB7nUi28viAGtswzmwYc/nDcZr7DB4IX6KgxwUrd5TMi2EAkSokK
yUD/iLAhXEhzmbQOPi/WweAemf3zz0ubz3HmuhJPXR5o5U3mJB26VrS0zJ0r
ITq6oiBSGaX5SeumQZD24aq2FHuOTlE6Lk8auHE8e+qltUzNQLedDoD3jCSM
4XgxZDHoFdW8qa/E80V+sQvgnJHf9b965GN7FvnYHH6xHhR6EJXtCBf1OW+v
ghAaOOJsDDQbv8Is++Fxyx6njoCUKDKVGcU+HwxPju2Bx/GD+QxKlykEC8f7
B8yF6XAK4ZbQmJQnQqlkNpb2kBMwRhKQ32JNzz8l1BvEKzVZRIouqeAX9ICX
ZfqRd8/SIlpo1W5KcF71ZrfVozDhx4tCFX2nYvrrsNSmZiwnVTKnRJAXCYNB
t/eQSyLmRnmWTIFRic+J21HQtml80vY9LgSoQbj/TdfpvwouaIbzkLoqOpZt
iv1wtKQ7OeavAB0fSD5KE0jO8aJfgZ/kh/q3V5PaCibWfURutgG1NOwchlML
GORp00PP4IBDv2gf50QWFN9Ioe2MJw8fzNpI4hx1yE2cBT1gPEXu2Ly9OZAw
bM8TIlaYSpmcOtp7MH5DiDw3l+9uAjRSzlmbzHO/CzfT85gdDv3vGGeWCui6
y8VruAOG9+qqhQvEaU09wD2FDon2vQr/3NP1aVCaYR5BKCC85+6/6FgtkHB+
h+Rf3kqg1WWRMW4v8zPOORn/t1bzL1j00fu1hhMzncQLZofV1k7cBLuyXrai
dGCmO4Eyzvhk3/C3kszhrvMV7MmyBejUJNJZuTbLdky4Rfwx+7dhh0s3Th2x
tpYX96SoddHxd7AsI1LpmufBpEFv55etRNz4ofk7znSIaF3ENkgPvThjhizO
vvt6dkDVU1QHY88gjyJYLoqt0pzjmyrkHR0zQ++hA2GkxMSaeUrZi3lQ+6ez
JsM4liTq6OCAfF7tk5yB1IOkvAIPuSWwSflOmTyt5d3ETd7fm5wXEkmUNtby
lrf1qiN1AMAnf878YUcEW3vGxPZ3wGlG1Od8O8dCjMnK4IYANqp2lZvMbxuB
uS9dvVoxRKsdt56EAuEvWco8yXWQ8j+0ABQMX0gtjOMssR07kSWAoYn9Z1hO
qBc0vyFK0MA/qfZtOC52V1KpOCtZy37phoF77bPgDJz488sNp5wYA+hdoMOZ
/pBiPWJdqDe8C+OkzuSrE8S9VVhdKLMO+lLv9p9Jmp4kmZqJ76wOEtcl2dk3
jO1j3YS20gGOdPH+vkHmryOXMBr4eaMdbGSmMbbWH/B5Xp+0Ua6j4aFz3EgE
qmwm8XCo08AH0v//38TCWtYAgwTjxogr+Xs/tPULYELRlLOSBZr5HyeGzlJ3
Zf/hm/VL5r89n//53LDB569fnLLwd3bejds/X39RkgCQ/UI6OLrNgA1RLzoy
GVbb6yFAlvIn7HEOcU8Qi485YAZLmwqPrzCO5CypCmwhgggYlIYHO8DQAl5t
OWL4to1RH4GYebp25Vzhn2kIsshrFyWm8fvTB4nVWla4L+9KeUQC1pxoYhC+
1/FQomPMCCmg3HHEgH1/hDXEkcb4uphqHlLWU36c4UQvCxVZUqDlg9qXmasC
5cqI65P1WJBuLnc27dgFSGGHmHbRp3Ea+2QIsJzFWYvTQlLefjSdYJlj6r3s
CFnoBjaSb6mrOIm3GceqnptG+uR5VbsrScEfHTMGP9XXxWj3DwQ28vhMvv/i
jUH5Woy3t20v73Kadg5z/nfpVIMlYOfzEbszGwaI5LBM4habvKACJ2CWdGVl
8HRWJ/NQYZTSyidZ9jIYhbQtKNXVpOz332GhnE0GWguuYZdrn6pOuAzvbL7g
K69fbhsfl79AA1VwmORN3Faj+bg4uULMECSf9FNauDAlKXjR8fUppQCaAV3i
XwxlLxNz7BG4F0RR4Goq/fyrM6aPVNbmre4mZ2+ujBMxZ5vmaB2MF2drpbWo
tVfk1dvBPr2g3n5ef1qNh54E3MtOdZYPbiLIG5DVU7w0y4H/7kHjVW+U6/3E
2tjzmLhiKynlR4dzXXyH0dN+oxc1VREV9baorneKHFmwiODvNHAOb8N58OBh
RxIHnXZOoUWwL9X4H6/0Io7fRZgf3O/Veh+IineRmmq+urF8YwHeb3sQwPTy
Y7miLHYhqbXXKlsXvCkmeCdyJrpxZYEJoRHvuJuZ2DGN+mWaYC3c1xDLQZ29
4/OzxhjLJRw6GR8TmSIH9mzVD4tt5XwoKVr1lQ9Gv/W2quivUpYx82PWDFwd
EoU6eF44m4kDox9wHNTTByjyjrU3Pdpp1ZRdk5urjNt5fitL6N5e5KXTKY4N
0WlRMEleXJfD/rUyE9ZD+bJ5lnRCUiEjfql72d6UW5goFF9ab+nLAKTuTn2v
O826ZhRftuxfArdWe88VSu0c73S8XcE7IMSx1NSXix7U4V6l6L5EyAuYhGdu
jBKMNuQyOjwZfIRe7fqjAEtcK94a4yYuyA7ISFv4p2OFkR3Tm/FjKwXbi4Jr
5pQKF4Npr0A9yhlQu7YUVxMyo9EVUL4qgJddM2DGqXCG1oQ6yLrZRksO38XP
XQu7kCmXR3RJQRhm35SKBERmODdEglgmXfrmwrOWtznzogZRqiw+ynZHz9fC
H/xERlsjsfmWyM2lWHOWEVr0HHcV/g+QRfh1X46e9U/jJCNe/6dEjCBSpEQ0
+iHjTPTP8t1hLiyZjZd4b1gO72anihHit6RxxDSi+06B+uPKFOnB5pkGOzt1
UCPiCSGj0N7cuvxRNa4Xcs3JJvL435xeDXK06i9hYnCqTaS5jVEU+5Xy9AmG
oRWDrdfFOrwxNNGHTbSIe8HyBZk8tuoAHrQxNWNGKoPGFTBMu2VK9qhMDfNP
khgc2hrIyBL8BdP43id/znlYz8xBC/CXCEGbYRPErFbKY2tKI2wWkkOS8s3q
Tjlhp3fwlA85BW6t0xncoCplc3ynCDdiLcDmHCkbk2L3dtItAB5K/mkU+tVp
ZBXxVhdPAJHiD7EmlgsBf+CNVZidUYAQ3W4qet7V/MgfJmAl4MEp8dfHVACo
UzOZZ9gofHiExydpJtgdnNkqEmEBuWGCmxuaAFBQYUuUe4jlDKQAycFPhcEe
Aj174jSxvx21JSMiWLKYStyAurSY9bf8KuLh60ez5CYGMHLVdHXrVgXyZhAn
L5mcKFiLtyQqPPBhbqGj45XbayWEHi5yxX3RSJGGEEmV8JkPX+/2ltuStQPN
0XubEV71/roKegszabXxah2IziAyJIUtoPPtMH+jybZo4HM8oARPBfBx6J0C
nuO7n56luwJCRZKx7sbEQbl5MnxjLKXTmJjxAOAf3wFs7aSTkd/sVROUm+nE
V14SiJqAVbLiLloAemXGIOjOQBQNr+sYnoWwgQsQNo9zlNBKDjZTiV8lRz5z
jTzh91tZj/uCJb6OtZLVuu3XP3Co81t25HMSNOjtladrIRm05tc1oobO5UuP
9+nQSiuqg0FSuTIx0BvdidjPetIRaxxYEqAjj7o2s4QtsUBqrXQ8q5TF8LG4
I6Jsykuo1oz7Qfn+C5ct1b1uRcfpU/PTJ9vxXY6Q6X4pZDK3TSuJTCuNQIhr
daNO/VSwc5zxNsFVgcQ9/ekLiccIoXcpNgfeEHOQLInrrWoaov61l2WlR038
NAQ1i2S5/lhiv7UIfBFl8b7qhyYzwly5C+CAwpjyJvgs340LHFYIVxqV7s5c
0cvqiYBoFaGxHIWGRryZZSRqVI/a1rpByxmdN2/60+8kgwzxcuIBNBoEPU5m
kyagp1H9/R2bNc9ZdSG/zLCfzeEXxltZMxZEXOYqcZBBgZibVdjBZyoN2LM3
p4TPyK5w9yksvwFg1C5k2n0Y5BBgzMFsQbGGxsX1JPT3p8a2Vl1J3t4ui+9a
JWMPKn6GX1XpRTtr4EH1U+1osSmuXVaDSVCsMdUv+yNoBi8ygonXYL9G1VW3
nFgUNDCWhSs/hC52hw8M6DP49UoWBsTGOFkkCo2TOI4IOyJh7x3H/s/1hIbS
ejA/s1D53Pn6upzp/glA994Qhwfwjsf9zI5uUywQPSpr2VIQ0oq8YMo3ARSd
j+ynn22O+OHrE7JZz2KPXBwf+++6OOjeEqSh6DGOGozF9sEMzaVOTOPbf/Lr
NwOSNACjPFGouJXKBp4bHV3KcluUekenab7rFh4j17jWXW+NPqqywRfAuWZ1
1vT+M1d7WF9mC6OmOcpP/ECjbcKwZ4yuFyNXcuI4GWQXqB/Ub1iJBJB49UyX
D0n+YznZKncj0PuSyjshbpwt2NKylZarZA8OYeMAlFwwdYl6qm08SkBtEP0K
LNdp7c1V+jij4vqYcBoV6QGJ3K5TbNXw50lTYY4tDfXWJgMLvfpfgJU+aJQm
A8WMr1+2NIYO4I3Lk3bkl1c9L7RlzGm2r78cQwL0gejRkXzqwiWnFrkW8/k3
z6FPb0rXMPcq6iOA0aslqN8QjuMqsPf+HZ425LgJ+iPSOF4kE5cgrBRvxNJp
zGEYWAemsK4xeNiLORC9pLNCfvHEreFx8fqU4E9gNdW9tZY0VfA2VK68rtiO
oPspZbKKCoUZ9j0lUKHfnkZVVrs2dLOClA7iTtgv9R1zHNr+O60bHnGT1hU8
NOSf4grgBzoQU5yESi9v4PvKN2bJx58GIGZltCF9rdJFufrYSYgePEUzMOK1
X/+UdjTWUKpzRosWEXEbkOTnWfs7sgCGB9f4EnJ9z2DaOArV6ZYpDnZl3Wb3
RXIanCqS0N3tq0kYnfkbvTVR2RLv+rGMvnESjYBw0UDTk+9yKYbDskb29xj9
Hkmy1Crnkevc4D+y5i+gvEgj0SnAFyLrQ1AGrvRcjnUkHOMO152fwI3xm/sZ
er4Nibnj/iGOXvTdyrIHHgMvfuJLqAZSpZD92w85m9u3RT3r5G36Jx9FP2yw
b1dNdU15yES/jK/XTrRMG5UIqtjjWzt8hbJG+tDZF/poEpK55ErnOis0R0Jc
yHjWkW4UvXNJp9Bp9IE9usfikfl9k/ANIkb3xp6gIEvmh9VYOVJgXkyoHcJM
PSzePkIO2rFfRKup/MPCKaOVi7W54DNH01RhqjkuW4ZwoXqUkBkBhfB1OXC8
iJGKX8HMKPiFk6mgaJgCF15SeI0vb09kj4h9Oa+QHlsBQp5KB8BtVyr9CwsM
/X3EzHyA9l8QxESflLnHKH9ivaWDjowPMo9GBlzP1gOWWcMl0XzTM5a6DCLO
hikI4MSTUcVUO1xMNqJZ47/Rc3aoDOkeTYVU0uVyzmMxo52AMVY8peRVT8uY
wzbCgRbHS/mD1S/5qPeiOq3dQvbPWWNdGgu3BXi18c00aMmMRIQ1G/zpzEn/
NhT4Z2h4WXXwgof9KQOQbn/iK9E+dT8iI+2vOYvdQWDVXa+X+SnHLuU2rU4O
L8OGEbHb0czzuasIWJdOATVRTJDK1jFt9ggUBB2t871P0fsaqK5nA6CWdXnq
LfMkZZ7gmPUFL5ApjUbdfigIOdSBUgDwaUgDGfpQx3HOI6sx8EsE4JR1zn8s
u2qzxfK10yGEO+vtgWWwnqoiWrRsARhmzfvzdmdOwyWY0n6qMezR4FN9Y/Ig
KyMuclsCfkO/PZI4ekfdktwMY9CTasaXXV/jB97XHUF177pevZnyegDnT3Mt
eDqUyFZXCilXEQnQtcdiBtFjKL7PObiylmgPxEIV7ZAzVUmQZtF5YVAtkSwb
NQQmuUD1ZCqP7ypk3ET7Y2uoGJBNkU53+vpeekNwc+PuMNatvJoMiXBKkXws
xuwYZB9l+Gkc4PrDIDli1Hiwjz2FwHX86QdvC25PRhhtSMzpitzflhA6UyGp
hiSXovoncMgOqCx+gZw0siOORLiIUxXjxEYUlkEgKntGctC17593N4f7Cs7s
sM6k3EvXfqMicwsxt+2ux9xDFq6KvfyPROCukI+HKd9K8nA7W9WdRNOCzYLn
xz8pwFb140ch7EiRKMe6ov1Lu4YxwbZ8zUResTeuAIq3A7co9bBpEjT6268T
OJsVNShMU/CkZ6Gxm76IBiaaVaeD5KYukU6c3cJvvvc9ta332TthIvqfDFc6
ZOlC0gcwxYcIuV8oCzJ6yvBMiRcX5GpHE8lo5BJn4wjxFeuR4TEzTCvpBIa4
4ovT1HMSyOJybDJnny/uqfzs3qZKyOOtqSV6kLqOwHBynNRzNOHsLnXn4RbN
8w7BRjrttMJLKrvw2C+nzj7Szqc3Wup1wunCQNM1LGgy/Dso0Bzyj2htDGxn
St2MHOzDKhHXqzeWHgx0SpbatszwNO6K4yk1p1uljI4OLPrdE47yVY1W1ni3
gyE3RrD1ea3zunWFg8qfU5Zk95xIiLNN5ff84UJkikXmXYgcTABS9sZcLOsp
QJN8duatAzOw07eChoNjrgRqCsnuTN7HMd+1hVB+Z1097d8F/T3SsFCAcx0x
Znx4rIe17ZUz0zQB77gwtMO3o03z8iKTYlMmMHfKBLXw1VDOAhro5RLpfG56
08Ob1h9rk0MSD6RWzIw2rF5wqtWL5lNbplS41GaB7uH/xaMw8HOe2oogL+3n
nTf9QQyVm45oZ37/mF8zcisrMbUrpuDo9gGbrAjNQAgHMEuwUBPLcZx34I47
EFv+9yz9TvMYtRMZ2OsduD2Ajfd9ZYQkzyaFtdXk+HbnlbJnoJ6aPPXq22Xj
MMm638JxIasjHONszVbeZFRvYk1AiPfLz6AMF/cd7i4+Yb+BoWl0KafwDmkP
eEhHKxOrPPDk1TpD/rU82Um5y+lTrfDchFiy9RTH1zsDsJBuskaRhoYMQFup
1LgRj5G6uldm3CxnUFupK3mNkqaKo8VW6VHLY+7eBhfnsPNwjxoe/bKNZa6m
1t3nF57hhiUbfbQU+IRgW22bXvZn9EqUGPSvG8zlrOl26Z3RUrIMsoVzt6OJ
nuzYMcjtXPqmQgFDGnePaEX2xLl7a6eIxAUw6CaS1k4zMyYWVFM4M9QdOZaC
WBE1niizIoBawaVxfD59xrZ4d5WM2ufwcyjMmwblGO8mkehYFFxNjSFEiZyl
V/oEPzhnKnAdXGXZiWWxiz3a1vE2D4JArn/49Wc4i/ZNmbRxUGnAbJRDPAEk
tCVPopTS1hMfyyERlno8Klsf/LTsvpo0VfWk/UMih6YaNSpdmfrosq+EBTqf
UK6uMZedftOZgLA8dYyy+O+yJUIbSXC7nf+qWh8p65sL2JERexpbNV0Bhq3+
0T+va44W0cVrEqXS5MgSXk7f5K5lIRv2xubRvQIJhd30yZ7qpVE6ExZGRwq0
YTQzseG3LUfg8RH+1pKAKNHnWFszA6NlxD8FX9iCsxtAvACCUm69CE1ZMOy3
CL5v9lMf3JXZiy0XYsgEhyEfpYmRRMUw19IOZRme49wq1pCHeBXXpvgY9a1a
8+BlMPpTpsqlsZ2u2tL/HElGWpdpuQiPi9lvWfo5kT86av3ga1iaeioY6h1t
TN+o5sZJCUaZAwoz7GpRErgtLAs+vas3eVzD6YxBgcm7s7Wb6qB54R9l3hbr
RA9BIrj3Wi23BpipV4TQzOwGMBAORiq3stjtqodECX1O1VDbfNRlu8jCcbf7
KAGWK0PdI9PV/c4/VjemZfLws9bcg7SN8Xk5qLFV4DfI+DkvLe+RkcvyT50V
7l+2Z5ukmln1yj9KX9Yzi1ZbaZsPNgh+l5EyNq+77aNigOGHRcCp8kP8XLBi
UC7yWGDsffDnZJcip5D65LZh+wfRLFnXyoqjO4d0xlGeMTZ9w+8fHrrNkKEn
QUX0wYpqX0C1eE4kwLKVOzG/zU80lXUMDzOdLGBOw182ykfVJayaHCEFz1tS
JvgOK3uC2R8483b57vO9tLq8jW9pWsmybzToBqEYFLDOcE1a8BYAzNnHH02Y
HlKB/+eyU0K3gn7U/zqhjc03ZEwx/6yOsPFhSG5MVeJvOaRhR501XLfn9AVJ
nwYKwfM7w18kW33NhMH4SuDTWC2eOVbZrP0TLoA3x+v9UThgnnTHmpZ6V/vv
74ItyLbrBkzb9/9iDMP/8xJ7vRTQciB6jwRGQwQLtAP2V0apjYX/4cKJMlrZ
X1RdMlPiexZf0iRpYRcUSqVTFuMhC0Sd/+cqdmEcuzVjTiOIkocm/PKPuQ4U
gt950yu4N99EFNSDl6OUnbh6n7a34djTqOzRrE1EJl2V2xDLT76Q/J1c17Ou
/4X3kMghGaKeAs3flZEPEJ6B7jexT69Wja3hOUn2GvRHk07g2ZMyFJz1o8m6
HIqzWUnIQRqTvd7wlBr7QXGrnuPJrsXgwQ2L74vUcbiT6yYN+8ZTnujhXwSP
sv+1PqNb94USbXJVuYhfx2PyNC8ye7QdHcOHGFRl+rkZY96qBWfjg+4LSW1R
8Ak0c0NkPuY/WJHX4ajGgGE2DjqfZG1CK5juf/vvvG6oHb6S2wJHhGqxKIhO
0aj8adtWqTBn2LlBgvtCqt72uq2ou5PIdoLBBGusQMUA47s+3eE6p3dlRvBA
cGKZu4+mmvKhOqL4+PbebOXRLS1N9ly9/dW+kzzlq+S9iZNnXVS4MJOq7a8n
vTJyqIAjst15BSKvKbPY05neYjCbMrRjQ92eeXsVi+viwkUzXFkMnBODHWFm
B3Dmz+6d2h+9qZmCpTYmqxJx8LjU8zyjBOmVLTQ+9i2ojd6ohZ3DMbUjSAOI
Drjep9WQX7busfzHLaEZKTXKh8SBenJOPhvGRIQt5A+BjPHvrYXc5UkH/FRc
zkkeO+k1O3Oylw18ojGuRW02SkMVkjDEreZGIyx3qLPPcGp9COdRhsY6oYnr
/SlQhe7xR0t2K3MCfgLezYRRNMUqycHnbGjlY7UH0s+OIxaW8cujjgvcGY5P
hlJSO/D70zdfHiAB75uy6Kn+Aw5QKBkUUbSOFoLkX5VOW6x+LSWGZh3byKWR
KwCjC+hoCmT792/HmCWONdLvHI9aAzuuzfY1gcBbA9Zwvc/DSiwue3rQ9DcM
WlGhwvd/hGlJIEHkU1vLBV5Lgn3Q+tokhWRgrH0nn6kUoeAgukZ9Cwi8tsX1
FdFtpbvnVFQpT7/d+SYJ75cNF5rp4zRCMLnWs8kdUCQUf8Ys5EkdnweI/xwV
zsaejwepKieAJU25j6yOIIgqcypzVDQLxrLZVDK4ytCba58ZsBEB7BIxPRRw
qL6CavvNKn8nQ+CZudiIg5zYgcJGX6Qwd3zkDjFtMrKryX2d9Oc3ZcLyN+A1
yTncWXpKXsDnpAYOxQ8+gWfgzdXxzrWU8j8WqU8pwZpA7wUCnRc2XD+P2lJo
QiDZLCth/OpGx7r9FTTQQgajAhLaEqx8o+A8H1WG0wlW/v1WyCZS2p6HzDgf
uFCJIl/k7cLAueN3aEu5raFe/AkO2kv6TaJfCu5LWL7l204zBM9Xs2oyRV0m
S+vONG643TFZlyHpyIDwdbwtGZgmFTx6wViwL7ezT4LRMM6OZrYOxJlbvo4o
C/Mo0VoJdyGQoMRW0fQEbwPKmc+JV3Ul457fUsi9UxPpaTeHZ8YgFxey2lmU
/ayTi21s9WhUwAeGqT9ZgGvFk5bjEh+ZJmNZybVRiD+GYryz4xK8eVPHIDT0
pnjR6QrdQRhQ/s4xpE/i+ea1WIScRsS2C9KeGB/orFidLVzI5aU/1jtSbLpZ
Xq/pIVGdI1sTl0S7DJU02b/VJf9W+LKmBhurVyxSvWdxOUQKixW81PyagH7A
jcy7CYtLTkZlHMFvtjkoBjgrjTQtleb5O9AI0dbbJx8oxeustpgqgPZ50p0z
lAIw28wQjqUEglxwAcSEgi3SmZO5cquwH9NNkLtmAUhfwn8QHthwckVOy9Cn
sufe0PpPZnX3in1SLj83Y+Zybt94OrEOe9ymIHB+IN98n82p1LsbvATTLimf
XsbqICAEhJH9ZNiN7j0JOQkAGMT1GFRCdv41gFBDq6jpfhXN7bkXKl2w60/p
ZOoFFpvj2lHk4+hpHPycyFkppxquTNQJxkYYsKJGAHVzv5XRSDE6dHh1yY1n
4MThjm+NXluuHPUAnhwzr8MPucIBf+6Q4OY3aFcvTAPCJWs84QRswVsdfBBD
heDF+RYwFNNslu3Z9j5ctAeNkykYdA9zH3EwGgV0TM8UPWzZbH0DcPXLJA33
IAZbWUz3K6FtbO+1P3FcWIR4QzPYdJ8F4xICtL1Fpr2PNqdKQTyNPKxkSLNH
g9A1f8PhEcROHJYCubM37MrS4T3jdojY3x6CipHbEp/8GuoXpJCUwCO3y0V4
9ZSe6eiyk3YLWnvIhgZKA+usmjB5nm3FuV1m6gl3N8cUrF68YDQlH2uYLZap
WuwqWqt9lYcePU2+DXSu82muo+PAz3fgNeIWPayLxLjqxzrnpVfhOKF1B8ei
wUTN9x3Cp5RICERE/7NO5IjiQJlHdzt4ikeKCQqiRFk3cSWC3+i9pHaZwMgH
DGqUMwCU9yiW8dabziVcGyTi8NS5L5Z7NYjHxyPJgg5Xl4655sEWWrrPlsB3
Y3Fe4c0M6LqLa3uRDaPBkyufn8jgEF3DOvQh72z7VZxNLIrUNoUI4D8Ldc+A
rId2qxuQrvNpBX6h8O9t88c7b09D12Zf5z4NnqYIru2w6EW21KM6NNblQM8W
UDhABILvDKICzgQPqnQmAB5HtErwgb92CJEd9dc0E4GaFmXOZfFLArjQoX4g
0RgiRKkCuUFx/YosLBL3JPK47F6AJPC/ic+tbo7xZP1CoFGY99ucNGimtsRo
yJa6w6dqgR6QLCX/vecNGwTjoK0aYUwIlRv04x9i531UEJ/+y7ha4QQCPGXV
kIiUJ7ZzNRBfvNqU7pg7rvnEc/uVh05S9sokATbr4Iek8hYzhLKFLMBtvnV2
w+eL4xDcEag/oxVxhjt0R7KfXIKTpuvjFK2cC1lInjNG0HoellzRC7bxzp00
QBjI1h6rfy9tyyS+1/e79aqXR6PBqOpJ2gUQv0QlVtJ1JgtkNNMdEf7cuYsd
4QxcE911A3PnxtF1UyCHdH2e4GzsnAxGBcG7o9H4vfovb4zNmmQ+I3z5bt4e
EQVT6R1sUvV92aDjme1gNjlQ4O/+GQhIU8yYiJs0/5EULqdqn/teVdxEWdao
SRS7G3k+wsmggpMIcLWVMZL1jAU4y0rEPOKA1jqudbpCwjKofISxSqpavDUo
O4b0YfinEBWHyR3gkabdQXamSC4dcPDdXp0nmv/CT1LFEBMi4ZPboUUQG440
lCd47u5p1OXMoZJZNF0cVu9upEFUe8HgVe0M0E1eo/6ec7HdOfaygqBf8Rqy
FbjCrAIfXxQUz9Eqkz9NvYThHdeePsNVolST/Kp87obcM14k6cNIGd3Fttwx
y5wuxvH3/U86lvy6WKMqYd9OGzJHLVgeRYn3FdEWImtF870JdrkN6CDphUzp
YX8vVuaYDWc9h159GS1uN6KNt/zF1hccMtJLGCNDnBd93lc8YGLsVrdQCSjK
1GspVwsAlXAtF2iDyn7Nimx5Bc+sCfZWIywfKOIQi4ZC3ZDt4+JSn8JVZIgC
f0HnE3NQjhytWMg3fTk8f8c9qQgABRTAplRA65Z4Ayhctq4AqQwdxl+Isku/
5T99ATXyw/slx0DyWs8sLuy3wZ2ksq92EBybz4NIvDVDx7MHCTgUkfnU7UsB
zcbBz3SJSzKwfb/o8R8Y32FSuOfEq5nyaN8aHmocN1EHy/Iz8g5tp5hHP+rP
+uzy+ufv+jOnIgpNXGljTaRvT+eDL0vr6XNt9RNULbUWhrc8+HIkfxxX7cve
aK8ISXYtF4LoSI/hVbtgxFBhf2D1V0Bzok3SZaFdrDFFnCR+gV/CICTOuKb5
IParwwGJNXyNs6xZT4UPb/Q66qpI5khbTyFhlm+cTXUzeJd6NmvfSvpHZVZE
Nzj4HtA3K0Y/fJGKCV+QvPkzI45sPRJ5ddrXgiCI1gQf0DBCQb02620yFTKB
9UZ7Ko6d1F9EoDXmLoVqKbNDkjGQXeIJdDkIUV663UBqK7f9bBNwVFzYFV5i
v3Kzzlh6lxidyiEWLVRvynzx9GIRPwXdceSPle8rPSTt0v/qya425cUku8yV
lNXGcU8/AiqPiycZApVqzfxwgu1s/eaw9z50FLHfIFblTMHdHWlIC1KRKmlQ
OlG/CSQ24knFm7yRRmXwRAYBJ7x5Z16Qrg9F1K8J8FbZXftdudLVt4asbzm2
ntGrUb8bvEv6NM2uGQn1dGBC9ZlkBiX9OxXgD5jkTvCOx8wsaPSvRdbB6why
6dcR73wR2N00+vZMKaWGkGMH7qJN4WXd5GHjzysnNX7/ITsnIRPgxmMDhHVz
DjhTVDcXiq9lKxk/O/wgeTBJiyNjZmI5k5wuji5nq31imm2GvhnJ1anuF/b/
2s4bb0Ezbm64oz+xakj8u8b1X62hDLg/J4W+rKSkGDLRUcs/d+LeD5ZbNscz
So4340MDUTaUjvz5GLUlJRSPUeqHYZquscn6k5QXwVfbGchVYjdkwGiSVRd+
3vBCUd5fRvzva48Yctig5bXEbNB9RMFa3kekOVvoN1LCNxOVzhO1WZMCRq70
/sVKvduX9KsoQvWrfMHtx0l+EfUSFM5AX/7oeohVoZ+4Sq1jdw8WgyKSm0sg
LxAM/yKShZIa9fCijBNZQvZHh3dLPrXEFMwuZnBR0mKbrdCoNoUR0seiCMba
swAs1OudAak81tHj9tupQt9bnSyrBzoj9Z1TaCSCVvpX54g6KpWlIjD4v7uC
13upW4slk12M6r8a6vSE8yYPgwcyQfLmg50rh30qRdP/qx+oopl+5OSyH9Ke
9Lu5IvNKwxoQsYQyz9fTqxIJOFFQUXsSJ8Yctjh+z8mXMEA95OnM0mkwmK8M
W37cLQy+dFfLv+kRL9qNiCAZd+M7+ujM6Dg4yJdlI+W4htaBlMPzyyFq3SB8
Tu3Cm7G1LQqoKUZ83VFbfhpdeM07qzbWhrL0dYD+hFIW9QfOfgBNl9xPTVgE
jl4we+4qm09trOUqiUq3LOCicmR6Cbo3SGVHNbtDmGhdzbSwcUWoI0gwgJAY
iFVC1u1fMA375dQ9FSDfT/QZnwtrRbBDONeckoeG7JJOTRYEsIoGIfuyZAta
mZqo/KMtl5EBjyr0zLqUGoKgBKBfGECA5mxhDS+AHQwbEAd1DNwC3PU8MDxb
UD5W+TGBksYK/BUUaQNzn1nsDkm8S/9+WeySv1UjQ+nbDuvg7HD20M5wgZ3m
sWwsRZWO6SJHy/UiO8/W/+rbz4YZAaEv1/h7Xl/9b7pl4zKjH7MDtRU8FKFn
RfxEw8NGi40O9VbgNN+MCltxdVpcOiUWo3FLWLazLjC7+FdNpUs+BHLZ4a5J
Pfx/bN1eKFSG9gNqqHtK9/01G2IJMRD50IHE//qFlZO0u43NgRqIWb+ymb6/
HjxVHh0fIt1/6XZ92QrH3BhF+gxp4O3XWZmqlL63sDi5O66azLL2vyg3WZZc
LwuVGvw9oKa6Wm0QMZapHTgQ6mhclUhbOl2NSxH/NPgAMQtlrcdaXk4fqXEg
nSPgI92iI8xmziz/aqpBL9KKQGyPVDuALqbd+a+O+DJNpt6YjFvfUImvyBnZ
cLI24OIeT72c/q/jahdHUc9MDl5tif4GWaK3UVXCcJ8EegrIfir+YdnmmsBq
46XkqzgMfB9Oqy+EA4uMOCWcKcpzoziGB8AekXi9yu1evot2y036zSUpD4K4
Z0kG7jimC0z11MN5N5z5vuJzkW77WWa1UIdf3kyZU/Zpk3XxP17d3/+bHcMt
paMaVn4xcXtiseZgQ+Phyl2viXfOh1Rpg++iJa5dF2MPtx5weryZvxBY7+xD
dtFVjrvwMCT5YS6z/GUdHmwYc5Wan47UqfZzofPI9DFQVkV/rjI2CkopYgUZ
jwbr8k/PUFvrJzPajfko11KxzBAFErw8XoY6FbBO37aFcaXatoULLa/Cwb2H
9/8sqbRGJZhVIy6wRrPnAQr4Ka1J5dNFW27UsN9Y/LEO0HFkiIw6LxmCqpcE
AlFM8yOz2kKdPw3a+3aOu3n6h+yNsfay6u7mE8XxEIzPRsUMgM3a4qQyRKpv
4wZ1avK6HHwX7qh3NhnHfNmbmM440MYQf0G7nCt+X1IDU0vrukXM5TTF+dlP
fpqafwLuEkohhpfrhXW3w+ymZmJuSfPNG2iYRhPo0gfY5r8XJTSuMvvy+tPJ
taFfjuRigecuG+A96c6Ekp1CP1nYogt1wqpnb04VGTg/62U8Egfp+2I89kw7
7+MrpZXUUSG6VS2+y+WnK+aNbNkhLEY7Ose7yRHjrzVEVT/xsOoTYe9n09ID
kocDdNHrwGM4sf32LHsPtQFZ3hcrC3oCm3BS5rmxSAy3fIc3WFHUeWvJya0R
xzr6YZAeJ19IwroTJKoXctDhpo4JHzAYnWnunDaaBjp3PLmcDn/SENHV/hrS
vefL09Uh5H/ZmqR0tdwFN4odmFBlEu6Km5Bo8poarnbz+gESVd7mJNmikatq
EWYXUWQ8X8dw/SfvO2UkXO7A4NXNPqhifiVMKxn7Luwh9H4m2/X5R9qpqguV
vBITPvuXXBYaitgeq9GFJxvR7lC5hV3ftd9C2G56CAGVTxWpsJSKTi9vPMOj
CugfxrNd7QE+W3T6jOkzvlg+IMiu+z3SrRXoXeXKQp4rAD/LmjQsQk4RU9K+
6aoDS71g6TFNVdDr6Vtqa7kFNBQRu1vx4BngNrKC2FNfc2YwJ2FeP4270BUo
vufxLYs/kplqIZx+3Gdu2zRDhX3DRGCWflW2tHZLty4kqhsESrwS3wL8GhsS
qAPlNXjfr/Au2lfp1PtDPBQVjHdc6pU++ncjfW6fF7vchrF/AoD3yfb1+HQc
KevOsRBhgpPCaGm4d1OU8QSo++VHqfwpMV+oi0/DkWGbiFxGRqemIdJoXYx8
hd003C5ibOydBl7UzGNq5r1wJWAdv5dlZTyHnjqki8h0hQ7kdq40OUaY3/2b
ng/pTwGLodSVogtMDTplOLsb8Q6NKg1DVX9JV+/Fz7l5Q9VUCvnPs8RA8ORx
0dSVUJ/r8XRAs1orT95/sB60Tc9hCsojFDFzkRpj5aLUlShHknSy4uYE6P78
Op7pfJSShMSO3yJ9gSoPVaJvCsKNKgEQlmhhBmquVj4dl5M1AX5eft4ycQL/
tEY2y/NK2v22RwmeG0T5GfmQQtxquzEJ3nJpnL4VmGIt1zrdEbjQ+0uMBPY8
bLNGPd6FeZRpJSesSlEjZLy6/5WeiCFbve1x2KuovTZi9AOo1b0ukFX0t4nX
CEjGNwTbEbn7s7bvoswtlu5BTIXlfYFKlGDpL1R+PwB9S3AYPjdCuJEU05Lc
1FNXFVBb8DLTmLl44zARGwjtgVYXldA92JF7DVAFhZetGbtgpUV1Fd1wnHRo
jzPzRYiomRzqcqPKyPT82IOJbrLXJjRCWRW4fZE3nxngL3KNz6z0BEnQBVpt
rBEfP6wF0o7uVvX5E/1QHyjfVW7x/mA6WxFFxjmscGJ/S6NeeJfMyaiPqJQy
jdWznHeEwivkD+jkv2Dn4aaHzJwnp5ZFIPbEp+59RIGZ+Egu5p7j5T189Tzu
NWh1LTSrER4IU8wauyqzJnxMTWt3V+dm32aIe74krsZNMer92FSVJuYDpXkR
csCXQZgKJtQ51A9QOAffN9jx9O7hB/kBaKZ7veyi6UpDg0UXY3+qE6Oz206r
xBBq7p607YIGPPUYuwIYkFchRzEQ9qjUHR9tqd5b4QB4J+7hQ6zXO2XyRKLI
8nCzJG8zRbvjKZR+s8qcKP+rQiSDYxRjX8ASp32UadS2EKfgjeIOpki7/rKd
6fuFjm10MxU6p0UnqTasRQtn2KaTcHzoYM2+ZoKYs9cYXcaLo/5JfmHTDCyR
Ld9X4JqJzvZq0ELYtRu9sA9JRmcoQyNuyxr5y+sz6MCFMHOFa0c21MyO9JPo
iDURUncHM36V1b1Uf9vdGAncsu5qMaSfBxk9NqsixAzFokBF6ac2wS3ir0ya
vnv/znBe+4jn6nANTwaqsC9jZvJpdO6uenwXFmTnZCIYYVznhIsV5u4596qB
oB+F/bIIke1psYlWOY6V2OPJCVzrAdO7EQFmYvzTc55E1ZdHyjIfu4h709q1
Bmytqq8Id7FfTvWJ0C7FHOlp5vordD4+e/0jXzsO892uQKv1U7xXgIHQ79m4
AzP1lTdCqLOObrHY8XnGU+jBAcaRfTcoX/qUV/v0sW3aEoYosFEDoWB0kdZl
rJ6U+fYN7ZqlLDTNAskzXuh1hUwdWwWQqS1Esk1Bn+Y01lFbJYQh1jEDRIa5
/RZr0akJGDBxi5KyxXE1lpBubLTg3z7dMBq094rAqWDStr4l+iOKdl+cy5He
h8jxShNke24QJf79/Q0lLgWPlOEkb9gkBc0aWTBB9FaE00vbCCgig7x9z/xF
4iWHOyxcDkSFhVAfecd0FWQy3glUycH14f+sg1H/b5BBpycB2FUb7ABCdSSs
ixKdhrRfb5cM4a+9vWRVAPCFnbN4nbSQlZIXT71DbrZe+0Y3iHtrP33Go9d+
JdyRjnbXvzJLROG2m+Eclnt6rRK2mEIEc47jQUnuNKhc5gDlKAmcvIijxpvM
rkXVItltI+Yk5exEQN9NMzzCo1weW1W7k/DRoaa9J3C4Nh6dzqKVqaGrNyB6
8hiCMBLyD863Cc3gi39Uyd+/BJqu4brOoc/jZ2kIdiimOulTp1DMtZ1lJkcG
ESA8Xj+drN0lG+W9WmQuMiuADXfqzcsiIi7vf7ZSSM2Dq/EHlBOFrxStbzbA
WMMAlWk8R0EZ63CW/Z4OGac3Xrqo2andh3g+1K2HvdKneG7z9nw8TMwaFurc
oIFcEE5hZ6hV8bzOygEYxUYjv5Mdt46febcetJFXaQQ/q77IZMpJ4hEruVMv
p7YYbKS/BC6qtoScNR1L8gKQF/YZ8/iYvyrS9MOw9bstRi81Z8Y7vEeB9Ib+
FsP/3yICgn67vf4saToZmws8i5TaPdHp6kOPqQwhm+FKEOERnASPzQJ96xup
e3trfvdiUQdzGjD4QmbqysFy7lWOfFbeh3hAtj2t0awBk6vuAUZ2FBNqeNRJ
+y0w9k/Qg8FZmIummJYUmT34gIXiCNN6WMuiC8E3DC/TUUFV6+pbBV38LzzJ
n0iNm3otwo3bHcqt5fQIORu0tB/uR9K7LnYVw5BSDSVzt6oHEhfkn8F4cDPD
9hBYgmLtAmB5I5Pz2JsN8sNTeoyanbPh+G7EQKDCLCdXDNd87B2GlCrbOvr4
diOe8Nt2O3P7/QZH4byjz7M06ZmQCyEtbGbZ9rjem6XtzsMhwccnhTzyi7Xz
0O3FjsLI9Pcb+xkGcdjT5DuH9mxWhseifJdEYuA+HqTvGdoOXXz7x5jmC571
PzGacgL/sPkTOMNQ1PPAzaqyvDilx/tuO4PmQB+X1B0oRJ6F0gCvXddDLM40
TOJKjHU2Cew194ftm16evDKiT3FeCw1eAnSEuX5n4l+eqAovrg9HKAaeUHOy
V6C+mj/XLR9fSOa65vmBT5rvJbBLUQi1hmzEQ/XvLbPVr3lSNXMLaWJZUYfi
6mIiclvODQpFpwjgNhhASX/pijU8FBGh2GJAX5vbZ9M2U/tMzP1/efRdRQnC
DJNxDMh6VN++6+ZdMOjqZh/sBntEOxXx6OyK6MYu3i45UOtvSwDGiYGJuZMC
4nwrJeactc9dgrc7FT9AuA+tx/1CoH0LVPEDMtRW0MONh56jdC1n7FLJMNxy
ZlXb142ORiwfRyY7PTwHFnS0KhyijCHWHja8hX1vvlfZcdqA4Qb4vpW1f0Ts
yv14Xls9TacOWqpmkwXSzjVNNIV1MWI0PaKzU7CNijiWAhtYb6+QttIUUMoP
7hnMwtvQIUDtyipG5Ua8D8o2ubthMh3zD9HIqUSQviE+7AO8ryKp+CYvey0h
DvCVNKx5nNwInBK2NaVpEsnI0z1WvnzCtrV6t1YrUtdl9A9qURJw/COErsHm
uAUl6zYBKQe7HMJGRs34DQYKhSP1PUQ+c1XoL/1l2KJ99iwtGCg1T2Yr2skZ
1wdRBIAPYH+c7KZF6gD4vk5ldl+BFCl9DoGZqiAT1XhsQmOCxANkrBcRObnX
oSw50zgDZUEF9lShKCMu+H6n8XdN95RDFWMOwF818uPbZuoHGANsif1Uuq5K
ObZWdrLo73s+VeAx257tnI3JdHNLn/wlA9jL3nAFcC9FxsqIA0aEzz3xAe5J
VEUEkLfZGijRSnRW8FnHArQTWM0N3j3D9Ck75awTo+FOfZcighxAyvK0CYe/
6XIziLgqfzkq65Rfa6czQNWVTdKYqRQYrV3luXmiyEknPnVGMCKwjB0gt9oj
i17sr4HtaQ6hxaxrBicmRUJnmHwdZdPupwPZ05W9rNo0V3bijn9TGg9JW6Lq
iHhJdzmsHyOpPxjfum/w1DrPiE/MezjIA5XRtvlCeH6n7Qp0D3eWhYb/2QNX
f/YZ71q64/533QLcpWJqDZl1sUz7XWbd1ecMVx3GB6hLjNxfvQL04sQTikQe
epkS6YN5UsHZKkEsWFB4k/v/K/hQiZJrRIyrdYD1ys9Viadm6c8rWJy0ULWb
QMy7NctLadq4XWMQ8Ay2HTQIdCF82C94Q1unqPqQdepEqGz8wOEOPFw7EujJ
zMU+uvvDTsIjPOX8u4UFqNwMwTaZ+uL+8MCQRcQf7J64dJXOOqyY3vwTcAOy
16KQtD6oigYSoIc1TbzzbBUaSYLbwGOvlmsMrS5r9gZwijuXRvE+A7tIJ/QI
yOwNt6mqAle/4+t30BnsbJUsudaBMkha9JeIzJwpS5nv6/69nFED2fMP45fO
QLTbh+OhV5wCKp48K5wzJrdTpZB5Na/52z6dtw+GnLfpy96yVPyhyoF4OrdO
MQ08kNTMQFv4v+Zx0i4ACHIUWj31Xu/QDAUNcxI59YNDF5WvnP0zGaOJ0iwR
+iq32mCjNRFjdAlIcOABHe1VnO6p14bfIPZgKGcNojPT+WkF+vU5+GEyjY+6
9yF9XODhPAcfCcXk+pYFknitePSSdpUJnl5Untnd4PyuMsxAqLWLlEsnxEPh
AuHmfreLOY9feiaOCD12GJUekGLX5wSVCyHS1zi98idvRleChb6MV/KTlX68
yMbxsMTRvMPGko4a5UbZwNSFG/Jy7GeQaPvOTxt/iGljoCSMqpDvfpi0WnAD
Ez30PcTgNijqDUG9RTuq+lXVUG0xeQAWoRcuFChjovVoaPRty760TejPZz88
HmvxgwvBv1kbMw2+Yvte4qdDRpk9f7FrX24q8cP9Tt8tWwwJHXX/Mx0Y/mTm
b4Am/b1hNcuq5uIiN5z5Njs7OkTKyS6stIcD0HDblLHj4VgKkOamz9IBIYiM
N4lsgXXIXCAZQcpGEodYg2i6SF6EyzA7PxuYSemLpaM1tEWo3dXxH2weHA1s
oiKFDm7KZ6YgISfyIh/y/Eesqn1AplpGSkkEownOn/gmWrgUCrAy+/P1g/kh
P0tozsQAta47ZgAR8io2NhR3OcMUPkd5JrwDZFj0lbPhxz/5ZGg8cSR2Ao31
VL+OQ3wqlS+Bfht+9LbFx3dZGUfKTe0hHo95TdpnAEfyNVJG8tyTZhnPfePD
5uAI5n6Lv2ZRAIbMpFF6SE1wEOyDZ4STZiOP8BqhCxzd4ej0Y6FVLSKJEzJC
I+90ZE9A4SbUKsALT7R1gm4u2co4Fop+eGemz5itT/m9dx2d7Nldt9NFsHB1
Qij2GsWSBqT/y7DV8ySedTEinN4atLoXc3Q9+EP4sUG9IyBws8BNL22hqFqb
/5lbOgorr6iA9zh1H9nq5S8ph+p5yBEV/xVILBl5zIflyZf/lTKRkntzSsXp
4ZQMODk9lCu+YvAIA5HSjfbyNX+Pb/BTsvhK2+93R/K1+ynuBVVQZj0GWw9k
nu4QVI+jvrWpJ6BsGR9DC++T/dASFqySEmoff74lfJSwpAtP9hKEqDxxbnVG
Zc48laCvdW6OWxy8FV9nAQfqPTci3rlKK0udfZRjKguGSjR5Shtft9dRUNGR
wElatyKDn8zkSaYcHfyYFZsglxLf376w0SQ/pjE93TihoJinu1NJETzrXXgQ
VMFfdPXwuVv0BtJ3OEogO8k+O1IcSe5EZfW+NIp7BXIJ08jaS02A2//4QjNw
h9VjdcQ2rCxwtuUdvUE/mqxlf1BZBm4lu+EzL1j4HT1AaPExnHyu/LurnEOG
zU7OjcCJvRiA5DACZpS/wpkJ1g2HpHpN9k3ZibSDSS5g4KUPFlQH25gnCkYo
cMMq0zgim/S3rOdvvs2lUS38hppJIoO3f/krABaw9wElUmskJXIvAB3A49XS
dpDYbRwiESnHE+N4b6ZbmZZmbVt3jOt/H0JZE+3gy6R4ryj+O3wId5D7AYoy
bNHoJeXCxMpa0VqgJRqKW90l6MOsOFGP+cDQMvAsROW/ejBEMWfOmk8TtDn5
0RUWvrGabD0KVfQJpYoDGVzHUvZXmiuFRYHdylVgl5MdZ2HV9vwt1oN5qBT7
oNQuF5rO+0LGqoOoHHELezwQFh/GCoNoLQwjeT3IKMLFJYDVg3/2WYYBTaMQ
HJvZvJacOX/xKKzVPpLn/TtKWAWo2jJo17U6bl2W3i2FCvlIkPYJ6knSkCNm
gn0/vdz8g2Aebhy1jEOltbKG4nX3wJHhk/Q0BlYyqlwwc1wfmw6MbPlFfIkW
2+9+7XEYyN5QrKgyf2IwmGYna0JP/zHEEG1DDNg8VFJ45K7aWLwAvY0HR0Z+
UOQGrtKEO4eZBYNDsJvAl4at8U9exE1SNZ8ARi2cx6fsLyoRjgST6zaiCoH0
IPfwzsgcQLTKeLFtrft6p/gBbLtBK+lSXKpJjJFZp9UZbaNHSL6bPKywh+iD
+8zXHWztkOcQwt0AWcd6QexqDG3OflTQ1EiQpFBuBETEthI8hHx4jC9ZzKnj
7XNtUMhoNKw34/uyeJUU/cb1WDo4GTwBSWmmeYHkK1pkyiV+LVAmKr+a01hA
e3IuKX1B9gB32lxQ6erGkp+Ze/fSROoIxyHHFXzkvrEkR6AkxABotsberFhk
httZklXpXzG09PAvxDsT5HYYODzFrQX9duosMjcVyVZD36p7YUeRYy1yxjHU
FBl6jgxSGi2dKg3sZ0X4jsmSHelpLDC3+2c3kMKfyxJOKpgd47a/NpKiHboJ
CUdMWNSlL14wefxrO5sE7HctnGMlICeL3BF+AjpLgNdgu9eKDO58VcpEqNnN
u3UzZgO2gRrsvs0bGM3MnOL8Hwk/JlMc56XoQKVHV6oUbUGfOMk/f15XOd59
zQ0qEiNtZZpBlzmhLT/8zc9Y12v8ENg0d+KylsFmkFaQ640d1E7ALWSZlvfw
vNUI212arAy8caMVDFEhewu2vJgwrIZLJ6Da9o9s12I9wiTZvvcf+acet1xb
PHUV+aiKXalw+1AmQeiSWNUnrnBaR0OolpE6uW6papfwuKWEfXDKsZ+AyRe+
YROVY3gzWELyzsZbe41VG+PZ5KjdXp3h7MGYqedOW+pHEmK5VJetvlIB8Ir2
9dL/9x9aFilkgHGQtYJonA0OFfR3tp1g2jx4eapZ3PmHJoKAJI+USuiKmEwD
Kj1G3ZwLBDw0QoCkGgj4Mu2SzZgmJek8xiZMbs7ikMbFLUjPsX8eBDWE3VT9
cOh5QVvDqLseki1CudWPliGceELM+42MGt5tNsrxF/dVsmmvxgkcZdczEbbz
7C284VpDzoJEiSszNGx27gi53vmynsZdQP/spgn26BF+vSc/jluFxSfh1daN
4aI1VhoAbOSuUtEdvMO9y6Xnq9ZhTzUHHEUX2TIXP6i8JBqyeh7koprdslTV
lbPgZXHMYgCqmWlzqzydpmwFIuA+dFWmy/Gay2ZFnan/n6+qCi6BQfSN3wW9
1hKF5efgFTGmey4MvtRAxxYPQaLI9k+OdqP23YHql9MYrQhru76zUuJsRoL5
ljZFRMWHeIrpZy4vd9HkQyI0y0VLWZ4HldwzZr5B3mzYtQ1tGwWKS12X7ccQ
JS/mPfkVuMOKhVfWeKF9fvJ13Gi4iAyF6akvCDGpHTbhe2k+zzJY9xOUw/WG
mkc1e23UJoZNYX5OGV+MUVhIKfdH8UoV0oItsaOGNJc4QT7L2a2Mnka2EW5v
F16j2VYEqfaQnF7AMKXDpXYUPZ8Bx7OtXg8m4fmkzpr564O/AyP5a1N5qjq1
0s/M2olDsTkZMOfQzlF07KPnMf34zwrmMG4P80NyLCID6ckDKj6XT3rABFAf
JGMqsrkbK8BwOssM0KZRLFN6ZYBuFDdG1BbyhWQZT+GfQvWMaO1bexlIiThx
PU17enJ5sAIBWOO4pKxuz9KkxNmpRVU2qAhrpbRNfZtK6zgn2g+a5dN4hmDK
qUAl/ZrOPZgLFEpGCwODfUwK+WbgYnHZP9EJEvsIORS1Mpo3PSNJXeUQNhsO
ML7XQUeuHna24U/2stdLcPcq0dnkS64vF4c/lDNLQvopBgKe7sfqT1mr/J6N
dWlTMAvVPar7hP7nmfimfNskUUYgpDsNORZ77cx1wPp6W987eIJ4EvKpKwgH
iPOgHBOA6OcM/2SxtuR8SzU/naxJ1w/Mr5byCPrzGA3yN+bISNPi4vGwoEuR
NtK+L5o3sd0e3uw+YO6SXsPXJxZuaulxI6+9BYTzdI7iJF7Ble1o3CxFFiIN
dpBNjcQ+H2DmOhTL6jY7vHwxBy4sF9dxOwc094H3awvYIZxTC8utMIMny/Qo
OruotKUT/3t0bn1dpM3F/xF8twrCt8LMAX5yiSD6adSZlWo00Oqyrd6783gM
D/RwkzOE8TuSMhI0+jOcPmx9Pl9o+cL1ken/pITG9lRQbWO1tbpx8Mp6woGj
JsowfkOQrafWTIb7v2sYMFnXJeksX7R7zZlyy3LXC2k2DrF27CFRp6xVbp2C
ovlN9lnrQkfFSf94JY9fwrIe5Yikc4Wug05V90EGtxmRxYJK2uhHDpKLC/j0
4kZQTteMGv+6VJPvHNc0xPmgxtwVgDG2V755tJjiPtnMLlZJthDzK9B+qr7J
9XA2+0TfT56SflT54JsceABVmYQVDGOTW4uwvHiJmfztWXiA2zHt2rpo7trC
rp8cpUeeVAxvA5eVhsbYT1q394BPftxSlNAnP0YRsXiUQ9FwpkT2ftBxI/Pa
ylR837IWvXdPmoj23Wv7TW9A21CzW/y2msjSfc8iRg6L9d18zLxn4iHVlf5R
2e2ZgtAz9ZFaHU6cAu5AWjsHur/hMCQ2k1oWzUPgqn9bzlTSnVfn2uIkXCnI
I+897wVwDloZ4KisexQz4PyhUP8kKJNa3lQ/94BvtPaRtid01cIBnScR1Yyr
IiFtfFeRfvbErbQJTSuHpSIg4tjARW8SQD12nvmYYYFaydjqNZFWc/F7zFuS
Xu8BwNaSIyRpW7ATeTw8TonMynIgaAzFMkYYHRWoj8AOJkWvu4JuHdWNbTRD
JmW7eItrh6sBTg4/RGgKInqx9bf/JocKR56N5sWQw5ZUuVoLhiYZKVxNrhWT
wU6zdz0moJxA/+FAX+Jr4XcwA0pLcEX4QLmsJDJMnhpM8leZf7sUQX1TgmFM
7lzNJX2iS/KDwie48z8DTEv/iR8js1loM1RvhHQK3YYiCQj7DwrZKhbi9kUZ
TOCN2HJXmt65exO31BrchkYI2peFOQ1Mi3ZrBHQkIDv9ELCiekZkHKAoPBRP
/sdgybidfHDEckNA+tv11yEUv3xFfdSOf8B/HOQa0HVSc1M5pNnMGd5g5+DJ
eFVEUjGsNgDDuw401YxV8/9XmftvUX/sb+aINhaqQd/5fRfyVsCwfzAlv8nI
lnxOvvhs2m4RIplD5Bzpd4esxKxvwfrzZyFczy2e+EO1NFHWGTmKa/cJ/eIm
Atzc7Mf2Xb1ujzpH8QWc2bYk55iTQnyIpiV24jZjSjaHYm20WaHJpo11/E0a
2EpZopteHSa7gzjZqqGN47nh3XiNijhWQXd/JLDK6I8HeSPH1vWXx070TnGE
vcuBX48Jv/H96UQlT0k+WoUdXM2TTE3+4X3RwKbSMKKggtvfRrNLNfbvjsdL
M166mihnqL/op015y6gCbY7q9AwDrj22ZZDl8OBYQQb+VL3PbYm4SlH/tJ3V
e9K58eJB9rOwJyxZAqbZ6nOjb+jnMJfUeSZhbFfQmu8oXIC43QI5MZ5Uk+vZ
dEsMJiD8HuGzjdBZ8GollZdpqvv1+eLZTWLX44nTJ8IUXm9jXpbRyk3ONvid
Dyf4jQgq/XhdoSVXZPbBATplgSgBJ8OiCsm6lkDyjHT2Ddg6g9PvSQbeJJw5
wvXi9UZh74GVqoFy3vYgQbmmrG2jx+YqVZqwFGt3BmDQW3kALgzqjVCtcSkD
1ZoMtBJe5/ACuwUfB0AYSERD0Oqa5jq4LO9RpN2eBT4cO2X8WzXYemK0fyT5
niAJWSXSMomRJsdIi821lL//CN6mvfPHYYrjBr/bHFElDKUx1AUNG9w6e07C
1QQ8g+kVNwgZF3cmvJD0hCnHtN3gUb0QmNVy2WqHguJMqFGMLr1J37YSkpNG
AmqjxPcH1acHjHDSbq1xTHvyk25AWLgYKOzusOfykOzP/PTBc6BcTZ+EoN8O
AhsKZmpA6gT/fFwO+hPuACMfT3iHibQS6n4PdJPGb5/CGIRUypnzq0RLDY4/
XsuKJDjLldt2yQprlCDcjijg2L7mn3RrZbdm6XkeDVFigqgLI+aP99mN+zKt
umJhOXeMrScyh9TUtRGwlcrMcRp/isi+BMCSeb2oTCRNZ0oV8AfRyyKm5pK9
FVRKiSMNhi3ge02N3PRJKgbZ0PO5QSUFFWwNZYevXzQNWvVMA0elyXv/BeFq
Uzvzbu7S/yyJuPHYw7xs9tZJA1H95UI9GhkMHszSbMFM+qrLyejJUGwBm2fI
kfJhChFqLKhrHlppHhIRwU2dPZp0fFwbLwH1lRo1/lLt8BjBDZXKf5zK3CcS
OR7oGgl71Hl4AlUk0JpzFEXTQR+hs9vwBbN065E8dwJ97cn1pbVGHy/vQBlE
6/MBZ2GeirDCkbjjOU/UlA5RJEXlJxQ9qZAm1PtKOOSuQVU3S0WeZt2eCC6U
NuG16LcDcvnh1+kBt+zJK0+SBkj4fUSyW7S5E3BEKJkyiAtHlgwTtvAtE8Gi
oy+FI6SjWw+XNYGV58K1L69GDpDI4/Jj96jVy8h36/dTsA+t2qUL27M5ZCVS
DylCVQYNiQfLbb5j18+YGkygRgPLBiG+Dbf04zccZe6JGMpSHQixG9Sc8YnJ
hbNQT0Bhw/aR6w+v/7ci+QGGdonY3XUz4cZYS+bYlkIsWA8cjSoG/4lVszjj
1IStgIVkc+5o53/4h5ZU44J1SnF8nqrqbeL3iAMyoIWfYCYyjxVQwnoICHWU
oeZwkhdIcoxFcCYgVu98aanRXLShDSmds/gBzsitBLt70Ulb2VyRRQ2VItoS
cV3qvZXy4cm+dVioM3kllUFe8GZLn1OsaVn/qFvmhqeiIP/fK/+CwNxiI+eZ
oYgBYPPijBXF6diCWb25u+AvzhqtXXQdZpfmOfcXBJc/UylHSADneWfjzPYz
sATrPTIXZIcalvmrAcUfGqS8b2j2/QeuasLL08HH7f1d17+kbpR9pTUuo8WB
jcwwotQRreciBshxNAoTFjTHVrggutdtI0TYe/7xgky3r5rEwOOiTlLuiyRH
mby5lw450iY8mH4mhd49oXBmcUfCEh7sl0Vt9eDbRwS9ggK8f8rI5CNBOBpP
GQiIVunx+9bSHIJceT2vXWN6ydi7tWpk2G1NewPhpqc3RvnvlI1SH5HHJwPD
DkWv3saIOQ0kzVItGmARNvNM4a/lDNwbFgzduBwKcS5awNxxuUxFYYxuBraR
0w2nbryqRRVLUp81fchjYzQN3pQmXmZDoBfETEmcWTBb0U+SmR95WCPxZc06
f11oSyIzTAlj2sFEfVlNZ4KhrmfSGAZIp/+vdoob6x5TEVUk4pw98KDJ4BtM
c5KMLjTJa2mHNYUDGImI2lIcGFD+ou1eIynINpZrSOqAWtuGSZHcuNqLZlgX
CBxPIpQecNmfFSMxZa685dZghGJo3XuismUZAE2zmk9RJJS77HTI74mQTxiC
51TcY0f1NQymsTHvV/wCK6WbyhRaZqWnXRT6GLtjATwQtkgLVYhbt7ASkyQK
QD7SnEjot9bPCvEKW+8K16l7PA6YPew9FFNjNaT5ZMi9SA/i0YsSTTk39D09
07xsE6F8qmBRQT/IAUjJbYDbrYwLMbngmxM8OqmLzukRTRWFbjWSuyUMvVbh
pet/Zf6ZNv9pgBUwXTq65R7/QzCJocwFyu2q6Cqe5/kelK8y11VZXrZOP2/T
42hgc3SkDloDHpWp8JfXXx2al7xZk6fSCHNd/KtxgrbnH8/KCTxymqttEhy7
OH+0UTX9UZt2cweLZDWxwmfvajXcevOqtSzDUrbZFBPbcIbywnbiHsw8I59q
CrVKhfZu7WMOy2gpf2rQJ3kIkHvCARo0Rqm2AWa7XS9hiqGxpElVpb1pwHqw
/3/uMji1rrrIzPOnJsnjElBWDYMPuCSC4tqJIWMAzQTNXIxg7Jls3q/wAx1n
wqrUWP/5n9NvhQU4nt6p1hleYlRC9MWlWePH6aBWGnS6JQ1mgRgswIziBVTF
IL2DovjYemDQuHDwT4XpBuj6NkJc82LE0i33aS0MrPl6upKGgS8QdSNEThoq
GzbsLZC7ZL6Bc1+U4U4el2/oJeLhMGbfZsB8l4b287c0WdrKF2kCLgJDTw/a
yd1FAz4V/cGjrCBg5cYqubuLgQAlzW2h2bIzFHkbCkArPjJIwkm6TiVBveNM
zvzjpH6jGfTizuInUswNWcBPwMhHqzbVG/krvbcZBxJB4p2IebMK9PpnJs2M
QUUqBHp6kYzTCFvOJJt7XoT5Q/1XwUKq6zYQCrC/3lQdD51hQQT/agNJKGre
RLyckNTUA/uHW+V6Zn0nbVdCHMORlJ5lLxb9F5kUI5+sw+E5/6YRXp9F3vXM
kFQoNKSwsz72VJzX8CYuPr/aMD8GBvWR+rwKw1hkBK7J9BcnnLlcgsGYYN4W
rNHpri9iCi6MuO334TddLXTm9WSZggeCiL8OKUkCBWplMmUKz2FR/+BQme4G
spZzo9utfsdog7mFG9xS2LW2dLTYJ51hsfRDzFH5gL+m0l8/N590tT5kE1YJ
VcD+QSl7z21iGFTYKQ1O7fHMQyMs0PSf9TDk8wbUBvwbfgicK5WQJVonBoA4
rlhn05BIVO80JvolublkMsWxbCCY4TmLhDEB3up9sfFriY2QDMRzgQ7zN2w+
pvqSQ8TFzFS0g6DSSzIhq/hDBMTqbcQLntRlxBy3fmLG/4zhr2BUd4Kb0G+h
RH3nhpOdp8vOuhCwwuvpaJeV67UMdnKN8kqTXq4NHtXot039u6W1KZZiFmM4
QkUSowmtdfejHEEr59HW5lbs1+KsxKx4PpJb2jSDGYV2KVp/W67yWWuszx5t
3oja8KAE7iQ/RCTuMxpRmtPR1G/wuBTUihqFelKTnIDJlfmJ0uLwKezSuCQN
hPhDGRjsPF6DXj0ajOKwsbzK+vbVx4SGlCJTGEzxk0FuOAsRENq7MIUDTOXF
vFr9q2/xQ5bj4N5gUhR/lp48aELF2tialfpan8VwfBfgPPqFQ84W0CYluYL5
FGPyDDOz1YC+QGVLBibgHFYFex5qOC/Tfd2sk71L8d/AMjtZv7DXU7WgqK+W
uh6xre3pwIJXf9M8J/s2h9OMZatVn49hYybc4A5pK6Ok8H+YrXNyAv4ELDQ5
9pzhjP87Z8muZPdBfSVm32KoJcHlYcXEm5vmmGSwLYJwZM222p042DM5PLEn
ZFiqhALOLlCzUsUum1V5ltE8PJTY6hnLBhyq3K8pJjPuSLJJvdx+uB1xPrM5
bFMN+F4vJPUHTLHZ1tisYMYAWgMoENBZlAuVDKYMaG2E0sIjDLPp0KFBAdOC
3YT+6c7eYfshUsyBHI7SrpSmeEyQXMYPJmruoi3Aonz6j4H/R4xs0+l6+Lic
1DbkngjBI8lB2qmSw8iAe8sKjrF6Y/yMqdAYMUJajNKq88Afd2b1CPsafFGu
1p2c2UTUtiPVBKOFG/iIFg1nX8JfdJ89rbjnm3thURCidoREJqBxxL+dEdBo
ykDE3J29KEfYypeSAwvF7QSR0o8pNS/49+R1A4LzU05PPTwFUcRY6h+VTp1T
PYNK4nuFA9aCJYBd82ihjPY4fCNwHaOGtXuXi0GkvH3XJfpKCCoQlIi98q/V
wvDuQ0TSqrKEgR0tCNPCLxcKPCuIvxVwKYJdL32wd0zVTZCMovDuz1MPwvni
mihYMbmW5WkUp5uDD0D3ydjdjiKEHL6QeA4QZQm0KpAsAgQ1up6ouk7fZlqE
1rxmyxJKhO5Yeasm7ohNttJgFxx6J2hRyTwOlGhkbDbhABqSsAvlZyGSgXnb
wXSdgSULHT+zDAQwhe06dDT68/BnSuB+6Ni5LkTf2dEgYbINRNkQPsSPku71
kpkqeHMNd3lGyT2NG2zbSWn+qifSLgC2LodplHc+GUPaKf72Pz04bit8LJqn
zvkNIzqqO8MA4gAxRf6cUTujkSlihq4D56/BBUwkD9/qBBtvv32+9zuh/3uf
fvDiO36n1Ow5VgkQ97ma/TqdsSIaP4gQlstZUHC7qFQzOG8nBEj9jamVnG6k
O/LyH7vAZ+98V08V+rcaDhDG719PVbG9lrTD4aSA24l4RvinR3MK3RSXYGww
PbUjKqapdO7/xg8ZFHRfxozSbr5fZfaiCmpPPdifoubTejUA93lCOXAKd3tP
CNV1r4EgyYjrMOpV5R6ccusBNrSLJ3JodPS/6zRxoaBuKoruDwR63jubYrtz
C8Duo6EdYtfmRJfbxbgDuRYt5vjz3wnxgfjqU8sVKNbTsfz9oTGm4Vdqq2Q1
XXwqY5fKLf43oLkIfKtoNjrC3wskkroWp4GHmZn2jxsxUCwo29/Zgx3RfuDv
LEWAuOmK+sFuIhEpytxOqxue9jGFCFKnMhFt1OuF0s9chMDG2AG6ofSsACN+
N4viy3EPfcuNfy6T0svjlnr8ClOheA/FwmicVIAolMAUfJXe2t0N5HeZ/+rZ
q9pMF8w8/bLG8A4ShStjmz1VJ9InAFFXclx1ua4d1eWB2DfXWLxpO5uub+6E
8hluv3aLl4xInxKCWnriH+dzhHMHRqSjk5wxsuEhJ0mioC26m0eA+TsDvq3/
S30vPhVvGm3cy/s/NCVr3vpyTnkZbSy8HWvjjvAg3GH3oL0QmgZBmCy81xJp
h+XHogYNgflS3UkWhgHoau7ti8KOrXZ1wC/fIDKONnyRCAq+RxSAvc0mTgqu
oz15EpLk4zx/OTXGggZyTCKNakAhyBqDl4q7HsJu6fRY3A+eT77TlAYMAH06
e0TQejfh4XtZogSNA/zylJ8UaZNp+YfZzAgWHO+om/EOOVoNCQNLgN1YNZjM
C1R/CDcieLqHafY6Gflvo2sMSgQD+uPzB64pWiPFD8lRyAnEVOYN2IWXvP1g
xa/c6YJow/QLV2SKVXE3c9IBuLPQbEovo99cRSKoshFs8pq7RIDjZdG9OOCe
4osMIIeqHsJYq21Ti+rEzeZD6fSABeK4t2qFyC6kJ2dhDsaG28p4wTcunIBc
xeHxiWRCxK8WNN1CGNGbu0K1vkNN57gNp8Uh8VUEr7O97UTmlGzcOqOa4K0B
kDtftNYJcEMAFdkypH5zlw4pcqACoAKQjG5h0lVLY3nOSghGShcEBnKVJkCm
QibWpp10EN//quTUXeLu7G+aGbtGmUoJ96oCuQfRXEoC8X17xZXfTl7uytJN
LZTc6ofdbq3YAcx0e00k7CDP6JWgEImtCrQtZvR3u7J+C5+aHkHMwNledXUM
xeb1inBd1Mr9akyFIRLTX5MBzXHfPGGsQRLS1Gv3iFKMaNo2US887DZ+niWQ
2bEgCLn5YmvKDJTZGsIiZcnc2t1dNmL2MEgWjR5uWqVB6Vmo8cYS0xGYbSB0
ydWdhbjSKj4AI0ueJLxzWZPZJqdxXTF5g3+v0SnBkNdcWrlV43MBFF+Rd/Lp
+lrBY9Bb/+c/9yeZqDcP8+yRrImZSLjhbJJjOa6QEqaxdJSP4O21oCfLE+MD
WrcS+wHCbtWTMOZvswDDygcsosJdBXOMFDh2+nxpjlTdqKuRiPHVPcBcpq1r
4fLI3GKCgOkBhx5ZCfd61n6qJXvYB4BrKwxZA2229lXKRmJ1V/faO1vEGzOu
pCElYh9ZUvegpT4EjEofyAWaMSDdLBIVk9MzkopDtHqpcrT06mJwaA9tZkEz
UlPeb6kZWccbcOh6tW5Qd/8gYFImG0RyAGQnTPYOLQtO6pOM03eDEU7lH/Sg
eC53JnuNTPIoK15LZifQ4/vkI0P/hB1RziLEOqT0SCqEXZDa+bNCZrCid6nL
pWS9vdQqL10Lqx3BUWJcFJ99n6SXjms1S962OHijvxGrh8BZAuKbHmNbLzMG
6/dQiniGHyioWFEhZOnkRymOFv0hjPKeRVK2HhcBIVMT6YBltS4PLZ1wCRBp
0z1OFDX3ddqLRfWwaTUoxOVx5NDLKBd5BcaecbNlE+Vi8IOzZl5PMKvbQN16
955HXB4MaxnE5amdqd881Fqkd5D6bwx+BnXXH9O414aoUJ3/MbsuvLnMbrCF
Ncm8GZrp4yp+UjpaSnEgjMficKecOoen/UoVZq6wXBEpCXO2PsJx8VIYtFH0
ppJ3VSQTNAvMJo4fma2/pRWdvcgfZI4k1BlnzvUNUK2VormOimu+ES12YbaN
WkVlncqoxhUTEIhFjPAYFr/pM2CJ2QkPbSmvO+edei6w1/sWxM47lV1Zi9pW
WTRYs5iaz0p+6DeO+/o6g1CePByQb2Uo8gQhwR4ibW+qGSm7g+IOdODV4Jlq
GQSMxUF8PKxVr3rJfKqdVMOxe/Dj9D9ejjhrlOkbUoGytKBYThFYxlEwzho2
OneRg89zNbyvDtTp9+Ey8QqklEyN59p6Wr0AxpyGSpJCzRlTqMdqcAv0Rpou
avy+SdgmkD3SP/pBmFiK219tVLPlAjJz3gTlaSytm770MGaWhFSuh/ykEyIU
Ov1Z4Q6uauFuwJ8qbP9uuTvQHCJ0/cPTLPZoe8coZHyNJQJbGco+0FLn09iG
I6rrHbRBxfFBdhsd+ekZ6DHoL9Ea852F9MLreAAERjt3kazmyrquuueb7wOm
9AWAtWZEidXibYP20/MjqflB6uVhcKea4xcRdwoQV/NTL5+W93PboRUu5HRQ
EtBVsYKe++x5g2FVMyxbxbGlt/RP0U/B9d2tZ1A9aH0hlAO/SUrVfRmLcK22
WT5T82h6K+FM/QYoDwBuPR8/w0d4sjJB4i9EfS55wTAiBKspe1KH7sVHileW
Ze7LYYIDGSlBP2O35nepw/PPArN4dVnPJVExwMdxia5Oh52ME3jvsnNJAUOc
MZKE1q6Zc2CY3o20VtKhHFpQS3NJsMsaObd48fCUT1S6NIP3rWwWYPntZGD4
rIUsjiCa8hkaqb6NgEp02hjM+r2thqT4AGa4IbaO1H0K4yzLOp5Sz5GL2Sh4
xf8KWtPkx40Q5FcoXUwcPOAVNZNfvZjZHpFe146/OezTAlzlIVOySp/Jny/X
UTvvneBPEE54CvpnyRhhTUkfxUoAsXOnlzZ0g7OJV82+hHFdRkD8k70f5nX9
qQyy/kv8EdnyqIhg0rDmGaS0ZYIfHhYTEu7BvmJ965LaSLMv2ASqIhu7sQ9f
nU4r2EtdZ8G/PQuoMNacy5loGqTZSN02ntoIRCmY6a6IL/yN9CLJb3eQktiw
HhyQ1GzwK9BK7bl8Ec3bH16EZMMdIK3GTNkLZM+HzZisl0fLBMN7o70IkWUK
J1fGofXt82Cr1Gh2l09OtQiajEfvcFa9Se6cLCRGcw6fvTUz2w5af9YQBKxb
sVIWBjMG6sRPymMD3qx7mxQU0vSRT7TVnTJ1kZ6Qmx8/4DK/kT/y8+HvhMSB
dIF8tLHbGRb+ULRrjAIlZmBRH8BVpC/Q8r13RFp3joyw/GYGZ792Za1a3Pl4
z6XNNYyL/rHoFllvZWX8vuBoalRTPidNyv+M4FrQ2zkdAnvrLdnx6JHvHWmm
BowdVRCuyJGbdcpDQMH40UkQYCO7mdT+ECs/fj6a2/6I/9yV0CMWuqR1mftb
EnNaaAhcVoUq+IdgU8vq0QaiB0sG/0XmbA68CTIhfVG78aPTXeoKzC41KBIG
bryufucRfYCFDwZ5sbEK+FmAgx/n9fd1Zb3UJfJ3iFFHw9hC0qChJHTTxgsb
B3/F6a2UgUg2+/V2U0rif7ZnySQK8tcKQ76G0A4bs3wY3al+OJIIkqSKD1dx
x6ghLI5lB+YegVdi4rkpCxQw05VKA2ppux1tb0W4s4wFnQsqGhseYNOByZOZ
1smWZ6VfGyaZaXLfDn/Wk4O5AcvAnUc7N5HvTAKTruaj3XhBc04BxM4POGKY
gNpD4dYuV6OtwHIGkLNl03455o+QEJTjlJQe1rXQxN91U5WrpJrqji/HwGV6
67da4pM5j4BKKg3vsCVzqPtPZ5HgUo9mcE5kd4CIhm8EoA73uBOhnokO73RT
aOLxTc5bOtW78USFqaYIAzHMxrJzX0XOw0jSluNnMM4seRMAHDc5cTBRNVHP
Wy1h1U14dSSjQFcuxehZ2+85oMug/XJc9oY5APiqJMeE7Wd6P8268b5m01z1
APRI9CIcRrUnBPrNx5HhPZ9SMxLlibL9Ffb77j/pyipPVTeCD5OfuBMP6jNR
EmsBGRuSCu8IkX4j2MDBrB/CfAMvPgsrw3E0fuLA1H/UOnsRa3AmSIpKEv4F
j1zr998B0TUaqkmr7AyO1pgwO3IQE6+cQybpADaTt4mo5eflOMVkJKe+PHgp
G5kJH/DYydOVvyiqyHaIJGiX95QO2kB7hlHRXzujyyNIk/s63zFViRIgGQWZ
zDyc4qqZ6WNKFi2vlAeYR1neNjBuWYlOr60occLToC+ErYONNF4eLmI2zc99
ps/PwkyRsd1Nva5MBr5jpA09OthUU9yP5NSZXMalIzz/anRe1QmjTbaXxKm6
KcZOSmCWNXfyiaAySmvSOXBCY3HMohDMXcrqqb0IfJVObn/AGZK0UTl2oZvl
tlBDOkdZLwakYuH6290MTff9uUvsB9j5cDYKADLNuTYOs4/J0yN2czLz4k0y
ScqxPXPGHk23R18javJqX214kWpLvrraSCUGl39Ni5N/SNyvsp2fxNVo0Trs
HVvbGVK2I0cIRgP4/pnnBwvKp/i05aT+8qX9to8H49uIBy6lo4GPik/rgoHp
bkCaRw84MVRaQPucvg18bVS1+N5ph8ciN1VU9wp23KbRgrKvVvd3te/3QpLX
I7cU8RnGC0x+/BM7zLclcGKtOYfI88u9XIqjmi2eWG80DHnxlQPiKjBoY+SI
hhFe+Tr3lPppugJ1w4PztEEuIYCE9kW7/hqjGxDq2Lf+qjeVpbv1OBJo3iYU
W+G7ESRw5369Ru/Eq15FPmv1M46miqkBkMpnIeDKaWPU9YJMu9vGznq9lnnp
omqp2mwHpCroRm0dSFaNLxTD3LCTr7KPPHGwfPt2nAJmQJJRUjNUG/FzbMu3
ZYZHyA/EQoj666/8egHHtT/G+XdgChB9vvIPK7pxXkn9s6vS271LhvZ0WuY5
kCpcqeys2j4YMxIhWFFSXe+oAvDJ1xehzQZz0k03I4F4H4e7XIXrn3evmKYJ
MG4RsVna2mahf6OIJIjvCC/Vsp237x0a2EZH6kTSK14bFrdU+m0jTOUT/CZ3
y28UTnsj2VjZxwPdCq+269b7ipFSSA1aTuwdvLjWunDSNUq5eIVHGlnn3lNr
vTNAgWcmunpnGD7+KiOrHoFK1x0ntbzclN8+me+3mVK4WTAaKj6QeBPr/mez
2+5d8M6esi3qJlrmwYr+zlOSgeUjTZfwJkaeo0hbA3UjkOWNXlKL3pvzN08Y
J9mRvVg9Lq6wy4wZzaWqMbxSL0557kGkyaNB3YtBCmG09b9mACAwuosdch6/
xJP7YxLOaMBd6yYEqT2T7rlNLeLMNZWlxbfg7eBgCKDRLzckyupDdvmPMQfP
Xeccvb6ZNelLZhygqrs5SExrrvL58HQjWniXYSrEYop5JtQvfLUgt1vLP+uy
VAKOCQOcp1N/NiOsK3Clqr4mF+ONyb2wje8dyumcYnw5suGfzn5iR36yB0zl
gK/rKc5JZj2Au2cWwHapIS9ZcuKjSbZI9X3bPVxBAQ+ej0g0kY2gIePooIa5
/QsVEovLicE0E3JYaTq0gwJCQzO/ZA0/4sOdQ3NsxSN2PEME0s62aL/Jh4HQ
1DCkf8TP3y4RXT7MvGvrJUdQwjuizpFXSDfBCRC3gZCytMy6Wf1PkhVSHYAO
UFUh7RdIELHtsdOuad4UbM+MNhVhcTXPurACYcc+i2KnO6nMnpySh+XxdE75
w6uh9AwQ9bNGk4mB1KvYBi2Tv5OZbIdEXB8hbDPyVqlEK5lOnQBDAjASo1Uc
TTqThBxx15i8x06h5yzLkJIsMvWHXa3903hI7XQgiV6fZDUVLUXFkvPdbKkT
ooMbkB84Qi33YvW0cIdowJcwp2OwOhuIsgQGAb+kftrFTK+v5Ss8mZjFTtJu
xrbKPXlEriViUNUT1azChXqLosauUaix5OgUPhMHGJsQruJY98TkV1hyZRHH
z7OMUnLutWVmnRsZeId32FhMLEGH2jKE7iijAWizSbTuTFwrJgqU7ZJWW7tm
HqVX+cWmfxOYYZGa5XdxPq3CNzFkzxtCwZn33UJC6IlDp+f2hwk49kfpA6om
rUq0lge+j0wFCnRdhqe8cP7jNVe69THJTW1RyKsWnf04v9hnS9gqCvSghG43
DnUpcJtjACznK3z0vWdWHaT6QR91ED6gxjo8C17KGdw+uVdjVT/1gk42/4Db
09UPRRHE8Od5zqJSdKTHmFDYE7QEQJBVz99Dd7yqMWDrkU9HfuIFrIYDUib7
14SNDbLkCP71/xZf+E1+gL3/VLW7bYM3Kxb9siknZN/66PFluUiI4ITAH86l
YrB4kGEbXP6ICiJ7jiOrNQLGJtIIe+11sI/dhb0fONilH3MLMveQRrvd6UKN
gWLuJvUt29rSiJc6fFPpZR1UT/mahgVmyqgFHq7Xj9IT1H4YR8mbXbl+uElC
/j52E2aN8pBkTHDtzPI0dSnZvozHpqJiSwFCR7XRzIKw6vNTPT2szULMknhQ
6UTw3IMr8pFU4H+4fZj0Gc/BWfYXc6vwHQ+WCUityXe51HH2cIanmnO8S4Jr
zrwL39MyI/DwSLcM7mRZ310Sj89Uf/Hf5CKSHDZOa8eY4aV47CwTLpCcpDgU
u1q7+eXaYsCPrYsikBx7KtYsuC+ZQjt84oUwse+GZvmntD8g4bLGytHPLcOz
uM38yzzWq6/SBDe/ectMqTQfvCOZKUt92oVByDP2jmZ+Nm//yHzT6GdCg17Y
/zFKzvb8R/oUSygp6dV2KBK7N5j3FKET943rlSI5kOk+1HaZ4Ol/ooLBUr/4
gbCe92dcZlFpRoskp/+rtTrBIIFIPMM+Mc2sFrWwZomFMZwhh7Pc8HV/BB73
XMb5gcieFSgxqWumzjmNsZuXMUrAXul6bB85aBtHCnZ8D2Dy/Z4F+ddoxXmK
vpvvtmym90ML35FcM8hspmu21IObLfERmxN2MNk7y/QJAQhqXdiWOWxO6lba
pQ44hzQPkdx7HXL8g3ILg9i4hN4Dn3Wu5m0ytcaQpDWkizVl7D72qfdWPL/+
09naFXGxKD7Zk/IbN3rC9kagA7C6gj3aSJbnmP/gMG+CssN/Xjf83PgcHGC3
1M6psRCUBqhd6qj9vSrJRWFBZTjpXpveIXx0vp7ICYXZe3fcFhIbA/ZvaGL+
BlYBdMjTNf6gBOhTwUNh6rnvPaCONdi0cMfqMN8oMH2MTA+SYO3HXW9t0iVq
nbpMf3Mn1UC0TgXPSEBpbxTIZoDbP3h2rXtVvX8TLY4uvNfSuC+J5qwL/ugC
5PkSxVldle6jJ7UmQCPuByQkmT4D93QvP1/6gB6B5tFf3u22DCMti/mBEYov
yAcRBVUW3a5GJiXXvprX2l+VhzG/u4j9yDSwWRqkYs+jBq+0OQViZ/9uNB5l
PdfXpByGTcFOTUqocjcW8fYNR7J49jffdWm0IvsKC34nEOS/8jHAMO6YXnlq
1PdE0dKOJ1IUZpkL2Bt0d3ZIHyjlMJHv0dMEN0JzjmhdvVScMoyTGhlnOGE4
fcE94mplSQaGvZeffU1TXTpy3XLB0CsG1dP/RNkGQxi1jTVEgqYQB/V0ScgL
q+iG4b9uwNV+X70WJP13BSvTSPsyY21mQMxZrK785kalo2VqiyooFKFhv3f/
J6hJs6mSzYFHzpsByWYs/K+4AE1lQNDpwLsOHC8/WB45BssD0ZSWAW4Rq/MY
E2YtBbujwbVCPQH7I2Pkg5AuCWDIGfAAOMzE7J7iZ3o/rgGkaELcll05ESa9
NAJHjjgIUhcnGM7tuhwYuhEGtqRZTfb6lYS4nPhNhwLLcMyeZx33naQ/AkqN
bxseyciER0H84w5GGKesolOeEKaMLLZ5KNzLmlkwbS1kyTjV+1YC7NfeKTOg
4gf2XHfHRV6p2jz9yCPn74wFqAhCI+tEx9ejPN1cd01FyU7M7moSXtR327Ve
LS25/FTh3iDbtzGJVDz9tVXPzucuLFElqJqk8/Ro4tTXIrqfMHZWn7zj9QPL
49uzpb52i/XwoXSV8+WLufmHTY4vTlP7D1O6taeevmqNxdkYn7cdGp2PPR5b
3wImUgDpQooKJgBtcSsH4GGz4nmPN6AHOk23SqVEny67TX3jj7jQnxp1Kl4T
tXmnx5aFZTiZ/8Jmh7wvWAYqTI45RwRFECry0efEbyuC051vc07POqDYUGP0
S8NyMQys1Gg3/y8ckjLI1uW2aNYIDl7bDtQ68sBVIo2lPjX/qhIatQv003Vh
w3QoqM24OQcYD3H72V2aZ2qQ8yZDYon48DrIEs8kBIXafts/Nwaq8ZQ14GaR
+O2R03r42PLI85Qk/5zyLMQKQy+RPq6NBG997E4vebemYhow3iZ0djwKj2+z
vawGak1efnmRCbwbC/BL7My2KrbPhMY3ONiObrk78AnFWSul9uUAhGb5saYF
5ayIvj1K86bbOnCW3u8n7nyq+hBmp7VpySrfxm1kX2k/oJ6BzPGrJS4GOMoa
wscH/Gj/bPHY0C+wchkO5Ha3PIZbvCjEIPHZ8MIxIz+c+lABWrElBqchGffc
gwB3acSeTkOiGnWMN8FjZgjpm4FJgRArutGBV9gpf1hpB9emWCaaeXbrcGGH
v/aDfxcS8is1145Fo2RVd4717jRJqHN0XTgE8KIHWtgFFbBTKYBH0aeroyU9
sv0pSnEEyN4kThotnfSK+5bg6e/kImMuQux6ua08/qYMOv/Et2rLaa82aNwP
lw5FCV/einol8QuUiLiM5d3D1DD54Cg9uEfEouksxhaO57XMtvLZGWQv1165
kQkQelB878a6dkPamuNOrRTJoPDQp9M3FhZQXizM59HvQAR9BPJlOb1091W6
hBVbBr5dj0KEcu1qeqrea3FxJm0WikDm81VjHamedCW43BCbbBA9aMQ6TzEj
aW8oDTHTwcx6WNGyX5C0dz6Un0vA7dThb7/E2DYeLuTEcXihXp+eMbePI2E8
Al7L/XbvWXKWRMYLsg/7l7RAtfyhpf6ZdqBDNB2v3IJSyD+EpaxqYpRqLlBh
fhXisrWD6nFaRBI0dcJmLTCWob8BBweS08dIiORl311WIkPuln+A0I+0m75d
gSliR+3OzysAYfblleQkOGLYjcp963VPEpcv83YRxDioQM44UdDKnX9r68PB
2ICH7ErVRcjyT8L3d9zBDHvbxWJVSFWgdo97TWQvqE4YN5D/6vauP2ITRIVR
XUNd8uYPQIgMrtTnlf5enfeADmvMAQdSkR5GPrQQHZeVf5uwMAACw90I3B0b
9uC17fwJLI4SeJ2GI7teXlTz4F6BjS2L1MNj3RhP4UwRNMdE797VgwbabKHC
cO+JnouxHkqeaMnkkCNbjOzZlbXLSg++DYaR9gqoQE605tamRuqBncOG0T0V
qTKlC1kNeGLHMzIr4LL/c006rtrrRLtkoWLuI4nYjvAoZNnYNeVr/7fzNFpU
6YO0mBdncmtbFe3mU0xKrLyITXKVaBPTp0ENkXaC2G4Re/HSqhTAs6uJaBrL
+FPYDu2J7h80DmOnLwp3HYiO2qy6njN/G4IglI4BQ344aGp7B5j6D8RQq41+
YGJqZYrphI5wvC9v9m6R+6Up8SHYrrt4yJRtDDggNQX2fCDi6v5dUIN9qcyj
TI0i+gUaCpvtnHZNB57ospnvbzEJNo6JKjHQwA/g4mh8E14i9uf6etxaCZc5
Up8rNz6JMSoFHz46ztmFAmxsfT6ku37XwUT7+PfZc5Qa1fkcYeshSVkF3HPK
a4ghYeWDhKZYuNJhCcZQNN7/D8MrJi3pL4ejsS7YxwqJfN/PP9F0/RivfxTo
lvmyehI27P15UiBcUjHHw/5jjTc32hqAEp+7CmwhvG+h4yTteiBPQZQdxRRi
NzzkXrsoEJU5VRn10TGQtEC+QcC9y1ZYKl5DlUF4EJC8ZK/dvTA+nkTCW27c
hT6k1fm+85MDIvUNpvjov3jk7F6J9yjOH8F4zwie/N+55W3icIipuSBNauTU
qG9lkntrHzBx06p+IbDpG6Q3FfGBP2UZxh9z7bg35EYBpr7pQJkW3or7a+fv
66nS19dx/St6r05ww46sSPf/lhGT3DpMG+WmLAaO+ZKFou7yqr+wgBOmhY3b
04scuTQmhqhEYtLJVTWtXSrGNDSIlPbtO7kKeXDoFJOTy7ML/TK0MEBMtEup
7dmNuK8i0dsUYuEhPlif/mIfFap+gbJ4EWg8aacRKanMPRajMa8Fc6l6JgHP
vrYt62/joC+Fn8PhebzaRLUWPyMIwhe5WjrU4Gf/ygdOqaOu+cuzM9czHxoQ
e1sotloGRYh85kF0pA6+lon3IEGmJDMh9kHBQMTlNbt+76vAUg4YiHIuOofg
QwOsc0trxtF/IOf7QrEtU5JSdj0aR5TlI0CVRjBp67oLQtqn5LwYUvt6Z8Tz
UU29Xii4ZgHFz9sUHMoB+jtfOh3aIO6CcJhL9nkSo/KmPg5OY+mKz3NrRFnz
ebaSf42DVex9fmrFxQr6HbX30gYV6B7GEBf0SBdEaG3lBBY6lNYr8qRWeeaT
VK9I4WdCSZqbCyboxDJlgKSthc62atSmzIaYv/sryE57Mmq2+iG3/1rHU7E5
qdnkKoH+h+5/brsopIW5n8TxXu6vpUxFK4ck8FvkaTEW0Mmy6LSvLXE+/d0M
nsYOuKE0w75sUS7ZtBJ5Qr4ALXiQh+qINIe+6sK8Xt71XdxyFFd9ihEOgyPC
9ppeWMzk6CUWZN3N3HFWu9uZz3euhessaInQE39h48RvA+y4rPpPfvpIuZgd
KXRZ73Dljj6uht0V2yrAQBfcOE+JLOqgpgCBT1XSRfJhg8uvAqPf5eoL/vp+
MGacszq6PVwBnEfy+4/7N8wxQmINZMKUO4ZcOklKnxaeoHfYKybsHmqeOqQY
nvW+yRh8ozq1grZlBEamhhkamRLOmbV6pIRab2cnJXJ6Ahpyn0fWZe3uSGUs
mpn195SSy+O8C+RuY90sO19QOEi6UGjgEtW9uExCUBi6wmNOpGcwLM2mOiCe
HzV9bkE5ke6O75Mzcvz/aElxNjNZJlqDCass/YtUxewfIjP+8UXjsSNfmJOk
3zk618bSj9micGdHjRw5/JVsQQXfsHmwXuvyoR7v3C0o7akbzmFMVbsVbwFP
7doixMu1GH5BkR6o58lGeiKXk3DcngjCROPWGkJ6FjCuzdjJrNd56A/otbdK
A0ybI2mzTiSTea3uHiOeQpesnA2YPEU3aZis0VTSddUKiomSC5rsqoFuUKzV
kh3zwNrKh7YAFWU+TxynlzLg1+Q4EViOvqQmPBSIQOAZY1v4nVd/qknXWYpO
27nrRtvkBTN/JBzRfOIlhp0XJRcQhE0qXX1qvDzpTBb9uXXUAcyTHK+TjBIv
p40nYFg2oFnO01WZ1wuDD9OOiOTqlzKuP70sD19WyberXXk/EXqK3mf2aJDz
cGzjWZX9zBYclew6k9k8HmheZozne9ji7byp8VfPT6A8yt7NQr1GniICXBum
uIQSCOqC62meA0C42lbI5yeIWrM77wT0DAyAdE5E/ezJnX3PSzrHECIPdtUh
QWOJL4o76DIv1Tu9EiZgZNtX9mD0fAGkwJvHsu9ZfQfEW+vJ0NJxW739ho1B
OJsQjCgftRYu0aAUkg6j6QjYl9Ny3KHEu3J0A4AphmFmbVu3hs8BfhKuLry5
yShNS02+0c7gwyFapV2OifcdL7A8OavQYqpRfbhDb8pseHeXH6D1a86/eS2u
lkgB/0ZICRt9WsNbcKfefSZDrUKF69dymRzTa1sxpHP0hSCcBtpwe9Uzmxz1
VfMs7IeFawjxpnUYXEYWdNYbGc4nNLgINJYf5kt9AlhtG6QzmJQY78IZ5kEf
rw+zFagIgD6lxGxN+zckN0irm9GaZ9Bi85YC9wzfGc4Fr42tdoYHmD0JvI0C
XO94Y1Egx/gCYNP2ODv+oevP1aU3CVXGtrqe2C927P/YNTaxNq6FA6q+1wUp
UvF16LxXwfU+xxXntVoDnJR+Ha59kiADlCFbLt5xbhYnlMcgm3BKyTYBSiNm
Igj8p7gdspnVbKQDcu4vZ5F89lCbRfxuNbt1AJ8ECdnLL90CCOSF8DKnh5S6
zpNZL6brpEHgpd4pZ5B0H2vaPoK83CHMrDwyRXdE2NO75IjNjPC7ca3NeUjp
1jYJlaYim/A8cYaF2R3YSa1BL3+KrMO7vuIfXyTDPnwd+y09JlbKkcEQLMm+
lu35lrNq7MLo9V6YpBGyO5z967RZA2FYhZboB+O/lQAtyvCTZn9NqiTlJWSl
QlQtkMPj19dMCECEZv4ubhcp7TKPqNHqkjcLJJn6YtxztCqvjcnc3Q/BbRaE
MEB0NzmJHwhki4XCtKY22RFdvEzuQNU4RTCmBGOwqm9Swu6UwVjhhKW7dyyi
qSr+vVYUSyoOeaTo3JOYwTnvg7Qu1WDjK+jA9IOm3nzvMV0sZjCQ9CAcOrAi
dzmBhdhv0A/XdYP/kC8ox9EMAErciAHcHmkS+q/YMOWW9wjbYsxa+kD5erE+
nBB0vR8A1IN/vWfQzVlgjG2oNWIIHsMWPQACtli9V73fz3tX9nvlgJDdzHK0
iY9tf9jFNOyuozqUy/2Jjz5Q9G/0jSY2M4T9lZ4gpPzqko8uSEzAITYC9XnL
Unr6FWxwrrtLVDQuZyaLpTjp7xmiBJI4rkM9pZsaRHPIbxw5dEaMnNxlvHqf
V+Gl0ze0efKopjiMAaVU3yRAc7HQ8yZDtpzL+7gWYuF5Jr7g5dwR8dFMeNy+
FxTafgz6wk2Ouw1frKbCAa11o0VKU4KkjF7B9yKqhnI3XZOmJx3jUPKjb0Fi
Ixhn32kynEh7jKUSqImWEhZhvn/vtsDqQ5f+CWU4XLTuOwRIRNx8t0bq67M5
h5Rl9URRv/M8bDkxjFTSNCOxh5fKh2CarJIqUkRVXI8yix6f2yj5w+6IP5q8
fpheJ35T9brAtuz0vAIC6TpNLPIUD9408UdCSe+Oq12SFmxqmKyfXpMfcAHm
hpaD02T+viZg4CoAI4BRZRW9tHxp25UZQL8g137PhTfHi0QaaRB2VgMz3G2M
rrXNqu75vX7Kzcjj6R6+wwZYwYVUDkHShvpJ2WC0MJJBHK+TbFUCtiFBgjIF
6bW7SZ4ch9kdVmzfgQzqJx/P5c3zV4aImVAVOc1NCVlJjksGkl8nP+J4bwFG
VLqNlRUB5xzxXp5iez7VqXA44IorNVuPKmqChaf/+OLETTZXKol4x7ojMXsW
0ktvewEr8sdOBW2BRt/jegtA5JZ7AvdOhxk6lZkoQPtqoshnTMSx/T61cpPb
7U+wf7EtiM6HVoOnxKGqGrO+CNj1M2d3JVe7hucnO1b9UBJfvbnX205Ko4M8
0PKS+4HWP7TAxcnwuR08visoOuod/jGxV4Q4zZprKSZ90107ZI/zl0fUs6az
psrdnojIT2guGymGMifs5549Ib27vgaUnxQ7aS8nnRZFNi3IAOX++t+VSVhS
DKHnVsH6YlmUNxJIS/dpnm1o/rX2uloU94Y89Siea0jk+hq/4YPDY1v4ZhYH
meLCPLaUXJ8EvOo0kURJmfqfJHpDKXkYVz5SgyESc+Eb31VxeH5ij5PxkLZr
Z28jXWg7+8/CeY2T1sphl2YVFMvwDxIq0DgpmYX4rWY0BG4Hh/z+uhp9LK3H
UI8hHpHXjwz70JCDYvBO7e7LnEKaToHPbIa+IXlBO0JKgbfoyvA1A+8t5XBN
UnKHiHDwMAcpgJwhxfr3WBQhzYvubZH7LWZHSi2qtftcsjgyFuHQwEcbHeet
6C2j8mVp5wR8isJaCDC+BdgygyYvGP4MbyrDsaeYzWYPAEdS9qtPVl3UU8Q3
7tDAvTGxr6WbWiEXB4GISQdx3zuzdPJD4n7pkNcDFpenTn1qVJXVrI4zngxa
YrsYeC21mQHY8nZbHVu0D57q4EkcKtYdw+uh+R37Q4Oavf6riRb1gUmJ0d9v
KjWz/DO67999k3n4l66DZvUHIOKWvdHqXsAmG+FcUjwyKkVZqrfGSYnVS7Oa
2wY9SlVg5tW2Ra/qNXSyB9/OG9b6MFxdFI9CrPVFCxVcFCgbtNmEBMt4pQ4Y
7qvnhEo2qBvOT8z9KqtmXQ/FjYFdKdFqSb57c6ZKGDWHrOSc8TsZEsw3PLdu
9ccD02MhxRA9eyHLWQMuXIIXceHpfRThwCjguBB0tbfW+GnIjhMEu3hqgYMJ
qk8ku/RMaBsbdexIAuv0JF5AlJ/66YdeGRyxAhygqMhe2G2uf3NSf9FYA/Nq
9EfVtzf1Ji5djeA+wfdnR7X2CG3wXRYCTQ6jDzeQ9m9lj+xG3VBcVNAsgt4D
PWb0p64N03WIeBtAkk71RXBzvWNd7HTM+FyBNOECAZfr2q499sF5zpZnKDXi
1Wrac8RR0WBq3t+yLiGVpQH3kjMTl0cgRdYGlK2bkfSpXIjL/Pd9oYgP/mvD
YwN13NoMuYip37XSN05einYSSOd+y/6CL9LjePLDpC8vy1tFRAlkuCOpKFWI
bRj7fMXAF/4fpCOhzLbZfenHwF7Flu8QBqju/vuj7BlfvORXhSjXWiD2Q/yK
rqMVW9mkYb6m1+0HIrffn8lcMSw3S5qZNTZF2XQ6hq807V25KtigCJTwNYCv
dlpWjoWQIHjGMpi88gPTXPl6Tsk67imQIPnnk1mVQKZj9KEa6HMJ/rfqFctA
PV0MI0e7he+/0UiZiNGmL10MHBywba9RmpBph5Yv6lUehlnCpK8eapelwCPW
2reH3n1OA+ORTnHkHqgfGvUJjxRkiz1HBkLKynpDoYZU8alHhSIoGXbkl1mO
4je8hdcc4ki26jFHyMu6fXgHvVkFZRIgvurWv4h50u3VNfzb5t5r3FBRsdi3
LW2btk+odTnx5qumS85kJPU2D93+aCuPexCT3kqgI/R30R+Q5xrTRkUyqz/m
4L4rYujFmRCcDT5LZJFrEWT34eSJpjju700lQ5GR+uAWDZe36SBcF3s5nDQR
ZYPU+XPCQ//pRtOIy2ZJDRY++BVAfbJhtyu0qA6DboRMCrjJVtaOkVOGCRUV
3RUf03++1paR4hnfXtN1iica5O0FV/aLwp5f72Mg3BB+iu2uAaixm9IxObVn
3wZRn0b4WNW0InBvhlNLpPuu5ZSCHyywYvMZrmmxpX/vcNpMHn8bjLSZos8Q
fzA+Pu7CgBxegE2uPwhiBRi4ktjKmlduLGk1Ah18rZPH21+jiPi2tcc4Ibhj
zwG1vUvIOLWchMHjrs7MSpV7OTm3VqutYffHSuAuvBs5BcVTUXuAdNeNha6k
3LnDeC2fDWm10S4d+mt3eF1m0m4TfUEPcGXj7IVWZrImyxo/coS0Tk909O4D
OHepQ1EVLIu4sCe3EHQ1gPi+naVoFpmNVNxt+HUGs7Q7Ni69TKJ94aKz/nTN
ph8KUkVJrhh/6ldyJJ+9YxPUL0+ggWmRg8Jqmy1gRP3eTO1TY43MDfN6Fo3j
5ivTHkYFUkk+1Ug84+pqr5dgzXz+5xXiBGyhOEEJMeyD0wu8eVXMKoJPDwyh
/tMDjvuErQMElSymzXnzDMBlBLasOjvhjV7qWQ3nSp79F3X7484enzfVAxEr
Z+YKmPa52LbfMvJS1GHZkXsc++AgBquLG+Q6/+NzJTsHwWkPY5CEmY2gE0r+
dgoCTubmheydsgLVQLjul3i1VnpqdsdHTKJEj/fh0JOU2ICit2vYrt56pXoL
anAqF6O/ilXLVBq1+fDmLRIHb1hvNvxBp/ODx75dHXdX8EAbHjCUv71t4CBA
c+lvS4Vahy3Q1r83l/3zdUzw2MXOcwWuQTMkD4VIZNxGXJ8LpSOzii+yAgRk
Cuct2Bg1ocqS5jbu2C2yBtE6bGJBCHWBx/fgiZWQCcXdlogak/wjcWSkety1
S3XtrdY1AD1CZyNdU993oQQgBfkvqU6Y4sqqe4g/jBUy0AyfPFhjzPyMqjw2
6/deICGU9x/sZOdQGDAn8qPq1h3ccw/40nRT7NDG7hiMRSov0bOoJqOpbwjm
IgWpa1WPlhAcx0QwRVBMFKxZ1C/tAulbeE2MwklwfT6CLgNXMnzYiQH1YRn6
b1aepGHgQYlI8Byr+UjX67Xe/3sJP6mmfxmd3JCO8H2Jz7/dw4s+6c7FRRP+
MgfxSLxfk1LWg2O4ld/5h0bhYgwxDmsebr1Pp+/p84LrLBi80GWX57D2OdY8
x3q5pSdS8YqQe6GwOpUrm8uOpcj40PYbLccwM3FuD+bAHdvf+TtvwhcXNLeE
UdDF43RhUVSXIsGOLr9McC11JwiTjP00NPoNqg7BiMCHYOtoSe9Rnin5jUG7
XY7SlF8wj0nBHNMuUdnHviOZ/yJ3NBk8Tmzldoc/2JJHBG126ghWu9VyjIfB
rRJ5UP64qTesUyw5CgpChch0e9mrJXGwwOFIAOpGFs9z3215q60yw3PYIGZZ
M1cxjUmcUJ1ipLBiLz8u17dCf6XjsE/Ac/zREHkBrsQu2O6T4DNMvcacvZ2B
0PPVfKVzCX2Q7UpoYvRanELFk601dC6GJJ/J8WrIFMOTKoaTZi2qIEAWR6HS
Xw4ygowbe0pdjWlVcMQ5mnI2cjfOF2uCPmibABMOTnWum3BgeVA6RnL0mRxq
CyjYioHffJh+4w5WIrNE8mybailrtjxHyB240RRDgQNs/F1l9KBk7tPg8UiF
+FG4oiw7obcPmarj/IfcQuiM9ob2QbWSfmJpOvkFqFCIsm0+mECICxgDI/KA
4GOnf1KKtjZ6/tW0Klw56ofwq4v4hEEz6l3sr9AWT77N9ymO7lJwcns2OhP3
JiDKLtuqvPfas8wXxGkP3CDVSPZO6590tfJ8CmkboIH+k1xwgdzPC6LEyj0/
v8N/B8opGYVGTNPI1mHZbvLEkR9YGe4UAr7i+S6QlG2/pjSYgfOBX0RQFSQh
SKEJpj5debyP5Xc3khX8nkeiNZOCC6kwgN7jgKVDpDWalyNk38CswD2ynHoo
Msg0I5gJrJDzEhvTLsEVaG6uAK3r/1eoOt7kqOjU/AxEASHVkZ98T6kR8/jd
8yxsZjAc9NCtwzgwBwicWC7Eke8+AOVWuxplVdO1Kiigsh55RN4E5sGEeLIC
+7tg9bKK/CHfNChSaX1LarqpH01mInxvClwHwcDuLA2paQlbLd9xI2NnbT2U
0RD3vXJMJ8oIJRiProCCSCFP6s31+ikZ8e4aQGyQkhTnTUrhPcFBbuDvU/Ue
hMkcJYAiXeA88shNgZAeEDx2jDLyBxCrHRTT7AvVuhn+VBxbd6wTnba71MAY
7JnkzJKvwTsTtU6Y3qn467rIjdDgkJwVHB3ndnANigjpAcYNO2gHMYvan7Eq
1eWrxJzOpJX4e9le7GcXLtLQFeIjPGY5hhmMbE7EmZTdOQbAFVwgLBA/Yfar
W3Du1xIdO06ic/3TlbLZ7aZ6R490df3MpEKU9vKlbwkw8rj8dmcNzZ/LCghi
WeQZV+YznTM93Z/NVNTkNzZGrqIqZ4rv7/snRqRgr8I3W+0ypYwSvAac80R5
BbqlFfvVbxyMoUhbotJHZBHEld8snGQIMcXb1OabCnb7lCAHgcY0u3sf2uC4
YlWMvzUlcf5FW20QOWUtWRCbuhO1jv6RHh3L9bd3EZaogtwbcD/N97YatmGt
HACiFi62I44FGP22DqykzxbuYZsqPcC7zRtr8w2YFzrI+UcenJvK3nxDRoYM
nxo7uWp2P5FrO2L9M5IGalDFYx+3wjOLtOjcskwqx22y7yFYPTVNFkMEuSvv
nTJRh8oTX2j7mCJHmjozmGObEzflBYGz3a/uGXGYTRjbfPmFOJC//E4t+eSW
8Ns2iPzkrdyRRu4nwuHSD0Z/CJr24ItEP7kmrYEBupiNWGEpwi5+UZXHISSJ
xSr6Y9YJqdR1ITY3tTPHsBLZKO5MJxkBASOc5Fhp/EA+n+v1mOvvpwe+O4JE
3TDMRXnq0PCcAwARaZeTWvcRh4CWctv7WEwYtD+vu7vs02okJK5czPat6OLk
ESRhkozenBUNO/d1G9+fei2C47XPccVAxXtytGu4SToedrpUQ1Tsl0o3vPbm
aRZt71OzRdE/iGcwOm86dYYV7WbHk5bxqMeOyVsKThoqc87Z78r77NtIBCUu
Jtk1U3iWGpL8RpbyI1fRW5OVBQfy14juOXvn5+p9fycS6kP5zZmFiTfVsOvk
JTK6YNhqA447I9wrOfbeQqqxVIvDyN5Qo1FoS2XcpTm5Mr4ia57efdZQZ4l/
NoSfqnpaTGuAAqWQEjvaROwwfBPpCr9NSufczG3V/zUk+rS9mOzQ0/TFJjQm
CnDOqbpD7Wd924jqDYRO9ntGAb/uF89eHNl7EhQY++BRcqeLCjaZD8P6iZcP
rk3f2n2aJvC4hp/rcaOgfhDysSncxJ6kOQdSFG0tAqBNJGw6M68aqZlQrWn3
4vhCEKb47K2O3MLCKfmFv7B3oom7A1mP7gV863MrqKj452l+A7amBqcweyF4
LpVCgnKf3kEbFw+hI+mv9S5/PcTqfjyzmBy+DbAxYS0ama8z2g3iJd5wjvhU
B/0bY4f4h6EuoR1lWYsoitg3CQkBNQ+AwK4WrfC6hAByqGxrV67xZY7bmg1h
DtQ4O0OtiM1N0uAWFeufTDFUsdRVK2Ce59Q4pfg3DO3l95p2vANWwAAu3FKN
RLQ/ZdCUiwBQz06sNsjbLL1UtuMlmNjn7MA+i2b4Yxa8POuycleIts1EVfok
hL4KodxA5S5Sg0C48nzjRrPoq6QfkUeOi8GmC/eVR7Ch9U26HK5fxCBDk3jE
Qisr8u5j7lfkPGHogkgmh5rzpmK0+msvoG1c0dblnPzmvNHK6f20oQgZ7uOq
xl1Os0INxu871a+YrzJn14JcoS2NQN1OGwanLZ1/awEhKKXKK81SV+WG1FLD
EJk0dRbsBP2MAzcHRKJuq2sLb4OF9E9yQ21l1kN4mX/NE+D2/pgIBWR9IUp6
piPg6UZTx89WMuKYDOWiFKlCmb8U4Q7smIiqxC8wJH/4ikA9E7WhU7DksEKm
xiH0qH6ge1Rn1AnZHGsy2HMCsB1uhig/TWWCMFUYF2gj2i9AxtBEmDtub0w2
CnjY7N7HUToDXWIM18GTD0b0UqRThoeZ5sa54odUJIFSckVEARc2r3BJLQsy
wgH2m00sBuj8903LI2hSDimBZE2YyE0dYNhYta8Rw08prJGdA/1N7zgeWTjr
VNWYEPkY7Zmq9sPUAgpnNvvRN0EFzaY+eru2kL9/JZ+Y17sYHKuXtNXRCyPQ
3Jexs8VILt8kV36g/sVJwpHMOavVRJsIZFV/MHoWJi6DDbonp9CMHOhxjIXG
73xRXOCZlTfIoMmWJ5iNgoyQHzrrN8/EFlZ5EBhUdKMil9a1UycvMOhdHcbZ
APnEwoLf+3oVxap9yei+dY+OR66FwhAdsCBuIW0/n+dj5wfwCkt39fvRVi+U
zCMAp8lq+jDI9iQcqMqZZOpn2bQpShJtKR09QRlqgg2w/DKIDHUFNlfb3xBT
+kwGwZHZE8L6zHxtte/LQyeMQDsfICaCSEJbiLyGm3O2uzcZatokTb1IKgRj
yadkovXbjHDIQKsC3ejCmaw2Wkd1deHz/j+U0mE7ay67UudTD6tcB60u/8y4
ePk9tcTWbB7fquFWXGvkBqT9eRLSmLnOyKhTpee0usPYRAOCIKMJs+qn3gr+
bIfnocP5OOp1NaUbIYMZ3TRt/21RObBIlUqb3K5y2jTlzFBcmFdkrixSm+3V
EWcBGSCjJlez1TkE+MrmiEaDe3F6Me7D8XMeMthV0YpQb6E+eO0OUyg/SnnE
5nluldeI6QOsTIw+c1/irv2galkOntoous4LPzoL1ZIie/m/w3dfBx3mTL83
BbBBPCGy4qp3CF52WSMFn+AjtvrcRqgNEjzzXD6tC4ghQh9gZYX4a8/psBy5
rDXr5IQ0dyrzGOKhsbW8Wf+f68/jYBFtpn9AOCoHSamVAp4gZmxMcmHEHs6o
fJ1FKos9tnDGEBfvjAbh/H7bREQnGMe2nKxBhD9Bw11wWhpNj1a9UuGDjvLn
kphGv0noB+MHcHH9cvuGYNV+PjLW624JJWIjBCi+Mn0OnH8kssLsxybhLy2x
5JfxZ+YIyGqhBAg+RaGG9ZtqV6UOf4lYLJiGLz4vQ+DZc+2DhqYInUGTMVqM
+d4zln0TW543TUUNqTTEzJ3qzHVPLfdWnxzXz2k3GtsVMgKQLSHgjM+Dd4y/
+m9mfeR5JAggTBx+0isqqIiSvDOmomUpp01K0xvd/+3DmFX5rCT0hh/kDFmU
0kVM2CFbSJtzHT0jQ6yyc6IIUy3ix8ryvwPG7Vsyv0/WliLj7qUDIAGeaTy3
zCgohaPJIwn3BDr+oZszBl3/AiunpILIc7my7Y4cwRAFGzokHmrhODtaDgfq
tx8FR+jWE5KthZUEeY813c3HGab9WMApZNMTaoKZsNL1kG2dAuMkAkiEOMlg
kOB0O/aN9SLgd2JY28j1xWuN1fgsfdQqDX8MSmXiJJgmdLYi4Yvkf0FqKCTe
1Jw5UIEoQy/4VBuEF1qr2WF+3FcQdWMQ8phO4RP0woffvLmKcKWvBCsmpKq/
m6gwEdmwJS6YsLsNWK7LTsEYwjuYC+zeAeByhRKaDEYoomdDQBvpih52yQqd
ChtLyKtUp0XckQpDRn0NhNdzTCE6yE13n+SsZ52lYsulMQ0BiyEwAWovI6gb
wuEPgGpAGOfjhgKFvLpwdvluwpxIWcrnfdvYt18srovcucZ7beIvvwzTKu52
0jZDdFlTXQPtpkc3R98WhZHPpCBPjFIHLocc4JXrwfDvRELM5+cH7tZN1Hav
4V61N7NdoKIt+NQcLQaNx9r81KgQfZ0WKRZFS5s9mPSbRbQpmh8/Ekk1WYA6
LUURElugc030wYQLeDFdYMJxWEduDWQSy1M8D0Xtst1gbeGj9xK/20YppEN2
vscGo00OnIsnxVJ8NYS47Mfja+qSUn4/MQ+mB9qyCNdgy0o6Ul9AlEzIGCvv
x/ZN7nMQb9Xa9zYzqcff40jR2gNNHInltu9NSI6oQZwk5Gdffng5pIUUPeom
4K/PopCkj0XerWCxnG5Q9amYkBQLLX6/3V7mUAEk6jH4rn4ouBYukVQX9ZSl
rwTA7PpHh9e79XTeppNQgdHF9CgoIEHhFR7fKvNc0+hmMSuPPr6DDgOyZhFz
IYeMKhZM1OMG3VdV6GyQXMHXEbBB3g1NGR7IK0DLl57g4RU87P3gtKfVSKDe
I81RCT/FMeQz/zpn3wxzXi5xDaft78JmqULL2FqSH4iMQRgWD8GC8OoxijdB
m2IOPqfwXwbqhqFopRrhsPiIBmZ/BcmrnHABhlf9vIF/1OPKytfvZQ1DelGd
kbbjTIZPqld8l05h6whME6LPzf/+4oEoeOFurjwAlqK9fTjp+VjbQlR6aHqN
0I69S4mxqNPFbIvIpzC88xF9zq7NB2YgAkPvbp8DqNk+fTzdnPZTpD104fct
dDsZ9B+hTCXH7e/2pfSTm4rShglhu8/g90fzdLkeU/jUgShK4upVmohQxINX
UG6IbmDQtno3ki+m8NjdGSemehy66l8AhJenGuFR0aXO8qTuY2pTvYOoBdPO
gbM8Q85RVCNXe1S/Xe/8J/rJqk6T1dpMC10q8jEsBBThGNF1kHtj3PYj4oJt
Za+8Dk15koMCSvvCy7zmIMFVBkcLIU8wO2/ASF1Yg61zDNxYymtcaWqysI+j
/T19G4AzvmvCxxHXiMQPxIcGIRXeCqu4XVua0PJ2YehsYY4+/q38L5prO4/K
36O63CNVKgQ4ktGu2Zi9ct5T7X1EVJOMEeyeslWAOSx2H+YVWA7NQQGtqHb6
oI36LTrJNNebuOoe5dVUyOZgQe1cfLp1wr5aXjyKBme6UOiDClOZt1nFNRPs
r14TP/UM29QCWaxdxkEPbkeDT3t29sp1mbjZy++9y6tL9WkQywJkNxU6REuX
gFh/U4FjyynCbyMOe7NApXn3Z+LilwCxIR6gE5p4pO0a91iLsHPs2K+3bNr7
B7cmS0CG1W+Jz0VymKBxuG6sa6gYpEaL9KXoJiPJfqD6wffUh3x/ObLFAFbR
tlHbi5sGcl8mSP5L82u7o3ruwSG0o1kcFUkNXGik+6lUe9pbOTId5EXqlZBy
fNTRT8BvQr+XRMGYtQcYHrBsSlKzm4aRJNTtxrKYQIfzr+Yg4GbZSl/VDwwi
tZ2iDOGE4cmT35mU+Te+Yzjo4yLVPgk39BSUg6Xpk287JS9+i599InE49J89
I5k3XUBCqPxgkhuCvb/3NtcvpeAd913XVVa3vfQuAJFWASArd8Be9QyhjxEo
CiDbHsYNVRWXzEttjVt62X4a933Utxl7DgPYNalzts2W4L7WXlGaeNzmoG7a
MRuH2VXdoRjY3gQI8+gDSZHsxM+7hihujlThEXUf92iAtbOl+kYFQP5C33Hp
vUuK9sHkWlN/G87KBZLGTjc6WCuv0BnJPNU0WHtUGSGwEfqmwMVoVkSrH+Sr
t7pGynVa7j+mSOmkaKpu9fPi5bYM4kQvvrDvANzIZAebIUZQUJwMoLui8ffa
rvLDMwtOcQsEjA4DQV93Zq4gSZlQk9yZW/3xiydkrQMupbAbt5G4ZcXeFqxy
UCB2kK1VWYZX0mxccOVjJtLXYtV8IT+9gxNr7lDj060N8ji5q2GfoFsOqIHm
ji2dUgmcw2wHIVP0/QGJBgzmrCCR6sXwBJCjy7Z47WSs4TYetxeNIIEk1SX8
gKQjf0n8b7PAWiOekhMqxpkXksD5nYKG3PSAbetixWQ+ldWWXyBGG/U2P0a4
7kMT5YG2HqWgFtHU3MRXZjDdxDkd+xuCBh/YMTdPAEqF13Ms8ZBZP89Ji/tF
YWOa1ZYfjpyV0rcvbHXZ94Nr4YLp7mcqZWeO5jEP+xXYlKQcmzxPPlaaugJ/
7CuiUz4k6oA09j68TGCqvBSve0u5Sw/nuF42ac1CtDObuNUDQqFkThf9+yAq
F3UMc0iNrO8/PZuDOokiIvywjcr72PHwBjgvg3oEansCcFWM0bNWTeBkeIPu
hsdiZUOrSPaCial2lW9NoNRHaJQjY3sfQlm+ZNzFHxbcTSxgg2eLHd6Wx8za
bL+1Zg9+byHiKRJqMLJpJwUhgtgTKiCMD0oM/+WvKN+arY2Ty8udHbqrG5Qf
tz0+abi4LQ1WKzrNCWObbCoEmQ7/jYyxcU1Xgkeh2mtrCqZrHk5lZJbXncpr
J4RaWUjehIUq9u7viqHuxxu+8TUjX3oqCHh5IX9sMYBzLYb8oyUwctG2gvxA
Dnk6UVZ4T8sg9KCEFHvnMl0v5RcVUGnyoLNzowlz8opkmcUS96x7gOvcgGJS
Ke4fYtX/IvBiUtHjwTs0TWbHQ+xvkx/jRV9YYgrUXuqldfmYuGgqmV6LFFAf
WBmJ92aMRkQjgP7Z5FlHuxvcT1HugkQVLN4ByKzMChhSWz8x0SuWMa4azkP+
ce4fDACH3/NAJcgaF76FT8/BycpFa8FMA5QW+36KwiVSwQDGJzYtttl4Z2ec
vI02FkpPzNxdNakCMdYoPbfbVYD1iycSK3Ds+qIajkA42dh/Z723VwpC/a4r
TI9JfpQ6XG343yfVah5lKSCYGmNT7oeyz/UlDbEJqZgHMMFX70StQWK2m73y
LRvveCroOM9C70vkYD6jyBpCP4PX1SuevOwS72zGFYNa6Yl5bxNgNAytYn4g
J7+B0fNjcaK38sgF6IkZ9oYoM0oIcHyGQk0DWQ735XZDlmSlCJHNFeLS7qXl
r23N624H+L5n/V1iSwAd3RymD4M/ahTgAwTqE1f1Ien+mY+bYTv93G5gJua6
wukZKvItBywnIhafhEZVZ4n/+lPWNRBW6BK99Z0m7AUWynXoCOTkd39ijSsC
Axj5rWganDcg3E2Jsx/cC4KflDnHO+KQY8j4jAAZHoeBkIlqvXO19Vpinvwo
dOs9MOS2tZaMwsvKAz1JmUOxsDuB1/LSasaIyoT1t1Dt4aSd3U13hP1DOETi
u96NYXHekcPFKcq+vtYLsUfQ2ZEhO+sLoAc7S2VGp5LnlvIc7QYPCKdTBpG7
bGmUmxI8M15Mro0ndaTLKHfpARohEBisvq4aWtIaXmhs28kLjATLglUtTEPW
z621ADKqxlPkXy7J0BbKSL3oh7kfESqTyBN58gUr/3sEWgf02BARw1qqUDnY
ptkzRjOcFQL+2wjGo/J+kyqoxp6/JPQDmPgDrIY1iOacpc87euWmUs5hyE6M
NlQL+cG8F/dF7VLAqhX36cpDjBTN0a14TbFRn5m9KbIsc67/GchPMUfYxfvs
MpgIR3gFu/0STV4uuegiM1G9oZhA+P65MlDn/DM0FMVK53qPNhw0OJ8i3Lqd
91RbMOGr3D88TXWOw+mH4uQySiV+V9PneT+s2s1zcmrdy2tn2fGEm+dvQJLv
2RpF2aPRqcJVvDgL1Pjy/Xb0KUJWfTYXsrOf2UStMmg6YE66wTic2H3OlRO1
/yuQw8mRxyad1Uo95I2uEEBdMSrNzEsHWSmV7XPdQ0YZkAkZ6VlznIcUaJvC
QUleZ0rOO1sdsnv44vryRp82+sVnObuSHAMjoLIE0hp1xVm83p/+oMUKXRvN
Ygw3M6b0gY6zQ2QTC5BLjNiuffjWQozpepb8z1ur90+Rznt5ZGoVvczEOG44
WndH2dMaStmLZnOiZMRtOEtG87qz10qTu6PKNqI+TFzB4buYzsGy2za4Nmz1
87bAkKFFJoq4Nj2ZCICCRpq57CXLPon0pIk27vBpFD1Hw+BFs30JnhlFLJx1
2QMiHy3b8zlAYt8vZzw7kM2NAA9q4ZkSoEYExC2KOpjv/uBQfqdnoSDwSo+9
ZqFDI7LMKe91iJt5wDxzoLTCfOG1tSjGlNQ851CATARKY1tsHkcoZfoYo3DY
CRHyI/MMCMHNPkHTOEcwuwqES3CF825VOsq0IvOFh5GrUlTOOW8sMecCKa9D
sSjcWPDmwwruz41QvDJVXTzgKQebUPWIINHl/Rl7kV4kARFChb5NY4NmgIQD
y8EXYn6XksMBWpGGvcM1d8ATa1ZtdeIfkLojuFvIxiHGC+ur7OrM/sTdQG+R
UdUk//SwdbRNJs8oXFIVMbtdyup2wx6F/V+Jcz4zuTREn4B/pM0aE5OSUskW
FC0ZGDxtZFlr/2gToAkmBz0bVq/wgapOF92yRaOyXubBKPMQBYSL/sOs3kd4
0b22T548L4oWjhxjI5ezHeuPPKVXynKuVjGY+shTCUpIQn3fL5WmKT+tY7Pw
ZJqH+kEhdPuXKmlM7Z65/84EkYWyW5yWnsVt3l5CijTVu6gcfg2z1aPvku7d
f3F1cMH1aIk6Qqbik/5IqTL0UwGQuquwvXVbwYa4w2xrvYBvGJF2mH6rWvAY
QEP3mxXHbLcKbsyaC6/0J2O0qQlT9Z197KKYnJPlI1FOfO0HVCypwiEcm/EI
QAHbZWPmnB1LriXNXbve2n1AdpXSQ8X1oKXvYjBb5GFZS52QthhoDK1FoVnj
aqc4AuCFeA+ydffbrhUW+S1fxX0elNq8LwJx5ajdnDPr3m01Begby2QlRhTu
G1Wl2frHYP0LKY07DUJLUMdD4zCBFx1IXqFa2sk+U/eXx7CyIBWUelJ4mdas
UsMaBI0oE/B5AHWaTaX3sUXWr3WR8hrRq0L96EidS0sRG5Tq8i2qRGa7vbLD
3ZdXw5xywiZ54bGDUpVa2XYVtH8QPGdXip7b+Qs0zk8PPlzLqIISXBpia8fu
Sw/8igVd8BDiNgbRgOuRJiBZnk8P3YEdXClDBsP+Bu+DGFt3yfvxLYPywYge
v46spVXuHnNqeWHSPEB5Dk+3qQh/oAZiULEYSz6qvqPb9DA0HXPfEY1kZ6AB
gaxuN+IP8ZH2Ir1Cq+35TTdTA0Q5RRCyDe/urVPhjnefgfaUlyOkClSR51Vu
Xgukukoyx/zSF9THYxX6ftd6wez4AFH5feVO2IOPxKvshznspgMh+GpBWBtl
qxAOWrc+VqrTJtuBTZLx1aEk2u2A7j23n8QLEp9Lbpzeejp3bx57of8+7gdM
dxLj+yPqrvyEFFWLADHfK0IoT0EFNXmonFedm1C+jqW9QAuaJnQLneL1r00Z
mmYbg5eluuoE4nfdHXYWNyWkHwtCh4QAWpsX9+LSdPKqZYx60LuRdjOihQKi
SgSdGQbBEp2jb7Cl+SeFs4RnteJHMDLsrcEWc0Jug4kw2vPXcQiYShzKZscd
37drGrOePuBTyt2pWcEavi3uzl8uHrnzdgrRaI4kQz4Lrvp/HinEc3T1rjkI
4jOIV/eaKlrgw4zTz9mR6yPiIzgl/KXr+t0yI2AI/vtwai93AGu+IWW9a22a
0RuQFGgEMQs+17ZevOBxmOe3sQpzW1f+7lX8sDXHAtTDaDgq2LAzxe/j7pjj
s4jF8R8mGRnKgUn+Bpl3nAu7MUYAGKTt8g809qDo5YDQBXluUHtRPsZ7DyC1
L+CzWE14aOl1A4JcU8QBWhA1H7P1PBycpRTKKOsmA+6CWjjMHfIhWfnmb6ZR
jG9C1ayV/TJ0VP4bOVnAwijryheKpRJmc2D7QYYc8dwOcHPBUGDOtcSbQ3RX
0+1TbhjRFNnEqtakBFUoyLs/xKP/VOEhEUG7YPOkr9O+xRWBJKvPOxArFXV3
MC0P2RL4g1GPcX7wYLf7pkgaADpdD39IWHSfAI21PR7lvm2/JCZ2zmPXNx2Y
LvehrmIv8JkSJwQjXtLxSxipz4l7KjFMIjD0UQ1Equ/M9rodlGJZ7O9wraSa
OTJIG6pkdj0zUAjSTYNJEKtqA1/Gpc68UZGu3GTAXMWbRn8QZrnFb+KcW/oN
SF3DUtQToJXvgV8tZFd1QDhq5IYweQuq6MDi7mjlG6IHcFxtL++NfFlDpZhr
ZazMb4kKXCISkejZ09X1RtkNTwCYknMouUujgWLAbhO0JIOW2ZF8sNgKxQDW
eTfAdbBHtKAxhsoJqFnBJYPI2ObXnu+aM9Y/4vGSemiaxVgjV8ZRA8DgUwIc
eLXLKAYI6ZM8ZF3OxW8bKEEoW2ra1I11XixvDJkZ+JI95auUe1M9TYHVLSbc
7u1GHSlgpPl4pQbrYYViIoVWTRuDyuB4+8cE363EyVE/KT3l4jvxbHL6maEq
ApMRTff4VxQyFsYVzHjqur8wahVKZ9lMXjAWI+QAnyh1LGA1CPWQFiBli2VT
vd1AHVbBFVOUbN9Gecso+1tx4qHxWcr/FfNcEvdeih9zf7S3N/AULb93s57P
QWx1T03gE3KKipR0wwtbsAXaV7daGkOY0tqCZDT8NIQyMfjvze7ofKgHa2j8
+p1lg9h5eVzj4h0HWSOoFZ3+x/GVRdXux2sXGYd7vRz6XFWCCcWDmDVPvW7j
AxUyLSFPaxsjnpcqHPM6PpK9A8lTq2WkoXejg05qY2oFpPkVzzV2wF2x6/d0
6GTjY4g1YkPk0PI5fV8FzIdmgnWyacansgSSOjZT8BG3MUN8Alw2v7Jba8RO
sFyOX2EdaHqzT2VtRw0FPAiG3ZxeftkL1pxhbVuN+vsZsCsqVeN01Qcx2qvY
GQA/U/eJSIFa6z3Nm96BePsOtCS3kuQNSJf7liN0Oc+xm3uf2FsG55KnBWfk
5Tfp2xPS8wf9wva4GsFX+7qx6R/urPB4HbFl/cqueF2qRoKBwDGgjaUW0r7J
4YBEIqryeOpKimkNosmOdcAwdbYXEeW3hJNEDJ/LvsCZUNtS6aV44ObInj1n
Ajj7nCdUtI+cx/kCNWFCpXcys/kCPpUtT86UtC8Rb6M02UfuKXPnn1Ri0Utq
Z0M38XV5RtPLkYtNWkYRZ/421q3PQcVpsPxHW9na/CLbhxc17skRBlStzpVo
/jo6MES72NmqbUIj9usDmqr4Hem29Z/kMfPtJXLNdlPKJ7mGObq8mcuEyQ5V
sUIReCo2dVqtzOa6eQ94a6cNbq9UotRovX+BEBo0p7HMoQ1YzZGPcZMoyWh7
MDxdPNoGn99OlcQibqO1dufKGKbipmRY7iHI+WmmtRzHfYWodCXiSYHnRJYx
uUZliliG3LhOqRdYqt1pYVnnpRMn2kvXvW6u5HXBjPjnOffOh/CLq5ddOqoh
RuYGBsMDvaTC19e4aHWa74I4hmpbegHVGXQFkN/IASZMu9JVH+PnSYE0xyG1
ciZehrG4w1RF7RlSe5DS2RcQE0NKhs7ST4AU9pywdimCRpZuJmY1BBkzl1Mo
JHNeo5FRp/gBqAFK9slt3JciPDkZprhOAQZP5lvOGJjxVbblrYlsZNaP+ghE
2QQEHnhkbPrDKGP96oeTBgeRvGVF/wBig3e47yIJxsJ2oWpgIYa4KmJZpSYS
S9LEgxhdNaIIPc9sY+A8ljUTAdWROTgqBnSRBAMjf5FPCeDufmtVNEi9E/JQ
DbsLlsrIIUMq1xIrBlvOkvdEx9g8iEJXjcqtiso1fSAU92cWFStGBJaAHIzZ
N6F1iTidunvNb5QVeUwGLIZvw9zFG6TwRIcCZTRhk2MgS/Chcdzc+4WUN6AH
YTd8c3FPvmFqB0dplvZZiaZjHwk37x15yujEi4Jeby/K+39Jg/UuYiKlA4rN
CjT+BoR8hxfPOkEI7/HbgHnDOsDvZL3uSo9BaGeOuy50jUyQZPFNtP74+3tk
0vxuqMrQWGGF45xcZd8esADPIuZpnZdMZViZTVYhLdfeUDns/fF0XM0DM37w
OA4yB5Vo4Bd0nD/z3prUSFm8+OECMnJC2OEK30f8qOT+oB1mtBMO1Rnm1GA9
zfiK6oWUocEggHUx9lxlCdwCiiMd2WBOrZTWjYouQkZn82fG3d8XjidNy6LJ
LziRO+MFgrUMCKsACi4/3QBBZcVh3DWuO/gniBEfrOISbr75IzXu2bikq55I
Rh/NUWJ2UWKr/aK0H0Ucgahan6ee4wD9RqAgn8P6WBTwTFtkZdygSEz1Igsq
LmxLYAgb6hLdBQ2iXIsZBAK5KLMtcF8Qpm4gSEFQi1QOB0xOFWdnRjf0x7Vw
Ena9xV4UYl+V5g41yeYRzAf/HfBuCeiMvEoViyzh6f2SOgbIPLkGpzQjU9PF
IeGpW7JQ5XaUVSoYqCv7Mv4TNlUQppSeIp0N9zc9VJm55WEvhesgZiysMgU6
OMuCJRWCXhvh5IJOxDgQIcvlbZf1BtidXY1ZJyaoHI/OhuaDNrxOA1lllIW/
Sr/Rv94y45BBO6OqRMTlwJzvff0qqV3VXnGU/ODB4hs1u+te6zwB5dJ5UPIu
VLTHal12O8Se0YRqOoYInFReW9a7kGc4baq3dIjPCF9MFotdJZnox2sQ3Keo
xcF/iDdc2r09D/SDYvmsky8085mJPH7FjJEqucLi9pxwG7Y/AAfzJhVIKO1B
6YLsvYplDNGphM80XUo+sAL3IjobLMq1GQTf6TsoX2ZA5I5ar1Czad5wzyLa
MwzKost4IYYaLgkL7rOi+RxGrpk8MOfzgDlyURr0YHQLRVVzB1ol1OftK5DY
jmJaBCLHXEibfrCCtACcQT1kp8qCJ/oqWHOzs24saU3jxFLEDvctlHvKognu
ojud9XkbBhE7ABSsQdlJk4hN/pNwMJP21US5So499qvSQkW3rmoY0LKswcm1
ppoyrGZ91fVuNeIqFljnFUEjxJM1dDU3LOTxEdtJMM9vJl6kwaFGxRUl1jr/
zxISyeCcJN+XiSucAKBaQ+RX8N6oFUxPq+fEwnvfRfVO9HTdPquAtQhryc0h
xQhe3prYpFxpfJXk1PDcKnmICVDgNYwQFpv7MK+WVB1F9ZLkVMDKhiLrEaDd
R2HiMBdsmztSzhFKH3IQlu2pDkMA78B3AwXppcv73AZ4O8oqV9X1LTuLON8q
AhpECYHqEeScMLJhyJeg8QdTZVlui9OwqD4ED5w96depb610NvGeJvd5Z6yQ
CxF/zOZm24pve6n+VbZzqi58eofnyNc4lzawHVkDhaSoLZiKWcG7p8E9w44E
9cjnPjp7Q1bhZMUsPA/3kx1nwXaGbqiRtFyk703R94sGOj4HMErjW4k878jJ
iA/X2q8G6ldkwDWI51uDAVWg+ozczDq+4YGo9xNX/xtkRfTn0IHxTL/wlj1J
2Nw6k12E6wBwNRlq6KmiTUVj/lb5IJrLmjM3xFf2yzF/YfMzEV0/osTnaOER
s17P+yy5G4+i5s5+rYsKw9187OJoc2V/Yr/iFt8SdNXy2esgVAwWXaA7eWii
AU3uSWQj3U3mAd7h0bR00SLJy3I7vqVb5/AKiaIebAavPv7IjHDtjtSUxeMo
5OueDoiSoxJdM262ZJiVU6lHyF8vQNqQoCbI39MaXyhAyu/awDlUC8OB1TMV
tb2ESfs8BWU890+GDwRVxcUYiih25YmqpN97wPymScZI8oGOUYczwJeT4wOT
5/as98sTP5pGVbzZUfCUnEVAEShWGKEn88d3IT3zH24U8GDReQUhK2NW46xU
WcPtW2piVMi2MsG8x52tDtUkjr0CFTpeyIZz0bg4vIyPbYi7gsE+Abmn5Dok
LMgCYdxX99sLhpsVHyCwSUJHOEbVSLjZvtCj7tXuX0iotCg1A+r9OXuNlOdV
GX6oA7bqATzrmYutMy3uX+focPwiP9lvVImvS+/UNF/nrYdnV/8S/fbQyOej
cmVX+AC/mxzB4wGGu+iGtanWD9S0ygK7Hz24kxcFXGFBCPLj9X+4FoGnezvQ
JdOJH1zJ4PIZwLR6+kqfW0PN7UcGf/BWg4+pdrZr3rh65NtgEZ+QL4/vXAS7
Z3RG+v7S17xmAwwfdaI5qOYzR6mvsgkJCfhoAz69lhCSWVMklmk80tIfSkhb
yESgL/nZbeooeLzHkXCwTgqArMaMMUAtdGcnP5SMYwkqtpro4I314adZIOPG
sqHTTG4JyNC7E7yenii199Hn1v1dTMvecFBtZ0ERE5vDJx7uWRzLJNM7QaFT
V0Kx8IkVUZVrpq6S9t3RAf7CThG6TNyIKxaE/6y5kU7B0I5cg5J9w0krUjlp
6z1/DTSal6FGOgPiGP3ID/8CpbBLtvCw3vKvfHu5lo6oVk9xRZjXjNiFe7At
wJxokWkq3TUQgTmQftOjltTkFVkci8gw+Jp3gft6I5jztJiV3O1qWHFNYxxn
9gC1E1P5DczFpjPnQr9oO0GdkfrPPBxvatUenKWTzMAWQ7n2TJ9VLJ/71UWa
NCXe8Rp6EfxNV4cBKwlXz3c6i1MUiN7C69A/D1vcZ5jF2MUIyfxMZU/3EdX1
SElIV8bJ/rneeO5oX+lirx0z96BTMIELH9yevEkMri3N10OFQNnQQTMxVjjD
l3mO4nuRl9mN/q9Bv2uYMlC0LaSQsJFIpz2NWuhLgejhDvxrTk7dRxqvjdrH
DTOB3hQA/lsFemijK3CQPkvpQNU8gZXmxaxn4lnXBzl266HTXgo1Q74aOu1m
szmLitvLowA5D7bRWk6AF8kr5xoWjqHl9ybp3E9UMFwOCSN+rA5UK4pucQt1
kkBWtNqfZFTBg9QR+Xa3Oi868zGZCDI3ShXFidq8GbicdYQneBtMC90HnUqa
LAOW9/KfeH4or+VuZzD0Um1oULploIBO2Kv2pBlafqZ+h6AFlZqz7pfCFKd4
6QNBJnxiqWYW4ikZzQu8PTLVJW6jqbwpBHTKqVd1ZyE+KZKostUsuRVs/qmK
ugxbDqwomzNfU7DVCn97NbJj8Rrp5PYZ25IofjKwcFm1YA7z9dH8LghmFMJb
llqchtEca5XrEXKiWxDYo/4WFV+sIdEbu/1NG8uwa8acUf1s9y+iFBGU4S1F
VX3CFpa+14MvvAAZTFLhgJy4Ar/IvqzirhgOW4baGMg6xtg3aDO+sJqDFebB
ET3qZWUzQ6sAqKjd5mUT8KM/UHAfkLjeDMaMHUdn9dqa3hm9i6YZ+xkO2PvU
ozg2prodT2CO/ndELOgfvzAm4vg7PlHeheDzh/KXe153Uilmvb3wQ4TAN2tg
Zi0EIFB8yw6AmLmyKnMDXnqM/jm7sI+FD6+g4gL2XcW9FHmP1yJfhnSGlhGo
Ne3e3M4og5ZfKPJqKpbLb2MF8C+XmX5FWpv/YP2059kSsOFqV5bdwqZtU/pC
s4nuiSWimd2l9k9Xe+yGnE7SUCFPj+S9dhekgtBl6NH0Ot9Xk33lOEr0+na3
jvivN7kj7D+GfXCLqHDIyrGswEdWt2/TvxkXqNp2XBWxA9ZNlqGl7Z7L5boi
V1BDC/rMvVVIbW9yYZOBW4pPoGKbS+dgwCtN8fCMItr2Vz7ZXvs8Dl6E98wx
T5c3ft3IKf87nwb666ZQXlqTGf0JyWzZGlj10E47BCVTgAs4oPGJSiAfXzsB
fd2athiPckFtoheNuYoqgFFif3cJ8+IVo7EYI+5H54Hk2nA7y4CoPWXmX7gY
M/HUCYy13YxEMkLwTkwWWCQoY4n8k2N523uzDtO9MQholm95LMJuCbXxYNIB
JX827DbMxC4xpkdU0+Vu6LcyRA/UBGF1UDcnV7LqTzyXEsX3S6MnLdyh9ayB
sOx074NSTolG821XW4kXaSeJDmXNOUvmDyRwWttyVOEn5noumQip/rgqYQB4
0Q6y5nDXPGU43vf6UDZXeC+6JVLh9Za55/0WHss9YAp4AXu20igPLtXdzCiv
hu7iTo+NiwUEMBoBj6pMys+mmdTiDzmtlK+DxeyhFUBF9BSutMdTk8M4254t
pVADRw4g0fJTi2t9aewPjdqkkvvyjw2A55R6vL05hg9F9VcP/qeN/+rPspD0
GYee+R0rBDgJa+guDf1GRkxdHeurBlQ42Q//3vz95VbolYYUX7xgNmcko1xT
if/jybIrT9r7yNkn6bGmdjHI5PAAxFjug/GICVLlYKlvnaIiteWYq0K0UNoV
B1HWoVIg5O/T3kCd8MaOy9gnbddNBuSVSAS+q7ZxfiACrIFANRDGZZX9sytX
Aq2yBk/V3CXpPK2jh1Kxr2hGYUCYn3b2VOukgT2ehdbwHaKtkRX61PEzSVdn
fdtKzAxpC7SwhRCss9LhNBRFK3CIYDwo+dEugM3iXJzlxIWKG+g7AF6Lp0Bq
oLi1XW+EolXp7el1QDMvcRXeMLBIQIBM0F5bGzKFO7zYeo97fFHg3/lgd18a
LWlOdavwSujAx5Ao4bvpmtO9xDyK41AeUDKNdVpfr9bdTcDThjfXufCZWzHf
VAXP+pjaXCdODbcvfSqiAqrxtvq9rE2v3CNX8/EhxB6Z/qscpSQ4fiFVEpkW
HdcPWVjf9bPS4Jk/18RBAFbw9waFc9MiWL2bLFYsnIAtuUuDuvhEIi0dJFu+
dEhbsRdf94U63gdG9tbhbMHYZaLd4GErZoGuZFXhnEbEiXOESOqNMq9f/LdJ
v3dh46rPy5EAfAwiTYH3zAp4uJ0yYRgvFqZJB6DT5xw0vN7rCtb4mUT/dQN+
49csva284Zg0y42LMNWo7Peiv33TtepW+wGAgnJ9lHPdxRlG5V8FRFAvJdCu
ldsaSqxBe0vxJfyvYubJKSY0v2HohmekK/02fYj3rIInsZbW6gndvbbyJaee
XsWTO+6Yvct7Xxw5U8dURPjfbldqSH7Qzm/RxX+SMLRcszqSZByDwRuDD4sd
9YyXngeHW4Z6Nw1MhThTJFgSv4lXQJihHs7iVNYUxgAWDLaeXFykFjIJ/6fX
QVwBi6fJBOPN7C2PaMqo7JAsW4L2+jSwzFXH2sHmY1/uvvjVHMb0iioyShYx
gIn8DVUTTWrUvNaxnvJSpzvRbDuhD1dFGdyA9u/SUdvRWtTW8mS+DcTqjG+S
rmwMq5uBSk8mcp8cid0w7DcYod4A/sA2t9Jp0mzvt1luV1827t8lh+pZm/lc
RsNDSJc4xq3kEa0kHfFn9wZ/BOQEw4jY+IKkCXixfl0lPiBom4jrvOmRt399
5p1VvKzw79QFSGszhwI8hd2mUvbYW/PYLDMrfjSOyIXu+PNx1rnJI0ssMoUV
0x74IWVtJlzuaiMuSHTXmBDpwqh/BXr5UL5FHff/9st6GKjD+DG775Ll7qON
q7/KQWy51/FG4qmEtJpp3Pii98MiAO/Lj7GeiJq/+NuTqPueXUqOePMa1UMi
DswsgL2CJP1/iFAQF385RKhiuoeKvHRl6fqpdgSttPdlUgdHU7lkv89fzrgu
gBfZYkSw3mkPF21AH2dydsA19+3Ziq3QmXXsDN++s6OMhWlmyYqmkhZ4PfmX
5KtT7cuskL4/QKJKEwxT/vjP/0GBk3TXGrHtTMejAXU8ZdD/SufCXV3mmfsj
2Kk6i7Nn3kQhNAtbgDf0ah+htkP17CnrOn8SMHuwb7CckWqSviyKOz6cr6uF
QbFCpIck+s627AS55gIfn6rnK8hyMExANomTO+RZU5wcavuHL2Vch4gz9wJt
oTZTTuKQU/NCz6mSE7LyglzKVkvRAZ3emqqk3PSUWWoCfypedKdBwwES3Jnb
FUOY1cFeWt1h7A8WkIipcEPj3z9NR8ZSy6rCa6dlirYVzPKxd11cRFjH+gjz
8ZyNM9NjCqOsO5AAwOKkp+YjYXRWAnJSTtbPoQyiRyKNLfSCXGHf0JURjvqS
yFo4BgwdJvv+ve6sTEBccL+8wI7v1TAXq5377ZoIchvDA4PLkJbpOHqqStfV
XV/sH14Ew9sBWUzzlVR+LwmFndTEpmR5odgV6v2HN23TC4aoxH2dtDJ8jcsh
63HnS18L1h9/sF8ZcYSC+wAqcJWqxRv9/QqcOjfXtTfK5bIhTAj4JVODTupL
wXcgylgBuHxO9QkUGB9Ao/nbnvNvW42zzwEPADOS5Z2PtwGJmcer0pa6fNZu
REc6VPL1fZYRfo0mVoGrDEJw90rOVTfT87qnACfLP+SNDnrjXKneKbdoiM2k
hygfXxCvJKTGnaJO8QnzRptpe/SKmhtR+mMA4Awl52oyimrYvdUJtjKSXaTH
ZLpEUY9ZlwsXF0kEF7l+fp+/Hph0/Hyu9f2Uv0remX2YuM5VQr8BBWdO+7tk
00fIpaMkAHgMwQlMU5ZVRc5o3w8RsfaLL9gnAY+6Rlrx2Fxoy0ZrJle9hi88
IW8wjpL42EwOSCTVV+GFOoWDD35P0DKiYelfMKc6pmnSe+XzFGWJH9EUUtQj
C5CMwVcZ+sSAKLm1vh1W0075ouNuBZMD9Bvt36mPrdaNxlcStJAoaV6I84Rh
UMh8GoD3x4p9MeXvCBgUnOWMZHoSMPXPKbnAnJCK9fyeTM/JoJCS+QpSk7dn
xgalFtJSSan813nAecRl/bx4WLgHRZaE3tSWgqyNnQAyIE+HSqLJRNHvkGO7
5UXKw9xNiQsfDylyGCVrOpi9Khx4nozZSBIl3J4w8Q+7yvmxKw06yPv280wt
NMQUlhBRRsbuUOEC1lbAAw1cycENdpTNJWNS66HiQ1pcqmTMTRK5BlhVbw7v
DX+9NJLYXw2Z8PpVGisWMcvv7bisZkIxC0cdpxHWM1c7XLoRmoj2EIqKAbmt
GR6Bnni6FV0zkn+1L1jU2GBIOidRxVxpy4spPS08vm+po06CkcfNXEgnqQeE
wD+Hp8os2IdLPanyZ0ZLLfngJ8GpQBAwUeLfV8xBIyZIt760uSQdqc3JO2Ru
Ft/8IKJEpGmfMFfcqenMy2HsSv7UwAm6bCOPZ6Mqvh8G+6QHSId7Fp0SMzXn
V4V6kNCL0DSy8bw/CxBkHhNDCJUNA5anUfRVMmZIG2NwNWsvZusLf5t1WCTm
NrDxXRA9eapAvwIh6fvxSWHNBxnzF7OlkN0ylbfGl1h3y7TSRjWNRJ/BEIQV
hGvDb/WaTVJ8BXZYP40xOzoNYWmBpI5snTKuOsfGbHzK2Hy2y8gJjjX3lYTB
jBvuUsPmFkE44Sfkd3gg6G7kSAGtSiC+GDhkfRcBfh3I4GF7he4hEEbiFqdw
CYEQ16eEbVIek2Wi8YEPniO4P2nqQ38DwH2kM0tB/H73oNcURazIbOJ8o12f
mVqbZqCPouYkfXe51BLBkWhV0NcYZokwzBwIGr2ssTaZWLkfTS/wVH1OE2OR
Q0Fx8ZcRZlMKB2ockiuxZQ01D03ptB4mrjpOfnYUvlH2h9PjX86yRlN3d2PF
hlXyKShHomCnQ4/78hqrQ/f9Grhfap43s4YFs8QOPQQaePrU3VqqtIz7m1Py
Ml6lYzC1l6RSWXAP8Q481/we6RSCM07J3oS9z5eZGIdec/OymWRwN6VzihvG
g8Kw5QxcirmXrlEubEY+gZawQmdTx9hpoj4u1GeXZJrstUWkkyDxy6BguXRZ
/YNtCfR9ntQlAUigNmRQ9wMHuWzIfAhOmLzApUhNbS93kPpdBU7lmYqBxsop
qKMB7zvhypJG4Ikou0gzxrlQhZ0LtEMGUP29pAUrXtnS52btqOdhX0mwSEoD
zhBzgGB+nH73Ai35iUk26yS8K963WrEdlILf8MG1gGQnsVTXJFRD1u9sjoJs
mV+tI/19KUkwAEJAWAj1sC3ygZ2iMX3T6QCqWPsIv8TuDbE1GaNYrcl/y3Yb
6zTE8A8Ygy9l4svHLCNGjqh0+yLvAH1cheZeS/Pis1dxvr6zrah1ZI2TA1vB
qEE/ixs3+bBubsBQZFW3ON/CC9yfGf4+GkeWBG3JQG7gCODMOdvnhiIGW6JK
t/Yf6lrE2vOLG5aorzAe/SXnAEWOa09DHCIZVucm/eM7J3TAWhTWIBC4pDou
ikFn/DlYzrsIjtigYEhi1s1jB8XJqRGHcP17dLdhpDD3/ARoZviP07K/1+m5
AaBSv72ln6hNv51C/c2dULVQsqN3IhxCxTw+jlssuEIl3Y5Za79MeE9SW3Bt
D0eLW3dwNYxs/+xNcZ3H8oi72qshBYu41r4t76QyIMlDrqooU+C9sDgDpNhj
qtMwv0gV9rOrF6ZPtWoejFvg+I+LRhnmaFgqBAb36WA35wVzkvFyYygWHfm3
gVb99V0ofruyT6AYxxnG19dxWuRnRQ3MeTXYMJb2MZKCi4C1XLsL6TwIBpFM
wgLwk5I4WEotjkVvj1s5r3JNa9+XHcIYu/3PkSBJZIXXykGPIecq4UjI+cXk
Dmgy7uLkUOxfp2K/cOWgLTN2DjWCotLF89iKWLxAeC3pfh9ZvwfzbiFNOjo7
nz3froXWVjz/JGC1D7//qcW7ho3wNktoMgg9dxsQxDPF2v53wuALWGq95ITV
0uWGTr+/Vn/i1+ec1a6jiye9LdmHnWlOD7ON3XDNFhFgG98BvXp007USVtPQ
TPYEm2eAMzl6jiD8hMUrBpsgMuan+RgLAHMuCpouvfXWkU1SHVZsKxtnbFL9
9eihXOwOknD+rgquKx805HGZSmXvKvEZZ3J73ms8pYVFZQg8J9TmHe1sI04l
Ukh5Y94aDW23cpvYdXCqI6BYA8mswhgqxXfIc+aMJ2x4j/NkussetuRsAzNB
WtoJaywnqWx7SqIUjqoGyckz+9er2OXTmOf1d62eNtw8RapCT0s6//L7T3wE
d+55YxWFWVSrUN1K5TmvkKdZJ3d+vXj1yRa4Z6jNfEhN0+9UgE66zKRwuD97
FZl5fe1eVnlSN5HeQbu/+FWvUA3DykLvVV5V98+mjb8BJEtOqKdtFykrvcUF
v8fOdQ21HFIBXmZtj1LQtdGtUfHfbLkGR2nc/oFS6Mxj9yKmDFjgkCAT66zc
L7mbFvDqTRDMe1bbiN2xVz9pwU090GP9FAfd8ENImm+8Awe7E1MprHxwSLyZ
XeV7g3oLg1uaQxWxujpUw0nnTZuq8BxkIDn+xb2XDk/EOjxKM+snzYTgqq+V
puiDXSkL5NjuvJMHMT2s/28DGodywG/vN1sZibhW6E3xTLcOmuN99vnT2MkI
VekUvmJawwCe38CpoAIrRHaCclxbeRVc6MdK1c5IHy15PNiFk6g+DUbRDKg9
YL5YKaVx0XV7GpVsrVVGx5O8dHuvHJkg3DEssgfeV1q6/GKOpMdO5L8FS81Y
ilQTNqIHuq7E1IBZTo1iy4ChOT/aGf8ebYgT9KRukX8F3Epk0ChKYtGRcEtV
Xg4FvyGOFWZCrkiS7U081ONOmN0AgMHehMUtHeacwgujRLbumvg/nhOxHfNs
JtzzJymKrSPqhn04Etek1Rh0P9x8WE6kz3iOSLbIDKJg0WNmoFrqTm5lR0lX
gDGXyJTKAMHO7u9ct6T1C0O+OoLEkJDFnX4DepmGsU1SutdpYP2wshRFLC8f
xWCFRYXaXdoXkLrsGQKbA5hqjAmanr5qg+AkQIPb8VP25SvTxMfl+xAaq6sV
aLIuCT+xBlx5uTk09p8QTYiUvxh/THc/bhQmAraIeJ1fQagDZabYVY941+H8
CJdzXG21B1RYryU4ehtSZJoJfn1IXgZM7GhV6hKT0hIwOz1b9gKHOvgJ/pKS
qVxuwUOPKFYwmjGm+m03r84X+dGTEhRmOtZmyKErvFn0+9zC78hQgKw9DENE
+Uy7hBg/FhSiUgsQjHiVpShNwvQ+/a4gVVfHKWjnqh4vfshiyMhg/6XsMu+B
nIpRTdusA5pWH4yauscloMoIlkgHGRieGZS17JLFahtabRsP8yzVjKJJgNCq
FDIG2jrE2AuHqrcTVxIT9tWOFnRD7tOHxj5/s+dgZpbffSQrxlTquJErfJ1f
VkpNaIGkFI1+v7wkYocP+YLZ2Y7OGRaMq3gWt3MSgM3ytY+bMDkN9dx58VMG
y5L7MpQkRWGMbqohOZV4IVNMEh2BmcXzmZJ8VIZqr6TM5kqcVZ2VAmCm6hH5
6Y8ptTt6DRPcuudYL8Ok6go1qfkObkqkwjacCcSmMqhyZVvF0f/qEmguzOzP
GPwJHu/kmrPKd6KqiX8yPu1rxiY/zPzmtmQIqmY3mqdnuhDQR188wqSJlYWA
dTyWyTaicmpkGc4xVKFMO/x7rMoYTqga9d3GpMAY+0IodUQ4+9hXiPA2xe+8
hqSF/DNkm10vuVcSUYKGZ+6ykkbrR8BeD7l7WjMdFqPYkheR7QCoSFfV05qg
EPPW0aOLdhZRRErMEhbusKoYA+fj90nlhTV3KuhbmIiI7xISMtbKL2mVE+Tz
ouQmo4x75YkETqPfaf2TNNt81BRISAS6IMGE2gl5I/Act/Td56IE9GuWh6+5
ombNTWhCyCAHiuFdDsaQe5SCG8C3JR/a1sm9RtNFf4hhmrIWtcKvdkJEK9Qz
rUZT/HtxFaDwqlCUrK6oFJfbvPZaa16p3hx8mnY47hqYA59sWnqWqGx/Um0a
zz1iwNtHTloiBRvsdFd/eQrJFzQ9JogwMIVoNUOSPx5GHEbl1a2ReRvohwkf
z5IP8G2SdYVq4yw6NoR/dnKMmU8WrgcB6olMT++CiNL5shzbDhIJdoymoL/e
lQSGbRQhqQESExFmq1IUwq8nEpyKDkjPRT7fyDRHhDY6/5DyGRW6NBfmmxZw
dNlWpkkt9kUGQrY8q6sXNZtjsnhK8qi/MOYwYJwmWMq/kP3HDtVWHePWEZqw
olx/nv/CnJwwonFhl0o6vWzmJxvnfMOyln+7lad028ZCvtOY9KjmELtZ5jWP
ldC7FnyHjpt3bL94RlyXDBtpb2VgksOSrHCFCY/kV4giTQNIt4kuoCUM0ELZ
9h1mgUl3MCfOJuiuTj9loDQr+1tVBNcuge8BB3M+WTLrUThZ+XwR+NnCwj75
2RAUXnhe2VactrcJqsvCwlahs5xjqJDc4fs3VEQGtjI8lQILlVN0sXAuJ5cg
WsjWViPeqVvNhUNDmB113jXeOnVShWOQ2rMm8A4XjcztIyEVB8TXksMhh1NP
1DHPx2f8t2M28dBAhyXSD4zuUAvfuD5g542QZoEE6FcLlN3rCexZGFMPF9EI
wjuqA0nSy91pUxWmOjANi/mTzmuscTJcwavTtoff2XyAjFVIqg55lWCz0KvE
FDAPbGyJq3FTpjnh8hfwOH8jwRIY5RSsvvqczerINt8I4T+/U2RePY8rRzvw
DYdcmiUC5T4vGPTzszY+8sNCsocvOJAm0FTHgYKEWyhZgSGuqd1KtEn3NKNd
D2SeYKqSDs6JEYe/Off9s8y/YIOQIBCVt7k4l/Wg5vu+/EHW9e3qpQUEZZ0I
292c5jDPWeClxs7Fji7cnx5cmmybzT5drcJrQGv5z04fKj3IShoJEUPCncGP
3sICMGqpLAZIBj5Eczw8pvHejPI1GMdCGQyi96A35Lm+lhsznvA3NCHCtlwM
kD22KdIOCUigjAez7Gd1w14S13YWGcdobooAVTyeA/Umubs+X0/oFo6Tpho8
gmugATXzdCl9fBefHRSrOfEyoEFlDBbdeaYooGHF2q2CQRDgFvHqXU/M2Fx1
V8bllu3jO1CHN6yUdGyclTIU/Rrj7dBvA7mslG4vdnhlZn0189DPdx8Xc/NF
4WrcKbvI0OzfV7lwaOi1hyA4bsTqNWWGzUBCxuB8mDke5kKaawn8vMMa7SmA
8zJZz9APYu7kG9NpENEGP8Nw3Jn661cCh7c/ulLAbYpOQfb7KkqxUze8vFZW
Dmb/kwgb1F7EnqGe0C5hp/MjDr4cGFcLbKapTWL8gYXqqv2d74RTrJSllcS9
kuNd3drRc7o9TW1sMAJ1+TeBm+xII98oN7Wgf2+41HE+eHEO16sVp3ivEZgR
xH6BQZVe0URbY3c7sorIihVhPKg+KMbExl42pKFRzXOBDkYfEBevfpUvP5DT
QJNp0qP79LdZ7YMGq1GuPkJUqgaDafzCVfqTlMoVAIobXiLHGta/djRGPPVv
hidA2dEEkmQbz6NnFy5ICYHgom5t3RrZ1A2fSeD/qqe+BqG6hXMMjYu0EMsh
R5f+I3afiBdWJe1nLMeJUCnM3zKK3w62Dr7e5L/qEt/fsAXMs+KlHkfXmQZ3
4MWlAK8PC6+YRRdiNBhtlhF1Pnx/1/6dkYEmmGm/hGIL8ZOMVofXI6bSUR02
ILfyqgyW2Tg6fqBEbPOKMldExRSf+nnTN9UsQhe9z4cHZ45D942uGtHwSzxr
KvKPFG0+HNc+Snq3J75dAT0QyULTXt0FKC9jEQETBzhuEASTnqNlSp3j2cas
YAvoGBK/xskrL0eZRvd3zIzgrr5QUXJNPBcEobUdNKIy9tOwX5XYk6+tpmYA
Rjyh/Bzg7X/U6xRpkRAGhT+uXEi4iZ67hK88gdf6/g7zkOX4HJd8XOMKTOGE
p4CJ7VKyED1bXjPrP1O7mLgCybpIKNZ1ZjfRHT4LlbsL+J2W5g1k7trIszy4
RTN2S4SeLFszZEnSf03q0yXupCxLy7nFfiotjp0x6wpbnjQAuOpFEMoAhBtE
GFtQaKh4oNa7NXzBSHcCLzJ1hkajuP8KYbME34X1x9R2I0yMnYhjGYnqAkI0
t53E840ay4kBjAgR6CkHUer4v0Y19r28MT+JNqpxcwfbR2iLvHiGvvP5mRUL
+/Q4GO234kvjE4OqKNTmzrKxWgE44feaMw/PTCZQNZAdAvgbrumWiD9HI+UD
alaE/QjywQRdAmprtBdUD8cfAUxp+RsKFA9CXAahN+TqzU1TIjvd2JwNwPNw
8Q2hAAj7UctbA1p+1/YDCwub5spId7jCsL1Gp7il1oPW6ozF/i6AIRsT+nyx
sgwtvITYK8GTcVUgnsFGA6yZ3m4xYPZ8vTfrWnugTcvCF1jhXniysLOMbsw9
vWwizWnR+abdYYBPieP7ei/FLmXFn/d5S4iL84bz3glQmJVE2+7mXVuROHay
Kg47yJCfBV/yDxVKsB1NDiL3Axvs8ERhxXtFJsoM7w/ojFqolOLfvxjnQiiN
vYI/vwTG37XSZrsUxGbtCx+lI6xddf/u9WLM2IBE8xiShAz1s0sTGTY9KhE9
T56gnKYBdwReYBQzeCxp3Xjsk94hoz3LXopeuepZVPIvBtPfrKU9VHurHzNr
Db62zGzeKHIVpqNCS0dI9AVrtETCbSR35PIQZpvTx8wVEcHHQvWwn3ib3ZVN
gAvA7cNrUo5diPIIp9hGqaz88lcINj6iu3vR7bZiKIKIB2X2J2GFRZNf5d4W
0YPbnqqfuLBrQ0SVnXy1D4739kt+kJskjnnD5welrjhCeoyxHEsO6FwbDcM6
lfTtGXe3FmF+VaCZ9gVbRPTT3a4U/cY9/YSBMfJEfUwcuoepFpRF9YtzH/ZL
tSq1WvfcjrG8T+Gd9fD9i16ZsaywPamtdxF9ZzjFhv7st8znbon4KKbwQRN2
F0O91b29JbVokDbIcspBVnTEYda4pXDzk2gVP0N/0VkoR9srvnPtLEZG8IE9
KeAEfoU7mq+6XNk9WlU7+7sFrTQ+szoke/Bq2v9oI7U7L7nf6RoOP8G1zuDL
s8kxwFydEBq2tDLBgO8mgl/0Z3Rms9Jwg537Hy3smQjnltVCxKeWWd3n42AZ
Ii8Tco8aAchFpYDia6baqyxkNkzJ1ujJFNYSz8DCfG2q0+LJmDwUO15+XzYI
aNw/YeGdr9x6QeqfVjD3x7Zwq5NZDpK5BVZTvvkGSDg4m4vJ7EOrYHspZcYS
VmgELd1Iin38BcM65WVemiQIwTU4Qhgqi3uT7Jam+U6eVtzY92JX7V17Tuhy
GAlUMDBM/vUOEBxsX5kAhF4oEdiG0vWOUdkOO5MLmKJeHs0B4X3NQxyxDAi6
2ddtqKPrUBDBlv8xtWq4dKH4VMenbswjftDn3iBn55CBXl9E1mPIj0LZWs6A
bwMM4GJ4t4sqEbT4FZEfcsmRP6zFz6X7PsCQOAurezp86NPZsbJys9sJqt/7
xmErGVO2tO4XLfzQO22x0WyxddDkqQeV7GoJP/bZ0Hi+r8CwoYbhL7SkxbK+
gnnOT66Du/UnVwhoDrwRx2BxD62Ua4iijh2sp+VyyitGWd3/cUc1Zjjw7nXb
lbWfIHQ4hPNDo2ivGvr4Ff0GhrJfQAF5LHIaXTtWjvcHgXk8agK+JqpNwVL4
kupmJimSoLJD2OciXzmZv53JHDTMLZXno6UOfXcQnGP3hizUz/PfiDkTa6wh
vSL0RtEpoc4hSNz6/HyObpO3bAlxZXFmLtwmWPKzwCB88aW7hOsYcEA/T7G2
ODDU2GZU2TiJseek8cB9iFlnM9azuj3GcsWxKVF0As8LlacIJDq5WQlxFkJW
ThiarZch8T+krZmNKOeZZsrPp+aK3fmz7jCLM6IKTIqb83k7cvK3ix+O00cq
4OsDBoULEifldZlVkwfF9AS0w/82LRpa2z4O7tfoemqeR7w/4UuNmDmnwX7z
x/INZowgP9vlr1iExEN9R+7Se57GXer8LwMkT1bNC1opaMXGZZYdVoI6VAWd
/ArJgp8XVU/eZfll8KshnRfx1h+LTkdi8swFrryxMWE2WRR8nneMJOBawI0s
yS1EL2TvKF3O+eSkyNIFU7wpA4Uxl3cBHumTDlx1n3brPRi1b4RFqopDdAWR
bw8P6XyPKfXCVugyODHVXtEp5ekwhXrmc+oUM6SUwO4VekDnDi5JbN+79rSV
46G2zF1NKe0kJBuvxzacYr9fMsbMQbMoe+hWXYbDBYBAIK8zuZC8K+MvALA+
a3ZiLoIQEq/Xr1QT/67ZOkiwEiAW4nuMC1N8lNTkdYI7UPZZFNl+Lvz9fITE
BlrMBq+375BAfpD+hX+u2IubNDvV9TeR+nCIRKuzD6SmqHxsheIPPP4JdQkC
LXT/C9stkTQAMtqxGQfhRdouli2OIh83Zd1XUmfJt98kx///ia0qkuCSh0W9
vq1w/uc66MjnIVuvHGt+wxHOzSUjI0GE+WlMrddN40u6aTOGRTOSW+dosuXJ
wM1S8wamXzHuQchaiQW6C/bS/tVfoOR+5tnTQJ7hdgorMgi3Fdug1iPzrm8M
5scXNav4xWDjoSTcvi4x7yicEt5aptyNQgb3hNBuSs17ztKCJTW9Poo1P2ye
K1MUrerJ9Y406mvPjnM3+J3O5J67fMBFgCqLY9eVg2rYpwJgjmBppYTMIwWz
waS/d8/5d2wi6aFUtnVsHcaazVPvPi1iy2HEn7Uv4ndZ++EX8cfvYW5kuZeL
ECpHd+T5kMdoknesMRj4FSZH26tXMW3Q1GgIJ9KLic+zXKWwB9sLmViwbP0n
3KdbzEvY2zyx5GWwsRNdmnQRcXTn3QbyoLTexgTIVTmh2gJ4QXjhL5tevXYF
/qmY0eTvA+ofhgL3d01eygPQBOxmmUcZKf1wbIT4oxQAiVyR/ohFYubtW0I0
YVtLg4XY5Oj8MTiwlY6ThO2x+FyL7DUCzBtOtfDqJLY3edAJlUcacaZ+O/7E
MvVFlINYzrDristeadLAef1OoBYTdLUotgiDncY1O7TDtqqAPB8FsbEWkBUy
27pJs7VUabl6g3NToRBC7y83A9EDCqLa7Xx94bAqBspkgynNzQKyRddqLfrj
BGJGrkoKvclLKkHZDIxQ4u5lNoZKAcw9Nsav0EN4aXvW03AtdTicnZBTq9fG
cHc9xy44hGLNuFqVyM+9KhnHWOnhAg5jDUcYY/QbiVseW63rL6qJ9aHvuQyR
1S9LRmtKlMBDyJNJHGPDJP72pHczPQbXPwPgOESmcvSDJXMQ3GpYZNtl3NcW
BV4vTxijPyQm6FAL9U37vzKOFL7BG3TPjbzxwneAJ1rBzQiB/AboWJPruQj4
xrkZwgP6Hb7cu8T61z/VnjQvdLJz5psL9VHiOkGVJmiCjSDS/vFmioBigNsi
7fCM8LQH/kbgZrjbtdhO1s/MrxsG0he/tVztAq+5sLTojr/rq2KZrdObiiNZ
JEl3uJDP592C+J1vj9EahEs/mduE7IFiC1tXvpyENf+J+Yg2dfhEgP3t9EzQ
nA8wAtLOk00iu9PopbjoPvAO3I3TdhlOrIGGLIHlPzFpQceQnLLm2vw4uWBH
eRHe1YeQNCFyTZYYE0BqyKy7ES4Hk8xDqOwd8MNCHd8oeKongoxy1ubMZg2G
a6/Heyqu9nPXsDrnYEJhk6ahiRCq9gkffooEzSXpVbi2MUh27ViNPimwW5TN
1aViVdIaYOp+pjEKj6039tTak+olNg1lNsV7Tf4j1nTO8C4lDm+ZzFHzSWyU
NXRNfBO48nxjika4/fLVbsMJuiVmPNuuQ1heAPyJeQGo8SPC33RStd4Tsl5F
ed1Rwz2QIBTU+Uiuwty4v8739wI1J6+Gqdc2bhfc4S1srDmos5xv07hFivcu
2+pkuIWTHdAnvydu2WpsHIiqviszrD+zXX2xpQuJjQTHgn4rdfWJ7Spwhd74
3LS1xqZOZcTU2otF0TmpOe5klDJD7J211aHsPyQnhLF1gZu7+Yyqa6H/922X
qiMCe5jKZ6Z5h8HnBmYbOye7tM3FtuDph0P20fi5kkMFpr5RVD6GLvzdkoLP
yvIiwF+0VSgxb4NB60svRoyv91KXfJfGH7EFiGvHetA6WJzGwWRMGfFXyNE0
XWNeKzzuHIH4HKJk+hwCN36DQkuWxo5FBVblJu1/XE2/2NPzuP0mtbSv/GHK
fbTAgUB5RRupNG7SSGTzLXCGUkCEzjCISSMUlFrrTG4aIy7XLikd3Q84mY9u
WHL81Gp2ytd+XA8ERHazevXruQpDRlUz+PI6YXWSzM5HT/EFRa1bPo/SQkVP
ibG34aKCBfpchMF+WbYraeJrB6A7xcF06E/ikuHb6eBtAfr1zGjgUNJe1ix8
vL9do6jwM3K6R3QVKDWQlJuUWKJ4Q8kkzO/vXAntZGcUxHLvLQjPRylatai6
qhCUxvZJWaQGTVE0yvtirvZqJSDpMJIFlmUjIqi/UqgHsCwwbxqojR4D0/eH
0fOtPRDNFu6CovTFXTgiNh9DVtboeonhr0SbWneCT+t0NZtTWcVcdDB3Dgk9
mPQSTAchLv5xFKeDiT3XBU9/GKbT7iDlLjYQCxtcenf3sq0ZmaVGLdPUywFI
P+M0p1MA0fEO7myiEy28a8X0buDXjrOQ/RRbEZe34zG7UqKQPJk0WMxQVP3O
0iyT51jcEPaQgl8jgfh0uGiaaqjLk2U4/Mc410psYOmgBj03A4+03eJvKzS5
xAK7Qvgk5japrabqqPq+KSzY/DlXId0k8V+8vW6+qvBdDivbl3SfFjJ8tCWp
j+MQOGrYFuNuu2vUMZWCmLyTjDOB3VrC7QM6lamJd5Xkk/JlQo1FfqzKPiCm
tbO/zlL9bUTJard3HY+eGu+GMM1eBPShh4ie1fosVa2JnScQDDYd5zfalR9J
fTd+Mknl9FYavtsgukM4cURjzlNmMhFo+ybUvAD18bzU/Uy9ppQSmSiB0ESQ
w+zSgGskO2A4LCmKQAKGTvtrKu+nzAJm69ijK4Aa1li6oYnft1YYmYRytqqW
eiHnRDpGGg6v1r8EyAqzTyz6waw3yObtAGqr+xKzX1CpNihfkXzihOk7pAW1
ZsrYnegc1+MelJU++mPyBoAo+Oqyz/w/jYVoLl2gHtUY1C14H+2YxtS0SsLl
KOK89ZvfydmoN1JUl3QGv8MVsmo0j/rQZj8xi39ewduO0sg6NodELptbQLZR
PHdZm40FMou1Y/Il7CgHPWn+8pwoYqz0+6SlYkJti9CO3y7YMxl27Vc4FVT8
3/EMsYjCXN2v/GCNnANI9xURgHKhoEeTCQo35RxeOffDnSR8xPF0CWw+xL7y
CzVt1JmahMZGUZdI3ZT+EIzMyhi6/WKozru2I35nKTlmDqHx2OVFFqMgdw2l
m/Kl1ogpGdko4HpJFRERDXUDC5h329qr8YJtKPxZ5fCTWuy5lOHwxNtCSQFF
XXXfkRaieu6x6VHpAqBlQl3dTqdIQ7vvFolyrtkK/WZrCe7VEspwJDpQu9Tv
iEBKIJ09BE2cPgb7o37Z62A70z2uNJZF7rKyBesudSGzK7d5Ig0McLHjRILJ
45HM6JBRZGEwRxiubhAGTejWSYoLqQR+ZBrX03YGKHXGhD8bnmlyf60J3GXx
jCNVly1AyhcwFkW8wS6of9fcg/x52UJgPeEM2qV40Bh6DKXNx1m510ubr2E4
+d8lHbaOwVzmM9DIHF6Wb4UVgFNfA+AUrKbJOB+3q9t3xZd4byTGJmcmKD80
LldSxnOj/uJB0K+rlbf79kADM94w6OgEFdt5cxNXgH7yxXCYe4q3ZVjsTmnv
bY7GpT3EYwt5gj3i6ArwgSg+ZQrfP5pSJzzCSv3hhWTfMwms5KX8pgLsyMgz
5InoFHEnRGSPAeRg8LJLspsCze7q3S96qdNtQFWuJYBQRXrwImCOOLGpawyN
HoWSnveVd/FxfwuWp3T90l7dfD/UaqXkgNFZmTovz1lkou6ahei51X6nYYq6
ULub5t9Q4nnC+/FyYbzCHYrxLzvUi2u3tqlaDIxqeuBcxitSTbfVr4BiycPR
+ik9YXlO9kft50npa292VxxnQog8wimVBK0/dtT/FWk5THevzkZRFPSLAXIn
JiQGgQDPJapcqJy+UETQQDGbthUSHDi90OQ4XzDWpICPTc+w8WZ2oDzLQ+2W
CyGYtb/Sta8W9ftsGi+vCYEW25MByPfEr14tjpCy5HkOCGNrw8j+UvATSvat
qksm9dLgg17YCMir7gWByywoTParpLj+mLNTcl8zH9nW2uVGbIEkEvErzpQy
rkchWUF5c1bJeSPO7tFVamt5ui0NE32I/C885BWjld0EStHE26Ab3ULNXP9u
7TNmrPgUgMX9ddXGDxb5U2tQo8bowtNLKo3dFUfKNo9HyUlFIlwQALIe7Anz
m4vh3cfjUfhrB381v2gF8r9K2EqOyyFn5Ug+xdjb0B+lY7YhPlYUPTzG5s7e
u52o33+9Flwhbv8tA+hQXcmEGMio++oCrHRr63pTnpkqKSqRIx1IIfo2/Ckh
bPlbbgKIIVntSWU9SKcnr2xC+qsVo1OLLbH8s1QV7S+7n/P0hKVHmMxIQxic
pAD8tF/GxQ4fnJNdWuXpkynpc2nYT9++GVEPzi+zQxU1ix+pE2hqX4z973mD
I3ruGES30gqhKL23q5t8z1c2hmM//UwVFLQRDbSig35Yg6qxErdkV/bfVHVJ
g+PXqdQ00IfvURBBG8GOsR4rlVGOB3Q1ID4j1fp6EvUjE7EcVb6WGYHvH4xg
VXe9WR+nBy1SU7l2zvKmmNQyg5a3dlt3Zb239GyJu2Hz9S0pSsYtODOZh3Dd
lVZLLi0Rn8PBukV7b6WmbZeamqtuAVrP94vwnjD/NuKOvpSOm7/5cgyftPYR
IU3rWOes3gNuwRMoCOJlgI0XuSyWldivRThqhoTTHhwePylbjjeDHxBl6JJe
vDcCz6K/CSjC9JEx6HNDqNm3t/b8QZNdDwhLResyBXmkZiCJffI2uu9Bls76
KfEASdG51pkSAXKR9wVNfI0sCwDr+HBsWSG940KJRIjY+QYKBkNDuXaV9F9H
dKT1s8dLwtpJGf7y/l0CNGS75Qv4mw3pzq10fJCFlyK23q7n5rOo8g94CkQm
mNVNcrJdzUMSmMm91ULqo8poeyRtUd3iegRuhF7bhXC9uduOVPeMZVHEuGpU
8d3Lnrcwhvq8MFGOnf8+c3H8OUmRBWZeSxESVfXmmA8lhv7RIRg989+E9ByG
aDjcdMnD45T51+147/bafLQ5L1IdKqXvFpmCULS7Kz0t+4qQ4L3vUxZr1obd
8/GDKEzsYWP4d6SZ9frIdzW+FICKrEZrTkQ+3HmXiUZ0ifj/AfkKQeXwvIbm
vW1xMa4tw7qrGfGpWg81Y+4LqBe6r00yZZMROPdmIyd5oM60qqNwOV+OA6/x
m+0kZ7YMT1VbPJ1Bm+UDK7uPkl6S5Tlc+NZN5c6OOhGU+75YnJHiw9CL1RRj
btgZWqr58xGZqFqNsiwVhcAaZPbKitryU1GWotNUA+yApROBI9xu7GFCYa8G
y/5frYd+AO/y99H6t6SX3LXmcf+K5XDmXeGuWQrh9/Z+JXInQBtOEjzHR8bD
KgrynMuDMLPaGFAsODF5nFGV19ZkKSm6oZzEOFJ+qvwnpdbMeZDiwL+rEwKN
NFLrEndjFkrRkQ9fKjj7IJUhiP6v5q+zaTYU4LlXzFFfJARhfngONzIytXqz
wlyk1RsI+ZXkZCt+10etJh6M1x7UVNyfAHewfGN1rT/gjnN1p89uVzFrMR0L
trC9eC1tznYds7lgkpeJojm5Y0HPlp0UYBKlRUQUbywpPssQcslnHlacvxxQ
xSZ5oivbOtTohqjMEEqnUCD5pplVol7vwMhTy8521IC1Og1ovkW7nb/ENIrc
fU9Tc1MHzSFCve4BLgro2IkgQSP+lmCDGYsGeQjsyO+2goggw5tIfWan6Dtc
fKyhDKmMt6mfgCwnlxHyQoKu4LiqYUQyU9Zo/9EC9x74YRyIaBGKw7NR9pwz
0QTUl1vRIx/qMd4gGH8pbglBpNfVnsQFHJ3NRk7Je7k6MAgqwG4GsmBCZW4D
gARfJ77DhbRxBh85ATdq8weTAG3h3SgNnypSZ6ujwnqpskiiFx4+qYrS+3d/
vBZSUFiVMhSPOQwhsSRlWKnEOUBQjZx3sb2UPbWk9OjIhZlC3Oe577aHkXE8
rTcC0+sRKUGxxjowrK6Eo1c8fssJyshUZ8KABjeGQR7bo3+YcVmABmNfgVgl
kLz9phyFl+5xjmS0aRA3GaqJTti17QIhsILvwiNKdAcz3AtDnJiKNmISHVBs
CpeLF+gqE731etV6fOs/EBDSqQGfUgpg3Vyuznmqx0z/3VqJHHZmM4A2u6XQ
7IMDgaKUhmqHv4TJKt4N+gBl1Ik4gx7W3DLv3t5KPSX/YJTDL4gAGl3Wqxlo
BgS+9yICofGh7iJTEzRu3Vwscntm0oFkjaBnpVOBXoSNdkb+g0pAkcAg4hAu
1aQI9o578eFVt1o6Ku+hHShdlUKcUSTUgy/8VvsOciu0DHLnS6Esl4Mq+mXH
1gkxLeVl+G95d+CVmahY9dAi8Zi/SLTjiOq7c/MTnhsCbRh6bv5iO830PlHM
SY2h00FQapi8XVV0KyVWhnmDaw66uAwlle/7XPubj4Q60POAxvZCnxVVcDcS
7uHKPjPa6ZjtrMPkmKbi3M4CY/JtH66nMtrufbI4OzMEE0vm+dLLl1R7wsxD
zBDRVk/WCGOj0xo/9ks+tgyBc2wxDocWBC7+CtA7D7ILus0PUVyaQtsV6WBH
pbQZ2QagS2WzhcuY8xa8yB3dUyKsF2f89+FzNooo8G/AiOCBAkxyT2tiKd5r
4KNKre4J+JmwbQZzKKAzVVXS18bCAmMKy2HANTtLanwWPn7CGNp2HCymMG0P
oaOD5gSq5X4+qFwGmPkBGr1h3A/Qm3T3eTHk0Q+8eJM++V252XCu/frdUnpa
i3ZdUptOhQN6aHoAwbeNBqcb9ehhYSwUSwDAZhBGCITSx5licURFlQYnZprI
Xx4QnA6BzuP5B673wAZ5B86Maz+Bcy3S5u5SswSRYhXi2570/0ShL5XsW6Ar
3DZv/80KPtCGN2uwhsA3q9Kj2D1m2oHMSJ9Wtzy6qUqXR5t07sLI3DKi9miI
JGQexM7QNT/Zgi8Mm1K+ELtpdfP61TAqo7dHk8IpwmTRSRbZKI59qsAOa8Iz
k1PKZkxz4qi4E2usFScyWpqAVqzsyJAFjf+Jjds+j/bPr1V5hlVa5Hu99OOS
DFWrQg1vZfMHMQqx1JbzyZnSRHipEdmbwAWEUyuR50okIhZWHVUZAsEVF40O
5148HCYCh0f8ZHwWU5KmVsmzHykU5Nk0dEWcPi2KT0tIV/rojfZArSwmnkb6
vI7pjmC88tKk+TNVltwIxkJJ85lNpdeEPDbJYP+kedKyaBj5SQg4mcBow9u5
XJbXhNakLKMQ0EVNeDYn2sX/U2TOUjrCxEtrcRXsapx19dEW2vBgymjcewqE
N/A+meAcfpNvLhXL1x6rB8F/j0tcc1aKwOyduARC1zo233sFHVkNhvQ8Hucc
iR+nJIYKXfVmjlkEw+jYge0wyaLEy46sn+C9Sj6XYm0dOCYoGP3np26DzdGe
DjSsA3CvTbft5mka5Ns1oH5mZ0dS/2vXMyaB2knudUCMX4YSvXV4v/P6JE9/
/kX7bAn235nGj6KJLdMuGOZ6EAVOLFWj/SEmLvrBaR3fgA/eeLZXF7118MzC
lST8vzt5k/guy2vJlo7yLg7lYmoRBDAL5LoaPUtLF8ffCt6s5mU0FMgu1Dyy
CIQMhryDqm1ZbBMMHEKCBXzoKJRpyW8Lt6bSX1mX9gmD3FHSKf5oTBhYkY0I
xcImyu/u+g276bUo0e9XRHAJ4ap/7SiyN2pZnz3ZOYpfPn08R+neA03caDFt
RTDuCqHjsvNcmMn7Q/3OLSxzAraa8ZLgBZjYAs/Hhj05q+99Tcv6r7BZPmDj
uJqkCMl9BGGFKMhZ/e75HeKkxXvgMJapdjIoFYTbKXWwI9nQf02p/TH3QBFz
2XNo4uBqpqT3Nn+OuppwwDcr0/qBLtF4avMP43vmNX4IA4Whw2837TpwUFLr
AJKlVtBsvqn10RzuUFrHHzjtJ8G2DGFFdXGq3jbzE7l15/QmNWw8qLFSoZwJ
84yb+0jLTOhi/zsPJZ0YF/yDNH6VlTB/53OzJIUfKpY0uKPNV8R404xok7zW
MulbzfTPmxx8LRNpRUMxTA/geTbgizAYUCnkBx2vTTIBxp9TVIFVape4mebH
XhbzttbH7s4b9gwSlNVy8hBnaaL0PqMoZopS43N686ZqdxYLqrkRKxV0Nejo
qL64yW09IvXFuuI6arexZdoCmuD6bCyzOBp+p1dHgrmdwdgcyJycCcCpx0Dq
8U3jBCGnT7y8YLmRUqu02nNHQu6Lzpt+K79JC9YI//kHs7GBIAxiE9FqnZPb
49btFWg2JN2pPMsztzbRhJOArqM8WrtS1WIBJbGdeMJlKKe8keGwEYbBO08R
CXMgsOcUT0SA7n/aOLKgGkouUx7OnshKyqPYWCRua8J/p25GVXObuQZhtEwO
QDl2LjxyUjQ4mTSPWrfjfpwLjtoYRCDMJgZ9TgBCjSinRoDD/eM90lBNNjcd
8XybrqGK0CJW4loNmVsSWcRxesDN75IRWcEx9fr0l8kk/kfUGsDcF26pojpR
GE172rA5H+eF62QfrDmLtPe/9XQI0LkbEvIcjoo99TtdZMhU66FboJpyi3iX
dRDcURBs0s+DsFt/04gK3p1qVILlHvVR5siUgS5bevxS3PSXZeqY+Cqsz2I8
uCak5tlfwhit6DBL0OswkoS/KoLrEXcOxeBaT0T7R7TG1G7+ERICyFiowSP6
vD0PnRLsrLYKfZj0FM79nbgWayVCAv9pT/4VaIaaHWlnOjM67Ox/cqXtay+l
mSfJg5hL3OUi9fdNYGilC90hMQmmjCA6HfO6jYQVLgo/7ezn2Ptw82JKtcc4
4Qd/E5ov5yLdCpUFmHTWJZVW1Txbg/pW79kJRI/Y/hKet6RBNS3KdkZds7BL
IirLau3Y7y4Yb0C+Wv1tTakFeDm9AR3g6vdRFGyI4TdQfTugj11EqTuUvDvs
COsp7h6//q352vLCaUSpWxQtSN0XUpVgPOSbdEsCZ/C2x2ao+QncA/J7lW00
ZsZnRo1NiLj2F6vf+va4ULvxVyP3d+bcGLuKhfQN6mbgr8F9SeAQoMT3TURz
lBLevkLXv65jEeUKZ/YdVs7rkcMKFWx+2rnRgK6TKvdZQrb4f2WLyJPqOOn5
6rGfi3NcJNl7w2Z1nn3n96NqNgu27JXMEFzk/DLYwcxMS4y7goJMbaJ4ha5c
Na2phbkzloRu6XT/c09AVTe9oQfhgPNz+mCC/33dwvakT755aOz5xJfU9suT
NlOcK5i+7tc5XdO6WL6SIGzOZmyT+IoO+88hTXYG95dNojqQBRYCyo1mXnWb
Lr4HtS2HF64zafDU3pNUwM5a71hwFGhyQITT1pGOO+ll7K/gz7UwC9XI4uo8
5t/PNY00vCk3/U1CgJ1L1RUPLfZaM0uV+tvIbuB3GDMFJN9d3RfD5HWIj75j
eOD3JTT5vfrU0MdkOgNtTYTOUCqOafWL14ehT/L/UrNOJaNQCqL3YkXAGWtC
QUAioTdG+x+WRX54bK+26ECioo4RY1MDxKoaO/xLERqhK2s7bQBGRJrzeVPp
J7DBVpSwzkD3SgyED4Upjd1rfM4dfViadxXhZDzFCQFUlktbNaADQSjuPdWQ
qF4gwg0yVS/lbBd5onKh06XA/HzraDFt2wla4v4Vo1EOQ/qhbqvAuoNDJ4s7
fBvpgo94raVd5MasHNCi2Nf3kIemeF+QrUsjIb0bFobx4hKErrkgBV1mJQUL
Ris/FhD8ylYg70eHfL0O9Hk9PbDtFRK+LtAwQYFQMc77ScZOlZ4PWJmje5jH
peTuGhwtCQjl6TIUG+hsF989zLkinAyl2fblCegIZIrRwbXW7vKT+DWE5c04
nQ15vhzIXzBpCRYSwFU+1sEWULePG8HS+HC8Yr/PJ+Q9D5h9xLToetlgS57w
SRDN7Mmz7b+H+zP2AIucTqIBX/tGCXvtlJNtncxHd4/7hXBoPvuFd/PMmdfw
G7ibKLsZOre981FSjfSckanfFyD3eih8fXKpce8FCU/40vYqPDexa8bgCgIy
aXKh1ii9BWHzVZMqVYInr91UYF42wco0sxkbZo4QP8upineKt/U9l5r19epQ
51w5dFCWPsTbs/i8I/DA56BxPep7DFDlBTpH3DjppVqM9bUWVmd77V9Y649h
KVaNEoA8CdDW4FhWz7SeROjlUcHoLUb6wV9so3XZNpyUg0GmVd6lCl2x2zEt
hU7tvhfWBi0c6hAI/TO3xYBTblQWR3YKN5Y53UX5SJ0PZq3uZEbp6RTQs+bS
bVZdeiidEdP44HLGS+CeukjO9COgHnoaNcY9/I2YVoL5bw5N+T5zSUgDNaJp
ENcJyJjVtsWuM8y5n2TZ/ZvhnU0gtCwL+p3v9ksYf3fEqsFOjc63US+2qmST
HbBEq1SFWD0LUNk07TKyT4ccwoSghR6QhXUCfH/e89wgbSX317y+0Okryl01
6wSLspRjDiP9MhjRY/nGGfK7M6Rx2ETexp5BQYD9yLz8jEb2VUw9FN2fUFyd
IYFqAtZZz3jmJqAsynnY0hYacnU5icJGX2jU6dv+Arg2cvi3du6ofu8cFSqC
xopS6747RVXLSa2cKpAjSfPkgEaCw6pgdt0GtkxPUrK4vCJ5SVHN5c0aNXCl
0I7k5Tv/BT0AoKOhOkE1HEyv+RQNTU4prX3y2i3wxlIcoptR2CA89PEDaiv7
pc4tIMTeJGw8ajP6CmzVHSxYNGoQismyNoqb6f4PGwjN4BMT5D35n/B0Jltm
nPWMeukE7h2RKDPqCxY6Q/w0LFEG9ZPT3zLI8Pq+pNsA46Y+mJkiuljpusUd
/HPxkOqXdwH1F2hwjodXwz1OKBqsBPyQSaAFkPw/MZGjAkhU0JIy5RSN6Dxt
2LpmgqZpU158XwKesk4ey+KokeMIEaj1+DjRj0A12O079yZu3TEUK8fI++Pt
lWurRkaYHci/w5wx1IyUDbyqem052m49lHk84DOEzLFyyD3tbOEHkR6WoKxz
BX3oIJRsf0hWNvLp/qMqU6CN8jdzK3t5DzGzDHzpUu9HhlKgI5aRGfKP9u/w
iZZ2RlHyRkruH1jzHb1uU7BC/pj0LMAf311Jdj49QINv4jJWohPb/QM2Oq+j
waLFntLelhfAAksjhagE7h8QzthUOB04QHHLIshu4qZLJ7n7KhxdVjdb5sXW
wA+bFs8pBlP2pRAn1DhuTaM61hrFjpfokXmeN8SBrcy94MtKesMQSF957WOn
rWqt5TbOfd0X9ZCy04/j/9K61R/AfKQZsjzSnieAiFxlDcpqjjuDEspXtN9j
i2XClhMMdHPNN99/01K8do6G1q+Ujiq+bOHyUqrfAwcfJbG2f6bSSwAUJr0m
1NnaxoDwVoyQ8pWYGUunNfS5ZESUxGKjlCdht1d5Fu2rEpU70HNLPMuqDLkZ
VWypndEWEA3CzAoWPcWUfuYGG45oCxro0Z7D0Oh4ceaZiBBpGtlW/WbwJVMP
elz53NQYtzP8lantJlemYj9nNsCxxjKlUmb1SR5jgz+Cwf6KTYpMTtNHjX6n
AfQxvD9BNHkf2LC57yof2y1ryYuiuZmYqV/aqf26pcDOw9Ph7Z4wB+1CznQ3
RmIFtNMkrrFmDe/hClXP6sNymlweWgQQ3Gc7qHNTNNkDaWo/gHnUR4CEX0jM
Vy8qY4fe97p5NBOtBsmkV+AftrwKJViKXPE1HGeszakmkIPOtC5EhiQ2D+OQ
g+P/9TaLeHdF5SrNWvw6xG377wnDMLWBaDxRrv2txnEbbjHpiFQD5DEXcK2o
t2pGuVOfapDCw1CEHZnKIpnMeKVMNz+MF6jJUTMGCCW8+GBDFaYEqkkaZyBp
etkRl/v5mz9uLvWJAQxN8KAqitapN7r2kb/ntjT+NTSIXR50q2qyaIpE/zr9
Zt/8aIUBXJWDyK+ai0XldNFHPAxKMCmGw2V3mWyoFypsq+/CnC6XyJfGmREA
CV4g/fCfdWugE+hl6JE6y55oD3jv0NTldy8ofNWXdBhBitiA+0QF1FD0PopW
0PvN+E7QdwP/0EjtXhAorTROWCo6PPH9cp+uxrTdaLc+0rIvO1Fgy6d03EmB
JvHYfX5kLBLn8zU8DTJbBNmd6Sf+ah58D+OBfTRhHhB8bsQuQZ0bsLhUpiVR
vg/zJGrh9Vh1RybtE2qWHn4IvFQZu2bJXylvgaVZiYUXftwuzJcSAPBBgd7+
mBHHo5iRjTMLxY2GyFpLWPi+jj6ywBWEJxRgDCnfMHBjtCVb8HtZKAyiOFV1
ic0h9y/wYm4X0wVu7uGGwCM8b5aTYTdC12jRqdyIC5/toESJZm/t2rvHOSMh
O5T1mbnxpQfX62IdVc9twTgObSn8MSwanr1JyfZDha5buZX/fYUM1qKlROnm
Yg9vKfoy7Sd35+xOJKpyu35rbDtIgk8CK7qDodjDxr8A/SqFesKdZgaFd2VZ
485Yl32RhSTWlex8R/5QSfkQSRfGfcfuObxBFFtuMo6emR9U0d0WjuMrTmVV
16guwDpQWUNhR/ogPBu+oDh2ChyHm7DhVcXEQbB6i/ZBO3byAJCcIHHF9ro3
Pkio8GfNQ6Li/FrY85hoOkGxUQ9Z+3EWpdphc4H4UWrOMQPjROmdHiwIT+Ze
1Jf2WAFqqUTwZRsxfkoP6PA2y06cDPQwNcxfT96KP00YxPpihHpCKqvnm/3V
d4Mrlk0kg4he/hd1F6Xet3BWJYLNO2qB3o9M3uD12CJbXjo5rxGMFWgqYhFK
n6B8z7ZCYfS8tdce+AP6QmqDHtfHQoKuOoy8L+6d4xbIlK95/fW5qwVhz0r4
KRnIqTKw7M0UoV++HQgMt+N8ozj+L0NGqqeNYqe/Oszfg6faEI9wKiBP7ktN
Mis8f12VWHz9kvQxfoBcFv+BvMAQPA+c/OKr0qWrrLpYbtOK/OxLY1V7VEMv
exS0mkyLkkmBSDJXqFsdLyGBYdeeQ77JTk2MshTEdcT1CRzhP6ZU72+CWeMz
V1lb/8ThEKKLah+zGzPM4GCzsBe8hOD8pynmyvjVUO653UXMIH9F0ko1At0z
WARnA8OufMYsF208LAnPmb3l3iae1kVK1Pu12bfORkq724Z98XpdNa1mKWje
EqkP8yraXYnNSjtleOR65Q9jDaJ2iI9ER0Fq5tlFiwsWlSP1f0tFiinWQ3Rw
L+KGOltubm1vUZn3hBFLddd/zzpP17byAhGXHlrtjSHbh+KoqP73svsh+nLH
N8BL2h5qvaH2oHYWapm5vPQKMRsn6sn61QocFO5q/NWnk8w0hJ+d5h6fr9cI
obU6wqpuMEg88VGnEwWd/JUVAoHzANCNa0K43f1dmTYfUVjVQCjvXj1NAvK0
pxoT4j+axDxVj26Pqo8cDOJJpIhNPJkoob1ZtKvsPs76r8NWsHv7RU81jdum
1ftJ+mHvahkccFLUzJ+ZdLyVCrF12N6FzamSm+uj8FWKR41UcTgianfp4yL7
rNuYfEa1HTu/vHaHUNmBh9Q7JDNePDnYfHHPcpmNx8kAmRJTAMfR9O4IrCW2
9vlR5AcPZHGROKz/19Sq0D6SFpoWaPQUJvnXkG0tjXkMSxgN9wewvPG5zMo9
wXh57wUPyfChnCyaj+jLXfpAjVpUURfWNFZokE4Hp5VXRwDgS/E0BWV76c6r
J4XjcWBGSATmjPbhVu0hQgnpQK1OzJjjZKG3aAas4gcAKitYTVOtQOo39iXK
FHQ77KOMVJMmadd0Udv1okHDTx2Q5b97il7aBHDgDEsbd7iW+shaqDPO9ycX
zpSz01SK0eJPpgXNYh06I7hdP0Mf2w9hKZ/9aw+KIod/eQgXyjQk/O3eO8ur
OD40dbjfV+TOa09jgHXmV03y8kkPimfMEUzjt+RTdL1knAlUej9opVJU3BjO
0/RiZn0Nx+Wxkyaa8MoncXGL9JGENbd+hLLKZ74F7FeN3M18urd0l/eOKTmq
XolmK4om2N6IZ0vyM3T29Ut4j3tw0GLXy3K0Z+jpNjy3uIiGIBU3zyT7LdL0
HVhRzFof4DOGtA2i3eHTeBLasYfXe/4cbj5fWlJz6mYT4ZLnjKltLKmss35S
0B6PFkRnqhWZv3HXJ54SArtejuz/FhNdudUahGPoAHCTJsMbyRZk6zAeV0HM
O3a2J8w/6HTpf2mwGNlJKPAUmC+AI8StbWzc7A4voH2a4IkRSS4MlVA6HTbO
73wPX41zQ6zwZ7uIVkk/ocHD8NaC9mCgssvpC6eOulbVeHAvavxWWIZZystG
9EaGyAJKlcZVf3+wivnKd5NjYUV0tJBEdbfmoCtnUnkyz+J3+CPJjrJmTqhj
MzxRLjeNDLymYfEmiW55+p5yrqDp6vgeh746ZbOMjdgFNMNPLmi6m8qD5U+V
tkFl7YIY4F1cV9+DCwhER26B4zIbd6T12ONMV6bB8X62lx4fOQrkbE2fZMyL
GwIZYo1aW9rT3GS0QfgaO4tcBrz+y99ks/BxTMrqDUPqYi5YDebdlpTRisqF
CvrwixD3VsjcPTtHOf/yzn1UEMAM/qScST0qzqGPGeRjONwVuKSX+Q481k+Q
3C8Cswd59IXqRiRqE3wm0LCrXe1HHTxbWu7FUzUoNIXD3gvq2fXj6b0aQf5+
gO47xZg8MByRqVoNrvHMZzlUT7GCNBKoLz9KHKPniA2D5UOabw5ero9iqdGG
vRBMSkdjXzCuKg3ucB+yL2Fq5t9XUoo5mMS03k60pQLwA+yD1BM/A7w5l+Zr
89F16xwYK+RX1Qeb+w9x+WtbDux9azRJrneMYt3ait/GqswdwMZooRYlJlHA
f4IxNN9X3P0XByW3EOKablAP7LLefxjoiGvYwFX6luX+kptYHltCDyq2QpEI
q4S/OaLiEiJbddRNrOYvbMo+Jbsmi42KG2/fPoX8fdIzK9fl/sPUij821diH
7GjiKLMiKjMn4PmOCo4GT88T6Cu6Ks9FaM7J7cC62y8GxDVODAe8qmiVkD8c
P1rY+DzwiZSfsd3cqV4C/apUp+PLpORFOrgXhv9zCw2Rr0ubBr9sZhpIly9Z
b8ArGuOqy2AP/cx6+5FqMI1Ck1xolDJcNDBn3PMKXwv0VM5w5fNJAqD807Ry
QBtZaXj+AW7BVKGURgdAgMgd14MFwOcg9HDqdWM3c6v8YnNz8kK5RlwP86yG
LsePPXLkGF4M8lKEK4apTjKNXhL9PnYFrpwxcS6Ou7eU41Vnh5B05PKmalV5
2AeMJFM02MWmb8K5nFPQpqPvxZs8SCjPdWA9tsFu91Lp3X1r77RJJ5PaCPJg
qsbvRfr3He93n0I/EOzJ90Zktw9JaYm5JpLyyGYU2qeR2YWmyN23Y8n0Ll3g
i6byT8Lz+2DaHQL/WCCOKNjmpCufSdH/bpb5IL3eLyOwP4pn9MCAd2SFyqEg
1RdbiKEtTiG7Hp00FDsMIF9QFbL1B+ZTXfSz73LW1C9xqgHkkES7APzet9YN
1ivPQmDKlYs+D4NhQyOpcdSiVHQ5KfoZczXw+YQOLuXzZdJ9lnPE5pgfiea5
xurlSmLXcrXgnPnpH1b1G+pLqQTNYiZ+kcd9COYW7Fiz1/x6YtCjGKF3qxIZ
5bJyA9c8OvJ8qEeyYM/HYhhbiIb+G9Q5J8Qp+rK8PC+sXa6QARtnxc9aE7S7
ktM5d1WcU2Mp+z60u8vkPj7bdGlQ3TW1jT5bZdcjjX3kQuvSTlDMAqJ5cP7J
4AqQfQ/35nHkt5b+/P3Y4+iHut6D+bnm6+WZKvYqSVGePH48UVrom+BSOluq
MeNDeGUjqUIWmNyF6vCc+9C0+L1s35RL2532Af4DBnVNbfLb6Thszezd4cCJ
PGnzmPq12kxAwS1AJCs1JVctlxs4LoGDhxBy9iyAVV4gotUdHKSycXHp1M0n
2v09J5hdDs0bHyWmk6F939rlm9rFajydHFx1yy8BcCf/gIMbti0sYORmsYbm
L4E35xogKElGnpBM3sWXB4Ep/5iE2bbV2WBVwCbf/PILPw5ssTQ40JGOVVyP
pNN/bjvpML+h13EOJ6gB8TlwDfHCkrDoqfbSWPyqNoT2YG5rw8CEPSWAbDgU
pklnadTRb467GzQx+HHB2x2D+Qhc7p9LGWi4IgeAzrTRTu3hciv8JJ3Nv1DP
lX1ljGdhiUZROjZS7yNbKiUFpg1Mmmougw9HqlZG9LZ5wLSyewvfcW0bV+Mu
ZAKpYdLC/mlLQPCTZMIxsVlqeXMGL3L/4VVOD7hj+oZz+ONskztdYUHFQXKC
Lbkgp+2ZQ/9zfGZc0k9cZo0ZnE+xyAe57yKs04x2WtKvAAqqL+qJ9iD0RsOP
EAezESA11bh2i59JXgx255mC3GaAGcv1LYTi9yI5KYP53i6mh1DDY/VZx9Dh
EXv/X+2CJ1fHwxL/vDC8hZ/mS4wc6Sgdg0dpKH9X0CvUOmLoba8RXjD+Klzr
Hyj37G8mhyzzE6Jw9aspsbSGcwNK4RJaVkDZqf+6pswUrquUwhgYpJyRYhVe
LE8UlhJN3i5AHmkKGyvpc9hd8KCwDNjPRnPg7MFIrmaLde6jpCqkkmTFUYJV
cH9Pb9YTwzw2LmHr/I31CRdTZmti8mTSgjCa8H4ff9ZtOGnncgo5Www2QvxA
cbzAChlHIedBx7ZjOObDIzdqUweMMgQ4DbY4ZmklF1vX0vqjokijiNLdiWGC
SCN2Pel90Pe6TrZadLmO6PySwd4aotwRIPnncI/IvEU1bjuzZP69JGMQz/iW
zgYHLcmMu0b9te9jj8ySEZBPOS79/q349xGQeRsTCMlTaKRoZ50TflzKxxQh
MqdhGM5hESBL1Yk3DYI7VeG9Ne3R4Xe9zDuwMAELrHg9yNtphQVKHmHXFRKx
Wn6gt5As6qGgXceumvjWTgBoRT/fiHIdCFQtYgQ/8HotGL+yZp7VoyyjjMj/
pB4DNdwO13GA9ZHEPkDCHgWu0dCYGpEaXMHUVyDwUDxd9m6EF1gXAKOJHBAf
WfCacm93NCLBnC9mwwuqXP0vnURA3UJX/gZQDOwKShPUDjqQDDZveYnQDFQ0
JG1H87UEvAFg0/2XU/PuS3KHnDl16k2h8HNRgHmElFALZJ0FJFX21/E99Hdx
ZwU7me5xgFHpqQ4a3kYmmapvQ05o6IYI9R4JCvZ8T6OPmrqNEJSNaQX3fkon
nXm+CY6Hrcoj4w87iG0MmY/Jl/8MPazov+bIcNykf+1oZXX3bk7w1dC32h9T
PdDpLmYa7EGrW8bL4GyKubLXf6BIUr8gtUGS4VtoFY5zCbRCtzFJ5Yv3KZfA
ZG5T4L0qPOUBOeeMliJ5BwaleRDcz0z8uug9zhjlJuW5fXg58cqambSrRfl8
8384b11y38Swcsfp1xe4TYNNWU08whCXRT12/bR9x6qirGMU6KqK/S63+FP7
481iSbndBA3OnujFYpbyfCPPrSl9rbVhWhv748p0apl7fMOQVjO64OvtI6nM
m+WVsCcnZ4zEWneEGdajj1ClzHGQRn2gD2IZ2H61JNkBEa4VNaxS7mcaKQnr
5hQyOih3Dyl2Fe5+3Y/Or3uruZogl9CJ9QRjbZWAC5GkJ6CwRjmK7XUHsTTK
/G7OEGJOGHh8SZDuH8y9oRUowHfZCWRRgdqBIlBsTeEn7MN9EohttXt8hksP
6lQKyLRvvk7ythsfdSaM6Pyjyaq5f/j4jzuLQLV4Ml15OlTm2g7kyY9ld4oD
+UlFSDDcK30YkAPwPYn22UctJWc5lJQQWJ6D0ORw3/6My3cRUEA04Mx6VJ9N
EMIl6Bslw2Zo4KPWoXxPa34Y0q5+kQ7+CK5tFLvezi8QHnl6IwuAAbEhI8rx
2Ed4s6NSeRghafc0eliFft4T7DrxmNN3weXJaag2maDtpRR7pnm+NGqjuuxy
kcWz7UqZp7/yH5GEkshUgsJNJDblVk1ttGF0eoRC5i9zwdkKlUpvafcRDvaF
LoLm22wxXF0hGpxvJyUsh3YCJtPlgmLRRPx8LBhVmnCmeS1YBPEFcYBswpKa
6WuQygOObd2LLlMb+mTHZnZlWzxBllA7j9pujCM4tV9mHo16L9k0OHzx5BBh
gLhF1p+jA7W03QiOtGWrP7+o5Vx+OkkdAbS89MHNFRMkFFMsgTHXWn4QeVSq
pig8vQ0Maebyc9uiTMrkEH+weJltYnUcEGuO62MTJM9sZHAmmLyOQ1rKEuXl
0rJCNIifEeroZwmYt4X+P6E3ziFY5IZO07jgakyh/reWB+TSxApiFQHVd4Ir
VrtgBEYxrg+tCJTh9ZR6Uy+2pZtI544X5FdOtpwplifWNstImVQoIAYnuAxR
IGF5lEddYvmu3BewM7pF+8W79gpN4OJr/Y5ONowRcRNmrnw5D5vO6d4NQlOZ
XzGPFBmkjeWqhUonlwVq/YyM/CT7A794i/j5qKwnXfUBlPBiLZVJHIgTyAvu
TJmqAMvPvsRPpP77rUysBK5fGxT/8X/J6/CPY6vhoV/+wz02D7Az8Z2Ld+WC
kXHHacOjLEc01/WnQEWLEzt3lQt5EQgpZCbkXJJUSWMVONby3KVSvRiYFhRw
UYItTov8ThZFnCTg9y0eF5UdKcpHCK9k4iffQ8LyyNAS25Aeru7DZ2EPahPa
VEzq26awevGKJR4fQARYUC1SCacpAiDWeUgYRzUGChhiP9fKXAiF0vXs0k2U
ZlApClokdb0Xfbgdyv4cy++w7ZOsVWfvUwK9f4jCMpJpxegBx/DrUw1TepAa
Ts2R8jyll4OCxxIqmGuqkPH58sCDZoUYMqN9cYLvv+yqXR9htMAfZBbyGjMq
t584aiTqwKULu5g1M5rbrEryf/3WIxVAn6HFb1pfPHV+VqEQU/YF7S8TJSOr
mXj5k5RGnV5RD4/u37+yfoejCzwuVqU7LT8rm1k1qvniTGDk/gPPb51rWi3d
4vVgSBMKnQ28ecptosLd74r/ibPhF4md1rZDZ5xULilM/bkDOCfvIX+6SqyF
56BsFlMTPqwK7M1b7biiHbEgk59WgfLO0aLFBN/R97m/HNisLVSAXV48O7Eh
vktGRMxgQb9XQBdeLHu23LqQz/fb6D06IXapetDaAE/Paq5L/MDHv80mkKL4
uHXbRTRcA4zqgzwRaL7iYc4/lig4YPPHS9JRw7jvA2BehGXyEshdLJRrjW21
m1qJOEY/znWurXfN4c4Nz+TJNvfZAZNSNwrbhlWoh3aEr5mEmz56Z1QU+k2y
pwAnU8CGZprTi/cxqHRP2BpBZNbsVSPSVugX04MHzZ4b5zMpquoJL8t5GYZg
/MYUdyRsKDHG8ET2TZI4nblh6oTq3NyLMUdKCW4ayz+vuMRFRNvxEu9WLxJC
GFqfxiBViUSakd7HzYOU6ZOwHspxKfQ/rT+uK6Ql9A9z7J5Y/mYT7GH9YTWC
69LcnD2BDLywZjnB9iKiMiYNt9oywMCVE/SRKIUL6ZABXbKD5+mFoW6CEQEb
6TX2CkJjtrhEHrkWaOO6WFhaemr23TZ4ZMBv7sQr5jhvh+JKo3TTc6mKNK6H
qrRpNC3qZ99RKIVVncYB/lL4taaezHqVs8lRCqNDqFItLncAKgfAIBmvF9L6
Ahoq8A/cYYaKe0J7469l8V9Ih2L7MUHkEH72YkgG17ipsRtgyc8bgIJdz03R
RCmKG/fbK0VwYWq/0MhWJOcqEFq3ROrxEvTWChXjvFzGfyMI0u8E1L1XfifQ
OYMjmgw0OdS5m/4EZCBZKjR0vwo+0AUp9MoCvpEEObWyMGoF+tujiFDXnuwL
XnHOBoM74L26FuD73cYXVFkAqvk+Re1KF0sM6dTfIi9dUcAP3y44ZBc4lvGL
POLqE/8w0J3vV43BbjYSX0+UeGAhCygUiM0I7fyaJSdC78U3iTSlE8gkEDOv
QrM4LYXuQLiNZF5s+geA9B9bVBtws9wy8C8ADANyCN0MUoj2wxtBvTGDdzC2
aFMhqt2Ep1SYD/VZTqLXBCwc3uYYhw3MeRDx/RYvXA0RwjyfjqNdOCoq7q+f
gbvt1ZQOa94ECe4sd/2DLXy/7dNdJSkjLXESFl4a9rn6n7Tb3SQTc+XAQx/w
A2mAqGCq2T/ZrbgnAcJLLEi4yzcMGMTKRTiaEpZmeCBIcigs2OFuUTcSajHI
nSCU7nhzZG4bKOqK4MMJjm4B9yHXunLdWG7buwnZDyj7OPjUEM4gS5mzxJHC
SdrEYOvEUVAFhc2PPOZIsRcAUtb9ViA0jSbGyFYczaEDclVi4S1p/Y65lxrw
gAX5/QoFdQbbnpxTTbDvChPZXAcq2un2upWlIiVMRILUV1mnm7Vu+qyUpw6Z
XjqaiIemA/xlmkOlXQd0rz1LIx1DhnmGLhxaHIfIRoceX0qzOGqvQj3REaQ/
NOO01gqlsD1/sVqrAtHdjm1S+cX+nEjL1AvHfnqsIHBZL2V36bA0tsbT4O1j
kKYZwxHwx1R4rjlKGB5q3XN2uRvlazPhviJJflkYbh3IkaeNW/THhbbYkrG2
/2T+vzSJJYfttyFb2AZEiIr746uIg+uZPuwZlfkAl/v0qaX7UZ5hrsjro3cc
tGXxtI4aawEAsRuTC/IDr7mwkpnmlvxe7zJmxEFgNNPu2Su6Ocm5cRr+xhas
U9am8Snq5172w7H/XD77GsKxcWfhkHd2EFUIAJd46/sbZZcrpNdLTTHdYuqg
5FFeUh3UZ3OmcK8Elfz1+zw4BGMrYdW9aLFlxFIJq1l5Qdasgl+sXOVFkgp7
Vg7j45AiJH34ogTtGvWGkLKLN3+ukL6ADwlhB7dmqaCNxkpgkSijOD1DSl2G
WHv6Hyu7hfVfgkwCz41JBkvEZ2EmwGF9G3+mPt+6CPCpqkjUiYhJQSkotW9O
rBhFeeLhpjyQJBK5Mddyu0FB6n2isvvHPD9ie5CVYvuCXexCOYMJyWty2bJP
sYW1kwU37xsZAec4pKUWUW8k3KcRaC4qJ3lPV28Q4POLG228U/3cUjke/K9M
p+OneoscpwfCWhFn43x5ZZHNMDvHw3m90QLBPaj4eqVinyMceH2chzHa6P/Y
g6xv70Ki+L4hhXLErqU/ILi6WKiy3UXqMWR7tHrSFpHBAcftk5/zItja9lg/
dEgtOcnQMF32/BA+vcBdyPa5hfImTMzCvvKyCshnB0Utt/WBz/3QASKQuZ+m
KeEBAovJdkbXI/OVhdNH7CNuSGzi3yxMgz5YmHuKGvpDAJgy1C8WOBTcw3QU
7J4EfPOv/JM8RkIn+8QZCCeBwyEFQXOoKjE5F6rT/pZfei+njV3AWZj7cCCV
hQDcRZXcVVWwBHXAEC7Mubl38hWwCrHQwmpa1Dkidadgag+qrEhobiAxclEN
NNW3s7QzVlgJbNOa8sgXP5rtCOPF76jsX9TuwCj2xkauqVRhTqAieIBm0x8g
sUM8Lo1mRWxx6lK/LDnyMXdy9jqYE0kwD5CxkNLGfu/P/q6Yb9a/DW7dyyGz
KEMxMalHf+bm0IfD6x1W+pM/1UbkjTBSdsVu+8EDpsKc27PVLT5IMe01E5X/
IXQ1IOcpvzC3UUUg+2q/SDoRvuM33sFVjWKKh+A9aWbWOcpvhkuY8NVXfgpy
AzFV6JKA4zxf9FZkdFtiiAem2i5sh/41j5gAZPso0ly8gHkh4i+E7Y0JxKMw
iETmx/nMGFVYhBZa5swFBVBv1OHAHsvX13Fu1Q6/Lhjd6UR5oK63SojlgMIX
+aJbw26yQbuYuhj2WOowsicRixDv2xrYnZl2OZst7/cVDpiAjsIvoNws0/fd
PlTUXSe+2MRKJg47bBEMv8jYNy9oDqpcd6Qmho3aOQCY0PqntD2orNIaTWAr
L3hgR2CzXOuIPChd8gjlQO3OdepJ9XCFgRKw+PCh0/3Ak0T0Hzn30pRnPLMu
ek8iz/ydX3NRTaRXfT3el8z43N32g90xuqYFXPAwu6+5r/11D1zzr3TS45wB
Bqot7wjSnF2zbzx0FcqWcH/qK3r3bzbuzEfTb+BJJRi3rAfz/gVJtA5IWs26
Ovd5YCSEbkuAUnpOhK3UsQfcfFUtg9dE56J9jWNNdRONs+fvl4oxsweNvs5r
KwXGaY8oHLVSO83K+ahH9mHzgUK7IrFVKWz93eMZOTJtfZ/Lm81XuT8SXvD4
hw6KiHq5q1K1WnUlqc/Pfm6P0WZwBA/8AxjkgTCyDGHvgc6ccLoZ3GfvnW3q
RTHyMQ0YCgi8ELADaXumiqD9Z5x6bf+/HUtxnm2nEJ9BrpCD5TJFqKWuIsrT
2q72kH/vliYuy3mcalGfP8kBcOXlRiY2giYFcBDTInksoR/B+Avu9I5NU/5C
pCBxByBYnEG48P748P4CHCy9FvNDQWeKyaI9mtrK/QeZYzfpabnT3cQdKcUn
Gr1RVPxvE5xnuoTKLJNHI18ZyXVuE+XPeajlxawohGbQzwTOfQbkSrnANVxA
JTiEcu00jJ+4afIM6eu5eucqkJHyfROPn7jDqvR0HZ+aD5JgmmjwbeFKZ/dG
fF1ia3BbVktZjijk1SWaNsD4tj/B0nE3+z3rZ40sE9ls2uRyeJvUINAj2TM7
SlBcTcU3PviHXgzQAwI+iRz3kWKujxI22UUOThDdB/3EO0U2qKL4UXzNhzN2
9fo7AJDmO3kdeD29eTS5ptf9x0HiULcyl1TiCimFxZnRfVuNbMQW8OhmZ5yv
6gfJS7EjFyPh9zcIFukfGrRXEaiUaC9w5fFoagGtWg8mKBcgPpKRVfgqOEoc
EovJiM/iAGpkUw3YC0eayolbfdy+/nY9nzlZ3wSb4TPCn2RXFEEo6bSIwElJ
5ua3p+efeWuTtHCmwsF2tPQJYlbfMVmxa4x4voSBvtO10TNFis/QcatvJpP1
CMCxfZ2gtgOby+IGE4dnBa0FV2A9H2hn3Onuuigrj8FJ+AwVbF/6G8Um8PtQ
2D4DY+/qE9RCh2cs0z/M+TgXr/jgOnhdF0EAiQQOIse/eXIAhtBLXUPhJ+Gz
SaYzM+jt8iWOpTG63X3IwkY+3tpYl+aifT5GkvTYymAzonLypgWq6ND5Nd1y
q1zaTU7zsjrbLt7b5C58KZ15z+idIL7h6T5IwPprgDQo4pBPuXAq/Nbf0mI4
x4BAPlhpxGKPOLwhEmlhmhjxwf8flpoat9QSnvJ+3pkrih8xzF9SXxyvfzWI
k3d4IQwKWpJag9HkixYeiui14pQVMKOHGky8RhtPTKPQ2YnYxUrx3LsEKSxA
bIzCbdkqtvp9IUYtv+78J2MHFz+ICsDoLuZ+lwSzFmQN+Fwz8DSvwst6dm8L
QFf2n2xQWUpH86fGMkwrnnVmXopvExjaeZ+ImX1PRpV94Mz9jAEd5CbaY44j
0TMHC8L3DDwMnBuM04E+aZpaPkdka2FxbVRteVEzdT2EIVBCBMKcBgkajDSR
rNLyXnnRd0zZPsBMTJjESjm/ZYF2ZwU7a++zAbP7BYWBopOQHhlDsoEjq86V
C8XuVVZNMxVrGInr0djK6hm4jVrcbYk+cEQiDoxYXXoTKwowYbgs965QWGKa
ZoI2DWGsmL664JylaBv0fYEDhCBWc8ujXVunEieQ0tSCZj90iPzSp/3FWRp7
4JbV4jo63M0MXwYozN5xDLnm+/VNvRJzvOwvjoAbqbnSDw5Yr8VFkR7+xPrd
SFW5UEDqV0erOIzgArFWqbhBhHxyH9k16iplUAwkD1DG7SsWVaKOlFkmZUQu
cj9afBQXI3pdWJcjgV2zUO4fHt9NGQ+U1FLJye0wbWp42szqfCr2kRjfGVqw
ShyD3ueFGpxWJq2JRc2s9ybQMmwyGHVqn9dId+LTfysnZVTGG9NZQBaDMaAe
tLNORDCdNABg4vEfDbQcSqFSKL2WdPalsAXWfjc0B08Iv96MkLen9OwoYPQX
XFw8qXKoblgJILLIBB3r7Vnsx02xxApVRIFGBa2Vu3cfy0DTIv8RBZQpb9o1
0UIReFXqZ3JPu1zlLdwWYJSMXEjlfPbjWrqRRr0pIfp1hgM6hUKqjB7Nyfk7
w/Tn7jD0l9LCyvgJovlM+KD4FEiRUJ/WWFna79pvr5hV+zDt3BbRwVMkp0qb
Y4CImeR0Kb9LQZj5pE+KQwm+nLc/d1JvXyTj4pMqylDLbofk1V/9odi9jaoa
9xWAq7at8E0dNn4Lz9KfGOvc41QKMBqVknJ8QzFiBwWLvx5zWt52Ez3hq3Pk
aUiO6bnnXmANcOCUVmwPrRGWvST3rASzYyl8SgEoIucCJ4nTkRj4lekefrhh
u63XVKK8IADj8MHc0FIfkJLq5qjsowrVyebN5TQvcY5rQuWEaXwbO/FK2zu0
YI1l3N7PkMpg4rgq/PeHiQBUbR23uwpN5+4S9nZT1aZWlb0rimqXkQ/+sW3/
Xao8Ql4BgGC9tWeakydAyPj7AFphW9aup5BD/1kWEG/IRBpS44A+lQTrMIXT
UwovOlIsZh4LFQGRzwNL6iubQZy0g0rMNdKsUle8xVGj/MBkYRIbgm4ldDnl
c/6glBP90pJE8YuUAakLoMd/OZk3HLMSD7jo0SNC4careKYNsdpER/q3I/3S
2LCMy8RR8dsGs6LcbUwzKHuulvkodDPYvowTqZsXPV3FWT0J3ygsUZeVZJCy
3QuKAQYknGBwDW161wFKcGR0zvRFezsLXORETgwc/Pdz5scew/naEgbqRYVC
vf/Mc3+b4MhGv1f94AcbWQBNd0remXt+74co/hMIMhJN4T3jFLmM71hXLb4A
RNpqZfsez6vlBdgj6lzwu2gCfoE5jML/rE1EdUdeW7K981I7oP7U+vbdQibp
FBX8WaYmrLkeO0yGsrjKOuiIMYhk6kBhcEj8A5bA2Gwd7+cvVEc/aiyTlcEf
Inj9NjF0hMaR4fhGw5QowcQ2PpyK+ucS/cNKpcP3oc/a2ZCaQCR5q6noH3wa
UpxvtwFr9cO5lPdajL/erVuFdPzcywcaeE2GvoolweAoL4UJEHcP2jrVOeeg
bZuXpBCEkGU5Bv/FTgAtksckJbYiUv7K0HHPAxIVFdWpnyOn9IWH+nrMwA8V
OiuV3F1S1snbK1tylTSo8RHvlEhToYHY/TqyGxzTWDoHSEExjfI9b0tU08i8
tP+2w3hD/X3Y+Fa7TN2msu2Wc104aICC4+XFOghyETU3KciZ8A4YIDXmrFnd
zz1srIbpcjZKB0hoqmTZPoEU8RWWkS7BU1Ms6ZRGQ1NKRRS9oupMC7fNAHtM
HAmGJIHpsRS42p29JCtfeTk1s8nmPc9L936qzdrKUMEPwU9RlJaoS0Ro+UhD
CrECdvKpBnuKOrUGW5sb+VLpMy+NOTZRqhoQICV6xAEJ0IcEnCkxjST4Wd3W
5BGbYaPRn0/sCJ9e9XaFdw5JRRK6kOW4syoic9hobPKKYFbybt914Hom4N09
YFsTw+y9w7JxbBQHOSfk21FSypdksfi0px5z1NgyZpQ+71zJ7jcgidTZ/K3E
wEdrf1t8xbChuGmW5I+7rwaC5wfA2f0huRPAlVLpe+fLl5/5dDH7i646N00K
4/f++35h5Ou+U+Tbbtp/0mpJB4+Zp4TWzPcKbfNXF06OVO/LSv5YmHpm4czY
ABC31CkSdUnwTqiteonjA+6g72xwcIAuVeGVMba994BppLkWKO70h7fLuZaa
VRWfLxbRqe/9rqP0pSyf30JxLXg4s0pESjXq7fHBU4vBPYfVAqaGDtHXR5h1
ejV/mQWRAyoQEeopyy9BBTgwzKuAogFErnFDS479Zn/wjqK5b6BKEJGEMj++
W4stUU1apXpz9e6kiV+9/VZiOu9Ac8ZRNqoGeJwQqelsGy6QyT4wOEp+rQfn
kdWwrTMqTbeqS6LXofX7xmgIqowtX81EsFTm0hOVTn8tIa0thQZHQWA5oSqt
62rflAcDJZr4PpRZ6d+YcpCbKRqUhd1Wy9KJpZMFZYYOvmkcCsTpEFhPE3bR
vk3IwqnPqcbZjMSra9lO3FLv1L+nsign5o1nFY7zqgAcremUrEf9o/pZg2cR
cWdG5q6OJ/KZc0zcejOV336zp0ZZKLLH6nr5a0w6BwfyyxQqy8uPFwrnivhQ
NwjBabBggAgCLeYkR/jJ/rAJz6L8QKktWaKwa94GMaGnD3JYYb0jFb88fZBb
dsU64sf6jWPW+h7QZp3W8Z7+toH7wXer8sh6uJaxcbpbAGacZq+JmYm5gLHQ
jOAu7FPWyt7FQR+rQNeG9CNr1BygNOzcwEOPwZdlIUMuXApaIpXxq6nMEsYA
A+EdCIXPFW1rJrA0rMn7nHhe3Ujh7IrTbX/UF8F77flLgqM8k+XYkiDcuy07
mI10kg8khl3WVtLqtut8WtGkEklIeX45HCPcEK/YjVGLk5yqm5xpYVSeyC9m
M5AzUPMAxcLuxcHXwWTkZKkTxymFcJJhav8erX4Nr64Ijn0rOZDV2ollg0e/
TDBZDVIYQ4SSKNoOOp2R0xudxxXHlVlbjDNVGbkjdJh/0zKfBkhm9L6zKVZ2
tVtWbNjm9zJsZMtM+DZjxX+LmtSxZY3eNzpF6py85pAsQqPy5cT5wRf+FJlv
jGp7mU1pdQtzRkEs7knBCIaMAxI3/wdIOGehVBL+Jzl0RPLmGEdevb6Asd7i
lXba83E1X1TU+E6aGzEPVDSWIsQILYxq5CK/o5YxvIIK97tCW4EMeSDEnlaI
O7S/OKN3nUuwZvLH33CQkWYD5AtnMuh4t4T4V9i/TVQBQsU4LmLTED8mSzdI
JW8+ZNow6LB/NsMEGa6My57Xfabek5ZzN0rBl/OzxdO8Ra9Z+IfSWwxWjCAV
jYFpAiZQj+XF4vLx0M1WYiBqj8KWJ+N6dm85Qlkeazs3XASTzzgrBS7UEQEE
Tm8kCGkW7Z5GrUXYJC9y0AUmCYbTPfnY42vwCOKIa8FiqJoZwb0biW7A9X9X
/Ec8cDQwVPQ1PshjwcOLZROatAS8aBJ++O1+DJVSm6SMzklHyM6aPevUiwzC
+YxhF323Z6kHlfl0M9WLPrXCF+u3D7vopAhQuWLeGk89AeHoxoLKywFswe45
QFbRp7jaKJe/1vpigbRetXJ882MS56tB8A2d6e3XImCzhH5B0aT+7P4nOike
Q3fsqZsStvrZo+8LvEYdB5mYGE2qh72h1bC0817DoNEW0uNOSWXRB9tHPCMl
ykLv3rq1OLvQewztuyejVcwNPQsGmHfSVJueXW/rMqJPb1Ut8kARnvd/v2Go
SGIz4l1BbD2IS0619jW+47bXVIL1cJpkTpRgQ+ItHPOKr4Z+/dpdKiwajHO+
Dikngst1wEoydcFJnhpYJmfV/ODjxjKFiBBdH5VH0DfhiSRKABJxMEvPijHy
MMGffbGRHlWdTNuO0ZA2/4wjJQALgMi0o6ViKMfs5EMazaoQvRB0MOCFkGy2
UNWqPupxi4Cx43aK7hYMeee1/x7oD+xyAgDWy3aa7qkLtI64fr9b4p5Lzgjq
ynrO6qSraGcFQA9nB2jZ7/VunADl+nU9God6nLmzRjlQOdeC0/hC88PkNY85
Ei43dbQHBsbJMfCi4qq7Of+LTpdUw0UMxqGTe/gqTI4PQLm8Cy47ixAaTDRY
0cSdwLGm46QLKXEsm6kcMRoVF1qI2dKzc1PPqoJejG67oukKSkSJ+G9O41fP
PIo4qvMzJVFSVyo18s3zcdpk9J2aUmG6aZfRebl5yvJvrCpeUy1BgUazehqw
vQ1ZZApRupihz7p8OymwETtvl3FpVil20HkhU6XkI53HLktTxOQ6rBHMLXnV
t0FIk6owoiTZqtKzDggYraB8EAOPRozmpdCOHRZNDZjeyEvlaRgaTWhiA3vO
FQ4bCWPM6VtPx2PyeYyn7dEYLtWTpEmb/nQxQGb0GtjcP/+3AGuQTgi7c0j7
knON9YC0WaQ2quepaK9kMqhye5+s0IKfslKwoVImP3rZeQryD9kBJrMhV1hQ
Ff7FlKrEwkQ6QgG7xl/NGF7UVV35ju2IgX8ttRYw/sVYJeKdO67TANYyTlp9
02rNW0i/ixFr4oldE5OzvHW/lrJ38romI17V1iK5rrP1Asd7vBtTyGkd+oqc
KHIbsS8Ju61zF3iTFY4mH6ubRybeUK4a23yip5nd98z4i0bthHsPRQ2vzEJG
Jp5JNk34vXFxq6/Q7IgvT2Eslw9g4moIUUP7M41a7/9TxjJ6EiyG531l++cr
/wKYV81wDJwN9Hsky9fBZ3oRTwJGFFEOEwt4x/CgwR4giI8/YwaKN3+BwsY6
XHvHqDJHg4lSMmQJDezHnKKvjuUC8ZA07FzobEWlun0BbwWpJW7ctzaP0BrC
HDZD1EuzIN2ecXmajeTjyQi1HCTovHza9ufVpqDUFkUynOAP+kw9wHaSwP2J
1NuugOH24pPXVceU9ubcWPXybFuEMywvy2lo2UyNxvqv9VBpKJBU3DhhNkXF
f9VPInKd7HxeIc7y6QWeFA542jbTGCIIY3Ui9ElP5kJJpPJlmFWBgS1PjPUF
vcDeeEHq3acFLQZuCyqNiLscN33e/620t+/7i2Ti9j9Bezhs1DLQLjkP8wPg
Pa5q7mDjd5W+kKMNsH72/ASDdXK3KtIJ23Qq7fhvGPiKxgh5VZIq3k/VL4jf
EWjjw8W/rw26DYvShkY5NFK2KNZurcitW0AmPgaz1yzWEntmI7/9rb5wWEm4
vpTupsshP/Q7KtigUvfRd5SuAGlhQNKF9IbBcl1t8qCirJYjMvDDBzGOWoKI
U8cFig5cZIhDWg8aQTqWa2opqaSJL0z6oSItWtrlqhosfokfXCD3NzUMzjMs
mPavbizbx+YnGastAMMIHhSRGHlGJv9GUgzxLOBVo6larBwNmTdNHR64jM1a
IO1JKvvg7REAw2mvVGuBM1GfkB81wrTInOCZr71f0Nvs7f+Glpj4LjiQKVjU
j617bDBusC/4KBojgQ5TUXf9oW0m2pK+80jPQPTgepJK2kPSP4INMTvF5Af3
iOhhlVpUOy1ZFFX1nQdC02U3/hYsKBbDqgTmyTNQgKxtC7UplPAQLBaMN/Hx
Ncub7tUCwFXnRd3KntcQs3KNiW8PUk5PO9dO0mDFX2YaLnh90HWSTYCDvrTv
sOoTjINLkKCDuMIqQpEsRg2kcaHzddZeCOTOujkV2l/Dwt370Nr4HEsd3n/l
lvCDU2RajcKSsluXwh3CJfqGHTB8U+gzP7yr8W8/wjc404vFnUFDj1GmRSVs
GO7jlF169K5sz8pyGf69lH4jXKLfm6K4Hf69iXSJflsiXz266wJhj4orxlPn
tUXnj1oyXLMHV3LzAW9m744dQx9tF+FPJ9xfdOfhltx4euMsEGHuw2cG2yGH
9xwRE3+ulk2G8drVF3TysDYL+eNQCbOxtwsGaZ3keFGiE8HaE8YNtUgHAqKu
dp5qcbA4Jd6LwzvdoFDWIg2BXpVDj+IDFfSx4DddFPt9HUMBj9Cj77o8sUwj
fyLGcebZAt3ZPdSa9Yz41E2/5vGY3tZbGSilD1xxk7Ct8V7ktVGrJuHzjJ6y
Ypq1yj49gpEdRIbFhae4mNMpku5K6lIKvVs6Zw0vHwT/eWsJGc4mb9Hn1X1d
dDOtRw7+a6m6g4vMeYu86SjS1d9PgsJr1BJUS8cKQ2dE900yiI0n444CKzu8
azGa0y3tb+/u1uarPJJZ0SSMwEWca7AsD4ebFTm21hizOq3Nkl+1WiztPaK8
oSt4yn8uj+4/AD/Nwcqhj3njDfaiy/lA+2LDHPQkTeOo/uLH9QTGYgRFt5Fa
GMmUylReLXNC3BUlFi4dhHjzVmibD4areuUrdtSvg9rI9jioMQn2tSG/GzT+
J3R9MWaiG4o8gLClJWR1KKe/uKDoDaYR7NplNsLnibMsiEMqGayhxq1LAW1X
sW/6uSb9q7E120aO3nwXl+0AgW8Pk1p0dUQodWVhSv8ygvGytZwz3dw5Men3
zfmvO4Swzy+s6Zv9XbTJPZ1O5mYoHEbtt5eInPrCoQUeGR2RYRSe9wgQQW/N
9cFFzSHOfbapUeGvsMJuUGc0zw1Lqeu5CtjK86k4VCWrVIZ2CuAjocTJki/X
M5STufoWskNNcWHf6x3S/2pL2N36VLiCGAN5246+/yeqjMh5X+ZddOh4S6Mf
XvAAj3a3n01ANlfwpgp9W8PG2ce3wH8V9HExvFhSMGOGYgbrqZ+06T1xriK4
uekUrDT2E8YwsTTGsNyAkaYWd/cL9VpeRybBlryve7DiBusXgJVEotIjBaB8
L261dn5ccIDVjPtf9jJZPS6zb/EYoBxblFJ9XT4nFiIPPigulMbIDu4JiDNr
3k2fykftaDYcPrJq2WakYFrZuW5PX+1pdtbOSj6ajqOw8CbycpPJB0TqRLZO
sAR/DOua6DpbqbPM6nD6W3aVNGKZ2fHNHWFzwAYhrGNkCsvnH0/bf0jNBsXy
LfO4WoBucgVczuYzzi+v4RQIqUJKI2z8JnPlH/JPqUdDMJVf2TqaSGcBOEOm
2bAqmwmzwHY8xtRapqKTDaXyxMF5d8U60YF3ZA6067oz1Jm6DqmyMJrw4wyN
JVEVuV8rLftl2dSPiQIPic+NmMIshhaY4gwz1QD0CnGIy5DB19TMnqTdnkMl
aVfxHFk2cRi+6Dhg37FnkgWgXPQWVKuYjwxsEatT9d9/xRq+PvHJdmCt/PEm
C/sQ6zURI9V7ZrgkKn6i7rNnSjXCffLWaaWc5uHQiUgL3b1Hb6eAoMrEIqGZ
C2g0jVqhrn0KTe3dqnSI6l2d7L6gtdIh0ug4iO4j3T91rdaEzpicPPq+Ei16
ixrrwYPEooeL9wTPOVoCL3c3Bar9vvHqrhjm6eO84gsRMNp6JLDlJlog4nh6
8yu0ZQjZUYa1SCdu7nyeK88PWJZe6kUz8Du3MEttDrFDbTpkmuRTg5eta/b/
SpFpQHZGpu5VPxxn9ZbmOzMY4QM3EqqqHtvLGl4A/0rsqgy7+7X/r3Swow0A
RlktPe0clFH/OsImWpypg30qV+slmmdwJMhwEdiDKxHpvvnqhd2uOkeeqO//
p4ltFKgH82X5gVfOq04jIMZYzNr1sMPL1bid/qAE0e7dlG0dWZi0CFhKqZ5B
YDPNIQIMd6vm4+zC8xylOp7nCgGN4KeIFdF1fymcqlaB9Lz1BXPDmQ4dhf82
iAJrcCUjgzoXZoJq23qhSOcbnCHvETAlfHg83heX3skKf/yWnWIekHSLZGo+
NJoEt3RynJ+J+Do0ITIjcuVkwuNZkGhMSJiRiCVtBFQ9bVKIKTmPYV+lZ+o2
ZMGYe0YnyIiQdspI6fTEs7dDUkUObb6h+yzGbdtzgZhrLtMsMos4yAtgzJei
WDrHrS0SQxpPniI3YBlxOkTtgkAA9ibRE9T/bg15nMoIvhSx8Kdf/4FTGtLW
qjdF9n9ZZquN5io0psUbZX4xP7u1Hfb/hedx9+8vTkzXnupkrUsBM17u2o/h
qMGsh8XFe2x1vsrrEW0nufw/SHfvnNGe65G6X1YR1q2p8Ukh/pZPXgspS9V6
nQpFtoozD/AqupmV5XTWXPNQ6Kty3Os+FYWzn77lk9UEYSUUjQk5ZpuHkFo0
ieYHanhCwD2Z+wcQNX7C8FLcd9z7Sw/2S5noyLDj4DDRESxoLcQubyYErICB
d+SCzvqtDSeV0vYARdh9sLMGSMoDsukoIRc+5ltx2ODdfNn3+KDQJxSKjS0S
PqEfslG3j0zJG8FRiF5p/Q7hrgFIL+bHIXbzZqWLb4DxJvo8rwTohDQeSc7x
kK86hUlnvIW4YzD/P+kbNFBuyyHpiFHV2K8AmDqdbOCTo8v+GqJX/5ertvcU
y2Ve1FVcPpqkqCm3287odz8pqETdT/y9mIYMn39fF5USoIa6Mpg92DWI5anG
XNRBwbuiFp99Uasux8NBwTkLNgZ42UiRV751ZjSAxNOQXM0jTQXoO7VL6i/Y
XnjXrdkaLQ8Ecqq/rhTwByuYryakWDVwyT/33jBVs1fW4kybjEiZJbvfs6g5
O2F9AxZXe44ydTR0F5ZUtv7g9kTa8Pyd7rGCjnIa4osy4zVQVq4pNigS4IlM
g5K3bd8y3t6b65/h7YNHix4rf1vaC6uUGKIxYLlkgTXyiL6MCeeM8c0vdVIk
8iPnk4Cg/0Q7aiXojNpTBq6WqMjRxdgfjIuO6XEnJMYmyDWGyLTw21LBFY5H
kWUhQy8vFZFsKeKL1HxSk4vev3PjDq/jtbCHeMG8DZUZef8Mlnkg+7b/99xf
VzSYexbNSDU3L9v/yup9A5wfDprqJ1UIx6BIV0FcSK7nO2n9kNuBWNW9xwaD
fAPel9Vw8au/hAuhD011jL2Fr7g6xMsM8dhfqqb42I/fFbukYrHa0L1OVlXk
zUpKL0BtaNBdnzVyuyhizLjAYC30wEjki9XN5rpkcvdqs2aOJmuonWBEHVZc
oNS0rus9KbThmYAbNt6e16NcWlaB4GjJdjC63HZJ3qoDOh3FTjpjLeGNC6Pk
jNXtWnD4rXMmA8e+x7rbSFWOcc3iEY9joyPPNRoJA8tPtv5+X3DsMFLy0aDP
/vVpDNaJLZskN6HOc6WWEi/l2m9eJRHTjxip5CGu1JTeFz4eeb2r+YB6pHD3
/vGZVqaDwFem0J5Yy+fZySY12UKf8RTbcUmKmjP+FtsuqsQkTobDt3WSUVaL
JeV7baQIiZn8cH7VZrzk1kq9dmJSVJtmQwn6Qz0xNJ9hO6x9NyjkxKQ8Pacc
Gg7p70sDzuH16ZHz0YeJcu6OPUlOJBo2zeslRTidv4dql0TsXjMRgK5bmhTK
ArNuGkCjsOcv2Nu3lmSTcbz4pK4pjlGMqhKdifv7PNIenOCtoIdPyvZ3CU9n
vcefgSTSTBVCk/eEI6ZOmzIF4eTOqk9hN0cteCGrAEXnIP5BotsIZ23tbWCi
DIo4ht1CHon66s857DcQr3y+D+NTxWOsq5VO9lJeDqyO5fn1SY6q+Yfrw8To
FDc1gjTClJ8WhokqhD0oiuJU9C1W7BGaZ/FU8EJEYJYfr1Jn3Drc69kAEggS
SJWRpF9MW78N2GCKhrelijOoot3lU5du/4lzTUsE2Hb1UQUi+feLD95jR1GO
sTtx5X8xoTwcSgx+u7iM83lA7biITYze5ZMWIJZnuMkX5cgRYiGhXnSSyNIC
xg6SvsqL7Uz5iDtTFpqfBc9s0v11IcWvQBAVqiPO0id41mA7HmkX57MSHRJJ
HoIzVw848bn4AYF8X+TcYRP++wuF32FPSoQRAAWIu2ncDKItHpHhvS6oNyDk
LcqACFOwGoxCphuqui1eFrTFPEQYXjjzwRrluDszmOoYJlrk0YR+11gUmaty
WUtK/Y17WlDFtKja3wNun8KJsG1Ihxw52i2KtFY3FbFeQdvfEx8lgXovW8mN
fR3U+uCHqsCfYgrYo/D11yBPQ5JSCFpTfYGwk/0Tc1hODROzVfLJYWhrxlnr
QXF27PfI6yt/P5RYE1dTdLzhWneJ84bDmsJSOKgvdiHsW2YFEJAFdxzaFWGg
F4USYaphYVb0CZ/SgbxvWl7REfS6yEXzQtwBm5zZDN7VPx/at47gWQUQu1nD
ZDNROP+7S95Q+V0Tc6Nnek1jnnyFEPzN8e4aA5tP+fYWwpXN0sHVbHDpeBa2
/oRmMyR1qS2qT2Jp3p66ynTqfJgs1AKTSasmmvbJFIsmOWwRlm0SeJ6GPjdm
1G9sm8LyJYxMC3+Y2H4IIUsGElZv4P+GeJ+5tlSnIRu4zAE8Ad+eA3hzKrRQ
RGbFRY87eF3SGsWl4MQyYrbDyj7xXt9hmnAxmnYFO0c8y0jO/pQjd99V/Z6P
X9WNup5+pqHPFOkqbjkd85YbYQoUoxUriYImad5/gXSH8Va71Qree9lZtxbq
qHY3F4gpOWrxihXc7US2GZ5QlmZX2ged85rzpG39jGelUSTjWA2fQq5qHqlv
Az6Dy22W8tHIy97ObZVf5B05vq0qJAwSE5Zl6ADboa98k40CKJ97Tb/ZB1qL
4S4Bdp9QrEB5STskiBBsEk/ogjRMuH432VdNRqSoVmBXUqVnUp/hSo1OEqCM
Fexm/CB/A6F7ISM17H+FQFNbd6Yf1S56MCe4/XyhvQkZHO9cB85+1Vgjzzql
qDwQVWKPSknRDZFyQk6vu2LnBVgMKEpE6lx2M5jem1LUFOxTw+/eLri3Z2BK
TD4+7PaYLRib1QYV2W4INgdAa7nuT1KMzJf3jhzCKt74e7UuDFKK7eCf9d/T
kWj/tY/1RSJ2tl4ss8Ix7jGwZzhorLBjjLrB+QU+t/cj3T+P2/whVrR8dsV2
EjQzPRa+lUEqk49xVDqA9JTLRR2Otp0Oklqk9zsiD+GLxBkzqNa4pvbHuA0l
zm+Ec7KL5tNkICiETOsgN6tvSpwHCd12w1uIAab4yUYaGzuikUEmtsodrfOI
j9B5BtC27yCSFqqr/CYe9WWfwLq7cAPuS0UVo8q0XXEXWxO1r42EkzJA/hQH
RTvtwehVAdA3l7NDB7WLcWPp48FA3Ws5ob+wBYCYlCvbCjNsBf9ywr+7+mJf
OBDVINqx03WQrXo0/fX/ljlbHLJiiv/CfxjMK34yJcz7S3DAdNWbeyp686xF
ym+LY/eU5d1f6zqjYlhwYRF49yLOsQ3H0K8IZ8jLPzXj6JGH9RPbreWGeN8a
opV8v3oNjaeawxKWCgpje+vyGLrdSPKbjP3A4AFFEq1YjpkTPnfFsQVYKADf
5J0xx5tPvQx7et6hJi3qnf79gk8ToWEWYucytLihaBzhXyn5lb07fYkTmtSq
sJTYnIoWBH0h9+bWg8u2r2tMjlcUOv08XqEfwL27jINUihfZ7idvrYesmQIG
UgkufaNTwCZFcDpR9ZgD8Vuxz+fKaGPO7QgXreSTL84ydt5Q60ego8/R6Ip3
DBdRm3iij2V/3tRPJAwrDhugIQFZpcFhKpPN+MACG6iFjaCl7N6Ouh/SG+52
SZt9nb8278MXQ8nXbnLwrHOVAHCNmu1DqkutP1rvMyV9OTP3GUw0IIfOAkRJ
3meXJLQYo3YHyMtGyNhFdNnxS2VcCxK3RUec1NPDVDMrtTmeD//qwMSvWpHD
fYsuIiP18TXZNiD3wrsli+znzwv5F5a42O7IWv20pxkTxYkD6bf4AV1ZVgk8
k9OEPWUX/lYb6SMFobnwK9pfexk8og2PD5ZoIjxcOsCRgI4E5aExYnsi3uQD
oy7Qzz9QFoIgIu+Rw2uZ+xtUQChjF4OT2zrOlEG9oiV9i0Kh+aJX6nFFhauS
XNuayMdN4Smlv4+dpUJOevww+L+aYYoMYRC0WmP5n/mVyGomP4rlymDFQ5B8
E8mvTtBUxmhHGOcI1vYVnbtL7xmzefMn1LR9E4fxh6lVtCu0ggkIZ4yjkVsV
pKb4EAPBnwKn5Wxu8dmeVfJ+W7U/EpgLGlHX8NsyZRQt4PTW/5YtAvA1uOsX
3QZODcUHdzPXxu2zTt/QCUyQJlpiYUTDeEYhJ89SAnkKAaZoOUFyF0fgO23/
kWOVJC70keFB7I93F5nSkr2waXbtCu5X3m8nNP2QRVbjqeQEEst05GlTXv2k
EvpsUZR8qmp6wQHy6qjyTJWU9sHBRbZbGNJm+s4LZ20v1JuE6n1yxsldYadZ
fxPaWp1Jb/WjNBZBiLpDjE2XnRkdfBxbynzL5JchOr5sumBRdw5q46c7dz0Z
hCeDrI9TGPuhITkSmUlx28EgHS0HEMLG8FzGm6v9PLFiDrFE0qBsFSprfGJD
gLJptoHhym9tne8K9UmO1irceWKaZFSSajg5p6gsl3rghkjG7+mDjXV5QrAa
6hC7yRonMz72+lENNd9LPx/S3ik51E1/vD9VedtuqA/70X3lpyW+P6OAnzo8
TALDcRpwmXHZR0La83UjHWFQw8/1JaaLaexHZboI8dhv5bi76+RiWfA7S95k
PcbaCJxcFqxnUBdvmNXrXrDDYDdgZY6UDcnbfR6hJBcYCMyg2o8pj2+zL9Fv
Ru1xtib/7QiswDcpBbTkwekpKniIpkK9jptmwWGz57wusZxHADUHIs/oio29
DdcnnD4qDEEU/5ng/M25JQxN7WeoQZXya/+jIQP1xDm/lhaXea8Xn+bq5WP0
tGDiUwB5fuRlH5IVF5nDISKbGQi95G+/fGb57MeKppgH0qkko4zMktW9guRj
p7zeQUCJiXmvTpYgsnAWqrS3kgbn1m657ktLQORDKtc77G5QmMYY7EZIqqI2
WvJNXKymxmPrENtcJhr7XsT3z2NAIUNhohAM8mTJtRS/lrn9n1JBJRlJyl8x
euEXQcH2H2ZezqyXHMtyi0Rz8jzV21khcZSdDveque7urzBQHzO5HmKrY5cN
LOsjNYnTrJLYi1dYVFMZvLoN3+J5fEFpEdQBnOtPqw/e/FiLd5AbOZuzdcct
Jn6O6RjJB+wO51G1t6JyhyHRKdaoxHmnAcZ70KgLdb9ZVJdHd1Ko+FgEJCGb
nat9ZeqbaoXdmiVQK48QuWps8NI0MB/7nWcZZNxOqm/Iz0PnMXnjk+vOaBy0
oKy/1nG69e0fjpGYEOMomvAdX+AcxUD25zfxKSQRg814znYI9n8i2divsaiB
ZIRwYByDcZl1C61IyZ7VCCY00wzUK2gYgO+hDn/2N+lwQuCX6UoSLphgqccF
6kfMaUYg1bgvJFWWmBYaG+SHA6TEzjgxXBzUOcLLaGJVOP5BVcj0adz2SxGF
KSGcHSixdEdlu1jiZHRHYLOkapW6oX6Cc5kQcOKAjqrFn3G7FzvYFUyoRojh
7SXUZh68YgDQTXPASeKUe0BK++Nr9fLeVStqDvv1cuPsgDAIPv7jUKs1IWnD
6uczeBhEoxK1ZmAUpGaMLFjETZ2mAl3iuBd8y/otHe+QcEP2gOvrAig/AXb3
HydmAoHWsLRYigLgpOs2CVMjurR2AnpcID5d42784OAs8p9JmXIPmAqGh0F1
8Lag8YPUT7EzTszT/BO5cGy4b0IFUctQDKGoNKWtTH3AV9cYwCmONS+FA40J
EdyWvpg/DadISGB0oEKx8AmUUm4MOFmgr+jc13tb99fOUfvRlNasq/hQun9Y
5PKwOaeBEJzZrkReXhG+AvYDKt94pVjw3KPwvu/ivXDzkIpr6vZo4Ip9pAq2
ExdYzOyREmz5G5ddlyOClnxNuXiOt6iIAsyovGubXFmxNJnXjRiwZI/WO33U
3KbSlDWLqxhjXJjy1eYj6NjCljhPATbBx9IM+pJARnDd1/Nm4l67yRgtsX+w
wcyaQ9pdR48AQzpHyz5tOv5FIhl4e6cmBvU6SCHT6GXiCFfmpxi7krkqt2p+
Q4avZiRRnLkiRbj7siLSWQ8bg2LPhpz2XFr7dMNL9lVSCfItWxkUb8SS8Sx8
i+Kg0KRqDKhA/hhEKj9lO7G3/XLA+fZWkQyJ67orjxMflTFE2/jH+zHPk5/J
G4JftQikcc5dFI+5UZXGLI8nsbtoqs9xB8HwvXQ5168h3QUwtg8TjLU7isyK
O87u1EbHTEZxy0XZ/zvr98R0t4OEXb1Xu08h7yduOjfCH/evSFpdgHD57fEJ
A8ijb5lpeEe8sFtrZgxSOWRMvCkOkhzCH4v0b5whPydLIqVaiUaHiTJp9uOB
bgSKZgaLH6nZiqvFwnYoMAcukG4NovehPrbS1TlSlnBIjYVCx9AWa8ke9VkX
nQAIAFNJ6czvzo/L3aSpnLeg/62FKNQ8pmbv+uEMqsIxYrWmjbrdfS3YkVAu
B05GJyjYtj0Hinz6ZO++9FQU9SYNAP8X//3zdk8kJW0/GMseyQuuFYWl/46a
KaXFKIsOTDvMkm0j3kl7RR0Mfp1MYQoCnhhFEK/vj9AfVtZCSnZCNyx776O8
wHaalvWko5aB6AuTidF3JSYXoGxDC+vj5iW+Jq4kURs+hskg8XcLL4N5bzry
NhowOaBo/UcK/TgY8Bw/qwDACtxeVe0M5uH/hHoRS+/QlBsi+L2joVWmekvA
TvsOmopahuqsojm/plwCe5cYt9HC2D3aQEGUWTh3ll/KOUv09yq8rcWKQddB
ubkPhtFFdvQwXL8LzB1BbU0EbRLJ5hjUWvlAqIWx9sglP4FZBFW3AnRedDow
XucJ1weM7AZrvK1sL8PQftLiUIsQmU7JpypbDhydyldbzEu0fAhFA7jsQmWT
bhXOc4VjRIwH/qRJvG4ia9qfxneAVzZn0lrPURFca0mT5UKGJwDlc9ki9kd4
Rz+SODQeZD8uYKYk7NaSQaeG8ayw4kE+z9jgy41GqCwTGMZ2FnZUBHh1j3Dj
m+EbWk637vESC6I+FVp2MEbwVQWVdkOLNMAyv8PtovHSQY+hwqgoaKMTNEfE
AtU5ob7AN6EAKjPRwAdMd8/CA4LPPfBaX4kewkEQ6/kLGWMnTf0cN8dfhQ1W
aYNe8RJxSfbu0daXmowU+Bkukcl1cRLeBelkGJXZFT+s6IkRgx/vMPOzv8QM
Rn73CK7HUHaEv/3WvLcm/1I17DIzVW7lwqCBch9ueMOmrOoCvxrI+xlZBLlL
a9eTf39fBKE8223ozMQHFeVBqQHOik1yym1xXMqGw5teJN/eO/Tl/C7bXjN3
bP1MYHP4KH1+tCp6wy2i30qmbN2jhAp6w3040AP+D+fezIx1HDYpBt1dFgG+
U26quY0Mh41EvUSTFCsLCNXltZ0XYRd1ezgXumycrp2ywwozz+yKff4qxa9E
D0JJ61hY4szFa2h8+lmvsvJkY56gKbnyP7eBPOyakppTva3FlJeWUcL2Ha/C
VyDldUrn344zqxO+oLRAjRjJP2K1AifKFBpoZo8G2sZbt21bTKf2hwwL1Wri
d3q3JABUk7t+Xmy+g1hWoHcQ987kPfSFo8/ONow1+Ww448YUoWtoX2WY0UgY
PJECi+VQjJlnikUW6L69d3c/h6Pk+Po08JGDcGbEtnPP/rhzwaAX3Ht/m1dS
X+G043MKvRPYe8pMAudJ7trOSgHBfpl6322J9gjyesYr0EYzApstuMqYPOAs
dMNlwqWycte+gMh71yfdgfrI5mnGCzobEzjfdJuRpDVSJZgAlNliQVuYesq4
zGivjcW7sRdQg8RH3XIF01ROCr9zin/AaMenmsHqYOpPLR3frFT4K1BIhJBC
SJt0O+n+ZZU84SFtrTBVLHwuIcriSKFayXh2N0was7WfU0VupX1K5Jp7cf+t
2YkxJ9bK4g8cYtxqpp6VDu0njs2bl0W3w6jXwAgyJoKItkOguWmWV1YGZ5Mt
jT61bf+2Vs4c4zyGzzJw7BuCeVknNJYsV+Fu5XMocgfJNbCPZ3lf3QON1Tgg
xUv55lV7GWRmEga7wPzf5S2K23GVH6rd0WGlUojdOv9Qb6V2rQWSZeTAfOeD
IowTrBtaaZzlP6fiTIU0gjZf43qA6vrhU0k+geTRWCGvsha3M8aBTirMOgwe
Is0+Wh8TnkfQrCM9jPK49wHmzHnMuqeNWy6RD2Sy7kg78f4CPOW+2qKyNkec
B1dXiDhnGqhv/VtQUpQTo8o1o8jZEW7+uj3ODWbBlFscvyfBEVjIlM9bbbcR
QGqmXTd4XtpJ40AwK1HLl2zDApd196g6KFGWVUAwq23+1u2sZ6de8Ol7xhJ9
I4QBmXiF7hcp3uZdJF1e18trm4s2UWfmc8eiMm7q6O5aqAq6tK43BG8gHui2
H/CrZ3vsgCQRSvwVVonGIel53GtUmhK4epCb3/r14EbWO5eT4hOWHH6u5Lcd
3vzJhMkYM6QkcDecnLB6alDkxAMLRsE0UMbgD57V8taSiv9y5cGAyZt0S7E7
zgiu8VrIy4mtqFblSaf5fyKlr9F7a5w0MVlEKj6721FTOTOlq0t0Yt+TOh/y
L6+f/CGJr/zsSxyRf9m6XJKiHDjcfcDHbJRaOI2uDyznJKm73toO2cndsCE7
eV8L+LCLSudFnxVfd+mCoUe3OOHJlS+ZYJcmRWH6EpA9X230o+lLHsWtLkAY
7Y6wwXke1N9Jvv7d4u7iGwiZpt/P+atDlDbk6vRz/jZeqvYcetfeRidAJSbT
CUSeWCbQygukWugcc8qJOAY3Fe34RdEaUdcQaf3Wv1dtd4MNGWGNAKetHtVL
H9S32/CwNw2o+za5CkzrGuPzdzwvwP4WNMHs6cqdyzAjM/TwALqtg28oO6m+
Czfx/4KNYSh5RUzH1IdArjD1vecSCDVr0PV2wYdkp8ejeRA1OTjYSJelcgXX
EhFAsNhYzpsBk0GAV1MtdO71h0mojYsHDpHb+HB2rW9ONntoNaTw5rOmcY6+
P+SYb40FqnQF5fTCGMNpYMx67WB19hfKNops4wLS1zyorLe7H9aTxkdPvWq2
7Dxygcl3bXaOkeT29O4HKE/p9cZe1zlR/CLi20ym/HpWXh9LGsxuT6/5btPl
itnfxbrkHnneRtoXcHdvmEFSVegFZKwwQVY1EEmdL67l45w9zC7P3sl8hHa1
RCQ6grgqWJ8AzBmo+NQD+Vo10dvqSsz3vKGoVuWySP8tEBKwsytroptRI4Ha
wGARLFQzI8Ya3wdkX6wZy2i9FsseDvaVOxO5oH1I971yXkzIQqbDfzBnCHrf
S0X1/nMmJqb3Xhe5dkOtK+xUV0D731Bfk5g4fLz4FjDpuWmodW5ey0+6opmV
btcUQCwtBGiFHVm2AKaX3W89LcqSAEajsEMtMxegRsPWh/W7CxxOHloxCpoi
5qzZ11lxmRi33z8OEd0zxIR8UsW10kU07215gS7LEjUd2HDgEre54SJE1KhA
nbnYFgoJfTsNKfyLRf65I3zhV0m1OO4dUIKpLh7WLiBd+wP2tcPFIzrX0hzW
jo069I7+ttupRK/7WfEsKiIAGrc4nrzH0YARIfo+tKKHzXKR9diD5pFk3y7D
9ysT/ct68jrbUenu/VUrGc5JpXIcuDYDeUtYtZDz5wUD/90FyPD362/pRXmP
SbD9Hv0gCE4JfZ3LwZqSdPT7DqAW4fKZAiqpdNGcLgHYZijXKe8zMuawfugJ
r1LeSy8S+QOY4uvXSq+D15zTX1JPIUdZ4bktNZbFjy2mXvseNStPycmaNl5w
nlE95FamT8JSmivuxghbJVoRYBtSYX55VqzK4rfNfkLmqIrcoWdD/4wSUF6Y
/tHuL9+i84PZUbYDrPxKT3nfEM5wSvLx2oNsFASQU2H3nFqkOTIMcMMeCuLa
7b0ME2rYpRRPl5vpcK1jAbipYSUo3/D8Jlhi/M9x/x+misGGnseQ00KiC6MZ
MKk0jOqArdXySJpkaYkhhhipgTm6tXTS7qEZY50gUAQHLvUPkroMjx16+Utq
tFio8EBKkLzm+4G+Pu29RBv+DvrR8timUZbb6mFE6TzCU0G4fe5bagiPBbt8
v9BL+ADHSn+XgVp/oNO98lYl2Lkbr0gBplmVhrR+icw3vBSrHuM32Wo5eIb7
rlnYiYDvo3ypuaOHt+u42foWKtB5BAdlMBozfP75/TQcO5FIo5fj0LGC4NL/
RG39mZJfr4aDBbRa64A4jae3YOK8iqcEzSJWGZmQyeJ2RpgzpI1rPn11XCaL
ZTKScV3c50qdj+EYD1BlV1SOB2V5NKtISVMrF+k7gXe+Z0eZ9ziS/5zvXqHJ
ZcUylobROT6gObiy/f2DOIa7IRV664HRNE715wi8WyxjS3/0YLpNTIYqgT4c
fW71BuFNQ7aQefVAY/CnGgBon7oaEqYP6cWSa6M9aReDm4NI5Csn9B/buG9C
OGLsjvZvgzq+R4uTfU5RGxMZvIMLiv22qMPiwRv73J4T+Ts3XPDYXgNvL79p
U1uc0Maj6HfYfeGAb5w5dazBlb39BCx5HkUQ23zJy+K1VG99W7gtPcnnVZuA
dt/Ols4bIX/ePGfGq6TFIxX5pEUKamLRDrQ8lyWrG2tjdge3/FhV7G+uR8Qg
ak/7RUCEdlijRdt1nwu7XVmvuPmbv01q8L/tn4nLy4/Becig9pJu2lG9BmQn
h3cdKYvRZWtE4xMBS+ZOG7px2C0QXGH7pV+Vd+8LAonTBq8IPItZa2U5GiND
izt40QjoVKzlodDTEf2Q3Ux29aAg7sve8PiqNF3cH0DTZBpaAULnyJT6g+HD
nHnbNvnlShHej/uMlVmXZ+tuOGTCsodHWintuUw7MQmCUSIqcbCcCxZkz88H
xXwRLYZ+T/ZzGW6ipGrPrVbIBOr9EygtZ5rFGsv+s+7es8vjzEOvx3vIBdKk
N5XL5hTep/q3xXWStG8yVBe3fo5ICmTja/CHvQk3XvEAUfujypF4gmMLO1qx
lE2W2pCyYpfjezVofevcEUGwc5Lqg47tmDhmIMInrCSoMROD89aNyCtQWs+H
D0OZnXror6+fEX+hbp2lfD5adcrBnoccZNOYObqC/1oHCe/iZes00Gr+iJ7E
dvPWmVvf+PPYREfpYYroBpGr9+of59US4Yehv2f6teTO6pbIeCfoKN9VFRe4
Ts4QIcQDau6kScO9ufFnNuwQ2EuELBeVDOnPfGWWzLD0n6DVUXtA88vkzrUl
5oXuALpV+YyatZC9mMBox0lugSKK/HzA5Ug64HL9z1z2Km42Po9uj2IR9bGQ
vvd+Y8t2Wo9v/p5mPMouapiVV1pzfR3WYOOu0B1Czwpfzk18uoBI38eHmL5k
lrMj/VYhnbLXkeyUIjDhsIneUI+t8EC+fDjoM3t9xBxRX6urjBMuSSqMsvjV
p4l/iZfEAANBlj/A82tfgjK/CObgN8GFkmLFHbIE96oNzx8r006OjBHD11X3
xED0lRMh9bDcpOTI5pussAIxB990+lDp4rV01y+j8hdtMrXQPWuyIEa779WC
/2sPdGKxTeiOIFKH5dlgvzA+G6fvSYGW8PRUyMKPpqNiQXWuWVyN2Ksq5oCi
kdSRy8j1azhB+2eHdjWMQhI9u6leCMridWPkQBuNp+6Etidvh1O7FG5IDPNB
YwVx22MOjew7dqnAQs6sVwhrsm9VVI2w1nj9Nerag56lOPRIsTQ6C9jR6/bh
Yc2AIRXgisRHxHXY0uzNYnFdFEEPHnRIHqiAAjpAEjNpWDpyrZ6psE+E7Ube
iFPsDL2HkjlMv+fewb/AGu41G0iePK1/tKcQOV5wjun2/azAxO74F8OcIVSc
VL3foL+xxpJ0udY6zraG3JGU9ofHfeZaZm3Noq7pCi8rdZiPjb7Q0syEQqD7
QC/gZfuklwH+0iV01ooQjqZ2mRviQ85atwGo1bHegkafTYv4cIqFjHSjg7G/
7Ype30Ey1/vUDlHP0ILSBK+4LrDrLP1G/B/phbZ1eCvWmaaqJh5H2z4hrsu/
Py3NtVnAypUKGnqjpR9QZpKakcItkx76ZywUpTjuGDcgpkz9i9URloDYb0tE
7KnOPqE/Wt/TYsTyGTNvdwWSVSI8S+IFWuxU/knDCZwFdSij18CJLOBNybvt
Ni2gJnK8zgojmNhJRgzi1vWhb9VqPu3qrJ+5/iL6YOrG1Si0ZbosGFjFykaJ
gHFTHLI5a7MN2vs4ah/p/5pVpcdCVzbernGR1fEuBOd4g3krnKGVtKHWfWoq
eMY4vBpM0f+3304K2vSlAyuEXQk1vVveouxbG8Lqi2wpoPf8hefvD60MTFc1
lqgbGikco8kzspThzIs+XZS5ALdLX9mdF1XuxT4Srpsui8dfY7o0qxWWyBP8
wYjGdOhwvDmdgLYrMqDyGvTlIZAVs+Zxp1spY65qerhF0QPqbW2YflLwbDsI
UmX9/nht9rCU9mf7snaX79p4MgvSaS3Rp712ypK2dVq51KfIwUfVN74XcF3/
+y5bF4UpNmPAoYCFR50k/SWfAgdREfk9MzDKLFnA66RYYpbjVH1GHDtFcZ3H
Zn6ba0LIZfnhjfNvwslNpleO7PEu4VVpSI479LEDshb98k/A6a/ghkrodx7T
BQTauonxcYw5PtOWTJdXgEilUX0Il7+U0vq+L9QWIbZvcnrVe05WYO1l1fm4
n8n/SM+oZ36m3n7/IeNJseEOi1pXe1tmSuTYD58TN1EtWCuxwHI5KbFM5szu
+SRku9TNdFbHMdUmqg3i8cYboBCUda/uZdsV/w2NdJcK3rqJ1kOSXHkRwVZb
WEvTe0cdGFU+QH1bZIHe0sV8UT4CfVGj08O8vBNNlPEhE8VlBk2YoTny+7JW
kSaRHgiKY4RFoWJvqZfRnU4Hsv2Y6ef16HPoqda1yjcNp1voZ4aKB+YxFVIv
U8HsRbif5MSkhz2AoiBky2lFL1R4aFLHHvupWMeZj/LTnfW88EPxs8jdoRX8
TY2DlKPM++cwMkF66kw5XMmAQzyJYgcqocF5G5qyYBKSp7X+Z/uZWTDaV4a2
36VI/cPv71ulQcI4yk85YNl0DX9ZhFJNFp0YsAlofi5bjU3uM7LKKOm/Bfif
nfJ4laJki0Jf69SmSPxcyYI4hNxGnZNv0iiIbNozdagoqph9I1GYTXP68ob5
QS1wK/xi9ox9BLe818MtCD2yGNYObXSHKXeD4inF5dKyRyokb0y5nqGWH1hn
MfKpcF7COr38X7f9Vgr3Km0VSvYCHJJBE2fJs+9a6ADnaJWww6IZt3e6e8L8
A5n6+ZBS+re6zqPkbFPmuNyPGZrLxXhMCbjZtDqdwZBFV2TflrH66e6lS2IZ
5N2o5WqxUy11MvUoaHuZE/kN+ZzIxLD4dEXKetS7/ARMTqzwOuX66GpXKBKT
4ZDv5/3PRDE5csoLN1SYSa3jhZj03gQlZYTrYmmUsQGdIg8XJtRIIhZElvCw
tVaCrfkefcro9cgzuzX7RvmoY8si1Tx7qaelijGqZLRI8B3fA4RIuRd46NUf
kDn2Vsi3buKv6oaN8XJmQpBrAdzyVX6enioHcUvpu5nBAz8Apf2WXFJJMLRX
ZGZ4uglq0RVcH/ksrKJLyBsEJejdfUrHEEwthe6MUMO6/TNp1iRPli3zkM1K
M0OVrsfgubWfvRsaWb9W4MOPumDa6bpqQ0ZJQ5DI2wDUAoQeFUprV7NrfIVt
fh8VLf6YO4T0qihKjfgUTCNWDjo+lo8YyS3e400GXA8NNQzk4DbOO5c7jQFI
JgLBrd4z/IgJ/5vamGUbYnQPTUgKgiHUZl9FTyOniPgH48G1J9qo3mmryZqP
+mMENwDtuayMHdB5l2Q2DOA5HvOUL9FUgSuI7g+nqDVFiloiewnaHJchgqrB
wzrFVJT7u93dNGCpYwv/uBpyynrrdMQu0zRQX0k3Yru1V2ANf9IPjAcMnegl
QZImFcHRQJPTPKImrOv1ctJG77pIUPDgU92Yvf4RecwgWYtOa16DXMj7P0Sr
8+u9J/b2s46f3U9QI8VCqULsHDcKRBDMK3h3jc54P3Zin6G6P/ht/JvYWhQE
63DbMLBhFC7LhMSNh4yOHAIvoohFOCzBN08ohaJ9LvykPVQHkZdpwbQXxhb9
JPYzAfdw0jVcp2H21aSSbCMb6rHuMOUgX3Fo+1ZjRlIzFSyC11h6dLfofSPU
XIfm0Vtk/3Lorp8cuzMvImiYlIX14aQcICe6iZE/9Kifami3tvCwl4dssvFU
BDm+HGamVUVAZ1aX4CBJdHbtOD+aBhUvAj3daBuORzorNzGi9VLQQtbwqJoO
n37xPDWUe0xoqC/yW4KaC4MeB2nX+RbKokM8s4t3Gsbhl6zXv8Ox7qpe7YQh
ga59oYd3YmfZvZc1GGQx+8IzXyGmctwQIrBiakvHJ2OEPbY2tRf0QGKqbNeh
a0IdBDBbsu/gvL4f7cLawsRVHorLlio/HOVwfJj2nr2V/wXDymh5LlKi4kaJ
8Y/9LVDox+P4G1oCk+mm0YrTVkfHdXQA83BFCvYozfIXAu5kdy2Zt+wKScid
2EexYaTvXnYkEJHkKY2L5m0/2hNk1n7IQPFjpbTe/PKkFJkPR1ZobG4UAE83
wyDArULVCg7P6SfeqIIhRF67RlOQZMiFd4jTzHMGwqYhk3+oBc6fd3JmE+eI
wb/2JsOlYjw4ZcjAYGZ4aINKsDEzz/GRvM7ptrQ3c0+H0uKHza3dOb66YLzU
HrlB+H/pozXIrv96lupJALWmNtUap8otw5EQ+hBKpF3uCS2XanZ0LLRBEfBt
vTJYk6J8/bt2zoQ0MeRUjaVeZbZOebFz72cBqrc09tZGpeyOFy7ExAefa4fe
6XeZu7EaxC3rot/tMla1F7Yhzs3JbQaBubwDhBuza1Ix/C4xvUTqJSKWMdm6
OX1HPk/5JCEIPE5GI5K5r51xakZPdQcdOufd1usARB233Xzd0XyJJZAofJ7k
tBHg24ixF98Wl6LGnLbra4xhk+5q9F3kctYeGcW8GGZhF0B473qIKa5syvav
+dZlQVF2VQUASXn0aY4u8kQFfn4q/6zaMJBUaFChgwQARWsOxjhgASIYIAhv
WtSlzdKfPsEthXBsv6cXVWHeQUabNq5IfDUIPE2VAeNRNABmnZrUsIqudfOV
o3aVhEGMMx9wfn4IJUsW0ecKRt/NinnbKCV1EVJrHSSvR/7gHBRV62fQBeZ7
hsx6leglxuqy5+QsakNaLC9VgyI4AzurmY76d7X8Gs0VuzIrldDtM9zd3fwy
uPaDdAFNAyaCqntke5Au2v+b0vHddS7ok6RA4m3QDECCCYsx5UfaYu7jPiy6
6xgdWGtGbhD2r9fR3fvpChoUB2YCqthTb6EFHI6/+6lE45L1K9Oy8gegfv1X
euOkNvEiKmtqEGwFS9NcuGi2prh/qci/qxckQ4lAa/bg0UjVNOYNaX4Qpp3p
iWzAZg2UTHHzzw9a3TavTegge3i+QmX68pb3NIS92WkXFwoxQOavhC7tres4
yf1sodPhzROC/yGINoKLIAz1wOQmy/Sl1DLsIjthQm6SoqciD0IonkDuF5Xn
HL5urmsy6UjdAoLj1VJFYPIBtT4zC6E3Z9amLeR7UqjKfaluvzVr3UpmOgQv
18TZmpBfhGF9LCh6V+gwTKYLzxewFglJrNnVWH1En5qv5kNCDw7V33qPvg56
JC8fRLc6TasPzn2kMcVtdEbZp5qbebGCB9gjDmPlerEnt64uxE+5CSDmY5A4
/Ks4GQE4JIUI2zPoS4/BzVy38I9BJ8DRSRj3kSWC2dm4tik7OIdq1FSBVpVY
iauuvo/aRD0dUWrEV/FzHvvJpVIZbzM/Serrg0Rrr0+Mk/jrjRpNXnKm+XZY
VQwmrHOvaljCKMVbAiEhP90IxtO0RlgONJb3r+yyI5Wnxxcv4fOFX9HPkd7L
j9UlNtfuUUdAtMGPZRFQFqmez1gyaTrL2YOyLHbx9hWXA12swr6PvVXyKmVE
tLOT3GrTKgge0hjyhbGw6ymUdOgDVV7M+knxqRbzqSZS3duv2FunxgjKYu4c
P8c8pkz1aFaZK0NSOuFhZdj/Hi8aCwow3cejVgf5T7Vc5go6EebJirbrNyG3
iugWUxMTiCKK3v8wZOIQtiqqw4/VLt+k+eGN+uNxDbaRDolcDcFjQqTjCrn1
0TfmE1rcYGpoXilNXxMzBt5nvWM/ZSle/PPCrBVj2IuODZfRmD+Aym+x2RBk
F4k/fCICxJ+YiW0LgT7WmH1Gpp+BhzasCl16B1Fydu6M3wrtFxuq4UeIMwo9
QpexXVW4vK/kg1NAYZgURkoWoIGjA2ihRqMqBmhoaNVrzXZJmqXt4ViYgS9D
9oHLAvgsRftpJA/kPS8mneXeVvly/97Kxyfc5JER9dNv3gm6V2PKNRaidpXd
rvrtI4TQ5Nj5lB4MLT/1QCXUfr0YB6/vsVCwbW1YT1o9dW2UOzN7n3avMSVH
+w6k3oJq66J75cbbdLpxhjBZLm85aMuALNdNnzx+pKyo7jQgi9LQXXjJVrcg
4h3ekPTIog/FZe3Nw8ScBGE1SaoPF8vBX5PDfJefu8RIOYQWvRGY2nJ4oz9F
dRRBFk55UktQTF95fThckPQCtPgqwl7gFxyf7Km1pZDnSyoAJOWpXfemgSPJ
jKRvIJCWXjYJebn8HlnYsTMsKocn3fyZn3FnN47H3b9oRWiTexCHPN0IZJtH
1yJnDRSf3b9A8DoxWrQlVJLPRyKJEREeY8iL/q3Hxo/vArx9lVE+Rv6iJzb+
Xi3935jM81qJTCXjdis7vsKeg/KIa1IpsDvWpyn4ZDpizQa0vmGkZnCRbYGt
PNDnhwcEE+H0w4bOL1YF0WagEauWQslz5fr8h/TlS2jmx7+HuookwP1seKJY
E/Vca9whY5qaVbMcEGwwCqK+oX9/kuQ7q/pmdcXdeJ9H2A+XjYI3/YJk2gF3
vGE3H5WhSBcwMsoAQ3b9ZksrJutoCnMbp6DtxEAfTtev0l5SPHoEWTZVg/yg
jPNkIX2pUZ1yF7PVvs2XzM27Dq+nOzdkv/uLuiPjSAKznUytC8z+zVxoJLif
9Mm+BRWGzgCk98XJd/x5tJDeoVkyiMfx1awsNIt9c9a/shLo20NBDWjIP21s
YhzZWaQbSZGqdCG9WoNW+RXdAPbdT0c30oQY624cg9dZs6/LW8Q+LicFt1wu
uNgTTjTeXTBp8aTYbXVh5G2gdWtAh3mKuvAiYOgbH5qP2OPrlpVidfM4wSqO
y7u8kDV5hSmQ1C7KuPM0Om7L0r9cxPAFlaeXvNXM8yLAxDL01MJx4xaBOfbR
5fy9mD+ja6zLnFNKvOUszTXAuLy/eemLKkLQp+mOzuMQEG1iDLZPhRFHxejq
Fd9Ok5yBkbKNdKy+7aLEtMYwEVx284Vr0zCoi0lcr/MfWQsrjOPSL+FRvefM
pfVTPxSWd85itdR/apHyiijRKF/N9+wKAzo6BTYRY3bTXXyt3ig8KKM8frV4
v/YeAAtrG00eLtZanT3opg+tUz51hwSV9+nBQHBy6x2B/mHKNI6q7eJWsFY1
S3nPQ0iWAoNjbVbpkknLTB9SDxuCrkMFt0HTvUvBhaw/msqTChRtt2RfLu6B
tvpFCgzY/lOgJLycZ6La4Di8yDyA3e3LP2ONDvj5CmZ/je+ZLpt0+u0Z2vxr
l42BfTp4uZ356tkeATb9QFcbmN4hoT1lHwMejnKisUq1ijb5H7MrHny36VCp
988Gkrbz8vf3t1ZGRnxJXlujw8mEPILsLsLJXi+t++r9H6IZpF7X1oXXVQiL
BxPvVghnxobwcmm6L06Jp6oGk901JlgYVN/AYo+WGHlpOyYt3Ayxc6qnT+aE
ztzYIWD1CID3ssI+AzS7lJOfAUd8f2y6l4PWl6X3bHWyQTm2iu6K2FRaP8mE
f2zEawPBRB1oorV0enBnqSZeZWrTKtluk9LGVcbkJmM2UGbWNCZEkPBTx7Jw
yeNO+IezKfLK5l1fiMzuWtKT4njUlEOIgncWGDfXI0RvdfqCii5B8yIxn0qW
l6AH79dUT0ybwYY2q3yTsW3SMQXqCnJfbVd3vwhO9gxe3tRZD5ELs/v5zXHP
r9MYdgIJr+qKVAMFjBIIMj5hOYmn0WPbzHRJtcjImsjsgYLTQpaQuWKUekq5
IIFHCrDcNqcen97XB8KXwNLlARjdsck1wTXC0/tyiSam2Ud1JFg5GhWUoibe
Do8+RMpnZkqNIWAYg8/pclLJHikm03o0wCsrVxN33QhjLErr38l1nScw2wIg
UfjJoLPe4z49IHB3w1m39GzhJJPSKMgX9B8DcK/eJUrrciI/EOKNOKkxxjsw
PVvj3VEtJkF25567C4ZhMy+GhUcrk1J7e/k1jupxQM2TlHQFcU+A4F5IjQic
UNzwKbvNc5Pw6ynitJVaZhEIN76A5XnKoxe/p/2jLn+A8F9E/UcQ7cSWQELp
lux2GiJGMo8fQ7or6/YrFAqNWwOF5GpBeAxMymLCejXDhrAziMPsIce/OaHu
UTPc1wXWRjWTBmDQRuDG+FflvA35Q9u7u+9MvbrZTl6M6PpklUWAqnMo+UWI
PjzmHrGsRFes7Nwu1L8xj06E+CqBAqZtMu8mn459bTfFJ83k7Xw1bgSfNJJ8
rzIxneJkzM+9f7Ron6DDyHaKyGXx06k1kY9PW8hllVjYwb3LD7gcGH+cyCvk
sWR6myMuUUDrT6raFyxDCHtdOOR3XFhIovo+aU1ZLrHY6/MOSHsHihZzmaME
Wjshl7uj9kthm4bYnlUtATQuRJDjS71DAVRp80zeFfmM7R/vavCHMiF173gM
dOi6wrjMqEQALY84zCx+FldPaO7OD70Qs+YjfU3UZwc6XJRDD1nclpvHs80u
vJXKmsZ+DXd5ltOM3sJgNhrOsOwRoCVTYs8oGS7iys0gk0fd6ZRe0q+TF9Um
N02+TehUfLk7VOAOW7fp+j3V8LJsml1bvLlfobtDmhxV/Nq8DaGBj9RTafzn
+za79whdY/2whdiLNqe8yoHBbmhdDf/qjcZI8PJhOigktgbqEujc/d+CMylM
/LYKzwI1TV898uijW8cmueieniyfIV9UHbO/seXSejb+3RsPjqMnexQDMjw+
bTob3wcNorWqBkekn4r4A0fgkdfpxb+meDCUea+5kb07akRgbKf31tlgiv/H
ofMb+7A4WRSE0saK6tin4y3AO9H2TPgXnzBrkIq2vDlqPAHvbyZCdFC4drIx
Ys3qZAM5b6DPsDJxSW9Rqp6VZ3vbK91yaGvReSlAzG2rmVkmwFA0eKZFooxU
hMRE/YjnPvnvi5FdNBVVagYTZuDly5aelUoXSGWnZs+gu6HVuZsxRZ5OiRK7
TKZrZaf5VvhSIF1jBux/aIrOwnLD3SOwz5dRCDj5PkQ5LqXt0TMcQ8deAz/7
Zoh+b3DS1OXbzqnoon5pOyTvGETEdFmm9ahllg/9qrZF/SKp6MlmE+jdk4yy
3KEI4epFLMjUv4+q+aLxygNJZOUO2BpjHMfJ++TUJinJxY9COZPtCcPoacOW
IgBhyo2rvU8RPdVDgmWMmwvEcNKuG7zqsocMP/aGKvgLdiYRG8GXcnEId+Lf
fgHA3R2/tprYX3XufWrzfEyOu6GCgXVZM1BTjXQJXDfcOjUZca/mVFkF7JzT
pNzDXertfwJjGnI6kJo6e2nHwdeThtS/TtQpHS1CffKHxCVV4vtIDZtWn3Bz
6pFNalLMyG5a+nMzE4znozAlkuN00B+UNjw6EIzqdPkDgXNKDs7Z1FhejJ4G
PnMNr9qs9q+IGSrDTXa1D8SRK/avTId094b40Ag2sPDUAx1EYVQbDImRda8k
+X2/xubaKknr2QWX2U2yoCH4eoJQGq7jw1/sQNhlbiZyD2vgxnKBDxhrFrZ3
nER2StZwcLY5QstBb1tXutpH7gxAT7riLBGbsbCVG62ERUDQLOR/JvQ71TBh
ykWMWCn0yvSKQHvHhq1pQifsl2ZZZhxz2vUgcxmrSziPagPXk7erl1fh6HVw
Z5gdrh7lgVVJ+339uXwRhljywsx2UEXQQ10256xeA46OLXTUtplufDcsr9RO
NT+REO0DMKRtUWZIUU2tdBT/3fElXSS33ENB8Au2lwuTrR+tifJj3uYAAKUH
JfoLBgBurHAnVvQLOXBLocETzyYX/TZ9H8eRewsUfgqLq/gOtjEjRSydUWS6
ic+KaKb/+olOYwkPrxmIWHcAwLhae3HpawvoltUTEaQ/90iYUu6m8bbFdrIV
x9V1iv7s9r9XDrYpSC1NXPd62CI0CkPI2y9Zk6XeFGqKF3sb73CS03GhP7WX
zChF7/gadHht5rsCyxrPIX8OuT/57P8yw79cV3pfMwKJjUv9LUXxvnbauJvH
ATgMClA4eSmqVCzNHar9/dP90I0mILaZEawdWBy7QIKAKSSTTSmjPrP6N/Qi
y61jfjm/ep3bjUoVJCipgOdl+Z1UDfsiDyGG3g45K8tUYvFaX1FhbJ2zUHkN
kEYkeFvKzmjDn/Z8RXvhCYcO0traMp68cMEes6am/o8NFFjU0lZQrLpdY7x1
KEzqr57rsg6Ii6W20KoLm5DsoMKc+KRopNgOyNR+VOQedOIwEc9+JBM4svNv
d5yL0kFvCNzfU34xlietEtSNeTbAXfcbm+68jstTuH4jaDGYove3Hlh4nHdS
N9nRQimPjl0IDJDFhJC1GuWYJ4kLdHui4WT4dnxCDxB/ukoe7KE80sa979tx
42l8Q81vODsyu+6EZhJd/6Msxn3OeIgYzc4fqDkhPndbnJXWF0T5waY8ENqq
mV3JE1ulRbqWchDMr+vL2sUGvQ3dbyjYsNIG8LsnZ8Tors/8bINSzIaSabco
8RTzjQHY0SV8BChFFTlyjtG4KQbF93H3nYCqhwQjWyoQjM9ybnQnYOr8Ycnr
w2FyMbY4ZDCT8Ug3Dg8j4VQQXCztM/qZZib6XXcPYnf2HuNrRSNn6arrOA+b
3iPlpby65NorWpFAXo/OrLnHtFwXoTGePP6GH+jpvXOeXwVcaW3aUVjAbM2+
kVLBFMR0iwfN7pWev/F83PJ0MuJnzQIFG/by7Bt43PeV1kpvbzV4A+x+HDX5
1PkzSiUDeAYhNIDKxYT4fSXjvOW4p5/MFZrCGJa+jNnrTN7EIDWhUFgVLEuo
D1zlCYXo9gd/uUdA2WKoBfrbGQj/44WMaHgIq/+8EDcf7ZOCRZdmklfy6CW2
Uh5VEFkglIZtuIsfHb+ThmV70CkmomggkIEHZqsWbc3icKjeRCE6olq7oUpq
bg4bX0G7AeJgt0xfkVvBjuBkqyOnlVDQATJh/KqkSi9wDbA94yHUCK0/WGig
/H/EsyPz/jKDEwd4VlSilRipN5OrF9qIFH7u2Xi6iKEX/vYkiDBEyPN4x2cj
sW/NoYiUesjNjoVz/V5HyycmRX16SRoMKS2PrHzdM2il0VgrT9qANMy740lv
diZYmI0qUTgS4rF/P836uhA6Adv3rei9pX1rjCseiu3u2DWCx1ixLQx/K9mW
lJJjZG2aW1nnqwMhyMCCkWxtuTIcXFnvw+l0N96YJ+2fIDi33nuYEUwg716j
uD6Un13x+WQ/Hi7H1SVRsB6fxAILzLWDogj6u/hKk5PDDzwfLT9zo6VSs8YA
lMhX28XO6dzf0yxmt8FlNBu7uwFvhOu/41pVvu4/ZArFeahGeOUrCpa4Hul4
uZSBPcyR1uLtJOjMSvBfLF7of0gr8xrEOrCCkgIqheXtvxB7FAU2mvgKTyPk
TWlO8i61HLjWeVqLQqPoL+0PLQbRDdsp1ZqSeTqnjp1cIQrOxO52IuevkpDs
GQar8f+0l286QPJAdEcnkgtajBOTMZOcFaHEc1ehbKvRQAWYLO/cg5vdxmkN
Zu+B547YkGhIOTt++Y8m5MVZyI2a2AkAkC42hoLStWvhX3m1A+N3Hw4qApGT
6odZZmUj2wFgHcO5WF13kCMIo+opTxAK2qHaJTnCzybZJC3qB1QVo0J0aKG6
SIAuO1r/S1ckrpUNnctIkwvz09yzgc8TTfcp2SyH9FItFhfY93pFWxE2UzzS
OqiNVnv6iCCJAQcx/CxjC6LeeEfgv3wmFFHfw+U2PFERqlfqzNp4zzcezyvH
kN3eF/pJxMEkwDDP3S6NfX3XVjxR8p2BsMnM3cGX7YW+zWb4aHtl7pNrFzmw
rDObMfu/2mFq8LrMkiZW9xKuZKaByWNvzsj/n1ryBiUjgYdUU+C9+ScsGvfa
+0W1FR3HWSI/OEq5xAmgrWwv8lFLcQKVz05kIb5nUuqYdKnCjEYIfIwR8hfx
N3vrPVBpRP1dKWgEyDuswLKLlD8XhbVeew5ZOXModVPciBSwurI9nw9FUNsn
Oh/zb5VDBJjP8nAHabM1Du41IvxPFuEvXXU/9UxrxG1J6h5yZMrOR2chnR13
1hy78YOgnl/crETDRi355VrwxiDZ1jW+jhmKmHQSmGbCiGNyWJMpiQ4C3Y15
yOBuPJpGm4DPvp/UjfXZiQ2UA6ZcW8uW7WhNVEvY1LzAb5l73QqXuo0OcieG
z6FOSyUF9uXhx3sEKRhnKXoUn5+JmUP/3TGvNHoXA8YN6Fz1JYe85n62m70W
EpTKISNazi6zGcl3N3t/bXQrfIL1drdVE6P8jfJQjEd3n/zMXDzk+n70A1x5
aZ5ug3raTDny7O7jKeN/tIidK3HJrdMlsWRGw8sMTMSNRAiH23649ZZeApNr
cVRpmD3cte0liyKjb3fYj7o8qKUD1W2nDCFVDpFtlMddd4k0pv9xrfxSuL/e
5I6td1ddBTe+CztCY6Az6GTjkk/4raUpYC7j5s/XBxAKMZfdEZUs27rYkl7+
naY4JuBprHSwF+e2DybDQrZwBQUuLh2KNlZwrPJDUXnZJvMrwXcFmAWKOueM
OP0QW9ms61LSZ8Co7/goSrXV75i4HM/XjXITQroXo05il3nUm75w6psaYrqn
sOvq+iijcRsnld82WpGpV655lhx3Ok/9SYV4jTRtqaXkEfNsEuJj7IIaRsit
8TYRW9G2fNSOL3YtRYhfjignsnIHgfT7po4DL9F9R2Eo7Qs1wTdCG0avSiV0
Zd/elXrO3eOvVZEl9Pi2zrupkzSp9CHFHEdX1jdtFVN0nfe8/qiNMoFuBMFF
FgBktIpsT6Ct6pEiW2INi+AH5vKDfCUPUanP/1/2mL5Crd31mGbmNEbZmnr3
JvU32rQ3rn0rNf4bTby92+AyRrDfoVMWi76yUsXZd0+8ZDjI5wzTuJMAnJ3/
8yc1PHDeVfIzXJpg909mlsfGtDH/0OTdxByzDmQroy4waUC3HMd+1AEx59DX
0sKsH4ReIQbZal178Hntkf/1LTS0zTs/D3L6bpkInaado20DYSiCQwWh9M7F
MDQuRUfgi9M56LnsiPYxSsVr8xtLnNoTtUYB0qm8ihj9WNF7ERMbMK3/yRbb
IEbmSjdSfaQ99/JCE5223V+V4sA5T42tzWFKJN81ctKxU1HTwgIXoIsllEGn
JH5ecMo/W+2SsM2FZ4ZUuLbzZB0Y8R2rS6Ev9F7P+CpNzHgIKmMMoj2EOmus
XmZIWsjkrYhl5dm84RST02XqjNczhjtWZW8Ad7yPaXWIwipMjNscM3p3XvBw
1SJHtQK+EJP2fu0G/zo24pJNc4D4vxpWHs2Oy2lC5cFTAq4KUJHmGTmPrLXH
xtQGQrOYKy+RzEt2aPsj1IJnfiZBBNSNxI1F2eMb8oybaWfTVVaYfSGCDd+I
OEusYAGivsz5UtY+aBSYfqCkOrmldBKw9pbfpGhvR9zjg929wbwjUldYR4cU
iblylGrCcEeMVbnpu4PXOq7O9xJIvNbWSQQDFVp5Icydv2yOr5E6m7WXbgOh
6PGjqR0ELNCKqgsv9zmKzvkDStmuJC6BC1wuvwC5k7WpYvvDBUpZQVui8jE6
N+cCPdezxAoA6Ix9SxcS0yp7X7DpBj7Z9QajNGi+UNM4w51JdgRcbqOBApGw
OSPqgrA91f7qtcgxfDCTJt7JFQSimkcf8IldIcZB6ZaxLoEJFQ9JJobsZjif
/RzAUO8DGJwaH0TJZStNJQQXbijHYQvIIDUOQBh9j3pMdCVc/EUJzhWME5YW
+sCB2/3brX1xZt+lL9qWhSgv9iVU5NwtWrmeMAWXXWGdWf3hvq4fE0NAZqnV
14Gq04o4Zv0+q+Lks3BuTNQm2mujnqZ4S2Zo3owSFhiTG67XY5vBl/H/+DiO
Rn4QC4KvkVxkVJzU8wT1v8PJn+WuySsPe4vh79VP9jasOWGbW5UaCL0OZCn7
cg52I7OSb6lbQvgHiT/1GKCiTSikas5OFnkhaMOQgEuTblTYGeWJUUzTnhYm
bclIeJLKnVCRn9mMiUm2XDg5+4Kt1BPDYVzoY6uuYhJl90lYev5SWIDzj6q4
wWezMWsbDVxox1OPyLY3Gd3ouW1dzG9EdYUlrN9HIRSC2YCuXnZA0T75SHJS
qLBZyKykSXUzV673J4yerr5/pxqfw+ekxBplOleGwWRB3wkHnDgsZfhGBnWD
DyK824FSzpMeIatSndHHqkcmZFyXrtqyKrqBqbsm+Q6evRMhA3h2R5OyiO+v
iJxV5RrUFzzYzpTJzrBDk1FWrfCD2se75aY+EisNnpW0Gbz6dj2IuyGTZCaf
CvUXz8Nu4liAbHKHV2Bo7e+TQ6UcsBFdxQNu60twEvxbyMkb/0YudX4jTgzw
l+rXdwK0Py8i0dHPhS0CCZiqBiZs08IjQQfRf+jCFwE3Uz1z3U5Z2ZeRpMwY
eqMNeqNGuWFWslCT2VRUoaz33MAOoMkFvngemObhYsBnQbGcL632VWLV89VM
zoShJiTJFudnGKFnMVKtxvBvR83N0rD59gmgQYbgM20K+G5sETi/E8fo2Kz1
/47cMA+h+ajYIeIkeJ9PGvREtdzJFxNF42XLCTfIqn5CKbFQAXGCtzp+suCe
AZh3BvaUU9gdab0T2p1e0ckOUyGjDSJeM4tKeyJq1Yvx5zlEW4uDjXl0xPiC
Y1QGAYNie+IeN/a8hLi1CsyTotNNnIVK4KrS6lgJmp8EtZyU2ppguLlTp1yh
hqytc1ok5vMEQBaRcGpz0aZODDMeIdbOxiMgskakI7XQYYyOdsf79WVdxAQq
PSwEHz3waycN6moEklYVCRJHZSDvLuzIjQ02k2lkmlOkI0jdWCv0IqUm9ep2
wDBkbHwouu3qPwx0N8mtxMCobxJHzddt+IbK1lt/78nEVa6maWdWzVm/WbjV
MHMc81DVbUvsMJLnVs53n+snRfALUEUa6CCDQo1Th+hhz+q4NVzo9YtjT7iQ
3tpAHnOn2OzxG0nEGF8zs5uK/mOU8o5KKiklYZLGx5EYBmEeH8X99L+mhS4y
jh5ASHWRhMizA86nawzLDYI7gaKy6QHeqhW/6s404K5LzdTAMuW8FR6xlNwV
m6i43JemIkzvdJIK1rJXK/nio8hLHzV6hSAU/qMRd8uuOz+pIxwUrUsCjmrq
FMtRAjwnJ+6Do4jK66yrlJqV8dt7naPR8hhzqzCh3dxX/OFRSA5v/xxTPtrP
CI19mUVRBTzwrXRUG0eZX7DOgyGPvPgZXDulUpQRZlSXQI5A4fp6H7Uh1Tq2
PTp1XzSl7Vj4NyGnvqlRqB8Ft5+lKzRvyrma5naQTohep/G/HpZ/hc0N8q8y
NpGCMqHwmiC/SGWItC4ay578HG10fYV3TYpqEPiSBdfHMchOj0naqT//PbWc
mHFGsLpPaWJezHPHi80K7mu29GoxzCTWPKE8ln5A8BHTaWJclI0RUwf9X6Yc
SJj7gEnYS88RDUn6lkbpfA/BkCbkTHBknon8RYBuJbhkNhMjSE7LwKf0K9C5
UEDzVq4Q23ngCAiraUTF+Xs2acgflw1b5j3xYMBKZ1gmG1CjvqGusG3biTzs
fY9m+LbgjDXO+kb7QewtBk627ZOrRLpK8/wmr1ltx/SYa7UtYlMsZ9JBhQFw
dppyL1XxsiLOkAFDUeGkU8QqqzH9PIFg8yAIJWvhCndJdPf1F4WiRnOWBRPh
HsurAW2paJ5Q5xiLA9sGFeKssYP9ZHKhtqAybhI9uYEHBvtK5Zr66IR7xvz5
M6Ka8piw1IQiyxbrPoA1GdJ+Zcp9xeV6AaOIp9FbeuxHx+gX2rAyqIEl9LEc
iaXXJqmh/xr7Wm8XCF/iVTEr99cgKpJ3EKlDzO6w7cF0WObMm3iyQKh3OE5S
8llfymWUNN++NULlBPzMLkYYQyA4dsokaKEP4N2Kh6di/E/vCDwaKdSB83ty
deuXno7AyWxouyw/EQWZG1lzUWuUesCExQtGJHXM/AcYRHW/DNSY2IU47BwQ
52+1tFz358aJzUIEy5r8hzhTyFrEeL9dcF+Ex2ectDc4WNYY+qDGbPPqDIBy
I6tNh7FsHjMF/jspss0fD7bUeWcwszfr04jR/GcvjkWo/OIImsiOChDiWTIY
7u8tSmSJZnLKXsmzMy33R1StETds/z9CS+FDYJLZy5AmWxNKzQAKneJFWEju
8bGMicV1CLTgnG7MMdYrT/zQyaYtp7kxEoxSS0Nb1oLgXkNa5+JkMs7nUluA
LOBzicK6qZK36kAYmX47rlx0k488jQz+abN1rZmP4d8nOS3wJpHVf8AgctF6
AOu9TgUv/l1zvCoM+k7gi8JmtUWwjsFxIBcoMh9GHW/yCG9mAVl/lse7Gy4D
VYjsjn+CGivPWES5AEokUpWc7UG1oVavCxg+O77aOxMw4JCRu4unWHdtx9aP
gzk25Ch1PqxjZmfFp5aGYTzpSV5effU+NrIIawXv4WlAIhyzclWgFkTuoC7u
7/XbSJ0UJIPVo8W9tuQ3+O8ksvyqrDKKWRtLbhZPUi4dZ7ReiJYuJelSnTQ9
fpitt91ELY/pCcjCJ+XO8SrM7aEKx14vs4WbCGE8767Hzt20cNdNv7ISOMv+
tFdofgnr5LiQ8tkzXGZSAIiiVDGlhzcaYtoGVIEXDY8iNaPbyRXBuTLEvJoy
FGJeKV6yKfvw1w93twK9y+q0/Y7G2/KZDwPSKtiZDhYxYUR20Uc8Y5JjbTaf
1LW8DKh9LO5GEfolgS9GKfpPDIK/4UMZv6polbC+8jWPO7WwyiJzqwFMgWr9
+A5jkh0WOv5qYIuPW4X5TLXAlMjDKj/sU5Lo+zYTEtTAL7JdMlxPNe6yyblE
Ku2Owv4laLgNUE4s/TN2mzO5ESHkie/HG2aqZG6JA8i4nOIJvxO5pGF3MEzr
od+E+c835U3OU+Xth9u7h8LKNldGtHKicvK7KYljjddNnp0+nkFJzs8NB+Fq
w0xy3wQiJk0p0fuhosH1El+NRWqkZD/6xA60dZBoXshie78ipSlMASHA/8Z+
1YkXXfdtUjM38UsLdf/muL5z7tobMKV0HZB+XFaCOvI4E8E4c1zwJSXsJKhw
o8ApxvJkHpCZo2kf6k+QWQrEEXbfi9qn43s7/kLFg4lDnF8yIA0spYxSrq0F
i8oEJwp29GRj5s8jT7QCKUdrjOb/LiRJrCggz3eTqNfVdCeBEol8x2785/dZ
NlavKwe1netr78OGxc+GVdrNKosDM87UG2MWEc20ap3nljTas3Xw/F+lj/Mi
zSVaoUIl9i4H0wjqMNy3kNbkOBW7EyuM20Utk2jjGhf2d2PzOpbOvRrKdxSD
EB1zseIxfeuikWg+W9tfIWBINUBMn03wfQYnRxMibpsad4d+eSfvheHEOixP
lXBjthorEBDEaQ/DaRunE/o1Y+Sc8anZ60ojwxwbdH70f27+0jO99RNNcRM2
I2FLRp08ksf4/e7fZRCnmIHK9TAt1HCTlcS+ZLr4b6mSbyNcW6PdW/tOkKmf
fCceWjR6fzCraMkitaziIUh/PuurDQz7MhgJEqZUeqfdJnuakvz5r/IpV5nG
UGJXevU0uR1yWWxjKtAFfnp9Ay464Rvz99PMCzK89luNwnc7WTBqg5XhL/Vq
zhs+Gh4cWuDLrELc1kOOH41gZEGSZwmy8/FfXdvFluhyAuNRR2TOt32RWkIU
W/KVIzPtZURQ0M445LTUOLrPm+IxXwabt5esos8J1Irhwl1APg7BiTUiX0fe
mzFVcqxy+LN8OibnpsUSEqV/klBxUtaAJHLA6LUSultF8ZCmSxwsyZUMIs9w
bRgS4/95AcMDXxBn+IvU+qKyNJtR7ceBKHDzQfWQWfkC1tJJTthYojiBHteb
YVT8ObaSYB4Iy5BCxcYXFfE23GIuBnbKySlpkccpPDm7kHR1iSSW9uAjk1CC
2iO9yuy7r1aPFUILJd15HTxzb6fvf+UV/FpJWASwlXlzzAzAgVeOsUSzjklF
bjRKCnZ8dvKUYfVhgdyGxZu2Ko0lGVXilASF2gRHFMa8YrZANH0vNkonozfs
2H4ciW9sW1B7HuoWmaZPag5EgnZCzycSqscaWkC8uNhUiHiI4nTIkojcqU+w
wA5Ma+cnjTI4yEQ47/Wb/gDP4WxeYQ6X8LECDM5sIOICn2RNVZorqgjVcehD
IkTtVICA410f3Mv1YkzcUB4iR22nHFF/G3j7Mi6jUcBLjGIDtzdVNmqWRrNT
wAyHTCJJuP/wXq6zVY/G75Qz4kfl7dlks7Nt6KXVRupwcFMqMVWWZfdycVXj
TNl6EU4GFkz1VJ7uIZ6qCWs9qfwhogKrGHbk9IuZWdTKdhq/Y0NZhVIZ+tYe
fy5Il6eE5DKSDWpVLn0BqBEw2wRTNxBrCzKyBaGi4MJGku/U3D3xr1y6+b0d
ocatGlBjEtIjC09crWYHXLBSrD01i2XBg4uFfEYAQoaNW54ueTm7D+lU06HY
TDKrkrOvB81K6sNp9sMEp7o7e0iKq/1JVnIYGh/fJyh0w9foF9by5hNUZ9Lm
dkIny8iBNhPW1V1rgV46x5HVUWp4+4VezuDJbxlH80kRxiOqz5qdQ8n4Lx1L
gF2fD02MpqrWPdnQqyjuexKEqeUI3J20po2CNOx7dBqIQ0nSV3i92WkqNg4U
nCm+KP7gCF0Re/KhY3TqdPuxviO5I2naMrpRqV/MRVLYZptXKlxrqENGV5TV
r128qruchwA/Y1cvAgecYRv+i0n2FOTkCcG5q4haqh+zCWpc96qa6eJVnwmI
lwmDuNvcA+7sqQO/qagOLiog427SfZcmH4AsELUI1lN7JLFvVKWn1GCOI89L
Mc+QYFuhudT9X7xSKOt+iRpRleTzsL+ztOvTeN4aKUe81UXShhWSlzAjHH7B
w88K8te9/ofFvki3fR1eAIh+Mb65zww9SkEaBvLHCjT3LdVO24OwCfJ/qB1w
fYTrqrEu5CUDGXln7V5knnUid5oM5t0rTrkUkMkDfEL7fVnvJMpOr5ll61Jb
IPpoJg0tK6BIS5RbdVQtKL8XEKlJqrg3Gn8TkeSkJgqpM98bGAsIw2AEauvv
jxn43IBkO72MCzpxvw+Ktf99+wmFRUQs4IFloVED/WUvaa7GW+klXGP9GS2+
KMitAL3afQEJ0D4ImkdpTgF59hh0hA70YNxEJkzvFWQ44z9H7oxVOdrOn5r+
NitCoaRxoGOCcKp62uwxomfszpElP58nb/Hl/MCeeMpLneK1zuCElZJWkq70
Qe86A98+inBL5p1srh523nnN/RM2RW2CXvSFmJdQaB4gNwFl/agfDLoh1bFw
FCZtUB6wgCYa2sFMQVt1W46wt2/0DOYZPLBIzmK4XmtY1RNuU1TCpFQLRLZJ
QWkoI4X8Kn5/JB4PKlDSeawezN4QDPvojX5oyf6HuOLSCg+u+EGN4LPtPxHB
4fqBDYPIIHYFVAzNmL44Y7qVixMoS2b34mb+sdIhQ9SsL18/2GIPV2JDxD8e
RMVS3jDeVf/c4USUj+ohYTXw60GQijXVNbXdiKT27Ph25WTF4jOIGRH4PdYd
qMMhejfSH8J2TIJX/q3/zxOssGr+7mH4NYkUNonA6l6wdlKtlrbVFIATnuLQ
/1P0M+Vlri2dpBElfQapn73ujPL1hBeUWwJIGZyh1RervJK4YjHIwTOOSGBV
DHD4FH9kkeC0y2+DQZ5OtlUueZs2VBrlr95uTUEok5PaSBtna1qf4bfp2F6K
InZpn11UF7042MKxb47dm8m6aPaVrTJrMsF2CMU91+0HWfYLTGytxOe28tIS
SjmZTV3piDaEhDxR9IaLJAiFoTbxs4JAse43n6sDQgIxAPfxSTW+rFGTmGay
k8ip/rMbHoLbgSDXrjWMtPzQast3Jr6KCml2itPPJsjC4NZ/peM8ZOXv6RXS
03G9IvEK+NtGb8iGDCBILFRQuNBSSVCOmU8d4kU/hu3Ql6A3qRkEDKYEmRUk
IQPFSAYloNEBezreFIheOa9kkIu4cAgDbgN3jM1QvHDVzk6SY/2jalROo7Hd
F4sKiek2UNbFan04iZneUubScmr/9Y0/mcusMzz36bkI6tmkiFJv1vLOSvT5
S5QFpCsK75yKbwvR5GY4tqF6d2xWMHc74qLW9oOBXnxvsvkHnCABtL/2u0AC
yd0ezz1CR4NmbaCxnrHU8We2WmeGb+8aTjmHPDywG5P1tNc5NpjOldvnr2Ui
JzIqzXdFngo2nKH8L+EA5msil5mmcmiHvLz0dB4qB2eUyc0NM68mJf4+leaU
fZ5dsQCAbxylThKNVy0XpjQ/WRaiN0tP9mO/tIOIQq+wSNlPBnnMOULUO043
gjv6xblj6aW5v9fal7SlZiIoHhQ34tCWH9yI2cvAYJxXsuEYiU8jtNhWbvZJ
3aKLxi0YMegQDUBISTCsI6Swb6XW0LXiG1Uq6pC0yg+hw4ynXrFbf1WkyC+C
xTBXAKzmoYMr0fK+ivf62Mh/SwG6raMHsIBCM1J/H5mCYJqTM5KEL2UGSHGm
n1CEnl7GSs3dxP6C0LYqb2+QLEpwqgz9DTXkY7o9qGhT6dx8INC7citBdjpX
qO3Md0/MZMvhPxk8dfgtP4vu6hrT8618pJgCkcrLAIlKEoNQ+xpYkOTHtZDk
+7oDxhIZZ5KFy76JRqIN4ITvaVUmPJ0mc6lGmcBGgHoTXATbL9pmexKKLQTp
MLiJEtZBEWZpxuJ+ATcf0pJVU71cr6/6rZ71F6I2vCcwMU6cDADeKcDlB22W
xjSHpJEQWOnpytXFde/hcGDd9PtITtHXRtCPI9DysYUDdUHCeerbqsrfdr3n
HImPtPMyE9pYV1nFX7JP9Eq39nuCwXI8/l3cHznEDzYbJxdevnTJAJcH++vG
xFfzAX+btTrV7bwJZWXtY4tpiV/ywqsE1t8bpmAPHMCdmCd6P4X5gLzLgQfE
n6F58Ov1rgbtJV40oQ9uAh0h9e4Pj2rHe4Sl1oVjhaB6beqILLh+0WIK3GFj
Aan8xRKyoZV0FLXRaoRA0Xq1AI6lhV4/AF3uG+vhQ0mI+uE75aK72KVr+PU6
EIP86c635Uf/HrCxGFwhaz+2steWyX2N/qer8laO3af8IsaajY3GpVqX6CYJ
y58P9DK5HYxXy8ZnFm8l1vav/eG/9hl52SOy8B6GHRlMCoZbRRWb4jG4JiM/
swfphggy9O2CwX5CytzZYfH3T+4RbiBi0hMxbeaj+/jD/QgoKFpkKm6UVC5W
KbATlfN9jEc7P+kb2McO+c8OW9GT2MygGDBWz5W7Nnlv/7kR9JPdac9mHXS3
7aecu+jStLYH7VkAR2A9seivozECuulkOH9UZnA7rCA5mt7nlaGgesYHxeY1
x229YXTkK7+8Y8nobsVEDjowVZK1ONrLoW9m1bFPKZ+DvCg3WNunbv4axcGU
rV98HLpphpfZfAzQnGmiCXEX0mxwG5T7RJlhoiYNLNOkjUHewidccPhmp4za
Ut6kiPI6DisIEXn7oT24bhmnBY5H4GLcegIGIO90eOiKDTKWTAqrNhLPX4XJ
0w3fZkCb2rWbO+yFHFO0Q9SLcwMx6ScJbuPmJr2227IUuGPqOeOU4a8/VRFH
f3x+LHeolaOcPrh20sYBoV/tnpBsN/JwREutFM5+tlAakvT3YnL3vx/hW+mf
BMy0Y2yxFK+tKjao4YH7GOr0trWEGNTH90crCtHde3Iw/AiOBxeQ13HzUMkh
qx7PIeAWjtEiv838hhJj/x9D3tRTRdpu378dio4BnYoNN3fZwLcYLmU2S/OM
QGe3hGUGBSy3MUN2IgEl78QfRmKuFDxHXlW01v05ZAm4tWor5kd+lB4w+Dn5
9E95Srye32csvU9Od6uPLX+bCJSaevZpdGxtKHXN5EdlKlCc+/F5HqJ/N3P+
WwRL1d5tOdM5oVI7tyOwiz0kaNTd46lEUDV57lzcJ1Tx7wadAuN5+f7y0hO0
FpH9NrJbzoqqLI0XNUaFX6WOMKxY/bOAMENL0RhDFOhlG6vNP7/k+M7+2bFb
sVwva+I8MazO4jLoL2wB14EadNMtCxIxluB6Q5J3HeSIJAVsB8dQ84pDZUm8
ujruQhoD/ZAl7TWisODS6a+0F0jkxCa4TFZunAkbUw1C7FiFJPg5fsodiHiV
mp7a72rFPxYmc4Cv2GVfTKlk2AKE1d/O/XuFsQGM8RacwciEdM9bi3wE68tF
1S0zdJB8NwFcghpJ2JvMc8U1TOWUdUDm0YUzZXEUBmaidMa3wb6R/PAnwrZK
wuG/lYnZK5LPU44V0tl+JuRFdB5q5ghbByCOtMGGVktWEaBK63txHYYFzDsP
JIjISDKiTZzINSJTiq1hGMkSJXhddni7F/iJ6/daODbvI+Q8jEVaYKrplpq3
YQWJ39tOn9uyYkFyzJxYBlGnKrlQVcrc7FVX0eqARmJAKu3vkNSaU0jM/Tmi
Y77AxEqAloOG3DnV0lfn9RFTDNLNQxby9p+EmgfRLqfpCvF/4yPgQSSWAeHe
6bSkZBcQYm173cfw6a0a3t4FD48Ixzrkqbw1+Gy87JZyqLpXKZb5Yey6Cmgm
FFKV8lsIrvZFlQGdj8JEeH1/eEvkPsoYoZU7B+OJW7wpcYl74BSfBubJylyu
yff9i6eNF+O9TOqwiDIVpWdEN4LJ+aCINpLW4f9yzjaJcmdhJ2vt9uKPb/sI
AynBBrQc1G2FY11aWGjhmFaVQr/zN0t7I+5n0Qpo/dfCjE8eImsI7SsVJybs
ZZJPzcIfaaemEpLursC5PcgPTI38YQfvBQPIglZfAhnPWgEDjkhMIk2ON9VN
D58IphDnH64CphEgMmAnctnxp0IS5hfats2eRh+SkCOGXv8hOoydLX7CALz+
ag2WuwxdsEhoTDut9VaCjEPHDG0stJSXSutokYr9p3bdxJuMfmFLneujE+95
UikHKQXTZG/0N2NkbbMG5+QFPVKJdxm5+vAtAUmTbgrh0mTXflHUq3ZSRwOg
dpV5A8xAEkNoc+OrM5mcxOnUUB/LsYLwCAK1w86f4kNiLw/q7KtflG7pQ5ub
seah2iN2T3P0gmTiksh+09hRFn+nZ0qWtvGJJIQHEX49rEBVQ3XX3ZM9P0ta
Xc5alMi7BW48eW4oYo6/FPVjuuyAiZaFxN37v0d6zf9cqUthKaqSGOnrXiqH
P13ubClNmSu5g1TA7GnPUXXPnA3jMqCnW7dG06LgFG2RGpAMaw0lf2mQsw7J
8c1HIrueII0NEcTTR7BeB74WGRqWXf3LHnZDT5wnk02i9UwmRVOBWx/3oMid
L++v66pggMYZUMTMwTSZUmVWWo/5xXcCEf/wzl0QTMdDQYjLQlXALZVmB1h3
nUL6bg1OcaZtAbFTGhHA030W9758H4FyHwYn0kpyyU/ygH6JDnr0+s/3KHhz
n2cPTexQwcshgQ7KBx8Dz24gFpnn1abd0Myi680oT9xgNXbvUWqmEsVRHhKe
YQrCNAJfTkls975J4w3isydjDgyf9xATkjZLo3niuiiuqcIne/2ItkZO6DVI
vZ6+VfV9hCmldRErriboG1ZM2hQxZPB3oMVVg++OV9vzqmSb0lXWkThRrvfL
xvlMN3wRc/loV6dmzPgobNVJyHcp3UGbZwuWPjdUP/imDSnolLJPQXxsNuXS
m0gcaCwFboUAI0QCu70labOoTHz0gjDK27+ADf0DoA8oiDoK9a1hYexL1MM4
BjA/FNIOZEa2h+QXaiD6kJSo8rFRFaUdoiqSKREOGyAxj18FNHucblsI1aBh
iJVeuist3gxOhBEpEf4GjerXu/Qn/FplHBtMi01ApgjZ8/56cR7wzIWIHxEH
30cJ+onysjtM+Yz8hJLiEbUzFE0TkbVlZqlPHWurBOgCdhpynbCBwL6eOo3A
iPFnrRK5AbO+WEx94SYPf2kNC/zhNHIhK7jsjcpPSKd7WZyBHiqY1oH61sv7
d1lr4z1oR6bdOR6beleYzuxT9mduORLb/tDbpv2BlfFEIHKX2KLr+gvpBSek
EmN/G1ObsSYoh5dCA3m9dJR9fKck92NM7hsBzHPF6dfxVDm2WdZezGF26ThL
IXHXq6he3oJ1vfW3Vy6upnxZMTiYWZUXoOJjsMnrGCO/8Nv7B83VbiV3360w
yvwtZcbfffd3j+yLivLxg1U2hXpYbaxmi/fuplxEzf5Z3D5pGywVs+T8nVav
uKhylYII6trmkIsE5o1+FwYHN3h6UDDWtuRas2HggwgXzw/EWlPKKgPXc2jB
TGHlY+rI1doRaXBtGnWnglExLFNn26qj6T7JO7M/eW6iECgZ/qaw0kPIgvxE
oqY7SUJ5b4AVR/Ch/yyYrE3AO0yxybfRXmbx9iKu2bquD/ymG2u6jufgGi8c
ubLrXc1vUJIML7iKAZ3q/GJVWDll237ZJysjdCnYeDz76Ib/fqKkeiy83zC0
uJGFyrH8oohpVrgy/g1T9u/pmEGHYXsSHuipOkudJjaxI71MI48j2pte82xC
QFQSGRc8pdKCY7j46e7EwDBntfDq5rExNepws7LMoz5b6tVLwU4QoxZmeZP6
1JeiUKk/llD++ARzRkeeTej49xqpjOXS+0+R5lUeo19GQTOdlG+0x2U4o8PL
XVR5jjaIjGWqaFRjzHDZjaYfZ8T2eEtZLPctOue9FOejXwd0tCnp0uDu5YKZ
xqqe1huapQBUTsVv4TPoDMIrZ2tHgbagltBi4Ll6iwfJacZE0DSlTJHBJTHr
Bl9+0AIws5NpNSDpgbB7agUAnliW5LyejvOUtmZ9rljgFVr7nO1GDbGMT1ES
ImzOuTQ6QfA+G6QOchCh2HjYvYLUyLj+dzGSmUVsBJ3++lhm+C9Dt/+Eycbo
HCuaF3YkX17eZ3RxuZ1Wv5n2NptFqYCQLv0pMhG8+ehxs8p11WwvL6QI8ZME
BuB6n3cYImycH60I23bzWPMDiqZiklvMaR1HGjetM5sLbLlI7mfsl3GAL7Pq
mcT2YABtXupjQKlj6h0lwUN6GQKMwUwSiEK9FBV0HuUuydlhNK2bI+ir7mtA
xiV5RSxWawZl/WHyaCOjPq0c2DrUuoGmsAzVsFI1SLh8dQ6/0DHsLS6zR//4
xE/eU0X6v4TG7+2lLElSH8L+uyARiQvCZzUg3hZZpSTBsIpRDTt1luIT/frc
jQski0AJyl8/HF4SG826I+CSgrZ8Jtzrzid/hUKP74mCzmnEmDE0ykCbSh1G
IeBTq06Gh9fEFwX3mh2T6q70wb1gCHnjCLQtdEPIxPXb92NhFPQNI9IrABVj
eZXwRnsZf8qHAJNXFh6KRFMFcNbC79MAHvwpzvc4/8HwUiPDVeq1K/Y+Bsdr
OCOkBFTXvQA8ZDwdJ3DvFOq26OTLVe9iyYeo+6XaxOAOu2Vr2iPXN0Y3/oj3
XRpgfCPjrNgqi5diBVaYoWxTH458A9LIMgVy85458gMh3YBedTudk+lphwZo
o2YUOddC56cLdWz/sni7VTFXxmlFCXVYpbHrrBo6qdk3G4AP0IPWllnE/F79
VYzytdK1l0BKzgyfN9X0bSCvz5U5UlSI0zvVR9mPBNlpIlz6jSENCqH8xaBC
tPZ3tkbcq49+P9ZwQ+vVppokx6Aa+YkAr9FinjLFvK5EhbcTQ/ZxKYuuHXZz
d+Dpbyqxpp8dyoUeD1y24bfwGNp08Ib05jPWlSeJAuZqVVICOpEFWNNiNCIX
kJQsnna2F3PfcmPLY0lNb2CJ/lFctNrVoCrDg9UohmkKH78QUr3t0JLfQ7ep
qGhf9D+PzRsjdoHQ9aGUsFGMjh2/Q5tggxhkQqhSYo3J7d/DBLabskyN0GIl
ud5RptoqnuwVl7mw2V5RkIBefch0OX9UHQvTMh3IazG03j30Bd/P/RHmNsAH
/s9S9PGox2buG/U1oWwx4dIAtV82u4xPSSTXUZkQCejI6LabOSMKakjiEEFY
6JJFHyXhzpGi1tU4Qc+Ew8l0S0JfibIGRmg5fl4mpulHwtmN07/TO0++EkBU
6qE9UEiKahe6tx+43frVBzOfL9dY8SMiUkU7y+20R0Yp36w5dAMgdAxADtYe
kAQjqFcEBGjeoJFdr6piKpUPjj4l1WaAvDNS/7A4KeYFIVom8gqJ44mQxq51
wjKY979qNygZNTPWGtxhVlzeVXpT2G1C3vLlikSqFEfeKFvGPai1oCaIQpis
Q/uVP9gKaCoX0rV8VjIIByln5e3gExGJyE65MPF8sLsJh+wExJSvNDdtdf5G
zwX9gi6a1CpXotgyCieEEHTDOYBZnRQfItze1y2UmpWRjRwOLcyjet3MEWdE
FycLNAWACwKBmIEMKBSc+d8p8f3oVoF0QYyQsfw419I84VxEUaNoGwDNJ8IM
UxI2LhMdK2nzNEXUM+57NM6OA3NrffsHHnCKL/qePCOhpiraHeCYD7QJkDMO
aXYSfPnaQG1mwwTLj4+cL6bdXX6UbS2yhtls5OPZqdvYFGUPCMUmlHbvQKvH
20Xd+Bu4toAW3ZT3FNizzoHLmOMZzCKONOnP2zPhAjx8YeSHaeATotF0DokK
TgEiUV7Qeq/eK2Rzea30lcbSRR5Seg6/e0eUbR75YgSI+VxDY6mPrZq4XIo+
uPQPuZHQZkWWE4Liw334qqEv5iOoon5DPFMOAAnh9figIeUTkG2FX4NHNKgy
qpdHgNpjiAnLh+aMcyjghxRhf0LVOvfMSu9lRzx1KB6IFKDrxywGbGq9Xrri
NWO279NSwf4q/nqD3kzomzkqUkZVpILnmPstugTXrq9xFNB+84duUZrXqWsk
dCACUmVRv1yMvNxXV1E7T2i8sYMgg9l7x2zn+r3aZmik5XEAQ51ensOSmq/p
mYHjrx4uxJtk9E1U63BDXz0ojBTQ3iwoExwO951VdhKHorORn8gjJzmfaUnS
Jg3u4kmtntn5pw8BebD0GIFz7qnaXCBHEdBARFuPTp/zbT3PW+UxXuCbIaUz
HK6+V8Ji1RDBwDbIXh+c+iy97AVEDTHUhaIAGUhnSFDvWdoGcerWlp3Ncyly
xiMMgUvw2sNXWuMsAzQjru2v+kSkukSr+LbrGe0EZ7DhLkKwlJCyzHEeFHBE
HL42wY2zK3oJenaqaZAJ3mVHAIxTqK9DMrM68Q9DbGH29sHSGTO0UNkJJJBM
ttakkWcN4inXkp68asKjgwmZS96UTXyc1lqMrcpmJ8stDAfRnVnK9nwg1KlN
1/UYAkkeA8lVyA2zoK4uxnny1tVkfCZgXn6Sp1RiFshEpIzmxLA5Al2PIGFB
eocsYsSbbnHwu0iiXJWVuL63wpSB24uyUfbtqOz0qnV7MTNKYqp+2rGV4kHU
Mmm6Us05snNnWUwgxbfZ4oe48B0dacPZrRwGpoUZDHFZMcUd0HzDspAnhWKS
5hO9QJieacK54MIS1+riJOJkLlWbLCoE24rv8vsAzzD5/w0sZyrY06VIcekG
/uYHOCYgJJIPAilVUb+cXuGvn7wtmXHyXvS5NBPBhhn/2LSbR1iJfssnm2/U
+MDhcWugHIxbb+kFLq+aNvx/JdNJmivwTBty/RC7H7R0NIxx9XlnhDBffbRN
NoT4RU6iD4sQWFHFf9QKYVoZ50Pce8L+lh7Iigp5Wrg7vY2QMGyl+xCd4CLG
EiD1L8BHFPJT24VsEFHC0hTUdwq6eGTHBCceuTFttgtupAhGPLbywDA+n6Hn
A9ZSMlBnzy084aEhBTMM4F3/C0a9ypfL2wR1LwEmYCKLUwOrUZRW7iI/Z65H
IhWoUtopBqfJEP7XjdPqoKeofRBn50k0l+I8yPyz2OMDAzQ6paKtoxCgiZEH
d200uKrO9MedYXQXGzZHaFOG4+qiE3oO+pvdhw4H0v19GPRfXHtMMHpLEGT9
QBr1YqL86vZV5E68xonmOchwO2CR+ucCR38jZZG19c+Dvr2EotNpFD4BG5SG
H4ygkuH+OOtEdLsD8EPnaoEgmZvZJm0AEQ/SjbUjHuQpiKRidZRpCWVUaoWi
tVT2oA2kPoDGKqctWAHlqS733FRqzmkm+VmrqfBwH5/CIpt1teaoVKENMQFl
g8aIfV7XYQdIUJWMKDu4Jtuhk7xkWA4ZEf5lfdwSvGizmG8YZKx1ld5Mr2fy
oBxVEGckbiM2oai+BExM/U73M5aHXw99XR3K0MZjyGjYOVL4oEiiwklH2zy0
Rl77OrHHJQQy2vglwiqiMA+MZQRe5TfXlDwTLkEBOUZ2rkDqUVLyRfrJf2yw
Tpadnpj7V7uqh64Bvd6i2tp4YmpmugqNIAvBoMJ+AXztbUT6AzJTJwfcsAnB
m0iflJArZEI5ipRM1J7DvPXqEZMTV/Fs2YwAgXanR/h1xNWaE9LfApXEKR6V
39xs9m1ErgLsjqB5KpQch6dTpZNku6odqBle5Mz4V+tEf1YTfcoPbgFnlUnI
4cK7aQpTEEnqh8RiLGxzXKDqyaYHo1s4beZnZ3SBELSghrlnKIhrFwThTxS2
T+u5WzgylK3FSz2tFLDQljyG5qRfDFONzvAKEBc4ySoLL21vZmcbpXLhiBDu
PA3baDxyXtT7VLyeAx0diLsw0JSDhJ7wb7dguO0UKh2w9o3RK0J9ttYAFCNm
Z2bth0I30m4MWvNEhJH4eKI1eqhCO/5s7bX9qUEJ+MGP8vu+L/UMagoz9PJt
yK5+r1qDbSaRrNk0ExpRtwRpCYFzrpjOhkckoiynk06URdw2l0sm/vRqC7gz
T6mNG3XmxJI9OMmiIfKjCzohLOjENKfL2ndFC4KKufnhx2SY19k9zQrcIE34
QTq+ssymTCdKKZhsbtA0I1V8edbkutiyYjzp/FvJ8HeQ00eOTGXdQHAn4nFb
nw+UEGmz7qWTKnjrJ71eByaMZlz7ETq+Tq3B7GHx7uKZVDsVyLfB2SFokKHA
TeRICgnqzdL/5P7UZCge6kURDSY1G0HbkH6il1an0Hc3MSKHfurzEyX0PE7J
s8lKI5k43mwx4xYcm9Wl2WSY/xgY96Ie+7nQKw84vTAvnTrZR16bdBRTS8dD
Eu9vO/+4kW+AMOVVdo7wVZ0i4PfanCNlDLL7zgC0ge2UhQWx/RqkTHL4j8Zy
igs3IMOEeq1VR39OT/6/1KzteUzuUOw2HY4p6sEfVFMngqhCWqHDG24UXDj8
g/TmwPCWFiEaYwrNjk11WNO/X8lRF8QoWvwNaI+18NTHmj/qFlw58OFi9aC3
LI52Co9m7sgsdprCE3pI2W5azUPf0gSnzdiCswKDl0dZJK/hF00eOQ7v7vXc
gjoBu3HglMJlX19DIQgQA0+ABaN9HUxEHDHMn62g5lKsOVohIlAmcA248fgU
quewwPY7YKIMbFUpMj7N8xq308bodRHN4T9ZlVIt1UuiIbQWDw5S7GUkSuRv
AdhY04uOirzoQbtkTlVXlpmLxFS2QVEnMrfmabli69oB2wN+Rb00Z+UflH7E
tyxqkWnN4i9OLyqgVSq9o+b/FdXbKhJwAIzgC6uf8SAEYf6ZW7r/nRQFTx2Z
VWs3zWByRcPF/HL9KlzdavMtjYeqrMUSxyXkYPEn4V0yVYlPkbu/18WYajNY
ROY6Y1A971FpJZqRzMOVLj5S5A2HTLsWrX4Yp8Fe8FIOcvNlCE/KmGERMYzb
upwSON4mwZH0+OTVeFdW5mQDCvORYdOe5ceqOUg2kWXnl/cj38P94J2R3omU
Kh9fVDRM0jbdmdQJW9Xpn3t+yAXqJm6CLpou4Mk8aInc5p7cS7MlixKR4ueY
oI00gZDJB5rIVnBvZdXcHdzqcL/pGdGxcVa53AnDZ4Mygi8VNIx17O/Z8pU0
+SglgzS8jByVO5leehQabo+ObaV8VznbXlt/lbfJYfGBlu5SUrmDSUUYix+/
JksgR7g9lnwQmfh3GuDjgCDU+yP4ntLFjansUiiBZEOZ3DYDyJvu8XZNtCEH
9FHQw7slU/KaTv4RNsjWuxT2FAYchKw79Z/g/WxaxeLJAjitWHuZFYsyLMNq
qonGFP9OVJTMJUyrHfyALrB15szgZZhIjxXhAgviIV8/s4/QmKe1lq5Eu9g8
FG4TUwudH/rT+ZpyWdKCPe2fjR/G2Kqe59eQfnxcEUuX5Ix9c99rSpKwMFp9
0ux8LakxnqUB9qPgST90Gy2psXRI2833nkLESmTvrUxNEj6mAi2LZvPlZOQk
NzpqwM2zcS0AulOn/4uDOlkWY657mjViQt/+QQ2yasqpnHmaYcGbDfUJ5iew
p9WRiYdaHM2MV35TQ5dcPZiHu9d1ONUsKkKQkLqjk2wsYtRZ78YMk5Hflkfe
a5kJ8V/jkXTU/jZd9l2QA0/RCJw/r/CYH2mHZlbStE1TdxDT7XIPv/lfFc+z
mH6MbKOAijfrFrdq5n0xAhbhiNsW2BFvTR/lpkC4kp76BVJi/B9TlXgsXMDF
Ba5eVdj9KTbLXwKzoqTMzFdh3MY6toX/uJEXru9B8bXAsvmx08okdNoZa1KN
JmyArhe5jYooer0OCybjvS58wGMxqsHIdbjCf/oOfldv4SAwqm1eEx+TiOH5
aDjMf+I8/MVj5LxVkH0bo6CwgMqMIgtnQi8HOhnnVflAi1jB07HwFI1iiX8u
R9Kz/t9qc2bkgtu+iC/TQ8I0AS9sfg1dpHjsJbEfwmxPgCrFIdPdiAmVzPNq
SCR5x/HDmX+NX5gQFzV6Z50y28o1p585QfJQcgYnyFdKUtXtZB+OV6L4LbYK
6tSgRd3a/bQgql9y0sk444ap1fvQdbMtBDOHX6kfeFNmfDNsk7D3R97VwjaQ
ubCDhuPBxFMiYxwSTMzkWVVOoFJBRYDpxxfh2rpSpYbkGDZt69yWnSeKoHa1
J7H1OuirSdZGUVv5qRL6uZJPb8ZndNcg3PrKvu/O63LmqRWfy3arml/2LgYu
ecbRUe1C8TAuA6wfAII8wHjRsnt8CYrkNn0lM2cPdo8f6S7H7o0NvGO4Erhy
RuFomMr6w4JXe1/LFZwG4F41zRqTHksnPW0T+AIpISR1cbpYxk6M+GG18ZgV
+MM+ISsknEXY046vg3pP7rT0c4WrI5R+PxwQvw/YSxeuoQ/7ZGuBA/MB15sw
GElUHeMHKakd2ZweCD714sNfDQO/ouM9wMm8hkVYsFnJB95+D9IhBJZCJ69I
oZ1MDuAoIGUwctWn00twTDxzZkPUVM3vr53J+Pl0qaH2jo5Mil0HqyzCWefY
MaMgZSwFkEHjLNvLcUk/i0e67/ynYEeNwdvFCRxtnqFg6ghXjrAvimkNLNFv
CbuCYfC20T5UfDRzCJBEErqPSaXSbNNF2l6SSxNkKCwBTeVgv4BIXMUCWLdp
tjZbWZILTEYelAiJi7QQyPm6XiOfZUB3MIh6Y/ztIU4jsZUUANgYCYuOWO0j
rmY3jWeibD7qGqs2na8ZwqKwH88uShzNBb46QKdgU4t3O0KbftaqVMqjocrl
fp54tdxD07KD426FXTSxSAzTcQeXaR54UE5qLxHFoCD5EKR241E10n3XomID
tWT5YY531QZNZxAKFW8/Xig0Qzw6+t7XwOTf+9V2xEiP5kEOJ4yjWSIx/1cy
CMVKLZYjlVr59PTacd3YFJ+KukZcP2auNH6HPIAh+fA+DTL9JtlzW/sXpJsf
XnNT2th9W4gEPZrDpRR+IxTD3sqRQDddjK+ISbd+8/9sW4JWot8YvBIP/sE7
F4w1z78pUoy8FED/mziUfNht52GFTEZRMdUCUxfh+1zBTz6/mYSFS5sBZQ6H
XbpZZOme6PFBz9R+2e8NYX4grnIGr9JT6eq64R4LqPmo+Q6CtEQHDSrC2uk5
aOPeEYFmCEpy+GpuZWlLD7703OQ5GxnCZug75dmyM2qv2S7apGV4OzdsLj6c
nQnLax3eBC/aXnc4+bRhy1IH960ZbBRo+dleEdVGmiEp79jzCHKdpiF5my5R
KgzqDaLjiydp6NK9CTI1qT2bDyiaYlz0aMsbaPfY+1iMtfUuEaMhb5kkjU0e
dvmIwSKpKtwBJoVdKkd/YULNTHWvIl2wpsjdZUJBbnTfHhUcTQQKuNwClY8d
fPZggRIS5UQYB13Re0FQy13xlbXHsj7BNmi9JNRhgRTtFdQUm0vexL2Wb0q+
M3/AfF60vtPqVGgh//vRONbjK2uIp1tmE1CSaokq2/0cOLqCn7IGKCFaSmra
bJ5Svj5v5/1zOIjnuWcIrQMxx0UFlVMJnxb+ELhvG8rJk4i2R7T/0r1KYpHL
NwFiqKSQ2h5RW6F8QaPidIBde48nxjHtwLZlMz1pOjFG42w4y8zkYAEVhg4L
tVT5x0bujWUivRCxovjppK7wrZ0DAj7psTPY1yCb0qPj52bERfOvxJzTWS0g
mfEOpvHSGQ5MtdBbk48Fa1tURhwQIH7taLd/msNhj8TsRbnTtaVpxHy5/hfv
yWHGkkN+enrIIdtjeeiDWSK8jNaWEUaQcXxvWpzl8KnnDPa3fe4ez4hXBTxX
ruEy/T++zTY4ln217fOxsJkvAjkLnZhjLR+5DHBBgjugom8vkTeXSd9QnM9R
PvvscveeofmcFBJsa8alzk4KTKZKaCOUx0EYJWYFsau9KxNwUENAN27bVIV/
A7m2W9cRUg7LDKO9DYpICrDahzg5v22lmDV/uSuWcNLd0zA9HYj4dnZ9BLN2
aDWb+CFF6m36HyJ8cQKQN+diaQ3b9nEomXGzrunJpWuHvWZ/9GHZBGnaEiWa
cdiSSlc3Pdfz0oOjdtpkEUGlw0wAWvN1Cdcw6QFDX3VTKDVRoSRhVCtSI0Gq
dVqVIXuUCJ4VvALO80OgqCuiD6cuOuEHaCNLaViVZZPVlTUF19TsVW6Sn962
Gygn4Hkv6e1z1eOxrOIhXtA3UMDy/hkLqNNoZHFRLcuPJv0dFZGcp7CTST+N
by7vMOOlQwhaNreOtz8Y+pZEXi4Za4VhXwq/hLxgqip2CxfP2o7GdRqJCbED
1wPqbOmPQliACf/pOI6Mo5U/GTHlOmqGBdbPhtNu64MrLECzNIQmbwGJLYEc
Xa3f/3WZnp6nN+eFhKGWquS6jZ63/5XqpWeSnEm0DXYwwc7/k7B6GAQ23alf
3AJ0ZCKc7gwmg8+fOdGAQ0QIMNxvN2DQVR1IJazLFD2IO+N7JpAjHwYOtQXw
6gsdT90ZPBKi2T8OjXZ9sQTAOhbnI+FsnrdqIrRSzoiFf9uPRmLFxXPtAawn
/6RGu4dMLCol20gHhh8jGrh4aNixdBIKr84uEcgp/ajq1+0EJXehuPDQmTqX
Z2VjcsWPnmcbje8F8y5VyJ06CQnEHUzjOrwVzcedFQ8N9FC/1akrLKzeMQDh
rwchibtP61574HN6lZdhNvsQQBmus8fu2fwjg3ln6cWN+ZZBAixiX7Ay1qtM
ehv84Urno9W1rwxeqnQ/qCeUYG+BOuLZ2kDQ2wNtl2CvRGHpi05d2C/dZn/F
lYzbZ7FJDX7sIuNjS9sn+eWfPOloYJuR8ICk/LdszH1DOX0txSJZfmRnr8IF
W9wfjlc4ScJEgVrxtp9eZ9bgrcY1+igxpNUsFoPD47aQCwV9liAJ4Ippdhus
4/A3j0VbWd/jpz1wIRHN5FZiHvvCXtT5vNDtl1P38xc5L/9nlqK6OznMl1KZ
kNHg8LgmG8psQfKd20n/id/KHZ6sJjph8TDoCp5y69d1FW3PxYiIBdWQYXZK
O1eowXf95hix97Np7vP7z5AwJS9e1tjZW63QcpMfOD8qWNPMX945vr+Z8FNj
lyt9ICj2pGZ4KIdTjr7jVK7JUm6MsdSTyEoX3dLWlKZmv+1VuUKquvyJo8+f
0DniCDGqA3oLPuyFKJm9jH4q/1XmKZ1ul5VFddsn4YpecM9jCTiEzOT6Oamk
6ygOecK0F2xJ43kv7fGsO2/z62UiOOWT42+WF4cifrbv/3ZAYBfj2OT5TGDF
dFhe9DCiQ6sR4PPS5BA5TnxtnsYm5RuEIoHn4xa9uNTQCRDET6c8rF9HXbwA
G3iLRRQ+bd74IBjp4eokLDZTOnW/UZi/X8bHi+GmyL4OtahLCQBhu1eJHF+K
jtnyzK1St5kjSpUBFQsujkl47P7hf87m+DMU6YS7q0Ouc8AksMQiJzuYJF9o
EKoJoIyFEgTbkArvjAM6yGhvH6rMLtIf20nE1zl7BtYBMK56+5+oNYDr5RnJ
AD/q4T8ft82/1QPPVgs8/ip/OCQmy/HsAedy5z5TEF0ynXGCgFebu5raDT5C
GPkZyNi5EYEIHX3urHgLsuIWIb/vHen6EhzZ1ZIqm0HijKL9GRmAaccoEdd1
aP5pV1dJSi9ho4dIqBkpKNnPGWLA01/anOQmqN/rmN35dlAeIPCWWUt7mGrF
NGX5N4p3KcX7/Pnh+WLftnoreWRElyYoM+oYBTxNLgE/WgwIm6LU4AyhW4jN
zx2lGcU63iUrk8AO2NVN4X2ytQm7gE4Ygbk9sgK9Ifg4CYdkfofZ23ef/Tj8
kvBwWwjcI0MfB4oI4kq7wU+kkXUsu5/KUIGRW7qdzuRrYUDsnpo86oiZLfGZ
JuI1C4StxmLa/Dx29uQ8dtHFw6E0tELg63Jbb9rJq+j96PeEUR7K7ijGA2A3
rbNh4cPnebRhE0bhhdxlcRMio7j6RvMxhHGzqr0uwkI7J3ns7XkfducE8MuS
gp8rR1ClItc8U2JPNgHFP5ofuL6Hfujpb0zzKBOs+cmizgKAUBQUBnm7A/EP
DyolaFFFVN2Bx8l+dBXg6IJQMkr8IAiOlem13KZ6GVyUQIgYibHflhUKSFr0
WzCyIQadcUS8AMAK/6pyJHyrxc0TOuhrp5b+4ov5QPtRAz8IDZle6g4QzhB/
kQ4t/f/umAaBbGidvnegYjmr1Q64MNpkHJGiYwXPps+8X7PokEMKpWlgyjlm
gO9SS6bJNfBJfWvEfmBjnYoG0PBrc798gcmcvBzLJSH0IAwAIG0ZxQLaWkAZ
d+lWga14lXLXie/S82/mDpakawt7aDkEkvKyzmfNlzhmOp36v00mF6AhopdZ
VrtXyahrQu/FlS0rL8+tR8PAYQuoPjsKE1gTRihp6hpv3p716EpifKcCju1I
XFtxmFUNC10bBDEqD0hykx9IGLxQ4aunp/JcvdS6VRInSZ3SEk7SuBrKSARL
kuuOGbiKidismAFr1Spe93P6YPLN/OEFLRwiGfCizgrw/XofP8i3JGXWaKqu
bgP+qoUA3Ebj+sxfDowmTD/4888KQmFZddv0WAkkMrXguA1kXr3Kwd68pK+U
mHPp2ArJGE/Kv7OPIZJdLytusyse4WXCjTdP1WP5sByR5kn3AIhV7WBtXk4B
4sIzcu1Wc+UaVO7hyEH0uwLso+VsjswLhj9wBNz/NGT99IXBXXuyoH7ZRtAc
UlqmpY+26n8WRhHPSabg4oGR8dZnMvBFOnO3lhx67mYhYJA8Gy9ri+np/NNf
EBvSdkV8vA38R0HmLDuFh9uuPYu75n4ON0nJqU8rkuEv3vrb+ysYQaP+Uoqd
rks6yaCUROyM4U+VEx0xhCbBuvaww9v1ItU9kiAtZBpCkWcZGcGcQnqceaqg
tqCJ6fPGtHJOms7VhC1Y6G13hD5fzPIfLFUHYz4LPshyto497t/aIdLeZhpd
J6uNm976VyNvPadIR2chfV8YY49PkjKJHSBuul7Zge8W5qy0bJciTiUErL9g
3/czyCErDzE3PEq7lGkM5CvlcRetsQVUrW0HgruJwTrv8eUcEnqRZmz0HSjJ
05K2WK2kkMW/jESyezL1AW5IJxN8SF3/tb6kDql99ERy/kpSaIO3vegnPp0H
st32FCb7VCvOsJjZikiAIZPyYA78eJn+1/xi2YR2Vh1bnLuarXCQfr/8mCbU
Q1tIof5OEw/rtUv1ZRil68DLmY7z7z30nGyKbG0VLKXPzPOodHpRbuSJGeSX
A7tyFWN2m91vQGIvM9T2VVli7acXL4GmsvFDFZbvBzC893q78NAF2tfoSuO4
VMuCpXEPc4gRsqM6w7AytR0c2a/YieYqqJB3fGMS2KxCKif5Ur383bVT5jVf
bfM/xK5UnYZbKQtmInaAPgEDCx5V30rhC9RnpCh3AjTprB7wFrXtq53WXgxx
k06AZf67oCChfp0oLjDYmg7REQ0WiPVJGo+NN3Pq3L2oYvUKzdFq4pa4el8f
Mpn25/i4rLJwGO4PfQhCpjBbKrJ/qodw0bY4QFVRTn0fGsBopLGF5Byr0OIn
JDIXGZ7dKJvlZOn3QMl3yeFSmc8FIC5/+kfXOYv4ZJxi21L1mf4rEbvXebyF
jAADf40ZEeejGIIPYP8Ay0ehWuqndbqTR8H0iNDkewZhQYlKfJcE1yCmo40E
jo3aDwFlhtt6SEBRP7Pi8XmrwnuXnxea5GU9OkpDataWBEdfrb4iWW3uN37G
6yC1ZlPQxWmKlylpb+Pjxon439BIs2ViLJcH6ddA/xU5zeV2M2rb9Ls+f+aA
9q4R4yX4obCYkCP6T/uQ+I58TgwDPh8tjvzC9uoVtKJcKJr4s8E1JN8y9uFG
wo3SFP/NRfRO3URGxa0V1TaZOsgN9yViGH0/iUy0AFBqhL2wb2VpaIwzIxgs
0gKFeDv0TMO27oLjo4g6Y42tMfEbHzWHHUkrXpuy0qM557vxEgLssKA4pNhJ
hpnSoGPns5PCQc1mfncajqmwHZkudhjFiwnixo95vSaB1qMwZtCoe2o4DB2+
kdWbqcDR/lrTsMeRNvtY/EiWKrGL3qTQP/joLm4kK12ZSOHVHPdgGEnC+R4d
KOrCgPAp6Ea8Mb+Llpd2p9WCMqAHnQI0OgJnntiFS7TQzQlVfiw+qIfDG3vR
I4z4P2oTCZNOWW4VTsUNppV3r+ikQTy4rh1xc2TYTMNPvwGF2WPCRwpHhSis
kwQCrPoLz+bqmkNfROPwi+aezg5pXQ/eqSO9/vkWuAZggnP9+LEqGcBgj54z
4Sni8koFl933FHQ+NxLPYM0+LQz9Zd2wfPXFDGuK4XgPhqr9ScdAbops83gF
IR/ZxXb4P5c0LCzi+ySup+HML5jDAB5MYoHWIbtfEYY9b8jhWHgqov+38nec
jS5kpO0fTcof6lAmTmuDs66Fw05uGmtN54punbqjCR7K1xdz8DguMBEZF6Mc
kyNkYRMf/5kUninltZErCOTgsi2p6ndwVHQfmXkFQYTqQ5YSQiy7ZjzXPkYw
GzC3cHXUAkNCX7tlAKQMV+CEzt50brhxcJWEM3YY3b0OJx1sxPVf26AAo01g
blxaYBijjtC0W6APyMlMbw22iKkXS4iX9GFsD8mf6u6NDvdFwkH6VpxBzvHn
IMQcBjcM6vAV+pjORP2NpgkHNuTEgh5DA+ue6BKrofR0/qggBvZAkLjPnaEz
+tj/6AjlQXcYqJGwVx7o/lzRG2lus93gfFRdRg1OMY2BnzheYWZtnyyAkFco
jSN634JoFq0dwGsadYICWw6WO3887PMZe+8PNoSskqPiibtlrZ6qwr7Y3bHv
pF/QsaAPu60wG8qh+RczC4vfEJHLD3Lx/B8eSGnhiqgTa80BcCVquddROG5h
9eeiFn3DvtVgdOBALR8awD6rv+LoSeGvkOIBqCGOnBCPFvrYBpBVXArJjnpA
McMPytI4w+Ys4YYhPcxqtq9RMYasNOpgFY9/ZDfzoitQuYzbE4JBk2bqSrar
9/5tmOJ+qiZYl9yYLT+2/hAi/nuuEuRrdzw2eoMnkfb+a/GMYftuUq3jVHM6
TXH3Hp5Zr2o/0LqvnTH6xJ9nOZto2Yv7hfi4oEYZ70WvsV0+O7A6AfWpBMmO
rkWyU6G7rUWqTHBucv8esW+g0UuppQmy9/7R9GHLttdE74SubzAuVLqBNN2n
d6AxUdjd/15HbQHi5yMjEfMSa2JDOhxfLxRglegLM3/0opR42O9Fli6lgCXj
WuEFFMpbrX7W5vNjdBzMm6c3L9BBJm1TlFgS7APeEXNQ4Qlvd6JxPLoytopO
gm1GR/xEQ8YsPgsKRGRGKAu5i59t3etKQiuclrv1/XJIdo4h6oasRkuyHt3v
/3TbaJybg6EZKUeDijtFthwcmv4hZvwZ2xKKDIi+ieVQHInCH2vSKkB79lfp
3hdNNGFqQTn3VmUX8hiWd7K8RA/X7zUL9RPcpXvWVGAYZTz1tW0Ba3yx0RNs
HqRJYQ0pQJp0QoZI3ci7AxG6SiaupUoN81CnCtRUbQputoCwReKrJT7qJzv3
XOx86XftJe2wYfzSwxOkZ0F/Q5ngTUKfO68lc77gUXbIppac1r+8hF/c17eA
d6kDRUPN4frGEU0Zxu6Eo1eaOw4fRUKOKP6NRhzIctC/G9Hi6d08DaXlYcxM
VfgNTYpjnUZWzlePv/xnAkzOMbS6qBoU3CVL5AfutCAyXrBs+VAhRBmzG3L3
wtnNhN5ZEtWy2isapZ5RtQ4bnzwVhg6M0vHn7HJr2GyxPRtUmOty/WX4Hky8
/89qvt5os2NTTS9ZeMRF32jj4Omp9hM0t8/rQcwf5lhRJbjIVaks7V7q2jZW
YSs/QrLV9cQYELvGMsqCHfAem0muc9nnFtWnffnYl2w3xy/1wC3+rsQ2M9Bj
9twNfZNRdOYnATQRIae1C7EDUoHBW2QxPztxvgjHPP6zddCIMFS2MRxw16VK
3HxR+dvaG8Hx1XtnZbZp2ZUR9v/Ht+hzCRB0apyofjo1c/JPaPTvmPr4HBIn
w95eJoo3zbi1uLpPmvnOylV0qHer33t+0RHDvrV7m4glvd8HZzpHODTzWEYy
oDZrN8026jm79LKhAXJWgHZnw3mgfwmyM9hlH/ZB7rQ+Xl5CJkDhyxkV0pJJ
ICO65uPlSjwxcyXwdLvtq1dJajwSnlm/g29IMd+0GquNTTDk2U1BMXVERVko
MHLJ77Bc6Dc249l5G2FwoBSbzOZwMBBiVyVWEpAdfHHUCsaW8XtdizHeA2Jb
HKD6YYM7fNBE5Y1p6fk6X8h0e8+BDmugF8SKD6krRMDo4PsBjjlzUwg9OS1v
AHXoPpqAsqkh8sX//njWnkBv5RBaSFGoyRUM1JZn5CQEj4lS5dL/NkPU4rKm
CsIREN7r8FBKt8oh/0ippM3Q9lOcZyS3qZet2qJDOs/uE0Xq1et5kzLNV5Bu
b4K7u4qmtcYtZeFuH47flu3LdDVUr2sx56bytfs9vRtxrxnbT7ROS0pD5kv/
8e2GW127w1uaOyJ7LbOapHx4b4oop0bqNSeuKUg/R4P6QJNiXDDTOyOqKXe5
+jAuikAcs2y5kcMBcsI+GZdwCO1Xz9dw8fKyanuo1eyt3EmXn3XDlYF5+g4j
0bbbAZrmOw/hDhPRw+FJJWUCogMtyC6i2ATVCxnGZh40LOlag6CvZEJsloOt
3CBCABY6kLos0gF2WJsWp5y42btEyzqVq2FGt3ePCN/a8l+fRWUoYlwh9ZDB
aRNRQfyofnYti7JePDgZAskFoFyBTwILR/Syz2qRHfdLARZhyV5ihhKn6fYU
07EEYtxN1rOmB0Hju1B7EbxMRCXKcjSmJ8QnOJ3YUauVBYbCSxnRECKUW09F
+IRuVABJ2ashWJKln9JqhtUKQWNIZfDqtGvLjnP3nbl4mtOOI9xKS8c19/TK
YlWZ6p/n6DTsts0fChwegHeV7j/fKEOqfAtTAsLQEQbzWtRzOZPW1+GYaYak
8ZH8VHgrj+Fw50vedmBW/kPfXvPQEa3sRF6joo8wokRzcV5d7H9fRZGexu4I
vBgpWo3XxnkJdvxdTlBWvfF9v/FyyNBe5pED1IbWHNMuImAxY1AgH/NhO1Wx
k7IC31lj2AvIidUVVLhIbM2JTGOP5C8DfbonjFr1A98+CxMJnVoCHXqeStdn
gqDiQTY/bKRWJbjd4cEAFRFeYOIyI0wRMoGLh43Acjd/h4JKQCvDSTnuwZIv
9/G52NAlqOzi+lbTc+0enroD56SlPzK+AJh9ZdrD9PSro7eehKY4lwpJd6Li
V9rV7PMobuBj7Guh+vne0+qCCkVJItXz7kE+8jiRqqQbzyR0zd73M7J6ty7P
hUHbiDVP3xFboHp7GA9nmISJc1d5b9Ol2/gzj4pCoyzSpq82HP7/P7x4TQnw
Q/zudm53vMQ8OsOdb7bpVVBln8clxvIOyMR+v+KtJIc2oQwDQT77P3XCwOpo
XBYpoPBBGZGZ2c6oX7/QzoP/CW3e5Iy6J81PS1ApBtlyK7+xV6PnuDSeo4rr
v7xRLtvCI0VGyeII3ymk1AGULJVY2UFT2dQB7lM/vz1qCfh76ewP2Gmc16QG
1oPv8SnoqrWeuXIwlshlvIVkvwdsYAh1jm2G4NU6KN+uzfwPTTyfbOWm32zc
ZrTuICceeXcaP/iWncjNRcAHBJNqDjsWiKqLs67OLJCeoGTKoy0h+CRzeEkj
q/qXHgFg1MRO7dCJbUCYPN25RX/TK4UURYExh+vkgtsTL3cXD9rPf8WoT4pC
E1d/GYwFKxLpd+wnzflK62Ug3TV9XYasbUxRro5QVkRxT5zBpXdlHmiHs8BG
hhjgTF46ZfxuqNoRXt8Ktgn6HT5kG2mL2JC/aOF6jRAOeFYFroCAhdcIrncJ
l+T9KKC4W2GuYnggjdJ8aFt1l78sC1VHeWGm47zOJPLo8+x4zi4qp/vVJlrY
eVtxwETZgYdfjGxd9eYnGIQYRd7TKCxoZdvRMvFShNpYHv75Cmk2W2rxkZQY
Wz5qzH50DNA/U7yeDsM1x5p4oemDOapFJscdYZ2TdhE6w3s0+z8gsE68c/+a
MOXHZ5uiXmpA2KpXkyOBkF5jlZwhhtI/BVp9Y6rbe3Ql6mIWWhq6kAm+ahJl
NtDBLaxUULD5+JJe2vVHXSWLLimy8gQIj0GNxiu8vBYp3uy1aa3Ko4Vbaot3
nHleNZ5yHU9Ag9R8m0+R+47rwO0GdH9stHf7BHgHMyrpGY8yZTqvNoYSJ55K
05W850e5ggBc1p/G0FuOt6Ei1FYicy9esfUoGwL4ZZuF5OELO82lMtOjqaMQ
kbb7ezFNp8K5biVTjYst/AfOEDeY+Tbi+0nS3tTng1Gyk0sDFh9v2WzzkclT
Y5A09ok61uOSC/0snHvH7AdN4Njies3D58mkR6BsiGforZXy8KZaDRWmHE9I
I8fdZUL2xyZQ25RuLUCCsMPNOzCAGi4HS6glp/uEoSLF1V+2SH9Voe1Cpkzx
Sct1+HW9HeOkTkcRzzRToTi4jCHe8sv/3o5io/7V4IKCcNS1vMQOpnpTg7ec
c/QPWGbIryCNQ/KEgFAhee6vi+LdjSN7OLd0d0EzbCJ9oSNjjqE6ApMQRdMl
M03RzudyzfUmEn/5NGEDDPi9jVJBX7CHUcGTVmFItzTacOwh4C+3f13dGFHH
85KL7l5oA/mb92oJ8kGMD2WajWrzCcsPTsEof/p/9eIZ4qtZExmzx7IwWN2n
KM6493n2w5/QRtV/rVFEhY6E1aewp1rwP8nRdFq7bU27eI1O5QHFpX3TBzuJ
ERsVNkenKAMzvS2aHK+iPxrauwfxCB2WD/QJMaBidJ1embg1EuKSJQy5nxwj
rXKxMf9MWDLfBwTNaQbatCz/kjxeHuS1GPWk/eRZITv8tCChMrSlfycnwkS1
Y13JlrJj8rwhKWgUC2TlXSiWsSCCJwmEiHfja1iFrD4N4oEiTV6JqUUnnWIW
PZXbfM0XQ1nlJbmunSHQc7DprthGbi5S+naaKeEsr6uLZcfcsu8r4zj2v+90
PoSEsJ2e6QftgHW9rLRwHYr97WMEZVmy1sIujvRZofJPfhlrEkXfTwHEhZZ2
HR4p+2XwsT5G8qkkAk+I5Q14OXKUsbCrSjP3TcywyHpij+4v6wMp1TWLKWpO
bXPWwbc3e7wEaSbvkuVw0/FCFQUNhBe0JXklBcuTLT36SVWrA1vui+xSFlSM
uTwbjbFXfqzAU6yZoG7qTuUD+dhIgBNZZ16k5oO3/GxRcsMzpXcEnygAafSg
mjiDD0JdzFwfmrlVsHlBLFA7wnvJlnBephLMoBXchZLS5IW6GKicwl+Srxkd
u5NPU+6iAHElr0uBZYmI7nFZE9mfEGqZgsdpgRk6MzHslN+iZeSfpgmA5vad
uDtjUKUSJ5tUxiGeVtxRSTW8oRMp2jDgw8MMnXQrWrCbQWKdJVmLSoGWnnoh
3DNHFvAn4qEdluWpmbSckARDzkd7m6kxnf4Jxw0xw60xXn6dECTTvjcWs+lv
w6TqpVIKUEJk8aI25z8ZpwErnaElOaHKgTddp0Y5geuPoRO6VV529rkSQXHQ
Ut+LrZNc2lsIlzkwxJ6r5Qbq0aBhnC38jADYQCfY2VII/4ka6pWF1H997Mu0
NJPBbFpgf6LMxk1NkaEMJStgZzVAXNj4QWojYQ8MjMJztfaFddWgdQqq8jN7
O3t5nPuQIB60EcKSZAoBKcX954h6NmTu4VvPF9nxW3F3OgVbspxOUqkq+egg
cdEw4+T+v/SVL9ibOlFdEQK+WT/ZtBDkyTTVAta0uZ2+KJSYAvzGoP7gp6O5
a8Hjtk8ypY3EQ1opxt8SQxKDN/a/O6m86Xev6vCOMCCytlm2FvUpt046Wulj
nmRsMuUKJ9+mRY2UjhX9E/stj29zE7f2gfM2Mt7TyouhSnK3e/Hx1KcCw10X
9aqXHBi9xIqLYy6HjfjJxEUHQTa5oR2bDqIupLaK/XZLKpB9Zku86bokG+Du
CahzYcUelaE1A/rM1ghIg1uT9Z7776YTt+9jz9jpXdd6hlJoip3bFIzixd/k
EeS4YE0UrLuTugGIDD3dPfcnrkcDSt7YOm9swbyyks46ZWBRKJPpKOYX5rPs
WHFzpySdp1rYwQTtGrudm+/W+e6N+AlQBW6ase9kvkgQVDi6t+FNBY/czwxe
MyVaR9MM87kqrKvN0/rU1vluJ5uJG6tGg5qQKLUBJ0eOfavRaaiiKNZJS+90
Iz9kg0PfRSoPQ9BmG4MCQMkklIdqijrJL16nn62XmQhBLuS7mh7yQFPTsPso
lEKQD2Kq2KqFtGGRkOriprQ2Nj+YbRcGQ/wyBLqnznM8fyPa6/RZYUZ25JmR
7lxfhAez7SpULviIT2D25Fd0Sr6PNzP9eRTM3ueT77renh1FMC+4ZYtoBNw6
YGMWVrVt6lwMoSn4JywUjO5pSLSy4YbhE0rUsVGRMqPL+vLg7O8K6sGDQcWY
bILtBdKaERxe1irRSh/23MohCGL0yikE+QBLYtMltE9R5wMGFGGy3LrUgbXy
FqvA5iIQeW9uPQecpSd1v5hEIJP1dZcdewZD/9bG7oej+OatYKSXq3SEAM2S
MOB55HS1ymnP6328+DRQ9bU+AgIv3/ClFQR1en3oY96g90BPphKL/mNE/0CC
GPB2xJr9nDXetY5M8UfO9WxUd1J4ioqVpdaOlIebQIx9YRW46pe4k13a6etF
vP8xvCHMrLovw4bPKocMWrJmxfJI6RY9Jrjm44jwalkcM7Mu5dPuaMW+DZbc
SXA+XbzHbBNMS7wadzI89oFp6jpVxsw3R2HToux1TxH1I9vaslPMBfe6tHtT
AFWmuLvqEZkGkLeJ9tHCKSDE8FedEDdml4SgYyeK4Sa8bRN47nQmc9KhpyGH
iwE398HL6sfLZdZilDuWdROV2mHX4gkgjVr5gCjD/K4hFG9owQseHE4uwhvX
r8rKcN08tbCD2ayE3dZRbqEgEj+BoMEIue/JGa/0G/sx/l50hreQirLsdu6k
3prWQinuozd3dokkD9oFs8tQy6KQyZoRfcAvwtXj88XBLNVkmHzQNvX3spVV
jDKDyW/TFkNu4YhCVRMbR56pYhdOdVFFxeU/mRTGgIrnnfHBR56vH5+ULDdw
q7GOyTLaBLks4VW4WQB9RqsfTR7urYFCL5O02DUX+JnelwolSwPyCpp5beGg
Ndyl60m4DTHaVpDJbfSrc3mTFOJE8RYIIPKsthrlvnGyePT8rt1nqvSOy+o+
a7NC81BBPNnH4JrYdapx5v76ldha5o5cIGOCzC1ipMvyizT/ZAGJz4iaATWe
YwFPH7QfNIBo8GdLawuyAxuUqqdXAKf/be5VlYm+clqiFt0whyV7EAmihgNF
mHEeiNURPSjf+UkuAHuGmtN98y0ISCod6VXKXbqyocuH/DtuxfwLFEIOZ6UU
4FHIdekrSobose/wS9RHaqvOQuNSIH2lehb/90d0oNQRovcGlMQQ/wMBPP6f
KnlUVZzZUMhxk+BIpeIcNUyFQkj3gfMxe7wXLwcZwKLgeZYviCdMpATbHIJa
R0GWEBivyDEUx4kdVhm7lXHgbji0t7qkMzhZWVVGtl0aIztRRrJXnwCsTete
JwSigNrxNynudDfBO1zWZAL/VnjfImXHWKmynD/pbPjhYwu/xbtg4gJrtSnv
peGj5xhfkUSru45h+VOB/mOMZp7i7XplD/nMiUnqGiXf26jv7jC5wByxVQcc
py2udBmCi04cvt/jI1xLsl4Fyc1eQQfLX2Ym05TwgYOB8G4Y//mfJkSb0tAF
nGEPwd02JyVar6rGdwX6TCOBmocXYRQb2xlxSGI+EpvTWmcuQt5j8vd/qGD0
CIfI/UGZUg4zc9ynts/qAE9M/VrvPN0DrEBzLBE3wVcTWe01Nb89t/cwVJRl
ziFDJGE4IEmLn04KepBlPeMN7fVpP4b7+BYxUBJdBcgMWy1HUSLKxBza9xlI
e116Vo6wNo7vWYU5M6JbNwRlGoNSPQghEXR4xbknKnPQcmw588gE42pi6AZr
2nfP5gLEgbEy+HBZSGbEwomSrXLazg7kFeJLBVSETgpzK1QdCmQIBuBJ2jOZ
T6VdIbAWpx3NCsAakQAWzOQRvRgA7HpTOscPvsqbpkTyFm5Ab8IBa1NL1jxx
cxIZ+8893jfLkZU8X+/OW2QS5F/7nSFeq08bN576cjN8s/UeDLGF74UICu0r
znjEGdLyRjk2otWLrfxZLaVwBFzK0dQmlHC2KcgBTpQ8o1wtTQSNSdRNJfWG
LZEEF+9rYqoitRdBS8wIc6cMvMf0+TBl719WsEtH1wRVB+c70zuqTzxSFl6F
OING9+Oo998cSPNINm66tAfaGGVuRwc0dFEWA89l40bzy+XvcgCWxqhHr+Yw
8rXIoB+NJleAHJvVQNFafOKPhjtgFVaPk0YmDZNy4KlYoRKn2jZQUslm54Q3
DHMXYNJ9PAvUWi6nK0ZqPuga0IkfNADpvy7iY7ddrcGHia9RApd2KHOTxTqu
9IXzZvqgxSGMqQVTua0w+d2tAfIXXBjjWytrZlnw/pgJm1qPQ/7r7iFUv1Pc
zx7kLhqa8FJ5+lBxX2f/7zKnYzZ46CJqZ7+vqJxr/tbuEbArVlSs75gtGZE7
cOibj2Jd0pCQ309yMQguzE/w/ijgO5R6MDvKIFU/UaoL+bcGuW9L/z703lVB
ndboICVr1gDI9JXpRHdGCbcZasm5v0E92oUvfRYigHYAbl7L+F587zTAnatw
fejxkbo4nh0gqtM46zyJMBVFwJdXYRCAyAKYRN5BAzVb3u6jbBfBqik+vI1/
be/9L2idJwkRxwfpYEkCqJ09ykNAMAE2qrKbtvIm3txEtpSzsTMv+x96n6J3
5PrmHTBrTv8dIk4iYVpdeyyQuWbVA3lf72rqrjWlTaWVUJ0iXPoSpxpNK/sk
bKYybtMSqG54DnkmlsQvZ0TvzrWwnaq0YJNMUJcVZJVG33F4NymmHGJbi60d
K+GQFb7BwD9msUydDqYLQaU6l7ZmTPoggBWrfpV2kPVVmfrOXnNO0HRWZZB5
TcpZp6wNc+50wCJhZm5mJkLGtwJ9BCgw9S/ANYDKa1pKIDZLQd4COsNNAMsM
1qDwzhSFkbUs/v6e1cvnXNqFB6mGCKJiKSqkEa8/l6YXQEJkG7K725KjnsnE
NNm6FlTK+JsW2afZSMNj4ZNuiFpV1AXDuEgsEpDLF5cHjfyJKo47Dpl5onEw
XjTQOm/kvdyt00B0co5MJ6bQ0iXINLB0B6Fax+0SdSP8S/VQLt1R+5JtYk5e
4CR8hF+vq56Hq19Jkid54/QBVaiorBpwYOQktWVppqs7fIBTCIHpIouFZzIz
bfhwKmmPrlxX6z6UQV+68sCq8Y8PVNqU6skjWu3pqp9sgs9nuTgD6Ptl7pgO
Mky/bsA73zqLCHrTFM7OiMHPged+r9r7IxOq6UPXl0wfeeLcL3b/GZICnQTL
TxiutkLaDB5hTf2rtWmE3Sh8BmFNS+IMSMGjBJIos8/s1iHfXlLZWUmD8aqX
25Kh67sBUYVl924ssz+8dr/DMSxyQjj8hYAcKJUcR+WBG54JdYjTH23hZbfp
rr7AM3OM/9fQ+qdv1qEPP2udZk+AO3lIZlAJhLWdrkcc7S56Z38BZV++1bxm
Zrxy+kptA67IlW30COtLF6+I8aKqO5Cxyq9d/V/yH0I3jkKpROop6zVqU+wf
jFzcl6qJfacCrt5KLf/fByeD5oCjuv9X0XxtLiRdULeOYpsD7bX7Iar3aRLZ
Hpla4qT4z7kFZX0Jd/GU1RLeX2twbYitHp2WSwZIogUZsB3TDk+8kVteJ7/2
ELCwQ8pkRhDcHxlwpauAKne5TV5LG+WYcnm/UVO8q1+r3z965laVmZhVaSuI
yoUTM1h+rmjWRpdLsYNVnTDvWurW8dVP0rCoImvLFWG6OvRT4yXbZkjwUfT9
E619xXnjKyCkrwVPzNA5p59gBrrxKwye4IEzbK73NylWRqiWYORVRHMyV5sD
tvzGmHjgwtPR1yRMD+RTAyAsclTCTD3h2yHYzexKvTacvVE/8UwilrvZ4Sq4
n9FXRV3NGdrRM5lrp5pnQMNUgn9t2gA5iZ61thSKGA1gBV02GLQQ5gCkbwy4
ymVs5hy3NvT1t8AzQ/vGDeOHN9Y5+ynwabvYDDOrC1I6IPTkmi2EmntZ7xYu
3v032bVOIr1UNJ+JkGv7+CfkMBPJ/JQCmVfNqIIU1prBzeijRjBcIxs81fi8
mjOgniDQb6TH2Wg89DdzdNKI6OEu+o6UwgdtW/dBn1V/1gHGgNDdudVh4O3B
3L3qzxR7ttYeKMWKfJd8gSJu4SqTpjhl+vMBH+f6wo7WQzMyWTskH6Nb09CC
TBjHkb46PCBHGjLuYH2pvlY/p3DzcfUtB4Ne81QhGmOHkVMwguEStILX6Sew
UVWpvDHgUuDzul9R4qeJldZ98L8Wd7BNxh1dfH2oQ3gzbqmlA+v8r0g0AYoa
3hTHYQbwEOqdhTMQZrne0qS7woQ/VyAIzVFDN0B5XCVEBRDEheXoSMmkf/Wu
CARFyOlbACdcJ9i70sgVNucFMHYUwB0zkfryIJ4/hVs34HEkJF3pqvpf8maL
0aBdWhM/xYzkrvDoPgjJYU1NuRfPGCB3fQXcaPyVVk+kRYTtQrqYokZaqZTb
dmEezGekWCEOi6acBNuhkHV5OOw2QRFBUJEslymO95SazWd2Sn0X6P9IJ0+f
TX5YvvHbzSXi5iW4cOjMs3Q4dNOiJCUtvecAdPMPNxnvot16HGACdukIf5ah
fFbXpMsKhTXSD9uKJENDFX/HmQMk7Ia27bq8bcfDjeVZUoAtBYmuKUL0XHSZ
zk5Wj9bHGuOIVO6Wuv15/D3QAcUSHiVfOwJQNsSIua/M9HWzZaBq9Scb6Ry/
kMMwMr+QdUH3rboqpNRlma6nr4aHVyeoV0+FFm5mYpb8GdtEgyIqPMRhAZx7
YTjc8fCTDf0YLzkgA+ssH718MBKDwnb21E/bfEQXeKl9NZXDfzLSqRIwjaMv
zOUTZaLpHc932ZFzkb1gkOZUBJbA2nthgjA9Z2eum9wC5PxAES9E/bSNUhX7
zwn8ZqkwFynKGZbvV9w6pQgozg6VDNThdiHNNSLn3gfx1+7XCeifB7apFsvt
FlVtQcyXRNrsmvLmG0+MNgWmA4ciez/oveOtr3KEqrcGfJVrpvPPDzaD8idf
qv5fwER91vzhkEqzjaE1Ce1cl6tKi09Ucqmj7mUgp+Mj73rhzwNVhB98SVJ3
VrJKwTEgjL+PZUHP21JzbWeMW8JrdqzAl+8VkpE+hncyWB234q6X3jIp22Ds
EKa63qgDp0VLIH/0RXWqXI+7WywAMhFDm7M8nO2PA/qEk6jrKk8TGpa+BQ0n
JvIRnZ53w4mD2YNThnZbCr+ZFo1NxFHdVJUY4H8FsE5imTfpcTa4CoP5m9nT
RkQY4q0kRvgkfELjFQZFwOMOEdeA+9wfY9cOjaYi42wPZY07lkUn6/5OQeIE
1YMvv7LOmIIrpUh9DcPzjG3pN281DFb3UNrii0SWkQ65fsLUN/dMcK5BOdn0
YBJ0k14lnhoTdhBhmlSoT+rtPbWdCOoWWViJtY4+PKA8R6k92JhO/gQ6v8cP
zjwp+NAveohpYqxm/yC0bek9MmP59OK/3Nb8p75r0NBUSUbMF++s5Lidzcn3
x0wJuzMMH75vSCVQFzuXaEVDi+zPmhqMrn8GEWGSUswQpCSQDzTJ56VkNdIn
mDwEfLMIqhAjN1qDTl2A0s0SZWXOEUNEmh/4EeRUNVsQr+kq91kxFcub09qo
rkut0J2Iv/VghtI6TEbTYtBuTL4V/jVJxhCzJHcHfcOEVNvtl7yrTBmXdUSv
3av3PrUaUFtXQMOZBa+WEwV1DB8vWEf4vH52JN2NnuHPu045ExUIHNvhDpf4
WOKPT8tXe5O4zGsqYmC6c5IWNnGi9j2V8wRGdooGEd+0+IPTue6Jdplv5Izv
4iYXDpQmVqM8ggQkLeJciSJl9jAHKnyG+AwkXuQz2gyPpkItT3K9iqJjBkml
k15IMvPYmyOKtfBqagNZUV9/6wlZjSPa42y7rd5BioxCJhvu6Mvn4FbH14fy
BluIw4tupLEKIMfmWRyJJJpLGnULHrPTfrPDGnrI0E0bzuD0wgcAy2EO1sIQ
iHPKbTXHWAdGeME+xGrobDZhFM486v3x1AR29vINS6ns/p+V8DZ8OvfhizkI
XChY34TGyirvZsdD5YBA/NEbzZLxRPB1cGPI7Jsn9jSMnvSqu0KuYbsEFqhL
m5REEjyK1k2zyIVw5+ZJCu9vBBNY41jt2wr/KvSXhhUg9s4Y0vRsQ6HGL1hs
z+pF2Jq08+m1KL0tvuL3Co57VJHr+1Zvu5ZS2e94dvWwZBXrJR8mXZ5gijE0
yVMHFeBF3roBQWKzyO7gghadYSjsOrO8zFH2LEATecpX08QKirRJ6wi3M903
Vm0aeoHnOYYzbteSPYF5HNKKWaM2OELan282+Bae+OSnLEQ3wpxzsivBGfox
9is7D0ttpokqSdeNzoiESGM8C+BhcozZZ7r66OJeyo56GUUTVm13EMgvYgb8
Zp2mm/TBsaKvkbNr5arfTeMxSOLDqyJRSuLUTARQdzeAmxjCckWRzPkzltWc
LVwyih/cCf13jd/SGh+4sz0GEFxArvyFWbh8IZQagcV0JEYddVKbZUvJVTkq
ACCRoby8ovB01ilj7fzc2lATl0YmEvUcD452X9qbyk2wH00jtmStt9DRKe9f
hTsSpPuU4kAfHylpSxo8ZS1NoU8Y9bYEEDumyEZsh9/0Y5S7ba0e4pcQbfO4
LnGoJvF4g/K87U1y8J7kR74MOmI088QMyihveK137l+xAb2qg9mPEclOVrzd
9Gm83m1rMuhvzGTrxsNgs0Drvvimiw/G5i+PoyvRmlYgbnaFgaN+zN68+UfW
iuPePSUXFBok8KIVkB2mZdCQ0m42ZCbl0qsIQ1NnsMwvXWTMMF6NEfZ1eh1e
jTOJFZHJMt96/+4xroeLgk9ttBUqZ7jPpwiowUsQgSnEdyaCxBD9sAgn+XpP
F1FRu4pGvoDykH8dAXyCntbhJDfpg5TFxXof/YvWlSYPWnc8WggOBPzCjY+r
0qrmeghEacPFf/UzIbjL4G8lOLC3ztnNyJe/m0kIXyf/zSdCcFa4p5AsX7Xu
MyZdlGjgr/rZ6t3H5767pSremM8rBHAi09v/5K2WJQ7z7nQcDvzu1W+U09+l
QdVT+8/0crXgcD/dv1N01udiXuRXWyHVPF5mnyb6lTVY5a+kssr++QBpU9Z6
ucx/Th3l9cQnm+Y+cM5thitZaK+MxMmrq3PrGVL3qjFCnl6QysUqZdPtc0CD
2+0gwzCpUT4RxV8mattIDI9iyAeNQ7Em38TDIRNp/2/hSdZqTOfOEp7ZNeLn
CQ5w1Gt8SENY2Ldgrm2GLPnxE2yQQB+Hypq2RxNUYu5GQld5oWyAnvjFvPwU
+YU/hNh9zoZ7Qs45GIytdkmfh0LmtVhZMqIOEsAJY7kqAf57lMkxneAKmxuu
1F/L3FFQ2aGKDJcvglJje5ESBN5sXEINlgt/XLSfym1idlK1XjYES+C9zx+x
JYthbhQli8OD8soP2yvFsQQ/xDrqQnQKZb7giP5bYIvAw/OkD+MmWWrDUXTZ
Fko9u9BDBVuXkNGKWtsYIBkVMqmLiXwLldgxKznbD8e73ZPOVAe2J0EIOTlw
35RD78HqH8yfOL7i+OW/+cGIdrvMXlG924oH2br/YDVA/sTjUHg2SdoVygPU
gOppGXVRrEg0dhG2b4VA1wRhQexqen1h5q3POnSGb2CTtK1/bNCSPkcMQ+YN
4oPM91SMUaNBnMkpe9+QvZ+mSxccB55L1dhpUeFqf0j3GSsooukvsBSP77Cj
kXW2Q8CMbihMJ3Ty7OCMTzZELr4oAj+up01qauQigLHw4TmgforVaVZnl8Ha
Xm5oHXGQqkFfV6ca8v3m5onk6tAvDlqfgFz42WCr8ZDDSPf0H7fwewyy4P+3
s6geKSoXoTqhxeY6iiKGKwOrpq8GAc7FYdbKbFxviy2VXXYfT0MHsEAfAacV
aNiRYILD7091OfQrFnCTaz8s8sbAwsjUR1u9w0ASIjLEm+/1Fc/++L8k6yfb
pBUL5hilcjVYk8zrW5uLv9e9TOu2Yd0l1K4UV70YCKDeJXVTBYze2jGOkj/2
BCjF1zq/LM1rxAdJvQhw8rkrVYCVqoF+HBJZIAfiShNxaVsvcAav2akFccMF
9XbG6xLK3T31GBEFvEW0BsmVvwB+eLuJQdLA9d0H/qwJqzCIKLSmL9l8WRE/
TDjY7JJN45zLtc2j9I/N2vtCAATDZz1aXdJHiVX/S8OeJyE7d4pAR/XqxFge
WkfalVWtjT4ruIKt4GiTiisYu2p2fn1WLOnOPaaGc9FGH4EllsnYP9+zt1bg
1bRe9zOUOsX3L+Nz9npuOnlxQucHTM+irdaDJNsRQ4DQahtF/YINgt/6PZaX
rCf3WKgP9W12dMhHJlJW69D0BEbGca26ahhFwQcx1WyGw1t9B+z+B53Bn3qs
gCNdRbIFc5FeHHRQOt3f82yJvlkhNe9wJWg1e9X76uENm7o3l2AqiY4JZ7rG
JZjyi4GrPVGv4t0AY1nMQtztXcmxZMdujIQ728MTOnsqs12XMhonFIMwIdS+
ww9BR4ykfO/pvPlPE7I9u1466l8L1y8lz2gFNacUMrSVWIvEy6e2r8At16gW
d+X7cbbEs0SawHwylw7PSMIAVR58mKP9gqvNpRVUtyDmeasDXv+AddcNL8+N
XVNygnEHut4q8oFgEyndS5yFdRdjkZRRIuo5jtjuarrdeeqnv6jwO9mQC0kd
BA2ewrQhe+DPsWidDQbJQa2ltJZSGjLEngITRoU/XUCYFURsuwuN3W3CvBUw
bhtVETlNNfhLzJd1G0v7fXc718kazQW9f5YOXZiZYR4Xkp9HPdt9Yjp9t7FC
4Mvajae1oFWGx7cINiW7TanZ9gI9sD5U+1pOqzLHLl+0Sw/RboxwbOjOeaM5
Rn6VNJZF3NZmKvXVgQJOhVQDIAHvsgpzwRFLMWpANmZw14cccndIHX1oqaTr
muI8rUs64TVLjflJ2dX9ct5nBavIRG/lpxoY9L/KyHBplQ09ScSeCxjzuwZj
EvcdGYFzeUjyNl/N9PGEGfik8ihnIA4A5aWFAGjQ2QBi6pu/siTgddVjgkmk
bw0SIAilL5vI7MOjlsWA3uca+u2RlKX1hULuADB/m+Go7ykt9WRrqXfMPjV0
4xGnH+qNlJZjsvUX/Sm05dR+/phwZTjgtTd/AmfLIF68kS/tBbu/QMfXERzb
QUcroJ5unOoaDS0rUHr1DcPm895jGlpuqIQGpvrkyZAdwEP8qEb3vB3jbxCJ
ggq19r75ot1sZVeyTchYNND3dRwilpHi7pfW+AenQHm22U4UO8fto6gFJiqX
yii8kNJ/P/AztcMGdveTfF35PshD9pzZLfeo99wDzwbJLcryFXVLDRsVLqiW
qNLKEA5H8YGaCMSKKMFELy6LR1fx/ObbNIso5htDtPNCTRAtTxiyY/uJphlE
3D8rbQLELaL4+5MsXtsSd/Nr7HK1I+G26DwED1LuEz2lUwY+4Hyb4eupJQuD
mVQYvjhLhCXTHpUNe9et9fVHhcA33IMI7Ty3CK+UbT1dzeD2AN7r/2LVtz2b
Qgn0UZNq2OgP2so+LqNPoB8j5p2Hsz++poKyU09MLj+Bz7Ao8io0BCGKose+
Bjb1Uiuo+i7QZHp8EtNOaCTPd6R0fLdeL6g0hTUh5fv6eEWU2g/DodPxeYK9
tADIJgX+/Eiz6ZP3TAwZbxrs0rcM8e7JxmVQuQH3rvP3VmMJmDxw3pwct5K7
d+8cJnlagW2wFV1QVBYLWBxgzQa+6WyfyI3Qtmd0cOk1FKzlmGih826aZjdI
rMcnZ3h9xIk3B5XcA3VJh1YedexNl0Npy6jQSrilTf2yAnZulQHpBwyWlI94
gCo2+7R4wl+bM5pk/EJRrOPu9QXDnDL50bGKvUukb2xL6vX39wjvH8hMpfn9
FviT+0GGKibU9dqKIV56FFGxEBOvjw9RkQP6celuGUZY5B1YiZH3qTD5/WPs
2tpj/FGFU0Z+tfBtmETqa9GxgbVusksUfYgeb5OVs3lFBiQiBTtmEsNLNFJW
en2G0u6j5IQHVz3R1j7jhs2BYyYWO3Tms4K88owqSbP6k/B9lFnLb3Ky9wPV
T+Zs5MXkiXub/Y/j1FMtBGsNf9eeF1EP0vbj2p1bDnWlJtuQWTT6smfZHetI
gKlIUPnMPMIjOIIqLQDwWJfhJg69fB9P63tJS5n2T0KcTiL47cXzp3yi0d3W
zFNlyX7tu392CR95RO1vaZqtv/OG8lzBmtW4B2JPpQJo9mLoqc2Z+37BD3dG
114q5gTgkb1vqTYrM6n96jrVEKTfKO/v8W/xP63lWB8kNC1rvkQ4O8BZ9pyJ
yfzTJGGheMhjM8gE3+khzZFpbqG5dqCHMboED4gIoFlOPHOIXazVgWIyxrlA
vrEfNy2bJIE+NTbcdtZojGqXKm5FNuZj6SDGY/PDhZHIURrfUrrszejplTSy
6I2C2/4XJXoww0WUnCL8sKz/unwBny9ceQc8Ta1YYtvKfvHGhgd0YLZrn8N+
ZFVXwV6mQ5BhjQ2LDuskMD70ywEyhcqcLiir2rmyrwrPG67O77NrrxjHj/aQ
WBLb5AXzTxlrkBJvpgIQVadGD2n4cJZOUTEaLr6zxAvTtPMaKGV8HAN6Q+Zg
oqPtBHjrgUoUplxHRDpoAN8IquBidBCLlVcEsGrNKDCoIrE6Gnh6h/Y1eMGG
p+7hC1qnw3P06hAW4gQK83ng8xNugMhrcQyJw/LMEIJORNAraZtEdBI9JUUz
q9HVPQvQROaBADXgBDDUPx4/rYRFTOC/Rz9HZRQlU3ZK6u/AFbRbk1awFDWc
9vWf437cUvbvo37sR5tngPkVROvV1kMx9Ur3VW8XLXRk+Pe6zU+EhYGJLceZ
KyaHZpX06LPePjvrTsEgkCSMZDLoo2L+0An1X5N+JtgxPruQPKsgHYplBLkA
JlnM1Qu5kegL0k7xDu84iQHGR//MwVSW/orqN66Oq5zzJwipmILO9xUasLfs
n71gNuxgrpCrdNayA6/jH13ZAsZj0GyKKzEGzpM0yQ2pbCLXVyw2M/GKIi9f
vQ9YbldwFhCOKm4RzuyfO+J5vuRz7aCg9+ElQ+IbGIAA/3oy2ls8M6LYjyXe
yY+inXVRPYw+NdsOVN6+5Smo7mOzZBlCe1jVCF37EhGAAkDquMfU0ypt5hWq
rKcdWJ9WxjVfP99XTCZd2uUJq5lXDirEGRvP2nwJ51X03C/uW09rf1ufPh0S
+Aj9/hmVtfPu7xUNETcnB/LEWg8pdegrl7DCtkUuBm3cb/4BrDfJicplRWwL
8xFJtgfXI+mobvvGK11zDoT3DzXRWJ5nLJHrsqxk53hyJZDMZxwhcR82WOY/
f5jF1ewh6RT1DdnQxVeV4vcfxYj7tmOxFHVi2jwwpcNigZX5AE5Kjya+S8Qg
MfOKloyw9Dk1Cw5czTBVltojIQAuizwo3DWb7lkQrmALbrE0k1QEbSXI12b3
D549i77LypxHnFilhyalyDEmURIYSeLEakCpcnX2tKWMjxzj9LtGGzlb4qzr
Rs5j1nawVkiecdDPdM7YJSqMrTIJn2W4+gdt5SU31eLPm77YypdkorEmbxf5
nSNJ6y34xSVlIXyeVuexcu0h5STv+wguwWO2XMd4Ny34F4QIXy8JMQV2YdS1
HYcMjksuWzwPMPLRIMRK79JqNCqjSK53bgmXQoMx+rY6dlvIrpwH/AJGv+v8
/4nY7STarmO3TRV8xP/SenqfSdswFq5snj9EucHV3wZUtyRB49Ox17JAAzxh
1Jj/sStS8WeB+1fFoJ7ba1vkqJLWrqyrJh48+MPia8axzCl682+lkMAUQcuV
+dVCneSG9LpF2Olz3xiTcbnWLRqsJznc/db+dVTbEu6BWjZ6ExraSyJxleTK
vRY4pIet4qdoMeiZ342gxF9zR64MTbvrZtkjqtqSJzdK3Gin7qo8I8txT2Ru
5zdm7bwg+CiNpHpUWeF6HLpHr4hIbj2/cq31QPl4n7H9+F/5EuCYjonPHClC
cp+6v5L6tONgVtzaNsAxCR3LQCQYxwN5TRQ9bdK2hE4vyFiLQByEzE/RGdE8
DOYyqWMrfwJSF+Kb2Q7Vr1wNS0SBn+VzQqowtJC8ZsRauLujRtU3Lc1pqK+t
m2OH1Ib2CwJ/nupF0DTK8koGovxGS8ux+IXNZCHj1yvQLqqRLgU38ueNUtFT
Ltq9rMxJjqp3g09v2KPyNyInxeUSxpWxPe/z7sjmHbPQ2/v+2m3OL0b4V5at
eauAsIXM9sTZx+n4qN1fiXORPNxPpnYcGmF16uKDUKV+gYaOV1Bdrdyi623Y
QYZfmBGEn7J2UhQOnw6NatziCbf5XUEziVqxIUUkR10S+BL2Ser9eeT5Vfpl
iW7IZYqaetJfbUygfuwJ57K0gh42K31FqZW2EJRllF7t3U24pkCs15cxPWBG
b+wLoQuOtYQAcofGMoj8Bn6/zc1povOtqXGMUlaCuQa5VJxhJg9bKVm9OisH
OgOv3KDmdMtN+AxOCNziniAFK5kEZ35pzYGLsip9APyhmMR1kTc44CwrCZuS
oLg0LgBRHvluYbK0Kx8Tyy9OufkLGPNfjt01LSCOXPmVuHDKDK6SkLkej79S
mZ+Hpy6RX62neHrIaIJ6BGu02oMGzMCaUutPSNV5Fk4tGmu6fQEMAD+cpSs8
ewvg26ZnymEqV0CUDftE7MuQks00Fs8CultzRgjUSNsS7i99z9D6TUnIhCeP
2jbilvCVRgguOfDp4xDeFrdXRsVUoys6fdRpEKr4/RrBoFCWQ1snv1s6rSd7
kGjGs+W1myvUyvlwrQ9PUXrz1EPK6KTxa2sC++RaOG+9deWvW9P61JH0/U3t
jc9VsBeJwQogM2iaujM0lpVkYDm/77dEz1CKt6aL8ayZ/W8Q0lkT24YGxRT+
HuunDkl4pKQ9wYjJ2HXsNBxZLd+TA5NLA8mC4rIcmGfYSJxVOrf9RDeXwTCu
OKTMB0oNkGK1eAu4EMavwMsM6CWQbUZKZi4qASxYLbXFOzi9wXv3Xv1CNcFP
OCRwAqOb405f/9FVNGtLo/e9ghvc1r8HZ6O/Xk00W4vJ66e6196c+CYahZMP
t3SWN7basB8ewtdTLnU5WM4R9iNFbzu7B0cTQj6NCjsmIk0Trw0wUsAbuMLT
LJyCGk9Lz3NOflpxYxDZB9glmlNUKwHzG4FRv8WS/mE3wlwwjkbUS3qQPIrJ
e7aGuQB33EMIe0jmHg62efpglANm0ckIOW/oKeTEYD/HH1XBP/nX4rHrA0HA
2VjAZHs59VjsCQP47A9/TmxN08CIY3cz3WtNGkT4g57enXJZFgJtdSk3MeFj
mETmWExuqV8Kqgry0Jcs4BQoIG1t+ovHJBgqIb+WyXYl009QMVA295slGHuy
8RiZRzFaMAqdtJmT5lE+/j2LP8LLz3rITd1R98ufdZJN/R68NiQdtfQA+UlV
EzrbaKp2MnvqrS8/D3l4EEg43S8rl/O0HieGvjT3pK8dvIkZO+16QNDkn9Lm
yuPsst/R2ER5TkrXY210Ca7zrCusoQxePC5NLap1NbYoKQHlUsSx4B17hz8w
3UX6x8mw59Z9bT9Iz484/azDtoRsJFSzcH5W7wTRoQXkxXwJttgIrsx819C1
40TqzTa0NXHW19OVz0cbqVrBpitX/abQMhWehsPS1U4k6KOQhvjTwGa+5nzM
EfULxhgeu39T1ojSOD3AOC548o3TUSAtSIvjFWxihM7PEZ2H9VFzz+3OlQzO
CCvyQF9k75sSqhcdd/lv8Rrki2WpoHt8Zw+PDywA8eixg2I8vI0Mx4op97ht
3OmxVfES9+F3AJ4g7eUzxFmiSJXZ8RRTNfL7KDsm2lbjV0MR47WPi1z9zFwa
6Cx3Qkuqn+QsxOANQZcjqf0VPJLrrvqe6oRe0vV4TacyXvkviWGas2KVnomZ
yk1Ind3a3NchrI8npX2KdEfhekvnsKuq9PZyczJ7Ym58IERfxc0MCOtjdJjL
55KgJCMlwDTl4KuY/KJOsvjAndyWpkLU2APQm0DAZ5dyX4OdZ9P/Ugq/5a+C
CjW7Zy3GMn+nHhrzHalDVvAvzgmBtG4Mbrg697fHy5+5wem/RSHeexmWT7qk
+VX5gsGWay8bwvMbZFNK8wKBttgdA+oxqAjYdZgfoY3KyF8+yTfnFMBe2GI7
UhZMUXQWFNQWXSPdL/O3CQBZAgAgRIELYWsimF40bzsoYwImRWgpu3cjXiNX
ivYhIn/5mhUfK4l07VKEX7qqlxvYsmwjPP/3s8tsU0/ih0gKyd0zVxEYkMzP
NbVz57oBrG9CnJxqP44XDEgpaYUFWmogSYsydywiy/r+pLB3JJOiwGuaaD6q
1QqNVrxBtDZnBshXQVV6i4jVNLzhbWTSTA9w/pxh2po5Btpx7uAlESoh62Kh
W8mx1WyTf4+y/uqH0NCYOXT1YlEOYn5sMbnJ+P/zpWkRrs3+oOxMP07ugmlR
nKn5RhigCWnvQWNlYdTYxLLq1encCp3qOjVwdxHERHjfwMJhdF8MqbdXkaBh
SdM1OrEi4J4NF2Zwn05VhD7w+95d4ctSyctVOfXSamdyKpORdfppXoBitimZ
r7DJn//5UznBRAJdKYpskpMJod2e7gH4Delx6bvEtODLniQq+Nc7rWmKXZPP
HHDUt99rdDN8xTcPswiJGq+qGe118+5mGpdbhZuL2hBSWhIrfO1x3wqPc1I8
tQl02epJxJCfeERUhnDCzpbpDa3fEl6cq+zYnWbWlLgEJxSKCOP+FhqwybiB
M5XZbRx0ZcidHGgd6Yah6aTZ5cwpxIpHAn8wey1trNEX1heX16YL3iwQCprE
voWxFxT6LMGBvZjTDxk2Y/T+BRuH3t0cpCbxEXiOMqoSM1lR7T0yGWzHHwgb
lbgXuo5yxiwIcFvvuYia/yUssp0L5bKKhFN+GPVKqtg6PgbSo/1c4CQeS+2n
c3t8itxNTXXsWng9gAETLk/y9t+KTrJtbkxsU38U4xrpQVHGKzGcHV1CNJho
geTR893UBCqsqr5jyjP1R5h6tB/Plk7wJYmcErGH1fOeqjxHw8egYY/Ylrzy
lNLC2e2oIs49v1ypIKn0w8zJNbyiOMhkEKqMNYkzO0h0LGx4De9RJqLCSS8t
VK1L+sQIRJMWoMazyS8GZDDmWvS95v80lr+RGIf+Ln6qz/TPlFwlOEcQZV+z
Le2XD+DTPKlAlecITqMQev5QqIBAp8TFDC9qPSzbW+b1PROiXYe7jWcyK+BX
XFTxv1GEwxAgqpYwsar3EgNuWilZ96X5M9r4ys7YBmzonQ3mg2IGoTgslFQs
UbsWCtz7ArkT0c8x4Gy8p5sIzgwOpUMYA8AW8QA0SJJgNAzkWGpjLnIDCKms
IqOfTtoH5HxTUEgXBFUf1CyphVIC8uqduJFlMLFlTtJFrRLSavH0U1jD6vW+
/Lsj2Vq9L15snxbgLifp3dMGhWQn/eu72c7mKvvWa+9S+bLYN5e/WDjDV6iW
KES7Sli1T6Tyk1+nLpi9cg6ZqcuxDDobl6mtuTNIjKrfO/ru0bzwothKaEHd
NbvLwwWJKDxO5Q+Nb9sBt/BnqfKcx+LuJWNqQldNWAoeBucr8kFPRIGzt98Z
ItOcRL6yRqRkI45f6yifbQ4tRvFrdq5oNu78y2tHCzu0ioT5kIPpndceluqH
sC1isex6oTO3Y3bbsDONxhKNSeyBQSZtJIYGhu9shuHj0p5U44vLhNz8c/ON
y2wZkv7j9OBWZrITWzW894gkq25bd2APyhRcTPDcBbzmk2LOsBAHl5/7r8SD
HVzcJqAcPsiRWmjNNYsvj5Vre0hezx+DjVUghuVAYtMye/eaT2AwNqMPrvvv
rbCUoFod7qssOJNfZQLW0IbUvXsods6qj+fO8mBMe3LD2ivTkskxKse8cSs1
5SeZX9uRIMJXYZCyKjHldfmDINPKu4U9eenfM4cABPp2HwQ6rpRu43V0SlDQ
kjH5VEBWIAqMAeRVje6acCNAgeZiT+poU8j4cNyE0cAcOGXt1CUA+Xp+er8+
Uk0rFDYpMvMAXZ1NMEzUlbfTf3p7BHopTHzUw2mqpLLVjLjMvnMPwW7Lb1SP
YGdKVTOdYeu5GscTKCswvmXVRYFH4Hzh/LmOkQBUSe4Yy9RDndMyRhPCU36B
ylMUZQCCpTtF+yUOkpjs0fHS888gycHthmV7ye9F/R/YufDoj3GkRJ/PFuNU
eKYOAYflPXHOnGfRXFVVCgvcHNmU0cg+jfbNtIhRPH/82FWl03vQ2gCP/vGh
64xFb1j0wuh+o5RmSlvyb7tkgUWrhBXt+LHdQ9PoVLQT5BZ/UUhttkJfb0Oh
bRuphPbraYxw9yv3P/FXProL//V6VGEtHNTA3a/eSj5Cry7XcbJORi6puk0l
1nY+6kNvolhtNosuB4oo9TB4rFkNqMkGAVdvTN2wAyAhUMwHbFyT/tjd/ZnC
04GSf7qWvtiq7aYfluqUzBjOClqA7uUGktoXpiyFrQZr9AHnV0LpRrkk2caE
ZODS5N/b7OvK157cexFvtHL+/kvd5tTWjlCaR8/z+mCgcR/uB5N10K76BHPl
WeffP/uuCGIMIeHZflL4R6LtVOTIVYwNh0rUMp3BphUYzzyjXv3Qk5lCc7pR
euGJWqHZ/eH2nYSlrIqpvz1+OtYE6k9SaUXue9ilqXUZE2gAgJNqWC/X/hN8
mdye3g1imm73nj0x7s2xbhWC7wBj5/x5gknFsgMJu5Z+PXlJDqgPxp9iWHRd
7rsTXQlkSPnSgqvBu2OE3L4egTdizC73ryCTLxbIFiX/BwSxJKtd3F9pJBRf
swwT0+xbR6va+4nDP2krpj7G+a9qGDqNsKg+PqERDCvdIMbIdj+KDEk84+MZ
FgeLQoC0j0RdMnWdHTwrtFNbteVVLVk6e6nUhz5BzXi8mWa9h59FLPo1Lmkm
7pEvcZwzx8SwefqfD14qXa+GWiprUr4f0/OSXOgi28gwzIfO+kY/dcJb7Yvx
TsJBCI3bYr6azCEK0GfW2Idg4h+P3M16AV0S7KvaTsqIiprz13bCc7lrgFmg
76hA9HrkTHzxzf7VTWZTIx8LaOP9jPrLn/x08KJzrDwwiJeSR/f3hE/57xzL
FF25nC8tDJlULQkX0Ke8qyT9PRq4AE3NSmlrCpZIpNe54Aer9fhoinZ3MgC5
0UuL8NPWpSLvNYNfzg18kMx8376fO6294dPNwHSAu36n+UXY6mOmdShnZrXh
pyyMINpt6ffrm50ghQ7FGAqHrO/0GfueBcwrVM8JFDSliPXaSuyT5gUKetB5
BgyPj7+0kGiQJlzEROgn9nKaf2YsrZ/QtkOXdTUck2Rc3IPxpgLj9Aun8tv6
s5eXJm/DbMQuIYXqBxbjHpHZyjcsjvEURHYJ3p7O/f/bF3axT4WjHi/78d0O
99knH+lrIFPq4OcGF//4n2jGkZAllVn5zhG4TBjHaajJ6inTFJyp+6pSIaR2
G9I/rK/dx+Hbg4pOAwyo3yKRc8AtPUXZhSwHxudIHUIsTfEpCie1ph5SbMg0
sGFvxmEh8xafz2m6zwjFCaswYmyGSG0UQIkNvtIb/RvP3vn0Dpc6QSvRukeH
zJql7/bNczN9Mew4IvhYvlaAokU2G9opqyao4s88KZYEXg0KKSXg+S0HAWEq
AXPGGGhfm6uHrrR+o94kR7FoP84VkNpK2K+vZOE8BYWd/qg1mPeyJL7y8ITZ
HXUFyI1iF5e42DoplhoeUe+AswfCTJ7XAVLqebdQ4Wm28C5jzpc2Xci7FCid
aHeM0w7U2lzGhtkGEiKHvpqMED/5N+ifqQvUVNGqp27ZaRoz87roT9YKdYER
evMbIG9pfwE+UwEzFJUx1NNSKDqTr9RmmmHE/wH+Ypk/r+4IACVjg9VSajzr
aRyqEqH6bD7vEoRHaEdm2uKa6C/3dciqqH4xlCd7OdDRuYCp/aY1SoNE0U9x
JQ8F6Z1NdkqggRgdi5IdysMjhS7k1ygWoN0xgpI2vCjDjR6zkLK9ReDHrtcB
L6d0B95H2p+lR135lmyc9poLn8Y1pjyeN5Bh4sin8MIsjmyqyK++KR1Eh9AB
bM7lcPPWxBu7WQFohK3Asd2trIz3BKp1a/vYvDCD3b1VnJh9jscUiK+1dlmu
RYNq4X50pP+4JQ2vzwkMAgo0LVy0GaRlGQnzEs8GUKBuG8FjJjAWiwa8ClLr
N4yqKB0kXUlugTgo2LmP3SMFipiny2rvVRCbkWbbPEoHIUI9hhb2QLg0ozYp
w71M0BI9uM+63UekstappNHzAb6U/qr3HP6S14H7iHeSbD7WE/SoHKQ0hawJ
9KVHRmBfkDZGY6zxHuFW0TRHxlxhFY71f/aPuYscS0aweYemPdeiOl46zFKZ
g75q4xhCsQQMJXojxyFLm2g5TMW9vhvia05kNCtP1s4quXCbK8T/6xMfF88m
e0guztx2n6cLAia0gsfs8zcrFbh9FS3RdqTA8Wmm2g/DAX/kNNKgsurSYoY2
TF/NhaGjlWGM7BKpxMNDGxSDMznkJeXbudseNfiVU5PJ70GV7cvc/Xl8ZARO
sq3ZTaH1BzMHikBpGNcBblu+o2F4tOsoBnA3gROBFKLkd44dlmprXVfaAVVY
cvSF6F1Lgl2sPez2O+7Bu0KjGUTYIp64Z4evxKdaK6RA02nmVH0nDqSBoG4q
JqtxBmQFsaW8rjNuVLOknGw/PrlgfLS58DA9GrmnAdaPQRPH/kYuEvA6Jc7y
NZVKKavs9Q1fJVu42VTnf/eJwXoe/a7ONKb+utt1GYpOFhHLmnzZIHT7p8dW
jbDifCd24jEWWzZE74NvGOFNheHVUZUKsuQinFcx7ld069yZGwMPNuRzcd5s
DAwPDlQYvCoMv4LMILzcfqFywl8O3kuFutW79NqICpWzBaiUh6AxpU6rSYXm
UdnU5v6y0dC7LIlro5IthUZM1y49DY9H8PVdGr0b2Lyreh8eEQE0pfWMH7r7
58o/If4CGSGRaDtavR9AnFsu+iKXhRk0SsFoupYcqKrtYiEp2dQQIiKYYYL1
wCoztlDeD4pQDCfTieDTh7Y7KXx4/xijyFSTUhivqmhWKsVFD8Cd1nV4xaqk
h0Y0lt0PiU8NzFWMdS+PjaaysghFAfpJXsoTjQRkdX90zcqwai/SqxtlHxVx
H+jdv4+JLkzxfIOiJnPTlTk9Y+DgqTVdMPqcqZmHsVDFoQWJY8u23N//A6Jo
opgnmHmHk2qN3zXdM37JvoZ+l5zL2KX9cLoyJ09nMJR0HdgBgaeq2rETsLdx
oL4kVqCASPYPK5jX7piSrWgmPCWdxwAOxAwQobrDJ1Q8avzX6oiWk9Z5Yfyd
S5cOQxU0HfT/dpsnng3KCW0uuC5CnCNpcyKsP8hw99vbI4x+TgFRKt3KEKhU
bO3AL9a/7ORS7DFkgZHkf16jgLvJ68THCZtOIzSDrrtyUxVAwJizts6UCqMT
mVi405SbZS0HfEPlw0/tG+0NgVApFScCiafEJtl/Op3pszC4WQP0Q26d/ZvT
v6+aJ2rurMmiuD/t+AeHTpGmGMYAE4XPmjlxeRcT6OfYJI9NzQRKNMRYKmdP
2iXACgjDqq7Z8ywGUWwNTBtvW2ji0NsIz/Pe3Uwv7/LNz6OReFlar1pgLneV
numKAhZt3Oq3WIbKTf4a+Xfns1SmA/EwAS8gynV84Zeeu39dQngKGVFGUQum
AD4crhbVq16WrqukXdOXwDUAKqxt+qkhYk3YSPra3DF+ePm4l3uitEVeqT3t
2vjF0OmzL5wJCB6hGg1BeoDzPkDMbJsCoidzIllqGnrIhCF2aJbCzncIngQ7
DrLsloc9pmiaIbO/fb30j4oQWZ0XR+8vx9ipnK7T6fSxWBsZoJhXdFy+L6wp
L+4xAfoismH5JvTZysaRPOuTOcQWSxWPWSLST/nOf1PCqKSy9rCuqRVkJ1I/
OIIrY5jOEXu0HoV79yZXEHR82iXdqsRCj5nBpH3vAju8PM+pqfkPzHPlDtX4
edmP3mX7UqoQCS5J+9BDZGEhtF7X5KwbQVJQcRlEzR4H/s1FE+h7BChMPHDI
LitwwUJaVx6t4dMzWZ308Isf4y/x7RT/8LzE0khFpcsnm9ghpiKWYGE9UJAb
VjdbdGC5E/WVw9EPo5IimZWOFD2a9DIvQCm/2tKlvf84oAKwUMoB8e8A/qDP
w7NbDfB4vilR+p7pKriTX52R1MExAGRyXnqWyhIfYL/+FavdGhUWJU+uvjjZ
LLh/vrVf+MX34BiuVgGwmVDdIyV4ukk//oXZlSDiq4Fo64O0Eb4XinX01uj6
B853Cu9o1MUI53/Vdy+uc8hOixdJZv9P8HVkMBQgWdnOFLPq+ilezNUWn87I
gELHRez1g/R81ryGlLLa7eaO+gckK1Nz3Rn6AV6g6uSd9Kelhlc9HE6JGg69
Y5/q8Lnf4BRXPE3pDo6Tuou+MrncRTaUmmos2s9SHvWyGOnEInLov3u0tuzk
NfH1pvuWJ8HNV40BgliqOJzPpwniImaNE3lAhRh6cuwqp+gpepeCWDiAz/ia
0akFy9v9gh6eyBYmkZro50hX6KHe946bojCN9KY25SVp4a1AZIKueD9KbxVE
GaPNgmsNIZsFCtcmHZw5o4os6SlXyJQCQtb2Ne+PcPI36WQFrxDOqlEmmasG
NDVv1CW58a+2EmPr0OZv+izFklrAJWl9/OFqnl2iaBR8dlzwx7pzsJoEy77u
T5jY1y6/VcxOsZ4WystDDeEKWsiFbfio4WiHuIb63YH0ot/oIGdsOn5eze/2
L3R2gEXdVmbBJ2QBCh9h0P2DxfQS54iqiI1NyYYBNZY6nR6t7yMVSR8BQ0qJ
KTFOb3Do9KTm1lQbgKx8vpnGtuACUo7sWZ9TWQUbwWfMvkufeUkqXdyzKKPF
eyuKM6H1CNCILVGI8nr1DkNDBAEpAdBmvnbZJmzxfzN9EuzBzvtxucEf8nOY
hgsJTYpFFzDJLurAq6VwMnieu6UKZxgyzLENoOYp+LzWKDYRKj+6xonUDEDZ
w56G18Zv2VkiP5R+WhJbp3dZQX5JiIBvDQ4CVUSN/MV99ZHMBs26IX5DpvUJ
h3/9YqZt5lYPEETy108/Lwfcqfp7ghtO+3grj6dMEw7nxeSwSGBjFj1L4yLM
82t4bkbBpAPkQgx/DP0iTd9GcCqktrF7EWxF6hpC9sFGQezhnh6TxpU1DEa6
FMf9+h/roKOrdFXkLHnaI4tYm8SbsWfQfueKVIDCqHoqKURNzl4U4j4QxZhF
fxn1F8UgIAd4ZvEwYs12tAWOAeVNHMJV9g89wVouH0BR7Pj60/21HXjllEZy
vOkdEZjePpgwFhksWNLs+XlxhN9UtyUHqN7peNKAXHMZ7NX/4C0jEw3TurC4
Nw533qS5f8UgMUrwoTUutEy1iDs3PBpHlgfOPGSItISJKM7yCddoo1ebY1+f
rNGdJvpNUeiw/tzd99BtCT/qwsgf/jwR/qN9RGzoPf5ybJyijwlpEPKTpL6a
vQ7wTYYBgegMfeJ15Tgs5FIMHaicKhE8axEcFEbuLN4o11iZv/MuYpEOIcUb
HyXaG7zeTbGk0NSCyAgYaQC0PzO9tE5c3jQcnAMhiTQ4UjurgwOhMnvOnc6o
EQF0QDzbNsn8bnC0kF7I/kBQ6GGelZ/v/3Tg6hVpFQZ0EgZCqh9jecueU+Ug
eU1uy8b0f/iiFe2ulU7QkJm46VrHkz66dWSixK6nRd2blnj9oSPOBFmYtFzi
dcoPZEIcxMO9nNf+yZLzK1bak94DX2kofAMBBUr2+1kygchJC9rvFCWjZOW2
h93heFgyYI3FNgLgsyXyu54FwM7SqdjSueZCsqIquRD6QSx694/NOpx98m96
f/3ZrU2zXFDOFyucDG22Y5ycJApY9j+7dcAbmxS+AfDj0KwhfSGLzr0V9JeX
BmebWdLOASm/WcWcpd8RjlvaC3Dj8ibGhX0MjxSOs2woJGblZhGsMFfoDGo/
EO/KT+JBzjLvqS4SyY4W9e1gugPfHkR9OoyBR2p1mbI5RgvLtyM0JrcvL+aM
RCq++jJ/JkiqoMEuvqmbhfR3Wbm6nfb377+oHkmxJcuWkxNZqJLZ4i6tlMn5
Jxxc/esUb6HGJvoZMhKTzw+2R3TbXbQ+5y0/sGdekLb/VfB9B/OaYqrMrNzp
fPyFjgAWPguSYMon/YHvYqMZ+7GlKn6aDtYU7L6epYTj6D2FCnBhvKi/M5pY
051nQz95DZ2DCbqbwIvUY8Od9lHjXkCXN18CukcU/wzTYoqVobiYzt8Q7DAS
sR0+fAj8eci1Bz++TsFYX/Zml4xbf0O8LTHvftxSDuVSSjuALB48aTa5kyv3
HwuqKqYLi7Vn9HcFBJEenhG0zYuY7AhscGOXNZ+Z0uWgTNo2S42ExJ8vydfP
yJuNH+Lp1whm9YG2rEPsXXcOMbuaZSuuKY6utLqDBh9t2D7KfwfX/aybjZ7X
SMOYtV23hQpzuMAv2VY+8ionPPf+ClovNZ8B9uw/H5whRa6qRTjQ8KJhfOdJ
G8+nbZP2a/OG4sISm43p01aTIn6MJyQSxtHlOvKItdsl0Dq7Mws5B6JkksIN
4ApwoGwvHdeVsUR9eCQT10Qh7cHQdOTfAuwzT4DyCm5XCTbwHr1hs4Dsi6Vl
F9rqPYrOUsMhsadX5vpJ1nWSEFON6DLoUrgiDTcUlmXwvJzaVF+xtOPKRwUw
PUbvxnu3xqrgM+y1UPM7+N/VkX/6CYQYTCVMonjwSicVMU20D8AS5Dv0lX05
/moFOvAi/VrcYtYqKFJogDvnMxuuEtFBLkyvflvc8FFqUCPEnM/EulW1HP2n
zw02Ip9P/OfxVZxuD6nqC9onCNXrSIsq6WW+P4EdbywzMEo3yw5U74N6JLeI
t/zO2HickSneb04vE0pLXdxg7WlC4umpqlhsWDSkrXUQJmRa1EDZOxVtGYm0
tFuz57Wq3eE6E6pU74uY9irSBLFZSbwPxqFo+0mrLPFps4Tbs2iC7QLoWwgo
Qc1o7/BbIf3G4Z+qwfpDwfSPVfY4UPGWGCCd/yRgC+aib0uYJXDV6hRbtOY4
K2GPL/9Ff38McfjQ5h6lGt0Exh+QuIa7ZCTJAImODwFWuxfQobhTPJppIkpL
DDFu2Pg5poxFsiFZZ+hkHoTJtqIIbY9yxlgSa4VjSGpsx22CtXSP1kUOXRO8
XnaJzy27r2WO68cAkNP5u2X/Ax25Ct6fhsrDl88Nkalv8mvuTYN1+wPQXzC1
RqlV1x8RGcT2zFuie/zlOCz0mvB8X2ErA/+34fgX6GZBcsteUP4tY53Gy4uV
jxq7tBK6QVproOp2z+bTC/qM77ibTp+oZ/cjsbd3dRFM/Ou0wQmzQiK28IyP
FavWFMPpKJADiRVDFkHW1aTzO3hnNGpEUy2ldSDtQ+eI33LQeALco7XVEBTc
pIAR0P+7BrUVzZuag+oph/8nRE6v54GaudYd0VvSG4Hri68EYuW9YiE1fIh8
XnRAEXw3BCinKamIrzzNtNLFy8YBXVSa7pH0kLppOLsmugcS0LXnZOja/DV9
wIHy1dKB+HimIoasOIkeBaNJRrCs0ixfDFlP7W7gwKESnsqXedHEowMzghuT
N8YW44tOYt0Ut2onXt/AFNP+Kter3zqLtA2cS9OY60goWJpHfpFHDd5f7kDT
1JO1jFNM5RcmMiUL87zCv4/V0AqVr1DJDkamXIO3pD5pPH9W3jLXgkdliRCT
mbfl4Vg4XUfTellibs29OefKSgBQyp6lzuvPWoNtYz8zsUMjlsmEj5uodj+S
D8T8xNX3Dk6Hx1gQV7ZMR4Nq9mrC3Y4E9bvqvyM7MAmo0Ngde7hW8PPeCEF0
S8etwWYzhLhr+4rirMQgKPS3NcWpILS47+/mZ0G5s/byjkQSbopgRs0c5X11
8Ni9a9R9K3XBXYtTImV1DJCWiaj3w8blKSVvfYDPkGbIjZh+S3OqP4WzpyCj
yGE17sQpom1RTIEjO/Y3FrpWyLFNRXbXAWd7nE7e5ff2rBif0cyost6ZG9pc
oab0VPVjXWvHiIjFE8joM7+j4DrmSFTyPHiDGjQcBRupRlFoBIjG3vfAECJr
28+S9mpOhDjylUA1jmtxs8xYiNLCmIGCe9JEnVHa8+//YxVP/9NMZyT518j7
pPgJ/AzRhHSytYW2xdi9GvIBGCQHYM+CuPzevM8qhesBygypwBGtyZ+eD8sj
PS9gDHiqFOR1BoGG9B9JQBUgCeaEDJVJJ25hkCP6Ev+XhPMeRtnh4I64KLQa
hP/4C6UAweYJOq+xP23j8W9hT3TCFWWraMQOht1/l2xiGr1RVoy9JrBlr3Kl
xVpXvy9AA0NkPhuIdkgNgFt7ir4ORM14eZ8oiQozdLZb2/bcBP0o37zD5/hI
4eIdmYLBPmlUbKRsKE388XTq+1MJ26sve3ITd719+GDXYWuB8FxhQGqs4z22
dh7rsKF4NqCasV6gDuKRhTp6UopZaLxrIIcHFYD+gBQWwyiEQO7sNxVGJ1xl
//18uYsHfigWLZqhSgmHj2VrTmrG+JhUIMioOv6teOkYSc6w/nkT+11nwD5d
ENTaPwEfmLOXd1BZI7KJUZXwVTkbBB5gGuOEXtCicYsldzimM/dm0pAMv44R
qsWVwHVP1UdtOB54v1/4LlUIpLwB5509r2Lw5xyEn+Z9s85nlQ+MaLR0yWi0
+znpXdKethFCs5MoDg3vQYIGLUgQOkSc2+Nx1KuqK3ba9wQSbgSSosG9AtXl
QK5wzuJ8jRKNdN0kT+9qHTCJJGReeOZcmOP1R8VSWrA0qJXztFA5OI8/Rzdc
O2aNGcTw4hwsXPQ8dFyTC0lQK4H2iTMr5USt/GCB1GcpAdYtg+HlfMCnwx60
it3p987W8s5klQtZLXx619t1P1pWlD+Bjn1HM6HSJ4cVy/uxgWk9Pa4wGYjw
hfH//GHfpNUAIh/Gv0k2DNNJF0+Ra18LnVnpPfrjTVaNw1Q14AcKHXYrNiRo
XvbyIxgxd8ER2zptQySqhuf4Bg3Zaw2Npv7SyWkYNAMeKM0u/V8YD/xvmkbT
w/TwqfwXRFfD8iKwCB9JZjMqLVIqyqc/rKgcn0ZpDLqDX0Re7KEc5MIIpvlO
8qHD1MQ54lyH19Q6hNYnaYFUU8D21hoFBhN8oNJIUlmuW2tOQxSCS5AuXA+m
esPGK6uGzT5tQv9H2zlK1VXLNcX30EjNnEquT94mHJUb0Cw+SqTFE49YZpST
6rcpKfBzXoFDQSxw1F+M3VqA6RO6GSACflkveSNEtfNX+mBf3Xskev2/5k5z
RsxmNIfuigwG3whG1pgvzsVVKnQQkeThajMtSWpsEjrACQr6SImnmGj3suXO
2Dw0w1pzZrArfpmkU1RLxNGiLGwanR9KVl7QA0jN+zgSk6B/B25egPVd6JHg
AXGpnY7iUwqZte3kME06bI9xWm3d4J8bY6geXwRPvbYwQzv42/NUpmlzvbzn
Jp9fAjkPKL9iYw4BSkBbNqXhmKG4oegJgJItaWroOtvHKX1vp3dvH8WZTpPV
YG8YfawKczKXftEOMxtYy91KkxruX4NdkV2x4jRk/SNYkVRdE6RtLJjGpu9P
ZK3TKKLXRujFfVMx6EFKk0jkTEk+Z3BV5w8Iz9m3SKR4XLCBhzzoXZBoWPhs
ZFLSumC5ap1Lt6pwYFLZWEQy87vIPLnywIfUHaAu1Z7AjDvVDiZ4/7KubtaB
4b5nHfFxepWnIqscN+jt+aZNrRFWRfra1bTC35Z9s9HSxnQJMrm0zcgO2Hpr
8yFyiMqBtfX56n7Ul46fcvWDzGNfkafZf3cB9hamgGGayYh9rP/h439CGYE7
YqTr1ONWn9/53JlsS5LpnlVOHRFkXNASpomxVV1zqpYGXoet4I0zhBXqEuP9
PajtLqzJ2KHcwXGopDas2x8B/mrBqAzH/aak0tdoNy3H+n8LnwYosvNbsrkl
hSisfrAr795acNhozjS/V657rEOStIrfxHX1W6lt4Rz+dT0ey4FBLBWfJbxP
GGDEUchR7Bo8uR1ELMVRPsaHJypcxv+oBBnY3cdZx+LDpt/Usf/x5gGdAOtL
JpOsJSrlhUYnjMDSivgb6bEJr/fiOV/HaRMHSsTP1Oizqy6APUGwWA3IcT4p
9Dca9Tu4n3YFYgOVPWgigJhFywkIjx7w3OvRKjZ7xxjuNvY62M0Ia6CsDgaE
j0d2JmVGrOi6SLYeZHtMpcKzQvJ/d1YkB7GeMDSF1d1vDMXVIqxwsvJ9zeWP
NsSceVqp0ud26+a5w4iRvqdfpsyySgT6jyPmNbHck+nzqg1gUrpvW+0GMLVJ
9kdIMD7obXvBgQvZQsBiLPn4JT9Gvrwl8hT4j84p/ZVit52lA2NhBa5w2BhN
Aj2jpNdRMUj+CV4mjFGujZLq/+glQmlaFb4yGKygaBhrdxx+jESmWaZdXdWo
waB21VuRI98UV87ARWe21YxRdQH1AZoFwa/1sr9ZNkThqSzJsVmpR6za2iwk
snfKHWZcHULdzWvWl0A6+uKeBj85HB8k0bsZTFPQDEEguuPcdEQdHgTgQblp
dIZPpNt5qqsbCozXCCMUIbUhQrH5tad4aiUQH9FcRIWNg2oHK1Gq/t9O4YlO
C+UwqoxmuRFB/WiFTsQMHJnbQZRPHWeYammRTNehBkqHzcvUZ5FVj6Y9De3o
07ssjp3NW2/i1s05nSL4PV7MHGLpW+Y5BSt4vaIBO16drsGJyUPt0bbHDIpG
Wq3v9nFvjQml5w00zkoqMg8OvZZG4bMpq9PUP0gIvVlUsFqGDYSdmFs1XdMF
m2bk+KnLptKLpla/JG1CA2rnE11mFsnShLsbN1QorOWoShZg8758sZGD1Wbv
Sq1AiebXRjpP2n4oSmNiqhg58CJrgWZZTjzRv+Vd2DTgAYvfucGI559XsfDr
NYkobuADJdyLzNteq0O0SLbCv16pSll9uaHlgY7BbHoVPE6JrWbtx9AlXdDX
s9rUovuvMyZ+79C4K4YW8ikSDNPY9jZoR6GU+ICN9K1qrbMCk69o4PUX4yWY
uJbPsTafPnq5qklpG7lBAN58OA4S0DS1cSHSZNEiuSYufAZPPQfsir9n+XyQ
OmFiFirS9iY1nqYSte7P1ZNkv+X0wbvvAeXasoRxTluz9qbrMaLDy8RmjqMe
HV8QNJ1l2UFihhq3BFVkFYwD3nlJoqBtVR9C9GG5O6lVD/169oQbfjJnrhsu
Yrjnmsvjpz5RDt06yAP2P1gw7gj0Dy1hR36Qg84Qg+09zToC0qW8a4A8ehDf
kQ4LhxBJJnoGhRqWQOgfuoLoCUNs/sYMK4TBJJxr46ajKEqXaxLtZds3pmpV
WjpKKT3/NNkWeQrKbv3kJwyvlKU1vcGUZMwNSXPon+us2w0mg6yZoR7yqT11
4jcXHDLdURLvMcnWuhI5kzwdgpaEWCFy9QbiXjrM5W2cbMwL8FjVag1TasD4
+xawZ8e7V3H5AhzoBnagrHAwuivkC6tZcka2sv0UtAcMtgHEauEcN2dThbuu
pvvLJI6wKewMri4vQXwYPQBiV2XlQmfb5mcFXlS5Ct8Th0E4A/PNjQail7NB
x+7laePyfNESBpQwgvrTQ4TQ5vFRwOtV1Hmrp7u5D6htXzAww3YXsn5olmOT
OSd93m8t5lPkbFGy+7VLLHTzLzEpceE6+MYPNu9hOzqo85mrtP6JuYmtOlbe
yxD/syOJkUZHNwsyfuzLau7sTCwJvmh/EsRuT2Q6l8RNwgWq3Ut30Tugn47v
P9VbrE9nLE20vf4SuXaM3mST59DNVIHIlx4AJHZi7AzwceuMrBvAY30IGsJ3
0rxrhkYRqmCzcUHD0hHApqq2sBQWrTTAPSa/U2F/IS77UAVUGkORZRKxrI8Q
BO53tdDg9mJ1HW/lHAR/z5VKS4OyLokck5c61q+Mc2bRHMPMcettA3GO5m7p
5rxwpqOeoxBrW924o7U13m9i4slBuxGXry0hmvE7qe4NQJZOBYQQyvcqDsw0
e4x9YlgN0+7oiadcAv++EDKK5Mrm5t811ptA7q2dUV3LsH7ArhCNtLbHXuRZ
ca/mQ4phayz4QTDF8cnrGm+qXWFbUiS4hUHsjS69SkfCTZJ9SlLR/gAxpdg+
ng4X8aTKHptHEJOO9B6xNRhfYRNQPAJYAhvo4N84jITxbHSVMdqpbTsXNYKO
XjpKRSVvwXXfD9akQSzzfcYsA74rcPse2FVdZlkvTn/oC6rty+tnj/PN1OFg
gwtOe1405i8Zl0GM+OfpmkFRRIJe3RnUkG2oy1cgiFmckwacrfUsdU0qK6Dj
X4rKmNGWTCUTFnZJOkFk46zdO9Gx4OWnlhqijyRWSiuFfLhAJ+4d/lbsPlea
pPenSWdxy7hci6g9909sTbTR4kp8GfRQjAgRlw+WXasT+hW6jnfsziJQeksQ
UHMrKl+/4jgO4Er++YWxadoqIpK/Feag89pN5JJU2jrwJVFphVqGmJSIAfnt
/5oPR85KeLQ/pRlVtVsKJA+H0klCEe3Te0YEwmlHuAvRAsOufnXFeTIqqCCc
iTprUaCeT5OF2B5nlJ0pA/tP6SGkBeoiT/nCzPS8VFGEHEHKJwtpAuCcCjvb
Jqhb1SgkOgJA/T8kjgFgd552HraoDH9SAP55hhDGLnk0A3Ojg4jgca4caSuQ
MNxP+HLAF4MyeoOqjcthG1BjfaKFOc5q0qAlKn8VreGO9QTqf7t56EA+0pFA
Z6Jc4bnsfdd8BJ3miQo99uQQ47d1o71ovxij0J4u07ZzRN8NYoiYwGaZrKq1
i8XVRcBO5Fxg3a5PB1Cw5QKYhZdHRk7uSsMARikPMz8A+WGxP5Z36i4JlJ25
kx9/h95drmQRAf60lCsZuqePvd+SbljN/96wjMded2KxhR6MzCTPrgapHJQ0
7/x78XfhsLgToSVpL+n7XdOZvlPFwhrHO1gys3zs/E2Di2pixzYKfvgYTrsb
4nuE3WTQkRxaAs7lPrEXQIulRX9RAdzujfn8RLWFhHNaMTcLi1dv0BRKPWG1
pcEhmws9e1RQVRlOC5bE0stDQSgMENGYOpZwjCJOVmkK91dJKW9yHwwwIYGv
eQTlJFTm/sdwNJhL245zHrtmwY71BVFJslMEU/mUBmfxhGUxws03ywb+k+UZ
x52eHHoXv4n1AWMloDCJSM8asQz7qqp09vD7QtBp3W0O9X+zRVDL4BVB8E13
nTY4shZT++y7EB/Fh8UVeauZpBOMGnvkFGyDXJ1XcpDcf79J0w0K7Mpka6/W
KM/zMDA9wPVk9BgfxSxNBbjGx4APVctjDFJzcEG7Op4jiNCHBVNb1tFb1Vwr
yycaJ6uRdAXze8lxLE/hke5JDwhgi/h6Apb0gnaYe4GlB5Xxgq4qNyuzxHhm
6csX7rUyptu6+Jb+nJ2iCiF6znm8CwH8DKGxE9EHQNf/M8dZETJjLUFWRMyj
uwTQ4sozQcXiwA9M2MsBpopmUvJ2BXA8ZiXlZ5jbUKk9IW+KbQHaMzxSUWbS
ZY+15xW3xx5ci1pKxV7p+Kjs1D87MseJ9bx2L8LoaEnGgtwLc8+JTSRmKT+0
sJzUpir7QfD+ZHCS5kcSY0Ot+Bhc7rJb+OYY5dpilUAJH7b/mbJGH09aXtIt
buF/nVGGT7poZ1hFImB7jRcSS+mTKQLq5wacqIJLKhvlh+Zmd5hJFY6uEAC2
yF+wcL73Ve9Krnz0159n00b2UUjWSIDeS55bKcktaSikDf8I6TCZvEbeX8sS
u2ulVfgdsEPae6TgyEKMPiBbS2ts91/noap33RNd891z86vT1cbLMc3vL0tQ
yqRRQZJ0cKJbu80qzF/dCdTxpWG74zJ/e7fXXCLc8xMzQkGqH2wF8IVdJ5PV
P1+SDrs3QvUYMegEfYnZIQ9X+8iGEZ3yXv/IRtoVyenSR5dBk7P6ZE0QEXeK
pxD7AfkLV3qGMZH/CwCDGjMDi2wENy9npFWufzVHQA3FsXZhCVi4St9i/AxJ
6yhHJFHQFtZMZmx15sx8Idfq3Qm5fFuvsnZraq92EbUpg7mIg7fZeD1ZQ2Ce
4m9As4HV04wByYCyUux3HerNNGbTHHQz1IuLhPc1CUbIrW6wkEam6KDTs8bB
UIOGUwXE6sE+zBfuthUaS2/0wDtaX+pTceYZC53VX55ZjP8HJ4/dwxBfFfo/
T6shYv7xQG+SVGEhe8IBgJOqyT82fPP1T4QUISOA/qkQPbdcfz6k/VsnHFnb
8s2jpkTcTW0fsMomCZmKmsJLDSaGBEH07XAAl1w6PCKCoxxBLybxlToP+xij
bINBMmqZL8LXwU7lqoCOaOXK/qmjnhOTD3Bw2W8UFDqSMudvvVffpMmw54HB
RSnFMiwqyK5Y6bQJ506uZvgIMSPo16YxkMGeY3NogfIbDGyNNx/I3EWkF2BU
5MeTPa5YaqaTY3DMPlZ317K/PTADP7rRZnobF6v5k+lnMmnqoYpzy5cG9/Fz
4JtAOSbya1+uwZHCN8NAzncCCaVpsuynngbHxZ8cMMv4IzhqAktTpFTdU5/u
CBK4SZv2Zij0Yac2h2L1bySFwBtB9lXxCIFf2+9yIwP2k61C36sbPQpZxg2t
8PvHr58BF1Z92rHehkNaSWjkRXcuv5IOX29Wgv+3j38uGJcXtvIn3WSWOpDM
uqhgMlHDpNRK1eDi+OLJwgyPDwo1mysr6N7H/kqsUG2EooNy5aBCaaV6kwhh
jBNnp4viAJtQbhWAPR2oLCvsJgssk5wPV9DUeNhH2OIAkPmStlLG+Q+L9e7o
c0/VSUgD+BU0076+4yFyKMn965rCpM+hIiECfp6VzSC+xtP1kep/arnW6NZS
Z338pfk41YDSD+lUzR4gMxGavNPEgtF1INbkVYJb9Y1l3lkgqkiQos5/VdkO
D2vHDoUavPGnLl+ldTQLAdFdhZAZS24NWF7hB6R+IoIFp2+LD3aXUlVWhXC5
TP3ixWeUQwod3pBYPmRD4xjw6QjBv3Hai4bNoZ+k2QYXJdXf3vIPwGIoJa3i
hAmBMag8SdzTeuKxQdlCCAP99aV5A266X4t5AcJgS9S3qGLDapXLGVr1T5oT
KloeHBjDo2H5oZipJx1GbwiZl0fRx+vRcAmD2G/YQyYGainMaYWNDAMZYm/G
w6+hxyR6V5tV8NhImVXZ1LFROp/NcUqsRYt5R6WUl2sFflarhrxBxk7NS/gF
I+0F+g1AobWi2hG+pFUngkhhpq7O10rKbgiZmySZ/rA4elCvltAqEH0kZ+xs
e6bErMeRJC2uBZeeSYWPUFMQB+vpgzciyMdgPbJmCAmOlgt3hepmJ1//TmdG
PhR5HAeKTT6hyTb7F/IkpLw90NjwLtNhwB2MJE859dE5raWP5lPmECaAymon
p5Oelw8uyJSwhSE43X5/mohYlj9TBxhxJUY2AkxdLzVB3fuUdGiTupO+Qirk
VBOBrwNtJqlTnz9bWC2VejXxMWUkZbuERZEaUS8Hrzu7v2K30lWCVKg4K2Yd
v+ZFXqD3puDr4SSiUCEl1kce/JukOpMsccIHQi3ti8fC4s++0akCQB3Cj1bj
3MJS+8IAiKwOkD4WanG+D36FiUwvtFdNny3BzspZaIW1X/pAP2sLWkK05t8e
l52bng9W2qtl03lSY5jaBXfkZne5SbliCzwhlvg8sp7tBnMOTe6xCVbehbwh
hl8Pewfhst43NxLobLD84/e3Fu7Z4z3okmYBS3/Cx3YWLd4OVCSLMc6qJm1N
4z3CFufy9qNrDjcarhdQOeJ86CnfXnriQBtIKCCvT1fVHAty/UqUGizgr5d6
NYttEtdZfGEze27sZ4QC22sEvMZtsLWIOQAeCkK4drioF2+VVFVymXmzoTqc
v2omkRhXWUkjzk0a07GyI1swHlmpJsi+UNXwR0dwawZKmf1SKteT9TbtDUhn
9pa8JlP9HzohnjItsBXpWri40wihKSQ18bpuh6w/1Cx/SnoM+RzFfMa7VsTG
UsunPFq3FGd24ItenAIbPG3otIQwvpyOvvezFj288WA+83dl54bM/GF5I674
cYH5o92QFyGpjc8HuevMn9TtmSUcL43tZJc+KnY1yfyrUSIpMYyWKVKdVCrJ
OEC+bpVWI+6CdC3gsdKqk/d5Nv2qC2AHJdkYJGYFlq5DVfGfum7Z64fya4Pz
l2dZt7Kz9Pz66KT2MytF5lQswacMSGu3bDXr0qOr9A0s95xCeluj//eilcsK
nF7TIl7mc7sXmU5aSHfiV0sLloWSQfcU2/Ab7GH6Vg/k/dZTwuNUWlYf93Dt
y6qTAnPMd96VV2lizR+iORUGfVPhEQYn/9iDdwUF+U9rnEDKYOhU7dnVYAdw
s4n4YGRN0VB+6N2KC3nJRV4fL47IebIdYhA5/uLzkgVZxmLvSa8wbec4sgfq
EB1IMYcHSV6Fe6MDghYnJUkxEfDW6muHD4GHXHqmSDofp76UGhn2IYhzSIWf
wcgztFiLuiB63i/DTt8+JxTYYLJC7c36wYRPDWN5mnxxH/ddJsa6HXmCKmMp
Z5uHQYksnZd0HdThw3ygjIwA7eAQQgwRqQmuwu1C2+hIs8HMb/0lny0dzgMq
oLHMvckTasBzTUnpndJ3Si4Tk3UmL7Fx0gLP6Nqxqqv8juuk7Ey/der4nHiV
HXWmw576c3AEDzIw23oDKSom8rNYawdYduf3phEHATeSE4ajYjmV54eYkCAK
Oqz7bGvVGBtkw4Gh+DMcxOPB8k9mGro7rk9nks/4Bp3JYjHr1+30gEwr7zh3
jIZUr97GPaV2u71cEXzG9G91ZxhLK6vPRrDXNgcU7IfteUDNabCCWDFwY7i8
hTnzwjc8jS73eutSZdXR179bfbILiNX7UcmgTj4qk8VkVSvqCQj/vIclg1nm
WAFa1prnDDSCtHcWLA7UHKprS0hvzJG1z/IaksqpTz9l2rXedG8RxAOg0w7p
NW/S/3UgnNHOB9/kvmKXkeRbd2fet44o4w0Lokv1J8KTTqbS7DInMTZ+kPSH
Uezrs/57w+pPu87TnZzuHwmerj0yvENjJ2t0Oxr5iPPp5ovTVPiRaiPU6U3t
KSiJOBMq9SlM4ADr/s9L/O3LntSQO0TCGAPJTb9b+XtOcxxA36obkUFz+CfE
cqO/5202RKa4qEeMyQiCFH+stU/sboODp2zXA/QYQK7yOC1j+c4QVQjzVf3O
M2DsI/KER8VPZpXrVK6zrB1Ae9EUp2LhUeFfdXIr82k0xoLEqZwo8vogWwZQ
D8pzZKVYpc3HuVkNuBXax+A50dB8KFwKosnhgtTXB2smfEcjkR+DBF1sj099
Cut+bw8i/vVzvAMnIzU5HjiPTDW1jUEAdg3XtRwKJ1NVywJYeXpwuceJ9WqQ
Pkb2og8eqS9Gm3NP1AN9TWmEkTtLdM6L2K6h9MRy+ztQKPJIe9hjMp4vZL1n
HqYee2N1JwXQpS0/F7dHEj/GDNZjIpEepMwcIHFv6pk+hEmNGensTCYQk6L9
xP/6aVCXaHVRHhK6pcRDSj4DapJMG4ukQq/GcDkcpvgRw0dEB9VqBHFFTxMH
Pu/+gV19d4j7RA5Zf9q3e+egOm7j95NXP00q0xDaqcuG1WaWMB3zqXoau9Q3
oIHyCMfCBeGrw5AgXZ7GApoUH0tg/bYD3QqCJ9HY//AuILx6e/myyQNspBta
XZn3ok4id76q6b/+WwTaVch4V765L+W71c6ZcEJhwpo/5HJop7zJhKszgIY3
40lESHOTWl7PjiugAe275jPcZuSeHvyWDDyRAtzCZC1Xm3NhgKxzS4ZN451j
U9SisIh8VeS9vX95ZLeJKgJNnvPn5ADUf7We3DNZM1o+3RRd0U2q7mLbftM5
/OW1rW8Td2ZF6zW7NPJSfxjB/kmvHPXLTSgIhmORWjGiqmHJd+HFCcmcp7T3
wLZ5OCIZM3S1Ob2s5CDovWIH+EX4DKoNT85zV4gD1/dxmCzudvhLKPN6hTK+
kCq6KvvQL5e/MRn5CgPzkgYGxnD9NclaxDK1kkF0M8IIlINSLqjtwh7vpJXE
qMWLm9wNbcYP7md/S2+KsMNRQ9m8MEwzNpeY6rZfTvngY/z0I9OqTdFBKH0L
ts5jSfGqFyhFQ9xjLet7Y4C5G2HJi9O2szDsNN4odam3w0GE6QMh2hYMjcjq
x4z7E8owUPDQ3OU2796h91OEgLMYMmV2niqw0DCqPJUIdLRC6inL1rYgHT6u
1csUEfYtrt7LUy3VHCW88+hSuNoxGyjn/b0uQGIDdc7BFVxODGbjS1SJAtTC
efPaA+HCx3BbTkaprFECC1WJ7SI7R++8UlDqMGLaL6DWpx46T9Fjkt8ZQIvF
Bxn3nvJJtq/Xv9Bxd2F+CDguDAOjpclrWHHeDJkwjyF2MWKK/L90YkrHH1wi
64RhhGRfKFzCEg28kzGA0cNG5TTjIz89QILwKwKMYloij7N0FSORo2n2MJgx
EOZ6Yd4WG6O7WfZGKuZXfKgZLKuggdH15TNCiQpBTzfplQn2EUb31B3nbtMJ
UBdscr9qi6uJCzKmz6B8uKLlQo7Xxr8DERfsy4LyogU7WgALcZ2Zo1G6P+1v
QrWeiKV/7PJr5Xa50813asy2RU29QdlztORHEBThwO3fo/Zpg8qnCgFKK6AP
sFJ0ZyqDvp6Q3DzZLpuAvXibRlBd7qkvc98upPHuEim5TMY07FmFcdJ//rpA
z9ttLwegmC8SYAIOMFKqeo1y/T2imyDDgIEbelUl7mM/bKx2SGuOh03YDjqO
yHGcA1E6849/QF6UdRvlHUSpBVutC4gmg4FmpwEq7btrLai+n7cX6M2ghy3c
QrIp47pBwFBOSYAtEZ/mKhnJzV/VDpWDQL6n5aXxgCRW8u29AUoKuq1jXxG7
ETdGS8FwjV33T+wDfM3g+MM8aXFlbb7zNQDyz+eheyUUgasR0G0QMeMvK4jH
bLok6mew8BbVdzNfw+twXAeS2cWmlCxFwwbkb3VK6ahSA+O5bxi01h4Hkqc3
XpVS3roJ+bgAvQYt4gubBuni6fUP6sUdKyT6RVTCI0BZra7iDIyLbXvmVqgl
1ONvm/rW4eWDU651UA34VL5XQIqoVmq0RxHM9WJTsX2iL5i5yC5sAV94BMf8
5MSAi/60RBQlMeIzlnnEetNnAMsXTCeCZtuk/EowbNLMkQpy+2tvRndbX99Z
m28YzW6du0uTkEYkJFiSoQTWLJkxQE8sSLAO5relpdpkClEMfSp6NA4ULVqD
Ic/SNWy4yL1lEitXXsLvCzJMMIXarGddZVQdOFURYblgy9ws9NbnD9Q9FTxh
Ywx9Q99LY3nBLuq4P5Q46u+ZRD4oIZbK0PO0WX1JUDvniia/B1HTgFnW9Jya
LRPhpVniKcyBTN/zK4hMTMV0kDKs1S5WJQwNp/STk+HLIAJYcMRxkB3F0NCv
l/7fXuNhalbWFfPvEW3J+DwSYKbrXniZlSgNLa1Vqlf88FciKl1D2iAXT3Jj
GbjW9BcCtRXFIsfM9djKVIP7jlncdjU3ahjUkAyfbnnM52IzxA5UMO3mZ3lU
vaFxKIKoIqNt0vnG9w6DnOo8KoMJBeUhKszPuXDNRAktHPV+vF81qMtPOKkM
nm07mqv43gzElDqsxnwYdajaPMtlBHu7GuuWfH8WA3YsN/l8ohMsXGG3ZqFV
Px6vT9kQlZ3pgy7iFCmIDYAz+J+IN9EmWHU+9Tn7cooI2nF/sQIpzJQy2MVB
IHss/HLe8gXnownA/vMKnyWQSIt9ZiHG2m32SRE9xNhKL+RWkSPlbFh7wPoC
OPlqnB/InFZH0pYoccOBi21pyo/zcpnSicibJ+ZsD96PCpWnzZNbd1yJ/LIU
rjKOl/Z4fgbwkftpeSZ8z0G72Q/JJu2gPjs1zlGfFs0uXX8fdmaXNXN1aSX6
W3CIHW6NBHfdOyXVl+BTvpkCjvFgGVYp+1qDeEuUaiu8cfzr46e+DbCxVLMt
Q6pCFzH3Yr0irmuTray43iTPuaxy6hkWTVcpFjzMCghiZ1S5W/DszJojFFC0
EjHeLgW8WWuXtN3VIh2GRcguHsNlfHvULNCf2YpS/fSdsEbbEnIXFIsT6/gC
9QZASvjcm1z/BH57KB2SsHuvK6giUWDOuivWVAVpQDvguTTa3JgL0Kptt8wS
HSra3qxl45AU3cfHcuKb5ocugrbyqEax9FgAybRzgrruKJo5+DXR7XXo2iQs
TmLmQIzpjE1he6UnyF3C1NTxwvwyDvItk+xzS/RPCnYSSkJLzrJTfSatXGpY
lU7RfvGzStIDjBT7LIiRsa6DyV+F91ZQF9V3GTn+oUTFeVQvWPGkOh6xOIQs
LNYFrR1TjRPHpUWwDJHluRJAtmcWXUkq/pUmF9mDLjIbNVV0Vp7TIwl4xW5V
EKfbbOkTaFyAsFTdLPM3CGcpl+occzCAsoA2hJePjBA1p9C8Rf9cxCzCO46T
FD06vWa3+wIB3FjgC84srwRyuYut+Eth1fyrSGvNyz70b6BpIVKjhsmbcHwI
VTZ68DXFIpyg/6toUrWhou5Xfy4368gUHhYmJJAFnPtWQh1AbMUyOtUkUlja
ZcxTalSs7sbaDXp2haXz8JLIXnG4nop1pBYUsPq0UMhLnxzQqgyr3b+YQ71b
HGwQHVETYWXeRcLkcPA2mNvfpQx9wo3PDQ9tnRyD0EzsMAAploObGbJVGNuN
q9L/KO7y6LnBSZBViEVzb1hW8d7EcN98aHAkoUDiMR/64dnmlIyngfEsgksK
UnZxVdJAO9tHRt+FalA1q30GGHZKah7oNKvCrhEmvnL+cxQ36Ek2bpEOVT8P
5jXbpP68gmW6cFN7Sh915riRiWNmrPGDznOBt1HCqOXGHCnS8Z+RbNo2Ekp6
83n4Umu+LE8yZV0fyR5WgnJcrBAl5bQe+lJytaVg/WGQ5Ts0oK4zH5VUA7NF
K7gqUAgopl5J4dQaItr44FqzfQNUIvcieTfPz7NH4t02fvtwa95alvr7CXTC
qQlLNQUV4A6Zvq6eQqXSFDCO/+DFP5im5fTlZksKOnHm6rKLvtAL99qXo4Cw
y1dLnSpSH2ICWasW7o79qltj0Rvb9T5vyPGE8twIHWYbuJcHOT9kC8ncK82i
2a6O0pGT86zWrBqR8K1aUq5tCywLiUVIP9+DSotMHSk6JenyrFRX6ZOgU/GP
0sAZV2esvzBbChpvfDjewplligStfxAV6lmFIBS6NXL4NwVy0yVtNxfpz1Se
8JIxG/Dea8HgGyMeo2HnqGL9GVhiQoCjtFKTKhzFQ0HvVNVgKCjADYz8QA1X
HXmTsPa1toVd2i2vvDaqOSTmHN9mmtpn06MQRhY+TuYCu5tC9KuU4TAfptT4
jHvFmle01YDcWIwocA+lRmxFv3DZyPF6OFALkqIm+qN/9ooB8SC2o5EzMoIv
i67jZgP7ueIYx6olKQmaks6LLTE8HnIUvyu0cfmpoB2i5ZMilVsrYYuuDpQ2
uZ6SFyaEWo6HoqSNyjQzT4YA+asSVmrTojD1mmXftErUosDow6DD1kV8bFAu
MSiMIRtMyWX78lhV53BpoWy41G5VLuhl+y5hHm9tLbE3xOW4CQfnmbQIup7c
qYnR6IuU9UCkwELUTiGPpTQEs8rTM5bifNKxTQfbD7n3ar/HKxVp9k5lNrZg
hhIn1y8H4AMcjK2pAT/Gc3Kh/eb+Ld3uKP/x89w+mJ7agLu5DawdYZwQdjkB
Sd8sqSZP3ZKObu2aNeEevhlPODi9Q5rPsh1+QRnn3KtqMZv8TQcy52GsxvZC
BmtHTV9rdmF4hpF2LfOSjIFsNpX1ycfK/KRb5DO5kKSS5kz3PYXob0ke1mP9
ltsdY8nPMnnUBAmopbV0gyynE6HHgWTdn9Maf6cmRc44JCGpyyCERthCL8Ru
tdh9/bHmuX3WZnMawu7c0l204hGDO+m/irlmMn5B9QVR484FFkM+1JQMMCTk
GyPuy1QroG3HFDZkJtTz1u+m90vgVUeMOPtCPLcgur4mPac9lujMzoEFDsLV
p7q8/tJWhsCWtSaFOusmMX8fW2tDggDWuD9Q28Q4Aty+axPMVm8h791CGm0x
V4l+FOwR4pFsSdeo+I98cxBSIiEzsI41V0OOI9RlEt6NhqXYWNaIO81yZBmS
OQsK503s2NdY+QWmgBsddAk0PLOJYOiL2MzuadMPEP6AHCZf/3nE4TQD0BG2
VLq3n5FFm7O02RSgqvrSJfRuFGakAfCo7NbYVzW+zcif8NTgJKpQvRBuA1QG
NrqYMzRKvt8dhCf0bEYbRcJSYTaXGQYfmDNh0SUaiX0YJ3gwmL5tE7xQGBa/
gCijO69CYJpzZTPoVdxxgEHzW7YASONIotHjI75iUKC/XmyOeyRCrTJC4YSw
F9mOwgPqJlyVY+FCPpzuocqnO3lAU3Hh9d8ZW1qDZHiSrhhdcp+Z3oSArmyM
cY5Fc0TRTxbpPQPT0uRZAdUK1oG199fCvRnlW1M/Mm9qI004U2vrrUUr0PIj
3K5aVTCtvwSndbAG65+DkCUmoHS+J8fWQzhC+N3cqrDkSXNz4b5IQ6Hn8Hk4
uyFMsWdMJRibg1A+OAGMNnqXClfGNQkcDj4V0L5y3TBZuFR/qX1PQJIN5FZE
T7a1PgeXuBpScypdfAH7gy7jYf9W3ORe81qro2R0X4QFLP5ZqLiuQP8SMaep
JwMZn6mfTJHdrHqNcmsz+8HEFuk30uV3+aq/YcToZ7UeqCstlgR3dyO0RN02
M1guVl3/F6bk6k7SiFAzp4ZIx7BPojIp6zglHQsJcLrbSuI6Pdj7cl+D3rD0
RskLEw3d0IPk5bY4/QPCV0D0cCW2ho8ngkwaM45sAVJ7360EYEsRc9nGBkPY
JO2KqPwZ06SJ2qSntMWhdl/pnm4olOFTdDlULULFn0wsw58zDjfcVaHwY627
/QzIFJya86Pn5buUGfBxUzHXb3xI0LKgCaW3fHg3/QXAStQgsVg+YCC9zayC
9fBJGOTKGWLsn1bHwuOmpivwN9RRk6HdriqWoUrwZByzbnDST526CwhDHuaZ
G+Row7b964+TENW9tZrU9R+aCPFZ4fqzfmtjUNShkK93uEGz/i/EyuYR5KLL
9XrbtbRljYhsUnV9pioTkhJ2hzCOqJqqgYEmAwsRgWrQn6/cUXFAyvUfE2oo
YWVyUYvyG6JebDK+JkgGGWKZiRPX8MFcy5ohOX5uU5ffrlPLQndIX7tDqqk7
Ibush6QgjO8JPk41ewvXjcZe7lA6ttU5f0ogHt34LFWeetP9emBW3Tg/rIZ3
fwTa44OaV0kTvjQgBSnPdRwRSZHIW/cS3amcbjIAlPoAJblJjR5GkJwhVt2b
HPCulFQAJKAJIZ7nvk+dxFO0mHU15r7PPPDrr5i1kBETPAKWRYi0Yv4WIlti
pUyTB088yEsTtkkUPNIP6Uow0G4ZDCIcwTpXhP7+CLv6w/6CoOtGwLZaQtlK
1i/c6I6BpMnxSC6+WUzODzYBvrnieZ5W1TfKP6kxGkIdbXQ+JyXZUdDzxkJn
/gLXxWYMlIYFbzUGPPt8obhTz82sLDzUNz0sfXrlH+xz+huCIb8G6ItAARg4
VEG8Ep9m1b9dElG+0ExWZC80IEZV8mo8OyvXFDckVwGefTm9830edyvAsp0n
yCZgj4/un0OjjHKUQNGTKTSw4/NAVJAkjav5h3jThsHOaGnC6N8vFb4oK+2u
DC0l7g0WlESKk3QP3dDCy09w8IMI70WuMN4TX1dXoT2B0pvXcgMTQ8wfpLrq
D4ETGIWlzfXe55eXjjwtbpMBNerzR89vCT9eJSeAg47nGY32Tj8VZMo3VeSi
B8RaPeHUrOU1U/4sYSvqfyS5E0IziW75mUhCBzsH3sCAlAgULtECb78mONmx
7KkhyaKxKxnXThRDOICep/cEIhKksnHSA+TvnpoWGhpM/Y5+onQNqBxsa0X/
7E9BdSC0NdXX6JvVpJ3vDEUAOmJpFpcHHs9x2iPaumWfn6TTN4eBBQt5Xvee
tpT28pZ4FHZpOF6fiCu0nEKCO1i3L1j+712Uzvi5/u9J3DQnI7AqYufbQGAQ
fOSznYy51y5GnUihcNic8qdCul7EOgFMSznDbTlIrRMs63RnXMm2Y+WkPRq4
87Y7xyfIP0OjW4taM+jH5jBKk8ATbsTjCwTm8EdN1r/fKbZjzOO8EsoKPh2I
DcbQ9hx6Sz85lcxU2+91iyic1KzNbuvgggdRQ+N7KoM6E5aQ5Cku1/CI2gig
fvV1ardvhf8Od/rXIi+N3wILFV8BtZt98UO40xCEPBcYtpPI3T6ScmaBvcDz
UEQEpYLe6flE5xj1mpoV9Gi/nBFQZy81jc0YNMTQkmfea+Gn2FY46kaaRxCX
sSaY0up52Q3LS8BG4eWSpMaijYI7d0zRm21ZcUBxV7Y5eMII7I3Tr9vE8oF6
iR/3kNxGjoGSkuRzhZWNCdelpYgc0bkOevu9tcky/sTfwoEDwqWkWOs3jv63
thAVcaFly0un/5pzNcImZ+R5/TEiLA/qaHX9Dahir6SCKbM+zuECvHvigMhG
u4EwImiJVBlY0dKnWFM7BuAIZqYCMJ9IcD0Gvv5oW66GdRT0JqzcDCcUp0Fj
Cy1bQsV/PeuHzOZgl9QsazEP4oHk3EZUcTJ2MfLJNigMfacQuhVAZARChSUE
ibPMhr4AepPplA+ynr1AfItbzLhEYSGwjxBurHtecqdwwrSsSXgktiwon8zs
vvcf+LqN5VeqiEox8KJ2RFxxacq4i0tkil5xy6btGQZ4aN1M1KzwP2srx29t
fceeIAQmBgqNww1qOB6dSYQq52Z63cMFHxT8sETeQbKAPuXssEsmb2NQfT5x
+dJAusM7JNSjDqTamcGZHstU6FADqgd1Cprh0Ydp9H3fcE412/r7fThXSpjq
7hp85zoGnq7Updhgp48TOVl2N54oeg5SwhL+1VUWGEPVPvTEI52G5E4Brs+w
HC8vpWYOWlIjCGp4QMekIW/Ru1dJ4HuigiQPMU9sMEa+XSd7BGV4hLnxbjyl
GiYyk9QqLJAFkwDOJRDjHrX3RbgkNSpxWgBt7KYKhCI++NmSUqC7/ljfK+y1
YIi1828kBJJi5/7zGUzADjeIaM8CXi3nKQR6mTVKf56v5q7RWux0xY5yd7t/
RrFFVArO8hqvvj8qAkZ1xMRfdeX6nQBhr9dHQRT064UMfuHS9v3+KfasI4q+
QSCKGPMo1SlY2S2nD4C0k8EC2117Hq6vSaS2yMjY0toeFzZFZw5YD6QW3jkJ
D7tjs31zL9miaa4+wd0NqGH0hUo1klH2+pPqEqsm8vr7elr6PibdiaKlt0h6
DfMW7M3srpigJr83GDhm9QldRV/K/+BzPrptirT9iG1gys/X6hz7iRTnnY5u
OyS+yUaWf7r2iBkLDKq+nIwl//Lft86oVghXwMfcNcdX6QinS4Ict94NOD5d
A/vp35HlB2OLkLAmw+LvGvxaJXTaFVUtF4EUsd57LHB61YfJWcG64SDWkky9
14HD7vs/RFcaPLteHF0bqQA0OBoRRnjLjikGP43wqA8cjGNUVvUfduGPdyQu
IqqSWlTcAT9Ornfp+YrGAwmMDD42Ru0FU6pmmNfIIzsGjMLlrJuSBn5vaj1r
UHjc8l3OzPzH5PhR0DsYLBdcu0ioiJ24e25EpO+SD+afeWtdbYSezsi6dhb/
+FRcIVJWJNhcdRJ1GWF1ZWmQwQ5xoUm0giQyg8Y4LjlNtWP653x9y72eFfnd
eHAu8bV5nv/4q33AZPP4zgn7RGkxzF7C0GWPUjMDtJDG6sBcH7xNiYBlJOX3
8420Y6Nmi6mSd8CW2m0wJJGrz0kzDL+0WqvCPAGm0krn+Dj4Kpd9pa6NiLLg
MwJJNXTJZ1ztuX34VapQ/auqgqEO37dzRjZ9UgiKJmjYvfzuc5vuYUKIJo2v
3x126wZzG4YD1LlclJSq1S0VdCXqvDZcIR3eJeI9q1ymiOrlP9gRq0TT1TYY
zSBqjmf4nUw+TRNlnbqxXgm2OuJyQwlR5jLcauVtgKwVu01rE8MW/FF4Eps6
VN9FK9xrpAEt8nlzqb9mszKNDY5UO97CPS06hvEUH9ppfeKLZ6BcFh6Oq+Jp
tBA/oCoDtJbvyr3QIUZSHFlvYufMqCgkBSZ7EX9x2xCtIdDV5pW+vYHSbOrg
eF+ZpocSq8vhvKXQ1Qzmed3Y19XlKhhcnI9Oag8DBjvaF1YeomRRKDbMidUK
nWGwIHOCreVKN5uP8GrSMI/jpy6jHNsZflcSz20TIEc8yMRpC4nwPT60jWWO
eX9qgpFuipm9fhqJW3fi1KSTHPRFYISKcEISEd/fV3aLQ/6wF+oWd/hT8Fo2
fcQC4Q6WnZWr17Q7UO4mT0IFYL3valYhYsD2c6EovGUQuYG1eOsHVxpT+12+
GT8YvQ/fSwB1iyNUB4hsw2sL2z7LsMjRZsZxEHPeHXWmPJE25mw2TpJnVBXe
G3sJix5PC+NVa1pwayyewFrZqfa5O+Y988B/lA78BN2R6Ky94fYpeRf7z9p0
+4/0HHPKrQfOqs0z3U2fvpeGzrpgxCKwIvdvtGyuXeOaFScjhRLEponpHFAN
9aoGC5HiZGfXQNyAkKabQpjbhaZO8GtfscvyG+BsQBgohgLxgo74xOOQVrew
bBxp85X8FsZAEmQQ6mCsXsHlyTXLphL4WBkj4/1f4zu51y9GtFlIsv3RTovB
RnpRlsEdQKNccoNSvTPYlp5gq+va1ITRRe1U/zLO0mUA0voxLEuDd3zWDYDa
Oh9vD8cq+QKVNfWp4NJAbQ6SRQkbnDlDN0D7sJ83fcTdlinkD/jbAyDT07gL
s0sz1rdVMxms2sBpj3l5/yNWD2ZVzDmwwu3NF3Da+70YYo1YNnwskbimD0xU
OVJ9RXqKsVb6PHEOEbCFPTx/8kwH+SmkRG/hPcy0e4qxsq4mJLkBOEvdu7N6
OsAUW96K2ZF6+t8w1yPVxx90tgRJqw3riwrjTr49rLY3jkNJSQsoZWGAHvh6
UHSedEc6rrQhjNmJlB1roMm5T9DbU8bzMY0v/tbkDsw1zJLkX1qgr88Bw3aX
wVg/8aqVZV1dGV3pLMSkO2mBjK8rODLsfwJGJmMXGXkgxeBEogoSVS7fD9D1
PUL81GYdu16g3iinxpEuaoIzqGkruhEAs+EK5WjJ40IW9bfqAUkpbrPNwVtp
P4e8miRQO6hafJtzohwHaphQShH51AvD7dwdY7+5JWWg0Exeg9eF7AkvfCPA
2hLh3HK+Gg+ihsS2f8TQDJb0WVJB+rCodC/SwVXtqaV3OeFScfq7L4FPLkD/
YZes/FxiymkoxEvnPzxE92S1AKA7gf14wa3tX/RJWU6h/ljIVLCkx1HPgh6m
tpvKQtkyF75irANGOn4QVdHrmD2VyqvBmKKfhpdsrnEGWRz7mJCVrMNRHTPY
xsEvhZ00pVf0E6tGXhcW8i1eFyMq5AyC8l3u4UeKX0OeXEUC1eT1DcxCWB4e
cka0RZHAELwpdvb86tUHkgG7fPkGJ8wncb4na5HTPQUX54Ru60HzTVQzHzFv
CQ0fOEm4D+0ofurtYKmqUXnLzmH48QqhryN8t+aCuHjS6E//jo2oEFr7CTDY
msoTwGoNxH94gdV948iLfJQLNSn5dzUkeE9LANaqPdGsEtLZ9Q96680p4SWN
cBHnnRtC7rxp+yxQDgjxvD0G2+YV/pcyKzvrrbpgY0CxW/CP0bYpNhHP4W3M
3T5A291MWbcvIuw2nlQuZVCKm5JznIx21bmpugJzjoKHQGI8GAsWCHSJsi21
BAo3Neuk3CsN6mmMVspNRxf2PI0sTSzFpq6pwjXsF1uejz6tiKlhi/uJWK5S
/y7H/TWA8lAFt2YOTY2NRZ1fP8hvB6i2TGv6+f4TBRuZUnFCJP5IiOcmAcLH
sgqDNdJrPcoZrdCXNBwR2MZX3jILQHjUbPdjZkIJFmp1gOWhIjp4QfZDJxp/
aLuhogmNIilUB0jtcUkgtmZIoE/x6NbsU6RXysxKlosUXwTavLfQUHXzYalu
J3mUzsEJvMl9qGqGD7N/qdFTSElp9h4Bb/Z7Metx57ZV7ASsJKpYthf1UMmi
KsMcqX3O8UHNdL+h0jsaK9gISKzQU+QcSyFNAoA+hSsDh7BrGxjm8TJMAD19
rdH/VUcBTOh1P7e5yacYmtU6J5pEq5xahlhcEFR29zm11tbsCMRlYwaWRDui
DjXKt3GoTRxmQeGcovSgBKFQ0o11pis+IEsYO0FqzgicqnsTms9P0zrf3G7C
p+Eiz+OM1as2hJAXIVPVn5Ch2QYvP+D7EvyrdyDI3FzIAw6hff0RF6jRwTO7
hEMWMa0/YsXGRE3liqkGhRNSB8WbnuFc4Ztn1idN6LXHmhBxF+6sGt+HrwCr
mMsrNBGsyKIejAQyAdEEbQjeQ/Lo8+AeV7EPgSlzprWaFm5kGlp6kM8+lLYp
W8R3CPFfUSZR76SflJWqp/nVMu8SZESMife/B+jHBBM61FBYX33y39/en6SO
76GQPMTuoX96wsG5V87ALTODRdm8aIwlt1wN1lftptNBZVrQejKnmjKnsGGJ
uhJTqA/37F9KvYsOT4PRA7fruh6vQbNb3/NpQvT8kH9OPWg/8f2snNjO0dAC
zFEr+RWtzKK+uBaRlrv+dvLAzMSpQ0AScTjEmJs5OfQR+L1H9+79NYxDA3D0
Qw9BrHjhjuFBSY9ENp5+TcCFBFFJ58qxg8RtrTfqtS8x+Yf4IoOcCUzDHKjg
D9di1NjnGlsHXW53l8w68aeK4HNMcjUiqRrNWZjN3z4M4YA+rgn4c/G7xLsv
JzEScjgMvKluJkFNhlc1NKICrbbxeH6neoxT/ZTsI+RM9erTFuTBH6PYCFQF
72wMjC0iX7BAnyu8tKx8DOI96YAclYHLvr1FcC//aa/kJKbGhdMaTJqTTyrZ
uYzpnmDQRS+LyCYByecd8Q4aTsLb4tisUyh8qmfeo5puuf4ItI09ioxamkzl
xTKEfAof1rJp+myyVvZ9Q6nQxqjLA6NHYsTY2MiiWzQO3MUbAZk7cZq0sdja
JOcjaFSr5dHgi0g2OKoXkMKLbt+LMxwad/R26kodqHEOSv187OaVJjmjOAZB
t/9zjG2xU7wbUSpoyMtEeybNP3aI6nlqRsDfMSSph/0KCDu/gYM8ShO+m/WZ
QcwCCFcDgDjZxIXHYvba10HxLHVhZ8QWFoPMMbiUa2Iy7GsXa1M/MgkKyCb3
vmU0YnZnff3EIgY1GI11JddtW9nDUNGe+BKDQXQWsRk74B4XfOS4cW4aP1kV
grqh+3W7FItcsJuqtSjnYCVAT16mO137rZhkQBRe2qnqGf13jIx5hcsvimgZ
D4jcYI4y5rZshuvoA2TFjHT0JIqwcmJ8EGPBgnU4w0eJNBOPahHmBFZbfBJC
PNUcYm0X5zoKEaieVbLwp7XXUTLKyDVczv6YXVSRNF3XTTq0u3e/Ha9yrKT4
Kd68ox/fy4oyh7AzIH8hEShO/K+zy5+ShlZvLD2Kj+PE3Edf3Kt2wj+zw4fs
IRiZ0g9t6J3q0/JYRZIaI1heIU6eUsJ9iglWd93bllhmgV8exuZvmj0/ZaVw
uOTfgBsyXTRZA+xYljoGpIzh0EGBNzdiqtyrPpauKvdbY4z1febZeALhUakL
dgrLwGsDJQucQojsCMQurD/tdlNzQ8yspWM+rFoZ0IhwiWOYcNRD8bqmszOO
ChP5lfEdXNZ+aT6TBjDaURnKx7okLDE2tjhOXP1jKoMGRvSwjh4VKtAL0/vd
qRTYI+tE8LxF6M7Di+PpC8nbCebWFXhiETAusWzzoO/PPrM1KNFrIFuQmJx0
yE8PykKCnszyrTjfyIZh8Byh5RBMXhTt3wJPcpvfiPa7xOGKIS8f3uPBFMco
uHVFGf6rE+doXtVksVqFRz1fY99n2Ja/uNV+hXHAoNyVBfIs15IvQm1GIGTY
2wcXZAib7isOLqLcBiO0cAgkyNLZkATz5mMQauaYBQMBD49PIeSFtq1U6+eA
zzkTp9buJwjSU/0zURsCloGdHvm3q+7MM8VmiTI2cliGLvgTAg/4BRTrCLSo
Lnq315KeWyHudvqFnOz3LP2QE4qkznY3Der9iOBA2B8V87vOQI6apLx9g9+Y
L6x2sLRgxwvDihzh1kVfVmbmDuUDJICdjuvv2hoxpug3+I2VI4wQAKEzsBO1
x9Oq0RVa3E9FUjbw5VmSeQuxovHIF0UmpXS1mjHRMrymrcIARTF88t6ixtUs
q1YA12B4jgbvIITJUxAmbRG+WKXBx99e3g5c5VauzgQ2/mWYQLBUC1WVFaet
jHVtcAqigprWSmL+hquz+/Ad0Sa35zUwOPk8dRYJB0S4SdT0Y3Uxj4vBQy4x
oJZ+5FWM7iaA0dNRk5Q0Tuoq7+42I9oHRqq1HdU3hec+kG7BGf1KiRpJwzrp
3+a3AAbxb4UAm8lVCqm3qLy0LCXJlQtjjtqNcif1QlN4PCdpUHZMq3L9SItu
4s1zjl9/StfmuOr+3meJwRBr/IeXi/kReCB0eVnqmg1VqDt1JnHveyee/B++
orAwEYVpVe5ZNbWb5OtrdbJ1HsypV+cxNL8S7nMheEF8CVketV+9aVAiSbDu
FBSxHb93RtxEWlLmM/Ma1UpMD7VI4mbT9h7fMDsgYQej7Dl8eYcw97zZYkbt
Obfm6SBdJUD2+IdMLJ6ee2JG5LUzEVhUbXc9rUnLBPcuwGsdU3Ac1VHtmofd
/pdsTirdn9UUHGGx0VAmWWs+ROT9DMHr4MtFDE6qhsApml8spcPPijTdXeeo
ENvRe8Y3P68jn4HQlh0isMXbtkIn2jGY5O6ZwMrJAOhLmYoj2XtSZiZi57+a
9t+ckU4129b8g550Aer7NKpUY5SFe9OLk7UVWeDWLn5TsjsEEbM/Htc/YC7l
z9D0KI/IcUhORttad1j31xM+4C//Kdyyra2zQTzc8BLQOmhigXGztXYnparC
qvAUC2esmxYIyIj11Ek3/IVO1FEvC93FJ2DMVI6kBPm9+Peg8C5yuh05hZmX
b3sXAq1rRMyElrKu3GuenTO4LriDKP1LG9Zq8b7h5BCZd3MGByft054oecS5
1DtQUbptTe8UHTs/NAEnxSL6+rYGA4nBsYmvwkc/Uqe0X/HnOe4hKzl3rVoy
Isx9euSAhZfMcc3h2nkbrimLWeQzxbQJHD7aGgmljxAfBiTSxx108CW+lNdF
E63yX3rEt9UIMascUnjWrAQKhA+BUrg2lfMUa5VP7cTFUwyoxCSYKM5lEUbx
bnxEOIl7DrQ6zBxBqurnD1uPCT99LepxGEZsv1+9yGBrEUSf6smAG1EB2bFB
DLFyLN7/OzB1D9DFUVzTYmkp0RHCSt2kFcTXcD7QBjIME7asmTfCT3+CJPAH
+vQpMtk1VtaLUpyxFZbEzVWaRKiYxeU6zpg/nWB8ltXIvfForRoV2oADStjY
6mUBnMq501Gubdc3uXy0k2Udq3VK6FBmbR8Nt2Lha2dcdHC60wiaz7VVcWiS
D4jECvatv5f5hC6RSiQ4+3kZccJaDsQccd+ZzZqRPr/sG/dVCCSdnsMYgI07
pb/+gCcn7mPfvjWJAhx36adUQj248wUQE/TzGr51cyoqsOjEkoPQ0lYezJ3f
D4zWeiA9dvOPea48RtHorcFmoiU7WgxciQ9HseKDpiaIhx8osGxabdUX3Z+h
/82qD7kR3b6Y0iRUCmYih7hOfJebx7FOE9a2eLkpDQwUMyBYsGh2XJZ8B+/C
bTj1mnpN993cI9rNBBpdQrnX1ZhzvQCq1jXVYkWkJjD/v/N/MneuskfQl7hy
JXgGtBdQt1FhPRYaTatFpEd1gKODn2iPbkEQKt//JNukegGzitKLGmCJ/Srg
j7uIi6xDsT2YRlNy2zXI5MthUeSHCoaANV4FlSPkkKc5EIYgD8PQhJSHDhKn
fSPqFi7g+tAH6sV7NW8BV9xddYRA9m5/qZ7h52kJPLNmszqAc2Lc+mf81agD
bv2bR9IPvs/p2wTudgzLfACh1HGd7Qi/rtRNLmWS4HF5U6FPHuChJkW62b9V
C70kN1XcXgOVEKUtbYs6Y6Gf3FAWRBxkGda78NNwnWAEZm4oQAl3wXdmNxhd
6OKq9oJqp4iAwZD0+jsy/dw58fIAUuCpA4Td43dqrCvyw7LqKnP6LcWxpdpL
UA1z2ObemCovMXU+IQMTsVZThEnsMzAObyvsCcNEm3uSC76EIXGEhkCWX/N2
d1qlLPB9c0FI7jeOcAvi/m5rtVy+DZ4BFC0pHQATO47YfKvOSJ8sXLbrSjk/
9HSjCb6+Eq3JzP45wqmRwxMtiuynzKM9au0/3XNFCnE1iuzCKY/Pcz54yCzK
/6MB5e+GSClrrHdiJOgn4x7GifGX3vQ3XF1acL75GkTTIKXFQx37kXsjmM7h
gxT6VEYsnRpuohCYiTFMIRDo2kjHAaJfCuJQyu6zrjge7ET5++OaGWF8sl1O
gmKGxQVvXDqzQHX/JHE4c7AufvimkYbjZ6SWXNG23AK3Ta1+jOPiXfpxZGPB
jYfOwQHs5DLtTGctk2uv4D/xxbwDpkPpfQC/SbaqCaDlmQLiikNfGNy8mOU2
hl0uSq2s95QlcOfl5ke7bU/h61+5XrXf2VpF1nlL2T9gBTySZQj7r464MkH8
oaxbCBeaGvGvs9tWXmtHJgN8LrxzDBHhs0CF+i4yn1AUVbgSVYsPcQHbOEuk
QVU4x2mHpGIJnf1YlCqH39uV0/nNMiZqwuLRH8996fkjcpXTOX0DsIZjszyy
qYd7OdmKLJimB+kwpoc36bSKsJyE8NFHax/wu82hYHsVqYYenHFI8+nxhSkr
njBedqW0RQ/s9n0COhvFjHGh/hguuEsxeUPQYGucwWx6XiZjHwSfG2fZ4zAh
pw2qjQ2558hdT2nz2G1m1P6Xjsyi/qgYLYYCMi9R9d1X7g0J86pHZjqP5eo+
OnMpRowtulYPS1/h+3RikbPplt0EMOD3rpgMzPdRj7iilQNDEI4oCqOI8CDR
cqK+FT+IbyXacPMlVjmqDa0LZCmkEus1vsWmF080fEM5I/wpunMAvQTJ5Nz0
4IIgYCR/pAzCZJltO1G6Iqp8YC4aiwTASqoizCkbgM00BLN80FQctHp7tg//
2sL8OaScPXs9xe8NrKTqvCSrRqel5dwF0UFslnExE8MR7bMv/0QOjNvH60mr
B48LMxDyP4jT7SG7yy7YLaZzk1H/iZdyP/w7JD0VKA17nB35Q6MJCYtpwD5Z
uNK+oGMEplV0KqhUwxV7Ml9gsxNwlsPUqWDqvq6M7roGKcmyVSIQ544WOTPt
mkuBvcB5v6bJ+87VAJzHlF4o72hPQRAq5QD82VwPcuH9T3bmR3pmKqlP6xYI
Ha8Am02g9/rVHA2ha+r+aEMkpCJh1Xnod4sjpN68SI9hNgzD9ZRAibdkxHtD
/qTKFcHW4pLbl8iO3NRGFCsA7i85bkcTgOGOgwRXpRvGz7p4sp4IrJ5hz4FC
oxD8vYU4Eie2F1Bn+nINX6cnhTRNYQCJ0ZQxK+ij4h0QFHEcef/8itTVkXhZ
yWfKIne/tk02lY5abOLyInowveYawGh3DpWiWBSL7FyvMkTF3ymjh5DqZsY1
1B+uvp7Fe/ZR/85JkUizoIuFgiK8hpMICfG5VjVApXAmT0ZXefdwwGHP8rca
SCOlcnZaWWzYXklpWdG2shDh7u2LzPqD6ZYQb5/NODiwp3LLWBfFkYyF4lNm
qDstk2/O2ghPYiQpS+Joaei7pMAjDpmgaNftsUgc0vcGSZTbZ+Hd7/86PIIk
Tj+PjjLirtvbmDpRU23cBIZ4ejVwEnM16xLpJxcrHPI7fPcd/q6SuN/XL1JN
CjxZwp1lGExPeWUxrx0loL880jM+dXGOxekFbLpJqHS1nENOsEB3z9NEGXP5
jiL49+b0zAsxGbJe6JLpVs1xwSZoNvqIijjUPcDkyY5/5Yv7oCF3Egkq+93Y
jmXG/FWcC8BJlDUtiVHAeTh2cgAl7hBdY7N0INuBGLYo9N3Bw+89RsDMQ2e7
d4ngJ8+mcyaAujPP0y0046pn4jpygxnhezgwHTiGfAAHLzJOjIjIWMnnhCaa
vtesS04Rl10O5+oud1WSq8NIk58Hz1umRmECCauCBkE8DIIfd11vyvXjI+HX
vEnY0ogrj4UzOkwMqFZafOkM0v1c4LXa6ACBYPeWr3VFgzSBqC/xhcMDeEbM
zk3oEmPEPb4pb5Q7cJ7z1o5sEAqUbbsIgeJdXgM0vcPhty5AosuG4PLQjrFH
YgXlC9OEcYPtgb75Yxs4aCUVQMT9a1Q0Gf71px3Nt1l8uziHYNQLOWDUZSO1
cjkC5NIHifHXAX8P36a57FGMnY2x1gBZEhxssqq39/1BiaucyV3yxUHF12AP
EoB1fyEvDUhRswKXY4DAGJ/LrCb0liWyRGNo14NZJ2b/zzNR4me5etLWRcGQ
aB+xbYcYCERgfuntBiaK+hCVZPqlACx0BibAKAOOk2OIH0IWN3VUzAF2gibl
KTRE1qY9lEDNwqyw0XppWZcjaFsgDUjmIDnmBkD67f9XegJOVebVCW1xmrkp
d6TYEWxpBmXaDhyjzL4M+dZROeQSOBeMRpz8Nr9CFqoyz8r8VbODWXR98E2E
Rkoiwp6hVtT+V531XmrmCmCpnVvF84iJ83CvXhmg1n5+JW8pJiUpdENZ8QK8
/vXQRPKyz0iMLp/t1D7z8qpfimOwEn3pjoATOeefPmCLKU3ChfweeeQ/Q3ge
mgEpwQy5NDOaYfmlV2FFyI5oqpo19jjcaJdvRhWLtXNKCYK3j5ZWSTEeCSjk
BjAGyoKo34X6irYZEeJxQuPJltqtfqwpDSijTsvyeaTpF7QDnzjMlt8pFiDm
bc9GaleYrpdWnN7E+v+eHvsv8hE6Nf+V7whhXu0575ZGP+DtkO38bwTj1Nfo
hinA1gmElsTpPi86kQAh7NFW7uzbdpb6L3FULvwGbKHOOxu9900FS8kapTZh
PpwoMiq7+Hc12MBPkTbyW1cgYgEtrUK/yjT3BywRNAYrc8v4a5kgvwSSWtMx
b1oGcsz2XXexT5dslbvxwCR8ZHcYNc1//ahKRjtVI0QMK5abxWTG7UDgYKKG
3cHE6S5h61hdJdf+xI+ec2LsqlXPUtouO1UTGUgdymlGtVfWxizLPFVxFoAF
VFJC9ExH04AZ7dA4+A6gqMVw9gt9Yop0MmF846DH0FMiu2Pp3Frat9sXsdGP
nN90xzPcQosGqsVcSzAjSNHuEDO+YpIh0WS9lhryAysQmyHzaj2M9WWD43gL
qHgQZzKyWaUHGZKVUpRezYmy6JatyYy8hwbZ0925dxibJY6ERWNiqjKn1glW
FREtHJ4RyxIVXNKbsf38tWKq2kwkaVtl9DVBG1YlUMTQ0tY2cJrGNwR4o8/6
xujGp7MwrMXoQy8PQUnjGKAJJMrfjkKocaqY+1obMRtv5Hm0l0gNNsrXfurZ
KVILDqiTKYQVqRwqgKGTuqSmNIisGf8ePifcjioHNP/atkLiBIgvi0wuVPFG
EcsteJLIlnz1C9aD38gEeqNQULUSKvHQ0/Q+mWrAvgiq5dad8dhATaOj40Qb
MWjRv9UakGoZzez/YIvfJLFokECcO7gwLpLxGRGLu/dKd720hfnOL1OzBM9K
lzBDWVW74jIzpjHld18s/ObQs1l14atHliP1PSWJDj0G6zr7HAM/jUATV7SN
o0j15PcNO2Xjjmz3sDL+yF+rr01PTJyDFo8fm0KFWDevcdS7wXF0SHg67FdI
XJ10AgOOOAsGwpby+00Ubmm5K9fb2PBza8hlsiTBNzwefJpAu0CMsMJ7Pvt0
W/bkbmoW4CSSSQa37ghY5r/YJzepSXLEPI6D+fuCmuMYjiYTsKYvhtOWHaF5
zDsEGc94XKaUJSGL/wyJ1yrOTo1SyNJjmh8oI+JYi23Nqa5rSzF8FakhAh6H
1Jl2MNNaRwCNTa80f1qPEtz+EBx1RylySLPSSGS5yBIeYAN8xLhDVz4wr3HS
IiSl55WtO6ifgEy2NnTB7uaT1dEe2HaDsXbTN3S8qz97v7gVE37gCJ4H68D2
l7fL+vs16tKqGi0iCRwsf1P44Gh21f52v7qvG/Rcz965VVjG00ZOTfh/P2A7
hfQOBk25xV7wdr3ljxqUIEH3LXZSQHMYD/6/c6UjZabEIMKUSaIEj5yxJmmr
/cZpQ0mzwFbBSeyV6mjsc9+x875VssBVmoi5fkcH8rqEHKd0yKxYrikN5GWi
TpEL0UunJovzI+MlZUQwBOkkdgqk/PSpOzyqOFAyoZ7+CREfNr3asCOd+Si9
dRvOMrEIw7yVozjzAoO2+ND2jserjAPSs+GOF6TePRsWlVnqYUwLaR6MqfWN
eDun9GsX0yGrJSy7OMKfVahzDWfPEtLrs604O8PzVbO9ByQ3RASkADzuUW0M
QcCEkkoKG2mLki8Lo0G2aeAGO9HhZtsQnhaoYKZoVgm3YkOAP/JtnxIdKPJ5
bGFNCN0Kl7fmuOS4Hkc69QAZ0dHjBo8t5rbJebnP42qgmjy+Sv2xSfeIASKj
5kay/sA6CiLPw4fU++kZd3ch9wNvkdQHG276cL8AXiOVdb4buLAVf+zUnylr
EttkicVjC4Wer3ZTQIhOT7JM0yIlvvvhbDvzGJseLm8gKE1CGDJ55OqsJ8VK
qumP5C30Gds4Ihwx6Gd4Oqra3mkgIYCqzToQZGt0AxeuTQjE6SeGi/g9IQR5
YRgEF9Ijn9XS/dpOnJc/FP6zy/jAiQRgljkcL6RrcCJXXUPT75YNIjwfI8h6
nf0Iq63yOL4m2M38Zm96F1Wgk8Ppsxl9uKSNzBJOjI3A2/C+WaTKq8BotHv5
ncsjIapGq3bUzh2cBB3DKSBtsGGgZILUCeTc8TioMf47L9EVj7YowUbDtGh7
sohzyIiFsY4HWgCMo5s+lMEOZst1nN5f2ihb+kPZMn4lDgN8A5idbEor58Ez
PDq4+Vd0jNLwF77Ggotjy0xvdLeYQHCfx2txDC+L71az/BUg3PX2TtOU7dTA
DD5zesXykZI2rRABNyEB+J6GXVXTurGzrQAfBdia93+GYGvWmbofTHTxmLfL
9wOSMOu9qF+eveondQspD2N5psJoU/K5IZX7+CF4rtQq7jqEH1FsPwpdEBNU
CnzvNwtmTwB76dJ3HKlXkaz27+KSxfIZmzkJqn6zcjj5pC7wdSldBwL5RnO4
et+7KFDZ/e8HINXGRSJMCJ2XlA3hTJ/y6+D/krRMtr0lpopjklZCuA6UCBc8
5bwdD9LCouI/i/yY1FmvwqJ/o3X9yRov+Fm0TKiaYLCvPQKJdKMLaEoX8h6C
GzfKtSjo+isSKIHENIOzPuoNmI+yQXo6C3WUohAH2mYdIF/ihhusM+9erEQo
d1jOkLvEUKjvqvN2OX3KgdeI47dGL+fHnM/6yPinpy5VGe25QJSDBZHgd3bx
scXmDAFnwo+DXCIWTrrz311tp7P7WFQT0CIkvwY3MHCcwGsN8usAtxHkPNjI
x23WppR6EeISKOTIT5ig40Cg+icN+Vu8otyyNLJHjikuXSqfbmQn132CxRQB
Nqvm538dsY5EMUmGiKEU4WIbb957jnOl03X6VDHZqT5U33PZD981wj9tB9fe
K/3Nxy2QmpbrDR8+VBMmGm9nDOu3s5YlskjtAh2uNfbBdh/bN6ZeWbi+mVmU
sH9Lz1l1AvDEQ3eSO76jryLC1R7uXCWMraMKdp4WLuJ4Kv55/U4uEEeQMR37
VvKQydP6vhvLbp70POoXggBzevAEgpwyiOCHPmRv7iEx+MJynTMUPbcOQEBs
V0vv3PfRSapfHBIqV2JMMBAp2WYKNWrF8rslMWs/eanwmRbnW1MKHnH1YD8t
jHQWEhuBQvSEi6p6Ey8BthKsQBZgyADNEQkZHb9R19wqis6J1E6Dd04vlFz8
TouT/8ag4O4xCt2mk328x0JvG3OsqOyMnBywRB2yJNftnfjfAePxzahui1tn
02DzY0h12WDsZqghWIdaVobqobNiT9YaAZFGUGaWzDgkgWO4PhSXo+FgfQzA
2aCXi2uzFMOzFKMSyWJWbllYBiBTMsQjcAgObEklCFZg9+45ajKGRl56rtQs
E/SB2AK1fmfst1dls0eKRndcAFvBLcrfTKxZJkC78QBR1MSzzuZwCZbjSNG5
TRdAoAODueOWD3/eSVvm8dFGOSy3XcSJrL2hx7kP/iPH06HPhXVp8EkKNEyy
VnUh2u5igS4H/kkrcxl2eZzkDLva+3yR2tVh4sjOhf86gYxliILX4JPkbV+X
T8sB6/xl27U2/QSSNhHkMgHaubFBEHTosLjVhQ6xUOCQpIa6JsooJ1UXVQdl
QS/3oEr7J+msjU1I5shC9xiD1TFtKnQeV3CTIcg39f5ah3ZyCaVWuSylrtP8
N+nMD2nRSRFPKjIJmGdpFhAh/Ftjcv3gOzVjx59J+LTIwY4Jv+cGsQZhQOXO
Z1qVkEXiOsHAc8NzZgKp2YCX2Xe5ozwnAdXCgOBxPF1QFFQ7GY53KW0JIiuR
p5W/RL1SJoz/lrsfo+ie5GUE4Per61hFfd6/M0fwOIJ6BjK9igE1gi4dh1z6
77izzADPRwj0/oLW/GPySQwZYQTy0VArZlPHmgtNzsZwBneW6ROfgtbrjM0C
z4dUlqGpYOK2lrGxjvNyEHiPFnUWircWRx15GH8mEVjPLnEGM5/AjcNUEGDW
jUkwL64i5y/qcreJWv7w45b9i8t+fD4W2ruJd3s36DQbMWDXXAjshI6uJjER
RCk71We10ig8eU1Iu1ildgE7XMbgI4NfmbJYGLNZ950Ya5o7ku0xlU0bfqcy
m4B0g+jfnTQu7TuYLns/by+G7PfNTIP9n56i2JVuh9Wqftk9hmTet6+f6TMi
4nVHWuy3sLyZAOTI6SG5NFuwj0nvsXr7BsXOOhwIZSLOfeDiGP4GXddUutU+
ySzAxdQo/23QKH+OtznJ6KVrJEJIcgAbPT4hlfgfEk6DS5JLsqbHMlZ27W3M
PI1cTxpqO4j3uIlvoGD/o4qQoN/9llXnadW0hqREswN/uyh6JodrLXdumGtE
6KJkxVlEVjd8SBOg6NghSGYwTGeWl1vxBgTzf2wJ11IpwJeqsJ6mVcmZhTXE
are2Rs3fbB3JSXgV1T4PbkRcBDGZwHcJWTTdjLgzRlWFQ8HSo/Ko9BD6DR0k
nBTo8rO1qsn94wTOMJjzg1KcmAXR9+5WF4vaAzUzWs9mBCmKjp3OODIWgvYn
jdJmMCyb2nA8DRHZfBbRd9Ey5rYL5PIUgrIR+ZnGVS0LKVbjKOtWgOeeymcC
vdobvkjhZPg1Lpa8k2Gy7zRNiBIQKK6NIIahcZ8/sdBQkSqLg052cXl8xyeB
84z8HyafIlGfkghexHM3VXM9chqY7jA7fN++PuxQxmgZAw9hpowppY49QvH2
jTmwb4douwX/7Tni4Som/OrqQssj14xQfIHfbdzQVd3BkzkALOG352u5rxZ1
/jLjxMmMztnS5WyHICjFIbqpu28ScrmPfUTWsZlxE4mWEPOu/1noNV2ReF6h
hJuXAYZM75rm9K1rDXvWmhvWTkinsfxXheRcJmclw53v/oUqvTHO5IAfIqE6
ZoQ0+Nl4my/kghJXr4Z69ut7tN/pxprkxSo2aNhrzSWN0O8zcFzoOCo6YbsR
P57Vb1qEBrobBO3B1Dwkql/Tjbgder45hgir0zb93QKGIXAa8ZOm+qFe53Fb
EoWz+L/1Bwl8vsB1ux206yberUI6yPScymeRmnXoGtgO9Yzy/uiJ/hP0W76D
+puHmva/AW1mxP2ppl38WiWlizdEvs27YDpHebI+JIuITdoVX0dGN4p5Y51N
Ej4ina64fHVnF9sIC5olNVCpJmLEWrxjTEfdQDorD2/PyPfDLU37C3MMWT3L
BM2KEF9LBau++nLkjz4hEAOPCxtQ7eqYEdm9fmyKSnBJau3r8P+3wa3PmyTy
0HzOZSiq+k10t1xPHukVkPJYj3TfTg+GvyUqc8DFNqaNJbesgElbKJdIVnXc
MlwZnOny8JfSJo8fx1Uq+Sm1PpFGCL8Vevv0TuvlcAsCSrQZA7NoRg21CaaA
Vwm3o0lPABJMCTqM8vlISo5Uw2xCVyrjEzqRXxyG+9ETSU95rJ18akf8nswH
p3iyA3H8JEoi5qdAwwZJoWIdKX235J+PK5gJBPhpWddE8njoCYbjXUFCzfOt
ALM0LtoAIfeSKl0CdSwJy+ZFPZdFXB3DunfWUkanF4BJreABgVRsJkyf6EVe
Wdp82mZm9w7ndc2CzufzN7E85jLhFryeqYzFWS/yPg8GzQWpWz4dlvGUD4ML
uwLFJopV1HcQM3d83c3mfOJAVluCbtFwHEjFmIAApWr8hMXOFRub8UbvJ2bL
ksATJZakFp9HAJ1gIkPWKbDdPhPd0iIq250eCquphskHfhBCtkSazsPf0Pg2
GulMafW0joAvbOTN1mfnSG15TBERBmql8spAs3atkwi9jxkBRAuZoOzTcPkG
mXhkOOQ7EjZ04bcoI56ZsBZhe9Q/CBEmUKLHaD1aD+fxPHh5ske7+/R1yAR/
EJnDxlPd/VWQj2u72kQZr//LF489C0T7T4mSBQQuv3QIoKoWVH9iXBhovISS
1GR38jyDSV4aIsx6o+9zcbG23yAqpw5K+DCEskPbV9gqgM57+6RaayixYjIc
MZqu91j6b+T6K7QZtZSFzG9/SGx9bELtRGX/k8KqxRrQyeuvqffnYE3JfP00
Wm4oiErh5hPP+q2ezEDL4oTgSk8K9IASHwUnheqdsWqy7mzP0XNyXQLjbhv7
LWmQB5BxrjrnEl77+Yct3lIBTPTYZCxdAni739g+CY8kjvwaaexXuhmvpg+g
J7t3h+7Rh1Y9DXMYtJv/VyiYXlhPlvPiUS6ImZ1GL2K61NtWVVajA72Jy45b
ZRJQt52nzxetVM9dME0LSooRKnDuIO39tPtSLIVo+dCwi35ZpDPfxVnhCtup
vHZ7/levg0TceX+jA9Y+k+Rf3RYbAUSob/X9ilK5GzkdIYfWcyKbNfPoz/J/
3GSbRxEr2WPhV70x6/xEd7vSSPLSc+ffto2TFQ2Kr3fpA+mOCY6y6OhFqWvB
GgrP9rA5ep08j/vIOJNhC62rkjbczgigEnzh7a5VjBQnA2+rXib+ZTRe3X3d
cI1Fr437txT4rrcYsCmGeJeCyx7nTUBrMw1mAV6Hm3H1OPVvyj6tcbpc0X55
dhhBrvdgy6WBSdw3zUw5LfgBiaSeacHYcEmfEN06xQgboFgtTG7wDZUrqH1G
hIqGNdJGYVEarkK+NKL+3wfIGO1AKshIXwz+eMzf/DbKVwEIUUD0orRNqx2C
gG1TAfFmatiRvfoTIOsxUcGf/erI1vgTQBj7qYPvcCVqZJmtqvmveL7f/mZr
VknDvf33oAwjOSoqhGvmghfxjfZauNlI3BbTslYK0Pq9V4qU/Rm25lczM4GQ
jEY8OYj0VJXZMNw5MqSB7v4SEIQlD2WlznoDluRRBjv+R0YWWoHW85VKZ3KM
kmZYx1I0LNYk7ilCxEnACDNiH7s0hDv+2gGWKi65VI2AnB0epKC5a2H2mnLC
1t54mH4u+u6Apj1ndciQ/8U1mM1PnsmgvTmhD3d/nUTUz0v5904CTLAE0/B9
i1YGTiXoL1gY4ojopvQ0YwWqmbE9kC4Dk/dYLcJjzOglFpLvKAMzMqWV44Sa
Eny0wL70iwu+ZI+wCINh21VvSMHqsjJMiyyjHLzdo2Kl6lpqkA/8lXZbOygI
VJiLOY311TLLe8IkgI/A0wKpBZp7almhB+ZbYjW0uPKSc3+iieYPcNtS8ghe
cJgnsjuXYe3BgtsWPqnhRgMoPZdkIKzQBdOCXZ1N26TBIsF/XLw8K8n7xJUz
zHMtCbdJ48GjEkIlDi5MkfUK/foY+8WvZXeEgHaR6jHXaPdeoMGsQFhrskbd
zsd/6zoSjc3+Q9kMvUL/3apUBGHTTVXWR0XZFXKfHreA/yLXztUlw5MlVIiB
e9h8vwn2Y8uiLoh4syF4J2K8B1ex+muosJeBKBNh5aqwJD9G7XnBcvbWy8Lu
vhDCEy88oHJWUlrQ1kMVVGJOXJ3hh5fBiB0AF/6CyxxzKOjDRc3Ym5V7a7xm
qHkoLm/hmukBwK3Hpki3gObPVdxsvbXBU962vrhrNkOu+ZKnWoyqLE7mWbw/
5N5QutZXHHr98E/VgLYWcrb7T/BtB3Fld+u5u0q1ELgf/c4yAoQ7LGm70H2o
TNKUqkjTzysscfK2sUPg9AeTREiPmCp1a1HzEt3REIxml9H5D5KmVGvTd4uI
Xvj7X2a5/IjBTukWus9zJF3zYX7XwrcOGLfBjqlZkQlvmpgEbl1hquHZB97X
5Dc0LbwPo24qwMA9pI50qMTudP7cWbAznWZaRaqKuLu3EvrgyWNsUFLGC+bK
wm9aOXGl7H27iMKua+hswtrp0t3rLxqKYnbuouHC7qBj4R/nBfhOTHPdAdaz
BWnkOTpkZ93N8CtdQi84s75SZHkFkCK1A9fdG9O1A4j2+n26Xr85JRrs6pka
aVX+b54vH7CE9z4r+2NGIWmsXo3rPUwscC4i0oNxtaEMNijpMYZ8Evr6C5AN
Q1RUPKYYu0iW05ggCy+kIFR0fayr0AQMW5ro912Y7QFcNByYk+l2Uwh2qVN6
FzKDrkbN2al3qtc7f/WKOzKOmI19dcJbYl/cp/z222BYQDK6xFLTf2mavuLn
0zxuEF+VEWUJc2sLOgHg/95uSVF2u6xSc2QF7yxcaNxxZwrC//tTf+XuAbGy
b10EmDCXHnm/U0ArtuQ2Jljr8GhWodoC6E6yxhdET06OfvzK15vaat5rQz/u
/PHX4GyTDKFEfSmqjZxzaBDdAScRRJb1O6en4dI0SkQ7KMDV/fGlcxlfiJzs
5rqRZy+XrAHHfjCQTMiOMnd4IJOC+6bIR3AUZvypQH33izo0yHWvIfxJ8Xl1
XBESgcAdHugDr7gkn4BYAwxOUjFnFqVVpycpzT26J+Z+U9qDigvGJiaXDlAx
pZDHVUFq0FwzcUSRUYMbhcyRNuNPS/Q6wAyif1q9Hy4y3pdgYOW00j/guqD4
3LNHMG4f1u1dMC6d9OpamuQ85z2vqyzpAoekoWJhsL2Q3AW7JcUT0YY7L4eV
eFw969afD+MIGCq7TbeuFLxdgIv4bcwUy06Ere0JbPMQ9nxHd8T7L7e6ScLM
CPSvXKHhB2k29NzZ316QVw3zbLgnYbS0I9LbHAW5SQCtuVGEdssoZi6kJJks
I24sZZVq7CklJx6e3fSjPezV4UlbYybGOsB3xAPZDOc1wuioToKcQVTQNPvx
rwE5VwIHhmDCiuOgLmoYk3RTYAiEnrJtu57DeKcW5qfMQHvc1XkQ3N8ZCTmQ
WUxFdtrBWxRCA2LxwYR/ZzfCe1ztAQwFGkBi9/ej6jVWI5NAHhIk3nGTi4Rh
ZOnEh1PZjwg53LusUGXeSb5dQPc5OWsQP1ae7ZZ7uu47kgaVCvXweC/Dm6gR
CLcFQSacjUxPO+xYPJceN4X8URWHyfNWeYXJU7xAgn3JOycntOgcO0+pt2Xx
Q99f47BlgYhXztcQvBJ4X9YZgFL94wUCLpe4tGjufcltStrDmEb1A9EEFg+J
cbXF+jpubdj97tLdrY/ADI4iTnQOXDlzFKt40ZWpSdZ8TycL0jwtWs/hE9hy
nYIYsDKGGsv/WkxyyE/LtyiLe8+7EW8Z7qBVdRAYFEsNjoY+26lZ3SW/A81R
jB0cltQ8isaLFqewxq3CSpmNHc3/xY403GBuAAIBgGfjzRgKrDkdDhuEi1M3
c80r35IlQma/sx7GU3PtpwtzORhX0XrwBY+AFRzIZ0A10+b5Vkr75dxOig1f
ZP/uZentiur5D262LGOz/KXlYIqWxU9uV/w/paPpTOYU2GjKrIeQWFwE6HCp
ILUhIG6QPhmlFP9TJ5VSULZoRFYDSYPns54KhDofef85dJKYE4CtCUpQ23Cd
qFaAlGVPxZaq2HIqJ/1iU0YoakDTcBK0N1fLSm+uz8UsobV8TrXWdZqHN3Qc
b2m5yW7bvzHMf1gAhqx/fXFutn/8oOkl6dEonatzah/j3r6zHbJ99VDW3iT9
qAnHCMuOmszs5wBGR1VP4BtFu1S+u6cCm1B+LrxayiAe7O/SoD1F/lDJ2J6o
HjwHX+tuHGAnjIcYzI8CIVxNbSJioBWoXJk6t2WDH9x13ZmTLPQQPjwfg7Kb
91a8UHMmj7MwXN8hksyjGFoijrGsGGItYjg1Y48uivyiChmNlROGR9gZbOO3
DKUl3ZQYSyZHGzzy3HQWpZTMosgT7rpBZW/ZVST3m4QLd7Q4MeoD4DJ9pJe5
qSZIIy6lLuEv9c+TkqO6+I1iMFrlqMsLi9c+pLsrMWHEKniysTXs48IrZOCc
507YZjQirgt9WB+Z63KwPw8nd3AwljqaohUm+YhjKPggk8FjtoOpMtS6N8cS
+4ikHFXhFuN0UaNe8p5IVP/r9YkKQ/QdhIuG4jsi/FCOXCKBMpfH8j9qzP8V
LAbyGRRSqk0u1MYEQ64h8Q/g7l5GdWYpB4PohiC+038RcOfDmji4BbSHCHwf
kdTsKT3YiUfbX9S6BfjO2c1SupIpuVLhWR0aCvDakq6jMks3Uj0Fp0hJLV9G
NriAvmZmXbgoNfUuFiPoFFKP2kzLHHh/pRf0o57dsQ+F9LE4tobYe99VA2Tf
H5o5o7LwLtNqd9zjn74BNIi8FGDNjqZ01zxGLABAoUyylVS47r/PhfxkWOUq
9TqXWFYfbn+hkWUQf77xvnl+taCAmYhTW7Z3qFUXgQh/+7vjDHxxqn0UnRTS
7yAZU6nhvIzYscNhFwuDjj+zJwdpGwQ3RlOA5ywABdgHivmH0KwHwCsEvjnb
Y2WLLuEW4qMzXbxkiRREmiFtaxGNVoeK+QLsZzwy26rjf/8o55+j24SnMcpy
eP9cbQGOpLL2z0SPpK72Lf96FdnTByPcsT1XOZDUmuKxcINMfBqpsC+wdmL/
BgebfrlNXInSQ2FaKONzByJzUUnh1s3xDb3DBCZKfBjdMqHDwDnR5+dzSA48
EqpWRJ0P3vbgibR60Rj4j/JGOygMCsRpW6TyYOysVFshjkUgwg9LBzMz03yp
iHQ9q3CaIHNzuxEsy3mIzWQVlgWq6P964DnyzbZoFZfsrRcsIr0BwMyWPXdD
uxwf2GZpbZgyAifr+98UBZxMgmHv5gjp4hIoG6r8N1a1xjtbkIQiY6AEEkW9
uxF7nc6aHiwh+4AYJSKBTciruEcWt32a2dOazjkJifpK0uScYaQZMxAWLJ60
b2ucaeBIfT4W8BnrshnRV1y/KwDOPMjje2yO72TpyG17hgHFzjWcpM8n32JQ
dHOfDYRSmAcR21IfXXXN/Po4Qdxc64CNFoyi/dvhFHGGGobprT6UR5fy7Lh7
IQVvrfBneMNXqDKgIQ2psjuVIjQXv54vbp6GmygTqWTHnOEkRY0mG6c9H25j
YnvV5VSDKIVZXI5ai+n24pgvh6tvmb1WHoDeglup2peisTAAKGa8JsXFvFPF
nZUnJSlzdEMQYMQM/5J2eZVY8KC5rpbZxOaO+KsMVg3Kdg73iMH+bPHjZsdS
Pn3Cm5+BkSD1aDRlg8kEPNcjwPWKrvwzULA7SrqUTRGx0QJIzfDz6tvv4QhU
mwHuQmb2mBk4XNUUlo+t2mI9x5TAhjrsg4Quci772tH0k5n7iyWm662FX13a
AFyjSQ9NFBy8Ia43UIDJddyJdjCPW4m43bJdrw5hSLjYL22HYJ2Y3AM46Npt
eelkl2PGQmqlxUMg9ava+q1j7tLSLBEzVyp0kkx4buFWZqS6+7GcdN53ekKG
lQdG6kAiFfJAKHFCZmVrTLakoxPkdkgMV9AKZ6wgkS9QG79jA37hQp6KlLnt
b5sVQv9KJ8KUzpRvennTpic0JDTfhQTfAwQZzTrb5KIV6AVMdxp5rciIZJ0S
WtDNjLn1GEKDE2nam39n2laiDsiK7ZFTAIS1r2j6INjAro2Riky8+DuCpUs9
T5mVQlZ3Hrc+yt+aRO43vB5y511hfF4WkFcJhoYVz2Ma0f60faG66seXz97I
/t5btwXfzcYkTATabNjgaol3FCowzZezPqd66t1hMaiKCM52pmZ3BJseDKFg
vPCIP9BaqUAEJZHBu9oPRPZIwOb66r5bpW7wACqurm14hzJa+By2XMx+N/Cx
Fx/37r8iLunHpJWNtwu4dDZJCC+QpiYQJEiP1MGo8QxzaTjokxG1Obbx1wXb
J505gkM3h2Obd2lwuLfwQxs/yfGBo8RmiyVm32sBF6hZKURCaNPI4M+ZsPQZ
NmHMQ/RfmUWMLVcn6d2/Gq+qZrXvGDs9y5ZO/CiS6ZXmC+SkAIW5aTnKY4jr
/rkLtOQLqpsv7R4CGujUtr4MW9jUx4/Wh/CyhAUpJapsvsD//Rkg17UPV8Tq
TX5xPYKS2A+/UZh4WMLL3f2tS/rEFxWICsvwkDYKBrFONuOAquoz0u/imMZy
/0usNNXvd5IxA+urU/uqIz/wThO55F0MQDvQ9sw8j4tmKMALFVApkCLOzhcZ
t1FyUIXJ4N8jEYPaYiejxolzBaNA27tXETHXpq0KufapEqQQPGC4L1kAqz/a
pGCHI99qaSHh9UmU9NdP301EnLY7qwDYy6oBoJe9qWyW1SD1GcEZJAHDYauJ
wXx2MxixbPjFnyBoY8N+w2SxmsQGicjBgTSvAC805wMNSR8Uf83AO1JOe6eL
i3vS2tfWfL2mBWANabPbgxwxOrvp/nozzYAVz0rEnMkF/WMsw3kZHq69tlWy
szsyOlNR0xC70zUnqyNmAqcYAVfHovSIfntULXF0WznozSTLu0O0AWa+oWRf
fT/r8sLVIyBZCAe9995XwxGjhsHEX4Wg5HWL2TLZg7kiPbrQQ/SstQXTqRnJ
z1LayM3SuQGBpvgvJp/JJM4F7Dn6bw8NSb7uvYKIt0XioBeRhAUGyPIageZC
+C8ShdeJ4qhscljQPCi111nA2S7EX/nZuZdT6iK+i9nhjJe7q2ySZS0skOe8
GR8vW/L6t60A4moCX9IW+/Gky4zV650/e+CtQkg4lFOa9hhHJo2wWgniahya
GEPxvxSKAUvWQSqgRYYOy6LdZ251Hegdpegxhd9LHYxqigq74xxedAM/elCf
G6Y3l79HsXxeTYrXUjmEKmxmYj9PuQqzDzKrrEhrjF2rfQp/SPCn77nhjTUR
d/bCLqznyWbsmeFsekzbqxb4826HdLRtR4nA6M4iM/NP/mWvkM4dU6X4jtMm
hDNwJ/jiXDdw9gBZxVXVr0m90R9d8iacF+2sNStpkUuDxM9nFx3l+c3OlCrW
tH+beunBlbOr2jSR29vt+qx7tjHuIhPT4OhtCcp2vsxDXnHoUD2YX+4aR2hF
CgNIBdm8pB2+TzEVlNi2WReaLJQonh1OcCvcOEi46zMsWi+82UjAdSUElM/P
OY55aV+zvqIrWBfn7MiV9QbaEs5niQAGvJHvqNClJBi+PlmKtVvJKvIrQfO2
i2roPZRIiXkXu7c315eIgtcWf2XzgAzvZys9e/IvRNIRAopTiS2LsRB0gWbM
6ra6LZJ5pUDJADuxg7LHYggypsc+/j6OcmoqLu8QiCljh5eG2Z+H++mgwrmL
0m4TvXjJUSlBwi6EVfalNJvfZQKNDXGlnORVqQ/YHg1R+EU2EFv4gI4cIbpQ
1vvn+pkBdNWgXBs3TV/NifNR8hvG/qUaN8DqI68hbJiLEZHhd5nzy7MyCZpW
qHiKwSYoSw7gejIiMFaHDwZXYAqh0cgWYRdcs0CGJWWp4ZjdxL0k1PlZdUJt
gO6WME7y+2ILvFCe3cr3PvGOv8filPT2yk1d2GMk5lD/LQqmaeL6xqBjkrR1
6BVI9smmWtfam7axrDqNqyKJEL4geU5+oIFZ5lTSyn/gatQVXK0nr7t16ifD
wsukMPzVIsM2c34OmRnFfZHafhHBV6IpDRXRUiH3CtgV3SptVNtP5bOdPnr8
ZcCa/GXwq7hf3tjXNh9HPmdCItsdmUoD0dyyiuxATFkuUjnWAfArwS1BKIk6
bLZ6ggcEbZXQX3jjUsixQFqgeuJygpZXU870rdBCyVD5z/QnOkp2poUjrlX/
enq6rFtp8VQe9YnJaikyDlezHjuzI4ohJwE69y52Qv+tWPCIvyd8iiQaZr9d
YVqfW6geoTXQVfJGcyVEWkwVCodrBIBYKFwmF4GXdiXMt0if0L+ofE3ckFe/
45AMQ0CMN6bF76J33CaPvV8Em5yeOD1lr7iAy8b89F2p0E9SfyalUCKV3BvZ
SI+u+t161mOicChlvXXvKlAASTKxG32uoqJWERnDpC2mOUtuCKTKNCdDL7SI
1ttJCvVUtxu5cOAgDlZ+uOaB1zIj9Vekl9m+qP3lYaw05dlf6hGEOO7Vv/38
Axjby4jgUyYhjzaQt+sqGvTfIRJ5R+HVIjoHdh7ZIgL/6JqG9u8RMHgRJ501
HJOTbJVc+nCKf0H1nCL65IVvlOz5/jnawDAE2fHUx6LaZF17c25CArwHE/Kw
9TSgY5p6jmm/HnHQZ69uPVeLYSB3uxgjs7xWI/yCBMnBcT4qAiYHTaNWJm6b
/TxdFUfHj4AcOoGmrGeV69LDfF88tJIulGcEEw0yKUoND/DwcI2zKf/5xYPR
dbCnISz/3U4UmQOshb/xn1T5pkxsC4s2rpvzY1cAtf2lKiGjmBZnsVBUJSBu
v0eANPMQgp1JzxU1UhxvIh5Zv7KgMHlFePu9zwMZCE/gU04s2nqQX2mYLJCw
rsrh8Os8O3sntv/nhOEvRBnTdm7jV638YU0Us78Qmo9mShUvkuL/6uZtorKM
aO8W1HID4CJLG6DyQfdyNsXXy7OdFscVyyMtthwmsWKjXqLvDBBzNKjeJgHb
AOr9yYdYcrrTq6H0i9kM+IAofZ4Qx4+/Da86sVQ+qI+WHbrZvtXfgcegNBjz
KFIn/KUqIt6NnNSAWsXOwGDphEq+zMb1s/6Yg/2lkUoOZdpJD3jtOhtQty/t
9MulgEek65EsPdQi311ysGg3pxbxwxFvJ97mQuyy2adBx8J6ApfP1TvAWkC7
/YQWp4ArQMggCm6p3QioXSaS8kzVEVwiswZ7PyWh47p21DC3UDuYwD6mL+lc
kooX+cN/QVO7qGWv7nL8o9vvirtyhHhyUIyrIteoJFEbxv3vtdHNjihGE+lv
OBcJAbN2kJCo1Geci/jib9pne0YP328zIXGUlHUCnUfjfuf0IQWz/MdGECiU
ZY/e57LO+bEpa5KZ5aRK9U6yPSzpwbLEi5J/7SnskZGmuHRM5l5WIaMGJ1fU
K6ZZs70XyGIGsqFrrFpg0UfSbfW/tILAbNjrDBjybWTPOCjZIvxxGeTlut3c
6shCHxFLbheE43Hr6ZBD41OfgZF4XDKhaoqRv+ff8yWj7BAt7cMeg3Y2o1Ji
cbxUtwTAuA9y1XmwGM0L4zSdWO7Sn1aN7lLlMdObUY+rwspw0f/+0J/tJZil
8IEBSi3pBTzyALA54CK+gW2uBsv1LHlj3vNUtCjpJZA+dWy8l5qIScbUf2xH
wCc3o5f6ZPihURow839Rqtwo5Bd/eCUeN8mLj6d2J0hUglgFgVyIi1iwAEAF
xnk0POw4oQdS2mnI/IqGAPhNOFqwc5Z3FPmPWpNkmUcVn4TQonGxo+6fweno
wQ/LgBaSOQR5LfUk/DjeFwriXxBDFJ52MEPgp+76OihAlQrKpqD9dSpDuBT7
aEMy7LogCwTraxxgS8MHxYL3fBNNTNeKlk/A5r6MQql5oPdYmv74fy/4d1VR
2iZx6qjqoUm/nYr/x56uBkvIbl0cs3g/VJNGn/vIXm1SslkB3Fhb9MxlIKVH
I/79cApke84hofQfTeajPZO806JNt3tDegbNr9S6DNLbt5xvmh4Q3A9kNdBM
P3KopukuKb1DdMqLqpivrreogkX0kwxWWyDCtmLcsMVCuHV3FOZ2HZ29gEWl
L83hJAlckSWA+8IcR0Ukja4VNjADTGEA2w4rKOfCefQzNRdyK5mFhhYw51rX
8jp6V3hrbUuXk7TONnHBEo2fa3/fhiss+ChlOMH4ZnD5V0/ACnZj+Mc0iMlM
U+NciVoWQ/kArxtqqhadwxJNrpTmxn7Ckp7kqgEpEI/JpvOh6UNaiX05qqP+
uMSNZEMy6U+QWWmj0BsqlKcEvoFkaWXhuWxn1l/F9PJ8oMODgaDp6l2wGKKW
pWEd8gGKl1+qrOt2I6Ogx7UlC9FdqZ15AbkxknPtO+KRKWfs5LSx4LvoKhO/
XDMD7EQtLPC9FjDz84h6CwvHvq+grwyrKeMU3yiXrE6Eun2DTXrxUNYM91ct
OS9l/tX4zYmn+pgLS1UAmJG6vmQ+BOG3c/dsGpCf/u0jYYnbLxe1PNcLhtVe
yxD6HH6vIse5kmvppc3/vIgpImkeupEVQY1wtLx4x37Mx0Ecs+9LNS8NaZi2
lp4ykb9+b3+gpS3Wj/Q+ZZJqvCzotCjerQsVuFIqtQp4S7HPb4uLnPGc/j9m
omVuiAVJBT6xHXeEsZfjJBiFW+i9sqQTThiSEwGVrR3/hrB2VPXJZtRMb4nT
oJUNzSW8agd7kXbZpLLlRD3kVjw6y904OxPz7y1oQl0uDF4Xjxm7g1c+npDI
Q7H0jyRJBmOTN0mZgHQHXXHHhKD29Sche4wf69AmmgFDMPBpYbAdVSiEhoe2
rAX3OsjTHVcXsjd0wr1jRMD6Lc/Lk5DdzTuh4f4gqzOR2grsFdlixCDoRAhM
Cgfki9ne7QzUk1QqyGOHhlp1FzPbDppeTivuxhjUbbDxkgPafvMGPAkrBT3A
i4Su2w2NQCsYSifo+/+CSX8Wtlw5mRRQYU6OYj49PzltWEgBx4TKb0Axo4Je
4a9hkVrpOz+PIi2nyoCN5cVnsTrUhILHMo4TPQnvGwBxgRnG5fgZ1gtSYHcj
j7e6OCDdO67IzK/9f/y5/HKLVfQ27RluE4aU18QRGabp7VpnoRN98pdFa3qO
vXFxJ9PjGTpPhM0Twy1NUSyHmMWqDu+ROVN8/eaIidfEBOK1HTsu55DN1nsa
27U0oMeH98DTatan+YkgVKF0UWiUnqAxzliZj2n5WwY9M5LE9LgdSP0jXnsX
ODllS+XDeui//k5kF7EWDpb0UYONPsgxgOGVpScfl6vp4Mk0Z2i5Tni/E4KX
t7ClUV0bCwHq7bhxIXt0vTOonKrQmMRqeoPjQibQWDmzudttg7M9/OhzPeNZ
5uT35La5KD+km5F2lHYJCMa+vtCMrkyJH9EmcDKB4nlDYM8baCi35qTvTaqU
/Za1jd17HR+y+qMskucNL6CdTLHE2Bo8dDmkYaDoqcsaolues2DzlMvWF2DZ
gpmWYx5dpuPFhgLFJVbXq1BKcTVy1PIZZv51HBPgqPwSSgjzRO0xFMHgilLH
4Op7JJsrEsHGypGvtQLv7QfPRCOn9LWk49UZsaic6RcINl9zGnuvmzoO4mgl
CBn9HGCvGCJCI0bZ0NiNtI8X7tLNGmGQFxGpW29mp2YBuiOr9fQCAxYrwQ5c
AuR38ezzjkHDfs8tBD9iKfJXjhHiQS8YvZ9Ny9UaXEK3vCmrlvQg8LAydjTj
8hAZr9Urt6cMDXPtUFXa9sQoXtzzDSbtrwaOkxhW6noimNyzt8FctpoJw3hH
v0IDHsZq8f45H0wITWzflwIlgMcLEc1ZDQpCd+fBEXZhPt57xqz2toOpfDct
1Dqxj1hiXj+GRLiLA/jR5A+V1UOLKIzVdi8mLwxh+9iN/G1cTvLTvnYg88BN
4KnVzWwJYIxy41+ZH4ZTMyO64kNuiQBMt4SmGJOPFQDxuhBwA/FpQJfAbe5n
jXuuQxTQ1dOBiBP1pnqI+p9iQtm1vXgxhfOetuhUDNGcA7aevSPSxiX+IyRE
RyVNgcxljFFAnw0vSBcS4s21bwIVY1CH19ThwtixBIOOvAJslL1cBz8Gg4tT
vTrCOyrnlNLqyjEI/vc5JzAwAdxbVcQmW+44ngKPrnBTci+jq4pUtmHHsl+H
omH+mZAcFfSPZycgVA9eCbazaC7e4KbOrLrgs8WqExA8Pyoh+Nh9L8zZu+PK
ChVWsOpeNRFZDGqYf61+jRocNK0TS+NIvBblKmXiYAgusvDfRD+AQs7XOvfN
WOH4xRvTOjOa6KU/+V+19M7q+pgFNlyVKVTFTDKR78DOzO1ZqIpxVO9dAZwj
wC29pQH9l/9MzVgo57M+fdk/vSEUx5lwrt4MmNcNvkw7b4RetvLr8cF18nKq
MXzrr3e2fuct9NA+y9lEB0nE8ssjzQovLjoAw4DO6Py+mbQx6uaOI2k0iiln
4OTsg7wnDPvg96esS3tnTsnVBxRWfdRoqMvMa6jlLC1fULYVa5XvKOPOmvbm
24jNFTzFiX8fPwMKMR98oSIxgj/2XvaxhV6RA3judf0z2YwD77k+vpDYvq55
uNohK2WKfNFiBURm2x4dXOpVaVU4uS2nTXnSFPzOOPYcEQGztDDMf3hgcduy
UXO2R2NobjzMoEj7GRRJOz4Yz5kGXtkFMUuoXZCXnnOUuM8SoD35hIpj+r95
QUPGpYCBL2mwBo6bqvm4zAqjer6HZD92PeG/63PGNanqfNadymXAdhebww78
xEhR5au7pYUATiKD1W73ffsOjulvhB3YP97jv+L2Gpr0+Y+DUdywOWG7ZVLs
tSEsSP/wQvPuSwSV2xwXcWEr6JRVy3JwkDLopwe1fZsRP+VDyc3fPbRtMwf1
Duz8bCuSIV+XAFQxvRI960k4zUNPm5xwdvVkG/VujhyXvxq0JfQzhEw7pGTs
DZVzlBxqUqd8PCh2uYizXPBmdSxRVraqduuoSQkn8vqwZD6XkYM3wX+OmlFG
cosMX1HtFY3aDG6TkEBMCW9VhqcIpYtOahszNaFJKnGgbdmzNQhqUCbZ5eqq
wCunI1bJCJN5AGtUcZ4xIIdEat4gTG0bmCDe38EiIMKVZkdR7bYbfquoiFhh
f8gSF+WCPp8C95FZlA1eEhQCCYXPoRv6Rw1g7asHFFNvbiUz4dVVeSLH/agC
fj+v9VBwuP4+agrC3TTp9yZqc/L7SOUftxELBusAG2GpDFuDe24plfHdh3pQ
aIOioL5ZxB8PGJZ7QesFD0xHFGS4z30sINeNAjeGKLiPvyr0Y2f31YeUMPP2
kwU4yBg9CirXly5MNvuFugvAEAPTPTuleoGwwiDrUnfZMhiD5rRJDJKwj6Dp
VoJ8aOirv4iO1goVNz8htcFUOtn0ofmg6LjuN72tRW72uGOqqXuWP8wdT4Mx
idEJbzEXGG9+pi14nBEKJ7i0W3cHTbuyGh1PND0UjM3UAOG7nDlC5ScOp05Y
8QHK0sFAjEehSyN4PzqRHBzj31nZch7JBUD9Dt7GQyKoe6vQzsI10ijYlffz
tcBn+P+Z4xHyJQFKM6F4iNZENh1azKnjpivLPMz2zy1mpqHM9gYkzLLEtnYk
G8on1HsskMV3rTmnTCVb8Pq0WQoj/X/vl59vRo+wAJcewvpvYsBD8vdyEzTk
zjSFbclyrnTaUrB2nfURlN/wX5+M0Uz8uxfpkLGeoQMuZuvf0wZMFSjtoHhr
aug/9ky1PgGcfPqcvnObseDFPQwSpq8quMlUVWph7l9l5x8igwqvbCRhv9x2
oI1SCNmOEOsp/iVloeZlXIWuXK1jwWyV7BJWHSGf3zXoMfvkalRy0yyDetJ/
gPCJp6/nuNssLJTDDn6PW5/F/EjUj9fomsmUllYaBnJb3GRsdT82WiNr2ZMW
NXtiD6XXqsVQsGko5lZf5a4EvH7vMpUQ5xV/b6WDRtU1LPZbeb4sFs9gtRli
mv7qwcmNEWJ6z7dMSBPooxdvcopM5qKGMlxY9lZgyCfQoARFiGzApPzpitPO
sWDgU0aOPSwPD7VG5yvFB0lD8z+IM2FKKcvP+1gCyXK3jWPqFCWPf6DUbPrP
QymHYcVON70I6H7PPN/YckAWm2lFohyDvyIW9wzsm78yXH3kvp4bcp2j+con
Bh6fOHqtIQUS4thgu3MxoeI45YTUuvSBWr61iYZzmhUQZUeGwZKPgoEXZ+Ll
5MXriZom+9Rl6908BIybSVw737na0/t9PGQbDGqyalJl3D4MTQS+Q5W7oQjt
iI341rr9lvgw2iRqdNbBBAJtwq4DCIft9FdLtMAwtA4HQEicD1KNwAHToJrb
HEoDrgTw4gceTo68wZYwhdxSH3Cw0lpBV8tMqZOlTJm8MdAkeIHHThjvg1x8
oanMktYbCK/swPqYHq4pUe54XM91+jHE17+HlnRutTho7DO+/6odsW1354E+
2vA8m7rJp3aTiGSjlGtEownARQYlEnipmvcbd7DoX+11Eh1pnWfx+iqUXsaS
8V97jR4N8MPfT6nWRuo/7Id92kSR74rJy1/jVxbQqZli+lhJ0nWkWpMDZvtP
Wdz+UmWLJBysubHfvZA0r0U5b5ZQssDtxZjXsdOI4iZQqYR56fUdTHs9atTD
cWyh0n5e7JNWgNNUUEODiUx328tCu5uTVTv6g/PvvDQbL7ZpMO9BAJU1FSQW
yRncGBquFYJPyglM8vH0K5LGr6gR6pTRrwn7ubgldwOKlOYejWa6EDrR48sf
/g3AcIU8nU/quA3Y0Q+8mU2fyF1n/V9bVibaL4kDCGQZ5gy7WIRQAkG9ZXnn
HL/rYWHRASvVJW8MEGh/lbAHNNs9dgEOBuwEGBQmOvktQvy2qc/H/lkDfjpR
da8cPi10CLkMaf6zuHt8LC8+uev/tf6Kq0GSJ3NmJMJfg3KFucZ2P1NhYYkQ
QtmlSxZqeEEsp+Gnz4WDN0JOmORn0yIAmnl1qXMZ+e33lDcQKDxSvJIGxGrI
4Vp2RLyFbAhyrtGgQIMCEunUQk8aMcSSoWxI+/mSHR+CNjFpBQTQshCHiHli
uk8/A+eVOUzNo0lhnsqdO+7rVxjuVIRh50undsgfXb95xFrnryw1W20fMtrx
cysCLk0aUDsjbtdwAsyOAyx4aEHBH4dkwjdo14tczAvjKmMzfcMp4bjibseH
1kMD7yRpG+zN7oCicX0pZnIyltHHo1EuFgDC+Shp3wZJXFMv+fhKX8p6aRs6
7a6fBHYbcOHt5xXRbYe81cKs6WFrZguX5mD2T/J+BDCgIK62urdx3oNinrAm
7T9yi7CfCkfwLWLd7HK0nzurhplbMzc2aPZ437p7No3S4+Gjx5rTSV4XLAXE
gCTSna0kPxkxl2yK0HwjJ9HV9zcqFWRoi46PGIW2K26ZNJTYNpAOkJ+Gak5P
5UjT4wcolIMhy5kR0AeFoApP7/+mEkkCq8i/s9zD3cSsl+hR77udr7BFHW95
uEmYZLJlF6v+LuFtAlmvUTVitKbd9q8nWxQvGYU9Et5LFp4UTZps77kJklmL
4WLfp/ivz6lErJHUK7jVFmwCF/ibaS8IDkGQR74GYdPNJm7Ur3vV0Dq45kRb
yNQXdkatNnDTgXcBYXSXrNE6eUspFw757MFItEYBO61x0t3ILygitH7Ty082
NNriwzYvtXJ0O3eg5L3gPNY4zXEQl5xhrAcGh6rhtLljKtFwaf6V1Kk3j50t
qkr+n4/Kjal5ZREZKbpZ/gSxKWuM/1agyhqHS36kHQhGkhp/JS/Ia2fIV+DS
4hP/R0CAUlCpeAN452uGOvllrvJ382vNrm46dsK6YhrLlhruN0hr7irXeS2V
RKOkiEJe2/hkB/zZNFok6G7ZfbI3vNrVOZ0Pe7zb8dkCiRRnY+20CEx6HCMd
4zjcwK2KWa2prfheHCJy4YO0Bvg+iyQH12FRvfe/y75NjfwcmnI8igbCM2a3
myqDhy2eoNL5RZNsKousQgukgAu/9SBwI6OicyBEoaIyumhoc/vQoNTn8C+c
xuNUjr9EspG7QPQPfXXa7eLHGyrdH1vKVHNdYFkhGVykxXOftvnlqpSdx5+Y
Q2xgPYmhHJYHXzP6c3XjLeFDbZwk2EpLSif4g7Ow6yJzucOttJKT4/khdwe1
AvIwyFV+x+HLh5vwMgGzgNX25nQZVcyTk3i2EzDXlfUwKw96MwdZUu29ssOS
WzJGzX1CIREC7Poj+sjHM4YSfl63uNa2RQsHtc2rSGHpfgSbbr1mUrlTVwC7
C7dPIyMvWg+8qXyGXDqbBAbIA7QmUt8jZH1Geag0KrT09TlMg7E86Zjln7x/
vgBtM00fceL7f7qbMHBYwb8lxD2LGuNEbyHo1jXJsBKjWJkmZU1cSK/rtyXO
BKdJvVKCL3DUC03VzI/6YR+SMjHROhd80+73vUx/11YraaAQOFa0acaFPrng
OmTr3lCjbSfoLxkOh4ze5lxfAAvDkR2hc1ODlaFOxzlJ7JYs96wj16ZnZac3
61HBRO3VWNy763tbxfJseHlxMokfde47//wZpASfl3ve1njD25W9AI/DjGvd
88UHiLG6l/U0R2jtcCPMvzFrs5gbZAX0XjXlFt56mzyY9jYW7tANvbbIahVJ
o12ogOVOqVycH1LLWAvp8gtUg4wLzUdn2P2HNHj80E10jqEp7E5CFVL0FXvF
N4CAOtmr+gVynmCkI9Y53ijJ4kHx2aYzA8l6kCyGhbsGFCbDn0gvHS+qWnFe
kxU0TsfHt9FRC5ZR7igIFlv8bLMit2FQle75umkPtvx102ZuVdoD+nn1YgiH
poVwbSU24VSebYgh1qkNyKdybXRxgZA6BGz8hh4+3MoubpPlu41+O/Ak+Bwp
fA9zD2J9dQp/KMSzpVNIsRC2e0B0pI7sJYmCdT5oW+rvSiP8EKLMWn55V2ae
9bsvNIHOkm+YUdpvseSAi81ceEzsabq6llop1teehdZ1bWEmLWmqiiPEMF5b
JRbPqu7KMBh/WxkCjyjjEbMhGU3BPpoFDoOaoUpSRHPMAG0zJcVL9OBEaUQ8
HVEWnhWrRkXP+Y25ynMYxOgTHQPFAsh40PfK7OA9eGDVZlALnzWi3Jg0jSMw
DJffCeiI1tHQfvhQv1uAbq2LG2jOCmjWqCPpU7liyKZJC5FjcFpeaUAaBG08
sumWab4PdY4rD6EaR180aMHx/Cvk4GBOCLX6ici1GNbxplc5wNmczxw6KgX3
WOuh5jgdy8dLQooz1p1GGUL2a+7asxQdb3hr0v4vH21ZJyJfAXXMQh8OEcpt
Vsy57h3SPc74IxJSWDT2LVxLT5Ff1l7oLY3niVWirJp9ZLsWk/iHyjKENEXx
heqOnwHyjoe6agRI2weFpG5gBZrDEmyXiNP7BcGXjPaNxaKEJatxPKCrxofO
vJ2nIusUC7rwezwhNk6g8jRUJoPcLVPI4z3OEr23j7I5gLhn4HNZMh0aNbyr
zQQMMytoBcji8l2ALjRlja7BZZPkddlulh+KNW8y+HRPuHsSta/LaudNCUTp
DdlbaFMSIPv2nphDWpTZ2xL5eimf6OKoxqGoRtB4eY1I4dojZa6klTfD3T86
BwvP5YRJ6kmA0sc4Ypac/t2u0qhC/flPIsMJQrNMghhI63PPb5HvIVfqytaE
OZo3I5sDeWZrv3oLtkDN3qjl9/w2AY0Li8UYIbuqWF4eM1sVlqlly6Lq3QYk
Nb3yo8IbSZncTee16dgxdyd55VEpJ++pjtstI8qLwTFLPZsg7YcLjeMNG0Iv
O5J1kImcbIKJguaJPRM1lIL9e1MU3pAhuI7nn5YeoMacKrezxmwTKgGy0fkf
0WmBsoMmH73AzoOWDqi4vJU/3mo0e1biE9UEV5ftPCMnE3NxSZ8Ct+zttpmX
OyIibVUa6MeXOBIeVzFlxIZczB74FJ8GfLzcF7BwPARQCvFswK8PEMyT3Ls3
4NoJQt1X2X08TFH6mSVGrY5VouJ5aUkgatXFhCLlu22HR3cWsEIV6ukcZj8f
DoriC8znTQJo1mWLHf2jMOdagxuCF+nvCHZ87zB+c7HGTwdrp9vQt7xtKHQc
FyRQczHWY4Yny9REeKoe92Tf1WiECjiNdyZN0dxbcCTtYbPBXfV007QkrTE2
VTWUhQnl7hBym8C12wnFjjsGeD9pWLoDpJLbMwCHfy5me+6d/54J0bHESU84
hArPbvB6kAHJt8Z2F65+le//gS8ThCqGeklf588utvBRx4Sr6tPjw5Frql9D
3TyQu6NjY64Pj+zF3Z2HQs4cCePqv1keuQc+/jkgWuCSqFW75UIRGiGG0Dqt
mdHN1bZ52pMRfTJZjNdhI/vFGomUlGFx1z6QH3YRM4ZUXbxJovvlnRL67zk1
INQlSAgMgFz9k4jrDVe5yPx0Ypsrerp+ugwdNvb5xIhqQDWnkrBQ1JQvQzDx
o76e4iQz4eHlcqw74JdUpKwXBHDT6ixcA4kOyxh/ItoNWGXkbig9VNn/A/0m
XD0WRim/2KP12UtNKrN+52egsGtzQD40a3ZfOBJZpAMWY3YglTfticRAhHru
e/IAnlWe+wzi+bUFqFUG7wuS6Zk58EQbC1uYUUq3o866+ZIbWXmkVhQNRFpY
J94fhpzjjpA+O31vK+6+uXROAkmBQP6KKK9pFiSOxW/sny9DiVjFzPCfCqEp
6bacR4VwypkZ2AKEbfdkqf3zhTGO5cECrSpRiw3DN+hOaDxMPzN9a/LBVAKW
1OPYUGDZH/MH4wLN5dO/T5xVWMh5NHbNmYB6sqe0+0JPMpIdHzH5lo4Nk1f9
QyNijockWi6v1aJvwqETxzsIRGcYsBYsUSKzNCNfbark/QXniIdX99/gsMe6
d2KWMas3M1E4CggLlMxKQHbbrxt5PTXM6Y9Jgeq/wxTRFQkKw9FdEOWTq86V
tfa7xhjkI0wKzlInDNHDsVc1rA2LFdv6T262yK0XxigOzN2yJj0///uzhzh1
uOJYAFiAiCCsbQPW7S+/ipxiALq7Lky3eCKX/PrSCu2+ZDxf/k5COzd1hyhq
c92lZ+XoC29sWF4bcb3Ttzu5slC002n/I0lXlh48vLupIXNIum0pnacP+8Cw
J1FmpvDu15ZdZkEuIHaSsBhZj1wlK2zzaf8W19J65e6aBtCQFgLGdRRwJYMt
2f/nZgYtnAzl3lHJk1Rbdhj2BhSZHvOutEXbsAt+NM1NOLfURDXldAOoOGIK
xmaHxALN/uHMACTsn9ArauQ61pwvIaSP4oY77cN19l2OyzsLYunWEUEWZb/I
K0DJ5cpQUCwexHKvMmKD7LCjPENShL/Lmiq771R6W6tVm+1CK+RPIQMlqZgX
bg0V1cLvebz8++OxIoB3grks6QkSh+qg9Fy+uzQFz6oBdV1a6Y/lp0J1A+IJ
CkCJQ4r29TnDZ6wPPwwn0UVXskJHH484rF0PiMX+EbERaezVWp1qIlY2cgQz
RrukrQ4XyxUpIrWcZpGccSt9nbtCvZkgzw2rJdVs7VBX78bqxknoxfg8LYJb
VFnD0i+rvRoyods6HwRW8r6moJuL75knLYNYS4PcRYNDS+eV0KELlxXG74as
zIQY/fVmM7FOAWKiyXaFSNwI38vGT/uDsuRs1alLNxX2kjUzyPB/SqR9AlMM
1YgVdb5fXlFJipV58e49Yg8s5BL0thwsUTPvC8Lo4sAE1ZdndhdgzOmLKI/m
YHLeHh4mzpTcbItzIBL4qqzhbamNGSoppkxDZ9pnTcMeIJGbLt4Bxq19vP85
dAh/0SNls7xH/gkEdQ2F7roPX/5V2QWa2rLoE9ufGchIrEAXOpjC0rsnI6K/
MppL+ledWoSY+EfjB3XwuTMkA/1Eaxf2gBdZsLhFVSG3rASPdqamyl65HkRS
sxcM2CssztCqavQJIIfAZ8yEdlXAQ6RnjjdnJYniu/NN1xCAmGUR21vt3Noc
Q/g4sANI/WKQArYI1C2IT8Dc3opzM3P++uJGMF741kX6QFdJ/27AcctRoTyR
G3kZND8PivoT9aSsMXbMjg1vPq0oNNvjouT0g45uQ5sUw2CAAhcHWLhEkFPc
HGYF7Djuabf8hqgp1aPdQXejlsyJLxAvKLkaM/Z6ISdugXbvo4WqaxCQIwKZ
rRPkoiUxeANcKogjldmBv9R4fTRNCYbL1lYzkMuUbowKXtqhYT+NPrD1R/bF
p6TKNIbLtKyEGSZ6UxPSVbqg32nYEDdwvrfVDsi8sTjly0eEPlLOg386kCWm
j7sLxC+gu7sP98vRdLuDPWvHYaTmFz16/BvBsavsppIWDA3/DcoSULoOw5WV
BMISZmgloEdFkExC0EDBFl0azhxP3aaJyktycC74/oPJu23t6cBRmkK8Xrbh
orzMd+xNi1BKQffn4IXRfXOrG37JT0ZWjTfiv5YNQr0/MdhxbAYNOwdRjHEC
yJCo+P4D01/B7aPaqsHdXyNrIekVosJCg452rGroJCZUrYCyOuCJ22NTa3Yc
SKVILvkOP6WGoaoeZJhjT6RMerTDLHW399ui+l9/0GO5Pq1JCLHvJD/qd+BD
cfmSMG6LWAR1HI3jorMncON2pWse8l5pjvXxztqheXgcT662FLPiYVJecxPg
Q705Qm54mw84Zwu1UD0BwPOPtaKS3Dc86bOam2oxwPUBjgIr8M4CQLw03euP
nbzf7hxUAUF6ViBegB3xM9hUYBaYzbzHFRc3xDe5dEVY13kYQTWiKM3N/gps
KAoLZ4XDcAfsvt2M7Sfrqm972HeFk9SYw+XXF0zDvgLlK738XDzgAkZ/6jOF
6cEgLf4jhizp8tqaJgavAzQDCBPkEAoqPxK5cSC4UFV713mB2s1yqF8BXLCh
iChOS0/KIzTWKvREMMFwu38vVneRf9pgkr0EJ3iXp2DU5bs77RMq6J7Ej7Ax
NygKlCCVqS0DheGZDKCKb2eOJAuR6meRwyNlqfhalglKAAyPRkGj7RiHYlmi
Xn6+xQ6h7Arv81CT4RHyOGB4XKr2/NHMgQwF3T2VK+K/fP5CUsHAWAPEJGYF
QGAc9KonjrPVt375I8ytxfZ48gtRruu7JHr3Hd2KOSUCRi5uqdP82UdrrndB
Hr5Phu823/N3bZ0CjNHstQc6FBTdP8wzF89OmHKbIIuYG8QXKN5cyclcqvBc
Y4LsA6Mm35fJXYNkEp60+P1JeZuXfYh1GasbPT549jwTADni63fpG5yolmsF
R6v3QtUJKM/mYfIo2W7/ExbevApLsaFf026IJ9SjSggK35hHF98hUwgkhBBY
wHmXLTyhQnXVuTHGfSI+Nq8QrSAo37uqqs9ranX8U9wKkh4uMQYbHERRk7CM
9A8gon1qi23dBwMl61tE3o1SowMcx3T06SsGvZjbcOSM89PHVuJEOtoMnrn6
VUHPbWbBy4v1quy+hgwx/1e6aoqoRuR6ASyEisgYDDPHredlHCGAInmHUldu
Bm8iHlHtiKSSrGL1T5RIKLneUeKi7KXu+3Dqoxj2xxo5nPYk4//yB2Qur6Dk
pi0ld3w4G6k8Loro+gtAmoTMx+i+DavMNpROap5NwckMRGdBws1jEGfxBmgj
qwx4AbA/GCKHjKKg8gAygs2A8Dgb8MbLRIdhXdKNCzMaMrZ7He5cDu7oMAAJ
UmT80bTZ1iQoA68oDJw/JUHL8mcZ0jZNFdeVR+iudJctmq5j8M4O1t139kCo
5rLvQp3GBq20EES5/cp2SANVoAoDulOX1w0DB4C0Y8wC4X1v1JJKCFy3Ee31
s4PmWnbZB50T8ddtZwaMIQA1+c1fFZa7x9GZVQQYCZvkNFxfV7cWpyR44ZPw
SdCaNAbJkBm5z2WnRpKybl37QZTjk54/DOl8Rcd+cnpep4h/nIr+OJMyBM89
2TQ6yMwnRPCpvC1REtmWNoTT7rA89I7U7Tf275FFGP+ZxATluloeMxYWtpN1
RJAS/guNAGQCfyN8lJgbGmQAiT9/q1u2PbaiYS9HfBiIYXEZKnTbqjn9pe5q
UkSRSlfaEvbAB7xfjGMX5kXi3H6gFMSw4VjfVrw9v+bJCA8Qt6A47C0uJ011
WIwkqJ4yjLSKYLD344Tqfrg4F9eYxH8e6W1GV8yOjhtg1CtbEiNDVkSqqY98
HMrHZVnq13CNYFxMv6FAlGUo0q7tFYi+PjYWdYKvHdxC41O1DRNw0MBMl2cX
igxLCTNdZgLKQCAfMJqOGlSUxRPrpWLgD31jKlnNtRs0r+o0AswxL0747qeJ
hx31tILCqEnvfE143vI5ueol9xtXvG76hmC1IDJmEzgp88uAA+ekTGFqHS87
Ww6UI7cr43Ik2WYGkDliCnwAXdyjxC9MwXew47COSHt1LcvEVwvW+Y7Vq2ox
qBieQPOa0rAED5wpLXsIDZc8vSLEQeFWrPYlBFr82QmhFKkrljKkUVKHfYWK
cy5iJqeNMa74Xe2mdRTKkJlAo+ZFORlLlXWQPlx01ug/s6sRLyIG0fFZ+37U
kQAQh1VDhO9XkE7j0aiBxfiT6PB8QD8Ye1a0XCV8jaCXBDG4uOlv3j4wwTwk
FqmstI5FvumiUMURQfKi8kaMBybM+r8jNOeFvU7EM3s2IYaZvXdYiGOjNLiY
skMUu+MygyHRxhzyZCsZFJz/sGVT1z3Utanpy3viVhPzcv2DcOY4RFl+zzHT
8MrrdViDFsXQDmPRjttBEe5CU+X/OClTC6HOmO2ViMA9bte4+NtypIDPCHRz
imU3+3Bxnk1vpu5WLiqkybPGoaGyYZTZIjS7rom7/P6EwLFDidBdreiPkG5y
T9E7qWLuGjZc36yiwUd/yCjU6dLOtB1zmj65WkwTwALp1VhQQc4mcDI3pMIh
GiPQGnudOWYoNzWQRbQ/l8vLtS3qfOgUC4sxspaSFlhFK2jljw1GalNUCUK8
qXoSWCXgNOPy+BQMj+wMJsRazvJpRC4a/k+jRnPUdMuRD4J3TEti7R1rrotf
4kDr7zu0QJ5IKIOrmyzxv9LqcAzH6Lrs0JivL4UyC2j3mNUlplypz5tpKeUI
BHPi403vUuJqOlDGFTq61mYrV7n9XtOOUw5LhVTqcR4XS88RcgfF9SyDatGL
gHx9J10SUrq9hJzStfB5Nf1rlbn7v/9U14vY7OT1RIbIOXrl3zJiUZ/vS9Nk
UI5tPE3q3s6nsNBonmpnNUjfWoBcTycmcPDwulSUo1G45Zyma3VGvlS/P96e
kvKNm+X8HKG9ahmIxtOfX15t8oskAoNwiuDTV1v6wafa9ENlI3CImDoTt/8U
h7dcDWcZC639hilHZqD7QYowLPA/NS3ucx77Vc/lD9127YyEGheBMzEPOMmB
tgmJc/AHeCXaJfu7Z7DzgTGs8MuHNKxXipCccvN0aSmBySyJ3Eo7mEgc83qZ
IZkmIJR8V7kDo+se8DtXoFKXnteXI4BZI07z0e1rvvHGRFIvW6l4pa+qCIeT
WT5ceSMqx0RR3rT7Ly6YQ4TbsRJHwMh1W6sLpeRMRqrZAZqlfQrw26Sz13ms
sgpvVutNjxJclRkPQmx5emHWgHnHwlB7rdXasKtrIyMFC4cgEnZ0ZbBI2E74
19YVphnpwKGsTlFI8aERmKbmgl3ZsWA38ujfrEQPgOG00cs4G+a3SN6136VY
hJz5FK4GhMB6iAHrTsHEJG2wpfDaSSTz5pltoxmm1HyLFAQm5ZhLNFhtiLqe
0e4LJ8febA8LrqgZZHMlBYIXCKiF/92YlHDWgkoGLymjG8wKPfSp+80jDj8Q
rR7EtF41TS9vLq4UlpOIBx+PmnpDOeKMqKjYxaLZyK6tl222yuK25IZXzeIo
IkDPcAWDUeGZeqzajKlJxkgpIAr0eg7jOjMxvc3vUZuSlgGZHFXWcuTjfZ3w
M56af1w2DcYSyrmDqj/nH7SbBRRVjZH4j2IwMIMbwgHoHXeKV9AIlZjIL+37
m1g/bXrSimxdYWTremZYsPJPJHxCQxitvbiyZZH5APFnAEGTfTmWWeczIgs2
8Ayoxaj/ng0t6VpCsMbgvKEzPwHlrOqDC9K8Dzyf91KkF20VzxVWXzQ9mx5H
d9D45VBoyLDARpsYP73GOvcA8bK5SDwdhGh7Q8xrvg8/NFOnoZ0+xMY4adE5
TEKzbCqxyH5EJ4kNT3BHVedMDImf8QgXrk81GNBj1RmWF8C+memWDR6BxAK1
jKbzysBKtilfCAWDKJEzTSH4wDHp9lz2hUPC18oUYFrRGTULxwgoU30oZEB9
PnvhByxA6knejaW+Xvlur5LYctw8UhdfAhecyPqEDaivfN5+nAKjPuUZeqrP
xXspmpPwpqZ3KWJC0DEnhUjh33xpDWrTnjtRc/MrGJ564MXQwHlwg4tiuz25
4RfaaqDteWrEYt77habXWB+ZIn6Y27wi/XiGr1eM/zJIWrqsz8jHs2wv+7EJ
2/OzZgI7VBh4zVjdYcs4ippiCtO3Q/cJniZlEdIcZH/l1e/VWh7ofA7qoVwY
aut+0lCxFsVV62hsj1p81foiAcJTQt5dt3YNfJCO0GoJfau2is0ukR1IVBUB
kNmZX1uGWCCRA3/I0HWR3gnK/LMtXz8AnwmDfYDg3QCsiOfaaRZaIC7tGc5H
OlvBY+xuGg77MUN/7SlkKavBCTLkraJYe6Hne3/urABkP4M6gcxLvN85FuQ7
HR5hLc9EXQ+I6UhJLhukE53v6nxObLS47YTwl5L/OPwhWr0xXoRZpzZN+OdF
6JgrhABBIyPF29TmV2+CVxYx4AhyBmAFBjpe7TMbjh1SUmvbgQxcXU66TIiD
TCG9WYVz4bUlI7QXm+MFzcPHUnWWG9z5rTwVedyGdFbek3ZYXfyglf9cEJcs
/agkZt5pJ+z9ykMg+ifSziU/af7MWdt5rIX+HtLIzeFITQIeslkd0XYmRmhC
XwP75/61UAmazbsP/ahBmJhDf47yyIVrJJOtLGikT2BLD+L9XWs2mszWDNXW
2ZVLEfEYkY08fcsMBA+59EjqtPDwq4ptEGYfVF0TjyECXJzr/sA2qwbodkNi
OI9fgwMCoE7y39SSNf3f+KVS6NsT4Ynu0apNdFZItPY07dNPC2cjx07Uo5mc
+CMjsYKr/Ptjvh8/1TzcefKMr3xPhVjMTH8tYqrz2Dgs2J4Mp5fQEvFPMbQf
klTpZjtM3GMxJqo+FOW6P5o+Z8QJSKR9GAmHQ2wCgtJOUs1yB43expXyOH1n
cTU2STlbTF5vNsJoHLJiYvwG49Ig9P3/kany/GBkAkmknjNOlg78NTGtvAfl
nU1XdlTvy+nWkrgKnz+qfXMqH18Ct0U5jWxwBlpcbp0FzeFEQZaC67YpElB6
pdf9nMItpid6WecZCaOJYgNKF4M5ER7ltamCLgzNkr4Kc7yqi2ShcG+VQICh
FoCnYeMQeWutS67SHUbpFdlWl+LHzWN+kHjFz8wT5ZuA+Ed7LH6xbBsT9sf+
dL3B7DXbuL2XzKmjgl15M9pKgK3ZWg40ANXkTdrbmBP+9AEC/t4keoddvHlD
X7ijVl3o5+QUl94I6qZBtRT4B5oLjrzdQP4GX6Gld0LcqzHATSLwp9shnPqs
1tSILEFCMFFByhMk+Ceh8xKxU3IdQ4P4SSHa8BiWK0QX84jlGy2xu+sq84GE
lQs3Om3tE+hBQThq4EKE+LiaBvCzmcUSgLKLSXT3i+s1bSE/x4J6m/j4YKHS
VwklF0XdnJnryP8MV2FgU+TuTtpGzMqZ7rxj4xodD7KrCUOcKiPlKzRPXIrr
2cH8bwHEVl0Oj5KxSKiscCc+BvbzlfI8K0Xpx6+/eZ0fq0MCFWXOtyxI7WDX
0PGrq2GoyF8gKIcJBTDP9QYYrMA67V0HeQ7fkmyjJtS0CLZCeGJVCoTqT97l
WMdOeTDr95aSv/IzVnDvBOHwLwrngt4MDxJ6/T5/zFiuUOFcQOZH69fzPprg
el0WJoYVeXiO7mIBvWnS5nu7w4jPUg6U9BLLpdKCHKgWg4pOWJYXOQNycZku
0CNFPXqu8HjSR8tmgsTauJKIx9edu79Ezz2t9Sh4p2iTJz/ZuDat8I0EpJ4n
Lgfw4oChMnvsJicEZOUDtFNmqrt/i11AakPess5EAY6MRPtrZM3MbeHrTQIM
mCXA99ij8wcdVjmaC4Qf05Ounywei2fBakuVoRK50M1JIRiHOuW5dKqXUyOQ
3XfmaIVAdctgpCtwbLpwh16YiPejTEo6skfN4WXW4Qx113gCvQ+Sbg8nf71q
sMk8cxcpQ674lGuIolYuIcE6O0HWzDnJ1kPvMJ88f1w+nFcLjnkEshqk11gA
+QBeYmvuZv6uJ/PfIqcRo9O2IitYXvW8tAsM79s0l03R/W6qXgEVckL99lye
dzVJTAF6eKAstwtV0NdFD15clk+3BUOjgWNJJ8A11cdCY392HCw0FHCcCdPF
k0xRggeqCbM4xbs0MT2BpyUyL4sfi7O/cfIUAfobZUDn8KfN9dcopZrh09bI
bOWoAS3PEG7yLp2sqDZwkeoapcmDcUmZJjIK/3EyI3AdgvK0WVpX0wbs58TO
KBusuDpPRyQEmJ0hMm07wSoirtIQrTT8qe6iqvl4CYtr9e7YBBh6O5vy9Bi5
kE/eGTaC53PKrkWo63eVbifxCKuM+QnC9wVzPQ11SayzvWmMmQCONd7Xh2vB
UBEcQyO+Xk6HC1w+yMWUrHGltB3ywmYQ1nqqgEVacU0Dg7JLqGetwOg/+ZCp
kw0xxkKQxA6HicdcvBGAusR+4oaBAhfij/OzFHqcG41VVOP51B6XlsM/F3nk
CfLWQb8KhB7dCvzdehW/q12LPjLz8e7IjNkly6lKQz+sIE8MKBHeZdRd2m89
GVikYc2tb1L1QXBsHozS+gpWxT4nNKEkQ36TlYTrzpkDTsLR2JEV3Ncdlxmm
yCRz/V2I0zBZLPM30J0VObw2WtKN8/gWmSHj/dSDaorzz0qS5/4q7L4fpqXN
Xa8DcuXITBM7Bpd1RjzlIw99XwSG7gnh2v1vCzsRjxk4cyxYQUfsT8OR2+QN
+/qSXy8TdNPosCq1/yCTfQ+k1Xixkv5NPv11x4zYJiXR6c646pxzzB4/4LG6
sqwNiqETmNwhDLlQ5rFLxzl+TKxX/hFtER0c8kqY+hUwT/naVeJtbXXF41fr
P2fmWtPgLslGh7PCKp/xQj9VLVDZV5QLmAhTJsnDE2dxh4/DLmzuZx4kS1ZU
jiz3fVlK4mxNvKabldp0XSv74az6Rz6ywgndFE3c34ibehBIIWrNQypl2PnE
Gmsvkp/cFiSF3mmyu1W99ASe848CQjhq/Z3cgqTxHACTOxECHBz/wpwHTkbg
T8fcrPC4HVHSOm+D4I47wrn4mHvbUcPDyER7OuvTRfiLtGbmtB8I7JDDZEbE
m1wliErAnRRbRaCCagTQ1WyWxFVeQUz8opkXYat8eywtk2HZAdLXuCEDx9ja
gwO3OgH7puut7QOOccja8GJetD5v7WbLzvQIOPwnbEFq81dcymYoCCn4uHKv
LLs2ZXmmU355Ot6I/AUVud4MkpNEhx7Bo14ZUvx8reu0cbQ6gBXGJWvc2GjQ
OeTWSIEZpYZHx5YuNfLg+cuPnOSIVnWEDefHdQiTcyPNReyRasRcadR+SIkd
Cx3cP/X5yMSfHpSBBWIICVSzrJoecF76pAfQZrnIrUPDdF8lxy/4nTeE+EMP
kIj5rc5mSyqec8JTFYGWYU3JEjJYUnOtCnMvkP9GzcGkbYCymMcYr2eS1PaA
Hm86smAe0qcMizsHIE0f3wCFgmyN8MwB3LvrN4+nW3Hzn+ljlCcK11w5p/5c
eIjqx34m0R1XHlK1sKOwq7+4bvHQXFUavugBv66e4j15dsQuK8nW5zjxqpvR
ih9MQCatCwTaMFdO23zdNTjVZWo/6BKjrbBUMBVqcgRnAVix4x5XIWzpErLx
/Tg8jRFjFYNASmRzrfkw/RDF+6QGWFHE/oiQK/HFFOSkbyann5wcQIKndfkS
NhybmxhOFCnKsdTO6jSvJ7JON88gBSZuO4IYbgDJ2zfqI8/syHX5H0z9jS3j
mWSuMSPzN2i6MXVt3oaPu4dS5SdTpRAQpggoRptWwEOd5E+vg/w3yZ2tVOxO
yhIxAovlH8RUYw0+eKAz6Fhq28fgqZNvwtx/KXHYi4hn4FVm/67zCLCsrT4W
a7g7wax8ID+r7I4hrY+ITNPGFpQOGGmhjUYRCOCI9NHvPNW1a7Abl3m6C0Mv
uHO3Y0UXw+nE7/GtLq6j5pYs8Ddw96zvgtod4W3Drbh12qlmMKFPK8EQO5Sn
Y5hJy7vkA+RKhxzurwY2s4oy1UECaLiNcKOvvEWIanSL9d41QKjFo3qOHsRp
2q3nQnVpRS6fPlcwBxp2TFEnMEfxtSNyYw2F+jEDHyYJsivxlTeJ+9eGIu3o
x6j32JYT5UbyzObSzqQqaqIg5MB1zIFkye13vm/YZs89+TNAvLJsf1RdhZMB
kCRvPqBSQyfCuWygqyPhbwn7JfyiFQkYQk+fmswirDjMEhWoNLp/e7GMdPJT
nWo853enpPdH1fx+pZ4lK1pYvRuBmh4V8qrknE+tH/ZcqKVhG5DKXKj6JiRq
YJxWh+HkXg8qxgyJTCWcQzh2JAmgmW2xv638pH3l72xzftd/Okzs64HQm98D
S46eESblXYSKBffWMtZvHrfR9pMr8Vy6kJYmoJScp6NCteD9te/vdKXY9RRO
mrL78vTx/LfjwcbGH+qio0Aqa/W/VDGvMl4cKcMpKkPYn4jSj1Nl9u0A1rlc
7gl4Xy8csIrW+LX2Ok6XoaszoZXRSqVTBMKCN8Lq/FEGQunnGtiqErvD1zOj
D/++mlvtJqnmdgfZqBKJiIzELj7s3sdbaTvmcmJuBvxVuIcr2KHdAI7F49XT
gG9kthyw7HipCi0D1gp31SAdoSoMRoe5P9w/2Za6mdG7tebC/K7iBC5MEbHR
+vJ638gzysy1FE2uP7pRCClz8zwy6c9cvi0Rff0b5Imh8Lw+CW2TabFTETh/
bEDmj/V1RQOOYB8ChWk25AimSx5+h0lQ6sZr8Ry7zK+fv6nsjH4AOP/XDcd7
2bv5IvqsCZBa/Ymtrq2T+LJwBDdBUKKhY/KwxsGEBQy/uZXwOxd69KVrC0LF
zflodtDUbNGsYKQiWMTPZ0+w+6lOP7Q16Q/qIXFXgFfcLtjPSrVDPDc5NVYW
lu6TfHDkgc13vb4qCaW2ScKQcz0WsJ1Mqs3Q1KjmEUG3TNxhbbOXlpUPdoWT
G/X5yelMAq+uNgUOsyuOfjaWnf1Eq0NGG7ko2gF1XeiH5tpmYmR20jQ0RWWq
P8LdkvtpFM3gTWSUP+acwbrPigMNOcFd5vOnHFf2bsSYVqmAMNlemFrXx/nn
1qY9MziKXTZHnfsc14+RU6xr1qiJ960wJ1nuElyx5AmYq2jhXojHTy+8iewv
LbhbdLbPykCofsPZcQ60G22bZOiZecQSCRAoaKXZfIEG9lnGvrd37oQCkvW6
WTqsVI29Wj2wsXWW+ee2n31EZ3uc4eIm50rAAD6VSj6dnplq5Hixcr6pSD/3
gdlP7XKX8DIe6K0qNl5Y5Ee9yNtmjoMhtpH3pVFsW1qucdKBSblod5QBUtQ7
e4/0g1TRaHzMppnYoGCe3wf5fk/AgV9u2Pmfbeb7pboEHKLifuVIVXzRxyjs
WXopBMqZT/vPrD2aAQhNbFgs4v+3GhAkbAUf5wfcuNN8hUvk/JbWRxx8Hmn7
59iMRdEY0r3ZeOJ79c2pTCX1RFzVfOXiTksfuA+yXCX07LGbAiocYr3qybid
o2tVo/C8rQiohxZuI0Y/VNJCpsEN2AARqT9xHr2Zaxy7wLRLmmp34/5qZ+D2
nDJAMtdIoNjg6oUpXXym6dCYZPgEEDMBmmxKJBx2uoDaoyxs5+eUupV2AXBg
Rm+/UmAUy5gy/DsU25lIo7TCMLiblKQ+9yX4xcWJ6xgCWX61zedpWuNbVsLs
tmNhVGp9t6NPrUaCcS5hRhgCA7lQMBRuFwh6AsvlbGSrunacwJ32ZGyKP2a0
nmy2x5R0YqZ15bybZv1J66Ll1fzuRDARbHFL0okX5LQbYbHE13VjeXPVysOH
N2RsQ98Gse1RtPG1gGXqHWrKXK6oi2vmK7gwINT8v57GrngaDitLUW+uyTmS
qGnRF5urinbioIyZYkJDxeqNVG/fmmoS53pSBnwX1dy2XA07tw0mu4yZxHj4
YPzdL0PWfnKLL7lfll5qy4EgawVayD3QHw3nBQHALSRbY2J29OsUkhy+6HDP
+si6dFfFr3fDaMK4GchzC4FzuvUQmMYEDFQHEKSTnlfq+WbGaaZzW3chbgdN
EvNRg8cn/3dAka51dcktoltgf6qQDyMiNUbPdKLcj4AZGT5/8o03OY/6u9a1
zYxtpf94MrOUP/32EfhbFNzYcaJBgEq190ELcsftfK+Nd6nEOCXk+KgnVDam
FzbiAp1bAPTU6sxNLRIiK763bC6gMhh15U0zBKuhsNwFfmArDGHaTQGh33k1
XtwVRN4zLj2jieTOsuQJVvi/E+kbS1O5Dxv0ErbOC47XyNgX6jAXVB7AuPsn
pDWmupb2VLTGuQvBSeyTg1ZBp3RMbju4eqojAfWmN2ecBVGvI1k4QIqDTMA0
VVOderdHwvcylbM6VGRFleEDGYvymIcGJjnSdS5Wpko4eugSmYj3Fnkk9Xoh
3fw3RSF4h+sr23H6qqFH4l7Mj5nGBvYo5bZozq71Ka9v5c4w3iqjeBrXkhKP
i+1HgHUwzK6dBUHH4djgLM7ekys86V608nPaw1178tK9HwPqzy7JSeByb878
YmgD9bUgUM4YmClsbV0aIIlYdcZoAQv1J8CqwnI3+uJJkhtNNSYDNYdXTB0j
xUA6YkuQMolW8gNajTuTwC0A0aIS+RcJHIBeiH14VTz3zxoEnJ92O3RtNo8I
VG+1SKYkSF18eAUxopS0QDx6qdAuxLjGcPCT2jhPxdHpLUSlFM+Ucv5O71iY
sJZecmbgx/Xo+YK832iFd+SLf48OMEAqc0dK+eMTNus6Sis3hEYYrbthf2wB
UHfMkpyAonvjbXHdZUaImDEfD7hC+id5sJUlLvPWWvBzgZqD7YKHxXNVaFLW
wzcwpfg50h1U+SUdwWKQyetyRHw+mWqQrTOsm00RmH783waFiLQd/p4gisVY
H/Pf5YThVfuzyTn6hqxpjMyOgF3S6UqdQWrvUsGXjTGam2MKUaXxmUIv39LL
ZA1E/kGqRF+xOFCBLeT0nXXYna7w3bPqd1IiE+NAE5c9hjrLaJdjAlZ9psd8
1bAjJJNu6YVFML/Kt86CPjzbvIkf92eF9ysNhiuJhQi73lC6jIqY1mKDLnBS
XpJIKNq4T9Y20CucBfUnCTEeiYcWtc+7nS7VIKaHnytS3ru4Ze2Q3+lli9yS
IJUP9FIc2ichDpLFXb9I6la+Ua6eNjsUXvgctFF1wS5WAeIB1HamYQ7033Mz
j7O3Pe+ob0MA09DpB2QNhaV21pFfqGZnd+ngko5mRix++730YQRVVDxZTwzu
zw6JZcpEQD6NWAGUU9Mx4EEoVjvCuNLTHYrAfD5FzRva/vUry4Z1Q1iqdHN4
0662zfv5tTF06NV6k1wWeYg0DVA6OXqtXb0hVBjYZXdWlf8uI9yeyQo/9Gol
95WXJUWsS0PqPU1nzLSzXjrHxvyzNBQspguTvZEJYaFCzGhuAQ2SLM/Ine8q
Dzo8yPYkoYX+L45/IrTnp+AGqkjYgDU0mM6OQ0mgnNYvtAAIWKFPKcCJdkQR
8iNJw6MeZc0tD5IgSmGLqrYgiORCLD5iYIQkRtMxgi7XyRZ8LBJhDRpII/+q
LeMNei0aJrTouoS6112hyU0G2AlyREp124MmrX9AVLGQAZ2YJFsnHqow8TaE
wXUNHipmHEU4utM3PyqXiZJ9WohMVJL5wCL42ij93z6q7gmz+rkq4zLNj3/A
Y2Q7h49xOdzAyy3F5OlmTS9ggsfD2JrgXu0byHImnrb0wSZX4Un5cR0UtJvO
g3VkgPN1oKcItX8r3BdOTyUF2+1VT50mmL+eaw9e+l1h4TdKcPlL8wshFbfq
H4gRuFwfR3kc8T58fI3rWdTzly1RA9A8UmjLlbGbu0AVlVfxfd3sSUHrGtF7
2DMQeuAxRIyJOxraBbPfO/1YQzz2/ENfgW0vXmipgqi9tfxsSLvVPEKAS+7G
p9Oc6AIVVmBJh7cM8wo0WAyyj+prU7Vm6CUIpp3cmEOOpgOwkwVJJHqJ1kDz
IW0AXzTeC60cQ/H+d+1PU42Y3xVTIb8uIT2R2LWfS1uEzEoMTebez6zlId8x
keDE43KGfPd0p+XZiNuj3nG5TBefiurttbefGpGN8wH0p+9B3vBDd9NN9Der
3o4NQDrZcVDx59ASxSQbnZQgM8qQ29kt7ojnCXwwzouvKHYte8YwSnhvJ/pd
CBrz9xBd9OPaZKr9Y6SpEJ0crJzWVL2sxhP2bn75ai/ELP49YnDNS9Dclcd3
pva+hXNlxZ2L5dkuP7bpm8UGi1271/9X4gGqTF2u46gMmLpB7P2LeVgvWpBw
SSXUJoNwjUkpI4h0EqhhhiO6laEbKBCfo3iNEuv+8ZLNV6zftE2L5vPt8Sim
60Gj0UvccPZL5X/THJJMvJnUx9OtAyuY+qM2db3cLUL9u5NNAR+TzlhduOkS
WnCKydc3iBnjnUTM64oYVb/5taIF0fEICTieY6tNSPYXjS5g9nwomcun+FbO
6b3Oj26p6YUJX2FQME02Fss9umTXYkIG5Kqpp6HHh9xwQJTBSa6iGOP+TSxj
OzvpSYu41IKzW5fQApZltuhKJOxBDboFMh7bM9PMaF9hb0PSjDYuTedFxizV
4o/c0NU1jG2eg+i/m75ySTY3rhkuOHNebqCkOv+1KnQeozpshDKuK3bmb0Jn
bDzGQVVVH2mPF1WvQE3Z3cs76jYoqtjDSs/yWwOrXed8QQdVfVKYRf7Wf2lm
WdPLtqVzVecgstmkGLjNfkqnXqQnfBleUvRuf8xeMg8A2MZOl+SLJZOq8bNR
XGBr+2BpYcsyxN+f0TEqXNhLr3ilPD3QvPuU+DzNsWRmUrT0me5e6SFk6AiQ
k2OVO/85ClHQX5fvjhhfIl/rp0BXnSYykNQT/+zJb5O409kimKOPt0qFfw2i
oXl+o9VqXtbNtv3+xbUjNJZUazVFfJQUeinYgT7mtgewkl3GQPDjVx+/46Ot
PJO99m02V3PBMvA9KbDfxyPPyQ6j69cGZHjKRv62bze1AuJ76cQa8Y1Ersrv
dpqX3wN0Y83dW6fikFPNKG7LQEY9qqtw5uNzJIcAdyFTikia+1Zl7JAT3SrI
SZj6KEQOnCvJmJ5aD+XNrA6k5IdzRnBASfK/8Cf9z7h79WpBMqsA7Okz7BvI
Q7gBWO99UoNAKFlJtvNwKe4xfFmxsoCRlk9GsYDdigW3n1jYVgVOoJvbn2xq
0DvsoPUPS2/sE26Ebf+rWyUkk4In0fAQ2GbyhW7RflEWL7ROG3TgZzyHR3YW
qranXD0uLezSAXDvIuRvLs8cqL3bGsLv1o4f79t2f09aCw3LhgtdK6RfUH3/
QtCnC5d9JUazXZp4cUlKWeETjmHODgh/5sn7FqZvpUBdpepqMk6MF7Qk6PNh
/SRC/6tvN+PMpOz5fYL+0blRXlSfb4Li7yqYBBBJFCjllRBWsa3nS6Halike
wxFvYLia7hHkQq6RnEimBZ3v2FBaNbxPMbDU4bdXAmS4mPXxU8e8HLxnJerm
cw4wVzwQ6V+fKtdUxAVlfwJ6I+G32dXUGxEO9T6O+8104rIHnw2VoU51zLPM
RcYBIjSDsObNYrz0b0R4yOwOhviSgW0EML2SmykuUAgueLINDXSKv0F71UHi
R1dXXZ0HgG9cp85w5mH/ao6ga0287VDYV2/aUGw221n+fTUcZLv28m/fV81A
7IMGr1XCEp1nDb6Zc4VYXHHmlhMyV8Ovpp00sj7u8uBED4ry4+vuuehU4POk
5YlUG9aReg+EeibTcpzYUKiBGUTjX3JQuFVPUgEayiiKal1ugHTXC+vEmcSh
zUyFYBCYpnq/YMl0AHhOA/9szMUN11vcm0HqQvMI6BpjwowCwYZnsKL+HiQ1
DBSocTS1qlwIYNXLbQUOlNvyJzGJ5JIVifnzhJwNhAaeUZiJNNPj1Lxa++P9
A/pw+cgD8lOYtgspmivXyPApRLRlneLR5hlpJHbcV5QylAmb62MMdal9Ed2k
eSRlF2iQZR1MlRgSjOrMm4ZHEj/KI1VM0SNl6WJjJ7H0CBpqLPctHVt/voqY
J2QQv8kJMjpH7IrzAlarSrr7adTGdbt+jsUD1a/DUBWmRq3DCucWCyoiU6bU
0/LqzWp0sdSiWMdNhT45sB1IPTW19hl70+UIvUHXT12hAtTjnqYMoIHUxhh6
BNPXUcJCQgOig3+hiFfNjVKAZJ63uxpZnpqDnG4/hxLW09QKidFaQyF0nSgB
JPxyisU+P7WWpAFKyD3lq2gUKNND+fUk1kdTOkBKM+Yfy9w7WwxL5wQqS5Iv
lxQ1X4JtChqqd8pbddwAfqQhrDVPswvbdSTl+KRs4MaVDqCpMubLx9WyrXkS
l3E2aODQhYPjgeE/Ze2z9s3NvzwEbV0q3ApNo0GQWyuNlAFBwEpJvksaeO7h
Zk6kpLR2/W5nWxcMrE2l9XIY5XKYptn0OoKiNsqolTYR4Rchw2NVa6Jk3HPo
Z+QdlElL4rWkKCXjQi0zrBA1jc5feXCxt3x6WChpMIZnMPUcn8Kc+Z5AhnZE
IV8iFX4wdyKmBBkoFE25M/7NYimw1o/fKwe430hyLJOq3P8bss5OLoZ604eR
dI7IYGl/kxIF/iLin1u+iuczYkg7RDHj69Wgj1tC/Qe9z3yFAmg/KuWPqy8s
szNdOFg6YBK4GZCuHo4ssYu/jmm9zxGNmQTUcdPrpSu/wBZOF9xoSvAGfCYJ
6BqmFUIoE8rJk9wTC/5o9ZMzNSeGn0j5sohra5xYB0nzZAtebaa7zroVgj90
dHqpYGDYrGl5B/l0X9K1fPnRkCsNprnFXEagdJ0UcYpzWK5vzKQRQFIBD1hK
LnnSfOtyOslL0QfMw/Iq9PzE+LVYfGYYsCpXCZHxl9s+ZAsLUvV8JUf1GCBh
vi0g5sTBy1pJzppWshLIlb55WEEaM1vDIckQgCk1B1m5aLFQQemQCk3WPEaO
y5nG76jjdeFt89hCbSwNHybc1Ts+XEWUjvqrrv698+E8kKtyShNK+siCUw0r
YaAvMR7OfFCrj6GlxNTdddXEDKIPVJNmT/HJPG8xfrUa0CLfg7AI8KmfGVlV
amsO0HehQUsJ2aj67JP9wL8XlOrxR9AyAdz+Ry7bjfvLoyeMjoM6lddnfvNi
YpWyzkId/y2FeVjm9jvd0XvStc28QdpJyQHimC32ybzgA/+yuxL4c/heLLqi
kRfX/hVCbM34AJxMTLb7IX7Woh7vj0sk5DFFb7YnaqO2Ul/tMa4AA0XwbAqa
+f8oPcCaqRzB97q6YS5tRJYre6GR387z5adZMBOZLacYqm8ht/oOtKfXFMD/
bDd5tIb6KyOzBdhY4XnaOfjn6epcLlfICH0vQGoiM+EADRsFrH3RJ50cDrqL
fbVHw6JAmYm3na/TCRw62p8AdGbYl/NZZAxDEdE3ucFoo+OcpGQym42Rch/v
Xp2lyBWMzRLdCnejrnG7OFPfqsMwcSY+YU5cJerugTCfC9rUhGTTDP4N6+Nk
dUxcPYIQxdju84mrYNA2bYkrJJTeatNnaPkKJBU0id7lzFg6F04Eg2GOddI5
7v8gS/DL9IHyqHc75cnHuXWmzkBdaHyLI1odi1L5khuLVj7CN5h9O0sCSWLM
LOM6D9h+aVrv1WokkX+QYk64CuInGCRg4T0caoEXqFMU3p9QOJ+W5Z4HQod8
zeaSNhixOp1s7JdfexEdF3H+pBTRulzEAImap+Cy0r1MkD8ZXQUp8eY3/qKP
Gz8kah+08+DbuMUy+uzwVLcaHQjFoq1HLsGZ3FILcSkSd3gr3RnZh35OSCf/
zIsB31tFzQZ0JPfwbSSxrOkwfEyg9TIqYw1tMgtt4SYYIWh1BFOqSJZkmNyY
suVcAtqXAAT0z0yasN6hDnvTPmCzAT39TxdGGtQL6yxoxkDl+kLPYbAz5JJe
lrkePnUHZS9/hD4WrXL0n/V4+H3WRaHNyBs28RgJuuM/ab23jxKfTCCzRQBD
v5ckH282Z9b4aPlAI8x9oUmURRl0eKuTkWMyFwlar+G0LMrcjv7ezsltPvLx
9LVa5/OZBvC6TqoNUGECHo2qxXOaNePwhPZTSyCgpTUzF5aiFtB0+jgr7iTP
Z7j7cu/GEReOU/lVsZaQrBoZuIO0cwefHUWUTw8RjNZ4Q9XUMAmOASWoD2kB
cdlr9qC2M5iRJWkDx7FJH+uEmG7webSdg8ONdGdy4VH7zBE6s08Pl6fDMbJo
KIthaltI0THRUkuMpB9CqO8rUBrXwO47E4GtmKOmp+7IBgNyKWQ6vQr+8qg1
DJdqgvizLJI8iqIgffb9PV0XstYsCKFObw8iaKI7zhn/lT08hmppvB1zdvN2
ZWYRLJAVR1ldUcf97mUlvkqNNEfqjehqRs+lbEY3sW6bWAUXxqC7KvWfCdZo
uiwXPz5nOzXQPgz6+HvniX7l1NGt2c5zP4VQdGCm9aXiTsoew2kT6c18e5a2
fbduS6pIdSl1tY+I4jKDd9tIpI42Tawj7JKjipPUvpH8OTgBqqsigmnk62+q
gg94khEy0kijeN+F4HfnnVl/dWDzp0SuI9XqaE/X00g8DFJfFFtv7hEo81X+
+SttHXkALuDHeo1GNMJ4bp6m0yTBJDVXahkbERUftU6TQ6pdDvKyjHZWKSWe
qE/O3Kix4ONp/Ka2VBEt87HVL9Qeam2kuaA6AYldGQSDOQV+mukMax/jaNm6
/4fk4toopXV9Pj2K6wPUatGI61KIKEDvASDy1JdFUYy0ux/9DlLx2SAHXN2a
vo1SLCJL55PhE0CbZfvQkJCrTLxtcbMVN+vpBNtbzmUDdZ+5oEXj3v2BVGL5
NwU8Z+IokGb8vtXmfz7g6g+SJSerV7bWNVMA6m0HT6W40jYnR6kzwnOCDFZs
j8LZU1FwYaDEdRqwxLI960uF3+juNoUkJBCtJxDkzLp2C+VRqs6fvjRGJgFy
ccCNZB+oj1r/ijzWeig9qF3FfK6r+4XVAEE3lg26JXzT1MVn6ZlYM0NfPr7T
8qMsnHyRWKIQav8+d/DQDKoVsg4XlQd9E+mhWLE3nHZ8L2i46KuSkTLr6OEw
TUd2uinLpNCs3fa368uGOFqmHw6T+UUnjsCxnAtbhyVTSbuR9fC1tzq6XrM8
IlMmI8W+EDm47Yn1WtAU1JlWSax8VPZAGTXKsA+icOAhiUhz1KrfKdOm6JqX
H2ujnqwP4hEzkDhVUsK5P1CWs3iJ6VjopE9uiORfQQpToqrBAqqtUd7BSUNt
/2HEIrnHuNflKbgXH3Rp7E+uHiqtVp5Cha4HXcd3AWwTx0AWMnebQqulQQKg
Q5sODi85EFxka/QxCt50/0TTEkCQDGpMI3FzxMjXWFBLr+MFio6OMaaS8F4k
fZ11+S+eUX/lrxPKbRXmFB+STpSQUFxwzg0HGvwf4Dd/GdZHnmElC87FDbPg
3oVU8v7wsqZ94FIdExuQnKCdf9NOZxKJ5A4o9OLt3dE3RCssB4ql+UAtedrL
r9ef3WdeW84yqyQfCXq4h1FTBcEaSMOVfihG7GzTfuWEXcXgZuMLt0I3gQ8d
/7+3LOp8X0PrRks8UhKdPBeWHHpihCXJA9esM+leR0eR6cZoZPWIlsfHfgNt
96EytyrD2YvSBoo/geKrXdgnjc7EnmCFYzr1E2jD8cK+UjDLaE/sA1vJKuO9
xeU+a2JXXHNehs/tj8wELWomspUgMb/2PW1DQOhtmS+2JQrGZDj0Ybmngurr
6d+5cErRfUz6Cyk2vC4o0mszpHgcJjMH3fAx49Y4QnoNawXQBEkxtLhVII4x
p4nczmfkYmjYY2xHf8hINHJShpJDEtwSijHz4kDbOTwdxaw0MwpfIoJRQeBt
W4Cu+U7JN7zH/EVXjFQnHxXhcjZ5yuOzpjnjxhFJyFLoNDCcPb96C4fT/O46
Dw2bQURCm/mRqEQLcyOWR9MmUWrHmgIZYpulQimFiQDxxuk1F2w46mopQpCZ
B9O/AyXZ3fBL4rUPAtIrocBxi3TipGxinxTzezlOYpZ73SoCcWUqAZ9QjpeM
MGlzR3P4jsu/UcLCc3KEZpx8DMZeYZDX4qRh2wgwhiNJD5e/7FJRZS6d2GNx
RKWnVhgxmly+lvNlA1UQuGzz0HkDuJ5P7++Om4PznrFneZzGvumkzqRwc6Ex
O4ullD7dS3ml/34dmHXAEKVZCr6hkNl5vQRaMgpretO/4htRKAfwbAopSCQ4
QhJ9L9OY2fX2OfLpohZG9xD8QCFKjTzL1ALs+WUtvVgrJ9F1oPzixR3OqC5O
7s4Asqehqa3Uw5m5FmSn4wcs4BfHzAMDtBscUdaRxXkWhr6m/qfz9W2ZLAsU
mTzwFQbEKQ6IuMjO+/fVAAK6N1OrdlQoYvH3zgxugOaqub5GWxI+vhfqOZGY
B98R2/1st7tmKmwurpVyuSZ2riwUTZgbCd5rRWT5Owk73TEUgphF4ru5HlOY
lmoQQPAQpiQcZGxyLwGqbfhk+2QUQ42mJ6ElYH9RfHzKt2NXcOq6md/JIF/f
Jzjf/famgRPrZkXiP6gcTsXDEA50a6L2fGAMiQxVO/32hUaRQtyJUfRSObAQ
q9neLDVO0VIJmp6O+vhkAciXiur+g6Ux4RFI8zVps1Z+3GOszXayzu9+51f5
Qk+meONp4dyU0qhCSiygh45bmcyr2L7MGtoA/68vPzQDrIsCDly/aWfF7h+e
m/sHGcoqwlnNPu06vqghdk518G6cyT1SesX4tL5CVd9LltSzkdU3rcZIEYfF
7uZa1zC6uT2KhT8Q/e0rWXZethUREGpbZTj/hs426Mi3LbRnz7jcxOTfgUlQ
zBbtDmm/qyq+raQU8NNXND2us4tQ5IPbf5n2ZNjX5rPsIxVtQqF5BcWwaMxd
NIs7ZMaekuPF2ruW8VxOqNpAm4FdIBsiwwl3/wUcEirp9rv1oPmmn+ZNVh0P
U0R8g+yf0qoKsemNw1HoEXIWdDswuFPHzvRA6TBI8ePyEZ1aXEMYVJusnR34
6IcLaSFqDrI/Vaf2GYB99oqPt2em9m9kJMoqj0hS26eEGzbrf7gHp14oq/v0
o52dEYwXtGCfCMbipUWbgy46VUma6Mg4YJ3uRcmZr2t8xEfLR1eK/jwETuuw
/fhFmKHYq6WQ2WQz9YGy0mokZU4xM5Tl0cUwShCj7E3QChaZ4xkpOpMPtaUP
kVURGuII085vIJfevlV+jZ0xhJterysTefSeLqMh6xdLE595O2XcKnxoFIgU
2v+ZUx6w+dmmNeaaw/4qnk4O2lZUzwxYWRW/DU+wddP//OB9Pypg73VVO95A
3ZreU2HW+tRpmQfDtxVB8tkJrWhEYbI0jOmUXKMEChxyfnEvwmOaZjx6DKS7
EHzJhlEkYIk/xixpob0RKQcMNt59MaVT7l39PhAXIqu6Tqemhb6iMLy3qZ+8
wWeg4kJ9dCXjlJtRoQfgn4EVA2glO9uWvoGXpWOEtabH4BXvr9LT7jAmL4ka
GZjJHW3DVQMOyBo0vYjzEYCEZeXj8FgGpvbslRnD6gSaQaMNF797LzXfZMgL
pcMftRwL3ytTb8cN4Rg1B2ulUv30q5bufOj1Bp/+JES558ttuP4w2AO5O23x
/a8YIJinHmv3tRTIwvDihiTChDt5XsIq/tIebFsmRwJt+oyJPjop7gUWayPp
6ljRruZJraF5vcXKzkWdiw4LQqgtuO5Wv+kZkflYLXxCOz3mJgb5XAGLDtXY
Zt/B5In6XkdNy6XVF5iDDgy876apGm6YK/w7w1AWCoNCkMDkYInpbScz/B4B
dAmv300jT2TOWfYNxy1HTyMy0N4mjUqZLDDPbsIWe2MIcntFvQ/Hvx+YySDj
dr18bu9S2YOjtNozvnfSpNjLf15h8g9uyB3a+Rsj0cFPP49cjxShqaZlPmYs
ZOzpDvyQgUHsqR4iglXzKu7S35k6gvDtu1Q//ABC37H/7PplXFYuUyzmUBs2
QMPkzNmpinvsRIWhpnRupKQtv7iR5iA7UVI9LxMWfDKVcPMP5LwWTDOPuZVJ
g/35w+1EWjdEmseK2jAQeOXc1p4tpunRsWTOt8JC3x5vmnSu6elBETfdS2R/
QYOJgvCwPszubm2Pb91j3jeXAn0jTWXqObrIjaINWBUIHyHlrqIk8Od8Da59
0bRUDOjelEob6OxZXiEBb0c6V/1fVJDQCK5HfbLUywSJyziumaszMfO7aflx
QwEqmzigfbxEfHQnn14dmJaDSG8Si8EzfFcLm0VRxoRVP1ry+MZN8pBSSljy
J8yEnY/yhw8jHv4Qlp3ijmLQIm3vcc4JlxX7ojalScYR0upG6oiUpcJw5TMG
LoRhHwn/2F6Bd4pxwzEqMTMqRCbllph+n8ZpR4UzzqpgzoI0Cf79/RYIQmfX
2iFN6yg02T5rlqNR2QfZf7AWxrBxS14FE8DFmJPGkc/e4/BGHnFbKc+Q/yqI
hwG2ICgSNUJoVwMsfjjsTL62S2sOEJuFIWESm44FbC0sw/fSfRWLxdmh2Rtm
/+h/ojuktha6I+cOOmCoz0Dr/fkKEZQzeCpDf2RlcRRrc3lvPyCvXV+zTA+Q
DeeLqlnUAWEQToFM/anBiPQrUmwaSVybx2QqcRzo47Br+ypDjoXBNQogJpd8
qY2tnjiCdbf4+RfhqlT9xoi2TBYW5Iucg8SQSlF3TKJA2rNKvRBFw+4kto6t
WAb6/QBvoGpQbxpERfaCYDLLTDCJSVpH6TjzT8g7GPOHCXtyKKA14G0TXZMc
cb2jaGSLHiLer+f+V7RcktupbhVMwzockOEPpPDgA2p07EKMq0xtWVoYioxZ
4TaWXjN7NfR6UcZLKIXY65l93J60Uk4pACMcCskdp2jA6+9miu15SlJDehOj
DqVp53QBHiFIIpKvgDZGFLbGXO9NSGOVnWPCc7lVhQd/jLeAQRUhEw2bbgC+
fo48exErgLCz9eA0pnnTPx25kBbU3puoa0H4BmNdItoH3sopxjcH1V8Aa0G0
jH/QpbooLkQAyPrcmAKXMOdK4JFU044iMtaIugiaEypvUadsytYf5N5KLujw
SlfyvmVPX2yo3CkvfUI+dHUr2pR8oz02ETCmuCWM37lnwfINriTiuvLzmuak
kawouAzRfaawDexXHxuM3H9IUEodyyfOTUERM+/sW0VNEyMjQlcfK76AGy6V
8IK3D4Lt4v5bWpX+Se5kYpUw7bsw7WT7GjXSv5yJhni9ol1CjNEhnZRmTS6+
3ye392sUPcZOnUo5EURzK0p6krsjE4TPF0wBh+3Oe39xYWQJRbImUBH4SWX2
xf6OQbhOuplBQ6Uy5Z6+lxO167LSM/Hkcnr02qTJC5BFRUEcHOwQRHtZz5Ms
x6fmPYcsm2YMwtY8YO4KeNO0OdBRODPkM4ieMKOrTACJFNzKD6CapH1h7Yf1
1JVZhxwegO+SvY73e0BXAmrnlVcKwTSwOIKEKWTnqOtPZNm7Y0lwyd4l3Htn
D5bEY8oOBVCYiDVGuOcAlH5GgEmM08uKJ95UPeyNQ6MgSKSy372LJZ3eMLnQ
eVHBS78dbXYI0za58gIYwY+5txfhg8VoERzITDkW6Gj6fTQfZWjm56yxAa1g
XI7Yrdlh5H6OA+ijNJgRKE9g4ZeQHJPe8wCJcoFh+oZnotDoLn5dj5IEMX/X
JXNLh2nUsSesNhLm9cPYSt3AhbawjHd9v+VBIWGyuUP6csldzSVntgGDowuJ
xs0FMxKyvRduVYv7ehYZFiKrpE1pcBD86GxpiNqyHMYisBGcYA9unaoOBHXj
VKwMuNVfpX5RUGlZ553x1Rbt3sYDCzmenFN8fw76Dqs+McADwFNFwdikW/qc
euMCIGJ4vXcaNpL5oHL96JRGEFx/Plo2zfjbR2kK7teUcq+oP7vMoh98bGBb
7IDtmBLsKjHwMoUEK6IocYXlrkt4LCqe5TVcp1jyyqT88zNd7z9T0eRHEtXh
Ar8qm/rsuyg/5J0rmsh9kaPc3X8BO/v+DsntFr+5+aBVxctOYblRRIA2P8Ct
+ouCL2E5lJngpzTrTRRzLUB9/0fco7BUMsu4F/Wij33YGvY/sCxIyXlqhF9V
vCh9y7JiV7aKPVE/94busI2ZZYU+BeQhD2FUaEbg97wQ39ipMtae+Ai044sw
hOyMV2ERmNKL8srFSytaTuQ0JcGU45EKpjgkxKpVyai2/0jN/VqSp6VKc2QP
1zH0Gqqd1vULFRzrMN73WIv1momPktjy9n5guoMReesst6PA/bDP/EatyBse
16rXiQGIn34UvRQWZyf4n23zacsL6uRY69HPQoG8svIJZnHoBaByoKNb6U6J
+8mM6jd6ECu1cuFTPSDPnM/QJSXX2o4rY3zFVJxtDjE+H5zoqHDYXqByGh3l
u2SSxL/pF8wHSafcbbpdM1CTIPgTb7XF7rnGcFDw4+6NpvwfA9XrcOUiWRk4
TTmmDyYDLFUCO3+k7axfJCedP57fLrUJKU/e21d30j/2gbGdzb0JxVDTaGb1
G/j1CMYL4TKfA4ijT0aDc/uugAk4whJcv1pC7a1XpAFuDqSm8iKMcYbwhcpE
jejivrqXA3rni570VF0c6GrlavyG/w0ZzJenH1ECB0zDB8LkEgW7ROPZZK9z
Zg6TwALg5q9LxNCbEtZ52eajRMH24HzR/G1LHl2Nviq2aAIcxEQmu6HwigJV
vC7fkhQOTuP5h7zqmuUNTRXgJk4PgKRC8+xrNZm7wt2yqZI/NEWG6rdrAoVN
2mBLH4MWH69+BYBlWge94wfXbRTuzYm/SD+tSOhAwd50JPAklHSUwr5LjBsz
pvS3LBERteiq+2P7iigX0q7j7FHph3UaAFIRKFRstLAq6xJfHl0PBKqJDfBv
uoUiozqrvnw5E58S5gDqvLPjR1j27qvP4HXyByo9NjA0azjAY8et//mUmobG
z/odOdhQcl+vXwVzFarR7tyOjhWbOiEk1SqSieDutrCT2URFkN82+ZWvm1w4
WSGQE0bCD7XTT2+wnpQKQjK/vk3J7VOyydpKzse/lA9kIwGfFkTgBf3MjQFW
IjKOTorvK/eFksYCtdbmem5XRRcG2Aij5tLo1K891w3P/Psej1qGEgqvLV+C
yvJnQyCSWwEJHuW2p6ieknCGis1m4HFVaedgoVoK2WZ3hoyD9iuSrLDSd/zO
6j0m/ABkrpm02PWodsScu//4taQB39r07sQJG25gtiBVCwuSHKzUHPHVFRKd
zTNJM7BkPkIhMU9dCREELR4YhSw/W+H3kCDBeCR6EMKKGf2QQOCxLDy1XZNQ
U91+BdRUW3uVevdNkJt4qAE3nzfs3caqZSnHKhpYZ6H+zGRpI7zyngv0vCPb
f1GLuIvofGyhX7LDDShixwL0tKc44R9DRJRD9HqPgnv+IU5aTiNZPhzY6GAC
WgLau86KkJvVrqgO1Gl1X/TLoLY3+I6bINJjkX31Tzg7qtBBHTMXF93YgUSl
ULlw8RguEZFgywxu2LanEuFSsBBLHYWO2f26A8pzgZnw+27l+KM2DqWOs0Iu
9rT1QmrsUfEEWeMKc1jom2wSwf75a0RA3ZPGMyfRPgJeWkn35vrTgOrPFApE
7DsfpJVt3hWYX+e/ZpJjMtjJ083XIx8vb83gK5RzpLKn6vIwqwxswwtbE1oF
jaQP7jyr7GrQYkB2iZAFqsXxRoKk4t+V/A1pBz+u0c3a7sDyy3hRPJQkWMM2
2nPe8hBJcv7YZFfAhYEP42s/w3cK8T4Yz32nL4NVvGUDkRcu8jcJLOuPGY0w
nvnkuXlx1cDbJ7A9a7wv+11q12eExS2WGEBw9UjPdrsg8rLNe190YSpgkyRl
bLuaZuwdG7v52wEl2VnCwASdIwXfMTk2m6qAWrYF/kotvoId85TPtLTkA3XJ
G6UyRTMNlJ2H71fH33C2cLHIoff1fTT+RqVRm7A+TGNupBiHQ06Ko3ATrHGj
lccTMf8KlwC0rfqeysfFh4azbK3vkn22PKsx2CvldbFNK2Zby+GgvO9ZLrnl
+c6T1MWp7q4ve0E3Q/62eLY3NO77+5PTri1TrsIDFQ6Ft1OOqjNj+Y95IS28
gLf2fuzEehkT0lJZhiNWe52nnVT2m9ytFIk2ke+8dPLGfpgk4+tdIpJdaV0Y
7lSQRZCkRj5dES+malYJ68ljlcHrf1o2KBVgSn9fsWXVCkbV7ZCrKMR/jT/q
788BOXq1tP6UyZjys7A4HxzaNa15JM2RTMEoGYZAgHEocsnUY3DgIjQgjTjL
TSE8PVwxGN7OaapuKFBDu1iMVVh/rdW6ut8aWRjHPKU5uxN0TlG9lrh+Mc3h
YiFHphEV7fdS4SNC9Qylbp1fQalbUp1iPFkDKolp1qMfjltRz9x/dOXBp0Ya
Nl+OOrL9fwg5KPrx5XUc9gv3ZM2u7Ky/cylO1/+rTSV+d6+TgFNrdjoA76Is
HdaAnWZ1U0gvnxY+XFrqX3kJuanjpO2c6BtOiBtKh0RggIff3Oe/8rmVI1E2
/tHSlTXSMVGfVchGMKEqgifJlcXqi4im4/uE5laHvNN+NuDlG3pDheFP3tj4
DqocifZ64ZtxM7SMT49FuTPK1H9ys2nS6y1qpjeZsNhz2SQsfwhpePqzxc36
sWsSf5GuE4dx58uqYkljoHxAZU4JJaakYiaNRKf/t/6hDydk1AebK2ovw33R
RBICs7S7N5KAw19GWitgy8O/lvABsqqtK0kHIROmRoUGc8dlvCQwTQyH1cWK
RWCEox9Ivn6bZcs2aTDcFGqlP03hsgIRKqLJX6j8FFbMBDFEEVnT3M80WDQ8
1kSv5OIZxlsYTI3pmdWtIl7LVS/fPBTfuZcqJuF6HOi3ICXkVUG9BTkiLO4O
KSElGSR6H18O+rqxNOJKEAGtBba4nSzepOQ0omQMsH0XwKLyqj6MX6NM2+XS
3/FLnw45XTGey2ZEHsiWwGE1pw7/IZzd4Rl8c9aFI5DSXpb6EYAvgdk7U5XT
WaM2HTkJqTJXFDtVKZVDbNfzM+X1aaRHCaSse6DdHbmOGcj2/gjdwV/Tm57K
iq5NbYXHqrE472K+O/tZQS0aca09zNStX4sJlhWVTf2ySxN5O6FgHJTe28hw
Avk3RQ2kKNxIl7nuP9BIYeNPNC2gknJ6HdGvKzgbjNz8yQdJ7EvnkIdW+0dV
puxfRTL+gsueZMphwjHQYs7E0CgwPGX795oiKPSC6B8KkTiVmS4jk7QWF8Ru
42jQSUONm5IRpQeQm0SrNGc69oT5/pahvDO9FouAHET7DlDcb+o8KQ3J9JmG
iNzAvU+l/jAzWuJwjONufxYbv8qg8gscovbTYNNJ2gIixposyOL4REKIW5eU
IiEQ6xeugsJXSKkdowAYIC9UHHC+O3nyzb9G5dQ/sfulHw3BQ4rkL2uhcWxX
G/84W2E6hSFLDKnlE2UjfajPGAW+OKYKfcuFaNeXQQl0B2M8Z9vCn15/iM9P
dsrxbBP3LR3bW1Cq3uzL1ZqL3d/4xDQ+CLrOvjwMSgNgsuwRhxKpRe7lJm6J
uPXowNUPKKnKpMlnvnUiUYJe1T9pyQHEQ7KmTldZpXa+mjrlyfeMldRnz+dD
hnML0s0PQAaC4ex1FOeyQfXe4SHusn6Wg8Uhl/FEWL3WBYFew+bQ1M9v9l0+
Nn/LnPLlICsomRZU0aAQO1tkGI5i64HEi54cVdb5sQXBh8NPwvQq41ufs2SL
7UIKh/eRd1ImFEooitkH975mmMoQ8DgrxmZWtfNeUUsVo9b0qD1eZQzkdk3S
gDXUhjOfsbPIyefqi3DQnb2HrXvu25gIajQVQbz2kPmwufv7pYrjV6/Titbl
imGuGoS31oRb5PVcywsjl2y7nVVwJTAPTOiyBCjFNyYfuV102dLgErojzjte
MJTgY8dodaimqOHnkvWWK+2hyur3+qu949U3o9i32kXWUPSMCBAkHvdKd0ZF
UTAauWC19tNmxDQwAJrq1a9sIVZfe6XIFTlu0AFMTHhe2FhFPI4lkC+1YOs3
gFbqp+pM5xP0ABF5du//EJGfWjvvVya6PX5IyhQaUNfwUtLhAnP4X4J2uVeN
RQpsO+6bwCNn6KBnpWXWCTtGbqImRaIqUMg31i7SQ7Mbaz7M3Wjg6+5ocaNN
RvhpGG/tH7CCu9hkd0XOqA+LW+uUUz1NLqNN74HlHLt33aeOBKuVWBr2aMMh
PeZEj5BhHgO6ix3OTRu8/8h51TJrqOhUEfvmVK/Ekc61UpP3pE+mGqolEJjB
qWJoq8IKJsXH5WtV0cDrGQ0+OCmawq2N6A9QPzvFMWnVWKoxUrFKCFB6gLeM
+/E7v//JswkTy0rgQ1ISgk/kdlMPADPvme6Q2VJjJiM+9oX6a8D8s7G4qSWz
W7Z48Im3px4zKQZg+7SjYNUyKfpFqRTwMtFNAWV1P7p4YQ5Ee+tu85lCoq0P
Bc3i168iBfqQwB569HwVji8E3HGVITv+QLWC/RkXFXSSDPrP3vjE53gg7P8K
hHE961TRoVEH/BDaHsezw3qyy6ZOdIEucljiOuRsS17DkjgCO4EKZHUhhdVB
nzY9l+Mb7qFSK/1k6rEJ62r1gEGz4w9XgpQXdUyuKgz3XKmqknwq7wrXajdO
fZbTdIa8m+kOWdso1WhiDS0ImuZdM1Q4thi31SeW0khbgIGMbmE/oArSAQvR
0naykruyU6QNtxqAFPmQtikCYk4KCCG5ufTRHCgG7RsZrhih3FGkJHRID1hc
Jd+i00MKxDVc2IpEwmngmAk4fGibV4taBXMjdupSjxbcO4mgIMJlAF+T+mjA
0hvX1t8iLm6GvDrvUbemNgEBd0Tb8UYCCV8sWOWtuv3wSmDYC4qRsLddIN11
wt/K44bjWJvLyHA16mjyhlm4FJQcRjpc91e+E07zmxiwmmtSlblKGRIswf8K
HNvQAAFAiC5KdC3151hV/nVLkSTiox0EAb9S1aq7WEOmq42vgVlearz6BF9E
ATx9FXfdD9vNQl9gsEGpEQhzZWKLKp2eRS+ZVHf8uOVDBM0ZbfRyvuJ+v4TJ
Qsf0MoIHyfLc61Bv0eSNtbQcJGmgw5u+Mp4DAAHvQqo8+sBVe9Khh/Sq7vrj
C80EetxM3YGUGYqblrhXs5JGR4dG5t/nTbBCADktQlvamrfNF1rGPFN9uzkU
ZJLFuodL4zyTWZI4IgJI4CkDhdN6O11kO/Ugf9CKJ9iXl06xM+ucJFvRA5OB
pow++lwOL2TMxGKrT2zIyJsPSPuKPF8tFsFM6KB8BnJyKl5N0PcT8YOUs0yC
TWIXpQC6l9xLluRcbQix53GpsxiwRrsjRmRjEo8NU7LLX7er7LjwMHu5/gSP
rx5qNy6mvELe8EmxnKyH1IK0/gOAvOkrWTVGiYqkYz/8KC5UjcdatYqJ4g+P
ZN2Izf+sD7ORkrT0/3ydD8ir8Aux3+HOlXEAz+lo1X88TQbWwFqRlo1qmPo5
G5lzPtLjf/AYNowiFFVihQwsUdqW21SqDokR+g7PnCQUmqzMP5ZUN3R92kJD
+YzXKFe34/IJdaT38Eocw/WJbUzH6PG5u+rb/Q+Ol2pUDLZFCKRuB84nxBrc
VpWH4+1sqngmFl9CggE67vWh3xopyx8vQXUwXDoIsJpLXLz7SfPnYT9BxJty
Q4GF3OM7gUQrXIr5ByhH/JamShUNfb8QbNOc12xctXpfmMkIQyY2fDWvyK7I
gqVvSwTAurGtVVibLpQRE6vj9vFDlez90lOVovRIeNuA/glPVuOmAqi5ZMo9
/w1egAt+FSIvWr40ipNvy3yXdB7uP55K5akKFf3SAnB3MY3zLviPez1WAS7I
8/Lt8/IjpN0jxrmPFJj0uzpOtGvxkAzZ9L5m/iZwU3fT5tx0aVEg7X0UZPcz
8+5kcWye1bjqma/VzcUMTCjMV2qcIUJM8lkNLWqH+46R11l7Eo8OuJqlcSHn
G6xcolMPRdy/nziEnYKTiJn+pAUx7kz3zJcI1H1j+Z0uh1QjILrVG/KUcp6+
v3EJKfaQ7I8i5r7F5TGEkGFNFUaboCtdmXHun0tGLbl3BC09XsSUMiYSxmqN
OBpGtSQCO1OS84DVlTXHD5hb77+xqOMBI8A1dEuYsz1duYMcCpVN5786LALP
brZVzGcd1VrqxImyCefcFOnADk4JLa4ewEotJx55x5jIqUPl6UMejamXVH34
zA024JsuP6P8a8+oi6GEqbONdS2XszVlz5xb2sAq2MkMXTJ1ZLjZqXSn7XR1
5qEyIe1ycFXMVtj31ZHzF0219/MNIJi4f+q3V3eInvNVcFMurMI62f6vDolQ
q5U3ma8mBkqXV/KHD0L3gvHFtieLZPStWRp1/ENI5OviGV5Pk/wnbe0b/MZA
5jXaZdoa0VNvf58bZ5K4qhR6Gemn/n53LYiigGx5xkzlijO6tj9Lw/84LL91
+K0lZkEUC/m6kthjwxWiDchIAoSagxCecrtiuMacnWF78j7d0aG518gzEwOO
/DiwfJJUl5zl3Hv9PmYUg2q0ZQ1i+Dr6JdFds5D90HtGoUaQD2PJ+9zGjxOo
toOizvWFsLzlVR8w5EdsxiwW2zbI0tGLQjRS3SCOP3Nwro/a+ohkMdclnHs9
dtjnA+h7nxuRPb/xExEus+RZ5nGp45qwESpPSpsmzo+wz9TBpwoeZzpF1zcI
6TqiW8Y0LXgdXZ085N3djKrn2ptNerJDWvaMG3YW5gnbABxOoySNdBccymGn
WfT8aVIXz/RZmxWHpLWNEpvbbJkULjC90zp+L64Qkajssp1g1lGpTm+tlcoh
6HxHCr1xKGHnBF8SdU5LNFbIwSOqVhGlvuUzI1BVuoQe3fJMWSn5CmANA2yN
Rrzu/7AX+gBynyGouPci/MHpV0qGztIohv6iQtTHc1uh+yrxU3z7xCYVPay/
B9QBVa0uX7fePXoG1jDY+ew+1JLcVAUVDMkXzYmmnj/JLwqkPfNZ3eNuakB2
x5FINFOp4g+P3MBCQovS3sIas+7TXg191QIcPkAqBbyhyRC/5gzANfOslU6P
sn8gyKmWv3F62HTbC1dYenzvjtxkURCNdjNNlKYHvMv00k1NUlW9Y6RH69iG
Iks+4O6Vm3g6aAKbrd5VEz7QoSveVf+/38mnBw91uFhFUYBtH+krcNHz6lpp
gDORXu6OQsTbuNs47u0UqA6zEX8fmro8omKhnRDA4Sd4yCW19lGuxeWx283I
+tq+AlZeJ0ZcftkBqngEz5laf8qmPnH1FYjqMPRNBdyuZxc50/vRlwa0UYqe
8VWocm1V18YLMqp5HkDhuF5twbZdSGM/iOqMyOIRGq7e0uPms+fiU3Qs/Alr
9BuwFLZX/8IYNHGeryMA8S6V4tZBkDGMrRXXChaGCbdtwFLIH6JU+bdTqTSf
54yrl42yQIBaksPFDH/3jrEkDg21KYna+MzG1ovGvhZO/J4FjB/oCbqQbJoH
Xp1Up2WnRbWNnrz6z5anYUM/qimaTbkA+25i7VzcEK/Vt+m7VMeye8qvnJT4
OkYYbf6jRvwcszwW0iM6UeVE6BEICfMVfPhwdX/29T5KA2OKBbmQwKlhwTzt
Al+HUPLMm2wth1uvgnMsZZb4khaHebt/ysyVyFxVy+z6bOUHbpcchnY2l1Yg
3rJtl6rB/90+LBv5mHTW7DXoHbeXXjCrPnJ4Al0GM92xOJJ6E5nUJolBdqAF
pknGxffL823kXRcWpbHiy3KjzTc5cc9G1UL/1/lBL4HlF0robj66L0N+gttg
j+9GuyYfQ2PoAaaoItG1RRhUL+HKJE4zQ84Jy+d49q9WE3lBTjyX87fdqx8M
ImS1SMWReMPm2j3FoPZmGlsXROydiFokOJJAj6gTJUn2u2nNtaEjQqqdye9S
OHx70BWAkeTUHauwACpnUiDefTavYQ36aSduWStn4E5Z+FSUWdzRjmzwB21K
LVUwRjzoG2qKPGEfBzMLFBsc13XkJxg93vcHs8bEET8+efKKegFw68QOfRvy
qkGoxl0xgys4GCVTHJXZbOF0p4dxMn/m3BLGGL56GwXrUhGIPqp4ijf5AKrv
OEfsm2yk103KXt74avvPXMMYR/ank92iqDArvlIov6hMsObBvoS9eZ7ZcGNu
OXbyRjtXNZZoksa0fTi+k8U2Q0MKDSr+wKrw1ASnT34cpIIbvZ/bTM8T/HVj
sex2H2Dgzd1EEOHipwAKrMMW4uC3NxqMr5Yq6vDAHVNTwRWJSMfsM9+f/vyb
CXEQuRop8u9YVySHRhAGYUg0r1k2amkngsLJBLdX6zBdnKcUpZ4eeACXXCEn
xXzAKAAF6zgCFwLD5A0ejQeI+NAbDghNSn76PseSGWP+oFawgEDmAciaQSjS
jPdriwhhcF/3pXLYWsjfoiiVavOM2a6hYZQ9MGCxoJ6+bbo4wgeonJfG3nwU
U7iCAMx4yEsbAR2gK5oCDWccp4uzslnNpxd5T/sezDWvTactntWu8uFHGRSl
BXLPhbf2sy6rvCDjL4HbAlDKfS5UJjkka+z1rf5K5DN7vT0o/uqD/QaD/O4f
b8c+iZXCF6pHrqzsKrqL8mbeuepBUCRv34OUwFS3x+ia6QGEPNajjDJqz5/u
rVC546x0hNmSap9ymhpCMh4QMuW1W+A1K8EKYwRYsLuB8uACycK0HcqJ1/xl
lF8GA41fS+dS8WeNKQ5LpzCuzt2VO0fP8KLe/6gZKErJwvlAAa5e7+5+nw5o
h93MhORrOfmbllMxxhNRpmjwHxJ+ka1SZJBfIuFGfeK0ebQdBbVnZ1pM3ai4
m46ITUEiRcSPpQTBDnGiZnbSV4PR4m08G0n5yXhs5Rw5hJELC31JPVj7g1Ak
kD/MAbheBtaAGNR2clt/8rZTivt3DBWQNoUS6osT3rkKRB890CZa336s3YiF
N2dtfcxkw9vLtIeA8JZ41YJQujw1rr7/4YLhpEVsn3MbjXH0slr1QpGbJotM
82bAluZ1zRklC1ATnjl9FLOdP05HvvfnjSy5GtQXL8SdHeN1ArD7L/Ra/40a
F1RKRrGL7EhkdwgutRQNjg79IXZ+UymRtL5zHSNjI31PYvT+9UPNxmQ9aPzF
/riK8noGmNX91eWw2la+a6HDDNuCnD8F9tLvqqrE1BvVOHeHwboudIqE0L72
1bAS8WNwA0IPaM/2jCiVRILOIIzBE+XZa+VQDoy7Oda125b2kZEUNWIM3wOx
B13OZql2LbLBFmuNlZxDSUMKlb1fNOwMgH00BtC8oLdoZkxsjW8DqMSXegeq
dYREd/gUUX3KcRINpY/lGhD4g+xuO1VnxR2Y2SolAjxLf6Nq+mp1d/SrglRI
YsjZYFIBBRVQiwudIXjhR8m02dZb0V2IH/j0KbFQxSwn5l6OGGPNdmK731hB
Cb95B2RtTL1oqOpdn63DTdqvZawT/QSwq8iD9Kt6Ft6htS2AyVC1kd3dhdBy
G5N0Q+rtExrFErcd9H4ljESsGLXSpPVn62PFQmuwQB8vFC1GyYSIiPNi3/l5
2HxO/xrsZUH+QD6rFrOWzjkaRI3DTljfqH7VB14CSyL6SOsVsrAaLTWKDYoK
/+mQDZDu+VYLo4oj9Yng7Mr29ViJYDgYtKaMEghPNqBq/7qAbwwPvDgYtshX
9dQ5AQvVwQMnzCcXBNJsGaUSteSX5QT527pftbwWnhKEpfvAn9H+gwEdSP+G
rdzna2SQo+E67j3crTR6oTWLzjYEA+fwifn8yaeC3LWy9fDJGwPVxJiu85Ri
WYDKQte0SMA3yQ1ajdpNsCWvsEkEtzE9+OQaJ0xLICObKwKjZJxHpYjOLPRc
QJtxpjHPWnaYYZKdhbxWJcjiGTk0gt0A0r9ENJ3wT/3BSMPid7dEVrjVtrGx
2lu7BvbgWRTF25Prl5ECkk01vwebHu44QZMlNqk7sfsZQMwFh2PktVpSwTFj
qgVFh0EKpUXH7qCyzL6OTKMWPOrOR2OyYdT4mB6wyxOAn5rDiKGktUUvy5D1
Bt6vVZ3grOKNYwH6jMvjfp76vLCCUxyJ6Fv0D7ub2MLHEC52sXWyVSp5w04K
YS1hcWKWanOOUII/e7vj/Rk7nXHVlS7oARJY6WaprtpGqJw7ZZHCCd3xDL4x
xpLFaCdZuwTw/Ed+m8HSwtsmj27m5hgAaC8eaXM7kw/aW+XCNIN6PSUiNZ8o
Qd9KfIQH8ZaWw5TD/DcUPyxoFhNnJSV4Oxg89NbNizvkPOu5sYrMTmQ/GdfQ
yNMAM1lE+IvaqcSogoZDob8vLXGj4WIlRwq2mbT1gaJtneZKucOvvWBAlJjP
mQoQh3nk+OAhP8XomK2TsdYvPOv+d3FrvtxAXKXlh2Igj0Hlw+7Wvkx1TXra
CvycvScPE4zDCmn3crqRUrzUAF6LUitFnHiGGafUaZq2rvhD3s/cyygv/ajX
GzHh3XR/8xJ13frFtQeviWZGSyJHYGZn+SgxWSg5jKYtClFw8so/XTP+PlCZ
leC0abedsBcdIIZetFIEhTeVmqif1xDcwOBOJIoPSJLt75JMR2vjz/T0NV4B
oc0lMBLpAt5mlUeJzGkFBjdKTMUd0vTeHmQncIOCbviKnJL+DI/3EPiR0T5C
WeJlSYa4HRyDJ0SyWXSwTSy2CG56t3wuHCIQGR7AyE+EjA9UF2L5NDIn8tuI
BC3WbSNuZfu5mZoqa4Wj6IkfhvzU4KAPsUIGgmsTPrt8ijJ6DcTvgoubw0hN
DSaM0ptPyvmymJm/GyClXTk06YVXpfRlGrCDDXo+f3yKD7qCK2cO6VCmDUJy
wZ7whRy4I/AeMeEz1xbFITL63OOncFCBYMcZVQz22b7on+VbJSn6hLPRK6H1
SpyEmkZLITtqtApSYbqedHL6Kf5toawU628pR40YSFT9BGz3bxNOq3xZRfjX
2JfUZVjIyKTXlAvW+fPTjmJPk11XO+3z16lXIIylPT/bujp+k3OSNBQXu1Ik
chCDgYQ7kq+wOaqSMTaHG1kjh8231Wwt4LN6+M1a/qvET6gnJ1z5WT3TpD/A
D+nMEb8ybTjqmq9CFadJlAqcbRxB5Vt7ZsdhYdW4Bk7Q59gq+HXBPWaIIPiT
9dUHDCmQ3kA/bZccLa14mNsxzOtDfrGXFMW48VEEnyYzZhW1jclQBMRA9A/R
JVYZEx8D9CH6zAKrkSZUuFIv6Cc+YXMv1Cr89bRybyqFJaJbltj8OtzrtlR8
1VWfT8BWjmoeqhbejfPf5qYx3vvSYGlk/vODt3vX+Z/plbkLWduyF1IQG7XT
/3fEm6uUuMzNVEWU3HgkkKYiZDms+THD6BzSSDr0REsUoB0DF7IARqn6ZqaW
lURh6nd/SulVEgbS5VaiEb2cpTGpbxOPZppUJGtkv+i2GnkeTsMtHmjf5pYo
tlgivmoAlp4tt2Uzy8QPlsEFFwcI2K/nrOsTIwD5B1JC29ko+BEPh78FTaPM
dk67qTvDYfWdUvwhpznMVLR4K4/Loid7XH5cKVf9YV52u6eGSsVd5SMJiSXP
AnSJPFAVVgd8/FppTYhURnS++KHbnh8yXRS0nlXM+Ghn7WcqyeOMdS93Veej
lgubBM+1f5PCPoe8mQIit0tU9bp2c72e78ThX20YyhXkBN4lTeC5LrtBlqvU
GKuyLmFb61zqQzetxay3k+0+DJ57wUoQE7r0X4Fi8Nx2MZjs9XOT5+Ze2ATt
qIrZ17WEUmrDy6irg39HpjMWrZFpLFk1jbZvfvrFx1al0ZrPVxix6eVdCzme
PkloH9Vyo8jTVJ59CcRKfdexo4Kpj2OOg1NEAZ8qVkxIJRm5BGfCD/5E03cv
RVI6w64F76lxsXKnjj67lneJO8EpLxcfCgghp53I2cAck/gNAj1fSZ6f3fNi
J+1wJFegaAipo2ec4iOJLdcCcmvNlimYEprZxd74ysmgwwIYpW2xWTU7emjr
uw23nSVMWTYu9sGQBDHCYj1WUMbEGUmv2On+B14SOSr3W4saoxJ0Ycz+Yv5H
pVCplzbTiNUomY4hbGYtr0YpfaRxWMo3k+OSGdaz4r3ruRzN4ChmGK9PQbNI
FodYMN2usvVm+VIi+BQ0Q/D9ZrAd9mLWEVDEuZAoiY6aejFP7zBsfsj7SQvE
vPQ6W5HT21tYJByC829RMiJQG80C97jIK80/qiM8zOOlrZfMWTV1bT7pVnc8
728Pwa4mNZ1eqeC8JjxTshptLIS2KO0VFqwKl5VEA4MtosuzZB9lFojn7cAz
6Vt+3wdQi0wzZfCAF5HgEzexuEEWpV3+EoTnvRIOqsrXFvIMSnoUwkrRbhva
sayGBDgLf8dLNHjH9geCx/zH7QWPXZVDJWf/zm74mub+Wrdf6Qv+1ehxffxv
adV7uta5lqZ7iJEE1jZgtAESrFGqKxwj2IluReOPiN80IekmH4ENozzYj1vf
XVeYsvxutJx8KPCHlI52UEL8XTKqlPUA/xczcTEq6wdebFu9azKwg5DkwZSh
K2TlyVABmWKFYonnDr7mCse19pCwNSKaDtHW1vNjMwPoro50RtMCDGl19Z9h
sq9h247Vgf5guo0WxH+Puvp1moPb/h2NzULnXjuhtjCkhVyfic343gX2XlX9
aywWXd8932vl7SRJAn+gBEYm2VAGg+pU4+Q+WgRmugBGT1Z4hcCkIpzGnR2z
+md+/22ZNFsrzJWENE9kbsIm7Zv16qZ4dqWIWwWkUFFWmCMyZgJwYOpJUfDq
zpM3jTKbMlzcmxPPMBGhHYfk5jwhSIipmfrLXgg4cot/ppS3pRv4ippaoTv7
HzQiLPCKZofmb7iBtQ0YJ/lWvF2DDEbMY+fbZ8TiuhRNtiV9i3iXkKP+aFaf
qIUAsWR6bJgKEG3nn5b12Z3r8U5GIz/lmwEuzAW+VDofdvpj8doDc3aEfIzk
3Knag4GhLvvVbUGaHa8laIQPIRQs4ep41p4+hQxqyKRfx36+2fIMeCgtW5ov
5g4auzTdqcTlBTAleBxnX7/ejANYHzEMzi1FiNwKDtynwd/YoT++qzp1Ao+K
QUAQFl5jQ2GJo68+WfxeeZ1cvsOUYkVApguvWgurLmMNzZIfbxVxaAYi8wcy
3ZRkq0l57H/Yq0pwLRfiQftrlrA8HSKzuly6HtVMDgPi77DKemD2FkT+B/DU
Jj5HqrtVCIAOQR8Jt6uBzanDWISIylHnsuovTKFU9AzcbmRbziH+wnwf6VBt
a4kbo3sFdVyIHjWOSzFv506dEUqOv5pJURDFzz78kbrUnbdslf68oCiCV8HS
HuAG3vswDeojN/5aXiPDdmfwa9+LOisGq5FrILhJ4aA2yjpx56ywZkZoSbKH
QpajnUyO5kCOa90VwqOkqLjZg7byadhxetIKgfNTfyF1Z505c6XLOnZi2Zuh
EDZXfAEjM+zcIMekKsPun3o9zsLoeSh6e8Dt0O5ixCUVSESSd3P9zwAefkM8
70/WNgdYGR6hakk9INY4hh9BTm0a0EZ8CzdbF28kjllDQw0N3gwzsbUB3PJm
0oX3baciPWWpZp+xS3zXfq/yDYuo0Op2WVCdgw/9hc5sjlZ3NvcAN+4lJcnC
kSSttsul0JlLVbVmb5UagtcJTOyOyMhtOzFKif3e01NzNWzL20Iw7dhYI/2j
ezSRS4Z2TCeJ2tUuaMWxMBP6l6x2g4evptsy98aRznPmN5mnYEzNqsMlOmbi
mfLT3beuk07kYCjPCBSUlcdd9VPq9E8i+tYrOC9Uv2uqy28XbpFwHCWwY78a
mcoC1cFqOnoDu/84Jg7gZcZ4/sYkHdFAPHUy+cBCjulNVOortb2C+E87lEgt
3rusQX21QkZHjh0HNOy2L37ZpX6E+Ol4ep5x9QtIOcyD4dChSSzOk73I4NLt
5Dvqc0YxwXqvAlydpJGchUNkfT2f3QrQV88mt9YxltBD25EUJf1A5mZTsXKa
8r+EGGBPut6XGIfQsAcyYdg8/RHbxXlheLlwJTBu9umP4T6SZF24XtEYaK8Z
5TULfgG40y/AEat3fiuj0WDuXz8jsyTFBrc8F1fVEW9zFAlB3Wzler3p3i3D
T8/m6yaaja+0lgmdRsRQ2GcnpWARcEzEEis3FOEmQtbPv1OqzaF/yQ3bGgKY
QHGJOI3+uIJMMV4N/EaAB8dOdw8ESAJ1Qf8x2z9DpDLWytA+TW/PqW84Bz0k
h7ldWjTTiD2WChUlNea9nlXyipD95Ngfl8Bn6qTzR+AVAKhvKJ2BcMMNVGBQ
yW4VsaPE8fdsF64/SG5IFMn/fLLYQCtUPez9tznRc3RhBmdayB+JNll96iAD
UW14S+njhCFpzxze6ge61S4jqjrUV6U6q9tlAAXeYl11VRZu/43kzpWBl/UE
LmybznAF03Yt83tRMwVW9VhDrt5tOlacrBxQhQFOsQTbVcSofjsD+X7CAB1v
K0MlesQRqQx902LRE+jwF+WtM7L+eHmPlPDXJ9EfvV1mN/GlCVCdRmsK8LnI
t5KZFo+p1nn5X7G4WQzwfd5Ns8Tm9Wz3sp5oWSFdKfePc5smy2wdEWsrM/wF
T2CvkbdnhC1NHMOcsJ/RgxTHmJb4B95+qlwLla0RtEahEmOOsDtDzPYRMOFp
mrb3Stg/sz6oebI6w06yxfu02oXlAggYyI6IIA4fj882cq2oioSG9T96Mw18
FTdl95ih+IlUUffP4vDry99YNS1RWCMJDyVQ73wX/cIeAcLjsYshZoQ1POMW
jdCc9bbp47pY1qexjfWL5aLLJo7tepUXdqVFZKsgKMCKSRTqZpwMIx74pUAv
6ynssbmN2UnV4Z296yQGxK1t0JmYMH0KV//2kFpQQ9wIOfHJgeMbcbY2j4F7
GwFHgBYMjm8cXteYxO8k9+nozPDVjeFX5T4hJP8FhC8db2vdSSCueoXfaEZC
2LmVho9LGSp89IiBexUKqR5Y5xq/K5vungRDedsB05w69kcxR+uAPong1nXS
bUnHiBNAdZr1WJFsI7GOeCDAgzTsFFDj/UZebUjmCqeyBmrFe1LhI1XGKGOv
IB34KihXOMzlRAwmHYfw6cVLPjf/Jke9pcy+GOwe+iQnqR7isIRInysJEkLJ
FFzK0a69qa6Pcuu9htuCTDnsrgGn+ynhXnWJrLjbaA1LETjDjWJ/lcSEu0Bs
yAZgvv7jdck+KTbBm+lXRo3Mb9JE8HCFX3QZoIELoc/d8X14tjzkZZr5+QsU
DqXM7liSkGQQNWMtClMw2j9qsVd7ocU59ydtFqJUAbzEL96TGhuQbJuqJ5QW
2UT9VyBaXZyRYf0IqBpVKBcwtjLmmjPcniboAyUNRcMRXG0wEioOC5bz6oZM
QgekPivtC+XtEDk+YBYkpz8x1al7VmPZu3NwKecsSvqRw9uTrNUzdV8fmz9h
QGddeE1cCe8FzWssrhlRX6VNf5YeLT2nGDqRJOr1enMN9xdSHbIcQ3C8RYNt
4/lbLz9APAZV90SMOCNuWUvc4L4edEkcAr30FX+qY105on+zqB/S5SVftOE+
Vzk3C0SoX9NhgInQTgfWzPf376Piabe+8lgMZIkzlYcPhgLnvyQC3ydtWThJ
FQYu4ua3hy+sZ+LPvLTDKvwfXXH5VFp4QK53MDG7Xs4pPeGXK8+zYi8pKU+Z
1VKHogA5cHwG8S1YYUJm7gbxJAWutWeNnAT+IPtc2B/5906OfNCCefQq2hrp
omqolLVWlnTpKW0ML1VSVTBUOvNeE6rr3eLacGX/MkMKDh6VHKCNkqQja0a2
xfpKDPAw6eScPPW3Eh3K2kdQUvhuM2NyGhoLzX5C2taHgie1qsVLxwn7sm7o
SnrDZlEjNogmUwfq9F4iBhpbVEwpjkOJlcRJlXKNMWdth2BwqQNVsF5VVs+f
1dcNTjmO8Z2yrH8LvDDzqn61m2ZYGsyoSKFODLOj/3vUIy5gxFXO5WyF3jAn
vzoSRkG/N0IgCcO1eRdk1NrAmNxnxk27KzhJtUvmzc5vHKuMBzB6JlPGyRoF
Rv0KkGdLox+Su/pzULiTqKTF6vP/8AavPLr/H6A+t6veb/jqM98OktY0y1sK
rsgUJJa2q+mzYC6y9nzE+F5V9n76EDo9s0JGb+zFGUtQ5jgClheM0rXL/1L5
BQxj82QGLBVUB876H6znrs2zc3obdz/8NOkiPzqM4bscUplDK93U5SaYWmgq
UwWMWH6h+O7mblu+u2/808FN7jNss6I6ZnxTkCRU4X6j8vnBdOzsAiJQizj8
N9BNucQoMHZBIrCU0kJgWZwz855+sj4ckzM9eNMhhpgsu5kiyjxk05ZiEr6W
DKAi8FrOH3J7eiu8LHtpYz3LaqCYn22J63hFzAxd0WfETg3Jr9Uo8QnP5UQU
AcdJ2Z/PPAjxIfJglAnEuQZqsgyZMpRHibxkxuEj9+ErzYA+8LJETG6gqjVC
h8Ba7pLNvn/geydL+n/ySKxzo2yV3TqrvPZdRe41g816EgaO8RFucY/TgGkw
f5l7B2zLvxMnAWyCNv5hzq2om4oxHOd2EuwClURya3TrwdtqmUIdW0aj3wNu
U0dk4PhY0ua66lz/kp/BdgsN6nQglj0hqhF9/eonPhdmGXwLfMnWSO07QfnM
HInagvu8eLHzWNjJfuJ61PEDMULEa9jeNc2vNZ/+DBkq2x8t1C70ysKCCWxd
y8T7HcOHnBjNq/BqyqaSI5Y5zZmZzuZSEgw1gNVVExzqbxWqMJSuje9cQqWe
hw8jltB4jbmv8gmZvcnaV2DzqHz4P3yX5Sf7PPAUzlmSTSVMhFmfgYuqHup8
B/zt7C8T6p/v7uKiA7SQmm03CP/XD0j7NE3l6Mx+ZGAVEmiNIEo92mQTO3UB
x8hmk89UL7S39ZPlKm6awxf7m4he2xu4DfWot1GEhrOk1BdpH/I39ON530Pu
Ft+jM+8Us1d/3Eb0AtTsEM+DnZ1NeHjjfPHy+vSsRmB7gOMZVBfHme14gyH8
Nw2I28XRewW/GsS+MjwSFFPhihzkz/9jNoAp01tcZfrzdowm3XS71nl78S23
2zAZeLUE+CqMhSkzTTL8KUfHPFokLkiBhX/0/Pqi7CPDCePsn8XCVui++ESO
EqN0eq8GsUS/gY5IA6bybASxiFaENvhgF60l92Q2FxugNnfU1PdCwVou3X18
I1Dj1R2Wr04rGaalxn3NJcG+PIDxAkZypwBT0w4XXRTMBBG4hHw5fDIYzrHC
aCHQo85C6ISH6+PwAJsKu0TGwgnbAj6KV4SFLwBQhcRhfhowPDGYFCbLBP+r
VZ59rsdpPuKw9x4OHbGuSW47w+ppahliLfcoooRgG/MPDo0AZDh4zBxHGebN
goeuLmnKJqK8Dq9Vfwv2P6A4sdbnzaEcVvoSmirrGdsMkcu8gG1VKUwLjC78
huCPveaFw2Ut8gizXC5ADWKyI2FYA9f2hYkPzKTY41xx4AGz0B3bPhfNag0R
VE6bDU0Mvsn40A1o5XvxBDJtMhjwgq2PZbhvVa4RowYIXyKO1Pv/sJuElSh0
pdFVWiiJ4M6uKFx2CrKy8yQFpCABfs5dacge3cfTEqMkmlf8wkJMrkGOfDD5
4tVCNQO4/czxnCguh9VyU9AqfzWYFm5KjtOUcxbGtS6XfXj5QlsUZQOBws4O
fJMWrIYSSd/NPt7u6g5a4trN70FH14S2bvU530rCzqADE92oN/8SV4ohznVv
EEggdqP1307M2ULHKza5ruCEIrD3NM4FlRAC10ZPVZRgBv8pvePOyYlzB1T6
2ZmFIJVl0161FOQy5LUe+gchoXMmAoqJqZGE8MvDVibT2UG69eJZxYAUCMgt
Ri+GmVxMt4RNjaKvi76Hjv/Ex1mbdftLvXE1iCEocMYbHJKuZcqA7zzo2GPA
QN4tECylNTUjw5BXhBkMwn4HzjRbk6KECmPw3ewF12CYA9nyCOrRY4Q4/ujV
p6zNBe3ZK9VvW1/xpmYTrTHVPSJ4EUNOCjDa1mRQO+lJ3zj8uk4glid0poLx
7rqB5EdqYvwtEC4m98Fc4MYWMP9+mjdJ9eeTBfEKeKPdjRfDmDlbCQMM2/+8
y6BvbrXv+Pb5XL/X87Pv4eaFhm+ox/Q/IwLc0SGAI+YiC1e7WjE08yF/Q3FO
Tat062IIR10LfcD/u4uzI71651nwKim53NlSnVnDG2XJE9YXg6hAJVmjkgID
8P6Er2C9moMluLZgQs5BB91Y9UktVLYw6cInc1K1gmuzedXIAHyl3NIkE0fZ
nkKzDGPJ4qu7/XK9+E2rbMk5k9JaXN550Jp2CjhW3xk1tYuhZ+DYRdYvddtY
kK7ZxxW0PTIT0VzoVqXsPyMbzzaUleOHGp7d2MKUNihst+QOdljwix9wNljc
bbC109jfHe0BkFawxOdj52AFQW5CUXo5utMOJGN8LO+ERja1tCYFlMIMEHIu
eqJIt4MlgGBcEK+YrtcL59NoFLuFYppp7YJfINmVD+iWSoL01rxJOfLENFo/
p7vN4ftTVdvkehFzw5x+UJ6Zq8lLSLyZQwaKZuOS7ckXDjWtQz7srbLMSfC4
ko32zEPvDgKy5V3xjM820QTYrQf4nfxgJy1oTHJpWX8z05RvE3rwvTnTYPLj
HAAF79SOYojWIC/IJ2CfvzDpngG7X9nz0LTC1nhVhf5p8qwl226Lcyve8BYq
WI6+NAqAmKLDJJlMwNyJPjEFRfm8xAmd8amdNhrPvvYD6VW+zHAAja4TrNDM
65gaUyFdwoik0/JcxbW3BzSJ/RcDZ6FGva+6V8Fet8NClDjT2hMvZTRrBp4R
p+KZzlx+8KLyBNa81343rNhoTeOlJwt3AUXxx6hg/wgrKuB2/QqDVg1/AWgD
r31sQAbnhC8hXCkTXmA2rh2ZWrc5dX+O5iafZ0YBcTtuw8mTNmfxNNglPftn
gvS59UeAwEORM0nHIc6FPGHAC0GZ9TbzxRmCSkwGSHZbym1Fd6KOQlciuaM7
goy7sVCxZ4jB1l+NQ6tgvujRVknhiFOXc69uTIvG9JF6iN3ZsGUchXlGwUyN
Mw+dfjnGFVL3FflHYUVidXMWsnOEYgd9HITEX2TskUideLI/jfAXevVzPwVT
Sc+BKOMqsfb1psG08NmU0ON2yzyep3X7HbAb2QsN/nAFUvPdHidV9vIbGb6u
cPmrLmKEZqPoqUzjLQHuosv2RZXnOrGvNN5UDoTj4dcZYBAXx/0r8m6b8Rj0
FeMvQDL+5SAB5zdfTxaOwY18ts2FV7icd6fTzY1o/OwhYSseyaTQWZh0FO3r
Q2HkyvKZhA787p+8DWwFRXy5L2t5oq7mCDUKit6iwJ3iZNbVYgSQ/qjMalYK
tB9qiZLR4A1SFXyw62W18dHqebAYhIeGG0+qn3sLljwCDPHImwwSGbL4kvRL
BWGU6aUBHFPOId67YlpM1jKC5ddaI68fsB6gxNTggAlGdqvCA96UyILI9gUp
/95vclhXNG8WuhXme2ITjUh7WeEVlZVNVN3N3aNwpTkBMinCskUR3g8DmJ5Z
pfgDelAiMAGpZOIEgZ3RFg2JL6RBiT1z5O40vsPEa1szOtJN9V/sCB30zqoA
7AH7MWiAURoJ4Mhc/4v/0dL4jkAuAru/YYeI6kQ2Pewy/lMG3O66g3g+ZhrB
z5j6dADLWtcAS0FHcgd/JWg9zmTU9ZkRnJbCc8SDZkPhSzf5ZIi+6JEl2h/E
Nw8qMfYBLaTZqhxVMUTVD/c5KDRBbZ9TwjjKtbYodCKgbwwM8vQNAiZLOHvV
Y3Gt66sIAfAbohT/Ijjla5HrX8bBfUPE5J8LatjLJTi3HjsUgsR54+U2ej9P
ZhU+cxCQbcaeIrP3zyA1k/tckwVCoruoH4JGOhBhbvgnKTwsapFdfL9KJeVp
793GcbUd/lrgf5tKlzhqVAKQtLwyMpUfU0lrvl7p+lkc3Bu+YZcEXW2M01Lx
4oWjiAofxSoNiHbG+ShwruKUGQ3tGTc21MCQgtPcCjF9s0qGihsuYUr7cmyh
ifr8dUSx7M8dgEf2/gZjI9sEwqmMWfNVA3AubE8Tq4ifralsjNNsdfnhk+wk
7SY89aXtW0vNkjk49Z6pchWUOxMQhaiIM4+6gXd0Os/pmpATdzLI4eWcvQaY
rkc38ShWWr2eV63FIa1U9RRZ5tLQP5U7JhKWkOJcxxnoJfF0YgakW6oeXJrF
usUuBRDXTaLt1K3ZS2yxFZi+oC49QuGBstiWuM96dXI1Jg0x8D/FiBM5D8aR
/oI0OEqSz4nxk43JHXP1gaBSd2nAxJh1PxyF7fxtwH7jf6mZ8lBjIUV+DnvV
A4e5z4/2eijMfe3eAszkJvDJXuBxbTQCBoZD4nioBsktsmZbDecspNBQdRvw
6PHEwpwuXufb6rKUoMgpUIBIsR5S8wOAHDt+rmzLehIWR+rpUWxt0SCyf83D
OESL5yDZmGSW2+AfZR/tQc3zpr6u7Uf3wJrSmnnPbA5F5OB4/3Og/WUQH2fV
sK+147HdxS+b2YKaYDjheFi9APNLNhTqcyxPyo3OhX3YTLQR2Rq+w9UV45jS
o7GgpHnx5IzPWQ2tboH86qgpimU3NTXtvtGtzD8LPdZq8bRwPmhwHpMYPdZg
gL/E01eNdPDGZblPT1gVAQZYRmSBkLi/M8X31keUjhV/uq6NNGeN509c06WQ
VghVWQabeYcIiaI78DBHQLBrKhDaSlf5F2X79ND8+dbS53xXUZf9ydgU/2fh
pzkBPEMcPZp68Yxbd80JoMutHQCZB/ham4dtUL6oLuLYTm6iE7RLyhUcuCbC
GY4+OZhfxTay/QnmsZgxN/aZYWTnSbkodoSwtm4PBh2TA9p9lNO94UFL23W3
9Jv60ISrcW40rJVLAd9yu/roIjJhlKqoUvwuIeF+XTuwC8alL2q+QD5b6Doi
CF9X1JpI39ylsBYmjvwnXfzr76ttHwzwiZniSzq4iH/ge4cnyyetc1WCnaEP
QX0uLXG/RbS3C409gUkyt/wJhKzPPN+DxFUOUu3fQ0LAFJl/EiL4pBBJ1rOj
mQxUg1mSSObYB+fnA2Z2OYyRqhsWwY+M+UDEEHIezBcapFzENAi5aUi/xtUz
mV5F407JqHQz2ZxWNHWhHOuApi7uQu63wxLDsmbJrX68fobLc+XnPyILvXs1
lcx7+zGFIrP4cfIVGAx09Ju+dBKLmOoWnxoJ9oLQHuLoTRtldNe6mztWds7E
od5dIbV1uXZaxPsqPY0MHhEdIQEjPJUi9XfJ1wzZEBxU+u0Lp78pgqYMocGI
oQFA0u04TMT4ubfIEb92lCqAGECCtnwt2D8ioA/0LYB3+zPlmvy/rR+zvtWO
GHEO3QX6YrjAMyQZRCOXxTfr3QxF7LJ/zZwfDg5NgB2g+8p/IgucuRNEEm6w
nYX1TtEnPpdKcOE3fxGaEnhIIqjodEgUyy47oWynPuiJMO4hTgAHhzmgmApB
xXj5rce4qrM8Kq0GU+CRqS1DwrhaFY8ITI5Q5M3OJdrgnKiI6AB8QRpSIiJd
q8LJbswZgVNbJMHkAe5bno67VHslQHz4CNSgLWXcf7a+gM8mQh+K7RhbIacO
vzHOseEYtLwJHeB2aJ4gtihxQPKSo0A1SIF6WRFm3l0piqlHpo1dMyDX2XeF
0q7g46jBAWoZ2czpsWAYyYhGl4dTK3SNG9VboL50ybbYIBdJyrM6jRiMomNf
gt/Gg0tIM8bx0z2YkRHp9fPgvwnkpGSkT5ifVPFCvLaARjRscdEr7uSJLux2
EE7yTr1sh3TqfDapb3zdxqhykr+Zfw+2oOFj6uW8I5KSwVm78Gd+P07HS45Z
VYj4pzyY8sxNFx5spRjQ9UgNkrpk1oSrUzDQmdeLTNGXUZI3cJQVaEfBCu+F
Aoe7v/ZHPv1wKLL9DOEdOFZx1KgXby+rqe2dnDvq/TMFTVvqURiMBUudk662
hgJseqg/6tO/2q/LbNy1hcCxloFECw9ChJp9qICFV+q+aXLZbCJ6Eku8vdOT
Ji6fkWZM1GHdXwnaxoNpe0gMqs5VOwUHXXyeeIjAmhZMXinXhM9twonZj3hP
uriM8Mnq4mRZgDC/UBHcdcciAoboLwNsZOzmROOgS4y526YFf8Mp9Us+vyie
BTzl1Lva30zANxKrSfGYadEV/8hOOSjUt5UTVmhzlVznB0B6KmmGYaEL/06R
nfLbzF3XE2csj/17GUjiZltYXlsuoNUeVPAaTrZTzj9q8G1JRxxzZuPhice3
dOQh8skY2ND997u7jXw/yKFD0Ck1c7iCokUt+utRxUlWHM75bobip42iudVc
dQaCRsj124pb+e8yyBnhdHqHpAAGIM1lipRSD7Q1fH7/TU6bwKSw6gTzrfVf
vXNtg+GSJ9Pq/a3Twj8v5EKisjn/ctK3OA+VVvsGOt8TTGWTUepgG7Bxjs3z
4d6HeQ4qPRQbEDQJIwrndOBNIyPe7a7VOrQy/AAVdFTfOBAtNeLP7EDZdoXx
yqPgrHCyoUA0V7nshVHEQUTge4k67NatyfKSuI7VTq6Q42EXRY3CcAg/QOZM
FvqyaOHsr6Rf5NTgRmMh/sC2NwgbC6CMhRMw6L1pHMmv+684Z6+AyPL6HoBx
ryBK5eOINAW6w7l8BNUmzTdYF5XzBpCcGM2Fa+n/y7u0MHFEHBuuuT1HYQvB
IHizx07b4LBcQvEK/e5UIK3LeAgnHMS8TBx/aDnq4h37mH834yykvrn0o04A
wVXySi/w57AGagVupSdJdOskvbzPqEpH/7HQXYdx/Sx0I9UTx0LlogUHnP8T
T/G94FwtW5DXUjuYovoY0R+mTqsahs0Nk4fZoSL7JA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "221cqLfSQtZLwpVKjUxAj0azxWo9qWyTHel1yyBq9riDaTa7pjyEaEdGOLLz3wcrK5rHulca0g1g9Zlx/VJp3su79bVOdFJFOSZrof0/9wf6C4nAWrw+2PgJSzMMKpaFLO6gpDFruW5083aTh1M+Q5KnW16yLzHWGhpxtWHi5x5kzslfPRMwe4HyZUYh8/FwJanr1Um2jvkSaUjUKvojtHUTdbUpkWg93bqHvMIamsn0Iizf7esmpkf54G/62RFkdyZ2BdNRUrDkRE3oj5Cyy38/xnBH8PzZZCTfYbczWn8gsnVDYqJdh93I+m8XvV2is0Hm6fS/erTJRC4sW2DUHKA4l1cPfT7szFwXKbfp/hVrf6WtKBr/rh5qu2BGqzWC3Sx12nPFbrdx8YFkthL0ZYGgQka+oEdD5IyJ1y+ACwh4kWq0X+CC8HnWe1OURNktw6EAVmtOgxhqLK/qyuIo7doI/943lILVa2bqgQMwV1PoPA64cI1Y3AObgaVeWc0rsxFS7IYKcNXCvuHin5czOPfEcZ4Dbn43BhO+ALu/uEc7LI4RimEuk50AZF5fEltPz9y9Qd16d7mGfVJUJnmclP/npI+hEIxUrlsQZYsFhcloeTjPAy1snAk324MNzBFUxoodcPTBzCLh6xXoy/BonWZCfezpHtyay9Ccm9Ry7lac1VzdXk130Bpi9V6zETRlS07KGrPIvDLUJvpJbRFyRPdr01Ef3Z1BSiqOLNSyczPd3zco0eNqm/5U2ZUqDCDjbN7eaf8Xl4quD0NzbhSZEyXE5At6s8Kr09IJd9QYRlXiOE8AwbMjbb53+QSaAJcPorVGsupSUZEfpI6buWcn1ZbXFVuFZFC/G+crOxlpy/JDun2KSiy/0O5s24UWK/E6R9spWB8fZAu0fjBWkDWaHH1+GgEKbw0CB3CCUaC+Thn8GI6uiMtYv4h8IbWw483mWAldBQfAbWz3THb71IjVHQB4Ukbcq9+eV1JqnpMhEJnjQy8F1wYfkzkVwhhWTdJH"
`endif