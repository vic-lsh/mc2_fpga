// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
wELXrEpJJvS3zXyB43jxVvmHNvwtXTUK8VLpb5zlQlQaQvbrV6P+xAHVoadM
IKNEDWloG2gQ26vqxh69tO2p4dgLNKHwJuSJpAeFrO7/Rt5119Jlx39ZuNkV
81xfn93QKCCk73QsAMVQUkM41ppJmgsH5WTbKTHL0WqCrwHMHyo1nttetsC5
f1kua9UwpWTHcS8FSRZ1Uwomb69OcYgRXqypij3XdjNhu8qdoQ5rUBqjtWsu
DDHxmMlrpgfEFX/XQSvC+XywJBTuZrAprRuW26fZ/AiRCkbQT/aJx4shlrpo
cdN6ybULsMJUWzXoA2lPMLcvInSjROxkS+KyJa8ACw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ATbT/6mpKJ5xz4t90C6DzEV+FI08dw+Jt8DQfFyamfwx06PMEtWrHWtMY80I
ePYDnxGDFBKcqTE8rIetHsbSCicpDkGmVWmMTynYcsny666z05CEqihgCMX3
hAymK2+lWsnPd0+/hZv5G0wX7MEBk7AklS04s+jFf0QI5dcbFnMolA91bSWv
gd2LEg2/99hBjYiMIDvEvd6k2rduXqdT6nVGs1SSMYeKpVL+1Pxaxf4oAIr2
/cQYNAMYRZMSBCgicaWBgC6HDg8DSXSjn10f60KSaSuTJPiC+C6zNSf5+4DF
0viOqus4fVZZgv5Cig0mERDsnAI3WCp7yyjCJxWLtg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
tVuoaSRvdLk/OVJsqrWAk1U+QTRIkbuQkQm86zLX/x2fxx1FZENA82Uc+50m
rhkwgd3TWZyPjYKjTFlEiNehSjLPU5LDylp0Ahuiz4uKX+L3WubDAZs8AZyy
5euTewf8gE0k/iOvfC9zAhN7UhLClVuydpFyrVfaGtAWbsjS5rRJnIJh+eUR
fcxSrx8q1M7PTe4b7pP9RkxlnswD9T+Am2cjcXgOWxtNA864gMSO2UPg15xf
h3lDgaH9wB3TsU8fKHLwgLmxIKre16EHGNOp7XHoAFq7n+HuBCb49J1t1Ams
OoeYw442+m5/CeELtppKcooigz0FsQT/OyNOMdmJoQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ze6INNMNjCX3yZR/9DigivjnUAQnFYiuD3FDC27nY95tA41usfGBZXi1J4U8
rx3UV9pHhoMX1ZM4JAd+u/yccX2NS/hZjAL8W5KTaVOHMys0gnxFjujyHfXx
rAyXyVukQQdgx29CLYxwuaaZdradKpFIPm2INpGlmH116BW0ecE+sRIF4Kae
iUKtPzmSK6Lkqix7CuaJQq0EbrOpyrd1BbWV9gLUwbsCgchBDqE5ejUTkQcw
kmcowIoGmSSRotf80MX5zZ2dZ8tXwEUyeYJHcKqXlNYKaACkLP1sDaGsSAu3
i5ImZHkOMSCbDUgUM3m1+3sijDzc8bmnA7nCaY3f5A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cHRwo58VrvrtGynzNHKKIcgbH88Sd2tuJQ9fgCsmXZrKjxT7Lm2yUQ9uxMYW
BIUYY/aULz6kyzWDnq/ztkZqRTG4pbupk2BgdPfSCSl27eCP4p2OGzWAbc1z
6SWjUhZhFfa6EKM0BeOrfErqRdSw1x1nQhK1W1xaIsPRJNrVy3o=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
SiDUdH5eyK8N/QitQ+BUl/MlRVKU6p59Mjs5bJDO/7/gY5hyxYlyXBZsUB7g
jiVXcUy6zfBWZyUhqWTRC4xpG+bL+EyUHZLt/1NGapSybpcze74ZNL2wtm4P
PR6dqehRYWMwJKYGpCxxxgI7LEz8QSyfz59FPmD5lxdN6pAQh7ywaH+h4VGd
w/pm4XjMgCZrttB9URJKR65JBgMq5/Qhb6+XQz+LupbahnRC/QFkDJjOkbep
jOXuNN896pP4wd4a1loulZfB32cw1r/c6d9VGBlwTmWss7/9m53faRR+/v8d
KunL4qwssb2UeFdjNeYYrhfX8uQZaoad7FOmZ0a2/ggFX8xqdI9LJ2U7z5Sg
tRg3ph95tzVyRrMgQR1MpOrKR9fLKp9PnYiSfrtH7WOpuKERqZ/qaeo419XQ
pAcATxKgh+UJkqeuMtOHSBn0oPcLORu2UhmAUQtujUAFyuUAT9KwcmpHjow5
/KnnAnYQDSuV//sSJGIwwN5n45qxVEQ1


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LQb50R1Knf3HdyV1Pc6l9DJiHcjdagsFIDSbxezzIC5TqwHdIFbaHDCtjXLS
koQghHgifVARYKvYz3DpVHSk8mA34PInWBgiQCRSm6QGmnuH3hYIp6BKhQmk
4kchvSt5mq+apsRTPzSg6fJUGvEl0uc5OG67Z13i3VMjsZNI9ik=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nU9tCzXDF0TIg/RfnJNzl8/w/S4h4/SyTz6W9QHAF4aGgzs3+V7rVKcXFu1d
wkKf96auszzQSvfmRhC/0jlp1vGhK6Qr9jbK+tgPAXwyICNpjSJDYvI/bcIL
siYDfrfjQOyDUUzTcGxUNifqJYhz49WL6xhC++RG4KgOJRFQVYg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 46352)
`pragma protect data_block
7OkArHdEmfJ3UnXm5cjmDarB9YSJ3mArlw/ZQmNsM/gOCsxXFf/wqmFp5dM6
JO1N02hcqC28fgNYbc6xvq3Y5dSHWquHDYdLz2CpkJnYpc88B5ZxKGapAvEy
OWVgAxGJqeTZRmWVCHuR8ImbvpF3ypekYv+ZOg//rshPzer/jK3Zvc0x9qvm
R3i5cCB1onbYupICgmToon4y8I6I7MYStpfCErifNghYzmWb8Oa5FStDkwNN
euviq3VeBpy8mjfFWApOUAF5qKbJkyDgfV0u0mCMs076KIhH/9fzHTyeOCnZ
kEzYAuN+TN5K/rOcGO1/wmTI6y7qTn7/aGtczCyLjNx/EVYN4Jz7aBM5Rfy+
ElROegW2V0cHGFacKd8Y1kULepYwZv2FFxEBnb30WL34V81wkx0veNC8X/wz
jwcxMprWgpXh2mDx5u80Txh3hM6frTKhbN34jwstJGCn9LE7DxqKC4NWWZnM
paECmHBHePfAoRXY5rIJcoaGopwXTRBJhGpIWi7+8KBi5gR5tIl1c6bdSANb
e4iO5z23GvAyN5QtlYFR5ubsqh8BZ3HK+61Sx+4hpo23qaQIh5NgA63YEUZH
qNz/YzkvrRQySEv+lnTyMDW7MTR6dzXeWob0efn4r03MFp70hZIZAZ9rr994
bW5LnDyEQ0yTjMSi/TdGq89frP6mNj1reA3hJhoEBjj35GfsXtApD3w02eZT
kZMaaIm6GyhXG8FXA+rtKlXUbz3l5O2ioR1DRF7/xo7SwNoS52UL9fJckAM5
yCfeqdE3AbmMtlhj2r03TI07y00EpVvoB4VdAsjhzXgg8V/IViN3M4YvpXGn
o2pN+hkgHRAc6Yku5eAXxGbIqF8oIGWK0i9rD6N0arDCi0gbBbj326FP07Tu
DL2zerZBzyvBFpqSsSuc6fB8NZNg8ZSzQlmIZFG6WZPaH4GLtN+FJ+RP0Qnu
3L/ga3eDomNUhnbfxCaFeZMB2aTw31MzjTFnOeWeCAq48W1r0klWMG6eJw2k
ui9FS6EP2Njj/PKCWCkQW6NsOfq1930Ik6Zgk7MjJParhKr1m6NgETGOS7WT
kxu/kO8totszKa8RmTpQ84iXgsBbQVKT+gOocfGL9eCPRblRQ+0R3OWHs1pi
6oxJs3x5jtrtiOlKhRDbUEE9uLT5d2JJCWhpCzD279bxMaQfjdpM+qkyGYk1
NOU2ADNrTEo2WV/JH79k5pJPkKOpV6ZdAiITbnaix31pCwsWZrRtsQ47F2Fp
j4FrvEamrrZ6UgmZuco1v/DPhHoSS18auPW7aBGzTtJqGt67JW+Lp0nab2o+
7y5j9U1o4xT2plmEB/ksRFIJq8NKlOpzEowjg3fWAgCmKY7Hy0AEd+xQ3rwg
htMA96PgukdJ2s06CUVfN1w0+rpsxd5eVJNb0QAKO0M3r/+lI5LeuIxSlOFB
eklU0Ci1KkEedn2LL+ZCkx+2XEfgba8EPJhJXlJZnClI+H5XBqMzkGjMz2uj
htGERKnowzpmgL1vv6i3DMt5I8EHyL8ovsaKRZYJE4WqD58KYjQ+xBd2Vd33
9FQWM35ccbMJDReYsECQappkgCs3qhtWEwvPzXINe8+a7GcekUG8WYqGwR6c
vYot+B9kVzTGE1bDZU0hpjB3idcyhhFxeohGaCjWjv6SW+rjIfkuXPiP39mh
ub+O21y4n2FOYMB1U6qoTtqXUa3KkKF3JX/R6Y8cEQPCHY6lPsJ/PhEfM4xi
wK+WlkZyRNz5nj9QBvAAq+UYMccErv501mAtzjMeR2iX5wAdG/84KHP92+jE
np4xUBGBvWDE6Mr0pMjlBZALOU2s/bZV4Jc0T1uTSeEcNr8zEQZR1ukTR/H9
RUqulLU5jnHkPRkBJaZFBgFsUoc6LVje0Dn3zR9xwn5+R9PcRddRUQYVA33q
3qCneCXd+qPaOsT/L7/57AL1gwRev+NfHuYf5Tkm94ftUNmct7QHY3z3iGDp
+R0yjVtjLsRcnQz6utE2/1jVJ8N/7UzRWNMcirl3PQA8TEzTB6nObSdRRLPN
6SVinvt9PIxNYX1s0qrsIfMGAMj380R4eDB8S7O5QguaqG4fP3ogfVRnWYnh
/PVhYrIVTVo1WkZGf82FOJXYWnvTSvDWErBrT74iX1iYy+sfKIMkDnyL7man
DjVWsME79F+kwvv5yJNZ8z+Tg0Euct6gqxcbKmKLboLY6tJWtn8fpZArT2ZU
iQMEmbTvhYhNCmRNKqZAXU6ujHzwjadOVOjVFP6jAzWzYdkKx2DmlCLckoxW
B7KcFRivcWN/86/npUYDPDZ1Dn/cV8f7cRqZGvY3vvdCU0XhxxQnl6Ss5R56
GFQ3yWBfKqr4BoVZiIM4JNOJDHV31JyJvXJ97O4avvwKQduob0MW6+xW+MR4
z9LHzgEaHv+Iw7ft7bBOtyo+25OFaLUDe/w5foPtWZh6b+eGMPGP1UxZ/QfP
l735OZDsBfO/W3rHnsRK8pPthTzqjcPTvJq93pR6UiOgnYCMJnlX3NoTLkVq
ceIPRkkgtgiice+DoQLuVBiT8yTFMUR4v+nXyp1gYGi8KOSJ0KhV0WvRU0Ot
18C5Pjkv8+iQzPHLPNcCsmotxNWDQJg7QiFTCwAP1/JxrBfJiHCWXSBB1pUv
iOdy9EhJE/OsePEH0+kl/JNMOI3XC26SqeXOguG9jANPw3Lc2rlOy4El1jgh
mvObJyiewId7CjcTjyfgLguG2pZFGqbWLk86SuOjWHyocYLFPLTEG2MqzaBx
t1c8b58VpcYFfZUkEEfOlvKi0O3/J2JNSkv77X3QFxBn1ulWFmSVTUhoiwCI
DSItPhlN2LCq+Zb2J72bAR2piYH1ntBWPZ+4eYSy6TfKYpSoho9BPoFQvCzc
9kTgkY8kbNTp7nQCa6/e31foLfF8CwNvgivPMZE4sqPEDikn7k4ppnYqcnsY
NiLsHlzsGZ6UusExar34wEdmpzpnqEnDNg+PzPYq70fCy1KZuwzA2AZfN7WC
j8X3kqnuLLQTe48QtzrotH5RCIJEo37lURj2ks+hJ5DK09HDQL6OhJUmcBFM
wAuwx0UvhBWDYTJUL1H30/E5Jm1zkrV9j1XClA6iTLn1scKFZiTJNOj79hgV
2C0ITNYyZfivceOuKbO5lqblBqotXSHhfTXutz/NcyIzp5IuAaW3LNzlP4/P
5nQAuleunsGJjYNWGbsuvs822GUiVR1t/5u0GEBIxc6PKlT9wYnlOBrY8Iu8
vMNiS99iYcpGCzZOsP3uBnKte5Q74LHWwWrnHprTGTPXHvf9pBBGD6Lqfnda
ShBM79mZm8kqpSagocg18xE4mtSBu5di/y4BWAguq/nx9NRFrrDOAeo/4yFI
rT96toF/T9QRhPAWLFWz0rg7U1d7gGYXEo6h39e7TBRff1q8sUAxMeNjd4bn
as0n6e3fzM2gg3aYBveqWgUU6tVU7ZDR4W/ujweqAy1A5tiac4Dk5bd5xkJO
7LXf1L1dg1k7KnyC0pJROJmBaDc4cXXIwt65Z2qGGBuFstwrILCAnezmdhHK
VkBVVGIvoym4EHNqXgmpZNAyhdbWb7XJPimvf77dVmklguzp107yVwJuIyBG
xI6WmEcz12MTAIhhCQOf03CcnzOCxNWA1y3ZovuM6fonoU9cOzuzucF4Gi5b
cvo3cqKABvHxocCfQDuRTwWyzVtGafRYQJJeESZ7BQGpfr57PKQRz8U+oT3a
78m1265Yh6eklsxd8zj1LK0d1YVVKsU1+h5vOYD5tpUEVe28BLwHOOa4JrA0
20lInE1l9KPCZu4ANGqdN/5/UDQCVjeKdKrIkwbAkXPGUL2FXoJJvH2cqy0w
Uw7FK9BELBWtJH6RByOLI1CNwDeX0iAj3K74uWUakZH/vTd1hYY30sHeqYpZ
K8PJwnNsZ6bJDjnxNfpyAOn3HSLk5y5M/d6zNCvOUHO8QW0qZnEp6cbR+Hdu
ooq6fr8dxCd2pd7iTtLiv8G91ZcNcB1IDOR8FBW8vX7NSjsQzjruYgEuL1pB
MOeyfVWTRRdcIIdVEf6ENJB0Dq3McZiUb5yKHaImLYHAUkw2IhCPh2/4EMxl
fql3IH+eSuugS0ZeaDhhkroRvp/7xzhQm+5smjIqJgJtg+uMpYcgRuGiJQwn
FFqa5sPnXPEA9KhdmWdrZxMF1OGVeNaalnaufTeLtSTAwXwQACrQJVKTI1kw
nmEaw77i0S8SrHsSZvIu1BfJUpjICGYNQ2LKOd4TiCesxjhZwAroPq+suH87
T5Z9O9fEZ8Mvz0iImocGLpepL2aZoWzqjG00zc6VDVVD0tqEnjz17VkuzuEy
WbzjZirWlw1wpZ1MqOc+rAKyyreDmge+nA9sbY7LAbTY3mvpdMTWboRYtZgF
7q8neUhPk9aTWh+qMN4frXaMDU7waevSyFDIiZ+IkILAWmQPlwx/ralsIyce
Cj5RqDZGYn1b+qodURlsgknyd68bbvoqMr7kSNA9TWAk+JWl1eKj2SG9NkWs
BXsHbdkAQj274p6G7HkT5eBAURA4QDc+KwMse5/4UYKlLE88Sw5bSEOF8D2q
cespkPK9lLY6TyDgEuKYq0BP0f/9/hI8Y3PDGLqBqwx48JiEOwJGyWwMBOZX
eQGxecrDuJXA+Y1FcTjHTRrdFowQYtsx0FXFLxaIALLIQAqj/rTNnZgCT96C
f1FcB+ZVcKkEPGSIENTfqakPXbaa26gto8OeLvA9dnXw4h24ywpGr4RL9rOO
hPRqq0iN/mDS2NTuMce/gV4Z64FcywyurmaSzOyy0Atfev6Ykj96KeEPEcha
5T0p+X8h070zmxCgRsoYL/BjGL5tRe0/sPusWVxlW/bJC//K5YZep/QmuIse
eXTTUU2tU4zy7uANhjvqLSvWabLJJ1CclcCouWAnFVHE/ndCJOUwlNrb9SwP
Nk8j9cubpyVwf5iM7QDb7grpLllUGyEWSxXHXLTSc8W7NMe9yhfE58Rb2Hbl
T2L6QBXcK32gZnCFokbsVm6cscfX6wtC6vGrZYx74r6QTx98ibSZoDdSVnLf
UhpPTaty1gtb/nqvMULdAa9CiKVgleeti6chKpuZBxHYA3UNjpF3AGMXERkR
nliTYDOYmy1WCXjxjsWg3eJgzlJHkEJj3SVtaocVKA8dFOQxpKzb3NfNYAbN
5DarOVT5WNqMOO3oxfu46s4+f0QN9rhf+mSp2qn7NO8V7WfNhUc6GXe5ZnrL
/4O3uG3vEdadxSfkIawO1pu3zN0GkccXGiTXkM/2WcKQgo9xaRVBGoxkeQ1j
dLzhCNHalF7Jw4+U6NPVb31RGgcULKkW1GriX6laGcWm7wRYRBbHRut4I5DW
k4fPfpiGTwk39YPH6/7ZCyU0clDubrpo2496fLoQy56n2fVX23XxeV/H2KzJ
+2/0VGYg4FjfWZtLNIxwbaz8IeMUo+ZCV94tHRohd3vwUo6QQVAmkdfU6Yge
iRfwdEfPLxBzZtIeo3K63eOYosu1DaJFdDEA811BFgUKML7M/hlQHAWh35/K
2VfMDy1TK8abVHCaq2lSIwZAYDrfRcRhXbjzInjXmlcGemQ1GI3Ats3cDo1X
UpWwxsQGD27WkPQfJc+HBdAK76twcs4M9kQzY7BgDoqKJrHoOvMzLsWPLEC5
c5rMhvgNE0oRWqQKrbs1Fnv8EhLIBF3LiSQtb7pyuhmnz+kDguKadHhAl/2e
TJyiSHv4SgXb35R9iJRChNGjTP9pUJigpNXddLYEUm5kO/DdSZlyVvaYt0Wp
bJT1LMKVHrdpOzJnk2WM08Y17z8alZkOK+6Jj31A5JUD92njxbasqIGOMKKy
ohcg5JmmYjAIh5ixjKxorX8uyXeFJngC0RRTYfXjmNo53v66OC/bKj/7CATZ
l6YFvMEqU5ajyRt6rgNF+EcJMgJSytFBYQKfQHRv3G7EjikyhMwkx70gGMD3
phY70jy2sFy1fCbk9LVrosPeVZx5yJfBiox3xWyUcyZglPnBVR+87r04FG9G
OPl+2jTL64pDJ/vZRtr1uco0o/6fd1jZBpFC+VMIRJHLkv4wx8hNF+rb0opO
CHR5slM9yPq/KLvMHiLl54YEO4HrqlG4fp1LeH2IMb2vMddOnbcsyPHQuh5p
bVFRzVxpIsnoItGqNRcVIBYoJqxX8q5i7btkqRhibZbJnA3ZwWd3BD7p/fPQ
a0cRH+h2GtjMH3+tHeDGteL15pDaUTiZzDOBhI7asDH2yL1xiCbCa/cfiaMn
VCL/iYw0iJhHsRUlbmCMsNO93TFnwNgEM6sduWPCddv8hfARq5I18RHZR/IF
e4jMG+NflL6MM4EJSDVullnL7ZG2lTQ89lwmqXAPzHClrzZHdKwTkdmnCp2a
FHg5EqHKdtJqBaarfrntjXyf/RaOe4fgmov69Hf/RNGp2tkxEMN23Ufpzwy0
KTiO7593HqNzGSb+gD5l4Z+LHsQJi9735roi6DBztxvgCqRXk9X4lvMQh0f3
BxIFz1nt5792D47alRYpUMNLRPUSMRF2vz/vzUMq96YLqH1uRIh0Y9Tylaq+
jcBBkKteLUy5CQ522fBNaeYARRB76B7ewss9/8vX+pY8bMiUInPWK/7fW5Ju
amqhwFWdQ6FZV6eI0o6pMOb6/LN+KXlofX7agBd9OplDJA+ld52uyhcVdOBk
O0/aU7PxQPThdBpIc7xUadGN6I/6+3zPiVhgejD6R4GqD3BF7FEwbYg0O4RQ
EzxDf6DoN8AVRrtRpx7glzCVYIcc8oS0mEpY963CFdtw2q6OPIZt66R9tus6
ZedJOvodp2AhoABPGBewE/Lc2zCnY+qYRnaP9ZfjAGb1r6C2yfyr88Cpjdo1
xcw2caOMKU3z9EkuRstXHHrvvp4UHQTDKIm+a+/vGf1qRF/8aIJlGPlFEaXV
Aidq0RU4jhfnyeKM/1KSnjxNydMEPGKhkhlhDqvX4lPAWvMgJGadOgV6fg1T
cwNLmEkJjgyXnXOQlvRMSrbCFtPPeyGn5kAYCnu77Ify15MlstoW7Ck9/bvJ
yHXpIfoK0RRwP7mvgMri5vsgFSC8IcsxFDkSpRENmPkucy9TCpJe0+Lz2Gws
qYbG8Z+rruywxnbC0X9guy8Y9Dhr/DH4SJuK6utTwkFGTUNZJQCivBH7RpwN
QjETakewjpGM892D8ySwH26x/fe5MOiN/ueab3rSbEO1M372JmqGxHqPxwhB
kguf/4RBsuh9gMpTQ7VFcPxorqZh2JcH9jNUHHOX0Ut21tL1OHMTfl7cN2ZP
2UeMMV04e19KFgwMKibCJCS62W6pLnUPazwizA4/y2MCuXqQ+Eq/sA93A14e
YgFl+7DWmWkuFc80yGRjnTP2scUPqZefaXBDmo9s3NJNvrW80dsIW0LzbseA
ZuOLxpObmLQgr3YgZusKGC95ZLpNeaTB3khYs10lLoAz+AS8R6YkGVf3iQC1
h/lHXYYc/siFIOizxhkcMITMxV11HOLcGxlPqEqp7OvJzCq/xV9jQPFHsK1d
i41f7zGGpwPsAZwVQ4AHF9F4fiRS32IuHtysLbVQiw5IhLWg6yBBAjBHt/Ew
OaRv0w6ZIP0vphEmXfQ1rrIYxfGSSfq0P9NXVmApVv0vVvHeqQQe8vIq9ava
DaQ0cVDtxCzYKlZTw+Z1LMmZfSAPQIwsvUZO6/xrOoivO9RgDFk1LQnRfKiq
tR9PhzP+nJGh8P92n1mOJ18NGZ8S2/gJI4K77z6Q65cCgYG2wSe6+6xIc0gt
TxSq0WzCzZXI/CLfhqSQRaEXI7535Wdh+vNb0mOoGXXopthm1/q5rJYijwYe
b5rwMp+xbhAbR9cIBYV7fuT9h6+nKAW27WX9AgUjeymtJ+5H4tQDeOPISzOE
tCPNUxWvli6wfu+W8XEeEUveHn4KmmQySHNa+IxWzxDmAAOnLbsnqMp6copx
tCog+D+BBc3aSjvdxUW1X1GAoCJYD2j258dT3tC0IkrtfCTXoQ7vw25KW1IQ
YMDvpmSsCJsHjpqsi2rfMHIy8c+FCfPgWB+Blxjl3xm5bbBg6iNfRBXIbIX7
4evMoiS6exySKBO/0lq2YxjA0nC10DVozydydwDWwnjCQ5WKt01X0mQWE67e
wwAeOfvRGAc4K1t+pn8FZ3lmqVRLJ2Y/4yz/XUmqE2LbqjOqI+t2X7isaBoX
AzpVCWkMu+zKxMDCIi9KOVkHUPNpICrQZiL9H2DjX6RaZece0ATh7x5xLOIZ
FwU11hdSNmOvo2tGFYIl9Bl4GkC5sVg2SXeI4QIAGwm0vBzt4IeK+jkRGakK
SbeFXW6zq6veq1SxLfZKxlMPgZSbRQGVehSR1W/es6pqmMuXWTfRLbb5ktIJ
2zgfwhjv/e2A0ld9EpPXeVzSRyZmmNEHMGmGwCyo50kGFyYpxXHh5KckgWG1
F8eCC8/1XHZsPUV+y9Pqdp2XDKz4WyXzo0SIeCJJ8R4D6OuXu1TplUrloz8u
gC7YQfaqZ6KLtr3/fVxZnb/A9O1jQXoYqCts95SBI3902HevzVd7/S58uhQK
2dOnWOua1N5v95dCC7b3vQUVtI7Ho/Bxw4URYk+mtA6+AicqSSNOhvaq/MRI
yeJuVDH1Cj3/+ziN1/yKfj6sjAXLVFm1p6szmDnyoARHFqvBdq1eYV7MBOny
1rPVJsx/6+piozrdZ0GDqmPqEdmaZmpqnG3Itg6++UowvfuXz25Wnqc6RQ0c
H8lvIrrlyxeWXKjU/gb1ZtG+nCTZ3blQ/ieNg8wNkCYCpJLj7yk5NvrNfUUi
RRYzGIVSTbQ6BLhSgfUK8WnwPFvAOef/qfQZrqEbcySakJjC9nWFlYOkx5gV
EQKl/JG0e6PC1ndmmGA3VR8g+TQPttjo6XqMN+otfc7NqvUD9coh9+txPfYV
HgectPG2bhSdiXFpEmiqaxBLlWOwxihQ5Edg107m3Ax44fGBWd/vOpz6ffEc
03P2/pjr2xtYhFffFVrOkeKeNBojODg9hDICFFuscoHKCWO1poozKj/jaAt+
HOpJEgWNKjBUE4zdruQ7edFiwutmw0lXhgb425vzutrxW0fI/XReDCmr+02R
bFXn8ZTigO1Zv6BClpmF/tNPOZApiq918m97cwM2lYzH5L8pcBg3dJS8XoXl
8vbjrLvGNlsd52zmCIGC4Q+0U1DKoet4Eo/SgwTAWNg9XPYE1qJeJw1KuPr0
t37vIGO6x6wa8u8dGS3vVGACvl3cN9Jto+gBuGu2Sf1T1PmvMudDnXP80I5U
MV5/XDLA7NJCijR5GkRCxIcwmx/LeP3L7lMRRCJTogPKIRmZOfRe9TUrIRDc
zTq+94YNacWtyokj5JSzAHWa/CHRgLQQaJiLoqYFhdkbkD9LiR5IqAZZD6+J
6QnwAw8p8wV6KsaCD1miA6I/rKLuKa9oS/rzUJxSU3XTJ+/rR/TqfCjCgi4R
0OXKH0UjVgNpKoKIKadpnASAcVKPEmVbj6l46/h7HkNBKDUphbyMZmGZTshW
g2qcykjWXSs/Jg+2LeEkhW8hxtjz4q242TKf/FKianNdfxOzZmnZigY0tdUP
QnGaTEYioHYxxlLFvjAHBoTGrWTKJ+ZyATSOZwGpFVAMNf8mz0cDQ98J/fS5
abvyynPHGcSPUJfLiARCfd8nP3X7mtEQ8hBoC5tINspK+NS5AwMFDbWxBEvc
0n1SNsoE+SWadfW1Euht02iLSOy70behBS2OjExOG2bsQ23OUQjHgINL98cX
GzQN4YbFUVs5xv6MPA72J/YG4JXVHwZCWbR/xU98K4bStvGespoiE8eXmiQx
Uj7PBTNI8gKSRvE6UCGN84UJ/FyBcJ11xj2KxY6ELxujKJ0O2Esv2X2kO7m6
J7+7QO4c43D6RvNgDL5cBr4G1t4jc9o9gqUQ5NOd0w3zjPucf59keYDC5lNX
Xj3G23vuYrvSSEg+/xiVxQP91wETDxFradLxqy70kGGyoqazPw0VmY6fRU5r
SIBeMMAnAdPaOQkTpT/Id36TFYFaugjSUzUgHb1joCfD90OqKuTe7p18XZTV
rcqiVNDDIq5wIzkSSqLSDW+70gZtZP9hjnK9dcakz0a7PbIWc6AwaRAzw+Yz
GZuKANRIpLVES3Gt7ZTbjdeVSLkoV6rkVv7gZNXv80RII5+bQM2QCDPBI7Xo
AHfaD6fs8fmKMSKQAZQN0tQMZ0sN9S8D0HQA9silZ2s9SaityS7MgUPXGMyY
B5wn4/W8gZZAaFgl2/0yhyl+9k1LSGXQEdcyLibMPNe3TZ93SoscgwUfoyUb
eS41PSysVrWwd3NAH0uHXtjzu7BlvEfvBgoK+1FdaljiNSj9AdGqdaN+1cvX
s2R7EyQXAaLPxKvzqHWyf8AWP9jSHSc+Z7vje7mtprpZyZPgq2e5XIeHXW6B
O31n2lGIH67vjtVrl2qc6mKpWclIQs2KHL2v2RSAIgTnMc6qNtR3cqyZHj+2
hDPgBL/rxgmjYyuNA2clWMA2ryzYKWngD8wRBVDjwfC+TgoryrOBTAtQOujv
9GjD1luUiF8W5IPY8s2RiaJOm2L1N6Qqv9P0Eck4vAyvmh9y9Psg4UuW+dEJ
MJWt2fdeV20vq+tCCqddrBtsgxT+IJEoQzf/fBXje4pfyjnrKoB+7Bd8C+Et
x81N/kCiyvcz9Tz6ALCT+GmeuaaqVeZw6nn9X8MGQyh377OQXmuaOTTAposm
zfEZT9GhLB2tqavqbpDvWC4GT+2NpvoCyaj9/4NZbZVirWTrYJtbH8szA9Ry
uq7FYZ2t1Ez8rq33XqEgciyD6xHFShrkX9rZ1PRsvhZAhxgS8SBeQ+OI8gp/
lKAQ3cteJOsmq5wXOWuQR5AD9hWCg2H4ehAn/W3YLFeY3jSMgdaoFSvz5Dos
USRuSk++yCA+gOV+wWN/M5AyQlSVbTO2W2yhTAimEg6u6iPnCaEYxLPmuZC9
SmU3reCJD07zLx35D8OttDuy11WJtLybg6hDDvJs+wARmC4RVPcIXTP817uw
79n9qkXNrGdRm2NnC/1OD0pxpPLWlKOq+z79uMlJxXCAY8G6pWh6/NH877ln
lm0JzWjEsaEqsWIVSh9xveoF6hAAdVuKFJiHSRMLt0yAWrd9rxh+K23sZKYP
N7eaLy/mBwdivjHFuHcy5X9iJyWbKvOEMfj4VN6CDhjT19W4CaMugqmenFH5
SeO1rN192zoVYgyECHbnzkkrmiLUvPZWlevgW0GUXWNf8ruoKLU8JO2OejeW
fjaiDc6TEWX/W0MteC62tZC0wB46jRY/iGpmw0pky7VEvNqFqE5o3bK4CP2w
ihgmGRaxNyKtb5OPQVQjpmtIbeT77WqDxfpWfswM6JGgXP3rNswsDQWGOlIA
Ax/We4qhYmad7YxLdGDeA5BjCyIvpEqZkHc6JhLC56qHz9zX7C8y+YhYyhcK
+AXE+3ESJs7qzJU+1wehHqv4d8KIF6zoLKxufOUHODSYai6wqySpI1Lwc05Q
niV9uf21gCb3oFcQWNek9S2L+q0i7L/nSxwrSRzzXA7l/I4OrNHcgaeYTswm
9Ny+JkcY+aq3XRVtDlRn/ImGaEN2KuZFfBUm62TSHu+GGJT+nxCEelfS7jiN
qFQQmFT/qp+o1Sx/A7/JualACwxjJBfPwFtpifOGHSNpp+CncEZL+BkEKwfx
FkUqhNv5BqtUyWCubfYKeyrwdrvIsjG132w4pVRb89tqSdTvsjILMqJ0cbKx
Vczv8Ix2jJOVNpBpEXR15aMtV2Wop/RNHa/poiWqP0iMqMycCzJkeORTJYAm
vmYNX6DQ/vnLIVZNAvh5LrBwITxPXyBsPCi7vB3YcOd3vQOGZqPeBtNHafjv
2O2swAlPDvu1ap0J9rD1FkN3f6ciSORUgv6sAGH7kG2XcTawq2ho9/FGPmgp
YVgL1EYnrURIESf/6CtIcz20/bPbRe/Jw0gnh0vFru0psgzxnKAVMCyz8I2Z
+CR2fD8aM8nZpn84CRUwFsucIhFOfdyJAvMQksizzN8uyr5NkDyas7NbcHyl
VOEN13XryUyA98gUiS6mUuB3y1GFmQLr4KM4iRW08MezhT5TILQ7bacveKiD
0R/NZ4NvPHj/HVxKq2ga/RyMS0ZoBL9CRfHV9lc2nFf1Y1H9IU+SqlHffO/Q
O6ruC8M84fCu+myw6KGaGYD0WLCzX/NBqJaGIjuAdafiWgg0vY3MO4HOsq6n
t4E9827DHYemuGLGHP0TpoqkfGFs3KNiK8w31WdEAMBDKiGq3KYVZgDTw+wp
8WC7b49imWtlhmuGZkSmwRyWX0YNZ7RDMYOFgrFuefctXPwJmXraVMoCbL6U
p3nQ6su/6ajiGO+gHoFA0i1ES59pF9XpsmbpNMU1BtSgB3gtrodFDYb5c8GV
pp6iMJcfzYtGh3ZvXcMA30vTqUfngRpWIwdZ7Kl86xoDc9pHh1ZkKyUonjWe
VBpXl13lX9w1Q0fQ7jjj7JbbQi1arhoWezJj0Wa2hEcvlN9bSJdJcgXf9Gkx
3mFJHudeplCm8v4niwgox+2/rCRPmox3MYA5ORq4j9HdnkXSL9PZB6kDsnyR
IZsTKpPSkmIa1rviPOUzrLYz+dOO7HLaxWGVANeEpKmMv9uye6aMl+LMmUiG
Ukk1SbYH7tjIlCkFavDUOHZFGyRzDD4MAFy+2ihlOFqKaT/ns2ZFqFCWmPqM
YKHXFetNJZfIczaBvKNW8CrOos7bEA2jMdpc01OISieeUHvWPUi6PqBfWoMr
E8wDAool/Uol30o7F/BMHoNq+JrxPPMDv0mI2EdoSH/MEnkQe3pCwe44XtVB
WhSqAT5j85tHd0bQtgHgSUIKQT7CWdBIyPzfmy5OfVD+ieat1p/hjL6hREup
Tws6U0J2qglOvQM+cYqFSO3cYH1Uzp6vavWRVda7MTkUTHuwRgMKvGekJvIF
FS6PaWLA4PxYCjqr4LRtCCOufHF86GtsLDCL08SrgIBoP37yBQicrBN8Vg2T
mnEqYlmIAz5Hs5tgJlO/Cn6EZLoV8R7YJfc1MUQSULFDuVU0QlmhqVAvyxWq
bmAZLiXurfzdX//yREkgIppR8UVSM4HVkZ1Djd6Zdd3NBuIvuIcKNHx6AXAD
MrhkpxbFjgvN1Zy/EGsoBnoEAQtTecvB7c3/PvDSVN1r7dWgr/rZTP8KRAuh
RD6Pe9yxV6l+dNHy/3hKv/H0wSmRQa11pgIVbwA8qpptu47gZApBsHFG/+ya
bkh7Hy9LiHT1poZxTyU06/E4ZljOMhe+U20/lsaQ+S9jh6MO/pEucVM/SPFs
MLsBmAMwuyC/MGkscB4+MpuRYkrRrin8wyHd8KA57wO04mdfvNqHO3LcJXQB
E+xxGGm+xTFkAdUO+i1nPTunZjHpGh2c7rRJEooMcntcmJWH8myISbvhzOXd
MgJyLyJ+sTfeB/r8d1vkDfMqPxxkkKF4XJY2uk+ddN+n/8G/+/V+hcSg+kGq
0ILYAtLsfTkNPW2RLym6r8E6Bzew4xtFKyDFoC5vb+X9OiWJkJqLPkuNJrwa
be1GkvKwPCpMY6jYUetN1AhWPq52opZClNjxXHgLD0bKKQxvxPR7H5icB+25
dFj+rfnDywDsH5mI8THxHPkJnD9W8UXJT7MkXXNSEGd7uTx9ENXHsqhSKII1
w9hIn/vj6pwCx6k6flI/qVNDapeFezlgXI4lnrSb8UrrthOUKzG1on4pRyLz
bGlHNBGX7CujNK8VzrJSfejgNn5o/Yyjt4NmF/BI+gY/IHL6Q0ZZ8si/1XCV
0X5sd+i8LhWQSpeXEs4abkDslwKlv8t2kyowKRQOpvguqFG5QU9dgVao7PRW
1h+JGDgUtWple/XqUTmezsfx1nQR+2W+7CtejhIIa5gD6y/VhxqO4x69Ufnz
Z7zFLoayGw4Ir/eYezuaoeJJOQGcU+mPiEQPRG1u6yi2/qcjQNuN4ZdZ9yqt
zdJnz8ltppV4bsBm9HXO9YeOf+HEsOQDoEyf12hPg36l/WSfj5UbcOK5ZYnW
9YIc6CzBmKpkMqKf/0qngdOQDRfLYz0MQAqtFw1kKYnCCDEW7cX6WTC1e+8w
BXbMPRpWIlB8pqhC4oWLRLGEIFaVQkiswj41NZ9FnpDj9R460srS0PulcBen
HPflD/ht7pTRO9vMIRuxX9V2KWlsbZQ9ZQm8O//Ph03KKV/hUYrHQLvZg9o4
FnvrsOTw1rbbF+Q0MWgxjJ7u5ZxkeMH757oRBywdv4633g4wyRdL75vUWjM2
6+CnNzAToUyOclENnUwdMhdBfgX3DRx6hOCVyhW41YtOFeXYhDfUD1X7RFiJ
ivmI3JrcxHF2wtuYUml5kxKAlJ0MtBijsdySfWMJj+pCxyKAKyokANXgiXZ9
dhOIcWnq4SpGg+YTfHnaRex22uJypCzT0OXmt7K6yUFTgfd8LGf67jaE8gM4
f+oikwjxuCg3c8wbfvO4GrvhKJ2OGgBLFbdEaVt9EjepZh12f576WM26nb4o
52hj1MnQVXIKxNMJYH+hUWEGxxsuarvjAHkpnFO/+sFRkWht0A/wGh7Xd82a
V5yx6PpTfGa8QZ8SFS/jIljLkOo5Qm9HBPyduyFdVp2K6vurMzmbd3CSUHGo
vp9mTZQudFu8RswKBpZyFOtUEP2F0EsbiNxj2hp3RlmC2ZoxNEd7gDE0WaR4
KEzWr+/WJQz1ohxiuPWVAQP77HcrFGtO9QD/wjthB1yk0/vvsQcqYg0ii73f
nKE5UtrcXa63Hczs9AY5eiiA5BjSDtHxDy1Rx4jbOI6s1HKSa2O+JAETpGNn
ugmIyGd8xis4IqCHli9M7gA2AH5GOPnC73xhByw4bpy9Psc672xg6gv3kvLJ
E/lxLgu0tqgehXaM/54IIG0J3kYTrQalnsBzMTwezIUibqEZKJNLaG9Cy3/4
BMKb1vzYhRfUFhits3F3Ps4LSYO4iAB5nTzJNssVhdcZhHNbGUFn0FoR21uE
nnVQEURnVlcGpZNGWujjcic03q8GQCDmqxIXim2TRV7ywR+5jmAFvVOKNy3+
tgyDRGqQYQDmPCp3Ed++dgaMVy4i/pnp77Sr2iiMpAVN09MiIHbSfM/1Fd+Q
wi4Ynq0MOig6+gvobxU4dbbeMDWUnbGWue6eXD5UccYLG0MjSH63/eo+Tcw2
bF328TYSHC6cYUUgETRF1hCUT325T1QYHmnyDYtIg9Q7n5TbP/y8HopOTn9h
BYhBrDCyc/35D7xNZsO0MZDvyQ8KrhpH840g4/KMAzmqJHeKKAGvgGmeSw3m
xgXvEQamwsL9hLaQBVJclZc6weXgZZ/aQlP2H02ZFuy+PwK0w3Oktf4W3Z39
i0P7NJ8aK7HEYMlO6q9D61lUCiaaVJNoYvidMqrOHu/MlbDBmevkS8KaU1D5
1zmmANO6pbL+jlncMOyfR+kh190SpvW0ihSdmbhizee/GRYweW1wS9lhrPuy
p4K6GY65YeIKcBJsXb4E7DV9HN4X/ZuEA8CZCCSVHwgl9J6WWT8ltOnWcaXK
uQE8vFEMZNXLvn/1Vq4GGU2rr7Nkbfbn5vNvtYnJ56dARLI4kXd4M7Z8HVdU
5QdWkJmglu+96ud9DXkO5DbKM9/VHEn8iaAck18/XnJEGNI6WSkSstKrNhOf
Se7/XxnSTj8KQkK6GVwBUKlpeHpFdKg7U0Mf/mAtUh7/cHsGm4OJqOwmcgwB
H2lO+f1u1t6smwRBepzGO8xch/DT8W/DFIr1ySQpMtLLh0OHlfDIV5DDAFwA
0wSdVBriDeXO3aB8gXlihUac0C460jFVqBGXzOqsmZ8QhhHoLgNaYisdumuw
hPCztzVz8cf6AqRbkJYQx/oohLZAa9RJnTXwOc7SmGn/56lfQMpXpWKpSDFg
uwN/vAZqb4cQqmNRSPmpUOSAjiNIEr9fwEopbMjMQlQe+CdA93RHoc5Ua5qU
HyWzZNEOoYzc4X9agpZhO7VJxYuUgCpzi+w7Ak3rLPOfFd6H2UWDhMKuLKwy
NbT6lp8wEbuzH0lIn+2e8MuXCoMxo4BT2V+u5KB9CunMNe1ea0M7SYnVXKR9
eanFgwB6+RGxfv5PJCW6q3X7go+4ozYS9u1mwC3+mhJi2Yq1N3y8y+H66mcQ
OU3DdRc8RWlberea7aMZinLqwUUO19F+jreUGy/m7anbVh0On4CopVwHIIqS
koGtbHw4m9MRpwbBByA+NqotrGyEgJ/AWwKJLCdkb49tjFRB15H8Xhvj8NID
6A5u5kW9X7Itz/LV4RCDJIy+tA7VCKgsuM3SNEYx+Bekl53J9yHA1kICA7CW
m6OPD8oKYiQJIg2pnXy8MJFf5L1ZMkvf3vVCIfGbO4NHGFMrXceIToig6eWe
MNkhGa0kFMuSE2SccNcV7MsP5XWM395Tr6EXkOFCd/C3pKjHWLKNLfMmuTpF
tix8YCcknEYLd22QvUrF9NxMm+ernzb7sSHod+iOpowzkAVvO2z9vTcDfGZu
t004PThR6uKa6axGMFXhLq85PRDdfRSn9TBplmXSJMfq3N1h/FhIQclCvqYW
w9oVM6VH9OWmb3P3X+7pBE+PbIF/t/V2rzewXmziUS8f0PkENnNOkf0j+/p/
xWKyPcOcI/Pwet28Ht9u1Ol3aDPBI6gtIPwEGaCNcSCwfiCK9fcs085SoOEk
gUVE0Z/PUnzpUTHdcFBbigmXhP7/TSw/hoK+T5JxM1gUpqLCrPQSPMyAD4qd
B0RmqP4XoddFMVUCUy8BlJDfQhxQsV91365T4dZWZWoirMn4lP0xv44P3iqB
ZXna7lrD1RnZCf1RL08yHOAW4n32+KdRIRCLmwXh20nLHTx1DkxF89Cg3t6G
yix2/LWhnI8pJkI51xMwHVqsFfYXdlgxmxnUSebzGYeov/5OgY5yVhmYiHyD
C7mHesuacwVnjXJU15lbVufDUB2UxMFl+S2bmfYNZI958O742qT5eAKBomAz
1U4BxrafrVdWFqc0wSFfnTxfK5GUdk7Q7pA0f5kX9rJKENmyv40n8dv96a21
utvFRAyT2ZcV9X8JbAPtLlIEqK5dfWAXMkpRN+0ufqqbRaaU/Tay95Ip2lbN
e0W08HZq9x/03SCV133ke2/4y6B4VWBxHnepKWzkRr7k6s4XwaHwtWp6g/mW
zZOoysY0YkLGRDHrRXt3ojVF2P8D5UAkIf6VbH7wds7COUE670eAVPdQI18u
ncdsSuMMQRuSn6VYx9EuiXtfqc4/i8fUy0y4MtmskR6o6LEU+YP52Hsqo7im
caLXfiAwVba3LN8/FN11xgHGsaQgAwTPPWIM+mYP0wStrrcAugGXnjstt/3g
qIarP+aSVbzzDwG5Bk8TOiLcnPR8+9cRW6qfTw6naVh+gNfg6q817MHxsUUi
5ASPIseWC1vlFTAfNiakoXYc/WCKIz/Gxd/lWRQYEgMEV7tyCGzgn8Bgk046
RpifIluc5TUYe1SYFrcmRFEy+A3ORsqadQH0sNouOdWzrr5aYx3M77kHaJxW
aUUPlz9v1GmbnnTfSykchjrtbiFfVH2eJwOJ3hg/2TT8tYFEKdg625v5ya61
HLDYU50nTOhnwZ9yEzdPZI02HiZU3OGuT1zbCd6uQ+x2229l5prRomsEwus1
ezEJ/LaMJ21n0eRCDoCLuZhQ/5Tl0g2JwKFSqF4DUyTWQ94lbUMqkArQr0Kf
bkcOpvnWGHIfPvtR9TE1E4o+3j6exvlUUVTA6RzCIZkPieR77pQumrXFgJXb
Wv4Yh9nvdRXTZtfqNiAVCwQLOZlo5LHK90Ytao7iBo0H8LHaMGH+CCAilIH1
LPo8bFP8fBGt3+emCFZlpkLSW7jR+mvRlCYEm248krx5NWyqphWzXkQ/0pGf
/lB+Kgk8ho8sssktnConX5k9B0Sw7D8IdN1jSAUiwsLOtTcH9MW7mxcELRaB
fzEecD5/dpBebC6iAib8vixEt1uRV2MWpfXOWKE7bmCVPbng+4Wd0GJB/Z+c
IauhUEqHXtYvMaGUH5ONbTKO7/dfxDldN4d/IdxqV9U6z9qLdgc0vlI8Kkel
+W711KTXpbOKWfLDuzB3n0+GjyBMbMfOCodVMmUi3U4omc8BxiCJZbnlJC3h
FrpzAsAuAgnNioX3EZsQUBi7inscwph1QtKfmA8cqqpcn9j9kicvhZDYdTVn
0Sea6+KyZswTVMbwz/1iEvLiFQncL7VRyVaTdQWLdQuw9e8F3PBQY/Lt+xCC
hiXjF48rxbc1adIzFG6MOTyalssfdtGrxW30ymUTcKXPCgPyvPhuIym3QtaE
UdIBDxEodpUsuS+qz0idAZGbh0Pzy23jWFe1g989Few5pIDAPn1SHI09BZ5X
j0kyCS3T23CDZErihxTLjuhgILxO97P/c13lozwWjeLAen8erL1dJRHp5p0Z
0PqVmtQsns6kZpdD0u1pEKA638nLRpEoTJOAlcJCvCvl7PSsPnT9XEouP8v8
j7kdPuJYJEtg5dWMxUTX+razIb9ouBfta6K3cyOzaUZRwZttHqpeS5W6R6cJ
CIQJ9NtGgg6ebrH7xfMHwOzgwduhvnxQpugKFoa0462QB0RP23siAyPwrRoS
IFgLCZbx2op3i13X2gtr2xkKvYCSrFfsCYyHJXgXaoDyhNhvfgCPgULqY9Em
YtLpyCUloJ4XRV7gWsNynhsorXAa3c5H5AHpThBfhVrCpT2y0T/XbK03Fs3j
lDW4uR4DGldEIFajbnOYbyaCLmXm4ibyZcn/zLsril8x1ADT/msXUim2hbDn
EfBxD3ZXtf8SUZA1w0HiNpg0QaVaQoGWd8IzqdmPx97Gxn96XagDrlYOX/Ap
oiJNLavHSbspMhMpTsL6ElX74WP8hLJ/VwY8mFRiQ08oXaNRYFOh8zmOMjs/
I2KbsLzbliJQPm35+P6U9QTGbhfEPYAu+Y2wuWwNjhTIqVTHrZSEu5wH66sE
zd7/KBrkhs8p0Gpd4rgAUT1IemWihzpBpGnScvGa3wv/nTn+28QYGNaEXT60
ssWUWObED9wYjIYOlYCq+UEvnZ8p3UgDRhV0X/saaSnbvMFILqm8AQm0L08e
idwvlZRS2KL8rpM8qI/D5PwVpxy2lcUwSWplPUhro79s7KTJYI35U8kDsKOG
88CFB+Uq/28EmPwmiEwUSZd4Li23NK+jCHL0Dg05+oaxN6rs8ASNovfzhW9c
fRk0rXjYVgv5wub8sxRPDbXBXwD2t2IJdE4pfVtpetJ94EcGXncAwdDvNEy+
RErSZ91D0thaSZf0S5hlwlNnII8R8AU6zX4Gqq4/sOGIWh/xMZ2V2kNxsf+1
C39L3/FmtBSgE+2hkfipNc/dkWvXPIhnIf9Deot42ptdD50TlDug6AzGLvSt
0dzCwPX2gle+fj09L5kQWGcE4693EOKOTmA4+VnbWqZGENKd1y0q17AhBsNp
+J2qjZLbhli+ixzQo1rhOQ+errT2t3/Z8mUCVYMBJx2XWb4U/jF8t5vZAFzx
gYUz3gYvInASwcbn7chixm5oJxKPofCz2LINQwd+/45Ep/rU6XAEl0dboBse
sPMWnjYLosgI4Jax2wrl11f97vPr84T1CI4CBfrEEdLY+2mS9RHk3VgNy+8H
K85lrrG6kpU/RID6Or2TRwZX1iINkFvDvq9cpBrj1lu1r2xyA9qRsUS+JgvM
iMAqV1B5iIKS3My9CGHQV568teGvMnYFfB4N01r07XodpF/NcqkD7jfPu9nV
4tqtdGG9bRBLctoy/7UUV8V1FmM4ZURsrvAHL2LwwZchQQ7LBTkq2RddFgR3
19hwjrwRHLk/w7ZuUkMXIuetb+mbKH8hLshHEofznRQPQq3sD0Wt+LHfTiRQ
HKhKF03zWac7Tsyn57Ar3uTut6J3g8ymR2N5cfTJWRtjHbg364SvIDPhxeWC
+F9HbldQvmZ2bXdjVEVQ/o4ccCVxfbzxc/khpJ8wvjPhVDS6b4eqkk/2xUFo
PVabkDFzLZPGBywA11JQDtCOhbuItyMkTMUHpVrqbmnf+9xk8+gCztIeFsXM
Cf7mm0JdC1vvvC3ODxEaQDrAZ/1fXiTVafdWjnMnZUnlCF2fwFLOP9gWb4Li
NMbkpSMwCMLwB4XtzcXL9Si5wNCqCqjjqQugtVKoskFZeNVpmAzvyL7YrQx4
Xy2JpuDL9ErGKrcU/OWc62LU1NrtYjT5VqXgIODyIpXI6Hs3MDfqXW94Xopy
bw0NB0hMwwuahTxzHUpWL/Lg4ZQqcCCYSHtlpG7loUvEvn5vykzgByrqxxRU
KbIetCccL/vh49bY4D1NLmOZIWwKyrpRI8Rw/UzpcKFDbwhbsKDiHeyiE32B
vSXBqFNfxcD32pEgwLtVFwbL6+OsH6PIciGm2a5BxMNfzqh0jAaGVSxYpPy0
DKrpvbuUNH8MVwvypMmyh1CjKl9OIVc/TmP7K5b+rkpW5kiEApl8FiKCd4Zl
pbmyBM5ZwSeBL2TZELn3tBrZUFe047uKzWas8/9QdvLyQ/TL+TLODgrjP9GP
zVm+tI+2ghKbYnxDWtSNRpc4iFNi3lTqa4J3I4zhhZFIJ/n/rKUAeFiYhlPI
j/b5S10b4SlgeBkzUfUbkSc7BjialZ7ALFsW8a3IImTSN9x4DdgMhnQ3f1iy
wZyq3SiwpZybAQFc9SnNKc6szSEvyx47dDikjfvvlTVrBv2JgHHVPrCLhs9q
wghw96+rim3m6T0m6keuDVShmdekNcxETzDC7Enln/5IlZYwWQFwYBc0LJsk
nEyFjPo01zHTzdbtFVCnhOtjxNgON6f1T2cPgSk4E1Wi5zwvRwLP8O6NSPyl
dLfbHpniI/ogaNeGPaIwLRFkig0h0stOyT4usBXBGPZ62qOy20JL+8NbAA9E
hsJuHrenuvrSDnp+hs0a2m6hKua+JC4GdcA2cJp9aSSxhQOkPdqMFuolFdHQ
rDCLYmiZQUGRlz1vpAy4qiG098TT0vCBpY/fIX47U6NNPpQFTDQqk8Z3N/dQ
EqAE3Q/WGjGUgu9eg4BufV0WUhxqg6iV2IRuMp/3iH/xIGripZh7ZR3u5uQk
lcnDGXk4N8aqaIAzxl8swpWW5q3RYobodBv5RL+fNp5Xi27gNnEuquxKHYiM
mTpEzk3yLbSYHZtZ/QJgCAmV674lL6HtpODrGjiN0KFgoO173JSojEUT60AS
sbAsX9IVnx7QxvchKJ/yx8Yj9yo4YtU9kkbDHkR2SzAR8B/afhc3H14HIOlF
kF/ylJiJrKQNOlkfuiURNZyK+iBysCxvb7PbRlahp49t9qdJgLhUMmFOxBtb
7qv/3ixznei1g/rWeuQEFTMpX+acZAKTPajbGj4RF3h1ae+KO9SxxhREAN4B
cGlKR1ZC7kJBKRq8SP++El4oKnoFtPE2Qv4cPVa5fd03n1Y/DX3tZxqMTYqu
ZlLdlhs/N3xt4WBdPFRDu1oIdLr0waTr3+VDrHgmG3FrdyGxJ9sKBD25QFxp
oKfAnRff3uKs35Tgyz48wYOM+xhnvBKwp0EOQ5fFKfjancOvrg5TC9IO3cuz
iUl6MYQgly0QtcdCehQnfYEwhzY01AmqW+EjOTdHMBknL/sa2yM7p2YZ7O8S
Lp61R8Gni6d2wYMcy2wcfH7TnL1e7lWf+jUeiEd8PaGEGr3MF9Fl0Rrr9AUR
ifXthYUebWFFSeLGMU0MaRVGu+/Cc5TOQ2fk0KRRiTb9xgCuiXHkqQ/rObyU
SdizT4wEewFAhPdlv93miWkroF/3nswYPolmUPwaCwlV+B45+3j+ijlCrwZs
OJkzOU77MJe41XW7UCRXvYo194VquQjlQT9D82njfltfa4YXONpSD6CcAKRb
pbxEsCl5gnOK0ioZtPcB6E20Xya7w04v5VGo3WZC5SqPMwf9Q5o7pNbtYfNn
Y2hxd9P/xl084JyaItNGU+pDjkd85U3pasJjNLgjMVQghUI9QdbRRYtEQkxD
a0qyFKtB2Ik2Ve3B6Mw0YN5V5AoYD+/ctfECXsgDGUKyd8uw+vEolAFdBo5V
e/1b1BHT6S9Q79qnFjymBFCYganuXA0ZO8R62iZg4xgUAsNkqFuwaKNK6JUI
82XlDX6sXRplHsaFbH6U9nUaUtHep8F3nnNgKtZli/26nFdq8fdTIkS+Bsak
lInJYHYrBv41Kt4nP6CyRkhOQc3tmS6cvIjJVC2QjH8ofkCoH1GbxwP4sK33
KwpzoiN8MXBdOq/0TReXg09xeEvUnOLLne5KqaL13ytmkxdcQh75rYP2XIXG
agyRWNcfNKEkFEdUixnOtm8u/q+6xBOVji8LqkX9TInalNld48hJBX+eXHzT
VKXW+JkvN6qjYquqIhfXqAgFn/mZ46Rl2CENRXQCZ3aUpEeucyOssz6/cNzo
gwUj96i5Lqsx52twfoRINlbdfYmtv0vmSvBfOAemhGxe2FeyIdtNaF2/Hce2
Fa2V/DbOJlwHuuzKrY8g8rGeKjXwYn36TE3HckKyQ9XeCPO3/X1WIQM0RPpT
cRb49a52E7jHrA/wbojdCgEo0rB9Ud8V/8/miq8GVFZfcf5VCM122agiWdHC
7rxaUvtLbTA0uIp9YMYGOYT1JnAXZ28kg2Xb3BxvuHPpSEIikw0JFj3DFX8P
49jQFXHd3WzUux7rPMZwiceaae+5opAEdzUdGfYbOKhC7rzm++hcifRu00Ho
lI6VfyhiZnvecA0QS3tK1tBdvHv/4itd9EWt+Mjxd1s/oNx0b6DWTSW51d6i
et2lrLJQ/9f1B6AwOxW9bpIjAzTPsgxZYkvpEa5P2ZLXoUfdQyLArifyExLk
0Q1/kNDYCHh8jlbBNurNIGnzEl3hSX4gWE3jM6cYJ3h3Ixr5noIj+Eu4dwe2
uqhsbyi3e3R6sDOIsB/6itfm+ZcLdEjkGs2rAbGhd6Dd0NQHRd2ojv62NZAC
z2tzMWUrqb0S9c1ncs5ME9GoXK3fKoLXcOk0ufNZRYR9PR9AIYAtUuM6coHg
H9ugNwyhBpQVJlbioMvb5bep+mJP1oVyFhqkZ1fY6znyKjdgm2p9P9SgAYS3
z6hguR2Vl9zuymDzUgtvePkLekyosfrH5FvW2/2asoBU4NEJt04+8yKdRnjs
0kNks72Hgel/vfvaNLBEshGY6q9FlRWP/WfS12HxjnURdIg0wgwQWuBMhgm8
zWCkG19g0El7QI4hvqXhJVa6UjQBwDKFK/eDEB/lvwvWTqXwgNXu9t/iniD6
wh54kgVADDpPsOcNxTKmBiorPowGZRr3SACiEvcJcZhDEt11HmcZkKh7FFCh
uVRHtGkjFGm6j6LWIf14IAmeyc+/Zq3mQQKddR3UkU/UrPLpf0pmA5AZpA0S
PgFXyIrWRsGm3+k7ljDyIxg+zhjHQFsYh/bDvf1EQaO144RNyUSVWkbMhOiH
qdkSbJDEkfvPFRZeOXyKDZGXDGPZkFVhvD3hHfKeFJtEyTPO6yokxRRrt6dV
emeGtQGeXrDI6g1jrqWsO4XeNSE2s7eOvuGmNV8Hjege7eXp+YcI9vmlg3Xz
0fSdIASzf0fveKIun1hiNI1B6qTSPiHn4GFRvCZox6MzklMQH5KpfEqDPXUK
sXDe8x+IzRmMETv1jsZHgxkP4LvONv0kr439xM9DE/sSD2LVyFcTFAbm1Q48
HaGAic8sTkEQWZmHJdkMLI8r2kf/bECa88PNL7EdTOIFYS9b342r7tL822oI
jBlPc+s87D7tEQ3UHeJZXc97kbjsjNYaA+2UsSizc7wfFgD6+nEAy50OI1nV
hAdjaAfqOC0h8DqmEmZAjtITFy275qd/wHyz7svJOAeW5kTAQw8BGPQ7gPPr
DB9N0B9F8280wRw+Us2Y+syr5rno/6KvSHBz+WmzDSTgC6mRWC8rDnjysmG2
Q4Szf7j8WE33fG6uGLwj4QWIJWwaB2raxl02PbGQeZM/GfeX0OBCZTqSTubm
+HusYJ7LRuR1g2hFKZGf8G9buGgIY7CXSDrJwcMl3px2pJnAf8U8T3kxoE+Z
XQO1HOXEqtb138xQl904N95gK3p8GB3jbQwWLBc9CixK6+NwoKXQcPjfZN5b
cGvErdS1U6vrDhAJs7WnDPVOeOrjojnypstcxgd1/jtdqTit7+he5x0PsBG1
U8UNAjCFMXJjwWz13riAm7/rkE9THGcxrMTo4pYuRC4QBB5DUSyycTIj5Frx
wEQPj+bTFc3WPFT/jQ7G/1E9v/LcBN1hDtLkbXkUyXXZ9UrmVhK9axcoaX/8
i2i7jdFXGFAINu+PUI4dLU9fi7UP4OdFSdePAMntvxL+xNCTVZlEao02NHdw
eSdXluhhxsBzSPakD86pZPLgDpiwn7vni/PPcvJA9tDNPJJqe0KXeTXOI45V
O6EbB1hfZRridy81Rj5GLXjZ9YzkEwQyEa70L1pCfjc83nk5PyY22NBwMn6h
ogc1XhiBtIJtCdwYW08EYc0WRLK1SwlzwIPZSier3/VAP+iJsZJUwyR5OeMX
409WaULqBzDrlqrvCxLvxqFN5qjEF8Ta5iTVc/fmJJP18KzgYiDwrB3r+Jbh
yCTQyCvezFSwH19unReGOhLr65hzov+nC/YyiOlcZ4oU2J2v7/0++UptSN/9
Es+sXtj62/0ZAYQZGnHf58JN16FTVd3FIZ15zI+RaQ+dqhej+q67WZ1D4DoR
ximuWIDwJD1/rH4WMFBnATCW8jKT+N3DrJAfmzMyPrNLG2wHyMTM4ne8eqvt
wCiFpziY/WTIgz8eVIWLUc1qcXKyNWic5x97p6U53dITsLsb0TsaUJRn/JmB
X5hsVbr87E0ivwsawSMEJJnKhLPxi9njlgcJ33XknYGcZcKwUDyYWP9A2Fmc
G0e3MxvAXzZV4i+c1o5H7J6/Kyj8VrwRIjNay7tCuZxrHX4LuSTUfbLTBQYr
ULCzxnuBSaMmX4hyP1NsWdAtMJFDCltroVO0XIyz6a80pRj9n7s07P15Wdzf
nxD6PpR2GvKD195Sq77ilAS+ucSOZ7ZCK2gKi9znEDh/yeoPmJWWzxR9h0g+
N9WhtI5u1M9UR0Yh7G66vnXhVVS8hMf/DQBtXg8XdNKauMUnSohrYkqP9NNT
dXhPPYDj7Jgxl+x8w6WBLiBDFtptUKdK5cQJdoi7zZquKpPsQaj1iH9DhNqQ
KEMyU1IRBLnQ/FORB4tiOvwFXRcesydfidd0ieEneJ/xjBD9AG+i4adfWsu/
doncZ2EJNnGyo31XI9oLOBtBcZe5mIHwaek+FXEeYGKEE62X9qJ0JJ4oItH7
no2BkIJQViU8nuA3/WGss+K++h2XTWDm7YuiDd1+3GIN7lSKFBPpncQf8hry
0uoRc0PeLUC5s/RXNot6/57uOZuawrDrNp69pz77YpyAuhypVjsBuP0xU+pP
nnANJ0pgzlOhiUqmLI7xWgkWmaiovK6JFAxZa3bAcvCE90PyAX0qgOCJm0Ew
e3UdTeQDTbDEoseF0fbluw6Umqc2jggZ5OzVFc6rByQuEJ5CWC2KmlPbuUfx
EqIMF5Wt4qus1t/12mm4CdMo6KalHltBOMsAfRmtlfT3oebrZyKu39GTj2ZU
mqWVUUlq+FldBnuwdgB8ewXXG+Jsc6w6LlIOszC81eoY6Dq5o/zQE3kmMj0W
1f8KQe/u7AhV6ze0VbZfJICDcEp/FMMFT8Tc/YxxybcKg9RbdxR01Z4lCpsb
oXUPrGTHLffxFTRKuVlrOqJS6Bvn/JUvi/3goSfKqtnFLCsXIuC8tudvEH/M
x8WOIm8eO7E75ScNrbuQVKj+fKvNeGTaj3ui+yBk0c/gFxqJKe/7db+6Vq1C
FZ1ZlUzJbC3NTGquiwBV7BUNKpt16G706e+Nb7QGNxoSjl9GUkjcpz1481fb
EkHTZTM6Mh3C+AcOX7BFTYpM9PbhSKkl0m1nuzaw18pj8LShNn2WqB9UpXEF
CgJ40QJbu4/McP9X7Nm0xw1oZhla4/NvEPqlUdQS2AYyogoz4qNHsoB3OnjY
qmDZ7y+GiQuZHhuv8RU2d/Iq9l4Trrb83kEYueYI3w5G1AWWNoq6FXte5kCi
FJvhpw/Hb32NuXJoKdXz60EljbIpGn+0XYD6QUzVop8hKerj+FJ3eFuIpnpL
KqNH0qh/9f4ruQTDZlUVr9PVrtrFW75UJ9knjHg0Fqu2JaZwXGMzbY+1TGUK
wb3UIt7CgmnGD3De6IvCwJ/fa2ilIiwXCxnPzCQukrVnKdkxz64jh49pdo1N
KZ8tTmy1NChba92cn2H9qXuYTccJEhJ3kHkjuV9KTVWMpz1AjAT98LFgnAFG
LU3W3aCefY9qhu8M8QYLPJtY1lcDlDE2Zv9AtwS4DIXIwhdYRg225/U4vyWy
wIvsagj+49QPAs/c5iKn7lWmd1TAeri9MY+Yxx5gFDFpJigEtzGOuHWipvjB
MKrWLXNbGQHmf5d7BFGAfSQsdVQ36xC1dMtYo1qFe4mi4PS/2X63VQqfYX/f
flRDPM7sAHPHYg9fNDK1bdo6GDKlvbDMMgv+YIDqgTjsA+aKWPSw+4hDkO7+
xSXiR4deB/i72aL3wAULt561vRmcsCvN48J30ggRrzRJUUkYx88s2FvjmdJu
tLAFNGdi0b9erjW0iImt2bxP9G5dnway2/TWMUASzmfd9ZYlo0j9IwS+oD1/
CNQiR9ih6LzAAKHmUVWCMG8hfKiyLsE823ca8coUouUzuUpFvTsvEjQmnIoY
FGbyvgA8srhm/cSkKqfVVsbONVMo8ygy3Kx0EPUCxVGfu9pXlLQm9DtTfnDT
RDI6tlwLTG/bsZDJYjWPaC7FP3YnZnr5jWub90/cs0qa8kDpbLNwatHTS7Bs
ZDukAdFUpZhXNeDD5g+Zu9yC3rDBEkX9RKigSzWVPLMScrD5qJXW8TK50KOs
XooE0Oxx7UPxkAEezy+GvYu24UHB2Zd9hA7V8Wfp+3gRTt3DGuxRHc56rE2y
m+WRUEO1l0dn4vUKJsr4cZyZRzlp9p9iOq/ym+nTzGgh13VqCeC4MvyKdFeT
5D4K+JEc0rhF4zIV1reAV17LIT2TsI1of391vBR7hIzOZqkzQrJRtjt+tRqE
+Ne04N/eOo/4nL0KcjE4uy/+9cJHG4G8a28807HNsp4O9JNgRsXh71biWxO8
SW662o2SBQxgnjUAldCYXfXLHbL0SKM6snigkMFwROCSQYvV6ld8DQvfIElM
OxRtoNtzAnlXsGAluRc7jk4xw05FNie+mEn8gtUSw/Gg4N4S1g9bOAtX23Cn
76tiXoDZb7VmOUj7rYCiC+P6cjK5xVZch6ldWLWHVxVxjNNClpj/DKwwylni
qU/YBzLye4SLvFxlpiF3hvnhmcYERqAXYZJ7plEdXnlMmI6pxa6H+SuLZMj9
xL3Kz0701ksLSYy2YoA7CYNbL0dLYdl0VJf5cAQ1RaJgjGNgvK/OYcAWj8Ph
euJDC3FqA5VuZcadifW99okHmKpkHAUz4axN0GVQZKEnEABhH+u8WfzyYfT/
oV+2OJeqblZ+YDEtoNOU9Ma+5vXwT3HyBRerpoMJ+NwD3dA2GLKSeCh0OLAB
9F+mgIe0fnsh/XQnLWUwqtjy17o/zXojXXFxChLpam9uP9vOqDdZjOhSft1g
2LPEWJwubzPnI4QjnA0RvfOMR+ve30JoFf57phtHalFUDISj7syakxdLGhi2
5sxKqEe+o4rYq0s5ZLqrc9buq2onHnjoNWfaufP7pr7dace/qTrTxVC9Kd1u
wL1jLHW/NdRlFzNoQZ4FHkHMpff3hi8p87c/rknut25TXHasci9Q0NNivtg2
+7yjP5iyu485KH36t3dscQrM9Bit1IChvWnKQ7LW6pDuCWlQSM8STpXD+EYs
GZzBWGeFLcVD5fDm5lf36uRWsafof7qupfKvyN9l4pfdDq1lhYawOlBILdTj
W9g/ir+rZ3h2viulfKrIxV85hU9WuhuKUxNhnnv04pUz5B0jPw1NpuLEJPfQ
xz8B09XqNu4bRHHzALLP2BtV4b3Xt589E3eBxaYvBd0G8N4LoDYcy8Qen4WZ
9tl6mASbeTUJpftBjo0yKiOXpcY9Fq+tMQFtFchA6owGATNEB8oOK3GDcQfj
ModBQPvgejiCUeXLJ8gieFW0wjwhVOZ5qehr+nUEIylX4Vt8JVhvueiMKVWj
i1Ke3bCNm8qM5aGlpTJcKrSEv9YXpNohg4lfJQGSdcyDuyneAOcJx+nv8cRj
jH9s35LxKfFOAsCeKOQx3SPhKz/BtuhJH63ocbUhoQsRCDrJtmuBDr/6JtIu
2XkUN3vcBqEiCeN8R75EQrAqy6Om/jhP/HjQJwTTFKBDsqGehFopUZg7N/AD
pM0+4yVF8tLV5SrjlMqHfzqZJXZRxEYE9AIlqiJHnYcLgVM/+J89g+zEjnbw
qhqg//12RxPhlPHWS4/QpUSwtOEYktCineSeaTHOPaxktOL2qgUQsYF5W9QK
jZsGra/63dtYKFpSvDSx4U5AOOn94io1+dLM9GVf7oerttDb4dokk2MeGiH1
B0yvhQjXFwzwt58hh+f/UpOUEpQK0uvrRt1HDuc4vI1ga4yBjd/9yflUS82a
necFoGoIJbu2PT/JwthhDrtbIKOh0uhhEVfthS8JobvgP/EwRKvMY5uSykHh
tVX6PiOxAGtq/Cv0LORpmT/8KDeNsSCsxb1kJ3B9jmoch1dOsRDkt6cVkDlx
faAxmVDaIdzJo0xG34lCxr0s9GGdX8Okw9gH4D9Zgo1kpk/2nEqFIb62xusT
Ma11/EnvEbpvTnXIr6RLN3NI6vd8OMjp7lkOP1hGWRUkgUi2foVdCPgbzT1Q
dEC/OJYZS2SCD+Ez9dk1qhCncOAvmyQuahtYm7jlWK7ynb1HkfJShjkPw8ls
jYMJzpRS3XWoj23/HloM9lequ6bJEdktm12Obqud/nAmmnaLG9nBzcm35r5z
A6ru/ebKlwZh0D1KkKgdh+VpZhezNzXyTve52eRUMGxLSLOxXZ3ZEFiUAT2U
SSjPOKZefWBnC/3M8Ko2YFghlr+QvRU6Hcm+Yoi7KRZ1qec9qo9Owu6bxmND
Zb1jkjM0JCLz6DweHcgmExYJPO18frGQudI5JDiRm4HQorXBln/ViSs9IAup
DRs87ZRwJyP+6lhtNRUVLzl0VkCuMN7dxNovEhNufi6/E9jD6KcZn6ogsalR
y/TylU7miDPhzivrJ9ubWMF0+noSoFez6nXTxe+6yL5vZB2+VcEL2XXNODw9
Aws+fd+ORWew1gXhzPG5DhUMRv/JDl1VzIEg5rAzp54QGaLss5gv0weWVPYV
EGxX4XyGG3vKN/2Vyl6/KHfqTXjlQrA4JJioymH89N8AdJjWhP3trSkqQZ3X
AECK+Ci5oqvwUWcyc32K0UF9UO5zwF4IJPj+Hdx2qNvDmE8DDo330aFqvbfg
LXSUC+PdBqrzKSJ342Gt6rrUrq86KJ/n3OJKSQzQW+8DnZr9SYhZokehuPj1
j1O/oxusxKiVyZn1X8KLxmFkKnEghXaRKOvjLVFPkJg3Hp3jp+8TD8fDwYIQ
wziIg94AGmHGQXaSGrtsFnaJAgxjEKB2nHaBFd0lcSgbdImwAd4SnnE97TdH
C813tLnkpfw1lNn5wfPEZa3Faqb2hkafwZpKkU0dxJKCoF3QGNYTvRcwK6bw
hlorHN/ueqZNEBgnfQIZheFflLTYOZ/ow3oZtk18DTE+/2JhVHqWiLrI1tIB
PIrNAsFUSLIdmDln1jmjIjExDmTjZPBMl6atQVaQW4QH/v4W4a3FtEd8vNxe
XiCLbLbAtVkO4d62DyYHWLCzmslLt46VoYwziXDsmo6kgbxDqTOgsKweqOw2
PQyAuk7X2tENMf8Zoc2RddwZA4FVIrvlm7XIIs1TZkk06rbFC09Tc3tj4ED7
ydY5/Hjh1DCJ4FqieXyA/AOVgb7MbiBZQfoR9TLktU1WLnP0dqh78MFjtKAe
RZTVrJbwNeldjBxsUt/Y5aWcBoSvJNrNvtFj1+FTNv3g/R0TurXwIyL2+hPZ
gWNQdMa0COrzwB38OiWB8k/HiT+iV/cSBDVmVqva7nsfkYE8ltKebl48MglP
RuPc6pcC6QPBP+rj4oI4h6/a9L5aeevgCAIjmu75gRHj6/vRoWDAXtTMQosB
kh8LL3+NEpgdJ6rQU+ot0fjz3iAV2HLPyWESyiJoIgVFC/Cm8/wuaDQeGXiX
++yNZCXE+ulaxSBN+1Wtnx7P/AmzNhxIy1ji0I2nHBt3nGJZX/3oipC87WXg
iULSR7tCNaCE/CHBV+91ktGhGILYVOltk7EZhRkLM+OyJbaQHzDtdt8OeswX
zdQ0e4i7YDtRQ6OZNC1eMMnZL/K+ZWP2vuuHAHBRonCkrIqCmqlz8R3mvlQv
1cDSxzeaMdGP6sUyUYYxzCLKCdX3UfrA/AfRYfK7MUR1ri1p2EauP2OoIEqU
ysZ/bNLz7Rpoc7ryh3jY2FY+obEDxUn0uYy1iHRKDCjjwBD9BfSxWuoWUYjt
zboHMI8OeESOFpprRseI+M0YGfXxvntdwdK9KAPIXdIj7MGiEWBYerNILdFy
5z02oHmcVBEgam4KA50ldLM58lEPgGPjni8eMRsilkfpoRjreYFkk5CKWwJ8
kUbBj8xfu21EqySKt+CrdVhdG5iA9M0zW4PFf7EB0DZOItVsp2CgG7rXs8wB
HZH005FAYenANJFZvH36EGaG18gVKz5K3bdVsatIPRUPuNLw7Q0wT0Bj6U7X
Bpaav/sA9TM2S3XqaLzQI6P+vBSsroCrjJxPNK28vmmlatyV5FLreY6ptxVH
/UjsJ7nw4F3ao+r5ltResaHm4gqSG/qZ+tOmhhInNQob+ziPUz/xZgMaWWQ7
ZamEhh3mE6tBK5/hurCpyHPjQq8D3vjVlFFMz+RshslYaAHuiyPLhrrySrX/
hs0Dw0eOWg1q7PFF7JOGRHwSbwL7ErmKhShH1VLXl73sDTCsM9i5szzksbb+
ilUAl5oGOZppEfAv9Btd6W2mKXQR4OUBGyCUoCRaN6EOf3WPDavXGrYM81/e
Qr2VrLLC9Zp1P8f0IMrjDm6iAOPif3CvhO4HMZClgq4FlRhIIquyaZVQZw+X
IX5ddr0qwlnVXdIoBVA0YmnrlcKdw0uaGOxMip6tkbwNpIc0k1M4iIJu9k9u
8107NqsX/HE951VHKaesm9mgMqIhpDVEVZv/DVaAn/cT5+ab/cqcp+E9ggsB
R+Q/nPOAs+7v2tGwfSphkxl90XMqdQU3XW49X2t7bZPanGgY1t3XjZqz44WP
UPqDXacy82HB+hFTRIW9CPpB6RAzttvZLnajz/h7X+LJwX8EyYzp2eqX/rZD
wbJI2i9Il4x1ZWV8V4dE5iHuAa59mvYs5JtBzmn8Sd4Lb+Qu/V6X5snnpXXv
nTJoAq3cqwlD1MwaQSR2INvJRTxQV5/Hr+few99KP2HE2gQBWpKCpLuO8utR
78xlYa9IHC95gMu6LEpGwlQmCYSvKiHkyPkMcsPHYDjEbGNNrHcHhj2MShyq
oAJSk0NEdxJpcedk47e+vSBlTCtWwxOiXgZopWw21jNe/Ed36j6TZuOjAQFM
/efDnV9nRfBLQbeMgYZDTllP8gKSNJONNxN7cwa2zsqm4YAxj1qHRiT9JgBL
B0j3XXRprlk47a4T7ckd/xYEb1PA4DU5BLnDwsztqayUP6LHVhwT2T/Kw8bC
HrM5jln7qqrspUjjpkQmtkHtBbCC7G9npIrW3ojzbvTXvN5viAZyjOgfsoLk
+YsmOy1zsEqLwe1B73UpTMLfum0fGRhWAYygA3U/grJMrW3U5EapDgtsoOPG
eA7RvSmxZfgtByKmBv/TCGJ3lVJp+e7kxIm5PtvknlC+NVYV4oiptOeYxk+4
PKuqAlp7UlalU0Q3WnG8Z4+DaT+I3lHIwXawXzEkx38w5Bqk37sv7U8fUmf7
wSyjVqCrxwI3hJGnzq08zau9OJsKEJDV0owsE3ta83ziBFmhS8gi0RKRiWZp
6p8cKVNtZ6FvVTkyHq9DCSFAQZSJx/8+MUBiM1cCEEPOWJ02a4yQu6UUd8wq
iPvVp2acLSbQvxJ+8vX5q47KO6suQuevSghHATOavePiLBN5fItXI+K847J1
hpDYfBvJ6db8LvBMyOTUINgXLwkFj+Ck8rvHarq8K0vAo+0rxaVK+5pKi2a3
78jDpzKqGZ3EngOp7x+9UZ85xAr3fszmtX44s88QDFLKqBJn0zHte2Nw4BeM
4dfX22m+qRhTIenl7FIcpUWbzOgmFcnrck1BSV7Agd3kd+pmk+cTzZec3xO8
B1aWbvmD7IBEepWhXohj2lnagJBP5qRpvGYMQMhr2yRIoJu5vYSyH1eAOf02
LVN0BIAD5Xsz5Le5eab/etKyhnDIDWm79dHEBxPSa9BW7gpuMZK4d96lmufY
Lr+whyA3whE555n2hullZeF7RFh977tmzv7lphYCF6Hxqul+LgCApfqGceZy
OdJqp6J0nRpVLrNmld/ZQfwn+lEQ+FTkTdtKPrhVyfOBdqGeM4VqgiJ3aE3y
C7Psfm41csSZi8MqslV+/Tkmg+bvN//gEo6IH0b0U7IcJD3x42+Dqdi1ooOv
RFVs5hH2h5ahB3010cokXep4Yy/M8wsHTUKNpTyr7WjD61HHOa3gylI1yIoh
+2S00IVfC6Gw5ff5vkiiWwSrHOuQmiOfeYPW71sPHcsLaxay0Z0+iobjHvsC
RAkHRevQH3abBiIO28T//FYX58fYpvSrlt7lmzftDgUdqHmTi2Z1rDQvk2Gb
twy+uZgkyVai5/RvFOUhXLOd2WQzzdmBHGbF34Ovri3ZBfgJSvfNvYClfmAp
Uj1QUak83Y32A4RcHzFDna7zZe6J3QEVGuxQ60uN3toq5+Sc5wJGEUM3v0nN
0nD+LfYDo56hq5cUSiCoU3juxScvgu6g7nRg/HTqpI/3fr2Tj4qt4JWpKlqx
WaYZWcnMpFzeeDvHbBUha01GjNwLun2q6snptyi1t/wLKVQIlKSlB9q7z09I
S32UhC0bvVX8SrehgUxU99wCKmXebQYkBb1uu0q7gwEDIyNmCf8OLZK1Bj4D
qOwPhMDZ4NBzWaOHB99dXL0oi4z+9X5i01t9NyOCxBOMQ1K9YwNmtsdf0KKJ
vL4a0XoT1lUadE9ehtumyzg1EP1+C0eSBdvz1umqjzORc8kjePZkg+XTPe2m
5FLjE1mHte1I17B7vc2qjs/oBJinlhqogjZHiMJKwnXOr+ViPcQARkVt/KUQ
1u7uiy2hF3lnRw3a/B7EMjJxNckVsZc+TlR2AsOgx2BsW1B5DGVUAgBX46J2
5qxFIKivSOEqggIWXZd9TizC/43OtlvnRFwrl5Q44QaVnZYB7tm+GHJ7Xa1R
qnffxs22KVgIdQwbr/BpOZrA+NJatSi/IF+7jDBUOAGgSyijLIYNrvG/ethE
MHrv22j2V15R1ivTsAhCBJw5whtel8OpV3sBigB6YOgMhT/zerqDdkMu+OuG
LvRqKNUV4LbbMoAZq/22KTWuv62zRJKSrXGcxjYeY7PiS/z4REYn+zx+6Ggi
Esst20ZN5uNihxR4lQqiBr80ygVk5I8nDvGVYQ8SVoYfCsbD9MbrbwM2QCtC
78As19axFFjZpRjWB7Rg+zVd4jWZFXtGwXKSkiV7+8n1a/3lVx4n0fo2LchI
BgsQzhqd9/m7Ujr+0nsmoYSjurtCvY8O4sQ9+9MvCwkHtaZzyh/7FLuwo1b7
PMOuZYJ74icRTPQD4hDQyUblo8J4Jsm+r+eRFpo4RpeKuy4aRII8Fn/Nr5M+
nqIv/a65+WBz1BTIYxM9Q2ziLE5og+ZyGVxnVz7dPwFQeYLashttL3QGht+I
TCS738QhmuUxbwn2dxlsEVKBkCAulfqPNXUjVfjYTFJ7KxwX1eLnhxePHCnP
KQAtTmM4Z+2gmjZe5ID9wmfxyP0Zhfz8O6u7azCx+edSwhg6W7W/05rUWLZd
ciehLfeTK8AW8s89Nu5/9TimpaJU2RMfJMZOTI8xMo0bNV81bfyJXt5zml68
PoyZG8w8R2sTevQ6R3zs9lUoAWiOyI1CI32ryYqhQaH9Ya7/ory2hRYUbvdq
3TFbWUeE5phIgRp20LF2ugD/kl1pP6P7x+Hg7YWXUpkpEPlisqrg+2BPdRxR
rLMX88wtkWKDHQJr4EBLja1JiCscbhfMQzJ7PC9MFIo4K/YzFu8RlPonsuQi
XzlJn8bQNakEWacsFFHgTHBKjiLz/jKYDF6QTUUeCWxVaLioIfPt5FgY2SNT
7aonP3Bco6X7e8ntaS2WIihk8DWxuTjDwS86Rtr0ouqIKV/710C2Tjj9khNI
MgDsmDgiSN6G4HZeY8/8j3novvvxFiEF9JJYz63Otkx8RR5T7CGbQC0GkE16
EsfQ593OakbWSRQQ2sdM9Satv9uLEAu5Hk80YqahAGr/Z5yaaUgMo1a46v2Q
toEZZXImLqXPFd5ofTASU6RtlISgkKjfJYMeSjYi9DdBE0s0oC3lfwiK794B
ItMsw1RD+PDF8KQT2tu4JlGMGrCq8f0eCHSpDSY8i2Xvu4O42ZHZUKBUOvSg
9+lNQOXz0eHY4EDralbD29j7mzwM2uiJKaIyBAshRMjCn3qSuQk6znIX3sNS
fUm0jRgMXM8lVPP4b0FPgTkjFfaDRdKTNks6GHAg22SrSLANR1vD/RkG3lMe
r3sN1nSZyUayjdERa4GVszRkpdOCQAtedct6AFlTs4Av4gDMNoGPa9vqodXT
CHsErjPz8cD9ApavD/qVAx0YWKwzX2HxEKV2zWLijEwMb/SQEezgb7bGSFDO
MAyKm8pAtdDAXF+OVFUjTZLfzO0dPsvtk9l0AAD0ng4ZGYa5gA9o1H1AoWTk
vD2hPCkOtBw38l2Iy8soRn3IE/FgWD/RThOACndzKmVYfp+VQcFvgVzqRl+u
tN2vgsMZ3IefkfH+KWIcHaxPgjjGVrbeQ6EZFU6KceS2uVWGScBOHWeQ9FoL
hKUVTzq6RSm3Fg2Cjn15wNcARzuPE3XDkThpTKpmbeBvRHsHkKN4hE6zsXes
JUglGoUg+rKGuq1WSZBlcY0zBD4jhkVgNA0M47bHBFKMAajWuaNfpoP/X/un
V7+zGJKlNcYejafX2/fWxMexIIUEjuA1l4p1Z8t3e9JC69ayB7kmy4dONHsk
yQDNDJN/Beqgi3eNuOHv7oENqGihI1FKXCltZ7tpvI7IZ9pkjHbyKYJMT+s3
+f4fk5E1GjVsACYU7PwcO8AL1rxNtE2YsVMP5KdcZq9PFkmugnFIL5uY1NDi
TN8kOAQf4I61kQgse+8rYoOwAME46+vZtm1EmBud4cX5cLX1nXHlVX9Plbxd
G6tL4IXCcjjL+gvUtZKmvPVoM0GiHLCLuLCvI9YG/xxy2Zl8+gnh6jpKXMsk
ElrKs47Gh02mTtVUTTmcmTn7/dQ6iV/6bj4GMJRWgRtKGDF6NW/rPI6uEXDQ
pyZA831HB5rhYbCf0O/DSQnZpzM7+GwVl1/PTTYBQBpKVHR8wxZI5JNxT15V
gSk1ORDgkNP8dyamzQpL8HvABYQo5KJctOjjeb5fy5t8z20Lhxl2upCJZZ+B
jbQNh8z6C5r2JHPOyXC9EDBVcnpiFD4blixvfhlaG5yLNHL50SO5M1/qho/q
slcz7zz0abMn9BngJqJbL/LnH6FutlnIIkjZP7tJnnIp32cvQzABWsE5AKa7
fEzP30F9Vn3VFdXeLl1mMN55+mbCnwGLzqEaDBT6WA2gjCP28lGL51mAv/4p
d4ZWL7Amu9yQq9tjDB/D9iesIwu07x/FDUIvtnYkbxX1u0NHtAGrTu/+fVru
XjsASYLDWdq5SR2RPwb4tLxDsc6B+qXjodpkJC/F9uqrWFrQbcHH3ofoiT4s
m/BXEZMSIiq3kpSq40G/RDhrkqy9CudMofnakUAgKbH/Att16hfScjvy4sDK
U2Lab5W6edNKyFM+igN8np9qs9nisCqPBp50qY9T5eu0eedBlu1++K9qjHJ1
zfu95GCl0v7Sa3XE7JvCYNr14wFUcYbbvyxcqgDvQU3d660ZC6Mzjfh3Ih6b
XL+oL/gExKPyk1Y6ssxTqCFuuUZKurv37OijbHqz5jRInLZKS9ih9oOq9L6l
8CfmXFg6Uh4C5rU751qGc4iAGAw96+8Yd5AjsDdFlWRfeH06ymtlSuOffCQS
ZKm1urGcFStvgqPWp3woo/La5gqF6xhWmGk/kecgwkLCpCEm6Bs/CmmCw3hi
nBFoHlNL/QCemrHxntXJSlz2UQdRBO9IUUPd8148N5XWPMVquNFl7W6buZno
bLjL0kCez3AmFtIIJu7Pd3qtBiCiB7xJMMf7oz3jTFerBcNC7KtAH7r5BUpa
UFHLFe6jGx35UciJqmCzeWN53xIpivEBv7Dd2Ac9ad8/yYqzbQuiVX28Xp3B
DNc6JULWKql/NnHy7c72YFWN9F4Y0aJ2xXtnCHljWk/M/xAPqGvpMqC3GTaa
vBqS7z/6W8XDCIVEM9Ek9f8/whtuDPA0pOSxMTi5XcWsMLaY2Ljh83Ku2by5
RwR+u4PedsWflw2P/qPMgaEjRTGcRc38DnnlymrOwwwZFo6g/WQQTXYitEny
2kitRRs8cYwE1z0H24/x6PKNv3oiHGN2Ct9Y0aJ/DSMqh4/XIIGKXHu8bfwG
ZVssu728AMjezPsjDl5LAT7OnLA9U2+zoloLMf7l/OpqUQO+wvDYwP6w7miN
TDDd1V8PIhS1YQb3V3Gy9VdavWRBVMFAyLXfOmf/fqKI5Kmn1gAT/HOOPfBf
uorjDkVLWrksHNoLcoz9zQWd+3B+G54ziJcs0ZV750/uB/goTie8xBQ6PVoJ
DwOulzQkjscamjwJRwMxZjfEVDD99EMAkis2ITAt/qqCWaNOCc/hN7T5JvjF
pbV9o7GcKLF1BuFPY/f4NGMm9s8JjbHvOLpZEMC23YpbrLB+5h0cn2Eu8+5U
LJ5xK9ngyYtBoSbMSNXmx4a22Cc2asFKMJ1NeVjzSauGKvo3WLtKGKhxsb0h
f3kX/5qHlSB0wp1curFY3o8JKyRnsxAEK9mjQDfI6e+7n3X+Mmsj2iNt5MIT
SnE/I1Z7t+XA4Ev00/Bf3un6zNXySK88Bsqruz8XCoNozzV7FPB7IHfoBcxc
wD9tUIp3hj2vOswBgg+65qqF3u1xJ2lDcoLSNPhDH82wdYcciWbdWEXnmmBj
qOdBUUQA6d3eSAmnLwPz0lDRBZDvHOUDsmonVAAROH8xfkE79ButftUBukWq
wvYZLtfnN7rp5ValBF7TQSnzfZZa7BnjQxH+tXPzvfa9jIiIGnq3yVAvrCNQ
5ntDOhN8E1pNt96gLhug+RK1Sr4MzY8guEOsZFY2SThr76Vg4CpMGf2SEzJS
Q32HReqWRkHKCtkkUlWQ2zmDK15iMd7T6zHX5edS48YcmwCmSMtXMjSlyh/n
UBq3SlvVoEkMOtBwCgoy8aPyfJ26R3ylSupkm5XQh0qs3/a0btmKAxwR3dg1
RsL5J8qF9355m9bwyqO67poDsuwT87ZD42JFgQHl1lh/GSjcCRrc4Ov27ueL
Wn9f3zXN0Wv14XmtPtPlYogwOrU6LV63BpnOmIF+EZjVGGs2K1SD3kclNtbE
I20Pp6L5f4739hOYmwRbNIHtenx2oFBi/N54IIRZ/qyAea8d6sJFdcood+T1
SYkMYPhtG2ipH7HKQOWTA6xkwa9AvnDCAaEf5A7pRLw6ndhTIcG8BEdU2uC2
O57/8NkPinKJc6h2R5Xr+Ydq4CyKl9CczAFLSw7rfY2VeQXEe1QTrgL13jpz
ufBEA98jLtIzZWV+3XIKURu9l4VcXV3lmPVOdi0h7UDAmCzGZxEwZpHpG8nr
wIiWxS0pKZBSYh+1PTUo5jBYWHhqm1T/zOQXDsb8Zjq1+HK0lCu+6Av5TD2N
zGRTosgI2KlC3xAz9MKVRNeFZk3BnjqQPGMcK57ZYW/2aa/84m6xycFIWLtH
uS39zXIrjpICNtY6qOkBkoNt0ROJOk6ln1uRRmhrCg68nH/fl2l+Up/rUHK1
NpS4NzMKcmdGveIVleVL8Mc82iTf9rZRx6LfPXxfSIGoDqiW6p4jwptbqzWD
HX6t54rO2DwuWXepM1aeYP4iaP9BlsfTxlr5kjof1I61fP7oX4G7NAG4UIO3
imDt+Gnem/KTonptOyV7WtK7k44ClOVFGjM+Ha3fNK0MFBKELi0/w4SAwhjD
qhEEhShKrO8S+aPibWxnmJZp8fxw414sAmzT2OnUXy/H+DgVjXpCWdcXdxjs
bBkH6kTKZbErL27eK1bahaZLAFuOJLY8pB3b/F8RuddubsshUUrsmFwqFlyS
GHHfiLdLtkBnMZ2A3+RLjfQli0A0mpTy3CFL2tk3OPpSMA5V68hjlJwj448D
fxSCXchPQBn+Mia7BPdwu4cLbJ3s8NISOs9S3jc9nQxssxMsU9Nr6Uc9dMkn
wQ3gVVa+5MpFiMuGPQU+sMOlxLUpWBCnHoGqBBi/El9uF7CbTxbuebpAFFNr
LgFnneeuACRAzjq3XpJ65U4YD1d0WlsUV4mx2fvYJzDXRP47AehRBhAMw+2c
MPBJMuVeFI6T1PLmoOCmqZphKXreCi0oBYScCnDUWu7awHqs6KTMBum8PDy/
ywEqkAyWfi+883AZs/y8G3eWxhx37l19WwoHiNGE9V4bkk5gdVIiGCF+lCqy
/TPJbYrAXmXlWx0VtmB2wPj3FMaqQP4uWw2C5LLr/M2ZbXkArmV2r6On0ysf
gdAJ5x/BT6NWS+K7zcUDgT3i9fJA/3XM0p8FXW26hwj5vTIZu4FXkR7c3nA5
/nAY3xyFF9R1O2FmJp2B3Yi8OV+ZJaCI7675afXBbEygLqQoHtouRAZ4zeV8
aYNhYNhSn3XkY8znEdygKR1uhbwwDpBYdzG+8CMguH5xkxL17x/3tTIq43ew
glJ9FSFm3zE6rzPouLHIpQCl4I5elVMqxwLvro++RvLGI2UslZ7edxHjFLCQ
3NqAcxA2Sy522+xU4FK+J/53bvOmOYI0LPozEOvXl+OWJPcLk1LZp8dXN6VH
h+JRei4/DY7BzOds5dSt3holNCLBF5XwcSVm4XpNuTsPrYc5bqbcKPByret3
8Hk7D1H1mLNtEqgpJz6KJBTNi9kyDl5jSWv6R4/pdT/hu3iqmCSJkrFOXa+2
TrX9vzhDSrbJaQKkM/99Y0FR1u2hahjYB6DSfy/Vf+MQptdAzVQzZoVUH9fo
NTA8Fw84HFxIBOSpD4XtMEAkcEfo9qF44B1t7/+I5ZhRHZ2MzF3ZG3hOlPXN
BzbbxNmdp1605OBmdkkOS73RPm3YQ2TScZ+lFP1g7sPI823nN3Edlpovf4sf
xTUa13Q13mDPfteX584Qqt49VmdjdUFx5ss5naRwUyDc6egh8L7wwVPUtZus
dW5nwasDc3Qg7lfopHAROAT/I5x6jbpF3lR7es5ZqtMtEuZ2h32WWdVLvouZ
I4UbdkfE+J45LXpl/D7qkC+B0pxCBgxnpAULuxjWFX5Kv1x/rt+E0yVAl0xv
OKhiZbOtMmGqnhLbIMuV1WUdSbE0FGzllLsVP8mOU0VDCzVkByet5tgCNBKs
8kYxqPA6/zHpJ2SC6Fa3gFcYFgkdNWY9uvAhM4oVQaWQi5zr9EHg+ukgZdFY
qWnH9XwTEWDilT3hDf1vd/uWgJVs3mDGnh2/ZYAwLTudQlLApTZ94pXXAyfo
JXU4rY76zEwJnriY63b91fMgL7UdZfTvCVDvukhvJNPU7YDrhEAdSE9z+/z9
1h+n+0HZ4hKLlHvbT1EeEIiXYr+5D3xgQKpHgZmSB10KPX1WxDV+ttmq6wiP
m1kfm1jakSddlcSPa7gDL1cBQgeRy895PjxO0gEcE9MMA7TvwmtOBCkbCLt0
skcA+0A8DHAbhfBYDOXNI9EWWq/oAcu74dMlpJlekZ9ny/kqBqv2R9dKtNR0
3UxgpbHGCku4puJpVdH7b2KnzsxGbVdZXDIRPcPJ6HWDblPElFjd41Jg8ks8
usf5cO7oJzcbZCG5x06kmzsPlrtqKB497nWXatViaF4lWm+HWhKsVzu95pVj
HTgmUHgc8znv3BmqiPJtzJzOV6iPwCikuH7m3FwnblnNgnzZZcFOlk1zZVQP
pWD1jF1l0+rekwFN6UXjUocOqV8qhxLtr8CPF/PDCYb1gdipVEhBmiFT3IjB
/ytVbUf2ga/dckA9lNB2zoL5kZcmHV3j6pao38YBC+yA3KvH/mov22GFuPXe
1QYNuoDqTi28pnDo/7fwLQClZBGfmfZV3XFWfa1N9E1h4+ySmIPx1NACYGzb
HCLL5uRWDWkBS9FJl+OoEME6e/Gjp9kmbR4ghg4/Z0sA7s1khXJBW6smaEPw
WtUFUqL9/CHFp3j/wsqT1Y/oUgGFzSPj7KXuTfGxZUMcwvluK3OWHfoZzp/p
CGu7+gaEPxLJ6g5tznC0L94rRMivCuZXVR3lfHM7hP2Sz3UONdMQd42gpnYd
4G+dhzfaHDw3TzmOsKMxmD1uhUpXhOQQYvo9gIzV5NToVjxFz/BzxR7ykp60
h2YQ9xkOcyyrIGkmR7loWZlFNx7bEuhihUpxJaCDam7IxXgGHch96n6tfTIE
ZNwOFosrWsSh96IJcFmYchqMbG0WkBbsR6kUU+NYWLVanCTQ/HXMHLxUQG+t
uXsEDuEyarZguZY16dsZEpJdCE2ewVBu0hvZBI16NNvTGXMnAHwPoWlTF+Cl
9LSp1mj7mP+qDWHzhfV3/xquATwcBQlEF+z8ZY3PuutcyoCmep5sKSsC2uJ8
bw676mS5aN3p95zp0Bbb4+fIqG/H5AxoOpITg+zhBliDzbq0Dm5XCt8UXuHe
9FKhpA4Rwd+RGI2Vl/jO6e/txqudcQKOpZxTQr4+He9kVlCFO4urB/gghlvR
8Y7SxgRxRMZUO/jrprZPcx/yivsaIrcUGHGemX0yLAOrFm5Opjm5u/EXNTKt
jE1W9hb19G08PYoc+9csJaMEYJnzca79ehlIXH/P1KDdRARstBAvd1102gV3
nUUvQtOdK5U/y2W9Rhbwkjd0031CS7lz2ZgPLRqmDSt9S32A2Dqhp/gYFUrE
srabXOKsFdjTYsz2RhoewLq7F4hQYcYKCmt6yzH5oK8LzIK4KpePhZwECZXD
cJa7boAPri95uZNDp4PY+fL/3rffzTya32k4+ZKalNrl45iAPB+DaSZugy0s
2KCHlID94SGBaKt1tuIZkaNOEfFEfrHoMn17wm3qa/Qrd8JOdYZxCPWQVNzu
yFFdHfj8Ba4cQ6Ox/Sixk8LoQOWF2NdKULwYOR+SMS047bI8FdSYr/vAu6t3
XRWreNiLB6Q3bzRW2RydQIhezdlBA5ASE7DVYoMUSYYTwpsw7TKljq4sZ8OQ
8q2I0koBe6z2WNEoYLN2ZbfaLuPURZf8buY/155hYi29JhqBa77u5yhll37J
NlEXROBF6jroFNAx2rOLnGSY/fM7AZHgT2TtdkJRj8i9VoFuaEpHJHcCnWNc
MPs1QenH/DzqhZQaXrnozKObFT4nBshzzsZwaVh2hmrykIFCinD5MOB7b6J6
ieYsLl249nPNfFND4uI4aCZXRXrUKnotGCbXgti1uYfgF+U/XsXf8zAqKE5s
o3qw2xQA7y0JA1ybIBjB3p+RH+vA33pdITbwACPMDlhF9oPHND5BD8J6AAP4
nrBCCUUDLDU+nvv+nv5pbaqVM1s3S+s9bRRqXFyS/4OsdBZ4tz57gWDfVECM
EtnmheoXeVeZMYbwi8xHlVD8zSDNhwZgL7kEdEqpfpRjIgxybPdTlRZuRoOh
H+FHJov+y+YCgboq6hMvnUa2lxa1J/IgVr0sqzEUZbfvacMTo3E5/7F8a0cs
qXW3/w99eJoDr5mz/xlE2uycEVPD9UeJGdL9jULrxPhWxphOVodeGpDm/Rjo
FrY95yz19kuWl6fpmCs70rGleglh49Vn8k3ikYjvHzoeF3qe0P4teLwLbqYU
AQ9VWkTJUG/gh31IauOCBScpvuUqvMCMcgtdrvFAszRAS8nnEIgiZLXPZb7L
YgVv8Fx7HdbKCzDHrt+ifeVggpY/tgxSN8fkfxVYRJef5puSHmQR7xteJr6B
l2EX9wTbx2yzN6vWG/8IhoTeh9jD7DbaSK/RXtvo+M2F/g7SdZ5v6GKuZjaL
9cnKrgMfO3MnrDYMkrUQnAod57pyavjUMEKi5cDel6Rn/tlWK6FD5rF1bIke
q8GVCWXP7iLWAsEKQ42Jn1eq7l9/UE3K4/Ls1h/UXwxUrbPuypr9dOq+RW/G
IEY4+Ru5z7KDOOpJabWIoO47rQ0vWhFnrymAr5/0tEmgiE2LLnQmS967HUnm
+Z3Ii3DXdJUVqDvf7MJr600xzdgeC9nYq9MOU4yNw/6qoU2dzFjybRnhkKXr
AZDP1bzwnBIOoo1c3WkUmOqXaPaEiQj9U8UzT6lZqppE38eqoMnTDyLCWg3K
bDvTaDvYkP49b2f00AbjEXFmXwgDTrw4aASbO6Jq/qA14xBQvIJ/5Zc6Rgf0
xrWAhtfv/uSg4gHZFIp/ChZqOBxo8XdSySByoGTFVp9FNfKSLvnmCtO5vhBA
YvT34nl4xFfwDXx3SnzPa/1SynBL2fVgXWB372ROXBGGwvMOTdYuLkLuis6r
qHpiWR3WRToIG0sXk3Xz7iE2lhtkkNjoFrHtm0THLylAR7zvN9/3KZlz37it
5QWjvoVLbp49ZnswNmyLTRJbChfcdUHlkQ16gYtJV0kpByiL3Cvo5gp6xEgU
hJFNEBZKikq5NDNz60iyfd2o0D0INCNC+4OGx7Mv0OtjZDbmIMXevDUDGYGl
gB0lzOHZblPvFF0Zi5/NAlUuOW3jEzDDqyxHNjRX264NEYUQFBLGVffb668Q
856Z9FGpxCreEs6fD64nWKHpUoMoXwo6njUIs0Pxk+gdgoVbp4QRv+ccu1Sk
NCQ99fOJrsECdfnSalxCyWo1uFE8kH140LpuSejnMbhALLA7Kwv47IxIumFH
BhggN4WEvAe4yjuQylKFNg6tAqI6UX9HqTVs5A3ZttqDpmhdEVSCw0HeJyDG
cyksNwEqKBikardmtjU/cQZmdIcu/xRWzXKyx3xgWCRLTPN46OSZ6THRktIQ
wgV3u3GwJHtxO0ydhloKeUrX7NssKG5XmWYAA9w7EHFlAx7giqoMtwfN0QOJ
WnuZHc0NaVjIOdmp3J7dki9m2ckRDIUXC69O5t7knEnTXr0D6nWmCDKC05BN
B6e/kVKYNJDPLoZ+Z8rDNk4Rrfczy9u9K7dW2Tg/8d+J9dQsLt+8HFQVL8TM
yEEDs0T1j2m09OCkNQ04cmqDnTgQm4Igmv5utpTTO+ixwN/epHEvL3eA/Ck5
3I8V39OQTLJwRVxct+aEzYI7PisYM+6Mt1y5rmLH7xppDQ9tV2Jv7W5B1xBA
hoCqyiEmxOTNrZSxlGM5KuwENYzFrQPTx+sWzd9EimVg7E4TsdhV8/5jpMds
Ep5e71+DMhOGPAsDt1H5/KvQxocFQi87S0MZtP6gjn7vj+NkjWNQNCvhx2/N
vu6bZ4alhESpVyqdoVIxFfNu5G93vSMG8jpaN5jou1NSSgKM1V5Ra4F5hkZu
kf5UNmA6TLljNfSINR6bLrSFL5R6W7FCeBXA6ueLbd2DTzNI8h3Crrr+HVlv
BJBYlUWP+BobwhiQ7K+J8Ve75NVWmwKtQN0qAH4PWdDq9nxN6y2kCxE0OWt9
bbz7E0rxNr4H8FMFAa/V+b04IYLr1sgYWHHdxLenHRqv8vF9LgzYIUAUYX0b
R7nr5dIQ1EoKbR9k+8F6rZssAd4zKBYPU9rcE3MNP88lpRtdlqqckdfamEPS
0HiAd+SfLKFVM+lggoN3Zn20h7GxUIJ8T1FoqhkRQJrA5xLGC8wAqT8OY499
pWCGHMdAajay8kQSsO9CDogfOqS3NzZ8NB4nFDPB9T1sn5gRGaquP1vbJMmC
FY2QSPshJrCYeyRTrYMvHmE/EpiSevgLtc1xCiRUrV7IsRnpCGZoXPECW3l2
1AALND8DqseG3YxCTwUHGBiy4QvZNmJFzDl1OunSDn9bHtitJprMza+1hud7
OmugYzKP0Z0tGUh5kDhmqMxhTIpM81SBGRL9e64fv87GlQNbxNeb4fhDAEM0
t+KFOCzOWcoeGZATT1lKkHQu/3K57Kk8boSPBKrLDhxjhMKyQabYmqzUXjxz
OdrCOWR10+yDoDiI2zPJZjMqFYpcUHnE9AwcoZaIYPQ/cFw5TxMxoysdweBx
T5jTXqW9UdC3QDzA9GXtRq0m3X5ZaOlWeio6Xu95LgCDB74KSOxhP45BZWYm
HW6yjbh6M1fDDmlGJpAeuYibPuRE7g/taH9mYMcZ9bRLRQtvEhy3V4yuagDO
T354tSZcLhC3Nw5v4F+keBV8bohlhtHauE38CZK1SC4eW6T+U7MnqVD/zp0p
tGGa8TvgvL72s8xOQ/N/hvUOmZE46m3LOOSAgYeMCn2jwtQ7n+vn+ZJhvqi2
lMnENMx/7kMfi5pSmWI5OJsYCeNIvi8DBKUrKZBeFqFoGCjA/JFHoInuoMnG
qlQjiYqytcBIokcQbQJx0nK5nt8097CIEZJJTMzD/KIVdZdBrwG5iYoxrGl6
BJ2rkrwa4mGovgYhbKrJsiqUrTP2YAjI+728AGZc/Bn0/eGZGHKNN6dvoGKo
HuLdXtsx+955CGlBFP7g52R+t2lN79PT+kgWt+IF1tbrULj+D/FZGxKFeusj
j3Im/MmU1VVhoWkeMVf1wy9N3lwWS7sol+SEkmX8sgfDb3InwUnYS5TmIV3Z
d42+stATCg4Qtr3NNKmPWbtfSdSLlHe9xPBVlwUxQ9IanzNZNr9X5yZPDOjm
ki85vP2nGKLBdm+78ky2p0ByHcLgMbVCLZVCkzTpFfZ1yyXjo/bg6tu2WCSV
VgjptvYrdqh4LssIJzdhOTVOhCbuVNcVkqgEcVoGx3XTgg7PEDi9Rvrn71LO
5u+AJ817Wg0KbK7vmCubIAP2Iz8pEP8kEtYrUwGt4Guamn5BQUbah9aImp3v
U2WElx4uiLSEQ/kjHJcuKITu12gb61rISIAkJ/4RtzXWMSQemvx24D+ONhBB
6myhPhADClz0LKx1/UbBuElulzCmkMhlBRHB5pZErremsBxaMMD0ySTlbaVG
Tqt7B2A6rNkJ6R3xZwJtTVhX1b5ANZsfnahOjKqZHbsC4inMr/xEeFXKVXH9
Qg5LTM9Mlsmq8+6Nen3peL4Q+gwpWL0l6GOqxPyTuKZmQazoU5DhQuoSErxb
kaePI1ipkdqrkOcpgam+lAZYWY5PCIxGi1kQ+zgn3oG49nSxpkpOorgIWIVh
8rRkAg5PMNshLuW9ip8U2uiDIyi0VSrrlnnB04QHk1DXjicWcIT4AfJsvf9N
T3xT/udLGyWqLf3Um2iAO+ym2ltDOvYd5/XIe2+Gjs2Jk240W6Huz7MCEek3
C0tiQoQF+wDLgEVEq0deWRIDpwsb191Pt+qbb+2tLeimzdPlY4b9yT3PSeJ7
FrMxNmVdQGCYBdVspnxnF0f40Q+58Cf277Bu2zBALaMv7enzluLU0rzQ1fkn
tf/9VOLvF00oqGlyTHvLTpCL4iJ848sYYoGePopuTAIAs1i0W05pqoEO3lOE
RWCJfV0/cwSy7TPGJLo6thRwbkQFdW/scBZSIahrck1k7cZGaX8Z/bh78ew+
PCD7LmhQTUrWXnLi1tGVJJ8Q8TSIK2oiiOiFHcow4OL26q2Xm6S6sh29GE8x
Ql94QU4HNkFtbh0znLFvA8xry1DgMmcELczj635jiENgQJCp+f4vlUykyXjB
co0amu/VMOFO0BiZ6HUy0hF/CQxm+Rnze8nzP520bkm2RW9YKweom6KzQbfK
aGlt9vqEd7o9N/cs30+7wnMNC7QKS3Ltv+Q8SJuYhZWGNAfsek1s3KMSPZol
C+1rWDdkHwtHrcTxHSMzhtfK+u4KFvJdoriDrhvdYnlgEFtc+9SRcZksAVXk
4QpRHfHmQ4u9UMCDPz01xC4iie8qHk4BStxTWXhqySEj92SuHNvdmR1OBMLp
cwD8x8kHI6vF+4f3zEZIXnUSiohRpvESMahMG3rH87Fn8aYBTs2ySGjfQ4kj
uf7R4L4/Vh4NckuLD2VzMxbgx0qDvKZd6VNI+yFXCRpkn+17CnsMgdtt6i1y
jQLv6sdM0wYrnn1Snt+YE5Y4GY9RZBntxh0nIpmto2epp67nrzkPYOuUgM9V
8KMRYM8nbN0zMx0pAXzyBycPJUofqbRkUMhIdypj3qOfLzE5hvKJuhAcJeif
YqgTY+VeTxO0dwX9Ft6MlSGuToydAWjNdOsK6GtAZzOCgbGfWgepDg2PTSvQ
Q7oQINH8f65CPENmxohPnafmcUilmT89vchWpXVpg8UWQ86Fob04JXBeI0XD
hAgjAGs3ayhLtNB2euhOsXbRb4scLjX8VXwhzoHCDW+6tTD3bJSMUnW5cg6p
fgfiswCCjCUc0V74tZpjp7GvPdRZ/zk99v2BI2dnbHFNTHjqeicmvfcC+I0C
kOThpbKLnWVuwf4LABdG2LFlR8xU88dWmJi/bXHUZoTaLzz15MtMDEn/cL9A
v88VP6vIS1/M50rZTkEUwIRKrq/gtJ7tkGITXogi/l0PxjyPDBGyWBsprFwl
BL1nYGd9lF6r29YogQv9+oyIJPzp4h91VDJnTH8d3LHodkB8ppkKJM2bI6Oi
GyaQi4WjFgq9AxgrrtXNVRHomNC5rVx7o9BSEyOHhQAkgINhymZ9CgJht4wp
5V8tslbaMfmSUAH9Ux2QbE66HuqoHtYH062dTUItK6ZYDlCTvueCUs+xfulp
1GADL6Dli68Rhi5dFQchUfsRH+IMUDLMBbkWTEZ9hSNmIdzOL7SjPbSvIZKE
z8eZonv2zGYhbdY4Iq2e4DcHZXV2CWv6AnGV/JXHlqwrPtXsAuUy43D/s1Vv
7M9zdaI5KpavQ8BOdEvCwgSsAxKER73cc63FR0xepmsjqRwoM+CGK2f8NFKY
tCThXuT7xGsjup6CrCRb5erzwoXWUnauj72mJQ6gj+R4uf+IbT3UZdJEw4P4
YORKQdF2NG7+nd3YhSaBzuOqpDBgHknSCorzsYp6B/grjJDcvq9t8kpy5RfB
OpR8Fg9q2UeLuA9EC/sSsGBzczpXxstv3iMvtHH5UXDRlzBzpCMBluE7FXm6
1aX0t6OG4d9RuBONDu720yjYIKfVvaxn551978/Qrl2WJzw5XHAbCBy9koav
cvYwI30G/Fyjr0oevKTMJ4PPZBtRlJqNHmJYuzsqiNQ67ANZ4OaMPhdGVh6h
rnlMrfis9FdcSgE3seIMXGMefZnmhZ6OdUDaAH3ID5knDRc5GIhOJtBxtTW3
Jhq9pQ3mqTztgnkKfMUmtgdWjbMBB7gCn4lPMVrP5/iWjsGlbTfcWCGBDwaj
p3ooukiQV2q1SS2JPF6clLKuJxR7uocZWehFxmSXSDRngL6ibWlwGZ7RSq9M
upJYQ17I889xKdYuigXtriCl7cs/pEufAGucJqkqtbyNgSXpf+7M820ivSFL
cs5Lp/Nf8HKPO71mJPYrAa+hdmHGnoKUG5ka1KDAf+WTQvHoH6de3khY1cB/
Bv/LJuesNcnwu4YmE4t7fF2V+o5YiD2KZZeJU55vzflpdy+DvGT3ruoBHe3x
e944+YYvz1nOYH+7VEvPgAOr5hU/+w/+SPk5d5PNl7tv6WY3uw7orzq7LsvK
Q5BM3hk7zmQWQAoh8EN4qrW+PM/AzSnvt9qevO94WHGIx5Zcm3qR4qnrRBcy
KZfzTOGDrrVof/7oEntvYuXlfosxb2JU+JZWJs7P3urLvrpp/2e3DU3eE7ea
JoYg4Lir3+SBIRMzcTztngGFdy8EWX/h1BrMeKurnacvKFHT1GyIIWQgxxxo
U0TQNjTJG6dc8GLXwQ9eEhJwaroWhovex91EZPcxHQf3Sp46sApnAtvhHxHE
c8GyXOSgPy963VRqgE8fFSO+tIQYr+hi4Cs1xtvtmU/k36LaMQcx8Ray81Ba
xfn/QdNaz9eW3hBQI4ppuvedHzGDdJoQnd4PSScMXYMGWRH2coN99pg+vHI/
tiwWTN1ijgpyDb0cb9J0sLhI2V+HfRwl0yC9gfbRp6iv6RmAXf1gKYPCuV4D
XUweWkrfHfT5jz/whopWyC1rCHp0uGSyU7uieeJqVeU2RhxGpjVQ1uv+Bw7+
y269PiE/vxcNUZmYxpraSWdhEpERdhSVug0nGt/ljBCl/qZGva2JZK1Z2lun
A61bj2mDqNXvrI0ECv3j5n727sanSvYYhGghF4dKb0w8Xesc9sEDD/S2i4Jp
Q/8Z2jKAD5Cm61blEf4wHgafmv7Jroqi4xoCyxUlD5xwxl50ESd9of0HF2Oq
gvLIhVTL15vxSmmI2t4TNeYR8G59Iu5nAKuy4R4Pk9fS8rtYNboWjpSOYe8C
pLtC6M7rWfoKBuzqKcI+xXKMFywcf2/uyQT6eoFguuLV8lK8Pxbjj6eot4LG
FIGDSEqziq/yi2ZkdqsCA9RwXkbmsNAUpeH5FsABFZqrtBNmTTEcmwfkVssI
AAPSn0V3mCyEf70hcUTqJSWB+HKHCxm1I5M6GJ9NFYSlsLgNgKIPvq+1FxZB
rzO5QS2mNVrygfMQkJXTh/P8E9kfOQQ3myj9xi3uneSWpkKhhzM4x/n+wmUk
WVVott6C3xZbf7vSj6/QYIDOS02hC6b7d5ucmtBRm1RckjAl+PKf+ApOEPhZ
bmemWus4u2MiVrirgizTjlI4CfqHur7cvp/oEH6CHmRFXPl0GwsZWAYeh5FH
ieBq9oGKjeZw8nZfqxlowJXRsa0yicVM4rL811g3CWJv6H6Ogej/EFVpLO7E
kN75dSqweL0qeUrvpXJG9vMs5E3yikpi2FHJNYa1bSkHv8fscMLDlCbxQbe4
4ibSWPm0CbUxAaV7aQtaYbfgFQdPp+ATDMmqxpdKxEmzL5RptTqJj50mCDIM
L16q7Vp4v5FJ/5hScHtUuM0N59EvwI1cpcEmE6U/N1tmy+E4N1lsOYwNVftG
eTVocgVKbGjOGNdC5tebVhl1+5soT/96MITm46Y3+jx319EZb7HfjmfsfUdN
s3kyGhiD2/tNcawbWkOrg6oO3ok9wIXl1o9K5hfnNi3XrDWkCVwbk49vA6CC
RbHEiL/zLigBIdeX+9U+3nCohDuyBcFmz7R4mcrTP71Jn9aWXPeSsrcNgrgi
Px9V07mIoDJmv7qIATmkNCHLf2eDM3Bs0vYvoPUK1g6k1ky/IeAxsL7ckKYT
BP5Tqx2A8hMHlrtwwOLinCxhRnK7xbGsdCJqCP6UV9s8EvxDXLPJXwYcbuqd
LuhfnSOlPSmhjly/56H8nD752RRxFnkIl4SGlMIuGQEOkssP3vw7C5m0w8qi
DPwxU129cNCntyvVZrbsLXidfvJHWHGOtTeSI8VI9wFx0clNQ9BcZ0uO/7pQ
OZK37fIvAAxd7YLGIy9t753ZzXyjmrv49ntNzit2oEqPPXWzaPFx3JZOhCxF
sjJibWpc3CNIzOrhYf4BACLJZPe9ZMuPQ3GUqm39Yh7++3SeSjtmjLJCiLBl
eaDxF6FxsaeKXqsR6YMjAFb9qO96njQte/EYu+aLWDVLPMZ9ou+bvrnoJiZ/
C/lPxKaruGB0aG6jud3tlbw5nVJHpIbhn7De8JCiR61LPEpAlevca5mwzO3u
yAocWmAjCAJJMR8tWNHkxMRsM3NAxoOlyKZ+ZKmMBpYGujhzSSeKJMYjhbqK
B/ypb3XmVOQcnIi8jai3wluytjI44meshG5SaUBg7mRCFB92U+b5ygo3xneI
9a5CLUbviQfMne2rtj6xJmTy2yQSXbWOIOgyGAta14icgjAuVFVHxgktLUlP
HT5FoN4E7xEZkO7FAVUIEVzsF1ADntn4Oke7T+MANwMm5uKYouGZEz+sAk8G
276XZdCQxcY+UrpkOaUYRrquMmGNIxwHqGNJJUKYOdI6YSDJW3/gOzfpK/K2
6sZ6+axrlBE997bSd1bkEg73vXJC6SKq5uqxlP3uaHx9iiyTJ6BFjzITGoAj
iYIXXBL7lMv+sbYZfsWMBV8/nHL6QJYmJFSZi2wAY0pEuO3G9H3sNk5tX0BD
FrZ3KWYQc0g4PQr5ZAquKFdanzSyK1r/nUAiBPGFcQftxRWugffQvnLVgZfY
M0UPRCW9QL8ncbb8mQ7dikQy91sv6m3nKbGISV+Qw91zSFd0fjHmtUD64v50
yL4pY0g/lb6/AhNp5Rh5sgj57kYRkKLylnO/g5qJbxZ61sC3B0+WZNC79mjw
UZ6hz3/ObW9ieCLlU2TAe6MUxJv2fPin/PwHo/NsRhUCeZMHCBi18VV1+bNp
KqzO3XUhOqxhjZjCL/pGBnuT0VGt+Vo3zj302FFnhWbukSfnghTDFoPNAsrd
uuoPH0wodmsky7fO2FH0quJEWIaYtu1lruA035nGjBQmmv6DfQjazEdgmS6i
aRoDKXR5IJcHr4Jiu2xQ5wjcSuIv2RwJMQfRDrAhHGW+VklJXCLQJyIvRFG/
zqnnJFYnD6gvmWT+Nue+IfHMR4L0sp8lQbdc9/brIUhmzqcvCmRrnfA3tS5h
QlbhjS0qRDaX/SWIl1eJgMj76k1rWKec095UzVVB+v8B/gNv25xSw0POzyk1
FCmbnCn2N+aPL+t87eZ9503fZcIgK03SLmCg8PlW2HDSBIyPX1NbCp4KN06u
3Fxkd7JxqH82NUWG2/El9YG7wHi2kS92zAWyn2xUrrx68FS04EpP5RFU6EE7
yVcnrRc2S9/g3Ur/G278FEmJxUhilKcaFm8CqtXdWpw645VuojkoLsjyi3wD
RgBdIg5+zJqTZ7FyW4R6/4GaWLi9+wtZpU1+6I7sP5Mw6gnoG8kxJ/427Hgt
ODEiJ4ojZ2GSkkCROxQMoIr02kznvG2Zhj3CUOWMrdVpMA5uE/Uhzt+4UKsB
SJ09LM6G19q7Gu91JpZVKtuDNeBxYq3pSUjoVOneCVpLGrczjZhqToWm0zU5
Gug8/v9GoaXeuTBY/uruL8lDEFHa//3Hn4ptIISA5MwD4qZOlFDFOzoJnCWA
EI8fj8gFPiHgzHX5DsWHOcu9P2oLut+XFZNUrt31XjAJXvaH8KlTbK5sxsRU
Oxk7IbSqYqW94BoxGAsdacdZBz57Cm2MGDbIN7kJo9MH99S7kiD/ah+fcazj
uyZzK/POxK0fGlgPuc2wJmQKx1LTr9FzSDUokJrPOoTFq0/6U79ZfFVA3JoG
ttqoSYgCLz55KsBd9sj2I6V0Ex6gxYnxrXTrujoW0ZJyYtn2J2hJm63cDTxX
4TJWi8IKoaLNEXo+NlFcJ4o9Y8D3XdNMAqjNfJ0n/kgh5Q29aMGzfMCzYa/8
QU/PqKCVlDU+/VJ6BOSpELXb54BczOhG8/rIBMDHz8uEOZoS/7r1F/YiyKQz
03DotM26z9KykQqiJT7dax16l0xBAw4N9/uUcOnd6QBi2NYxvvF24I8EB//O
ftssnd96r8R3tddFYoSzVmp1YFRh4/GpuIjy6pGT5PM9LoZnovJZZie/G0Ud
RBMUMwojFV0nrhbmKSTiM1VOwccIG28MkPSz1fsuc85cwwXFmVpnrN0z/xeH
AlvziFzZUO+nGuflN16pJ8Z5fPvsOugjFmhVyJdJKzzAO1R7DXIV+ra4fEW3
hiYzEEW/Lxkk+Tpsk4AZiIA3+z6FsaTSnOAzx8R89ZqkL/QjncM1uEVbAPxU
3zRS9ZOuAf3TV5Uimw2Lp4DBj4RQNe5IUhDLhrSW0jJwL4dBvFScNsvWMBJ4
+2qWOHn8OkUkzFrzyF9UaF350By5OKEUjONmI5q78t1i2L4xGKTkAYnrk6J9
wkizxt3KYjPjDQXBcZknJKRaU7VoFXzDHCUpcF/kD6AYc1ZS2uyuVhV3dcrH
2AvQa3zMvRJi+jNQBw1pXjGEOKo0y4v9ZzAMLFrXB/rjitVl8noieYnc+Ous
O8p3qbk7t1+pY7jxCpNKROcv95rk4Si4EnRUdOP8l1GhfwA5UYJkfzAtOqYJ
DTYbamIZuRRvI28go2RdRxj0OiOP6ihC0pjQ2EErlJCrHfG0yttmewO8xR6+
88Hz0Tl71jeUFaX7SjpOZX3+E7VzgFn0cnvlzXb158lKLnOJpWR7kpf27OEW
+5CeXg1BAC7e//g1YIYuHgRCqjZsr/ERJ4WAjOVo7J6paYY2Oj8jnMlwiCG5
K/ocylJyAqxpo5kN6h1Am4immZPHwVFepilDH+6/FuXpDyC2ut1ajX87W6DL
dkDI+mCyJFyKpU47GdR5bz89c6rrcNz7OPJ36gYQooJoQGNC3DNHmIVG9xCv
Bx1oX1pxB1kQDOWRit8zXc1T9VXdE0p1hvhfhCtRi4QphP8eR4N8Yu326IJU
E1nofDK+qRpKNQfNs3ksoXlvfrH1ZtVd0y4sXBYCN/OZqNZkMHIBm7Idrobk
OAohvsL2sWU+nNPZ+P0kcNvNS8BhukLvB2CB0LbmaIqHgCzihr6XQ+3QraQH
+Xa/VwZY6xEcrypyuqH5+YkE1lT1ExepGtgikQql+mg+WUdE9sam50fK1qiP
/KIx1MsdoAUkPebUvMKK1EkFVuXEm82a9ibRO5b81epc+Y7xIyuUSkOH60fm
VIQWFsPpJTdhAq/igUe2H1q6Uy5ga8QkfJW3dHcxoiEqksn67xx2wwD4kSKn
8BScD9D+GWkm2jlf3NLCgYDUj8KzJKiRw71hCQ9mWY+o3QhHEF5lj8E+aiOE
8cBZp6FULAD63QlXeP21m12+ELwswgE9/iezLcFKifAo7JkYw2sC/WA26lDc
AEBJhCyQrKa/L/VuwviHDP6ts7nZhX1jsYD2H8t/qpWgv4BOLeaaHie90pr8
iXZJs4Gf3uaUHMYxAcclmBBVCdZ9ArflB/56yp3SEKC437tj2fyhzkwUkiGV
Iy4d5Pae2mR29qKKXXDC1PATEyFDbgw946t/JPKqK1LCrd5L8RrMQrbwQzC7
ouTJQkneMBo3Kf/XmNzmTZ1uIkK9a4a+KVQdpPgzVSp3Uax6ikwLsIaTpDr1
xg1KG9jygfx1DZyTaX6r4ec/4fOaYQrQeUCTHiUSPOlidCaMjRAbInjOn/28
r7rcvQQOkntZupQMym9rmuYWWgeNfmOUaHtCb12Rt8WzKBCuASb2vgZBbNvO
K6I1IWFQTi3PTJrY/EUPN5L8D3SUQgMPOKgVQZ5WfobHhR5v9lvXGx1/XyXR
OCl/SPps1mp5id32YyR0du+RtjHopBzouteopKfRy3NbGljGAAd/rNul841z
WfkJRdwVDULXFFLRonW1Z3vDSP2g+LByrcCQtpLrrSEOhrAoqaGl/U8Ek8OR
+O/N7iRhoBEJuEgP5uQ55P2qzJtDTB468numyQI428VLskr9CqynYOMVTxTf
udZ6skh0z4vo5ixrOOfNFkTkN3dtPamL6tCgEWCNjYasotfSxfuz5bzIkgNP
CCV76Qmhh0jfXVyWfm99/Qtbdb1fRUnqwl5ZAdknIF1pSHRRNz0zl/DfB7jr
UvH7AfOYI9+BAESrRJiEWXh4znEgO+P2hmlYG7k2w+dIu7NJ4unYixLlkvK7
6Ve0rL9gQW6xMLp0zcfkydngIJ7Lqicug+7SXf7JE9Rgc6s/Ep7t5IMPcnuJ
OFwyqe2My//EkcuxXLGXEu6/pctXRBqnqtgH8SsWUm2fdH7tXDrfx7QyyImg
c7hGTBhboZCgzoyM5oxuQ877eg+HyhS7zvtiz08ex2xyMfurQZd9+bkwBne9
/SGIV/e4KJFFZsxBhrr7b9zc0/7Hz4E/q8fgjphuFslPJF4gsDfK1nMeishS
a/6HT0nftF4if/a8/117vaEjml6O2zTjwo5y9dqw2t6RAPHXUY08RsN1GUW9
nM4qXtpiHOC7a1vu7nlVqB1xNnR7gJ0wJM0d2Y/3s3RAUDJNbUKHDQ1+6b0b
1f5UiY8n1Uxy3SQnfincDoLK2/eNlsb3jAq9j4KjJ+wCzOBf9yAlX6lZdI+E
AC2y7HRGmqFSC8rIj859TrLo5OXbqblMc8tLZvFGc4gvUpVY5qWTKEl5Hy85
TOpOk3NR7JQRZsl1xM3Gh1Z2Ot5llVB4W/ECZzB8/V//9ylZvH6J9GF7WBal
2wyk0TqhtzqRo4Pwv9OaosKI3TEVdUNSmHSqCTMSKss3/z3KbQB09Dwmwono
O731R5y9AGXfUZmriev6XdwmxDjTos62MrE6BO2lDfCgDnnp1mx0wjNkqs1s
vGJZ2NFwsCc5ElUUlyJa/I3uLJKUgrVul1G7oY0AgN6G0I+SORgzf6tdJs9o
5R2qor7xUaPSZObLlf1oLG0Zd2H8EYDJj/Os3kkBCd/gw8rwiHaxrfQabRVX
o+4AuhSvQdw88M9xGHnHWvSUB2Q+H8uVd08AHwiVUflIanaHGUBlBWB6t/s4
Fv7hy1c29sCXbIEHoXVdkm1oGsIdenBqUnayY0LMXit3RZI+RzbojSc4l7NB
RHQKwFVUWSNqgzdCk6E2nLIDeOuXAFdQiGMV16hvhWFJX8QAxmrxAuAd3j36
9KuRvDnRDvblAEULUGUYHvDCFp2HZ8Nnk075R1eVHC4+o9VeNYHVX3kexZua
HoKHjQGq/Fm0ecXweobuWVDXTE3xkWqiBJ+RudkeN7AtH7V7UiCTmVULQ0I7
dgVHHI1EqZNNemoHKLNjirMiRLaqQmE+kl4JD1OxhAQJTww77kdsEYQktZW+
WJ+ZK0pNQkKk+OMYmHBWWhbeRSgOI5B6W/hz2bcbtoEQCYqfHVeN8RzcPAxV
pbz2i9jY28/yUsjJzLLA2KufqxvCoLRsiRBP3SY14AK3qhG7hNuBj1N1cK7M
BrL99CEqZsSkTG8FK5XiEedln8FZaZMTJc/FFS6v/96YxEyxx+aw9jmq1Zjv
ZQK+o92W3mEZUyHe1Y18t4y5hwzwmimXQ6r460qI5KC3v0qKAu7gyODgLG80
aNczW1TUmTrWsN5l005ZuXGsS/CK6fHjlaEcdiWMMslKSGrTvXgkdVB+cETT
Rqc8XP5rFAmSwCkJSLBPjqL+JuhuEzLx6FSiLfNg+zytQtG7w96Xe7/MSH8S
1Ld9CyjRGfT4xm/v/mPyC9K28mQq7WX+qKcVlRvKPVeySSxFu9HBGnuDbRU/
q5qCH1JuNG0iVyj3kYDlUA35yowpi89gzVr6xn7GcblBqjCmAc/ko+t/0b9R
h2SitgYRH0wMH27W12nGTgDwNBRWz7QMiRs1PPX7ZDjm/9Fm2lE3xzQNdJHS
+DA6TkKANKPvX6t92ogOhg7c0Pjw/8YIxAXcQuOSbr2yEwNJQ3vkANAkl7i9
jWYw2rJm+1GPuuFUuaUWkRrzqg7V3vHhSWNztRq/45B3b+7rnPNvupd0b+AL
hfPybV8Z+S/mzjDTmIebVo16OJopidZPOXN0yFLTSO6v5NdNJfy2p9mGvCdK
Og3zuJmY7UlSFG0Cwh3ZWdLvt0KxzcnbO6ShpaQOyCtN4BSpI32LxALSh3Nw
fatQZjEd2E2n2zGZE/nHJzsdcIlOXoQE6uGdfqxLrigK/t4n0825QQH71BN4
JPWS7A01S0m5cbCjWcr/zF3ODVK3LtGrMDoruvJLjP3jJRlR6yQltImfF7G0
pSC5YU1HjMNtNu9bvp9sIGjPaH91KP/ogcRLNGzRIH4J4XmoBy33mk4yVfhH
AylmbLj4z6Tq173OFdZn4tP2ICOiOF6jdh+ai/WdVERgPNiFQdjzHTM2VNjI
6ZYxvsomo1i6IEy1x+NwVpc/yi/akEI/BAvuMsSQW35pyQmoDT5+rYF3Z88b
hYu4tf4yEkfL1TFJoQmtAMmjX3HRpUSShKCoM5kYj3OPCvfDOBdDL0YtMlWU
Krc06Yp3ouR1CG9SSCm7NBZEuzLtoufdGuXn3nLx3ZHOO+kSHpHKpSIoU3hz
Nq3lGsLSU603Ou+qPVGf0vWtmsjASlKFhOjRIrsNbHzyWlFPrgocZTn06Jxy
0eUpkbfv50unN2Wqa1XPHGwitXWd+sD25hnl00sVOOjOfc15IPwkLogbLlmm
rxi8eWzK81x57wZMKygTKZiqkbM+yWwBMSMTPM1usaYagssWK3dJ9X3DoWix
ohooYrja2UueBXijv+UmHKmec+0vLlxbHfi/5Dsd8ZvuIRG8u/Y1Dpr4k6At
QO/STGhNHkjeG9i9LgpzfLpAyvGFsuQCrz9zpl/j66oRa0Jmp+ozd5pBSoot
Vh2Wm3YayAARRXtGkcDKcFq/zIioSkFnV6waWhs2wYy2XFcLCf+OeBJCv4FE
KOX/EqCukHI3ThfVvCj/g0jsCPdOiBcJQXmBIHR0ztlFfJjih8JS75m+uArL
f2bpCmGXe9Vjhj9Y1g2JXLz9nypL/6MZX0qOm/o1JN0pT0DbPtRJlnMvttSq
urK/jmD4DRgffBXyi9JdUDJZGLFj25HvUll9gtfrNKQg2x8qShFNdb2D8qkR
BXyKD1xe26GsoK124xXOymH03h3WrJo94ZDdIUvpTtHL/IiCw4ebR3N9ARAW
HIIadKmdNe1ajjALXJxp8F3C4Ef7YtTNxVVAHyQW2X434uUvnXoAeawC6Wfu
c5vm27B7oElydBI6SkmZTKKOtzb2gBxLBMqe6Sremn/tvZr9lQggnvc13WZt
H2iZLpq0QD8hhleaVvEOEjUwnkfBbcZHs0Emd8umNJUmu7WEOiJODYJGXgrX
8lSM94TyAaTY+3OUarZWPOgoWl/xS+SoUkLTHDcux2KPJeCjYmp0FooXRcwy
y4btptnV/NPfLeO1WV4YTK2vpx22W5/EFROplWddutFa0MpZCCMSMrrWpEpc
YsWZo/EAGpCLO0H7RssrwZFhnf+cLgMrveb58WjlgojgqFjgV0o/eWb7MGdS
3pAQEe9FHGO3t/QPmPsLIPvCip1VMbyNAxE9p2qtfvPi87evlKM2SiqiUdYV
fFjZSRlpDcAaJu9soKuQVXM4y4hEOa+x4gXtTLTF3INygNrjfMTS3ijqKqWm
hIaKWaILaltZXi0rJhZhq5MU/pLIaDm0Ic8osFIET6pDQZJrOXUrubND7H1L
YJm0fG12LtkG4HuqPFeYaZaxRyFc0y0GdbjAXEvxXZ/TtUJFqkMkDwcH0Zjt
mvkSWKooM1jHsgI8tEzbm4A41784iuFUR0LuhX8mwtfKU+Uri6d00l/8nqEX
71zeywZjdrHfdwJr3Wme8uoPQbZtV34bd910AphIOBiUSjDXtqhCG5Y+bFMi
TFe5xr4PsiAYbki5mMD5bmljyQxU7XIEzxVmuwEcQVSOlfOoo7YwuF+eDAo5
6CYpLwBQ5KiEDUmV0xsNcBYpxDQMJs6VYNtbNGjwhsbeJyjADKuC6wL3z16G
RNq7/ctf9HNIv4ovh3leEmoCb1BgoWDKBzpS2aNUC0iQZasiNaUZLxb15UQW
30CHGFhk/PU5/RkLGf04X0MTMXpyrrBoWad67oAX5XjEeiN89GQOL5B/zJkG
7VLyE1uYfhHJCQIRWOnUwA572Q5/WMkiRaL0pxhDt2wuGF9XNQECTyZ3uD1u
0xL88ND08q9agaRdDX8cQMniF9o/gNwLS86Xb6ipAJIV8XUMdf8nX/HrM/2R
5/Svus2bP2HK2DEGVRW0KH62Sf3wHiycy3PNbARVm28m3tAEVV9VonW3qMYe
hvpDyNA7PzTv9JuFw8/SscwkG+JJTHB6iLZ3LuUGu+3KhfE5U/D8vi9YKLYV
E8q39JA9M/Nzkw71wfVr1hAqaZ71V0CzpkqM6fQWMpFKrt75nfY9ubC0xcYR
qd4VlXudCTZobRFrr8jeOKe3RBi2EfiA69tlLqrnMadC5At6ICN/17yjQ6QP
WmPSAGfsAux6V8DDwZBo4lh2DcBSc5UG4ZheYc+awR9dYhaMA4FNaRzacwWv
O2OWTi66O8ZZ6gDnmeCh1Wy5VJZm9s15m8C6oj89J4va9NgpEQr0mw+Wgupu
0SXaWe7KJngOlH7+urWKAbJrpPVy/0ff+Ezt/FwXM7b+U/yUsqHZO4kPqQ+E
TsnoJyo5FnmSI4aiVAmZLk9IVpiw2U/FlpFSQinGz5sI+k/Ng3NjO/HOtRkQ
XlNkrEiX4if2NJugauHL/fNf9u+MV/vFSuVnjrbWgOX4AMYg4imK2nmnq60i
YFq3ICO8zf15qjSG6sbpuzk/mHZMA9uZyOTdzR++KV9KyQ1TX7sfOPbl25R6
DG2ZxmMzxCzHqEeeIm3lGdz2NjWNUFkuCIGeXDXCzGO687jE/uWJ4fUj0eMR
OeNG3aDewpZvwc85DWMynjlqbdhUvS9+reBDY28tKHcZKbnFPVZUovVdYJzW
+hGgNc7dHzwl7bmrbAVZnB7GVgGOi7iT4ZanJLUAsGSAtuhVdVWoCj++9cvY
wL0TEJ2d+owSmWwejaZNpLhUWwq8QN3JNKtmGQq38tx5e+c9OPj5K0rgYPxN
bvhCjhUpiRYdQ1zFT1oEpF25krs3ZkRjulM4gmOaPzmoQnOkO1V0KDj83MLQ
khzTbMfWgYRf88QqcB5MNfxIQH/JDus9NAnMA6sDf+CemKbCjFoZPW5cgzfj
RnG0OzzegEajn51A3ZmTVQ3JXjjkZ+wnjYEGvYPJsTwP5/RlwwfATiBKvWAJ
YEvJyHioeQfxTEyP/j4iINcfr9MEAbVCmWPsVWyy4kmkaGknej1LpN3CW1ax
rWAAAcy/lJUX54MfHuM0I5LdQPyvnt6YNsuZhHwrdeKRsc8HDtYRKHp+VLeZ
+K/BNLFSMVt+GCFuxsXDFqg/NYbHzzwertBMjPDR4fNjhutS0rUzFbk0/Pgi
8lbnGIBTArfgUXjVkhxUUxgqidfu78dTtOVamPfBhmHlQmNRO4C5IZuqHA+1
au09KKnwMZMSxGzwME5ya8HMa80dkEm6u5g2BOgKnUlN5+hHrBJu9JnChNDd
r2b5/8R22D3HRYimSe2DIH8OP7dikDTHqmOtU7bmImh/H0IWzFO4kT49bxX0
DiYGD8JtO6ZC1AhiZoaP4E2j+Wc9MSVqUBFxTLtpXTpP9wt7yU3EHTWHF6SV
Ga6uCwVj+Uh8WC10mjx0TcJUQGpjKzGUNXmtKCA9UIgm3HNRvpkUDpK3ErTE
Q9J57CoWeiILN1RhxoPAyOsxYOdcFZUOWOEtfEwlLAEzWqfxwVGvF7POz07c
tm7A3AXrQL7XrLggMfVD8xhT3AP2NEyT12KLZ+bqkFXnO6EsozjLwOx6KKow
H9OZjbzLIAjdcizL8/cva1emwWzsEQ0IO6RH8MKS/A4uduhy0MGCG+iMxhLz
Ttf6laaFFnZjl+7oHTKAgzXOCrgw/YCcv6bal0+kT5xSxruTos76OB10Om2W
jeIvqHn7eQQyqK4hxraIv1HxxCpZb9kv9nWMCo5QY7mkSU78k8VNQ9h0eHpV
yxQQPVZy5pZ/XRIU5zZorTh7jO320p/B/GLJhgfzkt+LO6qpZ2GfHtPZRsRK
WeNJaeVSsJmX61syvPcxvtYKkSvIVn3FSG3OWejZnJo+8wsSWlEWxftjKZ8E
jkNSfJaQ6EusDj0O9TkhHJNZn5Gk1KPzrSafPr6T0q377Qb/pwmtz5EdzIFi
ZEO/IrSiq+vSQH3sQLI8XDNg2cnCJLJeSw1PfcourrpFt44Y7hU2EOsapeuM
aSBDTGHKZ38oQXCrtz1HGjtZN9KPG8U1GvHF8ONLKcoqmP4wdCiilYeMor4u
hWXTcxVMUTcyfcSittGt72SGw0ecGAuvSL76qRYsTqa0PLHtPND5XGphHwBy
8kET9onJRKkhZnYTReFCkb9MhtQBqhJAPOS7+sESIOKlsoO1eVy/JTq2wz6U
EfHgFyzs6E3ylj+6+u8WU2X9CW8OQYxvNN7JaAyCc0VH9iSm8ImD36oO4dbY
Gxoble9bwyb8KP6PLqw0P6PGjABqx2nmE0nUKCu7lKdiCEb90602k+sYSZA+
iC0PQvy7dII2zNkFntlX7/o01VlVsa4rr00A7B2mhl0SM37Oy6GZAGy72I9P
xroklpWP3s6xcltaHjUplRvTGIK5ji9UVtPmtfQ1CdZjGYWQYXvD5tDw9Hcc
lbUDQZz7JLVzEhQkX0QPV904EVijezRIwM8Xx8LzXiLX3BBKQv/1BrA2gOE9
7ytQ3Wgw7gFfKCakdgeK31nK/C3B5bK/Vdy2l0SocWeT0dK5sYaPvk29wBce
UD8t5mblH5f/7mbBaW2AG2VVHTl8yDPugFXMu+9PTyVJeD24y8u5rcXkOFyd
+WB6llB9VF0YWeXq8uVXyozKphwI36Wu1Z+1/CTie6SQBlfTslwDSWsoMvEY
rZoNiGsfPsqBdnC+yLC2k5tiZxfLJYhkYGcS90hm8TACadHVWv1KNGhsxr7S
hAPrD06Ed740zs93iK7kb0ssoSHh29NA5rE6LspT4MX2y5CEiNTYO+uH6Cdg
6sNreIPofFUoipyYOUX8RJHs889H14OPbuT4sTXvZH7uoCKZi1Ekf/mmrPtr
vG2rwkeA/tB9kMvZaSqjqBrKO/W7WtgBNkmlfWIfhtFDcZ/8ZEyMl7hvT+hj
pr/ldY+GnnJ06Il949io2EeSVTjMPlzIDN/Ki3HR3aEX5FoCzDdB11xkn6la
jQlrStU0xZ/fP3hALje3vFkaPQDhlXeyTl/PYDkKoZafvgOZ+1dle3KWyu7L
Ht9qG25Oaqry1JwC9/EU62lHazdqD0TfzfH8ZnNAnZehh9BoeLACJk2SvKaz
uelF8J6H+R+Ttp1DSJZ8dptar4I9WgJb6ZIBvhhoV2+FZl17QHfAmaAMeGR8
lgWUke0XfpaUkcS+OTW3bJqbe09+QHIsrf0EZuL3o+mqXhbMotDxJyMm+e4G
2B8N44AyUag0oi2GWsVU06fquE4Z31AJzZ6lTuqzTPl6HaajI4NxDLBkLsAA
LZ/5APjSPdjnsg2aowmvyM78xqQfhcpGj+IEvsSR7wlfLvQ17nFT4zHKno4Y
g80FHxL9uHJT1Mt2JnPo+22PM5BttPEZ/TL3dm37ghX5rLhXdt1jmPDUzAiE
bw1YFd9TyWV5LRJOtZ4ef0+1Jt4aJzii65efwAfyNTofK7TfpS+HpLIicEqg
t5uj4NNf6HzHXYq9Un2eNEgrACI1aEwgF/qYiYidfvjS6SFtXnSymzSUtTxW
4GEopvQEMV4Q2atsP9zejWQXOLfgnrZWa60CuuudZpS53zpzWQG8iF0cL5Fp
a+ENjj3d9Ax+jCl3GUa2VR6X9FULQrwBx3we0ABu1jkdCg9ePTkQL33wWvET
QbPR7qJwCHe2yeXy4T5g6KBKCpsmfRoaFgfObpmjd2c9gXMIIw5AKaFtDhPw
puu3XIH2K7FY+LLeVd+VsW47iid5LP+mte01q4bAVZFYD56dAfJLW+5FuuQ7
NzsIaOBU14t4ppTUnehYoFR5lGXZjwaKpm3JmIdjRsFQvDvTQkjM0N2Kvtbb
EJMSnhezFC8hpmKZaLvMZ/SS9e4/LrGjXUbpDZ038rROyGmzsbfltZPKHZ9l
Z1TvvBbT7W3rETErk0kV5dYvz/y12U1gaecAt03TUh3RLSDUcNOLtLImAyUJ
cXf2IQPZsRjRN+08jXTXGIpAhuhZOXa5sp+0mdLT1TlysTcX1J4aaEmU43Mp
gNQOpw5YekzF3u5+TVcaagkxc8YRaSlSzDquPFDKd9jufVd1x+GEBrFFlLOy
1Q8tyWh+b7Q2CLH7HhYfKGjCRDbFfyxHCWMzOQuqou+u4bcUIR6fUF9n4ebX
9+Cscezf7wX74yvqhxoKb/vH0ayI2O27tX9UxZ7DDofNIgkjEu52CBvAJRxb
FTw=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "B40jvh7ud/ahkCWXo8CJP0S9JYnc5+J2pwOdONjrEnmjRzb1YpxBEP/gM90XdEQFf8e+9j+GJABVN1VA/EUgHmy986oXHU6n9uJJjaeBsR8h22iSaiy//95eH4kKFakRZgkZDqWp0dX7AUTwRg4vZKk0rom9cx0xsiuc1Ki6fTzxDmmuuNW+yyxk/luKJogixDl7f05H1PhFx3JTfD9y6cRFGovJ+RtyYHOBbLpk0wgVQdQ/xcRbIkbM86PtUA7Wt5LLc47Ojn4KEAKv9fZmFbaAAXkEhKb82ReRoSZgk7VcZ558fUkp19FkHMMVJIudDCgQiPhwGZRNXAJW01pbeoIiu1Tf91lhbgzgi/zdX1xYAtyEDGzdAckFb2O/hhjpQtAjVQTv8DgjN1HpPLsrizivOWUAXDsdoSCxWUxwNgBPj3AaD9M53HUaN33XLvwu73kz5Urkl68WSk7MqyVmSUq2/VFXQy2RNCcy0+wkE2WMCohtkWDcN8G25xEzuRTw/3NEhnhT/D+gD1mClK2UKfKLf3D1IQBvOCJRqkWntZBiq6/tKWa5ugbgkCSoO7b1qXUNZxnur+AWa9hVcNoW7YTU+xcFA0cCFwHzb3dYz1yREgu3Vw411fREBjYkKL7+NBQXe3iuWEiJ6QG3ldpF7bmnexSrG8Nr/uKUnlO2Zk1S+jldk23QtUYyAlUZSMjd8vTnQ7UbCZ70OgsoVr8EJy2BK+uGD8tRi90cl90n6eWq3OWAG6Iz1dGZdeKs24z1NhgSq7NpEw23K4HkZ9zTX4+fuLuf4Dtri/NZQ5ZCuvceIwiUdDYg09LY/jbFqi6gUHwn6EnFedx2E1/0irICZeAI/0SBHPDOYJLaFXIp6fiKN39YGiH2XiVeGmhC3rl8FAw0aqdJXdHGat0aHheM+fzM4cG4EMhRs/Ttm7wAZYt6vvfRgFGdEFUmbtrZHY+5+4rBoOCN7T5UGGuDUwwTF97HG7yfqc1RhvrmYAsQb3mNfJ8s0KYR5zZPwsmqL7up"
`endif