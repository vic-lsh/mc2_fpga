// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ddga4g5B5Bu1QSBC2LWrVpgYSEMN/tlq6Jom9SranLAzagYhrIwlhL/bZyvb
uj61UBMlC1DEvueoJyc8BwhWNgQIERLhPBvyjiOdoa3MLoi2RTFPnax9vMwD
ADgUWAZR31OuIJRVYf6ZMBTESbm0NYlrY3tlhOu4rr70yxzII9loHnD+J7KP
EUm9MbAy5zR/bzKFgJCRflnGkBeiKBozYJhAzrgWhPd5Dhi1nLbdUvtayBvP
4xBuSOe9vt/Lrxdctrbk+yETclOY4VLz293szCydREcsomi8IzzxF3B7uX1g
/uKkDB23jwkV4qYWwBDBwwZc8gJXiNYCrFdwTr4XgA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iysoux4lx0edDiGegpmQHoycDkP27bAlvHOMzLH0Ll+y3Oh1qkc9x1BE3Wn/
MJVi2t12nIYJsBhvq72ujhon8NeF27nQh4e/90ikTrMdktOZ8bO5Z5OjpiEO
2BCsVG//vGLQJ4kmwQZq5K8Q6vdg8+DR9tn7RXREkc69yZt9cA3TB/TN9JFd
krchTYUDl/XtFMR+r52JOQ10yT1Xzg7gmniqr0FE8JsjYm/fvg3bUf4r+zc3
kSexOJtWPg58l7oncapkhKML2IpRDyfqS2gdh+UAugTZ8wlNCLb5gnOs8dPx
i9355PMLZ1L3mKosw2vJKpI6UETO+0lGWEK3L4Zdzg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Pzvm0sWAXxTBVQluJYkPfHtdlpA99k6YqmoRe5PFiJ+Fo1gybfmaLXMEzMmc
Nm51dmkLN+cKAAzAc5uEifuXmBEPXX1rWuA7YjMkIjtaNlP+EW4TNKayfNBf
IZiDq0+BhG/vcOMrXUfbksyngWvW0ByBkAbML3YoyPN9l4v2r5nBF04p5PLa
Fg0/ILVDZmrCjclyJ9y57Yh/8wCa8fGbvLAioNeqkdmqoXlN2L5KvZf8CDxj
UoCt5BLOH5MzfRifLkjuUsEazOllXi5Z5tNL3r848U5cs+CPR241gxkopGff
Q0V+mcnupSeaN424sTrbZ6LZBvCBif66hSfvsyWIfA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
p4eaWFFvUJ2ilZkl7TzUm2d1H6FoOeBfHHrWxl+uQJYoLX9Z9Sb1mKszWRyX
vyF8YReRDbmE1oEYi95N//aZDZH/xVQY0y0B/yWBmoPnOM2ARrND20MQ+iU9
ttjS8aI8s0Kg0eWZcjQEPh1eD49Vp4fKv9lu/CdKK6a2bRoCnAqHZ6vRvmyi
3mRVsYcR8HkcVKNPSmu6mqUd5GgVyrnm9pdotQ3jotlCjdMjjTWTV93zRA+A
KKBcupqPu3suXLHIJKxcyi/GEIvsWclG5hFM1OnMrz8+5k6fE77WHJH/aSt/
AcdLU300H55XTzawUNKMuDSjVPnsxw+TQWmAGHf9dg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
m6wowQi33Bj1frVB/XbWjh/tqmNUmXfJ6wHPHxooTZXPKuvcXHq8BLw+phhd
GVt/wcqGekwGBPMhvcWhx8GEJsgjzxxIVvD8C7MiVlq3MwFhx2LElwPm8OYv
lxsVJewQqLBxv9I66+zsZ1QIz7ZN/R9m4y+WBBZwSrfYjamUWro=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
hsIbdzLMy1PRz0k/x0lpJxrBroL7GZGGnG7QiPNo7dwKleCruNPxHHuJAeu8
eSenQpsMXHjGERZjAuQLyhJmtlWslVWnM/DEq6HxPG/+mXNBbzQGxuxlSWpr
5eF9yyRz16XiOxY+HvFhd49QMS9QEOzZOXYP/Z6/Rgi5X6Oqp9T2mn6JXVTE
tMDq0TQ6ea2z5pppanxY1aCgVEdRitsOw0TwhTANLxHUz8Wyb8XLTSu+Dvpp
JaXoPOtTssHY7KYeggE1z0jtapyU7L4uap3yU0SJfSI9HSlh81HTTGmHE8Va
PgKHQ19h/sWEq3Zb/1JAoE3xc+Q6gwFjxq3uMgEcbGkaGuO4lSCEBCAQScAV
Z2xK4oJxgIu7b3XnRGfSrUgfXhm34S0bIUV4Rld2sN9XCa54Zdo1RyWCMhX2
dNjaxEdtR18vb6sdxoNzV4luNTri8VaZOXBdCyaIfR0MaMaFhjbx6VkWVGeK
IKWXtVJ5NEbkXbVJSmoxUKEu+/lDWiR9


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LXdrtv2t2lGLEb02YQp+yN2+Ey+NiwW+UGSp6hYTcchT7ZmdPZJtZ6nT4Gxj
GVFwu2ZHqb+JM9bXvEmoz4axxHqCBVDyGjkaUWSLXsjRFgQr8K1vd8qjAF6o
l4frMD8x7nQJx9Az4Ncz4U/kT5i84Kk50D3f4Q8nuE6h5d8Jxi0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YRtL+vlTM0fj9No2NgLrfXHha/2QZ0l3+JpzAeljlkejNgm44H9RNbSLO4wM
EMVltHpr2rYowejZEyWgwkRBxMtJTrg7xSIsFmkjAvUGVQpWYUBzJRnPiPNO
hJ0jd4ZeqXtdbq00FT2Zgn2AV7+vtPHs4gHHurzHvap1/kKqnq0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 67280)
`pragma protect data_block
znKegXJbZ/cbRhQJ6YYOneU+JcBd5bzUk/Q4X5a1nReQyNuX04713PPDDiDh
1DGGAZEmz0Xti5WO4LCPOoeBuRDjEKqYt4gpNYESggszgPPRzBBM+P8Z4xF3
EfqBXTN4QDdDTcrdcugWjgyTKPHqyO/P3g2HewQB2v0cBDyZqat6Ed0AHDiE
TL1KeAZ3XPCmj8u7BEwURgPfsvNE9aaRfyB7BerMWO3JOtuL8SwfKM4reqdq
i68t/uaKFkFFNheVLFK2HLd3q+29bRKURJqB3tLwDoCcXH1jvX7zpsv8gg4C
ThEdZ701W6hf7UzeEU59tRZJxe8zAIWwcwMxyMoH2rOLhyKgnULcSpId/3sp
N53T4ZlxLbY0Q5dkS8ERQWczkfB4ahCjOjfPd8JxZ1vTr4+kv9Y1KEEx+IRf
6oqbFiHkZ8N7XC3ougxT+DbFj19/CynEOV5g34xbld/oKzE/uXLxWMJkggrA
RrqhpVrGuX1ZvPQPuBop0x4R+gi6ljGnoLRTmtojuSCVovN0GAqDnOQCNe1+
KhfBLOeMj7naiWUriA+0KmVWKocc9nereZ5HglQvIsckPV+Wojnuc7i5MERz
Z3nJwuj71Y2iPXxEpmiltXitc+thHcoH9oFHi5fuw6HUMzjBQqZrjhwSiaRt
eHN2VgrZYbbZZKvdvMR1oUWtGYOvY8ldeOddjNVeX2WtTG07BeDWy3YKXrbz
FpRJMKXhOiXR9ffmyxruIrXsh+vmpg/e7UFdl8WZ5c2BuIXWqfrgoLYdr2bi
j0Lpbbg42oGEg+D5F+cKYSE97Ctx0vlbYJMVEkUGRxi1kz/bCg+ufdWidoNW
XT5oJzy0vvEWtdYsI3rivt4uZ3iIW0d4jyXCuwiAi7KQdhToEBrpCh1BO43b
/kmzrlMKakQTuGogTcMFJeeVLdEXlwq3Z9gSy3FEs/fvJKMCLoB4ZDmYZJyq
a0seB70H3QUhfV8huk0urFPAxOICuf7I4lm//ShJxyx14MKvFMBng3jRQGWj
dbKVVE9McgFWbnl7bg4T3rfZbKldVPovy2/Vx2r+SA9ZSy/q2MtfXDOifkuk
M47QR350xUr8LRWX/TGTo2Bbc8Od+xiajqMWzj7el8izom6JlUpy9hUwzRoI
dzXVcNofu9nKsyZJPepETKTkPPobcG0oGi8bIO3RbyHIftAxAoKZVTcOIyU+
rC63Hmwcmrmkr95nTMEJCpWRcy023RFjTBDi42NbpI+BG+T9lG7YK/+jftKG
5O2beUsyZIjotq0PSc4OuyxHLrTITnTdg5mq6DDR5B82h16BILpaDyOkm6ll
Hy5C6cdt4kwp4LBYK6G4evelT1kzmTz1Y8xclf5gL/jtXTFT0/ybhAnlOi+I
QpMEq4SYD9bxYGKg8bjkXsEDnKuW+6+zWA68KX8AnuzxOiPU8wGoptgCd1Zw
8UOLxF6BojpzRk9HKqufvLxrOSfAxE1f4vJ2/IMQ+5l/O5eexjxulNVDYAIH
o+JEpzoua3HPwgB9ZzTVf2DZlWO3WCD/5poMa6c2kFNOXgWw5Qx/eHgO2Y+J
T7ieoHTdiMjDIiNdUFOxUKwQ37OmlgawBS2s4EgtpgcjLfSFS1ocubqq4eTr
n4dWTd+/pog5qlhs+lU7YRRQSA/8T2ynN5bGg3034cmFzfE/c8itp7oqf0Y8
8LytpNW6AaQDaL961XPdiMyo2lIBth5dkT4bNvLMKY+PIyId4TltzSGQGUQu
pdM0wn0VC50QalNZJuJTd+IEiYU8ZA8oGVxfifX5gJuWLF1PAnugTvvXPft5
q8lf1bLqiq4jZvLz1egbBDpmCMz36qE/omV3B+r/oZvPGo+VOm609YEmPi4Y
qnKU6PTQxknhE/35K3SPt+87FgUoKZmbVcuty/+Wdia5moGT4nivATJWXEtT
ENzcQutEvNc5l3BC7mdWL087RHbov6Edz0oLLS+Uei67MozDop3r5CkipdxS
N8KSx5r9hBaK+JYcnpmppijX4zvTHjWN9sTsEO5cawd8+k688u1L9YVDQqqO
lpEe8dp51vguTmP0K1JWiNpL6bjz4nKLnm95LJFQArjteJYBMCzYpfz7z1yA
qhVnTwIXR+PwFO6B0aq0P4REOfyiAwbsBwH++lOpToEXEPVMW+MFo4u85siO
ajlCa/cabLBUdMBJm1Kp1GlGHjcPsqiewyA2cLO9akYwOX4KFzxDT3pXI58t
+cuHikLDQcuJbUIV7rtWj3Eke8WUmDBdOraIgJE963p/04G0BJ4em42JJVp8
aTYKYUXcdezDjMhhHaKE/XFWWVhOkDbNtoO3MSMs7GJYnXq3LWyhT0TXU/Dz
ZI2lOcl4ZotAv/htrCVsPfnFXxsv4gygkFkAmTKjczIBEy/UUoLVuPyH7fkg
4TvxEr6OIB4Vha4JA4p5/UtfmYXVYbU9+W7UgFlRxR5pNRJw7TcsN12aExnJ
YgJwa0jBVQzhQCyIWd2RBlkXOgpus6f/6FGei4ztOsZw1WSOABnIJwccieOh
2MLeH2YtMibJQqvJ2od2nEtHo3CB6L3As9O/v7drzAkxLW/E8uRgEfeQV+sN
ZrFuTU6/lJFr1PNo2BhE7fwjKYEkTIaGX/rb7FKrgAFmy7+g0sO177eU14OW
8db1dY5TDuNZFjdPZ9vyPN88y35ZRSeAqzz+Vi8vM8xRLSuKrefSVDogNRvm
WvnuRqHwlK+R/fhXDQuAJVFaO06NbUpZAK94yQz9vqYnuw/fXLzWtDVPxs7/
O187FE4rLZu+Y43/HpaByDUKq4vMVngxNsYInMfBPL3uACLhzFl6a6OkqmLH
wCmAllooLtyrFeiWc0/YYA0LlGRIL0pfuFI0YGYwVcWta7qQgXx0szjavays
HUMvVcJleCvwd/78mI+cM6gj78D5WQy+s7CnAU8CJW1c+dC7GFz7pB094A76
jm6qkeW08N8462WiYCyTxv4zCurqJF295V5hrRjcNqOE+s+2Pq1wopnA2EnC
K5AoPFAbVdZ3Ux0ZuvMcX8a2cuR2BacvY0E4/ndvnls87Nkhk4qiM9D8JUJP
7ZpQb5bkIhUVSwJhZeI1KuQBuVtBpcyod+aOrr77JklgC/nKOIVHSi8mWDlk
p7DjCNL2nqbNpxyHDVYL5gPHw8KnOvSA4sFuKhYz88lGkBHlwOzyPHdnXbZ9
ZgXPgk2gNtm4GXQlrPna+5Ckdfl3p23S2Vh485pUXVh8CCE4cMah1MzR6Cdl
GcrCd35a0MbjoDJcV5HqpesHF9KbVnUUaoBqsR5+bRqhfmBL5g6+c1Bn5E5t
oNon2fwjegPfW1ZEt9iNQmvO4ooNRlP/CsQ//ceZOltOnEXmtDEHAmyXYmY9
DEmKpP84KJK2S5KhnP6Qqwe4ZeUyby2GqpSmueyQOxizohYf3ZMj2XQ6syzH
gkooMIgtVGFajz5Bijee9FS6IsIkbJQJeIuJSYKwsN6jWd3+8/wXxVvvbH87
ZdYDdRJPCo4bAvhHO8ek3j0HekC/EVRvlHvZSWxhxHYkF6qWBbq8gh5ljXgt
l4nELm5X13nGqvNGotRZjB5Krkd/Pe+jrixMLQTaF0tWaLadeaWN6zDkfpW8
fdcNttK4lqIIZ/cdaZzSxl4WK9P1dckS9vBA9rI4V8FtUOBxFuSAFgtCqBno
RhV4EWYsxU1em8ajmc5rKMOnZzLcbzO1JyvJs7EcIsDOzI1ZCxKx7SRftFsO
UCUwU97X7DxECGfx1LDE6US2ahWQkYoEkw18pnVfG8EaDxrVhtJsfcVHBZNy
EaElyvP0xHupCSu9aLLzbgvQHJ3bPFAObF9sOy4nFZ9WpBtIvzWSXNtj8wG/
EDxiGrqdm7Lni7jKkQ9OOnrIXMFpgZhbMPtVaOsQV7ZbNN3Rh4rjn58kYPZ5
GSeARuwf9FLEZ7kQNgrtrCMNlQbCV2j8q4m25dHsjDeJ8VxvedF9AqyGIA4R
cjdUW5mXYPYH1fJ5VNfwthnpaxuAqyq0ETV36XWNkCulceQ+/ciVVMtAUdBZ
lJRNu7FG2znvrCM6/3wgt4nwZLqTZuw/oyl/8XVZcCEfl6J2LM1T+g1K8jBH
wG75XGCBtqG49DwK5IvdzPR5fnFWy/Vwv8ZjXiUIpq8pnb7zWjo3RnkHLjrm
1ABJ1jw/TQGJG0nL1BRQWd6KoCcWGVH24ETGu5q0Uf6VzXxkr4acgly/KSOo
nu/c/TneERO4FaU0iuuKbFjY3mEqZIfrfBTJJwpU+TztICRKOkyqS2txy40G
7ODlv9aLxhAGQpXCAgALZ3o7YzAXO9BTEDX26RzmogzfcRXC+uiyVmXKD4Ci
VVKsufWeV7sC1k2qGu+YRr8KC8zq56i6N56c/SD8UnZXtzkmcm5oQ1c6oDvF
itjnqFm07NVNoXbIu3do9X8uZaL3NRIF5daQNllvim4vnomjHlj20naZezPY
bEdHsjpjiT2xMe/atn+LDU0M5MkFAkEY8wh09gWfAOZQPGJaEu0zmQs54xux
TRhJ43yycz5KRXbG15EXfNXeqsVufwomjqXWnKch4iLLy706YBF/bQCwAdxT
z/wtiWWenl8bR5emtXQQRKUjdIkl/1TsKT/+kaKtoC1/9iiHGnv6N2uzMVGk
p/sDaduPQh9tyvkIssu7hcjL5zuDdu31LegFICMle1gMAxLxu7SXlWsQlEGs
vVJ5kkmvhIT+c+jFsCJK00/KxZl0INmQMaFvavtXvdTkaZ7pyy90DCgyj1/3
aAqiHz+o+KaQJh/nzTVGq8eCE3Z1ZLvphYvTL3PNwcDttveBHkyjkzXGzpxP
zBU+RSQhPNjlyyhBzF9Q3iQ8K5/o96TPjpdawhZPygKFDTzWPWHSWKSgNe48
ndzdEFIH11nbr/2/SLGVSq0+eJP5gcuYsTWE2j92pA6j3oEtR7/cU7ShqJGt
MdxLiO6lm9FWNunwIbU1quUReYZw86grUmntmc4xxU0aXTg2AXp0uVELn/hd
VswhTb5SgBAkocvlTK/rMp8HiKoCCdXHS+AoYLmEs8CHAax9O8ihpVHnqPBw
OgKHPHlbZw4YdCiZFVw2I6j+l7RTKFOuHwKm7OHmadDlZQyieSQBeRs2cnkM
Ti3ampDZklP/DA9uONXsYEYLQj6Yo9NlhPrrTiYu+uyDvWTlxDztSNOxMAyD
bZXROTij5tvezw3jlZk/nz81EbU+V34J/iVW81S7OjQBJR3phf26nygXQK2Z
4cfHhWtmlx9TkK2NrT3m+lJwYGrE+XOIiGo/cNy2ft03ww3vA7XX6ObEG8pW
/ME6aWTiMHo6/JYDv9OwtAI9+qx/lGfKPsvsucHavXJjzrxgu8n3rgmY67G+
NHFC1Eg+/3ghroKaUhWAHE2/b/GsGtqyCiIpNuarUP5jBBRqWOReVQx05VBL
YZE9YTODDuQ5JuORxST5vZSYMgMn2X51wqgdEnFjZo3Uelbsm5rRzV2Xpmv4
JB6W+s+rJFbUht7CKU7MbGKDlrZ/7IOu+tBtPmZGDM8kp5sR9rqnPaYHPfQR
NC6UuSmyAjOprehT6vBJphPFX7wRA/bh7nW61AAOwXJOIeM8CSyeOMFOBQGg
aNWZZx/X4RxFbpif+CzdCKIREhuhTaPbybG+Ctb8ENiHRJ9rbPE/8/4bls5y
HWoPdNCNFNhMuj+mL2189/4XQ4XlfjQj/GPVRKsynS5lT/iIy6jyrMWSdKm+
1XK0V12XGwQK9L4aqtGk6xKHl5PDnRc4U1pNRjIH0d7cOAFhohemxtKN+t4I
1KcV2jDsgyfQ1Bgh3rBQ7w7py2sEebtdTgl1cUvmdRxE3pC2ttEc1TKXUGNI
DEXP8DYg7QunGhvUKR6POdE7B3i0wnO5vbsuULP7BNJ8V/Dy8eNK/Txl/X6Z
+pmI1nXVrdkGQqvRKKdg9mkG1cOtqSJd/evhUmCEd9wlnMrGa4ycEJM5ZBN+
TtDZSOyB86Bh0Ip1QyZHUlfk9UD3B9Wwq/GhuqI7TC7U9NzdT4ddv0hjefG7
Zy9Pd1CrEuwvL9TuFqzel5wHrmYIKk/VqjbFZU0/Biv2UeoFW+eMpTkNy7wX
vRRvbNg4zCIb1Os5b3fU0oTFcLm9Yxka+995J0L5uo54/PJQHNmvejM36rwB
/X2wyH7wLTmeu0yBncpjJq2S0pNOVRhXZ472fflk7Xbv0E/RB4QwXDlBt+PN
rHp455pYE/Vgkz1XazDhq1dO7xgMSeZwVLuVPlOrfaSYOStFxeaGHei20Y/d
MsTkt1P+i3YYSn4jjN+ZAH46t9Lw9QQfamGGyHio7lhcQo2ZOvze4wbv7R6J
VBpUoztSVFrqZcWGfcF4PyVNhEAjcGRflsbk1I/AV2E9+qKjX33CRCWQ1gTd
fT7BtefCWLO7poTbV3JwE3IqEK6Ny0k4zwN3RdMqCDEWBmFi5d4X1LBkczP9
Pwj57hyT5olkDQAMg1yaS3ckcc+W0s46EQ22Ibhq/sPqmU97jaYtxBI+7rjD
BiuCzxl2+BlBKEY7DA7C00MlbxkgMTxoxlWpZMkho2eWaP1l2aegh+eg6a+E
0suZDJdpJSHdwIZ9T7fXN6fAL66/wCoiGk1IWTBSkRgSY6b0aYeLUvhnlSrk
+wEO6WcAkJn67LECIJjdoK/9ZqzOfBj/waXzBO3G7X3oopCJfYlOAabN5e6C
F4RA1xFMd9guTtnsqYSxEsJEy2eQ6J1BgTHN0t8S+VgJsiRmhOBdy7YxR8ww
n00i5+EUSDbuMnJwktQ5BuhCHJFYcGg3jqc24teiuaDWz/GGT7+9Yk/Gb6BM
LIKbdWEpCz6J3xV3DwxZPXlwB2ZWr4UQ3G2lojkU7PYB21Z00TfiQp0JBDIg
58wUbvenyKyQwCY+fhtUU1aQbddyzzYJABdtO5FYJGZPeN0f2hSttQEdP63Y
3jWv2bZjROx6Qc0ZCcPIaApPhBgR7zonGArvgr8uuhEYBBw317yzIcTS3Azr
risXUt9ODfV8wFCHHrZq1eljGEtmLzQsFroRi4EMTaD0bcRgZCz1IoumA6SG
BGU9M1sQpOurkACVlyWhZkim1NlTQTFRkQH0ynSDAEWH9JIPWtKzh/8BcpPG
ByFvfrT6hlUQmIcqvVEwigDuwpHlsK8wN67RZKGXp7DxiCfyLWsQzlB6AIq3
hKSLqTYdMGij03rx0YoOPWcCsdant/YF+sNuECTS+DmVzjwi8qlR54oICBL3
SJbWLPsQSwnFgvG5NJ9R3TsfdC1095087yPKnpwnUynisAmglFLfm72CoVpg
UbHVV4hbudaMIcECq8z4gHUuCkT7/1ahCXJGI5zr6EYH+iINaRSKzRd2Z60e
yoSNKku+TvFfDd5DbzmBUIpk8K10Ty044x/T/6M29687oY7zE7LrCKD6Nvic
XiLnN9uIW8M4/osSrTljHVSDAIN9CBecIOoI0agUgvXSZgknVc29LkPviZuL
nbQGMLoDWHcXPCvna2rMLsymN0yBONl4vWG0xtDgU3jcpYT9nvhA8cyaaHlX
xhMl+pxW4m2/6w5LvaEW6brZokgyRvl3aGu+Vs4WxjyXSePOPRBf29+sMnCu
U5mKfrWfqL6y6gvdGesqViN7BZxswodUH0paCmVvZq9vqSKI2rKtUaNcshVb
mFgMtAS1hScRz7KvuwuSEI5c5thQhWPC6F47KmHzfbbbvwDysGATKma49LV2
hKjQON/6uMy+ltQvde4RoiQk6Jd40ecf0j3gu7oPhGJ0CxQZILuwoIWQyEFY
DHVhFWsKF7WJPYMxMw8y1ew4jZV0CmYkiicbUJDmgICw7g7Rhl3hQUn5WJ0u
2wqqAXjTopHgnz/89LbtS3LNaHidLKv8igCVBjAhKsJau3peCtiwFXY+WwGn
Unm1iRJetBnDPNFM3Bx9oC2rcT0LBKYMe7VskNVqM0hFyVmhxuWnf6+Isnkj
f6LZ70nSaQ8PTP5ShiZrLTtXS/4fuWE4EBNpj77wr1MB8ZxFynPdHYk+8qBx
tGBCrRgxMm0dSA5MTk7T4uoxrh5uz1b9g8T1XSBRMtGowav4Bt6tsf1cNAS9
caiaGDS6CMwXo4JOD1CaZNT0WmaNosaaAWh5GMz8glxx2mzNsWWwY4qRq3JO
cWjlT/40hKSifPus2K4NcV4GdE9o2eqAmJTUCk189z97ycBXPw+O4CddGzVA
CfSLja6eYxPmm/NCY+GQJLByB687AhEzbqKvKWlmv1VvDp8jQNVfQ0h8oYOT
/dwYyDJFllY3lgGz878C26mgvoImGW5bZll89wsu4fjRnJjvDQghHVv28zlL
5IGyDHQTde+8Aptws1Za4T+pFlfGS6xOhPNzEI16TK05TuQuQkQtA9TX4V0v
i6CuoEa3qx7C2VGi9cdoAAKMRbcS5rhR04e14XQoB5cmRPgeVMz7H3lIoQWc
7s9WPt/B0+VNbpQsKbiXhnBxXnxuHnBiektWbLWTKcwPn31iio/TEyrwbG9n
/HSuV1TfXjZoxSS/IcaZnCPByIzZzy31lOw67sD6rYebBaa+7sEsRz5OEBDm
gaeDnpatJO1sfBdW5KeBQxbj2BcIYmXt0vuSBf2o6M8/T1NVLwxVY0O2/Lj0
MK4gsT4yZ4sfkhSApeyJhi53FHSO5oapqAST5rhYfvrqKYjS3qVEjlB6oi0r
lHAfJ6gkjtyt4/TYhA4SEbQdNrqVD0if/oKH+JZXoV5ByBBqkMdlZS9pwe6x
xbnJkb3X/ib7s14t+nVaRXzDQJrRVDwrGnOHogFgeBLgRmG7GG+E9gV6ztwj
xbiq1zbD3ck+QxLxqzcULPlyEEQrlA4MG/GpW2T9xGiu7fk21EycPxEWDK/b
hZEZfTDaLY8s6lHZOwwrEICJJgo9nZ0FS7TOhPLQGS6dGTrs50+VOaAfch+a
3rZTvLU+NuetALm287k/u05zpQOyI6/41Iqu6vEGMJp7VyrBGKcTfORULizw
kyt827DfkX7ggnm6tiN3PG8rGqfjmyQuM4YQ6n6dcl2xNawr0Ffg/ii/oLbG
zI2RQMenjH7OQbyX1x9IFyzBgg6htpYlFCbK94JTojyMFzVeVru7sH1/+oOW
Qb0wFyeEBSjlBk1TpOmSI4hp+YfUW/0SzjXNpdlB+wIleYGrEw3uaCVl8vEe
5nJ5yoDT1RAN0saT/4lP6jVI9zA1uESHJRdtS6te2+GJGbI0XPoyz2X1mCgO
0Ym40iM1k1pk+QiOiOqUzvmxVkcZ+hUs0YQNopncyHazh/v4o1eaFrHYTakB
o6Db4+hUZnrLTE8E7sJDeEG66PU2kPj0j/8xA4B7KnnCSnU1vPxRxvW32XGl
Ei4iFMm4abCRFWJAHpqQVCHeKcvgalL0AweQlAQ5rAZKxq6HLJVFygyXVsGn
GMLwJrz+jkQ8L7IplMZwDS4/7js+MN2vrWWMBlFARDGmPsz//+9dNFsQ8zJp
MetsGZ5d5APiSgNjOpAq2Z1wY8n79mUY9GCIB9TvPZmM3XEJ2XmedeaO/viU
pWJgb5j09wkNzYCog4T0BSwPiAn0KyqqGbb76HqSmFL+/dH0wr0ZC524Ty4Q
oepLNsdaG0o77V4t4Me/XFxmRxbINndeojA56vFIcHQq2lb3MpD0D3VtnrXZ
8ezuDLfowOQ8n3ZCOFdqnjg49XjQOz9wBaek+voJpr9nqJvGqWiw7xMQpWMw
NL/4PkEUzijtdTFHGRzoS3hSMcHD5yytdSxqlxOKtFfoTDyBdd7IbUn4wfYy
fT2F9qcOHHcCwdIpTtg/Nu1yIwBv5zwbfP1tWvgb+2vhuHkNIi+O0iUGI6+R
3ddnlYkEODWBc7lEIZ2b6+fO0gmRF/I95bmJ3I98+/ckUhB0Z+Xv5WlD9yPb
2Xrwu1dQb7BCvTgg6H7gON/1n0HvHp9UVw+FIJ/YU4YPgeqCQZ99HVVJp1kE
PVnZUCtw0BV8X2tUJhlq/oZhbKUqn05ZB9a28GU4KVo/kbnHKbxh4abISKzb
l3xopz8YI18DlIjtPA/4tiw4g9IpBjC3DLnjRwvVhWOEMg4znAv18Gixn09I
PdPX1nEk+acAOuF8y8hUGo5BEjqFTgiQuT6CSRcBQOC9uuXidxUAXegNeQEa
4hH2SW0Hv10VCgMWj9PmKUuSQheZMnPz4SCFtrejGxKpoEcSrbAc9yYuIYu8
v5ruTIwnuItd1AdULmUZcKi6HGy0YdVMTo/UYcGw4aqUQNRgnZXNlKuP+Tnm
ODLzaYOV0KikfnnivW5oOmnEDtdCm39xV+bXHMMykpCFUNVCkaXAtbKdg2WW
W0//0UY5m1kaa9UAQVr2Sc1YcXAz3ZfTmiHmI6GIqI9p1iOpB/52H5VrlkB+
mkB6OQYzqEX7pIE3RSRFZtkG3587RNdUim3LddDftRmnheVYJ+D2lgi2NXN0
VbK9sGDuveUryuD6aZkX/rWBRKRYKT8KLETGbx3p/HN6FdwQrHupComDzia5
geuB4sEUzmqV7AB0tlRvv5hKMp8ST+JfrD8ETMlI7BGezoknUj4cJEFzRoR4
d1NmmwfvZS9pY8u9XnLAsZmYfR9tRTTJ0fkSaDE8NqDlDoyWpAURxBKjxqd2
bGTh0lhkRr4uAr8tu7MYw7UXCPRG16knMO37pTAk7DRmMDYAoTXDYEzavTHP
Uxc9GGINnZFGbpSS/2GYCJ1My/4iawP07DNN+/jl5bZ1aq+UdraYqOWuIE6W
hkDQAEGuO81nnpeDhJIudoEzzJyxEZkknzYFReBag6KYtgIOjYKGzvqTm3ka
UA9KBwRBOx02sskKfMQJDSViGx+4Qg7ScEWxo18644rCM15gGwR8WeBubk5f
v4D+SBP4bFsXcs7ObIvFNHAqSVNiQajcvpmZGv0rI6OQZNWDIz2zYvNbRG88
wbj2l3wHgZnjl8qDA7mddZnLIkuRADDb+gBmaubGHfIZaSg2FGIddeX3/U2S
a2fFOScmNs2BOWllEyWf0ONS7X46Hyj9iSBv0IrcjP8ShDbVvfsLFIVDj8oX
1+jUcZJe/4aLOfgz6oTpRp6SRHvj45XAuIi2h1/e7zTAFpNd+ZikvtjU5jrq
entsmUeLL8k8F/Lad9L2cG64x3z3QhKq8XYtXBbmB6E+4Gh21/QGUA00B5oN
qYJ8qoLDVpEVyyg4nvxdldJ2VWDSAqjIpndqQoUWIsCcPb50h7n+W2wwiK28
KTsMnvQc5KRQ3VMNc/zw8zBOlEtGNu1sJNExLlftA7rl6/7c8unoZMujq+9S
8pRJxcI8yQw+7Z8DSQfHaskogpOp26FcpviL4HCZW52BvCwmgJ1puyMarIzz
KemnRUIj63nr1IxTYvBQ6vV1u1U2wDEVbBKk1RN5DVHtR6JnYpQ+jhTAfKzH
0IXp4hNw06JurcZ6Tj8qJqurbEXmYzrtULCDKcuXk++vyuUzz5zOmYuHoItC
dWanBjGSYuYicdsueMSRBOOAHlSK0gNZFn2d+70cPj5T8gncGJYCFbLKSFHn
pMUqhDPt9/kVUVi9Y0JuV1dMR8mMcol4BR7EbPch6DVz9rxdOv5fBKN6WrUi
ZQYYra6cYWTgQimiD9y0dwBsfecgm6grIkfEjf5tuOkWjFlNxTRBE+twCiRV
/xR1V36QijC51QlQPri5GWDSGoZlIzJHW5Yze6FCKpCJ9VtuF97OS/hOVe5S
yhwgfNzHgzJTsnFexLvO3dRpUsdRnRrBSsw+h1HXm6XFAIpPeN0+GD9Qb7++
OhMvOnk+FVMcK2TCzt5VMtmTJR+v+XArt6ydTsiZdfcHfVAhjyeXTTcditqz
PHdOK6jih9y6WNX5QKZBdCPMH1LvOu6uiEzMarSxsqrwxhUeemv/sZbYRs3R
VCBkWyduDbAY2Rof2jQGcEnPaPyu/A64U0AyweW8sl9b/J4mpapHY0SEawk9
sOPO0GpA0IoMj5tWfNYhiOhcNEVJNGwj2/qzhhkxZ6QWZlk79roxv87bl9db
qxz+dAf27T+Er+Qj/Y2ovjdu+9/5tiGEbVL7SxRF3mjtZojIzazrwq4Nw28U
o53IK/+a+vQFGGLO8WOSjDlZrK5czN8ifzUAfuxWZKdgZvEsKvz0bwTcPaCq
W4fZrUnvGj90xmlReO2G79LRZDzhskZ3tLOyOdImoAEETOlHhJ0/vlXn283G
8BvJuK7WpzH4KiPT1RdrIgRK8Eu86TF+GMxeqAiLJf9B/riwCfY8RNlh+003
eCcDOM2AQeF30KjhadaL9w7yyrKXUfW6k2V2R67Xaqi8rsU9SGySVS4PavnZ
+vcaOgPvYDQhbxYh4yQWLpVvkAdtn/sEd0rNPQ52CGcz3K1RMjAMH0Rwsatt
kfSZ5J1FxeIlRf7YprsG1I+0HchF6HWE86ekSMyOaexc9bQ79OZHboIxWqc9
4n/QnIUorCco8OqEwrsdhuZYjPcWvAjdv/urmP130m+h5qqx8AbMva7GiZh/
LBatGZQmYhJXRBen9HxDbByPkaN49USVv5WrD8seSlTIsl2QccOKTAG22Dvh
XdvZBxafk6wB2p2WNaYN8D2BO0SqeXQOWzZq6kE4KMd32O/J4xLHOcVmFD/X
2Ku3HhIIqs7LOgGSZARprJwS8hO/3T4tupbWV72ke3yGaMFgagFsRd3KW2cV
jiZ3OIysQkdleqb7TNOUtwLpVXRzaupLdkq5C3T1iQYknb9Lqay2QZu/a2ub
ZtW3koL36LW3R68JXbXXyCU+u8JsE+/L3mQ3diauwHMvu0ohzNQPmvrpyjxN
j/ISSXQE5xKY1MnPIpcveqtpGtc+UUKfC5dN8p4yEb4qVvpOXqS5tiAyRoOI
cIAw09pbWvxOT6mj4Blgc6Jz57yKewIEKOmNxQiAmcOizJ4WnxvEgfj6bVPT
EVJ+1ZxSdbfehtWgc3Y9pqnoINfGCzZxXFl+xth4aZwXonyZzAo2lVQknfGM
fxXmS3riwALm+y3tQrRrIeATJqD5e6wfL5sTxQ66st3wv1XnJ14waWweaaau
xI4Ep/romgTTm7fadTx6cOxV06eYcYcQ0gPRk5bpS58OZhv4lbFBPe0N58qI
4R9JYSmo2oSW/aT4t/+yBAE18WkwjwYvQzfcYMoiixS2p8gfoTagcO/fWjW+
aOanWAXQJkGZfpxv7XaNxMO8o00meyyBeMmCVdrCj1LYbHtWX84XpeDSn+cy
46WWDg5jBRMPbEZcAG6YW0mbfdsTR5ZO13O6qRoH2F5f1I99wdKS6t95ar5O
SX0LuK+O35yH5AvC/8/ElKGr3Mr+8C0vohihYu6S/vxhDTKqfwKkp6H5vxmd
lPTiUoVUB9vJ3wUmRC9xv+bWU6UJib+3cjQuCfbrI/BbeC+AruqHf9S+4byk
1use99lFOyqeBMtKSbTbeydZ96DqQljoOZWbOFiTNU+1GsNC6FRWHlCXl58v
Gs4rcpEcAj2+TdDbBhpqBzoqPUWWZb6GTALpqpUwXQQNA1JdE6BLWk8IkbOD
hd+FV3TQpBJR3kJSaQ/iDsuoPWUXgLPVKEWhxfQlxYBmLiijd6eQSf0PmnLj
OlJcB5VrFj6X84FaBC6r0gKjWZyWhgwgjhLkaMgxfpmc/rnV70uLfMagKGQZ
HbWV0X6F4O05qXk3Se6YzsaU7OVHlbRurX/Sll5EVAsn08H5RMv/EUgeEuUV
26dPnN0DAtbYQDhohotBpPUqvUlFzrhuusrjDm6zdCfOT7q5Qnt7rISpc98l
7zDYMx2iiK1xpLS9iCtaAxX4Q0kh0Nm5KSr69YsntN+hB3t+Bk3eMllni40G
WP+EJDL3+98yw9F7il1uC9jLOu79jpfwl5+gGdmQVQh5JKuGdGL/gyNxgTMJ
dJqEkg10kN6vhro+nLX5yCYzvd96I941RjJka8w98esDIAAY8C7T2BVqZuot
CFoVd+045OBRFpz9jvCuv9REWtxO738pU7XvPagByUT5Bap6dCu8efUZz/2Q
QPQHjHjIVeQB6pMcf0uEpwur/E3eh08JDDJWiWWvX/UDzDXcC6VzzbIzvawH
Xuwc89c0UlGDn91AFPL5mM56NRIdtxBh0tLPkmNR/F3A6/sXFLgs+nCshVac
NXYZWE3qplnlRaXVFWgM4B9PbAHgAfyUUYI6XSPQiuPN7AZRImxJTcc8uXYh
FU2B3PL/vBQTbPXJVbAiq17VSLdhSKbIe9L4ZdXm2eiHsgMQWom2OFsp38Gg
pC8g5lokQOmB9nxlLfLZrwu34q6r1hwYEI9kWVegGfCICB3gPyI80yULGX4f
OyRFRkOQ6MDp3Eq7OELarxwuaJ4JRqELFmCZTEmE2JAc983jkTGSvQdZovnJ
Bon3KjP+AOIVCzbD4JT2LNnAvSxLg9ewilm890Elhg5/k4cNBmQy5EBnTChx
+KhHh94nPCR0q9F3dCLkrUWJ/3d5Zf7WeP+E76nJd3g16ocLzZZJYW+i5c31
fz6Fy+nYFPo7qmbtAna6GO33Jp9Qo2mhJ8XDoDKqqN0YOsa8W7P5AEmH89PY
WKbsc4h0YMMzbCTgKXBMCTqovtPc10BazIWpsTf0vgB33SbaGSq3ET4yCl3D
gMTsZ3dI6uQceSohR3KYMBMpYjc0bTifl6hP7LiR2dyYzqo4nvorS16fGhW0
FCiiyrUcbnKi5Cer1Jc7WrN6vqETGA7begxJ4ztbp4wzfnW1/gYpHCXHF+PG
C285uk/JlYebjxiDu7TBYYDtv4MHC7Wss/IpGK5CN8iB6PExgFJOKiyg5Bwf
jqjpmRpQ0wKoobEh0I3LbIIQ+8uwHHLATe0BbnGS/zgb6IePxpRqXh4mo6mr
tCSLIlrLD7nu3G8/baLR6K8L2Gw0v7aEuWxx39f3wVBts+/UlhY92hlQlUGy
QE+R5fWva2mGhT2Yc9HP0Ltkesw0x9CKpvZAsN9asSabIYLPRgapdXReYcfI
dBvju5y4ZNPfJDVki2XpmzCPRefz04F+TTzazaiU8FwyyXYl1tsz986/dDat
HrA7fH+o+bDzgep6iwhO1Nt2XcBIu1oIOF4CfdY41wSKd9uDzHmMkUn8+S0z
D6D91kqcPF8/IAyaFdRqHnbbmXCqgap9hh2VrJtkFLJGTB6w5JTejKvhd5gS
VLTXntiJt6R9uGApz2cF1NX2LoCKbuoImdAfW+PQLcY3amJgCM1tsJS/a0xl
+wK3yI3duye4r5ZHPyFeuSwyFEOiAz/7peNHi0YfKQZIJiobVpzDaO2kzMqU
8aSscb5XRnmUyHfDhbYlu3T1g9S+S6DZS+X/Xa5dYTeZl+61Th2ZjHKLQB8C
zlArhFOtz0xBw2pUHdSxIiNF39o3KV+8D7KpkzjCLWqycCl/0cCG3ZxZxezt
n+FxJBeoGvzbTodjFQzCDbGTnYn5et56lPcb5uW1tTmdikKfJpdyURe9bPZ2
QP/++xMQoahdpnayTS2w0U+w4hmBirPq7Nl+irR5jFPiIbzEDxd0PZtNoWz0
OAzKQhYyAkvWYzNgI6mRwO4ea3Yb466q+Ug7ZtbzrRaQ/oogrgQ6lsJ8fgx3
pduB/7cuEYfM1Rw3wgro3OCBBBGKFvG0o9GLTGWLtwEBRUH7qCMA09k8SMFo
g5zESVBOjg4NW7W64NmNyixUIa+Cq8DoyJePx6smqeZeWKayjphjWw06uKnC
bOTZmDWFfli2opG9aCk4eF2FBo+8xTIYWFetVbLX1ESEFnnAFjHfBgcHUUPj
QmQBx7CdSYw4k+lUR2ERBjbB31WD4X9JNY6LKvXO23WXCsP8U4n69Ygd5SDJ
rSr/If5X3EOIyIG4Axtziiz1EBeGk6kcn583IGC67dg2EsFR40rVZ8NlOjWs
nNeofYTmnJbkdn8Eoy/ZsoeyqK6mMQ+eILavjZiPS8NPtpr04CgNTwTTI9YL
cBFIKHcGANTo9Q5mVzPI1IXpEZ4SOZAM8GBYJSyoGZ+Ixdrqogj41phMlPCG
wVNiIYKXq8Wdz1y3Dv3Cv1k0g7n1uJhv131cHeSs6sAhwTX2bt2MVEPDWYi5
yHAk1TmIafhE5FpX7RhKAVEBITBo7NcFAYJpQvfsva3HS8OaEMKX/jb70uFc
uEaH+s9vrWlacW/y66DEIGhUIxTg2J8C+c24MFstEz5tLUbqw5CANopUOUFz
N9zAgNCKxF6MtP26eV8TEj+L0BvhW3TTyJXFtgbmILiDNNU8vQtv+POzBaDa
omPTjF5c4kWNIFf4+rsSfW0oLLm64nzqEyD6zuAZXksop4QjYfidFp8vmkPP
9VwGAAzbnhfOW0DEvRAnsBThX18VQwiLZwWq6zBnmDfs4/b+tScvOZE2u5y2
9szmF9a0JcmymYdKg3qxl2qb5ighLjN0ufHKhzjZ93/Y8APing5CSsGR31ZH
naNinXcsZvIG0697JnFhebRCEZpEdDptJAZkITn+F4ntR6dCsW57XxCVYe0a
sWO+Skn0qjv2kby70h3cjy05L6i+rx7HQXbdH24P7HaQwDnWTjtlkxLDBeD/
d3FF9rp10v5invhRQ+0hn9XvccFP2WkMu38HVDOc5SwMwQkr0dknxnLlmImU
m7yp7rJECRZarejFZiuBTTzWV286eWesNBPUnggijAD5OWcTi425JOsw26ab
AgaWGXlGn0GsN34Wdi9yKWMmegD9WwWfirYcj7j/rOZJaRdv6VcjjU6a5Pbt
Ghl48+bd/OsdrqVztgaflZjugMZUvmLcrm0NteHR2rsVzMRhsUCJMBRR+Ncm
SyoJFyJW2qDyC5DQlHGY/C/o7ZXnKEoswJaq/mnhE5+xffcePCUDLcbJimDb
WjfzqHI/IZV08opyEQTErw6t7NWr2zBkV2R1xLPOcQEP2YarOXu6Acdz/D05
CfSTf5jyegjfo8FmxUnE9iEEuBpFVXoVosiYfImkp9IdRZtQpndaXiaSYsgv
oIyGZFNiBcplX0jxXRSg577/njQoauxk2SmNgtvQh1yic+kTg5ieDSTfDuC4
6M0YlG5MCwtXwm1m5vxjYs1eTrHJskxSya5zp5K8j4UVmaDxxQbk6KKA0IuT
WytqcC9mxgOeoCc6niein4qtAbgIOOO3RLq5YGdTZYkb4uNTANMr1vH0qHLy
0KMI9gLkrryqRz9Oeax8H/n/zkVy+62CJA/tYG+VYFPbl+CEtk61VrgmpcZL
Ux3Wn7xnjNCtgcLmZP+Rcvd+Yr4yGa1Lpqh3u49mnZ6/d6o+S8d4zexmR4ag
iaR0hoOLWy4sP3S2pZ6eNnFyjtwXSxcuISgVA+yaTUBlQZ2SOcuvRaNU0nC9
gOzxU6B8r57+3sp9GwqVu3Vvlxh3kdCZWOTlnaFtIYb70aWPdQCsb1prlrs5
M5Yh0TG1WVGVlx223ijSDa5d3V5MB9s17kPYw+jUx745lFtT32a01epYZYCW
XiYvNn9ztCVpphGUyStcqfgj6sEbV8P3zDbSVfklIXY03Nkv5Q7+qbgpnF92
S0JeNtQDQVdfeljZl58sh/X4Zqf1VgB8K98twnGQ79fx5ZfgKlT+4gBRPBtV
crcJFozCAogCuZIqBK+anYFSUDUvn7J/d46ku134qQ9n/c41kSYYJ8mWFCmq
iHU1JxDGxyM3OSbKOfKczh3fRL+femsIot86QODOVQS1Y9FFobw30ikyMhxt
LxLz4A0UZIvRhGUiDSRd3KY/GX/p/7EoZXMUsCMe6+ntpGZ3L+7Rwg0xvZdg
uA775YYTXOH6Ly1tu8O27d9ELb+hSWsmyUt8agTBhlynC5XfQXJmuyXKnYIY
ar7U31JwbHrMZo0HKAqBKnNcz0gHb+00/UDecSJ3ES70s80N70FXnhUpAa8i
Eb/b1AT5iJQn3PfHpXBmkBrmGrr0cVySa7+QHpbCIlCQTHYII7AzrLceswxL
yE6A/LTILJYDuwj1GEZWX/vIiHt9N+r2VWEsc1quo+G2OxAwK3RH0DY9+Bcn
LA9faJbMafMji7INr1BFZupjy0SvInii4XS54Pc0xCbmOy0RXaQtbfjIteH0
iGvzw6+ONR0HVbJ8gaXpmEOAuo7+aXaRLtmDh5N8ZAkKCl5FbyNyNOA+d1Ru
d8+F4ILKjRz45GfYnFRETVK196/tfupI/wG2EjGR0aAE4YdBmkpH3w8ZzGXM
ebuAjmDnHtRuZEWhxbL7pz1QQI+baeolGmUNPxbdtwCjtb7pGuKxKUpfplp0
shA+QQZCYYcUQ2WDLdmQn9fasUJ7N9d1wxt5pFZMgRE+eUwZxHx/pQ3ypMMu
OOt7rEJzNBaTIHwdr3PnWBcyo8vXGmQIIOKXThiiCLGw4JIl5RG+q7xgssiB
ZzklXNZm93ZabS60jzeWyEGc1SCKBXtGN4S46lXXWJAMElyKUPjcJR3IHcba
13Dtui0ixiNOX3T7vTq2kXPFahEsARELu6PxNHl8JJ9YLjkbDqLqRnvOhfTG
cBIn4lwEEPy2twdCYHNVoQPxXhoVTNqSAxoED3ATnPxUXn7CMP4RUYOYNrnH
xh221UTWjI6JaJEK+nNcha4VJIu+mhruG7dqre5Lmc+OPqkcvwhvzL50gtH7
OHqe/cXY8fYrjsR3lx6jsV4zcJ/EayP0u8iCwGJHCSlvy3dO5VicVGgy6mfV
N2RnTDIDIx2HIQO6cLof4/WMkapxjCReF8YiCzk3RQ2bhCY0QnXFwtrzS2U9
F0F8Cc1S4TuZLPmo8AeLWS2IV+rwu8TN37uq+KKk2m9FW/Xt8x+OB/LHMCZS
G5qsyX0RaUvB3snPQdRuJ9Anrp8Y5QOvWho/0px27uYESJkGMyyv1tN0dR8L
jRGNOIUWi/xqIUHoWxIcsWlyRAWu/qu60asxyCF7QYaiGv8vW9C/hmMxn5r1
NMzpxZbFP1eEklMh0PP3bpKh85uMmrqYEBOs47iL3fq0FrnwsiPbBmBvCZsX
Q4NQ3D+lFJ34iSJazJaWMXbpdhjKV1mIb5xEEjMvcvD1vUTgweaWB71e0YOh
KV88IReymIBvzbn3J2GMc0K1sxU6p84HSn6AbXwSuS/Go9nlWLrsnjvR9kLO
P1hAtQGJeksgceYokNL3lBmlLZgpyf2tUpxSfULHO6dDxRFJmTEgXW1lpkaa
FXA6ySdlx01Etp97FXybbBT9xUyc3VhmGaPufCl1E5o7IYrNqfsaFM8amD5x
nzf2jzmmuVtGTdVr7YUlDEG82hKW/VKhA/t53y6pg+io5XODwLK+LLF1yIhb
eoMX1kd5upfl624q1MIusXUV5X1pzuonFM9oPGv3evUGvXP60RrrsSHK370R
EiXS+VOtTDjP6U/qnDvsvE2PElhj9kXDwrs4t17ZSjuoak793LDNPR69h7RR
3Llb9VuVWXIRuGMEHvb0A3z963SkBRdHKZyFKqPCVe6dC4EPe7FdFV5J3Onm
JgK/VDbmNy4xmGklGOia8cLUytamMHGMm2iPOPkYxU7h8BjOpO3/StENpMiC
yyHa4nDLx0T1bcU7fpqMRWalvyDQaWFDvfe5gCq8S9KNiKHL9K+SUccE3qJo
GGY6hfasJk4Z4eq7UIiwYp2KEkxVQ6cfrNtPMHYMjyXtagYk2mNk+8TboUKH
9L/IvUlN58BCSVx2+6k9sl413bqe2HOZqI5BqjbxcPqgBZHrJ0HMq0Q3/Wao
0SqLJrPEnRI5fxBdyRpACnQxuYwX1xBwACfV1oUF5/crPunR08/D/BUdaBRr
GKCyxElGisXcM/rlKmt2hf/aS8NDUwh/BuenHRsWPKYpO+WGSVMR4SQYl7yF
CwUdZr9xNulOgpnTijUzNmbsdea6SVye2ZmYwlwr257m0GcGDRu6HNUi1iQK
kr8zlUaLdM8xv9rAz6EAKcpy4ctXIWj43Pp1vVbIekzD+zI0JeqPzl25gS6s
AtT9A3MevJMc6PcHV6BZwwAF4rGcUeDQRDnZ2oG8C9abtzXNAOpcYWdGXYeX
MhmH4bp+zEAN90lv6chp1VikyAnJjrV2AL11y7Kr63UFscy3kOg0b4NT+V6t
QmI0+qr36H43DkVcIg8tnJ5EJLv5vm0DMfT0V3pP8bb52/L3XXpMQbuooIt8
vXtwC3HXdb8dglRJIyuCCCy5VH/XuCOmc1apPcq2zMMnEwFhXd0k+9kp/nvW
H/TMADaoCuKIOuvhM3kcX2qx94yX1nn+0u73GsiXAeKn8NV1/hNz5vv7B3o6
qcMswX4V/0Ahan0IkI/wBUEfNDPS2g0WADTLnK162XbpcfbgcQUo+xDD7LdP
I/E434nJrNkBX3iY83FRqRb9jDVLmVmU4d2Cce0654qzuUX6i22JG6skLZ7W
BF6ejuOqyBSZz1hG9FXZCSJzfjb3zELfRsEjG7OQcz+mIFMsgQGgLSColXQk
kAGjOomKUfKrT21y3pZcnS3ecwQ483opBKigr3M0DthtV0Aeaq+oN/6dECdb
zYCLEZ3ahWWy8EaOAqGhX4N3bTIq/D+KRK7/55PqYYVqU1UiWG8mh0oF8WN5
SdBYajgPsayI3O+knG2DS3QlNjgxn2SOJg4Fn5XRfF9PQkmstJD4ULB/Vhzg
7nx225fJiSiCKnp2szowunrAnm/snAhhdd1GjbD3smmNnckqq80+Z4LmbBK2
SB1V5Keo57rVwOjY+7e/Q8N7nMr2O80tTRBar9eHWotnay8ONr6iWDpMIy2L
yQfY/cs0wod7bYHs3jEwBaXCeGjqr3HYaTnlpLWrIfsvG59fv7DscK2YVQbA
WxKbgN6LRU5JkFycuuiLI18invhgZARIg4cdylQfu8QX7l1FlnrHLtp6gc0Z
FdfXV+UClRUTwooIXKrfIo0IvmxFcoH0/IRCfQe4PMWW+jGNikzVXg6pqNSt
5zxY5y7oeMkTjWIMvOwUhETrOhb0zcfeU+e5tjAWW5GN4emBzRPqA7zpccEe
/v8sHXd7FlexuP2CqBVeilVGtz/am+els/3X0hKzDiC4IM0cxamL7NaE9x8w
DfSB9gx4UPPOeO+47xKqKQUc6uuMCXvFsVj6WhRt5DAhgvH2UUkYP1WqpIhM
Bt3vZbavVpUfw7pCoRIdXijR9SU6iIVS3dmVBDVv0Jq3AQuo+lruHsdDYI4C
tUXtt+V9dhImIZ8bNY7StQByAm3Z4l2b+djaZnw/lgp12rEN+IdSe2uZ/v0q
nPk443W4SZfZDqvz1bBWXKlSDbELH9rhvop9bcky4S32woe20vd7oTVDEw3V
cw4vJUZv5paveIjtjuwc20AC5mvHKUvwmSboWbt3fMeq02sG2moCdk4ej8Fp
Frwg2Jmk3jp7r9DVZQckvo78mtXHtIaU3y2So4ahpD4cq+W0WDdd4PjfNWBp
hlGPrR8nfhNkO1dwyW+x8jBBsLVmTVMr4rZ/RC+0wlXHhqifP7D9gCiRccn4
wGYG9RoE8iLBv3q29ZD/jl4bCUWQbZ9yI2iZ4M7uU1/xZIgQAEz0X8iAWJyM
DV062wygfVbO8raZQmxEKRW80PY7ZUp8Dd3RzT1xhkrPTM5Z9lkyBuZNmr4L
IBloqoaGd76gy6TJuEXVat8sZ+amTs7SgZfEwRDb9EBg08MbpbFvTAs6rzSZ
PQJLJg/Fn5T+3pCYJ3y/zX2iBJGrW5sao/5p67uAh4x6FjV1m7y3LlpIns3t
kNQukFdScOf+k53zW3Z/sGEYeWYFXPHXQB24jpXBd5hDWQr2NEKSn6RtHNlR
7lWGcZSz6xWd5XpWVZgKdyJ48hjZul0sgFvmb+4ef2/XKyJ7hHuxMC36r/b7
CDEF7htIycjxS94XaGoh0QSasWeqc/dr/Dy2ZualsbFn/5Huy0X/ZqDz4R0+
sTFSLTRwKpc1RPxtP5bHuBLliiX5mg+lcaGVL7IlJLPHaGhHOamz0TbLKbee
F2Ilr1F7IifQeE3QpMnJH2y/qXJgpMtR6giGtTZQZauxiL9W6/lHAc0HD9Y+
o1MRunZXfhgGYvnz7gcsoo5flsTYUc26mad7nvAPEaw2A3dxTCRCkhck9R4m
/tS0fyd9xyH2NSDg7Y6tfJdGIFqLFsV39RUi4nDJNI9NF34infk1hOIFIwfo
e6RmTpYJrBZvVjwkl0nJGCeKAnbj0EZoLRRUBjKL/nv0SwkE329pMmb4HGjm
FpYUOV8oIqsqdIYu6NyqYaLSB0uxUBWFWP/QL1DwKO37dbuUy6yMK8KKsLLZ
AoXWZxSSivsqziRh5X+W4V82aZE9e73iu/AuZ00aRUIvi8PkH0+dFfYw0kwV
Yk6SXpJsZTpov2GHfKIl+Ejo3A/YZ5l6e9aBpYXGAedx3BzsVZs2wZgaQqxY
ccCmAo8QLeh8wMCVTG2OxMaEyvDtvGeyauFy6Twun6DrH4qCll7ImWKegL8x
N264IjwpRcMDz9BJHbBaphekM/PRans4fqQgnBfWNqZYwXVCh25hpjL/hXC/
1zNlPNAhqkx2fi2INqLEi5CoYlWPTDO6UjvKBnz7W+vkNpaHu6ZX0cAa5xTX
sEXcWqGPDTlss2riZOl7Q/6vLtebO9nNGLTq9QjBE2PNXq6HhMM3/0A5Fd6G
tuSMAwXC/YHVDLCiOitMpn2NAzAuMvmbYDlFjwa8KdxFrP3lvyEIrLYPDyZi
qMno7LyJLDYhxrzC0HYj0GRPFD9If7/TVNO1giumF9mtM8x0E0hqx/8Gq0HE
vwMa4zKgWzgSc09qXRM4uwhxP7N906MEYbk8tgBQ6kC2drYHeNXvf9xaQ9Vu
agsFfesmZW8soryrSeIStAMMpxmQXdWA9P/B4KFmkRgdExMcYFwQlGmjREaE
Ong/E6Oo7vf4xD2o9ZmXGjQxRFy4H7I/ARb/0QwU+VNYOGvA/wkQzV6M2+9h
D9rHa7sW74itNr3sxlIpgtOJ+2NLZg0w9jU43ecfZ6McaOEp9l8Rm/ulsPJv
bPfmHdbpSe8qwGSqGp6/bMOs/YFHCt4gvJlGKM3WGAPU8lSPitMbo5NKpNNl
iiOlmp2d6zjhwhx/babxS6++azN1NMu4oRd6U2VKwSydJ5CknuZOy6bRF5yq
ZNwck0B+Si94V/9Tug5f42FL4O4b6EAy8f3jLx1lqwXg6jgOlv+IWP7bGJyR
dysSpM9METF9c0ATlqz1Uy68kQ0ErqD6hyfpirHIgIA7wuFdKtjBPEY3vVQk
aGB5FBCwFsJgvpVa7XWiKBFIxTDt9LZuMY63TZOeu3ex6zI5opU9raBiJdrk
uLr8I6KvmIpXCJvbdvpivNIDhQPv2WBMQpukLffLfvmCzbzcwEcS2jC8ic+e
D0FFP8IozeIos/5gTO24iAyfDo2bl6l06lSbQnZ7Mm8rYwI2PLKtpSoJHpoB
QaNq+eFomrxvZqjAOksO7LTOX5D9eCuPbqbpfIWb48opKKbv4fVn0nbVxZZy
OUOwiRmYkxSkiWSKOeBnahzNqWdpDeKAZBk4yn3xblG9JEtrv0jOOead0yxC
jRNauJa2mqs7Q9ql+Fd1pqKbyfY9nOyTGHUdUimIND0UE7qUV4gwK5j/wgJh
aUMkg5MjPp5UXz1IMDWi9SSkuBr4qgWv5egAQvWpAjfp3gI18tQ/LYw3sJRa
ju6mWMqMaBZJL+DFsBjik4xpXAmtqtGqlfQ4mYSuX1GYRcIOaeWF8CTjGVL7
HSMuNStf9SwIUbIJ8NvSkIvkJQj8Xe//8q43YT8427D6h2lrSraUNeDHK+e2
n4p0+e5Pq3dJ1GVs+195+o3MYrQTUXNVOpH+IoUo14LZ30QLsVcVAsMKXv0o
JPyMPcmVklFJdLJxxYzQubEgfazzQnDOGJBEefbzBTI9j9zEo8v6vd0Dasn5
iUbnrm49czwTs5BcSZVR6Jr1X7CqJ2ivMKBe3/3kUq/tTC1nMlcDSSXa/5S0
3dJnyE51MVhV0PAfD5+kpFtWcWoJnF3gc61gAKLduro98EKp8YH+znhADenY
nNProS5p2VYIyEGu35LsvsiFZa/uXBMVtqbpbKeHUlq7ipRGTZKiPvqUPrJT
MFp47Eql9+qjFIK7bbYZg4MnaaCrvPicNgTwchjYmYw61452OL5ZCjAN5jm9
CY4g8GgQ+zi4zs45qvxuoe2qj3ih8NeDIM5OTmmugvSrz+/KpSpArvJZGgLJ
FZfgkyQbxZoHLc0oMUJ0TUN1apqejDHaQPQ2Be7OaLUa6IwpRVBOKBxJSXpb
wgjVVf0f3Q0w5ebce3t6z6UyYzyfrTOudm2IHDGfLdKJ3XwWInp68jG8MZFD
zwGu7gYTz53AR14t+rUn/nzvKCwZuW4j+W4OPn1HGzw+5eeFGRzlRHFw8pGc
3kWzB7VfXUp/C5LOThzPLSeGO0rkUYMxnsLaXk2Hf4PTESS9lw6PZHnpCTu3
UvecEL+Fpurxjz+bsVrLA2TZ2zY+o8ypH3uQGd2z0rX+wn+eaTmJaEk/Xq4j
7azTgg5OSWrUlSnD353P38jYysMF9hGBGCzlCy3K2riIFCBZA9eN+Fb2VWws
dhcEKAM/F7Z5jRC9hC/9e62uNpJxudFJwQGKmf9mq+YwvVrlBetdxYrMyOmB
mvvr/soGrw5rgzMB15BM9DE2u8G9xcvcLR8Pz3pPINPNx/6k0SrCEdb5LyR/
r46tj1+zVEVnOZauJtTt7qhiRFV06cMxxox/zlcbGsRe2pWYQYW58AV2FbWh
Uj0T0iRqQZQE86C6t746JUJ1MIy8SCco0YhQCeJvJL+q35+FMI+5MhgjRaJx
DLlMU7XBeQRGOomdOh7ePj8PBq98JTle7ChcC17L7Rxq2ok9a51G9NFOjEnG
rFgkUkCnTau1oXRG0yi7sYNEFckFJqxCfTGYfECey84nf+A0dRf1r/9KHS/B
apkf4eEHmCuXWH8fBM/zhdSlxQHlcaMe+js7gt8ra0B5vcYE2fTtcHPtVPiw
xvSixuSFTaosdMJgCWuWDcuZykPfuKxnLsHMqV0sUlvS11r9vFWEksCSo7h+
xULQLRhX6hzNJqerHlDrfh5J6qhfZ7YpD3aR3fS2pNl536Q9bRv2Hve9sFg7
gFFhNBfdFYRxNNvTesM8CDcXn6+L66CAaEzi6EtG43tyNC8fXqs6CoW/OEhM
kDcYFdxTZeXFtdOHiyPPyRl834la4ZOSpibDuWa1+TtHJDMEw646yTuX84rA
isWml+XePWvCrH7j7HcEJ11OdP42nTiy+g2IvW7GqwCJCIwxSoEnSdPkaRGf
7HcxUcmRADLLGWCYJgq+zRBHGofL5oc2BsnFbg//AMYOE5LrkgxTOE5trI8l
JWgL1d+HFIiNp9rGpG5Ht37In5zv+9V7Q7RxrHmVWDJGZ8NA4287zl+C8oQG
+WLhwd+zNLGbaDMm0Hg8lmVwaSQ5zAdwN0W8LNgY+B0JXIHFyFctXV/PQ/PW
01DqWMGCPQt5QhV3iLN77TZMD5zU30fiqn4p9y+h+Oz0Ea0l4C2RaXLCLML+
32uOH5otN00oi4XIPIsnQqaIoO2L3sVSzL4JI5d/A0tGwUJ5dUlF+TMx+kGA
4Q36aw6TqH9i/UCAJpYGff9sZB1Yt+qnmpWHe56DcsxHhxsGM52RjYrdsMgR
oSujzwjPBUgya8yGKJLq4DzQXTHWXeF7Zfjt0QGIHypplFQkQxtsr9dskmwZ
NqneQkeZwHivrxUemjI8lDP++9nVh9PV0M/+yYsGslkTl2jZVF4fS5GJ77Qv
jh17vtUItlz7UcsDjGc2LH74C2oLPoY/s/rH13ghzMkiUTp7yHsCn0GszFLj
V20+E0gCPRaGy05mlc+U5kOItpMBVU0PIV4kYCkWeaZUSlBKgYPTD1IsObIN
Ug02MQEL57xzUM9ZpXtamIbGHc7a5eUelA/NgVPN2dcsKD/WD85ER3oqtFpu
kvgRsiNPgM4YSVs5zLayFcdQu+vtj71GSRT+lu9K5LbcdWntJ02gdQAzc7Uo
scID1+nztOq4rsmA8CyYzNzH8AMcFP7X1yaDtTxsxs4MfBRTToN+Mg/gXUhF
CygEbt0pCEdU/zYp8rxQ1KnknZ1TTnrjWRu54jvRpRIBaKvS+siqjpsW/AVc
quYBIT5yol/hIE6xL93sh9wZwkvU7ebTRdcdsxdLsnbvOp3l8I3G933ZVPMA
0eBExLwZvHfOxC8EXNeLZ2chUndXobvPWV22pEsFTTTVZuq6u389x7elVQjd
Tlf+t6DglH/ku/F9pbbxQzaIDwVszZ+L8JIvwmBEvjzaKfIB5YQnt+SSg84k
9bLnCJhJn+nglM8HJtxlV5C5nH7VCU1bqhzqy3yf21f1yXHKlC7OZgplSaq4
iYUevuvqsrW72DBvXy1bgWDivGd9OIrP2E8VI8NBbaaRdyLtVIwJqLFU45BU
w8DvLhO++fObZlVxXQigaTIhhqgRRw4GSkVD3XaG6mZ7cfoiS8elbXIir40Z
zzx5UwxSowXuaWCvTmxp8wKu0yRMm9xQRvgW5uL7qzaVJMM7yiQeQP+8bnY7
W9rwdahOiOghb04s2ceGBT00CX80/YuYmANc3QEqqLHTZ8u5OYc9Xn+nKxrj
voWDlvNGLHvs7uMHcJWSIfmXgkpEU6rO5Vd2pB5OnD7KL+EKFxhyvwq9J+Sa
KoOkaOstNtNExAlLtwlGlCTFsoDlRsAUS+RMnGiAAXmA5nqzZ7PDYi57NTfH
0fo+PltJqo4TuK5jo5H265pvzyxTCLbA389G+0xetNJe6JE9T93453/iBOAS
nOSbrhnF+svjHW6f6nS/NKWIo3svP8utWngjJGtNZodnjDgjczrsYh3Cvtkp
zwtwo1Se3RDm6nVWoer/ypE6cfbLAlktdiFR246oC/SPjvt1ZIjnthofQBCK
J6qT63l/iRMt39ed2t5s3VCHZ0Cyk2Ortk1yuJtFPV9aiERvw5A5r8eES9NO
ev5gv912EXlHLRg7AHXZIoUM4UmhiRbVvInAiOFhNYHctQwkiiKRFxbBRnOD
/q1+lV+koXtbwS3M9fee/2XH/qCLWcJubT2TDP6OqlufVoM94NJCIYZt/qqo
lHx/zkEbXNJiUAo+suRd/9cu+baukN0WH+R1+bkKtK/uMoKxlNaBN8y3d/Sw
pWvp2AT+1YdtsWM4+mnnCPh/8sWoEZFungKs8u0EwQFlhu5wxMb0206fvsty
9pIJDbWAwXwc4qoABmTb49+FgfPm2RDxaLtYBEvtVf62TJD62iymfTkcoSFw
a3IYVCSJYT4xPOaAyJCcaYCsppSZIPpZ01TN2C8Wfcb1FaG4eLcy759sFjnp
Ui29OT/zdQ6br+zAFSq4VYwWLJeO+N6hqq6xhAnfVqqmr7xIdchVU0rA9V0l
/r8vRGcMy9N9HtjUN30uHHLtfcJjUfq7mur/Hg18JmmDccSg0NXzTJ4cpf0X
jG0fmC0hEk+iwilm+6dv46Q1Ii8RR34GWy1gKtAFodkOChICchgUUOlkePOL
oCyOFHokJMRDA8jOmYijuwOeX5jpaM2KNQJQgCH+hYSOzrKYyYMVraC3vt+v
Usr1Ugq2svrV37p0ELTtQy/9B4JBrD0IrxN3MocOXpr8g37mfjYmqp4jEGP4
abA51fZeIyGSyzbQO5KdqlN+iyxzgWVzosQflblnb+sAE0Si36NNDDOT4QoG
BiDrJvMmVyDh70faxYEwWoSAzlvLeeSHgJoLXG54ENA0xB+rOyyK2fVKO58z
OEH+kOKgBfR+oaAl4Ukk1nJDXGm0TAgiYSRrRdAf0DLw74/QHMoxu6YY90LN
FTAMkx5OGOcfTiOe0eQ1xuu/XqzcjPZY+KdANWtlZBhCtvjBrJlRU5plUULD
QMIP73aDjkH3xbinAp6NfpLU5y+yi6WoZNb7gubZVKnKFK4DtmqFfUMYNrPR
LqWWVJ3Ibnb13rJmzeDq/cjzqMi1P4mBovu5baktgqmL6bgJEe9A0dp7BOUz
lQYXftkMUUdtmGcXzdWiHZmk0Oq5jqEsi9vTYJmp2DGpRyQ8/Ca64LQUW5Mk
pYxD1f/Ijafxng4KSUr5u1xwb6T8IewgpX1Vsn3YyWBiDnuDW18Do0OvR/W2
G4pVIEguUyEev5GpYfG8I1Qp3C4S5SatS9OUy7R/iu2ZvcIBIO7fkgYCh3Vq
J/XQi0dV1Z3BRM95tUrBaF2xNk7M8s30kqI4Vies9rjkNLy/IxHFvYajTHeR
sBtRqSFCurk2KFZAQBGxa8wB7nsUAoXD/vstSm4putMWAztnz/664hHC2dHg
XJ9QbX/D4M4WvKG54Xt3hIB6K1yyu15XzjfA00pcXQn+9wfutpcE95p0XHyO
0VK9V8GfBqi6MJOBSDNkRn6ebmQTjxz1fGs0a5M2LM7rS3KP0YGB46JluTpJ
hOcFx3puS2g6ZD95XyDnEFB8jZI09uaQ22pFHYmBakRI2x6KwjRfH0gfTelS
SS67KnJODRrjFHp7wzOx+gpHi9Ml2+gOOFXT1fyVk6gx360RRtKf7pDKeibP
7p4DYuvGgI7XiIc5uwPXME5ZPOBCwLZOcU96iGS1N6KiaYe7b+xWVW2CuuhY
c9hofnTzSV4m1qaNWZ6///ucc2MXZnkLouKck8cZHPt/8Ojr8/F+ejkR7Dst
He9d0k5XlesE2UmwuUl2eEs7M62LRe+clYr9BMCzZmEbSSwcbrv4vltHd7zE
79w26S6H0tOe44TdOkzTMEAR1llINY/XbFJVF0NKepof+mzBR5p0cfY+X9oi
1dlpNlDnJZH+OnIQoe43aqLmPNYfzo4TOvOeSkSaeD6oOB4ijhuHwX0Rtih6
MbD2iJJqJeYUQk/cRQT1l5SrdsCMsvv32EJjvGjw6cBsKbUo9PzDjijZEApo
1rbCALVWK4czZ6rioy4SJ9I720GsYwJ+Ne8HK+mIVOj0nTTygfn1rTed7KxB
QL67IpFLUt1Jv50T9SKPYu2j/2wQyu4ddCA5+j6nGKNth02DwPGUKPEaLq2v
Ym1m3TJLrQDkCKgj/iCEdGpsappryeyawmnLrVJQwPNS0AKlysGsIpzVmVeC
+x5rX8aTem8bC+WUy947QSqBw2LQcUcXg15NIYun/GndVeXECvkWaiBgvegQ
iGQ3FRLP8N8a1NIULPguZvRoigR8Rsb9Ee6XwuR0hehf4ZHzBwaBXQ0FsW5J
RpW/hqSQvkdgLT+XN3JZefMKaD+Hb82xH/8GEARsHmz+RjqH7Zsga9VAVTOl
qNnDWnuF82sP7vQt+/A9heIiiKZm/WxAlf1O3lwuyC2wyDtR5QVOgno6e3a1
kSGfPPQNxW9e8+DeEH9VlPzuEvl5UvB9ipwRQgDR5XvDvxG1yrgA6k37zWJN
rD1U7JSWRlfjjHYhUQoaHNjkQY937QWjpWNk+X6H2/T/EZ8t//v+Gtoa6XdL
TWxxXpZyRHxp3BFeXRNcOHCC355/lXpRU66jjgxjesVOp1eMBMIDW/sxTkd6
phPN+bhb7sSJlw2AM7aWa6/PbdQOZgbib6T09ZDHGbByvkI7SOzo4a637kTM
aFPp6IwL0MCKUwWswdwaXt+GV4GTcJ7qBwXf9flIIO6ijv1TIOntnvQkTZaL
JkyJZ1dAVwHkWR2d1fogIZ0G4qqZ5hbCH8MUwVmjaAFt3rAqzGYZRN/5ylJs
Q2T9zkwcxCtC5C7Iprrc5/xlYKGF45uVw/dvzXrrNTlD1/r7q2ZSS1pKlEBd
+TJKO0scSzSl6Dcwlwg+0MRuauy5M/O+ibEcWOScmVveOD83mIvsMLx1YZjg
MGpLEwqtxTjYUk/NETqhVuowhpdpoGsKE7I2T2w57ESd1Y8XATNqDTD0iVfP
QraHNFKru8AuvlAXE4V21mpGuVCeYUb0+lRK8iwI/xQogxkvpoS/5d50j3uf
NQIHhdXzH3tW3Kcz3s2syRhWiEvpFZhvs0WAFpX3Dwrb84p+i2zaBaW4pd62
dry/mQef045X3QqwKSMABskT3IO1kFzGZ6rAUba+nyDnhCtkyDNRgDjBsHuo
rPTyVQtTih72in208CATNWDGE2QUtyol5T7FsUDVv5fWqcAoHDij7V+7irBZ
EaPmedhnTjy5dAdVsaAFXHfESoxm//rD2QmTsIUt+ZbvFLbmP3ep2sqGF0uX
KDL45S6hDP4MPK+WKOyCRLiqROmy3ibYRn16maiUjNY5SOcUvMTeDo7sTjvk
GvXdd2z2Gzk2Ykx/PFjSC6ZxelMl8vR0N6ODRc7O7yBPxo/RhPtJGHs0EApi
OJGyWyTFByZEaGjgKB7l53R/2SsA07ZozpRhRC4D3D9CTXWIYWqwihx9qRxm
1EmVxz91AvVkWPx6IkglzZkpHTwpKiGNopDqBUq8UpFSONaoz11tsbgkpMsW
qsBPS6klGGGsKF3HvqalKhV5ZIKoLXj0+VlzlHw7AHcw/SftnC3NYuraCSfl
vzfTq1LwTAbz2vG/P0qPPEJeetWpX8y9RoxIQ9rPx280K9iRCxaN2Lan6lD1
VE8VrMM/QHUVAYrzAGdMIHX2allPu0ROSyUx7ZhmiPW8HhL1+5VL7QtH9LsA
zKqKhzYstNF10Zap+irgbzPpz+nEgcClhNXHynMAB3lGgch/rRzk9ouOzPRX
gsRBCeATOcjjBa9/0+divb01VtM3+9rdwvaHNMIY1pJUxWkkXczvyTws/M+k
BFodMNmN0V1OO19gU09N2f27YyecslVHYrK+Eqktwqb/N+jlFRIjsssjGf2D
KEx/47sNUuJUX2BzqUXjx99UCWfQdoSiyMPNk4riEomQc5ktSwV6H1coTBey
ON4k7H9dTBoVHXHADHJhaSTldHMMxYBTaNXw9D/cI4VZpi9r3yN64b1v9/3N
7O0qiGMmR7XaqeXV4HeXYjvHHQf3dPtrj7z8/eN5X+V2UcdhELGl9ZmHkvdd
Po6cl/jRYTYUiIrRrVLbf8UvJiucpRfpTnzjOCtQ5TGQMG8WyJTk6nj++BWT
R6CuV8XoC9QqKNVWRYBZfxu4EazH7XmFbquCn0h4qP0Vh4LxWgkN5AYMKrm6
TZuxMoDoaXTLJK0bnbR6dQ7okaTAxbX9+WZpqK518/bduDN0flw42ghF3DMQ
GP1YJN0LP6F0KGeFrfvazStIV0nd56X6OrAgWCtHTIP+BCerRpqIjY8FXoXZ
xkTGP9x4ij7KoAb+T7dfHjJIKNmKqI2yLkocDtDhovfIfoDlGNB/fngFGPhd
mhjwnAte2ccwpfglNdKSvFssVM3711K7nJo0MzTu5tFUPF4tvWR7KBTAb+sA
wLYSsIQ0LFLWcnFHC2wSHbNUy7c5vaNShZluIfgjVNjYXF2rU6uIVQVIWlXU
NaTFUyYLij2xRU22Niv8aVZO/cO2IGq+4GWuE0xrHTtk/2yCAyJxRLzuHmSQ
2MyXJfDR2EweHKQAO7PjSsED1vYCUH5rxRDQRsCECJWKqpYGCR6vH2fMv+Rp
qa5dHg6TDbPZ8Syv1FrFys3IpQ1zlblG6AtpGAdHsILQs+RZYijP0GkDEIjl
p7FwoDpAWLj5JoJDnT5YpqDRP8GLwiR7BDapwqDziQEVof3BOrBvIP7sc/dw
NPNt9yruPTGOYyL6Rxdq2m++0AJkbJhofVmsNp7074uJpBNGGNtBP/sEgq4N
z6ngQ6EGpgQzMD0PIG3ft2Sh3NMljIKYw8S7qVBewcCAz8YRHwVaubwThmse
dDIJRU3DP+vzYGzxnUUaIgaskUJTwwi2PabpuPALxf67kRnm4m32AYiamPUD
3p86VDsAhY5hV8cr8D5vpDC+gODtAO6rxz+2Dc4tVY53fzL8b41EMUNyuJ6r
cQGZUjp/uNXCoHQP1En0/WL5uFLvnOJYoWxGIVoIE47DvKgrMyiICfth+GQR
JEY2MsNts5rRD8oo77MTh0jm6qlmneqGuwFBgZDyWcC+wqPOmYrwWPxjXyQt
vKXjj9tON8vcTY80I+jmBXJ8kCzNqvZwM2ns1hwemUPDJWZkq2hMyHykfCOR
W1Ib1bHJOuTKLhvdf5fz9+7YSy43PmYwe0JYCRKb5MQHPO1C6gqwIjnzVJg8
dj8NaYsbdyQ+TA1F0KceuGhP2HSvnoSEBn65xTXoUv+qHww3rj1H4YYVy5LD
Ulr5/hjNbzG3Cil5SP1VC3ktKZ+mUAkqGfm4WDm2gcV2n+kdNpaxJaGuGeuj
z5WDvM5Jm6LFqY5mq35kO7J8ajlL3PliJcJMl/LjVMWZwX7vT+TwqGlL6F0j
GORmE52GHaF1cv9pl49BO0kuoAyw2Lj1s7vR/42TyIjy1KJ25cbyeKVCERxo
pYvzroJ0kLoN9B7Tk1uYfXtlBiNkzZSTFOGFZhyO0iMIw82qNOozbVo4O2uy
NKeThT6rh+EJnFrnE2ZMbyHu2+5n9qRUvLwrqjmTOg3GfR1xU92mxYC2omdb
x9R/7RS67AbkEmWKBBAc0bZMAApD3H1u8kkX1bGoU90uukygZeB+yI7emlmr
t5PJ9mT6N9G5YbATrZkCqLAGpoUkjAkFZXTqvEnljOPmz2bxf03GTg3KqTTm
LC8DyeSaIbkPWcCYErWZjn0RnTW1Yiqg5ga2/XC/RJKS5vU3nNT0IYkXRRMV
yXZOV1bNW99NQt48iDOIC6MxUuwb2+uf7pznUU6EFuxmix8z22OjQLxRa2hB
btH0tRV+8KUvdPeydeW7MenTYjxaNqy+9JKH59Z/fIibNq3d5qL7rG3F4nKM
zw+XEXnqGG0bw63Kj8nxABr3B+N6OzDoT26nPE0AFltet+P+YLxcdHMA40I3
uzMpuO9UOtgdVEJ8TINOrURhflEEVpcmBg1sepbhAAWOVITYftBSr0zsJX0Y
0mUe6953FxpRSi3dymK0hCTyikabxlQFIrbd1cV7wQHKofMwjo8fmARo5uTn
q7JjjX5ZtTKPIwDP6RyFRovlYKQ7TQXiapyOezMEDFAWyuUAHTxS6uqd6s3b
YTIFvwCsbnZRc+RMVGQpmnl2NLzbcP/Z7Uluhq9yOysW2QKlM7AvoYgENOrq
T62ez7fNVsqqu9VODh6QcEnDe6capHBIiRU+gytWoA7+QL7QFxtLhk9LJ5l2
yB+gll1lvzrXQpB2gfxwiU66Jv3TtKgm5E9TtgyeWzmpyMWQOTtGXyXLok9w
ngWPl42cv1Z/6Uf0a2vns89ICE8PEZOalXh/nQq3TtHAXPL2myXickUCXhyF
EYwRim9pcMR3zWEteKv5LPy3AztvXVu7XBW4LPG+3rdXZpA2BA1sWe9tZQiB
hd6FHWUM8JmkyUpy9H68H8OfubJuaXhfTvjGHuj0FqO7TBSBJfDLOkHrQ/tj
OU4KVOob6/NW7PZyBZ6r4XjVK7ENfZRbOqj8dnCUY8ULYYROYU8+kGpr1qac
MR0wG3bwAivnNFduOJXEqT26SadQW3rc0vGqEILCpjxOMJR0mE3IuEiSRyUA
/KVrOT+o4TECEW43kRtLdePZTHir47wS2jmKcfaEEE6/DpghFAx0Bfppauga
3VhZY470mxSJdHO2Kud9PEFt0BtuWrgYWZFjo9pzCSUdU8oPgxWs4lmsRH2y
SgVnN26pKmKPuEXurAR+3ApemMBQGXl7EGUq9Iuh08CBTYNoD/1V386CcMAU
zPPy+0egpUznUZic+sGXb/KfyzPDLe3LSQBNkKLQX/eSC3z9wtpwrE1RtcY6
CnTOLSyroZF1is2OGH/vNmZUjTr9+Cw+dMLNybCiIpEp77LXO+oIbEf2JUn1
vH9Bx/zEGh74l+U4r9Cbzo3NFMbU7UyNrLLWb5JgRYCuyfE7o+mrPUekdgOM
TQqXN/RXPKITYaiHi/gO8d2k8S4NDwADO4cvu4GXrPMI786q+5OUI3/6zBc1
mrY/neQDTKiZEHrrfvzcmEDpNAqhUGEHsuDB8wAyJfmDzE2INxHcPfdepg2N
/+g8NHP51uqz+Hv9f9Wxm3ViGfVvC1tDJHcAGn5R0i3wXU1pgQjAR6Ux5stw
mFC1v5jcT6/HzfcH/UZYvMoRl0Pn6gsSmZM40XizSjsyObMunGhJojCVDRcp
l8zONnQ49Q5AXdYQsVhxD8HqUpbFJ7MnxtMWGFhhHGvl2QK+Lb/i2eIrfcsQ
0Cg2UBhGf588A94jgPXCxvkDlF6tIUg+2pW2l1PnF78Ovi1iu33xZn/UQfVg
QvsWY3p1nHWjtHPVZazTQvEY5eOM2FaEyypo5Mjtaqz5IBVZLGoAREwOa3TM
gkIYNvjrcZc6Tpjf2AnNDU+tbPZ3aO3zuhg1CShPxemjKTjLkveB1Beqi6T4
+7V2RBK7CfYDDp3EUUZuF2mKdqaZAjC+kewUvZ79KMvut7U40AOH3NdDH0o1
nxg9MRG0PSi6O1rWRBCAKxEGUbvQDPswvIxjLjBCes9tE7QXCHsFsRfzzXSr
GKbX2ncfoaUZu2U93UVwPJgTV5PAAJUDTCDcwUXW0wN1KYflQM2MVzOrJz3C
hgZcxushmE3Ig6CFBeMWpwWb4NAlMIyjh+jL81uQLr+aeQ8RLlFjOkzH8xmf
7zVk3LZxvEyVqYU4fRavYoZM7LBPcQCD/bEiaaTvgmiy7OqSw2rO+4UCgLn6
lUE2CYF/FLBCXLKzqee3IglFlCVLna53rys4TMvW7v68i5OLnE/XadMOhFBK
drwrcqi/KuLJZBalvJD8qQLeDvzl4alGWpJyxsNFRVKxWQbupXfA1wNiOMk0
DlJsNEwFlEdR7FDAftTo8qTsCweXAw8rVM494RE6e0wqLfqTvp6bUysSfe+a
s5C4HsDJyz4BjhOMyVLzFaHErtbUal3CyaOWIoZxWYLBAGsCECRANCGf9/wb
gD4iYda0G4ySGH40hakR/MIUjGW1P7PkAEs0uUnsTU5/JFTfSIvMQ61svPJo
90mWx7p2GRD8eReA3VlInuZKfhiYtJnk4PrT6LWx7Yke9i+zKKjeTjm+OIyT
uwPzdhkFilsiLBvtfQ8G9FAw03QneoEJqW4HtLkLsp91srvNL+4ooiaFd4qe
rvsuXeXukgCjcors4z9By5AMMDMr6RoEqesXx4dd9uU4+g/czHJGLVziGneC
R4+ACTmSijeS+thw1TseXEWROheEJbMYfEVDHbC56GJ9HrTQwuLXM7Xs/U21
NIk7vryYAmH5osdJOWWSs3ohpCCkAk7CbDBpgdiMRIuOAcXpHnF9lOfxg3I1
gTfCQkVHV2RVwq1yPDBUge0ltv3esc2N3FkYLnZHzXGYzyF8hNZZqh+Gp/3b
njwZVX3G7psiUOKXj64P3VHXFjEE5HbQSLVemiiTtde1YxDsK2yittXzvw0b
wwe3m661chTU2Ie3TzjZDsW4cY+FoqXoV9hCWiUDR5wYFt+U+m29eyy9fm7e
0PSM2/iFD92veRSIOArglsICAibRYHxEIqab76vkbfgwLyuxdN/wzn31kzAJ
7O8fw2qeYLtZRGG91nDsLPHiMx/TKjOFOLbIADFXLv3h81OAUFZwRedLx+2Q
Ni5i5NcuNw6oIFUEeXs6kuR7eA0zf4DVpWibQLAyy8IaTO5GmLIMvMVaWX42
wM279YIUMucyeVQGmyFC/+ZbnVbZJJzO49QsQmWwWM2dHpcxYy3+0859vkzH
jMb35LL/OjFLcDzjgUqC7uCu0r0AoMZ+3Jf4pJ+UVdiy1IZEoI20AOKm+ffA
FygX3SFyqNAnpX4BRODU9/iWt99UffGorQo3sJe93y87rx7MKElr2zYAe8go
Qb2c5whVzWEbb5BmaRfS46T9Q0vO4hd9pOVYQxj2TtNxDrvS2OYUQQlz1koy
Vc6bv9BLy9IRLKqs8/ukmsqg7sK5JpR16YEl4gmX/Rcl/bCuzItl8g+u4WAb
Lx3FMZWr1GurXKFGYK77r8det6DeGdv0z1i5Xe3SIVWCi4iNLYlwkWOs2GCl
79jYwUm1DSulwXGgsH4ulkAvzjwOswFPGQeZJiplXbIH1tqf8vC1HR5zCg+0
RTNDNYFMlt1M6fO2lVzQ/wtiHHDaR5wMKFErzahJU2lA7ZydGKsfOh4VNeBt
4oTi0Q5mFNiKnjp5tW0eWsIH1a7K+HZsBJS0MwmEZc+HiibT5kZpTA2SYCKX
LqM/3wmIsmhpEeCGG0HRP9eVVTZa+BobpSi8WADfiEraN9TuDoSijljimFOR
OawLzek+h30hJOQP5m8RdZcb8s/JQskxfCv7P1jzubAcyXWmrxItK72noXgo
WCByky3jfsnBhY6p8geA6xLnnrFWLtVodGoNwNfttMBAA5RBg7g1iCQ3tTS/
8trJTUFay9AHdnEIaE8eD+4qbm6f1tbjeo8iDSsPOn8LqELG5/3EzgEhojBI
CREVxnR0qj1rWpqSMrT2/6b4Kk6vxGXsBpGhrAPQcIAEIBjdJHccdIWmrmCo
fi42qEF0knAjIFiUaxBPspj/Iy3BvEQzu73WbaohyWU85rJQnx+UgJYQqw1x
/g6q6T0kA9t4jkxNK4G9oMmappFKF6I/EpL94Ki5UmiUhB0B9YYyHrwHOz6s
OqnWerISAJ2knd6Ajr3sWUHgn4XVl5N+rtN4VSHeeUyyPZFCYEQJVm1YmiLN
gGqTeKlaG3wluC0VBg+yQ/+nc+wbQT/NOGZUigp5ZL1J4v7tDeEN9q/jwm22
kWJewpWdHk+0DnNp5cRHWaSFLWjd4c+CsVjhN+3NLvqe0/K1P4de/LDLfnyP
hR0W+ECMimlLWzVVJwiaLryy82CrLMgtOuEvU3kTAguY2TdZIlyDcYcLZ7oK
nW17c4kmn1TuK4a083N3/pmVcMKJm161JmcJh3gQ2RKtuvIzsfuGTSq1PqLM
uGnhFxcW4ze6bJ8Ro7OO0Uufm3PQF4sn8Hdt4Y595r5aO/yQ2SljCjtPk751
oqy5qf8X5BCfTIMRRZ/nbbxUT0ZDC3sLkoY6/3z7Pa8S2qGTpI78a1o+eDkg
qh7n3DALkq9aRkwasSfG62rjNuLH1gi6mElorC2qHKcuNoqIaVWX+visV2/s
igZKsOGxdEaL2VDSNVhRBdAVRAp1DU+MS6ISnosLE05no2LrY+u/HB5lJRCH
hQn+XcvH9DXzM2d7c3jJ6S6zsy1Qj1a3PuAThURUIeHV40V/RhtHVSparmZA
gtaZj1UXtqPP2gRW/WD9hwJM1pc08cqwbRnEqGeCPD8RQB4sOfxMbH/bnocG
jNv7EKXNd/4x3LS8O1BBnRk+cW5AqW8whaKh6UBtaAb/3dsnExCEfXWMQ1dl
/1g6WDdMWsnI94s7NhTkcUjdzCVDPTLsggnDuMT6Vvm7VJfr0mVd1wWmmo26
Jv2Tc5kyhNXd1K+ct45rcwWTlilEdU5q6uZe9bQJWm3wTztOQx3UHEx7Tm94
cBnoO8fIbyF0O+rPy/5Z20acu0MCsDxWLmz2d5+PFtDWgBK2+LJBldAcW2Lo
nNcq5oe5en0w0o2iwOiRx/UO1gW+B7ZsQMyA3IP/gDIrqVkFgkIF8ah+bXdv
Ay8feMoNPlSbeH0G4t6esgnfqgCAs0HRsY8ENoRvBUFavcxi+ZzZm4YxG0I4
DWE09CABa3nr+qlf3HWA5P2XuWB0MeENmB5r0UWAr14RYTUyGYvFNhKARLw1
RRTHhuiOX97O94nLuAxdbm44XBl+bA9Jd7fQIcvtTjAeibDQGxBJtW2nsaCu
YbEMaCJI5Hstk8SqpTMSVcvAIDoAj4IybbeknG5cvOhcLEq3+RCoVYdyqAlZ
ZghKDue+iQSjoOS8NbXgLxuIkqO7MFk0qEy2YXWcdyKncKTLKzgQwwjpCIfF
5UhQhpkcXFa0fhWVINRs78psag2vk/Tiu+9k6oZJpitBlGOkJOL5Zhpq8tzV
q9V9aY9gJKR7SaTzWb5M9EfB2STH8rrwaLQiBOJk2tp5Eit93ACA31VDYhQN
wFU5FCZQar9HUdptE7/EWpW1pMfEmJK6OefOMuq11YqqSNoWwOsyHMEyFMXS
FE40QTaw9BZysbF8o41mQB14Nl1YpPrBeAb/bH62YRsALmkkeKm2NubTXTWc
Ywf7B4EADHL9iSVzj52Rza47zggZDEHzJ9eg8HFVIRqZNvT7G2TjLFXjcg5D
/PakZWUyYpVZ2kg+tBY8lijUNMl0KyVEWmd0wkd1rAOdVZaKccdVdcv8euxi
eZztutIEDBqmaJm5UEJrZdyFqBSFha5n7TkFxqW8ZU7H/M60SPYTfsQ9pOyo
4o19JAL7uI1bcasm6Rc19RgEHNosV1vKkTma9gyclts695kxyaP/J4qxUJ9p
ayKA6kPssfhYvvkOEFxtlvPcYY5jDzaLvB2SUs+SdKCrM6ldtFZwHwkTX9Va
TXekyKFS1PcA3ROJlmgv9oCACVLqW+JsdjchsFNo6sJdYDzRiaFjhJ8cTrIV
UsFv9jLKwWUcyg2/VWRAlh89UKMdBXvj8PYL/5i4ayUZMivzSwboN4AfxyXc
dxwH4jX7kjPDwlRLtfU1BKy6G8O7mB/H31MlkVEYysjJn5fLtIDBWCugLfNY
CoxhQXp8ZyBhjSRol2r+HyoAgNCwM7uuCr+OoC/slve4EeNxQfoVXoowU4HN
YW+1rl6S+elJaFyYbGtD17cGocHTN8N81C9v9clVNX2C+5XFKKHsFF1ysDK5
g9Kb3Rwxr8YmEjbYCbFzkFfHLuynZLV4ZuMRPaKteztO5f61Yiikj+pYkXXe
djYtJqNNNZSS23HCfkeFtgTYVZZkf19eZ78+ODC8KwfFvahwr965lPEgoVnn
aewDwIBop30h2cFaFFXR+laIpDYhR8YlQs7n/94fptY5xraJ/vGFPCsEsAPq
iqqXjc6u799iNJwCIQPuC0MBCjTcawlQbt7ZRdgdme6YyT/v6SjrUrOE+g/E
CK1SEDXxQphMMmiTsrJOuL6Mmt8gWgYFZfFFIeCP2MU9omNGjRkUrDASc7sD
H+SA89vteIkPCJnDsaTNpERqvRAE71tnC4S5O2dWVH7z77Rz2JiEeEuWxqHv
By7Cht4xFJTDeqTNqXUPsNmcJnckG3LEt+uewDaYFaYg+s7KWPBfwT8XUKfZ
2DuSu/c7W9/xP7/YTNFmv72+XEFzjsZU13WZsERR0yQesAu0zT9jxdOxfBnU
+1oweuRbwjAUM0m1dw6C8NxzVhNDZUrDlX5kpINiQqg633QhABgClq/xdqjp
ohUifb4nNbZ//ceQZhO/H1vVlXGs0fOYxj96p29M6BIhM+DqbdOxxaLuju7U
ZYAS9JolPPbUrFieR+mZ3IJm4npg2WvvFmKERLDUDufl0gS3lWWVuWYEd7If
6a/ktZD1Fz57yOT78MDX+xbjuJwkVlpwWuiWvXED9kjEHvomWYVB2UC+cvuo
cfHj9/V6YC0/WyMr0nBe1K4jnSFSPYhQR3zMnnS83MQtD+pjX/qhdFeyq2L1
Eds778o77GKIP4F0B2oxXBXyjshMSxevXZ6mSyjmROW54wWe85yEdd9I0uTK
fBmdSMpqN0Byci1CGgFiCskRu0jrXxbgwx4lhAEyHkLf3yxLP479QkgMynhL
5r3n4n6iD/z4GCl6QfsHi8e/96mZlrJtpn1Loz8N8yXzFmXAoy2e9sflIYXm
jvGLggXQ54NCoXdE1IA0H5ovzTlzSghS8DYFJnInSVa6RTBguG8SQwwuqTZp
PkZ/bn37CREMkxbCJmPRjmjr2jmishmNLD4ji/vQjKgP2i1YZCYyLsZg9oAL
IIVS/wYPMpiz1lEdDqF0XKBpMhf50ZGhQ4rlLGcKqVjP7ZarpEYl5tLapkyI
2g3kclHDhdsgrjMZ6onmxR8Fa5Fc6PnazbP/Y4MJlAZ5wR2YXVAvYrbtgiVP
ETC/DMJklWnQEMUet73DqXCI1hKIXWe3tf2kzoXPen4d/ssPz/G/AhP9fw9A
fGJ+JaEkq16NAOxy95W4ibRJ5wfIz0o7hvT2s76UbEeun76Xrqg20q3T5UeU
biRx2FaUo0MfMcXgK1VpkRluIrSHtbDUz9txQ7Wpct2t2+nTwBsj8nUi/tsD
/rwFGKdsnOOswil8gsmLfQ0g/scShyhIZB0NsfBgzauB5K9gw+HMJbIt7RxY
jVB96p5vLFE62vYGDrVGCIJvDai59ux5gR9oTriRoLO6CitJgOR5PpbSFWmy
DsGsTEdyFjAWWABWXkp6WhjyfF9ii8gOpA0hJvfvP0QTKQALufYYtonzrq57
I9FfMsfbi50aNvsFOW8R63kgufLhGjE9NNBEODz79YO26maQ+nRfQl8MnDyh
DKtcmW7GX4LR78t10Qnin+WCUQUAMS3pcXoKiDaAMb226YSdgGpf+G1d5ZXo
Kto9cxEvSjW4EpQFBmRYzDg4XwSwFIy3Aa9+60langoEzK2mGtYp9u4RGZW6
WqiDFvSyAA+fX+LDvV2H91Ptm6a0N+Dy8Im5kXk0bPHAA0bPOujEb/XfEsIJ
+XP+5Tt7ToDxGn9jqBfrrdQMJc1aMW0fNpg9dxtLAhKml7JuwWTWl1ycgCyC
m7iSfxJS5PK5XzRLWFbiqhBXyrN1hTleU038X/l9UAAcE0Y1eXubsR0ezdqg
vW0BuyYDSJrVeMQNoss79H70PKxxravWOVLcp0RNSoScZhSybQJYbtvfpsxM
kmWtqFLgQ4azn3/ksr8fpqiuxccQRUXIDwTk1F1WhPtGlpXe5MyUSyOu8XYx
GqQcYobzWaujlw65rzxd4di4UaezCig+Lv341A1LHeFeak9/KSnC76ct8uBk
SrRJKTMdNSl3/nBwRjoP+F1Lyjx+fMzpCGaimupNwQJs4i/bBpoH9aq5KLme
LsdZ5st70z8ML4MF06ZIDMVNVhp8kKTHRgM+TUWPF514+jOhS4KYdsPIZXPL
D4APaTlE3ajPQhsrDKDmwuRj3El8Goelmu8rahkhPVMoxY9l9fQKLH18+6Pn
giC8H4WRhyIQi2tLqIUnkt2EIFs+uTYoT26BKLTe2rngGGvve5cWDWbOCl4c
fYCAQRqjic47ZkeW8sfCZsXS3sBpdkJviRGX83DwJb4Je6bwHDEC51j8V35a
t/dJE82ofmmCdY+i6Da4k6D16lH+AueiD6guKEdglA21RZoME4U8NIrmv3OR
ioxjAWwcAW63GLoFZBKe0WHGz3Ys8XrZKGrqk8MxeILaZlvkC9nPCeCIWeOc
8ibd3EmLslhTw32Vf/x3f7YSvCkzU/2aKivjELjlzXOlkbS47c5miOuCqFvp
hqLvuIsv02rqG/j8qhtfJ2eusM2SV0bB0ygtk8mncSIDx2eULmPsdqqq5oJe
Aba/OMrCciZSEPpkof8AFgSFWE/wyfmSYjhmXG3sscKbEJBAXIdQTDscnKp/
AistnrENvUOLzKvjwbVAB03TzS8Q8gjLZQo1/JM62BHRG6DaBEmyLq01NVcM
TWcbjOQ/rFmgHKkytfNxdqe1x0Qc+rlTr4mQisRiPyL9q2ceCRa4Y6Ek+YEL
cW9cLDtK7S8YCu6nILPe7hVQaZUYV+KT67ZylS0T4heYjgYuUlix4f2XXQCB
Or0pRIWAYIpHHM57gpl7McUYc6nrAkBG7kW1wSJtwh2FH6/6ka+Mpcp4XqG8
FJ/wc5wIQdNw+T4AY2huwByamzzLF9tFgTzviQfvHOsa8IYu4coFPT8xULO9
HYdIsfhumIrv6xfWmHukEno4MoWR2U5hQFo5i0rXiNdFR0glPOpqPoTtxPRi
N+Sr0ryDxalCqVsx4rxMcl6BrwO0rESjHqnsTdYn7RW4qIMbYr8PNQM5LH7z
lIAfTemw1DOpdYS1ZxlgcvxxMFupzhKpWvvEFS4qv9vdEZuHPraYwwejSSdA
aiv8kWi9gY32Z/lNvoy1wqgSpEESqiLm641Xi8H+nQj4l4XHOclVRwzw6+qF
sbzBHpW4kwBxe2BWMNbVpbBSaNOjwxBYiho1A0cnTVsrrO0ZrhjYsOjaVM4q
90LvjEsfMO3B8n2ZM9i6VyR3wNWJf8yQa5EMpC0aOCP18aRxeRTXst2T3d5X
dk60R0DcB4Jlow1JOf4pxSeGBSou9cy+y21Qq584+bOhx4QDm7RF1brRYQxH
C7lFK0YC6yraWZAm1rJoA0EmHbrZUzAJUQtz/MhQG4aoCJVTC4QdQPwPupsD
lb+E6xbTgz5o1kOPRsrq1f2yZ+psp4iCyR/xFH1oaHsEhay814vjjRFUhTQx
xWaSZFvfNpdaeCfKAikagnfzjPn+m8C4rGqnesou8LiFudCpgh/NXJ2OoN3U
eSNIYxyQlvtkMGPFTjd9jDHe+zHL81txhVaPV//VAkXDvyLBUTfeBQXbx/xh
GwqqQbyDz477X5cXk2ZpglEumWIyh4x6BtVgj/eYxVCD6cGwU49zLJ+kqBGb
f0jenGzFCBe9ugoQ+EkY7M2giUTT5XhZEfLyfgFlfTq5k28sESeZVHDWHDsF
HfszyfGlmdm4Shn0hEWDby6PCspvqR2OU+nBE59V5jAWsWwo8cMM8D2LJlCn
45Znq8UCPWmslYG8kMK6S/iPIk9Z3tAU89HoWSzexNyIEapHVOooV82gKWIC
uuwfRgafxzmXT73Y3aEt0IZnBsaz0FlhcoQOZSGis33fbrlqmzSv4l3plV3V
wDDw6VjM1r3CnaWCRQeiaucQ8izrXj+rXOFkdfqlxzzOxCCD1dZjVWdKCY6u
Vg8abQWg1ERsDJus1tnnjj8ZT1swYMPWdZ8gwnve7E4v+HZwI1I/oj9TqLQA
h3QF6XENgQkk8QaTRMdBGj+xATB68HNCPP+VeMYyfbbB0XZjCnPX0X7/rFKX
THZ/jVWIVYLHAprAUXd9H3gv2JHI+M6S8ot4Mdrq/eJp+LiWsS1G0kU6kxHO
TNjQivv8rdfkKDK20jyYLMOR7WBzQf7IdKyxNSrzf8Rz2geNLbc3/pOSZ1mU
DzEIm9EUMn0FC/9w3WFU4L23p1DVmfvS5NdqzedO9Y6rDQS74QPJ8hUOh7fc
i2u682LGTD2UslZAniVB37+mvwbnKievEORe9z2qA1O90MC5zataeaKk9CSD
rUOd1uGK6TJeoXE7DNp7nOFuI+PQmw3fMjaHiZ4vxZIRJ9wwuerRYN5SdWCO
SG4WpAN3Omm9mh9otpu13cXxX+DoR6UfGn6ZNRWA338gt18qy8puHHrFPIca
JrXflOmV2JNJWzH+95UR/OLBsoCxO5VE4+1FpRsaYw80eF2OoBHsslCOyIG1
ZIcgUW0lyjmQe2rw7V9cQ+l9mtYYv//R5HfjI6jf/XEKmuaoVnGtUMGQVIBS
0xubBIp45gZ+qjPGhoRC4EwftjvAgEoFwckTKYAgeJ+fXfUHf9XmII6VFu4F
ISw/Mr33xO4yQ0F9i1tuqH7mLeJseh1aPNC/d5sRYd5qBMhJtx6ktAbT5+o1
LjZ3XL8JAoPUaGCNx4LOyQ5kfrIB/Lo90dTKIHHjFciMfvQQWhJVxLRR1AXj
0HWyhBE9QzUPZhqz8yyUqItJM3M7yFiPrJ5ougc1lI8Zr5DN1y9k8UsYbmRh
2CFHqYkJPaNJKMzAk8TP6xHIYlxvKOs22h4Nk6+5NevrTZZzIyHCYQcawoWr
1Av6CjBXl45DB4iafgkwtlSe1R9z2pgo31UoW4wiv4UbDW/uMVfrxqmUfGr0
sUSHIxgTNslkM2PNlQwVNIDum5HRMVwPYlmAizV1xFWCNr4efE/QHqOfVhaN
CynDWNowaoz6Ka6Mk45qAhZ+55S3ZFKp45fxeHhie52otF352wtvpjbRlGfY
p22SdyoDr48IQ/d5DUNOd4oto2MSW65rCrNpUG3k013N8HqDvAZDAddfw43I
632T5dTUuE+BS8OYJIsDhvzLbv8aIAvKMGyUd6mCC16E75I8B6/mpruH7zUJ
BtjPLvlBDpvgbzHCD4QSozEvBlHAElSOUihojgKdZWiEr/ctlemJ1i+QI3Es
MxDqoDzgi286j7p2D41Cx6QrJP4b+hdxEzSKCZESF1L5PGe1RRRzqVD7PuDK
BJZNOv30S+FCzCa4iWzOxmUDlURNskSeFc0xiJwtlpj8Jd9R93JxVwQpuSfW
+dcbncS66K4kZzyB1Ad2CdeKm15JRNBB7Lb/n//sQiCVTDe9/UEoigYWWR3y
l92N9MS3aFxayDLvEvGuY1pILJbOS5wnOVNBWDdbcpqUwXHSpR4MCR+vqjf/
4Q9mg8lNVN+Kh36n64OJ5qt1XfDtVORhphEvIMAO5ETHnYYWrEyJ6VqVPUM8
Dr4+FGKLIDSE7DB77BLriE9OFkxQ0Zn3H42Qeev/oC7iNmtoZppiFhaukwlE
bGbWJGsNmfY2FNbe+BaNoKQsepftr/E849+L8bsJxvG9TQZLHMo4knhs207P
XFNwMJp/mIivGIePsLdCu5OiNi+ULMebflsRxgnCN9jA0TvE94Tbr9Mrixsd
VNOMnScMDiK9Kz9F89clAO0Zuu1Z0XupnY7fKA2/kvClojxPq3/SkLmNt7Hn
rkzT/aUfpKF8UIFwamUq5i9//epE+r4aDxlmQgF2lMzsYTCNzWxERkv2iSvX
MYHvz9sXwDgiLDgZSa9IaK+gACAjMiLAOBl0Q0VVDyy+e6vvI54pNFcStEaU
KmjF7OuIXGPHDboCb9wE6sdX3F68Qnd8oqrAFZTgxQQm2ARQ7BEQn7sh4qhm
0YVqh4lEw67WAB3Js0wlC6ZV7brMF2YLmFACeAWG6PIZPg5GPJcPSfpw2oae
kpjz6rJ2Glvukv1chEFrG3iT+sLEnixs/CjdkNi9mb+pwMmTyZ0kyZN7sijA
QSpkSueRyGen2cX1yuDXX7Boa3ICurIEe6UmYGPNPwzW1pw+9pf868judtpK
MCLWMXv1vnEC27uF3bKQmLgcI0LZfNVCl6P94DZg2U0cQO5qF57VTCxUwGyl
BrGYA1TxgjkGvS69I7aONap/yt1zNt2ncrhu0W9VycLgzrG7MjO4rw5bRZP1
mJMJnLo857FiTJXBgZX0rMbtrl7dkILWdBq5O5eVtxzF8a46e/dnpEKC2aaD
DjAbsDHpP+eifo23d8tWrwIZ1d14dje1jhi6HYjjj27UEavbf/rsa8boEyuA
maYoHllhZiLuJuktrwBYWrEaHdnTq5uD115FKVl+fKNo56on8/iI8C9KV4V3
bBITl4rvG30JamheGBvUpeQLzV2dCZpBHRRvGXGN9xd+EOVprDTNQlsD8Am+
z6T0sMw/GG8RnFkZ1BhMXocH0G6FngUQdvsgvTQGAc08xJF81UADHFo1Nutt
QpApCvqrf5HS6qdWjQ+Z9kztpVLCEYWaRZw3+mv6lEKme24ZaARb1h3KBJqN
fLQO23vA8cwSwWM8G7J5k7E9zyQho6HlKxhB3NfTd9nyvbJo9pnJGqyLDoHt
Mra+VVKrrTcVycUf9QvZWppKdcjmdwv0YBFgWBzJNc1/ZpOHM+nx9q0l3FR4
SHE4DFIw2Uw0SEcMmlUImibscX7PxxqOzshuwXUbiMolX9haOXvX+m64jUVg
oAA3qZSzgMwolmRvpb6v08CpZHe+q0xSr78ubS87qr8ltyy2pOXck8YIo3Ep
tJWewmeFebY9mP2hI0+RlbZ/oBhFJPUbebdjUlPlo8CPMbrJVF231fiVTMws
GLSkyoAgrMAvSQTqrLcZXBmhZ4pZdohMdrh8hKyGV1J3q15nzc5MHx1XsSPJ
zaPr/nZtgsY/IvlIUUcN6IxPSTGNGCg66DGyfdY9lDLdZKDFqaLHfug7KTWR
WW8MmX/Mz6UjO1BHd+R31VlFEC2ouR1uvCh6a7eN8GoThWvGopjOBdWlWBwe
q7h+Ud8my/nBbHxanHXffKtmApoznNmBoUTTbO4cc+GLlwOXejwAUjXzaXFP
aaLlRiToiymc2WJjDqxlKKfdBR+HgRsR6YtCNk7vVh/XFwLMxaJHzXQyh2N4
+UYxy/kpbCZ9RoJuvhVyAQRkVqGKfCcEFN2s9xO4PoTkXofM+FWlXYE4RxiL
bmne1KEeK0D85INyRsYdUIc3XLQTmTZr1RT0tjBAz4g7TowAtDhV/rNbBt2w
yffbmHpvSpimlTOA+r9Mjaui/APCgTpRarAE/pxNMX2+UM5VcHS6SrZO1ZKR
EAmEHA9paINCoZhjHo84Rru7QFoi0ZFWw6FG7y9EQfoFNdxq5cCm23mEAWyi
maFOoFORaKyHTVoo8ahSukqCKzuOJh+IJ8VvwpSyb1KvdSrPNTEcfPClpK4s
/vqb7FhmmLLy7D2n+4GwI8NhZTZtxkR0DPEMW8YigCOLebVCQEvsVGCNmQYU
cZlFeP41IZalxJeDvsMmyvDNoCsM+G3TECVUaybS/2AxCWOt4BXoGaPvk2lb
H0IO+v+26SXKYOapQ5T5eXnW6JsDsx2JF3U2zqgxC/CE6nt82Spovxe7R3I3
8T2HwxwKi+URpVcTFv7N3OzYwOrx2F1w7OdW91THhNAWMQEkGf/r2HDEM9ZE
XG6x8ovAhlG+ewTgjsfd7by+PCcoHLc+Xyo3sSHXwOIQE3YJ44HD0LK1o/L6
K7e6NItsYVPgHiQpIwXnTuvTnMCJol3NXOJZgS87/nL81ZU2rNxlZiCUUQj7
A/pQVLizZ0oW977ywPC6JgdxZFP+sTf5Ycv7x5tvfMllLPkPSD80OKdCmoKl
HZf6GiY1b2LXyPmX7ESG6aYvkcKLnXD6H2YTvc2Nxs7xXSeBYz5YaYjnRHXb
d6EMN1lEHLgBXu4mIsVzck0LJ7zWfd+hI1v/g9DH9DUH8kMPD8uojGSWc7A9
lxHVsUwMfL5UK7aThXnWtHO7vaQtsa+UPeG0P+vOqGi5ctf7AYMZ9kRdGT3U
nGpLgflZkjqU8cLeKG2Nt0fZ+hPWl3ZzMl4lBdmd/tBnD1TE4DZhLY8crQfP
qjA1VLcRp2b6AlqXCTdy36SRFmCU+hoq3c08WAM8Qv9Wd6vzp3QtdiSG1Dgp
UQwQoqQQsJmaiN+2F+D1rq3HS4mJDCv8vusPJYPHB71ir5Ju58+iDLF+k2Lb
J7wXBYpuyat92CJKEYFbODC2utkI5amNoY9xRmQRVn+ynra+qboXKfHMJdIx
MYAU6Yf7MtEKbRpLGWKwm+gn64Swem2pbwYWt7T8PvoGWdF9t9GXcYI+fLfK
c5A1ARTxdkZeQzFWtoNksfrLQHCMCA76xOe+06QlYt+8dFZq3iKORYqhdIrB
DV6KDkOhj3BXXs+Sr2V1UrbNc1xT22Ke45nxD/5pyz7z/TzMGMXQqRzWUX8N
DdBBxsPD9sjWeefQcxdEEwHdJoF9qKr9cDIQbv12Hf1wop7464TTEMEC2Ra3
Q9TRLwq3N+vEjZTrCCvuilaZouUD79WEwxc5+PFU3LpTYtSHSMJ3fCQIz4iQ
BXwMoeA0J7EahGFoSB30l+8DCz98pvyJHtu2zaPc9XAoi1RBvEZNDgmnqp0m
y4ukPSh6irOAxVtdVVTjG/t5e+ISQb4OM0Vp1KG5W0GxA9X1jQtpqx4WEjxE
1RFv1qlEELDwnUK3Eo67XD7o/ba6domvAKFuQOvopcmVlq0D4o+/vqfWjiOY
/u9MEXOuHB0fg/5ymH1sjVpChfgL2bi7pisUETu4wo091xL8Gfp/xEdMz+w6
24KCY6aTmyL42X8oh5Dhyb+7i/T6WcSjy4/5Pph4R5Pxh1ruf9mc74D5si1O
GFVW7peltM0DDMIkrGDB/MH6HBx/KHcLYQAx9ZkxN0Djw5VNihpI81CoDZbK
Tnr+k1Wj3d3JR+SQwOYyOoDYZ4bcwSncg3NWKGg0FslSK6/G1MAQLMMdjJuj
KG8PSBoEULCv4725otFB+OScZhEnR9aa64x0gINH2a9p0vHupwMAM3LS3tkN
GhOfE4v4Z6vB4vIU/szwKLp0kIwEU0TXiFbaSo4AtRGaOVs268NK76+GuEj3
x5KVviaN6FHvTMOmOIOz3WNJNYhkfo05lkwxnEqXJ5aoYUMGtwQ0ED4/5WaE
PlSzS4p20uCvLaCod3kSNXse87TkHy0QfOq9GvLUoGUGZnp5+h3tQA8ToGjU
29hYpuEIJFREJ3k/1HCqmQg445j3vV7pGuPUupaKtmN2UVlBaJMB0VOQ+FkI
oxR+jJxzkg48pvOuxRBChVaLlJntlfPDCqQJRQm1wGdMb+ZJ6yG1SKTzB8Lp
Eetm9Z9E2FnWG+Mgl/FHCKnEHdhcz10lrCC6peEbV2dvSdWcKpEi0hG0IdKA
aKwo+7rUn9IyYMuVoAI28JfYTh2edI56Cb/LPaDW4NXhHhTkX9ticOXQuzfA
9Ji9PDBg9PEov8Dnv1Q1oWAscwqITnWhh0TYM4SAEb84Talar/lwHTlHnrCB
g8elOG94vYWnSSThCJOaK/OWBcGyHGlP1/fuetcp5R1zkwa596L4IPlMRAaa
1X9KSZUsU6hIOnxossXIOVvIG9KyhWSMmt8R15TtICz6wqEc+ffrKYU7hiGL
5Ejg5M/478nYCP3LQYWILCEulozc59AC9fEYHmTU9kmDiGAZ9tDdHQKwN0pA
83IZQDOVDob3DvgHQBBh/aD30v/Tz1QGGIHMLrzuyHIPTVeRwW3d2zhH+cSZ
w0oE6qfQhSwUj8Vv+LFCALZ9VuVdBARHyDwM5YohPr8OFCGT+sdPbKQ6FAg+
51GpM4DjROwTqVVDawh7gl5v0Hwu33wyT2tZDyE5uX9+wbf6Vu9YwyhKks25
lGZMJtd/FHabz5c9KAPFIXVGkwJrmrzwk6mJn0kQYtDC8fJDOzkgRRRF9Qzp
xyXsZJ/CKFM4QPFh7puSHDSS0nAZemDsL/AYEK0P+8pgmUTIIgNr1rvtZ9ui
o3EzS9kr6yz/72Bdxta2Lt1ehJThM1Uhb7hULVTd0G1dTR2MddACkeFILPR6
B/ak7G2rURwbtL9gsxdT+9iXUYpZJR5S0+kMxygpnCUD+tJh28SRuZsiqf1G
hBU+0HTb+yM5//LSGVxWsQ5Rsgk8HRxCodnz/sKH9X3maHMcbbHBHsuusgrK
XKt+BGRrz5quO0myeCLGsEpXaCbjNiIOaakJddZMJZGY68833jgefTfssrPj
Hq9enqdq3nw0MOc7S015EraIcWcrxTiIIfd6oANxm3N+SYLSHTwqJn7qs4id
GDIKTIRoXwHxRxDKHQVPl5xhmWqI1WacI3kVGym5XgBBMzQhvF6pEuxZ5X4x
1feD2FpoPC9BhUY4uFkwLH6VRFH4kQ9KYY1x9S+pzAic3L66AEFuouXA+51C
PPNxQDggAxvW9S+8jFMmCrbuzWsmsX7qCCzno+BWoqlNf5fO0JY3a9YKvmWq
GeIBor+FoFOsKo+1HkuMXKSVTLdrqCMhqWkI7g9idvTVy9Ophkcgjf4ciQXP
b3r1udsNdKdkKMkgeLQOnl+nlz3QkpGFcDF2BPuBt0PN4dvKyt+++bZHpS1N
3yTwjpYbSb1RgCpymSoTJC9VhOY+FykCx3mXzyjwXa2LRSlu4uLWr0DlBxMh
e8F3tf02yk7I0MaCQnZpo0ELJxn3ASVn9G4N6/HSKKD2gVwzLZ+S4ZMYWEot
0pWtZTAAxm5HWN6W+wnpb1YCROzakwYlDtqiWFmHQBJIu+k6pCTRUSa27cpq
FO6snE7exkZP1JFj1oI7peX7h63SVf4rp2PlSGqS9LCuuHkcwCnZ6m0NTtzS
mqthFXFNTouTOm3o7T0b8tFaWZzc43naGV/x5LBJwOaaewwsIgXYbWF2CUjt
9HWZgJHCkbJQsQnCGrs1XrBhd2CZab0lwCy45IPbDPgV7h/wxqirG6Da+1zj
Z8O/6Jr8GsLLw9Nw4CrIANiWxNJ76SndWJ257uLOhvRKfxsSlCSziGEmvzzd
+Ba/wTyUuWv6Kq3XkjbM+0nPl1fgw3sQHXk3jMlOa4ac06fUFWXDpf972F7v
7HCWASQtmHZOjfvAuWAIG21fJ47xw5cu6yRrQOlahL+n1S8jUVOYIMmO0O+1
R+k3ZrfOgqB2agIV+NrwfV/yNvVV2VG0bpySF9bxS/Qqus5Ha+TSaei5UP/0
wkKc83/y7yuQ8M/8ixJS2ExPYGXAexEEsRxl6FfvVbr5BwqirfGxGkdMzK+l
6mdf1fy/uaiCzjsnHnTA8EjytnmPJuHlc3V6Dzg/PiwCKZviG5btAaIPndR7
TtXSgWG1KEtkSLoxei9ZPcznlhhkOwwA9MnMOnObRO5K8dvD4Of6P10OsSU3
05qejRsX7P0EGQr0Jt1nhsZWfSbD7KUPVP3yAVESrdswQPpgGwiw1RuAm3cg
PIxd7GN0UxYCxL5MS+eMy4GQI/IDyyyW+3KcLXCOwOZSEyyqONrxS3nZ4KzL
gcNBrEwihnrRT/zPIsb0gK1XNUt+rqesKJaaGXdfzMXy26PeSXw0pyB4wZN9
Fd3imbt0ggztbsh7acBGJutHUWLEYox7fpzOvAIpBilzLzq7WhcbqijXYvGo
WoOPPRWz+vj2rtQ+QTRMVEYB7stWpkJB2ThP7C+UOsI/IEq6DBR5yN8fa2q0
LM7OzVZObgRQ5abE8V/GvyGmz3OnXIH5x+sFqNhDYqRF9+ND/sXHZiPkz5t8
OfPiG7t73fhx6gpb4WKnSUcERuL1acHVMS2rkYf3AZ5q2OMx+8FHqGhRcDGR
CeIPtBN50OvDbHe3UGq1EhchSq+2mY3TDuZcZ2TkvOYeCsFrz8HojoROdkDQ
JSoa8zwNCbPY4SQfQWXoYyalXHgtBP9sRosPcug4NvKTGjvV1bq20TBrw5N8
IB7wpF3Uo/HywWI2/vraZ2Fgo3o8nfam3sVuyZKpXlynJxzrUnzS6qur71SM
3vDkdPOQip843aR7MCI9NrF6cSLoWtq4DUCSpjzFuAR9JP90HA929vJS1X/R
WNiKuuYFlMBJq8UYD6gwxeZM5cS88DATDvJmULd2lKFX8/pu6Xv89ukdZBSm
EFoZ/jrK4rW+zm+cyCA9stzbLVPomaybHum4QioMFc2RxtHa/Tx7tuTFT+Vy
W8BOypa9mSqYc+ulapQ1dyQLjuwwvt29tmOfjyh51gmQhQZwub2d8h1D205+
JHjZZM9dtGCil2RqOheh1hLnzmDpsl2YmY93SOdBZHIpcxOJb8Bm3L+mGh5y
OXb23qv1Nq2yfDQ1piS5Rbb1mInWYk1THkL5XaOtzHPNm5lfEb6a9wbN2QWw
smhGBr3QUjWju/difpouwOIoJsuxMA2lIWZrWT6S+QwDqe77rCZsZcZEwHFr
U+pcAlnCRhH1SavHbOmB8ln6cxieswV1bPspAf/blFj+jytgO8nrcKhBV+N/
Om0ZyAI4p5z/g965lJL9AMTfm603NLxRwd5hIUkuqZEdTCVCI7L4/8lKyimu
iKTL2v0OAzKrzBKhpJjtwH/WHmGRRwmtLde6Tunp1XEnEJdkwwk5Dtrj1A/4
VZCh1xl8i1eHAT2vSyN0UknHxg8jHre0HXsGufzH9y3AbptWbAURQKOk+48t
Aqnss2ReSo/sDLHYn7LxFlNm8T0V/7uWEabuIQTEY2XIuzq7ii6lwsgu20mA
GaVCovrkJQKIhlLkAHpXsqe0ptmFlvU8dL04RAuvRjZFOy/M9VOj/5ub87HG
ifhk7kU0tkU4uhSs4u8s9sSOrQyQf5O4eKUJsV3uyTdKJ3NycMgZsAtuirRv
r8i3WZW2FyrizsvS67j1ER2twwtaPHwnLCbEp4Xg/8TAUJ2mZ51u+2rpyM+D
SJ8lHx7UKCKcAJjixTV93mu/53XeYFbqMNqP7vxYVdexll6zIL3rZDZb/ie7
hwp57e0ZQ5PdsbE1L2XAy0Ruj4dKnRwuLLIkzXFyzKet+469pvNzFyJ07Qxi
uAf/ILQY6EbNl+V8vYk9tCtnnVkSy6QJ8zcsf/mV4YUjtPvnJRQt+ahlTX0U
JRBai6Ccr0ijqZfb4Bw3xVsYHnfhG0uHreUy2Qybr/W0iy1pjUZBDC8V6gfU
Q0BlI/2a+8o4j58MniG9XvBnUa7Iww9ZMHN/8NRyRvhtmNnjnm1m00u6gQyM
h4bShR7X/iv28KYDfdz9VinvbWs/KkL+RKYs2H1G2wRwEfNbHE+4j+Gi2vKT
spihT05XcbJulZY5oySUGVbQxWLe6FLYrYrAOqx2RHGqRWKrTyV95KFCoJ5m
YW4fN0bkB7izbpFvU3MvefQSn9LQI2nzQPq2XY9uQyaFC0f4+XrAJeQzvp2L
MUG8G4/DR1EgAowKVsGGZ8O+tsWeL1V1L6YPM9ycLf3muJPu0d2ZCPwOqdOk
mOFnB8wsnHGOezi+CvPtzDpudULSraSwKZuE1P+3qQC/rH+Qth2Mp2qNfzxa
GgYHZWv50HYnikMrl5ZLvayrP+qC85HA+8dKg09R7Oh6bklRi3NEl3n1HIgh
2At9WqDWyJ06N2HK+BBhwlB2A4AEuPTIhc787d/64JC56lJycVxR0Hc+NG5R
pAxcbBEYRrSnPua7fyUKSoDKu1ZhT5EbN9XPnHketi5xZGfeZoN5VwEBYAXh
xIrSRtVg854TYkDHgvFWhw1cvZ9nF7NYt9pkfl+T/ddpxPm1u0E3oaZTYtqD
YP9vCwkYr8Lv1b9aF2r1Hax4FNxFwQeOD5epHx1AjPo4+iLLjHHZLK1CKSIT
G6g6DVL6+2DG60gjAqgboCL+wkOoPEY1N8egw9U90Xd8eV+2glIZXAm17yYi
KKcb2grw0Jkvm3H2eVVCsT//hGGwARfHR85Duy2QOYl1ydV1pkSb01KxQ+Ho
m/feOeGPrEDk02iUOx2QhQZL6IqiJ3ZHjoe/PpEm5CHSTUGnBc8BFVNyEZzd
FHSkUPccN8NzqNgnZj+sPP3XRuXdU81PmKhbeYwmAbN7C5x0dgJmvYBeZcUH
6YPl8sXOYuKMz6f4FtT97So+dbLPKTJ2R136iqECzndO0PlOztzEzce+e27h
yq329eoBpZsk/glbn8xxuio8ntCAnv5XhBu5SYQc463rOO6xzjn1CrVASJo6
kIPNSc1Cg5Fh7Q5P4oOCEHgHcLcRcikzesimJtWg3xFI2+/WkBIy25ZNHUqw
9hwr6Ju5Jf6BS7CeJ4++DMNrGN1GRBX3IJVIgQ/Zk3upBSn9JolC4lcbOV/E
HuyqflWpdfmjAu0ypDbOiBMoFu40XntXXw8njR47fxFQBV7jc2dyjsmrnz86
OZIB7wsUWDUIo7DMecdTP7KP3ZU7oWHSHlY1SD/1W16AmCY9yyJC9TOXswKC
PAjPjLRUKOEhqKGT5N4El+dyqm2BchaUoqjpjeSex/I6NEg7RaYW/4G+TRIw
5ZQqLDUp/feo3oEmg5vyP6xT2GR3YFOZ68wpY1X06VlihNrwqtjxe6hjapTs
wq9AfDkDP8qDuQu+3MLwLMIXwnHo7s867Dl3m4EOUXKtnrd478e6ij9MdDwP
P5DihNAuiNAJyXc/0TiaGYRZr07J+nn8PkYdO0GWl2/xlLjAX6srVpbixsoG
XveI59hOkgktwWbXr/k3sk8YVHTrZOJl/x6Bb+WqjRbZj9VvfpyunQ+103O3
CQRW7EE27PZ13L/1MpaxHHcZx0bsJ1IkgTGTlEC4PXcZAFI2cLqmlhkdqBr/
2FrdT1KKqA2x4mBPq7fV+0DIZGMJg1G2aHFhVftX3hIXm88OC4owBfTLtTqb
OUOObS+7WDhzB1A6c9rjHb7ByXJRRrIWe/BDyudnv3aZBRrI2ChBhRAl+eit
GIQvA1XVMBbtxO2ARxGKrmbab8GaP1f+D7tgJM+kxltn1XvykuUuClI/Am9w
ut7DCW5WHZaKaxX1R5gMRXGYz+0kEaD8qoT6PKLhYr1VSRruJGb+kyWuDgl1
5la4cIXU+V3jn2j/ocG4QwI96RmRL2y+JvWYuGozn1Gd/yWVwPgjiUFgkCbH
zh8U0Znl4J3XkP3CHqZWTPDU5cjyXJjZyOKuWLibJ0YDk7H33kFEh4EX2GTk
EbY62kz+N3QsnHnL575zensgAlmSgXCNFxwuxXwIbWnhAr/h6M3BT/10gIGs
kOIuj0tAHFkJ11WMEyMe1KK8yRLJDqDDVDl+gfGla1QufOX7YODa6e8J+wET
vBjK/Vm1RJCyPtwZ4z3MT6s+PGgZmh5MfOor2Vak7RQXCSIRMeBqExrw+4s6
wWbocc88PV1H+serJmcT7sxEYGpWBwu3QTLDV015GsBQYDKK4egVLSVnfm6C
JRfBUnVnFYmc6F2FQfBDIlCNapd7UoRlkQek/df4FNboW5AK7LBl6F4uwN8j
XaR/F8PF4+X1lt9rx8p0YYKij8HJNhr4jjYC7nCrlPg0UDmg3qGMsAsA4tC1
cF8Montk74KiTyT1M9CHt/417zEzRXQ09TTlVr+n3OU6gJfqN+30p3/lNbBQ
NiL3gNeKZMs7j20ViqIMT8DF4O4wQb7TNxvix11q7XQMkpXMDQSbwLHYF6+y
LB7fo018WW3uEIDRiJVXzMOvQMnnaqrp7rCrFywOkmEx4CVDBvfWjoZDVI1L
ifSKgECOAfeD7A+RDeDVqrdcoh5REY43UsE9Vd/VAHD/XkwbKPbJuC7z5ecx
veALPjSL1P3D3FP4tkHMB33XzVl6JzNkL82Y0avNOZKmBjZdnYvqlOpoNvDN
3ODMcKLqlKsdNrAQfiD/zIv1hHwEhSdneaoQADaFrRvGJPqyWKrDtVD4+xdm
55G2tu9jtOtHTbcorkCU5f4St4CbC/Jyegch/+EebyeE6O60UcX0sF66cRUP
VwF3Q4D8k2gzHRHAUbIrbdp0NT9+4JoFe4b/eSf5SN/MwDsXmoCh2VTRsHzs
sY7NPd0dKILmnYanUpZhBba04TjndA/wuHMN8hKJ7abDDKw5ehymBp1TaLJV
L0WKfFLHdzsZMbme7Ih3XVlShhzo1yMX1UTx5BkAXjUD5P9N5d/dQRsngx1v
bbg5vgmceIpb0nHv9tH0sydN189g+8a+8C/4zngvZaabBO08qWmI/G86EUGh
97U2guwR0Ki1QPXUVY4n3Fmm/NLS7UqSHC5whpKQi031RFkNueRYruWgghtX
50sPBUlqbsq42FZlPcXEEqdi+gOEl89q8Lh2dOJ6RD90W9NWsLmhHVn4n0YW
7C2+6BgPWpfozGSTmt1/4S+IW9hqD/lOcB0ZQ0lVkxndITEBxBX4pfchWi+R
qJcgY2dzzLcH1xSiI5I5tiuIGvMWt/qZkGR1NV1JZZQL3IXorgy7AwVyYPNh
P538bOALz0CNDr6UaMDz36+25uM4DEOxyFOx8HLJ5CN/ZcXjZTyThDllROMS
zc15bdV9noQTVJCDEjpkSVybslJH9NELd/5HMv98QDtkfm6Sn4BeKRdT1Bih
vUEduE2j5ANfVfsnJLbPci76UC7m2qTmjb5XN5N9BBDXTZp98H7km48oHWTQ
s0UK/4dUhV6bbqmrVR12aUMlCf/8+DYf82ux5FjnjyLlt5tN0pGYkXai8DZ/
ZCazqs4C/j2a3G5L69zai9AUYRbTahSuc9TSViVuL8oO9PaFou56HNXekjIM
HdWCY9u0C9rx8HngXsk2pUebj3dBq3oa91f6cJTC+bp/TRtfXEzWanQ3kFdM
qf2Hy1zBuxUNeeAq2AubBtnSlJqR/uFOEmTAH3pHHfRiArI9XLhP9Bqtn2zr
9mXHhsW1ka8ykyddi+1IcYqZWZpYXghBhw+YHeiLLxGb2jwOkrweM7Ahmt/W
rjPKdIHG0dbV6w082qndIESRGm1u7cj6XRK0JU677u4GBshFLTy3vZvFG9eu
yVkrOkTTvSO40Gu+eP+2SaWMkceKMHp3MlgBGojTMH2WOK/neih9AFfaSI4i
RGjCAqKp4O+JG+Lkcl1Tc3Y8XzNd/4NMEzqIjCZUr0t/7ZdTptAsX1pjqi66
dryzrdoMp9nY4xALaMvSIoAWM3TmflF9vYH98rKPczXRXIGYmHEZ8bhlp7JX
buhgMushD3vvvkNr9Br+YZjdEkaUxvy1b7MPF3xIbcVWHFM9rvDkWUYLYGc5
qBdvEvlmoUxGu+LN6yn1fpNRjvHie+FErh3mOY/rLS4DwSQjLt2pwS8+q7AB
a+nJekXeEqP2OsuoC7usVevraX4I9HTEEvPCUO5w4kVHTv9cknJ9MxFnUURJ
iqt1z/5k+NYm9OQ9sqYlbTe4tx4yRBdj1Sq85IR6CxjbVTo1LzI/Crq3/LCz
JeuGoMXMqhyDNNOFKPrXotEI5hea3R9/cX4sCWUW7jmJNS4cqM4usthvForr
9U5TdEwI1CmRhKULujkhMvwaFjFlp45EgpKseGZ0tdAcmGnykQKb/urxsvJL
T166gyOwob6c5FnDVfP6sy1si2Td1vQmveTr5pUM9xfudCjhbY5iaKwWzpXc
24EcuP7jrBiyfEPK8EfZZYhqwDS2fYptYuQa82/WByvcBNOyIC0HsbF581aw
gCxhMpOcfyOtKb9PVGabmlstDT26OfPQnYQRg0qfQNfe24obHXUOEXcgB4Lo
CJYGijrYiFCIbwPPwwIAhCnTed+8vTD5feDH7XwaP2mPZdLy1d9nE8tHvKAe
uuHjCwmTSDBaFQVQlSAVoegjzb4W2giUEagwk1yC8kq86QXVyZ2DDGvZROfn
nDxnsYPgKKFlH/lJN1zfSokCwlkxchmBLS8JXoyA4w27BpnCoVXXi03TDCik
o4BKMIWQzmtJLO9Hm1fOiyxTut55ROhooj+0JDIm7Cvt2ExwLh0JKb1u9WlC
sGV7Ar/Qrj6UuOOP7dSERETIoudYEwWCscIYebVejmOmlb316HCGCr2OqM2r
MVaLyxe2bwEP8mi2o6qCaohuM+nwZmCdaKiYNuDpnk+zWT/c4aoreKo30Y33
q13enFXc4nI6Jr2xSBgrDi4jYosOY+WzMcFV8YXN8nP92L+v0wfPqeKfOPU/
VfVCnjrbPIu1AOCEnpUSResab1+q4AWfr1SE3/ZQ4lHGAul9R3cub4OQPlTm
d7CDpyyRqKFS4uoE3L8NiJu8GMpOY7ND2qA6CpikMc7ghd5pUsirhtBBIpeC
lqBTopSbkLiKw3c11ip0r+T+na8lElucfyYDNgPJp3cSQX8JtzELwojOrv95
ZYqggA9TR15tz+SgoP6QHBji+CaZF16Y/EqvQGfr8XIneS0SczobfJ5eblG1
yP25eEPpKXDfCMD18thHkpqPe+M/26xkfMQyBjfgFHhGJuqdSNlXvkZx2vFX
oQo3U0IIGcdKOseeO4mgsxPfIyj+bLSCsszk5dCsmPONRAdNuyeVz71gNTdi
7roTLN2IRDw0dLuTlZ+2/QEt+xtdYECQ1avED6ar4y9cx6BA6MhhuySGTDnD
FogexBM8mxdoeJlIVRESDDTjXCAnEWJywWHgZ/iG2YytyP8zr7bqdxyAEFZQ
3qV+dlnYTeMK+YYfZcyblkuzXnH28eawdyyWuB6Kb4VRobR7pn/usy9ZzMrg
2HoFBAmhttrYECn2qXkCNyio3en8Cl878o2B2WUYh7KxXiyGnpegMAMkSQ4f
T4OBTQ5Vm617IkU+2oDASOi0LRd/oAbE9347HhIYDyz2ZKPFA/LQqgrbO7h2
rePp0R4KvYPE/rc6M8CXCOcmtoBW8jDzhkG0DWvEv1kxGb6ci5J0oIUeqRas
sn/xW5W9O33e6lCe5gi9+gZwJJV6PPo1J+fPOCwibpgJW9uEFcpYF4FyldDQ
2sR+BQzJkWM6mcLamg1YpYnPZFgkVkzTRzX5+JqSjnTseF0J3wYy0OC1lEGG
6kyn7xfwfuKPg8+U+qm4DOJpEej48QtfHkNs38sLZq9wFVyTqwNSbedvn8RE
A1wZvOWzRW0jsap3/11T+5K5u1NqSHoWGrApIw4jtSKASi9+3/oUfisWdsqo
n2SsJWd0cLrGEFG8sgYFyA5h0/zhN4npOQBshqDGzQm83YB+85SlYlTvF586
EVbtSXFtaQEeT26qJ43kwL2fUt8IB717bX5HFM38HnVISO6UW9CfOoF+wckA
s5QJdja1DaS+SkpxAgr48jdH/6MO3asLP5fCvZQGXagjU+0ziiN+LnJdM2Zh
YAgUPTEmMmSlFPSm5a3fFEr0bpSvBEQRiNBTANoTNSfRw9/yAJzm2s/WZe1V
rwzTX7X5KS1G0BKXM1+GmyYLhVByM9mrdDSodIUMYn0ybsgJDfRHRmTWnhqH
qQ0zsIrjD5P2bqCKElG3G4OZfE2zlHVH1tJIvabQYsvRp7QT7SX8r76DFuvm
sQ+ZORoUVg/Ry1wD1qUcIF7GU5a2g8vfDvU6KE3PW8dTrDvKokQDKfaEs9nd
kg1JWXCZ0KkkOS3Iv/N77SnBMGa9g37j9yTxUvYxRWQlJnC0tUDTVno6D7Ci
ZnvIezGkC/90otx9p1D3lBDVpdIdeBCBDFbPk/gjyOxHs6uWdRBV8BXSjdB3
KhD+umE3iCE37724WhElFsKpPz9skRXYv44g5oAZn9BCufWAPu3I+ViIuasV
8CghXcFXmWoDY/Zli8B3xHD++X8iAHVJdhzKujn45teznCJUWm3J4qQc/lVH
yoRslqvPfH16zta+eCq588pKMvExmipnzYNIQa+sGTrZ4R19ZQVXGzYCQZTm
NKeXECVZGxz1qoCOmJElOJRKbsWKjrfh9GuZGqnG/lWkO5yhxFOAuwp+Dmzm
beJGQnjH9qytUrZdhFrMeHsS6DFr5LjKMUHDsb8JZhRvrBmcTKy12GsT7cY+
fiYCyugCpDKXYsNUFXkQApm4JYCoef7tNl5J03prbZ7brYQbW1ORooAqFjqL
beeijkpjeTuwPgMVA1HtsIgv9JeUGoW9B5oGqf9vBhbWJQjFS8MM8+4x3cpW
ytua5vHxGx6pBnM8PG2LwJ4w2on2E8hwnmHKnQniVK1Pin0twe0armJ1i0Pp
sEkit6G3CHofwBsd0tfx7XQbGCfDw6Yj3dv1VOmpmPAei6QeU6JWXQRh8j3O
IFybX1G27bruDqOAin+sZ24tCYV87lWtOVJLzc72lkQpCekHLlNG+/hNQyXU
CV3EAhHZxF/PcaRfEmP9AG/Iag0U5wOJHBFz53ZQGKhHEb9wVJdp9PQQ/kU4
xIQeAuqS7b263iCteDQUlym0k0XPOgqq/VzNAQfEGAtoPGSxFlKkhXyUPAqw
ynX5f8jiFAybffQmWaG5xP93HLVcKPAqNCPW+I+nFfGp/BU1Af9bVhWU+hLB
qaEX80iz0Q/2x1HHOfFt1PE58VmZDJk/t64BRZJIhnljojyJBgGDrAXLwXU3
ryfHlHLYVMN+itCUJxSBRdny3kvMW7INfEOhJBL/TKbz5lCdyOwasTNYPDn+
MWekjeXe8eshfbFZQiwIogul9xnHaqOTth9WbCY3HIVCHHIWRD08WuuE7uqn
yG+0n75Se4oagTEs54SLzhqHSSgnnvNuQ9Haus0dRRFJGKNHWdrqoE6KscoT
8QvV9JpVIONbWUr+fm1BWafAwsOoLKYZHpppPA1Ersdie4+y9MRQKwSUKaKm
HbTVkv8XYLOUVUXDjuq4jXaw1+77iFt8+QuRHRzu4V8jRNYvZk15OkR2u0FF
jacBwAwkzbqfEdYO3lIKaGW3I9kuKkg/VVkgo+1tdI+9Mhi/7hwrRJTgWDfz
ho4w/uXHk2/OmxZbSGLAmlnpfzsrn99E0A3rfJaAb4ijtPg8XZmzH+SbByw/
gxKq6xl+x0IrkhWhrzq6rk/dvUt0Fp4s5RVSJcTL/4MeAqPdom3M0gnC0k2I
tajUv399+QzJ9UrWPAyOA5oZvYWr9PJkBTNF/VRQR/Q/hwdAQrsi3Znkh07e
y+ZGKHcZ5V5Dls3e8hXvWbrchYTBwtxC9Tyd7gkETlZTHHlgWAomj6JtG+R8
3cO9TbveyznQzJQW29ceEZ4DyG8KaMTZ7x8dprGtpFIsUhxOFgK+T16r8cXl
W5+2wGuQ0FtZK8OhGgw1cAY9n78+MVOk8Qku9hYxoiUdwz/ukEu+z6quJjNW
wI6OiK5NUmetr3y3ZgyjLTIgEIiyYrUdP9XkeoVj9cxvjhet5hA4TP2EgdK/
yCP8b6W8O2EHRST9VZ9UkkdHbVCMunU/PFNz9sW7l0X8zEVZM8Od9+CYi4tP
TIGNVGKJbLHb5P2bgBpX9Ss5syInbSo3fvJlhAw9HwDdAMrjPrCE56eQyRoz
ineuZRu8nAAkQaww0k99BXMZpzn/xFTmDfZ36xstyukZDIH9vkWXVDu6dIlK
sw3+3VU3x8Ys5wvnBOeOSCau8uroivhT62rx7LvvO+zbxG0WHzmtlJLeh4hR
Afa1hEbS6TonMU26tSPQ4yncoU1jinVL2eBUMcyA8x+QRaaCtppeIILQ4xH6
JMysWjKjpcd9VUBMBV9rdA2b0aSV/kF8fF13aCFrWz6ZtDxXaf+BXXCJ02G6
cNP233/TYDb9Elsc0reASBRxmSNHZnq4sGv0+DWA6eDGemjIDyzwMi1JCXHU
4wIVqCMrvxA9xCNQr1bvZRvLtkVn9TIU4miMN5ubORtz1/DunR0rw2ff3qOA
cu2/Ml01ERH0oaIBtHE1FfnomjtaZenH9fB7dLW3sGvDWHQH+8pfUUwQlWsZ
PuRJRDITT52Yq6+v90GCntsTQKE+OrFmTPDUkS0fYQVDSSKZpIWDoVLIPkQU
KgQHXQz3VBJt03GNhyyr/r+K2Zu0pFRZOBy9f6yYzILEln1HpqGWIzmG4WIq
redzlxiv442t3SyE9e5pWpw0Ns8vCPAH9h/3ZIZPu4CNGgfN8rNXtJyvqsFH
PJshlEN7kKFiXNwTl2gwAeoGVgwWcPY2PUPd7RnjTMKS0wJdzMWIWQj7x3pj
fNEz28l3cCSxIeNiBLj6vvlcrzdwMyZoAI/DjYj7OWAdQdmk6RaiAETh67b4
hLYUQJX9GjBwt/7pl/APhub4IBn6IyYU3Qvp8DCi4jT6Bch5rZC76Ef59af+
9nBj2MMo8hlKpr/mACFLLpTpSNYoNc5ANBvyApE5A6TWtN30hIkh1JXdbBwd
i18ROz5M/zx6iJRfRHzkijFxvxs6GYIYFByXsmU9zklPbpyj8A8NwOKZ6H0i
rPX36DFJrR9cA7yIqvYL77Cjhn8RzdL3f2VQvcJ4tdAKjymllGuXm2h1C+Y6
UXwqFAkiX8QEZwiA7Z7Y4uCEe9Z3YQDuisaedlYR1dQdNvzHXUgWJBDJopUc
0HvwV6YKp2P3jXcuoZQ7xG1pfFP3BvyMDWrBhUpJhprzztyuPOYC/iOZlQqs
vW5ow3y+TtmhaLUDrxm3riBXRQxVUQHMJEVSo5VvWSoq29rVpwc0bKODiCQr
tzRICLSojkIyv4ixt5yXEDkpOAV8BxPF57Eydkw5ccY9nyg09jYD5Uglkydd
iDV2+cAswQXpdFU5sEQfCVSfNKzwdJRCjO5hNJZTAefwuzcbsyR+M2Td5M0B
bADHJppWRmOXS92IiKmLShmYjQmQckUgK24Ekcd68dGNDqKGSvgZ7Ob6ABvE
O3Sy0tkB45GOjQbr58mvuH2w8DdwvA/L6/YtdvmLlMEp0RjltV2hRqgJyE+C
SBADdCuQh7FaQda6AWxPflkmmx+H/M9TzzZbPvC4jUZgLMrmSOQnY0rHjE5Y
a0r4uX7EOwvTnEpBjGyq3GJWb5ZXDpoZBCsx0wfTy+DhM8Q6jERy6vS0ix3W
jVt6XiA6TuzuUfz1JsYHz90NSmIDm1fDhR2hAY1m3VVisoOoFnWtoa6tdM2E
2llz9QL6h3QutLOd4mYsWOw5dtMMKDSPHqMqDmFvUUMOZ9y3cfzrjsjBfqDM
YTwQtALyvGfW9Iz4ooUCnWUGwb8xAefIvmRIdY3MBcC9j/vVWAa7JfvY/eLm
hnvP4XxYxEicG/e/BI8ZsF9BHbcs+3Ij18ur5QMo+UGeGYVtDlkJV/i2oSw/
pbBZBpDnxV/GURY7bOYI7On5+FhdH/x7TJY+R3hcxcTE+iv26hGkSWV6w58v
B0Z3Daiiz+PdybIHh+y7UKTV+PkooExwvwiG0hPVzVPiQic7s5TJL8o6dMQO
GNnUw/ooSjx53N6b2kgjkQGphxIIulPbpTBXfj5WSKYK1mToWerhH4er4DMV
9F4A/0mZXYfSbdsfKes9DKKiX3OkOXhc/HF3KnFngwFKpawAlesEI3bW9H0G
dIfDby0A6HuLSh7kopXEUAafx6BmUn2W+eq7uh23wpii3xwd7/F+lF8hTnIx
tL2GfT6LgUVa6Kc0f3mKTc+lCCUwHFSATDMFHpovwCpelwIFAswP4rKRzQfc
OuWvR70bsf2Mmikbbt5cHltn7YpjuEp0372ztprUVe2yV0w72A/zG7qhD6qV
HO6rK2bQ3ESCfVocCKlP8Ani4jrCZ6a9gQi8qC2pKIwYtIqdjJmmyx1+hXpL
SOSoK6VxAAEwj/fiIE1HRXzosP511PWnFBJjn/SmsGP40B9LeZ/66IluQRWa
9q219MyaXYfi/ngcbm8w9g0k0jcfm3XK1Zp/FH0hmH9XKw+Y7d8BUSXWzEFv
TouT64lQYlB2xvGawhgejfuPfwrEU+eGG1bl60HdTgSYIX8/bMabUYJAKdxG
g7F2gyFQ1pyOgZ6j9rGzvLB7o0etE0gc4xZvHAvnwNtvtQ265cQwYKg7lWz4
XcKIbBkdTjkwwz8MiO87N66GO289MOSkKjHCMkpu9tLLfXk+K4BqP9lnaPIA
HqHdSbkuQ5COEvBc7EXABZiudydCsWp9PJtbDx41rWRdMHt4nmaBJKOGRAUl
TzZQIoi+qzT+sQyQBvpVTJz+Qt6ZKRvkZeFIOt93xU1zP2WHAw1jVFFSZpLO
svnSP45cC1YR8cp9lplVhnLkTme5+iyh6F7dWrU2I00U/a+uFXGHdINmLjkE
DNGSJ7DDa+QnHlRxyYMLelVIxZbxvUbZ7qkpMJHRLD5PS9g7IhpoVbPR2yUi
zwYrppNJvxjVgTqJPM/87KMOcw7jQgjIDV36bjrFZHJeK9rbmLdK9rPHi8Yw
BsPN+0v1UsuyVMI2dW+AZkCq/QgB7VUkppiKET4tN11mXBWpQMYYhuZXslCD
ZJZ1xbuxnOaZA/u0TIZApqV5RgZXIh+w8wr9qHFhgVodk43atyjmaNFvSjUX
ISrFb7y6Q5V6gBNGMfpyNTJbfI9vlWdX8d3rX13To2/JLPeBVseDCfWrjivO
RddeYZzdD/vY8b9kzN9xalsljkwmDVytvdIlh7RsEMyq3+rSyBOqkBRShxDT
FIMNGo+gpoy8bC9G30iznld26/Sngaw5z8pZ0xo9qTQ8+eziZyhykAGCoimH
CYV2OHVjyhraqmuL3H0//03MHPKpTT3pAhae7mVGOw6aYXoUIlkbcmEbxMRc
2+5o7rMHDvLs/AGVpjDMX4coVS8QSKWB7hdb8FZdMONEmfsevSwjZSdwVh/d
XqiPcB1HKOMoxUb3CRdMd6uuX9yTkEAt5l3wZsREQBXOtBXQLLzNaJ2fbsTE
xOrOrvyXKcTmM6RTh+sn/jXFM5hWuUbXHqXJdnoOMSuLZ2iJ2eBnXU8jRySH
cBDBl0Ov7qo2Km8mGv7YFi/bhtu5JvjrZJ8WEnw6hmBSjxAa7i35IMtamKNw
0ziCmfJUFATyfHBTtG+ZbXzHVwgDZbMGVOQRF5nQ2FIQlExWk9/6CtmKDApM
TZ3syxSTAjCn10mfsFv5YbPo+/+xAsPv5XbSPJgT/y72EWHi5Dbz7u+gK7EF
GHD1BMW0kxH25sVJB/IQH1P4kU76QDQJ+P+alfOl3wCwidXX1r69HofyekZo
I/0H6Qg71JksksuRtBHtJfnhlemu2IHa4Wrds0dVgNTCC3AcAdmymZ5uq8c2
e6vDvixdjMAbNGs4sLovyWYaXk51O/q+oWkz9bSvtZvxl3GmJ5Xs0k0dYAIg
U0ILnzwF3Lp9cvllJCNvIIzlxaBDEJ9Lts2zP0hY5qruc2J1P63rovNWrzSk
0/9FSKBjNIv84N1vka9n7R231bUW6mdIKYXkLiwus7ScYSXRMq0ufMTH1m6v
1YBg5+IBRm4hAs0R12f4M9TqGbtHSmcIbSn/k/CD2dTF9ThulJP6uMjTI81a
4XPT6yNO3/W2QzzBTQ0Td6H8z6IaAhU1rAJUmEjjOy2vY5JFSPQcvExX8Z9m
74RvhPXdVMB3SIg8NfECqQtAtK+igJUXoFQQXsLaeIA+G9y5e7ayiqYn8sdz
tQM1Pfs5op6427HZaUqivx542XdE9rHIHSulhn1QybAKyf9KrX+tkjO4QIKX
xH8X4Ud+SowNjXbVXdzx0RztLjo2NpuYJbKp9dJ56FHPJzJWkieuqxyrtjG2
BYKhk5AJQ6Z36AG2BSv4Dz25aLZ4IU3ObP959BtXT5kkko5ab6leMJleVXIS
/p02f9XYIGPHB1+srBlAZx4DqwMWCUzE3j0AYuj7Lxyr11FcswgKQlN0MWQ9
OHreKskfO++yK71DgmVAvqvWLoslkttwRrixoR5moPwKy2SqbusAvsjvXxYn
5la/9vtGbS3BBTV4H2YaGLh1wuchFsnAOlQqvInZVA0rS5iVyKAhaqMsaa7f
O5ZLaMxbJFMfrbuvUL2UjRDoPXmaqhMBLuba27fkWoyg4UbdmGq6XtGWCjHo
qMsDjpYac9AoQ6j6+1iVi6geKWu1Kwe0stpCCTjiEhPAtolHKWeQ95Wz/0Br
isTKNnfyiRioAd9lzi3GpUd74JkVTXIOqXf1blN5/6pUTYYz8O0/Yn6Wbhii
bFkascZK7grTDt9U2/bvn0HNdq8tjcpnW5Enki3KN1LBIPrxqT2nm3HunFnw
Gd9LwhweJ3+/cjTrty2XqOybCChZxMZuKdjY83u0UdVq86HdGE/WDJJCBgVA
R1Wf489IItfITJRrm0LT9U3XG1YtLYxsbhzZOWkzvZmJOampv+pt8Lfdo3vS
MKdK6RQZbia5/LQVKifWwRxyIKskMEpdufFFDVxIwJIlnP4Gks5sELY4qdAD
Fbf2T36O0wRMTk1yRAKpcruM19C49kKgNH/TfPzTVi/fPU1x40ul4o4/QCxs
7K68cfUx4TFR0rk+Z5yEcXlL8HBSnpnpGMgjCXd4Sw3CxMaRunDbphN0X49+
WA+TCTJD85brc7678B0RGCjfXwl2XXhwGky+O3xlb/vXsS+2FydxO2CiWFDu
faLGLsIaPSeyJxs8HrDRDU9alit0pzv+scdkrxz2nu6v1O1FfIFU8MAsRcGN
CR8oKhKz02zKzP8yzEH7yjl2Pu+UAegi/BiyEp4x7YbaDwmRg8JyorI2Koen
Qt0ZeUWH8QRV9LCxholkoJR82dGoyWlKYfWGs69tOYDLVuPc7Fkkdmf3qMt9
CYDt9X1/JdTZv0XeX6BsT0KB17pVMAcIHLZWxT+tCNSGx40N5nRyXkpRlnpJ
HocbyfmgB4LUX0LCnbTPZpQ0aKvR4sfk5BN7Ny67sXzQkJk2lbmV7rjV1ZAZ
ApWwcOLClnP6FMmf8FwzDOichsbOgjj+Z026kJxnzZet8esuS9lfPKOef67x
FGR7Khk27QimuKLyurFa8fPC+yxRQoIEoQ8z/e8zzp5mkhf6wnMb6fBxK8kN
HvPooaPaSM1zb5peP9Tz6V4cdroDG+58akd6wi26PTTKmVHdWaTj8+nKgAMv
qLV9bG7fKNshmrtoOZYR8V5TQfRSYbr0WMjYdjLxO4Phs6VS6InODxmGeLCM
U+m2U6GLFj9J6WO0p3EJv5k0+o/3Vl0kin/q3M49ycar0EziKSItvhplV6NU
dS+FR/HZ+rC7SysdBh9SMFJA+5HC9tiOs14vBW4Wdq+kgC58PrxurNGYQoH6
Atbw5Oixp6d6ViC/quKSsgfBMiXiMz082pM69rAKqHNqrhydvi2ZjJRb9Shd
4aIz/47WdZ2DI4QIMtnOdwwznDpawgR+TWQFqqC7U+qTjTZfpPeXEMnKx89m
3VXdIVcD3nJe5qbaDZBgnUxDZ8/X1g2ZrXrEgiFxAvBKz37jN4eOd7DBUTZK
bp2mT8s3xUfFvV/Ja1RTyd1ABz5ByMbsMnWDn7OFKF0ILmLK0iE8oIWPpJ9e
8kpB0WUNRMghMn1AVGOtvhjNB8+bYsk3+M4U9gh32HoUBg1g4We7YQ4I5uA6
5Urnsl9WiBpAivL9MbeAIBisoU3LhIUYvah0LcIpQmWMiEiVi0EfeVrsJxaD
661lpUKafEQPK+20/c2NJjjtuPuD0oPxw4HlLq+6EUYBs0VcOKaPNmWlT9/K
b5wY5A4i+rEgwx8Pd7Gj4Tg1bMqYr7RTjAWbVEVNqwhD5ydVdcuJ02AMm4zm
S+GA3AUPJkPA70mQZAuaPz0Q0PXZAXVbKqVtkAHaW6U5sk7Rg9H+w2gQtUND
jDuIf4ngjIohcPq1OyqvXUMeyVWdPHs0FaA56nuDrWvNJ1B+QGQxSqVjQYKJ
3dqZ0Z+oCgPXWH7XAtEEoQo12yDelBhOb6u+ch5ocoPSLWIfsaRSJi8B9XJi
wgBkh4K7LOLEZWMXAIpMzaJxtI517d05anMpH8Avz3+Ifiaq9n2um9C1+ne1
3+69yEc+Zchp6mRKaVlB6mMZ2jbPD8vlPcL+LmEnlCMw/74+VhQsyp6kQLbl
0Mr/ipT0DtAUONKpuee9WJB3s7c2l3I+4gxXjomNuT2PQBWDPg58b3wC83lX
xd02+kZSnfe2P4jX324aEZL27QdcHrbTxtvMEEwBPLX4HItZhwhVWUTxZ/sa
1rV3ai7j87XZIJu0JoaZsYDfvRe+UJpXrCnglyi7yVE2L1jZjyAdTSBCUd0e
vhcnoGnPAiNNFsMaNbS2fx6fV1lU+jS4dVHtNAd1hYjtwd8AW6D+R3O8Xhiz
bia/sat5UemvN/3SXHFgvzY1GZPCkV4b3uBCitQPUGUnuYALCqWbnl2RXIAL
SxbvzmSjG/DKXnE57+DSz32uxQIcAsc/qhXHPfarTTXvIUlBG1Jp+iHhBaLP
Ajpuqcsr1ffq/ChDIX3p1lsv7Ieg35yqSbDr3OnxyVWzDlLr6bfdmGCfWjPV
x+x/iNNauw6xu5EysHH2Tziv0Wv4e9YDOX22qNMSVZ2RdDeDoUcfmHZ7b1lQ
Rw817nkETyt6+YGHkSKDEKTXY8Yqxj7XOZdcLVBlMcz60cS+M9JjCluBEVGk
w2GCyqHk0uvmbmGUYyzR5i2ljqbcLCEtNYP/1rzH+kmihN68Atx2zTK6I4Bs
bdG+LIZWKExVnCuSRs50pvUBgYxQWDqg2yK2EllDC+143JDsuDvhdVBX77w+
ct6bfp1B1fxU20VDh2teVnFcTiMHQXSGPgPYpRYroTqjhQg2W+uP0u52Jsmw
IJq/gyJl4QIB7l72ye4zAbQ7CKlzpS26pujepfiQ5KQwYr0Ict/N68ga7Gvm
702ut7Vqd/qpaU481JV2IHuPbRXkpAnFvnPfWFJFjMHofAksL6IscLw9wS3N
TL3JQMxI3aM3KoaSq8P00j/O9yK13+iFgFmkpz1VkonGqomvfsvzwlGundJM
lb2rptvk3kG0xrRpGKSYtT+m18eOh2XxnQGwnk1shsoNNeN6WV0ftW5mBvZJ
OcOaJQEahql5Ra1uAZDZt3kmcRklSeXoXwBsFac5xuiyN6KIAKbe50VrlA+S
YYk1tuNYyCA4J89Yf+7USDEW5aL8jjm2f2Tf/xK7Ck35+T/raXHhduy70PHq
q/Wbr8rxCvvOFBQZuC6wR9E0dPcbH3HaNCySsdIEq/Sja9zPTD/wuqZiWViE
ah/FMtIc9WCMPJ0aNAJV45zBHORb1Sw1dIerWrYsQJOUSNS3wS00CCf4ZuyB
8/Gzj7Ii1OGGeIGdueGfitHdVxi6trfZ9hIjlbTQcGvJp4nJvfPab1NhZPKZ
dNHhEGu69huut+dt/S6jNEhhscWP0xUF9UbzFwWkzvvVTOYM4Vs2mpHjG2ty
0GDMuN7Jpczkew1SzhB1dvRQKzjqr3Yx0q87vLKZIq/YhYzaN8PGKbQ7lVrl
OORRNDzJpCqBN/qAqNoBiAudddKYemGV+0J7UzxCLDfxxltweN/MgnuZyw3p
kBpnDUmoj8935xUNxy5TAbzjUBj82zSvxO4BHfix7ZutnpjdfiyJ/S5N3U5K
5Wg50rnHEU/aK/qSbVsIip7SR6ZGpoe0bjz5oHuGnHX5zvlHxFtlggfZaGLd
IBVtZH2EVXVQSlE/FPNXNUEVdyQYFWsoEOWZhvNiGdTBpww12R56Xt6CZpEv
caf4w19li3bhLdn1hqrXSSFVmKjJSKvaDZ+gZPVPdyFQQjGk1vXc30vmakgE
FpB2tH0uqnW29IFm5Sdje5AmaX6xs+F6ngKOz7EhrQ62QBAnepw7D19lQMYW
mkAjzhPOeCDFLU7hA7J91aPz+KZG97AmlkbzEFvVHbk0/iOHODIcrtTMJRuW
f9iwifOTnVdzdoUnL9Wk36WE+3gAsxATyXrJSMN4H/bjioK+bamfvsCbjrgT
GZMr2WItWve7JcSPeSCeeZmaRNrW9elOqBNR5yxo3ashwXfvCjTiZgH7MZQq
Ar3ibzoTUSWW1qTsVSG/CtwuXFtw99A1tXieen+5gADK+kfhJDLhWYywAY/E
VYlZO2RvbJVflZcd5H3mD7ES2SXvkW1VYf4uwJLdZmRsMMGepjl4rtNZUzy4
//SViiZoAfa7ZO3k10cEi11DANjzbaO40GMkjcChIjkUuwWljx683G7nb/at
y7bYOHe5vzb5KUxXRKz2vTSuX628trqinkC3j2oIpnoxsgqEAXd/PsHrY5KN
CpQuOsYS56UYipFdhKQXC6Ss6tFmG1099OBymMsRBn7XacNthaP0nE8uf4Ea
bVThmF5yF9B3JHuN97mmxCOUq8YczJHUeAwlcyFodqcIYsUA25CDkT/rBZ4z
4R7nly2OBnuzPCNg3mtwqMchRG0INQTx5Ch3s/4N5rKcnKOD3+tiKOlNiOfO
jNJQy/F/bFeoz0YqkdPm5VCnmAqDWTvC09QRYMRUep5ivYLy5K7EpnRorKab
jt32YOARlrVZEpDjNp2+OBHLY1mDeFZhzcVReJqWGW10SXbbSZTEwmH9oSzC
gj7gp2uG5ydShoFauj5UiplqlnumszZTzljBBlOSxeOYA9fEhnzN2R6N+MuB
EOmODA9Cxo/3aTqpSFv3laq3pPf8Sm1oiLI5Wd4wrKv1MoBla6QgA4hj093b
NQiFg27YTfLf52SSVGkP9lU9AiJov8ied8FWAbLV5emlCHZmdaedtb5fq+pJ
Y1NTzbTG62HRiSIzYKYLjurubsxBBm+0lT3kJ3q7Zt1oHbfnlz2Zl1Ao9sV7
BTiQ6TcDZCMzBS9ojKPBWLN+ALMgMTaKjjUak/zViRgBt2bb0gQori4agIkj
7xXGlWxPejY44psVu51GG6/9ofK6IgL5gVkeEPW29LothGZ0HMKTiLfVbEVN
fIGu+/gVkTcROWxk+bQ8YRxc7SOfK53XtLvDZd6h946i+vRCOcQXM3+3HpY0
4tyxIEKVzhrMROmEYs4JD+aUgxUG7xA11JJpA/tJomHjOfF/gMduY8SDGR+u
XqJ8/ML9ejlz/aVfZi7JvGoCltgVrKiP+K0QjZjOm9t8t71L6Ne1iqH+Hb4O
F79BZ/9knka38iA9iwBQMn7xlkseioUsf9QhgW3S40G5tWvyoLigeXCW3nIN
GtAcaVbQHa96Q5GW4cP3BvtJQ8TIO/GlR+CbMtFSBSJ8SUGRNO37yyPuv1WF
kPHMehMJLVJAfGvRA7UF6mt6+q9rwFcczEWck+QAQVGRngsFXrK3lsg3RFKX
UfgTZJiulNBOkVvZHoSzo3OTWncAlcCpZupv+Z8EP686I7P0fbZTAhw4Jb3Y
YtIDCjiXEapQVV1JsAfJgIkSJuyQJgYyhAZGF9lJauz4cgxvrOnf+T/nnyLB
ni5DEoZ8QAHmwr7sm/YWx4A3rhUStnsjH/5skuhPkmZaNtODSWy3nSlPHEZ6
qt4zAOSoI+28JLCLYfdXKDlD8naF/9cljfGnfdYJ81A2PoiauYO+ILSJF2O5
LPAlvjchEHdHmWINUneZtNaWq1ucWQRfKD+6iDPkNbMkxP4+B17gLxDHQrEo
JKIVOgO71EbyBZHt51E8mY3rR1m0iwanOsBbHg5OlYDQXarZ2FhIvQg8uLxq
p646oHWSvv6qB5vVE/MT8ns2QfrXymTSvdLL1EoRtIH75p23g6nGL5UzPzET
e8gO5IQqzpG9g+X1QwzB9h+xca7qNprqTRv84tVRfwZsKyGBiMo/TWigvs+T
EB7H6OiZ8suN0GH1+RqwmDOjotILPl0poVb+hirhXPQagtSbiU8WYXgpe2h0
YjdhNMdfWDmrqR9lyzLSd/KgXbHftqyeS9Ug5M0kzxObu6IwaEDv4HaIa0Nk
PF0VJ1HHQAOnL5aSDAGDU69Y6+4ZMc4XsTNpDHZijAPtS+6JSQ+VeeR+GwG5
biM3cxWXuPAOGNffOPw0Z4A12mZMkgXmqmGH2zU9yE8wE1pcUAWEclERhe6i
4wEV/3XXJXmahNT9YTVYyGT4tsij91d2qUW3Og6QNrBjACgODxgwI4/XQLim
IKzp2YshLQV12YHij94Mi7Id25xDwyDowXSleRqXfF0tEaKCnNljBsQVo3Fl
lMDn07BbrmPhE/mtFrvPEzCsij1Ii95F+VM5fs2hvbJixqwYrWb4W/bwd/X4
cfXsnGgTZzPS2bBSc2Blba0lC5LcYNMRoFZHjL/3kwXOCtw6O2xsTWvi6C6i
yazckMvE8ZjpB7VYUo/xIjYQxvs5+bf439PrYNYG/sCZYzS9G/PULttgISol
lohu72qC3+auLEZdfbnCPFTxy5T82DNPlpls+JZfue4l3LSsGHgG3N7ngqWU
h3fyIIJxpTcgbGJJ0pzdcEMl9+t6QBb6VebyJnLHkgAFvhzZet+JD4O5TgYr
9DtYN7H/EqfQfmrj7OIbLm6uQbh0Yj/DWfls5nVfWCPrM7CcV1RXtrthHalJ
gGLvJDh9HfKyXAx9VvtTeoMrMbK9LO7iBBtLDGo0KadE6poC1b/IVfw1Xjt1
rlNIWsTxfNvcTDeBjnpYlBUGNg12qh4QAbieOm6+2TR2uJd4PBYSzgAfF0xB
oK38zWB8PPTUcjCSSwA8hnRW6DWoCpSxZ810N4lfhMG5/mmW+sI5AsZrhCv0
5McbQUTDDok55EPWeXHYMMMTZFh/3vljS08FYi16Cr3Ib6/cD144Ha/I4RhN
L/xq7cCCWjZnXCA1c0kywmbdhi7str60cywXElzX/oWj3PlIzECIUzsZjEXo
2J5qe/aVvMgXC+H2V1GHPH3VPGnkNBB78rfznCIM2c8FKDss0pVL9ZgG+K/m
0XkYiITFQs8Z3UHL/pooumCo84Uu84TmDsu7dTJsyo6JJ0LGVH7nw6ZpRaHV
yyiwdNsxj1wNSTlelQGatghuS+4nRApMbPjM8KdxsZbChg9yH9ZRGGtkNSFC
yE9nm9v3QLlooyDKNXW/JV/tP3QGyu3pBnV4EOaREu9hpOjBQem9QhXW6rwU
uSoZi0JM5IyZJise/JufLWa5IMKs/b7PdKoe8lk7gR3Meld24tHRWPg7R9cA
G0AwnCCt0VC30elefuQdVmjJslJJtk2muTAcioe77hyVMVFHvLkMf4aSNhGi
1kZ4PhUp5U0Rlar7BoxVFuaz6qSV2nJ56c60vq2oBR2DexdnLsHgHj1B04nC
ogvCzVKjWa/JcUZdRxVXo47kUb817l+WpKtXhgoRqefOq1wWsLzmpUd1AhML
LFl9YycKvdCmN1jnHhKSyRFm/qOQwRYU5enfkxefpe4SbXvsaB/PFAf+tmR9
GGU3m+OZvngoWEbX+PGUOChr0GLtM+h7Ino9m+sHhiddReAd0tI/9CS2RX7y
haxqwhTlVoQ81EL6re29dj3ck1FoIVhNidK691DA1Z5JRUhcy739qy3F23R+
XO0u1RFTQ92sWiENPYAqvm81fP418Y7p0vZtQ47lGZz/EMMBLe6PDZeCWWDQ
VWxjREGikQFZP7GMp0xI5zvvN8l8G85PXeukMLCNh+QutsZAqsjvcHysKPS1
yTcbH7sZpuNcIOeFzFmTrdpoD2gHSDoiahHVAECe3yV5Kc2nANST/vogyBB/
kY9iv/QjpCw1cRqzqSwwBBqGaTV5vrSdlKezuL44s+Op02Q0gTCWy9FFwXwz
HwCedEl7ehMLvfAZU++yc0yeCy2qZkh9PZ4fevuJonxnBSTSigU3kI2ZMfbZ
oqOroScz0vyROqjzpY5htj2liga7w4+HyQa0kO1ZhQlTP5wD9d9ACnb/u1EC
LbvAODx5NVm6O5tRlTp17YPdpJuZuxJMd7uY5IjtaU8+8pLxUkPrEwmlencI
LrHdBa1H6CuYRY5tivPEz9m7jtNyqYUMVk3zU7nNdj+2hiu2u039NO121Yh+
BjpTMKQtQPqqKLVUo1BeLrkbDmepP8YUfspDDTwQVgc/YRwVhAHKaNLWfu1r
EuoPMt1+fj2V4HaZy1ZAijEJQhY4eZArng/gif3oXQSoiIbcKrhX5+o5rTCm
i0IuanEl7+q0uI81KcnJQu6d5zg6C7We2Qr0xzsysW9mmqr4JC6KTrv0Bx9t
Nwv4ioWyKtIcQ20QYXnmOEpLq6zdqt90tk0ussTQbMgw43EYl79Ck3iI0x3m
ckCKlRApy2HWC3LiHsoIZyEuUh/q2qkyI8kQDjFh8pglYlZpGDUTKwWA22Hl
ryTzCz8eiTHlfM14y9qmhLJ4ahRchpHKFFEJF+NSybbcNpz+7FB2tz+aYVOL
AKZSV92eTBx2JqcoIckyjxqcEwf5BHnCi4jQAuo8yOBdD6VEVnVEeIstcUhI
/aWqui2daek/Ajfx0ISyuf0P56/y8XxcRmMCICEYxMv5vBkegr0X1y/qZvFC
g2BGtlYgl9cU7RBFmi788o7omEDvgXf0+g8JGA5XaE4wiJ5GqXgXU+h6wSeW
HSAoj0Q8+v91UWutB6GNQLL0QhC1FRHlmZUgAUcUv07OYMxKHbgeGuVygH+v
e0QJbVMXradtp4pqDeVlWFrfEIUK8p/Wbb28/VY8HW/0xEkQ6EsZ3TOCN0Mv
2nxY5gYUxLHWx24ofak2zxNiNnPmuLAQSc75+Pn4pWmOD0EV62/7oKPkSd8X
it6uqxrr50ljZLnFkegESTcqOvG+J0zYt9EjhxFHzS72unxN4KDOSigtEH4g
w8D9rONCcFvGu6GrqNymWimiBobLiOAqWlPIDwEZ2+/va9W3AeNAWnNn+1uK
LYS/T4a3/G0/3+2dzHji6Aez4wL4m9PHl6LyjijP+VkMC0TXo4Tf1g1ddDYi
ESiFQ2bSOenRwotpwZth+7vGT1ZzXOJBpFzjGhUtOLCcDP9HnngIvTxg7tsF
n4f9LO0yQCopGlEH9PzcywBMpBTmK9u8uPhZAMm+T2BOmtZ1J7no+6n9VkPN
HHJh578ncVvKCS1iKi2kNray0SzrILT15NmYfquQUXoLLySgW1PNuPD/ZFoh
NWBnJddTnsndzRdKgW05eKqQURRy6kZmISfXCQbnZlU5p5zbFMUYGxmy9M9V
+JEXTdhz3uhCfVVkqEyBTQig+pvrkuZ2Ps/8ZtEQ5n8OXQMZ+7hR6gMXUfv+
J7llBHmX0CS5ochFhQYhDXeWAb3nk76uEcyGgf2MDlTB+F+qI726Cpkfp7Tw
QAcwitoiUqj/tAjVqPgV/EphXsusOROh5PYhtZg18Z66AwBkfWi6yrWEJZfB
3zaf9JUX4x8ukmE4IB7tZUSsukF3n3QoY3vV/XzJobua6Y7S9pSStoukFN0c
tGUZpAS1Z6AqITcYWlupEkbxYXYIAPUD/MWF2Mub9NAdd6RW5LLqp5h8hmGC
zoBseX8IsfNtI7iPL4oycarafAGo/KsHYW3TfHHqgUcMh8qU1ebG+1yyYFRD
bwPk3A/t5OCE5ghEHEWHlpJye+ZL5iVw4eq+bVpDj9U+cS54n8gHvGgqA+SW
UNGcz3Xp5DkDLUGps9xkL/Et7tSpx8KhtkAH41AMnxLkuK+QHTaQMd1fh/GR
scU24IKEal6q4aQ1o/BsA/0z0P/Q0JDDvTx5Az9btmld1ulwLagqUhaJGI8Y
3ssChAs7BL63qyoSK1qmPRG8eP83cpWsMJuCKDbTA/LP5PY06fNvpnMdTs9a
yCq0MxMNgKZXhVbISm/FnJ0MtFXmVtFFiubbTkk24o35w5jIJ2sozdYTtfrP
+FaLy2Q+cH4lQxpetEyUJUoTekPPBiJMPHyl0QDDx00L74p5jAbvgEKC/4be
h0OewFf9WQKExqMUTJPOk5VPaverviasxBKruwIqjnm9jDcQYbiShCpChx8J
LwwGQVqVwEtGpSl6jQEIEpbWikQCHiPj0PX1Jk4/3/dU03pULxN9lrTx7C6f
sEz41DTI5zYSGx1apHRK8IhOk5Zt5t8QkDwrwW+M6WnmMChTMBn0RrMOPlAM
E4vFkl5ubyyRYgpz6V6rxHcka9ybT6RAjW5/sH/V8ehkTrrPGo2N9A+24R4c
KQgsiTdQMLIHBgpwL95SRTYWfc6/3JJqOrL7PwneIX0cnD49Kd4vypwawd/g
/RFxYj3ogBku+tUXcbBqf0MVsXDLZEbqegtoKSGC1Z7kcEQ/tkWFYcXmA897
HYPg6luZsBonSAHGwso7C4572qwRDVk74eXLe4E73bW81OlJpQE8ZsuDaQCm
SP1NiSyHz/eD0f3bLsVZ6dYk1nLgND9SdQEnI/kta00iKJ961NQHtdcvWBT0
IgfJ+avVgjpYEd2QBR9e6h4bzbzWOOxN6qRr1hVLFH4ooXQ+lDno+XROtKeh
RI/gBJobvGuv8oKhQw4Lfo3gDtUxFlDuoaBDaEKNeOgAiw6csAU25AdTRLvH
670/iSf6iCphx980Rq78XpeKGwprPOXfieHm/NFWxwYc2xw2t/5W0gyNvEB7
4K5ToYSUMAdd7or5mshJnLjpHET4BE7qcpiMfJruS0NzH0f/ajks/en3tjOE
J5XqByEzVLOtzF6iMEnC30F6pe3L+I28DN4906vR/5tLLmDYg7K9OaJzyTit
yRpWSWSzENT1uVDSAY/kk8sW/nzZR8s8nKsYgtJ0bl+JyJFInTQ3as4mQYcD
BP/j75ly5izHVO5RnQLs3DMK/1BlUB3iengLff9BrO9mSiB6dBx8Z5SAW0+o
Mreeo/JrYjYoStLSv54+5r7Dfn1Q7V66j4tlgUoWBgR8aNlf8DcBZmSvOgF/
5Egmc09xm09tnF0v5N5KYuwd/2TrHOvctMesXbuppXqNQ0r6j7NvssBxqIAw
+6kIYZOe/r8cUhc44vPoATVIOetNA/RmfZOijr78S4jUBPD+0wwymcn8lgIN
HvhR/ofEN9ctViPiUcDCuy4GKzvQHt4c9MWGyDuRcCaql3dOOkReo95aBgA2
c1hsFQlPpKMPiXikrmWqyGucJjmPb8tR5VXk0Au3DxNMvYp/sxU5A3hRJ4wS
BeZdhcL92b3YwKTJ7ZdYggBV4ugWdMAlnQOdl2CoUZqPgX219+ZLTg9x/YVL
DyC/nldOORleAcDbBMwPvw7F6zQw/I4L3/7HOt7Zyz2CVYQwUaNQtD7PhOwp
mZrjIcAVbf5TpSWpDbMuS9Wa3c+s4/JJdmcQbKAQNEBn51ZCSUwNgnH7t/2X
maUs8B38sa3cDBQPPSSt0R3R2xbFnA7aONZ1EuTegi8ATXooIn6kicpZ+XOC
bmlZD+586g6nWiRX8dRWwrjVBy71g6AqOLmCwtwZkAMDfprD4UQaaJCloHW3
oVIQp/SAuRryjTp2SSi7NYPvUzvKdu0jIdUuBcuEtdAvzo8WjC28Uadau2y0
gPoGQh104Gz41kwHnszUB9lLvgyNoqfvprdUTXCBq/Qk1d3vev5NUQA+Y/SS
gXNwLuPpCvgCZuo6JSNcjlEScGWw1B216L8QEilmtOa+nqH6GTKFyLrYVvW0
3vBkqg8qXzwWTErBJy36UmF+lII5NmJ5dV3W+8IC2a9UPCqpnMCFhHbw/xmr
wTCyu9EfdNDv88ITW11Hy9Qlq1Tsk8tiXrP8k0GgQ0PzkAvUeGA4osHpZo7y
qWqeHBwD2jpJc02Q3G+caJBMqFUAv8NP78cxLI3JTS1DX/N9TpnfT0RG26RC
5IW54+wP3RE/DULGAG8QDPZ0AdA5JbLttvb7FdgjZMf6EWV+v1TnNHTCo6vk
WkYL50yRKGCyfrFpAAlFjBvq7kOcO4LzU9TDtemM7W1YeSa2cNEpD/F80Biy
JB6VFinIw25/k2TOG3/Ca6JhNE2KPszfuPn3Ur+dSB2UQr3zpOUmORH0BG3u
ieyz6+STIuNp3Iq2wgu+/vIHhCMIq/dpwT07oyEktK5m3PII+8+0WYSqbtPi
qEQTheDRA3A4ASw1ThK2My/01gGFMbvohsFIYACoSB20Bk/S+ylgFSkmfGmb
RsdIjP7S79CmEc/T8YfFDXdK849LL1W8oJtHgW+c245yhYZDljgpkl+f/L2r
pj1wCDIXHO4CUWw/G9rWFxFdiDC0rquhVLJA9OR3Npdb9It5YUbEvop1btcw
k7Ps+oXlHbMxiUAG5mnJVctT5wgqlK/uYWLW75O3lgHWyoQ758WBy3oWxuZK
EBdcap5GAmYvTIvG9Q9n+11Y6WHyeSbdM8t8Q5bGf2F3klEwfRTD9sIYEuqT
MGdu/vLGvaD7ir28FbD1d0Up8Rr+pIoOtAXkT+3mD/13th3nnX3hnnjQ30HW
NwtEZ9B4wgXdQwIOD13t5GCDY1mM59BrwX0lae5BowgkjE53aDltqe+jn+wT
uEfijluWnLvJWub81iC7CDyLpy3LfbhHxeRfrX/HQqP4aZUnvzXA+JxHugRZ
wLMUFR+AXo3En+Q/qr+wsez1r0d0MD5GwvMygbsYjo4B3F8g8wMV2JthXpf6
0KoD3XHv+Qto5/4nk+18dVHF1T6kNM0GlydtQTRWAfiIneJ1PdXE8uvmpV36
wEbo5G416rvQuH92aeaKceNUI3goVS7G8It+LSiGok5Fq9bDVAxclRKaC6nY
hfMGtbt8GBtuHWor/LBMVIgvwygmCNjiNnnN0fAXAH2xwjk0gddkKS3cUWn5
N+VaLrsEV05F89q8eQggMmo9bRbhXrJRW0H1P8i4vdqz8f+TiQ6Q7pJuhjhJ
idBfP5VdXOIzMWAYLwI6Kts8C4areDpOxKXa00uDgMVplUo6LFzLVusTgfCv
fZKxxdiJiywL9RFT0SqGhcNmhX+7QSvrGldf2ovzVjrlTSXsvpR1i7BfCc26
lBSxpa5I1AMgCSMb+0LwwM5YniWSAOVdJ99Sn/fhq6hyVaH8+8oF+cmsjITV
Oc54pHSu648u6ZC8napnP+d/hCUVhh1PhUNMUlGTMReBToagWgoHkZgGPi20
RRLzf1HAVtyRrTsAqdzzGj2uwscFaU0MxkAR30SWgtxNngMFyHk1AU63azIp
02QE8uCdJtchqxlh7MjTVoboC+0vr1RHxSOurUDbr1Vj2b9oLPGOaqvYi1UH
GffOwXymUbbqhLMMeUfVNr7JDSzold06W7lUJhgVIZKDbvNjTUD4108RaBVK
plNpzj33UDLr9HD9PsF20mYFyOr9hBklh6La+n2lV4WURFUPuhVsz+LrS8V5
4XJlIPcLQ3iqchKbfIU1XGH7Qr2p4ooliHbtwgg1IbDaubJOUccRUIVbHObY
NgIX1fYpZ7EwJJV4JSqwLO9+mNSGdiOvJZ4BdrD+AcsuJDmf41a/ocPItSfR
2ty2BToGotWcQ/FrURk+7M3I4f5DK6ghDjohk6XU9JsDsXuKKI4WHZG9ciKZ
ZlMgr0Scl0I6s4nXW9oNJbZ3xShUmoNRDxYq0Mzb6E1MGO5R+HjXp7jjJkRM
vi9C27YMnazfF0w0jhQ6KjXbvAAvrxndmUxfSU3se9HS/ZTpxuKvIsGs/1kO
sqOj4gj7UUnTOAijRDoqrgFB7VlQGq5uUcpiJwAB8JWCvFOIOtwzkrZhcEPq
Dn0M+J78FjLDckY3fqID5iFVkPwGFYGZM30CHMRJLzO3yr724aDo2nNJHrLt
kThTaF75BMWMXUN5X5rEcG3QpkXMqDMJCjxQRJqKXqBov2qe7FYof6h7RYFi
sVPKY61HSQ1hQfok6zyREHB6C2yMyl1/L+R0CvDjHV1hgJYaglqwGCc4xt4N
mXkEP73tWXI4DAArhPCrf0UtFXtS53LIkdtyOILCQg+8cAVx8c40wV9h8wMO
8UP6icEa+kYEnnAkvO+qWuIDviKE8CTHWOYpB7DU88ZFzFNxQwR33dgmz+Ky
5etCR8qHr3/MbzZtmT5qkmtemmTtgqi78xx1T+WW6tpbiEjf9t6wJD6PJ6ym
+VXaJI6MnRAK7ARSWjSguz0B22n0HahfUW2Kiu7I0nYbUkNusVNWOAD70ftS
64NYD4guZKaD+8pqn3oy2yB+3XZsm2Xbjy9akgvnrWMomKQnLCeJYQhlsnbe
9uU6nFE/CJYd45CjlDgSOt7/CrJaQIMuao4kn9ivxhQGyIVRR9OL4WCjQquX
AV3dN+etAiZ4MS33poR6icAzRm28aGCbHadKEwDPhfUCgfM3THE2Nr+HsaHz
MeCl+BfG/1WJb/ql5hWSKKQqJd1KImFIi6xJpplHNpNUZQL1oPl8U8EX5VzQ
PLSnmlbHLXy/Z3g9rk5uPVC/lh73JMB4tw+VfKv6Bo6ksQlBhmDQqqkyv4YQ
G54TjKCPfrvtYf3QBHeUH/VPB2PkhHYrjNIACbCXJhNK10OiVXLQzh3QbSw7
dw73zF1aIKJBYQpgbGLR7hHaELqRD853vKhtoPrwRqpEiiuh6wCWdIMrrLnR
I4j+CCv3IrHwogc+HxLcB9ukfXN2d6cLqnQmYqRh+c/o4HCbOynJ2gTFpOPa
T0/IFI7b4664YzLBTDI3ShMEnr/sbyFXhFxyB1Ei3AbTs7VNRKkzLj0/OxfF
1AM9Wmr32hPoDzDD9dcQI0JXkEKqqnKPK8GlcLqe+mOHZ9KZDDpZGx7DU1UE
Br4ywYQ8Nwx7rZ47ktR/NTRMZUQpYYltDxCHydHTMS4aMimVG9yKo6c7Auw5
TbTnAPcgvxZVj3rAHgESQRqRWOC5qlV7JbBgHMjxvM0zUGYLSfA7w8HBZH5k
0T50VwrSYbz3ErxqgwnqiiKGzMHlJ5zSv7eUpkhf8ENd4TD1YI2j7EjsJK5i
eGX6XAuuzan6kNBiaYzuOnw07gQqOCtUUbu5gOR7N58B3vH/wN/7DTVoCkiO
Li6yyVgMf9N2t+09dgMPPqVB5DvL8jKCCUKt3pvO1OuJeRP9UA/Nne2S1SYh
GnYCwdtC6zmEf305dgeYeknxDwl+3xoPn/a79jhk1KvcSO/XAA/IDg5uhjy7
WU+d9eCC7IxN486pwDV2MHtFuMuQXe+OIfKvwKneST5zVh8LvNSHOTdwPHx8
6uENxE+5pXQ3jr1EVpG+54+oInLk17iNAoqPvAGqbG58AyFeQ4dQcVf16Dsb
nS2IRS880G4yletYZH/f/HTySjNjbxNy2ielsTQ6dpj7munD+CpA/kRiEP0S
cPH0meiVbKdWTgihI1oBETIkn0KJwYllHtc+GAoBivGEPCYJ8pMoUMs10rC9
kWq5loYYyZ9bY5qMkNuQQuROWwahgkp+SXPLv3NptPIGcBQl4krXXZdDJvN9
H3SCZlQW4qEHyhCOxIiQrYHxHxmwYTzH32a0CLfCbPMN24s9KhhFwPeZpeBF
0YzxEreMpudkua38V1TwhuTbeDijlG3EQvghxEYrFydu+hcXAgpBRwN/dROB
jvJPx+p8Svsn8NEOqPvNxUOYsSKgc4K/mbhAlMEkCuSmXvbNzCq6PiVCbnJi
EY/mgK8qQcB2iFy0IjCnNYpF68iD+4BDNSxk2+Q0AMSx7uG3lYRQPk2b8szY
Ib+W5wLcadwLYSRGOqojjsjzBm8zMtYhqsUFVAsZ1s7miw7q74MPMwaMfMNU
gzr4SuAGzc/N+dr7ZGwHLk+L+hg6zemRidGQ7IBqGu2vZQl6xmEnMfvdXCO9
XkgPzVoZWFgW7SzggaxD30aF4yv9tiHKy9vKcl4Ob+/tnG+YfW661RxjHRki
wsK81VGJRUHtt0K8Bh0QgfyQV/Jj1hgHFSu91CT/PDRSNa4f0F6I2eP3busC
3CfAxPoaAHeOzCgvO7JDAgFhK8ABajsaj5xwQwd/XjH42cIhQ/ndyt6W/Sdo
aAwFFfS+dHLfHuUWMd8feZcRfUhFlcdejoKlXqa/LiqrzPmcrQp1CAkkbWt5
iZK+HC8j0EKVCPGhwP3z/HE4Qum7qz8lg3xB4NRhvb2P+zcnVmVC/ti5o2R2
MitlhtCPJJU4fiVwZ/g6fNQlKd7HtVxwYJD8cMnvoU76qbpZqq7uTQQLgI/b
S2M974vLxLgMb+nSOF7pt9N2CNjyDemiQHu3ERlVD64jJDm4zMJQBURsfRuy
Cr3se9gqomJcY2ahz9/vMeRpKw0XgWChUxa/p6UP3FTwOoF9kYHht7Pn1kiH
X4y/DhOIMsTZqUiTRUhH/o5CWHk9Loiqa+iQm+/vIh2bBDAyagaKL9ZA5wue
pVzO1/676B1ZuvAlvftGskyNFyjnpi8VEmYeLjZoAabwYL6C8moBffQ+M2EG
2jtfG2gQMDtJTpMrrodC+8MWvymUQ5geLmL0SjAIg3x4tgKogQZh+uNY0npr
mePnDBf/eZcx1eMy93Y0+eJzR3qkROWAOF9aYury2KC/cMR+FLEw0USDsWyO
jTjTlU4IbQ8KhIhMcCu/VCkg2h7LVZcg7XnpFHrFPdHysu6OnkMywNhh5V27
1vuh5eN9gAaosvOBOcgUockDo/Fbdu4bynRoC/pCtb9fw0kwtCHQPPomd/Z1
moeNnBhxQ2Ogum4vL0it/TLSPhCW8UsgZpHAKhSJGJ35APcrQxKSB34F8lqD
3D4EitoQSrsjUILkHiVYC1CvKpFMTlNELsbpvFIjGXci8ayMWpIGivN91jCc
eJiBJWqnjcdryX9qYqC0j6HGpuzeWT/Vc03q0fjIqOMrz42eH+Rm/SB7UVGC
rtos7s3PDAxn3OG1mapyOcWWyENKZd2vIPuGfN3py8Mx8VPgvqhdjywZWCB8
Xe91eoY/xj5MkklAI7a4RkQ3I6KeG7NdHd/IMB6/bK36uzEKrtmLQlYpZIUW
xM9M2F3fn91cycg3nRJYqIbNnVWFSkJGLlxJFvfUnLitBXDj0mF8pAZUk2qh
PQJ9EV45ofie9Br6lrScrp9dYuFiVMZFjpozNna63rn9MkK9vk8/Xz1f5ybU
kTIkz8EnHRDpi7P5WkjisDMGmdElEa+CBixHrkB0U8Q2fjYejAgS4GSyAyLA
4otCppLf8vwCxexQTQighc6vbLRytdzMUMBL4AicnZAw3YKMCTGXjkXl8ysd
vq4IKodg3bpmQX56Vz5gzcDDDt/xbq3c3pa+yVDmVQNA36u5F8yDHVvc9K3l
7Qz0AYUk2+y+Dm6je3u2FPQL5WhKxa9FHlFOcY3R+gt8uUFhvor0reD3tDly
d5jzczz+TMyIg4V8866Q9gmky+S76gnYKBcwoOxDXmLqrmFbL6vy4HHM6yB1
gIozalQ8yUeuLIm76S8WAuTZea42ndYd0DCm68kAOaTtVFZOki8J5724tTpp
uCZbj+fXteF4zVyZ7eupXlXWIArOWsI/5+bJdIOrr5MG/ETw8PFmY83Dw0nh
SkLECvpr1sGFandovd3CEcN3QjDZ0aTiw1RlRV7bjFD0kimxDI7ry6dkwb4g
HPpPL1wZs7HDjMXBv0uHGbAzPOnhBiLzKBE7eV1d/xsNzainTwxr3uTr6/d1
w/DLctqHVQg4lfntB2vuu1ET/a9WHcFwOJRRXmfdE8l/KnqgyHztCq72ysGE
PxlxF+VPZSR10xJZhiGRla4xqT0uNitPVHblk7s7rKZP021bbId0vdIcQJQG
EpoXvU7nxF3AuGkcy6DiiQ2tVWV7Poc1Cm4/F6s3CnH4/d8z00Knu4MgvTsp
JTMiDtAIiOfbjhkUeHXVwrfQD7/dKZmNhDz5r0Avyau/7qlHbYWpJTwueBUG
Q/nOjczGvchv+bLWM4t9AO1OU+LPbxHM1NKDQrWGrCSsWoISFsS1ifoutqBH
yV9eWQ8Ts3GZpYKJGzkQ7bufnlLfzSUa340XsPTeHdUrQ1BEIpB1d9Zqpz3z
Koa6DVfBBNR2Zcg5ePEkDGGimiADfzKXpuJxqEdUqE/eTLiiXD/BYmOaD+s2
gF4WbAi9vEa5/ytZJe4stykl86PX+HACr3mmCChq+mgCxwY3Y1G0yBCNPRDl
une6kNSJAusTq04LiaxfF6jopJDwH4fIjyL7B2yop5F3pq/H7f6I/E4wlYik
vbi6LNLrPVFgvCYDmmpfPO0ViP35dsmW+ySSLv1ZBHMjM3TfK6FLiIrEGuiy
Gdsg9bByirOI7PUg5EwuN5btuXI98qqyL871kesIb1o60QYg56O2j2+L0SA4
AJLTg+QV2tnLet2+v7g6ZUl0AXeVR1xxQAkX0CaDksxyxsfA9+5Y0lcG2JCG
8u1vkxcfxylgtcsiiLKv85amvHkzCy+BWkZKo2fmJzRGbGqBLGSg+n23hl3T
LXap4R6xggMtDvLIM1i5vvM1WIxgr/MG5W+NylOqouYdju4yJCqs7g5/GmFS
89SINEmQQ6xGuV9sBbwp8Sz83NycB+GT25kNeKis+8v+CEcMgaaiBxCuoIWr
teqTB+GAwI28q/w7J6RqI0WYtY0rwPMts+RlfOkB8qXfnTK3uug0AZeWf0CE
UdElKDGwiTgAqc1zFKK2v4vxJ9Zj+I3Yh10qaolp1yRF+ORMIHq/cGbp60E8
+Eg5Z0zNAoL/VMOmMlYrISQPU48kJ6g4gRjirb0PXOocCDv1jpcswDWxEDJK
9ywKLU3EEyRdq0AlmkhW2dvNL1Vt8QfOH8aQSH2WAzbQMBz4oRHumD3yE7dk
Ts5beuCAoUgI3X+q7PSqP/43g3EluTUJ2OzYTC0FsqXncD1fovTWqcO23EdQ
meKo235XkRF2aE2KXJmBqGBUTuHvDwPTAmc7P4p5ebvbm2vBKiMJ8sZ6oECF
R4876DUdlDEyDBYBWYCENcLG8QEdWcSMlXd3tPuWebrSFopmBlfD2OAg8JPp
oRufy1qiVeQ8H7u6Rzw/PoXCkCXMMZGbG2vSop7nKluQ7EO0Tb4pCH10o04f
yjh4sdNyBQpjlTk0D9eeV8eqViZIn202eCHE+LsmCAVkxuS0MKLQlqI0+iD4
YWjvxgE3BtDCJykEVsfBWEV7PxtevG4wXX+eIVd/GQTSTaizfl3kac9B3Tm9
E2d61eFXdWBzQIas6oBUwYjVExKbehjoPHZPNSspXN/ODWImItlHDR03Cv6b
OOKi9MAoB8Dvnd3sizTKcnoq5fvpkmrB1aJUNjUFoUVilK2uS2tzKd/TnrXm
+WvwbiNRZuasVr0KLEqKao7o69EKFSQ0vHo+6ZeN/FOAYHeqG9OOcLkbeQyE
upNtCnviEsfgN3lNxoqQI4NqdIVSo9gKceA0yYgAIGGpdHBE+VWWa1xe/OQ1
hTEuqgbJVqmiVaron7TrhkPIh2iiTTutkzx+ck6Sd+DOqWG11nc5sBjbGsUt
Pxa9WZKFi4whTvCC+BZUt8GKenM44aPEm4CPG0qp4Hz5yZr8IUyLspRSXwDx
lRfH9wnvyg1idTdn0+8Fbmz/id3XttxKL1GOVYoKQ3hvuxHrpbUsx2264rKd
Cvg+y61o98m5cgReT54Ezj5yoOD15xVvNCgxT3tuyDJdZtwBYymtmXst0CKm
03yelPgudesszZIZ0L6NB7TiXl5gQ8HMnfWGLUHCj77mjfyDf4/UjrXfoJQ5
IwETTapaEt7k9rbAYODr57Hs2VSm138Xc2a3tYJsM6pQ8VGL9gZO3cc4O0pW
r7zxUhTKzJdTkYqMoG0tMg/tG4cN/idd4ri9aaby8EnlViFpnMzYDDRlKrXX
HNmtw3zfKESHUJ5F0WBMI0HJ12NJeLAPidu/NS+AqBpUw13j4ZDirf9dPYgG
5PITIW2AfKzOmhFTRDXwY+Ld8/QbS9Z2HLgLc8+TSEvmgwnEDJT+dJsy9KG0
OxlS/DIjYHk0hhCHNWOsRt/tRnbrQL+norp+cwZ8JyXGW3XlR0D9d2k0ezEX
9y3HROIKMLPGP2Hd8YfDIpKQXkO6ZPq1GLvg7TZPn6yXQVeVJi/2kBCxsUSM
pYy+GV0Ox8P92/+yDu39eQKfkCh08eR0tvlm9qN8ajMk3sGsbVd8sub/R7is
JOhM4y62aQB/B/b1datbhaaxQbutz+PxvxuDm3TTMukd6lcSlUNOsYeaVOnr
y6a5EQZkyhY80sFXgyzzYv2Wcb0ZJIbzJBEK2iIi20jWXH0z1V0Mg/hp9itj
qIWhWscHAkLGwkw5AbNWgkTpwa97EBuWsgZ6u98fVRZ7yma6A6iXenac2Ssn
UzZnfEuRhOdJDclR3Rz/vwPN+Iy9eUQTwvqvvLoi+0sEf5r70GwCyCEMpRsN
awNm7qjNHDzvwpg1spJMgETkbr+OXeABH26IaLH7EiTBxq4I3xbuQMEmX8az
yZiPosrRHDUc8xjmNzBnSfjUaB7x45+lBUlssxaeKmtlYyszlTJuwsjCRd4b
MOnF+h00hW1gAJDVnLsX+7r7pQ9DtK6WmKJ+0zf6uz/nTm1gJgOfLkNJkG1I
MEmARRRDfl2rknQEjKzkIUYcKjk/hCBK44zDqafr5XCK9pu+sNQf+Arbekf4
liilDX3D7hOu9QjB9Fc4IvSa00z6V6p4g6RFmps7ot8cwtbeCHdc24e1o71P
sfT9j15Nk2v7/9HRj8/4F8ph+37KwXdrZsos7Mw/VlRts5ZO2uaflz8rKzxo
43yJCa6CMSA0Ywq4lIpCCclE+N5VQrg7gagt3dIk8elF1RLKhUe0QWY7fD9A
Da5kNyTeJ3Atlt86i8gkFyoU77JDX4yWg76y8wmxfr+NvVCMPzlbPLYsmFzN
Nk/4DbjBpT7btEC/DNYq1iTWBkrxFwscDfCg4Q2Oo4FSz76/rM/SDN746Mkc
i736mFY9En4uQou0iztlNnCIOnE+Wv0nI3H2cmXsbk40F8h5/ipc73Ui+nKA
PUii3YTbUYhQrXy7DR3oO6J/rRGint2kLzPe7Z4MqrQ+QxcYh1KJIQH/MW3w
DgRRjVV5YoekzySoKeF5rg8GAzEK1t2aknwnPq4ZDo4dTb5JqQmyBfT3JZN+
dBu0eoSdyLRiZd9vNzyWeK/qR1FFqfoLk/C8jnHG5TnymIwWbOIMq2cPPilO
ULXDWaDEuLgOsCy4+oesNle/Wg+Si1/qE2ZerlCWxNxiVNmnzJ4QtRAQ5ZMf
zwQjw+WnqdCze/gI3DNtqpIZoMG7hwB96kRRPykt/Vo8eNhkmeLsODQKw9fJ
J6sXK23w3r+Qu0AnTrr3d3wdVFq9ZhFMMSucmp1vXAtmz1/zCsPsPyty7iDX
XXZak3tDT76nqicZ2SiR/MtiUckn8cd9P3PKA4eynWqOkksw82Uhp+/wx6IN
oLfZC0YWIiJOTnH0ooGfAIfpl8Ys0XQhPmY8ioQqqucIVlMTG0wjNyHHA83M
owD85+aRgi4g8lTRtVrfGUoYSXGSxxGrOtINq9XK1BTx/3yHUHgijorJPgKT
7GjFH1hc+PJsd0DQW5GobvhwlIX51Z1g7s+mYQazY+2quG4CKXbj4QNdwAkF
n2aBhDyPnXE93BEODopCdW2GKMBHPvCwuC9m0ZEnpaYDslybjl2qsKwgnDfl
B3coXwE6jdHunacuIZpOWDJVdPrrWoXNyy8OYgXEjMsFb+s+zE9pn4ywP60t
SfhfPMTc4TYbQ8MTmLjYt8g1GBSqBaZjhc0EXcZXf8AOze6TeXnHjljPRZS6
1i7xA9Ahbwzb2/ux3ITiiTatLm08Xf7i3UY+hNqE9mQuNR4pIG47naCVvFvA
JL7x4UmtQ9gAltCSTwCTwrb9aKrmWyMq/v5UHPTTsBcbwpXKNIFgVHm/gfkU
qW40T8F/InvwnwQzdmrFiI/z7nQeDDVRMIXB77OFOXbKHgHM/jbDb9Qm/KIp
7pLDxKIxpH1WjNpL+BPQKQXZGlgmtH1rxo95XsWe1i1V+kUuNCIGr3gfXJtW
ljWQwb+xOrJqVgjYNu68YuHRFuiacComx3/JHbPYQJUZuOYsDRkwSX6UWqqK
6RNuNdyX41+VIQ30GWZro9R+90Yif9o7PQQg8W1f7qt+90+MdjaPABduA764
+DPME+xO6GxRpwvYW5Btg3/JvzvL/jwt+p2LaAbWJmDc4m+GAAz8hQWFZLQs
Pp0G3Ykyee6kO7ugYNXqdBKxoBv1BBu4CeHBEAyxuiwIA5tgyHuDHFCoZXC/
zDsP+SUJFXKkCmYIFIb4RZ8jukph/6N5JjMpxxZ7zHBm9QGuJot2tTzILXYB
VXi2iP/aWlMvHQf8LAfswczaYzh/Z0uajwLX0QObCOK1V8yqqkqtmVhO5ELS
wG6T4xI2HziqHHpD3BJI6u2ISbUSOxXUa3HzA9WrpweA14iYHIt+cEqdcWNz
xBcZ6pjB7UoMqgTQMwzfbGNgfOMaRJv9FGYeXymr8qm6wi6ALiELlLoqirAN
aBkSMnTp1dWdQskxTxakB2mQuUn6OUr4KgMlmtkmytFBVKShtQ5j4r3ixQDM
m9JB3pbiAGYlSIoHMh2KrHGhL+Ga3a5KyzjrEcIcGYmKF4eVY+Yqnc2mBMJ3
RiMuxeWxQVkxZ+1DceifAuH3lnpoecl0Cc7Mea9bGwJc7mcSdRMDIfZd3GZq
F7c8EmbNXuKMBosgVu7SacEvFVIZOrKuCXnuy2lOu5u0cjQWavUOphkQ10WT
q3rB594FmMAo+0l0DzIc4j653eakcjUs4nT6GdiHK2N6n7gilP0vk2c29EPr
zVqSJZo/YjOuJXz6kTVspVhJK5DVg87BOU3xgRtwmAbWlbyyZmem3hmn+AUB
IAh0aby0tX3219T3+ILJNla8XQVp/IAKzRLEoadLN5y88+Y/D3H4bxqrFuT+
OogznYt8hZYvqADrvdV0EN1f7uom428c0Krlj0h2GyfEKCiOGUMQI4Xibqnr
nwAc2C8mtVPx76dvYZBvBq4pQUiw/u4hFCaDduwEJ6INOqHngBkOSeO9+h8T
c62mbuFQw/eyUiD6n/YZfRBqeLmlmYhwU87DVs/tzQclqLXks/+CqQqt5jtB
2hPSvq74i7CZX6VILM4Q4A2t/usOLSyNZ6o7qcdm8MFwz4pRiKQOyYRgjHuO
hNns+bA9HmU/+Vd6/YoyFCaHaSoVRSlctMY8J7LG6Kqyx8yM+7LweiR95fr0
m5J/pKkakLn2FnzragArzws0OM2L0Y+GmPpjNbONOoTfwzoJRXlWcjwGbzgv
21EABeYnJ2H//4qRvugkOM08STGHASPgE+e4CUPMVJmYfXX2gMY/kAl5obFZ
/SSW4/iiRvSLHqEeljHra5lSiKA71KV2N6ZW7FSVPcXGjYTkdx4HKZBxlChf
gFqyqEPI38EzGG2tj8g03w7A4Len9TVmerD4XsOYfh6Ia+jy8XYoUBuokV1R
nDZkK0iy6D0EkyGlEQrQKaznF/IAEfDwcTDxn/0339gNkUv0el3FbnWvsFTD
MLB99wnYL9tGTbiAkb6xS3iOIFedmQb472v5qLDJBgIICd8z5th3f6CQ34zB
haSQEHnkuvHdfo/6vRfe1UJBcPxNO2c4Juf8GwE4tEpuRNGYRkfbaqqLyFHZ
iTdZ4UWdzt9eBPVTDTuP9lAzGkNE3Idnmp7nJbLzpUY/8GScOK3h+9De8vuS
IdOzlOo6v0sAAStqN1ttuvWJsyeCniVt+GxoProRLkfZ5isXghVE9O0gQxWU
f15jU3NTdO7GTk9wWQTuRBfk7OIP+YwQv61fwSmWX5qFSmlMFyQwUYB5zLzn
9fkCFgoMU+GIPl5EfSUgKLwDyPqz7RKr88Do5hxykMbQlS1BsZiW68u1pbaK
vMXPZzi1lNEEPaNVSE8GV+HHSVRGTdk54YVB8zzaPSiZY5dMpxhASS7nNFY2
3/+K5o+q7hGSFvQQzzOPog7/gwyyor5C7m/DomNCG+MlZmL0oPyXgGUMob+C
/YivCD1UI21yiotBU6xSceoVUxLvhIlcajEsyKIBhm5dyuVrCUQUXYmXGtib
kvdjVmCKJt0NYsnR0YS0marnIZyKLbJ91xE5wHOjroNjbMLbVJSAPzlnab+o
nhGIevIR9XJqlFKAOfn020XPnvpn8fv4nSkPD2YWSVM2xxH8BM3hbIG5kcDr
+RxkCbwLlUo1AjayRBmM4RhvvCsXlkA4/owkfygUAPI3rc51jSZxpUpUTnD2
SmbsLD5fypwdfOy8DVFkDXlRjqfN2n/Fyx+NosH+9cuAmcFYqwz8UHdSdg3a
JRNIvrIXZes4Bktg2e2BdOO4HG7bznqlPyuJjYZXH3oGVn5FSMEiA+LmwmsY
PQz4XhLH+6U4MEbZZIwsqFo7lqPl88BbV8U04vcKmN3zVFaA9C7D4/PlpgK3
pKIugiNn2gfrJwOo/qluXr0cOMnKHSQ1MrVCtUIyvx3UjM6xOMC+FFRLn5D3
koWYBoS5PYEWhfGG7VzXwghTq/IxhrcO2MVnOQVaRwOBSn1nAB1AkhzmKwEK
4FIjBpnA+gYlbhzvPYWqxIVDpDYcLS1ah6NEusbh0zmDQK1cbkWFZaYTyh8d
hRY/lpmH95qpzgEjCb/+izWS6POdK4hQ+4qvOJ54E7QMsx7wr5epi4MizN/f
MuvlKAlEB2c10Z7wx0hU38eIZlCJ74wxVhgheWAMH8OoJZv//ZxsMfRESFax
nATHy/6WEdd/R/yQi7Seb0i3cWQSgz64WNeXddxXJ9KXVslGAYTdfWCpwgnu
XXafBdIPv3pcEhmuovREegEZ0W+L3WDUP8CDhxcHdT+9o5c/MIz1iyKa+m8u
EkFLbnVa6kwd0haHS4BNFlobGZHjzvxT/vJrvbRqdqDnJNNRUH2D7RtTSSFD
44LUMopkw1JVcwl+bDlZkrnPj0W4Qxx7kmdwe5TG9RB1U8luIIY1WUwKSsTU
PvKbqcphXifTyYivjM5+CPpFu0OmJcicZogHOwni7Y3OlQAh7mRzsEry1ZQj
eISM/FfUbZjmcARyANTfrXuRZoJkGRMmofjvR13qfYcP5/qAJsrdDlzYQkj+
Z0Idxry3PeYe7xVBfVegtIeieydtEDjXJlhHF0YU2b+Q+e0mVdW37WcpwGqC
050SuT5Y4RooX+NHIIGC0j1iBGzZjnHdxsB2hoXSi2L1rSWq3ZuScAe9CNyP
o4uvWK0VZOVufmB10shOI+RS7NrNyS9Ua07AmLoAoKoTj3iXn4UCSo1bAUPo
t1THRGi7G5xTSrJIoURJ4YirxEPexgwtKDP3IwZc61rdFcWdUMzvK3l1c/t9
ybdGrLhqaa7cCSK3ia5Pau4KDbzJva7jjeSNjmJG2xmrheNjAEjTLevP4Tha
I7021g63kx8x/+uy+cd3HaX8uX9NPFyAWDgmxGMaVauUBdl8Xry/AWPsoX+v
bnYKpxC4cfHUC553cr+3T0A4U33YYFIavuz91v8L8WH9OgdZ0vXB6uxpfroQ
7OXllzID3liYh0Q4stKaURcMfu2oDZYyM94VofCRFWjE2n+EtnGEWdjaASu/
KAAbFHf9dy1Xh4eAi1F4yCxyUtDZqlIBRKbQErq9yDiz8s5yt1K42aKHVNxR
zuIZPbZiVpNeBrAwgE+xGHBWxZ2N2qeoFHWATJ58LsABEu2GyzojehZY4Nau
tULa0BUxUfLMb9vy3X/ASwmvRAnmRImPl0TDa/FlQRll5imNvpvqx5MNgJFn
CeAQbGKT7+IBUt2Ppe7T/pRMfqWseVEQAsd/q0ipLqlm8fraIAbnQcaZV4Uu
ah8an+rfQkJtV9r/zewIPnspzyW/FzLQY5vYCnAFl/nVDp505TJL948hP9DU
nXf8a95fFb0sRfrL667aos2FGtqJ3/yUZGKXCa4DWV/DoO2pJGnARJy+Z4vE
y7NJQdM=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyJHYP2MEJP9VwrhcI/saChRqOIyyXRdQC+/+8Zm6/v97BIAtJ6irj0IXxnCVeNlKdOQ88c+hudJvbsNwbdXcjiI2vLL9bN1CPB1Dyv7u4MaAu+WaxJHtJSrXbcmb2n/hCPrVTQTJWtVVwpr9/AobsFH1jwJpwslAMKSXB1PCTlqilf63qh9PLudFIYkdasC3e4rOgFuBPAWWAdWxdSkgf8Tkqv0N2NCyoNfH1KQzX1DPvC8hywGg0jGNawm+lf0bcN/7zqrSAfzsY0QyFH0yIoDDlH1cHrYF8lifFJfzsEGmWsyLqffgSM3LUyeFI4pBhMCzo7lhKu9Wv0na45g2pJvVwXMXYugOeEKAzjtEPuc+38Rk9cq2XJYftbLF1N7YA7bpeNQjOYKS4/sVyJi79VB2ST/CwtSeHtffoNZVHERLE7x4/n+UhstCK5kQ67XJ0Q+m8jFkvJcMIlN8dyxWHZtA1klT9vMG8fhc06DLeg//roPOxbXvVDpS4UBh0adHF1eOsRMeHsk6kQt1sCRnEzsBtZND4NgoOEHlE4b1tgl/h023e/8tRoZyRr7+m0uUEG4s1QTh6iCmBKcGFEDc2Hj8Mwaf0z/cdMku93BZJMNAaWmGWODIyyizgV+TKVmBwI1nmp30PDkEIiMadEmLg1pHS9vqY+Rd0r4I1BTZlvrpzH+rhoQdQiEPa1fKJfxEPGsRJsmj6VDbMWg0VRStrxdx3sg4izKXvnv4N7Pk63xTh1NKe9YmcIX8MOfo4ZPZB8g4TUJ3td2HoaIl7yJTCD+"
`endif