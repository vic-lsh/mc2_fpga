// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
K5jJeIdC1Pu9/GvXrl6PZZc7eEjr9Kpkl2ZhW1MGIHXbdsbW0fy4GNeHl7sL
ei46ytPDU9xjVqmgKQjF7l2TvhNJZ48GPBqg3gGUEn8t5mPbtCBYuBLbjNm7
lYC4o5csH9m9pmQRECOwMoyLY5u8sTw1oVXsqdr7wJw962+9JBc2E8jWdPpy
DnRNPmno1EAF07SvRD2mNo5a8r4bvwk7LrGvwVaGMuAG//vOVeWvINZXTcyz
GE3kBpp0B6CVRzZr7FdFEK2nX027EmIAbFcS672K0Ej3OT9kLAboKH4JNduh
Wh8cmxsXJO1NL/eKVmd+gjYJiXkQGWAhrpsAIjwM+g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NYNAoAxuXC4BQH+ppCX2hs4XomzxNyxo6hbQnua2JdhiDHZ6Kqr6RSLNpsK/
kThKB6ryvmIuydKhzdgh5lvu2UAiiznthsmGYO/76sJUQ2nvXHMHEpacHGen
ToNNZmqnVo2zhuyke15YG8D4o6ucUOLZ4iVt6y1NTmj6k8HMewixQx8ZO5Iq
N5Sx5NjGUIxXqUGQ3rQ6PMIGuT00NFWH0Nm0jZSK6QkT+NH3tnMPSzhWVfmH
M0Ol6DFueCk0DWWhargRqMeyIOIQYt8VpBJVJ3gkgmG/ckM1H6AqzUXbVmiZ
VtgYO3vEKNviiq85VHBvbMqKuvhXgFV3mop+0zVGrA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
c/EFav7axQVsDQI/J/A9phs+ua70GwKFGNeP8wYsn0OG86tgUIxZ3VkgQ1Ml
jauYFLwpgP65c4IGQVB9cgnZKg3csBt67qwyfjNA8P/1sdBi9Gokk7OsCXJB
8GXZs/6My99Di4ffVs3rHeDr2fXebygRzqTqDRi9CL9VKi1Y6DPCtIa6idUX
c6akAW7b0S/kEtXYb+PgPMGBRgU8Lj11Iturp6ouiUzynbwWhctWHDcdUzZy
On6W3OIMb5Of6fxJybNxkmKiMu9Adz1F5gnF7LKsHqCtO/f/TF8/78RI3DwM
N87LwSfg30ml/FQidNF/282W7RYc/FCv8BoXEI/uqg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iw4uPVCM0n/kwCQxAV8BvIBix3pWU7739KGrLEgovx1Z6OgXD+u7J1l/OkpZ
qwAo2T4fOSa2sl+78+L2bPML/UvLgRMGSYgiM/vr2NI7O4VeGigfAhbERX3w
Df8QNvMu5foDz0pVtKbeoS/6Vor04t0L8klaXPmDG8PeRsmc21ZQnLoLQcST
FXtP+Hv9hvWwzuFqrQU1+Hk/02FVBYTONDCM7rRhd0eb0YhpBOTvxm6GFNxd
ROnX0NICzVovruLZJPUce5r09neyPRcXl5X1SsAyFyze6NuNeE8M+CnP4Uav
oqIWKmNJCew2PX52f+UZKDBHu/gEz/BUkwIikDLULw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DFGLjHV2gexEw7GffTEdNmvVWXslPjOZzBhUndEGAPKBURyeEDJ63BQAp63M
DWYZeItv6WjhTfb9bC+Q705wKO+Xd57+zmGm8KISCr8NBDI+Q7V1bh4jOSvO
ec/AdU9nRN3XBUyiwXcaTCz2pqg4RAfGxXXuabPn+YnWtnU5rJo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
vwQ7TdFfzdxr88nh/qyW73AewZKafGZx7JCJQT185TMJGTSVqSWex7ytEBfT
EA+0v0MTW/WZpdRQlU5RxwdxbDrAGt+TF6Kl1+MTORjmkDoVcbM6TQo+Sn1r
IIhiktpjYU1DfCwG3nZKZiKCfRryicC4Z/JmqSdZqMPyrIM/gK2a6FbKt8FA
kCl/eZKzSJH1vG00oz1PKjqcnUQeOsClrIkDzrfWMFbZ6KrIgedawGpzqWxr
8nLfb021Kr37TUBTImZxXgZ4TdT1zed9CAtGMFhackGpBKnIlkxng9nkvS7J
xhxEd1zDnqlIRXIKFVOWvLVAJeFqxmCMwbRzQB0mBFsbQ/LiR7R7KncHW2ki
2WFrh1NaniWEKe7KQScbnibYHqarU55rM69pU9Q9QOi3annN9twvtXzSmQDv
1nzCBfhFDBh4ACnYmwtkZhHBY4+RORzx+uWfKUPpgRpbo26zBCDZPCnSaU3C
FUKSPUGc4C3gVScb14LaqCtjmuyCnAs1


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
AjIAwwJo0a901L8E/v9GCQAg6pj81AK9TJjPwvadjcvyAFo4a5oigchCbRpx
Z2ohbkYYUswoRjE7vzRVvuT1eMY9VzIzKPk0xQ16MjkiVV+EDTIEBfM/ZigG
v2O/qrhSYSBKM4f9MJTTnG0a5UnIRUs3WarDAow2ZpkbUoa546U=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jQ+/b1eRQEUUuHUVBcMvSSpHUCmVuMMMpP1cm1OOU6a1tpas+harbg7m25rg
nxJWRM2WN59EzyJo8E4j7PKK+ZpfQnefM21cPQ6YHxz6nlUJitQHOEr3HbYj
QBR6SJCuz5ctuc7qc4LkFyd67nGBG5O85iISyMxuS3rzG+iTAIQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4064)
`pragma protect data_block
3So6DyRK3E+AGH1PkEMVBml19kLeItD1DSZt69PP/w1f3/36rBc225DmZWBu
OvCYBUmA5LwHfi4A92J1wk+xiJW6QxTRm8yjG0HHrL84waj1rTiNZApRq8s6
SyXJqUxx2Ix43Dv/ueq0eiMF6ea54N+sLHtiNzctZME0M6BnV4N4cbu0mUrV
UaX0ajKEQzaQLehM3p8w0KcSUkQkAQoXp1gnmqvqmQDqZR3ck5ztr5mwyMK9
koLjDaCtAWACY2Okz5ke3KU2UBvGPC+RTXgLT8rHOCTkUhT2MYIOFhHllFH7
tKq+pAGbFYDBMC6Dd8AcvEewCUl2cZ7TOmnBx3Y5Tj7tCp/ziWu3qVpZOc9i
MILAyA5UOEhhI/bVZWhpUZHA5Ld71mIgywSFd5z+EZGsU1RvgmuQRWWm5a1n
ZgOmy75v8os6YtuNziIWfJWHFCAejAb88FTle+LPJDDAWj240bZWKyq5f/4j
jqD6mh65TQYX59GnnkD1G48bNza0bVaunP0pjUa471WLKZ+emGj5hJjKQJ9N
WrjhvDnfi3fCZnBKQhwKMFRSpGF0xb65NG9k1PKe0xOgCinxocXzTv/hX+uy
AzjNYYjD+QKCEH/ul3ZupH3UlycmBuebCugxoX8GEEypx7ZaTc5688q82fOf
4aGUJE8/PN2kmkO7V3kTFyWRA5VCOC7F0q5SPM2XRIUUtM9ryrqQ3aFPzFRs
2VTKAfSrN0V7tS6QdEk61uzxw2PYfMHPZzmiO3bas5C6gu7SA8MJ4ErkbJxL
MUiIvrwckWMzGvCYxvkHImunS5Tg8Zr8wPcqX3kaSsvt2Dfmq0o97GJG3Vup
JIV+JG2CwPKP9+VFQt/QPIqCh/OkS2jbCpY8f4JTcHI7Beveyj+lAdigrgJB
q4z/V7GcfeXygcyz3zPNs/vjI7jaxGLg6U7f6qC0LujRPNOEVwrV/6dMZ8P0
xixpDKtdNz65303VNyMRECMev7eL6tFzHPPYL11Wm9RqGmUFZHEXadh+OCIK
bfa0VTOkHXdXUVfA7SlpMHS6SPeyZstyjCuJ+lSPbeH7sf16VNUD8yqZxF2W
hsEPJ+fTHGdD41ifVKerTT6wvtrjWMRv/Uo7UHkaS0l9v3otb4gx9ORQFoud
/CYNzSo8+mX47z+niwck7g7WcSX3MtF4UnyLrdu9EOUhE3qbQk/gNerZBHgS
espnVYxt9WpkAIlCC7CcPR0HXTN7R5aLsUCm89BlwxeiBwLoxY7tjozshYGx
U3tZpEDBCQQ/ETdUFqhG9UHQNopXdzNOAMmC3u9FyGgujKIeHEh3mx648rHv
SSE6Qbc7UyYuA7YQEgHCL9ZZogrrYYoP5MQux6W2BALROIPEuC1ZkGMkUi65
dny8tsoajFnkuc2OndKQo5jKyOvCFHPNulgkk5xiIiBHXdKofs/jbMgZXDVe
ZW0KP+XIuR4mFoQpwRaeZj/upz6Qb1rN12HQgVHdj5i0jp0PkWFTYtK1XBFl
rc3T7rw5cUmfCcCu7BS0/099DsQxN5uaSwGsDpOtNHzHQewr1GVXyf2/3Gnv
uRjNBuqwqVkgK3lDPareJ/H4ZKhr+Blxke0NE6VCfG2fG/tpVEUTKA/pkKCK
uzxog2KND/+tqBV0/A8WMpVI45u1g9n/o/bWS5Wk9QpgfNEA1+36Ikd7u9Ai
mxoKkNxkB+pzz0qYEnnWxcS1UNwCpXnUzvO3laXbdTnWEb2AAFqL0SuVbDeN
E1hmTt1zzTU3Kk+fakwYEtcx8LCxGaARt2IlgVHMWmIEL2qW8QSjg1dvtsBP
uLUaUeOg2YWLXJn7LELhw4XUfC13tRzrAuBMQa/QtE4FAuTzbeT8lr+SpDqu
b3S9n1bSndHgS20pMzLmhTWnYos5ij6l9/J0sblTVAXeY2FsNyls0IDDyehF
A+p9xIxe30JYCKdx2+IgYErP+MmbifudfFXWtdV6y7EbS+GIgrNfIQ9Q0ugU
7f6GBfvK0K4Pw0EAqxSl22oD1w0qP36PHFbapqTf3zm4EeA5Ui668UOevGfa
8TY1bPREkHd0jwjZ5YZ0Y7+PoEUE3RVmgqVaMMJe1JCp6ZQsDj1m5hpo0EhT
2P7xivqnExztpr6w+EnCpcXXIwHr2R/7C67yRVdgiCPDhCs+vquMq+axJCIm
Kp9A3kADCWpwGd2hw1Q/wqW1Q+Vtkw3xZ/5wmk4pRI6JjCxN7zNgFN2HZDza
xvQ/JPQdP0UYRsQ8IVXBZdtwXWogsHO1K2+0K5c6uZRXu+DlyxkjQzDpYYYs
cxFfeQ48eXYls7qoOhkzbFeUaF6fxmExQailABKjUG6rrZAn82zo8e0pANd/
ly/DDLR8w1b2uZFWNU9LfzTZVY+yD+f5U6h9Zg54moez6AU59eCAQhbouZ+R
UMDg1MGe4d+2PNDP4YqWpk/oODHJ+Zx9JGIamYIgEsCZa2dKLKxDzj/ZvOYV
JihnfYq+u8Mz6oG3+PFRWICvSSLnm76vp/gFxVykXvh0e2BVamXus+whmCN1
ErXmCYEwl+LLj3G8fmevzLyNyM2nNRNFNhQ5jdqgQ68fkfYZdm2BQ1LZ7plT
CU/vao+uVzHJbXAWQzbK4Eag/DCNl8fcv5LA99NwKsAi3aD5jgYD6Coewwfd
BQ4flCpMw61EX/iI2rHYIg0z3/02JrZimACm5PcO4yYrv69IOloILGfaSYF3
rkigEcJ5q2RW9tBIbe38Lg4YObOE5FYdfLHr2xUy//svrYmrhSCfRvkpy/dZ
cVbu3coiR4HKThCHQ9tftskTSitnm0XDwGMFQrL7f/PMR7kXgGZviEfpiRwJ
GYDqZd1jaLcSb/VYzn4UuDBtb0daCImSDVkkrTSSzFrsMkzR13kZnyAKvKEB
bEiYA7HuXDBBUUHQa5MPJEGVtYraJQjL7sZI3u/KAoyvS4yw+mglenX1Zw5v
TvFc9XdqOSkjEF1MHwglz5/RV/6sV20CTSQ5BOfKwbBwJtA1sNKy8rGHZtsy
aocP+A8x6RJVl4yIPxFwL4nf4x3XM5w5UioiqEqSL8KODhNCHAxZm9nCntza
nGtenIcIcF+v63bx7BJthUG7J/vFNvLqGFiGTa5KVr7rNQkI2bNy1C+SthbI
uPTKuo4KLZdSySzn4Q1SEtjLaMRqbw30cKDBQnUeD/mx3dm9+JoD8eJ5WP3f
zSjG7qwB39xbTXFfyZufxPiWWsIaTP2jI1RF/Cb8Zwj/7ZT9mkyb7NhwsXAq
JKj7yKyKYDXnC7GXk1M6TFbLHBrrOuIdb5M27BUGSOQ/vDTmrCnN6Opy1n3I
fZd45pTAdsXWq1WBbi+LKnm41SK2b+jtpI5oUvkbP0CKakdQrEGwXPvAzuuU
U0DJDGpdmlnWTKEthxm889JKPPW9z8bbuR84PUNLiFGEDKwd0X3dl8jB8YLj
g6k9BPnUpk67j8MI8Jikx5EhMrqTNsbKw7150eImVSiDagQE/S8oNPP4Jkd6
o6kgE23x1oIvwkmFxLKeK9NFQMCKlCnakMAMs1PiTWAOHHYV11kePfPFaM9h
HP1XcxLUUhzU0qsDTtKGRgefh8oSO39GfwHScn/zgy3z66nffDbDmKW54MDn
Hm83Lwc5NlPgd5bLJhrdfM/7d/rZdyWiPI7e37e95r06cvCmNEVgR8+dcJ/f
xc8OBVTJwoaLTkxdnQ/EYqRglr7kR1OIwcQebl0GzpWrqLCrvHEfyrxiK42S
cDn7HpkpVj15YbxOpiw1IMBXNsgXHp+Enf17vi5KnHT+F1HUAY/1oRUe+2dP
n6p6kRlBjSlB601IlwEmV7gXQsco4cOnVlTk7YLrX/UQTITIxJMmBsJQq1tI
LQtpZ4vynSLDyCBVPMIUgDbELDhVg6RJJenx/rHFKe+eQqsoLftsPdV1uLkU
J32I3/nXmk8ZSuqpsv5VscfPTHexQZFC0YE1S5PuFqx1N5yUTn6x9dGzauNN
G0uv92Qc3ujUCG4n9WNIXrBVtwh6LDf46lrmoTNiY6U5fDDiEQ69w4GfvTyq
d2NtFLyqdr/ps6/ods0fmstLRlP7Jgnch9bLoZaq91cH2jE7/CoH92IVezLS
cdeQQtVlwpcEcKlV3rlIpi3+f0ih/dUlL+6qWegK0sNEO3fYZvkGHyird9qZ
aIhXGz0EdodruvVRHEDt9uFXGpcuBBq23yZNfloLfIBkLlVxhL6pmTxGy2yJ
IwbvLw229Rezyi4bjTWxefDqSQwDm5RdODgrpF5p9mWyCcWyqOtsdFmvRihG
Z1pKvl9jb6QsUOEKxZ3X6e4sAJ/OMVBHQJ5sO1YfBSGP9jrFtqCukq3/Gx8f
WWpD9fmh+nCACnQYvw9wjh4PguraFHNgVvLEU5wh1Fdg4vBPXr5VTw4P6eDG
7B4C7xGKZJuUnQEhlTlXHgO/hcN3P7GD/aggggUzWYD7I3ePRAW0ZJME/iBC
jJM+UXqqfo7GWisdB3S/IAiws2TxDJ73+1ZCUG4rPxn7LvRpIzf8rdMubvlb
EMcdMsuB3nA/SaqlsoAFeXZDXhEbehFGU9bKrTNfF1rAp4PSj9xhT5HwR3Yr
Z1kFPo3eHLmJryJAMHUbdNFLZO2y+DBfKxz0MWEXBf0hRiMQn25SgYZVC7mV
CmvCzj3EQgkFKXMxQk/StczFrphGTlQMR+sHFXdIZYoCTF7rfcoqWOAPSSwa
ojF0NRKFBNfadgdNqZ7cRVwwXnhcF1YPEmVaRequz7nn4viSwNT3o7FRTTNU
jEUOEDS6mvMaQGQ+iD/mYwl0tZvoZGciW01/PHrtSDMyn8AGqO1Cc2n+852V
8m4gNE8IwsXDulDp4dvrRho0z2+lXs9GIt1RqDnm7fBVU9a5OoX/MYHwyIWN
3YvBLPBY1TjfjhAi+0DEtPNowQVVUEIaw9QvOsH9qBc0HZIKPD89KD8OluoJ
Wk2MAqugZ1v1pvi19CNFWXu3IU6WUqADo9WIsFToVZj2nC8GqVPV2QNWAM/7
cA7Fvobw6n+Cxg/hksrT/kchM8CIwNxkqntAe2mF6biimcY3YSbdopclqAfb
eEyo+bgpsZdcAI58zJr5/X9XVcM5y6fD8ax2IKa1kTFq8USYX1OKcwsUj98L
ZHYuEANIZmx1X8qC4U92mZh2DBzqhxtWk4igDKNVftwN/ltCphaepC8fDuyz
i6xwo+qF7ZIwwn+taJ6FCfYCMjqPYfMHeY6RU6H+SMd+juGLnXyx40CorXUd
5J0qd076mRO+d4Dt9nTyTq7BPI3FjVkmckA6NSkdXnxoMHOJzVnw2Ze9ZJYm
a4wgayfKz72BiuBxSrKfM1bfXbqFjVbsfn3k2zG/VqQDHePuk+y7W6ilo3FN
7DLPLUd40cpF5V/BYMskduwv1RPzItFca9m2wA+zvYDq8EaOV8nScdYX9qLL
VYLRHylCWBeAi7U8pZM=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "B40jvh7ud/ahkCWXo8CJP0S9JYnc5+J2pwOdONjrEnmjRzb1YpxBEP/gM90XdEQFf8e+9j+GJABVN1VA/EUgHmy986oXHU6n9uJJjaeBsR8h22iSaiy//95eH4kKFakRZgkZDqWp0dX7AUTwRg4vZKk0rom9cx0xsiuc1Ki6fTzxDmmuuNW+yyxk/luKJogixDl7f05H1PhFx3JTfD9y6cRFGovJ+RtyYHOBbLpk0whSHRK2dYsZaAerP6d/76S/0nP7+fM28+J0/xrsSgxs/rcypKKVD+WBndfTyDludK7x6NOGM13+ZbWZLFB4DlXHVoK/dKgEgSxqTOd3BV6yAYORevHw3omrRndpZCdLiHuhvnT39uoIe+80PLelxOcqcNI90IehmAy/x4TxSt+kj8h/lXHD/hlJptWEwV+q1U4H1pVEM6NcJ3Q5gs/OO4YOQ0zYsKMnBT6CwWLVEvYrusd9+YQ6uXNkSxCuvhL5J6B3f7iQ/6ZvMtxh2wz+AUpvCmwkFnCWzpKTLhytbWbUHFVUk+vmgURPxdu7bwCd9RZ6piTjrb9m7YR+w0ESdXJki3Nh1/YuaZOU8O0Zwr+Jk8V3wj0lv3Quhatb18X3tAa6KEJjJr/koREvGbkEeY0iZVKTCoY7b07erSj7IK1vI6Sw4s27LD+Nt5wUWTl38dmtgtS4w8nxOjHBe2K2Lv9Gb2Y5v+PD3B6m/iD6CpfPX4EgpFifL6Xj9TCyX7u1eAeFSGnHp2c/IVY8gvIwX2LzVAPxkCaMTBFGZMjrAwb42H+95aNR94QO+RFffXoqx+u1QxVQIaWVxz3QLL/d5PR40pVm87jCfpI6KG9XcR0U4i2qJrtDL7jbBMns2LBP5l5y7UvbCB6MzmZj+fXUcGAoz3io9i+4NZ3BTXVWisiJ1MuJeFr0bh8mE84o3XHYgW4WF1U3dlTaDSynMhQZ3cHjFVdUWyB/3kUhr522+b14Lu1vnACFfZINgensDK1On3wyHO3JwKHH6fadKCbcl4PU"
`endif