// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mhiA8otHo2OTym0FQyPkuuqgDfjiAh8oycG5rsS80JXC+JGKqacZpPkI0cbz
NpiNo07Yoy+RfL3TCuSVfJpKFTwf/2j1k4CarFSsd05YRw12/Wj6bQnuysmX
Mxgd1h0nC4hGzpHoitGMU7GL++ChiWyUQNzS4BiVhFZ9ikUOvf8Uve7m9G2q
ToSddoC0kfaKuQX5gjyKuYAj6dH/hUwCT/X5KCZcw7YN9OGUc9npCxJ0aE1E
hA0uTep5VgE2BEdnwPyx1DeCF8iU5wx7pjcfWWervxaMxF0eN/xA/4qOD8DJ
FzwBwBqeG/Q6xM6+jtUqj0ZhbNBcMKIS7nY1Ne95Lg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WZzPRHIHIaFZj7q4tpezONPw62pO6dxNauTbiDx95zefED9UQK1rIPm8jqG+
fMF7tFfgqgyCWjhn9f/kL0UxT30v/t6mbX9vw79fiB+jK9krXZL3rzdJt8af
MWG/2cl0KKTmaEGs9J0d9+qvxIqrfhEo7ztoLKM/hyEdt1isl0QZWDHBl8D6
Ah/B+oWBBRCor9EoGV1cv8IpCYUdfFD3RUc5fSCaP+1a3TcNZSLSg7chrvvz
irED1ivWn4wQcqbcap97Yxl+acCaVOmDGcx+4iQZBCjdpUo9DjHTtRuzz0jz
TNTTB4DHnXiFLgCUhNaegXzeGnOvqgGLVYVo5M8FIQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RGR+Kz37g1jPG/+BDm1KGbC6jsU6SRTaeT+6m/2MpO/2ZxDLnJoC0vO7TZdf
xUSNBtohueEq5ZWslZHodUqjDFBw8Vglf3OfesRTN8X1ri30FTAYBZa2eIy+
1kF4GRwTitryA61jB0cVtk5ibAz/SMasDx4AirJvs0iFFxfUa/mqNrxWXjiZ
3GYBgfd965NFQWGT+5AkPYKPkS4KPtJ+2fjkV1OO+jMTwEYCs+BVgdP7G1wM
teJ/ofkYyfHop/9uMDMxsI8QRVrs25po6f4zZVvDoMHCDToPk42saf0yMVlR
CemUbGaGEvtGw5p3cL8EkSF75gmeNgOO/ZI9WO1CaQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hA3aN4gSSxStgsxZCxBfV55trD8G7qC7PZKtFDGQtyiYLbWNE/xQEoccXHcO
QxzczzB3tR1qPQiryAe0RGmcxnnAEfd0s1cIJFFHZAkW/uP3R3gF9rz+W0w8
5+iAGg7+JBP75X30BGE79FLEOC5/VQu73c5+c8echAdyTBdoJNWneF8aLXmc
2eG4IRNoFd8sJxi6wwwzZxQErfJqfVfunuP1U9XCLm9L3zHZhm52Kt56TogY
Vl1rBf9Wuv0cs/OA9nK8tpmMsAR/4Su3RM1Dzio7GTNwRvezqmbjUcLxddVT
YLRX1AV+pEGtAZr8Qm3SG1O4AZnAW0e+0RYPbkYsOg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dyaJrSr8irOzZtxERTHWAgYwjmkIgBs0EGhCV+t3zcofDHtQr7i4VMd4XDIH
RiY2F6r9ZSFgxyUVYANdz8wT0T+LB/3OqpVof/fJh6Bsf1TcW95cToiqWtIC
5iQQmUD/xp+0ESF7Lwe8T90PLUDrCdXkBOJLKgec+5f8/BhXVjk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
HoXWVIsllLZ9rBlPtHUm7/vqHKtsvHLv4KGTtno95YojLLh8fTe/KKSwYb8s
8wYCog6apbX4kdl3WzPcwg67qT4+fi+WHdEGEVgU1Ai21yzYCHE1vDjh2gNk
Uhs11ER8Nb5Vrez4bpL2Cxh3OsuVKZ+GY8GEjlmYqDPRCPqaNHEIFA0QRvOI
kKFoshcGKxuHi9u+NfQjVx1j7JHf3ntClBdMkvFWZJGkILz2PqzKvgT2oeWh
ENraZgPapqC84vzc2mZlU0aupbja80boUuHFlUG8a9V0WZetYT/fXnXvCK+w
M9sqGDBLsDaB/IWrzFUVixBqKsAgVp3Zoor7lyQUhVUmmfpWnXfKU/ePu+U/
WyUwBpFhvPvY9Zfa52AA2E3TXfRF+c9lgQV/WbJS7PH5aRHRdCjBDIphwwdj
Wv7LZzNiHrcP2HQWvGZE9af5Pj99UbGnUbiOxyr7uEw/eAHWsjLrOvJWi/tJ
m+Y4WRvRJwxtF0dujn2l3EMvkQoyAGoi


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kwTfPYBZDsxBhYZaMP2ECzEraSZri6OZ8ppYJCmbWyKQLPpGfaQfBKSo0qPP
RBNCHrgX97qDkHUWoVl6+J1LmZ947LTIN5OvGQOOyeIXc11+jh5tRSiA58eK
Z23eWzlDfr2v2J/R31fLa+7oYbHDp1kDmDY7IK1uun7F861AB/A=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pSUYURQ6QU88OUO6Uq4+IyY+GqdYgsKzHzN0jRfO58oznV7MpUcwBlcTzlre
kVeLqgCnOiu5UX8NzmkB+cfwUCYnJm+AjAj9sgZpq0/WZyiKj02/6EtBiz5+
aKmKNpPjwnh0LDPcntA+92HmYBB21F4RpJWVqfqy7+efC2pKITs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10112)
`pragma protect data_block
zqSMPPn7GuCywVp8BBEnUSa5Gnq/o4i82eIu58jm5EOt2j7I0NCU5NVzHocq
QgnW0KMUNs2D/86JE1RX2DpWLZH6/i25j9x5wdupKzdaAQOzZ9ceRsV1cUkT
Xewdn1zYrWsyNq35Oufq0w3ksYpOghpCSxCdoez362rmzKF9G6oboF/ZDLxQ
mbxUoJ5FS7YA4o/DTXjjjYsmlwH3snpu4DfBeGhgElgSssHlJGS56ySfEqpD
XeGz/S0hOD8rkRoGXggEbWISAWyht5Ho/f7iLqrMxEu3JsahnIXwpnNoqvaW
YxXIePai+coamYWtAPcxMa7so5ce/HtKhkGHyEkt9n69Ko0RrZ+phZW4pP3E
iVUn5nbvMjWjdgkNigH0UqcSNU5Dhdxl8/bDp4Pcg6q4r+nxjUKsR7WIva3S
vWG1CiLm8hA8YhzaydipU2uem2tzgkS5L6DzA+PdFv/Q+b2mkehJ74hEpOKN
+iuG8aPK/W1KLw+cvXn5V3ZNZZ1L2m5xov4aXjEJFIHA/oCb+s9eWe4bz/Dr
TyaHeTPDE8/ACeSwJABFkgUOgZrp742chMh9FQf/xbRJfyua3yE/NaZ12XqL
EXsr4kKVr/KOZmAF81rcYSU8biFymqGKjVSdoVHKAOqyvfBzFm5B98zq6nBm
n6un3W9SF8/M8xNtV4LxfZYX867JAl0DDQezWGCHPwtwaotbk6lUWWYPVgS7
NKBsns6rWdIniKp9sS4xIh6wt5np4XZgG+5rDBLERKEDHBBc7KqsuWpkaEQZ
+wjAW5R7KDmYO85ORhjMtqx9thWLCbb7rTUeLGh5ougLX9gjYLi50sM0MSWW
S5qiCDZudkMDps6R4RGUUSbGwLoFJjCSYHYKKtZOSOY9m7Ih7AyyrnlzpT9T
EvZyHl3q+WQNSm9f6sd/bf6VyOw+IRskjAJAj6uaQDDSWst66sn0+5+3lp7y
PLLDURv5hk1NWB2+ZimGKnX1ov0ywOzKLYEXPQBFM/uayTdxPbSn55dF6Qjp
samtR1TlGxvaG44P3Q5PqgOOF7kfF1PLGnapgPtf/3hlaJD7QHCaUdgPXrGJ
/Shf/6my9A6mKsN3K7oDJAxxf9Y4iQEeEehyh652iNlTcTq6NCwUWfHwFdvW
snPX//b/zcQ2XD0br2jmfjLU/7+C9JGqAbgcw97KGuX6tlc1KdpfTuGPj6Ph
mthyPUqCcbkQof4ovLOaO+68u83Uarz9Sx0DLYl3DiznTobB4zxv4XqoV+47
jN7E9Mhsxb3aLMYfjwA+IKbm3rg3pX1DWOuSsoThh21otZLvv8KqdZXW3QHM
OOpHrrpg+fR24PPBci88SuwQzrZF5P+Y/Zn24/qokH4nhzs96LlPCY1nyUo9
4UMbXhstM1Ica05TGN+bZLJa9YIUKx+nB1cFgdq7xun5YZxoQXms+u5MVULl
8U52O0XIU7Mfog8w2kGViWflsGxD2VBBMlr5lu28oj2wlP2G8j1PaLNz7Sx8
ng0Bv2sy5z15XycVWAB0gD1xJDp+IpXO7OqXGROTpElN/UbQ/+mynSLOYY1u
NAYMHJUWt17zasWgbr8xlQmPGk9rvf4sa+/cdgwLuesYouYT+knFauBf9j3F
7uwxIOShiuHwnUcDvvxEub36Y95u2wois/f7DGr3P+R2g55v/U4+XNuE8iAg
NIvAFID656CqG2VO5XA9nXOvECwCm2EHIYeOvlKuPfTmvkYSE5cnJuxjcXqi
EKYwepu1Jc8zEKpvZWIefBICbw02lFll/NlduLkSHz0YSw0sK3lrtC4x3map
zQcED1GDrQvP3T/Pr//8195ZcqjoGHqFMLB45JB9rBu9bftExAH9FrdxLh0d
b8hvTK67i7qbvkY6dO73uPC5SRVvJ+ev+M44zSDE+VrwOb0DzFNBXm3IT8lE
l06KGsoXCDmlShVRNFCFehNApD0brT7MAMxHoDSvZU1qBVKdoOAh5oGvf5wv
7LFKGWIisipLTiwcSKCU4ZC8jihIr9qI3TS/NW/2b9jakPKMueucYOnoK4cS
uF/Seh3zMOtvq91TfrUijwE2DMKZ8IVQlPLqO6aQAY7mXrETgyncl0eX8xmQ
K3ITayqu4cdAxM0cL/uQ/DGyxTwphxXx4XI+RZ1tbzk8rngBt+aKfLPUe8SJ
ZH50UMhbrNDnt85b5C8QdMJ9IAO/D8mkBD8qnP7GoREbkurMMb2HKvjVWTNn
RnLwuM+/WNPlLgr64YxccAzpLAzp6ymHEiNEpG9Kp9l0kToxIvBFC5BkcFaT
bokV1zc4toisWNED3+Me+gTPh1qnfUvVQ/ZiNWkV9EXONIwyJUv4waQTNldR
T4a1a+eBR94PR7ru2ELfcT227ofegJl38g/nVsq1VIaikdF+SWhhMgjmNZNN
1KyzgVrSOmd88Z9muKlHkgsIZNF/7MwTFsJfaQcoXzgtqzkvkn6h2TcSF3r+
GYKSxkRGi2AYCQZ9SgXhBT/vmxVvjLrg7maOSzPoTohxfdYdvoZ1dHRDfsYu
nNe3hGmE3MWWywx2mREHn+aIsoeht5kn40v4g5Z8flJLb5OWdUrYsB/hmJF4
XgD6AsXWX/pO+BqN5RuSlnnIzxtzA2CWHjMI05R9Xd1JVtdjnx5lC00MQn+z
LitQJgGg/180S/ecUzfazjYQrGAES7AtyQp+5/ztngzMhFOrL0fW471C2CXe
82Om/I5Gk1QNFDnWKRLUDPraYMg47i7JsvPlC+ymUDrIk4pSkIujiCGEwg+q
ivmvlWSw0oOcLWJTLmeWEQoFugm/A81l/SPhOuhbLwmlQzjdpEeg4yk7s53q
NBSy4a5veymmW3yF0HiU5n4fx8/+FyZcRBDnawIYv5126dWs7y0HbHyHmUco
Jv3kqG8BSEwEN1DyAc548fyIkfT4ci03VD8CE761VlhIueJh1nBwJuWVeAi4
hvzuekHG5CXa65asmstMOu2CnEvx09GexFGvesytX9sCtzt8mwO6mG+wJvMT
DfTUU9QAwt7pfpeeqaS/xibb8YLjOLxAoYvuKw3lX/96Q2Xu/Eqj9pbf9/My
KB4v+wPpQ+Jmc6g9PKTsnlJOczXTy7+avPhUkE03Qe89cOj52FePTJ9Q3VH1
0fHdf3jaRH321GJw9trlj+UHhZcX3d3OXNC4wvl42lUghrLzvEuIQ1CA+3PS
3FAJPWI/0KiTTL4P7CRtkveM5Pn5OjSxDZdzRddwzLhkBny1YcArh/Ua+puP
NrjW309d9dtRk35jm4k1yA61CLppMoOSJVTU7SEmaN6oTfHn356uD5tzpxzt
vbpCDj64ffFXoXbyCSKwSjaJjmR2Al/YgvMlKUvmX9Q1hoLmGyCXHxHYD30a
JeVQwdvsbBitsNKoUeMXZ8HZu8IBBTcVCrZz+GZwdGDbyzDdr+hfnmBihaKm
D23COfImaBVKJyvDwtyI4hU6LBKlZ47Ipj20hiFEeUA2WZqEj9IKHHLEcGaS
/lDYXzCgI0osSuU6A/l8EJrQcDIqbK514Lc9odq3PF2yT3WZRqqlNy2fRoHc
NThh7r/7gFIpgn9Gb6ZLQ379xUUI/Y69RSwCpW2H3u3MeqeqWGcfYLnYEpOx
ZlpzkOobn7fUons7KQpyL3XQpgTdi4sWwCV1C4HxD9pupUOpsEMMkU661ctF
KWQgft9hPAMmUHLCs3g/7Z8FWOJDwZLGfLIzNsri5khn1J4wq/gYByYgx0r2
fDxFTIQGSqdd/l5M8PWJtzdjjJLc/OsIeqLE7ICg4dzMbfwtVCL7H3IdkFSt
SS3INPDy9Ay4++nAlyK5CQx4myozKvlSSObCNR1KBJ5Ase4zL1XVnfDz3Caz
MeQPuywc2yIUS3k2KIVc3z3Cyd58amDHtTnX20yVnuEvJvhh03q4Wn9NWtAo
/19lRyUo5W6CVi1tyGpPByyOvYO05L7JV76s8lnG+pG8/4PrFZBei2K4hcZ2
iLbaZynndVhwsfN1oECckZ6bOQmu47VH4Zny5szGbjt6EtdQVWkcvW3kNeX+
1jjsDZufhZg0aSYfrWRcHCyI1e9wxsYmZTL1mVGxfonM7YvRyyJ0NvNtRCHC
zPE1lYODPes7XaLXajA3tOwKP30s/vsFZQHCad9pbJCGWnot5slXR5LRsWBV
hpsKmJwMukiQnNkihxGaN9tFtK7rr9Bxy6leOfOo2oTLXi0NpWMFQDHApJm2
X/Ddl3q8EqO8Cg23mL01eNJN2WHjShVeG0co1Vwm7fm+QMEsXf9MS5T8vlk1
ub816MwC4kva6pWX/GUNVJoq/bnfibU1lklZPjmKypo3k7m6EUagH1zPNhmk
ogf6mrtn3RTOkTXGjmGicXtViQNZqlULFU6Drhi/QRBGl5TFVztsYsD6OrG/
wvGFur/06e1Ru28htYEotxjUmLxUhQl+vSxuwq22CV1s5L/1LOpjHW6zmFnK
d3JsIzcIeUIRELZU1E/SO+UyYmhdNbglbMK2goa7MvY7JaVptqYyi3KIGXbN
PPvQqfmPBaA50gI6sE1EutDZC5ph0zDhmjouem8B+1tVktfwOWNlsi4Uj4WP
WnPf9yOBD2mJwWNMTbFTU5keQGwFYIJmZlyGUL+4AAYT+9Rm2L3kLbnYVE4v
QOOYl0Ca+ZNJyBD8r2T0nL4IM8uAz2EaRbH2/64B00i2/RBFSO0u1KXYyakT
VWi2+TJy7N8BnvPaVHPz/pH8JRJRQq0R/LTZGx+F8JMJDrxmINrpP6DdUqDz
p2SaCqgXYjtRwhKD36RUD8wSc3+Dxm1DNK4L3ZTph10hacNSkfrc/8gXUeEa
Gjd2pTtwc0josx6K+A8hNw26RTvXQaFHYxn8jRUk/v36PP1ICvM9VFSEQPNQ
DSrqid2E4OnmDW9d2qBmCrPgNB2ke23yh2q2eQ0kpQ8VKNZpLaaCA4zbb8KY
45phQshX4SwTi4HLfrMScZCU5536iI4qgp+/YTtWVqs05u/4dItuPYRocCIP
WSvUDSlVsvttrja4d5vNhvRd1shpWB0mJ2+fw0eEKnvGDKIZdqDxdGNLWPJy
ZsjBQw6viFMJ3kWZv6CqIzWatE1ffV0mVQp+V58Jlt4uFC183BxxJpluZUAJ
uhmUfTjsaEVg971RbkdwrObp+dixb6lAd2fHeKgvM8Jyff2jv9c87d8DLfQs
KkBuoPdsWFCL+FYyG/OXOTmGLnHf+XayvrXGOkCIJdzgHcPVlhUYCvoDzJkB
S5effkPhYnSc9lFQtYVl0oHm3EXmclDFKGthKI5PYUMeD6y8rVtW3S7GnsKo
0niKeYSJ6bjR/BGh/gHF5ENgPvnTSFPn5ER7ss6FmakbJx2sHB1SexOVhMSm
zTPJ7qU3Za7SkpyH0jw9u8knMIoG94u8Cuq8qpoKhGMj8rNHbkE6YTefsNGM
H0S66EtKpHL+0qSnlw3Qy7r6GqLmJ/MFxxqZhim9VkS6HIAulUKHJWcvR2xz
ZFhqSTgHtvXwQzjqCj5Rl4813F1zVyzzLwo4HPhUW9POT+Q4C28sno1xHsBo
e226g9KZRXAjiWlF6Btbef564yk+FnfVKtaTeMXdHqqXXLT6daG2dG4VU35z
Rv/H56T08D/zhWDpwWBpLJ4MFzD2k5Lu7Bm3RcpId9SS6laKYzvsiJgWApwG
8CzPSQvz4+HusPmeqN2JUgfPCDTwZkw50mNX4D2vBKTiiLXOFM4i4Tgd8KQ3
k2off/LniJ+aDmOzCtiRDPzO4jMA0d0grnqRSngpU6XmYbC6NQY0KbpUH6Q8
Z9QLLhJVx6Py2LZcX47Rz+OhDiDZ76pqJp9NB0aEy9VtVMT4xpiiotgKhBq8
jOjRWX9gwQjUu4yeGEED9nP2eBcfyZdaK1jcDN+H6M1xIEqnhrxggbuNvmE1
hVXHDSYXK0jbypi7MFqrODPW0gQppBqV67LBd9GItnqESwdFBD+bP3vpVWXX
b9rodp43duGTV0XHhMGklaBqvQsCSEImain1Te6GbFkqq1bVIqJsxbj8C06k
WgO5Ty/YSXX2PqKVBoHBej6PaFvMPiNE1reY2yDcbnWqGttMsqVeiVJhyhPJ
8tXSXYVasxRhZbyAMAgjGoAMyljzsy7/AioED0XbbBcdJvSbDYrYuVuGE6Sg
RwpmUybpePO2sZa70gNf38tB6ZfZjQVVadBD38YD4T7Nz68mqNVU7C/bViec
uLpKfU7KDYJxZ0y2nbB/T6dsXIyARP+ubO+W1DBq/POnuEQOWMycKHMYWFme
C1atUHcPxKAPQrxvmOmauGgoQsXNGfjW9XDAZx1AIRfZtG9NRnjRz5g7oHAO
5HSas+fTuJsSnGcsHRm3TP1wo1OKXh1Ufqr48WG0PE009mlys1cpAZ/w2/lm
AigJxrMGimOQX5CNOJ2BD1aoHWXHRrQDf5U7pI9GhHpUzP0i999S0asZ7M67
rjljqUMjzeKsgzJk16amMtJNGqP261uGenYeOHYL0m5Uk/HMkOkSzxH/tDJo
km19MfcVd9GjYQT0WJriIk3sDT4+NCfMK+WanJpybUC19o48eZRCX8ha/MXf
8+v1nyiscX3PPZHyw6ow4JKiR+dYhjv0zTM3dOQyPe/2/FSP9pvzhfbnrNAr
Wr0GjpY6teg+JFTXSSsk1rBkoiUFwvO4on9MSRIWB6D2hR+wA/VDibCg8vUL
a24iJLCRCBdY3fQJ/CM2uOlCIM7mCa7YvZde35vk/m22A0V5dHyD14LIvXXF
ou3hsmdlb3/cFZGVeHFjqKN0wyQJVAFrs7W3snd776ejap1o+HoTM+Qs1ZER
1Gs+mv7SLULVnwhzUUPr/yxbUsmP6qkgKsXMPMKtKzGpSwzAJ2OJAYRdWUvl
jaMh6EzwgOkehSKPkFa2U11Znm8T5cQ1xdTEsr5q5Kz22vudPyRkDK/x3JWi
go6uVY7p1s5O3zGHUqH1YVKZwqt3p0bOx8zmH/io8Gx+ir7rSwzoDP53W31d
0CK4I4FPKM0elHnKnJesBeUz/BNjDBW0uGE36v875ovrRh6AUpIHQK/MNr+2
X6udzjm0cviyFIDvtUn6GHm+X5j2+1lKfh3nJJRC18hHH+zULgHTrw1cLbQT
k9jrMbUbq3LWnqwXhqaL4A+pWRKpRDthb2rRZ1lVtMFUvgOxAqWIsNhllgN8
zAwofxrkxRDoUjbuCTudh7FR8yhMXbteNOm3KT/cDqpLxZIPV3wf0ws4JE9f
qqH6LDGMBudGDhgxnbhPrtcPP6WlHmirR9avDRFIPR94vRai4ZxiQmyqy23a
cSbHz0MpNNFWVQTLte/IcA6pWb4Vb3t0lRaXaQG1EYg6yglW8G+lN7slnM6Q
BSSA+twYNBSbbp4Umh1POVnl5CZs6u+etFIvaxRZHKIgPCB9Kp7yLcexroAX
/5vK/8q/xEFOUhmO2fjq7Dg9FF4i1z2gGtpDmxdRNveVj3NNJr34fOAEnOKG
bzJnuOvBDkGy7MbJlsAj7aOMD1SM/AX3vbE2vT0Yu4jT6aangfzXXhKrAv2l
E87HqwO5lTOZ/21AU9I/hZFnFMDWpS+GWLGeBruprktgZsiBEje/3YD51cR6
Tlco2ZMNuGaokA5ZrqjAyC2Jbfo7Euyf6iNuDGV1FRB5Hpcx2G9pqRXwGyHC
VlwMOKzBwyMga9T5Jul0p1VKb6sYQw2l1SpX7nhZBewIsKY7+SwXnVZNwOmy
NO5h+QIVQ7vnKwrof9fs9PbNFg9XJAm65WIBXEg9hyYsf+6DWg6GrS+cOfAR
olZPmDjxSAo/rF1dXBnhj5dETcyfQBihx1SKhDCr43UiMUXNhzC9Js4t45FW
AaYUqfoEKrwQrhA983lkY2PrtM9QGock3WxZK6H775w5JHRAdDx7SxSLx2Yl
9YrUjS8w5cT944jmCAInG3HCapGOb/ORl2JlG8k4IIfDrBbiUBBQQJNceE3h
U67dBEwp6gQ6ybZRdpz1nS9kABv3AvwYQk5DfLQrJNZ73Jw9LuayBFzPmsl3
BORvsm2kUKjfC3b9Gf4yX8HXmpUck3vvUhCSPPkegBQyeecbEPaIQegWnjOz
gg9rzqBTXoRNZi9PsOq9XmcA99cjTu94B5BoRuWHAONcwKa7sO0Ottr7GFth
PfXQ0i4Cb5nJLzkS/ByYq/qCF+zqdaqKw/aALiuHGORHBXuxtDceaVG5G/1F
2ydndUTfGHBVmGX9QV8yopvoWX+Vcdoxua/raNE5f2wR4P0nezIL6S54W7Ke
DKt50zBi8Qw1iZ931TONUu5BIv9RgOw2c69GZiHs8EobHOZPLKhqPGF1aBjF
o9X8IRapJslUtLmt8sYN0GNjE3myL/Ze38P1ZTEh/uK83F6Dw9ksz2vkMRFP
87ieZ9nSRmkXkk4OBlsmCgUqWdmN9omfBpSkKinuSlAtDLp9sc+Jt0C8ZFQM
cGhDXhiUrydihhIoXiIE7BsaQp7dxeT7oQuF5V9WtYwgh7JSf2wiFiEpAwZg
RGXZznad0ArKcH2idx8/28CZYVJAMhWAssWF1Ignuh7clbhBKVegoJjV5gL3
GxIe2y30cDO4+8ZGgnu9b+HjSq6i+8heSqykkV7SKeF4nyz2gWpraj+7vZKB
WUMlC98Lrm+DF+w3pfwyGjdzTHs8dRe4oIjiS05xLulWNCImm34vIDsdNlq6
XC4yVL9+hqBvz9F2Z3p0XSj9FFSubFRVTj5qx193QdoTIrV5mwPio69DlsAv
WdXxaTN8V9ecoSGNKno0M+5vg6GvlP3s2sJVZXQoBLE3sy8B8I3oL79qePeV
Drm608PWLXDPZirqQP1fdLWQ70buiqvQbOnnxQDW6fzXlomUclztBcLNZCmN
px23oeaG/iQoJ8wSJVyK8UspmPFwYg63Ui/QphmVESN8jq49t0hNwS0yK4KL
GVotp/1IlPFLl0KuywJZ1WwShOOcePFQLyUUEW5o72ruWj6ED6XxyDgmtkY6
htJBHxKuNX9z0CerUE+F3KBDUljBZg665fZ4CpnRgSFWCS+Uvtrd5ISnTA66
lSrrJ4AvfwzzPkugtX9Sy0tE/y4++RGMs5u0fZUgjdQgHDUhynvbrtpnR9+I
J+DqYbWrR8Fo3GheDpptpli0PzENwWeMQziKZylLziPoVAOraTzGaBUYJ32n
AaFGbzj3QeF40p60jQpXsjhckeI2nEa10dow5jAq31DmTcEIgfiBICqPa8nE
MYK8JV8rlxWcZ91qV//lXW5qckG9wYZRpvrtReRlaSfeqVTTedqR0Y2+/Lyn
ML1yn1yGB0UAlpcdd2UQHqU2v2XX+0XCY3goF3ZyRQagbuwolJ9DRO1nDC37
ec6jBhXhIKKuK7ll4Geq4ytWTQR0Pj1ss8ALRXFWdN62IIGIy8okLF5RN5Uk
I1f5WgXLa9hxtm8AOplxrbzOhK0MC/LmK4Bamg5p5iQ9urtsrC33BpiBu4Hr
lhhFeWR1uAiBrNgtXB+xW28zfkW0wNRvoIdVY2Omh0NiC6fQG3WC9r83xWe0
8HOR3MM7Pu4Tosw5MEZ1gSLowT/74oI+u0+7R8R0wLUvslAi4LOcc9lVzWGU
S2EsJ3sJ02iuafQhsXkAHDGJen3tZBfWuH0XV7nOXJl/D2RRQKZxjhgLQqd9
tQ/dcWC4qSDWEwFf1UxPdT4jk6iyxEyPu4cpzRqj0glhJrmg/N8skjzLT97W
3q+KN38UR/krADXjyIfgx/5wJMUaPMVmBXvmFaH57U22F5nHJY5BpmPNqNUj
1/+qv+O0wz8FdkaffOC0BtQYrHjsvVZvKO5MwW9XzKnoYtninA/A1CGse2HZ
HHTp472kiJmwp+yDTUWqFrCDNL8/7nj8FMMWriopCD60pBPbwxlJ6CmzvrLe
jmOq1Nu8ktuIHWC0MtboMkTaQLoj8pTVDR3Q0REffeLLTmwhFC237FLgVq+W
ZK2lNmazOpKYK9GhnplJgKmSTCU5OOuME5G8XrumRLIYX2hU7M8YpSi7bJIj
aTHxTi71jal/187oN4L4McVKsUnADp0xNJ5S2luD26Ew5MslKQukUQToYQj8
SdI2v0PCNtvQirUuIrAkJSUZEhIIAglwx4iRFbt/HbYd45HCqD/Y1WWQqz2I
n4R1JmzI8cOjrsf/2UD+T2tI6ROzC5Ql9PUxN13PGO889P0yja4d6lFuZEJK
q0+rMqncF+PxY8cq50ySwVQfcEtvSVMWWg17p36v6DJ+c7C9pTwG2r+CrIgp
HyLt0PECmKnvrnqNL+7vX4gAePFZdAi0faTkgtO6xozLxOGhf1afhqWq8mv/
29GF2BP3T0cvvJ8hJPKnzKLeMt25MGeJJDrQGIOE0NMWZf17ZEyHaNWI1bmL
nvu+htLwwaKndvNGNh2I8MLKy+2D0mU8pUs/eIqV4FvlyIzd3I9pXCVhAwCs
DKYC1hyIDJAL2QOdG66j5gUsquUmt+EYhwyBQ7yrMK8ewr1PPXfvycr7GSL9
mafITKDuqXcPjeofEjZoBrFX1+PGE6bvRlcSOEO4rnU0Ef+rR4zmAu4fxxg+
/K2/o6Vdq+NkTNfI4opZuT5dLUax9S93EDz15oKqbs6GZab3+Q14AUWVVrdm
FSYee8IrSmODhvQEqm687LPVKFc4ztGlt6LYM8A+HNxUtG+rxpFdcM8zmIUA
6b12VhsmD0vouBPIHMsMdSjnMQ1VjhLVrgDCnUYhTAIUbcL0LLw7cIox7tVC
fpYm9wJ8bAMt4pYfSYH2sIo2IfsLoi99jHSQXjQYM22lXNinu+QMVMZ8GZAh
V6TjNmmvxasOK3IQd3U98OZVTingxXaVdGC+M6YXXiImS5ZYN3D2wDnvJWna
y7hHoyPjuY+BFTtl8inTBdx/KTPkMQTbmTtu0W5DghzuVqYeObXCDoeZ4rp7
EoFa9lkApeppHIf/dDjFT9dNpw0kHKSPYIY9T0cPXkmjlUsLrxynsoQG2Z66
5mMcpSmfFkOfAoOEC0vgVipv5/jdcK0Qe58d5DGxQG5cQBlkQD4GWtWQ6QF3
zfNqa3pLi5fI1aq/WJDGQz1SzBN9WjovZwQTeWxYQEOoBxNN6n8Jhc+/hNc8
35kEA58M+F5a6OeyJXnS+lkr8aNajPu2Y3mLygP9mQvSJPBiy3nPcJM8iADc
d/QzFntmmLGWWpPvliKpSBOh8JJES1av97AKlQcz5m6fHXw/wa2lTQ31B8oA
8P8qH/n7RhIt8iix9E+lTnP/w0cGEuxEQ2MCrL27/DA5Ge5Oc2FtpTZGKDSA
tzmPugNBeIkZq9Cjpri7xlJ1Bxq9tfSriB4LBro3xva8aBWRMukC4fz3/qLp
CutcLzc/QKwh3OmY2tTZ/gtTlKjmav1uGLaGIGadU/ywUjhn2pAK75tQND4s
uHflg7Tf+mhNJO0mXDYuATXtXiccKAI7GPEA8vwC4sdCV5l+6rwEsjNDpJD0
HZ8kNsDhrUnvuRcvVZ7h923wZfU3ZhW7XBqoBlscbif00nsXfPCGrGJsE87d
MRAp+6dGlnJji+e2p8k0VCefV384cVYtH9wkZ3q40HyBRvTFzRrzaUjEnvs/
w+JyClp36xMYIBYD7bKK/CqXeNAWkw92GShvvs8Ng30AnjorypfR60JeI6z2
z7icCoOQdX3cQWsx8KGpCNF3BysXyg0OyganMKk8RKFtFO3jNiBiIxoQ66Tw
Z8VNTE/TRSOtLro+3g5hpkFuaTHvwr66c+vhQtFfAV77tkXXtcbaS9VAHtrz
Ga7yh2JTExIIlJ77PlOUQ8btnBTflulfW/btfkUaV97NgWzy9rR5c0KFX22O
2amAVEGIz9YU9UVVsOMLLWFYI2dG2fRqeRfeQzDz6PZV3bkm3eJOa6129fUQ
Y0/hjDRmngNQT9uChV+1OhNadydsFx1rG1dTGQ1L1MsBOspHAZxeEkk4PZSW
FmcTWMbvrIMksOfdyi7YOMqHhrgMIWb1EhSCCR9zq3tUilDbQX/G3iCzVWP0
23/qP3tC33+V3J/zv/WNEAUxWW2YCDNUoj9t7RTJ1Dd81ULmqPBV3vNZKJ0k
hbmUJye1YNLZGA07EnarGBb7TyMulWvsmAVcixi5HoUPAdKVPiYpA8KZwJ5R
Unq4Inslp/mhtdYbZlgQNDGoDbo8P1TRvO6pg/nJ0Av6is49rBZr2crmltGC
DZLLuYe8DNAzen33NOzIODK4B+C6sC1aAaC+d9qCvqKG4vSCweZM/X3wovfj
nkrE9sElwv6O+S/T66VxGg4YRXxx2T15LaIgm0sY3Vr8mlFDFMB3BxaA5J1M
McghswONNCEzpWbtdTbiEDfPAlN+i2O58HY1c3wBztCKjrZ6ZzmEKuiK9JKC
D0LPx2S2xOUJEfpoJJCQzEQMQQCLb13hm4r4PX2CSmJ825yducSh+ILsFOWT
ESQ/6LOlitTVnIyX5BFoLfjVhaOj7/h+ydwY9qJ14R8HVEAzllu2F/bdxaNd
TXRDZtkD7GjRZryuHRUgAA/fQOpdY39qDo/La9yl8ehwCDqq5n999NRk2Iqc
kSt7aO7Ycv6jHkCYlMEKq5r1MvL3yTKcPGJd5HRgo5/lf0/QzvSwhno0QYUe
3n1rJ5xGm3EcZL2v1qGITgSslJ77JuVKkqvtC4sWN6lovm0kUon4X1zzDUjO
SRiuof0IZj20vk77f4d5qELHx5TaUIomkYSDhrc80z8meZklGJ0KuIeUikGu
SJjKkhlPXXidBwPcNW5k+cJIiOcKs88bvdrjE9JAKwE6g2BMeMjGA3/AjV/4
dCYq1zTxLQJ2MmepT0SBWkUS/qWJvWb8mUC7r3jtuIUht3Sof6hGNMXKmB1J
WI5sSgG0RqFeUltMQi+yvdwXo0aS5wJX5NoyL6tsIJ4fTrQ/frXo/5zz1XLd
sc6pXerIAlsYf39pirV7r/eX/tlzDzDWfF5KKCgZn+knw9M/VIificJquDh/
cITk6H9FBKXO023nu4p3SjRlGrUaMPR58Az8dTT4tFhrWm6hv/K2vybX6xkT
qSWgTcAL1Hmw4WhZi8OYXyps8HIR+J1JmjzuhBhyovQB7OwE3XePd+GHC7so
vM0NKSgw5LUxOqfZCyaT+kulFxUbQKWpj5tP+Ik6dgCkOjdl4bgH3UNN0ePT
dD92rzSSqm1rS417MdDNxf8/69ofoPC024+atgQbEB51HOS86vtoWYBsdNGS
466rAcaSsaP917g6+smiGAygheqHijXYQoOFEKXgj+lyoOQZerZWVEmeZKhM
sStHDSm828/PLH2C1bBhEacsFkEXj1750GJ/Bgyix5W4V4+z2j1eceZs8Ds/
GO+kgrvlo8RIR9lLWyr3BwRXSc27U3hNySpnKqj1Ar645Om4FRMerEeglG4x
lQzr+Qbu8XlHGy4M00+vAcgglyfJbGiBGwKsK/7ugb0Rz2/iSpx85E1EGuGX
a9jUFg1fckoZYVHN4zYbePNeGNcROGFmlKAFv2pi6dY9NBgIPJDNiPw4d5hL
YJMhwIq8EKAURiD60tjPPNiZ5mFbFEEe3x8rJIQbV3U=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1JT2tN9iNsQbAdOxDd/VOqIbomGWbqGZ/gw4N5E35626G8Ajfkr+kz935PVGxuqV44+wM6avATYo8CNNvK98qV2nhQn1VFVOWy2ynCvW1tYmzRHkxxNUabcNB9sTg5g1/k+om2gA9Grmxgr7CApu227KxyjAYwcAmBo+8eQtG/vt0t7BG8goHoe/EkDqB+/eGpyxW+zRjWI3ZOgpMeLL1wmRgfq9zZmAzqN6NqPEuy+Ew0n5YNomVAz2SqsK07fTNopgnr2/mDNiKio2BtQE2VKbFRQ5ej/NRtFC02LdUD2Dh6ooP/BRtKKMJz8VEhRTL+1EYOZrXYtf9l9STDjfeJSPysgVL1dLY6Cxtol9UpQ5iAhFMR9O/5gb4CLNrCdJ+e9uW2pFvu2SOecGByqSSjBptkoOw6f5qv1Pmov5U8fH+AcnxAoITA2WX9NGNtecs3LPtbOPDUBlEv9NDkfzX7E0DO1+7UZLV1JRFnzszVm2J4DhR6z4Jbu9M0rze6qLBcINRfd7FV8fiZUfVujltkbVVpoxWUxYvzXWu2s9uB4g9RO/cqn7NL/Jd8AxFWxbBLELeabC0c7qghPxs5z6bDISprvFTruXnEC14uIS9xtym6JBhoe4gWVFYti0+JKYm4xQz528n6tmH3qVsnkiJYxKMHpFGi8aCkjkYErLUKRdxSmwQZlRy/IpF7y7fzSh5k6HokVwYhvlp2p2a3h+8MGWiz6o7aF7212qbpSiG25lXR2hAgJUsPbrxt1HEnThUoU6wJ7VR6j9KO9n/SkMs3Y"
`endif