// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WJb+P9lhiAJ/7psr/AFmgXboASrpFqkt6pY7k8hWJ72FVxLMMm4HdoC98rtZ
sV2lyN/y8Y05CqigHrKTZc/yFSsV5f4P1eXjjFwO+86tKQxkMbJPEkO3jmBI
LzxosHqL/pxC8UPFZHdKey9mQ4lhgAQUuj+OcwNqbeJY0AE6xmrBT1mMqE7o
aWXIDTcb09/+aZjXmjos5QZ+3ru/qADkJIPJFgb5PHb8lA4b1ldkJ/lrlzuH
bK25o7oSt647xf88irhCFO2PewODrwxff5VVdtE/TBoaWwcx5NNaGVY54yTx
PFl9XW0Uan6i8swAs3fvpVXnoLaICmkcAXP/m6e1QA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
o+x0l1LJIK9wjwokxHqCPPC8fjjiwOkz4wQd3u7zESBbLaRxNhy5Z3Fa+dIV
GyD8KRlktPxQ1K5o0goy1wDi5JuPSWXDhJGrjNyszP8iSTAh9vVFJCtCWqqv
UDjh9c7VtMXu5JGc1yfz7cuxVzivwKl/WB1uooSv36OCWgbpfmb/ICDqflWn
x7yoUmuDcED/Rp8+QrXWKHkSqeyfGmWkbhg5/qej/h1QUed3cdljcG06swrU
jfXjm1i2ZLt3I3Z7+5YABCsMfUT0tEp/POqrfdq0l4E2TcrKGxa+jcEtaCrv
11KRkZ4/nrzMF/fKof2mKS/zha0n8vw9i+WW1X0wgw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Re4z/xH/7kKibBSdfPAmWUKdUR6fLYRTx0wZlqxFW+giNT/sNw+/mV10uGWn
3trTuoTahJ2GeL9wnPZElmpwHA8aMhk3TiJg5R2taJuSyu1CEX7MZIJPm4LC
g9mSLIdLWTCwtggZJbwSuQ/8C6mmhMyiGqCDAOJ0ykekcu+XjyEIRhF3Xmvd
F35/n7O65nbH/wYJJ7kpLcmz4jfHP9HniFBs+HPOH8jRrvtEFMDN5qU2Q+dm
Qx+qpKEms26xoL0GgUfD7NO12fsknGtHP/wfe/1fLzsKDJ5upyduyeNfPLKg
eAkTEsXNLlfQU+YfifXyZAFqhuwvfuiNcT+sPcPrVQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cSVIeEl8CkHxmqTN6AG8OLnOyy1KGn4nRzfO6ZqfqsnbKXylYk6sDlbMBUj1
ApiBGbSsXeq1Vk6Fp5ZIIXnV9XhlJfzLorLGAp679iUGR4iM9qUtDbAG7dYR
c/Tlc311VbbAdI+iV7NBZsGF2zOHiIsMiB2v6yo33k2QJGT5ptxBdvpd6zYJ
QCoD4yCOSrtaf8kEzaXVUdF1yShwn2BoCsvZ4Jn79hhSx/lGntUgvAmHMgDY
0p9ZxiMJtEHowFEzOMKGIuOu7WH2vZwJmlzY3b3h5ksV9YcsUwpEdnXCb6rJ
96EmfV/aGMEv2IERNgqpzfvxBz1E8FWaV557i2OdZg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
F1Rf2gAv6LlS1gQpAZ0V7/U5lsQnX9jTLQlpOGfbmCR4/oCdgcUYTDOhCUU5
20aNRf3Q2Who3FFJ6eb35HpY7Fg6se1arGqxm36a73lYgUacmVDu/z3HCmPV
+abiq4/+WLJHvajdoK+05w/K8veP2ynGC/nlaK0GskguW8vVquY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
aOQH3GVGioaXejkNEh9z1efVz1h874aDHTMJ9XDY0k+YfLc9ZqrN+2M9mh3y
2WgOBYxnbRHDXrn0xWmLdHivs8YLq42UjrTKDehcRZb1Ki3N1pchCFmZ6As6
uF4SyBm9yeB4WQgWIEmVm0vxNxW0hTwEC8MmsnggxfsMCMEIL15jbsEIWd/m
+Iver23FnzUJfSIHizSo9GPJ7bmM0MX1Ruv361kjI55LrgJMlacBdoZ6p/mB
2sIHmu5cJb5Pa4sb7SkdF8q/95vchBoe1yW9SUSMyATNGbJjx0Gps2CsBunC
kj0YCrDY4i96LqXx7YUF3LK7CYa62+03axUI1crpIF0qFaFa+jmltUBLLpBF
Q+tai1BFk/ipM7+ALpWxG15j63E45kTgMylh3sLMTkbL88+lBIDet2CYkLqu
nHlH/S/IhcgvaRoacr5og9KO5FunpGyanpCnuKZAZc++Pnjj5LQbBLxSoESL
QqSrABcr/KZQo6eITNgUUr3gsAfIvBJd


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uyAKSksBMH7kCZPoGTKLoihMUx+EZgu+yve+jb72NAY7xMzHm/uES6VPWwAu
mP8P/QpJQkacH5sewjgWQp3IMDNQXEVT51LGLyBkLDsfFjwPpigAutFSOH0L
Ce5xMlTNwk7oErGsikMgcUGEMshEFfkU9ygzboLSZ3JyAsZ/SNo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tgrvXoynoSYB0ak5qiVgp8W36ITUqISwmL0AwMHsS7QDzIvKn5wvgLimfCdn
P1wGfIztECs6JBwvvdBEmh3MztLaqkxfkocBGeQoWeYk3Ui8jODDTcW0BK1k
99kQ0q7Sr0OUqY4aBQJNkbYJMkBoI+8NQfkrww291O0qKx5prVw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1584)
`pragma protect data_block
bVOK3yXfIbleQBZBCBzYLCwN6/NrEsK/wcplDq/nHMlfk9Hm6iZyoGkt0tap
fqHdxr+LUvDTJnvJ1NJUFPJUgfYVxkTNA4nShFGSQ8IvC16NYTRM5e63R2dU
TKieV9d3K+sGMkNIBizHHHggbZnI3ad+v6izHMsA2fdRYPunJTtWukMQhUXj
cOL0kU2c0dFzCVd7qrJjuLywal/Qbnr8enU6F4QEkP4V19trnaqIOVfNbUTI
9zA/bv+MbyhF2L+nY8VdarTm0ob7583XwmziZSAFD7BxMOPJbZ8mn6AoEFSI
W8ixt8LbV4wPaR0EnR7u+QI0i1GA09RA/+hs2l8MHk0J3CPoviTQVaQMgNp6
hrIG+PpmV1Q4f64CX3xxwehLR3ewfnkyGm4bLkjh7uHueiWY99BolPMivblh
oE+n9MZg+UfCX/Wd+r3IBU5Tn/hxjc0IeEP2ZYhyAh+SpK8w34zLZaF1y+yp
h4lZWoerXrk/yM6aDQQTCDsws9QdFRXvTlpLy68w3RmbK4RGeNE1Lrv/73Wg
HV3aKGLDgiIuRmHR3rof/zn9cAMcTphZA9RM6v2OPrePrpgP08wVrAz0Elc5
1f9Jx5WcleSpkPnvHGrRYkzG2Wu8sOoUaIWPW2QhNAX54d/4a0bwYgY/Cw9E
CiLowwBWmdvpzc6uCfLIDgrtpIYUV94/atCYMEqlthH3xpgm4vgYGuWVoB5G
l/R6OhWXAqAwZbvlvdvGA4WC2Oau4qQjOrVzb6mfXoN/dFUyvJrNt15k41Bm
gnO7MAx3Ymd4imocd2pEBXyAI6LxyLSFqjP7V7qPmI3kwNUDUV8GVO+OLNKP
GST0wn74zIBYIGbLSykD26XkAvy4+T0hMnzbnSh+5L5y60F29OgJp2v+jfam
IXW+Xg6Cc9hXY0NP06a59MxYYyhVEiG68729KAKgLuf50u/ZFQ59nnoMLNuz
3VHYkLF5zlMgKGcBQDUuigqZO1r4zb5sSAkqHCRkcMRw04Z6ybf0OFBNuXUG
sN4LyYxuoIgTsKsL7YVtBxuBIJ+smiToBbSqhKHZhCiqjlRVTCw2sROW0S+m
UD/eD0nOR+1KymSgzOFeyeq0OpCqOVz25aumdfB8F00x70CT+hZWduSTvKyv
tb/4iBDzuWIPGu66sutka8EzvQSjAsORtAdc0vTiu3yyOpMyOy+2YEGED3XY
WwUJOXFUJGB52+IsInUmWBrFoXPnvDow1XD9/Hn/A1YjyYNuvrWJ0xBEDdf1
FsIlVakTHSHjetW6OPMWut+XCgsTcSsP+/xeI4GBw64kPzzjvAWRufzTQwgF
iKC/GgFYzgJYiXTbH4AEfSx1Eg1oIb3ZjMMnE8GOXUUCT1f7UTS6DV5FS1nG
YixKRtXU24frwQwjTWzknWpoYVsgsO0Ol0DgIHxN7UXhOgoib3Bnz4y7/yMp
ATwByefZY0E333LR7UW4gVpz2y2p6NU02b9Sik6ZnTBzWPL5QliHJEhI1YSo
X5YMOTdvIR1FWgtlOQWgmGz+qlYIEY3i83M6jaWfrZOfYE2YH910WzEBl+Vd
/Zl795msF71Ot5Cdfv7jrUYppGNBMt3oeSY/xv4hJ5o8F4CpnEBqxsylCR+s
SY1ed5HyUe6OoCiLWkQRA8QeMFHt3Je3/UshBdzla/KiALvjnwW1aJ1AkM9T
eXMCuxsxbHso/TSPVmSpG1xqjRaMqFH5sCIsrr2OWVv6FlAfWPTDHumtgGUy
7HJLo8uPY/EBBdOLejdjIQrsvw7NL8iOoBDm0Nt7qNHqB/VwsIPRQ9XBXnwc
6ByUrwPfm1DjAb4x+N06FP3g0utJrxj6Vi1CQzdPKIesHdv+qXETyWA0zoko
1HztiTIfn/rZpwd90vVEHFuMz0Red1kSwnr3jug/KqRFVkWzycx4M22n+9J5
j6Lp0LtCvyPqH/zv7YFViJOfizCLcb5Ge9It8ttpi3iyRmIx87F/11J1R223
6fqtCc98qtwdeHLPInnf/EN4cxZO+DEYdxRibcXDZm21tA/eEN+eiwpqiLsc
C9ozsmL6Tfw4YzPXVrR6DvciTD8O2DmNWaBg8H93rrpa2izvIaYVayMrHchR
uf/Viv+rJjeT

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyJjGCcZEyuBpEdgrq+uOobByulHxPP+V7Keixmz2VYZD60Em4GisZBbqFzCJr0j/WGa7i9u+grDznxEpwwg52dvPm33caetLRriu8sY3uA3S5BSseQEFAUrBUkN9nilD5n0RXyb7XtJq3siFed7D3UXvWvuGuGQ1DC5q3s57n2WiJ0gy6FHuP4V1w1Y5ma/wYv8CaxbjqmytTKZwc6ixT8HR0GOOv3ZC2Z6wyOxNi+nFCi7sodj2xNnsHHUspxAR7vNcO4bas0fvajdgKuxHD/ibq4eb6Eg53HefpZ3xY6RlSvmNJUgt5ajPHfsuVTJXh1rOTIg6bgq0yyYyceeQNChqjtJJYnROd3g6lehYrGXPpTjfeipqVIYdTedF7j2Jh3ox0lwe4qgCydj8D5acg/upLC053UL8jQXirv/MS/j4pEO5mMxH490TvKngpmRLa4bXBFqwDQaWn9pGU8inw2+M5CnCd/bmhY6s8XwAj96MXSRcMAypBY/02J7F2azVMXchSbX/AQe30wW57i8Hkpvh/BCF3LgN+QqHs19mSH0YwRdnLlbv19ZlfqTtV9Oz6YCCBzOIgPiKT2ZBDGR8xsPIKKui4CK/3GSsdz4BiiPVPpUy/idkvjM47pABSbZenB8lCyOk0SGcg50jfL6V0A9KjfVvEChawJOxSODOmlhzMzK/q9zl2Kg8UMNZvjKVPR4U54fiKO8zlUhS76Yoiwdu+Oo66jWAXl+KUvmfa2o/EiQy7byhkdYKiB9v3+iPMur48nY2NnW1V6ubMJiELkO"
`endif