// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KxiV3O0MV9c/QRm7ShYP/mlmhH0LngbdTMaHPbxGD4IKZ38uZJEngrmp6x70
Omqud4s4n8q1JmUp7ObI+rYxQaq4smxOzrVlBVk5WfhEWwECYvTcSMJeYJrc
j5z/xkxCuZbvTiGpLN3e+X7TRwigsaV2RwBBdWnMiahVxxXSuoBKbx3bjEQW
uKX9GWd4CBLl2qwp9R81EAgs11caWWZimOAE1Twlj18HBqQEsqo32xK8pqlE
dT44Gqi/gPGjqv6RxQBJ3Knp/t5Pyi5t6SHW/JHhdJzD7hdUZ5dfoMxOTkLp
cfS1KLEwh2bLkSJkRFTHq8AoY+1TtROCteS54rjW7Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bKFcCvZUhkRkKd1RlZJexYfPURTeO+tznpXB/cBYVPNqPK70Yaj0vqS/1Z3S
TvN2t+hHDaw0N80bC14ROznwW17FQ84eeY3w//F+0y4+1x9ApN22Zsa/oDXZ
UwdrmynBFwaHhkPp0gWh1sY6+qeius3/5SwQt0CL5LL1enCkYTOcPeI4EABr
mAHRneggElGKyD2Q8sGQ60GT0pwQOMYlaTGWfrbLA8zs05wKzBqHjn7B+AFA
3EgP/7N94GbP+L+cvtKtHsN/1QcfjFUg7vAGnJxdwoUyE5b/kOj5wGIagc3S
K9mgK5mkSyMo2zFKWsUdr+sNlTb+Qy1OktpLcROwlw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
tDRbzftAinrh7qt1Zrlm2Hrfmk38joM+YWzG/iwDr8135YwVz10nWpjCdGem
2ls8WfzkpOm/cFU6lzxk6D2+bIaM0+wm++xnoZKPZv80oKhbbwcIxDNxEpxH
fhLv9LXbsuZc8BxbAsh2RjQ/HbPvC1aoPQe3CBpbBt9yV9FCVwkc1cvgU31F
OVoQlM79fkvsNtaG82Lxg4QQWO2xIIUE/HJ0oEWRRoNgJUjJahuv3En2VFuz
EVnpMNFDmCJRT6FTd6ibpzZliymLOWqI0j40aC6sN7vrtQXTuoaInNRQBSoJ
4+DX/NFuYNkILKeanRMt4EXZOkbkm2hmoM4uDUDl1w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EPBpFy1NYqEYWTpB7U9UTE9eyTmZ+OKCw+uzyKOmOeGLz01aEo9f6bs+OGVx
Cvi59ZdQr7seE1xhT5bMPq4vsBHjMsQDPvGLbz5MdT002Qsq1XbBOlaz6iTv
z5m0YfJCc8Cw076Dewu8jGX5U5L6cHUaFJsm/OXQGnbFG8OndjjaCy71KuEu
Xt2sR5gzwL4qCbGhOSUnNMthMZYuKVGVi/RbfGNQ0and969yS4LchZnolSR5
gYs09A51heTzImIQ4qZAdk5ft5P3dtETF8MBoNrMUvNKhxyozN3+OxhNKial
7Y89+x2fx9ncIxl3JatzRtjnDyiXSAKu7X3iz/kssw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BJC7EmsMVjdBgBCj4KiTg65L1YDGD87/aZpZxvwo50brp9Htx6164lILewzd
cx6JEux3vpWml6muSA8Y+wxBSHc+GFRxw02lxxi99Hb2IPSJSxFILdxfoELQ
BTR2+Dd/ZjGYmmHIASWgwvmO6Z7s0qA539ARTRKsSPEShNbCSeA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
NJdalSKgvcZeJ4id8XxECdA3I8O0eIef9HPRYFYmPAgcw2L8DsraHxVvWUxJ
zlG7DsLV/5H9kQjjuNN2TFpja3lg3v8ErVSoFuDU0YHP37SIz2GGf+lCV38i
IaJfMwmOS7eVQxwCS16YbcygnBueVYf4shtm97N5UCfHyEkUp450FIzCWyej
Ne8NibP3RQTXVMNEte8uZgCPrLY8+fEeFINKjEBA+aOM48Y9nc8/I5ZYyrqE
A1JUicTVTJUb0B59xmrTbSch2OpuH1DK1LEBdWO5tn7hEVQHBbTIvPbftBFm
vp3qGERVrYP/qsA6LUO4qJ6vY7uIHdnbL3hAlYEefJ3Vt2NVWIz3lpoAwufM
rXfG9Hm2s3JszNq3+2ITKIODtOJPjWSHcXvYWoDEGhz0lgzW2QKKniR6bvs1
bKUFEv6gyxO4kklZeg1b1F9Z/Rg2fYE++/qBQTNTw1JfxYH/AlC1nK40o0fp
50Npn1ob4onXdNhLJgswlA4XvGluvdmS


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
u7or7I4yVZAShURjpwlgSh7jMnHNoqj5L1XZTqIXSiEBKx+DywKwJfEj2KPm
3zUUMYTi1QUKOVLRkTgfcuwjwCsxBKxz+/pNHPHPxREW0UjVvYQiehoU+nvy
4mH5UUEkDhsg4zun4+4GIWv5HirohZpFAzoPQV5jLsIwDXDUeE0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pzZwQt9Npx/vTKtuzOHLyOyiGpe7d/6qubc1Cqc1cl3yXLixKKoqLToVXoMb
9eSwqTA8uv9ysLCBVqxukRf+YwA//OVgx1e3Dg4pqJaz9c7+1eCqP6zzF/6+
KX6LxUitQ6dJ6a42z1fdyQOAyegybfoxE4Jau58aL7B2XWnAlq4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1184)
`pragma protect data_block
N12qCFl83d2u5nhotujjLMynhAc/BdHuaamD8l2Rr+RJ+jgMoas81PMoFyYY
0ge5T8B2h/CEVOvrGUhErVVqBq403vrABDdoYIAdrHOTckPhmsT6H5Z1kHn8
tv7gO1aHVMfQ7vuSa6GdBFH9GQunnCgiuHnd+6dxtRbjIEmFzYbD6vCZs38M
PKuEu6D+qaVptJJAVBv4Rhh6eF3xFgN58iu8MdXOPPXygHtRltNaPb4sfeDl
eYEJTFVJ0vwfLLfdvieYSXv6hu86t22Cdl+Icv9ZDRfJuWxVRaS7CptHHHlP
xxobJBnPwI63wy/bWgFf36nqEhDEKDKuBOqtWIZACI6DON7WP5BNX2eNdavM
3ifUb+KdICu1f+YhzWHA88eRM3gugbdECwc768W/XZGcDyFuGP5EIG1JautF
bG6R/tl1dJ8uxUvzPew/48VgB2AULCdvB+253yrKe3ksAHl5piFDtH9HZfbo
t31Zxz0TznDzYBEcvveUouwfzuhDerJsIV9hetXX/EyvO7qqKrWnE9jtIhIz
83Zvs3G0XmjAjCiz2fL1ItOsiU+ORYfGWMNmRB8v31f4Ic2R7XARDlXsXQ1O
gVsYCcNlIgrOiendvk+JCDUM9qXL3+aWRBpl0gF+1EScbzTrvReWi1oEReg2
i/q1k70lCAk7l9nvU0hdLp5CpMfCpP/jqoeBmCLpJGJTqyGSJw8DaMwb+REo
WA30Q9wFHmbfrmgS2tmu4+EUQK6wH0ycLLpJ2rkEBIni5Njvow0S/TwqWY7x
73VTlvKPDIqfNLQuFKmsp0Fu9H42XJI12SMq27DRTBfAykryuhrF8ALVRYIm
nuoppk9xJIOtuW3ZbSNiVe+Kyl1FXSb3G6/etIAfFVrdvVnd92zrAMDegyjH
3JTHeO3pI9fFurqh+v//5DhN/5y41t8Db77ZKFGnCLTtM3v35RF3f+Cxs5gq
aO10kWMG0OwzLWJRxMHcQQXoIZ/lh0W4OhaQj1z17dl6ZvkKRPuzXc0AE37K
Ru8M8WG1KES9NKa39YZx5xydpLhcRKRH53w3sq3gPuD4KxJmTLC3qRFGm4ka
OaB+fJ47bUh4VniCK2SijbqMVzMefgQYummbgZQ8+2rYbOKoOoyq3Jo2pjuR
ZIit08/nlfA2cieOtREc/U72CQRu70zPTxuRB0+myDZO8M9ZX3KQ1cPI5N/Y
CHr/pSp+szV+MCz4/hZ6RGqjEMlggW2tVXQ+Pw/YuZVk+viMEPVJ24rqm6T/
mgyXH3lQCCy6pu4hqpbXYRppE7sWvd228KBh0CVNgDQ38cVj4SviM1cgoVth
BEnWGzZwQIhAeDmsElZ1oT3yoc/Z/MfPoFOiRADkPmvB8Jof2+D/Uduy2Iga
xX6kWTj3LyIYluF5W11Bbf+RkYVfhCvXAMG3oez09KERkjhZtwWr8z1lzeNI
F1+GjRXVUpw1MBFR8SrySyvAsB51oeysO11+2c42mmEsFkJddzyEmRYBB6R7
tqVsVVQFrUpwMpiIm9v7MzlKDtEEk4zm7LOIs18LH/NEX2foH8VdrfNN+3wl
mJrGN4eCicIP8RIDf9A=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqdYElYfsMAHK1qtZ9DO7ztBZbvUuQbMsekH06QuHu8SiU7WjN1Ht+y2VanWI0cKc0JgMmZ72cGWKNF2rsqQfU28tnsElxOM7CIV5dcjwhCJaDOyKtSqybwS0WPHjkiiam5VN+fuaFHP0Pq2smgFSCWBwmRriOeLKKYtxULn8ftjyep7QkoGyEIua8xUW/541hKnC83w+ZO1/1KFQvjh8pyKgHR5DWVSpe1HWa16Th1bgeOhIFUm6iYrzY2RpKgUImBT018ARTbiJxN+kct3ZcUe9R60rzUZS4bILYnvmBD+pzVAOXoTzsKZ4bo9L9FitHYcybOaOtSRTsOW6I/hJNvgp83CSG/KquDmcLscuhGDDBES3JWIifim7v272pP7oioLhlW/JGBHPtX07gyF0NCb0OQXc0jgLvsky4jmeHshRA1zBKuy66wYxNO+MN44+jgxcuOe5g0RKkwdCzpQDpCaNjpHrTW3cYqas+bD7Z/O06fmb7NhTA7U8JIG2b6C6vG1ZXKgh4dsIvZGFSjivC6IltMvz7LBnIz1JorMMSkh0bDxXupRXSCX+4GFokGagG9zK8freo3FI0bE9KWOecAWqGduRagoEmdgsOc7Sk4zZ/WC9jW7QED0pR9+4MB1qriN/D97yFjde/J7YeRqMWdex4bOOj1PYPsPfb4iN4T4To8/DR7aHunnAN/AJe5PUHBiame5PGTUhPecEWgADeHQwXcCnB8H9SLA+EqYJlovDyL0DZhJ0pFbVFYqjWGGgtQ541hWzDwm3Yg778jzKkQf"
`endif