// altecc_enc_latency0.v

// Generated using ACDS version 24.1 115

`timescale 1 ps / 1 ps
module altecc_enc_latency0 (
		input  wire [63:0] data, // data.data
		output wire [71:0] q     //    q.q
	);

	altecc_enc_latency0_altecc_1914_xfsfwyy altecc_0 (
		.data (data), //   input,  width = 64, data.data
		.q    (q)     //  output,  width = 72,    q.q
	);

endmodule
