// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rKAW53Jb57aWKs0+Q+6KgkPnBFf4Kr9JgyCPNf8IaLRUEvpLVHCF6BVnuhzm
KCUoCShzr1ecAoiKQOqsSIe6ppZdCSwp1zmQe1UvKXZ5NCeVw+fEh+s/eoRm
O5IY0QSQQoBMCbhBI/TJErwkpGg6RkzP43VlvUdxiGfDuYLis1naXhxQyK1N
E2P/R/pISjH6UZ5FW9qCEetZq6PRF3Cl6WBPBq0CAd1tundFOBcNCBCfHBvn
XOTdSn0pxo9t86fq8UdAuoCFe5DFw8ZwpjsTWqqoC5O1sC8izKHOfvVdAx17
J/xqNCmWoZQG55SI56du/2FtIPOQSczeilboMVeQwQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Rii6IL9kP43TWAhHG8+ToRP34oIt/gL2uaz9Wf2RB8+fkPX9QvcfwyBrCIvu
e0+U3ptir2pBRVllJLIQUa8WzBn0o/w/I1D6m6gfM5DskjsRIE6V224ZOouC
/NStV1swBPkhCy/P5XG7aCicq4wZBhpOx9oPiJ/m6BudXu4pAZXP3DyziBjs
/H7ZZexPnh2ZJrPxW1xFluFvXmNshRmMoJ8tYnICz2VWtsUwtxKPBhtv84VL
EkyNkg2+dyxOB85Un2Utgjhb10CIGDnst5qndBc5Kfvan/pTdFR3XS5hmNVI
fdSl7NA3kmffvM9/ejoj+VJRN/lNn5vIIID7C8VBDw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cg1WrFNSSxAOQjBMOx4J7YwqrmDMDUHGEgTC40es3hg1XqZk6/zb5tiSWdel
QKZj3S0HX61ccVFH653/gXdK2eImUjx5eQQ3QfAYRabTGeoyn8NuhXhRJvIC
J6i0F6Byl46UMjCVK9qndxqDkrcpju8+VPgvapsCO/0BEEKmcMZHb96XbEdR
Or2AKbOx6ipRizkb9QfdzFyR+OPx1cBQno7N8JzCXVRnsF4uFesHSoUuUMLq
HiWSgyMthRCkpLoV0GioXU3S2TFdFPRGoiQZfi98K9ofNkZC0mS/xCifDzDQ
vDZymNf4hTBMvDmRlMlOPYH6r8L8Y0Vru0ptxM9Rng==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NPcmo6tVVWk506r0HhJc6K2+Sk9TXoeMQCkfBRH8+AphMWvqWUtxwBJlXgMJ
gRUhUvCg/txbrwvYOM6xl3dejwzmxMD4NxYAMSaQwePilMzykIMTWZqKKLlo
/DMYfSpdO3wt8sbB4cbpf3M78BSV1XykeHj74UDNllsvYtLRAMASTxPgTH6J
buQKa2phrcUUWqaM7zQ58uMAZui3m+TwB3zMg79Hjz4Z2n9DG0gLyyelypy0
jFgcPGwtyW7PvEaeLGuUXaab86KqnEJ74qVQmeIp9oGXUdddMxo2pkhxu8kX
rsnYm9CeiQU7T674snPniUoFf7WxuwIUQZPy47xsMw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lnVLSDkxbjoWVwut7oecnUFTgqFucAHS/v+ljH/mJ3y0xPUuqrlZWwxjYix4
YqyttGwBZ/F19qFzgM2D2m72/y5T6Mih5s9f8Z18N2SlYPafBJTVV+o+2Cpo
NEY2riDvdy8nnjEh/ccktqz+TxHfP8BUmtG7tgK9vSJTSgs359I=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
GlHvfNOU8GCcJuSWradqQGRCFIWv/alGhBw2Ms98i26CkfnimeMd6t3qq4Jz
8k4Z34S9vFpB2u+RcEfHuoAh4gpPYOHdvysCZOIvxFe+oyUaxrE7319Wvgqe
nckfmWMyBYoiVL6yBrg3yTPaLkoZg95v1rijzpVOddbWYJinUMUcNnHPE6+/
3n1i9F9BYu6EwP+CMOQxxx99+XmHAFC3Z5Ik8YtGSS29e02aH+VsdIi2f6NP
gK3rUaU8kFmuX1y0NOzcL3cL/0ambo1lztUFJzIrfk4qd0EkdnzezEfkcIgh
r6gcFViPjoldZ+jK5fxo9RgalKE9TpCS0yCoaSpk1rgjdieH52FkxAfr5Lyf
k/nYtvSXn+kepvwLsJSCBnnUkRew6AOkKCUxsaKQoyykxY/fKhv8LAuoxVlV
+0rlfaIzTUTUlXkpN8dTK4YbM7AJo5Y/6TyUCjnLD9g3DkclcAL/MlsOYyPN
58xHGaO1VgEB6mEtKzSyMbeVZXhIIojY


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DwFDs1SB8OTQ0uQsAFWN0ln69zDgbK8USWa9pxVn3aOZJn7c/OgT8LRwLTmP
A+7lj6nElthbgIom3YCNKd9eySCtAGEcvIZYi2JIZ/UyIIRtKrtcvVw0NuTv
IF5MO0lRw9IEnJ1XCat9rPJ+pnr+IxnYLKS+wyRgyE0UahryoVw=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
J8hwL/cqACZd/pD57i+1+/G2RmdBRKOwgmQRipal/4YtQ8TZzxwdHFwYY17R
DM5TkQ8PqrJWAtILYjHkOutgyiHzxXFQI1SDiyYSXK24trj59ZV3PDbY+V3W
nEhWSvPlTmBlV0mGp4VqgcrXPLU4aq5fcXXi8bfZzy2oApVYgrQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 16880)
`pragma protect data_block
vKR2WVbk2eL4pN4tmmkDhATM/91wtYvkf02+QddhKskLZ7OuXNhCnXjuhJjg
Ko2y6tEgTr+UG4JJS7420yILPg8st4AlOX9zhBjvfPk2j+Fe3oaHQolx1YKF
nPVP43KatQCHrqEbvQBiYNzOLVFqnTGGAWBo7PXj7ZtpUpn52h/kvJ90E3Iq
Gy3nTgA5vPJ8iV1AyMue89qYF4Nu8DfLmrY+J+nB1S0lICQywo5fns/mWjM7
JPcP79JIlvljyTd6fT3mhnz2HMyK5EUUXaIXNwgv6L9XsKsGNzbNM5bbHJKZ
75iH8Lm2nWK5L02GDzTWls0ThE1U0v6XXH0PjbEgaehXRzKyHROyRUDJ+AKG
7KQzhtcHqgOPye2WPyzY/x2Qt1bR04OZAfAsheJIWxVFDYNzoOUKhkRb5Rfn
DhEEBASCeQXMjc2clEalHDxxirDrbe6EV44kS1CF2J0rgKOXpAyUMWWs8ppa
Ft8ilQVGy17ny+2yXwq898mHHYPbyV4/fSwh+kxjZTMS14DJkFKV/uBRd0l5
822F1VwSYts9/v/RfMX3MVCl2S2FsxyfW1bl9HvhPEMgyqWDzz6gtooS2mL2
o2zJGqXx3v24UESCDDPaGpmyF2UClUZyTwrR4UVkcCXro/goiQ0TyhpLTbr6
JpfInZj+V8gD+9xeCIkBmAlg0mquhl50mwkQXBiF3wEyme9br8kTjipOQtU1
Sv8bzcxgKKLwVpJ4f1skFOw+raQY1xJawjvkGKIzQWPci+EqvVTCfTh7WdUx
ateWRZXyMWYucZsTsZf0sPeBgb6V9F4UbUosWDduajOWxxqTabm3yNE/6VDf
TG2hGVp4EC55heaKFi47yKpD9mY5TCCkcPnw1zp+R0w0VQG4s9iBRFMJ94ja
uRKaWZND9m/XaHReLtTz9J8kcOZempua/z+gaz8/4M7Dyz+cbhstHWoG5HAK
Suj4pOfDrzAzUknBSawUPkHQ1gqHOTR15/c4sXT/yufUWkuGAu2vpa2p0Owz
0JgTuFvYWkgcfxXeM7u1Os9QFuKBVfihaVGpmvMUOzYObFMJcibF5HAxcJJR
jzy7BhyOj7Yr1CvP9Is9pxSlC6CWIyGR30ytQb3sWMmEqAGd/cIWOwCzX5vy
dWWYrGRsXKPQDYdGyxFPFW+CyMlvSVNpdIcXwNPO88304/E/bvEZyTlAEjZC
fH8dQap+hs7FRGZpwmKIlqZbca5g+iCO9lUXWYZLMmB1n+DxfHTL+T9z8Czh
BuASq58j1lzIVWLy+lNoNq6nlufhIbyt4JZJcHg1tMqBjZ7I4LKpUr4ojONc
YN2m4EsbQ5/JICzA3BhircHhinueNkH5KMsCH20kL1tD6FsN2SXMOCstUUki
oKBtjshRbJPgZSawTVhewPUt6r/UQgfQzUDIvO5NvpeDi+88pmDjD+4PjqbL
vZF+nj8OQTNkxdJ7SuySXiOrr3G0BU6dYwV9IsFUM13bXosQhDbT+mPqga5K
d2wNUxCnZ0gfrzqTylAM8uXT6xzn6aHQEKSVT0T7hPivRQE5RNUyDv8GqiPb
gdh3lVGnG8zomqbU6TR8jadBpg2BKZpV9uGDUkww7ucvS1KItClZ/4+/qvtL
x+gJKnUVxqXg9+u/vxQFfejhN7NJZw6ziV/EICIbZk1i7X7Lo4A1UEyckqBb
PVQspoTgqG8MVSgaKot+zXEBg8WzhmKps7Q5fbbYC3E3110j15Krrhnxlsvv
J39tuCmRUdOSFibGLJWTkXV63CdH5BB5W52VPIldWqwrlh/p5nGZUSdV+Udc
s2D2spu9m/7xPyILS6mgZQlE2gmAkwev8V8EFvbSLoAgQokNlAf6oLWVV33b
3QgzwWsUZskP4Q10TgQGB3JMp9il2tAQNPZlcuANXqzLdY283Dl5UYureDLG
shawRGbf2OU9aWzmX8Giw2Ej3+gKha1a+Sdxxvh8tBSjS0hyaWdZolrLSz+q
fTzWyTWUqT6OHEx+UbzXhUz4oaWjeQqGRETpYM1AKW5lIXgOIjzs8d+3riyT
5iZAY/YASQQ18HMYA0322STCyRGumTF9xVldmh3dfQhTvBQaOBRVio6ovokD
XaxUnQ0KSVZUdSX9Kbu8XSRcE1bre6I7wEAqk4RQ4SgqzPMQzRP0uLktehB4
Fg5U5pRGzsHOqt+i3YEhpeeZory19GZHxyAWBKTO8Wc6K/cyOl7EY198igUw
Y0dUrRGXxpZHkeGB53mGSV0MACWKllJTcXZ7g0CsTHZyZQzqtiE5czOi9TpZ
ELjaNAQ+m95PInSsOFwn9mFBkK+IJrmEtg+KaeoIsamhT8qGfrSvoho1nSt5
oWQU1s34aamcdiiSqKJ7+nnqAXf5AWdftu7OiTT6CMGRD/01K2F4biTxQjxp
IDvPre8FjCmx4VQpDyu7woafJYNBNLsffNjHcAoZOl3kp7y8veQrH9KBof0m
St0ZUDcfkt9+aF8XFvaZE5oswb0hFsv1R3vEq954gQ71SbAgAQzq+iigSp7C
NuiXWw3zEdprof5wdEyeC2LqrnhAfbLarPFitt0186meoCDOT81um8M9N0Kk
GeY4xlP3ekEyJnDzLLCwBkuL8GnJp4m+/g7XPneOrKcpGmBeiRvNv5yzYOdm
6maWqq7UeG7tq3zKA8g/q7XXu9pNYB/HvE55dwyhJavijevhGUTvsM5ht6DD
bw7JwZrITKzxYeFbqYShiGeac5heS/uIa8fMUX1Z1qgC2MVi5l4Df60JvxtV
BeGC4KcT7vAiD39+A2elEVqSM1FTF4f2ieiS9jm1SUJbExfrHipLBszVpqTY
yMf6eIvis1/2O60hbDYpfUKsDG+pXHKf5v7iaKSguikf9Obk51jDGS8rR/qk
ARUzFUipGX92zYUfhUDaz+7Mt6Qz6sTP3ljeov8rByxInpQT1J/wctw+wRgU
5D+GHXODJkFy4gAlNmOYwoJR2MtkcdYQr1e1D38mw7zC3tG20VkxMJXVcy6t
rn+Hthw+m3JgN/N9pwgzL2pNxtRJ03oTdDr2Dms6S0aKzxx6pNYZAAvaPykn
MdUdCmnlJw7imdV/r33/CmlMdRCAaQDp4kqP3tl1W6bayE9z2kPA3cNbEajU
Ari7fVoSL8ddnEKTqmOXv0H+M9+nZwUiZoA1jjcWi5WtdXqy8QmfbtXVHEoe
FFBc6/XCiZ+lO+WPc1NF1aFSA6Mgyv2De/YQ61GF9lWYLS+bPmG96EE41QrA
+4k890v756zfm8Uv0oeQ4Hd0LspOr2P0Lef79k0s5wPe20g4QEj3plwo3mXO
+kQ7gZi0INYRstDVH2505g1WOY0adiG4iBR0NTkry7nb20lqSEADmYv2krXr
Xc4pImwAdBJHN5vfvmLP/2VBceVkcT66HBwlsWzJaL0fpJ67Yn8vGh+A3GAS
uF7m+ClfJfkzloD/RDFKWECl0y4ZufntAJVZjKXZDZlv1Rk3aNqe6Y43/DXX
DyZZPvS0ppweZywjSbY0c5uRLhFEF9kvpmme+L1bRghfjK3SAJF7DiYj4ZiV
C1TU71SL003SFPl4wRZAyJk5+Z0LObq5NquLc4pvE41KQ8r4G0a8uaS7CR61
LF5xgi4hj6n4ZYMRtgR7VinlzewzePf/bPbEin/AAQ8aJTI/LM4j4X3olX/z
kUfwFcSRxJTlvoAKWOULTnF9P8qdR4zVNffTnB4pp+1/lLcolqlqse87ekFc
TK08v7cYnCZot4iRVtRa6RgLTKahTqu1W93OtBYG47RyrvGSpTdvK3DdABM2
dcNJZ46PjAcpoRukfKY9Na+MbOiSj0A5Zirva2l1n3LlgTUqUg8Mat+9Er6U
GOwxqr8eOR+PDzD5sdKrrFteUn0t6QoBKlb4K8BZBArcM3vdQ6rdG6R8Jm7I
thFkiuYUdKUi/9JLUaJybf74jTrnDQiP0lexIANaBRdk1xBmp3M9YJRqkYPi
U+L8tT1LL+hzVygtBzDk0ZffdDqt3g3vw01oEeZI1dKG2VW+xr9V9Nyve2bH
da/+C/QHhaWUkg+lS8Ldeln2LP+oNW0ZDRRPdBEjC6mB/qcBFVArwEzrbAeA
Jv1dHZsKR8ptmhfpc8g6DfQJjeJxxtvzZkwb9GCJuzmdC3C0wrbpLBhyzfK0
AF8hFoqBXUE5Kwrl6b8CEBPRA3p2hU2FEac8qyVl98+F185WSxTVbk0/48fF
1TWPFYzHG0UrUiJvF7hxT1WWj6C6lj4WrbOjfXEToRckTXZNnV9YvTzpyzqS
QEkbGdiNokFxEYrGLNHszbxDzqUlvKaQzdja4taOAxr+/bTiRwJKBKISDNiz
Kso3bCUDmsYTTOXVgGMRvXg44viuLR/BoxXy74qv7K531g9C5l9t0jzgeNix
eR/ykeY+uarWX1NbOMRmK+UtZxf7S67UzSZV7IWlfgD734tbP8Kr3ZYhRTEY
8ZgB4r/CCRoLKUpWCBYB1XjuBXnkEeAvFV3kExmawACBzBNtam5+lIq3B8Cb
vqNaKKvKwN55GuMvXoePJ7hGzbZv7Yfkefb52YVLuWbVwNT9tPC9pLhoo60Z
1RgxH4JHeNzceVXrcYNyhcAockY5kOMhAfTu/7k1PKOumS1VfxytE8Nt0d5s
ETLvl9VKjhYAfcFY/FJxPzn17E1VlrjCxYj5KRNledXYothRtVn6Jh+W4E7E
zb7T/hRoY5Ar7DXSiFF1UokLhlXSViHqQlsPdRxaFzJsjqzXbhMxSgy2RE0D
KT3zq+cnq6tPZCoqm53VrP6CNi7NhkDrfgfwJvmD8VXqZUKomOLwkyiWkv8b
mSoQnYWgctdf7Ys4pABG3noBMBIYOYdP728MQwJjhOPn1LOE0yQlL8bmZBp2
9r4wrpIn59FTeEY2DRVDlS+n1JmRfLw6qcdE9uZCqFDFxDJn9Kkkuylk97Gm
+h/Nh0R4qp+FU6Vbm5Mov6O1flSgW3ApJBTHRlJHmWbDBedcKLTK8OWvSGrc
H8LSHFrm/F4HfC1/BJDs996K81+qTKWRcKZhACbMzPq9Z9U6eZpD9Ijpc1gT
egQhU7DFsZIDGQ6S4uWrdCLIXZkeHi2eWoheOS1J7GJ7WTvs3xq4Zd63F6Rj
Yq2LVvEjr+R2WyHac0gNQabub3pZvsXA3M5MUppcxkFhDGFt6JgMXOqqGfef
2ZqDCqUNqSpC4CiM79zGiLN+aPbPrQ3Lq5KWErrOEQIMIod0q5mtT4IGrHi/
yMsDPbChgOCPwcihjtBvY95vdnYaFBhLxtF7Ui8EG3NBnFqbuGkgaWOuXMXU
J1rK+JVala5BrRD8D05J5XFcNwmpm0tZAJ/dZWP9EDXI7dEKoyWG5zY1h/S8
5H4wnc2tZ4a8QPToNgeDmyazi8SsA5a+D9BsIAOL2priU01Ob4H/V76/u9GC
LGOTtklG4ROawHkVtM3vxsF0/HE88pnzILX7M7vniF4PrblyCjWEkp59bHjR
skcGjTeyeFOD3YTr0TmbV7jM6tO2npBxxn9SDcxWJ+dnU04PHK1wnQQtle3S
2mHLrV/P0pRWATTxht6jMfog2rfUNBoclFXvZf1owf0aLvfBLsTMqQ7G2fON
vscJjf9FSWZ4ijejAC0y2MTmgb1SsGaTVGOQrAXT1eO2M7K8T/gT8aG2RmcI
bx8cZVoLvFadXjfQkYtd4q5DzTI4wbUvvOZW+Dk0l8c7xkcVyWWsfjhdL4hr
jLGh3Mo9PQvsgCv3qV7FHWYeY3c82juIQJW+lWRC9w+kUntOzuGXoQB+A3c/
0/volA0aceiJ8hg8qXSLJe6V8N/ecH92FOpS1/tmiF1k7RQ8Akd3T4c1Dgmc
0Wit49BbvaK+3tF389c8dEaIQYY9CUuzDNrSDrDPKC4YpLG1s+NBuU2yWgXN
g+Ypf5BjsF+NEfrn9rRfnYAmFiYH6ey5v8/MMO+HZHlWGmwK6GeH2T4kOiii
+dZRRx+3XvQLWzs7NFKhtqOmyhJXi5u4jjlgilNlflo+oV9GFdahlg4feB0a
QOGlkf+cOuipK75hihEA54yZ6E5WsSMrUZskx1GKDEcRahnLZfqGEL1eOEbr
Xwq0xGqJfjZbzSFFl5Dq0yOS6JZRHl+FMGsTliX/I1mWpMsK0Ew9w6Wq3nQh
gJdsJ02cJShKN8CR7AgvIUrEtCY4R3n4wR0trlkMvyImjL3LzqWu39Afv1Yv
vOlQuGxeQFtIIbS6GKZRE5BuahqMfQqMR4lDrA1nABgYuZaqfWYXgcbkfaHk
sslVoZCVt2wU6VyfmWAHJBCuO9kMuggZIv7AwhYzKfjB+6A5Ta74R+Y1wnUn
pk2nPDyxcAVHLCQu4n2m2k9F2VvQShK2nt2iCz5C+cLAkj377Y6lzuRMRmgj
GXsvPxDkjHi4Z1jFkPgvUVvPafTwji7VZFNFYjBH2bOgqbtKA1sD9Zzaiwzk
YsdNpMZ9PCg5CefGROMhG0NaoZ+pDqmuYbSoOyrBfbFpc7CIqNWQDsqAVobq
Cfd8jhBGK6FtM2RQ/P2v+qgyeKjZHYf5I3nzkAlLeUL0HvH7YtheuG9yOhtf
IMGgIR1qY8K4JPbHoE0YJP9uGOlGX/whvi0/1iqbWmBQMcEfiku5mJ4awzpk
q1zjetp4c40C/dU4WryBr8ZaprQBM5Y+NqFMO/vDB8oEfeeqFAIK8y36QXK+
HYkEZNywzWa5V8yTX+Y9K0bVlJxa4ayMt1PiKq01JxxGmx1FEO2eXi6r6xXA
kewLIJasbZ2aUKeITs1QVMoIFi6pCpntDgWaBOZMzsCBoVMXGfsRnwc2xgyg
ekFOlCpIcqMBU2pzasIUW0wsp1a/h3dQndaRN7ZFOnfqFR5XtuXaIHkCPC70
VqpTKOXNMKnm4o6tSPiiIEX3xRxyky68e1vFwFg48yHhX5sIuqrls3fU7T0Q
j5UtEEnvtbqt4ouUQgMPZp72H2h7LysRPTySXZWULhQh163iWyiAeQy/Ng7U
bV7ohWLOCSzFoM1oZGa90PL5KV5/jgdr2Wrg2g6AY8moRa8S19W9Pq7R2gQF
hS+N2025jQBtBfG9NQhKAhpX0Gpnk3ke2kGQOhHQoLwCC8BLFIbysnYC35q9
BWrbKzoysaK+MRx4C9jdbOhpZn1BsNnpOwSoFcR6QKupdRRey4Yyqhi7Fbp1
hLel19Ib/dPoIwUs7fAbaoZWNXxPnw7gAQ4ov/eKE1yI19jNJ9mxqCBktlYH
Ng4JGuEeP7J1nl1K9AlctyKtRgzPzYN+9zCWMujt52feJDby8GBOQ8WWZt4k
caFTlC9Verqo+MsoVhBTRUlbF1VvH27mJD6lxfC/k/JZzZl412pZLC57xdje
ymdy71xx+hfTC2f2Gt3MLVjWOgfcNiLa8eOjetUUK1pUBhXPxg3hdYsmIH5v
2cpX1UJZSyCWEETN6nmyResulqEVawZHiR00EpGNUIhHr5aFZ8rbxDQ64mzj
sbTho4mPKn6VqhXufm34zfDSkUZCHV/XyA2eaJho4B3o0hsWPfyYaW8N3kdw
80+O5EUlAqNAuvB5J9BkbS/qrDJOA02o0szJzmy9GRCD0942NBhHkTF0olWT
7i+6pZ5FNkgnDh2KwP7ECRPsyYWGdKrgge0XevSKNNt4267a+RlIhov1rsdJ
EXkTADI4TZKpRJeQADpHOlW5YKlVpFBfxIwzWQVaxPBoXPgApgoXNKlnvWiZ
IZsSNCfdGwJ9dx4JfTXiqGygObUtdgdrp0q33QpAQ+OzTgrMGuPR+F0cWKTe
OcpbEHzaJrvA/GSBlr7pL+EsnfPHDg3acGKTZbw8bkOuc8e2NWaoCTq4fzv7
j6vNQZh+TtDFwXUcBih9G019W6NY6Lwg60IWV29vdDWAkYI33ShPcgQsQjmv
fQ3rU4oqBa5OGe2e/uJFPtPin1DqxkNC1G+8XXOXJU9M6goOvhcscqiCxa11
JAQ+JOVDYvIE3AomqPcckFKJPv0vxirTN0aTPb/uYuNNPFbp8INjxRbWtX2s
KgwuZ2xwXLEKBedvZUsN14pzBgfp+VfopvzezSFkinlhDsANkNyknOBspH8B
Wn7LOU06uu3TZ9Vn0+vCrNw54M9DvPZ/NbTt9Z/N9/4mqPE/wM9ULrBg6ber
NMjoShH4xceJC1tQLRgxwYTqtSuQ9RslFVEN5cCp1vMLDDrLPCZKdEYZrJzn
IhzQgfr4lPtcEsxpIIeju8Po5c+Qkd3+Vg416p5HZ5WTxuRBOvFnoKTE+66s
iTfnIMgjVliXpn2cKUEa0mbx0KoYjwFyXN5J88k0JnfdsgixdIjvTq+fTFA1
2w2I1eVjXfylA8+Hx1010ktqbzXgCwsdNlMH00rEic2dMtRz5a1hSCoKORFS
1uC3U+Cmatnz8VMCweV6ClnQlyvf2UyrjuGwpZf1rnhnZPZnlqN8R8PoCE5X
JbED5FcaZeZTlHB3Y5F0kBnk72sHlHtdQcDoQRovQWR0MXbNBPAHt+8eLal8
ro3S3paKi4Y19FVfCG44gXR8otQt+NAs6Hi8KBSa6gvrCgZULH08k5pPcfyK
X+6+i4lnyighdBAW9Ufv3YCWtg3lmq0Ae5DaGtffeMCFo2t4+yX47s0UYd+r
QFT126Yxo7WnBflnH9j2+bm3MtSg119LhKFrDFumzF3kAFRhiyTmuHaE96rW
8ilPO32e93gQZ+D4NM6YyoSBCjldQx5XxkSCc0gnxOnnWq6c3BtoHJNP/QOW
4/v9vNzH69KyrI9PiiYkVml2xX7GiV3dqPP3cqNQtNwtlQkVnMEvnmm7LgYK
gr1KaEMsmRDgklnEX0m+zCjBDKRBl1eFNVoheIhibgAN2Oz25H9gMA/tGWYc
uYhatLrtABULyt95/NotXAt2Kvtf3hxjbEGvuem9b3fkravK6VJeLeRjTFas
fgpU2w7AMx9BB3oUh/4wWuPXC4RntrG4CATH8GAt7MQilvDT3xV2waLzb5wD
dcywgX20UNzY6ocwJar5cCSnP7QIXAexir9ZGDnqCi5Fwnid6jkI5s//JVGx
InsgyPS//dLGG3M9keH+Xu+dhIJltYaYIhgaoeILn3ChK+ff10h16LLeallj
BUpAmixsBkx+GeGMk4KEzdLgPyaj1uCzQcnk/Ri5ENTmGIay1yJuH7s69fAC
noiQlKEKhGC1unaguRrVYNnHIaWafV8DlvyVI8SA2UP1Cg2pUpw1w1J55JTc
qdhrHFP5EgNaGXOQ6OMwW092Ks+zCPYm24fNEB0OmuyASDyfL1JYj19YStep
OvMSIWl5ppSDwBU9vMtn86lDK86DhwjDVYdJ+BAz3X4q7tFquD+TTLSCbE2u
sjggxLG3TtmafJDsPT5N53NXjvaWnV3m7V3MVHYChtQMSfUQUs3Sd7JtCSyq
+EnQTC6bqLiK0paswnaPfJtgj6tMH7kMb8M6MHZ+uQNDpqbDmWNmb0dLcMhI
MMUA21ww9JV7GDq7rIytQI9+vPfbTBrs9ruv67iUi906YlJrRrAtlDEsbD9d
hbzt9hGqpphsi2sjLM6lbqXehZi/wHfXdJzuhBJR6y9dHWGQNo/qxRpE/LY1
4aiIidTFQ6WvB+mE5uAn5rqBQgGlmYdcOdWXA0E2uhNmIMARCZtAOW5aR3s9
GBLKNFeC3Yy5HfsB+sNkbJQEXx16ne+zWX4hft0BXU4f7CMJEUmLX1jDbFog
C4LQfPDs6Uk7gJVfMJVjlLzeFfsuBv0m0KbVAY84xrB+7/DMODSPlx5lw+aM
+6GIm/FDINWE/LSKSGRWxbrc+t4Vy6MrfuzaT32hC2VMPS/5RoFaf1zB+xSV
zwZWXCNFLa4+oHfuiBtT0arQusfUjfaO29cPmG8Aua71n6fv32aU2ZBckMdb
WQcDV5JH3yIVbtpN9IJrCsEZNH7WHn8Rggu7Puf4W2b2NG1ZP8vExIPPoFP2
tFzlDGFq2fH77Kh9lI4JWtMKb3aktw5ZQQfygwoWJlnqm7s7OxpWkrBYRdyb
J03VBcn3Qz07RF7ujF6hXqwh0MJjdLsZs59vqiDiI2AHMzHBsKXfUZXm6GI2
fP7vCgxDKrpgc4rilGGZqFOfoStWvEFgeYuQvGVTdoWcCeNyInxDU70qmcu9
x3IeCPHEqraIeJXsZFKyMpENeeWny9s9HBpsIQMI3y5v6V+4tRpk+RBAE6/1
EkEXoPZ1Ceywgef1a92FapJAU9Ii/o32VsEzb40PVECX/GghOMgw4aQsI7Kv
Y00hC4AYgNw6673pp2WXcjKhkW4dfrliwwFt9y7s3x0aWHBt+4xmFpNkgfzn
wphk/B6o6QrC4EIbwMnOo2/E6x9Ff9VgdRinkgmxo0e9HkRW60u1Cvd6PM58
6ntgwVzgZfKqw1H/TsjW25H4aYB/s8bBZ6x3rItngMPwUERA636UQpHI0uFY
Xcz5fZsE7R8ifLBtH1FXmM4xGlUf+1TpNcHUDlf+SeRd/YwqnTf+VDLokY9u
wEfYwQ+G499iBxPOF1SrU1P4J8KePYIAKEfXMA97eVmxJvx7Zza3fo5Tp4zj
5N8XHmCNxpsFpw0Oz6rjyddXCtHh9hQyn7aJaIkjouqup6J+xd8G7/yqYOw1
FVXba656e91HXC2O4X7tgSug7C/HKgmo/Q+Opuec3d5bZCcUfazMkwDdEhjg
cdx8jgOWPhMH0U/jczOvNF7ROLqSiTzwCLjkw0jbjjA8bBhbGtg1X0QC+sRn
fZIWbQ5Y0zFzLCwG93FYNEji8k8vwMjg8T28SQqz67Z6zwagARjgFWIC5BC6
YeFbJrqSjesSvMLdL0Z5WjhftyRzKY9ZskGt5684NKpNW8TDTynGmCBiWjSw
eaBtmfjNW/tJ7qFCUDbyTFe8E57/R5lsIJyG24A/S5/hWaW8mVNaEoMOhRqg
GdMajyVFbZ9lGWYTi4Ygj5WHyJCtXi5MYMjkYDOtVhX7VyjVVCG6AtVacdk1
96PKfFSEJd9Sxtaq41jhltPci/wKgVp9T8h0R9TE9ishg4GX7EOKgThQ2ZyE
bl7MJkksZPfZxbunRN5SNNJphOik5n4/VZwzE8zbA6Ly6DzBVICcc51zd2Yb
BLOOmQlV7k69iUFWvlTksXOVZGRSjyHdlEeWh0mrpD1qTLznIl9pFLQq9xFy
SADuVInxk+joFO6rbGoSTKz2BLkUiR/kWatxJouQ+CJVKftHJsFpVfG9jmO+
oVlS7l35tA/xWLmxQHhMXWFaYEtowScf8jeUezXCBm51SdmecBGkh9i3nUgk
eF8qXgdPMlS0JTqw7ZOvscfGMTfiEPbXUYXa0uv+sdOFXJLtrKbQNrY1b+NU
Q+zYdNW1UPh01Ie7l5zS3ztqJMV7vAzsVL2lGfzd79J+ZyLap0n2GXaaYzb8
wIYeuRM8KMFE6S6pgBQU8msqjdb7qDwWUohNC0XhQDmgOi3ONBMCAQ4gCsBX
bJijk/T/jeItbM6YJqDJfOCtYxBs+GQwZJ7n75wInNp+xJjAznf0zR0xRP31
slfJkk7/mKinVala5YbMybL2cP03qcW8+ExyW0zJyxXImE0olkFB662kRmHD
2FUn3Np1XLH58iIavrZ4SRk1mvYGsFa4M6Ybtvk+eqoJCbAUru/cCsmAAw+u
orljyIr23DuwJwhcvQ/HHnBFSBJgiS5Xrw8Bz0zi71yTSuouYb38xnVR4RUi
YimBJ3rOOdwvUlrYYUmAyr5bDqt2PHEk0uzsswEUb3OVAZiOIj0i4Iy4uyDA
yfPZbqzVxOsEkY42MRbtWdrF5W28Jlp6T9CbluVNsxivijQFoR4+ZU4b7ksW
CV4pB1+dGzhnto2R1FeUJT3IhNioiqbX1v2vmIS2Pt2kDStOjS49/nXZEcwq
UxRx3kzc5r9jvpF6E/LCCgzIbnmbrzd/l8aTj3e73rC3HAnW5G8y/uH27SSL
IWHG+QuUMSaqgwHR0XXCOW4udD6nS3J1t2yNRYL0SIWs1UiHMxsMio2af5xA
ynGdmHbGpi/9KEhq3WFoy76F2vT2mus15YcDsjD/jmLFbyjxWqY7tgpHgAy2
CYYeKd1MvZ3VFFdNYkAk/B0MqmUg0Q/YQqEZ1e34ya20jaYWnoOf8JXWJpit
sQDooHoKx0WYhmH2HlUjMRE8VDwu31QwvSdefXVOP9PbdKlanIpEbg9Wk57z
KQnhEgWRiRC0D0WiVKjG96x0+XAxHI8PcUI4nXjUpeBcrdsizncZvcJS4qM7
Cu9xNMrE4w6/CeezdCK/BfqogUyhS6CBgnxF8wmymgi9DRSb1EtH7HtCVXqD
UK/Smsbvo0TuuSK9s9yLTYWeVNDAyY/CSDBLkV+zJFhRxpr9C17AFT6pKntu
0r9kb8aJO85cSWLGckDi252g28ECsnwGgExLmLJMvscccuNiS2/2/Z5g+H6F
gbIwwSd9ZzKWv++ePdilrUW2lspFIosNh2Ku8N+eSUUN1zmFtBEjvCL1jAz5
JiGCE5727hhvLrR5GspV6tfh7NK6rgfgx4LkyxnxW3AzI2oDZHfanB4NNJeC
Vkcf6wf10EMWmqs6JiiRaYB4ZL138zpbARGC1fa4ivtiZY8KWSdq8OFGW2uD
lTfMYBORmDELkGK5wO4CcS4DHS4DwQq29/7M2z1GX+Oiqh/HrjblirJD9N+X
SlAAUobCYXPRyzisf+NRJqUQvq2OVAyb1iVSwBZjQWtz/XZS4Fv4JoVIICUd
xd7iFEuTyoerZIfxtZB+T2u5RaOBI580XYL80p/WUivztdjKZGr67y3A56Ls
l9NJUHrH5p6cb2DqvrR1lwIapHc9JX1xWcOwumekrtamE1GMIkbTonYTKxMX
ltcktRV32KSFWWt1LOhjOoxAvXwTp7BNTesmiU89PCVZLvlOkXSXSf+snfsL
u7ndVSuqkkk+gcade7WQRD9eElyWC8Q/gj2jAnrVICyFdjl9i8L15Sw09han
afxKXi84SGFGGFQoqOWPYxI1TdrMTX7RNJHIicHhE4QYOFI1L5GleolzoD2z
suQVpfI1B8l1hUdmU/qm/LA2oL/QX7ZH/drnSzedt0Kvo/SCWdZXr8ZV/daN
LVtghF/8epDfFybQEOU3xvmWT8qth5iLk/LWWXyJxKNOfo3PjgZiUBFwFHrt
Z+8Dhpfh7bhvE8ebfYyyq/jb86B8PMQBfh67r94CbkXYlro250gqXOe/NVMz
K6rETIQJURCJ7ip75Dpkyq2juh4D3Kmn9rvPVoF/QquqzHahfIig+OypesYO
6DHoyqEtMk6ymlgfrf2bItGVq1pDhK0v94jI7qXOuUECMNeAVRk0+M0VKMYx
UhZLpl54phzuX//hbDH7B7d/fQkpHimS0BLbT+bcK5z/8c5mp+8c/WI2ApP6
tA4TDdwHN3VppZ2iE2VvQFbowcIWwLFjlAZIxjXaGiyBoODjcSsh9UMv5l6Y
u5wBqCB/nZA8REfKv++2ZhMvcbbQxH5FKeo2UBDId2HRY00A9nglEjEQP6+g
Gl1ya3jT8LpiSKtjQpijFFFGSe2eUmSTqdIGOF9/L0EtGKcygKyo5ntHdfY3
ZfjlqkETEz7V/t1xH+NQYBnKERBUIuSx+Q0Nm56rlZrGc2n0powbSNnjf7j5
DtFHOq6QxSy1lNHaJ9mB1vDcWj/CHl/FrcaW1v4J9gU4JBSqAgw7QvWmkOY0
w1n7qJKDZpA6xmrANFqeTgmQZhBe834XtUKMF+9yELDLwKweT1SIVSrVhtyg
1zdYrUNoWeTBbfUXIGKK3Tae/ORjkyw1v5xSh1k470VfiR9nDHUs+yoH1Nux
lsueZibAd4Y9xkP1RqF+8ZzvsMcxXGqg7DZV3YTftAGkMbzc8HtkLK2rWarE
mOkTnjlo0YqFsiyLklqMR8H6s5Lyes+6heLNI5huwmGidODUWsUwuRO86hmJ
BJqAMpE3yA5TbIGw4/e3M8fKk9abo2NHwSVYFnrV62V6/kEU+YwKSqcMAHrW
Kp4bNa0d7jLBYBQFm5KW8g/z6HIb1+uQjpmySFXATDpeiUuT0rRk4n1/5+gN
9i1f/XvI1jpATsfzzC/QqZc5UOpTmfUIEi2sy9Dg2jY5iFV+7U2tKAT/sX3u
V07q4pIuVhNoI4Uq2vO2litmcScGUk+sXAdF5PPckWPTxSCdUWoHE7UvNBYO
u+mADmi01GubHlbT/+OPvQdygGSulaGKPI/o7ADRtlIZd8yaZWVcMVsS49xd
fWbpMqOJf3T3abEnYAwpHDQ5Pffp4391inarGXib/QpJcHeCyLWBIZ2diW91
d2KtT3WdWdtnPFtHIqOyScKAJVTCh8YQSl0fxucLqlMCciU+IERQWbMkDTDU
PB1FFfffdF5v1YCYpfL02Mn31IncLW8/2Ina/ERp9U661/GYX+DLtCZp5blJ
ldeklu3XmxaDC5CVu0IpEh3YA08rACXtk6aJ5OBzxir6bd0f6eIESTMHStFT
oaQvCAXroN0jBJXrNa9cWcJ+2RygmmjlavgPdYSwD4tQaNHjKaZAZI7b06Ft
6d32RDMprRc5l98oEmlUPjzISdwiKIQ+5ItgownOym62aWuZG328jAZMK+fO
mZExlkjwD1pBO3VAmlQGqa4ZCwBg1njA10pYcok+kDUtytLQ0trYij0134mt
jSusiCStRT8T/km8arNNA2TGm6ZmWwmm3HlBue0SW3AK3qQo44Jg9L0T4FGA
OVrp/dYOCjAtreZ7wGZeiqS2EWm8eZdclT+8Uy9V3JEZxGViSeF684iaQCDa
WQRtnMz5YmseoxuGRe0XkM6ACgiQbuLWZcutf1AKV0rVFiK6qujwU9TZflJe
BQ2KLEUf435IpYe3MeM8LHBJ/P/Nz3dq3Z4et8iKWXqug9hnu9vci/ToJItZ
Jpi8hC+q0rJszKAgD+e3fbrSzDJjCc95X596mSLjVU8x+VhwgAc8l0C73cEV
48wfiVZOR4h17H8cnL1emX1w9ZJI8Q4mxMxV0FPjIbHdIQBVDbYvfjeeKLGo
IoghtHsNahWrDKH4nFJJfZydCKAcDJrtwOtwexxw7fyb3+oADt3jajp/ZaTU
l9+U31pvOjNMFTrUsOh4r3WLpN+/QJkK8C+P1EmbNn84m5IQP7VG/9Im6k3D
a4YQ7wt1lsi/oyDQINe1/ktVFHkHt0GjExgmoW3yUsxHzR6wMlDTPtJQLWHd
yb6lnumDqv+dS+Uwvj+T8iYz92R6g3i5/jbnuZ+KTOKj+aMlU8pdNCfL3NcK
t0OgpiG3I4C7YQRyYvRKlK2CmAde3M9rRRSzEEZDFwCXExm7ToFoCHKekneN
bITTh9+6K9Im24jtD8wVhf3KPSLcqqmi4ksnHpisAHEeZfcYYuy7Q4slA32J
LNYd1drGzFGBjcyUocT8b7gAXDsLt5pSNA5Y5FcHfmzVChwmTxVjbwqeknLJ
9OZu0UluKEW301hLW1QSmGp6Q41hnV3ILVy1DdHSvNE9gthJ7stBVdrFW1Nl
05eE6otbgG2VDWePpztvP4EaoNjw86cF02e0sqdGnGbJx5RnljVgbpSQidMa
bU7sBy1+n2AtrORpL4WDP3Lc3xUIQEmWOAq5Dr7YVhIsDqeYZ+KzZclo5xqT
dtAWKQjOPfCXylIyLH+nZyvOFZO/w36eTQolPW5dv9vcRkFZLGi6bXACPh3X
SrWi08Mp7o5luG8X4FafANCHiu/Mo9kZTcweUfXWIePSuoUfRWMzZF3BwIWg
C09BuC9rrG7z9uekFYUn0LJrutSj9pykvO9dWqTcODbqfj6tw88lwLAXvkI7
3nFd/HVAzQmm34TfrXS3j8ytSzP03iA1QjFrvMzmqU2kUJfEvQVQguWWnKym
fsjfCDYCGjVRkf/6nOhvmNsIG68+JwE/xUPm3VFgFTG2lK+VKyTkGzcpe9sJ
ZiAVGLZy3xdNaxzZKdYo1BjtWff+brwzZWsYQP6uuaKfK2HiSc2MIVWVwpzD
5ofSHVtfckZyMgB+9qCL0aNafE5AhGdRhdHoNMAoRYTL9KhOjWCzLsh0ODpC
PeMvL1b5W1NtEBg+iDVLhzhMw/TIqBjxfnGy4xECvOIZeiN1Lb40za3k+9NG
Xctru1u9UMZmnn2Y9uARX6eKR5cSnUWs232koRmdlR3rEw+0IfZ3Ah/USN12
lmgn5d7Du+PIosafzmzTi9LPxiB2MjWdTCIXGsew6oFq9lL40xl6/oiCq43B
PxolAkNqlHTWByKjQ3yQUhqKiwCOU0lgLEfH23pq/jnDHsZhUQ/8MvNiVyNS
wcYG7qQYj9Chx1wMS+SRtBy3EZzVoCdN+C882NoraBH3ca58mouwperXMaYz
1JMLbBokKjeOkpZejcVICnMVYh0MD/gjZXcO+1SjJvjEX1wQ9B2TipeHSUQ5
oYAmI+EPeLhCnYtTN5oQYCRIH4zK+Mygji8vmYouVC4+k0uggj4IQjh/PrkF
snOOcwluBge1RbteYgU/ZQMZvhh1WVG3WcVgCgSHHWq6D2fQTO2yP4BJC9sK
Uq2YZy21+ISKTBSrbZUxkpn8u2kvRAZ/MgN6TJ/9Q6sCF9TmSsnHUqJngOqj
qCeEVbfeOwMlYLTF/1TPPWpYkubgj632mq4lq7M1i5rrYxO/9HGJLFIkDwif
gq6JYcTnbkX9if9BXwH/tOmHglrlQciSWqeYBagGvigfrkad8eZgSiTsNhb3
yX5btJsAcSAQybY4luq6pCMEFcGMvdW7cxBBFG/+gSVCWZo1IqqF6wiDJxvD
k/KjlW08Y3FZ3yL7doJ4csu4svQU3QlbLvUEx6f1clsQ4VxBrfAIEccwwJQX
cUmsbRmOOJXfJYDjm1mRSip/3GSnKnqPP7WGh4FA4U4oNvVZSdu0zKdcOWC2
yvB/q+2W6tlHBRyoQxMBqOKxYh2fNxzmaOR7YbWnG3pBgYRTJ/urrXOXWxJ4
lyShxjqRvZmNr8Cgd3OnhRVamslYx+hJ1ABI7PX/K9/SsI1b8AlceXwrnYSz
YUwEyyK4haj6neNXNvq5z1QVDT2sRQa79xcMlFVVXDxBcz3hEF8j44DK1Dqb
8/Pr1IlZfwekVoHB8wsbncxZHUxLdd9Lp61qO2YvtVraYdTdEQJKpR4BGDku
R7bPxAfzdPCMtvh6CjWCJArh5+hy5yXIH0aIqy7942YAA82oRxT7B1jbKd+S
8+mgrIc9Ir3YN/z3uL4GbDgZzkSSnAozVopmxF25B4Ga1w/RUNiOhIGnrboX
uM0zk8k4zem/77/sY3drlSWzX2cMAkfDtw+1q1QcZu5KnuX0gjk0/acS28x9
8TW7FPxWdrp4HW3F+Ibz+62IxFWsVtuRgZyWqTRLP6I6q7ntQvBKk5wjKmPQ
/cVzJw/WBsQsPCK8cYNbwr2Za3beAWpc5X8nKIJ+siSALoyzrEJTHBFRA7Ij
R/hqFbsHYoWF58D6O+6K/8NUtUarUQ6Ydh+iw+HWztUVQo0IfYwOTlytx+Db
iesrloCnvm2BRMzZrLbRuCaJ7CBLgTnyiNqvFAl4srTbOIgwPrFQMlDqnYTN
xFL8ohZzI3azvLKCz/7heC74p15RGGpOEDsxCM9hKC2CyUuibtzYjl1L7TO0
gELSL9NZi2jyDrRcpQ2MwbkMeNYf2SrbI8zhVRoHCFMY2nVOMheUY12iLXUn
4DyjlcD+U6QlRSR3OHzf+vwIHCHKpf7z462uUk/VrC6DueeYhnhSWPTFwcym
dNFvyHDmBvTDrWk6qiVm8jVBEMKRcz6xi4DtoNEwQAQjQGgQKcy9p4zwWNee
2BNp3Jg7TOpLu9Zdp33Luh0sWllmEhE+/bPKnlGsrNHl3xa8SvW5X7MSy0tC
hiy1/JWby52NnSKkv43VRWIrtXWJRCdTKMOYDz/8hzkiBmbYmUJ7BpM7tbx9
m5ts/2TzSONrjZIJMcC64a27yzQFjKSKTfK/7hoezDu9UJpDyKBH18de+ZSz
BVmE4WWIdWtUGvoZeL/oscTBbFcHoLVvwPwG8NoZ8Q4P9UX0q6f/mU8lNYBa
5SI+pRq3+8z2BN91lnLI2y5cCfGqSLwq/n7LZtsIpxLu8dOzGV+pAduhyr8t
lCzH8n17273a3hZ0tVYyA3oAm32T/bPI+lIoBB4WDNRPNuGBqhIDj9tKh6bW
v2HQzxNwupGPGx9sH94dRqRsqZFkGfDYTRy/2Qtd9R57W1FfLRWhaG25uCNF
bSpaR2wZvrj/psHL58E5MfkoYqcUkgschMFuan36RdkHUkP9ZnL3vhiRJXGv
C4axFbLvME6VQMmEPftgRNUe1eM0pQw05cH5/bpYMj+fyr5504cLNGleUUO+
YynmiKt/+SGaupqtzmBRCcNv34R73kHzpdf9sohKTtwbkYclUmb9yVFp14PU
WZXGVy8b5ZI+fsNExQqYDvcw8eRMsvJDkdgz5D8VDSq2HdaaH1TXAB3CVNlL
hQcst5+upZjTje3Jths8mj3HG1HusOeNGyTrkOSguVA4m6l8+a6C6IK6pE9r
P9/ZbAnmzefH61d41mUi521GRvvYiOO+KWUVLUSOKSQP/P7p515/BRMgYyq+
UqSa64j+mXX9vVo+1ivNwP4AF6U0Yn4KU1M3UvXLSUgSTjonK9bv8EwdXg6a
+00T/c0ByMECYCfVMfNC1aM+G8pyi5zcDaqfpmSLJqW490FbqSmMFff7P7eA
Ma5IocWkmxoMLIH/cDaib+o5AoWXKP4sqn5O5sQDFTaziL9yjBuq48pwgIs2
uKDeSq9g0OqV97wyaODtDWE2xzQ/Lqu6Ih5OhI0jRqlfz34gwcpOY14I4+9v
jUTIc/ksk3PYYvQ23AcbwsUoeO5ArdhapOdul8FqKUfIRGYiV1yJU25aS9Yb
UO2xvJpH9kCtAjRqerZCBJSR82yxH4I9RtOoGuOKzsWWnKgfR3ZzlmPR/hkH
tmVRt7v+4dTJXTJxTPvXTfxpIIAKc/9TTjy+J1wVa+k/Ezm1FBsg1Yn1BmTZ
HlIauSszDOiIX4KyfMBdOfhAj3AdtmNe6Owc0NueNdkw2SfV6XlQZrl2S3ON
UF4D7i0Ni1nDIPqLvMKa99tud+InuUJPwBIhuOIX6/pFn4VC8uhdEhwBAcoP
+qPNnslZMyrt68GWz+WM6I7k+bZvGA3phc4Yx6/BZK295nuaGuqHzZ81AODI
BUgJUdd9/2bqFI8jot6g2IopJf9x7lRV2jqxY5OyWKao4GPF2KQQjA3ycw4/
PWxvWMpTiX8EDZ+jel5OV0RBh41SG5+jObXQU6hyenaRcWaa8SJPNPBhJDHf
rlIX/d65ZmO/OrIn6EecnA6LBALau52BlayFFJP5HV8VhtP4zz2ayt93w4hT
rBNd9dWeJ9lJFJWqjqMXCGivHOmc7EjK+JxgPN+BI+zCiIBCSvEww+xc0NCi
T9f09mpCAjIbTbYD7kcx9Ej02I+Jbh/vQbPJM6AngRVH97tvVK5tOxBEUYJq
wiWto4f9nrL1v+wgO6c5/NUDrN2F3AfVa1kHzPHDC55yoplpJjufZ13N1+SS
LhYF0+7uv22dsoFx2VB1lihsJ8t38wc3nvfQK8bDfCWkzZF34J56DlSMiPZX
n2HcZDBCGHNSGcHYqtBADMR5qabKv6/c8nghGZOuR5kUO15GV/Xpb6HgAgJ7
tCSupEexQcdXUrcbsDrCV8/0Varo9JUYeUtH9k705R9ePrLogzJSRgp/e/XM
tBWQe8kkF/WUB/W4SpU/qlwZT+fDt5hqESbQAb5+DJVpa3vtdv1bf/kGgpg5
eJRlpyp9uYLfZWATcgvpeZ5aacUiGWSkAqBh6uTEM61qP1C201JitWsWuiwO
N+7ieCv3bOFO3Sa2xZCe8de1sZdQzd0X633pgRsl+6sJklb/MdUPst56El3C
zxxory27IvoHuHr4sBFBQOb7+Gj5gYYmsloUPB39GYHet3lWQbXY6J/ioi+g
O4cPVEm96WHiJocMOk6/eT2IKRmLqa0Zuoy1XkCyFYoeK9h/IHSqor6GfEPo
T4uOA9PjGlzsHOaRT5QE/3OCdsGJjVwr3xVZ9NDHB2UfyI0zLVDB7+gbcUo2
HNgwnnQQcmHNV2gMM6XP8m1CkOMi9CAVo0ilBiGgbvAhk9xo274K13tYsSfE
t3p1MAGOQXWUe/RVAgtsG5S7kWA50McZd+0MTP/7pa1XTHGFLDyUiWDykW6a
8UlmbyPP4Qa9FsD+DeYgcy1Hzj9o/71mqkldjMJnHbpbgVyhws+9+XPTTgSI
Xf3Pc7XhcmjDUWvJ6pYHQfTTmLjH2mN2RCTrKICVl3dTst3gGklSyiM803tG
fkSqpsbuWtwnUH6HmEPGZll0bnfSUHNAnkT2YrzoJ26ucR2aANoswy08k90B
SqD+KHKtgD7di/Fu3jFIzNqtiyU4eKjq/JfZBNj1VZYsT2F3LMZcwp/Z4ENr
4B/2FIuXfKFMt10j0YMbh4o2Zn6AHF8Ik+FPFCwFXDUqRHzG9RDh/sVNJfv4
3ixUb86SxbZ67qa+BVXSvxusTrKZEiz6Mvb0WPJlrwgFd85jXkpNHAGFwo+b
gm+ETBtVTQkrRr74f6b6dee6XlNB6wFgcI59/3mLg7qrQvLJusXnd1pGC3l2
fi7Ys+K5W3KqdedvzIENuz7W2TLGcSg3AVSpQPY5POPyvaUbpL8eVjU0UBqz
8XKPmTsy/f4oBO95mAhUXBa2Y2c8SGugKUMwtd1SLY5eFmiN4/6Tt+vpwLvZ
D5aDQXhjVoTmr0U7KqkKucLEPdsHMzK1mQpxusWoxCXwQ9Sf1nidh0hGRf54
0T5+lt0x0ikJcPVzUbag4vFo1VjqR7nh9WxNZWbmsgKRynH6IyB2y5SjWqHd
S+MIQGLR2+VXruWGl1RNXE8REJw3fR6FCvXEBucO7ln+3biKDi5pLy92U/Rd
XLtCnKxsL2QfHXRvp/pLYq+fwY3gjlV8k3pnErOZ8RV5j1rWVG9OuAEwyMbo
TjfHQuKZj/uS2pizZ4779eSm9P4RN47mbw+30LYyupPDhOeA/5MWCHKTbTkL
mEB+vmx4RLvcZ6v7sk7gYQionOJKt28gqhhMpnGPT81grOwH+vHY9AY2vMQG
Hl6aHS6EeGudBTpITmwDmXZSU7aV3gaZVSC9AXcBdx9PWK7pdn8YbF/AhFv9
+T0OXGD6MwUomSEi/yVcHzCkAfNLyOSWL8gmdVKYgyPX6CkDsh63LFH64x4d
+D4xZPdiGzuazjwxAa9Myw/pxIV0dwffzHhxqJ+VKyfUHcXTey6XEMRSbKPC
kDCX3hQmGoaC8zkdbS9dsAN/gabTMw0gJ2CqCXCg4ckWD9CPTCGi88NwSjWC
CCOHjzNEIiEIPNlTnJeWeYBUKCeq4KD87M8ghB6795zEGSfN1mu/uAlgWGOW
waemBsWRV1KhxgV5eNqKWs2Kgsmm15plla9lZiQfiSlM61/L/GxRdRP82da+
oknD1r3e4u7BBoongWEY+X+hVeHaGZ97MUSiFRnAm1Bp2Fahgbub9WJ/rpW8
uQEyBPrfA8Tz+tZMe81PICMtwOiLlF6XH1wfsl6IyC6khBGUJTbwsIzR2eeo
VuF6KIdgJD1NhNobuYV7uBzyN5i5U8wicr9goIMwrrxsoScKVOaLV7opwbO9
ZJYQnxikPk8fjak6s49va/9cDWGBGmqXfONR1Vv4p3Id0ACz27z3G7hz0l4r
c26PewQ6fLmFGNs/mx+N8HzcuGci4AUKq923xcazsMtKIqd2ImIL5aKkcKQW
1JXBEJMe36C+WCVJBcuodyWN0f6fdi3FlFuQSlgapUezv0M9ALp9+ksnNQZw
v6LFKoF8xndje2JYPh4m10hsOOG/u8YTjg4h/p1OGWWNl7KfY1cqCg/IkA5K
M1ruxS/1AJpEw2D4uO6OC8YrFPw9sODTYEcx1dJvPW3HJfVE71ytZAeLMXqf
aQnn6u36SFzHgFRyVWYkKnjcWt5zihUWxlj8x5RTfPrUoD8IgSRHyqipKkx8
DSwRWM27VB6cQXIn+n9n7djFbXAt7cp1UHyWfPZ53YS3TV58630oBtdUqK50
MMFwL8YlF45jP6B220IZOnTkZLRbnQCwkUwJc570QyxkPVReFJr4v7PLIXTR
ARoPkvJ8ELAsYc/Ir9bDkLyqLVLzNeq8H7CMbBVCDQB7WlkRVg7mCABm4QSd
0pJTCAKQeDiiVwYvEzKtVwVoBDbYjo+YY7UCe3/ccWP6MpAZv7xG7DdwOT/V
N5vsg5JG4x8M1q/OBSsj/qL3ecx4J9NvZkzToB8DSWPX+cK6UsEVCK7EeuvF
zeDFSKqDWX6hOYcUIuCRbEEIEmfmO72IU2lMlKujMLN28h4nldspyWWTmE50
BPJRT7uLhjOFomoDztM09TnZk3T6qdKsx48MaZbyCUgbtAYHjDXMOZ4WjjBP
hNn35lHwIckgmauu2n9eLFIEyoWU9ogXisjBFccDbVK+n+3Sj0dU3J9J6YuF
j2n4zhUYUKKBzM6OMRw6Zj/njN+pkqX8bcYjP23kx6/qRAyIjHM9ldFZgkBI
ZUQysSzXvNLg8C3Pl1bUIhRUF6jRiq0sOmbQ8O/kACRyRtCgySD9KkoQmDqU
ecTfHM0=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "221cqLfSQtZLwpVKjUxAj0azxWo9qWyTHel1yyBq9riDaTa7pjyEaEdGOLLz3wcrK5rHulca0g1g9Zlx/VJp3su79bVOdFJFOSZrof0/9wf6C4nAWrw+2PgJSzMMKpaFLO6gpDFruW5083aTh1M+Q5KnW16yLzHWGhpxtWHi5x5kzslfPRMwe4HyZUYh8/FwJanr1Um2jvkSaUjUKvojtHUTdbUpkWg93bqHvMIamsnkPTRFPpNCN4ocODv71U0D9o3pueeT+zRqXeH3te/7GS7ilzqzj9m73ibrVLaKXlAXqxcRaUBgjaQeBDpW9hO1Qm25tSpE6JkKVAUn/7PAWB2GIijhsGjKmnr1f+9e4cuKTEGiEY2l9T/Y9WB9cMSFh9hUV+bmfFcfKw2VjaP+omHgQV5zYZMuzlSgib5Ljj54542rSAytK8b0VlCoPvuFRCb0JnqEBCnztpDYlCgbN70AwrMyPL5jGJYwfUwikQFEqaD0NOuEy+zaATWUCclL/2osikp4g27RorrLOjy7bR++4o0Tis6JZhfttviWGKiE8pRgjYUD+1L9TCHIyOJjsN803/VERnKQV8n3VqUHczkKk05hyWk4Jf0TKjaDzXSlIG4JFR2CMunA1qBFAoEsHRSs54XkKjrTyM7khszJ9h59Iligekjk5y0NILtcqlOPXt2+ujkyrv30/5wgYbbhgBJzRYQbWCVcGiGKbJ0rp65A0A3zSxHXOFmGBLk4e1Lwk/6f6dHyHagqzxnPhFh8JHkJP3EImMFaGoOY89QZN0wZd6w2NmAps/K1yh+dGcnW5Dt1iAoETBbDiBK3S1KjJzjhxB1U/Vvl2RvWkILPR977RONu0qCaZydX0XSPuWvexAP2COMnHkNkzetxr5iJMKAVKqbAhmBqF7qvuP/In/7e/GVh40CzBarGHQWMUsIJItI049WGumLM+M0DeAzd2AAJay4bBqXZ8ddukw+AoZA2QJ5kCiGls5nzyWeFpVTuS+K7MOLhEV3nq40gBRCz"
`endif